`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hulrRGewxnypy36JMhQkyhJciTgTDxDanilvdgXP3o3OpxwVDHlc9J5R4gBNsyMQ
Z0659MtfMSqD4xQmtsfzA3vE98QORtH2VqgDvzV2duqlxBRjh8P+aBm99snvkdMe
yfVcc+xDOgnUXtMNSQkSm7PqetTH3ENVLk7DEtNH+mEa8b5efyQdut+EisM3PDNT
cZGhgCbibuysfYTMPXFtsqmQSAC3zWspYZMYmcpbA6H3Lnfz142TRLwIG+gs1959
lK9i2EtvlPZx3d3dibWTVIsaDyBVhbOpWH3krAB9sBE=
`protect END_PROTECTED
