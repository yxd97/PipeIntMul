`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yANuRcPBq2C7vc+WmhjyH/5nolMjymrg47S4ovp2KDFB2msEcWQykuQ4Rp06AYaC
gWLtu8v40ab5BjmKkK/HHGaKJH78aOsXjGAUT+UE++7AIFaBNjkcnT4YDlKLcoAK
iyHjrY1CqgPkpNCfqFJyXG+FNMk3bO1iFVEKIEv8pS1U2zP3bcA/Q/V+w5pJuMQ4
4cKAtOA3zioACiTLciwEKoZGMDsUegfyw0PLmAdMSo9qRJ2wKoOpzBnQCKV12UIq
O3EN4IUPCfHtbzlKq9yIavhmZDqOBcKYIFQqJrca66ljBKUxEWv3sJxODW/X5knB
RnleNGzjiGMmkleA5dnm+JeqcQ2jKoEs8fYNs76y9mTW2/e/vOg0umcBt044f/Cv
OpBQ7FWq41XB/ng1hGZVdQvjjkSW2enH1RF9G/ywxVzJAdSmf64OfXDpHDQGwBQn
9TgIQDwSswNtRhfzu3xAWQ==
`protect END_PROTECTED
