`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2d7+DNSEL9UGK3hlxqrJOiwkHpOA7nmqouAbFhYgHKTRnctxBXDUN7SEzSgEOhBX
qXqkD0t7OJ2GA8VVw+Mx9nVX4KEOn4jcEmvWknkpRT7Q4yNtgN7+a97PWRuErvbh
sYkag8+Fnx5QhmP4mN+api7Tyq0GTfTw16uhe+fW7/VdBpfWa8DjyO5HOKMNFEVF
3oHO1+m9zkPPumVanCMOkK9KmKFnn6N+QSKMJVOOrfJj49IgHHa/GYGiPSMvqSgM
D58LXfg8nIwuDOJhC4hra8P351vvZQAr0BgcQkT3kR1u0cJWWHhSeT2ccM2VArVc
3h3P5DN95VTbQ2dxNqFd/kyfOoSu4AoU5D8dq9/HqOT3THd18+rmQdOQYYx/nlXY
33Ll3AwWAFddmi4voHuWHZk4Fh8mDVpZWnAyh6sKtchqHnUkDSD096heg3oMG4/M
+0xiv377uok5a9s0qGYGMew5Alk1BIApZPlrpXe+m1nNVKxD1f+iZhCj2yFKshKv
LAV96oP+86OpAR/uY7rc0PVGUASpqKzZjzuBfFvEE1tXIWz+GrdJsD/ZtYB2vnB6
6tLUCadh4NbIIZR0zlEUMjqMuKKy6Zg2xu3gcgYuR3YeFyYV6dYPl+6wonXNrEW8
vwM+oFcEk4BH78bZg4z39hly86E2a9VIY92rjeVmHVdLyyu3yHntg6qRhfOxj6xh
2XPY2bO9sGNv6wDWvVPYEPC5HFrYeYYMWWC9pcVq4dhacJgKY3YPeqA62bOF0gBM
aPw/szJoS3fdSuLcLow3j0LIDqxFM1fha1R/hhSJdIKvLybjEJdTiw/Vs5JtqeRW
jjsRM77vXqoDzyz9QrncxLAZ01vTx4Jtp2gtMa/wxoM1yDmC+2CIHgdTDyaXMe3A
I92QoMIIk/BgaQwpVkoPgdXQPq45sjpuMEy0hx/A19kX5orpw4lB9G7cgryoWyvy
XfKpdkpPFNVFV9X9u6kf/rcw2soA3or+g57givdPueBRmzca/WFk4t0zrR90pbgP
XHRMA4fsxXW2tX1LConpZ9uLrsiwT1Ys/avadFZyyjPboraYvVZQDSXBj/zScPTY
WxyrDNocgHfylGFORk3h0YZmDwkEV0882NMSmEpw6fkpS5YUEMIM7l8GemWeig8J
2qLizhdxDmrR5zjXR4r8JxFceKqLRFlhFxRatPp9kRBoC9yd6ll85IjTZrJDt8uo
eEATozuoPz9YOj/6+u1KqAqBsSWFfvAjl+8wm0W9vwbPuufze0PCwCQTFbdBj6u4
Zgk2rNMOFIObxDuqttrT2EHMTef95BXolg5isM1qTXKe+3SfhkC3PKqjrxgpelO8
nrbsKuontE2LjdLP9F5sy557MBy/U3UCY1L00cOjIgBR6Pb0HS+Js0yE+9EZUluN
JK7A0Sr7u5PJ8qBZoHmGt8QDmw4xKalK6Lwhah85eN3qSQodSf+B2ZK+I3a/wrlF
bSWXpFeSzeGh7mFMk3s685xqxv4eHN4N5ePShi4uVXHT62ji3K7aG4pFgycWKvM2
yiIPy5SIFyftHMJVmJ5d0e50o6wj+oj3n6lliLPAz6rTIti3sP2/8dZnh+oCydlt
/lVrdeMHlFfGzq6Jg1uZTRSnGmawSGTSIuIcMYojxhkyd5Xxzq4SFgio/gWXeFqc
IuO9xNq16OliUksG3j+MmRYzFZjdA8KJ4M3Uxee+TwRy1yI0+x2Mbwdry9ETrpnM
hbRf7Tzvv9QBXNKB2+cy7NINkOhNHYWQDW+0oGQw3/24cgwrn18kcc26N1EIr277
BTvuqKilMSDM1u9ZN07c9lQ0/uNfrqirEfzPnM6kNkTHGi2FSXqSkRTsaEqegqbE
Q/ImzI5Kc0p82NCYz7rDqQbhy38CSkfVZGvw/o2plz0=
`protect END_PROTECTED
