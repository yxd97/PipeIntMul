`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BA3WInsjq253RlJ+egIHRjGRyapANwaQq/SIRfil7Q9hEUeMH4lLwDEZJWpPhAK4
y3qhWLEV3tMnr5/dD2i0Uy71Tjt1OEyqx1RgQvIIZj8ZemmE5ENOmsZT2M/FYOlw
H+3ZNoSeIKDvNaKgPGMsbeIq1KIOjF8rjPeLnM7zuW4sI1ydieo0JQRCBP41H0Ij
vRGkctlV9ZTfjZmkV02v6TMMfhgIpFoyCBapPShMV+eMNiCDJ2XlwdD4Nc016O/C
VKesOyyE/Cgz2QbhUM7GbNqd+PLlGn46u3SVsNj4NK0xTlR3xUmU72To1NCh1fT6
EfYUlBqv+/QWOHE5eLY2ziVjqNVwg1cLzriy5S9HhBAME7crCX4awB5h4ouCs/gi
ioMNm1h2k8x8jLzJWq0bYWoizyFVLYXpxOUp0mMgu0PvdLZ6JEZ3c1ZVCyq/I8/V
CVcF5snM3cdEckZQcpF+M2mUY5RuFAoVGWIL17aIR/ywXhIRwtWSXFYV1wjdlprw
Wzzp/ikcZ+8tQGN2RL/OFi9v8/IWCxKtoi4m1Ns2XaOhMwqBwXyOY64Kp2pRcui0
KvK1zd9MqDDMw4t98BALlVGqQAnZzzm/+G0aNb3wwmbqwUs7xp0NCK66S7/sakoJ
9/F4Tb1cNTsga6/L3R0oQ4uPw2COAmu/qfyfcnomu1vdHFTgcRKie0WZaXADQmMm
Fn8BE/Y0YD1oF9t5IW5CmSsH1ttZhyRSHc1J8sggoprporQ9cAbsYR1b9GzI2c8C
tmj9b630YzeY53OjHwQCmxJ4TejrOXSvKxsBaWjTlGCGjWU6kzTO/1vMQV6vofVp
shMgpwqdLNhR2AHe5JHHtH0YFEjmLgRY0GCQDKwkwkqQkUmOu6ZhbIUiKd0VR7Wi
B/61fCC+LqzUANVCHAxXnDvuduDzWn36DaU3HjufbUHdL+WCKcPTWSrJ6j6PYwsL
2xDYXbPdD1ml73XdFpPcjxfJb8ukSGBnzZFeIW1UoS1OdAkBug4reAE6LB1lRtfd
A90zNZqs2vkJ8xBV85y9SwYJAgqi/JXoM/kFNlq8mGc7FQrYXHeI2O0YzsJWCDTH
X6Ziv0AII2Yz91Idc8MvIsPbfrUKvvL5jKKBpU1sdcI7nRwDZ0UJNt2AMmEkj0W3
sISNWaL6HzaAz7qQNY7Db71nV8AYZRCzgunPEdh52U4CRL5AZCXjGqNfbFOogo58
BDW2fKMapWIHbYrJT3ZzDYl5NAFl3x86vPugBzcRpEqZ0i14Xcf+cSWC5wg1gs7g
VACxCM4TjLe5o38aVN/YqhKJIJrqvvHeh80ibjcYYKG2esZJzW75m3pWIVoiH9u3
1p+UU0uPLxPREoz1N2UB86juK0ZQtizIPvjRSehsPcGqj3riRmLPuqqsRftaUKjg
ERB5ieObQgLKM7c/YfLOEG0EVpF90+bbTN0oc5cUeiHe+pOqVwLATOhv4rSQY4vJ
7vxEIMh9NrefahVN+UWJujBFikE+Szbbc5H0UDdgqKl2Z8T+HDEzrVY6UyR+U9Z9
kHPyaiibOzH/Q3dSP9yFq5FFYrN0LROMd0jBYunIN7kpfMSFZxRy4tG/mBoIrnz9
5HPQR1z7DsBz1DPtLkNM4EVdpuiwRPdYKKV+Ygky4vY1uLM31zg8MNB0YYapwhEw
+hWhTCN6FT7kxH9uDdeSBCyd3HRve+p3hRnL/slUJAooXgAG8s5IpXEO76L+sm+Z
rozsJNC4MIf8V4CfDD15W6udQ7AItlLFwfzYyasWxaBLeSqt1J4PTPQDiN+7Q6Gg
eOZhNSRmcyz4aTTd1o0NeTZPMestEeNvH+pYMFhXFpPNc6dMY1E+tDa/PAh5pNOj
HnypXERqBknaKkqxrsMLALG7eDC0ubFwPof9TX91Mw0bfCu3jau9bU0owTOGAenQ
`protect END_PROTECTED
