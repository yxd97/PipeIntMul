`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkMlWJP8YbCMmrWjU76nN+5nDCXcA1AEeUkMqOFN3Gy+HxVaB9UczGUl3rxE3TpI
KAWDqP6+Gc9ThLW/KatV19Un92OEy4eWsOSpo/anE6YdHOePpQNTKxtIea8rctGM
G372h4JphjjPklN1l1zycbJcZ0o92db4P9SaNu+xYhtwE2+qB9WqifW6L5go5sMe
a+MTe0g46M+Cysh1MmVjQSa6c4hEdaS1a7L1QKg3ZPm022N7CqbnXGbwTpbp/u4u
snMVsRoVAcL/U4B5bxN4X44qnPHQwgK1y0nIv/CXbOOk/zXVF2ujShrH86w7Eyrt
VrOqQKGWvUZLpOMHL0I62NB5bKmUX0TkF1zZY0reDLvwSg8LSBXPXhW35ho9avvC
nH/1TsISI/4y1bgsUCmiAWEgXOWQA8dSJQLvgar0vlWwEDUzSakpxLdFtfdzMxtS
mjlrZ/Q3GUwzR0MMHOBuyrMpIgEHqEkE8QfuRKJ/QlSYNKo0XrCIlfUPHk7Y3Qxj
Q8eLKDvgSd75V3lqocyJ6xXC0lAZ/X6vBVzvHgAlcr8ubpOE//4a+ixEisbwxhKP
+AAYlVFTzF4ElzbtfN2HuDQ/KqJUil+ORFRlLsXdFdM=
`protect END_PROTECTED
