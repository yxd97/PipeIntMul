`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bv4NF31dM0iOxcMWoC0eyk6peuSRQZgwmQFKHwgc0KwEYwptGHO6v2Frz7bEjx/
wFsGabNqwmrfe+ABsJKHcgYg7Wi0mN8zoMTL2mH0910mGOs8Bd2aZKf/K0zI7MKq
jPh4fO8V4xPdFCV6ylc3O0TdMXHYbzIdUi+rdvTvUtsuz8a4wh6cbUWQO42QAm0x
6MW2rJf7LZgSJf1vjbb5Gt3LXQHI+QrblsUGQJEudCxp7XT5VCZoBm1/wW/GH4iE
Gs1ZQCp1Vyo+IFyvm625USZlDSbbnJsxVSrtLPHN5yVEZS9ywFSaIOzQgu4JD7TT
5EhOc4UUFZ7UYX6I0ZWctrwWTMYxB43GS3TmuFtskxwQR5FSJuKN13gAChQeaAaa
DAnl5h252Z49MBJGNlmA5r+oya/wZx9xR2a8t3sgpB2kw/owRmGPjiGshIr778aa
W2I5QMSZ4JnDNZOi0niexkjEoes5oWMX9VoN1vAPO8pTVh6roIrqy4PHopv0DiNS
pIuTOVbctiZusGf1NhiZDKM9VgTcw+x5i2snWIidf7BocH6hvqVAvYFf6wuuj7fO
IpsOUcVRWnvcciUrFI5+4SS0GTciQV0auFrD1NdlnfWTQxJbJt+8SUI4rXPSy9k7
G66oN5ea61vCHuiB5hE6aX8rkbpJhRXWzmUzZyIpDp4kby7l99qxMuFmKPaV3x2p
QrvP0tODNUZn6/syHIiZBFWoBowep+IzcC/NLtA+5h2LrKnGMK8BEgfkW4LJDVuZ
8YugdYKjXEouM2ltMPXuetEKL7oaWpo8bMKDfdQNL9HDBQ4KoHHPgs3TfIabwgp6
lwkQutusx0eRH1MunROQsK9wBAR+hLa5JxZiTt6KJG0nvvcLM2j0CrRDMiqZVgm7
F76DUPwbaO4u55/KWFvqEMEU74guGBYG94sQmjoZQH6bBTOnQ2j/6DRD8kS5NIAG
Z91BzI2uaiiwEFLl9pLeGoqfkhR0nWWM8XURkyq9FOs=
`protect END_PROTECTED
