`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3t7ONW8LKwa0yrz1QUa6Ntn1foJAfqD2er9JzLVS4SCnGtwiJOJqQUN+kBLgeQ8B
WeJYycF+8zYXOBwD6ay3mcU5XHPBAGlrlduZnxQN+xJOO8V8fAu7DR72ZwHTVefm
M07EZ0Pvv2PHHjT41QzSEzIOTgIn9XZwMfQ3Pr3qEH8sWtOkN5qHx++0Mwitcgk0
kRZmOtoX3+/6SRp40TdIKDDkv3mPm1OoT5eydGUiam8UUNMTK1s7xM02L0EtbYwX
Ngc0KkRXhaCtp1JQVscq3NrxEWVjydecn2bCBM7uRiTkxmpZY6EQVz3c8/hQ+AAE
DkRxq3XVaSFm2dX7Kl6b96YL5rWpwG98DtQ5TNlvxRmRua7Fb9s3pqJu+shwLJ7g
sF7kIMPt1f4H0vB2/2pHs2xPLx8vPN3yUlN224oF63dgrXsEdvFsaf72hgrSeJRQ
2VoiG8EbGCJlWzzCuy+NlKThKvs+kBMhQGiBhm511F/L8VRGjoTOp6qnsmsUMOIR
94tqXf5W9CVoPRY//Rt8KfKDyPllqlD5OZfhadRc3c0=
`protect END_PROTECTED
