`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAUQLKLSzBNTZHCnhBV56ZJwKvgyuEELapKxrAFlPPpZ5YYiB+4Lv8o24+Yk1pFe
kvNZRcQSFRM/mWmvnGR4zRdtDKtIomlyjQjngWicnBxNvsiKYt9CU55FhRl6RUch
o5KyyOnZnBu2bZErP1pxRdfkrHcERC0taK31dg5hptCwoushRdfrprFCu1LFGVnT
mK9m21aNoRA6PxVl+HdO+5hMx9QQ+IrU3eMHAquQ6W2SxsAJHhM7xRM8IYz0Q41H
jXzVbeMW5nyjf4ofVXU7mq8zcZ83IZU3opUZF26T1T2QRS/+riyHQJZnzh4lVznY
45+ZtsaPpQXTRBdNOoYlzWhSfc8Zee3j4qcVhe114NI2DiaWVihPGHlsxsba7Nms
PxduHRAhB0GnazrrlTUW9TModWNMQ7fSczV4Rw9o8d/Inu2K+By+oJboxDztEc30
cVfWQmFaHDMygdKuSN1vQO4J4TEG39F6Uz+MWp9cmRJz5N3NfY3/8TUVUectESKN
`protect END_PROTECTED
