`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YDoYh+ygg/SPIrxv+P1Dt3wQPXG0H9YBWpnzpk1tGpJyOyNPUMSTeimTPBZfxLI4
LYXaGrbxsRpuon4astpTn5Ay0DpfimBRV+AEAiMAkVl7OJRVH2tNaV/8SrIp1Io4
x0Wyra+V3tkRXzfD8EEM0CcUBGB0jaj1LfU9XbhSZ/0tsQI1/qXG8zvA327BGO1I
HElk3PC/ZwJnAy9uX/rnrp/kqnXMmMlYC6wl8rNiKyWxpElrwgmBYrEt3plB3GHG
DUcs44SKITfmXasOXYAsN3dDbNnhmGk1GpZh3hjptXnbWueReSqehc661yep49B9
NbzqpxxaYaqSIcBTWuYbhRddngRjTBLyAn6CgfQHuNl1r7ThQia62mBGaRxWfxb4
EKKR+/RLzWabhTtfBAhoj1KDnAYexQ+7U6TwMTX7F8nGMIoK2PG1umfYfbCSgVhU
sCifj9Tj2FmQMZvMF/M7b8Sn+BxGMjcc0hcOST+xmIs4B5XFiD1DZ9DOuwKg0mLJ
8pQDbhCG0y5VRNHdxXIUBBDzGiiBwY7EnsIAnYqGhhRW88uSfElXurcaWEkwfPNO
5AVil1TA+mVUQxJnOwHUI4kX+ZQtpSeLAGkajtkoWlhRp/+Oo3DMGy3Kj+Kr8T3a
nteTCP0l7TvhQSFXTLpeQC+1d7WGSP5MOgdlfGan/8aZFuERuS2I/G3o+N8aYSOP
HWzcEhXuX6CCk0F9RhQaIt0o7FIbOFy2dKcYFbYM4+djdPUop+7ObRR/1TzfR6wb
y3BsZYkGDzn5dBF2ZGD1rY5iyP2l8+cutEmpk2jBiGfB1fANplsTaDDCOJpx3HFs
`protect END_PROTECTED
