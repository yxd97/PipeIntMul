`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IskeaA7YtnraX/NY9Y5+NUow0wxmFGaRFo1oU21eFbc8WiDD5UYZf3zzPm5T9Yl6
98FZ2tOGp//RLWzEm8jTeyQlilDokXKIBKDGAdWQwzTXXM8akBFciZdqDfYlV68+
aOuK6UIHeuFhwKT1h7pMC7necREQgFl+SFyHtvu7y3FEWk16b/py9HkLBddxTFrN
xeNvl8NfhVZv92+AT9/FAJu/mf/xPLrpQ2ACCyvrMTSqyQtQ+pBKUd7Kh/fF7xxL
pbt4zokDXWDwZEfntgjuoQ==
`protect END_PROTECTED
