`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2l2APuXHoov75tAZju9DAXRzF7oSgrGhhbwmJ1037pVMsyG6A0OXt0nX2R1MQmc
QAv87H1n8sXcQlsM8ViZzSHGbUsmrW+nwEWmr6w8riTitTYB2dE3f80PO2dOtVCM
nFYzTgr8Xew7p7Hx+SXw4OsEXW4OKWSFKOXIcqd6ChymLDVK1aIQS2oToBQcqk+T
U59BleSKvNVrIf9mfzwbER96uxdg1485aNhiabWGRmKp8Dr2KRinkOWsd72W+uuk
xQle8gZVmVSLUZBKfbsGH3DaEU6vWHfsVynb8oLdF3PtWejYVeoym3To1BVROrpT
UU/wA8jJSnLCCQbbeF9+ub7BMvfglZ8R9kKT8w2SpiER1klVGroO9vLaxzIG+5hS
MKH2UY52gIApXcbRIosHRPh+LPNXRWTwdHSyKHlhbXnXqXWTJYvTuLHCcCF7XCjE
6NzDJ5AKtaJVz7yWnsidQWsdVofcZ7dxwUA9GTn3dL6DBHRWPip+DZsY+M2q20dD
XfFFA+GLkSpJaHZBik7l4EAlRuHyqUaBP/demOpMAoePmdm9eL/0P9pkeIOKNM2B
ZDUUR/E6hMmYpj1d1W+v8wG67dGs+IFw/68Y8njvGdzVUVZI2mjnHeiHDYoeRiTn
fCnJx7Hm5QEPwMXuERV+D+SZ9ILTp6yvMHx4jhBW9s7bP5Q73jcIYtHpM+/+V/A2
ws8ZuglZcLTto8dWCMrOuH2DZ9NxuTrICkPYZf5A8c3spsPXqA+mQgkDpGyDxESX
A3aNCVdH75TDfdCkJoMaX2i5VEH04DM94x3EEgJE7UUWU6Zr226X+XEOyg9k9tpL
3WvWLTkOxObkyEjl4NzerE80XIQKKo1XYayNqY9Qbw1EUZcDbzQ8pEc0PHPybNWu
iVWGD32NaPiwa+/rWdfd7CIa5zYsR6zKI76hN0VFwaxfUPrhXuLhQYFq4oKSVaOq
tyLQ6xlg3Tp2WOqx4R7W0f8l3Y+l5KEiapXhbsB929tjOit3a5Ta6C0+N7Pa1P1v
oelzFbrOOmt+K6x2Ng2PQuGQuI8muxt0VdJ8AnbICn9PjhdoL/BmayGwm+JNIv7C
Utsrri26XNKgJsO+dp5PGL3HSEc/4tS/DFpy1I5VnrwJqjGOv9Wo6ueCf9qN9ajT
/2+shRJ65Xca2cx9Z1WdjxT0gbRdRIX6ICEfWAK+wK5iBvTNsZ0go0VXWi76hY2R
8VngCLCpQ005NYfqHptmdP8UNNzcGmu+jwQlphRiJ30C2T0JFogevV8WoWsUDEJ5
coQQMWggu3IXeV6dcqaLr+vcOCGuS80Z5JOdirOCb/yMB3vmotvigoSAzKpLtYbQ
IDpWX7tSUGLA+FheV8IkBKMItStnWXTJ4QBUYDHMLiKM5RE9jHpMxn3At3V6U84S
Q07bGNGHuZBgqvMyqPmOjLgbL2L4VQWn+/YB4632KxKGk+3p2FClRuf+aZerJSot
q2uWTEEqv3vbbPUN05goz0klvnuGKYLs+So9SHAf+ZVSuCD6dUhgPtK5KD4ye4Bd
YyZal3dMO425oXLnHSUUfIAE51ikcJyk8dcC3Q59Pd0=
`protect END_PROTECTED
