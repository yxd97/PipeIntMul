`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T/L11Q+PDBAzpyoR8UKGZSyGcn+aOmVCF+ihzFC7RP94L1Pf9pNg2+5TiD9FEufl
6Rc/0ZpKnMfJwix5FYj6IMe2tABA1sPlXWEKmpqyS+ABcLfAenTOGIGehXMcM5cQ
8WqJf2WDmO/OytAvlVFc8019DokkpNT9STo/5EeqjJt8xXixrVQp+khHkBWZAMMO
ngxwHMc2xPVoNpRaZ9s10wV3Tm5QO1zqkKOFWdD5JDtgszPF35p4712y3NNmIHij
oMy7b14g+5Hh3xnVbCtRosVJmPOH4LScbp2WB9ngdHm7DTBUVkmObkM0YuTTFf5r
RUXGt1EapwkuQJvhfPgUgGkDrK3S0sgHDe2mXv1bXcxmZ2sVnJgvJZQyFmya1djZ
AEsnFNTqaUDoKi2lX3pQIsn3ogXEUzgQSqmrciq9Qck=
`protect END_PROTECTED
