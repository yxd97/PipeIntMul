`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CyfeJcdtOT+IbAl9OmY1bT3JDw4YaJiKDe7jEY/upbM03iGWkdbLffgVCYzcj8Hl
bJtp/PMvTKEhxInNQBj3nA4RUXIf6EjrqIoLWD4p9Nf2as4uQqNwyh5JSZTQk899
0FICyG+G6JZ9fAeVKbqKXPxm0mLktGP1i8OVzGW0yozyoJAjCtextE8vNHydYNmP
tSzVZY16DKj5IslN52DkKKT6R4xNuWC2ZRS+LCIR053TPO8lR9ydMol/LrSftytg
C2hxD1EXqtWuyGKw62edI5VXrN/jFdqwk12MgbmJFF7kzCm99hUF0HQ8ybcrwfhu
yMq4M6HM4i1X/AI4TMvyVatiIvOkKCDXE3BFK/5oVlS7Pt8QoofpFw/sRXxbtCWS
s9ecNX5lpS57Nx/mKgY6zGNE5X7hXS2VI0zAfaUfg3l78IjvU0S1WB/Os3oFzjnU
oHlNVf93F1I5+ju3/C4TAdPhLAlc9PTUN2mYqZFy6ZqDpjUn9hXPufgygczQ7eqL
723emFKEodFi3OyC2A+rZD33U/bYMVmiah+IE1lbHs06yGHzIHeTXNTxcTCXs02c
t19c8e3/EpaVStlLiyTWw8APPDSfQ7TONXd/f+sEkTIfdpo2gP6GNdjBTxYL2Lbe
XR0dtKPOSLQCDeQ2zxQACmR6zSnAU4VXbw1P4H4dL6K5DjLUMJlALcgHf63oz3fL
ZwFsiGlZKT3w8c+SSZSErdkhWqy21ctzfaf+rEncnbJDLlPqMaGVBWs6yhEqixWA
`protect END_PROTECTED
