`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXlmmPKZvCC5bnpGFrqlZQQlUCnliw1/7VzBohtQM8VY/3z7WvCincbQhvGiCauX
PAtvVJexF+kautASy7lG1HuEEd10g+ywJ/saXTqsV6vYKx1CzYsdAhOTrjDzhW7S
JW0ipHGikYbMsKGeK/kVlZSGBjbNvKXQRnAGZl1a0rK6lSNq/Qaoejm20m/zdhxD
amf5NiorKsBZkHODT23xVuNRvKTXqb6uipZy9rhQXEaZJ9aLUf8F4U48KvHTLpkz
fynUbKGZi1Ct0n272NMWZ28vRuQklOk6AmZCGy0y546DJY6jphF6QH7GFvxXL77h
UHPJTKIqDFzg+dquKCv+cvi9BcmLHhPt40EEI+ZMAjPTK8ula0BD887KUX1zcDUN
GMcMnhHgK8h1OA6sE5VsSg==
`protect END_PROTECTED
