`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UxvOZlbCaBsZPNpAAMnYG9PSjr4z5QRcUoBGYJHQlZdUJGeBuTQC2LgtPo6/ilpB
CZk+oZHGR2p0UxcFJ4lVDQ/yvOs2yi4FWBhUJ/NSeDSd3Jc7xsmsPGdcKk1p2nG6
aORqhGlAVmjkQ2cbI+SJr5yOewhZHKMhGKNJJ0AFxptVDlTw9qjuoQibib6jZxXM
g+Or9CjQyPwTQwyo8zzoaHatXvAy4v/CIPf6e9HVem2zOKyLr2k/J/iVCEfROMYT
Iqu6QWGeqKM7Yy1zi+f5CUnkbIMKlvFLYNCPMU4rbRD0CB7n8MVWrguVxsltfelm
19JZ2cEACSHWGpCI08dvuWO9z9imPpbY0iONP4t7DBXYuDOEhONRRZXBA+D1FmV9
Mbj5RXK+WBdUixwf+BY2VYSKo9y+N0TZ1HY4JMSlHTzLKjMdx1GE0aFtZoGyZa9L
RBk+INnpDBFhWcMLh6YYzq42y+eNFUGvEX0QUfLGHAiVq8lqOsKjdwIiC+1hxWS+
MaJdY/daauEHmsKM/8tk37xtEhwXvdJqu0gXU9QGD1pHwWjRCBJygCCF3AfqMlGX
Huwvn+s/tSjsI27RzUeARCXVKfEGqbhFRzQyyvVofcTkkiRZYxk1SZKAeDqNsxxU
TqtI63VtIgKTfOUuiriXPbvbSgO//4Jjy08hFS8nPl47fzJL70tdafEK7nO8d/kI
+xHGlf2iqlWCuZupZ2qbmSp26KaqIuHpaKNeo7dYoUkMhf35t79/7vafxXblUIKI
OU85ZXGG0ugztqBKV7KDC+be6qJOwomOFx3OB/UcQMMnKlQ+3m2i59ndqF1NWm0B
oIK6QWn3cGlqRalVbD9YGa0+PummfrxpPRb1hl+YfRGvZ3pV5iE/jdCHCxih3bf0
Oo30uKBvxdBsjqegORXP4k5isfr72/9WRvDMhfBB+L6Hi2GS4xm9c6vARfszQUxA
oS03VvQk4ie6WlmKjX8Vbb52H+cTON8rrGOk4GXQO7RDNqufsIP4T4dDG7NAya1+
I14+HhHeGetc4hyBY6MFfg==
`protect END_PROTECTED
