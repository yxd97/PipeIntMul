`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qiE9W+Tck+Sb6BE2p77xQzRlFnGelXNTexjw4/ivX0RtV0q5JhQhW0WR4S6JGkC2
4jzna/ua3d0cM6ephYcC0appGvdaLHx1YVCDWHStUgkD1X14u8BgbNADp7o4QlMq
P9BmjuCUepNo8uWwX6Kz3s5nP/kOrdU3XW7FuBRS1SkTr6w+7odmTie22yjAZwb3
eSB31fnvhKrpwrgA+oH0ZogdVoqF9ZZvaM8Aje1APCmZE1/PaYB10yweWH6BPvaC
GEd7AUqafeBim929USg8TYuuUo5ilwhYVRTiOOvmmDHx6TGaQuLOvHymzUVU0W32
4bNdCxpYBh90T2gUgZWVcCa6MwbKReiv7LNrCjdqpFxRvkvcl94nfdcv5p90ueom
w6yflffA27maV4AOckZnJdqfLWuqH7DG7T54PZ555YAbetMEKv9Xx65g6SAzmYsT
tzOoBlK0HChWIq7UR72a3qJaybjZEB4pVAId8xRsdx0=
`protect END_PROTECTED
