`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ui651JZGnIUoKUUzADRPT1h4M2JE5bqh8VKcL/3ESMyuYhX+kuC3G4Skuf9Qwui
f+gJGHikl1onlx/ksTM61/+4+HJKfEoicPZbVe95bM3+I10NusCMczyQ0Mcxznwk
oiQpP4+6ZcMDTEgAxJ9upNzPxF8Li95OTR8FK8FSsNBULhrh06R19ByH4YkIG1pr
qCGoXC8hzJ70Bpk7s2fznBupLe+0FlH9QfXjuNtaBJctXv64dPQ//7Vorcod9ua9
3d6M/KlKzjs6wFAHKw7eDLNg2mUqCoCAKdfxa9Kox8fzsm97FQZZSbmr8GMqT+iz
/fIVIMOHPnl3gNqyOihWMZHlzQ2gEsTcjZiBmFDhUFGJN+iFZoUoIdYlOv9buZav
JB5czGwWQmfZSlvK3DrXZg==
`protect END_PROTECTED
