`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXhUO3XoxVzu5Clg5B3d2Ylnc6AXN3jILqeCcg+0vfwljWmM2yqD+rB0oY6X85ki
oDzBq9ByisJ6dF6dBAGROWeKWgwe5tOOzvlAmOzAzyJ6VJMjSq8Mv//jj+hYT2Dz
dIACb8Fv4sEcnarTwn8LhUCkUhVMOrvCRSuuPAHJIFsy/p8qFJ38DtYC1bCjJE0B
OaAw5bVbGVP6wdJcRMhSHCulUsaMSaf/EO/KU+Hst6aJ/FE1NWs521+A0OSXDaK0
BOJMjo4R+Ayrq6a/pXhAAtsMEzCQ4WqiLsY5SRCufKqToSmK4YJqAopP6iag3ZV/
YqR1dWdYeLZ2fgVJiGNL7kNYI7vJLRtwKwXRvkJac3aUAWwNlpsly1EaIsVbYU3t
zIaIPHkcMVRby8mHPTBjVD2dYentwUobVfz8P7jDBp0=
`protect END_PROTECTED
