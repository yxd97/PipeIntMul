`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WrHZ61jPOT2Y1dgJoESToODMIssLdVYSRfHcHdeHNd9Zw8/9KRyXfa3vqP4lluOQ
FDMdba/Wuub2Wu+nnxZ+k7ECwhqGutaSOm9Y/JDtl25pf7wzMMK66khDwiSTtzy0
tL596sLBtrFoNZytx1iV8KcCGK8GgC56stVctr213+/wjI0gA6HCNH55zkqqQZ7H
K5CgyO3+sRH/r+MhRqElUlJhoSUWYy12DPXuBfKVk4fNcLOpEPRIxPlQgLuvEEfx
AzJAeHzxd6rQ5aepr6LKBH8adCUbggh2ir2T/XAVPHAJ5VAztdytw9kkEUTmFyvT
3Ebv2DjNXYVgAxIt0VgdxhQXtJBUcFmNz0WxKqfgIt+LoUqaxFUlJOOyBHXS7jIy
`protect END_PROTECTED
