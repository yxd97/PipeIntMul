`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ELH7Vc7io7fLcQQ16J2nNi6oMR52x3DzQSkl3i68DCarAn4TcCqdUsgGEpDQ9gB
5VEd8amiiXiwBVwL3jUkR0s04J8eUAr0BsykdVIVKqSEcZrdeTlj4FNrWPLEkAoT
zuhrb5mcGkqvjto4ICFYZVU969XwRDOSpqq/BcDNGYpFDP6AJYHbiOeFzrn2GbjC
/JV1/Ov12ydIjHtvKI5CL+Y8QIwk3gBkdrKvb3aeGp2Qwg12TYH+eTU1Q94E7/bT
se8jh+BYbr7QIP9LVbkGk/+A9m9H5quTIrzZnaE7vWss6sbiUwwhU8rTQ1i/hdLb
tnyM3G237EUkrQV+Mv01/sTd6Kh1Xj5mQvuEVqd8tItjZSyeCTO7s1NizxNbpb0r
J7TUwN+7P/GtA5Rza23WB3Mbu6Fl5YI2yYlRvb/MhHmNOA8JJlSwz5I9vEuEI1kE
wkbJh5GAKCFC/Nx/NBnU/FYIyhsFPesgz9r3Qdm/l62Kn8reOgFU5rYSZ5NwOSlL
ntahBBRipoZ0YX6hhaW90nHY5DZqjWuJuim68Qa5Ii1yzlQh/S2Gs9/ZJ8KARlTU
OaUH2YW7D8leYYsG3MWi7+/SfcA+1uOY6gY6qWmod+xx+36N+SMaqNKfrXptJ2xA
mNB94J5+QqFHl98zXW0Tu7ig/E3YIVIFi5Ls8+RGofDilGDVjrufU/i6Z8I9TplH
MFjfOI6UZDN/xJ4CQyjRI4xR+nSjHkvRVkQtL0txRI9IVVgE4pbLST55j9eezDgZ
IGfj8aTDfiguUBnD83QZy6H2+Tt2gsFp9QLDOwqqp4dXIO0KxV4X21kFj890k9uh
0ecmqTHxtqAiecoGpo0Z49XubSmIPs5hAcBfHRDfQcUpHII260L6k0XoAXfCJc1z
ywHhTNt7KN+Oh/1j1SEYm7sSINFTVasCYtiSdRMvymka4Vx1hRAbLLsXU7B4JAW9
lU7M1r1nV5Z1hK1qcHKyxk397C+L5UoxdUE34yeF8Nk8xMyjr9FDH3UPd8R7RaD7
`protect END_PROTECTED
