`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F8OHwDweFr0wwFdIbpWxYTsKe39/3qkR9WyBdxWkGe/QJ0wHK/uQbO5kTDEnPvPU
aG7YFe+FbXNOb7QMDAH1oHeoazKx+VkEe2KlcI6UoAz4SIR4ay7FQ7VjLCiUs6hd
bB0QHsC1yH7rQhbOshpNNBI4nY8fGAHnCce1QNM6t2Dm45DsNFhh9QR+ZNoCd4Zu
BoEwphuaHn/q4mWh+Ac4g6fa6WBzf+qiAAV2RiEW0HswdHr1btcRfrNdcNWNVaVt
SlN5vkfykXYVCjSxLSqwJE/mIhBAaayvzOsJXRw45Jk=
`protect END_PROTECTED
