`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pY5oq4ZpWbRMiIY2GLCu1ldw+izwkeVfRIZOZ80RmRUhEKcBSlk/rSOM/DDPnUWn
GL9mVpmBedIDKg29IRnVdt9d9FEfwfTRMgPqbn5EwAgCPAz6dxqJ9BiqASBKdVH1
Xb4Wb0fc5np9NwtJl6DXWJIB69RDfSQ4T4IEBq+U+3g0YmbirX4DbKICn6qDa6Wb
csaP3Fm8tuv0w0rl+72P69vOFURb3PcoLHwm/jtp7ebrDup6Ozv+ttV1ycjweGjW
HWcaummTMjkmGwdtYE7isk8nrKkMoTVqBkTJk/KtLeWjnaUusrsaCoITMpB0i2gz
nzLLdH4v+oTF7NeuCO0Gi9Fas+W92jBq98/U5rO00qqPnVWSUC4jZdog/XZAMPwK
Vfi/xGBZPH5HtNmmxuYra9D4SKjYxJqHRIoIVEgokfku8hpi9Vi4NXPh+FrWBFgV
aPT30FrS1HRhK11O+Vd5WIdjaS/amSQ/OLUpMEM0Pg9tXxL26KDf7Mu/GTzkKQs0
`protect END_PROTECTED
