`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wRAj02dOnTVKEIq1uAvrEYI/jzpHDtysV6Ejk72WtcrbzKT3t0cn7A3hJTsViir
pSdobB1j7XwU8vI+Q8aBFw81N8klv2MvSQwVgcz+ooOsaMcWhtZuXm51rME00GiT
y1L2s+wdNQ4+JvxvsgiLc5oGlRKcPCz1VVotvBqOxpO5ieZu8M8H/NQMbnTeJf+M
wQB8mBZZWThUcJbYSH25k0EwLVaCzKB6PsWSwXnXVBHknkWiZNyi2xp9s6Gn2Q13
l9O6LwuXhmoCZdAYLrJprfYDB2p7Sds3+Xr+ZObiNtBL9w1GZu/L8LY+6+CiAlaN
fcFhtojTx1K/XqOuc9pZvm5rZJKAyWAwfXeUnfPEx5P3j1IJojG0518dnlqYlx3R
`protect END_PROTECTED
