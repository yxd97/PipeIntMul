`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OdtR8hDEiFs9d9ipPrY4EFXBGdkJn980hbrkTg0tzfyyUX7ZcbnWZ5xBAtsWJ5V9
UhVL/pt7Js/Vf9ZE3yTgac6cmH+knpQnosY5XWl/HjT3ZqMMWDueg+Nv1ZnGSVzF
eqwO/th3B3MNL6twMXrwimF+cGT8ZFvfGvsMEzpJWEQEkPteFFTpvBs/8e5u6o4d
dE4YODz0uCZQXpTNGzFoGnI/C4TLZ6bDNbuftggSSNa64Iyl39ri5V+OUzgtIBWU
92P0P97X3Hbr8b+lCb5wv2qFBwAD9SbklBGTABAvIBo7jtkp37yqdjEyCgPyew9P
xHU2fGVNgrRpyeRI4dwRXSKMy7EtPRUQWQpBYWjThDQsB3xu0qpNcM78LlL8Snc6
XQ1K4PjZGjEJiUrcAwWwZ12TqmF2Ze+CbkmwGoXr80HWPmQnLEbGf/UdiCVHJdrn
OVeUgav5JXTjCo2FvreMoBwhFLgix/kUMt58YSDuSr38nQmZlpQZSB3lIfLPp4WH
DYfdylut100fs5HR9GEI4VPlJexLG6Bnx9i5Xd1xyCla6SXfx9y8ju7zbjVHqEEq
qrVGR1d7ocIg0fVTMogacIQySpc+R0ycEUSuBVZWqVResEhrS9gS8BJIt2ADCqLu
tJFkVVT0B5THJCpx0KvQkhLGJRIz6u0lnwWMGkQsy4oF9SpyefggTyIezM2jZP4e
SBAwpBhC0l3DNFtuv/2va8kLtTj0CTiUZoMqY43HMVXsWgnynt6EXzW1LaJGdXg8
TFFzanTCKmJJ+4vZf2WxgvVXm64KJNyTsPwo7jlW7EwBwD2va6RrnMLS84NXLJwP
6iiqFaGnjIGcHyD+egsHWlEGxo2r1ommVk+fvl9gDkBzGLiybnM5i4Z/88Q2Gbmy
f4lTffuHburFoA74dEul+fzGqBfRpE1tmVY5R7nyd0pItbJ+rny16jUNjCuMebbr
lPfKbFzB/HjEIrg0AL2gMPc2AI/MnA2kAY0uyXwy3uYHxCfTcQl14CqpZ8CowgYJ
yzUWJou7UatLrNZ5weWUSTRCpDeQ9W1pRqq/SnmRl9X9wsKvaLw9PFFIyTzkG2GH
Q5a5I3a/CaDG+zrKloXw2sS9vtREYAXsHl/i6iif9d72H77LXUAXgNACDsCyHUDt
NevxXLTgzEtTZVHpWYZlTKJu+c0Tj67S8Qc1XgzVm3lQO6hmOjcjEm9KpqwhXTvI
KOx36GsSZtK5KTMJyXUps2XXeYtJ6R/bkx4Kzz47XdupDOISnslY7Qy53QolcMgE
UWVeWsr5DcoD2TiW/yDRmKWzBc3ZemR0YUcHH4cgDR2iaM2MuuRNdWOZsmLxlWxy
oDxF2jq1xOYrmffcgZ3U2KiLCP/QCewQtcxbUqlNYic9KZNXS3PTc7tjwZd6kR0S
bvFxSoDlBrxNYctW4hV19LZXQTsRzwXefDxrxrS0oVQ/Lb4bkv9hfpTM13tVJwX7
X8cezvKGZj40j0uUxKHqRb+gFRXQ+T92UnrindjJTQi+bnpKVjBmOBp1932oD8Zr
J4Xsb3h4fl2a3sIg/BdHowDdQhEMVTwD8ou7QW7bEPE1NsWe9YIpV8BE+aZ6V91g
VmREORnhsPGXMPPNvTRGlFRSRiwnd52+LgE/yc1X0p/AuYbfxoVRRW3VBKIDy8iQ
eMKDlQIZYiZW/k6O9iJAouFlzF5hUBfKWWiOW7N6ZbCz1/BOnde2KwIjBhd+VpTn
Ke81yotU0Ru+GyEoOcPY5d0z+Y1xd+weiVJQ+p+2/kC8kPxhmthX0A405IIV0m8v
Q3vRUQRCFG3jZ7ub2BtJmslws78CZqnFH4wFbn1HdS66/UYpQaYp5OL8vyT16m3i
LmmeS02/c7HvpyTv6pEmcZpmQB8EcgePOVOFB0XmBKzsb0tgls/fDI46/Cq9Dnbl
UPiQWpLMeTr6xoYbCdyRAhpdhMdqdks9k2WaAGp7rX3ij3dLY/EXNa8wm2MqAVEE
AkQO8MlUBdr0QUzx5J4arhfW3z+HaDHToupkoeoJQe8nTYMBS7+jclRV5k5iqJMy
4+uDX0BLMMTCmvuhQqG/ibpqVjUpNyEeGsTvAIWSgU1fzWCBJtD/966nq8TymESa
CDd1bK48v2cWJqpXA80BTx2NUKuKE57I4Tuzdsz5gCbiBwFV4Q596Mp02dR0LEAr
y5ivbypU3GgmPUPAoDoRvzV3VmJAUcA1JET/1m7t6su0niQVFzAh967BidfG0GGE
vngV32yS/rtlVjI7CvxVVnAG250uTW8mQQN18j3U/t5AkvF1sshVv3IpmZojvjE/
E2SKcDve1hFP8VLkaQnRvIcoQJYsagnUQycFCtm3xKjyJ3VbQp4iPuzfNtLnKSm1
zoo/ylt08pHFZZJ32E1gOIINKTTBoGN6PGRL55lkzeEUXL8WWjDqibrwwWrPL7qO
8Z7wZ8DCfmc27QJ67B4UvMz6cjHnlVQd0Xns/Nu0jFWo3gC/9QrWJSNYO1dlrZrR
LnI8xLLJbzf68/AuVcP43Jhc2ozWvxgdkerZGnb3vzyHapKc0G3bhohfEAfMOOEQ
2Vddy1R87ata72ThTPHie03xIeI74hT8QCF4yp5h6Bx3Il8DZM4t+x9f0Pnj3KxN
cI7v4Bf6gWCYcDthkM37H86jdl0DyO32lFXRlAkGY3a7o1ggPY91Mx9w4rQlwF1A
y1pHjNhLYpHne/fq/oSDsTIcLe3MygdWzf9Q925rdnP6wjsPM1xQ4+gRf/0jkWzy
v9ZmdnhiNpQpSORsxif4A7QPV8/haMgt+vHZbTTWk70vIT6yQJHKG5bOn/bjTTZq
60xoqk2V3hgb28lJ8wokcm+G3C6Rx1RX+ABzGdvq23N2mY3aCaMX9+lsXq48UYHg
b3Tw7PLUhLJnh3OCmYIhtQkdwf4tUFs8dCs0PqBSVwswhA44BycBPT1AZ0JGrG4W
2kBZ2ZZx7A0B/wFToInd48hYBD9562gPN2s5e4IGIBSgonF60TJhyp/clewyH7u0
Sg/fZ56oQTeRp/I5yBpzFM4fWkk7+wH+HRy27jIbVWhnRJvHdIKkyKZLkgbeHS67
/0DLwYdjNftkWQnKh96JLH+UuiygLU5dLM4kBUCgI4FXgglH8Q6kk0HaJUswRuBv
Tumk6P5som8HMrsnC28MbM14s63LpGy1FKaD+SofUc1dtY/Wdsz1AJQUru2lkXwy
L5ygDrTVO4mQcnbsWht1g955fIq64u6FT97atTJjszr/wDlFS073/0vWYb2vChnS
oscyeM2169p/UehOm8RSTXhxK6gjRk9XVUN3nDbxSKIIzlf9c3uX3DEh19CQ+n6D
XyrugxaOe3BZoP+LViIZLDJN054ogZcvAZJWhj8tbSHkQs6sARcesm+mK1kd9Zuz
Fm3Zz+3TJq5RJIxAPttoSoM9e6fWlhppxz/sRj/iAOSV7NkszD9Jh33z1XNXcBEp
YERwpTyvHci3HogrNY+7/3pQyAzvqfys04XLGMrUwaHctoZ53Yl9qFQ/wT/JeKZa
p8WvNLrd8wqFpZQ7jN3bYcMCx2klWwYeS47FreA4xicyg3U2znfjJvqbecPDb8gK
LHQrHWVDNnMT53xPmgDMhe172kITx76cNTn0EvHZm4xf4d/w6aTqzlVze6MssXHm
L4SpojMyJggF6nOwyPZD0ig1ihmG9/e8G9qPi89/k3GCqUxpDpQFyHEk0Dpq9lQQ
R+ZDgYSO7WgOc4J19VZR/TN+Zv1zi0sz6PkseGKSlKR5B/rjQd2yk98DJbK2LMk/
SSuYYebLoskvDWOlHwxHQlYQ3GPmYuFofKFBg4SoJ16H32c3TiUzpbRhdZ0JsDiV
JtgUyaci7ukIloTesEKSOt7eGZ6r6Gq8dNlMgbstNylB7AiSdKS5iQZksFeoZT2D
zKlceQ82xU0PyNr606QB+3lB6FyFdQ7hBt5TX1nh9ZkpH2+2hbg2f8Xi/Mtd02uC
t6J5iuMLMy8KyiZOKVzf1E+9Rf+DFNaU/+WES9GoC1A31UErdeKxeGPVhJ6LJvox
Z61hZHDd0JmlCuVWBg5uBiVllf6bHfrKSDJS4INVF1suJyRnjXN0ew8dMpI4fz2S
bLC2UidueVb7EjEDAjUQp130FajcNy9hOtpgGwwQVZcRkyo9/Onlb/XGNwU4ges/
efzFrehyJurBveQfCoDYEEYy34mtRjerOVDJyGm+I12yxBNTx/eeXwyJmy/GkfWj
9jiJiB0W/vx0eOyA80a4puDxjHsjurtdyFhA2cMoMOnDthgkD11a5kYUJSBxfqie
HIUQJ+wU62I59ThqYXhvCOsP37gIm4QMUsbcO1Trw9mOIAECQFNsvx6BBdHG9+pS
3MHrRGS9XlZPs4XBSYXtz3WX1H942FDX9WN5GDVNUnPc0yim/DHztC+/paWnzviz
5QtOATjze95nE49MOpJU+r7ZumlWu8/WW/5VQFRxes6xA9EpN56WaASSd8Koh3vM
zi1SCa322Xgw0id9DQRlmb8dQyziKYxO1jrxsJUf/xdTDTL3RPsjwgPhHFyypnqd
yrUOb9AvGx+MIHTes/9NYksTHpUnpieoFq1Ri0cVfzoAW4L3z6Z4ShK7/CLkf7Uv
AYCrWNSwzHfbpeBqB4TaI+oRkV5mhFwPhJZeb74yL1bqnB3/6HRVZZImTsFOVJRh
3ND+J/dGtEsmJm4b1r+fLTEX4B9S9uAYoMjl1q3ePISh+04DPrLJoGXsPj1oRm3U
AVn0eKVZ4YkGYVr7JaKYFeBLBWb1k4cg4LkPfkV4Hdd1u991Wwvvc2Qt73ki4ru5
/pBfr64jwB3vrxBOWic23QrvnoihL6JdzLAtbz654BwcoXfe/FzegMXVkRE8kK14
+z4s3pCn+YligLMkCCMaF9dzNL0/Wav8Q4J+C3UWxG8sMyWYJ+BW29BcJKEVp/hU
nXkX4ywwjLGIxsDVfX7lTcYbUYl0URRVdbKXDp5V0cQvx071QYJSnQw0bmYAaSd0
we8aVaQjcYcI+vBQv0L4YfIHCMSu2N+Wb/E2bSJJhT4SzZE1Ud1hYEv6n8uWjH5a
BKNzvQdve8UYs/IuITv5vB2J7AafgRuAEIxchYkSYuNZz7KqtmmL/MY4W7czEWD4
gKgYocq6sPzwavJrPKep2gwxaogpKs7pl0Lvme79Y/sH+dsgbmdMLxn9CEEWdNUj
8HKLl6/TX00PWONKLxnoOg4yrfi+MEg6+kqLj4wLvIgpK412RHjZcwxiE1CBGnIZ
bH35ENUzBqzdswjAa21swg+szVy6zj8nmVt5Kdhr0lKxF5ahQY80VrZhTrqIYaCB
GPM7RLb9/eT7vnF6jAg8UIjLxTUjMACjjfA+8wxefnX9W8YyTshEudian6W9I5sY
EdwWrTIN8eNMTHlmyP6Dmp7aWdIWHVAai6sIx7pWQ6PtkXPYM9OrdY4A9MyxzxKn
yLqSk7cz8IgqgzlVM+1cQcBu7M8DV637vvRQ/5tsIJqrRlV83pCd0T4/rgJow8Jc
enSDokNws0DBwFLoDrU6SDNe4z034BVVf/4ca17enTeB4QnEXp1I2ya4F6aR8Ujb
i73TWMFwFZBIjrhpO+ClKHfBoNzzBsL9qaK6vaOqokxWFD1prkDl4pXqgk+dxfC7
P4FaQX8DJl0qZXEgcLX852Ks/MAgyO26t/RYNs5Vl21LOViWbyLWgHuUnrNSF5j6
K3TyoXPZFcGamD5nqivsGDzNnoNvJRLt/wI8WCxll2fra23+JFF91YDK7/R2VikD
BTOgmrhGwjKHnGZcCnco87pMx/GPBWAvPxZan4uDu4bwKGa9rhoZnzhB7nj22Duq
ViAXqkF1gE/WkWCWS+wM4IrXQuE//Z5T6OVtCCVix2BMVv9S7O2/6d3/qN6Vitdu
3ChHeu2vpvbRArYyI3Zb3h4hZeDt3amMgcdj4TnolJlc4vgxzlhYKwm74m4SlYH8
R9BFYb8f0+rRPPTyuToySw4YT/XxwSe6IV+QlTfE/8hhfp7JJIpodH6VrVlqPsdd
r/GniVnLeIoTYqcqBTmkA30ZUhPjvpuR1YB2PtEUvgFIcf37l8qbbmURaoaxcB0+
jkg3Ip1oS5CIuXzlD/aX1/iUIcM4aSulBEY4m2j5y5DkcSQ+LK6QGwylxxMnioCR
NQPsZOoiVk8QEnR+02cADQ16F5+zdsbrIS3dgVu6+EPkhV+d/vD0IYt0JO40UKhY
Vtdgue2WIIn+Cf3VAUR28YlcNpsdcWfBB4OW5Bm6xWidLRkUliahseRUAZGNF6In
fqNHyYfo0ezp4uYJYf5TV9rtpYlhH23zTe2WssRvPiHNyVLbGoRWOoUmKO3EmrhS
7Uj41IUEhl6DZ9qbyi/rOgs8VCywb4LJ7LpO4J8fszDNY45ciarZUjoxSeC8dDlb
c5Qat79fepxpGs/TuS8qXx2MXTJPlKEuPsbxygjy1OyxWxkb/SR1L8TgGiqcUi2N
SMbQvC+iA8cbJu9ilNdV+h+H693Auuq7kp8wTQDYHNFX3JkwqbyMnaSB+R6TUyl7
0BYYXusBB5CHscFLZ8Gwaj9bl9NTm9EvnJLZDi/4LGyAwUJ+v3tnh0PAsMsPcEaf
LsPRyMGdGdaVYESxjRdOcUQBgp33XQIQZAzWEazquYlZvNnsMYUT5ZLU4ZgbiMwP
5XfKS7U6WBSuYOmB9RO28nFG9dUj3+iphQQv/FmkpdedkF0Fu3xYyaXt+j7pgJQK
kzM+C/qHamZvKnz/NzcPUxAtVnJajGy11cvqh8eYpaLJDtbPl8o1STJxfcGV82mK
MWrZyJRk2tmghfyj64epnZPS+DWCOZqBi/IqnoTn5U8DF8yevlpryh7qJ2HHgv08
EJJ2kZWW6Vh808g16/jZ6s0y66xv50x7pcozqklnPxcHRNBB2h1m9o21dL4FIXji
1WKQY2Tnfdnh9iT/YoMDrWRA2cifhMZalHkvWGbTsyhBPObMtXCntyvbwgXjqEvn
Saa/kzxzHh6DqlcX8P8A+4bc0OIV+MxiLq9UDXgottIo0TyKJSziK0uBdqE+z6E3
m8HcYFz2GPDrETaneSWo08BEuwlB6fexuhW2IDdnYFVZ/S2LkvYS0ojG05HaVUqC
yN4A4yc6QhQHgG8ANmKeCZNoxM1tdNI/twTuw7pZkZx0sl2NU5kMHLybBSkTMR1N
`protect END_PROTECTED
