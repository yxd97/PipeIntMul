`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLMyDzWSrhtn8gHbb+lWPV/zlQF5FKODmxOWVh2BcbXmsn6yeocIrssa3epoYzmH
IFoZpa4U5zOwj98W3kNEcrYBga9hsv6OlmYDMKwiCo5BDdsAfObc6gN//Q034R1A
lzI/Hka0zgjTVtiVhTl9dhnDzchizdHE/wIVC/ryMrQ8F5p7/8BXBTHnlk3OfzhE
nb2LQw/m8oELf09bQX7Ssr1SCDNtVCDQ/AH7eVZcUvhftnDNtLKXquguri9R6SeX
Ki1tpt/NQos576gLtOlZqBc73hxFjnIBB+z5DE2CAUidCK6WInT0FgcGg9HV2nmk
5RFf+9sghhyxXnytCK2wWxGYz+WCFDSeTr/5kZ7f6/NKXdmV1aJ/02AnyMBvnK7V
MbjRgvMCO2vP/6nqDZ/CrUAQWi624BhEqYIwaAp6+cRaN6iGetCyHZv1xu9PlRvH
tnmuYPTrNupUVCbGanrNShPpJ/Wx2iLIJz3rwhf9C0pZet18SSfufD6YHnuXNQQ4
RJgBdbwKr3nNvpxDRUbmGqT+byVZXvZoSFm49LTjYj1ZaUT0LF/1HFt+JK8Xewma
BdPWP3bOpTFPBbgYP2O2az3F4v/j4D2JQDdCtcSnlVitKsii3uSCdMK43+4ECIij
kGa6+qM1ilhYRslwiRqcvTW9SpcymS/MPW7RqeMPnqE7Hyf31kfYa8MUrz59umFW
csGQu3iDvSXIPij4Xnoe26JN+fAZEAZs1jf30EDX04GM4m7f67CfXPCXobPF4Xec
NMvjU4LFgkqi2hEvsazzQdJtOnhaq3+mewOXzyfNLwzVHSbHYThuF8QHUkm7D5Qb
GU3mDGVjdODbdyEcAhX15gZA2hX1WQLTP8KWyV69eMvyevsDA5DoGDh1i1kIzrE3
Ye94V28RFnEzikxVgU6llokadi7b+okZb1UItWGCU12V0ulUUe+TUhYb7uN32ITL
eS50WeQc5RaUqevqwDsooR09x/ZRBbkjrluRksUnfhms0/xaPoB75IPlb4AdHWbG
JIUFu8niHsmz+mqxtl7B1ylFAxapq/gnjTnFpRO8bujb9EoTxf+kvjyJfT65GN9X
XJ6CcX/l1gbod5P9iGkzj+eLy5qLYpIjXGU3CEBcnSMtvNqpTBD2+48UKmVrlQJ9
ZX8EPUXNo8bxHwOBImoJqYHa3rsaimv+J9dA0yklxicV9ikP33YBMn21RP3prZbO
5GzmmVAA2CEc5rc3ZY1ntzvrYqktaRISF87vutNQVUJ76WjDYJvfr557x76lVoU3
oX9kkJHSc7uHLuakuYgMp8L1wenbVD3PtlChA3FEBzx5BjeU2dYeq7+wgHyNu73G
4VopP+iQa3Ef2XhplGJ7Md8SP9lq18aEqWN1x8RvwocN4GpBMkAZ8l0B3oOH3jo+
1k9BStgzYNsqLBtwF7c4EuxrNxaEciyypDee/RhD8B25RYG66Z2f/QPJ3zP/VhGZ
cR6NRpwmPHvZpsxeV+OBySaGfZwVKh4Y8N1rvhy6J1yLT5wXumQMP4tgd1i6sHwH
KETRKuXAlN1orwqs7viYR40oKqalu5RMXFZW8zdTyoC+wgbUO+Zi28OH4z3bOQT4
TjR7Via6QCA0eigZ4bvLMol/t7/p+kIWjduT8zDEHya7oAj/z5ECOQIf/LMdnRtv
l6BNG2iWT8tMpL7Mc9Hkkd+oefjqlwXpugqFk3DhYaxPv0tedfHk2Wwur5RXMvHW
ttljMSsYqEMMgoWkwEhk4ZdYEhXT7z49osY0DyHjvPmfi4j90kelpnXMzGMHNtFJ
HEOE6FWxSKbFWm/f6SN3mHuJRMX53Nsn+DnMQfbQwobQLSpE3gnvo31XO6cWvMWP
RIhfvbcZXC10T//aPa4AmbjGoetczPi13cBoh66rcq/E40TywPX+CHfMbRcpxIwc
mNImQTd8ZpcmTvbMToI/Qkuz0homETOg5K0oNTvGI2ENa3UDhhJO1rVaJfzs6c8p
jOj61yPSLviNvMsUXUm2pxubIAmX6Fkwi0z49ZRxKQam7dVkxr5baSrzzr6ovoOL
HbcH/rdo7tQczbAGTAjB1tFAQeqmiNEz9jUC+BFkmErrkO9JNxrebCqaGnru9TD2
JPv9YxRXrXasYBLncCbujb27MeMIUDl25R/E9ZWOeD4P+QDXjLU7UPiPwU1Nu0ZN
Ds/0YlDUq+SeG8q4A52U1a7doss1kJEwE76iHIOpoi3LbfuSfXE5KYEC2U9ahWiS
yP3Y91NGYzAOBHqHExRPd6dtm2QmQvEHeQFEAgZsFTXVswn84OvjcMco9m96xO8+
rCxnpcbFZkaO0V1eGeKwpscQeF1+C/2EOXdGWVZGrw4IeeNLqMkvg6Pwp6XkS6q4
N+EwOv47mZHvh00D9Ju33iuj9zv/sIDJuGfUNXpK5ggIfLVfAwPtNauoIFZzQI54
k6MxWwo/Ccd6J42lXDKuw1TDAnd/fdrCPKOuucM+rQa/gN0i48rNZ78D1mD7JLnG
xLbzDk1Tt3IPVACk9MX50662t3o6meWrukeOLOMwr1tR+SFlDKEKNpYFHr5CiPxF
zLD8w3qN89MpX97y7r6CnxI7V91qEcLwBubgjw5snLcEMfYGpLOD0BEB9LoA05aj
iyVGx9AqcN+5GrCT+lMFbvSRIgjUqoFHcymri+WzOyZh/IIpeXYkdbVqudDtP1Uv
5dOMG81PhCGwR9P2IheP1Ah+YYJIYU6w1abeVzO2YIM4DrRvoD6Wwgv4rMLm/LHa
RtnosgMLmhfYKREAxyUSevve2kozVW0p7SY90ZDkOHdyvsk2WXrCAsol/txtxx2p
IIoAtVyw+QcwPxzbgrzD7LxfIIjCjdWpHNdUijfRMpnJY8AcLO4z9c/K8VNLH873
`protect END_PROTECTED
