`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgagQFYLCNqEnGm3EsR9twOftSsDEyuhV+N1nw01aqy2qdym9NnEWP5EGs8cAM+A
E+px2+NiHJwD3qczD8wyueNNRU9sF83kOFF4WTKjnMBMQRGD1HGpG70qNAdygZdl
X3UiHS0sfF7/upZdRCmZPGe4S1RR9T6YYMGtgy5dqPUXZvoJNTKPPXjLMmPdiLef
hnsB9Hb/+17yw7RCR9AF4icwpKCqZ4Czmcu288jCibFVKEsLL/BOCcuqiA0Dn3MB
quJqgSYvO+woPqKblOnjAip89rplvahJpVZQLd2/uofOao2fGcTg2/dJdIq60ONd
NSo11GLPYfwGy8fSgwKD1zOgeoeD60zVx7E2yfTPOlafo4Ssow9Zolon2Q6MlQr0
WjjGV9NFRSJp1R4hzu52QihXS/CCZnz+FiqeQvdo3RUsBDZq3+YKZv6VJaXSqWr4
ZoregdZKWzEMNhIMnnuV7a1lVDgrjan3rowcTj+JyNpi2AhM+6O/43hLifqxy4qw
uxNd7F9hpdKYi4kItuUcfvK+b5dHQ0brZE7jkrLA3jkokEEANxzcgtmVVZq305tX
e5TY8IpgZ/rb8XW8ryqM9GrpRUH7FXRY3Ud9Hp8PpoE0LHJRhC7Wmx8zVUhJdCoF
Nk5N6pq33lKVw6NCdTNv9PNJbSUrDoQVLjobx5lkRldz4vmPtpuNDTxzCwiU9i5V
iU/hceDIqS5RkSpLdt7Y0ESgpfSM9gnk+KtT2SRay7C6iuMWCt726h875KedRmyl
`protect END_PROTECTED
