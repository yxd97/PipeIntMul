`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Spxi0be4WDLyE9ORLfWEBAMpWuXfcdgLf9096ubfSuRHrYbi+nPWLLwcSHiG9rOI
wNeL7W1AWCjRgC8kPmGE2L+IoYoiQvvQ8k+rYrtNbdLkrfcl8TzclBvQmgXo7MFO
ITCG6tcd0r6K11Ylwhpvo2L0L0S8H9gSusPaRjmvtLt2QFWpFOBYD56hVb8Pkap5
IGXij8MmAromM7tTsvcaPJVyDfR6WNRwC83lXU4YnFyQZ355EtGu9wpReTc1mmk4
/g4Tcb1Y7EIOYVkpvLRlq7jLstGf+rQ/+giUttIhpo9PuGVS+BNY+03R8D5vXhV2
9/bCUmYac2HGnOvR6/X9oaUkH9+e8oaeb8Jb3N6QjYK44bfa0UdI9kcmyuDpprVM
lfnznFNApOoEHpZuwQW/Lkg/BxqKGgMsUlD6rHLQuv/+PgeyQx7ANxevL082fuCm
pTleN3YbV2+It1teCEjgdHGCfK7w/YR1L1BZDFxhH8vkfkqPJEh3tNoq+3Xgop3G
I+TGqzqXZ6yVW5CMP7wUTmn2AUT+8CIU2JcfiMsIrhVCgLrIAE6feDKbBVsxqK7w
gZVd3xkGBFEJrdMcHwPOnT3GwrngSH9cMmExlorpE/gNVlbRN2DCTIS7xoEXyI/W
a5Lsmv9WeoglqkuWlMimWA==
`protect END_PROTECTED
