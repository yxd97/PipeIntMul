`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qipO7BXIJs1sMYnVypL8l4vHF5p2+0q8QKb5xTFHcZNIpKGAOq9910UHSZQ4qxIy
P/yKad5Gkwd4B5aQ696bRCJSGgThIRlTggemntXBCe5tZMpmKkPEIncxuJzMpALv
OziYWNw2ixkhtNR8owuPy0foWRNqtMoIEajwyB2k52SMHUQ9FQajKd9bhkjqMEyi
aKRJDCUGPF0ijX3G0UEbnne2XhYUCV2yVYtHn0r1na0NKTWCQcCDLmRWwrFW05QE
5wDgPj3dwvMWS1vKe2+ldg==
`protect END_PROTECTED
