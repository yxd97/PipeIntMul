`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Euo1xEz4cDb2IeCA+cvbiND6nvT8TTR9qK/Nk1dzGfBRUuac8bQ0O/0Eh09ldeYv
FIENXmcTIFoP1saABxfeIuDdGSnw2cenWnvy5n4rAssp2EpavaYYpWlSVdLBJhgm
UhFrdaVhw+kvevEnbjy1B2v6JknTrF9xXTS1sAca3m4xPy3TkA41RsFhUBh94aMx
l8se5uCPoexHGh30J5Kr8nwdJyYW8NcAevs4OcJxLGTS4qOhAnvd2jAdX9o7xJ9B
vsKgHZAo9CaEfIPf9KAfojxQ1r/LvteLam+lgMlHrCzQt+oa+5FXwX80oNFNYCMN
rMtJqFlfdRrhprbhY6f5wf+2zHRqrSJd9rnm7DQyHf7QtosAGwGHKxb9zvOQnztK
p7cXTivpTJIHOXULNdfk3AbaJM/851Kf0+m9KqDMyC1WREDUrZxxqC+Eq0kGz07R
rwLAGcG6O/fcrMPYqsQCF3hPyYhQ+OXxyZUIp5SfK3uIa1jVbLmcjPfn+Gvikt6D
RgVIH4AFmfStTvgNQ03oh/yySDVskT+1locAgBoonrnA7/gIkiOghaCnAC/c4Us7
0pJQ7lGe811nL+R4LZOwFhNJlW0rSbZAfAtCpMm0jkk/00X+MM/2AXFZeat1i+W+
lGoMa1+29wtm2HKKYr4Ah5lZ0Xb8AVFt8/mEtkZDUnQFPFE99Qs/2Oo4Uq+gsFAV
8OVqeIVwxkguoXpE4vckzKHHPSE/RTaBasv/pugSqVTLq/jpKXhhscnyvV/W8ogi
825DUqRIHD2j/JKD7aNpH3wPv+akqF11RWaIvY5OH6Gwxyp1N10WtN7GJaqWnQxL
t+GLQzpO/MLC7Uamk9uE92KdYS1iQTjEw1FlYTJMBLCbk1fM5kPYnls0cRSmK5oS
Bn1AyKiSVCVam1rhV4fRv2wt+H1f9u1VTLZ04HEIF0MOtEYrpqyJ+6Anl1p1JZrW
yrDcR0eShfMS4CEWdBBVMnXBWw2lOxx5ceWdJdL448vtSiqA5It1oDzKIVwIyhf4
R7h2iuGs8gS12FRMmL/qrf1V49XKKeCe4fppMARupgp295e88sN9sAY5kAm7EX7a
ETHVecFJQuu3mC9g1dXkrHBVqUQnCrsh9t875yY/6tPfzSV2ssZjM9K8auf90b6e
Ah5eiUElZQWZKw+evOWQf09NVG+Of+t85gnWGJp33QM2oM0Lmc5K0Bh2L/B/julS
xSOAc2oiyrQqRoxydNyM/juTtITkWNDBOqVJz/d3knKuylU96NIZ5Gv82YJVK2/b
5EVrNQk1bvQeFe+jLozcZbrXcex1rIqeBd4xCtvVI0LhEYZ/32x/NTw5ei6fm8FQ
YBK3VULJRYqKl6eAUkOdLo8CRWw26wu+w+kysqQs2nRisD7Jlrx+Qj5anvNiZbeL
7miDK54cU+QT3hvr0T7PvYyXlowbNGsCt1AjpRQ5w0ehRIwuYfgWuVnztEm52S1l
V8x9f17GBMTePszOl9D5neItaa4A/Ft9V4DVuXZyk33AGxrDztb0p1sAPNp9c2tA
lwM51wsuYz/9yNoX5efhwdWiVemLssvGw7wfn/tOPEtGV0SapYMP6L8jQ5HYPYEM
6edIx47Ljiu6RzYjesUCG6ZEp/IVs2jKNUTNtqf0O4HdIilaIvbl8Iuh5tnJZB6k
aCJJA/hT1Y4qFY46ml3Ejfp5cBdLrc4oZttXzcGUuYihSD0ocrOWhqcgiiv3HfTb
DzLWaFAwqXCXoPhm+yV+ZvFBdsOOR3XvIg4gTDVcnbrBY8ooKhP0LDtsr6GVnbXV
PsUgekH7TJpAejiWFzNQMkj1OYre+NTHbu6v/BvMwTxnF7VEX46EYkagOM2OrWlS
y4lRPxawqGTxTw+PS4EGnNxQM8Q2vj4Y0mUbtq+UMaJfxb7Gc9U64pj39p8whRjf
UcKaQbeU1ViUQg+wTrnqhmB1woUrK5QG4Hvo1TkX7OLNvUQXZgX9QFfPd9KuF7Sm
j7emE1OcUK7wagaUjVcwG8NNEe/JquFbwEO2dD+3wFzGBL+a7wKHiNX2j/2JnxSE
HWv5+KCACW6TgzH9PHfPjknXkbNL7fvLU+x+XoFSCU8dwLF+PXqc7mmiw9dz0lM/
SrLeUS/7uR2ijl6kSBlAnjTDIRik8FLp2aD3gWnCsqqIZNtU+JHA7o9WNlWWPaiz
+WNWWVgfPv2Cod9aL3cF5p2K8pP1TiQaysXJk+GqDILyX9Y/M05XuKxhEy1ZARL0
AIKpISKvFdcpBH24OOqbAVYs/xkPxIwvKxs4WN2igaErjqCTlfXFzrmReQJfj68F
IhFZQVivDlgnjCpqpYvxedTJMErP7s2LbFVyKabmpbupg9H2m3NqGNzVPuqop2ga
8o/7jM5BoLMFKD9vLulEnpATFvBezwUrv5lwNcBqvIJXNuZ6Z7W/1HR4t8HFK21o
qWcS3KdGlp42TIsCc+oSjOKva3yB0xWjpoBwoadAzbLf75dBlLAC4OqMkes/kZL6
INrP9CNi7349z1IBqx+PmA==
`protect END_PROTECTED
