`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lzYDiQb3xk9+Ee/e1JDvLMlYsdD9cSFXTzWvgbG0tb9Xi9JGMjfTSbb7CEs8g6w1
2z6x5859ucHp2pSCPi21SYz0IVe2r/udxuybrpi/Mo7RRM7u4r+dMH764aOaZ4Gt
wSSjMprIIAEAPYzJe0wESHJkiAmJielfykI6yyzu53R/bS5s4vKg4Hra69xXXOoZ
E52BN7qiaOx2ykFgV/XjPuVmKGdmxWgvBzupzDjXQ4ek4mgHFmBQXSnVAIWPrvk/
mRqLBbcSAEQCiojDdxXBRFriOkrmgqmRjYOBo7w/z5j+TWkNirkC+9nDKuCpHkFV
2/azPd5uJkbNXXwEYHoR3jyuLw4MjWUv8uL+XtC4UgjfkeORcyv9GyyKABaT0o0k
WbCEVjTixeyr2mg6jXcGuxJaVHebTianxp8jWjtO6rF0GfjZPddYzKQSorLvHcBj
unj6x7NN3rUfgG9X6O0zWwfuVllOVuDpGe1cPxhgGQZDwW9+HHW/pTiKlMWvj15H
ytiTFpbheN9u5vrWoLYE2JyiZ/s7NYhaiGmHiez2t8L2pDqEXP5DFG/6rp+095+h
tc1RdvIITzbHW9sFyerV63Tbh2eVJ0XglTqIJkoEPSA=
`protect END_PROTECTED
