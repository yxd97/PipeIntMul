`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gLkRPd/hI8pxeizTO8d3AHKFRY+trBAFgjBJ/O6h/GUvtX33VMbwggVNsMZPLsKy
e0x071JTCr/On0+q8FMw566ABNj3xDZWeZgrqkl769Cvp86PK35hNJgam/GC1ejk
O0zHAxQ2DVTcBP0JTxmL+4tweieuwFO333scohiFwLnt0PxM3/85lSp3JwXshLVW
xYdr8Ri+sew7nbT7r5rc1sAxCweV7BqoDqhCg9wfeUGvtBcjSPZ40h4mbCDbG4MH
aRKw8LlvBIFy90zyXZ9lyriFS9WOpVetzQEQdapfPU2shWbYSRvYFtfrAHJPiTPH
1kPQd9aBFrTOA+0tncAkIzs4eZRB9Pd1oJVdtno7htsCFC5IhqqfTZlGDb+YISQQ
`protect END_PROTECTED
