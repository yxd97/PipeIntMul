`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKOBdziU0mx+yB9zExEE/22DOgZMxTW2qVqgGYMxdtEFgkwNl6wWYLTUGmeXWru0
a+vn2qtZUAtbEMaotPRb7H2bR/4b8mzJ5OzHs1CPu7JT1zPvyyw3NTRliR9x4QnS
Bf9DPiJdE7lenaDIe/Xl1E5YyBc1nTWIA5GyyusrkKYS5e4KBvV9UZYiO58zoCsk
veqkZItlZKVkiAOD+BryeiLTBnmFy3oZ3XXbOTfGAjgBvrmSgaOlvb1cRMPqixtq
FDdeycylbcsYeFWvhIO90iM7ozLcPET/NghqxUCzSnk4kEfK2dJNt0DD1fKzXU+y
ToYUshSDT52MNtMYl38yJUH6CQ3mN2dJY1WzunMzzCU9ySdl5PIdfo/wXwz6dBD1
lzOKBlacsUXfcycDTS192+MEXT3ya1yNURwwzh9wFOssk2sA7yw7BbHCZYtW5+Bf
7QoR9PC2mrF718bg1uRolKRpnsT3IrKrXKexWhLAgAY=
`protect END_PROTECTED
