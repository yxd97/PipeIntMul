`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cRijFbf9s2LBQDNUpm6/c93OsUqRRSDWkdBjMcMhOM65v7WYfkPB9R3Qu41B6F5B
+X4T4qhGo6xwxXudRLgpvTo9/ysXgvKvutAyI5a+3QJbhQIfqgZL1VNcjhDsMrgG
4elahxrXjpUvSWhJ+RgyjvHf2UYkCEhvkQ4hBfUv+yKlQxwa/go+4EN+eYM9wUV8
wrbFIoZwaSL3TEn3g22WfYHg6GNpFcNFvL1sEzCY9eVwAMcpRN7btb9FS4qhqR24
2511xnQtFAEHSW5J5DbfC/kPAKwZDFYuOTN+/QfSVuo=
`protect END_PROTECTED
