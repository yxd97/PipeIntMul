`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SK2qp6DraADpcY/4A8aBvtwxZKuVN0vFDKZuE06Q4I8baaoObP1IdUo0AAAlvnlZ
BQtED/6V8z96zUlsdSK7ckLbtiH0IDJhaUiibQSOrPlRiDU5Z3q9MV7gU9ZO3XDP
KWm57oovYmFA7wClO15U//4t1tq6a9HJdQjZzn70oPPS4jhyEx84MoAMpQ0ZZN9D
Bv3N4x9d6ezsNuSUrZAzjtArEndzStnzd8OO/NnfDxXQZrU3cuvKuHrIVoKlSqTa
ziJTu0yZWmEz3HYRtIBGdz1inLRiWAVQyYtoRRuc2i47EXnkXM7ee6yYo3kcboev
WXlLyUB4zyLrUA7ZvcLaxlUSWjhBhkikR9z86F4rCsitKZ30IXEyHsTpRkH0hFAU
JZKXnooe6zdfB+hpSFzQj78jZx4O4VS7M9QFmrEomzhaRqTioMn1E2dsYJWhOI/l
foZ/sVBMYiQbDTEnQcZ1qJqCP8eWydNWMzsahA2NQ+rGDKuQ9dEkqDbC9O+QVFfw
dqHB1Wb5BG+VBpPa1CVIslT8IVoatbzOBC7rNXJ4L7hxUv6Ie0nq5U6zDUnMxjHA
kGf07Fp4kvRRgW/XgJLX7KRJ57PtNHhUvj5iXZvHaECJl6sdJIVJUwQPy1pOWh/a
akieTBZ9FcMmOhzOgOjjIZkvZdmC+5dpAdFMb9Q3VLfDVgHDrayA1kocENE+1O0M
euguBknI+qfwin5+8xeYiabf26a3Ml2v3MtCVKg8kihsqRx2SEShCPmddBnwWxlP
UJhcmxKlMDY10momJe78cjW9ozOYR91X201892Yv1jOrVdYQiSzO93lyP4WeJktV
eAfPlOBxIheyh/dTnKhxcNvmCornsZupdpBO0Q/JdDm6F8tB5nT0COJEsVH3Dai9
EtQYsQpjX9GOZTeOILXloOARzbnJ4TCAygmdd4/S0zAMPmw97uINOO1bJfoW3iBL
dDTKbQMURgaaIZpgKwVcL7+wSxd4ybn1aXZZPFFJgYyAbwerPuuuWP8Mx97NvJws
gBk/r2f7l0YRaKcnvzOE+fftHSHeXP7hQ8dVhbR9NEk=
`protect END_PROTECTED
