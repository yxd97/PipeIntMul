`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2bL6UdnoHhYk0Cy7h5p0xVTi9RN6h9HM3DwW6NAXOJBDMZcc+qlD0k7BrE8UKbAQ
JZuGTdGcx9DKQCdjc/kd7VmQ78hLBNmU6+Ua6eY8SZGO94KgmODFX2enFKN1YBbQ
vSU/ssG8LjimuA4hcwNxbgsrByRhzGsnjNLc0EddQloofwdr1KC3jlk9S/8CXCAc
SWaljTFInzQqSMuKPQcG4AT/0WLvp5OIYTYQA4Q/9nSgc6Sm6WIKNAkOh/xXDBSr
tgXoEAzAoxW0dffsJ+V43elzYRi+hplf2rOUPVSUOLiN9ndCTXo+7MmA3i2AjuPI
TQd1Ia0CjJ2WNW6QuO0I9Yrh68fvYu5gs5C/Je7RO8XKEtOsNAVItunWLpGSyx1S
qtPspvc9wHHImjGS/Wk1UBGNddfUawLWCFbMdHR8MwTKfx3knaPKq1HcalJhOt7p
jgFMDWx2NRFCBmiH+lkQt0x8AvOZ3i8+hieNNSV5jtOk1wNoP0Bo+gXdLgK0jX1Y
eTeh2i6FpCr0B/9DRvc4LoNGjaj8yFc8wRxjHkjO6NFk8vQwnVoaVMVpFl7ufiAX
S5+p4CgrJcXCtKIDxkywpw==
`protect END_PROTECTED
