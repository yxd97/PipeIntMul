`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lQOtdVPkIYXgJgpElC8K8MJ1vEaJh26y+7gpDwo0rkykn/P+t5Xq2nGOYZ8/i7uz
zhoEon/AKWAJdnqCezJiHj80Z0yiLcWkKEYkO6PaRDt7maPhrUyUoNmZss0q1B2s
y6dD/hwTktpP+b/MxzGDZwW/d1eg5c+z7rSvqxaD99B7FiZpQLV3kX8wWd3sylbz
pODLD9qz/s+p+Q76Z0djIStMdMkwyfnKY+gGwy0ON8OxGIVEEocRUFb0FWCG8xAo
XTuAql+SoTeQbPKSk9QV3o6oTwstFma3LmzRt0nyE++Irp3KnQD2worwAxAS3xCT
VLN37AtFL2oJzw7heUN7YgPeiij9qf+08Ko1CGCfrT6bSCH8BOW1jo+w6ED0Ius+
uQ0NMW+s/qWg6MKWm+9b3/o/Px1s1/sSHEb10FC9AwY7SWuyDAIUQnm8rA3Hb4RP
1jZ9ruP8N/NOEfxn4lhuj6y2IiZ63BdcdOMWp0KsI0Y=
`protect END_PROTECTED
