`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4NqyoJhokEb8WuDknkH3tgLCVMxDpEYdCPlqydh4hlXkcdj+M1vNx9j+U0gsEovN
wpL65ODWlGzBkJtbv+hOzwQmk8cucMNTQlN3vCjCrabhQ41beYZaA9veYvj5U8Nl
ncAT/9vun/jB9Tl+bFfSeo5SYqF4trCwyP5da1G1/PL1xuymlMpPa4hEIKJECR27
mAV3kv/JC0gnKcl3B83NdL3crX+AqOeHbpx834uF2N6Wz4SIkbrzfyqpItb32TO5
ud+NJGbX3vMkdwjpn2QQbJI3uQp2aU+cZVnA7FzPlNi2ryi+0H76aRlv3JiqMSGS
p4Jsn49klc+7gVHR5NS1Wev4yzUOpP/GjTdhlGceaOv+cDrpvCBKT6RuCHJ/XtcN
FqpEvPf7wrbcWNDt1j83kqJlSLInC7JXZQdYpU7ysf0=
`protect END_PROTECTED
