`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DR6UUTZYNEX5nW4H0Q1M2mAEG/k2UQhL2ymtT4UqWTsyt3AJmqLWXSrcYAr05wKP
R2kZetKyjrKrlFUAE4N1yIVek0LEt6UwLbqNU8gXiHC0wp0g4N02fVrSkW1+Tkhg
yzn+dHvJytZZMrE5Broew60Skj3CYdq6d2bsP6Hf3b2dz7NvfSbSSJh3dsQoa9KL
nwqQ9Ladw57X4X6rBj/uxhQCFj76CH6Xa+Fm9T5vkchHDSuzkCfxhKqfjwoHxypK
YznrjBjAq3niY7p8j7Anuo3AzFKyG/A0Rv3XvqSMv90YnEMI2GNP3APi9gt1iXA4
lG8TbGdS9wtLOluRH2FrmFhWi2ioNox8yhvHDeoOv1bhOQvlGWytDhYVPIQVX8TO
jH+F//EOkupGdnsfWVAuTDBrx4GPqGjgT/APexwpADAirCdxhPX2CCgQJ96Gnobi
dxxuAJQ0WPVeoSJmAjgqqBbSTJLewpAd7gpyU1IAKQCr2YlF4kX7lqLOITLwu54w
E/PVcMIzIE3+JFkX+bujYEJvv6iXEbXJJiDgRJh2LrkXXlRPT4jqRiEF6Kl7sONh
dekk3ezmMhHclIi9WYSJBriuz4YxYKfkcsssdgnlVUC4wq2SK3DwVDs5IWihavGi
zGCbNcqxsUxwBAX4hVq96+tAQ4WwCTW+IQZj4wowVnLcNaeDmvQ67zSgCi91OQLm
5HJsIEaKN973FkDlk6UTf7vnRjfUOcwaopDcu4eHkBqXGJZvAqHGuDnT9gvivgn3
`protect END_PROTECTED
