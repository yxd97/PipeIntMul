`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GgA/syNdulasXVKUk694V2xiHzCRW1MqCdUSvG4yZzP+bTFbR0PJtdd2e9JbDQaF
OU9E6/i7g5H5x15cVy5om0TkVAMG3JVhEU+16jZUk6Wiqs9VdHzeIrLvsWS53dC4
rrybfrHwxhpbJm0ENLkpFYl75/nQ7570Wfl27Law8pIAbOr1Scq18GqdDdqX4odq
Xg0/RZ4oEqnfNge2Ow26Z322wfMgHpSVDp8TbKJkrPkeCBVs1AjEiq6zIsavWwA+
36+NfAcCEoDhh8hksIFCnc+2uozh3ZOaYpf3xFF35qBICqUp8T5/XB4FgAxX3Upx
9Kjol2lMRhQoFNqaSNRfW2w1gml6zYQic46ub7rOLbnGB0DgOmfs19HOiS0+ga1/
YZ6IXTmVhpaHbDq4H3VTdzIIEKdsVScwQOVxPuqYAQqVdZa/lsePLyOlz3zZWSBb
rEzW883iZ4YiS6BuOOVnhCD8Owk2IgkSb8AN+BzjsGWpysO+ptBmHURh+QR9ApWw
SH1TO5uEEup6OwdSE3tuQQ==
`protect END_PROTECTED
