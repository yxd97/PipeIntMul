`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QnJbUIImZqzKT6htTHoVsG4XLhUU9bVTrRnLwrU5ZJxtNSJ4uT8zQjc2KyZkH6Q9
VUi6gDZGcHVNB8lY+x7Bip/og0lY0avIJGUFh4ulEAcR1Y5VJCnau0i4hOauhSW9
A+DZ8iyEunh+2F3o4nF6opiNyGGgwQfRvfPI9T+f6SMwNRVwhof19V6fu5S3tHiT
eVQoJnShEBNIhigDvieGGVjC3aJZDgXHnHOskUngwi16ADGyOQaBudT+BnsVCMaz
ovVhV5A5m+XNOf40S3G+H4pgAkuN4OkA3wabLg9exvrHpDR3Q7g6flfRNnUzruJF
7HqFw250Gk9qdj5nM1f+IX8z6gI0JYtfXu7K391Uh6e8Mk/R6dLCB9cBkCYJSzyc
uWei3XoGyM/4DZE6oDwvU1vss7fYeI2FlDv8J8SBqyVyU2n/lDmY3S++C+cJXmq9
6QlusFbQrJql/vP7jHxG1OH9I63fj/T5OGzFjb5YiT8UfanJ3dAvHCQ3xHooVow9
aALbI4EJuXIVF2N0Koommu8WaIG3XDgPigDWFDUtTYFcytZTUhddeClwjH4mtnvU
Bh8unkYdDwMveUgKMtMw0/4lzHZWGmdwmufjMviAyNhk4rG0hvLTSoovPprhqJIF
tK1drdp9V8FPOl1Ya2r6PZ9HDjY/w10S+gYWS/HRQnLj5G4qC+uwZhiWrQ8ZOiSd
EThOGGdld+1aHKd/iKA6JSCntGoURk9CCvc5SWZHeP0FvXS+XZBaCvngmHBeqnMv
9Ko4qaRY0r2xBJiqsLDdmolzLfVA02XmBgUmFLnX2HzcQL2921e8QWwUAOfSzT7M
XZfOYxlB3ZTT/lCboTM6pMGi/tQ0618QJusByIOtzx24Yx6BMmrUZC/F3TroHP4v
vs0iR8THfY89qjDVk52A8HYgBnWZICd7JCslH8r0Wl7Rjeg0zwyQpXtUzCBuvC1Q
n5lLfBWEkF54WDgVnKmgXtga2CaW0Xxb4p3BTPUFAu0ZZiD7WZ2e2mc4UaYSM71A
bHrT08ZrPf1P+WrXpV64255u/xpHYmq7sQ5YAX4jG4nxeUEOSeI3Z057ofgz8+Ro
MneCc+wP6Rhxea5M21H5va1GrYnSk3kV8zYpNQO35xAnydojgQmhov7a/K1SnJmm
jycTC24Lfi0d5dTs0dPi+2rP3h52eJnM5fYMBZLubk4hZLjqg/8Bzq/mEXmkG6/x
43dxPNhid1CUgQGoOdunbTkU5INl5wTulRaj7oPNDYPzQiTzaCFjfkIONtL5oZyj
`protect END_PROTECTED
