`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GmauVedjOBc+TjdOyVywlh0EdFfFWnjlR6TKcdHr6qCBNxcqbjkXpZ706H9ovLeg
u75RPmLd5hf1ZR8wc6K+rwdH3Bxtlf1ZVnk5Y39wx2fZSwrtJUf3jvKsnV+dJC3t
J9G7pHDUur/bU30fJ2aslKIjc1D7mtwa5wsu2FmHQhP96ff/L5PCl88JutcFEbYH
L+waMMFlHRBLjSnONHjLIYkN3egfm7GQ52z24m39GPjUySOfMufrwh5hqV5TIwQI
mquA/xs+OrpCKGBShTtivRrfCjv6fF8lVLtakdl9aVPtzkWXuxYp1rTjnwm+mJjR
tbbPtrGnKOhcPQm2UTbseLBy5YaZmuzvO7vdZL4gpg9cWcddqDC9Ba+4RQ4T61iC
JdTbb1lCsovRO/zS2tcYAyOEIqOvaqHhLov4kgVw8yMQRa6E9ipu7B2umzc+hNIH
RlcVlV5zBJekX3l9JzHEo2vZjdSpEC3dTuxrP9hqmVHaAlcyzUyOG4NeftiRfXD6
4anxLWVGZZs/1kGpgAYITA==
`protect END_PROTECTED
