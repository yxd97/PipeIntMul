`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkW3o6HNGIOPejO1pkT8V8t7LhyPT9TmSiacvTt9pbtPdKfoEw7UZIDFEa/zaMBs
vUhhm8QCFt1Zizb9AxVvMj/R4mqs1f52gspi/21CsYWOCK1V9K2cTMxpceC8nV2C
xmUHsPzHkUyZujvz3l2fHOcA0TaPcvvwDNYHgg2u3UFfrpIwDlRrSwMIck+9U9Df
mbWxhS9uKoGzOVsg0WQi/DvmYbVHcJ4mkqT08/vgB5SzVxM6YXyEBG02vPzIoStb
XEBF4egcyBe7qCpTz50qhTHtXmUYBgipWrU9kpIGoQQwaC7M41b1ZsFNkUSsqe5H
e9bfOsZP69zZTtvZgKvKpF8506KUYAAqhour5f/a4uQH63P7uLXVZeU3f6vjfXrv
cG5zsGtFW6AMWliBOSEKcuOUtCsv9jwmQVMrX5Q61WjuwYim+5G3QY6301glaX3r
PM48eiawGELKsAJfGcwTQ4nOwcu4YKLvVDfe/iRci3N+IEOCp371R/0bD5vN+AVO
3quBIlm/BtGfJQyC5y3ALQADNslxoXX7FJIvII0xu0AuCjM2UUhsnZre4D5eiHSG
tSXR80x0QFweTEFkO7HTcuruhpJCb5FPiKBNYTFwsiAqJqgfLXO673AcjAkQ/xyz
`protect END_PROTECTED
