`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lJSMp0673nbNRs7E4W9COMSvgSIRSGttTPSZ+eE6QRYgVZWsieglL6WmsuokvFt5
l6yxb8fgR0CCqTsCBhRArI5q3gxFzPOj+jWyqMMgR76ywtZiHv/fyEC5hR4863vp
wsJkPUjjPrem9xEunS33haETxbtd6VNmbscoLNvY19TA4qWO4fabcfPTkoLXeGSg
I7FTPCztys5IhV3OrWnSGMDot2bjT7bxAraA8DU3Ct9iXhwkzOCf/3t/oiG14aN6
mSTmV+dmaGP2+BYCGwrHiKbyeRTepOB/iJoqabJWgPpPIGCXrcZUDerWE/v4ugAx
LH3Ag1o0v4TK6rkjZOHfhnIzu1M1SHgqXTRcFNKU8VJyQi5vsV+7F5FxPHzur3Zh
lPPuKhEcH5w67+t007pY9NmHYGoqxY0Bv9vqYSIv56+kUW0QRGdC4cOt1hM4fUZZ
C1BtgDZeQE1SPI9g3GVc18UmR9IpkKX3fC2C1dviY/ZMWR17lQWl7KlyGl0sSPZU
LC0IToPx+sCmTsEpHpryVxVwczpjMngYDIzHWZAPIB9OlUOGQOsP6QouXepAJ82s
ktLRFxohYmTeVyFjnY9un2IlFRzHbHq6xP3BiYoDR/VLTvK4oYZ+I44M5PP14T6r
+8KYTW+QHKzKtZCI7v5yIA==
`protect END_PROTECTED
