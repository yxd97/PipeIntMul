`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
74hZwrwkmMzfPvMWc/VqCo08/JMtmJX+5WBWnDGnO/GSD84oHMzNWYzfEDu1TPQZ
cEVMCifXiD/JIfdAbHd/D9JcnCTV3IPn78bqxwGB9o3HDYgcEVBL7cxFPZcddfVW
/irRuT1TtN28QcvIUZP59BfcWAXI2j/DJoP1iEre1JpuPmccGu3UrRmU66PtO/qD
AJWnauoqegRkhK72QSiUYQnbLUZ6FUa5a5KKExNJ/ulEgmzp8NsjuqxqYNxF5/Gw
X3WcP79wbZuAWbisT8x43+1AJIFihRMDHZe4s4E8aQYRlEIpjPPYPCNRoBsAdgwQ
44HHV35J7tvD03ZlkvIdzgRp2Rn6B3JOIQ9F9SYCLz4iKkUZXljJl1yikcMPd2uK
+hgOoYVROcpJtVHSh8cS+VygJspqDCgYYEenygNG6njnQOpP+r3w1c8Km8I7MiYH
QObKi8jUUf+tg8m4Xs0CGK4JjHrtVfgzjdGLWpaxQyMXs3O6BbZuhe/W6wUTKr/K
`protect END_PROTECTED
