`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUEFypOrcPdNUMC1zkNArX0mg2XvZ/cFK2YZZOWMt9KTswcE0aLEIL4XFKBlvVM4
7ow295K/sf9ZPFqRA8l6tWpqbDp8xDIBTZG96k/5Uq5Lf3vAUB8yE9JvyC55tONK
3icfb66b5YrexwB3qQZ55uKGBhtSoBxZxEq2EDDKUgLlWf/sAhUaqHquK/DKMLX8
ltg7MzKK6TJA546YaGUo9E0jbCNKiCoXgSeA5rd3ASn/i0GkJFms3MgyNabb1WKJ
NfC7W2VOJ2T/zCvy4NhMRcbgfRj0+dYE3XArFRpMsY2KI2LcpV0IbxECtB0fpmp/
T2dZGSGlfIA7E9KSNbAuo/j9DjpdwfNRGqD0R1yzlKYQpMi9qFDLDPOAR2ifzMGD
PlYD2ip5QFkV39xFIlJxvsY6rTNsjtRU2OrmnKLgWnI31DqW5NVbTl65aFb+AASQ
N+zcNKVjr/ZWk/ZmGDpBPLzwAE+Hz25BfPDmxgtSES0fa/vI9vwJTMRfjCXXy0PO
sn3vErmneDBvhWrlI5stwZ00AYYLqjSPu1WMM2gyMBEFrmoS6t/g0bLAs+GULbk+
GkixiWgQod/IZdbxc3FX2QP89LVWExcKFivoL8k0SR6yWn/zKOpGH88EVTGnNgpn
0EHvVeG8p8txdm323oL2kJT7qSvMhqsyEF34dMTetNDX/m48JFSC/tf5/NC7GO0d
bymIPjRfSEU9+3+ZBpewPSxZtSC/gFPoL8s/wY4XPyXxQZDLYCjEjxYIZqMYUcNt
RjvQWFy8nf+rRNqIkFkUzFGFKaT0/NG1MdrR3jc3m9aQV2nH84B3r4rqfdvXmfSH
krP4t6qOulwZfjsQhMm4s8Kt/2rVmZmreqwWk34uSv/nBTN4Oiz123NoTYgnRTtF
qcyZFJL4aAk7nHhcwE3PfHF3taF4lhGPZ7PCUoCn5W4dEMZjFn73CpgnQPWo3wlB
YD4+91BpJ8Z0Mit6kitUCYsdlxnXsPr0tSXez2JlzhE=
`protect END_PROTECTED
