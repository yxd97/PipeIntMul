`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z3gk9EdKbXC+Yp7awy0UQZ16m2CcBcYDaszhsifyFBzFkZe6JotQO/3Xd1u2PNwM
Kk1hdUHTUBgnvBYxOVcMh6nurEAw3uJhfiOFG6Fz/2zWQI28WoDy/PpKaVYmQRUh
QPvkwRmR6geCwqfvnDPnYhG15xjNdPyOUddBX8WKLpaK2/bmBMGXAUO44KKKMhRt
Xa070DtFzhwOFNnb4K7eRY8nyjZn35UO2SV760R2Kq2DGWhPdu+u3FCYyDlLYMe8
Siw2Hii5qAjkvU2xtpMo5SwwUbjwIGAUbK1PpU+HBFawx6gTr4WwSJ9E0aNtqS85
Y5DjafdVvZOgL8O4E02GNCR1b4U2au3YS0RlZarHYupuDuSszxjslj2EIx6oI9Xu
hXVW2sN1Mn5wZhMmF66riCOJhtqbC3Is/dLu927+6RUmJ8O5F7DpC1zyIhp9VF1j
eI8Iy7xRmZue5EsNILmop57FP0kzFWQTeSD87zWwoun0oU7u7ojHqLc1SnVzyHgx
YE4sGqKqpNjSJySiaq72vHCa3imWm0MsjXA2jWohqUALxF5AF/i0RUAEEK5LZoBA
RRPpQEtzWi+xyDmln1VaScZN/Lpz3bhHPvABS3Hr4hDkkCGGJdtA1JslJNOCwgny
JqY3iI1vLT4j1EhCCGWAkecyrKZU0pN1Op2Czs2T0i0=
`protect END_PROTECTED
