`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VO+VMluzEiXCug6Dpwac+EsJS93NU2fi+PuW96vUWhGb0GPhHpkaKAgow9o55BfU
z1O8sUDMCh1OF6NSC6CfMp47goUjC4Gk6/v7CDUyML4WZMsXjF23wQ1kxT+u0QVd
aLG6tvq32t6J0mJoqKnYznKs1Fa1Xvc8XKQ+311+pxcDZRcUbK9sRJm2NysY8ifM
bJnTPOMLQzqMz8+TmI4s4u1UtFmew4rBdhPiGSIt59K3kQL2bHuWMIKXdoYTYrBW
MmSAWW+xiHulToV96mqWag==
`protect END_PROTECTED
