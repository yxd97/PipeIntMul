`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pbeD4DPl8cwIgBxsZIRpbBsGNDLvIWLSVs+9CBOHhyS+xP73YndvhEiJL8Lr4dgQ
Fm6sFnQ6iIGd5M/BVILtskNO34gL6/jQubAMbPXcBS98+QRf0qTxldQj2psTWENJ
Www0CB4aLtxlTx6dJ69Hyz0qb91v1tHrnWEFCR4ZoOSXpjHXOWVAoxYTxu6QIgRq
7ua2wuuiUGj0c7RZHTTqmxn2sipSU8Z1GWuvHlgJv3ZAt0j9gb0+nyR5c4BOU5SJ
`protect END_PROTECTED
