`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TX1w01/30aOhE45s3pHnbSORYElTiAlg/7phbJf4q7/aOhmSf1sfnJOk0B3WUQvd
iAQ31xK67Ua44igPKYODSkX3Jf+jGaXFFQSvR+LFDY3/PKO5u5xM4AoxUmVaBBTR
CsdeFOiR0k5oFaCqGwW7A+bKx0ZEHeAPq8q13RfUlO48f8Ni4khk+jYIgRL+MLGd
nDABUD9cGhai6fIOUAbtPzHSVrOC1VwzY26DS6QM5Ul1/YLlIvge7F5VtaWwhWHx
RUG6EgqvQmFvsZDBBUSHevxP+iGv3eEZeTxlX29vXHLZ0mtalaw9TKEnMGHRKP3F
2S9cU7YewyVQS0Vitqu9CM4z++6QgfGzdgwyFz9xbg9r70V2izaTJaV36x2DqqS7
7jklJs3QQIWGPS9pjEjbWJe/xZfHOuFu+XtP7udSIcv4T7MLanmLOnfv1yI+QEKL
Iw+JmD6VnWsi5ewub5km9emkEctoHe8aq+HZruQMhC0W/WpnPSnMn6cEA1lIwT4C
8kreqNt0zF2Yf5yEwOMdJuENBPi/BE9Mn91bA9hOczdRtsO4cH+HWiIsddmkZnA+
PGcc2e7QPwbv/oRiBB9udEEAUdC2zeH0HbhP+Rtthn4OSO4uSqFk1sU/9XKE+QWw
GSGzH2KA2R4s69dcH4AJ1YviD6uSFupV1iyYNQcbfBqRvosCMrlOIEdIplJsXhrb
XeJxHLvN+AF7h3JUIJZa79w1Y+O+F2cvgVjVcSnFcw/LEdShkbhFvtkf2V+ucoaM
aO9JvOTi6rnBriRsw5XLb3ihBxbxrDR+i7QEk5GRQ1Tus8HfS9ig8OyQu0Cw/q9d
Ry8b8I5u7jf4Ng+8EO8NzW/RG4giky2LpLEDzNzabWp55pfMaUKkGar9ZWMuSGpm
FSoKBLcrMrX5ujoERYCAeOX9HtVaPKVaxiBo4o+trLkbCTpPA7ND3azHMEo/8/GB
zU6t0/HaA+2njoTwaf3+MFf92/pogZ2SyvNwaancavTFOLD6vI1htLsv6xFAyK7B
rPZjkeJ5SWXJcG5s8WgB68CuoosyCGqLuy8l8JpKF9LDKmZf3D39Vuys/zZQPD6K
OtzBnRo8Ibkcz1WBvJ87nKONydVZdM0AoZed4GE1ks+2jCUNVx0WUzD/2/l4ESmG
zH2BIdJJfvFobJ/EXYSeXIhP7TSEFOfUd33I4c2RmkCWYsDl9lSzpc1oFWUqYifk
sVYwQTzxI9QLZ1nbFbaOYLuqLYfM1eF5wfsZNUAj3C/sInnyq014/CTHbF5G2LdI
pb2ND+CEttM1RC5SmE8uPyXEeOQgnqbV4vb+XKv8kLYnUZVYQ4p6zRGIslatJhzB
07ulmkrXaRwbhFaM9lAovPHJLqX0uZ/WJIbWFozoqnT+TbvvKFJJwGsgtIE+1Wxp
pa+vfiYiTyfR0c98re0O6McaSPYR4hxQFS0G6lFpVEToWOH2ltlyDpfcmO6tFagw
qVjs3dvKTwJ7iKs3hRB/VN1LBJ2XOWftOtoS3bYt2lyJMdfJdTIrLG0POvMfa1Hi
Pv9Z7n76DZ7CgWCRdnkaMsoHNUMzEZin7MtU6Vct8pjyHcM6K/7BEFm5iO4IXCzU
uTFW6yZ0jer4AgUSaudc83vG9AGhxALqvPchD7vC4nik9l9tVmOSYA+Ee95sXHQX
V8mSOI3SSftNPKxwMEK9iIgG/JmbgmjMXie+Z3+FEFxTGAnnEV93EpemV4ngdB8B
3X8sKwrR58ZcCCYNA664YgCRoMIct50B1Ztb0ZWAiQi6/SYWfMV3Lu/utpP7siKL
R3yb0kGb9iJleJmgNq+ItFkFvuEfKAT8S5rXSU5VKFX460BDnQ3FfbXBrYbgWkCa
askGrcqooLBVSaAYf+5Fznd2EMXdidRKn5bU4QcukiAVv9hW8Eqv+fQGRS97W+pE
ygeIefaiNoMnMqWIw8QrWcLquJMU0YMFYQ6ULZbmQlcto8nn6kOU7PlmfdpUfRPo
hS/hBvJ5Q7GsMIxEzjvcuhEfgVKcgiONakedKO54eBKqu+y/f4XZo6WXForLVRsB
4VKqxf0W783S5XeVZ73rZe8PXGmaxlOJauWXr7qEfBDwcBjAhY7ZEuSi4FK/uQwF
Cjx0mlJijloR8AjuM+xXVV/fgygHCDPUXI2TCPztn8vEISxiN2xWByILwqqQfO2r
Up7a54vwai7QLDXify3D/icCs2iMyQ4ZVCQFeys+kmcmeWmBPp/NzVPKD9PVLDGC
wwVoj7I+nXtpMVBBPXrskGE7I9fJOTa1eXcPQLWqAZtez5Hp0FpvUl62vF91gPKz
v5AC3oFMuw0lfNKMOiTShXy8EN87zp8pT3PTM9vr4heh4goDgWeoVxBuSrwOu/SM
zwQddFn1xl67sIxOQKpu+HyJCeknTUkZAPyo16/XRhDsEJUU+PxpGRb9EfY/eGVt
kmHSLVrVh+gbWpRVyG+fdvBykgL9V4zuWg4BRSYkny4uVpz3cr0VEY3mk+3TYEoT
5Joi7gE6qrTn6zdQ2FqhStxHDmEV/W7jRAdqm0G+/laslrlpVK4BCDZON6PoFqUz
Kdm+heXTeZ2YPmqlkToL6yc/IeVbEfaK8YPI7A4CDoDTp4ErD18y/MUJS68Ek6Ez
xiu2y62bw9SqqGFcqQp4YOA+pPuxA3Tgzn0PPkWSG6Gv24PKotcKpiMY1vMyTYYa
4vQkrsdHUVvjeykJ8ExxKuYvrZpw3ouN6l/fDCOmDRAoz756xL1DMyGxPpHZbbcU
N8k0w0U6M3USTgFuLwrmyy1bguDIz3L9gO2Bmvan06e5hDlNaggZPzr0NQOd1rZh
V4bMR8KnytsX1tWpi7P23kDgRT9phsVO2M1Xt61+jhPXeppw5vR9lLpuemXeqG4X
UEJ4G3rplQD6GNZ0iU9z3tES+MxJyDAgM9jO0We0vax86wTGFtAGiMSVUSRhHe3f
PpBWmC2kMZw1HhFdLJqCN5v2g5ugzgbkAkFECYnm7cWQCHrxKuy3n6jzOxr0p1Ui
m8f5wZJEI/dDMgsMKQ+G3++FmrpfIkZuyHlTd4XxL4uAG+wiekiSZLMxpJJnfDxC
DOFdrbaGRuV8ytpupS2AwsUdLgNW+k1EdobBD4lllHZV9IrWVSvpkxVWYL1JRfwu
ODGCn3XuISqTgu2p12skWlG+llr+r+cpQtkfknktATseu/PDrcb0BcBo+QUpSK92
Mb+UD4mlPwXeWLxBG21ubdBFO0/SzA2EneS1hp3L8Yyo0Boa9e+Cc7D7vi4zCe+C
1uDanA7F9L4Sxvk47Iy9vcl191hMdMhNTxeSTWvUw3HED+ykiyHUA1KbRaUp+8Y7
HyeXx2JuMvnqhtlCmgKolR2c0iYudqGgZZFqEf9G6azLs5YRvEDQPqwW4+c83zib
NLhacTX/rcxxObd3Bx23BWA4pgYptQKtfPmTfh7BWV0cWa0e1f/+582v7QaRfgq+
JYhY1zG4Fc3utMSRWZA3R4lW+QL3556mQ/Xams/pyw/4U+98p7gumjRrWDFhUVAv
5+7WkjyZAB3vcy5gxQnzwucAZpGxOlSyG+owOkfrg3j2H6xW5uCwmtNnTTpsUG4l
pyWfQd/HPCvo8r2jM9k86ACsZNUVI7aOb76G9FJ7G9k5CtLaymlO5iiJ93OwHgxU
JZwsl5kHa25xMoVs/QOnofvmVjm+LRr1+RFCuERMb+98+RMPBUxDNqn8O07igGnG
tWbP9WWJYBSj9/5Opz4UqC+o0xgE94V6/NtriTZM1TVq5myv+19rEawKMNv6LfpM
7/rbRGspkPlUVfJ+R094OQukDhhfi0jdHzEvx2+l/h8wK2pJJHlQ0Knmb0uDlU13
gs69ViG5FDs5OW7Xo5GHTLNOPFVZmmvw/6FUMnEyW73pucNcdKUZ8CQcSHhPf2kp
Cco3yXq0FBRcctrg7XLET8wVwLYQTRcrS9ttgl879lSbUJe+Vl82UtSa/LflPwtG
9WwtSmWJolDMWhnPW7gv+H4pnCb8DNxcwra99f/qw4SKlaUMXpL0HEdvpCkXCknK
wO2YWuLnW1VgiqCC1e6UQK3mBl4OOSfhj93lp0w5Fgy2v2A8YPtpR0GEQUg6b7O2
MjqLkf/beQdDL0f19NKES9C/97B2Vdbd+6g7QR/l/BjT3jnK1JmHoR3e5JZvDG7O
qSPmomEwAnTCHrXOSOOJYLKnywOS/VHszf3Pm1eDUJKkTF29//mclV8WQGgnykXT
CMDUSqkSTsiOE3jTNSmpkeCzHBKVCWvLOT6ZvXfu36whKjr4r3qZZmdn/7MRmUzv
r+TqvaX/QA/0I86hVm6mlWQDpJ0gRr9aKRd/fA23qR4WBUiy+4dwZpLkrYPvG/Qx
30ED74UQXF0Trd0ST8IiIf4Tw1CZt0f0GIqegw/cOYaPt4Pbwpu5801xeW0mTnri
sZJRryzm3ZLZoEGuwku2CROK/APGc+qYZCeT7KXVjMv+94oi3emXwP4nkJxQYm6e
eYd8re1mNxNzoLj/suxnhMmz9UvUA94mJoZAOEhLSiCZJOPH7TFqQvwShR5JBBgx
u7dyKvGk1VzFK/NSLzuF7QwYJnjc3zc3TKgAU21wTUtBZZGkkhHnATPlX9pUwl1F
gHILbLsjt3O6DnB7kjlQfw3SPkqj30pLinDAChe3JsuYi0kpOswbUoWJyWA89PIF
COgGMDFL5BvoRi3i7vlvLQ/QuQ/DNONMLbHeZ3CZuEeuwG3C9kTVuX7bbmxfqjgO
KDzTH8p2/8MoP6BeBJ3Sog==
`protect END_PROTECTED
