`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXmkVmRI/hFJoEV0BJWzNRi8lktfflHFomZ2tWstYEhclLiTAwrvbkiNrjeJ6MEE
0YGHDvbTtzCUzc6/9YaKHIQ0jokRBJtqVT1WNDznMXTiUWBRS/Ag6bgI1H2phLR/
yzeI/LFb26Gs/N8BNoSWoJYjHlvZo++lQ8ntvnb6Buao0AsUby/VJ05OYXDXRibN
zkOLSrWnb7cp4U6bonydYP7UEwhx6swc0XW5F+Kpf6dVLC1dETFwmSH0FAL6VB63
7K8EfWxrgP4bBqTLJhWmp3Qv3s8y+8bi7RwAzMVkI7PsARFbpX00p8lffR8Q7qsl
qR54N+2xjwAdOAMQlPfdnOQ7UBQ9cTwi+GMxZH4qm/sEzG/zJTRUzXDjVDiepl6Y
q0tNEqX8oWnX3e84VQerx9gqxiRliV+TIiq6TG8tqSgG0dmHMvIZt4uD/KeBkpIB
`protect END_PROTECTED
