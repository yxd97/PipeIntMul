`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEVx/Egcmiv7p3LQzeVSJpLQ14yuiuEbG8zOWvcb3cySbglrf5PUyeqgTiR3L5o8
roHIKSOEGCZeC7plsMIn2kQpISr41/5cpntX8Uh7/IBiLQ4y1HLwYqSJYjz7Zfwl
shBcwII9ik0OVHuCpcf1AqJj72WiUrKQJoxgMH5FHZ8QIo6LkNbJEmEjSI42E5xI
O4aJmOyoQeKxOq31V1/4Ov1KNUTAxlnVHp2YAEj4dExOHWVkMAUgtgBYkE2vzwMM
QZrFGwHt3JOa+1uIx31QAt9sZ8szAp9hK8T9O5NubOAfaDVZvjlnQiEW6fcowCRS
U4FfWleDiFR0vXw0v0Fy8/HGHJdndtXR/MGi4wp5BYUtIAQWN/JIbbQn/iORL/Pk
qZeRTNpk4yxUkots6WzrFdqSvSeAylRytwmYdq65nFIl+a0TrmQXl802vKZ8OzOn
YTE/9kJJSPbBktsJ91SjeZslJ8+VrSSZxC4I76UhD01981C/RgaCyRUaJJAjLSmK
2UlLtlUcENRyrbFhKZo6Gjl+g9cV+TtscxDSJl8gvwHZbiRV/UZXl1EAiooD8c9K
XPcDczmaTBf1hVU7bdaBpcI5+/IAzDA7i7qqD0hB76A2Dy9MKSBQbKK6HkZ7abi5
9IyDLJdppbEiQOmC24r3JxwlDg+2R0a/21SPz2rtMfI3QCJlCY+/RxmaHfgdW34Z
x6ovGjsRbIPFMzlfPmZsskYStHrjFsHEl8HlYRiE5fFnWGXclf8c30ztaRgDfKqU
fL1x9+V3kPszhFEruz/CEKj5Glf3Zv1u3JLQ2vxwwNGp3I/PLSX5mEwk+jNgZXbB
Nwjzjx/QbYXs0v5m559/oDtFA7ymnCOi7Bf9rGa1NVYCDV7NFspErQ8t7oJlFsrk
d+tMwUXQ5G7PtszinXtORpChp4kOLudpXvCPCmntcB9tTLJ4rFZF24sC7cS5wcIm
pzaFS60NtRWS5GZwgMGk7A==
`protect END_PROTECTED
