`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNKdMzxfx0c7iEXXX1eR1MBHaJwovMXZQiPQYertG2FIY19r6zpbj/SIMJZLqmxD
Ys65Cyo6F9u1lTJdpoCBOSxSmr5q6oLsiBCMiDemNRk6SBHzXgPtT8vobHOF5Mfr
tH6+9rEhXunvn1mIx20MxjiJvpJAxmMiADTGNMov2Q551HGceDh21GJQBTMaaf2n
rOAYMmmpvM9ERgTs2+mdCiACLz7MEk/aaYiLi358qBpEWvHnkJJ55a38cloB0gDS
YpAxag91QtyuHl/tcGTDb2RYguccbXniREZBSWQI/S+R0BIm9QvCr84WtgaqE02K
xb6RbNy+rrjHdkPBnDuZZgiBz04ALxINJtMaUGrqtzvq6gQPu1uSKCox+RTyBbAS
k8BHhdSadqQgyKBmr2gFxsJkk9YrFszdbwTU5v9TUqoetXEbCdK6RyWFXpEm+J+v
CkouYNXwLvGNE4fydmsCh3Ej/CJJ455QQ2xRJEsM8L6LwW0+jV6ALtKruOYnUTSO
IiDBBIU9Mf+kIfqjnMOI7hBOUSDTk21NkCxkKtTgecRXoK7M0gjEN31xu/ReZYyd
bmEDickwyzB090mMBEibfvRvd2V1Z5UvmksXzOZiSjD/aAE8nV1N07vwRbYQPqaB
kzINbaru+Rjy83tAtsuK3wv60DZtXZj9YLPl1immHSu+MyZ2XoDQutTdQ/gnVBSM
nCSLV/NIpJxAusJtuwwT46Fp+eiGbWIrv5VE8hHH+V19mY7DMqw1UTTAnqaKkTg5
9n2fEj+fxepDfTLuPPehuNJC/Koi8EpzGNgQ21/PdCcJWsmXcheXy+6r/iHdnq2G
E2BIsi1Y7svm5nRE6NEwyICsXKSWtm22rJk4uSnlwI5hoaDsO8q5UkaHHmA1Ls6z
rUNVw1wdDB4V6NG7APhbYd6+cBR7BUWAEIVMhrdLNMxnVgqy23S6CvvI28T1WEWO
`protect END_PROTECTED
