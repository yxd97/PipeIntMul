`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdevSfrHYSnIvK4Wn8LgcBvSWtIHkiTDQhHyWKBGVlifEjIFHPtKcQNgS8J+FqiJ
D8Ay0m4+uGJiPiRhJr+UKgISPvGO9mYY92dWxryPiVbf+hbgMrUSeIUxFgw7DoDc
ZZmdELx5jHrRSvu1cCmcqfolEiQEMnqL1s0W2Xoify2XAXnM1Aig61Jd96FjD4p1
wVZizTnUR0Qche0W0fg8KiRRQ5msOgWqdUAJMUbeTAGJehgL7S3CImVOImT+TvQB
C9mtQML4p9YQggDBGJ8UNGM2yTDzSAGfuTtBHextKMreTysQ01fOqf9YVKR34nza
C4xe8HI1AB7cxMDpsc6y3zFmvo+KNUE62GheowyLIlJwo5/WWGVH2egeYoPusv8K
H+Ld+rjOGZDMVFXzQdKWusCUTLLwEO9RfGhWGN2hljfBnsBOgtUWlGiZl2oX4U5p
jV9LsSB6zKtcskCn+FZ62VuNWSDlwLhrDg89hQ5faz1UdjVTQh89ogVNvHtXmqxr
UeCzvLioR0+uxlJBX2RYJr0WIe0SwYB+bOMoMAN/iQ00qB8j/DnosK7K2j7ohU5L
3yxGzroTy/uHTCks/D0Atx/d9UFtaqdJL/hz433aKVTDSpdbTSAFvIAxltMKgftE
TbPYUnGpNK5+yKJf4+ZMHqiwQiqd5GvgI/r/u+QNYD+k+h/5IBn/J+KpXCQm9P8i
WVyX4y/8GwjwBXMnGC+T09B2S3pLIiV4ljKs45jV5nMxAG2oJ/s9U1ZYFBscsVJ2
BOr+uVeHeLplm4Y9/zW96q51earshDnkdM5AKxXfOhlGkjSCBr6KSuG3HVb1O94P
gTlTldMoUi5EmW9z7DaTfu/AupvphJs3LfIsq8KS7lwyGex98EUQ0as7ClkeEKoI
FgzEpvCgCS+Zh1Nwp/0TvuYXvdSfO8leUj3XFsM6OCNIhTvuAgPiztzlRauK4ilN
Oa1pUj6y2P2gqVGcIOwGtJ/Lie2crlEnJv69V6nAdIkNoxbEGkNRfNFCAMIgXvXF
QDGAaCtYBYbnp/FjP/oEosOWvSxaWsTpFW00d5pDdzmG14T6CR0aNJ6cb/7tS59y
cDVJ3DQALrmMZuHNBrdMQo3Wou3BSlWzJkOkPneEnqF8FIA5Ks8oprNZkHqaPdQe
QZgWpznUfw8MiEIdJM+34kBpbGqGb+tcVfSx+GPor3Y46UKHwkkXhYxNdzBmwo+k
H6LAzEeTU4SS1f+Xd2ODXulRd3ly8+YccKjbEiqx/5xeDBivexV3POo3EkMOp3bq
ze56yoOQNWLiV1S7e/GPekw9NFEbpQ+nAM50a4Hc4+mbYm+k+f+/c62v1dsaa+AW
z3RCt4VAJl42ITqNR85hWp0UlK1DL0Jph80BMpcHJSwYSRqhuLsRBb/FM9UDer0j
xlpq54HM3dTxUfaaTxFkKeAo0DBkHHNusraNJjUS8E19KQZiu8Ag45DDcX9zLe/d
c/AmNibAQo9MPcIEk5Sreipo2he8KS8pf5PkYSQaKSZr6u6Sxi+45WX938AQRx/J
i/WEq2XslhjcTB41p+PRh2coUM3d2VmE1BrHAYFwNq4nD0N/Il3NfqTpFPzx0TcY
MrvCoeXER4LrqDUi5FEeem5XKgRNdiU7duYDgVbYVes3RHyczdKuQ46OmhYrbjRC
eymunRlgoMKxqm0L6zGOXks4wc/+p5Uu6h7NJxnICnAvoRIwO6fE/m6gxbvXJkGs
KKG0RBssgmjXsbl/ZpwvnxgqhzKFn8zK5a4FHMV6obo2DdWHloLL07YOppWwQ3f6
wam212Pglz4BJsbJ6v3MZKs5z/HkXnlKNwqKOssPKjhXbVBTyDoQB/4JbqJSIYes
A1PHSsPJjm4qsiRA4oKKj5ye2TcoAV1/kFUcNzcphPSFGx8Vnp5Ab4YdoXeSZrZn
1w0iMA+Ol24S+DaUa/SIo1PHm5QiGF6+PPWpxbYNjC5kKVtPntzWWB6c7CCyk54i
12UsDcnq/Lff6XeZdjxNkEx8Ntl3M/J+Yqb671yo4qsMaa8UFDpEbRYRwxBtOeWp
cwB2pLc9OnSDIZz2qbDQitv52HtDyQ8llfj/1ZPprOeGWAoz976dXYj3E5mnXXk7
+33sGBd2sC8T0pJxiZ4TybxPAa4GLjfvLYzM/v88PvjOGfRo4KUfvjakinfkbWau
xXyRwcuwZl/L0vi+1KDCnLGT1lXauJo4byIVBto43XHbGYtw+IX4xj02EIv1tBnd
xe3/4F185WMJdiBWim2Q5CNohprIRvMCamsrMFb5T05IsGNoGQ4qMCM2tqY/rJW1
s5h3MwabWzq/SZp57QUj+29+PZHfmmCBiI0oBjGu3FNp4E5Xp+T9y7lI1Kemtnaj
tRU6WCj04ywTz0ohxd9K0RBaCZvyUReiMZD0WtNxhzWG3F9/ilA4GCDiYTD1hIO2
bmO4s5A+a76Bwplppj/fK7mvpaQNv+TolrsRO+sT59naH7swCXdMSJw7e6qd1+IX
hB3AMf75T/7zg127rz6Rox1MwfESQNOpZZmCuUajMi9hpOiEPYjPCFUqwQY03Zpo
HKj3Hl6EAY+BB2IqPIJ+VvbYBr+LsH5ak5mg+oM1YbW0a9iKn5CehvV9Fr5zIUpw
7wQI6S1IKurrz8gJAOVNno5vk9zjUm36/jiTx2KVGEn0yG4J44ehv5kuIdwtxSWA
tA4pt2xNDT/KriDU1QiGtQyEPq9q9Wi8mI93n3PuWnKOJaJaAaOnSAWWKvroumw2
pPQJHR7s/QxbmZ6jntK9W0Z3bfjbJv9UHqmXrNZBRz5bSR6issa+vQdBbEPgUUvo
2YT7roZ9x7d3IDacuJrFbqHmayDnP2YbNlQqfQfRXGNH975fEJ6o0qBTcSJRY3gh
rt27AzMBRsODCSzVsGL2j8AxRiCLxlFddv9ySBKEc3rq5LWpwZqlBbl1OpRfOs7w
Yc7yA1QhZ7VCuXnuvXS3/jkhEs3c0tr/jDjgDOKa/jOHa308pxFVNwgq39r+6lKa
qo66APK2nOsBmbSbDE3AlDnvgA1zGgoMYOIgVH/XOzLnRWYtzHI4sgJgmpU7xM2M
FJQPfZ7mZgVENZd2HyNO9BXPUTx21jGiz4mztzuUdx266xv5JYbnlGkYmFD2RPmY
1CtEKXQia+mVUhic5KQ3xisULGA0CnkNjQOeNEM3BQo9KQAYVTXHKLyjFfXM9OyF
vyzmtf81+Ye32Cgjd9SNYghD6nkm1j3W4VjHZt8EKNK9HSJO1xOFulBaUoe+9p7N
5RLmrLloaXRiaWSy6uEumDUjn7EA8TfJaowkWs4icEpPEgU0ECqBHo/LUth1a8JR
GhFNvzCTQ2e0vr5m2lMKxqgsuULi4Bz31o2beDMNkMrqS8t0syw1/tShKqFOpxiX
S+ouwyv2VZtjMitcFLEkZkd/1BoTGv7GK6NNiZaa1dM/VMnNZml/ASVGPE46/Jhf
dlI7gWolmQDxugWOF/yp7E1uRscKjShy10nL7WnoUJjdGisxT56pIC8GP2yt0VXV
+dtf7DfChvdmjn5xwOAaKt/4rgWlN5fr6/PuMkUSXIJU5rHCUeDFi7OcdUh4i/nv
1wgWVzu01d5CE6X/1p86HPiaknLyqOAnS3zy7LzEvDZD3YYFqGUCB1LRXdMnpOX0
e+xZshGPBjZvrf0TbOofYrfNJOsANTt7Cdn0yM3CP3zkH3x7ETURLqJi7wBEt8tV
JWCsUX8CWUfn3UPXmG5OiiscZ8bHoQi5AfuXO72enrnIeckam2A9lXX9i6hExVeG
l/AQPwEE/Z+bIwCq1SdvdnQR1P/EJ5f1nW/2ID3LDNsy5nugin6x9HuD75eTD8ra
z78Ck1ZW1rPakE2bRUJ2rgvc83OMX9EcX0Gz0W/XjN7olxJ/XeKpl2ZbcIizxg0f
rRFA4xqXXtdZl45q7+7V5ddtl2RpvdTWTonp7UN9KHTpms+5J4XCbYHahy0AHVsG
syTZSUidkyd8tYUYILSR/W/3viBTX3+PGF8ofkGmmZ0ZmWi0k1cwjMIuP/6sMFBS
EZl323BowreW5ERZOqCvwznxUM22o9YeXebg/emYFKV1eESnBI4OHqqJpF3CoXWT
izr5krSGTv2NRYN4qkQvIU3lDXy75/Xiq69JyQR7ztpvMyal++SOtC39FTHS0JTY
E7dFCElzP7xLXhcw9jZwM7oyIMj/jWzDD+8RdILer51GRolREpRh54f4ZJ9uiRoK
9sN0GMOySdIfuG1Pj2K72mO6TqTDUEX4PilhrHLIgHtr8qpBHdbP4i1IbwiMOU6n
bAeuh65iiwGqP2GzqwfCTKnrlwOtojYSJEBIw2KP8VppPsQ3l4nfaFVP0/wGJnh4
CUb3cHGbZjaqvOqo2nQab/CMUkqHkBwrg8Em8nAGuM8gAGbz6jdWOtaubg/ZZgFp
hZ/fsTmoqAi1TSQaDZBn3KW5h2oCY6kdSoY1FZGlyZn7W4adxtsAD1kmXrl+8GJM
pTICg6XagbppqzoIxzoSFGgPEPo4G8tAJmdT7NseDbyPFNM4juMMIGNuLYDyrDTF
wpntOVXVKDLXY+fIq+9qhXmbclaVT/xaFMyB8SxvhlVj5lV6T5oq5FnPcqQQF9LO
Ro7oDkCIKmM3+3GoLgYLJQgiHVrtg5Zfhe3PtvupQijNynyD/aJ2vZINqkiscaH+
vAWD9ov/eko4oR4x00bDnnvE2WN5nSewIQG4VABjGFQec39MG4jTsCBcl4DdWq2W
CZRotOeTVlbWwcn/jhlJmASSC+H5Tu2lBthBTLUtuLPymIsb+ElZw+DJqlH7hfTb
Ndy+96bkYQjUhscTs/rwIyQErAatyFjiWo6KBGveTxcnDegKVDK50GsXctMCYxS0
NH906iM4nIwkF/Eq7HxLAq2fDQUvA6+tox1zqxvvwJ9MPZg1Nls1AoFQkc0tUcnN
ak46HJDsknA2OSUqHVJww0U8//O/RQoofDM3B12d1JxtwlqGKsaS7oH2iHRW7ci5
jpGPdDZAfiw+m/C7RUfMTuvpubBAapBkAjDoSMZ55+ittifft9+25ycrIeYoKBEa
Krx5N0Cc2zGxmEMQS3kGFg+xRUEVtFAxfeVySPYbDj7g6u6uXB5KiYgf4TxBduE3
Ae3C8/vjKf+0xtoksqBNBaH/ebhWjrL/3rd3B2WC4PnZPdmuzaBIviwBEdrYNEKJ
GqvPIxwuBoNbJwi6Vxke5gCFNC4Lz+Ty6ThIvDmaMEaAMpjYipUMb5tZB/RxsZvt
WEuvIYz+pgYTzvuAJBH+2mOpUQtE+F57unC6P61laEWfEgs47NHDDryHK2IdxsE4
rSO2SWUt5sNbz+ngYUhnKeXMZn60OUfmyuWKFixspbENP8bdIp/lXAQpJNYu0neg
WephNQyNNHjYLfW/nyhI3GKvYFqtK5GrckTm5kjDqGdaONr6aOI4UcZjUH+hSlNU
yPX3eZlMDibrV3QXEnUIHmgMgEn8Xlng1ok4s1PFdSEAJn5ls8Sz7RgVWRAYIzfY
t56186NVBv3FlTF7OfOgFXKpCsUHVWNc9QrNGBrOjkJSU/KLYa00jEW+Im6WhBmz
ZaNQdkwNP+kENdbjstV2tO0HEmjnHmMUtHdFq/UlSXu9C6fbmBUWSDOXIHG5DG6p
OWrEuuYGspquGfRLLuu6SCeM5dXo8CtDXF6gQm97rHfurOm20/fPZerO62Ovv/qv
HLLTsFF7Wxy1tjAjsDtSVDy2oE2SLxVdIHvaS28UgcNWyJy2/2m/r1ba8HBbSzSo
uPLKXQmAAkYkEiN2Dsg09IVFFd1oyxFk1x4TT3nGOZ3uNmVbam5YKsZl8oliKktM
vCWcOHETH/2fXKwf0+00MT8S65yYmwpSvDx1QkH2H14tgeBV0BLAvaARl/j4TkSR
Rij5nJ4I6hLNNm7ozB4OBafkSndzEK/XpP5fYqNfuq543TtKMeAtdFqxv8mhOCWR
6lCHjChJZnNatilT8TpGuKIIKB+ecJG0uxQJK5IwMmNJOL1JnB9z8366lAEV7cXV
/pRxe4XFKemGq7h3cTIOHzAid4x0QCbFByUCuVwieL+YcNnapv7czBOPUK5SRc3h
kjHwbekUsj5JYmhnYrdH9y+xQ+zw6G68hH0PZbO2kRMvTbrVyWq8ENpuzXwdoDls
Pn9b6n5eUBo1U8LGvrssQ5MUeHEw87ChsAwj2kIJVGGT7QgEsyz1HUv5Up/J48AC
8jrLWZap4IwyeOXUCzPOZQrNhnPnZU9My8qV1VzMllgcyd/UXCShXjbyT75M7/dt
DJM/dJh2Lutg61dhgUGsvln1rXRD/c4FE+93VwuaTXVOwkJ7sEijtx8xCv9c7MFb
slOTg+TxLEbyQtwCXqkWG1V8w6OKXprBZTn+fLcpwzRgsvYF9IWWYKYTcZRJkTso
eK57hj9DxMfEPjEi8HQiYcuvq8eV/GIpxJMdhDShrMS/Kod2+S+jyhFtuMTf5Lrj
kKhz9IchcAJ86Jbn52l3FnkS9wNJnEu071ld67G1eDUsajFGJcYh77jFAfprMolQ
p7Pw986pth1muutyFoctZmfQAp/SNyRvrjdq9zyfTfys9aJZLdAErU7i2MxtlfxE
xlQcw5ySUIfegRLg6r+1B/fEgIGbvqsN+nC6BQnTC7aMrIjsPTaODk4ii201g5LW
wPYZejd168PpLPUiJYHQemTyXTJ6j80T/X5BYVs8wNva1PUUhvh1yWVdcrV0DklP
G7y6PJgteDrKIfmrPBCWOfLPlA6UYnubUfDFkuRNZpXEswq5wbsMq8dsnWYok50t
TrbAWdWcOj4lh2ULRjRDefA0utyOH8fkj19gfwdf9fYBpxogy7C2Y0QZ4GcR5Wq8
BxYmbmScOAAHGsuzobMa24FOjZiMt6aWw5kgho8xNbpQG06fE0JH8V/x2ELeBfLg
gUXcmE/30iH5b1CtMh9DYdNOvvfoA79NXA7/PjZg6Poq5tVdg2u/Ke5OUuegTMy1
1Kt5xWEOojRjafkb5YdGZly62Ma2xRsdbcx/KJ2D9oOOCjSp3fFZS8o/sO8yMsyM
jOZ+MpJO17BpI2gEHF2Zt08MydmiJDsvSQjDpx7Oj/B932vWfvL9vVEddfLsSdN0
3bgri7tlLT7IQY6JmiPBRWb9pHSm657xtIfeBhM9uUMSXO/XqlkxDl4Ah9WJEGbF
AIxAsvj4IOurKOUUCMkb3BRbTniOl7DcM/y7KIQJYVA6aeIqxyyrNtSLISj4D9vm
ppdm2cRqvOk5tj7N5w6H0Sk6qxczlhXfpI9JksVh9eIRW8jPbqoYiCQYkcn8W9UJ
ty5kHPy/ScwyWM9T5HivnqLfa6tmvUmcAmjoCPtYsypR0yp8liUwqldnled+gh78
Rm83vZ812JAf469PiwMYXugefogSBEXiW0UYJjytTx+by/23kW3gU0y62qPcNlvO
kxNIPmzlK7jfiQgZrlsd+nTMNu6Pvjn/3A5Jq2lvEf4TDeyjxTMhNhv5lp3/7EQq
E0ZBBxsPl5k30kwg2KueCYVS//m3EeiHbPjxsdexT9kevOXuveyKeHsdBuSEHj8q
Vm3jPFb9NXUziIQz9uwoTbRcbV+Ye+tCimGGP1a2+tk8Y2PYY7oQpsR/2yy+WDTZ
BzRXTdvPuJPGhqhBzaaIvTk97LWI9YRzYvTmdtFoo/lJpj1Q9EIPBFYWKbg9rCc9
wCIA3ivViuoC+qr9/usSr2ycX2Gc7o+zHyupERO61SElJKz+wJomdq27RH0yvNuS
87xUy6bbw/bZtvbFqQzakh6ioF2Mst1VIj7puMguWel7IFBlxePED7a2OO8WThuS
PJRoeUtwJrqnSKCBgH5V4b7ICB+XfjYh86eEkjc+TB8KVGrfiBvHdWKUcGxMhvgO
TBneli3pMHtNV5rh6JTwsEQAvGw+9Z8nrK2mHgiXt1hyY5W3DxEIhp/sLySRMiDo
L2+LMdyPj96B85qw3BQNaNowZPHOC/fzDPYj6EgcZxEKUdvX0iOHNdx5WSgeQysE
aajbGLPtr03NxzHsriSnKFCusAWtQDcnxX1chRbZiEo11NExwLaQY1CF5VfTgKV6
UnsJW5Spek5PRLTGRV9F9Y7xxOAzQDnq9+BLKEGIEH39SdWRUf+u8eQWluBQD2g7
rFSihR8/PsmUiXB0Qng497oZbdjWERdqPArNnje8pCqYve3bHLa0tsyk9lnrpSrg
hYgWIF5ozD0+XT+WeeVIrV6bxkPw66YYfK/Isu/nLo1yxChaiFwpL9JhITptPvxe
rm3v+cYOK9uWB5l0l2RydT70XU6Rr9pOJ4AoY1d+oYszMINFhR9HB0JZAh5Qzm4Y
CngGOVmZqUCCXXRjEvW5K/3vhNfp/yryiCgEybO05XZUIzuN6G5t49nbFMjJDWK3
gntYw1gaYXLbearFapZHRD71te0sJ3YDTkShFtGGOlkPM/mn+Oht6amWoXSMmnA/
SfdXl65AuHK7M0eIDGbsH6+GdXqpe2tQV/Mf2DdDphy1cBDTOby0vW/Nq+nsEjaN
7DYjSQPhEDIxnS0bNxm/g+4ELjB6tI4KaL1s+ur9zHgle+JuZ5SB1eO3mi9Gf0kV
ZUpyPwCKEZXQVfG/EGVCvXKx6lbazww8+MQxz//T25xoVcgjSBHW9XEo64h4GCvQ
Yot5nTXPcL6q9tq+bpaHK1G1Dkpeeb0CAFT/EF4UCNZejf81Yb7Epu+YpRTjOsp2
pC4XofvDWL5SyTrLiniAJnX0IVHgh9o2foPhPnntZXpGHIWimtBBeCKQMjqEVkkk
CeklzhOhvOy2pFJgwTn5LmNf6YDEL5xhDJ5YWx6W0o3YMHswLeVO89yxafXcGWv7
kpmP5AXcNxA3g/PvuxfUo/laetJA3F9op73YWo/iHBkLEYj23GQPiVAIhYWbmNT0
32OjjxJnMvEeTsrjuqmTv+j84lZo16jZ6fHjTefAgt/25rXh+UTKA4T4nIBdj39z
pZXVMrTIKuuXehiouzXhVRh/W1cl1IFnuYNzkCkXxDJrnvmT9id/QLARApUrNoYZ
HwC/2CF/Dpdoedp0EqxDJDArs5k+SvzQ4zerWuTHF616ioZszMGznwu4BcklNcw0
itQY/gPoWbNUuaxRxZGvNOBuDhhDiDwAFg6XcDUgvSX02WJyRee6bU65lyN0zW3S
YdXCoGrFu7CqEyvOxVE9h05UNCuIFTrFFw8UVqYUbsSaTHhXyIQKyk/OqWtwF/5Z
ooMdB3FAXX8X3JvpWbJ6g8Qq5pFk488/ruHV0BKDYX4LMMIBR3dW0pKXyYdBGeHu
nrsXWXsZz2uhazqlCLGqoL+ApKx2/K9BTCJiOBxg6+f2is3MeeddxkepGAsN/CGs
FApEoLGfqQ4Q2QMYrS+n3rvRVMHpsBv2QRkwSPmQ1kAfUWabnZLUgDrnUjr6fAwe
Cc78p27lXXZAIsC58RLpaPC4fxDNkf7B2KLYuPpbYb4xHWnJVIWYZ0SSri9BOZDA
yeX/rE4HAhpvfGHcFngEz9nH9RDGvj1I1QE6hCqkiD4zXWT0cOUuUN8UONRDG6yq
wR7D1dk6qJWZUJAfC8kgjnVQaa7CrKQILJcs995OA2JR0imxIseMughZXzTh0ENh
talw3yUNjyMKGtkIg/kAB2kiW3PTX6Rj61bxAeNxsJcwXYUib25Fh7gvBXG08gpR
LQC5F4mUXY+IbN4HD8nQPzAxc5NwYHNZoeHO1UItuBg7s2oX51WXsax581pVZyP4
Z5xa2AR/BhSEubDaWwd7f3ZjgqKErWST+5CA4ioJck9IxPfEGY5KLsP1CKRKDS7e
VJKX035IL1ALW3wQDG5PmMXFCz9IV9YEILHr8/BYCFmHC10ydzbzwcACtAKoDBV5
C4P1CTrG08QJC45TkPkPUsapX8CtuzL32jSwfWuJqTPAOgFR6Pp9pZn+0B0/Q6Yp
mqGPrBDyYoiRX7YaLArRMyx/UN6PJHHm2U15ajj+qkRbmtLFWnkgxoUmR1k2I1my
ScCuLB47ayeQoPH+0YlVnKU5BofBd8jCtCCb6Ls0yVcnfRa+arUSHVfoMj9t61bX
X0BGWvgQyB64vMsIE5LbRdFv+64c6rIazWoeuT5bYKPDnOByUvnUpEx8hnyQAiM9
NOTsJmKJaHY3oX9xLZa17w9ECvnDkIOC99xvPQIkGOXpZ6jdEDIqyeOM85IjlZd7
Bw4R7HRm2Q4G2x1sXQCRaQZE0T73fVzXFtxF/tryfJWQsRzSXPy40su44wm58ipg
I/4Ab9QIwCMoKkKcgN/BTzn4bnTgN5+AU/adxITbFgNwRf8s1rUCA5zUpn1yGoJJ
jqtVoDiydtmkIDPfCNhojeXgC/SjgvzggxTuS/JE4sxOH+NoPvEtB745koRc2oA4
FYpxP/zloP0jfl2KTp+a0/SJVNlbqmnsdoJZScK+3vszu0UpsDFTC0DiE9eNm9ES
SFufWpuoIFruOiwFm/3GBfN5w7wadDVsBBm+M6a065olZLiLSQWMcCF2cmPCmxqD
2T8kVcWYFJ2CAuo9kkggludbitpo21BFNIyIp1jD0jftEmzer39WIuAQ5A6oBv1h
KIj7i2YZBSRYj6CqW7CEgHNpG3sQadGtLVLRwdJEpmZwWFpaSGvfTzXfBWdi1/Al
J1EoGoX7/PDPLnDfh5cM2TJelrsLplsai87X4nB5ZbsuCE3vo39hmfhbTbAvQiaU
7GiN4Tz45NSnVfSJd4u/Fqdh3+lW2SGqiSddcoCmemYjRTuMF7evW9ezr65bIMOe
Z2Vj1Ja81R9m1PCXMkI01CLT5NZOJFMZ38fVEN3GP8ZE8ZYs9IKTo5aZ7uE0lJik
S8wnICUaEvpNdCDLyr8nWIFle0sh6x5VYdFBDhJ8hWAGaq96T/NkajjYTaaLW4Pv
7hY0Jwb+hI9nQivaLPLD3k7ubzVQ/80r6OMt4+JSL9xr9yUCpJysAIn2Kjx8d/as
EI/dLVVD8C267AxQyq/uVkjWPAtmFLCEuppNhjAxeNnLlqSklP3jeclwduJsZobm
Jyjsj7shwzQO5Qcrc9htwYnTgwYHjEk0Xxv5RsB9m+9Fb5yfffAChpstK03J3XVm
GlGqV3ytueRRuTX+6ZaLxLlwC1Tnvbl7rDT0x+vnyEo0El79CxGy8yPTRxIHtlHJ
1MwlxLigwypUQyAX9ZYkC/b0TaiVb0//2GuZl6LY4dukrJXxA1HfgCmTxEQ2xBYo
gkaI0AuNtFnNXMNiZp8jkgLGkKoSt0KDuP89HllM2cabcxyo+vGMDfZaK2wphpGG
/IDzzuohtx+zUyoiEJTsE9fsWVAj0D6tXTNsJObWLrTVI9vs0MdR7gFdn4cxPnk5
hKdvD6rmNP87RU92aEENXT5cWoDPZdMKj7p4NiZ8v8WZxXSlgWkNNgItYF5Bucyz
TU+FJyWZyHhwLlhIgto7UPrA8aPP5TWKxaP+kEBPZR/CUJSCCJZ1G7bsPu5tPt+J
unlaQ1t2NsXve/6599YPlutc/NYoMMrMuxAhksv2jDgHfflDrEb4tnzboe6BxEIK
jZhnNBeaXF1Ju9bW68a+paryMVupSmJQQB69VUi9yKPmWncz5+RYojwfDI0RM39U
K7kGPQF0cz5xj1wP7xXI6U12FrDOF2zFgMddyutWQGkMbr8kxkAZwR40NcCQw5Yl
cCfkMsUenMwr/6lrLtWGyp2rrEc7EHNXGRjwM45YgZy9pVlp4lAcexi9Z1Z7l1Ao
UugsgJASixPhTP9z+xn3bULhp/UsnKQSWo2y1nbSyDgyWgyep9Pjmk3koiHX+GV6
J7uex+Vfve8vi2LWEFHIu5XTckt5cJdvf5ZoCIJQc1YX5Wh8cGNfN48v88xKj+hf
Xl53mM5OQrGuUJasxiLuuYbNxO7AwXbtF82Mdxc7zhQVS3XWgBzo0GXkEv+LxtUl
EsxY7u8eJmqAmFFtIouxeyWPs5NAG59/FLYafKiay8YTgk4l3Txa4Mk/wF9x68Zp
baVzFogadHXTIPc4RDgQUMYfRLZSNtBF/rbahnR6t8oS+jByiOXT4hwKfNUOqBxh
LmCIPpmy3XPUbwQ2/M3f2r0taPAzC9YtIcIYopweqhvG3euJVPOcu4zwW5UMxum+
j14G8fyP6E0KVwOZiRDS78sHprA3qcaVKt/jKV7AO4SRzxZDiV1TPCvtkL/AeXkQ
bbmZm/5TAPQhU17ZzWGU7quT9tShgexACIVvFvKf35qg2l993nXAplGBGtRel29p
3ERTwbVdRHVIpVW/bxnMCqvvhvgxjjIbM89qx+guRJ+HSAfwVxvTVPoh6D/rjGu+
7K60glrfyaxQ037eVnHVCZrzjFAcQRcxXLp7WhyaeENKgHu+UoIYI7if9oVXiJT4
Mb4+bRUU5eBCdS136lg0SdKL1jM7sePy0HV+jaRzLtWEPYVPR9QzYYhCb/YK4DLE
hQiFL7vSY7pld4YWcXoynhJKTH4zNi/XHT4BqNZSOYTjnxooi0iOX/hfv7u258I3
c37q4NNBvU4xxZaZL+7e1ULWAAHaBAa2vyWrwQO7wYRs1ckMRbRbC1FqLBlzfB4K
7KLp8Z7AH/EVb0JICru1dmadJ8j4PPVwhAeWW+H+f1o2d4NnWXHoN6/qpAYBWiuu
hxzNMZQmVSYPNEU0TCZcVus30Ylt5r78yjDVMuFXz8fVN036O/KLRTO11D2j/cW1
nJbeE+YEOJR4wJqisNwcxC8PX3/3n9RXEaSVjP2tgUxAhtk26p2XfdOhUGciBATX
tdwOoDBNw1scRBQ05IMqlRuCSO+fCZl30dHEY1UuxqH+2/A/EpVx8n5bs0HOY3hG
VAC2Uh9lz4aZMKSCftomCcDgbyKuGXA+syq+nDa4J92TaOAIYwOZ2fVPCF6I5O3u
NqQVf2s8762R78xaoGmdw/O5AMwgKUyl5W5jk+oOezAAnA4378IbVbEPTJGEEXxf
ZcrDv5HKL4vS0MilF5CfzTwncgwuFnhJfDNvJ1egtUyZkKcryRN5u3Sk5Ozz+Yc5
JlLFFsPoNJ4syma28NiBegKQmTF4eomij+Nyyq2zC3kZyyOFXEx+/gy5KfqwXaFN
fesI0dbLmZ2N/CrOfKMEtOIa8XufFxQAfZsCCEzUla+lcwHTRVjxV0ZWyOyNgS4K
PSVrjbyFBMGFku4o1fmNJoOW05Qd9iF/XObX6sZ+I+cLI3hc22IFZFWrCkkzttND
57vZWzC3CNdE7tMWCIiLdqod2VjIEQzyihYjD7x3cIE1TNGG7hL9jeB1oROmQlln
BwmEa8ru9Octxd/EpcZYNkc8YXfYc6hqmmMpda+xW5UKR5cYwSUzU9yFtj/NmulF
BFvqJPEXV2wsCAZ8fU59hZm/BifFNrgdNbd/3p/ndsobKW/fOQuMPkhUrfjk9ZoQ
mubh89PziZkMM46Rv5Yc9W9Vw+3ftCFr4xdaZ8yuXcy+d6JC/fxEAU4M+2n7U/um
YZNKwiBBxT0TFMDz4RSEJlwENUVbg2dEL6/M9NJUfrk3GkpHmCatqorKVhXf1sKH
BgtcAY392La/9NJPt+tiRUjH/kmfbtBGvDYOuJ5qrgUKdmQYhgOFdXVeGliAHSWl
hHwYjPbfkAB4VaOsmDjBu0nLhp4sAzvpR2nseR8Y7pqdJgUcaU+R/znKJaH8fPfx
/4kzRnTODXCoHeRq+p93KyZVQVqNAAtuNP5ezhjjKbQtsos38aLxyvmpftc34YEF
UxNS/CLFPz8xjoZleEx/iACusIQ0B+2bEr0sMs2yu+CjpjK8E1plSdjoJPxhX8aZ
rFyYxcSfRx0hCrTUxUddOGIY6CDPXUURDDcQGnod0sWBrpOpAXO6RTgmJR3MJzsg
/m8YMMi92xPuIvq1wSWbrrizplSuEjHI0y/tQPX2fOVGbAb7RPyyZ9jfqpqPsf1I
GRGAMzUnUxW10bJilU1x7XTPYIdR5nVn6efhr+kccUuUrBEZ6M1c0PEbWIN6KM0K
JPNfkn44CxBikOBOYSJTL8QgC5cDtvfFni7A4KifBl1oWERVCRVuVtkqCsTDsSUL
W7VwbZ3utGeUmZ6SrQV3yLvluso5wK0jSvt6SOA7aTj9mmetowMBvsORhI1J0Z7X
sHm4pwChK5rAcaGdhRvX1sQ2Jck9b2cc+4oi9cYlLpLwOEh5R+bi1LwjLXdLO0fw
wkRbjdqe0Guu680WfanplLWxU3HN2w2sx9L1l8ZUp5zy+z6ARqkJgH7UF2I0e7RK
w1JzDRJfXZMJQnKiCY3kwOhOfUHxuikUyFCR5gjAG+yAOV7mExJaPSupsrrSDIEh
785QQP/EbCbgeSlreB9nDX1MoAYnQOyRWVMaOgQXgCFSGf+9PSoFEPAfByKHUjr4
SQbO8PDSqx6Z84ewjfYL1CjtOJhB75YNbOLaICrjflyoxOC8JAcMjNk5credc2gP
s8n4mebk/YLqwPjmDAD3hRnlU3/dON142hiaI/BjFN5+bwsjbWFKuFODECD7GLjb
jnXT8X3sm0q2Hv+vGmXrxtU3iRjqsxFpQL71LS2JzoWNLbhvQwOPucelTHwCHJVp
+6r2JPhRIXA/VRjwu461mLoJeqck6goHQBMY4TjBtrv/4CtE8WgSQ+vSfL2GDseP
o4FY9PxIwACl8czBPGIAe6T9trCm+uIa2Rn1DT0UEMTJ6rwWcVzoS3GUYcot3LWV
Po9925lovRwU2ClwqbZrdShivvh83b3CE+u7aMkNHpeInN2peWtRZOTpQWvecST4
nDFPifrWR/RCuKG3zxPa0vXkwNYJzXlHA/uBTcy1EHB+Eo6QFqWYeeA+01jCHj+0
wSGsr5wCvYQKbEy0HBOjF+s5Fn9VO5ONCQfRyg6A8ruy/cXTNIdTphZzG7ZHpOhB
d+1puruWoO6aW5VVena3z1dHlqnsSCwWHhq4T7r9HFCv0AxaLRy3+37azlR5uakO
Ah7Vm2VjHYPTF8EbEMj5O+w0dW+9vfJCMIf2vlz66BnWr0k9uo4X2EA1s25dYUM2
8wSqPAFeooG7AFgVoFwUrzN9cqy8vgcvh1El8HgkT2o9uyfvNVXGgvy8fYHS2oWM
CvJaPwzQjC2laixCnS8MSCwvyCV0vo34bBz1h2Jd0R24E57u8dIZoKFSwvASXn22
zg87s1ioEvYG/pW5DGHBx1M3qwtO1oDn23KDGEG7aTaBmUpeVnEVQXnQgafajBeS
5TYiB7LDxtkVnF302fZxBUhqsd+2EFo/XHvEvNqp2e/FJtnYnZbQ7SzualE5O5LB
BvwQ3I5rSNw+9SCXTf8um9fJ0uUqZ6xCOsQyHmQ7c9BLZC/9r1VUdnhUFPyUN7iY
hJiwgJBpPAhH8k7AmXjwPqiqNVrnHwcQD56ND5qPW3JwmBYGRtJvLNrzOCRM8aSl
CHaQI9sXLrnVohZJpwJl3GlymJ2Mo+xNvOLz6x+I18COG/PI+zpsZX3lpDKT45kt
40WT7GxCqwmjjetNbbMGJe3VkhzjTB6IybIRbw3Hvr+1AH6viLrPi3o/9BvSI1qD
4oKeScJXZ/oHSYA+r4iJDYlNqfBg88U8nHuK7AztrBWIHbVZ5fsVh3jY3J99pDCT
HrwCf5oPiedtET9U7edfRjLcXOhdedNq7Evb8QNYevMOHyxfM8RQYfmfCS0JfhBf
ytnVlWj9ZnbAhD+sGDuy2fq469WCH318MZhn80+GFgXsZgttjnh/E7iDvZRJrIBq
VdqHUcACbXDhX/OWagSebz7hCyc8jkzOLn+LGegjlZ4M3AGnI/P9ZH23Bh0+X3w9
I8aSDk8vqDuRRMi/dRZClX/JeJmpihYh6F+9GCMIKMQz3/dxQ2Ns0ORYnnoOCOUr
b1b+pP0D6k1fNZf4joLpJEV2NBqfgvrx+u/j5D0YDGRXvXtc+rk2l0U4kerYNuf2
F861EwjnVjJi2+niT/VtIRicszfv/c8dgEW56cUDrEq8D118Q+k8EpcC7+oNOpPi
dLZwrqMeUgvlmjsN5xK617hYamN8hpc5PTXoX38ZCMW5/4ibe4tTXoAU1WjS7VgO
MlcHm15CipEVPF/pYaaydxdLzL4AD8EVVPxhxhv7Swb5jrRIl4Eu5soTgD+pYqNv
DdTR40M5AWGEHhuDm9bXfXiclWqmL6USLRwe+ZS1V6W+Xycb12XI3wSpl0I0cqSX
E1BG9VQyMhy0hmIXsQTxXKGmGEqqhnVGNgS4lZpEuYgvMDvZ6vjJf6/K4vxyP7ex
lQpejOetL+KOkBIlRyypS4VNZnBMAwNBgeKOBBQtQNFpjsD2539NaE99yIsuLy9s
c4QhKjLK5RGzSyyVU0dTVi7GlxWr2jdHGzr1zswHjv/L+PfT8jb88DBfQVDYhtaw
/OH4gfUHw+eKJwUuSHG8TOlQw9tAdr4unNAWTwHs3lCebCnSDd+8BGBdKeeFf5F7
7RDwTlr8u/tHhaVXb5UaIQ3GNWgcMIWlcO9htHx0V9cYpbQhmbRFBaZUJ10LZhWh
Mw1dsgEkEFfn5T8Cn4mcSMs/A6GHKpUiXpzchGVFEyKt2W4XLswIgJf1xqWzoQqH
SpPyCAYUxv0EZqs6OXqTG/NGN8FFGpITds2FWXB5RmeoWjKQfEMw7BfQpvehq8zb
el7PY7e+/yJAY+pEmjUvPH4ePY4usScGE0FdXNHtKH9t5v1+hjD6k7hDRTeBVRTs
CSzrCDi5nmSNny/2RrKakhrpooc0PNY8coLfUmreRp1gvxpbQORv22tFXs0coYJb
ddKKPllEMLoflGypYLKrXvF6k+ZKxKOpM6WrfLgWgBblgQ+bC1LDeguWSL7kolSH
QIZO/ctgdjOiKCFpt9lTH9zxMPDnJMoTBURrqfQX/HXY2HmARXDpvv6zcNQWQrL4
bs69cXh1me6oXpEmOh1u/btDk0SfjkXYUqL5jSElJGRHmHr66dVC3iDeZx8HDCG2
FpOsjyq+Q1nDwzV6XuI3TGmyYhTaYyrY2r34e4aYZXR0qLjGdUMsq1OuIBEaytSV
RDQk9LY7J4wHvJvpdJTFFhb0oTq8mBPqUj4Zu0n1HRuzENRaLo32rfs49yfQVvyL
WZANwI0uVJdnxkLCiwQNzYhjkw9SFHr1vWtMVz0wRGDThhAEmnfrgwkT/gGJGTqu
fFzqMkEbUXlLqgyXdeaNgb5cyvkeNoDhXq6EZ6auQ0arVvSf4pErwZlotiNbTfsD
ndmAMHjcRIrmK2enUhlJp/i24KBa8Ip3HbDwt5jB7ODau7tyDCY54T4whP/4Zx5H
D0zDwgcW9Wbl4pJ/k/EeGbMniGePtQ2Z2p9ibK0Lw7QB12dUuiCDazNKS3t0LFYi
2BjDD7KVn99yZm/NpuCoZPbMuWfyoiGCz9fKHySmJEbTnb7wyVyKTLKsCS0CGsNK
s4VNefmprz3HH16iwiOxtWccvoHFEPWizDUev8chko8hpsi8Lu+RIq3WOR8fLkuB
lY26KrQGg2MJrKhg2c4tiRl4bfXf0Y9GAvGNYld7JI6SSNV3Koamn4MD1ZGJyXnF
1Yq2FZIFMzR+SFAqi2iOgZrH4T0OsMrj5+ekFZ525MxeyOCZUocB409JdckjcqdF
beU0tp7tVdK2xjEHtSyBzHuEkxhuN1iEmgA3ibMZGavcncaxv/J+hwsktFPd1zbD
5jghidHyquVn0sIHQrpyj+0OJCbQk4ilcNxHARFStKaTRbzLg/d2FzuA+QGRl9mY
RmLq4rYi1Y48TYo2KFr1OYC0WyH2SRzlCz/N497doldhuWxzlaEX3g2DxekaVEkX
YeQrAUO13kUT+HR1AKZxLp9tmMRr+oMUyddUYcdAKdN3FUwUkCODO8wYx2fWbEPg
XUjNvpOQKuZvz/wLLTNV5pz+SIaLdQu0yUwS3f2wqsvlxk6AizLYT7P1dLLp+La3
cF3z/Lel9yepirrdIZt7wVGsv1Al5fLijJnnVs+QW7HgBEg8VMprOG5LdbYxQktE
no7Cwqx2i2JdFKEKrq40Xf0u5vYzrlA6TERnonW2uS0bR1ZfdMLvvS7CXxkH7ihj
ldGcezvbEeV0T4S4TCLilmH1RxcCTxi7fwFdlDqsAtR3Urszy840RxAcl2NrEiWG
6IZhoNzi4duISNjVqgxzOuR4qfdknPjJOCDb3neViqs2iER66/LDiwGtqazm6D+y
V4ANR88xmH5F9rA1KzXlBt7OBr4NF5KP3VSF078TI4/lqfDz6o6pQfJJViO98Y01
wwN5yioaNXgWUf2mgYoO2TFDzB6Ug+76dVzR51blQLsqvkKJVQ9n8dfEWdi0mi51
SK39lsrYmkSDMT0LJofeNFyHCPnRB8/qvudFQYi5NYoeiqIWafb5B2DeRAeJtaAR
CGSNd5XvX4VDFEGV0/AqpYRygay287HcmV8BfS5iPH0S3+X810q77vsRDpXpCJlc
EBbh/Rz5Y6EadTbHRCkOjXUEbRPb5pGCaovfcVCp2+FTz1IKUGzZqUTJG6ouVJsF
L6NRcXru+C3tFAmREWksJDfS2FLvOEyCxcse472ItwMGCKVHPSSOCFCE6ZOKVZse
tmmvIlEo2CISXkgQbLg/5Mt9l0IUaGZmtsChuaXUY2x9M5wkuKVHWIipeEGT31Wi
ORGHy9bN9IjAwusoVsnGs55RMEU8hzq/4NH1rNM6Wa5Wica5SmgyD6Td12/S9La+
pU51CMdO2+Tw+0ypxST6HVJduTH5/FSjsxnWETlY2qlYErExuzTxTvI5cFY4y+V6
ilCRCbCHBmu5uM50Br5KqD2XEGorMc1WHB/Y5T9DOacvLBNlZgTXt4w8v8LTZPfD
UPLfL4qMZQY4Btm9gGRd9csXFWgLkFuDJRfJAv38Ny8kttxVJCVUu1PR2+BRoOCH
UE/3l7SFgZvGMyk7hHKtiHK1MFnUr6glgcBM6ukDLer4BFfNgkXkTsbwInSnik0o
wO/YH3qNsWLdtuX7uDUqz6QXSf5O+YxTbzqCPyPExPVLRvZ+zn/X4KX5RQo8Ox7W
VwfAMwGs0XA4TGg4GHmA4atJlhfnTOQNmHeBsOzL7vvNb+IIvaO6dsCUS77Y+jR0
80yZawcqFO6ApFU1TdzOGTBZmvhwXOlwsOpOPtpYK+Ij/EjeK9UOy1kfUNmJw371
17ID8wc73790HffNsfqO3UKTLs8z3+QSt4GR2zeJ0WWVxoLnbk0Fe+ldn/PcKPtO
0GMT/U577BN1iV2zHDknfjx/wLz/tOPZsQvnM2WRWp1aKAgUN+OzTLQBsH6O23YW
4u4+ay/nEHu07rgOOcCSozzt2VLdVYu59n3yNY/NRJr7/K2t8T+Kx6UOOsiYDOcf
+dLBNdxlq00IHvMVdktbRXA3Y2ALbOcaNCLx81ntVMNuWR8pxKtXrW63V0UV1qnM
FZ5IYNpEbYRQ3U2x1PBi+z3Z00x7bM3bJM4RuaUIGN7C8b13t8wn1KVcZMduWv5r
5Z4+rz+QkUTk0ARYgk9cwpVChKjaOVt+WoKBhz9M3X1LIqHI8IVMRYpsxabc93XY
lSIqhDG8hqzT9BGKhWEinpC/5JuFHJJH6Yl81u/oo3gobALpKfsaaVNKscYO8x3M
6pc3Dm7ACXSgso+tY7yCrzfgox2DcM1/6Aj5G5mg/wpmXk27sEiovPj0UU1cFK69
y8BRUV9QzRVYz6RsCOnHkI3V/jDNkBn1GQTekmJOnYKWd/0tdOtuiSMfKThdKdlh
ekfgzmcJ+7+WKlZcJMZtY1BJwoytIvyns5fk5f3ErN42JQ2IU0Y5oi4cH+RzjNay
xd1NLZN/r8QRe8eJT1aQhwfZWZ+q1NjhZ++20YP6ONfjaIQBxGuo4qIlNlorGaPe
Rgnmsl+exZ2AWReFRAHpTdy3Cb99lv682g7XLBEjjBU42PSaaynQY+RiMUsXt6oX
7TipR385zRIrRuRWLmItGwE0igmz7kXi+2hzBF2Dw1wiHu3hnJP7I+XL+7+IcWfu
j6xr4FJQW9xB8ZLAaSKwQPoEMkcPBO7lbiy+1p+UuD7k3tVZNip+1itxDTz+OUE3
4uYE5BZ2oISCEeObJRbGrms6E1bKMMzLF624QhsVkOdlI481WVZAtmgbxisRr238
uCbdFEY7kUQaPMxzmAjeO09sSl9pIGqyZ1uuPOBM47b8j96kuDT24bgBfe6u7TJe
xe8P+Eo40EsPRHXO6F1Rl9vgeZJNuDXYMbdpT0fJQRl2eXFcmqf4nGQ0vBmYmNE1
CjvxxGL+RpuMJ9KJTOG6YxnXlJ456Cc6WWGMpQBQxzk4GFq+np9RFAu4TuaNgsPk
Q2wOFUcYkes4VzykZmVAJ2XtUSc3BkuztmMyZW56EPqanRMZq+2EEBtSnmXCXJVA
0eDV0+1eli/luAaJUtKR6RpOXarku/1S1B3PVwOpLlvFNzv9wUDF31sVgeYsQF2H
VBIF59AjG0fYiHieQKUW9NPi9mXAuWT7AXpRwMPBQc3Cs+6cKqnmLd603DWhnbAv
UmKQq60M63xTzbI/s1KLiGXl+P2HUIKzMvzdvWkFw0jshf6JYYVFZXdLF78RBiuT
gpNHZobpAoOcQ8wHE6unnkslkIvexoaQLwGuvTcyEyHajOGMPWSOn/y9f/iUNz3O
0TXH6a1a876zlk8hIaMnTL6PLc9b30yqQ0JkDiKEPkB+A9CdIwNmWteC/yRmzNE/
Qg/MRrdzQwiILLcngxVFPhlvYvmt1bZo+Wb+Dda1B3MRxs31kFUKKWiqoioXq6YX
SpzosuaoFetLp0BMliQ02+sD4iOIiamcWujCAaC0QpkxGPYXcA/kpnz1AE8VHMiT
vLkEncld5vP1J5H0cJbXvXCrIIX761Yef64+57EBite2daDPcq58B6S1sjkrSpzt
V6h5zhyJrO90RiHJzymmMulgiJt2xAyaON0G+n/T59toHLsySpQ/2hMpwVxPutvM
DnOZKJCSejZ+i8YWCdinzBbTjqOgyDtGWzct42WutKU8mTGCCbCX6rvOvA0GI7vR
mEoUhMNWRmIamlrsFbeBFrWdP38Y3nPGJNEYna32zpgeFEtzzxyhi2GQQWtzxjNr
IddQTY1/eHhK4Srk5YhhiXopO1dPLo0luzojJUk22zwbbztiqUd/wA/i4qjp7TQq
YsWLUw+joZt81GIXJUTsq0VEFrSeLopKIn4eP4Un3Au4zA+xyO+2G17UR8py2YbN
wEXx+5heHRIydPELAvaWi+tpbC3IBIIIUtZphptGJ+91N1auIe+bOcR6Z0D1m2vQ
BEqcFXuabIjbeYT1CMAwTkX0M9kKTWJ2lnE6bk6KOHD+/JHoc9IBk5eS5wJtew/N
/uLssJQ1l1ddwcfyty3eSP2+v+OmQ47/wTWBsxrsd+CgygJ1ny0IbXegA2xfZsP7
sbf0gPOjYXF400NSErLo6va6K2PYLbufWWpUC2n+V9RYUWC+WshNO2YkhotEUb/h
Dd71+f8l9Ploq4aGH1F560JxKIp+6HeUpYBPG3AbwnbX3ChftA5eruZgLmKkJf1I
Bc2BoR2dTVKHsTf7zbi2b8Oyz+d9djHdAZlFVN2NlIKSMRFpqim21ilotlv2RdxX
14wHYosp7a/VvhUFoTAQAE8/vGE8Tc1qH5s0UiCsOknavjII+Gt+BG8GHhIoVAwu
TnvdnDfCKHz+7WF+pm4Q9/tcV5FL2aYFYCw0ucf62T9OcBskYCnIHKd+4KpKObgX
oWR0P0Tzmp7ifrmOfW51YnD9fbaO5AEETxZKvrSrd5UZEmJW+6tmrxSDbxBHQZGG
V3wUIfoZrB/f2n/rig6rm/mJvODSKd91YWt8e8TiFbkXApqn+NYaPlH1ojSvmZ7p
QPywffi9g4Hy/7ABBCjbIMDGcQHpCdd/WRCiwiUx/bQYUwC0rQENZZiseoIz2+q6
/Ddfly9DVIvd1K78Qhi/T0bsth+7BaV560oGuxOLnzMP3QL7QqCG9q+rWoU6VSH7
Uz090ryayjVCIMbREbRdULm9MIS45n3fG4IteogSKwp5yCuQgpWA3IXj++63E8mx
yGAtaXmG9lCdLyUHfXuPmq2J2YDpKuq62MfIo8gh2MEH5i9BZLfjOdV+A9EKtay1
iXC3MvoV5aP3rPQuXpG8xH4GYuK1zo7Kg/u80S8xWUTwleDJ5NTQGJhDALfGqCwp
v712dYlD/xWFt0YkZSzZpyCaJLZ37nQ2+XgsAyXqfjm7uhwfmYh+2c/eaAwVcnf1
h8JGjTQg6oWGsZcB8lJ4USwIRdj0CIkCUh6Tyb0eP7Oj3QUN9FeTU0gyOSN+uHLo
/b5aUcq9ajqPKbR2CV4bRkfRi7nHf5FPA8Zi+UgNrg4ibWDajbDiBgjt4GEpEfJg
mXMYSyhpV0ioz+JAAGt58NVF4IiHxnbOwEmaJllvUVBvdENWl6duOhxEWPVhWl8J
6SpUt2HtWjlSoj1uM7QhObZobMMtIvZjTIG5zvd6gnqnj+WVQBe2m/+Eijirp/QD
jqKtvljhdmYqY69QCgy5fQephiQD2mk4wR5Cn/0lKdewkAFbsT4wrLtbhGcYOmBK
DgL8lKgcRy8TQU4Tyv+BIbpA6RkZbAu5AFrtElXJfMCKEmWKJizrQ9RAldSdH2Us
aQdnzGV+tK3UYzeJc5ggJAKpvt3AWNCwpgXkbY3BTo/Lq+9ThGf/J7iJO1x8y8+8
meJG/IEzCoMpQjhO6wXLstNbD50WkEOgdGh6zLtNH/XTN5lkoAL9ZMCCowAxsiZY
aYI53YxD25b7qrtsW3PFCS1FfO48+adtRg8WfZBdf+pbzfOeQqWcDXVEc7nJAb78
fABYy9oCdLcivOI4FV6tMfSbB0gjFkF15vYNYW3jMgA+MC0dk+u766FnHPy6v+3+
V5syQUExZXSDgk6UCmyKhZXWb8esiCdKEt0by72hRy8b0yJ45AG7uI2jC7Hpl4Bi
snummvMkYvJ0VEH3eRYD1i6dXqqmsBV4lY9A+gqpE7+aIS5SdXtSohYQgYIynlEv
waTLst3iiW7VigEco+JqL7VAbQsteOYYS3KrfaGKpVJP5Jr8ZdmBsxMaHkNEPdyL
T1iEof+fhf5PexYcrA+Rj+CD6Zv0awpven3Ib8pTD8IDKeYeeBdPZnk22J9LLVk6
fw1mCUXPZBuA6Yl9ss7QiOwkp/cQTVrdm9/giaksaEQnvH5A8/9buXxuXjnDPl4K
3thjZxFvpBkj7S8Zpw59kbleEy9puJ2RlyMrg1RMqNBWycrDfTOi29i98Yc/VVhJ
eVLRfF1uPWb4Y4nPDfOFnmf6qW2i0T5b64brg5qfO+xQ7ZrPeRE9xEkiC7cJH1am
eryF3Qi0HB7yptRkCIGsVY83/LjxkYSLG/1+2nsnxZAb8LdnxdywcZ3XE9/jgbQ2
U4+6V5rhSsKLGBkAjwsP+Isy9qpj/uhPUogvOnqAsgxgTTDJfNhv8F0rR77sHkax
DY5ABeIS+gWVIdrVl1Uirfnm7er2FJySUmGI98tkDMGEoTdHqrF7hQ3jug/ZlhcL
OdXAIY9blBfr7EN9r8NJoiUV3HQ4rR7TYeC8PGUWyawxGpx5MxoEK/oNHajo4jtz
+ibrSvp1J6iPAnY3adAeWH5x1YtBi/hG7U83WFonopEgAWqj2+0e+B50ylQKVxap
qPk0qcx6KcGMIt7+NM7rQfons2ITRBCJjNxR9atVILNEgGBTAOhVTDNY4q0c32I+
zyoRUoU4WygwhP+dYwW1aQ7r3rLbj9U7zkS7+gRatX3nU66cqcsRBHhr+tZoAi8q
1H8o6bD3TSsPv0k/Ks+2RIoMsn6K4QmjG1smNYv+YbSyqmRNse+tf/gIrkP3kaH+
4KV8ptH7lghxI6WVNZAJwMmP5IhLoMgQFD2TkkwYdIUyBOSnmQlqs7zZFveL5GlL
/U2PnxyhYjquMNzz4Q3sodm2JxBM1qgUYWhMR9iaJsfJ4PzYWn8OSJhptMw2ZrKL
xyl6F/gAkvwGt8Xb0N+/IZwOpm7HJnbxl9iZuY7Lo5mR976y2FZ+OVmDRjzu3uXs
3gkXCwWHjWtFUXp6hTTpiT2xmOKKnFI+9vdNlVA3BNPQXSoaqXwkLkKgx9aET+bp
10vc7KG2kl6dLRyIJA8vQkwvHb19zPa6KDKdC9H4M5Wc8xtoYK3CGb+zklhJKBau
LeqoZtwTJDBsYoe4so56e5aSbJvVgeTIAm1G8ilxto5P4dNYEk3B1gQYAIofvbaq
4ofvK32jTRNf3K+HWhH25b42f0QwpEdi79mFyQt5unirFNA2sHK3xKfUFOY9rSkE
8g9d4ED6Py10T4lmyD5uC0Tm4koIbp2d58kYNbLCSeaZj34pNkDDnQ0mNgjiaMln
CKwN93bj71NrnKKcKooKNoJcPmxW+Uk1IHknMRQ0UreHGj6gZxbgbH0jMzFF76Kj
X3ZezYblxfjBMd18nUUiNAm5+dbItA0OWlEVRFbxvNXAGsRC7IoLFL1oPv7wJzzk
T+HVmpSCmR/Lqs4BqOCT1+BO+RbJvuSrHRn4K69G2HakjtXH1H6jtjKp+t57VfE6
Si4NjvVjn86LdLYAVVgKt38MvBXYC3f6B2S/1mDHkIDRTyj6YfBrFsRjsbHe1JMS
3d5tiS29cAxhnREkx5B86DLZ9pw6n12tKI0AzhqhXwQcIfKflpKKAkb3pMbNzP++
lHKsxbCYxqzULGZLjfErEmjuVxLhOHmM6q9dl0IBlJc4UMjP5PRTVOQP/lSxnqa8
HjBCyRabwMhVzoGO/xjG7q5cumxIxWHhMX/GY78QD69Loa7Z+KT7BDdeAT52S8M8
ZrSTSD1ZLusbDUylXwexZSI1yq5SYi3X0u59HWPP1ZDy87HxcVKPDL8g+pKv6iL7
I2HoV+yZNbOtQZ7fmbJywLCsIqdxeC+g6BnGu3n8O9cdNtU3kENwrkxRr7VvJnkL
pIXArAG/vkrRHNfLs1LBjWVSoNJIKhhQba6rHQLYD87N15co3pJqpNK6+68qc98J
G4c5/udKoSwlGJ7DNS0wMhcCv4OmFhW8gAC3wRQZi8QpkfNblwf3Whbr1w1TOjYm
ETsTg4TUROxLNTiP+/jnRz36GxvUqpQHfQHjJiqMho+uLvcwsqPxOj2W3+bn7wr6
ioLiPH66BrBWKHUIeYVccocrxUaSwRhTPQbclS9ZS7f26sec7HYamK69BB3p5s+s
cjSbnsAOvJOinN4sq1dkNM+Izc17aN+zaK8en7OxVk/KvL0PHlax+KWkXGFFaf52
7iOOs9Lza2F6/Qvajk3zfuSrRNx54Wti32mEYlh9w8Hl4tc1GtcaEdQvrtq+wwxa
zI3Ct7v+26mAkbx6aMxKtEByIt1cIA8QNT6G/xyzia6DYgYUx7JTTliXaAS6l86c
XOxP1Re4ENbHHPkvWfIDqQLUtNVFeSDvhrkLsNOqdP4cWUc1knJu7SXa3svgxZtH
6vWadDcsZWPUP0luq+dSBLhWj8tDWDo1mMSMN5Yd0ENBmsv1DMr3J9YyECsEUGOZ
GfeoKhomkeV4FpVfMFJSTu8UgTXtG6Nl5e24r6UBj97Qq5aj1G44djj8LkmcSgqs
XRL3wOGzGvLh3IHTQHDKHyQjz4qf/oGd2bRXr5/BbUydSGJ4dwHoh8lPROAUQMSE
O922nDSbwA/+WvfZbC3q4g2VllBdQTw7xajmOkyqS1w6KEFc4snzShY1IS91swIA
qQaXjRfQkh4xMHC8rD0KilZTbaWaR+ovLynrtWCuVTG6e8vD6YerGcAmfijSGeK1
QOZHvf+Qy2zrwXcxgphxEUaEBJsFU98geFTsVm25wIgFqiS9Ms1+HWgqNIOltd4I
K+Wmp05+/VV4Z2/tsyNP2ucwM5hUmP6Da9KVKpYKwkxBI+LNeoXSBs6O+jR/QIYE
ISfTfp5TFjJEIBFD95OpbxrjY2DWt5aJt9fhfIBOG7DPbGqM4H/FRtQa1V6NNcKX
4cjnK4EFdJz3ZEX76jDeI/D70OSsTyw07re79/j/Vu6jn9GS7Cl535bDvcgwAi+U
ZlfxpQ7rEQcQK7xk7Oy+GAbX04YFw9IIW+L6UE7T2CbBAX8xTjjDX/3bgeCLNeZQ
b2x1lgQ2X1CpLU+vcFTNlL1PLM2rKi7nz3J4z10ncQF7ceDkTpB5RQKaFLW/A/os
XvIR1MPgbTH6ugoPy+fF9NhlIcBIPEqVZuC30ZOOUphNAeCexUR3EBv8p5RBUlQy
Da67Ov4QXNl8EgYW+iDTt9R0mqnua78bbe5eBDUeg/ZLeWtd6TyqaUBdN+pxHFsQ
xrZqc//nONh7vRY6PTg5kPOmXGDF/D0mUSK+MurhKMclaVcgQz0HDBmGUdqikuob
MG4HfhklxQnGFbjtUUc49+YQa942+SpamAhjCmQCJbs1gwQ7rudRBGR5KfNHaw9e
vYzmMldN6G2fKKndKzL166x1WPremLb5QKZTK+hT+b0/GPi3WA1KD0/VDt3q3t/A
BZ72V0JuLU1tfm25PdMs0JPXl+W9oqVIGsHratwzOtSxvXhoEcPHjaV9ucsR3e4f
1YAxOha/YJY4Ijj2g/Z3wymfUQI+8EM6dSRu4kbQm7rmlkCIYHyHXdzW4lBWHbgR
9pTazq2ho51rxMLdjSs4RxKcEdnZh/uUvYfjpt2Wf1FUQH3grq1zCjvmBfw9jCAL
t/Q6NdI9qUjPmvE8f1h6rFnX13+cKiIgUaGDFZCjFNPA5Hs8kHaqcFUDN1NgzTy0
vcwc/2R8Jx1wOJH3+zZKeua80NKZVSUmBwrwWPddVIROpGMYZ3GCj4rRl+aG/Swc
cR3h6OCgmC+RjX0hdlg//SqOebWP7b9FS9ZNWGJ3q/eIXg9VZ1CrZA2a3/o2nURU
yvnE37RKEzIMMlotdDFAa4+yc8DFPVNc66UwjpmU/Srh8iRFid2l3HqanZv3iQJn
O/3CyZhWnNKFzG9Ynhj15B3oGfu9PHrdEVQHHryElvJ2mp5HIYWFikdkLBu2v9/U
AtepKu9qiSBPiqKTMonsK8KWYjCqKz2/yJJgXWKyAKNQpr4ociI2HaP5vLIs77+C
tzl9zo/z8ZldBb5Ie2GbjKGMbzvk6Lq+KHiTpns0/0aubk81TSN/C4odwXbNcJfA
jnTPiJM2ulvYIM2/ZIuAcGtq3wF4CCJO/QlztFIQFt8S9zFM2pB6HYfv2rKt5va/
VGDDy+p7nIf0Z9EACvUyx2ofaMjtb4U9jZ/qZBFAwf6rts4JqxQ7jUUnjhpVv/7/
RT90rEW7Yao4d2o/Pfmz/TWIrDk9SnnObvn96Fp3yY0IUPpVP/mYPW+pIFM0NDP1
FtOb7I/h+2XpR0zNrtKJgxpfmdOXuKDMjSAKqXeWRO1ep2fNhM5GM7sOWnpKrmTI
8wnTE/I/E5UpDE2k8kOxoK3YSOY8dc38rpRgx3CnzK/wks4GyUogfByO5YduR7EE
vigODSApr4Xdt/Etnx0Bssv1HpA6X723cHawxazqZlvXcZe43OsuDrQ3w83zBnFE
Ula4qsWS4oVrzNj/hbd1Bs4+MqGJDF0u9p0CwUt20pj8CACsXBYjgRmJCYApOhbI
KZYfn+mmLnuE6nl7rVZL/xLkMhQtViJLGaF7ijTWFYEnfdEEuWwvBHcBeAkVbd7/
eRzQVsjku1vpzYCAMFfNVD8rmfYrqVnGcyOlenfe0Oji4kJoCUi/O5gzBK5PrfRL
b7/4ZJ9QITlLSyjviLNQXHX8xQJJzGH7sT1W/UnY9e3L4o2XOO07LTiflZEgBuRB
t1ESUSEfcAx9IQokMoJqKmzmIQCvRo5x5lNCy+rXeGq+04TJSyCEU1a+HqWHwSOR
Y8uhNfkFdGSL8pa1BnOVTxRJGXRuSkFSu1JUuDIjTbfV01apEmqGucdKrr4aflUp
E9EHt6yTrIhi8kodu8V7dYUYQwsFU0xxaP1QachyWqXL/K/5sbWT8YFrFE+Ulpy2
OvZaV5Gv6r9nUstQa/HVf0KxSPQKL/ewSiptNgEst0sCClF9Mh5ev20GeYUgB4A8
q09CO8WmbMNXDb4HdwM+gA/3UOqSmBuKPRKzG+hhnBogFVQypELYd+9mpOG7wCPY
S+db1iBYILkFnXza0Vdb1igG+W+6q2T7nUwZgB2TW/iCta+3suXgI7cTfIIPRhfW
K0mqUMLsF5z75y8M6g5dpWT626TBcC059jmA+3BqWVshVwmJsjPNwphsJKII4HsW
fKcWZCm9Hhlyz/YJfGb3suAYu94edQ/4RcouK5Xi1OtNqvFbpGxCOEtwMoNCV/CL
2Z4LtZ/2M/UmLbfldreYmjUk1wdQqEsAJTLzsnp8NH63WPJ10CkqyRMnbKUZVvFE
utDDMYCW4ALcewshF4AgUQIlEfNaS9SQBgyac5m96oo1bF9YyoBMUoQkLGC2KPYt
FJrE3ZtdeIQJng/nYSW6J2rq2+uzKX49mYPeSERNJhILlcqiiIxpUNReYNwU9WoH
R9gXBG5WPnPy6aXUGzuvcbnre+ENLYTx/2VY1hUBI7Rf0B9ff1m5LU4f1X9xjdCe
x0buZzA7y4Tq1vIjdhSj7mnbswu1SJcmXYu17ATqXf00eWTIwMOCxD/Zre+9xoLZ
otHKfjyvAvsuHVcL08qvVbwugxN5EFZkvxVqQjCMaAf4Ul2v/LJemi3n3soRiwvi
IaW4WMVsHqButZwPYEZiD4nmxloA+dzeAJdWlp7xS+N5seY4VelSgWlAcqkNvS34
QB/+9WzvbUpBGf+IvOa6g1HI7AmIKSxx73ATDOrE3fATe1xddcNsBgO1IN5ciwUh
u1/nPSwPcucNTV8qeglKhmzdFxB4QHg8ATapaxxy3zJPnagPYbrpLlIutzMR4fC3
j3Su/q30RRk+CBjElM/zSZR7tqG5QLiSezsKRDPhd5d/ZnvBWtlDCXfvJ3mNWsNb
CRI3jZmvDWHncWf7pujA0YKDzBKnGYRbhzEkLb2Bpz/xmL0eqJiGIvjHif+xAgcA
5OMKWfxcVHo7bWFE2EwxVFPe7Cd8cgqSbb907TJ9zoxWm228/DnQzYsYlOOpMnOE
ic9Ti9A+leIgP037GYfMvBwEanbjmSU6g14RgQYWnP1BzNNy+nokwXzZ6+aJHq/4
KtnycODGeW4SMNDWySZVpK02xa0m4rZvz2ri3W/hcFGApVkvXsypPfCZHtY1IQ/C
NfQ0QkWzVQlqZKH5hveiAeVBKDyPwy4BLM9BxI/bS9uyIdRG6WMm64DcJySu3c+w
LtL19sDneUhJZwW+qQK3K7tUXcrwkAHlssa1NjXluLoVugAP1sRv8Uez+kAaOb9T
2RcLnz9PrpwJF03T8TVFVCFrxJgcjeqWevjQLJj6ReB/KSB3KM/3JmBvdq8PwEh0
VQj9byETYwm/Ly07CMJc0wEVzJK3c/N/ofP9f4MJ0uivFkUMowq9NXlLo1Nu66aR
Eq/czoE9aQVCXHWfYzHmnx/ii25xXZDHiHShcjKw+BD+7uJUB9xpxlyBmcupy9zO
JA2p2RPKF2xAknQErnrlFap2zHOJO36OVMZq/1KT+UxhVFYcMJ5JBSBf61+sMtIt
hVBtTpPa6aWGZbr7+TQ3OhtcsQLtqw49OBcAMzqAWTwvybPy0AklYXbbMyLyCh4l
bhuNWwP0HODcDImBIF3Kc06QRvuXppb/rIIZ3tXUBYIDxD7O4XMGVPnKC7iZWnJk
Ap2gqUpBswXQo7O6+DFAHtsj0Flb4b/i/jpn1QRZfLBgw+hj3mEZNTSbGDVxgT2v
6Icfn8cJxhYpXjk8cR8KmgAGrCX9T5TdEikG8xem6Wn2J8z8xzD1EC3WCGe3k32p
1D+sAiUgWdEMk30dx90CmWbD9L7/oVTfKfLjSFqfZwYHZrUno113midvAZeo4LOQ
tqNLLj4QtbXOUwbYIG6oBQe0yBUuPsF4xCkaaPlzXJJtXfTrC8apG6dw83GqSDqj
3KJUEJGW/g3BvCvAcqdi/YCdnonid3OlUnDAC15c6vRbiZfkJEdNLzNN9/BtIamn
W+3HfMG0UiO/5zwP/QwDys4smy+afXq59zYstflb5UeIporMXbbr2kd9Qm35nPe0
/A7lg5tH+rNaZURHpRlWMN2khnY4U44oD4Xf8IikEE+p8V3Pb8v32uLjBOPes2cY
DZYzlwcsHSSyk+kG5pc09iJdAxcENtwoF3ETNIEwnCWncVAoS19KcFSPZM5VZ06v
JrD5Nn1rrHFqh/MERzKM1TdalQvC1BiOW3EsPylLfPOTh4PjL4xhXf8WcQIIM/h+
B7hKduxU5GdMNG5ff3eYOvzviVhOBha/npc0ZldOpy8VGMMW0ah0lBaUWGqXQDnC
xWXaLCxip8oQH03Lu4V+ya0vuRcC/MV4i9bebd4ocErtNW+QrLMV1QhvIsMisFVx
LenZMOTqRvVVUKO2ShFCCYn+/xf1Oy7RUJaiy/LGevGMO5R/lur7a8KMy/QA2zY8
MzveBRZa1fVRbdIlCa9Hfkabl2zwHlDSpKel/ZWaWbB85oi8Dl9uC8LpFJKcSUbO
vft+q33vNmUNx5Q7DPbo93TMBeq1j9Jz+N7H7QmrBgpTBf1+6L9KT6OEf8666zaZ
jQzTtumnxQrPiNfy7X4kBHJuMLsGjH0RIkm4RbCLgRbHFcHe/nuzPd14nURV4ixu
pby7yxzKKbPOZsefFM1fOqawGG5RCEKS7+QAA2501Q3CIVxv9nWUChCRrr6w0It5
BXJPUJYmgokV7Q7NRipU8D/QezOHgGjcs+2QlV92mt4ACsku9QYy7KJitlYyTL69
hhn+N4v7qBHXJ1TuO0aU12ZA5eEgNPD+kr7MKvYd1MKXRYNWpncO/8EarLEhrYOQ
32MiefGqG8CBs35Dg5FReyCYs+9YGIi/q4MvX2OfO1qUXJjQO+R//42hHdy61Why
bwdkUcqRVqdeF2CISs8qkjeBxi92xIBIATwQ33efnl04qRY4FkQUItJnicVRzbUx
x6rcQK0zI3OFUCUi7iu6WHNm/eI5JAk3SkD1lcK5D52QdyWJKGvJGwv9qQ3Jod5w
4meTEWQzBw4OQ9Y6Q/lDVF3CZrs19iaYIr7kp1AwSC1NqLG3FBDcfAddRoqyP6Wp
FwwTkzHrYJAHMaP3DnwRacQY3ySuzaDxOG/yV2tzyziCEwOQJPflKDJHbkUgYjgv
MCF3jRxUuMFRtATg3r+REoRK9l3zB+bjvLuVfSE/8dvrvtlBk82g1j0ViIAyX8pd
+YJIPoBwiy2MRZrh86lXw2Xsz8XiSSgsK1ORpKQBhFJD08uioP76RfL9xyGqGA+R
ImFcILAW0yStXhHQgLwa4TDMP0HJ+YIfxycQvUnZg3CAJBQ2JgJN5vnAy1rieiFO
HtJm/nXs7w3RrHP0cWiV6JkNldu0tcoL/FOqLjxIr8T6t2e6K/tZXF/4B4LWKoiy
+3b6RvMXOR794M7IX2KIax7KFr0nZ9z2E+2iJwlEi/ftQiXkuJSSmCXWfb9+naan
AnMISPT/bucAVh5MayYoSq65yM9MCqx6eAXfDucdKtTLa2DA8/jLCVazXnFCXQ8M
265RPgYp1pTdPIb0hVmDnNBbi09ElMkKJgQbwrKAZQ7i+oVv5v1xiHWgrCLHA4ma
1QijNsIIqlz4qxdV//ufph/7OQP/ISEzFwEfRVEKWeKJU63dxYtOTPj7D41gR55t
hQhY+x+JOQXQ9+KEtOXcYqPsOFs1NGdQ6E7w7zsFHnfcp+yMmR1V/oP9K+4Sjxmc
zoJjOEshDZZ2mMQGqTJ7Zy73Wzz/tCMJZEGZV9jXRzXP0Y7N6X4hqdqlwddxUq7j
ZOZOoxdrn77MT9QTep/oR6FzFrc1/B5tycBy/bFVuoybHpfJ8NghT6bSbbLEwXzW
LQ3WqIO747/NuM5oMf/jkhLiIbxGRbzTO7phltdGRAAl6H+sSXA99K1gK79NqD3M
Jti8eE52EOvQwT5NsheI352ICNaMb6l9nJaGJvBcAyZelKes824WKYpee/uXAwiB
yYd9P3n+0HZ0la/9pzHJ4PHjtuHiLDTYi9iER1CvLTnirCr7zrLMWD1pjFGii++B
wLKfvVS4/at8fYsweLbkwsbRQ8GzLwbdChDVH7M92GnYvK4T+Cs2fLWp7e+OXrcZ
rMdDesJyZyev8g4RihjPg/MIU6Xc92CwXdrhMCBCGN6U5oPAYgPgLWm7q7zUKxip
y7Vr8tUf1WpS23oeExPlaA8DumAYOj4UKrj39UV24Brc0do6GQlITps2wryQ7tX1
0i64/3M4PMOhTj1T7vq9YGr7DyHFkQWW3MezPLDmLYB2IlZpfsLiIKyjmKTkHk6c
HvtVxZjEn8n+LrNi7Ovw5MMLltstv8ZNERRJIkAskavJ6BOswh/vq4SdDzxHndRl
laq7DGO0QldJKuuOi2HotI786M0Q1qvGM+fPPI+G/+jGc9hJ0BL5azhhDodOKdvD
x0/5j8yQHbsm8f2ih5nIew1Xp0SzlrJUqUpJevwn2a0QlKA/g/isNVGDohGQCr0T
qWmFOLAA24Hu2QEPaTZoppbN1uN5xPIBh1NLwNFctkT6vE5oFGifcL93mdkJi8Z+
xrzGa93xQL/ZekaT2q14MBPdBt6KEOcMlOH0shSODOilx4CPzh448Z/ct83EH1JB
T+L9uU8EZDEU6m60mdVxqBkMNq8WQunNbREuuMDfs+OrI1kIm7Rr2xHv1hpssXuQ
IAtiA6pmY6cgbP45pprr6/HYU+TZLlGLiVkYv8OalvWh2F5Zbh6YBiCGBdFvdQ5y
dUD3ejimxV3TVP9UobEitCAJ5bdaHDT4iDbKiD6e5pm8r3kXOmIsZDBNhYz68DxY
OlPqtJGRGn+45yTknXintV9M0ij1zDmDJnFFmUYGEOrrKedJiKzf+aFbRSjPkC7e
nQOJ86y6xd+aVcMfBjD5rMjaev8av6HVOarJbHxqOnDWyZWy51tqhkFLuH7TdNhw
nzgVWfSLCaN2g6DCsRs1I9u6b0+ntrKQnLaM4LUsYj5yZakTnhvRCOyocnLq/IYH
mLTG32pdAhimL2oryVc2I7clcDErjjsuZUQAHStZyueXiRxXEvT8SoGUXQSK/VM/
U7oiYs5R9o/7g0IMJxkrmYdJY+lJxMNq6WLnzQtmc+IDVuv9Ba/RfeYmZRkQdKS1
sdFMXou+ZiOknWDJyR72TbdGxUP965bydm/jnjIgqBcyaBwlIl05qE+AVGc0d3aE
87WpmRlZ0eT3jtPagzRUoGG5b+Q5SrsY62yTJ16HIZdboRpUYBZlVK9eShlCG5RS
fVycjkGG/aHH7c7zAMRYL4fF8J90Q+0CBwAIierJnFkVMlGjI/b619sPBkDmjPhc
ZANa95SKWDxhBWL0pIhJ7wDBIXcRViJgFoQjPZO5t4TUYykf47OOeIyzbYEx2k++
1vFIxPMFrxbZmeSRMdgoZvtXLeuzd02t+FcjDEslw/8G+Amj4dq5WBmQPm/vhcCq
vD/vgR+0sa0hYMSKTpbZ9gFyofQUDxVURXLTZWDHOqnkBgr28S50EEWkkGX/pRt9
0hTEBaNGodAbfXpU3OlwsaHwfy8wyfmiSmdGxmfXGKhCsMyjornVP0IKVF5ymJFs
C4MqVRuHyJqcywYI+obiVZYvO/a4HxfJ6NPXCfsiRmMsOb7XBUl4RLYrccZEIA9P
bGjqZR5WrrHsJ/YLTnBMEf9M5vkSCENlnZQbYEaJ7wYBEp7aQgx/3minUqBplaoo
wAeJj373VuT3sENG4O3Dn9TdZNTgU3BtpiSQMP+KEShVUR2AV58+jCQzvBirHKAI
8USIYo6uRBoIgp7yVoWFfZgPrGiQqbiNokUblsb7xUMrHEZxstgV4ruTCvpmVPYq
dgsxkDwoQbvvMYrDS72qwpGsCLRCdEjYTdH1nuXI1PqsRcJuzErZBJZVW4XNDj8V
PPRRRtFne5HDdX0VMLTA5ZIlIEc1pVqL5W8/WmwsGhAQ1zO9hWKToECBgLG2CyBU
cNbh7bSJQCA6ctXs0zFZB8HUhfLijaoSSbS2QIAC9SW4IT8mcxTW5NHESAvzeJYO
PdRGFua2iiR/5s4QZEAlPH6Vizv4da3TsUXOvCIF7Uacge/0Rgu0C7axVxONzws0
ebb8qfBY/0caVs8PXwycTrtHcdNAl+U0pBOoiQ2zPF8M0u6J5vQwTQ1kn4RXjWr8
RkH4MPYSxGpUadD8LxX2lhuBUbEO2zSVgidFMGbYC5Sx7HfuA50NAQpxjCJogSUI
pJtJZnoIfR4ujsmEx92y4sRRLw/Pbwa1FNGVJ6az0/gzMzj0gAxKoYSpI/0oVs20
OUmwuCkzHDwtnDFbpXmX3vPF1Gm3gsqgcQFt3ObgUReRI9wE9oqI+6usgtjbCj/u
Z0bJtx6rJlWpc5UTduyUz5xDMs9NiPXWFbwgvhDJRTH5IEpnDuQSfwoOS+gV2Bi2
SZHzssjjtOcMdFlQhL5B+Ua7xYQsLHu08p9LiP6FpYbrFI4aeYEe7qdzMmsk9A4j
kd+O6OR4Ks8COTe7lotNaVczO74EAhJC99yvES2iccrJPVLi4KkBhA+nbBhnrVip
jiBP9/Xuu8HiSsIwTUP3Jq+8/tNBspmG2UkUXcv+F/UCdVmNGy0GtaNX1oBWqlQ0
++jlB4BFcQjtvU7e1B8mx8dS8mtYzpDotFtbzLqtl4zW3OuCkOY0QU+9kNbORdsa
xAI2bUvQQPzdVZCZMgycBfZB8bId69eIJ8DvmFOdQCp/BPgiKBgCE37/VAI5Zirk
1IrxnZQMYLrt6ooEnxNPWrrx67wNDDxvdQhg0ntVZB/5DaRcziByVUAKBBDrGq1H
gykL6NMCsmcs+VaWt9RFXTiG1rQuDyYs618AOI4EL4JtnguAJsx30aB4fr9fVHJR
XZS7Fp3HZhlsWWf1tJnP76IGrnrlRA8mWYBr1kQcXYG8/P5Rok3LOJ9AMVcyuCKL
FG3rfGwydGY0/StzPn4IQl9Jz2/HLqutUxPTYz02rfuDUQGtaVIeNy35iZRZNkJ2
BD/vAIEPcliWtBSQ5ZVEh8U6vhyCVxV/La/x8KPpX0fWfEzmBUL6262hYku5LvJJ
44F9eq7Lf/9GCdpemvTRD5cB1ZRc9HwKVH9R8nM1HgadvdtNZ6Oa+E/rz+PsT9XZ
Mf+3SZVFokyoDX9ht/bvis/Lhpu+NNyWdhwICIWFO6ihfI4XDyXFC30RBX8J6acD
WNs3F0d9dMWZnNlAN6pp/vJXoaT412cNSmn//BwUmeyRJmjvsbu0wG0FTvTj6Mod
I8awHzX8SaJ638LIuW63Z5+W9vh/y37jBKVh2J9X3YRDHwpmMn0NKqG5NnyDmKBX
QiQXd6O4IHV6s/u/UaKq5Lzp6SJnGtZ8SJxBaTjI8ozfH8ristiYHh9uZR4xXvSq
dzBk6RqexBwCUl53ZUL7dpVMVQzhvD3wKYnpQCzNL+75/er7fvJLZ9ttA4G9pJG5
PwKTkeXnfrHX3tnVfX5PAYspKg0e7LTZLLEXGiFyYM/54Ihz6/rQzk9cDSrMtAIG
CItXDwAt0iAHoyd11rAKFQkRP8nHK3ZeH0E+6Hc+9kBXgAP8l4SdQhPB36pAY47c
a4ENdB3kHD5bslykDNkwcMJyCbk7VYPtjIM83d/bAOQnLHaXo6/cujLwMCDfnj1l
Jd56U7UoMGm+DuJH7QfJBOkdjmP13avdNP2qYHZAxdDeZpjIVjSUEJBk/2mPUIuW
6Sm6ny/FLpK2L06GDLTmHdz6LcHwUsCYOyLmpfY6WVQaE/idmzaHYg9N92LzRbjI
dqKew1DnsayZSWOd7Y5PjQmrfdF4dEDOvnxF7h04CbAOa5cq7r0YyWyqB50ozKA0
mKTqa3mnGkrJfT4YU7MZsasvA+l/XN8Olebm2LLdofzONHhb4V9tIDfkqhrWkIp5
1FWnnSTYY0CV+YwzaUvHkvGFGJlJnAdak0W5YdoKkWKDZ72WCuW8kAODfg4WOcYb
XE4AtCT+REKIYETmgyqu430B6O7rboSlMmVEOUUcfJXu8jnN0/Zk/1TQ90+s4V35
lGOLEyuEIv8+Jod6UoUpvBaazlCopm5NISDtvvK3VbTCj0hFzzy8nmKWynH6J+QG
bxpcS66K6vLTiN7k2rS0xpg/O6CG9A1kEvMwaRLCQ9CX2dTl/SoKFs+5Xn3v4w1J
xYaAQUyUY1ke0mvy2naD7BV2AcSufh67+eAn0Qchh+d3bJqSvHqNj2fEFXglzDh9
ztmkZIkeYFLRg0v+x+sMavC4ycG+2Iw8kDcftsgyB7rbbtT0fa4RV8M1gkWGG8ed
sOKAGbxPQSxHg3C2HwFvDeHEP9JTQhzetE0Av6K1QNetI7SpRlCoZActL845P86H
No+g59yFireMVdM2940VOUgxDySHzABq/d08FjDi1+411c+maHSvV1GDvXQqmFaX
2yBj115M1lILTLD12B8jz6sXR5yLzfNTRLzu0gFA8oy3zek/PUg9TI3pB5RiG9bh
XxklKz8cYOJWRPOTHtI/qMnO8g9UNbtSEfeUd438LqIiemZniqeHHdWZt7s0rDFW
RoPXUSgTnkrv3aRA/pWojtoDhoenc6rDdnPrl/gvNAtGUzbb3QMiV1RNN7qXMnvo
bhqX0nWcDki4lFL5MIqlA14SfSTLJIaBp3YcFDUI5cHcS7/vmukma1G7Fj3cjYBA
gJyT+OxkhD4/CUfxyogUgYnr66K7QLJbvXnvtV2/lODj05hm3CwHm7KJgzy/f1YP
evRJuRHsY8kfFx5DJ665/6bXA8gWI0ChAb9kFYu6vDIPtbXe3fDlmWhawg1iAwY/
dVLkIkwGRyFHLcCas0d9nOX+LlYzSIM9WwQAIgd7oCbqv8118sXWshycMbt2cImg
t+8S1H88Ezc+sgGq5EXCwQ/QhzyyAQVGryV61p9t8RoZNhjUpLQtrPfr+GciG9xl
wlAmklSjdg3A7gcJ2gMArkqSLv0EsGJJn6/pb6dlUDmp6GBoFx66GZnJ8GIArOpi
M2gZrY4FI75Wtpxj2v0yzyPSNrEZynehrB+LFelz7ESfOMjr7OSrYDVKd40X+iBY
es89Pi80IKNVilgb9JqK/5gNV/WO9Rpsxi5Amf8YrE3lKOI06h/DaSD1TbznSnMc
C5uif32lJygN2WHLi42QBXIX0LN4K1ChWVeTRosfbH0s/DokqV0pM0SciA3w+vwj
6VUOWZvBn36pCuZmgzgHD6yu6VwsQsQ6ZMfv3/YE6HZojBU4a30NtCxj6o7K/Pwz
RRMlnrI/eZrGuRMaZ460dZPO0j7kjLKIL1+6qWMZ7H0t30DW/ZNg8Rwc1G9rhICT
pSVXsybw+jg6kK9G1bN4aukt1Vh4u79j5t51MXfO/VHQuHkrugvsiHfmrPdMxTQB
cWEvmPvAgeZQDODv6A+9VqAdARDZHfGXkoIPaG8b+g1GeOR9DJxaIY1fQ77uqrwb
Nc0uPLrlz7ApWJyaMcBqPt9OJFl8AseF8GPxCxykscl3334riWVlgN/wZVK4FXpY
HmX9BGWZ9f+/UkWCdpuOWEBv+Ki/3QR8t/b+1P5RCdYcOtvXzINYO7Rx2/Uc0NQ/
SK2DqIu5+ypVC3mkUlb2xR0mgBbhp0IPavxm2mDF8moiL5EJkC4xLRDQmn2QhDdH
yD54xcxkoNLfeKe5ooPtTfC7Ym4DlAjpUAQdWxPjJ0sGl7hiUuYHMD9Gb6jIsLdC
CNaY1yprG4Vw4FYsLhgi26Wv8cZE/ei+EsyOOX+oNZR52n05hp3A3Ot2RiuLFjV0
HwZ+C05x+kvFKB5YaRYA4yLWpTs9/NiJDzrVppPuIAPmjU6Xpvv3wKeYEHJbr8YF
d4IxsZP85duLwPCkOa7O+z+HMntMxMIfr3faypcmMWR68r8A/xersLdDYZ0bWLyt
RpFRFGnSUx9oPAgk4AH4W34AqpMybhIAekDAEZ0FWURTCrCt8I7/HpS6ivR5GkNu
StyqWJQH2j8TzoyjGZrgNoG1Dr8dqavq79XVmanJ9zg7xW98ky168l4hdjOzcACB
I8jOEtSJ3AyG5oCRaexpsS2wkc+ff7vZO3prNMmcvUzoyUVHvuMyiU1cnxqa9Tk5
2o7DOSlBpyUCGMsi+hoUDelqT4YZdQ1bfZ6yCS1Q+UCK7jhUc2Cejh8YFIbWZ1Os
EyNLT/qDTzIpCcnJjJpajZOOwfEqRH9kuB9OV3ftlV6KE8cprzxDJZKqsZHGmXRr
0GGp6zqjozPvVjtdzmK9ejxbeICzXiarRlG8Zxfj0oaM6JK5GOM0e/SCi2aP8sbo
As3hgkP1nMy5d6X0Wq5AkA8y2FvSXfrdNz5zgGhgWD9Ip+wNY2mrRcp/+2x/DZu/
QYS00kRKmpI/uznr375DXrZwKdlG96houtI12ZMa+HNvO01zm6aO2VJdXsr4BJtD
aphQd6yQPchS3STrcINrxqxKe8QoKK+A7QdIiIwr+3zvkA+cTecQuTXMse0sbmYv
yGgYQ9FF5pULTN8ijbBacRg/Kid4sFH/BgT2yc7rR/y4iU1YL/KWXxrZO0oJNiX2
A3rCakxGFKcRhRhKqEU1wEbvA98mJBXNYn0QxmAHVGuKrSCBopzOAtT96j2UPH1e
O1MvS+Ui+2pX8KCBQLqBc1rVWhMZm3vpln2LlSR9IwUBAWJZxSTAt/NEHv2dn5SQ
zsntqZEMJlpcueO1hKAhaD7cb1OoDXY4BR2Ga6QFudkxyo2NRPKRQSeGM4WXL0RA
6UUd+4JfEmmERaXhrzuQx4ufe3UpRtlJk0hDEgfk77dCxbECJ6G90Wjaj9jtzupR
ahuiUwyUohat911xCHUhiVVG/FsPaoyAA/d2LLxVMUGHi2rxOdU90QhJ92dGFjP1
2Yw1JC57fyWyZRxa83lWczCrt1Nn0sGTEm2c5uusYQFJfaQagd7Bxsr7SYbPNHjX
wAS98Y1ArBSuRsUKewRxJ1r+KN9FvjK123isYq92i36BzLK9g/M3YZtDpSXj0pK8
uDwAE5wBh8lgFnmWLl1T8aRM+LsHYD0v8qlPMHNL8VuvSjPYIsdKVuJQyQDKqq1s
TKVj/hLdCNm06LM00djTPyMECcjNXJfb5WOQZss4+x3fOKzN9gvHLatAiHhdFGqM
pNMSHhuCExtpHWp4zzq4x0avx8KRGOtVb0ndlC7w4/hwMxXEX7WjxVBo4h5Vtgv6
F1Zxh2veOsz+eUFjC+6SUzZT/tbMcNUXw1YEmKCfOMECJivxIjabDJE08v7W/BKH
hRXCC3GcTrWmkAT4tBwZMqxjzBFZsgaiBHlx0mb3nszp1qw18cafpLLF+nyen+54
n2IptMojAe6rrRfPwy8pN/nk9rlvRdmx526ZLClMjWtTh6rsrd/OYj2Gz18Zck3U
vNGYveKq59rLrWxFcfwrMOSlsmeNo3KwHwv/KIW4G9U/ZdQEJmHoAtFA2cuJsSLt
ZrpbitfcTLcVWjjcL/f4Thp9uMr0gyf8aGfrw1nVKNsqJ1pDncyUtI83QpsuKJx2
QmiPK2RX9/LolZeFt7pufF0sR0tkmFH3ZcdiGm3lEM8CdzcTqOsHyvBIaYcaHuOn
4+Tfx2obysy+OYG1Eo3bpny8y5JgugZHnpGUqVXHf40hTWATT8h5bCajKCENHOY4
pV1wKYE+zr2AFIK+OhpOBSA/9KpL2FbUTmWeGV0HYD3r+Qjj11FeXGWS8CIoOtxr
qh9QX6Em1SDiqGDXdDMEmjL2PE+++euYW7uH1L/KoDnmVPYL2+MMcMLimDRCdSoo
ehwOBwoEVFzyDQvEVAPzr5z39BBpDI2FK/R7TJKPDEwoBQy4TRoWB7ecOv+cn359
ewDE0nStl3VVgDwzpcoVKBROhgjbCK9vyd0ABMrNxmP3dHdb4jDVNsVZB3/Hrzjm
X4p3aDOmrlqrhOby9H6LPf32bv4hlzpr0WPL8EC24Serbt97ZE0J0fr2ES5ci0SX
0shxtjsf8b4ur6Bodg+a0IBnQrymVZgA89HBq0GiUgsuTb/RAKQORGjAw8UDPsyH
HBhpBLAUGfQg4PRE/71NpbuiO0z6Z3CdmwlxesAa/8nVeu92TjqjNndtR27/NOG9
ixne3+sNMoo400RMLdSVUje25ILGPK7LNGCacfQxaZq+MUuKrTnGTfWi8xCUy5//
HTIPz81K7fe8P4+7NOL0BStST0CwzKKorByUovC+Z8EhXWkdbv3Z1/tP8I6oUHt1
l+2BQM2tdNjOYoQWbft6dKuy13sSvwI/AykokH0gHNGTOzelpCAFj7NbU4nTmoWs
jZ3YuclPXNpK5gVkQTbOsZofi1KGZKbA5tqygi9DiofAzQlWSio/EfA/IPkgwQrm
p36FiM3XXMcGYmAef/VwRj8Bp6mQaYojNhYCzQktUwOvO3BJ0oaRU7wQrksiPPKr
Wgf3r1mK93AfBYlamg2iPhBCZS9p5Ryez5BFAWLa63SbtbRYsnT0d/MwfqqrcwHO
HKGWjVUHuQGDJT2CdEr/VuGP1HR/PV9JprESDWEFF7HtVntIR60pfRgh3Oc9GcQh
tx2PpErBsu5jA3axsRTma7VweFlUZNb3n9Zd3DBWefTmC0mZP+qimrezfr/tgfos
tcMMm/rQhTvU6ThxvyAf+vDFN+zicc0WbI+g0RDLBRKGzxhc8YvljnknJjJqupie
djXqc5e0SwNXvQW3esCjVeJRpa2+nVhSZODarC2UMXPKi6OgsWC4FufdhkvXE6oe
LUB3F6JshkocstwS3oSI1wDySDkGXtmJucSc5PVvHq8dUiVKkjuykCb7c6SWDJ3o
5LQOPwfTT6qqffSXy0KIQxX//6sfTTT7Bi84F9LuFbHgrl9BNA6PAf9OKry52oI7
CyeE0xckTSzKhgyaKoIDp+vMETZUsfnBHVcwi7sAlehI9BQdiIiq7otMatElNX+X
rKZZd0GEvlhtd++RQeEJpDPl0YA9T+CodWT4N8bK/kp3xqPYiaj5IjaFumbv1+f7
5j5MH5nBzn85B5o5Py5A4BJBYTV05vGXh6Ose1DgY4kYmEHL48vAiL6p6tvqrM4A
fd8HGvrpeHCQmnTwYol6+KxIKuAEQd8I5G9uNymJ6dBCS82stf8W78WUKVXS8KLF
DraPP8acNQQSlOJshCMFClA92vEQ4Z2lzGbBcGTWOl9k1OIF7WWlwKG6LrebnVTs
WEBX/nPfKlNrUS/k8EfnckPklIKAGyYl8kzHXFPfqBy3CC7/r7eSs/h4pLtd+0kt
YS1zXbeLye3vsiwaj2K+smuNFItoh7VBne/3ZULpUbymz8BPaErriSSibnK6F1jM
PfnZye0I6+Q0aAZQCTa40wM8HXgsWqd6FX/8a2+MmpAb8/5GhL1r4FPf7Lu7cwjZ
oa2Q799Y60hCPd6EGRKI8XYAmzZTi9C9sCE+Gu7QfC4SEnbzKd8vRKFfT5JbDNDQ
QjxXsa6S9tVTRtN9vWR9NfqoHSiAALfVMPHz864mcKO/37jJRPISrDRVwL1lSKPJ
I2hLUac8G/PysCxfLlHv+STyhw1e0NGbb0ifeO9z1YDyWcDuJo6R3dXnRdcxGCwr
GLyZtJinEQQxiweQhWrbRq6PcuYaLFmMyJG33LsMXqw1+TX5XacHuPtsXSDGrjXM
r3ZPUBOXv2ygKVgfgrWnVsSzHO485L/8n7pvpLH7TI7a09nQtIiChKjeQ7Ao8Hgg
szSVZYBfU7K9bmygOhd1rzuftir3pdyexG7ZHm9gJupU/IxWf36OCkxcxNKFxxex
hpWF1zWcEylqM95ftPvSBz9IEeT+enKzBqNfn1nykQllSNKdWnhqA3MSDcuPvEUr
f7D9GYkhEOITcXyYreDnnlWwuo4FrS4YSOTY+N/VTqYjOeDKfd3/HuLc2MDdN2w1
Td+n21EO+w0HzONRsyRRQBf+3ksP7Re1HgCGlnoIgU/sIe1xP5BrbfNMNSbJDmGy
VEtdc6MId5/Gb7mXM1Yq+bg1qXUGgWDDBYZVBcFB+/emsao1MO1fPvgU3PVC278U
ymzuzZTqZHtdgC4xzJUSNpjeBER/mWUVuR6c01YiOge70ir8VCArqhtCjkLCbynz
7I2KmqbnazEUhstyFHv+JDpGUmahvbSWXKl4P08IidPLtlOWTpTul2fKGG/ywbo6
icBeCgC7kjJnl2l0Wz7noZxk0bImMvNEQCGDUMlKHuxdtH4HVGmq39nIXuK7t1oM
Tio97jlMz9fKdrbzf2qCTQDbveuICBtfAax8PwteoUIw20BLHPGwIonKUYFJdNmm
bkAvUBB/mJnOGPsyhSxxjyfMMZ8D/yXIe7QEyNgkrKA7yCsnSCGeITRRNRrUGg4t
kfgDotot+U9lLHqYP/cnBFO0ecgUc8sh+eja3XZi1IFjXDRHaTStDHWWkIa+etUO
/TuJDPZC7Ey8TWb+Wv0U1ZZTrIXWV7yAmpBbW8EpaPWI0SdL8I0xfHeRFC4JA/Sg
3fftvHxI8XQzZAUgGXiE8rSvgkOVK+XG7CyeOERnmeza6io3qR0oWFtg/QO95h4A
u134KP1/P7gz3JYmEt3lJsE1cukD7fU0/dbxqLGNn7EXxgyFk5btdnKFBzEovY7Z
bsMURT55o2vBNgUp//1MzT3/SQeYSm8tF5JKX471Z6mjGaNBRFe8XDHZpttxbWEc
fnKKBl69QXCMsMpYkj3hfcgSJEK7BZO1gGtC3VumVRAzTZWerwhDKUVJ3bYapBGw
p07vXBfT8ilsX4S81035hvNftFXPJLuXS4AWcRnE44y8fgpzhhOmHgJWk3Y3fYls
XVb63Urce5jaNgVnrzkU2r1UAwmCDhUZhKvPbs/UuSz6Mf9tdOV1So6VxGkxD755
UfC5e6CsdHE8RJqXXh9qmB3CYVGK491jXSkIrNrrqM9AWM3gj0FXwOpnWcq8A9ri
yZSgxE8HuO9Mvf2V34PVOaT4Dszh+BvHSM4zyrY0lmQZF8kzEPPKp0drWNhmuLX0
/RCmUz1IsHbo1uSO4dU02Tj2PPfuj5bRELMctFBrGtATPdB5Cqt8H5gCbtkokxRL
wXgfkX2a/VXrDdAWxj67px3A8fizu1/VexufUCpBtzXei8lwjovJKi0gY0DTcRR0
j5jD0nuQDeYwwCFTQd1nw1IKtKV+CAfpc589/1GBn6AKGCKVMOwYtqgx9UGqn+sd
fqeXH6QqG4DKVpF7UjrmJU3iS0/57u9IhpZiMxowuk+DZenRtpAuTCa7B2uyJHB4
1Bk4/LHS0iFzOhwB7UD9cBDr1qfoGCvVfoEcpE1Ca1sHdFtF1lrYu/EGtF8TSLO4
Ra8D9wMS40Qqgxd+Z1m6xErkOg687RITcas3uu04l6ukWT4OhDnpo40eSXLg5Bug
lVuInqj6yPYCkldryMBZXTMiQ3YdqHrmOJyCCxT99D/jBCf4+kFG4in2O46VRTTT
y33+kYIKBfz6LiGUiVNFwmuiKGYpyY362x0gWHwx4bFqNgkv0pEejE1xt95LTSLr
2oLwBFKthSF4CcT8QeV2f8iUleGEwaT/RrI7E+UrWUQ3SbhbuYLa9ixoBNoUopVR
lXBi4dsc1sEysOZlrQaph0UfUKJCkSZeEbVLhNdt4pvXTjMQoVGedxLHFFgJn+6l
i0/s3ZOrKeDRD+gDDSeaGN9p3QnLgP3vF1/BzSdnK/dxs9BsN7dg/pm/PaeZzANa
2uOtVUZmJOe9Ku4AeJqRU84TpjYaGkiYvZ1j8lzgeryTYSIc/gQ0oL9LVIbVxMEU
fib/cY4GaHa7Tkgr5smxCARg5lM0vC+9walkyJMnd8xrN4ep6Rnwdrk7d1ADPhCQ
iG9u11CAv35DJZtCVaRY3YXwtgW1GB5XEBRfv74E1BMwhqFOhfDUqV2gPAuHQQni
aA5dTtwoPJ/VdX1NBRshxq3uqS9BbRwTDD3d+mrVfTxbuT2hKbtOmUfkVdT4wB9A
uE4fl3cbpHOv7/cRfk2z0edwcWDg4VW5wl1XCI/mxLmpuUi3fdwIr84H4wPP24l8
yHg+HGD1Ny2Exw3srFuRt+/HXLX4R5SnbuGII4P+7CqiZbLDJXfa8to6wht+6xGE
grQ13sK5GN3HduWtCdS9e7PSD5De1yBMiX6BpFmM+nq85N4aBfCmvopRFklTTJmA
JTr5rTkvgeGoRiXd/ScB5QBT1iXs7X16Yt28WqaAOO48U4RdBblIqe6w7nMfBi0n
lcwsHXBRsE2TPlJgE3mVlQ==
`protect END_PROTECTED
