`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BJlXMN1gGAv1di2t1wf+zCEGy9YDvINWu219OnaV1Ue5QUUApfDDoRu/4TOp22rG
vui7nxttXZWf+PcG0FZxf+HA7soRs3nsPOGpRKS7upgEvErDCIjWb+TI6kf3K0gE
SpJnboMFXqj52tAPZvWo7g9GlcR9PR37q7xVPZynu1FPr4s3lU3hEIIjYEVD1+RR
dGkU7ifjqUgwb1Fs37Co/b3P7mpN/SuNDcgrdSIrcthKTOWp/ftCyOZ9lh/2mkuq
QmMB60gEi50EoXlNwTWR+57He46wTkjXwqlSwhHobnY9LuVC2EfSlRJtBw3QnKo2
COuhNpwfpviptY0hlBrVsXeiQSNDFNoyunJ2r+Y4cYZWUoAbLRnsKIZpVclCqX6m
YWGNhRJfoLttcdIXWyZDGttNR6jx3ssjTZ7V7mtUSSho2k29YZQffQqUvDFXskz1
LLGded6gvcnyWMoCnd6D/IuuFIxyYFucGKWhK5BJGIqJVnG++eg/4s994J4whUla
Q4RGV14fcU9EZM7E/km5kEnytHe6+XgCkS5w8zVFkBjmsZANnxV4lnjj7y3a+yOE
mPVDSndsXaEWgovEtZD9O/g3jdm8JG4+3wEPbMtq2lJGeyv65yAuq88BLMaoBC4y
/yhfDqRcaeGmY3a3dezsZWUejGB1rkwaP7zi/aizaFVCE/VrGU5ZQaRG/SEDAx+u
4E2RkmmauYo17RlKGG62+LtJCSAHbv7zvYZPokpGNF1Jq8/yYWzN+3XG51Rr+Ckm
dbwuukMAzLtMuC5n05CUMF/Z6GIabAirQF/eGWJr82j0CQKw3QwtiP+MD5f66m7/
2xjzt72L88GBMK4/O9LA8gXARPK0i6NrnAYKMQ5qnXsKp7LSmFdjyGiSzNhM339W
xC8BTpbNkmYY0U+aBlb+juxd8IxNGUYsQUfj067YbHiebdW1NJzlV2EF0wI0wUan
32olX5JBfbn8marLn6XzM3vfcJPxSVnItMWGFxIu1qiy3600b6Vh8sgM0b6Wr0nT
6KE3sJT/mNZXQoN5df8SazFMYG3THFXppdKJpjYHScszjs1510Tj6D1qmOyhhgLq
`protect END_PROTECTED
