`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
faDlsw4gxFhfpHK9y5b88ozWhQIkEtgCmTObiTF+aiJEVJ+0fl/8GqZNVRXOP2xs
LCY7MdUvKb8afwOZbpgF1YDpfV9aDby6h2XoA/QUKyqnWAWgYfGrm1dm0nbCqhDM
9LPgjrbcVJu1TGFZ8fm2b0MQXyGpvhuQUfABLGLjGUKduQcyMNSDOj2Rbp+buELW
BjKZekEkAhwT8wI4WWmarLeRLZdQPIno1seHsTBAroNdaLWk9O5+y7EFq3AlwaqN
osWILWPikbxpssTnIOsAgnqMf6kNhXv3kgFXLy+7SFz7cQirml+hCr3jniLFydx8
BnAw9X2XcCRl74/HQCH4ehgyTuZt570y//xJPOslXnkwpo9RIg8tQot+usZiyCTo
2CH6Wb5dz0ECN7jod4S0/SYwcKdYXmc6udC2hZWCkAiR+tSQMDlIsFdQSNAJOmJ6
kNZQ19PGlH8r0jSdtr9rX/TzKFXQr4ABOBNY/aDL946buLoQ5toBuf+9KmGFOIt9
+N7U75snHqjp8D6ZE3voPFOHiOPPTtAEhXz8p2qU3+WtatfdOKDy0NGKxdL4gM3C
+hzuKXYrAQ08Q7ZNhoqIjkymxizGyGBHcZsBPV5A/nMBuwWoINODCHSF5E7dCocK
5IkI+vcPlShprJn124Oam6KigT6IzK2YTn8AwtBjR3pu+92O8A6OPS8UXz3w8KzI
ya5URrUf0//ean0F6Rga/KSwZiGssA0Ajf7NojWwVCzosnCeGm7rHOFwUT4ZuatR
iPdFYMSoukwbTu0CVALSp0CaCSFPKcmb2jf3yPawQZu+3VJYhn3ArRmlcRtlaOmq
BsrwQ6E5iMLPjJSdvVuJtXCD3clnPVmNbCuqWKHnp9TZ/0s0AAzCJdtrRhnQSj9n
wt7EwGTw7+VY2RWrtLxc6WK93SO0AIZ0TkHcpSGSf+WDCWsT6dYhdma7ybubO80b
UdaTjKs1IVO9o+HBJLUfKkyxADXGVUON92csxJIwGAB8cx5e5WjsbFicfFSY1Dbf
hrzjI8heb7l3gwFYaP34r+1djca38LWtDZBRxhS+sejlXKMqCb8H1lv7BSUigjUa
2FPI9QatNyOQ0W2OqNx93J06e0eE6JqtI1Etb5uaeXL0+fUJYyXRHZVnMZqZMuQC
`protect END_PROTECTED
