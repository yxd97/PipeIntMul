`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1oMC3Pv22PCDV4a0v2BlExoqccBbS8qawP+tTfGcY00Zah2e+d/JKAi2AmLwIuzA
CsgHJ9Pkt2OaiLn6/Jy/xGA3VDPsTSoHwDgLTFvXYwskI6LXr8LDpIhXG8p0ThtO
0CIWRxKS0l3shbiMC17hahj52Dj7GaLSkaF7lP8N8evx+GMdNYHmuEuvgIbRKVWn
212xzq4tisfskVyV/efbHAQc1RmQBrLenfiTbxlHmy4SESXxXEum85UDV9Uyao6+
BpPNjMlozIIPsLSal4AyApMT3XB1PJNFHn5K5emgv09z7AxqF10jtz29cEzkyxbB
xVX4//GWV/9/INPTO6n6pwd+cRWcTyrofhc2kJrUXYazwmbJOX9awXNCpF50lq+2
fbekh95WKj85NeVl9YqqeRJetxO2ajSoNoj5gEGLgHkGZdqE0lxCVrHRSdkf/NnU
tVI5ipg9Sfpo0NqrRplFh4YUgJJscAE2YIjSqgBqbi5YnX2m5XriBibxe5PqVapN
HPvrONJq87XZi1SUoG3OxW8jRcPj0iEXvEJgXOEm6D98dVUzOh+c6+8wmyX7tPns
nmbiabDk5jRpSgDh2TgNtQs9dCBP4r8ARL19syHbavsAVnuhve1oj6aRWiILQibh
Bgh2V0pwA4HBgc8Xq7Quar2tz1g9919GkU2jPJD5fhW65aMgjRMZ7K3Os9fgL2Q4
75lCS6UJCNWLS7WF7nnZXEXWaGhP4JwyZYzxVaCSWZcgFi0dyjMoevQa18wVVsWR
opXcv+aZLF3+qyf8nk9cgw==
`protect END_PROTECTED
