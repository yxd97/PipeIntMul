`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcn9DNFXgHtx4+SU8c6VyySTj8o929xEgacUj/CxzVqNbWuUTL3kXdEHFHEc1MlX
8O8dK4dULnOx4SfJxbL5raNmiNDWfouKxt0l0510L/9MV8BujU+guYEMPNQJUA1M
AB8CaRIy3+Wc/ijnPsBJC83WtAMxDuY/F1FOXu32Aiab31bc5XvXypJQad+fIHNm
O8PTcn3zkrJk0yUNYcKeS1bMeYP/rEKPyKNkBZ5kJDAr62fQrDNGmGfY1dVAJgEG
m/0GNSM3FBd7K/uNU3zvwpSu66U5gNkCeKoQpWbCwzrMyG4v7gsI8TYCzPyewLx5
PbSV0ks/lB/GcADdxgAg2eYGKKqc3cT3yxCwpSYCOe4uKQFAWzgDfh/r1M6ss3XS
6FX25ksV+nEif/jobH0Q69Gndezaf8wZFPOfvQwl9JgHWP8n4mVPFBdSIsXpIXEq
NeHqgWIYuSxB6M7pKcg5fxawf4657flMHtkr+hr+ak5fZavTo7tXgCOF+t5G/rY+
P4FPOT/VjzHjN7+SuYbMvOym6MfL2nDag0SLK0hZVw3UBe7Y5vKh071Nnz/RXE+X
hSHtkapH9m7ke9j79jImP61eUSDoJyIXgnsqU30L4m63U7nSzAfJQOquJFieS1nP
5rPY9Vxux7R4sZ3PYyxL/Li5ZYa06OJgD8V3qtrW4XB6S3XynKgTQt0KCrhg6NKT
/5ba00Da+9+cR5o8A4np6rforNUEJsQ8vHC7HJZtYlujAKnJhGqXCaT9x/KBTZVY
Xew/wi67nhU98Kmv2ZXcQ/Gzr71AFzk+M74iqDppE7XCnddmn95YqPov6MksL8Qv
Q/s+9v2YZV7L24+v4FgFBcfIH8oa1idzyCKBOZBJHZvq+UwhTUrylb40PTbkqmb+
8lXbnhdAFoOV5PuOTQaxVPj1YSVFPC5SjPnpkCrs8iwvU2ECKD20yZrimWEbaSw0
k5NM5oozdKO5vWiS973mEssxUApWY6ps4LR1OHEtVTwXSxoPuj4vsTBYIJXRwmcY
Dq1GOifl+rFOq1quOB1+3R2hb54tbLTVLJ0VSsiT/cCB+ybZ44m1oZuC/YR+FC7p
vCUZhmzmtOXmRV9PpgOqsybW+fM8KTAosZkUrDrcPbx2+fkwrjpr774pP30gkea+
`protect END_PROTECTED
