`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qaPOF4VQfsjGt/UFP0FkGIsO3YlXqGsb+q2iEXpbzopTfm2ksl/ezkP+4lx3ojCJ
t0fBnoJ3qNmVX200Ln/il9ad7TsxgdJFIG7PZO8MjeH7jWuZROTV5klcN/ps6mDE
wUp5jHC14nwtHNGZANUmFhR6sbPpAHL7UVOIpWfm4nQEQdKlvtY/xPmvlhPCGgTy
sCIl5Of7MfZjhc48b3eCcA18GPLS1t8hiCsrrS2lJURtqRKUeokJB87nHw7rAJMu
6rUPicDzGvWoWYbXovOXJqPJTxpXL4U3YqpK3GReNfUbyNTUozfC/tkDt0A+8M8/
8935N529mp0H7oMvwzymHCkQbvBg0zhY/8qgQ9Udbl8bYsSlaxXCC2dv+OYe7uXa
Pgo2QrMl2Ox0VmVODtIoh2UiUh5bRE54p0XmieX/es1ShcbmJzmDKH+ShJ73Ffia
`protect END_PROTECTED
