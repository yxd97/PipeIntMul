`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3yGWvs3JdhTAXkIjeZI4pYOrCnJwY10sNnMTmBD8CqLDx3yVUQmrOpJEw6iGErf
gOi/LIkzBSDol9hTlEIHq0Po2DXbCYOhUvYsfNfpnjfMKe3bEfP2DsIi1HlhWHPx
jQ04j1fPHIOAuhkdY+NU8txdu2inizXFsemQqHqYFZ3rDgC1OAlpy5Azbn4mW5YN
gCGVUA2D2fMG/m+reP+BltsmQcY9uiHfEK7NpPDXKEv4Sc//fiwrOxG0UI66Zik6
fBeyLH7In+fZDFN0aa4QgeVEGJrOP17b6NqiiQ230eQoRkEac4jKVg6KFHIAbiIr
JaVy2KrYGGvaALbCIQwAV82nv/Ky9CT6W74CqQF4M7gcdRBtRs1/XLZQBoIDOWNg
WazGkQTxhqsxTOlKf9GhJV7zulq4Ll+Ro6knV0fEqwosRhxl95g75xEslrSIA3yK
00CCc9tBbLrV2iNYkEOJfdNJIkS3P5jkVefX0zaZ0xPfx+p7f5Rxywhd6HCW3LEc
8dEbtufUf1W10gnaKAZjd22QnHWUiMBU6Tg5BHtNVWvymF8K+py4mkwWfwk3S57v
C/7xyVPgdT+zTSOAoc1vXhizZ9CjTsyPjLFeJq7apOxbmSnJTsx8hTZgsNhwvJaV
Kcwq0BteOdTH3kVFC6rFrj/kMU+atzUMw0UkZfuErLhEMTKR+Gp3ymnnv/OQFG6x
sjhXkrfZ3Jg+xyatODiJvjRMblIFxqfXyw22jdZRG0yupSdyXKBBnAZmk3LoVXER
OCWNG2Gk8b91c83im/6SWC6LrEPvy8uRq5gNcFSOaN8=
`protect END_PROTECTED
