`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68HuLFhgKLsPlCpA3VHlLe5w4eONPNej+OiaBWfgEcPUVsaju6w9Mpy8xrM9nlw2
8Raggm+pscKQsctJVHrvOAxX8NbBqYYtS1WKs05yedtyESJPCgi0N7MtQufIdrLm
yn0FzMrNqCjYq3P364OPbXdqMRbh4BaohY308qyhfO8gI3BLEN7qQaXr7lGJ+ZRv
oETlpJhqJ8EVmheWOoe9WlQN2+uy0HJW4BS1K0MGqRqw3vTD3aB8kczxneF/kGgA
tt5ux7AmJJmQkIQnv+77QRhXiUOp5+FiCbiNtPMFKNU3/ECox9UrLCHYmAawOpe4
K2/BmjslMMPlr9EzhlExvaB4hAUp5FCiR/DKqfzYW7tzcG2/SwcHpgmovvjgexwt
h1yPqY8c51wcZwY66O6BM6T1ujfvsu7AAKdwRIUgWOcoIJqiiRcancEg8MIHvvOX
PsA5zWeR5Aih4yywA5CCXxmV7soy60dRQPd7EN1bYn6BcWFBTn7E/dQLDwNhVC9l
yGsvjYAxlI7oiTZzMGQm/eX1nH8g5WTrlYRXn9DRIAo+Przw90StG2L5TxOug63f
stbbRXkMNqO5od9dxt6J977U9uL8rHI5CKgtULMe0M4Kr8qrq4uyIXBTuFIV95re
Qj9P0KHGGv12t4OY7jgwAzkB25erVqzdnNMrA4OnjlG0xj3Sks0P4rvH3TTfMZ6/
Zz6oz/oMigoOmwRg/jSo0vDcbW8ctybJ6oprd3D0BoAnJ6q2z/rt7YoA9iYqBgRL
DlN8JaajBJgjXmIcH+fcG7pL6z157R7OUcLWpO34PkZaMGM5sBLXyB4EpNEAnKjX
lSIRYx3kJcjRr26bzTpEmWqdZH0x820Dr3geJH8bFDppvdXf8SkW3h1/xeD+oSZP
esgapLCONwrhSorS/GP9uYtXq4yRGRA2NdvfVN7IuscfwsikDPZdZS3WHWdk9kil
pSyiw/+3J905yLOrpZxANw09XH0ZqpFrRRhmDSDREXWvE2Hdzt2eO+id+WE59QnW
067wfyDc6nHiNk+iBMZo94hIp3QwKyRmySz89Aoeis2y0OByGOY/edn2hE0dBAAt
YtzZdhG5t2kJDeXcutOJMoCvM+BQZo4Nby7SA2zTfJvI3S4NwJvgvJfZGcO6cyju
HpBdxvscL2VyxA8nvNoHq41yfa/q6FS15HPzKUCP5URn/VF1K3lHcjN7R1b1wo/z
Ndh2YPGSKHZRXGfwwow97cemVFWEqZ4xtEY8xLls68qYGb5AeNpYMZg/+n4yfc9/
PWlNky4a5wubyJeLzCMQawSzDIgwieiSeQiL6PIkWZD2KrZK3F4tjGxFUD3N1KMj
BG90xCVn2BlfUz99UtJJJ+sCzzbwYGk7rqzm7sWq8+EsD7N+OJ+PvTdLUBTTazzy
gV+rt+g5klFCPHDlc4e5DVHG3szwTbr+7fW4VjIVnms2DkJWhrNHa38VvxhT5PQ2
ECS6NjAhvvzGz7s0Qfz+E8aDBTbYSJPOrRgxQKl01TbkrFPN01Q+S+BUMhHrdFFP
7ri0/4uJ+kkmbyiL0s11yzedROin/yO0haYtmfq+jbD7320Uf0LyPjoZJEyJQW3c
wzvblbrVnA+kTNBGU2wCRbqPBmbqUMzOT0Y7Mrq0xQYtv3H8zaPOjFwpZIBlcEvq
U5osO6TN3nxgQnNd6OE7KbfbBZXHADszt6rXQny8DXwsVVGV5jXeZTFxSDFepTFE
e1HjG6QAhV0wQb31H75z85n3UAqXjfpVgfWMUqMGjEe0B3EPQUhyl4GAFpAHkIJa
wBwDNHQNOcNlysXZfpmG9NrhlYFmHuCuwU/uSbveoxGk9V0/SS1p6dzbtYPmVz+k
MSUD62vZ7I98hsrCXdQXKIplAQOzfgVVNOyfNOTYznhI6XEXGZP78P9nDZOz+tkl
yB5E/llq4S5pP0a0aaIKLRjo0t+z5L/RzdQ2+gOrTkTpRvE3CaLXMtnTiytsmBYI
SJRy9wUup8dJqz5WbH8O8Y0V5VlqaV1yXDy9KQb2DE7+ARslemfgZSzUZRvSKLOZ
DkO8IjO9WJyAIv9+FuK1x8aLJ7KBJSGVvAjxlZL9YFmlshqbYDuk2av+GrhfBjyC
Wy4fMibMPFrLt8x+DZNRTpJz08NgBAzcI2jMaZ2OMXL05Rl8S/Ga2pcVAwQWeXge
MR99QwGJ+JGE2VbjlKJSMrFhpxHA+TpdCBkCYIjGL+wkuocg+9nZQ4YNF22tZmvK
Qge0hT6EA8LT4tWHr7Tfx05ZbYHNyWZ+gQkSw0DVq9TX23FJpFvq8FnhyUSdUHj0
f7xFQJpnITmkl81h1P6JikOTfUEgoKerG2BI6CIe4TNh7q9UAIeQVn0Zd4jZeEh/
ugZpExTB8g6wNqoyzGBJBU4ZG9A6M0PIwZPJqVXrQrr4x1NgfKvrY2IqCS6APtoK
EFwQddgyTihoLEVe1z77Dx4pXwZ/TRHtysfmH9MtvpwP2RcLyYp8PNiVAaGj/xyp
sYQoMGn1uLlmTPE46Ykt8fmvyRK1xzb+73K3t/Ki6dgJnPPtXRfiljXfZhc55kq4
lHjAIzgi8ITt4FStHEz63AOk+Xs9N6uA3j75QFSK9Mum+2QRwMvydgQhMSXzES+Y
rdyo5VfaVanOfkNfAOdhVHVMEjX6ujG5lmDPFHAetEansHIRJPnR9fYab//CkMQ4
TGMARlUCDhIeJMhSTwXqrcTiIVsAOcQ4+W5BF9EE4zluqg677mbDjLIZ/2VgOlUU
4WvRfXu5BjqXdq+kCGlzsIYeUPBh70Olag5irrmtKv2B3UQb3U6RYfNH/hMm9y4n
e6ZvVlJgB/NNcrset2JzKP9mXF6u666bXKqEzfmK0LrQGlaGjrhLhy6FNueyLcge
OPEYl+iS15HxWLEJS3Yuc3eGwcTUEec3z0DNJ5FFB8Njiv9fiaMbr0JZawyxI98Q
ZyAVf+aDVI/3PFoAl9Sm6mmddHBETh3cDTuRF1at1UrpS7xP1SXKgicWfhG/TmSp
2hmEAP2hgYa1tT5FMoNao93mzRsS1Kn9tZOgYWlrNib0jiWxWyTZvB6ho7NxgxMn
V+nL8vpD8wVHh4DWrix56o8cSTvELxTbCxk5DCJM+NRMr/OiXIeZvC0NZqIOq68j
W+v7deqL7WGyu8kBWbdw12z0sRK9pdq08Lwf6glHbPnczARtAbHrSvy/GhER9tS1
sqX2y7aK3u6V+ty5s9ZQF7RzUIyrTz5pDPZqKF30boJpr1ab+ubPTJdTtlBmkZ6/
rA0rIX1O+n1AEBjRIZ0/P7g/sx3dBfyzEegfiPUYEvIBnFb5ZXYYDMmValmjfKld
frJpq+lbgYOlvx9zr6Sd4/FCwljnRv3fL4WDcQLVlZGHYqtgpJ7lfnPEXQTnZ6X6
/oPK1o4NlSzO+cRUseUa9nOgy7oXPg1QpKuGNZemtjxE1reU33cxLN5TWCFUH2Pi
eXVUhxVps5wfyO/0oEGisTeCT5YsMBlkWfptHZ9KJCcBbRFJ2wpXzB4JIoWq4tCx
dWbcRYEcR3Nla6nlVeyfJxihXJ9SmpWrGQEU+3UhYjrOEgsmRzqBXHPH9Eb6a6eB
pKogGqkAvuYmiWvYbbBgqzzdgHog/aFhjoe3PQPxD5u/3A5TbBLXkV1vgLE8cdsD
ZChW/s1OweQx+H93OEYLgyrPtS6OmxAxV7BUzpJDgHToW3W4C+F1I90WHGugd6qS
vy+3wY9vIlvYGhCGjUW08cTiDUW8FuH8BP1BATKPZXu6dj8ZM+3LAS29aqvsejC4
CJiqK04IE7LnK7Ko1gt+hH0FfBlYZRcBoW81iXa0TDICtBAe1C/IVNc0OSenYvaY
B8TbseFBh8KyYeTXhTdWft0AVk4CCOMD/nUnLI1DPmuTn2zET/slTz3tyIfVK8Lm
flGpvpdV+wOHOOQR60bOLG18iWiG0BrY7UdLjNhhy1GkeWCYMtRLQZvpS98VdZf8
XB2lJas5ZhPLpZzIGQW/n7a2yoyZhS26mQK+YPvX34uk5oz9bIvg0bNkjaqXP9qI
oa43zab+uLoz6nyWSaob6rJJ4sP/7VbpX3SfEY3TKUSXC+0IN0yBgOk44dYg22Ig
/qMlXgzOyPrvcM5O96juFkjjuqM++bdGukHsNUFh2DwQuOKqlRRv0IZYWHkdAQeF
5P2ahJ4TqHH+o0vV0QSk1AMfohi/+yCmzR9j9YrNqzrH4B3sPwjtCe1SzKcmpAZN
f1k4aJRkjNIy1o4DDwVOq6aiYGsDBG81gAqnyWYNKKrA7YCv9tnA85xyhTjzkUz+
h0kLJ0VgDn7cHVN6caZ98JEuq/und4Qrb1OWhci9fiOMVxT8MiSd797IdbIWYUIe
xSWTBv+uPt6wl1fEwViiC7KOvNoHwWBTyUaB5rA9o8pcPuKoaXRWDjrsdhycO+SU
ZEEha+hi/INLpDfBxHF5eWO1IDF33LVKdxTxKdvlGtLaAtRRiAuiaF/r0ArZgtrq
USys6w28orpxkH1j4jjDyn+/dprt0BWrVJg8y4VY12b497xLMDaDWuW6+avbPQAe
iejZsM+cmOfpZ06/u+zC2QickFDs+bPV6tcTwUFvSb8FIjMpsNy1W3yGokIk3/oh
anoqjzjstaPZKfx2PCAiDucb4jdwbrXFPJS9hlAcaQk8ciw0kEE4IM65lqeRCxnI
+Tt7Nd3LAs4VpCeXG0BAQx+RISeVq7xmegqQH5rkS4zX1nWBw+zQSfpL2l84QADR
7/kS9FM40hPLmq5Wsev7dhGJjZ7YcPwUdgvP9Mef2RL6YQM5co++L+/5izgvkbGs
u49fpOjsWsdxJxXKkQmrAegvWEdK2db3TtgcCqYohdJlcnRXkANJ7bL+4QuqaW+s
hQTORWDFBZoTbVmcNiazZPeXMSpCfcjGPLWn0kdCvKtjokJdkVrniVqBf09qbKEf
UQ6Hlh+yqp0KbKDi9+PDavHueeB5cm8f7onL8crHTAZ5v/2vfeALr/Ik3LVD5i/L
61xsRjnFq+RmTetnwf8uDWWIQxnIhjBkQWKAdC3HvtJ9U24w7crSDsHFWHAH1wZz
+nvj/s3zfHJF0xMFVE55u5kS2KFFtHLDz+LlNFaBP7iTO+7Pu5535uTdBtiGOBgF
dxLm1rIJdcsLgqSxqwnRjmuOyyxZbAZGikdUbRXyn7m2RnJD2FMCEpO3sJz7P/G1
U1gac/RGf2+jV/m53AUyFxn49xR8G4+SwqWz3Yfy61ExXARVpdUM/NMyNn/JdTUp
K2iYtwUVXi4umE8lksc1StgEFekoarCuiSUWGiqG7dj0M95pd+irZDynmx2gI7Sm
JtaqYMIADdZGb6P2kJVfHLRcYS0CTWmin2Htgu233M7YTPSFUSEvYXUhCKpahkIo
jfYeVOl/0VMjKXtfqeZq44i2mk9vns9sQPA90KZONVJFvoZE5wnCYmridRQ4XH6l
Y4mb4dx7ezTUYdC25iRdHRDcLJWEwuyJmKbEv0L4ci+mttoeKx3T4nF3amjNgvjh
ZgTV2ShasMzNVSrnYrN1lCmhDnWq34Vdtsn/tymZNgc8gLDshihhJmu3VqoLjEsX
1HcjBpZPXz+MxD5SJNrMJij1HyMfdqJS8f9+YSnrNw+JTmILH/Sskw2yhnF2jK/z
tEAP2sqDH6UEWbzgiBcQZCloYGwq462cJJE7jCnMB51IoAiFQSS94Lk+DTDq3+V9
+jZhk8/hyV9PtxklDfV/Xv4ldOLEAoRMX51xHMV6lpwK5cBgMrR7iTECqo2RxsWb
w4EZTvTTnnK6sFSwA0PYawsKkf+AA9xgS8/MIyHp/9LsZAsDN0yJZ/YPgHUXFUhx
u9XMJ/2F7vsEikvpmDQXaXcg6Lo4GlD/WYWp10gz4Cjp5DJwrpQ9Iu/jAMKqZDM4
tqUQOTEgPirkdcYmDVfs00nl8itZ0atvMeB26rGI7f0SwTSBgd3kReUemfJZTSvJ
1xGFSeP6QT29k36ezrGiAom4v90WdJ8g4DV5IWFqWvJpqDnSRLZJ83FaXx3d5++R
dj8gFZ8PZPituoifICHck4hfpf9vSD1cgQScxSTIS7eANCKrqhfmNnLa/mVaAFn8
quolyGdUGtNf6w0gThfJfg+CUgUrFd18IVJYT99g+SgrrZ9W8rwQo2rNwZXT7O+G
O616DE7+PCWIxqhzyU0balw3YTVaE4qA5STMvr1nyQs9O66p8j3fJNcB6JQDXPgj
+pLKieBeKbE+7aDQaqIY77272Evj6z8xXElY4Ay6vqAM+4cFaN1Xo1VaSYzVEMYE
ZQbEmkvQi9Pn0w5W+rSzDDUcFGEfZ0xFOPrXk1Lu+SEno39GHKt/90CGDmyxPpT9
Cfj8VaEpqsdX/PHfO1RZaNZT8o30XCloPGAUSgFDGYXeT/ZNl6NDnYksXeE/ofqq
aJv2Epr4JdzdEQBtn2eGB+B48zKaA7U/47ny4yilnaT/WqFNJsyPDC0yOi6FICZ0
MYId0BMbJ4FZcwjl7yIV/eslz8irTvcRVkw9zDKAVJLHwt9ePAIeSt0F/+ZV/cur
+ImXSFpssc/4w1MMvgZt9RjU/uZ8RsE3aaXs1HkTsW3E1kKkg82zcg84nnkG6hI7
osg8paXrtGcgB+kr4pB/GxbPqFvNJJGVMWB3tA4sTqSo7fvyvF/TSGR+19AVNuSD
YmXjXZdcEomL5f7FCFZVbrUGCo5Z0/P4Ml07g+E9+eX5EaxJZskPJJ/c1jMfyo0o
hqxXnyewycG+N/ttV4znHPP1TPtJDo/lHdCTbQrbZv2c6FcvBE11LtqUYQHXlDic
p+Nu55p6oXLCwLe8s3MYKz4NXwRJwJFowmDaC9OqVuPLyP6w8wiWP5lSF5QsW30+
u0Jjji1+Inos8+GnfrTRz2xRuI2Zo/N9tLS6REws1Hb6/lmTi3CGDt6fE55lOxi/
RDVfmCLDYRmk7FEzP2cKy104bUzGBTpFISV5qtPi14L4n5IE04mBzWvYLUjCWSQk
H8ZvRudSHxFF7sXJvAKlgPU3jAO1bgEHA6Kltr/qsqnaHU41tOFFEYl0UuQh0UwR
7NhbOePZV2GSebAW8pL8kv1+CvCx7M/ymPiLvpjff9dw6S7o3w/O4JR3+muwvfwq
6XbgBu88Wjp4rruA4fCtu+ye5gZLySFrGe57aHF30hiSS9YoCA7qzsIpnqihEMe7
wYlJUw0LuxwuY4ctNA+R26B56vr/Y281MtZMSll+ssP0U+iPfKi+Xvddt7+/R8Fc
jsncJPFKo/uY7b0m9RLJyAqKitEZInviMq0tvWv1C7FeJLlB66hazJec4H2bdtXL
uPEy4OxlxpVyANhiiZBzivvkt/+HtLZ6tR2WLo4r85ihLxwucPyaSOeE+91wZXj7
froSRgDCGNLCuiMZeOTHiawEuWAnZLtP51d8lZnejc8JWtmiZFL3k6oZqnwrYVMK
Clb+/qkrLfbnu3LiEUXz4Y0Qg+9VyY89XguZpZaQA1YXYNGixdr/7tpM5FqgmoMD
VBQKG3Hxmf3rpAfZU/jS98AsCioFiZhC2FW4orSyV/7NVfPQcLXgODbtVuX8ZTgx
6pvprOxpGlm24sapcTfiCvAyK0cfn/SLXl0fA/v028BBy+xbOgXoXrBJJ75KLAeV
rRFNuqv/DB7jyPwu8DQxcCbjGP15Eo3aOFsLX9Rqyy/QG8SP3D2SYz6YdvbGUMAx
lzu7DkhjmkR9eNGHT1qbMHnUxYMB2wKG5LrlckqpV/QuJLfXKY+orz75wNme7yF7
09/H5xISeWxdImKF0gy6MGPZEsghWYAf9o38kag6MTUyDPwfO8MKencL1OR1rJg+
XeLV9+jQxC8cqqG+vRskEK3u2AlDVMhgwXMXrMo1yXFN69+lFF7EEUdldC1YCzRg
XQRRKaPAof1s3WEXbeqaT/RBK3doq5mKaSDZgE1hNHpPqUnPSpuyJdJadXDmJQnm
iO+7crH117krY+eJlthTpUeQA2mquwSFs0uHAdMsgnPq19Q4DcyiYXlarTacmbTq
YErnKSZ57hyQz2cEaX5h4DzdyA9mkg7IMySWUcbe8FkXU2X1hxn0ztakx83UXbkx
M/uXzYWWhZBM9QGf+4Dxoc3ANLurtY2RQeEQzxMpf5phdCrj9l08WOMaQEiSKQnf
PiS8blYTfs9KohCVNd/MvOaI90nRu9+SBOBKAI6iKXlAKLQkPuWH+C5dfezGmKoR
g0mDeXeKsIfyLaPkJi1aeXC/grxx0TAUeD5kJ0D2uAJfhX6mLAm8dP+9LJ7TGfYY
DDkhiX56bPOXNVMSTPdZ8vcZErn6nMnR+iaX+oZmbfMdQqrSq9FXRsN4YJ+Ce1tw
ahXwZYvSkZMywkhb8SwZ7Gr/XamV/nz0AVvg85ZQv7Bl/nQvXfr4IE5n524OisL4
sTCqi7Dtb/BjFB0zfSLVtLSD+FdCOqr9Dqn/p8Ztd2u7Ax2s15U1jIWfVZhl5Efk
U3TdRpIfJbWOLIWU91K5IYyjq6iZFTaSyK6e1qnhzuPOJ6FVLt3EYgc03FoFzwgN
Hpt6QBTBezZ8VVvtagVU5XTyzeVVsn68JqQiL94xVkOwyWrpqTVF+G68NdzYdOXu
b7iGqvHhhTVhD64e12Lb10AYuT+4Ahq740Edrq1OZQOuDbjPlTItIs0C9R9uX3o3
3ZSZ8SKoBhxMnoZ2Lh0c/gnPU7INUr+Yt7y7DrYnSb0vwY5eO2AdAeAmZeh0m6K8
HjSFXrOF47KWFlXCSuuUtkhTnJMqQg4b1YkSJdDEsVNnPzvuQ5bOU/EGMX13U0Ut
Pqj7MQGFF4huB4olDshjj7+CXRXhtFzsCeEgd98vJgHM55/VoeUvdbcjteAIgHHG
AGO+W/opA//5HuuHp8f5cFzOwB1krVTF707fr0xgKOMLmxjSewI0FEzXrJYZhXjz
MAMFMB9GmjbH70GEyG38KzS3BSNzbBNss+2y1YzMs47OxG8MbuBTj+1UKbEKsXLl
uikT5nnbnnqgTdxKTj5px8kVNTikeEbRRpMprp1U7uC4264zIfLj+YdRQkCcA9dI
XJnQpZ5kNtliiGmvYfS/Y2IvooYt9KH8xUZRztL8bYtl69B8lDjraVye+WyjTfv1
W4RsrmpLZ77+EKAgS13vM1AEBz2m7irGygWloCNSfdDxMbUwvh88EYbXFNVlouBp
xkfabMAzmLLaHdpoxV/EoOZyXeaYgAMHnucfzDqEgt3subEBy9sz3XVMwHc7smdv
kZVRkgWEiRRzh7ZsFPXYFmOravTWwRoowCG4aCZpYf/poQ06jLXj7sgWjcnYrics
IsdF7koi1J8gZoYJKapD4Mo/+QBBOFsSBpVCQAcqGeUYjlRTcNl0uLE+bhQ9b+ge
jFbo2TNxSXpyLFg7gdV7ORuzVHhbnea/Mim49BYY1K2bA5dRdH4iJ0qT6UkTfJcW
7R2AZmyV5opOfTSuw2CjpaagapPDPWF8NZCR4UQRXhtYfO66TrG22cyRmxjigeMV
SC/EerpiaJhLzndVgxArQM9C46HVx9F8EFZqKKZXmUjgJkKMSpJg3AB5ydhw7upT
8gbcS9EIzfGkPaC7EBZt2yBZKDu1g6XjgbKaQzUSqQ67c3mCBvGSgJm5dd9m/LC5
gfh+TQCqImndr+ytv+b+TnAZaLSLInBiNa+UdyjwbCY6Z32meigG13x89cpaTihQ
V2LyPiLSMVs6pyD0B8oVcR4BpPLzhTggP6ro1xkvSd/BpqBZxqKomGkTXZqNJkod
WIvOreqrTqc8rOyw53y29yS6+kGVrQqvVoijMuoa2xrq6/vo+1S2Ie7e5O2Ya6va
UsM06IRWVCikVaCMCRVgxs3w/13qPkSGs9Q8ptDrdI1aCbBYIvQFsn+CC/KXQ6p3
pzaASJs0wFRq1yB2D4smxcjr+URJl87u1epDh2yR6T9xV+HaGtxkSB7+GXBCNPFN
G3rmHTdPeLE78/7bVCV+Nx/7+gP77OA9vYUbQhJs+q2pFJsjMzYLOkdiTkwUB+1a
OXeYp043qw31dvTkNhKAyyoNOaAwpnD+iGeMqcLghcCOwFtRfFglt/NyQkmg4Jv1
A7sbpevzaZ0m0++Psmk6qBo2T254KiTMf5mhtdsKPlHprha8NVmcZIQ+v5mqfmu+
pY+z3iCnyJKRbXMj9gCBXI7nNSNHCaXzgZ655/UMXLJ/HBMl+OQuYoHz4IBjSWXP
/gVDbpcKs2+nTM7e0t48lfivXqrJUNfaIeG1Ql205hHtPP6Q4L/j+IKoeNxox6Kk
x5tFtqrsswKBsnG6XP/Cm+7sEA9HxwhYU+iESrrYwEFccDxWV0Lvo9cIRmJSD1SP
YKxYgW5s9zx2IJ1mIMyfPawLS5z8gBT64oYkmrKkBTSzZ5cZ+iIqwFm1186sOubK
6LtlpnxzJFHyLvwa6HHHxYm8ukQ+UvHpK53pEH0VyQrNbmb32vSFvjIhsIp5E/Wm
acay60HmBvAp46EwJ+XsAClNzXwRRo3L36k4GGS9IHlR0tRlq4mVWYNQcGNE0mag
ZmqQqCm97qCuqPP3+S/4fLt3uqjoR1hv1b/gyfQ7+mTfdgfhraRyl6E/UKeRsx6q
uDTkjtuMK2sc2Emr8HRycOJY4+0B+D+p1CwegBSA/b4b8U8dntbM8V7IJJHuOJbf
UoD+cvVMmHhEWGUuEdYTMUHQOx1+HctA6FSYLh1JuzEND9o7yAc21eZyZ9fHfbHX
IZuXnyfrZL4FriSCfHyutmtvwoll9mUdG2uAI/FvWeli7O8DraBEzglB2X8yy9nV
zSHJdpz7sEIRjwSRjl9CD3FTcFLXtWLNDhCKpYGAW+W9w2O+j260z3N8u8yJnyXe
lIXEuhRLgU/mga2t+tYRQWDyqsY69+S80ipzofkLL9BI8CyhT/anG8QrUxQWx30V
+2/VVcDckBnKOkr5P9qYCol0ntx5VjoYL4rrYRF41vvlBsokJVSs4Yi0VVkDpWFH
Z5ih7MIfau4BSA+3qcUrhDNTNdNB+ORdeHQXdU/DBYPZJzJ1BslsArCt/TCr936F
9jCz7CBiheOsvh+jezgUicriRsSSErhSxX7qybw+/g9VflTNZFytcnS/5SLJtxeF
zq8d7PCpdXD+9klGs8Iyjo5wzAuukctZyHiI3D7M4/kNVNXVMqXo4eJ+X7zzOWM3
8lOiIVKcpKz+deKygDOqKouT1uH361LveQIVAbJ4Tad1gU7c996aAxSTwwVHt0k6
h6RuwrHDhpFtxgkZS+JFKk0x2TZzzo5nv5caWGv/ZMpJhKpQhd/dGz/2Cme4l5gb
iZ1fvyR+uph/YaaueZVTjyRy+IbTE9bZl4sDK6YlxNs8NRa61ff4ZIofsUS7Mft8
4oDAo7TMhS3vVwWNi1vyVSUg8ZHDviDAECm9rn4mwr1wHkdQTeb3DOd4fy1VLRua
88eNPuwcGxcq1BVDcmsK2O4zIJ3y6X3CLQFVDPQ4XHH4qulDgAHKj0Sqcf2ZC2pz
tba1LSE4cV/BwfTQOq9C6xPF6fftBGh3kIXINxOJlHZ/N+ojoUyqxcZIyzLCAMUP
R12hBP28EiACuqdeGAhKyb/5J/zn8qGZOrs8ntVe9Yo5oIA5GGqZjP3bmIiVoBx7
bynBz0XzrqRIRuottX399aIhoHEopRvt6UGi2b5u+HrrE48hj2EcIC0gB1eM+xNT
lK5UjJlnTJB2+ogrKraYF8GLzsexZ8VOo7ptRB4LFadY+FlppcluVUVGLWKZpM8A
1VWRgygWU5Hr3Q6HQvuWh+ibyte/yjlJvxlbZ48xMAlFgUnt7BW5a1MwuebCFpOD
sLZfzP7SKx4doTR421L6APX+KnPB4dhtB/iuOBGxQwTCYksEI1PyaOUGOUKnfTnF
ToEFA0JqwYFPqZU3RdzaP6PWqFSWIss/jDq3egeYovgj5DznAInDmhVuF4qEIP/F
yyoCkqlgf/tJ93JFfZOau/JDZqwGCHJu5EpLewWCmAdmSRnOItd8BvxxNZykT5j+
Bnk32wG/GY32z3PVl7q6kYwdmtQLPdWRmH2Ejk3zqOu7xsqO2r1h4ppVnF1m8SaY
5qHC6YpVqp6AWHNts1RRI92qJcY1AxPG0EFy07pIAlEIbHrtXCJuv7KhGwccnhuK
dN34bmBlpGXqNWQ9UxjtkXKerg9xe65eFvWzsxAl9UEAVrUn2TMKMNihCxoUO7rT
6HGQkFuoMo7A2G9C/gYe9db+prXj1FVvK5EY+aIsJvpDm0uW7hWvF70p5awGkVie
lNJuzFb8rtWcACMU+isqXDX+qhOp0pDB0SYrhunVBr3bvhNxw4Dg5eaAZbVLyKj8
M+ftFFgSw8juNJLSD/o1ZUSRZp003jBNMHm39RI23IBH3/6e3KksgZJpveAJqO/b
8MUq+JT2xE+qDY5w0OUlVp3pMFx7Ql+aNtoj2hKecxtSbMFuYziyHdYLkcW/3vkG
sf+NEuaIapaGE67kaWyvUbqZY5/UmIBJ9Hp/eymk8VblW0idLlGVVOVFoFK644gB
Q5dLPX5rS4N5KF35XMiva1TzR3JjKKvK/jrnRL9twdAMb/HbqjjsLbOtCZ9bkHKq
J0jsesBIKNhd6It89IO2BirMZ0mwyrClez6yHBmPF16OVkNHPe4MJObxpLnB9uWn
uRatxfdXUSwZYa8jMoyWaa1iHj9spmjF2OOrfNkgbzVNFdVeOPbvDHDyUYrg/XFH
5rxK6/datd/ELYy1UCDZwudQp23FBgNUKlt/2qAz4DWKZlLID0u7kb8y67Ul74jm
un+y8VsA2hWLY0UIWShHmiQ1ByT8/LjVy3XkL0vR80ytF4uBrtVffxKzJ3UvqIFR
haOMo3V4G+ZX0XfpisW5+I+mREfoxnOy5jgKvCXTtMWaTw3fkOuqHKEZQZkRQUr7
On5gutdYiLPIOS26xtooL2C61gzjdNrbiEMLohw23dm++Z/N7J/ahO9DPQKOu7f6
weH5F4M37e+F4XM2ifuw27cIs0eVtOnb2mOCHi4ZsdvLTZaT2evPZQ5KNpBjlgpm
KDL4jVk1KQvAFVX7DGhbl3r9wIvh5tgBuq6aMwn0lkPLmLlNS+5dNiRVoZpG80RQ
YhdUmPyE15VvDBJAuYCVWRKONvi4DdFbbZPjfiCgOArj5L8Ea+jx2KOsl1g1g9AE
2/6yQh8usQAvn9lGlkwaFliT3k/BOnwpD3d+j2cdjqpyUNkehcJOTJ86EwkYjPTc
I5pLcr3tq7efQ8P+nckld83A8GRPV7vizu+0lz5Ih6EswyeTaV3oA/kKNGPdNm0y
1IWDSLkOc7XDIKXSzHt1g6u+5ntOUOWFco5QL1XJM0hbshjdq+wMuTpiXgZdyemw
gditpUotyi1gvsoTwGaKqN3GRS0X4qsh/4r4uLiSqNlCTMKKoYffUTjlVDv3J4pp
qjOFT3AddPnInoyetn9Wrbw4Mexkxinm4rYqdCT1y5D/URZeZnDvHwHovS/PWSnm
uGRW7GcAPndqxMFu9OaG9bya4grWyQfkEwxjcZ4eC3bjI8cgimfc7eQ2N3+w3KvG
CtlLgKvy4C+B/hqFVP5kGDzMQsBCEXnVoxKROwQNlRX9xFazHpJ4LhPVwZm6DjmB
P+JFCs39ij+Kj5iKs6a5mEV1JbkRlxY5S+SZAtyvYxh9VJB5uyvU8znYpFe+5+dg
lnh2TIRqgedfgdJJBK5wQhLZkqmVyNhfnEapsUSaydar5s10QDiQ44IOJflcSa0v
0KWyDjyCOqs2JtAPPvbDkriJnYrYfEMl3cvwajElwllhq9845QeWdGz987Sy/XRE
0G2+6YZtI0oQnlYpFCBZy+qieZVOpTGp18Okjtp2bzzfer2tQ9oyHhwTRJRImHzT
Om0+cvnQZuUQRTD+Q7ETh0RNMbY4qJ0wDiBDIZkc2hB1z3+jUhyixnU9R1ASbtdU
iZJe59h3uT5ZBgmWNxSsAUIA4mMVPp72HMIFUQu0Lmt8hn6qH3wvMyozQVeZwCJl
6F0EBJi9RR3Y6WD6lAIeS0VjmUqRsjlGOEuZdH51BYJ2J5FiLR2JoyfUu1baecYx
bECPsg3rN49UsO+q9i00ci5Ev53yZ2XKBEf4rVNYoEMJOvDWvy6v3cQ1srgkujd3
zcDwR+LauWN9Z+OrFtrkAyPI8B5SGVSuLu15lO9nt9bfsyfChmhbm2E8JxYPSA98
2cshHC5I4pnvUNjdp1xp2xR/7H+KthGPyxES5uFmenisshEY1UZowDNZIgX4Zfl/
4vtf6Afc5U/36VCGE45xcV0gXXpsYU/z8kid7dHyKyfMd3gXWoa036GFzsWiHfb9
ATjBdZUhGokxFAE4znUzXT02s151ghDiKJgxC0emWkW20/zL8iIMP/rB4yKCEHpb
cjQMh2WYlKzhCbn3ZZ62x9bR3pLYf1GiybslXoVSjDhuzCMsHSar7dQnIl23kKFO
/aIGfixhxeG+H9JcABrCExM/92n933bclqruFUVSNL9LMcGF2julo8Uw/HCc8pwF
tHdCiw3HdYGqQjMddkZq7aX5svvQIGDAECh3zVdRvAI/hZ+YsJVXbSoq5+zQ/UYv
4ozB0X8yTQXR8TbCs3hRjqgabItrE/icrBu2bPypfQ1iy2EBRmW+RCDJFoFsPoko
8VacBWtDEfHFfNHSw0TzEc74NRuN8IGEZ1M74/8n0RNVv4v3T2G3DhtUTEHBp++n
pbIU94+eIP4OzeYJvvVPcqhEqHaBxJWUfwRGF+vIqehXI3ETRlPKKilGiUVM1d7M
AtwH5RVAJ7OKnli5LB0iySlucxnfNp2JIY2POub4HJxJyKKP0Ko9jWI8I7UuVov4
3ENyg14FRHk3iHIN1Gk4OVilFdO6r+Vrz1I9Ke5UM+OPpeDhV9/ayh8bVEYCJER4
Ma1WxlQ2cja7ZSdfzT96xUdgwHDFdb0hc0CpaTvesExE2Wz/EpEwX4eoCAUlvAJc
3kEcc7WhsUoEgDfzNEIr2KnVDQD88auKQ9SrL6gYdNSKMxbSvod2+s4aF3u6/QVZ
JzLkUox9tvj3mTcQrgpF6lo57VmIc+WdAeK516nx2QNNe4W0Hsvz+UJUzPvqM8ei
dn3/5P2tF6n4OBm8WR5MYY2pEyWfXxIzI624+UH9SVug9oZM/EweQuKnvCff87nl
7V14kk6AOULlO1Tmrvi692sG9B44Q1DBhXduG46ZSEi9eSTpI/VR+rzbMdoSe3qn
KM5tBrRsSyXszB0H8NHHM9ANhZz5p/t/vFaGz5XH7tV0r1bihf18elxU9XgIbNgZ
WBh0ryAUtb8UXgmECiSt38VZKrPAIAuxYUtFmvfWpsNKCxb9GuMedG7vsK9PXBBD
ucWUzkqjVZQlm/W6ANJiSfsRvJk5v1iYYq7680L4MmSBwvzp2IKKNb+oHL+lbNic
zKr/hacxHr+5CwDnONoWfylSZRmwmU8M5/CJ2M/6+GKNllidw7uBWEQgymoZrOVd
4tb2s8tiP5vz1qxr1adxNEpCxzlo+wSBaSNaR7W5xJnutRIl+m+D42tL+TDB0cnm
DsH6f0g/sS+Op04DjuczcvK+SeGOCST+uCG4hLZtyGcOBNN3Vzqw1uGflglOVLIc
bMHKccoc7gAnkDxfZ8Zcnh+RMiL8Vb5NHpPQ5gOBl0lBJL9+l2ZsHpGnCCeGkQE2
Xq+W+p53+c3dQFc8+IASlLEBxYr9Eg5m9/XBFhmcflj8LiYGVFVmZRGA7F/pTM1D
WunOisB2lmAPu+rgY8lat5V29e0oH2lEPb/UCXWCQ3hoyC0Uvh9weWRiGZYVMMVG
tIypudOg9b8Q5XzREa604PCkY+dJ2VYgz4X5IlqnfJ7JVMxZSSrSCIJ/Rz6PU6BI
NDnL3kiJxOobu8PF0rXajnCHU8716IHQk6cQpbekNmHCHJnouobG2h1RJEzSEsiJ
FUFoQiaSiOA9xqkGb3w69Ez8DfJiEawyzDtdk/eN4BLnnGhiLaKR18NUXGWu5cAe
tlnKGaCdSdHNdp9GKPj1JdwvHkMypf2uGM4vmONy1/KWyQw2W9/2nBY01Pe+OK2+
AatB1QwlVDG7sSULc22V8KkEdG1RC/8JUNClAd4k9ERXPIYQB4XXsocdn4s9/fi1
X+euX84U2ebBFGit7N/eu+ml9Y8Rd+KkaypxDc/zvkILC85qT4a0RNgy+CIe8HMp
GZHV/eAB/r1aQIvKqtFxPEx3Iboze1PHZgp50o4fRFZXF7QKJzba7IOzIRSWmaUR
abtAf91Cv1OHaP3raKdrmfpOI10j4BlNReSa1x2WR/02rJAmA9cX2RfqddglzdtP
f4iciGl36DjmEXrwqLb/N4uElZ0Kx8Cq/fwYVw2N01tTDYY/WGzaDYdZqbXr8tTd
/yBnx5GjOce/2yAT9zHcZqINX6qfE8FSGE5/IeRK1yW1gtw2L+h5c/M3CoSLHmBk
SqxhLSYrNtCuRa0uSvTL9HO5cgVOjgUzo5oemzcT1DImzpO34hlDcNo1HKJsAcJ+
qbUkt/XvmcT0KH1pm4aOthhCXMG2aD0mPInU4BAoWWF9U+OQyf7LBsQPhmBYEAfm
qn8ujQyD/5N9GxqOrjnMKSJdhdRHr48mNekGpSeTuL/fBdZPzERUZBwLruoyA9FT
Si6qx9wEmxKnwISpnLAaESFN2bbT07Pqwz+KrpxAt9NNLRR4Uym8z4KxCy5qBMpb
o/I04zorNpDvUdguxis0G20DWIHNJig7/dIr1NiSoNcDUYDD0SqfFQnKv8fMY1kr
nYD3SbSq8w/LMKq2gZGFDYERl8ZzWktoqWonrKRFFyRdd+Q2JgP+rqE91mE2sUv9
Iklx5oPn4LE0ksTftRGif4ucT1jP48hoQm+6HhnYN3mSs33AQdRb+YSx4q0C08lf
FhNSqyD6aslc4lhp4lF0XGhqQBaZC6yGxI+MWRvef/sFYSydsKaY5l1Bic0GtO5a
zxG/2/MCVvh5lWU2Co4sPExaFZaR+Nu4KpS51DF/wkZvUrJ/9n1yXZ+H54cptl8L
wpA534rOXOGK1YozkKcms/aP1Wdm+IM7SlwKaaUvxYp2toR5VKnQY+7zO3P0GaQ4
F862CqqQN5oFQgV8Td4ytfVu1tGlXLSfpYcgozk/noPJ5KQoWxu0PwNpeU2shVcc
V1yu7zWVqzeUzOcIv0symGZTzdvc9nYBf6hdCkja/MJzfWW+ax5Lgh6TnWvktr00
Kw3Wi0KOziMMhWCqxtknc8yNx2rAdMvHG8ziDhCgKk/sO9iQOx75vfW+BHQVJQ+i
JS57AQHeEgzaXjjqJ6KnndwEZWRjsH0TLe2UR/Cs1ZX4qwIYOjRk6VbmRHKkWNYu
fNp15mLyIaLmTXoFHjUfrSXJ2EhE0Zjk2TxydqyohIXpmv3lX5yiN4HjPTxfPvjH
ijUsp6cKD6QC4VJHbJ/tf2b4/nHIL9KIH2T0p//KOEx2jvGfjsYDsO0LIo58C1yF
KvFBBd+PWDt47AzX//p6mEphSgmxLmvzEcp//oAJpJIVJzFLpVxaerxXmQnAEaT/
BIyaATr8FJkegiwIO8uVZt57ZH1uB14vmcGgzTHM5HUauataoSkAWv0FuDEe5tJ8
BV/hVc687admuAR+/indzhVSPx7BNGlACgQ5YpMtjtXSGReQkZWWszswhkT7Xsot
ihy/hXFWJoXXAS+v6Hei6i2nNeWxRm8+dSl0Eiqyh5DQQvq3l18FJXbpKoC4vYer
ssUNPPIdeOJdslNwx4zOuKWTO+h336FO3YkH19JmCopE9KijHdVYgmzhIOZfzASv
mLP55ybVzQsK9doGniFg2h0GuvntCmZFb9qL8wRQwYTs+kRDoLr2Z03DNNIeIwb0
po/fRONwhtKEp/xwi0nqTbJ/oOU+Md8as1XiEpR6JbWcPss8WEe/oJwL90ePIMZI
bcdGBSdsFAHGLh6tssZ3Go/+vmjLHFJ0CmdUjgz1uaAhs4/4JcPjTBswSMl3vFWz
NY1crrcbiJmDLzB+M96bezoGig8VAZSFuGG0IcEKuc7v9zaud8LTCioQoMHDBEbM
0OUtkUPkKqQvClH6Ofuh/vJjMST1Lz93/ot4u03B9yX38J0RTtd7dq+/XH9lN+Bo
t3wsqgtwhqsYju/2znlibq90QOXTUxwsMlazC6Z1Iq26HYgFFhuCkRHqGuQE5H3+
YgTCJgOCjalIgqyrE8nB2RAebhL1KFWIMC8CB8El+VblyOA544FNg7bLSlTnR67w
cJogFDqMP66KxkQ79q7+PHRB7/P8UT+EoO+6JYbDUHksfLxuM1F8WXf2yQ85094g
n+b6/0uOl1BuMfh6WJy5j1PBW+BHsP7nLoChmsgbq9b8BMiYXRyXowPv/iQg9FVm
1/JPhy+6IhJgvwKoQFMQUIiE63bvpl7+fAZkNBhJTqf5w7o6U0fxJtxn6MFMe5Ou
1LAN1UZWubOFhzyFvBYdIaEPhKmKwYG2arKz5ycv5N0wylwCw2R63U57q8xEV6SB
raJIRdjlKv3SzG4xJBcvMgaiGTVrsgjfBXbd/yoYGKF4cnqUSV9Mat/JpyJGngiQ
3g2yD6DZbiTxaVSlFG429WjeAAtTkxCSUSWMj1Kn4aK5jwNJnZzByJXXmQ22eVb6
x2cqNdl/yFQM/FNWe1U8vqErRhwckSvc7gnW2SWTraPVfcySUvjX9olL3hW0cVrj
oZkyiarYu/ck0PiJqy0gehC69qdU4gX+h+iq57AHE0Z3rYu4XttAdPYx0bmNXW2a
pbvee7lc2vNRt2+8XxiqNEtsKa7aYraA8rIrrg/ly9GjMn7NI+AZYg/MlHb4Kibr
yZVxAv4VfZ9Es4qT6OR7NYVsj811r4ScwHP6QEZomUmKmHxfDDm2xShS+TriuuiZ
vSqyQjFLUvtBLu//PLDVH1TOQm6uqVbLNEGbqHOHqUcKJLuCLXeTpPk92b+jPOCh
FglWPgavJfh9NijziePfDCM/pI1ge0Q29EsVoohs3ljlpIrF0lezxvYgbQYMnAKA
1+AqhIHeGr2JvknZgLse5EM9dxsoWT+KvinO7Bzd4EzFZKA7h1muLhqXqk8TxSrJ
VZ2T/GaUmx5e0uVRdHxOE20fHxSrUL1YK2j9kfv/fV6KRXX2a54IcxWuwE3swyDB
UpColNCw/8IkxGoAcQ2I9rxOcS3NKXQ/DlK4Sf31in+bglT4v1zmKpxDHSYIf7Yx
p/D1zABMTNPKMktm8I6cOy/DuCxB28hBYq/iGsKesT/Xd1xmpwkkIxSG1BM43bEc
f4BRb/y6tMAChKhijJjl99kw8SC1/i7mg4UqG/0XiYJh/IKlSqjsTc9qGqN3yF6S
JloR9elTIxLUU4FOw7xZhXJ5x+r/4z/3cTCw6vgGyLAGWJ8xSbf09nOxLdBdxXtE
/S/zO1/uAi+NirFfPV8qfFXh0lIcMk7ATfP4Uuw/obcuOK72fklo9gqRIv3mMvGR
njLUA1WpM0kqCtgqY1td7pQAtB3JPpkmSFB8BbgMnrhJh49aq1b1M3hLD3d3HS7J
fuAwI2rFHbZl4mGhQ0koXAikqObbzCA/iXFKS73j8tFdBZbngK+BeesH80L4AsNx
4Ud4WLr9lgQQOyjbgiEEmFbRSIArc6ARfVLUo+MKP5O240nAilMDzqlrZNRs62v6
8aD6P4ulg+ErR1YrqzgoaD0Vhe1cHuDRH5mI7aF7x0Pm9NmCO9HaBxg/JBWS3bB5
RsqwWnxrUvDF1BivulGwrWof+sRq9qaqhTcbMG9n+6KPI2XEtfU6OoRO8eBXS0vE
dM+NDv4SChwBOKFp+wTQJeZSLfo2Lvo+3POemDJZUavm2QtAY+v3Yx6xvi3ggSDe
ovCP+txBC3zwxBM/gY9vtLVmItHP90UKC8bI64DYnRgZVTJFf3axViWuJMndfz5U
mtSxxFHiJSCxhija/Qhgpn04eYfeFJON7Qg9JIM+M8yEBESrxTElTDp53f2i2Esf
0pKI+ABTkr79ZgWT5mWXfjGtjAVH+PRaMj4qDZXXPGRZRoux1eI7aXb3fqrLFvga
oyiibThpjpeahOaVlhIVptCWeAQQ50cSg+zeyMAM670SFfiFaDk3MDlk2/1yIlva
fF5j2QjJjkDiezRuDW2kNK9ZMxJtI5ivyB9YympQVwkISykphkIAcKrbckhjPd+9
X86BTdHe0uKEcJWCusprFTQKjh2ScujRCgFL0gv8wPXRSCYCG6SiUtZycPM0u44O
WAq2VkaPJiHKZUHRRkV/nK9in58YFHtXex5HCWa3zpaSXySQ6Pi70pVyOwpMr5k8
euKbaqgLk6nLnuRhki+xidjiMl9Orr8xGDJbHtqcA3jUGWb8Eo6zzffokEbyU0al
g8hq1Lgb+WXWXaYzW8kTbhUuh51k3Qk5ecPz4j5X2HN03B/644yvbg6LXVF+SIS3
rAFG8DC5XqSPlf6RflLgYzAHAJH2KFJ/dTr/QcMPP6GfBPu1HzuOIYox55GuUiaj
6Yv94IUOrvzpGmmBdsVtkCea+AGem09/F2oDIyf+GPjBvmFYLidug27t8lsdoV+0
jffnxwvxv1Eil4jAJ7K0uCI2XzKQy6l391WvJzovQFOCu+a/EhWjjxdpogxe1yRX
dZRsO6aot+SndXNCa+kXMgljs9OWXY6FqfPKo47TxU05br5soyFO+4sn9sxzbIco
T9xZL7iPRNY9PChUBl5Bv9RIUfGNSrWhkPSVoteuercWQJP8hnTv/Gxrc7auUFt6
KkixmTSzMH1zrjDTlrrUCVR1+TZNJP3fGP+1f97X/pjLRv8lCjQ5RZHEJf7nm8Is
F22uL/hJzewfYsoLkml5DeD38gQJ15rW/zL5Thq72L/F7bzYGr0atYliK5eh9/ZI
s17KGoEsoJRfgnxu5BebiKI0O5ihpWKSZMs7CVrgaE4zwKT4AIrKEr1WQeKd0KEz
TJqExao6G+GSVY78bYYEyTiR3VIUkzzCI7VUcEGvNGlQzi/bXiM3C4QT5rrJkHs9
lnNv9oPnW9zcyrhwHO9Z93QhVhHAAmP16Ox+jUFShj5enlXuxiXmY+ydx0673KxF
PzsaXP9pdBSfNVpaKvs2/n2Tf9WA5j6bVVItGfCowxHQhEjUBsfkyP0pWu2D6ZNB
1GdX+vwCDXqDUHcXzN2mRwVbfQkH8eP9ym11OOUrsoDFKVmax3bqHKbp899h2XqB
bimKVa0N9NxUmqsgUXN0/qaYiYjI8e3eEEoFmZl3OZzhAD2+t4fJaKOzXIHaVTu9
+LRzBFYA7CdMem/NMKiiyL7ig0RSX73Grn+Q8oZIiVF9/5UTQD0gQv6z1D/2mBq3
oRDcooLm0CA4XB4NwR43iyuJ3ZrptbX5z70Lnt0yqgXQqcL1sHns5AovDBu9VphG
twjfosT0Z2lAKWPr7uZIu4riJmgtwk47Lp9dlwyuSc7zp1bxo9qJlKc+JxS1XH61
d1cAfi2gino3YLgKF2agVfmG3maKSPrm+vrbYOe+k9ZeYIMCgXeSFl8tqB7dh4e5
ys0AMTHG9Q6OH+hUA6MYKXEEHn5tkVcwwx2BP30VIxHCLoEuyVxjxze6cVXJ5Y1K
bc4p7Hue0Uz/iJ0b8qV4rmbOVXwZrTk7qMHjqLmxWiqytBG85BO3EHFqutjfLH2v
D5wKdx9y3cs4vjJLIfkFY9WqNktBfMWyOlmg4GS2NCWI+AKDg6fVFTiQFPHdz3i0
GCNcwrLf3XDPra31HL4+dLW+Keh5doyncHec/7PpMj7/vK2K/ZNPKbGOA2peLsmv
qj4a3fE7rlse/0x4wghmZlCRCehucLqSWtf2w04GxlrSXAoydCq3d9tFq8kwOyjM
+YUDhYT6GM7Wod8tpQVcTf31egCOia4SPqqT4lpE0ZShC7dslkbayahzhRZf6MJe
Y/CJjgyuXP5S8YBIw9f/c86iNJQwFizXttnmjXyK9zoxIzVO2WhIqJk7uKAK4E5B
itDaexaCtACbYBTrog2+YY4A2ab/yoUaaFQVQ0G1bFjAqzv/zBJTG7NWhEyUAnU/
fvmHNtml5nk+MwkSsc0OUJu3kL9EFGRb0DL6aWBRXmkyBXj/s0GMnzFG9hM3dmrf
nuTxZ/alFpRnlHKdvftZUAskyLatTm9REg9adqKiPAvm0CF0RrNhdRPHVp7YZWnp
RD6W8zizU5BJlJa1xGjhZOwvjjgcgn9RXPrDbTNCUzQtLM42c2gVoiF7sOAzKFDY
2R9mzUw0LkkPNXH/adhdsbl5OdfYznQzG6PaVbAxY+rkXiA1bfzoQZgZg/Cp/cg3
jMTGFEvL+6W8JahPYmKCH1Nqp5qVjittwhffbsCFCdh56ah2wUFVTTsjXUEPyMqn
936uNdw8xnJ8e1nOc/sAdoZlBCTzV7+LuTndfHlh6KkADZK5jNiQ4FYnC5yOXkwu
Xjji0bsFOVugtkvTazq1KpnM3EUVtSoHTmigEEEuk0kR8zeWur9B0oK2znMEanIR
Wtjsmzo1V2acWpM2Z15BLDzRz4pFZw+3gUa/cRj5qMGF4s490jmHhMKZuZJpy0sP
zb9KUUpYwlgl7s9n53fHvAt8Tlmpom3dl9W4YdImaJ4A4sFCmmXBUqXV9Wxn1JYD
JyQ9pnJRI6n1smA898KgHogfJqc10MI+HtiDSayEGaRzSmnSl89P/pYktlNrPsm8
Hr7ODKxTDlQfh1Bx59o67OVumRhPDoT5FZ8bnuiwWjsor2+Z/KjwuZbtg5WsiftE
5Jt+VtbTfkLa59qhN8el5mLepTfwp9soYBDFmc2kD9t5qqOTkXPxno39IAwLpJE4
JymB9c1hZG2aat55zjP+n2+uoaXEOui5hgxiZpyH6bSpnp0zEKCQiG8cjF/Q3eL2
TLquEo4S3fSRWROeZF7TvRpZ0jJf6zHNv4wmGMlP3d3NTKftBXV9TF5/fc7jhmTn
hWiP1/lT4YdlWhkazSWeQ82lFm5mCLOKBAPKtZ7bYJ4YLb4yFVwkoecBTbmZ/za+
7ud/i8/Kg8eZxxHHLn4q+C6gntinAvIuT87D/lFiOSKxUdcD02kksudjXNuZKkS2
y3eRegHBuGsMXvIFOlYo6ubo7Cj8W9BOtEbKGpopyy+k10BScuGmlVdlTq23tZZu
I75JiMil6llhELGQKoW35MxF/zg7+hiDOKty79+xS5GKTcowsFhuR1HiLvglw95x
j8jxzJ2mnrOCQxGqaihZwp/LY+LE/f3mqrSC3CCAJzzgbfxK3DqdwXdBawHpASah
mOezpHjSw+J2+kuBUxvTD5G1+aI3/1mYj/fvH4UNKlNIdqYBJDyEtLzLR9aC2abf
0w7ZDF3zY/Hj13x4sUw0U6Sadh6mBalzrG7o7AwIZJml6nqk5KCV6ZgGJgLsJUj7
h5loN+MHwYuGWfJ5jysPv+z8WIJNzyTV4VPDxxh4Jnb/R8hOP1ldJFt0I8USX9ED
JL6ZFlH8fr9/tZjJ28nlbpKG1w2c4xXJwip+0XgXKSPGReBZqlQzFBWOIINoWE5p
vGQUoxd+dsvmimeC92Jtu5LTKItw5wtiCdZVVCIeI7JhHEfJuYHglnQG1aF7ZtBt
7YxkvBqJlQ+40yOFJYVsWrEySxzk8FA8lPwG7Q02kB7YWjZ+gZBNATHG01HgfObW
wEZVG4qOk7H3OYsb09CbWbqr9GFvc4ZBcj/vxwblKkZlRoInb0IXoXiIEixt2Jke
vxBE4DyHtEoIHLPjcvZNQWOGYME0vyjcPr3na1XY9kC/W8VFAFPdAAGWx12I6mC/
Py8KHU/Tmzuvdy2BhRcueFJTY4aDNvQIirDRxDC/VlS48vg5sVrAK/Q5oJq4dpOU
ikyCRuI0R98IOJCuwzTGkyiG13xnn5wzk9m/RvyPre6k/tGwWg66+hNdrO7Wjbmr
YxTPCg+9MF+D+3b0MpFoN2tUYdANH5PzGTMOiRGqdfQRMeHuDiZamVQL0ebdjuJx
8pS22V0FfeXDR/tk7ZULaNZ2K9iKetn4W8E1ZWUZYIazejox4auni/pCJvZdU2n4
yfmJYB7NS9S6Cb5URpKgqJH7ZpkiwtBBSpyrI0xpdZi+Zd2MFXvRFF+KmBcGc/uP
um3dC/R0dzTi0Gm3m3QaZNZ1JrYU0obTQw55Wy7EPnt6PilvJIVB0ku+oYUIMn68
SfbSolgDqltjfbiWStsM52/xl/02FscceH8Zu5ya1bwBcpr0F6Nh3R/5/qZmXoLV
qJ7r9Pgp8hh8EWUWNbMWAfY5dxF2lDbeWL8oZ6lXW6ezwB1h8i1YWZXmBixgdcY7
G6Pl4Hlqx82KIbl/MQyjUrtGirw1aPu1Tr+5+fhVLwjoi3rDBmVQbJ8NCumDQuaU
t9wwoCkNCT3pNZ2CKUXnMG/ya3C/ea25SSiIrICwtzPMU1TXRpHm/LGo5u1vuAKI
bUyvZ4yv8irp7JUw49mBXJ//th3mzmc1eF+v673ybgKo73FdP9Ol4tQREDwMbXFR
0ZgBEp5cFmUzCY3noQsSurbawtJFG80ogo+bzDTPCSk51NwxYIEBVxNdz8XWS5OJ
JXKRMGzSusN+GQP6tAEEYnOzIniDbijNE9NzjTOKNvASqcdAqcsqpJoXTmbKXsBZ
NnobUUurL/toP7kywmRVnt6wB4beH2LF4KIF0rEKUXLm+ha7Kk/nW8H/H8uTLOTd
rzJ7um2DuXp8DX9FezL/ER6lkK9ngVrvXP7jyls2a83N8XWO/aIHqz7G/P9xxPEf
ZL2/heJsIla8u4T7PiCMxyBf0e/5miPCrMgH4UEvKWvJ3uY9cF/nGnaZfXyPu6mm
mz97yQwfs5m5gO12Ge5E4Qfbe77iLGnfEoGZiUTmdKeklnBj2Dq7fc/cn6D7Ht8X
z1ORZqP32zzuBcRjKhrVrvoGsXSusMdwJYHInqnoPkD8HjDXg0KnSmJtWqtZh92V
XNrIxsEJ7Uzb8xcpQZadBQEgpUHwrYovX3ozh12UwR9AUxeyZVU2Z74G0MSoU7LI
EhFeOLqEGHHCD6nC6NLDA/P0GPXTE/DbxlU+VBo6xLPmtfenLM/Mg+WbkIUsTvbU
iTkiu5KOzhP27cJUbpYLoA+x3BBUH4SSJlHvxiezAg1dj5Z7X6J+7S8WMS+V6NAo
PmBTtR93jXA0XFrZowSb7Mek3vARQvuvM4RVcqU5Dm7oSxxHiqf6i1Ex6mf69Ap5
xcO+cP4tU5YaU2eEfMJ9g3pjoTNhWynTzfaQiEqHPpQRYueIsT/hSLvml/DgzfUE
bTr7jHXJRWSSldU5HcCXh2bVanHI4Gxb0rH84a2NYeROyyhu8Io5pVaWQUTEHHnr
9gtQbYFlSL7UMWIL2nsKAXBipkizF+2GU3ZyPOREhVLKAmk10lqMn0OCOJX1gVZQ
phwrKgVv5R0zJgahZX98D3dezY5aZrV5GSeBmZwdK3HTaXlL7vy7Yv3UnPpzzUXB
4/YFQuseKTkptM+IldSW7+luRdIdMTnp3U67nVZtnWCKnggSORA7h3tJjADgDESK
Lcf2db69uEi140dwmd0ue2HVIuZpuYMFt2qkO13iGdT/faylOLJLJkjycL6eEyVf
XL8CPEEZA9S/lGPqM6SrpP7Ag5Vsckk54WsUiRsWMbM5h/oaRsJI9GY6DqK7Ur8U
rdq+HqcYTBMzCrOr8Wr91hw4Wwh/Fg9Pj0cTARP89wzl8nIfbDDTUK8iS8SIXOJx
5laK+ypoTrpepg1yjFtwbPDD24tIxmcfUprXN2T937buDbHax2HQZQVZkeNtoDMk
ZN4WHqcAElGuODGEhuqxX3+f7bcnyrYjHNudoW6tQhnBvkn0GFNbeRqaH+oj7Gg8
hj4TR+myuY82Ie2XnWaZGg7xG1l4SQw4P+6cqB5ttD13hYNNDm5pMmIaRgy6g8jA
o/YMWdPo8qe5eybWP42IiMrSGQ+gdpZLz2fCdpzl1i/T9QFwPKkWx0nu5nL/rP8K
RMZkqwFI7GwVOgnNF6kcWaHvmaI2YkY+C0q8AL8pkbtd/RPS7nPg1d24Ut24V1Ss
UEEoGUDSbfMRrEACFA3Q2fBjcbWfTgmr9UaeUPo0MXCB1OgvPVmVHyXFnmUwjacz
xRR58dQ7VGi09VsYu/fU3q/Q2JbvMud8UHCGH6klKd41exaGjRQVt69wt4OcnANX
cr59zPyEZbly12SFjpEMJlkWN8e/sz810026HcCvQXaheYagShQxxatMs+1cQet4
nvC4L/fJUWx9Dyb7Q06eXBR/Y8kzuNyYqDXZP+7zpGrGSEBm3v40hf1gRBo9MTp5
l8PfvaOoacUso5Ihp9ZLva6lSnyBpfAdlgnj/eVCVU+myZd47CWTqPVObY1jmWX7
594E5AKKVWgKXyo00zniLoDCEMAHNXzxizc0GojpycG9XL0SVXKeA1A1N5q02gxS
v9CeCcxzquI4ImICH1x71XgJntEnmk8J5fYo7L5bxW7ifohryTwekeX6zCy0WKl4
1KUz4IyMnAQtBx9922/s8H4P3FOLEzyyYmrU20zJUswtt9XGIKgA5RIb/pAnWK5V
3khlkysPo8vFtiaPLFcTYPp0oq1jJmIQjQT/A1/N2ojeDrjlY15S1FMIrcJoD/SG
Xb1weiY6eAuu69FN5RWqcLUkG9ultQcoaEJv/DoCC5E7/naGCMbeRO/xm/DLIUQ0
TxqGudbgSYlV5onHVL9avPqI2W0kgkXNxxtlB8tVzyN13+VUyFyGnoxVteh8yQYc
nHAeuDP1qDlC3QwYLVXHA6lzmRQ1BtThVnuDKUsIZxdcWAEAsuV4zMdeZQaCGHfB
usu7V+fUPOBSTVNa/oZcjiCU8Em1LuVm8/1xTjEnqK3wcqCqrfxEgmhktIAyERxJ
b6XZDv7t1EiIeAMxIuhbRBgmfn2x1Nj7+mp1/aKHcCohOtt9KnKSqqWDkusWLeiO
kYCQEmeSym9ZZsWD+GRkC+uFyB6zzH5I98my7z360RDlrv/ah2r+Z10o9FuEDESC
L+/GS0T7GJ10uArumEjMvTTBmxRuLuQ2lHuMpck2K/y2Ct0iJW8mExsovd+RdaTO
aMWDgbJ+pknrelGweCyKpcfWS92H8AMBLIVIgbePkomIleYSl0a2LjDsJytgEzbw
d1CXTtlWEhcjrLDlsDWzs9UUc2OgfOElqLMWAALLpBnaTghRvoMBWYKjlWVj1GPa
QDoOW0oRJHf8LbC46dtiQMzeR7Fwtr6CMD5K5OMwiXZgm2zTmgou9yewBaNaCXFU
TyA5aFTURWB8Q32zmmWTalDxA1gPfGwHbQajilYQlI/YXFnhptHK9XJa6ZxPvdNx
R+WKAHHrloAR+sgelJ6FNKUNfETJpNVt166eNxJT8avk3tOmDxAAXLeD/9V9LEdt
5IRjOkAYhxD0oYS9IdpKZDzt6359lP5CBY/qpAGMzmaUMF7USegHVrEqGWYd2rW8
BiOmWPe2na1TDGEhxrHKLFO3eOTpB+cmoKm4hElz/Tu+vxbHDs8Bh41nJy7cK3xa
uHtoeil3V9NVbrzguSfbK/F0FfPZYIY+lOYOBODRlGB2j8y4jybnkH2W5UBOEnu+
QtVZGLL9BBp1Bc9dlNO7bRgTsM/9s1R0l5aI+kaUg1ytaKDoxVKnVJLpVKRcT8oW
sQLszBIBXnkFK/NWpJkYYvbOHoyH51z79EHrcGRJrG0d9iTEUdr3blYg7R/vcA9B
Cd8opMSVy/q7sWGlqHsRYJKX9s3Mo6sF7MIoeC3tlzuYyp2FeXGxAeA0P7ovbpDQ
Q1mZ083PLiOitbHDIZbsHWu21G3bdWIv30nf6Goh9zdl6W1HxmjTzzFpgq5vEviE
Hwombd1uabyP+UHl09s2/Rf6RQkqKvJ+943h4jUsE0U/xak0rGrzh2dGggogwUAo
jO5u9d7JnGULwe27ECign39YhbusYy8OaVPjdNal0o8hHggmMqRTYjuJEZjeykQH
cUVXAD65lYvLjRtZayrzBediDCQAAl+BgGWiCXWNezX3/C2QiSAkkh2qnf1vNIYd
PWfKaAxqBjLtoDY3Klci9jzKOWluu838oMHLYsr2T3iD6fvJDxX3D+a70pw6tkVz
AcQRNceF349DJ75jKHjKrThZX1/23/FZ0z7uhzo5IAcvwTiVlQJYyskA4y/38D/w
gM6t/THuWGUDTxY5qvojhGYUfI/cYlWKcGcvMxyGOGONzYKLfTc+ZljD7iVKOrRV
6ZHMlvmiVvFVJqTC5OdaqSxjuuoCF4v/N9bkDyESC47WFbA8SEO03UyGYP3ckIwA
IfEjAs9T1JvW8w25LDdpYN27gcG3AabFSWyVMqe/iTguIHEItz7qakIAegFrKOz3
YVQIA1VHKtweDQVaIZ5W0wxjEXoU9P3SCWBHWDHi0XaHKWw8zuJL1OaSpAXM1ukm
ItnLTM218AT/kF4X+Hxq0cjbDNcLCtRzFlddP9jKKAldCLv+ih15sop9dtEXBn/2
GxshjJMzuxF7gRAi9aCTlctC5jZtcVU6t2cFwyvVayxHikNTr14luTzNoO5d2ebZ
wHun+YSQnCh5KSSCSsIwD7o4/j2OfAPIKxMyblNej8TMUQhtRUW2NTGcX0msC25u
ShVv/DxMfrfWhIQfYV0UPw2fAiEsfu38hd7d/x7Miip7KjyQhhOzH/ijq8nEd8RT
yr1KqMr/oUrBsCHbsJ7JFkm7aUfiSP1Rs2FtiJmAElxgZAHFlaA1tuGf2J98kXnr
0uTCLUjQLgEDyAXcxoUIUqRzLTYdvKUgyqhBCq/hVztJBWQVR0L0mYzvqYb9jldr
8ADFQDR5BMsC+/J7EDVYnIwO/jqd3c8WIlExAaaCUNPZDfOCkMDZfQ4dSCxkJKIq
ru2vEkNnVlfKj8ptu6ty6PpNtmcE5NSWPdTeb42zT4a0SQMqGmCtQg8MvHY+8uIW
f5KUu77QkaC0DS/DOOW7RR0XggHgNWsoP6DOs1l3Jhs9SIGcTjNyLoJnb1AMgxAj
AsQUubUI/tmYGsZEYAV0niytRm+u6K8Qq4PBzWgKFh16VpbBb9jVGM88Cip8oauP
usHXxE5m0b3pHz3NIgNQoZ6TQTuw6eV0lLtYfXz1PGBkRxis/FCXBA4QzWweA+P4
MCucn6hfYTod9NZ8GhQu23TCEM8Yswd6yu3wMH5R1go3DLCCTZ6+FCuVxwbX8dOs
a/3Gr4tEtLiCWqtH6u2xoA9H+qaXXsC+LFXEhT0sui/JVA+0n7PO3S0IXfjRLFR3
wpwgJnRYrvPyFu847g19mEMsjXGpvTaKAOqZLk3nA3KoTv+xmfxDDu9NKxihRnKo
FSFUEWx73uRKPGTqkR6U0uuPLiAvuE6kOAExB14IFXm3w6P77lZ92fGdZU6emQoO
gux1FnzMD6wf7Ac7tTeLCXwVlj0Mpq3v/4076QdPFda4kHOUsvVLSDW1sLxX3qjV
gDaEJo2CAH8FrBgEzLuievmtgOSOBd1Ud4E7db+E0J67So4Nzo73dts2UwYtwfEC
ax1SMYgftAtiM5TFMH8wHwszjNMXD3GlsL0n0aLUaJIpM1bY0l6GUSs6ISt/XHS+
TF8ASie664im/e9fT3obviBV1gtfy3nV2B3SEqRrshKZhVpAFb43hoUfkocFOeVz
5UJVe0vNzmqgO28oxxgKHa5Fq/hNYZP0Wy5CdZVat9X2ssF0UU5odRVQgvelzVq+
37E+YHS4L5mLKYUBg1av8a26QNA8TquEFCvEgByjlbWS1Skeb/89GjUFH3MKe8jG
6M+0fnAjeEWUms7+yY0R9D5BOWfDq4WWdq/78MePO1GEL9TFlJCoH3WbAHorG+3j
4bDFFB5y8TbQR5BBpj2NGh5Xx/aBqlqyWHdhCfPHHsQoEY/+h/oiv+MFtmzsuYqO
3osReQ46d3xl/TRDQG1HR22ij8kBy+l3RcBgtsgE5257kK+MJCigAjUkWtjzvGCM
XdMtJ7YZLMzdQUNennWfLt4E+VnY6qJE9oZtLUL9ViL33u/jxmGpivnNRy9Q160D
rfkdX9MGCEOJaS9+zyXuE8XKI4S6EwfQIe4wuDFV8bfrZI6TCDsWwX0abfvH7Sx9
8nM3HGdJkgjhBUAPFiv+AkzYP+Hk74pwfqOyKTja+WjU+Rd0c8qdp/yP/h/DWguZ
pl5RL/rZ8WfRm/EGUU1jYlr1rAjisoHnXIymyiHUYAvbVJEcsjhPsrZRYbwvbQTl
qdg9uMOSDKc6fZJirm3EEJGiV3B3RtMrThXQoW3ZbuHSX1MRFtuAv/r/g96gFL+o
1KO8GLlOa61KnNpy7ZKOSAqPo1eMPcc337WalIdyPFn1XG8CQwISldf/y+Csu/tL
Q1HWDm3NWq2eQ9K+B4bq0JafuSh50fkq3StcrCTeh70HIfgoUQgISSKCuR5Knd6a
fzsrOG0T0qYkjnpIbCcd1emCKoNENsXs5BLzausf9OtDgr5MUhpq05dAmb6P7HTz
YHPq7gfzzv2sPLQTSRi+DC8iogexo1ugRCeS2ykn//SjUfD9g0U5OXtZqJQ2l990
mB9T8L4anI1WQ6VbmIFXmoR+iUqDLAvYTFmCJv8PKqOGR1Zqk3RnuoOX4qGyXGY2
TqCUoNTXXYfQUkDIAgUCuYlqtL1wo7+lAO6yrPijzSpOc+4pvaDlnVHvc4EdWkAr
kiOQIZbX4ZL5A1ovztUA7N9DVVnmyKJRoN2nxTthTEtaqujXXUhBPBGyyaDpscbe
Qnnd4g2IqnrIZBXFDcYzW00DkyZRoE+H6Ia5PINvK22LLtDEj7JgHMgScYPKL07B
pyZzsfIzE9ERfvgKMUEUCJXOqrWQ+mIxZFM4qPtLHYSEfsOuLXhSISOqhoPW3jhi
CjM2yN1pm1lhUeF3YbbvayShv3yd3UiEUvZP91HI5s1DkidssJ6CClxbqBao8s1x
DI+zu8dn6ofH2BkZrUKvidGu8e3SV15eJzyiUtPqQYskMZvDt5su7ILG4BCwtVNc
sSehs3lT/1xRhvtbMU477S8iSw6w0Y/JQDf4KhnwZkKSgXj1upXeOW53FV4kfV2Q
dD2PVPio3ZI9OoxGTBXqMW9eoMVu27qpBkO+oYCDVX5TinMjv9km6KNSboJ6BbpV
iya/JOE0//HdTSvgOSUTaH4BI9tSL0HjYx4YfVApK4D13fRhqOwVXBGpsLmv26Ty
bv40c751R1zVXKo58cJAFAJs9FXVz3w6yukDY7ZOj0K68r9HCUTn+kd03z+6cx8d
mNBphKuwI/F4l+ClGMA4IggLCmOLPeuDQcufKnodixv9Iq/GopjmhoZpA6j0ofPw
IyjhxxSFRfhMqAhAotEFzxSBEYrB9UPOxFZ2b3D64lKX4JKYCAznrg5PJUuCzsOp
QteobuwcnmnPbvm6smlLq2ThHCGEt0ZeMVnPpE32S2vNJWANvtV4g0s8iPkBTtVu
mujsAybRNxW8n1DAKJdAf95BpXMYfUdMTE030B9pSYMcVMTrnI7jDkj02IsFKlZ4
AQOObRs3Ahw9nmBYZ/l0tPy7fwfGaEGms6fzdAOeWK1/wxTqgECgVU62by/ypv66
Kyy3Jxz/x2ZEXmxBLdY5mpVxZHlCjfIJNx+QoAy3LCdejKialCyvvAojPK8Pddu0
IfYW+W67TwFO9yzEbkqrfb6FEtb8Yg2nbZxXtqjnovMGpCgrRRfNXBh+f6cUxK/a
TtoPiHtEu7J4B8wYskXkGXQiwIUb9zsL7QxSB3V465EapAnCc6nLrFgSKfPE0UwS
5vY3gyt/R3oJF1xfuudrscigCEjm+ZVvWy7mVyJQfZlBcv68bT3U0Rc0cNFOaFSx
CB/iov9dF9VRPWnSnPc/+MNHnnsKO7bKTOmXqqNX7OzvTfrP7NXYDnS7lkL84emm
ftya1+SZbqazAPaAyEIQIyrof3akKONYE/CAT+Pp3X/ro5/68OlLAZnYqTy4GZ3H
wqIBd64vu103jyWh6HoyLutWOFN0RyqaAM5ZiKttRjmZ5RsudZzGAYeV9b7PT1tY
crKSEeQnjaPLJ/rjMfDCtEs/dnC58eDejm6CIaViLHo0/aGvqlouCNJu0NxrKtNy
JW2BFmdJZcVqxj99tJ65sp1Zn6JskHMCAmn3Ex+Dv9Mej8XEVz8FktaOcPDUvqlq
kycXn7NKs4hflvnKYZ6wr47lpn0YEmdfnp+76AGUy8wcoEtIekqzTU9Ikd5VXpSC
0HBKNVTXAO5F4tpIKE5mRxpxptlsT7b8LZf2MAdodMpAo/UW2ExK1X4348PHuTjs
AxzaGIcV2tkMBTXD/Cwne1viwHGREfGG0x36zsM2my3Mv653jBOwOp9rU0dvtCUi
4jAUFqsKYclTqNbQXjeBiaSuEGM/jpb2e27XAR0LV5gGSRjjBuTNCT8+iUsnmbha
/oQnJSJ6B8sw3cVC0owXkNU5Y+4HFzhDMOlZq87H9rbzsVwWwOrlBhUUSjATbjyZ
Z0V2sHysBkqe5IUO4AXPe+gJTWkWg9lQr/hJe/alohN88GkiZvbNgDCfg0OwM4Fx
+bSlXHKzLpYQsyCDbBg0vF4vxzzXPImkv9StWOW0C93ect7Lfvei0aJyptcpGtsE
KV+mRArRgOSuizKlgHiJHkZYnQ/ZEfbf8DL/3232lwNzHCRHNxg9XWyoiVfS9nWP
l+oy1lDmhvS+vzJ4JxxkUIQ8d8UXDP00q4Bv/y2TfO/ATD/KgaOxOdKPVz8Fo8f0
G/wyMxB9xfxHd6VKW5Tk/KwBp1sDmcomiSiJ2/vpIZIuQ0985Xgomf1C+1w0HvuD
8+OTFESYuP3o6uR7CjOPXVAioWjw6d3J36r+MrxTiJC3nyKu5EVjsEvsz6phiLsK
W1y7uXHLrt1M9CxSESTK2UkrHvYtmF7TZgg2T8jcjYajSbLH3YD1RGljybOotQxb
NUpM9f+EDZxA+P5pekhWsPG99OUu1H5+m/otia0OuMj2jQ8p2Q2SLz75wv2DLQOx
o5fbtu+gvZ6YkNvPO506KweFM/EP/EtiRbVUgoX85b0291Ah+pwlSvY0o6/0CAW+
x6h0La5zN2UoGIfyt1Cl85KxOksMCh5z3nCN+uUEP1krW2zZN8+4lqQ5JKBUCPYh
giLkj9pwHVQ/1fxD2htpL1W+63556oAZKRYFHRPqPOz3q+CwFHh1cZVzld62Fn/P
NHlobwTxtlkjC4PWw5Fd7mYtL9HmmKKSYrjWQdpymRav/xwsTNqA5LvxSAyI9WGE
UrjZdwvKXOXUxi8FxZe0iGDxRFEY9sOzkGojzNZXmbd62P1rclGAgnodNRcqV5iq
yInnxVEak2ZqE1t2AchmpAg2jqZ+OWxfm5RRAOcV90MRJoW/8UfG/fqRKCCVN5Gz
SuJVa6Oc8BR9zkdnrPrWWs1nnSNwlOjG0/+CwE2E0O1d5sduYNhrFr15T1flOxIi
ZQqac5hr5EZatTfoB/g7/mNEQ/VAMKsGAAjo7qwnR2IM4sqyNcgmDMtdwNlQH+9/
8aMqG00FPLhec4v2+ydJxAlfcJI+t3Goy3fmajirJFCos5K28ZZi6mcM1crTF4EF
CTWXD3z0w13Y3RKSheKuPTflrZGPdG4pBd85ethPULykiAJ5gBjNnKVL8TRYmz0n
GH+YfxH14XzOum/UfwPAsuv4UAex9PETFos56opuEgWZ7/k3OAINXBRuJCF1oCea
DXhEUT2CDM0fLo9ZY09vmlfwKeD8JXAnEM/tgG+cXIFAYSBcuJsv0ik/AsOkvK6V
k4OO/f64xsQqaoKOYw/rAwL411HIDx+HxuLOO1zLvXX5jeQVz77b7amtul6hTLXR
y5oKN+vWqb0S/7nMWR1T9YHsR/pl6xaI+XmNd0R7GCMzscF2ycbkS2zRgRqu+MkQ
FftbKKVyKR3cNv7GIWOxD2PD6cHPPnAwNz34ZTJi0VcCQzP+pV+552r+KyWAQ0xG
fSIh9+BhvHHGiXiaPbNOtbYbEpBcGbVHOm2d76RAnAK2JwQAUrEkpdiZ+4+QhHPW
ZDG5MdVfPA8oqRyUVIuRnFPkprMDjpfjY6cpdguxSOIW8tnTpFFOPD7Rmf+0SfyQ
zYFX1TUkUvquW49ke++RSJdkV74xEZnuUQ8U/te+zr8y5KmaXbVdaqvKSbqEzLlN
EtdLF12maViSx9Txpb5jcQznGlpU3bWdsE20XT897tuU88ZgNiKCCO2AW5pdMC86
0ChLBTtBXzY31VVkKW1BfljNAGltPB1+X5d8VIDBzWdv+KmrNb1g9hNzc2hfxMoW
Cr34o8t2Er+po51uLlcsAJRwoQVFjcI/jRUMuQ9kVtjNpE7OEyOsW/j3iMCWBR5v
XNCAgw3o1WtxBYMQQOhgqZ+FAcMYvrH33mfVTHLX/w9XdMOHtS11eBMSz6+j4nJL
ptrc8mrHgkVOMkdeFVoKynysOr8sRK1g8XLsvWzLW6p76YMlYsaMdsJs1Z1mdlyE
Gj9Lju1cCHOjLJAs5KgKCcmHOj6OY3rLBE/pBRqzg8Q004UhHpia59OwzRU2Sjdh
1xOfyI8tKpalmDraQpVRokRorNBKxBxatEZhzT896SlmctlCcSo0tV1C8iKcJtYy
mHw9FCmB+wJ2KH3LYdRDrznq7yuAKXQX0BDlrz2ehYSqTbaWxQenCq2NltwP+Az6
L0AMWpmnV+1In7QHxL6C7AmTYpFnegbetQBTAUGJa9EBl1hCWHdxo8KO89hOwFwD
NTXATvAbHwHiu2YiuSOhuipjLFlFlbn4oWBrw3k54IqfA9mtboNX41uJzoDz1SZ6
hqbI5dCYFe2yM72S1q9270oCmANLWq/Ajrsm6Qbu+ewy3/D4dqV0gEGX85nQIh1W
i7KAzlLqO16RurNfX50T7BXOpOuhZ8TpOHKqbWOMLp0yq46GeF9Sy+tw9cZR8kmk
YafRClOtL4QGZqKdHSKM5d1gcsMLBSpFyTgmGaz8kRfjv745PJsuP4pNoQUB3/KN
HGIq9BrJqu5p3YOVg/pU4bWjXcUwfQGcqC/SExSxPjO2vvEmcPTLCXlzepURWJJK
7L6+5iDj+pGH/eESECggmskdzcKnhFXmktm3r3aPJ/eHFwSN48ogxRr4XkFW1Nsa
AWbunBTHBeubevFOOl9CmjH8zAS1RN3V8bTMKX5qwJSvr/MvfJnnelDGu5kacWYF
ouITztXsiixv3GZDRN/ykjn+29IFnTeyinhJawV/NwjqcFcClsz+3QJNKcviniYm
XVjd9J9fYQJMux2/yXGUj9UddCbqbKCNwvd/B+H8wPiF9Y3XmLGT/9X3R0ogAuLP
dziqh70INrLL2qv8SFpKYmtuk8RduqrITwEoYxBg2CcncE6CcbQShgV3C9ld9TpK
J/MAUekOC0LchDlZdh0YseWVLakUnD9hBzhI+Too8MZKGjUbDmJMohpgIU/xY83L
dqS0QCiyHMfG60UDSZdN1XlRPewVVyOz7qZzbE2GrjJbdzRZBC+L/IQhcyyBygLZ
nOioiCWE2C4Qkjvt0BRtK8dGln4wBtCrsjEIiiFBIBdpos95Zhq5D0WXIYJy2QGY
C6tO0fsGJXLOg32RP/oqOQE02ecvNr5mF5xxmsOzrSVwA5Ep+N1C6fkGA5JJTMIq
jfdTzxsvHihM77dbAP9nwPDVD+YNIOV4Mh8Z0AUYas48ndHYiphIz5ekcr1MMiOQ
DZqw2lqxJady+2c06rPXQ6cR3YNzixoEs1x6f2yc3P1L2oxsH8HJUQMkK97osRDf
WPokKp0NF7mNQmtFsgo2iPVQKJFw70SKUqH7GoHurxisPU6GU6Vr+u13uf1cSL46
goFuiI4vISoNiCp4ROsgfXskSnzOWPGoUa2Yfl3wPhbYBwmrdhSmipbwTs9JTXKW
oQWdQWX+avcuv/wRl72cIlRocp3ons1U9AWKTAlBquXMR1Bg7nw0ydPEopi5Ppan
FhRMgLDZirUO6JE80Kyg0nmMqCEeVrfoPeGWWdP56XxmR+oQlaADoReWTNyBFg+8
3fEpmOnGS1figAN2PRtalNTlWKjkkbGY8gOb1AHke1KEZIgOaBUlJvTzI7U26AyE
ybRwSNX7LW31bcZw3xumVZLksGceqK3QIljc9mCm5gEqgOyk8ngAjxKAOasBUkU4
JkiFASuLuJ0SfoZjAEozcwgY5Ew13ddd/Zn0IwZYOglDmx+mJsOtbOG9ArLKN5u2
ZaCdwpIVWldFOUth5GbBJzlV85MMvNh9NDKe3L8FXfozrrS2UttDksg+l7QdIScd
XKeM36AaTPmbGKNokkpEYJtj6fVb4IoSZAsvLrjk0+aWttit9p3suMvp5yAXcwib
6N44fzaH780PCdUK3sUtEBDoPXUMSZ/tmj+Ju/yP72qvbgMyw+PMfqZySnN4wl5D
aRIebjdQZ1l9VGFJQ0ltnTJnnMSQca1YmFGkfmr2fgBjXVDiK+hPm79wHqEaVa+N
2gG+00RKho9iqO8YdwMEX3o9rd7VQ2uAQAnvK4yE8CZJVU5k/SNt5gUG+5fw6cSC
470NGiXay1U0ZVIPxNAEpwuLt2nFZLK0PTty2zyUn99a0VP+0vATsx5paT4/BP7+
m8pZvdrDqp9yWCDPFyKMBGIyzXrUJs5+r/lDiftiA1991ugl9XkD91LbTL7D/H4j
QTAdymc1WQg0P1cu5CSWkzsRjK9dIfdbP+bNL4d+s4SGIzYpuLfYVxCImVT3HO6U
vc1e3opg/xKE9GCkd/U30HzGgF+Z+MIJEEQSfhoorUwAWTfz7khYYxXzM24JkJfI
w4DjvInSFo4bWy6RiA8/9pKZu5XuM/Fzqyz60Uv9BokJk/uVygyuRI+H+RgzC9Z0
34JWnD3ku/f0eQOzAcnsI9hODtnNZFpSvv5XdeEYzrQI67w7CJ8QnIBLjPVGhLH3
nwG6OIkBXriAMsh+LcV/0WaAONSNUZx/+b4PUPnbrLCnfmi3IS46DPsVo6emPGPV
UZtMQ75VUWIXVgw9+KPXIQmuCoHAQpHi7d0/eYzw+46SKcGwfTBl31Ab+8+hKjKC
5eEoxQv/2WnGnMOqP6ZKcY6Xu+c4QfulDjAL6pEIu4/py008PVIx9xS+ut/9oxZP
LLYltCXuen8UoPbo0JaOku9xE5YoD6TMjEClNX3S0RDLY2SdIS0isZlhkDNtZ4Xp
tCVfyq7WNq876JKPcbc8EJgf/xFA7tO6u1O0oAlTSAr6zKACBRkcolp3RWjYbded
mnkr4EN6JKqnAQex1TGssFC9IM4zerhdJ2Sfw5jdCO2DbnqprQ+5dzt4rSABf/zn
bKs5ctbyaHDZY1joLGN5fhAz89wqc+FC/wGuN7CCfbmu7+9WPenH9pCLIQGjO1RC
SrltdrCxgY4b5QkNV5gUk9pciT0AtVy/aFS5uaJaQ9IGUARU8GmWfy34TIeudto+
r6766DJuIE33lEpHLNlJjC4h8KNz5HHFdLy51JIh/gWknv5nYEBiv/NjsTvGvnct
fx1krxE4iu8WurjFpGS+7hFd8Fx1U4O17bOhXHfQVsw6lEzKEm1NO10olhoSke2D
JY279IC4Ga2l9KrIQwu27VlTxK3c86ot2HnTGxHu8uPwbLyJ7+MpkjlhGB1b+An2
HRay5fNasPp5FIo4yJVJigBdj6t7/XjVKl0bLu66PmBPzL/rRNtCayUHYyX/c4G4
OlkDARf1cB3cPzYPA26ovIp2aZ+LF+HaYg3VSrB3oOAp/mTdm5Quk3dQYcJHcI5d
uJq6TH4HzX+5YtYNJop2/u9X1wAjjNYbvj2UNZAFu4t8TWjNkqA3JsLJ+67xzls/
a1Ly0nYXQoEtnyUVLovJDhCHl0TPYh0ri6lihyA/srdYnM1G0fgJnJNbnLChs4d/
qBPVsUSQLe79yembLd+nUBuJJPdZdSLV8Ln7JUfSLazUSsfHjrj0PEDnXhxJ7WYb
MGEPvIWJJ5Lr/lInUP8H4aiyIsT1yJD7X6k2wLrD0oVuMPyPntJX08TQdfUSCEv7
rSvZ42jVryJ15gMn9Wr6Tmhv7ignTut6lkCVyG0pAo72rdJFvcqlPDfBNGLwq5SQ
LjlGRBS0zf0pXJRV1uP/Yk8ZvQ/0Z6fi8zqe5iLDsng90ByE8M3JwZRA3MvoXBv3
x5gtt2RiiB4pO/lFoPBUylXWI1s14DGnITppu5HXC/wRANgZQbFL52PZTEW1nDuZ
5npLsrKL5/38raEECsdBffj6I6WGR9pe36y9gLsCncmsS1WpzUzn+8P9n3n11aCY
1mGVjQEi3qrBlJjC1EiVfWF5cxY/zpLYboXww+vLY063BtvJr7HpCCkTcCmhQic3
+uYRkNhdYiA8ojoKoy0m5Vb3RsYTgmzrX8n50l2P+50FkIH2b5+508YCTTyjdhG2
TLAPtpUMJPqYwniFwpHctZzgby77FjOHandkeuNgCw5gdEkaoCI0LnkXTvLxTxyl
HRbO35TaBFBcDEFbId1Ul44X6OOBhJnueclfF0/7PRBO1bq1iBYeEmJTShvvKNDZ
0Kf14u5dW91GqfqR+dWHl07/uTJtixGvT9AQG4pGOkueoADKSlZouyJuWS2Yvm3Q
A+b6AWErsu3tbjKONEi9dyXUs7gT7cGSadyKhEAqTkpdvKp3Hs/CjSA5Ji4B18Fa
nmY2vqqJHBMyolRPb5ZaASAz4IQi1oPzaWtH2laKUbkr3XN7X7vqpcLGPd5M+Jk4
lRbhzjLnwrPkforP1uMlJCVVd+Ovz1ef0Gj2Zx6aiT57WgPDdjDJRXSiJrn5iL+a
3Lh7fqpMGXfZaqZ2NIil3t0covJ3SPYaDIiMIKYGPfl2Wwo8TUPPkXqkg5OrMmX5
Mx5ITBs6Vh0OVc+SXHR+k5uPCwm87VA6ledYoFcBFRpOmIh2iW+MnF8PgFulKy2d
dmRmEv0NL38tlAY3zyMBlYUgXMfw1lZ3KUzoZFjzjQxH4sMK0op1No2nqCKy6Dy7
U/AF0PwiGRv9RSH5IBvBVlL7ucYnC4+Ncf8KydxlvEeo7nqlLOKVqJWtSYbBMmPu
1VWddyKZNBKaQaT56OPBnuL03T0dTJEqidmbSFU5V7yaXjlIVrQIXHlgMCv0Jd8O
7qoqODJAOHpkAp8CEVAfMOCefNhMSYrv0DckeOUfuidkOxg6aYLiA9B3sb3r1Oun
dIzIXL15g+VMq6Kixpp8JyysiKfb06IlEmu+W8jASjuyDrs8GxtARrp3sQIT52sk
Dg6p2pENaPh9dBtI+7KEbol9TRo1VYyRlUZ9b5+fSmdsvuyegYRf6ufrIySFDN8t
bWMmjZC5vyN1r1ldrBIB3ojqiKH/wIN+V2wKbC/yEsoJxVG2jdZQdFKHl24O8EGM
lLENek0jOm8EgvELMNniEDYaS7ab63/ODpGW3N5CM/vUcgIgeeEFuEiFXbpCPB6R
0DK/syz5L5ANrsyV1/iDHBJvRLKUo9xoBIieIaIizwgHem21PXob7Y5IQxyNFoQu
yFw7ExRVrsSuYAjTg2Mn8fO1gliWJq2otHsFIybWfGdnwL/1mbGwhdj46BBl5R18
6iuMrTBuYWOt1RtmBCx+2G/YANkN40ozrCdY52M16YK2aGPXpC2J/Oa96k8+03Ed
Re2y3F7JnFH4KDpEaeeY9ywgIE9MKPr2JdemKGVlK+4sl/s7AUrORf1/NF+4FOYM
4FnUijdNv3X3m5OaQWH+xECaS1TTdEktAgzOBPp5E8V2gYyYzgjItge+FrHjC0eN
pX62DvpfmdCkyFomTPrscOS3YcantuRHNqu6N2YGwa3+ByUrOuI6Eu1ufPE0EYOc
9xjj1g+PMYWLEx2Dea7Xz6tTgA3zXXaW76af6kHdhk4kbEM/FCX7vH7688V5sJ5+
Em2GXUFvVpOrKtjzViTL5r/DwB3Enhb4j6nfKveq9Q+x9KNN2TmsQLneXxr8QpZr
5jWmD6vIbciyu1DBF8aojFD/VwWMPshFkxSgJpkXQh0i64epcrJP80cDRc9lvIdS
zqlxbWsACy7ElAk7qFU0G745HLexQ+7tKnIE1O51ir6SHR42U5d5he3CSRlIRhRF
VvRtMrRT0t4CjCOS9JUOoU0hkgvyFXOwSysi10DpabUWgV6qhCGOpKv9sTH5bBBr
sjyD8R0iMxBqYmPTOxN0XqHwuejzNdscv0EhkQ63fj7ZnuGt142Drl+WiRW2AlxK
YE/bv/MJ1bCGg9kv0R9nhOheGqDTr5P4Du9Qay2ptAc9q/e0jdr1THO9PGfcH3uc
kdkoZhIz8z7vhvqbS8FPZTvEcqPPJ/cBI/k4xCJjYLDlrYFgMh+/MstROlLndZL8
Nu5+b1zWV76vK28FqERjS5nV1fGiniSj8iwfscANPxD9vPDdVBgdIeUjdSFhlydD
fIRXVKtoWLan0GldOAK8CfwFnKyat3K5Pb4P2UURg39i44O2/xg5UQQzG0wzVHgM
uXW9FPAZC/jFUuCRO8V7vsNYyC+abt/T/xwtAn1nRSA442Io81BNa1UoUOdEySW1
KS5bARz/ZMCk03T3psS/Jp3DGuPJzbDNljIL8JAgCbdWrNlqDKYTd2DzmO/j6tOx
7kONz5E29Mb2vV4Eu8opt+OsWFnDx6vNUAhqzGbzjP8pT/8KyclxWm6ttVCsGN3h
h7tCUX04GHC4/xJV7aUD7GAxjYCNOqjWTWV5Ik61y+rM42GVOGLwvQlRXMYnpixi
ZNIK7IYAGij6bEqWo/50LDF06p/+uEf357Hp31MRobmGMWKMieueZNUbQ/OsRop5
aY9QOed9hll3AEBbaA9rlRTeRpZem3nZOB9lXbW7J4BfIrvNEHvrsNO/pMHLMB0K
5YYEXau/IJzOezmNq24wJEQ6tDTAN1viocz3tuO/8+hmC3FbENrC2qfN5eA3kEYx
sTeAGh1ObC1X9ePfWgrvZGVZynMz+0Xcsk+htdkI2Db+l+dZ9PQ6rvMjORpEtsKy
phaDz59AiVI/o58MEvQmMmBFmmFAN3SnzRcMRaBxegpgHRIhNNYQxa0fpiUhnDMg
a507AB7AxiJUjCjGT20Rrj0b8oN5LhcdnejGZu8zIk1yHIXk0JuoIzK+2buOVWPh
CW7HZigJ8P8up6764Ng8I6tWrBZ7XI1ta0pr+TAG9xf3cKLejJS70xXEfPL/EEoi
aYujWvmbDYzlQigrFU7PJQGv4RJuGprAWb6B+Fun4w1NPrG5inh/PYBMrMs5b/Fl
ikJkZ7+sh19P80woZEWfUZ4k/5fZefGtaGlbbgtiIenMKbVJr14juc0ycNZTQld1
4WtHz/WEYDiNuhkRYonGCiN6gN/aTpq5BGck7qpzig/GR6ZfZ8J2b8/3cNImJPlY
h3pFl8B0OFZqAQ16ULo63yKim39vvMXPbWXhHo7KGi17Lg2PAiyHjcFBOHAqNf3X
6tguuyDCxZ7DpxpB0/uboEQ6tzJlC7Ms23NI9tip55h0k7O5OT+o7TaO1Zl84XbG
RMFuaXxVbpsC1ZPv6xKGSv/bFGy8RiyHZ9jGHhuDIRiCzl5pex5pxffhsJg7usij
1/RWPVtZGUlPTfvUWbEPDZx8QTcz7VH+0K0bVDoRVrpqKLzETvUcm5Kat3m4xgVP
A+VnjvKVAQUOxU02ikb/j5LThOcNzhtVKdb2WFjkqQMi4wRqR4i/3w8BEU5W2/zP
TkvFqc2eHB++i9GXqp7WXAas+kI/3TWHMTqKRQKKEfbrncoaToJI0d+p7Dd5oQy3
gRVAEy2lS2Yp/YDAax8QccWCTAEnq6N099hn72DicKgtkDeDaIWm9y9LSQH8H0wL
kjsMPoP84kZDu4M9yHuqq1RgLe/CBcBaAjl+q20r2p+j9uQleWWx+lE3gm0lp0ET
ubrpQYdpvrKxXM/8GBvzcF82ctuDFj1OpLuOEQaXL0YzvcR0JFkkx8YIxPlymLl1
CMcplQaCilM3W/cbJSzC+J5f8yQ1VeE6r67SbV9hODChSRSkvkaF5NFZMu+t6jgg
Nf/Ce16MLLe3OoNMPRaAlrlGSIlHGQIYc6X/fUkoaQ18+BdeJjFypeY6oTGEbBz+
RobFgv0Rgxgndnhv1sFCJAcvHGJ/2hGWO6TIc/HOe71E4gwTmjAiVYR+bhbCfHPF
5zfKhiYvIwR/j9H0Yi/H2/TmzNqkq4XEuXrNuYYQzm6nyQzttCkHFU/KkvSe4n5p
BTSQp7aXWywbDdUg+1QNJb1Ur80Us2g+dZwh47STJnAQtbxxkJsqxAOKtLyjD7ub
s07LW8WvUneQFJQ453a4/5GmfYvuD91RhrHBIyOoUJNlhYqGrr492dw+1A5WYBZy
pVwLA670vXzkmxtKPcer/CjRXKFb4QgaTWdBPjZyKUPuaFGcJ9o2hGyS2RIKylsk
z0k7cBnh2wbO54jfpKbkV20XYs3nnCHMUQYgSxyeYGV6wW23Mi8XeQiU55P6RHuf
NCVYeyMmS0X3oQV1K6cERJryEJMWug/pUdclykyI8HhedBkfIueJKV+2BZI4P4lY
FaAWlDuZBkNDBmAe02MTZD+K5QdRV2DAg1KXxfGi0rbcA07PZbgKJ3t1+thG+1T0
lIsU1XVixb+yTpyb82NWjc90W/X5amBQVwn0WKQZd5DuXchcRziPQqQA13PNDbW9
oKpyB+3WXLEnwH4lScTrtKHaKIO2G6jwOB0PSMVouT1+18EIgizQ7T5eSy5jqnjL
g5T/dEQb5IOOJ/bL6AoWKc2aUNdruTUhLo1LRJ+vw1j8PwiUh0caWYc0RyHvdyXu
Lj8yLE5PJ1Qgm+uGatwrikw4Ld3T8SJ2pO9YyVGS8LOYoIxzSdIHr/uD17LJXLOG
tdwLOlgZki4E4qk4SlEifdB5Sr2YCFgHOpifKpCbAvdOEm6xtkPMjrjHRhwTWzuN
wm9uexRYxGlr6Wm5Wiqf+QW86/zf56YWels7hQzIi1CwPYquob9Ae2cvgiglwG0X
cP2dhbTvKLc5daPfOuYV1TQhsynCDkmSTT1Nrzgv1Je/nQmTmFFrfAY/c0UFh/z4
0oTb605P1OrDW4XcPHAHZuM7opLaP17RC/XhbQBJmzB6gOowMN5+04uyA0SdLpgC
yGp5MbhGMMRL3ZyAUAkVEylOmdwE4n13U8Gp3t/L2VEig4BriPUm2Sx+E4Fo0TM3
JdMjQaWjLM0/AHzV4oVIgh5aG/OjayX0Gw4dRJgREID2pXZ2cODvhIFAxR1tfpiL
tRjZVQBgzEubn/k2xM9UyhutxuRqnYr/YPdHu1Q4ltdnld1DsqODxGvjrxF44PTq
amNZtfgaaXZ/sgHsBwnl1SGXtFJ4NnrvUqCDNMfI0nkIOHW/37CMNGUcHFcqo+Sq
bERu8v7blUwtwXgnwxatpFf+hGtSxh/dNkBR7KfPKwX2hBiVdb4gIDJXvCVo6rYP
PqRE0ZODSu4rGEeDNv/lsoj2DSF9BtJ0BAmcH01lBNQSRFz5/exik2mc8UTyN4Bl
VGLo0Ag0Nm69suiomA6afYqYGVGJVZhzRwCjLtTms4e+q7impNIkfOewXjXMPisW
djEslyyYj3c4csq+wB2DiJRex/8ptIJ7xvcwzyNn6Y597ATBYyv/g0VYv7bE879o
eZsGigFkZ1szYdajPD1SF2HIoaGF9huodsvonSwCxej/gvvSq10Qc+tK1qiLtDVY
xQ2fA+IUmGnT0+VxkVGOOnXasOCT0yjkxAYc20CHz+lN7K6U3tE3PW275lsUDkGB
0J0teu+5wSolCU2pfr4FfMXqCuzk90Z7mwN3VzBd7UJozUA7P+bQxLZnoVuyqade
JF0O30ub2zaVH2whwYfRTzO/JSehizYAgF9bsTM9hHZdKjVNSAVqX1bVHXwRS3pe
2oSh7LvTCQwQvdluVfKGoqmBbJm5sh8H/o8qpMjJHPn2Sf/SVCIuGOPFiZAjj7Ct
hwD51S4KhO5M//wryoiyCRgWrvY0BH4k5fwjD2H3xS4pBcKf/iZw0ZfRi/zh30gE
RdJURJ/LaGkCNcKyx4zC3f1+ySHMA2XhzJUBtOoz4FBq9C+qilN6O51wtMfhA/MY
IpNnsoTjgSU0FT5au6W8eoQocU9WdBtsabBXJ3UB9+3Z0epCie0mixuIxise0qTd
nK4nAcky1r6kg9Vx68zS90l+XhMMD/DCpilg1Rw0lVyltWOhBnS1tCjexNOW8Wv3
dqSBt0YlRvVnuA8E4ct58MQYolyHqj9ck+Y7YbbG+y8hNmzj7+U9KbdA7kbNvkg7
gb1ZetOK0qG/5R1Rnji95/mNGsBk0kiHeaImAuDBXuZrBNtsUT6GsJsWyR5SqqUK
a/EbCi75YDQhlbsTYBkivlpkspglp4m2T2fzq4u4AyUaHoTOH3EAtkIRiMQScQkN
QaCJZGPL0gHJRf4ICUYMSP0kA+ORX6VlAT/b9O2audcS1q8ZbhztaKp8v5FmkRIf
xFyNfdY0fbGj5Q0SXMJSVtwIqKnRdT64ijMIIJwDUvj88k1dEafUkJxHYdRU8PUG
PTZfs6fGd08wnwCSeMp3bmqoBWINywaCxv0JMfDgVCyzMh3zm8gMGpUK5z7QNS3V
3BDMiMtWmmAst8SIlkr7lPn2sf0yLsipDvsO+sbwunnpa81bBnl/fddAmG/fynHe
MqiBAYKa3+Koo2EDF8sPbjgSmOI/V4YBxFeMwmWj9Rxsq8GpQFjK7lI7InyFN2Fm
a3DS46uKSitQgPhvjKBthpRI/ORR/4lnyF39TFvtm2Yo9DXX+KbhieNB84BBeyBf
mteCjVDG8ZxUaFJvCwQEjfvRVidCSKYU7mfUdbtxkidRZQQwIYsKCQ+Hg1qv5peJ
zt3Ye+qr2O5mFMT+SMzjCQsrcq5V/OWbWkCuQN+bDMse0w4LnibVlh1CG0rPKmiK
zT84lqFr+yOqHK82mK8bhVZbxTbjA0cCoerDj/npBTh60dKQTCFv20y/gaKw1mre
xOZZ6ZLYwMCgKXMh0REYuWX/d4Ge6RhPZxeMVX6sJf9nKErJvMw7CRbbq2xTzESq
Z02QX8994fljIzuVyj7wUIcpQIuG1sFzGbekuooYL2HxXpcfByBLYiMH196SexLj
S9E37xe5yF/LfDMjS5rRUtdYL8zmjmcI8YLIoVmg3++AfnjmCl9S2b5w0feSpjY1
tbQJ+tvWUynxFZpNRm6+kPtd25G9fabd0Jphb2IcTEaAqKFSWCNMmXoRtKQf6A8x
k1AFkpP9e1jPeKn0EmpQWHvF1X9qyWyWBaiFVjjZIaV+Nu5bxa1fYMB7oV926QVI
Fmxc7MOQwAmCMH0FOlA4nKY2T/fieoef39XhO6IfETnFNPGWxskroKnAMZL04t1/
qlHIGGxbC5bE0Sjzz7m1mYOuK7QrFqLTemTvmYFCcOV+f53i5jyY3EHdbwi6ycdJ
dIeg0dcjjFW2LwimRM1ceWJ4L3MnpwU0hMC1s+Inc05vesPCCsKq151Z4Dhn9BnK
9cE78DqWPWg4YMD3M/hYveYtamQHPgOnmVGdC4nBwPDvsSvPK1TLnCpagdtaPVth
xAkdV2WShtyZnaiZLtymUVqUaTqC936a+Xl4k72J4LZirQU+tutVNq3OEXe6gDf3
RyreVkzhtnfoKsg7sZ8j5dwr6krOXB7OAr2zf/dLdEG4SN3iqz0HemVtgilEWy2M
fFdvRJgzgL8BDSRRvybSJc32GymJQkx3XlsCUYu8LSsFcGlZem8ODUcALc0ohn9u
V1GlVM0kOvesQlH6kzNZtRgZf7vgKB2bi8RV5Kh6ZIvvZ0cBj7bTieYqF30it7zc
fRJy6mLAHrgf2B3bXXD0a1Q1u84FxlB1TRN59tOVYEX/LPmbAy0d/belwk89NYhH
0ZuxPPMR0iskt1s/ybFt/s4DpM4c3gqCGCKTeS1pJurNrBsbeLTBUJqUtbIi2ifi
ItsdMCCTnJoNynds/zBpFaiRSLPOAn4KRTvjFmP8ebkXJbZKrlT6s10OiTcE8a7c
vs0LWwgw3F2+sJw5fCQi0sk5fdeitiCaYZJ+y/oos7bPiQ7iWh7O89tFmZ/urWCa
6hhg8n4zRkrzYBjkao4iwbf6S7N1fdEYK8OAVQUFevDlj7kI03gAU7vpLEZIaiXy
NZOElVLDzaUOY+jsTwUO3NpJiUKTw6J0vxtx3Pvw6nDqS+13UrWLIZOD9BG7w3Cw
NAfzPsFgJ4Z/ZbPBmWt8Pumz0vYmaZsznnYIi+NyCSxruiWqhID8grLxOKcHPsW7
ZSSepwp5tnwti7eqtg4QcQ3VXZ+eHzc8/P7z6WMsMhDpKhi9W7epcY1GdjCgFb/H
LAvrKjYvzQpoPKHwoez5IRMz7eipw4aGZVA6DoN++QgIwCZF+8WOiTqynQwlm7rX
BAvNj3awgEnpqysKRRiMy/Or2YIANrS37owwBFSCYO7JGGuCh6DoFB5cfckLRrU7
uwsRzi1dx08zaH+9A/TNIy83GEY6/Azx/1lo7o14v5ac53THmWGD6TmBMxA1NUwj
V53sGRYHW5rqgZQ3F3JSq9fepGpCWwigb/CjEJUwQ+5JdCeCCuVUKJTT5Rk8qQyQ
ZzWHrxC96Gmd75797PLAE74p3+nqzoza1pzswBhsbtqXgi1IBpOLMBnxrBk3k61B
eYHaYzToh655i9YXG7vVCLtOHUm6UyFxNDtqob3RCDdwGoGoxKv/acGB1i8vtivU
hbGm+7OsLVzxHNyvxHBonQG5JFEUcqilvyhYzKa2cMU6VzPduMR1b2mxHvuUFG/Z
KkCxg4VARMMMObEkmKtSc2otuNXAMuMJpgP4VZSIiOE0/1q0KNn+7EG+kzQHf4cl
ummeGzLu1tFJVXdZlO5AyftRunnJ933lA8B/jP53OMTs5che4R0FZ+jSvYsShlWx
BdGPkLgfGy8aXOS1kX7wZrdLkyTj9vjJzEdMD98yZJ9OmuV+qKq5pvE3cWvRPHiI
YyT/VD5XVdITxmLh11poK4rtwWHH8wJ0b+au4nrMUy/9gGUMhhStO5WI6MkJBzDt
antu1jSS7uSO6tavvLPx5jt2ASELGGl90S8p+MXqK5WWnd4NRZK2NFoBfW/lwswg
Z2zCCctbEYANZ3KI4xn+vjjgcLDQSCcGrsMOEh6UpiUA6IlRIAIRH0jF/PQesZYx
snDnp4DQQhR2eb5Zt9HMQrA+f2PD1bh16y5xhpMye8U0b1btb2GqAUBuRzafEsSF
j0unFf8cRGNtji7JtesI2zNURUVhoRkYHhoJf/Vd4aofJm2/qTxlWdn+2dM+nST+
qfT4mFPaAa+YYLDoZr6LKM+L7gaFNGFJQO4Lqt9MgPNEYe6AArMIGBYkIecLnrOA
O0jIbnTzDfl6xMyOoskTw46T4swxIf3TGTd2p8285/zotc0YTHXpIlGaEBuLFhGb
kb9XjALsGxu7wuTepsVbsCm3DhEeau/g+h8T/cUd/SvP6sr6tans7UgR08iVsws5
kdV3ZgNwOAqhUkbUzE7x/9HJZ4MGDrYBOGt2IUk3QESfMu6h8z2NohcePhJ2tK+g
wHoVHGgvU/+7AvNljYFvTrCnTguyt+SqR5FCApU3qpCshs6wCym58X4OziUQJ91y
4z0WMJ752zqgJX+QQ8880aAgImd3QoQ8/ejQefS7RAA/hZRewhb7B0bpOiO0fpfk
zPjxR9xgWYU4N9Jxb1eWKNAIHh+me2w6x0FPZm6fwQl5U21pYKteahFoAOw//Cg9
1daINOtdRhWcsES3Ut9iNuZLqMQ2s/cqcDoEwuflZuSF8NcrYZc0lf9c16m3DbQR
j7J39V2Cr99GES1K39LVDhZFX0tya+l/GALwnVRNDz2PZisSb9g7vmRJ0nvdNrWx
9suTzgFefxIFKU0HY5AjM0ClqObkgKsAdLksas4vT9ZLRsOdjSgwMENgy1edJKy9
xSdpyZOYaGphLx6ISGEw66yoPkzGZQ9WDjkCjoYITZE976fx8Sc3bn/Fjj7spzlu
94cqvi313jQ7n8asqAavYxj0VLLtI7nII9oznKh4DPK8iQaOZzankxz2IWgfgQTi
LitJvJgJCns6Bk0vVS5+y9z4x3xKbOU4h+MEUW2TMzyUbZkFF2CIWEbQGk1qX9xO
Ksgse3k0XtlKIum1ZEf+1T0QaO8U6Z4o/t1vL5pfT2x5RIHDvBqzSVh4g7+KPrX3
kL9luQnfvWTjtBkyl6k7kdb7C5VBxE4loftmw8mAw33BDTHGpmae/cXPXkYZ/ltd
Bcb/1aBi0AIfkPYYhV+RZi5N0MdkUj1+Nd5BCt6M1EroxLpaG8IAisMGL/U8TA6z
MqRa2C9gTuqJqBwQIEIxAmvLezSA2LrpsRLK0mKpYFKauHI3hmNi1BVkw5wUwDfC
iXupCrApPZML8QbRoiSvT8zRHivx84Krx9P1YNIy5Wv6h8WfzQLBZCJCrs1Ox0Y8
Ikj6tMvdSDN8e7+PpPgP4OqeZWu+ZWVPG2Ve1M/Ji3LCOlDwkIm7lI88PTCbUbOu
jtgT0bgIPJVL68GegO0NWxEUq8HSVz6gEa2YHwFACI6EG7mjWGflL0KNEI8pKBGx
t5jEewLjmxuk6xGvZR2NfwF1cseX3H0CYJYWixMj7xC39yiwTQQ8TuReJ9YftEKV
65ffh0e/jky8SF4kZSSxnWmji9qKS/0vRPmJQ4jkGCxeGfuVYR2gcIefySzyUyuR
WfBY+p6FBXDr8XNA4m0BXsVnBX0uaQmP7Y5jiBROaBihd9jT/nOBOIRwHIDj1L7e
t7r/9Cq7wA3jPShwyngzW7Kb6iN6iTezFV/dqKCJfiPlEGWWrOEUYpuq3uuwea2i
NfzzYM/PwY5Gh/Qn2c/kVDZNU8D8fRYzJBvQlvIe0Bz2kv42qo7B1H1WLws35d9M
D8gczmFvkfgflkwG132m5SQH50Y5mVOkSeK0Yg/Z9IjsO2FMy/YoBnisk306ZCPP
9ktACdp0yv3h34xa0DEoXe8MbgnGTuRglVxRwkr0N4TSN+i6FP42h0Pe+NPXfLJy
Q+m6bFaJrNapFA94T2qyrWWU4+IFgqV87UvrQuyFp5NFoJej8rlqJw591vjMcYGk
RpteMc4VbqIjnAiDFMOnSGt9jCy3n5PJFMX1G+XjtnAU1M+1YUZdShn5jEwqel/3
+kUTqQkaAhe+Xn4RESQEyxfMWq42gyIlhqDdr/+ddiZIFSfb6uhHtz4iyLX2BjFL
pC8y+hz3ASH2jZC0HdRKgCHi/M8niJe0qneDNoGSmbD4FiXEklTpWOVGn8Ts17iJ
PQ+gVgrpPv5QZSEL+8MR8iQJT37frvl1ch4F2YcaMmAtaRrsgCrPb/sBjE/XU2Px
gk1NsCyhErgqsr9AkE0N4plcONEWyvEpBiR/qwPjJ2mG+U5Yto9uo4O7J1kfnGnL
d+QCzN1hHKklK4pAg1tt/5s4SSzD3JVuG8+BEcZA7C5EVMhk3a5rJgA0oyZe0phw
jVfpM3JeP3QiHubX8dKYB2z8fB6dOj/YD57N/hmekTYKNhsC336zEWJYBNnVfYW/
7BoLX9thh2gIginhKLxcAMjmVuoJLILmYwcSKYkQWXyZP+G/kptl/cYoiS+TjonB
nFQzkHhVQrXZ2Ji3/Yyr7HhTngkMR6eX2vcKjDaiudlIsU3M+plPCrobZpLmzcRV
bGPpfWCW+SZJrZKDHdNTMDFlaTY7eXQAxKnDUSynJONQXdiMLc0qnL6PVAgo62XS
dgXbMEN5jYiunRalrQlh7Jv45VE1z+vyTukcY0B5mn9/8k5CMYuuFwH2xFPE4Dxv
X9dkxLyQElgJiyEn68Nh3Ye5LnTMlRDC/1UEnMF72NqEkfmhJCOa4bASYxrKH4mJ
44qrsr7nlJY5Ccm+AT1bZnkVPKuR7tvoGLmDNId8GrHHhs7Qg2PDB/0uXUtWVjBX
Yui8YayJ//WGvMbcwRN3iExuIu38biLz9IarJymqLTxknJhqKePox9mi+v4+qfQA
92kowf9VYpgo7qF3XDCRoGvF+A1HVv6k3SXK9bVWHLPJd/pXKpqk2B1ROU4qkesJ
By1GcgIAio7cvr2rTTt9NpsXI0RBbdz9usJFYpcOZx1g7DKWaaS7ZDQzBatAtJ1M
ZxxcTusG9/RmUCm4NW57tG6TAYoIzEt9gBCeTSJffBAsls7Rk52LRi+q7TFmvUnN
zogNIYid8zdDOFxxTe6v5F5IKkIkRB9ll7o73p5JM2+evP4F8oXHOQDRUmDCv+1u
hHb0bnoX9cicVcMD2VE4Z66SZksvRaCrksI5h7dPEBF0wS3kcRlhG+w3BE1JjLjm
SgVwKBV9iJHLs0CP//1vd+JX+YChrdIjtAl5RAwkn77EHzSsyt1U+W8VCWOCaUOm
Z6wMJaMniVi3mIAhPDa2UpVQ8WkEV1gcknD5uO2Ccmi2MyJhb7mb0mInSgSy92+s
1XASq805xb5VkUjEkGGJ9mjxufyOfxcR5PItGJWtfT1Go94HpaeU0FHZDQK6u2qT
MpEnmFBjaZAVOR5arj7Xn/gOOVhsG58DlyU7BrSc926XXL1qwCaZec0O9ZPZt1c0
bYolqDtwkjjK3CmXyGZkVDwtefBRxmaj1POrzLBQCajxqmRvM7wd+cR9lruLxxP+
nQNTZSXmNn2z5ePaDKZIzFpp8NuC7n4tCfxXGB8S39r5dytxKNf9tWnhNugm/k59
PnQjT47SlGbGEwlGHmf2T9hB5/DNRZlyWYJXw3aM6JCRIdYMWXy91oFn2oHb9Zd3
ZQwSWB1fjOwUSs8YaJDNLkIgpUCqdBRaidMcbbhVQItc7nC+od5H751StCIjn2cS
I8kaJLkjZaEz7CjV1ep+NdFHhNkS1g7sfDBrs/A1bfHTzmgeY0n2lMZ2MQZ+mNIN
sdPlLILucN/Txcllx2lAOS7R94tbrv5GQgT8TSTClrj4pdEIGB1fZ5CGIq3bVINH
qOTOefvMn2P9xXEcUeR23fxpCGxBBrel3wZ2W4AGeZa5SMOthPFiJR0a8U3Qx8jd
d79lmXwXGl7BFl6Y7b5yVq/H3r4YiCKh9jo/39u2iSyLytslH6ZRF1cA3yPp+mi6
cpsbBFNwKZ096xXbL9Ha/qJNZiK4PvpldPrEX4aQ6ZJuDiVRnK50qFxVKK9fXJxb
XE6FEGO3kMJ9GlBGmdcnzgYBFgtabWoiiFhC3JOWZ7Tp98Mk7KEZfXFWPZHZSRho
4jc2eOCooDqvmp6cLxpfFzmVgKqetFCfZsp4VFtOnI3xnn/v97jnqO4lOHbB0/5V
ukfnwzas4zCd7MdUpfeGNRSaegb2wxxX5wWQpOaHFpUkOTjeVXkzPCVIAC0q95EK
2KAil3vRxQCJ7xJb5laHYV4RBoBVXsjr+LOUUlP88x6hz99t2OQevc1wwibhXjk9
cV3H4jGB4u0HDFfKmdmnjYPIghGNSRRVxhvBTX4rMEdPLjitolOx7/sHHrzNhcg2
5iPYeVCopncIpvHU7+CuxkufKbIZlHeK0AuwG/u9PGykeX4fQpc8LJCA/igSROB1
V7ShYiDVwxlU+OiL2wOk9cPDAdSa1gJJ7QUIa+mUeR3DVRXtv59aYobhK4Yr1weo
QWL0vID0sGE9U7/Lx1vO9wvXgBHSvFh9DyZQw8VsBn/3pXGGqHtP+JnJlFAJ4lOM
MTHT7IpmRxdmAArH7oQjuK73dHvqGbkp07KDXdjsk+BufMMTLwpJs9mB9iphVgVB
uUypJK9AWHaBUXArvgr5IzzTkrNwPY6fsjyVn5v5nB9OXu/ymo4llsr9/8+A+EzN
HuypQGl68YwqkmGkwH4DGE5taLdtl7krQZPJ2db+6oDeLfltACuqkAgfTLsCRT47
NtDIqZltSEBYN/WFxC9lh7FV/ipT/aomZrwEDsqG5fjvwcUAjyBP8ZtIY76ON2au
TLKs6NEfifEY4o9SfkqVU0Bn/39bk9bfiS7ltWiXb7Efiizkwv9LsakrXoveniYt
aT0Clrgumaidr+b31VwmZJ7uG+ioJkju1cb6RWSV8vFrJBKHtLby4llsOxeV4tje
2oZfa6d7Y6f44hAXsFBSMDaVe/aiLI3zFpnUEztJD3kuGsnGZRmSpJdfsALMd+eq
12fYvgU+vn+ARj7i+CyP6dYtlX7ok+Kw8brAErhX1XmX81EDAhBSL1hAVyqi64Xl
ihDxxwXMFOn0sBuj/XJ3zb5w7yPGMb49pOhFJSbIZt7dbARUQ8iiu/Hu+8O+xGwh
lKTkjRctoxdE/U8CE7/Diuttb/vRsR+Uj2MMP56vNWi+KutHzzOsuU9+HfOTMZ/H
CcT7708Dcatsjw0DEdBSYUwR7F7aSQDKu1V6m272FSdKBYOCe5nmecrYo5J628BY
jcDbk33aLhh8XR8likVL7kdkXnH2eCU7CwRopbld5dB1HLSp1sByRWGje6pog5Rh
UnWh7Vdrmt/TbvitRnM90qctJZv6oHeDbQvqWG+3hsK21OuPXRUBOOZr+7FDoNlR
i2FJYaJzrgxiqg28vgqE/b6A8B9HvafrXLPH5//Wi8gugG4hRjNrrtyG5iPNPcuf
eY28C8fj9IoBIe4O2NIREgRDF/TD1HZTds5CUQn79UXZu3qlkEgRa38wTf5nrnXB
8A+xABw6RnyzJQU6KiYVAJH815f32JPNHxeZA6jp6g2XUphm3rPaxhodngb7mlNI
qfcAsFRLnuAYXP8UxcvFSZYXIB4qIHF9m5REvA6rWPOKrJAzaIXoxLsEDJo51J13
b5XuQee7DeFtBDTJXA6LVFCFR4LZr3YmfExIm0XMatdiyV3WUIgxW1G5ahapv3M3
YN2BP3BNug11KK2LwHBdhOyPTiPB1qYb7UWZgSkugnjOLEzyBV0+EvqBCOJADUWt
ZracChUsF9qWxkEHJOkMauP44GrdJqMDQMAlRFElQBvVCgeXo6vuqqKMqNcbEWVc
K9bhCMl2PwUPy+vlz6GqT5DzhmxRl6kmu0bHU5AmOPG/8J+DZSj8l7ln+S+xVruz
zIDyDiuPEnEZz3Z6J6Rzf0kzTKkxViv2m9pBlgizGACZqtgL3BSfNE+hMWjUG8UQ
dNI8CWq83xum7BthjEWsYKqtDzAN2rsK3A8wXgMKMyqDvvHV278nAfi0v+XII2nH
ZMzC5RqOfYNtBgxizie9MRnGVwUnM5p2Me91J5GbWaphRGs2OJW046dvsvtFAIyS
UduhTRezNXmopGONM6+fSjvHOhePT7M2gCMaz8yfsMllR1MH46tkhZDdP7a9nuqR
O3WuHKloBxI5kduERUt/LDos2cspKoFD7fF3e90x8L0tS2g/XcUO1tH2QkG/nL6V
D+UhQOuxzDUpg35hV6eGABs0hyJv0KxCV2wr6NGWwDKxAUdFjaSuyYgDzUzRD3Dp
qefdoU9dZQorr1uukWhnIzk7h8VhHapuBI2kw8whvFx2y1ZEwYQDyy39per/De0y
ZJt5oWgit3F1rFU5U2UyV3Ml40VR4YbcMVuB8XXPiTtE2PGyfIL44x3KPOYB30gd
DmlLFo7mFfMnVmcmAQtL3cM3L9fmDYyu5hg7jU+hIegWlyqxvuieWix2MuAjd0sy
6xrvyNpuiv0GVX7X9tGHwCnXCOI3zHdwDZo6HOHBn92tDpLhU9NeohJrPNqGbyR3
VRGSuKHuEIq14b5uqxlTBdhLgfPmHUnIUZccsxQvR9FY5bzPQryaJB5o0NNjn36T
Ye1yMz6D6ydHLRg27f3OlyIYxBTpwaMgDrDjFRtAppzZeLQ1bZAMj5O881WsoNwU
AI0Bcbs6t7xHIHlVKaFNboD7oHGaZgEY/6yyrNvOmeAr7KFG93TsMHaSjjmlIZwL
T5275jUx7Hr15oDj2PZMloJGviLCGxmHCCJ2ZiZDUlcxVMGyQaNm8sNMhL+atE/i
KE8/VkWGw0pN/hzpor1ROUvuPycgcH3azZcgP9zT1o253MJ8qsj9YLO+FoR1OB7Y
EuI0Rn4UUe4MCD4BSE4DoXO5QvAzaFo3Y40rvGbYiezL1bxCIbTY6tEqr91U4SqP
aIw/7HrsZ5FDZ1D6bh5OMiO06weOVYOOvc6VqbvM1UkDvK+P2JxtFIkppK4KGmXL
QQma5S+JXQvOFKGWUqgs79tAFRIGEaNVZjG2k9+24Td+p6qq6zoSebmBAg2VrWJ1
zY/WVtO43m4wuz7VMziqLAnDgcdNiB+JrKEPrRYFJ0q1afPHtoJF1bhfTbwmdZFr
1aNr81JGp7Sukp18SDdyVJcImQQYORpX6CBDdDqxlFJfF03hz3vI5fFMRqhbP/8L
f+Ki6r6ATh/1NHX1ABkgYTjIrf3QWMUP/EApz0aSKJzE26TKw3O1yiWyn7pJNl/I
yjwXG2yewZDL1Men/kbPUy9GQ22yy7eq/mDZf3Q/jhwt3LkXM3UTInZKxr/RsyU9
vB7HwWc+iFULDO6vzLrllIVNyhnNTJP+Dvu1YFzjJNoxPe8x16jzEBpP6xTBF7d/
mbzUv31TALdJTPM3lx4XsaDvEApcWET3p2UT+R2u/UPrDjP3oG9iBWuDZaygyf9a
n4hiFLBxretJitTcjkdWTGWfM+gi/v1uOGvPc7arhkIStmBORls2uXSStox9S3dJ
imP7xvBKc9p57iDT3c8XjcBfT/wgXhFG4Xse9466XkfbKMkecmB0MGBtlAfW4z4Y
tTUNxsuHt4HyqGCq5dDFpoj6EstzWEIzF2vDC3s/w9w+/cyKouUAvSI+46XRgFhf
3Le84nZPzd0+9uBvN6gy4NIxR5B0v6+aCWlz9msYteTD4JgT99UpzL0mBsnrvR3F
LDJ6JPN8dMJX2B609YNyqw5a33eTZH1b5FozSvvLGToyazOM1Q/jDt1yCk8kL/kM
fn/on1GR+LgtmmhCyNAQq64rdLBiM9me4G1ZPCnJZn3EfN/EYWP7bCVFAG3ocpif
buIst5lcLDyo6/NDLFObafQoDfoYZgKkftEHroY6pahtq1MPRdAeAtNsov8DQm84
zX6ShlQRG/SIwVLClvNG8LbJ202V0DIzdzmR+EMLYDcFS4t+xDSawAqtbY6tRflF
+1tZ2GcQ+6YkhADKWzScB2YDPRgS4jyAS/IaBhbo1Ix+hj3wtpsrbwc7DbY97gak
050IJSNKyN/yyJ7B8fu022GuDvTXY2OJQVoInPic4+1TGnVK3rjcgxwTIjgLsGPr
4Zvs2qCyPqdXdRXR9ZdzMZZb9e4Ipv5vRH4OJuxf3Sf6XvNqxiZ+KwEb1jz5470B
xdL+uOBe3z8x0PDm80JYTrHGyo+IMl+9+cLN8zVjYygp+zzC6FggJrsAWhS4Ol2d
bDCpEovo0g8RoLMOTmIks5/09QklblIwQ/zwbsB5+Q1DcYR0vc/ZeXAAP38LUkhV
675/9/gGh1LsmSt/r7QCdrBLQl4LHRbdAX1qbkTlRAhwV5ALTtW2dhocnUYJ7vzr
Hu4Jnc36Xee0tQjTXGpDRjomMo+GIZrjyGQpF6vBNeQHFQFkHyiegpaDBYGSCZu1
HeAm4kb7aRAeAz1V7Ypi2bo7iQ5XHaLnF1EzVCfXrL2emqwnnkqzPlaFglNhgl9K
gRd2zMHtJCrlp4DJ7Qs1pvpXiDTCrxW3i7bF/7/uJ0ShK/FRBHDh+BBBfxmhCQZk
vE5f4RwkEh0hwHBqaEM3yILtMG1d9LMEJKLG76IwOw/h+fVqQcdxPMI3TN8zbrkx
jAx63Lxy29lUiFF9CDPdUaY9B0BJw+SnPKioZQzgW0T4xFEd8JAuYDG5OkTqbhrF
e/P9QoyzvWM5zDVdB31B0B3swwYBMJHbSFd/ep8uojX+quX+0E1SAhVgTo10Rj7X
EBlif+HtHTep6pR+we2cE7JZtkSX+bfZDWg38fzpbo5yvmGwwn0/gEXuvrcZdDx6
pOV3hHLKx5Hbw1msBBT+p+RVO2VU0Y23k6WTE0SSrdhMeZ3m8G1V2GQqRm/gHxUm
eG8pRPBng1nsaSpR+wVMT+jgMqZFj9FjUHqR3t4++hRXF7T85qFlAZdcV5ucVwpt
/M09BZHCHMTsMUK9kE+yspPy6JkyeM+PI/nJCHCJksoAnfRycKPgAF7HqBYdrATM
QEpWKMlzrSijrmVl3RiP8qba6HucU0B2SmO9Pj9ogR/hu1iB7S8px/kJXHaPZXFo
wfiDijoBAtc5TWK2PMYBw3hyNiGL1HdTFeb9pZA+QgM9ndK/kyjSN4kPcq7qKE6P
cXufTCqZkB5z17irKUDH+XVRP+Lo8lxrSGmCS5QM+n/+epN2Olw4PX8DV/G8RES9
Np7E+gFhGdxGPzdFwGf9SewMkgcNRW0ux5N7uktOu79rPKoAt8LLUr0xQXoh8d0L
2130G7E0HEk3zWYU0miCxGqf9ybbD+dPcE95kG99V+jfwz8HRhYJ761yVbri5nGw
H4Nyv7nh4vM7bgBWXU+/f78/kRnPnCECfPZmYk2wkQA3KWGJVdLRPOIV6t4gr/mc
aBcOPslNbkJkr7q8Ar1m197CDNb4tHdVdrMgYsAeaQOalZrLFwXGFS6ro5bf4IAH
1581Q5MPshIy/9hjZY5L//dCWasCr+wfUCYJsr3ElIoZN9g0aKGBTVveZnptxMv6
Cr/jdS9lL4rM3dnN1f2I5iX1fOdaUy17mxewG3TwVRjxIFCCD8t5ahrv287ZYNGw
+u5Be+xFWSb23LZnskahb4g/Fks1mgq4NoACq/t+FtcK0TV6bjDHNtpAIJYsr84p
mvSK9b26ALmL39vAys5uR3Aj+FAl5ywgIKdQHj/V2VNt6yVAH66+ylK76JJYKoB4
iWdipyiCslj58tohRSYRV3Bj1MkYAt4PiNvFRlN16VaM9yijHHracDzfVD027xhl
lymGsB3423m8ixAL3IkjXvzkEdx10mauCtAAtSQxprYXkPdq7dQ29OOIe77YnqMr
w+0ocDzoAae2sNiLRxXPEdsE9fWabfyydTPBZucVslJ9dMSvp3vXQqT9rdrdNv09
Z5lUQahHy8946NOKI/OwICREmk7+xrQMKm95ipK+DDsOwaimwQfBnxDt6WF453KY
ZYsdRNeKVjT2jNQb6jGvpL4uRvCzKjF1CqP0xjggyGCoVgLbHXL0vwfKSxGX5JvQ
+pBCvcJN44qdhS/agMFOz9MoUV8lmzcffgPl89WvFrsEDV5Duv51JolZKhjVmjRY
1kauwFnKjnjO5VjcWHWVurX096NIsUqKdc9DbZzZ3LvHHw0uqzMfkQSuG+9v5xJx
xOOHnDYcx8WX/z/d1uF94fviKYeB/qkDAbEzAwqaTP5HULKZM3PHC35TlGdRZjFY
H9UQRE6GWucf8wM9CBxnaVkTPl9g6KKrGgYPGSUL0zjjTio8VK+/XPe9AkWQmmJS
Xbrt4pNa6Al5ux5J2uKIFGUjKPx31S0mbL0ELoYV0ZuyJ9+91Gy2n7xTxGoPnR5o
0pPM2j7siL5G2kqd1lk6HtO9qUY0mTb0mQsA8lN2a3dDXU0q3XEugSsz3RmY07CP
i07v/+w3FnWmqMoXSM3NA8gtun6aj/OgqhbFo+u1/9X70RH/cfgY3EncR92DptPa
huK7NLqh0oNE90CtLVFmsNQEIBP+AV77+7jnoMv1ZVxkreCeSgQsk1KzomkvI/M9
+0R2ZLHbF3a6F4BHdam8FQH4bsNYT492a1XnZREU3LgpSUzDniZhS53Hx6Ryztxy
axSVfsb/LhZWmApRNEqZUtcy3HuR2k22DqVemDlzvC+YceChjOzqDW5ozFig9b3v
qs6qkRXi2rsvMUY+ASb8iAQvao2/sAr/g7PsIBKXIgQht2rz+3GeYpbJYOehE367
cHDVj09UbwM30BGl6wcct5ssTPIJNsFK99/8Zl48vwcx7vGHwXjmrEed1Ch0afy0
oqxMLJKunx2mLuLReUbgUgJqbDqPSQNf/QjMHBAYIdwsDDWddhfFhCrdJstnDU5C
wBbMKigHX91UFMlYELlRigLc0L5ijPtcHKNAbIJDvPlzOFqsyG8HHtud7UfV0Qmi
NviK616anp84nv9z7mNJI/DmuBVrQ67/Z824I/uQeBFm25ln7RClEhAOYjow31k7
ZuEWduENS/DyznYdhk00VaaA7xoHdEetYzGK5PM953GmF083lib7j7S9aDeAQhvw
/5TnPXSO8BJ+0ynFYrqQ8K800ETN+z05w9HIeCKt8rtn726cz8624VdY+UaAv3PF
Cjeg0/rrvMbz40n6/CpcjLFRMJ6sa1jBQMKoDz+rr3ZwoonnfJ7ggSIGUUpaOypi
wMGHtgHEZhCTDnH7YLVlWA1dD2JaYcjtq+WG7Qg0L+Wz+3u6NOr4DoPL/GfsSe3w
A0kbs0+IO+esGq1ppNdWZFTmbnn84XAZufbgXVjN3iEr9bAE0DqCC83W7rqTqr19
YW9nk/zhdARcEHKTDNfh5QDfclEE+Jk5dS5dlMDJrHR8CTPWd/ClC2EklyM1Zyeh
U853w13tC0L2O+fRZgbQ0ci2m1sG1zpn0EfiyRgKFn/vGandZzOK6Li5g2JT6mxR
7XmP2isWQiqzI6qrZNRjawfDPhMM7akTlNB+lfh78IH9iVtNMkZKYlk0DmWHFsMI
cFvWeDkm6uzfWj74Qbl83SQbrQOjrLceDumsd3PoX7tvpA6AAyoeo1kQOPL5RSM0
vh93fpVAfp6iIzfwRjI1DAlCvP7E3jpk2py4SVMbXqIQmzPlF2TA586AFahgTPHg
hkAQsrgx8BxxyM/ziq/Abx+JcyGkHm/ESdfaHgPYiFqH3Llsor9BB8rnnKoFyAwP
PwpHnS7UQQWmtPVfoLoe4G05xnf2jSx+KJ+lb+6IFIykEeNCLIp0HtEiWKciHKs3
zALLLE7urZPeZ2NJ3iLeVPIVgqejVVuHqQOUtfJMypekE8pU1TlmR8VjAoKiPK8f
n4B3fabKRsfRLM2NQ4AMPRc2oM5hy5apGGWSfIFKYkBpLUA04m4spY31X+8CtDyH
UyURwdy9pPvGASoTQVqUOVp1e5+neBQxeP+jc1lIpYGhp7hq3QaocxQjL7FcenN/
K3j51dGa3J2Kjd40kk/RMoOl4OKO7O24FfC9w/wT2khjYbSV2alZz67ie1dHH1il
sMUgapGymynHix71hYHq/4cRisaKBcSYixLTHa/oOHQ1FaCVaXeg5Nm2M5RFrEVQ
7z636DdIi/tekHqAKaNR429lBdOgyFTalNN3we1TbtcZNaqo66Fl0M+N6RyMPfcV
IlIsFU3dzMbxZyvzatjsnPElmLy73E4cekDyDmpRo8KyXUIJAcBBGDUjnZ46j/L/
wAZk3pzn67ZbKRAjF981vNy/E388CYAmHWiQdcDNdJRz5lvmiIjDdd4nfdHiNvFp
pZWaKRFOPJ2dKt74DeuiChOAxYDXqdXrAEL2ICbuNv5xU1Z/j2vb2Qc2ZDWKBInp
a8PdA8137xkTnyWGl6E1o2DdjxF06hmLDY36uk1gWXLWAMser+FGhTXm4drFRy9F
u0bI9z5tZqfjXM3oagJgjqIWvSkuZidT7IfNVidd4pvuNBFTaVx3JWfBDOf2NoGl
lWxPs3KOj+tRKGMteI3rinbulyInINP0fNcOQpWH5nsOJlaDX/uc+Y2RFxJj8LNx
9ONrNL+KOtUoYyl2UE/rCdak+qlQ//1uhymQvlXRphj1Ozqj1wOY4/fqSTpTDU/x
RC//7e+aYVuNb5vPfZQtZpaW3BwQScfyG3Qy+A0+8OKkjWde1EHJnZ0FhjGOEG4i
ZLAnRU4BiX5LMOWYhTsY5shimAR77KuNDyXevXa4HF1vMD/DNVsAnbpi+b3wps1v
dAZjpQ7UxmDkWQcBPGVcCQiqkdxVeooeJrsrgW4TvbMWWM9qy1XWQ7udFpDCl7Kt
XbBEOMvAxEFwQu/Fs9PUgXKzcPDOllLof63uSE0a4lYz/hjUhd/nQ6KVBTz0F/te
ULyPmk0kpQs1EB1UgjvRxVsQwwZomDSnhlt5P5cytByFCritEM4m61pkyNg+iDp0
8GG3JmNMxtkLbiYvFZGPsipeqW0UhyKNTtle3xlehs/N7S6rLFqmu1dXkp9zW4wE
MSKK3JJyhz8oJSn66V+2UIdx1Id/6ltblnzu5B4VRRrhODnIpXLtUtXGT1o2kX8M
U8JU4XUoWZkIedlBqeDdfdUHEFaXNtApBagMdnZjsQzeIm4jm7XFep6NJhIJyf2V
gut0lfdeKTul4a7ES4kWfF0LpqDqfEJWoDVZGSHTxM7M78OcZD41HdJ24IWuy3hF
MEeKaVUZPPvM41WKZoYTqRvCF9cGGYs5xJH+CqMZSLHCg6tkN60nH6xKxF0Wr+7Q
4TGO7GQJU4DRjwm4zsCsy/eWRTVhZXtTlz6S/VUvDdJmmlQk/AEYwMHADlwMp1GI
dtBFfPSc25iegnrhEvCY5+PRlg6/CzMC21iQQ7g/ifY+7NvmQXhvhAkqd95w3VDH
wMMx2cP6YoA4hvDJgl8qetpoPCm8M+BLTlqanD9fTvGBjCZ5MToNq/j/C93M7/qd
ZbxHUrA/7QG7fzkbKuGDyiULjpZ78ztRM1JwCuEWK0zIW9nBfIA0MuC+jgarjEW+
EV2aiGklgBvmdfv4mkl1FXJvuButFLITX/HHZuP4YyEJjhfmrNQQ1TCTsrK/r5TI
KZ4srt2RMxyhnoWJrp5yUciDhonnvLoUOkA2oDAB3jnX/iQqXhSapvgQkhAMvGZw
rICdQB347PjE5i8lvHEZrIj/Jz81KE3b7uAJ1limKzyCqBLUZkPZpcye3SNaECA9
+97MiLTjgGHLAenHXX9S55gCtxNtjyOK/+13bda8DlshIeMc6Oh2UhOZGJJqJ8hF
2fz3tj2wXqnqzF4GbMM8eJuX5LFwqNyM1R/VYBh9oKpOs68KIXWz8GCVhx5dQ8vM
EsK3w7LXRY6nDaEy56B2co/oF5X7N6fMvk4lEZUFxGPvarohMLvyw7QIj7yeu6Ml
YFbnsvgssX/uHvNg5dbDYMfrrTzWrXVub2Qxh7ILkilUTwVjEsV3CBgAQX2NBnCV
w8YoUDd3bVM5bRe6PQF74U9ghVLrMpyClRVUwrXc5OxzepDwQpQM7ee9embLc5FK
dFquJ7OxRvtrzpGye0tNHgvztJDa3jA8gn4kyibdfoLS9qmVHq3oGTV62uDqWox8
yvIXiI/DSwUN8mzBmLXMVoxJFJNmVPbeipRdOt/hEWCrmvQWqZP42832fUbOg8V2
lqYrHRc650+h1CnYr6y6JlubYSPOc9SVhXUozjOnYcm3DEwRX69QL/CDVENjtz4n
R/TMxrBDO5UW/qe5sVT8QblrxWxR26UxHasRJxqXci3z6pcULhd+zLxgwKuoVJ0n
n9WHDq7+KLZs9CPrxwasdeUKQd6H103ybkVGfGksYlHbk1+gYlqRGdU82NRnegz6
ZZoBM0XQbwPyR5XyAbdsuUNeeufpk4EN3rndt/eoSfmPUly3JzO2qliV+s5+9V0S
5JTlPMSJrrPA2slEIrkAmoGIepA3MKPZ3PAb+ojc38qWRYKGLKMAYqaKu0T7RrQn
anZPq+xIFOW3x1yzbDoPL+BeTLoOxWEV6oKKpU41FPzFiOawtiWU05YBFyoGX8HI
EgOe19NpXFGPGZOlUqg1boMPhP3UZPq+iJlLd7vS2ErofzHFAjKCI26l4mTyrtcc
IMsUmNsogKMtZqVoAlnh1QkkUwTbOqRtUDZ2QQmsuuoWxIghmy219/VnqE4m9sEk
61fglJtbhLwNQM8n2jqIoSR4M93IOhXRAdLWlF5tHEi/1i4k54w4vLol9BO3fZZe
o9pvfQ6Er2ijiRLsw8H/1OvWlESMH7iyhAfzTB8wiywttu0cX6A0sSm4LNbM3Hfo
XSfCKCwfJt/YcDQizjlk21g5p851pzwSJjH0/RGVNWSrnq7dCZVZVnCGCWpzmv0H
SNplvi0AXw0wHkiAXJEK4SN5Ezz9X3FG1/lf+q/hRSnk1CC6C/kryJTreMQiWhgt
5D88cdUgPrgEeVJC7BZT1vXPDHfCerdWQfQ0Tk4sxRFsYL0NMuP3s8wCkAcBngSe
I6H223jIzgfc+s2WX2d3y6WpI9GeMWi+0RYs3uG59LYR3AcEV8vzVK7HNVWQLOF0
LF9iaEj1ESPkyR/u4czISHSeLljXwsf4REvgQ550nenHcKJ9mnnzsFHbFOChiUdB
qzVmq4sQxD8gMMR09hwKB9tvqGDWTeawDCT2F7wxEx6OrT29eP5d4pRRgD6fWdaE
p7Tr3hEe/a8c24mTAv9mte/oB2wD+oJzIvYWubVyY2LlRAOSLQs8iDIoiL4/nGUU
WzrPqHI7cZLjY2ISIGhr2+rrJRjdglbZmCtG/aehCnp1deUhKOadeoZBQmn09o/f
ExnmGlNiFKh/uEbUpmLyXXbJvSp0/4uaxGTHDEGg63aliceQjFyk5jdpbM7g8fq7
B6zyK7SVx8yn4ypkKrrS1HwEAGnvz0sRGSvkgxiK3OI+lbeupWOMfix24VX3R1CA
sToj1zHs3a4rye590BtDmjkCGbV1RUKhzT4bVCDyfkk/DkpiDhQafZQ8SROiQhIa
1jJf2F0FMozFekmjPPFIQNPsQJMyO/kp3NhzdtvwfjcAIcJ8pyfJkLqd4prtw+NT
LmWAs6+Z4sxuKAPC1Yy6PNh6imcTgl135rlMD7Eja2+2OmLNhHnzNTs+yZAuiu3s
EHoCyW4qao+94w9kJzU3Ah5UysoshDrm/0IvV2e4up1OTWqwlQ5+ZlDkKTfenwOG
+dzEJPfIRp/xQp4klXYTAraHDHOnEmXv+qveeCaZZXcYt4uAx1O8yFsvfMZ1DLmJ
O8cL35Ytaeuu0YiiHafRl0tQW4VUnEDLnlQOse3ZpilUH9PlmvKZONbQJwHdxVMp
+gy+1E973xNF5NRyGIsiXrFsH3pnuEjifAbWSjxSFr+B8b0N76XkAM/czV6BdAq2
Cn3EJ91PO2k30Amdtcn77YVmODHNX3bikQtNuNPfs3XpPLIIwpS1Apm0DutCcCh1
K67b7g4IJqP4x0XqEqikBClLt0A85zzMWxlxuHKeSO8DnIan1Ui3zJwVmK0TqwEX
nkzrOgiiNW/VFm9z8ePfWK6uGn+yh0Q6atOiR02R0Hw5l8uM92Phdc/KJXLON1mG
ENUFfXTScmCLBV7Yo2l3zvyQ+z/RcWkkfWOW5DUktGAskon8a2xNrfe1V78GW2Ey
xXaZOCh5Fs9i/3GrA9otvPNCPZeS6cjfbOsoM4v1vo10AVlQxeAE1uVUG1rn2Wux
YyJDK3QQ7bpDDH1JTUOlY3OxDJ858bPEVJMdDUtcWC6DbAr7Mr1L5GXztUEI2/sf
5rCdoub3LfDoyOeJKFu4acMfnu41kLEWdu7fLUxpEOqEg2ue8svby3Zsp5JaIABB
KIqctaOK8cFie4/kV8AyTwrHkCu/XTug6WKG9YUBi4SPd3piNgqPX2vDScrY8zwd
keCC9pCRtQHKVzCqPx7HxdvldvpdpmLb+OQ24hpNQrnx7t7yFcFh0q2XzdK+H2Gh
iJSi82cSdwTXmZFbDD5CkPVMY/wVKWRW9qqlsBXEuMW8FaSg2f+UKDZE5YM8Gfac
kpNGXtYwSPWMmNCW1QhbVINd9/LtYTmJg3TdFrFOQs/VSA1iyNPeqlzAcl5N9Bpd
RYMxYSDwq+ZDGnan7OSL1wAKjHW+SUNqZPuqVwbUlMxBxdFNMgvGGXIiuDMIfmhb
PARWTuHE9k95KjcCwUMVphk1fJKlLPHdrvt6mgs3irxELyV/gX3VIe9+PuKGnBu8
YHO7qUd1rdE3YITtU/mH+vVGUFI+rVpNPAAzxDv19+WBOYDUyjwW+rPIPuLcAzC8
UwfZgF0aEIqok1lfr4NEPEIDwqs2u+WLAJ7bhEu1BRyZFueeZB2I4j/oOD4Lsnk2
94gtypeAYhFgC7W+/8YpENIcs3RxIDA7dlCuMhFK+lvfCvGfW/mlYWkcRR33B49C
ZQCHLwwME892PuhAYZwExnWmgzbeAV1eB/3AfggEX6EDHsUw0fa8Faz62ZRS3biJ
NjS4mSkVohCQnovy/QgsA5BGsFn0/xWMA8PYV8wCDp4IMBKdxPse1AP7LHbR5Qmd
0zdNORsoH98qX/OZBR4sX+YqmIfU5/ihSEeCRMJf7MtYdmlqlHrUDPbbnpJE7PW3
FYG5oS9Avwfk70Ps4Y27Pmw1ihpMvybx8PA8gy4uddGtEaBkXLCaLKxVDg6lxBYu
cw8OTZmvCQI8eXPM++BRyqmyldoTmvL1LIbHIElnH5ZbWXkZv1I7fVAqB6d17ZXl
4COaTnfZZUT7Hs19QgPvKDP2ebsq5W4F+pzJmi0rm4mWGqOWxoFwktxcaDG1vXBd
LL+4wzXPl6/9k/zHexswIvFQ9fRIjCCb320cGwqbwicztGT3my2mVtmx+7uXUREH
ZfAFcNKi+4f5fwuVyAraVbOi982ftA3xADCbQJCzS/xOjLmfgR33aqxKa0EC5N3r
ZsnXVtyyZP9F8WcMtdxPDK1/ApbVt/rLD7fX6BY+90em3+83pFVsQIs4ASh8WGBF
O/ZKmek4FGL0OQrBmPC5AYyOorIaLt5iHnBl0kf7KOX4c2ZwNWSSOdKCIwkI4dGh
4vC/fGNhcM5sdE/97lsCsfIGDYSd23zjyABguLvMEVNRsbC/MwVLL7Kx4pg4/8++
96I3eysjiDug1sP+PVlKaM781ZNHLgzubSycqPjGDH+L+tgr2sJ0qD+96MUYaOmj
EB/IyWQAbRFHtus7ZflrjO68VFsLcrpt5Xt5fLz6KUdUTjecVDVrodbaquVc5ntO
2oIfpRiQSAS93iqJ3oa0omHXxbIQFgYflY79/RmKnwDbx8zaq/uv3kE5Ierc06DX
eScOGvec+KsOHv04X10EahExmzy4UyP3xyY0z6U1fraWL7Ae9aFEjMV+MR639UlM
SVC0aGil7QMVuAAOsiIcGMKfGBllUKzQIAN4KmruycbNMwhOHnMWGtYLs44weZkf
TNZo4yE6E8Ap1y08/y+FbSaYEvAy8wYddAkxW6XePvyrhA1qLBQrHSZhEBvfY4Vn
JmEMzK4P2qSjSxjnshtu8J+33KQPdeybESBNpV52EEODsYBhRVGtrs0RzWYxGnHO
HNgsGBUgyN5pUx/QmVQgPG4mgLJsghYYNKxVsD2kUN90iGYIIdkfMT0a3CnXss9M
x6MPxm9zuLaIXIJCwsdKntpgkPsSNSkxRnLxob2F/CLePOS0c/EAUZH5+wiJFnDr
gsLcsZ+VM7zgi6S6fSM4ChOSHTaAWNkdxjqhEkBDP/H671A5ktacRlENKrOWeEyk
n561JxwPSSB1/0iQveE96M4aCRWaATuq4+wXfQtfBM+JzsfQSZx9kkRKQGCcIHVL
W2lXVAsGVBVxZRrYehUGScFWHolo6qNWrIjjmniLh0bJw/4RHidsGim0F7HeOHc0
wA19LZ41xmC0rH4ao1+RkbMO2PYTPFZ8WnZyWFsQSlE9Ec33p0rPsjHZXGZvcIrN
KBzcOdXUk7BayKqXrpDDHOio2fafAH8XPO+A6l6CLC4X8WlkkPwmJ/S4wBQ/SybU
j4kJol34tzmgKDTK8jSema8JlyG/6qFm5L8Vy3tg1hjyJducUpon7l5FvHWR8MdQ
bxCdASVM6+eDpXlJbfDoMz680vZtiJCl9o7sX54KlqFPk41pqKkSSwHIsFpJ2AAD
KH8EWNQcj77ixqe7dc5KEjcAAeDk0Iyj1zcPUgytvHzvjFqE3NFugPNX+e00xL0w
tiFBUN6OGn2X14grZPD1NdlBgXmmIHWKajETpJXS4mitE3sBK2dUn2U+rjOdqnR3
CjmZmNBH1/R1sg4BBb3c1AfY8ui3h7Q61jrFjBRU10AUhyFX2/CX75aLKZVEjX/G
QfxWa6rpo7C+YttM6/40HE146tQq1uRG5QfdYzHGGEiPyrX6iOAaCNX6NxLky50X
UvEWYXstbMKf7ChlF9/R7A0XtOXT6dZLJV+NjLURBhvxkmLqoi9bezvLtkfRwB3u
GT4vg2V/OwBHCEIxCvGaC6XBmf4FDZF0m0P6/8arLAmGXwaJWS7Fm2HUHspTsVlu
VTQfuqQz6+if/Unia4GjJyV5cJEkvZSWK4hsBI7I72o9sa2N96Hav5SbzHYdq5Lz
lgrrhW0lCuW4kQeZzV+6KIIT41k6++iKabZTePTwzs+MUZ6oyvNdQn1jOl/Iak/A
drj1XwMchFNIXBuQbjhSHacVXd1Cupm4gB3ed3g2NqtAcsH9el/CrTHcNnqHJ5iO
7x4qRnZ+GaBn6Y72x9SHBWyqQMKui13bigKgeZ6WSLlkNiVc2y+LUuwtaoiLSTM6
qv6do/mTlbn6lZIlSbhBAZC2lhNjvdqXhc/KyaFGFFlALPCwXyB0gq8vIQUxa+kq
ImKOBhURxtesuY4A8VnwiYwVSHXCpvrvNyTEANiDTZwRtmrLYdCK2FX3dMOQXbtM
VeippREx070Y+XFub6QFZHDczf8+roWtVO+t27J5opqyWQh2p2AzUs4l4D4J2x6R
fAbIj37bevrkNyAsf2Usgg7bFHw1PgBFoY7I6Y0YzS5ax+0RueIEEc0lIYlVuWfb
g3zj/3MpIiLJs2BvvsiBpMl2LDXzHe8TbQUsFHPbu5KtLhSzS0T+ZedDk0K64R3Y
RPwQGX8K7nx0XgDgoFkOBz4t0ucBr0q/NqryqSAfzG6+kYgwJpgoLIuNtrhblpHO
CF7yMkqHYR+ui0Vq+kiFIJOrN1qJVdYvG+7plb9uVaH2jPR3yDnfKSF+i8RNF5mh
R3shXsnYVc/sOC6DoOESNaMxyrgZ6zvIKAnidJnZrQEirtEAwwS7S0Bc+TZvyzIz
X38aY1xMRfk9rcuckYRaeaduih9APHUx4uWZOzQ2ENLTsods5PNfaZy0JoC2OEkl
R2vNTA/09HdWAUnNixJUeLo6Y6QKiIFyADDrBV/65coecfXuKs9IjUzve0KHJEia
wReG+wppefxoJI6WGzRz6X2s/ggFSVjASrdy9dxIMvxxwqnBJsJyO4Bai5xIpthE
QuahRpJDKRI2iYHbJcwny/qBjbLHAQD/kmjAwj+makTK1quDR4MmgYYw/oAnLskc
RtnLvl4CRVDCs35MpDBC5xtBoDnmwxJ2TzlsM3HoXkKeaGnEy3/RfnDYMQDnRW6B
h5KdS4v/ZwpQnq2wT6INRUGfDHk1Fs3vkrYwthGXnUuOuoaYNw/SJpam7J+epj1n
k9x0t59dHlU293Bff5kUEYs9Fdq67ZIJoenjyXv9yx4HgKkxr+UY2u5o3a5CLsfN
jZYd/nEOI8LGcmimxrLL++emZT6H/kqbWfC242ONT7O4paTIParyRpGsBYhSI2rD
O0a/+vziK4LE7ypvFWc2r+Z9Ryo4FR4qUeOgd8TjYqxAYgm4jFWKNSFnYpeSp+OB
yaOu1D9k7o7HSD16u0/TeyM+lfo+5xH2Ut5VQt8zuhe78JZ5Hf6BbVdZw37aYLZj
M+PqK+M0Aj8gGdEh4d0FlSOh2YkLaPNCPiCFDcYcwqFWNOLhkyy1k8hfbVS0KNRJ
iulpJ/5eZkKBGxgbOmzhNGKgjtF8uxJBdDwlkWRyH6PAX5wtVe+izMBDVls3xCyb
YlytgV+yEpIazLLgguNXt7irZgtVgot9eYXFGkdFbxhvX3S6sS/OMXOr1u/ad3cf
gJWhHPvTjzX9Gdj37JvulgaPp1oDEicN1aTq+hULbUCE7R5i/FqSC+TOnnRMdSbF
Em/bDpg2HRV17wBjSgeljp+FLCcDHgAaaX4wCqYf96LZrSf34W8d+ttexHIdi7RR
dwvn5HtsepXvfpwQMduwpqIFcJLZdh5NpyGzyeHKI36JhJjm/hm9rSrh5cX+gkzn
u1zNPqYtyC0s511RRNjdc32J9OwIC91JSoZeikPk1HWolchuyIzGYmoZBBTpc3JS
rvdu7GeSYdW6OLncjkpNF6kLcD7ZxauwedAqN61PQMTljavh7BfWpHrN9duNJG8W
9tRP1cpAjvH8pne3lcB5a8hfPPpuFZJiipoI/Be0TGAvfin0x+ZlP0kjsLaU+oFe
6ORAt10fY2b6NfR7GUVs4eQi/4WU4H2LSTMxE5c83iO9kbzsDsXo/7rdOXWOsTaN
/Y6tOUU2c+5wf0QUwge4FhCcijbAQxaLmS12v0ohylfW4f2J8rbiK5ptUt3PgrHz
tL+9kmL/G88G/8mFMIVF3c6QzII/BDKiSQc7tI6MNoxsOHu3o7ZuizQQhsHc4jaZ
wcZdwN9EtAsou461Rs9b6bXZ5IDoTebTTZ4rr8UmBuhIarY/imflWHoZiZ8YDmYb
nFzoBz21IjIgbsszCc23qXGvtWzMcjwDcuPGifba8qpR6Yjn7Y7vNdZeX5KfGhy2
NsG8bhAu6QU58qoqKuNaIOEMxZ5kl7asI4tA/7oPf2KgveNs2FIEsKueC0tHpc5t
vsPX/5nXYjbBfifE+hXFiwFYYWcYuHpXyPKvBuQIOPU6NxaMmqLhOHzDs70XaHnW
jrmCv0GF80MhIxKYjLgihKvAtSOrMiAuWenPlpENA/QkStny2vYA4u3heSccNckA
l020t38ebZ2PN3G1umcIV6Hndrrmmj7NExBjXc4OtcltrCogwgGK6eibh9NuiWEt
OG1cqTTRaGqIfR1hTYmHG5fDaITIVVi06qwnuvJWxvNy2ObUVT5ZUj2RbWzO5TAP
jZhUeOiz162iIZCqJGN9Plr9tuGjSE7LMiK60ynxlNvXGZxrdw7nzTm05uhlFSq+
yPggMtOk1NeXBSh6F/MqojU+AHpweQHV+wrk1Pd4xB5CRnmKc9+M9GMB1h/GUqrU
NZKSECccG4h/kZzIv6TAtvivu/N5KhVHlEtJYQqz6CPn82HZBZ8+ONs+HFWcpy+5
8eG1gTyu9Bt+AZ/wc5BzVyoYQMGCy3Lu+4bv4cZtOpPheHbU5b81Tovxy7n5Qqzw
LKCcXShJH/jzHmmeuldQNKCDc52EaWLzy0Bva0x14UxBVHklSglZG7zWdGqDfRYe
sjZP7iDdDb9sHv6fbQCzd1V5yi5i+yCMVjppzJPLE1amNfZ6gwHAqiZNBg99vOdp
QtTauoP3D62R/sFKJUvxADJUXTuULeZMX9hZc4qLyc3HTkTBOqUFq5+2NJlT9tnC
TNgxbbcmmK+/ZzyjvFsdM5FVOMYNNdUMd+NHCHzUy0aF3D5F0V/+ybQYa7W9uMq2
5JZbJQDFk0CMkQU3/AbtFipCmdgU+NjedR9tyRcvnjtYa/IVuqX6wD5guqqOHQbC
nk4+GBej89eE6TGSdcwbdIespsklSknuKCwVkuF0NdK6tedY2IAVdTLwtWbShaq9
KI9B6NHbDHV8UTrmfxikOPJS5F+QcotD/sMHTuFV1JAa4FCaEqqiCh2bB0xEX/jf
VSXRE5tZdcmLnPWV2Hxw2lDrX36hyg+Q0bIxvUezf2RtqlWQWyU/cC22QAHnnGb+
g/D8TEQCYuLyZfm17NUwOLnlkgRmfyZ67EIVsFChyDua+PgvX9JskGMLdtDkQfhJ
Ytphj1zi/NNCM4aoTm+ei+b5wN2rYi56jwo5BZ7hBnbMhoJkZl4sI9m0bH72VjV9
RKWkGZUzJAMkqp+UDsB5S7iGrMkvqO/c9tRD0mHdsm+dKpqbELL1eXf5ofg67FGo
8esK/8zwo7x+ThgHzeISHzwo5Jc430kF/8HNRX+XXnzPc5K3EVJdgqahdXSZtvbz
m1c+38pz4Cz5ITRTHHttd3Omo6DbG7pbuGAyJ4mrZ8kw82btYiyxFdh36DTwAqcR
uaA1VAyPyb2EYd8a94MYxMaXL1znsgLRzaJfSRL7m4/y8XfDOCWo8zykK5hQeLvS
vtfS+3YrOLncKRFV4e+/xfYuv12KTaGv0QI7bs2ihgj6rBMLjoz1HI0YAQ+4a7I3
Pn1nBzNbVeP40093bxsSQ24x6Ac+pa+Gg3LUMPZaYOfT9t7Cf4umeOki/nCSThLR
dQt5mY7O9wfVLKm++HgLCMuXYmEBGZ0hrnetbOWZeffEYNClQXM09G/Ltt9kF5/m
iY6F6y4tJOZ7KPENEYiugFCt/Fjjeix4eYHJ/n4gXqQuKPKtzBnbr/O06UMMnNsm
rqu6qj0/+cjskGoKEOYNirc4LmMIviO6Oakqx9cVbJsI+GB4dZ2JB0+zPRki6H1A
siRzgORntNGJkQOuhVOXX8KLFNnoCP1wCfwhsERQUCiG1VvOM2CEtGVH7RsPRMnY
Fk3vvWK7DTGqm44cfuWKOAfF/ATCr3X2T2xP80gyAtYiV182kaCIeF6wrR9LXBfB
Pw0bbcx6joMigdli0MsQX9OsPkmRyQEGTkP4XSl2KkVsljIqCUb8b9x9MJ5UHvyw
u4LPsGmB/wLpg8Y0ki6RitJOar5f2TlkY9JH8vX2JAb5hvQ7pBoz30y0gaLIUiy0
hBvv+e4RrW/5GCpkBi7PrRHImwdSI5w/p0gnP6lygOGfv7O4ZhmiLYPh9Yv1wOzA
OmbmYXO0N+wF/TSEPqZLatwX70T1hAwLHQOLyHxD8rTJuI0fijxw+pdLBr+VIC3B
1ByN9toSMqxfa7ajFvNqOVS94STCziRVJODCCLf2mfpS2S9EpVQ77t6tJO1o0Nls
cUxQoCWjUUz3dvTVq7WPQCzrMXc5ajUtaJIk3sM6Tt0AvPfTiaUf7ujcyiYSNnmc
Jec+6RtcbXy7t5Y1Ws09WCWqiW+Iul8OvKLfbBI8Y8MNBgEeSYqm79eQG4z/bL5c
B5rFFKWKMpcYydvSAk2eSs8wZRbRl3ozotmXLx6EkaMMjGLWC5aaTliwHmYKEL4V
TzslABSyW6TrxVY9GzZuP4j/u+MLUaCAUUwoINKM6HU0o5ucxJQNS5payfuIKavY
N/frB+jXN3RIojPNGj7R12lwzSEYwqInqmrUFerNvIUaFGbgEcuudE1ZEnmtCjJb
sMDzMxRqwHsIS2DG89iTnbp6sVUEvbua4RfTmi1Ulrj2Q3qexpdIFxUYBZMlOf7T
k0GfPx3MZOyKpPO/L8LbeTqaShtjA9MTAjIsvlR0xY2BoreOra5T0HcP6DgVegj5
t6FjuB83JBe5uIUUJH0MoGImmz4LhG02hi0J63zUgAcyoeW8U8KHF+XLxsfvjI13
sopVpgeOOfEF7exVgWi59BpU8plh59q7U6XnPUsK90e+6yYSTbmTf9Xwptk5wzdb
o9CX2/JHTLxJ9FpAzSkid89xpq7ZgQgdDR+rJoDjqmI85eM0EMIEQbnKAgZu0e+M
2Xv7J6g6nkbrdW2POAsS/8qG/JWPfnyMpaWaXsVQ1brpidi3tcHZXKtfXKGLMnMl
YLC6rWiYHYbSOkzWLrGaSjX5myqvUwzaEqjdRrGRv3vsZuYcpwSK26LPXPl6E/li
VJVjaPNkUk5rU+jEWdmpzoSC2C09y1p3vjUEHUqDmQCWbXpFc4Ecy43kHlRqgJb/
72xs68x6eo83UHroGmep+szqWT08/qu0XRyvmlZ0l2NHmo2/yEo8cklWNYoXAAEw
RIkTMYzS4v0grqG42z0k05mVyP1ud+GNan7ZHUNOsNzRYfYU3QXuh4XNJ5MKkPk3
wD9vqLQxuhIoNGkIT7Wcf2VAEJOnFv9p9j/Nq+ifcMgew6FAqOPSn1jZ15JYwFQW
OKHUqlLeA4aPPewVBcPnaoOxDhVnf3VrXV3CXniQsegug7w0sKpeuXzBPPJSQeMB
wmMh4T46OSf9lsTSCCzVcKBHab/RoRat0zngPPaw6SE8zzspHitDFUhh5KsCJGLI
gTPURoryKGtXh/0FVGt246akVyBXuyfspyqphDcC9nzYACpz0s43YVM/8m7wKqPC
ZUbNxcOJOBatfX4uiI2bHmTdwzznaPaxkeYV9n15+0HeQ9F87xd8Qbx3DBPBNXvH
fdSFPQ419kL/uFoqW2OJWnlKSzoA6dm4978t755VB9MSssWsqkkuofaXy9Dt/3A7
Asn+GsarMLtztJ77ijUTWW6mzBMIs1YmbgP4EKIRMJv7isubUrsps2SNVZOjABaI
EOnpvirtBnUCMRKv0uPq/XikPK1N1c+loMg9tLQnmHtnGxxEpbeRvc9TYaLB7x9+
BmsK14ofXQLvcxYszvDZ5VszUhoyYiVSfYAeOYDdhOEAIZsT5+CfazkI3j1NEajW
nEYL2zcKxeQjww6vRkPqeyAJpIX19MPGB5K1Y6JXSxF+CIZL1SelQEekfsycPe1t
rH5TEctExEM2gDztR4k+sIKdQ5NpHnn+HTGQr8Tyrx3fgsPtFbOQlSfnsaTraK9t
f4V3SA3tK6IeOHgNtYDIHl/NqOsEjY6XJqE0Cd1Xp8TLvNEwFN+CNDZg8NvIonLU
qiDkNw6lS13NShN6JLgxespUjnG59pYjgNzd4u2qWKFNYX5B6H2Y30LJtQTE+5Yx
8d1ODHIrKteKShnxIF7Gru34yQ1QvxH5k9IOl0UALJOT0/WvIsOvVP3MilaZO2VD
/a2dmqdbVlHL0JJPiB2vr1aJqjkAAr/VZzc35569w6iv8Eljo7Xk9o92g/t3jIWZ
jxYll84tIlaMDMyE7fEcwWovfyr9FQQ4mOfCv/zGjo0aHbeluTmdDqgDDu+9TSlg
Q2ZR9N/sMJdHyH2DAqaXe+ahei1MRczRhdlIx18j3c9EuBP9uIz4w3BqBRsK3A3n
jqkoE5lVEglDpVjaOV1IyvqWaGd7RNdyzsaly60+N4oVR+mBfdXi1thB+Bkl+b42
J1QaraVRkGjrnPeyz9sDKVVbywuGvQ9IIL/RvnN4bEHpsEFoQV9GUJ6x9GwXrOck
fiK7Da2CDXwWA7PrPoCPgOGIfFOh9vRaJpnMp2aUP1kPGi5vtCCNQfeoAeXx/U47
+hIDlVEPYc8jevTMGpkcMUduDvhJcINwnhcEowmNwXECxUgtg0YdqOHKzoiUhxvc
Jc3EzU0F0CRQqbss5g5YnIVrRKKMet76Ds8b7zsW7js54uHF8cMlA/r4vvc/UGu8
LQxkHmj2ynZveMnegGTE9VdeZAN69RDVkXA3OLor6YZNfPO/nf1omAd+QAwQNzia
gqtKP0lJy+Or7uHGx/XZGkaTbaIOeryReH5wj8K82d38iL8hg7i8/2blZKpBccrF
7eOt3X3BI+gYy3wrOdvr7oK/94/By3bK1IHlMbXrK2bj7HPj6Q/YPZAS2TB7qVwo
SCNpjRx4NShFf1bAapjkuTd7kel9KsAj6yLuz1joDEocuirEI6m3RkbpO7uLwZZP
HtbhIFlAbardFWMLGEtkddA0AzsEPpfWsD6fUC04yLzhB057O0r5MKA3Fq9phaZX
P6VJIRO729swqnDfyBl634qnPw3Cto6H38POfGg/Or3cg93zaKqA9DCSusxAI0Ga
tUDYeP2BDHELJBQgd2hXWF4IlnbK6v3aNdwBgA3nu9Fspc9QouAVxkLURyiZRcJv
OZJFFviM/FBq/+oVKllZof9OhFCo5bb/S1u2jJlz6g18QzwPgfaD1dkSFh5Hvt2I
4ClRbi688H42EgrhpGVXuPtMucugI7BUZi4/p8Y8WfhwcFTTscRw901nNZ5j39Sd
MaxNn+rl7w4nWjZnobFh3CGhwNrqGhz5jQDFfesRdAiZ7cNzArNu6ynCUc4daYrn
EhJ5y82BN90NvDBac1J8la3cif2p9ORTEvMgwfAMlqLV8L9rp8QZm8jRN720aRMl
Q7wLFBCUbB46gT50fHWiljLHsSseP7TQdQLrZzKlPYD6RZh0vU4klrx1o83Fkvi5
YEyW7B4ZO3wvUFWIimlZMulK5I7R4uc/+7zPymzdj2YBX7NV8OEUl1jFFQEZzzCt
kR62LIi6FstqaeOLw+M2I9NeuPtIrEeiiC9QfbCIvf/8l8VnMImWoR7RJOodbNaw
WiXRomfjca0P5n2di7xezGa0jQTG72V4GAydV7TM0Nk7rzj0Ursz86YU7k6zqEq8
n2MwaocGYzJFWAPfde3uPJWk1vsvuw6N1DkVMkK6VIDVF6JgXooExTPlKlgbzbb3
TwrEK1vJyODK8Pf9iPNzOVLpDr0qdB9aMhkAkVkQ76rWFrsbvC2k1SHV6ch/1YA0
X/hoTaXuAY/pPQtNWXT3AwmfnlsLZeoaS2WDOevHYniBTcm+rXto6VfagtAzkgUb
lV1mDGaLDgmj+4y+fbtEuqZe16DIpN/rIqZV0ZEj/ketxNtmgWknO87Egqpn4433
y3ZsAtCyXRYK3BY+HkF9XubxLgua3efKbH2i861zCEOn+QT30qUoHvGyhLDSoGiq
2inzSfFXGlPYy4AHXcPOeP/NMRbMbkukech8zvDyBi133DkDgcK5lTbiTN58Sr1h
GU7h/5ikQNtkh8DAu/vLNE6NF30qeVzqpKBnO49EbNRdCpFXt+LLys9R7hHvtOQB
N6cWqCV7oJx0pPxINg/+MuaAip+1tFp44gpUwmB2qJ4PTeqWzUYZwqL9ute/q+K9
na7tvW4dNF2zFt7kWqiDmfHw3OQ+TdoZjqP+CFpjjYByWmNdOUofV2K9eGkT+2Ko
BKg2pgn8hFhyek+W4kqiUPHz98fZwDefKzuIaTs7tXsIksmSeWoRdzGSPiD1m0kz
OVl/hWhiOVlasufyzrlJD0UP/Cx/UmlhzaHo2mpBqKq51SOHFxRUgdWXVhnpQsmZ
7VW8A/p8f3yk5teDpstiGSz8XvKgT5RqZxzJPznlhIKm7iNkpe900Ibn7hiCX0Tm
5txJ2QEDBt+1DcV3jlEqqoKwtcbM3AW5bdmxptPKODgFe7Bhytl2TRRmTRL3oXsT
o+QQ7Hk7vN2Bl+7jgT6rRykrDcSIenPR6e5NCLVIZq5tQv/szQ55S5YOTyPDm9wb
4KLpKdjjpo0JYDhrzuDRo1pBbh10QIrFb8vTS2k4Ur0jrur+/XdA4IHPgY+SjPTH
dt0FDN1kZHdm0hd489OgTB2w52eiqs6nJ0VS63MBcI/KkOeWi1CFJb6HjUWXr/TZ
GTOMmem7aBMdGkmRBrXMsUiQFn99egcicH6oILTen41ismVyQ25kmKZ/awS7rSQE
Sg+bHvtqAYqOZ2NbW3WZKlpHhmhHtwV998ohHYcqCljfvGM+0hGwVX80KpljEw+9
tx5JhEXXtJuMShyhlc3OW9xwy/fPOLALn2VEdy/uj6d4gsfbd6aB7dK4KAjTSQ2R
oi09CNbz0G7EV3vwWEmdEn5hNHxTeGB9SNVpK2mijLsyk/XBVMz3sofoMdKRH2rg
/EgY7QXEQsGh/sAqgL8nxZA7rIFGnSUgWLxCuOWKao48KzpXlTR0+4Ak0zRJ2W/f
FZmnknS00Z1eaZrIoiVeODr94kdfLQf+BZPTUe7PbKWygqqIcws+FwhgUpLFDe6T
fZLiTkZNpTI6vcnKjNSlgvE/05iDW9jsU9zQenk+2efitDHZeCqX7Ec9iu8tGqYX
0kBmRKl2O+WyH3hSeE6i9Kq1XWULx4JJ5PXvELzMIoNrbGEIox9mlEW9d4DdodA2
kNemWNinfUoC/xa2+kE2Wh3oFI0WK6vKb/5dcEGzJypSy+9DVT1ZtTbOOg49ISZB
C5sBVPRlQGaeqhw6Zw/gfBLpAk5GqT/PAVh0cU3NJWaC7RfVc7KzDmjGBQMi1+T+
LydD1gDEpqM3ChtbSG8c5XqcgeiLSpuLiVlFxSeAbgjysHWGRB3dbnwSd1zSekkU
vGHyqL3afWRwh65TEa2XQ4wOv8a+KkEwgYaTMGF6DvXeAPQ3xqwFJll0BpCaA9aI
LGBxMAmsXqICRTPsESJAUtD6Ml+opaPDURzPJ0av9kxmQO6klTIBxW63PH67xbTf
rsPaGqpDFUO4odDuKeGWnctUYVFqdDsY4tFa33P+2RqrZPfcXLQv9O5o/naEu6np
WlShdngbr8bYrxEXDVAeGRCsBewB4OCf648DrxMPPp4rzGvBCz1m1nmR9N3HDPdU
VIelrNmIDxnbTLMcpyWgTxVRBy/5ZdnS6bUWcKZD7pmI5nD0IdSvvK3/r5hH2yaQ
bgNpzeOYp7cUf38dm8huK65V7kssxpM7/W9nxAe5wAA2wEkJr7Q9olasRICUV9x6
Vs1oO5tgOGAQbIPK6BOzmS35gZ5UK61QqJ7+0IcXsK0n780o4uMw7biGo05LskfE
J1cFX7qMiHzZdWgYHskjl77J3OP5zlCJb4nO6pqe1kTM/3SXoYCAnfWX8m3iJBpw
qoxV7C78bGyWaIcgPi2BjfuKzhLBcRD18mwGUHBzMudB61cWSjMMUnVUOfFX3/sH
X0Uiv2O0sNUBUwRM0Xo6Tjoree6W9id1TdrbQx/+AWjGieSLvvZeim1DXa05kBlO
fPRCDJR71ppbT0grAf5ZxQk0VfYRa4lMWPEMW641rJSbk6CpCLPs0zvdfVbuD3+/
imXT9otm8tvgzRZ5fDKBjrGiTXe53K7xCIELp9xsQUXmnHXdBsq5Tg6b1RrvfkV1
Ju7CTDZlOOZHbk3ojlS72ZHUROVdGvZslmX7pbtVwiYCe8y227pAXJQ0k+5W5VkG
Yubdkr3/8IXi+2rMBUSIRpOXnE6gEOKjV2RR9HL/afQTgvS5otMkTU2jBmzZIkOJ
stOhML5ligfSqlaUgam8V3fw/Gmll2aWK5kBY8AF+ePkqHYz7eWUuKM2kh08ogDr
1lyLh2GpWCq6FklaULfWeaGneOS3lyZyVqDkb6voFqa39uXxvx2ZR8AEPGU+mIPQ
7NTPRm2iHvZ+ulp4KBhFoiRByI+Sh9tHIGW1QMIWRAVUnEf4wisqEYnoR8oGd7w3
gO07QHi77mVxYEjHDjf8KwdhmcZGK3dGUTRhdhLB2kzS4MlRvofqGX9x4s/f/6V7
cv1T/al2r+3YfPNP3nDBYj1l9ASNXAdvlB6bSBb5h+INNxqMmnMHDk7I1uzOSQiZ
5aHoGWxB7SzIr+bvWnRI0thEkJv4nOKqNNWzPrsqqNLmpUfrxSjo/GSzgc1KKbeK
IgEZDGw6/EmUvOUDHviHF6Cpx1mKNWh3S7XR1w8DJPVX+NR2t8Jh10ivFcDp6yFy
xYkDxUSuB3yJ7Az0DbqSfG0NlQ/ueyzGfY2FUiKnmh1B2r+fDqGn3HllQIF7VvVU
ud8WYUCTqFTIJFBHu+Vnrb4bh7bSWQ1xpvsg5m4gYQyHOtzrn9z2YHW+2o2nOwu2
TekXNHPjXUwT8/YpN0oE7PVNKdYS4z0IVHc6Rq+QHT+EmVJUmp+cvsKfyTOBTWH8
XCeXAHod1JRFa86omvvzdOu3bJwKx6ovx1iZ1Gse8AB9s39wan8BoSEPb9geeS3C
P/6iC811srEIQAhwF6dugKUP+oMX50enKxhJsUIYSshFXYho1HBonm5m4YD6xMzo
w6AmQBIlPKf2YJCwMMSEURWkC6dVsv/5YebWSQNSy/JWeYXcFVsvOc/pZpEIdkQZ
aZpnpsk75hoYp4PV4IA78k/FVFPU30j0VEdyIc4MqAxk/ZlVDep1b30h02sbm8mb
O6CHpK2IEfsbMtJLEyzWquOFVNz6QqtvtTog7NdpUibY5+3oeb2KZGui7g0wWjZm
JnOY+ZZJbGEEimXNgZYWD++jKtuN+041DI9mNSjztB0UrpwP1vic3Q8mpiwothM5
KgRSBTuVwUAQumAIHNLEpuz4AtFiBy4K9BMhx/nyMql5r0JMXzr6dm5+9dB1B5+j
H+0oKz+W2ZhFF0AIL9w8DcelE+KJBoP6OKgJYruNKAXnDjkAKV1RZfFjuFC31Iaj
sySZ+c3TVI276m87Jz3KOYWFiI4vcP3yNg5/V8mQY1MYErsrHUuYiFYSMUsw/la2
ohIy2NAq7SYxLYjs7DEiKhNX8l8GQbCYySAvmw7/6X6aee85xJe9j/HtPqnMIYbW
0ckZ3Zon2exQ4/xHGX+WUS2rVFzD8pK3OEbfAP2rS/Av7nwAYvuIRwG/QonnHLy0
pvq2f1sbk70lgUMHjHI4ZLBwN68wHayTy/BUxfemhCO/wU7tmlcvllVyOBv3FUqq
CLWTM+u4bUMfhvEqNrCOZodCUUBML1VNMpNldlPvNCk1BMlPCnUbvjgiCtkS6gM/
jbWgwhe46UKXT21aA4tISOYgL++ovYnCJ7z2O+wJiKcB+hl/Xx7cDyz3SvGAfljN
EdIY4N3VfYjbxzgny06uM+BJ5fMy0q4HekfDck3dxcCUtrmXqXML1ygLATrRYwLr
D+dctsEjxeQpaLqfEXp4Bdnxgqa6exwH019BT8ylgitXVJSi0MnH6jcUC9/+vTp/
rIEzDJWaLTNx08AGNjcNqXez7Fs0EXJ9MCj7ckw9TEDUUAdqfiZr22cNPdsfEczR
9bZHArabrc1cow41m5f31bBx6QFuTdAc/si2DZxvmK6auuSwGkR99qHVMNUDI5de
Jm/05lZZMfRne2ziWphNyueCM9BRg4le7SbAa+MVdvUSbDaqGHqSiyEy8f1k4PXD
1dnVfYVdz3x0ZMvQEbhWL4Uj9ST2YABZaWBb2/iZ7p81kA60YrGqjDXRrw+eeXsJ
fY0IjkodcGsd1Z3TC4znJo4GhrBVYaoUwlXbPU5Wz0pQHmymHP1YyUYmekxclrzI
DWns+NS1+smIyq0U+j/22vNr+RWpd0uSmShMSKk0e2ONwGkm5ntTBFM/2DjtrMlv
orrZ7wRPf7zHMFi9wFPoxb1QKB3jyaZ6WoSmhAq/38Fc9QfnsROoG5iOhtJE5yAM
Roj7dvrG1KERMIUC4yge+xyyg0yT6JYzNn3N3Xu8q/Ojkr9QGzWhVUpb2/3QrjkI
v0cuNOSIMw9gdCSCaseWXVezALzUd9ilZVPFtJHDCz8GKm0a/nCE6PZQHZOw7fJW
288elHP38ScgDNaX2/wJ3r0ZjoId1m3nsoPBQCabjXyf1kZm8/3WStK3Oq18G0z3
L023agrSoyzi8yBgjk0QRvyu1p89y8vrNZxxR3AP49stmJZiD+Snso3txlnwSVtn
4vKmm3O10iBgL2iQJVCcJfLKok+DE25/fZI61vgNnsgOXRrStJw7HN63X5pTA8OG
UO47ArOqCOaNbPz38AQEmja02EE7vYDxsu7Dxj1NmlA9vTCHhJaKFt57rlEmlu9M
i8XO1aCKFun+GJcZbhkmA8zPOIiHj9KtvVX7z8YWwE8mNnWtIMBj3L1DuxPk77E8
JfAvV2cl505GhA/k5VDwSK4Eb0x1cpq6vy4GL6cKtvqN36+Lh+JCtMgpPVnON7ur
BuLC41wGnUd5fXlEEglYBu4NmCcuZkoSiRmc4cfnJpu/xvrFFcQGfwoiFOFRWDLl
Wd7s5/8IgR510mDq5FrhuaCW7+wIWIEYpEgXU0eMi4S1u1tX8B/p+KVVGdqnJrY7
fWOGAO9wuLfSNi9ZV5lIbR69KWDdUuGBjdPvio5fE5MjLinrwLNHLP6eXq9OwZBe
6OPAN9MoD4wKw6zg12lmnRzos4w+cylIzTo064e0VFQTI7L5fUS+6+U5gJjgaf58
63ykChoftQ4bb/xgsxea0L4JYcCv9eyZPGCBIrn+VK+8FeBH/ftxvI16GRWfTrNW
H1lXBmkpEufuFL2tsBK8DpBs3h0HrDFQbo5ZZ/l/44X7NzVEx4mOxTGFrUZufPrK
Z0LXyU8WuoA0jO/Qtqfh3m16jEDqqQKAxZMcEaI0/rdq14MAPALzkbvGzIyP/Z60
Rjd9eX3GZqRUhEV3yvFRa7574rC0md7RBpSRSDRGdI6RfKZ1QOK1Y53VlN6aCGAF
hEZ8MbpYceLW2Pon5a9eZ7T1y0Rs4KVQJjTgil6cOxIwvxtsmmmER/rS37Hpxl0Z
snxdOf3h3rUFK3rkDB8fd9M7yPVbmLXnl4Ej0MwWaEsVnLQOPjXIk+bvBtLQctRD
LBm0h9w949isMBsKxadndJ+CIOX/QoQfq8c31DVVLOw/rd1umUWBPQlsyrVfZYR7
wBKDgZ9GCQ+4UslzSwhkz7xcHFChdOvDczsex5X0644YMhUvYggZt5o8cxFNV7Pz
DX4N4p3vsucPpw4N9yYD/T0eMPGRoV0va8jSnBTlUfS+2yt8uAyeJ6NHFwPwfCsI
MLGA1g6q6E0aE/JSyJWDjXpAS2tix4MiIYr1NYrADikOBNl7eF4x8PaJL44x/FLO
JT2EyKx8iYmKZvI5U0NZyWBRxVxKMOvF/70hKd0N95CQ8z4CSOwOlywX7Zsb67uk
5YNnIKUd5XraU16H3ulHAY+xrXAqz+ZnVeri5I2H4bVJREe/nipcHk50IlI2gcJL
6socXN+5Ozco0dVx8SZ7vd9UBP29WCrm3xEywfF2CpTj9t/qP33mZKfagPRVfLPr
3Yc4dLigjqGqPfUQHwTaUkW4jhdgwI2QrWolbZmXJU6GFMnxUJMe10EukbO57bx3
6pkg97IONewzee40QtEC41QqcidyI81y0OD0Q3Ce6bJeeXD6rGDF0gPMvo//0Vvw
ja7jhTeAY1xcyuHF/XA3VlChqxVQahGX0LIyJmoewXQQm+rP+Jf1g0SUWdVrsF1D
+EeWBRgmCu28RraP3Ru2fhCN8EgOc87bocr1fGeA1mWloWrUWqj/P0lHIQsh2R4F
hLIepUH0Qhkio3dN/yRkjsLu/lqnsJtjY8hfx33DtfQpNMczvd8mSJg8SyqOjXsG
JrX5yqIUUtnneditPx5TOhAesD7J8A+irZPzdxEba5Az3ZaX48dgH/gaANiEGo34
7IIlNjlnrt5E12ef7RGE9hloE1zbSZyYUdcAHAucqhrulose/Utv0rIvjbO8KhSC
rBx9SdpBgdxK4r6Ea6wnJTgC0Mp9dQdEBmcQ/Z3CBelTZI52k6OJEq3AFkN5R9g6
1akEWh+bc1OSxSCrSl0mzukncVEY5WSD5U7nIdxAWiHuO0iC48cfAFdvrVBL+Pfe
DLUB0tnHfH5PQooR1XPyYsOwDw2URsIAvB/LrdeifmiR/ke4SBd++VMPSWsDN/TC
rreUzxAlM6cWlGFBEmmQc222wDATs6YsUC13r7FXN+YBq5TtOkJsHgcjS5OzyImx
LhL/WEpJ5Uv/sxL8O9PCL2ICHeYKesW2TNipxqPgxeTs8m5h/rKTvUUKoIePHdmQ
B8tpIrlmp9QaBZwHfGSgJUH+4zagvL4VFRTCAsp/0KsAMqvidaAfbnIg33IUNMZZ
b75RRi5qDe6CZujKM3y+4nOCzmtgF/icmeThoXJ0sg6+XifG3VIKwxMlhTPmOhJj
0wPZc5WwjmpBDPLEKxupQviHnMlMWMU3JvcjzFUu7h4QHghXmRwJ/WcUhYMQAq9s
2WI6EfbNFLl4WYiTa6i5l+81dXtM0xuiFAjfGytxiBMOd/nOOYFCqnN8v/iEBoeW
atvgjswZ7UIlwBO6CPDJGgiqEw7mW0uniBK7bE7Qr6WDndu4ygFnEBo2z9IBOQRc
8+5AANF26fS1Wl57ekjPpUbkZd50qAUHwzXI48GJ4+TKWRp1T3qa/iMZM1q1CpM8
wN/2/KYMFf/eYIsUo3m6aU+RHa8naSy7NkUmBcvDd/FY2MBNfPmD0AYC6TDvGs7I
1CjJsmVYPwUmGuVU8+/I214uaFK72vdpbJDmUD2ufRLtf4+ra2gMAfUsnPWP96IX
6VR4rmVYzjC2PQEaccDwuWzNUIrNhOQIs48tfwFNqujORhDlgFPmpoQvKTryN3P6
mp+6OkbMBt3P2uzcmR0jWUbqVjFaUFC3HzBlBXm5Eer4WcyiNgs2wQV8yUpf5FHN
npvAai4SGSnE30ogZoA567N3zsAdebk11Jz6FMZXziNAXt31FGN1QpwbRiz5NVLs
KHByGCVJQEtnQnJEGY86xmIN0wyZOkt/81Z0quNWYV8e4tnpW7FuFXozlxci6/DI
KVA67aO2a+Ou2hE73QbAxiBc4SRrrdcosDzDFhIMXouUMRXhlXamFyYsJ/DPKeMd
r4uPa7EEAClJ+eWSbeNsCkPTPvDPLyqkhCnY1xoyC6+357+LYAeJIcS3goU/uDaI
a+eo5ZAFoqGnQdtmjAI6FA4qgsbJCC6XeQWtduZCxu8DAnOJY/09AoW7zEei5hav
e33GCu0mYmViN8yGR63KXLpa97/O/et5m0iwvULa2BL17tnrheRC86nE2ng0/pyX
N/nneSckhbGV/KEq3wbBh41a21axBvF3uIS7rWFt9wrnG7glx1RNsaYasxZq84Ct
t45IH57rOjCVlW3AwJmGqDF3fhfGidZrwy1twICyAj/qFRO83J5K1OxEsx3EWU9s
7QI1YRErrI5NGtYNskXMip0V4ycz21EV47eWno9Ppf2I9aAkm/Hw6HIaCgeBsu2Q
le/N4ZThY4FDq9taowb0Nv+6TsD9NV1ZE4f0bO/ZAv61FjUR7kwpgECY+PEz7N3N
hbCm1T+U8iZxG3f+kUEzBw==
`protect END_PROTECTED
