`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vj4Nn+WE7TDgbuUu2h9rWutKtmNR/3kKKwluUBthYvi4HI75so/eD2rAfLQWqskH
4iHO8MOoO9x2mCO/BRDUEfApy7+uHi1MkP4CzVdwSaol5xPzyyndKgyS7fIbhMdj
nN9ewTSa//bMChkQHDvcZaSRfzjdkrSKcnFWGCtpT1uKihPYmtH566xpVCV4YhCK
HGTau6CRiTBY5txDyvY2oH7X3efmpHrOI31tdZIdK9GhWLFM4v0aKXzNEofPX3hg
kiwsZt2gN7zTJzryb43sJWPGqmWe/LmFrVjmD6LqPK6TiA8LtLDcOEJ9rH361Qai
dzLdwmJB6z74bLSJkcEWTehhlz0wf0MEmido10hlYWdqyPnpXx3i7PWlffbUKdgx
RNKdbLtCSiVwVUmXYxzYwZH34E5Lrudw+y/j8JlyR/ssMePcwA3SWl+EPpctAJ7M
AH71Flv3v1P9tFOhnG3qlJjfRYjmDVxpjcPm2sYCIR9fxvpDROu7Jn9hBBt+C5ji
MhMBRHByzzdCtH5YOI90DNUtWpq+2RurIOKH1gUQvOK+QQ5iApTYYw8mk18JaU3P
yfWsa+78cZp0sua0bmhxwUIfCPuTOnDNblwOMiYV49MSuOi2o8w4Sgi73A8/5/ar
+XN4/IO0LrfdkUS4jW/6CgTgS0gOmNK0alzOpZyRpTDbyLFsZEgW5jzEjAUyvRgW
7U5OCP9mJ1V4XwV03uQ7wKQowMiHph/QNohDWxwoydnHfxpb8m2ZhF8wfnmJ+oMU
0qRMXVdpucQJ4ucJLY8B5CgQdlUMVML36Q1iUd03NFEemLOk5S2qg3b/czQHLM4z
vY1ZmvOt1H0kGKF8HWNW8Zxj0gGOaJC8brq8TM7FB2c7gE0HlUqvo5ndbqIWjHVK
L9H61eHEdtAM3Y33M+EK6PqEzpocnrPL7cWuFnLB6pKKIIyzVkWKPNvC51jf7ui+
`protect END_PROTECTED
