`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dp1owA4xceUo0paH1JfuU1h9a4bLUSjE+ntO7LuC260kORw7/lh6kSSJL5h/spzg
vlV4tw/Zy049csJaOnCDXqEDi9IIC1yqiR0GUOH1qzowpG0lpqcq8WLp9EJHOvPK
9Vi2MnJexIORqx8o6SI5taQ8BfblRIpdQOlFARrO6+6M6qlRS3eQ3GTCtQLXUHMf
K5xyAVXmoh0FRyUMqs0XEPXWKvZXcDE+HXZdgVhH0DEu1zFBzMCOVuXGs+3lcfsv
KYdRQ1eivGOESE9nco8rXAJkHh4yNubtR3upMLknHmm2LhkSKEZ1udR6j/vY6OKD
lKG2hP+eNxTY/7Esx1gMEGVwu0LAIiVR4vGk2YQMtCuIYN1r01RrPgBOR8jboSmg
bnqR7Tn/T8gJzYpZ0CBuXuzEKSfzrdIvIXwFEtWl2AOREAQRGALfdeup8t0uMe1h
EW/s7kl1lWJ3ZmVoOiFbbSn6/fRFwtTArbVtSICatArnOVVPIRqX5xY44n+StcTa
VAx8sdnCiOulf/o1nbycuJ2bASQ51NoBSTaPFcFLNbHgsDOZ6tIV+VZu3C+4GfRN
Ye+C6F0ZE5jICrVJGHMTJDWhc9XVmmjfW2B4UDr1kdgvm7g7Tr6va3lMzc2ZakBm
pRaN21QC6hoADQqs6riy05FnguQFwWK9vxuyR8On6/LU87P9Zf5X0NHCreTaXnTq
`protect END_PROTECTED
