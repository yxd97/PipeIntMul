`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8I1tsKSUO5M7vSykzwlJN/Cd8m0oaTgV46Kxd47PncD2HySYE5/KhKrRjYVUqpoi
XJCDAED7Np4aP1Gy/5Usi/zVQazhga3ph5aytRl1fGIH/McmdJrifC+X4ukGG35S
syT9JT9vP+YilZdTJJjNhjjSXTT6ADXoVADldaaOILZeWo7pi/w9QuOpR4mBoLAh
Xh1rk2DUTyfquE7esVpnSPFHMlnuKUrXSVUI2HkKWBaUAFSeQ5IznAD2N6J/B7c2
LlvhsFLsjBs+EKl8XtMp31lAts6nQ9lhM9fAHSBWjkIyawc96fa5UmxZJeeRAzeH
7tLzumLXqfIwVIWbCQZdNAOQetWVpBRLY3Kw4/LKRMW4RgHb8R/Y97MfE/wOCkvX
OBPQRXYBwOnVDcK96drHpFl1qYn3h1ecwn8JuTnTei0NHIiFBBLT2Te3iSlU4K2p
2UWKpJgQnQfR05cLwQ6UEVD2AXfKABZr3kfYzqlOlFUMCWfM5rjaf/G0Z4D6adxx
WyEanoDLzIk32jQTN5ibzQCALxz4zMhxuXTrid0ccRdOyoFazO/IKYyvM73NEx1g
vlXtHSfpbUOukPJT0lpTkw==
`protect END_PROTECTED
