`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D2BOEYEocZX/5aKoq9D3hGLTdVyq1nWJEVIGRke8LsUY4f3oHDs68CAYoovgM1UE
joXuJEGmEoikB6A2U7LGwx1jFu6f4Qh0wEvdd7VWb25hacDWGx8Ym8CqHCWexH89
s41YIuKFNKnqdjL7FStwL/L0kWbOg0yjYdBIxs6ObnOz/JAcXfEo+bKg9Q3pPbW1
ueCb6q51vtsINyicS7Ct3T7GzA4mDRbFiUypXHZW7RcEtEEKsHQPrhTfAdvUvwl0
V5EdcTT3J9hMLGwf4y1rdRL4p+qa8tSd1i21mCj+mA/VFMBOJv4kVItr3GSmbk20
ymlHUNItinV6FJ8ZpHfKtT+ETM50BFMjJ5SHvCVBleaKUZVI8A0bTraqZcuEoeZh
qjOkq/FHO9dqdCJOPoec2wUnl2vEPLpgifQIcnt5NQMAv2ZArMfmrdOJKYTZEt44
nEoGpPlRHutjuiKeKMzxsnDyvVrY+xhjfot7xTnEaoFPbS8+LDAZZqR+Si1mPoNB
OwQrEIBTMaCfqUEv+FeHoKI0O7OvF7nLczo7pJrWiEM=
`protect END_PROTECTED
