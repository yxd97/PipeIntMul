`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2nTylzv2giZw/9IGCMBhuMt3e+fEctbpwJukx5Bdag0l/kUVF+GbF5Ly1MVG3ZN
e79Hhhp9xP7+3ykTBCZIiXNa77KNpUpCa88Tw1KqCkgpYigrRYfo0+NrYokuc4xC
dlOmQiG0tRr3fAa9WFRu32gXYoW265bTf3A/au7vHUTQAzOhMIY/ZFhmNbNByn1J
v2yfQGKLKiNJw+2wwqUEtC7W1dZUC/vZbuqG2Qlsc+WGy/F313BlIP/kP12gtMP1
3Pi0CDRitmSwQCkqgFtpgRKf/PULxHFfyXmBvZQVY1pB3mYPkzCglW5nSfME9lJ4
iMdrIG/nIzx2xGjd+HApIg==
`protect END_PROTECTED
