`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qj0ISB6wwdew+qdPi412t8thBJHALHnOoIBKwvGfROc5CvlKvjqVFVx5E4z0yilw
tQ8bRTf8dXBrtTmhyoNgameaoxygxmy/q34iZz2YVyNz0pPb5MDFGnwxUl3tKGIG
riAdXhSPh1TLldISd3qBybYMoTsIQKXu3Pzi2y5Tx4UofImOnlJqfeC2l68Ht7DU
FOu1uVfvqQ9kBvpdyYvjpFl5lzPMvscxlbPvqvD1SyHhiLxfOiBNfOFR00rCMPh3
H1d8ewEHlpmdEfEQsGjvE/xPANEOG/Jv3Tsi0cw02Sd/ZiD+WcsVwTtrnkxOCjLE
9ouMcxLL9s1pO36Kp/Er9kFQ9PYyt77V/G1v6n/+Wc2avybO2jfNeftZgu07rj/7
6WPgbzt2iqAuu3jC3wvkjkGCU12J2Xic91/9zM3zVxDf7qumwFaOZucpSeyzww9A
dVREmI6H4cA7B/7RvsfVpqAOvrkqVannhRC8wfY5T7uhQf21O/rVtT8Upcpb09JU
xjWxlEUCNx0wZjOmjsmyR2Id3kroEThOhsbCOQq4rBc=
`protect END_PROTECTED
