`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zOwuhhYFp8GshlX9EVdlChaK+lZlpzKBE2hawfJpSbeLzr9r8FFaU4zBQ8cuKwI8
l6pY2KAmdl7ZsDcGr+u51npQ6T6iK46CcooCBvEM89A5rfGwjdNdwGy42EP3tjKF
zKYEQw22Z9wNSvp90TA4brhmIz70xZ4BHCZW9M/E7r8hOLibHKliYCGHmhZB8WF+
UyZazHBhyWTLDrweLi8LnH8e8NmVxeHw6bUe99za09MNDr1q87tepz73n/8VvQke
3OehjxCH0m6KQikupoLBE4gENR/XVaIOHjNAYMPaeaY=
`protect END_PROTECTED
