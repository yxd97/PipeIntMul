`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NK2eG30kFaWoExDdNltdQE85UpEXiWaYOSB0aKbaSjybm/R4Z3TLSqiQKT9Z761D
UlDNw/hdiPZ+0erA1hDUS1cL6O9HP+ERXpRw+jt5S9c6BhKtaE20T8vjTdu0l5V6
98WEFvVjtJNY8Uk98D1Z1R1fRvjVRDHDHopwGQrWehu96o/MbM93sF82xmtqDG1/
Uv0JmkqCA/VjksJTOZBUnttMbWw6fH9jWhkfkRRFHK9CS1u2em/kPmSWSTHEju3Z
mbpm8eWqXgGFMOt+uiUD1Odo09lSZzDMPfegHxTRZvDp+xEwJ1IoZJGNKPn+qYAN
VNqoVKcHDpqmg5He4SUftG3Wcbc+1fFqxxrLAJU9E7OWdlSYEcCDDMPJqCjILZre
Vv928h3JfzRBF6lmUvh/25fFksyQK04UKdHFy9ItR44=
`protect END_PROTECTED
