`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uv+J1v+q+39QFa+uF0egFB9YScq0rgjV/fUaC5U+qiPXKNivZD4TYH2I3xUEoKdR
o8ohV80Bw2pqOnhTxWJGJ1bnDpzwJEEmqgcw7E1l7b2n9Fb7SlLsazR+MaVkZcMz
SgftWCto8eBis1hrfn0nbFxCNEYUKoKV1dQMb0Pn9hie25PIVSGSBFacSU+Fkjlr
ZKOaVT42zBSRrc9RSh7vbxyBWjdbNxbldGExLlfr6FRgn6B7QgHarbDvtppgClWw
AQ326KtcUFbolMLi2DNXE7d+wmObrMVbN+lPVwmBgXAURyi34QVg3TCpXVE5rTVn
NyEGXijea2sbLT+Pp3ZnXQieaV4q27m4Numerf7Hpxe4NaiekzMLeaG2ADcLpzic
L8lL0LmKSQH/Au6jFbUDlADuU/ep3IqwOvJTaXzCKeu3re9qlTGkjT6/DAZCLbfP
1tgvUO3KaH9nvDqxehpf94xxuuxg7KazBYcuzwuq3BuYO0rQPRi6dw8PRDDh3spD
P/3wt6M7QkGNoK3lFvya7V6Ld5BClnyTfm/1zSnmLOVbj7IKuuui55a4q845p2TZ
CHWkNGJlr12Nky6v/0WFplbBar2lGb5p4EbN7SuMYCKQ/W1iTV9i9Vx40cSBLU63
gfg1Zf+Vt+ByNhC432wrM1DqvEN8WTxyb3MZjbBeydMI54/a/Bd46bEC/dZLMUqS
EzYIE0nCBD5viGUknJzOeF70Wcwyla2aLClqfI3BKKs=
`protect END_PROTECTED
