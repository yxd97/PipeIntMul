`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z96lawfBtMuzpmo1+9kyy3sDUiLB1nj6ala+lERxXhtEjJg0Vpiw5vyRrgFyPThw
sqQ8wQqF+f+F7L4ktTG7QDGZDV3d3fulyJbYGcEX5r6dy29gJQko61l5EEtHJaAE
+QmSv+26rp5BNaYLw0hasZhafoogWCg4cju7wQQnbqk4x6agYy+0Ls8QkT5aTeSG
EfgQvXJT1xritFcGnl/naUr/27P/GknQgtLeSE0eX/cjR/Y92SXeaH6Xn0AN7Azs
hzovTf2TIdj/SmRZEdbjaWLvtfkm6HG6m3EtaqRy3QLJ3LG1EPF99xucNgE8Kkj4
AJ4Fagka4TdRsCrs/XOCCTVnAiO/3632YpSMKRADvts4AHtM3UI77p/y2O2C+A0E
KmOQAULne0d1e4BfqPx2EkBOhAiIsvXOVfUk3dU+spDj00ShgqDXnDOXkJ0yinHc
`protect END_PROTECTED
