`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOoCFwds7yTBlcNPNWPmOwsMWRRXg9GCFQFOaAIJN4w7vaUeXFfULI3WKi66RrZZ
GnIMZZ/B7vXKFuPlvEcMiFrm80wLRYPuUraOk92+XGHOQ6jkqb8DwHdVYXmtcu0d
bGY+PfD+6Rv5zzwEUQRm215DZmwewOKpnfppVb0/D9eHn/i8L5neGCgFemNgftMl
S1iTpLLhf0fr/DH8oj7tFyiNAKmMlyCweSLGhveOZoVhnNsyNnvInJbui3I0ZmsT
Z8/CtsmNba4LoPJqx/GPew==
`protect END_PROTECTED
