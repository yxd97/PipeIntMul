`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8tjKrxKbvCzm7VThaOZ8Wt04tNEHlzZN4YS9Q+oKMUyTgtQHlcGf+mgTxG68Vh88
euIVcr52yxliep4fvJyXOTiK3lS+Eoyum7Wr8x+uzfTJ4jppED6N5Ll9jHvK8Oxb
2UjVDJXCEmOACDO4yAyuDCYMM/6gXe2d0HM9o1eHhJ42sOz2Jy4ilez4V3WwcKzT
vZKCCTGIreB+rSz6VlUtQsdDD19RaIAAT7ZQ/ZSCne9yc80lAt0Z5bjbTIegXLtc
OU6epG0XoNvrdty8cOY9XlnYy5GmZgEKHoPd0ZHA5LU=
`protect END_PROTECTED
