`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FKUSjpdfXUeU5s2rMtmaA1Ot+bmj6aZr0FRndQA7W4znvqGktZ3X1MnbgV+pJbl7
XqWMewuPMh8ukK9mBu2Fhn7OiJzd80UAltqBjf4JES8TY56Ff/FvhwxShFp8jc6U
rp/GAVR4gtMxteBm1A6R82/LkBkj7m2tpPYBgrWT06L2og7a3wFgGf5UwP+HSWH9
Io8+4L8XEu1ik+MLnLiTa950HTHzOqGW3rlqCww7z8sz0wil3JbpXg1H8mtfv/0O
5yWCoSk/dwASCsIWYHimBgS+fN0JUcoHiZr1+/ZAATrEHRoKUDieC+KY3vf7F3Uj
c5Zuq+BmggF0JZRkWcYeblYcvZv5mNlLnGW+2Ca6OVI=
`protect END_PROTECTED
