`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sbc81Oyqai9c8Qur1hT9hPH6EhRoMcog+IBdqu2fypMvTL9B9FNtvpyQCtwxPrO
7Nbh+0zNDYTrAETefmEcrleqcotMFojqZVteGXOY3EKgcYYqgfkueFBblF0R0qSB
4QnuzGrJZ1t4e11vuPelquzglOUfnGkd7q3YglYLrP6lP72Cb50ed2WC6UhkW7/D
plBJd3Rg1RFvZzcshNipcTqYD1r5GmGyShoK9RDG3Gj1bcORIlRVJJDFsqdgk486
++WMOiPk/ulRkJyp39BKdwVvA+ahNkfeis5trZP7KOmaqrsoa8xS+EoJspoOCfKV
OXTVPxehchAKX6uwZ9t/pxFGww6UWaP4gPwiS2V6Zd9dmZpxc7LuwGnu1ElV+zFw
5NE7gjQL0i9Q0fNY8EZirdW4XUb1jUBMKND6ybJDklbKYyW4NNVaUdYtVACNGgGC
OHPf3SQeCctObQOu5ra6Fdd7BnWYTEbnaMpZj5RsEFYyt7xWiG2QqpSZXZGPdgsB
N7rgGQ/XZWFri/APy7SRGzVhrURIeZ3QLDgEkcHaVkZ0iUZUUkTEE6zpgk6efjaS
SxZ/OMOhHkSbSTaO06S/1K7VD/7yHPnG+F654XZX9SlbqZWdXU6qNa7kU/JG9iL3
XSZZZlVw03Y2kyFK4aKeJ3E3EwDEzY91kU518/W1Am0=
`protect END_PROTECTED
