`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Goa0HreqV7mfmcccOq0EBej2Y970i3BaAcKWNtpZCnK1lxY/i72KrZptrkRz6ypP
ps5ST0yjop/gfr2S6eOwuSvjWMHe7kppW+VV0+5GlN4qPc9IRfQr/+d3/p+qS/CY
azmRbEeRToQVNC2RyDaee1fGBO/vMyLfzyoQuTyNYKPpBLER7/g78U6Kh8wOatCT
qLN2PihJT5wQ23DFpECeIrqIKgwlqVnwtQfPL2Kkp6Isc8g/BXifkt6ntmNIE9WT
Qj8ZB0F9FJjmLf6tEiFrzvxdfbVsWud/gVhar5XcCEH0/kZLZyDS2wibKLswa0u5
4rgp/XTVdJ7+24K58hQo0641VJpyLXMJyAP4sqr89TIKeoc3LnCogiC+1KGWMuiU
LRk1N4bgqeeEYajYCfCHqjRHA9BFf5yOLC6YatqUf8lKvG+s3KGrg+1c2ehKoZY7
aAZfclnVQXrzr/QvfT5cdleRPpn1os+4DFSLB6uy+cEaTr6r2sF4Etc/lpdeCs6r
XeIPsge1B20oJpDOn7DAM9kr7z0LMYgqH6U3C8IczDk2v6dqkt11EN1wKYrYCrvK
SIPejdPHtXX9QGAcPSBck1fnT07aEqFrxptQBYtaqxqLgDFEtYQ3BNw6d41yWWlV
1pHOJtW9rlHnD0UIsdU6t7eDvrCG8KTRsUI7PYqoBfgBQEP3p3qkF3JAuowsh3QK
L1Ow3grWsfq6vtwAtr5Kcu3ygEyV2iJkWkIZtMjq7Lsf/7SqSArRy4has5yVSO0y
jl/PLVlqZu5cZ+Xod5yktpA16VDe+mkT4kkpqdZ+RCE4AYaCwKFGwe3Gm6jFCENh
95RnNjTKwt1ZgVe6Zup1E031QUqr+VT2TvF/7lGlr96PyAPC7BzhdCU8tWlCaoZL
khcFnaOd/obBEhEOlGaSNZNYtlLSEJZ2rfWXj0ZZXTrBdO9b2JhWQToLeVpKlaIM
`protect END_PROTECTED
