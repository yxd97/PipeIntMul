`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFBTrUiGHDg5kAWPTpRDhPxurJ+ruH+JLndFN4nU3cYe1MR2kbfWEoSfvQiZ9LuN
C+3k1gIQwT9EM6G+NU7+CWDL6HkXgwCCxXWMhDbS7b+1gZvF3o8JdKF8tq0SAGnr
dNDkij3CM5BoNJeAIlwnCd0U/E3qcV8k5lh7A4At+nUbvKys0llMkYb+tyAqYng5
QbjPvnWqrmU31sBl1LsdURvHxwWpfCCXmKhNLyEDoBuPoQkSkN+9KlXJ7AoZvhA7
jhnOkPlnOQc9mOy+mCu5NcvIqs9jiGzjyO/c3XtFYNE5cUzEl/tC9bDHLfoVuCjH
80TLkDPQFeaZ3qiwdZqLEB6m0c/knNT/Z4AaKzM+RUVIEoIQNjOh7hzVzWDGQKSV
h6oNhjTp1W7b+8jShH2WYDMF148KTaI64imHCYZql8GVLDpEnRLTDS3lfcjINlzs
PqVO8Wcf5aauF5nPH8E+9GjKczU1HAVwAK6J/FHERG4imf9bReWUUZ4jj6ysQQX4
WkOBo9uQyo5hsn32wCi+GMvjjBaBwp4yhkBDp3nHCbdn7KzyObP1YomLiHmqbsVJ
76MQlBrZdb/JkPfctK6tw9zN4FZ0tBjgSiGDH93pLJyS1QCchMrE3iY3gNY2Ynxd
AXlkTFQkuxSzZ8TJmyU7MaM7KPdj2reXP88xFKIwmBeVzL9YiYF7ZBiB6EYzz3OR
hnl2Ag4VQg8CeS85lJ6+dn5jNbLU9KzlQEqOfCoYd8FbvPGiQQL5ndgZbxRirput
daD9gS9QexgGs7IsphY7r48pdl6T6yZYEgNRLHdUlqXWi3xfQNfheJHWSF+/Ry7e
c5deA51e06Dhdwqta+reecSqdSI0MzEhy6pzZgxL57Y=
`protect END_PROTECTED
