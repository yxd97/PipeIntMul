`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ptK8sO4wpKOgM871bY+NuYdlO+s3hS/u7rBBg3MwjfjBcpxjaljbxgRhetTHQKYz
Mmfz1J4Dtn8cXfsHqUgJ8N+/7K2MiPKT51K3+0kUO3sulobYpKWhYBskQZ5ZScyO
UgT+AvbOR4zPa4Zt1xeQGNS214bBI/+cPcIjdDe13185+L02e492RAQ5w406GxYo
SEapCHJpksPr60n3F3yGWD3rzQ0ad6RJGDxGVbt/9yqCsprzWcOCl9mqxwKBCaM5
ekYZJWbwHVz9nudpfwir3TNwOKu1fkury4ldlFfPKX2b7hSph4M8KEPQMRRyvpAf
eqmu7QbPpuo1Yn9WWrsbfnIQkaeAF29N9zZcHJ3v2/96JINRS2ie04OZKynYFQt+
`protect END_PROTECTED
