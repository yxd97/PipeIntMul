`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUybnuBi6g7FiYnsrSghNMjTQ1fP4yo0OMxc8lWZnamvpZ0UAgdYXEQru4liNlj7
cuXXEufyDNkostWaITgI6q4/MXBTReBaK6BF+fK+rxsVoevTc3ZGBPyp0ZYIjWwH
mLEyQPWjqUV9YGmuQ07/ebbuce36LOIvtHWmTj8QmfDZj56xJDL8A+t10q9zxsZP
IoTZJEnFGCJA9EcQfrUYu6N2UbSDEenvBU6D1zvIHuaPG65OoFxKLIUZ4O5gFal5
RqsKbYm0uKKlIt8yqQd/+ti1EsagYwvhkY7xwAJJlhYRjljPH2t3kY8csLJizD7F
PjTfXK3/x2bZQS6XU+GNWS1kVbVaLRukdtBt0Xm1ylDeMZAYUDCw4LUdCSSHm/ro
FTnLaK4DA3yOicM/Q0KnYzSbjPadgVoGN3BoDC0XQ0fOpZ4SOxQlLtHx9MN/6BI8
rQR7qiPW2boANc0iTN5KjFSNmMz1VZzW4ik8rpV4ulfMrykzFvustxYvs/ybI/8D
JV3fLZ+4kiFVpRVf6OKL66WDZbhm9IuAczEDpf0vfkWs5mlWnwOvPGgCq1l7ZBK7
AZ3tNaQ7Sbc4k+s8peURhi0D9BqAV0i11XcEMgCE6BgEQ3DqpZVYfEutw6ZHL3XK
Tv5puOPt2hmcdHNdxYiyyL5O8A7ds4V62nBoRias1ybirUJaBWff6cXF6DSICF5s
uvCQ1L/bb4ge3UB07RIYcmDqDDscpmiHLrAuZmI6FG4=
`protect END_PROTECTED
