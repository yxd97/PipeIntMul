`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
90KqelnEx4csHaOmFnwaAuMcAa0lufAUrr2ScpCZAhnoy2ksmGzpTmX6gh05ism4
t/5u2rxre5Y9xVhSncxmqd5dydQ1Lqo+gStgtbg2G2FSvNdinQSgd/84H493GZVP
isFjOeR14mnKUPEP2lVxxRXvm1g9PZhIPZrcfL/e/SF3BZsJfHaYNcBF/T7BP7Cg
Tl/3tRc+++UY8/yltvX9a2tJlUwx4LlxKEzq4KfaMrPpUqUL9gWaiJ9QLaUkRGWt
EQ93G1s24ysZ5Id3z+wnBmXjfuJ9GdM8XfeZ6lK9piyAcZ1EH+EdTwHK3N0zxQT8
KfaykRaWO210RVzpZBNFQjriJkt94cKBFIJGcnJYN5qQpAIFXlObNgO3DMhSbbyR
l6fG4aHv8m0Ta+iUdQPUqFekYaB8VlIMVJOXcVmdDf0IWrSgFoYwt/Nng5oruwfe
qIOiNuCQlf/Oh5fYpBoM9UIn8le5DHMbeOPhlQH9R8XIfXB20Zl3x2RdFpHtAI52
6lQ5tzj8QN/o31t31C0ABxMUfqa6Ly0FHe6bIuShY7szm0ARzaoqQx+NzcQ+AbhU
NY/nYbaGHG5hw0/o/r8XB8opuTE27z3lhQuoj4jG37WliUKFiOmFC8xMIlOJRkes
kVjHrwbJlS5utR/fAjn14tegKfADg5ok4nyH93qFZZc=
`protect END_PROTECTED
