`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWfVy+TiuHqcYNTQFnd8U9AJfgkJANSFG+Pf6/hQHAWtPG9CnZfZ9UKaXmeZaJnl
J7pv8mbdv6p1Ic0CULcuwwDc2PgKsDT/YZONhWUM96yvMDfGeFlGL/tR76sSTKtk
Ok7bUcqg+XWMOcLsQHUrjimHfgXT8XbE7oranlZoej65ChTxvHoHVATsCB9b3RMt
tMR9VxtDwCNVeqZUyl74oqB3WsV7fFIlS84IgDvwpx9ZI5F1633qx3olfzSMVY0I
9bFToBLl2BX7WZeaJtHTWZZRIUhr+x0NluUkD2sqqXXTTpNfwNni24Gqf1QRiile
eNWEnxo/Kz16BZ4A0SFbzeLJY0cR9Ozak1Q9tdyVwcytP//FgvW9JLFJUg3cRmzQ
Rk07LiAOFORnkVyHK6I15Qkw2uLf++0euS9LQQiQ9t5nBosr16/HmZg0IOK39wva
PEsWKrpLy8zNdnFxOoWZnYmKh3tCb/3pJnW1qTVlozZUK0/U2kAiT7aLfWylXjaC
V2a6cySjsteIBtx8M1Vin7pNjOKdo/r0VnxoO9MfPY2OfQ5FYoxb6LX3XT3WHqfi
FbziTyi1KiRI84Jbe8VGZ7zm6kkup/zTpP5/Uu5sqYY9/3KUdh1iLpTgoQIpGsTd
9vDQwcLpw1UoDB+izC9iyc2X2gpAT9MQmjNxKZFhl+9BKzFy7JpGvn+3ZR9Vq0/C
6/2HLHT0mKUJPiwCBBsYRh2vOjzVeAhSzWh4QcLqeMqv6HW7mqEJgtvsj7A2dZlW
ctWZooYAseRFxlU5saD36DThVpDD2ItgHBgdMKIUXfBuRjKPZOeyvjAEtsGm0bbp
Prc8Ywt5WiEqfKr/ZumufwwlLDav9c96JLneEQHM12fAf4ogBVCL9/fJG5163kfW
g8kGGKa39pDhC5erzB9YDkMrevXlzWLVZ9cv52g+xzSoZR1CRZonNcrnbq6koksu
`protect END_PROTECTED
