`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8ZWTtUB+4Uj82rSMpbafEbGKkeMRhNPJph81wdlmKe/FOc1AaNTfm6ikTO/6wxB
uvidhJGUkZU2zekmW2mNs2fSWjEnHiha54TVYXwR0gfGosuSNf/Nbh8qOEUikJZB
PfySkHDfIwYQEpDTdGnR/K+Kw4nL0HBleJ+I6gLnE2zPmSUj4Gxh+ikICClVjrkO
aTNQu2XXEMESl42DCv+zlJf/d2EHBHptXvY31lvpqZDenSL1PfCSEMoZ6GUY2Sib
A7Ke/+tuatRv25AcfnXP/rrWrccK1LMzfwslD+8qZb3EV2Whp3Kfq/nc2CcQzrIU
9balT5351muJNBvtX6bprhXatQK/J7JXWdXBdJSfVFRkno8QN6SXivqZqdLWMrMf
7z3fZJDjqtjvlC9PRAEmESVwDOfc/Y4sOpRKal0a0ps=
`protect END_PROTECTED
