`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5WVkOqkctPRSllUqHy2bmwtUMEHOuLykY0DJxTF5z+Aik0IQ8s/VLghN8EQSo3E
A5YlHy1sqrmtvUIwjpfnz64FEoQc7bMvOsC6F3rpeq1oulssVbsIE7afduxkBzxr
6POj344bM7k1J3yOuOoPE49EfogDJMiIhrAaAwh5L1TqPIpRH8RKkRxESbYg8c6r
i8EvEzxGZ0SYbka3AWn5h+vp9+8p9+yo5lZoTRLcgoh0fmXkash+xTthpEij2RoN
BEuKLlRVAfH3CaaEl6rGNsKrJoCeGzI2HFEWtD4F+uw7J0PJNb1/ZyrGL9M/Zddn
t951SH3I3m7wGQk7k9DGcU9vOk8DRTT2bxIehDPBjR8=
`protect END_PROTECTED
