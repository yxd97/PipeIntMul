`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ed9mZlrmbg6fPWyWJyHcLw/+gOimMUPDUKv/yelD/JeYWYfR5U/Oax+a89A7MlgI
qbhD8lo+YF5IF6HxsQfuH2KuNzWf89oNesbePo6NxCyZjFefyNOIiGcLkXEWhgbU
j3Z02T052weo/C8sbDNIG5YKqg7acQ0nRLtMEmuFGh2dDJlsE/rDNyfYigMcbFQ2
fhXZ3RR9z/Lu/JVOUxTCQ8O2H3WIgg6hmjZGjCr7j/CoSL64Gs66oQ9z3cVnS74h
SgPOc3dOUC/8HjCAyH8d8nAn83fyc8YZMekE5iKoDYfp3TvCT+qwcA4guAxjfK+e
ClWGAtcL1hbRzqeG3LXxHtthY81pz6+kLBzYdS+CzexY3HhcE5eTFgGTqNrblu1J
+0wu6C1jUnfTGfaDx4xpUVqIuUUqWbqq4+SqfO3Q/9r8SYaLSGo7MZceXhTHTQZ+
U4QotYp2Xygk/i28EeaZ/L58Lobq5eOr4tnnZekLAP3vT8uwChZeUzTaYYyW0qGE
QCScMkthzSYfBwq8IvbNZLiD7auhEEvv3lw0MupL+Vl/UMKI0I2xQfhNDor8roWq
LvoomJuztllVsXKEXbWXpY22/S2n5F4n54sWjRdjk91i9xMcHiw/XwRp6bmX3E+j
Mds3Z2yfwjSp73LKHh6BJSmso30YDv44216aButQ/JzZJw+BStWa4YnPSNdU0r1Y
GjLx3te/rUmWbjRkS9V9IoZvinOmqczBjZSPZwlE/7FE4wyMFnlqR/efZIGpyXxi
8LZyLQ4tw3r8/Fyr4uMwESqfu77LyjgcPhAjLtvBUUbCPFdtRMpwuZtxbI2cb5DO
uwf9WcHug6ddV9vmIiG8FENl3gysijHlz/Iq8WNT9hIQOY6lQ7gdYwiMHKp8QHuq
x5sF3XH99LegXfrkAe9xViyC6MjARW5UYspX9G+MU1MWNxO4Y0i/+2OQyvcspDvs
2x6OqskU4VHv4bsUwDQUkZ49btphjtMN7/vq6J6qyA8l3ygpqFE/hn2ClnFvEk0P
vafcHKjzAYGqgsI9g4GVfjKwUJCGLcSfe6gspcG511HOUwEXAO+GBOGEXzvS5UBn
EYxj3xi0kbxOijyWZTnpqf+WjHfvWAtWkZi6rdRmjEFD07fwZ7wasujn6DFRLb6s
BjZj0c6P2V9VzL+U2myQScnydxiQVMCG0Mm7oCRukP/NGwUvLbtam+K+64+bl7qH
M1e42MHB8/f+8QvVVnvrDwhR+y3Lh8X+b4ThinqroNcPu9TDrTAm10rrOFJ+8Ghq
H/85eZFMaVbpCuFRx96AEd3J9PLCrXNURrLOztrYMWCT2ez4nMOnFf7Me/Od9u6P
8yF1klzZH0iyJh2loSGBBl40N2XF1jhjDLXFUvXm9iHWST6k1qVPNnxs+FFOOnOv
YFQJAeWvwxummthPiD9vUt6G9hDC4bIqFmeUn8qNsYLHemIxjhLoJsqb/fLQBe2/
+CTJFakW7PFsJSNMh4dmNwJOY/gsnwZ2yrSmqJTlB8HcB4XErZ13tH4KK1KJeSFI
OQQ8RENQOHhVH6vWOR20ta7ZDOo/0LtJXoR7N3wBdjpLqKwGURy4xGJawBkl62qB
ARi8fOQyHj4tTOtKqt86SikuOfaGnoQmucdOEhVZZ2TeOgAdqPnXnCefm0vGA2g9
Mp5k7BzpLo5jEfZovSgzvM1mTyy3ThuqWo71A2RQdSis3EYAIZP7a5SPAB5pQhfx
D4l+/bUtsN+xTcwgPpB8IQKev67cRZkXmUr7Aw2P5loL5GXbSYNnimeOWUaIjWio
VHFj2lj+yYl6siR4QxN/AGTMD7CqyZ2oKzhTfNgDixKSbTDwFVTSoONQ+ezrdzIl
9tqT7JhT5bgW/ITTsDGc40r8PO+oE9XxK0Yhj5HWGgaWjaFi0Q9alMOqNK04vWcL
3AnMEk3OlWcUo1jnrf88hYbbAcFYMJW0FfIY+VhrXTm0PFMQiw52kJRNdsrdDuwR
FrYM9VuiDg5jaf6M+xqI/O59QXHbXeqQpwp50XspbcmAKSXjGf2aXu4JxjUOKk5M
z4rO0vqzIYpi3WBMpaFUJYRaoqomqGIxvviWhfNrO+4d0LXyYlywFU0UI/PSJF1C
m25kaOAMBl/4WUXaQPbeeY4tL0pGggbjX19t6gOuPszxXbsPmoOy7ur2IpgQjCop
W7N2Ar8zygWsakGdv5IaAnTjHAIqUQ/H0JKeIVD+Fg2I7VbO8ct4CyEZDUuPRWNw
SRSsBgEBkafG88ANeyg2Waw7oPJfHVItnJHzmJOlR0rIolIlxwHJJ2XaL+v/fDVu
npz8io54e8KstcW3cQos/dZf+HZ91SB3UpFJXoXXMXQcw00JFxiNkGRQd4We8qUp
n4506l960/gZRXGcnz9lDpFOSYpZI5oWvAp398nfFNetG2Pc6NjKbT/0JvlNdtUj
e/qo9MHEfleBQ2kHLZK5Th7uNIm2F9DT2U6oM4MJa9pAz5kooEPz2mdfDdW8RYNp
1U0ruhVZfNdM7A6l4R9u9BdqTXgdYmhfYlh6/GQg7UWlC3+7xK4yxkh8Rwht7PAq
Zi5XrjlR4gd22endWkvxcUVuqNQMXYZenVoSGYkOhHtEr2C0yuHcGMDJl3nanGon
`protect END_PROTECTED
