`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGXavWK6kARvrg9V3jHSCZMsafPAGLXdtZaxjoa+Hdj1V2B1uAs5NPUiXTauv+ee
CNinm04DIgyBMtsrQXfPaFjmJCHPz1mk97eAQzZeCuq7PvTn+2k/F75FLHtxVv4u
ldMX4G/Zay87HUyNlAz7Wzw5KEIRTiOT33vRU3ajOG+ysrEGCrkvlxPMryPbovgS
9xGGUUX1yUWAJZNy72pU0MBJ5MdAlH05KYhDwuHGbLARpdA0zKruuq/oUgZMAbSI
YixgFeknBIojSkNF5r/D8JW8EfyXa2eld/OwhyBdgeE=
`protect END_PROTECTED
