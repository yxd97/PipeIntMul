`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5x92kg1J1lnEa1PJpW9X/EExaNAz5HuuCFMYRY35a+3oCRZyDQ0tN5ya6fWMh9Lz
IdZQEbASuKj6juPZJYVEbaBy7p+oIHU9ZSnMIHWTLSYmXHOGx/NWjcadPBgG/C89
4A27A4wRIQIuD4T7vOjhTuU3TJDIX8tg9QGcKy7vWAUJaCfKi+czH/HSUn6/o49R
zpOffBK+qJPArVTVlDFAdgaqp3rU5R0ddBV35hvEv0Gmzg3OJrvXCdUhi6g4H5AO
++/EX2YOeMgHPXQhMIto7atQNdA+ZXw7CGGtRJzX8TlKnk/AZ8AQ2ahOxXiYRJwY
RvlsyNIc+MkzixVzdLdVA1CEEfyshVPAmysfeRyZ8N40YgM4ITaJ0TjKRpwo8jSS
r1/oNcHmz4KFL/RXmuSfvtLng7H1AZ4bPID+yK3R5wvBPahiPtLKRh3Fm78wKhvX
CYUD8x2YXsb42vnACs/+26KcaGJnVHrLPdSFAl98zY4R4AomKqGiEUvtkje8RaY/
4nH2wcYXH/kMdgIjQON1m6LSC8VJFSgGWLKBcR9pvA2rno/Gmq8w4p//cyK3/UqO
dLBJvWeY+FMFfOfc+10MXaMklrOIinUKDLH+ldjOdsvDlboRVh8cpL5i7V8FzeKX
fIn8wNnA8gm0lvgYVMD65R5o6kpXtRJaP7EgPSiWNKQyZ1QMVZna+kd44Dn5YFqd
NuM6Vgno0IHk5N8Qdl/yMqSwXWwEc8DZkdAi7rIxi0idtbwgvt/KcEAvX3MzqKwn
hNUhXYZRW/hjOAK5j88WLampOlxsQp5CzlCltd7UNl8=
`protect END_PROTECTED
