`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/k31xN2d3vnrvmMc3pxZ8yN4jFhupv3CV8wqzdaLaFyYQ9Bg/zs89JAlpwCMYReh
h1xf14qZEuBm2hB3bttntnkbZtcGFNjVNlUlW4JC4sXbyUmICuY00tnDUkW2eV+X
7l8vU6mxvj8QwF1NaKD/JgIMzsIOe7CBEDBTZ3GCoHwWFQi/oQN2fuIfkc8x/9W2
kc/3GrlpUgph2FfH68JH/K5uo7b5XXotC3G6TGU5OLbLAJo2lojGgIGIxrn+7k0h
olc+r9tkOzcZKzugE5RGVx798+70fflp0M+WCSXWPQRPkehE8GLjVbaTUEQwFxKx
W66FZV6tzNTNuE3KqWP35i9Rf3B7Z8F9hiFWOOhjT971Sh3t2TIzP8z71lKTwfzA
agQ9n0bObrGigfjl6z/lYOWDoYsXjmMqgIL2r3HJB7zVJaG3MebslOU7vyB/9zyr
Nn1irZdlq4hbkTxDTpEaarzYie7E9Uv9ArHIDn6aQd0sU9XA8xhvSBDK42cuyke9
k0zr4DydUocwlEAI83ij6y7n3qAUq4ICeOA8vRGdl+NHfqBjvxgmW86+6Fk+Zrtg
4+H4lAmGInE2ob9+39d0ExnXitV1dLOTyBBL84ABcZbaEmFwApwI/H/x88N5Jqmd
oeqS/ov+N4JKsu9KGN7bMkJjGxsQwuGxcrYlxmyNIUXMo+XLpBbZf+t+zhVS8EJj
U9ZyU++mjxv2VkJsBlnCw9fSdKzeLIEq7nS/7O9GwfePxFLwzgENFcakaHYcb1MC
lOaD2Pnvn4SvzTTGhrJGItMrh/6YHR8cSgE2m4ywj88RGWwVNO9ik/Q+z9iUxB2I
eNPpzwDOBQbYWixPLOx06MqUZXaM7GVHf9ggeIiy+KGjb2qKI+bjVzOhu/wkBdHE
diAE9e0vzEwKVybqEQNeJLWgDr2H8ZqB4AiZq8urZZRSmuDvhNeI7SjWJ/YCdIrh
Ey0bSHhtThR37Fd77smBCcRy377RTW6nbA4JnACR397sycT9fmTjfKYBGengH3JK
zbk2NsnZUTzt7GKua+XqOEnfDkbFs8sOFpHnTM+Fmu6pfOYuP3P+Cp4Agy6bQ03r
C+0Dp137YEwJ0tYiX/y5dg==
`protect END_PROTECTED
