`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NUTIU3jjc6WP41hzyQnor5YapWkwYza1TDiQobbOw8nSFN+DI426bZFwm6fOpS4X
IIVNMqGVweIjClZ6Kf3bGRscBPGpmr5duHAyhO3vHxFJmgAgREn3RlrNLT0NWlqw
4cIoBsBa1P6UsuX0fmvgY6rHZyhAf4kNueNCF9QuXqrSPGTCG8r6uaH5EHQM6xac
LvKPhHknsfWuzCz5PFJUxzAGHQ8xOFfGiDfxLMux72/rrPmggi0RlngIPsJSfgeK
/ySz6bTbz7pTekATJlXc5IzuxDBpFR5WqNye+3JTSD9A7nvMw+P0ieFaRGgvHUvT
ikR1zFNbU0cZYfGK0MJxIZK4ESOvPtJsnnFAbyhLvKNNKEs6GfAEfSjoyOFvwZwV
i34pDk1g7JA8PP1HOQiSwwtEOPf5aVe1U6itbCuKwWdEcZhKZ4Qkd+U2tjkvCefV
JhHCqg+UjDT+VvZViBnjVt+HZzBh3ONlVVbkfyNQVk9lqRcCz5Aa56/Zcc8qM1Mf
CZMh9JbOHS/nwlRvvQtTievBaQrDWO3TSjhyi4Zc0Hkq2xtMU7OHGb0n6ZGPr/Rz
MAmTYt6yfraHK1qD9+2CwInnz70nARKmo3tBhR+ymV76QDxE16z6zsdZ+2vckIgV
IZmRnzKzDoVLp47ImsZYsX+Kfflr6gUuC1CwoYzCUiSGhyWhxvwsNbAmTw8d6c/g
QF+rKDa+NJXX6/5VKhPAp/e4bIryCNahiIhcetB8t68ILwmP1IlRru4ZsEUaU4tS
2JFAGaC7VACE/LIssrIIhSKY/VG+8CUyqsM47FpYc59dGII3z7JusPtxMa2IDQLH
y2tG3ti7t1I7BI2SR7guOz4k45Z2l0B1vWilnbn5bXaytNisnGtr+nb/wRq94aEB
5flWqXvEZwlF3AbdFgctrebYbLmT3EwYU+m6Qb+OtL6+f8sLnchttbwk6uymniYL
`protect END_PROTECTED
