`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m828fIvp/iEBJO0tJ8n5CKm4ZF4zDFQxnH/DmQIx3UqziEG/BYY7FsmR8ilx1fhj
ggF1lLroxDLIAvgFtIuDqxlo9RLfIizm+NOO/iTfTpPoxnEy4IXEgR7JqkgAL3t7
ye3poRruNhuHU9QdqPnHx8AwscXV/ban3GL97eQwgRhUunnrnABcF4GXPLvIvyBB
N7ccTC6WMjtiP5l+KelwLJYqyEHzfBD1wle3MvyjZ2QiUh2Ml+O7bl/NC/rdZRRG
aLPil+/fL+1Vxq8p2g5xSPxaq/j8V0ChgRar/cgiaAwoz8NJByjrh5hooa5bQ4md
rKhDGEmF9v39LvH5GhoMvYRNn6nc/ecaRMBGImnZNkD6gt1z/9OcJS3ifWpxg23L
EjRGvBXJX6ZW8cip41g3W3QUjNocBvK/GfrWd7Dw7hAsZczTYUm9MNDrwR880mcJ
inPBTkCQpN6sucWlm4IVQ1HTYFpwFGpQBtYZdTDj4152mpCh/eqZ1VesFvaZA1RH
/qgdNuv4qip/2z71o94N6Gu0QmOv1G1d8vAP0jHGEJj1icr4gjfFHv+ZY4W7uXEO
`protect END_PROTECTED
