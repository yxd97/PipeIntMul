`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4CDMCaAxJ9I6+5MImNjkrjFLheb+CQIsOib+8KIqZ4LCBEGoV9tk3HZnxYTDrvo
ZM0NBLE5qHByfKehsyaPwHB+IROozuofCjYERlZTBPK137AVLKExq6PqLXukj5D3
+lOhotBeNcGX5ZX+239MeZEAm1TOFlnTFqvU3OkRmAXymikU4jgS2b10sl/E632c
HaXoD+JlasZSNVodSS4VusTiDgZKvXhn5qsiemei/lYsT7fIEFYxsVP8mSCFHMdL
FZL7mxmzRgGJmxRwgasyzZghAbvaG8/e/PqWSsUEC/iNB9KKPUWre0uZ+pBpYfMb
vlT/v1iewxnC4+a/+DXVBxR15ht3baThdgueZ8adZ2OtlzPpltMNy2t1XrrNwVaS
4lTa8xK8vgMiJqkYeShvJZ7uGnQyAhcWR/ABkef2MAuTxbwLj8Qv5EzI8NcoG05B
kj4jezBJbXOwLop+4Nxx7g==
`protect END_PROTECTED
