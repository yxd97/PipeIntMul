`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HARzegLRouIjvi7AU97Z6gqy6VPDyB0Y4v7kDYQJr/SGYGLR8VA/6QObKLUCKs7
IgfNw9AwDAHYB55XMUrpw6IG56m9YJb1A9iohjGnthHZ0+x0C3O9W9J4dvqaJFXh
DGw7guhHQtKdMtBZs/T0+t8a52fcmFwe83h1LlZ7Bh76w6P1r/G7fkD4C0iyKzDS
oRo4ZJ8EOcxH490MaXCjc+vQGxkNNgwGt8VAbKh04+btRBos5QEh/1hEPFD1tZic
1e7VKSb/lmwxoV6QIfd/aH9LS53wAXuGa/g+/y7nlcI+StTl9LWWwVLS49gkN37f
ka/p9wcJnRlbBWpYVXh8UMBcwlM+j9FhasreX1Ypa4AENAKYHU8wSkfj/lIYtVgl
cOoBKH7W9xa5A+EHrrfPbydAactSaU6dBlm+hUDvi0TFBQ68oMwytssq4HOd9PSf
g8W1d6FNyNGC3UG1bvaXbLbROl602ifjBmbiF4ulVQw=
`protect END_PROTECTED
