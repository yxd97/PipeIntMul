`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AMwphXW5mnWJznFKYN96igZ79o9hBN0uW4XKj/9HoLe2yfgFkH3nZ2jC1OekIG65
+07MM289F0jS9Hs7CZTU6ax7FPciq8Oq/ykHUrQUe4KIV/BqXUTt4Pmf/+ORIltv
IFZjaHgIfq9boSS1a8Bt0GCk2URwvaTug57c9HsWCMPIFLmXtYTApkIxYjleTEnW
FhL9mzyCT3Y2rPBMxc8MSVhtR2Zl2aGgoBhgcIQ6+Tn+zZp1QCxa3ihRy/w6qUEu
VtYcJ0DFqFAvX72XlEQtvJacXdc47G21ecFw6G05aqk3wt3CD7fbVnr1RW3rq+Gy
eJWvUO6Bth7VOdwHQ2P0XkR0UN3aWl8h+4qidWV7TtmVvPW3r3bAEwgDGTSl9jAt
RZSJ6yQIOi/aIi4LO1mqkFXPxEelmSqoXoTqi9WrfkBHx19J9Lqo0tQDjE2nZr6s
kK+er5+lzs5fAt5tvxatdX9jyxsJQ9dN2ME2KkJ/ssDw+3DDvKEr+AqAQ0Im/PWt
Qj0K80sP0w4lrBCfTYPtvU56PE93dftC94Ws7+6Vkel7eDMFLRu9o5KxlPlFwCpI
0S0qeGE9+3Jv1t/Kwe44eKAC5e8DVcIsGmbxrXi7Mh54PDorcCJ2ErzW2AaOVV2B
5tzi/tbZmkwJ4bAFvEUNVjkzsWwrz7X1z2N1Yux3DFTUShlgqJtQ0KggPZlGuOab
THDDQQRuschiNWLa2s6DpZweuu7qAXX6yVqeRMENYQk+snxP0HqOg3kw7GfjPaOo
2rzL5E4buHCYK0gT4OV9BXogrwfo2lYr9Q5MDAqz4As4+n13wM8N55ClTCUN10UI
D60Gl44UJBri/Z6wWLf8AHZr88XQx1CvO9+1QQHPmYWisLGVo6eCyq9tQuyypdji
3GjwD5+jIwxP0uLn7fIOyEWyHFFT6wgqYZTLeXG4xQ1vVpKPKeSXS5Kx+LDFEXYQ
SSklWZF/cbVMRkvI9QedjBTU2NrRv70ZIncPda7y1BWCNK2969I7r0b1wmJKDAoa
iTRdzgSrt1xzQNlgETEO1k3vejsv+tBCbox8zMh+B3o4zq/omXTrUaUQ0L5ihBUA
kvpBtZGtvfEFJRcm/HrTIooGIb8wMlhv1oNNNLjpHtrr31yuBqBz5vMnmr3YYY1O
x0vr7OqInIvb5W/RDkzDQwP9fg+Y430yzkrmAdJ0V3xYISfsKfTOgDwCkENf2SZG
sUYItc/fSf+5D8AMlu3p5vtPcmcKhJbfp3dUPA/hOj8p6PJnqldkRSo50QQpWVYi
`protect END_PROTECTED
