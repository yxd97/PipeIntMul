`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WcNsTII2GThoXaLkOgiZYhw47zjk42JdFTTMYDZjvT1E2+VG3stavSAFpL78j2cu
0oXhmo6N/If0TYU8OVHi3um/pCGNxZGvQKMsQ6iECgTbt62HHUBkrLqm/J3cHxA0
OINDCNxT6kBKPGGtYVETGkPRuXSU7cjl8+XHdR2pNi9tkt2w7uq0Fy4ZdHZ8pYYM
V8Ul1DJmuB7YsbSQSnr/bNV3pd2+ZAyH1ZNLAqJmd9N5pZqLyPnY8UluCcXwIYpd
MgL7nvAb61h/wOIDgH3NaNeYATt7VJVbDWUd6CCgKw2rutbbn3hGRZpi/m+Ik0Pc
Y97XLWNKyYlUKA0di8Bw4gcG5Ra27HiO9BIV7+dU8r/XGLIKO6Oi8EiLr5L7F9on
cKlIzyS1cmhQMugrlIC2eJholFcf7ek6UfzWHgeYOcIIys8nmR5xcEaL2H0YogsU
ZAA1/DXhqx5pvtuNFpa+5t+inrIJFBu5QYjUxiVybyfYxy0B6DyjB+C3Y6qesMw3
`protect END_PROTECTED
