`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fbL2og8IDLGBtLuzgkOi4+WkFpLg3vQP5lNHUVFbeWJq73mzCZ4UZKC7ucu/H9Ok
XT0huLCTMN3DpSccHaqk5cIwLUyqtBM6cAVYRuU9XTNDYvEp8832arqPG4XFq2r5
hOLKKAaJTY7xIcMrjmBM6A5yGL51Pjnblyq1StVHxK4maVjtgq11iL3Xt1akLw/o
IYVGZuUIvYAjjilM1WU7B4VfGigX1cls8vkQOnyX8tfYWMZwyntKondUmAjyPU2H
TXzwtlBukIqnN5W/vha9ghJVosTxrIkQnFLeaZV/fn0=
`protect END_PROTECTED
