`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bD4rlyhoV7HQ2jtmqzSbaWu+H7iwcLF7+6C4aeGA9LHpIXBTgTgW09PL1Y1Ubz7N
L+7763yV/YWWS5pPZbzf3Z0i4EivfmM1T14r0gOiDZ4OzCj5W5f/MjAUO2yujPKW
7TSEiyW2FCkUHGimivkOS3nyS/LAgK4HFLYmObn1S7UefKImyl5qEA8JQ9Xt+9Kr
ZT0ujLURbJ1sF/tW5CMT+xYFL1938L/MifEnzUHY3xHnYD3vBlOMoOvfgvxNyx7C
f+JrKkdMAwY9skOwAA6xkV54jKLTj/PImlo2K8+/TzNJIdwV/mokL5SJe0qly8y2
E/kDjyZeYSvhWZpgM5M9VOAXaONYXY8sShmJ29VN1Tnwm2stewcFgZsE3N6DJFgm
7hNwAPlQmt34ScsTO4RlC/ACszmarahahaFlZOTtstolkKT057Iyl3eSgFjuSjAV
dFruJTF/0D+vqcxc2Ddt2leUPmUP3S8Fxyt3/6U0TarwJ65Tpv4T37Bls/NkbRG3
`protect END_PROTECTED
