`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ERMp/b1sV6Xcmv28W9xCqVqjoPxVq/gKAHFEzwEhgNyJ0QzijYQ3AlhCJZVYyl/D
DKTALeR8RGSbzEWEgwIYMijyYT/h3YDDXqoGotuFD7LyXKX8bEIUaYo4kc+saYZz
uUhrb+oqKiSbkUV4UmRnle4r71NT6LR0Tz5XzxdYVsnpzuMj2TYEo/4rVAxi9rYb
FT5UqLguW4Zr8K8coSSplFDZcBvXsiraVQgaaMMEunSSZnPV5M05pnNc1VnuedO1
tEzurGSO+89wmgntFoSu96VvQ7cHCaUlaQKHva0CRfM0HyMM1wlgR/L9hR0JazFl
5kHqPUncQXD7/7Dp5aNF7kUOfr9srUEdOWDwwNo7DKNrDqxSeJdODseWA4iUtR4k
EmUoY+FKhkL+hxLpwexz16ssFPv4iEtyGehNMSg4MmJgAEjCfABBQ6XIgrtz7RlZ
M99px1CTV+myC3yc3NvTuptr/pLvArKPwgaSgc3QWCV8uE9qF3hXooLK3IIkSNlv
PD9LuQbFF69zA+RUn+/y0Sbw1rAoAnmjq2IFoD9b9ZlA6RPgJUzqtw5ZViEojYau
XVXSgHSBfaRSNUK2WjC4pk8Y+XhJmhXI+C0ZCoxQmT95LNQrL6DfdIhcBTD02uR/
vwBMorMa0MT4CfJstYDOPUNh/7BKPhN3mww32E0aLpD/4VR5h4bJJuQTcZbdmKyc
1we3sO6rh+n12mk3xxQiLH9kfE1FYw23hWYxTxouF3rF+Keg3bQytIyCHQ4nVL4Y
vGGYxFwTddzRAupppzMYx/51bStURtAlK/xX/2yyQXVZe9gh6AauoGVpJiU/7z8L
5vqSI5qJO91MbRgjqPBk8rGUZ5QMJAAwhbAx7BXvMjLR99IiSNCO+JvAGx6wfAEc
VM1GFlhlrVWG7SjxnhDKmkiN/nDZYjiKCaPAcd75zQd5l+FUp9ANmzNL2HdhO8n2
XtPb8gFj7DDo2Eusu0ANcUYQbiE+kYo2zzpi3ulSFO89eS3R1R7P1+4JqxbP+pM5
OoaKZb0f2vqZMZJacfeqapFevUYoM5VK2c044lpeYlip2gsNVnk3Ngz+qMCDRySb
oT0CedTROALhKUahfmWleGe9m0bCbHEXs/sg8kDWujY8S9ft70d5H/ulwSFZgX5Z
JEgZslG5U8JWk05bghbB9Yb+8pAq86dm+70iEbtZqc5/Z2oNsDBpQhCisk4oqfOr
gbBcZRU0pjh3yeQ52Dp7z7XtQ4Vb8OkoO2Bhn99M4otMIU0CRB1QU6n6rB8fn+Oi
0QujbRmbbvEroCV4RfNJSlITR1WNiVMd5h5ZCzeyOxYxIkTPxJi1CxMks9G7l2Ep
wv73OYNxD7e0QugCphoDP1sqEynoH4RAGLKilcOEhUjSK/PqdyrUV1O+MZObMh/E
hI729zgSVhQDrmkTSH91NtT8rFY3zegaXn4TUv8yOIaPFoxekmEUM5EpOpQ/NnFC
F8HAjyICSHG9ktDmSmX6lp7pnjzE4iUKfQQsqPXRekp9HjGGR788/Ukh1z44mgm6
faAKJci6uepjUowvFxeHQ5LMvK9hwY6RzpN3Awll/mTNg6jR12GHLjaKBt7cg3SM
xMpuQpo8oG7iN+Gvj6VLAcy8rER9j4kxb2kOaHc680yjh1AtCfkvJ1oSGEp6w8ol
BEVUnsbqJ9KrEIBuK/txG7GyXAriBqb1sy9AMBlLhMOkew/nd18Y00QQGYT+gN6M
lWt+C9czbXcOmg42Um7ZDv5wISrToQoWINitU6zfHDVvxEDryVljIo941jxQotRL
+ByUYyE/hewyWGbYGPR+guHmKbM56IzBiqagWprfg1TGJRpIuGSPw5JED00jf5iI
d9Yw4ZhHFUzJ4KrOrtwzlXcyPIg1FR2xSJZ5WFN2oAMqv5rlsDgUAnUHM9uo2GIK
TG1jC68si4SfbzYYOhR2xK0qes+FCLPhnu8oiK8v31OdLCDIZg3YVYwCMnp9tiY+
WLSHQqTMJYIhmFtvNFeFv2Sfo9Xz3sMLnon5F+80rOZLuPjTdTpBkYtrvNSIoVXt
rKqa3hlk/JJvgjhqm9HkHs5djIl9gS3NTN7VUauSDFo9BjnV+19YQtF++YTdzMLt
TXBISHijuzKQNPaRJTIxmiXS+vkpoFlK2PKOaq/lj1UIartxNAQVdqYFQLVOOJHj
k/wMl4udQsmzIssu/oEpcN20pj2ziHjotiUqUEEZFBBMRQSpzOf1InOZ7Q5hQzB7
mQ/00PENJEj8kIFijB/20EaMuXCy3ziz9JHPCK1lA/yd7BMNRZXGYgDD3ht+i/p+
x2JVUNo9xrZ1nF0xzcbfom8Zup3PFVjZ4fGTj2NvXSUbR0jmHvjs4B+oESXeY8wf
pCIITaVnc4pVOa92IduTD/AvVl9SSZQ2UoQC1BagDKXPbEfYQsupgU9YHOhZF4Qg
jAokYXO5c7zMlaygov/lyaviO1NcwwRB/T1fzV75m3WHXmBvuhYgPO5SGUtfIQUM
lUlyl6a7tZJgQfxYtIp0hKe2eabLNgW/dCAh+S9ifBS5lKR+l+2VeksjOOJhhdL1
pNQK//s0ThazokhnVGG1GSxYnmVvyIu63VJZxWgRSd1Hi0rZCaI1o/Lgc2oCWPpr
oy+tNfc3R8Zyoaor70sF80HsuOQ9zxDPsZXFEBdBdDuW7Tv3/Te3Ha+pts9wad0p
B8pGIWl/kDCRAdcmf7niqXzGMZVSLYSw2DuqjF/BvLe3IZIj2XjuC5Tq3x8YqbPr
ZsID1n9IqLv9q16BAxeGdFxspo/VBZ+yVh7Mv48LZmUweQaPJS2i7EGoK6NjPkOu
M+BpacOUGRwEfa0bPyUT4hRNRXjxuRkPLNbButeHMqzRxWHVC5mf12vNYKkBopse
v4d86jmUnXIJ7IKljesl2RszpOUR628wd0qrfydWdERWkQ6+Cia5GlBQeDnasoLH
Yx3WKF//C+O1Thazb1qG3oGRaJ46rR9VTv1mODaKfalMpR5sAdLfnHHI6Y4lwGO0
vOBJAGjEZwBZIVAyn2tEyWzk1ow+pPHvqcpSY+y+aKkLKDkEuzJDmpMyW8IHgUNL
B8A0fXCEOYaZ8arPglEz0ayPEBp4QwpVI+Lq779ZFDfA40mcNV3NGk3GdoAk9EDD
9ygO8xueN9YdNmGpNQjF7U3KwQ5hL/wYAFpLK5VrKggHhygoi2gSUXqULncHNsI+
Ck6/JBFWf8jNBSex61nZvlkej9+/N2nOZSGdTOcjrx8g/AQYStHelhurvRxyRQBU
xLvtc64B2KGpKN4C4EY619p4e/UYLN55kE0zL1YN1mEGQs7vaRziGypq9cNMmEAI
cW1lFaqqVNI6pSM21u8RWE/yjuG/3LGMWhNVBo7h/Ma3RQXfFZgD2rqhWTcDSH0L
w07d8i/C3uGMwBa1u30Vf9pR6cuOfi11NHvgcEJbYvAR88YGqaAeNbUOif7zFaSq
vl8Lr7NlfEzYm2XH2JW/bzb5zTL4+giGGsyOu45QzwcNFxbPStepty8+12W/bHh/
tHPv2Xk3SMmF1yvVg1/FrUeDtwGb+Go7hEEunbSkqYLOOzIK95r2P3iIZwVvNZqW
7x+Rjw1Oxf190U9+fMn2Yh52+GIuUBTvDZwNAkBJ6o/E4yFcPnOJ7bCm6YmG1ojf
xq0M9Zl8LQwDk1HFbX++PPYlhdXwASvYwWlMFmG34gLTO7+DZe02cFNKztLzHKTy
C1xy/yf7baXhHrceOL78n1j81Xqyh5f5EHOW3eQ/XcOu5NSpGbWrsaEM1D4KBGrr
juiQk3lSPQt5Y1TzigM9VJHqDMa9/HXgY0AathbzMJHeMmGcjEP+eZNUTmgAp1/n
E/IgXVV9smwWGYFkGGZVYvLdgs0p9c68QMrNI4gf+uttCJM3N6rZ0zqDz8SB3i48
SG4u35PBehz2C+fz50l6zBkCxkXc8EoIKTSWoEH3w1xzHN9GK1dpILea9mmKErLi
tD504+ijBBNyVJUlmG8lKzft3QCTNeCRNVJqdzmK2MUSY2U0W2aezaXvjdVwvdPE
c0U81CEyrAUUFoGbLpnuXuQUYBBT7iqsK148LnGTj9V/3cRH2ScK2lAgL/j9HRxQ
mIih4GsggJlaZMc7zpR4zvhA+R2WwJz1VBZpD0WSXf5+P0KeXqnW4F9lfJZcY2Gq
tmHIJrzwdMzvZKfQUjplc0/G2Wb6Oajcfdi34DmWBt8FZNQf3bHPGg9RzBp9OkcO
y32h/9ZWU+MggkXezrzmzkn17E81XWLDHDKzOvhAyH/+JBLUSjjm1P+a0DCyDPDP
xcAgq6khr8FZHoEp8UKabzJFciJ0gTMmgs2zUJTrOdKIeqSfJdGTjdsHXP8+HG3L
KHoviNW2oESrMfPBnD/GnjVQ7kFkNRmvuLpA0Fuhybqg7yfbRUt4TfV3V8ZEHqe0
a3wrQk4aCmeJAzopcyJbWVNHRUQOpdBCmQ8UFsVgbPYUB375omSxUqBKBnofDpf6
vkkmaV5iJCzJXcpfXizJnEc9cNwNW/RlFrVY9PXOQ2EKFDq9sWs4KiTg18rHVNmm
T1+2KgiZjnwHmDCVLBh1Dx6+UHclEkZQ+fb6L3pxQ1pPqJt/ay9cLrRtey+PrNOp
ofDvwRDbvZ6VM0unlzioKVmDa8gGad9wJaGfNVsmth3azr0MWymhtI7SbD+t7hA9
HIjVcuMDo/PwfBaJXGtPKYJLrUKFyK5e4R4WLu/RvM3A4xaIPCZljOrcloVI+r8C
nAKY92lDGLTR6+ynqL5sDcdoW1GEC5xRlvP6FRFUFdxgNUUyYyYVDwKjOQX3PT8k
6Yy0wtkBXqtcTbS3Qo4EreQxQd7oC0WgaquBoSxsV2VBopYpe1QEE2HbsbWNrO40
1s4HGDKss7UFYJrVVt4UCwxLnfl6Zh4lTeTDjQdOVd3vMEvOu7laJtNfB+7Gj1Lh
SzlMf4B4NnBsaa9XLF/zxCtHsAK8iGLH/jJN7iB04XfJ9zMXAgZ7lp8z/JMIdN5T
6fCR6vfvg5LG+nde2mTx2h0JJC5OxxRDsSnByN+2bEUF3w5JJ04z/jRWILGx7wnl
yhTQRWT3i6lWIzmngzWRkEwADW1p40LXcRGBMhMLl+g/PWL0uZFuOOPcp1mP6yqf
3K3HOnraqnbOuqO8kEwWRheVOnuwru/Q6EMhm6UMiJ9ofILM9hy+7HjBOlE2okTP
jzoDr5GB3YboilDG/R8gLoKFdHxwizZqsxrTrPuAr0eq7ma/8BryxmctJF3G/wBP
zOxCButtZWL1sRKrSpQb1JMpTH1SqQrb2e8fys4X3QqC7bFgxuW06jdZX0Xq+KOf
moCkieyNpphBDGIw05tFunyDstOZ9IbiC+0Ky/cTUzM6+dO32UB1+xxCmspQGNiN
YANTDtduixJKEQDCNQk3VG3G5bRX1wtic3Bq7ZROFh6r9G34UvdhzAmRcJgIsYVl
qqybsbkMPIetQljYADtYJeqFlmGmHpqFFG90k2zJvlDggkVPeO5nPOc/Ro7aJ+N3
URG6TEn2p/vv+dtnOtAMfCQCH6AqdCC8uSOnSmJfzIenLP4+mBbXw6Xa120RkHr7
SgROCo/KLKKY3mWPOuh9Z1Kdsvi3xwx1FwxXlwNi+0jD0hHP1IziUsnFUQ1eBxg8
gOsvPvPp4HJxqxrIhfX5FSSmblsnqLu284L6WPBlozpAFnwhQtDPMpg3hAYYwYYH
V5L/OhzqUwSGPJk9OIgBlkKO9r6OtIZuCVibodUKb8F4aAh64erKZJUeqv8ITHX1
+nQ20SsdwtDRRM88w/NukJuBcWW4TphOjT4cjyjx1T2tb2VbcPNkf5BgkCezYHty
9dTtjSGdr+GGL48XUASZaBzKx6xgaQZJ+km5kySyagW6b3P1/QmXcJIxMK4vnt5G
u/4YIuJTMb69jK3r3rY0Wpyywt6oJ5P63iourHlkw7IdzoNUJTMnuW2ChicgAWsP
dTtwX613X8f9iEE1tHOs0EXD8Y2e1xBS7p/dS1KnJbavPeEXOSY2ZI27TmfoIoBc
QBfmRuXIodPYzPTO8TOyZbzcpjJiOw1k1IHTKfvdF9tGhZa96oLm+VrdiwUDZlqi
lxUKG305AOaUpiGWPNms3F/L1spzrGwZMgkrojrRr9cAxqjcREhWCaQfQi8vsQFw
zHzYndfpAcmUo6g+3T1lRalQN+nFj8GnbgoIUv97ggkjX5T2owH3D26N3ZV7GHFC
gS92HuxNLyptgtR0pJWOOUXpOTVC5ho5Pcq1Nl54FX8h2cjm2C0ovTHDr/gkk2D4
nkKK7V4Q0cohcUnndoH7CtsXKilN8bmaKqU3cK/XbbPgtCUw5RN+Vb071BYOgOAo
5W8TtRxXWrIDmPlh0CmglxOnojLyoB4QC3LmhYZgd8WB2rpYmBi7yMZIiAmYQ7zC
MrNvL5g4lNoCvHU11TAKYA87+kONbP2pCsDdNsBbjBJnV23mJf904ZwlKweq95VK
KAFt8OMw73Sk+EpXPw+ptUTia+lyY8gZdaV6n+N/0FMfmspZiI/o0dEHxbwQg/ZI
cgrOiY67Bl886QRI4YWtLwPPS/IC41yIwOXVvNwMiKgLGoWp9sGKbsP80VjqBmsx
Udj5w26snK7iv7WQw//PuAx0sos29naquh2K+9uEkle0v3efB8DzzrdG5XgXKrnq
IfWIIgvlgQAnpcIccuypcdKoH7pueA7NCCWsHl71OSXgcVqP4EGJr/9fKaTwPnbO
jmeLY7v8xeB0T1x9VSu5RVDP57ywOFZroYavoqe1mp31WFWal4d05ZIwI6+ds4ak
m+nCNLN7uSNdc5GAD/9eS6bUoFPB/kDm379N6IRpA+Y+uXyPWqDaEhZuGKpiN/vh
b3rehTTxCYkDSF/QyuVUcWwJdrAKC944A3ybdpPkF6+/En5kiWZ1RTfXL5IlMP6K
Ybu/vCm4LGzom7xELNpe91YgaTENMUlyQgKzPDOMinW9Ads8cFr/ee69IReUbIAA
5Ql1qeiDGPdcsz3xjBn2Ajz26uZ7G27DssPQbYDX2ZgSqhJwkjOb9d6aK/AnXsdo
U5lRGAk5nOnMUMoadrltYnFMn95I4rTudRYd6DTPEYgui3NXBduOZ3iBfjPBK7E8
gcUAGMy0r5P+oh5HgLll29sk9koh0UwAtr+811FAx/YndUTA/U+AZG/zp85rsGtc
mAmEQEI0ZcjwUfhRw5VvaRlePSNzlXIZzSmQHhYVWuwsqFBBio6XCuzLF93gyQDF
P2EappHc2y1h0pMmhXkf9bmO7M9YvOBo1zmJNcyF7oStcSi0GkjK1yBjcLcqWD3B
nafaFo0tBhrAv5nkl80j7a0pvhjfanqWH3nqBDRpLbPE3B1rsLhNn6/XAI4Dl+8t
2r9T/nz60OsQzGMLH/oB/YG2O3bi8398a1gZFIFSpgB2XeZsUOM/GP0hMqXlczUq
mqUGbEizHM2tFgAXj6cgkoTElUKw60GF9SwDDLNZ+zmvHaMnRdyhgvzZE9/uMLbO
VYsG2p0UZeB9LXYxXPrP14pYcdW1Hf8j7aQGS1vjRZHz5ZWPm06cBppkL2QeHIRX
U8H0e8Vv4R4WsN2qwfI7dmkGnaCQ/CC9Da5ju1KRWzo2wtsaVAEWT2j4dIN8YluS
f+cejV7pDiBFjdAyHxe4BKWo+bAScgWlH8x1ImbOskJaPjgHwur3yhtmxrNJkYos
Bl0uzVBUJbjej6N459i1heHJQ45vE5ty/JTCqdmy1C/daJiVyWLbCU9/AM8f+jC3
tMqQBDHUN3/D3Tw8bPhbVI7ZT7ZttC3Zs9dlXNvNpSKYIXaat7GFzgwAuSgfzqGp
gECiUP6d+d4Vc12HzalVptgchzwBFXNVB2CyHRFOCWj59wzujnpLQkZIPd5cSRkJ
hrwqACZsWrRCN5FhLSUzLQ5R3cTlyL/8ar6JdHOlETnwJz7I3cdE/LXAfTHQu+qj
tBlZqrTLq07V3estf3aSa8rAm/x3X8lFSIcaAUnU6IYnKcGkIp1ekePSeNy5PFEr
CGQPrLH2cmFqhFiKZlLJTFJzV2ozY/9DowvVxj+RR4AxzRoOdwwTVdC4czlLz4wN
u6zkhgcoKZgqVh8rxWpWBESCt75dj1+wPXu+Ew0qNKmcEMFPrXns3AH/9VFoZIyZ
8zfLD9TSgzSXKekUpPkvZzPTIuGFnvoWEyL+8JC9CHhHfTvU66d3yIvDKrc9h+ww
Ib3oXt+XqJirfylAqPpLm/TH2hmLJJv+Bxyf93znVAUml4z1eAKvcAXwxZAu4Z9v
9oSbmMOgm/5GlJI3rgrFh0f86eiULzDbMtUbfoTWKa+rSs841XYkGSexGS2CMIN3
qSV65qxFCxSeDoxZV8yE68QL0SdwWh0hZVZx/nX490jh2fYGQRqHo0dNnUrZczU4
SmdhhhMqSksZ8ewk19NZU0I4wIZ6KUD+bQMX3VYbhSAjDUsPu0CNo7MkNIk5HxaO
hgjEQHUEAn4TbnAgOx7OFmcQVRe2if+hedcVXnnT5wQ6sp6inmd4KZiyV7wyTqbI
lp3BjZnSvcOJL+NKW4t/Q7a2aqlw1i8Or/Nc+BQ2qIZchGMIr+kV62VszK4jxcnm
FFr3FC9sDEH8uHo5B8kwgZv9HB9iEoSGCVqrItGAYds1D3wZ2giFFrIomf//HaMK
I/9vJx+80C9KEu2hPSfMuw0M3eY29GfuF3RWKscKLt9ED1vlOVPV9YPCopw+mlkL
bUOs4EGOLr22De1wSd37nHOsfGdoA89ozXQ8xa4NLIVCEq7rnkgfW4yVvmkxK5kh
d8prs67CnnZ0/ccW2Hb0tD+VrJapifgRV1r58B7aRwWFA8g7xezqWY2MRJifxQJj
Mtzgz4Kd6Pdx1/YQTHYB1HntsfpdniadMQnR4SbjKC1R9JbPYSleGxJATEOfoGfK
qlki3XNqfLw/2ANxIkTYa45b/HemBiA7lA0QLXxMUVPzM3XfmR8KLboD+ZYELaYz
8eSMZPEVBfy2z3tNVZWVMMVHYimoGpLETGBtbo25II+tbb2Z9Gj5Ppdz/tC6Yscf
Fxxw+Et1Ug1qEiqYAms5iKWTiGfEZh5gwyg9mPcarHWbIZn5RiFJYI/KBYRnjlOV
ZMdXJQPDJhIRBX34ZgOffsaQu89qFUhggeFytZvetwvlNmTpERakEvOvooiLMo3g
9OcAlPIUMKwxVaQDo1zNH0j/bBIRFS7UxOZkwD9lVRAk6mNCt9euhJa6c8C+c98u
HvpiSAuLVEWSt3xQE2+pbDS17Ef7sacMgoa5K2jSGZvKu9HheqI2w4Xh9SG62523
OEJ1B+QiPsREwaVwkeWIrBGbwznGSrTD9b/OY1X2TFrL407wmTIIcaUfjf6LKHue
JBdwyfdxG7c9TEnQPKoa0UyY3/NfGnvSp4PoeeAr7tfTqgILdDNkIW0eD67qWr8j
KDXdllCxlUz5zgxNTKv0DowKcJNYn/F0w6Tc6ku5yQfB1AyFa1iIeXyf7gt7J+LO
RIiG/EcZHWe0sUiZE9JnWf+r/ydndtl+qeLhgCppJO/l2Qy27OcCSR9b9/LHZuzo
N8dhoKsGxSDFs1vH8QhjeVk2jQLtnCPHwSMRit0YiOJJ03cNu5w04dfXAReg1xH9
VgXYWWblp9iLc4I/dhS8U66dw+OgxTO6z2YxlcL1INs1IMZlWrL11sOVX1aKVZOX
cnlp9swmYAe1m5pSEPTu5VuDHIvfUnuB2/jpy8K50z/aiyeMk4EHTMxKRxkmju56
vAQk3hw/fwgfOY0kzJNQAnclbp6os0yzuoMQXkbpz1vrnpytdO/Blr7QPPg30kC9
T6z34UAlYlzkwWyWhh4GX8K+82cRH1iz/+aCCYSZVhUQauNdMdo8Ltn4XYrpCuca
/FeE23x9P7vklgmDOn/vEwefjudbTUzC64c4Ubf4r/l87kRHYh3eEApNeW1+DpTo
eAJZJZja/IJfFA4jYLYXnRV+5WyvkTdga2vDOjH93BzoMmSNETfSlPToznXe3Ien
sJJoqWKDt+ijHP86mb6fBAdfAHKPiP9Ft1ArLL06q/evLATOUYXFbU/QCPTMG+rH
bFlL1xKlwdOPVszfrjzaTnGvw+p31eLrm8kPw0jagp7GCCrOtpvhEsF9n3Bap57m
NKXOPSFNJ9uPFCXPosdc6rXD41Zpy7EsMi2pOeentA5KDTHsCJaJlg0ByDu2NyPS
x/JMgQ5eKtOfYvBRdB7yX6qVhPR9QxAEV2F84JOrTKe73N2aVIAPUmjTD4YX1y0E
wHdKIS/gLSciJ9SLtFSgLeuOSL1ysIwKxZ/BXE/+A1ANGbfT/S+ZsUhO19g2xjAk
rKZPWYLa6gud+AZ98qX60CCMtZtFsjaCafElkzQA5uph2nH5ma+cLYKZPAajEF2B
ZXNfJGKXUQGfUYE0oraeBq81RL8Onjl0ErdqM9IwADUeG6zCEtTdMAkgAj/EtEFJ
o+kJ9RAAc198DS4tbKRAgG3eOHx/Tpwn21LmYa3PWnHJzNt5koWK+Q3Z/vyCzvzV
gpryQryVajOE/5iW3bL8hMWBrtxQh1zKDGiBqKTASNnhwSaMzGBaEykxYRrVFdYX
CH8y/1MSPAr0j167OcKOX873ZtWmRxwYlSNFdX4yXjL4WUw2tgaK33Md5A3lfwSQ
wxFcqJQSne18K3It0aJ6eY+dh4JAaA33ICupVusuknKUvWcDhTMeUOxBn2t0Dcnu
fTi7JZKXdzvTaQt15w/UtNkjoE1OI7Z4YUedr3V7L5UdtWsJswliVX7gskVB1Mid
hw1/t/79ED8pOOFWg3qU6xv3pUFXPRIboSSl0UmJ6mu7h4NLBXzTSPiqK67HvYfN
y/9lRpL4XmKrXxVEyxmH+KYsvjWAIwEPLeAlnNzlx2JNljjUGoDGJV4cmwUMyhdk
k0DgFoT1ozvTmnxgBzxuf+Vt9zE/J6at4pHWziR1pseVAmohytCH5EIo7auQPVjO
ISohzD9us/hMHeJ4sNqkz+kMRjvG3E5U4wJqILcWOIBsAVw5XmOLdeYaPUVnhgj2
G6meAwtXEU3925iI5Z1mrU3CONka3qPVGF2CvL6m/m/Zt/0zq3x4JpdjziC7SFLe
/25DKbiEQ3QMXa10fwQ7r5yo/MKOnNkrY/Arlh0rIERKqp3AIiRtw+u4wyHk1UU3
R+ZWbe+kimioVvUmiJ3OS0QimoLtgAygqkPCQAQakovMOfzFhbh15yQJ2yYJtKnv
RhPK5mwjDckyj6+kaqtkTKYfgY5i884UBooC0lQKLIjSrry7aq0HwJdOZiqKgPCn
9N0zMsJJcU5XU9kIfce/ruzn760lgD3dA2LcKoOOTEijxgSx8RRKfeGVuB7XUWct
/qGd5gqS4f51S/tnBS02ZlCZ+d+k7lrhE26YKoktGgP4bM2LESih1T7LRZkZk+W9
pga08QMF4GWQMbXSt8oD3ZjWe53CGhI7Zg3S8T5jtsQHTZ2sZj406t8ozEdTKGEV
/82I2geFsh1ShJPD3OJZdxDRo8ZY8pu9b2ausxHJbi3F4nNhZbY23xklMdRhtDqR
O7ZEk+13XyeManteYtVnYDwcLE8YiH4t9q7Xi9smDTMMa+j0X8jN0UsMA6/Io0V+
2GN2qYvYHduqIRSSSWR8jpvIDasZRgj/C6dEv2rKOqwiBzifQVj8rJ6FkHtArAsE
7o8qEB2kIXMaTQaXbyDhayae5tFma8KW4JqpUwTRDXTqvRH0Lhysmfjjcje9pfM4
K7KOe2brC+N3OHSzBPkjUVpYuD2Qnn+UTcHyHMidvH6oeFc6OTFhP5oWdZExH7lH
GDVZaxE6p5T9d/aHKI1/KNgcDzkDiOyVYykPqWfywCZwDKHLgoLbdlsqUqhuHJkT
yKb4jRlO2urA8JEEjXM0ER3c392hLOg35eErC3Ax0lDhgojKzZsFoDhai5jK4b8B
D4yMqu6CMrrkyQPsJun3ZAjHn5VGuvEza5A2yenA7zcxWm4D0f+vzrCW9gO+aGnF
tsMT2XjapxJiNKl6v4UwjpTplmVSMxU1pwG435ONV1uUgix0qP4ti82OlDVbiCPc
TsJevuOOv01h47KgS9Wu4cl82rM0sDHJlmZehokJgK+pyY9gJ36amr8JJhFDLesg
BM/DYsj4sWCKUd74Qwom6qRNyDWR/G37UGp0RTJSIYtlyN3MjKTp+i5cuJf0E8ug
Qp6Mfb4w3RMaNXTp/VO7gNWHhdouiy3CAMnbSi0hLr16qmtZAm1zot6eUzcqgXLF
kVLH5uYl/JjJZsFM3eAFafD4LCgnCNmP7JRcWeGdTYQsubHXAQWZeKVLl/DSl8be
XoPeItRyWZm8MDuun2U37M/HCH4ETKvXi9Fm1sPQS8Vi3BTJXFOJN/JSTyu+mAvM
OteSVw/a/5XjMOaN6WCf2PxJE0/KW0QbpEwqKiL7KwQd8/IN83S056gDnDIIq3d2
5XdB2eTWm42wz7DiHSeSc91CILK3KiF44VVmbCRcfoSVnJwmUiJdubpbXcaodVWi
gA4W/3iJzuUmEvB0AH3MNgmIWaQUomYZsZr7bl6+gC9g2U9v/OwI33OqUDx2KLfi
TWoOyyLqsX4qBznj+cm/Hu26J+AL0mE7F0LPDzMNvUTUxbFEJ5ZtWbACA+4oo+bp
u0UxFyoGyaKRHt3Maa2ywH/AJXSvtDlSTFrngZEb1/AKCcCOSvafzJ/E5iNx7sio
V/JSRRg1m5vbAgSmSMV6u+4A36D/2DEy/kAsCAIK6MhOjNH0V7va+dKSnv/B5orH
RxiwJou6qOVxUDZzXXVUjzIq5dZ+e3teBeDUhuXmQrzTcaaKiGawhqJafVaOcHpd
nOkSZtZoouH6QW2z3puJMKDs78MTwdSa1ybhIjfeYKjZHbs9jLigF3fT6pnQILuU
5OMvoSJ5cWqsOiGgRi8fdqTeqkAuckRGGVVcbP4Twl6yj0NUEPaPUITAaOmdQ+Do
ui5yNyh5yWMmihIw7DsFfvW3wOIypKU+SB/q9qc8U6FXGXiTHs4TpYJlvw8z/jaZ
4QvtydqJsR9AzO/iPxnbiv3/ZKRaXC7cnXAf0HrbWAw65HmyJyUD/BSetOKIkS+P
pxmHWDXuOYRlWS0N0trlEE0YivvB9gHf/LGzErZlu13S8pBjWhn5jXyquK/P+mff
AuDFXw6IH0fzafpag4N6tiPe65i4N5C/eSoWu1xKpJi5Xn/UaDOJ99imOy2lYupJ
irRv47nhJtPdx6IP6T06ioc9VqKlncASBCcXcF7XiQYMhQr0qvfrJKFskBb9lSHR
MNcia3+azrsp5ThsbZui2tl2RRm++9YFxOAMWBhUdhISTS3ZxClmH8VSIt3mqmsU
c1GxXasxGepSxxOpUI2i2LesWIiG4EPcZ+SoSsnrIuwCGKzFeDStbfB3fnfil90k
bTuyOD+REUVCZQxhOvYRCUNyVf2cq0ik5NvXSfLlNfisafJ0X6clkEdkNoxEPVJb
ws0cXJwf09R0oOELEB8tED+EK/znjIxYrBqXynYr3W3jtdw0Xn5bCzH3V9C6Oc1l
oTEH+k0N7wCcH6c87AAFHGgnAxL9vKCmcd+W0x1VU6+eXuAcayIj+0AKawCS7yyL
4xx7lGpFbfxs81AybYNww3q/Anbr1mQ0GAEmfGzhnXCTCYbmqwSzFUZcGl4XCM+Q
nHq0T13CYT/qlew4lbZD2YGmpjDMHkjG431W7pvs7aXPTtqvhZfzzfYeRrB5iyxo
CE52c8I6+AdFrexKQjQ/BrxB/zHkdthWrqvzBwHgbT6l8Gn0VkNmWthd+n5tUMBk
tqVfH0M2CCZzLuf3MwkohduUtUFLliBMMm0jSsvCRJ7gjjw0DMYdJkE+BJfDXb4M
NV0wXW1ZbxISMNhpDcpkbfkHYr1apmPWiPFkV55sdE3nn3ys4e95/AHzdNUK0J6n
JVlEpDloXtoACC0KkXjujhZBaKN6K9fq9AI6RKjXwquREDETEnRxs9ZzhCgv+tY+
z6hFFSVKwJ4tldmU6eqnHFEB+pL7EX1hxP7sIZUsKvCfTpW1aSqRx4vwrJW+BxV8
UqCWyHiNiGpj22FT9pAGGOFKqKeFIiSs0hZP8CcYBbJFpesF1Cymgosb3+DWaKFX
cgkzYXpgtU2HooFIPMPjY1JwwwS5r6XVroQCqGl5XaJv0/BPlkt7gYFmoDBF9upM
5OdwD1cC8e2fa33igSQ0KMZ44+MbFNbwKMcnVL2tOwB7Iq9gWQPHDfoLrVu99QAH
+C8C/NeMouV5KZ4TL3XqwOB84IjQ630B9fb711dG/5zuCBgEK8DKhh5yt+69nNfN
dq/IzZpZsWIrDgOziyHrP9iti7W37TyFH+Ub3pnFBuvJ9bhV53Jn804JOMIPF5Id
GC8jvlNe/82vIyksn5s3fxmSnkxmfH7X/wx4ODmn2+qHmpDMsSOZ6DGqvFz9eIff
8XK8gcXk+FsVeMbbH3u9/DJMdJsSFnTEtqyfTmRnuM6IGRPopYgaUJl+vk0pYCoI
KlFfWq/geY2D/ZtHoUDWzjClmyfz53ERnsOa/7ZDgemMYAL1Q1cTc1jdQw2pYnL+
2UxncBjbBjeoEAEf+kJ0I5lpasUIVxodnCf7Z8oxFO4zS+TNGRS5fZohPYW40XXu
YljRsPdd/ihhwv4j3W3KDWoEhDlgz3wVAwPUIqqVvtCp8aXnKu6texQPTUUOS+E3
rX89bftn3CQg+NBvkEC/VWHeE1xYKPxpLdBCXo1DQemej/IeReyPzirGDFBmyAEP
ro/dYrltIZVYzVEImFcMMgKrswT3fUbShiX+P31ee2mUaMOOE1OIYZeNAJsZ54PY
R8Mfy4UH432d2LgpNGBrKerrU+6kgTTlLcbGMmsyIyHigv/9Xf1lioNyXN7V+T8I
NlB8dLcmBuJ7Vz33ABiX+Akf7bw4qDNKiv0Tni/hd4QTNZZ/1l58INOaemTNOSi/
2l0iyvEs1KoG+3EtZIrseetVtS5LarCMAOzml3g6tEEGGVxeBbAuQ4rycwMJBWyG
2NEyHuyHVbhx+0uHfAQx8wzcHLIbOAAvh1y03IA1XdiePBAjJNoAhPxvjUGq4vie
pqCCpVeE+F8T18ooS/EQEZ28cbllACIe3Gd4o+qDG2tvV2O0mEUQwza/e/ZS+ETo
XazHuueB1M7WVl/B6c0z3u6gDIH5BXMxVz7ir3b6Zoy4CWmyMgujqLxUF1IqKzLc
36j38TX7UrTz8ne8VB3ssE1tFTahx9wgIgi+5zYe5Ri+4E6MHzj5Y+F11mZM1yxy
dPjmiLKFM0MOOiSrhS75u0SXN3gE09wM8P0YgoGq3/dRGR5OV35VWVP3SKmePMXv
R5E1khaVNO5XJ7OnzjFYabMVbaBaTVjAzDP2jbbyd4CrUxM159K3KrLmiHbeI8X0
DEdyJLFM6G2HfZ3RX022vHf6ImGVUBsMVrwd38JoKCTxbvPLLZy+RkvhJpLsuhjH
MMRDf/VyHzNrYtcfTbg6YSQD8vNIdM3plLw7kPO4mCnl85CKYUPxYEwB1EKSc0WN
YmG7AQ8BWKZ5KZoSwlY7z2s8Iz1zNfQMZJZ5lv3Boc77Xa2zM/MJN4oVJd9MMJ7H
AoNZNbW0l47VP+LXnmzYXzc6GN9szAMzBI0ZaiKu02BwhktiHD9FuI8VplERWf+6
1ztjB/FeVQzL5WrnpUtCaT7KCNZg3mh1jBIQBe+BP/v/hWZLSLlFiKXZGxM05IfT
vjVWWmoVzveeh7Zcg0pNkq9xMZh2sgExP0hdx5PFjgaHWUkc/A7+jE2ZS66kfYGM
XxnDR6G8iEP2J8jiGUF0QzsAk32xvtrBUjMPdDxBGmwEL5AKxObkyyDbuRFWKrFa
mwJddqpKPgQ/rKT92qd2CVYJRkGRR7LeYfl7yfYpiHpBYnth8tjEOsBcE8zj71lC
C39c3Ja4qYflpHNfI1yPvL4CwCAk8rQm2tCARVNsfS3nv+4UEc/lgs7z3hHXNszj
XNAb8VWGR/Il6vqTJBSn5O39KmYiExWyIkZk4J738glyXyC2qLgwoiuRrQ5IYzfI
ywIE5RiS5hLFccKJwU1Q61ZfAz3+V69PzDSQFDaKt8Iuv6qGTpfGW1GmiQx2DG2f
kD4ywkYn5ZjMM7R7GkUodac7CPVL4gdNvisnUkM0DQ1YPjdsrN+7FCNidA6YZQUK
41J3ywA15RwX3W5xZ/McPuI5aZFLX7K2/sTlvZROhRGdSNUTxTcyYDVpsxcaS6LW
kQqpQc0I8vUMZc1kXKDgf7iLh+vj2hk5OrYRBx2jyo9XJMdzvs1/jMe4cOb3o/vv
LGoUqBWFxhcW7FS3yWQ/4A==
`protect END_PROTECTED
