`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Y3mHfYgQ597nKVxbkJMv5+gdkw8ks+WpNzowTGbIvPfKHh28fd9ePkf+TgTJLTx
jbfjnD1pR7WJIBchqraOgl7Y424byiFI+U62zFWY1dQIZOua4j8hQITnG1tMvlHp
RJTWjgJs59AyYQXK7kv3MJ7y1kRBJV/Dv8ogUEzpavWpBEPov5AjiXUk1dwYt0Yu
bZp+7n+LcgNUYhX+g9KqRX6BvFSo39tnak2Yamqb0wRe2mJkfvK9nD9Ym53i8Z6H
M5Uk/55NSuEQHQnv9ou3SPaKjOh7ICm/0PNKM3cuw6WHfD4NHwJGHUTo8iJgMYrl
rcSFRjTtNeMVsElgITbbudcTSRuHGq2cXfkpXgBrRdh/G9l3Xsjw/WpWv6RjTQ2p
+Z5PhIH60cs+Jrsao0sRqyI2IhnGOqNjjVLhwleoycnPfodontQpEN5emwiyA6ky
l2IHg1Zn0I3wdy6YzMQAqVcdrS4xqEhZfg3MsEWlzOs75idHzEulVuBBh/pBbpgn
ZuN5lwucRMGjkvL7AkNWCkMJMsqKBvI+kjMYrc6FZdXTtshnO8m36KCUK2+CG4nX
Tvz9ZILpk/kLCMsGv52ZnNh4a89M/MOkurKwayfyaBV9fvXfovhMoQXZFRzElaGp
o2cPMAlK6VqFoHczVcw72H++aU1VKBab9qUEYtejDnCgTdUpVSgM1dcq6J8Qq+cq
RhVAGJRZSlI7MWOVgeJ/BPedTQX1X//5xROndRthuYvakziTdBpx4uGpbLXJXs8x
vLPZUiu0ZRhoEyBAsxDYsIrJ8p03q5BDunt8S9Ffoi5Tev3BT5xhpvguY8U2n5wy
Dn06odO0jq4N6cd+Z6zQvzmvpzoAfRBJfumeTWGuKE5BYzkpO75VN+nv+ySfrwlk
DxVE1+tOSh8ly8fIKqkzu6v5ymAZzfj74ARjTzOdxSQEcO7BGCCXTgHFgJnmfqaC
lP9g5Lbocscddyyqu4by32q2VgpbX/gddXjrX2T+/luC3N3D4ElFq8il1uz01ayT
DcpgnS3JeWfHFOomJ7Mo2A==
`protect END_PROTECTED
