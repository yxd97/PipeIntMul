`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NSKFmG+7nRrnKnEYkjxeSeD5DegaD93NFpV99HQhxg15M/Dzdvd7MGQWdEBit8Ih
Nae2SHuZ72gFSTV9ldggoeONe8ZxfvXgMHVmfpZI2TCrRSmGmx8WVun8L+1ioY2D
oH81M7wzG7l4RTBx+UvLv9cV7XuPgh0C4CDHM6uzpvv8yiv0tjXsT+nd91oGTy83
/LZwDkWRcKCKKOlEQlZDd0xoSeoTgXY+EImE+BLjI8rc7A04zBmpd9IRZErPUyrX
8wdBSBnMqRReq/qbwCT89zqcTf7Q2rrbpfi3KmXJMfexJfPVvKJzGK1bU+27THIC
NPZhfPzsbnhL03G2rqiXoM4gZVOS0WY1NwPerhI2JDwDalVs0CWZ4OZ5VRJNo5f3
SGMz1Qs6DF6WQcDPxO9wWRlSDwFBSEn+EWVaTOlHTVmlxYZ12F7R96bZCCTQ9vi+
`protect END_PROTECTED
