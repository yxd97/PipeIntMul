`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pkFNPigdr4exuv24GbhlZXPEFy2Jz7BH246VkxXntMqD6bKhk5KUbIpr5l74DJDN
k88Kb2/Vnq7GDHhlIYxmCV9RPE5dUwxAX9F6jj8Uv5miROqnUeQvGFzNZH/fG7AK
vfE2h8+fHp3ZhC4XOPainN5VObj3X4piJ6pj5y0p0/iKnFQjQ9GgK0AcH2EFeMxd
Oe0OHEyvXXflT7VkDzsC3YyfW2nq983+9O67489U6M2yJzn+TNrp9fGZ0me/Cjd5
VhkAJm6tSsUzsea+9NWKfdNAtLzmZaXLyFsX+TI4E54Bid5IuAZdmHs65kfFvz8K
dEAPIwkDOTVFctCRAIjp5HsiCyBZLT0c9e5FAtgBVuvAUWillGf1euGPSNkDwad8
+inxf0ek/72iOjtm4gXSzP47F4MhldZDekog1MAUWDxkTg482hUBubYoPvXUHacM
VOTScwubFXH/2/T+avmCuXd2zjC/3A/cX/M1K8TXAgpJbLVQU7h8H0LTxPB8AvbT
8rcrzN0yil+aQ7EoHL6k3fPuYyDnRTqkVUsIwGMh6rL+6QW2s4kwJirnYUyJkJlR
9bIV1uGQLzxWWcpc3je3p7ww7TPzME9Etsk6UOurmnY=
`protect END_PROTECTED
