`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
169CZWVWcWuDaxnAwG8sZETpRFxRUio1PMFl9lt7nBzsa7dcrib2okZitev9Wv8J
Y23T1uB9oXsN4YH3eWzURtj9KCMl7LsQ9aMGykV1Yu6pf0P6WeuSwlsuTOuTCx8n
kUW8fL5lNUhks3cOilq/w/sWERn6ftJdP2BNoIohSjQZQ7w2b+AnM7b66X99G04p
3vHfiskUCif9DDTjksRkQZanp0y2kYtGHQZJ+4cXziHN7Xq8HANjYl3rjZU1IsM3
o7rKNdFmRxjtFzLLpfl6rv1PMG+XoxuYV9xl+2NeP9O4eUYAmcYzpa1+KClidGps
HO/3RppuEL5B7CifdMoRyGL3HdQ9K3F6FaqIyV+G+cKYbut4xa0Iyr7cRgK5EkIW
G8pzlCCThYmsl+vjecS+cEKZ5Hz5BVh4Rg1L/FWr1JHk841V5dN7JVczyWpoggTM
xpVjnjF5gy3rBDdvtlOr+QtMpNKk2amQKUKDIWQ1evWZWea6RP2tPMgHi8dGagdk
sbH8FtZY/pa+WOKOEGs9xyzrTUuQaCQFMlR25ag7Jd5BiiCyosVemOgsNQw9hDnZ
9AGo5JdYZxGUXe50GFDsCQjFgla7FhUuI5bJVf9N7Rf3tjabNV9dVVtU3cwInQFS
svDUZlWmYQTkVZj3Fo/XO0ReL43MlWvtnSlarNgz9d9bqTvfuwIu3Zbi2JN+Dmbj
tF16iXV/z5fVfhULkFhWFQ==
`protect END_PROTECTED
