`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7kFPbbP4nWscgOPc2mJBYYltzVhL/enHMNp9nlYmZlGGmn7fnq0ecq5212rlOW3k
p/VgELFx4P5zruoyrTXtw0/ZGlOdFsPqF8F6QL4UWVfTqcmqMMr0i3tA64tw/22U
I/ph0FR/sJJShHxb9SBtsfGr0bxJsStgBXxUmkHjA/siX31cV8PwybGif2yRi0KX
PHX13omLgtGmuM49zkyFbeVN7LpbX2LKNguZBQHL1EEC3OFz5gWUsG1JZkWZAx4R
Jd/b0Amg9w7TvDtDyxIVHrfl8cvr+gUl1oi9S+raGL8ICTSHA5iOPyaBfGuVuMqB
gQjjVICRGoE3QZ7+8B7vtojm2oyNL8Yy0lVdz82bWZXXUfeTXC+QpHh6Ctcy6oIh
bL4zGk8uF0V0RnU4dlAnzcZjSpKXPuOKH2cO1X7hCRed336tSrLVwQH3SWK9UrBW
BCdy8Bdnt3t/HPrlI6VeJF3DY3QP6yl0SoIukb3AZnOEm40e93HiGF2zNEC9EnwL
6bwJFDJmyxkiTc9skya8Ie1u6f5bET30G/sTWGQZW0LgIJ0dPr9CbujV4+tvW9Q1
Z6mMgQ+jnHxcM1PjAeeEQRpR2buGvYkMG/sPW7dJhQo/jFwstmQaMcPxZ9YYaltO
X8MYtIzjysg/qH1hTVozgw==
`protect END_PROTECTED
