`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MX5iFIE7MMPlRG7JZpi52K4ndJzrfgsULEJmbgh4jp7jfzRtS1PPxzk8jX2Vzh3c
fPmglMSux0lowDt0DpLEMGZWGLtq01sw1ZnHC2UxLGhO2kl6BdW0b+pAPlZXAtG/
jdlDtV+7fVnRlXtadtZWevgkG4KUAvrjY4oHKLRsCu0KAtfqaszk2FR3rDrWbzmB
QvqmHCr4vufwHNbc8SbeXeRWjx32TiRSCv7MQZ0YIssYNrO/5DcIQAewxXmn6wMG
jHecw8kMP7nq2Oj2L934maVnxMDGm29wR8gi4T99AYcxqPmGwWpuZ+/T75Yj4sVR
sCVUdN0dhehbuhfXDA9WDMBBr8qnqTi0tMYSoCdo2KlxK23znU88VTkdiL1zyK03
kPpewiF+nDk6D7/rEnmOFbX9bM7FGlO7FLC+ain9JaljIFUnxP+S4zLgrrS3eEh3
TY621hW/kO6504XBQpl5DK2FYv4iUxmOURsWHYWbmcsOamgZJkNg2s/sn7UDxRXw
+Yyi2jnsdO9mlwDZEw/b89veKT6rMBG4u7qC7HT777i1svlze7Rn1ywsGyyPLW8D
HxWCJN1TSskOKv9e/ZHU8mDlIjPxBkW0SsDym0yykmZH1lJhb2rvD3Gm4GAX5Iq6
0LTJUKdaEeCoYkJ1H9OZW4CR/U4Un3sN+UsgPTXzxEh6EoDEYk9iU01TIIfWQaML
Eemarg71I2uUr2DtPCOzUO8OEJf2OlvrysosGWohkI2U0uNCPS72klAC4+wGloXz
g0SNngISckyhzvVwwPc0EtsiADLVZym59rt9B6pUxCFPQ0u6jfSVvujk6zupIEMs
+8zSdy6/6Hrh0Yvbsp+hRI4pdAsMfPTwjn+zfyO+7TdtxQJaPg3bnS8eEgqHDKss
GjTvZ8OPFULbKNAjwRiLwXqf4sTSbAMRuQPyJWIgdoSmQjP32wOM/rgCoQkU9sJr
CMzHqOnLvVnJVGFOL7zC59850hsqmOGsECzf+HWg+dYclJQ+SReT5bdqXqi1yR3+
bKRBnVbTsp/xVO8ruU3rL2jCVPGQQQiX9yxSgo0TDRnSiwCnGAIbAqimNRe9t1/B
Ro8K7QF1SApFg8DMHO1LzRSisOFg6gpPQqjfKx6yNLLrZ/KFF+9ntTd0up+VMMxQ
fT206Oo1/YPrQBKAdP26PSoO4N3Zv+TGIZAF6B9z3/zL9qiJ+gGZxKRLm2GQyBKJ
`protect END_PROTECTED
