`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPoCi47abDV1RlUp9M45eNVzc4VyCJGZuDWi0ce9hHX7F9gNDHvgtEwV6T+1Zsvi
Y1cYF8b1fVqbS2qinKyloP+5G0z6BK/qr7rAkCg2GkezKklh1gLjY1UUw8Ia8G47
4vXrWZ9uQfRKIBSqsUOyydx67WWXfPvBOKwKnidTkOhFdSWXsmW7pdNw/ZLbcFdt
rRBm9kpqINcclLila1cVYSY42gZwH4UwTZZ8jLe5aJURXHBFliQ8bDDhs7dxgPXn
DqEwRHMkdHWnLaKUtnBeAx8J6NdgUI6DAi0r1XTgvfqMqE9lILz3ry4PhsdUg4VQ
hpkjnSIfn6W82UUIpt7DGAepMZ0vjeggbFXNN6RW96QwxmzCHONz+Z6F70SMJSFX
52WrXq84jPyNqy10wU8tKHa0z0efJVzDFp0X2+WRms8=
`protect END_PROTECTED
