`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pz6tuNv0i84FU4ZT0v7QHmgs4pYnPMWGuXUMQ+GKtXjy/ukun/TgMZ6wKG1rVYLS
nXqM9J3Vw8B56xx/zzS5qY6BnOrQadDSdslcU8urkKM3mIDHlaL09Gf5vb1ygbVH
A5Uby34HpWJ3EC8DwX5kw3OWzEnC541GQZGaUNPCz3kjJVGJnTYRYyqomfqFbD3q
NUmgK5NMl9sBk5gm3vvkyQ5E0wpdVyiAVnVTOlcwX2OwYxE1ftp6cgdhZrvGaZZL
eyejlrW16RzZ2bEKcWRSipk8uCdN15AthPw/l1nSxcAWCg4KpbtdYiXloT269AIK
DIDzToW2zssELnyeTovp1oqJ0LldSNS/1XaridTyH4+ooq8iI+SGm7ILKU67opWJ
ZsK/A1SSbvoBzCd8DDNXwAOLtYbPaxPxRkkMXL7JZnq9N3U728ZZz9zsRT2YhrJq
S0DQxATY1dy8ynU4t1zSbRDLwQ6Pn03bCksjBEGr+rKpD6kDHqRKLm/ttA/ZRGD0
`protect END_PROTECTED
