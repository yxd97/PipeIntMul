`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0B/CjvGbUWDQTLJyv4mggmeTpo3P5IS9TLft2FOp8W6QG5I7uJpzvYVd8Z147cH
WiT6oa69BrChaslNKEkLHXhQVu6yhrPJzv3G1q7LVWcKTJW/u+nflKHyuuqqg9sS
zy5qQe4nJTenK81xFN1laUn2+cp7xCXkJylNklP0YFzQCRH4R0ME+4LzfZ81fVgq
hfn20v7aPixwR8cForCVVOtt5ygMYaxAZZeEL7bIvGPoxajIHGrtlSjiohz5hRfm
xruRjcPyliUtrakRB3np1BNUfebuyO4oUl9wsN7ICOMGd2O79mn/hUIwk4Ms5F57
RC5yjMduNY/Jrjum5popW/fxAgbNCVdtbIfUJ2R60kRCJOsR9wv6Usbxry9sVL+h
c9mUJx2J12YsujagoRqBkhdgaD/8v+WBXwiL2S3vXf6eKDED8vlTGnrPHU6vu7UM
+63xCCjZCbLxLmJLUIGvnpAiNT5JGE9hlDMYEWwZcgs=
`protect END_PROTECTED
