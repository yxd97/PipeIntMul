`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RaLKZUmbPgKvyQzbFKm1SSNzvKj3i4zCWANcyMJJ4gQYmnVaFWgtDN4pIgDDfbS
Lko81ST7KyCVmTtX86I0TeXeDEuYqq26Ip800C7VXUMR4I4+h7DaNPrYXPopf7qe
+uhLYjUNqf2b22ltVZoO+vjJ3wumYprVi7ob86HCfVbt8VxyqcWRskAsc+usUGvQ
nmlhU/Mz69yeSDaMf41Pg9HIJtXFB7i4u1guL9QYMk9TnV9dPD1PkBmJI7vorf1w
qK8E+xbhAG6Os/JPaPthuxzlnly6rZEFUD8/Qtzgz4MVwPLNAOonX2Fi6irgIOeJ
VhqaDYamllWBmaByLkBN38Heyly9z022uEXkK9DNQZTouqtGO183pJSHAwd8mhAG
WLDc7pEwbF6ljJzkGnh4Ps2Fudza3zLfOupx2J8GRTPxk2mPQzNauxiPMPFtCD8h
ooMADM8NNjrXMFFbRHEDJ/cRaV60FpicdX3TVjQlzAqBwKrFUJ0gdqAn5YRgG5JW
ILOpFodNpiGz+G3bhVUZYn7k7hRpwtJUV/esNchqXg/ujRI+WK+Jmz5u0CnYBbFQ
HUc6hcze4Y08K5vVmMvLIdHeXolB8Y+08e/NlKBf+pHBa++3UVILd2FMWIRtYpax
6J9/Qs5QO3fOlwQtGXB59rpArOUG8F6lfjq/kmLJ1k3t9JS5xZy7gO4orFMJ2Cjn
RHJmlqUAnl5U8oB8chwUcTfvW5A1S7cx/qSZaB7DE6fbuDwO2Oma7CBYiCFGguEf
oIFOiLke07ajdKSSMYz4RNHXbrdkpI7hl9p3TU1TlK5T/S/wQg4WY43MuHf0uA8l
+Dx4h0dD7Pyd+RXF5WF9c4BcoEp+T0EsjEsFhZ0cSnpVLmAHMs5HkYoEd3vypRsl
yNPCy8q2ykjM3/PajwftsDdD05rtztKtQ3YnsNkI1apSWHPKp6GHMI7iSNDJvqnL
6U7Kuva9v2mIwuYxG/4O0i9+SIx7WnVIGCLmdjrEqtU=
`protect END_PROTECTED
