`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4mPXDiZ4rb0PuxFgWMdZP423aWj+nESWMuFH+BtGMU0zh+rZblLhYIYPqCIu0uv
ISzSVrw/emqDsCMfvFL9qMpO/KCjUunADIhCwHMIIYPr4FEvq7G4GxZ6JRndyoQw
cSxo4wiw1WOhSMA9g6s32eyCYTLAb+ZT+m9iEbb5DoDYiBvoKr2tKXKYslJGVibJ
lQDS5QaYuq4D/rDtrYsab7ylDUp49qXJsriUzsEHXCStKgvYHLQUPyNV8h4bAR7s
+rJjRXb9pcSN5AW0JyE3QV6A0azlpIC4C/Gv2/QKx81toCjapH8BS2kZYuuIUW7F
Ee9oVnnYSaCSJOAj7GtNNYaOMtL8WjhfqKhGkj9oQafb0o1XF8IdW6Bbgyd3la+P
X6QtRfm1gQqYmDQmykibrDNU36SOWfkAT2IJrVmc5IASEfDMWZNO3t491DSdKuw9
`protect END_PROTECTED
