`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UszUKBGedC7QLw4D4ySXPp2hiTQXMPX8X+tRRUUE8o92Ujkx5E5PW4U9pkWa8Jbf
0vxRWDR8EQHm7X6E8Hs2pvzCnqZGWr6ljUmE15HaTKmZ7sfFybbe3G+rjjRe+P8J
fubl3Hke548TR/o058fymzZbxPxZhhBsnWJoxWt78xxRxr0X9xH6RNvKmIOWykBg
NirH8Yq9TCyl0hHZGVC5cznZRdVzxvWC1i0fuzIFeiF1DbjkVcp8BMqAq8SEe4wi
7awXtdQ79yX5m8bHM0TSp+KQ0Yo2H7phZdZ/rfoLhnaEO6b0xiKuE0RUiPITbz/m
sLkz6GDEAUsHgXF4wlIXxpBck8HqhszPmv9JHoRs8XJYKs03YQUa3HhWmHV6t5ey
5uEiHUQijLrJk/aaKfEuDS7SEgmykHdpl07QZuAvJkEWoj402MtSMjqwCXbjwc1f
w7OHtAWgtpssIlROeXX8E7yVPPQRdUjYysY4hkvGRsws7oRza3V1IGx0mZoUCFCM
AiTtmcIfNMMJMmrx72gOEYEpJ0ay/Gmff7Ho/oIGA9pFydYv0yQyoCdIQkReMTPt
stTJmX+sj7jyfoYsWQbg3RmBi80kRBZvDmioBC0SrRUro2beZNhH97NtwVXdVanD
TAr4C/HCdKjgeVd14jWkyw==
`protect END_PROTECTED
