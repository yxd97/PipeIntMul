`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PASdEaCdcefH0Z0Epe74/du2X581RC7h4TMUl4wejJVPlz8sopRgIYI3bQdaG68
8y3ia0jqW86cU5FqQ32fFRK7ayWtul6dwEMdqAe7hQiu1l8MER16S9VMit3e/K4O
8sLOvP6zzhDh+GNuG9nimZFQjADb68RIO0PC4oyLhiGOW20B3FLM5Ben4j8h8jjo
idgwZZxbaqFXNoCTRAfInEZnCxQNBiU+aw+Q/pgPLzIWWMCiQZJzeySiiFDAHhUm
PiWrf4LmrqfoxdL90PV42qn+5T44r247l2KoYSG9f8rXngybqIHprHEVfFKb0j6u
3gzcRotGIwWE3Z3Rky5gMxPDSSpHSUAEZRg3F1ZzMkeNcg6GgUKg0oMpOJV9SDDX
rriaw2GrCfuvg+7uAgG/fUIPFOruTEN9hDu26o4wTdBZRyADtIC4T4lV3FMvkIaG
U3lbLaKgNdA6k7MJkruWmAiMpA1zcVRSwb6IJBio5ww=
`protect END_PROTECTED
