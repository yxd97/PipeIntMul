`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NiE77Im4mnHfIPMepqtBm7i+GyGXzLbi54YachUajPCmrrAwWEO1hxQyrqWaOtj2
nXr56uvEec0i8fYm3sPUHxUzlN6pcAS3iy38OZMr02iEgMk3bZr2Cs8nca0xzYTF
IfOn9vVpROIyE9RBdko8YVT6UPT/meHGXQ19eem7vIl6BkJfc2zb5KT9Z14lSmIc
m1VHSAxw7zrzjxuoMvk5JVcvesgUyFVsmg+vrvn4OpsPHpgoJJ7miGWTZWnS3lg2
N9OdWQJVGuDtCmlHl3SQo71YZC19hy3SjCHL8OdZiYJm+b86c7JZTnRSyCPEYZTv
PbNUFXdk4+01kCTr1XNaSHrnXV3ufX99iTeDwrckSXw=
`protect END_PROTECTED
