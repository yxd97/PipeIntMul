`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oe2UPsF/QVa6w1l3GJEyMxJe6ilkfUuBaC28wsbZRPf7kjSwXR50xRw0yqDbtSt+
rtwu7bEmvQ60yi3fMvSePQfuQW9fBZIQj5Onsu1RxHmRWRzcSTAJmqA0vp/Jgj8S
x5I0OqeD+OaaSSJWfA14mS3KoK2RqzH5LzxsoHwlp7DinhsAR7Pwu18dxrZh6NaQ
3BtwaD4DHqFNGlNw9Pcecc1irxq1v2eTa8WiLnLQxSJl6ZRNtpVsD80JnXri8Rwl
HKp6mXRR+y7Qs0wDwhGmbT2ZS+LmpAy22XUzBQWx/FXjZLJEKBZtwh/mfD4Ftsj0
11Y7t10l4RWS9wSlyNgqnUVWHK/SbM6gl4CKrS71cQh2ciHjQC3zKu1OKL7z1aDs
qm5gVF4BgKhGbTjzkfHw9CfmIob5lSMN89MGAXvXecqldPFeO+wxmWNZ5XYCyIpG
vyqN1e5VpA5GH4foDleZ+Omuslhtb2O1fPciM0KoRewsUQ/c61AxEpMXti7+D4go
nLvesIvllydtstldz7at7ps2R66wq/Uo9Sa52sTE0QrmMqSvxQXz67uN5WDd24La
Rx9YT5KbNfX0FoJh/k1dCO1ZyVGR6M0cUJT5uyHqY60bzz75ZgwozGwkKc5BvYiK
2EhsyFP6Awo40ahO/gJilscdd6GPDFiDAyb8EVlxR7ftYs4X3bCbJ+hIundxAznE
W7S//N9uVbZdFskVv0nKTAnTj7YLfJ18lDDAWyvXdNm9mNdkLXYbUTe/fQFzInbx
EB818IoH1hexaE11E1pMT5CzFKpEtZ4UTXeQkx650kHPZRl7stl2yQbo2G1VEnog
APkVz2+PsF+R1mf8JT8gFiVd7l0EaevMEazDsunqZf91B9sj+myRG7uzauNs27ZB
2fZ1QMeTdlt2TzSOV3VgGTVS2MCTTaZB3TyekownN5SWja4HvOGBPlT9MQhsXneC
74fQ3teEgO8igr7ztOzk88ZJc+C26LDlu3V+FyCyIBAcGXtODJKu0u8zDB/zxojB
yWTyDXG4gB4yOYgjF7Su1iuFaQgxXNu6bkG5orMMjJwRj35JJQAnIKwf9Q3gPEz+
9WJ4Fg6yp4+K7sKdu21JhJxmbtGEFla0nk8MhAFwHm3M9Ug9fMGe4dfYETbBuNij
5My7986thiZ6VpW7ftLgmU+Jp3GzTg4L2HRwiJmRGoZnkC7j8wdltkwBWYmdaNWA
8R5J21n4qubW6zh0Mynv9TMyTApbVYUUp9My6Wpj7hpr6pSzabZdKVmFGYdN1PNk
pVMIkeuszGiwARqCHkmU7k+YVXLOLGnWUR09pTFEzO3RCqYySa9KdMvZbHThZE7W
`protect END_PROTECTED
