`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BYRv0pqJMN8/1DU0d9S04xKW2v3v7x/iFfXpn7Yf7SMCStJddWeEA95BQlozpEy2
NXlzqzip0eRWrkkRjlX9YLngxSE5dE6SkZNVFserYEfm4rWEYucn9wbLdCaKWvA2
NaNK5p7dX+FBdH+9nsGldtHN8XnyLEo/eu0jvFVESkLalAqkJtNlxWHy9B2OwPT7
3lOFX+SIXaQVRm6GoQOSxGqSrX6dps7VT8nPMDNAkpHoacQ/uoxz6xb4lJzHwPeU
86tkJd6YFxXK6kD3UMDg+C4DUGIb+VS4uL11O9o3pL58JO/bW1jk3lmJb7iiMET1
GAy576xi7IGkjIEy6vtRVk1NtIMXNYgT08941PqtmMrWrSwpwq9G6Dd35fFJQRv9
g6tSTSuJDmnSRUuDB5UJx1pFrMJ1K5Pp7eZORna/sYLnza3WoB+sYxREOwadEgWC
2NDBCCsZRAcZjxx6QQ4QVmYpgb2tt56QduRp4Co7q2OekuDKjk8LsXCbrakYhU+E
+I4QD4RS1cX8HqZSW2sDvsg43F/nNW2J0hY8d12HDSGYxIrDkT/KsrMNQvO55mUt
2y/8QHMHWzVwhNhXA24rotKexqmaV4Uf8I4bmUAf9Fo4fJdMmhp96HkjE8CCUBip
ojYXxHfC373CjksLpWz74Q==
`protect END_PROTECTED
