`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ktB3VXmKGO8/GOL+YpTm6ux56Mk1HAONFur/9IiSWQgojbGB40qCuwPfKGC6MW/U
BiPgzaYRY13+TxLZWkxoW3A/RJDluVG20F3a5KmvjC0+31FvSUK+34e5X/c6GXPF
0tiqVQDAIcT/lM01YBmQrXjEchDQApDWX/AFyOK6VA0/JbjswWgfw+DRdlhpyhD7
1cyYYKdEwY+tU0noYlVvJUbpOVygOxjVG6qk8HM13iwDfycUYLu1JGNQZgSJM5Jf
1VOu23iVqsAhV1uD4KKmALEJ8R5wukMmdwVd8znepAG9h1XztQcuDa8r2hLssh02
0dPyGRvFDasRwjet8OPCBlOt77l/pflN7KrsFHaTdc20TVplOtqS3O2fxyt/sl0J
8Ut8nMay9pAHRTIFz740h/S7zBekNrbvMKWQcuP/fWTeeXNDXBOBZ5rtpnHV1Ox6
F+NxX9hwXfcjqKvI4NJBOPT9RtXSLFts9tuCcfQVaQE5uaYPwyOhpDb+bcWfjgro
hjtJMGFR/UyTWBQTjvtYSeS9BMi4fAXY0L1s8b8rSmmUiMjNM8I17CII3/V5uLRI
bBnoaCir0GU8ihqw14qUJY/LaXsgKdh6K2EOyaet0QioRfaYKzgOrNt2e0GPAX9K
4QeDb6dY60IgC/zqKBBLVZJWhuNEAjClnz7vyOtrxEC/v5iEiQOSXbvfjJPvSp5d
ca77ZeQAyFVBOowUo7FDPHWa1lRHwrbLTt3iTDiLJluvI+CD7/o1vh6NDbjg/qjj
QN1DdMvxD44XmSFZ0fKIiw==
`protect END_PROTECTED
