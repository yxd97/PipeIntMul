`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQOYqS5OTEJszzFu8C8xQgUhF3a1/vWvCtYg7bZ3GkjnBg0hHq+dBKBrAhvPT5cV
tKD/yWV9ETs9hB4m/HOIfzuI/tQT1k2dbK7hYjVm/mqv7BOLy0ILx3A94uYCln71
JcDMvUkjJ4SO8T9hz3znD8qKrx4wrrAMVStaKs2AguUI+YrdCNZpaG9SPQke1FZM
UEX5mPyKXa1ZmdahzR0aVNJOKcmgHB8kviGRiw3c2u5IvRYFgjXbVU87PBeiUH0/
EGU2p70D07clL2c8p6lMY+Hl5a9lvlBRTdSbHN2gtdFXu1zQt3g8Zuo9U7h1iT4e
RZ+HqVrc1/xmpofuLFwUILtKNq2EgvmL5P5libcHCGNswuCvf0DLiDSP6NxbuHyC
4Gtk4Qav+nTBTxqAN1O5k/O/tm3hj7XK5XPMm+NlPmU=
`protect END_PROTECTED
