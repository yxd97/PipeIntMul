`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BoURnc7agbeJYEfECXbxflntIXZuPlHOXJHiNL7aXLG5+/3e6aszlXFsU1wQajw0
VdsS2pia1BRDSNMZociHzE2SXzTCoOiE5V5m+w4tOlz8rAw/X99EVfknMoqWb1lb
mA8B2wIVhrrxzrIQi+7qn9Df4mn5TDJsSUZbmcHHLa2c60wO72Zn2kr1by3JGbxo
t2wIVhuVvyZ4fUoVtOrcHCt1ys/ChQcrd0gR0r8TqimwGCeZWVYOnEc0c5PfK7WG
cpv4+S03WpW5fhzAJoTkIX952XHiOnUUU52DBa6oWtPFkdDiIxBgoSICEt8QstRw
lRgB+gqK5/7XrddRtNy+p/crm048Q4FpECe2Nd5oUb/eibyA/BMmic6LpRJUGNZM
mHVe4l8f+l/+RAwe+8i0tRL2CEq34BrqSIEdrM1BwptzU3TzpF1RXw/QvmJdNL16
9e6k7RuG5+WVFhXQSQl0CUKpMCKNj1j4ZCJ4jQzPIcWtyyLd4HfT6y/JyMUGzP6Y
4mJcoBE22fGowHPZbAjohTldWb+I4tCnMtNUNU97DzWNPJ5xA2xv3XjBuyIgkSQL
99EAH5SuL4sTrdfblK5/vRmKHZdp3j0dk7k3ygCbao+6uwPa22W3soCbw/8jcpfl
kuy94dFKKbhlxvJQlCF8q4TIsjD/tJv+eKbKxE8+70OUVYGXtNv0JynMimOVzX1J
7nLwQbgIVcsH1vu4hLTS6ue8vI31wHY0tGkIlsrApVnYZHoVw32sL5YqbLNf2mXn
fRUuOLDSr70Znm9uouRFalmBoXzm+5cQyjb/nrdOY1yIyahR7aVG4z6jOR7+GqdC
pawoh8du4lNIN/MYbSsZPtCA+od0WBSIP7Wsia3h7hbWuAW3SwM4NfcUeWMhoHFa
t8MN8HU8QRxSD7IHrOv4jfdUM4RJudMqQlTtcQ4FickT5F3jOuVYTHHLC3a+Qu9Q
qtk7r4H6eIiwLJGlzu66Hk7FGCqIyGGRpOk9caq8ATEwE/2ExwkQSJ3qA+uUoUKV
Yq0SiliRRafNkxndkMoRbTol6viLVO8MlkmHF51XVq+jklX9sLYxW9OXlCfjk1BL
/r32MWms75/lFyN0uRl9CYIJPUj3ENbpIXpm12is/RpN1zOfSS4IoY6BDhtgf9di
YvX7rCUI0PHYSjB5oyk0AhHUtmOLRnjLJDTlLh8P+2UCkhiaXZkiYZN18DE3a8t0
K3YbaBMkFEUl1ukxsOhXMaNN4O0OdGaw5/N0pwYoKgiVXzhjrG0dhxr4ZQxY0ZfD
QDl7YGNg87CkXUNaSk7K47vluX74kl88X+yI042Hn0f74WSnJQt/Uq4eYdKgsSVO
fcVzaW1d+oqIqqWeApA6NewMvZBqQgixBQBqDN7f3B9HNY1sevQ9UAdtkq5HtZEQ
OST04IqCNkeCiV4jNvSmJCfdGfFuyQqcbknJ6GSffYWR4VwKqypfVJd98ycHWt5r
TSpY2gZ7t8E7hqfqoLq8ZnJ4dQCcBwLWoMX9MKnYkhr1kmCjBuBOWOhLwcOyFora
DFRDilzfniqJ7v7ZFn2kVyl5JC6b5JW8Uepke9T7LcU+IliOzv2L/qBqPQpdJ63F
p8mGER9hTL1p4C4aIzo5eWzN0mZ6ea/aRfZkz0gNlGc92Sy3Rxb9zP7ZYX4ZppRX
W9h+ig/OyNYgadyjYMrKWFGc15xWvQTK+bB2vOTQ6DwktZh7gmDUu41pqbd8VaNX
CDaUb98Tfsz9M7cnq9+TR9hCiCmC5elpEYT1dQ9GkE7LwBRlScZ7KgKT2jT+b4LC
lRdlgRGxBeJ2R+rYnnE+Li+a3egOMB6sL0mX9Fb2nMHaJ4c2B0MNf5KF4K2DW0Da
FENtXCb4ZRFt+opToMu143w3korWSbu7aYtPDn5qM03x/E737kRQh0IjiILBu8vV
4ZXWQLgulnUTb22Rqkm9HQUqaA3X3F7967sFY+YE7pyYsD5YA6dPPFwZIKJ4TBpz
JHr9q23olWBT9B4c6OEB06M2eHxz0iQTFJ3zTNzucUg3wz/VefDl6YbtSGXroLeY
Mh6IiTWkLi+W0eXjVhyGsdLozhJjMJ43Sr71hBOrkMJ4MWpLjaIwCzj3RsovHSMn
5Z746Kb3CJIEkEJMWAZe4jFx2TbxHjBeTjjcpv++LX9bnwtx4RdWyHfn5ZEMT+j1
Tbj220hus0+LB/Cv/6cpz2/Zb5VXh+MCWXgCVxoHPZrE2lUtrT5w1odVBMDrUk7g
mcRFBYFoluuH1pBQsUczfTVEBb4ViRyrgCyRlPz94ellipKysa0K+NTT/avq6/Ma
lJJ0SjACSRkUVUSGWh4Vje89GYKNoJ5sBUSNSJk+dQyOKOWL7DPpbLC24Zt12Yz5
Z013fUSpQObtSom4pL7EQV0MNLRlednowzQQL6NEl/BTbL035Ul7ZtrlWeUc1Zi7
575RuWW2b0jKsBX8PYFnTcWnCCldfloCv2oIirYJoiE14HH+802gg0OmFbYxtVlh
RfglO2MVgsEWpdA/W4tYW1ftznMbdZfn9YLm/VH0wuyCVX2YCn7dsAq7JogttTC8
VUHwdn81VMtODVCOcWTJEpSUhKLqEzO5r+C0WoJw6wT1WQ4tBwM+dJ3O6PIvmpn7
W63ZHF5yjE9HaI89ConJAnpsJhfrrLWyKRdizYpsRfSSFf3NsulYfTS1T18RStKu
Zxcy37JH45OZHmaLi4u5Lm61+wJWo79vf66+Jg+wq2We6YfFPG79BnsPvAtj2gdM
fmTcp04LiAPdBpxA4GV9Kd72qXL7V90jmz8/Hd6zbe6muvjNPuduy4TwLsZhfb4d
PoRhz/aJoK6t/45z18AGZupI9RTZovY/5im6nBCww1NeWtV0ZSnEgPUpjYKbx+dV
uNhr3vyClHPUBc8oqzP9YYkDe+wP0/RdlupWcWK6Pry8GQ4oBfDpXT2+PVOmXFBI
4noRTQkvjEhYFylAJPcxSnTqsUoTiZJ4YUOlrHHpnHyH6OVsMiMuhnIs7kZ+rzjz
hUocpRqR6OSZNpEfGkvXssIAdGVHOQ9G35PYCwLHFtQ4kS9s5oyHl6wFXlS8vYA0
5YIdTMsAd3B9qkXRhoicp1uDSogAzGz4Ag5hrPPn+U717tzr9QGW+giFRFs9SWEs
+DpwbEyOYLIbH6GJoWXKD3XcGEIWozGqOMlesfPnl/cMIwdgOCAW1ncLs3Kblaxa
5qS+73aQo0uZ5/qh5DC5apjb7USDDBRCU3llobUTL76n2I2Iku1qyVtXXoV9xR7a
Cbqg2cRZD9wDMbMyxA7MZd+MVmnoNFjvTsRdC8mKJyfh6hp7j6DzifPNo8YPETKi
0IJc8UvTgqbJ3p3j2Fv2eFN9pzV9To2U0eNslFQd7DAWYgaqI9IsBzSFn91T1s6G
1fkskLT9ngGJmmZSXQdimR7sPrBoGZoeYeTt+xesYqvrpy0ZRPftEG0iCpR+iSIK
V1TzAakJ0HGD2fFONhK0KmF4XYEYOPG2m74YhFMKzGsIrC17baoYdgdhDFLGoenk
lGg87nsl/TzUeprvpVeOIcZlJCoD0qi+VbVzbAw3dTntec+3ITZ/2MemuEM8ELAw
6zMhZU6U3Ugu1+wG1dH/pbN1aJEywrmEQg5qJ9+RDMZehhBP6oXAON2/+40FBTLu
3AyMf4qbahXjo+Uh6eK/FSnt5yWo3FV1CRbgBgzJFABmy4OZevsyTVyftNJ8jZVw
Beb4NiygLVK10KlP/TYZVcdmWbVBndd3VqD+yyk9+OrKd9Oh5/UK/u9Rgkl7XXeG
5D2Q2UqC01/txr6J14mR60HcR0UYbpia71MhzjCSg88=
`protect END_PROTECTED
