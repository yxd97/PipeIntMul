`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6J4pgbNxABjAaUSL0F0jX+ZwwDE0/poTYini9Rxvlri4LvlswSUB2fygyk+Es6U
gjzn8g4dAjuqsGmWvn6o5wY8NQ5lnep9oxooBFPwuZshdw87zor74GhQZgyoHU2P
SA5JVQBF+o/KHZsWTs6fHL3GU/pOSrqMD69CiV9Iz7K+k9ViCXxaOgNAy39qYtGg
mOnpTjYAr0+sAqQwrMqrSZOzbLu/StLu4f3c+D2mNxqgJ8kQuywRXekYNBj1P8ln
qtXLKSB+8cMkGhWGwIKEYuJsgP6Be8IISuB4WovyUu/pLtaOuyn28FMaL/Z+60Cs
77Q5Bs0d3CT+pwYa96xJjQ==
`protect END_PROTECTED
