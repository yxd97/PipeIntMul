`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vAECOL81BBlYaoLL+6TMDe8tYILxPurr39bAGOyzGHeB3dE0jHSnVxVPzO3vSeaM
/5xmCmAiEJByMDcZxnXNGaLYB3RFkxh6yzcjvMrFV+5CPD2SwO1GeP5zi9zCr+n/
Lq6TiX608HHAHlwFz/TxL5PQ7QfUL4UHyT/LwCjX8EvnI8DvNvdk6k00iCdUcURt
e0PmuTfFM3OP8Hj7emQCiSc0SVaa9M4GA2m/wCXZTgoibTI5lRNd10AO0XMhh3is
dGgX0BCdNA/HVOq8HYfJOSuv6GelCZN/xrLYeManInw64Wb+VlccEJKplOuQC+/P
0mbMvkR3ErMXTVYZc/jG02qb7jk6d+Vu3SypmFbredNKUL1z3NqtuQpuHWNFyqN4
YzAflAwQ8C+mHKcQCRZtprLfX8OvZA+JjqPKeZQsThrEdS7wtv0yaj7++cydTEtZ
Vmm86+Vs3HiqqqFFoWHA9EUc/C6zZdIxPulQ8r3axb5eRvoshaqcThObB16kFIoH
726kE1lqm7Jpantlcin1wbus/ig4bj3MxwesuxMjSrCJV0q4roiusnjwmsBkWxRo
OIy3vPCTVsyeJbx25TNC0NRwryUHh99bGCyUA3tdQE0/Rk1aUsOhFeubrwGAm8I/
pj/BoL0xeGah7BD2Dcx/cRtlTvgfcf9HZc0KunQAMEYvCWZ4H6PZiVqT30uxwcBj
t+MbGaRcu5zmxYTGj5MJqKnlYYjCR9I8n5skHFCisG+jURbB15sIVVIPJCZBh0XA
zitHDcektt0OaAR0g+Pvc3Q5SwCjmT7DZ5NpHtaFbKWSqjl4GKKCTOeGtSr4YizC
k5ibR1lohGvTrMR8/yBkE/fG80jbWzKA/WlBpTpghOL6bbeVodBvSySGRIOPqqUQ
n1hkpa/C9fvechUUrLvX2d24ff0vwC5hM2UzEY0I7gPuzmcPTmeS6Rfs0+/arUmH
LF/sTdzAX0XjskO/D4YvwqzSi3i9Smx/mZ7+835/ZLmgtnuGI0yxBFRD8BL3NjIR
YHvtx1P/yS6hzcmAbgBywJFr57lOcJxbEkATdXsa7lpy4KPNZCMV9vgfqYxnes/W
gVe0oc6v7zs85t0Sqk5Jli1FXyibG6EAjMf+eIn337/Eeq37TekIGgRThvCn1li7
M677A6t2jl9qVR701btdOUO9J5koHIPz8xdZz6nr9KMQOP3MOBkamUKx7i7clCin
cJ2VLbQy0AVmWnvDLBZhpMQXkythCAyjHNZk9ix+ZyKG62hwV7DFa8bWTD04PZ55
Qll6+Em8Grtd7MbgAv4JQLXBCm2Otbuu8QW8HdAT9cFuZMT66h8hyGZgOGbXMvzr
BZ0dT69dnWUySowXW+JGLs/b0BoVTLpzbOM/TWaiPBayWq9Juheqw0rnG4iKaWPj
QX3RRwdZENDoEnliPJ5imMrBLza5mv3YSrNMCK5fmjmxzNKAna4G7kplcOnS7G+6
zzFWacujqRaDcmdf3nGpVJD2gcLxGJ5pii7UloAoV7BIYtqAAPXagNoxsejflYBM
eqwNjfkN7xcBJItGS3ChwgTIByWSeCWq71dObF9rts5Ee2iNpKYHbPiSHOW+tWkd
ZbnEqL1NGTpCEOAY+NxxPLybFL4sUE2lHbWZs4w8/Q64Rq6ejQuH0WNyOj9OytM/
3Jbiq3w0Qm1k5b3kIptYJT8ZvBeBjEFXKRqk8T/jp9wZs4pzp23KhfMGSSXYb/eU
TJnPhEZxhZb97+atRWL1XhjVnfo3IjaFjcoJ58WRDeu34aw73cIyA2oLMBtg6nkN
O2n6zeTFl4Wka7IUwWfB+f11/c7+duEaM/F4p2EojViPz984VqH9xkj0bQAgt2mg
kxbJRYG+ngUlBw1cdSP9fFuuREpQEMTmboIM90ZjmM7CnGAeKi+HnbfGAR9fCbbo
vkjpy7p5kv3sqdbNYk/D/plmpNstdbaceD+/WLI7SYL7yLNVu3Szvmaov7Wpenwf
WhB1lLnrpU0D0siqcwYnOCS2+6b5YGjoND93BKZAT0kTaqWokd4+u4GXOBNN7qfq
Kn8qYIYJOgt5SRQg/4Vz6OJBDMt4rDC/G9wvvU4ezPJcxn2CWkUWyx+A68jAoaLq
e2nLDztaI2SfFySk+FvTthHvdYDXIX7I4YA8Kg+sWgSBPjL1YEhglISuRohU93q5
4fEiGiOeCdn5Q96nCWk0xBcCcSdxu495EFTT8yJHXKMCFygIOzvm4TeoqJl/2jR4
lkQnRSuQ1jV1Ue36MMzfFyzIOhEn7Iek/c6oyY5sKFOAmXnmfDEsLb49Nl6CW87b
2FcV55TjkaUha6jD5LaiYVJrIIjZYqabZTBlzLdM0fugP9L/3hHmj934LK5p9v84
vNYWy0i62oVGh1rGvr+gxvIDw84KiPn2m0wx5cRbl7SAimIRDmJohWZpT+xPiuUU
uRKWAy5TYl06HtgrNs1EN0/8fuQHWftDOuweTC7sojg4aR/X5bno72QkflscqNz8
OruaAXTuKcq0S2g2KQxTIMjriHch2+KVew8du2qsX4U3pGiWDNq6zqrKE1QKpOgz
gtP92qFCqpELGmyl47B7YVJYHaVNd7KaBsMnTgM3rKsm0glJHEFsefD9iYii/hpo
riFc/+rinWpJckQNQrnlc3Czjb4HqVdbdfAC3/MditvSVKFjH26sKkZcK84bZmgh
P8frjm0ClU7nvNk0xJBDjDH36ohuGLK5KJ1h70gguhy1x6/nAOGFPMX9S8j2vrZP
pKOrxK8dp0iYssMKtJVbGEHsG4DJnoBw4oPASBOg15ajQeP/EfiOw1BBr3EFBofv
4GdZYH+9qxiBZPBKf1XUdSDclCiIMe0DGr2hDDJFBGUe9a6DsSUQ0atyhZeXsdd3
sC5ifpwZNikiASvIOD7W51J5MdzbHTHG2li7Kz8bd1RqZp+wuUVYzaEqDf7oWRFt
eyfhln2Kc0XR4PX+DCN8X/VO+/OJMjn9VuD7sINdE6sYSFCSpWTn4jbnvbfzdPjd
279y6v+FNBzJwQ260z2u5rBBmJDA3CTeZRtU8UH2NMlM376pXqzpO4oKcY8j5zOq
+Jjgvt1n/UXSeplKCFHZ+EQfgfPYGnshHp7cwnUdwoe9wKFIRNO7YB5vCC7y4brO
snOkcVRstnFOX8zG+3CnEywdeHxc3wPvuiAKOXTSE7fVZZAWa8Jv/6LNnhE4ytIU
gB+gcXiDhH465X0pVnAVdLWKbuIxw6dj7ZWjay/VCwFUNW2YfDZBD6Pco9NjQJQI
ZWbt8fPais7eg15/L5WL4wFWJrnRg5WkjDDDleARE6WE+onyHbDVfyf/GRmkzLAp
SAWOnP/YhI7+nHAWPC+Wa101AQJq6sXfMKKJmUzcbet9p5p/lEXZ9gy7hnS3pArq
9Y8JK/jcX5Mr+QWjKZWRW56PseFU3EVX461Kmz3ruJWU0ZSW91Jkq+D7Pk5a9JDY
7mzECa84abI8GQPGQOt+13y8CsKORFUOiuv/TvEvIFak74f3J78q51CnA0LjCm8l
nUPD/xXaBBr7OKVfm2m4cbfEh83OexUIz8F4gmivgwkyqHdN4S2bEG7GIqxnH2ZD
NQIRhlKVfXy5sElKMsegukmIVE1u8Po9ApWWPFahcyy9oNzz6x6blwvImKXF5H+f
JiaVUPwhuSBEcBT4XJvFez1772OIF7dMnCi69OBznagkuLuhVfZSels0rRs3Rgi2
7U3/i9kFIWJ687abpIx5rG7IQM75ZnOku+RWHNaOoIoi8OKov/skzmEfsaRADPvZ
VwL0Kn9LFDxaKCeb2Fqx+ukVtJ88EB1rh5CpukpoKReK3S5FuqZ7LjQfwx7eMmXM
U3I9au722uNsu6f7UvlzpB2hqQ8orhlvStfP/QB/5Yq1kTuDhB6ACEff7Fs7RYGR
Dt8RscUYxT+1JaE9iq6TyUAD3YBlpIrVoboX6doB9GsPxDPOaUggiflMd8r5lDX6
x/tcDw3V/mLGx0aYpVSLpxvzjA502S1CSgzsjMvZ/yAXfsiG6/C21FujA6tz69xq
bYd0k7OD+Hx9hBScCfwViS+SpPwnvdB/tuurJe2zLDl5ue1QRkGs9t0lINcdUar/
FOQROYoSj1fRNkHNUuh7Yj7Qq4HRypjRszrwy9M+/PYoh+bNd+caliPBfSsi5HB6
hT2LKEqiJDJxQiGIM1bH+S2ZU5/Rt+ddtkzim47NiiWo2BKnGQ+mWyBRLbiennXB
0fqIWuNTR5P6IV7dPrDQnMXNtIbAvUMfYxJn3HHcTZ1Qp1QCMvkn3Q/SuK3PHxox
b7lyt3mdZsP6KcUaO0oj1uhFcVYISVbzfmdaBa79Ik0N1P1OHOaKmR2gaRwf0Gdn
co917kKpXbkbGQjiEBfMZXh5XnrYWmfiSxj/WTlb7Q96iQlHvpIFUbLrguVW9Ncc
yJJVeZqfJGgNaM41ouZjP7if2+pOXr76+Mtfx9hakxn0eBd9M4KRJl35TeiWQpdj
XkuQ940SaRtrp1xPrsH+9bU2rXB5At61lUxghCFGbySrK0MO6bD1bSXDrc5Ir7Gz
LMV1h8nU6OxBS+DX9I0pOrPumc11oiKy3TVFX8ksqeWx8Od3yI2tzrKRb8G8+HrO
zbSNnxFz42QcT7vBqc8ZRuWZpoWg1NV9yfvUDkUfW1FkE8zYA+fB5NV4aUlW9qk4
KIJHpaPEwiaGfh8V3VNiCvFPPqYPRgfqKBFbgT4pyyujlA05N/8HvEPc/ipTjoqC
wjOkahBreUg8cAo3CUU6Rz7cAVjKr6deVpI2Dwj/0SPKp5OgoWD+2n1prgp2dbCw
4U2Lqd6Bqh8hUAAjvCNLIyluVwhUkuWIBEVSf3hH1trLwWbTEXiLajWMnCRKJEtc
Mq3DbmNwjBtqek0SNrM645QhkLGa/GMKxfPmSx4u5bIWsGilBPNGHUjUAy42CMSI
bnTs4nN32YH+04mTQDEgegMFDDYLWfSAgBBplEAGC9KQ32x++JFa6FkkrH84Hy2r
r0GyLLqspN5UUlg0pzmmfqirq6pliKevY+LzjIXbg+VK1Yy0+0s3BdBGF1RdOaf4
vwRIcjqsAz2iUsWCVamo8VsAOO2MjT8PuGnU28BkzpuGpXYWBU+GMbStvxib02Ci
MoXS0F4eMNOjUf7aYPbcflcyZeh+ICASRmI4d4u64MgDX1Y3SUqlrRSUklB5mWcP
4BGySc+yAuTQ3/ZKSAcvcisTqKs717ee4hAWH/FYRvAKMPvP2Kk9Cru5FTDHNWRz
WdYdSzhpTygENXOKJOu6nZBVsApAQjjvUSieZ89O6Ribv3vABOwFYKowQyjwhYmi
XjxjuzoQwSXQzBmSiPvICSJlo0Fee9PrFrU7AtC7b3N0cpHHRzQP8xkMkRi2NFX2
GypsJfJWJRVe4FqpVUB05EaBivkcOAqDJ5kAjYUapuq4lldb1z8ns2BVo+VX5mZw
KHmD6CqyfCxFLVENVX2KZN+6j87/mv6nCGTNZtKJSyjavek/VCSY5IlAu6XiM/Dv
/74X2hM9h0K3ik2s2OxUhF+gKzyeCldo6+FSIQIxqSGZNs6U3EkQ/Aeg/4Kw9ss1
mLwiYumjhnqy/g7TjNXki3DOC8tjwoZ7CC23oq+zIPs806Sp0+R+giNoDnWdZQno
G07Y/vGPPGbtMARiwvb/WWJz3cUNLVebj13hfsEIjR8ko8rWaoYuGWO56jUtH7gg
QgR712MB1+OuRrQL59epKClLZYKBqxHtkJx1oXve8Sjk2J10zSiO2oC+Q6c/89ol
ZFZdf2R9f9+ipE0iJ1OAsSG2KweFhN1WaxEKE1NkCi1+D2CIePep06AgxSZqn1SB
HygjoE8pKfoFg2JaeMPaDxYY/tjPtJeDEHvJoD3NU+EMZlH+HuH76DXoeDFpnUNI
Q8QNdrC3uP3/x58tZFIYQTQkNF0Xkzt/g6XDv9ZL+vS5K8tXcqi2tsCPErpyME9Z
wGjsMdFoIClhstR/z8DgxzWspU12WrWzl3mNS74PAeXxpff5rd5ioNN8YtR2zuM6
KZinQwGOorYOdpA/4mHSNvYyJRR5EdFJSqNBtnTflycLfMtlQYtDsbmVmPJ4dcCg
/lwobI4tUjZzE8+FAsY1yNnBLBIv2l/gB++3Htnjy3NPQTwMUBaR2lSvCepmsMcl
1FJJ2hZnDhNM8grggZpFF5/b9WNULMwE242wFkgosHUi6OK2e2SYLFlhTaNP/PAh
wQx0QVJXL9Gep6BH8+Pv4QlUqWkcgdvV25YuqZi9TcsPpxRrM+DcntekLScCrdnw
kpZsP+Pl1EXkASw3M3o3RY1iIeV4vNwHkyHZXy03kSQgeoqwPpBxh2QIlFaK4+lE
NdhnfNFkHt0DU2YeGY3Ur00CpfwKu+IufWit9Txl+lsHLVpkn26B/NOkrVP7QX6K
8DkEEFPu9CL5m1k5Q0Y80sj5FhvSpFBlVt2602dc1rESEsICjhajtzCyIh2DIG9E
4yG84gVYzhpEDOl9l7Ikrqo30KPBMJ2pH4J7N9WdF5Q3+o0j4KsPR28wSq7Ss0bC
FF6a/JPk3peJttCdHW2qa/HTqwjdHLmdAFgPUWI+GacFvnxYZyRmCldLH4eNTEU+
XpMMufD8W+K4TGOjacYNJHrwpL6DXr4/6+zW1jR5SApHa2IGQyQqIXxmfkZPauLg
9+sbuSGsoXy6CPyPljrU3OoEKfaMYqMp4f/xQ9PRj4O76GDKSS4sujljq/NsAhDX
APhfYYtw2Yh1FNP/TriFE/EKcvzSZTIemp6kYcl+MYmuH8FPHIX6++uiSgK6JHKW
zXkkXNmgsGG7y3vEeHJ6N9O5zJFAVUKH45D++ENHmsIon+XgH5rRew/sFsmC1zCB
ctJMZZD2EmSi4hYe3Msq4vXBzEr8HdqpCxwzwQ3pq9A5bjis7x3vqyt3uwscVAhi
wTDpwCjw/sBtFYt+DuU+5tqHAMGE35FDxkE6++nHKbhn3YthiskgdzH0H6auUoGn
rug095BH0jhTx5xkr15CeM4HUSPv4CHeG1evREKCQFDJ0ETHFMjlqjdrYzJCmBai
JMbCfmpMY3T7y0MBgFUfsEmZossQR3FdYMARfiA4bVCHS32ybXVBnKoLCq/pZx0a
4je23L9GsG65Le/G4qW8aJZZzbX04zmPCsg7UeEaMF3zaXEI6pfkyV8v7feylUne
jGiY5w6YExobLv8qRZB+vdyByBuQuerjrvzYJgax3e8pG9sq58SYdP2IrTV2WfkE
2hhbVwA9rKgpQcMJiY2lLf/hRJLy7mNypeuiu/6p42aM3FC/gNmdkgcN/nVHENG0
tZuUCxb9+N0Sb/WgIBrMP5U6/+ZjHZHZSd2EVrXV3hy8zi+PL8o3QGOpEIKlZPRh
NA7VcCi3gFPWL4VFWRFBRDhlcHKGjDIrY98nqxgirbGJkrISG8/1suP2KsB2hAPK
5vpLSdcDZJ9+VHQcgT0H+82Ty7Me01LcA9Uo9Upc++4QCftE0GOyy935MJZKg4Qv
aOxN6Krow5S5s2PMZuVIw23W+Eyfir73qQSIzpN2RbmymaR0skRoN3t+poIeZ+oy
VDj16TFEPwQk21aSbHMarKWFBEC1lBASwmVhPaqdRGaoRvO57G6XKwg2EXlmMvbF
NCLAkmfTxrP5LKW7Kp7G2MvnrZzQMGhJCbatIMxH2JzazjRK+dZod+mVBK0b9Q1G
6tO76OScvDqEU5r4HS+I70wK8n8gpjtKbPZ7zEtV0YICHNQNGdSqGfyQY2p0payn
9t+uIv7D894bDgH/mgWcdnijBWGtu+RMQzleO8ONK3G8VUbLhevzF5QEYB8MlulP
Xga9q7oW47VkBJ8EaB+SrCKk2Cf7LvvT6lyqtuyyIkIeq2PCdNtm9d25yzJuyUk8
hrJAe8pBeTBSMOQtJUb2mgqAswMWI2btFxQp/ff2uTnbppEoTQX5kZJMC+wd8dA8
zgDEJK7ds8Onen5VdUv9XfqQ3Is8i/QL0/RxqrwcYitsYGRg/zdu8qxm13MNLZhd
k/3Yi+9rYxQYQcvYcis1dr/q5aA5jXfClCSUDfdgeCQlyB35Hl4OXYyrpWzmsLOg
wa/FpbA8VRhg9jhJuB1wy1Kt8xvj9iPKhW3ZzuPVvoLf7pvnLOKPhhYq2ek824O0
yX62f1tbPNhSL6VBvywsegCz12qfcyq3B4FS73+1OaAdIZ+90D/3CLf/MLAv+dgN
fybCz0urznXfRv5yuxQqkxnDFm6sUbqVwLv36a7uUyIAav6DjnM1Wi8Zl+LSTVT2
OdXmYQtv0n0k4Lv7vW70btISTXdsWaJ7xHow/t31X545cfX3DbryxxtVdA8o8YC6
K3UvKqtZbrvqjgs1UnBPxy5t9+nATw1VrZoHNqKpmS4XRi2HM/3JmSy5nB8gVXB5
1IVWyQyWxcp8hulkee2ljYIu9UspUQW88X+ay4OKlTmzCMMP4wZFj3espU6WyLY0
EcXe2v4jmkp9HpnFlYQQInLdqHoZiVTTtLXlZCnH5A1jUV5oefASYsafmJMqKYGW
hA9JuPUJnWIqye4WZR7rEiUgKxcLe0nGibMLs0kZwZUX7irFeirRobqYzuoFO5za
5v2VvttlZ3D4kbOJgUMVdQaESi+GUfUBP+No0HQE4umQ0DzqZMDK3GbWruI4Wfou
IlkbIdzjdduaVSggkWNcS8XfJI4O/e2dJCMk3HnqJUurXHTHuWVbsQrb3G0ZHcKZ
+iDDn9V4Ck85PpqlLpBt3axNyWcF+fjU25fMUrVeKATRmm8odB9A9mjaYeGp9wsC
2+eLGHrBvavE0jeCsxeSKe4aXQIbpK153rgK5J7Ajgv8MuRg+Kb5z/uGWIMvW/Fa
JQfJMlO/HHoQann92wypG/sQE+PfFCBa/DnLYYFGBnHLlXdOO5uY3P9pc0AQDh4n
BvQ9IwvJRp/6hZ48FYNESRDX4+iDxPA3M7+juCm7Rw7F860/08g4myUSdVU3RcDO
bOWqnTGGCbpUJ37tm3zPoI66UK5LmNGRyQHKaQCJXw4kvaZesJ/KQULavhVr9Kcl
WJvKEPPolg8Qc/oHXBVo2swHEpuNx0PxKiSZ3B97wlvxFvHmhTFD2e6jEPuDFvKY
btVsqNN5O7F9ZvdxvULPiGoqrAc8I0LLELIf3X1DBUVnjL/eqEq2tk5bGo0P8geG
620tbSxhjA7iqKcopAUOtxOUs+75n6RrI7PE4QpwkPIW1x62sSc4zap0QpULnjh3
i1/dCQBbTMU/ZM9wzpqhe3tT8KrWu7Jt7Tfu/83dt+ujHBJ+3g+Hg7zi9LCqUIbd
PH8f9Prsewv6RW0xIuauO5tVb9PblWYfyUcj2WzIlNpAadfYQ7PREx0DcbrtQcB7
cTXJBVs/V6h+AHoS2/fXWbzIbySWeeJ/I7jlIIHs1Bj4KcKZ3WuUdJlRWyDw+Mmh
hIa4IL5qo5/p5g7P1vcTitKZu7Nw6R04MjrfFeoacaVFXvUt8OEw3ZR0bj6zGJI4
47UopTJk9fOCPLuq3/hHoJ/3Lmz50CzXp06pgp0J2TP4AwSmmoyicfflzXfq8SvR
DMEJ9+fwwfhLx1M9pQqZF/G5+aH/xsdqP52ycHWAwAm2Ym2FYyu2u+2RBv8pWwt2
qLphcrYlxxBhwM35xeCMZBfGQVk2XoFC4N24UQ1RquaTnEoC2eczM5D1zAL9xz3/
mqJktb327bniR3Vz+djtdQn9gP1ZoCbmqjpHapQKbR79TbhtM0M4BgaOAj5IbpBi
2KAyjBFa025M55eaJGD60lLDBhXKAfKcSZVNusu9gUkq2Dozn1TcD0YI2meI0zEW
SnsTxjba9/y8IR0lPQm4R7mHuk1Pb96Z1yscHGsIgWLeUYJ+ivesByjyy7FYsNGN
84jAwNzaaiguaLID2q3vtTgBcwfOPqeVAfUhdCEg5r6At1RYJreiCcH3MbNpsccj
bpWjyv08lBnQxjVUZuIr9Tl/FMu3gjWhTCUg3Ku5AiJ/Pw6BiRV7yzADiKs+FfRo
ZGQOlqUhEhC5VBu2WcUZVZS8r1RfCkdTHXccdgY7SQZEbLGGLZUjueo9O6tF22Op
GjvVlmdZr1UC7fvhythYScGWkx6qhplqpFZArkNQjmfdasLKiDM50b2U1lUfmOrh
ra12ZvsMq5nUmB9f7ViFqsMeY5D/5XO5Xaw4Evj2m7Jy+IDCnrll+Oi/I41W3QrK
AhGkItUWfcycJ3CJsUVhNniSWxcZz/XE8c9xt6ZE6+k63tyRQyDRdM0ExBloAHQU
cVFwY7GLt1iiKynBJ/6ySRHfUVFYZwtYgDr4uMVb2/c7ewIKSPJnWWc+qxlZeKDj
N1pWDlZmT5kqzHso07PGXU8WFG9GrWYYf6qMuxb9eRdAmlcA059V2PH5WmFzptNi
TA0NJXo04YfhEtOLsy6zK0gerUfgp+8ZMXStYNpOx9hkU5jOAJpuXw2fTkEM0u/u
QJShUON2JuxwUwJOtuI+mfuFhk1vJwWMOvdfHgjSOYolAAy9Sg0kZQQRdsbprgYT
kum3eFW6b6sLl8T8tSs170YhZ03sYiVXggI42GliXusd7Wgyk7XXfLYWZQGrrCTQ
hIO4CIYw5JqFs9BIImyMIUnnq60ogPjr6s0wcRlMNxDiiasNHAS+ITskDJGJm2LB
sfOIjDXjuyrNzgNXzPkA9eFGnl0NZE8XzgUbsOvd2lVpnKGUyl/CB8W12K2oX4Mq
tkAwqu/TiLGS5nXI4ZTgkXNq3SuNt35zvPV9b3Og8MDt9tIIFkLOSg7xdSxRJZdq
7oVSEnV+KuVxyjqhRycYwfUE9mJ0aMSyq+QDEzucWhLDKZ0oxhZ6pQiAtkwByi2t
NMrL1IQEI1iGriuktA6x93PosPx1vrqmCMDZaRIaRMv+dJ9AN0OAmx6BixBFxBe2
pMZPADIU5ydbpfuZrIkEe3/spxjQnQh4kMALynDTBBma2sArBtRc++PQHXKVsEsu
jdiUFRiuue+rtcGRDQB7RAhL1RqCjSZbhs5jJWkVY86qzzLKEw4kTKLEd9yLIVot
kllmUg6UkP69PVA5HFI9q070Q2OTX/CIq7oluTyV3B81PDD7tKL4jBV+nwTz+5li
SX83h1Uj/Qc7k+HFRMyArpT8q9PiB8IGFkTfOuzMvqT95sViWeP0X4K+2okt/WVI
HXM6Eol6gvSIXSFCiU8RXdi2S7LdaCHeJCVBaZnx8g5SiGJ+lZPksEhfpejOVp3S
5e87X0EHwakyUq2OPRU5+VMwu0EcQUG04t0i4mcLLoMjvsx4WyN+NYjToLZo1qGG
muFVr4AbSKNjOvI0momc9r8M+ckkL8nOcPk3oXDhwbQKfWrg6Gsgk3hhzRH7bvcK
ZCk/A3zvzu/W7xEeGzjhvNAuUjZV52w1R+jyw1NjolgF9e8qBQsV8Xd3yB7ruG0f
3I4doTjt38CgxDhaogZgvnaXIjiiNs/7nQFogRq7EmdChi06J8qN+KT2E9WbYRk+
I0GOP/WW/cRbxcs2A2xb68xbMhJSYABvfcGmVMI0Hs8WtN9G0tBKhiFLQfWGimv2
N7jLEAN82w10msdujHoxF49xwR0wR+YbbBkbv0PP6MRPT3ZxXmhWftaAFwQrkfZK
vVcr3vFZXDdyX4IV7rkwoo7l7MOvzSbl+kU1Pu6O6SU3gk7Mo/1awyRqcPBGRU2I
yJA78uvelVSz9HP0YxdFQ3pVxQ1wq0/TQHYL6j4OjQIHlyDzJIp4//XoZZmZooV/
dfihs4pz+1byBbyI7UkUqnrD3OMNXN3wLizEJgdBG+Ma7Q5xWPqvU/Xi3w9NYFNU
i38VleaACfPsNfavRdVONL9AAjGgPLrAZZ7VjpZjYl6YgyKKdSangcaJU/vqTHjh
9BZG6hHRTEEwnWiKEkdPYR+3WISGpGUDmaCN2AgAXKD4aQN6wCGAs6fJdwrW8A0c
ujR34dauHleMFmNdnYP+IEgmVjrtaWAOZ56F+U0JGGzV6Qwi2sGjwZlggWCAT6ub
61bMXbOwQOekaNWJS8wxzr57jDrK4e8rr9EJ/MPhqZP09hfbkfgK/f47GnWqF7JE
BTY3pvHYFgL/yD8dHcr/ZMVE2AXAhochc4W68Bl/V0lRen8j3v3KKWSDvkXeHm7s
k38r4DdKIlUh3Mc6TJoWNDNCG/EAwLMxEcm9O/+l766bbpWZf+1vZmTnIMNe7O/p
NBJBnY1YlbjdfpJ9ay8Vf0iip7iN3TMb0kMgCn/qvc521RMD22qR9V0MWs6LIhbH
Cbg7wZEYNzoGIh4RVvLiBUECPejP+jAcg5gbcdGODMbzY2ELhP9mp8cgKptzkgEx
pBfn/YTWsgFzUuerUkxf2erIxDiJO2qH8GGQyM0wj7EWIcl0ngqyRrtxn27iUcsq
bAlUiU5uV17C9Rwnj+rj74mJ0qS8FPu/5XQ8wrDaBjISI4L30qI5rfOI+3MwYQ6j
0Xwo1IfNqqX+pmxex9gDAIlAe4fiUvXtBUi9/hR3DWMDCDFTpzpBzT9ytKjZMd++
vtAILisajL5Gsd9n+GLJoqnqMzU1cHk/U2BbuyHgkj3yp6ODASlOVclDjVDKl5cT
jpoBKzo1tdMIMxkDyDYOjyBgd34eCkQgtF4bH9fznjtC0cgRn8fSe6kVD3oSly34
dCRhZvg2+PDYLrNfp/i/gAyzs6CDTKV5axdE0gQmM396JAvegzPtjUNezEjbRwEb
NQm6ABdcP4iN0tHP7klQIKWP4ueNJvdOJK6rvPkrR64abUKVp0slT+Xoni9yTnw3
z08cEITfC4hV9K9g8Xw6k8MHKwHBJoZSZ6xtgnlhHA42sOhe2r0LJB0gsi4EaZwU
JYPoMOBrPa4B40A8N8+Xh0ZKl4DBMV5wL51lXL0ONnPl60eSuOHVKERdhNS53qao
5jzSMyYgymFrvSF6Y8BiLhA2vhR0Cw/ZBfOMcN9cmp2Z8SQAnkURPSNXdfrr+XrX
WW3NDC8sBSyvufYPVOe95yjTvK3vc+UDJweqkKuJa2go5Qgm1UUwaiIiHKajyDqu
0Aczb55Ek92h6xDa5um8tQu4eqF5GbLuMYBd6ExAsTOQZPbNaQ/YUEdbU0dkxIvA
Aw1RD+WIsEeG3/x4HjhkTCyoNKWG42qP+SblG5cEL2uwCnKZ/tSZxqW1RTqjj/v5
raXubDHC65lOQChcB8cI5+yy/i6gVkpkQsc4iaCByvDCCYjlxpX6q7idx/rjS00H
SSuPI7p5BJCELRENykjT9HH45X3XnSeyyM4uwr9LjqNQX6ckbd1c1mNhbCYBm07N
/6TLYvgtacwc8LjJjffuys314UfDPRuxv9ht4KzjezaYq8RBRPcpdnTXaAskoAG5
OI03OJaLbaSfPYAhbJttWvzDac5q7pht6RYWVGU6zF8q3iS3/1J8nv1vds8KrIJi
lquEn7zOBwQ1WoKU0ZNUosNDB/qIWphYVymJI84qVhuS/ACZKCuRWeN53yuBa9GV
etiZ9lU8x7OkqvZsrbGCq0d1+8Y58pMqPI5neHm871Q6VThb4QagCgZ2FeqNyiNz
8g6Tpaft39SbqolOyqgthr/Sbn3Km3CICJKoEqSgjPvf/zgv1aMaQO7l7gUXHhfE
vuvXjsNFrBHmIxUao8bjqXxVoJToRuuKYilGC1+m8CCvfKV+mek2UvnqlfKKPpqp
VPAUpDtqGzxVJz2sziYyGz0Q3RcBwpfRH3BWDHboF/QEU0oI5OGdu52qlPIYW2DF
bQvW+GEIP3o4nZMX1Bs7cYwrQAs9kMJDQ6x2egykviW2n1PjzZB46vJzhPryeLTG
R0WIg5rBESvya0N4rUqxsyLtyHzA0JriT8SdWFtk07idccmGO8+KShb/4aHOyxkj
kkxLOWuh2h0A4+h+HMGw+OWDxff6l33phGubgRS6cXv9lmugrHzpDdzGKB7izeFL
0zyIF4d9Kis/4ucxT167t6qHdu85xkU4iIU2t6Z/sPRIBqExBsfSZdzR9KEuWIx/
i+5RqVzx+OLqeImRzpHDLyMI55JucKfgsU7AHM7pOU+IQPWRxdZyZxUxCzGvfLho
xRyKQlVHRwxzkyNyE7McmZLdbaCisbYnX4ICgK3ZOcqYjgIQSGVN5Rzzij5eDNWb
pzmvg+ORp8vNiunSAwMIDLO6VldejpnCavNkCJDnosaNKX7kUHuLlbL63VhZnSI7
K+3tQVgqsATb0x7izkNuz09CEv+I3DZlFw0ZrcNLwcDN/lBJNmUqr4TJgJ1yJnNt
qIRN3c745N3MzzvJaAw/eSiz0gHA7uBlO0bYE+na70j00ABQ+lqv+Ma2+/hY3XaJ
QudOSMybl52XXis2LQnHR4LJnbLam5oznevKKtZXI0WvBBLP2fMVTFQx7nwgZRzi
5NgMsiZ/YgsIaa/n6JazwxjNSXuqt+B4t0sgBGTI80p9hdDCI1cGkfHF8aNxvbgE
M4FLAVhw9v6gc8WIWKzOAjkwyBTMqGqGm41xTMQpcJHcewBl2zZe9ABJ1ddMIXvc
q+VFEam39cNUeycAW30HPZ+GGT7COGCR8yYAyEvdiwgRW5pFWvcYpajfl6NITOW7
e4/9xjt9Q5naM6QJXisEsHcU98b9cH2+oQlY8oVPGPXdcmIurWROo/c/ICfzvSHv
RUSciUVA4NL5oopdS2nCSKOF9ZBZXlthIMUzRZ+KtkvrptFoWWgD6pWktbmDY86A
P9noKtWt9PVHtkeIpnmhGUkVqHkPz9WATyn+71v/BLh3wVUI6Gm706Y9AHqR6jIr
rc4LgArUYMsptykjEIftupKpQ1Fu6h67y1sD7gcFarMrhoXuIosRORT0rWa8Ehod
vnvDODb73PxQA6rlRZw8DvZaJFGGo8fUUO3Hz56KKSxwPlXy9Wi8czNuG7bRK3/6
sGwAAxGi8Y0RNRUvzxpQl/sm56LIusv4HG/rhArqGaTclsLZBDwHmFw2c1FBux0t
gUnT9Khj13dBaEB1cYlS85JXYw6Co2PVlX8qwdxMg1iVG+M7r+nYplRot2rEq9cM
Re5KXUjl3+p7RL7u0lxx6PpmLGyNA0FjUxbnbClKVkz/joUu8O3MKJIhltOb1ru7
AdugIrt4K9DzFbuJ7UXuRlUeWp1hVAGEMfhoE+NvjzibdXUjHr5bEwjqoBZW4AiG
hLtmwjJxXTUJCIV4Zo1/T9j4+ALJbS7jW57wjlzV4/LTpY1B0BYVVf/dV2cGGo8n
2IZzahv6jzJxtlPqXDrxS9rgpDmf4q/EOiPu+W5usU+E7W3mJ3ZhuLkHSYnChrzD
kcNcWzCppqPBhCxnQ9baSomQBEQ39y9tweVPCUjL7b8aQcrqoQHmda6AQdXxvad3
5bWZZ/Xs6DCllzRJqWbKvFsIvtotK1UqXy6/TKrFCCxsxM7oyxjbFWmomH6uQro1
1LZCyhfSwijTvB6tmoIvrPKnc9t66+B4K3v6WPDAECty92a6n3VU7UboZsGHRWRG
K9IO0l0UyoVmbLo7rMJIzC4tYwU1itAUJrTmnMe1ifpjNODKl3EWIZmYIv15u/N3
uTYlA0afm8UDlr/NZ1fBTgSpTjT7pZ9Zg2yZCs1bc12yoXufdoCXCMxg/iKa/JiM
1B5gWsODLinN42xGkbFiskrbKXfRjdrMjmfF24TJw4vPG4VTi7CMXnSL+pzuweO3
/TZajbFhsvr6LMk9jd/FANxHPB7n4/vmjwext+pd2/qf9vLSq3CAASWl5KrUIf3j
y+hfznx3kxM6IXOkicflge/99WkhOrjBH+n4hbC+GKzBMxx37p7m7WWX/yelMuAK
j1k+6p2j0oww79OIuqVQZSu7Lc3LtJJom8b8WQQkUitgGSX9Ed0S6F1chLADC3LC
QniGk8ZDOwhdK3lOD6NkiOuf/oYsa3PHcpS2cN8UOA8aHLgviP/vibFI0vOqV/nR
ldo3h7HheHuKsLSwxI33i7uGPsCkWVroDBYaaO1PHBPM1pI/4EK2kAwwTuo0nPvu
02T6kU99QsQa6BfgxLoqKWVWyUWtw8hQDK39SbvQStOnkLY1iOdnYtKvPD7xH4E+
Vntkgbi9ujmc2ceJ/DCrW01kAt3+xdYXxypVnINwpZM8imwnWyjUm+50I0qRbBmI
/ZRlS1lGYVemGA6Odc6ODkvC5nRQwI4LYM5Lss36auGhow2C7JQxSYCmLaEXXTMo
IGvb0q74LUxU/FJN4ZnaSoW9blU9fHbVI32Qdh/jYHVKQ7UcNaFQWw/noacAQ12V
TRKqcOASU9C7V7fRcN9xLv9SnR1U6eN9Dp0FBSMWVOE5BpODVGKeI0qr8gHWr98+
zquuW9eqAV8CRube7admNuzXO9ePrY94F99IAqkM7zDcAE6Y3jRaurY/fT39BStH
nx9E9r24S/qCPsWzINFSeH67Wrm3ZZZJMFi9pIdLcfkJgN+beecxUI8eJwT7Zvc6
+U7hZWrjOUcbH1856duy86O7wtmCf67sdkLAitLlViYRSdXUf57U6p34DpACjM35
MxkCKJJeoDF5507ONg8+Go/n63eVgVMLwHX+b9r9z3GWEB6lGXvpRYCgUGXanar0
XLAKXfS3PwYfNiTOxBqOWTVJHQgmsB2VRM9f9LtFw4KPxA4XHL5r5lIqWPlRYM3r
WTLP22XmuJa0rBpQYhVXgroe/FLm8n+tvNDL7SmilznRBYHAwRNz27nbvrgKRmTa
yDoyhPueLzpn1us0TstFk5I5ChWcbK6Vs9Pyrd1BOn7CZa3NPuNdINIyb/DSiPh0
Yo9rtbJEuNPDks9aeIAXItLnb9dkSuijgXEPeRKcP4/UeUzZCuJDA6n/wnMur1Pu
6N41Dul6QdSsmIep7LP+ntu0qGtpftbeSHjILbyB9X+RvX2SWzvXDKLvUD6HanT5
hFt0FAbCdvdaC/JkeT7xIkfR2vVY42aCgixohIrM6JsIOohUyjk5cN5aR3eRkRi9
rqaOzkN5trMPja/3oZ3WQ9mASLxHzdxi1YPRoTFvS9zou5S3zrE5I640s8M9bO24
lrYjv+aSfl9hFvv6aK8s4rjriNbQvUXnDRZN3KN3sf+qO2VpQr5ly7shDbePY+bI
4Mnabj2z6+aOHxxzVDBhKqqG5B8N0DG0GVKER6X6YrBk2kqaVGSzPyXT1CGXD22j
vQCaRXNgDb5xYXwqwEmk5+LyT3rRKDVbz4/HfuXmWSuuEgBER5SUnGbZafbUzbZZ
goaIyUz414MgokqHrSUJ20aHZtFWjy3b5Xy43pXZsCrpMgLHLtFFznmQ+/5Bru2X
4n1prBs70sKBlc1aml/zvOJjya2K7eKMHMX95RFC6YjubYPUnamaHGK9UX8dsvNA
l9NwIdClMsWJxJmd5JMSDqtxfqZ2Z8r5AHIgjhPUzgz3z6Tfp2vZ9gRnkvBBlyQp
s6wtlNJZjGVAzfHjvW0LMCTu6tQIQNgBMNng7sT/AH5Yq+phh+vaeTyjaH0zaxiH
LE0zoO465fNn31SrJTaF/ETmd73k/94uQ+4onZRoWFblVbxqJwb9hug8mqQYbqU6
+UQcqmusXge/KQS/nAPTYkjgiLHqRAwiocJcQPBAkCtsV2q7x6r34gVEv88XXnQ8
NWG/myK0wFdE/bfL/tIX/QJpoDqZuRWBPd2pwiapKtawmZ0WJBktSUlcwzSmXsbg
9yKNOItQxb/6BQlk83AqigpPxDUSRbgN07oZFWxnvt8IJ/BCAkha2IXidAiZ8wye
6s64YH2/3qAXDFhyKQ/HCsdRJ5q55DOMx9v9MpeBLmlzEQByLfY2sr0sumgefecm
/LcSeP9VOvCQumsJSxVwSCOLgkaAx8qzaXk765vOIsxNQzerFmq1J4E12A8h25n4
GIXsA33grxMFheV511P3wUt++KO9/+lfHn0EvMrDwbDg7GAymsP2ya4JU7jp4z3d
GEQFcYwKHpY+FyY3aocEAMKFSmo5Y2pTdb32EpNJzHUf5Lw8ZJ7qcx597Os5jNGL
rwbKqcICyCDc4lmni7GA86wu1XpcpzeGwbozJAH+e/D7hV5wxPxn26Pf8qvN5aE8
c5Vauy4ZfQpEGZgRVT5SPFjWCBpSprPNbqRtB/IAVec1prP4JVdFOhreiby0vOel
8zE8pvM2p8P0YzBTcFqpTfEboNU9Eq0+qRkRDa99LHCQzo9M2VusMzn9k6Z259bH
wBv9wKm/JqxvLIVC3pNgZf1zuLxJCzPuqqBGhkLwOeMogjX2HtUJoADkrg1Nh3iN
QdJQQy24NQsRrI5ttx4O+Pciu2C/cPmn+13Xma38HBrV058HaAcKfy9ToccxFlvm
oB9RPZD6qMp3qQO65Oo2Ao5imz4lbcB67tGZLFmIE3EvMBl13w+N9HvTA+ugDf3m
Orw6zfmows/8o+trFnhoicv5DkryUfN1h9t6I9h5vWU2oArDJEzYrtHDT5va3b+M
b1t/mIwJUQVMtrQnzvojhFDN7CDrS9S5XLOBatN5Hsss+v6UOm/BUQhcEz7UuJit
7W9DjLn17CBqvfKVCJ+pVBp5nUxa3jPeDXfpggph0NC3KfTu2sUz8knK86UJpKDI
vl6XpaFkVhCpElMFf2O7MVYY7DdHcPdbNZthwy6keTzkYoG9J1+1y5PJzXAvNvCk
9Cl+r5TN0eeDODmaNrmC8bFHNpsCQvE2ZmTILo83AvxS1kvMrAv/eCN+SFkPD5it
Dtf11CzA7YeVfm+5aCnZeXjuQQO6mneH08KnrHMuGmJMRBhXB3bFt+bZIxe4pYIN
FkZ3NfojVJQczq83hSp42azA4bryY+SmLyRMwfNbj3VNMGtoHvDJDJ9IjaEPHutM
Lfi/rUECH+1ad3GjQ+TaF57IvXjVjIpLIZwCvSfYMwku1lQ6L+elKgUL4m1GxyS0
KxWqNilGSimquqJPRDV8+8AC9D2JXciiNAVt/C4Djof5cyGSd+KcSt4pG1Pi07Pa
247iDhVJprunkQvwReAr6L5+w0WmkNjGV9qzLc2Vg8WD71k6dhNLB1WYsSvaiUtg
AI3TcSXmoxIOz/9OH8AHcKlbzLgCZh09OkV+1n8yrvxcD2mgDaTH+p+ECOmyDBQW
QJcICqYJis17vZ8csxYywK9KRO51DUiFIreOB9GkU61MDd5UUxh1vq50Dbb/1laD
SJ87IsnTSWp66XV+8DUbEoFVMCtAVvT7zuW1OWa+N3JTq+LhpJPv2cfCIQxuuyvx
KKyBBhtAFZ+hhCI8U2b0tFBkDm8QDn/7yGqWA9TI7GP+gypGEXi3P+hbDVU6cPte
5IkT0lSD+rFYS7dI5k+m05gRSL3NqYuuEmwrXV+B6vRzz3TojBsUzjROMy7Osq9z
1zCfAEa2Ux3yj5VL/SKkwRiRUyfoP7DEOsBOZwSoVek9uKRvaTaImT0Z7CnRUB40
RypREhMZLf80M2uA7cfi+A97BHK/sjicyK40/t1QShdwmFh3ZTvttPWo/AVXE0qK
IUAjtWyjJaQfNQODwspOZezUC0ooUHPZxX+FtOD3xBL87WLBZdI7+1EXhqX6WPpz
4tNlEWT7eTo65ge+Vc2e03pmH6Dz5yahgZyEUtTLRo3m+qaCTz7kqoo7W7lGpxnv
86wFQ6CIt9W0ufzhddVVP/NMIrRn9MvBGVoPTsbKFi8Cb4qdK6Iv/3cb8mFZ0urG
ZXEMRuJG/CBdbTmppWzPQxJZJHvqJoKZ2CFHYW2iVF/lvsGWAaqQPYkTnhRGztpc
xPuljMoy2dCmwgPxpuCSOHnWcjQLza431tZE5CiGA1YVhyxUohBUXWv5ANpEwKOf
fG8TcVlc0+IhIeZKtMD+ld04xw8JDZWPMH3TnipP/SGVEiicYriT2+9dDTRo6oSM
GZfVULr/yoiOzCy/W2BY8bfa7pFcW0VQnR7JCzSRjlZUESjpJupGzqwXDmdc12OK
9ZoqdRHR9YN0/n+U6pQnJQOMCjPghkzt/Bi/A/tYDJeWpFrVsFljqFhZD8hkGmOa
X9jGcIRQcJ15Wxajqsd3fJyD605ljaokv8bCYLuvV2a1sMrPC+me8Th5aQgod45O
FHAZsH94ES1mJ7Qee7lmuT/0g/mIdWErFkwrb1Sx+T76tEj3BLcW20d1LKINfwKL
Frp+zeyiu304xg5O/TbJ1XNRjK4xCrhfQz21lWOQOWyS8q1dqJ/9gG9zd9WXmhbz
0rYuo8TkNPEDI2thSJe50NOxtaTriGZoFY/bg6YWe4rgzBsJJOa4+6+i7wZFaNO3
ioTVWB3nlwHJzPrRttvCVSCrqMa6xVe+4MFL/UJ6yGkxHRRdYgng1oI0yezTebia
tZEB8tL2PEWwImKjWatWyMbkmSm1P/wY9VIlNpnLbXkDBQQqFuqJ7b9d4AaYFjIv
67XvyuwXU0WFkto3Hy7UMnL34LIhCjbRX/IN+lAQApEyRu87e5t/zsC0KZ3hQEUm
vvncWIN7SeOIXlmdwYy2shVh84LMGUQU3UCWqca+U7vRba+//fFMIvvVznDxNfBk
e87WKbdVTNLWhnOYAlyE2NyGD8DL4eOtynlE1mqk4mCOTSHoU23QCBF6IM45moJQ
CGOCEL31p6pQNPVYXGBmqZ/EhEjjfo+zTFG2ZRNo95w9CqClQeF7ZCiccS2OGRVT
AATceaH/PLB2NYkkyjuv1JUiQ4jNKjBqhKteEtZvrY7++HU1jZtZ/FEWDV2wB7ez
wMZ6bYidrl+mGkWxma7Wg3auEeZrwKFUnpegR5m72Ep4kqR5JQlWxY754th0mmoP
uNJcTJ7K6U9Auwf3UOqsjhttkSSJ6dNTAW3DstuhS2N3VmA/KGEJmAvQniqOekqt
z43o3/a6iJv0M2VT0+QN63Y6CARfAPfXCEd3jVRFWGuTNMJ10Jw80fCYLvRFzJDI
uT504KcizTGqe+RjzXFY9ZzOiGfY0sj+UI5zwW32/Lggw9g532SE+iKXSRZyz7kA
GZXXCbfq2NHbdFGuErTt/VZ0FOty5JaQuBGJa8HteB1OWona0TNMgk2yeJy5F5TU
2XK68qWBaWjkjfQXLkuynULumjUzwrGpwvTQrhQ1QnMSkzsII6Zd5Y/bxL9dji3r
NlTy1VvvR1ypPtjZhqyUuuxLDKLDgokrLcVe+rm4KT7TRR/8lkn2F0JTNH1SVYoS
Tt84vI5pPjdht3auTwdrpf4yeN2kMMf9KGUUaGh1te7+r8EH5iBmn+QrYykDTHIq
afMm7xuRKamM5QeD7l9wITfHHBX9FOGZWHXhFh2WpowrHsW/z3Jn5LzX4YwX1NK4
jYRN3FcLUfQD3xV+Ce7RWbb24caxcOMaCu2tHuEPq2CiZsbugLNfPEOEkKwgJOaC
sIEEF90UFFBQXLRkxbtyq1t6ouTKEQjbzhr2HAm4DzRFMLduimPeTOhw1B3Jbnuk
etpHQx8fcVu+AB9TnNeCcUu6njGYqbf5u5nt+Wr+vnGHSORKTUPWR3vKiC+AZRvq
eKgmzO9tfO5VihTzCVO/uu+cM3gKo2FK6jPDPHo8MxCZZUBZexslZDsMTBMmZSYn
wBXJvg9QbA151a1wEdYDDO1/MYrU2B4bNaRumSU2nTzVYCsMQpIOsgqI7DSsC5UR
MTWCGlblR80efdFZEJcLWzDRO88CP96IVtGPVKUYS1TPq2A8xG0vb0sPPIUu4q8y
qT1d4ySnSVERBFRNWe7BxCHs+N1y00rJ0Bju3VZLQBQ/GqElaqT8U7xEDTHoZhOF
O7+6LOi7p0KneDCsFk3iFXho+CVLvZLIvxTE30fQgFkLYPvwJ0ZlatLymEJr3qCM
im370k8uUVpg1G/yqQpGSKEMtgGzhhAN0hFeonTVXy32u48ucrAM/O4rTaEMTfPw
+W2ZXMQQl1xa3SVYQHeLVI/Rv3yJOfBnDf1chaWhjOFvsMY45/NelwWdDDoo1MP3
T/QMzd06pi1L7hIal7QvrGlDEqFzm5+7MgUHq3s8nSC2Z+ywAanaJxO2271JEDty
hlygVwdxXwKt6GNon66TnxNaTWLGL3bN9zcJLuvrdoBJt94E2WsUggVqtNytKFR3
RqXJv7Y2ECYosyirUp+DUmrv4NfYnsp52TVG1/iiAqZsuLjPMyZxxpDXWspxcEZN
VOKE5FBAexgqZAl6xEb4Bpw03hQ9Hc1/A7O2oUAEZzaSH1IZndjqlI28Xq4J9vU7
28u8M1iB6utfLdoePftcMYOLPUESF8x7pxBkJ1Fd0IllHTqv6e7t8+EocEMQNomE
+UovMnKomm69iBd0aylEWwFz7RaXALlo2NOXj0opayKIpY44WOFxXtCDnxJ/RpBj
l/ubE3+zpfcRmEQSDKVX104HaSTWtuRN3AG/1wcQdJKj8O0P7MYzhnFSJbXqT+WU
eS3/bFa+CPqs8tGP+6Q2Fs67wzmAxlHIdXQpzRv6dfgXRQkNogoNIOCRoPVWEuyt
t4sHMN/9VgHM7/rgRn/qY21eXBy0Id8CVoglowD7tgs/sN4w+59DWLBZMzQBFJma
YU3W8p2nibwxa6J+1Zd8ajIhSvK8G4tKqU+sUXz0gX9UtR3wd8VExsi8rIALatHm
licyGszp5M3lifwMutqE0Rdbmj1OkCh7b/w8T0j3bLZjyyPbNyYdpXmNHjzTLpQM
5JlV0IEPpDwpyqUPoY1eC3NUzB1yKwichIcoxDQjK+Dzn2CjMvPhxr0sRwLcIhXv
J1brJUjDch5binJvx5EyjoCQiKfoOIjrNeiq8/ukK4m8BFo1dE3qvXBeJUrt/SI7
rWcJjUYOF4iLVnvPWKp+50Sh4zZgotZB53guZ/+gohSJqYQEr7utVPlHIMOr6xaA
hLpttb14gaKzlJG6v03hpNP9GrTTRXIwrRC+Pe+jYCJwpBb2FWpYMZacCsENtn0R
W/b3Vc9SgA9yoSph2UwlQ6Hmk2H7aDB3I5Fc8asUfnJp9LVzitn/ueBnuNKds1bp
BZxPMAt9st70c8DFA1ZzwB+1Lk1MJi1F9RBZq0kKrm/XLRbWMuEtKOcEqLw1670y
No+XogKnMr6I0/qVEqO2MKA2mmC45SkC4lHbKs6bmACVmPvguye78kxCIqczTfT/
M601IKLl8HQOIGHgsDqXea8hFXrSboT+Js1XoFcZ5iZnUoUCAOtQgjmMdbrntVId
h6NZYFJ9Z0uksWcaw/MZW93lCp3+tCK8/QIHSLLBiK7YBpoR8WAMy799K47tMXce
IdELE38MvqK3gIZvAh7Q/XcZdTj4CWEpGK8Cy0PnSfPbuTHXcl4DRfek2VqW/AJE
YolL0jI0xxgTnuaJxSphuxTEnTn0S7R8Xd7gf4IxTNIr2s5esRcNuNoAdkJlxtVh
2TV5ABDBgOsdkVxGfQCt3vYflqeuN9xZUgZFDZBagEMgwkZK7BCLXC0NUG+wShDb
jbDpSiBd1l0xOp7be1fLgYxi3JF+lEK70SETNJOv7ecJlayrWu/gLjdTF4ND/mP1
BUqWl9gf4NpLGzSRhSQb3Wka/Ee9OdgsfgvXY0pU3LAAgglSVkBxDNFcF7/uqUxB
aQoDAOOketon23v0d1c9cyrClctjASG0e0kOkpGKK7m1YD45t3eV7WmLb/1imC+w
SzjTRXde8TKBo1m8HjgJsHqzCW5n1hYIoXJ/6PRDTsxelJq1mqe5FWrG2fImPjKM
RjzYm3/YlJhVBgIZX+WLP6NHImpswnqFsvxESpKQYAkeFPHBrruv2ejY9O+G1WRx
N8/fNjCGpe3fQGqWEXIHncLhx8LxiKRTP0AOWXJU3GqO+tTLS6RptsBhlCN4LBSf
dbQ3vH6F+cTu8dsO4+OOjFL+C6nxO5RNXkCXtvCqs0K00tGRPZO2AW+9MhJ6Xqm+
aaM8ZyytcqPnJNJ4AAvyPZ/cPFMEbThxvCsQzG6CE6+/HD/c+APdhJnzos2g1WyH
MLoRinE0CMHEXXSQNuLg/0Vsf0Ban8u1q59EW1mch8+GKTA5JSeF78UXaLdga5hn
4m6Bp1OMXKyGOLoPUHsmV/rIug8T34Kk8u+EZv6ZwoM0CrQ2a0sUqvryQ4P7ENDS
Au/9y4SrTy6p0cvwXAonaght4LcVQje7dG4awMRfL2UatYo3FSgd3LeFxEPKOhE+
W5VN3EpEoqcHs1s6xz0ug/4/kfbxofvL8G5G79gkj2lkkL9qs6kF9g5dEcO8NGcU
xPYqmt83hnqzJhZmJ4o3F3sNFOk2+IrZUKkiOhT8a4rdRYCA7ijM6AgryRiYQUCO
Yr2ImDQxOsn8IHhQJUjQ1UBomx+IlS46bHJHjdU6yhawd5eu2Eao8DKA48zGWz2h
EMJNo2JMkxdVMaSGHwj9K15TbuZbRmPhWMoom8GD8EbHJMFFLItV5kClWAtbu2t7
4vmMDStr+9rUOkckBLn8WNgZ00FWW7FeLxNzCYUySpWWSTwWoEZobNk63yVSaITl
J5WYGCNMSwSSW2t99cRMGCn3pdwuXWklyDs6HnOSudNv2/dPRy+LHP2E0VCMrW47
/eVjTZnIlXDXi0Rw6gbWxernlMlLHgq5+lggELDi7oMWiSjict9R+042u7zxgQFc
5wghY0CYa1Q3+aE4YSTsETisSr6ZIJjcAUQe8Dz5XD69/qsSp9pJ+g8moQgiuH/i
+ul93jF9AK4izb1HvpzXy78VoAJwmtupwlFm0GA3Mlk0j26TOEyEQUWbPEPHDUZS
w62xUyqa3SdPnczLweOadow59cJJP3odbbXW5eCn2uXV5OWT8alPqQ1zpPQd6baK
LL6BXzo9dqxRbfuoKL9u8FgqYYjcKWTbMk5RHW8GKmFK7BZFjpSdsOBONzn3XncE
ORFGi7sksdysJm1D46SjVaaDU3YUra5NxH5+o50DzMZ5vy2ujwHmzcrfMkftfvAk
S4e5oauvUa6Qq/aN5gAQUR7c/csfBiw7EhbxH5JGrt2rN0dFlZ6gFpwccn5/i8Ze
GB2l81/tBxp59GUzjPLeAtdcuM7l8yLmU4uoLl8SZ3E3eJwRo33v2cauDetN18S/
A+p5pPYx1xIOxOXzsuDzTlTLCVKi7ILPYyQVG8iFyLH86n8kOsaTarDOkzOquvbY
lCaFo8Tp4pXFaKaTwHIqjAFb6oaUEJsSj4wzjQ+Mi4rYmUYUhamY8Mui8QwCoFSo
0sLjOK5ezUAwt2dABa52ggmrrgM8B0W0FMTjqsG/LA/R9U6XTRSe1kt9/MgPBjwk
ngV+pJNtATa1ThH4DC66VRwGTPPIn5uJHL9vw9ZdIVDjrKdLKoMTK+V0sngg+shB
ihHzYsG7kL+gnEa3pG+GD8cMOrbyyxXnerV+KyQwhnqJA6PSIKPg1MM2wOcUOU/o
AjDpJiG9JF0hb8HJ3e9A0kM5ZRAUGfG8Fe/6kERjy3kK139StndC7cvfGaKRewoK
+d+g8HKmc8+So75gMkrAJvj1EmWb5ZgAYRT6PYMM/JQD4yQoYZKdq5CvRbBC2+A8
UZ0J8nw4nfpxmuCTV/2SS7s+5S0nkKDaE8B33mNmQFOOw7WPivYOiDymoKRJxT8G
h6YhPJTSztL/rO6RC6btZCcmzkjWZpbzdCN0O3kjlBbDrs1jKK8cgcxhdv5oNnH5
ekRL1wzQMryTlY9T3NgtVnTvyhYNOZHlXEsh9w+myoGMFP/eqqZBg4Mb+IzSyLjN
EVcrVWi6Jcv3tPph3MwDqi1rRHTcPdApQ/1W1VKTwJymA/x3h9YuCJ3LOzxPPh5C
TYwVjSa77dt29bOVzFI3m16+xjFaEyM4y+hueCsAqrLYg2v2PxSNdIbZAU3hbG+n
kZtP6rBsH/oo4ljArzt9cdP6eAkkM6TZbStJtHqj/RsBB1dKMbLBQPfaoghT80wb
dQTRjTiO6TYqIiDYvlOfVzFDZj6oG+A3ID4hvRwG9JC0HW700EK4df42cuIohmXr
cMQNjTJbjccbJutk2INWe0kkIF2GPm6NGDqXx/ks2GfkSxpAbW4xAlXLPKfE9fYI
qxAmL9UJTzc18QkUK8Ke/wJfe3sGmrjdnRfP6hG7AgF3UFrNUBXPD5VVNnxtymeX
EVOkVAKGKQnUHu26OhxMtWZCX0fprqrH9hrnUz9Uz10NwmJSKHy9gPvpGsW0MHrg
YQH8kxCdXjl8mqWXbJQztuvNBqDpJjSMdAl/KBkCKItfE+eq+kf0rd7I85a5QVkG
BN3DVjpGDgxBzp13WK40bFQ+cMMGpSADA9dEb3P96ZBsZxEIoRH5NlGp25GslWEa
JRolDLrlzkO9MkMG6jpRbIoHVSXX8FR9+uPIr0RJMxXQrh3DqKWd7DdtSwsMBFW4
HNLIlMEhX3VgFAkBEaewQR+e9QGCi5PLqsZ3ExLO7fwJRMcdy4FelKVZJgajk/Fs
/IOZjSAE4eYZ/7T7uRxhDa8BR8qyp5gDDoo2IUzsfde35EYyX31PIVZ7+jEquSgH
X1oHyvKMvjh6yi9lQrB0vuL8ThgANJTrU12vpWDKKZfynEOFMpAYCmO5WmAKD/e0
33O0c9iZ24W9woGqfJuV1puoR2vnJBUZjIk5HQhvf6ZXlg1Enyj76O7eAkw2L4zS
LL6Uhd4+MIVib53mDlQ42RcvcnAfPfFzTib14CQWIxPrR0XdAUqfCqALdYKPjHH5
kg7tW/Bw/bVUbCdDLvTMebGT6mSe7FJYuJtJTZJ09EOluMcHO0d+A0+JAIpYLzL3
zbAUxyZoPpphYB7EZD8h8fdR4BUE5zCXfQRc7BjzJuxUE1fWFBQIOak6ZJmxrs7U
RUhk6az8tBSNJmt1LHrKYJ47yrMrgTA9Zp/THHb61RmZ45nJD+ijhb5NGbn/aocm
OvUlPbS7KxiUdqueJQfYHNFaygDHvHHdW0ju4i9AZvmoOYeSVCdaHlIYwByb3PT5
fgNs01YE/qMT0fTCFOSkXrvVcb1OfXxc5ymKjRH285p7FMQxgVnmJv7V0JOX6Xzp
a+fC+WlxAvslQ5gGgMfa8luxxNanVz6nGKJcAJ3m97pZw9myh6l05NBfE4JywCZN
ciMouuDxGKtTESwu+YrHYZo3x3gXOy52PVTV2fVfsUthkjOSWKjFfQkxpi1w8XPu
cAxP06dxFbzI08iT+d4nuiEdzNzWaqYrB9Dd9sDAkpPxb0z/fTJhfFp+Do0rWfRL
bbwGFi98Zvm274ZQWmRjlObwdMQSMQIzHUIc7hf3rScM5gTdDDJxZ/66vkJ0rjrI
fsPbq+sn/KaDPqVRqhoqyXNc+sPle95LfjhSnWaLfYkS8Fng5KsW95PwdJdinmON
PBzYtwX/pA+qDMk3aqw1BSv7xX7YuJDCpnOLWn45Sn46Meqit1pbhh35hEwAShfb
/80LiMimKLw4P1BJV6fkgsvtVMovN67fjHqTWDV8dKrQD5gvjegpSccOZN/UE245
zU4YmADgtqYCjECgOXevE5whDZRFXXGy/SOWn6Ne26zTdr4cjcTSvaRIF4Z48KW3
Af88fQ7E4/+7gKQUfCBA0WJeczMMh+LFQe4wpnMSNlUuyWaO7rfB+mE93SgeXkUq
//wv0BqsF+eBPzcmgIPRDHDtHreCfFwTQf5GWl7NNOymYweFl9pMfrh/1A0Hl8gy
QrWLxYpJhzlTPDqrTs8XmV/rCJ2/D8X4EnPJgGqqumAnOyn2OBtkiqVQVMXEPAnS
lbYXjzh6hqNkNx9E7XELYQwsl5oYLjCg6tf4dp7OvPFOqdDrHREcaAu9ZtmpBEyY
Kcydrs8z7smuNV75vMyNDQ+8nevDWZbegH5niXtWMk60jLX8f3NV9QLmKhv8iz/3
LDnqTsCaHN8JwpjtpAI59wVYUuAvipa0kvPizQYrZJk1QK1vVsOw0oXOW1aKM4Ux
CGzlSzu04R/24d5XZ4FzJYMGzO/iR5TWlQ7b+F35IbDd8IK3Yo1MXbroqrFbCTiz
3HnrCerRYZIdQ2t4dfj3RUvNY2Kl1Ri2zRvKPsxCfOW+J8SRcjeS/6f/RPX2n1ow
5gbtBAZLfZQv2cJy68xxlzwka6JVnwwWmu565gI26pqsmj+1m/e9oBehnolHzNq4
Wl3pHtdxFcAUSy8aIzDlG/ejUuiliyUmJD3I/K7A9TncusWS3W8X75KDh4PrZvAR
tXqZL8RWsJqxo+30ttaXLdifcnOM4C4hhpFqxxmurE6ZqdZOlgepcu0ERXnMFgAf
FNr9c9AKljYdPjnDjAQpUiKB57OLaJ33L32CMTEhbICAv+5geRqUgh0LaZYSU6db
djldZbaHo+IlLyWZAl9wrOi857pzUYZISrDOFUeboC2aRiLT/bFdP5gkJFb4dLEb
bV8AQA+3Q7mf3nwoSInHrjM7HbxHUI76tOOXmYjMq04GjQRUg4nwqHesQ2CXgQ/e
Sd4uMhRasGogXZVVsvDqj5iCn1af6vCUPAcxppnkznSvWhokIM7fcVr7Jjijtxlo
TMAz35Kun5yx3XbzZKlK34F/iger/thB9N/zytBz3LdXOFOZZRW7Vtnxoxd2Q3bp
TLfx6p2lZyQ9EIABKXCSVJqp25AThT91+Z4MJGb6SljH8uqmv20DKxIqdvEJIbKP
kNImfqyuf/0B2w5lAYiYl7gfQVYUYHV5VpmolJdSgMjizPuaelPs77m/gaU8CQTV
7wci68Kye92wryZ8QXbHcZku75WTCH1Dyfpdbc3y30zJnZ+PdTBUpgGBklgEfaEC
F2PcZooAoXKfEV2h0ox3euMIv/toV19Kw1ezBaFnCPr7OXtfEiUvg4Sk73JuP1ST
gOol/rswHkMvOx8Rr/L8DtjCajjyBN7Uy4TjLup5hcdBz2Qn94tJpKYKcWCx1rKV
Rt/NZMz6ERsZoOXdyJlKlreUBl8DUYC3DCTawhnSr7m+7+2V+cR8HIKswSQr7YUr
pCodfswAXWRRD0LQ1LMWEHWs+7zQlrm3KW3rL18J5wGDvLRhCPiTkLHWUKUsWuB9
YcrGki1dGnuOkBcjYHCJq9AZr1UZUCc7qE1mVtALYqKiFPrv2lYhRb2Lpm9V2PIC
+sLHrht9Cp+4awOMDMthpl8Xo7qKhyjmBW7HmN7Meomr/uhSK7O1AreFy5Ic9ecP
y64V3GnShfVg855mS0NwmZmFhNLk7Kgkk3M48M3PfruESC27zZjw1ggJlRUYgrGL
hVTNIWUSy0rjIWXT2tQssR9NKdaJ9x//7go8tITy0pG+JS0r0Bi0U05BsDKopMA+
l1qpt1mVnpoWu+AlZFHpBHOsEIkwj36HenJRshFmW7k1eJ/uB+lgqtu0E4B9MNgg
zxRAa4o3DjlpG9AzxDvtge2Upkb0g5JBZshIF3dE3BxGhyxuM8baiEJG61pFJ75+
5X17trzhKgiE+fgveTx//S84EnyKOxvqO9Tw6S5XN6eh+Qp+dAKUijOgUinjBiW1
vjZYcG8PFh206mQWv1W3SC73acfBSOxhM7q/5APTampm/UGQnMbdDBgRBxtjwX9f
9CuEKil4pSXMzoqIE9csY+oAmFHXS8O/cRg3ug59vbyKaxq/rhAS9j+oNSWPidnE
VczZ0IU/jAklx5lt92LzSVXkkkYoq/bz/3ebOhgE7fDp+exsHWI1NXvAP0B7iM79
irvT74fr/A+Tb/ZtFmlfZ3HMjvIX6sVOQhD/jh0vp+Vv1zW5UImYBROTcPCpi8UJ
f3q3dDRJtTEy55toxCVXCmoSZRfDZctSLkG4QaVMTYAgYU0azjQuFI83W9z4QlIY
68IVp5nX0AJUc5DduUqO6FZx1AZqYzN/p3U/7P5tM9BOBNEX5N9h5FVceJ6YHXwf
p3W9tplBstpgcrRENq+jds1BVFxDV2fAkJEf94P7w+NIYkUCp9aroDXJVDwc5Jqw
Pm9itIrcvEDkvEkZIyngF7rcDo4UcvSC0O90leiHiWKnJwefgM+yxQk7hvT/pixA
146lShelQIw34C7ws8Yw2u2UvAgHRVJww4BDsgCE1YZ43ITBb86SGWHLkAp5onxC
RToI2QL0F5anXiNLa9BbQS2Lk3bPhG7t839TBpVfRtQVTfwSebNgJdTkC899/MET
cMMVK8lx/kK1TpNZBWPEq0eiRfFMSzp2VI87RxPcmCYSaht1UgNnUhR09UCmrpgo
9gXv7nwy6tqljbB9aTgyIZuu8OEiJxTBumj9dZAOfvcguErNNW9AVubqLT7qgtVo
+R6pIIhvDAZ9sVgmPxZsRXFYfPUlaHPVVUVfxUcmyoYuNLzyHjCL6E0BitU6Ll5v
Brp0mSMcUSnmD7KIjAh+7JA5Ba8JStDCVeu1Ju9LEKe2q4EuykJbU+dDHM/QWXt+
zCKZKqLQU4BwZe5TrbYLuHYt5piwLPfUALp8EBdpIvGaNkKzQzeLs76+MQNbW+dA
W8XjxmhAt6PW2FObLHxKkRTLsXddmlQ68csRdbv+K7wYniB6ONvPoi1/Zuj8MTcK
NsXsxg0ZiVhP1KkKbjwlTjtsDV5eC8xYoX4gAyvtnh6U9nhSroOg9ISI62pDzkoD
B2CKTZgAEHdoDtNFu5e2IMNqYi2tTK6g1R8HAFjqhXrO4Rue3wv+w9mBySdXOEmJ
jjstICV4Di75G1RT09rzEk/MK9AM6yy5E/M3K9v31UCZB+hmwjD+27eXyySg14Ag
cnPbYyzxxdg54SzGi7/LC0glwBt2otLxbObmyWWUCMH+h9hhagqORvZAGfwz4AJT
Gvpk+yjrzB0o9oWhBZJ6kGFdgpv11OXb7NdOsUann0eJF+sQqyf3pXcPCZRiimFX
SXOMa38W8K26y1mwZ5EnEVqZv4+9O1dPtaISxt6YuwVLZ3GpvgOyzY3lQPAOl20w
tIludJ1huym79QBG36XPCdjDoKZv4iW5a9WUh+89/DGYKFnI9WMdeR9L1BW9UQij
XZ0a1xCATMT4fX+zobEsPWjXc1cQ3WD7aokjhiSnFthjntlx/MptzA3pHxXf1BmC
4TrPBSN7Gdw9S7b6uKsPBv6JqkOsOVjxXJu7ih0YhTYtgS0FPpAqsZiEcF2GXIiY
+3N+9RbcWR2dcSbeERvJLYjx56Au+E2oUzzg4ZcMIX71dZ2w8bpEZxqtcIjHiiz7
sMNzTzcMTEycUvCJ5WoWKJ/oa72m7b/XG6zfYBwSVTpGrEKndqFPmx+/RsLmSI7Z
Spb/9Xw1LDhfl81K9caeYrbPERWWGWohdp3xzUHgO0kYf2HuXqHZJT9TlK3ggfll
ZpERLYWHyF15QrkJpfobu0sdm4LjqrPQF5NvM1exWig/o824zAk+EEZWKo2qUyF+
d0oogLwj73eopqOKoeQiTt1XYfyTBUjPtnsTp1qmHTzQXNKVM0bC5mN8664sh4cj
sD1/W1cZVyZiVRjKw/xtV27YMCPmap9bEcx4Rmf3wGtWqUEQf24qDqiY2hmSQm1K
5vK0uw1QqOi9dJ6WzChOdTwLkRAekayzs5/pjOs4Q6nPXpVKaXbggNcoC7oRJ0Ir
NTucLTqCvsYWnv7ROjWxKf1HOiOGonQySwxCwQWgX8RxGdBhIy3rts0wATw9B8+Y
qg7voPreDk4Hvx+UC0Rj3/IRZQV0Vi+p55REX+s+6YuHsgiPqG+ELRyyXU+E3lG9
ElMkGaozTqeSssu1KEQpumbf5WHD53d7dsDu5PZjpKXA/yUJdV8Uh71cRk1aeKP4
50HkUpFT+Wrs3U8xjo5euS4YThU2uTxJUwt7hAezy4ZT9+dc62xZX3Q/LQGjijF1
jrQh37z0VxDYjInhgUAEiZdc/AHstpDoSK6oNdGYk+LsJ0JuTA9TNOP3GRMZ9kjk
7bsc+kp+p/OrNKGmbywo3YrhD14Uhp5Tt1GUbzSJtXaeWLElAfOMpXsE2QvE3IoM
3OSG1rSV9u/m0nkf/twu+jFR9U4rwNCdb2g/Zw1Lic3CwdvS8P0tFoQYAv8Wd9Rr
8g4ZM75167Js6NIJ51VfF+DrzDTypo1YClSt8d/GUirvJVh8ragSnnoS+PoJyUcY
ei7Abc/KOPwmhDPDQW46xxog2zEdt71CiTdsJU1749DLrIis94rT9DUCxKNocy38
lpQQtJtXIOU8erzeWBzPGKK0XTHOU0mIsqrMyAxyRges4aZnp56LJTHN1gKVq36R
Jt18zT/QFwb7RDkxwvh9NtKdnO0Yz9w6bJoRa7cAV2c/1cTqx6z8ctvZq+p9gkxZ
UyVs1hc5DtT3wlqNIqCzbcgKT3MKQPXJIBWTLdZfi0OoWU9mHfHbrBjYqZmET7Z4
fXnQYRwQmva9xmzJuXmxBhQqnBNMSa0pvY8xa09svV1Lfvn8vmqQGoADXqZR3f33
QNiiEmU4oedsGqKSFZsSu/amHC9fvYsmXrFw2Giy9f8ss8pSyiJgI8VSanPx0Lsn
p01yuDLuLBYgT5fT7gUSwaOlnFh79fnHSePyskDV6e7KsbNmycXGNzFg5bJ0vzx/
7Y3UiY4QuINZzOky4vk5XZYjQSBQasK2jRj+pEyvzRh8C6RqB0d660OUmKwnziVM
dFbXEJQG9xr5HH8ycS7ssFxhDGe2TfAh1X4YP370MlUZLGtzxCFILZJbQvaZnCL5
uDPVSEUPhRIcFQdnY5NYBImTKcloSXl+DDtdmFdRKUEoWahrEjHuxAGC2rbn61xN
nOz6SP2hnl9SVC5R6wO05swGIT8dOB0qFCjSGLmRWg7nW01ftvw/Y3aQOuNdG0Wj
LDyLlyOU/i+MF3p8cCRDKv0lvZspwkXh6h4ekBNu/bsembxyKY+kk1y52hPxh8Me
gTuxWvR1c98mZtOiZt9YcQlvQnvngSCVnIPbnFZYAttkQzX41TfhTAS6roV+VYfE
javlgujt2eV+ko3fW0IELPBBbldL05z/HgTgZBgNMMua82/3I3vd3MSHs3i2fkuB
VBzr8FFc4JWGr+ZGU3nPX/56Ziuv67GPWyXK5ApC+HEVnbqmAJlMPIbsZyj9Rcu2
2wcsH7b0KBqO2lSTBwH+Hd6owYFwDU5WkDIReMOQKOwWmSgZeTi8XPr6B0K85M39
Bh0JKaVKsu4s2dAA6LnjaCI22rC0vySoVlH7FUdtX215VDL1CdAHsHW2DqZy5Fjw
a31mxYmopRXuOy1LEnJbjzvL36VjmegaLpT2evlHKOEQhD/xuOt9wnZ5jGKcjufu
MKDk7dv11MPKY7BgxKPibNZmn7UQVFc+eFzyolhHb+kZF6WJDMKFbl8HyyONW2jO
2akeFpAKU8Aff3Fei5dPFLrexSEZRoKmKO7D+TdUWd7VUJnAv2CGvJPTu0n1MV6a
y7BgnsKP63yKiCylESE1JBeESp0Za7Yui5Yzqx1J9wXY0KtDLTyUVc4DCd+/za5N
J1xy+oOCpb1CtedfBst1YqixVpWRqiJD4G5Lk7sOzJob+XwHSymfgASDhxKNyL3j
0nEOX2FejpE+seHkZNtyome+21actPe38i/uAV3cs6O3ZQdtYhXiazamcIyjK3l9
yq/PY8f/KokmDT1JpKRsrBM7AB2oYLT0hS48uCg9MhC+7Qk2jwxLL7W1FDZMP5Es
vJILmVy+r2UsbQxq/Cvct79ft61PYbOwBTHkBwwZfhuHN310jOxTCkFx4GUFxbXp
vGUlLXeiX4LB3AWmGD0Qgz12/PM5kvOsfjaX8O9Gp/ggJRawUSDntAfqnbxj9vbv
4PL4cA/xven/Iccm+EHK4KCWsyhA2qZiyV96rtCEO8bFODDBiXkye5h8m8bxRQzD
TQCJqRpdUBXHh2GYPaaEsxB/X1PzigUH4eXi03i0BEpyNKhq/1OF5aSdqXQfwRda
zZSeyhPdT3YiPtV4egCitdG70A1YrWj9y1XoBaZz08NR71Nfd3e5ojf/xH+YHNVn
JXARdPKiO/A1NQqDUaDFO6NlAiAeYCJUjwKyBFwTiUzpRE3EbFe4YO1V1wl2ZjWZ
T8gNInzzV36GAOJy1y2La/yVb5sHCjZqqMMQyRefLhIZfoVNHYJOK2UfJBTvz3Lk
s1y50yVkkjGFHIJQEB4L1H8EvBgPh6940tz9oIzlJWm6hSlwe9hyuO5ZHKFR/ajq
G2vacA2HT/H6bftFpE1CggLhIAWd7NXVFB7vyxwin4K+PRYKd2IMd/SHmQafId4v
cX1sUYcF3kIXOKhynFUhXl9/1jMFQPLHo05uzSRgS+klgGAsbFqFQCXVw/eFx0fI
AgGbpIp5lICQkntoYZiMIDZV0x9DDQqgWEWnTItgOdkOAtqR1n2dapEthAfh76An
6FWwhDncYQnR2NMj+cFBzofar1ojBse5H+3h8JcbcrgzE+ZsXfs2l1fMXxT+y90t
MkWTvYwPgyN1Qy8mhKYkrL59cSk5SOTsbs2feK8bF1HTj/EyGH9/o6y+asnGe0/s
E7IOIrfPknN1YjmrkeSIUXUv0USBz4+zit/TlzwRXDZF1QgRXANPt9IQllUtRChK
2pTl0UP1dlOVfbxOTyA12bKFrIzR7CWnTboTtkUXVjUOHYGA7kjSwx0GDP7zYswz
b1RVh0OED9qfLkuqeD8/ZCdbA5PsMc2WYk2Iz7N7rRT9O1YCgWtea0q1HRw112b6
qh/BXFlT0MluCMAyU4jqKBS5hYzSZaprhtpsjATKCLD+yJ4YCvvUlKrVPFEHuidk
I1Z8n/n8VZtBT0kz1k8faf13YDZrSScIPzfxry+v9dzMqgaB4m/+yQ53bQ70p90G
M/Q9RSoHCJu8HvF+mLnpp4D4KIjbTdb2RRDcJbwy1+GSKrnvdKYlBjWakV1g+JXN
FTY5wnkFRrnNey6S2R0x2rkXXXnzRneSRbTXjKJYdojFhfhn4EBp7Mni0bZcnIpx
yS0hDePM1UlU1lk5FFYiyuct4u4TDye6RszxSJw3/mGXY7pFqXEvdopw5HRnZ7mC
sE4Lw3FP6eVlLJzy5U7EpqGNc46J8SL/MP7N+EPdXCFiXrqWFkZTrQutSMEx09wq
sh5myIJx5hKs6zcFhKziLpWgaOv0Ot3dg2Uc6yIpxRIL9XDfeqgqidOpOiTixmFZ
BvjxqSGM9aIyrIRhwi9mCrg5gFhityqOTwfb5u7bZrCceIuFGaPnZ1yZ/DQQ6HdX
kroJF6BRk8GH3o+ZEBVXJumWqoDOzTzeR2TJaAM36kH2HLMBMU3rKCwovqBSG+7B
gaSiUVilq2UPjfvebfvivMyEfj3oJ4tIDHnNuIFzFQRap+skwry47HPX21Hq7FUT
k0zdVEnbwAfXo1otmBKNDGuGDSLsazUco5ab2V8CxzL1velJok7OHg+lcyYk0z4T
vGHAzLHFzZMu9180YeXdqWHO4yT/Ac/gQ/H16t6P8/zX3MtoRksJ1tzJW3FlBzli
6hHe3o4x2WqRC3XnQHvbHyLxxbQEjuCdpiOr5Bb88SgckkqD5is8cJFuYBDwRnvA
yq5O0mbHgr1XAz2P+Ep88hnyhtBsQ6EFYZimSEmMYDXv6M7TTQM2RB9t3jag9Zu0
m+Qks2WQCUGeQVBvT8ur2sBtzI3CTIas5FMyfdJSBwCY0PNbRBe07gKnUqvfg4w6
z7tphsZw6Do6bW+yoJ4REGiLH00RgUv9iw2rmAZY1jP6bicNvUk/9PgIwyEwyPm/
iQj1arY7ML0m0NB8OIg0ysXhpsWcSkjt134sNyQZeMnScLrG+XdznRUm4dAE+Adq
eH2T31IsbZ4s5ZwyWFp5vBSKXhdf6LDElMZJyaSbjmoQJiF/5EHxPUmkY6pwV1DA
BvuZd8LTs48dF/3mqGLoH/llJi3rFEs7T89cqMyBwXRLotAMQ/9i2ODnrK5DzR74
HHjkzoEVsEZyH5I3m0CTJh57x7fmMjf3gMKzRSvqB7t7NeYpsG38Py4wLCVwoGQv
vAXGPjlHNsb7qNdVs1ANz5T7j+PUmNQb3UgAz46uaswcljviQL8wAAx5wDSIiRlr
gUeYulxAr32RA0K3Hi8j8dxpWcWMhPi3oYO6lmm//C4CCssZmTSHY2Pcqd7vbSKo
0T7odQNB7Kkflu577DS88Q5ArNgXbQWc71uR6g4zx6LAutCiirn7vymNgo2m25Gg
Qz2FXRNNaMDuu95qnRwcwIbFwKFYMVGglZn48myMJvb812Jws0qrJ1k0i4iZ/JNM
DjEb7+NQbq1dlISPBXONCn7beRsNGEBP4hny5evbGkBWWbEtanD4NI8F12avhDmp
8IUR4+SK9hvSE86rN351krI2sSz6ObFktxi721Cx7mCEteSvE41otnbIf/bqfEIX
87CMnzpJ6FHLZ704HaC1ZSaBybBd2+HFip+FSDxXWefNAj5phXZpuRjgUk7ZoFOF
f2EGvcOYK2jvnhSw764q5DrajP5TV1/KThbIsaVhHMHRhWsJMsuxrCtXrB+VaSdG
+kkX0gxoeZUWPYI308TQnRoDJ7KZ3qR6lDBwEANQ0geJNsUYLeczpG/OXwY0lT+F
7RlcL2BEugNGmSLbhCSnmTOE2wL7O9TeuLDM+37bs3RcAvEAZGVUsxuHH0uOHgAp
VXfcQjXQv5lBmj6vy9OogSTe81e+95w6P72ENB/hFfzhx9nGoWXQrIS1WRBT/z3h
Ry56cfbC6ToRv4ChM/J7NTGOXsyhmx47h5tVjdwtIP+3iToY8aoSgnD7jnaynRTZ
V3/tpmdjZOO3L8qvWxlqTuGCMGcTVPnh4xFvGS6U6tV2PdLQYl3zdBe0PTfX4F7D
2le4b6LqVMSZaZzwW1QnWHZVx8Ca/0AKp/mBvc03KvgCcsoIPWm/guCnzi+qya3m
g64SLOkgI7WmvRV0oBGb8i8XjWjSSuxxd7FFI/uQfXfEP2dGL/onR8VuVS81H9LZ
RO2Xac926UBZdkR8KR1HGhX7BHMLwYJ7kcuAbldswuH1eh9UQJpCl94yzVJSJrfz
Wktj1XbaLcFnCPuEHAk+jSO3SRM/xLpZkdmpASEBP5u4g+O3fKnOzZBqmCh8Bo20
8Sdjgb5u62+1iazT+v1UfI4NsKPL2ZO1l5FK16IpTO9YGQIh5AHdRdlG5wAyeQRH
Dovd9hwrATQZdRO0ioULoVzEn3RjczJizc5vNPVjW1Z/JEGHQMNDtvCGaowpp052
2P5yKjwhF9isALI09bBED3mWKh6JVOehlZgjoX3sy3P7v2TZvbMhEhucq3kqajcu
mSsJFtW8oR9imfgB3dny1opsYV2vVLMzqCDnQThee5Fo42FZbpt6C6pTOue/hTyW
g98am5zrqRaPJng1wvqmS9DavMV6N3sgn+1YeJhpjBtK/dNwsStpnrjAi54lSswH
PGdZwYoBbMqFEuSjMFBQsd+f+yXyyVh8l2v9hLRjEWfX2gK9ytrYefJErlcs+tcI
V3Nwi3UJOg06+egMXVHZAKxBPiCvgzect0FR/vkG9lGEHNiUA3ht9UgA7JdVfB5E
QvKENB6+4H8waNnxkalJMrvCgwdOy6w33Djv/7WNyqECUB2W9AQf2r/rPRZNg8g8
rqqGNM53rQ/7LjE3fxBkdP3BRTMsyqxS8a9l/CsbcatHSnZyyo6S8EPuQn2hSTaH
NHbu8sS1GYRbx3ZhfNk4EdWucaxyTpadweJs9V5EHzfDVVItgolTbqq8I80sj0tH
HRz9gKmQs/9P/Qu/3CRhbAfmJhL8z4frDrVPXVzxL56Q0UzMjN03zKps8h6Y4yBB
24HASTQimrSiTlE7eBgNBVtaTxsdaWUugCRJIh7nnlLVBGgihCqNRQFCeoJ2l/hV
syTPyH08gF5uVoyP41lcNmL4qbArSqljvkPHiPwznPOa91XZttxpy3T9T6t0LIq4
PXXKXBv/QOKdRtu4lm6KyOK8FKyL4y1fSMcX/B2Dk/wB8uVQ+h2Nc9oCY0QT26nJ
6fwntDIQ4gwJcSDm7iQ0B13kFqhnSWvX4Luf+zD4nKejuvdio+turdEipMJg5J3q
QKiXhdVTwbk5w1iipgBSzC388TyiCyID1Vb/Gm9TZNrYFpV5/bPh2nGT8F78m+nU
BUGbYKvjJLIlVFbVdOn+QT3SUxZwxY35s73tpigtRhKJ58rGB3CyL77JZk9ydDU4
Mk0twvS4/J5Mrm2oUi7OcJQ6nvoDFxWoaWIBhQad2Iy+h4Pux1ibl+7/4wqj4jVS
b1RP+T1TZTNyiR28XsxwxB7j5buk8RVPAjB7TTNaFlfPuRgqIoMWONuMEbnR8TGy
Dn8LTwa9JG2/mMxvPcF7wbSyt26rH9tz/o9t/xhMIK3w9y1dywf9ruNte9cN7/Hb
2Lnx9ejCUuXSRCT1iWNJCuUIqJ3hQgyOrvAY7lfC4ldbOqt5yW9fo2ojN0xac17I
5y1LoCk0WtQ0PJWjcN1Ylt881deaS37u6Xnuw6trd+n8lYdcVgiW5t+3YBxkjlr0
x5yN2IzHEp4kJai3+whuJr2n95hrUlWGLA75wcXPjyQQPPQ7ScdphF1kpvnyGrda
GQVqSowvnrqjTp9C8UTtiCTuECvs/ezGo95BgJ0koaugRmZCBTZtYMLzfcGpytZT
HMkXtoNLKaNdaF122AL8ZO8CsIkL7qdA1phtQ6E+7jxl2Azz4m2Tc1mglYYy3X3K
y+voyFnLkH+Y0UgsmCembcwbxdISU3LQxCmjIbHVbxfs4RY/xnHWegg/mNEnEFNB
OB0cPnqn4zObkgrDFWTcni6aMBWlPt5KskPNO/HmS2xr7ywl5bPZaY9Gx5PPqPn8
oI52n0jSfYDB16+00f+9wa38WVzBCFIffT4nuZ93vXb2+yj9xRonF0G+BEf9M45I
rtDpJpp8OmHYvbQKBHyYj2apF7F7i9qPs+LJVhfKjs0hU+1zC7f7e3S5q8ZScVnb
MfM84OBv5oajLSA3uUDh9zlyXmvmzcg1GUub/egcoVuW7fJJPKSLgL0AtH5Eer+I
+aqNXq8xutKXe6PW4hfOov7d5BfSAPFBo3lGZ48nViJuEvJMdqtKjopGwoQsbasw
Ph1qB2FrNc8fPIQEskp46ucEjTts2V6+t65Sr2Qr5Mn0GHB5zDFMLDwv2mV1N063
MoVpnIpTaLL4UAm838qSspdDzg+E7KI7STK2lyakaRTjCM8uHaTSFzxzHyMGO+zu
TrmB4yhZ2grMuMlw8gUyHPiMdyeuT5brqW8Rdlhdwmhw/T7OnZrTAV3ywLL4QZWh
H6+tUzk6A+themF6o3H0sGMv/SBCWsExUwAYDI6zqek8Io2nrACCETRhaZF2aAEE
oetXe9t6z39mscbr4jas5tvFnajtfVtsWaoOMtRtUalvx9hnB4Dni/LyDFhMiaJZ
Uov1JgTcTn9e7D2+RRuGx4FEE0PPC132OwfJ6ci9vwV/XtcGK9xrnvm//K6IE4KD
X1fPlVi3MzUpkETVbJQm2kde39SrynAHNMm18Dc6jPn/8BjNep61JhdZZQe7TSUN
AQS9fJp6tCRBdavrl0S8k/hH8kKwxpKcuqZ8IU+ey3U4mA9/rIEtqwnLJRgPKLhU
XXjdcQfNntFrzMhnh6eEC+5ghiuaHIR3Mmg4ef0ydbDc4Jiro3cWt5Nvpt33QwYs
QkzGvjUIc8dHstbUhMs04ldsi6GZGHzQvJlRRNN4f7bZBaE1TysmrDnKm0aBPx82
+UFavpytV8VIlh+Cl+Fd9QD/meFjFJ5RJ0wuxvmyi0mHdMwEskNto8WjI8ljKMVT
+OetiASZ1q+2L1IzhtsOjd6KpsglkfJMITJkg1VtkkLsEL/BkQ1rISQRAIcFQveX
gOKPqxlJ5hRyGMJwVtzytULainLmZEnUN/SxndvgPiEtRsn7yE0FYRt/rmG7xQK1
Gf3sqamBgsSPZbAZ0c/Tr5NJgwQhCeeQ/PpkU9FHs4YFJtUk7JP6k19VaSjyCIYx
UihYJ1UjGyCJBR7umBcI2nX4f/WPRqGYwOlarrZ7IXl4SW6ZRDdcHaHvMQsLXb+g
AJh41BKQMYBJ7Q9tja7NhOJfLxNf4yYG6c5jc3n2k1PTQC0hJE21c7Z3VUlPdAua
nosSr8bun4UwTEWILSsBXITJLoHJM/GnWpEsMJ6lGwnDLudkQhNLtUQ3ESb7WHB4
VKzrNUV/YMoZNftGMVc7S6y6qQNsN9/RtqmS38mtslrA2WDTIgZqKT0T/oN8P+pw
w87VmB/kXs+QfJVSkWl37PFZMc5DgtJph1xOwnwiZLRzEvm4OK4SmDvmQfxQ5Qjo
bZslm78oMLJXMQ4fyu0ZVx5zBw1RgPmpc7oUzUoBQCSjsFlDvc6UZUOnp7u2cdLf
H4VTAZJJt6ChpRBo+Lbe5jWjI0xw5a8wKsZF4PnJQ2LjPmKsYWTgd7Ad7vfedvAc
/UPTxkqukpHXYYN+4+AYgAsoTBb1qLTOGuh7iGUEboG/bh/6Nu3MgEEaIvwj5r+8
bsmvBC2bEfOEXny9gL97mNlJRMadbuRVGo4ymm5hCaDg4WrF5y4QC1QRS4bQ06Pl
o7sD4iid122J10dg9fWn/GGmvdBWPiaQ1tsS/5rdNGK8TNNht6tbXAWO8iNhp+qO
Tr6bfDYKnfanp2PQp2T+QytHfLf0WDwccZ/rOzs+RQXZEOOiMQTQSKy0eRtTmIyW
teHTiqy2p6hD+ULgD6oxkMMQqSl6pbbwuPcdZPuH0Amjiq2NDYp8GM6hDofx5+um
lgxESFwuWrBWM7fRRI2xGyYIKJIrkAtsmnaFkXhOxwsQms1vSc4f8ZGaJjaxazLT
xED1Bg/iCVzyt35RnxXcN+ee9J345/IUuSL66/qqHC8Tj0k6M8WJTTEhxHaIu08s
aLFKXFUDF1+A7tkLQgp5Vs3AmRhxvtggj9738x488wtkbt5yvU6/gVkY4RZl61yy
AOR8PwK9POEupCtnBCkksx/ePlTnJt+Rmcl6yGyA7mRNtWHwMdjZc9r0muLQo6Tt
2lyJixTTHYePmpLUXcVIdFp8XJo64YLO2sQVpHcOPpcxlcLXrwm0m/pz16DwLWGi
SrndD53n8jv5f8HTzdyeoV4aAQWUu11jJC33mKPIEn6+kUX+HT+aElNvtYIgDGJv
GEdUntexUGLK0pu33onjhl1QKwhJhVJpZVGIVpS9fP/stGo1JnJyGLIu8uE5Uu7p
2K5QRcBK7x0Emv+ZVu7SaWOq7nQF4cx+iYqPmmCtjWSMxUvtwFMesY4sI9qzTu4K
6ylPHMxMNwFLVdZh3a1ipxNqZ73ka44LLVY9REBM8D4XtO2O0PAN4aus5Ki08yc7
EVqJFSQ3LhtyPT/8Q1GLaOkJh/sWzs6M92S+R+pwyXVhwlhLAsr6ruvx+0mFeu9K
pVfQVG6bXD8tWq4R5QbZpUYgW6Y0cIlZnZnbvBqJJXtBsIJoo+Rmpjwsro4wxUMZ
zf0D0QI1V8v6IbIW4A5gX79JOs96HWPLpVlcp9sssdAXSTdxHiSkpuTaAppzbAym
EFhPlWy3kjFR9WwETAdQm4ajTKH5MVS3VmsAAoKdn2EIG/62LSLYukpEjqoU1tW3
IOzoSE3h3vUSmAOWiB9s5PINMxwN0S2uoFmc1mpVO+cHyAxHDMZFVBykY3HNwdIF
C7/fB/8mwpA79jy3Pzl02sPihD+zL74jP9ug0AZz8U9ADDU6N35a5YBvYVx9rM34
T4y52NU8G1/CyWAQxvXDuuQ7KfdN0mp1uQvY2VUYb5gxp7hhLlE2SBf4bf0KPEPl
zBs/q+GFo3yfXlVBI4NmY8ri2i8lUJLgwFqvJ7jZBOpjFRCw3h7BhlkaKFR7c6Lv
//jeLjJRskWh/kjep08i62dUjwGW4LOYW6NVhLVgcZVrHIDlAM0AA/m5fx/J3Krb
XwBLmFJBzrGd23kFY6pY1K7+VGLGUK56QVfUYRB+CHQ9s5KcOTrnyY+UOcapZRZv
A4EPfRKnKDuGGuJ9UiOP6KBsu5RYRW3a/ZD2F+r+CtxLXp24QnOnuCyy3JT4fFeB
iDrcr8jBk3+Kkt5NKnKABJrKAYzjuVSsd7b9ClXubMUNPwa2WsjiWeewXKfboihM
dLrA7kK8h32TnkUTgD/BJxNjrqlcD+trSGwGBewOxQNbi3KaY7TCcq+cRLMX9xMk
S2TAMG6d4EWbdSpV/8IXe95efpoDakjN0B9Ad8Q/GPw9yHmkexrGngLY3VSbKKI0
qKVEelITXSYR6ha6TgyoBulgiG/kD5H8xqNQ1VUUBSbCQBVG0M8Et5T4nSDzN45j
J9lxLU8k681m3682pt9VLpqEha+NjdJMcH/s4ww4hDPR/hLnZ2rZSImFvteNXztl
q8wNOfxq0I7K0itQ8Hv53s/UQyJOT2hljDXGw0L+7taCRs3B66dDFkZg62bajGtD
0zIsMY7zrE/t9xukPkbrA5n6fNn3ggXDZ8UdV1WpeGYBk3zSTzz+m0oLWwCfDnUU
1Fq/McT0Ceff4oko1hi+ctCkk195EyKk+7DM0OoXrPtD3w5UfhrzULdu1ckXBDpA
zU6igraAH0/1icSXVdriod+Zq0gz1IvdZXnHYH0ecBBMF/PVl/x10sxwI8tKpgQ8
IH1vE3EfdZzxZ1yQrEd5tGghZzR1YocYekeny7Wi/H7BhI12N3uIZ9hv2WmHlsZR
KWnaohUUfj5DbQtvKDVRMjxifB3gz4IWquJtpmqvFqRLn/sdQ2pEPbGrDpmwWCXA
gcTWIw4YhkXcWcHyMXG5qVmQTfag//VcxuGacArm14y2LyBdlv/JMJvg9hEhiQmy
EBhwKbbQmZWFPEyokhl6feuMq9gB2gcZ1fZ/IW8uo+7h18SftQ15EpSplLbaeJnc
6cRTorvPiTneZQcuGM2GTqza16Y/lKLI6MeC5L8pe6YaXLHJBXX/l68VM23/ETo9
bnABBwIUFVGRNcDHPcnlbMAhK2bw7Ty54Fc0dE+wXDapmVhBqla/DITRLtELDuHJ
gz5DGXVpeifLAtWuNKLuXPS38yqrGGONmY7lAj0vJH1VKAfykitfH3S8E0ce95qK
+uY8HopqgYI7WRWp4BjdOYipBWIfpo9MOryjUhiZInl1izGiKh6FyKehaTSyZQA8
/FGfU99Eor2PptpKJ8dEulau6DqxFbWOZ66cDPqv/x13YpKNaqtaz2+FF8J6g8zi
NZydUufjQui2sN5wkAdI8l/FqEkZAu8mIaVEIPBWpLXJMGDqWUivmrLuUxFuSifh
5iHt0nKInfwfRAtZJRcX+f8z2s8eYQb1nYgBnBHOcodl36KKP+dLVM5nZ0VY3Qwx
WuDYPjgDswk5w7EtZ5piumZWDHMtvKXeZy5oUtifBv9Nm/UMme2oObeu1pCL8psr
4ZIQ156yyGbW5qu//ETRlR48lPu+VbKnYUJt5KyTgaan6qhESXS4CtofA6Y9ksn/
a7Hbrnikgybn0yM9g6pQ8J7TZ+w9pRi1K5A4sVgBYCrJeFX6lNPRimARwfWJB7HJ
QRNfHW1hi7NdQkVNKnxmqKaplms2+0zyfCGqc+b7+N+Mm4JJofMf/t2SkjK8L/fM
WMyDTlYjv3oCk2trDNjpBXgfg0AIaGX3EDH6k2JSt6Z1z0PNvo60oooUdFDoI78d
a2S+Y9+XZSZWyK0F7wSpKN4NhwqqhAYFolHjQQVKkZHXmcq9vs/ziSlDIbXx+0Yw
fcubmrC0RLDK1wAcuIJZsgW1rsNY7phQfWhBmw4YXjhv1hriLiBTwCmxv4w5Af/M
b6fVZOWJU3OR/qi9eIomfPZZwTCMmZYp2wFzSlYwwBPJljnaAKoiN4zNCaZ/rsPa
qpKrP16tDVfAj3udxGWcs3JTXKjr+FTpfgSMiLZVtxRbyt0xNkPBUCXzf0T8XBpb
lRTB0/2koHyL4yu0Okg69ZXDtZpAuyufp6nVuuoQntxISquFbFl7WX+ieBiIPOEU
vCGfB7VdX3HJbCjAESBXp+bMZ5otCgS6+cYtiQN0l8nn1C4YvPwpZvBvhi/sh0ln
rzQUVCinskG7Cs1cXVfG9TMLA7KqjVENU0w6St8lhzcDj3BlmyR/nfBGycDyZzIy
M5izYU19v5OpQCshxY9G31bu3nPuJ76hucoSFgZQguICiNpZDXHQDWnhsbebq9/J
3FTIIBTBYbcvG+KzxVyJGHZNyI/DkPnoLyrwYDXjKM8+tmFDxuY8BcZNPKaki3nN
0MK/bAUkHK7W5G5S/TndRTZW7Dqrisn9XVrF1sdPtkFL06Kj5eZL/XVJpuP15T7f
p8JGIfFImoWiV+W/vPeHTvznwFlfZBdtBr1HRLW8h782xbW8eoKC/EDtwBxjSVqh
hOTOf+wa4DGCm72DLDD9UcEABGAQj724fSObafmhHcgfjVsGDJ396Og1Ffw93iH1
2R3f1M3C/VougEXKAx/zhpiScczZdUCHZC+ABVEI2n27TOQztWyKezAAAnf3uwuG
3fTnyC5+xymHl05w3Eb5CH0WbNvVD0D4J3QtWdzHglO+KYgHAO3IVPz4fRb3YDKQ
HTFWQKF5MJQMWfdnq1SVLrnEZ+wjghMq5xB3csjZzwJOg4XIVNSu+s4TOnNDBzfA
LptT8jRQJLnndHN9K3PZdVGaZT1hBP2rTjDZXzquvuzfJ8pHOf+k/LYO8Q9KPg+Z
dqkBJFUgFU1gLZI5ATYYyOUE4tLf8MG8S7s5cah6lJWmn4z0WZv5s5s9a0vTDIxC
f2Up0WKNX18s7QhlHE/cV5FloF1wUox3iBOAGjS7euaQFl86HX1o084KyjcuiPVH
6Doy3LH+UCSV7PvPyhW6pA1KZTRMwLn4LTpkcAyFJN0c10vx3spDI5CIjh9T0i5X
STpKdOj5UUChKxohu420q3UJtDtxPB6gX/PgPPpVQibrBYUXs/mU1BdErdNaJAtB
k6k0fevy3FlbuPhpKBVr2gcsJa9XJujQL6tnmg00tGyWFJ7c8U0uPWbJ9jGYtc38
MzHfYxaX6Yc0NYtyb17ipzapx8JEJvGrVB9K6ufNoHnzB+oZdsxWvF9kjQ3JpDmv
Asz+HI4h6eKuMn6LlQZidA0PYr86dodvImwObZQiNmCnjLdkRDR8ptq6tPSYD7c+
4pby6lnbhn/opbH4W5aPlimHVQTD9NbJ7RpvIwF1TwdOiodI1dCIYLCDGsUXCLIH
kKnAoItsnf+NH13gtCMt6I6uuUjnnSiYHMqXY/P00/4StAUFiTGseByBchLwn0az
DGBvN3HfW3esR7lHKsvf+Psad4+qrnVysJPZIY4pOh7dbket+jtSbSFcHkMdf4Mz
JkhCAtGMS4wroDwzk4e80baF+pdzeMy6VzrQUZ8va+7wxdSvsTXtRXNonoQDTYWE
6JkOI2CZ6cab4xJviqGeUb+md9H8IPC3C+yyBlZHEaQrYeiehvnWi9ej2arYbBg4
3+a0PTLw5r1Iwrfyr9WadNYD096unFAeSSroog587BWOiQjPqrQeMntx5a3tL1JR
s6tBT9nr3qDcW09vaw1M+FrmB/u+ZYNceurs2E4i4zAyzTXnYo22pXtzUuG/N2EK
Ngq73Z3Jfe+9NAGpJlgeKCUeCUTsHo8aRt5F7zZ/cFJAp/+O4XRczBdUxtH9OAgr
XhQTX+w8iBVrEoI0xnFM609pK2Q1VKe5guJC+f0tWHzJdHFdrpKLYk1Msr8qpasa
ZYkk+BiIz7Bk2JuyiVoFIFCxD26J2uGjIzgf016u4qbmaLEq6+npzvDodg2r4rlt
5c/tjI5mIzv1Y0FDfF2hItA3DVp/OvqPKfR+RzvVasQmhEPV7I14LT8O71oxw5k6
Y2GC6JeGJegrVNZ2nrMgBEULxJes1XjZ5Z0SXjFtREu+WwsTvMh2kcOiZh/7wqXq
D4omZeyZPcrwcMe30a19br/5wbSgj8WAvrciMCSUePqAZGTfEN+FypfBYKLZ7ChE
19372qQ0ub1rwdJs8SFPK+zeNIYd9WrW+DDN6XNuN9zCmAmolLgaqVt4YVuJ/MmX
sv6NEXaO0Y2GY1szC+QcDdjTdfqx6e8V3XNtD+/vORlo06b3tMJT9DsA+NiGJp3s
JQ6j7Zjv5SOGy6tdRzKX5Ejuzk5DYH4J3WWG2k2/ISHn/aBi+D2CyYupMTNE4Nhk
moJR53F13j+EnQd3uyvDLyiWHLpCMNBoOHYRgwqJ9d42DzUCWXifeZ5VkFWa4PjF
xTg3Fqo+P0LH6CxS+C7uUbS6AMDoCtdrmEhNU8q1QGYO7L/2bxTMR0MQncQWwMDp
ww7LObDtaDI4vI97vqHoBYjK7h2aZGBXlf5kM4jTT6hq68LxNAFCn3sMRvWZKHrx
Q9Bq8An3fVtplZl1lapQMw+7X39kZvyXnHIPtHnw+gwy3m93Mm8mV4S65ySlmkHA
dK5BHxyUrPz1QG7EGOFK9e4y07AZdirrvEwp0J3kTkeyXeaStKsRhnrszrs9WQkx
+IZd2xO5m4zK7CxugSHMyXmqGlVYY4+ahaehF12CF/hYa5XbZxlyl8gcdaPFfvcg
ZtI6fkwhNlsukWgq5W9Eh+jVOmguyadPUIZKT2/EJDP+Nd1HxtDOS1jEeRrE7Tmy
EW7NYapGb8NDKXgfHmhOeml1qmzfmm7qK4D5ZMmU7UBZBMx9rqkSIHEmszyBsWc4
nl3eiqu9sZxb2DusqYT/cS60SlT39kktdvJnK7DqEinEegIWBdkcXgxXwpwxHFk4
V5MKEF/Ja3WNLU1gr+7emam/2zQ+Vw02InReHvr6nkBtgq2pXfx42c4qU9IMJjrl
xYSUpTh3D02kLlZ987xAq+NUE4WlXkZ490TTEzNB7z7TXwiwWMApml3vpf8sMyD1
aLL7i754+WOK8e1DtzcB4/0MY356yhMY7m4I930niSmV9md0nfAzv+h50vxd2tFU
VfoDJnd4O76BLfZVYJz3N6Ww7Bxj+G4R9Q/nSnt1kq7Zf8s0cHyhA3o0tNECQ7gZ
OnEabh5Ma09UzI/SO8cXqwygIRNlL+oIutFSsAGVFIxmofjt1PesGTzKUwOnJFpK
TXlCEwkdcfjPD/kkuXZJ8oyNwfWkkL/PS08XaLwZf51RR4XXCXUS5gKLVPB/qn02
vLjxbo4Byh+cHn7toCfX3JwcR9GhBn/FqXR6EYsRkry3aUcSeLJ3woJEoMwmktXK
Uix552AeOdT2GAb/IxhyyGS6tCkFC4vGTf0j2qHJAq0p+6x11x3WjywlETV+Te5y
r/NaNBK0jKGL6HSV9ajdmBgGVLWs2Uo5REM5SbHC6Hm+zeLwbGARzB/60UqOSDeN
o+PRsUl4RBwbFki/IpL10GlM0fTHwgxPkdS9wRjboIypT1p0Qib9UJjs6rKouXPW
aJ0yDgaI4TAtinzJEya+drrEnePmMFIt5cD+I/PqAt4dlSrc4R5t6NGlX2+633rY
2BWa3k2JF9cGxyBOdQGfyfphqzIK2vIvNYG8gEPGjgZIsGpMNhSfy6WVBTicAgtQ
KO1/azxLGk9elBGLVrMEROylSHKaGLAdU1WxO8FgEYe5SkWpNkXFFnYqyOAS5rts
aiw3tA4rwuPt0BYysIVXUpPKhAVHxYHKtTSOkW9NkmiU5QdO4M3shogd+1691AbM
d7KYoHP7MZ8ZdaTLangrenFRUpNzKwkBYuJ8sPgEyf//C0EygHGesO6qvpdyw05h
FQPx4GkpyYYznBxKGY/xSu1VKxUW94/h6j7pOXtXIJPH0hxr4FkzFJ3BkkLVK5wF
/nzDx5dXWOcjMhuGVGOnwCegwyqlmVL+fFj4z8beklK+/qnQ7Ohij6HKTwqFiRjo
JiRKP5c71oKIa0s7X1Xpi+7GyvOtJF5cL0KNt/VYzUA64xASSPwT9P2VrU/zbu96
tilzDMXSR6UuUQq/Dzbw3f28laH7R9pdN7B0mQZ1hVLX5CKDxH/H3MsllUqkepbT
yanOM0scGCCu3DK6UOppCqiNCBivqWRB4Mxu0m2jWOH78dvAiIs/HC1MgGAbk77b
Z3NHVwmHx+Nl4UkqZzJ81MGEUla6InXS0rO3PtlgdA7E6x1hiZQCdAJLgpILe26e
IoPBZEeaNBmeEkrtQZOpoodr2wXF/OlWuBqTlDuucKEjvYA8GYkx5JvaNP+VEMGM
3xM7hy/uT69K9T8uty/Ulo5XftuW9Rqj9/PAFeuUGWPOMePHtvkxknXz7s+Gf51K
sn9Gj6m+xDVzIASn0etBLpbf/DRWRI8/gSotZzSrMnb83KiVIHaDkXlJKyeStu/e
Oy/0jflUIA0KQ+ojn7SgaAk+3t22ci6oE78LLR49qA53K5s6u3Lazv1esu5VN4io
A/+H/J5YQeK9fKHt3BiMQurGSMym1JvQFsJhJFEZ8kg+RB68CLxqKvmb37h42Kgh
NVjDVgB1JGJWqHHneCcVLAusZvSZlPKSc1gtfwCakuOlDolTSxZWpnbceyEvvP82
zMIJfwYdfF7qvx4sO2w0Jf+jpsmEnhV/52vSRS7Jxk9+TpbfCGoJXfjVg8ClwTIC
GqbelbVuXFKGoYcFoBpBnW8u3v6RrAgFEdE629KERFqSyEVIG0cKy7U3fZAV9Mv7
5DpZDtY31YNwa07VRhI7mabSIrVtbUuuJVlrU1oUU56tE0VTaQnqZPIm0uCxXIbR
q0Yp73YLWH0KnDp5XJsFWShGeVPl29xVSjnX1fgNQw3FxicqDNWB922u9nH8qzQ8
2g+Exd1323VS8gszvLzPhLo9lfGf/tzFGzY5xvygz3sPIGVA0W8OZ9bHjDE349Ju
kTNqWw+5FWPxkSYVKKaCsVdh8xvZ6yO98DmzbTiS34jdOH5PUvTg7D/3Da/kQ1oB
3P8cSPZ7ejWFhxnnVEyxrR2S37CXXLX9lTpVJLbsk4rP6IUlDIih9ZUvIyPjBfPs
wwSymQkrTR7Mc8NO7NYe9qn237bSEXMg91CAAIswxiC6jTsYXlBikcUU+fB5o/aE
8K1bonOUcm6x59nJdY6wEsN43fsu8MSwfQRcaNmm0sZ6KgW5koFmnIYq27AjJE3d
9tYW+Rvt+MsLnXZuw5cwaTE9s4bVhdOz70LkilHD14mc6UPyeObGQmGpXyuv9St1
jhSu31m5ErhUlRDpxa/HBR6sqFMp+gouy8GybyzUrAvL8H7dDGSiqgiG484isMBd
fdj2itlSrhD16V6yfCUPvgxla1RbfTWrob5jaEyg0bo2nKsjsauMeIaiz6hSTUwP
lYHDkl+Nmj32SwzSp3TGS6XTGZdNq/P9yWTB9LVW0Gydr4UcmzyveFmQ43rtkO5v
FQFbAEPwhq4W3MLV29T/glMMYbJF8wfMnQa3eM8NBHwLf0BsNoMsWLgK74XTLu8K
Kheb7hV9k81KNaTCINiFgecCuqmwIc6+FO13gphp4CjNOU4/U+QXTBuatE5BJtQd
k3LpLT/TZwSebeZ6ttY38Wv+EtbyzxYX5qWL4BoMOSucjCdAdD6ve24Fq6k/z+ud
JZSlWVFxTT5sSn8JPNK1Tv5cpaecvKVclKHbCe255/pK8JYnmkYvoBZxt+ICyNQN
YQgrsZJh3SlqiYlkMcP69el8nyIMe//7/HSn/QdorsfPo0cMO6TttrdiTT2th5xx
g0OOrDSFTZfM2VzVpR0Y+miCfePGqmW1WScUjF468IYW04p3WwYna10/9DYFKLck
Hh/BXuE5lPoGo4Hl7m1xcLwFxticC/ejFt3vYfeYmC+bRX9yCT87v777UzklhPun
eUdoFOftFUVvkB0xxy4BQc4fAyI8oH7v0dbIA+ZPLTybN3ltGffxI9owf1HhN1wa
/w+SpE8WzhPJCCrRpUFK/BLOO8FYCayV8+esK+OmRKuF85wU/ec2ZR8yoO9OYbO2
pt2Kz+cBNirEoZFNmKD071xW2gO+LauI033MwHMVkeCEaoqRRdKDrhdyEcfuPYNB
l6ecR3Za62Pul33A4OpbdDEpmCaJTTH9jwMKlcSn8axEjtND2dT0uTqVpQOAMRP+
RCBFfiSYyrqCiyP7JpwsRCIkQtQjhMRwZroDYcxKS7PaWZYl6HS1QsHuX/vSHXNy
cuJVHBs6ILke6NGdGHndUlvbjIZmk1K5v+kNCIzLA20VuTqRuu3g1pL+5L1yaIdg
cndz1tG66I1WtQjLqG+1K5xPUjx8ARCgR/D8ZK3iLbKuRl4q4xCgPmFhntlRP3ni
HljrRv2HDn/qovZkXHu2LWtMgX23v7SBDdL4FPF2SyS6N/8xxzRaQmEWbUQ0XjLi
LTe8K/huVzOD1MI1hztoy5QKDLJwFWbo2wxAPhA7Cd5eJw1Afh73ibLyIf4nzkr4
eHxlGI6p71g+mIbmmr6WsEufcfJyM5HWNHvKdrMuW7aLYsZAZp8ULaQlrHP/8jkH
xbCaP5sdgBSxoLU/zJU3Qdb8W2sUgPDWyivsBAyvdG/kz5f2whouwTzaiw2/3rzg
GnlXmRq+HqD9+Pz/+aTNbKw58rV98ADGd+/AsWOUt1VBoFZIbyoAngmmejpDg3F/
KX7NGwv8odtEG5a1kACp9pRjaXbsfjR8w6umTdujnLnsPVDQ7mrAd6xPFd5UcyUN
yBSf8WI9ykPdk+/bbUprjc110kMVWdbeM6OpArZoLDIALp/+KIUSOroFSNr6uj99
KtXm/R2c3BSnJ/uvv6a2qAEHgrkxU3zMcoNtf/+ECuPmMF7evIJRevpdG5te5X7e
za/igGQXcuK+eftVdkRMLRBHMo+lyCX4p1vmbEc8grxthL97nz/mpYnPnPnghQ6P
yXIGWG6uE1mE2m3fn09drTMjjteODlaVNwGfh9GeaLIAoijL74fzR0B4jQCbqVp/
lHoyzxwYO/fTYHcitS3FwaBbWho/ZSwaNEl5PnmTCepu/h4FX0yp499Ij6mm/pgp
cX6BM5B57FT+QULtzmnR/GZ+o6vUmGEOXJCDSV+Uh7tiwW5jGERpkSik+aO5LM8v
g//Rm1rRoIyMeOfBKCZC8+IMxOYviK6pcdHi9s4bnFzMjwbnPxIg4b3Lx+eUjkuo
8qc8jSRr/hKx3fudnxI5AiRjUtRgwe33HHbbpyol1kHSifdf3K/jVTumGf4Cqrag
5dZj2eVFrs0kgYPvK3nPwEVtEqdsJ0tmwkTM3JEb5HR1cSptb8NFBYiGPl/JkHEH
WG0zKIKd3InCVQaWYEC0QnortlHR0yGw/KKFX/YOMMsRo6D0fRQpltsgbRcseDAv
7PPWv4MYoBhvqHHz0UxLmkE/Xtk8LPr4jnX4QBI+ggkmMrlZoF+6y5wnG9JIqrI2
gQKwa/CbuorXZCE416PjYn8SQwnDq7Zjsla5z/Ewj3nRH0S/mUosAX8/dKI/JzWL
qSAP0pSxi1fFd/N+KtdVfNjtr7OMhaF8M6OYUYknuvwDEngvGy2vp5WtMdOgdIuT
jgRC29jmUTx1zxxtDDZgp6giAqrrbQ7STcx9R3+hA8ftkz48YoSm6kVH6XlwRgeF
un8BQHEYMtgcefvS9WKUB92cAV/HZ2+/FiSC70pWZ55EXF9hb1Hs4SrwtQutSneB
gkv6pfc7fE6ohBIp9jdsHY236nM6UZOztInBx4qAaBn0fdl4q7EHkiaCGEnzapx3
20F4xFnD42sOBnZT6m12Z5CJ5W334+9nubnRRpSR+aWF6jcSbn2QSds25VdDONux
fpkNddM51IABcC+kMY4cOBdy64lTXEu1+IgjL89OSn/DbH3N1kPOOXss9+Yc2aKM
D6323GEUVa3Dr1Q/P+3mGMAPljIX8hNwcPaUjFC7RG6Y6hB+MHP+1pLPwp7H2Uco
6k5W3NZ0GSAC4Ckm0MgaunhFYFSb9Jl684qZQLVHOwSgpZzrEhmiu3TwneeK62/Y
4pMViJ8c6ygeKfmGwq3zEuIods++ucO90OVgmpMIstUBBZImlO+OIaBbudG4w1Gc
FImTfI4fEbIXwlDIREvwxk5O2h7Gd6Cz51rnBzJVbyOaQxlr2OGpOmiQaiqlvn+B
GtcpthCthza46hp64sPBLTppInuVRwqPs/YmrEv6+1bac1guOyFfZQN/F4wPoFxi
Xq2m6u9Qr0iD4T4q0FYxfZO8pYLuedeGbjqbvMzZqBqZq4ikp4K0c7JXe5nE0taD
4D3JPFb2lzXuO6kgC9DQBJJpcm0QJ8TCZJG8bAgFevbxsP2kP5vUsIiKcw/woNZP
27P3r112PfKLJuLYYIfCCERvVuOI6t5Vv1a1BJcO/2q6AXTia5A33DFMZdeQkYhO
yUeV8Xt3myDIWtFV+1ZrUDYQdN/kk3xGTOeHluPb7YwuvJu0w48myyh9BGKAifOr
lkp/GUs+TnOJMQrn72wXDG0lP8/+oSIiVM/XoaE3JKg58JAGUhjWkYtR0EloSdsF
bnWb0y48RqTm8EjXM7tW8PmFNs4nl9mvqfmU3J0QDor4tLk5e4rnKJIdiuxhxG4w
iaa1NN17FMZ6xHtVRg4RkzPHCnN3qMQlJv1IQeM3AUndmMZNx7exYJM0C/N7U9bw
ZmdZi8symVAGPpwjPI0UK1aeQM6HbyVTW+DSUCpeIlQEWGe90vkyHnfvJWLcbKsL
aBs2sLvuzz7ozs18grfNJaQVgst3q6AuK8vlYKRHVzS7C4b4/HFSsEsaumQt4d0B
6Y7tTAd+aInE1bp41fELwSd/7aieYsKDEu+dsOd0/dZfZj0e45RToMuwj9fVa3cB
rIK+ah9fxUHp1xxx4otSRTNbz14MeKJGit9sbMv29u/lk+NMRmE/1hwGtgmJ4Qt9
LawnKMLd73Lr3tYftwVwSgTrth5Sd616jGJq4OEtdEHfpQ4V6xMlk4ng2JXKZbqM
4XDF7TM5Xttk63q/Z1hbpffSkorukSaoIGnNjSFy/nYIDUXa43CBukbJ9a8qC3TX
OD22aqIjqcuXeqLYVBDGBMkytr8rMgteQE66ZXI1AW/ChetIrYU41U/+HBx5mqKm
bRpZaBrkkqw2vaYGKrULscdZ/cw1JMHjlznKfzUiTffvM+YkH4SZ+MSVbiMPTdxq
YDTvUJ3N9ol3EQF0m4w+g8WCNwabhALv0u65eZ/ROnzOkh5U6jcSvD7JA/qJOs/t
TDUSybM77c7IOUGvKXyDmST5FWza4ovtVa0RRawcA1hrr2RYpWz8HnOFQ4fPz1ke
7BE2kYDdrODW0AF+azIM6UlNuAn3lq8OChVenkAI0aI89fAHjAtkB8qy5H8fpcmu
wVUvm+7WjX+nfsbxReB92ED4TGKHXshbSCOVdYzwQTfZ8aTS2VpsmqSDyKjc/v3W
TqcqSNTPAsLw89NgIunBm6xJwP78rk9n10Av0geMaXbRbbmRb/MypW5hEs0toaWu
WLtnLX/mDON6VyMA8V0nPck4o6vX+4QlYpmPNeKIfsYxW/IhYBwP82lDKm1XWXCZ
20MqdnpAyZoynLzdQtv5EDedRKZS8kA6KQG/9RowViuO4McLieEqXBOe3k5ADMFB
JBHgLK3a+ARcnVPZllI5h9c+PIj/J//rSe3BVF+3AnBPBZlm3++VaxhVoxOpW/12
K7/vPauusLrT2E7udGtiJWHEnsA0QFcxxuqDPy+oPwlk64b9yvpm+QXlYfLXfWsL
a7tC3tZz22vmxJRq8FohP7nPA3COaEo6qF24pd08POKOP0H4B1FwCRUneGkGDTti
j2Pv2W7IplR22Ad9F7DZ77rJyPaSx47Gp8xq7cyZGnsIBt1gAodOJkb3nJvulSYn
+qw874KsOQddYusycETcUGj035punsl057d+5D8mDTzf5ZxXFyLkJsXatpZo9gb6
p/D4upC6VvpNq5bQJnH5H2uDx0i82nZwcQCsR/AWfkwoWlWkEf9nL7tP9Ra+URM2
U3HiUoEjNqD7qoQDsWSc3ZZDoJbTHMiZcG5Nu4bGJPZK/I01xvxSKr4+qz/jJSy8
Qym6w9XrdU1G+bEvmFbcaLK2Wm6LxDaZ9c3pjXIyb132mpqYjyJqUYdF0A45Kmyu
ho/en3eqUNgfeuV40fVbLYzD5T5a0UYaU6PZfRnMTozSE+iwsoG+mlwN8k1uwRQn
FdopBpoWFuVafqD+BO60A6YULORI9LEOrz3kCaEpWc1ocXmAnxkShVmxjyjF8ScR
C40aX2+gLnZa+FhF6qtOjVFU6z3jTVO215PC9CXUUMEKAbkpTHeQZt/GMv+Z5c5d
eA6ZSLHsHhgP6pyMViDUF9+raUuXKJ61I2RwAhBZH3T+hDXFVOT0hJc/PhyNzH/s
bq22n1mFX6CF3rbj6P1jYEtvKs+10wuI6pygxNla/n1N9ilXWBtxtvG+UO3J0Mc6
dTUDBCb3onIVHiioYF2kj+6PnzhNqQSPR34TZWyXY+A968F+kMpkhfpLEUYm7DZh
2kVqbj1ZpJOyEFhvc3EEQ0lQrGYs3Yi4GDuYdR+OdeY3UwlPs6Iu+SgyfB9EKYOH
LVLSnQyonHVct//BlxXyWdxsvcI7FX7muf9mVyzBu2oRzOFkpmwh/0hRd6p6tYlW
HlX0GtWDJqYgWc7krkdr6qsPuGw8oQMdjZQLbObWwoPLa7DZPF1Oy3hcGJFr7f8/
lT+ek6ynpEPueUNvDWSj9eoLplg47kWRaobg19T70gdi73gf9/ajDasi6TF319CP
W4Z5C276i0jqKbCnmnlWVRZ/mZrnoMbFe4UnZ6SmYyz6u3KQeFc+puYf4bFuWpAA
dOaHG+r2ibQ51CuA8tlIRxwswGLSN43P9F23bvOStlhlEPTu+ggoiDPlAudcDV1h
1lElIszKX5oXygz8YRg/LeHPHdWgJEV7EjMMB7iOCUt9KM77xFvQzNmkg8c4pyuO
rWirKzozlDKj+RitmTTDCeg0Tch2IgqtipregOUEx6NrfQK2ckWG4frY80sC2Xzm
2l1DcWTXkcTSSBbO1vXERXKy4Hvr1iUPrUMKsoxRvTQGL8dQkRRp4XOxTzu+8msM
BQfSjtZHqoL7cF7+56OC6ywIE5EJG0klk58kujRGOT7Y3D1FGfRbqdifFH73V63B
bF+YAigS5jWmixfzoy1q8HUKww2gepICjPErgm7+9rM5eX/cP1g4OXuktL2NZ0xD
BFXtjZu1OKund0Kk0u5irU/JLL9jv/4JtKJBJGVSIvCkrxOzEX0gYdeSBtijoYX5
qIK4JY234kF/B/Jtdq7v3XpGjhQ7uiNUrFz0tU9ddLXqR4fXjC5yK7S+qTYkK28x
zhAjCtE9isGvZRlc4F/CglcrhkQGfjv0SS8eX7lAPsS61xGqDeqDQT2Wp6Ug3EUY
UDCPL2vw6QWt1ly9NrjbS+w4qV7LYK+erZ9588pCKIV3bARDqIkVpmpogtbRp+G4
u0HpYetnWpmrsQyhCygK0JKbUEXuGRgbFC8rMm8SCX4Xao5VodtGIdcxtdl7LA7m
XrpVF/1ZLS9iTjfgQrVDgX9g3RBXo/f43di66W9La0T5/hj/aevUG56a0oG8a9OA
fUntTlQnzwBuiX9oS9oGurBHpCgJbRq51tVwUibvY33K1v5S22oDSXzJJesuRbMq
WwPJLRRmzAcuc1DLvjZ71w5jvy7gE2gZ01ohBddw+BN50pksoAC5PjOZ4U9Jbmf7
lPQg3PKr9tdIweZdUcDpI7VbWykzHrRHFTsldQHmIhcxy/NMf6uw/e+AsMOgWt0X
ukjxggnGBI+lkGrwHbpVKW/6kXvMiZjeA0A9DTsnjHsOH+HF896AbIfvTDcrRwm7
5qKpee180jIDayhhiqGj8NikOb8qjzpwcd2TG6iEmqKZ7pAcXHM3yMC8D33xUCTH
7S146GFgDYpb/fIV0DyjboVIpAG+Q6DeqnmP1YtFT3iUj4/U2LbqijM11b3d4UU9
df3a0YMFHS09Vi3ymAZ5EmtQnQSJlfwpwq62GC63ZS3hX8c43Ni3MYzjwO5r8/u1
sDcN+uVKOp3XzvwL1lb9Uq3H+LlVW/lM5jgYDk+NNwvE+oJfXwHnomx2b3BYMnro
5lSSF0LRqIpFBsRIauM3vptopVHS9sPKisHIrw3JpJQD1P0Sm2NoRf/De10sTEhU
zCb80iIyGLMJw4gtmsOLyG7R+CYklG/OXTsFTOoLFgzn8zUZMMAfIl7iKCM0Tij5
gmcpEE3p8otJd4LEO+9+LStg9LFKkf0GwxkrRHMB3059YMONix5oWCZQbVTOoQQy
B3RxouLPGmfwunnZM1NSyWu/ZQ5HpcH2AJVIoiXsunl7ppLfX/+xm+Vw9uKDABrF
jRK5Dw9P4hC6LYNMVSRjrBUaySZwk6UlToPUUjCsMunKZOER/2vbjPtFiCzyhQln
AD0tBDOmh5C+xiWu/g7IRkZYNeIROcJSiwzVc+VnfbkgdFLEorEq0LDzFyKHSYPA
RHpYAKnqXfDyW9RhR57wwUSUvopUQt4QX9MmbX6Bt4FylJgohz6gcUy8fFixYMNO
1DNT/JA4bjI+VLl7tMWqefVdqZ8qB2wq8yu+2jWNbD2GR5n9WlrdTom+lzJdoX+A
66+b5UlXNHlGrj/1+Y9jrl9e6moN32reKt8bbD9zPlcsFglZLcQo/fseDqpD9boa
0amHH+YCaC7tl2z/vC+6WJS8DoX4/BLeO9CeBXF8yVM9VTvT3wswriobWjXTAYDP
Qq0OCQTfVn9yR+X94I1gSiJkI4gAICeX23SrzVvfuKLlwJxw2ZWjQ0wMuzeV/ayx
ErWsGUJD4lChE45/CoRU+A==
`protect END_PROTECTED
