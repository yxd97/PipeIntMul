`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gs7/2YsusUaCxvxOozYqkMt3uXFpIjohUpHTDghJOHeHmU9gH0dRZKZfA7qUdBjt
AcZaOwSQkhsWxxujXQTMJqTxRE12kAoqIS/0y9LPew1q7LA5gZkYGjcHHJLh7z3h
qarH0RbprS8B3Vhsdj31J4lV4M4UWdg+D1GQmWpQPCzxCo7UzLAQpYsZAoThBRLW
Yk1WjOkTeQJNSglITbjO2UG9K/UWnZwfpv3mEi8eMV/Bo0mxY5qplJgwkUs/9PiL
InkpEv2raeBk7db+ZVZ8ladBp6CKzIoGgr5ABGX2BmJ0DurWc35eEy+RcG4Q0gdQ
UYDyTX0BPEMiC1IZIuV9AUhUgDsqkWaLg1KKuS0WBwgKVN5a1LQyESiw+FB7Xj0D
+xGmsP8Hc0PCLMGzsLWfe0OT6qj425kUav1BmdEHi2VJF5ektRs4gAR5jw+0zH2g
m1zCiWhxNHhoy7n9DPd+RprD9fd5uuD0ruAI2/RoE+wpuAXvcq9HVcarZIqsel9T
uoftkpQ9aYo9S6R4agBuRlMAlwa8NqzQG+ckhcbfSOh4iR2WPPsRAWX2Nh+f80qq
huS3063ttwcnjNFgTJ76+A==
`protect END_PROTECTED
