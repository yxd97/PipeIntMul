`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KU7pedD1bLUJzYxrnrI0L6CbT/6iz/s8yy1jzg0adTbVNMpCkNR0DFS/yjnfxvfq
gBTmYWKClqjhng4++jtUXRWkw5bypziqh9nc1GYFTJ07b6KLHqr0NbVMC1Y+SNh0
jR7t3XNgwLU9EbIOjNFfl+DxOeY6EwIX9rZfP1tmEUNnLMLkwHvUBbOhhMRrnwEp
teM36j/omddvSYI1m7r0+LgdVLWAe1klLeFZCwijEhSwEUbP34Zyb0Gb7eCAxDD+
SW1Pye1vSnuWkdtTZfkiObOnjtT7DAlH3LHQdl63yjpXeI1JH9jwl+oYe4vFxMhU
p2GZecH5qWpy2DrXTT2608mWqalN1kjFKBrd5/xnZWmAtPdDlS9iz2HqmcPI4EWi
fYu+0I/zJ9Wcq7XyN+iqMZu19OqMD7UzKVzJmJsnFzsFDM+Kf8TpUcsZZJ0c7AXb
7MFOCBB8YidDJo1ho97E0qLqsT9TgkbiTDDZxHzS2RZnGYcN8vdwBw66QorsoINT
9HjdUi0dL2rss351TD0pofbkcX1dG9Sh1+K07+gQ6mKuyx5ZRgzYX3gyVvg82/ZN
NPSFFQeykodV8lfSlYwbKzL4XNpyDbbHqu2s+pfDHVxve9kttwno/zcTChxS5mK8
1cb9W8KwsdxnYysCCKYGfirGftPOy2kDbC+CduiktZr1Fm43rYVMrKNgIccKsDZ/
A4su4wEreIScF82oLyRQKIidbWZ5MlBH8MS993du37EHncm//rxg0RDl73pzkmoC
1kbphHuVmZZfWWzVUIFILfN3U5TaGMvogjlcW7Q7P7BDO6RsNKGrecsHvUJC2A0q
NGRnI3jlabrZjA/WbB6ycIXV8/lXaAeClAnfEtbcJXH0hu6fmVPs9R0XLX28/kcD
uclwpjdqZcJFY0zUXyrtFYupPjB+bwSsU2l+YN/5U3AVYOkqQv9pc2DPf06RjKjK
ZTxzArbr3tndDcpcHYULSPcpZZmLh4JPmd6ZCtgO+exX5fmf5lNDUkphVYuL5/d/
`protect END_PROTECTED
