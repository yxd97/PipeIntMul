`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eK5n8p4CuMMemU/Jt24z62074VGC16pGTnS0wM4TpqW6Ylqltm1j3EJC6X0432NC
2gu/teBVMoVqfUuAl+RfgNAZnnwRwA98ceVK5XkWnstpPph8pe71shj8JQt2bqiv
ZHfHdL73s+6C4tVjQKnkoeicYbvZM01l/EyAwzmOFXLr/FLK/CsIynNN+Ese5jty
XVj7Int/ifPpcdhMnhboa3Z6cyu/5KPoiuq8l4Bxp+YwcvPjtpnJ57IRm4wK4h59
D0FA6YOy/L5yUpUpi1VAZdw2hI8tVZN7+7CqyEcrpDwXgD8JYs9dDnqXTFswiG+O
RqL6ObmO+aAhxc/BtBHxmEp70dJJiQyQFcA6OtiV1fbRdlVFExw7fluwwOcTdJMa
bh/hGF+xUgWZZh2Lcuyr6AtLDzCJZLnGSXmcV5vYwOU0ZDPt+DD39qtAGuk0YN+n
g7Eo55R07TzRRe9NXShVdsf0x1OfiosMzuHwc2jwizOk6mdmH0IRMyk9ZtQGmFNH
pYfzqK04pIcipRJwiXx+KMlM7gcyt5J22QsR0QucgN1sI/qkAlZWKFEQmpVLdjlK
WOi5b5wBlRz5P28jclwLfn9zWBf2kKboA7socSs2LScSjVrrWfyc45er2anjk9Q2
LRYjFxeZVlZIpRjVQTdJVLaAocZesoCI/D+TiMnIOAE1JOdtHtW6RTc7OEzSRnpl
Ri/yNas4RTF8dSWexjJT7Ugi4NqQ+RvqEDCvGIk/2gpPPK10+GkXhnpxm2IAzbOq
vxbqvmSe/1rzrMgII7qFVQG9JzUgQHrxUwj0Qb/mAKtSrKc6sW3W2LzvyoGwtnAF
8Q/QWQfFqlEuWYln6H54Jw==
`protect END_PROTECTED
