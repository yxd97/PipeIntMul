`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PAn9Ami+D1vIkJMiGpS1HvUaIQ7oa5jUCIgrhvUQvi/eAhutXQiXg/Nnbjl2mDvw
69Qx6xmRIyqyfNtyVjYG254lBvUR4Ydd2a5CNegdGzx47fhAVwBXAGRFXUs1zNSv
ZKKAhxATN26Y9p6ARpEbMhGSJi0v7uDc1QcMNfVZGLFM4Yg6BvNWadbSZw71AwVp
x+tAxHaixRc6phplnlqdjVLoTtER4fD3wI4khJI2f2Qrskcwu7DSTBvponRW3nOK
PSDDLw2Qb1xMJf91S31rDFgWIoxAeuNPD+vLQM5nQ0kdX3bmI7/+bx7v2/239QF6
isgTdX76QT2I0R/8W+QX1A==
`protect END_PROTECTED
