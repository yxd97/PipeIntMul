`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qjudk/DhfiJ1+f5T15rTcV6gGmKSUOSz5780VDHHKGiIpeDxMfg2NxV/N0axM09u
SJJoS72s+lprGit++9pkxbq7vOQMYKrDIH4n5PaZR7C15etvcwQ/g8G6eKWcdI+7
QwjofH3OFHQlhY5srDc2MBPxQDpJPkaguvKADJ9WMZlWIKa/kulrej+KUO0ka6Aa
dz26305GsRgfekdqqy/jpHY4WA3S229G+NaO3ta+Ub6J3DAZWrSbK4iJE7nQL0Xb
GCBBS1ZQ8s6UjfuyeMLOxkNjyvQatrmlxKPCeYdsQVBtDjjEuXl7M6sG6co/IgMN
uNgL/IK/B8++bii/jOPSErqRaKbicaiVvrMBYlN8P+/feVX659m5eq93IjoBEdS5
iYGrtNYfBPuU5dAvqNfTKWXMSR6sR4Ldfnn1gXUAPQ1trYNMsXlV01Xsuz29ZAKt
pl9USUnMmHA5+laf+Vb7gy7GUae//swgZW9IhnAnuxwJ3qZ0qVQt87PcZguPa+JP
p0Zz0MR1WUUKXwlLvglE3f2N+FGT0PHQ7Z3DKI7q2HjXb0l0bW+BMAp8jgzoXv7A
`protect END_PROTECTED
