`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLjFwMMGO3ZAaR6TUKUtiVnYFQCVrwnesCsnAbnkieAazaabaRx8VgeHdKc+9op5
PQn1sQv8eRJEW2zN62SC2FcgUUfOATHtAyOHDJ/LyUBEtf5Aj+IDSWiVHP26ReB+
G/i/IlzZ4POd9f8hkq1XDKtSDlT3FOKY69HNt97rdEGBB08s/XebkWYaHEgUzRLo
erVpFB6UgHEs1ROukRXz1VhHZSNh37oa81vfbpIjyRdGDOBtmrSMA0gTNs/WP9Ik
N3v/41ERL2yWzhN4dbBqk3/PNy1/BwnodHXEjaE8achd9YDYceBS1Yf54sHlkqKL
Ls2bAy4BOmRjNmIJ0+rzMusxTOamYEGVPmkHDHx+yep5FWiBwGTKlc2q4zF/g4cZ
/p3RQ/78Q4HAPA0ZYAJCW0DIKEOk7u1WvWXUhKcLfb8la3zwkoEa85tzbTsxo9OI
AdpnIUeOrrx4KtY4ig5g20dg2bgNhYBZo8Gw1beK5u8=
`protect END_PROTECTED
