`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7rJlJ1rScUasrjtH12KEMtjA0S+KbUA8RSyk4LnFJ0JUIpcnr5y7JxDkwIqNe8wS
rPABlFKYCs3lGwjRKhr5namUfn6Zx78lx6qGoKea3tyjh6mxgKnvU5XjjDfLVkpO
PWYCnWXhlx5CQierG+AvzTJishhrP0Q8EvLuddBYe0iImQ36DAngziJlSXq507qW
gYwAocFaE4Vaqr7PdFtrr+vFEVqTZHYR8bxGT74qVz9YUckL633t/tAG9aCft8yg
NtiNbZhrTGBh8tWYt6++ogtxHtagdyurXiP5sx2afBXuMn+ReMzTK3TP1ceTToad
DprMeqXo9zzHV+I3A1NVevfpV7c+I0HcaRxX3IF/U3WkDmY0DQFONflCkceMnnY+
nSlzvKFk0e7HcRa3ww29kxgSoD9HnlFrXCeAlprmBxSjSZN82LkKgMoqlht+BP9m
hzm5ITGPDz7SKacLMfVxFPUwmTTou1wJJMCEs79uvqVEcs53f4r9pfIbgLFBH/IR
4qnowrt/pJY6kZgRehBE1NpSOXd0W6tfJ8YhJUiUsZDFK+jtr6/ZuxxjrNtKxjZ8
EYcoi4dinOuKYvjDs8uI6wHys38Jwe3C2iLbAIrm2nE=
`protect END_PROTECTED
