`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3iuRhFOscwf32wgvfaWgE4hGHN0dRnVU5VYDNKh4ANtTMPyCDCn6BfQbNipTuQ/
6l5Zg0xk5ExWoZ87d0S57a/J/NRPVSqg4Yh8F0zyxhNuvaBlyz9tVDPPpVcIjtSm
RcfDkevz9AqfLXc/5sbD9jhHXEnk3522N+oTFClka7pUDEO8FoGLWuotoWiIz2F3
qyIB7Jx67Eu9RT46nkrj2upJHUTYUlMsFYB1fBdvchw5Rw+XH9YQ0NLmvLZ5Bqyg
SFKTeb5am1VK/pGxqh5bTWfD+IJ+mzjsRK+ywU+DqhGSH/9mwk1ihaURPl/pJHjp
Z/lxfjt5qOQjSBiYyba9228nSUchHUiQmt61QhnRNpLOte6qL8gqiEdNUb05guN4
TYCl0taeRMeNjQurbfnhbw==
`protect END_PROTECTED
