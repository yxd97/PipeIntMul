`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JtEkQAKFJOh/R9nm13JXjVxc/jvDe2vC/afz/H5w7CfTrUPldkN488uwSu//dZED
O+5tpeyg9n0VbsAgECtmzl/tQh2tE5wpAFisXzvqYHybBfTuRvBmn5PpxNaYg9Dv
aMiMMBh72vd4u70mfUXyqRqyOO3rD0ILpXa0yLStOlK5ac9eD0sLRF1ANuoXBeKS
mvEEQKFXkGNYy9YPk86i8Jcc2cLucJ61ZN8blbYfILiVhmb2fehVTK+yUVJtnHTR
b8EH7y35f2CboK6d1B+g1xuX+61cqKGK/oQNhI7JRXMKrz/wW6wQ2AFYfte6UsTG
fV4XFmUI+v/YIKY9mqfuJouzYzN6lPThRBd0nE1QubSYrL+a/yNyh4TmZoJoS4A3
5MfS3QbrHh+Gw/I/VeuAr/Gx4jHCvX9HIlYAH0UZhi9h5PJIhoyBwojWodv/cm4B
QnPXqgGWs5lG1gGbvstGsj9wMGpFHgRuL9Dzs+/dvUk=
`protect END_PROTECTED
