`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2YYSA/am6+9DoNm+QJHx0T5FJx/KZMhHqbe6f2btb5uF/BFpjPYOfd2+PDGw/t5
gNlsG6W3v0cvyjGwkKB/Rn6x5s073julQFMJnCiSMZovHn2QC6iq+w/fenvrXkpw
ZRof+w5DbhZK76tU4eeDxNIdLRjN5rvnYgjXRnD497BTGTh8qIUYxHBmxwl4wlot
8htiAR71NoXt31OmD9N4ZY8/Aq6J6v6AJfhQrYqjBzCjNoSnoUPoULVYePPwkNTg
5KEXIvIgL9gaDeGv/XAzhjUbEu9KaegE8085U7iiZ8cKPwY/NOh4oOewagjmKfVj
rVKPFRq/kqvVHg1cvdJD9C3khZ3CVvLjrSRQofeKOgMclcBsGRMXNcGTU7kah+CT
d9cWLH4/wOxeK6YUFHG/avw+u6HY4z6BA2VH3ASQLmI=
`protect END_PROTECTED
