`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+WIPKYJPeHO4USKaxEKAu3yt7Qd4+ZIQEEwmRHnNasFVbGz8fsdn1jS3RRRYbC7
JQQd0U7Ip9biD9LhnLaKx2vV++EtT3x0J+9njIhACNrk7QcL+Kr3If8rW3LNpSti
VPwJnTqwfN/Q0Zsc6HnAQ8Sr7RfPZxyMnUpwrYmBhaaTe9f7xtPt2/zuUtoNdH5U
WwB/tldUPz1HZ2DPKHjD6MQntt8zBNoNEvw1QSF166ODrPeMtHE7v65U4DL1tK9p
xE28s+Ke3WbLg/R4GGpRsp555zisap5u/96t0gYh00APvpUpxWvFAexjDQFnyYdD
JXq12inEw0C9aVB6pMvKE0BnXMhDlfEWkSA+32qJaMJQNNtDVkZXKzElg9QBRxoI
eM6Bw8UPXpGPKYof4AAhLAar4ZQX7m3ypD74DzBzoqnwhHGYLKNKVdXhJCRmg2UW
FjtRnm0cwRtWkYrwhUBMWIJ3JLeZ0vtJ4LWhah9WYmmEV98YB2Jsc6L26GePf97O
+HNGaSYuoEGnRXqfdsSzc3Vk0FreFkty+R3EndW/FZKWrFVdhEI+IGOoWGlb7yz0
Ets5L1qVwxtci51I3ATO2CvAfo2LwGGwoaD2RTSOms8=
`protect END_PROTECTED
