`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AtDmuNLVYz8bUiz4OUZm0D4Pd8w/lo8Hvqom2T4Llhu1YsbxaVpHQCwRYsFENnmp
eMcwc8/rfbFOzEQj/dMNgFrbQ76fFezhlAX/vmJM0SpO10LKZd3FfvEKPbn8qE6n
0O9B6Xx/TEnn97SSYfMhIfyYszhXTqmseopaGusE4VNZMeRiWquRIu7B70bRntc+
AIQtmoMdtd9bbMIRLmZTS3h0uCAmfRu7N97laMDvg0mygZC1Ng/nV3Xi5HbymC2W
PNpGUeW1Phb0CG8yBlvImo3p1NgfyzifBhVkjAlxJRs8bZTtGuSaQUF9oyjyM+N7
z0D3hjXZj7mb9iA2bKGj0g==
`protect END_PROTECTED
