`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCT6END5BkNnzkUe2eS0eJZSvlwyld3qbNT8UX1u/+5nOo/v/5QSg8p1YEecZktO
Q2rwmV2D6RxdSgir1CgnIQSXtcfMGc8ajxaJW446WqVugV0CbzTKL+OtEKrMpErR
P2DrrDGO/z0UsOO0EWrf2bkp+TWdqvMc+Y43JT5KCjpNppnnaugzHULx5xF8PmcK
lr7kLV1XRBuQ/eTITPFEIEtXt8czGocEGctr9utbxgiQRdEYlTg/GtIbbOeHh9Vz
osxgD/eT97avuutp8TU0UwYCUAvpA6IDllRzYoQHXTZGQSju/jcsLOPEpPzqPqS1
u/DKjicyzsh9O8mJxkaRIs+7scFS3G0WXPwcUTdarTfMll9XC4Y4mI94VKZnRSc1
W4DOqZPHVNKTWHCTszGSXk6J+WWaEPMmMOloL4Oa3zSr8sdkYHNPt9UqIgidQ3TU
BoXRf7UisF+lIwSTGVjxFGVj6cU2VFbqd/O4twV+gbk=
`protect END_PROTECTED
