`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68hcz/S109kfgaULev4kXGtRyy4yuqfrhP9VLiegZapdV7vsCO7UOT7azajml1a+
nGrO8LFRxiDf7otz4fYYRAsntyS24NJIbYrQt8u+hmBmdm1IcryARhPGDKYJyDRa
civ1ma9urZvQjJFvHV+5FTbhjvTX/4xVnI3Qswq+Pgai/vCHEqoFw8YEP86vGWAO
jFwjeuv5UTKuJhsI7+QM/+l0VhKRsAEjDr1bArs+IoK5+Ypbxt07Mg99L7vNrCer
l7SUWlERuNKQje9KyfZAonuEYC+5kNcb8H2ZJGmtMAB/nmWaVT1cGSIpH6/ttBh2
PCNChRR9/OY8kthqxdfBDx2YiHd1+aFKq7GHY+vnvcNTdqdiAi3zmyl0ZlfbZQMI
zkK18xF2y1z8Or+0vnvlJQ==
`protect END_PROTECTED
