`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9TnTvrNw+Mhao0MsP/gb9TUswKSArHqUHCzW+V7SwuYEaUz3uLnHufrwe9O7DKkw
Hv/IRtSvg+b7cCT6bCbPzAuui6pvC8OJryJr8MIjOzLSHy744vgKpX6LkgnjTJhp
vKor3t6zUKYq9/19ZlIhRi+lgtwRvrbiwm8FYDVcB5jhbkpYALHj4MP30B3i3bTw
4FDU3QC+N5oACxoMVXdlk4KeJBy87qYIRc9toDa/CGeuzkz1kNZpPTEBx21FqgII
RVOBjdKsNKP5T9qCVTGH0paHmMFBMPZov62XOL9puCnY17VjerohVyM+UlAaOpnc
7WSQvcIMqNvTvQaqu6OsTg==
`protect END_PROTECTED
