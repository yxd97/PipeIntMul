`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6pLqQk8pDaRnYNMCS4lx1Q3qokUhxez+1Ge2a2x46tjf+sdZMzGhe0kHLHS3se1
XYhlXRXnKjbemnUTdPLHklAAarPtjHAFXQKSb0gtEMC/59pd/qxsvxy8k13Wjq/5
/c4H7ADV0BEj767475e4fcxDjjmV92zxcM/+nDsRdCITyvCiH4ZBhgyFrs+ekyXC
JtVUlaMkoFgYb472AzACBnqS6c85MpLRK4KYX6RzUao4FhcumrmA2Es0IaTU8SP4
w9JZBA0Sm0Zr3FgEIteGyXdAzqzymehlI0ukjgGECs31tqzlt90TX9fWd3MGuIIE
56CyytEznkFpU+AqE9XUn5FeVUE7iYZQ5EaDG0ibsDQU5pBZqfN727pfQMpQ5KHX
6rCHLpaGbVBC6Q4XhADwOKuUjuFxzbEnqGlzbh0/cJKcOcxrLd9hwCtqK0IBtrrA
pPdjF+LSsjJvl8viKlHk3HmL4mrRDxjsuE7gYSoNmFpAMuIjB/VqfWGtKzQipLoe
GvzlCEOJhU0TmcCeIsYn9Do3O6Yj+UQ3fv+UwpXW6Y/CMNg4gumW7ArPzgGKB8sl
NvDHj0I4NgnEbYoiJBbPKGBh/a64wK6VTsH8KbxlPVMTB3UFKrtecsLWdn7rWvgX
p7EVfmHHh5nPoOMAGqiGuoDOuItObj/B7xNODq4iNPDBLsdF7Io+xUnb6slU3Jn2
xIirkSpSp9Flb1EbtraTtNghW/Wl3Tk4vWpFvsjwp5fwGsUyWGYpX4aiSQ8v7LYu
bOK4sLcihztWry7/GzkjFzd00Eg1FFb32s/81r6CKwCtjagPk6BcrCVrxHlR3aKx
AwkN5Zg0Ztg5Jqcwxg1Wtk1RssRCn16oiG/7x23PN5mTxqgfQoXQLrVku6vvWLGs
E3YtHUcrnXDVaeZ/eHpo9soKp+r67g1j39bTUDYozJF9SWQAX3pTDdz7FvpsJi5d
wcWX8ucTq5c+ocFcfmOxKQon/o9YVUkxD1RZMa/lhwaY/bx+mndKxbGKpKJ32ba2
723R+rI7zTJ2bcV/B0aNAHfAc+7LHd5DnBBWniNKmnvKra6qnQROtALhK5jrjsds
jbMeqg7QUrbf/AKi6rmrB2jMlpBVJfjLjeT0dK2RoXY5/u3NcFXOvonWqmZKwJN5
Fa8Q9iNpuF0h+hXSTvUmrzREYb2RkuP1AZpWLkvC6T1+htHzEFDAArw731J0gjSq
3DZLgEFICi4/VLg9Hk9Ri+6KEqE9E4nyfmcgaeQQzvu+kt/3V8hqV5a6bKjBV1OC
objKPamj7t3eUeVbWq653RaFK/MMOH/c/1GEWHUHvbj+atk9lVeqphmwUmbUEjHi
R4STnSA3PYBJS1fBSTGABWYTsaMkXtsrYW5poTIleJJlEVlzCP/tkjT7bLrtZNFr
3S2QehOs01xlT1xiIrTqI/+m/yJDY2XiKbpTg3dFJd8EXdKYQ2BhyCcJ/svlOxcY
cuinYJxIZHBeNmcCkdoIo6xJ2R/9Tb38QgaIZoHELaR5hReajXJPvoXt3CAB8btb
rPlhSdS4o2mFxwALWWNQjyZokKYDZK7QuJUgmgI0rZd6ThIUyG1xiraKR3eeuyWD
mL9L+WWCBykUWPbN1ag5NDce+q2MkQOHhwVWQ6fgcxD2ma0CwXy4yUhwllgdFzi+
NEcwwKjEJ+vbCgZ56c+BtfWC6ZhxfSiWwoMDvi3h8VXFB7E46+6nYU2kIu6qTZ7c
H/AKhhdxpEgboLRRHRtCuw4TUP21+nFZu0+U1hPtR6zk/PLsNxoqWri0bl7/UbG+
vC/GYSUx/R6zr8JKE+JEyWgzJwaoPfzV14KuUObPBB+c4RGWTH9kROoSlLcUhjq4
9Qd0giNZY2IciAEz/pxT+xvgWjMGwvMgT2dT4b/FyqsEv6a3yeT4E9ZSuwlkr7Aj
DjngFwpcRLi39K1S93ra5wsh1v4VRpyUEEINP3evJ8ujkBDBMdiY9dStm8330be2
AEGiB34arw05AckFOByTlq0wethtnMij+38MH5my0MzdYtRMXbY/pzQkSIP4B80J
aiePtPHBWqSj2mIcDV70ZeMNIwE84kSlnNF23MeGnguADzWMOjNCZOEUPUi5pV3w
ecMYRuq04/vTeD+tQTOHPKXG9lwNfuDMf0LcQvvBZWZn9sbGjVEEPtDVKY5idFbt
nn2fi6BMUcLpaHmx8JVE1c+Udg1Diw9qLPRGFLFA91WFGBzAeHSilAiG6mqqt9wy
aqCAKLAbRMjrpdvMbiSnUSEfSpairklLgb/slyROpQ0Z73MWwBf1JvX2UQ+eJgMg
EpWG9IY3j0dXuR4baOykL6aAlQOnMd+u0/84t9TV3QicywWWrgYIUQF6nY7MXKyT
sK/H+cAKCfiL1JLzJOCa7dOLrIY2uwS3gn6zK/eogOz2FwVKk9hIpUnypaXbRtvR
/Sk1AB6z8f23KKbcr+wuOj9S0zUwfyqipuiHJRVjcQ1Uc4w6mGOdt5b+ECIrkVg/
Q+bCiSTmQTv05NNMedQYrRvsAf1tHOp5fA/RGARTRg/gC1XyFlq7mCEJxpuUv/ns
LlYe/KTnuxuqUxWu/HJdi+ip5AA5IHolPz62HhB2yqtSgkyt4KiD/cqMmbfKwcgP
KtmZom5V86FKmK577raS3H9c59vSEO9h2iN2oSb3kfJoOzVzZ8ZUGp41abq1YHdI
v8jkj4GtU71Nc+1VmupQkxfsY44ClWE0O17E00z/tfRMbgIb8o0RrE4GmwnAeyVC
RJXoRYI/ghiYCYclcX9OKmMSKPOY9YBI9gZaTBFVcAK6rQ9OH7F16zCBkluORQMg
pNn2aHGF2S/BiPn3sFg2+5NcPNT2K68Sqltjk3pXMpqTMks8P52ySc4r8NlAh3X5
3qsGJetfKcrowhA4Ify+NByHLRYyMThSVD1Azenep0hgaP5FpWhxbVmUW8FaBT1C
hMApAQzsEDmfwaPK009CQHsiXvP6O+2XRc099PxspL1VsOf++yVa3M5gh2C3cdOQ
QLEeY2mN7256pRAFQnfQNJOQHkhVpe+OWlFRyR8FooPtuXugBfXfr4klOwYI4tZV
qYvAbctXP0RLEpsX0OLwSm8bZ4b1OJi+kYIJMVYekpWkz8V4aMZRjzimD9mBxsju
KGMvkhiiTBEp8Rpmsn6ehGnI1YiO+NKhS8kUvfXiW5G6OeZdjulxJ1wvklYP4bHg
ImZ9ruzu311eC4IpvDC9wPSw4AopS1xAGwZZH9uC0stwhcTILt614El4tCXVU1ah
ukJDIBGbMvAYiBfQNF39ZxBLQRIiWVsYtyXot/DxoUk=
`protect END_PROTECTED
