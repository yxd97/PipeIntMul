`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LYbspDCsIWwra2Q6lVoGf8o/4ee33oI7br6zrcUKWeLHWdvr7HFBMMthCP78QryN
/BeKbi8wzdmxCPgFElo2vDZZnGGwumro+HkUrP6HZLrLUTjzEd2YG/fo2ttKx92j
hEuZocd28a4JxCvI+6aSJAMMXtZzVw3bXrATRcR+Pf8GxhHjXIFG7MUTckhcqQPe
mg+qsH5IiMHtLgXVu1ozMd22C4aLZ0smT9mVXG3CzEslok/IDdAs49LdOKH/2nA/
lS88dphZGrcx6kEOYVpwOSnX5lMGqJaKle92/R+DX2FDQHszVqo686wYthIzkMOH
IefFikhUp0iOBHfyzokeZEGDucZfHo/G9dggJn+ck4yaToF94ebactP5UNrV36Cs
PTpvtrIrwaXxSyNBQKu9oUebQGy0HMVI+L8mKoapw3hwhCVlQto/OyaM+ULRrNuB
LDDikkb4fQcWxQqFzMPQh1zaXwyxJQrByGq0Fg5W14W39SOtoE9ngQsb8hvZmX2u
NhHigpIPtX5Ge2l5aqRwqM9iQxMUx260wr3U5a7Ro7NoEYQ5DJ+5SxgaNx6zvY5O
mJttz00U4dQA1b6X87MX5Bm1x3Ozxb8DgMkNDfl7hrafhCC4wdVO/FUyR/vucAWZ
yCR/5FchpEUfu81VXFRbNys9IwIHt/05IBgDuU0Uf6AOA7UyDVRhJ2C6VhZEnwD8
L9JGQJnvet4YsWvFnvACM7kUpFm0LfIQPs1uK8eFx9Mn3WVMv0vXFAw0FN3Zpxnr
cBD8H7xyyoZdngB/FPxy9fPakmbjwyio8CYbSc+w1rooavOVpwW0W3Ganyf8qQ0P
f5zlJq1Lk5naTfWmezrzp6ZmpmFQSVHC4xYG+edGZEmXVxnsOr7gW0uK1AyPy5VI
CEcsOnu9cUHh7DXXILrlBO9GvVANwSx3Bd2+O242GIJ69WdUtK1g5uH/z1AWJB4b
fUCwq1hjzqOvfN8jJUKapY9WgQVjp9nIgQ/42w8neSneOt1kHMjDEXMCcZIKmlWK
g1btKAXWdQdMZMINDM1UYnEZ0RJUM3shnzoTZ003xrsy7VhC5Iga9wLgfZsvChxL
pZYx8c1Zaw6wcymUoRUZis8tkL06JGIkiIyD6Sr90Yy3ne5Y7fJVxx26tP+FQf3q
oe59/zO6nTLSLNr+2+hgQzoMECha/ClqySp8+S2hDnBKo/bGFz0Obfo2Dqp/PCSJ
nXrXGAEm4yeKozVV2q81gBr3k46yNr8cELtR2e+y+2dOwtnTe2BXlk6BfsffOADl
t6PIDUtACnjPt9btUUH2XQ==
`protect END_PROTECTED
