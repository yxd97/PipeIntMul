`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZc1nJ0UaEkdV/HeuZDgkCMRWz1XLrBwsXOBXLg5nXndr+aqeZry1LUvfaqk1JAg
F7Xad9uhVOJUA8P+d3+1HMGSzxogX4AMknL9c7ZhqMGyBQCXOL55DIoMacByqobb
qXsLsxgMV/HXrvhl8AAvcR7xHKved93QjENwjL6vftSRJHQqz4hoZGP3hyQnPU2j
GrfmZljmE8OZH/GaDMnSRhjr4fYSiO+RmjINj64KnpFGG13kcTvqgnb2XRCPsSX5
IhH++T/1jCccvEPhw8zhHJXE6DKfIXgjdADjAGa2uZWqSI+luoFBztZO3nBVltxm
mWad87EcGx6Zce6IFoFv4QJwL48wtRDoG9z22khLLsBMDwuZ2Rfnx5WOPaOEDywL
k+OAPudezoP9rSnP6n0rWaDAcxNLZKxTC6XWs7rKa+iOcoS5aKxNazKcTe+0gA7/
/PEjYw6Aa2/hMHU0eMwHgGcNegu3qYda3hV46P2kYU5u/DkG0VQrZEoQ8LT+MUvO
RQnCPuatvPu55DPKTSFYbjV/8P1gdmqC1wlH/xctYE0vdmmAkEYu3YpPidFSi5U1
UH/2MDlv+9D0+sEJZU8oScRg0H6UpGHvZy71ZUqx0rY/Y7s1NYEBsTpQ8DalUXDa
LaUjZO9Ilvvon5VTSc/bBxxawaCblt1L/eSBn4XH53KMUhZVHuUsjWAuv01ba2+z
sU2XDL3gtd0NdVlx925AEvDnMHWRZK82C/xnFOqmXSEXy4awfLhE6M1kOmnHhtFi
6Vnfcig0igKn/QITEYaTQpYDQ30lxUAxqONJs0huALkWm8zBv65AOcfT5+pLqhOz
XxdhlsCP8B6VMnLCt6M9RW6pUXqJFLVMwpaw9vcnzm6z60xDzx5dansKFHInpRDl
Zh/vG2QD4DNThXxhuNEoaSHIg7mFA1YobPWMdh9OKKPSP0hvUObxscPb8Igx4HfM
uv3KjurMx1B/qM/a18nJ7mch5NI4B8KooNOb9lOEf2Xx8eg8HuDJUSFrtP1JrQas
Cd9Tm1BLgodR4zOv0Y1p5ffqISNqkN5giwYXoJhu0Rum6GebxDieLeueKpe82x0l
ZHVw3RJdbJ8rYfxvOJFVYn+MYPgHOT7DZShYTibb1MkIHvvknbZzaQjMXMKKQv2o
xj865ryyIw3Fs6P553KHsqlQ1AgP+wRfhdvQnw8TlZCYisrToXYl/itfp8PCHwI1
p4UOQ1jPpCuodo4mM5Rvb2vfAVRvt5Qs3UbgglyhokkmokBEtbZpAZBDxZcBDvU2
CLxAENRgsQo9HHeuAAlzw6TuGeK/5xSPOXUchhI9b1bltxb2Hu3/LeZt3d7SzaGD
wwbKe1xZ4Y9pCSr2RAcWBu5MzHxh2XQHn6h+A21wxadr3SlqiQHJ/whLTWlmyUNG
C+nsVCRKmfqdavEO/3XIb2dB8dJpgXDWA25P/VBQ6pZ0jgn5Z6k0P4EVeFhugd6+
SBeM4H9uI+yK4YLaRoFUFPC7PDbxVoZNPEmuXLRSVe7CfUNHwlVMDjc6iESkIWuY
XtirzvYVRZGb04gm+s/4fodWQiVw+QhgW9FfYbqCI2nJr/irnS9WjgXqFIapg/1T
MfgwXAo+kKvbWUYKAtuYJVVjIYsMBuOkCkWoS3j3mevnIhrPdhrxIuoteuSbG83i
AJOpiShOmti3BeIUVrOT2XcDoootXDK8KD4Q13ohI1UaG2pb5nIzK+AnCeWhpP8D
hi2sKVzcbuilN24c7LpyzU0onQYsKrfoqjWWYid/oa3WO33cOzq7HLFHFblOHjsy
e4WLGr6uwukA5ju4Dc2soTOisbDrgujPDHrkb3C2DazMwVtHkx9cHaf/da76MgrB
rkvlQ6U2aiNzJein5apzXm5xmvdKqDZBU8qjTAObmt967hnQGjduLvfT4fPaYwYw
9Ta9tkypw5AgZt0DVaC/X9PYgFWC0Ql5V/sw1/EeXdTvUcISX2kZEy1iUKDqqSmR
+W6RX7r+HiVjDGf1RRoo1VKUbcBdA7g6tQjQQu+zWTe0KDnfYaOsPW/8UhyY9Yvk
/UdlIvWRfEPQrcKeYi43a+ng+GKuz3GL5o1cRGtHwX7Oe1UGuvut3x8qJEm4utzz
Bro6Zvyc+PYnuUXLNtmTMw5poH9cdgc7LjlksaQYYnfZQSvRXQdgwpSQ530NlenJ
GTCLIdew5MhJxFNkIZCPHQD9Ve9136G0kO1oum/bpbWH8QsT586NclUZHek9nljr
FmkgSUlvlIzO70HHAQK1C/cIrntL8IO/JfNViCQnzdCoPFkIM1iBq0xdR3cHVMnE
+m189bDYWTZ3DV7b/5v6Hx4BZQTxVwymPp+nc7ZFiV5HnFn3PRDqgW+1fjQ43Zhw
ZhAgASBv/OKo4qzpc0ANoUHMjpCbh2xi9QIjzcZnBlpSysHFg5FV8BWxdcgyv4ZO
F3oTE5YwidpaMVoXSRJbHFfl2+S0iKRfijlWB8L9Va4jLOLXA32HppucuCUuUwFm
`protect END_PROTECTED
