`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JMRTZIDrsUbh6zedUF3eV58KDMCin19zeJ+Pg3m8fYC5D/31mhuH/D7krRFQdRF
ihvesLSTU/64McUhuhblsQcCn5rY7e4GyX1nN98B8QbdOXB53mFjFOa4vmOCZ+Io
A1yK0lbGqEGnHfqJz/IFuK4hWRuk+/XOYW5KLCVoGeT5At3gtDGW58IdJaLCq0+R
o/9lQo61KRJljoxjWfNy8lKcSyKHL7l8unM6mM9FwCYFZUtnijXXfBp2DOFr3jNc
RA7L2dionGeLKxs3xPXZ9ikoJCHup4h9tfiEeG/Q4p18AYR66UqZbU41BB8hrvVP
IHJM3wEULyriUadCFLiJBDzbsZyoIFUqg81unNYwtnS+7sXzjLmXtdNJAbJix62c
ocuFSmuwk7N9eI8bQud/6Q==
`protect END_PROTECTED
