library verilog;
use verilog.vl_types.all;
entity BLK_MEM_GEN_V2_6 is
    generic(
        C_ADDRA_WIDTH   : integer := 5;
        C_ADDRB_WIDTH   : integer := 5;
        C_ALGORITHM     : integer := 2;
        C_BYTE_SIZE     : integer := 8;
        C_COMMON_CLK    : integer := 1;
        C_CORENAME      : string  := "blk_mem_gen_v2_6";
        C_DEFAULT_DATA  : string  := "0";
        C_DISABLE_WARN_BHV_COLL: integer := 0;
        C_DISABLE_WARN_BHV_RANGE: integer := 0;
        C_FAMILY        : string  := "virtex4";
        C_HAS_ENA       : integer := 1;
        C_HAS_ENB       : integer := 1;
        C_HAS_MEM_OUTPUT_REGS_A: integer := 0;
        C_HAS_MEM_OUTPUT_REGS_B: integer := 0;
        C_HAS_MUX_OUTPUT_REGS_A: integer := 0;
        C_HAS_MUX_OUTPUT_REGS_B: integer := 0;
        C_MUX_PIPELINE_STAGES: integer := 0;
        C_HAS_REGCEA    : integer := 0;
        C_HAS_REGCEB    : integer := 0;
        C_HAS_SSRA      : integer := 0;
        C_HAS_SSRB      : integer := 0;
        C_INIT_FILE_NAME: string  := "";
        C_LOAD_INIT_FILE: integer := 0;
        C_MEM_TYPE      : integer := 2;
        C_PRIM_TYPE     : integer := 3;
        C_READ_DEPTH_A  : integer := 64;
        C_READ_DEPTH_B  : integer := 64;
        C_READ_WIDTH_A  : integer := 32;
        C_READ_WIDTH_B  : integer := 32;
        C_SIM_COLLISION_CHECK: string  := "NONE";
        C_SINITA_VAL    : string  := "0";
        C_SINITB_VAL    : string  := "0";
        C_USE_BYTE_WEA  : integer := 0;
        C_USE_BYTE_WEB  : integer := 0;
        C_USE_DEFAULT_DATA: integer := 0;
        C_USE_ECC       : integer := 0;
        C_USE_RAMB16BWER_RST_BHV: integer := 0;
        C_WEA_WIDTH     : integer := 1;
        C_WEB_WIDTH     : integer := 1;
        C_WRITE_DEPTH_A : integer := 64;
        C_WRITE_DEPTH_B : integer := 64;
        C_WRITE_MODE_A  : string  := "WRITE_FIRST";
        C_WRITE_MODE_B  : string  := "WRITE_FIRST";
        C_WRITE_WIDTH_A : integer := 32;
        C_WRITE_WIDTH_B : integer := 32;
        C_XDEVICEFAMILY : string  := "virtex4"
    );
    port(
        CLKA            : in     vl_logic;
        DINA            : in     vl_logic_vector;
        ADDRA           : in     vl_logic_vector;
        ENA             : in     vl_logic;
        REGCEA          : in     vl_logic;
        WEA             : in     vl_logic_vector;
        SSRA            : in     vl_logic;
        DOUTA           : out    vl_logic_vector;
        CLKB            : in     vl_logic;
        DINB            : in     vl_logic_vector;
        ADDRB           : in     vl_logic_vector;
        ENB             : in     vl_logic;
        REGCEB          : in     vl_logic;
        WEB             : in     vl_logic_vector;
        SSRB            : in     vl_logic;
        DOUTB           : out    vl_logic_vector;
        DBITERR         : out    vl_logic;
        SBITERR         : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_ADDRA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_ADDRB_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_ALGORITHM : constant is 1;
    attribute mti_svvh_generic_type of C_BYTE_SIZE : constant is 1;
    attribute mti_svvh_generic_type of C_COMMON_CLK : constant is 1;
    attribute mti_svvh_generic_type of C_CORENAME : constant is 1;
    attribute mti_svvh_generic_type of C_DEFAULT_DATA : constant is 1;
    attribute mti_svvh_generic_type of C_DISABLE_WARN_BHV_COLL : constant is 1;
    attribute mti_svvh_generic_type of C_DISABLE_WARN_BHV_RANGE : constant is 1;
    attribute mti_svvh_generic_type of C_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ENA : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ENB : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MEM_OUTPUT_REGS_A : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MEM_OUTPUT_REGS_B : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MUX_OUTPUT_REGS_A : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MUX_OUTPUT_REGS_B : constant is 1;
    attribute mti_svvh_generic_type of C_MUX_PIPELINE_STAGES : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_REGCEA : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_REGCEB : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SSRA : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SSRB : constant is 1;
    attribute mti_svvh_generic_type of C_INIT_FILE_NAME : constant is 1;
    attribute mti_svvh_generic_type of C_LOAD_INIT_FILE : constant is 1;
    attribute mti_svvh_generic_type of C_MEM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_PRIM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_READ_DEPTH_A : constant is 1;
    attribute mti_svvh_generic_type of C_READ_DEPTH_B : constant is 1;
    attribute mti_svvh_generic_type of C_READ_WIDTH_A : constant is 1;
    attribute mti_svvh_generic_type of C_READ_WIDTH_B : constant is 1;
    attribute mti_svvh_generic_type of C_SIM_COLLISION_CHECK : constant is 1;
    attribute mti_svvh_generic_type of C_SINITA_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_SINITB_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_USE_BYTE_WEA : constant is 1;
    attribute mti_svvh_generic_type of C_USE_BYTE_WEB : constant is 1;
    attribute mti_svvh_generic_type of C_USE_DEFAULT_DATA : constant is 1;
    attribute mti_svvh_generic_type of C_USE_ECC : constant is 1;
    attribute mti_svvh_generic_type of C_USE_RAMB16BWER_RST_BHV : constant is 1;
    attribute mti_svvh_generic_type of C_WEA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_WEB_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_DEPTH_A : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_DEPTH_B : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_MODE_A : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_MODE_B : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_WIDTH_A : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_WIDTH_B : constant is 1;
    attribute mti_svvh_generic_type of C_XDEVICEFAMILY : constant is 1;
end BLK_MEM_GEN_V2_6;
