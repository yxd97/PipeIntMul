`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSOk7RK2ZdILljP1/5QH8GNVT4CdTJgOuwDgx5TMLp5j+gnwclrwAWFY6PjPjHK+
q3DlErKeBwPR3yegkQ9pGM8hhqRg8GAvLFj5Y0O6c3QU7gr9DVkD+zLca/IW9A6O
HkZTLf7KymmogGMJOcPzd0SDfglVe3wtuj0C9QzJTlssnFBEd6zDAnOcF/RhyG6x
es5CrycrkZTU/eDVwVnMOLiR1DbgE50Ys6DHyJRygIFEDaXoCrIs0L4OWZfhoG3h
MzTSF5/V/971mVmpwS1XvbKoYc6e7m/PkDRx7JHJaxNsi0qYRb+F2DaOe/ucEWJz
iUbS5hJxPAqf698XXclKdznXTgsJx8Zid3xO3BFLtwDdXJu+mtZUJTHaCwUKaPRv
x3Agl2JOSHtmN8AcKKSErW/n6swXPLDubfUs3UOkBcfSYpWYDazrEd2l9AXzRHDf
EUoh1sJ5sjAxz+icVpP/QixSMobW+j1dB1TecTy92yAxjNJeR3Ag40DmbzSbCV53
vhJUo4OWbw3lQsKfuIu9ZtGci/Hm2HrbeNIOb4OeMu0ZPeS4S6Tob8UhPs+dD3yv
UBr4ZII3oN7o81lgrjYfD3w3hFw2iAHbWs3zi0uurvONq0uqlhIlkxsnKsRxSXN9
wALWDuQva4dVFm2tbUurRmLiGtkboBvY4mqP0JZOi8CsT83IOZoNZiR12iXOIwfu
0qj1g4bnjWk3BN8tg1SifaGobiY7VjTQwHN8O1whDydn6DAwh53mnwfBlkLAgh8a
SGgLnD3n80h3AONO7g77eESqMEPlsaPshDa+K1vltK0=
`protect END_PROTECTED
