`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hk6QMJfgcCPULAXUt+IxUvl9bHJsIHuc9SE4K5W/WBeTR6+BBKcF10urdE0puFLN
VINBHh8UNGkeda2p53MiunbljlaJlimcMbHNHsXjrVSB6I+6NkvxXxsf2aaPh7e+
GO34CXy1QckgMr6eLgRvhJENdQW4oPoHTf6Ehi9mZiTuxfcP4B5RG7Y1JRYSr9WU
lwnaQ6dozWg/6gOI1IJ1XJLs8FWj0nebW183GUbuh468tzvOU7BeH7cD41wc5fLF
wc4OY1jdcGA9VrE4FrLiwYrYxXm0B3qRCzSbOzAO3Yj/eZNJghBRVBW6iwk+lVHO
+U2cDWYjg8DofTdd+CP7/fg1K4YIiIEztEZ7oEaGiJjKKb/+k6qH0xD3pCs7URvX
`protect END_PROTECTED
