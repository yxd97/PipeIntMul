`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eCd3FcRu0Tt7lG2RtnTYoj1RqygfDdtmZAA0ZVGyvGx/mOPXOCbbwmviZJ2snsjp
Wwt+SZ7A0KMEeVFFtPaEpK22IcBvwpp3t//ieWFcXK3JUhgBEJAf5QHoAxzT1HzZ
a5dIU18Nouj2KYHVbh7DUplcMOKA+PdiPltuWmtOU4itKF+jO74/3NuW4QEEo0WD
qBlIb9uIhdSriysgTKQld9aBlgNI/sUq+hiB1oJsAgbEwzxs6wWRowSKX3XToLX8
dzO0caKhfdLuq3Wf9UAc0QmO6X93kXRGZz3ycAYdV7Vy9bFQ8CdCfMlMTizwnZ13
s4JhMS4qxpNlIIXgL9Hgv+Q+PYLaUjCCcYnOeW6pMLj0BgRF1Y0FtSY62qfdeHSx
vCTGRWNpG4Nf56n6oKQYymqXS7ruBiTW62s+l+/QwpFd8eSP56L48Tp/TVcqNSk8
i9sYo6BunjYy6L1y9GOLVOk7/b7KOp4zQjjdAppb+CEVPLSFjfnzQmW78tPvBagS
`protect END_PROTECTED
