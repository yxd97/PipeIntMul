`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PzbzyAx+krCq25q4FFPIMn2/5zt32r56EyvARhrWaDbD5rOrHyjukNjfj5N1Dq2V
b/wqn/KT04Lnf8k+LocWf5oacVlIh4ScbJh9CC0A6N2STtDY/YtuauVlL1qFeMC3
TVEqhqfjNwRtonIQFe+3BHvNqp9D6Q7BvWo5UZ5gmBLJL3Viitw6oo2RSef2O+ah
nkMEw4fp82eW5HyqPz9+c35XjL0E91ZKaNtxiQ0yJI8NR3snyn2l59zxSxPItLpM
Ux8BjI2ohLWAMrH/AfpErLTpS2h/ZIrvGiADSrbWDxTaNfC0TJBJRxyqUd/Utq6O
tnAGvpWQLB2W8LOFNTozzJhyLIXnRY9+ZC0gxUhKw5OeP2YmpR8zmI9uU6TcJJSx
FTU/bWPycz8lztqc+N9anQDLTLtvFwgsoy+gcbwhNARsWIApqpQs2g2TuiotOzvL
aJKW2aXKrI05a8bGInvv5k1jjG59CpijMZUMNJqBhMJx59vnpw2Z3uvTPUS+v3hd
l2J3RYInTxO0N9nEGZ4TdA==
`protect END_PROTECTED
