`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iIaXsBrvgadzw8deiw1EUDCPOeXjc+7sQDpBG17Tm0P8JgTbAklAASacWEbtCnQe
ea8pGTwj3te6u4VPBTHRNmIzstowWz2dudACZrJ2LjWz3SvESOTPJTkvfVlc7py+
N2KtYpbOvFvahtLiKfybO1x3Q+GbYnv8Nuq7Jo3YUuYWIFFX0Y9Db/SojUy9xj+a
pNMvkT9Wy4QaXebTIR3aJ2vNT0/xAVTf2vbNfcuqBnbjFpKQi34Vv8Fc5eam3lzt
T/pfBsZYEC6PyohZygjFb6L2M1AdI+ivB8oPN0EPJVu0R3JKG0ey5A3Wiycrh/Wa
4r4eKjpL72pv3lxhN2JhKg==
`protect END_PROTECTED
