`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4AhAdeQYwhjSFPaHabaRWjjgX4KX5D7RgbHnqw0LpBSqa7HZzyiyqnzm96QTyQ2
45j2Jd0IA0yz+3TaBr8HLxGQG4yv+BdC8v9dQ0nSpvXjBEcid1ZixYJM0094mRzd
WXLTcjeSBmXrYDX2roxPBS/KbIqHgBmlXxugsFQztxULjDzyhIREfvvt2pDAkDGj
QlvDpqCbW+7WLYzXMHeLvJg2Mgfn3MR4faz+zsTKZgz/fH/TNnRkTvKg9YLXEitY
G2p2d7Z4vnoT0gvwNUQOSbpJHza4lpd5/doeIYyASpCWIt4IZTS8k2gpCNDjv8W2
/E/8J/p7Ai5csB4VaxBBmAReLNneAbW94yfyx6/dQ/J7NTHdGMKaKSnEwftOYNEu
4v6qmm2ZME15ResqQM7CA4elSE5VHcIdYpG4lEDEld3wUilF0IZEz8GvYddpobf4
if1Jh/Gql9UmvU4YPWe5EvhVc0qZV0Llt8LtABroRV/7nMKkI+JJlElvH2P1CEpB
f2ICqN3C4yhP9Yo+4YaYm7yYZJghGPEknvFsxObXPk4/i4+eL1TdyQzJrfDMiXMN
bdEbusFMW1r/94lj5YXErozAtmOsY9NiH7T5GqdaDbmhTtIuFlZ0OCWKbIkZiLon
zLsL4itszNomm+NUUQ4CwAtyEjkJZq0vzC1OyyBp5TUWQ3riX2ssLFrpGDqM5t6H
BnSWTIB77VlOt3cxg3jDtPknA1ATL19ZNTW4GjSpbbhE4t0aKaj6M5RYEHRm3uoE
KY5qpIBtmSzRHqFKc8HmbkgvIKysExnvOO8VNei2L/GeEseCcXmvYR4D8yvlx04X
N3aOTFVeyz10eg6bmlKBo42HuD+XnvTIV13Kq6jwfDSOClgn1RW27Sz/At+yhigK
V1SYxdJ3m5eL1gFqlakVGzhYlAYDA9HqOvme4YxJGhYSxK6ekXRYtPdt9owrlrP9
jpUzf8J/PvX2eBnGqkJXMKEBhljyisQgJ56mibEEWWQV6WSxu2ZGg6UzyHFkio1d
h/iQ3qOe9fzzLn0Wvbsq77cu4VFI8I5xXsXlQpSBtY3gg2wvU/5q4sa6MfIctucB
Co8Hi4VzSVzMpE4FFkVdTGO7skqRXhY5jGYgsOLtvQSNUpRULOz4UZ1SQJHjzQSn
4vFKiNrUuks+dzgmj6rOfHzK1u3FTe0cR5B5Vdvf5OGqBw1Ug04PRR8CMgIGfeal
1ndPE2YdHu02hM8ES+SXBQ==
`protect END_PROTECTED
