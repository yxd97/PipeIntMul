`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMvVwa3KSEhpf/5GoYACWzBgbf2QvkPES6ycKjq5N2+Z6+B+AyhACbosgGa44evq
TWKvHcme8zUET9roBQPO8Xn1z6nrZcfjRZWbQBXYd6oVNohqdqE0wGu2iYCMPlUF
DuomL2ObLnjZKnT6sKXlMbD6gwF8YMZGSb+RietuUxiABtfPbufE7Otb16Uaxu+t
ZAQBwIXeNsMthofy59auXHYa7v6c31pUBbfJc1dfCF5AByRZHHg6AggNs6ulscFU
8LERI5DKL2XEu+Q1znfBta1GRSe8tnawN1KddKD80oDAuJUH5HFSXt4oX3CMCMiC
7OFYZ9bDGvZS3ybrAUohcEdfhdsulHPE/SyZcbjOwFpz12QwQDBUxylDYfIhk9KX
AogS1tf/ETjWVweNBD8i7A==
`protect END_PROTECTED
