`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2hxGSYlQE375RAo717N5LEDfvwGg5Z1s1m9dihyOZGQSzoTbq2BpMjokJRQQ1jVb
l6G4FY56FsyJTB6k+TDfXZEIuF3HwP/auLyC809vWYvDAPlyCmPLMso3uCo+KDVI
4p5TIz2Cj+4wmnvoxTD58VHOdDsBMtPSADB6UDcndh14RKhEnEYLZSp/5/P0MZr5
DVMB0haN5bjrqV2W6/H71eTeHkk6UxyvWfQYvKgq/Up2viBaldVtn6P+5QhZswFu
ZFSYy+9U5x9TD424WRPHwJSxEWEnmNl6ewX1QaVTlB16v9hRngcRF+AglfuBoR7J
c9XQk7BkU1Dq5c/XYjZ7Jasr0XpewlhYh0AutB7FFqYtRB3ZiWj91pFmUlcwyzdY
VMeTZfK2DDwhRjciln0gUBHUvvPCIAJfMq8wFBEloUXizhQVLDJPVenpB+4fWZpt
1CT7ToIRNtFRvz0L9pM8QQBcOMQD6y8Fuy0dISTJrakcOtJeW/B7s8cFfzbsBbas
d0bEQ0qx0Q0e3JT1AdBYUO8V7rJe0roLWeqsq3U5J3TJf7PNKSa6djGoDlemIvVS
wDOTzdPtXBT5wgCrtBlWmprf45563rWJOGx44r8/72F0mEwHFL6FLPDUMiaySTcC
nFWfr8wbvZ4QWJgr02YnH0iv8QC7nvBCK+etBOJLORWhdbGqTtwNYIiNq1FVS5hG
C2D8Gwm4wDZ9Bh/IVogOIP/2GfaRcngMcAnAJTLdiODPRIy4g7x85ZioPZQP1f2h
XI1kKrW6XyPYPwbGpFn4v1Zf/j09Sm8gCB6o1eKj05rBwlgz61cbMjjf/yXRbY2x
dKK1CqvsmtK+aCyH1DORxEf0hvdnMOLDlRQm+Tia7IKwh0f0RJkIkDsf9LLl8Aec
OTohT4pBYGei5fBGH7L2co52EuZcyh7mSCv8COrZsHqWRqp7qbWFhGlKKeojOpBc
`protect END_PROTECTED
