`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5hx1sjx9oCDOiJR83gGOZIjNjynqP9gvpK7559c9Z06aWFu9zrITLMlvq9kt+KMM
mFpiaCr1oItsxf1Zhl+7YvomLqe91g+B9vEBmhwnjbJ+Lm9FRXQbY1yV/oAL8fnN
Wzma9ZPAF7qjp+i7VLEAjnPw9imbxdvydUSx6LaAJzfGK5/HWjHhjaJcSJUZVjuW
9mbaI1LQpyEIWpoND8narFBstOEZGOclmCjVUPw1FfgdofxRkJX+dkRN+S9Cu2rM
l/krOc6RWZHuio3xlK+PVoXPnhxbetQH7heaWO9dFfZ+sxV4U92NBuqB4bSVNB4j
n1WVLdTy4XkXTYo3rCySApfwHn1LUrqi1FxLRP08Mvk9P8ynAY2bw0+mplzPKEI7
oiV+9AuEe1voHqFbTYcCeu85yViCJQtcmco12Uk3fTBRh/JooHouEu6B9+VNqVsC
sS6OVyYrEEzMeNwqAyQJeh49BaAn5M4g5d4e9wsv4a4=
`protect END_PROTECTED
