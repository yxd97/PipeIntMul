`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XYpajowoEz6ToJh/ooaKK5zkJrnP1Abr3fXpVYxzBxK4tiBlX4y1h+HL3jU/apAd
sX1HJ504tB907q4mNa5P16EFRrgy4o+B+cP+ZSqF4rb9o3qNkk3bt7cKCOcaE5v5
RJwbc0Y+nM9yyiFMmOIv6Zq4igFhjn3Wr0TaqF5ZptpDuZkDE41fxZkYmVAUKxRS
lIE0YQKeriYwF2GKQSnoKZYZH3FBMeIT7PLGYJLeBiOvkIbkaM+ayAHOh183HYH9
QnAw38FolPygDUdZzpv9JjzexBh12zqpnpE2D6c130HSR0nd+RrRx7cSsBlg8NEz
kShzAJLnsYSzfebk49OIzPRJ0xxhRoNXhmR9R7GbzV+3aR71fM2oOnaFdU/XQ26o
M46z7IXiMuyj4TPmyXiFGGyQVX4rZD++XAsc2pDswnWsDNO0vfPZVyrlTlg9xhkT
KCZQUmwww/cZzTJeGgcudBsHzr3LPpHsh9JM5qtKEL9q5seMOEiY9j7oHVVkunFV
PFAjNuWj4740ZRXmKb4SQLttN+GyzYE3MhpOYISPVGOraVyh6GZTrEz06bZuY1Zh
mfD7jGCxPeBZjJUrWE+AG3ViT1IBnbfwjFPGxR90s60mjJJJaLnUMQvhX5Htw9hN
OfWekyNPc/SMXQw8LDFR4U9OfKxWE3psTydDv0am5bOimveUaw7a3vcnQPNvjonQ
SsIj3/leQvXrYQ1sdyZfzMvPbQhrtEeszINtBo6bLpJLwE1HGBGIcbGVzKK64vK+
dEsF6IGRowv2uImyPbvLXQsis74KGri+xcQy1NYRjSRA7PR4fo6YtK+2zA6lR/M6
iHsE3f2zaPuIQ0YsW/Rar/zdF1cQx2AwaqhepkIElZdpRl/BJKBWCT8DxBLcK0b1
iUX0HJCGixJCArQ/WrondQgSTRkB9FVkKCFksjOCPCt2jLOVMx6IySkrtWuPTvaE
CpHE4/2rSE7Ys3HzkhIvqqzDoIcy76seKeCZqc47CqvQJTiuz7KLJmwYG5TQ2mZ2
9Ms9G6wGGspYHifzm3EOIfRP/VjXt8uXHH1U8prksV6Eoqu85pmRbbvIm/FUEmia
P3azWmvTFd2xLfRane69SoCS9Qfejc5FZLdjGGmoY8HmJ8K43w2zPCjuUQCRu4g7
pOSJjI98qFOqYVlIIikEk6PudIY75WQ7zM+Np7inYpm+O2zf2cW1y8L8ZyPOSqmO
+/9gBPhpI5eG7ndeFgvJLpSNyhozGlOPG9VGJtoPUGBAhDJbG0DeGgcNsh+2eBpg
e/QxWJTAZGaftYV6W4xjOkKBkt4ckA+NT6Ea0Ooe2GNmvSziulcaWwcJBgRBWSDP
CEWYY/xVzLS636YWDsrfQhOAEwUvIsv6bsNwEs+hLmKPC69zwS1Ah8I+9Lv+TeFl
Oq4MfhR8d+Vbk+AHCsuSfIqOCj8gP8RleFhDcBCYJ34SUvQWEI2GRf/KTpVlUcIR
OsBPCETXuBjHZepy/LPjlMAcBTNCohjq9WqTDhq47lM/I1J3oJ8NITu8Rx8x6t0G
I4eKiSFnwRaFzReVpmxxYhggBCpOsE6HM/WGZAo3Uo2INUQJ2zPMW+EfpUpalW7s
hA0neTVzFLxCDPQc2lESO9mLO0VJyybXvivK8hzTQFRHkcpgddiXOoJP8PR3VW6s
7+Zw3Uya47oHKidKmRWFRUPEncuqaCrR5eEZmfU2v6omuP09Ydi1Z00Ysb9QGnzK
3Mmm2dXhelsXdoIvTOpRSHj6CdjssyyNkDdVzs6+AT4eNZ5Gtr52UU0ZDP+V7E6u
ztOTowLbgJMvg1oHBseDfU2YhEb7W79bTSdPV/IbOkTvwsYl2s07POTVbpGlqC8y
YwROrKErzhjvasYAwze0t2hyasSfi4ZBRZTadiXlf+RO1X0eoAOmWZNPY2yKgjWd
5OJKrD3N6xmfQ3DCkikH8FpBb5XpavUWY/4G1+FNkG+YGuMZoP7kTL5YuD+4Q1b1
OO0BLBkY2QY+9mwRBPfQS18etuHGCxs+t6i+bf20tMVCNwLOve+EluCWAPl01BJw
2NWUMM6Ej0aHDfgeFnPQ44bhxBa7quA77v9uRwaN0/1sPf17hAyhTJYRQgkirECo
kfIbTgw/60ZcTTfbcKyqzZVFgy/zP+Zcn3ltjgUic/sc0zfXA+DQ/X04qDue/Ij4
h3f7dRl4UZcFnKVzJcV9ipDL0XHn4oign5vN2GaZUpx/Hax9nqMgjjdAMDqaQcGx
mcISV911i+Y0XUuKtBQpGs4Z5ZgR0W8osgfvoxS+uqI/pNMyJz4h8iin2owVVO/h
7laRlAE/Y1pNARp+sBjt3kunF01Vc/cw/DiFATU0OG4kNBUyE/YmQJ5OAanq0pmB
m/F7ruXKVqUeXNjPrPjn4ot8o7fXUeYmBQR3EVpLS+TBLo8EoLYTSUWU+wooop2A
TOZ186HKXrCyDcCRD2isqQ5b+HxZpdpssr03d53FcuLI3hQHkU3/Pn8akbH4KIIE
sqm024RleqiZotuzFdzsX9BtoXauFTNs3bfVCdgkcDLznCH7MBXAapAUp4mJh2Z6
jnLSL8MQ4XxrjH04tiyotGn1VfRnzTDhg635YOXW5oZlIS49zxi+sAQu/yRoiVUb
NRcfuVzfI+xH6Qygk4EOZYE12WeV6TUHkbQBcG8ESLWraB0n37rUMtBUMFKSKFh2
+ztxfXaaVFw8esBHi+Sxpe1j4lK7qFRYIcBFjNAoKQpmDYSdbMvP1gWd/oynqHpL
IL0nbla2uKBbVFC8oYtx4RvwTvjGEJgAugc2+7JaSKuOtJRDPt5n4qNuW3DPJDKv
ILLe9/sKs2F5ajqatwsW8LHnJQ1wxiYC9/UxcajQaXEcMLGLnDYx2d7hdScgQyqq
HOMGh06Yofm6cRJPhQUCWW6is9OkaqNPzIlj4bt9ystA0YctiXLM5IRSG49DtCV/
2df8emXmNFjtz+ZnCJBVWg==
`protect END_PROTECTED
