`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMkyLr2wW5m12a1mPQYgUkg2vGfJ+zN+ThCXJpqY7LS9Wox651Xthg2zWIv2swlF
76K04B3NPnkhiEnLowDnBUf/bxlj00QmK8hm7oP9Jh1RgnomrZM1yG57Qs7pABz4
xN2gHr17kE9BAlPh3732GGZ1ZAoGMTzTP2I4eaOVQVuiI0O8DswSVwqhaccQrr/p
YMIIXTOUnuUB7J7JzJs9fmCXTYi+WgZduK9ffaAMZSEt4WQwH7AtgWpuHSg65cOD
chU1Nb4GtI5STuGMnrbsljcumv3rq6fsF+rwfRs+E+2oayuk1sG+e2Wn0o4mRoL1
NTPenemT6dMseqkZ7x0qrV+LGpE/oDZjoIiyIjrdke3duxBY7RrDVKdJrDVEI03P
YuxX9Jnragazsvr14sJC5rnUwvp9pZT2ATfXSPDFPJ9zYG4KdoucU9tltIFvGhTX
DS/p11g2WIN5aV+QjLR3pDi/gYXofRGBEGDr1u8/pcABLZ6XIOkkBqLAqp4mAA7l
hcNsWWH8BB2WztpnMHjCJryfqfF2wRUm3upgKXX3Qm9NrAimQncduOolFNFO5R2a
io3K88pkPDoKxvUvqT3FJL9DODWsIfCDWnYOtI2Xxrin2cSnAb7Q+4C2cN27Nx2+
ji2EJcH0f1ie5YirWxcex6BR8AuV6d2Kv5mF+eVOb9x14/T+Xd9mvGxsSvO5bOpQ
IDxcEoOiuh0BqS2a5ZiOFedmECOt0dJoFO/cGy+9tvaUTkOkdJoa5Ro+eEMz2JCG
gEmajEVNnuezbAOKDrlZCIM2SFMOU8/yaXBtigJuFKeBK+/WWzrpuMh+OO3RrLbE
T8Ok6KZ7a3ZPWIm2kJjxfa0tWIeA9rramXTZgEp8fMSi2MwV37MIEVJWctDBvd4i
D6uqx3DcmTs+1H4Yp91F/h4fK63EIv8hDX5fvwW1xWJYeqULZ0JpPTGT6ETW9T3q
PZDG9M9QboMX1HIcOcHfgxtjVYD0b3uqElKkxuJHgrBNcCKn91KIzuVYlJ8eaUcN
MG7rlhoAi3uUhcCZzLFHYC6acjy4AOfMIamEBlujfMSV+93f07BuLAK4/z5TX+2U
JQtwqrPxckxWQrd546cO9zylX6Ma+kbi+k3HQo3anACUkJ1es+FENTyk8vZrT4N7
Vh9wtETWMReiEZCXG6vzxUubHxyYJJHs5l7LkhGWcMmvhj0zsKDG3gP2XWX8bEke
tJw1xwZR+/Z2OKD9GzU4+PevyhU3gnklC8lLULSXgEAHml2kMXmT3JRNvHRb8dk7
Unrthm3WUR0Kvzo28Bikj4sEAHCc28xobUfs8TL72ODKRuqyLFK0ppjAiQq5CGSO
efJDXBfoQVTDxyPjp0zhWg+5bYbYlUOh329+VW0eCge+MEyimACzcZgXDldXUkHM
rKsu+nRRy3W+cTfAU3EohaSbXvTowNjMdRNy2hw6Jgh8G4f5P0dLHd8sv1pspVrE
35MGWw5JJSCm+Y9/Dm/6d+BRETkrsoyCsGRmL6Wr5DcB2tp8R5Tya9jnlLHsHM7G
msHvtDb6OQjVZqgbXUlu2L9ChtzGsH5GrY+jJJWlm4Q=
`protect END_PROTECTED
