`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0lyIGgBqJU86JBRQ7W0WTIL39RsG1Rf9FAYRpCvB8+fA8mthWJERl5uytROJkxZ4
dOyXEIeSgwbQMUlNCCwkpsjVs7ZoAjmlKsqTQ3t8VlcfRCLfKCPXN0CSQvu1VHHf
OmmVv3NOQkKiW2qgFRkzw9qft/xOGcNyF4L4Py2wP7FTpj7Emi/uzHDI4X8T14SS
+r3q2WZp33isTYlTimxuuQaUXK18nHaYOZM9B7YiyEdWR4asrDsD+edl9xxOZz2I
hEg5BHcXJCoACwjrLRoFKTTUfAwLr8YaLBo3ZQltVGPCaUmwOhr7QmJA5pFnC6BE
pde+gejGjpwZlfbsyxT0zrd9jpMu0pI4aKQ9892L/fa5+NX1PMzzysKAJ0MpERqe
SMbPrIBrC4HP1g0FjzAuYxPk6qlQ8GL3culvRJkE5iUyaANEQrqa7pYy7ZWJmSL0
O7+empXO/8t4p4peZcINRyj3lZwSORlB5kCZJXifo6xkYZPGIGvBWFP6NjhJ86Bv
TNetCFtgeddiIHiZN8G+mzhWOn+yYiGIz9YXpTqDLN7zSZ0Fqt8lpeqe5jEsw8Ee
q3BSvbSfFFvyTrQca8pXD9GRQ68BV4KlTvS8idBOhMQD51PGKHDSKIB+G/G3Z70C
tu0V/JUQApKOmTpxHBYQ9vZ+dSvNB9/T618RK7i/4Wm134VgD4gFL8jcDGN2uVee
FoV2mY/cnGVFxH6QZ1zvxU/punyrmP6Ju+iRTDdxLt193DeCezXHHn0GOMn4qOLV
hq0fD7tb70XBT3/zGK1cEc2qC2rOZtcQgnJO97xDc5rkElupixoDN0Rr+h928/AY
1MBdLGaTtxFi+DxN+VcPPtHNGYW6NMx0F/zQ9YtYwhRpcZBD9jKYm42VAs/LKiId
wnVSSdMLrxlIq20PqNjimcxQRXVXJR/jwW7A/Dj1r2WWDF+mOJCTTuoMyXkBEoTR
xDGoeStFS42ntFenf34LaihgPVPKty5ERH2bMJJgKhAdwPENuJ/wVe31X4M+5uim
OQDKkAEbH9a/Gu5j2xT9f5ithAiqZiDMxADjYItcfM5GwwXmMsIOKnvjACkdMl9F
7nfGYCuAg02cwGZaXygR4G0i95z2LKW7ym8n3Nbx9mar89nrU/mXL9Zr/8pn3coF
80cVcsws5UXsp3fwEXkuTCp5HpQqD5wZHbRp4zImPadnbrxwRvUhl1jKIFPijh0/
/ytDGrkhhxpXHaoIz3LOkJ9Azo5twHJle+1d+TIR2qeFf+54Se8r+DdhXyiur8mt
OWFRxOcbP5ynSVEF1QvYg3bN80xQ7ZDdu3WArzQTjcRML2N42RCRX7Xx3G8S4qZU
J2psrYr/nfc8J876XE1oPn2ummVFQqmdGiD1dYEmtXrT8QyGhM9AH+VdLpeT8PL+
45IIxuquvBsN/fnuwmIJlLnqiV/VUlZ6i/admBENBoCKJRQUg9zDLTPOJgJCldw8
Nm1MhYBbUSungP50/680hHaUXeEVAFP8GVttKjY+KLZq7AniNLN4FVPhdIlBAE7g
HR/fkwHih3eQhYnZVFUZ4W6BbVLk10QIYsKabV6qfpLCRNSeMS8dLKpIrfXPFugR
gMzttZmaXE0IsRufONXws/K1IY6Ls709WjdBCY5VC9rAlMgJUNtjHFeH6YkuH5i5
tRizdXaw9ctICMY8KvOadfp9RjqsXr6KctfQpRUpn9RjMfhLOhmW/Tjq53elfw7z
v1UGzPfXwgEIiCETVVX0qZYJKl1DdUrb8c7vy4CoDkduan1t+ZXKB7tPCBPhQ3ud
O7tBanm+TzgEp5gxkje6g+cfvXrpVVayUkTKYfXfx6QMnq5NIObY1ldSkJzRkwMo
8/IcEoSEIzgieuwaDdy+ZQsnq69Wrp8DehzNaKz2nZohy1IbbiDFug7XCOp6PL7G
pjZW1CxMwzpbwXdW0Bgni37xtscRJvNw+K1NOK9p7GKot/VqXp27wfZmgmDPNRjj
r11N+kamCwubzyAtIWmA5ONntUg0DVhYPY/bmeIXpgMkZS5T9xwgqcl/vg3wXOBF
gbM+PMspUhvoBeh7StxmvgHCtSCl4AwDrp29fIx9WIAF4xPuBtp6zj0Aq/yf8n6v
Q6RWxHR3C404vaFD7wyWk2rV47Wj35sfYjfD3c/rTEn2xV6YDfaSVd2AkKm38nO4
hDogxr8Ef7EbpbSOEQn2IA9jms2YfY0Kal/MTIAZ0mOdIbyZ2IlSRZxXHBWtoxmt
`protect END_PROTECTED
