`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exhzUYmJVht6f6B7W7Y1cttvL9TInvuTIjyJeVqN462HXCDOjEz5uj8cB+GML5Lo
KURyn3/7z7S26eXoaUZLBX/yHgAkUFUZ04k8YVmJL+RmheHKl6qQB9b/KIl5TWV4
s+12DK1hkS784bsst2kUAOXYvH6MG1d/4rf4xiztJfbgwpcwNabQ1n/pxSwnQQPw
rfPyy0j6UloZ7FkCc/3ZlWgIqBtjai8FJZHthzDkDrZzHDYntC/sSaj85t7WTLLS
EHGGXq9mgNTjMAd7/VnYbAl8WCV+d0NC0SJcFQS9z7jmzKFobGkW3rXJoCtGqRWF
5Vt75LiPLCZaDHtql7yapw==
`protect END_PROTECTED
