`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GEjDoEN4za3WJ+pVr9bFjFR/JfVUWX1/95SvU+ES39VLCRO8yOiM0FQf3CT8xyLu
LG8y3O3tPJfHjeCkRRDeGaoeGF0PPSm48e3l8xgoDYATA2cNcQpD9PvS+chBJpiq
OyUyMP9rJU1PFbo8QHveItfkyQ7i5ES1tDXEgHvovsKpBQhyL9Uw1vL+Zi36Bu/r
2KTqJ8206IOyfVBw24XxfUs6qyRhkjK/TBWdQbt2yUeYkSFPOoeKPpTw5x2byK6a
8SBu9DeuMgUIAMD9nG5y/9mJewnQBBKaHlnW05nOY9ca6HhKLuaRJPhm+ODUPAZR
vQfnNbUR7M4U5nDoIkR1sEgfmFKt7O5aNSXcXh+zPN+iT3kgxbWkp9m3XTJsZ0fY
`protect END_PROTECTED
