`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1KJiLaVxa/ycq5OzbAo3a5wskT+y9XRMrSQq4fOX/emfeeBGLHPGTSwZbviarAko
8RBiKos201OE8PXbNag1GZqhX/btlsULSeNZ1IeICdZr6UYG2DLbs709NPZ7VIIR
m1EPmZV2r+9GKRTvIuZ9agEoTre7l/qlrxJR6RBgd+6yuW1tyYpHCb0ma+f6hKQt
jbvIaOrrJLfJrOj9w6VF3+yoaMDJsXB+BsIO7vpG/CIsGOWSdjdBSdPeOM5CitdP
jn8l3RA+pXS2HpNMmqAa/DqbcgQmoeRxg9BEITqluith7p6Ye2N/y/BPkzf2cZVT
/AnCJVJXHQQzKXbz4bVqm9+BIxkLfjm9klRgutBXFVkphr2ZIXRoxkUccu8+N+Ud
2mxwRN87O+tfbsQg+xZUkUd6vkJJ5cpPapsbXFr4yge7tgNDKRdSSMmjF2oT7sNE
jGcmoR/oj2JxK1H7pDW0J8cXO3VNEPgh8iLS9fAjBf9y/IdzY0wXji3Q2tFS6bJm
kXeNRHSN1lBGukOk6dnCZLlr6ESVTOsRlT3bHgfKBGsWfcaQXpCHhAF0RqM351ls
LGnWtw/Owh7H2wKg9NnZ6Wj+dhhYXCOhXG+jAjWnqjbabMv398yvRMZoHjuGS5Fu
8lxglZSqU1Nh4CajKdtCkVXKS6UmKwKo0fQv8GRLOlI9bgsVVjARnWvH3Tss+aYi
pr+yVNl5i2AdcCv50G9laCFfvrdXm1ymppvC+6BxA225kdzEO8fmkKDq0zfJX62C
/lf4UP5+8KQw9XOfHFgm7b5w0AxIpCPPIwci+f1Rpgu8945vn8kU7r0AsD6qx3Pa
J0rGDNcX6XdwnTZFycuKiY0L52i4H9HVM31GwsFizhLovN/xj11LRFggJf2wqy8f
Cv7dlXY9kDmS8Q2mIbaFWrBOZtZZMlrZLmn6In0aCgfCgdoJTWa5/WL+qfpM+uYo
M23TS23rCbOsWkHkO2knCFuGngGmH5mfNxf77gIpn5VOPQ7DAeRv8X2AptH2X0Lf
KWopmvfx8EoYOQji3J9j1DN08oxEJ3QlxPNQG35Qyt63HLBgOmWgbEpREIiBXqsI
`protect END_PROTECTED
