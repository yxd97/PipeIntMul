`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c60PeTBTLP9CmReQ6AZPsBBl5YgQ4Kk0MMkZVSvmNyBXNp+TedHgrYwrWP+A2KYa
KUWMOtHcpbBl3CibZWtRE2WP8Thgz43QZSqYXuSgBNE0+rss5EyFBjAhl+0es3m+
mbWuhe7wd6ClX1aNnT58oc49pbYoCSBMIqErb+XdCxK81IE+LPHdQu8apNLvM3UQ
m265NKNtF/+LNj+oth2yPkC1qF4MZ9sHr8ED5SaPjkET3/mSYoWPwPyvD4mrlxUc
yofZHOPLjeYQRxqUmeJEQ4AOuY2Y0hS7QBqpu7VfSAMdzGL4Db6TC3hMD1rxynuh
QltUWt38hu7xYHAytSLWCtSU1S89Oeuw8uRICgAJ14CwYI3yqVqW3K6CaG9eNl38
/GM+i9PIfxqDKm1TdcWkXqA10RvkUtYUpjkDDJJGLUanEU+3ghBuTAN9P3BG5TCp
iTrf5iq3qBmuOHDBTV/GjMut22bl7CLNN3/s+5AOeh3MN7z19eupCT2HEXaQGfU9
lopRY3V6KY9k4Zw2stf0LXgeXP3Gx0eO0gCfohD02igmWxH/5i4XZs2l6rAF3Yq+
qOOiieonp8sUxkNj8OAhdmcps35lX5RVRTxvXhcjrPzRH3we3KDMJbBSZDg7W46X
s2WMdzYMW5k+C2C2mSA7dEUQVZkCxKp3k24Qvh1qR2VdfA/yd712ou8Ij17zOtFO
3zdYmV0XG/2Ep9qpiH1dLXpUwZM4h4AICcaFlu1TpwvtZGirbd7YmLkdQpVteVcZ
xZDPQoEiwQ25OqIfvLFQ/PF/t09mqmgP1BuwR+v2GCKwTqd5VAdTaKHi1jEl0T61
/Husy/tTOC7QJJmHcA5S5l1e6JxfRXnceF4jyQR6bCLWEQWoHB+bq1RkdbsjHGvL
oQ8Hx/Eb/5WcD/+u4iIHbq4m/Kzmr3nX5GizPPbK6YYk6uRX7sTzvsXD2sfk7cj5
jS8vUUXSDY056phJeYBOLj+yZcqjer/VfV0LAtwsA522V3bByNbq83a9ohhJ0RFt
5W9SBT4u57+rcd2LXuCJPSraXGlqqiCeAo/4eNwyxnM3ZJCSW2tG4iI7ESHTFsWy
/qrGfTn6cfkeZKqQ4xmH5n82sH7nVBtOmjsigcxsb+iYEAY0ZbRftex/4xNZfO+0
5E/yRT3KkVdgs0BE/6AiI/rKuF1Ui8iQkz4yiySKmuyfsbzMmFVuPrp+fN9+g2nN
4pM8KQlotaVM/hEv2wrGsSSUTyCqpaFk+cwHMoQ/rClcwFpE0bxwL0+oMLNw6U54
q2Uay+TomzPDROoqPIaRok/1sJEbrRqhnc0mUdybJomb4Gq8LJIo5Q8nXG0Qca8c
/je9Dv0m91JlVRT1uHE8w6sbMAq0necsMyQ9I7P7Hw5bo4liA10Vp8LlHxlaiaAb
lcR+wbnY81N50Hg2GFXOc70eOUprE2ZpGrbIE9ZtudsrKL7bqNqJYdkYlVwmJGuH
9O9pcf8xnaq+8iqXB+Fwqi5epuz/YrDYe/t6ub0M2JU2qJ0UD8BEeNB238iHHPnV
fT243YPKFAE1xMrZoriDyQktqK3ZObGvIJpyfYMyt6AbGDAJBpLGoGQJ3GXfRb6h
HXWnbIy3rquBVmOHSC3DtM04lvffTHEbIhqT8lBFTErGbd26MGZC4uCEVMhLyXQb
l+tHxNUcaw5TL1Ms7xpEVh/SH62xDG0k2sKRb2ca+QnRjA2gZQmEIghZM5a8CFT1
iJV8lCPStn8RZpH3ZRN8ZsdFp/XKY544MtJXy2ZTLHEjwWiqGJguWgWxMcjCbnrI
U9kyer0A/XmOIxRS3rhtZ5p8tV0KMq9+aFdFkSNjwc8DHnvhZuLPtFsYaup0CGIA
Xy6UsVAcYvHby8Y1bkPiqDnh0yVW18hXurhyHmPmQJQjl/RdMwP28Q5FCWq2f3qP
60H/u7boiyxQJ05MBEArMwYjDGHUDxQTizP/0PJ9uYCWF5pgE/51rS44ASqjPmHG
ulDVIzTIcIjEQJ4WD2WN6RbGAENUNzJ+xgQ/7Iu5Dk3kx3OvIq3bY6+taT42kQd+
vTxziQes/bDc1ksKhKHSEqPWMO/t4X71P2qZgXLxBZT7Rjf9AetQIAhW5tAabG4p
vcmpyW4iZ4YYpGvo3kiaWTyvWb+BqSFiLup7HHenlOJqkDDEejosNSxptGGvaeaP
/EL2uTPy2PyZJ4CByEuBIdXHCVUcsRymwVIYqj1SKbKuRKxYa7m6KZJRu9e81JmY
OsIHY1eIGKFdwy53vjsVLwy7cGe5avCStKHGq0IywOjgsSSnuayfWu2S2oGJUoD3
F2jsqOUSI3Rk5nyIqtIfE8rzOM7vpI+h92cZaJUnXZq+YuqrmOl9DuqLDcBPMjfl
2DFup7aJUhkIBVCbPQCZSrMl0eyEdgTlnU1q01xMIUmQXGpKGljP1vBNJyeB4x3t
4Zht7Ez0T+lyZLd0/FqPh5mOux0uirIwWXKqqLiw5RJ10s1NL9ldjaTZ+Hf28vVn
VUfmH34fAgsQInC1IzoFEh/7cbTjHgyRrj0fBYsVoo6YaH2HjO77wOsahWX7E6vm
WOlYQ6m+OBYANB8+sVrAdvVYZ3VKor1l+GC1lj1TLu8c5wkCHtvBXENIfHlEG4Lu
hbHkvt6JdWog+lf5B60JQNOzWK7G+x62KDqGOU3FibYDp1per/nf31fI4xkz9fDp
Q6x6opnFZSLsw52uVqmqVrmx0EkVTQPz24RI7CX45p53MHu8jan7gRVDHTL7ofV+
ZROakrwGVIavrYVwAiwU3sfPwMgp1Fz69bdxSi7i6SwfOjQcszJM07dbhU5MFNne
CwVSEDe686FCr7vvt/4JlvHFVhcVEYlTlyfiq8qTzXyOFYjwsCmrmWg1hgpWC48X
oPAwAp4ckHODV+Ggdll6veS75uQqj+ZLXEgmKTuIweG+rgCZfUcAYxK1jP7VGoxv
rDWsVI6C9Vx2kGhhzcP6bv0pXVk7UAr9245D6wgazdFJ4cXUUxPHBe5kdmz7LNql
F1v00p94ih5HA43WDY0mwsQS45u1F9sIv8WR1UDAjmLTBJGtieOF/7ZpN1xQBr2y
1qCxdNCqD+mBaRt06rmcOR5+lJtVoLP+XVYgTzN/Vfk/A5WB5myn2wqshNZ3YYau
+zJMAeDg3h1BFxuJDB3VgFzUjzj+LRdP6oD+rNYh02qbe/A3st1WrSCQG/6D3b89
K4NWx8z5ml8b3uYyzvCXRscv/5qGdaWOu631CO5PyxySVqgVbeEY4SNFvWKjxqGJ
l/uO+WVA8H21ZH6GqOYjVNAzziGA+yl1VoNbjz0tHEAznKQwhww9Y+xS3exQSuWf
i+Kv5vFVOYyQVD6TN670siMWWW+nyUueefH2knjLQIWx6QdVG5sOFrM/9dSNjnmb
hb/laLQJrw6EtqcFM5n876lWvU+R7gKqD/DIvDfURj7kxBAje1X2q8OI6C+B9fxi
EaaTT8kGia8oRb9l3M6VxJF5vSzFab7uOxchToiMe12zpGZ9AuKCHpVrT1EytDiF
X/XaO2I3HO6W7AQ4iGQWHFjd6zxQdB6i70chONaa5MpAfi83rhUaJmMwRACeLxGK
iFP8Vhi5zBiGAieHPJRQqZeG4oltcuGW5qjUCPmql/rYxce/r5VZVES9MPSr11sU
CMqjJMnf/BlwgEAeLkrYtdOT38KTl+pdOFf55Tbg29cGpNZ5xQyVs1DW3kEYWKPv
11P0oim8EV3NM4SpOuV+f5v5K/ZOm53uU762a6T2luV6E3cVcySbofMjh8XvPyGc
1htDQdXQVtTO8pDS2ug1/MR3TIdNgO8AmchyCWEmLy/UMGV8OrUIiBxxCzgHF07V
Vd6bWLPYkD4wTPcGhRTDvA+/uavubaB/uhm+4D3dU6H8hqTm6OkqdCO00UaABG9Z
2ORwrTcdf2gxR6GvTLrwjiIsXa20iVNLxS89O0ObrMM27Zl7H/emNroLUh66qSMO
lmCAsDIyV/+VPaESD2TBDXRqT85NxJAzuH3Q0Lfu5kQnbs8OfFn+DSx7HwR6c2hj
opokp9cFnhTJChKdLEASH97lMv5GGrUWGw0oNnkDWymumaZUSEoKd4HqaXsl1Ryq
XcEst9+/W8mI7RHB9oKyWmAq+VNmFqHJAnP+kGwOt/LEv9R73SVrzq+nNZxgiOeh
V9EJOn9bOtbHVaJJb00x2VaOXnzTj4DlzSp2lWYDFFtYEIZ/NTm1GbHq3aPs8RoX
G0fFx1opTTKEawweQs/4etB9dN57sa/vhwnF1Q5CscagcTqxlpmhottnbG8ymxVZ
ip8dVDJ41lQbPjNoR6roEJRmjNbfrqqi4ZluJhewrJj0usLcEiZwnbzR1aBjLfKP
Jjv4CYILyKY76Ug0Y26bhJ4LdWzx1wQ+I168rZX4y1/6gKqxwsudi1tLiyi1cot2
7cCsub6p1BGFDNRoPBJJNFkU90Ybrub9lgB4raRHukLBfQD9wzunBvKvvyLuKeKC
Agp9uyQtvdGtFHEloUCG1al/9UPkA7iKmRbrAcj82qk27y36inV481J+SERs5Rwp
baYPP9KcNSqJ9TvttDFzao5ELX3seote10Votsd7iZWWGTe7+MJngdFv+KjFv2Tc
r93046rg5W3/BnpEUWy+uic491dG9G1GAHs4/LxZeCWYZaRK44IjcD8ErPKhRCvk
N5XiTQiJR5oAeBLgNp2IdK9N2YXfmVAgPTjT9IL0L8EpsgeeZ6h2xsGUR9RL+O9H
JlRwSbr+CIbOmHVn6/1zZl8QKQB0NSbNGqxs+hTePtuYI/jAm31M53+/4V9rQ/FE
CO4peeeIXMzIPrbLKg9K9BvWu2vBYpqOCcwdTV2EOL80TRfzF87lxArh/WDSdIeq
liRPXtRYz12EDljk0aF+x4kSmQfRx8ZqgmobrKGFKUkO0uKxJETmEeWAVQywQJXw
WdSI9bwQTZKAggMOMsbSLE6NAziHk0ntGsDE0TnhRzb2WapOqQuHeK70/N1VE01T
t0kFomV2yTO3qJZd2SjIRbdM62LhT2ImPTKK7ncyeFKwoDUjBefJTeCQKyglHqw6
UGxejbTmQQxqiGRNo7YGBEpiYdEVlLxDZ848cmBsjb3B+MczMSOHd+g5XqQl3XWe
t9ScjT4aLxbuQIbBfmQ+3sqwBjR9mUJeRxCBtxvOG5DEaxTIzGVpS0XAqi3Ecavp
AR/y6Et4Y4MJgQomcVXk5/mp9lcEKxnx3nsObRYJSRsd24hEEORjRxsRE+pp91+0
Ey563SIaAdOEEgXRnOV3mCMXCRapiIhzb81awFDDJF26BvFtesbDhIGMHaEXoKzj
/7v21rYX7vDImTh1FqZvsfCslGRocaG05ohyC8qb5TMamlTQhveYJpEq4lln3zVR
VTrZF4JSA/AG8ig9uBBHD5dw/0tqrzT8aVuEn9dRaNAhrKqSxqKv99ExS5iWZVXZ
jI5EkWFxiVS2xcczxIJ8jfEXJN49rxMg1Im217oBglKEo4jUaWHzqgAH/FJ3O538
JTXAttr17MefnI6UHQmBuRX705div9Qi0oh2xDasL6izq0o9LE1hlTLwlt8QqmOi
y81G4Go9HB8XVBE6TcpjIk38YYkyLqzYqQ31vY6gAj1LfWXG4zJQvMN5MlscN+fV
7IGVFO7wEJu0LRpV8JZ0fNKjZhDTcy7fhdlVSBPAnFSdIzkFowxaHOEup3NQq2C5
bhw0ogVX+ErtPxUmcA4FrCQdPEbfknMJhPDZ4Nr70/N/hvO2RVyX4/54WaDsr1Bf
0b1vdT7kFhExhdMI8MyLT8KHnwdl70RTS2fNzdwPqFIh9YpziUfossUrtmeGFDyh
7FDzeqG5O4/UoMCZa6I7HkmjCkaKMXJpC8yyhUZx41dzKCxS9G/0USP3viheTZb1
/Q1b2SsaWmoHClgbf599OQZp1SFysPbLrhEWjd4fF9fNvm/x/XVlnAy4od8U5PG9
Q7GoPQ6Hq6HE2A5R7G4+/T7gYodMmGmHFWYsUeQmAFjfUDKzJIIrn83O6XHRrIjW
MXDQLsdRl9su1xshUZoRXWrIDTkNwfJhiG7EP9XlMMy1Q0xkvPjp8ZKV+JQS1n53
oo9eZjnTYZoTnsyi6qtOBXATYs7FXScciPaTKZrN+9z62/HQvZoZKdwJFUJlK8nO
X2alrVZiAY1amzPaXMoS1FjQj+udhnUAbsvbPKW/lfxKf1tfEe8VCkz73+UzPfJi
GRvUdM+fqlTX5SG+xf3E/MM7fjSVDb8nEbirdFjMZMwbdPba6jokf+NXu/yeJqPb
mvRgdxAfjI0LVtCR5gj1K+zJ6wDskfuXoRUKLTu7VUJ6E3Dcb8u+GX/lKdg2KrxZ
pgPwjiJp7k5d1J8pXAhhF1Mhw3Ak3lhw9kWngcgQD6H/RUfDqWXpN03ZiBBmbw5Y
BXTVv6IyzY+S72TuX7era3jirhk60JSLBNJ5Q797mTMy8hxiFWXy2wziM0nzES4p
UPMPieREFvAPWZHQqXidcyUwFwDJxDT3U6x5+4vsKIQQooc8AS+azkNngQx9Hq5/
cKaXldVtPV8UR74VwPmlc57qiMBA0Yci1a46FpS+RhOu3I2hxtkccsMyzaPWzroD
DcQZN9IXlo2GgCdBVty7D3XzCGKu8tc2E4S+8zNP2Ymq5Ltzwiu8q0HzF8eJFyki
P/BUpXQU3OvueNJuJYBwfLbyE0igvkyUXRaPYBBMTNAbspyhwHHrdUAykPAK4aAr
Ppdj5BAhqvkL6/Y5wZIL8OCjug9XI4dCbrXuZasLtH36fftS/NvYazyTfRQ8IMGs
XK18WcHECvIhj0UdplmS6HMMvMNAdH464uXmHpbUwkopX9sAR+isR2yG8S0leTiv
N6t60C8cFbKxKe25hszZpgcoG/ZZsvq9Nz7uOFIebU1JLJ2mWzThsmXk7u0WwOx0
IUTRHDMEbV4r8KCUWnUIxgLkcDe8asPm42FXtMe5S67KLtEPX5I18mzU5ea0K70g
62TEMG1lXETsA8KRRzThoywi3v+Nr0nClHVOI0JRbfDS/0t74FZh5ZJHQhYvD2xk
dRirQYVQv++eI/xgP+Aec7RtbfjHjrCCPABaDUjrdbjWclVlLkQwkVCh93VhUiTf
6VtaaAr8cODgjROQzirJZf+kbpaPmnhqlZ9wL+f9EsBMw295QanpP7iiTXobYU3x
rYeBKouZ4L//ussF64Rhc6z5hCWy7Xjaim2gyNmLGAxIsOXfuLsX0eGLml2kmlkx
ZUzxnsnfqguyE7lOj22SbMeT/oE5ogNi5hMJYFSyXboGI6OuRps3GcTAXLb+Mjre
k1D37cVBcytef4UxG4XeYAeU8k9vQIaAvRHaeGx0TkdZkd9YKPnHLxToUaZH8PRf
BsR0JrmUGXzOPCTq2kPNBvd4O/Bgn+K5UaYX22Mr6Eda3SoUI9Ogl/8LIWLg0Xs+
MWO9zXFACHrhfnRMeEyqyawcDptIM2kffB8qRngCDqcWbnn2KoB3ZFaym1TcvB5K
k3To5uMMYz5zrELqx4sycfEpD5Ys5loHMY3TgdEPkAriRhORPuhzAtV5/eqBJYq+
zaGrmQh3N82Nu9igqxsPqgAq3qX969IPQ62kiLkf+B3qOGen0ereF2W0JbbOCkyN
vkk15bFFNfnvFKjB3JEhjNEQbUuWuwNfd+2+Qci8qg9o/CGZpI5Pzazv1Rx5a3uq
c2qd32fSA2ftATPNsQaQDB5SuAw9MKgX+DrFO6JW/dY=
`protect END_PROTECTED
