`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSl/6WUPbdZC0qF4JeYbpMROXSiupSk+OBf/Shh2XIqkFR65/h8q6trWsG4BSkdr
NYFgfkNWB5U+MUEA5SdzofPSPtSIQLfxSJRqL0B5rpOVLInQ9eOp/w+b0VZc8VHf
i5LVAXvQ+iWhQouh2qxLa1ale8jU2xThfuSCiatGou5da1ZBNg1OogdVHuVSmm/s
Veszy4LQa+sYJvLnmgeWhAoCngRhfj/ae58YyI1Li0Ni+aUM2td6bkeR2ZAzeLD4
eCW7bhlID5lgNRYaQ0iQdDMvnG6gLqs5T+TZU+0pd5JbXD5ufqj2jGvA6acMLwkj
fNSk+0sVZEyOT0HFdEFFt5Dk4Dj19LYLq1ag/dD4J7hL1zbmUhdVnMahxowYDeuz
sNmNXUPOH8e8Bot84Q0CrgRxA5W7Bh5xriCbnmXkw2MLQIwQRm9GyzmWVUpE0tQo
NsJEXc65O5WQOW1ImH+Je8WJQVTXSotf9C/W/Cmj8/qxRYfxrONXUUGRlMeXl7GZ
5vpIxxFjHfzme3n5ZQYfaPICbkopyMkPJ88pC47Y577kL0NFEQ+hTGGwlsl7zjor
ou67Isomns1KrbA6NMyRQPDH/FZ/WOU1etuxs3DKtPkHmL+3vAF/QVkiSuuvU2LB
of92Bd2aJ5oPpswXXP3EJEEOfsbvfgBiT+P+07SZAnugPiYMsrRfic6IUMkwCQQH
xfV0deeCzLSaNfHs5ET/+/F0sl6U1sYKBLYTpt7gcAE8rL2MS5ObJXveXavCNZew
SQG96XPCs1OhJuBjUmeVZJV/RIpHSCq0mwjgiZ8DVPxopvk/ygHz7DV3QSvN0Kdb
hGXClz12k31fE3qJ+r+ErN2dPqnILuZ3zLhCdZduyc+pfZoUiKAxsa/oIlH3PMb/
vXJfSXYAusOXzKp9ROrWJOnD4qvT9nHBJ2ZdzlU7Xz2MCZ8HL2lJpFFgL0rFMsZR
OocshSHPyiIKi9njDadz9jCOnfh7lCvMVxHh/fxqsjyfBbEKyTNApRRc204kCdIl
UGwpS8aDeR5QdiB3CX8roA==
`protect END_PROTECTED
