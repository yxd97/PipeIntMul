`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+Cqb0IKiiEG1BN29Ej9B1D+2IpAM6YN7m9lKDdruLxdqinzgczu0PhloBJfBTn1
+WrId1OPCUQrhjzqKJ+Jc+jHn7W9O8FlwC75CRwQbmFstYJI0qCxeSF7zDQvOTiH
ILqhsykAeSPc/YSAmHSVN8+gaBx6D0QL+WXERh0uj6E93ZlA9mc271tURkZ0EStV
1nywdTiYUt9tWra4IvXq4jTjW6sDTe+qyM3naL+3QnMP9H38UAK9B29x1JnaWTQK
TPzoV8IytUdR7L4UksiWCcooo0YhTKf8aG7gSjZqcXpxtUr1lrkhu0L6kRSUy2F/
eWHUfnVCPuPRBOMnce+SPsKL8dHu4R1l7O/1EKnFzG0=
`protect END_PROTECTED
