`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ilsJ4Pf/iLmju7cArSsMQ1xhdTN0nymrCnEB8JCsKKgG7i/VvA7fZBtMvtc8dZtF
+RU4S7kn/9sRYbIe9lWkY9Sf+DiOTmS0Sbxd4R+aJd4qj97/Mn2nxVHQkR5ZjSS5
Q99KixKl0vIYxqYkE7cp3IrzUzc2G5R/AJ20iSTTNOmqn2X3x+W+mo4QI2uhHsg0
6+QlnjAfnjN2O1m57qWGJjUfoHKTktWnAYlI2DEthzYmYVhN/vhKG98QzbK0AUSi
HzHRa3dWJHlsYr0mZRkjx0VJAtUjBmuhGf9I1Sv52hhHpseEqTGVcGEUbOEmOooA
hUZMtaNuzfuxKKI1m9X4uA==
`protect END_PROTECTED
