`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nt/UBTFpAy+HeTbVrUQltOR0kfTYpOcy9qNuDbGFYryqwu9VF6xvnrL98dDc7mFH
6lokSM2uFkeUAlRg+9Hw0vvGOi9zKuYMuMUOeBLQCWQY1f6g+/47dow6YSo4/wU8
J2Rwa9Ojnw/Bjfw5kON1LaAYfObuERw+s2Yr/19KSYt/pvDEsnq12R8UgXwmNCyu
HrxemfMsY0aZ2YSFaPCzR7KnpC+mAI7Vd8mV7J+d41RogdHnZPCA4zd1HGV544n7
Nv2mGlV19oqkVqkH2MchzKI4vDDHdEH3WgkTAkBu7RuCq38CddrZ2DO/T560EROl
NWQTQLguncr/5UsilqXyS3h6oPpKTZYiRA8zpg/HkddRNx5vJrXyBtTU+4XwsgIK
0xbjGgOniKLMr/W2ItTJYg==
`protect END_PROTECTED
