`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0FJlkqQ7pZaHoI0m2OqZvzwmMmKcakcYIcYOsjA+kMegTGFJ6n3eiK+9k1lCUrDg
nDOghiwnlXym5fDsq2KWoDGPb/dAdG8NsMV2e5zVfCaxS6AMmG04+1jh2TgRrdA6
mf5dWAMrbFqEDbyl69TJhkhVS5nVhP0Cql09pAOSC0Ljjn+qJDpd+hNiS+Ft2TqS
qUxgAwf7eF+Q5pm2+fRdffSNGNJMx6JIv6rnQwiQKNwkKi+WBt5v0Zu0sgs8CUNG
maWXgDWyDlz/TbwrIrOrBd/AED7aajF5Ro/TCQgPILvbjxEahjDOcggud5jUYRtb
OFmEYjWr5o1LVzO3sO2Je1o8YkZjlPFsm08jdkxH5hXJUL3VwlvszBqQ/vJFmqnc
u0bS1fSAtQ3fwtmGUy1DwbYoG6s/3Yw2FMvbPjX1l8oCCgNz40UDi83WTrUokLpy
CBcS2jmIdRo1ntxqM+4smV0VspYEuNpXha4qYDlFueV8f+cqO7783Mz1V/8n85N1
7oFdXh7GYRHNWS2k2mxXo3zFEDulySK9YmSwYPNrrOwojMFYWrzXGRhg5+PA7VZt
pPg2JhGyymUIS7QvROL9ITMfXNzZ0497C66ntnGOZP4hycXl/1w5yalDR6zo0cpb
8EB1WAbieKAqepjTyw4y+jBv+UnEZsfh/gELyaCG0AY=
`protect END_PROTECTED
