`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EBjtEcXosmzk8B8KxLPfdLs2y5tPTWqzcsFPCSG2DnpOv4JN5rTiecnW2NwldV/N
nbgYiR6gNVOZGfhI3x3Z7ppzvmtg0BsXN6hVf0Jp8/8KHitniwGdyBALhtZS3vA4
5GlAXS1pyc139fR9HRhgc7h9YnYtjmCPc3hEkq9hc4Pi1ThMYNrtfU8GqVJUOmvY
6++2YdKDi6hLVrG9Bw6mhvGkJUcDPEcrSAABDgWNtjVhyhZTDEp6NyBW0I/qBM/G
yZUR1KyvTW5ecpX9G/clhAQkwhHJz1Xd61OljYQ/kQYHVv9J9LfSFgHFSMrq04EI
ABN8aujcArP50IqEQOGsjSt9WtI/xfCmP+bBvlsAEVQ8+RJwmuhqcKY9q47130QP
RL9Wh8+2/JRcUGNIEJ1GUFFdK1mWT61DN4M9W37ahbTwQdX9fMkxuxtdcID4eN1m
N/UfRsbg116mqVHKVHkPim4bEtEe5VkdCQNJuSM95mQDk3Br0CSHspDwECyvut1G
B5VDAUGQH/iHt0UVwmiNFqFPILWregCeAy9ffXwRc+mc8XZv87wgA0ZVabe1PLY1
3BF9CpwJI9+86uVZL6QJV9dyr2zBe9cwqxy6oG07gkiK8rmsY0zOumzJzWQkTHhb
FJTBYvkzWup3SZIOWejGzUvcbyOt8BIe+JENUQrxktI=
`protect END_PROTECTED
