`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxBh4LbB0kDKCIwnoL8icEmbYTUStBRh09cJzOyMvoFjU2ULh/OpqxoeBGO9CQ+H
OT5+y3OojTrlsJnUp/PIVJN+JPFgylWrDE//oiTL/7MX/Iv+nX/VnaGuXFn7Ginl
A5PIYY3Qza6N/hhBZ8K94qMjEdNh7UpRCbDGtcg1x18o07/D9ctr/2Tuut9jqaSk
8Qd+z69N0THLiALPjCQbpI0CV4NJRKZmL18AHCjdrBW41sthQZRDKma5O8IbUlQS
MQDBLaKT9vfknHBrRgifkuspS+eSt12GRBpi3j5RD7Jr0HxAJwAxglxNimV2nDu7
+kEtRDEsUFONKf0SSB7gjNmtNCzjdTMWw5drp1qRhDfgfKQjQLotpRLTkVLJHkho
5jjOS4NodG6We45JZWnT49L9z5wnPfZmwEs5sN4owXcOD+KWwKwwjRoVL83bNWBN
gEVs6fpWDLRby8UH10kNYg4vhOt5pJjk51UpcFWCB751my3AX2MIkI72B/ZmrKL+
`protect END_PROTECTED
