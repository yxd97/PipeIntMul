`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WcV4TGaOb3gLMUcrV1MLaZD2AbVjAfmoQKvtGwEu9ApRw6QiSocWEV25flUhfPGE
abZRXBghEF4topmxh64FGQQpJYat1Frcc4YiXhKLwqGpgjKWofjj85nw+I3vGCJ+
HkdWeqV2+Iu0p2RJOzfjKvNaVm3GRhd2XmIpvaZn3o7eQvrinHNJ+Yzl2qKVD8HP
3HY76oW0igWFB6cbE5mqdSFk2uAlvvcRpys2T1a9OZDSakJPvLe/vKY+vb3/ofzt
bcQaM+R682wQpL9DMIHs58nb9eEUwN+xxuJjV5vyizrG5YJ8+CTDntfAvH2wXvmA
+02DubmYW/xl1Gw7/Y/K47+NuAqgIfe4trLNNlCfAwProlz+y1h5m03iu9+56Stq
`protect END_PROTECTED
