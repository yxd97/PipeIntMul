`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gexkcgj0dtB+ou6/JjRU31rPfDduogjKTNSE8RVU83XO3qtytThfM3FnA+c9Rbh5
wp/vbnQjjP9zPrUkEKBZCAxCx90jeC9/6i3Vm0ckRBgL2BZSIvchndli9uxrKfk+
+IURkKOFpMCt86ustQ3dvBLDdCAud+lkp8SQN9Ie6Goq8JFpALAGzd3f17cgdkwc
6yfZ7IxRMfiPRjow0PTfwo7kGNwQLfR02sThbj/686qxdB+zyPcBUOUQtiqslijp
vjz00S3unnskd3Lso/0q4GPdGcI6jCftiteqMIicY3gp2CzZGhJEH9mvqrY6o7xu
Jg8YjKS3ARSsN14S+E4fbl6Qt57GXt9PBP9RrVEYxx7cVbQ8tSU62u7MNaNl3cjo
z5EJ9gr8+ADvqwME03EaNEGgQnz7yWJML8mg2KpYQzdjltJoDy9egC/CRiT4ni2l
P3cPo8Jq6+F85FCRfetD6xal328fZnXQ8BMW1Rs0Jp52FHc5NklBX+oGdubKgx4X
nbSV78hSeHqcMPmtR9H2wgKaKO3G1h8xDX3AzA78kENNrQfKVe9oxBNoahpCDRqN
Df2g6jCRM8tFhxfUJlBMyw0RmeaJOQtzRch8Oko27fvoUh7NMgWRb2ek6MjxLm6w
cikTF88Lus7gF3L2+1Flmg==
`protect END_PROTECTED
