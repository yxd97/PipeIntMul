`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+JaXScdLXqWK/bXsBWYGLe7TeYjEPBxTMnwBguqC7RGaqfwwK/eQbRGYZPSi+DHC
QSMhZ9jKMI0mzlugbLX3/0fiYNtz7VbMFQxUHDTT9Pgy3uX97ITkA4NA7g7BtAUt
CXyvpNvDs0rWz+4dOcaGZUvIu5XFr7tjLgYUMzjRJJWOXjVniMNw7dg3Epjk2pvF
ao4o1rGipENErznHd99OhbrA1xrJ+6mV7AGOm3A6L/4=
`protect END_PROTECTED
