`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5qY9BBDEkFTcwqdVkX/PCYoUYOJsXtxdqCQqAPO1f4zxP7AlKc61M434+PUxfjH
adL/KtaAKBAVOJw3NbOz5mUKPbcJsZPOJQW8y9dBAnyRrl4tAIFJmmDlp3LMLx7O
FB7qq3oSDN8b4BfafIY7aSueAZ7Zs0axre3KVf48BHHFtUeavaeiBr57QX/WYJKu
AAviJXfx7wiiQC+raLMaRXTf+BBjGW0OtefrOdJgOhbck2mDYljwOWfP7Eem0uin
R6ny4Y6yQiYRDhA6gUpk3NMUw0Nb87LZcu8hfPurb2koxw+PcxeUwchr6tQj4uGl
ysSZ8JkNyvNcNvDqVftt4y0PIQ7cFnGvK+is7u0CBUx4QEkzD0BgozxOLMPjCjdw
R04n9RZA3xE6jtLGfzbNwAQhmvjMds0T4hha2CLa7eS9Tin51NHNrKa4siW5X6Kf
0ndIzfU/RQTYwqqffPMZCgQ/85dq3cYB3uy2PF7dJp2jhU3DRh4JGSY/uVCryRa7
8MrHY54K8UY98hdhgX4NXBqSa0QMimX2UutjmMtXHH+cn3nkyBAYC6m6zFAbQUYN
AQf9O3NXAUIFFxu3AULgVskeax/KVNe18/+btHMzHZaDiRt7ludUVwhtLU5tPMN3
xS+u7D6UJAeGZINtmp2H4GmL0ItB+Ot7ZtBt2pR8nPgfnvRsTb70CkNLayk8zRur
ZMIQNJ9s1q9S2vls9OKIKN8FxbHTqsAylLI/r5eReWGaDTsXWciKIJ4/dmfk5HRX
AC23l/t6zd/ohzx64IW25R3ftnpHitiG50/3up6hx4IdjbI8hUPfcGzKUO5FNTxB
OgvKKcoI3dqag14a6FdBdHfbhi9PB6/VFvVzNKONgUXUnUDGMVFV4XyOTxMjpxd7
CHWC+8x9fwBW3CF0VlMVzvJfgkdpUJXr+XTOKOuxAoH0rdMc4hZsmE3Gl18UU2tT
DdKkeDK4NOKWPE2OGJJu20gG2XgJ5ACcPYH7dZgxPQrU07yJU2cd/Tun0ElgVhIP
wcMkReyWtWtqxPAYfpMGMeqHWDVj2sqUkI2dPxRm1/AEWsH9aXgLQqulFOzgMAt/
mLFj8GtghGBU8sYHqkjoODU2EXfgD8OKulRzIx6h6VMuBJ3YBI0Qs2/aZWZvTTUL
rAd+q/0Ev8VeMUYkXOrunFxkqZUtS4TQ8NGRqtxKZaGxsh/lPk4quLcRDVYREVH5
sBhUS1EHmjgYH1CCzgetaednIB4+gBQQ6qPMrwKR+FDTxKChI83Z0a1Ex/m6jLul
1PpXdWR3KLTsVKGGgXDnIgRes4B14xOc8CmFs85F7wLrLAc3cHshOo3ioXvY12B1
Eg1KguvSnuQec6wnp9aZig==
`protect END_PROTECTED
