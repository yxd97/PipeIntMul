`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R1YeBF+rxcGlK/bi1q3Wn+EdKyDVre6+im2aoLCUv0wyQLFsMk6UiXnT+ow1gDfx
hJ9sQ7NIc6tZxOIJ/dmXg6reQg0Tdcwr87q1z2L5dfKZsLOSXremSdFMBS0jx1B2
DMAbsU0Ed+dfCPFYPsn8F5o1s8wkmqT1ZroUXi13dMpPSenOOmlgjCya1ULWDqPk
TX0bcpB/mE/PWJj1A8mrcX6awlgrINvAOyCXU5OFr/ZonEQt3m17kcRfbFBd1lLX
gnSlWEpv6ttpt0qP164QLjcHyr1BmX6whdMqCP1RDrnNtcOR5e326wnliAO3BAjE
6zXIUXxrGh4nzcdZHzSgWBs7s02aNQZk7bgK+ryCQHE9xz1JTEmI77dQSvRLdBh1
3X0T+a0L/XZGyHqPWsQjj+1AW9lesADNXmtC3NCmVH903KLYXAfktbW5cTcWwrga
PX1T72Xph2DAIljW5N6Eo8Fm3Jlsiw7X1toE/c5uNVMsWShq8CpXNbb9vWlPlcla
2+NqqOgkyqmbyfPc9OFtNAUHBtPlgJ1aAeT8pun7JNI/ud4QUgABrqMb3cD+Lt6y
tYCCDRUnDrqbfdwk0SJfwA==
`protect END_PROTECTED
