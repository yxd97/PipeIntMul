`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xVvvYaLEbnVVqlnlPjx+rE63WYpZM2X91leYERxz5dQ4g/bI7G24CQkLRRRr52oR
R/GvhwlpfjmWFK47GEndAbB7gnMdlHMqOOUkBMXM0mDmreGSLCvF5Wg0qLNEEKTT
JHmfeSzTCLvi9HIhz2W85j4W4uDE7OCZIkHk/SvS1y2aQhLTw8B4MQobtrafSQHw
7Jh1oIr4GSdCnKD4YCqqirLx+zDGaGcXHyfnPD9pw+/qc87DaTBrr69jUj4dfXA/
jPIHuMlb/G0t571hH7lMXZsniZ4RijeD05lrb7STvfxqtWnq1HPM4YgKKMugM7Q8
+ydwdb7mLWgFPKLdoTlCAn/e2JYhVZSWFLUI7B04X4zS1cOSJytQpStVP0LeZXLX
iTkMiVwU8PBemagC1VppWhNo2NXcduPXKJ4HlGQIWNgJO8s56herDijmUOukNzoC
fx3Zukv3R1tbtJDQF8dGF7IdymlKspeCm3RgMcUuS0/KVSaYiA5OVsDVosPlVEWV
41Gpb/LjuHim91c6orRV7EIg920q6jWG8CbaRGDWPt5ygKinV4nc3G+9fP8/mX0W
VR0+DBsJz5aQ9twIy1xHvJFbNtlNfl4qcxQowNZgbXuYm6YZrYQbG+NDE1HQ6kAs
l8HtSTrXAgjB3Zm2i2kEs4UvtXI6skK3dOCiUR6RsCHreaAeCVbQjHSeQg7kePFR
R/eBFEOosAOb0A/pVfwfArgvvxPHQjIoplQ781oe+izf5wGG761yTIIIRX9Q1Qap
hpT7nEN3R+3MniJIoSZNUJxBwYhZ7i5WxvhbEhPCELdo5/MtcTGRzgGsDYDw7y5I
ahByyM/e2juVLv7RHAvZOJI1HxXuzQ1rez7JpkIw+hMZM7puXMxAh5afbGxIysYr
6jIJ7mAReYHn7Em1E5TL5yXtSMWLSDbAUTRdQBZ4y8A1llTGRwjG695d2ESfTThV
FGyTAO1tOZNoEgeyU/WLlPzsrGH0M3ugC0SSCUYFY7wk1fe15yTjVAKktIB2F8VQ
m7Hx0tOEW6SVdaey0NgipdtIdzLRn7Lr1/wOgjHYZms5BVZFMfSvf4tfX7SlqrfX
3JxjHJLhy+ISihlvbVJ8Q+bBYmx0MHFeT3p7hTR30UfiUo/8Z0dkN4+zLCm/iCSo
4xPBTkrq3+aECQgo2R4GTZMeGDjXg7zYLakAuDUGyZBLhSsWAn9GT+n4DEy/Ox3E
ztqEnarXZN3y1kRRBGSXzWY1SFqBd43fh6cW10y9tuNMWlPwosc1UlFlisoMOcQb
EqQDcwXD1rQEBm4XmgL31ib5xrTBh165V1TBrR4Xz//x7ykOa4PyQvi1jc1p8PQc
AE87845Tt3/Lp+6Gz2s/b31aR0cBfj3ahomNFkLUGmpKvancJ+qYXQ/GS6Ng+RG2
cVWuk7UE3J4h9KcHdakYmGPbSiMxQKhRjsBUxk95dLJfZGNazBBWBYYaLjr3T1gl
drZVW4+ETd3VPiUF9bEpD83PHVATL3mvnajYWzlTw8b33nRhOXSG3nriDJPP5drx
4/XFJ5fqx3+haZlql0tHVMYrHC+3awoMtBLcotRHzNBoMSk7Hzbz094TTT9Y/fhU
Hg31i3SgHiGUigq8HBgDpqPiaPYqit54Etcb15xqHWuFunEot9JIHIhU99nY0NTM
HFrm6QmXyucr4U8/Ic0GxDfmspDXGD8G96Xd8ZglBSaaEeVZCJqrjU6o37ghnDd4
pxhIBI/cB5tkjrs7qP0ukHvJ0+yUSqLLnCvlMmLwFrGgEw6YF8hITvosCH9TKGAX
9ns3c+MxzrqCiCCFDtzjLtehSSPtCY6wXPUYB203Zwgh93M1N/vU0NRBRCQmAIk6
STfcrTM0kC+uJHj5AEqVL+7Ql2v8sOYQ1uiqUHohQwlyKw70BzJtT/vLazTu1bJX
nPDEwMJD+92Z/TZ1mzQUVImRzlAqDHa5OJVerww5zmOTsQocbF5lmS2LMW2Wq6JB
rZsqxDwj1WOtp+aJbCUYoaTs4KAzM/Wc19i1Bucr3P8jMa1WBpyKLH9WfZtEL4Xw
/DjFwtXotNgQLMGcHuyfH76MltdjQHM+mcuCimkg5XGVRCT7ZMXfzTiLWo68XjdK
KN++293i8Tsi5YOPQnb2hyS4M1gzy0zkYXsL5xtJARXws/HrpXsR5kKqKcAy4p0f
NipOJ+FP4OGjbzp5J8zfxue+n79nBelp/eEC1RIfdXpjUQLleZMDBbmavhIB4cXw
UYWBWXtSUQnZ0GtpIF+/ri7nCGUXgYWshepoKhNWo5VhBSEHQbTcVb+uHXQ9ReOL
uIAyZ50zx+aL6FNvliUcv8lAzRxSvDtpCcz2yl5oz2qTYWerSc9Rz9sEc81vf3ja
tRruc7Afq36csRoRXc2rBGgZu3c4a6kF1hWGoC9uCmnKc31KXn403hir2LwoLvPQ
ehM/j0EB3DAi29cNlmGbU/Lu3O6CfcTCyIP99UH3ofkinD/Pt/ivgAZzyV7RCOu7
wRfFpzg1g6BgyIYJuaAFrC+LWOOm+6nBQnbnXF7XsUe3ObIS77drRkOoD8fqXgAU
xarbwlWdeTB8ea50NUF7DycCDZBBFaQ8SdX34OAUEvmukv8RWGwSmkVdvLV+mmGf
hRRhAKRbSAOzh68LVw/rsus19tiDIOTBAyJxTgeW25K9wmUzn0qBRNwQXY9UOzip
yASdfNXqCknAASb2ksstEcEgS2yH2P5ubokJwa9mZNjBaCz0BStG4ELjeWyLgtZx
MssVnB74jLQTvCy8/L0NN/Ezan4Q9mWn+t9Z1M+vvw1fjti9BXhIgQVWX0uMwhTb
NNJ/n/L6FwjdKJhkhysDO+mPCM+nu2aCD5lsep1aLOFlpTIHGj13lAAh5LsboU9s
cYM6FChX1DWZOuWTOb0OQw1y3IfTRvwc0WSZvvP1SzUj9IFoYUhBoiWy2MziNbUi
PykYu7QycfaCu/EQOgx8jXXMSFx4e0wfEZjVJqNMVstm1nCXUaFUHPSo70svEF9e
6xePR5gsmaaPZd40T2ffoMBSsuzoPcEeDs2h3LAU7VxYLQFdGIdAGklhZad17aUt
FQyAM/8aUn3R5u+RACv4nKNZwgHk0jfXu92Z+z/yGsCnWuHocRzGjSWEYpwrOaR4
u8TjxEFqCXb57DcGHoaZTJEOnXGvaSeZb71ACD4qoVJy7WvB7X351jYX8UKooH0n
/6AeSJlhoXxhHazYITllZGyvT+Onx7ChHi8rRTpiTQpfd3I+XVdY8j5cvt1EGo0c
sdZRaw2qRMJDDTyLUm1rhdLJVCeWvyqyy3WopKTs0mVwqJwb2LfyFRya7GSDF6lb
XJHFhnQfpMf06tnyCtL9/tyAmmFoXuqGjHSG+ne+h8FKGoHayFQHVD4ZiXW977pu
cIFYuzUJ36zSkN9sw0qOQ4zw855aeuRcZQpE3Jf+miIGFHMT3HAigJEjzIKS93YW
y1y5Jk50WoLaaFIr91Gtx9qZYhh0E70pTR5x12/BWppmVRYEJa6+1wOw1jmXvdYA
NcLTFY7iq7cDLfnfLQBnsuodrn+XqGNc7g38sav8PZtPCdBYzDmHoJACHwnXXWik
kbisA+NJQw/aMKm4El3Pi1KHa4Rph1/cTPyTfHOtDl/L69cs51Vgn1GeIP1bDuOX
6fShh4dtFOudGIr9wsTS9DsD4rBNNoMXdEjDCJf1tfdr1yoOgbR2HIwdaQQJwo0U
EFO+9C+qjz/Zt+j+EqJsgzeAipe/Gqpn/ul0SWCuDQHMpCmcDU6+tY0aZ3aANm3Y
8P2awGngeTEbeSLgfCdYXkOa/6dxmLROwzr2YrEakSH3gZH+jA54Uv1+zaTZ5PbL
KE7mKMttlvLlAh3gjX9b7bkoHSRa8o8yVRuAXS4ornkNKXZ1Fsraplq1RBvXIqJP
F35Sh2mUviQj5LaYErFlVqjF0pJjeML6cX07C1O6aMjtA7hbainOA9MYAqj26fJQ
6cNoUrSPZM4bbVtmkHjvrx+oLLCQkCt26Tyc+xxkvHG+8uChtD46GZJ7266dc9Qe
zPMBO3XbQWfhb2fZcA5dFKwRwNIZJjI6gyKtL03wgtM/Y+m7D9Em0oEuRuIexwNJ
+QMSu6owSpIezDEvG8U5IM/0Vsu1+QEeJ1t4T3OY1y77DE8MCbqEQoyhNZL0J00x
fqbwoob4J5PIBpQiIYkIB22l+E+BIwU6Fk7WDlDfWQ4M91De4VzwYNzhZPN3vYgh
eww5043Pyxz6H3fkm5vQgaWfDDaUM+bYLrQu+qos1vuT9EgmdnumkwJoFLU8cCER
jTHGVVqaysog1wAwPWKHXObY5bwOuxtXepKb9kG5ivWGhvlBZ4JXufjBZOPIJaqm
KWnduERkQKEsWcjefU22xP+b0i2lgBKTHrA/lcixk95ZZDC82U46ORetyBpvPG3j
uUfznULb9kBBdFPEitGUrNziWT+2+O7/HvU5SLuD7pipIHlk7cJQ7NxmWqPmAIh2
2ys7wv7CzQGIKATIqI1OOl05GLCZmXSYUS64CmF3uxn8U8Z8l+kR77M9oD1VZ/Oo
PPg5NEdvLXzNy+Gm4GKPxcXy+ZZhJ7JbXnYS0SW9fZyHuyEY2yC9DE7o3NtabyMo
9hYRr3exShhstA9/xEMGZGJkcmhJUKy62ApXHVOrogDLsF9VAClSCJHtFbPer4rn
dabfHRk1oT0uOWvtFTZYCUWDDpdL8RT405FOpUB2h1skNLm0zK+8Lei9B0VrS80d
j9JqBAGYsdliqyrEt3aT3gUSEMO7h1x43LejLm1QeGKFLAKZDpTrLKSVYAHDZkS/
aZjm+Az+xrdIHrxPBUQxS7byDH4plS9wlVqU65fefomMfbmvT5PcXPbOYqZxcy7e
ZN150bnEqlYReP9Dm/TbonKRpLJURWvo6g9mcV8z9uH/4H/dHBytwaHaNvYHKO1Q
XGpHZZd0XSuVtq1drplzJPlLgau6BrpLuEGD1zmvGE/8hVJmpt2YwGnzcAv33K8T
Mbgv9a9ptekyAZPCUkrstzYNofcwEhWof9mlPQj3itBmFLXVYbrxH3EhfiF5RG8x
JzEd7Gwa+WT814+p9TuahHqYkpPuceDWYuByl6VkJNdMuf3+egaofCsbpkYaQRt/
c8pPUdG/tDq9FQIID/Wu9mtoJc90xeoZ93bTpXb0Okr5KSE47x4jzE/HrJA8S0Jf
nyPR8VEJVmZR83aSZz0UXFhRGMvtXPkowkmdIuM9AtYtMiDcne8NFI0PcjVWkbMu
CMFwoydRgClCus8MO+5FrJJJg0wZwfeSSim0vELRKZsOgyBbw3kCgqxTQojIR8Eu
zLE5XkPsyHA0HnxT9I2r9i3DOBj0vliglERohuIYXbrSxZKbITtNK9iayu1QeFkU
h5lUaw6iV55ETnyV7B+5ZJfQ7H2fdBYKze9ZvhPLll4rU3IgxJ0KgScA4ELo4SnT
2SiElQbq3xzTHP+0Wj/+Ebrq0CTimEKzn1S7kXYDKYvBIwNXptHUJonpAEyLdkP4
iYjYiBCSH5TwjSarneKV9KwDVB1yAr+6QedewKIZqqRtcvWus0wXVKkJlSebV2Iv
a/NPA+Fxr7b7xsyA76yqtA4E0+zhoxwlWkiuvDZISIJdDOyAREUsjzSsntg6N1Lt
SHjVuJ6SuM+Xpld8z5haFzHr6MDa2RTL43M6oIH+Lhrg4+nHBI6kuUkYmcvas9I1
TCBdjUOaFI09AjftPuZUeYmV9ObrBRSIsLy4OXpO75RHFK3jWvhpMhG0U/j0X4FC
mkmVN1Sx3VvA8TyeTOF1WZjYwaP0GeHwRfivV6LYqd2V4NoPo1uJ1JOstVnt3Mn+
Cra1+N03cr405HvgsjrgrKPSF1JAG0yecOZpNEkYhfHONKtBOP6Y5XNTCXOhgKx7
oH0TEwiz3e5dyItmJfLeG4KUlUDdyaggrCT4lMjuYgKUivzxCd/odRdQF7kNU1ww
BqRTCFxJghTgQhsxSJ0eSZShq1Sg+VqGN1RvbXim/yDgmz+kk8W50JmVTIdsddtD
Amie264WWJ3ph+Jlx6/Iyi3lzkmMPmYcix1sUvQzRrD8nkdx28QrwYpbCE/nSVUB
gnpLh1zhT/YLSQkRUJNLjAT3yDK+fMsLbXBHjfXbvAdGdCqvixkNSlMmG1a8aG9R
rt9EE7BTuge1q89gn9BzQXjcQomVyrYS90/1zR7V9vEKzbeSV/MSkDZy9NPOl2Op
5fC9EmgCvNtsmmqQMpDTO0WXrtb1mZ6bXNFktlposZ/pNFTjLNBYx/raR2ZOytNZ
f59wHkDa00T9JBxz+JoGFVc/3pCs68fs0eIjUNKj4mFO24osCmQUCtDyBzw1VBhk
AkKTfKrmm2CUMYnK1wvHlmAhbAevJoAlSKtwRRUKlsk65KbKJ4V4Qh1/Suda+dz/
Kzogor1vZ0DzArKlyKMozTk7DTKqzd93+K5fjsa9saJgcNxh7ttnb6/clI25mxw/
fzERapbSup3svRy0q0hPYZt023zjMHGdyk0+nNkMkwmLLXC01n4BSeFArLEqjbfM
7bRDvmrziyvnSOLWN5BBPcljSNZDiRn/gIFnuA8DD+nYn521EYI4ettpJKTh5irk
X2qWJGVHfcVez7jWfhUOwpePx8xlEfw9kdSkc1/JUiqfYXiiKwcT6VbV877RgJB7
Dps94zhM0pcoIzE6IWrFCc8gcKNFfRUHPztkuVfeuPkwfxXsvoG9keyATcYaMwsy
1IIApaOA6BqQahz87z+Zpn6IA2RrvPwfYe4FWpGPvrsccT2mlzIsxzVmNnHIk4ct
kad0zAYckfk6+fs1n1gH3HcU/LtB2HJlWVeOREieXuFM+Fr9uCxQ/NUv37GKELhM
bvpfhSEP46hBleAudZIfKReAPNBGXF/3tJGE4TzsNGJDD9Yr0QOQeD4u4SUoF3uk
nEjqITA+0zNkHF5tWoUmVxVatEzy8rQDHYFqxrFX5fiydGUaRDAqfe7SK4E4fwP+
n9oemL9m3yXN69lHLSYP9xN9DMjPWArUM9a90jheBugrhLtsKWx8+APMVw5O/H3i
GNqJooG6fqGheZMkNh+QGwibE83rBeiRYGF8ot/3Of45A6sDZbwe3MIHu/oABj8A
vxgw2qKJnCrWT4RH6ykYyAJNWDfqJEeZK6c6P8Aib7/5YkBVT6eKndAqLRJi1Bur
U8+Vzl7VbWAVwaAB3SHBS4psAQXJ0zp7Hl3kAWmkSDY1q/TrQVdnFPred3jgV+st
hFZiYVDB+/CNq4qIQHebaAG8QO5H5uHFIjfJdGxkT0Vp+EcwX9tcKaKFIWtPl/l+
6xZyE1ZQsLFvMPIHsZTTOFJyvXw57cdGGS7bMn5ZxHUhtNO+eY9qIUsHC4cN89yc
DBANruYTrixljSVx42HE2dvr6BEtPK50xsarpe/nJSNqC77+vMcqtCmZLYeh4r+D
qbQ8fMCbi9ZVpoaU9M8evuNyhGMgZa8qvH1Kw2YnwiJ3q5e0ZShXq7sTmOUKD4/B
8LVDeQF0hPjz1NNXI3Y3C33u4S6kEwJFDivim5gWs66qtRIAoT5yLYnXVK9HBzEE
CIZv93/SQ4I4UN3JLzh50RqKYH7rt9I6STnNxKBsgRpu9jXI6c7oxNoOOCwnQR+3
XsXoJg1TthK3Xa5QvLZV4nIKdIC/QOOCJjdALE1cJVNBA37VkwH0z7S+yEJrzbK2
VgS5CJ6FHhFmSMQFEZY/1kvFLfVJgYw828k5u3CXceIMtEXAM6W1mWBdCvlvjklA
JJmg7AymbaDVIdq1lMtsuxG79871g9ZBqeJ8f6kwODP39hXpUXd92IuLELKQRu9U
VXBzBU5PxhU7mzf28YlelDRHHfleCoHhoxl1ayJ5KF6NpyTbhU0I4s8lzTmBPYtk
arNgyuGjp/7mswtnrD/3dFvoICNjsWRtsZh/RxHMxSsWkvJo93F9bSuIDe7Fqswx
RPk3Nejl+ews/moGaZv6XkXWLhlVq2L6uUtY+tnRS8h0cWx/YVXW/V10/B9NwmSB
EOYdPv7UTR54tzN0WjCKE3E21zJfgoELBygOeH8PR3/wVfIcRWpBYo2rADZ2XHHo
19mwulHgRDfXiOLBnTUUmjv1kLqOiLlushcnTkplAsgj9tQVbYRA09riCfzAzrDP
xXKoZLlw4nvbCiieF/Ye4NEQBtLLDK9hjekeeVFiqskrLidOyRhDTotzZ1Kteiba
gBnB9JdLU7fC1uaDJVjsc4RrPK66NnxxPl4mJR6veCi1C1JRCZ4CACTJJqAGTTlZ
XLOxIdkKCe6gR8C12c+gOW25jRyqBehHeFJarPBj17Eu8Kgh1VOuIA3wkvw4qtvh
x/pBp7gypCI8DZHnqLel3U93+ewO0Z7qL4c7mr6QgGyqTQdw1rb8D6otrN7ECOhM
DQCXLz2LW/l11zs63/gEWS4yPQ/WS2PGsYCY7ogXNKU4rqQG1IkjhEe5nzP5pWGd
N4V34ac+9b7WyC8XwXor8QwplTvUXXsncgukzj0Ki6A8HC193DCPAZryKAbdzOkN
NAAtpKgj7i0CMSbKOqOFgY3oPVv9ah8oydZVD/KYoMNxuc1Fwn1A/x9sQ6vS98dZ
hJs1A1LIxDkMvXoLyM+nAbN00PxBE5aM/Om0ggQGFbHwxh6udYRnTMEr4P4L0Ywl
5reW8RmYGvBjVU0iW8axk8iew6XLbMrvsz+FP8NPB9nQDmnCEG4wq4Gd8V6NKbFR
YDxB3Oecniyx4OVILglI8f69ZLJEMh1FtTkV1wC36cWC+uGMyMecxb/K+O9Ss4ey
Omfi8rP6rqGJ1oFwVj350nbAg+BYlmqgaB1h5RZ/n/wPrVB6H/k9Nkor7zFmw+BP
wLiRvo3mEjS+I5/IBQdoUlLKSWMcO+tUQljy5/03P2az1y4mb5RQFG0rGcRSfnCy
XnIXXlRCn41wfOGcDmvad3sB6B8YpS6BD9sQ8TPilB508+G3znaskWhJB41ZhRtW
WsyMxrBbM9p4y5RLIcVFIj/9ZrFBV6quUE4MsgCKZVtxBLCTdvMeEyCQNCkrbjDW
e6X5+IV+0F+9VY75otlwCjYbw4GrfxwpS6ugJ3eOdFtfFMcHwvYA3m8onU+yFgCp
CwwIMVLmVrAQ829RDxVRQ66V3DezYGwX1Ou5pAimGXWNxZqimt5jETspCDpGDOgd
AdYOeq/KFVmMt43nY1ljuxeT9l0Uj7ZqoSIFmlvwDV5Bavy/gyVp+H96dOzKWSB1
sln1x8zt1f/lIPevMsPSlzJkcaiNvYeIyAYgtWd9qEd4PceMOt1UBpdZm9YfMSLc
NoYG1mTL87mV5EEb9Y0FoNMWg0oQ4gV6ryTyX9zwqDcu2ihJW2OkiW+WHdqiNgQe
cjf3mbiO5uD2yLCJIJ+YuK/LvKh7jstV30iusyp+NyBYrWAuxQVUfE4cxiAOILXl
iqabaR3Nmwh7OWd1LVavIi0t+9zZRvBr4rfDvKZ9gV2+1iBnagENKRigEPK4sP/Q
BjprcL+QggCdB8qecDjpLEKYDOUnEBakW6OvgMvew04TTc3+GvoV36kk1nxSw4ny
1TfJyQu3+e/CmPBluRK5JJG54KPOqnA8LKXI8CWz3TRRJaSPnW+lIwhwjbcdXOiO
R420CcWHHrHWfFlE8lyTEMn+vPMryS5NHStKwu4Aw9U7p9XF82Pm5kZ8yZKQ/y/k
iHrn9LbVAUsjmVZ+G6JcgObwOI5pBTCQqhMKHoO+OLlrEJVwOpt0+g0CPh2p0rjR
aF0bl9Tqngo7VG3RyB5erDdE6nm9Vmpgmu1lC2hiCDqAnR3NJ/53a1F07av+QfOs
S6nB9kt3RA8zOqjinC7ioz6WiVC0FO7kPDd7Vi2MjoaaAJXwhMomDnBw12g8t/37
6cHF4K7xXgCAbRnrJS/+D3yECs69VbRrXnuoXwvfcaX1M9bsE4Zsz0krCzkKGLtr
q7YkhupYP3hQ252eDQlD/KkJmCi4MALb2Pk49PUVNNwtfYcwbvoVwFcGaTyQOy8x
lTtlrJsTLiE2xyytZN0mzF4MGNqxsVasvoTyQjFbor+Q/G0q3w0D/l9LIxOYKc4n
epqqAxUB14WkrHQdeSd4EEp2IobvDe7Wr5z8izuR0FVr7rcJKnckynGRtE6JPxAP
vbNFowRQCKJBNNfsaQTjTmpnv7yZVhOLKm20N/eJdalOp2vfju/sh+9U8cGjnxlO
tLeCbJiJCid8akSj+YDAyTAtB1PNR60NwR7TpzaOGDHCmdASeSbWFqNrYcAsVhta
WY4Re+GD67WGqOezG96JMZKp9VTU7eRm9ZMp2/FNxXEKgoM0d3WK6DFhHJousnS5
+kg1GhBg6gh2rXEitRLaNsEWGMmMMbefss2i4IfH26pwCWGlY74EdGoqLKA8ZARd
ZpCXNq0tO4CEfci6LAqbrL/TedNdH5xXS61qga0DT841MgYl8tcW4cz9BlXyuPL1
97KbwGD4JZKXad044qmM3aeiivvGsoMy2w2bcNL0WU8sJEL771K3ZbFiN+l1RBrK
fkAlDCZhhXnI3ESAHJA+FOYBv6XJqP+LYkYxkrsZPVoOw/WCV3mLM0kAOM1MrEWz
VOdMBS+w9N5t4Hg7CpzYTcv6pSmifuZQ57vDQJA/qpmjorQ766J+SzhLPRGTw5Dh
zqIuBFTX25B3j6oU4bWQDTK7Ay3CaUg8wZA4Pd69deQ5h8ptoGYHhqY+qVZmM+w1
1nBrSR7wD6MrxgdNFNaS4iYHk8pusraadQNy3Ks3ztS3LKDMT/taUXDHq8vaj0VH
EubnyWr9fFw2TXy+voH6S/GqyHhY+v1TY6LrJR1UiU3XbnyG0miy6FUCAvV9KOws
13su1t8B58Et967z7TNkrwChsZOQEDZa0233quzX/x/U09uahX9VpIIrekGlwQkJ
katjrlvO2WmIfSH1hU+doqKcLqqLv0cgO7WVnqA99LUShmL4HlcLc/qVx4r4FQrM
f7Tzi3sTByqBsDBdiriwgw0nodU+DF42CmSES+jCBEyTT1CgUqPAXBiJ19acmIDR
ZvLTzS/oyKcIFDM2v9jsRD5SoE5vNc0ZK40SWmqBLHNtuRLHNuz/oHatzFFlCq1l
H7j17i0f8mzeHlxZvuCd7fEY9+yvcrxS6S7JXUpZA/ESgglACT+fClvFXHS0zZmx
UDj6zLDRha5z11FYkhIQKFRYzIc2AOhLmjPq7aBHfn6U5A+85j2MFeVvnesr7CLu
T79dsd00jHDAsRy6AvESyFcnhlutuKYJYT9+txpHGt07ocj8x0fUBJgWapQuIo9t
EQaLlPsiZHwsdaUOeY+kB9nmmmz73pWErzilfpSd4bQcs0JWgOxW9UTNpKcYB9tg
yRtiKIJ1nWXy5YXwsg99Ueg31tg004djpMTekUlqO7hBxXxnbW6QvJ5ue1wiO2qO
KOIRc2HhggWSuJgkrs5BJRrmkiwqOeN124DF09SKaYo6VfkRfXZnl4CBEJ49hwr3
BByoLK7RiaR7yOlhnSMzqOZC/u7IiScIfqrdz6TTUev2N0y/isg1zIdXPKPuA25B
OwG/2Q4tJ1s6cy7NQET/xT88REZW+Nq8EYcu9yoKeg8iwC43tg+G/aFrK/wCWDvs
JL0pw1Td86sbPNVFsmkM7OlzRVJAE4G3ln8l5x2C5KtZDLTgnp3wWTpkTPPyLWIL
mNgapZ4HqrG9AlpsrqmO1SwxTQCmvFhhLtSyP1nBy7oLOcZ9V+e2rRy0htT6I6iP
oj2wbRgUerQt2WrrS+3TfR1jG5HejdtRyjflkG/hUg8Ch5sAntGsKApuN5TdLosh
Hc6ceq7i9D/czgkAIzDrPStJqvdl7SR30rjbeTcE/HHsAVdsi5nD+uDmNMKU9eFJ
k7PkN8VM4rx3e1LSIdXfJTCi3dxfcl7i1h3XID8os+iHN4JcAPkz3UOJ4uwSgdJi
nwAzgDXF1DHr1gk7Bb9ni+CkgFTJ/blFY6SrCAE2aQnvBAe5t3354AVSq33C0usW
5xBoqcO+Dg0E/+hrXGaQd5GdZni811yp3n4cbyWTxQuZQE114qg+pen9eTcTISUi
Mjo3sTyblPnO+47P/h+JVuLuU+FLrd8eTVq6l5m3RN7lhwDEMviaBHM0sDy9uJm8
29Nygy6aBQzi53C/D0uQzErwuOUq39FjKG19jiULJsyosAUlU1PyDwYZX9dWvD0K
FLrz05v+gOusKPcNYG8lo1CjKW9rWnJQ17Vu7nof+qplaO9CC4OyxJcsOB+H62y/
vPL1gB37ZgIjcyRJWjyx38zsgfnBm6m3pVLU9gRNCYyGqY/y1TP1oKyD/3P7lzLJ
Q204zu0S2zPn9GC56uvNQXl5maVAk5Akj3EOzD9Laqoaz5F/bVxfuSjv9XxCGYDt
eHxMXpR5WF7BSVvIlr9n6tTMTTKZH1h76MhK6Yd+cY1Vg2qe7teJPNQONotvFFHa
A4Y+a2LhaeFNzTNa7IMufHAPifaY5XBbfec/oXpkeI4LCUzEJKPdew5S0Gy6jGJ5
Ue0QWg4Y0OONepoxH9K69pHt4rMMp6u5BkDIMlx3fsfPrZkM2FnDXZRnrkT6nS+u
UYK2GlRkkXJiqChnBblpflVlz5CoIihPDrpKEYKYfhRZaCtYbZV0cFVP0KZkHshK
fDLPTGmZAdVTF8kBi34tRXY2rUFE1Lr7o6E38oCgWgoFLIdmwOY/OdvIOmpwtS1+
6JbREIQj1NgKGILj+u54D3BRC7ZSsDsyZAuIzrIQfwMPqzF/LPm+DlQ6GiZet/3H
y8pBlgvnYPWp+FQYUlTBFDMHT2hWj2nTjM74/73d8XPvrRHCJRCemmcIFbIMyt8x
7RUZr6TyKCkangcaC576Sv6jws1msX+/FmFWdCicz6JpoNYRvcoWk9OJvKIPFWp8
J9dXOAOrtTFBl9igBMxlA071QTqE4SI22pKR7qDJdxiwI5szlhwwTG6x4CgKGK3B
0ELHhbBKHhiaLVpB3HTmPA5a6hxYmM33h4HDQBVMSJKDxBLSQtNyHo1MGxBjka7A
33AhXgXuCcM0He+fu6KBBRoJbba1JwGacuLYkGcb+gOPF9Ol/1xX8LU0pOtTBIQL
zMv9qm2XEBvwqnU0ODaP+XHEGmb/mX9fn+GuqjF/PLDQPalyJFHSl97/D6U5pVE5
AyE2zuyfoefjE4Tm5GgM+fVBg+nPXmp7nfR8FRXbPL2DbLi8qOr3Bt1rjtajIz5v
2FvHnzroZTaLX7JUfD4XmqUiO5bjFQiHjQHbgN+YmO7oyWWnmOOZFUpebThto9DM
JJb8o0/tYfzeZn6MXoav6BwON5/y1JhcaN5OTTRp7XGlIcdhYzT8E91q4VBIES/3
KglpG1OEm8aSJxTep4+2ISb5LCrtm6gLlQ+jF7l6udajDMxSnnj2epMFVCr4ay6U
I063JzPGZ1USwYi25xJZsc8SRd34XWS0Ur1E1+WeWQb2QMLDioFCUfm4gofm4KZ5
EIRf3h1NqRCVjxWIxjiBD81Lu1oLJjW1Kiy7LDonNJEHYt4IsppnOnUPTQDTFUFW
VGbbq8WUk479mbDaaJSiCr5dcS7mRrqRESaj36Ka/+cqUjWwSWSObVIic3DtB2od
Rk1nYpqY6n+ZATNlkNy+e3SJWsleAl7DZ9xFroH0fOJiNJ6prG+cIDodze/UOcmq
Trq3pF0ZgrihJUk65vvtwIGeVBoGOVlEn8DYfrLdMReVGWh5ClRFIau4QkX9ps+E
JuwbiI7A+XgAX9eARZsGw0K1e+PryDBhdH6/ABuVSeYypVs/KRQY4RRTCY1cJbxP
n2hCxhSeDYgo/W8EfdiFaJFTGxZ5MIpQA13kVBtMq9g65vDw6RgIWi4uvsJOInHh
Q11FuUV6fqFXdn1lhRtKpkbyTsxrrT7Nn0t2vK/SYfEXynQVqdokF91xNivDzEdT
1tvTH95/e6I6UsLqg+ggZgeBLIwezLvPqWzK7bh+6u3Cw4CX7n6Li6uSc8OskrQM
rfaO/CdVsqA0lxiEMig9tEwbDrXqJENsflYeDIZXusD421BTQf8s8CAsd192fvEm
8jElzdGKkUiIk3q7fCQlhmoUgD4R2vuCJvHGKnEck2w=
`protect END_PROTECTED
