`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3YLBT1QbJ5WxMtpYw9DAd0B74H+t0RWZvbDaiA7KDfkWGZWaDaeGieFMc0q9mRXf
v6b5Tv516iL7X7Aj97luNCt/vf1CDfOP5ze17Q6bxmoMXgsINg1lA9oYDPqIUovq
4wz73DR1l958/lV/Acg59RJiTnAgxLOz/ljCNeakmCzd7PSPNTdpnVymuemyhZRw
84a0wNQ1wYQ0g5oaGnmg4PK3aOJoXfEcR2cl6+vr8yV5LLBUyRgzhodk8CXdn4y8
xSKzTTz4wf5Ie6VampOQ+dqZfV937GBvXIEqPFo78g2Xnt6zhygOwDc7HVUw0fv+
`protect END_PROTECTED
