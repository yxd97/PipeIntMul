`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UqHNhv4ujg3eOpporJ7HijXN+F8vjoDYOLXAJF2HUycY1tNDBKuKOzNZi+iKvGn
0ehGQ0b2vZvyOuxK9H+gxWYUbzcHMNtULqDFsfTjaYmJGuzZ6oFTBOHAVFg+/Xjq
ie02ALmSXTg/vpfXDej+YsN9B5v2xAlWU9KaarxBndJoIXEJxOxTTB4XOgzGrGJC
HFgEhGSmaCw2bp2d5ZMLR5xfAw6Xt9NE4WzLfG8bF9Nq/23dUKnFKvUlrSDfkqn5
DlN4Ew+Edf47phv3CgtB92Wp6scJ+BM2tpdTMdtAFhJ0wVqk9ayusK/SeLR6ITQ+
B3dY/hdL82J+8LPgVNJe8vBU8Hn7nbuUpaLeE6Q8u3SjJOfJPWehdMn9fz9aFwt3
74JASunktVdtZoJ3Bwj2Wy4HfH5WAx/WP8GW+I81W3qdX20BhdpDtdIZyY1QiEGg
D6c0EPj1XUGcLORk3L88xZPN1sX5adP/6diQK+M0zYVT0puYsSKrH+eJI0xXipnW
FOlbL0IwdP/IV3YF6iODTRo1CZrF7OxGbSBR3A8VSBg=
`protect END_PROTECTED
