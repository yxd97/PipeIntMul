`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rUJTmMXYWE6hwphrTxLbevLAAvdyO9tTE4ku8mg2ENCkt8IbeAXnqSJgJ+GZe32
HP8K0lM9xinyrcqKKUBnkugEmvQCLJcnszId83488JD7pF/7KLyY3cfgiRjVleXB
EgVbVlxnNqIHj9EkKdvSA7xlI33ujY06MNqqMzs5UpI9ySaoLekII+FjbYBniFR0
7OGHJuBwOH6ovsQaIwSPCog71BqyjbrunF2md0MK35EZbYOzovUNn9bcZNZfqfuR
JN6qdmtcMHq8exfQAjpuusS0Ej68r2WpxlrByPfu2dQ7jyWJ+85WLBOAqVaCB/A2
e8podoE9XB9SOUpOqI5EoSR6QZTcJQ1Ex/2UvB9V7yvQH+4VPBXERVsY6CRttLyP
gDfX8ocBjsdcpVEJj2l7Mw4FXbz+REb5Jj0lS/GKudJOolgMiHXYYUUg1QaUIvTp
z80tkbvti/F7GaG+O7rydITgO04eST0MU5ju31GPTctDWAIGvAIPtPrX9OIBcUqr
iX8LwOw6cgk/ROo+WLjgYZWuVCjgM/ycv9MrWEEPEzCp7sDJVumr9ETu4P1DjpXs
unncHnD9KhA1Awm2xodo7eawGC6pwncNy859vh512dWADgJwrnDnfY8FRGlEhN1d
0ASKXR3InAL6dihxOfd8tsWERCnzhZGd08WskI+d2ALZXcunBPaw7aWbT6JfFxPT
huDBg3bakaaIFr5kZPgTIEM7BS0RVlJwGVdZ+DLMDZmVe+HJPxhyECPYAVgG/iBD
SUdXwbF+qBjRhwU9rKTw380oDhmls2485u4lIDAN2pi+oES0MFrhLOJYrLFi/av8
QkFbn0V8lLnPUcQfppRx8a3ZPd/sLJOmulqK1UfscTRkPqS8HSe62rc9EAku01dF
iwlNgHAGZOsTQvKNLYTzLjELK1nc10MvrSbr46yO4Iv3haZtlTEZO+EBVOBNqXqD
RulknCb1ljN09UpAmGYqJapFZEoK1GLDPYLeiaDf6vCcQy3EmSDpQHPezsrrFvNt
4OhLSN5DHi4GieUyTVmo6SXaZYzPX1CjmSaqlzFxw4JD2Xwt+LuXPPfXYPPPIiVN
yXKqL5Rc8Q/VaVTkpXBFKDW+dKn8nAF2WQ3Ye8CSEnYqTgM95t40qFZBic80Xf09
x7Mh3/O2v7lUaoP9rcrVP6ltFjzJ7NrdxcQl6ytoFCGeLVN/O+vjJS3axS9ZW2pC
`protect END_PROTECTED
