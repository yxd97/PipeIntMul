`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eKDk5XhP8jYWfi2oT7jkZcZEQu3F1mt/YaJ6XWqEYG0MDgU+NtfRF3/E1US6NLlu
zNyZhgKeUPSjHXBlomsXkJVO+PGeyeLSoOhp2+ylkMPh1df0VM0+m5YeJyj0c1do
Ie4ys1gkq5AkGEZwD/ppJL42wipdaj7Kvu6iSmOHIQf5wG+8KSgze/M9eyUsuj19
KJuH8vPsbl7oi/jnHfxGD1pAmY/Lsc1ud+OcOZRF1603noEWGnidal+en8S/0Fph
tKUj9LJhPI7RanlM1ZjNc5egX8t++KOoRAc6ytqSCkK8c8w/FZqOCUcCNNdaCwJf
K9qYl6+tmBEyntvvUkshqW9JY/I+0jkEYRGBLIkssCpD8D28E8AlQe8KXWb86Fsd
+/bp3bB6uU8Hu2ShblgXMWUnqpoWDpl4YZEu+KUeLpkoNHqsp1wcZmc1I/Ndm6Sq
wKu47lGb/E+TVKkkdMyux44BMif9esTGKGr34qZxdeEXgRkw+fQtyMBYBjoavHYq
+Npwnl/Lbzrvmwa4GOeF+fRh2n1UJK99CYW+nxUYb8uqmzQdzLbfdG4SS+6b+RUK
1BU41ZDiqEI3AhUxsJyWBmc9lKtSZa7CJ5vFkaATb571gNFC32NDZgKhsSLhTP/E
Oukvh7SUmRna6KmeqSAWHh3PzOITB+LbVwagBhYEYUY=
`protect END_PROTECTED
