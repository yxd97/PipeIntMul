`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQnjjqlSKZcZy/OEvdAm9x+DReO03kfRmWff/OWXjE9fTypr1bkFSBQdDWf5Jseo
bK2i5GxPk+qn2kd/SiV0Hv8+0hML/YeBFv8hdt/i1kBGjf0IKj8KvobsYd6NTUUp
v9BJfyIzZDrCdNjmAwbslacNF2R4eQYsMVqCZBQ+mLG0rq+BdbufdYikc4/4te5T
6tom4F21O6be2Y07F+xbvi+OQBK9jS/DhLvSLOWbnri5JXef9Cw+q4LYpzcvLuta
EBHtOyauC+MxvpuSJuqmSdCZAOIqcpCy1FY5a3ACYAVLaWe/X+KihhqSKm3W485w
H03jkV5mnetFgDEo/nNNRKwtNtu5rLe3H1Jecz/6phAehEzA6eHJSWUf/TOheGx2
xjScQo/ddOm3+TgvGHNina7OgJklo3Zo9Z3dBsQ3vGds4brv+BLIAqxLHgIBblzz
V594RDTJaZAk1XMJlzN0AxAhXlrja69fF9K/mViN7VEq7R8uaKfkKIlmlDerjsD+
VeUmNlJXnFRVDUCPmA9FaP3PbIkQ8IsL7XSdy/ZVxGr4AVYgW8Z7v7Um4J/kdvaZ
IkZ0+g1/7IfRcoboGx4cyAnKLSpe8wzVOotXIifQPJzWT4c248UJJNqeChHv4u7N
4Z58NnL6HT4tKOS6rWoteBt407gS3OZpsrjO6oxJLRP8Djj/mvIS6Kg2ETTsVSen
+orCAmIFfu/JWQmYzgQNmEVdGARbf0x/3njIhszj1yo=
`protect END_PROTECTED
