`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FC9ZByNQyfa8cwD0Fg1JMR1DVfvuJDUNFeQU7Qg3JJ4BprDWDtHgJsJb1212BNR
iluushGbcZxrGvtgpIPYyBWRjuTiYqZLu8JYjMKQLKrzzJX8YfmEDr1Wgig3jGLt
l6ym6AvrkxIiI3u5q0RNAtUngaJQy3xUgRt37PQhGZ48ItuHnhOHkKiQUC1E4ZxL
Ti6ujoZDOsNqLWIINJWwVWUC/WcQ/KtGGrjCQf37bELAoq0xWexFpJR6d4ji/DyU
bArhpPtUCujHi6R1JNzdg1iqFc6WPkpe9ZNODAY1Or4rwtp7WFXnchWiLI8QAXRo
M96FJn9ojoGBqogOe1pzK268GjpjjWLFjgJrZOvFeMOpm4eaUYcw8fdsAHtSSZpu
+sZmvRQVekmB3n38MozGkP2up8SHq9G2iqPrz1SQkckUJLg+ZpQBThfzFr8JK+b4
7rvH7mmlekLIHZgsPlT+UO716tCdZtJsYjRbXSNkKsELgdWAngBl99wsU7uwvhmS
1Kuuptg+hB7s3sh0rvPRDiT2kGWAcqL6HZVsYkpV+L1SiDKrNfEtz7x/doSphvi3
7sZvjxlwe4dG0i0/b76x+QTTEvz6+TUboPD3nnWkMyO6vf/YOX17Qs9mKUOcAO7j
kIXWhAQ7SUnXEuoWLvlfa9hWuSHLzDLdwT+IsQcQ8QLmP5lJLYeHu7Yn6jWmIDJu
yqrG2Zy5iGbBHsvdWHQv6YlA0VGM3qQ2MdUZrCEifj+Yp2b+o03w0OvZjB+XMFcx
8YTV0d4Q+jzxw9/bHZqU53dh3NFBoSwj3pPgD0v7FemMWut70Iy52znY11YAg4qy
Dyn779aVKXphKIqmVgoThevHIbHHHP9vhzuR//IVhAmb5TeLIEZsJdy8IsT09Ylq
ykoOmFAxnwTZicxlJ4CPMhfRNxuwOhXvLbZ910pTRwWjHeqJZ48GYQJEjjcUVu8R
XIy+ZBpBOoIu0vb3cHLdxh3oXPLC858JR6K3M7lIFwVUf+RvCa4LzJNB8lH5hgDj
7VGlkX/5xer8N6v5DiXR/ADSfwGGKPVuFB0ZsUaI2yT+ZxdLibveNyttbF5i2XRK
d2kWWJEdoiIfzJvOirP2kn5JKELeVN+/WHRhE9tX56cnOX6S7B4TvZ0ORkg5ZWdP
6sGU+E4GCQ6Lac4tF98XhmBJVkIwSEfcaDdQEe5tKvvYlSAYVAk4sTs9sGIBSwEL
dWOBhMPbBsdmz5UM4Z7JQbHFZlr2tOgHZrMCnOPKR6vn7JAsH9YrqQk5t7ii2+A0
ADks3bTIB4AsFlmLjBKsIt1T6CaYNPEIDsqwb5ExGrSqOLmZ5TYNhl6wEP9R4xZy
8ke5wGKGq8p1VdSXQ1i77Z0J1i0PP7qY29Wj69Hf2Dro7teGuQs/ruGu1+4FMOTc
mFMX2QHRQ5tF/glKxba3tiPOXi4zBkV6wwcqZXelUWDM65bntQjcQivDc60aEkQm
tVtyzFL7UrpkXyNTm5PODdl3jRIXd5Lgqlyn2dTa+6CMXHT+yh51aMkPXW1pZJnw
KLTssqcLxoBhsKz3dOY+LKUtR3oDTWLHFp9/E9vhSXkrad9uXCNtV6GPOWfPf2qZ
GlSwmd8bxcngXLv5MefSw2EEnt0VPG5ktVGgOcAnKmnbMDYrpOT+s0GzESKY6zfW
qVmrPbulUdB8vorNy4t6VubbYCeqHJ6UM7Piu2w/pyJMlpt5nW0/VwiUJpHa6ieL
L5y1IRW+lGgmiyOuWJqqAB9It2iYZwt41Eub29yn49lii4hs9inLL0mAejh+3Vh6
zmLTpP2qz3l0XEuqX8dP4hS2rcVd8S6GILV2+VDHDK+G+8RFeNJ98O41IbsK1KwF
wleO5EADoZgRAiACInO25CIQuhbOuYSCGE1zRks+eEjUxCA8wUyPpk0Tj8X0Gybx
sNnJkBSs9F6E0OKNNcOOCOIBMpMXD2WmjOCCii1PsuBXYPPhdbrLwc9SFCqpPRTQ
B+VkR9Wz5SuY/dSuFa2oVPZoED2ZdeqK/50q+bMDIddHajsHF8/t8h8orwlfg+8e
r+PpKS6/KA/VqTKlch/Zi2ot9jbpo8qg24JTFBjWeC/3y1nU88+TTFYOGt0wo82B
cOMeB9hvAIslUEUMSGx8tO84ErgfSwUBCBAEANjiEU2zrFamii/8pjLiv3juaSS+
`protect END_PROTECTED
