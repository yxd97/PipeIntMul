`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIH+yK0N5FwNBJQVnOXGDxk2soScOVNoGO/IXNgYffCFqDdnxpsEL6xogo0XwqJG
msuCVhQ00/EIdmiYjsWLRWiGxet5DceU3ewwsAVD/pvK9vNR8xaG1z/hMV1nbURs
j9gqiIDHgCMQROq+tXGzUdJFSoNu9Jx4jWYcCIYJdQValYmMUGbn7TJ6lES+R6ml
Sr1QDui7GsD9TUMO8lyrf5TWpHH4XbQaGlLPw4XkKyfbkOtv+OfI7+81vbyuUKY7
`protect END_PROTECTED
