`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8i939VY4Fqtkzi5/xKAkHkTEZ3JvabIzXfrJbrQbsTuOfUM+ZkZ4sdD2k/JK2Gg
XPmCsY6VD/irLXS0pNZY2t+WFXVSGYYVqxtBqvFzB8ih7fQKrc/qK90so4JdTfjz
srNdVFPbzk6beY9gDfIItG4jQfb15T/EauBK/kcim2rwvzi5W8t+9NlbV/jP0YLU
8OsPx1PMAwHRjp7i+WnBSHK4xd6UpMVcCfHiQvvGLNnuOWvsQcE+eejwHwP48DA7
2csGCoSOOKGlRV3JMnP1D9wrv7j//666WdhyGPaJ3AdVPVbHK8CI6q5uQqRPsmGy
`protect END_PROTECTED
