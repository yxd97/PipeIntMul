`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzGDtGVK8NF+4Musc2BtGrO6ZdmrRAeDdS+s+zplt0RLCYrekM8WpWvafA7tq5TY
jbmDVecgfG+3QWGWUWFapX4KvndoQ+olNzAEMNW2kwyDhexeMNXL/VLEl20UcMZf
MXgtqaTBMMlKbZzrmmNHlYFENqOBjuACQ3wmaBjRZQw5ondUHKNtt+dVVvuG6Y4M
GNe6XjJTvb3rju8BwDMAioctcvHjkKmQEl4bVtC6s71MHB7GcwD4B0hIwbtCPFyF
+uUAHcIgSmr6b173otZ6jcZdAhL16NloEcm3CLLDrU2W0UuR5esg36g99k30NvTQ
Fv9PtRp09KKn/x5yuLuBs4l1JLjZwcsCuwEiQIwsS/X+26Lj0azDvwxD7bjY+ef6
`protect END_PROTECTED
