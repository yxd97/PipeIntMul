`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tEJswg5lghmIaOFskKvT0Wt2GHWdOuyO0xK0+RvHjtkSWcgj8ZO5zCSwIxyBUNcC
pQK/DVVf0ADl16grAA3jrTZhvLW6V1wFGXOR8pzR9UjeuxX8kDZWDmVY14QcOhn8
jEmIaMtp7Wc+h4QqCvJLtCjKRhcC9YvxvU9vK92YLvd9hoyzKkjoqkiOEXZv4XKK
+GPAZAQ97VAFQNDG/A7S4+LAdOGHnejVMl6HGf6wHL5foKn2W/1ks+TvjA8G3X87
8nEWkeh980DrGKypC2K8c51t105EGOrNGZtSZ6KrtDpC0QuI9IZcL48b+R6Gspta
j6M5j9J9SDlMWMuDmpAZYrzyYAHWJ2SD0eainmCC+bKKr8NJHeK02oCoqnMqwEvn
Yz1t/zVfZtrWPH/ELe3dXW1IuFTa1J/5imHrkLYqGYR77YqrGqyqkzwJ9qx5xyX3
Doy47JWMsLb5BEcgnHJI/qukU5l+kvf0QAJMDCx3YxBbJO7C7+T+BVu77QW9ZqF5
BT9C/55WqzHka2Gz3N/bI3IuxtEtZTrgyKqMex9KpF9CaSTewGCMEMu3Yvwnpd+I
pI6LoOQ8pXMQFpxsPJLZVr7RvV0FGOg2Ot0HIUviG9PXISsVpi3FIStBIDCRnh1b
yWukbdu2S81xAIM7TCUCdmmoFww3FNlNv703u56N2YshjsPiSW5EVTxCzqtOWAAA
ClHRBCtwpPHpEDlzYRxS1notD+oiZwD3tOolawpH0LcfU48Xqqlb6Ia+CLj0cGVM
26X7fDwgJhGUYt/iolzc+RjTOZ2gOWXkV6m/UDkmxKvR1scz0ZOrhZ8l9F97B8dg
CYTaXc0Ma0r4s2+jroA7uXusSOhNLHp9B1x8HK/3CNmv1EYiowfAPSDCtVRGrQvO
Q77+Bu9x5NtffnfqFFYYWgmHt/3U2f4CY/78uNxO/ppqba9IKlRJY+UwN0S8vpPj
qW1qsgeZAW8P3mab5SgbLPUuMKny6gNwwRKB1Tl1njbUF/jyJzVggIURc58Cahaz
KzrLt4slHGNg4XRS4wRS+OG2Pl99O8RGztl9R9NJQHlOuq2QcY9h+ChaJ98PfBiU
u3E5hVZIvgPn3u5ZNTQup7owrgX0h8PZl4Dp4cM/uXw1BIxVqtEwn3zCXy1XoOxg
zO6VX2aw3rwzWegS3EcAiD2qMF69M4PwOAUctD8Iic0GGpsmwMDoKr4NwSr6l8z3
EHDuMWUOlUwqjeNeibqDkqqJMpBhr2SSQab+lLufQ42OHbPhRySU5UDYz1hFOHPm
TWYw+XAl6aW5NlXwKmRYBv+aW5Dp03rh+LvvFPnoUXwYLEgEQ8oc2dkDkfNS380V
bfjcgkyP7NhgW0aF+SDRPFrKM6w3lQvv3g1AzG64yVxEt1f3xpa4Z6uFQOuRS8+F
45sN9vrxd+cxnVQ7wlaD4rKdduzxsC655DiR4RL7bP9KENrkC6MTUe/5TY3EMa+q
mZuFYh6Zn1gWaJ57diPIFQinvl8PdrW9OnHfjdbYedn6LQY/+apGgd/aZ89+jTpa
ej6HL3ziuN/zmEUHEup+1uMsIPNDvk8pEYLrOWGihczRi2JgA0auT7zOHCnFy9eM
jncNeuGAcdpv4cmMMQg8gO6/kV2P5yJtff0jm/CnNn28oNfT3JaESe97vifFdJAw
VX6tUSzy5dQhLx+yv85f6ei/UifcwI3hdb3TAkclATkr8FmyDuEUAOSU2GQjNqZ9
aOFwXrygZoZllr8zJqlrmG8uLYZRt+gauGTMcSLaGoIrsilNtf2m39N35ijuVN6g
Up98nx9Y1CKeY5YnFhv6C4VHUhcM8K3bMvZ4u9QURSwfA8fCqmxLKLebYhcLw40u
RRF7P+d1U96gYKhoZmaZAw==
`protect END_PROTECTED
