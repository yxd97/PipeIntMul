`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TK1v1Cq7fQFBsQ/TDcAr0lNGXkJ+QG59wgolp9FYUbQszpyZIe9BJ9CL4iPM9drt
OeHyXGNzoUWiDRuqby9mzFVDnJZN4Y7AnhHvsAuHFjt9/KvO3gZ8/I3ZbO5ZpmNO
TeK3VJPE1xtY584PS/h0pwdYxXc/eFlD5GHS4sBQ1V8SFqeX0llOm4CWLz+gVzXt
sqFtySJoVv1Bmy9YS02RPU0kq7fNcsh/U8PDCfTn6zlmIhCX94VmM7FUsPMhrN4W
jteRYUrKWy10lkuHCTa56y68iXVVs3RIJq6MdDRVcWYHExjAsYGGi9JAKlvXKk4/
GJVEZYLm0SyCU57F7CfaFtGD1KmRGgwgWc2RY54cVWp4yXq6ITRgHPTouulx9nnW
K7fjTY1TvETiazuFl9tVOuHdQ+yup9sql8+t27Rr44QyueCyKgB2qUY0bYJwqY8c
Y6WOUrVrXCCD5FROmRW208PQHtMscXagjfR4sBMdAhug6fCXRh50j6wMTgmyK4MR
DQzFWPf4O4y83qkbSPaMLe6TrVlfYRDrVHFrlEGGNXznVNJ/6XgdRRn7qHEr9AsT
zxkNEiBQi7hNPuOGr22fu9mbmgA0oxZ5Y157CU9oKRFhQZfakkW3Fpz2pFx89yIZ
a/TTcRP3qgCvTOHYG7PrTQ==
`protect END_PROTECTED
