`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjlghMsFSTsQVHOAWneJgKWqTRkEo2kV0ZsVl0kAJyP5dOXdyBMcdzuSc/T11+nQ
HOflDczmweh+nAurj+UvWSktFvrfeFA+DXhw7jrSmsB9Q4JJrjWEN+8YEVcb9hPD
j/CG7P2bkNYn0E7776mUUvIdWAofK7QjUjm4OKOuFMuMe0sxbO7sfWn90oU1LJmZ
JmlK4/xUdrBij/Z9+tkOFzU7E8vKfb+FBx3nqjGYcWep/S5qvOS7BGmvT2bUfImP
A1/5W0zwXz4oIO4I8xdmKXyGbEMn+OUrU5BB9iQOFFrtTSlsDZNZjhkyztojvQDB
MfmNW6gblBFIPk9kTTom5u4usUBiFqzqvO+DkQ3982ymlzp643QZGTK/TH66zM8L
cUDrEHuatj8EKK7hcjFiA0NP5sWoMXDmJZ7U6tKYzJMsm0X1QF6qhYpq/b1liZA+
vzqUeQ3zMh8xzXrEIF5nMxQZVTP8IXOf+9tKzw2gPJPP/RRQHAFhW99Wgj7Zqx44
JeCGsSuSG3xgSFPP83uPNFPUkwjPdiyspHZseM2lvVjHVcmt0hP109Fzl6CcGqcD
ENfJgPomVz6N6oTqbNYQ+gsWnJ2VotPOw8zQ2b+XyjT0tYaTI5prliO9HKK0kias
v9Aocv/2/AejoSgd6DmuFdkq46WHWhmvayqIcy5qO4gGbzxvWvcF11ozMj8k98A9
RnAF3tJj/wgN7pTi/y/N611g9pOcUK8asgovWpCkBDs=
`protect END_PROTECTED
