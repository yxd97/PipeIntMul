`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHv3KDm7CJnbzBNwhOv+SK5rKZ5aEqZdHGOQFhSNnapgZJ5Q8pABeljbt+rqOkLF
hyYQzfarAJD8Y6PSDPT9Iz3I1CY2DYOojwWH/4Cb9ienoqnboRmpATtKZcz3H+87
G/5bt6TG5gkACjeM8io4BQti1PJ6MwiHxC9cWeFWIlo5sD95GUheifoNX+SBFNQx
JR/Mr58gFO2Jde+1stsdf6HqSQHhelzOA3GkzfD537hSfLQvxtHHs33jLvj26FWS
9tuBsCj40uCwybvhDl7+4vztoamh40Iv8ceYDWlApeYpMu2XLbmAaGw83LaOds74
gpO+2f3f4kVVS0GL2H5vCQnLWoJDQI3pRpeDMQhSa3wVYcYHnlvryqRzipnQk7D1
n+b3Z9BolkE2Da7rFimvZQ==
`protect END_PROTECTED
