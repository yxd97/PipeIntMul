`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FkTvme4i3WkFU7uEjCpMVWrr9aXZUkXHluwDmXVaaXaNFaf/gHKtbm8kIvkMKnOL
VR5kBK+49FkaNcI+B7AtjFZK9W60G1E0yXoat9kvgmvYyPhEG3mJzNajKulyqjhs
g/CCeGkFAyiUTNFa1ft1rV/9ReBJxtUyIFHqLe9rr/N6MNQaKhMbe6sL7NzlA18d
4K6FqYaXXQ10kf90cifLF1ePvaVibhYnJKmEMQAJEXAZsmDs475+9c5iv+vDRoaR
yyLu9m7+L7zM3IQN0BLw52Q3M5Qry5r849OYeYZFklfeLN8y62T8yGu+xb1N+y+9
GkUZXw5AopSucJErOaUT960MHoCYu2qNT1x2s6rSzcjHf5mIdLxNiOnjcVDyW8Br
TlgHoLsTBYFQdN58+ou9wUx3LtSlPexhQyMrE4NpbGzic9aFvm7avUVW7OU7slEW
g69WIdJBkZk9HdGBtbws3kNqzYmMVJLYz4eLjQgyRUbnVjLcp9o3Rd1tlZ4SR/oI
+FWjO7uK7gxHmsv0/QDO8+Tz0XDkgWNWitIxYLT3cLvP0Knml5+dtZkrr+LwC++l
T5BvBIytQzRv4TnDpejV5ccxNg6YGyTPExZFBm4mnyFbYdhVWohM09/1CCYCuWEn
xafHlWT58WWSzub3GcVRwVMyjxEyLABKcT2MmJc2yBWJ1mYnGXzPcyUXeKx3A2sX
5YLcWaCFsfwSpAaWGFHJgtj5ef8SvEP5jFXmel4loq1fkDsckrNllXPtIVIgH5lq
RlQSDzbMkFk45O66Xst/gg==
`protect END_PROTECTED
