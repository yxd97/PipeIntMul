`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N8XgwtC9SrS7TSTEvR6aSUPjlpbkGDwbPFO4xpz7qZSCn+2rO2jEIte2LOFKWLfy
++07Hcgfqa4EGgKALayhcSbvoSYZoSSvG6oiqs7MV01oqIekLVP9KhYBfPzMxT09
VVyIOeDIP6B4Jr/3fzjywZPM+RoKk6VFm3N9tLMErGLYrWuSTAZUZ49sskslTjUJ
CNUO+VTn3aoJJGFZCSwJiK3+AFPs9f2bUNXsmW3dEZUjbySIaGJa/as/jQ24I7Iz
GKavbgDaDcZJr4HvvSSDGwpSfgdkv97wXIhG5xX7fmVx+2FRP2aXk3M2NueAzlTj
2nF7KX1wzcc45xi0o6qBf1ejFWaMHAW+4KJ0AOP/li21i9fuvWm42kvpcvhL4UvB
U5h7p80it1/cwjjF6gqYXhXRDg8yE01OxUxRVqkJsV+SxV0x51aj4yBdUys7JZeG
`protect END_PROTECTED
