`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ManhxiRbbeZzDbKzR01x+lN0zTOydzKcQVSuckOKML7JhQqhqMPhD543BO1m9XJy
gDG1yUZseoWCYfsH8uRgAIsSRleOGY6AXTyklqc5w0vIz9I6+IEnjaGofGPZ5AIW
mUnppGnj0861vteSJm//chKrUSCI+VHdgEoPqOYXvAN5mhBLUW9CMHBFeiwTiHwt
AADiNj+NeZ5BodFEKv2GU/ImghRbtU3RwOdofsDf56gK1Fq9mmH/o0NsykwDjeCH
0DBGSTIqXmCezCKxpuYR1/9dIYYo2YqmwAFQ2D4ktHcm9nPyS2TEA+FCPEIh7J0f
HztHvHrf4m7Np+mkLfpRHsuACamfg3RlVtM0nuZU24uQFsk+LR0BTJv04iln6h+P
2zG+Sa0ktyqJUSOP8kiRjlS/sBCksVgrlnQPzNAYBVqJRfVnBUE5RCEwRYsBcdja
Q1bu2KIOpcSDYl76iCMfjAMDCLfewEUckeOSOxWYJ+y3ZSQkZEwBfwszU73fgEaH
Un0qnO3m8NRfzLqLXDlK0UmXPn9d5EpMG56IOeJokVTgvI/Om9O8wfkKajPGNcVo
Q+Y/T/QXONe4rWLe2jOV1Ll3yP2bOaBULirzr66OcI3I/HOTrHac3mvUmdnLFojH
Rb0FiPkOSecjxnzVHZRODg3B8881Kveqvl+A74pUD1o=
`protect END_PROTECTED
