`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gRjIu9PDig7oh+U2CrjkeK3GhWOl5CFSeRLAi3ybAOlF5815u691WQDF70vSELHU
toLSQPDRF6IfsPnHibO9j+RfDKeihwuUVRgFxY254KNn1oD7pi3TJPj1QelmtC6E
IASQUnCaNbWRqGQIPFjZgNV40/WlWbTDYuoXj712dioXaEQWHaTwCpKRcQzAXacC
hFWniwcvradzYxMUztaJTHq2U39Hb4jZuiE1dbZuVdysTQAW5ABo2uO1zQeDBP7r
QqY0PgFinzf6zaepnScr52mStXIfYLdSAO9cvx1m9hlrCmN3/2M+ok4KRv7jSqJ7
uZwoP9vOW3rra2eGwILZLf71IagSAVBH3L5AEqqGW72PqIdQMpaCF+Bpl39pGk7x
k4jhmdpGjO7Sd2AY6dx4X6Om5qgHTZeNcgwX9MRfds88NQXLqdhGF/T7jRulaE6K
HxTnpXIwarL9yBZCf7F7ZluNJF2Ccl+eDzmx5R7Voz8PYGW1EkfPq3o38GuOW8L9
+j/WjS5V78gtlSy9h86RemMR1BfNhDayA3IO6OZrRBg=
`protect END_PROTECTED
