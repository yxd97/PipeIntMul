`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afwF9ibka6+XLKgiVYqhJYiXgxhHoEuyRfdVy/z7Jl2UfkQl3rDRWH/9fOBPvY7K
otHu5DJf/Mpv7KAInrMsspNHnWsfjEy98jErv8iByCbyn5YDt0DCcsa/Z2LH399Y
iExZ1V90GYzsXCdsO19f2xxIwRt9o8UO9MVN3gEUK6LWWOa6q5XLQ56GIwYslh7D
8c2o6i7adqx8j1FUdit9ciEiXAJW89S8kWR+ExERA02UhmMI0GCllAeR2KdKHsCm
B1r9o+nDFvIXlAdZGp+nWJXx9CA2cuRUHhpOSdIxtEQb2VX+RaHhgA7+uFMIQJSJ
RcM6Fd0z10vAXKxs4FvkWiyedubFf/SzWNZD02YsAWNZkPRVKR0ngUYMVTuHj4Ip
u+cggJuSLcEIpcBH0YiYCkIZvAoPrp4R8PMVq5xly2lwcdnwZFAPBPO3b+hD5vBw
UHRemShs/Cr6P9XoPzBVyE9vI28yywhdxo4AvwRA/q8cQrtTdLyTM+gckhWk1ESa
`protect END_PROTECTED
