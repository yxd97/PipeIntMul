`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hX1Umz/7E281Tzvqdrk9PXX5WSJV7GHwFG1tZhSVXiSMOSXx+1d06fit3gSdheFz
SM+hMDOD0w7K3Dut7UrEtxyiVF5zymax5bprRieHHo8WAF5FCd2vt46BPhAM/jhu
e9b1pHi95rQJHL80Bh0rS7NiE/H10ObDA11/6doMJ6naz0AIh05HiAJD/kJ5pAfY
DoYq8CAmyZsbChXfapTbzbyOXtAEWuG2mKe+fFIIDGaQweRs7Qnbgm6FE5xQclOE
wfYtVcSjHDaQSd0t8gVy66Pw2VB58oSTHBrEqX5JdNVTc/wDtWtOBmfz85/FvWAT
92f4VV2NMrlZLkjcxfc6Bg==
`protect END_PROTECTED
