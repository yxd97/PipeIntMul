`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4RE+AtPaOWWa1SiQ0JQI31Z5qi9FVzqm9X81J0SgBc69WPy8eXY6Ix2zxDUKe9kS
6fD8lGNp2gHDh1oRlekauCVJGOrBfTGCy0onr3L2VTvjWgG1E51ckVdBr9nVOAkd
ANrHWtlV8x8/stssR1KHYWVtm5xZdMFPbfynZ0O6LKHq0JfArxHLtLlx5hlFT3Tc
3HXoiUyg6S/zqFLTcib1XAjhdWXi+Kt3/rYcst0qe/xk46UCIPHhNn3cxmnnx31v
8EQtKIgnTLispnFqbMv00JWETxHYUXUTCihY7GVT1pH9NtL09tXGxdGvk249+LtV
qFdn0mtiEe+sU90860QBDg==
`protect END_PROTECTED
