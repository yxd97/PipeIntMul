`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38Du4ODXKy+fuPzLZdqRkbLEyAMDNw8L/xPpi0BpKnQvDjgHaYFM6oW208eu0SKn
xGsoFp4F8Mij+QIJ7dEt9siI/TncZulsyavG0Q5umxEVtxHygn3PwMhUmY6Di34Y
5N02AnOrwxWS9gljcqfbbeF+yAHkYieA8H0mSSOd1WesRKpAuDabvyYkQG/S9JOh
xy2PQXXhbZqB8KWwUhHZfb274QWFtDXtJAOQx6ov3uFoMW93GJyKkZUH+jv86zhz
DfZzfGl/GJBcRxg2uwp8BoCzzWApGoIwhJe/0sHI75BdwDQ0Jqwe99+FeXjO93gW
sQ8Tx6rxLWCsPGGpr7T3u7oBybckxhHWCDRlKuMfjRf9sx/7/p3ABRj/+4lU+6j1
eQjCScoWgvYvXgZ2jSrldPbTjq5sTrJEFVe9WNlXW4cUoMB6TVXFDr0ezJprGa9Q
6xAibWKglbbEII1akB/LfAZV8Kg0QQUEUNAcSWZ4dsNc1OMdiTusUizk9VGUkH1E
4/lOeDizwHy8CsB3knVVoyTrkHF79mkKaUUmGgP7kOPlkWtBGqBUocwaClvM7ntq
/aYQNG8ypuqTTcllcUWnnvctPw4UFtRBoMfaCDSL2BAUmXEKafpWIrp/rVXhZ66L
I5DiQICs7Ukh/yfH45DP4ArVJVubWRLt7G7dfRmQeEVtsLl1ktmnldQcW/NiIVov
70WCmDBXn6xPdH5+Uihq0zu/cpgsR5t5nlmLxZq6vZdz4lzE21nICfJ7UYw3l8M8
B3TJrickvK3hT5SHBHDV4tCBERtGzqi9izfTf6YoJiGFj7GkjCCMD0r1XMqU7Hyi
PgjBiD0CU5fbCyOgpMim/4h196yw6Fc5EP10C08YM4XYJ/FlLeYPYzl7bK6ULoa4
RKGc7na1imy7gap5pO59gBIGUTQz9G9VS65f2TFNMZT0ix5WHGbDespudb6Ehfgn
RYJwIRhB0AtzsdQ1YCmM27pb/1c4AEnVf1tGoxrwk6NNIcS4PvSqIiljrSL3xOJx
Du+uBtDb/2JAybZ6ALwTtQw8Zrl/nEDnp4HeVroU0p72w408R5ZzEcTTs/EfZVMo
/8fUxBZIm+OTl6p3N11qz1NfNQePBN4MXMNFMMb+9AO15ynyES43fj+IwWf4zWB2
cyTPxqkJrl4Dcw0L9zrcHiGfqLO1Ui3IUTf8+KNCUf99RrVLPz8/pS/nPQBnh2XJ
RqEHY3DDujNsI3T40ZB8rKF0HMSX9LSXH7t+pLC7Oujz6dY/ftCR0WsfiGwUfkJM
Ny/jZcBa0dseBvETrff+LlQIqy6KBaH9RkdnwoMjTXykwSZ+3qbAWTwZT+8+ZoPw
exgAcqbjVvkjoEvGBH/7Vw==
`protect END_PROTECTED
