`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BgUYEFz4DT8S/jy9XdQUKhDUENN/R5ZCHAAnufASGrZqS0PmBurhmYCmo8ap3ctG
dJ3fWmxiORc5c/6vicbls/oN1RMLfmKBK6nBxar/jbBGr1+nLIZ1x4m6hTAZhrbs
XPzNeHyJMcWVU3xRy0fyoEu1VxHA9sSXx/mgDCTFI2vlhZPvA/V2VmSBxM8NbVnH
9GZ6i+055LdCO3EKE52dt1qgr4PeNx3/xE0hLBdOkuuMA1B+uDjZrMJka8dkU4Os
b6p87/qlqAJ2A2ca+oqdXEFCegcaH3EoB2NOS0o6zxMkY51n/jo5kRil4XhdZAjq
a9nXKG8b6PMwZLRSvBi6LGOQe2CElSg+PeQgzQqGk9n9elPxwVIleE5zDXKk4EE7
qhO8CA/dqCERNHmTs+Hzpg==
`protect END_PROTECTED
