`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sl+lV1GVKbF5qQte/SXW28qD3uX6HccqBfgnVAVa20W2OfWo7804Maov7Uszs2ZP
iS3SSoGLuJozo1DijZoHBgVlQu6FwCtvHEHfyASxWCo2NcCEzpsaNooiN3Ocjawr
YuXtU3ykG9JeVBy79Q6j5N5ivlRllrLPGVV1KBuWYE7FWIJ+0uebnWDQ63gFXgdy
aFfM1ThfrnO1RcZpjCsaKVs/GJ/G4vM1UHX/0g4gxEol141n3I/bYXXR+YjaJyCs
bB52D4foDb3prmjsYM6t8m/w1pbwUFoon/sxrGbdWMVNtG/WpvKjyvu3iaJgLIRA
0qTjWDMlxHKfGGOseUi2GtV7GsKlOK5omKYGrnr52C+V5tYDcWzxK1yxSmnD6PGE
7HDjziEyuNan5ruuOlJ+/k/JBNvwudvFa7oxDI3+1JvDYDwuFqw9UZ1xE+mrq3DA
P+0ociPd3NpZoC6VWXrLLUEg94F9HPUytQJPT3b2c0t/kMRieoWSK//TIGFrQ7kA
`protect END_PROTECTED
