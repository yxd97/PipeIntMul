`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6A9D+iedRAD7DWFerifhz9RAmX4Ea1a8zaYvgYeEukzEc8P79M3wSqtDM7NXvTVp
z9oL2lhlyiCvU0TiX+tfj5e/X/DgkFYiqK/0ZpP4EdxYpxa/Lbxfl+xIgZzVZtf3
umHp50W47aBqwsd+EQRmmZBczynFKM0kjMQh93RmwAk2ecwojhUqJtZOw3mwWeNB
70zIyKWLP1ave9qvqr3CxzqCqnPPe0LvIcjmWV8ZNn3MYChUpFD0N1EBvr2jDlxJ
7DCIoHYiGODXqpI6Vh0xnL7eERESRLx6UTpRGoc9Nm65xBiS1kNgH7PsTd1s4cBL
CxZ58xk8T0gIwimOudDLkyZwDTW/mYRMnnJC74oxIF6eJgB7O5EFdD1rtCLN2mxP
HuBd4EtqomqZ27R4zvM/i5AqO0oFZytTo4hTm2mcJY0MEI57L+rmo9jEJ6aSlrlD
vhgsMcalopRrASfxfOlSWrjqCGs6JMgViH3D4eGeMbc=
`protect END_PROTECTED
