`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgYzMEDMw9Hy3P4UzprdlY0UzCYuhbjYn6h4/nOn820GV6Tr0s4vj0njd6fCbeCR
nAsEGCdAQgtSSMGffE3MRL9adyym6jl/w3QtNAGbkfNbKmFP885MNxYRBEQhRW9B
a4lAuD/QGzj9+u/MzBnAHY76CrIOH2oXNQdq3sc0cnBgJPJFYcOh2AvLhcJo91GH
qTgiID4vvmKSD2dgBeuvBYDSk0s8sjlkwJ9ta2uPUYcocRudnTytOZ3hL2LIm/ot
x96BiduVc27q0VJhr3Rp+XGrFGvvCsIUkWLsV27rhwCLWFZY0PpnuElmVmogxZbu
RFxdVB3pxAdgjjM2aUiQhscO8w9ANRRAra5i5uq8KLUfREs0xUB4GcY59FWoV4x9
BFgbGMXFXbonVKPvOCHJ6fT2WkA2MDk/usmhhZ/iC7lG1vKuXmZq/Q14vncqEqWN
kIbNRrusdAlIOzf8BqPMrfcfzdKbm5GQhK3ArGSj7xO0YLJtymYLbv12S3JnWe1i
Ev0owN4StHbLdWfIvoU/dVUrq7UsbQWcLhDlGdImT1H4oGVq+kjR0lucb0ysF9wd
gycp4/qz0VBFWhhHaqGA2T78edsw6WRb9OGpso5enIXLEdh640SsU8pmblYVQ5hi
XGwy9BWwgCZ7vZhcShnKX0Ecn3x9asi2LWHGnxL+T9HbCmE8YTBHjnJjoc4ZwgGd
sVYdF9KZI1ce2IlOOn0Rb8BgM9EJB+4HmyBY/Z0wH/ZjanpWn6lzpA4HPd0dUCX4
CKyqSTWJCoTUaBEHmRGZb3TViGg9tfNAFgln7c8wZEKtFRxjXQ8WtCIJTVsI9k4Z
eLo3Pe4VLh3glkNZrDmWiOT01v1tyANlL2H99TjMPYC1jQjW5HkkP9WT/NsYh9z1
afZSDUjab0W21qnS/cotwnwkmrCm0tEffNqH7fnC8sa6f91xjmClNtzFY2HpMsRX
GyeqN6hGlEcacOc56tbt513v0WzUnESecpk7R9GxCvc=
`protect END_PROTECTED
