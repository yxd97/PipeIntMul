`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qE1YM5XPSG5m2BkH5PS5njrQ+xg2ZWT6ZvTmTyDKpRhzVCzyMvfDqY7axLSM9Liv
Zyhypp7sw9wVEb7Dn9YW1XrYQMdt3HWqLMeL+MbqkM8Ea+/VoNDFmr7E2Zmgclpc
4kXaQgu7eMAfj4LD7Pq10/ixzNkzkUfvTgfruNy6mSHqCNP+lSoCf3jHQphnTsfu
r5pFVpUeqjPzRtjQjipNNoldyv/DcP4nS59HG+a7HcS5X+mto+uBGuIm43ma2fZD
8h/7zWNek/BWL++NllV3QR4Iuslzoc4W9Qt9SGJDHbfRekE5wnYws7hj5LYTUyoA
6HDMBLji2nRRsr4VRam03Q==
`protect END_PROTECTED
