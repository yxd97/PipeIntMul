`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S0shpALHOwG8hn8GIskXHJUlu9NAJagqI3h9DAM1ul2D9iZBa9t4en0S3+ok0f4J
cWsdYoY9PD9FJM/SJDHUzF3hTRsGOWKECB/Yw+CyFmYWG3KDhs7/Vi+Qi6UHGIe7
yrbPdi1HPApLq1qjM2meo3uVqvwmvNxLiG6vXs7mKKMEs25nxrz0DCzMVONHJJC6
d9WskXEXpQMhNGXlHWHfjjRCh6RVOyHEIYqRw+mH63QpQRupqQmpjNpEb2KYwbm3
/rJFo6eD4oj2HwGi2GCrbpVGUtbtpW9PLAt3qhzlUqzALvxeOEt4m7GczmMvl8RU
0aPu8/Bs8Cc319Y4jgIoYCyZMH8wWTOaJ24ufSOjjPBjqCp/EJIymQEYDMCcP4Yt
u4AsVXWfpdQqVEvf6051p3rKUgArflfEYfJPky9t64nhgsvx14aLFoegSGm+ggxk
RHrCOVDuAqRvP5Hrb8DfYqKbeu8iE6yrxJO/D6qr8WU=
`protect END_PROTECTED
