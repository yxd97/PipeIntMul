`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
48gw+9lbMAppHkAWnEE32xXXPuLfg7+l5IeBMZ/2to02NLi4Bl7xJOK/5JA0kLDf
o4jJrnrjuDXSH/0ViCIZs980BZCfZoivxwwaQHwZJ3lRxBx+ndOpb+W2+qYwLwv9
1tTMO87fo1Q9igbWeCOBVj6iSZWQM7GNo33QiLfFUlwuWHrhWETpRdI4EGGTLABm
dTELxGexUZtSO/r5R4FzUBsgLB6LelJh/AoUIrunpiz34flbJYQSU8Bi/32zme4q
wOcR80t6cnBp+BBH9ZsM1ZKtTrbZbanNxvJPgyu3hmZOuqjAmwHoJm1xVnNIgbQD
7G/PqgQiQJEZupJJ9RuJmYTcmCwYBuBphCmx0JuXdbvKaMBzrR9cW9bYXq9cvpDB
1fJqLS1U6PybLi0xx6fldHuEyftFpNbzkxcoK/K71n6F3JTrm+5kse4JV7IfvBSg
ccgYBcSHxzCGyvLBz3fTdEOOwN3IphYVLLpPe7qCUvSU2l9gtQA5YwCKGBi8RiMB
m6AezI7dZLqItPhsfV7kl4SsjRRiz+XTFxg1hVHnGOfuxRmG4ysWl3nxR+2f6Kz2
SXC7Z11AL5QTJ43vGYrfuauiiNAnyaXsy9rGATrgHLYbwzwZFwmpxoSCIOSlEWYi
4t94DvM+ifYWaidZ5AhJIzF5TwGYiC//ZRRudzdVhP7etDQxzrIuRfGvaDe8DlCg
ALkW/jGMDjsmTjK+s8djgwP+cefNyS/7GLvEgFuxR/LETL45RRMPQq3g4IcCPMCr
JHsEeeqP4uyvU3NyiMvF8Rk74Ytqk7JWkOhXd9m+tjRmNKxFuzyYI4sXe6R6ANj/
RQsJZDaIxE1tkr+t16k2jGAgCEqCG8m2Zad011E9sDIwwqv5gBHpLrWtn85cNDQS
lUNTqu/XLTKC2sUJ3VoPWQUYG5aBgbtaJxkV6cEcxt4Tn9q8Qi1Unzd9rI74+7fO
vVL2kUHbJEoxqY6KQ+YJ5wW9mWrCKgF82S4nM2mhK8biMTE96B1fgtXlKs2ZxvP5
4TXfpXVvZlubYljP/R3/mUQTmeMtHEVIZmJ9oA/6tq5M3reEhD5jhpghVF3DMKG9
098tFXs/W/iZ+vx1rQ/EeWTpicR4EPm+Dm4pSCRLjvbKNtRL4Yx6ZXry9m82j5ge
1owM1NTv15r/6sGXSSamjBtITiF8TELWK6d0eQbqjTFbGtGq/grx1DeNObVXSgpI
NHZ8jMPvCkktAbncvt/PXwdE9XeWCyU7624Fic8b5mDb8Xswkls0H8oK7lnBBfOB
jJQpXfJRW/F+bt9/WJUyOgL2OFB6Zdq2imokMnjTmWHp8AOL6c4x67uIPq1TcOWx
Wav3Nm+cuYBx1dA8181HO18T1Or4euAWev9U4KmZzfT9zOH7AtqrxeieedxWm5Do
`protect END_PROTECTED
