`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBeHazKaMrqEcF8j+ZWYQQAk0zdIXknG0zxiUJ3ngW3dDodIvcn4YaeC5D9w37cf
zdn21t6xFADYUf8c25xzeMcNTEsLVVTrT7UcysPRq5inMp6JjI1bOCjfQN91xhMa
h5kUElsvoT7g8waq+A9h28tuYqVU4gn3MqTjZoFtX7C/jQF25SxmdCU3ODW0V8ny
S8orZSvesJZrIxzdevY/fTl64LX52VUkiXyiNIpQi1dFq0e5BQvpmHBwDlvAAG+o
oebeVGS7Nr7v5ER+LPcXuF4ist40+DAmpMvFqw6gtsA=
`protect END_PROTECTED
