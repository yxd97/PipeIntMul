`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y2Kv3oK7dDp2yV+qSdpB4OW8zrjbp+a7aY8Rpq78Wr9cxDkXYJoDavzX6G1N2mi2
DFbP+2PtKxCBV/zs1g5TiQuhJ98rs1hnoc/YkkpnpMOIepbzs0w5H+kK6qcTJH6W
4LaDTUX+TPDwLmGjH0pN8SFBueEBzg4i5R1yy70+UsOomSsv2V/A+hZiGQRRy9np
TQYF912kjulzX3mpy4RgPv+izV8nf/9O2GDibPxk9xZCy+6MDiTWeSSUXML2atG3
X6IUc1tl8QN9VWTzKBU4S1UHwH3J9sRiCrZ9dVE7XtEqP3+J2+yjS+ugOv409cDn
BOHvE7PizZZlIYpyzLUzH6Z3UYmMfDm7OSchWtwYq/7Aa5Xj2PwUa60Wxi+2gohC
qInfHpBp7sUoAfPrBoDwUs2fijnc/H5SRW7TNiA6zexmhd1ZGw0zxX4XKtOcptGI
uoWSX1kYHAtoWqYS0hJTrQ==
`protect END_PROTECTED
