`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czXQ1c0llzJoXzuznGA5t2BHxC3twAIM7wnxeNH0GITZwVgye7IAhQlinRZGPWum
kRA3wfLrXrPuQdXDiLrGoQ5iVOsMNL6R6z0ItNnE/Q80fkQvx2+x7GEXpqBWMhN2
5u7VjU6Wcwgv025XXgnIiPnQGFuRMTOR2YgQJJ11GDETYzqSRkhI3KspJgtYbpy5
b4JWjw1pAFYSdnDzo7HsM7iygrwUJYpsa5cRI0sM7ussFE3+rz9OTeLRxYw2jv0h
0PthFphm6R0PjfEz74T8z8F2Louz7vtx/rte8P9m5Ju7L2xyYj3iUA7ADDqO4NYK
7nzWMEtvnoXngMvOMipKIXzV2FaVo4X7WPtUK8xiPb8lw3GKpGsqPf+o13Xuwb5v
O+XRULPfVbz7f/zjabtyVSieW7E/yeJsNAiJO4hrMHU/mo25K/uaqVQBrb4LqwsJ
9U7x5mAL9sn91ZjEy8b4frsKSz8wQxzHw0DcQAqs2Vm3fBZJ40X4XCt7UHrOPOES
3VjvAPBImVAD1kLtri8zN3bBEeBIbU7OK3V+217CFTY=
`protect END_PROTECTED
