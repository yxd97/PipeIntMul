`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B7ZKyJmNsedO7lOYsLKDkSdBOVWgA+umhrgvWn4GLNa3SOmKb35rwSEGcDnTDzXk
r5NlRUIscjHYTdqqXH1zHx72MtmV0RMRqOktgULyY7u5B2xbSYsqo7NtJFLTcQAh
y/ytEmQwkM+dnGYthyInjwVqIovZp5/+Mf4p6//hN8hfeJ95KczcuBIchQ4BPKnK
l7NAqHkM5UIWV2yulW6pdeWFtafZrzPobNhxFo1cSuUgOHa6H6tIu90ZrLemxgnZ
nZKeOpVh8MnKa1iPuvHql9LzybN78j7ypvRVMr9xtAaJbccUtZF3iWdoRTTMIN/2
AnrEnaIlDXlwEjXqno/+YbPm6eqwH6FFbVWEZ0I9UWItCq9ItPuLCGoxaoEN2cyv
YF6IUHsJDhXvg0QTqTZB75qjrdPk3etXHXxR0AL975c2dbwpnKMDeJN1xaf+m9wt
Br1mSJrkYYNgX4R3SI9/Qz/rplx8iV/e4KRXyeJ8it895SXyIvD2IDcQb8mnLO75
ZzekRydVcoh/KQF9IMsDwqvmw/1Cih6gS7YW/bqPDv55fGNOgyW70jF/AeDuISqM
lGXphXq9wcx6HmyFx026tRcPXfnNtIjB3uktvuntbQxvIcUQaGhcoPB6oLYQJniM
5n1I0899869mkohgef+8Pze/LqsmUl8NTfbFcfFjmE6dEXPMJfEfHYjW9a6ynWmX
R+wOu8o7hMrdBcXqdwIPemP47iJR0Pmxczr0mUjikj0VpSc/7rPtVLO0RjOMlv36
g2peor3QX0fzGTaU+Kq+BOgcMonHHLI+iLOGC/w70SGtW/YgpjZU7SGjjj6iWlQm
mWKsof3N2aWxxREpyIlcDitGqLwZR3U9nZ05DRms2MMM3iMceBkbTiQRn4T1tcRF
aOaRzoB6WJNEs77ECQIvQDKdqGMEKwWD+CjhS0enHh0+sJ2hECMPKWN46+EfPDUh
UHTh5kMct3FHPch1kuThhWFv/5TgTmoV8MkHP7sDfCTw1pyG6EfD+38FmyE3/gj3
yCXnrTjQj50gkyaLe0MxF0GE/si9cQRf9UohEfK8woR8apZ+KGhwE6SR1Kp/0d4o
OOUxqCioN6GzHRH9JR1RsfvXusvi6AUZnt8IQINZsZsjNYtpCd0n7fwWjNjAXvt2
d/RRLyYQGllD0MO2sc5dhgfywQdzhDcDCYl/x0VhYS7PzsqZHYoz3sH6mWaZ20Tn
7ALR2Q9GukZCm/Zvnu3jFCT7EBncLyOYC2Ga4UvQL4DI2XkFEgz1bt3q8ayqfzwp
gcUWURukB+0281MTPawPBOpxUhB5fWmLGJnLI0+34bmRM1CAGr3ttriQBiLKP1+Q
1Ic7v+BqPI+Alk0g8MgGDdKkce1nA7WMmKaANwsprZnQk66dVu5f41cyp3jbEXWW
yMA2FjbUh8DPce+OWNpcFRcubEbEkU1NiuaxjIVsqSWIMTaYgLHPFN6KBguXp2L8
gmavwUw1qPZ+drpdOcs3j+/eHk5vi3udPTDHXIoRoMObUL4msqozdZw5gkf0/lgw
gslqsbbGd+hHq+ZMx8dxlSo8P1S0MJDRWvHVnLmxuxGkMS5+z7H5hKziSXEhnsnR
h1p27DfwZRlWltLLpm0e0uE2Lm7StmLl7m9a7cP9un+F38Pmjh8gb0+/f6rG+6sg
+fi/dbxjXQ/dPjeqBlo0kT7SjN9m9m8hOOvfBwAh3v3CLgnUEpKI8tza+XVg/fst
5O6x58fq9Xw+FcV3YBDpDlPG0sB7i9zqoKJP718Y40PydCIF35Zkz8fkziAL/5Mx
iEiByn+1P89ojqyoR55jnI+esAmXQCfl859RA6CDDeEqtakB314iicEzRIgBQAdl
XJ2odZwVWWyAVYRO0LgVu2+ulrJa9fl9KM/p29zf/IN49bq7mIrYzDnhb8xtEKxr
YuHcUv/DOGprJZ4L4gQmF0uCvFxL9bx6oDLye2BvrSBdFGKpNCh2kcNzDdcaTxw4
bf0ATteCgueq/Ktop+3HGUMkz1E8yVRDnVRvAOGXMaWcdXVfDM/YcpRe5vSwwtJT
7OnM6PYtum6P5/Vt5qmSMZl7egj6BqKalygjESmKmUBNiJnJMC9TjpxxBDt9r9lY
e5mt7xlWqu4ZTKUs/004w9UxGMQXmLm1YHupw+tOPVZhm728EKWL4srtrdYV81RY
LulwxKnii98psz3jksUfFWcVz8MBsNEWUlzlTNNhfLDKIwT14MTdi9hMWzkgAKsU
Xww6krMzrpGjXpNfXyWIaPnai42ansTENHKs4PNbnMBQ6GZV8qP33cpu3xKIoAJC
DsrPXn89L3qpisv0TAaGhmMcUQOc90RAMB0RvWYpXEuylWMGgHDYjiEq+4qrZ7Yv
ykplXsqF03JuWx+/OeJVEamJWQQSGNgIGkih8VD4hYRIXPbW5of7PrTMjP9L3Ydn
4O4jlKCKxozDg5oQh0R+hP+fYXrSi3qoXr6FJ0QLWObh9qwjWQ+shnoYlNhhUlZI
BhJFWHy7orGD+RiTRXCED4XFrW+BSKMb4P7beIeYkVmGb2V5EE+M3eMw/f4p7nzG
llwJEKmIYI9AWEGiNYIzcZmU5cwzm80C6VDJFlN5bPppo4keObSuRf6E5zpyxv7Q
bfGgLi8QBhDRKaX1uL2ToOKE7A+LvMdbMbP6YxTl5u+lUvSGSyXGcCImj+XuSAQw
gDmi60tWzoaiYM+lwq3pGfu553XShlUyaE702FVG8bs=
`protect END_PROTECTED
