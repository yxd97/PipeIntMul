`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGQUzUx1v4Gs6MqDBQCfkYBtLevH85BUewvWy0JHrljDzZLiJ/1gZ0oB4yKQdNX9
SPXlp9GRc/ZOlBB99x4Cs0efKa30+GjG4OwnnHh+OzT08cGO+jg7W5milKo0CPqF
bJlDpB1Wc23rm32ws5WBBT2DRrmFzMNRzu5MujxoliDhNBuzub9QrBypG5bn9w93
dG1VZUjDXH3bK4LqjGqKWcNz1P+VtjgbOqCx2mFjViEKv3fCeCoXsHvcPLCfYTmi
HN2mKVJW6/7lMQaoqY6GBwHOIHgj1tcc9Nky6/gOpSKVMScFmwulD3gxa4jQYnll
WFlb86kugqAH1qImMBRdMzjbkWIAgBgpyogYzFIwz7F1ecKVqHmUWhTQxLJk7d3W
EaskHjCctSheFBtycUr3xvNCWpjXTTyPZE2cHl7GcPmHMWf6jHEt83I4+hNcnDzP
bkC+mhCAmecAQxFjbHDUBJ7hEDG1znWQOFuBiRiQ0NCdG7kxNYYBZPvm0G2nLyM5
8eJtKatIJhTuDtCx99eR6uE4pmeg8xXr5q0LlmLByJA+7rWbcYsDm4m2pG1c2won
C5yyoEtFsm4s0PzM/knUv8zr4boHBr9oHwqMIPtdPoMpQtGI/1HjGBzV1uxcy0Sg
tB59OSe3/cRGUZ05/A2mh1ZvxGtRdxdlNRHMXI9EdIcdDGvSMl4zIef66/Zpbk5E
RMYPYoqMe4UdR6F8D0jECojkRK8t0CM5xChujKDNJDocZ8PszSC7+fJ8G63iumlW
azIFbuP5uZj1aiMo44975Anj/mSMGUtklCZwDQ/oof/G32byY/9gsW22TNTn2ZUa
pkzArpjWo+RoVhOsDIw2od9clM0HFUc/uBtH9jXsO90jBl2dLu/MTAK7+8nUeDqh
9Vn3oFRtTKC1l/oDxeKHKvCDOsDYHzMsSHE99yoPZ/ZokkXDIIZsLnytq+G4lyOG
l7sKnFcQ/o7MHbNWNXybJm/1aanFA4brEhtEMuEj4EkXMNexpluXR5pSf3jkhPwZ
fukMMlXNInTGlG6yU+SDVOKDzJvyoOeK5ZuTkw7FwMEOow7hcjGzwDkP8UGt+CMo
FodB66ujSzx8Ee6CkMrYT+vg8uwe95poUI8B/9z5VAIhTGwdiq6nlbLowT5/03l7
ZjFSEjY+pIlhEKXQCzpaHkg9DqbUOn+Zhc4RZdHaPUDIhsMmm+jfsy99H8smAidU
Nt0SsVoFsXvTN3BgcBQTmbebdwLFa2GI2VDiIXl+Jf4rtT3YAkvUGaDDCdaIhke0
7zKFHFfJ0k/AvLM6qlf475f7dCZLzHFje64o42TCidGD9qg4ypmWysgJsn2Qy2Mq
lR1hUosMj3cn1nXAl7ywO2l6wyp6Z5ZDwWBYsSmw+iDkikdqrCxLbfGwjgQ8wiWl
TT4AGp2GanljiC9LzscBXYuUb7fVEafGTRvuwCbX7GaGXaI7G4MN/d/44i787DWM
ICC3AuNsk0sHtr0AVEPOugn7P0k1WuVZnrNDa37gYZ3AYO4duVNDyqRzVAHc4HkJ
0TOMlvIhObdKRveAU4Xtx5EhQE8iEFDxLpADl5qGmMVYimaVsb7XPFnrltsVch1v
flgfIoLwaOgcMpG5Js3kzbotVM5R5RhnOLyupRnRZN7k/sHprnl5F4LrZbleE9PI
Te45qk0Dza4z9KrFIsQKZX2+l2fk59kurbXrExUhhEHRlZrFXELNefPTqZSS/IdF
1AOatK49R+UMgeiGrgLeV6GhrHJKIgBjFPDfQ9xREbb2PE8bNgUZXDZIRVfv6q/u
oH4uX2q7eMAuX2aMjtLBlexP+yTygWck9Uh4sxv4FnR7qWiD020xVdCshUZxi2ZV
F5WngktSymVMfpzlXrGwt+CYJHDwtRntTMtKfo+ycJDxCcYlhK1ExixTmqsyS0ay
9ss06YBxFCcScKtfDF+Ig8BlNc+ms05PPMZWUIbYCa/6kOeqHQOk738Xn0Fa3OYj
tOnUoYifvkML6hYQkoRtjlFDxo/j8972+DQK+yt1aVmm9Z6yUDW0ewDRTleINt87
O37kzwnIK2tSoakJ2y8xtjP3sE0hTaMr3NUIJlvwDNC8MIA+ki8nd2N+VOueiS3e
biX9XJg7qT/eZhQMrNkLiDqGpSDrKWjTp5jrJw+LfO0Z14OTXBkA4v1qWt84fiY6
/h0xZwqqrPqCbAU1zPQjT2bgX32eEgwALERuRzacUbwf9kw2YT/LstSOS+SKAGCD
w2rtpQKQQ7HztRdoNdjTYayB5qkfBOL4eIqoR8O5tPlV7HnIl+Uqnxz0UozmleEH
NfW+GhjaZz8bxbFVKxpyHczdqQMGnDird+Wpbss0Z3sudeD+glSi7l4sjN6wm4Ze
MBXNU2tM2SDWa7GH3GmuIEzidPNBV6NnQX3gEfjuqY1psyWyBqWOORi+pL5G95JK
4yuZtR3vAOeAhGX5A9psseQcC7V+o+eCNCjwidM4E30yY6UzFz3gKvLsw8TFROf+
yaeiSpxcT4W1zwmyP4/VX4uZfVWa0Q7a01NKrnGuT47GAs5C1nR8+k9WYplBD18h
cokKTc77btETuQOULV3Yd6r4A1N71O9KTcvzQEWPMTvjrGX4BMLWMyxUY2Zef3c+
4HxIUzkQwYFkMPOB9RhVVqdcTd1xVm4D4HejTru7r9udT+pP5iixZalFKkQIzAig
sM9YRC1QLqNuCLRhBDyMmQHFpIFYm9RBZBTmkTDdznKQkylL2rQ1wZMPjfqggk7a
HnXnEdz46N/Cu1+E3WSDWAdU2daNT6rbamJxeKj6Vgmsj8EVzEKQ6fgsXZNoQRLN
FbSqvRSk1gFY3d70hzeE5QGi1qj3PEq6pL81V9EsJqOpjNS7MZ73JTFeHe3ou+AD
IKi1FhiblZu3bivvuZVlAq5UTvfNxHPKDury7y5awgkFQl2/Xd1lTGwYt6e60PPp
nO4DmC3N1VEgvy0RpAsvP9qvNd7v+RNhV/ZmaF4LPftFA6UQhYbdCrTyEMT5N2TN
4CBgN8xJo1YPxaZgduNOQKVZkuRzWE39IC/qfY8Vm3lTaYoYUaj0XPKxcxqYNy2s
A43csmMmiVZbBw7ivoGDLkA0RN3X+dz/JDTp2iHb9zlKzMSOaTWjzNAgrDjYvBYg
TrVm1pVYTjqDqit3QRrHez5bQCa88N9CAJAjrrO5qmvLRodLnH970qY67Z63D+5W
E8EMrndo52j79EwpQT46cXlas6RlmJaK1y84+7nd+tKL+13bQwR0lnjajHUdG3CP
1ZJ/hXwqFm1WYTUSa6sLVHOZ+RdtQM+LF+MBzaXWC5pZDaX9XTSTBgrpZ7FaPJdT
MJqP/4FYZ+TBoPlVF3jCDs059UXE+cUYOhN0Ii91p4yGh3VTrOiMopOJdJjIiCdP
By4c5svMMz+c7RR23wmdoMvK6XqM0zPdW1F2y+bwbamWEy1Wgwl31iHopgOHVZmj
qpz0Ealbgn90w2gieSwnk7oDE87Rg9nd2cn3GpxXolGvPgFtonX6ZrK201GcJqrn
5sN1u0KKke+qRophczJxCw==
`protect END_PROTECTED
