`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogDU41aPwWtppMuP+hWBmtLRSX60uHGzWgr10f/cYCds7freDXJQOEdaULJ1PFMO
tS9lLTmHpjQo7jBAsZaYRm1Vx1VFUMENHndMeJbFjASoP09CGjrjrwmN+WC/cRNY
DjfWy9UfXtZRx+lunAezAE9BwAQ+ABtQA964d+/wbLoxuRPtx1zRnUxXu1qMmqPI
BvcDrGrSOO0OIKOYBVG+EqsQjTuAZYeZSLb6sxMUH/pSpPrRMEBkR6hjRwrd8yCk
7/Gc+2gnBbDdab6cg046VyHwv2OFs66ntGuu3ozVRFlZlgJKoLZnhwBmFUlWAsOp
h/cZSZJwJyxI6Zk5Faoijv4lUyrgE73LMmVRrveb45KH7wSYME/GBFRMSPauSUzk
9gl+K9OBPbzQwQxEgOmwUjNyzSfsaA48ORgcdGdGMS6GCnbOM8wKe9xIAW4sLRtX
T7cetM/JLhKpwZngTEY4ITQ+vdC962StpEdKMDATpeY=
`protect END_PROTECTED
