`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xj6Dxi7w/NPS4VjuCMJtyHixwPUVT4mUwNb6VqpzGtLmNSLnNQ0ibAThTNl7LAwn
CSH54tVehRn0Gp1V0a6kz8czayBTfBtSBgM7WxrS+L9Ag2MozUA0t4IYoTn8nuRt
mKZbjNXFoHvusRDlVd4mXjhrnD4CG2eqI1MnVK/ntR4AbiNc5T4YVlhcTt4SrfOZ
O/c0/EVZxjziaycue/OiY18PF3lhNZRBP8T6qMAaF4MEw4zr4AsuUPp2eVFowkZK
MRUt9gJKg5kbvsWVtJtKV2DF3+2YOt5dh691uGEEp201yBpijrlm/qC8BzNobvay
u8vHDsysREG2rP+fWxviZLXAAcUYXKG3DVJl91BjoQ7ZW7KFIUSG314BDrR+ap7C
YkFNcXqqtctylB+fhEs0KiLGwudiQSlTpg4cY0YEpOBQPtXQpsDvT4YnxyG4ilza
hS7bWKQSZOy6Cnd0NsU2FBKgaNwi7fkS7DGIM+AlsoHkoFaMXnZrsrnGZlbXIlcS
i1ytGdoj03IxgV+wVMIRtkdfpOQz+A9R0fRiQZWZupvz9lGsWfRRgdaX8a2QC4iZ
IH0FkJwp2S5+LOvv8IpV5tOFR/G98/uw9wuNa/D0bVo2PUto3iBjbOuR5IBllESv
4PTxf5eg1uoDQlDsHBc8imapSfGUFkGXR4TKmGf+wFRg4SnqjLZWi54OXOw1WdFv
QxPIWZSLre7MkbxBnXT1tvHssarMR/CQWT8N8ZtTuLgFhDwBHqC5pTJkzL24UMFd
Q2O4gqm5IMqWyzRO9/ikYS56ukzBMcutL/VQADsu1BhdEFcvyZs1Uk2SkBHjBIlM
HZXI9efEUEQmMCe9hhdJGT5B0f90atNf37xD4jbZvnhyo3xqOi/2I2Q+mR4+7rQf
XjqncYSk1hQe6n+GmEn57tCdHzSyWvfpaV+mG5keQ9FuJdyoGZ3An7nszfuzhhK2
sHRf/3UjQvPio5de/+nNvmUw87phArQ2ZrlGVutGfvtLRF5zGu0V0TiiOelY/qN5
AZER+xYVrDYTNbFjivQhh069hmqGPQdk8thZgZmSBUL2ExNLHDhtxIGtVvtph+yG
W+6q9tgdTSot5ySwEFqWmK+Y1F/TCSeXBz8s/mHIKWeJ3/IgqljLxDlJPnZ4qrgk
`protect END_PROTECTED
