`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dihgVa6SAFGUqWFS6TCjp67DtJ66AfrSF1sRI1G8y71KE/ZYjW4yps14dz0axbaA
/UuX+rD7NSP7JcKVmybAUIQ0uOhMDzsu93H49O7ryTI3g0rKm8WWpjJ27Kuqvrz6
iv+B8jtcD8qJDzJckfLoH5egFfe910FL801rhmhbNcd2FQtKUZJcCYNlQyoUuavc
e046td+TvAF5ho5UZpPQsdADHyKoB/V2CVlcLJ3/kRY8CzaP1N5nKEXrDJw8t0Y0
nsG+CWWHqIwQjZJfEwFuRhdX2VmCCbYD0f0qT0/BEmEaXdkKt3RaCl8eLSB7iWzw
5ZbvZyRt620gvfwOeaBOLUDZ2g1LGK9VvPKCjFWMbBZjJslWMs2+qZ5z8/pJ+BV8
T209UcUi7xgeHKtlkIAuSxyBsZMWe8Mk5ClyMFiKKRIODP3wLLHZTy/HgiQIjklF
t/pVce2hNNUlhjyOBHfOOXYs/kRRE61dR5B3/x2/FkevJKZ9cRDc4yHOawoTOr8A
MeFgGRQg9uBdq+S2hCzVzLM2Z4hcVVnkjjy0x1GbgoGBXtO59AGUwv/wGvB4QgJt
bnlai9dZfyAS2Oc5p8UCbWSKs3teCLAXOuAQjjjPJDhYm/haiWCkRbNhZYPrQxVG
IN39BwERNlMSIM3BG0S+DUVvvCFYL2l3osFJYQtXbpHVplXXHQAK7mDkAh9K+JYQ
cyzVksItFuCZLhC9D3QhSA==
`protect END_PROTECTED
