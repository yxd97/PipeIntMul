`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99l4WZOmUj7h3qYEDNuesGVc3007x7qrl3JSzxIpnmr7uRjSln/X3I8UXkZgLQpA
QnrmB/ONXYGGyS6I8KKCdUyVLQnzeGb4vHj4r3gFZ6bpYGvMH3OXBDPUmGiBkBUP
Dab8rg7uMSdivdCvQ1pzUlprGyTgtDgIORtm4S+xFni1/MMWOGSAekuwH2C6hoVC
VYWgzu9ylCLnmWJsL+H+Y5lCKett7LoKOZ5j8g0bQwpwl6UWpls5USBzjIAlQuSg
SFM8JURAhBN1ul671Z07BBK2oRe7BdA3krtll9Y24NdfScJ3QhcE72gdwxLndqZZ
JjcwaMddDt5u9eJA9oRPREKBxk84HE3X6Zga2d/lzZin3ba/h4qzvm6hbGtbdGgq
`protect END_PROTECTED
