`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ubqcUt74BqYG51XfhArcAVz7QdTJilSV4ELSgLBfoY9oumU92HYl4nr6xLA0SMK
cDRBnDQbBISu1q6NGehOjBzUph8fElcHlkCM/LG8RBmpaz200Q2XxS9CujKnuB8d
yVtUfSIPmaADykIDWPpbCzgS4TswCe+UChA/gYY990r1rV2b7kYjRpQEbv66Fb/d
v3cLWhgjzWf5IdVAgLnXQPwtI1igRtnewPDoxb0Ng04gYT74B2LuAfDyp02ynvzs
PebMTx+joH6fCHaVXlA0qIkn9y7J6gM0/OXhL4TS4KAwpmGj4u5eUw7zLAb4Gt9/
DHJRTJ0iYw8+M4OQpmfyBCtwOAfqY1HOUw0rnjpV0LJhqGZACpR+/hue82WF1L0E
88U7GJNyp6bkNY8wx8CO0WlJ5BZYfmigCLQJNbJWdp3PztBsn0/uZMkNYS92grbY
CjSkmF+Ns7XHwN1UUCFZlpSGSkIHhlhPchVwPOvt+6l/gdonRRn5AZwUDKCsF17p
6bQGUJUF4iZoUFr+GiTKTTv4sPRbsj9UbBPJH7WD/JDd1suRzFt8S4q9lEyK8VEb
GpPhzgn1tAghlYH6gE075aAn7SwkKuxbeSMQCSVZ6EWyO60ERaT9kuaCVEieEQzB
u+p+FkI1dQxkfv28ZrNMFKDLB1PgkITzNL3f1HGd3RzyKcNoOorQZU/KuPx/8K/t
JQSNY+8dgRQEKlMf2aSyXgg2EIa5GFal5meaEYcl+OiMCyNsW12BGIh8eNZ5C5Fg
uqyR9LNxV8xfhdlnZMr1U/v8uMKHkeZDsFSEOFEk1lJaMCwBR37E214tD0VIV/ar
rMBFjQA7SKQxbM2blhWH0Sq3zvNXoM9PpOFs0lipO9lr10RghQQg09N0vjofMM45
k347BDCMuRio0T3bpuJ/2IxmUq0xt7EkyQjBkey+3EGwcsuZ4AG8gNtavR3kUACu
r8OxK18MagChzudt69RbO2x2U/Z+loD15IX1fNbYZS9hAIy12xwfearAKs/f22JQ
4hruW8A84zh8LrBDT51tpM8wL3ZRllSQhYROykRBd3CTyQlScJg0sPzr/CyLT92s
UNINibx8gMcJ/PBycKNlz2Gz9Rmwz/tpcZcZBmb7BnvyVEfGFN8l2lu+WagEHyCw
aFlFg93k7JDMirgBFZWIdW1/leKup1/CA6GpwyCR+9pPV2Jy9WqIIXoHz2rTq0OH
htZpHAug6BkdZ6AmL/MW/6FEg7wXpQJtqZUwwGYJA1GHPmCk03JRsrENH+GH2jQf
sfcx82tNH7RuHbO+g7uXGVb+xft9qRoYJ+i/0LC18AKQ4jpmlB/9AnyEgQ7e3pvM
9NPNEMdNvYdtmf9ElskX6ulONnZL1+yUo3iXmkeJkImcM5rZWDKerZQPOdh8/viI
`protect END_PROTECTED
