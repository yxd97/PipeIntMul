`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ULBMkBLj9Gd/92lVVE9gKtZ1yQVHP+eusbq+n5su0nLtN8Y/wFjrUGeklb0hAB4x
psKXhfJsM8K2l5bTHTCcS3Q6W/gP2xhwpdh4s/gJYvc92SEfCjNcnxfDMAcDhcSU
OlQtAYjY434aJKAhx1m+DHOSgKFoT9OHvTEwaLMubniYdPKvrbJYXMxNzWgGaxoh
uDthHEaPCa3rFVNKxUxT5eQIuV1GyO7TERkxBEKYc427nWURqFPIvTopV7g79PrE
RYBRcCgTTnOYfaNhTTjQE+MqvJnXItXLfNlOhvCTol5Lzn02hBjuuvuoUddpMBTx
87Q8bJUv/F/Uv8ZyLxD6XgOkXNV5U8YwG+jezXd3GYlailWZHlAcemjSsWcME1nW
LJHLOU8ODCywwV92+aFUshebsWUoOF0W4TT6yZ3XSjzT3LC4nxk21PlifjS9ZPtO
3+LvTeFwjZXirdRfdT3MpUTfSXNTHXbrqUiPNJe4foQlwBsr4Zd581vqL/hFuTGB
oN/oQOGsVMT7kkmUg5DZdVTSzU3petkuT9ANuQRaVzY+6XXLXupMcNCn3OcWOU62
/9Z4DknK9ODOliJZuq1STA==
`protect END_PROTECTED
