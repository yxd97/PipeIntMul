`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8p0tcz62WaY0HlHWHR1EETmGtLQ5NBCWvJa7J8QOBbJCSBReA/ACDaeQQ2TQv2LT
m/85Y9pCQ2ydLwQ2PIz2Xhe6euD0IN5AH2mzsemF/7fwD6R5XLpDqMDBPrauw3uF
AgWwoLT9Q/WB7AMj/q7Yis44817UBSV6HZ7mUCOL4R08muN8qRTCX6wzWHrpSlHV
sVNYO6Xtc5btQ1e3jbvExhmV8Vt87gzFThIkP4+iV8HEjl46YlMjpvXu+R0bza6h
yu6yhbNOHdQDWnC8FhEtUn/bFtH9vgN3fdV77w0hPP0KXLFg6MTwgJ+7w8xICnUM
`protect END_PROTECTED
