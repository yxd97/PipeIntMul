`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YP84npMUDGiLhzcCp1NujlPD1RXbWwJmBreFkR6TXwi/pR+ONGaOkt09ULyPMtDY
F92NoxqHn1pUbdPXyzp6NUZusw09NPdM8GO9r1V9hpFgJ0/IO0szIr0FKH/6yWps
dlSFyTS0r1KDzyOVpDb4ZLIxeUt+h7YOMgHpqn99aLmhNoQFJ7DJ56dp1D5+fJB+
548lRguyOhjMEcUg8RFH3eVk4R+DbLqS+VXRFRjNhldFBfxjw6lJa5lICKdTnFWj
3/VjJgsheymWLd8XkKfWIC17ZywjYEuxa0NDjwCQetcuaJt2PknXzR7mHqiIdffZ
KXfBoip9MqyVWPZQB2UsjbbYdN6mlZEQETzCM8XS90GNAP+2BCewz13LqPRoN5ML
zgUJu3amSp3LH2/KkQVw3nF8AObwRTl2UHsb/wDpQRxrlnvDhCJMYUYLjpd+lZOM
DMXbMZy8uXiYnqguQqsYqJsyy9nkQysH/MvgJB3ETqb6VvS7R9CT1xHsMtQ1nPFR
wnZzi4NpRyReXK8o5CprJ4NRWcQ1Yd06k1ujUUtFasbRm1iJgUCT355fnyiBsrXX
TOdrLmnHqW4FIV/rSbI5qtEtEMC+p8aWcq0edV6VMsd0r0te0aLi/RroICaKW88T
rTnHPjLhYo7CBUIYwFdUKnwjFuiMEwVFOtH3ylBLf596mwlD58amJ63+lzlUZiL3
bkl178TmPhK0gmJFn0IAeYBq6MZ4eR1/sTfZN1XQgYSEkUv1m5LJfpczywGY9Qvj
aTEiFyOgqzd59sg7sCI1ZrhYivI7u+6InMEB+5qtJ/6ysLaEbXjcRQv64kXCA+/y
8IgW5rZrzPh/8b92BpTavS549OvzlmEkp35YELrBnjUaih9SuYq5w9Ov8lsrYHSy
9iw4kKEAw6UCh5Cu1HPSH37Oy6cMi27UlbKimJ9wS6fn+Nr7JimjMG8Ta0896ZwO
`protect END_PROTECTED
