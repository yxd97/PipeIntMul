`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SA5AU8mfZK6QaFU4DcIqQ8mtOLAIrEWLjoLdxcfn/FkT8ErpB+MnXvbmHQ6/GJxV
OG6yik3aDwM9hBdyqvFmaZVUz9I0CCjsnsdptxIv4RPCn5MU578VAE8vxIwRejMR
0sxABcizOP2VlhcB8x8zmuD2ejBgaUB2zyjEaPPTTfjc5pmUrtw5DFf15v6u0DF3
mdGBn32i4PbAJ4GYO82YSoiWyCag5PM8VtHWQqcpHw6pQzhy62dhqMH8bqMd0isd
ibOVOqdo2aKpjL0o0x8qMMpo3MosVrTmqpLClcUkjo7XZ+ZZs/TdBGPvmE6oNGTF
N2IPR0L2WhcheqmdvcfirpBX/BX/b0VjVI5E7iztHRhO2FQ91srXH2EIAD3R36Mc
PR+C1dCTV6JyLLsBkq8GkOKpv9QiUBMmm9pt3GpFykcNkGdm2Z79m+bKhsM+3IyR
vat+Gr9bapJX1l625S2J+aZqBAZB94nVDtKWFddEM9fE5i91YUyEhFObixdJATe/
ympY5QXgENRXmwSGJwhvborOvEAQ5JXh+2qC/i/UUUhn3W5CLM8vgNrFTIkZ4kD4
eXlsYAohMdMPUzgeoJq2uQLg7Z2nBVUE6aSLVdAfSHmzZ23btQhlJ5IvMyRn9V7a
ku9vHgaVnjUBFaLj3DUp6g8bNIfW3M1U89hUfx2xMqyIkYpEGemXDfXVsPFsZlMy
/BZqkjBAHi0+/DCSjFKYeCChDljOuemb+oMkO6Nm+qIzXGiMwiAxMvQzp5neOgYr
5VSHjNFhf4kFGjeprOXOdN9TJGpG1haJ8yP+Nz2em7R0nr8VGIaA08MpYdJqF0U9
2MVew31PY99HIEOQH2Q7KBRAvmEUHhezz9zkSyMRtaqLXouhVVXPZfItb9BRQE3S
tJegcbMNQFW8Y+n57WNzQRO67yX5YNFVUHoKOykC8tdDRf45BoPYcFVvm3kio3/u
I8g5RJPuKuT2f1rnuiD/lwNj4GLHrfBy0gF/RA9+Mg3nfQA+I6Lep1HzgMhTJXDp
Td+O084D3Pc7Qvw29RijK+t/peKGoAWvvbCme3tcV/7T3piDCDiBHf27BhI7A2cd
MrxxmZPCn/asNqbLWMTAGgUD/jKkYRp6Ub0zC2sSwTaMHDV4oigVERjSc8+m510S
0l2EuDfoWOdrwijJgP3wonCKxsz8E3xm31L9w4u3vdR6EVLZBQUSDoZ+Eq9Snm0f
9q+npNXQkA5HsR7fk4+1jCIAlmTJ7z8xuOTpYDf4KUmQfs8aDnZ1OPSuyjyCuvgk
tYnuAvdQKqw7Sz9lMUNgGt+xUXk/4GNB1XEJZR+n4k33qYuhyX7PqDKhf8ljVni0
cVS01e194W/7VmfKyI9U9NefZwHp7vs5aY4IB4JCDisB6dWFsvAY1X9L33zyGfK6
UnN7s2UIkCT1ww7AIg5zgMY+RPNtl/4f4cF3zbPpziLpe6FGX3kcDsGAJDfyvg3i
9783MTBRDRhfVs+ABT7WnaXYBu06phn1MXBA9jDu00oSBdPHxJYTm5qCoJ3NbOvB
959NoEX1InF48Qf/baYndKVLDfdHl+qYFkxXkQwWyssp54XT7pmw3tJ641pCt7b5
FhZp/H86DN2JWrS5hUdiX3L5RUxQm7XLF55qX9Wq08+rYupHSSfyTn0oaRMDgQai
h9UZeroKUEBHcMpzgppmwyRHdbI00rVLgDlG0lAmzcqpTinGZql6b1K1J4+qBBHk
Kc0cYOiTbYnvqhr9+NGCHRsTpBasbJBIVqkCxbh56gIT/5iOkcuciIEw+J2MJl+W
udRQSlzEfNwUN96TE+8ICwzQZr3iDT3F0qfBs1ojqiclOHGV7+o1+JWK8g0vPSCY
NknwAEhDtGYTZLGA/X3k0Vq5/Ha/yy3x0QSRHG9vLTyNjB1Sg8XI4nElXoIGerJn
ytNKE++yGWU/h6PU+Tp4cJsZKnDbBqe/6HW8h0M/G1e3ZnTHxVyjL9ev7gd9qDW6
xKTG6z2dPtTmM4Bp0VGQsKcrxO+88CsX9vXXO2TMTEX9CJmcoleL7jX1DZg2u0yB
xvZKI3o375NrDe03cxJJFM+N4LWfvMO261lTBGOGXxTXVDkQJ5WMVUbthyvo12Mj
oWpdThl2Cx2upaDcLpLZtygLMfVdGdX/6mfzy1CpRO75Sy9EPpRo9A9HYEJow8+u
EvA5X5eR5LjJLAmE7KqWk+pj0/acTp9+8dcf916EW8bPyOBrc2YaNBjEBEHYM1Gf
fdU2im1MlveQfK+h4j4o/zhXUBFvHJeJ0oLsw/a2m+9juMSqV5jDG+eSiuZ4qRmm
Z3/KAx1pKJZLbv4ezvWjWdDDXDhsQyuE/eOwZPznn7kbc32MIHoEkm7PdbyrIHBm
tWsaO2jorLF46R975FgTSDa/2M+niKtTu/B6Nai0zcFcH40IpuHFTxoLTIIWxQqI
HgpUDU73dMFmVqgWbqdBnCN6tyhuqh2ZHdiJ29iRZ+nVn6sX0arHMKEKtZV+hSCI
hz87BU2qwmogFLrrpnuaHl1UwdRJJeUFq5AHvurIkTRny/+1AY7fYkwFyHD0UPBE
purequuoNTOskUFXSvviXEJ0ndC//DDgI5hX4OTEPUCr7kaH3qgGCgpgymDLAZ6j
0IzKGbp75p3odAccQLKgFXCt4WIm1PKGDMP13ggco6PihoxVtysRogZaiUnF7Bwt
aSOXa9fsyJDKCMKWXzQEzA1fbunDw0KtrSaZ9zUb3mNTiDyapDdraqG3i1x+joH0
6t2j/EZpY8cwWzYGefEoBK/5pgp6byopxFnXv3JcMwzlfW0HfMS42dZrXtBG+vJI
8uOQT/gpZzjLsY/lcvDYAhIpP9gwq0QltBskH6icV0lvw8nr+ZdBJAdbPdZCvsFB
XiF1jp4cQ9TqXj7LzfYT9FKz+SZqJLcnCOs4KXA2mLP4jb4jGC6+i+dFBYiD9ZGM
lz3/388OEbf/2wjh8tg2cbFhlNM6b/fHiXo0iFQ9jZOcuTHmoH/d+ClkalCbvza1
hfRbooPTzddbhLjvrUo8DqfzrvzF/5i3+B1c0d02E6sPTqgjzASWVo84ccNtFM7N
Ctf98b8csOJJrKhgc2m0VmdCjM9DA0btbDlgKI+vAUXUhWj+IGwD71CoYNrbIRbY
`protect END_PROTECTED
