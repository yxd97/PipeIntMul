`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLrEE28FT+jA93FCD7/arxEEDSc/XBGVaZjD+CD7Wt/OGjav7nllNPjmzYi1w9JJ
NmaWwEwq0Y925nbQy0NXofmbwzBUSwuyMyoK1mA9f6h9z0cNwv/OZEhG9g0aIXAf
nxOJJVLLtm2WRqCkUhC/cpjLp5IaNC3z1uPLGbRmSIQLbCa864kSAJjuFPV81wBe
1geueKLPvEKA2xVRlybu6jkO4csqKgZL0HE0ivkn7w2mxMLgY1ppfcZEZHfD/EVd
FP4ltM22KwA8jJSwvNNj3Wc+bk0tgbAd92iTY+YvWJt5WreNU5GdT0/RCU7R3jtk
PQtYn1MDTIOHXG4bXCNYfljq2ZtwQTuil3VDl1V5QF1mlG+68ZinJa88eEn0FlHg
tRr80eGvtB8YHXsR67GoJwbepaZYGUlURIs+/GTZFkiNzBbPrH/fsfIRoR4/UTrs
Z2KBhCfWQoDhzIdX0v9i6SKFUsCadLAuG0hnNRrnWYSYfxCLnPDgkVfArJ3ZX58w
TrIK941pQ8jmcNUZvW97P5NDXB4rYIv0QXMBrsskEUa2AevX0qvIraY9GsHtMgHM
b2PZLeFJeVv+XtJu15zB+oRkbKBzxqpfwQbspv0/2ioEoml54vu4fy5/0MIpvR5L
MpwmQXgTQ2ZItHkf4Kj4SypBnfU3MHbfuW4lB9s5/uDR8WZ2cReHUyh8XvIrSgZM
LDPmOc2/nEIhYIVUQoylvFjyvjtNlnq3OBTmk3JDRmLPj93EkRrOfAn5+xPzzOn9
+he+ysehpFB3/Bhd/RFOo+orDVLcstUvCU1pKdCFevVPhoIZ/qE3oGIPS7aTtn6G
XfnMM28KpmrPEAaUq27Se4Sez35moRNa45xA1SqOqa0BDmFiksGH58JBB8KI+woR
hNKP8GJ2PDNlaj/5oN0D3gr5EySlvZQDWwK7oONMlRKyJBr38j4uOT+kr+oFAkE0
BomyOvuc7l2R9hyh4McsLDFN21+8hyOXTquFBPmvJpwvPCd3eFUntLi0OyyImBqK
BEKnU5y8QcBUOK2PRUyf6xYuEWC4cdpcxiHOobisc9PvEsubPvXRnihPWuxVQeAi
HxRkBpFAPXG+cKqoXlLGO9zr2zp25AYIWUtvXl4vYxBPZYvVo7MVj3S8axNJ+cr3
jw+J6KmsxMzBeRN5TKJ0YZgV+jOgfWQYgREiluEUAYWkUjEy8JPJDqWBZhEUEmPx
SDrBDw5dDS86OcxE9gP6qOfYmckJ33oJw7/vPwEvTD3nx3L0g+uLBO+eiTu026bb
e0QS5DX+Ty+8/72/BNVjChrRlTLwYn3Oz9hOcibUVfWldfm3ZuTz2XG1+nrUWiE5
PQvxnS8AYWAkQcVAX78d+Z/tRcMm5HW+4Z5c39sP/vX+Ci6uMX6avTA40Tpt2Ab6
meaJl4uTK2cd42QBUtD5eGjeoz3sbRKEPYNljt/3W9muikovsC0UYjIJKkSwMoNr
x/qmUZC1GoemYJc4kuY/OLCwopmrzIfL9kpS2pkoX3aTywhO/+ejW24eaUs+rARj
FhTwH5MPVzbdnmEM9R0qkNE4R0QBcyh82jrpAqrrG7ooR/Y54+k2kOC9dfxdnNlf
4jO0Z+IBBNUNzXPjUVxyye9QoXPw5cqqorXvnI10zs69VQkNYq8eD+tZfZWTV4TD
U0xFcM7kx35oKIQfo++Lp8kFzjI7I/Mo8WRgRs0LtmvqcJ/4SUAnBg9JJXDVu4/L
ATT9xRYz4X5vgjc+R78tM08hAkRYe8Jfd+KooG+HYe4t/DR35oQ7LYuBB4u12MFo
rv6Ph/qs8TA/Cg0FcnBWAVRLV83B2pNsy4GmulZYwzgsCHRKQ3wIypuxSZHm0BYw
aPwlHKmOJRnxhVQ9E2HlnzYr8bBysIBpfWS0a7weWi1txjjKG5ooNtjoqsC5dj+x
SB6D/G7OJ7aa1TNPYENyaD4YWxezKo2OYtY/9+N9ex4aNuF70d9pvLIBj55JZEA7
SQeSv/FnAPKPwITGZIJU7S0st6X0H6+M4GFc4fk65HOiXe5bM/ZM/7aBJq/h3Eax
Tjtu/Gp8pGTVmZEe9m4c8g4UCrccJ/8UAcqD+JCspvjjRDPJ5o72SqJl041xpBmN
Ax/QA0/EPos88Slsb8we6n7BsIZo6Fww1G8uyV5FFFBrbHOsYr7ORFcxPEyKZRs/
I3+MUES9G2AW54PdrMu1ee0Y2rfUFPRIRhXxWWBeW21K1uXp0byHesZWV3/8dwCV
+7VwR4p2ipa5IiAwtotKYPV1GExfuP7Q1uxeT5b0SlgB1wbr15FhOWCM2pjDKkvo
CxApaLOJVwOMb4saFPubIG0fLle/ZkbnyDt59btOjpE4wSMEIiOcCxkaw9Pr+yOX
11qxWE9ZoX/naIjsuMk/hrxM1MUZc26fC5Zbc9mwGbMs2WGQZNM1fGrIYevaXhrj
4161w16nGz4e1SmwNygn9+td7Ev4VDaLaO7gH8nL7ncx2OJLgx/t6Q39N8um7ejT
KiqzqwP2GBwegN2+JsgwFRWUqZxPNzW6GrwdzuOQfREw1Z+S9+G7xN05La7pc3Lk
yuTzKhDkkH2+5MT6GufdWCx/i0x95cxVO7+yHs/3foPEk0594Qafkl/hzcdW6lYB
QJi3B74G9t1S5Uwx+BN9qQ4mDoeJWi0kBcwGh6dyi3tGEEwHSqZ0FqFewLFuZcTe
CTFSi/5x1IMxx3991+Xc/93ADQH24zaELDIOpgKF2sef6a/VyVYU6fYlfEWLJTX4
TA4fmzxzyx5ZOnQukU5E8xHrfuEjTIsq0ltW3R8PI782/0ZUKav0/sGyUx3AoB8k
nonzTKNZCpQYVfzwKppfVPZ1tJIKhEWhTja1Pjl1nzCl8jT46dkdLlK+08LpDU7g
1LAvlhSs0jsNO4hCSVLgQtiX14GLIYWNaKlxD5jYdvEW73pcVWNjCpPJMwMfP8wL
S9pRDvNgpykSu9jvu+52fAke+lU3tdzvPXumqkPhLl8Qm8wHNFq7992WuYe7unDh
4fFwa3jefYVKPkg5HUDGqVfjqGubBNSKhzm6h/fIo0JG9X8KAcqJfCUR+XLkzu+e
gLjsApQsI3BZh7db+bB2WV+3/lySzNRCoACU8EYjjr5aVtlN9Rzjgid9Dy3MPIP9
QK7N2JXP3LAkZhhsgFjQhZ3PJfzdHBxnDA+bTGsm3ulPZN7NILDY0plO34NKVG7C
cHmQ2X0a/VqpbmNPjjpv76LogM4J84tX2STJOKohsItkMM0FMSd4g0PM7Jb8+vM1
POY2qCak7+7fE6LTJzwkUAVsSaxVmt2FNpGDcgKAbTmP9JYbtqHdqtUGIXIFtqc0
uB1RduBDRwkZTArsAfWDAwbInwzntncigsgQkbl9hcHpXfQ95tUtUFwUDquDnttL
zCEDwGjzHOSvy8QiUKsL5EQMbLKCt0RwaSG37tD5rVkVErGeKZHgVLdRQLYpPq2/
XhVNCLR6b/XaiAABX88Rc6d+udt3yj2XSB8HjqXUMPdLB2kuxe3Zj3oZWCtiSYzE
Rx6qyTAuS78q/FLLhvnOHSh51qcu51YFqK2eDPtzhPkqHwLIDfbiCVyKNlRE1cox
pc0871K02o1avon0S9a6noscvNiCXe2CWfGnS+OewGtQIIPSIR/2IbBBBJPVerTE
gdZJTP6JRzumouGLccwEGIZszcdHzu8vD+jVtcH0nbNeBfaDZXBQVT/4lJUeLUdp
L8F+5vA3F2Cs23JU32G/zJhBqZsEwQldTNYmVG7Y/n0=
`protect END_PROTECTED
