`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJE9dhZllyXJkVYhMSTTJBPMdCc4Ts4nKZ9Ii61WMkBqned6SAySFUiM51s33Lai
uqqUpPoGg8NS3VtasA1y3gPKeBdAOQlp+hq/CgtvBYUcsU84xefXX5dF+PNafh8B
+SESFDi9bWHPP+ScMLOJjHdaAt5kusiXcRQFq5aclA/xb0sNeHYkcr6saz5gLCHM
SXb6bnbrQ5AyjMmuk6AjwCEv5a3q+TI3HEeaq2XAHpxsVIgdMTTLzMSZ/yuC7JHv
SH3qTgvSW4X+YRPbWpgIUYsowIsTckhXGpKZSsD6EOeutRp1DI8oEaNExIdoDkKu
tmMVjb/FBYrbxiZXH+e22Y2H8IhtAnMkMxtprD5ZTBE2+/hpqP/+Sln73TSxlD+j
JGX9Pcsw6Y4c0I08Rx6gqv0nP3wRzILvCoKK/+bpaYJaevoOz8sgu7XHu2A5Rjri
vtaKgJCb67HJE55cYGgGTcNCQTtYmdMhZGUzAxjtFCrxgk84O3MqhbtzeyofJoKO
DhxVYbdKeau3aNZTGG89eVUKkuCa0OPn8hCX4yh7T2P35jUWZfqSEhz4bEMUXzBW
bYzg5i33Fd/MNQ7L3FAsnQ==
`protect END_PROTECTED
