`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RyBo1agaMZK52Hk7BnH8KvCMg2MCpIliBHw9Zw9+o83mCwy8WSvYi/jTqc5iZJkE
3j/ezMqlQMzDxCRJYfdsJk8dYvPhi2wwCQOXQTaQLkfwMaJAOyZ9VXsMmHof2Aqc
dYv+/8SVx1SSiP/sktB0Qr0bM5MVk/SVVPQczQw69k8oRz537QLV0J8H/Xn62n1e
C27+fehGCzK2YwDiPMixHfDkG/Kbf3kbXUzIAStAe0N8znM0qvU5XW8CeINIZzGj
GzosenxMVRBL7GQNTAT7+EIYWj3A2V/RROBQCQa0rGo3J3jwDy35bomUov6NWt5n
6dLIlOtiM6LQcBpFeUnzqoBQ1BnsworYA/1sOIJwYdQEG+ATdCEQ/VPJnemHLOH1
ECo9GJcdDpMn8bBYg7gnqmFV+aHtp12Iq4NPSoVeauS0OcM7TBcsEB515+oiDpXa
`protect END_PROTECTED
