`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJboDmHSFSwWi0oTfeI3kptN7X/qHq1eKKy6EfT1sTRcmdcLWOWDlbp0O3+B6u1J
PvrM58lebmnY0RYxlXRmrsBoW4y6E2xlod16tiddTs5/dFGMyqxYdpDqVoFjgdv7
2Ov/PT7BwA3sa45zg0T6Npd5nH0bpep9W2vjl7ya4aBXSTociVGkBbDR6i0ny/dg
4TeTOwTIHxGvmKBUqqHxWPWg54Ee5eGSuMP+Ww6iQ3gj49e+0zL90eezNAYlMKCl
4W72fouYHLwOfoR+e4JtQbTXcEexjl9cSGdluKi8lC9O5GufQvhiBs+r5Rufh1VT
3KXMSiZdATAoF7H2nqZ5E956pzcpUrDmpp2y1PMEr3QxQ7wBEZF+hzGJteBQo2xz
by4QQ+hotSI2T/qiCbpMSxLmNu0GYFXevmf+jlBbMwuAsyc2psruq4a3ybQgSdeA
LgglK+lg50nzhoDVk8g2RA+zpIbUNY8c2L5eFzFISKr/mqIou6KCuHH0H39Itspv
F1UnKlHdD3KQNfL4spSTKkBOngXMTsj2+qsNn42sz3P3BXviOUggxeZDc4CUGre+
RpDhoZrBYe5lY4k+BSm+GZahKZ6NhRoFVpMKfh1L7YqpglTHZ1lBrmqvYS3jnVE+
qjWrHH8KChzd4/llQWIErAbJJIN7UXlzcmPoKwWOuktK3l1+4b/nL8FSi9edH8No
nT+n6kQE7Vo45DopULsTUTx126R70arGOjvncQj7C34bexsKlhQdmg76G0zeXBR/
/wAbaTr2tv/mBBEizkP0/NFO1uQcWmzSZUkCL5fo0mzpNmopNVdSUTYUV/gVf0gb
+LGgPpwruYdbnWjPum3+JrKOzHFt8zJRqnqwQaxlkwrU5QeA444W+5lPdJSCcrx1
35S8uDVTyn99syv3x1hQ3vffQx0ICSTsCpY0b2u7fx5aUXv5PRSU07ZPL16uVVYI
ExB8qXjGWn4nl+HGuhFONcdsMkEAtSn340ix4oOrGr4kPEwAJKdpLU1DZbB4GcI1
9Cp9jL1h4DuFxW3V/w6C7g==
`protect END_PROTECTED
