`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0LiWv4V74uAWaO/DqIvJV/rIYbWebFsVjE3VcCygn01SPwrh9FvQJ8eOcKnLK+O
MGJKAMOgAYOTY7r9jR9WuflMv8Sne6+/V074bBv3HUJeD3tWBsgnk0c0ygYNKFkn
ntH5K/F30afk9xVVG1argiKZYUp24WlyOJtuQCiNb+ImMNO9SUn151rzvpHjAx9g
inHrHcZH+U9Ft01uSIxNlzuAbtmATL7U6jYabLVGpyYTW+5tl7oPrP+WXwAF18L3
85k04d/jlCI3Znbarm0q94BZA0dGJtaTxAqnPPSYgEFt4FSFasvsTCcPrE+iKXu2
wqb4w0I11xZsObp4p6cte4ogX8t0wTiivbXrDGU0E/DGB/FmDPmeVaF6k0vCSSZj
kF05354tNL3h4P2QcW0FQTv3VjP+tqmmTczsMimGoBRqqc/5hh1wtr2DInPCBWLi
KosA7KHCejYnH+IX/EwX6W/FPCD+NNEo9VOB0dedJR2k9GdrqVthrqHqmsfMLVeD
`protect END_PROTECTED
