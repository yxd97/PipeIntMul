`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1NiGIYeCVskUHNGcPw3yTv37jKWIS+XQr8CoCZiJoVwutSNHLcshMiTHKVVmaDk
FtFJEtGdkX9buBZcVdqsALOk5wUo+at0geQ6K3rQ7zAFXAr+/r/zibze36095qzz
NBe3j90VyIn2/+bGRNqFBZqYmNwUmxIjIGh4epr9yxjGj9QYfyyKECWlYaQPC7uv
5EdiSJQSOWDmq/fmfcOHUbgyUQCoONSxw0h1YBVxvGMiyQg4rEtaKBqByfWSEQjV
25mjvBAS8xvODDMmHyUsjllsSCMsVozoM0IEbdwgzsc7bODczaEzCOqI0H8rOZPr
CuJ1+zRxdt+NmqPhyhDRTsviC92ekckdC6PivM4iLXGInyTCyr5aQrhaQzvVyI3H
da71hBeiaVrzr2UY7ChPf4FCyT9b2sSFo4tAbJ+u+HVcKclPxnhIk5NnvObAsUzQ
YMnYQCP5T2rhuOpTTMXTA05AJ2mJqiij15Kw/GreJa9j04VOj/iTXI3XfQsVcOkl
PteztnZWZLJ83cObHBZvFl0mN62Uw22qH1ceBgtkbmqfKDEKpIPfmgKknweFA3Fi
NQFer9QtVC28+yCTgaPWLU8rmbBL6pNLfbWLzZ4NE3bFJ5q1aXMM/IOa2/Wfxs0K
Y03MPQxi+NEb8kDmNoC8WhUm4wW2fTloCq9FpcfNqM60Jr8RAeBi/p+uIemk3Fln
0lM7Pdf91850uVLmi/fiFsOTNRWYCyVfCWe3pz70srkTiZ2DqatsthD61OAw6R9S
kQCa2q829W9Kp0esQUOYHXoVcW4YfeZoCKQfT84zaVnyI/p5LPMtdIZZHVAAIWNp
L8v/1MdmHPQ0OsqNpVXnIqt3y6myhNpoJjbol2J4ZRr6neS0BSyoVLCDWK7WTFmP
NQYHitMPokW7xqcOm4MiydSLJOv91eHXoAzndui56EtJT4AfNpTdzVOuGUgvhPJI
RsMc1MkY2ypRsuP+lbvm8CP/q4tzr67aG9aamY0AJvUECKDR8cXwrqRu7rtybsxr
`protect END_PROTECTED
