`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nw3pEkveXvBA/4a1BNe8Jcw/hT9HrGki6KOd5/pbLcvmd1Dd32wnC3vD3BiVe6vU
v6EWSNAglMQDOZST7jSN4YyBtO9/ocEpyJK9ga8x/yWFlr9OIQpA3EjoWuJBuyY1
UiDuiyH5ILL1TfajicefmE+LGixMBkmTWdhnPzOnfk2zzja0hiD7LKo6gLx208FZ
X4+SiWs8BVtOhL4v675LeEdquW1cs6FSEgdx+1wklTtudQjgtSKd5lBMJSzcPcyM
R3uU5A0I/uURBA+X/HtMYu+bEOnHtnOfnqdHnWZxqe+PG+91rMfM3RF90D5aTtHD
O7FrIWjW47IopTFqYaOfMOEUlrtaGj2CVQUD0qomPnWHf1uKQpBVrOtWfMJzhg7f
FQeDmtm9Pu6vmC6VLGivhJzgPOWnctxHamQtbdRpjPFFB7QPLjbGK4n73lfDp+4G
/B6YGaKr8Fyf7e5r5pLMNYDj3aAGtTtAVvcYvP67zHbt6h8x8Ow83HrX6yS96zp9
RhDyG/DLai10iKj7bzZm496gzRPDN5YDRKa6z5Ib5oeIeHCc5PeIheR4XGP901dO
axxjEDIgaRGfmNfE0s2uls4g5N27+yeQNmHiltPNN9FFF6M5q+eiEaqlFy6RmkOC
u62yxFRx+GP8+NhH0xJAThMLd01rNGOq2uAaojRvQ+9xQXI7e2NBbo4fIod9W3Nq
7RBZ4uViuqw3fPut4aiJtTOLzWbkS/Mjf9dSxSUSOZBI64Xyt/WnYrlM0gD3gnzx
7/z4fxEKRhsi79pRJ+b9vUI+DUKxmR5vbJgTUKi+fWR4cNuMxuqyCL7UzX+MeptC
qjq+Qbnk8t1fJudBZfbNgS8CEsTJils/0ueMlzUkvhIzGvje280/SlFcW/i7+C+t
gkkurqCXN6lseDteVemH8EdkXJsRYbI7I52ZWqDjVp3PyvXZNYdzfbv1ii6kC4cf
6QhKa+EKndUrwMh2X7+T9Uu37399pGPQIGwsdDlemW2dXuPX4TFXsHGOZsmNeHBl
3pM7zZWEUseV8fW23NXQ5UrDZGr8/n9XTkwUKTObtNNvaLAvg+mLQjVQaQmtsqsb
kecuH3o9tdO+xb3zEnDsIPao99ocr+01+TIrN3Zmkfm9kCVlTNyzTq0ISR/h2L9X
aFI83sdSJHvYJS9EsmwXKErKv/HM/YVDQ/x3aBXDAPuXIYCagbPgGfYcwl2D6P+j
PXQ6rpQaY3qKul47UejKnAAzwdrQ4QiPoJ4oauQIcpDSOX9ExRFg7wGNKyG1ArRL
PlbzOR12DXp6yBha1xSfRK0x5GPTK5EDtJkhAW9a2x8ReBNe5Bd4BdRtIQRXeKRK
lqN8NCcn+SmhE8mD8j6BOKpT8xGUyUK0j+iPhcmS0NK1ZWypoC6NWS2wrpe9f2sg
ZBShkxyU2WGIcTTN0dx5/yzDuewjc708TbwFCmaFY9UAc/NMdiFjxFLXJdipu7pD
zsJpBKJbG4sJtBmYVVWaNhUgpG5Y0VPTTF7YWkpOQ223UdmxbDZPcaBwe9qVBPzc
u/ZMm1VWCEHLsf5+XKupx0ckOF3nuyPRshhvjY20Y2bi9TLdkxf9EJW05XutkFrY
1zVAhDtXFg++EjgsRBZltMQvkp0YlC6a9y6HJqtsYEtYWNp3KeV8ZRC5Uzv0SBxn
EJo/xshV5JxHuiKGIYnG3xMF1FLYdEovi6Q8wwOxYwITJTgqfw8I8SACtNZTrXPa
MfYHboHNVbMw56yOAaXPUTmHraO0BEwnJ4zijG1ofG6mys61ea7/yo34PgQDr329
vnrOFlaM0nowtQicrWeyrbFnyU1+pHvMSbw4h2eEB83Sthc6rgu9YGxUrpdQ9CPV
PdKLqGH0Wr/AYMrVf7QJ4yM74VIfBRIfIq1SpSvLobKEBJlxM/GZfjS9cL/KIFIz
3EhVqKrQivTWbNKRC3xHE2uZVp7S/YhGs2T/UYmgkr6RzOc1xXWNcJywd+HGTeFS
dWur2pCcM9tu63je7W+9G1MEbnM0tEwy1g3DOUM0J9j2p5X/Ep7zSuC2tL7lQH6H
bltdRE2BKy+ypNzvEicQhxD8O5QMKGBJGyUJsy5KfXrK3NG7PE6pQpj9FT63n8MN
T7RhoaJoF8KSlRKCJJnfVS4FkCXXwsxXwP7nTY/LtpdT36fcEIVVDfqd3w0DNzEk
C5aofTMUT5V9dvYccF9U69PjO6TNQMpSHWcRosFabGvL1G4Kn15PBGWGKY+r5ok3
LO1JQJ3/BKkFNXYIoFyINikMe4O0SNAPu8QUbupXVJnLM9vSJ2l2b8VaGG+vEj/6
TnxLbeV66BjtW05mQ0veq9DStwSbTnmPTb4oIxiydHuFWIOId0oDnoohJ0gsthB3
GTNsc2h+CFkB7QK/hSLcco+2xpkaDI/EB/M5Wqjki24qu7VCbo5FjEiezkjWziaJ
RMjamqfKXdwfMkcBpC62tErUX4d7MCnfR68F3QDLZTs9B4oCsHQVWKWP0lYVqV6+
ZdoVmk93FawSIlgcjFvcJqD4/Wu9eNet0mcbzvQugTQ=
`protect END_PROTECTED
