`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
amWNinHIeDCE58A3PzFbLoTalq+j9ubwmKZpR2FxR+YPuRr8vAYzeDpXg2uiM/JE
Ppc6gshlxChIvIwiJr4CP0N05dLK076WczHqYurbZc0xLRPJ8UYr44a8xkuKbK/e
cjosgADjiD/1DuQBxG8QWmxNREmVeg7POZGfjipIMuK50HZSH4QX6uNF4aRz65jS
1LzgwSjOWNjgmKDzmrNJDygucjtFLHQPj88heZu2NePjhaykfohzqJ3bZ56Obi8D
mvj4w+aXiKFcenaHGOK+UVNHdP7dV7ZwDDzC9KbAJiVhjnEjH9K2XQ6tIuN4RHpj
ip58oLSsHQlwo788cr5yuaGAzfxeR6DSHt0X548rxEg0uShXuWgK1wFVQew3zPxA
wJRh+sjAogU5Xs+KIbicazeRjcN+H2Ms4S+TsDxQBVtHmrSM+8gJCXDPdd+wJW1H
8stGFGrPHixII7PYKQ37buevoe+23uvAaDQfoqrbsdY=
`protect END_PROTECTED
