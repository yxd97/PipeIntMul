`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m+LXL3t8KHohBdpK0A3hOpNMU8YopnUZ5jybdxUNXRDcIPN98MVe41HCVkufUEcF
GvphYO5lvAF5McU1VoodrsF8m6lZrUyUrNguhaerQa/r9bar/9iZClef1AyUDUZt
pdJx1OjOdp5J0CoVZ3Od/7vo/uFX8Y5k+0SwVAp9Q5AroezEDBJSd+oR2SZnqbJF
B7HMN4aRJmdCJN/iGHwke+INYHqN2V/8W08jktMCl8nlHIcpxZmiv08OiVZARrKW
RwMgEDzBebsVSKbh1QrIBuO2/23RMJydLbkJlaOOodrzyCCl6fuKY9889Bsn1XM1
J+Si8VI/ICGJRXAGdpJWJhjUnc+M8zvkjbcN5MDDozH7yhaMA1QoDRekMwj7mboG
LVJA4MyJXoMYIphMy69tg0J6pgMG113n2iDfAxSNPfIcoDJ4BlPB/yuPzCo6fipc
FZn/AcPupyj76SkagqA1Mn7IIwEsLEP+hd3IS7mQRVP8Joa/okOvRuQT0GWPKQWG
Xozfr/V4t/wts+Rlt6g86Fyf9vLzDLritUki+6t2mNtm8KW3dgb7c7jFEg5FJr5O
hWtvNBHKU4ANwat3ykVY0QPvNZsB99P1D2JQ3kQIgjc38fIRIIwdAZmzFITuFj5v
j7xkbNGwAAG4X8xSYwxDUvla2BGlvdgZHKdy7lqW7yOR4XzYDuWN8cNJuM7Kw1Ee
HIM+HSvneQQVpl1yHAC/mqesbwJ3o8iT4kioiWEZErKWIE2KzUbrhqKGRQaCLOBn
TmRoAHlsTKr8l59t7zqK5lYpLhOCucGGioyu5Rm4zhads1zaDTq6KyTRJbmGCAJF
B3s50k5Gs6j8iwgUxTUbFqw0vpxygcjNasOLgP4Msr7YskIIpTeBjmL8QrNVtxBo
9Ib2Z6i7PDr2ftXLa8ZRnCQpBRLRsijBWBALR+RB4DEJUJsXbQ1Ln2ZfZs6k+NmE
Ee1ZljrxNvrUP5KD9QWJF2lGJRyWFsqBP9dvoN2HrG7qvEILK/vk8J8XxteDyeJm
PAmzUSV9LwVKaQWb7EPhD3Sc8vqc4u3q2NB4tKy/oiNmSSwFp8JB3Td+PrQHGW76
X1TYaf1dBvjzmmyFknfhaT7aW1DjCwQEfBJZIYiHmV7IVnU2EgYRJiwTRQKmfPB6
cel+LWQEw9DGP3HmIyoBpJseiIVgIiR+bb2h7GYMT9IXHpWWWRHfINe/lXT7q7EY
hktRV7Ry1HI+4NFyHHhzL1uJCAGMP3W0GsQS/YJ4gQq06Y74o2NLNxgHV4UHwEnZ
v75N4W0EqYfj5gUfx5Oxn+y3Y/ugCHLo1l8szWKRCT7w3Dm4S7k3+A27bYsHCckZ
pBwISAo/UkBozVf96T0So+YSuAdB9ISr20bdrH5Z6qmpNv7obZ/cz730RuVVC5lQ
1b/ZzVRACU327NzmpYnavoV1ytFnyTk3+W5wL6EuxyfFvJJguLtLJN2FQ+n3n3Sw
mP/ZtYWQnPCydjHgMzOn7KCytAY1PYHT+SA88087oZjTAdSfueiEbXuq03eofVfd
jzem6QJmqbq4tD2zMufdm75eo67/OotR6De9DO2wVIlqIoXH81kZdVLmd9Z/7khp
W4q3u/1xyP/41Mbez5oFmZ3BhRUp0lZ5LBn5qcKrfUSb7n4PHuCk4vdcmZhNFzu9
1AEhSV76Es4nWNJ/usOVoBSulEPAyFUQm1u5PAUZbIJ9/eMDjEm9GVgUf8h0l9Gn
yVk5jJY3fPWmVL3lSkU9rxN+wnaKhzdSG4WpwK53FBwByijUgy8QdpVZLgFUIl/G
FhbwQ5xW/qwItGIoAhs8Ja15j4U2J91IQT4D8Ngk9YWNsKKUpwuOeFHo6SqPb5dO
OSTL5HWBGuV2tf6nrvRog2a0LtiLMS9s30R44e8hi1X6MuBMHE/I02lWdAJHKXmX
mM9ko4Za9urKaveN5Lu1+cBlHM58+2GoDk29YaL7rMdfYVLHyvHOAVXO5PQb0NzT
cU8arHXRX3eaqUl71NUmdUFh2hhqHBsVmZrYAFthij7jUmXqUD90OK2o9st+Iv/+
F/Y0lLN5K3utZEM3iXlDwieptIeTT+Dzm0UfX6IFQE2PlQrwkGHbW2Dgf5dV+irh
zNDIHGoNu70B6eCHq7gqaaQT5UUmSW12T8/YoaJlB8nh3aWlDjdbTd0xURn5tq3g
p2de++jKwwkvKl2ib4UzS/vMLHPs94xPm0gFJfrWkalwWA18+Kkloqh4G0lf6DwU
zPhsgVDdfF53+7QXXD6r6wAiV+aMrx+IvZp8RmoF6FJGRAWqE2HINFlYrxhD6CF9
RfBUcNfVWOfnviwngnj2YlpXp6dMm1RHqVntCnPTsV1HnFAqv6EZbG748d7n9hjK
KKHHQveCXHEhKwQ+XdIFd/8qpGF9w0MtEEKSXz997YGDWjsaSIsyhrXmSvJfSeEn
OlJxuw7fMt7oLjOjGIbqDK3FjWgBwuQweXVOXkktWo9WX9ULKCVbOnKY5n6o+5BA
3jogsu11BKTJ9ezOiaDbc8Zp3csfEcOzBfw9hjFmOtIV8UtnOem5aLTwPMbpSs1r
L46Ul5JwzpBt3EeRh36rFYbYCuHdaiA2+h11qn2OaRA3gGyIyKI9KWytsxfZJ7F6
HhMmkw77CtPVk6Uswaut6xHvFyR9JhqoKWBW5Hh/UfrMCgENfJ3RPQBwG3S+ZyDQ
4Pw+fFXoC0kc89yNhe6f31pImqpTwhxi2EQcGZbBfMYgFkPuG7i+wY2mVQSfQM6Y
NTfkIL88sGZfYuaPFU00gn/NLc4VENTCX/MkTwRuqO/XKaKsKaB/Uwh65JOXfF+1
GOF1KVeC7utR4dISfztejfJKZK0ocGO6fjdx2lK0aDJV8G5qx8kG6l3iv3w7NRc4
bHcvgeMwrwDdfllur4fGAQvdWTJRg/f5liv39mvP59iL/OZXRtq1rU+oSN3QhTVy
/U58PYFJGjYmbp9Lu4v+z1n43jPvCeoxLFpiMcK178WDFCF+1OPFxx/3/6YJ0AZP
V+AbwXx35FKs/QQA2gltT1Qz8dnO6JghKQwI66o612wFH6318fyATWuj6kQcfFdR
a89kSOmCTXeP1Pw5sEvswKmRS3iAlNi6BCMvjQE2xzWpYOmC/r+qqXGUILJ71nsN
glK8sIzAtfWtf4PAdnhW9hRS55bkisdjamm/1tmxcZsJrZKXNw7qPf7ZALcnSPpj
cArd6TnOH9e8JkKTYxV9dkI8+Y/7Ps0QUEDMUuMczfJkFbMDdblyUf+1QRt5xdzk
02+c8narSSWkHeC6ht48V578D5YoBa1QGl6skawxgw67QEEc27timW5nWXxgEywm
wIKHuuGRoRTJnMKcHXBnuTmzxhWxmUFKmtasXmFUAhJQMg8giIPaWVA8bxDZL8KB
Hi0BDpK9C7AoNDmgHMsFbSwHL1GreeFTG63I5PYuBcryn15GtSIG0jmqxng+l93j
UmUk3i8VSKBNH3zZpyMm1lwhx1cCUmZINV1ihhKc3MUFDIUMk4jCYQUOyZqMGPvU
mGYbhXMuXeDiNywvPooWENjqejau6jmStDFJ+fMe2XcAew5Y5Py/HEyB25sRRQC0
um5Xvq6D2T3aleAGK0lqDWdxoKVYhlwYyj3OkytpWbXF7u/QBiW6HEryzfn4mk9Q
roitOp9pcIzywX4U97yJv66onlc+pgvNcQ75qDKi/GEKCE/TRkmcvuRAbs9nOafz
6wM43fYulC0nZY4nqwKdKrBw8te3gwbYHuFkq5wrARttPP+y4PBoFrVpPp229t0r
RuOmei+WWnyi6666hbCtQp53YYsCyiH2/ulxZA320d9FaVYyY3mJfOpmJQSCyEFo
FlU6KYdzwTqmWnKBJE/iwAcMmNO4eYcZUSQTHRJeoDeYkoumOmtKinS7ItDtJunH
y+/rH6lFYsVkfI4hukYm+FL2W40LIdGYN3ffou/8+L/hZzYebog34sA4OxBYsEq8
Xe2p8LAdaAm550o2kKL5fgYGERBPrz5y3qBo4+ie1i2zsaKj8rPd2BAgFTXOAFzY
cws0ITh9auKU8eC1rHXyA1KyBXMyfRY83yl56y9/P1C+yhyfYSnAILq/3rbS8QpF
3UvJk9Q9e3w3DfcAFwtrlqBNdwzWadriWdRdpFUDKsm42ozdav4D8hWM3Vgt9ACK
ZrKob5hjzabctuWC2IheWNS5BoDCynfM9odgb1FBhX0gkuSTzZsmxf2ZrnSwcim/
tnNTTQS998cVK9z1DY6FTkMJkHRLqKVVKkc9bFyw5ShIpk7mGUlBA85Cob7W33t4
6uoW+fk1QY4ZBqYL90ZA+pyQ+1J5lRmi21eYLZz1fEdjr7XmL2TpZBdhGTxd22wo
5OOR2onTeWY1S55Xxu9Ke2FDz90MO/pcDTJkMvFOFRzsaXetRenl4i/rjGfCw1qb
Sz0/d4y652aZ7wnsobmPuTlFV8GkHwVpQIv0BQBAxHcRC4Fskq3GbOeAOCKoxE17
FPgMGCMYEbwr42P3U2F9j2WddWpVrXURJl0BlGj1UYWzMFzr6TxzoHY8H64RsXfz
LCzCzpyt+KwFTJs03jUR60/i2KxpernS1mXV5+hjaiF3R9QCJkhX+e5JrQ6H6dAe
Cqi2XLF5hxV+MQ2NWVuWNmUJYa6xG3JWtyH9LBzpvGIyxKWsE4++vU7lnCCFdcXs
PRsD2QDy2ZKmcUOHX/k+FsFT60GAMBv8wuBq2Db+G1M7Pxew+ziDwY+rsPlNmEVN
wrEgRk1oZ9yCSTBFvrh2T7I3Ds+Ff+DA084OW5rSzJ+aQbekK/APSAnvpfMxJ86K
DgQUCUMV2/4lrrJOMeRsgFXLe0JKbbKkKgq1GM0OZzLNcSNYO4jRM5GlmOzGo0Yc
+dElQJ+uUuRn7hJ8HKlwoSGmUOaDv7BPxFIMq5X6AbuKVjeVmeydxpnaRq0C1IdE
oB4Y+SZj579P4oZ+/6Un0L7MTStKtn0hqQGA2ZS47DKUwMfWNfcujBlwfahO2rzs
SVeaYAGv8rTCAI6TMfF6TO7XfEiwILn6b4CT9tDHeboZmTOuM4tNJvYX23ICl19k
QRUrWwGCx3elE8d/p0G7n9jKrs2PwrVZTGjxfKsIFodVqvytWr2YAumcZYJLdN2O
N8gg3WoocP8tiKNYQ0k9WDV/o0LuA5dHM8A/gpUBQqDrpSDICd/RyNOTIlTOhgv2
QYM+EtyAhgySny38mMFXX6RSUTksLk3XRNK6wBXysNFHKujPDCAqr5sovA5MU6W8
zF6KtqWRPU7WKV8D7wG3BiFYy48kbjrNEPiCmHB4uskmADcjMW1FEnzKzrElIqDZ
ZEh6ERDXLE1GQFBOTx7FsvdS3sQ+zt1RSW9htEWNZJWvqt8de3UBHWHTmH6D6F1b
ecG59MoLBLCXdtdNrVqojowZ+jNdCtZkMJy8qkfPANY=
`protect END_PROTECTED
