`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4uyv7ThNwKq1VFVIUHrfB3Jbi7J7uT5Rx3/AF0l/EX/Rk3OVoDN3kjRX22SMF1f5
FDHpYjEDNiLljJu24uZMeA/9DqHmrcyvCb4xyTb/J6YjCUPB2XXUB57PHHR1N7Rj
SKNyyHM4iELmlruFTN5IeRgdU5fH2YjlxW67ygjM2xKucsHp/J+n0ZckQX2d/wC9
5nlBsAQ5B5uKojHtoY8/zYlUldXAfruvNUoZ1raFl8kB8qMRu4OPvyrKAtg9H5IK
80O8wqmY3As/1l01u4MRiwck7CwRvhPKh+bE/Mt1h/SfCGurCeAHMfR6xVhxnYOu
5PDuGppA7CDcqXbN+UCsqtBXEzHrtFF/DAwpRXa337BbrahjkG3+YvlCN9iHFZZu
S2ySb1oq8I0+Z+O7W98pebFOBPmxdMEoaFqwICq2nhmKxuCl6DPwv3pqX1pbs74V
9I8V+//HY9XESBdq9gGMKtj06MMvSh3y+xKn66zXDdwpMtuoOzIH5/J8QI1TZGzz
dnTbtrhWBdK31KwCQaTRfhUwOQvijjhKZe1xJ/dRR6L39F9VVDp/9pmhjHowkLSL
f6UxtTzO1Y3G6UOalbNl1JiIL4tECg8A3hNIUPEji1wu7qhLwVOaLnU1dduf0TQW
MBZ0+yOAc3/SWycRHccPjFGH7L/dOa0c9Se0AcoQeuBCF5GKs2bUZxOl7ZrjtE01
WYKlob3/oMS34Ws1KT4obI9gMMo9rxQ9UHITFTJ4aPRPAlZYeCQKatkheVyH9t6C
e4Ne0FUer5wed7bmPMOJVrx5NZOpE/QJcTwx7E4kH1LY2mMkh3CHM+v8wHQ6JTBE
v0uOMfy/BATbkbZvXBi3USB7Ttnwge65TkcOSjNdEC6IxBR+HILUZbaAi++MSYhd
xaVS+J2sU0MmaKnoAIUy5AitHPgQHh8bDH+YEkXVTOzXaY2SOdyOPJLBhecK/Nmk
p4GoS6/fBmfJIZ2Ch0Fxkrxmee6c00iVjcoH/jmypL9qql3OOv3KqYh7hPNl2hfm
2ZKw5aTe88Njre5iztWcf/GgfeRv/Xc2hzW6AszeE0HFxyfor/FOcRCo5QBoA0Tk
Q/c+8IErol6CBZcUNvcSndAg5FZmFi6FjH21iO4yc1plE316GP1bmx6SLSN3Jqsk
WKos19JXfnCqohMMW4SPn8EfUR9O9WUvp+py1sFmcT32Gkg937oNXFK2qrsGBVii
bI+17tEsW/yR8XAIsF0I38nAaHPqrqQqSFwPp4j526MrXCG2ommsjh01Jup5c2l0
4p5isKBE81faF4SaeLG+h22mg7U3KUrZ7pNww5kVkUE0AKEh/zo4kfDRSh2XgAkf
aQQ/BxAaybnLjEYkxqThqconFQW8LMhKJ5nz5QAgU7ssfzWBL5ZOgmcBTPWWPtv5
Y4N1FKWSyKCCHt7/qkxqvcIAq9G4sVwxvjjdHOAGd+o=
`protect END_PROTECTED
