`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FjBDanZCH2Kbahy1is9Y8zLI2zWYbES5284NR5WwEKX7QZ8fz+FE6IkrJzRI9vAl
SR2LWcmHnGU295ZU2lITLwcofKQb/WGe+nxTHwXx32ZhF6vULFs+67N58OfbhCaD
GA2/BcM8euQ6xX19wUfM2Seziy8gGqrNOEeNmvIlofMnwmNsJAnDU9MaWze7hMzh
3OuRb6K4qWMpgMbqNkxJXE1Lw5xuTwSGncBU2H5ZBbDi61Y4KicnaxvN2TU2fbHy
ci23WPMuIUCfHltJrxyZ3HCrv8gGW4JdFP+m8hzuxFIU6Yo/udBJEGdU8pOK8gc4
PnbEBVW4aq2dwoL0rTkhC/CZB+VElcw/Wrl+tS8kdYujwx/ifOpo7VJY/1pSL0VP
dPidkxoTFRq4aLSHX2rj3RpsU53+bL+6ZDwsaw8dAF0=
`protect END_PROTECTED
