`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYPb0/JRvNdpsUYFMAhi7z4Ma8uSnX4/cHKBU0Y7uaGHnBYoL3ORaJS0C27uiH/f
rDLkl7FdsNZLPYl8ONJkMwlXcTONEcuRyflD97FLWMFG4IS+XXU3pOBrXUoKqmop
kKSc2pCXjbL+H7ajvp/9liv0R62j0SgxgHB6ldMIA3/zF5TgF1dAgVJXKY1lyY9j
f4wpC/NRutiP9Lsa50k8en3eO+iknk8d6PIJg/OQx/5Alcm3+EVEiIBR8tPrxwSG
eqylfJZIU2Xqm4mbGLpwej6NigR8r+N8hQKU3TlKfTIJI68gJJuakVgVk5m4bbnz
OkmtUqV5YFAetvaQ95AEdRfFoghFvf95uVADUx9lTbNE3fLURaejUbueTRKwPAsx
NypMJuNC5HrzjCtru9EA18PVQfXMxMsbzK68SaGY/nOtncNduuF8iXXWsjqLDYb2
ilTT4ECJ1EFMoSs5aPOv4dixjH8TOY+4muByrJK/p/suSQgut/YTSmdnVkkd1xL0
vxCEtOSRnxUySQcn2vZQUCCOb5ZDoCx4yZlEFTdAVgQghfVszktgI7vwmqnQUtP/
D5PyIQzbYjmwFwpuHNs5DCGcd8bhy9PfJUi2nSi0BOzteJMmc58CF9Bv2JnPbr+l
fsChssvhOQWwqtXd3yolPHXUPg741fXoNJhvzcW0eESA6Yw0MPrdDprplfRzRRDz
dQhaMkIPB3MAsMlYV3LZGoMbpIrqb0/odWGMulTG2Yla3ak223sdXUcazudXOfwy
LIRsQ8aPNG49+3IQmjTqjGfRB8x+WmRxl1+EMyrWJ2KhT9Vc/CND4LXWA/JF0efj
shKA+7OJ712vK7fDvosjHwO9DncWP4nLGGZ+cV30C9i9NpjwGOSB48Uiktyr0bnR
Jsuzq1P1uHOTxx2ilHWFHQ==
`protect END_PROTECTED
