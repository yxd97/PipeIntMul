`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AQjcoukCUrTa2WVd1s98DKnlQyLMq7ZQ13nZVGd0otN9rrV0AfhSgn5DP8xcWZj4
ioWsvudex2DAC9SFS3rGUBjAmvVaHtw+kJcr+dZQiOlKYwOnNU8UF0ftyRMB0QKj
/TnDteDMakkMetu5GZQi4rZkd2Bu4lnFDTi5MGI3katz5D1zGJjsyFI+SV4wac3j
lGs8FJXf8NLwYhm4DgQyW3Uw7j9u7PPQJtNzs1JOolsMn65cBn2uSmVNJwQyUoTR
oRLTNToXMqp4rRC4XUphT2pJsoKze2TxCEb6m/xQWCwMk4DaoCNQPGOrcTdCs1FB
pA0MjQD+OqrBxeqpL8KJGD91Ks/OTee/WdZSZJXljeVV7KVgNrgdhmW07tr8EjRO
nho3DrTAyXnYgleQQcx8QQ==
`protect END_PROTECTED
