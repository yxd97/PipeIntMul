`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdbK8yBwl7nS+0JPhWMAGA4RoTFcBZxDcgs/cKiXoAh41z7p4f2R2iCeay2RM7aO
ly0785Js6woJ8MEZT5rDHlOsXYvbYpcZA+Darr7kuzM1IF/VQiF7L80126zBDeUh
BDkphhmzRRLJskUv/bsXGZ4/UX4tXzWjFNKa1frJv7CYN+flI1nIaOMarvaTkbNp
oIS7LfbOpFfk5GBJtK+iz5DV2W6ZxW+871pzksq9y05rZaxkTFWijZE+V0rZOQvL
26tfsLRk6jtvqtJJN+4aP+bAllzgjS+MpoSZT3QbI2/LjtO2SRlxTS9hp53/XhRJ
YKy1mjEj/PrtWU4DsFH6mFadtbxlN3aLVWRCVYMnumF2s6TXy46kLUHGWrAnNkVM
vLmEz1tK+j3en75vQiq3gKJAWrFUo2v5KOgRRqE6VoVCmWE0UEOxdzo13anacQSv
WsPpPpCByG6tChL8N4Ir2GGHdQJcTlLsYeBTn4fqHOw4S/HfJ8PiWFfs2qXYkL/L
MfkDrqL//n+HnbGZsmqu5dBLQ4QQaQYnHGzIIFu6wJpmk4r4cyxG8Hxz3zDcXxMu
BaV4X0reIoDMClyORRPmGXeVS6tEznvEYXkUVzsB+o17r9MeVgqoYNYD4Fj2SCa1
5hxLMoT+fWw1AxQg2b+WC9Z3tTH8fCxgnbvgImkSW1D7l05L4v5+wp7ZVLyAVi0u
`protect END_PROTECTED
