`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Yon6EP4AHVJ/9c/zZ+6Z4OVWbmNNoIey/YuUtm1hHBBgu3izbxyoFJb2WadEm8A
fs+LALfxuFP17WOCT/ihXG0wp/NTIsnmfZNnj3LZIOZoZCPAXGhDza2Y1LEmYtlR
de5XWdrY9DqtD88DLOWFOm+sVCFl9xVEZKoWxap2G5GLhJIT17T9NQJqIdVT/Mbq
oeCMa1oIx/6dYcfsDuOr+4CDo9ZYE4VR9e/fJmlH2IiOquF1pFby35FnoET+asL1
+ZUk/MOCwQL/9G2SHRNKwkUBNeIX7c/EBOg+kfNKFT9cayBY2Bp+JNLCjyaEiLLE
QLZQT3rsLbZ85yxOu5x6QqJUNsk0+9TJlJhpzhgnmCFsKz93ipHI6EY+pox6h0aF
6vM778stbf6yHE7LH4Gi3jLu+MyHBOaV8ACDaBGHE5MAeGQ8JkxvVqhvX+M3uby9
AIjbJFu7I6tAW8e88J13Z9bku2wvp3fb87cYf50rDwJrbS2RrYTcqzJ16p8V/jih
uLd9Ix16jbWCWHNd+ppPHikdKD6s/FgOtm9HzIxP4pYPn+WGiAx1EQhH09CsvvmM
m2IqN4mP/YdLHKFYJLKtpbTdM8bEQ+iTAQi3sMex6L3jKcjF5i+tBKbwq1Pu9P5U
JsBiMWsSDQlBi/3ncJbUn8XAxpto6C/bfbYBCopioM0=
`protect END_PROTECTED
