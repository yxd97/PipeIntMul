`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x3M5j/wcQEsSyfc7n1dBtXp68Blk1xDeGdSUEWO1Juy1hQip1IDUGnk2YOuBgDJy
VZHrgtytsGML4ZiZqV6EurZwmMF1yx4tJubDTJcsF/jn5alBWOEtvxfpxrhLOXq2
F37ZMBnBl9Y8P1bDrVkr/4wjEni47Oq80FAJQsmwvkRGolDVcot3VoE2b916yVst
95+u1pW//p/tAm54Diu3ripGvPmR+UJWYe2TA/XKUaB+oDLiTQrG7OZvItEpLYPt
bQacGy+zFP0UEQBuhRkxtZjebJcNbxU6rGzem0B88lpCzBbUFDWuUmodO8c++ICZ
p8DPmF9LPC4+gQnyaB2+W3BnUGLJ30mJhoQAGlYlI5dk/c1ZMvIa7nKQeswG1YMy
XBl5reS4gQjzgNRQ3/9vev0A+skie81VaAD+JKG1vpFfDdswxQWAfUHQgnkg4+DB
CwC7uQ3VTQ/Qeq9iw9ikcPNCRS74fa4zz0E/LDXnymnfqCSW89DosmxKQIM+665B
OLzUOxFUltan3vp/VlwDDuVKVfxeX0ep3iQExuo48eFTt+HsvWBI5SAksYgvtKsq
`protect END_PROTECTED
