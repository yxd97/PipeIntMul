`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7NUluMSkFrbrLDvU8604WAjjNYbXqrb6S7jzBQfRLDLagutmhOrMUKzs1sM1eK5
c+vd0EJNsdbi59PIZ0g2ig6MTltySdudh7hwfkCavRtb0IN93mE1kYTHaktOWNDk
kmeXQVhrni1rgyhFbgziD7hqMQ1uLqWrykKTDSPnfyQOv5YBVi66DA/1wz6jI7l4
ePnlj1QAHZevdxDD+Cq7v7O/r4gk/7Ell4XwXuZxKvOjvJ5wWw3TdlSIsomN2EU3
C1u2npDYEYj5WzQX1Jq7b+2hl9g+2jiGsGPgmASsO+x0aHXbHQkyC2lLHtXUewd5
6QOa9zVnwbRS47tws5MvmJf8ztobNWajx+3s1lpG8E6PlZe0YymzsBZZ8ncqO3Q9
l7oB6MMRc862Zj20q3H0Ysc5uOeZ+MFQSZ6EiiJJIxUblGD3Hvo7Jz8NzRcXQHbc
`protect END_PROTECTED
