`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pM/P+JikirK9vZ4S9kN2wPcFIlRboU2O5y/Innx0njd5dV98ob/N0BcgOvF0kVn5
llBt73flsuKC+4ov1OBT0VZYE7ze+2BYltru+f52KTXH2eqzp6wt5zu6ZZrrhUxI
340wKh7nVpBGyZb7neeLnwMU2mkIqFfVJi+ZfxEJYj1f4lbdSCwJ3mb34nwdKv4t
BzZb7zXsFAcOPGEHlvoOifhOR/Tz2/JBxg7cM6c4wPJ6mvgmCv8AOcQMV4mmYQuI
T7m7kV4dKepF6ndcErKRJJhPAFVFXxgjgZYp7V4hdGz0jC2E1l6MfB3zCole8VmK
BVZnNA8jmwSeQLghSz2+voGe7PSsVvao6yI959SGUSByD4RaGatB6URlKq8Ah09Z
BesURUNXKnxPTqpBGskuLzf8VgCloDhU5KmDXL0buSeNXj2MEe54JZrLpjDKHef3
KcnhzT8nFWTO0boCMCMCq8Cg5RL6d115DFwtR11aApdbHZhu8bwmQJxpNYKFXdpA
`protect END_PROTECTED
