`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/dcdQtVbZfEQ5opTHD0dLvE/ObJde3mAMvsqJj3M9kgGyhUOovJkYoynl4RlO+/
qDmHRNk5qe9OjkD8eMCwC44Nu5K16hgiVpeBVB+mh1uSo1IN0oh6Q9jGTlwNopeX
60h351LM9uO09Y+DUymA7voJNYluYj0EQTJHz9CxILq4TRIPpZ2+BaQ/V7r4KRob
rBDJeoDisiyfCP36uH71Ty6tQ7N6BVMqsqm75T7os/Za4nQ6IpcfzvMgCZLK0dbO
55P+9t5xR4pd2ATWaWafYkRFHBya0VSjKQKbX5rlUQ2IuVmPMK/CFijj5rbrRrc2
yybaQKY3eLEqR6VkMYbqA3UvN249h3qKiPwWFH18MZ3EAURm5wgd6A0/H7zpv9nO
M81ZEmvLpdCDruvkERCcI+n3XouxgAbkme+iBpkC+KpfGL5FqrL+fLjubLCNGUEY
UOaIHU3kW/Mva2tIPD8Pop0Mpt9Hh6/ELCHK0qnxpjXrHAS4+RiW7SDhRWZIYroV
VuoE2Kew3ObZt1ke3uKuHOtSxC0RCq+oiNH1voOVLRRntd6Im3m7Y9XY0HQoVqGI
nCDPRbtKqVw1aTmPXY0VcGJeZ/wMpS0SR9q54e3x2TzVh0RMbYNu+0P+x8XlO2hY
Ch7nOnh2Kf+yH9aSNA379422r0W8KjtRnE7V2Yiic1hZ1SsQjhWIvS5wDZw/+zTV
SX9GtZ2c+LKFwB7CrdQ/BEaVt5TERCJx6XZai69PpOc=
`protect END_PROTECTED
