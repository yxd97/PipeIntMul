`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yb8ufbn4M5JkIm96gMEOX9wPedCACQ4yefeuBrYUDAXJLOUzQ51eWqE25HMV7UOn
o7wlHR8RyRT53KOy6Nc4sy2estNA31G9J+sbXkeEMeAMUW7Uurx6QHxV5R2n/eZH
6q7bMtrPu3dVms3GO5h483YUNn++MZSK6uNfmOMuxs38PKBFLVDHdnYmD4xD2yY/
iB2H+FxVONICugUPfl/9vJSNLOXMq4w/snKaHR4SAMHSr+LnrxAFLgoVnn2jpGq+
zx5TadKwG26JVY7+4dSA8fXy+Mvt8NiSuoDh4XIMG8c/mGBT1Xf23wxpz2tyK45g
RCiSCUvOSiEnJ0P4IrVuBQfvUvlPCN9snADSiDR54RIl85TcMCHP+sJe/5oL8mje
QKPvcst6cf4lOyZwhc/CeoOlqbhhclttSWT6KhyYtQ1YG46pSwM/bJ1f7dqWkwgc
uGa/x+LZyl6acrlrNeO8hrwmNF5+0UnDmwy8JUJVb588c14LvRAb7qKg+GtaXeDA
PKwwqQv0v9Vvf3aj/fpHbtHPvKbWiihCRUzeYwqSe26NYMOLZdO+AdudKvSisay7
HF4hSjUWxzuC2h3L+bfTTTil1WVg0XdBHjOtNOf6ugQY0B47757WeOeWiBNKgeQj
P6NXoo7Z8nQKFrsKPeJhhGuHv6tBRbTWo0IrolqgEHU=
`protect END_PROTECTED
