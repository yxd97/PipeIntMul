`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+8mp06c1J6TU8+yXTOwmduYuZu2qAqdrqz+8lxfMChvQfnnWApXQU9JS2B5uQqvc
+0ZicSHSlV7udnQYkKnBTi3IWj0PZ5DI4wDhcCKRMV+zvhnmTFr7u+SRqLDJyRY5
PN7UK/sjVSxhb1GleVWFwuPgQV5n6u/5zCbPZEryCYQw+izELAtnF8oyUXm7hL0e
MFkiwEsUjYVEKwFqFHXRQxvVCyTTPz0g4ktY3ZxWQLgoJL69Wgv7EBWE8SIXwIXP
92/qaoRLpNUQEnn/P963Jjw2TW5ITltOzi5ZB98K2aQZzHijHsYP2CPI5V63Xqmr
RWUgDg9UazchTAYHBB62uVWcluqYwnsgpx/0Av7RyCdcYSYh42La8kd1EKc7L8b/
JbPd8KzB2OvviEmfcLloenmiTUo+9Pyj1fJDWCTqxrMbNu/3Sy9WujjP8aLOMBsA
5Kdlb/QwSP/Z3LkMiO5yP4UNWHT27I0hTszY38Mmaw+aL2nG4fqeDRBOQd2jVhmW
53dKBmGPG/PstIm3tWLniM0Gp9+Clss1Tth6Q2NfPTmpAOmMfKNmvPfy39zAJR2A
3ZZzhWMDWSRn6a+pYjNiiRlNEQuAnWDCCBO7jbxBr7v4CYFeousCZMARo7MoWjfF
x0HIoFdl+D8sam44MezVzA==
`protect END_PROTECTED
