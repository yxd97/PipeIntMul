`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iCG3z1DYCSt697JbfurdLg77bGhnVOJFCuDiwTg4aJjpbdbBEf0tB7Drv/lELX2H
23wEM9jHznvreJVKPcihE77UKddW8OCR5L8pwP7J/SrRdfzdXyAzmNaK1NyIIwQi
vmrRc2SCqwmd+OXgTq+QVHkq5MM7dU9iYHhYr7jyhAsE/TxtIJgkGDSX6rRRfB0d
MAUzsw4FnGRPmpXHiwfibe0z1zyfnZKKUusXwZUSC23aAn1viqd/VBKeqaw+JK35
Kez9oVrNPMNWu/oMyrmpWFEqy7axcfi/CeKeAHtws8ijBfP3YqT4eJuj9NHLxdTy
`protect END_PROTECTED
