`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzK2Vr7bvr+TqnfyK6DNhRsgjUck4u9RkarJvYWjJmIuY+7XNo5Da4/iUzvYESwi
/JusZkWHlzconc2Zotp4dpYCbLdEtuVbVrfW630u47neUEzQepSxMBjV8SRMI4uy
+DpdfCQdM3v+JH8jWWzN8cmMn4nsPSFbNrDeQYI786MZZCCmtA7jkZ8ngk5+vhR0
jCYES5JS3HVQekzBY2LR7Lt3/wxGgmdgaT39ddC8A8dJGa0CYA4YbjsLdAJcuXKJ
PnWaq9CSeujePaZk1pMy1gEfRFBUk4YwY1hD9T6ebXpPZORCIZbU8lTAb0wZO+aI
j49G+5nAYqq7se5mysGmoFkbvuSFfOyb+t9kFXJKNVQANkRhgl86Q1GUkwjP38dq
6o4TK+OUCkvzuXZt2A4VqQ==
`protect END_PROTECTED
