`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hm+ahtOJFsGBEnbFsTTY8L2V02EGR7NTw7rk3xgCeEoCntO+ETCWCMHnGiHu4EZB
1BokvxjYHasgYuWbNz++7EMvnDAhKdsP/aGOcbQ20agL14S0pBKcSuirD/CgUac9
eCLPQ7Pm9Xk3bECobmKPhiXXra/cDCkIOmD5FIoX3+KWpot9z1DNoUvX4QrbCA2i
aC2Gk6wJE4lvlY5JtWB4pynKvAot+pJUsBEPiKdhIx+0+SRCHzMii+AdxPv172c7
lXeE3ErYVtmDs8T4g61Y5tjAgRLkwXzYmpO0bAs5Sy0+NGdWbtEE9QcGAAxYN+c4
0nPewQez6uolaWAhmU3A1HCzvq3eCK7BB/FoEbyL0hwsrs/2oPg8T087u57+/VE6
UGNUYfUmfrYD6F/OtwyoR4fLbDJBXk21ajBjYm4t0hmmIFnODFm2ZB0NIkP8auLl
qtlrcD4wGqDqcBHb08ehVV/cmOy6EMBDL/PBOnNAsGhP4lhJCqzScKJUB380MVoQ
`protect END_PROTECTED
