`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJ9QXfDie2TDDqRr2Gnf7Nup8kdQz8yGm+FxOlRybtR4p8YKOTswiSu9ZQKokf1i
17rkEVil1Q8Y/3WibGp8zUlUUkH8mdnLSqoNBdKarthTFPfN93i9/S3jfJ8djWFj
vpLvBJkWIC9S31Q6rS26gr3O/qeSY0D1HMrdn3o+rV6a4388wVF+rl30WY8tRdPN
bRnXtd0uKWbyDC3P5RKo7CA8zr2FrGLMcUycDWfyifqJ8rK1cNL1x9ijT7TW1CfX
D0bNjgy8ZNwqSQlxuQCDcuo5bmGuU/qvvBc5cDyyo0e+xzvDDdUJl/1fHGyCBfEe
Kt/1tTzEWqgnYRcjCvhL/aVouQtEeRBi40mwxu+h8LY=
`protect END_PROTECTED
