`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhHPyF4LNgPpCEk3z0dhcEoaLhxm9ecCJAZ3pVO3Gh+gSoY8BhG1og4jSVUzX0eo
MfE3QkMCno82TaYjHXsZPGaV8mJDE+/HFujiQovaikyZtvnhHbewDDCy7MAM0JqT
gn/hJD7KbKydXcWmbjbs0pAaPS565WMF9z/e3KS1W8CoqcfF0dTfgEnGTaYFSbex
96wKnUvGX3gSAATq2oULtPyIl/qFgEDj92I1EQiC2/+AOAUhUDuaan8xQPwg0pLK
IHObbCkWDRw6QjYRQfmBVDHhigs/4mK6unRhSxnEVCHleAhpo8MKhWcIVN4FOkI1
m5ImN+6KZbqCB5rbgxm6BA==
`protect END_PROTECTED
