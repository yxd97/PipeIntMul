`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gLlcl3m+qim2jvo5RPHOW1zMfjKQAB4ZBANe5tOaOthllQd5tURes37hZODvXqu8
YpXYnaNo7TdOnKaiwMAKozNk13dnPIM9n25mRRqa1kDMGwoy6TmY2FqVeeMJFMfs
sH5uHuX/nRwShtCPO7QXqs9/3YKPbUnvKEwwlrAeD53jbu5RRTFHl8Duv0nrBDOm
+zKrYeUyQyVJwQP0Mf3Sly06r8vEghU+FRL9t+k2QJU9y/ZmOj80OdmecfPd34/b
TfuDrOqMDsBZejJ7rLLxtNQG+qpIejgXo5+uC7f4i/LMpV4nAO/Cbkh2Iiw/IHpO
5aQZiSaI/t4PzYNHTQ3m3QxtpCpt58QoV8ZqbuWMS8XTvbdSOlgtLda2JeK/x9AO
R566BepBaIOjDQbOwqP+0ktqh9QbKGM5WA6UK8Qc+D3kqEP0Y2jMqQEPpbYyPwuH
lj4yG2Pqob8oncQKhPzrKIUI4WQPV0ofYgzUt8Yl/1ZJtdBLzCT5Gwu9evgJb0JV
+CG/Nx+jRLH8w+4vBloMHjq4QrIGiRVEBqHJSXDeHvZplJZMP250h7fVe4tyG83H
Z2KLKF953hqVCtwnkONEum+NYAw6RVpwAzZkyYAvahE3K9I+E0hI9/li+5htTPuh
plkb8wfafaCJl2Y96Z0fUYXTnX0kjbBkFviPhwLZpnJM6kP/9Bx/lKAI3hYlRBbs
quY0LxjcuyW/0dyOXzhsr6C6n0kSe2rbQWBGddN2YZzgJgunGQ3A3lncr59TTUHr
DTl5NcAKbuYUuA3gyHyKlkE8ALfEl1HP3rTK17eHEjNty39lvs3jC4+DwXRNCoT2
AfaK1+P6X3OHeVR1u0jLn2aEeb4UwU7KZcRzW/bgplNOLo5Rk9QZyHOUORyzkgsA
sXvfBNs155CxhSxZ4day30/zPjkzKSRiRU5t9wPHPMnycKvARK83ivtfvJYN0kNG
ni0l3Qg3+QdB+/ryLX05vyYOXfbl2TcMTrvE4FWkcJYsi8So8fGYtF+nsf8lPggP
kLtl2GgNqHPolpl6syAjbHvJWsJTIYqxD1wP1RySJmD/52MFYvtKqd/c+ZfoWKSt
ynj1Q58WGS45sOGVlk0UotqzXMFW53I6dYx6Op6RALrHVRD4PWGkO6U1p4AvVZbf
yLDeqkE4hvBfLHGQkesmPJze+pso5vGVvpBvLIu9FYTGQJit1sqn41VAmU7zIO7+
6LZlqWo9JkUC96XSreUwxvGAp3IFwHCNU17aijfe4ktaFNuNTZHygOgoDOvAfVlS
ipjFtZ4rJ80xJYQIMRQagg==
`protect END_PROTECTED
