`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfnWr8rSSi8Pzjt0vJBCgKS3eyNRnAstke2PGLZ9t9TAj85Inwrk481nKeoM5uo+
wUvEbr7EBKLE0hwaIIzucMV8f5m+K2S45K2xcoIkbYbhdrJJe7T7TAZF4npKJDJS
7Pf1TmuzVdsgi3aik3VUMj34oMm7/BN9n2HfQqDAuWij1JHhrurpmVtNiPbiMm0O
SIoHb9YdvLYsISwRdNx5VlBmNi80kUAEQY2FXGrb0H8uINssaNJfkkYgkSDOts48
js/5994CbTHo/XxEf3gXxQ==
`protect END_PROTECTED
