`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zxqHPlYeJuUjBnFB0w6E+FJFGqfD8y+OLjrq/fAZZbFVwARlap1AilpxmBpdK2NH
vQZpVM/m6j4GtRQ/v7SPiW6zMNd2/DRSX7GNaVBBcODVrkRqbQ0WSSiEcC71Rkj6
30nXEZUacbbXyhk/zJSCkjl37obzG7q5JLhaiMrp8SEhQeAwnleuYrY2M66M7Ypt
IVjBKRsUryQ9chk1NaYsIV+r+7NteINbqEzYRJqfuWg9bosHsjwlNLQiTLO4cYHx
AXafDvrLbP/ZBNFdFWfgJxBJG0hCgjwJwVcqgtsXWxyHVtncoyeYdE5aCqj+9ZKY
Ax0vpgpIJcGgs9qnk+VCPqR/KJj4jnUlPiZjz29LDLJoeMxuKGdoC/G8TMET1M4W
/uFvHGvG1HqSzp29IhYc+GPcUJhND5MTJh2rlZpKLGRYrpmE1gnkBNgGqPeTPJeb
lRWHBQmGvox6/ck05pbQ/aBUE0wqgXUsTQsY5LFW9udePT2hegegQQ+TbyRkI6/O
oZiXhiWjmrKKwaSiYuEFzDNsuFV+q3G0GGM/VAth+aqv4xacDpiaa7rVGeSJfkEj
Pz1ZfN8bRkB4ZyPm0raH0oaMGA2q1k1/YVmqSEXBrfgcrnQWok2pImeHMo5RQOkS
8YoTRW0eMj4aEIRIK6KLZiz/zYELzNmKr4UbpANzzbNnxT8ONjUVKBL+xXHDHNUW
3GO8wwul9TamjhxvOM2drBTzGI3SdY1Uux8dscE/0lwpm1lkIiCySN4+xqMmKDPm
B7wDfAMCzAoCrNNFsmvgZROY45g/tdf3dfG/q4lSLG7bJDqzjqANqBOhrMd9bxWP
H1fJwhuKPmLYgT/O+6XyET7I79xJL/Cw3bLH+x4G+k8NAdGo7eHtril5c0oMzp0k
80rQnCvhIYDPObyZoO7uD+slIidOSX7/i78pRpmeqyfoVLWM3Ep7s89vLj47TBQc
9X8qR4/JUB538YG3ahEysw==
`protect END_PROTECTED
