`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
liogvAlm0peaPZPqw44b/oYWwBGBw3XxSsmAcibLMUbEEpEj8Mj7fbNdu6UUfzpe
I/8/SOeBOvcIOLwcgOeLRXzITpkngHaK+CrhR8KlwkbhnQfNEJQFMA/d2gN1v95i
9eeYYLjXuASnHwGzktex2mESoMVyBYRzfDlfEo07Dn9isjBw6yUKw3E9Y7ZdEhPb
d/XpR0asxecfmzDJANsa19pf1rCDjNJnIWE8fqYHM+s/n18Zjt2ViRZ6eKieTk6c
FHHafRYBXO/Mr5Ta0yCjAhagqSMTPGWecQeGzC2z/GojoBGOfgTyA5hpSkGxdtwf
n3ePajxGZdAgXI9yYfHqeMDce73NMecgunRUsc8dXXIH+c84EzF5dtWBwJYuuuEx
4KMpAcRyWb1c6lqK+MscsvLL9i0BI3es2CC9GWf/cUQkc9javG7aCgdtrKNR3Zgp
b6PWsXWzdbL73XDx6XJgT0qZDHp2ifghJ5KtcCXRFumT8aI97xWNpoWkzECn1uVf
ejTim2BHiZY9+JuTzxAYtGCVEMCv6KO40/8A5WRDyMZeFYZU1Umk/zHSgGkoi3ly
YgAY33t2gukElds8vAQCwag4yR79teLBqqblJ6shfDmuoG0HYjctzngoZAhc3zu8
yDrKAxTrL3X1WdQD29++h2iC66YrHYNI3nVbC9SwwwOdBIDJeFTyAI+1ZyqPlfDY
1zBbRENEHuQboO0fjzXSxpE5QPOQsrg75s7bRxIIUwqHU/KsV9U9vOSIvpRgFk+K
kfsLkDiJr/gZ8wJbuytSkZLGjoZRezfq/m8+dRsU5oDDLj4hjLq0/AIy8ilN5JFF
80BoHDfOcw8GRw7AFNbTunmUA4q6n2I900sQl1+TF59fp9Pe2PQEn3vhzgaRWQgX
j0peq3D2uEhtzHhtZffs8gX16XareMllblVwLeiyKMwDdzZqAFp1QlfXxYuS6TDm
RggzYf9TRiK4QPyPQTJskQ+2/ntHSQavZiWVVoyCMVKZil4Jl8Afp894hchkRaXq
aiB++vZC0SHG8sRwJazeRSlGOEZuwdxw1Piwndrvt2BMKF0gcX/oe0GYte0SBA38
cQ8LGSsyOxylSsqlYWjNtAw6RZ+PD4pHi8uYTZFF0Na8GZf10w5YGSzmbv6We6F5
DbWcEx4ObdqjsfpNNHaqW8i6oEy4YOnzYV2MYOIEDo0mgoyP1sS0kYG9SyfzYi+i
gZn1KNg8o8QeYKlJCp7YA7YLVQm9KzkHCADP7YSs+dqOWwMLMHRJEht/mM0kYVJh
abUBab7KMpTKhN66BETWmgMYTf0usaM72dvSNyxiB6/FyJMsHU2V2sI2ix4wsIIH
eBx0NgQblDW3WOar2Qkotbtjf8aa+/44q0yEHC1xtKMo1ODn9JoM6ZUa/9ocujCn
QTE2ot9O2JUmpHRAOFjUKQTDjBXMQx11rTh10Li1sMKgpgUnYzSUQf7nhlE3ClCB
Cm6Se34xI9Tvmul6TizpGcXzqQY1ZU+NVzxd/feXqu5Nc+Qap1c8rwPSoeE559qv
wgMu3+1Hq5zeYENtDq7B8urptGqnayhOoFZqMkkr9AQ1KsYmvyLQpL5eyyjJQnHo
NDBsstaAT9wxg6N/LvcisS2iOgjqKbsmI+ewyTC2AqQrCfcBQckL6BSlQVlSjAuW
4XHZzRSdln8+i2pfxKKGDqbmmfjooE75XPX7QuQvWx6F4irwGXKGEMXFWwiK4hyi
X2+Dq17mqpPSbT+JK5jEtuvh8qizbZ8m/K8tpl1EeZS12QtDC2f6jIK/gb0XjE2A
7gpd+Oi3Re1b+WW/8+TJbmwVezOxPLvPdberox+tfcLoUA56ITnHcIsjgk0GnjE1
RrsYyhRMCRFhBJPfnPAijhJZgXUCTv2iK68uo5VDwUc/1ngr0k8RqMqSbrw1O9Fh
1ipoZv6kHWUdy5EIe853i0YJlPTuTgjQKaF7HuWpWz3fxynq/ROFeRGujnxrOq5p
JMdD08NQvS0SsClPMjix4eOBqcpSun7SzeIvQ1AoI5CeIzizbFsdNq7b3c398YUd
etbM/Jbo/6AYy9hwUrfAu5EVQBOPq5yWNul5mumLqFo9B3lRZ1YKwJwKtRFgry44
rOQPsgQdxViluMgCqgeLR0grESF3mRL2lsj0hAicnOgOHIJivXw7wpv+16f4sa2F
Ax/NUqeBQXQFrUOEAU441Y80bEpCrUiOdIaG+Z5NejWWnWNTGJ7V4ugXO2/5bDgx
lbfF2f3miqT0iYbkbV0s+MmGu7vNpC6+4YaXwipuqq0/l3da0CMB7tooFKAZ6DiU
yv4A3KtP7V8Ll6rAjFdQ8LboBumpdtr/U6QrAaAVTMcIB6WBKYhyBHT64QlJj9dS
iHq8UlzJDwdgqmk8/W4T2G7d0nouxDTrQ2TCGTpqRSPIE5cgFgLkH3RQeMdzEtvM
rpQWkT+fmG/xAyrUK/3ubz1yYnp8d2zrtzZs73hhKEoniOsH+SrZvRkIk1L3THdN
Tg2+zBZ2yfysdouhSEHnTeBH8tM7nsKEUQJktti1S/7vV7m76u8w8sWOJ6ScIIBq
XviICF6Xr/erH42SKKfEBgZgSGYbvlvmSXEFQfIu37wdA7my3/wRT3ln6Spsv8fF
qQY+Pugtu60YhyQ9y3gcizvHXp3L2G3PuNu6FXeQM+dIevhRjty/C76EyJTSSlI8
TE7VWIqxO/6NLSsqaT/v+J+v5DF2fV2/ZOs632oujBKJDo7qWktySW3DUn6ylsju
bV/i9zj5+GLLVEKQRy7iD9iNBJkS6cNb9lvqfQNtA0pCsq4T4bKyyxraGFwLEcYc
am3O3+TnucAEyBsYzNkrfVw/HHpILRzFFtjdPcYB9g+mwZO/d4y8Xnt59FJeyJaR
Cb0inmhihMxdledHgc6YlhNxsK/KlA2MlZvJveL6rqaeRnTKo4FI2C+QLBnMahjO
oj7lIOp2z1b7VIFVluMadSW0h53u0Lut/l4Qs7zXu0uRhR4O9TH/N1nOrJ9J3lv2
uuMhyKkmJ2cxnBToImJ2sHIe2ra6+85SXdFM78434GySKToatiVq30/X1yZRdAtA
VOsdqH8Xo2VZr4DGymgBJIojMy4+xbDOd/jtniS/aWGBZ74wRX6NGLtbvSzI5Z/g
LDM+iJS12lnkJ8DQjPNQRdSlh1cbRU2868k3bgxfWjOAGJ0bUYlVGka5DryG0wIe
9L7US2jIk2rnSIn/VC/jdHJUs9eah86Y2HYXFeWyqnw=
`protect END_PROTECTED
