`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfItbAT8Qans9viYuDbzr8WsUG3b8bMA6EaM5vFOTjHzqzTxE1es0bQYbBMYFP/n
GNlLQI7qIVfzkN59gc3GrXza/HoWcqccZ4sRPskZwMLLaRuTXBMSk+wiBPAaxDZp
rJvcF/SsQ41nSTd2jwWSXLdBQaM3N35l90v6dDNbnF4ay0muhPe3H7WvlNIRNWC7
MbMjsDxS6x8aUZJ12ZUaLtBSsFQ3qvC/7DHprIbHGJ2v3XzKOGG/lLC28SU8fJzZ
+tM3dOZ5Aa+TZnrLRbUPZr2QkATEMdvQNPUeW55MCAVuH62AD0WQJiCf/7Z+Acwt
dhtsld7KTUvSHqT/XZ3mRMdVkQdsRVqDCNPfwolef+tGkk3Rf8DkyU2QeR0SO0VI
k2Z3zg+JCdW8R0jRCgQKxcpQejPuJpXsI0yLqHWrv3/ElIOIHHOTEc+CP3tIjZSm
Os3oIATUlADAMdXuMW+tPT7Y23UaQNKTvxTMMDttKuBo20/4PHAj55cr1fVuD82e
8lQI/wM5dDyGG6E5iCCZgk5Kch0/N/vPTCPUDrYeBtn4hnVAwSE300gRpc14tcQo
jSEOcMkS1Zup9qOeyB4QeL9NIQUBBgFUz+ConDYC1VRdXVDr3FRPigcUduaOQIjL
Ne17pQFy7u38PVVLH/T2gUtSrJuKl9zH/hNRy+0vHS/oh0C9vG3u+Ws72h3Uq1CO
`protect END_PROTECTED
