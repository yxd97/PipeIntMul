`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jtLBkDCHItMKAfWoQPImjyrg5t7cC8rALTRywaIVACCgOH22P4I1bbe1iFj0YGs+
gSogSnc7+BnqkqwkDB26W1BJYuQ7BDlKsVLW+QXR+ar9VFedfVbxQM87GZJHCMAg
GssH5ephE5fV1ce7IOZPuPeMDJeylGN9m77bQQJNbRsoZUwMiwcyq9OTWkDJCjgu
5BcKmZWzffWV0mLj9P2vZ8XYynXRoh38IdWt9QvwSX+cGGll+LzRpF8Mo2bU7dG2
pUUWU7b0EiKqfoHUrvIHvas5W/sOJv1GCWdqOu6HWKP9yM+/9JkwItGNQi56KmRc
hpeX4tMX8KZ8l1LG4oQZOthVm+3/yCsTHbzF18rR/u2V2NuMpR5l90Oi9PXbHoSL
CjEege0NBaYkrI1oPiVpiSmQ1pYPLqmFQ1aOMY75vGWTxD4KOppLGC4LD20blMIc
EcGwCB38bY38Ir9r9YYSnZbdzYd/mHZ6gpXYYk7LUHRJM0WNZZdYeoaOsbmtCDja
qgd6nALxsbGkrTcpxa9M/yaTGUEtqHGYcgSKIvtTXq5mBc86hH55l7Yo0YYoPITU
wmk6++YyVgJ+ENEfUoKFIcnFIYOzuvmWMlPcP5x/q38v/N/Ea7QEZ89a7F3okCQ6
uyQaX4sCW7v+3xThT8jVRasxKtF1kZ0YoJfD25qt6JuS21LZ7kB3fxfIabksdRQa
cpJnZWien3Qc82kO1x6RerjghY//v7zRQ3uW67T19DSQAP4rA6usP0mLi462rikl
gNjgQsJBe0XTaNDEHkem0m0Lou7j480FL4v62wtVRo5yQOJKDFa3gpSKQ+OcbWLA
+KgZIICyisgevXCW8z00USr8AJHRu+OsxbyVKY9DqOs=
`protect END_PROTECTED
