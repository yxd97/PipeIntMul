`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UxzA+xmxpZZiCavP3mnFnmTjAll+5qyLILHMhrFLHIs9HYOIiajX/qSLn/pA74QM
zafOe5IwapPv6vGDQKqb2mZBYsXjTDp+eiiAnAvitPbpI0DFQreExgeWt1U/mJ9z
/kUx/gBBnEIEyDYvFfZ2jfmWN6QJOl3ah/P1pC9pY/vxpKQtqdMUHpHIgoDf5Fls
haRfNdO5NAXHoWvmp0jEfumCnBIIkLLluACQwUVtoaHBjyw/pMfaVpN87GU9dZe4
5gpgNmqemaXYno6RNtjImMjRo+7e+ntjkp1ocl0FwtQ6i79A/beBc2LCq93YHrW4
81CwiX47x0Y3/x+HAfL2C5U9BYkp1tmdLWWOUOMy3B+RHuQk78jhub1MbbA70yiX
oDz5FGlVwFj/XemWa2y0BxhFlKmiMq3SAVBh6LIYRHgqY6AFHpagcy8Dpi7zS8+x
cUWk9Cu7qDD4MrQi8DYuTpjUQBYGL1N9tUQNpg1pBrunChmDBltemxaA781NyP0y
`protect END_PROTECTED
