`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TRzw8agwuW4gKZU0NccHiKHKfZK4NRZ2URvifcAnpev9ol0PWKD52dZSyzsZMDrd
w+YD9AzW+DyFmgSLEH9vu4tJMQntswtYfwIS6LRTo1C+v8fjztRbhX9S0CxUdzsC
6oWGq2oRS6mssN+Dre5pTpj6dT/zV10buLl4CZvW1+fObwsas3rI65RCD9Lq2X+q
Gej+1raMTWzDgytltI/EBGlqDFDIdo0eEdiR1geptd0Cyjb4MWN/alRoYd3Z40tt
`protect END_PROTECTED
