`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7DrzwT+3Wo8tjcwfoodJ9YpF1LlKB2RTtJiCCFbbMBW+0+c6trgOqT38/KqP7IH0
WgSOkTK3tJaMu83wbQd2anpeeErxAlgt81t5bv54+uCG1YnCuoIjYQwlQxrfG1kf
Aa9KNSA8B1BCZlAYyfFLrNkx/Lz+s11wHcByuTc/0vEKHtq2fg8cgGEeC9nblKUg
hZlNKbkiWiuwg/CzaaTcoWIM3cR4+Somf05OfQQ5+LT54LE2rrKw5Pe8ev5BPttX
M20KVGso9ihEgngm9dDuR4KDYT65I9m1nyvsBwzr8L5KuSUSUV1guDWJEYnnNirl
BMMBXj8ShrxTllTNwqistg==
`protect END_PROTECTED
