`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzWFdVIf0l/yHIkxRQCwTrI8iDOyV3XwVatcjYqPDVRvYpEJH0PloNr+NCKwRqKI
jNtoaheZxEiiEMPe7ndS9u4k1BmPTEOmW9vLXbfstbcq9chyazyZpsAG12dJUhbP
wC8lfleaZPPuDdCrBvXUef7ru5u53haLkfV5FMauDFEvhHElhVJzeh2AZXTFqlOU
DlNwoVtaQyYU9BHFt10tgZ1REiRbWG85h97LTdUwAeHYxI3jYHo6lHj5rL07bQIZ
Ij2tPnFeiHCqWFjh7aI1lwiOGrmB/SBn47YaqrEKG3uPEUtmMen4iVGdu7DPbGPi
dpqLBwVTUnJKegVTFj4Zfz32ILy2cyXuZOotpoLf2wVACdKFo/BpEqfv4/QzUx5W
LRSGxlK0xfTIDx7w3Tp2J/Wk3t65qePkZt9jalVQmYFQBbo4iO4pcxR4cM7hCfV7
w42T5gBxb+H2RpASHae9rzFtlnY/ew5MLjj4RWegpKVF2bIXjNBQkJat6D1ddfPE
blFAK8YygTD6ADfiyz1Vsg==
`protect END_PROTECTED
