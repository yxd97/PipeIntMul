`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHHQeC+xsCYd6VdB/1Up9SCQpA+ZhxzIY0QnskVTe17OJrVu7CjWnu7MKb/dX7OA
+NRtpKasVDbkiXpq3349BSmDlzcw4w1UXubrYvA65wIi2Ecsec8wvOkra3bzL0rW
Cvj//hNjjK4qbFc4jIqtoHamRAM6e+Ek/9d++rBEwD7k87t88ZvhjYSJE8NsDrRY
nI0faSnNsQqSuV+e0vxP+EO5TmjgrAnMXDCS6CXYQSkP77RcP8auEWqBSNsO+j6U
7EjgzBuZOzzfsJlNJd+KwaNc1qSP/u9J+FyKh3dJ6oQ=
`protect END_PROTECTED
