`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fbfod/4zy6xWxvKk9k8cciWoX0gdAcBlvp9RCRF2M76PxE450EP7m2xuggEhGzgt
XPZqAiBLdmPRcEsC8l8xQU1MzvScIfl/ZEPjlMUjzwCYODOTUecMTTJOjRxwCvxn
pzRUk2Ivf4S2lMgUrNYMaqkak7p0bevJBC+s4Jfbz13vl3RAl1g6nRX+N7yXLixJ
zNhGb/8hg/JhuSsgFBfoBc+GVU6rUlrfJc+PRWhHAam2yDcPOd17mcBMS9INJR8R
UZ6hJXRRaDbpOYWs1JWR/ZqlUHhFf4fHpUrdG6awlpi1a+lbgtkTAbQX7sNi+Tw6
OmZo5/F+AOmLGr57GVDDnrS0X5dJnyPO86tCizJnKdj3vcFx8ZtQ1W3lQqz2D2RI
ceemGbt/lbKhRlHgGD5RXxBYAhIejvXKr00OUa1SKC3wkCCXdKePi/h1YHVuIQfs
3lpGKwR/o6fgBVoGrfqrv7uIkqBjLe1Zo/SFL87DUeaGNl+KjbRj7JD1ix0EUOfw
WxRU4xO6sweTWJU63YRS3gmZ9IgPTTUiEX9AfRhtGP3zT/iWy9uqcovK23fJnqeE
kdK1ZrDvfmYnmeyaGwjTRQpNTNjL2qj+VkAXE2zbJKg6GHlgLovFjci1YDkiJTp8
CP99KYRjD1yFa2fI4jM1voTW6sFMKgyuvFzPwUDEFy9cxgJu4H5UClpp+rAgYqYV
OczytcZi76nX7i8ec62ipdD+s7Ef1vs1Lxjsf2OQVbF1HQCWIqRZjjPhSW6SSxj3
yofB6MxUYqvyZDN4koRlPXVoRsTUlNq2yEjNwCTPfYKS9nWaKAYb5r2tp3uUy0M5
3Cu/b+jCh10g5HvrFaPqk+8kD1QAGNo8eBHn2TaFipvEel9JJG3ogNqTZ4LwDEBH
Yv6083qC5DIwxDNxViKKo8bPdFtMhj8b1rY6sFJCcbes8L7gmB/qlgrDrLiniONI
`protect END_PROTECTED
