`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DcEEfzO4ITJmQLN7rztHMvhshTZt4Q+7rdypD6NErnCe/GDWOWTU2F+xEDUD+YB
wvdOIz3qsqovshviWdSmOGbSpMUVjzS5HC9ephGC9MhybuDeQl+ZpzLbHJloM+5b
HJv1sk7vw3R03QDyed3Vfp1Egm3sZ7ZS4e28yvPxxNuueEAOhGM80x6ayalq8ZFx
ZXDAzuK3FFa5AgvI9o0KkSyeZlOkiIk1+DhVY/5Kejm0iDyo8WDmaS0c80g7w5Bj
g+FmlMd6oexpFxcBbLniA2rltjKXPaMAQ6q2LRLlHEa6faRDQ1wudGwUTZVAYna9
+HO09lsL2qSZZDl5Bq0Jw2/SXjSFRB4pFxJzeGZ4e94qisa3vi25KEF7w1Gz/Jkc
/a1PLZB68godcLcYCB+db/OiSo8yJ5qDS0pLWAlM5Ei23tZkhWHGCXH6NsH5p2i7
D9yAWASbRNs3dtN3hJf9qxUWJpV35iht2yI2yGFae8ohKUtW03Bqzdkz2hpd6iEj
W32Rkj7nYEJD3aeK//ilWKcLTDyS7QzpC7c+NNL2gitY3Jz8N03TnOIl8IM3/Oz4
4LQ4z8zBX6x2+cb+iCbbIHVBVKWr/jQvNthwvbTyCJI=
`protect END_PROTECTED
