`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sajUGHyhPV/sh4zE3yz1NbkZ42RWj/YvtBehXxl2jrXiw8yoiYPViKqLm5Q3mb9p
M88ZoFx9WH2iUNoNcHuljZ1g3Lu8fATBOvk2oBvIpvfxM/YSMDJGyYnrnv5Om6eG
bZwwKccrsvTyrdoX8N1bazEqmB1cKctX1ilFaVXMkhTGcbTzmVlsTa4bgDjbxn2p
VtjAd8ss/Yp4P26rvUIMCTHWFmdlJ0E8aZ4Gomk4PUjC0eMhVtQ6BBaMzzUdSrUk
eEJx6D0XCFYmjEkT0M9I+drHjRtfCn32HgfQjWjmmXoj/5gNcxSz6fUcGOdKXKDj
Tecj8Kn1bb9m2AZsIK2RCBIOrH7+W81CkX7+A1WXPP9+PSY8UFNu3WGLhThaRDxD
mP1D0Fo4TIigbGYgTbYkEX4gkRN//YEm4+VbRrBTywLNM+fp3bO/X6z8+i35sCcR
zxKJ0nuFbe+CkNSValIGVQ9VXXz5KA4ECWYRkHV9cjaEefaZNCirfnFRSTW7Y5pB
2HDkIVzWgLkgYyy27Izix0KGZAFBgMxI400n8IGxj3+uQDxjybxemMukv1EaqVJW
DEZfcKmE2386J6rvw7bYD9j2i4Wj6/6MZwOdK5oXJ8hcbQURNwwEnkOWv2aEYtVO
jm3AIlc3E3pCTi0jwfxC7Bklgwa07jUlnJzueL4CGdkAhr40ukTHZHF6linPpDSu
4Ci8dMpHW+lkV/cPl6YCR+mwP/k4soTQ2P/35kXcjjnn2yWbZ4xeoVPpFHSatYnZ
Y4wBOwYxX7/VVP/Ic3lfFt8nY4XK7gpGLZqf4mC/YjYD1zbtqFQOJy7lTH8jx9eG
KRaH0Yj0ZEJjfaC8HbjxCAghOP5W5lDp1NQRQB0xzqwJzaUEXl/8EHNsKSOyxWYQ
uw0S78aY53+ZqivsxMf+7iApYMWXuiTHqSkvuOgsqTfRZnZxVc2BsAxoVZNmB79P
Ft0xCE7ffQMvA43ZN7RJWEb3EsD7L7VgcJ9/kjpWjYaovEcxV2tF2+6KgvR4hzSq
XZWTpLRUhZqX0GrSFDDeFuZQeCLljoOeT1PQShFJspwQt2Q//F8cdmnWiH1WTj16
WkGet9aRJe39bGDgjYxVJCQu6GBMA+3sQ4Kf3b6CWRzqQJPxg+qlwKx2t9XxXd6T
pEJte9BgXPsZ4aIlVb26EXN3ULbqcYYmIvbSVbN0sGWSZKpZqLcLd2+dS8bRpBvd
S6Tu/6YSbmHQRdKH4RS8feUJqO+inkft6SCq0k1p/PsLkcjZJNFHbziA/+ESOebV
KkCaxE9paB84I4rfl1wc41ybUuKPy5NA14O+flXblCJcVz7nCi9VobEnKlxXuz3v
9YxAXAOn6uv1+r1P+AkQd0O1aPnm+D/dDD4hFRgmM3AqCh5rVSezvoqmNqbyjRBR
t76jYpXf41fsvvWrLTyMqM1GMdzn1Mka2aL7rQda6VUHMW/u+hkg8XW9iO6ojbr0
GKe9wNkdJzhGorP+7bHE6/d3HdPiqJjY6XC4P54o36hAIlb4T6jfvGMv+PAwWsY6
0BACF71bq/JCxMvkp27K0t88l3vv6wHSOfkKNKaZdQG2sWPJnx7mA4mOpXf+RPcX
H7xH8ZyfetloZ3KcKIRx5qjP6uER072Z1ZAaOjW/GCmUzGYxxZ5T/CeyY/2Fzpjf
mX5Z/fsaKwQ0RvAyiYROzO+7xpoZykx+8REgaF0aHr2wYy5ArWMWmAjMj5BUa9IO
wbN079jk1UVp3UU54I/f+0AXqy/FneUybPWwSuf5uF7R/ycJtmK3VQcblaIENNgj
Cv6m7d0yoztrP1AcqpkNASdr/NqA/wDGr+gD0/84HnWKGtRxq38WE06Uq9p4lX2C
sQ8hVwfTBBwHaYyQBNZzI6qq49fmz3X8dzG4mTl2K5KUM4JSLUUSbzQu3Ex1CV1Q
T+JAfFEZjj2LvvzQn3KYIs5+viux9PQSwjk1OJCnUPNKal0nJRPI1xDjXaBfcu0Q
bDQs5cmvNxlGmBR9TwAUKLjw+fXvtc4Dzjhju6HNqRBHzIvoLOPBMv++uO/pozsn
BoJ0LuVQfHV+axZllO39ULyyAN2EcI1IpmzJDEIZGY4HlpBvFdKKR2SCiRNw1xB3
iZtCk07xLdu52V3kkSE/D1mWjKsjtPA15uYlcsS1QritAEzVM7uGoIlX7rHyWCgC
h0179f79n4gNTusTTdkQKQialzIKm/km9sfUCj/Iqm/12TDe5lrYFtr4+NLqfM2W
MlgM6mtk8+ByqG3hEndMk6+dD9z4ByoRj/Ef4aJaaOpcPhE87mshB+tNA6xcWCbv
nx2UvdrnhBON7leNVJaePUedvj7AlToWv13F/c4xkQSVqCcvMGcpVc9DgFqijDCP
m81WDVv7xSAq8Ci5N0/3pMl0lNajrcimN/4K/II9zmShnQXALYzY5dauIkD3vN4W
HQZeiuNeCAsRcL2QXQjNxjjoaJ/5vype88sc8HpBEm+ahY+X6jyKJXUJiFC4nWh2
VOEu20BtmzanOgFzWlW3BDLhmamEGPNurPeIQKEfY4FDTgJ0iUy8lidNMbmxKEwf
Q2ICdyRcpo0khiYKIPhLpzKbLTqCxY5GVhkBm+cjzsQXLnTMJ6KOFMUDEoVWV1Dt
3QADPsNiJqHgm7+jHnE1wGcJtZuW6sSZeNggwO4XrpUj16AgIU71nWnGbYZa82ne
uN6NiJ2kZT/SCrlE8jaf+MBUWDdlkn8V2xUsMvr2q5Da4uM+bVrHfZgaE1wRA+Jz
EeNBOC1NdxvZjKBni75NseD8Segar+7WnmSUlb6wG0RHRoYpLjvlnzkqgE6+itQJ
2AW2u5zAy765IcIFmh11kvI7VVkb7veyvbCfuqZ0m9jt+DSK4adNRQYvu9pzZTUA
r3vvUbx3s5S6KuZ3Dw9Y1AINMe4eli8SB8Mal3Za84MJ/llycX3y/QP5xM3tefIb
AigJbWLd4fCuyUIIAAV9JcmdffMW1Rf+rF/1Ychg2vr34yCwAeIuqmpDGUqBZefD
Mus2Lke840v5dtz6dUwi35NXnJnaSzwA4DP8EXUoEvmMhs9oXMEgQ7Kr5V0fz8rS
bSz+o01EPX8umiul00OM2QK5zqKmZvR9vVAXgRhFchqNJgwh9n4WOH1GNdf62bdt
TLweKocOuxCXC73Horenmf++DJ29TE330JxqY/Stt52SGMWVCr5QNjlPzoqMnT2c
bqyEO2w47ztl9vXde54n4DZXyXYhcTKNbzdXM/in3NVfG4i+VbFKGXUkY78IL8IC
dAb0JAUo92FzsrsXnVVBB+PG+rUtmL7GAwPrNaE7KcQgxqIV1fmEVj+9FQTR0rgy
+NOUYG+lIhg5y3+ZdLjw4p8Of4yCQ4rKcP00HTaKNg+MY+OkIQJOEUK2PdGzffMl
IqgitFgH65en2rstBlPJAtw4edgG6mNprVUuUu8QrSxHixWLOKe9FMs5q/QNuj5z
pRLgepVBC+hU67cjHc1eq866MMzT4M94Z50Ns60mjMcVfkXTv3+s3bfmXvL1FT6c
2bu9I6W2wZ/iTImN7ZsTnvGvV1XnAw4VategR+eSziRaLtSytrcmzTRwUvkRldkE
TGOZAHbGSqFyy6GGWEJb638XPR+7d0uxXHSAEZ30yxTcSwzJrWldsrjEvyIJ3oVg
CFuN7p7tH/7z8jjceFwVT9qhHZ9LT2nmMwMy6jrvs44V4++wiyGJl4YNSPWe8mjd
SVD3WnoeZYb9hMKmzZuQPrI4tUydFN6GkUhJ6XO8tm1gTNg/y/UXM4el4tga+yQu
ao1k1gH4MNT3PgJBAB9W/FluymZlCvkVUAaoEdFR49eAblQB0ZS+pDl8KJFsGdof
TzhbXAO4ElPMIRFHxw7xPjV+b7DLGfwlJ0CyMY9k3I7X/QBpemooIX6hfn0rA38e
ETqX49zmgvSWJ65j/z2WVBFwiLLDBLV9MNx54yn2lssGbRsfSBV5twKMlRlMeiIv
yn3D7AVoMk2cwivGLjkLI+AKc3mXGGC67iTjpBmDPANnxiuBvBuPctvBtFtIaSdZ
2pnxL4mYRkFmk2hxJHRWHmL+5Brhxs6Lpbm/onEFfSqIFlutNpbwK2OzKR2imArn
NLrztleQXb+qvYCHM7fJ4hpbPmeKrACg4/1DH0k53kFny5c9BFsoguJurI/e3jYz
RqjEiQqawrN3PBOhRohQgyLl2XFyOtAcOZ6FCgQ87pjzPeZ91adk9s9Zi7WWdEgn
c5ViaDUYFW1VI1WvGzM3RW4I0iRZKLwsMGqh65g+GxrPXrvKaxN/EOdWkKfwnNsm
x6Sf1aT49uZdjcwE/L6aXYwWY4N61t9fOw/fhD4r3JeCm0EbId8RTRTL05bixKco
04bqCiXn4GBY4OgClV/nhOuOingViiMhpe2UNrXYxXAXztq7y7uBzfjl6hR3bafO
SGECxKQRZvyygS+JToMxz6+8qt4lX/Iam5+q6gwzbyqNd8co78xDOws3aMt+NyeR
2wumrceElYVf2VDLZiOr1v1fajmZ8v7Dk6F0Co5Y0PD7PeL4Slm9nGMYkY7qfus0
ErdXaaDiFITzMli4NZvOthQD0J7YKu8MgYxvOJFZa4WHa+zPcGGPtcB0XhQGg5sR
ssV22V60udkqttFZ5VJv+YUP+CzsYoNqM/y5L3WadPWL2y3GMsfzWcavTucOaklO
oq3wQELnUwLmSol3/YlxD9CLhAFidij9igif+ZyLfnmnn0jyY0sPInzCzjPVYv/a
r0mmfvkFy2RZwftXBWGmjni0Fh2QToRY7pqPAmZZ16Tend/dsGSYRkqInsp+ko2a
5u1cxIoPEhknTjeE6CP8V+rwuc8rITFHQ1qUf18zhsOqdFe+XBRN54wALrUPTC38
11IDF0e5XjS6BpSWs0Zpe40HJzkKue++7mP64cg7Q3gsvWdVaBfMSwPmJa7IDfsd
UlZewJt8CJ4ycn7eiCR6shBwRbO/V5ShKTZqO+gzNC5GcigyOl3ZMyVYSmTGE6wk
l6DNNVo0MptVuA9b38QCbDFKFPC0c6R3/zxUuPBaovtJ11mpp+iIXAKH4BXTdTqb
sZJwUiPlw5QHXAsSISSOf1KKmSFg1bM4jRUqBYTW2rnoc41fMQBmtIOm5I4xUQha
8Rkzk+ie8W1NlHwB4szlQNC5dsTSO259UPnbX+3UDW7/ChKHA5DSESZntkVrMHvs
Pa36Np5r2Ws5GlauMSzWQKH/H3ZLJuRIXHY6qlQgsMOb0tAclAKrb/GM79Fs859D
ieg2TKUpBHDI2xtC4TGaG7bHnkElX5oDGd+Nn5lUa7IQhgC5wk45EfR93iw6PHbo
lq2ooUcrIZ/+9lvVGpiOo7/212M8eyyXuTZ2hsGmG5kRUNXb1PCJsDyr61Aqg/ad
mfNxdF0q6TzuDV++OOVw+Qu2OCcxIFXXtdNPSNSrK9iL23iL6a9THBY/8+Y9hpGU
0nwwkEBbX8hozpUyr5W2uO1FyJmjkE5fwII3A40elzh4+2l+FPcar4NH9hW3u0qO
mQBXL2GyrC7/rFcOXBxY8Z3RqupBXN5yXCDVkcpyM+KKDisPMqRuI7BVJa7z58fD
Uot5Od8QGnko4y7ggsy2o2qLuAvyz0kjveKPd7CaoX8zmrgZvqqF3jRy2e+ufy2q
0PIDsfhvvT9iSylYHvGCtxz1luZsnR/V4qKjRy7FzkBSH+xdZYEN3VgCgVJQjZhb
iLftzKCfRiwjF2DthoSv3kUdttpwGtgxaJ/54BMz0iibLhg2h4x86rtcVq3rJz40
tqHKPII1W8uceZAr2iiPA5g/sm+jXC1Us5kQunaiVqm4VdVYkq1VKQjF6riLv4Ff
6b1RUcwXdzfpQezr8lST444U/A8OYqS3rUzITmrd8Jhq1lcuLX2BxR5e3ecNgfJX
2uyE5LJqAsQgloWkZGOR87bHA0hrrw3Bq08hNMCLanU7m9cg/PZELbshdIBJiqL5
qj4dKCluRKJX5E+oEX0nDONeh7x/PCbYaRiAHqA/eDXhjARzK9PootK8qatiaZGz
dCZlu2gjUdcIpTJAGSvFJ+GjWafamg6AzDz0GYrI7H8pen2QKJa6DPgsYqJb9jiO
3xzv18+WhZI9lcEWDzI9B+4WkpUgPPG9CzzMfCgTjRg9ryqt/lOgD6An0b4hP77V
4sNOgwOArfH/iCxdpIX9XL/Sl0MkpypaHXOinDtxWR+0Yle7kdIUrSK43WxG1ClM
f0oYewnHwB1EhZOuJ5BN0JL6eMbF3/mO82Y/H/88wsaY/TfRclBy51xmqrJRnUb9
+5/IPmd4m3bfeUK09MkOoBd92HvDPevDisjY8e1URGrOQQCuyxbsTclFXq44oTEi
6nM0n/LdNRxJ9QEkGSK6vEi8WzcVWUURu58zK7ZtGnvPWM+mXsQMiCVFfD/lgU2k
E7WFQUE+7knNe3Z8kOJQgwTKwt/Z8tds5iPWKKBHUePEdBldSG2UDHO9Hvb9naY/
vKvXqzwmCog6I99xVernTTf9Aaj50uKAgho/KMVqXxH2EXE2NzjISFBEomA6lLhq
Pu58oW+vsHonTOo4Z1EKzNm7o0aiCUoh0eYYpvezbAgl7cjKZJOK2rD/UthRwFlo
p+vAzwr+68uxZHyxzYTT3FNM2OJ8ozufhX8yQhGYNWTWLaR4Y/WR8+2tngf3xSOD
jHOa8g2v3+F+sybLbV3p9cUDr4ztAJm+aw1PD2lL/y72ReYPlJhUBTLx+YPz/yvi
illYup7B/DAnDhLXkvZVtz4w8+8i1azT3aT6KaTn7Kkgz5StmadkIIsIXA1j29yV
1osZ3pAnQGj0MN+NCBRHl6ZJIPk4wV1D1bu7ylNWU6x0o7DqP0XeLuayX4NIoXQK
BEswFnEhE3eOkce3C3wYrxCw1m8sMK9HmmW5/Wm0HLZeLHQ7i37gRs8CiVTDVdG1
BisrQ1rQC2eet7TcS0tDqgB13TvxsaFVujdle5YK0V0QV30uwAswVMk1CcxHsGR3
J23o1rKGoRV4Sa1s0wc3JGpRRVDYJ58q5CYvJzukBqbPpjEDXEZe5KW6riWCUC+j
nyZNcQqwWokB9leVHx5hbR0HcNFZSQ5pocWe7qkBj//+69VQilXhDgDN7RiB69pL
oNc7LrfwNcnaGWDT8AO9ahHKPbTAdPzLPIEP34w98v6sQs2xxvTYY5ES5H+Oz+yL
mWPtivranCHG0N5ycstHHQ3C1Ymv8udI4wOAm4xB22PrIm9BiCf9L+ZTBbuF6MHJ
zTOaV2uO0mvs7Mg9Lg9sdXzVnFWLbTYDsxFSu4j7+KVtQ3TjQdW7C06Qqm70I/Bv
lbKNkSccN+Edc5CqXTEU2nRJY4Ejon9xyG1HNW1gqDSabC5lsaSoAJvtk73ugjup
OdqdRWhhOV50O1Uk0iAek6qILqmThMIsM4MYbfa26cohOaTbeMbSbQ+AdsUVkWRt
32Ghssl+a001uEuf6xb2gXiHH8YomPjYtgYWB3wjW4oc2umX0f9LNwR6LCdOC513
G+LuOWOn7nTO0QXuQwsH8lG9b4Zl7rbJ+7MMPD49lNROi59ZH8qDXEfzCx6l8CZ9
QpZ6uVtetLnTxeWeTsplrVSKpQRW8wvzCbbrSdLFBVHmNZNq8bLiIyI7Kt1jhFIe
99IabTnzd+jmTGug4Sb1jIY4/Fs3i62d5NAUBhEnfbg9zrBDPKtPuS/cEZZFaydg
91LvGDtHPomInnHPRCVEzzJ5ho4ccOROF578mfOePBRd9d+WceIFVNqlMQMfII9r
cUJ/012nZfOz8RQUt9IOa/z/iMWkqeRTApiTsMqPfxg/WVIMgpno0WIbuXHoepnv
zqjg6BJj0rPgyj/+wH5jn6d30HXz4YV2ag5/3CySeu0TTAbpU11Ljav8lvUS2s0N
ReKn6YNLcaxKnmM71oVE0rGNoC6JK1hu9E4Fxl+IntTdah/djHAXHNAlCMrrOih7
ovWtYTXg2gvk9k29KjcvpN0wqf8VcmU/6RvEYtmxEl3YS9+iHCvzAYVKtS1Y5+7g
fLJy08l/lWQaeb4AvZk3KQcu1Uqd0wgM/11ipPAQPSaePRaRbbMfZVpvNj1k1qt2
9Ef9fv+lFDZVwzT6wfsd+R7KMs5/0BiCc9kxfKJLRmBzViNU86jmiYIppve/hSGu
nOkdJNSEyt3tfQOTXwA4Q/XM9e5llpJByrrP4zFttSxVVxA7Cji5WO/wvP/wLnd2
E8w6PXy8BZoKlOIhEF5OTjt+eeAgEdjwwSzNHj1laGtGuA3aPu2QJC0zMFTMAzpo
GAy9S46uJe/p1J3wlsYkSr+UNli2tI5je/UjyvBLbxxH5T81artYdBdHHpCCznaO
+QFjFugssDUK1vubOkZ08m2F8wEZUYUu8f9kcNBrgacMH7L/3YufTWIUWbc40ogX
5oJpa+d4z7E3sKMoVnAOhyaPs2Ef0t1GNWm3TYdpFLRplUx7S6aQr8VlrM7bR1PB
KhX8xEQYi6uvKdXImUkFvGSJTTiTQu4nW2vJuv0xeC+PIj80fQdeypvKkJR+uSso
8RtM9vNjbDTtam+Q/7zlDk3diN8jidYh9QO0cBkhz1H/GNqMpYC99q+UqZkvErpt
WS/rh+fssI2YSPfOioXawHTmr5dLXgsZ68bk7cGkcdxIpQm100IgaGUvr7K2MTDe
UaJ1nSoQdOImlS+Fg6DzavscjD3TcxruyE85o/esER8JAPsU0beqqEQ+S8i4jn3F
/FBxzxmGWaguI97yov2v4xwexzC9OzkF4cWFRJzXXvtXM0r8MMKmcOJSrx7SxtnX
0rifuzd1yEczSXqWHyWWe5pIi4Txxq+x8BOgb+zz4ky5TADLr52ICZw9663K3UVX
x+Rvsz/t9K35r/DfgjjrtuVrPMc1zZf2Xr3FYL3cwZ6sSLsIAtPu8ZGK7vY2+8lu
4CUP5EH8tOUptKlcyH6DRTz8HphPrY1gZN3qv2h1Pd/IGw15rbYLJcriSGl0h8yr
KeyTL6fQM86AgFybmUCWuNjAHzdqeL0b7yLfWm17L/mu0c2/MvQ0n8rjTlLgsaIw
NRTctTZDgT9WhPDYiDx0CFFQoAsoFo0b/EdR5Es1/1MlX+E314sBrfzJDmSYV5LS
UYpbYAOqMsQtGZDD6+1C/VmHChmTFK2fL3CX6NvmQ6vT0RvS2eM4yhXu1ofsyb4c
T4Flhniae4O6e+dUZ7PuYMozIALC1t/Y5av52KVkpBBALWhd8iWvRJDXHxWnFGMT
W8D0a2xpBYzhODrf6x7Mg+ViwIqZqF61GuTTQhzb7EhTY2WwwgbI8S4nMGaN9max
peC2lRUOkayV0oO710WaQALXAAIurO6i6VADBuWEzE0QhEy8JqgPQlaZWpvs2b8q
qJVpZlfSa1dKr1GOamyd+LWgSfXiQBOjJXO79Au+RlgziX2sYdy58kRPsAhlj3GE
el5Qz9HRwRNm+wNE67bduBQHqAGVzcF3eJeKxManrsqPNYXH33J7DL3zTsPxT1yR
bARtreYDcffYJfj0pVJc8Pz6V77Qm3mF/8oFPHYT6v7YIjnTLdPgEs6FiWQtMfGK
LisB+2AAWz+FBlsLSoqA6UYdbdXAwRhD06AV0rMr0JY2cOhCqS+VU9/rROszyzkf
awaZuI18/jS0tWim3WvqHxApngR/ebWaC+WK7G9uNha2j7gJT9LA1cXx2QfntVo2
yWDZCjAju5lBeVII5UD0Dxsuz8tbPLM2UE7pOr0OKP9qrgKXpjGomAnEm6CzOFII
C9JhQHQWFBUvLlkSDSJjiQUJ7B0+oUwz9H+zWz42PSID5ZeRIXeBuJdfbx+E8Kov
gUDQ/fD+FUYmH1SL13S42FX2UGnW35s1Sc5oLY9ch3in4JambJXV4mx3pbpSbCNF
GM5RgvNctKlXXtWJ/y1jra9rF6zWWJrfhjAquhTkdL36lFwj8i1cP4Q/OnhIr8qG
/JC8teu+qSriVznrdB7AtXMlXz+A89nkS3zaG5JxBXhfXbDdUdKP1Atw7YP4D5je
xMIqJY1K+33WmdAch+SBrm196PW9gxUyqV+a2xnGI66OpSAPp99d08EIoo4eZOBa
4eifhmWY7Qv12HhX8hWzyUrnuDdu6dsAKD/LBmiQG9BPyTlEdDpl29KAYxzB041q
422EfHPHbEidh/dFFF27Q7O8GReDSV26LA2Cx6rSmfnX4zqQ5bsd66GWElC9nlc/
yefnfjlsxDS/YdU34V1r0DXugxH9wkNTDx1SNk9xIEkX9lcm2f7gzYEaRu1EkoC5
aXAyKsHJRxSHA/A9/N2sKva7u57VOTuEVWvtSiig7+pladqQ9tolYInnyjsxkFco
JZ4aZWNSLDeyTpFY34D5Gq3aBzn8YwukLJOGy27CiKGtwsCZifsH+19dhMXsfVrP
R1aaXIw0Mxfv9LZ0/D4j3BTA+1nIpOToaiwrf7xPD8WDig2AwMHpy6YXrZUhCfeA
2t/Pmnxiem8OZGk51HshU8Mu5CrCsiJwzeJe8wjDl2T28mWiriDqFuYkjMqog2mf
3l5/dg8NQmF0rYj5N6TX0AFAtMqHJ5cYbmNQepybWYitCzd/jTH9ldPcDp7OEbcV
/QEYRvbcRAomVMI7E0TPooQ+wmtnXnAHEmgxZ2S8nz+l1rbkUKhedyNJG5pf+Mpz
v95VRyL2NXlmyPD9ds+hw8GpAk7mBkfKQUSUYX6JQeXOEr/gy98OgxJLw8lID5oH
PpFJlF7LvWeCzRhR7IgN4WxtrEy41AvmyzSepIIqURh+0THY/eM2jcjy4GC0hlXz
GKQX9TjDpgo3VsIwxi2HP/RriEis8qD1h1TogoZSxqUe2vPjg4l83Gj/ouQNDbt4
nF/B9H02zbx0Id3dMTGkvWFSQke1LRcgaEGufWgIXcIDUyCX8GefnQ74J/MSH+8k
plN79gDDzTTWQ3/2Ym7SdZiH7mPwX2iL2GmwbohCjEOns3t9A/PaquBjL2HzNHwR
PgeBvQfWn1u7XjdaecqsMnRDYHS+/MXi/D4QvnnC5ofe5iESn717qBQ08cMaYUbR
QLrO1J3neCY56gHLofxjctYGQbzHGEUitCWbB3JX2bYNsfl227awCUMe85i1ZJRm
oVVNImWb26ujh+4KBvwi0c3XerYM9B+ZwGctrnz4t0nz6jagDP7MLzowRxdtEqnV
xzanl7CqufZjgFom11zMudkcYKxMzch6MIrfOMOE9x1kYvxtff3wC9005V9x3A0R
MnELxfADkboT75f8ZCbLDRjcM/h/0oxDGoDEz8xcDWmJzra+JwXNdmugf9nP5POQ
2Ci8p3es9Mm6iQ97O2+Fw87fMCIjPFny/XZlqYtbXcAByH9tfpzMycj7pWkedmZc
ksHNdlsCu7dEAiaOZbcqjVLRIBTI7DZeUJnegbJoJuJIK3h83Nal7/K2vsn7S65N
90NlJEveys9PBtk6oqpt00hjLz7BofweOtanPWnQzO3fOS79VEYdSDvBvmiAeiYb
Vc1rHRUVSiffEWEomD8AM6GoXNLj11V8lyjvCHx87oh6UTtsW7Un0lut/aPIfMYE
rEfhN1AFj/Y9YB00iU8dvlI/8wcdvi4FnrWvuKdoZr7fhlNTQgaeFJGoNsHcM0zX
JYYHanUlHrAh44lzNdkpsmGV/CUqE5ztqKcD+gcR71eFA0+MNULm9NbeGKHH727g
eU3pwiJA89V0N0sf1yOje24B+9JQspX1neq70JgcW/THhb6svc1+U6Uu/6LWDXax
HSXqTQi4/T3FIBDj4p0t7Fgf08kx3RnnK7NOaTHnQWMJEvzjGbYbq2j3WfuwaMAx
hmCu71UFRz15qCC+uualUctz+6lkJH3qMDM4EKiF2wbB8TU51GNwRQx6RJWRTlpS
CxPqDoJepksw3QADxQApUcTthUqMvB67zujnk+el1iustG2iBcFw/UTOKhB6Gh8Z
+fBCUv9iu1lFZpSmqqZzfbq7wXKjIoCsGpkE/1h1WdV7KDeqV6mpnyopSHa9gEJX
IJPhsewgoKWOWkupio9prFGCF6PvHw4CRu7MWdKyi9XkKya39DoNViQi9KSx/iwY
elJoDcDskw1BjEaoa2E3RyHwCAKlihhJ7OtENfOw9YRebZ5SD2cLQsfnLGpBg9kG
x6k5qhjruS6HfNuzCMqcQBSWjvfWh8mtXtlbX1T5bKi9DnVGZyC0WBWYlRXuK+Xk
lfsXAnoGor0YQ6PMlLwFTYy/QtpUYJ5atRmeSmtFhSoUwqoNqi3m51Yc1g2SmL5t
TrlNfZrlMYTSgxRtRCeDPTbBtYkoJi4nTcsLAFezPGZKdeJ3EtHrtZu/DVXEcvmI
RUpCq+47YYlsIM6ghX924+KBMmwUJ9IMIRYpkJOtu7n+6HbYFUIukPE7JFor9e/r
BssWeLuDaiMUwHD55dW8Aj2fMmIy+Y4gMrDIjdAEreeNugGCfNrIm2kTuBS0G0rV
aOguHqIdPnF6R5KlSCgcg2EZ4RSIOq3W79FdhRyQ0LE81rdCKPFhHba788guCvP7
bvTCi89ZmQbRNXJQCKyqS0/bQepvaZMenmIyxM7DJ7A4iHjHduvZKHsaufU21GD1
KE22cnMNxGqbsQ/yk2HGhV3eeEaLXLwWFXDMKZjWT14aMOGyndLu5KDCqBZBlerY
2M33vo7l1Q4SVRo5Nj1rwDycGmtrZYGxX+IFbvFPO0zA4Jt8dLlhqojzDAUwN6Mb
eZ0eq6c/ag14Pv0OID6BQn0WVaVCZUKMF7ID/yQAzb4z5fgaMkJU1SKQmKlYdZTY
DXdO5mhq2e4c/sPfhleyZYodLTBtRv9JJK4TNTQ+fZbdCrtZ856HqqNDLV7bfGY0
C9QVrpFAKIQTsMDc8GTYxDOG3sLES/LUuS6TGm61WUCP01pZhihpz0ts/1LcVIwR
1EAxo4GNPlCRybWwwFAvjoNCARVy3chqdSaEbTYuW48z/02pdKHPU6gMrpPEVm2X
e8lnhpQDOu8dkHC+bdJ8o4df1dIoeeEsmt5AalaXVn+aDLWEwOGYpk7nLmFhNbEV
xgtiuswHxsI3Amc6IvH01wU3J4CYM45J6xQFQkgN2a9svnz1fOhxtGQHmvWQNHSZ
KW2t7FTRnvlqvXwMYLQ643U8qqKAHJP/YBSRUWVEwCS9dr+diBOKgSzDCUCaXjTm
2+xM6wLGE2UAUWKRP9U7//nz50VK79zCHSyPtONb8nvgIXwTCFtAYmISKstZg+gS
fCuRlV0aZ3o8SGhCKa1UCkL5WO8rfkb+hcMzHm9X9G5DGqHQH3Tdjr18tQAa6wxF
2bPDgpOh5185v4CNLvNAwuytPzCYNOxQSlCEmG6G02vvpLp5ENH3jnJZXDhf/6VB
G2OIu8kTnQIJ7g3Cc6k8DN9Tjg5DfhH7zHkysyPVwlAOzcXXeezK7Q978qTlYh0k
VT+HziE9MTqjQZ3ks6GNnVDWoRwFh96HuZCiGj00EinzyWPb3WkEIPq+g97UsmMS
Ly/dCfhdS0rG+nG8AGB7ewfyXLP3dsjDaLwwkwkQFksndUuwyRgEJProaVagqvcU
Cf22fzZKb4CzWGw4qb5/g2/mN7bxcjDOlKzEx3fsFV/yhlK3H95B3l3CdluCnMkZ
TUlv0O9ecbbC808LSeZDx03gr+Bt7HWHUs2WDprJUu7ELLp88QqLfFohNfFjzTK2
GL3JVL5qBk+4U8WReH6ZjhGYrIABVA5jbqIKMk1JFL8tgxc96y9ughTXvvBujq23
BqB12yRP25H+Y2sCYlrICzKTs8atObPmOelz7DCnKNWhRR1stShAGxXQ6vU0xhUs
sVlB98gfFaCVTy4O9IwuGKB9B/VJ4EsrhfcmAinoDnmh2TicL0/62giyN0Q46+R7
8/jG/2T0mN84V39QGlgTWUC2dxVaNOkupIPB6kyGNbqhzuZvWXlwW1JL3L4xJwxP
oTWBiOQqkisDrrePLpctexGRLepOvPZaDW2f4Z632eXIxFr1KOtf3JghxWlRT63g
6aPgWva8sFFdtUGTLHfdg/MDfJ6q5EMz46z6aVcY0zYnXU1NpkHpBZql7sMdO8j0
KnFdeorKAjwxwAwrAopIU6bF12qxxXtU49LYsWqTNcIbbrUTSyJojWCK35cNmfG/
kOat+zcoRcYfJcbDEPIbaPFGflOwtaPb267u/UfI3UxFgADzTVbi3AGuwJn5hOL/
YjEAHRhOn9yLyjk4qlqt74cCgqYSCn4xuXCjlzGXP6Te4J1/qOnd7CVWXl7/2iKa
foHLaiL74LpRl+cJPAk/MtUaILL5MphabHF8jwCVAcuqfy/qcOA23WQcBkms4MVo
p47CibejLksP4A1qTJ6E88K0xWI3UzxtkkaemXyGNE8Ltn/byE9pW4y999rp52PU
dwdfljgec33x7tguoiE/57k9EFsktwbXeBLkkWkDa7xnHfz80B2vq3YbXU1vWojw
VwNWBqeCelNXTL1mRoDpFEVzNEayOtjUY8gs3RMY7vS8L/1IUGB1CDpo6mRXtzGC
KpyUKdQ0O0f908nUu7MkVHYkfctUnhEMyyAZsaUJsj1ALeD4PtQmZ0bDTL2tdkrI
p6dLRY+6sLhdAR1GkPNFkiyFmqrr6+TK0xm5S5CkbZXcZ2+jbemCMr1LVbdULN+9
7ylvqiZkK9Sbbq3zoMRJsP8z+LbPJMO78yAKRd3SYjhf2p0fVqtGwN3l1OK3cb5k
N8JoXMmoUhC0pkouDmW6zTwJHFoUVu7K4fdl1sfCpt0BCS3OTe/CY9sUmC6oDYE0
ZGNUa+OFFMG2K3p/oGQ+V134+B0AompTXJkn+Te5aHn+SMO1PjZ6mHz7PeOvuWnR
d8ccX9m1rPg85jwfnE0iOWKZHs3SjUkcdfPnznHneUodOto4ssy1XGEabOYhZ9Bf
wpm/MPWORFSaA5TQdOxj8QOiqDPEEtzsqByW/K4+H/Kub+GGdkMuKvhpbzo1w7KU
Zao6c6cDyFCySG46ZmXJJ3hmLJ7uf9xDQlESDTqgml1dbyAwHNUVY38PbJtv83wX
4zre0JQ7hztAHZA+XIBojHRuIy8F3MszfuDT3WSwF/1RDo4g78xx5WJOdhgS45c7
1Wno+/hHjtjzpe2FVaG/KCSF8Wm0Q0mqtBXsl1qmXT4QsjxJ3uJJh6hFnM4yDqtN
SumE9TpCb6BwGjs4p10n6jjmHmDQjcyClidqU50PFepH4iTGnHvQYy+Ws5AHkf34
/51J0F9oxTGLaSne+FrOy+kRxQeIqSQYFv8ex9S+K+iEZfL37zBpbyITV3388QiD
RiLORJumiAetxBNPnn/OwbL35VWtoykWB7CHMjklL5VHInJrLl9f87i8fwAXGT+z
h4vxMLrMGwwl+sb9CtxlRw66sKAT7sXweCvjWiTcInsiTJbdsrAlFi3FrISCCHSI
pqdcrJ7quhWnF8h5fe1Uu3p+2MedhbRDSrPBopo7aO6YCS81LzQLIRiIJ1hsXrHn
4uayZSZSKBX6W2JcPK00f3kQ5Fr2OGT3U+/88BFaWB/w2gZuymgC3a6CNn9e8avI
QbZhlT+3ORhkCgWzMWY7vnR9Dn0EORhgoSlmex0zJKGTwGrjTg0v+kx+JPyvinJR
80Nju+mv529Gc0rBISZr8utxhkZmXbvIoC9ybvpG9mhIZKpPotVnQmvdIhl0pDYF
gammT12O5/0Eapn6ALIGSloDEunrQbhWsq8SciIGvNiAbKsDUTaMNFWgSRNLOeCs
hOoXTvh5hqe1DkWvq/LhF48t2XHm+wQ+FqrfShieOsyXYtCWYDJbOIBaXXhcCG57
4UeOf/FRRpbRZYvt1UPwt2yqY6mLRwcH5uRdi0iqL12XUBRPB1/eKhklnuiKYyDe
ZBhfQLg50DoyyaYtIXhl3ARPc1dN/ammzzx4NvNOLxkFShtufNPIPqVEMMrLjBu2
xbQklm03yAU9+BYUGbEpEVuXVA182mVSfYp5Ty7SH1HvivH1760b3EODT3V2mxN1
sCq5kRGJooT4Es0FPlJAu0CfKxi+jC+UpDOKd1uaQl1oIYOnGAD/H1n3cVkRgreQ
+dvq0WF7Mxiw9AL6YcshN0+e2tPvDXm+CP5JXgv43zjd50G0hb3TtOJillNvjcTJ
OleWcz37WmewILlOEk6ajIgWPtg1vM7qXjEya6ax/uQstPpmMmeK3AKc/MthijQb
L5e0PbG2sbYmFdowvm+9YXaNPjTDwvrkvDNkJZHUrntIsxse4HjP8KhsPwbkfcEE
ksMyefwehN4qGfXMlyxVqbcHtNlMJSmx/342LHEFH6SbcxcpM6LLGCQSuuuzkuIo
g9jUNfxK/dw4RdRfmLqIRWqgWv5sKeVdmQHcv8oKiky9wWLC3cFmzBnJSiZ58jGJ
Hfljm6bj73GCJPg8xB9gfkt5jJxdmJqZsBevz9+zXa6Fe2iFUKi81C4a++j5XFrD
1Be6EYJ6xRPtySOGBU1M4QcNH6qioT841FVaxq1Orznbfkx/qoQq4zRqM2U6VeGF
oQyL5tf0CLgzixIwBqGkuhpce9H2EaE3/3tORRIBrp+gc1lhYXp7ocqbGTTatOVi
nAurlEUNpcOXStLaHF4BpdfZ6Uc4pxsPoZWyCn7DGO8D/JpZySb6VGXWhnimXbBV
S/Yk1R+ITnQRyBaZ/rtO3IMaBnBHtzD7ePSRjqtMauh2H841GS+6erycAPSJ2MWH
PxLzGAixl8BpGd5YOAukh4AFSZf9zuV9Y3qm9XwHTF5I81OItKChPvaPjiDd9NPc
TDH6xppLEupeZB9FSw03bho9Wdk3hSuVVERdIThleAET+NK+iwmQrdIPX9vkxKC2
hN64yodsHhUaC+dLQyeXInJ8iBd470VBe3I9mavZ20dff9LLfzUKl93M6q7zqpfm
b5x/chdl7oarQqLht+BWK7Qwo05/oL8z6J8781PrhQMw6y7O042D20mrMiArcxjU
xMAmezJjIanHaRwR7JtT64FdY5SpBCss0gKHduUMfgHRV2E4HKdm0dl2+fIkhCwI
hW9yyxiwE3yrYKFVxdW6TL8jLO3NLGsHnOUizQLyYEMweJ6GnazhGwxiUyAb/DRZ
D5Axn+t+++haNgS33BViMTOipxS8114YDlxUSdCaH0GiA/iys+SkqnUDY4zxyosv
0+Rdxaae9goG2MDGgAcYzGgAq3e+QniQOgBBmZCdJzh9jUt5lCZLz14jignNoDZn
fu7Fe3CmYvNZ1c/jE7d/69O7AJ3D1769mKI5YE7S9paQvj7BzJd953RnF5VW01BO
gvbOhAu/zcjOUAtzqQB92QL7i7GVyDs1iNtJ+iEyduFVT0v1atU/ouoRLnkwbOOB
7tiRTGqI4IGhUrK/gGL4aO63YJSRyUFcljJ/AwsKfUWLUL2iPx5AKl4CGZJKUuZM
z8GPMOkvfrlItVUGINkwN6vH3VUjBANdqsk9FOnCSihb415xvsfjjNZyEcp0OUP2
c6syjnIpze4DHYM8aQs+8m1i3E5sKyloSOI1yHodtKRtwsk3MNErOdj5Rfkluyzr
/Re+4Zblq13Da+vzQk2UgwQEfBjEtXbIADVYw/6Dp8pzMpIsT6bQKgsdg9DnFJcp
Y2vhwzxV+AdnXvD/eN/pXPEj7VjAVjP/wYWqcyswByI8CdlyzXOqkoAw3pt3i/XF
xeOXiG30cf90SqdlVFfvnYla/LgXfw2RSuqKRWH4vel1iKzdopzDxGHbO6Jsa3Hf
dCtS6l01aGM8x1qN8HiA0AihMhgkT5f4M6IT6COCD7HjTyTmdLryZsUosKAflnSq
e4XNFz+/KF9LBn4KR1O37HW+kwaW/OxF0TTg+2Xh2yGoluNxKYbcBomvAblCjlwX
ibOOw9VfxCMULmhA5EjnLpBm5cLYUxsrSi64W2rgUnEj3WxjUh2aPGK266ZFU1ZC
FuN00S927pZGsNES3TRNIajzuy50mkRPj+uezQbLupvHalokNm1c3yNfBf9mjG9k
GlsMJlK4+jjT+MFRHoatzWF2jx2jP3iPXAqEXCoCEvgaNb0NGlDcDTK8uLGiASfu
/jBbePtJqYMF8mVWAOvXRMj2LRxxr5b/wr/xujlMOrpvvwdw3Jke173kXd6VehCB
Mlyz4mCFzryu8TBVeV09HlI7j+Wv0ZmSMiJr5FHJFIoVUxkS+NP86Y/u4u7dhVBU
gflYjVv6Vkdywd43prhArGIMXCsSzUurzqQcvOFf8xeIAWVIx6pHbvzj+FCizXrd
4XgUwHbG3iRrSDUYH2dwtQvjBXqH6RZ8Ei8LbAHcQI+N7+7BiHFmHEdoONDHbZgT
o1gvMmn8fsJrqNleSNYua2A7D+kcYJnKOozKun0BXEJ+pYKlwuX0jsmcJBZam/FM
tvet+fRLhd5ak0ZFw2wvBKAARZa8qzNpdH5Km0BBI/OGwlKuhTgYsJ4id95l6PO5
zHlpTw3GdeAMswcwFkutly45lsUKF+R8Hk+U/xeiQNN1j4n5Rv4LqFYasuEDQ3fl
iKHKHWw5AuXCdFRlqFixwEM79AUlER5pWx5dsEtCSOXpbol+UoSwG2OE21jg0cDF
uvAmD1ZdTBMejPwCWLMOMf9S2BJy0921o55t+z4JIk3Zbxg1PaJEIKY5F5V9Ob60
DQsEvqyTJaaXM3VfWYBrtA2rvl+5esLTiAmRbyRcreczBTLmhJBeyjmPTpdiAF41
C1aeNbDAjIroCM0I4ocdbvFQLIV6qLsp6Iz5Gy6Jzt1qoVMC9oT4rG58cjn3tH/k
zDUpamceiTgpfExsXnsfwxlloXbYOrnD0vWhDV4QmsI3VB0+6P9vUpNpTMv/yipw
TLzomMHJ2LIcQLFbEeEg97S4vBsAAe6egxGVFiTNM8YeyX+TcRpCS+zHpIzI/WIh
IeblTfDfnQH6NJnv6ZYqMzSFxSDpmWqmdncLkYVV3aXwyUs0kuR0lECV4Q/EQqnM
SrU5pVQnebY6gAAaAXepeEP8qFdzwfIGucGu3kVvXuXLyAKxDEeHKuQ+ilZfedW+
ml2WjolSkxFMduYEZZf/vMCix9oLNJKfJiZVnOyQRW0rDHvV7GyB3fPnFslbVx5O
IG/OP75kviPu0B2qfNGbvth28xFsZkWLN65iycJMNUozDvNxtBXhJPbCVOzXNTdt
d5wXO8Q/AL4kCKwb3k4X9wR3dAblSDnpUduo/7QHX9IQu3nCbI4SIJq492r/QoMx
KjAoYn+ljC1i+8mXNe5bFlr13bBvytA8eYqP4nAKVixL+CMddU4k8881U5bD+5w6
etAjiEJrg7mcWTZkf/2HYTEwlroxspJNDcx/a+bpCSDXA4sfmu1r/xEWn8v9Wfo1
DkW+ED6u01Qr2NTE0b/yerwGMGQ3fEF1/evmf+6zRq5PswmNJFPgclVB/SWFjVJA
PfZkGxbzU0UtRxWKCugs/PUAQ0tCc5H3JS85gxVZFO1qg+SiCFA47Coy7UYn+k/y
k65bK4RQLJ8y7jyc1vPc5nlnerkwv2wKi0Rd9n/WVJ7LowIQvdOmsEdO8X3Q1xFV
ncGCm/6tj4VwBBW7n/kB0zjwWb0awEqUc3zn0aR87c0i4ZLiqXN9JOPvte8jlsZ0
G3BDRkmyVbIz4CsPc2zAdF7/HlVDHC2oreuC93MJD0x7Ldg2KQ5y/WTVdXy7dXlb
uVUZ309KAqOAwEsYsXdQtpAghnbHp3L3V+rwL5j+u9M4rNMmLJ0j3s+0fO8oJCO1
9bqTmFWUgxWJr8GvKB9TFqMnjJKoRhRT+MpRYD9tWqbDAygSL03gq3SwA3a5EdT0
slC9RSnyiyurHeqvJIPLuclCp9pwSqJte5qYZtUkRLfKw9vpcyPMyzkepedjBryT
eVs80FMEVpbEJlUDGD1Y1hFrxPaywjMMINT/DOL+/1UufklDeCMWl63JmXl+ocox
1xjNFykZKzJdLAy3WabDYT1cKgPwbVF1TQKyKso+OUTwabCQB7TjKxYqG0zJnoWe
XrTrpAXvdbhX+nU/imBzQ8cZc7s3dS7l/gp1UwHq3Firu+ejNHT5J/5UI+5Br669
42QTzFyBVtCM5XdsrKcS/hyX5c+ffHv+59rSrsUuyQSowugLlVJdiVJP7TRl5abP
nN3+0sm1dZhU6GEpPCVsbdUzwiaFQdEzKaCEjnhDnNgoeiFc2D4TCPya1+Imb3hF
UZcFQH9gv5JdOrfbuQWI+sWWETy8AmDhjykBNzRhVbYzha3Ff+bnLGAqnHBvr0Jm
f/bpM8iV/GwTd305Kzmdod6ku+owyPNz7BzI7p/9SxqQpAig+XiAnp4h9Y+orXWJ
RbOMVxVkklEV+KSUm2MAuWxSQlIsH3iGny+stDMgovJWYl7isBmaCRt76N6D3dmX
Ww9uHGyOqQ/UbxzVmb+4ZYY4V9SuWPSTwS5E2qcnZ6FloNiLsI9oFS2nzTV2K1AJ
i0ni493hwca9ya6XetAMfHzfMserqMP6Hw1YeabDxOdlguK89ZfU9XBtHh/IQFLn
6GI8/ALgKhwXQrWiP5dS/4W2peD8vIaCEwusvwksLlwqDCa5n3Q3WojaaL4gGICd
1M+bPzZGoTjTj4LTBOfJvZkXct6jmif+hJhe4ywcZHjmzBoE4OS89dtfLnpsxTZZ
b9ZBmh4v9iPMT8YN1OjMeKlzy7VPcb3Rty84dfdzK/7vx23/udnCPQMGD7UkucB1
yximq0TDmCb/nAJsGyCfRTdwavR7gBUh30rw2Q/Dsx0yNThFl3RsasaZVmPWo+Lq
Vpq4uJSIoXRKsFlgeDPCVYLRKVk922+sl2aqCKFnZ6veQeKS2YoYQsyqwswfpzFL
9cNpt8Qw7Qp2VX+MJgYBE2yCFmW6nDwDFsw9Tai7Rti3wGNuqsUvB4RqLplKRQaJ
km4+a1SpPLg0akMhoU7JE0H8TXX6QHPKpIdbfs2pSQa3HmaqWJWzGL26rEeR8v94
IjEhQ8C1Edib1dAqnrCN2uANs7GZS6KV/6k4MN2jp5n4xvOZmL/0mN+rDGm6JNe2
H1BQ3vluQ5dIZsHsk9bV1kyvwp37pOFl6n+llSiphSnloecrWOLOgNsy4O2Tpb3l
4qi7swky0IK8x1r2A7jM/WO1ItueKjanTyck04I4Qm3kB/d18gU1AqWkT/CNncXM
UcJHL28H4HSah8LpJIOpYtye/RvNiMe0C8A4x529hj0ubaXPeQ04LLP9fbCBM+9R
2uYMqtva/kpVoar0AMOTPn0T0TEi3NFxpLog3SNgsWjxaxnW64f6JgyoZW7lJ2F7
4VEKZPZBUR/PqdYin60DHkDSXQxOILG4Dce4VRmkhpsCBPU5Klr3Ca/A7Sln1Q+5
+1X2hc5u742NhRIJqZgICavass3vRJ8fegKp/kJ660N3G3qVgipAidFH91VJO2LW
G6bCD/oMvPNm4uveWEAwCXDON5mthjiD6LAqhkeTIw5Y5mWMIX+MfkZL6JOhpdRc
iiRpQHdfnQzU6l0wAXmJSJE1v9HpslFkD36fAA+6QwYm0YwUxqIpAai6orVPm0HH
xGsZ9OGfO6ShrqDi+vr/b34y2fq8TvpHwW5Y4PJpcl+m5FpwaKcHQkdonvjFOjbt
155Q80jM2liqOR1RvRvB/ZdbzQjMRpqMOlUVnsI/LPxAuEF3p2WXFoLiQGMnts8v
H7X760ZtU0X0s1qaIj1vDHG6SC51uozWLhH2cfIAAmZmoOkX7Yl4/1CeQtNnisJM
vBiFrAOkWA6MlPuUwaTPkSXLAhVXhsit1PT09GGQ6RgMg/3KTiCGO1/FTS0sqhO7
Zp9KjfKmpsaaeRCONueCrYHGT+ROkcqTrES0eUza0ItkGJH1yPuGrJcOtNQodCWy
htsnIEKex7G1EOoaugJN85JOxNS+TX2xr0lnPbHf8DugTvxb1aUd07oPb8m9wTM4
uTp2EQyX42JMVFhb1rlUT/jn5vnRpFD+dpZmD9RtvJPnqcizAeWbgbLrpTTxVMY8
2w96gxkwNce0qypHpUfnRnuoNeiy58F5RSbKo/YgR8Wh40KBT6ejXfpXLuQloSA8
Nd6ODcCwjBzZ6uArRw5E7qo0oJmsH+p3Ir1UW/3O03mXf428LSUbrUosDbnPX5a4
ZPacH+YzD+z4GE+AgzuhX6qy5eKrYLh7aQgDiEpb9tm76Vu0+h0HxhkNVIiRfUa7
9Lc6o0jEzlg3R5lF8UfjHvZ+rojfXNLmmCb6P4rNjgwXLhP5uV5SonCc4aY7bZZV
vkxXR5mvme/xWbBq3oNyZGhnMeVwcwjGiauWIDYOYsgDblMTJMkp1xKqTixSyEwl
WVqVab9n+XtLb0PTWCQIyLZZRovEyUlqMxigJGAQMasuq/1s7J2zNJSO11karBpy
R0qZT9s1eqHB039JOBGCot6bvzi/bLW6C4T3AaxukS51OgezP8Zu9HjJDR7i0Vz2
LO8cOhQJN6V0PyjGNm2iEfkwnhAGAZ+CRzkY5WkkVnJWaVjCEAUqw20ewCi9rxi7
K35xhq/dHe3xCg+hmuZoa7DeuDEWgWIq4bpSQrc7SO6AqgPIiMICvtLj8qER1/qS
KpeFuWeUjYId/79pxw2FY/peCyxF869UDFezTaQMGYKn7lHpyeOH32Zjtf8jlN6n
XF2LpRtGXQSCyiRVevoqePASz01FpLXnVEOjYY8Wp8CaDTA4rM+gzDNNu0BBDNUE
egZ+3uf536RHRXKVEOxFS9vwuDa1tQREoxLFdNLyx1ZTnnaMeYD+ohgmOk1s/O/Q
RelEY5JDU0vACNYwReqQArUS+l3P0iIGJk3Gg6fZ+Uxg+aUh+a6BVxU/boyWPAqA
WIaDnzLiPdR9vzxjxdi1gt019ty2XbqoZnUED8KaRKrXNntg/bMx7y/ZX0z74Cba
9PIhhxawEogHJLLR6uA0jvtnDtUSoHWvz8wiABkGuRcXav3gAIeQKoSkgPOPhk11
O2LCGPdvWOaf4T9v4Pgs4HR8TTocukaFkntNSqi+rDIYt1WaUd14S0vFdrl1qG5x
jkK1mynPHpCgCEkEdBgL6tYqV6GjOrybq6o5DNpeS8e/intjs0OCYIKBMkzAWntP
/h4IjiqI0rMuF7nvJMaWKlgonPLosmVkQui3+j3CHOyVLI3ETlACHs1MmO3CFxLW
V40ipUFebxStiXQB6XLtacTUIchgVcWgZWqZEsFoUR8tT+jnKU3PDZPmj1q/xk8a
BAUt8qmAGpG4I17YeWk3A8lcAzEW8WvEl4JWS8/DFtmAncl//PV9zDYw3QHCVIkh
fV/A6GMhwE8N6M/ybDTfhQX6K3wWIkfaKhqJcoIab7X5dcbo61fVfiNSrJU9jyeB
UYXj/lDT2vbcSGkzg7B+ptakkxII3D/jp4jQ649jcEb1nz4KM3VTq/BEEXoGT3ZH
ludM/RSMjihVQwMr+iOfpeFlBf69WJzZCi3Hz7qyGWaO/F3a3X+TXsFr1dhO9cVp
qkUUciswQMK3ij/TEbHa3SuGTJS8liuIZLA2/kZhDydKHPrjZ8bqpsIj8ZR+EWbF
grP/I9qEbOwyAlv3ixq1q017rnMfOY0BDS2YzmIoHcVsHiCO+n1Wd5VaobxKGMiL
GRDh1KiFYOmV6xBa1n1BNc8e5VXq6X8VXJoVkSeshs+iz2FIlbkkUrRmHo6BPJEG
jN+QLt5A++t2oAp0Gj4i/H+hobppn5hQWSvZEGxIpfprSlc5htvcKsnyGK/a+usC
5gp+6QqVBAC99iuxSR9h3tVve3IdWZBgCfBeJxjiPL9XD98pr1L7Rh2IPzlvP+s0
AiUXHCi95FR5Bo3QlJWMj9xnHPKqf5q6nIssWV6VQoAdT+xO00obTtB3ttcWFdem
GzgCrPT6Tq3GrBf5aPfPpJzwy13sHNJTWZ7cVk8hzmyFmPvmLGZlfw+PLsQ+56AG
hzslF7XdY5Ptr7EDGxpf6kXN9ycDcjiyAvDQcVC9ovxZ8LbroPzzJhIc/ZC1TQsI
z0Py/PCvM9ft3J66mMqnScHjck3u0kEII9HQlFEvyLn7l3TR2efbknPNHMmQ5O5M
rLjwVGxaDbcbEmITvyeIEP0UZaYMnUySzvRxvrJOZ363lCvv/lBwGWy4DGg9KG4m
/jBq8uZKYMSJNcYSfaji4UGrknKbgXQVP2S2A2LOTYm9NeACHjiuojSlySTCX7re
LBoWxK6GC4Acj/IvBbygN4ZXGtSkTq5Af4T2V0D0ouEs1e3Y669Dn4TRmn0Yisk3
PxJ/ozuiNkB+ANVbN68WIQiSblymQMRNj6XqrKnAvKC6MzDMPnmRh7dXV6YANhlf
cwtguX3zh4xhU6xqlTWfxR35vrCcTNXVk87HQDTKzYUgt3D2crFhI1EqlsupOgDu
D4yAiFsIRp5CD5oZ8XZTWl/K0ZH6L4i24tnaZ26J1lrQIqGSm0ukZIuIZ6E6mtIE
4ywXKswPGRNidZDJcLnA/y47DV6lNQ4dAP237jZsPLnsCleGUIuAR0wVSQYhxxt1
2v70/5QogyqhRZAD/vHcod8aD58Q8JaZXddv+304+KRQxXOEfg4o4zA13bLrZVya
RTOPLuT+kvtcUjtUweeh2kQHxTEXEANBXUESk3XMUgp7B5v22D7K6qayu4WULD7U
phmpH9d+xTZ34HsTZdAeZ7Dcuqr1+b9zbjTsbIbkKM+jfRYgX8uTyX3948LHO7h0
glS9BkhQog3l1qijy0tpgEOkxPugZcpC9gQXceydzn3s5NjjotMglybHZpBYIV0O
7WeQB5SlE8w7IcnIX5RAi6IlmujU4o73xfaobpjYn8epO63u3+cusyCYF3+lBImD
lVNizQt7De2D3xrRVCGsRhy03mR7fFoVytkVGXZSCzMzN5bcKyx6S9IZqOyyDIcI
+zUI7TTdbiPwg46to/nI8vuoo24xQNdm74pgBfNfpZMxFwnDXCE9raeXDg28pewr
+RzCRxBzkwZnHYqacy75lxd/9QOloNiGmw89fRjC3NZ61P0R2uk1L7gjF2XHb79S
n3xEB147dVGsW3jHPw1/0nwcrj5dglDQdjhSJOuJ/lFCOnMWDGYrKwW8a+2LBLI6
EFL3YnLefQceXpxMCvG7yex+65JkoHIWZ9emTZkR2NpfFgYSgsXqO3/elzLz4DrL
VvXTIpok0htvFPGxcWleOpaKcypWXZIbP5RLU4XQu60R6U6BNxA9FwqVVEmLzPV6
ga9ZpSOW+jLa07hy0vbhvLOMfJHkmd/BzxOcsNJ10ePLDLHvcEVBjACdLJV2Epdb
jeoZ823bGz2e0Hyl3aFV4s6PErnGjCL45j82uFQE0+06RW83QB94mdlGw9/P3WF7
WXE3RizxvL2q+q0UYX7QFT/5R0jOZMnN9+h2NgR26OSmQxPerKhj4H0u3+oAtFju
HgGe4S3SDGsK7DqvjjEHejgNH/z5dyVvTi3ehUMwu54T8LI3eUTOdAPAIO+iPHA1
1HXt3ri+AgcCv9UcolDjd0P9dAiC+1ZLrIwPc6scFBbtixNzhwA779scUH1Gr2an
ZBnegN/k1fCkZCtrSBvBz4s9kk3OE0JmyZiKEX+i4rreSNr3OkMK9vET7hH2N6jU
WHYAnT0CQRR9chrL6V7RG7sBOMQYjqmAOKWEX688xzIMape/gXRGrNTZfqzlWw80
annVA2kQQjbciOIZgNhnweiX+Yt9dJSNZ2FaSBdf7m7i5/8TUUEd8HS4H5Myoy9W
UlceSCUr1IHF1MFNVVRlAbmzUT/0PAsXkjQmK0V0aMT1AwCbUMECfmy0Jaa4hClx
yNvKwJ4G+DbqVn16lbWF3La/Qt9wq2vTyi23z0UcGpI5nCmaK3/jg2KkCc369wlx
4iEJXc7xm346i4kPqR1bbdNl7EPVJAUhMDMBe8RNmW7cUwjkw8GeKr3oE2wZQtu4
d0NvDr5ItnR3C/MqpyzVBXLkaTCFAzaQfPdoj9Z/hPffuM2olso5rf7qJhJTCMIT
xauXUPAMHhgdGW5FRl4zS8ns0krzaaTDyAz9Wgyw1d/+nM7kN750e58dAbj+gWqs
rwPhMKQlO9b4GfeUiJSt96uhsIygGf2wB2q+J1PKiRvzSZT7RQDD00fsYV3LfJ1t
wRR3HO4iuqizmR01Ol34SjZ9mqGTOUkuAunGIXvteEoWrv8pBRWCtQyFg9QfynVS
OIucgrYwj8jrOxLlbLUH4NVGpsvyLS3l/1/jS/ZmiV9DiQfWnlCcU6/KIAXSrMJb
yMDQrCD6LdH/mb6k391v334M9aj4TlZHCiNOfoN2sm6Uzzrc5Y0NSX4aEwoBF4tB
Pjy7cAb5GlcaTtkrFJwh9Zr0D/n6YwhW6jOYGZnLF/IymmMClKz4A4KnbYDQPCkp
EKpf3EhaIIhPN3ocTRpKAfggwztzMV/Hh69ifm25CPJHIQ/li4enuzEc5NyEUhcD
XuCbZrFJJKvwsKWz78fVKbgSsI0Pbe7akOL8hwA8foj8WRGlHfRRsL0Uk1oWr1ka
riM3fOlkt4A9dmJ9g2dzp4R4fxcnF7rhKTYXDJmTtMKcOS/Ra3hKnXeugm6ZgSah
hJxCt7ZX8Gzx9lx5PWVQIVLly9KjE0bjkVrsAdr4vI8IsSdUHrVwl8XYsXIeHMmC
MgUNG9RP+notcGLh+uUOa2Z+KihhPouzqAkpLhiGNFRJya0F6aRbFmHLvEFW6N7M
r374/6B0tYDJJwwl0MMDHidIf2d2DZIxzVzdJTpD9FlUa5HpvR/Rb47sKjE4bTEn
CwSsCZuCfUYJiLXH/Sd2NzY5U1U+vms5nX/I6PBbriIteb8Fz8eL2WbIQP+cvdky
SPko2bN4HBoNwacDvlGDX5uqCWGw/L/2ilGCofDG8pH0zsQ4oxacyzyyOnwCDEEj
sN2FBxM74JFQhsXpAPg220EcOTrA0pOAjYvxRdGQqh1o5KV8zdZYjWhaIT1Cadjp
auqStO0kfnG8cD9sj8tBBc00M49a6KetSVN7k4/gp6/7jcy0L/JUTlwQon/0wRYo
I7kSRMsB0x5cWs0yynlPlfz3JKEKxtinfqOh4hSC89B+eJ8h2WMBVWibSb+o//nA
iV4CH4YfJzbKrhcrJrCljEkv8zfRIOeuS6G0BL3iSxGch5HesFzIHf2X1/V9/+dm
qiSI4jlu0Y/BzRP0mghpIzLyDrjL5Fw6wv8A79DsLGQxwqwepbX9HGYRspEEaPvy
3l3Z2iWWrpaAMPbcTWNpM6yygwkFkJjFHj0KpLAjpykarZH/tfEZ5oETF6pOJ/Fz
SSTnuRo7ZM7wgLawnOrZDNrm663+3WftpCeI4UA9/5iKo24dkYTkyUDIThuI0Ale
oFZ9iCb+J9MSsOWirNCB3vhV1w8yN9gAfN2FnBhH3XTonSPzWNWvMucGm+6B1tyW
KZlBf/tTehvnWTr06GuXbjCt0QJOMU++ptAhsTFWVZCiZaFtEh3vrrPMK7fZCIcI
mk+/UqP/ZsGpHj0caiOg1zVIjMFCyrrs9OdvRpuhNXd3pIKCf0NgzcVmSnMQ6Dnk
fy/USqmLbaqhb79F1o5sy9itcEUS+t8sfGgwpk0NEL6stOVfhzsrwrHjRVh8wLxT
V5UN8VzIKzarVc6JPBF9qNbwaajCjU6zBnofbE82YELSP+DqRmpfgv7mIYvkQLoK
mDFu2dwVnYh67K6Oc14jTJdGQxljTpB1YVe4H6mS+b68TINqyk6SpzIAtpQe5Vq2
A75QDCAVeRhpUryijxlimoSfhoW32zhYNej5jNjEcdQV8Bp94aYgz232w/O6JP2C
r6YNy5tqPtd5wsOdB1gNtOSDPSxk+5MuUAXaQ6DglenM1JHCjmEQ7tX/Kx1zFF1U
lOk7z/+wafB74IhHSJ6z6HSMtWl0FvqMwe9M1WJyT6c+s+Dyve9inkKmZIh6REYD
4GbavxIsEKbEXvoGFKDqKv2Q5KPURAVp/HrqP86lQtmFE+NpEA4TglFbu9JWxpfz
BMXd4XYxgMO1IyZPHsuOrc21YMsEQefMWe4iiGEDvFnyZMNnE3UmSeFgl1XUrMzx
+3EAgdf1c/tP9cs4P9vQe/OBvKMDhK2sLUxA3RIbumwFJ42f1RkXT7ry8SR9uxt7
QyhguS7dhZFq6Jkqjl1MtQbus0HQ5L0eUSZEQ/dBO5Sm7qAj3mxpwaukXl5vSSZN
wbE+dOSz97qW/+W34I+mwmGU707yuqosN2cfaZZnzZpDCVQjLFcOmv85jFikiwhL
ZUMth69kT/eJNmUXbTpsePex08FNYzfohP6xJ1hNjyGCFAwt51YK1H+/xpf//TuJ
yg7mKmgVEYAzQDnBpfwUK/rDJaTn7SJUDH8NVOvtwe0cX1MDiHTF4cf7q0OtMY6H
mBy34zpBliWV6nfbfyna/QC11SFxZqhyF1UO534h6Ug+RAclGusAf580DUwmzTaF
c7lzijdDKvfpLpb+umbQyo5VO2/PjZcpDbw1tOUvAlfRdrwkJwvR6+Dh0idiNY2B
E5xDLZSGR+cc4vaOksE5E2cOH/xf5awt5t8gPdTOFmvvRxvqngAdZeWZosGaE36f
JMa3yEhaiaLoprJcC6dh15JlHhGy5cyJ1xnHDRuM7ibeKElmTVFBFxzK9McZI5Sp
Jypfc5gSJ6uwoaDsZ8VNdt6PRIPSGLK+kzQEqNPDPyfoH70YjqOoO5c3Clk4t539
gMR5WExwu88Xt+8ehsIB5ug+MIy1QkfGyriaP6D602jeeWaHd+sTQZStkoDyzdHV
ZXhNVSkNf0Jb4Zwww0JDm02Vq9cdZ4w6g5qPBI2/QBRVlRAP3fm1u9p/1m+w0uHA
MgaLVt7X+GBaeVVYeB4UeVfVAUkcvLS/7CsZfuLjjq1Tgw5sUhN1DMTFJiijcLvo
rI3bxda8dYvUOSLsjs4waU4LSD3ka+zz7Jd8wnMLFAaTkG38tgaBSoKMNRfBaft8
pcXqUF7xQ9mQy7aoG8r48yynB8CzimWaIbXi8HXvSkpUTPuPxaWnQawr8ga9IH+T
qo5yAbywD+7srVG5P9BOKFsZ3kiobNG9SiluDdbWkG7C+B/KsnyvjzKoRFVKuIKO
MViX24DYYmggo6yz2rSiioprswmBNHkqbstkwFziZ/H9/Qi2GD8SygFdhNCR4Y7V
2rfsnGmAj19Z1sjz4Id3S5n33sQ7uCc4LQioppOKf2Puovr+vZnusfuLhgB1FZdl
84gpItz8uGvXrcf0CJv+qeyx1rS1WY06mT+Ua7YsH+xoZq8kLn84HOcOpyY6pElV
t76Y2MKHr0vjaGF22sZWKIoMKq4EGTH/mhWPxQLXpDLunYccDKLC5NYO35dyqgOk
nzmZ1kFN92fFERAKVziGI4yCn3RqTkQ3M/aSweLJzs7ZAhoDX4DgZYgONFnotejC
N3xt4pwoegKrzdpYex2bsE7H+bfC2MKRhzyGC8Rf9vBWAp+uCBerdjKNLSde50ei
1sqshf2hargU2IK3Qu+B5YcVpJF5f5ZWSYVGTjSp9jw4cANmLllvYGsNxbsLRsCT
Nz8Mw4spsWfNzjmkNEreGDimvGimr9uvT0vvvJqx3upccEKBxeShO7Xm0swjDIzl
M9UoRvqHkZPLSsua0BdVfI3BOLrhhIQ0qoIAjBop8cAkuWxf8yGn43LtgX/8dUUt
UsQqTzmoQJwDq0l0X8vOkZBPnmY68Oonwk2njoe5m0OaGyTp6uOBI3PmseLOv7yY
H9oV/1ZoBM/CdZ0rlgBy9tOkA5aMo6xIcJXTU9yrxglM/GnBom/wVPcUcvqHUdnk
u+BU/1dazT+nUzWV5wVrFIxpbXeBLD1KIkQhTQWkjsDeX9sbEXPEn2hLXBVSe9+d
H0f81sAHQHRJ4qAhfsDLvwf9pTbvEUYDhVUNMtRlCEKdxwr+6GaspBbwJZa2Kl8W
S9ZqpLeQRol9bMryw7GF/4o5nuiRMEZWF0RgEbl2UTIjWWgtyeAEhtMmJR2lZTxh
FBh4BSEHTs10ahiziaUCs/LtY2mVHAOOkvjPwRFXBXsXJ4R9f8zKh/QQ1LrnaGde
Bc2qy1Sy8Lw+F3I6Pv9Gsat9R0wKS5T2nA7Wcc9gqrUUPRuYq6h2bqPBnMENNAme
/NRBFaPML4oQWYPapVtiSl+wcMtlH6kPqYe516hdIyx1rzcqv6YDzXHAJ4PVK48C
avQ5OA2tl/Bz/IzSdxZokN8oxtvdqVlJx06YlXY1+g3eBk6wbPm/2hIt1oePhNbQ
CbDmVVeOadgPXiKwo5vJanHn97ePJKsE8XSKG8u1ixSIzzvMjPCOja9QWmY+VYOm
eMbHljjFcX93tYxqkWP4wY7j0m28QrYXLIrTuI+S8azD6dDxbDiqFm5J9UZLuhau
wCccqwx3m54zAmVabXwNAY4y93A0yZx2QMqRLE1bR+hc7tQq2Eu0VhMMBJFqa/+S
JdFJ4qzfZ3i7IiIPCBjS7z8xCSnCEJQqdkZP788H7/VEv/uggHYdDieRzqJuQ+Tn
IqiQNAZHFQ4EDx8+N/37z7SFTLTuZx3DGcZwbsiwf6QIi5nx8vH3JMc9jweE22bU
88MXsu7V0IwY/gtm1yPJ440VRhr/gIzzIyOrSg0HDPo0E43XdWzHHRwmeKcDg2bA
P1MDuWflA873aKBih4ir9Xwi2fRP1DtOy/as7NdkLaKOsnybCkC6ie6ui0f4VxlG
h+QPQT/upq3c1NPBKaEO0sA/8EOyBryBISSqlrEfOm5nTglQsf2lBBmyYjYinK2+
YkI5rjASe3G7iMsxwNZf39cYfO/NbMascDRq3BJzrKwKz9UPr5k4oW5kDdp68g4/
go7Tn9AA/CULhcRoUc08zzUvNAo1NjelLDY6Lw1/j+NihcR+E7tHSes4gffkh8Sf
fmO98RbihMAKTMdLM9yPpbWX1mqwNoz/FOp6mYZV6Q/i+IqIgaUlpZbjuk/bZmLS
6qArRGiVl7UOE3EZoCjqguqg2sYM8gE6fjjTtzPfMnSVpIyJjKxgBuQu+eoQ5uDA
0HPUdPABgHhKox/+1YVaLuXC8qPk7jEYkVJV0Trn7scsL9LGVfsrPodo40It9pXF
tZ6j8Ae1TOIWZkHr0Zp850tMakuiDQWmhKVlwqxpxLzei7UwstEkM3pZZcK3ZR79
NpeMQ7lCr06jnw85Ltp8PhDX9pzy2fGpRMEyAkdwi7UHOQAkRqihgx9Hvz4Ays4C
esH+dyPY1gjWpxpe0iLmWoTT38avNVuJPdDHUCsLBAIiXti96of/RL7eUAVJx4pt
HalkIq20II0//44VPdyjBhK3bHMU78und1s0gmbF06m55UYx05De80QjfgXA3b8i
15L15YrOQ8jfkqv/OsobI4Z14UERZELaU6SnI35cxdKlKOXZxB/97qgmyVtL0Eip
W1CRHLe2hK2hrL+2BdawlShlyI8Oz6WC1g3DvzfI1mr4hEfHmCyIQpazPDdc76o6
Q8G+kgCTZly5VKbZFDHT4ZPgkJmW0g5zu2w5BjAo7enFL2GQPmsaidVnnEz7FVII
ZI17KDbaqt4/8xdQ1tnhyrgr3372QlKiBPvd3eVCEPWXM6T7kJ9OeCr4Rm5FUDxP
oJ5Mm9Qj09AJ65l3dHuaWYyXvweA9Xh8gttB5UP3dZ2rJS0P49z2poR77D82e+JE
7rEAdzvb9FXWQ2fBnmyE3iVTqs+6A3PEo2+7n3mG4hiLMKJ9ymkCirF/RpMT9gjs
qCdM2DQXql+nmA6psBiWoED0sQReS6BnOz6bcWGExjJ6Hlb/95eepaE+eEwhnwvi
adb1QZptAWH7Vrueybhygj0K51ag2Q+xh+vDQJLZPF9HSI4zDm/4Z2nga8acM+l2
EKWz4zlCsZgoVEDz4o1De+kaW4b4vqisN5l22mhatd6BXCcWoeegUa+fJdXqwUkT
BAsS89fATrv7Py8v4XEmMInZIr8j28G/SNTHT/mdThMxSlm+tXpPdOY93DJxQT/Q
+VNE/r5KLSefazcIs6v3kjx6sRlzl279PrVcaCy3rsKd3okkai5+DAZkBgzwdZa2
cJFqH2EXjRR3uyBRmErXzAqQs+JQ/nt3WLbuVD7j4mCtAMDdqjwtHPhjLKNHLF2b
6Vl8LGqY67XnuK1KHJjeo9rRGLxSerSLZeJ8aSV/zFEF3bKaMA5qKuckEFnWxG/G
7o607DmPJ7X/Qa4iW234rstOcfB8DLtg9oXJ7goHBPsZQSWMtWfh5suPRhkloA0y
ltmdWe3Xt3XxUQfMBOGw2HZLfkc0RRIOBiTyVjNKEwNcv9w3cupzorx1lEj0uigP
mdHz43KF/jR0JulvJQB2WUwmR8+mCnyGuIrj3vNGollqGfW2qtSqa6vtucOX0PE0
68sTtB6/cjmCKavfDvMrnjXE4OJGVLdGsr+nXz7vvy1rUgQXyDdazdJ9eMQtb3N3
UJgUZnx7dAfHRDMAsaGBUTRBULngXTvbnlZ4hKCATIDp2kyFs2LXvSe6GsTMAeYL
hKpsLLQIR+FsIM74Lz6qTL7YPga8v6zVigcM9b8mwB/Gh4VUOiJhrxFPXK+ycHe/
8TPLVxG1U2vIzfiCBNa3NKHIT0tzVCLEcAiADuOhWqil9N96cExwEJA5YaZz60ZF
QXjMLVniSe5A7D9+7TdFaCQETchze0TVoo2j4Y5dV9i0CjAfFPkym41daxP4Y3JL
jYhnF/gctqqiYIR+/hs4Bc27fgwiAMpfOGy0fjhLJUTYO3pusFcgXFkfRpsTo76z
klUz+UcXFQTtBJ62pj5CyAhc0W5LzhdyulLxttq5SLK86Ka747nTexhxCAFSVWPm
LerUn+4CEc8YZ0jMzfZN9O7DGf14Sh0PZvi9Q9cRsep8dW3dxET3uNhiz4O7nTVD
G3aBwGVBq8XXS6EBCNR08p0MWEf51fLyYtWw3tHezfTDcbe7mIrc9hXvT2umzzmN
m7ccKrIVTuLIR/l+W/uc8eJCVOITtu8usfGBRB7EXdNxrW3Ml1+nzPbO8t85P/ap
qWTDo+zSrNp73fKdiihxn3UGQewNUbfCSZae1wSNV9wdFYrK7TsSQT5Bl8L/aeAf
Shza69XJVpTI498ct20ajTHZ7kz+JGzhoz9cfZN+U5buI4YvfkPkx2GBYe3I7JVG
wxgTbGtJl1AVVry5lSipW9pZU+kByjIcxxYmLv7mE9HeKBK0gki0bpOQSoqZbFcq
graiRN8cV+CoqCNv6p4YI+NInvuOauKCN8X1h0c6Kx0IqkwBwws7BGuynSPEXyNa
ZrHpBBQW/6Nj6HXTb/btP2bvrSn7puoXEY0GocekzuG0+YEwX9rsCoRF2A8nXM1x
AjG3084iHq+69C84hJJ+ga++gsyTGEmuRb2r64Nq8KssXIfLHYTxBfbhp2gXpyq4
6UDXcmuG5iPzPQgD0N5RHuZGLRu9/vlbp+vwTJiSKoEMOLfFbVShlF3iOGazkE0O
Nh3lYz7eoLu4CySiFjpGeiiPyS0bPOcvaZPVv0ldy5fUo9mcZgmdhhRpvtRWCPC2
ZpQYOdk0p+/T71g0v8hZPHMjUxdVUeca79cRudILkCqYnwWIF3Dt2IlTrsDUU88i
WYAO4yymnZ6vr0sbGigz5Vpi9/6V1aLgsVU4cpYeTE73jlr4n0rUN8cQHD8OBRgs
TqqNaqBhr7Xq0Un/S1axi1/g2SEa6LWRzFXx4WlpnSJcCsGA3Y+Lq00DrBPWojKA
MN+nGSBw8kA8HMDkquSra0UlMgROE3K97QXVWYnUqGdncf1vg/0bNh7GInmPihJ6
BwYVJSD3MxcXJIz3miqxj1Kg61D+VDxWptRxVvhSqxYdoF917PTiESwWw9BphMfH
ENpj3UA9amuCGOsCxG5mI1nC4sb/RYFbXuF8ZUkC2X+g2n/RhaxeELRKpd3Utabn
zKGj9NFkNDlxxpnq8NmhknBiMcWPcFx086p5d9h0jUYxUUmEU1/cjeP7L8wOdpqI
gys5WqC7NHMVDk8wvsi20qPVka00KKaZAu1Alsq2WlyymQkKyECtx5wX83ES5jkC
Og6e95hV9CxLA/g8Q/rX5yIlvX639SdC9s6IKaXce+5kMJhDIaPPAVlJ+yGStCgu
Iql5m8OBov1OpOxMFRrYaZIni1AWMwHx+aqkKIvLbCeg6qghXUZqFf0+CB7XPKFO
D4ec+sDorPsI3jmWuTugGzq2R13YzfHGFYABdThYjOBjDihMYpD1ltfywz1qj3UI
NrJr+8szgsWhKUXmCfej9f0/uM63gCLAZsfqOnGuKhffKo/m+fShu86aLBQobwVI
BOE7P9PpqXmZgD23ZIPWAfk+UFPmaZCCyVvX8SCH70WU+rJQcDFov4MEbTYcUCSf
PRmRa1kUAETg9+0oazi8cqf9cfijgG0ry/3SPMmT6qlnXbyzFOPF6zrGEi7m1QEj
dc5zWJbqF0hpml+Z089GIDLNVwCqT9nKpA2kKTqQfPV+A1mI5VuK2hTHP0WtFbFC
b8CVXx2mw66QWdmrH3HKZVPken8j321aG0aCc54hyNYKxW59dxoAHn8yvgJ3X6Ue
DqK5nJI9tK9A/e5SgAFLoQL4nQX5jvzYO7CjmLvRfBTEJKqpamoHXMB469RhcXd6
BmqA2MI1CQTj/apXzhe49dmceLlmthfVyI3/7b4sdltDYGfqzYKYZ5sQdhOaArPT
zdPrcL4Ex7+8QgB9rzIbCterf7FiXp6zHfGOOZcU2KlVlTDqeiLhPncnRBgNWLiL
Sw6yAIpNV3fdcUvsq8BgmUg5pw9kaFBt2RnYtY8GItw4aXtDEFuHxGwC4/rRKrWh
oXtyzuxdN1CE4ljaKwMXxMoq5bWqTRxRzl9MzAFYN7D+39i+yb+rEkLSi4Pm4gWx
3AmfmdNB33Bg9zS0rXBkC2wNtHcVkLnYW3ab0QCO1N8V6YjPfhJ8yn2iaCkL+f6J
QYSgirLIQ4E0xOxbD9JrRa9s4M/672PxoQAUzufUDNF5g/eU/bESqk8n0ikAqJwB
SUT8HBeYzm1trqjVuXGxDzWwH12AoF0PThclBUBJBgTMLNR1xTMSu9oeOloGcOJ8
rfjI6r6P8q2Ujq/ejCaTyJmcU+JrFp39ts2/+s6pwgGY4zTpCUT/l9LMmE1lSrks
EmE4+G5Dv5CezgFQWeo/2zaHitTUEDsQogsymbp4aoD7EXVFKcE7DccrZcnww205
HvSts7bbj7CGA0/DL4n6BYrKFzTwp7xrBBCpEL+u/uV0gEWeoeCSNjrbsLH/Ot7i
5FbYBKgiNIdbkE+uOcWjcUJAhSl6z6R+I5BzY7rlm3hzTLq1h4f8ivg9/vZEfN/N
q9etZrOCuzT7MabpbVaPnlM6t0BjXbK7UASxKEcAPWd33UQ4DVwYpKUkcVnTMJpQ
pjVcORTe4RV/tt/FNUTaHpnmgAb6znkrP7+Lgtj7z5Ziymho0LOg4sRu5oQVCGiW
qyd/hlmhkJe3BzERZaRo0t0mqChOMCV4qSbmMGbR1RWEPCFr+hhxOFiQAfEv0HpT
dMZRPcyBe3mKPELT/sfwJFfo27JcMKl/yXbfqahghwew5hwkRguUpsA7Gw2ixSzc
HtTTtZAT6U74bztIlOFvwMi2RDusyZ/3G7LY8o9WZ/EL4JKv9gBoPJaUlZxbq7sH
B/IZA2JhVZa9TGbKDVSlWIP0vFGYBotAlPuL+4v7AnSwlHjb8THlFaBqR0yG38Cc
3197cfQYLT/QzfJPdoz7i3AXS+fQJ9Krr7zzyjD6/YxMPSN2xydElR21QxrRHMOo
dcbe0c3SKg6ALsNIYWxGYk/OemRi5XXFD2trPlbuWmicnS2Wb4SC0m9YeuB3Xn1M
p8fmDL4txB8Qv3fq3xj6sKlzILd4AreayDYAPRCqWFroi+kxdQpuqP3he9Cha8HL
VnSV+qygFYHd1Q0AlOeAJC8d503Cywk94d7GbGOVCp6D3TIjjACGz9nd+GUUKuZ9
MZGEVDVDBUrUkGdvbqUZ+FSiX9EOM38IwKJEc9EA6R6qxV+LAg7erlfSSzl5qfHr
KFpBs9O0OLeeQhDsXSD92vYyktlywtdNTdQ/nDLwp2clQcMFv+cgs9TJXeAfIaZq
9NJ9F7ZcP4rUAqeHTgR1bhqHd48CgPpr4XhFjC83yfTAuZJyAtcVnuQW1Ws/ANUI
5gheP0gUM5mp60z5LolyXhhyUaa63a7XrIjIDNKP2uy56pjHqZUWjHqZorRg/eDf
1y2hbCN/MxehCngBmJJUwNNoSGOOpzJXL1Ew94SGeMKc0SAX/rVpjEBbY3jjsT87
aAUVJikKQ44nlNApoDbEfso6bfD23r68Kia6b9rW2+2puTBP1gaAKpdH3HnVy7Ko
CsbCSZD4FmzlSgSVmeZ0++pusOAcafW44q9WsxyzjQlafW6nU2hjZooVQpUd1OFT
vQ8ZAmQDX/GOuQSAkCXtNgRQCLW9kOAd2DHAkRBkd4QiFu4bqFCjHdHx4afNO82/
CWAaD7Xi50lPBNl4nO+3RXR5bnIbf/2N2AF13LtNkX4ANPROIx0zdZG2XchHdXpN
pY03+vR6K5zdAKngzWGrWi938fUQe+M2gmcnhmoqwyQH8kqsuwQDzFVprxXMHM4d
DVUuSAVVIDsnmcXVYHnuQrw+Z8uEe92HE7IqhrbBKTOUUfnEYhprkb7+HV26T+aA
lhctlMfp26jnTWTYwxJeyUrLi7fyawYcVMjY2r1kEeiaHvY+Ag1u3hOLvZOVxvlx
xt13zzcO38KAwgSIctvV6zfDpescWVEoGiI649obgQirf4MdecnD0yhTqNuEcJcp
aDN0XpmcTiI2UzFjQF1eYy9XzUqPYo8cxGiV8KpPRTnfQ9zZFEp9tqWpNVTxCORY
UO/NUtqAMWeQXDRzEKHb0u4JDgbqoKLDnm6aokpiNnnJ3oKelo8jfvB5bKRuww3J
1okYXMLip/Fz0edQfDrQ22wEhY35VzzpmtiUTHVi0N3Zmdm48yahF+BNAoMlswIK
MvBaIwDAPOdqI63FJPrwv1OOAEMYo0e/AlqdjN4r2ulwdLvtNioJGj5T44pm9lBW
3kIvgOeY2V49z0HcpjzIdynEPn4pzJZlezTdCG4GX3lN0054SXWq6O4rjf2xZ0+J
a+gVudlMRxGCliJFAaJGa2/ZdoeZ7kBl8DDpkzCc3PBxlxKszjG+lZTNQsTiMD+L
upd4dWKmePlD6iJY6mmWsIT5d3d+GB+EzyW+3FkTKfnfBJdK9D7FT4TalZVinfwh
h4qEQEy0ercffwrVAvN4cg+PmtYMVETkqral6y29JrkAxm6TUZBSmmdQznSgSanC
XaSEjAraUPfX9iUGauEHl6L397TAsityeGtMp8Xnrbj2PUkJaZzOYopqY1O+YzG4
pzGMFTJ/pIY28+OsCyeroUSNTzegU05TDXBiqcX0bykHckETHOBWEtHKkPjmzPi1
/yj+SYt4dvuSthsWVR3ZFOcxP+9mFxbUbq6nw03wbQKgOSbrMplOqrKLMkoQBtPD
bXyu9iF5Nv12kcI+uu9xEPP+5uNc5IMS/12EuO6nRI+6RiaBgjyE8nz9WZvMQoCf
/VakAW4IegsIkKjzYrnIrMINwiChGwIW3F/pUvJmvmPWpqyJxCB/qWvdeenNJ3Fu
xIHU3s6fxTlate8NQ7x3pGqdLJVHGDJeEKSoO8Gz0VI0WqTjBxtsCIHPsgazdvwS
MR3JR23+2kFXjqRWEGnti3IY02ww7NZJh+IZIk72M4lfvYH/9ydi2BVdveIV1xxj
sAjiJ4ECMrw9AGWVDLbF5WAZaudWEXG1FbbAAQ0fM+Rl4u0W3pcqcJMkecknyj2m
wTL/UbrOnNfHefxkwlNSfgkaVEZA+YAXXJ0atPvyuH3irnEwFOORRzY12vzd13Id
H9jIhOGBJk3FU64zapZPwHIRclIGQXzrJlFsvT4TIFjTmn8EECRSZWaFjLUlTuC+
oQQj8k0ZKjRrGZL/Gg08fFLWQoMK1ign8G9d/x+BxbuFeetruPjtkMSxEojj2HMd
xWSPAjA8sMHxLPbvDuK+YZXpQkX7syo48DqqBQVo2A5oXNzzvULv5aP65onJwu/w
SgkXDdPq6JV47eWBs08naXkviEBF2M1eCPNWfba6INfrqwF9u9OzGEahklLqrohS
ePfpi+CKXISNCaI+FD2TB/ORxbbcWb30tW/RcmYpaBW6uYy2nAqO1BKKlgWRMVET
xwY7C7pRYlm+jtpR4e3BqKOBPZdf3VvsjB5eFwq59Yese8ghmJCeigiqIa1WZoXq
50d/WvXlEdtsflBDVsLnwBRXhfx42W/d+mmtPodvbH1IVrzcLezbWlL5kSChakkb
ABlsZXzcVpLK8I7sJ1VTuNoADp5AGNnea4acoT6nxHnjwVADI5CFHGsSAuO3Uctc
XMeaBltNCo42VU8HJ0K4byacpI4vTLOKsWKDXUtqruDNptDO2j6WwsAFkApoA1wT
Y4kdadO6qncM7YjbnlsfB9PE9BIAaTIDPcDblto9lL6V9EHULLACOQvicS3Kz178
kDutlPJ9z7/NdUZuIcqMnIxBN16fT2570a168GcPjd7D1Hlgs0XdHiawJBTpQMXs
HZ/6eRHeRQQCKsOeHR9NFpUPUyRKJRIbAmXXV19bo0IaO07Yl0dWAPqvEBKFeGzK
0wnSeYXxDiLSVtn7QrHpc8WJqC/1jq5CGko+l+aPTrbCC51YoLvqI24ZS8/egNJ4
8eSFgyaV1Eh5wEoM/lUA7xh/FNNYjgqHR1CvSi3i0qFOXab6r3PRC6v9Kiqd1qvl
dv/829bgf5MLEXIgwKMx1oUXcvMzCxhVgddDzWrsJBcVdgTjkFgXJLu4/k3eO+4Z
9giuLg8cG/ncK7pduh6TrJITwAapASodIlxS+cH1OQzb9zfqgt4IL74Tv4rPwxdV
o0RE4kwiaH+YqOIAteiISHUfqnhTDqIxzoLiamuC55Z+0WDQapal+L+uJsZXr9OJ
1axvIpWgXxPcXMyeyGqZ8Yqlw0cpxOYNFaV5iXDQQfXD0BhBezEZNrZ5HCbiH7Oy
S/uJmMgXUfyRMA1EH9YXcyDrHTB6wSjeh/KEbwvuu8LlVs289CdT/skTiHlIPxj6
bEoaFo6JfIKKSz6+UUOoztkFYn0G7xVHBj0kTwwTqUhmqhPXfysUZK8qbKzNy1hJ
2guBEQFMVn7/uQ5UdlHw6lcnD1RThDcJsiiLbrL+7E/exraQoSyG2hD4iXfN5DtV
BOk9Rkl6nbxn8bmGj7bsjxYbqjFugxBigITWZbsSFmlb7adJexc18UI2PiGy5/oU
eP7IgPnnPn3ITt/RgWhMl6JsQhHslMYIrOfNttx5zyLSrokPanZdzh2687W6p7X7
CAebhp1il3YzOqHwWm/XSOQg8PVvvE0MUMrw/2E0kUNFpoHiSFdzLc5Dbw7b6N8R
EJgKXKIFgx75jiduulHR5zEHf9E+YAgA1lOEqCTSzu7uuRfQVWZIJU9k3YZo2j3C
ehlG3GXUd+1Rn8BFWZJgpONREHLs0bSyM+zZJguvkynAhQhVLJe1sWx0MSX0qKn5
7EodTrRr8ie57w9lxwHQzD0zZZs2KkCIIItvZ3iTzpPgrllaQQH9UGj1c6zN3oEN
TsphnIh3V/VfoNY9nKWb8BnH0/evI1TWGJZIGNM+qQQuCmlm7B161ZPRJvcu3vUZ
upn2hm193qyf9SQk/Aumn9gQ4Auwem5KQDevPnLNFtCaoImgMYcKPbfjgQLuczoB
vsp3Z412QzPUeKqXwUT/nBqJPE/ea3bRXIGH5IRD2lK4/yROg9tI63o46b3D8B2B
nY18UY1VZNIiFbcVlc8lOXpwdsxTv/77iBNHHtSDEUkb6Im6pjT0zHwQB9BqinNL
52V1Awcl5vjmP42Ui80cHMb9e+WBjkscJIjiD8k+IZ+YllU3QQm2irAhFKNGjJWS
NunFANJnKCzo8WuhPciTbzZ+HOYONyMwGAfd0YqxLjSWhUvuaMtcY4bG9FNfheZu
54NhWOTl9UhjaZwzI0HpEHTZLpMxBOCdna5QFI30ha4/CdtIgUNsQCrM1+1UNuKL
3bAFkCH1FnY9wo8/kmswoa7DXfeI0THRsC03WIZ3kxNHF2noaDBWed3WnjpX30dF
rbFXCCjEVY31racr0cssS5ZOj1qOaMGObEN/J+9fV7qKMOz2z2cwakXOEiGNKXZ0
4cjRKtw8vgYRJlfF9m+8weOqMTX7dsO1YPKnfea7TyU56DPcKiP4ZVIeNTzZHfXX
jwQoMCXKgN4GHXV67JI5V64uGKcIBeEkuGLQPDmZior6ytcScH99kT2wjj0glD40
BFK+fgn0agZB4f2tT8+HuhKjAMQk5dGFxWlqwMGtShtpt31r8x6f5Wr83cvrim3G
aYi30rPJw+AjU7l1kwpGy4Lsnm9xUJ121U2OnaT6zHgX1pgR+P6yXgDlnLiqZFGk
+sLk2bBB2dkI+bAtdKioknacFZibKsOg7+5m/qwQheCUpmJwDvuwQ7TbunfQ79U1
rHj2aA0VyRJtVsGQpWYkl8oQMhfqkNBCOSfmh9DUNagcgsMLkEWUUfrg2IPJp3qo
w93L/VtfGouXR9uTatCzngqU2F1eGF66yjYMZa0hJpga/xlLJd6V2eQ65AfZEhL4
2DM6r9rdKh7L1A9dlToGKf2qJNBn0XZLj0UkhP4hFXDaRaPGOdpA8APtFnHnY940
b8c7GTDyz8TSqPLeLS+vjtwK4I8Yak3ZKmpzT3J/IcbDCbdIBtS1/1JibVM7c8K9
b9WntuLvQfpstcn0oeIOmd6XZGJbO4iZtBVyNmecMd/OPg9jnXaZU6yV/pDB3wn6
/y2BUdAbRSzv5F/Vd4K07fT5gbVDJ0zwCpVq1fzZ74YW4UMP9Z2sdfxw+79yiT+c
EOe1tWYOBxuKf9P0k9aouUChcsalLFQocGNNBAjliV2tCIi6iikKI3qrxHgowdV7
ArIh0OHZxhAjBWO4heRSg20FTXNedYSgLjmUDuqMDMWw+bOqWL/k+OJU7T1HXI8x
pttv+JrCFdeuBRtu0iJ/q/E3cRkU3C1DxxYJR8ZRSu/YOqM5sz/nSceWrv3NCclt
3kaN6HmR7tDoiasnrRvgUUlxdDrVqAhjzWl8U2iGHVKiLPB6Z5UetHH6at44zlKP
2ROwGsCRmnwAT3ffsvNvHhyDZbxYKELhthGKHbrKLRg7ULniQ4dgmjoo6IRexi/g
W+o//XMsmXG/E661LlqOGcBRz+EVb8BjprrJrTZZS5grAM2VUo3/KQwhI4DjXBqT
b7Vnjp82nf9+7uiCnMdBRMcK6wUJ8ipqW9XHOlsETfojM7jq/TMz89bVjGHnNVU/
tSdyUyp1nYwRk9ND6H+I3H+NcLCAIv4hgdItwjdEAF+npYpgN03UYzOe50qSJTPB
q1kcsCB8/slI8I3wFSaTGPKtBz9lzeG9uJgOUxT5rhcyM6ZYaP0KSxi2fb3Y1oyY
LkYlxAIasiAokq95V1zcIBBM370qHPDJK7AJsFFUmVrFFYOo35oephOPumD/WP7b
4+7dDhb3yvMANJpiJxOhGS5YnqfGWosXJKUMNK4tpSSsi05cHDxhNEBzS79mgAtL
UbGLtdYbV0GgLy2uJO40NSehDBTnbadPqwMDBvHh/l1zQhBtBh1ty6fJ0qbVJVsh
J8epW8Yc1amhga1OQrSkC2HqZK5g0fZzo78oX+3REbnuqrA2sSqdn/ESR67qh1gJ
J35Oiz/UWhRpjml0HQmPAH6KUtpe2fWf01p2x3iCIBjXlAa9ZwKHOezMU0wx8F+H
4qRkyMWxrSZxCw44FFvzJHqTs3tUcFkUTxTkpWaas4BUs+IbVSBMG3K3RhQZ3DoG
tNnKqz5av9GaFSlB0mHUf3K8SXRpn8EAVt1sU5QQWy+z6hYrifCl7eVzbqcbYOys
HbP/PQFEOMZ1/RPXqb1INV1DIr2YPTDxlVmy+X1RwWzIXECcDhKAh7e5rxxUzOq6
YyH3dKyITo1WI1r9ajBjj5STKiCdbgfCjhiAvYZ8HoE/Xj01vQt0vK2pd7Mk4QEK
3XOnaI6U/rIXptZHy4mOgQLJFf1aH/s/ctJBYc/jflfRM38Yww+BZOCRE2328rHf
m/UAYVa6wt0uW1sQ06x/8eY6j31T6+wrDB2rs+snSs24jALPxYnwNjOdyXCFXOzs
tNp98YkiUxHpZ+/gGZGC0+KIMh/rSTJa8BAE++7T3pxTh1W0sGTgHYkSdWMW02vT
VLHlMpIIr2fUg7FTi+IXq2NjXicb52bnowXsuVxq1fwtxVCSBn/P1dOh7Y3KaHiC
txAKO9Q/cDhrM+rfilKv5CtCIrkpgvJO9OaG2obpocs4GLZ3HLWfqbYNz1Axeumt
DL+h4eXQKa3xUuu1DovJScJyM2pknT+ODE5IEmexP9nItSDRPgWb4nsIDr/4g2Ya
3S/QEfffLy+ggeSiabvPw80UEom+I6GFNsNQyDxI5Wxo8EDUEAsUy6Nscan5CSUW
TUY4LtnKf/mRmh+OPRt1v3WNxJxxY6qQjs3E8uOAbO4tGmWFNb8e4JjscFe4YOMl
/mlHd+20mvwYkqQ/eCRjI40xtB2/KWUNfhQ6k8sz09AZeXkb5p3OJgkuGRdZSbT5
Luhrxj25uB4nAZsPZ9r7QALAtW+55AsqPscmeQqt9PwqN37JlrWGhAFhrt5wykvP
/zGmT41xxUsKvpJnz8taQ7qh9h1vrkCD9On0Pz48UBHf+f4xECIntMxbkznErhWj
xz0y2P1Z8w9dqyEFyQtI8gnptA4O6KxImb74uTW0/6PVDO8bxouO/caPmXsg412w
IANNatsG/PsFQOK5y62vpVHYkGLQ447wc7GPON4FXRtkKVm+mfE8puqS4pps2zsD
gsx7o/boCcnJxi8pROD0i7DxiMQk4YUTctTckY32IzzLGnsziwQibFXLxPt31grE
jQhKLpBY8U+/96LA0NlJkD/IyLS+ctB60Wthtg20YEjhrVY3a83GdWuYobOb2qmw
rwoENEDBzG1Ixrmnr29P81DHhImMuzWqhmktaFf4hCp5PrclqyePJfpsUX5MXCes
dV++Yx0rGXro1B+CBkr5Ezn+K4KoaXUc6wx5HtcNHB0j/8Hqgb4AZ4aUIXZ7sGI/
bM+qx3qj+CwULhDPevMIKDkgVUFGn4N8/lXM2IZmzFzqGHd6b/j1DA+UW0/kaylg
whkb5kzmAdbIUQeB3ecmbMAue/lbtsBzYk2tv+uYK7nOJwgEsJAYL9rUGESGo6U8
vRT5g/LX1pIOs0MqScTMlKvl2dURvVmnnpnXop0aLpKXr/xskw/zwI4EbsN/xhyR
u4iBoIPr+G/vFc+2hH+y59syADPfJXrLMhGvB8sYfKNkkUh9mZsTPGZ+UKvJ7FV6
NBebd78DiFIyUFpkMZWQa0T6o52DvZhoyqwIzITSrqzOmt2VQS5VkNWjayb3CRKu
`protect END_PROTECTED
