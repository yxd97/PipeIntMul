`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJeZ4fu4x/bem6sboQ4xDBupBhfn19Bqx0n5T2pPZ/MF8huge2Hb8ouUtyAwQSSZ
mkCa/5VaPI+kku0x0LxlDG7x3SHbPUh/v0Oeyzved4rYAQnbc6yysOJpo+BBxr2A
52zGHSyjCfNWxgH//VZMija8q55ab6l6TlwEIr0zW6MtXW9rnx+Ef48y61fWc9KV
Yh/1ogF64AgU/hyPIIbH6oxtXCKnojDkMkNHuCWZqHxuuLFak4DXbUJIsE7RCqAj
vqHVkgl6jIW+zZCY5wTAGlW1ciKOUpEU9hbYAuhm1DLsklGYYO+NOfVTIxLLgguk
dy4+NUoaiDWwIfKZAlAh2H7yZB1qle/KHTgtEX8iSDQvU9F/HOaic3vzFP+26wqo
Qfnb2ALC5NREVW5IY+Fu4ODsrYVlJZ4Sbm84f5Bns8rNFIN3V0RzY4k2AS569Toj
IKGnQkurm061vLUJBcd2h0NLaNKfNANS+/tgai+54b6em2GmWIiseokjuMWQfInw
YPqwF9/5vGWWo3zkeRxOpm+H2cpzDUxPZFSmr1x+UTEicXwvh4541A7M1hgj/mQ/
IrszeQyDeW8FJKS8hFX5oGFnDjYnon+OUxg0PGwEf9tPfn9aIILFDUKeuOo6DW+o
Mrko+84S9KIBJ4wH7PxIX7rMfsst69K/e6AxrEyD1Jibjaz1orssMdIax8Gc9VDs
dsNhEWwhUWfwA/t56Ivbi4BgcpQx6CSylyVJ8C0QuyopcZl1nBKeZAsACzjL6VDE
VjTPBI3BDyl9A3NO+fn4+MX8OpJXCsW+AZO2ycXiXGlOyGaumLW62FQEJJRe5CYX
hlpIp4gH42naPy6x/MRA5L+XTHbiCjKfc9c2+R4dMQPrVb/nbuV1KCU3Tzl9xply
yoFYhW7aHbrvr2Cc2wOLjioamLUx8OV4xeL4XxTeHV0cTe3DpUz3cgFapqRowTZu
wVmGW98i3yxEL/XmObr0tXQ42MyFh182tSukU/gw9wREdeCuQBgceTjjZe3yJ+72
jRhzAXXdHenvbaJ7aA6ZPhyCjn5IwyjappPxwB3gCBGc86NpqEURBzlbDkCYYjmm
Abgzik3qskXVeNtQ+ldIUT6JOoDMldE5Ko7QvG0gyngm693gf9B1Toh/12T/wTjr
pJqCZWyEjb4XB4wyiZgXcWp0CBD4T9nwe9LdL+m41m8Oyz1zJsqMYAmoYDgMdS27
aA9ajzGPb6dG4o9wWfPFbQPn1w04HrWnzNdqqTiwGobAIa56cwNPSqDC1LNXH3Yj
`protect END_PROTECTED
