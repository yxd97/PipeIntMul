`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqxbKIJIOYkFv4qwGyL0pCUe/smZNJP6KWV2f8iAd0F/dssAOQ1Yk12lPkicaYYr
O7m66ea7+Qw9Jtzh7OF7hk7Z8TCui4+FDs4G8p34bvfrttFHi7li6CtJo6Fpl0w1
Jpcs6Aac6EOx4ABV0H7JO7eq4xrP0Ipmk/SQfs8Tg/w0dA8NpxTfbzjg+lXxH0k6
AIB2GUeXdyHtZWDbjeGi4OZbQd/YBIe9rnqx0lB97WgVUMggt3jnu/LP0NtAhFe3
oNu8oZOCKxrvCERwzFEe6F1+c3OvGyqEpFha1e1Q/YhIzhiFm69idSyTPYgRGgGn
CWaVjkSiV4g/adnlEQQ/LDheqvcBL44QH1Rmvd7z/viD+n6otDNwLEtghpIXGqns
zxDT0iawMH+DpqTcfAZ1nTtmaNjDDGelQ+D6RijTTLcOVw4tOGx7sRi6urVIfaLn
`protect END_PROTECTED
