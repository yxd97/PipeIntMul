`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/BtOIo5uPUi9D6+JdP3Pcf8nydzoInkfmucvO7N2g5Qau5igtSnCuanlaP8784zg
EErVy0AdHmzdfFztkcoXidAk2NUhcJmoGkktqRFlQVRf5wbknM0lvOcvXZ1K2U/5
4f4BftJxlCVuspnUIzILvt2QmIlJSTOqfSodXwWVTSbyhNMy5pgfykq/+Frnak+Z
KoioYLcoBS2yuE9imWH4PY3CIE8L9kuBJo1TBcyByB3srbTx15+PqVmN3P2mdFy3
DLbz+i8Fbiuiv2cCgB+LyYbGxRag4YZiBPGHQByF4rvV0Cc/ojqo99tazO9J/oYp
FWPq9AzSKTNRYVbyOoyEieDX9MZGq64C4jrp9BcLcv8JQIGFCSAJjIxmaQPUoPKf
vFqiVxhs0EAYQhcB26GoIT3XQkJbJ0Aa0pjQY53TUChNwT9ak3aVh22OarBdbQTg
puewGg1KBeGuBtMKSOHANkybQMiVAl+H8ulQQoQ6ydO5ZrKzeZBIirqEmJ/AKsn9
I9GZKaZm6Pid9Oe2Dl649znP1wEeWhiwqRm168E3/GCMolX2NAAFRMW/X9n1Up4h
Q6jxKu3gs9Kbkhlu9y8nXSS7vUigbUPXSAndK/fyej+agZFw5IEcQGaBR4iZuw2b
GqFMliSWNInJMUDgBMKSNw==
`protect END_PROTECTED
