`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swyYgkM55Mz0SVMFQrAcbNORiVSkInchQQ1Vg8H/qu09bawh3Fa2ydGW6KvXOSSK
VtziIIDyQRTWl3U0Nd6fAY+YhGakwEqhOQ/4AThjApMSveHIqGTamD6JNSO14kRs
kRtvaNE9eEzgdiAII5/iGnUlC4acu8Cj2lrVbHzKCcgNehCSYWwOl0/Ibhhf2P72
pqEvTIz+OsOIRsnc93LW3cUboTJUzy7IaGbf6R8Sb/PiU1YCvOrwR74X3G9KNZ3R
ahSoEKWztUpIictKjwgxVkwSf8s3Mrq93eQO4Ohpap12DDmfxMeCyvHZqQ2ng33/
6bG2JoEoqdSWYBUFAGTjNeC5beGobaom5HdQgxl12HVZ4VRQWcZwF5wVAKSlf1hb
fZfPrRGp+kY8gZfs0TYNn/hUY/uId1QwY/xebZp3fphzAXHpE2UtlJcTmyTKcP+Y
PUrh5bNmbjY2SBCRHtEPGO9RW7CrLFiyJ1kierf83KCykxIGMYX9cIfB10hkktRu
HN2jN1Il0YQffj+7l0zN0Pv2b3ccl8Cvnt+fUdN3YpuH+BYgJuuteqEcgat9LQVZ
Cs4j+Cv8/WkoqN3fiW61jlOSbqnHeX5jMQCGOdOdvNaW6GS9JQwbN+3Qez2JwvEj
8LfgilvswBslWapxbisZtznR9lJKLoUqT9tVpt6MP8o=
`protect END_PROTECTED
