`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4ZRdkXDKYyAhK2/ILpTwZ6Il0X2zi6qZS0ewr/VJoe5IJEXOLz4u65nVDT2xHie
VPsoa1XeXpfvtklyldNiCB8vkMUL6tR0GpqlW3GaNnyNOxk6SyEbgWjWdpx2g/22
gsnltgQ6rB3nwmlrDKoz1SIhNBmwlhTAhsFLSFOaUwBjTcnD7pF1qLpidgwu4B+l
kBhUgD1EfdvIiFM+VlxzBCnwC0Byc7FQA6FAQJUl8VpoZjThLaLv7+w+HcReZu4j
oNyKmBcFqsCtSWYQA0LFvo8Sr5JVC4l2LiLazfknFtiKmMpKkACLxWcT19TKM4rK
N2NlygzwEi/PGSye7+hWuA==
`protect END_PROTECTED
