`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ui+YUp1iAmahZxUTXyouaV9hyVDkNqW+mpkFJ9ZsLEDiy2kZMXGTl2zbt2HVKjvC
iGFcbFq004zQdXi5gFrj48M/4ncywJKGMWzvI7QpOjgXjRBLHfatydJQkOWDENfQ
/ttBLiW71Tov7ZVdTCgo0GKVn0bU5y0p6wd/IMGwVR5d+fLdY6e1+vFrXbghriev
/prZFWReO9R0aJttOvwygeiD4VSKrfsRaLmHOEYUi//ZvMLnzrmgINTwkgz94K9z
c/pNqumGYHgSIyRdD0UgXVts6c4aQrDTOWbp8KSC9bL5yUcGhiWyjczetcSxQSBm
Dv5JRXzrnpEMni6RyGkf8AhbZaymKlQxxgQ78YYwX6YCFzexQjQefNkyAw+QSPx/
UITz2Obtws30ahNiXjQ4kgaQ1tpJODs0npunW6DaWIYE1U6mXKqFN11laE8aj+P3
CPjNEO7T9KVRC/rDPJSpgZXCSCHU8xjaE9pGQ3XwYW3zTe/4U/yVGMZ0gls5NgeP
jzVcuEVXwpx33bpvqFLldGFIiWZNA/qii17THvq7bwArOA5Fq3XYFxcMhMhUIRvs
63LE1vzK5XkpxywU4Uy5aZ5h3phZ8t6fUrkOJNEFt2v5gs1VDVxq4UMlFY4Lc2Kl
khGgOScVtGubG/ttlZIbOvLVXP4ARQMAbu8Ke0NRVLBGM45gK8nXJkKpN4gbyziI
Wk5rCK5Gi4oOEYpMsQt77AheoNtojOvIMgL1+vH8eErnHE/QG/XuweivqRa4ifUh
vzzHkeR/8vwZCPSENoznQnvzzugqi8cnyGoPV+jInNPTB7gUtgUioiDD4vtYV3Ce
UcI4TaeLQGA8/5M4UlE3cvR+jhx0fRhWoJxTGhtbLLKoU9pPMvpS13Emfg2y8wZ8
RnLKEDM0sE40g3NWGS0tvEwrwYirucw9ZYJMheS/UF1s7P9acQEGcdEhF+7wdWWk
4V5BFUSg/o6QpXPg+GimwuzbYfnETreWWGq2mLtPTUEJV+Aile9E8zjIYMSujzvm
dBeFcdMfHvrvd1NWZcBtY+ZeBZENX4J8WyjlGG4Ilbtkp2YkCY/OxTWtjy+axcA2
tIZXnZtfLIIp+IPBeNrztlRoZJZFNwB1WZyaV3zJduu5vloZr/RYJMdL/D7OIKN9
3WbVQKbOq78qHlj8Q1Cm9Wk8HJpGulz2Rrc8apzS4t6L6lY/Fd1PU62aydJLmsSn
hr04/I8oVFlta/KQFLHAhNUPGXXQwq260Asgc4FlRLvcX/5jl5AMgOrwtBSOggm1
oX3DC+/D7HPIyZZxBL1b3PrxT2Mtt/Bjkv+pQIu3+4grYJ7QlKOlsduqMQ4A8KF/
qsdbysVqo5kPp861jDeacJUgOC4Qwykixji3goYqZzmYLO+lmbdx487YtUQiWtx3
aWFEuI6w0D25ZulnQ6ULGJATMZBBpgYoE46eYAcvdTM5w3MH1pPkceCiK1JwyBss
n5BtUUfljsobQzIjZgYhvQ==
`protect END_PROTECTED
