`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HR26uQhty2INbkq1qkj61Wmv/6SDTyHduUZyFe+cd4IvuW9XIdEIYUhIq/bWUYXb
FKqVYiokpuaP7q+WF5oUA4rFQSwZxxaTCPMEO2ZMviXYtMDkn8ptaJCko2JNFe6D
pAQLHC9YJu5pXa3LVWla2KV3eW8IVV4fQZSR0zooZKSLuTFPsiq78Hjxokvf/i/r
IwJ0Gs3X7MHBYQZaR5zrt6fVAXnZMemAlfLKJl5iPRdMvWWVxnAh54JeM3/RGNBP
ie9GOuWXfGHwEjP9vPhDow==
`protect END_PROTECTED
