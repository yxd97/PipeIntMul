`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/nKzp12XKZWZJQFwXTRpugFGgCzfwseHw/yRqmtbx3/uewF+/8UjTlZNf/r3OOQI
aBeH0da1QC8wO5/okU8E5MyQoFVvLdjhr4i1Ggnq2JwrLOIjVns2wW6axQijGno2
Eo2cPoQfkWaIJMVemhwtMeKCGp+So6d8a2xOz9Tnm3VwSHcRqJVrJLkviNXOse1b
9c6Wjfheo9gg1tjBm7+1u1Qs6tLPsh+vBAZY54mSX8u3l7HwbzlYUnhFoIjXdSrb
L3h/VBsIJHbmgSJU6HnNSh2ozQicJlstqxhkiBG7cOMoKNP3nkpB2eFFLq1OTg4Z
bMf4Vq5vruFJA8wvvZHw32Wf1gTcx//KbqP0Ayw2RWM4Ow8AMVh00lPdqJl8Al/h
mCZcnFuI0rvte/+daO8XpBqwAO3MSMa+PjMtmfh8kjJoTj/JBbwt1I/l9ubRbeOA
h13gxadL2XUIw0a2EC56vTF1NvNUyJ0f5X0+FGS0SC+377l+1MzM0kLyYU0V5deK
C7IR2v7/w3+ezyqzrlLzK+CpO4qw9VLTwdn2X+awlP7EWvsVoz22Uyxh6xIp7gzl
407dV22Xz6i+tJToNPmnzMrGKdUxNZ4yEbB22w39OReiwy4w8xJVeZA2cp/XXhUH
Qi/Qlqnkyfhv6wWb8hLa2cIByiwAnjX1XNpoLjaYxPUlI62fsbIS6xTiEl7rcgW9
8xyHbdJL/hCxHhpU6gp/KQ==
`protect END_PROTECTED
