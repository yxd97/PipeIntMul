`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7OBHaPOc+v4keXvWNsk8XU1HpO53pmTz8rLBqngfnGQLK4TBuNyqMg59jKnDPU1k
FrZnDCqY23mNezB3xyKKmAOHlsutuaeshe+U6DUUTowEsLVh3WRurAwl88IzXuTa
pNYS3nx0rTp8zMIk1r5ip3LIgKpD/Pc+P/iY4UKvw154PxHdYnUes1f31dAQBsYf
DL7sGAHMryHCTMoMyko8VZILXYDEQZCx8WJxr+hQ0Wy3IU1/uuH//wmVkL4O3/LG
Qda/GJ74DVHuZweJG4u6TA==
`protect END_PROTECTED
