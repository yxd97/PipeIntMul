`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Y8oN4AMS71pet1Yf7wZBKR0OqCeJTVXyZdk5gNdCFimmMYLR+9R3ILqCeGjOHpk
1ZSw+7SDB8Vvmyw38hVQUN9s5BqLisrc0JH7Wwtce51fn+cLODw52ynqba53fFoG
iwSc8crlQOPF7PXZZ7a3IPIlCPuxyLnXpqrZBiqA27hXKoMXqa0ThdJBHOjwWv8k
aetSxp7uexuwVoYmAUB5B1y27F1EtpPLhxU6P1eBvqKItUtT6/lEh+IERpBcUhtP
DOv6ZIvmTDy3NpL96kdfXKAaE1aevHaEBEA6unAMwYWV8YAD2xbjpAfzjq6jfhK3
9v+ET8vQL5rlj0Rx4ZoAScBO1gvbD3mBPlVkFeX6FMhWhAbQdvH6q/akfNlNpmRF
SoqQF2RJ5axEkjip23sae8TC+CvtpFYCYHMBa6nDyS8=
`protect END_PROTECTED
