`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ItOSNWArXDCCw+qZOvlJAzta3AZWHqURuyExh4y51pdednm0To5IFcNp+gfZoG05
fnRDewCH3GpxKND6ueAllhujRoIw9nD5d8marvQ7sDUU2JSEvOzTVi2n7Ea5gyaC
lSoeKl8w+WGyzTfrImzMWcNwvx4gihXdUAmgWme3loeaAJIb85q1ZnL0BIrBLbgK
PtRZfLJzHq0ID5K1SEIOxurp/liTlTXuMK48WUv4Kh0aTPgHO9QmIPpkdwkV2uGX
s/CRGWKMwDDimaqZP1dM3oh4cwUMJV3DMkdvaAVh/qZ/WKw2nqbqHMvuzDGhHe13
hhAp0inW1KvKW7wWa5yCvani60SG5ukUQAZDMELa+d2I6EYixzf+PdocbOTWVNGY
MakgGdQgVJtsHP6oX4PVq8aR4uLlNPptuwVApIV0AD18XM8HDlYI+JrLwyjE9N8h
CX/Mz978kXxGh5KwrltRWbCNPfx9CWB0TFuw/9t6YiucGQvrkff2EscmZwBGUmna
P053GIpC7mPmvZZZFm9y5S2tKoPrt+dwd5gr25kaf7q6mCONcUSvUF2fazkVK/mB
8iAXpwko7lUqrLFOtLir2t9Nxlq/TeZkZd9V8ZbRngBA0IAJachFSAioK1LjXcYI
`protect END_PROTECTED
