`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rU7UYj1mwDkpacdjQt2nBqWkwjgqhnDNmswEs5RrRxMl3DCrutiP7qyvp475qjFI
y/LYKSlXYnW36fMeOxpIsracuH/b76VjtZO8+xac7gAi2g76Wha1b0YE3aTSVMZR
8tHz65MRAD6EXzkxfYIZZElmN2dd7rxfHrf6AuRJA1WQq192Pvi4b+gmfyOYvMOp
LlGjeL8Z5RJfdo3AKuTBNb1gzYZQU+LPkmgWCpLrM1/5sEPU3p2CkUtuTpEnAMGB
JFZOa253j4FHTBkhgKlLo1I8qXUb0OBS/63A8jC9rqwVk3id1GnjPvuUXODnSmRc
6M5BEisyRv2IqJE7zx0M42j/jrooWvlSupIh87WjMLtpJuBWYRzNA9lT7Q2OdL7h
6UdUqho16btQo+uL8MDW8yXHR4Uuk3a1i+FqQ/yOwRNlrK8S51j17PI0RGZ7bKqB
`protect END_PROTECTED
