`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rGXksa1+dLbKbcSmmq1qM9Uq/Dw9gUMGnx8CyOSnWypcecBcJGPI87Y2aKLhdjk
c8rRMHK6hFsKwpCP+MaMezdyykGWEe62QwPglJyyHrRCmA1OiBXomdH1LGXU6B04
XxSnxjnHNSuAwFo+1JnwVLPUGoGfewAhzaS4ZSZngbqq0GpkBlduRfCR9ZR+U+rq
fzbuYgtJ1axBfRGUtUcozMeojtUgGgPkYkSPmjpoRgt6srk4Dt5Pog3p6cQVKCJ2
2IBVi0B9IXbur4B+wj6sQTei7iLAy5Bn6OPnoSwa15cIMapr0KuVnHM3boqu9/FP
+zzp6Fk4oZHboa28KX4yFUh5W76yqrpskJlGBtn0lJgkI3EOmxwRnnkrzn1zt1U9
2aHdKUjVd7s34Ki/OqxdAhjjGkkMJTaKMsjZ1mfsYG4iGkOaQyBG8ZY6kKUt6/8u
VjVJhwctKOlvhtTyd0rJ/4hgUAOY8uNWtAnwoEh3LVg/xwXJbysLBGO3a2nJ1WZ2
1MJ0rHrHgvr5BMRt+ko38DniCQY/407KAPSoV29CIwHfC90so7xjuOr+c5InNBE2
INkCCF8uu4wvJWm4Qym0eaYhb9/4OqfEq7mA3N4bwrwfrgwLqxqinHaZRet+YAUv
uKEM5n8fOvgX4J2tMC4tJ0CAHOt5RmBW8rXICLbNz3ViZqSAHKcD/usu74C0bPjw
82b+vx5o8EaZgz3iPFyxuuLIGyAaI4e4PrF8c7LrY2sheUsBlPnUSTtnpjugUyP6
LCaIQczcdFQBIwz/4nY3s35W8P2ncG536ofWH56/3fKIYbSQ4D5EizRVHYYY1C5Z
VC+br0omjZ9Lht9ka0n4hRRh6X8bj3F/90L1IJchbYkduUpY5R0zhgJEFeKUqlm+
v361oEuYjw8/qe4Ei9A61JkW/IngkSTAgOhn1krj/KtMe0mU07CJiv84DcqbxXZE
cFbyZJ+oxMor3Ia2EPJh0048UWKsowe9tf5SyPp1ysKy8xV0pk381Xf5RA67bsXl
5Pojs3V8QU2bmOsn1fLREYsDcSeARcHvJPFqaXTfkm8tIT9qDtp8I1u3suDH14Oi
8on5CuJ5YeywLkseARXjKQGRKhTwuuv98DSiRMDuUvEE7BQXJlxwb4bKw+7PGdTO
mL5Om0+wm2KfvLVBtAqcN23Kg6a0KOoSwWpX92gL1pQm76gicVlEgAdIKU77X2FZ
BoJ8UEpBzjy06cM9m4Ym/eLmAmWbns/rr83w9/dFhq8+YldJ/2uNgRTd4dC6VijD
XPgHkv2z8Bj4fRmHRJj807D6MpdbSeruhJZ4snuxA6lLMbsQMthsQ9P1stOwRt3B
HjF+A6mqM+YHV0Sq8EyEiuJRBvutdS38zP8ekvIt/bB0ErR7GYIy6ZfeZ5bheGBw
NioVa0yBDvtQ9EeeYn2C4dg+fnM3hqmpgpX8Eb1pq0dYa3zvnO/tHDN9lhA9OUi9
q1zXVnDMITAWyPTXTkCwqYibAaIAFIWDnDWDn6NDObBzG0F+XPTLNZJXT0FUTHER
RARhAKIV9CIqTvkqGKsqUUIF5zP0CajEDc+V1LOBvppOAyp+SeY75nzEihLnN2rn
Mkw1OVN88UUjJ7ho2qYHnzUvtB25aUwtNalWw7qaXTp6nkaE1q2rwDtDb5cAGqbw
w+KRHxzcbIwawasPVZbrM0qI+mHVC9IPttf5wyEccUl/K5VSNx6JXqyWDMNJOf/Q
hmDpS8VVuptp9j8XieJDzw/3EJLIJ6aoyhuVWqcF0MbOE7KrF2A2MOYsxKwEhtS7
28Ht0UP+oJEE0MPAIN/NxDPiChK6oOh3Sdps+ZJLAnN4ge/SRd6AJEAdIKYK+SiR
Q9aSPN/xOTPBHdho+eHjf4+e5xYXxzI79HMeXoJfFQ5RTUD4X+oU7Dx7pjaUTtKy
GdkhD/QBTexKknjGKJ/t91YFmJQjGLerdtbpZeflo1cA3cAybPp9NrCovti0fGU4
ohhSyOZ98g/FoYPcvMl8+nCf4X47rasVxeB0WoDqZSYC0b5HRAiPFxQWrO5pYqyE
JZA1A03uu9s+3qVgigHlxMTduRIMaHZWJYSOTL4zksK3MfBMoZEzvvCstdm/DhEV
EpnnICnROsCA4APCvTkDYC+8HT7vvyHnd5uIKREFz4JhIf6uP2LoJqd6tDUQbsFn
3XfGPyA+jK2uv/gujjOWuOypcG6lyYi/plqimMtRi0KNCQtmuOPyzJvZrfQrdkdy
mgdsPMFQtSICMQq3oPv1AKWxo6Q78qB6m4tMcqACPsWJZweoUtpMPEMPEtD+Wke7
hVkikxRJppggYlOtMIpwhrO+PzmRLilcWHGHt1z1pfvMYC69J/JSKT5sHf87jL+r
/ZcsuJVnGPgYv2ANZzjRyGx43I/QnhCt3CdAu3FIosInCVmiHYeftHIh4PFaiRhA
kfDN7fUdW9lkY+ee4ZL/6h9WbzVibpphP2hqolgjp0RCb2anbdNZG6GW01SLpiXg
ItXlqsF6GMQAvs+lNDH5W2iSvafzd2EXKBT0J9w8Bx2jRtE0L/f3gsiiDcPVWyEh
7iCOT4sHXiGQ5rsA2/4Xx7OheM0NnnASx1IEAPJkNEsJrVPYm4naeLpzfHPaXnyR
7YfrXAdg7F9dfJnWprsGm3jiBIn8k/kZOVJsTsx/C7kVpK1MHK4ev+m8y7dIf2JF
S4aZqMvh81IPNSAXYfeYhDIPhfS3KzpDAnHuRkIJHmhj9K/LPfbZL3rFYHF5qwg+
TzBoxuemaAxc7ZvRJq8PsB4bkFOBz7YyR6nshjWUK8icEtl6XoSWBx5sn1wvKQNm
AFLRpzCGM964cvRSyCChE92qApiFjYsaqssUCkQifJvqr3k/K6RH91RnaokEV9ye
64uh+hHFlbgUKaFCNZls+af4Oysi7Y6Oq4RY5ZbhTz7VUWE2vGFQw02eMUpAj1Su
s1Uy+XWWuHeTSZ2VtkrwuXOp3F34nwKTbLPRKz9OdHjyIDdTCRonshmvDgmoS15o
YWTVIfEOElXEYmQ8HpYjjVVSHCE54NfxV1FAmiEbfpaYfbSjoYvOH/ocDKccLRGJ
w93bpu3YYlMM4U7eEaQKkAcmZYZQbJDMjIXKXoTYx+r50YIv9aq2cegNMOQeQrwU
a5vyJsPOoSDIUaUU63d6r766cS49txULRFrwodAoULeauAPs4F0IJTFuiYalaXFP
TWOJPT/thSgmjc6g6VeRS2FmP4oTS0hQf0wHu3BoRzNermsCY7JP2+YFUL2YWcIn
xDasDspMv1xf6GhauGzGX4xTAiOrjiCaZfay6eKfyf9HrXu30A6S/q8ckRCqz1KX
401ew+J8X3kzFvzPJeSWUGZMaD7J9eBcEb2F+pJNVqdkD50qbvahueoMKi+4Okxn
Qq8RXhyWpK3wC42KSbKOITrzFZ87VoXQxpw80nPkaei4MqyL1kdJcAe6k6CllHkA
OsUpk1nfpV6JoZtuK+yIeXQCrz2yEWEEkqufkDWK9xaWKPGG7zU+wNZz2z2zfjXa
O7nHOi+Exqv19vYkxwnU6eLbCXAFVcpDjcwyhLSkdUwMTwBPtr2gj7V1KrrrJgd8
jaKamqnfLn+W507yCsKopb5noGfridUIEAAxd8xNC7cmXOms2F8gnVejXKqIlUaP
UlQC5T9yhEQC6gAtJZeZBs6ZqGY6RH/FuA0CmMR3MI3JKuCDXUKhLRyxSHc+zUgl
rTp6eEPP6br7vFBSMvDhnaKul99J8BEvo4zM5CKHbJIriPNCMhcOV22V0+0xUKNH
+TPvI6RVuc2AH2w6Oght7dMLpPEU9pkIcEgWUHGa3BgtyAYPINCI97EffV1ACRCe
Li9uLgkiT7xIu4hHi05odTZNpMQfavnnkVP6TPp2cYiOrLVLxmQY1aOlT/LzdG1D
zdA8zO9T1JwUoG3KNEpUeDvI7KiuMum7o2RN5e4ZXbFsSLNXLGxiDibM9qSq8kNU
k4ucfOe0FYfFzTJ+NYrszmwHd9jJAO21NRx4iLI4GWagEUDIj6+Y3JdfnEuOkbNb
ypFTuUul0eofHjqShaaRuW9SMoQvc0kHF1KX2NqAw40rcy8cJN/30XnwNeCYbzv5
eOkjxmmxlt0xBqaNquyQV0ApOeygapSrmn5QvbYgNGZmaSQvtYOA/D4JRUqljdDm
9uc/DzTDf4LdKvCEtf4i2H6m9vIOfy2/YsLzGdN/nDdBOxW6wWOCZZVbtCTl7mFu
bmDh0v0iAKokkGinwWA0YYWPpm0dZuVFWnhoM4NtzrcMqVy+Yd6jokBDum40fueA
PIYi8NQmX0BDXfPY7zcZN2AprbzQIa46+HJghKMcgISBfCeLYVklhZ5oIqZuDibC
tG7y2iSMrxcyoLm2iICJiKVN66t2olMUHq8ZbBlRcSCz+j7xAtA1gMRe2OurGDTP
ozPZhg9vUCX6z0pOP8GfeplQG1RYhoa7ypl+n2Qq62zjlvSVXH/TJ5A1z5GiKR74
CxJREl3O8VYEiLbjJYM9Jqz4NnFe+c0Il6P0oOKRWNzVJqTIebKmxwYVCifC/e+c
J02gH6psCfmTSachO8qL1qLtGms7e4xaFu+wJ6QZ9hipOagk6E639Tl+/uS/55ax
wXFwBx4L9a2FKb3h3jE/+30ayBnzKfMkT/A6VBs+JxIxYXdVeFUGEofnckKTkXsj
8xNX7uf5sWws9AqQv5SbRA7c6wv2xL+mo8GD5/a+N1Ai0qFTbPYRBuRHNTjcE6eO
5u0nWrfk7xG8fE6oHT4cyMcguYD8cpH8bA/VmnfzpAo/Zv/QoKeCB77MqvDrRvKT
dbNT20FfcuDbB2K0cKsZCsttv4AI+rE92InZfd481n4lUnt2VvrwzhhRfpO9wu1J
dk+1KOM5WmWnFfCmNfwWlGTeert6NN1qztVixE3uSH3KGaabFHkNBAYwTfM5AWcA
dl7QsrZ0hGqzvgrH4a9KPm/dULBtLQNBsHYKVqQzPZKd+0uX4F5WoWc+XL6gVrB4
/B29bzp8DdauA4JK9XLI4B/dyVLTePHGB9QgwRGlO/UjGQJYrTkDdolwokAe5gFW
/XVdMM8ez3E4sGQ67IQwYPtI2J3OP5MOPH64n9S4VWH72i4JDCbCbAppm8UQqYp6
MF75jPLAbNVhWVsEAIyhIeOXEPE4O20voIa1Ww2MdKCf0utw42UpkG9XgJ18PGOt
uEHJg5UELK1pzYgccrvz/zFqjiIE013Xw3geuPvfCgeMrdVehMYyAGQeihhbpQz0
h6//9fmXy28gQg6ywYmsF8ega8GUeWqkN1KgrZuyInefvjzItV76zB6TpiWZpZQq
YCiNoLNzHGFfNELixFx56q2StJllNxHOPjpl12JwbRnv3/h37SojhxCF3zvQQn7m
6BrKl7xxApsxUS+FVgsVbLYGTjvbbWSMpLC/7NbjUCaII9C5vY5YT20VGVnArZVs
diaNjXUj4zFJMhe/6mzHoKRThKcw1BFSZvH9On6HpyMWcjx8gxxvlp+Ze1g9nhGm
7/gBA1bl6q5lpLYg7EVg05Jpv5jvF1NjEdyAj/3Q9sXKdN0ojIXRoJ7QDU4wYyWp
88xyNDUOJ69reB8Cp3cWdzKB7sY4ovrfo6tByJhYHvEaLNLwAsxYzmlR/lMvEVpp
M6mX0zLjMtMkfIfO+y6IplTsnHMQp72fuVArw0qsBCFougQV2XWWJ3/JyqUDxvRc
LBpKo7WHrcvaOECij7aQRD8WCbMdehya6Y08TskFFgEXEp1aWPHR/MpjzncvQ7as
E8KcIpHaum0kA/Ryln/2hisySWO/UpzOXBkgwi8kCrTZuo1A3J7io0df9mico6cZ
0vdeu7dCgs5Lwi+sXyheCKhMwSRNzbkyLEQeBsGslkDdal3oakiDf/UujfPlxMS1
hsZVDQF585voxbDDLO05MRsZSiFSV8l3Zsx8aMm4JadHa0qWhmLVkhUDhJY2jkkX
Km51017E8j1uycT4otZkGp190ug5UGSijfMkr3IKIOGR6pwS6RZ0XJucOjQ9mH27
ud431i1tba+7lZ0TvL34Yb5so4goaF4+ml+GJEY4LT5rtJDh/WXTptd5DCmNKC1S
36PJ1l71uFKkHzrxAhDudVXlgdMOJllFnPZh+E63cj0KA3GKQagp7RAu3epXiwd/
pRnjLDFD9GKLKYaL7HDmuNYiu9TfjiUKqYMdXBHkPbIeulY/7pvPCgVS76WoWUCs
HzaZaUQ7yMyf7yX/pj1rHQkRuJJy1G/w95hdFqCG7IbyIomc4nG7RNKg9//aEv9Y
ItIBkncd/iIi6eS3U2PojKnDe8WSAmkE1GZajfFeSaUUMMG8HQRaQnSIbvKhLi7l
7cHg59vFv6h1hx8hSIJhN9LMhLL4hNfM1cZUqkckOmhTBspxpyjy5kXUYhI2FQZv
4FpO0Q6zU8PwMj2s0MFbEssGNSQl2wisA0yzMkjOJb4WqhzDkV6jFor+jPB46eBR
4TzRW07HtIT1mWKhwIgiDUubBb4AP9hxLxwiGhxBz+Szd59IIHaSWXmDd4MWmPnX
57tkuFarHaNIoXffozmPULntzFnvjw4G39377EqkNm04pNYknWhFzr6AeVbGpxzr
isgOiYhL6TwPaeyAucI8FWA0mfIDYfOKPvw4tsAX8AdU7lbUgo2G+BW6xnSOLmHm
93WRLbD+DvysekDXZxCIt4OjsYRRJ2rnURJQ3nzZul/vjceeCVLt9I2N2sz13Yu4
71YDKq08HDKE0DQgZznJqlxJRKfeuWSL0dxR7aPitEcO2RO2O2C5YsS6mkCzg5lO
Kigxwjj2hMqqyDlQ/dG0O6MFSevnMQzxp6gb2xUkHkQ7j9GnC5KRXtn7pyoPZZyl
H6xH3yfxDuBvY1rzuppFmWuje+sNq7xL26MKYJ0uP136tHB4pbUyUawC5PwHQw5X
6UPts3f+21Vl8K1ScwLPvaVJrlj2Kbv3pIn5hLXg6I4fIcMRGsBYkJD1uHpdUj0u
fKayFTs6MB2LkPWLHZeL1522cV2HP08EJs3tOTcuqa4vjWiQW4Ue4lTWgfqBCftm
uiYmSjO2f/n5kQl6pgxBB0paXZOBlfeAXUzTVploJe2nZu+p6e5hPMKnyrKapbZb
N2DItz8aR6g7W7KkOuT1qGKT5ZjQZgnOOX2cKluVp+JixWPetiYYrdSF4m34GZN7
k874YzNy0I4sYEBoqnhvkoQhiF6XjaWsWEjTbhFx6S/JqdasC6g7CXxcHbEHD0w1
ovM3RrnMarnjgvvQOosfWirRyurqMLOEx02Ttb973TLpSP438v4y/huKQtpmoPLH
OXNdcSYOigfp68P6Eq9zJIgqV4AH73ctDpOfw5E5jyFEF1TS+1RsenvFWl6jtisO
rmFYaKA3mEwdAJug6jMZ9P1lB7DHco+UGRgqlFuSj27O63i8md0p687P59GRvixs
EX8gidq17U+dAyPQZCWDgUd1QDQcETz+74BGiJ1YMbFptmAjvGOYqoi8vBE/KgmG
vbGc+45lWW0kIfvvxLuwZIdPsnMGg+IX1MmyQVdtllArN2sQrk8FNUuF4tV81ETN
SDD71tstwNxafCq70xEXEaDHV1r3Qfpwe9/WJaqjmaULUr1C7fopVK/68FIKKtLr
uBF3Wmv7cm0b9j3sTCA7C7cfpqAcffe84vhpUiD2HteU78jsog+UxcQ6nPrhAyI/
o3yaxHcFNj66+iwQCw39pdMtiAWoJr/8Nyk1fh4UNAr4au515eSJsaDQhBeArnMK
81Vzyc80zRY8ZfWLSiZOadPy7d+2Es4pICCVPjzb5bmNYIWEeZE1m2kpapo4FvZM
lzRnwWp+meixaJ7g5XwidgcFTCcjqXgPU2w4Cqn7B102pOqCnd/Hfp/iy3tRTgNB
z+7dyEZXkmyhrIW85nzPkFsV30LUGogDY0erCl1AWrwtlMxD6iKxZ4uYDsfMhAXM
WDImmyUwgNJGarPQByYYnf+FOSOA3Q8sYFSdfFL7Ulq5etSxoOyPpkWWZuf9/G+v
3vq6bkWncbJk3VeuMfm9z6WlSMcw6vdWNsW5WQdYMvwjfh6fbh8Xn3O0w4IylpFk
DVT28vOnTD1PuBpujhIuduxLXYwTHIPoIgi5ajjFWZawMuoZNEwqBaN3YpM7PGaQ
tbFIBy8Vcujy5FtJ+zde9mYAGT9+l55hP7xuuy6/1rbrEbGxo4SattBRz5IPZcc9
Jc/3KjljF4XrpgWOyxA67xyXEiAoOhwduHXrDW/5iJY3oNLTUM2EuCGdZnF6A6at
wWnKgnlQ5G6X0apPgssU8H+P7xRt3r65+3Se8+NOUES91nkH1FSd23F4+bczwHyR
M9wasqzQVJ2iy5LK4vsmZ9GudjBXLHhWSfHO1HPjuHqEQMn4hXjZniPNeiF8CYH2
2CszFjg2u/p2GDYJuBS7DJYXye2cUlqFnLJyWpGEn3JKUYeCDx8B33/6LjHIWHD7
rSJyYozd7MEFakaLmrotB90wjbS9qVA/LAKga6zgmlMVfo5d2CX3zCeNEHBiVbVO
nv9r8jcj6AqjfdjvfpVr+mH1FwtbY3VK8mV52hhSSXHobprpf1UpZxPp77VsJ7IF
Wu6/AhShYTyhYUDeQfhjdC9bM5myv8bINP8gzcy4/van+inR6aFtXgqspEfUx45K
Gj9k1Q5iuwlNonU6CuPTYhU6A3TuGK1zmzkVW4rMu42iwe1OK3M7rDRPcckiHs3Z
fsy+U+SsAiFDhXVDwkAMYkCkzAdPm4IY4s3LJR2UOA84AVGBhuFK13SxmsRYQL2n
SFoz6Ccra21cHYb/fAI3tFjxSoSzlXJZZ2fgfcCC/oK9szX6OyrcOgkVxUgI2IH0
fWKC/YRTvcEBbRsjOKPhHet+oCl4JLh1lBtwo43glv1sCIkxrQKed4SFlXeIXNh/
UQIgHZTWx1VRIRDL5fu9jEqwsGq6PHsOSDCcIRGnIyIRMYIoTAZ4a0lwH+U3ZGpF
eDUTpdk0BtLzhnIdmMaV0ESEdYUCpDRPhy9WQkSazUCer8yk81dcZBgKEpGs1v9J
ou9ih6pDvGA9GR0FOZHH5daFpu5wrlCiWOQKD7gt8ztrrWIQSTaN8niWyJtlecOe
6PJhlsggTQx5KqI9+YULL/9UUYTzO/U9CRRynal21xv+eI607a1jgGHGPT9yw3Pc
1M3z7G5kxiXKsxl/d46MLlBsybOSy9f7uHfu1Lgrh3nceYCV0ziFj957Qb++LW17
RFDHpYDwBSt6Kb+7UHwRinkbpF4lp+9nLlAkN/89PI9hY+S7oZjFo3aHZydykvAM
4O8TODpF4TlR3FYD3qA3bFWWECnaOgOflqvBYN5ql8UD+KMH+0svVwMpBEta7/yC
307MiYr5camd+5l8Z+Bggsl5zQBnjpmurR/QNxQST2XCMnwuglv8gw1hTxqz6LYu
weoOuAoPln5Yfb6dLT/EHXioXbMkCOc1a3v++xt9m6Vhk4NR3v50topz8PYkc5z/
74ypatEWTnyJ0CVN5rA8cDYZdvwBnmqxxsbdV6Ns0bA=
`protect END_PROTECTED
