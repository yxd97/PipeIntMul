`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lc4gZr9E1ISGPYdl3/K4cUuLHAjg7So0t1qavAx8dJKtwZMymSUhoJ2QqS4dfbj+
Q5PEQQh2mMknDnPZYbAtHZGdsOiVdQnL8B+bYeRZEqpIxFfBAgi+DteaYgwqIft8
BhTLWoeULsKOexuYmEaiOoO9QHkTehLMmzSpj312vQ0Qbi0xQ+EyVpT0rjw/xKZc
GuxzMhV68KwkSV0Hh4NDyZvX86CnZCyqEby8PY02KoOLIqeW2h0E87dt+mSBYuzI
qxtANyLP2KaO5cbHSLNaPth8/JQlKvY6oE5QnMgNuoY=
`protect END_PROTECTED
