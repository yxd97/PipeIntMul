`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cnAuaeiEn8cKQGG73d1Woc6yxGqDJlSFnBlRnnzdDDU98gNxDweezpCg17Dd93lx
lib+Q5o9QAGEbqO9GP/L0qRsbLlJf6RYb9cLf9GplVRig3HAfCwz7t0LHywzJ5if
pz2/8ntUh6EDhMB3mHhf+Ysc0eX3Mx1ZZg8wuwrKM7dSonk8Tddphzy53eUhAWJ7
3e0l67ojMmCH88xqJYptPcWMmTlsGA8+N8mzZ2M5oP32xUVMMYaOFpHfNOgjPtY7
gbbqHKBEhx+MnKfsrQgGVH9NPQgbw5WR+ySgSsr1SL3n1jeejXRARNyJb9vnRcTK
3lZUVXO8n3g65E5LheBAxPVG9xrrq4hTirYFndrX446NkZ/iyCDYQcxaN70qytB0
4IyrxE1rZpWAvaD9i2zpuaxVMiD7pzFspXtIqn+poaKRg5RQJpRQQnCM61EFzzGZ
OqAOCkxYTGZSP5EJwBAzk7+iTNimxSJ2zGIZMsTx9yQ4CrpBhtYLcKmlCb3rNjsz
k9IOKUq4P0A0ZwVpeQiV9iAruM4XML9dIkMhZVTqyBMi5q2FqwTElygnEd9c6+TN
OnbQuk/awAA4kNQcKnhYGiKnlKX1teUtcI078+pNuqkcwjEnS78eWVsErKzfYyYm
b84Gi6wfdu8mtNqUXgIttsCVPKU4p8vpdKaeu38Ad3sq1+I+a8O7sg7PbFclpIun
Luy36UIM29HND/Iuq4bO4kouh4Xa1nNpzH2XMk2JXMtSII6KXfGn8nUpAuOl0eUs
F5XnzfJftfsNU6pGAwxHgKmhO08vQDHuKm2eimhLzHsXTq+yvVqCO7PgEvK2VQOQ
xMACqy8bygPduvzFusVbHVbOB/MGUgcfwbm6NL4HPBQjewQEdkQCwTEO78eeDmBn
IUU+hy5xepgmtuaMTaczNp6JxTbcs56IxZZwD4kuNCwUzk9ILJG3jVH4GSarbK27
`protect END_PROTECTED
