`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
juVpo0dUYyJRz6y/xxMwg91SoYUw6tQh8HcesQ22xLSzNv6/5jcGl2aR0aQb9kT7
3HqJY69PgTR5d4rTncQDWvAC6HUT19PJ35ag9mlTKuiQSY+UDDLxDIQ2/FG5hW0u
E2S1+xmCqqOAFJ9plpFEJww2yN4f+lhRXSEjhoVeTDBDMwU4ZhsuTshXnbwHQz4w
PZuBTefzPTSucjV+9EAP2PxRd6d5wSyEkiqD3iWiDwMlDB/WtVG3gDeZxuctOPjo
MCKYkcHOj7vKpHdgqORXv18CvA8ILZOaabmzEN8872i2AiGnbZVQ5HwxLqRmIrPa
qypefO4chT6jpfkTtIAoQQM0bXaruh32brDty9F3kZO4d8hSM+AXVX7jWv1PVqFd
`protect END_PROTECTED
