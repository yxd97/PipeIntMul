`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9UxxxQEwNW6x2oTB1ADl1IK8UDRCXHOwcj5/1b3N37bPDLo+Au3hDz4He+e/u80u
wpMyCIEXy6SzEFnQB3aBAFxgV0mWtoBu+YGUqablX0fuAc9mZ6TW84VkJAWDJel2
Zs9sT+WW4IID7HNW+O262J63z3Dc9ZKYLRjE1q3wjTjamqJG8LdZFCRD8M1ShKEz
DTiJdmHP6tXffTQijrl5C+Y0JPALww/rfUSzUIzK5GBuaLsU7AmbtaI7Z8pUjP7u
xFmUiDcyInI26c+2wZE63TSqYKK2CX+07HHDGOSbq9xsk6MaDAguT4KcNSgZD1H1
Rd0uv/d49AX5apUI5Irf11LpOne1mlUPEMVL9Lgnn/7DiehT+nriUckPvdGPvfik
b8zroP6oog5WXfHUSZ0AuvmT6Mu4PDYty3yKoDN2e/1c9ET7Y6GFN32ljeJWD+KV
oKiKU/6nbrGYm8aGiXGVH+65QiNyoHD9XpdjSXim5Nw9IamQ1yMCQ2vxqlO2WEUv
SnDg2FtcSKOJ0Y5KWpnN/Pc8+zZIQLMqFTVadUvWarNybtnUErhwS4nO9KtgJFIC
N5gor7uDZ795F1nGzu1haWbIOkxLBcqxSYEzqaREK7Ula9zeNxZX08XtTIVuO8o1
zIY7OMfhmtagnPRQJLLwabyGLK0EsOVzkWWlii4lfRvEOQ/TmeMqbVRDUg/CaQra
`protect END_PROTECTED
