`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kOLsV2vI6gYP6FNX+eaOTX6bc8rxRyVVwz+fUSp3Vr0QHBuF4a9edJQ/w4h1Vbkr
9KntXvdvcJVsTCwroO6nv2LIuoUs0c46NQV9gf0UZeIQQOQ7MAtZlawPQM8xMsPd
vD9Y9Qz2G60+uY2OR6INecZ+tk2hARwoHNgjWMnjSbqnq64ftYjoW+YkG/F7yXLa
NBherAwJDWV2h4lJxirTtZafrOIAKa+lEVfY1FpSLVRyKSNshdsZW+3qN0z5K4mK
eNocabEc8WEgTQL3JkERXEePHBlQou7G2v3VhveK50ITo4ktYRrzH6kHHVJnE3Hx
wk43A+EfCpzW/HM/T8/VbxVfi1eepWAXG/lfBwKgm1WvKza9rkiaSOzX+yF7fRoi
qJ7in03nCd4JujQuCEXFJVQLdkbzzgg5D/45O2BDgpu8nXHgFAcXz7UJL9oyoQs6
miuJJ1pKfKhRYUbqlKhIkMt2KVs3oZ0zxMbq/q+QIUrV52lt0k0vx/Kv8Aco38J2
Sze4SXLO/e7y4H/1HVRSdxhITgljkHCLU3vr+MhVaa1cbxVOYHhSZNWYwz6db4Lr
p3flQsyWFojfh6LYxtbiZ3N5Y5gbU3spRZevAM5+pZsK0CshzkENKlydJAAe7uhz
sXF88Uxp9HipqbEXG5Foj4PIFJ1+JbAXnCnnPDDG990xL1g1Yk9TWv5rnB7F547L
`protect END_PROTECTED
