`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LyrMWvZB7/CqfXHb7td19yq9EjhlD5fAh4VtoKfqg6kt+KyFU6LoX6ovoRR9C2/
CwyUiiD+idvM2xNINTiiEQYpbgt5Z6tgYm4uZSOt+07WTJw1zCaG23vMbMg7lkvE
FRGGRsb5AiTMKs6Svvdat9TnITIpVNC98jx4QvKic3HxEMJngUOcZf+KOd6yUgbq
hVHnXt2bq7Uu+ZDJqCpw/6qh82o8S02d22zFx4y7zi0O215shYmft6L9liiN0DQX
oTkeezHEJN7Lj4aWqA+kibAXR/fistH9kOz2pjsIOXc3uvGKW+Uw9zd4V73F0ggF
2N9QJUysZ0yN9auLx0GghLNUpJD7OulfjcGXlC99m9eQV9kJDjp/pvBfvBPVU1Jr
PV+6JEoHo0Z52p4fWf80NA==
`protect END_PROTECTED
