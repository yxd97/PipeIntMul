`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SSmLMVfZxytcBlgqtJrbUVNwyyEzLwcIM+bKsoOYDU0TckVVfDZ3QTt1VUlleJ9y
1BBpQYysqjd3r8ulTFeb+uYlpIGPAajOu1BjQmzA2vrb8FdIjDQ/MAX/qMNMPQmV
hTc8Y13JCkD24b8np/ZeVVhm4oRVbOyBoIUYafVGkgd077WSqmHDBiA11WF1L3a6
m+F3eWtMhsU/9t1Rk0mqAie86TMc6MB/kXd+a9K2c5/sI68yXF+uvzegLFtELHbH
22gFODUQ8A58rKHS3Ogns7/eAaz22JZi4qrcC5MYnaPDLdLlTdjQB45ZDblU2cCL
g90NbZn6Y6aDxdUgrvofzYnZOqeEl7zPsZS0JUrTL5uV5uO+qbnRRi7ajdfIruPe
LiiGBDbsNpxleSFqaS7FvQ==
`protect END_PROTECTED
