`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9GiNNgo821lZ/w8j+qYIqI94rfmnF8iVMDWU4yFD4pJ2lZ/kWMax/+/AL3jPWT7
mmHvRhQg7B6cW3MWwaCA24Hebs0WqAhUhpubQh/5YD+uUIVZrDYYHnz3EQ2VxGy+
P0qhnIQ2N8jODfVtFS2EGnURPnoTjRX6L0CQxGqJfNyvUb+m0iPqVn91/tIrzyp4
/jOZU/3Kj1GAqNQf3oVHw9Rsam40co2GAA2cpqjq72FUesq1OxrLkfBhnwW7gFVO
yKbFYkAZ8CrcylYuqr1D3Oku2rpVB5UjeEU96Hk56EuZEDI6tkgNizHb+xqstntw
HgNt+s84tfSsTJbDXMHdbR1ACJPe5YywnI64GUhwTNzeh/eZFRb9/vxQXCOEMaPM
jyHAJhmgAoTqG5wSqqXBvdiKbAKikIsOW31OvdWrB3X2A8aIu4wzkDlyWZu6bMca
xJw1oDj9mVF8MYo9dh93GAxitBNFSZ04xj2HRZ9dFPxP1qUIOzSHNuMRa8zZ9j9A
5bBlvqmIN+NKrhFvcliSIV/NklNT2bzkv7bNXdvieLQ700LErSt0OZ7S3YfGUhWo
J8eA/A6RDH7E37lQqxFiUzr5WXU70AlWuftGva8xPuiUuD4wr71AqvM9pt/cd6e/
ZrTtmt3FGEki8taNd1dx6CLlQWDagVYiL/wFrsrFroqhE15s5Wrq4KzA0jlvmu23
M9gj9Q7Q+KHDDaoRlAJttnih4Jsmk5SBPBoulVNJBcbKLw467nTxzm/jGObKDC7V
K5c1uv2fZEfgwiuBGdGK9FvtPQEv0wjBtsMlqe8/L9bHD1awpuCnnWt2vUcNqAy3
I1vJvxbhBXFIpfFwe+AS24WxiLoNUGpkfENT7uftvYg/AOVKA1j8OljN0dUKdIIC
DkagvgHUWoqhmKWzKHChaB1klzrib1CcfUwRlE8YGneg6R8ECmiAekfZAITvyttf
2+CNZMQcDUMYhGglgITAcP6PxHkycoBvsNPvHfjcwlJ3N9OrHbe3NuCki0ZoILMe
v2uYlY4fek+7JlYmEPr0DQ==
`protect END_PROTECTED
