`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IYF8NjUCGpPdJufHxumrmKRUZ2pBbKbuqYcvlUFvx/VjeUAyu0XPkYMs4vJ8oe1a
2NiaYWTwAemapD8oJqmDlQ7eH+Ru7UzBEOmN/i0TUTVhWH2FqSeKJqGYCfnmLZd8
xpEXqIv9m35vtMgn4SjDYSosXFF3J/sFDfJDs64Iz3SaqPuhH5yQe+P3U77AHDcf
B+VnLtSZFBZWXIzMoiidtjEyshszp02oxe7ydd18aG0IkiK7S1f7w1hket455WOF
XxElPeoTceih2X/rkwXkITXl4iB+jXGK8kQqxLanMZJFwTD4ZhHw+ERTX4P9AS45
vKYyU7kKYnb68gAVA9y1gpkq9q0jQAI5NArsZJCSVf3EsrKGLWREBZhAdwgNzdHP
oczRfXkFGCM+1+hrG3kIpux0KO3t+SX7+7cMr38HgmrKHKXYgP1+e/7idlGTVqMd
P4CC8PmQjcnG8GGANGFPJxSvWqLKryVSYflSGK2DUxWwEGMuaFQVGzts+WBOGgPc
XXvq2IbTyitOOvGw3V16RVSMqQLcCnrjOrR8+fGI7Ro8gQzbSydj9IAaMDPNQfqB
9HNDVyRi5cUpar3CMC+xZ/5YLGx1ElO072AlGZzMIhJJAJ9DMuMaslJ93dKnJ+0u
bEUvYR8KE+N1FNSNf7LcHm66AMgknqbHQA3SMCTicAKn7cauXcJCR3hELcFDiAMf
Wm3/jXUW3k3gM0IwGLNmDrs/xN7gH1/2avqF1SeyWwGrKNt4kuDjPIusYy+3LQ3a
dk+1lLqUmxLrPB0UxNels0R/bn6QwSnfoRhESAEAD1gRNqQxfFaB3ZNuk/4pw5ZN
ggyFJuIhhLA0AkNFkXOxWYF7pCBBI5FxaG2asis6uguvyj0lVMOzhdcvaXC0xPnz
jmkwKu7Y4+QQr90spd3IgfcocO4+7RrLPPIzWTqR0GylTg/Z41cLH+WFHBBYgwLw
qi5nf3/DqhhAdZInAF0vSRUyKSB8keBzSAGjShj58wnhazG36FVjM1/19hoyxmLH
5HuDu87N+s/isUObbAU5SkNXpHGmvMjxRKJYhGRAUucecIv6KCqAA6fZxdEtGujk
mwMvR9KsTYJ6IddZY6j25h8yhRtWOkLrsgqnOGDRpTFXHcniloNciCrrcRkgoQbJ
p/i60/tgPoVpTc64eG2Kbdf7sJSBk/5bCZNWIpFjWPEG6vi6Szx4cGeOGGT7wGLW
/AIK4ZoTGPPzSlLZgi74drA7/sF5lWGT/hTPN7jjC1u4zo5OfuesKVSxcHFZ3jeX
G6tyN8/o653XuVhYQX/tv2BZ68jr8toN0FzDt8jP1molT4jpwm0S8vCj1mORU+je
Gu65rk00BdljA+MyXuVF0FhmX/ISSklaSpXWCBoodvP+l/T8DgSKVhtpQrBdHdhX
byMYyu3dqDu/yuWtJnFGBw==
`protect END_PROTECTED
