`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ulVpIv+eGwn8K228nh88+1Bdj+najXm9SZ+s+6maHH1n0Cz51pMBe8dk2uLvmXZ
syOBAnsrQ3+/BcsCU+Y+fzfaNEawOsPFGvg7oY27rRIcuPd5sGZ31JLriCBiavSZ
7sHGb/rk11hkvTMDo27q+jOeYVuTQCHF542DJ5xqpfTaAX+4+GuqI3UaglOo5Vrf
vgMoRTX/wqunYSV1NJFVzpjEE307x4gv5MZPFcz689g1Ht7Gnr95JdyHKtYVnK0q
hC3/zS7UI9jjxnaqUqdefppO63V/AbOJZl2lqRiqgCRGerTGQqO6dm7xIG2c0zGU
FoMaU/Uvf4kNtXe4IF8RWk7PKh/Le0nX5q6WhbIbGL5JDti9f/x4nh7kxI2ru69Q
L4D6QgleiN2jD67xloKa/2SHwQttCL9wqGLTyyFO6R4RwwnNa0faLhw9hvCBAG7h
KelQRrZh2WtrToFdQKnVLcI+QiIXBWNHqc5YrT5yaLiuPiJBYqmtFDuCS9usdZzb
eoIyHh613LqVTay70TE0gVDrkAx6d4yQiC0sUeXkefQn1CjCTiCKi/yqT6duPZxO
Iy5OtxoJfLv0enNxlhc92ybENe3DI0TX8iyijlRF/e/fFJ111KEVuJOGBQatCPln
P2h6weQ0WcOj8hX/nldCsrORQlKibqfsrVFTrV43L6pklNBJoHQECV2eK2+81XTW
wtk6EpHUJBdXRDJwC3QiRtVvv26Er3IKNdEuddGIhQWKraGjg8Ch4sfObJeNR9Ma
bLhVW0HyCXDI23V489k3LV6m7uUvcr+Fu6w72Zkb852gpc4ulNzpYR68ti6bxPWN
gyiKWPQXKG4a1zX+7IrwEWmayo947cUDABFRZ/Umaa0=
`protect END_PROTECTED
