`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/z74qdtNX4+lN2Y7/xIkIjxzylJxnhevZAO9FuypMzjCwAe9xWuLKcLYVDByKjw
v/TP09wv6LmpVKxm98U7BVAbcRK1GmAG9f8SoEwGtuXY21IJ5B7AfN8+2O/3qxto
ftDYg1V7NbsIuhg1Vt7nj+BFwIWthlews+C1zvbDPrfshmMuXZ5twSLWOjXRhK/l
6tmB0UeRKFaN/1TrzhDhn3TVoYStWOJjAayVoUS7NHml1SBoLeAMQTBAuwWC4mPU
pKhgnjxe0wFPEreA4hogvBmyVQjbatdcs0vHyLfGwv9UJRfd3FU8DTIvHCz3dNoC
cOSDksNv3WCofNGiuc0Udgfq0yx6B/ZMGmuqeTpKUoeFT3Dj/Ly1wqE0lKPCPH9f
eSkOfj3CqK+45Y4R1IUw7jaUgOYQNkZvYV/ypJHsFENntF0ymo/AFg3lyZB7uudn
jy4QT9gp3VlrlUYMkTB99049lpWKwPdWLnUHyOkuthyCgrABa/QbDWB9uQIPx10d
odWRC0AvQVS8Uh8JHyape4kOP9IaaFkl9EF6vjEKPssF3Lv1ijujbPmbCVoafVbB
4It5rGLAoaQd50SdX3+g5BrhQIrM7tDCoxiezl4yOU9YK5qTUrueZlrjq9F0N6I0
QjuucBgCrBTCDXLUcz0WAmlZ1UCHXIV57McIxIrf+1Dc1iGiWGQ1UgCtFBD054Zq
0wohqCy6sQRGfvGK8OpLLgkB914NGPHofGSXCdqurXvSBkYCtV7zAaxQ2pqyYe2+
CRzJCxWXSE6nO6QWxFNE6psheiefPBQsjXPPdqy3MTO5DcFu7yfVUwi00bhII8Fc
CV1dCx+f5HOr88Zk7GJEZ5V12HkpRlZw+WWHwDJG65en4hdKrssyjxX2yTKMxgap
nvriYyuf37dAt6siPl1S/vc7esU6cMDhtjuPVPlXQBA=
`protect END_PROTECTED
