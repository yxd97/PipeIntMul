`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3b7QJS3cTVLeHC/Gmym2YtEPOl41KDLDsTNvLsSW8hKavItKJfrFSmh7zZoTPWO
0S6A3QTo62aLE74CWUkVy+A/Bh2uLtafsJqtGFkCiJTNna6J0qia5dDiFYafepC7
hyUD2IVg+tpAw8aHAB36p7/SSGP0PFPE0nxNL+gKOI2CMG0s72ifFVps4qel3pc3
VZzDhL8QKUfWL6jaIs9YKgumSkPYLeL9/ACCyUTd8OjY+eCeKZh022uFAqIgKg8w
E+AoPGCJMN7ZmYXGi0Bdc/1vaTPpsx6QawyremP6Wwu7wqjnRXQtyTth8btgxgxt
HN2nlCxYatWTQxsgjfD9Cjx2fLQLVeLBVpaNlc+IkkAykxRRT/EUq/t7jwZWppZM
iBk0Qrxn5WfBp4JngSqgPhtIhg1y8ZUqIxp5zUJtCCtT4tSL+G6n/j3Wuq8JvjHZ
QesmIS1ZuoDgcDfu55jgMxz6xprvGNQl56QP/JXTwq4OQf/+EwSvzPxD6E/TUw19
9jQv/ZXqpx2IBZA4p+k2liqbGrbSOoN+BlmEcMFAkRPLd1jYCZvVVv2sJ+Gx1MDe
P5yT/nAJz41Am1uIQWYQ9/5lYUC9EXuUiCnUZ1P0TDiyh80U28rIqOde+pT/xGKo
afOhESljcNbtvGOfQ69hbGpVBnvin+t179YvJ9GqMGM=
`protect END_PROTECTED
