`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YLva8XSZM40wrCbcyRu8t9dc2ETjveu3D6P+3WhsX7KA4S1Tf8VEDHRI5NBiX3KC
KtPHoCv7eOB9wJyML3XFMmwIYOslTOb5wDBXJHqTuahe65a5IC9uTRYLN4klgh2R
B4rcFlBbNRQHug8KWZXwItvilC9kukk4P8uhLLpmDStCOVNur5DkD/pLOpNlA13g
xYlIQ0Rsw7ljNcfGNwUDLxRevqVJ9qvoyte1mXTxI67zdguSX+hzM+Oe4YZZRgYC
rtV2jfs+N7kI6hvsRuKddTryPd2jrPBNHZe72OqLsaspLh88uLww74e01lLKvVpR
ShQK7eQJqZMlgfe2hxrsxUqss1/VPc6cJD7pA1q5gDo=
`protect END_PROTECTED
