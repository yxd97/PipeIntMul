`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCEatw9mJb5syRB/BCgOGr1iReMbeDHtEnA0Yn+ak4xcfkto+6fZQoPcBBtDad/O
PATlaA4YALH/tKi3n0QvqChsSpZgmv1iPxFOOb7KlGKn3mqzUlyLBjWVOXdpqFpz
AJJdbHHyZfPq8kOsc6pyIUx8+MqVM29QK3UIeoV1tNuLxyhm1eYW604lmKLriOCo
Jb0ea8G/SQ3SvvodrsgGQkU5MxmEXzMr/krOchq7ajMQe2J0VNUDfrjoigMm6QG7
64W6FMlSljIp01iAsIRMxRUknfvV9cjPdKc9O8WZ/+lEYFnDt/NGCJiO5I+Z4PcJ
uXNVtcqKvM1LLo5HRggzCX+kKS7yIxNJNO41UynOzlAr5ibijDQZdMBoS+0CX35L
qexKLNnVgl99FSpl3AbTqrXj6Ei22wd+IUHFTbUarpGoV5362OddOXtI/6uaq9QI
obV/YBIXSd5IrOl/6qQtqOvb/gTiap5ivgStsFG9XXumPUH4Y8lQHtSvFzO0+63V
`protect END_PROTECTED
