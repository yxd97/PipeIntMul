`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jy5DfwtJidEButvVXdNOwEUeWDSQXNXb4N1f1k6Hmv3qr1fwJ+dO1UO5ylBH9nUZ
WcwBw+daSMs2MeZnwoyJlE6ijTluIDIpmV/XKREx7/Wo19hplLRVoKrvz6WfIHjW
fJbcBDrZW0p1NhdMdM8O3L11jJzs9zp9lWizy9xgt2EnLorHOkFlYMv5MkSLOyt0
qLCwg2YT+VVDsnfyrjaE3Omv2MmybFjqcp+nEIzfXBv8gU4LCLuSxYWtRe9IUWoT
6ReMjZC8YVFoc16fVdhF0yDY7xkvzo4tlorpAgpsVGPLSP4hse5DJBvAPqSRsm1v
W+AISCvlr9nFDPantROcqA==
`protect END_PROTECTED
