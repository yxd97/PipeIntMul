`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNpG25dTsfOKmkpWVQvCgG3SLQTKLPUb90YkUpK5wi7TxvzTM0NOUs1szUfJD9uc
fdLpxiMfv/DlqhVYjJ+gE0kKN4vA5HQLpUqPHzrVyYYp0I7hWVp9YOejcwiTK1VE
GRAdvI2IZNdqh9VA9OVBaqtsuLBXFUJKyh4aitPff8ovmXmrE7uBP4IypP8rm3IE
4cC+9t/f0+oL6Y34gTlPBwctV71XLUQxlzs0pdN0CNOQWwYepwmx/ebur/6GxCbK
Y+W62ppZZeRwacSyKCdnZqvzmDptu6l0gEw2UjLDRoWU6gT6t/hON9kFxrU7BHMd
o8wh5i9wsNw/gyx7ELiFj3yhN4itCG/QG/ASk4146q5d62hPUwAhgw9031FjDVwq
S5k/hTV0F9q2b7jE5ZJi0KfH/Oaene+ccwrqS9VN9sAW0OdrWxVzqfDKfdIuwk8t
mapOCNKILX4tx/897YNhyx2/ojH2CSkjLF/Kkbn9EZgKrR9XpPhpB2PhGgShp3cD
ctSyPFL19kFsTOBqLCA0x0Ul0SQERI3yRd9lXAyythKA0BRawy2dUK+d/RE8MG0U
MnULa+suIrFsgHIbU18abQ8aPKwajMKEnD1hkAGru7HGph1mFRW44O+28pcdhIhD
3y7mfL0mpp5aNI5t0HnjzOazgzWMSM1rfSdxsvolSdx18opPP0uNOTvAkt6va+96
Fd/LB9ainYB4+4iPlZNxLUnV9AUMunQOgpiz4d4/V0gf0LjBMp88azfUeJV/W39J
QEOYGyYjnEQKfnrJPOYKJ3QmFWuzJlviUPkIW5va0ublR3Y4ZwohQrmVFnbcX6Q2
JXpEBu2aXBLj7NnuWEnYCDDhoGEN0Zy8k726BIdRxx67qknn+ypqPWJHUWCDQVvS
fZrjSE/OpjrlFdxuRietA3nkEBoldEoHGafLvuOJCH03ksuohHDPB9dUFbaBrwTl
13k5ZQtk+uCWz1TON3nql20QTk1Q5E0z73uE1+08RVOAot4I0wUPaDXOjt3KlzTm
CjViowdzbl0POZQMhtEuzZscYZionc3ZYrkLq/MG7BvJpPAcAIbJ2S8IvehoVhca
/rFfwE1iKI9PDZCS+LYMcYyC8XTWR+wZhP4fFHCsDwycQC5yCDTAC5f3hmsrmsqm
MWnt3Oq74irmc3GT6UUwjlNWWcXghTodqaW6KRhLA9U6v0wx/eEZaYd1MIBRvWux
ORW2qebTmTZSy6/8hBQyzK+Jm2pU4LdeILyk0Z+HMzaiOH4jmsdUYddsG2A676Qe
591oZ4NX++C+d8RuwLrb/HAUyBLWuvkx3RRTYBAq1XxfM3S/7Y4FhU/fXgwtmVHT
7LO8emPgNEJeEDD++MFgkjEyvKI/Qvzokuygqu6UkM6d05VoQRe/ZV3uYCgAPnxw
c/JLtRYKvbH/HjwtkNMVC7jXBD+d/AI3FaOjXsdumLBufl05pAJ8EMD8Xk7KQGMI
j654mtznrqCj4v23E6tyDHyyJv8yEF+XbZaUSJTaQ9Of6oCs2QVKNezv6slsMm26
kCTgpkaosyXO7KWmQsEn/08oRGR6Pak7gy0VxktXuKqa0gkAUZao7mWGfvnTrZw0
acAk0PdPIIXPbMCW5Cr3hIUyZyClNe3/Eia3Dib7+yJqa6YBnSri9ngXX/Jsa2De
hwKjgSFSHQCa3cxrMnJcY5RlHYha3Ff/OAq0KDDbAUn4nqQH+Nod7ELgl2JWZhkG
B5i7plxtJ1ltupQ6CyeytG5yx3HpVhbXDIS3zret1bO8fcthe+J/BUCkLjlCe5NI
SupAwWUrsSF3DrmpQJtTdUF35m6IdTUOtU36KRtk1saNKjv3SWHl0bGks+jNHd4j
jRIqBtXRmrmnGkmeFk8qPdmVZchfVXelE110bTF7uCp9sZSGpVZst7cqFLaFsnB+
nxOf2yGdemU6KXah7cd9VSD57gNVyynZx0MM4F1nA0F235//KIs/andIcpl0/zXp
i5qwqfGP4lBqMv2vEqBt1o446ThKyHK4CJMBdR5s8lkhMfex9Istjm155SASF68H
UGRaotGyyhi6HoAPbzxgoWqQxeyJE7HfofKb+x5PwrWT6tioDQr4wBv2iIeO8QAh
dcluJ0RKA8VWPzZaHtlpozYmHAyNflFxLm3hHXerFqk7V0qrciErZWoK/J7rlpEE
ksWh/8Wdb9vrNNTyj43GL37qAqS5xMJ4NBiiQMx6o9qeecmvqcI/lZkHR5CczXqK
TjtvnU/CLqYki40H4L6q8meb4mv/ig8qQuo7s/hfvwhB7CtdfPV5IT7FRp5id0E2
VegnQZhEGyfilc/QH5Ir+FEo/NCfyLmPdfQS5HEFTZvdi4WVH0CiDjhkKfxiB54T
aTaN3IMFzXkyT9UpSep1yYJDoEnGXHj0Xzvg27bU5FZARdH+8OpwomJHd7Cvy1jG
1nyXBMeGNPtDG7b/wGRE4/aLo94nBs+fj3eZVRD97zLcT0HG7gL7x9GsUelUH1ax
D7xiJTL9RaO2v8NX8HLK7hvVaidQgKlmhac++63tdU6mY0W5sf3NApjr8eQCiA5L
bnH0pgJGXv9gEH1/muPfixtLCd8mVcFhrGpgTZSuKzsX38e6Q2VnBFzCRx6ytnOb
cFWuV8mb0lLBQNAQy8Hyy/eDvSTc9D5K2jGjl1VZdeCpa7ZbN/98lDgGLS2vIgIq
+/Tkea4xOV0li4s2NYcRK1y0jOVRfdqWNuX2H6Pet1qbtaFN0FeUyKBXEapjR8hy
C4xUl3ucyWjKEcSRGfGTw81hkRYA1hf1u0aLMI/xGeI=
`protect END_PROTECTED
