`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DkKKXBk8/0zc1erYC1h9rW8WJVvY+Qt9IoG7s++GeiouO59kIWaNTScf7/Yg8xuy
94nfwocypCrFiSAAx/uZjhyNcKWxAwZdsnc4tHl3Zyszu+xdk4wYrnoEcaIpRRiZ
Sb+NlbDkX9WbolHYpisyS34pIy+8JITa+327RdXZFDCoBfWV2s0WscIuQomxAoEt
fr4BY9+rTKzjL0Q1AbaSOiH/PVXKnXZVbBPKUIBrhpDhZLfwqhdGJ9CH6StxpEsW
6SB7+iDbQQKqp9an9isALM8GhAhnnYr/nXW+yUznadsiV2OnCwYGlfdoZ0BMMRyQ
BZxBv+ErUFrSTmF6J1DPU2zUClhb/ERzlpwRX3UrrDGlPBLHi4Cz7L6KFVlnVjrZ
Z1aNEOUOFb8G4giqZ2anuv3wjL0KFsIUQXW/TOr4kFg=
`protect END_PROTECTED
