`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Omm8omqVs9YcVDBKEomlsFq73cdetmciJiHPP6M00IH3OCeatJYpeFM6Tc26Nuu
n6yZ1qPvEFri5uN0ciLwRKKongz2OBR7FpqSMl+pAPN7DgDCWWiy3ixIAiwUw+pS
EgaueoCeS7mF/YQofERCbOLqC0wV1HQNjy/m5cGwSel7+FeeHv7wngsPvkawBHh7
T7QMQkjX4IgUjaKqglaWBh0+JiOV5gUC3oY5Pv/go0JbrLOqBaPs6jcftc9ggTyE
Gl59TKDTYNfGtEDk3neFoSE/tQ66GYgf1yhNGt9mS9WiTTyGNjaTFLB64ndTZXs3
Eu0s2CytqmSj7QSKMunewo9wNTx+SEErFyNMinTppl+vasgdoTmS2wX7mH29mTct
/+5uqDQ8FOhta5+jKqxeigkS5Pbosgg7ToBmDDx04M6qiSE+4snAY5iysZvUtT2r
+NdwM9tIdaGagk3gn1Hi7wcQRcwV+YShW34035uyX6Sy9kk85RuNk2C5cmVnvYf+
c+Xq9FUZHHmgzCt1cq7jD62tjzcB8akUNdBy5BUq4LRvyTNHTGlPGAa8gZcg13ER
3wdyr3WXyURlVOtPnDkhfxOKI1RX+y+R/9OKaNnML5VR1s66fWVqqozDKpGOQa/D
2zWSCPGB41wNI71yoOgGVK/zi4qKnqiFKCALVg7VZudV6xSzrK0rKZFoiRrBfTjT
FPiOwJ4mVUQdLG9t5EDNsHiuTJUzcokEwhIRhBfy5Vlfn8mGpV8PJzplPtxaYagB
mCzJJVzYSn/1ooOQL8QydGTAyrCUszKVfXVanPinPbaagVyfj+zZKqQuiGcsgA9v
8YgFZ6KAi2Vn1Gpxjs7Oqw==
`protect END_PROTECTED
