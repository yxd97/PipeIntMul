`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VK/OnYaZ+/tdyTZJ3wZJvFrfLIJhbSuEErbN/oIyvnYwRSV/ciz8rydikKxLcOkB
xtQr/pdGT6QFzuENoIV2uWFLVXaf1ogkUIvCnf9NL9dN6LWwk2zSNUrBF2+gLrm+
ASRBaEkWzLio4q3EY6JC9tm4fH/cnTNOhemfuZRHSEmkc/2Bo0CiNgiBiHHvB79g
A3ebtjb1nSRHI15xS78kzCsTUBYRrVBdjkAkOVeYYL3xpjZXWfMxjmmKdRZ3iZo1
bunXRCMbmkEn+/N9TsikVw==
`protect END_PROTECTED
