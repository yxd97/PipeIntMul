`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HQ/I8sx4XUDL8B79Nkb2mctJ1M/H1zeTKDALyfR9xk9/qQlt6PElNTtbEWX9mcaf
Id76stoKIWHiXOrIkJlaXen6TqIttfnuLWko1O4grgFYkaGXo8TH64rCJd8aPLO2
YOI7zPLiSbIdTfnOmn67rhJbn/46EWrrDQMMRl4mIeotq/LxadhpKq6Eugy2Tz3G
gvR7WZx4HoH50uanoCbKALgu3P3ODT+1d/Xxras9UEdyxhwDQIk5wa6m4YynVAdb
03fr3MT7siAR87h8TsCll+C5HCd+GBubOcdznIije8AWomgizF/Gd6mR/SKf0/wP
G0F/lcxFVQPysvyleGc98eyvFH3ioLpBvwNmVAprG11ADjec51449afrTaT6gGLi
i7LRicAgDZCywk8aQHCng4/W1IQtJc7LT95w8vKJi1KTZlMHhlBhHJ9sFZTHmXjH
WRcHCg6KffomW7cdBSaXjustOh1xgvn89tb8uTZXtxLshQw2kdOHtzmJ5Ys9CJr1
Ubxa/oDnhAP7kYM6ARhSiQmkwhx5WzZ/knlzeJPrhmyi7N1AGKvyD/TO5ieS5APG
jX8tm+Ap7QAwS4KWC6AsMcVmh9VQoHyIUKG2JWl+mw5VR54IHhRXvwgjarqsHH7O
tmhLahIULZO4kdSWsEoq2InBtU1qcFsFMT30cTHpi57/phCcYYSZkud7kulY7LpY
XhvVNU8mWwpePZhTs4UPsn29M5QDb3EqqhJb19ia45lSFgsdLDcfPWMLwgRDNXNv
IhWjeefaMa3e0ouUrnxJq1E1GVea8neHMr7MuAppnKAUA4B3DkOdlu+8T6hrk/9v
5X5dVRYrn/dGxU+7IakUpom0YiYag7/J5/5Fb4VO0Z+y59VAOVTrzPmneLbMYWQq
d2D9qilbdv+n+/0mSpFEVP6OuZI4XZCANba/tts8vLPytyuCp9ZRzt/GkZl1AZ3o
CWG2C/gQfhmKrJCVE7JXmln3h0jPGV2OYpOFm6nmT4Cxql6pPjdE7/4bTU03Atx9
UAahwBMVLZP0SsvpIrF+Fv3e431c0CPwPMgtTN4kh9XxIBQOmhCReIIIxU9HdU0e
r/wrALXQvtfP0OnSqOAnG6DcQakayO+45/fzkLbAw55naHoItSvunLe7KQTcau8u
4SHUOCjOXiWH0ROdcHnQyCDd6Ieb+/pSqMRtB3BnSvgxCmlOswJTmjqGDR+xrwp6
STctBLgGHQ5E3VgsSBR9tyjVNlNraGBs1OSKZYvGU7XHg5Icc6631KiTg/rV8Kc2
tCibw36FSRVWg9bV8JwKLJUcVvRzndiW79ilYmq992JxyfJtGYu7JqBrYriTx6rT
VMZkIQMENgV0IVjPy08Z9hJvkUqDulglUVyN1fgkGfalGh93vdOIDY9KGHNKyUuP
azIgECjcQcDzeW2znOyCMPJ/AJaQj6UpvU/kRVUvwgzgcuEbzeMY0BQGJfNJkIWI
KAsviTeM/ViQQyEwCyu3l3JS0xARBxIxji1qK/pKV8laEiTNrZpLPLQGDyebJtbL
PqUMaSyjfBYaiy5Lu8lXsy4ZnMpBiT/d8VprN7Rgsdy2V+7JfFZKArcnOI4Q/0q9
U0ed4Hu9KTCWXrq3XdSVFr70UfKluxSsAvhdeFUhP+KCn9LF6Wi4XumMBoHTn1jG
ojSi6qfptr9VBuG+oQXzXNGxpoRsljA1+Ga/PH16mgQcN4S3fKUp28foyq5yyyqK
rv6NezW/Ya4K6b155msDNrfWYUNvHpFWZ4u8l3PyHFZQ/f435mUhbqv/mROyMw3B
5CVv1XMqpFzopzso+sFF9n07xp/uJBLse6yFpqKqrhtOOS4QOT3ooFv31MzbVIeQ
/K0esuHn022QBQdEl/xdqKZvCBPJYdKo8s/v03qyR/3VlLHg9LeruUSHciw7bQ/w
eShjccPhAhuDErJ+Uph449mxCVvDsnVy/nSrATd6aPhFJAeZspTwtgoEPAo408Dk
VB+JW7wnn0rCQqr38D5tpF7D6AMTij9a1xkg1J/Doa1BTriK3mMeFLoJFWyR6C3E
8p84PcRpr+GczCzUKiDDwBRDQJipkHUw5tXPAQgzZR2BJmiuWQtxhhP2jT9zmU0B
+Psrs5oo0Rutv2cFF7Udk6oPEDqhrlKoH6jh98q9yVoAtNSSqUM6d9mgzQ0YhUkV
yxAi5XmSjGa92ecSScWBbIrJ7bImLplqY8Hu87xsZjP/aGvZlYS8+DEheOWzeSyi
inm5Rc4OflsYV8RGg/F7sIMSpwihKdgEyJ0F5fFJKO5LAD4Tw3p+jHRaeOV0En8N
UOdOhLA2yB3KiIwFMjcnt8Xldb71Sg3Y9xL1pZf5PbQjJYpXHYQEi/2KRL30hhf+
Y2u61S4yAT8kg33Ur39xTZadj/PoXA1mno6C895sugsBxQLhehrkVXXZJ1viYRzO
FGCS+08Yd5+OMNneMF1GSev/UAKfmKaf1ldrGoXV6pVZm6Qc+d/ykaWFJ6nH1Own
zGXOb/u++5VjdYXIvaZ3SOsKml7xtf/AGLOMLGM3XxlpVsHsjTFD5wHII0Ow2mRx
mWFSgk8oZeXL9SvGFfdQQ7S80t3fvpLMlYnGMXiiAGlQY3nPU69UG5xtbfMWUgA9
IIPQYo6FcL9nxiKudPKTtmp3UtFarMbnMvr4e9XL3eAcVqgUfW3luZxnO3oyEHt8
4DORzUAjMgdsZXSl8bM4PvZIsg/+ThQTg+9G5oGCb+p4rwsqQXTEOUZnwsi7GeyX
f5iZRym2sdQ/1cdWj2xi+HjsqOM5nHkmKJv2YMeXfYOXtzlTB230hxApql4Qgguj
SsPBrxqncgcFfNY091USGBydbpeAdCh6c9vLciwEEF31DK7zpCTTW+sP+zh+vz+P
IovohQr+t64mXoKUtWJ3CzOes4SoGNiopdpbgKxLmyN9/q5V9d4ysITqwUvi1hzB
ZfSbeqkcSsvk4VhcpqDl7HVLGP3DLNm1mtGrL8ZYPDCqCZyWbszQdUnfquxuyyIi
XqkiBDkwkJN84byFPVbSKNuE+Fxy4dBlRX5KzaLyGPzbLuODfnW5ouYqX1B25leJ
xOjMzhx096KWiXHsCG+GejHZ+o7IpK60XtXs42zM2wqs7DoVnq9sNDcDXu/Lj8fr
AorqtwkwX6UVMBpZvnzXUv4kuQjI/v28Q90jQDZHjfKlnTzWs5NPTFR//uU7r1Ew
EAH+iq1XNwTz9gTOIsTOG4TxYLBshOpTomlNbuzY4XTg0QT48Y5zYu9SEtXxAw9a
Kcp5N2nc1Q+kclkqr2Oj5rdHeK5siwXWiPiHZn0IAowbFUQlVjfHxKVccbIUzX7z
Pky2A11x6eoGImW53rNLma+ZrwtjnRVrWxWnPjbAmwwF2gsvte7iDdOYbzlzEUxe
z9TojCiBYj7ZcdUwY8a+rvgG3+zGgTkPTp+TjC8Ojqb2hLKqMp6tHZjFUDadFKqz
Ov2/vsBgJQ43cjj+znKHcpFrDG7OFC8NtYMucXI5utTAZ0fcj4y9LnflMpiKqwsn
CPaX4vwelAe9u+4jvHPg9iJrHULEIQWdaEdyMv6tlfKiesv+IAsjX41V85qeM+lT
CUGjr40vUih0zG90IHPrqm6jru7SBdl4fi448rEUYuB/oWzi6bqYEivJJGT99JD+
8OjCOjsO6WNqvSo1FOiDngxaUd3NGtS0Fm4xVo1zcdAKprKrr7dTl2MwSeT4M2n8
5zeNIADmlNh5PK6ihDbJbdM/PPtw78PgHS4pygzZD0/97CMg2KU0TwlzW+QYPNFP
JV+zoQ5IfFJ1su+S57OTvMBmxNIySD86dLsP08f8ErQf6bp5dH6kW/5U1XJ+0P6R
VZMDKnonPruSdJM5cXc/AACO1jQ5Hy5/5zVSzhTiSa4cCGSP3J5+tlZU+6E3vyvB
w2OGn/ElwsIVpKpQ7Iawj9YTAMvwGFSHkim93wl7QUN9Ft3kSKti3DdfpgiotMAU
bpk/dExIA87fYy7ZWoMnR1BKt4BgYF1Vs+pXkksSWo40Jm1MPEiAVk9th7dChv5A
1sLwDkj2Z7i6S1GXHSXjHSfPrk6sjb4on1ARBCCbOdTwpF8eVdIapNhIXrLrLGCT
EUle9i5tkYJFFd2GzGdKwaOC4mM+9KEJwThmo2GahqMqBLoqSD6tcXu2ZvNJmM+U
7ha01jrMSaGJa6sg52OyJboDqcOKV1dz4LyLfzFUCkVkDCRfeUHdrgtcxz3GeQR6
BbZua5nwOR5BnDh/6Dy5gQIq/NUHmhdTKPjt0Z2kb2DIaYRj9JcYFTnsgcTvF3hf
M2HKSliZF5rx+E7Njex1toDSNam2Wbl1va0JTzI5rzgDDRZde824q8puNzWHWgJI
sjeQoCiZhYd1Ui8gTy0FpWktX0Yn6CARALf2s20DbJT73nfcgbaytmuaW9+1Tn5Z
mjdkYnJUVBbq4ioyKix6TVpG5hsd8kHVVKIfxTX70myUmAp/5MWNHgdZR4b+WMQh
vwqgl9dbDYCdDfAFGwRinsATDsftJv7eyYJhEVmgRofYsVkDbKDXaxtgl/i7JAKJ
PSzMb+r9+gw96cqNNgEGkNgwOl/EJIqGSU192UKdweMMk/ppT3LAgebZU0CIjqle
giuEkb0UVCrj0sJLQc7xgaCZHyfYVuqVvgJwViIlVSE=
`protect END_PROTECTED
