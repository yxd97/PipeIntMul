`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evRzm8aKp/3Z7aj4U8ElINW+rDtLz33oUd7mMqW5PJ6m05Q4l9AiCAsCi402H8Ks
ZVMOBeU10EZO7EuOSuyGCR4ZCY2KaaO6Z3L18kO/VbXKVCrjQbBezGua3fyHcVyb
3yk/gtWcJrkrRS6DeJBhhzN2XS+X33v9URx8yGEuAh0u8B93uCMhk2av+B4Q65ME
YI3l8hIK2v6gjh85yLOulTPOw0E7MKPq4/nB0DcdJPe5FfgIIuZla10gb82V+WFX
3cKauarVE9gNHeOjXmlhIaSiProEsnzihYzi0bJlUAWOsLwX29xEaRZ44NZIjmyt
0dX4WX0XMHobzWxsmU8XEUnvTbarx1U4PnaN2SXPaWLteVc9uetOer/gEr0wRQfN
GSuDDvW+WKWDMBY75UvucWZLX1uY61zGcxk4iBBfytDgTB7eQXdwStukTtersMvh
aFQqsW0WsnWC4aWc7nAA2sVxpTa0U/yXcfxF2mgzxxXGk55h3cKlmTfnzSKkVICF
4H+N8BFaqaqqHxuldBHcWlSXWFMEBuKo1JV2H0sxHAI5gI3BwAizYyD3FIvNAzbT
14HkytVGgpXout5I7gNTPLNU4MtIlmWLl5J+tBxmcRQ=
`protect END_PROTECTED
