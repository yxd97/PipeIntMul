`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rDVrBAaxQVpuXEg4SJbzlgyZ14l172bL4Fdy5+RX67ZuouTOVcLiyCgg48UyIHg
EVBf54HrDqHIhXr+ZMyZatux1QfkMjLzh9M0CswPw0tcoT6jI4uAKCKuxyV7lssL
n0Kgr9EkIqV1UKzKOW/AX/3sqUOus1+9/kliLyEZbt2iKMle1q1sT2tNMxkvde/7
c6VbQ5PKaAOXnPUejn5nQZbNB9nP2+GvlbGTruaGJ5gUNaZrMcpIj+blD6hEnC69
VR7tlbvF9oo1Hbm47NpLLe0x6BGVow9uVfYclF+z8+axSExhvidQzOLNrpbaQmE5
8wsTnR1N/aVIMtd4p5Uep5c6Z9QqjRRCMZbX8pledUSQ+BndAiVwUmpzj/XgV9Bt
AoA9Xz5YGBSPLINyT21snwYeo4w0dehdPPeO3J4qHLvJBw0SL+ruWawHWsiHk2Al
Jcn/9oZsNnhKsS7O/OYOvz8l9b26GZEEx0x2yFUMIzJrJVzBdeqaKr4q482s6dDg
PVZ6n0zGdeA7Uft8D+SAdNMW4eucxQPwiSoDVmUB3ZyOtwG5IlGPX0aVgEN/julE
lVGPqfbcxNsfwgP9OsK1kLhh5AkN/N1rz9DVioSXqunfcMOHPuJ3YCDNjGCPL1Cl
NIi9WgKdKFp2jxM3uB1BzWkJwfG903Vsao6Z1WhvoPPfaKEJuoCwY1871yEmmfdZ
EvwEqK1wuNxnv0hrE3vjFs/CF1rMtZfP16QxnUoo2jm3QqITy6hDZPVee0lNzQTK
FpMvfoP24AuYNoWOYOD571opu3tXSHItBxU06lTythCLRUD2ZqiMuj+cWjmEmLNz
CYaw22AGhQdFoDVlWMQoC+jzmRGH6joA0hOQ+WqdH/G+9bDl0BuMSbJJpsxl3CJF
d5uhJ2vem1kex5raJjfBp5oCUsaek3L99TNWadBWstGWDzL1BhN9QrkH375WBcAQ
bUomq3m68ykoofEz6FAPNVDS6Z9a47TKtDKnQ50wbZkxmcABaRkyTKQ31k6n9344
5zqaed+Dj3FpfMhooXx64Tq4RTKznDRrDhefy2wsMTtEzqYWuG88G8ojWPD1yTyW
MUajf+hYLjjqdIvKsR6fgdmD7FPWu/3db4hkEIvPYZUXIdbHVnyE0tbP0moOd9fU
8lVjWppiuC7kmShPZ7gkNLxXdixej8MbgGEU+pnnm9lThcmqqq+8DQXkJa0FROHH
I7sPupYH10yd11m7UuyZreiC0c1E38FzJ2J3uxLFNHiDr7KI3Lf5Ma+6A/wWH/zn
Z9xwM5UeouyshG4GxsOniycJVZP2MiH0izw8tH6Qa6jAM7hFU0l8Qsz6qey6mMW/
GWMhaVQeNCUTWn8jOrBAAy9VKdl3VXnJq1/xwJEoEApPuPGTSMLXIS8FXICeUeQY
7YAgYvpno9hHGVZTUsmwyuRO08S/o3OJhV1ZK687+06N5fU1YYu0kxvDGZXQ9Miw
iqdeLVFwimg+vz7FeG0kzC9oJTz8G7u9MGDcxJQyXeE/uXeMUHRQA8bqMeuFxmdd
NQMDv2rQSUVcU1U55KpYiRtDzZvVy7Zi/ldh1aqfCPj4Lx5aBIC6MAXKXXwDTer4
30l3flgh1hV2T5w+QGJxrPUO9iMQSF//2VW6bHTnLTN8ZoE+cNnkPabRdjLFRqPU
VXWzRPDgTGSG/7Iq+MhkVa+n2D7LxgF7Ck2KNjKViMrt+1QJ92gvKNasy2NuzHQY
/YyFAWpk2ymrnms6xoIjol6ftKm+oIRaOMX94vYu3xNyh9XylhiVvFsr+RtUKgy8
iNDgxubAJevZwzcOoTqBX/DmHSw5uqaWBNA/mNw3wWH8tN0Dv01aaZY+F0wzZDCD
8Mf1p7H9meJXIAzkf07LF/92Mirz+SaAOpef7RmxAFQjHROqQBJV6XwmMesUGMS6
Ga/czDYaBgqc5jSoFDPQvvc1XulXM3zgI+25ywOjbX7JwQ2KZ+5PYl/df8ZT9gz1
QTAV89P2r8SN4omB5/6MSuPJTJniV8owcfJ/LNQDAm2sOqs6YBx/tNjj69/dp9rA
ei9U7roeYvJS6XmkpwdQUq18aNNLKW+5mzQLV6cD4JrGomtckmgt7JVfrXpFFANT
9eJKHGhuDyiZ5tlgtoz8qavTgPrQhMKAbhz+SH3gU2Y=
`protect END_PROTECTED
