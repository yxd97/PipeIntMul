`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GotGBaNnFv0h5BvqRxOlTvTzci0rj9sqNT0SE2Mh5eufSE3LYRsrzqj1Z2M3Qikn
w5f4NX4r3KFcLoAlocDlO9+ZJYmZrOZlN/5q15kVit2mAE7TlhxFTbApcSW3SBP1
BJV4N9KwylN/tnP3eQ9WGBvZk8U7/WZzbA/VOEV5k/B+648NpggSL2zI1aQZW0Kp
6KRFFnhJ5pWx+330jdq2lTcvBrzyhlF8BK+fxH8qxHT1rhWDbgqdNe0nduZSs8mp
eaCUgAO1/cmQ9Pe6qdu4FA==
`protect END_PROTECTED
