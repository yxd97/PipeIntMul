`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+E7ezbO2f7uHHIzPPRBdmLgBcTrzVsQFyCyxteFAIzamR1VjFxquavQpmqGQLnLp
SfbApivfkrc3IwnFBNttcJyhm2xoOMxIk7Ezip6VRM5+3cmI9eb3fB7TJwklKsa3
VHJKzJVJJm8yod6ZXIOCwidxOYVm4P5L3OSb6iDBylGoVapk3ilnS7E3jMn0ULRz
j27jsUqzjSvoRQNVDLgAORo50PlCtvqTVGdM/WvfkR9kX9XmiAeXjri2LMmahaIq
4ptzlGrFUIwNNPPlCVbigdFHZWSvVt8hvcCIwX0oOXN8VsmfB6u7F3eNbbnbKBxE
q1QwZRfe9vUgnaoVOD27UMEm/Q/PwNaRTUb/eI+MbvOKEQQC+BpLDRd5g4A0dhCl
AVannFMYqVEpzQequKkaA4GwIhhdlKg51K1mqlWzL4nN6iiwPaVkKYSgVuvS5fk/
fv2kWX46NG9+TdOrT20VLHqkEcpaERfZaQwYFy4dPJ99KM4mglKQvnfkZ+H87IVJ
U1FHToicQho8id0ovg8DyTqLQVd/rAnaD0GVlwKTMp93SLBDoWvuuiLMS1V3sTNc
tJDojGMmg23ZIERT9nKONL7PWMaBAZIS5s0akrdGMPdgejaKwtKpR6vGeliJamG/
j0ZKdKckKTmHEJzpoQQK1QH+iht9doOqAZ4dVTZ+ZTgC2gHzlRcBf+kNvwQBXiIm
BiTj8dtaVxFFJxc9QDOeWfbJciDa7ChXZcWSQZFD0cFtwzZVl6E2ZqoBqBqk8QYF
aoxPPiVW0ZFlOfe5EGmi/N0iUKgdRKm/zGjAn+43evEGSs8P2qJII1K2dN//Ap8X
Q0o5zdI3TTFQ4ETc8+baqx5pdu77FYpqBZKrpGxAVHiN717Dvnmvl9MtoyEsumGD
ovWUeQanHoxr3Xdl6QuHf9V0iGc6fSN/9UvP3RFmWzDyOFuDE270g+lc2DE51KH4
SNyQyO612T6KPnRvQFeKPio9nQtWGltUEpijV4R9Ts+vcakf0EfB8IwevrzHOjRm
HMd9xatYm4cCNCmJgE85j95I4urVePm9bib1NQYB8qWctVfbcRX+m2eRTEbWRkO/
3PIlNtJ6ZBO6Kkvv9OFnAIEojDPk7oohHFaEdalyDHNPeiALAcdwjjTJxGNLTZDa
TdB50705urSKd1FvJaQosj9tBeuS61+M8YKU70ro+6sHpk0bGjQ/6N+5dRn+HAbI
ehpuHpyxTY5g5m5d/b6wUyhTdrnEsJJDRwCUqVS01773e7Grb1a3w+6pPLkvSG8l
oJ5L12KVWAC0pd6JO3yMFt0daBXNBlqFLm2CzpK2tJd0ZbTt/LVkMrG09i3g6OIQ
CaGSYmo8HKjyT7I+Q3QIkcK9Vzdhb07LKc9D4aITnT+V5MFbk34+kkp+arFbmxgb
uvRRawnHurBJynLpS2FexPgAE4Jx9B1n5bqFaLRfyuzkthPY57InLcbTrckNojTd
BfG0B0/xWA/jU2KjMj6W4e493E2XUfJbykZPCQZT7oAflhPv+iGPMw5wOBTeARon
ONKbW5XpL4tXK8pcSD4OFm3DVmomGTFeh5xVdwXYBOcW6t0pF+1GND9RCGqtzxqc
yi8C+LxmnL6aDYseMZX3FD3nIBg6j6VBEVvhSDgJmsfDdcCql/WumPMphp7OP8ch
z4JpukyJ+esHM/Jo+/r1h0y4Y0GqPXlEDkhjumuk86937KdloXlu8n9Wp1yC3s1P
ZFe4U2v1XCux4VXgjtjtYy9awLj3QDWEy1VIoLWMdTSYTfnDNq4YH29FaRamGPcz
zAuTgwMacG6UD9b9IDBypgSmFAEQFJVJ2AIHY8jBmf1LwIaBNum3BOYkbJm9Eu1A
rbxNo5xbLO3fL8HH5/WBlhZiPQqKSWqeb/J40i7GuNyqKxypfUWiU9YQg49r/E/q
slDgerX452kyx0KuNSIwsu+L/FtrrIuwTIDCMjYFgZuMleNXyVp1irocTuCmylU+
Qeo9UcBl8fMaMULI1PFtUkcUsnbGV0kFiy9rfzh3ujqELLDop28frwhRhHtwcugj
iYf5BH7HayIFwsqMOjm+bEO6hewDCeA4ES6N/20z07sMzkuN4GE1PlAgOFqvr8Nl
G3y8cIAvkWH95Tq33usDGX1YmQMELWRQKHVdR2MMPcmdytyWrW8OyhHftkXCSkXL
MqIBGKPxE/b5Ck84GDz2BZQ/9lRTFZPuPI6dXB2JLnKZ9Kf/QK95vmw1Y6fsyk1F
UKSAI2FlxlZJJqn/rr0kBLPN+IsrUr74ZopqwW6Gs0JeBV/bRR2BSMCbexVOZiQQ
BKp4PTNWYsHQIaL0RQ3L8Z6gh5wPT/2xD//G5LOoEGGUZrIl29k7spSv/YlQ4zXa
pH50H1jtl/k5pyl231H0LKxJdWFH0F1sUekhOdu2YF5F3V68IolTWRtDc0uu+D5e
mv/fnBjMEdDFvK11oz7m2d5IT7uResfYK9fNPtThST2hgUF3L2+IWrGRn04p6srA
swL9PHlH2B+/zATwZEXTd2PK83QLxhTLqPNet55TSUz8hShRM2ZzC+Qh42irZitV
FAvsFcObq881XPPMgsBiYZIuK0cLwZ8aEYK/uVfbZSOqy9HMbhUV+FIurDFSYGpC
Wrvbw+k6i4uSttiPyYzd2F6eBRWSHi/xS3h3SO5ryu3KRiHgRMFsAlpQNkMPzmXB
jESff4+El8fzYpmHlW4xs1PsSsTz2SC0aZlhALIF3st+7lnsKI1DyPXZVn7YpWko
orPS67SHuf3/RC5TerdvcmygQZtfF3rR3G79SF5nZoqK9jLKUsY602CKZ0214O7r
1EuAtczzD8iGi6+9EQzDU2PGArVK6oQGLj/4zAk6T+sonQojfjJadbWr4DgO8B1v
Dhl71zHt1jzBIKLS6mY633pXz3SJcYrcXUGPOUU6uduMJZ4kFY5aa2KjsOgcDm5d
MVtVUriCdPLLwYKpVikXxv/LSgs3JEv2Xv10NLKJ29nRxOV6McoIx48bdAsflnPg
M9NzWJuOhBZZ+EDTv0SB8OIHk3Wuav28zGMpX9IQjrPymAwZbApK5laU92E0Rcv1
tZXk8272LEDZLEroM+I+hyM6LdHcHgq5VhCVUrn2CnbbU6LXKssi60ioqbb2pWmN
5v50XIo6r2CaoFMQ5TnuCthTumTMMn3Sf7Xer6AyDm/NnSZia50jwzwDu9RfbyUQ
lq+93Q8Z7XxYRlK/8gDrlsHzaewmeFmw1pwJiLb2JSMqVADq0cFyLCRU3rVnXnx7
ZvfsftbW/oyz735p3AJ/iVqJwb1jbfVMad+bZd2Ot8XRoftI1fYQGW57kMkJ9Tse
miGbK/UJzpeVwDRiYiQPqZL9AvaM0xWODlE5tY05NYl7mbOo1/8JjFd0+4S3k5sg
zvsrhdN7xKx5COxOneeK8CLBLl3kIWt8UGhOSjQ51eGYrRl5KJBmGnNoDnaqRyVs
76VrcNdbcqZDwcPQvEiQSNmlamUgf6YKXL4u2Kowk16BOveLVK1EhFoOPmSoXE7O
CSmGuySYpoERgL+Kcvs0+/B/8o0cFG0WUYry2R/Plp1KAw8nQiKFIEcAr59mtGQT
2veiHlN8JQIjW0YX0krYc9nlgGkj3ssbAUje/RmJ2KjQ2rCd/mJ6aqA1SBnTiJfZ
WYgUSW4rwbTpYXd1/TwI7I+2gqxqOE0ZmIzT+GRKSEWXU2o9+ttipQy/RB6WveZv
gbuAHbQ1yWCTpfW1QBLW2dZkLbwaY6YUkW48XmkwYXwSRyPkplAnELHqA/zSkspL
1kunfPlGiJaDrIM9BNs0sq4ZWekOzAUxQ24ZknZeD80sO5IClw1xDFbh8NukUcsS
Q9H0oXc5k/9qi3ESk1KEwv2cduz8QXVtoLplijaBnEKdc0pjRh+qGIuY7oVWhZ86
83IXZprPGw3xArl05MkFFJPNVPp/1MPB8Eho9vWCOEqZvnuge86a/pEX2n3Th6U2
B0tu2s12NcGUVgzahfjyl1KzjMg5550n1xqBODbNWSKlcd35LFqJR5hxiyS5wU3V
zI/bjwAxGAKfDqe0+n660K5MkUyZ0U+bSTh978IQQIqD2x/ZYYmdp3GSZzjGHfJu
R1PzQRM9qRrDHC8WipvMqqGLOKLJRAqTuUxGiMOxM1X108JwUA7sE1UHJwF9hPZj
d85O0RUwc1I43MeKA9v1rcuR9TG0FFP0A5D9HyYNyCqHVI/+0bACx0ZLY4ZsJbUb
AuUYl6psH8AqGu/n1UdFWpDAB/YWvxNP9BtViSFKZRqPOifC09A/skC6gr5xmIR7
2m285CVg2c1oYbM9KBXnBg==
`protect END_PROTECTED
