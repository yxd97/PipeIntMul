`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IdVk0QX1Y10J3YtjHKNnClZYQAeqdWvzzz1g2ZUquehhUe9aqWtRlj7GWvrZp7BO
m0pZABoRAvnSrXhjKgWIOgg7qvStNpti+JcKrHB5iLWONVjdzWYgrJnsDSyyoclJ
MfmPRhpwV7wBV+BEtW/s5/Ajr7f9PRAk7Q7biOeUXxwT8O7g+dEcAXpRak8oD72+
aQEv9mMul2xQaYs72JzNYkHzFi0TTy1geGF8HiXd7UOMIGEwJW7wZSRFkqt04cVR
8rcfbs3yd8wn5LMmQyBc2UlmtHzrlnE44pMmOMAW6pVy4ifokgY7MAYx5Taby+TI
vjpFtJxdfY/9C6+1Qt4l8A==
`protect END_PROTECTED
