`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2h+Gq8BRlMhAVaoWC0hpu8MgClvowAMpwf8wyXRwK3hSdxYDLylx/zMWEgMrBKor
ND6yKxH+GrnYPUrtCNFkAkVkTjhB7H+EPtwSJf+U9lSPCXxZCL/wh8pOx1x6xkoh
4PC6ifT/7HbSqzbQr/cQ5Y80FII7NBhelQWkhH5mhwyYDmLJGSxF80Wft+7loAI3
dN13XTpBb6AmTUkYWncchH4yiGxUnY4EVHWyL/5APgwjpkbCovEJqDFWYK9c+FfA
Akqx4mfDvnW8pj0x1qJS5+HMI22T+uJJQ/vOx4DREcYxnx4h92v1lHnG/jF0yxzv
vyASMbz7PiwsNTG1SBjoAR3PhA6jJkdM+r0Fo4zUefT9gCtmAANv6QeAtOlC84vI
dQapVlMXJv3UMLym33AKHbgI3lWzC52wAeNxlLQJFs4muwcdxdjtZTu4+7ZcNVXB
C/5w6FktqTbsd/fVWAQsuZMfsNy6+IjQu/6PgxCCkOD66Xb9zVAt/42GYtjuKBRp
B2DSLEtDOTSLNIyYc22QRpV6tgakQaLG3FfgFJ43NqVf7ApzUhH1azwFb+e7c5Hb
ajVxS8As0rJUT4MYSSKVKI/6wWRAJ7cJvRsNuEax6kbWrI0u9k8D1HGBR1YRMBwZ
ohKppuL26+x0HWqDn3OM+g==
`protect END_PROTECTED
