`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I59KCFdPANep4TPZRzAEj/j5+nhxMxIHfqpK+BSX1dhJq2/BAogaxOruip/GiZqB
kwiPC4yj3YYLoMiampnqVxmNlkQLqcuY2Sid0RAxBkKExA7OAdteXJl5e7WjvnP2
ddCgqjzP1xw6Xnk1iYXwKiMe1hdWnV4YKqrcJGof4oN2mOcle0j5YesDahKHOiPZ
Xwk2nIEcXWDuypBCB6Q73LjR2Run6CtaPAJPg9BJ13Ru67xyglKI2E5G/GSpjxGX
5Qoo+CfILszDJ6Y0cH0xCOI9O3o0m7almTZ3WRg5tP0NZQK4/jKzIGDo9+7s4LQP
ZTQq9fmsJk6fpCs+sgBePhMizCk5an07Gcb7GxVDV/N4WhwtUVfeje73GOPy0KgA
Mc3F+N1vLpjeWvM4rSCn69+RMaa72NRMP/hshvjTvKXY5TJA+UaJGKhtVvDszTmC
hJdrjaPQQGblB+eYK93YFwBfeFz06NNMzBXZBwmVB9Ja6JsSb35Qxi1OX519HnK2
djLmmSOqC/pZNkZefxtZJw==
`protect END_PROTECTED
