`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RiVSpfxejsNywhFUwm7s42bmCtTB5Z9cPnht2oG7QiYj9nAzXjsCRwUvL4kfiKgZ
11kOdHxTx7QxCcz8ojvIcz6RYucit4mrDZL4Kq+L47fo9cgWOYgXDeKZOsiC2C9R
DM2pyKTNEKsZ6eeZPVfyy1bFcnP7XQ+Q1BOhPIHr+xHj1a/16/3oDrfkaTmN+RJ8
cSTSc1d7+8XXjjG47Y2q1jyCtael8cpBoJaQk4srR7Xv5dPJtrKQlNRFHUk0ostx
ZqX2VxewDDYJchEGJCCNYDfKDraTF0YiY+qoYeos9TI=
`protect END_PROTECTED
