`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ChrGEg2js8ZOb3fsMOXZ/uZ34UEKJXs6lEVE+HUBRsuV7fCquxl1WK65tarNL1g
KfeACf8GxJgSOxc2VYm0Mg+3aIETQmZbjz4fh/j/o80kptQ7l0pIBSETC5/4qtKE
LV2cPFt5dUDsPMQR8NRGXRX1NXGrCbRZlvkL11IWXSE8ueVeoLHQ5Z3M5ZOScYv7
pwmgwP1X64Ld5HZq4EAk0ACJEJ+/CGBGe4J9e4fCmgRSXJtv618xQslL9Tn0Dt24
6J0iMDG1DPQtqIK2GHjoxIH1eEgRxtC1LJJ3CHf8ozvP0BZB7m4rWXaGgtLujK+U
XBaotCRUYLYkdQTdq6aNe8zSteufMtOCrA0vgnrRMRj2qK+sW3qt/KB4Cx8T4xpb
aaf6vGFqPNJjrHhnag5slw==
`protect END_PROTECTED
