`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QKQBxnv3VAiXvuftfNLTajmdzQ0IZgCARdoJKfafbpbXL+YK4UBagY1LLsun/HpH
FG/4PXyQ1s3T1KbAiefWQ4xLbQmeRwZLlB+fIJXuVXQOY/k3LN9VhPvwL6yAd5Zy
Fc3b5fSYHFKcTdqINgVuekO5BVe4IUOZbjN19GgdkexIMdsFFLH6G6g7CGKO3TUX
CVW4v30siqyMwT+VKyHaVSE9QTOqxLkPJ0p0t7JBDRXD/ofxBXpphd5bBe5VXAAL
eiKkIbSvNnuxgGyo9b0VvCU6UaPsUTMxCS24oVx3rgcNMQMUvx6rYC9Gy6nQ68gm
3BWNM8pyGov1TJyn+XO10EMRBi/gekgML80dYPJWE6fdbz4ZEL/FtHFpmgX4IIOD
OqmEOZFkb9pY3v2Z3/ZyXY8P5y3Zg8fUxl6e1krdSEQeafs9DNXVmzKfeInNYpda
1q1JG1c+gdpyGvRKakQrhPjKXT10j6sPLTTT01VXzcqyAeV0y2EpsIJ6RmCVhx3c
yPkB0sxHvp9+BJ4Pv2FJmgnNlLOf4vWxnMthhVv7MryqJyiVnp0Xan3stSuq9ssA
VTuiL3uWZFKxJ2XrjO0BUEVZ5bD42vjuNs0TVUqJSodPhOCJ5vCf52f3REMTlOFK
UutqaceGSbjl25WJkLv+DT0GQBAZrd4P/hpeg9DSl4r8NFos/QlSZLR2DExCF/6z
pPx6h5O9J6ZsTIu2EMkwYd6Uk+h34z0LQEWrw5eDfkdMPIy2s3YK1w6ZdwHFxcT1
L3oSJ7mm+3nGWmWJyEgfcchHqISY4ss6Pqn4cW4nHsz0UczPhD48rGQHDszRvrK6
xPav5+mGgcPey+djQPIyrqnJNaA9Va7ofL1S8D8a4BUemw5z5TjNV6UWQpTfFRdJ
u95LjJn7KK9UDaIQN4dJmuay+KXgBUb+Fn0pfpzXQr+NDCUKk/8lYt4olaZxzEBY
hWM3yRy0Pyqe+wSFFepACuCPxyYwDFIDNfnV52PH2vz99YLrRB/4bZq57v25cHii
R5/PBXbzs11XszCxTqgeN/Abxx7nJiWCXLzK7vchnfu4b7PM/UsEhjRCD5nlCwx+
0UnwjIaM1l8FKHhjpwZepci738b+2Dq9TAoXSd6Uxs3xj2yxo7+sW1YWyONBJ6Eb
tN89369CvOB6eVC6d12UU9a0rLrLoh6jlL23gK+usnhux1gE1wUy4DIcXli/vMSN
XNlYl78mYlS0tBELsgrpfZmfYo85wWKluZ4kOjIgoL2HL8511gsZoN5SFvkPMKsL
BYHbxBNVoskGbtYxqs++U7msI5MGW4XoV4J/ktFFxWzcgSR72uKXwojGTbFb2zBr
VWA92Pbnu4DKM7BSs2DUE7RS9Al7pwKlKZ2+FZfcqKVGLVVVsiIAEdqx+8q3Ki39
xS1trUdX8Jw3XJqaab1C6XzKhJtsb8JEtGGd12v/nQfSIyveMyahUetabrDs2SQo
zqfKV5BlatxiFfNYOeaCVBtUhtjkcUfHLEkEoJeRuIpObw7kxknbhP/5UH5PXGZz
EKfqD2cClY7tuyDh+n8Wuxhg9h45uhyw3O+8zjRIkXXbAOp+imyoqw0haXYz/OnK
REEX7KUxmhnCBveA9XR4YFsaCEKa6HvqRtPnh19TJIyQrI8zEOap52+rj4pNKHhF
JgH5WrQJD7z9a1UpcloqDY4a5tfvO3+ynXyfSpuYxYEXnSwQ7HMLwMH76DQ36n47
GHJyKv8/o6UOue+dsA6ncCCvxE9EqdzJiy0I6wnCaoyXBDwlR03/Y0jzkIbo9p2B
YX7//14yDYn2xrkivox0Kbh8CK39eSIfuYS6lhnwGbt/4sumU2Tu2WTKhXgngTUU
GVC0NPgv2yU5u76VTRY81fsm2YQYbm63C5zynzxdDeNZpWbvPsgwEiHofMGERCb8
ov9WxLVxyOivdl941y+E8mUPUV+4oCww/BjVY1inln7kjuC8ibpmX44gW4msBOOW
oHvfAG/dHynYcq/5ZylG4/soCMyGvhS9YZnkFrgNY7rpdM96wgBg9DTbVoCCH+Uv
/uCpLOSNA8qBtCGi5UyDlQ==
`protect END_PROTECTED
