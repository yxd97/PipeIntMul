`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZtUr30hle/LsQwaEBaNnHkSPY2lTOcoyrrXn1nxoHjcCYVLSojlLNWmulukoXbDb
1t3FjRPzv3/Y4o59OMMru7i4c0VjNBwCrtgemqLN3CkG8fuHM2kq3E8eYcK5k5Ul
Y5/NJDw1rovT7cIWUOoaIESh3SOLiWtyzdwaAofXebdiMUk6ztbr0kG5XPXax/yt
1AGiUy06p3l+ZcSgiPfDwFLHllMu2zIN09f9C8I5NLEKOKCH45BcG0AdbnPJmMSD
NZwdFO0X/GGhRoqd7sX08wp8UQiYTECPJsbOo1cthbcOlqq3FfZoII1wziMuORAq
RqXlYIeu33e0lYDn1M2/TQWSrnjw7TCg4rYAW0ZZA/DBC97R/A39LsBxZNgqZ6Tc
EkOa5UQpEwJNyMziPD30K22EODaNmanmaxBdLrFKjKZdfbop5HE3/Ho9T6p2IoJ2
`protect END_PROTECTED
