`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
snui+h4XmIhMJ+/ze/bkoFdSrGVGkGUphqk0YrPfPW08cTrL2mXkKpUDGKQrns5t
u6mZX+U6JCWY4/SxsG/RVQYz/G8WtN2W0pAJRDR3E5fGbHh3QUGHudnjmpqATyxI
iB7dV/585uFJwzBGQJ8B4MoMYQL1JU3If2ivbVqgmUtgjne2qQ7JdJ0uoEskcCVc
P1076rhNu8hK7nXlrPwFuiwT+J9XVCEaCsGRBH4Da+B5YrMMxyb6SKXxxTiw+8J8
c4u50bkG6H9w93elcxXVmz7SUqRDqw5ldGKzzaYQ9Vb1jzNECt6nEog1fGGHde8P
`protect END_PROTECTED
