`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k8zsEJE8uNZeTgLIdzWK4sYXSldQxAHDcj9A+3vD4drbTqsbZ3mhO5WscJwQbUBN
rwwh9nhOU046UqUYHFP68+XgvKF5QSexM6Nj/lK2xTcodWHP/RxCGGZlFzUHC8zu
f89h2RIez7kkUVZyog2oZcitBaTKW7d0MyL9+AScbG8f1/EFfEPZy+fsOYZcyhg6
zkmOfB2GBbLMcGpxD6zRZ64P1bMJ3RlohoMsxcx5Ww+eOma3lSqMkJ7BQr1/5Z1+
orHkpvHGZPUL6rFJK0ic020fUDh0ZT7Ycjn9E4onemkXrW1FUKK0OgitC+2X4nlI
52ZV6EkcRqXEjsW3BoMMUtHZ21GO/FR7BnmSHA0gjy2I/PDXBBJCSK8q/mifJJXl
bErvLEp+8iBe6fQK6b7sV53KxEJoj5v9/GH+KEuPlv8=
`protect END_PROTECTED
