`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+elDpIVz2mQ0y+dhspd9yDuubbBm+BWF6d4Q/G79epwxo70qA6sV1GneMW+fYN6t
ECAEJLlQ6wyddyn7pncXPXIPsH/YKvznhx593e7BtcncQLoT+/qxy9DndjqsceVi
oeA045+/CR9+CMqlyoDcNUM2mZ6hB20q4WOTxx49SBjnwUJZI7bra/p4TKEC1rfQ
umgwJAkPiTI6j0kYIsV1VV0npIrgSkReBt8fSdMD09DOjdjIUjSSwGiX5RkWtUe3
alUZ4DKuvE3sXcvJs83dGRfDn3nCw3ti2SpOeVhrAi8Wo5hCflCCoPn1m7EHJqOv
sONPc4YvLNhRpMOu7LBEftzUK/prkTIEsRaeGD91XmUqX0T/SznGlsYLN67csRIw
1+dFwBnasf9e9itohu5hHhWuii/FJXH2TcGt6B2LXrss1CYEyJoW1kg0i0GmYPB8
7oYLLzvXFXsV/oxhr5wNdFqwatvEEFlN4T8scEbWRuf/X4Kkc6+lCCjdp5BCi7Go
ObWtMx7aw+dx63OaTout+C+gM4y6MNCdTI52HMtQWFg/4G9H8YPzIG4JYpKrba5j
dQryXewgLZC2w44c3/DQ3kzVO+P1Keq9aDjsoTwuqVqddVP8MXHtHzSVKQwlmdBz
w/1T1/rED3IXQ3BHPVjmucVMgZpVNdncrhXEt+QGxHSd9HMxiJWqKVoF3qp2YMC2
elnsrbyPdqR2WULw5WFQSELgNlfLw/OdU7HY51b6iTr5pIUxyqNZxiLmx80GRx9Y
MDp8/J00FuyR/g1y9xg65QipFxh2dtl2ZTXHx9iNWUPaQUlNg6DK5yD19/si5xHC
ye+RpZURP6Dm9l6ITXF9lrD4auP6dyC59elpYtrbTtmoP2a5gLWvnddfhumTKS8D
Vw1MV8YgISGGfR8XDFsjGrNKXI7Gl9smavN5a9Qej7lbS0/CK5JFMSa3I4CywvlV
w8jIc3uWhKGN8tPP8+YBq5hTjIT21NPcl/r0kZKerek1suXqqDd6Xx0J1hBSc8hv
81kJHoVKV2X4cFt7vdQUsq3Cwp6sap8yZrmgidNPEVHjtrZIf6tan8GhW5qDbDTp
SGsScht43PUnbinSsVQaUi95SOdVs3w/HqHLCq6feTetQZqLyOT8xgueBYpkY3dc
M+d3E9fdkurxGHqf2/Ood2y8cF8YInt4GPIAggoUDENWpOecAed7w1jbArBNCDWp
AsmDe+94PEv2d4w6X/ZAcngivnqdLKWkIh/7/8Ef7UdgzoTtOn6H+U3h0Lv+Urv7
1m3iXSWEmK0/8oPq1NIQC8GGUhutmRdl65qdsiosH5QIoIDdjyMTlL55A4CLCqkq
61L4z+I8ZaPJkwWCxxBRBL94vNWlVoPtR6AINy+Wc3P1T+qF+4Qo8JGRWrwTcnfs
P2YgpYrJUPPgXy6ENldoL0aksHOcBuXvkWlUvwo8uCjwbRSOCSuEKTPEEC3w+cvd
dW7oGAWzTdWVZgTPZ9UXVKnaSTr4abBn1Vejho0bEBe8JuVVQcBeQCNPx+B93Nm/
R/RYv6OVitJdwf7P1RoluHFYbZIyxCHe/LihqC0oMSY3AalVlfBOS70ICuzqaERn
dRD53wSvexYG56AIugb0ERtiZc6b7v2yzfG67ou1CqsI1GYYOUoURXHw5OM8r2oh
Szn5zykpqEu4ZvCOqlNuZOrJtoV0XeQ0sFWPuuw9zuzw6z4pXcKLKg9YAWPp9HcF
Dmhv4Kn4Ki1N3OQLWe3j4KAxr8TL0U1C8bOqszJfHlAdKNddRjeQwIc3QXipakGi
YbMzLdCgfXt927qqjMt54OeSvPZr+4vzZHmDG8dHJRFwyvpv1OUmoadp5cGRCBYZ
k0XjJ1ns8PrgBkPBbyslG+toTe/cRK9S5MCwH3JLzx0=
`protect END_PROTECTED
