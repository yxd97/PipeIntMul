`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RUzwV7warpfzVw105SSVh5UwCDmN8MHGbrgE0wYBCE+TxfpXvKMvT7SeC1HC6vIs
msL+jteJ1bhkhD7Kwa7e2Iv1r3Xsvv3TZPrq//IhMJfdFrI5jf7w+ENXj8g4H+St
Egu2MOdrj0pxsk06Ia85pRZiaPG+oI4dFMFnWNOLATYunTDiZkc/VzepGh/YYyZs
ILZJgPwyB1l9KSknm7fpswq4meOwmirK1EFqozKAe/eUNxFe0myMiUQrAJvI5rE1
pQi35SL/D+NY2iT3gDV+ElxcEnFmCvnWFhP6075alDPpeeYofJqeY2b3ijSszilm
GBC+jTWG/FsoFnR9sHFRAwiDfLTyyLYSH5xnEqWCcPyZEhcwjmKU39qZj50n/F6I
Zc69YuetOj/S8XNygNmrtHitk5bDcfzyf5ukzPCRaHor3vOoTNY/+wtShGyMkC9o
FZVvT9L+ER3yX2HvPvVf3sbifxoIk5mFo+3Vh+oxJuVrnWATcbWdnHjL1xoxBPZH
T2f5i3XytMcwk52pyMsf3ChSmLLAge43k4SUfrDVdGpHHH7/u7/YvYT39qyxlcVF
ONMEvigUnUKxA2RPR3NUopl4aVKCj3hRkjVKQ4tBQYrLXWhW2s4qraMgti/b75D6
qCGjz8sOWTWFnwyXaYIbuIDTCTUI+ossD2+q5H+Kes1tHTs0v/gJwBQAKBJW0Yfo
oW0DDBcE7LKmXrh6qJr8Cg==
`protect END_PROTECTED
