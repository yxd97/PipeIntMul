`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFfF6GzCMtIi14dln8vLtkl+4JROeaHgiAEisjMkmyDLG07e4WQUJYavyjnaf7PH
/kJR7L65bqJeC/YuOTy5kU4Y9LLsgVK74jPniOqu2zQ6vubYATTUGih0+ND+Y4cz
6/og+to97onIeCb5Rf/uCksXMT1LDT1LKdRarTx+v5zlMv/8WIO/oKzhuZaUPbeJ
VS2v6r+PpKHa+h4RdMPgx4H2JNv+dkNh1ymcHDs7E0JKwsGxU26uMyuiciaB8wzt
PGoGj5NjIO3MWpCUFgFTb+pZyR1JEUs4ITxHo9dy50aJPySSl1RolChznRCxUYm6
ZnSKIPamtB3RRlHnQlYbuXOZSWqtTltckZt/l0+WAt6lgIM3mCUdwtvjrKPvNBX6
KI+dbsfA3jLyLftJZnyNiT7r/7kLOylTLwvaFp28FMZ7l/+lKKiWXED3JfqZaA3J
A2F8ezplnd16p+Xew9aZhg==
`protect END_PROTECTED
