`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7jkTt8ZztdrvVwm9cPQ4Th30/W39I/IFIf2zNa/cHKoHIeG6cRsKaCQOwW+pUvB
t9yCLnG3OzWF2jWbajbcfK8YOZ7hKFmT7opQIfS1LDa2+WgRxJa7ZDYWCIP+ACb6
Wf4nTz0zwPnwTmQ0s3E8JlQBkbDUQjWYXBzweYF6xCnoxFh/xrSgJq7QAmdNVQ5H
l0afk37aCaFW8L47qHiKaVYSbH4iT+2/EqPVhfMWpg1HsQ+Pt4lHFB5fJk+8kdf9
NGSUhCDHWDJfxWb9Q8oPUPPun6Y9TYROFWp0k08F3aDDIfIwQjeHlOgNbjb2wE2n
H6drIkpo1OGPCxW4Si9mmNoFJF3J6CVA1il86uBxuaYE+NdDQaiycoZ8xGFY2uvM
K0P0UKqY0b9ntReh8X8hs4qPOEbj6CMcl1kvtN+qISWHUqiyIyMqtKw/d8Csj3ax
p4zQKLOXMXtk9MGLS5pn9TeY1oghckS87QLx5ZWmDBQ=
`protect END_PROTECTED
