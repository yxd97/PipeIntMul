`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YoZGz5W4rG7L/3nes/ulPP0118SwjfSUqeOpOGen2iMmZpswmiDS3gwNxsnOfKR5
au4JmXU7wImLO7XsPnq2g3jf3RGweQAHCSymJoWB2VowB4n4JKN3vNC7gtwvCaQy
Qh7tX+1+0nblYjU0qPaMYVaEpDG4dogOQ2xZV/xQo/PHyi/+i+NxpzDUHDe/0lH8
/ve3O3Tq0+3SaxdSAzCAvNRuinU3ZoJJ1BSBqciYbVZSrFL72MIR4b9jTFg7ulJV
+zDqc3uJdwRvMRloVDhjXQC7JtppRz/uw3Fmbjjk88OjUL9yaFGfz8XOmmljqSJ1
O18Oa0UWVobZBgVgXgeMDa2RNAloMDKx0ibRjKRNQ2RV8BEhZdro8+jf0c82LWID
biczPjfCAUj7uVaprtF6HwaBmNsgtx05EmRXxJPgm7f+Ko9bMxD+Fiia1V41BzVt
8Ypbgd7sKcuBCc+53DyWUD7elqQFcpdU11fSkr6Tet31Gtb6GKpdVrC6lqR7BT9d
N4yBpBgA1u4fvGQyH9YQxKoUpd81qj3G8pMB7Zt7hX5zdlDlIMOFQoeQqmpckrzO
nxASq9bcrmKZ99G5Bx8DEjsrrpyshYB6H6FBs9C2WVUPK2fxfB2a2fICqujhW2VP
uwgn1emCNasbORVKX51bg6ELJkpa7T5ztcT1KZm8Dsv26+qRsw5wcM9RvGGWhYGW
IF27b05cnQI8t7YXnQqbY9zffTwWCi77tfnT4xuNoyyj8tpo8OkZ8YFlP/Y1yn/g
Pf3ZJ95HfdGFzY9wWWn4eF4WRXLPNTHb6VWpjEz/tH1wUubwD7im4DIibfZ/8W/W
DPl3PhZubEhPLEF6Fuj2IYvQ+qdDJKHWnS9vVSfx6mZNbips2HAb30iKL7kFVVoq
qvndHBhJCRBaHCb02tR41+zWVChCCaurxnlItwbYBhhRKRCD3eo2lGSkgCYj+mbB
CPBYk+GfyhnCUuEVb5tlroK0TMpx6IqrIzbyKnQWmVVt8VWiAbehhkeOCNrnaXNO
pJcIKaqYebz2qS2XtRsat/piz8ggeL01cqxYnqWc/1jx+Uh6tdGrRo4ZjnBJASh6
JoZf5mmD8h2mPRnLfgOtglYTdvdBDYGG9+RunrckSLoxU5Z8yRNOkCTk5BS0/u60
SjUv1d5nkrBIT3y5XAonyJix6Y2eOQd58SHQr2Rjt8FDSaykVmwo/r5yG//RfFCc
LWlc+Eopk+uuP6Em5MVhMWTYOq7jBqGIDgRkmN9YHq2NR/KWRyBVxKkx8TNJ5eIN
uA/OXVCc2KZizbWb2XZ2/Q==
`protect END_PROTECTED
