`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSXdwLmB/P+yidvP9K5Ni+4dqS+BYHtrZ8gls66vjMEq/TKPEQDdk8ckV7pCjV/x
bSGf2CRCY1NajoqXJoGjgHfNDqTVr9HtMnWu92zUCq5jjQUH/KtL5tVEAM4PP5x6
XzY+DcvQJk62TVxwxORc7KX2zmk2z5+dmDZyWh0itsQxgAuuH3d+VZWr/+sU09r7
L/ojrDzoS9tyEfbnAE/rc0Nzs2oDxW6L+VF3N7NJ4ukbzDPsJWqXvFMBfGOmBfxQ
AXUwE9KgBuSEwm3L4pVjHY0lCJHvMQa6YxmnJDIfHZC4PYUPlRKXBc0pS1MjqaRA
AZ9Tw3nMO8F9W9uA4zy3bR+ZcE6GAci6lxRlr43v5aEZs1ArQn4yWa69rQgvHXsj
g7WRkziqVSk1Muta4Yep8i+b2lM4Givpa4z0FWgGbmh93+aVhRZAUFC1OyBeg3hH
L5LqNZW157aPrZMiVDPwxxHXOtePJswMRsINfmXSvaf/ey3uqirk6P0RBI1uXwKR
3cjmLXuMXJf0qcuhmOfd8HdtpWcqVd3+TCFlJ0JjeiLgx0OE3en2HU1qfDRp8zci
9NhNLDVJo66uEPVUyWQA3okxGe3ww/t9l8NymtS1dE7oEbPvFHm0kBiPfjGNEzB2
8TOq7SE5k3fvQ3QBBo2KwCQVmxMRXGQ+Th+b2uYbhZcGmxq2EJx6kWaKgd6DO64W
BwlaiIzbvPgIrL5n22Qa9S6Lks3jKpER2s81yiLKHFVAzQWF7fia8E7OCzdIqcmD
PQA/JIVovK/XiFi4hs00vRAYzfXk/mRD6ZJifPh3QzAQakTHOEpUsh9ZZmlzrzt0
UDwOhBqwJcPZ3nk7a0aHPXKNY+M7pdkg9RsBY6FhEUbodmgv99Cbyl7pypx4r8Ca
CQJsVLkjfIqtyk8i9BaD0F0ZhxL1XOugYhl1iUsd+7dgdWqtL5S+h8ferSXqnB8H
dglFwTG/opoeKmi7prN97DovJI7yJXU2ABMWWlXBoySfs/H1LQ6JcqEYBxGn/VFU
Z53VPfemmGj/6R8/MifWgeDrSWP8dzPMu081GUW/HlJsPsRlia/dzQ/rTCFtEiqC
KGmAgZEdtJeouOluDWsqQJt0eYL0/ywjKP7xc6M9SSXSH1+eOamc2cHjCufAmiRY
jOx9gIsxUVsGzjLqUfkzR/SBjRNmlyQ5d06aCObTnyuLlE+GGf1a2zHam0wcS+H0
fItiSz9JT2/mMxsU6V9TcFJVDK+9Q9YXA1J2yNNz8MRVf2+8nQZSNsNwns47Cbul
O9b9jH66debHD6z7cOnUF5zbrL6SZIx2MdInJysKPJ0kzXQYH8zbRgvZYrkjBdgt
9DZCuG4RMZFuN3mi+79PSsnl/pPeVdM5/CmjoSj9Vi5zfO8tkd7A73SPPh0zGagr
Dm2dWMqdMwQf+E9WwUPjTw==
`protect END_PROTECTED
