`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eCRmTNu//lkiu3LCUTGJY6ocpqhsb9yPDSNLtt0ziaVpBJFlRXaOtgx+mHrXt89M
+0qPKQsO1Kbb7koffjO2Bicx4dOumDalzfI0m6Vlf29NB+wEGszjG3j5FFDNtOkc
V3Rovut+hFe6NE8EAoXvDQr8cI6roI1v91u/8Jk7zyv9Xtg5lphZUGTzaOcnPJg/
Pkw5D08P/3tfaHfbnrWHPBEqGli0ZSRU7AtgvPTTYgIkiM9QWak3pKNdqTkp80aG
Cg8Kr648yeA49jiNFePu3gmbHzhbizcbk84kJPF7AVZEs1T2epypKuHzTkIettL+
lI1j5Fu60FGOpN2/0Wl4zbNu4v2f87ofuMgUfAL+BUiQFMJ761+z5XYElVASq/hN
3rvuLyGC+e8bjQ/wMcMW2DEKpTGWMxG0eL7n2zg6wP6V+CEoiiE8OOljGUxkHKHH
BBMkbRCIe+Vgs6/CXZl8A8yUrt4qjJB13kG1BxddIRV0Q28cFG6nPOTLz9B9ndKo
yWKEAXe/Y38cx9OLS6fVtUOho8cHH8oGA6/6iq6d7Mr0/IzUxj1x8W5ziimeP4wK
DX407FLjHSPQU+pW+SlKzDXZ5W/dEdLAVVA8hF2Gytk=
`protect END_PROTECTED
