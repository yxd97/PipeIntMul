`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IM98ApTlaWOiUnZ0ezz9GhHQjN+79zdDD/Av7PFO3pFJF2+XkZfb+QOU+pJt3vru
JZsRAxHjZcMZCJWacN2xZD/vAAFKtBn/X6zeAUqWUfF7ofBrFSqrsDqW1P8TtlbI
pAtNDQ4A8ex6vq0Abw6Q7NDK1Ta7wHX+IsfGZQUwZeqLOI3cHuYd51GfB5E59NzV
+m/FhxZeWxUSDpRzYEffb2i7Bs1Yj+1U9Uh1/LXbEpl+kdGVlFfrQZKnm9HTPEYz
/CIzdQjl3pwtxuiVDvpl+q0ZgMlssvL6iE1iqCMOi9BZk9BX01rNJa5dMLZ59BXp
KQiX8JDNJAsEnELhiSZKMmK9/sYqybil4ePtRWMY1vkEv3v2lAGP5pb1H++JUHO6
TDJNSx9XjlQr8fokGEBcDRZgkH7yXDV4mgf2+l5Eb/v82K5SsGo6eJpUbRhnP9UA
8EwL2xTgkFgTpZELy/vprLtS5lC9cOhzhLK2iSHNwoIkW0tNcg9i1WKXWMkuVrIj
WNq28RiW8FbS1vjkEGXNZnYGGIMp1BhXw5uyqQA6TYELQ+ZL4Nze44gCsHAc5Jtm
bXR63pk8mjSIkVH+AWQKPBoBjmhw3kgevlRHOzC9jHL67Kh135D1Je2SZCYkuonq
+Qb/Pl4SzxfoUzbG1x1U+rB6SBfLBy9cZZXkbGkcqYQDxp1HhPBqfCilUhxrko1z
sjxYV4/+w36CzaQWqGzxE3xrtHKOT530reVvkCoD9rPSGW/udwd85MgwAc8x/Xf6
ouqWzpZ3tjzvdWE7Bg+vTgeoQtEPqBTdhCgIi3X5fvs8CV+38UILG4BU/vbf/nJH
f4oI55GraCUtRisRr1Jc2SmE2n1gXTIg/1WfT5uV3HAFM1M2kueFsRT23d/HvhvF
Wir9WnUZ8n2FBxZTqrETd52q5dPTCsD7PR6iNTFMsI2aBVhBYtOdgZCCGNS/o+ys
1zAa6dwTp04PtORWfD5L7A==
`protect END_PROTECTED
