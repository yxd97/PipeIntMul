`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p3tvemkj5mMV/ymXPIs7Agt2QlgdBP2jhJGhIhUTuRbxY/V0G3mas3yQhcpFRhzO
uBdVpOwwzl8z0eeZbaE+8MSoxi2iIEeX/cHzVaqHNBTzDi3MwezBwN72G9Uh1g1j
E7eMzMX2FPMOWd9kFyYJZZ9FaJiBJl1CysDDYmB5Jtobk013SW8mPciBSIhvfggO
R4k685WXFwea/wZLpaTaefC0623GgN/vhcmq4KGI0Fb5Bj3cjEvETsMakiSgLMh8
Wh0yD6zJin95TxCTqVoYQX3mtqBkAlVw1NAtliQI8VK2Z8NvUE0CKFVJwcd/RoeB
0guXVFUR9fbgIYhD3iDjloYGuTLtWeTuHEcypxgFKGRtzJIu4RG3RCq/4+oKImPG
Mc47+ye11ZbP5LRggf4lWbks9J/um+DdqLMRi/o/YvusOTdn7WqKWwocZuuaxL3M
`protect END_PROTECTED
