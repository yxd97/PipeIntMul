`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DVHMaH61NUAuV327eI+C2FxjCop3uhxrFACwegVWE9KzfNcG1rxo2KSXRZwjKgiz
RdzLn0xMAE7xDYFIzoxJuWkkPQpkAhxBXKQ/9J/1YnP7ammUeiShAas7ebBHGMd0
v8X+cDYqr77YCwiEwsrMO0G0sxWy/i4FHyGdyDBFgwgsqb+R3VwlLROotJ8lrv/o
RQvSaSgNyeg0ckLY5z6/Ar726HFanYKrFvhyBLcl4BDAkrX5nmquKTH8IH1tqfI2
tTXLwjAKMC1+1djHFYsa7ozeJgFrdH6u7funzWcgS1x7EEmHRXO7SVlb/PkXG/fV
81VuSTiJH+VQZTZNn8M8Gzhjjk2zOnWmA9B1fUmVOaSVw6xMUG0v+Uo1Yj1jZaWd
F0a5+GdHRV+fwx0XsuixjyO1dkgr8Pyaiq49hKp6reA=
`protect END_PROTECTED
