`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MiCRdgr1jQb44+yC59EwH5RqIRhHRJ8TMmTIg7Ekn8Gbn0cFWudj3o8cGk9VDfpy
YPUWnmmTvviYn6rrX7TvtAVmSfMudGBpwCwV+ECSWqCDf3gVNrPcL235PHtSrqmm
P1C1IsNAXMeiasfX/vekIJ38nGAWCJ35WjrssKRtMWjwrYcIxJW3H6HzE3PnigLI
XTfevAdo7V5R9T4VprU5ma+bKLe4is4R2p6M/mnzqulho7n0mrU/mYYPTj9xrbNl
3rBQOd8qgamNHxS3GbUu2sBvrJC/wAIr7bbjVTIGMmGtGCzMZgUeFIcNHT0Cxzs4
Fqa/yHWd/quFoXq+qGppmyZ5IFj+KAJgHJL0KQSuEeDoIzA9sL5vaoje4WtFaCyb
fDLooGrli43S2tqlTAChS2Zo+LJ+prN41kkyFacURYM=
`protect END_PROTECTED
