`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gYjNdXhysHSJAn7rSvRVxoyK1OXNj5Nni8qEj2FuTf7HrpaxclSa8aOJvcpOIuPu
RLzmMU4R3+JCSHgMakypQF1a+BsoeNui9g0by5MkjbrEGdFl2ur/r+ioyatmwFFj
G0V2Vz3ixpsx+nUeHn7zm9DR93W9kdSdWvPwiP0bbf8mDAQwQ8nHcY6xBqtTb7m9
IMuchNZ+bw3jCRoGMskYvQ3nBSLn2iz5emcMmVm+EZwqeRGZSU7AfNEfugYwhK9w
6DaRVXc0gsf9sjYKtIr4lLp99/+RIDc9RjFLBVrHqKs7tgfVqLB0v5lwbT+m3BqA
FfnVaKR3wZOj5nrTbKywdt6RzwkQbeqHQpRkU8xQyvY3q/FOKoJ0FtoROQFuoF+i
9UC1dBZ4MchoL0OzNgjhvE5OSTLuIl0UxL3wR9a9OdqnwK/WNdUtd5nsWq2gk5Ud
9G1lwiq3h3H+ujWmxYmuboO8I3QSXRnAJL/Z9CqfJVUZEBMS2NvGpffnXuIzmnhx
f9vNg8jITnY6fRokZY4KLVreU9K/MbsbYijJJF3db6fN2VO40dSt3S9Nt1u5DROQ
VH5s58y5Hh+1Bn1DcgDLjlELhE/vwGFXbDXOADxGSR1gmAjWTuAKj4jLlnH0MiZf
6yrezvbhU+uUW3wtc7n1rIqU0wF/BYTU4xTctdKxbF0yQF1tdQSsu6gcKyCCl1en
1+ALlJoA/JjOuDSGV+BKoJlKJItLUywnrTvNvuxma6+74erSS/7rXDhGitNHlcMd
`protect END_PROTECTED
