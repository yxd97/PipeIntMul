`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9Za49FweKgyI7cLkH/c6v+TrI9hbbmQcX0F11I/NjzVeDBx+rNLvs5TBtlqp5pF
ausn5upwWXBwzwpT4PPFl09rN9M+jupqHgHYjAycLs2dx/jU8Ebxnxt5aFfUcFqU
V+Ha9zjor3u6xxXwMvlL89MFyiVGDA82Opuv1npyf91OGdFmCwVA8P4TC9V5u7Wo
rVw5tg01hCfzLK6Qos986c5+TEtUGbxzv5hoa9em/iF2gZ70wIpSiHYjswFRtMva
7GhfH9XXKhopfv399ZNaUBgm4H42nzOXGKYNV/H5rrJ6hL9lI+JuLXzxb1jfpCUc
59qc4IYGRv2dWlDvpI2Uz9+BtynmTEJrYDTgeOSApFJ0E/qzLkEvmpHrQHuad4Wf
WcQVEIJDWBmDgKoPC7ubJvrLCLPXHr9kNrQ0emhlSOgzHCFycxhlLSBibZ2Oh7+Q
xrJ9RFCdKY0th5Phe1TqcGpEWD8hysyqX9EoauNmQKr8ue3y006HZqMwB0SNdAH0
Sf3JMxiCI8l69loacM6/0uphyo4BD9JugBlWDQpPJIzjgdcFfX18Pt2Ts5xvVXm+
nV8I3/tMw9vO4RsjXpi77RcM386Mov8a+fzbvn1yhkWe3eQkx+DWY5G3O8SFgjEg
JLaH6ZtXsAQBbEve/iRljw2UAXHvpihXpIIQv7cArBJysWcoZIxrVdHewTeLtLgT
iyLDISjllhIEcRselBLjl4VePqrEOmTAjWE1TSgl1+JkBkVBcmunyqTewV/7NmSt
6Tle6JYpduK/m4qnbFvQI/kUGvim3wVEESxvsmWFFPnF8nJgkPu8TxrRXFznj8th
1epssgDOmQatkHcYvjTMi9BEi/mu1PKi7p1HY7K37GzHvGuIrbyBtPFcglsUy++6
sa+zU149Im7Wr3N0WmfFGJvgMDfH0VCg73LtJC9Oq9HvLnXRNtLPdQp9TQbDv7u8
oI5ji7KA5HhYw+LoP3XcyQ==
`protect END_PROTECTED
