`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6z4wziQvWQPhdzJhY8l8bgFb6DHUXXQgXIGfIGaOaUPnLDOliWSCvZFQaOaYaUc
Mt+ojjBcqDRgIGHYr6LHnj/zKBE75ghVWe/Yre027hxKJkoRQctWSIh0ZXjYoTvv
ERmi0JVxDfRmZQsXkKyPZ/wXYW9Xa2FSBf1F0ZdmoPJHz6uqOhsltaBoBocZQKL7
kKfrkDCADJfeV0cF5/fD712nhBoHuNYF2Fw0M+9QX+ruj1Wk7aJGpplTRH+3fB9G
E5soXUsUOlLJACJfwRBVEx7JP5oIjs+2E2hQfjgrxcZGT5tOc94WaPKPhqtcPMDC
a9hFPVONJa4dgPpOg4+CCOHH9v+SRI5Nka6y8OY62kgtI9dMVu8bJtvNfAU1h+Aq
44vnkXy5PW1y6UFMBMHfj/KIb/CL6dIIDihcT+xglGGxl15gmtEybvUbO0OaeJpM
b0dCUU5LoPOaSYf0wlXLxasbAkJHXxiv6pZf4TXkZhh01ewdFx2esxgIi60Ghjx4
wfPvWlwNcaLpO7tZiZS0Gve06Bz5QlDEMlSxSrNpbCcb/+0nimYsthkohOxb/ank
DykyiFUl1LFYcZSTzgzs3Ptc2/kBSNJw6l3tQKXF4W4rQ6VfPiKZ5HOIvufGu16x
wHDHvk9oTSO+YBX6/Ta1hPJUzQQ5FVDtKSmcjOGv5+QUVX/U8ITkLDjWYwncmbAC
dY6gFLXFfKqD4GkKRG/PKN2btxEbXLwRm2hIXXtlxGTtw8vhiOWQF1oHWHkY/z51
Q+ELkgupO9Gqszcj1IL5da8z9PTUkjPFVCWKpQ3WIL9humoimQuM/A91xlLoBopa
84yV4UzTHbGemWNu58RjKz4fw7NY1GZvDTjoLZ+sz4j3EbiPIzrE9epO1pGbHzNG
qH2ezb+nPzgCmfFblpAai9kkuOWaEr61uEVsV6oYDj8JDKED2PLmuErZSLci2jbA
6IFuqxrXYoLOvPk+MeAIEh8PH28WmOXtFip07IQOGw4bXFA3SPUDaiqlFcH5DyQk
WiONpVg2cBHotwQCVkNfCvncFo7OK3mYqGRVWep66CCLdPsQ/DhSQUvkpuuLry+n
yYBE5CfSEkFy2WzdLve//xvI6iRoNTPu6ztUIh2Mt55B52pox5lC4vySF2cTh6PH
`protect END_PROTECTED
