`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dOM63Dgj14vmQ0433GImMjJMhwYkryozFhlsBvDAfe5yqVH8h+4rGkriuU3vuJuE
7oaZuGTK0rS9E0ks6tKmSTOTznAhV1vsfogWLTRd6wCqemodIbHEBy1KYjT5K5yl
eD3SfXY367dVc9OKU34e53mRFV+NvNkJoDmsFvLdzbhGpmP0btWrF7KDqCm6duSz
lJQCpr02gG5wEJxKW8JlAA/aECbw57GzBlXDIXBn1FV8P2uDeoszdpqOUoq40q2k
rfkvl7EgWcG0rD0q/bYCyynwVkIE3bZ7HqAjXMkOG8gwDbbFsNlFaCFIl2J+qNrK
YL9CHNF24XCaJqlWIJB1P9ajEt3SWG1Juer/2Zv+Tl4BL+nChGV1+7iWwYqJgy2S
ihxVA/HHO+DKcrSk21ubQGwToUZYRrByp1Vo4vxJ26EuEwd9Uu0E5qerEF+qRZnD
tKWHMVtwF2sZ1cPI3X044fyjmiDOmpdf2s0A+caBwNBAtnj/eNr7p1Fp0SH52wM7
dlI202KuyF5+4vCE5xHn7aq8jzecKyhONCBcoIYdlOpSuc7QQgLQiA5mnDN7X+x7
vIWwIbAT6S6uZkaxHV18CS5jS8Y+XzNWpnDbKJUOP1fWRmXtl3v2BfuYPNvSKfLD
PdjOIm+J1izJqvvrJp+/3J06cKtCFG12+gJ4i5FFXm70NgtOxo8jCpCIFLMYG4s/
Z7IjV6zbu9eW9n7drJqn4uJFxltw7XgN/zuEBeBeygg=
`protect END_PROTECTED
