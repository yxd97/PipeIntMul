`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5/VxIK9o16pRJrhR4PPDDvAwhxWRkpcvIDtHzmbdr3rmJaPOTRl85AYCtNK69Y0
K9IRrJnY6DcOCJdcQNulV+IaeIReQ5Mn3sR1o9Fpuf3lrt4xDQMfXC5eoiwx1t5e
iiIATZva2YMe8Q92aFF+JtU4PQrO2avuDMPvHTVzORi/eTYiXOg5I7mhfqWUH5KD
EFYXbZE5XhR4D5Mkuy4SDVlE+jhC+GKbgkGPWjt2RWuXxigaEr5cffYU2XkoAfxg
qRnIlO10duxAMnNpmYssRg==
`protect END_PROTECTED
