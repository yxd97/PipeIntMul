`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l5NUDmqikVoSiaEamxr80BNOChu5+fdipJgz9Y+DKnPUr3keuSQfJebloUvU8uom
RjpPPP495kDzrYo8Ved30RpwLG0VBiKR+Sm6+Pd4zIFWBFBa4hWAJOVCY44NmREu
zUJF8Y4xw+F7YXhz7Jomduw7th8xhX+SO50BgwbBzjvdaDc5zofHPcQ1piZOeP/h
M3YQiy+skYEYKyELUIZ+SKdxW0sb0dry+Vyu460J+kzlsDzaFNZYv3t8IQGUb8tY
Zi20cdmBrzsnpjvTXN5kh5nTH9tbFcfdy0Q64j1fzKdMBfvcq3rBDviV02X9DduL
qAJTIsvh9jV/7Q5M2NAKuoyu0beNCulcO3DeBx2BFng/FkN2vcKwbQOAJYhkRNPM
`protect END_PROTECTED
