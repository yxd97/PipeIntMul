`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4UF5OlarRQ96d7PsACfmicJAfroUBZA1/dWvNnhGLep5jasJ3BuS4x9oZYX9U4F
+W36hHvMJtH3xuQIvkyjxAiyUOKrafyBcRZPMbMwpdRje88qx86SmxwpWaK2aQ+J
vQHyK7oaeE/mf9S+WbqiCfcsQ1MsG9jIn5L5cfV6uDs3bJcUeDy6S0Yo+q2sSU7G
wLEIzjc/M2H4yLUyLxtxMZfodWcCnz9FZpXju9/qNw82Vc1FuJks56Jw696D4wh/
AV9VHhAMz7oh+x7mI3XdcAT0SOfDbzOhASpTJOA7VcCEG52GYYDDskO4FzxJl7ka
mHoApl3vDjEyL0AXehS6CQ==
`protect END_PROTECTED
