`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
azmp3crD8Owp+aHg4eLkYKj16haunfgZDvroS/wD8O0kX1itfnYrNhu8Cqs5o6h8
BfMNotHZ8ERue61QRmuwPXoM9dNg6TixulxPsO5PicEb9Nxy3autBBU2fic9xu9O
NAweNzYyy2kUR0CJjFQ7slq2LL4L3uhSUXdXW4WOsUDYGO8BIcUWIfT/dbgnLPM1
mOU0+UxEWjvnUmnbyW4+rHAUTa7ZZLYMTDZaKUsJkcdBUbkhvHo9RSo+1NzB7628
EXlhM8FGWgyI2m4+kzwQkZ7q5w+vI9H+E7Cpy+6gIwjK1/hdkXlY3nXVggQD4O8J
rb1IXeZ//+TMbRoO10xxBLxgogDRpOqwmsmGOl69wKXRmitjOx6RfRbNBVOFAowQ
NxIURc5fw9YQqdtJaaiF7VUiYswefYszIK0JWN3CT43ju4nZp7QWxAOinoKMnezS
lPy77yptMZZ3t2A5ZgGCLlWxGgKyORAaVkhnXiI5znVkrv2pS2EHqdw5TvO62AOC
`protect END_PROTECTED
