`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrwDSjgZQTkZsHOQlGu4q3p2gcHg6U8EjJRr3S0HlfrXJfXhT4/Bfc7fxdrzo4rZ
gcZEeSGTFxoz32qIZPcyev31na0ewBfkoiyhGok9sJNpJLBBrnA8cr6Cn777yJXU
J0J2row3VIDookdDItsv2TuP/zGHRYWDscuQQCUKK49kXA+YFG2AxAgcGdNNhTtK
a+MB2PuzLu4leeg1hpuxq9KFeAHJv7MXzQNiIP9BPW1N5jRuB2t70a0xmSDDD/bU
x2dcIVVvpTh1ugveUUnKqIrZRwyxbkracXt948pP9+3b2hrMsqA7uL+F994IDls0
aMK0fQup/wdNLhpD4cE+T2nCFd7xYBsCxcw8sCsp68dY+xBAhOOStV1AIHsKCVBC
T1LmCE1rjmUIIyK744Y5AGWAmWerGAJobv/1vn0Xc/L9U2nBydsQxX8d6I2leHde
Sh6p+mxHll3MKY1nJKZqAuoLyNFxeshnSlea7RESHCJ1kRsgbHBldf0MBrxGYyEG
ytvLu3Cgem1eb69XPKYBtaD6LqBocAgC1Nf0MVUkNg6roaLx/smQChdklL1yURMc
YBhEnzc00UY6Opt0vEVUK2v/8bN+1Pp5n6LbTilBBoxZQuuPbpu+4z31MO3vfLtJ
Hu1NtNZMZSXZZT8vW5+eDc4P94Mn+G0MxtJnPW9qReD1RL/Gh/DJpLi4SI1pv20h
vnxXlmccIkPMPehFMPxVCCbpUEbuyL80pGvyokXKOGmzEYgCyrF+p3CS2VtnB1hK
qJpYvule+G9v6NLigy1e186w3xPxJWSbutq+w7nJMgG3Ehlyp/xbpF18gZppCbiO
4jI2lNHflWOhBwgCeiov8g==
`protect END_PROTECTED
