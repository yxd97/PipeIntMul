`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/QMJzmIwWxt4OD07lI/DbS4PXq6rzvfYENug7T4IaTMz3RmuwZwyv87fUITznOD6
+Ajr7GVbaru4TaJNGs5ca06pF0C0afPh4SYfjbI1hl0HnbnwUfL8NSoBg5OZ08Es
E3w2VN91kYnYc9oqJrVvph8isxuSyVTr/r3V3KXrbhthJ7Os5D75u6mazO4DjWYk
/7slkBHrJ+2ZxEtvmSomlviDvWEPXQIFvdp61M8Do3J3GUJMo4E0ok/vdh1jaFsL
IsKVB0i6yL9pe1AVgYdixZ75/jrmvNlHe3jals6oAjnNseBeY6wd4vqFguUzkwHc
7364MnBNTumAsXFnjCI9y7Mn/shC/FVGNch8CFhsEMSzUthPT+dc6XHEX08QnlOS
KEalBcifmeCCiNZ+ITmMiZgHNaLH8J0Hp6k+qI+uqpQfid8m0BIj94sQCgByN6nq
4/sY2RYNnJ9KJgp5nQgLMsL8RAQnLzh3nES6ahTmnpjA2qIxpoO0N7V6DOMngVnN
wHcH+oMopuh809PUO4kfvqW9Z3BWhw2G5KnD5wCArTZveHDTcLNH0KH+kgdocPDf
8zxxAcpFyloi/A2rwLow1i+kC0HhstfJMFRebJ5lRj0=
`protect END_PROTECTED
