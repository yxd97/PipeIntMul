`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1QoDsvDVLxeESa6PMsGag9SG97MoBP3SSTEqMJMM4u0oB8NLgjuzLIVsRJYXnx8
ztJ1uzwoJ47a6W0oxIbYcMMx0opsJVN2gcH3r+s25Y10y4GCRaiJk2tL8OqXPvHX
dgSLjMYlxZ645IKPmUlO/yM9OTPD2KW3pzhbBCrX1geHd0i6tzAOZpFCqrUUKRDX
Os5cb5ECYdfJuNAu28KIlr3igVlMs9LKwshMzN6WDdrHEFTYBVHXGUNlhT+itx8m
K1hIotjwU+pXFmBR2Nsn2rPCXdyxzliMW6jBkXQKKPJimPu4DAA69VWWIEN89F8x
NrLZTu7Z3zCprSJlLnmvvI4Xyjt8uSLOCm4axLTsjh2VCvvfdDgoDyzrAT3c8AWK
Uc+IvEa627dGC72jQGdUr08A7KYN+yMY4EOsWQ+v5zlkMn7ejZzqLB+8qiS5zZ1j
ud45/SsxNXFRymCBGw3186eydrUCmOx/JMcirYFnJ7CHxHqVWdEot/aeXvLIE6n9
`protect END_PROTECTED
