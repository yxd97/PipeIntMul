`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dad+CScLkOH3dasGV2sbEIwIfJ4vhxQ1DW32xTCXif4JHwylvaqu0RJDJHsPhoTO
ilp6mtpIqsDOgbcarg/Fv03r04OqeIiU2XXtKvyDo5W0ClWJlcg8QUtzfyPQtei2
6F27C44v4im+fFTyUXH0HD7j113W673t1hOBI5w4ciRIPjPyWguaSkwnxOm3qEY0
ravHn31jqVtwb1SCx8ITO5MfMdmqLnqNXD9ntiP0/EfHQkCaYvdbFHRIYYY6pfqM
1UOjsFj5qAWDtNGpiJexVDxyyyDjzZfw00FLpD8nER1ZC7yg+L+Qki/Y3F3d8/5B
7/WQnbkY4hqkDabcLAy8PJhjrNx8TQKTXADGJ8ANDwMrR2YqYEX6ml6lXOGlVGH9
v0fryOQnysh5KuWnu6QufA==
`protect END_PROTECTED
