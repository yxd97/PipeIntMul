`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKRGx7+oK0PBq2pabLkNIFdV16rF1N8ZV0PY1+i0fXogJchJhPD8KPf0M9u/e3SK
jYZPA2ETtKpT8qG6ieaadwO4/GlILV/OoFiQnZ7wfa1D8sb53oLgwes2GRZy9PiP
dXaikHmd9X/DJpBXB7Qrz9bu9tODicH0igkwfs2F7Iwjm2F7If9OsLlbauU96VaP
OvYbXBFwvOBfN9KGmjShUOR/wE6S16mKa/pyGcroEyBIjXV50seVileEEdi1FY+s
G3njgswFPDDvPlID4lnNKeqlUJEZeE9W/bHPNpe8g6BzAWm+LHC8mOQCEbKnFSWy
cgE0h4+yqmZounu6wrM398LNhc7ZDwO5jFWdOaiD7YkeJ0L1zE8H0Yf12SPFzEyB
0SOOoKvzRHIqgfTX0V1hY7AigJbZZi1x80Eb6W9WU/Aw93zFag8q76V/tf3qU9Hv
J/OO6Q1TN6Xucy8d+nIbNn4a093zZTHYgOaj94JFACQh/TQDXWgB4MwygwOScIvj
`protect END_PROTECTED
