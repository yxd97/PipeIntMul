`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQ0zDf/X7qF25Al36dkWtrbuIhTLpnTa3vBVPl48iPx7VMRJ5wG0wA1qgJtIp68w
5BDQt1pRP4TvJlajCLznrD84glDnTCI/kj8Jhl4gyOb9XSQfi6upvXaei6+K4FPL
139TEl6jLbkGijs4PN1wlJYMghvW8ZNvZ+8vxyqRLoTu1aEYzSYut1jQJGHd5k8o
N4MP0IAlyLz77K6L7quXDX6pZ9bAfe9Z0nIUtKpvhH3mEDZECF0/SbRCAYvXtZn8
wGNNfsvj0A++Z0er2xM3x9HMqD0ddSKdHVFZdilRNhzjrG3Jz3n2yNAGtZSVWKdH
VXwg+vxUXkAfAVhKSvQBjhGHP09R5dtbD3n3Yoyy+kUALf9+E3lEC36mQxch4a0+
Sd9WJUjQq0lqMN5HXYXIncpNmysGNP5qDU8hRuFmsMzpVrbMk0TxnQ1kGH8srYKm
TwyYQFm/7eoi2r9F2cASK1HGm5ZiXC0PGw0778rzb5dj7910r6w+8BlQp8Rfu/XP
v42EphmOTCc74G8aIFwckXakNzRaZC3BsJU7rTTwNYhS64qLvHfHIuaBkXeVfTlQ
s/Z2XOV9cd7aCGBKD7xSuQ==
`protect END_PROTECTED
