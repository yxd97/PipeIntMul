`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p26BH9qeYGiDEqjC0+2RABvKKaglIF7oiOxwrYUTnJH1FIZzd5i5bzVZcMb7TD8T
c9dw7Wz8WyASDHAAOzJQN1bYJm/HRIfTyIC6KpXnX/x4YT1HpRkbQHLRvovaDkKa
YmqOQMA31yUgWgT6Ixt6Sp+8vWICtb9LZCBFcNMyXqAROdMaBKxsLqY3y0ZF5FNJ
MyA7cACKa3tof5fVjsoiJeFZ1LXQ6nDSCy6byacvZVIL1y76muCReTDbkSFi3tjw
P/4CH4AGjOu+LXgwpLJzNoMEG8CaED8RW1QPD5cnuao=
`protect END_PROTECTED
