`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Io56lGuBF6zLXaBNYu88LUZBwnNP48eQ1Sh+H7BXocuQcwraH0MlyCicJ7ctJq1R
UDWGb/4PBxW/m4VAAtwb2qprq3F99Glfq9Q4mAlsv3btv1hSsYE2fbJ+u6Dbk0vl
ZKVrOE8IH/cUYog5a3eMUxRx4GKsTG55X0WdDMRskKLtpi0Lirs6hli4Ovhay8RK
Y2nqs3gbC1mNIWgealbMCRcml3gSSbvBCiKAeHKLPyQJKmrkt8B9JZ6/bzQoe6AC
MEnHiYPRu2s88JEwhxK3OXmFy0PiTS2Qkm9nQvLW35Ozl9PrIsNv2Tkcqvsvz5EC
EMTgSBKQvSR/7k7m5924ModavUym3XFQ+ClPwNcR+/gNU88igYBnY/7Sskf3lTpe
vYYF7C5tqh0RVCW/Z46q2mgFSwUbIGmSdhaGk1W4Mn1972wLxCFlNOn0wRqGVUVh
gONrCUCwsT5QwQUz+fyH1yrlCRrc6YTcDZXYbdQy3020n8Jq+8FGmM9iR9eS8k0E
kvL0ZrZNPPfFacAhwy5SMIiF5nmVgTq4GUij8E6v993WUjIYcrhlNgb/d5SqL0g/
`protect END_PROTECTED
