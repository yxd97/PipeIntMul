`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LDLO2OWByzEosRCVka5YWx4lhk6I3DpNs/WGSt4Xw3TBIdGPqyDfFPSEQ1fmEvr6
IbvTHhIiaKwk7pf4FyTHa+D+ite0E+KV4Mg3ka4MZC9M2zeYaR3ozI6PRE8X9I5h
IJqAxU9ogSYivK27jM/6+XNit8r06/sxenOQmYuvPcrzbOhOINfJEAxtMFOLTWwd
XSXLpNYrlSbdyH/hglPRIdG6QUf/C1Q9R4TowCqneF/iDVyODZxddT5cfFxOMIqX
fX1rMtpx0d4MRlpfHpW9ng0iCF3qPdLkWBw+OunUBQhGsxlzJqbp7VWmmqluWg9u
1p7aY7T335Jw5q5DcIPT0aHkALPdO9dKNbJ4VCCr6jya0XCHrW+ML0VqguZMY9gF
g7GqPHTtdZxlW6FxATmCbYNsGempv08CNoIdO8SO8O+oaY7H3cz4M0WTg0N13Szv
EBvoKovLypMxqVHIskTEWP/4GDmyAUivNiUndlBi3VPToP2EuOskYoMRsW3w28KB
LsiX2cMCZ4hHAPLsFg8g2+w0QRRGmdrhtJXvGdUf1Rjlm9cgCffgnTLNhnGvY+ye
qhPYQcfZsOLJilAltlZvj1njdFV7XQIGUMBv9JZ1+bq4idKF4Pam0hr+zvRDXKX5
Ad5b5ftmiLI583safFLpbd66rGU20QSpT//jdKN7dw+ZuTG45+ATofuotjNndRwV
/4S7xMtr+McekYSQLI9+MuC/fuvhViR1b0Y3wkVjs3i8RgqZdI2CSOiePFfsuMtz
+fhTeQs9koUWtCjPuDrInycMV1TVdin1teLqS5htg540bWQZ867+osb1+uJUrmQq
AdprO4wrWC9vY4IIIhY236bp34qnttgT1ZhEdTRKWVlDWZI3Bg/4ggRC6Ssnz79m
AkBTcjEixLsT45mqQa4noA06LLfDy4Ykz64WkolqgTC0BTh6uNUamd47wus7Xe5J
g7pEm7Fi1+SgcaOgRxgbNkRZVgbaNk1/xTbVUtmlbjhviDPEjG31HNTgmkAyJ3qs
9rwCy1DOR94wi2Oe9jFAIuWlP5NUVhOdI/lYL/psRMO+ZyUpufl0jd+VNp1x9G6+
4bb02tlffTJvFjUyXQfvMBtEUambCwJydXHg1xdxygn7Uf9FFnl8ctGKEiNArPrM
V66vQt7Rzt4lg/Lfpp1DnNgnztZ0kiBQR6MvJHtkWR8YcF3tvDB4V/8qzGv3RalZ
rfwrjnz1at5PvNlSesdDhQbfm0OW4QkpqVlo3ne+Yn4s0GE6CO350eH3TZWhcTst
uPNVRjbupidpdsVXKKFAfmVdziyEPU2gV7Lb0g99QGCXbKY7S8J9nw8AUxFvRH5Q
yYcq9DXMF7IUHXVsJ+dN2IKktmkP+dBDBTdQmSNl/SpxVyqqODQcUlBhA5iEU6O2
SeQcg0jDAr8+rlDkwEHmTIAybVOO+ph97lJY4kpHIdnb7UnotfbIYqDFQlhhYm7g
3q4Oq8TFvcgnMrYLiyQ2g/vtlPZbW5XTDmBBN1jM/Pqz5nCPV80GloY84/nQBWvd
tXvo/UXasvWKZQCfiPEQIBwFSjKD+J4POybffHHgzV4M7ABA1cnapsiwRXuTH5v0
UFBY9+XIJwM6Xci/3QkMOKo06Dyo5vgLmr4nthM6OZ3QJdGxxBKQM95u1vcHHzk9
eRSpxsrNo6heETn5RX5bUSAFlRldwCJmdmr2/erf08A1FxIs+3QcBDerB0bqoj5c
DK/Zs9hLGa2uYzKpADX6xgn8/vff/SOQTN5YKETwiMQceMEWvtrp2S3rggo2OIFP
vqDwvU7aixIYrPO05Ic6ysIoWWeQpJ/WdOAtc/McCXAykqKim7VYCp6XkViVxI1H
m6BqRfrcbwnGInhxY/DrUS8+B7TquuGa4rKmvod78eiZWxuM6XOgcYRB/Gju7k5c
rbOF1BdD6A6b6jivzdM6ts5nGLr7t7jFGK7x/LKDpg+VvZnRnnvimo8Qn3t0URn+
PqxzM0JRTONVS0pHMR3MiQxzTOP0SOzNlWfioDDDWrRJWeIxlIEU1/yDe1LA9g9w
3aFD4qRRmrxIZdZW6ZYssXGTSJj4PT3f5kIO/pM8yXs+4c1Frd3XEhMu882x81du
2te6s8VaxRwsDNb9pRzVbpFQlwu1GxHTHvcVji/PB3I9W2XjiDKFv5ctZDCUSbbo
V0K+FvT75Tz9OJSJJOJzUYbk79ut0+cu6CROh4naiV4/f3uMOuGKquLtgzxVySWA
L/l5c1jzLSXkExeLfBX1Rc5wRdb5hzqFNSMImctKvwcbkbln4yJVX7kMX0ApgrF/
Hawe1jr2V+dslU4ejJOus0SqdyxE5sdwkqByOeaVr2Jv+mFZtpD6YP+tzsfbV/Rk
UfSQnNQL8dMGimoNjyJ/RC68hkDG7l31U99NLqePUkcs6gyXrcyy17nsna4YV5Qj
pvst3oqXis9RYjgHPRvLwpWQ9sBRooQT4stTm1Ij/SXfSCaBPSLszQPOi7+7Xc/a
0DzU7fHtQZPD89cv/FqqZvmHB3MPVMc/zb1ZEb9/ROBaC2729qCCo/FqJafkWH7w
KOit6T5747KPpNzhj2ger8E19oLLvKrk7HTTHxWJSjmcJtHPkXLRPpxR2IXQ57yE
R8ycQneUkExNkChIKU3+kdhZdBS2h7uKIyjV9z7An9QOdED2YsTQzSFDmuI0Mek5
sQRYvTG+VEK9haHyzjLSbUR4OekyDlkOjZUtv0VmUPArhJhFoGOUFeePG36+6le4
fP0rORO9UmVNeXZ+UFhowV0aoi5PmF+BTEJXaLey6fZ14vuGGiveSXhsUqbo4t7d
97rZYQ/2ABw1sfGnpR7mXgIb5DOMFV+ces5jkECy7tB7g5warOAGrAcCCWDOWrs2
q9z1GUjMwPMKo6VrE2vFdoS7/g0UZ/n3ijhwdV4usBgfmu0kkACYdh91xGF3fLNv
VT3tUmipV8oygK4WijDh9C91SAmZNvD3KOGipPG3imURHBzi3BuvDlcZBBIJY1EL
iiZLmvE1lp4OM+ZUSrbnudlZV1HtztW5w2YXCRhYIAi3oYco/Q0JPVQDX5mDKhmi
mEloTXbY5TGtkmpDUKdTnmqNbcMbzKpjFmlD7C8HWGhPlHNtttQr0kNxSlB5AbNf
v6dxxFEJUfdLhAEeUsJFjW2Hy2y/WRZFJRT+MDgISAnSJXoVU8k/LTWtdZejAr7+
WeN/eKhrqbf9tbkRs0rVRVMgWGEDjkjYiYyflMfb3o/9rAHMS0LrAByp5W8yazXD
z4mn/j9Iy69JrI6DfYHguxVZ4UIgX8zHRh0Pr21iqw4ghEDYyDfXkH60cT7WeMXD
PXxb0zV2uhsPL9w7n3RT2hXtjrYDaoQLAmrQ55XfitfkQrqSTNjUjqC44l27U8TN
qkV58jZECMNzWF8lnpk2Kt6rMscuHIp5MFaHvbXi1n6is84ueJBvQDTuJljno/W+
dLZIA7+xChAXshsUM5LWyoNoVgIPM2c0ZVXf8xYdWg6WoMwvbgaCCO9eqh/N3fh4
yNAYGTaTL9umTYHYW51KBTdVudPlJD/s+r311Fs+WDEHM8d5u6zZ4QX70qzDC8ni
1qj/ptZecrAGLmKzYztFhhS8HbwrJlZCbyhMNWwrd5gG4vMRIBxvs1TB+0esimSg
lGlrQ+oqVWMjgEF7SR1xVz+59uLi7782L6Umzy2YpBJIVYjrWAt8EG5Hzkk6Blbs
SRQeAyf7NJsVto1Ok96Y32M4m4xMjDGB6bth0vQW+6N4Os9n0SwnK/KabTk7JP7W
pMUV6tBAkuKDw6Qq6wBEWR9z1f5G/90ttE9Tt5bR9WbBjSxMyOoLQgZrGPfzJCVk
mnri251uF+eH8JjI2YEXPv7IM0Hv2wqLSXNu8ttPg2u4LALqSJstj/dQ4ZYuBqNP
jfVTqRUyADMAmJNNohqWVXicdZ5iEY998FS5Klpbj71pQsS/RPM9gzUKEDYuDFIC
5s1XmR/Mn+pnebwBGnpvFrY8RCrQ6uDZM0aSGDpQL/Y2MvGh5aiKURalpX4TxFna
eBC8wIenqU43JpFX03x7gRYrxLc4UtQbvool6NvQ0H0YPL3Xsi3U6rJGbZDyU72v
w7tMrumcjmE8KyWSZ2/ZeUUFdyUPNtcm9s4EdqM3oAFGTNhI9uQJ1vZ3x4H+vNbc
zxp5Tf1SdSE1+yA/pcfxr4i9tSNM9cREkExnoNbP2NSuUds/TYNLb8hdh/xAWfEi
Cn7zfWVqUT9eeGSHCxo1YK6ejrvTTbjV4lyWXRqN6Sp2NyQxJ8I1PaR7mZ3KWKzz
1hU4KLy3/TAwZlht2q4Cav8si7z1LKp4qoog4nsVo5PNEYK8e6OeDR2K4MR992nO
znAl3lfZa9AvtUYYYpjFZAhvmQ8ci08zDJgH95jv/WS38BzesmVGU3ELenE5PgpO
0cOCLTTBuzwW6LWtOUCu2xQlxUbfLqJmYp7rjogara5gyCXvC9xYLGKS/bSbwztD
B/BORQ0YXaYFLZNmm+n6SYYSAGxExFVNKR7WnLdVoXvy5ddfgor2YEVFQ1yrGvvW
AE6mwBuCsSigTmlfebRcuDXdVbtFVdPyqkxhwRFoyZqV8EWNg4s6gTwvuhFjhpNz
D6OqiRPZxq7nKV14vcu3zB7i4368SAeBiI0iNBvhp9uNI+0axfKb9dbSQel8VMXC
jX8tdZYlFidaqTX7oKHA1t4iBeQpjHzO9r2nsYWCQGLQ8ch9MJeal9q0eUH4dWhx
1zxJ8gz6QrU8CIhLxr+5nJJTMnPZACThwHLiQUVcxWSFM+2gYpgXJzRtHehoGmzW
L1ARKbC1volxDCRjg+jY/wENcjurD+M9V3LD2gWcnkNmJ2LxrNT2doguoeKudyxg
FMVz/jFN+kN1EMMKD96HZ2dRCRcaeQEksj0+ZSU74+wsc4vXZF5v8renx8/SrNIk
SAachOkONMwGRy1n/jbg+tSBYs3WZhx96lrohp/DMA7GxTTQynsydip+P0qWKlq9
fAvD5bYZbUUeLdHQP7nHBDDis98pDvnSiHzCyj9ng2Jm5CknjPi2TGecQHNf4Zm9
2Lnx5ZJoLU2K7SRgsJkqncrgf1hVoCVRDXYtRGCgnT1Xggarmnqng1DD0G5eWtBJ
ISXVQIQXmswuITDuqLvM/D2kJtRJko1hZfB/pK286v5J9wjlAbxNUmR2ubRVpZ+l
dhagIUF3g4dOy3tfk3EzWQu3Cad/KFtoInW0V04Igb6j9qz8WmqtwNhuAiuubuO8
0513xLygiIrCH/67jyr0q8YQ5/665lhUwfbwP0YoJjgwVmxvnCV5BH5bOy/3n08C
eZZGcspPcnnnVGpSM41rnGNHyrI2zY0jdrvYtBZZpzJqZQPgaL3Q0Tnh2hthUG6V
l+7wIXs80ueJY4TwW7zpppeb+eoHBPOASpdxtT397ySXlK2Isr7T4rPNR841MSyk
Ahe8opmtRN+tBmKlz+m6PrbJngvVIF6iK/9OZHOe3MB9v9fk+H7rLuxfAIF0a+DR
jLoakia3V+O7Uej5dxC4b2tp0Vscl2OM+i1S2SXnjpw4RHZqJB7HcLVjsFG1/EoT
UkFeooYoLxpfaLN5QOaRGevO+/dFJJT05siD1+rffXk971oX3M2bkqYVjVoNxpu2
1iPCOe8ri2gJhzOysa9JE2XMckSFu/32yGMgW1oPndlk3qZ1pg8QlcLj9EsvHU/p
GlBCoTmMJx1sK9R8rriA8Tr2cwYfII/H3mNScUqpymfVMenlic5fkde4y4bZKH1O
ltfpr6eVwr8GewuRsyg3u6JVNQD0sZ4z+2NSUJbSLiqn4nAhiJYtdigUtMeh/qhw
z44NOx7azPNUydwn3WYjB9ruIrPkGc3BqB4erI4v/GKyiAW5b9sZ6GYOa7pQpsHn
0rwIYwpYmlnIef5Vo2XdPALVzQKPyw4ZvyEeDZA3waKaOhTk297KypDjNmsw6oxs
uVHX0DxIni5nSeIlsCtuwBjHjtv6yx7PWJRVN63bBs9mM4QgwHlPN6wb770uQA+e
SoXjS6ltK2LUn/GdKvhaerp2dM4aI99L5Yk/JX7MXGwBLeUcT3b+3bEuqXmVwPtQ
FUp2b8qdra1qQ89cTUlPUjXv1z5ui5fRKx8zYKEnPvM1GVth+zi2YgdunucBUGW2
iOI4wKaaFDG0HfGNwJaZ2RqlVlvAY0FtZJJyLdKxUmgNCgikEa6it/mHY8TjlSn+
BfQC+12P5l3ozYK3rNGBBrvqLyIv7ugSbfSx3JmCPjWZJfKV+1XH1h3EnBVgKu/o
bGH0mtbHQ49ChhPR95ZEgY4lWp0b2X/d/MYTTbvC9mYLnh++rc0jF69YbBwGPWrf
F2VTcBWxR/zhnvC4cuYckXFtrRHcswDJSw0yesYjc4r9nBbxx1ZdIcyK2rMJmuAY
KavLxlRlU6bNL+0ILFxcFCr0zxnlthEFK59NGXVxA8jRLRdRfcAVmK6X8tsnDmgG
KlTSsPtiCb/PHlra26sFDENZvaLZkuJa24aezuuFWRN9y36CRk0xAmUFkCyEeYPB
kLacW4bPPcEKJNIvmZ/yiO2mclH6auO9niDAe57uHFJ0OvHBVQYK9tos6qCNHRZ5
CwJzkxJmUE/qyL3XDhvlwEnhZdxa/fhaXrzTSMyXbXJbQE9rmmOWcP1HD809VecQ
rqdcw50T1LoDbxYn1iOhxlvwY671UJiBKvBg+EXBq8lIHShXuGAmCu9YZAAsjove
WPV8W/UwlcEFr8HfYds6MmMob6hbV3ZecppYWoqBizR07X+4419/BricPN0LHGaJ
DmsWHI1qxxWU3gTRJGYosnJYc25qKZCilRUtJToIJZ/LZerVvN/G5Rtrrudj1B5Q
+NQsjFMsprQipwOjJX1CNOiw86v9RT8YyewE7dqZSc/P7ADRConjTgm8WHZNg+i0
YFt2iyBWhnDj6ZEnPh6APYDQ3YwEXnneSOG9HH5NeTSOCJumCcNoV97+9T3SkvKy
56TVniAE4VT6mOzXjhx7/JcGmdwROzBzRBJtIoV/0B22Fme8fH2wJciqe5VpF1As
1W2x67N46VmnOqHlFZMknBsRUD0TcRbqfz+W/JVOLkkTJsyDxC4avhEtP+NiZPrW
FhKBX2zoC3xU1DjJXu0VL82O8L+jfFPcSi9AwkpLBAdj25hV7+mhd4VGZomWYYzM
JkqGV+1UTqUKkr/bnl/q/HMo2V8wxy0N55TiqsNNFElMHAByQ+i75EK+3tjCUtZZ
NUkXEE6hgYTJN76+tBOkVhsPaa0DSS3VnK8IfMxdZNUUnPENzKlI1gvUe+VDrrtC
COQ+tvVepbNRuf1PYkMGnYVFyZzbgvdJYf/CcmINgGPkH1RqUNLGFRHxxS8ZRDV5
ooZrJeW/eXMU9tH77qSiVA/4XoWQDRE2UEmkA8Zc67Z8FU6JxD6rbmN3ulcImExD
40YG5EqH+B8QJuI+ImDzleWCoK9zmelNwQU2pe2wT0o10X/hmrqfspwoXkobstvj
e0Clz58sPJKWLrr1vWUd3a/KCtffoqBCOQFHIUJI6YcanV75v6/5tCpyfl5Sey5u
G0UruE9JaB6o6hD3BZygvPL0m+5vpG4N+sACag5vCpQaZvMx3RPY24CCG61D7Ms2
Mzzx2LhHKp+nK3xCBu+xAuTJGjUiDrYKkG40IPWSrQiVmCQxPHml98cMyNYx84CO
Bmc9J2XAmhTwjHjRvsiN1Y6FsItBAcuVATiwuGY4JTNa0oQpVb4wPT1fSeNA9is/
kKEX1d/+9sI0MV7hlFjYVrryOlQqn+1ea+COwmWwtwjz3FOCaH27DDkgVH6dmRgj
Zoxf9iSx69/IMWkz0g/5bK7SXI348b+/lj1ict59IhzXzLnSzQ37cnxQiyoRjNfZ
0nOCK3xnFWye+7tRtEvy+iuHSJvur1FwnAqqCOcC5nEFdxLv2yGnmWOdkFLhSg6U
y8050TKmMad+wXdCCcv/MrD45u33AiFfHz1JsafPLcpCgSPbT7H86zAeZKERBqRu
DmfRT6i0pmI27YReF9Gc3mNFz/P3mQDgfTeJXN3nQbMFMGhTDol4W6m3XmgJHnfh
V2pLXI1BoTRF9V1s7VGnSS8IV/OUKPpUEgoWDaFHvoIFWp4tJwyVt/XqhFLbVPq0
miimti/8m0r/6E6z9XSuXgYmBy9UQ6iaCgMqdINJwS0f0jnpcyHh/OVBYa0jdCah
6La2PdFh2jTthnWzIrL5G82LMJISuTHrHKl6ZTR+gEoQVf3cWgAnvOGJGiR86v+a
ACGbypQ/yjVfQbLB3/mU24rpi04GCcXARnn5wYej/GLt6hTGnerL790rRhASQRJK
/q7h4Ngfv8zKR1atBbx9NJR71wZvPTbXGxRpyvZeugH6mTUxsI1UbP6+mQf222Cn
Y2lT+ApKySyt2uBTTVFO3DP2yV0JdKQQtCZ8OoUohfaw/y+1coeSKdPdD69ZqAe3
X2W3QE4KDqG0vYwj7Zuq80wQpvrnI+4vuanfTtwkajMRAuKUpDkGF+OQ5WtZ1ZI2
X1uSw32YqiKKNLgbRBenta4JZw5MZMgFyORfe5p99o6cHyh5KtmYtRwwZihHrND/
B0X8+QFVBcluONwcYfYTOr863+EDUMeSDI+rk/S0dn+TJLBSvfXBx69UJLzV/2cO
2XHwDnz7hRDZ963aq64xcyzTvrW7Af9C7oZQ7BV9W0kyi2pjtHabfjvZpiTWxW8m
CORdOImj8zXRyx7TMjcUbBLi16jHDLtHvS31F12a/o/UtAdspbpJlC/CX697Iexp
ivXbBwCn4xQethPSLt7LS+ITU7lVb0SsoMsElhtTk4L4asKYMnupztPSPCHm/ua8
qQjm4cQVLqb42rZQsBPtUrQJJoK5SQFnS4gCrH8ceqal4wet/dQvZC63HaB0oW6K
NaYPpJ9nHhltJSOZUuxXBdl0tJ7USuV9KhtKWeM1Lb6Ss6SeZ9WFX6KeEEb72oe8
ueKvNMS11If3Pwu41V5QZeCQ5e7l8sugRp6r2FI99Gu4nX39LMi7DX2XMiE7R+8o
B6wb/4RcXrWQBcsBy11n2C676qaBFTSsaOFRxOqdYyw1RCq9q/pvB9izlCRsSCNZ
YHOlrPfg8zIlpagVoADPJM+ZbTml+Ig+8XrxukCapy91v1lcZcoxdgTRjfKSSydH
iudvq649CVBz8PfLfuc8Kos3tdiYElzbg+PokJxGK9+NCGlP5yaoyZBFIi0b1n/m
1rK48dhiaG/MuJrFkDKvtRhcgzOha9NaDLBFJHE7UjbzjBGCqjUNix3zKNvpGNPZ
/sKm5DymUG9Mz4QJBIvIGWq0rp+yxyWqL5664gLmU3pMERpYo9KchzzsubIBfC3T
+M5AuuBb2OqVnwAWUQpjGaJ4SAQKddbx3AfN0vOE9XqZTqGKuCOWzAx2rj+SV7tv
2Dk2N7BuDdvQMaeiRleJDakNV25L0Rv6tnUd+NPIM3o/yVtQiUOM0kXepbXpmpDe
pognjwZYlT58gR933nm1OA3Fp/V4gozcT8I5iCkoyzyxzMwQYVg3JJLx8mthERLx
YdYsdYhs36phniOlRvIwS9tmrxLPw7n78FW1YBN7LGO4+VbkY0T1oHcuiiMwUFKz
UEKKLSkaVGBQMgHWt6dvM+x/xnVT/8oU/NB6pdGh5Lf68v5VuJJ8f413Vr0cf3Jy
yI8Q/AqmqsWNnozPeN3AKyb+hCp1aCpfUQK5hwQ8dTBveSj1oabR4n8eZtnZt/+C
emGlJYzCa8TmvzDfvrWEVQn/Hy+Q+V78E/JRXrP24k9D2X7AGUWw9K2MAogQ5k9i
fRriDbXLtwolgciopKYYkMOVANXXMZolpUc2W9xpSxbTkrD8OQTze9ypVyfEeJH8
f9QXaK4IYbAmRAEu93SGIaUgQerAFjeT5pBFKyZ3qxOrFhucT2Wqh8MWcZ/ePED0
i22wmwu9SjLBX8my1kx6kwLyn7NcKrgUg51Nzipj3vDhDXqe4UP2hyWeiQO4ss6p
CeNlymbLxYLRLr57ijJhFysipCoM++Czmp5GbwAMSUUjek0MzUppnwqi/g1IIcNl
cOwU/U0IC+ywnI9TW4SdrdzaEDYlifgVtKkmREvL+eXyUuXV9tl3kbyEIgqFtVeV
12ugjiooRhH0n6H6NRFxItoKQKdax+V55escfzEodSqyBgeJG2iZX+JDXSfQPbrH
u4gOvlGLey2LuRp1TjiIMPOCTRviktz++P2yg5jy/GwVTEfDKjb1n/OQ11QMASZq
mMau5/6SCIyQ1r3PCb0r5q8WufFV5VDIcmrWYNa/qYhCOw/sviP20iFTqFP68NDf
rJbuiPO6ZT0/Iiib3Fs2gRJ2WQaBPwRF1RZ/N0rt990Dx+ZiPUxYV4dRBSnYxYeK
1/ednfqqgyUm3V8IcY2n3vzyF0GAszuzfK30jMrwxegM/OMkhRjVucCNsmrBbSLA
tK8P67TJlIycaDCf9jOL/3lk/4K4xj4vhXNul0CRGxggDBIxN3DKy38atJxqi/bf
Bp/7mVrzFYdW6DmInlg3Zm2CWHKSFFoBKZ/oNqBundHvtXFbjPE5YKc8WwXWH/eE
CwGghMRcX7qCTBiZ+eDTcaS9xEaaOCtLSJhb6eYcTWyTLhQ3IpEI8MLVSDosF5cA
Vm1v3ssYB+iRnetOGl+Fr5T2zfu8gDQzapGmeUXXgVFGQy197xRdiP/lgsH5O+hC
vorIzfpIERrXC3ApDIcb6qU7necH6Y5/NCQl/mD7LoggnPj+xLmPpHtsT1us5xKv
bRyJc5V1RjkJbRWbN8e5BqxaFiPnjaZPW2EvH5SfLYLe5LJ2286baxvViFkm6c3g
6hAKiNUI/67zHKo025EVrxsrYBPxnPevjggBvbzlSoEtxnrKo2YB0cWJUE/twER2
gSQoyL6Oi75HveUsUe5zG0E0yBJ5BlD2vIVLBfFyAWt6kY0/PZ9CwzJZ/fMejl45
EEyyWenM2LsNI1vrd2ONZziIBveFT9SZ5MHbuUGh001bRNBo8Pu+DsOGUZGzuXPA
BULYynRiqxEuw6sunWMBYNmZfY1sSw9GUX4pteK7IWyZTmBFQsdEfisY9EaPqcjp
I75SIhP5/vRzCvO8tudC8wWdjnOfBaPD4YEpurwfq8CvrAejCuSthxy2hOOLz8B/
HWGvqWtFTIKPkiEEAEy1VgpuZGkhVv9yE+980rSGvJwNkqajvMSRhAbS43iHcTFY
z5BXoWxX8uBDFPkC1f3toaY/YCMstc7plUAcY0lFnosJPVJuauilNqkALASB2clG
qpr1pq7iEz1HcD7BV4FwN6VwqlAfhQWbp+lP4kT9nAQy8b83LoSN4WAgeTxbXy0z
pMAQtbCUa5eL/S5lEPHHq+l5AxeXqWzhwk4aceeSTvTULlGXo0wi3XauLB8bzbnJ
ZCh9TNiX4XTdfBcaZ9IN8Oh+/Vsdz6MzVKTB20hIa67q6m3R1uOQ5va520+l/3tZ
DLncllg0dMky4YMnYtVrvHUU0Gs9o5569Qo+7a70cehDTANJtyIah6hK+5OeOfON
EZvmLlFF/c/0iCVeY3MecputFd3qI4eGWIP9IpKELaPsN3fuIGyaVSILlXz9ThEm
q5rre9I9fDbicHQIGOTp24wZ0xuv3sD4OYNTy/SyUC4WL23k+l7/nSrfor5rmQwB
G/GeeHy7q5opuCj6kZsG63JPunbg2jnRDtpvGVYT66VeHwCNnaIJ9tnh9LY4eFz2
tADLXydEP6/y1IUBIhJ9yMVtf9zkKYCmMqsCasOSxgBXdbPYjZOOQA29e6vc+FPd
2k6RfMgWePvuUIUjyW7JpbazehQna2iUOOEIdr/hrqpv1bwHCOfAC5148qktpTnK
2Ym8vYgFCmDZ7yWVYjVZUnWGz4bhq1/TuAsGi9LB2iDt4RZEGU5lF5W1OhHvxije
XVGywSkVnkQrsItA3FQec/YrVK8yDuUwtEZwrck6fnAbMdRu05ySdsMoNJVjAPGu
l6ePPa8A4khyBnm6CWzxY+VBKC1xeWd7NPVmmgWBEzB1xAqfAH2dD6spHk8eyHl1
4++bFWdk9AOKjU7ucAzsAmE0+83nIQ3iUs0lZiRH8/d5wXjw8XMlZTSB11RPNNk1
+mYpT0wlF/a0RwYCTPnPov0nZrSlB9hTpLExGQXdzWvQ/mD4V20FZ/0IOvVw/zXK
X70Xf+Z8kOsK0kX7xNAWkEDZwZgFbCvC2B/vUo5CJs+O/6VrP/by3hMgVyflf557
NyKjOWzW1d1XehVuXeQXzQt3zM9jXX4G0HT6rp6znG8uwdOk8rFej2lgPljwLQX1
gb5YDkXEmbqLnWLywDA4BaBLyES3UKvo3dod1KUPqN5FDissgCLMWSBjo2C2e0+4
Scwn6+SaGqr6IGwbmiqAs85L/ywPS+0iWRY38erlGmLShbvG2kyDmRGzmND6x7SE
D5LKNg8qX+uUIeDxeO7TGxmJgJ33hr5Z/BeqKcwDdQYhZx4l11/OpqTmlJGa5Y4J
F767KO2jmcUGgIfg2Ea1leAVyGAl3kGXVuaiR+xvLDOkDc6Fnj+eqtLcH7iMID2X
KQSCAsAfibPKpKqyUvkasHpgouR9T1Pvzf9+9JzjYkZAA7gxfCzKtGJqCy8Yz28I
WEUUPlNAZ/J4Z3sTjiTaeGCzk4Yu8Ce0pnpdcVOGKV612IZ7NasoHl10EVe2SifG
7kcSbt13NskMQ9SpY4yEyR2XDDAo6HDTVrrXFmGNsoKRHGulyOiYo/XvHbfetcID
dN5qZp+7gQd3cOngauwevcSROnbptzQyImEdcqyOPKxWoWfw72BrgBG8SFXOp7E8
NPasg99IW5383LMXIGWPVgkVyOplKU4oqy2ULoZRc6it39i4ilkzcAQUMSo5Hf1w
9t0NdZfEdWBAX+NunYx90gKAfKbO02Wvw6m0yUQDdQ6g9hOXZJYiqAWzC4lX+R2Y
4nfcAODRS4dE1Gzl/f1YMhorgYOg7BNR0c4bkw0loKDI+qlIlNVS3Yb3RnEdPi8F
sojZmjH0csw2lvwt3zMr7HkskKomPpW+NCZwiMmYR+854AvPLy9fArx7s9cBYwtt
7wBLw9k8oS5Jxizqqtf0GnfkG17looHWV+DRHsTZG7hx2MWrTyN+xXy6N0JD6GSq
bL+WIcH/Cfe3Ui2qx0nO9Pf7eFS2JS7AuuxImzTxxBgMbHqift9oAyOVyl5nZ1O6
6cjmAkshonTUi7d2X5IMgGlel3axGSCxxAZf17aqQAIZWoC4AkBXZW2VaLOb2YRn
VB8xIz4nLzodG9j64DRnL+jpZv5MwbntoE0kV0xeWePeZMNBE9nuDCc16egaZe2N
sPj4b8fwLadVKUuXTMWqi43rGOxJpPvqXBILXggLyMDEjUq8d6UICDao4L40zk05
gXTMHO+hQLqoAc4rJgfR4Z5JwqqJYoWUljcR2TVmoe92QNnVMUq8R8w6pUhWByx/
ZUQF3Ph6sCi9ntmDgCieancrtSEz+JWg7G1QaUp3hSiFagIn0jS+yxK2gmojrfA9
Y+XTg8m/J0astVN0ZOH+mNVIP/UiASQyZirwqzNbZPmc5M6H5JJ+BbCl/NMJenMV
/vm06Icgs73S+xA8RZbJ1ocQUZHZwaLh0r4jmUzheU/F60iGWsWNE+ksRbqr+f6z
9ohvmb8Xhw+iASU/SIHKh0lReQ/yxl3gFs6Iqbj2f3M/JFx0JXXVjOP0F9Mf0y24
C1U1VD+nGf8y6NFfbTz5V8Lw22N90FJcWvGdunAoWy+lOIYUb2SEDHufw/7iVGpQ
FntagueOWniSrnduV6yNCosm+5Sc0LMCweK6EuXci81Hbz/anv1yPluXMBi+YFhI
eWuhTegkK6QWNUeynsX4/TR1NmLeS8xu+8EqDIshLvpklhkLCYI4/i048FGZ480x
1A52FLc2FYnmJUhQQw/k/Ldc5ULFEK+IOYNXU0t9vCmIo4J+ZnfM/DCsjISvogst
DAaTkNr5J1WNMq3hWqFVPo4F1+A4kR+S5/iGdCM1Vq9SGXZxkGgqlk3XlXfzbAaB
fGXsRmOIdGWW8grzTnCLzuguvVxJOgwIk8xbMf2ZTvEsXQDc/OFWT1/OWDB589q4
eeVmFsspv+88DYe8S3VlIhpVp2FUAE8cLPh3kS+wNb4KujnRVYQ/pBgXPK5R4Oae
PIbwgkj4U3J18Io2bGcVu9EyadUbfAvvix0l77we9U7222GlhQsa+F7MdqD3qH/9
FPkMP7anNgxq/HxtjDO2yMSTM1pEtnUz1W3xA2/rjuFvCpz1qhzitIfiiavmTksN
8m3KhGLGftyjc0dIzEwOmrfKG0Dpr8r979jfZ5q5sR8XIijqWX6LMHE/IwMt8Xun
89QMqw6pFv7XHWiKR1OZBg27ycLPOhh+9oaaz402aSGya/ZEvl8QDZIVoCprVN3V
YEAoPe19PDqOmFzgD2C39NWztFkT5dSfdbww6D3Z/HuQ2i5q5ZZdt+4n8DSJciSj
umAfUwvicn4e5uTVSye0xWeyNzsppCnFBbsJ0TVUwsgxMgEm3ULIxrbySIWhqGnL
3lf2EDr0axK20RuSKMdRFMXwR367dRFjZskYdjo4XTjvcFSecUTyHIVXooF7IYC3
2Ft1vM0ENpKaUt1M4JYkEZd0e/uudf9r28iAiLDtBwml+3+blQGsqj7Lm8wWIVSm
9G48hCZtrNUE+J56e2Q9aekQPfm0GePwPDNHdIvNqhI=
`protect END_PROTECTED
