`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sPemYTTU4Tyx3tEt7WSjcjcA2KIXHy8BDukgN8bz/LvY3MMkrM8ji+8cPTi/o8rL
kr6Ji+1K8+ybU1fhx5xHcZDHfDjHfw/hisiylZXQ3CnI+zVWs5y9JuV2YzMMfrst
UhnQq1Y1vwikVKMNEz3Vdj0cODLahrkCG0pTgSW0dIzV4n8VFhV/G51QbuvbAka0
GL+h5tOxbUMnJpD69DJvu2dMG5fAWO/w4f1+nNoYx1cQz8nzLJ4px5r4eikB2cTQ
HM9jF/vnovpYNRvzds22IxlBWVZ4OVR75uWDDmzJ+g6IoaMHb5Rt8vycT5T9Hvv8
eLv7M266DvC6LmgVvleLF50wNL2XpkdxpSxzcdAI4jav6C8NJ3Ko37VQCPFu8yqm
9oJHG2v880W1TBW3WxU8phcuqE4OLYAht1ACKsVm40aV6rtCqzdvmicUdQ66msvi
pRL8U4Fdp0VYLsO3dWtS9TYCLcbBplL/zd9/k6q18eL5hTLU8HqolNUcs99pyu6B
/secNORGbhJrAzEReWZJ6GUYYadwU3fZiNofRBYgJTwUPACxW+5NgUk56jx+3YcF
XJi1VCcq3IT/SawPgpnT4jaWY9SLFMwiizq4zPvV6RaFu+V0T5a/EHyWOS2ZKjo3
+aoT5jOjT4PbJD50vgahwLg43mgLh2xAsVlWARl1G4CVaSyaGsczfU5s50ZSRU6j
YHaIM3mgmXwYNxUfVXMzFI6KoT0aFkUfatSaxQoH/NsAg7kB1I2lJFA0GmP1Low7
HpwmJEiCuIBVr6z9DTz2t4d3RFn1JCpxqUoOzePM/AJChMrcbG44Li3huvzRO2Ls
glfPstvGHQOcqYltru5MsaCuUJUKFnpQs/udupfarAs53w6ZAMY54B9LqOL++iRy
bDESVlePKjw6oHnqcglVRA7I+MD77t55x0Mk3+IX/A3v1vA4lJ9Rl6qxB4GqgvJj
dV5zG6ZCINL4HHbM6gC3XSL3LHDrWrXmM5hEO8fLHSiInkOkueRxislxahNRCWVr
QOfBgquCvX4h+8MhItW4UOo56vCT0XCyplybWuoYFO4=
`protect END_PROTECTED
