`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1MsKxmwHMFfhEiTKtY/XJx10oyiVjICcfFCmEllARFl9wo8Lp61lVX9oX64uGnP
5YRVBnGHxLiRAovflkTIC+nwQdcpfW0YsDp61Cs3YQAZFoZAskht5ype8d2R8QXo
133F2hHPzYwohnnebXfTx0xnPmE3u8mzuL7nUQuhgsQDQ8tJg4KQZD9uvjzNRwA7
ncxV8lFW62KZhATVnuF4QJTNo8m2M/vfezySL0RSJKGBrDl4E7lJ2yzHS7fwdm+K
jt97c+NGtcnCgpKGynFPbbTfKiKcuq224ai6XvO2WPXEv2lMVq46zwG+05iflb6+
HY7Iuso1wXaPEVNCW+TtOZZGKyz0Su29NYOixfiBR+qgpQYZu0TYlGU5T5l5SYqi
K3Ey3mM6H2nbMNTqObJRfmX2DG+GNi8n3QPXGN6SjgpiTECDNIQMV149m7UPzQOq
QduXEwctpZsRkBfxQX1nJXe9S5Fnr1WbLVpn9IEgHoU/e1wvmliHimeoRRFfhGuA
HQbiV4DHXjvs6YuqsiQaWP4TC8ZLF99n6Kt54DDuIHJoRwVUQlwCKuCP1KkCLWta
9nC5VDpK30vaPLZ+es1JmBzX/BCCmVRBWmF4w6tnKEBfX6AVkOh23aXVH6jUolKp
bUUs3JRL72zEmOImMCtdu7UF66gsOIOV6M5YcZbj4OtIIKceW1GobmN3cK7mGWNz
gMFeurK7ISyBWY5c4KwoI3YC90H+/UN5N8cqmWSJNKiApqCTCCfhE8m+Fyb3zcBK
L06KqdLEr+gk5If0UFc8AmuE/s1h/5iTOlK5chwUh9e88hidWNETPTQr1JQIh8hQ
JZvm6y66zSQuU2cKhhARVTT6H9y6MbJQAxKWdQmekWHdC5qJvWwgKXKVI9ezzQQB
TxdfBYGg9DcRHFpSnYZEu0IXL+OQUuqa4G73xlvlrdEE1x9l9BrSDsMNGV5kt4h4
VeJ0hLWSH0s00o+W1K5e3dROIHKMkbiQlrk4BtTT56XClJ26SyKF7ipSSjO4NJFF
5NJcsWtFhG4GYAjQTqaFnJZIMcq58zo+G7/1RmAq8pU6SlTQN4koDgZU93X9AGLU
6bAa/kr+nOXPFCV9NdNm0jPrCUNByYC8DlcbSxRayPxZhUbZBmew/xjg9bqpL6lw
HeX1mQ+q/cty2K/W0LfNGjqtruAJNqyvrVcppkiazHjejD0vOuO2H41NrKMMYHsP
m8togJAUO9W8rJdK5MQXizUHiLUUgsTSc/aw+vQ3pr9Au2X3AM8csiOwF25iLdH8
l5T1KFuLP4fxlfiy/FFKTphS/bh9MXW19c3qBZXK/Hjif8TOuxBmD+0zcf2WquBy
gTnNhfblqbOXRXvjkeVbA/HsygPhuFnyqrS5csn9bI4fW/c+3FZ60H3vO89fTS9O
/U66zz0lsw4SlfW2L+LOgwd9hL1mx5dyzB+BBRwvkDv1ZIroZO7Hj3ow94ZtBbE5
tah/5IRCkWlWPJqV+LYKhrzjcCV0p3JTZNLiWib2iY2a8jzsMj3KKJgscNKTYWe9
I6hsmdydfXHGdWnu6Nutfa1NK8ShYUrozfv0ArqTjvVonHiLITosDPvj3J0hGbb8
uxdjOfVAGEK5NKGCtgrlqFJ6kxehFI7Jtl0XWsOUfTFCsqflHsN1AKOx784rXzfA
4xoFWW6BZ4pBruWw/CF/aGyjrnZ6Dz8P1OdWuSqS5xY/7zPnGoa/45Z6s784qng0
DAKTjZ2y75dzHoz4798e8lP3DWS3n6fDaX8GHKnMPErBL4zDROlKwHZp6m2NE+Ya
XCv5NO+8gbXelcRP+6DTYF5vwJt5EW3IOc3G1JvIGkvyFXD3d98RLbMRwb2wu/sg
mUqo8z9fo4n171VqfkavG9kmjljyZ1gz3pJXXt/00YkJ68E/uP1miHXxZLCzDnpg
AjFlHFPnnQ9LoonnOW+c2z1XBymlPb1Gt/bsE0gR3DqHXNQRo1HX0neuBM9DwDWD
pQ1aXA80901vtUvOtbEVgnFeAgXO7gcOlDVZf47BKGqullUdCN9qVhFCdmylb7OA
t2f2OfdCnrEo4HFbnNiTHN4T7sPJP/c9e839uyDZ05ioTdVDWb3nKehewFLwMMtQ
4H5XOmPBL246Wk7aknU1e0z129Cw74RYs1KvPRlke4hsYgOELjPrGzn8r8TpDGJV
yDke2X/43oCenxh0SAmEINT92LdVDN7SPrtcBLT7u5VOtso6Nulh3UAPSbvPBrC9
xkDNaUQ5lsdcAF6UI0YFi/PzjmPEUxLULv9NxX+znzaJWRv7FJGEPFiPsGjDsE2E
tk7cXFjMZVjyRUgn5HlZ7gjVUkR8zXvb0PkqOM1kgPrsVYvvv3g0CyyvIuzALsm+
vDSrQL30owOU4Y0O3Akh2non0ImBenTuptkF45OibJBMuXFLCE/11YZSLPAasE+3
m30xV3Yx7RRQAATxBCKw16XZF0og3dzZVYKwVEfCJHGH9IRGvz3Kt+5zqPZsaB6N
B2UH8IiCfzGOhptiMYo516iKqlJJ8syZFm0yAcvAaQCdiI39cr0Cbyc/cAh58pF1
qa5vA5eeGUDHS+HOaMGvaPMNqFTfI8pA+NKJwQofp6Kc0k8wXWYwR6SLxWfzT34d
vqEEascOQswgPvefXLbF0bQSixHxAu7zIP2qKTqogMeUx9uUMQyK5t/AdTj4KhLY
LRWbjE5s0SLc44pRJk7F9LhDsrEki5ay1Y2NlTetw7p102PsnK+i2K2+51Q6c0ep
AqL1HFlUBBHNQAbTRjqDcpWTY40koY3mmW6yYNUKvcXMrCAxlCaruSYpPz+Eomov
bPmIeSyQ08VWjVDByZV92hYroAvfp4WS+s5ppGWNJWKmhlZYEQGkfr4W0URElKVp
rPdTS1rAtJ8vAxwzB6ac8FeOK6RfefITqJpwQL5RoLRelMozwUnmszeEYQ1bZoan
ZMWWhiPor6oDBcGuqrWqfppOqRoep5jskBohDsTmBJoPwRbKjrXATb8fdU6+Up/L
EDdGA1AYoCLItmKZY/ic63f/OxGBj+NOoE0kKqIFK4HaOfjw1yiP3WvvZtWWNtms
ihOEh7QpryP9ILQwODlq+Tdt433kELs2H8xucwC4H81VMVQyYGsWp43N5f1k47UD
ul//BpiYjsydtk/k7dfoJX4vGAiBfU3j+mbWT6ZdDCwJ+KwlWL58G+ab1P1ogISV
tDuk7ffP665k5MavVnKSIROnVA57141fLLIEND1cOOoQTAgLV+naSqrX5Sel1Ntg
GkGmQ1DGRSDcuVfNk83tbIm5KoovZFY2DIrl/LiG3/y1w4c66B7nyTre01cwzWQy
x9RaicomiAkv62LVOIOibxJyvoHazQnj8vrZV8ByU4yEeG3Z3IUuzT/ApLYYoi1l
KlDt2MlHj6cp88WEtjcY6iBtkamaZojjGFnpWpJVpKrEpYzsQlXStogk8mUKDv4G
TM7tyznaCvmisTs7DAOeFlCCmsarpuJaYKJYxW0ZnWxldiSvHtEE1hvlzU2AfC8j
PuouxhxuWYWufqUJs63nps6PSD7xII9X9tnDOQ+tfF4oow3KFD8W5BJfS5uL2Gqr
GeVy+FdlDKw1RCGVTAOr7V5R+hXZCnQUDWJVQksRzfpWvxptUyWEKYC6Vsi9Zvtz
dkILI0Cke+fj45XA2Ui1CScE4GF6y2AZi+wc0deqgL2GTVpPcSt3jF6iu1VZYgX/
aR0wpn+GSyIpyfAlInyl32ibIX5LIueaXvz8S78ONjk/6DHmLyGXBEdkCYikIgMd
kGxOLzv67RHYTNvfbQ/5tqntrD1nxxYGxsie1EuGiQ8GU8ve7KkPhC0/nOVgLr08
EvDIuUv94qXCzBfj7P1Kf1+FX8NdVtnDCdRaEy/+blPBCsh8hFJHrVi7n+z76usG
Jd2lWxa4VmSkDwJFOXJKl77CQQCP2A9ayBJR98ZS3zL+Tw6jT09kBAHyaRObNzhq
xnSZcBRngPNi8Syh7TJJb0hVB8YhH2lEG6GDezZ3WaYKUXBNHwdjnbPEdhqENj2V
QCZPpKWg4ule+rPSFWvFyxSCDbI6EIS9ULO66d4FtpOc8NLimAp1c5KSw1+UZdFC
Y9MPYs53UWHznUf7i7njWwmQZN8RaK4wOP86xXeOTLZRlXhwvuJAbhyT2IJqGg4Y
wM75BswRvd0/7ggE9CS0lCSebZCEtApXjRx7DtZ5GodL8f6EvzofiVNTR92H2j2s
U+ifmUzuoFPk5714JYQEmLMBFv1RziAv5Rak5Mn78OFuPoAJBCbUhILd55jg7r3z
nj7wGDKXiYpVgI9KxzysBbXBJ1YYt/zAVLXcNcqHRyJn4Fqz2HEaONnx6s2uYyDg
2AAJTjqrJwxQXcNUhckU+QIrXukuLAhIIJZUH+ieRk0xIRgMVTZvh1E5OxCSDx45
ba2yp3WcxGUNyPbODBwdID/65pTy5kcWRa9Ar7vdnm0M3PfIaES8X8YdQN49My+0
E1UxfbmunoYzij1h2CsXnSM4o1rj5WSzVg1D9zmst8+FtsGMPLNy2B/gzOsk8wCd
FjZoBLQ2u8US171v+NitWAXUIwGfWMXl5PuZZW2vyacBKvbP7GY+Tm+0AW1UnHnS
aCM/zU4UOg1L1g/KBh3JTX8F1CUEtZuHFWQM/kfr+2uKIkZ3ML3FTYVNkbM0BO65
oYPSLYl+D8Zu147SLV8jkUUd3BeIudPSoHMKKPTQyNPaovhhX8Hv4bY2A8MBbMi+
nAGeNiP2ZUob0NgkKZ66QbMc9Axz+qSfQ1KMsY8OIUbhAvYSfncrXmrr7AvN0cUp
Yv9W8p6f2VJiUKcPK0awDSQfUKxjyfdYZKpmkbZveadK9iO2Ax3+kueMumumbKgS
PCUJZmyMbGdVmCqrSBpKrp9VCWCccRImGrjz1AWAPOpaCKz0PUxiROFKdUJxDD5I
ed7g49MocUMtxA4MQNFaXmjUmh62x8gwd03OzAQ5VWe5unZkObKyUr0fC//AzQ1n
OKdQNqL66WN+QksdlgUnPdxOQbbkqaW6ECmX4OvFJ6xPkCr2qsdNMORnq+rBxdpP
ZGgLaOuZWz6f6rVJ2/ND4Q2rmHvHjPjb8L7PI+A65nvAEkpqXEBxIWKV140VIV3B
wLFZEhDtAp9lOXUdGCJVrSW9LB4uaEAM3yk2C4jurTO+rNkl0xpkCSLIbf5s+ume
JvpGAqv2ztc9l3pLIpcgnFA1qpLhf7VNDr6sWT+DCBI+viZTcwgNIwSojLrnSH1d
c4DVumJ/vo144A9tCLnZVSrbiSgdd9a9EXunfN8UG5sUlAg9lVpHZ/ZIMoGeZmrF
ZSQRy+cDZv9dZ5evykVqOcnNld3eMLE5QUWKW9sEx+HEt1YYUSbvq9KW1/tiPda4
lLpcTpvx3MbgIWSbelEwMkdBp3rp50OzXFq59V8tb2zVyckiEavrawRXCmLGKfvg
Q+70JrdTIOxLQrKb3HL5050BfHgkKt3b7Leu3X94nthPZZ09BxB2Db3caUHZdZA4
nzlsqFx112Oy5Lq0eVcYZqGTcBVTNr/V7mjodoI2eRG9w9kguR3OYrhuaz9QPd0B
uaBupKPAlrA7wu1FVETKtibOt8Hv8KRYllTQjoMOV2esRhNKxH3XBvS7NOWRIZTC
+WxI5VcBy3eIFqAEKKZJpEmRKdsmCHtQ4MrZkt/8PI6oRlnMA6X6dQL52uJImj4k
pQ7QDjGdStjQlYquRbeOlQMltzI65dKmam+CHXujomitNB4ZZCwXrB6GTCYCgQlh
9uBccUgwHgiGIJRKEGDvfF0Xd4s+88JIg5pPp/lJYRakw3CtLH+eGbob+Dy+bZTD
YslEgZJ3aCnOZkpPrZG2BWJCn0lbYdSTIuB1JMjDNOsuWUir34iSHRzN1nexewN9
zxy8pPSN6/KZdEQWpejFtVlhGUhOzXeVW72ArBloHcE=
`protect END_PROTECTED
