`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+htGpnD/aMFuCgLMvR5vJtSQbsGgXAQzgEjuUT72az/+hoVl4XQyouwLvdlPvoR7
dC0WzeHLlqcsMAp52LA9q1azuRWUNcd6fjQO3Jtzsgo6t85H2DmuHrOK++0nMjJ7
opy1765vlCu1M3UsHRVzd7lRqJ/3IsrrhsqZquDE/paGF+0U79zrVXkf2WmXwk1g
TkBN/4P2nPKEBF4trRVmd7I+vLjFTkARCy984iZ8bLu01ribF/5XzP/ab3A6KGXl
gymQJoA4EfmVPVZs9/3elklz0YhR6l5kxEc/OTSdnU5ppJSFUQaBcYxd1OqfiK8T
JtGXk/SBHaE278uwfx0SUEMH2JEgRSy/vXVKt3EEAtvgdlsK6P0Kz9qIwjWu8vhW
f4i+87N9g580NHmgTB1YZ83G3RfMgRRavdvXyp54xRxfcc7aZu8bP0EVsw9bTRtH
fdnbl/oh60z5QkhpclTIdg8Q0mVWMWA6XtV9BVs3/eIUTEtmeK1orr3INaIKmwPl
GZGPlofKRcFPcGjGAFjrBNKM+rPUK0s7kAH+U2VzyJzKwzpwWMmb9PGczWIHoxap
mWbr35uCbIyVGhrOyhlDDoxO/6pwOiEa9b3vEHyZO2cbijM6gtMwxG9qS5Ol+Ulv
8YSgwxPTLc19Ml09J1RQqjDjp8l2ynBSdZcOCRgFZrdaTMGBtMj8PUhzpf8YEQc8
C4VuTsNdMxeh/bHY5Fh8G/UpbvdY67uT9kGgdLPV8BRqT/t/+KET1j4VNMYQZGTf
Rfu7LyeCnQG7dRO8bckZV5hfKmLKxePy9JDz/VdONMce0kimfuwwwMjgHXCRWlsE
u04Tzcn/+bDjru1ZTo34N5W7jHknhkDgg/FnpWqJ1HMaDq70ZxTqdrl6JJInvXJn
Lqb+FwN9RPzWmEnrhPpDWxaVZbc6+ucDQAGTQKGIQ5MTbjw3O9Jn2eN5yfSeGFWu
ztNYLsapL01/yy/ve4XQjXnHiyKbs7uj4YGZubHtkTRuJ1YuGp96fsobNXceCB8k
XyPNvpYavxjuuUwWKZtrLfsLuXBL/eZx9pbOWSenosY8N6EFlRxOOU/g6yCcGM2a
9krNKNLJtwZZCVL1KVQ1JK+9rqTheDlA8ZAbGrLTp8uDjYy1lnZTx33f0dkilPQQ
`protect END_PROTECTED
