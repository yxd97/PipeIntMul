`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vgPWDnQrwgVpjI+w3xG51uDN/lcRG+xxAZlFkwlwlSj4SBw6IqO6YAiQltZHhQvy
QmdvDtRdcpe9beXkPK8d/naWngJGlEJFHfcurZtW2GslQUE4NVRZp5AJsfI22E4b
4Ipyy9CKXxaMuZaMsY64f9Z6LQiAJHuyPmD0POMl51qIH+JewErK1RFm/1/jGDXW
jWr4eJF+JDtVIQGIM3+cxyOYFTMouRocILNMxooLHQrs3h/UzX6K8epQaGg1Yv2p
0EvMamRVDTCEMo1RzSyNPqC1+y8+Uf848c7H4mAmXPF8Wk6rBOj1tFpe4IKRNv5e
2nMhqWt58v0+h+BmbFq9Af4HcIAzcWlepI4SiyAFNX+G0aq5NjaXcF3gGSheeIxV
+8RwkI2k+aA3aSlhHLUyoQ==
`protect END_PROTECTED
