`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sp/y0saaQgBpBK1wVsrVVpqo0TYvr/qfWpunWz5c3orMNwQHAFmP3RetNeNyMEsx
vpY4WbciSABq0kwSLQXMkZXtt844RQkkjIWW1p0iHOCnrBPPROTS49EZGxojOwZl
JdzP733PpNyQDZRKkvIqRQqEpI6ESL8sdWeJrsOXbFVYn/3Gqn2gZnW4OGeM4pny
ONcli60E7t6ruZ/i0scDCAJ71XO2kcK6OKm0oFhyivIq4y1FzCaj2Y4x3ECJN5Dv
FlrS74BFvZsgLU2zPP3Ak1pzxbTWUVo5qwQNtF/bwH4WDxHcR9xnYqrznIGToyxF
atQP3bpkmkzzdSdnV0lFQyO8L738t1cLQhuSTKhklBX+MD2Ng0hd8SYM/Y1Q8m8w
NFeS7rM2/DI6FTXKLXftyu4lq+gqDWc/U7um9QZgTcBKe99ZZzxzeMNl357RoCbH
0zE7mQX8Cx7Y7+KQEGrCjpyHsOIRWuztWXZyXUTq8nzbIdjpk7UhtY/tTSg3YFhZ
UOc/Vj9SpPjSTXBXixjwhiacTzeCzvFC60W98HlNQW3hTsNWdjPAGaqYrE7hYx/S
ixy6Bjhdt1K+lSvNzZC0Jhow90E6kG1NSFkNF0vYr8+vz6tlQisTqozk4rgXdgYO
xkY2Ed4UzbpLpbP3jpxDHGSbGhCW3xUIDi19V14phujvYp3ce801nvf9vJ5j6cFM
ZcTYbik+fZEc5V6HcWMeIw==
`protect END_PROTECTED
