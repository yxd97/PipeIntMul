`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DEUR8T7X4/F9BP6inZORmdWfJaCgjkOISFKzb9pucsphPPi0uMscwXEmo8D+C6DG
D2ZNEpEKrxakdc7oI55otKjKde+M6XCZAetryJsejvlvUCz0p3JPXcHEJNoNKz27
6jIejloI8nniJD4geWX5bbM6kkrgisPTCMkiHertIXJWtcnv5TGfn+kHlr6Vk4l0
8dioAi6Bnphqi7we1eE4OpdTPoTcvjjWqfviYRBtUO/1YYQXWcpnwJL6/MMgy92z
6W+AqDvyM8xguAiYKmQHVnE8hi5kx2Q0inbjsIqpu5DQFjp04PACQVkWokZKo3lX
UBHMizr5Ei1HeeUFWD8+EYAeqClahihOi7N1kMT3XyhE98GWcPPkjSos93vdVYcQ
5YoZZhEVupewE73Y+7xUKFnVmIqBpXV4yxBotX2EhmEZRhmcWPpdUZTSqtW0uZJI
rY2+BbEHqTm+TUZcR7QZlFGl4OtgNTTMBCxfFSgwnGyMAt0wqXhq9WpRNTvLCpT2
xctOb+cCMJPTb+h1qUandz2vIcQpY6pxC0e+XZ20BYqK5NbpUiTPyNdvdjdGfB0P
`protect END_PROTECTED
