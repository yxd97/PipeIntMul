`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMeVknNAZ7lxeRPybIABdJRPHoHg92PijeXDoFYQAqboo0l0chPF0TX4gzKNXHrJ
e0oPTSP61aiuztjEA0ndFWcn+JJExaUbUCxJV9nkjOfp02ZNU8HRGOPQNEMShJfg
+uKFQsI1hfQY4lORKSnt8wzS/GSTNQYbgC/4SBBWxavBb4Zr9Aod8TyWzrr778mm
GzbWhtwdqEcKy3tcDj2hCCcNF2GdAVGU0aNZPTh58Rp9ZbVZlP4ADtkD0n3tS5LN
2D5IpWL/Hb2FqZ0vd4HnC7iTLiQXgMgdbW8zTstjZo4in46Qe/DL3qDNrXY7kKDQ
IdT0bkCtWepLn+U/hEqbfiomA+nARUs6xDnF6wz/WVw=
`protect END_PROTECTED
