`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RrHotE3Ywo/eY1NNqOxsQSosAVotUZJsiYsmSspC/7FO4CkFgMAAisgtWH1GXduY
xOVtapOzJcqJiWVk5fAKgShLXO8cIbPBL8fKMnzTjYUyFv2R3KpmFMGag9d4MNeM
qTpbwnJehG/CDHF7/fF4TF+a/lQa/JQL4MCyxYH20LdQoH3A7egkfHY6jFpy5HhS
TaP4Ut8Zg3gSoR+ohWOH22CfmWsdcmCjbxjpJWTcvYkdITYlGJjNqhJ21Qz649HU
bZsjO/2w4aBqgiTt60Sh9RHZGG+0UroTdV/9bsDgV4k5T4CYvdBmunzGRq7grJAI
VJw1wDozYmwxwXmwrOgFwi7BMlAR4Xu728pUduVbO4CIAyBGstXP7O5tIoP/4iFx
lw13KG8vDy1TyuNjp/1z5pgS5SC+H+DjMeyy0N+7DLCcKFz0gp2gaZq8+/efr2bP
icN+5f+UK3WqTinCM6uGl34wGHOSjY0WOTOR83NcObJEk+1oooPWFgjLFz5Sj2Yd
u+fjbd//fnW0wNQYnWUzQk0bdkjz1lYUW7cxf1vrZ+ip202hvY4XmyI185Xl3t7Q
5BofWIzKlK5lulkKzjdF4TKAGVGkwYfyQ/fOHTzs3AWJFSefWiPN3zO2ohtG9vEv
R7rUeh7HiMSyYKl7A4UnOJhJ4d4rKE10yaoFvZm85WbKVQ31ACLKLInwyZU3C1x5
5CZGltlhC9bYAyAQ7do5aXb2np+pFiWSVgFHh5rQIsHtpaCAb4X5XLDZZM9g21KX
LyCaanqiK4GVDGNXy4JhEhpQYmeVT+N1iIZbmlMmZkkIzMEnlO8tcYVaO+5kqX6G
cxdgTjFDcCH0tJLzTwqASxjy2yslDyXF5d7Isx7kr5xvRxCvAajjLsMhuGP4ciId
IXumerEURdlEpixSkvNN5b8azKcp1XwtqDYmMWtJps8RqTu0VKn3dFw1KtrmJI8+
AMzftsZrm8rxbrcBnqkIO0UwVIs0IQihQ8cmv9pTSRhs+btRnwV/vu95N3xUtwSC
SXDOY7ZB3U4qIzcthtUh8gRGh+TYtOBT6/nBM9RU3qYJd10cGKIyftAUsU6ew4qQ
Wc6r60OsX+4TcKTUoGcfE5EgWvW+L31TZKLP/7p/hJ1dxxUK4I0FPPnTmZ81Hbmp
PZebA2Lk9QKPRhisTNC3lhhkRVlVLPVDXLZf6Ac5NLMI9H7D1143AV/R7da8LUiZ
Q4NvMVIBAxRNH0nm5hbVHBF4igIRtjZ+OsC9XL5Pz1ini9J7oMEek/4zh1HuXPty
wq3HuD/Oq3JIouZ7LcXtNCUzWMBdsOJQwuvXqX7E8bWqNMhRunRpnsThnXu/7+6+
5kctlnd4lsf/zPmQ4uRZ0q1Nz8cJE4P7+6K23Ue7mvLnoUYXrUfxrB05o9FQ0oI/
7jBRF5EVo8ATPQokRuCNS6c/na8oUUNUfIVJAnlmRK1xK9zq57PzT6+XsprVOs8N
+VSa4ySAUD4A2PtjgY4MryKK54zHYpTXmSqCRpelVu2fEasFw/vcZSVFSZ4raa9v
ilnJ3ae2VAY6zP/GJw2GIwOL8NumQHtfJbiA8yzBLIfatiRo8dPr1LAqsH3RbROl
uuz5Tnq1U0LkdwlVi17mNSbErIoUrec/DDNnr+dQvq8CWfb3P+4WfUNiePRjbS8R
NiBj+7ORi5zBSJ1ZKwfvj2yeWTVTe8CEKPHXIwMgIYicfT7H6I/36pvmRQOlPv7E
2AkS1nTDQFfT1eobJDao9lfAMjotraTyWL8eEkQXJy13U884yRVMv2eOMt9lHELg
kWOxzjuF/iBxIN4qnNBE1Ypd3m21W0gT/ww45bVferO/X6S4jpvKDuqwaxwUzpip
7plCch0gHeXFlyMHZdoO/NSWLNHPiHVTjyi1w0tGAB1VwEfCyXZXilZwBbiMo5gh
M6jOwSiuotkZK6QmXo8EPU54iabofHxIjSY8rb/eBI4GTrEll6z56yqZLE6tIFfU
RgJjKPWhmsRnUc+TJPdWbjYD1xsfFa53Y9O/sPcRP5jMbCK+ZGc4ANdD9igUfKrE
ON898QgmLHU5yodI7h/WRrzykgl0/BOSC88XDUH5JPzAOLdghfOWt4QUZqSgbcOv
CdgUhZ+FwLFZbwjb2moHt9H1WbgypFMDa2lUySj3DOtvheYQnGkjuPZR3mWU+2+n
X7JoakOAkGBboPbQSrJ3bKAMWd5AFp+nTE8ntR0qE6ZC1rWGtKoaXTzBA4zVCAAq
ME9Z2HipmNtm3b1Vhe4AUDIWs7WaFwyyXxBW8bWX4C34BTjmk+gA0CHV1qgaxnnp
HJyVNrRSzqrH1MhZnChbB6mNlHjfql1iwwbdV8EwJyC9EZEumVlkUN/lkeE00NDF
JPnU6ZrOTf5eo0YDm7/9otpMypAbd/+TpJ/W1eita4sGSR+jzzf78Vf4EZeakJHU
JuLkdt3s7Sd16QW+fscx6A==
`protect END_PROTECTED
