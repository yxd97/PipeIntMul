`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAJEMydmxaaqvdv2Nlp6apCLHL/DcSN8vZSSAdYHyTaaxTVPvgmWF6SA1fQSDv6C
ma1j9j5mLIUcigF41Gzf0YexNKOKuEfCSwQ9resd4xQc38lNxY5WOsvx/GDzVDyn
envTMeL39WWjOP+b3SzVVvAv7IelsvMZjyuA7xTOlxyZeq3np1WTUWDOTakCDPsF
mk6dOsVRYDbKrVo7wiZ6ZcJtUm9wzRL8ZuALorDk9HvTi9r/uh6OX1za5FlK4zeo
kukovbKmNlvKfwSbHLtKKKdTPcLLHUe7GfB4jjZz2BhsbKX8SIf1Z0XVqoiV4wT7
Sh5vvo0fwLN8vaD0QIu8RIB1Yle6BA3mpBj+G5B0lYHUbZZRx/jE7axYxG4izNUG
UuGKw8ODMnh/T3BQlB1nl4JGw7S6sY9wT9woBLykbfNVpMb0dg/MIrmTaolCNbvv
/KFyfhO2hgu00vNXHnp6MgGQbjYT0hjhGZMyKBAqdAVQuv6VBktauXo2sQ3icO4C
`protect END_PROTECTED
