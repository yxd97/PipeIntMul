`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzHOo2IRp7RYBKDhLGaXM2xFOj1TWdnLr92CdRjaHBwKw40aqME+gJ0Hd7ZtS/vm
gmAUqFHX2uRa3OMo4oTFEuhpQlw4iVFGxGggiCmSPS+prDZziJdXBwHDjjMpKTF9
ded9cuoy+ze+nc/9DGRNQZpFlFLGNpSbGV8onMWlvLKfbfZBxfLufBCRbq9j0xCT
ZjMRh3gfx3JYYaliRCR2ZDI2Bu71DF2r45+bl2EMFnTCxCquomveKjL5IkWl5a+N
xgD+zHlXoNxsjurLONMSmE34/Fs7DRc1gwpjbMuA95WACfixb4UhFXwTbwFHvj8f
nH1GGakyBrqTmrYqJFpnqWil5SPS45IhltSV5FDAjFpP2h7OpAJR5dNvi/4LbyIy
2ykjW3+xfpbV4G/a+IRBJg+vaxjD23lIfsGJanWuON4=
`protect END_PROTECTED
