`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHkrH2IFCsv916HD/fpvOZRPf+s8u2n9szM/VHNlO22yCh+AyttNb41/gNqdWKx3
JfNiqE0uniNfeC002B0GRFNrHRax0fTXO8hhpPkMYTlAyJz/u1L9N2bCtf1yP7V2
mhgWzkIJPTDFrteIyRc4+jds4A7dBY+X7sTdRhtKFWigzt+LhhftZvHztkcAa4hl
Wk3y+XHgYNt3ODukk8vxX6WYaHiuA3TE9mx9vj6BZPXSzCgXyu3zDaV3myye5YKY
wYJ8fUMZAwVvBsn/o4Y2gKE79QIDt16qQ5tBkwEbxH8wJmaENGXJQ5Z84W+22+Ir
EI8D6qUE+Y4adkcyX6Feyt5mE+LZAJSRggXGKhG3iXLOitLsLAso5gap3IKSIXkG
+SJkw6n8Bds9vdH6WZX5FE6JT7fJL08KQR/6i6OHMeAP4n/udBQ065mGXXaMWAt7
jFcyeL3fPHMrILVMm+RD4w==
`protect END_PROTECTED
