`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JuZ34972bDiRQqkpvWSoDccXAWMKz4DIOS/CkbxCl6WMbufiDbi5CJR0YbiGJiVc
Ko0VCtM+DBPsFKwvzo/bLKttbevB6ULsnsX49RAvoGEG6VP02wo4yqUPF7bdWIAh
4XO+7i3kP5EVTUNnpWZG+wfWi2by0wDjoAHgHHnL+DWWiPOy/M+Ika7MKQwhu9rx
1trFcf4XmcdKU7SAQRjKjAeIFtkSNO5pDMFaUbHKJrclkicjkp3ZIdM1n+f5kZnr
e/r8p4XJdxVJrVHXtsPeuZcVpCuQOkIkO1EJ6KLzH64+OB12uEMhVRKWacS5+hm0
xJ2pOo7HY9dqIbYnrTLYwJiQSrP3csjx4VsdU96t9kicuJ6OatGTNF0d0EOlwMnf
Hv5DqCpogdLC4MW5psDr4NSZEOEpMKR0egRRd/uap2514vtfrAKaZ3pYfnuFj943
jLcDWZjZJKvDyt9lsGgEH40+0olQBBVZRCR3aDCPLrbwLIoJvujp1xGrlqqgvsM3
dFH6LHw8j2TiI493wpNCUs6AAWNpmEf6VOmo3mie5uOCpd1K96EP4dRXuAEDqiP4
ZxpYP6cjE4U1isP0i4/lFLlFwHbzN7ioHRLJ6l46UkGVl5bS4cEIe1p28u66RaOk
0ee/MPbtDHgfEq3sKnYAOdSai2IJgZnDk8rRPgYwKMdFSaUnvwU1MmOAX38fkQxk
Ox7fbUb1py3+ok7wg6kuLnBBrtbE7nhE0IOB+cTtGzQVyDsy4FOffmU2vo1Meq+H
NrsRKsR8wQSBmsRqERFlHqBDh+rG0ElNJlG3SHn3x0dHkk3ozL7fTcBeIo5tZ5Fk
hKEb2XOPY+2gbyy9GouvmE2HFuSlddoQXCNgesrCaCEFNlm6a58xPEDM5Mj/C1ym
wmw1GI5xwNtVNP4XmM0h0zYRp/n6T/25VPOHR0KELXAQcm6xRdwJIn+X79xF6E9L
hlLirIq8tctG4gdPKDPAOMFcbykdpxHB1NlMsqjIIcSKvctGRKbTtO0uyjN8Cuxk
5vLbOpEJUEmh5ecA8FITuCR6oMpu5h/ivmZ8kAeCU4apgsMUIx3QgKaTq22BlNX1
35oJu3kdQ4Tlqyvk7+Jg/w==
`protect END_PROTECTED
