`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kei5y24S+jWyLUx77359KO5njbt2vMfPxi9Uwk/KYdXrBTKympiC7/jdzWRt+6sA
5YJ/4nD6EMsBlkhFTd0I8JNpNY0yoDJOExiTbjIK6PlXbWCPJQrfQyLRUakpnI86
r0quTzmqgyR4wd6uWSqWSFgnYTV2H0mQoaLR6nDRZI0uGCkChJBoN2ir89nAj+jJ
pfYP9GzzHa3BxEIxxxVwwO60k4LC0aAHkWkPBOaUT5FdKz8Rjg4TQD+2V8o43cAf
jg1rqm49QQ+E6IzVsnBc9g==
`protect END_PROTECTED
