`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YJ6bFdJk9Mwd1Aa7pz2jr/ROoGAAHb1+T2qkCi3muMegAZFjuRx9OekVvXvB3NhX
8Be3+buo8yARgdXH6e5fKOw8Znbe/ZNUyymWrOM7LyTTSugjIf7g47yfxMerwI07
VfLIGzSTQCH9o4+8M9d8GS+GiKTCR0XwWU69giu0MuLfbfNM7IMQEG8N+awSoUks
GHCt6fYfmWNIa5cKN/WGgTjep1qNEskjdWU39u2zd8dgfs/kWIlR5MiKQBm4pbxO
tQrY5K6ZyRFZdmYHrD5A/VQvYR8ta7PGEtyRnNs2OeUlYpqHk+YcFEuw4MrXVLwJ
sTYF2PPirMrgq4qnHA4+BveRobuDU9IKNfKdOO50d6/WxlgI+5gUynAO0npGPJYx
Y9L2HaaH0XE7S1Q2bsRdBQYiMYSX+MX/2nqQo3QqUj6UsELGrAGoDBkcRYWmEyPc
0Bl6g2fbm54oRLbNNSeekw==
`protect END_PROTECTED
