`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A7heza+fia2BMcvt2e9QOUdYv6WKe0dtObMcdq/NpZx5pIDfDzVOJlsRAUR0Fb3X
6wKAnGZRbQmohCa3okZ0ALxZS38AgnSwpq+Ey0ZXDiLLTUK4edfc8bJjSjmOcgjf
9mvubdQnQoP+DTa2FjQnV5PN0peXikmZjI4SahSdZikurmn2Axhy7XNt/v7BJZp1
Aw8bO9OiMCucsWFChCzLvj8dD6iTUasqGcil+WX/YShXAtEWfdRJYq22vK+Xbwm6
4zLIPWtx7mDdPbBsOSBknoUn2ff73UJvPKNPomU1hqxm5kwM44SwmvL1kgQhtB66
HaKOZlVM5biGBa3/p01aeVarY1qldPXAceYkgasD7eTiL05z1qn932yRX646WERL
/FDKU3ARoIxtIPOcxYET8bQEONLU96NDUFpv2E+EvYTcQS38S+vnbtvhKuFlHaQ3
dNrJCl9LS98s12tE/dmbdcW2emJ0v21tyfBGo9gFRbNgymQu8BPDkCJ3RJ7fEkED
S8WOSRVpn7WurUZQJXM7Gg==
`protect END_PROTECTED
