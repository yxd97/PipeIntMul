`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IyvnxT1EKa3FMCE5N2422gpCy/g2ws/DkZRLJRZ31zLml7WDTDWtBk/g7rtqCXdY
WnfG6ccIfqOiyETEDQhULCcf2MbzDA+IEYsir3eDsZ2rrhUDD9ee/dfxNrCP5+p2
2nFlPGi5E/0w6AFNLyFR2CSqE8SC+gPrls6R9cnzKbvJk0DrIn7URANPkTpqVR0o
2rfgwBTW+3jl8bGyokIxzESJRIi/8wAyS9APukbx9Q/f9gUZ1a+JQSmM6gokOf32
3vxbQKCPTZenwTLxbKhjelWLkTIy06nHZ7eYQk+a62rcm3sePuDpSrBXpE7y3coa
39anWhDuw1kfZTQCKIGxkERXimDGXx2pgoZvbJzigeJivIBnlyTpcra4hqZvlzPY
ScEgsWADY3sRdj5/0/nsc/hKon3XrqZtaPXBJBruanAFucyEPSxocRGt5i1xCME3
IvoaT6gxnRk6DV5Qmp8oQd4E19xCzgn6LMNkWhZS5Az9R9jG352XcgLCpHzJEbOq
LCrYgUN9WKN3no5W8bUq5vs4y3YbEXdGcajOHgtoCS14a2PiTfguNQN2Y4X/bBj8
4czJdjFpcTuJ/4S3rmuM0ZNZI3+bH9ZoHTwWZmBvzsIbJsiG1Q60kx0eDEKee2U6
3vjemr+2noly3gZfWGeCT22VVuIe/mnwHlKhrWBK6qTyhDqqbBDD53onQ5KYOMoc
ulGYt4B9LlDNSHJ4QhKSUgBxMPZMXP8TdAe+6cbifM1xqFVnsz9CWGRyB5UFiohY
tb++3k0bjCTvQjJk0BFqX6kzoHADR0sGdAoSGCVWid/Ykp4bWlsZ9uUStf0hm2SI
3vhyiwtm69KhDDZHEnFBGx/S+F1u76wtR7D4xs2gPvAqtM9hVs2f60z6xsjMoJ3q
YqK2xluBWwmQxHi9b/NOY0EJlEzINEJ3wbgA/Y0I42qVmduRmrEuQwx2p+F6bfpN
GDoGgOHX46AshZNXBV17xEYkUfaC2ExaG72mZ0lfTpS5H+dO902XSq2WgyhhKUlw
yNfvs8mtdQsRyUHJj3jlVG3ANpUupmTK6X5v3ep/765z4WnD3XxVn1P5NvTqL5bJ
/jGTqb6K1hTIAqE7XZVWbLFrYbCs2RxzNs3WusL2FyahekUQKLaproJ1Xtrrbf0l
9joaFEK6QmHMwfKQde3whergVaF0JZ/k4ZWtBB2QRDk9wezbgdZXLsvi4m9ZsDwS
2D8c5vTFoqsxjslIlPAXiIWWvtXev/KrtTfDipHi/DJNm4Vv4iKWz6wFJoqW3ZQ1
7yh0vmVIK9/QdNVCB6FVULg5O9sGVFhoirIt5vIME+QNo5QmkSMqkPmwwmXl58o0
om+8ixID0pSeGuwcnrKNiGTegIaMFBHKaoNms0hvlND+pOrbVhkVZ7ChMnJHVXea
nXTa9nP3Z2P7uNV01cwBL6k97VJXKWBY+z0oQOQwWm9ddnrVeh38Xjgk1yUL7hNq
4vixe52Mn8CeQKY9hgY+fSNQZkXic5/gJNzbPOxuXKuWxLGTmj89u9ecKkz7jYfm
7mUpaRzoO0KDphK91uCVTwbKGtHNUlZK52ifYkU/B0CToMAY0/FU2uuOzUpPqp1R
iI5fYklcaTYxukI0ZARcfGbgNLmredKxgBxIMDg0PjcT8eFVom0YZqq8QjITxyj7
znD9PULV6DFIvjdGqpy0WWgOKo9e8k4hlCTSnXkVQv8p8lraywNzAKimbQcZz1rk
FvReSGeDaFPgLeZ9tcsUXNjsYmaQxO8nPq/ZUm2yuo+EipEG4+bpEJrFNzApIhKg
1/s5bNoiin2MVC71uwe4j/01krBLITiHn0zPXQqsr79jBcj+rxSeiHQvtU71KVO+
`protect END_PROTECTED
