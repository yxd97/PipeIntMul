`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIAZqGd9HKkqSvQhSFkgi/VAuVhRKefja/pJM/v6yIS0FXz4V48vrLC8IvNZgKcV
zq6/GWPV9OQBPqRBfO2BVOU9CQvJr3GrPMGg2rKnzmIRpVM+K6J3tHRkCUkACwaJ
aYRbF7oCJsEKjg8N7Ui7TaC7vO25w/KN7j5EGi+qEF/LOtyJNTyfl9XE85FnbSY7
qwgRbwwJKyAP+JwfOyCpi9UdnuzqSAgGeEMnI7B3Tj27XMmhKKMjZd8e5Q6GRoU7
5DSUgclvJj25ul1TNo8aughEBL6Lc7Cg4640r43KhdLl1Ccj33Os4r1HZvqEImwE
GXlQ9XB5r4/1DbYFKZCUEUlg9Q5e1mqAMTD6umXuM04v4LEzybhgwBlJlYyCZ2Z4
w6P5xvbWsYTMlW1lkio4HSBh1/Iot/P2yt7yJ5O31XcktqFFedaMlwg+AD7asvrB
Z5Pb/hz817S0mUEPzOacllYvZBhjovKEKsb69pIhTHWXVz7LzMCLvwtCKIueZA0k
R+GzB8mFaZOAsBycQXF9v/IuyZOaSd7VumgygliSE1kK6kIxnUgEc2NNSgudIcG8
I27cUf3jgfapC3sjWUazfmry+2i+BpejjHhG79b94ds3EPwL+jagpTGCyyufvCd4
AZG5n8yEPcBmKDc5VQn99G+VVP6yQyTtZ+jkvBUKQPJoRq/uStKV+plWYJ9Ew1Lq
SeJ4+uy9ZQcjyBf7aL/PNoM6NVpJXHDtZZFvbPwbHwMsBD9jIo6wgPDqp8qYPwq3
`protect END_PROTECTED
