`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oiyD6G3nc4IcmWNV33dAiP45DQF+vKgFPHrzfweSzmGsURDAZCb7jlgBsU1S/Wzq
pzBV3jQr3Zv9MBxYFwL6S/KZQCLq4yNBcNDkH8OEw8BdayYdz43169aKY5HLLOkE
BNhSqDrPakUH5vlOfgNgaQ+Leqc4+P2x4j/uLu5RdfI4c0zbMctwrtKKHJ9xdo+9
wxELitacPghmh//le0n+cmgoXuUXsfcq/bXRO9Zl9+s3wAOZFYD+qn2CGWNtORi/
nUaVWTQOYxKClFZ9Zu8LAUVB2/yv4bw2VcDXLJTep7b0/kErA6ut8kGvKhcs9Y1G
beRuChaob/H8Emph7gaecIW2gHiQfqnT3+V1N89/LdDZMhgxznSOvQ0LEwN1/Ay1
CVH7vh5j01QxbVDyJkmXs3ER9o50asL9YThsPWnKZoc421V0D1GBKxKu3VreCiTl
VkkxY6Zb0biUV8C58adayN0G9Gz86Z3Owk9XiQlKdp4YEPWnOfBnD/v3doTcg515
FGQAE+zyXOrFS/tmK+BlIcOrwbvTWG4hgRuA6VTxDrU=
`protect END_PROTECTED
