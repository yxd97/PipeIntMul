`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYRRXZQHCK9ofPq+rP6dukm74riYGHAtu6P0DODKv8VmLhZbzutR1Tramm05m46t
3hRngM4VqPbGaHQJqnRB3U+f2NAAMIuYFQn9J1dPyEe4EnZ6i98bwbSEupYbN0pN
7vewjo5f43tfAcPvB4uL3Q2eGW2Q2W+rjLNYjv7M7v4eL7qkvT9pDRrOp1fJp2IZ
H5Yp7Ba+CxnekzLnEZAaFKZTh2l/quiQ4XzIqYRsKzSVBQJkwaMjteS6AbyzMkUF
in52qzwrLAXPVs5K1gf9ur+E2ZniDh7GqnvuyZsS/dpv6e517z8Ugsqy02JKgRFU
hhL7hN38U9L70EWvQ3F9NefzNw25p+NQZjEhCRCtzXAOjhSOCCWnLo5We8X5Myg4
`protect END_PROTECTED
