`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82mdqPMli0Mw18X5htlwqddfxyOsYimeFrUXTxciq97lDfSdWflBFGaP4dHTtiwL
z3Vh+MJcvaETZGBt6EDw35A8tcts0cQM2Xv/a72ZwWWjvUHhOF7/sjz3GKyzQj0l
Swvfy07Eik2jdOfWeDGoFhwZI9i8f63cwGtIwi5TxW0jgJWjrBJ5RG4HnDwQ1kyp
ClYzYXDtZ8hKNGjJFt4FKDVF8Pb/Ji0hWjk/pIAP/qVEb5k/owECjvV9kpCWDNh3
e02e1KCShy75HGtV8DlVT1djpuVsg4SDkNf+eFmwp5yuyukt0DsUVvxxEtFdFs96
VInMFRRpbzGL6jfu0eqR7BynYU7duhB3ynPzyFDjncA4BG9WGQF4cDJmJcE9pO6j
cF+VVVJxTOYztt9fx1DhAArdGjDUm8Th4T6IDgBaQPk=
`protect END_PROTECTED
