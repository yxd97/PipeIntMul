`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xhGuDTGNZzzeVyYcDCCiJo+nwpBq5/60sJ5ZnSVLpakgUhJ76K1dX6FT+6g3fxG0
90ytUvgeIqgZ8VozWyWw3nPs0SJoMKVewKv6Sv7FCJeXivNnGl2cjeJjQh0VzL2F
IbH8GNqpjwC9yWCtqVvx0Qp7ZLENRbuFBru7t1l1M22HqH6+3Wdj1eP7vN1D/FSJ
3/yMAuoZI1JF/V5HdwY/f/gL5+qDHiH6Ix+QgNSGo2BbXsm2HvUrE7O/5co5xAXD
bv/uh6epBVTO+3U6wqQp9qg34QBBKyt6uRvxCh399XhXynkh8zaBceGcNKLST6H7
PKi8u/58uYUJEPjLP1jrh5bGOQawYKIhbYdbxiNwtfaiRGeie1OmexH3s68aAbay
yfZZ+xouN5ASceM+P1u9CcpzSekuEtresfxZHOdOuw86s43uWddKnSSz8UEfJBOo
b4N3DxOa4zRbJrwrp6BfbdJKMh3t87vvqES4y/tOsfkHkc3IF9eJ/zAlJwIDbN/r
FFdp97PhdVqmRsxsIfMLWjGYJUbi9EVMTY12xsRCBfrhWk9i+5vNWTAM+GjyoIwJ
MsE34NdRmF7J91S5hplbSCFhMdzsBoH4wrv6/MJ3VeGzJQCnqaeSsmWYuNpvlfEH
Xe60s4ZoCVxmEseMothJOR2gLUgRNqRcmvZBoUUx7fMpRRnMPcwPi3ttk0YdBddw
4evzVnuDkBG21XIxsjzMfQ==
`protect END_PROTECTED
