`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fzKPOasNGLQDUZkpGSgufJlwdG79H0NI2yd+s9aQzymaR2pQSq8KBsqubzD6bK9x
pG7sATRDtzfK0Vh3qf3hvvctpImHyaYS2yoZCAGfIO7ywqRdkXXr1qDGTVdSX9Ex
zqSdgEp5qep08rDW0OxPG+FxRCDIZR5/jaSb9YwAuz7kHEtkeXusJ538dts7um9y
cOMzmOIemat8wZ9+EM78rpws3Wkd15+R5qJ07VG1AYbDtSW0jslgNH6U6o55J3B5
9+Ars9RIOL2XWVIFwJNBUdjfc2FgqJGH1a9XASn2vb4hw+Or4un42WkaTi5eNyNx
NZekTCg38MSe1E/hdHcX/VAykdI6qt5YSPhmv3xWF+J6ZOk5jE9crc3KEXbyLjQN
0TAdoRNzeIwDJSK6e/cLWQeV8lBbuarvwbCgpBpDYEgH9dQmrgRd3UyIwKkPWmHt
MAtDXNIxvhEw0Y0aoSEHCrwN4Jg7EiJxC7FdR9jN88ClbFFNREtDzea7knMBYx7/
S12j2m8jDe5awetGDHX1bNajSlTRvUFF2x4cLA5MCd+Y6FRpz+xl+ygFBuBapVln
05l+gC4ZUoYx73TKrQkjOBxO0yp5jZ6aHo19050ba0U=
`protect END_PROTECTED
