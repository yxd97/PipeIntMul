`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/ilrwiZuzHdA/aUK9FYq6DP4HckY4bDfdM8dIzQaXoxJV1wA5Y9fyUS20f6tvYZ
l8AV9ZIwU1Q8P0aTLqRQF5hDMcYh+pS7wTiHh4MYbU6whNAskBfsJbaKqEvsTPRO
UYXyvvzZ1TndEQn+x9F/gIw+ggCBR/Gcste2seoFsprg6/B6CaEui3iIIl6tIU/S
3W8OkrcGl9PVH1TbMcR3yelHubjGrf1hYoGI8Nx8pE6vIkP6m3i2Nze8KMWex79j
NwHYheqPW8rypyL/8FGGWlCYmn0OylQRrDTOwhQHqPk/1w2XEYlHqyFT29+K2Ebt
9GblCJ7yu1esA9widbcArHUwN84sMlOr4OBrifLwHeR1stnGYNHXRRQrEHc1i4Dr
JPU2ZW5mq7/iGmExYXQ/aVc7I8HLNZZtIq0Bacj6YcNggeGhWpT2UYRHUKyXradq
5bizWV6ds0YsIfqkhq4yq9+2BrCqIb/Esn3JToZK+kbi8QXqkg2i9aPePI20v+a0
SxcWLUeRM9OhNhXlQ0kMmZ+0Z8tkpvVA3KIYXw+NUsetTFzrBPjWayCFtr9rr5UP
sMdJQVtANshVaJ4pTOb817fGZN6BnB3O1kL6jmvnzzA=
`protect END_PROTECTED
