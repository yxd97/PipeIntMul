`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+q4kCDfR6eWpq1G3C1YOrdBP4zTYxYVFpDnIMaKRJ3Yeote4StD9W2l/oucW3mRX
KprJ6bCtk68ffIUNuvC6HkmTp5ozylJF3xhqvIVXGzUafuhgOyLYUzoOaeGrb4QV
RBM0NQ+heH9c4MpYP2Nl3RYZB9OCEJOheUkW/pBNxso/mdMvFkp7XaPWV16diwXN
bWOkkgzi/I4w6RP+c4rff8SYcTsbrPxqfwhrihR6mDRcX0uJXKHqNfiLdn6Pl55r
9A+EAGuifUK9T6uS0dNpgQ05uWOK+PFCqi2rUkcJX55mL1Wt+TtZ6gGbhjZwjC7g
SClSuu8iYRPC1RQK4iZ36vwY4LIj1DpPSOdfrjpi+QvwXJwwfuE/q0LTEW5oPf2V
j+nQN1bpb3pS119cOjP9smHbSroJ8wIeIkcTjrY/R1j4e/ni7+fJOG+nY5L08JE5
bQ4HaeDgQPFQjzJBkovExvsEXdDiFHt6bA+J+/U3UARcsdGogztP6E1y8Rcd/+R3
1+JU1ED8i5lzH5H035dVPZZCsp65D8I6ncNhMKxlzlRzCW4Ri4Q5EywlBLPlwPGb
HU8Lkv33Y3I7KEsm6wBJ6agC7FvPwQ7Hg8fDZrrsbeaYNjGYsksu1xOdBLrwFwfc
0g4SHoHJn5LES/cYewSoEoeo7hVuNARgPVYgUXRD3OPxxwfWtyrQwBW619T2IoJu
RZZvPtpRljxrQe4cfC9Qq2ipFdXPBAPKtxASv6PP1zEfDIZEHVpH+I1vJ3uxDgEZ
POjUpiB3IzsqONSffpR7G3k89mTFWKZaNLSspzCSRklT36TNigup8hxWaggTDp8v
JZiS668G8ka49cnbbYAyhRezeFpI+8NfuAqQun6nLxpqlQXHyD5YzZV60db+hJTm
dHSUMJF+owNn6o6gAILdnPdnN8UDE4kHu4sKVHJZ22Bz/oSx9jIb37F3ZwK4J+z0
rOB58Ugg4liE94lxXpx+ykuwaocOBGWbbT7B67wLkZGoA835ZFf71XHm4TvsUdxt
xyMkZRIJG/JIXrc1nZ2gZlyAqm9OyvuBbdiApRUyHlXmlXcNGUxpobMgxmmBr+Xc
/qY2MTBn7JHNe5gcuA/Xha6+fCjSrBIPffAbqFp9zDX3JpggryCkqSAkybNmSoxc
Juh9vRZZtyTAWlYRzhx5qQexYZ+QHw9W3zTUodvjMoSDdTIB/1oIh+SSJMWfYyMy
e9TH5cdWiBcThAhv/1PK1t8wCjvcnZVarn5rFiJ35NY8/5gOa3p2HayyClXtiNs+
zfbOUpFZmNHAmbL0vHrz53YXq/N6RVs4SBPGy/yfyC3kVboMIHI2VNn3TsCnZr2m
uOc0iJnkWFfEucqQKAr3TwiUCrhySkLlN8xnhUGH/4jUG8l/dw7eY8DXzGBK/S/8
stUJMC54Qx2yCVDV5Sv3reWNgjgeWTC7qNncKI9rMM07CRqh3JPqHAe834V52xlk
RBWDhNs03o0C0jYtUbHrqnE9SnMTaFB5DRSYWdEu4NDYKF/ayEVjpeOpg2sW3vpZ
p8ABXjic3RXtld9xZE8nPPDyV4iAnwf7UoXVNm+ul2xetK6C3c1yu3/HW3Xm4MbA
8NTipL/Y78CaKXQFkNmuvJCvuckJAsugnYALE3aTltHt5ilPhsePt4Ncku0ycdz+
y6O1ahSZQtpcRgNVYDLQaLZIQeqsz/LnL8p1SehjVe1Qa1FkzmsXgIzHUaIFCA0Q
rBkHrKMW7UlofI4VZ1jOxrkj5Xd3GMBkWPOVa4JItZylZ/PvOyK+96OUvllbC8zh
l6yEcHvOtZHRNpKJzwGOjOD9VmTw0ALIxLxSucSvxd1c/Nkcog3Fm585YYkn2cuP
FLfUpbnXmfL2CYlVJ2HMj0QpExjmfZtLYUCN64roktjenI+/p4a76c55nqj5kWnf
Ius5FBjcH7LXX18sbO1dD4G3d7HDYdKZx3eTYy+VbO4OsIqAyBb25PMEKqslXfqE
nhmG+j0j/DWY4GMR7RE0aUhvFSkibHjpR4Bl7cI29+Hhr1irIoED0OIxZVn8WA7u
LGk5FbdojaW7rhGfgDwzQ3YAVjuHXrHxDdvGSS38vR1rTsCtrQ38vwpCAuXI7KFo
S1/pNDt65kwBWILQ1VwyUxx9RJEN8hHmfNJz7GCIwu4h9hKx0zKaU1W1b8MF3xy3
x2hZpOJ0jcl9FaNPdsBOqNUMV6bJEzGUjgrmeo51GtwEQ4VfpM2BA4ptkvj3HtL0
CMBfBrtgjgZ8CfH1ePmxX2FC/BQJG4mmz3H703TSWdC1EV6j7OuZu6oDRX99aMBF
cU1RtRA99IOXvR1HVexRuh7dGX16/x+K9nUtNdF85nrFSbLXSKm54vEggNjETRMU
ONw82OxVaYqqETZq6IruiNhmXvWqPpkPQqJI9SkTqOJXFq3ja16Aa4gcVZ4yGTga
nhkkguAjKmH/k7FQgM8gg+mzbCY/i8F0ec+iysgWMRC4sNs0TVzpVhnIN1499Rga
uda2ikUFLWlcnKIG2G8MH3XDsnCWG0YgHR+WXLzHkdSSfCvfknP8UMY/SsXSfuHd
XpCfNS727PrTFoJwpLBKPykow9a1IFXBRjXnjfP8K2DGsLHmehbbYYBqkZlvbvus
dtQJewphZtYmO371HzrH/cL76AbQz43Sk5+iKLJAI1HzqdVNRgaymzSKyRyDidLQ
S/Vkk+UG+9yku+PEY2yiyWB3+2f9pFCBNMIigTXi4zTKuoHxwpXVUVZ2k/ZSiCcw
zZY4NplLDFznhHWT/oskx6Ze5lk/9cP2tsk4ktu15bzLuFZTVuj9U4mhEWnhKLne
AmUvO69bdJ5zlTchsQZXKCYIyygL3BWDfZTAdw6px09oc4mChomUDhJbbapxhn4v
s0hiObKEiaXLhFru7GN/w8P/Ov2E2hKqVTVc+WEO+e0IlEt8bH7H40iU07n4z2hQ
`protect END_PROTECTED
