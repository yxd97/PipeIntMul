`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dw57HBBTrsZ8QSOUojQCu0pK+RyX46OaOBKIWH9W6/Jn7WKPf5g0vES2AKQ/TjRo
ac0VOZu/nNRLSsmrGzeoljojnrvvyYx7IPBzANxVmbudT36XruA94yIWL4xRXSRT
xftODiI/6Q4OfTIWaI8o+6aAthz52y3qgND6ZQmgi78vzNbmOTf3bf9WHDJSoTcc
IFW4nRz37YvLPG7ASZqxyOffhf6XMfqfT7I2iCA9u3l8SvXsOPqqgNGbtB8CJGr6
Csomr79calPjAqeN0uzPAkkG60fM81/4ApzQqkqdDSoh/SGnEhzV4NjulkdY9SQl
ujDkbh11+cwgESeXMU/mTE7OrHAvg6IzR1HG1vemWdt62svRTZeOgQfUFEiMZQMC
9FBslpCXoYV6lP23pWNSWKRVp8t9hCLGVYqSZPVPeiUFSqHE8/ZWXcVgMj1ZYFzk
SeIhjUqVJIYrhq+nO40jEg==
`protect END_PROTECTED
