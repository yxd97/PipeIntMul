`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qE3hhv1dngB6QJUqsBCtweQ4mg7qPlnLSylIYIMZYvhHC4Hpj3ENJy7hbYvmG20a
3uE2BE6/nIJ5B9Bly/Een9crUdrOUspGqV4lSHt/VuokitTRL7y2ENZNZpc6s8S7
NDhGLTXEznzRpdK3NVlT+VYgTru1KU4qH8PzvHOyYyVI4tMQVKAGJGcLujzfZ3Lj
A+Z/FNWrMusIwruY1ElkLhTxxZAYgA4oqcJGzcxSzVHMMseD6RmPAIyvxFU1qKmR
HuTf0KX+kcmQdpJWt03SqTofveXUIKQV2u+9LWOgcLW6rXC/AfT2nxlCYgT1V8ht
RO2rjMojqO7nzLgXpndXB2j4H7XFvXZQbHtbQecxoWozEGjlY+ou/6sb4YZ0LoEg
Hk147DRFR1qhrJbz+QR0GwB9r78kZ8ZBDFHEwj/bKrg1+6ScgF3xpvhvxpwQtXRC
NnRrlc+Z+IBSX0J6cVmgMXErw5QRaP8pZGi1KcIXDOwFOdexOPukh/RwRVECLUCR
CuJJgv+Ar7z5mjJlYznMOXCM7SscRGuSpwC7qCPrBvzd8RQAGeLbUFEL0yBrSoRj
I3NvuQkXgleQrbBnSmaeRuZoSzD2fpFGYXufDpd8xZxCERmwpfYqZagxa7vKq0qp
2rM5GXL4cd+y2xVtJvtUgQX0TPD6+l+uf8V9E+BHuBv8QxgRy5ZgWLFmzdcZoECc
DrIV7IERqL2y63YssU9BDezuZS15Q7O+46XVDbqpGA0cbxn3FzcjjafTAnLfEw5U
xT672m254C4W7HPFuoJluDRXkDKLCmzSQDoDu9P//gac5VvOLTc9m6d+dEr48LOi
IFc74fCxaxOeo4kYHKjAtLBoZyoOlcsVI1rqqH1EJBpDZ4qV4mHDJ2CriNd6dpKh
0ZQXqHo3CUZvlHa8YWTfVge+InKkl7WQfJiiio2yg/cltcxfZtNbmveFAu8MHaJh
F6Iz/JkMmZjNXb9xka/DvnpOXu1q7DkKj8pTi3bsGo2rlllfKTnHkJ07KcpH1K5J
/WpgTRc9xbRxYAG5WAXsKJ1A1A0Zh5DUwmvkVu6GwJyro06Oq/lE4hVIfqHY5adN
JasfacLIRmiECOpGjzbUpvZO35k10Cv202vrSV5CCZL1KzOm/E1l9xaeIJyPbSoo
yD+VicMPmLvWx1GPEjXBUha7cikoKKATuYYZ0tE99ynmbs3lolvluyxMsN9nU+FT
G3yo5JpFlWnKCQ6a2PUbumV/CagpGJ0Xpwx0aN5hzs5PJn6AQLpgmNHOMXVYonOp
iVgGxmwrb1IxEMIA/RSkQixdbygmHsgBqRWJGhV2oxZqta9A4F6v1iCTwrxTvTw3
C3mduedt61GUYyO5kkXx+1cy+9WXLmLOhWRaNCZUa0BbL/stZ6O3lAF09q7sGGZ7
gZeH10oNP/q4sXigswWUKtZ/2QyzIi90T6YQL4VdJv5mBb+Vlnb9IBRWnuae6oRd
Bz/D2Se1C1G8WEGS/GBttTn/QBOWp/3xmZ3o9UYqcwTh1z2S5kSzjx8YS54pJxaY
ZMTSttZYmsi7JTQJ/hdUtg==
`protect END_PROTECTED
