`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nf+4VfexuGzqB2XGyKsA3VntUxEOvZmWsV+ydWdkehGuBJxl8AEF1FHdMDTa+Zfn
vH9oGDqtMyjwUVt9JPsdO7av+hzCHH3zhb3ftZFHLfz/d0tX/jSnUZCa7Zr6yTRC
BButQjLRQ4dzapd94wy64M2cwLE6UmtiMkysa6y3Tti8ZbWXMpb3KrPkTtF/uidu
dLov0DskReLtAcSutO2GyP1ge5BuxhV6ZVcNk/LKC9hb1IOlJqZqEAO7RgcjPYtD
iWS5omiILFcyxdYwdLMKktvZc5f79fZ0LDxhnwIWbdo=
`protect END_PROTECTED
