`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LtcUk0FrBsBHLcpM1+ry76GTotGqiP14MmI6Qp2+tCtJfYO0S8AXasHhisVQn47o
nCm50WTD24rnXAkhRy7poRq/A3ahlbfIvKCOklmj9/c+lhN4jtV+MDPf82wPXenF
f4srYPLGBqNAHGszWZRzwKKJ8/ie0H9hIsQWVvBToi0pNjDZCn4gdw9UntKYRGNK
WO0meouwiO2QOiz1/ixjn/tlkLhJ7taZs2iLb3oqJ9Hgu6GrDVpurGnB6U/kAQkb
g+J0Tl1c/D6PO5WRay2nngY4ZEq59jili3duZCWaE0A1lMmQg8GvcoNg5ZG30NMZ
UQH5m/kCo9xIb93owy7Rwv7PXs6Eph4Dvx17K5ffH7BSADA03fXWbgEw60RkhhHp
XF6dJHoyBZoaV8tQymveFMrYDhTBUfqUlxYZOLe9EhqchSpEnrVIlGongFocdz3M
ewx7XO3pYW2Qd3qQCgneUQTPyueDTRnAFjMSEv/axL1Fq8yXqvcKcUjquO6A5oTt
02h7Rf27mfXsd1uxSMCJyQsP30IBnucRfzvtcFVM/HZtTMTWLLvm1NnUFUBtN18F
FnYcpGbxwKUJHl1USTZlVu3SHDVWilxXmvNeVuLxFuII2w/tTTqTkYYWaZcBqNsV
5Bh1hY8oQIvG2gLmrh7bzjUhUGX6WtZBRb84HRKelv4DDQ1/LuiCs8DqZLazRsdv
O0rt9vBGZJ6+4JJjZkODA8jTjYCyN6ZIdESjo+8ub1aKGXByFmLEHyYDz0TDOzu5
lPIZjyAKPXH+UmcvQBVfFB5x2AmtP6BeOJ8Z+obZDrdJBYT1bv0R2Row0SiZ6Tgs
F9WyGs4nEKVp+GUpXD8bgaEDnO0EDOmJ8yzjrID3FBmHj9rFwPSYYdbMIz2ev2Ko
RPJ2yVQVrHK3/TlR+7CLGcilRtl+4LBhmZxR+NnTo07AgwapcnxVkfDPk767QBNr
`protect END_PROTECTED
