`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xp91U7QSZJM+10J+zpAfn1tq/m3AUoRNEYxCqnvLIo8pquFJ6HyVHZ/eem1G069f
T6wLjouYKVgEogmMzzmCSgGCXosLfpvu/ZXNBqdZ3s09561+iRSpovm4SFxkA3Pz
/w2t+IrYt3FxpWzH+HuRnV+YfYgyooOjPPf81RJp3EIJO+5uIEaNdspTzmzFiSSV
+d+ZtIA+l2tiYufjsWej1AEAXYYTrlUKJAFH9K9H/HptsciqYHnp7bjAamOEXcco
Byowo5rOnd+02I7kCY1oH7lkBbej07/piellQaLyBSy6wAbW4g5vuOi8IZcLq2Cd
SKsSw8rkA8tF6pIiFihxcTkYhvQtcNyYOaWlsq0rXwt7kDf2dnYLMX3W91OutHqi
9AQ3sJqEPtVx8Y9iADQrNw==
`protect END_PROTECTED
