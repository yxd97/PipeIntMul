`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WzcXHJvru6FX1Wd/1gb5fhVWLT0Y4qRcIMm4XFFDz58dX+GUzh4Shw49xQ4QJbA1
PE5dbhnTzexbOQ1B1F0/bPyYm1SfCsgc0NZ+Li8lE1lNsi871128M4omwIFB3Pj/
ma2hfaVh6Frepou1ziiuAObGF8roY9ZGMhKJJxMSwUbNFpRVwnGT80OC95fDXsJj
VRHj5/+rbzupkM1PZX9QXgCFis6NbzbEKOzP78V4xYJ7pjK+53SCvAlYfMNIb2Qt
xBt4D5v43rgB8vudYMDFqugCxMi/ORKH8PZNsQ3ZUZ943MVnq08MEJ41hd2NFyfC
kmeVopYLLRP6ilWYOU3mIjIrX+egB1PRYpLAynM6U2mEIHbXla+MQBPdwonPBeJQ
2mZTlY8hBVnFevtGvhf/feDE+o2uaVM0DgsX4FG1f6jFZaZ1seS/MWsW1ySAouVn
iv20456r/JcejUfeBxCnioOmI4Wc4vb3tN1xa9MBz9RDbo4QyE+PTBvmkFoXoUGI
IpD16udy82LiYEYJnZj/8YCT9flDiGjz1/uxeW/O0Ju1TUZ4EiuCZMj6/8Yfq1rx
BN+DjZiTMFWZJIMxjiyVHTmWI9RQ6zFzUKRde9EaabU9Qx9OuC/5qiG2Ftypi9w9
LRo9lXnSyKjSb14EEmCpDw==
`protect END_PROTECTED
