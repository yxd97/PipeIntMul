`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3lxZijzSE4tjhLnBKhw3JzihVzj1cDWuagJHC5yGln4AVklVKPuorPfoZhrxyl4
DTZcBUpeUuz0GoeeqMVFgFP7adM2VF9L7loM9faBRcXCSkgrjQRX/8fl527iZnOM
qfmWOi4HxtHsaZHLTqDJZILZHTXhvlHHuAm8f/zUyevzUTws0O/SXHnj4r6MfxdV
4RGcWLx3lgfZeCox00lGBSGBUnsdjfAaGoj0dEreUXzem71MWXoLu3hqvF9L6ONU
gOyNVhnd1fVEkVT3VO++cOyZn2YsO3pYTyEWpnnlkum2HnZfrNsYyxzXbPyzIT3l
60GSgyvOp0T7oyqHTyDxU05CdHPifAlr9Mz9hHkmC461OYJjYoQ0xJCcARbtnA+y
sn16zQGnkAhFtgPdr5Rz1Bz4fetaHWzOJTbQDbR8tBENtukxpZnfYXW2J4Ue5GXr
/X70GO72J6fXTArpYzSlfmR4BkNN03Kj89Hp4r4oDaI=
`protect END_PROTECTED
