`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/e3TbWO1bYbiTKPSXwnZuhpcnJxUHHJLHuAd+p/6W/UDG3EYRCgCakBxrzhqBIIQ
frNA0e7eHu7AwJrCmlwPvN3vQ4GJqvqsLMZM3RlFwwRx7Elmyu6H07TgBOF0mulN
FNelSdSCX3HmHLywzaDOSDCGgnCdNnCrUEqD1gBEoTr+ZDpsSc2WeJ3M+287rqd7
0cjxbm7+QqQlJWH9LfxnOSMjBa0Yr2r7FiOBTVZJGxQ=
`protect END_PROTECTED
