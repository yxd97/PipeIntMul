`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
avuyZ8nmYkmTOiEWttGxDxFXnS6+eCizcp9qIo5Xnpw/dAYgBGcrsrdjcVaM1A/I
hKhHQ4HTcObSKp+wCZHIUqsd2y4PWJXYyX1SvsFkAund6Z408zTPBon1kQ1P9kjh
M2nPyM/yVcJyDo+8GdA6vzf2nrLXqzWIAsvFJDzFrJr+ZuPFtBNg0kRHXdmrY2s2
GIuPkOnPfyiG5UbwoAhMVozR3NdNehqfsE4EYmYd11f4VKZveNyRV3FAor1uoOjX
ssNJSU73ksyoy+2oNgCK5g==
`protect END_PROTECTED
