`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e2bjWNDD0QQW4pgDqDt7p4BLoAWbujEkzhNlbPaO9jE7CWeLQhzk18IZrsdPr0cM
7Z/EpAbiFmAiHV9/nnhIH9KEob4jUHWSw5yUKtbSX7fkFH0SCjIgwAlKNvcuqx2l
4mfxpeo/dXKeOzL0GOrfjjs/TM2hV8C6XOzW3J39mWVJ/LHFg86H8JzKpxpxjZ6W
m/5ds5ygLmBjgSgSf8YWZJyNfv4wszvF7QIGR6R2OLQ4g2XoKXhF+2oMnL7ZRVNq
epwUgn0eXDrZQs2+VGQ081U7KDs2k6slAljOlGC3HeeHPj6z5UMWF9d6ncWXsDBf
BhmWYF8VteW9SJ7Bz9I1wJxdRmuU7LjxOxAm2CsNr9Qrt50U0U6t/gg+PEzR2qnW
Q8IISlK6BQURFND1UVm1p7fMvV6jM2b3vo2rLQC7OGQCkl/1O01tVn8N/URdr/Sq
Q2Y58C0yl0O0Hz6wwD5glpXl8F0FixIFv4PIPCR6hmbLZ7ZMlpXM59RDGCKb+Ew5
ZvdfZtMqNJnWnE3s8QwXKYRlEcdXHMSvFdwYzxjgDxue37x9amg2uHmk4iyHO4Z8
bAG55dZx2IHfOAJNgrVKV16LS/MvTWVIs3jtGmtRmQyoP46WGwaQsdsYa+EhgAYZ
J4cW6A7Z+3Df81UemMa0FIwfPXKjuBarBYF9zSnfakdKw3VbDETWuQAu5mQf+vcc
5TZjGs8LBwCm5pHC6ySL0oKS0Me3kMMgwDpNm/YJd/CycDIj3A9J6e9yz7mMDYqm
0zOyoDb/fjUz8N/Z6S6O3yzmyKzjzM+bbf242TDr+vTtkOMidQoacj6KJ5GIQcL7
5vkQ+OynZDYpRwmvNMD45lAohl0kFb3L6ky2alVyJQxRjexZJdBJ0wJnRpHD/Wik
DHaVTNDkFVpzICO2iZ2E/i2ek3k7wb+gy7sf5UJkuJ2VetLLoaELn1AIPSt4h6WZ
8I0G+eAuDMA5aOEi+0y5Og==
`protect END_PROTECTED
