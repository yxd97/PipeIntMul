`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQHXMEYMN2erfg/sxyJeTeeHB04ZigD5z45cdlu1WgcnX9wCMySvd244D2BALobw
ueHMCuk84/HbHQb+Q0mHeUR+9afGYLT3+NXJ/qrvIPxpoEWBjkS2Em9Kc9nW+c8N
i8ezWLHIl8fuhVDmATD6CW+lT3lcJpgF35DEbJH1s3v4OZSK1R5EzNvF/32r90qP
0uKenE82nwsugo3YYW2MEhQ3uppb8iw9QsWQqgt/idC9Nj7hXDFs7DTL0fSCCT/D
DlP+jKGOFWLuTCTqpUO5fCw0GeeQ6XvSF4O31trucA8c+W1y9fg5iegH8ve8z4jx
H/vW2VPt7XVAZjBu1U2Efl/Scelj3q+ah4XtDX6w4byuDIlqtri3h9zam6mgxZwV
vOZ4X4pFntklslAlk0CUHzJaoB6uErO+JIGWa5a6lQsJyXVJN4HSzb07vxUSYON4
iGg0kZKHfBl5aCudsNq6zmHjquFWV90jlQBUV/YwvJ3XYbyHkmeOVA8RrKw/2YZb
j84eELHPSXKLnz0rL3ZHja3sEp09fpJylR1ZqxhJKBtxJ3lKM+R4csq35N8nnAig
UdP60Oyd0Pb/94k1OCClVRWlQ7UaRRJ5u1gfFDxbcXtnoYg0vIIYBXW8b8qFOqpg
67TNIl5uhi+sGvSId20TtXWqZ7JopR9zIlM+hNCb9CeCsiuCvXCoM204TzL1zhjf
WcZCxZhk8tO5K7Fax7ohfrxUbS6Fs9xFRRcXBTWZzNPDOtNFYCmmopvIYemkBL2X
hdyZ4TBubXaAhDxeMSrOf69DzmsIZEg8iaiwpdzFMvAwqND2z5BYyCXSx3BsW+PO
UiyxgA54qXRkKOpYlPC4wP6XmWcm7GOsEGUgydL+Un8UDaT+Yq9wiKCkiD8POmqG
hgLFgaFgvpPOLqYWjuWwfK/Qw+mrjhhGTc7A+f/SUZ25MYnW3LrUuPZSNdL/qCVJ
NP+IlUo2z+N6ZM8XhhbqyA9bVYtefs/ZEg7bbmHMShD4IIuK1sOSGae9dpW2wa/8
aSTRryJCX7YFpmqGCnKIOHxFOjIbY889YZzbBt5I6R4=
`protect END_PROTECTED
