`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vfrhxiefxirwJTHZlh8L7FvKEtaykZa3WBK45gnlRTRa7vGJ2OyQwhF+JbCJObSh
97k9DNKuehRUxkQV+5x2QA/fxxjuYEPqWvCpERnTzW9O3MWXj+m+5sag4ce4gP2z
yuuRa52Zm7WqHoURIQvzR2nQJXF6rCnEpFkirzQ0/tRbCA0sqwtbNLWBGgbRY/DB
o6ZdtcWppzoGoMy20d4O+KKaNBiRZWQI3h5bWbXU5m6uLGD6PkQzE7EC/q5/SyfQ
sHuaYVdaLKWMbNvoGOE2SEBgQCsnzsJIaZQH/ZwzlIF41tuy+fkgt+9sBGhbZr12
2+oY3uvqg46FSsVAu+u3wA==
`protect END_PROTECTED
