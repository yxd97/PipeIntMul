`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8xC88aJMShQDqNPGdGK0+7wUjzkXXXpvYY8O+c6j6pPe6lQgtUtzV0/B9UyEqQys
ztdTnj4Ct66QhL2TsbIYeVnQPYKIer202K2oF6Kd4JILukXIINMUA9H9O+N4OYyd
lk/BhwS0Hwnqz/6uVxVTje+UkdMKTgItDBPB0OH5Mt34NXF74pSZv0KEop36v6wc
Amorrq70LlUaUVdfpztpIn+WX0y0k/KqJASElzXqjO1AfeaCZOrULoUbcnc2Pgtq
Rna7v2ZQ/IMuPlv8igoNqX9odhTFviemZrsHDhJ/Gzf1uR8In1YOpkJsHmRvreuP
goKpG/AmOt9D9a7Dy/+9GMKR8dqYGRQERS1iStqunTcOp4RhO4ZXHApRMLKyGh2+
/feeTITFC29R7Ue09tDzAjStrKZVYJ74NEwWo9IuyNCteNc5f1XkZSxE9/IWXcLi
n3ohlclozMBUBmemvTgYXkIIwfbj6UN2au9yC+HwZVnX+JsxJNEH1vma6Sud0MWX
0tvUJxsmKPYdkfVhEOmUAWzw9FZTu6lUxc/pIdyy1ovXSUSDhVR1BjM1TCtcW0Fz
VfBoyZxKCIYPGI+WNXiLdUAAxQbvYQKpfPgcLkE9QLxYSVGRaWvS9RexhQwI1bBg
Ertq5JWmzh4pjg9Kcz70jg==
`protect END_PROTECTED
