`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sb1HVARgg21YToX0HAGYJSpt2PhCQzRZwcylbtfDE7W/VXspWtWktRNdz5ttM/Kv
PPXh3VbbelgHWwK1C+iAaAgSquZbMcMBgPmYCLv3ey+NEjfIqr+r/kKSoi2twj0F
BevAJTGQnilaeWckjwRPHLRoGdKKHIzNxXo0mBIQsaJxPy2q/1MtCVVCPUf+oyqh
lj6rWWc3tnEJZlrXqjOVUihy0A6r+U+D9z4lfGm0NxDESXVky/oSLY+7Nt2qAoy2
FVmT1NZjKybw8S6Uq/QYN5xAaWWauM+mJJtBBHpr9B2GFt27bb49rgpX15PrW/G0
16RrQLfQD4/wKSVPFh9wWNbLv+AwUCw6mS9y3G+9dZzrirZUM7BRlPDDKvDZ5jif
3DTWGdFRozt/HuvjYB+u3SINZtu1XEF7mQmdsmY+X0b4RoVc+eUzG90/qHQCT2Sz
`protect END_PROTECTED
