`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X4fjcsh5HRkvuC/rCDl5cw67mb/zpN9Y+EEinGNOpq+TuWK3QKjO+aT6JNRsO3Ax
6Oq1sfiEUftJFA5FVwfKGeo+3DGvr8gd3C7EGeed7T8AiFdrxoSKHp7+Q14331OS
lpcma44EmSfPsPqIGjoZ5S/L9E9XQr/6SFN0XGrgh9hWaKByXUQPYmt8Bzb0lXUa
6YI5vBEGp9Prz1i/KQEn5MOMFPINT7QI978X6gjLKot25FdY0wcksZE8QgcRKTL1
ZODBzSKMCSzCfFHhbJnI4321OlLq6Q1THiMp4J2m2+EEu5BQqTyKGfPzBHjwPquL
yhBL3dXr7xH5apUO7OrisMr7HTduHr1oNLGAJELAqFrn4QbsfUXdjgK8eSeauz1k
RwKSpHbxfyV2L3Nj4/QOQP48BFhLRY1ieo5lfVyoJFQ2rFMwXQozOXdEH86f6oqV
WCcyrYkLNig6vDQ1jeM9R1oDwkfDTIwSFZErhQ6/adZFCD9JO9pHFUcTqv7xvD5l
iGFP1LrZMmo4AsbtOyH9uXmYcMk0kvyBmuRg/bmeL4YC4mpyQvuO+LgCInwTKz7G
zIp6zDNjncdDEFS5RroLEdGBfeltkVOg4oUtKL2IoHbJoOHi+z89ynS8XV1NZOvI
ATNe3HUtSWGaxq7ewMxQ+uz77ytLa/o3+1hKT0mZ3AjZZITDJIlnXaqC8ozMDjTH
c2+UFIQaGYZtj565RyNNPgZKTVShGNVsNKHJ+9/nhY88Z//B8BIiKTZ2Xa7xBoeD
5O2AF+BQpIQ/ZA+l0L4lSk6P4CpfFhj8csMO5Yv8ajEILVBDvtarML4If1wnVawr
DZk585HgKyZt/qWp0nhJVWP9SjBugjLbm0sAZcZXnsBSvzxDDh/OivnOidD8fa6d
XvB42Gecry8VUxmP/yfgPBNgcg7LZyV8WxM9NpqmifPOVzggjxgE8Ed7/P69XZQh
MFdCDD7PSU0WuiX0DBvO3GQCE62qLAgrtZ94nVBhybhideFx/Ky6Ty7kn9baLBtL
xMb2sFwldW6SRwiB2Kj6Te15K0wRcCx1WNyYROxG4YsKXIwt4pb9EqNt5EpruuON
XZvuoeLtd7OGsoqTYPBCf3l4s+yYa3KU7xAsSoFj77jpb4OEGrjcGu8YRcu0KYI5
SuJ3IKOZbEcqu0wVBz+ZgRTUU/2oUkN2h2L6PhCjRdNEkuNRVfSVEB/PyBMo4e0n
icjuNpRr9FOz0ibRndPdV0/k8Gb2Kz/RqH86adyeAtSygsfrhcv4YHYw4au4kt4E
Y2C8q+B+k2wVO6H4MXZp7SwqQkFSZ3JzmGsmDoSlhcfcpsJ5FKuruoMjdKACuK6H
v6XEAy+itf3JNRfYXmimD8D821vrUvOHntIQWZgNmy6YuVU4HoNy+nVpql2nPo8J
W1y1bzwy4lqcPFm0xhRhBSw2LdcKsurDrhy2uS+NvPxE4JLhIUZaP63xS6O9X8ON
zDPTFyJad0CgI8Z082MDHbgxlOmSV7LRfFE7pd3abKGUU41OjAlBkj5HYPPbHwxU
Xkc8pPIrW3FxH589hZQKz6ZXtrGjN2S1DaN5yKirLRTQSRz1OjTs4QHPQhha6Eba
frAiZaNq78Wrl4tDduvO8rgoCqZvXiv46aBH8c9/EoNckMyurvVqSii6gEGM/brC
1vPSHSb55r4bshJRL58cHqds+L/IF3ZvdVxYJtNNnvf5BY2O8+/hROhkzzVDpR1O
HuVUeg76R3igndT6JG44zfgSjohheJET5iRYkFpG+4VNkFfwUnJ0HtcRbkA6ZfQe
3m8hYQXLkzKbouF9eHYcmgt19O1F+Xg8PdhYPhA0gjEHbJ0l9AhLgC63bMIxb58q
EzPcQP2mWl2zic81oiPXCfXpm+UlsYJm+OhJCwtqzp0OPHIexC2GdBi2bvnCEo/6
Ff6PZ3hvtxkXt9KraER+7tOu99tVMu71WNyFr8jzymiHpYXuBD+WuJVwdCbL8lWE
3WNXpnfVEPZi3Vd8r5V/ABgqtKbLbjwFnKcWXau52W6Ss6rgj0kKZ9qQAkg7Gf4h
P0k9LJKVrjmOMs5pPK4Zcyn5GGPg5LajIXxXUvRCdOYSSQCbZ6XnRxnS7CMrqYPW
AsuvUj+ZvDMqvGlifLxr/yp9k4Ee6gvLmrljkCcW/fyMlZJ0kiFtB/U/fRm3xDgs
Z7ViZbG6f+r1obLXieQW4GlfUuWiJjZomSa0MdQZTTlCv506Jy/f0ReOynVv3tEY
+b/nNXJZVLLXgnDYNTzJ/3AYldWPN1wH9jqbD0IbZB7DQx8wsrnLxfNzdKDBHOlo
49I+zXQ+7jARLfgMUVnb9IewJ/Ar8Xa16EVwNu6LaWw=
`protect END_PROTECTED
