`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdBPaFVkdGWao3BEGQ37GBAiPvem8auiwxd0Qqnq7I43Z7Oxf2WnYLPN6V8utsgI
v1V/ztvCipF4A4KVWo9hFoE4PS6m0ycVPYmysdllE5Yku7a6ww5MsLkilNf73u0A
SNfmAr8HsMPY+WsLxk0X1coBvwPw7GjpLTznVhinL2+ORyIP1VyBo1g7hXCoNs+4
ZHC4D9DrGrgrSVf5gUxxmgmeDdK4nBNDlYAj9QAAYWa+p5Y07B9sqWBnzKA5dhSm
+CP/2p2qe8EbZWO1OaGZQQ==
`protect END_PROTECTED
