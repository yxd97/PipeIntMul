`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9OX3bE/DLCDobnU7CckfWjsetUfnjU17mwwkPhKPatYqQaK5kHPi1xiyIxbWL5Qz
xzn2uHh7MCcsx/jFVM60fdhR9A7iuLyB3ni5Lvlv7tjLNUxSfLl4zk4QRmqsDtMV
Kpo0+/EbCUKK3JimZqHDc9iUVaCuFle+SpydsPi7UndcW3YFJWmWxJEUSynIPtPl
4gNEW9f27swwe+yXjNd2EE2tb5KRjOdWDNdNLsJ9f/Qn5t7yk9BKEln3xBaBl9Rn
IpHdL27fGy+7RyjldULIXjkt3gnc80RAEFIRgthRhN5YY3YHOifCBS/FE7Xl6bBF
HHwTNhiP8SOhBZKCRGs9diTORFa0CjQR6JHw0c0Xk9jhxEOuI7TxspoQrVU8wOON
8Xvyz3SiQ9ZHaF10EG5DZjrGl8YTx9fOM/T4J4UUhneIplaBKviQ1mGrodABTU3g
/H1GmpEtwPO//AafPp65+062ixfbR/MbOxpgKTX9+otQbDbqRf6fD+Y+ZiEZau6D
BJl/r4JWS0BKALZeQCK1qpZYupucLH++hkCOJdEaCFyPS+zcQmlwICgwif4uFjLi
XLvjEgMiP/sLXIsVjYb3izTdiwBlkakECH+d4PXGf8kXKFVT5yV3molJ6bbwpXea
6QVA3vCWycn5nsdUf88GkQ==
`protect END_PROTECTED
