`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fLA7UFfcp+/tpwOjLPB+qlZN2j/bXlCSP8/wu+2Kcm1MgW8WLsLEUtkmafbfKhUC
Jm9zGzvT7ltFWVWFzihOKkP633b7GaxMuD+ZWCrieDMETKZUKnaFCRPDNE4y0gYE
vROnIIXRZ8+umweMcPNdnRfjPsW0etRquTnOEYrRUs0hTsgst+3pcVsEcb/s0T/4
E0L8cjbyWaVo/fNAg4WzvPohH383Fo6Cry79lTSqq2FaB6mmfm19iRVo0REegTUN
8Yp3xAaP1B+eB/fSNNgSFEzkTCds+j2ssbfxp7PAhZ2cODMNtNCX30mmLx6N2nZ4
TCZy9x8HwyJqqW6lhrcBmg==
`protect END_PROTECTED
