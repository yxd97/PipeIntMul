`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HljjyplxhCMnUMYp7WEuh2QomeF0U+Kmk8010xl+fkximQ9r32SXg/MTDxUMbSAC
SdmVQBBqhIa/2SnSoRGciiyPw2gV2An3DOrYS+3Zj/0w98G+JDUWiR6NeU47rZnj
j9pMZ3JOPAKMLoKRxDtQQeS5O9H42wszhmtP4yn2QHIcIHtzufBxwlgDyAYqVlhc
3HhVV9YJjsGd6u1u0YqA+8suxwYTnHwarjGaLOikZoKjzm9q0ZP59r7dTzXuEXCc
/RwwQ/baoZYIQUNFCgzlbkA53IHduMO4LwUMlE2c73U8Xn3GXmKoxuGCslnhRTHh
4NNPPXi6VwLuTlhYlcAYUF1rSvZHEWSdPS9zr+byYyHYRalI/WZp+3H95q3eTWSQ
1JSy6FCHXFlhAyrF0M24fQBEMKW7KTDKd8rSXXljWELO6WRbbr2UhKBigKPZQJkB
s93m1vzf/+CmG07iPgzboCPq1/2Q1VP2KJEnC5N8qvuCQr2GtnYCD+BXNXpIbjCi
l4PQ+yt1VRAfidm8bfR6/otkdLRe3BqbbL/eOt7WiPKF2CscxE9Ma8Y3I+kWPzdg
BfyFVBxtuhnD43pLtr/lzgtbJjy3amT1niaKkK7WhLVY/ZVVOkW5d+MqJsOyPnIQ
0iqlpNKzwsxbLpnSaFXKRPqKKNYgcKh0pIJLt2b/C8Y=
`protect END_PROTECTED
