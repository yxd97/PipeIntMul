`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JePeZ7/gEDpLK8j/rV1FOXQ5KrSsTYPKGOZXGwy+yLeQ99pzCIOpdQvVzg6bLQ2c
tjItuyUhJ5PhHAFz2OwuCe+X3PsK/wFYgXCeAo8QpGVM1+8z7BL77+9bkWvNPeSk
77M1lozLG64P6oe7aT7lYYEIJXXcUUwJFR3hNH+WJlGJIWh/otsiPQJA9lPc4JZJ
flZ6c6pbjAGSGTSK0tC636xi8oZ4WpJuUD5/0xW4MXU4/0sIJzRNWCq+CdutRTd3
gS9PTaVoZ52QNiGjejTMJg1zs1r2jGGD7Z+WuRgp6Iw83nVYAx7Qo2vxxf6enHc0
1tqCv4JNsOjQn6+9V8ZsWv4Cj583mBSYhJkFP4wsGqSVeSl2y6tZ+1TDa0KIaRxo
Plhwz/8/yMvI3G/pYjRObZqPhf/WwO45JYikTG107PF+cUcn3tfejFWbmgtrG6H7
ZHMNOqhgHg2kXRaTDdqUB7W1jyIAIog4dC7PSMVkj8MSxes/TkwE2awQbySNtYbu
Q+zk35b10kJQk5RZ4Ixt6zk6iN6XwplMfXOPDpJW0fOrn/LZv6jRQkcq9lVKDc+j
pQgnCU0Ut7liylB34IbRqadjj+3jcrMkWIGGbCy9wKmm7J1KNE//EMvvNm4YpjaM
9mQAez0SYn+EG/OK509T9epe1crm/3FeI/883mARWdjBypZTs6P93wPZwg6xdjwS
PjLPeoXpehxIIRm3J259c3u5VVofPyZ/u6Fe3ClLFjYe6qzi4hfMjliahc0626yi
oHW1JWdQ3th0tWIoXmR3vA==
`protect END_PROTECTED
