`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sjlJZPPoAcVNkqWD/AHtOdGTiYiHbPWT07JWIECymC+M7vFv/1VqPNPZpSbmG9W
NdIqOqFiOwJjtJ/LZdTwIT0vryIwF4FTtnS2NjfMgNJjODC/CEWmoOmAeXaQWCnl
5aJdgnBEREHxMJz0S+eu5cMmyv5PExi7Su7+7WKEjfLHry6rBxF5RatQAGiPctze
oJF8Wghs4tX/+UhknbXIg0z1Le6ArHhwDPAcGh80JDjT4Vdhcm6XBeeoqQ2oiILv
7fD055J8fsFF+xC1RSbM81LLUJ77LVXcMJHDsKjZus1ZGRPj2RfShLoMLZ02xNcH
1VpzEH3JPJCxsX/FJUw7ejtkTYlreF97ZlpAVxGPf6ODDANLtorRfZ74x13HT9/U
yPrQ+vcHYm6uVJ/NMtWE2s5QZ+GU5gr1WV3xw6wxyp/2gro8RBWnuhl4HojRP400
O9t1adYxc/2G46GktgR0UUi0ALHqCsvLFefblfAIvsP2rd65U22CeW6I0T2C2cmh
se2VvNC7STUv7igIu9AffG1u+eTYQi1XxXMgCo+bt3BS4IPz9qtlTMT/ndgpG8Of
1RkKyHHSA4H0JSSbOniUGQ==
`protect END_PROTECTED
