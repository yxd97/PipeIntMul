`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cn4SJnNvwPvfv+FQwGFkrxaynRHVT3Txb0gXKJW0E7k0fJ85A1yKwNtNt6/CMGHz
XPsBpP6U4WqeeX799DWCRdTnATWhxS986fYfAmGedRc4mEOyDqQwomGkkR/JEK5Q
odTSBVmEncXiCxhNQlalAQfGnP68GfQIQqChfbhVI/IgvSBR2nEKolm7nM8HptPh
4qod1zPmI9DgxvsKSp2xbyDR6rwTZYACf/JGIimt4Re7UNx4WNfX7arF5/gG3/e2
PdUdhMCWVGQmy86KepAdOg==
`protect END_PROTECTED
