`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQetc5bOGwN1tgRYZVhZFi6EWbAGKvPChh6f+mqSKEHU1nVbSLTtjYmbD+Hmys1x
CrKPhqCqusrhaVII7QkiFw3sAVpvZFjX5wApYokOrE24CFzpnTd5pkQnaxSe1YEo
eJPkubrvkv0gm6XTZYLAKOgxipjKNCGgJqpzbqMTVO9s+TzxY67g1CqrRptce0Ho
Ctnp294fY1HyXnuQl9u6zh9hGCkpQtNYNxZd8BRzP4bzGh/99HRX2Zlrp0SSuYDU
eR0KPhSmbPH1iSRuf5PeZg==
`protect END_PROTECTED
