`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THrSqkntdxJsLG/q2Y62ibf1RYgSxVIEitCOGEBq55MvPKhAcxTWNkM+j2JRshP8
D3bNWfugqHva5Rx9mI2Rm8OGqk5OGul11OtZY2JQ1hwy+ElVFT1AzQa1UwH8uoQK
KaF1rgKLcfmEJizS4aOkFIQVmvJ241jzHSB1sed7kjZ4ZJR6YhA+S5ENIkNco0ZF
qV0WPagjPl55S16hX1mNaCTNBw0FLwz0DJfWxtdRK81P50mu8MRsfxExEeJRh9ch
ohOE0xpAZjBxBTipxPwIxNOhz/Jqzp8H2Jld4FYjfP5uI3x0IYcJlNqbyj0yjHdm
+Z7n4h4d/C484ejRO8dFwm6zBnAK/9akepjr6eZnkHzaj1dbaY/nyQDRCgwnjunM
1hVs9fEOwT+4MqtuZGOOSmqwfvAoAYFQTc0MvoXWIZbZgTlnS31WNC7oKsiqFbdN
hmpTgTBdNzyLwVOD+rARn0sHVkT1VHapqBtDzYefeWH7vVN4GcIsGM4nePZwDj4K
gaqxV+XzWxQD1itmYcrXjw==
`protect END_PROTECTED
