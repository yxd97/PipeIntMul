`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cak4Ynt4JOLSWutopiXwKl5Jq7jI1RAIHedOy9a6EV0Yrl2A7zj8HPlWn8ZQRlqU
fTJDgySbM8oxrO9cLZhxdtyva58QYO71t1+mfEtrKAxYJ6YlWWHBseXIJCseL7Av
fl/hFc9kjtcI8S3/hr/LtT4LU95SEbcClNKHT9JVHhM/duUMrZsjRewm5Vlblf8g
+nRwyPsn7EElA5A4Ay7ZAe56too13mFw5jcwe7Ah2SSfXqtQIiodwlQkC/LTXfhu
PfqgAv9lEaMtrBEhG0VkATf5gdF3fccayPmSe/ktDvU=
`protect END_PROTECTED
