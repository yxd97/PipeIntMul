`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOlIjlNyNWkzl1Ox5gzfwiKWRxEnEsguY9CV0jcrP7KoyAhglvMiqbTLoqePeLgg
UZm9ItaJX3gLulv9RS74dw+Wwd6AjUykCShOwPCB9CgzK24b3rRe8EF1F2XEFlNh
WKGlZ6Y/MoPRCLeXg6JgALhdTDHdI10x/wUXgEtSy3NAuuPO7liVW4uNwMBEU/T2
CpNdr9m4mfdNaPNNH6Kuoib+5WzHQQ8PbC1wss4gg/QyuiTxhGHB7WhwECRPnqeL
FzdEfUDeKPE4xPblGcHVfF/kb9t8oBsPWTIGmovFM3T0htMUFPsRTyvgsqG/PK0w
D2Cfjx1/BmzbrOuQNs6NI+UmqyxWqzHLJpSyLI+clBSHOMmxzZ7BdNqFwSG4hipH
s8eKwwe/9F/usuUnqjWEb6YgB9+TEjg4GPQU6FQIOJc=
`protect END_PROTECTED
