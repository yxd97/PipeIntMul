`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9My3SfiEjtHuocv/+mdBo/jV7dT/dHoTD/qA9GTyOlU524MbqzRfOPtQxeNY2Ce1
MGz3x7ymU+VDNvXwLcHr0XNBdr8GjtX6tfXJPrkOesYZfMs0jDoCn4U8JQ+p9Mel
sRjDsxmbvUIUalR6F/AkU4qAlol9e1T5Mn1rLg2cFuW1P0GvD6OYVAVVIdBhbDlE
HFMgxsjbDBGhLntMT3FW5EN6LNxEPAouBAYN0iuak1CLc6AqpmRAhuVzDKm26qC+
M9EdT1jRJ88Pb6wH47WiWp/tcNdaqy22Vboeujjx/aSJboSLcvpn5F2b5GsCFP0R
JvjSaKeelEHoSXXt7wgq+nMgKpGpeWY8rwX2MqB9WtSmpkeYJTDgdjPlLnPde0f/
+9+5OibkvsEGD5v9CIgbOufA2aNJUVoUX5vSI0spuXpntEEKJoOEIC7uE6LnhHRK
taYggf1uv5Fp7ie5KIpmFGhwI4OvUSbm4QcBSogXDVbccLxZvW6evrheNHtOK/BW
5FYHoYVUGDRSscLgBBSnZ9qwh0inDetYGI9AKuKfYJPiOlTtKhNl/dIA7h3flIOa
eAUTnl9AvjCfA0iEVL96lPZxj1XD0sCTBIO9HAiaq/lti0pSEovHpEzPIwNnO0TZ
ppGJ0Iw3h6vWIj+WdGV7oKlEsyxUpOgnW6zvHa1yc3d80pkHyL2n0OB0zVo0F7p1
2S4U0il4KzLxrxA26VgrI4ty59D+eIbIST89TeWVGicJrOZ1nfD56sOddQAUlrWn
RwTpz4PrgbXMzn7aga7ykr7zPLeEgAUPnGGB24oo0s+5ssmvnYkeIYI7qQ4Uuj2r
vTPbF4uj4DQ64gRIt2DCbeNVKd44nQResBabKEysKaVYb90sNBkvyQ9cvdz05I1A
89v87yy++cxgU5jdJ6JZJREqAVmbq12JAAOIEP9VKDfmzSQ/WI4XbEyt3pKoS6A5
jTJwiUO4lndqvtarqoi5gcXulwQC7dnjOTrYoPLzLOwFKOPvkqDtHm0Kcq52l9WJ
qkVFm6iNESV+PLhWifihFrVIMx2V7kUVUNf2HkbeIZbJXStIqEalYQOK3f4LFJj2
Zq0i4qFSBqjOKsD2Y7rcy60GuDtbAMQxvLcCqcVFiIFGZktXABRQ23CNHCeNNpMk
O8FZOL0P7O4V6tk5fR6kU9LsGYHx5/eqiJh43+MD4e1DmChvUdCK3aeVVD6y/MMY
7lVhXQXPUSsnlrSKYd/e5QV0GyC8+9RC/r8EeixoQfyr3v2d0zne9s+ISRyCAUDx
ZglfJMoZkOpSOl+SZp5bkXMjbKRyko6bV7vLQQP2CcorT5FUq5I5yPG25MNb0xZR
7PNldYYcD6UpLFN1bQzMecJrdLnUnq1LscKK94JUfVwMoki8t/2RezrEY6vBifFh
93I1X0KAZCyXmHnrmeo1V2Y3CZP+01KDvwNj4Q4q5w8JHmd7v18xFJ7MfcLNwry5
8/f3HmKhjxa7jU8/5W4FY2jqjKYws9Usxh6KKjF4JIOKlRj1fZbDp08gmBq3AObq
7hQ1dge5ITd9x+ayB6PVoOEjb8UhRqVv58uq/O5k51wcF7lFEAMJGz2NA51Zvl4K
GtPV043mZaP/73tQyIu1tzFDUr0n1zoRpmCMDOMbs3k3FJ2KxHlC7xkhCoDwYimQ
wN1T3eqfRBSFMqxMFw40jSEyzoo5zWC2oX5mJm7LE+W0G3HZQL9YQqnpphan9+LN
VHfaOyBk7zqMuNobxQL2AYREIQpnDwBoxm8N20TXybruedRPtzFZWy5cYI5UULk2
6SfbAlYtZeb65E0AOBWQCuzHvkb4nBlEhYQ46tiekNCdhfYJq5BLD/FsYr906tNi
rQKmbMV2hfKBUbkyWIWmz3uPL6DIURv7FUUtjf2vFviIr2BIaXB/PdzK2639r7B2
NDSc8MD4r/+njS1R9Jcp2KkyoUy3ErBcdsIHZU1wMf0AndNNA2kysxk1c5Xovmce
PgXADj4eNKCBAb15j3D2rGzssBKIw98fq7dsEM9fntkWfbO/VT/KLwzqaapFO4dt
LDVNimPdIzOX3s9QCv98eEOBaUqrrBcLVyeGvTQIFPekS1x9bIvWAplVGiNYMQR1
rtL2ZD9PAveUlmFGdlzBAeQhFnBU08bQDaY1acHcCv4nDjHNLuqKBENgtAnfuhRf
QIyWovayn9pnm1UmXD7wftYrDOK9HvIE+qvLh68X8Il+Wesw/lLYs10urKM4BFex
Xk7ew/hQ6MIU5BzTSZpCBRwKI8qdLN1Kh3DIOwq6i10CokNQGTHKZr5Oc+8IsL8+
KijKJ51xpUW29iT9uAggeagNJl56RUorJ5zagJGJDtyXwmx17TwYjYIJsneGhhgR
Eftu7RngmyaVYRquYdk7hYk7/eHbeN5bKyG9qmfZQMeKrlXNgHIN6fW6b5u9eKdT
yhhIBR+WUft0T/lGs0l2ENT1x3avoGoO+Ej5m9R+sPlPJ7VnoZZFR8TaerPrsu6b
w7JrTwkjU+DdsMMLrQ4Nn1kMNnd9tZg0+a1/Zqi+/WWEyUt/eyUzOEeT/uNz7OeQ
H8tXqr2t9GIeP5irNPj62+DCVl73zvaouSp+MwyK09mUAO5SIF4kICnm0X2rOYGc
EhCSJTbUMPdH9t76FxI+AudxfbDEXsQCYkwLqBvfma0R2yqaz7sRYoD4f4uHzzKY
GYLK9kySOphxaUe5pdDQK+QT9+BNuM8sZKKpntN55Uu64g9ennTEzl8xsm5p/ApU
09ogQhl7fPpGKlHsLYT7h9Xp2vlwjUX5JnAmrdL3oIVgDBS+S+sUxVT6p6nJVIVJ
LRd2SgwHW39MWntFkP03bmGIrs0M7V7H00JJGvubLV5u1m1Gr1+/uzDhofD3dbeG
6MXXUXJMeWA/Ev+wAEpRsWFjj7LqhHNG9ghLVBCQbYbo3DuWxucH6tLyYO2iSc5L
Lbt4P0n1iUUxvJnH0BC1btJDHQUaTcY5yXqyERJoosnrcOKAyq2IwC32EX+9x2uu
2Fk843lxJDb/rfNoKvhioIjzzyklroVH+7ytb1AaGix6N9Xnxp8qBWC/ykZIc+mY
bOH50pzDdggizK6O/DsBh66wjp1uygQUIaqfKQrdcjluL1jeOSfzU0zhZOBygWiC
yOxSlUXQn75okEVtWKAIfhxjVU9Jt71Cz50rytjISEr0+Buwsxb6W1WBxjHfbqSZ
MnsbNvjJGoW/NWGIWbGMlef3sGW4Jy/BotlyYL2rDB93s4Ya9SkqmtxGA3ur6a9s
fNN+Sz0qIIaU7QML3ynQj+8wghxY4DugpUPzNb4i3ttPSmsWaj2dv38U4PwoC8NT
7+eqU/ZyCXOc3eiWcgZVoTK0j0B+2ljgQ+l5vvL59HA+tI7yQvOIjJ8ngZF8QR1v
AD5OytWahGFvJtwXBL+rNdNxY1RAlOJycyruzqQOoSiNfUxsjEeMk7hbTIBD7ZPK
iL9J2AZeRrGpf78zvId8O3cMiLMLy+aOHKo9wMdyK/MgiKe3ZFlgAn0euI9WiwRJ
3PoD9EiF9jOWwYI/JQWemw==
`protect END_PROTECTED
