`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vyEqOer2tj4blkZPpRkW3jSUlSFntw2dy+jCOM8tiOfzE645ipCuQZvKisjvjbk4
jQjLjGih3LsOgmjHqqSyM4h/jjqI482D7nrfVAC4AUNij46G62Kb8rT/QNSkH0ea
QZpWeL/ggV1K72VA32VPRQ/weQnR25TCPPlvUQYYQP0hSSLTt68jND/lZ8/rTajC
lJ1Szep9rHsJbF59JALA10dV9le28H9Fy+rKwdbelnZV4kbA7Pz0ZNR8cm81kJAB
wNQddRX3KSDgFNFM+CAr6tjVPKd3XJTn3F1RAemv9UZVwtUm5XD1rIkChQT5MCvl
q5k0cqnbNZ8JWwwuB/9su7cFIdY2+59p8fvxgSdTOs1LEpStQ6UkGsWUdfSctDR5
lUfRUH/zjTmm9cIBWh9NjJ0c8KNRS/TRB9QssuXovpTq5iXgxweSsvlIzOrVkwfK
H5zMBU0oXdKrzIJWGSPatPUiBFD1o1RACyr+JNjsJ6s=
`protect END_PROTECTED
