`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asT5x/Cd+YJEfJK4w4GkbyLD6GL0yFFHRW/iI1mQwCkHAt5rKFogY75fIAWaCLCG
cEF9cV5kuQv5Z7w7vlvjyzx2PTZAV3uBVaEFyYHFyeMRdBtp/YG8lswMIEvY4WVv
Z6Pjyf9ezsRAJ7EmvkdnJyyq5R3oorO5YtAOJzf38haIV0Kt4b34/XBvC22I00e+
NXTD/S8hgiAK5y3lvu9G5spgCaBY/CmN/aHamjhWEdjPSyqBAWGmV+qJ8/+3q2dW
ljfskHg4ggns0RpyO4ZJ5Q==
`protect END_PROTECTED
