`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MxNJFGgb2Hn3YIbfL+VGSqZiBJBHbG7YETGCCb73cw4xv7kspvFwcwCqO5XlWDfO
o0ci2jhe1MB2xKfhBxqmrl6kKw3+C/boHn/zC7+ne0m9jQYtcdlt2VWASTWDAVPX
VhN2TDpVmv5hyyiXEuTMTyCGPQo7YEJuTyzcHTPuU77KGxR/jIVBfttiROFWuzho
HdNmGRaljSA9/mW8ko6nVJa2QVH32+lzvD1O5qui7Cse6bYnbQorPG6Ie79ycFRF
whNcDyGr0YzS/fLhoijr/M1qSpPyn1ysMkNQwewMMROzno2P6jIx9RjpnvxhPGkm
jay6ZSYAuv2kInCriXG0CJtoSnT18wYd9XgyKi567ouKm2Jvn1Yp90I37qf8gwbl
/8OxWN918RadYAZKDHLuEQ3bDjYK38otr6k0AxARuduEBzpEcOOdSjWIwXbxhyYw
y9s9HE+0OTz+YFz49cQAuC9A2hQcMOtBj8AnEPk6aDUjEz6OtbC22e3GO1nyUG1T
lhVQpPr5VzZA0SdgHuukmaq9FcaC++q/83CbXqW2TtejfWVWvg3k3GGERwfx00ar
O9XTdPSZ+apc97dEpjDSKnGNTJRjKIDN19XfnVdKJZHfEjVrt5sWjk5Q87ieHoNS
I/lzv/g/vCpSYZi+z9hq4se0Ufh0w2NwBEZJovLamw+8mCRaI2KmL7SXQ5QS9sTk
utyXzb5CMP2UIUHvcmjygNkPSzG7i6/ewxzaCMDfB9hBUzqLCc+BJMH5dNckNHgE
j9nW54LC2+EfBmgE+MbzE4tKIVZ8Q9f+Y1RnQrhvfiV9DS1n3JPTgNWM6eu8gwvB
L68TxSpJfpdmc//JBHtCiCkCWJtiNyNhJ1k9ftQpJV2EmRp00NwZ4ENwZLwuFBTL
ILrM5bqQHKDzAMhF2S8o/MedzDMJ0Dh8AOfN/s3bbiuJ8C30yemQAfxJ8/h+Evyd
RGMf4aMj0PRd/JsDLlhaIyAdedxGZmt5kMAk9bKUy+wLap7mP+sELzW2uxJTE3/T
SNqpA2U0nNIkHi6nIGfMdFP0auIzJZO6hLSmbFXv4QLjiXnfeRX1QcxxG58Q3s2E
Sq9PQJoSFSKMTDfZwmsGZ0d98eiH3LsEXAhpsXdD0SuPYpc+rI/u9d1a/SyaisyB
lxTLo7vyhvg3yumL93Xka3wod3Wf9aKZW9v9qWx5CPETnSg5zOf7/1QvAGXIjP4R
AIJ129M1L1/Na0ldDzfQ+c8j+aPFiHGcrYiFUmkV0/nC5wlHICnwrN7VLKZHWQ7U
YyjPdZWk0LblTVnJnYE5GoNLHrNwV0/Mz75RxeUoXd8VNgJR6gVXRIFusD7eraRC
oCxs0Iv+t+8uV8HGOnaock7sOZaQ0xzuOxKa1SGg23SIPjyQqFNAgYCSKkAuhTrT
jllAcn3WdlAh2R31E1AZ92FAjozDGunUNLLw7Fq1UeP654/y+HOhna28EasrGJRA
gc42a0VGWM0wIw1th/BUJT8lFO+tIw+Jq1cMJAmkElXE9GtRnprG7XHKJigWhcjr
mtgYKshcqoYztbAj01NQ9kWYm4ExUy4n/6gtg3IRu1UENhPN+AXjifkITfQMVwnG
nHIMAMdzoVfbB8XUTOSPnveJmuWIY2V2QKfLT+VLOa6C79IphcLm4wdUviERk8hf
Vq4lZLpSSX535O8Kw0ZuHp50nsKZxLiw8wkaRjGzfrhn8bmG22ClDEAd8ybQSojx
0Bnpl6poQKZMotnkkllG1kdXeB3qPM6/PzdNTluXQI8Enfgos4eZzc5Cr5cp9Pp7
x9RejH1Zb+bPFMwdnBG05ujcdbGqz3eoo2ABwry+z7aRTlpDw+X5V8OTV8zyrcr7
1tpyrUn+cfYhW8zCNpXhumIKknR88vpfRMdYV8j+mNY/YIIt2K/GC0RVDDrLuNII
Adz3kUS9lEIXbRhmiOkWHlybi9nlgN3bVWo3Je0oSxrHCz3CO7fiDR8uPRaXJfFU
LhlrDX5LasRVQYKviEepDWX4tUE8GnVEvJrGz740glz/AAlT7WJ8eSKaOBb85iIU
JHijLdJWkm5ZljoD6o3grWT7CZr9DkpmQ9W8MquxPl4wabl/KhfCDOiiH5W06ho3
DBrbEP2wWKm9TG9vp7sWKWSHjZ4iVN1equMdFh0vHATa4+affGGEQrE+tF8OYgFh
ZpA+LlHqCEXMp86lSCEAeIJIXfvWOLO5njIx6/se/KkgGPCDDwvANq4QRJXJSB9z
NgJ6wzp+XG59ofdHyBkDE+oBAOlQKCoSsCG3LozjZ0xibCnOp0PhsEvxpQYq927h
9uRAAy9qb69yTk9rRLjdq2rzYtyaHNjT/7pWipviCuvEvKqVNIdsfZbePvHvIrNx
czef1Dd0+Om7hSCC2E6rVxps850JwsIU0iKhWHHXzxkhIT0xKUI+J49Xe/93KbBb
Yc8Uvnx7qWyPegtoA74ce61UdXrjv/cscw1R/jJF7T/QM6fmytvRcwtV3mj0Cr+w
YIjYXZ//9URG+dqJguAQxwrIS7s03r7kTth9rsbPw9X4VcV9bEyNjx1gyMzR+Fh0
+nvoDCFYzmJLpAQqVtp8C1ZxDbyLu1RLTfnCADu1ZdBDoN1SQ75NkXZgsstapwEX
TxuKB7my0Fw2AUNJqAT0MVDKRXR3ZGdA5mPy4bOVj1QIz/YteJxUeuY5iC3LJ3Ss
pQEtlT+fLhUa++bWF+GXUuaebBdrCqTfha0Jxbvon37sQt4e7sXekRtDBC1v3QVQ
Nqu7mjGM8639WLnLeNsmq029puFxVDdn84sK25N8yr0kxkRcoa1DF2HismV5LhK8
b2vZlldCySV6oxXengoAIE7w2Lm50LCn+Lma1BPBwshupHXDk0j6L5JDj89FG3EU
g3YDtkpL4YBwL/IdrsNkATFNt5iKwWG9NsDh+aaMOuDMeIo/8cpJaAOUSzzVdcF3
Q4ty0xFBym5LdkSWCaLFoEm+RCwpFrMMm8t3Q7ySzeFFzx5BDZsPN75j7ZQfUdsd
VOM5NQhKDKCXJeZuoEoCloCEacbvaD1ucLBaZ9m2iygrPJVuZktSesi9f3cwmcUu
FXakaPu6ZUAp6JjdFUx7Dn8x14DBInxXllSJx0SWmHhBBy9USlMabKb9ecSWDe1q
yym1TYt4001Qvr8XszMsEdCamkVQ/lwI/jTQvr0m5WFA7gl3xH7cjy9N3C7jaeCR
WLu/Y+Q9UL663oB2mrIzEw==
`protect END_PROTECTED
