`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hASvoHsf3PLy/S6TFz/g/aiVdN/jzjf44JByAKx7MJ1Wr+OyC3BidKT5vao9Qvot
LLybQ3MQF7c58sNV36g8nBjQwLUWAW7yCoP6Co5LFy9oL393caKax5vhrRFPwwlo
yicj1uQaSy2GkcDYhrn6m25DFxQTZAnsvyJOk/XIBOXDQnORJQ6/rN1RLr5ezF+7
KdJz4DX+GUUg30tpw8rFeSWtUrzsd7F+JkeZ6iXJXvi2c6OrXNIu6vERcIX2pFMy
vLMFcl7/KHKMjb+LilEbJA==
`protect END_PROTECTED
