`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ylmJB6GTNev1zQq2gm7gUf6pBbHIgoqdddmoJqvnHQA766SGyQoYXq0zjllvKrjC
NYKFZl4JWvB6O1fMFpvQzukDtErQaivE5Pt1+8fbXxSilHfbaKi0tb7uWD7jf/c6
bWg3Qen/H1MxmDaBlfAA30g72Wc5UX9Fayg1Pfu5o4uexfL/dtmqwD+uabAERaRn
Q675/Yyu9bhNyLiqgfO9uvmQkRSw5SK5UyXNPWwYZZCe6uhMIcoWAKqHbrxPc3hn
kXKoaSxQbotjnMmQjl79lE+/ecWQO1Db5EDD+UjCyopWVQ3TOUNOHhyeRF7KPMMX
ZXe22As7sGHcneWrYOLUniKhaHwxVr+zxaVpzrD7xIioO2uRlXolyUZ3L95Qa0zU
7ExhqAu4tI6g3sTLPMOFXw==
`protect END_PROTECTED
