`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zoHZHejLBkp9La1hMH2DcMNJsoZ8ThhyPOiEICX4/RM3/+nQtU9LMGgEiR0l0G3h
UbLD+qwnBvSVSsUnrPfHoCYV47gp5lZtfK7QciiU/AsbDx60eTcwG65pJ910u0DM
K35im35sZhpRDbuo+nLwuGIFGcV3uSZc9TmlxyA81VFmJ22KHwxtTZ0xSHHwdEPk
ek8AeTOYxDSmXCz5wToR4iI/iYv0sjbGaO9+AksIzkZ3D0GiKPAyRPr2HF4NPWR/
DDr4HjUBe5zJXy/rtSu0X+N3ZcxJPY2TqoVFqgf/dY/ZX/oSC0T4spMMmklaHR6L
0EeCinHQutEkoLz+EWlKswg82I0Q64gsp4uTiUrgLmkTKzWicutnUR5pdzHReFW8
zkx3DOp01BbIGbrQ07+3Db7MAW4XUP94aipS8BDttIBbNI43gQHblCL//QvWPa+X
DaxVyr4pamw+ZXbHkTVXdEEp2GAf3LHO+Bm+bAq75K8oHk4LGIcqG4tdSvlznCCn
lDfZt6kPV+3W3wOZfHnwipBMEcTgLxgj49xJFAdDMYIVcMAtFVfLN4hgj9Xw+5eY
2IisTH1YX4A6lEjLJz19FpvRMgniAVlMJoDbKvuDlionYj/aGqV7ADMsJbYWZIue
XNLxqr5tFt5z++f7gJyd+EXkL3nIT5Oo+NEeu+G41vtubqH3M2/AM5zZeiyACR7R
pImbid9N38GsFD5Tvv1RkeoKPALn2qmfpANp4E0TqJLacyj/FeUxW9WAAQPpS+Df
tES5bBHvz46HCZ/tot9SIPUxJ5drg2hCY8CnrSmqE3O5y4wOGJdVuLKRUqX4UKde
RLStYfk0RyWtm7mjRZ70Y3g3mUBGIZ1/oE2QlymqZxBs8HF3A6MRIXL3uG8m7cxo
jaXLEZRFWw237KEiaFnP9OOXT9NUSS/ce4eVUmMUP/7PQYX4c5BAju0jCUILIi5Y
eDz2zaPJPm17NE8SXmtSiX+56WKZIqftdVW6xJOwpJk6evrjOqBaq86NDmQbSfd8
X3PejjKHSvglllCjCUPgNafPq+Du1xpttJLe0zGkaQ6F0mYAUiv6LmXmOo7xe4KF
aqCAMHD/bIHO8+0Q9nQg6QEgYTv4EXaiRzY3sNUUgOEgiu+q+2Y/PfQ2zxd4gwfK
YqD1M2sGp+x8vm12SuPN7wxOK+z2Qkc3nQPEW9b+UaCHV7shmZggjt1Q/cbuBDKe
eHwzJSw56aZjJw7aXEp+1uvA+rA8y7UmKHsxogqIgnYXxfqdnULOEl4hd7cJGPAu
bMVBNoKUoZq5+78MjpCHozklLgw3GuopSmO8lInqd7Gm71bIXmH/NsiJR19IoNV/
G3ywHOunDfGcuLYRVEBwDVGVgFMFp11l3gbP1GoWyQGpeeX36735JFbYfAlSrR5K
IARQWwmf+b1nDKQIFvfnYLdfQJ2vJQ+Zcd4Wvv0as5kh0Q0lm1cr9XqT6atyaE9d
1tgwEEPX2O+HjlEB2T1dCCzmXXzrK25hqgAhM2tzTihc1ggff6vmWrxiON75OAjJ
18dSZ9HbR4xhb5AtvzxXpAiwnx+ANiDmOvhsnWMU5LEC9Y+glXi3fy/vmEr1O3Cc
vTLIv3wsImqvGNuEe5fsdiCo4jLX6FOTyndhPnEQSaOvUmkcSzpv2TMiXSelAcBN
eVGR5Bj5s+lI6f3AEsu5J5GrCVqNiRCvRI+3Gr+q9CNs3KzDNbpbUWdPEoHjfH65
Zp2g5rpJ4QEnoIM5sxyCg+lohm7FVjPzl+2JdfNkt69x4iYgMgdN39MgDRD86j4U
tFZta0bJpAipwxit35nm67So/Y0tRhsUYhfUNQxWyQ26a9nNSCWYT5Qqc3ixSaYn
8N552ICd+DLiAY+NrA+p3GsBNXPvpsILsEtsK4o1xarmSprH+3jWS91IJeEXQ9Rn
OMuL5qA0aGTmxaBTSU/5SNfE+3TKq4YYGeVjLTN0j6EaImoUuqS6c1MtE38jTMMd
l+pMQFlky3CSq+fhO8jwjw==
`protect END_PROTECTED
