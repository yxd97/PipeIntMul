`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AM1H6+IRRtr3LI5XTWQiHVwdnp6EE+FkBtWPmTnZ8pAQWNXFhRFgx6qaC8XSR3Uy
10Ch+vn74PFds8hh5Q2z3k3yWigHqrtGPJQc6L9uN4+L04neYHs+Kfbw0tELsDE1
Z49rLdkJVRJZOetM3HE7VCd/j2PRjOXX6wl+yHyELi3LvEZW9/hs13hIwiSCtDT/
7BBEL+MHMX4Sgu88/aqSCCzTqu3PFZ3weZm8MU5w4j9Pn4GjmOdUrFZ1aeHIwmU6
so1sILH8eir9AdrNKoE94prhRWtvfP3P2VmkbT7EoYEmjHMfaHEPWRqeQKKiiqTW
5fi6SxD+SuhnXTkCvfm1LIdocZ6HxoRR+tCJZR/NZkSAW+QVi0oEBNMxNhrlG3jc
mskzLZ47fU7FmB1DkxsukFhz2td+ortcZfM/sv7GIUGXt5yoknVzu72VXgrxC4FZ
FeHv7o9dmz+KxwLEcikzbEKHO8yuemQNNprZpttXUCvjbKR+XDIJwCVLqprPZAKj
0jN2D7ws095KGmUmiBk7WSyxDOrHxMjKiyJneIWzO+0npzhXomYpH8lyFt/27qqS
PcDkzyjgpR3USVmkR6wY1pa2Wh9FBjBqnK2bTlb9m0rYE6HGkTqbkWbLe8GG+mUP
hZ7W6iFv8vDVE19N4WgKsg6sVE9Ar8ROCG7VtuiDsAcWSydjeqDnch59XXs7ddW0
wA+fPe9yDgThDBYtPRrQ4403RuDKAEYGrHRlS2HPSLifVZWZ9pCN6QJMQKYOIFBG
aFzVpUcFt5FkMHXFe+YStcTUGe18AlXr5jLBnlGveDKEkunaHcF3gO+EigPied9H
reFgEH49f3pdI0anQCSjMCtm2QpDbGHUaJabAabZkQhPRd5KNNaUwk8zRvb2M2l5
BgdvXE4/+LacoOsc0ng0bFg0Tbr5hiA5T9h/XHL5ZXYaufaN+82DAld/ZNZD0NfF
1GvjZjKwSwv5qnUE4iJOt7ETVzOTVYy/bCBpOcW5+NNZcHLIeP3Q0EOYMBta2h8P
5ysCahq3efUEczZav6YN6hun2qJFAc9zF+WV3kGMg+p0NzuTnQJIA5vI1wZKaf20
SUD9EHTUVKDpo6k307p3ldmfv6x+OJshXZ0TgGLkd/lk774dPOhYu3GzMwQfEAmO
vDnewZgySjvvjcPiyCWgvoH4rNJeWMFiEwF/EyACnFuGDskH8Q6/gw/vGwGihsDY
+T5FK+f4qi2dMKt4g7VwcgTLu2XHdHsayHPgKCPTpaD40gYHQuwZZ4i8OK1V6wGO
udS0btx8L7qFsCQIw5Ik28XGkfPKjpBzZY6fACEk5mc63w563CGJH4aqTspr1oFs
C6zdxdmONOwClp8NpB4NEI7GO0CQlOTZjEhcUk42VhlVoI1W2ec0A+7fiMNr8XYa
uyPd/KqypkDeWOKIFOuN1WId1mF0tHEoBZLq88E7FZCjK6KwlZRGv/E8Z36oqN0w
v6hjfYIdx2tnHsvlL0hwjSg/8jEH1DGay/AEbuzf7vHkV/6uyOh2zRGh7ysh6w6z
FTUCFubwUrdcJ2I9KCqtT0jY2isDOGy9QoNiv71j90rTbDKFMDoQ5UBe7+A50VHN
oUcCC7zqU7CN45qd4xjs0649sRprb4d3fbp+WSY1bzm9IzJFceBwoZ/jCyVxCNIf
MP7zsBAIsNogIBRLMa5u9NxAhdU5saSw9bd0N+9iz2XA/D20D59K+1jz4kgPLJxJ
0bQlLkomqSDD4oZBjJdsdcxMccja0cQgK6Z5XgUNlT10MVtNzP8/Gzc6fU0orTPd
i4YS3iob1DzJUxsUvmkL6Kix5/qPHFYOKIxovhrV0E0CVaxapo9f5V+dYqtrdFOg
6p7rg9WqCU7PG76lAXcUmHQswnu3gxCKkPnSgUTa4RKI1s/FPB8Ptn6cOK0EYjQb
C1itoCU4/qoeAzj/nP90tDKvZcxrM0FTxBzbySvN+sJAoGbda+BRzXpfMAk+AQeN
NoRBn5GC3JXln5hSeeZn8MsONUhuJncRHD+Arz0bV6C9VI9SmyAMHiIepo8YvbIO
IYoy3yaKUwAKgfMhqi/LezER9vo63lZDmIRFxUrHnbthyZHFb1O/xRNuf2gRvlyq
NiiWL3VqXGU3KGvtbXUUrA9lJMdxi5H0m3jYHWkXWLfP7C9spyZJ+I5Gs1/DP8Yd
ySNESwZLg2jjxVs8R5okmlWfGuB6MU7eAoUnEEmDNoTUCTLxD1CbGbE3a7/WQJIi
3p9DcNZMn+2HL1ycChyJoOSYhzzLCubHi/Z4Fm2R/TfWWGqg9Hxe3R1a4CIwJOMJ
XGCsRovedWdPkdYrK0RJcDDCdy0PHeKv+1kNSBcrbV0XBjIaiH/k7Vc1Kteh4p4j
n1Is6q1+XjPBx0VK8rZSpQwzAV7zzH6Uk/RWmAcGZ2+DI7cTZEOXTpYBQQuhCwT1
aAiFGjgreQ7O7kliR4tMPJxm1vhBP7cMzg0PBjEX0GV0kjfL5rhpzpsMMb3jrIib
8mmDaJYCPkfNDhP+FzMPnMzCKcTv9LnbZH6M1uSNxu3aK6GSgRwNZNLMQPyVKGtl
JT/2mk0VKSuSUsUmql3yk9ICEChOfejONjUK7O67Wr5rtQKW3DH/VemIrn//g/ql
lXdcjYNM6ChR+vlVoy0d/GHIvORZy40clSHKJ539Bp9kdh45kHCnp+9QkhXClKVw
OlXEcimxWRQKfzQYrOgwDA==
`protect END_PROTECTED
