`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n9UQYqECDHaflSNs7O5+lmETTf8AaugaakvxI6BjDMRRnyRhlMBdHedcb8nFQ+lS
PyNIZ0ZsnLDw0aVxBCyoCBAzAOF3zbWLS7qitKfLIVbFa2Yajw5goFAp2w05aN4+
QYPgKqNPTE6LHarVuDOJYpqYRhz3S3uJZrHwCelxyTF/WtH7N4i3ASr493Vk+Fcv
ZJME97YR6v0HIsRHPIjayUlDb3BLpFMeQZGLbbNdUaKZw1nECT7+8/wFGXNAKdoa
A4uEjZGBtmrmDtRjjR7RrsKj/ETjCL3PiEyZnz91D6b0QNpPKZgi5DhSu6c0NPlQ
VsmHVH+tfLM7M7v/PcTpqWfpkH2k0KFyp71N2a61N2XZXYDxkgCbk05ffeSNUPrH
VIeXhQ6OBxtpqFJ2JfCQitkTOCwyHd8iUvzd571IElcnJEMinvpjQqzZLUawI+k8
bpJx/8fo/erP5jvqMn64ZNEqfOOh7F+nfHsurkyjCamwbLXQy6JCxsSTnMDmjBN9
LnY07UTWtm17tHS3IG0XUyCE6QgTx/nyppJg83XjJjAkLJeWkjRcffv1nsrcVOpz
J3idOPEaVXd2pjj9QA2eDLHMgQelaipMDKYfj7hg/94+H5jL15QKDdw/OAyTraTW
3DoKsptRXXyGhTlofKYoAU01qkFILEoWtbNJDWkOx8f0c81sTA8WLh47ua0u/h3+
m2j0zpwUKBnTnGQoG5bvsELIdNDNT68InOyR702FnNLxr0xoTaJmY5VdW8dmfFh2
tdadKbiSrlJihqB685f2UIeq6tsupT0bqb067A+aVOT6IHM/bdmOob9CMq6/7L4W
ucuSIkEthgEB0BXrfFH71qKd0uk4flPA/I3Wb0k22bMQQ7NmlYWem//ctvOtllDQ
aZDuRjpaLotep5KnciwgEk1xhuglVkCXszgDaBgE2GagICwjTNnb4MLm1nUOJX+J
sE+aIT43PUnSttPMlsv3Fe/RIAYHLzqrl58u6ARfcaxMbGR/GN3m37eZSV1zSbOi
QgY7ZK1K/VtvTuktaFg27IGptfZS6zIgZAQFvN3iNCJFxpO/GMPY7GzH7e6rtNNt
b5k1k1oykXQGgxibLOSCR+ObC+mcQPPuWrXhsy1trlfU1DVw00WdqZx3BdfJtc2X
qhSZpV2sCEG9R0HesDfhY3hCUFWRjnp7sjfG0VzTJfO4P8Mtv293ufhKIT5EyfUb
ZqOta7H39UFlADgT6M5nhkk17jJemF6y73km9uzCOMQSjndbhCtAPjBm6ztTr0zQ
zYK37U/RAfOKlXtpvDavgLap3tW98XkFelv5lPJq1qxQ2F1TLvdm+li28aY/ZVPL
eMMjbKs4bAbtUbnEXmbXrYjrITE4SNfgjUjq2voa4sWlGkhNWQSB4o2UKWdOxGta
74G/g+VTzpQkRJ1Tb7MY+QZKpNt/WLOIZMc9YEbLo4FQIFy8c0/wGT/NhX+vWxV2
DC84gszrlKrX0snjGk/A3Q==
`protect END_PROTECTED
