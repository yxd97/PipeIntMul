`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4vkxyN5R9yXpLGXi/pI5erO5fdm7C0JPgfgPyGLSuVzJgZj+LUPp3dM+rlCsf9r
iqiKAJ+6dHSPEpuUvlOmWMfbX1rtWvlirScf6h1f0fcl2/ltP+2ng21lDQ+jk53z
DEEM/iwY2D8NBpgzBtkpWcLeGv3f0fZcoOUfKBfGtfogVm4jUeBw9g8bYVwgRUeo
D7b2DB6cYpjUh+Pfc4YV4Vt0s9rofG3sNYG0DvdT+U5xDSZiQuZPBPncghTybutC
PCCQ67cYaVTsVtnKytON6IOZpUZ3baqQDj1lt3rercRVDCxnPiZOSccYYtZB8EBE
Hax/Up24ZiFXegqf7ZYPNaHIVVoV8n18vs1u+IKhxHwH/8puyqyqimvzYoYMuBYz
Z3mtEM6MdpyI8XfZZdgbHU0FlVZ2S5qqu1IyR3XiGirpnGr3n7M96iBrfHtAoIXX
wvyrFHw1C6dPpQ+AyfmVUjn7bbEBS6lIc5So88HRmVv3edIWN/pWoTH0e5bDhSr4
PkqDJbv52KzMEZUntL+5Vi482JtD3hAwTdnucVaqwZjcYtich1nfHjoDGGXZ9+xS
L+I9KsLt2Fet5ox3Y4duEamgs18oMXG/WHBhq9djidCXXWfHujkklYsD4IqfQGff
5eX8vx/KJboA8CbQ75Kg6hwl2lgNfBh4zxyA9bWiwDc=
`protect END_PROTECTED
