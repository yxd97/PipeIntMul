`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UjIeWFQs+Meyqw854Kpt4p9VrEB2NpV+o8VnD9IXGc3pAA+5kyta82TgzIAXAxf/
GdqCOas3ODbUYC+v4hcBhHDBfO9gfBpKul9eq5vMYSslU7ro+WZfr1AkYYXfLj1T
lGyODoG6ArW/FLX6V/qXuHZjgia8MgC8McabrNJ4ulSdvzs20nzz70iuLcHcz85i
V5ZFbB+6nwzVwkqf3llD9PdKKjRHODnr/Dk/lGPO7wHSnuVQU2u+dIslKjndy2D/
1izeL3JQyzmIezTx6lNvpCd0OVv0eBlW1Vu1dYnUPFd14DzVJBCQpMdFoVqk+bVM
75lMODnpOddfvmWkAJPhBpJz+q6pflZWtT7bmfvye8jZ07OUVy3FoY4Uo5hvBdrn
bULOdeNc6blsasBRaHwBcjBs98ttC3WVCM7v724t1PAI0lHW0Xzn0NE5zKdyoZCb
5kDUddHqPQTNgvPMjZup+aPOlF4cGj6mK6dh+HKuYrv823kDthp3AR1IKlYoyjfD
`protect END_PROTECTED
