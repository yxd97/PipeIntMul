`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6SJMzipjPDk4QLba6S2L5gwd0W/d6H05983rtFnu1tPA2l/ZRzHbV82zNWFdL5+7
ZZ8mlSfLVEzO9k9eRn6cX2AVzNPDIAA28A2lKgJ/I3fQR0DbHm1mzMNe58N772+Y
22jIE78vKXGyoYySSH86NGaMa8MS8W9SaSga32Sj3qNJqElCqLMhQA/DZiMzKypk
XrdAvY73bf2PfSsyn5Y1ULnu7NQ7goezJuEzsme9WInQDDmNPzpcrRPfryFgxBzy
vbhR36d1MxO04iiSK4xpoLKVFG+HDD2iDWDU3ZeQwZKWmzErc4KTyCPfWFjT5L/L
bMFASKPOAvkLck3iFjWRM1b9WEcbB31O5TX4QiqPGAA3WeCd1DFvnSu84k6EqUiN
5hBRDDHlNBKA4Enp1S61dQ==
`protect END_PROTECTED
