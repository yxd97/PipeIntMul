`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xl+KXVPmTKTjQXtNZhPmPqmT1k4pGzpeQdjSYMgP1yUQRAaUy2BqJOv3qGwswlPN
xkoUsM7Vvil7f39O3Fa4B1opsFmKLQV4iDZb7cqjTcm/LA9RDYIV1i8pgiLTJqTE
FcWEI0EO36LwTbEhDEt4jbf/e78Y9TCDUItPeIV6F4prO31nHTdQ4swk4vivJe2u
lc4jrO0QDGsDoUie8zEW7FVr9sv7ZlNnFbztW1EOBgshDQaTv8wkyan1VQRRrNqx
GK0W2pMz5+IafUPBHYoCgr1A6PR/4UF3MUXfE+452GSs9ywx0So1D+IbmKfj+qP6
Xq8mCh6Yd/XLs1gsREfBxXJZCaajtCCsfmFYhZ67gUmqirzw7SCL/xI/7QZLv68y
cLRDvzHom6GrySuj/b5RT4TgvrdjFJU7oAhlKoRo9Jvkso2wDSkzTN6mjEZNMBV6
PFOw/3LYYFvhtVZ3AcQ2nZUzyZyFsmQRXgLyZzO3sRch8yORl+jZvTzjm1KobEc8
wyYNs3bc9cPLu9nQlldBjI0Hb1Q0cC1jYul/sljk/V9EnNPHW3YKLQj9U3J5cKMm
mDjPBY+67G0YVCMT1i14ai/LGULSWn1r2PzA9dXdT8oQzJLqEdgFofZ3Ftx+A+iW
wQl0gYGki8inTWghob1raNApU+9KCrnr37rl7c0hm4zO4JlXhgujc2cco+eNL0dN
9iZwunyvktYkIgqSKkwR1g==
`protect END_PROTECTED
