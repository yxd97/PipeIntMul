`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h72G5XsdKjEr6bknHoJt5LUahuuf++kBulpXSDtbyz2zQbMLiUKjLYQgy+cdntrI
/gedHI80L0pMipOL2r613fOYX5hirAKegkeLWmqA7ux3FbeDnI2UY73WbBj97fsV
zChcq/dhuZx01ma2ADGbAUAcHVdgc5Xs3i83/vgxcjV1ZFNtHF+STgufKbfEqffw
4tO65Zw7Odu+/b16zeU/5Q==
`protect END_PROTECTED
