`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+unzbke9NA/aAv+YI8hhpNu1pe4rf5X2lFeBDbhMjjp0oJ3AEKrH8E35EGzGOMy5
kYmjrm3XV7D+dqAr5z4BeLYZinh9WC91sPOV0k201GzK9EoDM5NMGkCc2xNBQDPF
HFKU1NGimO5UkMq5q2EIsIXJOFU/NGu2vh65FRKxhMCZBF91DfzthdFl8dY5hgPV
Tr/sWsi6rpOwLl38+Uimk8EOclY7s+92B5vYqmdyoF/viMLS6cuWTvlIB1amsiu2
WyuCiG0JCo5OGu67+lHUTsFjRH9gWFEdD0l0+j82youe+4uLFJughDAwegHbg3aE
Oji9/+toJwWM/nLh9leTg7gElyZL9fJG/uP2G7omTkPPbNgzRVbPbvhCUkEH2ETA
6TrC6KMM+6gRhWhF51KJQR7UlFHbJkyRS1EiArj6dgFGbDrqPnmHScAZwi5ZjXjs
31Si1Q9BZGneyOmMq1bHgpo/2VlrlLxWehFPFgHLl9bzsK2C94NDL7jmPHhG0nI+
1I7msrEd6oJ50z3QUjUGEWFwGZAwkeNairEld4J2BWolMysaFCMhdCAe+eCGVwO1
BwZohsDKYUISBKVxvjpWeVXR2poueGZfSBTrtEqxxY4s1+LltCLC39efG9Hny+yZ
iSOCxniIeUcPHPiLx5jllEHGgVtw3PaAiqaBYPFCm7/cvadMcusxQfQ196ZOI/Su
NLpjg4fiIoj/GncQWxBWiE4RQRKVrAuaBMRo7rXegLX5ZTyN+CvaYcVQ/v6/GrWf
i0yLH1NkEvMKDMuCBaE0Ow==
`protect END_PROTECTED
