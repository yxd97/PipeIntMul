`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bUBTLm8zG3e5jmn28nCWxqXS1PPXkeEaViTAOhIMlB5+xkf4mw1kZZsj8qnjj8k
o67l1Rr0hY4Hr3IaR2KPfW27xhBUCBXHDTz3mx6Va0aPRtHulDrYbu1kTSeZdp3m
uQsW3Z4VpNRkjNoKLgGuZGlnj/RJTTO8LOGH25NnfIwNjJTnuXkY1/9Y0d5r62GE
qXhxPJyn9P7H6PU+ReMaT5IxPpvkjVN14cQasSXNO0jj7ova8Jw2zltBu+yVTOh4
6NTYfz3ujikBOJuy6Aa9bqugkk+ineX3rv8uNTj0SPf40YA8N/xiyHzugK55MyM/
E9hBv9ej628qAQQ6No4UhtUzNcjdM0mZ4dKSotAUMyNzafGF8Q98+el13GDu3a4R
D3EIrvgfFCjld7pfa73CPDqvvgcZPikyN87fgiOfgUjZtO056fDHPiphaAVVEfjr
GVA9yzYho53sm2uFu0nzST5txrLEvRATOw0c01JFXQsdPFxblyMo0hliyjuRQXtp
/FbS8w5VDXz64Ua83lYgMYxeW5ER5iixxL3xlb1B0CZpKtbKBhYjn90J/kGnXXsA
rggSq5L/kiMyBuYcNqEKxBcQH9ZMujbKbo5oExFvjBunmmaeyXYzhH5EJGDc2eWh
CTT+RfuqAitoA+hdWAC4GrS4GuOfZOpD5oPXNoxxmuRKQb9+GIVkqPPV68YciIUY
3vaFXnsFiPFFg13YHJ3B5c7VvRbiyWuMXGa0E7wTagfTGo61xBqfSWHPOfoWvUwe
7ZWHiMvcmdcnd+0og6RAaCW6gya/uQO9ybqGz9nae7C/o2OhpQ+OQc3IP/NXKutF
CTP1RP4YVx47fD9PgbNnnAYiRfbzIrmZenwVBhS6K41jK7K/GyV2QoE6wLcBqx5k
mDDgS0+7GnWqgPVDqvAdZ0OUBEVlYo/LRTgTSom5MfVN90BrJOAwgdlJbpst7Mip
gRaf+OfRxtjq9ikQwQvaJrajt30K3Rmp+zr7l+z8/n2MRK/Wak01eNmWkhejnxG1
9o4TLkn8ROesTmIMpL+k6gFZ69RoBb2ZiJnOlyoBfu7IFfthMFvOcrsnsQOFEC5d
`protect END_PROTECTED
