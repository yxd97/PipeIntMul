`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFjjio9pbOSQ1rYAAUlZh2qGLYikBDzI1G7U9PYb1Ea89utWrnDJLH/tE9Xpue5b
P4yTDEaSdS3y4EV19R8O8yEbxKE2kFK5F11RG1VyW+zzzolFGnoERibXQxumms5+
KVrfw7VPTF0pS79x/gfV9/K0DDAK6SkExrAxbbShV5ejrAdZUyFJtGnuAilfffCs
9pNhtznKQHQqAVzydEr2BlWsG9Xha5zz8CMKAUPy0z3qqq8a6MOc7hVJ5dzNvOYL
LoEwcGwuqLO23xBxVoBgBjHC27RrJAhod81Mr9oCyNm4AfDwDk8Hl/cdJ7JDZhhB
4/ROQFZOG5Uker+6QqDwGC+6aK5XPjJ0PVBoLxuX3pIKJWZfzRQT2GWXUNsmoKvr
P51tkYoGEukseJgQfZu/gTDrPJmXr33l+BhW49HMe7YmOBcIvFCCJm8BPqVx+HlK
cY3NDnqP4M1zRso/u6EL7p8eweX2G2VAW2Mm/9JIMJMFsjy0DSb67gl8LSQpHJfH
8XWsCsLvwXFmp/HxZjDt+yF5fS7HDm2pMGUV+GCgzG6L25P8uEr5AkqRmsjdY2Lu
du9hdhOP/sq7DHf5zNhM+ZYFgowWjsJv6AW3wMqphYYq1F2wS2G5EgAr64f3eTo7
9bxlfPOdSIZVE8Nih65zbKC/c253xKSaDJJFPTbRnbJdgTtaRBH/xMZYjdSzbVLa
199lM4DLjIEP4lpjTOVggv+HzDorVisDB0ZRoDUQX7g0HlSKkTrTIxAJgkK3fbhD
rj6+8c3VSpctsxb58OgstWQhh/9fCkdULeW25jRHEH6mjGsEf+m2pt5X+wTDjqq4
3cnMdWb5Mo53NReLkr5KpdEwDZ6cBhBaVDcd9AA+HXH/dsACmZjSF1RsKZJED+wE
FadbvrVgjDQhjp9YV0NtbN8USLPAIhMRtTtpS0mkl4t9P/ClbqaQ1hUMBKHfQR0e
rucFY+wa92Gz3XH8vMzUPw44QhXXy1dlbgWIu3tkdiUygls7iEhL9kvS6kNJYyVZ
A7Xbz2ZwvXPOViY+HJUaAqANVB8sdFvREl5OYt/T/iDhBRSgYRwNg9RLfQSPTU90
ZGzd5BI6xfqbladr1c6Tm1WYC5wRHjry2GknHQn5TMgvRZd5rGWcYtGwBlxq2MKI
JnSYUs5CZZDDQZTO7xpIxaN1JYFgS2VhIlx+AoDRPI+HmPLtQpN/uGK30M0SCZCR
3d94rwjc0ujgesIWD9hFHNonacmcE3SqjHETC1vn4bwiTcKyy+4wv3wRE5q0iBeM
u+G7rIxTLWBgycz6v7ify3ajj8rWWHhSG3GNyPxfQqkuo8AKS4CYlJ5qGq7e37dt
SblFnK1MdEGzTVDvsbxEP11adHvV1XmbjF8d1UR2qkYSCpvwHVbVKQDeGAxSn7VT
o46S7XnL8G/HdRhe6XDbOn8bHO1LTLONOp9qXQQIKHnXUfXOgakbgPvtrhnixR5s
i8nuRKgsoj5+a2oFU2HBOE5+s/QQrwQH+LGn2g4lUcftzudLvM8CufjCECT/5OTs
rijIAA2NZ6MR+EChBS/t7DF+NTMv3QYT51z7iYDZYXGFajz0zINhSxXx7DPPXbjl
vMMWmmWTRsq8/2H5KMEH0qOKXBcemjZ/tbfqgPduGCVzCRFCUC1cLptekEEUy6LZ
bgehaygDSz/AskCiJpmSpACsgW9sJKy96boNyJ9OpTNJUd1FbPFSomg3q4nX0T4Q
GKhmwPt2x8YXayKqFB6KFOpX5wg3AtqD3eisDNW4ZHaAnRLs+Yk9SwDGHtMBpe6s
wgYkZUtxf0Z3BM1mHANU17isREzgTrXmG6d4kteuSzj7ZxXOksZxuJXt4ZXKgiCd
UBFlyrFvMcoKJgh7gUT0aHtB2LWidmClRtMFsVSOeznEg3TGjafa0yYlJ8vxH+dZ
cFAPUcRcScKjRXb4ZgKbTufQ0jsKP8RixyxFVtkc4jrIGMLxEEa3oyset8TASL/b
Ywk+8V3gt6YQOuGUlJAoMOAvVIuVLcQ91+xbYRy7ixjsNQLHbfcY9fd38QYSa6Gu
xv+BxMVmYrvo2EDUbfmeC5yVwU+/m/ss88Mcv++FszDdX/ZF0giCOB1E4/d/2IHF
YlNFOi4kYTUwlMyHAywQPxV6R+qLSLL6pkqI0kuywMjt36w6mWH8tK+Oa/VpTEML
dw3kBpx8CJ0KJYsmAg+6OHNRHStCuq3FVQOwPeNBtt+DJjNVUqxEC/lCTeJTSKcj
/nx7+RqPKGmWvZurkEXARkI+plzqfSW4tqOUGOykrXp8JDo8jzA3NiYyf9paRfjd
oSnuZje8Zmk9txW2VvdSNMkxAth+YhwP+h83WWqHTDVKGTb0kB1qQWwuzk5PkuGR
lLbQG4jHlpQ+1FdFsScAgn888oo9V21dsHrFF1zwzvKDCZpdZtW5i3E1V+QgpGOb
8BsmlOC9e5gRWxeumxuqmz+4FQAtu6FoOf2CQwI24r+GMff/kG7griI1PDo7EmOy
OIOynoSubBQRWeI6n1FXcxorhVHIF8oRt4g9nGNhNUt5X/NFL9YHduNORCujaQGf
edwpKqXYO9PxYnFF+vsQWqk/zpHQZNYSCoXGRUroQ5jGqxzme9NQBMhGZwwlAL69
c4kF+09PYRG6knyPf1QfWzkKHbIu4rWUCLVqJyrQVVTqFBQYOOjMTAPT8+yJkR5c
sJqZ8PA77CAeHhOxIDTSxceU2fWaplS6Nw1U4RwwP51+KSnGkgSnWfodXgyCNaXT
+vq5zOh0JTVakw0uyC/vNYeBh4KRpcupqJvnNuFCZ9kctY0HNk7xeXNug6b9NgVo
P1TFNwzia23JTmwbrVcW8D6MCt1KkpVxxQ/DY8ovYDoe4fGErRvbvabrE47+I94V
gpVBBck1W993OWu7wesEA8g5bRt4LxdkuxXcaRoejw7/CqXKAUc/3VLl/PGqt/K4
jaBx9mCxCcSgN8A/6re6KovBxKVz+qS+L3G6eAxR9A4IdrVbltR4bPqjp2F2lrKn
qYjXnw/AnoOiU0xRpA/mNA16HIjMHptslY9GO3jbzZUgqtF93XTgIkiDbv79leaz
JBafQlNWN24duTCTJdYxJjlSUtFkZcVX1jLTXGNNYRY6ytQQlkd60AU6/T914xiS
lf+1iEziAeUIi+gkndOwfcHWaiTHxF7QvT53x+JSV0WiRZAM34NpZw38q7CmUDfi
Ea6dHdZj3PoWAyBYGC06su/+XOR/gCXeXh0atoz5VY0Z5fmujXxwixdD82iHffK+
XIZ5Nx+k3LVeMrzJ1OV+PBGzFgCUptBJOGFfkBFAsdy6N9uNkiAgn2PUvaUm/2sy
fGsmA8uB1qq3NaYSbijB7NQlu2XqhicX7TJWoXaD5aIM8vfqSB5LwXRm6icEIpIk
Y5ud1CasKG2vay9YlUJx+YW88RrqZspyp7GN0NapDKvcI5M85vn8YI5M5jrf32Ff
1LKZg0X7RN/ElDbWDPIadRHCHmalgQATskG+GaqvyMfaAfB+GYkVotq0Ig8RKvYk
fCbOkQzSKIuWI8kRuRXfjmfE6hpoZ2XbMKk7Kg6gYVcJI8yGZOvepiP4ydhetKaC
/kWL/T43qj6ZhWjuu/cOuBdvhByLnZHmQKwjaL69d8oPuUnvLFhcG05e59k1ZZZB
iblEUqDCk4uABPu8v9yI86bVvFgk09xxWPdKUK4HZMQyx7BqT1UxzJRRJJsdDCDm
qsIKqv/IidBuharsS9CEixTNoudo0Y7FOfK/1IgiCn1h018w6xxFgSHx0fVuOR1k
4lJaNvI/KhHCd8cuWJmwlPvmB/irsoLKwkaIFOJ4neoe7LsvchTyixMEtvdGSxJP
C5NHI6Koy09Qk1zaC7etDHU3UJx2lurQtGQF/zbNfbfcEupNKPCNEH4d10g6MaEK
90p8rIm4C0CT6ULI56UTy7MXQUs+pZk9ZM3W1rv8CLhG56kVNBiZ8oecj6KmnDct
sjh1pKV+8kjX+8S8DKf4a2dkaZAqEvTbyMIsUgnX75GCP7Qz/hsoOCawkTn92e6/
dfOtNFPruUIkAmdjJcX3ZXyxJOu5ogCREL26tZXAZev/LekxRNdoFMq5FMOPfb1r
gdzmslR2Rxg3QV8DEG7R2htP+bFBwATQt53gF4864YEVP326MtL1iSq4c4XyoJR4
meGyaFA47gT+rmkAR67prMr/hMDlj3spDYtkV2aQiip/Lsni4MOv6GEGvoOLdy73
VpH9zG6/LBKQkFMNWS2zti5XFgYY1hXlFXJWLHu6DIjMPfa3QigeXhyvZd2TNJ6r
bdzGjvg0Qm/T50EPcg0KuWg2F+h3fVz4skDAwQmZBtyrSWfylFxqp/HgQaVFyoHY
AMAuqL2Iak7KOGElBzFBTDQdN1WKipd77PXOfy7DGcwJAiGIkl5GhbbX93yyt9Sa
x2F6ayux50XF55uhjUnTlOqj/iAvCXAp7GXqeMcNDIHHDTF2IGVFNwyp8D/N7aaI
yeB5JVmQzfkLRPNDSFbD0axYdgtDaQ/1ttwLdXLbmcNkKZdVbhj3TOiONRXxoZ2I
rL/P2mwDCIHuLus6+Dv5msuzR+9rOjtCT+SxxMMIZo3vuwcRlzqAhCRvH/L+BpRC
nyqSRUiri5mxZbCT+82LAZNCMtHR4a9vrvrht9zBEUUFxZlkE5PDCj0DkGIt+FUa
afNccBFs/OmFYiEeKgradaI/IbH8ru1XGwiwCkTTJRn/EZ6w7nPyrzlz61ltlhsd
Im24S+49KmB3wNChsdW2P5rJ2aiAjdP+fcgmLX4TAvP674ePhcv0tx+Ii7SfTRy4
szRsXO6MfL85/mlOSYWyHzeSFrmVvlUEGmFlVSXl2OIIW624FBMq8S65m91CXQu/
wXJ+2Sc8//I8YkIt9BtFn0Jk2zjRxMGiUYb5i/z4F5UwJt8wqXb0TNeytr4Xtx4Q
VGXTDsKCDlFkAvbmpd9DaxFUNGAOysARkhbRvZ+LWhX/E8wZ+C//DfjBrDaBc+FB
zyjat1GZlt2pLFZdrz1mxlu/h25vNgXZ0EKeTNLQzk2opgV90/Fq3Zt2ZQdn5zFt
XrN0swTDaLKUkbNV3Ubz5Ub+gO3JZRwumk2q4ejkBv18F8FiDaFmo6Ul+cQs52rE
A3tFSL6VyMgyIwOz+n4Mt0G6o+z+8gvCFfTIMT89uYpldG+8bWmWl37juxGQduY1
5F5WyYPq8gjMCmZeVX8jzKWiHHI5+ZmWifK7DR9nwVpA2df2Iabw7JcofGeZ6G/p
AbqLxLfcdnu312hyXsBHvORI09TwoBHkkms+JaCOaz5qlIsVCuKzbecW53IGWkLb
Yiwd93cuYzCvzT/JnplJfMIzYpM5yEz38eKju0yiNHYmk2qyycy4qHghdSBh4P2S
rw58hZjhCge5JQYBS2qSqNq+TerkLXTQV2FhiIk9BPIxfs8ZP9GunXBDLyy1uL7l
JlSj59nGwmI1cbjBG4NXM0DDQ5mp0Xa9w7HWPpiBLGibr3QEkEDWzHc8BmZ3SBNK
mpKFqi/JudTMpMRJfeo1FsnS3B2vGAKDHpfYo0WaL1sd2/DqchrQmCVmh+CFPmkQ
2UCFxndoPt8MC5PPv24It9S9QLUgIZBdvmHUT9jZ0kmUGli8uPlRVlGYuR60yHzn
MQmTRlQXrREpSRuEDD1praX1TrQG34UXirLUr8VupBFXVr9re9Akt4eEII/lAxeX
B/uX1bjSuCxbipR5NmYghDtq4TVNh3LATA7BnQHY2GNVsQnnEoKzW/hkq89QUfb2
pE88o/a28MdwcmI0dw51EsO5sBBmaM1WTzib+XY8NKsUV3qBS71fBBaz6JKhd9Sx
fWRe02eN0U0Vp27AIx5wgwUii3kml2uZiKb5o+2RMWHL+1aXvb6UtqHrZ+r9xsuI
fCIeeIEdUEH/G4687ramQgpp/Q0Rz9RWLliDMuH3WhFYplL83z9qBDLhbHbLVfj4
uRM8i0KA7+h4R5rLMVzemqhV+YTw+HvRas/8VimzZmNh/HQ65MBbkl1iod6F1aQI
pKA2ramTIc2JPsOMH3Wpc/dv00hma+t6SoG5OApQyTBJqN7yVdvkFea/HBg0gfJX
AJahNZRQSl5xTZlp/KesclagtUvme+ahM3Z8QJrOofT10P9U5rUluf7zhDJM5O6F
RSb8v/3NqEHT1NKK/RlMncbF4MxRKDsBYVLEU8eb68J55lTWvTMbvHSYKe6GBPBh
MsVEICZ7Y5msmD+PcxxeKsXx0iDdIMZ+A6ipO1pXeRyR7vgGIm6iU/HzdmurROgl
/6Xnitw5B/nr69iDCB9BDjqq2l0SKEfoGBCUqzcWz0iH0UIpZ0IFR0QqPiaSxWXP
5Tb5BhnA3VkOM6wipv2PUhVUlbbw2ZtdqTSS9ehiMuG6wPUQ9OJKM+Nu03H2UetX
lmITZUbx1xPskU0DfhUUXgt3QDKNZ2fjy5IQzx5boGLJ2Sf4p8UTRvBSkjyWXsjm
Txg+kBMJMnc2exE70FvhOs+u3G+Ja+u+kTp77FFfUuK6W7NGOgwUZZ+6ux1eHF+s
PKbN3trkjp4NAX1vnhF80tzryvbJcX4DS2rTU9fIpoUzshgNNfvd+dzjimA+Z2Hn
/QfIjZwb0lWhLFi3xpYDkfppEGA8MSa32fi5JsiMHO3fyx4GEtc98PeuWWIkcMj0
g+8AUICU2MQzwei2tu7nN5KClyirCUKpO5GWAumblWYSBgzda77YUxHRtFytrEXC
0SIMzQEim+evJVZuGk0dQrpur4RdvuO/ectqsgMYA0tEToW6+5BFzRhslxLa+n8y
gMVpe4HoTKcyYZJrKIjN2UBn+rRNC/MT/nUVmRemqhA46p3A2F7SBgRnf8NyCbhM
lCU/vRb8hp4EQkjLFHc+1ssL+xPBLXXKSc3eTC6z6H2dDuCVjE4fSPioXzBOr0wj
bfv0SDfL9et5Pd4SZRm+5KzJi7TDkOqFbhHLLswCmj2OZgBvZrIEjItGRga4fkyJ
3AVVqglRf7hHaM2w8eEyAvzvR70QbXUwIxkA7gkMHE1fSqeSIvSLpktlhK60Djab
fiEcvpsjORi9isGeNxCcsYN35+fQE6nwKRlcsFFva2ox69Yn92SO5YgExGsshX4O
wrkOBXEiaWFgXgQCh7Q7buhN58Kq2Jq/oStQHkpc12UF3/MZNHprqGLcvsCmFleW
+4fVg4DPbbGy/Z7U0AQB3tH+QZMk+uZIBwOLGg6rQ/Xhsh3EKkmJ0Bynh7oWH+Gc
TrwONXDVl/1oTSp8r7KuMhIFH1sGJwRGxokYtkvYt6kDIi+4kbhhqjnEu1W50kWZ
7GHVbApWqjd5F4EkunfwXgeJ87Tcyi31YzB/SEyOI46PFattLPqCqgcwdAm8qywZ
2iYmSxj4jV45ZgA1hqAFWLza/2gig9S3Bo35fynMvJsD0nXwVlNh75SEYDEC6Tp3
gXMF4IQwAmlOtZqvQL+fAmlg1qOZ8vnsOcGe2wN+oxk9cgNnyRlLKF/PC7Sv/SpB
/uVPfi7lrIH0CzDiUvVbrIkQYpB4bBVpw+BR8qIexSI8jcWeDNabLZZtGtHXUGqe
+eSfpMukikgFjxnhhP5rRT9inpTgdCjxJRsB9tF/lbrKOtL+FwQe520M1C8vNge7
qiN4p5ZBTZBUhh9mnqX6FqqMiloRyNS6JJnVGoq77BeVoejfh7gToWAsIuqgelXQ
OJKQM4JC9ST6UP709K/wbaub5spcYGf76uNIxD8dmBHUabeBNjlP7m9tu29VpUM1
FP1yrKVTvWznf54fymzLjdRsPdXY3knn1BTUaBAEWaLWSYsvfd/jsOQSRWdAArax
vaZaQ/RApxJoPPt0joXKmOqC0QioH+Gy7KUihS6PQsrGbp55T/GiVh7GdbkkOVEk
Ab1W1AxxOIy0yNKeD6ZKnQAA1bBA/joJJe3UfkICSkr1wKJaFjRxVHWq6UWNehmS
W+OIvNw2DqgW6ru/CUfLgWB39zPpkZPwF5SLDx2AJxoxZKJ4ixcdfVLJ+wyjHRH1
Y9uiuexs4XKjl0abtnhml0AbO8W5+2ElThv1taI2exv1Ffc83d2iEmI93ETBbbXO
a2+PCi6m6scaBEnfKv38pSegXmthral1oNE1uEcddKyWFuBS35jqfiix0Jw2jaa7
hC5Ffed/b4JeGlJosFBzDUC2p+5KXPQwgD/j+GY/hK2/QPLSVwKlOyW1N856cyQF
r8RxelMChyQubPqy9ZtsyjdiJJf3J5fxP6YY9sp2/vMlroP6tV0lYVgwJxjhE5kL
nZXZQxrA+jBPG0U2cMQBY28WX7IkcoZtb7hT8IczLGMJZf6M0Iho7rSpajteW41U
CJJF+c1uexo8n3bcR84vgUGLB9srjFNp/l/yBRiNdaNKtTrzdA0cx5JK1ENKHmnW
JD7Fa981GFLM7OUdRqGx6ce1GNEgZqsZzpJAfZdgzsPZlqzuu/fmhJ0XTkFDEdM+
JBADJNQnxLBtgZ4v2I8xTXJ4UoTQkAkzkCjOpQrs+tOXVRw81lC+WUGLIJLTO78p
8wv3G324ByH1H07D4XoqSfvB2W58RenPgg8PaFKhf1SUJ/RqHFel1mIEVRUPEEpJ
jfBFYXJkloR2Uk4+qMd7E5hwgp0q5rwLCcGnudfPp1CHOXwPYNcFRiHDyKwU1MTq
ln1BuMItlf/a+QmA+KRbh3RXCGGrZPSYDBgMGxehHso5ys8FhXhH8Iay5tLUn+vG
BhVMXQSJdC7TA9Tx5rY+4tXPoew8hoCjA4tDMvbNfIoTtQu8gaqdB5XoO4l14OOG
XkObBo7vS915Wt5BoGc4TKZkLcrlmjhjDQT6yzP3ublKCoVeBjFkyyG95Eag6nLR
eB4CES+2HajTm3oqOzA07Ib0NuOX8N/b1zBzc1oqPQQB9r7QqH4sZ6Qa99XLGbUI
1fOM5ZfS0LUkRaOYCoGm/m9XB8BaxuZSLKqLaEzMQ8fuoEOxos5ja6Cs4XNEYIZe
fC7mgei34BRZduwkGdwvb1m0SNEqyKAHY4PRNh0s2ia2v6n8wMtoO+QQ3A8u/zws
1bpC2FR4bquBkZzeU9qIY/uUrGHWPV5WZCLotEnWsVw/Ex70wNeo+gR6EhysGN6m
XDmBqADxloQcnZK5Fn/9E16l30u25lV7wHunexU1Jz36q6/58N89zq4tTiYV+rJl
2N+gBFwrSjBE8DYAAYZpEUlo8aveBysRWpJ8nFclmqKZIhplHZpB5hoD6H91B9Wc
pRMiswfE+S2zt8ivBwUL6LAE/9PUcUiJ8cU82FyaJ5nNpYBZGNXaNe3lWgJxK2aK
avPV06YGmOgQJYApExlNzurd3XdaipPTuzmj73GyfyaOwaLtK0I0e4uGcnyws7PT
WdTeUcm6dDEuScWtXzCcRiuJzgVV9z5Lw/htRzEIN5N/uthF/Br1px9mGYhQh3Sb
NM8Xv7tlGywc8J+mFJgl1kiasPWXo0yVhWHB2dTBwKT1OjICxdZUGhrPYUgzMZcz
kTjp6146hYLHDd+gqBwqogGiEnt/vKIH4mMY4eP/PxhB4tXIPWGAeFfkL6BBj31S
gy26Iembsl+fvzul8+8lOFl54K4GNs83rPHnm2pCweFkgV50X4ZTQ9W+dx4GSGab
zFUtqa3X+maNt6QxJ2J0w+dmZRgoxcUIz4wK0iptlKm/3kXlpgmbL+RxtK+CFYFy
AllSCdbmmwfA23YPp/DRknUvbxl6ftiIL6PhkhqgwANj7DH+DOeeKPLw+cn6JRjd
7eiM28Osyjw3WP57tJdHW9kHmIauvwd7ELm+oH50P6ONRPRNsYPuu2yMc2WnrWHa
Ok5d+t638RQYangtiCPyHkOVA/ik8FyqpuLcbtypYoJM5u+ZYWTVvvN+KdlukwiL
1S96XYvhf+ipilFNbKWJ5v0Nz2kziMEsGKeiLZoZiKL0g065+OI+ivGXLVKNSlMn
faRLki4irYS1MIrQWOjFqvYyBIGDetu7C+DoW1csCTvz7fyyWSFn5cHEr8L+o5rX
85+myJ1Bron6mGVG0lO0DxaZjAgYK5cz/TJyumAwUqU/VjA0QIOHerl+XueRsCr9
svMBgTLVKXSS3znblT+Y4fpo3+2hCmKr3oziT2kk+bmkxpz+wdr2fCUdNnxCc2xq
AMw5dXDWN5+P99ytTkgi7z+/KFQnOcy6alEYz7SFRgU7YNP7brN5FAnalhEIEvmb
XpYwXpJZVkInK2MEXLNZQL8EfYpuQvOwrKsfBtj82/8Y1ZClZd2sqgYa09uVlDrE
VLBjpMzpGtt891FruaZnhli2KAtg3DDvzps0YjQcph+4HIl8TxYzG2KXN9MhLW7w
LWN0u2TjZKWBDvnF83eW8ogCmoMn1asbb5DlOooD27N2mMmcV0dChPq4b/fgyvKX
T02AE/PKuMjxB+p7dI6rJyXJlsYwH9BSpl61qqj8ut9bDSoRu+KkpUkGnqRr4+PH
W8UYu3pRmyb7w1HtBsoDOHyG0vIpAFAPnIYHUrXQlfuEwuX8W8eafTPro3SlEysc
VMTDpM8KE8EHJVNkoWNgjKkeflBGl8x6R3FN/5YKPhGlrkZ845ch15PwxZVR68wR
XSO+BgdTJCp8oO1BFEZ3RR7sGXn2OSGxX0xlici3TQqgd9qi7FH8EayAIOrbTj5F
/9tNJ3JNbXjUAB0gb+jS4hCzCTPG6Z3icMH9hx3bo5ByeWx4vWLQAFX9vDByOi3f
1tlOcul5JxMpdubwcXran45Rmeyr5NjLqrGYwu8JmJn8Moaoz1oQ09vTMj52/3Gx
8mlRX1M8U6FhYqvMNMErVP6MXy9PPsyQqAyqHsTa6df40sWWdHzdkYx+2mDiaqxN
dO/c6y5pRcXnaS6KrMqb54sbANrlzCqs6o108RzXYsKj13g0HCFpdnzaldiYl5y2
dw3YwQFj4G8ZnrnFJ2xhm9tGMB6Cq0yjI9kUaEYcE9eoyRkPtFP0ZPZuLhPdrWcK
SPYbon4WkSKgzYeRunFs2CVcWh6NF73jmw4cUp6q822HTjpRIMKx7rSc+jDM4fhu
yLrqFFy0Js8k3U+sjB3nn9R6xpOnhxxwgeOlNAbZcg4uTXRW2QzCEPRCzqTWTmSg
LoDWjXh7PNYr4ggTwsYkmxOCgA7zvDUpSan1n83deZYRSWd/VyirIT35uw+ooRdD
WznYNY1l5SqNtOduGY8sx/jpBftsAZOY+9Zib3VJ4N2h37SvCmzO2GrCGKS9cPEj
bvthTLcSVM2LErTXUi0x2lBhnti1CZJSn9a67T34LdxDVCQZ4IP7hfo16gPnJpOA
VI7OPgHuVm4lhNGOd+W0MLbj0s6L4PrCOPrjNH+pAnNhHoqSatgu/vifMeBVHJNn
dTVNUZgnsn8q7pbmhjowuawYmP+gsz0EZFmZNvww4pBOWhFMaXnyQkAoHa0YfmYr
AcwOsD5VSNg5/HNixiW/Qg0akihr/tQuXRzVxksXl6NOSa6E+5fO0nSSCvf+WvIb
nGBGjdF06Sop4YTVpj8ESMWOQteCcf73qma7AG9eSV0Tc43Fu8Y8/cF5aPB25G2c
e8HMS1fexWbNcxC87XLRN1Ga820kp640ytVIPkVy34ziu8FWthWHJ67z7xUjC7dt
ndRpFAUrPTDSURt2FcKmXofvX9dLfckRheJP0SPDwXCHioIA866QwCxFd7FuQrv6
GOSmbclR5Mq7PZFE+30iEUTswKGVsm4YkR+qnrDHe+22zjB+pncYRHiypDYAN924
XxlnxAfc1FpbSbeKIgnt9XeGKiX3bWcJEsrczsRHX9VmK5U9oP9d0UcmRpE8gSt3
5RFdaWO+PCTnGBO/7C0Y5f3pVumQ8r2NjhGN1MehmnlCku4ndi7YGs9uzhC7pYXk
B3jbUS9X4Y8qBb/JkXAtJY74uh2cna3khva2ghAoD/DzV8psdtKyskK4Dr1bbIde
ISd6VOOVhbu4n9S3qMb+2jR1jTAd9gkv61as8MsKOgKeKXil9ydCt6DIO+5fFEPp
Gkz3skuZm/x6VAWzb+NJqkpJ+Uoo0dMWKnaztj5YgDhkIlFMAU1uH/5evQAZ0lbS
cUJ/OeUh7RLGHDnfqDJdj2MzbUAa8NHJ1E2wuk2BDV7W5+OhmZtWW3ahG+6PHtS3
G2ruOJpkmUBskzB/A1+wGM3gIw9BDSbcYl8+vq/XQktqS+4/xhVQBPIPEg2ZxI5z
HdK3CyFgpLhxyjHX2VLyX/z5HbPFBKWKzmehNiDQ67io51cec/eGGfAdmQp64n9P
o1gh3KeJYJBRfFcuM+/I/rBQ465bbFGeDTf4Y6Clxx5O/OEsun57V72A005i0bfB
lZX6lFnCGmmPreBZMmosBH7XFewNON7x+UnlezaaVFfwjrs0TXKU6rKedd15pe0G
K39Q/na650SdU6SzFnGuU07/hQVH9bIy6WT33rpfOfDEghUQ7f76aRHkyZ3GGEZB
r3366rJ+lPZRGLQzTKwJ+8CCiOPmC2G13H1CoBi+F5qWFcbIRzDJM+bFzD/Pe3Kf
ExlAjF3lcD3F0C+BE8MkbH/Yu4tCdZCOoGTlnxaddni6Ce74GT/R3wrC445I90qR
7e0BnWyLDozleJKl+LBIFtk448RAYrUMiSvhu6X8KgttoGfXdFuM0M6YkaCs9pd1
nXzlJvPJ6SYq+I4SxlJkmZPl2IIGbRv5g9UITjDrqYxG5F9ISPiRHytR1X6jBVjF
vb68Pb728lvrZ96gQhuklEFsMP1w88oCZFizCsYOI9LxkfSUo6CGYZzCqWJqSVix
A7v/qNwmEp0To2dsYMb+m6REUAMT/0CVSBvW4budlZwXNMc3duo53kqi7TLLWnMj
jvo1ce5XT9YCguj8A0rPn606DuqEAw3zb8iC5QHEEZ52C93aAvOMyN2f3XaFPYzR
thTz3u77TO2Pz5sDFKwZGQTv+EmmPuqE6pCE2locnQPVycTJg15yBbEMg0hpplQY
hF8z8yuL7HM+/X/WbdwIYdQcOPkVXJpBWCSCyt4JwjAL8shfF5DLym0Mj/kFfLxs
74rgRZtUccB6IGHOsx1Uu9VMKxlnhGm7fljlXXsoYKVKwEMHdqHcPRTjld0vor17
T9Gfxc2HVPvR5hPVvFQbKraBrVMN2VEwgrjRBT30TLwtFiOuQxiVQAnj1QrP84aQ
y5sb3fXXGF8SJ9sRgOyL6KXAMzFG+jWUbii3d9qUuhgIINDfnq5w9UAYxIFsSJ2Z
CsG43JwfSvMOUTSH8gEAOpq9KzXXAvbu7YiR+RJcUwp4YJG6CCLEGO6uxdlzGcqW
WsZmQOJJtD4wmzd0AzgNuhpG+k2Q+EjFngabP8irOgD9MdQwslLFW9JjGByTqtd9
hfd6ftMT4BqcxxECHJ2uMcCBZlQgWJ6UteSPeGGowTys2/5i7CL86NTExnVF+vA3
kf3jlvAIKX2wW93lBCWSptnhveB23GjJ1ih7N9sEP1+iUhD/DBUxmZBQwDmcYV5A
67Nanpz4XocaNuISGkEmihILAtdQYb26g8exxG1sLE2497A2I0hIY2T9hQ3WvNLR
U1PycmqyPhWVoSgUudGZzi+4ZffSnUVdSiiPQyfYj0OBE6hJgRjxz+KnU7WwAtcr
+BgXL4FwL+cdZG10190ATc5/10N18opqbioYqV2T2U28CGkSmkpad6n8QhSiricZ
8HW7z837DHrbRMnBLZFQNbXR4c1x6anDVWAxvut7pAd98FCtvLC0iAt+AJt3uAL6
uklaxzjhnxU5m2+PJb7DJJhBcAx7F+iDg1espySkjuf4iR2gK2LxphjgGPS5ag6p
gBRet6TKGSANZqw39mo7CGSHLawjatPw2y5581W5nuGw/c840w+n/D1xkSwJ88Xy
DBi5vZgVoQtZVvnf7DISxpspyKd2wfe0EgLfu0x9aCkiaj8o57SQn6ynmpVVNn3T
gM2Tk6g2Hisvx9HDf7jEFJ6XEruY6erTgJQq2xTgcTvHYy0o9LGwGoFZ7i7SS0i6
3it4uv7F/mYnmDVJJqo33DIsrPZgMATcHbEjHHkbj1Yj1LqyB464GCeKssEhea9E
mea9lTI0C6+j4S1TgcHnRTZ4cKmDbrWL8YaXs3h+rErnQUlm5jViPm8yYKA2/mPG
YWu1ahy+Ht5MrAQKIY0yrWRhbXrmL7bFoPgHkxHb6ea8cVQfMnQKhltCLZ04eMVZ
kLzT3+iGDsgLAqg1mqXJHGHlmmH1nVkv08I2BgYOxRmVynqwVMuPshBDEDBi8IEP
88mQDmMArnaEkfXxifDFT7RBTHa5v2epMvlaN9oCoDXO3ByXTXSE7wPyfP2/GBA7
LP3PYTV2+zJMObgbpmCPvfdXE4iE0p15UdROBTtsmzwQYiC4zJEktJFTy2gPtPQI
iFKI9sBJYvrGmxly2hrpVG+zPfzFuzTx/nMURqrPSDdtzz3CZzhkAbOlkfbP9CMX
FwShRWO9001PhstSqOphwKBOeFyBeY5nIwbRcmz5RBkRuQ11W98PhScI+R94h0JJ
DgQZZK6+SFZnF0uNNpQZBnZKfDxJF9kVLpxGxkZzNh0i8YUbr76+j0sPcCtXxNML
wbwZHpHjo5X1R7AGMBE4U2rpIyXzPoPMILX03V6Gj4xtb2UwmfnctfAxL8HJs+6x
0N5ExxSc8T3XAuWBOTYGZ88q8fSPeDeYEn7jDfMyWSKcipdl2EWSgNIqLGBK+kKx
qntkyKi9bD7yGrLkT06mvUKuG4f+YS/7AKzdsXuyCHzOInFIxKJjWVUlCenNv3Cq
PGNeOOf4LIuyUpC4apb0W1xN3Z7YopFgIfZKnXnWlpc0/vc43mPR/YgKNQbJtX3Y
a7CxqhZvuPYvIzRIuSVf44SYf+wy1Pxaolyl+heKos73jOcYWcHE0XHgn9hCyIU6
Vnnlm6oTRbLI3X1O0Nkoip/MIp0FOU8y8E3Tn5aPmFzaiqKPlmKVJb/Dv+COzoMO
4l6IIzc5o89Hwt6xFfhkLHrPooVwAZXEy6UwCZw7pS89f7jyjhxH/LmNroiw6y7J
gwPpHrKNK0MWk3zS+fv+9gdeKGMQ8UrWxBXaJONDDHnw3qH/BBrRZFgr8d1zCNkM
vfgoMQ3fXzJbxDLiWxHkn0pHURgoud1hZ2Q4vx7TresUPwhBe291l7mWu9R8j7fU
60rp9DxE0u5N6eo+yzXRIHxMwgz5UyqNXVaU3f2hG2/1v1FoUHaS7oKr8zS7RVXr
s9KKGSUg6zUxeoakmAc5MhPZc71BGzeeyeIn6LMXbXYoI9YKjWfrmolBueOguMgb
c0q/tjUYjgCJHqyreuTlBbxM5/o/5IsOhQpwG8FbHKmFGs7ihQSbeD17lJjwHycF
7gIC66nb0fp+cGtBm9tzi6x2rZrh19tjF2IXr8BgWdY7oy2C4X6jE3Jj57QxiYMi
yMAuqlCnHo28CdRnCua8dufphCyFl/9bMUM6t0A/TkyQZuIJcN6Amkxi842c9dEC
nqrfyd4QiB/TdLrd5mljA+tJ4+v7hobbPyrV+cRbtx2ufhSyA3WSERNslL0DuQZ1
X8xt1OpAif2ZXzmigFg9wPkkCxr2Yuz7V1h5BXyAhvcb4Wyd/S6By6RELffxgXZT
f+qxBlS28sz8txnmpFgrJs5rnLswhck+abocVFSQqcTMGEKVotwYyvdyLaCXdP0i
e847RIC/5BFVS2sn6y6WL5xieBU82Ea1oSZlCHh4JTEGeyy4ME65R2txXQpXlBmU
3VQ3AMgwoNHxHn1awWgHyMq/xE2QT5dDbIQsYIbg0r21NhuHoHxM1Q/G3NfPQVv/
XDx+GOA3Ry+bd3bSqO5YUQHg4xl/fVywgBW7wS0xL8mMJundNmYOY5qdb3rKfdg/
vX3foqJDltRj8JHN2QF8EOJdUNdadwt6sS38LFuM2uPfvNKVEzXdUf2rDuAqEXsl
syIWfLc0SHQpVu4/rN06X1tpf3Dby1YnuJz4jrsPk/UGFXnULOwY9gmpPP78nKSU
f/TWQ3mEsEf5qRGkDGUI62Aq04nqXe8RGuTTWEhzdIgR8j3/lE78dBpqrWqhhHRv
5RO7ToE8CR+BQt4BbyRgIka8rqPcJXxJWd3KJJ3VsPjlreL5gdTvQtlunVGBEJuf
LIPkstIRDtYuyQUkKiq18Xq/o0esOxndyR4QzKAw/oqz8pZoyHkrkyRaMsU4JliI
pyfuqPAAH8YZz8mojxb/DV/ZzgxQj72KOY05r4Vq2oyM3IcxiKAUmhZd00iiM05X
qGx87WFoaiJqbx1OAqpogjJhjbjRnk0mhKHdWRC2NOSsEYk4OsJbFRzNsHFj709I
+uDPErEB7ZethYmNV2ectDyWPTph9Uq8W87Tx3nuLULZ6usz6nyqeGRL/mmR8sGh
rFlhrqeYbi7dypoNl6w/QqSVewkKuab1zbEN8LIVlShTYYiMtCNNGY8lAtO/gfc6
ewKqa+vMoT+cC3ATGGpwihvcjWL3Z0DmGM1NL4uw2hvU0cljP9B7uzC28k+pgIud
DbxCzFaoQ2qGC2X0mM8H4Y+98CEut5YjuB+MzJXr9JOBuAT0CwhVdejy15YUTCcs
juI17LDUqnKbD66jbJvfGVXEePJJbx6sfI5TMYlc5rXM7HZisTge8gjy6UdhQQfu
/BOX2m0vYlWMGMXeI7gz4ftyTVXe9drgc+NDg4G4ZMeg0K6OCTvLgORGbepouRpG
9cSu4YlUn5WBVpWmrbdaGo4wH0pQMkXEC7qmP2Qc74Wb9Gk6t08c0Sb/WR5kgWRY
Ry000c/1HQ+X8OdboVTHztaJA44ftYC/oPa1uxouO8aMcN/FcCHv/Mq7UlVNd5V6
uNv903MZWIrmfglhieQJK5OXv+YXjFwV6w7z+oba2dKz13QZXXUB3ZuR0PqtgRZj
zuRa17psLYb25y5bqS8bI8mzijp5QeT+WC328oDgfEcqOD1RPJv8HRdu+Ec/rePv
hHk226FtoCiXSbeuHAfd+oLyx3SRsVhnBJWdJFx/3zpr/KKKSoX9booIca0VToGy
EbZ+LqEzLTdkCHQkxyVlZequovZhcoy1Odbpy7sypT3edtBsz+1A97+t3i9pBtJx
T4TnsuWzbJNEamoz2nNRe2kP5u5dmiGhzphM7pdib3fY21Wxp3d9a4YFJ6QIZ5Ao
IaYpNekUTaw9CCPSZNsTGhpf0o862ImOZae2ySN1PJO8zSqdLMTgQt5waXOuktec
jar3Cl+MwXl+TCvE4sbrwsVIlyUJcAZl5G3pyg0dIb0ow75hsTO6VSTI8/U1ntwM
pFA1JQyr7looty4WX04PZjhiQsQnYpd2b/qJz4Cy2xyVkw+0Nk3jO92bkZCh9nnL
vhFCRZZyvJMesgnRGGuecGN84ifW1CM7tdNTnzooF3Q7xnwxQrxe1CljRQCoMu7/
vOBt6d9LHQvvco78ryry6C8lNjjRO+d5IAW+4tmSRzU93Tictxe/zucwcPbkiCUe
WwBFMKAMVrX77kQdWcGyuPDfnfUZJ4U0At8gmtjBuL9MYhLmo+mEW5FWj/MruKrs
2Kh32Ay65erWydSgmUjLuW7SNlrzjQJ/2jKgfmB/vlb0WuDWbeNpE9SxuBv8oniO
tyZ19pQyduklTX5MZ8S3jB8N9Dm1JUc2reWGkeZkFSBUPDd375tU89qx/8fYFpy2
Xv8QID0efdbeWda4pPUr6KRNAeaxvFX78otpHbJjQTacoF4cPHRv+2UnGjlyAB31
+cVhSJEoO08tu4NEOgv7nSd6Xkch7J1qkDjfKEsIdjaLaMf7/6s+hj3kmO+rTgMr
nEXDww7Lp90dt1oqKW8l+w==
`protect END_PROTECTED
