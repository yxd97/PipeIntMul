`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuzuhLiEYkk4ppr8/BtssCf/1kBC5MzFuO/4ATP+AoQrnirnQ73Z8mDQ4tMm+i5r
HC3uKzvIhqY+X7lKdYFeLUWwZDnhtLahzUjYxnsWd0kmeL9ddh12mwmjkIJLaTiV
3AY3WlmCDb7XJdQq/UjiVc5kJwkb7kyjeozZjIhzpCr4Y3ESmOqAvBHUeLH4k4mu
vsoxIGfV9yuyDYmxU1FrcYUsYTvk7M/kx0kzxcyickEfnk5UJv+mWyk+U+2QQFqv
0LhdpG3nK08YqMFRBEDsdBHVJNZMZT/how6yJSnRFqzwWMuPOOBqNY89REWQXVh+
3U7YjnfLHmaJZPveH1GsDAM0idIhX+bzuCZH7+WCaqTMAhDFXP/SP6ElNaR2trw8
UXucvlacnP+To6c921E4QbeOg8cEH2leHOlLActGfMTozeizoZb3hr5A/bLkNmnj
MFZztTkK05TXUU67tec7gDtMvx9ZSgSYM7tB37knJS9Nu8JuGNu5xNnc8+fjN2yY
AbpSkxvrNqZFPGDSxjbDj9JFuhcQaRlL6GE8nFSkdSt4oEr9wAI7MpFX+L+of/Gb
ExuYA7XZXrgIlNP9nEZk/rtSEIUohzUvArk2HWgsZXw1sJLykGRKSkaX2MPbGCc2
etlsV0uNMVjQOALZMOgR45+sVTTfrejN9RZN5CC+GttTxYIj41ajBQM4W1yfJ008
OAn8UeqM0F5N24uidpRFYyd0bS8l3ugFaaHzzaomE2HHp0OExfOciRR9GVFzYL7e
59nxAq0yPxh0oSazht8Yci650elxd4g4H2rgtiowJhiVxaTa6+7SGFe3mRTdIO7V
s8Th+FWiYLIOuIDm+htXJgbgkczI9ERQntn/++9sFo10F7h+Arlf6EqSNPP6Tc42
WA9khh1MfQT9xqfAVs0TnSlLHHtQEmbzbbwCGIuk6VRjtLb6g12bDK2FfpvygJGW
ZdF3ludjHCuLwk1YJr9jp5EBb3TgU9ihDyeIEOKT3U1ixb+Xv4kKVH7e/zNCcmD5
3rXWOGoPkYuVxpwQM+iKE9F8U/rcNFm6beHPyBDeuvbWpY14WXf7xL2kS+iDI5o6
5GZjo73Dw6RHu7ObUUQLypuWFtnUBgTUya4N5itwiIJmfCrAnucsOzMcxs8ljpd8
po3LRXEdIfLvYxO4FBYtsXW96hZ4OdM+g7V1ObmayHJO0vVUpj234ZJiylHpIYe1
SBG8AtMsPDC3glBpxoH2p5bY6bn+78CT6zTe2V1atME+EddDUBxgmmJMZupXFqOz
UHOE6B37t19EU0z3BHYnRotl7yIoZKf8X0y+stOMolu/NefskU75jS0C1b/ckXqP
6wa8GtoXEAt3S6EDRHc9kWK76yRCDTrjMPJzVWhayqwgaIqrzdjHq1c7zYRLyKNq
VYuurN6tlAKLBjKr60CNw/niOA7QBSmi6deMgxaoP54Qqh1GLCuvK1cJxHyVdCmM
SDo7Tyh93gb0dgDtBzrVYMY9PcQ0tjfAIGJ6hM45i32EQ7WWkfwJ5He2ahfoc7k1
JCNpVN6DhbUy1OpX9xM3p5S3ofEoZr9r6OTRpF0DrfyV5E/KaNqfEH68tHaGqMZ9
Z0Ag4EH+1PUh3H6iLpKmrTXTWnBeVlPTBn1sd5Tvzo7R85qdRZMXNss43574ux1I
NwaOAI0uaVYJcEEDiUX4xbAp5ouAFxo3IFI/cXLguaYVeJ91LWZGwEIboo/rUYXW
TmqdIEx28jDyBvyjnMni6LQJynPAq2tO/7ihQVjEJuNdcqgpp/UMWk6FvZmGq5Xk
tdurmdMsQMkJOwMymTskoUEJEdEoMyjIB1AioNgvxFr2iNRyPCFE//fzUu2pxdBg
rU2nkfzWEpMUgV/PEN76BMxHopd4dRumdQz2ZLlqj+9CCAGzTNtzX4UJwm9VTHZx
EVqTPHBoWNp4RAim8aewRTOZMqODdO4mJg+RuJQWyR3naf8bX36cHBGRkU+L53zB
v7jXy2a8gIpUAjnUFRrBAUeH9roz3ssbuTb9F6L9LXSKrjmfFNMZgFkwPwrM1azt
nnBq2shPJwfD09k+ebUCCAJYEJMpcT4Qkm57XL3m0cgZEmRfteWXMXJKnOuAZ5RA
DiuJ2E9ZEo5HBUWR5ICcheU0kLrC+UMNWG9EkRLtxCa8kNLE3z7AA6ySmpUWe9GF
xZtztaZL4yYKt/firfQA8tfK/KM9B+miCwi62twCSjF73GHh9Sm7rTcTy6BNKSgh
k2XLHCVm4jDDrBkR+VrfrlndMh5V92NkQANUqqyRtE9JUlBXmP4/r7xbbMk4FRsS
1GiqJVKPbLmERCY5JO2GuGkTqrhcwa092iQ710BZrhngA0jnarRICqsmzhsODbpH
1MIM/5P0CdCO7okwoUcvHCeCY/jwOnNr2uqHDRMhTh8qH0vOaqa/Nsw1YerQdUND
wrG9Ol9OrQTF97FIWeCLFzOi9ghI44XrqckcVmpTU20KNwlg7rrm/vERTaPzYaJ1
6Yb1kA5BvkE9SwN2w0fpNlUNTcteP266DsXU2jlbgvgH2D28ytvPaU/he9k7jX/3
eH2jFu/yzzV/vqVhIButo2rQk+5639nOCw7Tu4+vHXDcINIcJ2Ah9FmMROfZPkHg
gEtJAwuEl2RgLggpNn57tQIA8a3pH+u+nmT+73NW3mW7Xrw6R+ESs6eMLka5rrD2
o01bsRXaax+Zt0vAxd17wUzXxVin3t5gmJ1CwcWaml9jEzhxWHLOK3IPMUSCJnGe
LdctDLwD8bDaBPo5CsmYMUkdxM10WxrR//TBwrufwvy+PCtVqW4SdfCAPOZwibsA
D5pVyDMBf3sDkCFImNy2l8++X7Y4p0DSXOwwf4zUI7Osx0XvH+Z0LoOU5rUBIFAh
eAYIVUVBlMWIdJNf9qCKckOjMrxWTNrR8DwQ7FwAyi5aWNdZ29N8uiAPJxL5OHzf
NlHnzPWGJGjdMCZekcH2EHYVim3ZFEH6d6wfsKwLBouEfR2uIW9ASBHU8QnhLo3V
PE3ILnq9cB8zCAdhDpD5y/hFEv3Yl0Y/bJkDQQ1Iih+pKWNnIUzaOUwlXJEsY0vE
/ml8w12un5PT/QktbmqS/yHfkGxpzLS08Xvm13hpPTF9goPCKWsw8zVhcrgMW2Rz
Pq17fbA5Bh58rGH65l7Giqe72vLvoVN8pbNZcys6uw6HKLjaQN9IP4zVSB7/1lTe
cA0lRNkKG9yVr0mX8WdLMjoC/bpwOTv8/JSU0GkJNka9P+e8bEft+RL2tR/ljGO1
IOyjb99VfRpiNE++LJ3M9EagJXABwlCimlbuPoLwYEhBZjZJFoZqtTu9dX2x8Sf7
9/Rvv/bRILdPo/dkFgH80+llLQuOVa7/OkOopvsckbdQ5pWjqmxOjtPcxSgpLWAF
qCV+NH++xKJuGS9cb4ouD9x6wOfECKd1IfV8oUrjvhBZcbUgSHZPWpyi8NzhNvZp
xmQQyim1/xreoP5bxJipk+O4S+OGCQYhrb713AETQlnMrjHDZiR7D7XA8MCy9eLF
qvER+BD5JuJTgdF289dAYKE2I4faYi5T3buztKmFPfHDAMqyL3kPhBNxVo+TgyQf
sgAFj4FO53AwbVtnB0AVMQhMNRusTpSCyI2jm8xiTIEXpSev21bgeq42haQFc07i
ukKAlnsqrPBGwSXmZMpTtb4DJMU3GZ2iAy/w4PevZMwZ7fJiFrStRx4OavNcieI0
P9vFaAyiJMP8VyAl2Z4LUHHKk1QjfTBINHII6V+YdRSUrz/n3sjKfqHLItsU4e/C
PWjheEscl1rF1IA+j3v16mB7OduCBih2/S7G0CwyEFBLP9smTsT63PGW9Uru1hAb
bQtfqO8Bk+uiEPSCxhrTn5kPtxCsLI3eSEXtma2Y4Ulz3eno0wAYzONjP5KMJk97
rfCbeYOIdLrqGqcSUP/a4FB5RG9U7hy3p3/3I2BfgtAWeIkXqIB5Qz+z0kBlfexV
+4f9c5ufd0aGUY8YlFhT2jBqj2W2Ljht4g2UZQYf5A/avMedxY4Fwxz4I90Oe1kO
ClEVBD5dPLBcLjOQ47B5lD0vthW6XvoEgVocO7Q8TW32bosIX+e3/h6QplecK5od
LjD52Ja3TMtaslxjskJSsiUDKUUt772H2Cai2jgSYPSO/P0FIRxFxjUIiJz7vIJW
g6dlo1qz6WlDYBLazVHt9mIPlVDvhlEbEb8iiy75HouZAtDT09yv1K+CWcO/n9y3
VGPFZXwc57oPkT4Jk7mvUlii1pRGuNYrIY1sT5WhQvdZ2zvwL2IOyYQzxL+tXYOk
iqtayRb5dU+JljZmKDbDOr5LESG5yexWTg38eiy2y/a3ysJMk2vtkbFxerpaNDi/
DHqT6EVr4Al5VKaZvfezZ+MZ0gw+hbZyjQK8AbUBBJDK3mqJF+7ZKGzgTKDEasAC
L641n7+Q/+wx0c8WlFxZCbQCUAOM9K9E2qd42W8n2DpH4oM1r02v7Zrc72gyldtn
mHqpIg/7ulSYhrU2nb//tCpkpq51IguMdfeZ04BflRs8fyaih/9WuBOna+CX6X26
7tJF+MC1Muh2Cbms083ms/yTEQU7rydy2wIa4IvYEc0u12gjTNfI1IilHYg3O+t4
dSgTJrjjc7qCNSn/jz+89wy89FwJj3xteGnpZ8xQ57rCXSD0/JvXmTowNFIhcDyf
n59vq3Cm80Tq4rBgxj7GepdUgrCsKdU7RTzQuTIXickyn+MY4dlguC4+dqxvbAcU
3elvbSZkgaSbmLeVyiCT2qUzyRI1zG2HHp2PgodQuk5udK4AHjcPcIDfOpiscvev
ZmM92vlO+kun6xQu7Fh5Npbxr4IGAe5OCWDic6rx9a3pdiQY3DQksbGNzbIphY+A
C3RLXhKFygFzkzL9L3ROzumlHwoo93l3R8VVFdO6vSb4CuISuA03in2/KQu8qZIT
MehmYqm/yWEEc9qPv6PbQGoxPkW5bNkKfQcRhRjZBeDN1qXGsT6VoLHw93GzxcMZ
YIICuzDerq0y7FTFns2tQwH2/fOp5awZsZs4/i2WAOpwDNFwkTvSx00dkUAJCO1z
KrwntN3xXFvLhrnumxap4YKZMe5xh7G0vnSlC6Krbilzggbw1rpb2vFQn5UFTWU7
X1mlAt8QKc394IRn7MSt+hm1vbco/pnuUXCR/d2siwXFxzwlzYUjbMuibIjdsgqO
0HElV54uOZG7eBG8MBWbafp0K2bFUFi1gpaNBU00RPOAQfVHdHTJGhxC8eMaOZK3
fxK779ukB2ZzJL46dYYXBz+ZWQWmnoNQ7KeX+8/pwquKIqzgaMO33k5HvQCyv5by
cnMFrlAgXPCYw6IiKOuR52g8EW9kY6apSDIE50mC12ExPjoZyd5qcV+k6LpTqg9E
QVdn8yOS76alrZa3ao2KaMOyTV0Yppwn9y3yxUQuPDc7scS6kFc93rYOXn579xBZ
3TBFquh+jZdW6OeiDnYJOl8/ryafY3HkxOe7QUHbWFgZ33JLnxHuj9k22HFJ7liV
XgcuEAdTY32VMZdFNr85GV3DmJZc8A63oDrEQjo/kwQiiWAbSS6Rb2bYDt7J9DHl
LfAca/Ir7NPiOEx10FS2bez7hcE2VPGyIhFRi6JY7TfzLGm3Xp6J1GAtMjNf06Tm
raCBoSTuFhnN9sCm999jlgxvfn0TiBtU2k75ZnJvA8D+U5QSVmQ09wbRAAyMQYfI
HtWZzJu6Ab2dRnCuciG6rZUK0440hqdD40St4ohe53dG7gI/tTl8PBcf6ZxnNw0+
uHF6qWmTR+YFQynelOzAJjk9Fr92oOWFrNoCwxui1Iyn6lO7lQkL8MXiceXvciYH
WQ/AHnpvsM7xoP/DbbLxHgBW6qMMXdO61Lt/t3tCwnZRHXCtaea4cm6SCE8DMrP5
V7rqUQBxdwRZz7dHW0wdAdQ/cw1eoU8KMtwCR61DqaEqzoFRbjKr1tpPlAtrxImD
fj1XN6+dvHpoiUnrxQP0R9jZ8huCs/yC7cYpq6sqZYcU6bebJNmtbtEwNA39pkLG
E9vaixQ1gKsPh9GpV1B2pHOk+M+3guoswh8OsqbBrYw0Z8ePTADy2j6nryHWKwdL
NzXQbXGGvPxFmJkAU/MJSvkrrq0hgOKfB0ZNcZZd77wQPmoiV2BAiVuVyR0xEVgr
Sheb+NW5nX5cQS+0Y8TjL5wKWVZp4a1uKCsKMvTX9wFVWiRmhzf7q6zgLbNbWm6l
9mZdkt7lzkfQu4r2D0debNzSzgm1CQcBk/YMhtfPd4LUq8dNxKRVmooRjGdlJ/SC
uHXftJ1/ncRPBwA7Ucqixphtwufu6UA9+/WscYa4lRwzQjY4Xe7Z8iqE4LctEQuw
Q84tumMhEAR4DiaHdPHekAfTfCyLfImwKNiU637BSUukb/OCIIFKyo1xeCZZOO5q
A0SYffB1omOkgAxiIYHmmIUUdZq7ww2yYcJ1KqbQwXlzEt7Q28FmnhmLIdpVidDK
2eG2LOAAWOnD5H1IDX7YU4O2kscQu14wzMjdBRXQJSxYneKtaTZ4/sXcn54qc4Ye
j77Vw7OT27+PKJSalQ2xW1J+gxXZdlTFYCbnJBdDbdbLiF3hqJWpDgiICAe1Dax5
brMFI8PeTfhd3FpQaLvmLUbtf5BXlHRTJgbR/u8W7UHmNzdiZfovYEtOQWW0LvE+
ojRjS/HSXrhUVMpvXKlWvq4zrg8ezlI/YddMzNA1V/YnsK5W1GnXeuMJJkcg4rG/
QOgm4knVFW64jZo8tP/m0HYEdHURPwqJJBiv0FFZnR5FngbUOLruaQ2M2IueL0q7
o/dQPKg30pMI12iwqIMtfnaVoRO/Qhx739CM9AlJf80BZL1zZkBs47CHMeUXIeBZ
mL+k6JYZRmYHL+zrOWZsPxq2Nr8f/JJZT4BjiFwqGDbZieTqD/rUUJQ4IoM8ZDTU
rIMj0KcGuA7R1jn8scDckUtjXoMGXq1bYQlTs2D92cFc3kP0NwwcOr9+Na9C0YES
G4cOouPqBE/Yau8NegdkmWd90cPtw601f9cvJ0ApXqE=
`protect END_PROTECTED
