`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rQE7Y+mI6RWGWR7oXN4KQwurR53gSbay3NATB2GqU1n7q84zppo1QR5VlWb+OFau
4ITH8o2eg6JaM3OPrpfwSygToscwbfXZX9SPWSw3jXGJHTgffn00gvTi17O4IP/F
KE5mLor1pT56RrYRrD1sRuRbvS2yoVvu22vJK56v5R/JFRr7d+wiygl9mw+uExw3
WklTlGGfSSJXhfU6NUxlcu1SSAPNEA8Hpgxo+3KD+UauKDKW7u8RXVFkuplND/QP
nZ2YK1yWfQGjvZDlPtcFCS/l+rgszhVMBowcdTNSEfnjsfk8B/gRin5sPxhh9FLA
UHaki7vtRRlRkiSrLC7jaVCfZJSs+qsPkUZEMypiej35QyJBheURBt85Cn6niaZH
xh2d/zUMzOcTma+t5nuX4skVzrL41QEbSvV8ZDQMZ+wC8VR086RFO6pnrJnogjDQ
ce+Ov9upTvE4A8j4VJ1e2yvoXz4Gcd7BijCf+r2CBV/H/OuLI2NBUNb7Yfos3izN
W5FSY6tqqs1jB4qHTWWQ9HNBwuLc7n2a5ZVVEinHZxI3FVsmlUQGD/nBT7XluUM4
`protect END_PROTECTED
