`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Rn+ykwF0tc88y+2rYOG/uYy4yWhaf4RyKcIWdT/72yqJnoNUBDHfLnu0hnpihDF
U0oXQ7nGfZO88gUsZ3UsAJBxIrvxYSrOHrn4VxPRqOOU5LBkBr3Zqo40sXi9alXi
WLLp0n7H94rfnb0UqsB2+h22exJJAaXTrACvUMzgM1z7gJHzs7XQj8VELaoCEZAI
an3fQN+TOspRgl/WLnF88xpbiwTfgJZwlIWsCVtGZDLQ+Ik53byEKGBQ5ChC32wf
euw5v2tJ/FKW7YLUdPWfZmUoAAq40rr7+PTgX+SxlLjsER7n2c9XpTR29XZu1IEQ
+bwryIHuAME0gQLBjGILUl44Z/3+1iJQIKdYdYvgpwW3y9y0ZPbvctZSXGHZWCrB
SKrbHnF1FTPKaFCdWhWTZtGRGffRf4GCjrnYb803MZSHCte6z5h+1K3coasmJEdo
oWB0C6rc5hj56XT+uMWQB+V0/BxDn142VBpzRPNEYnnhCK3cDCmXmxXTW/cWgHzK
`protect END_PROTECTED
