`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
diHbiiHFCIZ8CtaSbdpYm9B1J3V+P8imZtMF7ah6sDo+sLQoph/dJkDKJngUDyjU
c85vpXqGmAG87YAgHOX1wc8FgEKAk4n3p/UBfX5TRqOXHLKzK6WLFzJGmV8haRM3
D3YuQ+1RdPEiklIWMQTo/SYvl6Hk9UrVdHrbe5H4KPiPcqGpaIxwJ9oaU7e3hjcl
Qaqf8+SPjpycpCUU7IbnhuZur0finOJdzRntEnZ8DdynBYPkSfngvk8yWy0YeEFz
rv79p0IYNDgBaRPYw3Is3LCFlOuqM1vEMqr+7DjqyQUjJip25ezCeJmEw7aWjtKG
9ULCpvSfkvyWC4lP87NxfhCmwsZCVlqv5Q5rZNspxYGs53zVkwavuO6SDVBb9tz1
kZDjF1/Wf74WI0+LlqMqK37fmI/qn8LaMKcrEqlwT1H5S48Hnguj+s9bjN58g2J5
CqlqedIMwE91pCaRNzEgK2aUXBwvHD5PJodSRSMoQv2hYeaKnNyi67yGiufYPZLj
uDJ+Itv9bSIeQWRM96J8WQcTcWrUgwcNoxeoP5mwp60=
`protect END_PROTECTED
