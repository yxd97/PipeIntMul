`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2UqQcjLH1tVvXUT+VIqkUHwKJe7BFtUayGaE3a1voiWVXmraQcjhZcLMMPU08iE
oN0m16QzlGOkKZHglakJRN7leey69QmpomesuCMd29uVyVpU87/5nJp4ym0pmvka
QNjS1A2s46ennfQ60v/4A1Y9iySGltlyVz+ouXVGfPY0uo+UTwxDAeiocODI2JO+
yHpNvGm724Rr95gmczIF3kCroc8pRmjZ0gM97vjIvmCPqK5FXWjVSLVSka3CKVpL
gGgQ/H0WGoXHB4D5Ff/Pww==
`protect END_PROTECTED
