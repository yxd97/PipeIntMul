`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mtLuyMDGcSn7oghgApWOKbPYHgVHAoy6fx7W+gEt0Wh50TJJeWjNHE0mvBcpQEGm
6105nkJ5vVDkRhhdnJ78F4Y9dN0Mi2HVKrYL11UQEOrvErfxTJMj7YIs+WCBoltM
CSUdsLDy0nTjxoR+AltTY6WdlFop0CEZ9jSec18U74zrx78SO7iNXOhZ64B/6Xb5
70jpdlNb7CCQ1+pnM3osXB1FTaIupN0m38hJsUHukDmoUh5x5rcUuwy1rYwueRUO
0k56jiGaqacdF4zOTvtaY8wE0dA7ZZnMbbPde0CeI3XoHfwom8jb4N4KXeh2A9Vi
3/+bo9TF8UtwYydGp1+nvKh0SY8tSiGrL50AAZq8MrGA/HVaNnHler+PWJ7sX9ko
rsJwdjXbM9Lmux4I+nKsiRVadeA5HqA7s8AtjwcP5CX/F+TcfEw2TIC+qBdaPm8v
35/l1d0PJ8OV0D+HkjeiqZo14f34Q7F7bmtrjxOtzgKpc6Dg0tqg8o8nwDVwGo6g
q6gA3O5hhxaoLFUWYimo2hFKhSc8w0/JZ307dJN+AVuVTxKpNGI1L8bXD9kjdQpC
JF1t7CbFcH2roqY8BIdTYlnHTNZmsNHjC0UmrMS5olgcXlXHeJ2qRKb++EhrhNyU
lJVtVwiWdl/r7Tl+v9bJ6/ZbecS0Ofvl0tBh4JnX+apmYY0EbgGlFhe3CNWnck+5
B8m2NRghaFcfWTPOB/O2H7rW9n3lxe4a68x9qQH9VEtGrMYyyoq9NMpWgdPo7GfR
RfwAA1uLFId4IsTZsxrjGocTqeHmMNDiFmbioNoE9goW+keSRibzCanJ6V/NSQda
uj1QNSfp20J+FzVytYmwavqQq/Ht5K9AtXJSl9oO11T7Sknrvmk9qvxCbIrA/jjM
jO/sc28VsnkwEf6qfMvhSs+xhdfRSEzEPPbgNI/q1NWsLiDIK2rPNm3a0F1NbIAF
ao+SPtTmmv/E9/VeGwoz8g==
`protect END_PROTECTED
