`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xgbS2qiqpnHGW2s7yRBWgaeSh2HF3w4BpnNyyO2lrP7LfIkgDYF7GpMrfDOPRRFU
w87sul6bju+NgzIDlfj2Jpkm5UFpl3egcrquSuuF22ubtkzRmaVlND1U/qTsg7i9
ENawb4qxT3y1R9RFczeOnPHY9RFEyCYNdqwtTZECdaEqVClENcRHgNf/GQlZKUnH
9djKdNgwDZmm/+B4x65DaZTxRN7rZOR+bj7AR7atIDBD+TCtpI0tjzKdYQc2lj1K
VN/iXMbHMhVmHV1UfviPMtE11usxjGF0TI1uT3xuvfPAGLn9XkyWHEPr787t4aZB
wTtd0AgUG2TB22JgQkPIO+I6tOcVky+Nt6f7UUpAMx8AZat9wVruWWB+iBkUrRz+
6EutGAxbQtcWdVolZyBFggkoguKvSVcYED+9aGgakzavE1cL3F7RUmXqeyR7djXT
`protect END_PROTECTED
