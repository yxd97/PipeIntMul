`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ciFNslpJ9UiPqxQvwmg8ZvfhSYCgL+EdXJ22wgztk+LpkS6MFhhD4FNrIFjR4MnH
/ec0jeNR4H90HxB+vg7012p27XNhp65j3XeERl/WJL4CEg/ftl9yX7CYGu+PIJjL
rxx+9X7OdNUwoROozsYtRfzYdaN00KzxjnO0ty8rTXI3w0OgbwsrTSePRSjMJ9+c
uzeQ3WnJbejlmoDuQ53LDC10sh0xg428LdntmdU2OaK6kHPXKqoBxvoOvj6B7uHh
qogSpLHWxkg237HEi1z0+clqke2CiHweWm7Wqv6y8pAM3WfmCB0X1eSmu+Pqhj2Y
RthNTEbtVD1+7SZFq5aP1o120PlP00e0CaYLgOkfp1ZqUhJt2BVHtgsQvOH7TAAw
m1uNpgq4vBCRfjmMcCStd3gvx6ZkCh83DRaCDV/ZPTA=
`protect END_PROTECTED
