`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qo0lfixyCTVb/Xj9rn016eA/UZVf24hWS3Zx0yrhspZ+q0Sd4T3eZCHJIX/3vedL
M2MoO28ocyW68c8hO1ZYWXpcWJnpYIKmFjTFRT24QbK1pcDWDIjAwRGqa75bt6Xd
GqojrWQpNHtKo+H0FV3HE1hxZED2Ml293VC1BslRBAn4snolxC6PxNduUN4Shzm4
Obwn6OACu0QQfxPHbWOBNIHuIMMOhyTZWfAJJUIq8B52VmInvH2jiaUQVjnKN92n
hwtnpQ563Gp1hn3XWsjA/hqsfVVhwI+tUqhq0uyq/VG20uSUEtkkeXzppDeod9D3
OwpPWMVMCZ6a33n5NSWCbsJVThda3z0ZFjh/Hu1bp7EDV3bjI5IMJy4CzBeV7dNu
HjXJWwaWkhhvHKkLKD/5d1L5QKHTKoaaFO0AvKB47AfEeqnhKEi6OT5uXTGtUoue
944erG27npHUmwge4bcUA9rUhpfu9mALH1Jcnu50Y+IYcV79pPKM4x8wQh7j+XrN
eZgzqInBO15pfCNbVqAlglha8cz1zxF02ULc3qCsU7aRY6ucYENl6wwWYcAQPx2H
gfozQAMrygguD5MzXP/ZgII9y4lk96JjU+K/gNeZdKi1WOquEUYPbrVvQwLPGdCe
7yeOM9LVuSqaH3bn6UFeI1Lh5yJZinWfdcijxe5BZAtqajm1GP+81HE3RT4RqvLt
QEV4AmVCyoIbKL2wHAXDZ4AJuiQC0A4dnnXKalmVRLu2RrAfiZEtrgVeOlHcZGB+
5RxPMm1+1E+ihPyNThSvAmsAxe9dO9Fh8kXMcb7NR5xlRZaZPCXYELmQOgxWyd+5
WDGj1aNtdqYrfM8QwKIuRUdLdHAIG6vSGcX3cKqDVtN9JApK/gosPIZRlxwAJCWu
s6sqnoqomY79+6NChRVGChB9o2eJym+539xMA/Mk0UEGQmlMw3BrRfobjiC3/BW2
bugFz8nYX9M2NmwIWwNQ7DHzsO9KdEleklEdl0UV++TyDhvAsOGUZP+jkB2IAs+u
EHAbHifZhtWYdqscgfRyOigg8wuCE4refirJaikbc4VCjT3oJEmD04jPLmfHdBJL
IcM4CZMLorLTCS36kZgTvsXZ1BjHMbSwnXQ1KQKhGJEPt8pl0P0YHbbAm1N0CE7L
Ewr3PYqnBmTD4Cc6JagTCbU5C6yRzNUefGfdV0N/JQtobAGJuZiIARXm3vM4+ge/
qrWkkVFr0XXEgGeo8NItDURYXWsgJq4fvuYtKC0BD0QzsoRDh6RFBT1X61aRYtdF
OF7aD5xyQm3QnrC1qTHxL/KzfEvNGHOtO6XZ1C+9n/UQF7YgkQbQaE/Akhv5st5c
CopSNNX2QdzSteHWZ4ceHQEyc7IsTTXkZ05FiXW9DGoJUsW4CIw9MXWvyMPH5kEK
kyAMRzHAdPRi8QLMP6MRkOt1Z00r646dfi6m348h175Pzs9g85JfTcjbwtfROl13
DcIf9UFtLITQFuQao53zHY+VjnH/OJBr+R/+k2lo/hvn4Rfi1UTjVewGPSMiN+9y
hCTUCitvYdlEMw4cm3Se/YlhpOb/YBKskoy70HXi3KIusmsAahWx5F8psAcPERdM
2B/R+fvoBrakuQ5CM9DCTv4WVBABuKWcOdzQdak0wE0WRfHnWRJFa+RrwCSj0po9
1ZbO/yr3y5sJfplVjqtqjyb03qOxdV9DJI94rdaXZ4GnttDtebLgJziPXIh4qZ96
`protect END_PROTECTED
