`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+mSHNdJRo3+2BnoiEOkiHQkyAMo/LC1tb86jvg84HwdCyx0Oa2k7vN60fCn42O+
KbO/kd3/odr1fBF26qfjk/l84x09oNanhdbmv5b/g00V3vDrZpve4CI4eZBRieUP
RV89TV0FZYgx4yGvHllDo2EJ11499/3KhOxhJD7+wSGgn+OJz77a3k/tT42qo0ho
PgDAYCdIL/sTq0NHt5TkLFXumkpZpxhh3OgA42keUjKQJYV6b+3EZJxGHejOfBkb
jlls2YmFHlkkLrA3cRyaBJ/c5QJYBm1JD8Vme17YfJ4SkzKHPqLER4NBlya9hHiI
zp1Daq/WLIXmoxlb2ukwF4uSVjgXEMeCL5wyiehIjo6sdZNXpUcBZkEVEJVR6sph
LcHWh8XEpDvzucWLDL1blAfH3ekVgBJqdJMdrKZb1w0=
`protect END_PROTECTED
