`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O5ekboOq2/v+VZefDnvtxIlRcfmtzFWtLCF+pLgb68850nYdqHZ25xpQBJMn56v1
t6uhSON+gYlPSLbogjfTewi5nfc11bDprPqKBvBJpVE7atLP+heZHaIWomctVpDZ
Cxxr0+9L/QIq2MFNWn/IqPt+Xh1zbGJ+2vib7J2Whb+jsMpMZdbTp8tf1uSRDn4F
qB5+XOgqYqVijPstR5drSi+8nJwb/uvfgdwj1hEjAiFfC9oOYftvaQKDN5/kE+uj
tq/DP9hJ5AKIzmXaDtY+6TH0tspr23a1TnmR5aIELWrKItl/Fso84rWGE4vhNE+M
B8yT48fSLNKqwOZXrsGUt+8+2hVAXkJthBEe5xe4A/+xjMLlEF0n+Cv5ZmY9EyA1
G+YbSPjPtMhW5tFqQvSIR33w57nshNiRBcNLsCaBgSE=
`protect END_PROTECTED
