`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a5lqX/2pyvBXLp+rfURHmrq544kWhkTGC3xYQGoQy2qfMdy+0ie9zLC/mfMYDvjG
rOgG6q7Tz2JpW/5V9JCquLq5H0AUK/JgDqXyHirZCX+DY2xJBsy1YaJC/2agrwbj
r7NDpRXFwvHy6ZhTUCM4hZroj95bN0wClnjcT0zRhLfki0UgMEvhcluT6muNNY98
/LOHmhMYxjcDPV9dZ6/AiZ68ZlY9kTlIE+G9dmTJz/IRCmotxsN2w+zPXwzjd167
Z0lILKznWkSryRJw74GDtpczFAHDZ1nheFKM6CNexkM+bTjhGisXayxK6FMARWK1
`protect END_PROTECTED
