`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CzOLWBofUt3PGFx0xyClw+zx0rKTcQM9ilv7Yo4zUsJkC0V+ie8hA2GlgAi7EJhp
Yf153gJX95k7N5HNm/0GAfVjMydKdD4K7HiE0PA0mAeDk1cK9FwjY67W9MjE3q1c
ZdWqL75xtxlwqwhFnTjbfvrBTzdywqEhC1rPGgpbfId06g5YhPfRypilfVcFAIM/
z89p6kO2oaHTKBAxRvl2ZD4OcSbGCrg3+zwJj+QuWgeUTO61J/6Y6SET/+TE2P0O
TLFG22fVSiXE30DrAHVdIMvifaBu0xHvZsEUJJEqbUulk/JBnguzTE9DryUj1Lxi
P65vrVmag2wanqh+cSmhhaTPu3iiFo+DcbicKD0tRcydipzFvAQ/MYToB2UOx9Aa
TF1OK5pq4S/QORqJhsefA29QLZ/WN52iX3DegqCoNAoOZjxrOApchgWRtFRtQSe6
idK6Qp28BcN1HWyhh7mZoQ9UqCLMxcwtFRbl3bR5c4XF7hteUpwgo7Cf0wp8sfVC
/oiIXLbkNzSEMF80Jj+LY+f3lBPp4rlhX/WiXrCMqQVwSmUr2ELWt5yLr8sbgGBl
42mh5lBnROF2p3yindVULA52o8oZeetzXdoMFx3hJiYiTXcA58+Vqkmu5XWTnytZ
YujwuyTWlVg0ZSiHQxXp9T/++GGqzDRank2VodQieDKQeKmTIt3uZg6xBnKUOJUM
9UIdRBc63VuES5fHNJogMPyn/4JaXCgUjpqZNWpkSbLlzuJQJqv2vVaGmPJz4EqW
ytHgu3HkdIWIxSgUDqo1YLI+Cti1XBDw21TjeBLRlHVaGt+30WhSHSpOiF0tOKqJ
0NY3iB91hvWxEWFgyPQC8FsBrA79dNbDUTrrq8iSjXZFcm/j9AYF6xZHpwBV2sNy
sLxb2dmPJRBnnRYlwiAqMd+UbG5ED2wSOiFKF7t/NerjBbpxbgdHTXB/Jk6aY1QT
4aa62rb9wtQkliFKbArB2AFkkFPA0kJX9XHIkdLNatxReSqM0pTWbATkF9k2SrSZ
QRBIh8RNbtYYHrTlYW6S/rBDLFNYAN9omOVm6MMC9G/ytwn5WZ9AGJ6B/SBWFenM
sIwYMzWwtb6AVUQ9S6RrPpgqMoBcMCdjZRoobMHxdJJ4a1pv4J8kVJ8n2dGBLrWS
rzAhyg+BpxMs1gP/DFOmlrdzSTG62ExsSl/rwMzxBlIt1o8iTitKRw3qzwBfBUkb
Be2YPGCQyl2LeIyCXkdaHmC7kqEEet9neIdqYsRNNpCg6EfO+KMsKMVXG+TtgsP1
6UMu0k9HNrcpEHlVbaAFQepNShsuH2CvuhXBbHsk0lbjNUP4TqB04E82QQT1+Rns
rBj0mK6u/XZi2Tu/TcLmxLyISgOKduvdUODUuDT6hfcqoszKrOPHLgPXxq00cvcF
jz5e9L6chAs2irJZ+2HsU3FBNWCQdTQiYKZ8ByYQSoAldzTCthqGci5xJb14iLW2
h6nh8g1GykvZ+cS9DDvuXaE9HRuadWJdylWmlCd90qT4N4thRLzICpLiw8UlzI1Z
NSF7OnR9xBq0POnpyjZwEMCR+jg4/OZaceUbI3TTAQY39TiUNAQpKIDBLE8wRDKH
aP8W8OQtUUcB5p01FMc2ONIYc9bydzHnMfiKlhsofWAo0EisMiAaDimWRio7/BJJ
PcfA9SzSKf/rF0j8YRI+ozwdQ7sy+/kAeTpXQHiLd3elzLcojZllHbFeNZv+3EE4
XsL3YP2UjNngIYuRpNfrbDCBktVucLUQOeMDGQ5gdNcyqfUt5fYMc1rWDnMAO+dT
`protect END_PROTECTED
