`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frqvQumQf/e6T+GhOfObL9HCGnSH+0uyR6VU4KRX5q+Fqw16ysCiFcM6+s25XUoY
2Fs+PQ7mNJROQKKlx+RZB07M7GeEIo6WQWMp6O21aoUZSCES5bm2NKbrJP6TO80j
BwXcwkkMumk+4VWNu4l3dSoQ3v+3/UIeRbsjrsPKUOD4ZMZXeVHQEigrchIdlu5I
hZ5OibEs4IT57g6+XyoxAkqYkV5in36lqn4s2VclXJz3ywu7pnDlufzFCf+xDGbZ
XerSqi+R+L54vOgul7rS20/gxd7hHnVxWRpBoqHnPWomAxFZ5cSwAde3ym1KpUC+
vR5fiFHfLnjtc9ldbpXfyqrEA1iedPfYW0nUEI5XzwzsBybKmusivBNtJSQF4v6p
+/WLAPX87dAol2dWHWYqrCUWFZDcXfB1ObTZNi0uOyy6g9NnreCFFcsMlN/1pHwp
DtcT511y88IJN9GayKVlWQ==
`protect END_PROTECTED
