`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9UBh3zRX99MGd9rAgR4T8wytCxp3OxVZYjH9JduOhvFy9dGRb/x28GKNa1M4qpy
AqV/q3rumhhOMjB8L96yXdraIPFdPdM80IWki25/yjR4R8ExEC9qQbvYFUDPDLCd
uRQ2cBx5s0J8M8m14wJs0Gmx2XU33Uzu0/MuBg8WVikvrnCMO7aVZDsMbPC6Ug59
WL02CdpR/Yn+CMJEVdOfa3ybUaJinZmvZAx9UTmjXWzup0CP4rcVsSv66ne5GuHm
zxtvMP2UoOSPL2junSOn1Efjii/EOq3xdGq6RPaAY0c6GtBz9YF0/rUST7EzvCZB
c+V4K0nTyPDbMpnSmwwJsuG2nMhQp+haZhtWJCkXOpQZSQG++ClSOptXYcmvbQsu
CN0gn0pedJV9ZplrBVOThQDZuLo/xxK5TyPe7IF6rP8Ec0Jh4xAKJD1rwBOiRpOE
X07CKg7IV9zxOGpeUi7n+P5ixZ/1+Fvr4mapFAqqbm4dvkRlkTHu1+63Rc7nKzqm
jMGwOZ3yutKeHJWtnS4ILvgxl/purV1i7D9C0d2bg74WofldkZ76X2m4QEDfMqH1
Velj+oMnrdgHxJHwUwEVqPLfCto5tmze2ee9RQMpCxWkD9UfPXlXpe7bbZyu6esC
Bs/x8MTbGBaQ8iX4YhMh6x4iBB3WeSOS/GQG3jFbhGeq6bL7RSAEpsRzIhmDKDjv
A+kDgReGQq48S+r/KwwMGns/7fezP15zYk0BOohg4ytvQgRy4tbJUWSgaBlML30P
pCUvJ0jSRN7B8TY/d8viRw==
`protect END_PROTECTED
