`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lA0hiCOtGgYKSE7cCq1zihlCMILkDMthF2FhRlUM2sABhtUiCPO6udjgfYByZ0zZ
nQS0vSCZUI+mVLkMReAebnB4QoiWKcXLCc+wvYUZ/SWCp+QgQAcw2fkVe/xwHZZB
wEIM+Y4JirJRJgloZWFjlflwr80K1BPoDq2c8Ia/FLiuCo/nY5d29tG9Qht4Y70O
hKMHCNHTuMtyfKjDIBYV0+yuhtLDIzVEbVNI84k0Yj4WlgpIhdoh37GdLOLxBSE1
vUBlypaK+9NnoDNlCo/Che3wCPlKw0qZNq6pnTGmWgTLtCW8zeN5yEWhfhFly6w9
HyfyUT3oVQ12EpNSdyST+CnfZM5aef6IN4wO5TtpySCwfo5X7svUAHY1q5MCcIZV
+qoFEKu4LHgY4JRPX5LXnq/w/UvaYMNmgbLfShrmL28=
`protect END_PROTECTED
