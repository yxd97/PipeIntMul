`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7XBEn2gUD5Fm7m2UvlNcDGdSFwxbxlax36hYd3lQPda2iSSrONqDJfb8mKOAM9as
VDZjOmelwxdU9sluoiW362tc5Dbt2aYMl7kGWe4pJJdm4SPWbfBPdTwM8MeEEh0o
wFuZUVSccTsEts+we0X0F00DhziGBhp+21KOrQrqHvpvEk4ZNaZQ1Nu/GF5A1M3X
6/jvXnClq9/R7NG2iqYTx7a/GQK5BxM9GNs+TFkrw29oJPu6imFu0ciSF+/WA+8f
GuGUOTfPU7KCohmDV+k64Rr6zBwg6TPXCEKJCx3exk55ydS4p7u0rrLEjYs9Ou8k
FjEw/8wf3ow4lCZMF7adghN1Y6uEp1o2nDqjkSt07pBKxTverKjeNRgsOVaYL0LB
UAPbYlIOzOs9r8qwWFVBcLIOUBZ0l6fea08uRxglUlvmlyE/lx5sv/A/L8pxoLbP
x92tN2AofT68YWhcQOB6kxaMm8Dl7GuBJ7KQ5JwdymI0NRcWkPNslV3ZZt4jO4M7
l9zKW1F6vudDxm1XbnjH27Ynk5W4RKrcms6OK0LSSKgf+eptUM8mbb0UHezJiXIx
wZSz/TxdksIAUPzg3PHl7RL7tv/7+cdch/BWjGOSMztWMOZgr51QfSZAfsabTxFT
pcXWIr5UcyqH95mO74wGle9xzVpuoMgVX6NWHwRS5LX+gfJQCCX6j6tJD5hTkcRU
TBIsB6nRplSGAiQEADD4e6nk/PsV3pGqmOR6+E0/0aoF4yndt5KqDThbclmy/vCI
lGff+ErqgUMLuyK5HpJ48A==
`protect END_PROTECTED
