`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o7b99jhAJQ0MMGx/YEL1P+sG6d+eJoGdeqIH188dwmJ96AzJqI3zWri8xGuKv9yM
kJUFk4um9+1ET9nFAqFOhJ50/rJ9Qju0zPLOMkmpmM5bji+UIrixd2Oo7Owuwec3
6b3UGO96+8I6vkRBWz+RmErlec8PFkVywDtTZSUVgAYkUgoPVZEUwCad990lPhcT
MtHwSWc+20yMVGe4VWLdNg14JbhjjBDgvvvi3a0tvYN7leWhKfEiq66Fs6Yng+NQ
3F4MDwWuQkm+JlvsYKMmuR6hlKitnuihqPsHAjlYImu3yGQLB3E0sDz04fMo+sOs
aE8J4NceT74KduTfq1YLFf3fcYrWKxUPX8KyWIhjw0WeczkyCBiAtzdNrD3CAKXR
CXdgZmoEoeZjKswa70BSQd3D9H8gOQReUwtBsiBcGcKoWiG60mA6JiGm0FU6kjMk
ElNTKZe6cJX2jO5fScTdvTYf/oJldsUnknEKLcZOTOkCdC6zQmEP5WIXHj+CN8T6
pJkmZ6Hb5RiOgSKLPQcKwqZV0TIc4Ii0tyWmTBo0GJ94yfvzAYZkWJ/TRfQSMlP/
3aj4NqcVk5vvFoUGi+40cFBLhPDip8TD0+JSv0JFL06EQ6kdMcaC7nfJZVi5hIDN
kSi3q3owlDOKi/pL4F6FdsoeEom6hnQxCiqWlF6csLJjQ1+aGGoNFzgRYUpkBLvA
nP7ZxxXHrvNBPteV1+d6SAwRqjhAoy0Plr2dfHnjFjvbOneBfhTw9+0B3A62o2AJ
oADZgb7OFSb51PFCcArVZA==
`protect END_PROTECTED
