`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ag2LR/xXY/jbchZ4JJi17xCSnsw0wKlgHCNQQobUCDbMuO2hvMF1S/8JFgwoEKvj
gpBUJwqXm/TQrp4vbjHDIqfuBmD5mJzKhhCFLaQy/G3bgQXgK0+fzEISeO8Qko+V
MVg5/Sgxi6scXOZZBreFBbEKqm3Aj3qM19zVLvSvWVzqh7h68qsLkdlwjcimN2dx
j5aMTUfcJBuDMjvW5sAE0Ag2wzDCMFsXFVv4QdJemP/aqjZqeKanDZidUlhUn1WV
qK9EN48KvCjYj1jDlg7qS6O16ci0rUA4tXIDukk/AaYPLuMJmfORWfOvW05CXcbV
II1zpvvNOcKPEhDKEdMECg==
`protect END_PROTECTED
