`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2xBdGJHRjOMeoVewcCO7TiZtoMK+CKBJlOLZ1byTcfLKmjOWxxxsvTQSQFechgqP
gkfHSpFUgCEH+DXiHv7W5eyfvA5xFiitn5hA/WZKKy8B3JaIz86OfbL47LNYR3ar
6gVvR+LZmYEFoCimoqq5YvwoswkKcJdL65kNCgGaVDKkMzwDY24+WH86lVM38Qut
Y2Ozg+j515gUS5ZQqDDoJ2EkM54sRhjXxi/hUWI3xLnrpmvwjW1KeJlVSY4UtrJ1
`protect END_PROTECTED
