`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cc0FjsnokFabBEzlMt6UNhWtOEGrHv09TFV5V+c/Nf0JMz43CgBMrLpOMvXsfB6a
+Qtgzrzd0lGUIAAwpgU9aAuKMDAYwKs21jdxwfYPHkYfMS7ySSJ7wux0ChfkOEgU
4ZJI8oYkiGSGEOd02D7GfjImRaNmQEdxgCR/v5MXiA5JlOktxYm+jqWVuwxLHAYn
xGFmPSjf2ret1EAqBKi92fY9Zykfx02kh1dTmNR8fEaCcxWPIT1A5ePTfI6UJMKG
g2kyFf9JYo/B61/Ugp0sEg==
`protect END_PROTECTED
