`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QX9UqCpQ1dKIFGZSqo8LQex9tcDX9TMNmJmYsSOXsus33Fm97S2OKdw6hxqGNjDJ
+2ei3JxvuUrY/kuQ2GCYMQLSgAjWoAqh6zacR8lFLhMfGhPFFt5zKgiqCU7y10sb
2QNf+pNSBhO0LVA5mR2H75IvD2ZmAPxSCF3TNCeKO/1dX29/KWI+BAhn+c0vEoAh
0YjqKLrCWy6ivesRBII7FFqrlcpe/46kAx3U+fVpNueMFzlf3fq91j41nW3QDtw4
HJTvfjzMuMcm7xO1UhD0H1MyA1goGh/FAqskRnuLKOA=
`protect END_PROTECTED
