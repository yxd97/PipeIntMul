`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihQupy0GG9uLRgfO/HNf1K7kMhDA+TsaZO9iZy6i7VjW6t16kwBnaZzyYHn7BPC5
n4v1Ugnj8JOTmAX3RrhCxVOO73h6dbWaOmCKjDFNs0kvfMXesnEf3zJhADE+AEY0
aGk9chc35pMyF+wPBdu8t6Ml6AEqVy1H4Tw3xy52g0PfXAKBfhbuCOUA7jlC224S
UwlvwMwkC2Zw6A2VXnDiH0/o3EkL1aiR2lJZBvhQL4WXowk4FjBGmTpgRqaiu/oN
PTDYHDUnStkW15RhiVzew2wZaFZ1iLFHQD2qq3AbhCbSQbL50h7i//ppT6/ShYMG
aJKS/MpfgLXleWWGu1vDVn9sK3p+0fu4FzRggWsk6KEdcs1Bi+pZUtTG7BdRS8KC
NEt+t9WZZMnjZGSQVFSyb3APRifNzwg48GSijDdGYNuMVxoN1xp7kJJ5LpT0Mo2Z
`protect END_PROTECTED
