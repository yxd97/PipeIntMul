`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eXPm0llU3RzTOFhLYBZyHeAnEJpLs1P6IACteElQBdrCJXCOq1zczqyYyDhzUYVc
3cq0MRB0CR8CxhDPEqZtBlxydbQBEbO3sBB2w5BKWcvQlj8M8L8jvWzt69yaq2R7
IY9wxmpUUyGAufMIL5zQNQh4xf2Tyu96Gk8DyftpbR0OfcWWmiPo/iNtQ4lUZabY
j3A7Unb/Lr8XozaMwWRHTAqPVmmkvTrohJAD5/vtxokQkjMjHwj5O6IISonDnqNG
a4IBp5GOvUxTcP8fxfK4HQw+4vJrn3hWvqTrNciZm0libQ3C1hqNwBzwg+YC8KtP
MC9AuGZOLRKQ0xJWh89lFgn5YlYVnq6Rg9hTaasl3mYPbHcGbJEg2LtoO1QWxv7K
`protect END_PROTECTED
