`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DkMPn17AJk8+JPDiXN6q4WcH0XMysguq4kQXAFshCmvToQtHtOvXcPuNVhJCaFm
FyoNYI0IuDWI7ZqKMIb/xtTBahD42pnenvBP09jB0mS2xikoryzjMVuSUkIkCx7X
sE/WBdS93NGKjmS16W5jz0HVQfRqDR3vYhdMpJx/Iua2Y9SaVZpjtrnBLT6262Bo
lpbr0KEL4/l1yU5Z/5u/YGjfxJLJ1RnOhZQy3zwBshvSKqA03NJVNlvCMOCTf6ZH
q4lh/c8XmE4T6PkWL/dVSFoaW9CCwFaxNmmZvnubrdAm1oUlXGTYiVaU2Cs+QoI9
XYhtULcs3fWMsdPOlmEmEF2CAXAxaTq063uDU3yD2hYwR4El/onQ/84jSSOkNZHK
EbdzHOjeywPpCPr3aoui/IRBqGmAkLtDOcX1s/R3jfLT2SF4Y17Xx1gxKdhDXTR4
7wxDIjo2HUFB7wDnENqWnT0OVoqs7mn8UNaQmJkeLIxIEFuBuqI8R8jSBJSxTmum
8+Ae/OC32KiqmTfz1SNXE14TFFg2rY733z8Li3Gq20vIL040dPStj+pYy2dfYMkJ
Gxgv/YsmMnBB2NpqfWyShtCXmqcL2DUX0Dvbsw8JkqY=
`protect END_PROTECTED
