`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JoPtgZpeuFEuvrEsJKBwum0LfLztcAPK9RGR6pc9Csh7Bv9T3CSKUJaCyftI7Nm/
t8Sn4AANAYsuabaibQv27rX2fe1/h6rhWifKtc6QLwnkuFrhUwh80lVUI4ZOCxtV
0N+aUP0hWn3OwaFLbSAiDmF9adG8p8kkD5Jm+emLjJ/Nm09vGgM+g8SP1vgE+GDo
38lu3o1G6WdS/N3AT6IwycwjFqfdB75CkIzuUVREM1wct3W4GIY5Vl1nY7Gf7j7N
RD5eg0wLsCtuAusGQP5xxlJW2ifbivbWRu6pRwBjQk7jRhpAHLJlZOq6rDk6c72x
kpm4Xd5rr35QSPNmGtuQTQhzI/smvsDBf3s5v26xnZmJ7WHVI5BrLlsYG4H7IILN
6etV9+pbxQYRcygZGA6sdcp7iGZEU8gVvS/QkZiGafE0w9G55lNIbdudDBSF+40i
GVmA4hnTAM/iF0d3tPVf9rcwBgDnT51WAWg2LrCPbFnscgaRrDJ/gcJRXaTlaGT+
k61zVAa47ALp3/Fga5lP0/8P3pDDmM2WeoM35G76OBvpwc4REiW2NePECwtW2VOr
oL1aSHK3ey3YHW8eTuN+5//kTDudIQSOz8k2Yj0fS3lZDClEk066QhuzT5o66CXq
h5b55SARN4zzN7bWDitpmW1N7PMpER6Alh4BsParrZM4R6cBzZcDLBapm8TSm0xe
cObz4h/xOLNULIZ3uESbM/wsOd/eHyLhQN3RmVzDHYStaE5UKDUJPxAlHD2IGyQb
nKekNAfO2cTwmbkjLoluW3j4oUoecI6mlp2JgowVzrw45rzOwzvcvpsvZEtnwuvk
LJr4/f1stOO26Sjj4dxGBQ==
`protect END_PROTECTED
