`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NwWfbg44AoO2au0sHCKxNkCYYe4WrR12RuFFsA/ORZllQ9WUz+qgu4r2akzurX4q
seQ1/TRcie2USG0S08tSdFxs8fqfKepIisBXj6iE8L/3lhS0Azqv9ojjjodfnanQ
5Zt4XdywnZyh9cLXSAK++W2luQAxquBQBMwcNIEuZDW5bt4rn10/NpbPI2Ahqyxq
ZC73ob+1V7Z6IqRxfY6gKpYk3jAef8AyDI3NJwoCxIouKCpXkjAnzSdYWq0qJrvg
ueBMhs6YMFu+9YMqcYpAHrPP8A5Pp2/kuwrNPUveAAIbSpdx0tvUEWDFsxXL/00Q
qlNlJL6BxgNN3L8nBz/LfFCCMpIxkzV8Gn0h3+vpTMkncQpAfRAu1j/t9HyjR3Oh
lZX3h8FkJyOS4SJh4fDPwulx061eNOi0qVpfCyKtxqbfJFNxHifVAY/bumxNvJZY
0VfqH5gcvS4eRIaDQWjA0xbqINfflyIrCcm+bh5NhPD9CzUdnh8mN393y6WhLo6S
cFLX/+O3CjcS5h22pGQ4X1G1NECew1HfA2ijunL96xKWFX8yDbdKfJ8bEkGxQ1qG
nXnT8jyHxxCLtC7OtetMn3S1YRqW+XG8vDuz83S1uXUOAjI55xBM/xB9m3ac8ssF
gFbE6WIZOV9hEIRQoaBunifeHdZYWJYnhODSHxZ4ZrECTzY7j2iDrPRymN23Uk3k
XIALFtovr+idZWeG3Twh9+v5es7T9e2EsY3wou2a/QFymSspvAcaQsBEtOcfOw6L
afPx+DFbAxTGMOaaDuUHDmU/1kkQKRs3wmFz9E555pwXlnKHx7yjPC06IDESJLKE
CJOYlsTbcgsl8vO2kG7eGYxMwlJ6A1/WZH+ESuLgKEIeDQGfzIl9uYRexKgojr1x
KdJJJW4MUij3VehcCUNEU9prDVIpdHwVzYBcAdXBjKjDFrcjXFFQr9OtAycDBoDj
`protect END_PROTECTED
