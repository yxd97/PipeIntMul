`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lWYqXyD0awGahZbvVxI4L5CP3/AwjCNQK8WCtIoAjuQviq8l3hqxDRls0R6ZLlT3
rBY1cqWgjWwUI3ciTYsBmCDAkgX/MUuJLlhJxLxhbfZ2a4230p6Ba7Cwtu+qX5YC
Qi7QRh0dJCp17dIBLeTLG9yecHh2bYurAqbl1qD4SD8lSAMDNbqmQ5C1RO0ZfjIY
MVlyqXb1beCFJLVk1sA36lx7qLcg4QtYAD+1y1ITGieYK9BU7oXJxrMNDr/P4paJ
n3HsBTFmgit/DFu2M2vXo+h4luS5pRK3M3dkyvBVGY7OKE+TtiBg09DPqMUK77Vg
EENDxz8ziweTU+Gqtr9cQeaOlX7r45sQlEIUlW6OiKDoIR9PkmCjpEsWqyzZAPbP
`protect END_PROTECTED
