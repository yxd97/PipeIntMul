`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEvwLYn0RjF7TVPCi1amENbKsC0JZGGYHL52WVzROqw1c09Wk/f97mh+RlenosfQ
b5hw/T437rv0ohm/MJzdaJElsTOc4g0dv7JuKkxicB7xKQ3fWtC/pdgcdTnq/Wtn
Ychl7fOJzrYdYCQcKwMQJfskyOQ0l7kkP4TnGELBJayFHAvI7ERktVa6+Si7ogod
pJqoZtYgoezrowXJTU8YOXMIFeALdiKSGOeAgZHgm0I6ZgZldbsyID7SoA80NEJ7
Rd3OJvvZsuBmak1Xuy9rLEmri65bWwB4zW7NUYrDmulSZJdJ65zIgPyCQI434JAY
HSyghnpeyWnKkgRHZm4fZKX7Fo6zBFjAFgjkF5bqAS/Tkze7jfbDIKwh+l47qeZM
nrkKPzsA3hCFS9dgdS771dU+wv2M0O/h7HXMBhuoLflT6UCnNgRawfyK1gbbM99I
rcx2TiTVl57hCPSZqibMwxgFL5fRLfjFhUOkT77FiVtNXz1pXv1aD35j1hdd3cDq
sEsxq4kkRNBlvKuq6t0S7TtaHKDPgitwytoAu5fFhMmDe6YLZ4VADzickjIAV9OY
Mi6g4jav7AbpQgt0RfB5D/sTtcOfFOjEHWbj2J9vZJjjj7CtirSN8LKGxsaKLvwt
55oC76FDePIqvej13rVCb3zD3NWGZfJC3jksRkvVdlIcqweNhEWAvAb3EId296DC
jTNxjnw7KJbj+bGEeC69uisKsSz2/9GxCHLSnGtE7jZnchKDT86g3kz/NDaQkrty
4g9FLAFCKrEHl3Zn/fy+QIUW5BHfCN3sE/y+ptOg5lFg9KIucBJ5/nUaU8yjHxtB
IQi1gufE3Vk01m5NgyuSsmuawBWP9i2aOZHIe2lRxygjTxohJVvVfbuQBDmUsZBj
TfdPDIzBUOplTI32tDoN/P8F4Q/+bQBtD4idX4gBuRnP+auQiZsCStreZ4xw120g
AyBh+AERf1h6bVly8W1mq03reyTG+doXR2tx2jg58HFbCHBdYN5Qs7K6+5m9E88G
9fGWAB0hVvEIRMsIe8rjTPQVYz0439YA7ngC7aMyeXC1q81uI0mIimjLz7DLwQMO
j2Gdng3LfC6hncs/P7eReYIY0hCr3a9CQHERwDjWGJWXPJO8L+HlFVYeSXTPk+s9
NnmA62VjNAIv65jd8Jp2M9lzU6njs4/xl16VbPf81WX/OoHhmoN+C/valnkE9vxy
RvvX5G8DQMym0aiGgVJUsVllVZvCJxZubAty4wO3xWOg4O7sJc8L+Z05+nmqu6NX
AGUpLpHST+ZyBzDENLDf9eCTdUSBDW530QML1t/54IZSObfIANQt0bFQCfbMQu6r
nQdBO0EJb2XVoEfljIUwtyAIIxw0GuOwUq+HkRk3dx3p4XOlRDxUv0i6avU/RCIG
1yILu+UimC2yv/0VlpgPHUeAMIOjUlAJQ6f465/77O04D4d+rNjkIvkyFOWopWkW
Mo6/dGRQArn40ylBy5L5jn9OBdCVIzvsTXEUJIZb+SfFhTYeCVFwm2BAUoMkqWxG
KKq12lp6MWi9KxFc0UnTeRd/qPG/oUMGwS5+Nbj4QBQ/gjsxlOrGuKzTwAGG6yBS
LcgiuBAknnMCkEWgKVKzYP/nxcQ/M+2hr9Fc7nMJzY/txfU+k46EzVw4jzSRaP3U
ga0XDrkEVJpr6n+PSdFU5z3vUxEM2IajaQKvpQKvFIrqRzekvFVn72dCrNhioSkA
DGBgWOIZeD45frSx/WtCggkuyAwzW8LwXntgG97bKsC5pJnGcO9Fue2OwCKjgOwt
K98g51bpi/SECze2KJEHO7B4d4xCtPlCzywqdwGUTD73PnZ8RHY1B/ldYHiLHpTr
8XWIFjt1glcB5WrRAT+vCen133e0b9fDvSQdSLSnN0l4BUflDhWU1N/xp/yZiFzw
cvARpNTKx8N5yL0uDREp2BSAcRO53W8VaA5MGagQB3R4T3UNLiA1gE0vphbWjyTl
APDW7QsyZUd7PB9I5mLsPvJjrLBTest1+WpS7/vL6MLB8ZaIBKr9ulmhQQYg4x0J
sFLVkAqDifa+zI9Y+xfeDHpr9Ug8aMQ18F3wahiE8Sno4AbNRqGSgokO+WpI1ZEM
kLhd49u62XP+XNd4OGM9NI6Tiz25nEyU1fBhUw1M6D3nEimeCi9R4wZwBIyC+yrE
As+FZ7LGPGU9r+rkFC8O7op1R1ZA6JqkWHT+SyLeZvbcZVX0ZpDvq4vA9VL3Hmnw
VEI9lAVhEbuLzH3JPyzWMPt8wDVGeHMVo8geuj4t+v0VPFjZiUjWfsbhqMFbHWB+
Iu03TChYblDJ5E7v9LyCVsqfuNMUrLIoa6WR73s4Y9ZMrqbkpEwajCw+eWKKLwe5
NOFndqGxEhW7wLLUG1E5ni5U2LQ574XjT+9MDtBLcErbe55vrCkkJE2lTOZn1e7E
FjzgSkad9WPDa6BZkdmjNIJQjZkGG8vxYC6HrrgyG36YPslrWZjHZ9DB1jJv6QRx
pEyyCbqEcb2lMXajpgTv9QqqOy3rRoWxjDVBcB17WZWAaD5S4OCm6WoQoNHK25M/
LMGqEd+rACBM3EuKsSPRw+zYlapKiDS4YRi6ypJw/LoK9GBzpgy9kAB2hPzCJLyW
av9v9S+5SknlTlUuo4yd7g9YbwLZN5a0MkCdFk2FVtPdszRBPxHiggfiZ+vmav8L
bCRsr0VvH+aR1aazS2ERgYUtYRakFpZ2YQjD5Ds3d1c3zXi8yOEuWEfPbzk9zT+N
5elj0fJV3aerTTwqKHfKoZX+72yPnxW9p6gEw+HAD+B0c/XaE4BDfFQBaPlsEn8r
cjZpHviHptrxLya0k0i5BvJKrJ+6Zr+vWE7zJQpMRyNWSJ9ytjWLUw52vtoARMUy
cMRUpNj0KSf8dSPIDZvFYT9GfkQJ7bpOldc2Ldpaqy2DaVYXMon35Yj8GcCmP4w0
g0zc+0eMG4M/C3pb+4JK3EhVYjPfuOZxgFTztv7IIlr7aDHbmJQNl/bW4Z4951wa
E3l/PG2ugAruZYjEhsGNIxwA7KOOqxlYouLOhkEABz2eA9m8iAsXKO8ptzByHbmu
GoQXZ6V+gtep6Q1Xi8W6OjIjeNa6qDS4yagxXm/vXVhy9WMiZOCdn33ZMhddNtdP
XpEb2Rd2qaO3UXSqRm3fzSnxHZi1JkjOd1tt/bHMmy6+/ZERMnLfx1jlHjfSRwJo
B5+ImVT0qadKCUBT6HCO6w4qiqTQEIPxNSrm3CvJznHRJrnICmCfgwwnO94XDM2L
YbI7pD2WKsywAruMvoFYa64mH3W/yZoMnNbN4I4bTyoMz6g5VLM3mKr80F1qLCm0
yE8x+FDq3021cMpoeEFOa/MaIX8jc/Z8hUz0OXjQP/ja66CSEZ7rcYamSN4yXXTj
c9Hnjqo6l53IynzkqZjw1otLQdN0RCPW9CZQW5dWdLQ0pvGh7r1fIYtimmQH5Ae3
sMRwJ0Fp9Wo/5WKaE+Gf9D43Iu5WEgVbd7WUhz3qpidmiAJ6BtdQfjuQVhK5LfNf
q8KHebtn/LtccdAoxVwVmh6f8mJL3ThOb2sbAkKjiKkrw4Hk/qe9BG6hVCB+/B8M
YAo0lycQQEPA/BaoA/M4xU1r9sOVi7PDMShrHtp72xDZhBpeC7ylX6PZssDupfzY
gfTatpgahS3dT/jd9hwhPIPjb6Vbq1KQXJpbevKRo1lEvlidMdqll3lowgh4ilY2
ICTzh9+jTlI0SE/Djhd8rrxZgyJtG5EeHhZZDOwEL2En+qpu/8gV0oCwWge911hm
rkc2BbTL8w2hNiiIE92Z90sMZyMC0hgU7zOAs0hKkjDRdsI3j25Mgy8rA3263n8r
souGi05pzCvB7JzX5baeilNRfwScIYj3m3QbqOZ25eaJRtjlpcEZo4ahfVZ6WbYa
BT3VPQoU0c8nw8OhiSPkr++a2Mh1HvE9AKLlrX9zeN0UmorO9BVXgkYLeaTKl2yH
2tldboA3HTHXUm46vXdBC/1Pv6WkZreq+ixEtgxV+Qc3gmC+lmyO7RK7yqWT+RdE
fknXfUzZNKocVRvE/rdsLdCFGOepR93rL9rv8QclhghQb7FYQYXkgCs18S3ytyIz
UngY+26mZBVrJerFo56PLu7uf3baks6uSNR5B+bjfzNO/l21G+UOgspwwMktXnyc
bbKZRkeZJ36d86CM6UKrUvOARtHVJtAF8dZEWFudbWbyFoN3xtv527wltZMwR20c
xOP8DfwmRaVIetQK4fp77Gp3zuU0b+U+sbG1nWvPnJxhpqGgctiK0MWB21hiQWfC
5eWjPf5mmwbVNT8Xp+NrjqzmRXlyyWuqyOQzSndwopyygRux41FryvxF9g3U3nBf
bCPfQ4RdTccH659/N1O7nXFf0iokAwLvvcfgm+sukOchvKJtJsqNTSpiQAV1r0kS
V4/MPdediQwhu7gn9cj9E63jdng5792Ua3senvDdPoUcY78Hs6/KJenMpD0rJ8Ag
utyXjBrARITcsl/Bp/nBPjdjCSlLUXXY8BzGKTUWpjqXrk2kN7EKNa/TBisIuVur
4BIpZhU9iSRcnxwbl1fn1UJ21FBw0J7Zbk5+bcdEKtEjMUa7RGOVbr/34RUWjmgJ
Wm8S9DzsO9zEHX+Pao08afg/okhQT6BehRSiw0TCiLHGtaHnnIUF/6I+17uAFG/9
PttjpqVKEEGjHYLeKs9IaFlmi/Za4afAm7VxEeOwQJQxQAfvce4b2aF4AQ1If2T4
LNsUMjnmkcQrkas7AyQEmy/kK93W0Sa+XkvdwUyuWOyZGIwdZk59h9M/U2SQ/MwG
yqq6qgLCvhjPFunzaz3/edsOA+4y2qf1uMMGa+g55AegcZIZHk+G4xNet94CxB8E
DdlyhxRK3JRdFnFQE/5VoiUWH1U3/ESUl+cFYMBcK0/rPQAsX10IhTNul+EXVH+P
3osO03eiBrz/wRhYcD4hEiYImIzBL+iCCiObxeJLK/5VQXCOafI91GCgEn/vVAGy
0CIOotDiQ5eI0P1ZFFD/oGbHDbl3vqC7/H9NwiH1qxMnXZ98q0AjI6nrig0V5QHl
LIOjPfZYf7SyzemybZOOAEZmJxb9pHu2SLhoqYi4ByHCGglo3Wiui9imufWcpKrV
Rpu3lQV3fud5cwZ8K51DPu/a5PB8T4ld7x+tel27aaouv5aG4WmZDFkZr48Iuakx
1AqNv0oyCZVc6kSSVkmwvnswWsdS14+28FKWzKlhhMLkTLS9w7dHKYufYPCbr40j
/fJEDANA9QNMR6SsPdXTZ94EpY6+75Das5kuH0icV/+cvX7M2Tpkitdb6OX6YuLq
rgmQySM15IEa33NZRcrVq22VfdeOW+J6QHvd4GdszWGBJWXX7QHxktY9+marR4YX
Ct4xASel2T68X5UPX0yKRY41LcfLmCvcYsvAt8BWwS4ic8RhlDJqzyMq/i2T9rk9
1HwpDwIvdwZYFGYqwzsl5Z9VMf9E8WZ0PtaTmjrbo813AAqOl8SSFf6VnqN1EELx
sG+a26iCYR/yLnOqCqSmSA7Lrh/yWfdeWaffhInHa9FxyOUDHI9o9bEUicEWukcz
H8wyMzsIWKN9WW4/0eS8m+614/G7rURBXnBVEA3XXNQP7zjAdN7J1o2i0/1siUfd
CXWvZfKkDZje9mBNcBGLX/RUE+AKzZevfM/S0Jr2esy3KBgNN0pPPir4sE+Mg7Xd
+U2wWDYkQ6k2U/QwzdTA8KbkueLyIH4sOS6bUcPA43OM1CanXCbHKD1PbOPFNYUv
eZ0GRE8lXkE9m/w0VyJhnkGTNTvPJnr5IsaylyFu4GvJsbU2VR8ZmUf/IJNW0mH9
i5/OdxWvb91ZDHY63gGlza8VP6xc/LudvoOr4kGDPBlHmPVWpGvsH4WShWUuyM/T
8P5jHFsS5D6mhdoyiX+rX8JTJINIK+QlbEEXIQa3i+vTJBJ4cupm/X+MQg91kFCL
kKFdLm8qOrAlnuN9Aj7AR62dTcTN/UnLDiH45PM5iIgTghaAUpNEaGv5891ulanE
CU19dcAvhsOtvrnEMCjcMJdIegJfW1uDwx2NQwQh8ZnEirtzQFtZ5mhiZliwx1mA
3xKS078yiJZdj0bFyjRc8sVmOkAkcSbVmDi60NEIySpTSc310ib7gbKb1WCZ/3AR
ftYteqZfQjGJ3PxAa8kJrk8y7OK6H8b2rpX7x70/WyQqjyMmAS5/yHJaKgO6tSJx
3z3BoSFEItAvDzvQBBWOK9/tUAvWgDZ3K2l2CJ96EmzxNIotcq3/yFJx9MZFneH3
u8zIRC3CV3WLYaOoTIAi/fTCEfmww1szhBpTRvbrL7DXMAmJz8V4+DYKoRa+uW76
Qk335Fd36JfTUggQZ5pY6C4plIEE4VWh7gL7LEUWYRc0J5AF04bSRXzwabMtHPWi
7jPra2a/UCDW2fNz945jWdhVpUrWMKQ2VmWzQwvajnVIQJCx08cYwUMN4aWsp0PJ
B+aw9MGWv1OTS1isR2pO/xuL+HeDJHtBSZZn9t8HKS1mD0fE2exge/n1S96PG8j/
e86h9Yd/r+GMZ/wLK6XErWpetH5x/I9Ifc3MSU+WSzCeIMRere6JQnwne4MlJCDI
PbZ0hjWDYvMh5pjPWFmq4svNpNi7scvVVwDrwBvJ2+jbXgYi1sHcfk2zsOb7O6/P
COBdnpoEAtJes7Anes/Br/z+XVFiflh4YI0Kd2sZgUHKxrA/5zHhK8MApiAq92jW
s6Qd7kCP9WkDUZOzmVGPujdVTdklP62RrQf7sMaMnlOLx0GouzaDua14xfRHzDMO
3Dz+G80ITNeqGpNnnj1BaQIDury0xvdByyPBxyyoTC23n/gwz7kqunm7LeiKs5Dd
Hz/ErbsDbhVJQz8rzwWYb6pQmH+WCWlkoiqRScscLZaHrjASUWHZ/K83yz4asFML
9u/QT26La/CMWEgqewXkElQHpGG5HlOv+ILxy4yh1aWA54gQVwHLyxf4HSLLGO06
ZGFVBMYDcnB6JxGuHk6Oygs4K6k6Z2saM9bYJN1lQSrY4/rCDlzg+PJ7j8m5VYWy
gDbpFPi6d8VIIc+yl/jpCPkmyu5AINThhkJ9czT/mm6WSgIjYtBsrA9GdzzMHigy
ujinm/J2VbVaDaQUq3uXvjZXBzBx+d6/PH9q3B5qRdlgdWkDyUXNX2NSCiZJbMJp
i17sIHEwnKi5dNYvqNHuUK/AnR5QsYt52usywubjdYU7h6Xw5Aa3kdXhHlGoeclK
oQmp+ZKJANc4q4mnWJtsPBgkKR8eTKNOec2BB2P5VF1QBjPkU7Afwi6BHbA5P8JU
cspz7utxDvPlZGC/rPNiM5KsvLcVzgfhiHxSu2LkO+HlQ8o0jpHSynaZedkE5aSt
hNVdQUYfJc7SncypczCZYIP8/2HrA1/R/gSxl6sh76RvCS+oJQLOuU4I+KL4/0aV
TLCpul2FxxcbDQWNsC7CTKsqmljLODGX1CPIX4r5zGdahy0J7gnKprRkqNY/wvIL
8McHB4e5FGfNH+7eqXDZnRnoEI+gPKNWNT/rmWLqtq49K8pSUmm9j8G90ICDpLlN
TKwWFFnB1hYpDt6t6j0f28s3VyJLf/pWxfcCbPiACyhuBVcvb1Pa+44aHmCrT884
OU54It2tr2NBJ3vV+FY0mRQSkMD3RU1e7Y+31XUZvwpEYQbTCSs/6woePenJXpTM
N0e7CweLG1pQN0FWgYlBPcgxav9EBBG/SfFfcG8oMHq56IFmtC1lfU31myzSCGDa
+Xj1ysGWqw1AtuK0t9LQjgzAFwVfaICgmAC5yPWeCLAAsvlvxXcZKa8ocTivB8mv
C2UAOD/79dqFJDpTzmph1fssZhuH2XmpDpqgAywceagP8kwbH6HchYWZzjmiBq50
fYeWSoC3CO/6RRsk/U171/Xl37QAIENNOITILl6iJ1B6Om2XgqwOQuYvuQigai1y
y/v3wYR6AiJLubWPmjWWG9dIXoflXXhZwSNaTLiA9wEO+q8w1GwqCqf0Y0deFoPN
kjw924JZDsRYz+2SXRd4XDxYy4QmBYVE3YLMjqL6qIm0W2JLj+qnaK3copdNhdp1
Vvf0LfxgZH75GVN+VpX2eNXe9diWniIIs48SuYeAp9SnhdOXKG6/CPB2N9A7EOnR
m4g3L1XCI4R+Z6AifL57SYLSDnC7atTNuV/ki+NNf8f7vi+RnharTXfsM1CW2Plm
40kGxTmQEQcs4NUdYR/W73Yc/sczlMbuHzWAenUgyyBadExsGwRAfw5QIO/8NWAQ
sg02j6KmbqUIWbx/3lyHPuQqbFmqQpPx5zZgJkdmQ8Mv0mmL7fmwBemS5/mKk+Ei
hYYE1L/QWh5TGwCmW3aFaPI/fsthOiyglKmNVV80L7rT3xz3fhvxRMtfe9vnGR1N
gKAcCiDi1Pz+lUBFZt+tmawpR634wwt+5BewA0x2/jjrDoIQofO9FmJ/SjQ9Mfxd
dyR8VWZd7tad73XfluvpV1SbLM2rT0aR05hQCNaF+axzaYNkth4th9rekG37fRIg
fFARm6oML56pFp0hfWohkoc6oYHHb5zN7ubLzo/23kVubitserCX+1PAKv6FK4Rx
95VGodEl0xMwEdF5qF1VV4dYNsT9wUYe/v9vwBfDa3G2eozS/xyqkjBVmEwriqN6
7RagDZyF8iuBe3jsBvWX6ExpDwxA9ovFJpCc38ZOl45IdfLS5aCxk3FvBfIALZQp
awB2f9wpzuw+YwQtoSyh5t5rmmfTzn7/HU3tj/zL4fBVjaZRAoFyviRKxruPttOt
4AOZX96hRNcyx2ZeMnifUotPYu7fVWsxwqwoJ4Ymm+Yxl8YdF/vV6r/F6cFLU/YR
sGNedPTfr68/9fkebK86Od2dH4Cas9BrDi8lBhTsghjlg5z7q2h0kidjgLv1hrK+
bMKxUXb50bBm6RFVBdri6cTQ+L17bBXPm+QHJV9jrR4laLvKpeYPW4tfPc0i9H6Q
ZeTOG24ve6GpjQ/WV5l60a8pFOw6Os8mFMuDKYduyRx404YVA0ZGy83UnfUvpi/B
mo0CMBMm/mXBwTGI5/N0AowCCc9Wd+WxOJZeEJoyXX8Wy6zLebpNIq9ww8qYnTKF
Pv+1Un2APfZ3kC9OrwLZLbXT4d8gTK3vzVGaEfJRHa7z7ra6dLoUA7kL3cg5fPRh
0hRoq2jo0EAQOGBQFWasjw2p6qKxKBgVA3p9E9jiChThUQqwby3saPIfLK9I1es6
PpP1f/5sYybklK7epwTnHclE2MtWvfhLzkpJnfsLj2ul0yf54gn6egewPhNa4HQu
ta1Nc+eZDqPKme1ILHIyA2Fzc3kBYYGPB8NuwGxdeLpQJptY3ClmF25nhRtG6tpI
pRraRrtALrI1bJ5jl/1jjIkzpMPckdBbqBbr2Tlhjq/P6jThsl6EqXWnao3rd25y
90VWBoJ0zCVjQ89dvqUHRfMPF1L5xk/3M7wFgWKI4ekENSEcKOX23RcB5dvNmHH2
9jEiLeosVteU7kHyrZz/ns9nqNOdgYddSqjHdXs71G78hdy+3n588jKsT49AovdX
HS4ZFnHQFIFyCzBVUXK6qzu76Pe8u/3EIi1P9zcOCANUtzxhJ8uihVQT8rUOtuYe
4YIGTRAI7Lx+66vMyRfyI2ZWJItQThgH7lzWrL+M0KKnpEzCEQbuPtMWBjzSWj+v
J3SS0AP4JTVkmegiAHL5A5gweQ3GtaL4QpfvU4ozd+EtRabZtUxyGFMwFmMkWxhF
qtv+3oy7TXM/CydjPtE7f7anj9sqpEPNcF73i6HNJbO/pkyTPC/6fDnUgYe+nv9h
cC/CXef5tqjkyjY236BlCZX0X3zf8JFomx2oJMgA3oXPusMt3xEWZbFAxBRVQvQN
c/EqExcpXiVthFyg8+JPJZKFgQuVFkpR3+9K6qamLVo1IH2XOfoCpHYwiwZTBZOw
ooSj0/a06iX4KLX0MPX/oP6pDDQVFzSJY/yT9TuqoWKg0OtKG7HJfCgw0ZBnVXg9
JG8wM5AxWpr09ylorYzEsVrTXnwO1f7f3HNTUZNUlXkkmTrPUqKZAMw+hOAHeLRw
c8uLcmRRoZrfx1o6laXHUrHRn9FFFHAaq/q9mXNSno/b6fMdOKvVX1nzcp9adT/L
UQsVJMJnvgj7niTa70rx7m5ylRG4TzcqzfX1/Oh7+9/w2LPlaP/0QVqz3VcJQIu5
HiWWgn21rbO/jd21joSELDu8HPwXKFFcPKeIRbXB9yufCXwNogx2HgkQE4ewTPn2
6mWnd3g6JRg/004j3XSb/nNP1aNjgVcP0lEiGVLHpCUcWYo1Cq3Q9kR+zrbKUBON
wmKlEZUyQb2zbj8cmrTSiz4PnEbBE6r83+Htv39Qo9dbv7i1V+hOfK5Xxrp2S28H
eNvcqso1sDaCBp9VdemMyFdO6jMiKrFm/PORFG/+6UeGWidVCU+T0MhRifYRHuZb
Y9+zxu4ktjFU7tSFofWHlpZXYIW+EZlVuZNXJh8ZXACyLqJkFW7HhmylnWMyHX5v
jRLUNvQbCbAva9rRRtJS/Xy7/Dl7Zsf+GDOHhaw4WwsX2ueBHi1uMEtol6QgcRNM
HC8GsZSTv9PSZAE3QopfkVqJ/DHDd2j0FyP6V+sDHP8mChZ5daGNosR2SJVPNevP
kivV4MUn1Xq1RL5P7D43tmq2le+fj5pw4mofhbCYDmusa499syptnzDmLLo4oZvD
M1Hb2kQ0JZf7XjTtsHoJ1w0nDez5H7+0clxWIFds/naz/PuRzkDTA/pRFtBE83/l
7d3wx7FXnczqZU/P0BoptF6zZ0/8suvLUOtBQHx6Zy1VR+NYYQo2fEZnh6O8j5mU
DPfrkn962pp0NVlqsO/goioRlWeJouYa63hWI4SoNw3/djih0ygJC9iZjkyxZ5zu
ndmAJSu+6FS/pxYNBDbDAGdmH9/x0uJVquMZwiawFl85rfqtltNi8wcOxFFaspOB
MC/prvykcvZ4gLUFXDeHg6HbQ7ZRoe9zE6RtCma6a1OiRaCdUcaFo0zu3c4Lh6oO
PKI+rhXRWQ+sqs3UbY8IdU2XJzOOZJKRhyRtMqDpnqvieeEyhd4FB0gBTDSulQkr
W08ATHXiwYnhtRsyml0F7sRBFcE56VXiRPo4vbQzqMt9b1g7zPeQmUAqeFWZb5Hs
WZ9MzAEAxUN5isxuqDjvVwYVfgYxNSvnHX2zV35LjrInTVk1p1OH9/J1qatP91A4
OOzOKwMCxp7UEKesvsc9Z+iuQjQ4WD0EEHwVau9eJFeTA61J5Qu3RJgEr4MZjzYg
MBO8abo/RymhjCayaZYuSG3votgCI1kjeg3mTZKR6dpJuSW6Uo/AeYk2ULhkFINA
/dJuCp2jxUkaSvHxAXMrghCPA76Ur/+qjNdrR4xRkmgXsjtNKx24ToaVis3SCKQE
wWJKHR0wq2ZcWT7UFh/a1+TFeRQ67eh2yNMajjgNW8hp9CjcLzDo+ynyh9KAKOkZ
u+Y5CktJQJLLOpbni/klsFceewK9ZA6ikndT/PtHK4Jy61Krr1scKZWY0xwAe9zg
TxOkTanxNA/d1MLWiXN2sh4cFzMGGt7L1K26rnyRGvpnPWP3u1/pgPuxKpFFnmsE
UuVASwBpgpZq308KOoi8NeuDu5sdFp8Pel82sTVVsFsC/QlxQLNqMDZ6fQGyf8UU
ZiNxt84Xc8dMOQkDWfd0HIgobkbZ+RXz1i6ZzxVx/AycRwDfeN71P0jp3qg8fT/1
0MBGaeowmvzm+JTiqnBhx+goFfT/YxVc0otw9h2i0sqZOWaQEjUwqC7sahzTUUGs
G8Gmh9CiqNDn/Q2dH2F/vCx6hAGc1Ds4eMhaaRHDH2MsTa+dUZJq6oMbCzPEkVhj
P9BfNelQhCZ7xhKdzYc4ZmUcOHflLpi5AvaWn/9XpgSfFB3vtqgsf/280FoN+LJg
bfeG1FKvjVEmygLeshY0fgYiTQK/mLxPga0CaiAw6sv3MUEhxOejdyRUoOlyGOwi
5SRq0yD3brDHHCwF4JS/yCicUwPJ1uR0aK2qoLv5/+FP+NOYNKB6pcN8L9bDTz2J
6t8IOTGKplhYEo8bZY6J9fy1tyiAFIuosHj4LHbbXYYgXx/fQDMkr1gZP+YvJFjQ
yYLxydZ+prSYiMfdz9cvTCNgRD5WjVLJANZmH1EP34lRpgW13btdzhei9F/3f24Z
DusAWfY8dhGzxCDCcqjaJZy9drYfKhHlbgUVmA/YFHohoYtufZwGWmkwdngyPqA8
9E1rEaIe08fqWoC3i/qzG3oubyrsKRT7VqgAvhkzfWpYxauUfP8YSvcnckc4y3HM
gFSDbrj4CthpumDPRbuiSqDhKj5UloSPP1pu/b4H0tWuotvVi5l2EsZ4prDciliQ
sLafyzP+iS+DHKMJY8XdbP4jSRw/HigTIKKJciuhCYl6d9eg9Mvb1xPbdhEd7Scp
+ZP8qICUT8edTs7TsK96VrUFy45SD5S2AtDE+vrSbsEcLzgwt/UGSMrkyPL3zc3T
r04OzgAy1e8sOkhKBR7RrAyqJ45ohhMMD4Y/Uv68R9szVlVHDX2AYxqiSbhz2k4/
NvOsh/N1NT1z6ZA2Nn1NCtjhVtMNI3YhLiUSdYy1/DJdQ5nNNnn3PhUH9rruF6uv
mDHwgNCPDRwDtFXNtINXOzq5VCOol2pfvD1NAJUZYIkrtOG2BerHDqyWnoMZ8GI8
zxA+o4CA/RuTpUxARf6Qpi9Ntl/lZE0mkCDNr54o/bB/9UOPmR7ba2Ibl6Gtn0vW
5WVt9CranQbGO8OqpllM3GGbD0E29v0qcel/Bq+i6l/X5i3JTTPH82ursnfFybWq
//wxCnVH7d1Xi7Z+0wxFLHdKzHNETWuY8yv7827NU29tDEvvyDmyX1V0rnNXgiNZ
f+1jR2PXYnkg6Px/Yz+zkwAk6H8jYR3LqwAD2x0ajRs0CCnHvkZAUtryYVzx0gqa
fmwPx79kTcS75GleTy88Gfxh1pQc3C8V1Niiv/onvqKtQCJvhnTaedVz2nlMh8JO
ZILgLZj2iwbFtcD5Kk58z7nYQMsyjrsNAx0Vtk9KPKf1omZ0gKO6NTk/mQlqFEV2
CeKHbGrSBDDNYfC0blW/XUARpQDB3BIkXbo0H3nVdzITxDrmenUoTe7/1EReglFq
VH9/8UFdyCl4FbVjIBgicfpYYy7DgSPEULnUo4SQLaIp/G1+OkUQOz3DV5Of8ukD
xfRVP4WAbckuYh2WFZ5zhVayEoXYvYPtTJz6zSAlIbWSvKVvCA8Co9Ivz1txmlQ6
wkVwHUgcRUdPgnSo0oldfqG52oVBpDVK76v0tO6dhRwcWrgMGwqo5myU6BpBjach
MraU410OUiKZsCHKyH0mJ9WGT38H6BZl2ukxvC2E8qONZAhc8Zy+DOXkbgJRu4if
L6SX8r/OURbeCeCFnrmuAoFdNVRj5YGM+cRfaeLHczqNoRS0n5CxIAgbzHbtgLJS
inOETHQ2uDrR4V1WkXGF95wpNRK/fVuLvKLRSUTd/2yCYNlPYbEZWNUliExuCp4x
zMZhkmjQr8osTBwxFq7bujhLa9tLuYciej4QeTNe04NWHRktl+m1FpNWqss+QCwg
sJq2HF/w/+cLBYNJl6szDb8kq0c+zARW3ssfcswVLZKgQj8Di9DXYgeVEqVOxVup
P0XTOqZ0Z4IkPrXdEF8AqeGtYz9i3gDC7taFrHTyi3Woz0oIu4AWDMF4wzTsya/Z
PRaplhyowzyHHwjcB6mSKx8aP+arFT85m+uN42MDhM+pLBQ8DTLiw92JJsPF3y7h
HJR898sycjQkeeWJwKSS0URvqfvXzAoJ7pdMWiSt920jQN/D0i9iAfcClpfmtEIF
/MKEgaq68lHzJ4uJeyVBgfasXri02YpWAQIzyFvr23HfoEjFccaT/FVIsQ57Er6K
vH3Z5roseUGDZ/FKbjhTQ6H4xqkaDbUNA8WPVEDsphyWYCxgrw3D/vEw50xLR8ht
kigJSECADG3bBUFwdJ6ZwhgfgjmZHF8RgaVYLrkyJNmRVop9UcTUAL0g5y7C36wc
1vVtF9Pj9usn8wzW2T7ScKAcRYnySHPOG7bT8+0V/maU6oJvF4l/HH0i5fKVm9G6
VxBTixrp9av3tGLdJA3z4jZimyLRIgjepaVRMlZPxbjI1otBu1ZrTDfQpezAWhin
z7gm+E2MvfjP2NAKz3Awz1UQ5KO5CQqPDLew99TjnblAbw3rTTPLCOFNbf5R22GZ
vFAGuOKBT4a0ckA7UKdERdqUoAIIRkQDfhcrkUZrY5LUdQipIfH3m3K0n65OVD6+
MSNVL4Ksd161tMcdztR3Zt7kqcJysdCJiajzt87dT23QjIztKhHhORX0La3CWVlF
T3OYKf0wUIUnkK1IAYYYazDdzDkAbCYEUB5Um/gXOKePbzLtkdyI9Teab+19mxea
YDL4HzK03UUu/P4CKHjvIdBc+pvkwVwmMDJuDgIn0DzQ5jO3G+t5nbifHgbGFLBL
IF8LSnRB5pq2PYu1DvdoZYQVSuiLe4DnNhNXDlkKEZt2prgMoPofKpWR8DAkIBcT
eH49IAVkHtm4grrojNEjuPiB1txLHsKBftUekR2saKTeN4ET/A4vTZeptIGG4z9U
x5UBPTynHfu53E5q5GnKl9efqZeIBrETaxHviFBZWsS55IbeoIBWc02FxxWL9I4p
EOYFTDOH/XmRo6oLLG9cZCXrzT0JDxMFuVfKaaCiIa3AitdTW/sDHmm43DMhl564
0yWPx9T9Ma+COUV/qNmJ7peSBYzNOQ6bwXwTDM0fz4FsD0X/d2RHwewhPO0sPJxU
rdCb9AE8YCHWs9exWwW0PCXogLEyZxyQg35DjOyoEXc9BzHOkXNFuC1mCNXR7K+z
uiDp6/0xckULe/A6dcTC66nF5HxRtFM++ct1zxevXNP58waaeonbTToQNGJGf9Rf
qm1uG+a+eF+cNreiaFOhWNP45qYmCvky061APF4NdWfvnmcEwJyovnhqsdqcvOIa
Opl2Ol+rWzL6X1NlmyQbFd0VQi5fkHk2iQwCA+HB7VWQLzxpcajMof5MOSLpYcF5
oHGmGr5v/y4yU85yFGlGb/CI7Do4VTlDfiUUFmRGw9jRIIOaTn2EtE+F+nuejfYu
4UTYOsXB3DqHJau1PpXuQTBXsZF/9u20Z4yZa7sjrR0Yq5+vLHTqPhaDJj8jT1B3
gdJUWxXNRBLxtRyw50xryeMVXcEWrQlHWYCrnym0IEcPeqJMasy5rMd5vAwV4X7z
x7CsJ5ccNa3UjlZfuUypFHhghGPCuNfV3GtPcNCvl3hHawb/mlJG5eY5oaJg3kcp
ocfipPvg1xty0sRk8aSKWh/qxOHXfFQ117kny83NoHmkKRpzMKGS9C4wmXXnw6TC
JLw+KJPte/6Gpk9nYlfZ9PROd7yVpIx+joGKHfEhY9AgI9AC97ejvsu61PVQPwhW
zn6mwSAEw5gP1DkvQsBhrHZLMV4/2zWWKcwVIPtMs9m97S8E+TOa/BpCqF6p8z1v
buK9VKRr14pY+PAP31QxzC7hQ7an60cGcZnG5HUBvJzNetSzjCv5zTEy/WQn+xvg
IqRB5aNMlPjNcNGZZfB7ygKV+MPtF+IBpRAgp6u9+1UN5w2SQZSv/lMAVwyT4aF5
v/DRgqBqeF6EVDPzMtZOMeOCeFRNC/Ryk4Z0oyabYrD0hSN+i+To2FxiCEqkKkkK
iXDVjfhwEnq04EUt35KxvvmKNXfFDkKaq+8piHuQTO9XTy4UlORCmvJKeig7yT7g
wSf6PGlYHux2adNz9fEOoBOEeHL84DWE2A0ytXe+9ScVLwBE4V9fuAlnxFyaNwQd
g/4WKBfZywvoW0WRhd6vI5XJi/O5VamRMbiosCl9kz0/+fZb4RqV9lIWQdcw+nw8
a7IS0Q+6FV6THwBCRfafDXW5LGvFrvtOxAwfT6P0mh/Lp3RtZqvh0KCUHdkwyvNd
eEbtm85O3h5+2WL5N5OXnspENBDC3KfVXhOSEbrlPfAwU0tI1NYfQ6mQR6VOYWW/
tREApIFSmzr3g3BeJVW1rePalmtJXwLUfFQTI+IjeREvmDZEAkQEJAW/eiLSZjbC
vSaIRvlczWTwFMBZjgstHyZ7z58W6CJRja01R+l6awZNSmVTpfoAgbGBkzjyIS3l
xvFNH4rMhqD32yqXy3R3Gs6CFGvf6eOAuMxJkjW8/Rv6PER6ttJd2euLvepkO5fc
jF2IhH56c8oRb05VOxf3igNP2ToipHhMFtlBtH199tU8JRSW2wiRmuE6ASYc3ere
Zr5NH/kf1XX6OMVuUyZNckXYu+1kmerAcwxjPItH57r2N7XcZv6B96y/gEl4Iz39
O//x5wfzfSFNPxnq3yHMlbS8BvzdLoTkbV4wUni0fo9IVcA455Ng+mio7LFxjqd3
1f8jxql2ZccRHaKxqDSLoH5HZiBJzsEd5Th7X2feTLgyu0pbElp/yV1ja+jBgrTA
sf01THNCcW4WgDUkBBNgSjBX6DwDKCOFFTyOMJlNZ/7/vXXSI0S7faHidquxyfkr
DVE3Dd3ZSXPLWer+yV7VIYjjuWeAvZ1LNgIhQEjk7OEyvWFMYbAa0Y1JdaKGn3Uz
qTLPQy4sRsEIvafKAQL3AY0riKRMfgAcMidz3ORafBjUdlGMpSKnRvZQgTm1D89X
/xcO4tYBte7dv1yza80rEODPNJyqsJo1USxPj43FiwnmwRNzGE8BGb5LVJxnBxD7
8UWQ51xW/mGzuU3l1mvIB5JP1S/bsFM+FUg8d/Zu/TAIuH30wsd1RiUdGWnRmI8e
WZH1E8SUQExcZbDHy/NHj/4lmg7KHvXvNlqHFNDKr8woxabX3lVyXV26EivKoSuF
Wfho+UCQgNONQJktNV06o37u6uvNJfS3iprN2MyMheu/UqzZ+IuzXT8ZFsgHJMAo
fOlb+nZ8kUJQUVudlC/9rUQCfUENbal/ZBElA2uDsbFTEZh5hWbAImryaQWxYYqn
K5pWjnZJKwH+z2yewjw1KNuo4K9wUAy7R2mDPd42vCV7odZUZ/wgJ48XiwwEn0FV
xFRZ1D21ibup8ZF0BC2A8CCte/nvEvosTFtdCRaqDIDSd/UDjD6DO8orXZnuZ/xu
Z17q2Mw1mO6dZLl/El7cJbbQjweSib2Uj5YyOLKc8omMnu7bYFYtsazYDMcv5f2h
Pcraw9Fyi0aQ1q3zKIzYuk81NLCCV1spAI2seE6aRVCENaFQPbGLOfZ1cJpdftIp
pCoYVcu0bu2LZa9F18yQkk9zjSAGaXNOPtea3kD4ImlVcbrDlYoNJ5PTYwagiykJ
aqoT68FhJrYPK/mK3SWo7V9sN92exn2UZ188BaUFKsnLJXEMmwlXpCkiHFmLsHwb
Bsv9/cjnlMoObxeUXx3kXBrmqUcUIHQwYWVWsNb8YPllUipgjAHIemJ6fvHSr+/4
vLDidSj4Hikj7ZeQyfHs3o096hGSPxcEEAINrVrc2Xnt4KCldRiggVDjn5Ma71Bq
V8JjGd7qtl3hJuPpAOWVZGrYyIIbQozmBDIk5bkDvOS9nVI86gO/FuWIUgu6+ENV
ApTrDdMoNg8hBa83cA2pYd+3x45OPamINNUeAKUnw+dIcXw3exPapWWJjzgy441i
7IoP5ehUZmSMtmv8JziED5VUVrHbP1+52J71HnH/fv+UxDIhWFpXOxJ4M5h1PLiK
6jRx8IMa6gZ2jgLwotlySkkyg1TwUtVUt+Vrm8Jj5wm/bRA0tVTW74/mUuFuYism
SoqemgNDUCXtsYr1mBXccUZt6f9KtJUfb65m/H+GhHy+9xU9IwNsNvg+hWIMg8jv
F35fqVuSXmS8vzU98fdOUImF5AtccMlwfb0eyGnrJTko5N6Uz1HkmiP/0Mjw8HIK
7Czgo8kENuCNWzOxDy954kxgqW9PHraVQcubFijT7lfFKxhmyrGb+zqNNazZ6BOP
FGmeMlTc/O5llc2M+XiTOl0F93LbIPgZ+JDtcFvQeRltKcCW6frVnJaLIOD528BY
OOZsJwG3RU4/2LXk9jCUrHiwe0ISc3ckq+57M+0Eha3m7dC+VtKG2xBt0KYZakMn
h8zS39G8Xh1Aq3qMxFBVWSK9/CpRMHiOm8PyJDdLwB7te1MzIqJKPDSZfWPOJBd9
dCfw3pdolc62xD8kiDMDiMz0YCM20wCBg4qpnTlHgDFkocE18U51XOFP8mwLRpp4
iiBY14Y49vpvl2ki8yDtoJ6zRPNyXL1/wjZhjKH1aBSZ60eVmwpOIuZHCyqrECce
N6n+usZP+FdS0ixqIXsLMWrjhw2xxnpmUyIPyNFAF0fODIUFOMkzmaSQKPJpoHww
A+bMgcGOjrKCda1F7dPOasZvSBQyVcWb5Ve72HQVVhhWRlNBYNTd+CEa7vTRj9dD
CVbVy/ilxIvEoC/W22qCV7AyeZeg45tJfGdWoifkVJ0mfWBJMnzrb23n9LIODSLH
1ykZpOL5lbmFo8NB0lRG7hTgcpPQT4NLZB2XxwLuBAjwtUp7GhIGgY/0p6nfWXNg
sBLVoaDCoX6aYWK6TgcVGSBVFjfRPjIwBkeOCfwg5Yexp3cOCSAFo5Rb+JzDd+ny
zhmvdO4LcRO9jWR+CSBFh9sqBNLFt2AJJsx4KnU6/KWN5pZqJ1IrlYF8wavl5RN3
l3W6j+WvVK4dsODdy6C67QPeQI2IiNlo/yGIB/sE403+ukA8YDof/7nnS2NiMTCF
eQjI6GHW/1HIM//4HcqyXZbPlytgZtQMq+GvXNyaQn4UHaa03N3ReegkhC2g3V0q
rqmU09uePVqiokgcPQfCUbx1Ru0xk8ZZsBE/oAoZFtYhRZRvugaqMKLMdH0jTquR
4Id/ljKu5lyZm47PJISswk+sTput2z0jF8ju5Rr5GqQaoYoRrL3tRLTqq3Q4oZJP
ahH+d5WPnl6gIYwhpntiGWhH/SAR4QtWuB6vrb48LaHQ/7HmqlBSEeTEuVXMjHJi
N7h5g4Cj5v0KiWA5Fae1wGD4XjL8tymQd1jDLB/FUYET9jbzK2oUx/fZDuEJ22vr
yONbeRjC5D27BLh0h68EZAC5JNV7nKg+ft2BH8cJfnjIfQ/4tgywmZu123H+jnNh
MebqllOocQOpZnUmxa2VCA2ZfL2T5r+2aBniCuNgusrgzQ94vaj/VA6rgAKjHfj+
wwtHrxGVo+/CjF46Lap5DmpYVppmzQpx1hn0+p4S/TpCBpl7MZ4nQrD9mCqQEXco
gD09E8nEoaKxIUsg/mqmVhDSX2ScJjay6UaM3quyZNnE/Z3TDX4qZPz9kmYZUZXc
7Yr1s1zDuXLfywKHkXfOuYfrfzc94Jv6skiC1Gzm6e1etNuFPdGOpZmoGMvRZz+e
cmhYLZCchbAJXwXUlakKZdxX0LRms/roIe61oNF99dWtvppH3moUS6JxdpuzMMuj
0WOaFWopZCl4uCmv0VbIsF/KibSI9/kTPVbhs2Of9YWWEZMAGs5PrUH6IjW/R2/C
XFwKsG6Vpfj7eyafsSZblGk9fBUh6AkPbhQIYSLIydPvpgHTpa0KY5PBlJcRTIS4
/KWkesbp2h/ME0PXrEqVKcnhDV1YjSGMwz7VhvnZOZI1eGBCEczpFH8P5xDlH5L1
cxfboFwy9xfigSMCIh6KeEefqzoLmD1KmU9c4cYznBs/wZ3EplimEa+6jE8y23WK
XrY4Cvefleh/RhqqWD4gig4wmyLZwlAkJt9FdkKSFFaVSp9w4VJj92rgr4vD8Cbg
Dhpwzkg7qVMG7cjIf8PXBiOY2DHgPZ6DamWef2tVY/HnVMm8WoOthWBaPVDF89A3
t3/AWDn1gCPXkTW9PPQEgEvn6q14s0rXJqhB04eV4Y+7WLlLTMKaBM8ukZfIo0YQ
xRquM9rYQYAlqUAYZgnkesSmqGpSmPoF1lfQic+TNU1RxJDD9CLqI5yCl5pnoOFg
s4LLj1CQMWJHeQFVY58j61f2MfuRDZQgE1MJ2Kx9jL4Z58kMI0/0wrrrXGX7N5Ru
JqlLjOu+jbQR5ZVHQNNcmw8QNXoSdz0gbC7uY+UILXPloeztYqVKGSyABzpYDKfI
OmEb/gKpimaoFhVw2i1DndtCnv1fKHziD52OXRM09bKu2MGJiw2Rf9EwSH4MjALV
RooxNqkeb11ed721Wa9YZyZKCHSe9l4EvLsVQRSK1622fZ1uWHAy6zuYYEJTpjpe
XBvPVTqkOOM2ZnNdvhukVmdWoU6dnOOPv67Fu0brKgCmSe2HDceaS1OxetPjEsd4
/smCsBu137sLR/pW8KWO4E5W2seyO0e2kQ8RolOXinNAnxDSsddB1G/xWYglptJi
qpCE4aPpniAgHmuHcAt8vcmB9CinOhenSCksG07lbeR1JLmeGDeqmiGn8YQX3ebA
FUdHrkKe7UhdgRZZbAG8l96hahhn3vD2poVolLEMpyl8OCavuEGkO4GKF+yxcZW4
gp85lCR2z322lpK4TOJFFAsatVU5h5wia/ZToFuKraPqrF6V0alm6PnwxZuD6K/S
Omj3BKc3uJTQpxypiODOaLgSq9xS3WbkmZO3gk6Qd6m7s0MIbZE7Omr93xglyXYw
BuUzfJKpmY1mX6Eq4dr44jv6PL9sCBM0K3RYayqczf4LOqHYpUkTChjDwFm2L6C1
zUtRsHhBdmPsF8ZCaxra+ODWEXZplfhqCvkHg2SNHgdzGHSF6cpG9sJ48bi3pnaQ
fhu1agaVx78p8NRGfDIYxfxnf6gE6evOVmmEgf+mfVx3kQq57W1R0KxwTG93PA9D
nSTIOe44jYaAskdO1kphb0ujH0oqku17iaeZM5R/VSjFSIN1cMbs8vRQjwSXLsgr
9j+M3AV/uRkX90lmsphY8UZuHTUviRSqfthzHJc36QbXeJNeDrllVXdHL0Iks2kr
Uc1Q1IRUhYeRc7ROdI3nhkR7m6qLe9xQEjycZ7gLwTtjVnGs6oGsaZs8HB0u71vP
Mvfft5P+W3q96R2Mje6H53Y2DDiMUOZwFo1p0tmCAuUs16pUabo8Gksn76UYmsmL
OGUu/ww9PmqcSOEPS/WgPDCAngC+2qIMPXrw7n15YqN/gQf3+Rz2ChNb8/D9SvWy
lSBmK3PUkztvnIh6rUAu1BILeLX4ueMOjxcoqoTpXq0RsaIwgxTzCjeV1XSSeB8e
3qUZLGH+5gkxmJr2L0pDCLbp33thua+FJ0n7K6uUvJ46YArA/t+CvXsbemcuo21e
ctPX3ydqZS7D9vS98PHLbwaFOfdoMAGgO8RkoIkwEvgjCM83Fx4UWyNlYX848Kvg
U8V29i8OQHpe3zEcIsS8q3O85VN0Wm0lc7IQPR+zUhFHfFhsPIQ9w3oHWBkhHOMA
BLUyqXxV8N/BS6Qjl/hrwwSUI1Uj6tmhQUXZoWKal55R3fNrK3eVBRbMPJO4wCw0
tTfZgrWi049lSECqrl6PnVJVtc+xQbCVi6pL15TIcwqCwBymOgaG6YUU43RWng7x
UAKcYezekT/uWaDUXkbW/8T2c5AV8D+PLUJtZJ9OHVllEANIJVl35A5yNuTF7gNj
`protect END_PROTECTED
