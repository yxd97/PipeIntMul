`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHnB+YsdW/wAcjJumo5Zm3GaUXLEBlcnhm3ngOQo5htjhYjRM+Buof21vHXGtzer
l/hx+pwUM+QgB43cmDjfYWnhJ92SlycyXzibNjyLWxap5aCg67Q78QjfMqSpaQqv
JJfLliIiywNRXZTdIpQLHc5M5G0C1kUBHuK30gJkxbftfbJUkF0z/GNBIEXzjCna
xd9Fdmg/UMBQiQm5mBhuA3H2Q7xCT8bx7JnyPxQgFKhK2iHfJ3XowEtNgq717oV0
zRnw89Qd1wLOvYBfcqXhKs/trEzet137mKZrpmiURHnjlI3SzWw2bnY8z4MOMgp7
QaR6WxYSvgq8N2KfLehIFSednctxjrdEhyUxeM/hw5Ou0vhDCmtlRs7Gs/G2iBSr
/GBiQLJhwEyOFihGdC6Tsl/p+bKj7HK/ccWSoH/lRFqg2oPSiX7BNgXFZaKIZnLM
hUIoHJGDUdhlVKtB+8YUMIdFqExl6RooDJLZszcpZdht52iLSrvBzsZimTa8kKrF
Y76pqZ9DJC4Q6sf/SlNJywwqF6XFTUea0lLqplcVk3UGT/Khvysimj/Zt9SuQwSf
ESKdIGmG3KdN/KAPsj/o5sBiFrtSf5gib7ifMe3OpxxccczaGn/tZ8snWAdC4RTS
izy5sjwNIt5cvZdPFQAu5HNbtbA5BTcsB42IWZOklNZBcs9sWmScITkGQXUszQsp
atqWp7k7MBga1zSX8qvCRiYzbouD2aXL6Bh0ltx5upn2BoHo6C/B/GuWTafnU7it
VgmHuXX3RTjOEpJfjgMP3uDfK/uQzwgmE8NvhXNaVnbuve70Oe2DkY8+/j8ZEXt2
r9zd/21nzl3MUg1y3rfuYPHUQdVxA6WzCByG5sQCQCMkI1n8WxHmKb5K4LPAoLrj
0dCoziff+EOFSEy3JkHDYaz4nA5qaUqpx76OnsfzXfggpwNBswtqBZw4wWrckCnu
Cwkoh5lkx3kyvmbnVN+VD75YxSPwCnJ5HA8+M4NDJ7v6tlQ7nhOgthJQl4LtnlGn
O5I8UZrG9wguhV+p3+6KvmpBAITZ9yZU4XgcXCAc60a96SIwow5UbRvYWRU2kOM4
MIsgdqfrof2H48DKr/vgRbFVyF4vwOiFGzoPveCMG3zCpEoO9JLR60vU1fPxJwxq
fkO+04kLsfWkTaWIliHioYz2PfOfB+q0h9t+7hDfGOMWyFBdA5zM+FJPx5v0omY8
tIIJl8qpiJ4I4KYWP9IHS/KWiQC+ep3v2an/0aAEwdSJ5+TXuPhUR0uL+g2RnWkz
q2zKkvPsT4Xc7r25Vt1ZoMJpizUOMq8MrTCtcnzJy0ZkrD+Tk8k6hwF0pi4O9VoX
eUZQEYIn7D7f8GtMY2dXtsOybz0KLsrlRbCf8gw8FGxxyXyUQIbKMcVAKsqalWrd
oTqbp3hLEcNHVaiBMM8nxCKYS9sBW2dq791Lr4eOU7neiU6mxhlIOl9VowguIyzY
wQe5915uEv+okXagsIyXK1wY3CK75DkBPIyRYMlFU6fMsld19dBWd6q4NbShnxgp
dF6aL4UJLt0rjqzj6JLgPz1tX/29l86m7VibDsWJx9eudtDY0BJVLbrDHW/MwY1d
76T+xSAVyjP6H7Q4l2UXLTbZzvB6iwzvnlkxCA38cDHmg5U1eWLhdKJ1vIr6JVmy
vkgFor1T4XvdEAenqo7TkaEZyVvYe1F3e79a1Kmpzd/hcqIJmfT2Tkqiki9Dppqq
EfUnkRiKafhq5c2cfe9ijSLVqin5eUrPi0pjzisf5S+9oeYLamnie40OqQMA+z65
ObmJRQdyecBy2sI8bVgtmNiAE0hJr//hJDUBGVIoTEIfdanKtnJUCY3F991grDK6
uyQMZLEkAag4Q3dbmvN0NcS6jN6XkZUAUJYQq5twKJhFBjhJADBwxYom3aDbdie7
8RTr3QMo2NgAUq1IpKa7SAYBi89rYO4cFQZiqpj42GimGXi6kjO1TRNW+pU0+KDz
m31SIgPfBKfzMRmaKymFM1nhtorXOfcgXOkTdVCGluqDnHdBCGW6NogLiqqYutUZ
bollALia5Jm5eYavc6e9bCjUMYdPGOxEbrRbzPl+Gix7I0wWFb/boDvT0nXlGjdO
shKNF4WtcxOyulTO4jHt5Bin9UI4lb5t2a+6scH7Y853LppvCew2+4bT+OF/YPKA
Krg8OyNiPBh/L/eDj+0eaayTX9HRSFML8xJqbYCDxCkklvHPZ9v3U2U3goZ40bF7
Xp/wVyFJ/xOJqbjhLASnBKCpSI3eQaRliQyGFTt7dsensgaGPVfpgSXCL5wW3dOl
CFomF9jIz96TRPzjpv4RUHjyhVQe4APsBbpz2sZIjM7YmuzQIwsKl8SWQtg1qMVJ
8gkF0EpmdHyA2x/Mo5esLBoZ9Ccov5IPtBHvZkCshBc6cUnEtI3NZIsGL6qfJPrA
S5EFANXLILeVtVssCKVxtfdL1cyrdTN5buffznchac+wCm56LgVFpp+EDlrK4r2/
MtVT4wWSfec7KZ8whdfbxKS+Awf3aULnePY6xdxpbRqEIU9IKRpLhHlDKTwP50L1
KeUKKJsor/9/6KOfPJYvXN/q/qfRP6YJrFb0Xo0By1jlSWyAC5mLxDgODue+ikrj
9DFBJfRcOKthu2pERfmL6RTLVtXSdo+Ip05yzj8xlXA8xafS+R667cwSDpOPL1o/
G/K2D5OlYpqDnGvLMh+ID+Jn40G1f2FF/dJIkGyIILPfMaYsbILJJecpG2wN759m
SoHd/UGDQmTL7SYuLKfzov+nfG3iqMAYGXCclP9aLNbfXCGkLJ4ObXxt91vVF79q
QwSf9PwgahkXp0X1LmdOUMsYgDXbd/3xPWddN80PzpJLkSKk5BHgHpvaNczaY0hy
HyK5Jx24zoXKrfjT/B8e+5QswoFScOztzAkBkjeyH4/txZjFu5lX2w5ZxqPnBqpx
vSB+KGVgAi7uAlXQ/gyMEeGkRu56bLGr7bKi1VmEwuwflT8HBFa3yJ3+jKo2GyFW
FUaPh5+Eip9FCkNeR3shC+w+ZGr5t4bNUI3nWE/oZWMqnpXxVTeQGMqTzXzKCDEO
qQ1r+13wvN1AzeffKb1jemtZuwHKG/FeUC/2I3uMAvLcnlKOpLtxDE2VwwGWD1BS
Z3XkAZ+4MGpqUAtb2GOdBDDkuj4Pn2C06H3vBJX1W/WaRld2SdI+lVPPOHJWOAMB
KAAf6WlObf8m9BNFaeogqrOJ9qPgs0mtxSN7UQQZfpieyifXA48jJ/Ca+PVJtCTO
KutkHSBtejv5RSuRbFfCu/gCFN2Fwz4fIdNcBK47ZGvzYHD4L5HRhIL3To/OcBdP
X4QUt7UCERLO9XI3uMtDeYadCTF56Cm1/l55ajrNUfqU0Mj5L58PA/+cSDlqdCS5
gloaxm7uU4UjsueVHU4VnYg+q3tnc0e/0NBh+3pr+R7p7oaRL3fjijkG5qWhnG3f
vy5io1Ataq6Xvi4gYfpbwC5hsWJ/hVQUwdOItsoI/ungjlHU7PxX0QHKf54Slivu
U8HKOXGREBHuLFVTWeOtw987Zl9b68wJlKbJxMq+IW/0d6wcISdQ1f8rKFfvChCu
gBMi+ahOfI127raRVBW8s7pEtfUdOhqWKDHL3Lt+ZLtXKDt2VIkSNPIXu6T1TXPJ
PXdu7MrXWz2GjouRXEUQEI1zCTaeCTusxDhxV3+b+BYlbMU97KS669fMsIQp6KR5
NUuO/fKLSlY4nCBq14X3Xyoy2a+dLpfWPwkQBpC2aZDZyw5aajoWJGM7yf2PePAC
nqYe987R5MhSvxriTa/b2GNN1mXhfAy8jffYmdKMzd4NHJimUqcQMFZ8Iiw4dh32
LiLh7/Y8EZq3wMpTSpGia/7jn0LB2/YlZVyqr7LUeznnvaIYRYfUuM5/cNYfeLmG
RZmOpiMOZK/QrGxELsaK8wUKOe5WQrlVfwtBrDNtudCLmS+aUzieZ+qvpfrBfdNh
4fFBlgKLgHv0mhFMUlCLXKnZaKYrdEMtmJf9ayuhApCb0I30VZQSxYV1wwpmnltf
qk0F20KMO6o3pr25irq1Rm+UTEkf9SfhPXyvK+TNFVpvRWfK7q9d6P474ckF5+1g
npYC8mQU8r0PTWdDwQvCjJpV/S77rc3WZEuAh85Jex6umF7MZ1NYKzw/mSU/u9jo
5Yo+F3Sbg4Gs23DtX+OM2M8ouYTtxuezxQnHWBWYK8gcYpVkUn72dmv1aJaxmM6t
CeGqDBCRhE9CYBYeHWzx01/2p0Mtw1+DvWHVbZpVOm63YnVJVbbD0tGrbcoHOOmB
GgJkB0xA26hHwhL+NL+Qsi3FGT+F9jbCXxCP22HEssuRfiZGisjMu9B+7wIS2A00
Eyey9ThEUOQvdgt0EuyBEibI3KlR9mYJJm1H/9T6piBs4jYfRreSbnu5IDSoqKVv
FzGzDEDshnqA05Y7Eas7bQ80yxt93+jp9U18T9pF8sYEzw0+1ECA/qzedjryfKH0
+BXNU0jGKIrtpREGXyFNDYSbOebd8thNN4CSyMc9lCYdqly9zxN51mc4vkrnwwxI
o0A0E+Cmblvcc6e/mYTKK95vf8jeM2XggZGCrliSK0YgoLogVXQ9xWUVLCdadZbm
rKPd0tXGLcOzvksF/TVCfLglubqEeB6M2W6yAZ4rAKQaRpMJ+c03lFJgMptgT/Qs
VCrA4jS1Ooc+y4AUSAzWr7G8vEs+/WOhJJuhQCRkuqW0kLy8uM8s2ER31QPTm7Ys
6ZkGsOuXb1OfDE7Bg7SZUKSk9TJTuBRo2eLxG4g/k/JmGClPwYzqqXihXvKK7t2I
D2B3ykSWXMFWTpc8hNc+fuLjNsa06v9TMMCrZ2048jJ4oeTVM3rPpMs0wH9Y70V3
3j70jyc/00cMg7M5919EZ6YCENxC9Q8ZDzxLwB9HuhsXK41cp3dNNkLlz6bXruSg
qPMYHd1XPtzlYY3EyfOqLbt1Me7XnJgxBkKEmYPoP8E189B1S90i7bIkGbAfp1QY
acmDOAR7QSDtri/k7MME26tZt5qszyN8Ghg7OtDGPU9YaNQkmCaS5XP/c/oWVziQ
rZgjz+H+c64F7HfOCrmYNN4GSuFy8IPNPeXKne9kcdmlaGNCZ+7cNZOP8yW25dUD
zYOwKugH97PmboEje4rjcOkmwZ1Pyx67Zsx7/QHJgWoj6kzx56h5nZSCTMFsm3yO
nRbQ8lXOFM40lVPaSzqO55p+ErANURG4uaDUvzfjmcaz0gzk4YovTvhKIswa6tQS
TnU7bhOvY9ptv6dzrbRCSGso6K4PH7fwQ9tTlqbt7rgRpS28/M4fMxt3mIHtRkrc
C0iK/s7ZOOotlArBex72MXnn/pX56E//tH857zVcFzu4XXlEMVEgTd/oaFXQOLSp
Myx9qG9Z9dmBbLWA3Y2aDmeaINVtx7NXuFoNWRyC5KD2HHmpPX4coA4IHg7cVDpu
NcTX787hI1S1Lcp9c36NvNm6tol0AsSSHsDHIhhADIvyEOWaS9lcZ9lUT08uK1yN
raX9xn3kIhCkylTxIWmtaQ0ymZGclzsCrp2IOu8Lrm2h34vQjMpy8AiqGOm9EkO4
S03LRGA5zVe/TucMxcXby+CemQEF6nCi51w7b2paWc/JgnFFaSGSBdT+GL6PGGJw
0LMBMAHsh5bq7gzMArc6WEgtjXqM6/G+5beWgHRMNTyubuv5TzdVokFt5swtRNxh
64i9kataIVxT4s7M6UHAiWMrNSQ3oT4IwIQhu+Zoo2XqVEth3GO0chPPpwfM3D4Y
qj3rMRAsr/WVTESsEI+8Qbup8IVfa8hMeZpELkeXisGLLRDKu91oBu/aK37sSuBv
CaO8i36G5bXmhOfPnutLV8QioaBpheLpJWtJUiEZ8kyvJ2ZQZ+1Qz5ig0I/OaCpv
1JzV0kxJ9uybiT1FgI1zCOqecIxoekUyJUgf6JxqDGXAXGcIZ3kl51h3ZF09kQNZ
dd+9thhwJgimYOOPkX195lvQFOtGSt/e01C+Aqqmd2NhzbQKuSK8Ok+o+ilLGaJw
oyloWWcwTiu3HaGoc5RYceSAt/1QdEHhfhQwO60v884sAFYUuk8rcytSfo8HPB+R
WoiDmvFXHzp06hc3kPdkGSYMk1YhYaQoZFSoEnSnjM14VK1DkRXBR0WvIXd/UT9f
ZoW+BqfTJ7E8UMzXB5L8geFIdrSc/OJPBVoxdElaUWJjCQNSA7sT0BWeNsX8fdGj
m2EPmzMTPS50xu9Gn0NozYuEOMYxvV9PyolzGVSkiELK4BGsUZjQvg3ZGu3OtSjN
i9Y+1r8r2N4FXAqrnXLqQsXQW9ndCCZAFUAlAWSlAbBiVP1cRHT/LFS5XdTseW49
orXX/Yg6ofBiNEysYQ+/ibfZDdb+PGrUKtEPtIuZ1dhRS8OShQ3edYvbwJhJDzD0
faOmnBgwqRxqS5R+zlbJP0OXuTtN/weQ6d/LWLv2Bm3xpz5Bx5V5CFgbGMUaRwnG
sn/8lNFtQDlfYahRHyXiacrVFeTyxY7PdhWYWTc+mHuaZyysxo20aDRS/vKFl2z6
u1LsCqypSXDze2Lo5kROqd18j3HT55aD+e/gfrwhrfEtt8r55MKjCKZo2VNY+e+9
yOlFecoGJyJSfYD45xQpFhYkv5f3KfmrX8K0SHvC6CI+pLiM5i9aD0D9xC/7S8Mj
SlPk4IYUivxchqe0siPsX1IH+/gfD/MMWMJocVdIKlU1uyAG3URWWReyXBItff5b
cWE0IsSxScqNOxb/FjR9/lQKajSKsQoqqF4kVZ4fST0mU42CroTDq+He4Iwz+FOJ
fiXjD9zWfMr5P88e3BlnaVZaBPsD9RHAciwgMjCTP8q3gBcLdpB9jnIeWJ396yGg
Z7vCM+EF3IJhTrAgqb8TKu333C3zCaFzYLt4TLNN1MEF1GlsFQxf/hLvB7g2wLJh
xFMtuQV5aex1aG/ucoJJQ5fxwptqqk94gHEF8eHs/CL96C+CDq7vI1Lu94lXLE6K
IWnXeASQUfoKvuFhTI+Jv4+4nYZyfY7dRWQemKUsElin1tgqA1gVeCqYgBaHpACo
WcleA4YRQjWQM5zkfU98cJ675uBq36c/UrSbbrKcS1dgy0pIafk/hTtUpDZ0oE2I
9wXrXPwuZILnvd8PJWbAZCto85Pqv/oGGIQLXvPRvwhPJxUMhBNn1EO7cjUDtrrh
QBPe5Kq68pNjFmRRv/UT8sUN/6Zj5vBVbZ6R5Gi/G7+0QsBAUQsQDbtZciIda6Iz
y+ig/dqJbh8BdI+4z16tb6eLCO9V0YbRU23+Io1yUVIS4eiQl78M9GWthOHMMHvv
gRWv8oBRXY45sESxvyBnjNxpACBjKui/r065Iij8n+Pnckt/dx29st4j3GabtGeQ
t7UtuuxwKh4ZIkE3KdlXBJZ4d1Am7psWLbITBT0A6cs2V4c1G5Zw47MdURmtr661
N7GBeGGCTUpUhdd3138jug2n2/aa5sxAG3zKED9z6OgUVq562aYR22v9WMWe8UyE
tvouFpcIhEOaczEUD3IK1inNX6224yCLoeXvf12D+9l4N7werDPEJ/s28Zo1dAe/
1fhuA/APMYm4iHMt/ZCtO7rTC9JZoLLxCvl1xXEdWbxTscILsSMgBW0sODofwbq2
dV0kXa/O4GFu5ss7CIqbzx+ldQQMK0At1/GmLHFdTiHqrdK5izRiBEq+emd90kdY
2QKDmaB3gGqoh7Wpm7QshcIplZL5Eo6la8JuI7tlo3jWbcT1bbrH+R4jUxCXKDSv
Y46NV7T6dDJwJ2dxzk2oqciQWY9pWuO9qXMI8nJHir+cVm8a0cLRoSlPp7Agzhiq
+n1zYLklAX2aq5eZVjeIvsvglmfglyXQdn7/1S2F0NQGEhK0MvWxEVuFwRKGuLDV
HMJGE0JZ3DioUENKhMx/vwoliezOJOQdJGtH+AZEoQphhb1DDitEH7QUUo8Rd5py
nldtYwzgL8Y0CFnnSdKqpv3wCmo7zMCFh7C595CZ+EIsOsXDzjilDsPftYnooZQe
U7OmX9NAFHoulhdqdfGl4+JxdNYrFNc70BEZe/4ATRD778jar3M7sz4yIRkNozL5
C6jdLMnBYcq1gMJibLcxBGfJHjv0bEWaWCGDjDFUVTr4gYkAcNO0P8gqeZx3yAq5
rXdX86/gQpt8YRi2bRvXZ02xe0fdtDekfWEtbvgRJk2VWKQ/oPNkWgDYPvPQPJkt
ZE3EwhS5aTi09nRWxDSxpTtmFeVQ5QRS9OT98WvVhA1jS3iNQl6a89S0Ll0qNcbn
owCPFbAuhmkysT0iDBZ1baAe574obtuDg40IIm7NPEVLbMiGFmTP0eX5U8A/XA6a
gl/40SmaqfWg4Ks3SSQiWL6RlBNbZuKz1Z56tlWP6l4xmUUxty84XR13BHgJjD5w
i9Dsb6A2vF5G/J5hONl9FRR0zEGVQAl2RnHvNjnM2/x5XgkArpgwDqtl0J1Ey3Yl
s2Sg38v3QJEUDXtd4+WAqG1IV6yBDemvyWLbUomL3ISeaqpt43UWlrYoP7VN07Dc
s+c8WboSzfxoAowr/Xnnev6TCUSE4j1MdDVjnF9e5rE8/4FeozThJSOl8IeIzwjM
nCI3gId4dhwGA4UUGobJlWeogKgTLLm+D+oUeNyDl4JykgwmXjjIZYgs9if+hiYb
qa4to9dCdRnTKeLeuZs7Nr+Sm+67MqNVCGPlRHrS32sww5VARTyhdz8DmsSmqDnK
gNtLa0vUGj4g+gQ4xgSHsfW/qQmYE75eCi0BIuw3gFu9gohqescg1C/0D4kQ6ttQ
JrY8OYjI2YEE6Hjjxfxm+pN5UMW9XdVYs3vTdNiWz+LpmLI3GmcRY2cQcSBpD/CC
Js3KWtmwF98FeOKB8UCIdg+nDC+mW5ywD102SbnF1q/njk4ec7GdY76ffCx4G/zn
kr5lRVZNs/Nh4DsUImOla7tz7adA9G+aUI73ysGZi3HQ29NuiwRFTxbJUo+8CDl+
Z0iPZcmPf7GZg88ZpY7+iiW61GWVFB6D860WOwRrpXvdyi62xR9xvtXyh4I4gfjJ
EurRDm+Tbjo6MGHTdNaaCut7CzOP5uhdyvEmARuctzq+YSykX7MvpA4AIf+onKEy
qkvpChySwHr8SUzHzT2iMivlXIe+FVuuvgrVxpv1/pmDdmwJb0fO1CFUdpRRPE/D
Gdf00CuIArB3xBt6Q+aaeGoIPge6btjchExloV8CawMlTRveydoJGZLWRSJqBnG2
CPlMMuhG6V7RPISwTO5yc3vpZUS1QwbdQ8iGCZGB7pN3FHWH3ZcNSG2iuR3mAVNt
qMyO+9wj9Th56SDrzSauU0UhVrijE1Pn5zHuQlnZcmuWmhXjI/zHEvdmLBWsTmk2
i0O1bpJr6tX39KmLXnEvdxrsvKbvftizFkaP60UZLob6KdgYbYrk9zOzAIMTUEQJ
DkXElt7yNMOD5rdu3tf/sR54RU3SApgfBwmm0s4pyUjtp/cpanEMZZ3K3ysoiw29
votfupfBgDgSzeTiQA89bCz1v1R7AfMSfvF/Y3SkqtY8UuKAX8I87fBQEpXAnBuV
hPN9AjcLYT8TZTlopG6rH58Dm01AeWNb7kcFG2F31Vel2k3qHIFeXEWvWGzKyZfx
U6+YDbWpc0lsSql2vGPIiu80+f5Q36+rzuKzIFZ1EDELYKpY0huag+yuOHcpUEje
Tc1TeN82uw1ej5Tx+TB4ysJXY+ae8o7T3pj8ab80HGh/LhbpBHbdbSPVq9FHWfUH
zTJmzpQnIrIlqYcVR+Uy18GfKkTSo40VnQRz+pOjfWqV2FMTl3nuUKcNNEavVFig
Bn4znAL0lJEAUjtpqAUWWqGV2WpQz866Nmr15cxceVYh0M+B3KxqCAnCNJvO9ItT
qIL1Iz4PKPss0j17yxxaHCC2xVnekXTxpwx7pKNeqSujCJplkWZ4NWVsXtDe/yAs
UC09aYYiUOA/o4Tlap4YfQJ4X9DDaKgOR/TJqwIkRiT7pZwC8l8+/++o//Ei5qzP
HjkTESNML4g+QqMnrLYNctTL+Yny/jEWkHZAj/uZiIlK3FKSBed1OBkJooXfNXgY
C8SHv3bphQXtcETopnrq0L5JoMeINchoAGUulSCv867gCkAfSV7X8uSMEuQEguxV
Tvr+mKaLwG9sLhOF4Qg2KyNwDqMixRzt3r3riZhsM6JWQCfeTQXaDcZs8We5qgSk
QhSGNbNQFQ06Sp3Iw6qFFr9u82T1VFviUXKyxJ2UwcLAIiIVvUJcgYpP2YVp36mL
T3SfZPSlpmQNIvYS1J+1gqYx+5HYahBhAlcWd8Yw4ehFhDCJFOgwond1tb/713p1
jjwIuKmKGypCDl4en9ttb+wCHabheJn4/ahvaBQHFlyEc68OQ5/VS3QbaoywrQx7
hK3/8211xwksXCeTMd5sP8aOXRv8zcszEegfD/RLE8uCogUbWaC8apaI1PjOXIN7
ka6DDDe2xDSh5wCI83PO9MadTIwY1B0ODwoHolBofFrt+2Ep1xrBD1mWjSeGS7EO
NuFNbYY5imVLq8FnegDeYYpL6NQk1f+RTzijYQx6MqemzonBMp9883ctPxxR4KEk
dNvI1/JM7OR9Y/mbrlFwjphjNLFGTysPA9rcLOSwYKYfxOgFN1hBaHnyXhthIDBg
PEC6WokBH+eG28VNKNRDo89TlFvy/xlw5DXi7xC8EZJot6S+2fVaHst670V0V/uR
A/nSecwDqCIZV/SkIDbz7eQx8T2yBCacET00v7Nlaih4WXG02jeWKkY0mqFvZ0Ik
NeaguNN8ce+sjALWUnL+Crrolgk6YmQC3o+8g4wRpZA0cly+Vqyn5uilhK8uMxaY
c5ksTK0e3kIonCfxiqVS1afRNVDTbAJXi2rRF8dLFs/f2y7AHvLFaIVVq74nZCYB
4L7jqmw9VA5UZCDqQktepg4dkXDnFpNw5r6Xo4XMHw+MtRVjZdp9MPtwXntqM/4U
ZyYF0JooYN+byGqZKU5xlWH1oWlH94VmSHJSQpfoo0yqbXMgqwWpOSFQyA56bp8j
onryZ4MHIIp1OqEYsqEG8oEUaBcV2LWKP8Apdu4sL6jlf+k7uzeDC9kh3ijITZsy
PpQMMX6tI+iiZDqalQsGwY9ED2+w7wHMvx22XLUrS1BcWnqQK0oKttSwM3iDk21U
CLkwKawMB2n1TAIbifD49LFhOwON2f9IMjHNHmHCA3MWv7RbBkcCofRBrHM9AZ7E
iVPItbxEuKvMgSXMsFOOL0YuL7fnl4a4xOHKuc7BbtrVK/YdZt/syKpjNeUVqNxB
78UVU0pnNe874I1VewPea5pn4DnwvOxi818tUJ0iWP6Ex3do9CWctVH9H5eWDCYX
ctugeg876cBWFJclv+xf5PrHM5T+lROzktNzDeuXhNtxDbYQqmdFaQawjAwvRnYG
XW97Q3lmXjTELQGU8pXQoxm2y9+m3i3j4Q1y1x7yG1cLROs8tRrH0qS5AWRfY7nV
bkKZ3E8F5kZ11E0sQTUk/MxuY1AjcG80jpAM0+dpe55cV7XiTdmGUl+C21ngEqKt
8pYTooBPeKK2uqH7J16F3vly7h0iPRWTRf2KaPNQ5RFYgB+nKXJ5di3D6a+w6jpn
0GbZOP9F08Z9hujKWURtvCFsMU5DRWe1N3wKPIOq27uQSFW6bGv0iTOgjhP2b3O6
MHmpwN7dw1ezuF7Kth6dge+S0cb8hYaPirdSDsRixMw/80HarYXfTrmS77lIl8gO
GlwH/HdWNao7niaNRm9dpxlleW2aAjZGMPXLfz1Of6iptf3CmW5Q2CTqZD+ZWs+Y
AZe2cwXLgjYh3ZcyZE8S2awyCnofPM+2xtH1zF6SFIaRvW8K+0ML4tx/q+SZuJrd
/m/nqPri8aAKYHOsHzVn7WBvc23aIED8V3qL4/oriRBMtqb7gAVbRXEc5cDHKf0F
twcfS3+affZw2jNjobhCgNgd8VMyIu/RFqDx98RUDrsj05UDp2yyBsUc7MHyORxq
A91q1HZ9+PGh9g+b+rxaEYmyEcZez/MtYy3fyTIgRDRvAPn3l+3tlUzZ9vuJmiVf
FJVinMeKmZrsZyjcZlxZI1yL5EL1e5bstEMKdWEYNxAdyRe4OBYJZVO+VffPtNhP
qtLUIKex8WQuK1r0iZaQQd5rCQJhU8AyMoOdkbB1XCvExHTeYEr4thz8iPG+J6l2
Ej+0zC4SKxm/c+2JeGW7yBCu2MTvMF3V24F/t4BYW2DJIOartGp0HtnhDzQ9dI+A
Qy4iGupXCuBgXXdRrwZyoFUS8V8v9/UF8AEg06fZmbEztuU//xJcLw+7QzG5RSIe
hVnij7IIAPqj7HU+ceWJSlJA7Pk9Wxs5I9ehISVCGXsdrYmKRJ/iGwnfXURZySt+
AaUOkozX7NIwvDT+j573JepsfYfV6J9F2yEDDig3yJ27+Unu+TQfA9XDh+9yJ4/J
TIO+QGhUEPE2SKW7xbYvvA0DwXPvZEvpeo3Rs4VGQJQL1q+q4RI8TtA5nBZ0gqNB
X1m9YjlTMrDGv9VybgUmCfKGKuGK4wm1xEIk1Uzc6ePwYhTJlKP3Xno2uFpD04ww
RoinYXZIMdZkkLUlDyQHgXwl7PbU0ButxxabSZWc8/aDUyLLk5iEVpPoUIic3goL
VxSq1SzMclNNgnSiihIHhjf0+yM6o2JPAINrBo7PhqVxc3yN1uxexSzp678WFBCR
RgFfLtrmGLD476gQVTgwDKF+9/FavxlXOhM9oYank0y3XiInAo+SpJB8epx1gI+N
gihXCZtlpAcMpiBUdNtoA/23IqWdHTJhFoBMNv5yEjgz5YNQ2c6i4raLbCcXz3yZ
L3RWqSEdP0Cg/LhR2Zzm28U960WSjq40YKHgOLYdp9kD8UZ+bDcruH/Q5OrJwYwu
Sa1AzkcsAmEEq9RA13mPUugekCyKdI4heMwCPuDuR7MzAq0qqupN+nxc5N2PZBJN
iPh7QFrwPUQ72FlZaddHVn8XtiyWN/8cfM2zac9ni4JuUOyAjyBor3dVILx7pzFY
uL31l7ACwSir6D99lJ7BInFLMCupjTdLzNWkNYRFhyIIqy75an7JdBM/RK+i+klL
gX8txr3LKaI+fLyB8jNW5H6eNU2gSBMruKuWujVhqFBoRSl1oJdl2Y6NHsy4gDzH
5LeQahzOZKXGeDZJ4cQvDw2rWN7SzVt1cql36/B0T7EX7BMx8CabAsz6/h/Ni1eU
q6rBETn8OJMKqXq3nAfopeRHhjgXh2pQ7gHriP8aV0ZHWTXFl76TyQHnMgrZa7aa
rRlXv47p2iWGeWKvVqFhVU4I1DNYQSwOoMOwst89dCAJPN5I0iHt0l2guPPmr5Qf
FtHPfY7CNna4uHTXaLCm9SQ2UwFOdLLm5HMnMgY9/XKBPl992GfVKha82rjh4kFH
3wohhYKJQaflnYp00I7/qin6OtP7JG+x6uY8t+rp+AMoJEBfeRER5AfxfkxUSbvM
NwTtzmiqKcITI57g0Mdz3cs1QfP40L9qYKQWh1L+aw/t4ibF8nJIRsYas9EVHpLt
jwODz3Kbj4Qmf4KRlqdA2sBKTNa9Uzr7v5V5+VdhOvrbGeDYtaPwIEWNC3o6ugfG
X54mkakdoXbWC2S3OOocLk9mJVi419BqXW04VmqbsKOT6VY4h+rXtf95Tw7KeXPG
rXWNgCal/xYBEACflVH7J489YmTbX94qNglImMMnzSDVFM9YQDdwjDLgCrOA7Kqa
jhrKXLbRV5vDG2GNEtZWCLY4CAIbEyKxkhKXKuxaf7xdnhjKIxaxUqaibatzEJj/
+ibmSmIG+q0b5pJWZYz0y7dupiZcuc+9mp8RPi4Ju53LqZExuEphATPaBap1tJU6
qXpqBrCM0QZGd+N5Vq5K6B9bITIF+l5kqEqeGqiMyOdrOxKVr1jaWVt5gEThzRFB
fLhBCjtMaYBub9pDb6xAJDPiDAIiXWz20+uB9WXWt6ko4z7xN8p/iDjdH5tuEWBg
y1c4yOaaMMfp8nuYJXycCeICdtBw4xvOgyzaPMH+eLqHDN+HkVC8dfdrlJvLaZ/r
ZY+CLrZhaBmfRXeoypZ8IgcFg6hd8C5nrqjpitBnCE6hEHdxhzvZCk683hnEXH+/
azttxcmSYe4qGsbiQZ7/+DiPgh3MEjKNY3M9vF7Pp5RxB4FYyWUbrVMjhgf9n9ay
gb99D667/Avl65As0gz5d4OMWWB1aqPPdpj+ESi/xU3JyWtjW6BBNTBSqq2WHKIG
XoDNe9UHcG2yfYP+kKyTj4wUxN+qAQmbwqBFOgRdyWBj1qYG3yO8RcygVYypM5sD
4nF3d2j8ZQttnmGUjti7ukdU61SIqCOtQ44ODJSUMKV09SwNSL95mIWqOYzhpHxa
1IQx7asMFS0s8kooPK8h+fpbYYN0r5BoqbbaAn2gwv5nMo6XfJBQLifT8RiYJac5
jezDVEiBjAt3vUT5US7dk1gwojqtUMWshTp7RFOZnVJLbqyDePcprAWnKVEsQz0a
OYjAOjG8CFLBhNmP4q5B5+P9L+6hhOQxR1FXd57ESbSbABQy0mgUkJPtFi88iCB8
tYgQunza8KGdpkRdsA5e4XU6nZ0FwMd/xDml3gIX1aYyA5jBixp0jeaUKSdQGv0y
ByxdH1aDPISql3I4e9Mz8k0cuVHKdWO++JUNyP5srVoyYufN2hQZwSPg9HBC3oD5
yOhk0fZNbkmCMI9x94qVlNj5ZaQNvnAIOR6+DCtlwwe6EcaWbuiNWizv76Imw3SR
/Msd7d27a/DZAIzjZRYZv2U9U66pcqPgHCooS6ZvkmKFtyHfamVPWC3AbpNbdqIc
SXRs+xzwCFk1SWGI9gP2+1rDiKN3ujWEjA6zVI3Mgh6VZ42HcEbr3mXncAIFYy/2
VmwqP3AoOQPHQQx4cgDd3VwUtfK2Ce8+se1hTUrWXgEU+BKxmbWumlDG5Lt8m+d0
ip214i9tSCxL7YqAwaNeFi2z1nwnSx2xS+ALUeQDT+jDQkrNIfZNyRDpyQSPE48I
gOUYy/nXXPtl81t7PqpmYBYaOBkGeEOSG2IcmRvTyf5CERRXEqly+xOpXwOsZgd3
Jg6pnMbaoNTDAIo4LIy9A7My+5j1HzbWS86JWvMyAqDrBzQtfhKCiOLDbnXCJbTf
8cMvCFN5KVbse7VhW7D0INWJX90/JqVnYKe7vCYxv5iaECujSWWMEtImgTWLtiNh
gzMToceY6IPZ1agR5ebhcdHQGmnqkeMgYkbXclWkfS6XPjK6xAJwuQLXXMbF9289
J5pHoHf5Gw+K/T6MBTSJRWS5zKh9f1+IP+cn6ZDPNZxmVq3vuaaKIAUMKMZEIlPc
rogHopuzCljTM5ZWFReWmBZVMIDXqyWZ55gAv3/Fsn3yWujIHuhEIL7gI9+Kh+vd
UjFkTAvDFIIB8r9VRGx3iT4yk4K1mxEWkgKbLWq0IYh9QMrsmifneFJGuGcDoZm7
VhKOKYPOVrtYDYSX0z5qkley+V02zSTtmS3FenlWegC0qj/Jo8/wG0wPrtE0BYin
lCZsAe0sErjflA5chsjPeJtbBjyx1h+7n/an6M2Hawzq1anYAzbq8HiPBNw5EBe1
vOnDxkEn10kKdutageT1rBCq6oQdJUuCFcxQTa6SeScR5VZzjqHgJTtdZe3Xz8Yj
SXC81bndDtHG8xo9wYFNM4q5/LdhtVuRah9+d4FJf6zAk4tLkbUfTKVKGPUFOTzZ
XfLK6cFIkI2iG0v7rfsegX/wL7Bh+TOJuDSSRJYu19N0yiyrDawYI0ygvkCyrX73
aTJEfHbPkwS84d5rQ4r0vm5NM99rQPzZ3MscNazE/KVlqk5QUhZsJhQClePj+tCJ
C2VeHbh6A5Qb25hsJdfnDVCcFBN10d+so7GprmcC6U9pTEsA6jxnhR3MCapUQgLU
6j/37CgsgG6dmhnFDnDRZ/zsasleUCbjV8IZWg0G8y9N2bgQG6Bhq70jzBvErTa5
bo4kIG2w+lo2D25jOR+PR7D3T4o5QtkpP/qxm6L5X7iktkBA97wvJzRT2g/lo2XM
kUyFW57N3paHSfZHWiVaf2l/fRUgn3LgFkxdjVRlzY37b0slZ8ClTCCxtvAptvvm
OF2EoL39o8PnKtgDxlRyW/EyvMGWYT9TdbcgeM/+qXoA98718A0CwbwQFUo/ZjAg
RUMyBBQgqlc0POHXgZblak9R9HkECrIj2o1YXC//AsrZG/XR2y4Kbek+9F1It4sM
TD/da0rRDDi8aXdPQYj2IHnmPiRRhNn919DkfrX/B2nALuxjwBTxBQ0HdX1CF+4Y
opkdai5XKGGkqbZAzH1Gg7e0Gz2k3KqMJ42UEFhU16zfnlXWJkCTKpx1DtjRp7O5
WxZjWQfnuQdIdT1VB3nm7SLfJbj6b+yo65eDw68BZPRbLmdRcn5A2YbSGKMQS8E3
6aIHvF+DHpNONWxOChsQZi1s86vpcHidS5KPEUit6l+h25oZFbYST1QUcLMQXKJ7
/lskGSbuYf8aWZYf007oS5EI73DrP8L83HEnRSuuFdVFeFUSXCGZZwMZld9dZPh/
I9R2XpmY0nTLGdlD4bAt2PFHchX1LU2m8oyN+YpZTn3Kuinagg1VeyI3ZfBH/vDi
OPzbWknESDBM7ANsAP8F09c6aUAOnl67fc5iHK7rn+oCdbNbTFHOFjdMrBaxu+uJ
lzNpFsHqeZNVP3pLA9/MBlc/m4LHvbAeh5sn8Glbblq3r9Wz9g5NYNWaL1r+vKCg
6LrN9Nu2ER6y8kl8IE8wL17ATDQWXDCrkxgSOOOBpypMI98USPTn5g9UaDkgGUiH
S4QOpGWuMeyS5BZRTtoxZdKhSsNYGi/4tDEZlOm8Si0MXWSQqPAxMWiT/hVegY/i
Fa4aj3MV/VhVXY8A0+Uf62P7pY1gZ21JPA8/SJI1jdRewkTdbxXidsachr7/rVTi
mHWzzE/rhT+pWFcgPMQd9n68RoQTQCLCr44QSW2z5JRl4lRSppNHO6rbhFDVF+0p
2hUTx6MF/IRQKEiZjG+R76MJbJvD7U8WAudu+tCh8w21Nq8W6C+yxwvC2GLywhU3
yqJutWNT43dA+3bJ9WIQk8+M2gwZ3bIUYoRmqUfvnlFQWRMCaP3rDMZTnCrs8bWx
YLoDw1ahl+pLccyVbb/VlJCQCh/Tr0BLfqquiXv1R3kA1qVTvxQla7jDKzgBq4IC
5Y68QBHWhssv2vVRYUtnKkmWihA64iZqApY9q6DoRL46TOelmpNioPfUmgwz6cGA
Vtc53OVsPPt9Wew8CCpMwEmMZKzSxgShH30sLD/wfjrLSCfYCm2rS9/+yXSNaW99
7H3DLlAN7C2jz7aaUqcT//6WaUdDhTSwfXpKudypcopjMAgVedgvMY4g99kZaMPq
Tbcx7YPcX5jeAxDJp+DGIsNklV9vNcdNLP7fsnUxRrivGnLLXRnvJDazsfZVF8dD
I0pLdaI7NcOkDO4fN0ZbjEBjEwIfrWDtylNMTp3tne1jX7bSbO9MYe7OPSChEP4D
d9YaC4QR/KEeU6xwnZNhVDpVtH0sjaDCNYXMhuzipefVfhTuSuCpnfsyUDEbi4br
cZPxUgZbJdVw9zqIZ9nFpnD/2/SBg0KxxUIEgaPa54GuqQmVXjjPDj+DhpDyUhf/
5lpoxXUcDjJOyQX3bBOWWqIR8/SPx8p0qCjQ/GT2ZuFirmarjLtLBBO7LyMyIT/J
tzKQSgAHZfQxKxeR0tPZ4/Vif11Vh0J/B/TDA3TpkHr7Gj4QNNIHUKzXmZ4Di+EN
IMoPQpsRGDp4SygzujdvHEvx/Il6nzGWYm1bvOC/0i2T4/GunmPvrTfBCfFgaWyJ
7KMkvdJbq1bY7xVXW6Vf1XzqFLq7weU1q830HUTIg/Imo94+fw7zc0WKPPCUJLJB
6PD2mcEJdqeOi0bGgHL6wOodXjqUHYPf4igeq1b9+xdFkhWcBasTbSmpA4B9i9/b
rZnQoRdFWyjnc4BT5OJ1lPyku6O/6ewIqOtDpOC6BRRP/Avcz+aID3OoZuKZumQb
HzjtgL7/WLhkoNJI3bOlnhuhaJ45FEQ35eu2S3wpUcbOgccQsRkqBTgT+O5KzCAL
OY5qde9r521Nl43gqPxRpcp6uotoi9W+6tFnoDHQYcwjFHRHw8GWXKyCxrqHDx70
5xY/ENJtz5yi+FBC4vVW1zbCC2OIOz59L6liThuuUhPwchwkJhFIPw1467lBUBcv
1BsHNpTb490y514nweEP+NaaZBcnrl6otzdNk7JpLbwuxRHQ7blJZHNI1Mh2GNEm
8tiMnKxDPWa+0yQeMWuQwJPx2P/F4l6j3okLmzv5PJSnhw+d2FpomV0wx3HY2NOQ
neGFVT2yzbufcQeF/WBTb1qjCAQTuKMcHC+4mG0JIz04MBlPxTSYD2qV/8+T0Chz
t2qRcuC1CizTvj2hVPwVf3ZyOvok02LRgy57BRXf5z6T33jlgLuqXQg/S6idP70m
FLixKxx8Hk/rNwKrR9MToPaoh83fAX+9OrkFiAZGzPrU96qKYeKlAqWYmv2i7ezt
dEhgru6jDLU2EV1nchn7ruviw6CtFCo3u3iImDuJOLPPJ/UR8gMbNpYgQMd9ER0k
98JBBmMRCtpGNeFs4zNbcdvFVa6gCckNs1wMq7vXH559Vay+rTsVNzuiHxVs/aEh
eSD0iAcaf2fNN8gHkPJVq3Hrd6P4PzOOy53HA91NMcPk/dqvoYDJT12VIJ0rPXBx
4XQg1zfZ21wiCrNttc5Q+5e5Zw1iaqveAadZFeBrlqTQF2SSUGjvJ0KdqPYUzmez
dN+lE5E/qVdCVMfguMnxf6pKgKNc4as+fURc9ez0ugBcnEi9/spyWqi+/0dF8+T+
5BPsdecQ+XN0CiyUWDgRDD4YfOnfdACbhgV55R3xQcZltXEGEx7L6qz8IhiIUS1+
uf6TXK4DSsFtdO51zLZpL7zjtJZFVm+HyB25d68KgUVHOOTytdWkttDD6mBYah+6
EPpITIMFbOzn74vAuIQy6qaH/UW35wNkTKUlv8PMeyTUjmuJ3SkkwYLuLr4CfmDM
69HPY5WVS+BAqYRgMAHCy/p57VHmVK6tsyaKWW//IBBjXwqkQisg+7Kp0miNN20G
9HEJGYGF1J7lFOPJl05OnSkqGZ3NLgEFmvi/Iw1dI83hsFcPBrJFn3w4bQbTYMN1
1nQYyLGTQubeixxsxAvoitLK628Gtu9oQsLM7yVuNyudqQ5fRInV0WCUjU7oIlZ5
Z4cGyAbNo00CBckrOdyxymAFyKfmLgTQ0sNqiIweMwsmllRAaRw/tV3bb+H9sp+C
gXf/k+1PY2fcUSRmfcoOMnycQ7/tiySJQst711Mw2KC/SD/tRHfbB1ZKbMwgnEyX
FTHqUE5ZSCD2Bpagq+u03SZ+o7iEt3Ns79VRljoVPoX5pOaPps2EzJqOPY97pmt8
dIFEz/qsotcj98vQt1JwjSGI38/0zM0m3ravA7hCNf7wneQeSymwbqVFHWHyqhXT
BtBC6S44uUMq0a85OZlvo0N7WQiYowG75xtWpO9kw13vUukc7p+SZ8DrYy/A5Y0i
WfpSgEzDGPCIsD6BOkNhbpE4XEiZmG1lvhthIdnuX/jsFNaOf+XrlKX8HN3MN3le
mDhJXZ7/M51OrnK33E+bvf/10qSYqQjpqfQ8J2ACBUnNk9LnCfg2XlVaimd4rzPE
DXbNDhC6CponDm3FTxxcykIFYmqt5vRMhgf2RQYbsXh3tvpVGmVu/Pdhse40ZQG8
nt8EZl/H1GP+kKGc1gQq66Hamv06iDSoc4sRzeaB8z1TCCZ6XhPxm+MetXdKhm6y
4+/h7H9e9hiUIGNWoGhoRGRDNhhlmwcEphMFgpWlSpCdBTK9t1fwFiclKXt4v6eV
8H1cU/1+/tbXhcJyHfpiXv9VSXTfBvr4t+8FzUSne4tCizpK+112Ezw2IvVolxQq
B3fr5XywS/Pzu7mTmcmKLCcaTqUDF1DSzkHkBHxytZ+5fbnt2Cl+5MLSci/TECPa
rhlcwp3zsO1pHgvQdslcayf5Y+7ijxlOeOdnhTuA+AcOGn17mV3Z1hoWVkag9yCM
Y/D2jDgbCp0dbhYo07yGywCi1djFjWRsnlA0vKE5cceJACknrltPTcDth5S8U4ll
vdDzn1XafwC9MYMq/XQBruIzKYi3Vm0EvaD5c15ZvnhkzIZpJhC3fANHr2t+fyk3
7vuyCurn652bOfjE5gnOCyBs+Ft5gouB8g3pEJmZaY/tLNPMDSTGX66+R6FlIDyc
bOyWw4hSn3EsxGRJGbyj44fREftbAyVIsuKJ04OSEwhJW9ca2IQDOuiyNHj/VC7z
o7ZZoTIlmRo1UFCF7CNW25PYYMZThN/5YWU95bxy0B1q8VYTGeiMP4IXDPYyfkF8
elIXnugjGh6SPq8/KcODI7Cezm7h6giSGsbZTSmBZ1AMsaPgvciN3fPAbk5FAs/S
x2ceLJsRCysnvVfFixI8A2McnysrAMT3bJM1YuyX2UVqEVZIlnnq6AATFavG/71J
R7hdGjRLgUzsKTxrEaTxa/Hd+1mKbJ/qCIz6SM4FjybhGFo4MsT7+NVZlmnP2I5p
+Zoqv0+z2wSAv2qr8l7I3Ke2cHcF0HqenL8aiTmFxq3gsdwzCOC/Doa33fHda0m0
BmnoJprciEFZcOR/mo9CEfzXh8cXnxdM3F66yAZo4T8O+HDYWudyybcEeFDNddQR
2AsYZFEeIQS2PWcBkIvghMhR1KAaaPTARfJeDbcm94iHlD8QucL/D53ig3bh6uDj
L+72bJzHjWfRQiEt/Kop4uXD6eLAEI6ZGaw2lLSMogtmyB2i2sZbUIPVTn7vHsjc
Savzh/+sK0lppischIZvYVhAcHeRagwKIukFLfducrv+Ankr/xldZ81RibWmXCsX
BEgs1cKUxV1fwLSzd8eW1Vup+SmO6QqYNwtaZK+TKKn7B58a8m259pbTyibia9oh
wY2mceicR8c0apViUl78vlNsCPJ7hiQ9E8u8Ee/nPCoLymZa04qo9HsCQy1qPWjj
jnyS/c8BdIwicpuVPBNMcqniG3Xnka0zT+tD0M9JBEUp6QKSvuZZYP/10LEkr38o
wi8NA7dsFefgg+econXu37coP3wDKZDGtChjsEBVE6eh5PNFovkssj6QEQjZCOIu
joQ9mnBaMyoqm2N2XTrRqfE7LlNP7cLpQ5gMU4B+V+cYeLFuDAegWahYfzYLIc6h
R9Q3Ef7cxr9rdPdyPRL9zW/SILtrPVuZRKGx37GVdgEMbi7jgxn2sTJcFK41cF+N
0m0mmddaV6xyG/UPT8vuhv2JY6L3MsO0/Sjj4vwuOLa+yUeJjK9uWvBFV+HdXsL0
HOjwRzv1lhGvL9xI0zeP7mYckOJEM/AeoDwruyXAxAz8AkyyX5kUvgo6A++QhvsO
J6O1k2Xy/mwvU5zcgSoa4Hu6bfcg/ufi6NVFP78DLUnR1/v1uEZdhCgrNbTAQfWM
zz1n+s4uZG8nrNN8+B5LOA2RgLmKS8JIpHzaE8Ahc+IF/HZYZ6e/3vIQdhfDY8f6
ax1vWrMPWhZJ/l90QZjIoS1aixtpWeB1Y1pIUL3jnS44HDvcaNrsnrm3itg27T1X
7+kZ5lOOOOX6c009tDEypcjXdSJIBJmsDrqJwoTwYyF4axxG7rEQaVe/tgyfQro9
4f1I+c4DQaUGmGpjMDB2UTV5zo6Q8YzhostL4viKiI+qgMvkkA52Q51UyhgRBhTB
Jusf6vn8qPNX6tIHrb7uWWb4PoSReutx05JVhFtQNo/Y7y+UACOxgUtMJ7mKO4QI
yw4HgfZBvfzHJlpHDGsiC6ADlLMVB2UnNvtb4VxwAXKWz/YvWGuBN0tJ3sOFTF9V
xYVrz7Hkc3m5UkY/YoV8BvutRTGncBShzorkQMOnU0vUnyqye79jHCkCH1Fz0tDl
eCs5JanAPnQZU/uezSvQzQoD3/yAWwo27cfyH5P5A/IBHK6eulEj5+xDUq+UKUOI
XNYZt/a5Xo0IbdBCwwdPkzhXDITEsHlDNyMjbayZMpmoUGkisH4jkTPGx1IF1N2B
PV3TmHSLk5pdAqCPZ1CK86IIcH32qza4iVQOoVspclZKA41wtsrteI8+6aQcS/NB
hBV4mgQMcxyl1cV1rpvZg55wkhNZp1lbQa7UUBDNfzvBz1NvQWJhhvSVJiOfwGWe
HaYaxHl8WYIj2Jfk/tEHnUUc4KWXieKgQ3ThWRXLqT4qRBuhm03ozHdQy8NL6Z2V
xruRahoFGmVSqezyWiSjihRFMY37lQy+Okpaz69B5roS1rdB4o9LfHztiRICNip3
0rW0yV6HNHROuTqc2+HtgYyaUJoN09MSgWfAi7dAaRHxQV8a9xYKsEvpzn6jE1op
ljDRER2jc7fnM75R8CO3Kkpr+XqBRVZUfMPvEKGJ9ezvZLSAuWv41sB3spu830Io
JHZS6A5Ju0gRCrX/lFFK41fZ/ZbMBQyfAo9diIbpnPsQ51ubES6h8DSd9Y0Y06eC
jNumhEerWoSZhSc6S7FqVFkE3hudcH5M8NlTum7l+5c3ZTHjltxiB6WiYmgSIkIt
VyX4/Qt9xY+5A2wzSasbplDcK8tduN8hXqTyd2JaOV2sTelzX3C9ilykuj8/Ebt3
+aIgXA+JZliilSxACB5iJ57kCs7d6q7A3QQ90LD71BOKTIavBIDR3MP2Ex2eb3cI
ZmO3wgNTX2eHLZT3uEkr4bFg+UrnR9DfE6fRJPf2dM22PsfcCzPdmelaHApOaU6a
YC4/p/i39NHrFkA2QeM5d2kVMSLkGGMGiB8ZuRdQALwVXiBMM4JNlSzG4z2ce4rc
D5qZ3Ma5I2O3wVnFnI/f3QCfO3DvtR9MaCvUpK2AzKd/GE/RmoaCZRcpXXQEXsRR
2lN0TGg1qXvKz5q3ipiQvZTuDypmjnb0xu5vREl2fFMJ1qd7jXmbyUvlFwE7kkuk
qlBY2QbpyGOaEodzuvC9gk3NJc+H2UdhklA1c8Ds06vBBlkdLOzx0L3dVaJbLwiH
I9PY9YnTF2jInrMdXfRnOmwW2i5MTa3RxNbbyvms/DR9b7voAxQpYM1rl9btOOja
ybxxZY/k8A1Rn4wYxQMtay0cgAcTEiVzuCtl/38yqPMGVd/LK6sdTiy1VITac4gq
dFclp/pXQETBHnh4kecLe8lhj7swAIepVM/cE3sxXol8Ma7bCBArW+7CVfvSifpn
4y7KshT+S62SsT8H1EJlgUb7/fUv4wIRU0nCUkduWnvEoF05BNTe0TfC8aDW8fQN
0PEgcbXlVpfsmZ9hLjbxPwVSE93hainPxAf9KqLBod90l26zDDw6JCS5sGOrJ+87
aGdAKN6NFRq/3NCPd3H4JQK7TNCJOWIXFh2zAr5soshr4kZ0gOKfPp6BncHw9HEg
GvtUkBWxfgXZZY+9pJtS2v05GQ2GIT9TutOyuC7NicvrmnLGSpuu9qX/u7pEVJUr
AdHrxKk7ty7NiRjcGoJUe92Evz0IYMNBsZ7T6Vo9NtWFIZHH2dJdwEQO4bmlqEBX
GffO393F5LIBflhRLVb8yREOMeWcN4nMwO6Bb55vshAqkunfxaX6/o5b/2IwEBhf
CHuM7IypnoNKmQWWJkkCtn1deTq9EKRKlStboNQ2Y6HVrWS5Geo1/drg9iWQPzcC
zRA7po6dFFmxV+mNPG6crm5zY4pfpZyskODwrHqr8nbLazC4tm9YAFoi95/uFUK5
NNDykI1L66iVPR/kczASQmqx8ayMV7ALp858PmMvJ+y5BJ7u9uONVtWp3fWXrE21
qvt7LReCNlkN4qYO+lC4OBv9FlJuZJ3w2sKn+7XDeaHb60xZP6o2B26aGnclxSyw
qCuvhPk+sn1SOqv7KAxjaQqS8Sr8nNounM4pocbn1NRkCM9pEvkhnX1Yh37cYY4v
rEe6RVLTOSrgplCXnySa9hrQbOjM3xkn5ocRzZnVu57/ezxLZVgeEoWBBSsnDExA
EiC1G98u11QTpRbVQ9ah6+1q5AYogQgNoHbLOpn7Nj/3tnJNfHy0RNmdxMKBYd9T
TwGxwLYsoMlgN864Ei8UjN1oaq8fbmLbptzq5t68PkpQxFQGpWC1XFCJzUXr9Lm6
9Yd7zW+6z2DhFNbNl/HaQ2QJMS1owWUxJVFnLYwmDaAdrtS6LIXxIjq+/1ZJ8s7O
4Px18sB4wuRWMDqWz5qwxsUq9Br8fj2ffBJ6oF6LgKx3gr2lhS8/HYRGKmn5R5b5
fopak9CfBd7SeuMfpfzpptR0KY1Wxvy2fe0Bg67DSAI92+9SKwZFTE1YOP4/YysF
waJunQQkJ8f2r1JI/FnQH66jEkXqyoUHYRiI/88nZpFR77HYpjp5MDP0EO5jvzBl
ECNNvrfD8mJsHk7f5Ig1ffevIK7NQcLvgC9WX+uoLOG8cLg0VP7mbjLfxhBF+pHa
NpW+sUHNv3+M9836Ku22SihU0kOyLGBDK9mvg4FPSqlE8Br7hsrgx98KKOAbI3Er
hmUkcvw/lCdMB7kiRr+yCdP3tLiuMyasYdPxL8rx/xYOKCCCN4AQvzYkyHeWVONt
BuWhKsO1cNc3jHXP6o54FKz4fX4xqQ89GeuG9172EqZaixPWP8T1Mvydz+DB4Ljr
i0AC4PPAyFTm+s2V83MC2Xqv/fD0g3PDVvSpIvS/aJvepYGaRE3JhnjrDm37XGCD
9j18IGuzqdA9QbWO3nRs261V1fHiUpVmi9AcLyyCOeUCXt34oj798V5u9YQE7a2v
t7bIWD4CNMeZacMZbLtGzhAQmiPgx7+yr7IuK1op4l4jPJq9s1dp7i2ZIjC9QXEY
bFETZZcE8K7C6fuJp0YC+tqHIbRLPv5LQL6WwyORf27Dwf1gXPm0UNWs5LrbRlvU
1ziHbm1Lcyjr/cFW576Jv4sFlk+duMDviistgKAW4U2+RXfMt2/Tk+gBWx5PpwNe
TKFLKDkByHwHtonn9T2ol+4GlBUJlB8d/Jd8WFPXHJHGdwpz4sosLoRirUPE1sUi
SWftm80lbFioFQ+Ps3h0HB/0DRuaTHoryXK/scUSLm97KgjYCSq+L4MVl7sJaOkn
K6CD1uAoY6I3mAusmFH7yam/0ldxg1O3zwSJkxSlgWFHNmNAA5a+mI/MzcvAl+0a
HCSdNuxfGEXyu/YUtOq4Fmeeetman6yWmsHYc0rUC1rNXvnV/P3NCWYtq8rXQR6+
1ZMsYl+/8chYgi2ytwNM/cybM3WLTWfKhf+5r5yvVcWx2bg2gXgoS1MTGRKL5IeF
B1CXFLBLm8dXbBouXFysvtRY+kP5s8BDsBUP8FKOki5XW/lkcdqBMw0y2vAHrNX0
L+vk/bDQIivVEZ1iZuXH1UmS0Qv3qamW9/kfKkOVMEYL8Oj4a/NLdVb7Gy+da6Du
XFU71FomsBPbd2301pkL28/ebgfbEiQS/yC4Uv30CuBUmu9DhRPDzXwM/lk1xhoi
It49O1/udvgl85+NnHvQjrd4uUz/RW2NYu4gfi/HLkmH/atDL1uGaH6lqA1/iMIK
W68WKLdc53XCmNn717QQxQh0s+eA7I3Ghg9O3ymIz5KuGNxz+8ytcUd3GuTtIU1l
xfRjM2PaPi+pRs2ejJcSNOyQ5T0md3kBNCRn0KgFVpHI9kRZN2WpW9GkT42UCj0n
poH9mav+u0Upfcjt+Oc1sJoLKluPibHYAiLP839uSbo1CvfEsoeRrNg7aKGIj8tX
TuoYdKi+FqaDQWZ+mnHCJJC9XLyDQ11zkJ6hM6UeGX9CsAPSuJ9koTH5/ss0SZyj
vhFg3yko9ZQDXbm5UhB2cbDkgjAS+znoHGhm8wlA6cTLTNswHg5cqRxpOJg5rh4d
C4qTl/eaBVuUJP99G287ViilKP/uj2mYk39b6AHS6FsBcX/CYrBjxEYxqekuX6kd
nf4zf5KtQ8+DALlP6lCCeQ2H1ydXLvwhiHpNvCKhXvRZUdONGchc1CaGm8u8f0GX
Sg7z3DYF++AW7ywWolGRiNS1ruWCoka4V9B9pHxjNjkBD2jwqoiGKl6JX+1XdAx9
AZoUs8wC6k5pNwaI1mj38RjLXjKeDnuzy2oIjsovA7zdErPu94L7hmpNXFr9fOG+
9kIq/S/oFpw9Vizz6M06Zin6PG/QHHa5cZxA4snvdw0c61vVg/mOYJBxPyw4EISF
ZPwOaKHcbLanbQ3357MhmC3l0x3hzic6rleiBMOdxR0h1qJP/DEhZrrriq7S4sSO
TTS85CjCDAcl+VSnWaSIQ/Y7lgzxCqXcfCiKcYFcbRSiJnBDMe8CEKVI/pikUXB+
/gHPTiD9+xYyiQAT6o7QtNy8xNn37lMvPfZ4RfvWt0KoCUHaaeS1OuBurw1YIHTF
U7wH1mIO1bwFMyoz1nh+kfCVSd8xM93PY1z2NBSUldfS/9QlzvZrfbucOMRgs5mv
oq+4KoQ3RKbLqLuHt7OAoPUSFVedg35muFCVrVMZJwWJQoUE3fOVOaxDyzLZ7DU7
O8Q2lUP6rSiElzptjWC5EyrOoHEAL1QGn5+04SuJkSvq87dzfxdvVXraIgj72aj/
+1VnhFQjFjWm9nxHB2CFrb7gQIPueIFYTSuNwVT6pRdwCJ3d2l2TCjepm9ZEEN5K
wvjyjxO0Q/9Aa1UX47wesx4fcvaXhzbHl5jquUv8C+yx7yazL4MSFlSHLRTeaiFO
PRtNx6i4MH18EiLakqzRsAgmS8IB0y9US+7hpGVfSIsaJbTsK/NMYVc8VLwly6V0
mTuji+zLz/Qx81XQR9cebP1RGTGHOgdY/dL4Xp8wEOljNCREkf0sJZHEgnBwZO9H
A7lfq+Uo7ai4tZ3UEfD7NHGIP+To2qKiJLzJCIwxkI8l0NAOcco2FNxXC4jcHtYs
sWfPCpwCgp0s+bz+0dcVH5jsBS60oPQMM8Fm03MfZbNL9+jBn8mHUJp6kboeB2d2
nWkmDMim8Pm4hU2lfvCiqYrj7TxzMARNwFykNntZapNqxgLEtt26ZIW4ItsS3eVo
caW+E7b7WsuLDryv4a1lLk89WU7MR7hjy7dLBwt+mXn7bY2I43L3nIwHiQRiDCnj
iLPAlzPnvECEp3S3JpVGFF9nt5fY0YL7K+N4rrtwXoFra5dBsXnNP6XqYIbxvK2W
RJM0sH/cNqonlmIAyEbJvovgfFemRdFeBHlRI8My8uxv0OYb5Q081TLrrhVJ6ovt
u5kEPoqpXMl2msML4DMWB+cb9gR/lAD/5KGM+OIXsnovEKqBUM7Cx/OspzFggRfP
FEzOEB40ugzfUGgZmG7MqlxpMjIOX3FDbpdlP1AIvOingV8/fBQKZuaULnV0kj+F
/eJvEpBoaOy/D+JbSdSypVV5fWxy7ex0PZshWgfNUzROC5b8HMBCeIBPpHr7FkDQ
xXp4RVUc8YtTKD36GSYZ2ZqemNV3Ux2MlzAJVHTYqys3zBOm/PqGcVlJWQ2e/YSE
HhUTSwfCkQEtkN8K35U0KR6qD5LjmuzDHXQX77F711IhkdyaB+6ykFaSekeJI/f5
mo2AWulZK1Y92FFMEHJRDoFrzRi9Av1a57+59za9Ru37OjmlIf1As2fZO7WZqDSv
vGdgQdArlS8D5oyKB5EmKovsZZMTGl3WkweZhcU8q8fd+L1NFCLIrXgaUNVcL3QV
gbm5iQoE+ww0aaUN13HF8VsjI3/N57EmxsTBKqDSfqznlJmqOWJ9uzoB2nVM98dM
2CI2tZJhBKgKH8zfkq/f0bCZ6g7+HpeEOpL8MGu0/8SPIZ72C8nG9TatEoQSAQYw
LM8/q4wUtsBJhfrh+TRf7K+t78IAHzQEA66GMtZu2IgoOigQb9V8fvJm029cRYH4
Jrcq4c8owcTa0VDRFMErrq/c683ohCUB89Vcti0i+PUlcZ6jblpl2bKxF92vuGMD
IoUt2EWkgnLyNuChGH794xJCCwB73ddOCopmKy0iHwxAnPDGlFXhfDKLkGPBD3fV
9nNGlUaaXSlKY81tszvb8QF5uCQn1BFsYj4rUnZguopUVydmKogDzf73DHpyY54f
fbqOXKOkw8y606YL4q6JaKpFHXVytk2X4vBpyo/T4lf0YE+YQglqTE7k2Baxgq13
3m+YSwh7FMSMbUttsGhH77sTwt4bk+4Zx9Y871HnmdKesehiYVBmMwgbcmAkDX3N
SP19810j4ir1In1Nbq677SFjLmEkGo52zPh8rsJjxi7CqBF4TshJVQzRAsn0GrS5
wzcdZtA29COnZ0ZGICDBJhVLM2c+sC1/HDWD5RCSHqlJIncaTO0qP/uxB2STlJE5
k+08O52va0/KFSEIW+W0pNp9/LMgZStRl4EGaCLJkn+9c8XHkfbgyphxpaEpDTW7
8iwvOyNE9ug+mOeM0BXoKhxZF5GjEY/AWx7TtrgO8TxsrhYwFbXBFEwsmulAzAIK
PGEXwX72yEWXyvyweQRlkl4lMvSVs8sl8LJsAprw7AwJZVqXlc5TUFctP862XDY/
0MKERXY0IeTNnmsI9WHCP55e6eg+WXIwCVWhEigskZY2RmhtdQ4zG/lUMa4I1jYP
pkr+hpZMpqnwwHDxHsND4L+BXZanE3Coreyqv2OiKiaCM1beWaSdCsUKBquFXTht
Jd3WDYbbYyL/DLNGhkL8Ry79pTotbty3g6cL3So2JSSlZd9EEx3mBvPiCzkowWnw
fKSBVj7CzkR/aq64PAuWA8URBShW4zc2ioD4UOV+RcApWERvNINk26DQNyZfDM/6
soo2cAvtUCwP3DLl95sckKzy6gbGQZBxPwtDghMYLCkeTMqDEy89cO1IMB0ihvKI
8I1Da1av7QKiHfJsxblenSdUpk60ny9jgJ6lU8FYWCMJHuH+kF1+l/M4kXtis2tn
mMllsKeQhoH8yZlLqBuLz4ab+YNUB0F8sPgG84BtueP+HDpOjHWTsi0wpp5aEcQg
TvhG5JmUBWwBZ49FfFkF3ta96rvWAfhjowoVVZac3nV+nja4rS/WNpded3U8OxqE
TkySNhxbhij0RlXNSk61EtMJiCNxM1pUomFzl53hvbVqS1hvCcbE4G50FjDJKIEO
rsrmqeyOrFalrEitRVD4Ykxu+6At/+braTmQfXR7nrRE9SUCsNVLk6dql+qSENB1
o+QrFP40pP3jd19iO5WHdBnb8jfc6Fp1cJGVr4BrgTZdAHiz73opbmvvd8QP/G+k
nAx/sMZDJkZnpNtel/+qecmR8FVHfvTPaOe6oE0aRCKkrnFKLHQxlZT/73AQsBSS
Hfdlfx0oCMUzN5m2FLh84NmnUtZHXYg6IeHAjPSF1tO8VOydyo0Ws4NQIxqAvMK9
Zj+ChSbng41TMWXu6corIvx4haUH/oHGuRg4h3h6Mb6blEEVyZdyMtXZtO6GPII+
seTb5DiiQIhIUQJv+t/Can6qgEXlHi0jCAZ72cQxfPRLF/A79258KAvOaG/Sk5ZH
DobbV8urVoMOhEPaLJ+DiM7Q+eyyhLL6heyHlZL4PMzTgdpAL931RLsqPLCp3Yzi
IAxx1DvN6IBf0f0fpcnfYwYQwOkOkVXrD71AmS9muUDxumJ+bEaAQSad2t+BqaS0
ea+dBiqC8K3nU369e9QwPhWgoTJ4AcA/KGf88HV9UR4Kebx7PB/O7cIzVZNpUprn
0fQNk2+5MzUR6BdLfN7WjXnhGTWFkgZWxkPNQ7ZIUhruZUJFZKSXBs+Gn5GFttGD
E9UoDjTGciBqVoLNMt0++FG8OibSIuQPF2Oxo4MzF0pTEhLp21zOXAG+rPtlE4bT
A884G0TrnY5T7fMqmUo5q8sTlAByPr8mXptoDMhyte76KKRjwesnuhWCmNvRPhjk
bgvmaDd/IfpCl9GDsobXAUwZUxCh0YF3JeZpSf8hLyLF6bhmalBzGXJX5auaV42J
bHhYz9DQMUeKjPI4E1Ry7Eu2wXvIhDx5H1noTrysLjM08yzvI8XSsIT31xPEdLwI
ikV+dopPoMEai6SE11oVt8DW40+YeZNTuXxpTtKkVgEnFlsCQt3/fnDOl4J212ro
9nHqh6GxnCkWURyGNn0ARuA4+fH/6ut3NxiS0m6JFf5wUglaYWX3x4v1vG2PqD1r
9DszP1p0EoQS3n4bPY5AR4pfTySXS60HUcU+hIFR7Flxp4sTSdxEDYDfEJDjG240
Powtu9cnpIZkX17fyqgoYMWzB5VI0s2l8XSAxHCBY8xbSwabAD/l2AW0DkmAP59T
rYTUG1TCdVmsvwcPQn2ni6LNCCyz9RcjvmJBt+jIfACSGnmwSF7iYOapru92D6Ad
pE+q2HPQekuZOD4Gq9PJ/+q3hSeRretlI7Dgb56lY/uVnQAsEQF3oXe6m7R8dlXh
6kJJOn+kJCRLPAaw8YkaDRD8O7T1ehrNfctNRfznqm0LtlLMJrO/V+WpABWA4z64
WRpaOuIBz68NjWUimvFC+BDMNWZtmeAsOI3pZdLwQQNUz3c5u43F5vyx/nyAzOUw
9fSA8x1Y/nwu9nMovnM6EiSw3GdB7QeDFkTnuKdS//MZ30aWd7qjFcr+Usssenez
9oBdD8km9dODKhQkyHYt9QW6c67uN6CEHPtdsAewUUzEaP07DXd2MeUesk99+PvX
tJ4cSvth0JRlMX+n5x+WUSSfH6ofJEb2C53CJUmvZ6F/yNPgcqj1g51NHM/yje2t
AXZ3PKZfkGl2E112HEcnP051kwfOci32HpPyrfcHkYol+/09DrqasU9ZUC1shk2m
eP9M60RVGlOl0wt1hsZuPga3eNN41gNcefH/WvIke2ebn565QtJYJaq1OHkOjKvO
jm1hI/zV5rgqn9etfkTmhRboZWP1snIV7WDAsrPA6zsHveopFDNUitEygU4qzUA5
1GPqq+NrMC2jliqv+9pxUw+bBXd89s+yRiZJIo1e3Vt5KJIS1Q8g34IVG9wqYWcJ
ocuQ3yvgetSH+amOTKVAxnbPwqRTaBvGyXvJBwI9x8y5uGhY4mk3D4tBe+gYVMY2
hZvOh1tsy6ZibIBp0pP6XLaGT8uDqOb57XxcWCvOdkuamFwcWBue3i9Z0Eu9dZRe
UpNsszANvsrrj4sRCzyPUcsVojRs35S3wpki6XTOVJP23zm4LBAv9M4oMFHKdUrL
N7J5ief2GyGDsiigWteT9mG51yOVF3QDk+XHIbwvCVOl3dg58cGQ+Yd55E8QKZ1j
fzL+h3jguFXnIdcBrtG+mxj5FwAHgTjfRx/qQTg9q9gRM9D9b1fSxdC0nKb4YcXZ
ofCE0UgEooCYACJ2khJC+GpwOz9s4dZAMEgZ2oZ96mApCDaOBfV/C1kic4L94goR
pskBXrd6MRaLzrJ+ctCKdfQbvP8+Ppvz3LSth/T+oeCDw/aHpphS1KhmoBNwQxkt
GLA6BM9c7dOyMGAKWYWfpN9wavwZdRxd7e9KZtPctzrciXiD1aXu3M+wPX4wWa0v
U6Jl/vONpaO0H4BoK3dzTrGrPsiREkDlNxVna4tW0jRKakPC2gDstFdG2IY3fVRQ
g4XNn8ujBI5F7bXjDfsW0nMNsmD7vXVU7wCMZ4VtmVJGMgJMk2ZVTWSQ0tKy1NtR
PoIqdDeQQwJKu6xMEwy6HjyKrpPHD0r6BQaCSwBT4a0A/C7xZDv+05qJFFJ2F71E
hKUwzCEmhmGrZiqm6Mv3aCvvIfwKkHCHqV7WMBMBy2BUs+6QhwLMNn4ocqbWT4vJ
v6UMf+woXRUGL0luu/lmZelZHf7/KlRfFIrkFzwB+hktfPK/K575+BJvWHaN6WTu
aJfAdxNQgTwqLKpEVFrGU9bnZ9V1MxpJqt9uy0wwGj/szVzInfWlYe1Qvs9pxAuV
+yU8j4NgqJJ0I1s376etWDxk/S9XDMkWMGsoz/LwJv1a/uA+Bcew1il9BqfFEj4P
uIfVrHefKzgC3XBfgbIGBNgB4tKYcV84cx21iqo5EBXToO/cy7GPqYDQoQJdhwMM
N4Wi/ZhKug8KAz9Pk6mi9DjZpSaaspKi/3o+BQa5j/hpMYgHHo+eHUoaXYqAFPFf
3F6MPYJw49ooFgVVHMtBwSRv2yifHc5D9zXY7SaP/hTNqIN+9Be6RjGkGULZn8Hx
JvrS6Fxv+YnntRKAaWgJuvF12+gO2A6LeR0o31aKfDfJeAKCs4aPl3hbNfvSXLPS
SZrd3VeVNaBBd7rcXcTgFtHPNpLmo6NueCG+G1um8NhN3h2GiHDlNgBvtjlF65bS
rNF5lxG2Ou5ZkhK3LSLe4XGDNMFiTTbSGPF0l6DdloROGblTLGACIKpS2IrDW4L1
lUhDKYGkUQkl84VkXKrTwHierE9BLq9kDd0b6RtwZufyCL1Oypt0h9/DhgdDAKdC
xDzS5YphMip0yaBxPgn9FIntzYZ2NYmq5uM4heKkrKGe2qan813Gu6u9oVP0Y/mp
jKUXqrLqoriwxxUhuCmUjryCoxd4LJHA136CDA8s8Q9xcbhHlIOSPRNt72t1/nMg
+zDhNwbuAdDdPrlMihGiIzmC9SpMyw0PDzrnJ/5y8KC/d6NMjHummzNm/Q0GYglX
UMAVuTL2jihjxEPxT0dWv191VgAewY6nkGVHKA4n6/OKG4E6aloMHj6bs3JeHDB7
euhaM/2SXRHK98gcnOCsaCOqnM4/hlauG9bLnbuX+hBEdZz5bBMZURqdgqZywpg/
Q6m74nQ40ltMjGAd+16F4YLsE6qTjzTG1IabD1mWe89c85TSvYZdqu9nuYjW8c+N
hN8vOl2YxzalP/m6PvOhrmGHSeuvTnZnH2GN+NEiCfkcCPQzfXtebqhZMM14BpUz
A/BHHFbXM73YSbfZyLvYcL2pmhEFouIdRf88SuVy+WEOoQ3T2xKcei4GH+4lAro0
w//4kuvPfNnCWqKlWC8dEzGgS8fgnOlCCK06/H2m6dJ4nAi3tAUXtvzVvbn3djHx
s4BXTCKiZpsssJeokhB/fk9nxyxaO5vd/XFQwYMNEKFQvuigdRA5/axFAMATnzhz
5FXEmXzeQXkfWLXPkMEkPZrm7YH9sCI/bjRjb6rIRhHTdzqE5+r+vyMISs9pkGYQ
Nl51AJ6oCiPCljn3ZKiIhQWj8zvghYmkR46CRx0t9naq98LlRVSzvMvEHOMJSCOK
IjI4I+BgPEIncu7E38zDRJuUQ1b1OWx+Ksleo1ecu6A5uGBEfnUijnmiaVCYZ7Q0
n09d22mU2pxhxWIwBRSrFqUt0/VzXTushkKQkrSWs/xXT9GbhEhgJ9U+rbgcMrlf
U/SstVhuSBNG+4OTRDqAGhtQ1ZWQGvtk0YqAsdKCDZ4CW0sidda0Y28sFzniTZRR
xphRp6LNnZR1ezB5SJvdyQROw1lohZMuBIq0nXQzKKtYAilapZTYx2nliXk5YvGg
bO7mUbgG7rh3gKOEgTUOKSiLeESHYg1D/uSP38YBvUhFOwDA9p4plWLhsYkoVw2L
HITF79sEQhfHCmhQHedCTqwOy8W8pJeN+Z3+/KwKH2J+v57o9k00Dkgc2QQiK0H5
xlkMDNctLMSPMWip2Br4r5Lrr6efakZPG/F5EQ9gtpOLUK87dn8y2dJ4rDocdZbg
HLGJZMrWF2YzBMKWtcRlFtxcG0RZPfjWzNREpGWrfUFYlA+LbE1+6YEnTzcq45i7
6Z28JKhoVSzs47bTrRjxwq5AWhCWb3sMKO6BcN7K1IxUnaHdwKw+ewaR64eYCeuo
c2l55JdX1d153BPe/hqwPGHjshigVDf9jnidsPvT8fUzz4GxMlQ9J3q/lch3FIA9
gVhNsZWK9vcUDH0P5zj/N8qOiNG+CNgQ8ORZkdIP4gO77DreoHuH2iMZe2h+fSmL
/Prq6zZobhUczTpcm0GIsE+9ly36rZx205VRvKtjJCFBIu76U88CKyx488GCovJT
jkJpGvkTLt/xyVxsadEGhyycf6HZUvu6UHacbtTUnW4RVV4F6PzaAChEWWlM9aXE
KDLvYpRR7T8rpOwTooUSKWbN/7ih56cGVTbxRRoCD6Qc3xZSFo+cPKBpRTqoYTWe
wo4QuvuQC3aaYUmA1QHRccBFkeOOoGWKrKMvgSwBNNbkiVbpaNpOkp8JkHcaIvwt
vjmaHnHBPxcXGebS1LlEzGgWMD7FNwGr+izjdi+V5aJ0UhvdFZw/+Tn1wF4fkE0l
/1Ja0WOBo71SZ0VriQgLtTK03dgs1ZiHITM3qbZaroyFMnjq/53PX0GFaeyMLbI6
5DXPQ+ORNcIWXePH09VYJdNv06/oT79xYYNtkkMH/3JjobUn1p6hxkb1OBnT2tB0
Go4tN0BlBpXEkDxQ4UccKRtweg1r3eHzGKL+7Nl2+01tV0c7VG7QrWbj5wh8VA98
KeAqdraJH8wWw6VlLVDKJjuqdqAfumIVdj3o7Eu8MOTvz3qRH1LuMXDOShOclqz4
PmyWjsq1BayXGRbqWCfQX9viiJEhV2t6kVn2eLazyJrZhZRVtndVFiEakc2WtQ+F
QiK+zJNaa4b/WXcM3O/wHajA2TNgezPf2ADiw7GlBIpC6sCsnWQn9Pc80/9SDvwX
rPV35Cg5yR6SJG47fVrXjHqqf3mu27siJBj0JKMtc5jgVIatC78xEeIUy0ejuT8X
qOcNvmHfLkE1Nyp0U92O/U8Wms0vP5l/qEaoUGh+uPc2nlEiM66h2WgW1mSy7E0p
X+GCI/WlwOTF4XFzzZ1uPNW2zH/rNjVwX9BS2fVWlArqgWboONGlUcYZ3BJPeHuT
e1oa8sBC3+tIqqiRhj0q2Z97xgTRRcKT8HW9aD0b+9K/AMnyrUotcQAm0tkfsr8J
91m7Tclj/xXQzHXZRaWlnKQu+VNk/Sk4VpDIXCRsvhTVPyqF30XzwAEHm3bDZAEK
0NjPRiQRH642kLsIn1OK8gJrRFBosWdUTXATqe9l+1b5IJ2hDhet6P8vF7TvwH/n
jZC3E4QCclDxoENY+Fp0zj1Iq6TWyDU2TpSueZFqdANEpfWFpkAyCp4htU/z1DSj
BhAOU6YWKcXCrQCH8ooI1EO1cR9BDapATeH8tbLBNXv3uWFSap053Odsf96nYiws
KBEMwEWi/vwYzss95Egn6987Qz6JGa2sX1SLTFE7J3LO65NHZRQ4VjKSRbH4QVj1
vM1jkKDomo+AX64cYwK9Y5DB/RMSlZQX5DVln6tXeaWdXFXgtwKC2s85uWHRGyij
PicGohQufNuimDLARlhm08TYvsnttGxq+jalNxTCXOr+m14SO080ZGQM0GwSW5WK
IzOKnEbyAjcX7yVHHxOykDcbUCPEd4R77lNroTOvFKe178QImfKBzEDjvBKvZLtP
LrtWJUoEDTNmxQFzheWhPjYkQvuHmvHpBM2SdVq6ki95gDaAMZ9lErOm2tX2dS8m
69rmc0pP4Uewf3wWqohj91sxQ9imC35yjVClko0C1eWxcQllUbuFX7afX4ohOtKB
tNAHIcb23Jc6rwU0Kpzx56b5dKKs6C+Bc2Xb2+oLRAJq20qLSaeJWNDzHwvxoWN3
PGk98JxZuxLZzeqtMyRYYPq2iHnaaqTHc1B7UGx4cZsgQjMPNTo7GDOh3uZ0vPhr
XXevcY06wekiz1nxiFzsGPi2hxHy7qRVIhD98uih9k9Hgb0GooEWu+4vCtLXOxvb
NCiVxw7Ul4fWE8mrmjZT3hwL0aMRxhWEdV4EzEkGsu1PxNDRG5khpu03zRkCLRpO
fEu7TtE0Gos+aBYvrLzeji7ke8s/UV9OxBLqoooYge4zzSztn55MD17QeuUgA01S
cI2n9Tqwmo82XJ3tEz2bJ0xy08m4kb3jJ/uQE9TpT49DE5rkID8gIl48ovwOSInU
1Xmrsz51eAvPDxOiCjOQotimrF3Im3LJGmTdd2uaSJv+7xzezg61tbLgLQdVxaOR
3IewQWWvrr73o4KgVDd30cEBqRRZVJ2g9uFek/owAnb7AzK6NjvUSbuh0VRDlHth
Tf9nOdrBFc6YmUW25FzHlQ7I6vARssbAyxVGLBLt4MiD+XqEb35pqMCaw64NZ831
/2fGZUsK3L4GjoIYziLIBzsvT375HjXRcrCDGL591Wk7dWG5cVOH1XyCDtf7qx2t
6kqx5ASXEpn5U2lvyJujuAYj8sOwzLHsntj6u8Q9BOnEu8LTX1bZwXJdCZMS+ADg
ZWKg8Lvr3pz9QV5zRmZ3onsOunJpR5s4BBxkUoyKDhs8zD4Xtg7V1uyInPDyGpVq
r8KKaNwzumGyhJvGrft6qDgeFd28yZP06LSKo1Opqn0xNoblLmjnjbHM8ygdF8mE
VNds6eAjsF0++DS3kKUYFq4ZPKVJeT3PG/pwuqnU5A4qDpZmWyGodRLx3sBhoWJM
uaMCpM6qax3tq4XvNjjG87WIKx1pdnBOONKi7pvW/2Iy8bcRYoyU9reh02iHuI9s
FUxwEHsGEvjt8TYB6389/SFZO9ZE7HdYCn6gsmwI2QXPK8dx/35AgMtnEtp1gVxg
BFC8HYabqqcqjdO0esfcTJWioap1ohVc9B/t99MjXJoRTMBzeRe5JQfbzaNCV0kj
10I9ddPwnE373m70TFz23LbYjKgvK/ZXiGL7dXRMcbJc7DTuxjrAuwgNNeppdZ7U
8rFXlNG3l2MQt/+VEje6zpqbICO2Jpf9apTNQcMwtrlycKQRuM8Lo3qBsGgW7L8P
kXB8kA/ZDfaXbV7HqJwTGTVjv/r7oxyV10oOsvjXElL7bNfN9Wh/O3tFCUwuug+7
WmnWgzfkYwZ1oHNHn1raydjIkVoOago46Jk3TcuV640VFi881d4OsGXkq3hIap34
WaS8cmtOMUCaq1aPcM2hsOkHdHrnlhY/XiogS4jrSqm8YzUZZw0VLaZphm3zWQIG
VR+L4LJiWPAC+HblKZFlwcZFma1BrBmatMKwDSLg8CGoDrHvlq2vmpO8I4z+LeVO
miTZPjJ0rZ1LtYuJJnTIzFdWoKX7PA8Uyd0y5SWpaFXzPpMStJugDMrqqq051Pow
ZYu8rVJH0++W3F7bFCnJDaFJjDBv72WDCSJtpCLdrR0FrFaVoyFiVqiMQCNbj5L5
YeRq/bgOkhEo9boXrAvb2BUHFMBGMiX2c9cYcDcW9LVDkRCNIqttwY7G/pxIWHmr
COsAY72IIstTpgOUDgoBbkXy4sS+R1NkG2Uf/78fidNse9vYZjVwgKOkpONZRFMq
tS0ejRsTmD2bcMJJcoZv37qKv0IQ3a84IuS5qpu9/8GORjTYIBcOYgvW1PIZhwiW
HGYnWKzJhECAUqgho+QAn8OuOLZ9FMjdpPKE8QPVkgcG98P1v1lbo+30/9fNVej9
8AjHcZrbm0297/s13dyLA41C3WIPa1QUMGKr0shDzoVl3PVQ0HmtORSkh7iOg5IV
6nuvFLS0qa8EC8kvqvk88wL8cUTKlGf6Nqs48ZC5rtOv4vGtfQhHh8MBjaIR9oCa
d/LkyCiUvmP3nEZDbSryoG3D7f2gnKHwLTKK1uubqgIevcTf+r/m11SdDH+ES39P
8W7Hj3IBZPQ2ULobbhjVBCJ+C/M94YD94BMJTtmEUGM+MDhYWpFmDAcWR3oIjlxA
yfq68LWNIlxVU0bAwqpPeISAcUeJj8Rsc/tlRs7sZhdPUOmMdUsItboCp321Pekp
5JrD82QMxLmDJ2/X6rHhCgoGWwPL7nXZihvbOU5hkm1L7xU7cc6MYGlEB+sg/B2z
bTLBQaN9NPQLiAnoZ/kDu8jYVI4uxxyVAKEKrqr6yeZcGXZ040yua12mTmOQ4BiW
Lx9p5vCwSTlJJTuqk8cZLuSCHB1FIsFx3m+5ANaNxw5veQK6/H7X5lGi8xXLhgCs
Ez8fOYZoIA7e3q2quBl4yEiELWF/WBR//912eQyPWyyaeAXJZUZ7S4/zh3mmQvgt
wsGuaiUJ25zo/czYB/akSfgrh5+R+sS/YpQvNogPJnJkjkaptJr91dQ2dk7xdqtZ
9YbVivOF16bID26WNPVDwrL560CrNUo0c8HmYVTDGZkXAADcExqVoQqxidrXdTKw
xnLZmSJbYtUNECPYSLIhLIz3BVYkce88qatYMvGm/pZGTT1lckQLlUme9S/3vnNf
uBhr+ZrsARjxBmkPAAllW7oxPIjjsY3E1I2fnqyhIe7dJ1wtastEAxy96CAVSkhB
5mhY+cdhQBMMgo69+RgOhBWzViOdPwQsmgvOoCsH2rkKp/L4egPBlDLqhtcVQ6TD
udls5jWYbPKz6ts++yLVOkVlf17xRySFbnUO1jq3sIrOmFT0w52W3oaDPhph4SYd
/pL85k2xo1jYZKFBw1OuQP/9k0grl75sbbw4rEhEPp2VCdpO4SC+2oyaxAbfC6IC
34dlwayPQvqeGN2rGjqtA9o4JrCQz+wGEeedonIYSmsTeMePKUPeo84lwyrNGjG6
Cw722dEd69W3s34rdzbnaOjREXb8GV7n/KMTCRmnLhhNQUcOW+Z1pkUao+LZXvCr
9QtFxEYNpqsIvHaacOqAZkMlzWCJl0IJB3I0z08ANw6Xjmqy3o/euQBgEM7JSPrk
YeafLHfbRhLVXDMsxuhyak/DPEcHofVwvQMZzDjglo71JIvWzd6ZTGaiOj2OKI8v
6ew5zEw+Jo3W8GePT5tGPOyQp38zzy5n9hjwlzzx2/aqy6BpzPMuBt9YvTfAdSAe
SWLD3ySX7sq/FPjVYKui6yjuW0LzLxv0cigUGCyBBOBRibLDgbZ+aWaz5EEUSHXj
ECLq7Xb9iBux9niyOZH/PivuQtssAXgOEUUBlRIfOKr4aMi6GEflhbWtjIlhNVpk
8CdsyQO3MAPeJXmisSugNg+U337/HoAAlmciek+qz0ylYER9Ce2yQy4+AbjW+rBS
WBdJMPfvFf0d6w6BzxTv99k0AyuHlOSDBl2ONEvupJqRlHJco0m+9H2B8i8Vpzs/
eOK0H2KkBAMxMz5qgh2s53apk1BcKeafKV78ylN9uNic7VmH1G9jp7OqrDDsMdw5
frZ+EkR5/5JgLue5FGMFgwSKXN85e+TnysBvR8gDa/hmyNuYja9kMRMzwVGWz560
eJUJs+ifv0L3cPc300GNq1Rb6zr1VbHelDbFuklbJcTXQOvE5bq5QzecDi2P1zjz
D0RLq/vr0kRnJagcNqYtZyH6cmWE0Yr7J7vju938brWBtpHGEZKhpnS2950wEOFk
poGxbLkgPEcNwHOJwSNBw/40K43PDJZCBxe7pbLB17OOoqidG353ORla0/adPooV
HPrwOisurzLyZMauQhdqpJeC5X49zaxZIKXnh/HgLuQus8GpiQf+TzUzOSJweIUc
B1yAAW+xNav+C9CtA2M0+WAoZt19Nnbmf3A9t7FP/SEdJoZF1FnwXXy9N8e4L+pN
lu15Tk0iV0bh3Z7DA6h8rxeXB1dE2bCcuNb6gjs3Lf5AAIMmMQeG9UCCM6vv9/P6
LjuEumjGuyKOdf4B1+2eJzHgaf/EyQ6KGOWYIA+hvzVtdyg/Ccp/hrM08Cb7xpJ0
vQa6XOn/p5LBkduo34OJpAGbNT3+dNchSG4mvqHkNO6fWjguTk8SZy2ZBWKGPn02
CCNWJpLSQzU6D7ffieLUALXa71CE/d2uSn/bJg9JaONzf1Wm0xHAkmWNmA4QsrDo
jVMVdCH++WruTlwmxGuM60ZIE32xk4a33FUKTUCeJ/xt1s7m8A1bD3gRRFBLJUEl
HMP58PF3wt3j3X50qzE+/Ffdl3ZIdERpBbBunO/sclda4M2pv2fgs/5tFkfTQe+M
JLapJrV56B5AVPTkIV2efHOnIxiyZ4Rq6Hg4VxJ9mWFPgbgy5mMBObyWjoXmDnEV
QtfBmQmW5h+lPXbnmv7UctqJmXgbjYCGwrACGZ7emxiB5GDJg1J8zkMePWwXGvAC
Uo4dMI95x82Ctsv+X2W3YeHNuvYb4nq5fSZRgHABn5w75vDInIq23Mha7Zz7Wp2L
W+kSHRhvHJJmhelDut39Ej9MlGJAWiUVMuXhjykOIoPS0QH9mRR28WXD1ISmloZ4
3A37JkfZ6z7/OMearP7ld3Ub0p0O2TDrasGcs5LXH+zVdUXVZTfVEiGgJGKhrHbW
uGvABWYElSNyva9IgltWf+iB9KwLsBFbH0lzo5wMx+Q2g5Q8iao0BJPKeU4Le8U+
/Pe0TfVRLEBbr811805NbmJhfRmLiZZ543pLkO16UzT/9CR96kqw8ujAnQf6ddRE
lpBxLDIaJt48HVCNrZQdngZUptdKh3+3vWT8QGSXYu4fD+98OODqczycw2TEkuhX
l1+vkVwyuRuE1v+P4gc4Gk9iGmneJxdZaBL6RAFsJFhPOxB/F59zp4KDOFuthDxX
9pbuOSwbC8Qa/+voEXjLaz9n4qQ4RFyxJS48+T732xuJsgGDMN2JwTCIZICOwypK
3ambMwH22/bA23cdWprioM8cKseCEyc3aQNFlCukPI4Mw/m9WcdJq8ZbgB87L9Ni
EGC+daPAnfZHu86HZTL4QRbX5J2/VsOKD+0/aQx7eDVF8xdM5SFvWh9hP48dJ6V/
hGjoERtA6s0N16MpUHPQtFHSRemxYWlw62PZSRQcWSlVEtdmtIyNd7pnDNNHlCNs
8hFl3H1rZ2hPinfKFxCny2CEz0KNB779WU7U2btR2fE8vO6017j4zgXOEjH7p9fg
lIOstAwlALliMEiLg5W1A/bb0zEPfdDpSho9vbu5hfhzzuK+UewwiTiahxcNT7E1
yYlgMonZhkh0Boh2ZqxBouSlEcOAu3qduYfzihPycqQy+BB5GsXRlwNzg1Mran8T
U1kjtw8MWFGQsGUtRakNSVNUhAHlx1cZ0RdG0dM1Jp3Es7+FL+omhbQ6he5knn39
+tK8jw3KYWDCXRTyNc0L6HWefq7mHe530C8JyiWOc5YWBXscKHsZbQkl4vcEYIqR
+ZyiXNkGDpDxmZoaiOrkkXYkxUzVwdTpP3G66BauWVUBhBEoKZw3fousGc1mxKS0
9w0/I/ojB82OnK+q/UAfhQe6W1PHCHpLQmlLDc7Epj3QvSNkrGvNsGyDYMSShoZO
xQHf+87WJ7IbP+zxouiZ6NWRcJjSq37Wps4jEI2qZgR4YnoWaE9/KYwRAcglgQU7
2HZqbNXl0nBqJP3o5Gk2SvKN0HHfpFNlwdo5qQuu1u86GuwPgeypWx8w/QDoHdG9
m4gnLlQgJMr8/547fbc0U6H1D9M2jZeDXRHCHiCs+GKp5xhqxIoZ15fT+cNimudt
7gG4Sq6DgO/IEY5V0cVhq1QPYSekeqoyiHenimQN6wFlXBOXSYY5HoDANQfIXcca
5e3EX2ZhvjU20FexREkKN71AXogfUJ2UGu7KQ1pSD9/UYCvAo0OMABLxJ7TPhpIc
qCcm5vHudnwyfCYg+yjA6TQa7z2kAgPXsIZKHlnuwhl/8eBYmDVuj25gGTdeBF9K
XtinKT4m0KsM+iPBYX/iokphd37BjrinbS05fboD5tB+6cjpr0/Q4i4gPpsFFHrM
IclDn/s6PXNPU4doG0/jODSEu5THO7p3qTsYiNKwY5cMiyjpkkn2C/7jdV+n+z1w
SgNaBWdogprvyNDV7b+PCIE0RWcXvLZpLoa8TrzNXHmUeWUFT1jtcgZg7AKDnUV+
VqTcwGoF0nZ56yEv1Zfn4nXq8gTxAMWDItp4+BZNr6r+K2J7TNef+mdozzjM1yCn
DisKuzrl4uJTuxPTM7KR2qwdXsRuP5Y6xmB+5D+Kr9bBqZw8PgtWZU10CyfoBzFw
CFO7gbKw0rDjSKOaG02pejHoFPHI6a44seMb/oFoPesqAGdg0QBE3EuMMa4uk7RY
JkQvm2+q/fjfCqXuYJUaRBP8tdWhXoC+npHjMXbkRs2VB3rELiSB3PySJok9NFWb
9I5wLgQTg7e0llcNurKLCIr3BrPFt5QbmP+GGLoZILJj2sjrLkcisD20uz7oA0Nd
Xpt25DNV7XTbmWtTuG9vUIeM1WtGfYxYIvblry/VmqD7z/nWWfQA1SUjCB7jB25X
JrXdKuw4Gwa8RlprZk6yKhOr1VwBP4DKK5qYKfMBp8isVTO3iqI3Q3Z+BeAOT++W
FIU6zA8f+ZtOoRUvAYt4FxHHmWl7C5MJgECvLdLZaSAYMtdcDO8SypFm0opDgl/d
HFXWZ4tBin7FsQVQAi3fq1J2So/ZEX2ToJjrf6uL0Gq/z2xr111shAJV6KgrEEtq
41FQlC6oTXmkfKITelz3iBGwT1J/cwgWUzHDVa6Uuub9BbQMENSTOPobx0H4/Yqg
+amQAnnw6hQxk0u5Jan0m33BRGd54TcELBw4EqV5LE4HptKH84dIdAqnA2tmeuna
IZYquiJ29qWASOWGbeRyPQ4rSsyj3a0KhGNStwb3dNs4LrkhHLGv9eEJO2i0HJl1
DPSIlrU7axy/7iMc+oREBUdx5T5ESZetOrOIue7nj+09XXgUY+lnWOsnAPEHIu4v
uL8kyRnhtTuHXArQlwII0tsepuklaL/2scf/koa8oUJZr2nTAv9jA+HwVgIdMJRN
BTGyx0dSv6Z5x8jJQ58shCMYopWBa+czHiBSjRMbzSBBVoN9cWhAj3pKg0nJeTAO
Qj3WGjRXvbS6xnBOksXYgBci40a0hQEsM67snipIQWlzwpQqJN57pvlvALnkuz+G
BQVXl3icef363ctmJTAgJwdRWMqpNlT+N0joJoahuKYrM9kz8ig6BtqmA7SThd/B
SS+y4EnOoWol8hrofn5wsdNfy4xZyOO70+JbiFLtIk/+WCszFRTXmqoEw41pVAm/
1cwrzRCXe++zECDA2YU8yoOiVtBzph9lwx7AiJKrcOvgtWfWUMgbODp4qohYMtDA
1PSRRUS8EfhvBF2Vu+roqiXbLZ5q7uyVn4eLnIbsE8No46LGDmso2avUET21cMMc
onLhpWkjNM2w3k75jy31jvjwSO5OL4RBESN980yF9Nb2lSI4W8rhXfuX+4LES9Rl
zSaZNb8Eo1HXbgr95HktB5gSYJIxhDClQynXV/0KcG3NNSIqFYiGQU40j0yFsL/q
iWUUGxiVCg0mBtRMlzCz5ikSvdt+gQlSvdAF31hmFAhlRsC+tMPk9sT1/iIukoG/
rUAQ/eIZdnv3vFwvoXskjmVz/qMgG7uK3htjZAI4K5YrsvSi1EFBW6Kh6eY1WdSj
ofOHkzSFGTs9oFs+r5r9/S+zVUOQPeba0gk844Kbi2ieB3LoOd2jMs7fVh/6EyUU
ZtKDj9F32c+t6NwkHGjnBVnY91ZtEE7BfGdAQtPxqyPP5XmtIHqH9HicU14sRxLe
bmN7u1qeWglWFFOv/O8wb+trIHl4NKFiNOG9l0va9wG/26PkvHi/u0IBDXZ6OeAc
koTcC8sbDeodi8dVagK9S8MwcTT70/RwfvsC9qRfy82lK2Mr+33ANFUU6zNSUfEx
1fvdKFfcP53ioAuNoyC6T+WFbyKeivQySg//7m4aKcsGez8YThuBdIqLCTU9oSdO
5R/GtfB3712bm1G8WbJrfv3YUTUXgWr/mfSxvcpUaajLlkXdOa5BTo11/P+cMy4z
nO+H1fKvXYdoqKSOm2l6+epU8nLb9s7Twf6IOt8/Zl5IN6NpkOPzuUbyCIEOc3qs
9B+Ub7uNVM6jEsr0Adkc6PiaWCRgd5qRWtPOroon7RBu9Bg+GVpjAkrLMUToTanf
6SuABYdpjUN9zAIrWs+2uUpr/C31s3I40kamXBXF3Gm8mWnGTgp0xJEZi6RR8dWI
ajXU5ily6dLfkOX1X5OoTW7Hds5vJzNpHJpCk+tARwJjNzJNRsAe7UsnyDUBDCtv
gV/GMItHjwRhvhF29F1SukcdZZGAQH8Oaz86EUfcM2x7QIx6ZKj51cnpJRftVQrl
beZB4EGzcy6Y/IDTWwgURsA3fj3R8ti/L4iUr729dgbMdU3ciYBIjDdvTMLEaai4
Z4hBa+tbeRTqXQ1ZO8f7gBBtOLo5SZ61nVF9Yx284S5Fn9GJ19vcluIW29Zt/dIi
Of1BwHfFQiZnebIlgwrYdyF/oSx26C96HTE8MxgJ5fJD9/BsHMaXNkE5Q+/kkWqY
88qEVuvlVTW/bVzduCz3u3ELdx9k4tL3iSnu2aiPdlYxitFwmAMVkXF9AQdKgvBP
FOh3wa+cyrhCpSKvQDTVBuL7FFN3B5DujzXdSAD2WTY73/LLNknLInmbH9P8PA2n
a1tmQfqBXcW/Hl3cSx3KHkOCwKJ/hTRBNmDJeIdXiL0FRUUewiU2m+RAPxt0qObX
0JFsCSnjBv34FCZ0WeUso13OYJ0G8mmCT7ubeI+4L1ae8pG7N9NlwMvFa4CtE6q3
CxM3O/6f7DQTGAQvUpYzH7AKSXvj1kFyhpDrsv5CUV1+CRN4d5DyRvd3hFDvXBQZ
YPRxgTFP6oyu18g1xF1BMHoOFhxIys732i7N4s8+uurmFL3jG0Qm8ozrSGpwC3uh
6Z0vNJTRNB8M3vnjOAF55VPYReSKsinPkB55ZtNj+6/SGkIIoKJ2GVn8TkLknEAH
5Q/2J1NkRsSiYXRBaOyj24ERmogNprdk0SYy78+MmS2Lftq399yNyj6FPrfyyQnh
XaJFTjgv3+lfQs/Z66+jU/WsP/PHG5VRQ/2QYo3OfNhAQ1FuDLTjwRB07z2rIeD6
6MHes8f/izGYESUn1R6F/h7cxp5OXbFi6DH4m09YgR2tQZIC6Lu+qsOepRZIB9+M
o1s4Y0ixRKfUh3DOSoku2hHhIvrew6Ku06/Kn2BXtzbhtIVbvmd3vriaCHg1BGrz
XbU99U95ZQDnVXJPZ7EyWZ9H3D6JtWtRd2CeQpaUtqPaVRMIPWG3Xe6EmIWIZMbr
IbETSZ7evZnVE5FypXksrh7lOLlOnS4urgLPFT89Ya82e9MqI7f5XSqxXRGxgV+a
qm/equQfKNu9/V3HUalhUPKXuC0KrhfmEuUSKEBph0QAsAwPUyRg0pJtyohAElQb
86LO8CM2yg4QUA/Nqw57etj4CCOekrGrpTYXr7XIztPGDwA4dVUAJyhYbr2iH8IV
qB52g07cf+iD/e3c7AlvmMvstL0CZkEGtgwBveK9q8w3Nin639y3HhCepwV/F9r/
cFHVNNp/ccpeiAAT4p7aBYbh0xwcvHqm9VHO3xrTiheHfc/dHZEOHgjy+cZl3qnq
kMgYNdpS5CTjMLApb8E4pC0MWaR1sQvLPQUij5mSgr0pq3Z6buZRohTapNpxwOh1
vZYol/v8PtyD9mAS4ma2XrAB1iZg40X7w6gxbJpwNCiD84HyTnK9y2hKO4lbQ35o
5BP5Ey7NRlwRbVE/dBpPbvPM+SN10Mv/PhQIBQS2v7rhfGyANiny6Dk21kB8mNYv
hakfA0ZaJDZH+VzdskspzVV/0hjceyorkqoqOeOK6t0XC6prHtCPCSCLIrPpDQ6p
/IS0An9ukXSQ4YUNqnkv7rgR5VdAnM478ZTJ3Ms8OxJyCODKtWoLtfgE7b/xLT0N
YI7z80O4fydM1/Ca7XceHZ4BC9uJr8hj59FYKNURPvP8QmBCtH28lvYJG+8Qrxjm
z/WOlOyfDwEHEfl2V7XCI27UwhZtFxuARqedyh2SPAaNT4O2eOVrrCAxiuwmgcaY
/SLpVRZKxBj3PCB5Yr2PxY8E+teVjyeokT7ArPjIE9SBSV4l6RD4Tf4KFB1cw6zm
LoD3Y6zVk5QpEYn7c/zODOv7GiCntB/G0s3iscKH6MRsbNkcevb2M1ZX47xlQKto
Akf5WR+Wod0pn2h3BesMh9EGpFj2PFW6RSi+oQHRPOi9G7f44aW98aYWGYYIcEhi
CWc30hNKjRshI9irPXeC7tFnmdVw35ScKNz9Mk2lXJXnpBnOqs8FY4Yvcd18jJAY
RDjofQelYWQmTswdGkADUtez5byckg/ITaQIRiTC5WY1dnwhT/Uurbv3MrvJ5cRA
KXiCZS7juUQb3WaPiHhIIhKE/FjGsdDFE5R/HL1V12CRo9ABBGpIq+uNbQBIsmO3
7B6/jKJ5VPS2OJxirLLO4h0newluKOrR4cz7Pwns36FsQGI9PXnSp2MWqP9vDzBK
PHgGsioBUkJAic1i5pnYUpndH42n/tTFuH5jX0NAcjJsC8nVfCSwtutONROKvXnh
fwF44V1jb9pjcM634H2ejbmY4sod/KKZC48zSaMzTpFw01kqiajNV7VcBCrD35Z6
+1BDimlaiTLam1wvfhYpGI1jpsdA0xowchvMAQXAGrLEul90ZyLGpTjmgx+97AEe
TbUvwfP+/bZkP6USdiZ1wBtL12cHMq3evZB1LvBKhKs/csPCHE4g3rJNkSjBkg7P
uLNrn1quqPZemguC1NTvNqiDLnHF1Mn8qToEZ5BMXRhDkKIEQSMQJyVUgjfWs2hq
zLXHVJm3oA096zQlELsWwebw4MXlrgeCiIB8AyVr+DYyrZ1atMJ8dXhIhmNctJEs
D4Omig9rgP60l9fbepkCv4LzMYYCHhHOJzPNMQy6aE6unzN5JixssUbgIkY7LF6E
3Jhc+S6lopuTVpSlDnpQQP1OWKV5gxMUfDArWj/CcGcRjLuZYRg5IJdiB1y0T7ZJ
YP1O3a32PWeGA3wKJINc9zjhKWtVbJV44IKpkNvjnWG7kQD6T+OhZAn3yCrPA+Re
SInqRX7QdJfB4TbaqzWFW6qC3C7PbWL1//9BFjDAGMen7UX5eju3Mn9nC1sZYDjB
7s9q4d++ApC72/Ps98htjTDXBeanq07M2AbNxFEYM22u0fCGiXJmbYEPWVw1WlqV
kAUAzq5L0Y9D1wDA5DJF6C8fqe6i7itVNNSnKCba2KKO33tKzN2FLFJQADTYWrjc
Y2EoktaTF52ixfT2Dj4wSl+ATb/SIouSxnU8YUUkOvDfhCCpx2gO5+pvjfOAKoAi
2GYyGZz9mzWtrfeESYm4B9ylLTlmgbmKeIQAv63DGCE2RpRovPqDSUJdg96LKWeg
ZWK98ZFo7zubGtI24PYeRS1T6S6tJgAcoA8lwB/JCQtxYyT37RDaq9FQ6PbY8ttK
SIZiiac3oRTksnNMxp64BgM2Zn4kc+FV63q0yI6uORrM4B5+Zu4nxPyHSim0r+DX
fIoxZznCVblXNdxUA7dnVnHMeNq2bewLGpvtAeFsdi/SST64RD00mD0PWMt0WGsL
pZIMLFLLjqzk9hNXFifOuvOVgQd1tKOk0KyR2Y0zx0UCPVl0/5LHKpfqn5vIK67R
gYZO6U+qk69LdDy4JI+rBz+3MIeOXCuxg2n/U9fspGxTgaz8O9q8CIb+FMhYLPYP
WBVz/TFGG4qNHBlJxxULMcqanxYjS5ddcUuzCUzQhF7ZMu4oCF+i+ZmlfHyUT5ro
I2bjJvveIRZesISiOWqRxLrvcYOwF9pQ3lZr7zbi7qgyfTcZFoocMABgRQoQIlcL
SnsAcuUTSJljK8aYEVTJcH+XJCi0ZSYxJvxK3HWkMteqGCyuPbYvh3fJ1Kfx0pw5
IsxOHBzVCi+KSAXwrT+wkfFZ7lSDxsQagaUF8O8OW9itcHgMi3n6aK3PnqF7UR9V
nkbWyMRJoKuKgKIubFsBpwTK64M9DGpEPG+iiI4pcdC3G7dGCgdURYjEysj8qNF3
mOabqHIEZ5QB7RYpNt4RRZDobxIVzRiFuu6i63e9Ep+F3V+Q7Q0z91PyMf/bPB3Q
jFNG+PQUdr0NZFc1oJlprjTrBa8+vi3H7/uYEikvwHpS/GFqKct/NaCeMU1pw3Xf
WXrK7xwJmFaMR3PKLzbuV9JnLm2Q00jSCNXKS/Ltp5hKly0E2t/8HHWD4/EXSjUE
k7p0LkKlpfePtt/F3R+N06+xFzoysbwwrE9jxdcBErav2mD1oP63nhYmODxRA7eJ
LR/o+WqtPQOJilBNgsK7nX+nuLVyDfuDwb6MvZ6yVMthm01pLt/YQAcMv97Pdkx7
/nPiS1VjyRUDqFmDpXE3+IueX0eg9UUsAEnC+5vITYqggcB4XDc1jz9957MkVL3C
hbMYT6X+amynMSnTiPkYwPYR2PZ15W4xU45kEsXKN9okRhIHz1QkYWZ80YZf8RGy
mM9R8kPo7lWD4k6FIs951l2c5+CDeFCB2c0Z1MTmh11Nb/3yg6y5wXw3eDnDfjFp
qLEGw3nG5/vk6lJl4afkcQhOVKa+lvWaIeTeA/2RSDlA8KU1RPGSS80AoBNcm3oc
p3eO+dEV26Ncyj4tBN0IsatfnVBUdAavx6d5hbARTpORN7Tju3X0nvD1Kw8DGNTa
GvWC1tOCbiFTpAt22ecFsEwJxjjb5cL2rDTSjbXeIxtvtp9ywEMurONBs4g+7eiM
NtWfpVI9vaNCJxPfo7giNXPT/WFEqhxd3ZrQEjqAqNEu2NAmpHebfzHE3K5ki5iU
YgXSZpnxefv6A2RufCxYr6+sTyd7JGyrsPDkL0G/Han6feb5yTgE26Bwdp7extLH
E8JMvBFhxCED1dw6uHgjihL02g+cXXtQRh8rSL5mYST9mQrMlGdAjwT+ucmE4l7e
YhYjK3ujCXIDBEWYNLEZVRo4577VFeCjrZvauqcA1eWEJBFLIH9rUWLd7OEsoWW+
9wH4eGhFSXi3fPIQysI7hJwyUFiPCQ1Eiw1nURGzngeLgCIt9FV84IUWie50S1mx
p1kiymLcyGj38vsKS/iVayfvkwetAUqd4vQECP6U6UO/kKUZCdG512Wndn4DXNLA
8J+6qjmK9vf0/flWBVtYnoZreua+ke8xKjhFMRQN+sDj/qZcWgKQUuNKTiQeHokb
EaHugnw92CTkvhEMc1DgArwaXPaN8ph3qYVSADj4XIdtz7fRhFK+RZJY2Sgsi7xZ
oEkZNou+J9NjDGrUzb3mKk/XSUgXhnlpdLh/IQQZq+0Xb15IiKe9jgrONOBrmYwH
UP62/Q8kLTVaqeCD6v94HyKhB6Ji6lMQUAim3FgtV6zFeYRU0GA48zYEzMwl7c4C
kSGEF+BKT81PDeYCzbpb2y7ItqiRo71g84ICFS5JHuWl12CSW0hASsekfJ/0MECz
ewi3HEGpcyVJdUDSGui/GhwvuKdHFnQ5cwfFj6y1zHnkx09espU/pK/hBHMJS8SD
sVwlG57IofAzrQjusFcDxliSp5Dnl+kPOoMC81pqw2bcA6Zuu6PA8BSgla7b+uT4
WQKhS7h6asQYwvZ9JI2X/te2Xj9wXBbsVMHTaz4WmctFZppOA76VIcAmjT211iHo
MRBj6kqxwHR5v/aHbW21HF+ceTnEL2vuHxkwVBe5jGA5WeXgu5PGBt2XAKrM4KQB
e58UUSYPKpcypYTFq9agI8tnNvUvCP8bEBx/SQMWK7uYSP7TmK0TAL0g+UZtRB8z
pTG+woTJd2CZpTt3nLWdFymYEi8mKRLd26WtjoyWmgG8aYxVrMEaVbKbNCUr90Gj
OfzD630isVS+O7DXQsH/NQ9sA07o9lv1cM+Fl9mCRbM7a2KB4p8mj3vx4DVfhiN0
G5i3iWGX2Q1lTeVMvMRF4136RlpLO+Zn+ZBRs+DrA6+ge9jD/pui+I1YmOYRUWGy
Y9XHMJT4zJaufgU9NXRD/3IO2EO0FAGocg6d5OBdCpzhT9bVtMfF83Azoz28pYmi
OubOy+l2UhmTXPEJEAG6/G6p/gWFAt7qZ28enXxjYjdPwRK3hRIKziwdg1rMvOwH
QlEEsqPzmws+ZRob/Wn51ZjGR5UL1SvLsKNNpaPIr3pw9bmjgixQMxDIs+0s+ukf
KQ0x4Orkrt6IsuwlAAGmS5usk2vH+Ze6Ibfe0FK4VQ4b53ptU+F3pfQQm2G7QIjS
KWFj1NX4y4MyAiorNJMFdZmPSbdD/Rs3EG1nQkXXwRB1Idv8fDfT/+jh8IFlM4wN
2jTI5Tqd/bCVZHnPacIZhiF0cK8nQd5q7+/AqMCwLfa0ZgfgoP8nkE/TtkrOlChn
OvatjsRndlH4n/U0vRwoMvSF557E8w5AM1AM1FEx3ss/sWDtvVZON2IdZ6Y5AIS1
2t264bdpQBQrrrONi5RO2LlQzmu2M2v+2pbYvvWfcHbncGm7iJUfaztPmIcgK2H0
wdYVU4m+NWo6hi6Rasn5AUM/cSrXmWeVE/v9K2bclf0AXHckfj2Q+xW6ycpTeE+1
WBI5+bTpQ3WV3GU2+dqfkJcdgHFjGz+r9J9c7xMRBPUCTeV8YEeBxvGaIuo0DDIc
TkBjInKT9tG2+uv3m4wekLAxnAomfa2RjKZogGIEVJcaf3wpIxl8gg2koY4EIzzX
194/Ad8OXVciUWUFv5nq+NTRwAFijprpquHcTY3Pg2yb4DLyye3cdGXLLOUv8XYl
aWIHm/Cy5FfPIYe8jIQHjnI/NJeBol4C7pqdfyy7hIRyMM1hGnrchNxVRoyHg/cS
9zRHJUW1DBm0LXpOy8sYNAgQT5LbyrxNuOqW4/1Set5vSKpX42gB8aOT80BgP4rS
X8e5ZNOckNLkWGuRP2H5etDkfJNIwZ0XL43qPlSOAHVMODAf70QAuZl67I8hjo2u
jjRx153G8Bk8RQDcZm7fMyCM1y0PIyhmIBDzQWkpROZhgx2gOAVgxkfdVynFMU/0
1Mjv9whgrk7tRwvd4QD74TH6UKvcwSqgBjIKARN2Gd09GrqgrS2nlBd4Ncp7UsCK
6j3JRziBzJVBUUKC8AN/BeGQCWbEkk2tvNi0WqAroqyKHvmnCKsrSsi7vuKihVCH
RFS+MDH1LhrDEnZlrSWgp3t307vcaj0Kifxt7xEm3LPsD1Sgpn8m0C6IdeBsS2wT
mka8IE0u4eLFQGQFFKX2lkB48zBP8EPn+C7PJhWDDhkxU9BDxJFP+NChFePxE9cU
kLiSjp/VulrxSwJGVc5lkLnv4SMEVRqi/iMSLL5Pv2GYL4uO2prumN5d7qLqxZmx
6OgB+72RyC5NUMJPDSUoSA6Ba2M0J4sjdSyX8PTwIy+Y2AsweMWF1Wb1lahq0GnV
tdEblrU6gSNURGFK8Vp36hTM7Ywv38xxShy9AbRh8etQd1Fij3wG0WPEviG5JKvt
lVo8kh7mF2nv+VpeUrGa8oE/QrOpnG/FIMpDh5I697ZaOJUZ1DGW1iU9poZG5hZW
yrqTDUopEfaaCepHz81llJBOlrW7we6PYpwZ+rsylhHMiuyBjFFEkgT/nWQrBDs7
aWzAXv+H9GPhK9ClYmrNpCD3rOvDS8FlM0CH8ts0UAZbPAohrGeRh3eHFQOriv6A
QR6E1mlrRuo1d1IsBBZ9FhR5TvFFrrdE+70OqKHaZIEd916yYE1Ky5dSwA/YNUHV
rkEUkeqqvQrqK4sUZ4TS2deTwcpa5XmpnnGJIiSO105qzStfJsjeVhL4FaL3iDuy
WVo44eMs3dW1/UyyT/4fy237tl20WAvmsVDcei/UnNKNpjy3E/hZVgqL44ie6KAT
aFWo2vOZSmB7DfUCYKZu4Ag+lD0UBtPnrqBsohdn0Y9VOpQtE4SxVsIVbposnEtM
2GERhM1FXy1HMlqaiPRljhsoPz/YdWuRDWze4khXgEL/dMrNvZkcLgbfeqn9wcrG
lIY1kO3h3LRqV5ZC1gLYhvAJ81jMhaKahuyr/R/SI6uG6mquk7r49NpA32YGuYBl
OKHyM44q5rVLTqibZqiS2V208RGkqC0PVU/BvYxY5LRZ22k4JvNWGejzs/f079sh
HUjiyTVEg91WX6SBDo3PHOO6g+yHrSkouTzeXNkvwijfPA25aMqOwkJK9zCWw6zM
xWhOz2P+kkmXynGTN9l8INQuSG7kmd9ycAPhJMEiCdwhsLUfHoHtj2vGQ4ygU5Se
aEwUQoiseIEC4f3yyKfi6SL+A8Fo85zooxSCdJ2CSjerZApfdQPUiOPuxRTXC+EU
N2SYLdILW/+nApRkd2nAyIeQ/ClOKayoP9JGZepaVt8qyI/ZyTy+WB1MMlG71dkZ
aQSkHpKmNtNcPC6KXefdVK83b7jOy7oDi63JAguTvxl9vuq0RcG7gOPkokZ6GGqE
k2HEfU/9d6mp3B9Umgfh+yWbK9cyK6wMcAuvyydlih+9MI7cpW+Tzwe1OsCrbvM+
/zLHX91V1r4380elnmRfLYRA9l/Xj7sfey0YvSbTh3B7kzOjJWbKiWyZ37OdnNk3
Uwb3XQ62oJkX5NBDR49U3Fcuk0uh9GeORt4/dGxkin5X18e++zM0HAzeiWg6rGFa
GeMDttd/DqCVELwNa+61/PzMr3059aVTepfr4S44AJH87RpkEKQ1X9A2/Q3We6n+
SBiAqa413/kg6nk6rqcDcp/U3pAckEhV6Xwebr0ArRDXSTvkO3CHBbYw6lzT9h6P
9Asz++6CHIrSWw848NxXCb6JgYiC/4ZSNkaSXSZ0c73IxdZphWJxnRSTMj4i5ktz
MtEyFiQK4e+WYDzeT1GnaNwYelR1XsW2Gs9PDemRbvd3m04o4y55MK9xub4WBbin
V1wfjBb1mVaowNEA2rFi55SujlE6zh2SQ1czqy1WRgIy12g+rwLHZ03vuP/UvJZT
wQEZh8TEuN/ikmaIkxiMqbRagH+IUfTn26y5KCj/411O5pf62JOhw34MIhhlf4nb
9Wel8yn2DkNy4MUvsYaHV5VlJQjbp1Ge0ds1eHQghsJv3b3bf+5Gu46/eC51GN8R
2XHHZghqMxKzVKhFy2HpzNToy7P+vZP4hGvKl5Kq/vflmUa+IL6Y1/5K7H/Nmvep
ru9WbMLlOdTRxEcIlQb5AlMIBViiX6/p+6WFOsccczucClErM7WdxVd1wldedUaJ
SUoXfjiek2DH6QSxacNcyfd7d95rcYbXh6PKL6wg0IxSYT2FYNxEmLMFRxk9eL4e
fTE7NLbeMp+U5Aumb8b6j5bS4S27HBMcEOpwW8YmHr0+rsaIPCgi94poGAvShOgi
II1mZ50gdXbKsBMPL9qvdei2M3zy/byEvspiOSNr8C3eQnytD4Za5n4z4Z8d6LO8
g00XOWVooftUY0h1GAP1Xie7Ll+7A46JpZi+3V4RLZMM8Gg0DBY/Cu/3bcZMDnkt
0o6rrlPSrh25k2KWZz+5GlSxQDxJMT/F3ZdL5P1gNwhvpDxzeeD+x8LexPjpokCt
Pn95giLacjSd+OXsv9SxO4JjJDLML57l5rKoU0LkyWZ0TauxW0XrZOg/vMHfXA05
BvGYDg5+K2tMv+sTD6OZoMm8hXtJ9a/9K9U5rgXip4yjXfcM5vmQvyWCWGL0GTY6
o+iYs8K+gbPzQ2H1gGwgqH/R4FN77vuNrYooEr1Vu5Pfsl6UTlzr4GY7bv8B+rnB
laJFETRJM023F+mRiog6vi2qJDsp7hRPa8OsPiDwgy/0HLB2S9nwvSPGDgceeNr+
bterekThI3YMYgfYDapo0zc30hqiClYPcsjxeiVj9nfCfbUYQowzbZB6J4RaRMcl
HKycGNEm6+WVg4Frz0Uf4csLik1nu1Eapn+lP2nka58TNH/7jcTHD84sqy78QCCM
rVKbffoKVAj2CRxfdCalXxQ7GrAkYiPMlvccItGRLqAk9pbt4qPc8UuGE20PsBhZ
P5Cp8lKgcBMar+YRbwj1X4T/2E7QpkIeQP9RBwUgScWi5yzTylOz/sQIOL/agaPy
qcc7I7EQt/cIT/lLKHHFSR9q2n6mVkspIXCZIjPfq4TDQE7mHCOuUUXVHcKJOdld
wrw8pU8fhNVqX5upIEc58EXdI08DAlNFPcxl381e8LRHrWb1sfRCfwD9HNZlv2Zs
XlxpvftNjiuwGQr9mIoZ82eKh9D7jGywHCGZlER6DMezwEFCazrW0AT+ILIHNeBw
5iHLd8FTggVK0ijpIzcvG1mAy4OHHQGvH3mv+crW/mQrsCLbF9pRTpQpLFPhz8Rm
FuLjn1FWJ4y2osuXb/NuAVyJ3/NwiDj8pJrKw7cFhb/PJllR0lU9vz++xwGUzyPI
Rwa3g1+QvhBHGTgzrwYWbB1SfEcU+O5TCWgXm6Q83klQF8vzaTvEsq52nds4xC2d
pXUxItHI7/UxiJ5NSKOhkHRtJu0blnU8PSh/N0V+yX9U9TbRgzKpsbiU1MD0V2rD
9lAoV70S/cHOPX59tdwtRfcjemENpBWMmCWGBumKFKeMaHE/qTydFUNXXLJa/iwU
uaLwygrYkvfrwrxs9I+bJ+iCXw40iDT0F2LeAjz27izsTua3MizCe7tCfT8GL7ND
WSioPUd+2gvBuppciQUqkg2muuBlXcZiw9LN+kSRylhYJOSB+KwSQfdhI7FnRV9Q
HGt9ewgSACTbts+wO/mI1GmzJD0W4DNExxgevdWaOcZDQZnk3+hLLahje9lMLubs
nw7szTOpYpntOU59rp5Nvc2XpeYJooFrSiLp7S/qafRmryu9Bsdz5iwIYxgdTcHL
bJK8dufzYw6lhTtpsB9NzXOrZ1YHB4DHE6LUGaktVJS23Rxmt11ZsgQmrOTIepUb
W7tmNpnHCewp9Qr3VZSuV5qyjJM79bFXYKdU+OLvndmKst2DnWelKqpNplMMsvvR
K+iOcbBTzJwOhSO6wHehicB8o7MW5DmaV2pfpgtyG3/fLlmdebJUg4FF12Z44E44
vYTX3ozZd/MBQQ5hm8EUpsdfGxsKrYSeNWRI3KnnLrEUj4PH9s/s/HJwMCTcJ/bo
/Zl9gOyqgRrx2i5OaXaCvpmiQuc5wxxb4+E4v5/Hms48gBSfn5pBNRh06ylC/QGX
v0ONsNKgj5cK6u9z3BcMbFK+/e+hW/pxhanKEbTof+zr9AzrET0hUiginr3AqWdc
nG+yM/jyP+8+MFNShq4yY7haArOazq5jMoWUpzsf7qr4S6tz0qHy88XlEN+hi5eU
GKx5hSDLf5DOJLDQ5w2NpeK/1EOf0oRyR0c6vnDxXxcpLT62VprcYfWL8nKP/emt
5/pNvpQGJdOHul5BJGDtgW42UPNIpaOAaZ472alJ49GD8UguirZ1JuRKYAv4CMCu
I3A0MyNrMRsV4LdfDVTijS43KHWJw3BeNJdIxZAYxo3d7brnebnMsqQd9wvy1Ulp
HI7EMab+poplUrFTP0O16GyP92yLvPoTcsD60oZhU/3PomqNg1BeHWGZrK+nn4iJ
lDYjRiSp/YRH2E4Rod/og1CaixfYgRDfqZR1XzK2UdnE/2KBZZmqKE4ogZ+4vEqn
U/B5jIoj4mAp/6B6yWhV1lj8YjBueMmOk2osGDm09Irvr6aJwrf18Jm+wRhTB78h
n9WEflkVV4Ed1TH1OkW2qNSvlVIrMLVNHwxEve4yCQMq6QKJB3BgQF/hFrz+Q3UJ
f7Q3iTKK+1UP0p5J4TGyxdOijitwMOjo+l6KnZZ7J7jBiXCiXlJDaawoeser3Oaj
5KcDluZSwwTzhCvEsasGx4AxRV7JtJkmnHTdtStK2f/8yT8c5PIVK7+ANCxSErW6
DzW5TSCDeEx9pPqoU6tXS9utSV8qYZoce/ou0DsiKVsv8JfmbZonorlFX/N176kT
aMV9iHVBF647+1iTJLDKS6R+8/qmpz4DtMccLiibUicuyc/OXkgjR7fV/MVBsnAZ
d9cLewh/He089eNai3rxHMpMlnb//u4otZF+2mP6iSz9KgVqYFXUkB0Mv1f0v2E6
1JRyDkyk1Qba+S55HfRv7RxFRHygnEDUzch1DAd7EKWgPJW9uhulAV+KliiWC8YR
JS6KPg19kBZo648H1nU2F6sFStFM0EvEyXmotsTecdg70ZaZGi5WFy7BGz+oYExW
wdMb/HthBNbnETw3R7CBSm+Rrb+6MKGBUA+PFvQ4BrdNSt/a1UZEEPqjDh0lTWAc
YLJwW0cku4T5PQXEJNoAuWr8IaN/TuVek8t4fFs2VaYL2QMg7dMX9inxcjF6l5Tk
CFHzrhShSvVKdm85mhVeRjux/4shdm7NURGVnWG3HZqAYtDd8cImFmyz4cDQ5faH
w7zuhfJ/N4ZJtnEJvthsGx6YqenF4NyVVhzx2f6g3GgfLdTcmUxrVkHuNUkj3t53
ocjWmNSlmSaGk75WgjR5Ju/RRKXkN7Z6pdRVJy1FQcOkj46KkcOC9FhvU1Pu54h6
N2echgH3yNFIwHyFpeWDnbC1yEA4Z/nGeeWpL8NkNf8gA6qseNhMzBaLIA9lIFNs
/cO+yygXdEuIvQxqifVQtjnPFnHfLDhydX8TBZCyXEO9jQWIw4XDb3uo4ZoUfgJ+
tOu3ri6BGeUJUbQwxaXnmDfErcGjydKyy4N9GaQt8WEyTMgPzPoqWWq1bB+riIkE
n5So9zbYZlWQOSFJVLL2xDtQZenWR6Kg+MBCWAXai9Xb/syEbO9h9jwl+pxBLYLq
s7ZgcfYFI4goqNNHlg5B/15wiqOG1aBGEEe5To6cbatD338VhnKKNislysEQnvMx
J7jdxH4bMKs0zzhbEHi2YtdgUFP5p1L4ouiy2r1qTyi9b3Bfk/5HohJZJErVICH5
+KBfucvkBpM6xQJ9FIhjNTMP08cmuWCbjPNGg1OWCfDvLxJEzk/r4fWPuggZQ3NU
251Fj8J3EYsU5eoP8925ZMTpchmqmHHeQOaQt7B42fDhQ9yGiM7O8/VK5LshYRD9
k3ctLnlH6D9hOe1iOSy4NJqLRUSH9kwEzrw3BiJJWpRb70mPiDPqLHevGQMEDTt7
g7jEYyv91ocCXnHznBk2uewxt54WCLUaUgd7pBTrXiT5rAgXBbFz7NcxTb4diVDU
ALuOAAQnOEvWPgZuugUDbi8OHF2A7S1hFzPx70eokCM/VNmP9Rmg6Gpyp2j3ue33
FQcQ+wL7eOkrbu1yBPO89eiluEVKTYcxgY7EVVvSeB6qaTEp/Bw9HJkmmFhcWly3
iV+MktZdipvlArVHQRS1haz8wNrNPgCRhK/rz66wuvqoVD8mrHmYutP+EHChQGMb
BD1FEI8xLEo3El9BkkQWIluDAK8OJvxK11Ql3CC/iseHrc5Z6X60ByOorcB4uA8A
Tg1lE3d/cHLPSV9TbwxbMsomytG5X/2J3gA2o72DK813OMGOmGS9W/JUtsuL3zPx
ZdPogiN1lTdAqipgUGKexvpWxyOctlM1aXQJMKfgpASOqPLcS654HztMKWClZEga
+GFu8YU4Z3vqxykRxKeaVHK8vvP7WnSIkI6nyeT45um7x8dKwPWmMlTBF3i1/rXI
90ZCySlUqJuok+7USILUc+wl1dWSTJ4OlvslkzbVKqj1W6gjg0jj1otGlaoXd5vq
xGOBFYF/lOn933OvnOh/LpBKiy0te4TFueHRz5F6s+nlM67Rm9fyY5wd/ntSdmsL
ENsxBjTDEMFsrLaroezNpkvAvvj5H9FY27z7KprA0EMEjTycxdB7V52EeZXdZ2Ec
RP/nU5yDZgl9XwR80h3Dcbp198T9Eg0CFEVd47ZkoG2AA4Zjp7aaJBLFtmh898LK
c+js+0crYh3e7/5AWDnE1lzCUo/pE36flPlD0SeOBfiIpDWGEVQpjj8fIFr0267Q
eThj5CFJrgUQuc/8OIagjgHHk1oaDBOxo1WNkp8Vml5K7LGAOomZ0duXuKfMieOt
zBlEI+Xo4Mug3xWFijlQ1Zu1rrj8mv+Rg9RiH3dIB3ustU6rvJ+y90Ii/xC6xxcU
hiKn0dIUwyuVLqXEtK+MMtrUkX4712xWK8A+WooO1kKyAINMYr3ujFT7ow8BHknz
DQvAt2jKjN9rVORnQ2TPX6xYE2+R784vEsOTArByMMGjztlFp46a7fXFFNqpxI+p
BSUOZDV8Erfh6V20Pihvj4a/YHr3M5fpDalXMU2epSj9yxkDt2BhrcZp1CCq1Q4M
BbmMox866zaHnykMHVAa+BzMy3xQ5L/9ryVLHYfV3WwYzW3f+mMlEiYTrQF9lcNs
iIVDrn7gtkeJk1RK0zcGwE/rD5A9lJcS2vs61nUAtgm/N7Y8Jo93dtOWMKaoSOM+
84Hm3KNHHTrv6/y9FVOfitL5kVt1/JGfukG3xdZzv8Kx5kmx54fHFLNpsOhgIL0i
61VOxqGyxCMDJFLbri7xaLkoXBQkjza0cJZ01Xk4b+kdMjIeuWu9Dwym2CJ7Gvk9
CGRv7smbw+nRHl/IWWR18ylKMwZB/uE64rLWlv2HztJTBxTjYI2wo6lPtocIpWw5
2Bt61gvfcpILsFEVEKktxDJxCGI3NNWOO1EzFk+J8axBLadiQVV48olHzsGr5tn3
FyE79soBVhmh3kiok9YHylu0a0ATot7nCoUQ4Gbk34k04kTd3DVC+SQWkrHB0sRg
IIZShgy7Zf+B6LG1N+YghNpfguKh6RiM0NEK62QZNc9g3v3S80w9hJ3/MxDa76Dz
boUHASnvoj/hXwfvqjYMSBoELtjNLV9m0cX8cCnU/EbmcEhRpOrVfhh4ebgCrslr
V4k0ezeUAhvn5u9oIvhUjh3H3SWip21Giu9w3q6DDziq/6bqfCeI10NM1Fy4iDlV
5sVpg2/ahwP+UaohmF+JYsrEJhN/4Fpl6niNpOmRk07AGM3nAY4DOndPDSoeanGk
clQnkkVvFIF7CTkDwZJzULzEj/QZuamSRYSh2CvElOU4rkNW4oHn6JfM6ZRV0A87
sbheMJhOYyhU9u0F3p69d/jCAD4kkHu5A7WsVwrNVEnK51+GZuY/aRrJs1l8ufsP
nzBe2Mir0aw08Tn72TYpTefuid4+LiLmJ1KmHeEUOMPYE8wS25gcnRXWp9oWJR/6
GCPeJHXxCHNVvDlgeX2KBe2HgKADgFLXnP0TVGDeh2LtVEuoXF0uftp1vXRO84hK
6SegR2gC3t8gDCM01dUcbeuqxzUQfsm9xwlE+GzySuxqrI2361RSnp68Ygcp8O4G
TKroRyakt3XSXcdoElmlOGY8iZa+KpBctfSzPi44NixhxFOCYp5CoWOyxwSgTqqL
8kR7JwiphyC+oVLjLt2E8azx9Yy6IK39nE6CDjBpL5TjKXJZgadKv35rA4sDXY3D
OEq/lpV9rSWSQzZ+JEvHhgPK6uaLSQttQ5L2v1Lm9gEO4JhBkP3LnsDreyFv1vt3
zouVbnHhS//6mzrahlh/ASbp7woCm9vJU1vHGG2xHA1DXcwEdFVhUEwyUrmJLQmt
qcM0RM1uL+J0KPTH5GF4i41sdhRci2Tas9G+peLBE+GgtLGENUEukFC9jZ2zAkGU
DF0fdQBODK/5dsdcEt7VPIvYHBW095SZb4OmGTMwJO+Ipycg7bM8JskZ0h2SHxT2
bwKIT2G0xP9Yo0PuziD4ce8WokNshrgevUyz4b+L+pjXAuN8dEk0AfSDc18i/LZc
rld55QPQ4NpPvF4pieXuoF7JjBeUPgFaHheGZHsLnDfSA13KfXHqAJKypCPq/Atk
C0JPLtV/kltHFP53JuyE0+aP49V/Zhw5SlCGCE7wEbx/sA28vuxQGM5ByhHyEIUQ
EMLMk5pPjy81c4RIIAISdRiqTwQl3Iyk+/6Tr7taNndIBXcC+C8eEKPA9lZK5dIL
iWx+4W1PvUAU1FV6jwyG6MuOslxrjDCoqW8SWXaCY10g9Ch1zA7sQE9hwww1sv/a
EpssJUJHlWY66O+sXKkzpTLvZQ0Zz72LkDOmSQ5pO6QAxZtUZ889/770QkeDHHMM
LfnAQvFG67A0TC90P89FjBYndlTgwLNjRmGj6dExqFRLPnWlGB2AFjZOt7Y6Iaui
QbZgy17RgYwOslsD7/L071D5zejQRkcgUh8BLbOBwstJzuJ80AU2zsHvDjALNDGF
fEX5RVGDldaONNaC2dDdIt+XUj3h7GIaSkpxbDSC9d5vbif3u3y/nmfIk0xPymvX
1Tqyb1YvNPgF94FREg+t9QhZPffCj1b2/zxrrZ8+Mu1L2Zs5m+7glbXfJfWxmcro
w+n+CulWYDl33rww7kZYyQ/LnREFMDuiwxIOH8W8otUTWBOnY3g6ylP9RGoqACK8
YUiEw2JoKuXbJry4OagwnNo3BPac2HvnF85WWzRpye/4OZywxhKwQPRJEyh2JdyQ
DkHJzuGxhrDVqhWytk4xCshuJkZ1wdNvLEQSSrM5CCb6LGScoCphIwX0ICqexjrf
CG7nhZ9QbXLGmw8apZEtiltUXEyEFzwwVDYcScJSNmOBbSnKA+/f002blFRSaRBQ
FgfpCDCpNu1RruklAXX6oAWSo+qDnU54eYiGJCRH0xkv9e9HPIID4rWf+tC9qjGI
5ailUz9PimKGlAsBzDlB2Wfdz2yAl10l7nBT4wbFwoazB5ZNN6j6IZGK8Y6ApqN2
rrTClyWyNNG1T+JvxUYsuwOJzBJNx/9e2LOljoNFYcQLWhyVkrxIN+1UHfeM/oVS
OowbOABcfgJagPQoeH8kqLfVERYlWnH0PuV42NjyxABL3JjHdrDi/9/sxfL0r5ol
X7KlJbILd4SqGDFI5a1aoI7okRWP7wli/OB09iMEuQLZEoXzDsTjYmW3gftTAM6L
BO61reQQJXc8ChTI/CtcouHzdhhT4FLZ9l9lGVffGKgq9SYZWIUI73lXMMM6n7M5
1r64b+j9KexTFrgJXk57qGbsEjHAVPfJTa8YNShdnlzUWuzBcVaMch/WXqxRyMhT
pJXjqKx5i3QDOtbMliEkZV1RBxp31npuycC0xzuz4nfCDtf0yCt1U97uY2fYAJ9e
eYNYczkfhutK6T1L8n7eWvur+oSeqL7ojEyNA2SZGSM06UX0Y4Jj3T9SWP7TbGZB
C4dsqEFpGwN05G2UWaUSR7eQg8R1v+Jimne1usnD9+pMMuWvhhlt30gfgS+7oBUT
bd9brH5Dc7N/MnyJlVgoA4Q6VAFidORMc9ZjHmTmoR68yWjpg5XjI5FVfVnluiGC
bZsVcogjHW/nQQLutGy/y+FT2dg6S0TM9kXFSrZ6/5I294dJY4mRbTsyrd0UqS9b
Stm78kb406Ndkt4+cX06aKswcBfTUvk1sQWyZiybXxPQU28p0shP/Kjf2YkTgp5+
OHUJO/zx2zt3N+/Nmputt/hzV8jHKAThlvUhy931QkfSerxIpRJ8uphUzh66KSW7
VkjR214kjM7HIkgbzZv4OoPductRy5ZDpalU58K2sUyO1nxZA62Z8rcKyKOJ9ZHW
JtBX0XcKuUZVSFCsxLb/aXIDXTDusMEy0V8yG5oC6LTvSvuzRSg5/Vsm+VEMucss
7SEElvcHCSclsIY1L3IudQyW8BN7fm2KMPFtzLCEX+waBMMsr8+hYrCiFKWKLGsI
oIX5o4Nh21FnlqqbyDqUmC5BAgFs/1ziosmtkLqHHB/Xp9eWOk/L/6nQauuPfXPt
WQjkDWjHetvGUyPzQyuDs1lk5U7x0rJf6QO4C5XSJKGtfKsJJ6tCGE2n1IjQR9u6
8bWr0p1sv1/8uIOXUvHvx+XdAcMb3zlc2Ww5/723j5H19zhgB+c3Q8Nwo/2Ox6Pq
H9TdP02MGo/2WwWXvWnb2jX0jbZ/qL8nxmpMyk/vaKjDGr15mLrbTIDmwkUPRAgq
+ZpWFWKksSOtm0qBtcaNesfPxCxdnD4lKXXustka4ITnOrzJmReveuhDowg3BPuf
zCPVs4cTe2TTbiAg45tfYB4h+QXgcIgsEDiWuEWVJAC4JrbPoUrc6oCDLx0JN8hF
HqdSTPBMrHqLWEQxy7mr1Sj7hB8MX39qvT3lYa/vfEdqxOXk3V1ZErogDgJFIIXV
o3cRe//7NH+Zjra0iTND7zwJu+Jj41linrDZcjb7yKH3260LH+AtlRZDZQdftJDV
CL08PuFvMRE5ZAE9y/jAxWvuiiyDE1qIzJYp78oZ8GFA1DpH2T4nTnKrhdlZWaBh
w5BB+eLg0AlQTkO+MRCIbnvnmo+U+Q0RorYJwW0d5HYvckKXngQrUh/Nzs72/ap7
hHY0PFvEaRI3NulpLWvJJoq9GBPOggh9OJXBfrveWXgZCeY1nu7YukRUY0nNimPX
dwkTV/LWGw6/i2hexnZT91sKo/jU+xD9XLQ4K6BVUnzjJsYSVgEFgGkx1hyFdOjX
VXC5Xioy7nnhpyYWu8zd9Lt+HqI2ZeGvHgdbP1CxDnnm+lrnEc0VNm8KuUwtTBhX
vMrGkM0z9OCi7fO4p2Xi0lBJ/f824+O8dhKzYGYC51jPoTMynEje8JnUfT4S3i3U
VOg8CYaFoSP8s1y50BAlLn4bXh/sXDRLzY84E45D1CZvanfIuYuVUMZBCsqScpjN
vjPArdz9snyskTi2mT2D2M8pNcYanNe/KJcmuN7NAUnfF232TxvLUEzxtMuWUzCy
NCCjExFH7GMsX6dlueS3AyCfliEXcdwhsIFc+POf+26aAirBKAMgYtZwXPtxgnrw
9dUO3VSj8q9/Hqg6LE4XT/B5IAr1w8X1TORsNkfAQP3/LEsRT16igoLzqkY2lEdT
SKI4Uts/hNmRebiKFlBqOF2SeaiKKbDIky68EJEogAMq+qWax+qb4WntlVtaJ4Wu
CYhz43A/tZCPRKP95C82y5qSIha/h6/O7iaFccJQ3QIJCKcWXHG9im12gt0iEkoC
0rmxKAB+CATKQFK4/KbMr1z0/qS/tnYyagA6F9uo/yLbYLVRWzqRjqknHtyRW9Ca
qX6GbjWgvCtX8f/9FzOvG6hK3VGHJYrdqdwgq+Wy/O7+6IZu9a+F/ctOB0v1+Dl8
Yr+rdTyN//C150igByz6zG85wDLGEI5y5fIRWrtfXqRjW3Vl/eDBDTHefESeJoYd
y+zJbSJMI0ELhIJbY7avRUIvLlh9u6TbfhCLjZL5hwPmhHAzgojp3x32UdME6gkt
/mRwzHa7AXjHFdJ5dx7ciYB+oO5XaFO+UWUL2im+pfpIzl58ybTCWSoa3luofvWY
Bm7I2XDEndjqJSbW8bKhDtQEx5GZwsBJja9jOjAlL9YuVfQdrmewgk5+KIhdk0G+
DFjFXiPiNSEUZPiu/QKwSN8TSULmC5MJ2nNLY/VlvZCvjI2gFwRRKNJUeI6YmWrg
hF56jrwQThlJPXNnYCimIseGrgcO+DeqExSVtGZ+EmabNBKKEFjmit0oKkqbKBNV
stsota6pVCJgwJzg9bG6F72klReRL8b/6rLd9fAB8AnQq+JLreNEGXu3OFBomLms
bdXZoYtSvBBBbqCxGr47McfM1ETS/T3oOZ6iENsvh1p18AYf/kvo+MNhTw4/0epv
+U6Jxh1KN2EokW9xmWgLIFAJewMr7fUS2cdRoLgcLRsGlR0TJHMyMgmueF1m6RP7
/UpZlKj+wuMLk+zg+o00znJ+uZlBs57BBBe9Ky2+09bP4rNqC9epDgp1AIpegP7Y
ykspfZkF6MRzSbt7vp49Deq6Xr3MehLKtLv5F3NDZ+RIXpG9nakuF+QdV+CaKceB
ECEI/bFKqVPCxOw+f2lxCKvxehCpXwNtlE3lx2wpLiQjsaXxLY+0YfKlA6FhlRt0
dC8JuVJdvmWzbIrJD1cJLeZMJ11kRGaV4nCozArke2Sxd5UkveTMgS2SgvNtljt0
6XtasZPec5W4e2RG2uvRb2pOcPsKP5b2GsiqyG5VQfmlpsABDdHqryfOWmI41Ok+
8b9dkptkt8fK3XB12s0a+ggNVVxsFhgGpR6GRQ5PVnGgefOQXzK4GPwJ3ZgZJLjI
XUYqbLf7jSaB/XiyDI4N1kJKEm7DBKQ/U8z7OoqD4uZzDmyXXLGaQAi+Yon807Y3
sJdaF1WAYw3EAzdsQGderOvdD2CUMLeziRUTgauyE3MefgMmBvsPOeBoPB2Twmd7
jXFuuhITvc7cGTihwWbfv2O5PNm1/fnJe5EZDWoy2ZuTfx7xJ8PsUSR2rLeXZIt2
Je+7psQQCcfvleZvEWzX0Q7Nqgoiy+QJCaq79sOjNkwwrNqJ/itcl/awSKfk5d18
PMM1m9CvALt2vPYeIA8k+uI4FkAI/tpduaQvVavyGbQB43RfOn33/1kGIsDSTN7/
aX3SaIL/OBa9JCsQZVRPlOjsuKORXdB3Q3ewb2tQ+kgQPB8Hdvnmw9pqjX31qD2n
c6XkJZhNl5dM+UR7lYYkgyOaHKaTo55nNm2RuYfg/trxLRyHc7MQXnXS9OpCO5EM
Goo8Gc9CxLt7m2UbLnORRj05rnj7lgMVfh0muQCtQMOJvFDrkTx+Ou+iCHzC8aUR
YEMGH3FjYW7QXtGIMiAT5up21rTSLLQOgsknHfwoklReqWRURDYJCnMNZyia4dq5
RSWL7rAfoNJwZzT/kjowlw1lPoQ04Wv7yO9KuJIQP8VtNv1Mpn+R+5SlwcqkAd/X
mkQWkOxNiwUSKtUEOhExHTEQy5E+dwLh4b4M0LOjoNvxfsRUAqYyToGlUzPJ57Ea
hQGVHJ1KxLnoJNjf1/6SC5MykZzfxPT9ktzGv3z5oy7sbd0rQC8BtP9JZOP97WkN
R6VciIZ2saWQTdWFtWddNIy9XU2qfNCiC7SAfkwO8FWOlTxGszD41w9nUZggqs1W
mEXlMMTnDTQ6eip5syorWMqNcBOT1bVJg39X/xUB35hFCaVnEiOldSOESGnUMX8q
thA8dayrimyO/cPYGJCEPD/5hJZP4B/Z6DFnlytX2xMAlhsGJRghdIFTixIKqE9b
LIO3HUQHbN/L+xANEhoIh5JlJjnFWoKGH5n0fp8QH2cbE3rScNW8InYV1ePth0aE
OLr9ZD+YQoRrZ5MhTPLyZl3CpYglZfS+TeqwuJlt20iMwqPngzDu+qLWIk+k9sfa
Y86fY1SKfuwy4MwPu6oLqJtyRMc64BgO/VGcHEOzClMg3ySj33Pu4LrkZA9EYyJ5
Xdl23i7OGMHiFPnLbB8kHP5b9apnfEhnHBerNwqrZpfI3eJNoJE513NOpE/n0P/A
NlJ7VzQnAr5gwkYpwi++WCuzD4SHzZJDCV/zD9gLoEskBw3EiGhYZ5r4wq8Wj25Y
Y1etHwIM3rRa5dyJyqs+siMI60aAziSjoo2Goa6WojYxKfSF2KAD9EReVUiASJCH
T8s0DxgUdMvLVdmsKA9ULEBvR3og9IXlBKZsUqIiwdChEcI24q0og0/LlSO198WQ
b59x56kIBgij0f9QjieDKjhBqsaty00unlgak4PyuGxUBoJ8EvLFoqO4CpjNiYdA
b6SRO0lveNAjgzvhxwRutUTq/s+NycZCVza+dhfhI61W9SEySWB1ZbP6impVTyfp
uSAcFFdDA0YgCdiSFGRUuUdUyEoPqk5crtJNgZ4jw3bi+g9X6bm/oErU0XauiTFl
5wj1/YWKKDDrk0GBcg1lJEXbLiI8jk3+TrXh27WaebkNgHrj8HIaoXiNjoWRqNXu
xtFxNz4AHvl9hVR2hnGZMAfFstINf4GqybpiSxHunqcu/a8NgXxn727SILSks7K2
+c23EyUGKDETMjsNj8II5QmpUf+kWuFqdpBMJP5X2yQ7JKOxjG4t1DQY3xcMELJg
4R9DZPvKMsHrCQCH1Bx252ko2gY487Rp/ZwBh/k0mbVkfOlufe5WfH2TorAC5Esw
Hm5J9qVKncp3ghRI8JVq354IXixBcchejfPuXZzx2Ub+fYji8lcw7gN3PPNllm/P
U1vYSHxfGCaH4Wxukoa8Rko3/1W8bgvch6L0pFltiXS7yMgZyhYAI+xC8SOu/Q+q
7aJEFFg1nkFOK8y5E+ozV8qpdSDIuKIRIA5sep5AQXdI5ctPRQjFXMkPdmpQaLIW
P1UJ/79Xgcouvw2p7RCWA6mNJVEnFwBiVo4kWi+9n82DaMPkFyvnWgYXZtgxNNnh
LeQHtAwUOEMLGtm4r/vXzqEcWGVG9ZTfCcJTqkWOzWu6yGrFi9JojtuGO3kOrWFX
H25V/QIDDd46bn/JeTIgyRDHa+vqaIXnc9TDGitns8WBTPFPY00XVW2sFzL1jS5L
1+3MpzAnFJfVXcewjBEBP813J84kZDILvMZh+TWXn4itnoFueOcpG42LItRa3NOj
eGceLqfhXwqXjsqF981ZohHZZuGK7JToBd5/VnJfxg1D7ExoZcYIkSA/VSB4Oz+L
xQMt4SFTWH9XWmW8GRxxyzV/pZVWyOUs+dc4En9ms1WQ6RWB9pCu1Lfcb9KmyCc9
ppTVqf8yyfUZ9lbzYUPUQN/Svyzm/ig7b/36QpOZF5dF4WW8XsWHrSe/PWS2WoiU
27n8Hqrzfxj1zEtO5NQXLWexKZXdwgcSrItGgRQfMaQhniyjy737Rw9W0SwtZlBe
5FcnIUsnvrTDg+IEQT+BqzBjA0rz0cGrufomJZ0LWdWr4Up4b41QNPR+oZgQqLY5
w/PduWE7FtPZG+tPUbrCcyErADKdhsLtSwpZURCB52xFeRLgR56hbM6xrO/LJueB
CfgkFrGwra8QhMUr76bUaaKNPLV5EkC3QQh4+G1yQkl+inffR1fg/nBEMchAcISv
11gaEZ1+H3GRX8P/ZJL5Xb3P8Rkr5rHT95qyArNNMKfp/yjIjGvDmhilgydZEHTF
vnaz9REfEpmBk+dw+QDaQl3g33BfrrZPT75sFoWpSRp58PAYVjGWUyAfr77Hf1wU
/8mPzEl/IwWHp0DD3Ms1yJsye/5qefuIrQHl0vLaSdb8C2X7y9JLXw9rU7+AjmEl
+aFn1WGI9tS4aXGyMvkc+UV+0Bakm+WJIF9yb+kovVuxkBt8HYX00tlczYOtfyNt
M0gX9hBRQAPF/hJy4MF+O41C8S1cwB9/yvLkKamZVDFlxp3dmCc5jdv/UrEoRank
phF9qdB3LYq1vBbXalEqUEn74MUEsP+L5poGQ/pVwMo1QaBdpCcc5MywErEHCDUT
dsGamTErOM4PYbsDLtaiguGSxBE/+HMB07vx6LJ2U9A5LtSMvLZA20uypYqtQsp+
ZqNCCCbhVGyx87/O9/t4F+TMz9sToTQnCeI4ni3AyIsbGa2Rb7NzJ+Gn2Auqok5x
kB8z3TzxDt/64iDbOlM2MgksehPqybPYo9hrBAA1QA8Gi1QNY+kTsv1qPrvAMsnx
s0LyLmO+zQDq2DU06+Ax6givwQyqXhM+my4joiLG597h0a0Qnfpd6i6pWy384UmV
Md4wXQbFOn5pCaqTEp4lhO9Aa5Z9YXtEoPIXAZ2FfZ/B02gP0flou870tnxpFCfN
W2zM/i7cINLIgOqHkcxpoVpdoPILc7yLkVgbVYsiB0lcUJ87G7vv65LlFQiNBGUZ
+a7SMif0cWb2LiVRQUbV2n+uFfClfZ233pF+YG5eCPWMa1kiEqq2kNPxsuL4hCsz
//eQnexTRmMC930aSjtqhkkvbKLMYfD3PzyuyfjCir2qj/ozAihq7fd8Tk+Cw6P7
rIgqRApoub1WhoRE2A7EZfsxmXgkhT9mnIwGwTITny01EGgzn0G89ZbtMi+U6UVf
/jjzGAXO2Te6IG2l9gsVBk+pYN/6dJaY+iE12aYJRuQco1GbxGFTAt8VrZh7/OG7
Z3G/ikDnBYIG/bVgyXHUGtYbKPW9mOI0LeKceFJQkBp+iHR3RnF2rCYOTe8dv4a1
VIUYorwngRffCVY0YLPHRyIzmRFCXrfBYi8wNMnf+XPmWqp8Q4hyx2PoBZz/JBag
+IyHrbqB0eKKEqNzlMMC5ueV/0Zh/t7iLGzj4anog2esUELdSPdM6Kk3SQallLrc
dxcbS2gpTBlUBsqZHUT0Yd1DecAwPhO4rimowlIu5SUiflqBbjsxzMAAxNcXHEku
Hilv8ZZpeH9dFxvUVSeK5bwbpGqgAx1pkRRrEe85OUwhqdYnV2D0WbhPbCbcE4BY
3iQzwDhq/mtxwyz8SW5HjBEijuJqlsm2MCOfjOKvjRGRuTQhKkH0DJY3f5iQGUOw
pVrESGz9Z0ZNBIKUFyi6etKsDOx6w4xcj/cq6yePKKzXhY4TkTEaTZqnFwb90MUV
wHKaJ7DTqx9uxPHuIWm86MkStLmqF36FKxzvZuEg9/wugsr9e4b3QEvLTmrw89AU
S8hitXUAKTPec+jfZMguxX61RfnSGPeDgaDbuCEGLHU31XbnzVNRpHa6YkIxuRrp
4vJMuqcOBGL7JGHN6g0YXQxJOjGpqNviRex59bOJoLSB+OMX6XdgVjJxvc3HJ/hy
v/ifiDpU2Cx64Fy2T1Ik36U/wSeIeoxM7zPbZDFL9MOUN3tTCGFvPTSG2fMzCwMh
2W1vJ/0CIsMTwoBiYfZrTgR42257hi1W8E36g5zmOOWKylz0RvlbH3IA2K2QVdDq
JCsMEORltVptlOQBqgPIxWBlLiX3D7/f/1/WNAgDYrDkDshucgHJYu73Ef2LFf1n
WcPzSGhg5a/LeQ+v+eHEOsS8M4nCd5YW3cyUX8lJw9rl3pVEUccWNf5QcG14IfNN
gFosJY5wozM074K3enrGHN0BczVLXhzsySJE3daKUHvys1Qhmt8WWQhg19yMV67q
jQVPYHvBcyXymmapYbQzWgEJ75RGZYCUTwgmEOI9BoB7x1yET1wYlodgHHr/aWat
sN0vaJ5aZsBmln7XPcSKAdVDIJcsq5iIPUZ2JcaH7Iut+JSxufT9tW2f1oL1XSc+
AeeQgK6xyA1mvOdPPCjWEIZFJ3hLe3JB/SEQ0/I9tch8Sg2rVmFrYTUMgXdf+QFG
8xbzYQcwMxY3betcXNRI3b1qEKHRm8BrTEy30OApEU3ILwj/4tbX+1lz/cdjpW3o
pTS85ZS9WqQKwuzv8wGw4f9a2RLT6PLPAvLCVGF5Y7Kordp8cnmHh++XUP62fFf/
Bo18UYqZ09+3CzyBbyhqBjETyQ7vcl/yb/O0GhNps/SOnEigi/Y6NlPkh6xvsURZ
cIula5ISqonntRnDUYErb15gPzKTI+VnUQA47IhMuoCf2HEWqRnqFOpiVkrL10JG
M0YtP+Se4FJs8zZbU7SK6FbqHRFXI+uCmdPfvZRmD59wC6BNzYpMmKpDgfwRyrmR
3D7xvCTR+fN7j1P4o22tgIL1CtkYpxI4kzIF/mJgy0KoKa2NxrQgIpJpDvrEJHIn
zzhGRsBW2OAvOukVAnQZ8Y00UykQIaler1XtomGEHvVcHqw5RF3co5XSdA4sNfsw
r8fz3f3xCdKNv/L/EW8CKDOQE0owS9RWvVeEgaGeWXULYlRZQxnfwk4EXriEMS4+
f/cr/zWoBut59a5MlLSMcLz53HGdPnC1Z6wrcAfjq3HSoTeCYTFZNJ4VWv7+8DWg
cOH/WWebqBsm0swql1I39hOn4ldJ8HSgegsad6QpkB8mTyzHJdFwFsngHHEQOKk4
mXd9VTkwDIdCWzNflwxDugi8oKnk3h/AGmw0/m4/K8IpWvyG9eRToGMTb5aOK2fg
x8VjHp47FPQSaWsvc+dHX3Ri6zLuQYryKkElssXWvu5R3N+tf7GMJSmC6uYup9XK
BbO0uhDXEB1fpB1a3rGnwddS4N0aTQ43HBLnoj+2LG1kv6huRZRT+o1DGCIDLenC
oNJivY7b8vWsUh1uuY3Mr2k2tBSx3aMvupPfSMN9u/iUmbzU+SzYkLSxnu1pcz3z
/d2sQv2SHDeJxhXsUrAUTUIVVbFBOHxDNGksjogoSDpiR0fqEkSnFC1fiJDN6fqM
BvbGfSRuITd2esmMj+f0PgT/kYQBIjVc5l01oy+q5V+fO9a5lvaJcDdRzE6zU3p3
rKzefQR+JfdgZyid5k/w0/lsI0tneiDymeSVN40J8bhuNxuTyASIQiSm91iqdCzN
7zzrSkjnzAM+F4x/Qx1UHOhN6QAMBVry+jB6IawQOYZpYoaTlcqUx3KPqNoigiEY
wvgWTn/XLQ28GaDwjyCVjmUZoBGpj1RULMaH8ce+dmeAS0tK7BZ4GrwGmCwhHQCa
NjnyiWfLszhtLIKRx4XdoZ4Z3MmbxaxtZ4r6IpZg3mcFvprLiaaUXQzqbvWGeEEt
43hT3np0aCT5DOiXnbjaoZktloGUPXDz8kKd7GMt0DWwkI9Uzityvt61Rwt+dK+v
uB347lCzPWR1o5cdegYOuGDZQDwInSe2YeCaeiplxuj6qg3UzeJMwG5NVEPiLwfw
etU9cPtFUcR2JycnkK/8btN4gz9qQs5O1jtndjFyhkd4M3CfmD3qCcdIU4eYKffC
AyPVVqqn1z7eUyNj9mbLQJ4TtcWdZkf7ZO0SS9cZBsue483kALt7RKdSKB9PudlT
YuifbmFzDnU+7zMFAAbQal/3zwmEI4nZCQ1InI8O/K0PTnT3SYU6+1HdgqPHLIn0
yOn8hH1nUpV31Sa5G87YnRbexnCgKaNTJEILMK9MP/Z8SqZayv8QFdLIIHDYrUwF
DXvwek6QymOXUavxtBVpCeOfjEaIOXqXIUQ0ChzoE1/mWT/FkOSjS8a/gwkWBHkZ
/ZdF3AX90/AN4ZRZk1BhsMeC4M23d+IiBDMM7Y/yGWpsKL6btpjeatZst0IAcMDR
8bLpEUlNaNJX67lNQncVM1GZKf76WaXuTyrSyUXBBo29rRRlXEv7fMJSHBYJ1qVA
MAZ8Jy8tnwzLStgUlcWZM9LFRm7zh4GVwiMHjQJFCHr9iWasFUowY55daTuMWsTh
D0rIbur5si6eVlHoAOR+Qg4UKetvCyiaCb+x42XC8Ini64vAoYVM+k8pi1tbXRBw
bAz1EcgzR5iY4euDOcX17ynKPAMyx8QhKNeo5YXnrwFrXkqCcEyRb5B4dwNz+Asa
SJ8kwuRTJeCIvaJWbxaqg27NTpI+qvQjAZ79t21MQuCieb+/8oIBrcuElFH8zPC+
5016O/Xax60IpeN95x4qCLdr7zfwmSZOkYq8FyRW0r6u15wwn61gMKYCFjEcLsLN
PvkEBileIFyAW1WloNRfefEph6ayqhZncEMOHxw1vzAyMItvYwjXZvYwmmiocgbM
5nRROUcYjG+JWUKGEeUmTuyL2QRESkzZHFew72fTG+txoKgMteF/Bs7q2L18aqzf
F++Zzd90IyMYbsSz5i29hroq/EtRmXzFmNUCBG9KESA34N5NdTEUxAhPXh9je4iJ
uPdC7N53aWJ38N+1JnjjYIafo1B620mdRzF8EYzWw++iBB7usdPqIi0eSRswBUVU
KBPdCsYXbIG+YT1028oPOFGW+nUPgC9yCHj47UPr9SuIdvpQF9sRHgtWDUTjQfH7
01FssicgVJmhKzPg8vTSIMPcrN/Z1Xnxe7VCvoFA0wDxDNO50cizwkaOsJlsKWWI
/1bcUIAO4rjCSCnbLY3G2RbcXxB5Qo82WPPg8yxtodN94UzqEDJMEnvIVke3syu+
JKZ+7DxDlT4jCy7/A41js2kp7lQjI6cEAumdI1BLI8Pt/ZHuSlZVbOEjL7AHAaGc
h0+FrEA+qSsO2QRbmDeG7+Ftelocl6PeXz9n4IEeH88JVAvZ8G4jb2dDibe2s+bn
Kbdphozf7pdQppUHT7NjRqawFJNRDulPXBa+bdur6Ye0ykOKWc1b91WPdWEvOLsa
6Otu4SB/gBMC8nPo1K5JoKjY1CYsDfVfgovXIGJpKIdjn4Zcv3IXmnqDbVg0Xmd+
FVY9UnwuQkxX0r693zraePcrhLAF/IhOD0osvHK4IkWHQsT2PjKXCo0cJJlKC0wL
kFm3/qE+kY4q3v7EKM2Z45UZEnCfre08wjDeH8lFMR9g03/mMwna4Gku2uFofVF3
sXyB2xde3CTV4nMnFxREundEroZC+/LOkBDytBaxmYyBEtgJEltanG2siSZS2fKw
rvaE663EWcECKghW0x+h+IkEbsentfkUr7gXuwvFiZgTA8y+dTj0WkB4RjeZ6myW
Ana5Y1QVCoO/c3ML7p1ZkVAODJGycaQ2n/PQWM7k2R2T2FoIw/0r4/qny6vhEKTl
Kj/0PzYCVJLVsabeqzJbVhuPsQO1IzKfkxiolHa8U+sFksrmp4LWcUQi/KIclSbM
tDD+BEmtq8t6Xd79aYuMqyW0MZkcDyb6F/i/3SdMfP4CdhmPl2gj2wrG1NlpS30X
6Bd57n+dYdFutD9Jyo9CHUPvj++aAwux74CjH9etBtV/lnDJYwzR41iw/ryykB1D
KzQBzYFiyEHmXQcN3dPxVrQ3v+q39FEzIA48GPtg6F941CyyfPReo8Ndt3pUA6Mo
4q2qsMmdjwMV3RFPAJKc9wnBiy80hgt28WI9niFkZNhl9vsGzDFUYLJscXGXhx9k
0IcGY5blx8V6lY4Fk0KSRFscpNcej68jvNb5GEJoKlASCwwGMswQ0mm5AAmIRKVe
QAUstAvkD6puB9woGQjwhD9T01omIbBtwWSfzQ5r917bNfmcMlj4+0MihdOa87VF
UuxLRxzyAtohbxe4iphp/Sx9ZjtaGxL9X3kgUYiIis0/Ow+HBimUkFGkUoHXauQw
31r6z/NGtlvctueXRrLkU7H+7ITmsc61sleDRXD2yxoecuVDlCWiAc/77qTBoIy+
bnSTEWTFGxlnYt4o2ZIF3r5NcJH5CUCxtWlR+4ZFIxJJrop8AVWjEJqixUHjC6id
psBZC/QcYSn7XHBsbWtjNcpz7fR89eVuapGVo/tobR+7swPRIo7Goq5r1DaFOWZP
vTB7W7+MLgIUWBbNRAMZ1Ix422MnBoQUzRcF8TnZl+fn7j4FQMxJb3k0xWye6F/w
D3g/9q5+q1u6owuSjdXjR+4l7k+kfcLM+2RJHEysUVQCBCC6L1no9Voxx34bUhWF
Lbng4WHkeG8PKumtsmWVlXDYzY0XkD/cqEHyDW8GbCQNMBV+dZ2Q/aZeLlsjG/rW
Hj1cXTfLKx1lVDZEzpw+I3Wtq1FWlSA5mKErEf6vUX+K7kRd/zn9hR8F2ZmMC+W2
b0faaLZtGVx9jYbiuTSUwL+Swe4HB/LKmqpS7yWpnSiYTglzpORaWw2zNNiOzGZ2
gB4JzQdMsv3keMSSfPgca5mnYoF0hEjNI0Y2YUxHXyJjjMtHcfPPX/UsRgLOtu3g
ImzEz6+Ns9sahokxBE4JOxvTTS4gsn+Ew9rB2XXyVEJZ1O93B5SVnShd+6J0ypNe
vcHVC6f9AOHkhHIWWv0DI1jM7Xo3QPD/rFx9TadGPsvFRRVDTHSC2iAi6Jwn6LWU
rCPDI0DnTZkhGUSo1ae/ZZUvn25vWWMGinJJWRkohYte7p2h3ZfUylY43WZy2E/9
FJ3hKlxcHlX1ulSFynvVvWf4OqwcX2IZtqdlbYaCntRfKWacytQMy2ND8SApuFzH
m8n+YnXrjd6HBZl+3TPoVMV+zO8Twundrao/VBXu3MmU+NjAMU54+Rj7qYRPhecM
IbYMPo7fvttvfTcjRIjOhnWqYGThhbtucCdnltrOOfmRrd7HZaqjbw2di/ShrlL5
Kja0Cdun/IRVMyX4kRD9nYMCKJP8fHUdaco4v3C1pIufs4Nx64cv30+ge96MOV4Z
F57kmiqrgkdlfkURueMfHkNZiFiAFacHX4mgmXx/xwYw72eGqrVDTlsSsq5tJiNZ
jXtYCFCe9PMgC+HWPJEbcWS3W7On4tzowA4LgStXYnMPb056JMalYzB7EcSui0PM
04NXinoeEscLPR1wiDW7Q84iaihTsakLYCvpavK4FAbI4BBoKskoctElvq6QGClI
nM25g4+PiyM2ThJigqkccX2yIcMWfq13F5nu4B0Lk/j8mwPR9l/2/0NZlk+VVILt
dOdvZegEDPrwq9Kgn17zeY2uEwbZg1HrMdn4VMr3L7zcFMDUMD4LvMHH03vTQTXM
Ts+ziCJl8w7IZwf03E9CgES0F9suLa5AiVklJ1lA2YKZJHpUP9jmMDODPdcLV3I/
hZoyiq1Vn9Zk6+uaSK68xONrH8DlpaexR7B9nBN4/aNJ3EuKCzBR/gXa9wTs7nYp
R+TkE6VolCxBVpSHS1XBd7gSgJvReRUtErScmP7YbnUwnxgXClGw1hTbLIMyxzbi
Dv/VlUiDralcevS6bNVUlqnZSEV/JyOYqmvuJrx1otSH4V+URU3PCznNBB4rn59a
3onfaAFOz11S9GLH8pAyqxAGKsmY0Te5EpyKz8vst/ah/PGFuxBCcgrjzwuMkex3
tXdHCgXJk9+IZomtEWazzfR43YHBIQuUZaofkep9k0tG22vMGRae60ZXkePTmUvk
PELthVPI1j06znhLOWi1MX0DONaJ4Rg/SN2KnNrBlKSNBeslKaI3HlBobjDbH9yV
GuWU9DYUUfWiI6wczfX59HhlkwEIUzvNvAflFfCMcsOEtBVYMWi7Ctf+nnQhDKE3
Mqrq/t1yqlNfQD+APiZR+umbi8CbGE0D21/zKWEk41ODoBMxDAIlH9MdXlKjAyDC
xMcACDNmNcqxXrzpdacA79NPa+tBzyCobp+W5edPsv/V+xmKirm2KoTILi3Irkf4
I5bc1PMQ07fPScBFXTbtgFElF3SJjLeojgr6F6lh0RvHQGFKZncFISzG7wkgbR2m
YWa8HoE85MonIrUE34dLrW8jciEsJZFI9TjSmQO4lRKU9YDjILURs1W2pOOk7i99
jd0Gx7lOBxNb4NfLf1hkXtFpnQ/ANu44jPcovIfawbSS1HXSN6OLG9HHqz8gLZvV
sGJuCj6FWO2aZiQDLSyDpgq8v4ii2cqR6HrHcetHmA1dUDPu+r/RtEQf9F8imBLo
/eVFO1zy1SnoW2eow79vo6pXicIHYM29IWYvX94z6vNSdeaEToi4uW5E1mbn1BLZ
N3mcNndAHjEKyfJvkSqx7DwSTRirLiH6ye5MvYqe88CphbiU8CqanzhRz4UXGnlV
RMscjNsHL3pvqsHhtKtRkGC5+ixMyLUM3jnAc4svsLR6MLCK7QJvQwTo1Wxl6Eq0
NntMYvMB17GNy7aQMPO93mfTSyrgAO3qGijsaXWeEmXMiBTq4KU3Lu/zg0u96A9e
KR630a+pVsH3Fshn1i5iWqpztIavgKx1MJgJHibQRcKOrTGe9mqMDqF2K9Oq2pxK
m0syswQoJivd2hPe70rSjP4ehq8YWY9QPg+zT3momS+BrF86KLJqilW96tI6bBTQ
jVtz4CI7qntYRF7wzQTaUsOLC/pvZPCYHVRzBl11RqlNOJrkMxz3bEYV/vC7dtS6
+WB+Y/nY0YPtSETmtUFhe0bFqwl4/KJvu64sSV2CahHlmkSiluzwFHeQPdUL91wn
NwOH221MUBDroKbv+G3lqmWt43vtoEvOIWH9BsL1GKIABtcJ48zT5tmKJN1FlP1a
8BnYrziaGvZ0bGWbw2zkF2IF9o3ULet9ldt9I6p9121NwI3nD3yOQY8MTVtaj+Dm
R5tgLOUegovoA14eY58dCuGnyrx2vUNbuXvbwjPPQvBAzBumFbRoy7v6Dl/alI/S
uEyWB4kNqXotPkCHrXfmIkN/d6uD7pfHW763Q1cH6QO+6bOYFHPDjI8J1ksIj/qc
Dzm8oBQ4jBd7MJpb1njvY8VlrqUd/+0vO88Gb7x1AG26aEK1EfiKnYWKOnd2LdoA
jtUjo7GJkCVYIf+Ol3G4h6oX+R+AhyrDPg9qXBhLfoQ/4AjEZtx6MA28K9XaIT7o
mSNbaVRLu24rHztPdSDPwPlvYzAdaG+exoaItLSB6Ne/ifmdIEeD8l8t0hwRafTm
6AqC7WBM7zU235XQd1swC3BSlfdtEd8pQZMrwziDYggSA9KAnu+Y2NOGcfYRakaW
WFE8VV1xtEseAgnflaR8PJYV53UA2+nqlzerRaxZZw3ePNsoCWoB3auhljnyUGrL
mR6+OixA8aTrJNqO0HyDltkDiVc4123s+ge4nnHP1y/rjgH6Qdw6RAMVImqyVkRL
DY4hSXBcoxuo6al4gY6UyyAaC8oRDMSTjoYBb0juRT+/lpbkTGj8thgzJgAgY6mO
lmljvPLasyralHuLk6eFR1INuYtmCOLmA9gZeXOgfKr6Ns5fxxYbQfaqiVRAcwgi
sBHtOiEfqPTeXCnqs7xt8rAsF3OM2aIQjFD+wvVayqbghbtscuQkwCHKuOB+ERNW
Ei4B3mnQbv/wS/6ezBDGl8Y3jpfjpDbckS9ppHgbhvde2hXHLocyKdcjwny2zFQt
LKfGnnbaI0I8CQxgBINlaM3YbH25pmAaDzVRPZZdFkfXqC6YOZZDzcyVpWGATOMB
iGg1hSVfB5wQAcuH63EQJVI6yB5RUQHInssu4MTUGLD3+wWLv2aYU3JN4C9dd2+C
8npfExDrL44lBhANHCaAAyefny6ns1z+FPQ0aiy6M83VAHT0C4vyzHwakCaln4uH
hauFJhd+s4kU7fEYJ1Jon8cK28uEkCeg8nIhLzmhX1Xr0C0LTVBil0DoE+yDAxdB
y5zW6PdoHvwMNs5XMCkuTj17b2brMXqxH0YWQfo/AjzN6EDvCUDG4NopWGpPjgn/
IXK/ktu3J/sgSChT54WN8Xnlsdq2ZcBNRn10GswuwaOyO0coAA6zgur6ofTueph0
MHsUVFGxvOGVZSiW9W9/oD8RUiYI27cLm98AA+CES9BrIJp35+OjDgmEhaCOQITt
5cTaNyqmhrAepMeBtUw4CQWhsP3OFGMr9FI0tIyNn45Y48kY9s53lqFJvA+PfLqw
6fVR+bz4hIIeulRwzN+p4YzJtn/SU+Igpasu/WwyiQ+0ncCOYiWJy7UTAEkE3SY4
kla7YKwII0BL9qbOR+/LLhMbvy4t1QD3Z22TnDBdmac4rtZcNHmr/PRgLWNXpp6+
hFtqCsbAw9Gv7HSIKMoWGgg8bNsm91yGzr3SEgfgxREeYuvZouSDKjCUOp1LOT8S
zSe2KRPZZAWEQYuz8yvXF8EKkxFgVmumYeji6+QwBdNcps+PGfrLzG9dqJufxGs6
+i/TQdI8KV4yiZlLRNcWkES95eG1csjp/35bSJE+38lmhDtdQwQY36cFQXiw/byM
G4ztBPyT6ncP3rSeDf/fdwB49QZZnYuctf72v2BKSpC7ecpU1+kXEDLqYlm2QPN3
H82Gb4/fJ2CW4xY0cYaGr48PHqGPLP0kavSmWtMYXEDOa2U1SlmdPd9sZFCLfqYg
OlrpHDurmAjjuJF93kuEYxS3rxdXyRogibw8fRxruQkL0qaW0o2s1wssxYE36hZL
J4Cm+a/fXynAwySUfeUoSJ6d7EukllASamPDrc3QiSqSjplKpLccGZUIeoHsB699
fe8xK/CniOGjtmUyq13liglhHcig1/jCnskQmF4rgTzqwPRDDZwIm9kPjY5kgJrB
/HWIBYlU8gwQNkECz7H4cp9gQUNkzXNDwAuSA2xqJJRDpcnKVKKfBbMS5lK+Ih87
yOTeJ3EGLNFSU1pI2IEl56IJFXtxrYHeagGJWxiP9k5TmI2wa9WlOvtU94Bioyqy
fL69fwAB3EagQIvgoOuUJQnFzBebMrL4zJfyoc9uXiaqR5tmd79fYwCfG1Ivqxwb
M85ac0TJm+kaukKF25cWKsx+LQV0IbIpxsjztfxyxbOiD7WbMwI9EKbxzG/pJXQG
QmCpOf4w9bN5lCAnVhf6XGO/lyy/UdBYv1C42Emmw2z/Jgejw6GF1LEcZL7/ZHOk
B9GkDyFKfGbjc9TT9gucNlNB8Yc5qnAHxdQN5CPfN2JCfzE21kN7023C+xZNrzBg
R5PRjY+wk3hfMIYIHVrxE3ulpnWZLvmItChT+IoWihwniZJhE5bVViXTHuosvje2
rSWs+4P34hWBe7cTl5qhkNpD1mjfy/p/h5roSkYfX+wJi8QcWqIXHrTKMbK0jWQC
gF/dFQztCjTruwoQpQUstkTMuNxQ2GGvmJLGga4z/eiaqMMuPB72xJCL/pZmXOli
EYeMMnYVSre5KLBShc8IeI06QVTRQjAuPQDkE9wNyAFApgYZDE8N9o7v/Fjf1qaY
xq17GbkhBY2qlzV3loFncrYMF9POszGWWQtVYAMn3EMmvDhh7u5kMrWG6cM/HF1t
NtM4SJbpWQUEkw+d2KuZ45DmqGrsQigNkbVGrAYtnWY4llmU25EW3CgO85xYVcN/
1ZWS+Wj6AwdnX7GPSa6bdqKP/SDdbsi/mkhfSoemKCWBTXiE6l1zTmafYr76whTH
3J1s6fXvtN59Jg/yjnzy5ukB1ReWMWQzhbSmsw7D1IJMA3K7AV2FGi7R/c60GHXK
TzIuSbfglrxmN667V/SV1MqQ12qV8Ms6NMdjO97p80SoRwnuuIRCPbQiYvP7Qklx
kV7WmUE2m76+ePi1H4SHH0zXEzknydP5gVtc+C700cIT0gelEz+ZXidSTe3+lnil
QGC1z59DRLYSR7EaqocSZvSBUBlLP2G4X7294ZhLbWK7NI1IXtU7xhHJ0hiwW1vI
98qR/G49LyU8JDHwbONfow89rxzXYOjUh5AgaOCcwI3sblMHZ2+ueKXM1KhxxZY0
vi1jjB4qvhDsAwdoLoUUaeTLd0wg3bosLEgdMjacMF5XsS045lLBgKGIIPjOALD6
m9tkAquUgpIJRCmaAyUosPnuOgy0+Rlk/vlgDNTUImxwA8NlFEJBNC86xO1CXtcD
E67cXr3jnZz2JAPxB2PLsHU5Thdi+04PDZDksYqBGiPSpxhHPR1dWdik3QYrR1WU
YqQYY/fNT/d8k6eNADQ7QGUql8IaMArnVQfOHp/OfXqeCMW0YD8v3YiTuK8eN5ll
yjqot2dan9QnwG5ddu/1bPWeCe4Kag0QqwbnqZCpmAAUBF9I45jwlxkoEJN80uET
BTcQJwq8v4ZkOZXoAY+G53f4JA1WqpKeHpjC0MDSfYZSuz35qkePdrZbAqZLi4W8
IIQXpzduKS+gZ6Go13NuTDbnBRmFMn0TGm9/5xr+ppioOKvpBxyGtf8Vu8KYMbRU
on3hKA6fNfmx2V0AbR8wyvONhkR9t04s448k4ohoQPeogNLltMDpmoudI+E9OFLS
ARRkLlrCMwLQWXgJsdmAUP5HBfbjif0aOsGx/7KnxBJSAjNRfrDQ+n9O0WDsDM+L
E6h9+3Y2xMZPOpUtpHtyrSkVLRuhcaJnoyjsH3/a8bdK4CBjCFru5HGx+USAKdWe
1tLOvuvrWLHwy9X+2Pz5VStRME9nr8BTbG5/RB7/K1Jlc7XoTzs/9f7v6BKisXQv
m2oxKawVOnYPoaPYt17klEXyKtAlJlWALNeu2NfNyKgkhZchR2sX7tkd+bmuudej
X3LGAI4Nb11/gPhH85GMuUPVJOXosbumUY6bgiv/8+so6+KmSCyZJgBiOV1ILE1b
G8swiX8fS8ikaCiRu/humPD7wCZ2KTmTKIh0hJub56uB+VUVmzlLM7nI6DiXqDHh
dGrO8ev7uGNdqDCTHOdQtrMHO//EsQfhPIjWoTp1v7OkGTmVwlxc65FW3JKJx8Np
idWXNHBEn1tvmnz9ocdWk9A/f1K5yIW/Gt3fX4O1/OQHS8rQeJiYsd662njtnViz
uJJx97uExIJSQFgrMCLdBk9bF9lEMndbUkSvp0BkSrgVs7iLp7Ur9QMf7BBNK9gc
lQyP3tkTIvH6HreVubb5E+xSez9tIBQkPYR17eAXuiZocoQWM1+f6lKmpJuNyN1E
IEvYi07oStLMp5XpTyPvVPD3Se3XyXRMLQCwWIx2sWWJ+FPc8GFaquWf2/nOnVXX
SOzesMi7wm2vxkqwswTmV/qeKg534Zat+wDhUZxPOo1/vuctl7NDPeH/PXPyKKfg
/loCOxjWY7R/917D2ijB95/cEqVuTwgDcOCCdogrI0vlYyUq74mQWLzLifBxVxhS
EAdWPlWGpcbL8R/mjlJuYESFfX9pH//BZ6BpeobCA2WLy7MxInJv7ie0fRzWwena
OhZIF47LS0vmweercE6oRMY+NOERL5ZyxuO1+Rlsgt82KyDxpTf2DIvsP6F+PC0I
MAfmDlgojHdOTWnQj+1klrl1GpkOiEKi4+kasySgRfOdXb/DC5sF900OlnlS++K1
85zpmz4sYLD1vHL8ADD+D93nFFcTZNXSGS7oBdEt5XiGLcwlwVAGu9ktHIrAiiZP
kcH5omTt1GJZtH9Zhe2wnuklaRiyR3YdrlQAVQmoFl+K8C0zreL30tIiInpRYVHK
v+kkWB88D42K61qB9VwTRyOsRRR3cWch2R+ccI0LjPcUx+nJP7No4eFiAURqsxW7
jvPm1alOWxdjMpt1kK9D97Wi1ug3NH/Qeb/lbY8trUPg3qs2lnB9TuUm4CRJukGL
Qr0J7BM1jvz4q3C/Z1Et0gt4Lk1+0NyHk8B7eBf2N2r7//NMhtQZ+IaG8RskQ5TJ
Kn0W6du3272B9PvhacTin4zGEm6kBW71gLvjrSV4LrYq+DHuzioe3LGBLAnpsmRG
FXiouEq8AcGRQ7CAEuYyjnIxFb+rJOxVIP8xB+7wXb6M4oNnktIWVLgdxUILD00v
WmQmF7Ox938RmWNZ8OjdbzID7zubsNcrDJ80b6R9SM0bIDFyBQIyJiCdbpNLGYpw
w4Lc2ltrslWxSBs5xPkLXPr2dJ+Ab/cU7mpLlMxt6p7CS9O5voNRgc1bpL5zkl7L
gr21K4x3Swb9jf2AQQewFRceCTNHHQ86vmRzBK+1jGnuklS6KQ8vUiW78lf4WWq+
BwaIVjQIhlqmz+ZCdoDHfEM6MTWPsslGLyfitm7pSFgIKfmUKi2zPJwhwrD9Lp8k
3ywI0SSf/ISpPiS40Kcqu6u4JoYvgtEL0QIcl+V1TragmVm/bDRw67x3KfI8Z2Ld
LdcAly5daL7Y+a+HYJJUEO1M+oOyBKuM8ga+34Z35C+Eq6K3afTtD1zGLuNdYJbq
deGoSSDcDwPTnDcBk9YYLug+ZkY/dHz4oxaXvLhPzIA5jFyqTQhQ/Yg3U3g6UQyd
zE8YQvbGQkVNvjXr0KfLPZ790ZlGjQJJJItOCfaM+Pq7/jM+IyEXio8XQeCNkF3I
JUyg/qIatP80gFG9tJ5/j0slJnYaYJQAbqYVNsUPJE5I80KmXZ/2N9Yed8mQqZE7
fND06t5eO1GXDxy+WLEsHMcMz9UzEPv8N5ifJG7bgz6mpkWKq1Lb10cvOsZUkyVu
9uD4VuZqFHisJGDVx6GFKP3yUun+ZiwXpBvGpQEBO/ZCX5747bL9yLkVslf7suCt
/VeGVKd/OEmN73TyXRAmx+67H2lKt3H3SUX88Mdgeq2C0hoe8Af4/pkqR0GsDw9T
cGDILa2oNBxZ0H7Q+Z0rsHrgnTQkqXU4xDaryZdWCuJ3HL2r2m0vLX5sLD/26i35
yUvd/KBawftOCtHTmKxMP65n6wz07q30RKA4uvh0gBBKY1qyxXiFmdG+bXI8NGEr
I6Ht5/XRUF6IWBivRRQzwFAMxES7OdYUwB69APezNFOWDSP9EpQ0RrnsoLOiTIF8
8BdCZqrQLx3r8yEDGJoIliMTI9tEk+47/gzz1X04tDrDN2DGQ+qV3SEaCwcLZI8+
frIiG4U8wWtWdgokyVZJrzmtJq3dax9MF7Dz1oe85pXY7X8oqYP5TX8B8bqr0exc
PyJom+giklZHD8+E9T2oTJtfpRo5XKUdYR88yG0iaqFLCWvyfm8wm/SA1Sf3XFIZ
FEWsSCY/3OMNjUZBJabytUo1qOFTnEE+NO13zGN52nQgPjvsyc5hkPcXjVZKCwBt
GjRdv1nJFOg5gSQyXOocNl7MRhdejCOuhZmpKx7kl1/ugoW0gDdF7e9Z/fNCt18F
7bDS3WqMVPhMD+O9k2776P1u7TSCSvPZz27zwzt1u9xyTvxDghQPUGCzrSLr/0Oi
NgbS0yZXdoyqsQvqdVbcfbtsyBl1veGOLOJfjOMFc8ETojTgDVGFKsliUVAlCfkm
np+e6VC/9OU9LgiipFdeUHYzeXdUlYAu4U6GVu74lrJbbwYS46MfMHbeaSVoDnsV
kLfwchcRHkxmEgRP6I01u9CxwHLzc33U4lqVVUuRqPoF3uiZyFkkjZ/bnGeHo4A7
eGOG9q7KE/VpB8M8HxrHSFW7LXWj4bhqyUSTXBfU0aam3fxVLKn5IZZpSaQjcFKv
KI/h+68tU9g8qTomuLW/EhdrBGPtNqUBeV5n40fwln+3oVoHydstrPeEt6UxLV/h
zFZr3qPWpGfQWvlVyfqwccGMKOapNiV/2ITdCr7cZPt8qsZkEvuEb/mJ560FcHcR
qieF5hnlU488MJtwWLsbvOZzWXXSXfyKm9ZOmOgobSk+fFIfXN8cuzgnmdJAfrSw
4t1oJkmqR01r8qghdzgDqghpugTaNESSoPPAUyDWCSZZwO0c9EbprAVia0GHw8NM
J1HxyhqqhhhBKILy9ZFpjht+lTmVZ3xrbiOzVmTj8Q4Jto6vGy3PX9W2ZAL8oAvz
MyTEGoyU2bS0vRQW3Jjl91OD7KeC7Ex7XH4YJvDESs2PWT+m4zb9z5fT9aJj9bus
TEk8+6znp9VmCh9L92vnjkym1QpAnAqd+0kRLEHAgEWUPgw81qvU2dgNjcrpKoU5
JJmpBZkZapgryXyqltDo+/zmcSds1BaGnHcW6ruU/4PlKoe4Phe7sI+v7Ah2jE5Q
KqXKgkaREXUH+FX0hg2iZT7unn2H+xnN6EFp7NSRx/H+aiw8eEph8lJwm3Ryb4aM
4kVh7M9Lgq3MnfaeQCBxk1BMaVijUGvsgPgvKCa9ZlxIVmF4t70Tr7JqEHiUP8Q0
Rfv4s3SWIgKlfRuqkflk61OK8Y/29d8YW4/chdv7SibteJcgtvUyTxyb9Jc2H16N
khrQ8fVWr8ae1L+v1+DEolFNIhmFAOxr1yiudxk18rewjPVbbO1RmviMFzSso9Mg
o+EGcEttoGP/sYrI4/ahw0gXu8Fda5npFrBA0uVwrcvd6WqhE2LWtr4bwrvwCNFg
hLA8I6D2GwSYgLw058r+LF+bWC5wPNYqmLHLS6Ip2zfvmZr5aZqGessC14HWaxFo
+P75QcDuZlfKMEw+7ushrhYoJrc5oGMQQnUjHpY+fHKMpld8kN0G9oAYKOkyxPBD
lnSSrZxgs8OCuQ+w3zLmm28biTtC9lOfG9Z6gIrK03tlwUKzY/9CBcJadGTGuLyl
cX/lbBhZHug4LCIjieIBxEug/71XAQbBFhGcB8JdFRMdmhco5SglPxvkvCp/8V4q
FPtV7/RXKCh/1vxU/tCrAdR9ooZ/vka3XH71I3JRhwJeruMCqcQwuOtxVh0qs0H3
j0R+iwV99N0JPB3TDXbOeWJYpiC34l4eqJCjRp8EiLqTEBqByyLhDi9u5i51gW4h
owoI0XmNliM0+1JJustJPBCUVvxIlTKdD5KIN5v/K6FcBU8ulqStRy7lPM1b0jG9
9YOlvIZ5BI7rxSxjioY7fNMV803H9/rPFkZRkYIcDbLBYjOL5cDKhB714ZXLJnSR
qAZPfs2fbBESHQrMTqsBO5zy3KhtnIA1E0l9K/gY0y7x4MdVvnQMPDbQuoFKg13O
g3HhdFfduEx2IKiOEdWnmxx/ap2q1eRvJcW4MSN2zLBHkjH9OYcVlAWcsriqshWA
EGReC3oVO0xYKGcXS/Bjo8RFJZiNvIq3MJLaCul+o9LvP5sSFb9Icg4+lNaLObof
XuzVdpBQGyeP0q+ecT/aAfXxrNiWegLuv2nkQ7ivfrZZXlI8kXkOVc9Pioepo3mK
N6Yss6KpmlIolyoZo5rGdhqlwHwcL5CTlHGG5G6Re3nX1QvTJmna+6b22N9jHoSo
LFewMOGeuGxDEfl4plHLpl4Q9C5ARjQRtB7rfB5wh/VeK60HYIXAwYOwnh2aG1wL
9NaG2oW/Jq+qisGHKIv6uGIwAU+shyAksjKxSrWEK6ZHFX7pSUBS/Xm9llIWuBfV
fLkEqyK+6i0s+/RiB1PDRD/clidoLNQmaaK5isWWTbpFtfDBTb+Geh1BrDdFbuDC
EyIh4WKsuW/g/7+m3+DiVLeMsrFyO+w8zawC+bi1vhR5hLyC2/4vo8zKHoi3t+0H
MqueTomNANGEwMHHrOSzYhiwNLVIVtD+NcahwTbnavU03yLTUehulWA/qgPofCdP
e/F0DSEnq09hR7A6iqaxGjBMSWYVMInUnP9I2UFVvBXkrDxvpAKFTr6zSSySYyAu
3CwrT3muEf229iQ9wIoF81i/+TooJ82+ksS29hFzMFbBalHToIHdkoqjm5C43Em+
ftRSTrcVsuZsOf1sqtY0p8oQ66TsYhlO3n6gG4zTQshpRuqaScnYkrzlw48A8QGa
dU9qL+N2pdq3v1Mk5sQJAP/t9+ldgDAIqNR8f2CxHHAa3rBzmPmCo7LyuxPFiqRO
oEkHw6RcNn9uuGoJ5XP5Pk1HRQZlkLp7SPdLVU+GQbx+mkE9Tn2UpRlIktZcDuiv
MtmDPZU8aEPhSck1NqEvNlze8WtvGX3YD3Hhy8eT7SgFde/i2R1sqlqVjDMwdK3Q
tivp9wo0RIuy6kyfAaJRMFilgtJDOOScjhLfr9RbSeFZI1B8tq5zQWKwCNCrpIOD
1QMqA7D4gNWjr8o1r7bgjyF6RanElNtjzxM2XzLo1Bqg3DwXw1B0TNMhR9J2J3yg
nmv23cCYPkpi8faoxQUYlJ0N7aBuwew1zNp5Eb4S2l9iBOYjjVdjyNZAv+cX6Ewl
1W93BUnRBol7Tot/Z88ZzQD3OaEKn4TN4u0Yei9H50LOuJWA/QyhykOefVVVhyku
sg4mAQ39FImraPSvUqWp5xZ5579Hfzb1fcgIq5iBeevRQ+H6sUOUlhqhLe/r1ytQ
tLU7zC5g89d2GulBHdATg3oC1UD6iLcfBx5Ho2kHjClBnmZcc0As3tUt7QyiVpJQ
WwVK39aq4l8knJEKl0KnYZ9tqHFFK7DnSUMdP5aS6ORPwWgqN5+HGtTeqMmlRNR3
qCxfZDPir2/UB7rGxVt1TEb3Da6o7LIMgSNRQ6UObCLBel3AXDcHIoyukG4cNvqw
7BELc+SUa4TLSfoGzFNgS3MGWveFC+dU1R5sodt7K12heXvFE1k9X4yzejqhXGB1
Zefo+XbesElKqR9wq/AWNhhpEgqaxQ9buV8Unk0VObjGLno8bZXGhF3+iYTwUVgP
rsvedMU2xoqY8xeX41yLbMjogx74+Z8z6dHusFcWBrzn8vevX1Bfh83j2WaBMxU8
J8uPWVoUKgbyzpCpwI2f2iXsasQsFuMDO3RK5ZD5SdsbAycgf8UL0Bjp3PxK8rxF
75r3NpzMaPxgsuRh2dBCRZh/a8aTEUYZjxKHhjJHJ+5ROYa4AX8tOJ607sR2e1Au
IIjz9hQrNnbcoc/gmXxCgdHouhLaT7iDJDj0ChWYS/47IoiAG6HZR72iqe9j9zHd
c87uaAKTX3kcWlobjituCyRePAxfE9pC1nEUjWBBE4ol4/mStaFFbjyh/qHmtvDn
K2wn4faQgPRDyqz0P664d8FjCrLHzVu9MCxxral/YVxkQ7wa4ICTUPYxdEsMYcO3
uCSdyWH/N4obgWtkq+n7keHf0OBIdNEcLIOMVC6uccevTwm2By7EwIvUJOrvQ/Vv
GTC2MJv0kF67KStq46yVdp5nMs4JiGjVoYOARG7pNjj+8X71/OyoVD/4jUOyTkiw
jriZWZpr8mYypQzm9Hf/xPPCV1FL+rKsMxKvJynP0Tc5nB2dOgWQ8KYXXZdYeXPm
iqgA4oAbtWKXbCFWiS4Kk1Hoq4ixKwDTaXc1w3eo8T0hHf9lx4aEBr5bKcEEX3CG
PDvPaMuF7fjJ+FdCevl2mqiUqveu+DIgT6PMb4esBFwTfT76mkSQy6f50Ktrq9xY
BO/0us1x7CvrrXCGi/SXWUdTcXdCvGvzFn6OaUW+U9DTorYTIp0iwDVsjPBQR8dD
UQV4UYQrxqQamQsHhqQ4ygq9tdJdno6FgCI4cDSr6RpXNePhyyLb64A1AEh6OonV
ssz1rnfAFQu3JozDdU53oUy2yK4e5uXurLns4m+pYcdiBcKO4jeB27wrb81gyfyA
VUQvpHUx/oxAso2cuYA66RzoFE/X2JHlNk/hJ2RKPfJ1lJqZJBpEaoLiMtjAsi8C
+K4wcuVtaUetDUEWMDRDMJwRpaGjVezQuhA51FTMFFIMBmomkFOPCrdPYAw3Cmf2
GYcfBkBp00hHB3Lmyzp3nQtJiFNKlay9ISiESyVZWNkftSljlpZ8WeqNSv7bx+lc
tKCVaidFxWVZeytgiQTPGMvi+pK7DIScK8rYagYEa2AroK76EpN0D5DInA9txkee
spJ6uEpyvcEelakAIPAorwFVcUHJXzUOitv8m4/iY5o7y2eBdQ2rBPiyf3qPbWGu
vhJH9VpvOULoC4pTptPceEe4bGpTQAMFzEdU9gEgw73XVwwXfoSq5zpYB9cnhNCx
qMa2k7IH/fXk+3EoyZjragcJymOaTJ3jaG4OZyeHECtFwwXCr0+zcAzEUvdGUN34
Cz7UW/A6gcI9AEgCJHZR3gw2x0HGkY7Bf31RqQYqRn3dKm3exsNQO62kjR1lAUyS
dmuzUSECJtOK6Fzz0OYcooQDSJfczTs6dOrSZHE6bU7zxgMhqiDq9MW5pSPTkT3E
feOmJuC8OprkcwcLFlQd0jcjnPsr/9e5s29oMzMJGotTUZd6OaH6/MaOYz77ZwsP
F7UH8ymPfYEiaQ3j81wfinitOTu1xL1RT/LOI71mlcsRhQP76lxsWRDse2NF7b/g
Xjkh/1trGdWm4/MdyaRIVvUvKVoYOnwQTDhjtJtoEy/K2WWPZuqNVY6ww94saPOs
WcavtCa7XTdKzYO7NGy/TTj4yzC5W2rvcKBSlCwja2JLJ1PBKQQG0GSmQy+Pna+I
BSeTYj+pbdCEyOl2BEcuPNXpYcxi+QyQq791imqdzWSAwiY1TD/glHDBdqDz6+bf
xHO0SWJ6lyamBGbZ4Fx7B0wDsHV+kHokDdtX9Fynia0Gmyu9jnmOfr6OTTVzCQLZ
PjU0PXeYDf9jeyS8ZvKuC+Xxpu+UXhc+ZeXkodSZqjaVG/otDqcGKyy3I4dZppvm
dPWcqSVPJcWQPfnncIQibP7ck0X8bgz0IsSj+oa3SCJiNdlRPlFybD9M4xFq5wCw
I2V+GsaQ+zCDjLRmjKT29e00oIU77r/34cB9ciKMwFuhYnF+8UwreCZYp7rzNUjv
SV2Ysmzm2vs8PAiIxgZxO6Z7RedsX2yMNBMLnZ2I/tWnYrmdiCfYvmH4IYqPyPF3
z12hgwnPld41mYN9lF/2c9Pl/a3lw5OHKUWxhVBVmfHt5nxiDomZmGxJqnjJ8t8t
votkGNpuyzmuVzJe9TXQI9zWCI2wytGxP9unv/IOdH+TmzwhZT9J08474NBL4zJ1
Nhr+yRQuR3PI2UdGeE/KFNGHb6vz29XHabk2ecgLiDlmQgODFqjhxUKIB5lIuou5
KznzwXmpIBM0OrIByagdvHr3gzz5rSZAV47cW29BZPVYx7fe3EGr4f8cVhO8Xdwd
YksScz4OF0doWTaWGQixBazLZEplJfwrFKU9tiyY99g4kBBOO1vnG1t43X7k/t4k
3BCBDWmgeGEyQJeJRFZXXWL15UasZB3WEWmm3u4o828lKreKkrexRKf1GsiEE2/D
P7nz6o8j5HzuUA1AWN+wJqMTTaY6lFienxjEEvCfllxeOBJW6P4YjmQVcX/5KC1F
L0khKgBsk9Vfe/hyr4jmN2DsGEezfGUowsvq4wgp7vNQkL8gOcfDeuXulihKXDiS
Smpl+qU9TaVpMluZXGEb2fubwUtgzKvXoh4Kgmiuzfc8Zi8PS9LOl/5Wfp9Uit+4
QIvdAY6SzyAX90i/GCQZ3sA9xekpqSP98RuocX3WQu6up1X/wz7bEbx8lwSG+854
gAfkn4g6hY6Q9JbtUJzxyLPILnTvjtmKavuFn8lHA0oa7T45IgAP0gh5QlaR/1MK
+n0VNjOz54QSarTYFznzdGZNEgWBcBn5MODgYKdEUksM99dWf9QFlCaPbEVth3DS
bQDcVq7PVT/P+btgut+v+nCfNN7AruZDLBahkfLY4o+Ylq1qOkOKHvk1zVulS+q8
f9VKes5LSUfd13DcDPb3If3+FPPg03JGgyjH2BGOstQwlrclfTx9thbQyBzl0VEn
c9TrXg+2Lxx3ESKtoQPdZpoT5CQgq0miosJeHNs+HEI8LvTa1zODa1degdRgn2Vo
eeDSUoPgRSGgrKkT1ldYTu+dYIf3kE0QqPJMPaPSk9qpFOrxNaTl1muvRj0h21O5
FfH3VokubIup1p9/JJs5nmWcmTsRs/LMWX+wBUxqHfyjmdoTp/jxRsYV5Ri+n7fV
oCMosM6Np8EtIvqNxLDYc9Cmh4fDvOeuKHqMbNdPhRmtW2mit3Toracfyf37A62d
dtxghgla+3w8yTgQ6ppntTA+ef9RksjFBHrFg4sUAiCmv0NQVkxiMBPQb0RfPZ0x
r7jmN6M42p9gHR18gqP6xPZa3eqw59ucaVwi1Gy7maij7an45WtM0yvyGwO9eyF8
/4Qur1lwqJ9i4xgtpkoFUj+T2JeBeYmpaz8U+ikzNXI2prYuYQiZSCrZiQLJfG8f
cTKhqUL5VkihkB2+ucj8oSXjfC6SeX0+pa2mOaPal+k3T1XBxqafha/++jnw6fyg
OQoKn3C135pWH7nNR6NufAs5JNASSDEQTqPT2yxgZY6AE/OUl3LjdEqxzq4dCKsY
gNAsq73MV3j6GaIqodzYgYUJXRabSQReQowWAL7I1SLbmGpqTynSejKYmy5X3kFm
DXrkQ50epZco7N6XfnDLT0mBzPDSjN2BJDh8uXdhsKhS6oBbeOdYRx5THV0lNnkd
moldNSk6ThymBEI/AQI/A2tJbl0LrCWz0FVQoeHr5YobpX/tR2yw3WB5/pk1nV6z
i2i//t4OZVezVUSXZwQr+mbju68wpTAUUboasQWLSXIpv+CNMwruuWAf8oxsnFcS
al3Ed8NkrhO4IkaWHI2ES2Sbs7Zm0Q1UZy3UeNQ0aPzh/KF/KMNuz/05in0vdQVa
hhkuErDbrHhNqFBEmYo11blgJgtQ6DF1BPQOn1NHccBr6XQzjMkbnLc6uE6Is25M
Y9hV6l8YM+JxNulWLMAL0uqLr15s2pKX56ICzr4Q/NxIUyI8HGYLx5do56nIHJrG
CDUpHEqxbnvlIjJUql1+wolrPcmHHAWzvZygkF2mAaEv2zya5gR/myqk8V31fMPB
4MI9rmlf5keFFVj1682R5jGTOtI0Nl+FDLh2NoaK9nsyKPiBLU43nu+VuzHa/yxL
FN0jPgNEiFT60kbFqfzFwDGwlwL5eRGQSVx7lRT5tUV6ZQnN7KS7hX4T3x6iGCwI
UyzumUZd1qKbhh/k0WgaEiLDC9atXkCKMPht6pMC+pYwXwPK2KucxdriCdioJHWg
Px3WqcU6sIB5PS7QULnNtn2/VsaEFBeNs4kVrpV5sYwC1xs6ypDI0KABDpYWk+tI
IU4wHKdABdaJxzxxqINZpEqy7FtJfV6hbv0WE9jXrcISYT+lyjGv9iZx7iI1AjGb
+pgCV5MwwzIg4qLCnzwMm5VqXYAmOIm9Sqn+dOILZD1jrgYsvYYXqSq0arDIYlQ1
algyQyd7fRJ8/0MF4ZUAWQQtNmkOlyHCWG5WPEm4O3IdsFoJHk++Z64HRURhXle1
7x747kPmsdUchmJAcbvr2b9Soxn14AJjwiJcB7HpU5CgrGALXKInQg/za0ERl0T3
sdgN2TQ0qFHTE5RU0ffxBUfuq+PvqqZlFXIqFMPxC5OQqaPiSoEuxFBC0dG7Tny2
kI0r6Tf1eTHhiTiS3O3rVO+x824VEGxHT1zIFpmeNWb+bBiYZLQYKltqcQorKNTg
6x/LUZHkuYRlwNYZj5TL/vIVsE/UktpwQm6DCd2nNvEHt372XKcq+6EIoHP/7/OB
azvebHZMgNC4NAit1SFk1PbnG2NOu9M3CuE9TgSWYeHqXVMI9eMWDErsQdasgbSg
jiTmmnoWhQ0CWDC1Iej8LahzoKQHFIC364tw0ehBWWM3yREzP6vPIL+mZcaZ34WV
gKY890hNFQmey4VNf/xJvt1dmxQ4ijjdcRCj68UNrYMVAVhUnSDS2XWWiLqBEEPc
grS1sKps6/VDzntCpF+uq1azogjbKznbN0M9tPKjsbOyIX3i8UnZp3UbVBZHRrHJ
+DpHGaIeUMXdkL/ZekNceUI9w7tCg3X1aBsb66if240t2klKhesY9ccobDQEqFvV
e+HSCP4bUwYuNm5KW5FabPPDU99dD+8Hg/f2Lwsrahzunn+4/ULWhWF1iJGjtGjw
UFr3lMzyRdTzzht/9Lbzl2Ql6iYkS2ILGQlttxTFsj7rCHJLhja2IBeLp2L27gl2
qFWvO1TTbMjttWzCq3DMaBqTr+wmw/cSnG3U1KRpp/A1nG5TgCY+pVPshg84Q8H6
eLqZdimdRDizK4eyInEkR0/EqlWhuFSc/3BDmeOZpZWLo5889k0dJlr8NowlDq6a
Kix+a23nXDIQSXVauYtpVl8/Lw+Sn0i/USuDqgK+ql5gahpSFiZf92eGqmdAxlhV
bPczVplvpKTRMVggQFboI0SLLlmOznUw8r62I6U8WTYxDeaccuIg8d7Y9jAPmPBn
nbkonqsp/bvUnHRNRhc/17fse/t8hIaxQXoAcbjD+BkXeVA60KExOvGQHBI3ngMM
7CFCZRHr3wKvKda9GV6TnvpuumlWg/fS226HEgVcp/trR+7Vi9SDY4WdFcbHwtRn
zSRv800hVGlUpxqfXvRDf3pn4WiRXpIlQQsG/tOA0O2YbP0Zc/56NOJVC2ecDN2w
dcsYuT9tTWDBHkxiwmjzVcHuhwub0dt5ubb2xFlt498n2bVEJOxDuhnHddp3JNBJ
OMp3D835xkhVYDXly84ZO3daoO0/b7Sq92JCvtWOtqWJwAOXBLHOeATPvsl9pQvj
fY5DgESGzPr2+P+wZ1dqUWWHKc9M5m865qz5DROYHPm5VdpLIYMBhwqFaa36t2p8
oAasS55BBi/79+WGszUxuPE3gXjrtEeqPBxWuoA1m/IjuDIqxy3llfWrRdHI9bVx
ebrZmsAsV7USajyjas/54waFInP0DOSv3VvfxQkLROxVghpSNhHHmh+KBQoO2kLn
qfSYApEva8gDFtirVB4LnpuJ4519j/wl6e5xc/lX1iYzG5JStV3qJOL8b3VJCZEB
/CvkSzkdLJsxEhn/sBV/cmv4RuFLHCgkw+yk5M4jsUNClbFWIuNPprUuz2ofx53E
fiNgbyaU9unsZ4wy0wH4+KG/DjEaqPv4JbM+Os+HxINPnePm76D1rqjPw7YMAnux
S+QrJNErDRBZsrRwL9+uS2ZE+kW4Qm93xbK2GivvbqFkXE4HqFCL8L+U3m2Jm0l3
2g9RkkR6JMhWXgWG2yyj8c4EOUw+Oh3ZyLnLwd1c1CHXbWWukmrp3sMLQ8beB91w
lLMfEUtgV+iHbRXO4p1FF2ZggspVf1h+Fphd8EMufJ2syzX3oa/c2ZiBckaBM2h7
p4+xTB9OhUPqxsIjzSRMEFIbhSfX1IYOe+KL39KDrLWfJZJZm0LcZtA9DSgjhy4M
vgjFUky8Np6yZ9cJ8EniV3ml2JJN3guhLIEf1XwKuZUS4H8BG44aHKk2Bu1iaxAp
bDvz6U/kSesUG/BCeGJNg2qLurTHSZIrte6oKSLdaKdMZZ48L3fHuikPu+xzJ0Ou
TtJVhZWQskHLSQqVpsH9z4/9BeUOKZj+AbtLMKhhYjmq09R2XM90gqSncucx9gUu
f8c//BIX6tQjdSCxf2HNyOCkhlD4r0sKRVtGZ4uYaI7zhbcI9y1BYwKTSzkXswlO
aRk86OuRUxlBrUGoFVpQ7eZ2K0MbWs23INVWM9cpacMl/P8SpwGqAffrSKdFl+SM
iTdskLrNoOkZ8b6BUfwaNFCTEuIoNaHA/45uz3HbdxlZMXqgzAIJUneynN95LEjz
zHkiZszyeiBL6f+V6Tc6dleL8KA0at2r6kzvhcquG914glhkH5WsTvSJav6O+sK3
cwyPktNdEDIqNUJX8wXnYlbXMrSC0WSSf8Bys+Mnvk5OTcgv174a3+O35zJa7X57
+3RNMukNNxYeuwSWrDeJXi0Et6iAyC6txLP3O5luT9x/XwFNLjqnurM1pQpKzGVa
jaLcTCiO3gS9x+k8iL+Ekwr0GKOtma9qmLf2V4Q+pABBrGhCsR9xtaL9PtJBiznR
ujEdwMo/PjOIhRr2RjBXMrCLxoVpn2HjdahRSljXrV0hfDfcwSTH76HdjPCHpkem
v49c1tdnaVH9rNlOD+snKrbr5zlPjZEpgUQZRCvBc8wXtcAUEHm1WZ+wkjAoSRnt
DaEfWY/K/82rbnISQMOUKC1+KAmlLU/aYxPdfoCY2sd0rv70ioFbzYLIY6IhxEJ3
OghC7x9sMcLPpx23oAQIKWo2At0tKKKBkLlB8jieedmpciYyG/0BrlN2QV4Smn2F
TisklqjH9X+xeGfVcYtI0HT5iNgcoNGInLHc3zCysZmtp9J5ubhFRgOuhUCRIvp0
IxRubs6uUC+fZT7eEjnVed9qQryjB+Qn4cCW4HdP/FP426eEENqK+0NoOrlPeJaV
FOlDvfyMjY9HVKtdGShOw0XcTS5o42Nqi5f2JxNfJlgL6CjBlcCMImmkjVVB4GNF
AxorWZzcYN8dVtYI3ZaXE162PxQz4xWkFHQAQoobtxtTWqSwHX37AdhsHVwK5daT
uwzW8ssnz5EAIkU6QxUJz+PLWyx+awVwfAZZAxU1V4LhNcxEKT0dbOsQxsqJQgmb
rxli4vHHob4l7KSCKQ1J3+26l5Q9WG0Z6d+6LIVe87YS+xhyR2xs3k/N49JEbiG8
AWX1fPPIJ2eFlaHHhZ8el3S7IY06DXZey9jYUFzhKjgvfOvnrn4XJVw8jRMg6RvS
5h4sHC0rGbtHW1A8BVB7x1E1x2HpJ3thJ7nrEvhZKf/apuc1QgQLv7CaOCml8+Vu
ITguTitfwskAAMuZS9OUsjEkL76mPpAPf2fkbS47uNJuQRO2Eu7B/1iDe6f1tobG
nElNzDWx6m9DUQ7ojaNg/JF0BPKOSfOyh1pRP+TLWXD9CeFRKDNU4RmlGcIl5Znk
uoe3j8ytsvDFoYxEiXeDqSMypkjRhUHOHuvZussXoo82BP56R7VFGAmGKRo5MIQT
Sguw6efkSyKtPIY8vTNJPPfNuLzmmic9xDwgKspx6VCXR2KgTMzreLUp0/yCX52/
KpR76VpKu8WqiGnc0ac3HcsKsjQBjm/FCF2hrK0WS9Bmpm7dn47Zd0AjBKPbQoF7
SQjkx/rAPeMr6xFjEYIHo/ef2GVm79fflEJicpx+Il87EAvULe++nRaVKonKDzPO
3IcBaed8Tf4F2xjwujNvUsE6+QiyAPk8Pbsv5/hP95osmRzVcOHzJmNVgIPtKALa
tl/XCFXaKzJWOoUO2snMbJee+ll+5H5sv7EHaFXUmWE0q+/wjjq5yZkq4CUBFWeH
pk4nkiCvpCW2qYTjVIY1jqyKQonaJfAe1QVO4jKXI585kBnmIweEETIj+/GamWbI
oVdprCrB0YBKelpJEOZ3Zd94icfqYk2shogwW6kFqXMxtiG1GRc+i25pc/2ERg9P
w0QnRIfymGikgCq+I3VsxHU0HOlA4oDxrwwWYKx/l2/9zea3Pj3NFdFTiWcelnzy
4iTZ1Odv5U0GLP2T1W7bQsOdcWvZYs8afsu74vnW5HWMvr7FpHwvBrdDOgDz0cm2
4GMT4K2C/sBK64Ahpkr25Dez49aFBExM5gcSRwGBFDo0dtQ8pEEsxVa54zngtFkl
LULQMFniim8GtXpEaLmYFuSYsDeiNxoIjhwTQFyjndfK9jW2hMj8Thuy0Q0Bfpvo
V+10lMc8+vcVbKwB9Z33MchsVKyTW5jPoF2/C2LMKXaEnr00e2TcrR+09vYB22xn
UTZ0v6Wfr9MZFJl9qqpS9q94OoLknbxs+o33eVI08W1i8Wz4KHLGvpkl/A70bE6l
lDLvM3GCsDtvIR0bVurCxC5uN6tdvjxDxW1Z5Fbt4szV8uz80fPdtBO45uTCe8f7
Pbxp+Iugisxg/Yu9kn/CxbbU5iBoX21Wc1I7H0n2vjW/o2ziI/7weDZ8entQfWB9
l/6RMm2oZ5z3kyqF66meJcQLXnzFpRWdYacPSzWe8z7wjWeWlyevMz7CtgmF7wSh
OBdwE/zfRjyZXAJcmzVBvb92hmkZdz/xCvYK4ictvr1H4z7wp36q4mN5J1JQbF77
dcGnjKo31yjSHyrsg8d7NIzDHv2uytZn3drduz2O4sOXarsExGLQAzZKU/hxDbx7
aPA8Vn4nf4O0vAFd0TA4a6z38+dgHm02pps1fK6uv3tD8DKnZQ9ued3nhEWshDZ1
wVq1/f6x5A83N3ZtjDWfZpc4XwfPeYnW38osPZtmss8F0uVZWLETaNNFZiTQxe5D
VAi1JoH2Np1Kus9xatr8cFVpr0jHfp3Wha2XOtI+GCijt6+Nq4VezDelJkuaGD3C
bprjoD62Fy+sP+xgQ4gBmzNUWYXl+3ZAJRLFu550tuk+3foIMhVgIYXweARbpQBO
RnCvVZmqSrzirKuXXVmDkS6HJeKeRPgP931KVDGnBJJB6rtdD6W1F234lz36PbfF
L0sMyTUHk0wGdjwTcqgUYXsKWR2tdllukoEavVFy8rSVo0WOn6lidabY5xTFYCeK
uWeR2WM6WCfYSeZA5cnHdTSPCeGgj0UMvoCq2YTKTMKUp5ocTlZoeJsnUgJELOgu
QmcpntouSuwIIqKsHduVC6Eydkx/khWHrjcAwQql6AHVNbxbZt6gJN12RwmWH+vm
fINByQVGR1Q/SjiWOfDpgIUnt7HsN/SeHV4T9xNQ9cW3fJj4Zce99sy1hIlLqNmj
u8U+5lRoWLLVJ5FcJLDU2UyY/kEoN8dNhj1F09pRbJtppXkqVegOlcLG6oMNyOHc
Pcy1uWBqIExO6djqbXKuIM4nVn3p3S/fa3CwuST7vCXG5QDCveWE6opfCWZFNUGM
MyBNuZ56YnwIVHljiZeoNJ3wQOi/1tF3RIxqqMrtzzWIaZehuHyDFzRkdlI2S433
FVrRiQoKhbLRHnUTsJDmuc4ahFOZRg3Dbm+D4RRM8r2ni4IV+8aITDVZw1/E6vm9
Nkt4FcRGXClUBZaRws0/AQlZi/i1H+iqLmhSBhvECSW21uVCF2PjiUvjQ/O9TOuC
B/RSznzyAd/LXH+6KjY/H7Iiy8DVCKIqsKyE8ONWUSyuoLP1kWxU6egsll8uw04z
R4lpPyYZb2/ahBki30x+CuC5owXz18T8yqyTODNuXOkdVeuZY9+Y71yY5m1cO/sN
wC2Yw0pHiic85wW8sI99SJx2LxWGJQ0Wa/DvroHb1ewnc6THlGC6rNiWagY96WVv
huonhBHTe7lrEyuCUw8D8OKItrwA1pr23i4XyMMK8hGxgGdXx7B8o5OUPMD9DtVI
bkrSzK9UGUCA6InVaEejRJmPcsX0yplkicepSwtruiSNhiz/02SVH8jgag/h9d06
YGNlrUChvQIAt8ncK0BbHGFJFRnbNkWhVIvL0Xzmlf1rGS3KJLOscPwWiKMrvsWP
5c6xyvuIc3+4+5zU3s0KYcM6sFoGFVonPolHH8+qh4+E8QVb9u1IX8XabwuWwWUv
dNzsLHEkPJXXuSEojrfUQaYDJjjdseLfeeQ2nXQDyE4pEo+W9ne7DEGWNs2HEpT2
swJ3qVXIL+BD3YC/4zXoRl0y5pin/flKk3RHLbS2Rvu/0pqrSJIdYDHJRl+r2cGo
38ZgAyg2ys63KJsLuvgfO+mX0k3/haXKXoWAet0FTJ4YbpVXhfhuEH2uUSjvPYbc
6O8gzTeuyPKh4UZlyoN0qB7Y4T5BIkeqe71i41QkYgFihEAXwNPgMXMTY3MdTDk3
OHg6pqB1lJhZy+/zr59qfVJYXCiKv/PaZToRxn+DkqZ3JNReu0ZNx8v8mc+UQVUr
Kgbh4qVkKrnzTUh0NUw8gGQBWSq62EoUkVFEbuw5YeGBZXim3Hbo32i+DM0GsTTP
z1YdsvlhXJZPXaTImfzDBuDPV2WYmnwNGgPRVdx/gK7Ex0WEdlhCSA9x/XVM6sXo
+jXw9Q4i2ZtMecDl1oAZiX054wCbS04BCz1ShEluuiTLcdF+DVVoP4o/sSiISN2O
kUdJT9gzfUEGDZHxPz445eOviMG4QravtjnD9MRDP+ydjqaB8Iu8+oueaxwXqiWv
d7jWxg5YZXCCEG9nxdO6EWdWmT0YF5Vol6xu/+vM2DPVf1NRait6oAx2bKuleSMF
Vi3anqPUcmlML8P6enknKj8VZfr8PRlhDohFynXWgtxWS9+1Kfh2OuG6lq/J6bqB
0qpJ27gN7luX0mRsUNXKDgDlxp+5jcrxXUn5uHbDVNS5OlymbB9d2P6Zr1sWIEaG
2ijt4e1a9x49/nO+f8rP9H6vVmQPtRkiKTWY6GVY89Xc6lwpumemvjEOUlHT3HT9
IKUf11G2BYLC6Fi1iwMpXDUVKMB0gRKDapeU7Rn4YEvpdH8Mpr/WHNtV8Hx5gKEG
k5Zv8V3vr+kZJ4jE/C8DzOb/Ou8BK1tDr6gzcHv4DBHN6zd2Kp25kiyp4HZJ0SIN
isfbST2DpDFOyB/+ZaQ+igoHSEkCDv2mHnVa2ZAkq7N6r55w9TbzHE4D6P0LomYQ
8TFeuTYpJpYwMSpyakaiYVsdjm8t6fK5DcSg5hP/qk3TODh90jn566BlIZ2KerZI
YAza8uTC+BW6ADVAUu2BsZrXAILti+2fMXVUPWf4gfJeN6/PIt6K55bA5AgJOp6A
gu/Lp1wwyjst/CnsQVKHL4RT2HDCVW2YSlp6qTAebjBqBXOfXLftbmXYa1BOcFTv
jl9LIMLbNuAlx7j3l0ZaEmk+SWP2ggQ2I1img64ht6RMTGJeV50yQag/WZh8EgEY
a+ApVmRoHIKCVMV++Xax7+nNKAffbTUYKBD8key4v6LWcGpHMH3MH9ISdZ3PF2as
VGwa9K815O25snMtivWkf0Nx3AXmwYTjbMwB9NTXYEra9UAQsfYih35AN9Bm4csp
p49BZygZ1gdolF/+4yygRQJi/4PA+nt71GGjt7wKrF8YHaWkY6kGsQ1Q8NBJ9hTz
7xs7dqzMmKWwDMcfeylA/ZyanTA7F2gMU+hJ+hgsJH1S0H8stwi0Tx2pEBZ0AXXu
rMKg8RFKgoLnx8+pFgYoMJtKGkIK59UtxH8KH5WtzKA8gNaNe3/SlRX1L8mUMlzZ
JP/DYDQqZ21MiKGiWu1vzJT9tgfGRw5KfxHrp2ziNMKotJFacioMsThPbRDOSvE5
p+ZyHT9P297Oathef75ChlxfaPek0ZfN/eVfwrZ3tvT15P9H2VYFzG5/BHrte4FE
gR3ZXSNrubzdjTAdFpZZqsYg8J6t/R+70l/D5iT5NGWLH4bG4LfUBg1LhjBUn9aa
m97Le1teRRfB6SY7oxuva4fYeFiVmnx/HcCjWBUO6WnsXeY/+3AqvW6A7yqRhbDN
3mic9zZARHZndP2X9OHKLZKXx7pR4gIRYGNmn7W84w2xHDj1+qHnX3DCNpLM2uqP
BPo5t2/Y5c7aa9BbJUO8dFV04eybLKG7sO9UsZgGVMKfumVuMWQJ6p7wr5Juq+8i
AHqMYNIF1WYNF2Jxc33l7uX5vUTXfpr0pUG/zmEUlvLYWQBtBtixI+moTOEZKs9y
NcxHSUckJmzYg9YFgu0jGg2zCTitgznybMc4HRB1LeNiM2eruNApa1DwUa69LeaA
EKJAoi//Sv7vR6akLBWIegoJR0aJNyPBbM9sy0qomFbfxH6rUeb0Q5tpzo304rfQ
kpGkn77Scd7mU+Kwnk5267ZjIS60F7XpZjT7XplAU/xNvN/eTBWeiyFokI6bYL00
bOFToMh3u9F3/B/9FVQYUCA35eeWC3EZ+6Q8Y+mPSaYetekgOKunSPzKhk7vwZ5t
AnFQv1LV5Mk54wnDEtg6mWPn0Vrs3vl8GBqfkW472KGfRyutmYFjriRVUz5BUD0g
WPT4W7c35DvE5DVJXofdBewMJWH/j5U5K+nnP/fx65sn3cD+Nn9I1c7rrFfg11MC
L9Uivr5gHeokLExgjhOq89qZHholZMzINgujQXbQ7idzkAgjQ12uT3HqugAcDUNU
ujR/s0YswScFz1qs0d0sNlTwMiIiYAHKun9FLXg6UU+Nn+jAoz78bZwA8Nv4B/si
9cZdPnIWpfsn4Jc2WkaDx5xDjHn/ZktnRXx/4pJywuhijr9dObeNBUdus0U0JH44
7oArVVoDUlz+nzQWuoA755U7cJ2pjRK12TYfgwdcK40GCZjGV/6E35wIXTvJL7Sl
LYHEq5DjgmxIRG1xcIjFevBmEmYyBlc/EgjAqMBGIwq5QQm6nD9N0WYMWVvEvNiR
bOjdHRAh4qnjKr2WBxxO2HniiGRZJSSLhzVUT4M/2BR0/zqcbVeXXjQGMoFJyCKN
yt0LPOL7AHXTygbPtD1NcmhIZE4yg3Lt8oEvgbX63H/AQgu3CBviuQbagwe+E6i6
PNsMpOoJhvlnUqX0C+SIo7Q6S2kW6xP8u1c2KvAceluMXwbsEfIt5NVRsY6/RjPU
11u7wqfYXKJIx9NSUPDWQVhSDtMFkEaOIS/NNPFSbyewGQlbR0ko+NaFKwh6cUU4
Gb4PCKy94XHyVDKu07Y9afrZeHF5MnXD/e+PZnOFdf9p6KXu24SblYArNdDQxUPb
BvZh+iGFe7MgMuoy/mP3FaQBjzPGT9SlNoObAHldwmMzX+kjOVXC/gNy9yKab4x2
pNKoi3srPFg25mQ/m0Rj75UpSe+gZEYjz/fxU5jdeHqwt1GZE1tYlVj/japDWEgw
AtiJuBGAZN5R5T5Ykg7I/BSDZKl8NFMeEf/MKyLHw2R/EPV2ufph/x04sra5Mu7p
D3NbWqYD2xtF6qJXPMFRwcf71IjAI6XX+/RW0AphvCSUjzFunxvykqzD938OtU8n
5TPeoDy56I1tNq+SgMFYKqsj2iKZvI3bNypwbW8ef7lJ+2ckMMZmBu6QLbJmgIy+
R9WR46Bj0HAHJkn7RNIbHpQ6nY/2KvH2UJ11Gy1sQE9h5z6h7gPPV1zEVlrLFgDP
Be3zuNx9iI60kRR4krAVdl2JIqBg9s9J4G0t1NkhwOms52K/eIk71wvRvBwq69Xj
IKjslGigbJlBXCNHmssZKUKlRquYZa8bAfSBTK8L+L8Iq9Ct3sG1TZNZtLvEK2uY
UVZH98PSP33HhvriMvsx6veVJ1Gd5ajbdboKOxtUrmHH6ihzvxvMRrit+P/RYKcF
ScMh04wBME9h5nNFF08lqPWYsvIuR/qCnDku9O5AxPBxaTUp9PoTQoRXrOlsy0Zt
2U4FdfXqIMjIRKJg5SKGp1AqqeUUJYbsxGon5kqg0r+W4goriEjvwS/xEAhbDv2e
Ghvm9DtjxRc68OybZD+n0T5o+YBE1blxV4GBBzO4AFb1dYXR4tV71R2ALG6786zw
EdMpAuH8P1VEj33UlS3z7du2hrBqh3Qcn9UWHEl4TPBicszxIgmA6Ekk2175Anqb
MmEpzEmvlq0FcOhmBDzUtsDdsWUH8A7HcoX4/R+fQpbpnLyqKpQQod0Of9hD/3Bo
CCDpkXeDIOc0l4IbJ+foP4H89qK/bJlkz5oXhHKM+e3eVAjGo1Ees6E48rKcszn7
+JuXbWdbs5uI4tedOkvUtgN9x3d1C34sn8o3auIjBvAkveMv58aSz7OJmcwRNx90
M/XANLLxU4rvbjUwyO/dagpKYqM64E4M3L8lF+eetos+ES9YgGSEbPepurXiB2/V
MEpaIUjCCRlOyvGMV18Z3xJz5gVxwXZ/Dz8J5oE8CykP6tV8iV6oio0qZqiGXqCJ
GFT8ln6ppzyo0R08HEVqBiJPquOjn3hUtark6hEHlekOx2bRraedJpMFEvzbVQ36
wbv+E/95obGMJdsc6vDN0oFYuemxRhFiUfIrFeLPPfvB4QyK5AaOvBApL29Ugz4+
dvU76ROYpGi6Tb80FA9HRS1ctCBVPqeb59itBcSsSrA/UYBcLQqh2MNNVIS7BUWK
CBVo+oaMB9Ctl1INrOMYX168RlSz9tSmtFYcx4WBfIQeQ62xUfDBcjZId0oIlA5j
ifyUe3Dlbk3iKaPqpA+6UP41EPiZPsjfpUWVj2Ev+MsuWyC3qiSLz4dEEm+swq80
REAQVyKLBcSDqWiCAq/w5m+KY+0yGEsYzV8hlyGXf24BahDXV+2wtFBt1s4A9O/s
aXEY6HvO5IcOAZllc4VmCwLCx+floTMajFYEm8xiCIcJLyu6grtFKK3hGHkFYL0W
FwWY7HtTPe/1i+rxhn8nChozuE/Ao7U8a0rzUFnsQ3TfRkeActCj4w+cc3W2wVTA
TY2HShlx+76UVTMRPofmjWJ/M8w6Iu9BKmHaLUxNhSlXK1lNCLT8LQQEU7c1DfGG
elrnd6WNt/WS2zZFO92/FSuXSVFRAx9JeZhSqZCBBETorLm0jw6VLcbCU2gq0YMC
D72d1N7PojWUvJszcK6OxfUb1Dn2+YF/nYY13ZqOR9gLJsWdPA3UYlLg0FiV0CJZ
P/if/pQOeNLUm8blegKvytKoDtGqwBfsKENgTe/rMcmz2R5xnhD2vBJwCBrLlbOn
zEsmQoqZNrOJ9VZKBGxoQlZedy6JUa+mZp7Aog7K41hD93bV1d7FRENFBZ7SKtOa
7SsmnDhcqNcWveJUSMGIITCNuLAdamDwCv62C7ZfSqAMQjcgzOuoRJmZ67av2oRx
9SFP0kwdAqd5FtW8mZjFO/Lr9axT8J1kGC6FVuiB9DJOSadzjHxdAUEs2lXthHyG
VYRA/sG1B86x257p74VgxEVQpwHxxdjMZR0ggQy0bZ2Rk+bdCZytOKZVrWe3Uha/
yOXQClvoEKRfKdH9j1MWKNTG1XAaqJOXA/lg3D5Bc4Py+L5csUZb8MPp8K5d9VUx
/SWr6dgfzQu1kus4r4J0eGMciw4z9DgYZtEZ3TJ6sM1ufWf3U5AsSkOfjqxehif9
+oo+bKDD+vGLTASAhHIeNowBShTQkQ4JNzzRah4nkVUdwdVMqcgGechzbnqHw91u
dbSmO4282JHgUWnHNf96cIq3RhpOSC1QJ5dy0fkZ/k+YasaEi5dgh9qOUrIfP4Bo
NkawGaaMjkE3IWmx3TJS8AVgHkOARXJLukfReWEljZHNUa8Cq7ZDKJ7vGc1hE86C
eSwCD4gohIyGItzmTc08BQH/aY3uwBS/CHsc3HezOg9QcV785DmqfIlFIUwaeZW3
ubZcqI1fp3l5c45vtd4X0GEhAlagshxrzPWC/XG54wt8mJqmac/5JDydgUC8qxdC
h73IGGRIy8XhK9+fYPryl/bZ69IpDbjtIaSdZxeOaLrOiWEf6XGfcOx4AVA77VxC
RczBVQbAfjz8hK0Of8K9miwnPG1eXzYiZwtphyhzXwkojHQcA4pnVVPHnWrhHaJ1
kGhAbK9whVdmoyCmYDR/NHQ1cmtG34MdhN35jcx3zlSuGtyqjNsi2jOsaeACVSV3
Sacq96WDAN13wOdbXQezYAaoh3H/um2q3K+E5d5nte4CDsgFVEgx5KsXtGB9DnJ2
+IcH9d6I+YJ2GMIg/IY+BW6eVXeWc5Tzzr0bwMUXF8603TSVdm+7MkRAc6ItSfWA
3gai+7sXMVAy/OTEgThpoTPop8XFilMX0yRursprJzHGQNd2BGA+pWOTZOuU0w+i
tq7nV49GGq1t6vzvOkZaL7nxPZkb6NQhfZcWnmpReKdJLu1pDY6MGPGbU6PupAfs
pB2PYtE/FHuy5skiihUIHBWNs+Rr5+GVXAZcBElg7if5foU/QIidBrqCBvk4A4Ye
XJYVeUHvyGcDlgfPTGFvwRB2Q4JBkRsV6yKfg+MEzx/zECNaXNYTxmtMXeW+fPwq
aDim5ikItV6X0w6sdOEU0OyPsliFNUvO1sQdJi3eUP2oBld2okUTLlD36p9r0VGn
h35OaaWwjSCbzb5zhRX3MqkSB9i5bpqvZramunmcmxEacxOdWcHlSrrfFd13vcQf
Zo/u/5wkcLYwbghmvlWSO24bWWOtsNyiG7AAl3C69wmKbSi1oBcveTFE/cfwM85y
JPdHZrEriclBu5qBhW1Da60LMbJKIyJ60Lvh7C3ZUZrRe8ahz2HZGxvEHGTc+IFa
VBowUcsphCLjZILPc5KVJ6Qse+bqTW+s5RPW2/NIkPDVAcY6wvNTuXaAoxDbsDki
nBPQ9Nf7RF7qIUBipNP6siHBa2/IMiODfQDlrofG8+b/wbv4A6+201QIsKhDUtyo
2VfIk64F5nXqYsJAViC/ByRRPvaRubf4SG1RTQTApVMKWoLkyo5InKZkk2L4Bnsc
+gDIekTjbuJoEtLqoTDkFfGvHynaPP61pMR+M/GT8ruzd5RamycMaB8L9FzTTfOa
cNKlz5auTViwWw8by1dz8GVPZ/W9k3NnuN6hEjWAK3jB0gZquWMm+xP11ycGBDNa
dKcpRvVfG3ESksh1z5I4a7zMwXdDGMiOcE8Z1jPrNwfIi7HDpvaVJ6uc3Wd225xl
Craf8G9wO4xmmAlv/VPBEZOZV8d5Z2ZP7smyA1XYH0ySseAKRx8p6T2lLq4csqGP
l6Yb6Mc6/1PqQ8vxCx3aDQNMW8D/9yZXt4fFxC2MlVco7JFqFb+/OmSyHpQrRhpW
L8mVNegXa8N19F2AbxRImREXwSKpW9XfDKUmWrtGKjuUl9p9p+rjL4sWkQrDLYyT
8xeuSBBVt5C5NoPLqnPTevnUnsBmoP0n72PpqECS76/FcRlf2Uol23SEuw04mJq1
wY6oQhDai5dBTl5H3JRIG4obholSzfwFs7Fxjy0rL+IKFSXRDHB5Pmjx4P3S7tnh
RBWcQMeck7XIfvMkQvettxoU6Fh7mnR7cjk/Ey9FlbviRLMK8fzcvB+r4Jx2+t84
XW3abjsPerLXck9qlQJBWI/cMU9OSdbr7fz2BNC29yYZ/oAu6hr84SMVlW/vDlf8
96ZBrlIpiL4UnnecElxUrxNji2I/VDuMgfLrG/qURNanO1j1vJI3S0pM8E7fmF/e
t95+oqdQ5A8dkOO8ne/4k8dpq1cBr0HH/QvOF2Oe0xsO+/pobMpZKP6wLzr6C2ok
zcI60sMVW3X6KfLNjRby5kEsQNI3LBkO+2eRM+p3ApulEahalgN10c8Oz9A5OxVT
psUVh5rYoMFOFKbxlQYLp69MBTzUD2zunB6UXgeribGlh7zdlnJD1MpmqxHIfEQC
E+shTa76l+5dxI0zE1XaCnzQShsnIDzo4u5ASTbUhNkCbwb0lCTFTwjNduvgQ/El
yEf/uGFwQ0ZoKf8KbXY27guMgPjV9At3FIjCDCVE2wZiaUJONhzmWTitOhTR6KJR
p/irHUqM9NEzwmsEepM1uIwet47AgEn3PaBuBg+4MFffnXncnWBbnk6aQRXm3BzN
dsH9/I8RByvfS+OY/JZn/FeSqwHkTvEFr1kzcOw0MUuQ7QM/ni2h9PpJon89YWGt
gwaTsSaNcSOvtViyjoHLjC+XpiZxrfjbIUM7Ikw4OCK7qcg3y1DX2LOFyU0/lt23
xO4gv0TGJgIGG9WP10RD7+1bnm9B7NrDI9nazH4hxTOsXe9udIRx5L8h4N06IxaG
G1+TEjWDx36a8bLfeernQyXDbzDP/RYlSH0Wogh3Cnxi4/q8+O7D0va8F5V7jraO
KkDC7EgatWXdT3s+qBxcdWBg973uXGBExBB1jzBS+rdnbwhR/hnmIHDPsEe6g6Ku
KEMqZkcDTkoNpDKh2O4xZwVkNkkCLhqb/v7x9JfkDShYfpmj7/+9KLKqb38qbn3y
AUPKH5YUjh6EhBYC0Vh6o/lfpVS1sbsQupEaqpXTUoaIsqcHYuBi8nPJui02bFF/
abJljtl9ael58hYOLhrVoIUYbHmDUvVBsc/WHJQT+FKwGzM2XunQa+XeNj7N/1D8
tnnowhmrycForoq6D0B3tTyFhDjd8YUp4tnQR+fMj1JkW89d25o61n0uwicslBxn
NSFtdiK3u87OBgq605aO8/HVrnS0JYjTACU71tg0uYI0PVrBW5rjrBXkw4GT+UVe
9rz9rLcxEFXSCD2lBt1gDtSX5YecqQ3AW8N0eUX4O5jDvLHbt3IhfzuNYRClFAGL
n7Y/9kofdSUNa5qVTVUV74QXI2HkQTQOWdxv7eUeBw6aWlmWP2ptTJ5WriiynZ3J
uvNhuixHAhBEmhef11PtEvnEt9/+YUdz5DB3/WeeeAiSm+sif+2xv016XG0AubyM
zSvHLei5shwyNb/3vP1iP+v4exlMQYudB9s8yJJZX6szkMwGBbz2Sk8W5J7yn18p
+tnzOQr+fklxcqJF9doHknORmZlfR+OIsK90J7ROim3E1lm6PBaZvJIxkN7in32N
xuGXyrOuDSiG7ODfGkt/KHvpJbB7dWRCSbYkQYkTVOqs9e8DqHFRYwLZSr1PbtSj
CMw1JUejFw3nH9g/FtzPVOQ8w/akXOk6/0h8HXkEpaWFLrJwFEknwoLLlBZ2dgOf
QhL57NkjyS+CkLbnoZAhRBakAtc/jUj+iR+aFqqw8lSrOOWolVdkop6gTjG67jWi
ECuPntXcImQkxKMYxoRlz0a2ApsgQcKWrpnfBNUrzBVInImfV4pF8hWVfWD8m3/x
G9QvYEKoNrfAfwXCuoZX1MOwfvgnIG1Q3T0ghJAb6kAONzsnwsrsjGo8Gfhtuxaz
2uEhshjxAW900WONq7UEqmZL8GEfPZuB2UI/F7CBW404Si2alRrMErT0CiUyIX0e
4G6vXsI7sE/O3JbxjsgenIYZWD7hcuoRDMIwqnxk1CtsDClYdd2VwoomevS50Kqw
6s9UEeGMSLYfLB5jOcGQ3p8F2YiRuV8Gn86Iu4VqlgUe4pDkVUhKjAxbXADkBNFt
BoxOIstSxX8adS84G8d/AE6TLxOz0EvIVBY5UFBHZfGUEqDu+3STI5nqtorskYMF
ee9m9wU13xeD+Uc0MUchahmxiSfzc04OcH4GXNqDZDevRTHPYEIqI7vXNKd/VD3F
CqziqaLIYG2Zkt9KLh7iTD73WoIqwFnc36bnMC8LhvpiRDo7C9T1a+ONCDdMXYSP
fSGUtyNCx8xAybWzVOjP+tDO1uEvr/6EHh+8OLUd//lu09s7mj+nDJEcKfS6qHdu
uQrCakyw/OGEfUOR7g8dHXxzr3IsGbm3VCYk/93OU4wrAiKfkguFOoVmIPm+ZDyG
u8VQ9dUhHLRQn3V8fUhCULTyHk5wLPWreHu3kp+PFxQM932MfjE0YItPT6ZZ8bMA
WQ87STSuuckpjsdf7mADGAOvrKyTz1WdvgaibLpOnuwSGf2avYrfeiCDJH2Bbeqr
anixNYf/7cHuH0o18Try6HmmeBByZeOymToHz8jcYSM+jtHHXYJRBmR6mQSZ9Cn4
PrvwqCxs9ce3W401TJMXuq3FLuv5zUk78bxMAYKoBlwXzg1Xy8Tw5vnS1/C5QjGd
vagLdO9K41WyJgFE5RVNTeQ5p5GIe0+24jZQHLGMr3sdo77mRCne9OScdN+qAk9U
61pl5J9VV+wsYF0VpFMUo1cx3PKiTmRJu7BRChkUtTbujevMSP/U37lktXLaebmP
KOpHjTtEWso58CSrwZ2kjtwQ0td/82ANY5/1wSvONpUZGzCpMmsfK/TJIBOsDyZY
7QFyxuWNi0YtgK06a96afpl8jCj+90PGVpJzQJ2wBdC7bkHFCzQ1P4+PBxMkhYsL
sabXJ+E13QO8iqBeJ4CP5sNKzEk+L/+B0ucjCTshDOwwAoX1UPmE6h8I1Lw2yP/+
yblvicGiabQA5X5BIN5ty/c0qKFCFlseUXZ/xo766zLeXjGW6HFa30LL1IC3V38A
U1ajzQLjlraQe5DwhlwbjVbJzM3OyJzwXwl1pzL8nXDbd73vJy0N6wzBdOWlidwf
luWADKwBjSAS6XTm3r9iTdk5g3XGXCGr0ILXzz2yMdvm/v+FYftF+F6OLvePJ4ja
kUIr4bfl/ktTlSEv3XF2rklFvipUyulWbdWQXJ1cZDDgmkNCl34PVdShfjtv+JW2
J2dPwU2M7zmSLPd7ETjaztI1l83NEnvvFIQWMzTqdp1FZq3svqUmWgzjzZdcu6fM
rgPKEId9XHxDMHil974I0BTq+ImGFsmAkvgKJQ1yHFh3hZx9g0Sz/3TE0m1Wi7TY
Hk37/UYxmCkMTqKkW4s2fzEDjCDsAKFoeinA5UE9kymrMvfA5iV62ilIHmm986IE
HDaOb660ULyRmngMjgV5YnCDz4cf8KIERZcuMLyoeXQvqrQWhgjVDUhmXdMBFLoA
wowwGV/FwOQsXAY91RVkgxxCVa84NXUALyL/mqAW37NMhMPmKxNJzM2JxHeHF7Fl
OkbqZC/gvyLdK426rJWTghdijN7eDjlHb9/BzWl7WJQjdM0eLlvvsMzN8tbdJgbX
CilR+n9UchBObluzpB80P3i5sslWEIZdNUJpZXrwS2456j+UVZNiK5JwwNyV3D4i
QTgeVI1vVlXKG1yQmYgfS4i1DusfP8FwksNmTPaj/QYZUxFtolvfGvYeQc+kP9IY
3PPgtl6gtOljwkIkvR69+CfSOJvUQN7ZDOtVCK4an1nHHYcWKFgsxPVJtAC094Lo
7mIF/UzwkgQUMF0nvqMxiEatitDpS+enfxb019un56xe5Gunrwdk/rJyqWQh2rTW
Xz0LsMIUMETf0nn4YiBWvaA2akcIBbVwALXM7rMoP3GXfDV0otuJVBkQgCJthkQZ
BG2Dn6SVjL9uHGao9LcK95BMzONLk6DiVqmM5RC73EbIht0LkYyyERpi4ZSaWljW
NONZS+C5RHElB8gx5DTpcrUlugBiQKC4ktfqvxkjCxULe/tEtJ03Tguv85AIIZsF
7JcoD8yQT0HdzVv5dRAEM8nQsF2GkjyrtYrrAKCWwMuVglwrP14jeMz5ivsT7qDT
T0UfNZxnMXV0jRoGkhxLAXYwTk+pU98suHyZABhjkPrElqYQXgyoxl845BdtHYwZ
a9ICj26zzJHV0AWm2bp3XwjiPEF+XOYv+5fyE+/y1dT6Fqd/rR0gXmy772o2hkYk
HpzbdfZs5oj3aNb6ZooAu4+PwVosjbyN7Sh37rNN2JbZlvBI7xVrlS6fEXELZmCM
Ktl5veCY42zp/6KaIy80mNpi0G7CyeaL97qzR6sdLp7uPgCgg0+jsIxBP3OJnK7d
VWl4vZ8xgQ3dan6YcFtktP7mW5Gsu5f4ShzSGGdbkUz+ODJNf48dpZ3HAoMFcTBB
HVI1gXDJ1LkvgNATHk1J9lh83OSIhnHmoqT1h3XMyoMCjxj/E3Be4Z7N26ZmFtMX
dPWCxaIa+SSk0Lzk3J2/xDQFhFQjz5KoN5KgoyasSsq2dd0wO3t/Bdz2cwziiFiX
oN187O3dxFcXciIA2RCzxQBzgyAQgs3MIdyOCIARuFp05xpGAVk0MA58+LaGMzvf
MsfTmiCUvQNBWtIAIyPKvT2Q2Mpz/fE0JTR46Bfw5lqIkoFg2gm5dZ3cjD9BPWjf
L58KkbLyrBnFdlcuLd9UFI4hOw23D6mLKD9KJ7FzriEJbf44yh+fTlKOCtqzZPO9
cY1nR2LCHLKrjoCRnkC/0WhxCvtf1DmyOffcApilDJNduB5oqc87wig7bemWUDNV
atN5qqMZoyXDW5wJK8GIy1SVuJVqv/PWtnxk8WC1VBQ2Emki/r3xAdtaEc0aeTzz
NX5DAtVTDu6o4RurDWB0B1BYIJqabWiLrO/0EdTppX+SvGG3orz4cI4wL1s7NiHY
1OGV9v2Bkn0IA1JXxGZJLjPsDeptEDgRflel85FPToZgRYoFcvVJims00TD1Zx5C
Va1k73jRGJtr4y5zBx/x7xAGxm2upukiM8JF+Iu6VCPz7pLmUohSh80bx3QFz8WJ
jrodWpknpJR7Y9s3BfcQUjVFcTdzCUN9WsWNLAVUeeVYg+xwwRAutJvhCWBsW4ro
66HF6FqLkutsFK541AGxjQ4uGsZTS0CWaTQb7EdHwOwxhS2+27JsKpTW2zuqB0Yg
bm4rvKearUHzZn+oaIQASWkxgxEJBqMMXK2n6P730p+FZGgGvXl2b3RYKKlWcpJZ
MRjiu2R8FM5z3bIJ2W7QH8aDZSZEPnfm0HN2jJYEFHQgK1dj+jq9fkjGAak1UARB
vodtmuu1PU1VAnP/ZfHbn0XUjIhqKcXxzytw9FxdHXrcaxN8/Bb3PPp+msr+qBpQ
1tJd5I2+YVoXQd4FXp9ODu3qWl3XCdokE4SbTrxaZEFEyTA/JciiKQcYAZUbrUAg
3lRy96HjfknfaJtRFVlMisgpNHF56+63ZyQ9UifwaP5bVV6M5uGwkMAOP8ct6ZP4
sog5GZkFf2YiSBYanVx2l+073Yki6m4X2OToHsYCGtHYeVdtwmwh12zK85bxdN0L
UOCmNC8EqgOlRoT7eRI84bkT9faDKFCMMzLtdwh1Ig5pIBIBhQyKdfNJdhOfD8BG
CCIYg37M1cpj6vBV3lCjlvYt8sUMjEW3L/L2AeDXqjoiRAulZI9vN5GTONiMwb71
tcWZkMNl1fLSnoXG6jM+7GRd9v+pmZKdtRgr9NDasZEVs81cvuRlpfDtJsy5rMkw
7JiwedsUrYn6jvBDV/CNrePgrIGSTY2Keoc8UAqQOiJd3X2rvEmlY33mFx3wdAAs
zHGGv54tBbceH5ggEYzDnTDXPHlrG8HXBiNwM9IAFt/bpcvnTpBAJKPWsNzVPMt2
kX/4MwBhb8wY0otW6YQpA3fK5h6pRgMw5gR82C4m3hQ/HqKeZuYye/nu8Kzo3SUn
TFlGqfRjJLE9SyF++XGanJHrIsHzQBrXmmAU1W5nYtbel1QeELaHKuEAiJ+/Zy/Y
IBDiCczUlaJ1d/cTPeFsElf5pugCQOMqls1yIvYxrproYMZX6vgebZ1olE8jJMtP
4X4bZrmA+xr/NOigxpUseMSsqdto4VhuAWpJ3OYtAEeV2kpXz+GauB5tG1ttGBo2
fxKp6teiJgKz1VeeLPQAX6isv4ECO+8TcyntHpfx/j+V7Qv2RnTTvuaCPxwKqSgY
BEs9K4+n9ZMLXe3YT7445zltMKZIdcFAEPyRKPs+2PlQRo/qgeh5KIR8tR0lUScE
22/mTDqnKX0sLMqwDMyaJIuj1JdA+wmtUvLq9LyVnY/CMsV4Q2s28+5c0hpPXBLj
LtY4KpLrTiTaIkLdld624h9ZlOuMaNPu7dzijvyMAgtTY7kcJVXu83Hf7x2/zD3M
WrLyJYX4rT1ahxDBShKrqdc49rC1aJd2wSg/9+lbfuNVXP/56Baghqez9UAx7lZE
nzSie9kLNsn6O2PtsDCEKT7dextzeY+qPeT2SWt2q8hW7HVRzBYWySxrIhYYa1tu
wOKShR13LFy4nFLpPBBkUk108yN34KECZm90R214pJ4s7dJzB+eEh7ygQDT5YFbu
szNbPiO25RQNRZ2mjxKv9H4Cfvo2CKd5nPzbuPAjYAeDTJt/yO7jub2g+aJy5TKZ
WjFV98o9EX8DwTxlCjLFiEzU9uGhCvEE0FpVsGrxw2thHFS1OW3jTABcP+/HPin3
j6GeQ58UzxnDTRWOPmv2yLwHcGS2oDS6ucROU9gGSZ0BCPmIIWpBRSZpawKRYe/A
HrCQqyZyPU7WVA+1sCDyf+q+R89LTnQL1rOvQNpvjOXSVjmGHzhdwejP6CfdM/GT
XnFfqn0QIUS0w2r8QqYtVUluchXc1zdT0K2YhsIbVGHcfK7h8hu0ISB/wW2zzP1S
uzwJ7rDlblFvVS9QsoQ2nSTGvNm5lf49wj8bdm9Cx1t3woHJdw2s1eyHIchGFeiD
3PCxyaR7FUc486Ndp1T90ma1IXP+B8CE4HlVVe0zauZB2r8pmXSD6syLbOrs6oDf
Lnq67W/sudKwa4yrEe/BSsJJZ3pLdpu1al0rxP449eRdQiCHC3fc3z/0LOTBChHI
GpO6ikhEpd0tcVTDK3ZY5DXbMro7j8Y5WxFrNZlKBLwJJIzTmZUF70AyQk9xRi+B
bKwOMTn68VKEcGd9XQOsf7lwF7H6KJ2mUQ4xU1mqPt1NKa102YJHSM6iaI11bxF3
pZvrtGRd+TBaWito39S5u09VwsC90ILlT8fko1DWHYAqt3Y0pPTm0hI90btUzl5Y
WNwoeMd2XZSTS/C58Iblh5UCd6Ly4z5rpjNUSCLTLavqvnJUddwnosftyEBF0DdV
fePbxcXBZH7AxHpjA+/FjAhcPrgbRshYx9SdgiYYmS/HZP4pJgPje3IDH9nRA/Zz
Wd6t62AOMBE4Vg3UMr9wkTpZU1fDqnt9cugzyDr699qS0SM/LGotWy3+/eqE3KKT
lbXDGgil/VgeOhv/64x88Yvb9mCV4ZGzqZ3vTlNlO4Ye9ACAm9QbJfVG7O5Pb2BJ
+/h6K+nELMqU86AHGTYYEdqCXauMYFvhnVEE4FajfK3Mxe4WvDbGShztNzNG5T9J
yZcvDH1Z4zrcpRca5anVWHP3M81rWlPnzNoZRFIPcQ3FcnX3Uj0FTT0Uvl/tGyGB
HlKn2su/5TcT86MEvE1GKQW3VOAST1ZBJ4Jt+VUyTpQEpGheFH4TJSWi8SY4u91Q
70cUVP3MEbjBPaUkPLO0gRIj0AHNsJ/MRXbVaE6KO82HnK0p4A2DymfrgQzVKQE/
3qtbVMfslo170zjCi0U8PcyDCIE3+nm9TMzNOYIB3c4HxDoLOKMFpjtJ6GAQi72l
LBH34qEz6Wbey6LQn70hIi7d9yxK3vOzdbJhOEEB9EW/qIGR1uBZ1WXPeydgpCsf
h3oPYDBRIda30ozoHiX6jZIJ7iRkDIolXByL6Ou5wgsanBQAa8hDKhqvY6e2a46n
4mUDI/GX/CvW9htc3c9x39+l4ec8fKdHDhU0xTiVyzj8kgllhPjmwbumjBmpomik
W684MMkqCTa1ugjAg2MTtODSs11RK/J9KlMxGDveGLULCbNDi86o034O3fIkRiN/
odAA6pWnkwvI/oyGJgsu+54UU3ZcUq/03SICqr28J3luWiwsKtpg0YbHOedRVVoy
S9oJDG0kjoOuuIuwG7HpBFChtToEGMS1qmN+Uz7t2WUHZMx55x4PRDgBNyeRohAa
60qJitnSwHHDzKiB+xr6VPD+SlmKZ6aMYOqsqnp/OGfN8D1Exa42zTja+/JgWxqd
Y2OqxZBcvqdsC5UwH0Dm2l6V3ma/TI6rgI53kl6uDyTiMIj74Q2OfE7eTuUxyi1K
R6gbvlWbfRLj2sKlyCtIr38zk4TQIDa+BAmFBHZi/wS+z2t5r2beE96OJjrF2dMu
c+22T1pax+yWNLMZm88CCT7C3kU5YOyvwXbsfRUNLtydvQGgMjACJAXe/kmWtmHG
mz7QPCwm/EBtkXwPePaIpDM4BvuYD5vwFHT+klyjiGT8ULO4fMY83fX+HT9jvfbK
RpsHOVXm/LE25Xcv1IsxMA0zhFcNC9Uuftmmxvjc7aJQSQ/ZtwCbqU1kcy6128gX
AEGDVYHcvWytI+GM8pWi93/TthGJMAK5V3qmIYaNvo/tydyyQncQ+vHONtqCiH4W
zpA0+2qDhZ5FFTfI4L9mumAHGIcroqIFAFrmBG4IWsm9HNjIKC+GjH+1dHJVSPC6
6bTkeTa7zPznNkTyPDtmHI9Lx9w8ljl/wdvj7XyQpv9Mkpvo+YsKMkDHVsryHeJh
7rr5gsgixvEvHrvEIDFg4y9xQyh+MllxKLY+18QJM8jHhCmMAIBXMJOyyfF9d9j8
kHJoOk31PGGKgPvO3pKWdKHAfcE50SwXH6Sp7LM1CW9p9yXwLDos8Z2jtnksfVf1
oBOHbH6x3PED8LiA2dWx5w97yBJMd/0oN4YHegcirfLLp9ZIbAUcqEhi0IU7Vnp5
DjVVwY4JObCf6Pb0JNmyTxlA3QSM57K3+M9ZOy+PydlHLoGa87HnjC2qFWbMC48b
f8etHee1y+ltUwmFlhL7IIrcC7q8bONGtjqBqT65t7Cf923+HUtnTilRqJoSnrry
7bx5QPz5YfqHiMEnk6co9KCkasb1AOaGk9ZrSp56h97c0kuas7/YbG42yW/u5Dp0
E2/YaBux2fEaq6AKPmc2txzvQC8X2FLks/acUAQB75//DeZX8sF4X1eM+6d3PJW8
j25mPqHvqk2Lr+faYcL61rzoN08aUUj0rzZsn4UkAdXpYLG+qb7A9I/8pZbiGPLA
jkBKdsywL7QcVFbsFfMbzVpwhtga3YCyOrejDNXITxn5unCgrEFcD9iQciCRLMn2
CfPWhKp57qeeLoRIPMMG87amqRB/fi84FW0sK5/KV16ZtqLiF+SOvx7oNUOsBFL9
7dbPuIqcaJ+N/EhloaQFZUai0/PEoGQTOv0KbhGbc/ZKhx2NCku19F1fYysFH/SU
Us6hzOx87c8ACWD8hY+5MfTmSkW8AzAoVKHtezh6J+CUYWqbrQEj6l3tMAdmkOyw
Wesjy7w84fqfHfYJUVTQWAcUhXcWh6Z9pa1361rfXZeWXtYVfMzvjV+qq/GZONfQ
ablguREXT5yMWKKbefDjoKeSN53H8b+GfaM73csp+7mHq5QENw41ARPRHp/2HzZU
hsaJp4pdDYNI8iK02vX9ffaTlI7qKNmO8WCMadCLirLt1Bg7D2yRc8gC3KiIdvhB
wedrof/MtKuqHMeAhnh2NJAsHjTizayWdjwswZIe0PLohvPh6errILZCpXsGAdR9
5ej6ZN+3UmrXJ8xbogacOShUXz6aGCo1Np/iIJom7vLP8rccVF2Q5lAYjcrOEcS0
b0zIDxd75Q2Bd7NR3ERaKurFejQ+uLi/pfz8MGt0N69xqNa4i9j1Zce3sM8lO4+W
jHEkDog3GlWw71R/RM5L/CVMo2grbQtld0MfBCq9O59AO+CBODZI6BfXrxyXzLYG
+2sMRmGji6fjHF61uPcuiFZKDPH+wSOsHU9n3SBbkQ5hHgtMFJGaMg9W0r6ezNOV
CsvtkphqsyrgCOwjlLd32/ui5+2bFTRlNX5OvDnfBa9aEupmeOau7FnOhhT7WNeT
RaIIkfIVSw7M4fd9bxRP8bqtemRT7IFnmqku8v7QaoiigqCWLerIvorPHqS33OlZ
8RRLXzeocda62UzPQDX4fAbfJ8saeovDsr5PS7MNIs/kk4Yg6qKtOJWRAxSpYH23
SUA2s0vzg6/gtKfTwtFeE8aZWd7UKcWKYNFE4VHvEtKywDGzoWStxRBC1QY1EY7b
lNRInK6EooNZ2ijp/xzAi8bIX53znJnt0bvwIrK47bjf+vOS7FuDASDKrc8jwgGV
iZoq6m+aHmRVyx/u5tjfQhwwPLLmsYrkxiMwdAdT2Y12UW1YN0JyZ9tvqpxtAWlD
8MrzIX35sN1uLc7G4OeeAI4AzR02LKSGyriieLY0YKvsacK1koWQWpL2UAN4XASo
I6OE7T5EEwFyQGrTFVZO8N5x6g47qw9zmU+DTloa0SgL6xgmP753wbxWJGlbkF3w
jvu9DOmXv5kS7e5KECbbBeSlsMQsy0BUWFZMUduo6T1RcrqcwymArHrl+hskRAA8
4rN3bFeSY/OVS4ey4fCu55fFkOASX9XbS/g1hbnewXYEdkBWwChz+wQ8bn3N/5v6
QzmgB3S8KZ4ajrbdOb+vaNUxCb34aI09i0bGnI5yYIaSJSy0mgZr3y8YsorbHbZy
j8TkXnxuuxXyBHPSzeTy239zrJ02MPpUI7si8QxVcDe/YP/SyXSFQwCU1WFJV+aR
OqFywMEjgS/J/SJ2ed7BPzn3wezhLGSczQp6dj3LUpvmOXV3nAHUuA8nRAlkGqpA
1IbHLDXWdILfkBV7AFY+1YVTUNR9MN+QzJGDMRA0OyN55olX0wKK5jWeh3EaJT4+
zXw2hcLVVbBAKfgXToQgmC34DZao+g/Jg2mdoatpopyHDlA6QtTwdXew2pQ1TNo1
a0DTsMKQ27ogVwteKIjiPITij4dqGRBipFjz0SKnOg7K8H/EGjiepc10AnSh3xga
y0mm1TFNQhFtfUijBZ2jLa2BRDDFJ5HOkbnNkL/qr3aKF7Gl60H5qccwxm2xCu1u
awekeuT6c4dH4ZfS5HEs6TnHpdgJtmLtk3/c2JhhqXr3+Kz+pKViV1xxmvh0mOM5
ja1N4hTijgoAJaIEO6yxBxfAT28D14ergnR5d0ympcpTM2bjXd11Sghm68h2oKqh
eYv6Ft0Tes/Kk0hoPVakV+CpHvN8JXxIE/FsEDaxQnLBise99oE3YFZJH3BI7y/0
DeOk8WGB0n0Oe4bPxCK31zw7A6Mk1fQX0r1TViN9Vgt/Jn+dAzZ6Uwnfg7iB0+91
YGogn8Zmm5XH6cKdEfScG4zcpq1EGrJKy7eLJvzf/JSDtx4f2/fWiebLefDpmr1Z
fGw13z54VZW5KVZzCw28p53tHcGf0XP6Bs+Wvblss/zH1abm4H/fKWPn6FXB73Sm
SxsZJIBrOJvxSqF01TW+T02jZwx30Dkg78d1cz4rgTqc/dPt0mFIpdGPm9WvbAlU
iy9BDko8/oUmv4ViVbUedP+8ZhsE2FgtNx4wJGiBHzRzb216uv5dbpDmgbVero0I
t3ICRxrnx17ubc2Mx0L38H0SwqXahqD/PvUHUTD2e9RGDq6Yu28wnFP/Ebo6l+n5
GsuhSamdRNagRzwi1lcQ8EQ6+Nn9PCRlQSi0vfs1SmL/cPs2FP6bEKAUhTfDCwZe
aLPpccWZLHjqaPON8/ryvICPNhUkqumlfvBb73gqAbhYKZIpdNAA4hVlXOywbepc
AVM+y/qF8j7zIaiWz9jQ40oDvtgIMGtAJVdKcw5u4TlW0JIMY8jFpv5QZo5KHprP
hnpe1qnzb+y5jEG8gG3tP1w7yhUw1pugbDXgpmnL+HN8ZNHrpkr7RrOg5GSh2cYM
CpbyEXF+RKbBcsBpDQEM8OP4i16S6M4vW9PsVHNhMxn7Mk6YEkVSeFOnWmTdTocm
VDRGCGRxthrtMC1iSBUoi48c7ZARiH4LWuduUI9W0ndkukNuL/C7QEI682jpobWp
8IKZqIYpt0pnOLZaOizKEMOW4kpHpNpaB1EpJFZQeVv7Ki67tJqM6g5QnKc/EpWv
W346JuVmNvygiNa3IdoAsWd/ed6fYvvbZt9gjaYqBUJiwJznT5dUxhkkxTqVrCaI
Di2fBfFirGI5fuk2qaG5oAXxdtUCd59g4/6X6DSIKE6EHXJogcXPdod57LYAziXE
zkwwFkQFrsNY5DvIEu072XGhH4MWFRveY2NknS4eQibRUiQ2erWvxQriAWhY0eoP
oOLHSHuU6jpJ68sGKD7R1y0KsmPKQOGbZarwBBTCY1xcK81nzrOHxQfSvlaEbvQv
Nkc3d9AOwnU3FcEcLY1YWDj5z5KOijsfXqsQfa+zYBXGf8/tc2OMvr9waHOVSHTQ
cuzgB0OBdnc3/xPOWefBPsnFURdKkfu8vCUonkK+sgODT8+LDpyGl7z+BjR3Ehqb
A8VVVJSl5rphgXLz/VdJd6RTuQFdD4B8fYKPmLO5GQPfK2T2rbOgu9J5LtTaTQD3
DBD0QLtQ/tTK2XMbIrAesG2wPoMsOeZjgLgqKaG2dRE8oLy4AZMKOz8ypFiyCrxQ
KGFLWvewcJi3GrQRDbtlrBbtZaTmC2pUi/fJyETyUkX8yMwaqlIXDcBPky3BHgaI
+WGnfYN0RUpJyVdqOMW5rG9+01dHgqlR9wsq8qEGjtF27nD0sohcfkhZhfk5VGA8
sM4umvHoD/4QlrTj89ciKMhqFSPOcP2FVgh/Qv3UXNKnZ+bRY2XE3hAJnZVpeKMj
ncI93apNe1jILsZsY765w2ckTx6g1TGHIgFefWX+d4UO1AUXjzvnWx35VE6DJXH1
EAXYy1TKE2VUxGCrlo2iO7XVP4tSv3lsj4Ue/TUFrd3203kHmfwW/WzaQWQdC8Lz
m7oaLuNjV9GzIwszZy+vGSKkZax3STn2URcRDwJaJIwLzh/sVUtQ7FL0yxhvInDh
nmZXkORGK62qhY3i4+kohZ/oPYxP2WyB1BU5d6DBriWxch3bhc2p+ReAMQwsK//H
fqDALLte1r6MBJMwArZZm5U8gxKRfJwf1oikgGmVyp6pDGEWvvCXrfMmzt/7II4t
paC5oEytXLZmbJuEMaBASZb9yY7AeNpCj9dHZ5OTBeN+N09VkmjKT9X2tJpHTTsG
BsC75D9JgBJLvjzLmTQXtOdXFpinsJh1DPfo3abtP2I6lxXyZsaVa/CiM4xf+GMr
7AzisxBAuYdrXAidRH2xgNttYgBoZpHe9YIsTcpMKaGNLooMaAyct3xlDp9/Aw8E
Q5I8fIXHOIzPvEUkQNWGhImtwl2ybZh4dItMECuFauYXs+E1nrWhNDAYGIPSWP7Y
v/n+uqkE9POaE4fOvhVFg6cDK8Hj5XKtA2uL3kJRcuk+FcG/PvsuZXQTkLcZN6D/
8na+ZM5RIs7VtM7AP46VW3n9Z8N7RHu7ztnMl6raR1KsKUa1TJqoArI/7Xv3b/i6
JsA7bBpX7x3ebO+p0hfr33iHF+heZSN8BCblvKTmsCt1psoO3iUxcXsuLBFNqYnV
ieJf9Dph0O7hRHGUf6JTuhSw7NwXryYj4ipqeyZIPJZYBaDbGIPVjdcpEezNC/Or
8AEc2wFu2aFwP4itwd2Xtuf0tlNGyfFeP3JAgi9m78yKTLvuXIWa8ydiOUQdWp2x
oByphf+BwnhwshnTomBJas33iy5iIeaRRk30hzz6OF3/2i3t+cuYxU2PCEfbJ5D0
GJpArtvNSH+QGZ5WHn/IpEn/+qKXD71PVW9FRpukrwPz4FDf1acH4hxqc55RxuNX
H2oZV5c+YgIsBj5YlNs20uzWmesekv2tHvkI9zUBGc46S1+LnbpF0UtIamF4DJsf
b5QKGgZRqGjt/6bA/MGY77P41wohSaGpJVYqlM3AILJe9YkG+RspyUCxejCJEM+K
99oL21qHlp2AuKsT7vogzwifa5oafSFyV4jTByIqUC25+qrexO32D3iZ6G3RpZqo
pHWJSAuuEuJFhFr8RKRVCD+M2rRfDJK87xpAPdbBtIodIuxfKHblCc2rIuG7udJN
xcO5HNmWusLpo0PH1eqkh8MuvlyazaMFhUV7l4GeRQjtFDfQMyKUHV8kY+jNvl11
pQ8JSBqw1g19eSvrSrOFDxBA2X9eTlE9PMASgAurM79D9LA/hy4AlnUvhABno88E
BZ7xw4m3KJEr/ihgt2E0uUZ8ftQd7AAxJxGyWVzXRkjJ2SLB5nfiIUFV8oj4wGKx
w9BW+L8dr1BOYsXSA+buYeHXJvcUwkOxzRfpSE6XYBx7dUVzHAnZPU9eihAVcNe+
HooHuFY4PS8agcPg41cCarszqU5tSj76ENiPZdfCG779dMh8j/aEALtv/1ohrWiL
/yRmWMLewU6i76AJ3fQJB/Yad/9zYjhTYSaNb7LXBiUV2rFNS/7651pyMLJ+aeW6
OtfgI6LFLAKqrTuSUlbQI4BAlBVuOtvlOttjnO7G1JRoKrCf2DdTzKLDYtjlPZQP
16LcaEu12yKggnYHbZSLyNgqqRqx4dFDw3Vf1LDSgOe01ANrXaKsNn4AT8YCet55
3jJos5b0OF6PrNz0L139SpslmziEIlq2j4dTuqb7zCPqcCxQQrLNsdJw13+Uq5UH
vzllt5VSIl4vbu2ek1E2Q2WWHncUXedyJqDyEIbHwNmecHkfp+9eh6lNJi27aBJi
9M2RF8F54skpto7Zq26EarxZirvsgG4TP2adHeGWy8uGC2Y5CSWsikOKZ0XdE2Hw
3uyfYQfN3oII9u6LW0iikw9xRckbCNvbUdOuqsR9hFmI+3YwYHBHdSHesxJrl6Py
tU5q1EgNGdsTdj5w7fjBtZTa+Evw3cb/aukDzV8GQJHZTbxT7H3lvwscRr3T1TU/
jpBvQ7DxD/L1onsgzbmS3nQD30EkFSlWku0DO3GAjszkVmVi8piv3zwrROywdCrv
6RvDIwcCrQQ+zcZGalwuujSgTsxnW3OEYrCvPO7RsLya3bv/aFd8NJQnaJhKzdco
7Qz1tAKgHWWHaMUex7PAftZo0yJSf2A/FJJPSzsul08pETM3ygKGJxpU+xXLDq/A
CT6P/kdocvhIX9eb0urgeB7tSVhJ+YlSgWoabD1YjVy+LaRb6QRYldXqXnY1DxNZ
FfEGSY8xgAhrK8ejbDD8P9CJCHO+T6FCSwe6zm2dINmQ8DgFZJpozhmAR+9eJLmo
mKOb7SlF5sNKJZpIfnNTe8rzl6Vty1YzRqEdsRLXeBdSPlwYH2fNdG1ALWuKVQRr
Ck8Qoc2VHCOIZUnogQmq46KGyjHenjSzLzDNbhAZtawCV5m6IqtmYbwoUc+6cxpV
N8pOreom7TfkuQ+Yfs6VFjQokxk4kXA25a9OQYV+ZnoRkL2xddI8nHDUBEgsyGtI
eGvos/zITJbXSiqb5lNuhqoh327IT3YFnlGnASl0ClnMY5Do9Cz3wMvdKE0o8Ber
K34pOCI2FkCnnjiOXjDr1M9ijdnJfhc1GJO23Hzk4YSo4H+BKshOA1jXYtdjDntD
l7xwxfjl7BoT496uSv8iEGzkJismQaeaqzo7Utf79UxZcztGIem2Xwo3K10jQT0w
bGwmexmP6YHEGR51pTOFtySmd/Ydd/c4J8ISDU7Rz4NehPqjTr21IRNC6xr9z8KG
84d7XMQ0nW0jT3KtWRlsUwrQfrChzBH+HNKrVaNhJjKZzTP/qBqX4c8D6G3AZVu5
WsYTt05XmhxE/AGcFBkCC/TZKWcqXQhe2hp4HZ7HYmScl5sh56Vhjb4OsEMpgVYT
OEjL/3EKtKufeIVIGTPBze7rE/cUL9edmzvHFcapAlVF9KbaTqSBjLBQ1nkvMvRv
DkZonzEs1ybfBvZo+g3ttyathCdet56IlzkzFMpaZt7DcHSiq4qq/co9jXJDTRvH
XrvGTZm4Q6J36q8u7jjIgCeIp3G9i+GeGvNylH8spIYUM+gqvI7S20bJTKTfOdT2
MrFsqnozc4eN2oeMXYW3+iR9C+278QWVQKfcG8rJ9A06SdcFyJHGZlze5hW2R31K
OeFPinPL2n4YJxxM4oUJbpQhl+75KbH2qP9ge7/5OOr2asP9fMeKJeDwGIjBpvM+
fGvyJ2pOrakoniwk0bhNgT9zSB4Pfa7tGbTiY0X3vDzUon+bCxb5DrPeNa19/QJw
HPeX7mfgWuD66ZVhG6yh6RnhZgVCHIVkBrt+3Ks1pkTopBJakz15rdestMo+3AnY
Q4NyW94tEIru6KipCUU2j07q0PgQ3Ou26Svy2M8jvqojH8sIoX3gSDbfRvD6YBzr
bw1f6z+Ntkg30Nlk6yqeQkyKZerzDGitaPItrrrxFYtBVAbJtwyP67YwN6tlyHCn
QQtZ+UZlF/W/JdiYLqamCkIgolvqzK9OF2wbDkhbmZ/WU8vp9OuhHiF5llEogSDB
wErAFOI+rPIfgnNJ9GCeMSzUl77gpveROEdlPXIgUWqC8KYfv4+4ykcZ6TinFouf
TVmGj3ma7qImdZeHBcK0kWxjbQ5qRFZooh+KPSpMwKeG4ygwDTtNoNsoxT5Cfy20
YsXfdFyuUGWVEYMiAy5khA9O5Z+mFUy7ihvNX9zy9Ydu7IV62ZUjExRFKrMiN3iM
eYXwcjrdbhO0Qk1Qj+QxQcQqlscshkMFMWntXFEJqnelHUbvCbNx7ddtEFQIIha4
ozD7GHc44eci1poOzJ5tyyOIkQLVlJfMiZsDEegUf4Gom79dQ4sOGodplnFVMt70
plGqVKgAHS9ll3ZdwZt7iOHGubBVfNtTf1Nr9U4AEazPaaFk1ZUDDpX2vedMlgbn
vgl5fnvwv3knAgMvx84jaroJZTHIzINOBOqh8ac/xEJxki4e9eXAcVCXBQFzG5ab
zPBpTnFqtqOr92YNO4WMkZ4OYQrZ9hYQ4GM/jWKuktNhanTzc1sPIkqZnfCMNOBf
ZgggCSHy0A/m3ldyJAupbgXCgJmOa9apuN0KfM1d6jcKf5ADnBY47z01xljNQZOt
/yDUqbZ1495BwkYRKk2d6zGwXFsMyRij9AT+jgblFPa58ec0TwbHL1y7OhhuNrfz
DXU5VybYQrnOhz005SoetO1l2B4jDcODRT8LAVDoxx32fFxYLjoD5ZwJbM0VSlZy
KqPQ0E6Ed04z4rJzcvlCT4mwG8i9I45bTdeu7qJaa90N5CF3vgd/lz+NAeEBRcLT
L0BAcQXEDeOuTzeHaDSwPKc1vb5kisxEWZJ0v7npLzpex5nYfj6SubTgNQdannrC
SDgYzAJBfis/O40/4c54l3bXatozxpStQ9+SZ9tP3Qqz+7MwVPWx9zLhlQ/tnF2E
F+OVjAFFIEl0gV6jB0lu/yvwCml7OxAnLefTtmrsc6/tbbY3/szaSY79NsZw9JUd
B+jXN4BIz2AVr+AvQncInKjsK4r0utgOT5nuWQVjKEWE4LTxgxFi4bb3u7JeASeI
Q0UdjapUx91tB//u+5VyfOcc6PcZRGO8EZS+eqTUbdnOIbtiKtAKwPRN5qoDW3jK
a84nmBx93WhIXKJyeSbqA2EoxI2pIXl0WnljtCYBdHJYA44gd9XEuh7D5NfVT9wu
esKszFPitWvZ4oaCSBEdBXyicVqCB9Je72oRgddOPoVljIKv750o4DL1HE+igoYa
TTVfVW6/fl6owZAd1az+LcVQGvOghxXTBVn4Bdxm2Ip66lmTrJpnFP2tdaeEsHME
X2wHpY2bVOhigRHpPoiO8SeCT1zDQ47oqyimEQTRxKbUpyaZcPPyuKHkjZnyViG3
kHyIGEo/PPYPvPU7yOw/cR1rMGJ4NZyKF8xhUQ97FSU3bjnZUVVYCccTNXwzSahv
IRvtNW14XYMGkSivcWD6iGCgEvk+38xb5gZOeEEh9/U1SIK/lgQBnfF8Xgb2TcYE
aQTmt6j7NHNerDlY7rxjW2ErGYWZAqYkNJAIC2WfdzB3nsGcu9zivdMl7WBOFLYI
9iQBO2e4b4BVTupP8gRt2YJK8K6A9/Eu1EQYvA/WeHfCq0Z4LkKqz6JYm97IwGKG
6N4j07MQM80+JONSpPE3mf6dC4ErtRQth0ipR6/OHcvj3v6leHZpTpmZnTYFgID3
hxT24jJ78i2nJ1hCQaR9bURC9jwz6R5m0Q8B6xnj2of6MRMoll7XUfUe8Ln7WAAb
YfDPinN8/skBncM6LQjCXE+lhTZW+LtLXqLBQB7OIVWE6JSM7XeOk9f1lG7hpmAq
ZpKb+lm2uMLaM49XYvCyqUcpHp/MSU1giMDC8eel3Rzc6wpg3as6ECu0CoejePUb
HzG15hbKWqg4eLMs3WiYaGkF3+C6fjsg9Y/bAvKn2kQ=
`protect END_PROTECTED
