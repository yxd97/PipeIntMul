`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TS6NgeofjkejgcMUmG/yK0+gF+fZrHSWrvjW4oArpvjFOhiHhP9F7I6/JjkmG3zp
IcNY0ra3WZ0nwIxCPfmo6JBmRXom1n8t5yv7YbEDfUHAJRNWHOs2UKhwHiIk4B6e
NXJZUcc4xX8PZaRhZhTE1NEcsaajRHH0jlJmIkX4lL6sTPakUBaX9jaF5YUnhnRl
BNTBVKr3gw1oqAcaG0Bi5OsHeqMArsPFJBuejVIRy1p8h67PwxYUW4BWzSGu6HhI
H9FWS4d0rhjxv6u249JP/sqKiJHJI/UxnXNp3lVjj/Bgy0fZPQd9Z5sExPdlK4o/
iRF+89VUS2xMVyEuOPKfC+piGuzwk2Fzo4Op90NslRftkVS5Vw1+LW3281RdV8HW
yyP21yYxqt7yYMF06CK5YkJ4hjGtzb4W5lUIZcQGrm3GfdW63yjm37i0+Nd0aohG
supRTgyGwaiZe2sCxadqhd8TsAN5tlvd4s4jBtPxx2YIk7o0eDtnb1mAtfxvJK65
+OZwBzk5ryysRnRYnqIoZ7xIa80nTxFkh67YvE4t0kRtOO10J6QTzi1gBh4XcYV5
BQsQJ1bUoH6IEn0FBn2SVUfXx/DCUk+/dqbkH6jXfn3BetiYmHX6q96u7XJIDiJR
3/nPQPC7HmWgXcdsfln/Cw0h9c4RBrQW1t12LqxkZ8AA4rsVRprN38bwl5NIScwR
K1KnX9srF0aQ4cCYy/qCXoOaHasnobO2F1R/uons+fvP78mu+H1C+9PoA8FqFiHf
Q62Qbze0JqJG82rUwCSRjg==
`protect END_PROTECTED
