`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V7a1Z6/kxjbC46G1bWSnd1B75t5PjBqE3Q93uTW7L3gMji0xh8PNpnyhQe0vBc9A
m7r+noEekrfEitSoZt/LO1VCfbLQrkMsdsnZ5gxrv7M9GZmAZlA/q3EOfhjlBcb/
A4VfSyakF6EsdUZIYY38Rk0S8G2FLkup6IIYRJddLxKU1feUh0NwMxwK9maSk2tk
dTxZ5ck/qK6/ERFo3EioDRemgPOIgoCQNM97Wmkg1aYgZs2Ax8cWUynUo1ypQz+4
AQapQC5r142zkP8XQDyGwmwB31ZmTltOocaf+chf47g4Y/yPrz6gP5j34Hjt1K2h
87vAEs19NCJHtLz9nBjOKd94RpPB71sAU5Fao1FWSOGL5Xf4YL8/Po9pyq76Q9Uy
`protect END_PROTECTED
