`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjp2yun3G26k3dWmYZOozeaiDM8XxBVFepNx4oTLJFSuQaLefKwU5Jq8n+eT4dzD
sNVNXfQVVArqjvNq1DFJA/AI2g7Q/WZId2K/d00ZuH9n2lxPw/XMKQsVIZf4kU5U
FLmjFHBzVZ65IbWO4bwVo7L38YXZk5PoCwjjTyXWW7MzlER7Om7my5/eZnMye5A6
Uhp+G0JDpnd86rrcN83yqxkBdMRjbWFtgttFk0np+cUBxFPuaN1lZZtUWbytsLEN
fpuBCyTwaFfx5dRNUdqnJbvpqqKKwZfQhQ6BgMw80BY3iQjYfB0qPU0PoxCpRYic
wcUohPUPhxLvwnXlOcD1+MLQ75wPMQ4qqKmYPG8RLlMPzTDevTrJKfRbObIYrj5M
VmjdsLZfp05yRUYMdcSxoA==
`protect END_PROTECTED
