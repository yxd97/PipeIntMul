`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGfER/bu04SQNaRAvTrg3xvtpVXLTsI4OmjMmy9amYwRhGjOspxwWPWye9t0DRW+
skr/4pp6PbTgxqDU2ZbVYai6r1GSii7PNdibwU1UsuI1jOwMOp6E0KgeMXRcyi6a
Gd6oJ1hq+qikmeqFztDoP2FfYGObTA8EB3UW9UpRBA38NzbFxFvy2A0u0xfJiRvr
sVAZezMb3jfJHXeOx2JykA2Gr/XQ6BfYx0ZbtNP4Jo3/XsSDmw4dI5o5gCr1mAIq
p2vznoEiNjY6MUTfR1HafCvMBdP+YOpIh6iE/hsKoODSTE1MzKG9uvJyiW10sAQy
jfS4ja/852HGAplceQv8zTj8nxQoiQpG3+H0ThtaNY7U+CcECT1zQskHdiab6iOH
EnOHyr2KuUhqLkkG1hftqjrkFFRLSzOe+WP13y1j06NCktVsrUh9yhyJsuR8l0Rl
Wjxuj7C9he1Zj3ZlhSzaNvZ2ELT4TETfxDK9ntrTMoJyHse/p88lzRd/70Ir+K9m
Kn12FgQ7K2G+5eXrUjBpmjZFCDWDKSQCEdiZLba2xkyncllGC6ENzVURWvVP62re
H5pqQdOF7+TMw0mkCzsE9L9aMZuuYwduP3gpoy4Ext+ej4XetMyrrXn53u25xzs+
PLh5boh3I5GOCQ94tNQ44avKBszq5VVjf4Sz6L7g2YtGl/R/bIKh8qdx7FezzZFR
Rz7cTKXrlMw7hg0LelfikcFb1DywFqqBaNtctLK5ujGUVTSMvjjLvn6iDForiYAu
nmzxz0d/z8CjC8qNzbuTUGNge2jFelHeCeyrTcNH7Fc9E2bpid+U+Tu71AQVdiuL
MBIiG7xZsBuS5h5MLlj8j1vPELkWidhMP4Bm+O1fuBd269Hm6Tig5CjHx+0XTSnf
akbjxCBUnrwyjhRf/7NgbIJ963QmK1/Jw4Bo/STCIX16+IXzjPsxJziZzh+3oZq7
+dEUba6MZA3yq+JaTP72BQpERxBXQFmEILBykZO1aSasGTQFunUuh6nT5ZMiff9y
gK6dVaOwpDkYNvZrnuVkPmcGbm1XdZRvG51Cp5TGpV1KI0byqiccgIeVLQlWNM+X
FG8Us5O7BGiiimZDb2IRzohudAUagXVuDMeAJvUVbxic8g9nCDKNNYn6b/gZ8VVH
0gg9cKLWEUrI7669YOZs1ymIz2O3GzOl+Ym9/nlenAnwRUTfwbiu+V1TuGz3lsp4
yFFwkXnjg2hoZOq5VhfmH8tWab2sCjRSsChQmZ9VpgC5EfF5e8QmVhVr+J9iCcMl
9+vzG1DmTnGxyJeieFjDCD/tAuneZEzgDNbvBz28epKcZUduf48dmEZRUmOf4GMR
RAdoKOhGc38mtOudf4oExneKrqnnt3/fu5K6kAar13ElVeIUe5VyeHoKJK5QyWVd
k1sZ+q6PbdsDFdLwSPqaU+ePkAYmUZNZnP/b+uyTUWa68HXVrilNHUbvQbEMaFtv
ftqOTrVSGX1/H8AubtDCHVT1rEUGjlQOf8g7yUOl6tB/cAHErhCPaPchesxNRrlU
IzXg5TvoetTedsYpl6IGPFZPwACYHeSfvpzufI/TSwqBlGonxojLZUvdwT7NRnYx
ODitPlXIh5Yal/X3bStqZIvTcNhEkSXHoAKOw9h6DofcWt1kiv98n4E91D5+Hn1+
dIkebhhtC/TWwgxqGPdyKPVztGlUoTLwtqo165MddiXBYAHsU/+/oFut9TNwz+ve
m//vY3aJFDgTbIsKYbvr4y8zKn6OiWB4PtL8Sxy9jLCfKUQdkR0at8N1zF4k3ElB
7vFtOHcpKfXH7A4sDy3CvqTc8aIpK56nO/+LUXW27XV8nT8HvVberKf51fXKMF3j
I8LeReP30USmT4+WlWL7HUrLBuWgSqE5OwtUiPnprs4FrOFeO7/aauN9NczAAbHr
xXDHXMdRBa6BwdKQ5d8HC6CB1QDdIYWWlbevLignpsNmq9rvauw36thcYQMskdHP
eQOeS/Rb8B8F6f7vl1+GB9N8tLJniCiiWrGItbLP5UVtZQkoGUymJEZRH/eb8G6S
d1AropSsdF5lUViFrzbBGXbghBBL6itdQuDltBavIOgyEk+epG6DV8tOCK7AKNy8
qB3a05mr+8tb2cwzrFGl/zgV9Eg5pp3cRM6NBZ4b6+r5wVp/Z8boboqAsTX2yEyg
UEt17EE8rzwEgwYTGzlnAfV+fTOfioPctiD9+3h3tE5fkpVDESQhb0h7kB+3u/is
vV3jtBNl/1bH+djw35utnJzAp+yeB2dZ/wdyGGpkp54Q2Br/WJPG9VynHhsvlN71
JIuXT75qhJIH+rk78/Miy9whoMNTJ/nmFh9Z5q/b7AOau2nHqXDXr6sCQBh7C7SL
fw3YNpAzLlxat3N8SE3cxRNQOYt+hrp76nq8/BK0un7EgrRpCkCf7rXM0/3rgyel
uGnM9zCPIXbtIOMfVuLkT7Gc7C4V9rWGCKdiNOV6YyE4uJ+zjoYhFKgqzuMjnWyy
4mDgMJSETlDqp2ETjtV+GqwJo6t/+zW2zsE8v5jvLXyvGxZiQ1/rZazBjWsn+BXD
Khl4dx2hX+EnT6belX1F27sTfyuwhCbL1OYBzNpPx68/oB9d19RkrOUIAJ2RfW8+
MR3HhxwMcPnq3BgxaPpD3K5IaG92vgUNBc3Y7qafNfZBYMfe79xlZirYO2EQnwqd
4NQgrO5j+i46TgFKRUGzWedwOfKp50rr7htwCr/Ayfan8CnGimHWIuxtU8vaeAMv
sK7p1htAOSqFhR3FYaOk0V1a24SlllT0jl8GBsWvNyOg76pwRE/BgBynzwXHEZDT
NKaSvk/YXJA9fZIBZWdL6R0f8s8H93qa1QJGqsQfc8vcKhaI2ph+cKy3748D140t
uHz8/8Z7hRST+QsFnQFCybYJxm9RPtFNxiYSF7SymayDHSivu2hbI+CkNLT6PF9/
G9TVIKx8OqXDKOiiOkDkLegOujyPXUV5oXtPKi36im0fiYaEYC2flaPlGvzEFUm0
lpUiP4bxqXK5kSqn1f75ve5KlSo9VU19M+Y25NmLizPeAvvgmfhiXsFHHV4oSbV5
h7BuFXkH5FmZooRp8EXCTdPRRxAAgJnzDIwC+n9c7s6hOgOJGGYtaKIIsdgJj4Nx
pRgr9pVUOKJZa64MiEFvPIfO31J/eci84+if+3t3m5RYS0gPMoNIwzRuQlf0KwRB
ap8E35Ld+z3DJzF/Bn4BA6fmSQAkdk08g84l7nOD8Qw5wa+grm/72Ld69QlozQp5
m0AhJv+6xJAIJB8Frl6xx1g9bQvnnawC2YhNwhjIw57cdsqA6Xsydln0+ePLSpNt
4pAIV4KEtB4ANefF7dJPT7/GYRdEPGjnZeyJ1lEbs2gB2GOn4zQF09yKY8PVpjA8
1pMeK1X9saI1kRYE1MmNuYoQs4EeI2gtW5Zgs3clAESVhEtGr1VoBp8oUX6CkTKh
B0+bvuYbbTLcbZPHdknjccPtBSSjtc1I++ZcCW+QcVuwuzoo8qGjJwHSr+DTzu9o
FB4RFv4NFJ9sjXa+BGLqLZ/YSQmGjM+O2d9iuww6wzm82xL6CK5tLSAdbBtiiBo4
gZJLFxm9DhEGBXlKblLi5CqVxwheIhc4zdAt1L1VZ1FEVpxsevHR6zaUaV9EHbxp
/Ef9Ft76mMr5LnAv3ur6/c7l/PNSgGvGM16g2Xl2zr3HumUVqAi8g3oJJka7WjBv
63ToGVtyDbcVrYtZ8jrYNFS6rj1QeuB4UBwRYIKauDww+SVmADPPjfKvVsbwrd50
hhhoG+dApOCS6CtLpn16WvKkIwrtcsJxhkoiHPYOl8v9VWKAQUJres2sMzaIGT/W
/ol0C1Dxdy3Fsr/1qMArE1IO0dx+QtMk8R9H936KuUwR97fq1bwhTJbBsIjzvH4y
BsgilhTYQ4PO9r0NoY2M0P4zkb4oZp40CXDX15Ydmyl0i2pEf4D8BQd4Iis2zJNA
mMwcMOAWGZCnBT9jhuHSbzX8P+IQxe8bb9hlNQAWXeoEcInGoYpjs3wPxNYvjFhU
zncByrrmocikXhkihwcLN6wr5XjsAojkQxZE9dyNRlXAXQAK0y23lNvIgeWoNiSw
viUqoUOasDC7Y3VEFN2R2wCHCNqrt+t1UnlrB27vMSz5Gbp+Ku5nt6SiHRJL8hGJ
VCYP82qZED5leNWbkZoV2kgUDYS4A2+R1qnjXTDCWwSvcbOJHx9RrvKq5jva1vrS
jwoWylVAUx57bRNJbAfE/nz3k3hPWA2jTJpU+2giXJvugwSJQSIjDPsA2wUye/ma
ACo++Ax+UDvDccxerbx3T+nEjeQQRJCVq7jGw+HJ8v4IRKZVUpUZbHesijRkxLQU
BJG8wirpfoiO7Viai2o/PaZ8ZPOUpr0Lzdw7KfDfNihZKttUkQwqLfYhfdKwH01o
ecvfWhg5mio0nH/V7pnksNkH75H7ck1F3FvXGpwS42GOFitJ6K4VPN1faLxdmEJ3
XnQmguqxC5o1FxalQ11YghvfiK88vPuSZ6YRQPEcJPeiDcIVEBUVH1xNBQLjlSOK
jZQuaqaXCIaQEm5edmsujIAz2elzAGHUUWpKVey03uNSBWvyTkUm6z1C5bTU1mbG
wtQULAfAe/JgOMe9PgMKnBk7ai+nydB4v/9jWkEIxOE1yxUgfnltVWWdak/Rsvxi
PpCmm/JPP18fqeCxBI6TAaMP0VvC9HSaJllzyD6bhy9ma6M/wBtdhpTQGlij5Ud4
Lhpi1bGMQ97RBmle7hgBGO9oAkVWAP2M2OTBcOtV9XGFET9w6ILoEK4y5/1gRMV9
asRL+KIdwiq3ZM48UViQsDUiSgFljAqIzAO7dZV1km0Iv1jJTgwOSs1YhzpGwNrn
emWTqhyQqDJ3pqn6wXSlRYCYg9ymq6JrQv2LuG7EK00wAqp5R26evKugWHJTPJgG
MJiURDvoFol25kRWp28Lv/YdDRV8p+xgkgrYKzOkmtVfPS5gfbTubvODHg6zowXw
DydjwMzOOO82fyfCgH4+SNNxCQAtP6YHelG/yVOJDpLnuhGUjisVlZIETbUD2IrN
eiymg8h6FmZY4+DjcWIi/9apPV604nHoICTrUQSAU6HOKtSBCalD4w7Sc96OWtJT
0nI3BrjNd1b21j9mEia/L8872hsxB62/6RAyYwCk08c2s1yGSMa1dHKWFqjZ42qu
QuciRYDZBwbYONvfeGk5lrmAH5a3g74McwS9eYyLcXncJQXMzX9Vu3vEAvLU/q/w
oapa8LEMf5SvVJMk3D0rzCI10dMybGMP01l3T+79RbghWHfA+PBD1xM63ojPB4jU
NQfCjpTfFJgm1Kk+LQLLTzZFnt79FwZSXxhb61tFBVHhH2x8AFKIOUQwfMP4waDM
gHU4/ZONIVn8+UfGPW4ceAd4MTVAKbBJ5bmydwIGuieWhfWtUGXgCCqEKa9D/JfR
4x62rZlk4UbkcwBIu8eXqNv4zyw1Dqit85C4PTHcnlHQe+UeED4vzFe56DicbU7Y
0sTET0Dn9w512KJJzSnvqpKmGH9Iwy9rPf2fyaOUTnD7Gv2g0muhpekwDMjhwmPL
7scWwJy/9B+QLfXoNCxfdUAAa+Da5smBqmEW4p0aSs4/YZrJebQDiLZs8jQeoQwD
DnXK5xJmRILj1FpbwRPnPw5LltmrVYtTH0MGFX6WBH9Cj0YPqU9rOMc8YQyaLc9D
LbKBE1Iex7DKib1XNnAL2BgyNGalJvVB0XcNlR4h91m5yb6f+Sd62Svq/1VX8YSV
eDakgILyQ4LGpNBnKIV6xykoWEz4Aj1mnXNhSRsUyI5I7O7PL0Vi9vLWu+hBoyoZ
pB+IVSl0l0BOS5zUH35DVg==
`protect END_PROTECTED
