`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4gNpV4+lWO/+DkNYPeXo1nMxqNrRp83qZrDsQDkLMWdLVcefV883YGq1kLN7p0C
AnDeksJWDnQtqKrb8JVMFn6xZ03FM8jDSVJ1XAjvpYXrjYr/OvFYQBOQwlAeouJ+
/YJ+9DfGZMeM0RFfOiZEuz/4dp7ekzgRw02442LSfVzNG423/SOGGC+LQTQxuBTO
+oB5fINhqw9jyXmpUppz7PlT93JYfRem8jGMG4U3mR0HAtozAQxhO3voEAfse980
gna2T9gCSTK5wTsD2T4OYTIV91FWxnlYuYdV2smNp7nm6Zzil8I0Fg2oNYpPDqRd
kaH3t6bO1Njv5T91kXg03yOS3oZQU1zbwBTtqKW6lvk=
`protect END_PROTECTED
