`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bD5bm30bgDqDI2UsGK73R8kjnwIR67cdFq+YtfbVOJ+9hKJdygkh6Fh8S4Lvzg3a
7qUj+uSPHZMVpL2JCd2J51Xc+PuwJPX1BaUWo6IjpbrdW8oBF2ABQ0jRTY3vv++O
nolwuI9lIEOvEOxfZgL10PNCXK6PIpu8aUKPsfv5WBmcfT1PSEkvxvCIkvBwZ8W/
J4291C/8FtrEhrBS7GotjesLLZYWIRGxgm70QAo4D5h7lB0zCtuVz8URr+Aghpak
Dwy1y4gsbY+u9++0VrUInp+ZQ6Q4UKXuCovUtN+TQi+XOYx0lC7UZzx63PqUoceF
jzjfjn1ZmsEAISamUVDiUgjmprg8sJSlFJW6Cx7fPNRimW8hxhFgzyxHI2Ziad7R
QsI/71guUMVhHbIMYN4aG9pST8y0hM0/SMmll2/YenHsz5wQklCupIUK+CaIO9hO
15JMndnadjWY84OdtcHWdqxopb5AFJgp7O4C4Ktp2nDQj5vBLwHVTazk/h/k+RI2
`protect END_PROTECTED
