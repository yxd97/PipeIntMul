`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rxbR89oIMibFOMTXpOMwxzxIcJxdguzo3Q5wWq/3nhczYoIVcdpyEcnd7TgylD2
SMMKD3aG+RLKAm8lKLCM0FCDtB8FiYSrJOs1TJr1aP99xRQzOQanP2/U9NNsd3Ds
3KbzOLgmmvBhSdZONXxmQ7kFxwSZ7LhGkElTzql6H8Y9kaWWaIZIKPYRLlejocCK
zrr7ADkuqMdlPapM/Vza7l80/qR5NcrPYKhmC4iPC2JRn++lc0tdTB83fWm26C8+
5i4sL8yFGqXwd49Z8SegLhWKEumYjh/8pxCxnJTn101ZPk87WAmGRygPZXNZlOg7
OSGheeIcY7VCYJR0hBVH4LLrqe+znr+ccOJWdlVRHwAmw8asjziM7keLeu8h9AI3
f9bTyvDOkNf1WICKHlFTQC7HKaVnxddFChyOst3uYsQvWoVwAcs1iaMoBS2LRY2K
decVmwmqfKqVpykULfbE6w==
`protect END_PROTECTED
