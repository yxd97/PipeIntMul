`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
07eWwp3nBLPh0dz/2qDJeMa1UU08/5Amk24E5eof0Afu+/1Yhi7Hw51ro2cTG+wc
KxP9p1XUTxr4TFZC3KEklGIBrbTrbkEm9k0zlJ1r4OsjliT6i/mBehZwwg7u8lbz
mBggUy4r6gC8zt8pG7EHJJk4pxBfZtelLRORyX0M3gv0dpidWBrFwIrU7YyFZQGc
XtMxBdxHTrRL5p+EzpzMfxAimk5WBTWlPppyuv8dJzAZXCnh0097Co+zoZ0Sudpa
yltZOXgikPTYJN35G/rJR9wJk3yNGs0tsw7JVck0Ju1K+DkU5V6KpSwYRfiksn+f
r6G+KxZZswIQ17IEBlhuOI5o0sqvR3nhmRb9FLmOzSIbpDlxjL+275/zdlaDkJDw
bKhdeJV+DBzrT5DvmQZFgAl6+JaFFPUAVeu0fomXlAK0SBzn40rHWoQKsPL6T3An
`protect END_PROTECTED
