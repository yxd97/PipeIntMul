`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7v26PremZacxU02oJIYGpiCe9RwU/waiEoaqkTpFjs87hiwaUz3PzmV39NqIsEkJ
+RD4P+7Kc6bQZRanMG7F7lCRl0e+t0pRyoKzGaGxCYVq1sxiWGOERk3ViHLLyHql
OHL2FTTtNgg53db2uHSu7ieS3ROsWq3xJKJpkuWj47nb0TDAUcyLJ5UGdkP8eHHX
Ngl1mjNH3Lo8vKJfOO8CDtGC0LSjkrZrdZTCC8sWrdmDy/krC68bJ1b4c8hlIX2k
LyfJ5RjMlIFLC7HdUzAtUKfJOMOZCpqrK/YKuY+9r3jOz400T8R4j65HY1rnWuGj
9w2l5tdo8kkqwb9qzNPVTUVNp8oqPBgnaM99ukkFdReI167RYvHRzUgtiDMEO0k9
dsBcB75OmPHTn5NjMtHcrIPb//ooxihiJY4s3x4kB7BEyoEM9aMDhmRcsXYF1/37
JpDkrYxH9dzl8ymKGFGR/z8Wb8WYzfKgyLe/agqM3Sb5aKXwNko28InbS/OSV+HF
z8tp64y5uc0Uwc9dwe6RLRUfrQ6//8lIWvefELfmKpcA07r8SsxhbMY8AcHkyF2E
qP0t/Dh1C33AK7bL1JSTHjIcV3g9UUPUV3YG+xyRaUphoTHaTWTly8+YqAtyzmHW
IqFDAMCGPJrpWXKdBcmOz/rEq2Lx2ustZ5iLuN3m+gD44wbNob/UCskEH76jGMuE
IOvjBKbCgYDzt4zWEh8lTDefjQ8uTnBoT4bWvRyJRsb1w2qOyLoTLdbfsrz+iDhi
hsbg3w/5XUSgQBURLFCEFuX9etM6tJbeDQAcqKI6gtYOzT0KvCKDhWnREKWgBwc3
zgw9YLLdFJXhzSuA9L4OVExGm+lk/hfzDlwHdkPvZAz9lWHtu2/YzoaRjMud3sl3
ztf+t75kTxhyLss3fVpzMj4v8UBoOiFL2jZNAcxGDQqnG8CGEriKuoVBFCJLjx/N
U6UDIT9+nphI/G4p/zq11HDRmC3ocsx8UddONnKlesHqCNh1ip84tyIuGHomoDa6
80romTcWNpU7E4OEnmNBAZLVNMMFtsSfGcaDd3DuegzZbx/OsbVkQ4ki7nnOCl8O
O815v1NsXSZgVnlIpar7O8crRuNCFnabSWptr+1OwUKes09PAuUo7iIZ29qCkEhe
KjO4gCGCbw1aAWNEVqu3ZmiHv7JrXqT7P/6bQhgjtx+FggRNhmgqhIyKfX6dkf5i
SMZLHTziIr6H359kjSvXhg==
`protect END_PROTECTED
