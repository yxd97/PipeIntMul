`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zIqezYPHnDmqsge6dM8m1CpIDm2MlwrB2CXwGzS/88sn4sEcTiN+ZysvQYB9s8v
nRRnqfXxYnjAXQnSE62tiu/opKeykKQykZIK0iU0B8ksaomZwIWIJVUul91w1yQX
/KSWg9HyZ9yYEUdsom76ZYfi0UqJ0G87EBWHQX1dg5TZBHXoFWw1/BW5rt8Nequv
Dopt+Iz3hCfL1RIWTAjOQra9jY6Spyx2Oj+i/7X23R7giAwdwSSb4DqfjqaKUOgP
NwoNa18Aiu7QROOmqAYFQyvMAkIJ90n7orPQIpn5ocvRgoxe/SMRPgCfhzC4yliB
TtevGwFql/iMSxVEUwAdCPdm577Ko79eYlMZN0wlNR1yjfSkptgaoJGhZAsgi8lq
5AdPbjNJ6DC7DOidjqBFZ0uXwfN9xldhraSKmStuvV+STSAnR5xhmYSfFUgo2U9Y
Ab8Nzq2y+noaEzNnJwGjkX/EN6g+pGoOSLr1KZk3rXaJNgyl9SK1emwWrrZ5tK6g
kTzeieTDjNugE6PrxK9A9CjfmyGDFLg5iyPXXWP0rtFpETRcPAkVDHmgVk2ewuf6
nqJYXKnBpnho6RadnxlSU6E9ayyM0Efsz2jqEU+tWFqU9SH0NRl4PTBOMAeMutPA
DvMY+TspLkmTPG6LYLB5OQ==
`protect END_PROTECTED
