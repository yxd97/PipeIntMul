`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+p83jKx+6fP2yshI3g8/1m95eBcIvpFuGBkPEdqk8AyUNnHpBjkZYExMEKAexsH
KRnMP7yBatJa/PydiNGUKB5cDllwjNEuT+uGuemoOtZg7jP1xWF4kWNdECAVXRYI
iv3dPjxg8FhlQRBI4n9BKgZQjxrg7CvZv1bGDs7oSQGtsQlssOS2dQPKNm5l9l9G
Ks2AN/EK/YU0Bvze1Ro6wPMN/FT3WbNvlcooof2gG73L9frXcc4m5Kzvo2u87kKP
`protect END_PROTECTED
