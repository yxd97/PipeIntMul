`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TbvLAp6sleIOYkhnh8r70cEx2z93IOfWv8sp0spMSiugvCwuAEEhOGpIRtF5/3DH
Xg1loONEEiZ3jYAkb65sBGtICFrg4V4dFfeq3TR7afLMjrO1+iU6Jhbfb60ma84i
aM2LS8JerTvMA+mFYnaoPdFnO5zvfTjiWGsrSQopQoSD8so4sVcr4BF5JCrEs6tH
m2k9tsNr1GOi2PfL0Eosi6XyNoSpClC0EMmUfZhJDw4GA6SN6cdQPHPLQ+qTnuz4
C3YzRVEgv/HmzcQZWLouDA==
`protect END_PROTECTED
