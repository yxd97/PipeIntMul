`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z539xTzCMAee0nm6xL8PBakM4qku630feCUcxgpODAy1E9y6BH2fWEcA6Q4wcm9w
XU1jC9fgTfClsu9fQ57K8q/OGdyFj1POM6g64+FzlQ+9HbOy5Qsv/Dgp02sBWBhF
aKOpPXpW033lIIXgUGAk5Den4rK9HN6idgm+6bJ0ZqAFEVx66LH5uTJ9NwFZSy+o
s8HuE464S42Q89CGCC7P9IQJJGh2/Yy7xuoG5r+aLRFjy3Ya9MFap8LoscQJ5uKl
GFAl8qTIPGsKL9bbLyRdMKSbOkP9gzwGsKSQdnnDZP6JqSTWCoP2UtajkfUfKZ7Q
K2MmJonjF587QRPvLhm23pdBMlRGzceosvQp+MoxfGAbh1cRD7Zq1+8WUa/8z4uT
7ZIF1rL3pMuXeVV6pZA7Lu2XvS41NM8byM44G7nUnLv586a82Vc8LyEF+gSeb8sA
K3ybAszlVwMnVCbbVhMjHCPKg8AXyAvVGxtjaPppGduC5azu5I0QYc/HeObnRbUc
ZsPd2qi15g362THpRuL+S7fTnUqXfwNwofX25cmWILuwIVV9cAFwYoyLmGp71Xfc
piA8zWU9Uc6EdsY7Lf00+JP4BRcQEW4xmIK9huZPdAEI6XD+77U916dtxcyINB3M
ZZ6Q4CzyqcMOttIoVB8kIA==
`protect END_PROTECTED
