`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0i7IyB1MlILRs2LL3j3TI8xlqCWqTQsOJ4TsW1crm2u5pYJ/+WogwonHlUehT8NC
p6N8fL07nBthy9m3mfRi9Kehq0abXiqrmbhtbQ2qNEdInZY6FjY50gkvnF6ZLewt
5nC89ZIZoEu339VkjND8c320E7KenXyXYGhgwYzmH9LVu8zhpFu9T5OTeFDXWdNe
ByZOf03WRAUM/PBRDH3u0l0R44QqN2rTAQ80ycQkW+6frQZeouVuPlcr1Kjh9b/w
2HeKydTs1+2ji5ZuRs44kvfmtCNbMJ7najlv0Ofcj9U=
`protect END_PROTECTED
