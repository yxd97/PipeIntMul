`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBYxIGc62uGRQ5/vHpVSOMVrk7oV0V7r49Tva6Fw11VvXJqmzk9gmh2kCnjbWYkG
n1aHOPT1WT7zeGcDVUDbFlSDMyDFDG5Wdgy+Lh0BaK+5HWJbXQniM3KVpQn8GLtd
xkEKdzkUw/GDsKjX8dGjXAfyObYz0GBC2DOvqWQxSnNdgepmfcPxPQM5oqfm8hsl
MpYb3M9aEb3nXDIhkpZFVoK9bAPz9ZwiXEBnmivDsj+NEWYH/wYTKeNwhaU1ZUhN
aUFhoPlw0NKXLCy+QIyk6aehNTpTuRQwyTJUjZOSB98fjtdhf5C0rr6wvtfPO/PX
030etA6iJdJMSBC6pAtPvYoLkvBeiYqMPdgsdzraFCzXAEcV8Uhom1XWkdKxJROV
gTUdL2z3gu2VnoIEnsnNIvFEedsPyr7dfL66HvvQtgC+KyuS1RZRXWvI7eJtxjsH
`protect END_PROTECTED
