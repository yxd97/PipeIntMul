`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xhnUaQH/9em+18xRkSNaBQ6sgSTU2FwS21acFGlc/Kc79jCLRzd5JCQl3gHp32Nf
9HQgo+Ht4zQDb0HGYwUVAx/YiuvvcEdnjT53umeha2H8j6+my1Al+yE56VoN4haj
mP0zeqhImcZoEpZSgERU3V3T+L1LxnZjkKFEprWYCF5S12D4uniwdKL9P0+XBLGG
E6Pjpq3hF0S3uQR9bmAugosz+2aQoVFNtRJGV1eax2AGgrO4OKKdtEbUvH5Jm1Yh
8AzCaCxnT0a8MxZgMZR6tGvpnAdI07RP3y6PYtgMhnbTNwh8TvwNSto9hJOQAhuG
DKckI098WytpFFAfA15uM8x84o7UU2uRDmK2ThCyjx2deV6/WJo1XwYriorEsAur
LEw55vSO3gH4Xwo2A1l3vxdNXjIu21CrWkjvFTmvb3dmb3ionlAX4GOS/Cpmocnl
ByNLHL62wLdp2fJT3And881rG3DSA339WsshpCXjiRhEQkLVP7uPS9egayn1gggo
`protect END_PROTECTED
