`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mo2tV5B45VUFHgGYsSYGErkFDJdS2J87noniZiLnJK1ULc+9U2YaHkAh/BiHFlMK
pbMFzdjSodgwcVoCEsZQXCBPqdRimLvoQBKc0juF1nGsS6f/tOl2tSAXyBoTyp8M
8Ddpygoyl2mBN1w7Ou3M4Ki8xsMkNkj6fhsEo67DN1II/0LbmjiIUykUcmAzyoiT
2Ackwrs9T68qfpxAxJ8syMFqZvvQe1HO7qj42Ty2+NmYLlh4BunEZ0OV0iOSqLpU
MJSydHhTanrIOQAjuYBFMWgoKfmVDCnUm0iB7JeZTGj2EjQsqXBBTrqxrUTXhCTj
lYkDNbA/oTnGaGxFeO1gx4vVgZ6dcjzh5WTE2YMggp9Ba+EKIMyw/B+Dh28YzFCL
dm3T+KhCsyBlK4EzAT2E0aQRkMgtjKRe4CTD2OU/LDqguv2LN/jVQmIoc7yB3O91
/b0zmxUha4YSBpFoqR2WjUmd/eEd1BVS7oVQ7S/8HKUGa9RxFepjugpwCEsRXaYN
Ds1lPq0eFMCC+Z93CT1Xr6kqjU0b31gxafVL5qugHKd7qKGJWecQTU033RKbKTPZ
+pv+zNtMKe685L/NG7Lz7zJXSYnUk3fxXjYiI13hYAMhj163qRmAodkVrOsu1cDY
r/MlpHLpxNwrz9EmVlF1KgsX0teUJ2KWRWwX147AG23mNQvxyJt05eTmA26MFysC
uGUOuzLuN5uQ/NNbJQwREHWzAz/LrPjUtsQsSvNsuELsJI4VwO4jjUC0XPGYUp3a
WpaGh5ocVTvZsBsTl+2cfgHkrznqXVXq3dPbVwikm79rGpgVou0zjQRZ5tQdsOMl
EjkYY1k5DPQNt0FdOkkp7ljYncPyYH/46d0Rb6vIJZTracRnwI5qiuF1WsVTFB2R
LNZgCFGsyQ49ZEMt3mNJvA==
`protect END_PROTECTED
