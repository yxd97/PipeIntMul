`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGT8zFzAeKPsIZmFQWAd4QTOT76WKLuVO1Z5ZPnQSvE5zcCtPv58lTQetpG9aFff
+AkV5OdhxeNmfza7l39setwTh83PUm7p57MfXzfAAjBuOFjDLlwFWRGFcEsPTMR6
zBGr1wb3xa0bkjH5M7n9iLzDLoy6G4Ht8K7BWv1yJGCwfrOh9npnNml9s/s7hmxD
KEmK83XoNcy3zH7MFrWjhBTDe/OKCW4tWQdfC/p7x1glGdhuI1l64ul7lnXmUCp3
GSPZ5f0ffoo/MRmvYrBdj1r5GHByuyUVcm2g7jy2tDO6j4PJPrl0llS3KzsQIQxw
1hFCgcIQQ9011hJ6vV8KFA==
`protect END_PROTECTED
