`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YgeExN6Z0eyiRD4RFB65bJaQcXQT5i2PKt4TsLSvIcJo/ZZQOlwB6whEuLyhS7mo
CoF6DkS7f7a+yQMTrm+NE1KJuAJnzdtYC/Mbbnl9F4CrrP3RNuHm0rXU+TOBOjjD
tl3VfssMyIDPEadE8PHY9wHm4CC/p2253TS0rFJp3pMFO3ayNNnM4btAko7nlm1Z
A6HB8v5YBK1WVXt2aPfQ2U2E74J1g8Jm0a/IojiKfeCHJ2uCm061vmcQzc2cLfI7
roPsO5sASr6Ke0rfwqgvVWv3EMDLRRZzyg3z4Y8R54IplEmMpblDxbHGVwvgJXSj
iEgFpN/7gxBb7EPGaO4ktkwj5NwRwpVjO9XMF/8AATM3ucvUyPc22Tp3LLvnMEbR
+Pgi/WJYra2UmS+0FN5sPUYMrYmnQi3CzNA0vffevqvQD1AGDvlz7eakDYb0qTmW
x8WkjNz7gLt8UWGLnPF8nPEnfIN8wi4xQiaTakJkJ9RFf2UhnrEnSwz3fbs1qHGt
DaaR+G12SSY7dZDsook5Ss/RqKUhPGUmfjbG3rdqmta4ubASDd1/HojemZBdbMJG
AOOlkSE90S/IAZ44lwAJdg==
`protect END_PROTECTED
