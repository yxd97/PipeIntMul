`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRB4Vw3Wdsu9BOIPj75g0bADwxegbWN3ayq/f8O4yaiZljlNLtVH3V7W/vWh753b
FUiVKhP11CXupMa9cCe8nB7IGBngBIhbElLZ9UPvhezpj9K/AbIeXCsCc/vT8j7x
gVriiTtUIlbr2q4VnM5uiCbTowKFNAL/9zmrwwOkb6dAJUS1OQTzJ7D1qTyQcwMF
rH5K4MqztngI17CBXf5uitveLERjlWPxxBG+eURotwrotGjrTz2wIqL3996KgzBw
jQX/Of5LqOIAJx+6KPxKIBZQKpqlA81wJzEJArVSKCw1hxfLd2VoNWgkU0TdGqVh
BycjyIQzhQB019AGGcsnDuGzdGbul1dt/Z3dMu06/ObeHV7xqiU2DoT7fo3AQ+U8
Af/6MI9R168kixFq5p4Q25VyBjAe7jgZ8UkenSb26X6rmrr8ovQS++F1PqPHknG6
yKIn+F+Bg+5AU4YuwTySz8AdYwyEox1UmL3CX+EUE+Za7StA6O/heorm7eUIWuto
Mx/pHbOfIxquKUfRijsj/xr7pSSIrkt32Xf9cIzUI7ozDBucp8W+mjzYb/o5JIi4
C8gYwIvIRtbUgY3078jXDalPSqhbMNBhu4uz+863jvnR++jWtyRVZDyk4emKmc87
o4H6IJu+drGDQdQQbRQ7nhwSO8FhoEn7hjM5VoRcOI+Dwpi8100HN0g6iqk2736Y
uitNYxWRHnUUJE++33J3bAAHjGHs/8gkJIxTwDt+P4A2W9L2+lf/FWnDO6ih5AX6
5j4vGnPYCFRQ+eyhK0hr1kD21TDogtzxWZ+5H7d3gFC8f/QMq0cMGyU3SOoMWCCS
f9tn/SrGAKPyphyWarImFz4cx1YnCbw+j1rsprNg4y9exCcTx1rCXNRO4BKroz1F
yJMyb/5SLcXvnI/v71pKTnIk+eDTCxIaK/uW0acdt4Jgyp8RCCO+9t1kQDwhtM4A
9WnvqhyXeCDK5aMGAxjdcOFJvSZKYr6xuhvJMk2qUK9GqHGx+XtlcnryZ7lukrCX
j4wc/SkoReUtJy5c3xV8GwfkzKK7jU090w8t34GAO0K3CTM1dIgvYeuC2HQ7J0gC
UD4gt6W7XVt5pht3O8BlFGo5KgYwZN3vrClbsP9xE0h7iYotoaD60UK8u0RjT9gB
4iKMKhecDsPdFgXOaZ+dhkR2fXaHwRibRiGGddm6vg035X2ga7flQrszWEjLDvp1
SLlT4LHtebhCXza7cGS4XSvfW0xNZyTLoX2r/gLtkfP2wGTiC9l0kPXU1CERCBPj
ZBmu6kv9EhykJT6lEGJoeYJ6uMbwKpox59ON/k/w+A5eeATFqNc39kNMOdSZi9EE
Msyz1Uk89Crj0e2ViEONLK8VfA2xqKoPpXASk/rMEf7cMZ3tuj+HMInMH5sCJzgd
9NuV57osoW4p+nJv6LFslZUzvwI3w/ELoV4CyzvKIzAAvIaCmarozwR4MBHThI8T
QaZ1DJpvj6XzFWQl2epNZV52Qd7Q9q7aHxlaR2kXc1jpy9rwOpmDReo5cRis2cLt
MF4U+zDGw8YMDcY+J1GIzdcspzCIA9wJGeAfBs55DYrD8niI/XPkrCHi/r5p81BW
WLpxKnrLLjjh1YfbivnxBtOtE0I8q8uK09h7xowwiTQF0IZVGCU2nXszXUcWGAEz
zGJr8DnRFYvzk4NFcBK66enyLZXz6D6zU+kJ87al/Wyz3jAggTXtEk8On9k9Abwh
yUpiaQacEAFrXuPF/pag7c3LM4n3nrQBzzjXdhcp30OugteA05A/blwetbnSjHk8
2hW/A6m+1QPa7OZ+agCEYnOdBE8uZmY8/Xx+ACSC+H+LXjRaOv9LcIwirgJxGcM4
ZzMUhOR9rUJPfX9n1Cz3vnIreupyIdW223V6LAwxvlmxiStyDz42QPNaMqVDjaLI
TIn/jebiYQvglFIodwtURxdFXz1so2yH/MPpqLfWwE4Xqo1sPMJOOiQUY5o51yGl
6b81rZVk7JBp7VsAObvt/rA+h6QF2Jw/yxnotDMjSRCOv90C8yNOo4+sznXY6isx
aYKjqn8yrPtj9QboSQ+bfPrzK9vAFAxF17F12kFaJMr8j6qYOLwVo1xwR0BeJv7M
R+SIjxMXG2QGp7BPB+pnVMqCPd9yJq+6PdMEa2//IAVAzjxxqeAaRp+LvYv7wqCH
Gr1J4L1jDIojRa90soIJcGyTTJcAiDHiCIhBXLBEdfB2exH0+WPeZgzNBRXhmoDV
vJw0fZ8CiTdhS5ncdWxfQCy5cDoMd3Oo0OkuXEW9XSUh8HzG91HaQnzsUsLnw/NZ
2zXkK0quWpGYZgA9j3keohfxxmD1qlJKpt7QZUUfB4kFglEpZRmp0XYGy0XGjFxK
bAF+CO/FUaDexCTldGeB9e/FGuHLfqJupTykuj+ze0pM+hhZ1kxEMix/4wHiAAkF
sS4RgsnH0KJhRG3kU2RkvQ==
`protect END_PROTECTED
