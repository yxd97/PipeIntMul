`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X4uGWcZgXrCBOVKgTXMi4hrEuxcEW6Y7Ho4gk1Xq6TkA9sQZY4gbXb8cKhwcqoCa
tbMrvAjPjnLSco1Zu5Q289nHq0/wicmUiAMTx82KVeZTjFWvq3+hod+hyXcM9/Mu
o+xxUIn5kHVeShFK1a9v/RqD7R/xwUjuUtOVwiAhV6wq/M5eF40PjS5/XJzBo4y5
T6wISkj10dWiJy/gaea6UDXZiikHFc9NTMcC5LqasbkWxjDV5ntCgLX/dZdSzJtP
0Pa0lZ2MMjWdwhkIlaY/Hcg5phWvDJ62213mT8M/JEo2OwHr6C+KMDHRQLg0ZUS7
`protect END_PROTECTED
