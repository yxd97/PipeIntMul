`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bqv/KAgTuoLIjGEYQ4TJlChmRBrNS5nsN5CcZ8ozy228TE57kMgTynfYkwPz+NEG
R3yxFtIjilyC59sfYvTIgP9j3lrCDM6fvc2x/EpyyPgVXmkfkrSAec6XHUd5UPqG
eGDd+ei3uD2+iGa+ZbLVG2qMhcO/+EKgbJgzajRagDA76T7Vt5H0/Xs4tUaaHIn8
w4uoWKRZ/vmokmeZiFNsykjDnQ6FMuqw9vBLmVO5b7kpXXmGFXwDgbwfnwO5qh7r
jMqc5F5CVe6SLd0dUK2Z6Pz6/OJkPlSpCcZggSI6YwiVMY/PfQ4O49N94WWZwkc9
huN0LHk9YykZ9MWkDERWWxWApvYk6Pg3KtPZRlMRUMa5ssDNHUjC8C40TTvcUj7g
oTyg+h7aaLDNnQo0yhfIpx8Sdrh0kh4cpiL7F4IcvapcyxuWS+KowITL/KiPaPrt
dBQyKw6LUy+vPJVcN/oRzNoRaZcBkSRlBANugU4gRrkNXn/O5OXV0jzAvuEJoHvm
`protect END_PROTECTED
