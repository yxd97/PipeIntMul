`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ma+Ql6tzROGEWN8AqG01Wq+lCgPHXbot644EG2gwWJZr6fDTzOBPNHwKli/9br8J
6j9wxN1Ji2WMEcjj9GR2pbrm1wwkTKvrIKJ/L9e7ct/pQcvheliBGTVjb4yfw3SD
Sn/4b/nOsDy81JXicFnP5yjeeQCIhTpGrVq/xik5qwaQaGlzhodTxz+THoAOK4zV
mTDuE5/qvwEgAl5E4ZfI3rDtrO1AFaDTtzDg/oZgB8n4p+RwDzmZ5DOIVdGBGJga
RjmFmUgrOogX7BvQqVklbsFPOq9Mx6MpmHcoM5sCfu/Gwp1fzfHMCEXc8Jh9ocup
g787g5oewyp0P5EbRhy2Fz8rD5fX59GF9i1Jdls36IF2K+QbBpPYFKTTkIKcHTG2
saAqKTiUkb4R6NIe4pUjhv0M7010mvOGR4lFsc4j1mdmDE9eEQkdjtsvXg+h6pX9
C23C/e2YshiML4zxq6F1WExlnZUmZZHiWnAgAZD2EPafrozKfKWe54EvSM8RXeMA
AJ4CkZe0sBMRqbg3mfxbB9COFnJrUSllCeyWRSaFgpvyT527Wm6V3/4LPvc+O1xm
nSHZxXxbSiaaYBIOP7K7YmWO+Xs3+zxlf+Dhf7uQCr5+uX0D9fS5DVR0kL4IV4p6
fd4Qz+0ehcvk2pN6R/jHESQHNjcUooMQx7GPTepGVzpN5F/hKYCmRASvEbrMy9rZ
32BB5pOx3bVyuEQWzlSW+g==
`protect END_PROTECTED
