`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kLjxKm5PWmw/FtFgW/TJ1dyYw/zfeuKTkasb5nFDGnGYlJd0xnzlZgMHq4UcqRV6
tOrf2wUP17I8Un45paw1edj66L62Bqbr7c8vnp9ivrjblc/rbQWGAQyiUEnKcSbQ
cw6HL+duicAHma9gTEgIxw47BNFsULDeIzYh6tX47DUaxvlTDwDQ172YwLLXG3rW
NRJtDX/BeYl62/F34C1kTBPR7wBo1kKN93C4t95xDkDvoPqufm0o9gd3j+wSwepV
bgG+BIZS6fDZ2eof1MGzSGfyxI9XyQgh7lCyovGGbE3XX//OeiMw6jidnA8DtkTo
zsDvGRowo2Jb7oWr/7MKsla+1T4gJwbRzc+ahhV+3r/uqflT5qg4xQ7VAI/vrAE3
uIHpqPtSeHDm7KTsT9mOaqJUzYePtLY3Bpx3OFxkp3UQ9fRNLkm55illgoHNGLHx
HIV3E076t8dsDgwBuTt0s/5wXlCb6eRD46zgLdC/ttEK5gQnJcgcdoa2U6+OjVuF
`protect END_PROTECTED
