`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85HKUy/UJgX6VlsuJ2HKr84fbp2Sw0zEq51hEpaztvh2mR3X4OtyKfux5g4CH9ER
3Ue9pz3OvdCmxLg17AJMhmY1lE2y2tTi7Vy3tnXA5aJQMKIXa2bd+/B7BqBJG4/Z
NQF8epPyClIZeq0gdg5lK+/tdMr3gcy8ma1tyPatexA6scjqhay+voapJaBOMWOL
oQn5/c5VCevOuw7Om/siCRaQBA9tQimqcfrrQBGbWSVQWd9ngLyLsFtkJuxjMYtU
fFPoCJmRp+qpo4Fw1UYaLk7JFuN/dXDeYGc9Q1AFQodoWxBt4T+kie7o3BrbBJd5
LRIIp1BjY2FRzXFe/P7cSNnGctd2+xxVpJbWTUChjsWNbMpOog2qZnfFh1aSND0u
`protect END_PROTECTED
