`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBhth88oZLoZXKe30iB5+Kt2NH2O8n+z4AFVydJoPxyEa1+vO8siVdQMobQsq7vg
PiG/DWlSzYFQdQ5ctQc0BSX67DGBmjxW67FqhKTc0xrYqSMYr1ZyDtU1VASdbGss
S9/lw4nyhV2cCLm0X/kqcp0XLplYSdyg8C+e7ZTyHU1DSidMXL8+mkZWtzDPo2xJ
XKh4+AMcKlHZiLUSoraDNUUXd+MaVtKpARKIxbM70R5dZC8s0zc2v1d1IgURL3uY
i2s4vpaR/W6rL0zOBaRDfsROyh3ZMrMK0Pg1rShkk4NGHqH8prkfH3hpTQBWZsrK
1TYRKFzK+f2sdQJ7N8UtRjnkhQ3v48nRMxGrr/GUkc/kRAj17Iq2aTB2HY034NU0
3JFQ//nr2lcd7ZRWzoTVTNLgKPM/EeTCimepwCQ+BZ/6XvFxGdPjo2F7s3xORgZa
qWlyte15fyCwH0kd6Y8XSHRhLrYoMHIhHBZYQg4SR8lm/n83RyP5x5Dk3DS9HpX2
hl6pNVqsjzzSu0+nwb7DPZk5uekjqafju+d5sgW7h/NCM9w1gak6Q6FhDJY3AEAj
6qqZmE96LIf/M2cz9yjx1ujqNoSbnBbU5AK5uPuNbtfqU22OrlLVhq+67B31tdYE
seG2nq33RmZqiqPudk6jrJacWvAbr0ei9rbZseDKWeohopkYu0/ROfk1HuRu7ssK
YA+/GKD1QVaLmYMXMHAHchQH5BTll6XsoVUU1Os02iCpGjXXdeeZfK3Iuta2/4K2
zPRzGixSb86Mxfua4ddUc10+O9QQY7rLV1YGnEbuWfdT27uyTfOwHWinLR4XV1Ll
w4kA5gTmcV9H4XZL5nkCB+Khmr5H3Phdj8fzgQ2T1EkLpHUUAYXVLZMAI6cuWk3h
`protect END_PROTECTED
