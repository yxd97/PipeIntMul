`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zg9FqI2IMxwI9t57CoFagP8e8ohxKZerRNKN9y6NGlleTDaim0fPVL9JkbPLSkWG
+BVqvDcVwDnclsEWi2sipk3stciq/x/DBIsffvryAWa0Imu7cM0OlgRvQIfrmqBu
j1kZhZJ3GsdUZAThMxvujhA3hfLV7GbHV6CO4ooWoNeVmTxOog2DbBsHwgrBZjMu
iF4hN7Lb2ImveVWOxv25sEnfupbjYdkHMc5D3HYyG6I4oadFcJnRmMcrtF933STS
fsQgfbV3Hh9UA3mM7E/OlP8WqnmiM6QqpuIe1k7QWBWGEwpvhpOTTetYWWzSVvLM
ig3VMmEi9puroFChMto/UIKxm88slKylwkOQaL+lHRPaRcxPl2w6yPKgtitONNu2
SwFm7YgrW6Q0JkcmYIGNfLkkRxUIIXQZIdYgN6Ci5NH8ZNGubOuuRHU85PwoCYv+
mr5CM6+ZBGJ4Dul04v35ag==
`protect END_PROTECTED
