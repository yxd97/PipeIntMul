`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZZgLmm1CdsMf7FBE7gCSNQ4TjwE/q75gtHhgmVXRs3Z1jhHnTFQ5y4T/Ujgg83w4
FACfJoVrnb2PyvfdfXq3NoEERd745jCJl29I2hvdyj1Zvg8b/tH/zrYY3P3hBWx6
wNUxOB7hZMMi7bgrKoK2NS/v/GxhHqSdx9fFy0DluG4PzBzGzvfuV7NOQgCu9Uoy
CquQkVEhH4AhterN37eQhOuRqDZEE2H6w2FSU0uHJTVRPkFt3bYmUOLPCxxxPD8F
Up0Nt3tgWsV1rQah0zyfesUHYey1OOMozTDZ6Atov2DSpabybDFQFOGU1sLJS5mp
3JfP6r2d89BWKjibF6VGKpOHYgNKqCxnM/afe09SZDtZpkymF3pnCwsK9ZBjigVz
73C3UJ0SVydrZuvg0DvC2ebkGqKKL1kjFkJL+taNOiy597hCWdpG4mJNxhm2zCZ5
LjE2l7li5iJkLlZxBdqDdDyW1eDIVgwDFmgGoBjISG0AMejhJ9OTM0XfR1x9YVvF
V8Bybtbs2QimfKadCICssno45NF0ysNE53HppVzAle3126Sa1cYWbBL9rWkboYjf
kQrn+NEJCZiINA8qWa/J2OCN5NyrHItst9Mhk21w9VZTA9B04o9iIhQfwKdgjQ5q
hFQYzw580p7IIVuk7Rz7mDY+YuDQ8ErYfQ3UAnfXhIDx1q4w30LFlqFPcO4qmLVd
AxwJQfap+npKkQtSKc+q804TdVUUZrRWidpe4RLwLfKiQAXjkRj3USLOEfP1QODI
8No9RIh1tNQ6hpaSB6rWuY7Hb13bdxe2c1pOMOleH1fmhQ5jc0niNg7zs/tU1okY
LZJTGdHM3mNTWEv9nb/ZVJ68Hd1fvtT4Y1uH2RVnvh9iCzD1dFuiyKiJH1QG0teH
GbeiEEenaoP/jvYizUaJlNLAIe//aPsYGHYMlsKJQkQ=
`protect END_PROTECTED
