`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xAA2K3FCvgLS3/mhtUvT7t7tjC+MVtrmRyMn97JZMFipLWIeN5V+lQ4iJlgLp/Tr
D/A5kPEGKu1wGKVp11j7QjdtBitLq4w5B1mhhtc4y63kSO6EBXwix/3lOd3dOAy1
djdN0Y6z7KWwOegzUL7kVO+lHilrxt8PCjrBaaCYxWrzcjqB1k/tqtnROnSnm81W
NDP5qOhPQds8p3AI3kIYXDytqsVITr8eO2GZBYceTDeeH4WqXs6gMeZzID/YJ9KS
irOSg1HBvSQ8/EV9lnO0xHuVYW8wOYhFqU9iZvjAATA8QoyvibakjttCp+9en655
A+Zfp/eczql8+KkWTHRm4lBL7PWFEzYGQWdHcRNybRqSy6wJz5iIHTGU573Z2p0t
Dwj0IIiATKROUaqGMERi/7M9zh1Bcvgul8oJ0MA3Co0=
`protect END_PROTECTED
