`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xWm9Siqukzf4dyISUGwwOuPxYFHK0GvQFQCRA1+Fz4HatdT1qYcj2qWeZ3Q3abFz
x7Iu5He8wkIMS8k66UzUV31sfDh0qfaBtz2nRZbDaKvjAFZ+8pMHu3HF1ZJXPDVY
9mzsMVQnbmk8Oda3+7xrhWYKPPMg6LiMjmPt24tgF1/vxJeeNi56oWUfZYAFfTpE
EbYhA2gMNlq6ffuV56rLoiPy5L/U8+Eb6n1TgISl1X6dfB9L3Za+jVMBOsLMsPSn
VAuJZNl6dorv0kRZgCcOFw==
`protect END_PROTECTED
