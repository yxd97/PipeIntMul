`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vr4eUK/w3+Kv6eu6UwPmQjW+0WGcvDxFm53o/daBAVl06cNkMr25S9FWexY2I+R
YoXOWoLpQBqBlBWmLF5yM1knGtsIS5FhEOoCbpK7MssgNKzS52ejw4rOrUDnFEbz
mNqEjPsKSRveCyq6KpAYF6L8ON6dV+I4tJKFm48G3qKOB/qj5PfRrDc/LIzGWPh2
TkDJOyNKmRcz1kcfwVRgu9SrCt2SAC2rFDrpMmoE0+oMvmodaXdUXqZYJQ7BB3tw
szEuDKhueItVl43qqzi+OGBf9yZk+YWwO9sKz5cUsQJN2I0/eLXS6dyj0UDarfec
OwXwBEXuLjlZYXpS9NQCx5O4qxm0PuiDmafLW7yXQoYJ/3ULjCcK1xH1y21JQAPx
jOC6cok/mSBM/RsZt2HR2uTdM6jARe3g0LHI6Cp98jgWAtqYFsEuTSQRe3Ih5qyN
FU4BLd2Sy/zvj1cyqmoYi2yl0DAUgId4AoX/68NTl5+uUQfepqYC4Q7K3P3DJn/R
XW6zKYZVWBfhDoLNGk/ySQ6E19nbB4cVFQdfO10E0Jj0GGh3SYhHHJQWdHPOQC0d
LqH+UbMXzqOSDS5b0PocDsPFTUe5aFfWl8JDNymfguP1s3RagtJ1Uvs9tkr1QzGq
UE0As8xdUB/zm1k/Sy+XdQD84E+TyQCtL7hrx5Io8X9fs8EpW57WnQj9Vm1N0Bcz
lcSB+PDAkmsH5Ne2shoFPwZ0FSxFIp9jK2/zONbHNEhFybb/X1cH+6oBPxsU9oqR
O3w1MSQbJLIUod691AgMauCff/VqhZV+DARTRlyif1eYJpAo590En5VINXs3deM4
5WcZOcUFv8bGbpAYIYOZbdvYfi3hza1qkAuMoA2jzPCK7PTCEBPS0iM9XEWOiMIl
FbFMmq5xMg92K8Gow2SgQ2hlPPAzgmN50AGi1RXprVbMONCmCLxKwhOx+vaeCPLJ
R9AA0Z8CIeFzDkaYGooJmLC258Xwtd1Vc3BPP/E0iKF6n23y+RoZlWCA1BzXwpFm
HrCqwYTlJob9+3Y+dc2gCpgCpOLnGuNY7t8tdsHjVKTsMFsdHjlnYcYaNgtxNddV
GqNn+GKE07adnBpccLrGi5QN2gE6Qh+9IdmHD/lsnM6Atlml30x+CwnH0BMdVf3N
8wgH6GRTjOVYMIw2sxjv7peg9yQYCX4rUgW6wXTFhy/2NC0K9gV1pi1RPdRqDK9v
7OnxRJRTkMkyd0ZE2h2JvLUBAEevOvBtkP9rdrnbY2WZGEuXXnPJeDv4tpONFjND
EiFCdjLinp/2XVOH/tavZQ8sa18SUbuqwm1V1URv22iMFilx51hzFOXVuU6I7Zyz
8R2oVlXhHFmRjhBT0WYaTyttP3tpKqINwqeMGRW7JbH41S4T8JOUUvH5bW6aZ0zW
So3SblOrv+9UvufZ6LbKwdlpAfAp6keoBjeA1crX7cqy0A5YLF2g1YrxIpNfqPDm
losG1RoYU3OZDEkaToqsqv7AEbpSC28zjcBvO9urQ7Zu/aPMfecCBFqJUED2h17b
iQ35BXFMaeW5WhI2DJmlHLwxf5Yf8wuXXJWQZPz8WvKr6tMRP6YNAG9hva6rOZH6
aSySF1vxJWP3Mjr69XEWj7f1iQQ15CVR1j9aod9z7WiT3s4QCL0dLvI7ntCL0C5n
LodHF1O/4qR1iN0alSE6XQ==
`protect END_PROTECTED
