`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X30UDC4HS9XxxYLDXo9qLgs1NQONZVaRu+ETNplst9m9uOZUAhAXL9UA6D8ajo9l
S46g2ulz2rCslQJpplWcRr2gqT5BBiJwfcsDN0RkVcLwjSYAicDqKYxjt4j5LSIy
e4IKoDd76O01cVK3GRNcZp5J8yvfqbsiQjDLlwD6ZTNM4giEjmvOI+ZlvPl+yUzM
NZuD92S6Rhx6dhS0kW7FyyKVO4k1qMoVel74JEoGkwFPXc3kKV6J4WOK+bZtHfbB
vw44Eexkh+xVBmyWM2Xf4n94tCIC3eMOct4tEKRcbmkCoJGuRsru8pYKU0b1cM8G
HqVjkVJGO0vrzuhdmaxgczeWMYoLEY242g/L/T0kqIG06MZfVnCTHA+YuHEYcyRE
`protect END_PROTECTED
