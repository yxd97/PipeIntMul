`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mBhaYkNxOEGiZbgSrOfhOZvpQ5bDBxBxvPx7eMflZgWd5a1xM/eKoIplVS2GRrOB
S9OEetzF9bLQa6DTJMs41uSEiAR232hnab8F49fzaViDyh/h6AIlvzDQgwNsYkWQ
Qd2g0v2tpfFEV1AgIhLN9tMisedXN/gqMUUGYCvNB9K5EToBClkPDZ/MyOeZZ265
B4+dnql2M3JzcCiqBz2gSfI1dxFg2Zx0pYUFYF6pyvZN3XzUKfOBCpxVWyJDl22e
nRzSxjamnKke9M14eZaWz3D9R3XreVFhBh97BmLiZV5YGDXSFIyN6P8m7Q7ufsqk
5WIkj/JfeIdwML84/pyczPJz0ht9jVpIT7z80WYZCyqk4WyXm/yaIwHBeIwLQ/kx
XZcjvN7V/SaVgZ5UquwQC+gorsjne+o63i5MNzufQ5P3b9p7eoeab8H6B2neao/V
/+4N7vPoiwzmWgsr0boSFTABDZir16BVJEB7h7e59Jg/MryhcqA+AgT+kn4Q202m
T5bjiI/4exl+w6tG4fb+FfJzq2H0e4MqQsWcAkGL12mFxqXyqoXzS/iUUzqKW9o0
g/f7xDpW2TjtXMvmNNVAkrAiGSBA6rlpqlowDZG3icnp0tY2isR1JVPgrWNHoput
XcU6Omih9lKMCvLV5fgvqwn1R4ocl0kCwK/lKmS5F8ENWImRxYTQjSRuuIm3GRGj
7o2nQ52ZY9gMs2KFBrq/gX0glvXBhRQ/QjErNvcxabIqaUEhTcMg/YAfUbls+Wzt
nopXfCIsI8sPW4w/mBbcUw==
`protect END_PROTECTED
