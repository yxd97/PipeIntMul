`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/cN3eSFvCZ+zD27z8OTDwaOF5fdV9f7LRYm3YHfifOrEJcCFXgz9KXCayWkyt2oZ
66L116XLrAebH7qhYDEmLFM+PYty5l405T8vD+yYq/dpYAf9Sql4zpREho5P0WtD
DTvW/SzmdSOKhyAWEaDkzbwHtE7fOGIknipmDxT9yTaKk85Zuweh/2q6/nGd0MUj
9TeublMSuecxuG1N8UsoM2UiSeD2bBlHlmXy7q6P63z8e2uvbS3JzK4mWzNxbQgz
1z+lGyzBLNyhySW7X0Bpcw==
`protect END_PROTECTED
