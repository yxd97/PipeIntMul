`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JxqhiOf9B/OvvS3DKhHrIUfU2yw/0DgdTPb9VB/25O6JqBDnKQHeLF70gYhoy6Ce
PgBAn85OVTAnaRILkDjfusSfMaT4PGVWGpy/I62fP6698aYSW8VodC3KS1ApJWIM
+S14PGhg/VcstZ3R1LmZbv/6WN+6NYwB6UX/2bbzqcmmpWNDzfwTDaa+CQetfqCU
IL9ldRIF3V3oS/jlQG+QRb6QaLTJvwyHpRMwhzpejMhlt4ONcRlgbyB+NhexIZJ+
30TTeysVKCQmHlcnajke5bv0lwQPsOJgX9zay50AQ+sWplvZneSHzyvmVU7YeIhg
uphN49i142oV2X5C8m3zrPXzUVx/jIDv9wQOB5syNUpKfMvQD2qvwqFQQYizJn6O
gWsinn3+nQzZ7V003nL8XFZGKshnCW2g+EqnB8nomOL4fKaG8qohB/E5VSB1ClWQ
weQqKDn8hnptIoMoayL+uUolmXRlmYffZhcZ26/fDjVwFxQDiL1e5eh0kChE0utk
O10U90+VyHKt+1Qsl/sAHV/07cBUHpD3PqYlUCSXVI2H4efY/7umTkPn/o9MDy7T
u1khDL3eIdSK65CNgRVlnVZ3WjoScAkgJGJrNFbbReg=
`protect END_PROTECTED
