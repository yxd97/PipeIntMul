`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XM9dZz/fDOAe8NO76cTmU5Qv4rYgwYRrgvu8Lj1i4KtJcuaTHZt4z5p62mBf8t4t
/yevpKEZ2Kj+FA/F3eEeMJA6TmgakHeAFN+ltAvS9Q67LeWhwU/RqCXUbrGPeUCd
huqmTLRdy660IPGyovTP37Kbe9VD7KGAWxW4CuRJDq6mrX10FczkLUsJf4p3dsiR
W5PF9homj+SdhtkiXoPsR24sAGGYkl7YYx9p+VQB+hxPmLmzaoFsalD/oQgKorfG
hhpxZbT/MEHJ9eAkgsMBCUNDAj/jZB19Mm5Sx6cabgyNfrcMbdB78MVOkWqL+prv
sh1/mRRZgklu5y7pQs4EwdRRTKk7UUoeGLWnVN8olgsaRwQhE7s7QDKoOofzhWRH
hbdzB+KtugFqLWMpD0v3sZbxOi6q/gXtOWPeg69zv5+qvHYsmhzz4JpxL5vW4sRa
`protect END_PROTECTED
