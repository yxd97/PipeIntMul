`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v6LPh0u8aWM3Zl/hEfTaWPnJ4++bhZFY1WPyglXrYh474MRCrVve7PeHAUlQzYNY
apzW7Z6b4qAo8i+ej3MajmQp+swcWmaqr5slDzn79KgXMz6UlNV3fA6oG9wVTdWn
S9MhxwoKeFBR/N+9lAZFUwnJyAoYMYRf33ENqk8Gh2TsISVZixERGzKPbFOTiGEf
LF8rbfpwG31S7yTATH6FzBVTvP6aAU4Z7hkSkGR9hw8BTlGnGlkT85eXCUujXSDR
60DySrNPGwmRbOdPBzJJkg==
`protect END_PROTECTED
