`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xqI86prwrT1Q4Q4wKJ4nITE9e6NlfJHZtZCCKHdVLHI5LpdI9jyZ6RNXLduc9G4
qRNP1+35wRhVwtUfu2WA67lodHsTMAf7G4/F0+O3xoLHjIiSHiZ1gw0kcsBdY6mK
jDtTw/iS1FplsQu9FscWcfCeSgbwIS04Uotc770/k2TkCawlgEkoc8xv4JvWYsso
A2UIT5Xj+Lra4YK8erTWlPmhu2hLxa73af6rUfAFnLuD1NMIx1qmikcqr6QFitts
Cda/ZOH1VzUtqsSiBvsvM3drP3R++hyx7XfrNe0n93FqZ6rkY01qz4E9YY0ZX4X2
1vqV/wrp0B2NhLAKLmcONsNb4Uji+maBjbUzmoz8qnxa6UAa563/LGyWsqYVFHYE
pBNQLeQAk3Fcwy2hKtUQOK5A1QEt4npITedbwKW9Vtwarct0K80xJwbC+9+JBNtm
Kv47vAlXCSWU5LywWfDsiqInyNA9tzHwskv3x8mYF1h+/AG26HDQ8HVJmWl8hN0e
HDtoGd7ORVMoDXGSSJlQd9GhWJKu+MCOqFkjKtA2ApI68EQV6DRkEGq1/JnkXNJ6
63q29hcYcj/yafyh4B9afeIJt8ne1viYw+W9Filr2Kbjh4653P3jUyRURdWMDo3G
mYbUHtLDw5DkcKCz6a5oY0+SpU3sU3BfEgtUpw/+h744XPlr91rCEsDDwx+fUkrf
CEM8eOjjOkM5y7f6OWzWW9ocpfuXbo2jKinKWn0Hg56SIyE95H/LrLim245wpEki
hEthey9aZKXYdwUbVQeZbWWbzoIGw2li3sJ5e1VTt0QhaM+buHemjkLosG1RLZxc
l8xNdLU/tCCU6A3eQMmDGI5XzHbn1O8IWWpyWrZrmOIy/GDtqeR0mMCE9tQI0AkX
UxKk//h72rzz7xf+hBusrTsHp0NN0qfDHlb3jpO5rOaMVYZBq/JRofWI6d3xlrJc
H1QfciS0JSA7mKgPqfwKnAYfLH/UisHnCfRvQRGUeAXPkItj+IpolJsUNBxM2d8r
WETGxT9lXCgDAqYN4rklbC7i/RO8JDmrHNWVGATdJ5P4R8Kq3Tn+7ZgRwtjnZm1T
FFZLPAeo9TV1MGNzW9LydnfKRUPMfQpoCJZwHGSlDNLH97AJqUfGV/ydmZrjpfqd
2ry6Gnce9qIcCmpoAABVz+ueQi1o/2OLanG5EeGm/rlJW85RwVNCyUYlrL7cyAat
tcKWzaSBCJ7yEk9Dkh5UH2Wtpbpi7tzvRRCAlfXljtTeqt184CdxPUuHuFmEpoBW
rtOCmo11NgJWPpBX6zsQ5nOB1xR3a+kxfYSNwF19FT70ilgOHcQZLeMhn086O5ip
W6JKdzJP2U150pgz6IK0nlcI7X6lRDT/RojgfBOcqAabhCaOg4zlXiAFs4l5BA8g
Vz3JFfRXir36pUo9SEA5POdIR0Xb6j9U8DAAY7Ba9n7sirEXEzuuzc6Lrld1P82k
kcwYlKUqKr9FQvadJFd4Q16FHcGje70Ik2rpQY4S8d8MHysPSE07LjNNYmCnmEsf
ncuPXiYI2zjHJMFhagwZSCJqReZfvhiuZNQiWVsYnwtrtsup1r4yINlWCQgcgtTq
qOhav8I35Nkj8Rw1v+BegxflQk7pyOj6rS5YW5TN8vS2Fj++ANueB58S/KpT8XrQ
P8GIFxXjuIwWTFJ6BijB2GpRFVElX0y3dQzJ3tx2Ck0C6yJrctgubU2Rf/MbunXC
bCu851c3xuK/hqOBGEheJnK+NDVFAj8kPO4pfwQRz0E4cOq7ZUMGPWWheCOcd/My
5Zyu8JlLaKb/uyP+S0KKBUe7mBmzButxhU1f2YAU6SEOrbdsoaYnxAVQ+5pRSTYC
frGVY10hhvhvuSZjhU02MkixT9+fOH+XOtRSUl2UT+e2aIO3K/hucEZmzv35Eav6
ncnqSY35X79oTcqk9g9CRq34X1YwVhW+qz5ogOVW3ExYwl+qYe5pz4PYKtGvWUTX
Mqu7E78EXEX2gBecQIcrlD/II99YWucEQSqzkvagWt8Mr9gcovCxnBzbRF7U3mKU
jfaFfu89GW19aRIUlWkdZiutzHyCkyl7jNOIewR9IZdsn5v56BPCw5vc1UCrxPyh
0bAgKasI8v4op9jhzwrRH8UKrchzIamDY/7HRqyIH7F+JIvnInnkN4oFDNFp5wVh
G+pt51aGBKnfV3t7W8XCiBkwCR1XG0lcGMhvFQI55ekMv7YXK0B75yokv/Wjyw8W
YYcNz7t9kTK5IQvpjEbFDgZzlpeCXIgGYn3X8t6yL201smZf1CuayABf7h880bLR
HE8d2GecEfph7cL+05N9mp3Pl2JY/Y3v+iQ/HsZzArzSnyfeonZxLTBW1iYpYmjC
6EK3XbFChdEcXL/vFYsi/O+/ngl2tqWlg4uV3J7SX5ZqDuB7fiLCFGwKhopRbcqY
LNezBpJ3g7F0oS8UzLPQIRLtu5fJhofCEunGKdJ6Yd8ITzCnS4aD8h0gyM7yquks
So/GM551IyxfBZlw+kypmQywlnNT4xvEmFGJrCNZ1ylg+ZDHrSAlkEXXIXGK/S0G
5ZTDE40RCdqL813pljKJUOcQ3M59nixeckNbjoiAa/jFj+q7vSpdu8braMT+86rp
IhzJnzSlPJRFhLPL1dwbiUkb9sBYHyYNZXDRCLzvT4zl03iRD8aoMDfiW061OggM
n9+HvygHvevJ17DV7biSWIpXPNF8OEVvRiJOspwb8nGmfwnO/HYz98ADRVbqzSs9
BB3oXK86LWS0rDUwp00sNBajLFYCqMRk2hShJFLEGkEwOy6D4Dz7i3VU+5VkHjiy
Tt1B23rfkW3jUH3SiTk8r/6D69fZi2JkzPRPtUVIiapO8s4mZKuILKR4h3T0mEtR
QcOxaCCiIyuRs3/umU6uPf39xV0aXX97Ba/9+4jDup23FqdXLlVlYtWrGMwoBG6x
aKU47TmCYdwB4jBcvXczcVdxffFlufBgzIC59U6B7CanYpErtRIgHLr8r+bZjc4a
wX/XF+MF3jsW4JC20/PYFVpb+DVIgPCJnkHFVaNgKjIS4/aptg4oBZUhH0kG6xIL
SV6+sjjXmCfAj+rQCzUyUbUU0Na/6yGjJwKPjPVyrQh22Qw+X3EpctBsxIysGP81
xRulDYt4hGkyqbMiG6iGAn436CBpUyk0mxe277P2Vm2tjSnP0tk/Zf0gqv3B9rLw
JmYWT6y0hlH0PgzCy2sQsFyrYu9jKwWDE9M0grKLXgQmCE3ePl9scqCKao/vg88h
k3AdbsIKZOFc+yWBauxfFpo5tKrRCCxWgkt5EqioESup7rZQTCmCno4FIQqG/lZj
tApJrSTlWxAEft9FLA+UeiE1RK3Gf54MRL6NE5bwUkhx8UU3rmHElM7CBo/LN5Lu
ugGYBS8Hp7PCQo+WfS85db/yecmyjuAXtcaUVcJVKTxeiimZFnoKYQzQyjU/pTsj
lqJC/48LEiwRkhtF9hC3z9ttYKnDcuA4+4lg/kKV0RZgiiukIWO+EmXiNAH5wtp0
4S2ux40yVfUsA0SlaXU+vNiPGMNOgJVMJIMLmghZVYbfmJXWYo6kiLYBUU4FWAdl
we/7cM6k8xeEOqwert2ytwM1zTa/4w02Gcc3aziXoKUD+9tUEa+4sDb5yeX0A1TZ
itTvVQVpKLSIBtlab0GsxiWZVJcsQB7sxtiO4miQvLSJHy9RCqX3rLDaflsb+Vw6
s22JzW3U0zyWdRVzoxwY4q/Xw1T23fwbMqBzKOb2Hb0BusHVYJoRiuK/qZHnV1Ws
n7vYjy0B7lFKvPh6unNTjizl/Haxqxvjq5UXneg7XTTyCmWPRK/lOjUxxUPzDcHN
BV7VqhhuW2ZhN/iBc/Lte9OMrWgrue8z5w4s44h2mmQnFMy7dwN5LhOoqcZBj6aE
euvJQ3M5Cy/q11mvTcqyL8kcbBXoujltEOhSeWbUtpML7qTHd5Ae384EaRyMUA8H
8IbKXGoKNTQ73v6XyBqh/RnA2lK6ezDw0xHJofc5WS1ooO66FctMZ53SOrzKtaMO
6AetR/DsoKyEhSQA6Z9j8GkWmarlPnN79tYtK7rFfBBgBa2JU8JVFUdM46MOhMyw
nf8tDxVimrRZYVpL9RrH17orz/1PcCi41nFaBEMefIt/znvBmyP9oBopJoPx4Qb3
ZPbcvo7Ma43HVSxuJ4q4yfjc5bTXGqcnT/GKzAlDljLiO5alJnBRR0qqmDsgxEfE
tz5BhA2KpD0wcd6JILocmyEywkhM9XJwfTi+Q2OkAL1Xy6nQglIwJxlWUx7PsmK7
lr2JJV4Ajx0XiRtZZmuH3bxGjCOsFkbHcPjuaC8GbflZXIldR3Dyoxw2cytKBUpz
D7F3PtNx4kHOTHhg8t18axsodSVecnjBWraGje8RyyHzVxfQvy6oGjWiUzw3UPRY
Pui9g3w2NXlkFhFGiVuLET4icLK2+FSY5nMoqn+cWG199j5bvH9MBQuysCmzI/9+
qQL0nBhcYpA+Ktt2KSSIM+LP2HBqevjkiaHFZUUJciG3ydtfDb9lE4pRuDyyP+sC
GOVcPYl9mmD+i13oLNc8riPQKJqznsCYrQpasOQtxLPWkaNJBwWrSP2yknhVjG/w
RMvPeSVn3Tb+x0KkdirY8RDHM0inoJETKcMnzaNsHdZrsHa8A3N+uNhmbnJ0Uyq+
9wwE6zOrYKrjDeIJ/bBNa7lxMT4LxCstIUsUx3u5Fi/xQeVBR26W1V1/jrOkwUax
AWDfBgzgX/IjR4ztCmZT+Piz4XWLyKa+ezrS77+TpibO0jVrs9aP7UbD1u1DMGiR
OAhM9wr7ac2sijsMVGB0lTQVWgSu8wd+BmMzf2zX0SpsgltkLot7WPOeT4LzBqfJ
Roe9bd6qqek2fsOzbr74cZD1SAQ/mktWd+OHcg4Cubg+zu37rKrwpM8pRH/+wHou
nKs3+34jWuegzN3rLqxdNdcd0iufptO0s+ZHCTnpiQukel6ZpEVF4GwOnkgQrQjt
fv/IaJTl9BBSp5v8dcnE5zsHryjkrt+jIvzyceNNncNjjlzosdMvH/RpqfOHnIkh
xKzcgLfbrd5L64sNtXmIQCBwKoKggxMy46RAlyO74cNYovBrJKoFx/MLM5MaWrFZ
IzzTqf6Oo0HUGJ9O1COUZXRcAZT/jgLw/bwfCGOqR9oMu1mD3sH84W+zV7KPJIPU
dspH4tB8OhNy2CgR15sM79v6bGbiVquDGvIRrd9e8ehr1YtOKfDRRiMXUfbszff9
Po5ctSaaio1uJv4lY0O3zuhBjo5lbbzVodUa9NIfoc2RvdkNvIl+BOSx/wt1dBNe
MnsTJY1ZHJisgOrH0hk/whFhXyFRzUMcya1bwkPraP5YVOhXF1RWHzbgUpeFKeDk
D5Z0ggcPsxkbGGvRtX6H3qOnz6deKBzMNWPQf87l28umYdxK1wlAgDKy94daw4Fk
1EocDkm0fNSf1R/+F+xqh0cxmUnhn5vD3dqLXUi+BCYb6heIiiLtDugi7f2iEJ79
i0IxFvKxlm4ZjUUzNRXwMbGi/ynGt6i8zd7Gy602f+txM3cRvgcCxOe5IUxHQVTO
GbLpLxx+PevafnyQoPq+x9F/pMP6lxeCT0N77+MAhTlfKo6tlbftz9bqXztVtf/p
bEQp4ofPUjekiWlKQdPWrNtUIzUqQDoDvLicfH8a3mXVeVP297lSr11UtnGZ2C3Q
pc2UZE+1k7kTM7Q+N3rLI6SgrocB8e0PPfuY7o7vsW3lY8IuqfUJ0kfp1GFOCoTA
8KoU+DIMMhdY50jnZk5uWlv6aVCEdNm+WWxCbfgaBkI6McKx2IA52haN5PbzjM2t
1ykBv3xc+aNlYPWmnBT4UJR1qT9zT9fLPyFLMpno9jQlbLuZiN4pKc1YKdTeyL5K
IjFyJEy+hL/j48wv6L0BtQqYAf7coQo5UDmDeHjQOIACO6tS4Wd9P8qm56YnYVvb
dCGKQVGmV9upWHPTHckidrqauVGZzri4s8AlJLUuKPvziSpI4DxQvwsQbUi4bCwD
c3Bh5lMxw4SBViMVvbdwkK63o+wPFgnoz3ndd+O7ZZdSLaH2XFDWoo3uM3WUMVP5
wFWdsoQPpGV93Ksru3NwBQTtGkLKhTIh+Pj80J2BDs7AKBkZdFLGB2WRv6SY7ZdW
0wmOtSeDX0ihZy3wuZhT1Rd7ORRM6E4NrxZMGhy4dj5MtH8Z32NaDEfINapwmVcb
QqrQWuOs/4LAyMUdvmJRKJbBSn0izC1SpGH2oOXr6Rrkto8XIv9ezjIWXmDjEmY9
g0L+qaEs3w2F/MMsAWdmmfNtER17w0MeBGua9k/Lx6sc5zON4gRo628C7Jluqrl0
uJeUBYHa2r+1rXFL7Jm/MrCoKUBAJ98t529tscTrgUIn+GYuqrT949NNVWKzJ64K
wmmYlxojxvqOD1am/kqks8TtN7fgs0J9u+YP5sZiDuq7RP/3BcncCfeNMbR/eePm
Kd6mKR2Tn9vTiqJro7bk3YTvRwSupq9SGkhRwNRwoUjuAvdLWAXUveWYjvPWzxOV
QHdlKTkOC1NH1ArhVpbK0QQAhItDi5DWaK7Ka87CNyVwUoBX2bb4DjAlnihx+Hi2
AoAEXN38w1iPbgMjBC5kmu8+qQHvXj+mM/Nt1nMJ7wCmgyZsxRcfnTKZlNox+xWy
CMvWLMd7LOhX5xzw/Vy8wfDyYNwG3Xr6eujUSbjGLwhJaE1It2lA8JPT3mr/mCeJ
2xXSpobDV16y87PMhBXC2seJkEbk507sfL3H37Bex5yPxgqRU22IWVY0+q3WbRRM
Hu/rPSD+sh0cES2qT7X5bTPeryZKejhW7yukyg6xl4itnjlV9Y5H2VG4LTLLCxv+
SEU5kE9RPSZ94HTfyOTIO6nm772c8s/hfT7Gh0r7A1n7ATgAjpVFICZNaHrV5F8y
QvXCjNWuWouEVJift2E00pP+MxJBTV+/rWIg2d3Y2VboZDEfToqNqsijgiQ3U5jW
Q5+iAKmx2qV5ULQHg01Arx/sTEUC4JMYvRjAVH1WFY0eqcnAY9KsUP5Bv9OEq7yQ
FGI8vNuFsAznB0bOc3qv6WvFomM0jvbrool5nVjB5HRjLSqax68gk7ufWNex+KEc
rmpVY10BLxzkjNJMxSnzYfhRlIMhhrIewNvt3TE3faEdj/mf+qgHnT6tj3otG23e
sem8TZC6TWybyAAuTwfiOmVnvO64NarchCSixGoZEakT8vwuI34U+W+R/5vDnc5z
ja49WLfxWxeTtAiAtAG4BklxQPnb5G2eDZPF75bKInsARd2KNw+NyiDHuLjUxnPw
QdIReMwoawnTpl+49rYzVWYEp8pP+QJorEWeG4dfKpB2G5Lf1XgCshHIZHfFiFJL
gLmaW5xddCZlfaqer0XfHjFlKZOxo8W146ac/9+rbtlyNLEb9BkBBwPLa7JxV+nM
P5i6NfmAqXWPRX6m5aFXnEoWI35kqxs/yNLQFVRK6L5zEeDmpH7Nd+G7oieFWho+
HbbYhnSm2AZHEUppx7uN+cHyIcaArXR5iVVf0mC/59Z55XZ0pzE0zuvFfFXARUiG
ZlxNpgMe8UXyFOkrHxSQ5Mkw1SEeQIb5stZSk/OkQ173YBPpVSwxpLGdK24K+3fk
2wYOgobwnf3bvwHtbIoODDeh1gaB/3OxQdgnPFJUiD0HFFlUAp7vYjHrE3ZS+Mw4
5JD52V/PShGbPPh0tW77yNJYVNJP6n1Za/SXJmwOgg0Phs6f1bp40rI2tkSMdWo5
Tkt01fgDr3txw0hA5BQ/BnJtCPLSmFibLb1nKEJNFHHnbcNZGZ9IFiXAzZmDYx8n
sPlS0WV5ys7mzOtnSfNDXyJ3ebVtKFTZvxSgCD4LxdACQH3cCYzMjEKazpMQuhjg
pYlWMnLJL+AqzouTq/ERgy/FbloHOD8P9BZx3aqiXE5aBbnTKkFLJawdlJSw9vj9
3iO8vEsdjyMiMdqWV1HNfMGqwpHQ/Ul9Fi9x4UYD5R982rEZvtNUNNgkqcsdAHVr
PE60uCsel10gfHLeq7GJUvSClLMfkWgaL8oQW6m/p7wwuVQLe8ePEZOYHFr/08Xn
32j37u/zmbHLRlKQWTKk2oNtjVhQG/JDfWyxzWJpY5+g4RS06KUUKp3A4SMES1Fu
yt260ufviFMXX0QR9VGeKK56vbotA4wewvval0jyvpZr689te5LBtdKox43b2dgm
/qaAbl9x6U2JOHsVipmvN+TmGbazpOXNEds9hG71ESFBQEq0VLLyPP3uzJs8ZZLF
+q2amay4+Bw5C9Omt2SpZ8HKquxtgjtFRY3RcqJbztVhY+ZGpGW76AZzuI1LSIpQ
cwQRuNDex/Eucvc6UyCXkycWGq1ocG7ViIXx+PigwJ3yGkAkoGQhnpkBJ4AhWyUl
yZLBNbGpRh+NgbM7/Aju/zUZnx8WT9m/PfzT290xeoV1Gx2aM5H377g1IGRrMSEm
pjD5WzfE5fX2knudmJtMXhCPz4HCVHUjw+seDPekkTh5q1tKKtuhb+PK2ji/8zqp
SnDLSzEh1310obCNx2Ctwqqy2P/w6aiLUVNGmn1yLdxCQiU2Hcq9jYEdiQVIQbSq
JnQdqNeJDtrTv6w30JqpCmfTUkKdhZzerdTlj+0nfyRInURATv3v0am3HjWyi+jP
fUgWfOUmHrGm6lSZG3aQ9JeJpfoJPB9rqP5Rww3WIDlrqUu9T/5V0tReux0YCAXf
L0HHmMCzULC/rO8Rvzzo4lhILSj2WT0bHW4bPXo0RLilrEsU0ntYo1OmUYHRMpmJ
9SOM3i3d27DRI1zEh+DLexbwNyt3ecPk1kZp0v23/5HLpMLF1k8f5DnnN84qsPTM
Kx5Cao+jlRcQl/w5+UV98OTG8wdYChtuvdbe/GdNDYFzdiuOMq3HgoK9vjRwdILs
TH/T+Dv4cMIkyVyxxoZzM7Sbe76XAy+VEtPBdeN//H0c4w1YRjOfObwO0JM2DtG1
GDpg8e81IOflMlDYpt83rdIS2hWK0FYNL8eT6994QMXLhyxkp7NCWNffmNJG0TlX
m80YSnm8RMREyKO/CHn9xnPrkYPtVMyttXxirxXswMYclkqWr9z+wPPgCxsWLIqM
GE9e5ngfzsi/qoNDPc0gSkLZ3F6IwUtLaoe42SzSN4vhK4avAwBgZNLOxH0G+96g
mbssLwtWSAjkltSvMT9TtVmo87d5sgRuzsrt3j/UiGrbbj6JU6KcCmeQmRaAqnp2
lCgL8sxhAt15jyPgCGWNX4jhO3zBstg1l1PlOMckjQuCgMX3mKU76qbqFGxOEL/G
ak7tz0G2SpRiV1ELt4atGD6AaqeOFtsaB10LMCTcdVrLIarHfgmE1swqJ4C938/8
kFPtB/zW6EDuDv0NQelhyznZ9WBXdHDzCjRwrrl1mbAS0lpCR2E4ipWyh/swiZId
HqAdvzDKclOHWEOvGMU8Aw0w7pdIdt4jX+fTXTkBT8clkN/BYoFASZpyy3O8FGHc
qBzVf3WMRl0hHiGy/Hujn1uUjVIce5w+odOlwfUU8LShGDl5TEk2yW8Bo/C79Iu2
H/qLZvxo7j025PtGhwSGVqFQ8oeCUysJ0BtJ+EPRezHuPm9SkVncE/n4K+Lz4Jd8
a4WZauVKbCFpSZRvrCkjUR1nUoP2lGITlfDWqa0Omxsk5TXekNLcv/3sRaA303UF
blcQYOO0faTn7W2Y1N1RM8zWQTVc4nvMxU/cOZdYLJOdqOrSqctW7RkaaiDYNdHk
4ELkaiW4ZMntD3SU4BxTWFcWm+QBK66itScSsOd+dAy0IgZUUKDaweAlSArzI6KT
wR6H2ZYp7GfLDVF8V/YL2t0Hd0+KH9g2dhbLJUnv+/H9lsrrUGfun0DI+g2q3HPA
IMEHyaSVbfkbQT9ZNoS8xD7njsKg44XjDWrP6ya42/kCp0mFq2O3+83ODtLwyRYi
Mii8ALOzZWpRj5ZHNKVkHnKw3lS5z795a2e+SaeDs99fQfLZ4fNMMEjgFqz9jdKI
OZ8WFI8tRNdQNrBawGC8ELOoMz/exA9E9WliFEoR4/Ee5pLgO5chvfhImIiQovRw
zrant5G7Dcb5y3XmmiVNUfDApBsHCHOgLCnEfKwOet9XDtf8cfbfPmXven1Xl5dD
JUglhOoUWNhTw70ZqtaiU5bC/f/w4G7T8EiktAsZmprJklzDAYD0oBmhbLSvZoRe
XG+s3gMTLflHE7JjCuFZeHmPsJRwC3yE3YvRQsHxkVNMgHdcdtor4JONQD7wmbgC
oedEUWFTrqVepLwNBt74WE//GNJxkSSvLuTsWo0DMPPV2jvVbltSFPUDiny3LfIZ
ySGT33dHX7FkyYl87j4HW2rJa8ZZ6ZAPUyr79r8hOKboRxfZjTroRnkhrTwYRf4D
jXc4AgtM04a8lphPLSrUY4i2ZRgcWyq1jGvv3/+vrm9DY/80KFpd5Gddx2leFyC0
cKbKdfqdaTqxJSsRPkkcsXXwM1ueakbt3XLwcAkV2FPtB/LmOId+dg8R6weLVrp2
qHdFUHgi2kBOz1s71sDtGZStwC1alUeLA3pmngyD3kCcNVvgLlgPeXJgywoQqwBq
JsWh4n89+EVWlwewCHENl5bpoK/VXmTQEbBoKQKGTGry3WVjWk5JnT5SpMpYI7Ey
pm5rycq4Hzjgvqtbtyc/9NXP7hejrU72LXXOp2K44+90YfXorsDaElZThYuTXykH
hnq1D/Avf+6ht+3R+NW3DiU6UZdb+0Zd6ISzFUJKVf5to+pqOrA30z44wKBohZvx
8kxLs87KNc0Z6Ypx5xSTvCxev4glqOCYE53pQ1iKzlrKXKkQ1em7rW4Qp8aKGU4Z
2pyTpHO2mF5RvKQCsnqA8PrJa+yQiN66LDp0j2fkRhmArar584y+yLd74UrnPncf
+GM0ZthX6sB4K+/1N6g0AvjeglFD5Zs22wMuFtL0nNFFfaW/FKBXqIiNn/GGavq+
HSYLsr964o8M50fKdGgI8ymKtGNWnpKUQN+MhqrLr2TilKqHmBf2xbg40kCNICay
B6oNonsLXDZDhVaVRvvJtO4NdlYttjzQrZA6R0LiG28qBkx27NlGRwoKzME0Ph3O
71vlGIw/BUamqC1KtrcEhXmGBQnnqKFjPIMnPksu+Ddtg/I8ur6+KP7bfHjieyUs
IK5e7rH0fN1L2c4/ZWgZ9jyewdG67p9UL1PnKfhwiEfaxJ6ygJhQq/ELdhpKgyx/
w6xnEmMQeqnb97ZlbXf8kgh32FBEQ7h3f3SATH7J7VOC+sV9/rQfe3n2B+3DJaBQ
1NwifXrKpoYwPJhsGV6z8XBlUJDGJFQYRP7f9b3JHxtQHi8JWvygCV6zE/9dpGdG
iiOqB3svsCKYB8CVYRpIn6TNYg+V0C/2+UZS3+Lx7tj5cpeWaDhbg1m4UD+GFkiB
U+iulhMDDu4vU7OReSuu9Jt47vZUXiwkVca0/HTBTOBE5j1GswKp9YppxjHasuPF
2RNljNk6DEoanoHgm5c9JhKiCdy8yoNP5WEG0t8xzPFB0nCPX9auFbwsj40C6cAH
QJzbhuN7Mn0nfMN29COUtpsbLDu2FiIifct/cQJ7N7wgyI4i++RMJXf1PWEGa4y7
DtcQMZo2zmx6DfxqBn8fLKf9kxUz5D9HhKgvi9F9ApDXvQN1GZhzfYDIhb4i4mY7
sYrJm3+QeI1Z6g8WFj4uO8EUM8oJ7N22Hust8vPu3UWw0RnDZj3zorR/04Jepyog
yO2L3GUBKUTWAilgWvTmYn5FC+65zOcat8q/0tLtbbMVgsIUA4muNg+HWOxcTHcx
4qCZ0oM5xc+49OPR8cKm9zD5S/5ay/9IwLTuUAcfiMrZvtypjmbRZPgLWGpMunGS
bHKLDGwBp9Ay23fs9gwiBKQyAsDNn12OMj16SkRW6E8p7gZtJQgvRHeRL0ObcB5F
TR3A5JcpkJPezTIZERX2efZI1al0CCUxgDthbQTwCbWmgQcDLhqVJPlmWPm5MnHa
Iaju50Z6nQQY2CylXv+yT3apqjOKRvChHgt2RUM7rdbyJgFEIHYwnkwFqW/Iv3Ny
pxVNFETNDRHCVPhDafQTwD3xY04bUHqlM+5p8otWx6crYd8lb6ia+YsUFB2xYmqE
X2VTXvgRbSuNIu6q9k+rjib/3WNIg409o7ehRiFU/49GLvIWjfZCjY+l6UkHG6nS
XOe4IMCfYOHqK0ULTXV6hMyjoP2ylkzetTYi8M2ysoI+FlcC4FICs4mUUtOhZrH5
BfFu+Wx/hoqLMxq3gxLra7RblreYMcQl+rYRbAx+pJOiG58qPmNw3WsfZOuGMxir
gttU/0C5lkO9GcH/rLFIT4UoONSYjmtkTFLFYp7UZsBkvff9ZH6s5YDK4P7NfHX1
5GsgTt4RRLRl4Cc5x4yEYaSFPPICJCwuxBLZfSklzUK51FlBU+P+Xp+nMAKMoyRm
5cEGscaRI2Tw9MQFQpdPmpNmiRWGHa+UNMNzVXe9JWVzIRUoK5KmAWz8P8xAl/7E
vxFUTaexzyrcbqVjb+YYO5v4j6HHHmpiWo+RjfWuewJZDNZ98NFbHaaKLX3axbKA
qRfeVuyjxAbdwcJHp0K/06g20WA7d6gvlsPxJ4RYOHym1X3E1Tma/NtU1nBhs4zB
mdJHDkZBpPBCDax7EaZkytDMAUwn4sURwFOXkUZgRK/FvlMphme0hki2WcrVj9tj
QHuWdyIr++6RiEILPE4yyveAD8tGxiquZUiH4sufwFwL3mVF87C2P/mks2NZT9Aw
/kK9urybo3UovpyH2sUadmYgzhs8NQmNAEg58NZUYy2A8uYf6pelmVSd0T/kPT01
Fv/w50yd+UEGiq66sT/fBQHCG4GU9Jp2VAckRbf11ABbBOHbSVNbWO2qQ+mZupSi
iGNBzC7q+ynAXjEP26DP8ZgWAb7qVebgmiod9wCq46IS7a3oSCnH0OhTXXRLL/CT
MzK1Wom15OOzLRrzzaGgPvoJHfl6+l7xiDIacbujnOBR5hzTq6bqQ73hIZIeiSMU
s8gTFT8zmXEUKahc4oSo0soh/8uEzSb7ZEq8rmPHQOhTA+orcs43m5elHE/F2d8R
OQBDV4EEg0sgHi0s7OrP1kf4qaXevPV/53xcBHXp9TfSiFX3As+YuQJ4zAYj1knt
HCgnIyLXZAPXF3umUXww64RiyA4Rs/hBwc7h/PhxRGMH3STd5BSDNHK25+vPN+g7
F2ZQXPd6Nxnezu1KfB7ErNF4mz6BB59efWDPjm4whf5NrqfL3/+ZZ/6B+jte8j4S
5K41QmrZr5JrI7bt/XpRqiglPbZpSz5nbSkhiprvofDtd38IUR+jaCyd1lm9gO0I
H9On66CI+04HgS8VkXq1ZAPxdNW59WwmenVrZ12zItwwBEB7MBOBshDksZcK2wR7
AxhbT8w9LM5nsF4w6wFukCB0s+Z5Kx/yaRMu5ZSUocQcm333mEP4mX1ngLblyF8e
pNNESOUd0SrPCyeZIeTMmlxJukoe3OzFeKLCyaDllKjOIv2O85jftiUtEwFXL1e/
E8WGHCJfjM6sj8efl6zS0F2jVN4ibbZjLjCEh5UBvwlcqPt625GrhqKmOjG90L0W
b3Z1ojdc3XDIhcwlPOyGKPn577fIaSkcAx1+R0xd2Zmdy2iCXXz3Rm/fqedEx3nh
WmLyXTZvt3467wCMc8DfBka7WDhI6nE5DG2hpuKTJjCjg6CS+gXDFNba6deCJBBb
/YhC9kRwOsl5ow3RlzPDno5EHNnwrsIsj8j+zJ5NmEVeOHRx0iD/u/sYTxB4VOFz
8wSRQQwjIYm6j2yi9c0dQqT8OMJtgsU2QCpMA4IhfBTI9Z5lXQaGD8j4r+vK+DKe
Wpgz9XABQDEJU0jEx1v1p0hLMem7Tv8pNdoVgm8Z8boLTWZsGYWBqwfG6jqCeI+5
La4eHwfumISek2b+B+RfITsezgr59b1qJXsHR45FXjuY59RyzZi0+wd7pvmZtKZt
luMkeImjR3OkkPG1HR4CHFof3cjt3fyOtRVLqMpIXy1oWqdqHOV/KyeqZtHrVsM+
CRyB5SXaBk/4Y1KzJwsmmbksrDB+zut6UN19kuur7NvvqPeeZKBq+tigZJb6f3WN
C9lj3gWNjFrVi7DdqLrJSC/5k4ZEPWV4fFc+T2VdG534p18o4FLtfgSHuim9kKT6
zHPJPTX6CMAoj4aLA0x2ohajamLSfG9jAhEcIGBbG7u2Wy5wGPusrNyB9HlhTj5I
HhzOrcMCp7kJXabeaHuLCMxU0Cw9ytMJjzwmnyVpBJ+6HHSyhoKPpbhhSBRrPEsn
MrzmDUXlu39KFuCL4a7gGFII7nT6KdnSzfraYoP1BHAAmJE3f+3kscZ2mzzPTvJ2
dPddEP8Ij623wEtGIsACW4b+2LtHvUBY2iF2LQZ8rZktrIudiXaBZ2YXh1pXfNup
QQ09bycWr5xgcMV/qweJ25uOgUuhUpcptL5jTPH8sQdAS7fjlYetuSjIt3S7cXpW
/QSBD6X8O9BjJHfnzVUyvvBndREEyPUmwZZ5nOa0CD7EGs9M0ymJPjUPeAEaAD/1
7jL525qi4tISQIFzf82qo1mwniJVVd0Vym0/051uYNTPLYx5MKr8shgK4uN6EnCy
3lEjL5wTO10mkj4vHKLVCItRqFSv37iEKUxessqUPE0tsh8I/9sRGTyc0GmZeVp9
84UBPqcVQRlS4EK5LtHwiZyjycKWhqB+V5uhr4yVL5bFzzd2+unmCHBeFWavPBFy
8j7uV+Vi7HYPO9xbpvgthwiJUxesIFwHBaAHAXySe6xsItAL8l26iAlaNF437d+3
FkFzI7zO6s5ovlTkcyo2gy5R8QP2oc/760/GKUUPAkwLiiFVQHvfvmYhKTeau1mh
778SAMUXWF5SiR0lfZAzoMPrFal9WFUT59wx+XYbkGf6Sas7fGtfJsgBWjyKGcph
GH6MdnIImxr8slRYLSMYI24Xj5q2l8sp8vwRMsuy0GZ7cURG8Vnx45XLOGdMYXY2
KLKawyO+rjg5bY528YSE3liejwZgG7Ln1QIa5c2CL4gBUnU6OuN1ao7gIt+Evdtx
tczOavguKA0Q8zUNZEv2cV2uguR3BIFb3fH0HWSX97wRK+NNMQnuB+e74b5DtoF1
4OqDGUnrAtFCUFFqvIPHthC6IQ2o9PlXJMZWXkFwDZJwWd6e65n0WXfTNQ/r1CbM
o11u6j3hNV6D5XGOCUgnVHmJ1BtVhZ8aGAnKOEmS5PyzZIaPGLEac2z9WXpnzB8x
uycxLaSd5IPFjtVsFFCeSxSmu0ttiIwYsA49q85zw76D4Ky+G7q7J4T2uufLjvYn
tpOztflEIxjisRjA9wnHCxxn4K00UaYB3cas4iOyRWCJ4g7bPmjbcT3CBlx24C2H
bf4o1p8pwv/SHGLB2q0+iao++ep63NlOUCbXLJzZJPzBXUnalemuOzh4TGKs3k7H
rT2QsYD8mY4PdJiwdWQYvHN1Khvdtr9yi9Gh7VFsQG0f1phBO6a/7svDRrOOgCjd
A9KlUefx7idsxbw1j7nY1ZXqsEzsIa+quFOzUc11UhD2YKP0zODq8QbpY4DIgHHv
ns/24dYxBeo9pT6mwAEwWt72WDI482/eqj1hTwUEfIkwLGT54aCzmFNusCl8j/Ea
PqfkJOHBW28bM0soV+Rt3Yg38N4FUy5a5QyEswUt0VmVXDR8qDwMakfCuodDqO/o
qGtEWWb6omRbixxpmc1rQ9mTQ8DQwQtOxrr1kyFt9245rri8LCAY9Y9IXTcO5iQ4
g52OtookuaAlkFyWlFjXGjloUh7yczMdN0uWgXzVhhbAhRuQARVvNxxykr/sLdL0
MSLjyivXI/xLAj/DQ7t+Go/eO6n8HdtXZaWGYUrJQRQtT/gLbuJaqSXdUFOiMm1w
wdBSMCHVDWLiKPYYdENfuSFeq3QVrfR3Fj1tYw3rMOjUkoKN1DdbESPL9BBG3lx+
P/2NX+6F0IurEWSr/5aBR7jg31PCM4GatxFUo5AkwQ5c0g2On0FM8cFDD9n5rbTm
md5oEE3cUhjeIZmoLc99+kTJD3LM+SqRQxMkwaW8UJJED8VAUf/YgT0anjIYg1+s
FU1nr9MDzlnNpm8BwYZGMHBgrKbtnsfYbt4F/8OoQyHuSzvleC6I1EQ7htfF2T/N
7JFuCOcEv7htCuYV6VhC2wT3Tg7fktjgI5LD+t6pqJno9bh0kbl46M3MZjApIArX
ICAeN5G/tjNiXKqp7RVYeDaytgX0lKZAY56m+zrYQWiiZ1j+NoTOIo+6023jp4R8
qGJw43lK/5d/ewb52pNgIEZ3Pie+lKpXwb8wt0W7Qfo1FwY4v6hFmERP/1Cel0PA
p83rDrkl3cHQHsUHNvBJ9JmZ1rKQkw1mhwRlShjX0FdrUAnEV9ssZvzP/hLFp6ro
XNkUgL/aw7juvwiYJRLwbzuqs8aKNtjWra4SRjQOTfMfjj6FjoTEBeWuj2uwPwhN
B7xSfcD2p1SQDNCRiYcUuv4xOlKRmAo+mOCHfxsIdiOPpFxIlgJ287U+NMSmGqHR
cgNDXxGDE2tKepJMcI1JgZUvBcWYChXiH01ABiyQzbnjymTDrpo5YjKFHTm8daYL
CXV1w/RDUMPHjUHKmyLdgSkn7L7K3TGVnRKgFurJ+3aGf28XoErCBWDGvM5CXNV2
s6embvVF0/71OTtSzEUyU8KWLdJzt/h5R/VvagNgMrJAIzHNqhegAfXELqQ8kETP
YaP/MPlaIGXtm9nTQMKpUfn0o7v0W6e3ZbgSf/kjpb4xRvsehQpFWEeONmbkVPJQ
f1a1W0TI8dBtjv08zlOcFfpC3GaYJNmKFx2KWDLhKR7bWetn6kJzHgbV4TmAv51y
VCLrJPKsp0wTBAtSEXHBDaj8/1asJese1jmBCq9KxDCpeavnp4RCNbQ0BoTyKB1K
ujgA4xI1lmlw+iK280x7DPZJGcJdTQ9RZvfi56iwREq2D8rg+TQrpjG4Xa392lZg
K8Fm2huJ2F3CKPba/0REMXPC0XGk/OG8m6V63XZzmLndNX1f2UF3wq7HHiiLDwev
ag+fFbNBoN+YT6u/JmsdGhacOnoVctW+aFmNCqxcln51BpI4+jhtl9osl/6+Tb/2
gndHZdzM7+Lt3LRJ8ENcS16LAODhtqH1bQfs8241HntB2qfiPw6sSlMOwE6f6AC/
csnYenW1K5IC8UXnv2KlHMz6pk8NDviSu0B8khAnO6CNpv7LApgoHNaHjsExfcqm
mWxsuHklUAOqAjyab1ModgadeO8XsNnJddpT31Ia5qZM1PxvcgMAl1hPhCJR47Rr
h2xlRuyRmlyhuE6qPVBp8PNaHrogCUJ3hbD2zVjPs9K2nUwOEq/v1/jXES7q3t2A
Iizkw3WLtKSs0cSZXj3zKqd64STTtFvpHS8zk1q2JftoiA27ongt3dl5W6t2MA5n
mlQg+ilOK8yE3F2AGy5i3tH1d0/Un24LWD5zbyFtb5z9kxJTSVDDedybJ39qG34U
3fpijxyiiDYNKCjJqX3valdr2XuYOSoZofNcHgz6MUnMEeom4RSTHyHdA1GBAg6X
6tH5YKwlinYwsDgOvAtKD/czqT24aKWnPad4WdtfgE/JP+suZTYz3gN6fR7ijfg7
F4XZXDIGr/PE3ZA8QUmqwqsukifERLLWkE5UH01/PzGRuL+V/eAVgcSFiuQAyFAU
0FPT6ZTcwSsX0vyIEv29D6nW5U0DpYxmwgXemlkhN8CyBfiUvuWHw8bkYYvPRPya
lrCB6MMIKx3IALGARNQNOZeV6bHny1m7v5ynDTm8+uOjmimdPL9x/+nViUQdo+X+
j+rcet7SkH2EN3uGNSTUn9gIzRmHqrnbWKc5UMsUd06wEzWT/zn6YJiuWdJXUWcZ
pl8z1W67KDNdCMgX51CbNLLIgRUnY9rchZ7wMbRrDzjUJlULPE3S8HBqOyYoW/cJ
8/UYHxTSntWD5VaomOZILFtjncA3Hb4VhsN94CVwdeW6zhGDpr1tOJWpD9HnV5W8
9HLfEtsuab5xeBcm0WeUSPf5YPr+NOkC2dLTwVY5OqUraZnffFg4bukYhbsG/SQi
41imWR3VPGoTcXTsN+45l5w3Pd6i2JL0U3MQ7MJa/upOjPr36NxzEwBgZjcB5arV
MpZX9ybdIH9ScD0ELYdiSPnLR5JCoFFci7idpSSvMXBNmxaAcA2W6dWvSl0pMURH
8LOCxLWtQ0yb/NX2+hhKOhPOYOtu49NTz7Vdlh6DrpDuK0GJyRgzYz1DRXtiGcxE
toy7uJhMyaCLDfrG6JFe2kzmOvBI/TAjwcHtYguLBnSpUe0OdKbkGgIUjfqagUBs
t7shVaKuxPNX/3mcIRM8ML9XpCw9dhxi829VsiNUizwGFTl2Ia6pxOYX52k/Awt7
nLL4Srpfy5iNL5FhMldObDp8qAmhXsu62CwTG7ZnlZRN0BYMJdliBoRST76C3zT9
oEAPQE+mrwwxyu6FqpKDqmIJG5qD36zKjfI7q+c3WLr5jdmy6Y0biWVL+DnoB9KP
s7U53289pSxvDUKXbxn+Nb/pF+VGCLvNIg31GoW0KAb9kXnci4RlMcQZMJet/nKm
nBjLfb7yqsErRXdI4Q6W60j2tJnJsHMjS13rrcHJsstk8jILgHAEocY/N0kLERgE
mIWOGUAE2jjl0Y1fikEvOrbQ5cAEf9o496OzaAuIe3uY5+DkMdKaweTxfOp7h1cU
j8osJFdLSA9cXo/xYWzWsf1udkS60xsClMzqf/G4Opd3Sq4GUf7sgTmt8SAGOjUl
nvXwEbzl7sDa2zWqXyTy4ILOd60IfbHPheSlULuNS1sPCAXPvee5Iduwdi3WXwvW
07vlW3KTLu3x8HaN/nlZQ1gb7xV3yE8G4r9pSis31zRd2kI1k97ECsdjP4Wl9rrn
5fvVjyojBkNRaprYtPn2NIT3XQglAwd0ItBjpUGPkwu+v/kntYUqhjKpuC6ba2uX
BbVbkRDfgLkcV+WuAMWKZp4nnqqJ5hcy1sM1scv+ISOJFmo1bUVYCI3Xivfmlc+A
+JFk7od2UVSOAdJ2OAZBXXseczRSbG4f7rlaG0vFRsgWrIfdl1D8cLFbyLyp9qmc
tS1t7ABzobe+lVUf4+G405N7rlIjDfBUDjCdfP07XWNYRmgflCVIepFgRtAfirYA
ZIYxSKVU+XdF1UZDDj1YthmxEhnl5FvfsOu0IctIVRbplqGgM5EWhhk25R5Lgt0q
Ymbm2pFVEwepyvEBUCUZkhWl5PyO/EGxJpfP9Dq+qA+UJZ3H13FVVtQqdaHaiQ/e
wYGFvgYpmP74zo93IQN/ouKswT6/zJPmG7Uww84/MxfSerRBlllvR0Jon9G4Hvbg
pgCvm7Y2WyxrCn9QvrVrOQW0h0ZPDmM5chEUUm1I5kvdJsEpk5uCbAepADQpVU7N
e7tjvqEUWkfZMy6ZX9J4ecwf4Uun3kN5bMa7FyqM+Aa4CfgSye29XgXDiHn17uN2
AOTwn+tHOiHKnqNcPpVIx5zJ1dcmiGxc9Z1V88PnStv9yPSrgyWY9JenliIm5Tiv
QcouqPKGJFLXExv5IVHNAjsLdHnG+XeeLI8Qlo3DKpHMzeSEMANbgde6w59gAco9
KAgiysMCVVLuodAtClXm/sy/EWzdUvqw8AlW+yL4c9/FCVxnPjfjPnGeHIg+UiOH
gkH4hsNKTDjqHaz77cgSHblKeDTYpTA7jFc6VcVrANtlA7xeK0yyef1YaDucGypl
D9KPLtcO9spwDB8P1+p36YQbigVG4s32Rtw6EAwQHM/HXPIWFFdtJtK5iTzpTfzH
DQquI2z1Ej1CTp7+Ea0DxySJcGteqbrX/ofuG05F4KC3lNkS/6DsSFFHYicMCH/m
na2devYcoE/VBdhso8XLv4iksLpPBEGjXOuC/6y/5LZqIUViklfpJZcydOceYOPA
t3xBCbekeRgHEXShZM1kmSLY7iNFiMtZzCFO8Y5Ko8HXVdOqG+Gu/gd0B72Rk7ek
sgYUMn/qGuCCGhny6CHE3jRznPNswG5O5m643r+cJBEYaPZ8hANDkCRtiG0QHgZS
VfgQFPNyUHplnSL1DgLmW7dcarD+6TsB1T75XG7ZoS0r0UqTzMHW/O6YWQh8URE2
BIFP41y4A3HtirLqjmtfXF7p/AGz0VA0KBkoPXpQT8P8SpWcFR7RYKBcWOaHslh6
OAsImPee2ilQ61zpKijNJ7hxgdWK2QR/VukTfnG5BLIkctp5blmrNS8iftCy6a+B
jVQ8Yi0hIzN73002inPcmm7eHLIdQTn1eqmOCl7RonIunc3c97YmJAs7HHCfIEKy
i15GJQ9et9R+/CCmEdcguRNB0N8lU3YNskL7NugW0EnXYeibxdaeO80kHnQZCt+l
B1V35hrZZESEzr/NaEsSGtnKFQenqoSm0hHicF6vtyX9x3HA0Ql/EqAGA0ObX26T
uMM+nM/K7yzenSdFnjG1/F/9/iLka878N+1kJCwjQlWxrF9nDLzipW5hU89wbLjk
Kno5LBDxobXzCSZSJXpA7MVq20nefwgcXtz+tt686OQyIfe/MoH8oA5x+OsAre8w
bW3qE20shXWI+DrawddOI8yif9+dlwUx5dd4CkOTyh3mh3ivLYcEwlUsSzYpYcgi
oCyw5PfBNatLISXMLQwRCzysHttZEl1HoqLz+NZWZfqPSikisp2HAq7X9YIcmknx
ahkMfj0zGN/GdJKZoReFeIfoTMprzcY/lrqM1yK/slfKB7t96s8DIb7OKSaymWos
KfHYwZHhCiFav/pIygOfsMtzjKjlAXMI3/n4Kkl5xKfx8F3shF+Gn3M/PtvP3tqw
iFtY3lSGDG/+fj7B3qo7TFTec7VJ1yPZby2xoFBJFguyfEgV0H3q24paEWw4vWft
VgxEUEABYqnm0fndquFx/1dXQQVxzj4/J9lNlPtT4+fE2KeGDk3MOx9aD/vK06OX
tVedRU8JSI8jghxW6Pxs9dSLjU63Hqx2cAcWcsXp0Ll2UNZO5UuWQlCa1oEzChL4
JDFGuQLjW9sctTSBOsZ0/t0X/kmZp/Se8/gFqQsVY/6oQ5Bw5V3V+Wad1rV+oDoC
MJQIEtORwvZQ+JvxxYFN2lNNkM2RR81lesfog35zh7uEjyyXXzizgNW6geuwfT9/
CfoUVw/3Ld8cj4DxEYvuCrvAMebHEFSUbpHM3lzeGiTl+g+wGLf7k0CboogxX3AO
R71ZBvJQMbQW8l6Fhf8f6359Oe6UvVWc5882sLH2kGR5n0DCgR5sqB1UO4gwXmMy
keg7vferu6Sc9H9PtDB7hoAFGx+VGJlvnUeylCvd9DAuLE552asl+H+mmgW7X3/W
ZJmxiqSJ8K2yGF6JQLIDsb/94QW6x6KjKOZwR3a25jdRHmaphNkrNVQVfw4lI7Vc
JJaNTHp79cHOeIU2zM9CKfwGYYnFDwyPnKLMLbyTN6K0sVUwQbQyzq5bt7K/G/bU
F9INgaKfuTQIa+KMemch8CEXDkV/EM6Kq0nF2x+ftAM5+G+rLJqlrwkhMTmgWwv5
dwVd3k3oAtLsTQam0jE4a9HSFlnGlDXbfXMJfCfuIVaB/hcJRngKednAV/BFh4f3
gct0GU9DGDO9xwyrpPBtsibkEL/2w4RYak98dof2hdkgH6TXGFltSPQyHnenFaxY
VW7MiIb4kib88wQn8wduaHljK+Wig/rrZVnPaKYA1de0pcavDGA1OM8kPGlpofmn
YdrrLXgICvNmA0PkGvtSuZmnPi6NYZNyN8Xw/AEDbNgZgVctEtVSck1NkNqrRv3v
BjS03IyQWSWLyS4cr8dWruZs2Q0XFrBmyMxletS0ShsUbRxGXkLnzcVi9c9QwhE5
uwLCSMz/xkt5CN7hs2zYgjtvbuOb8xL8sPmjtoC/VxMDtTi+aG1ARUJnng9tc3Za
eq++SZHgWNQ0Pp27tyx5PLoZ5Hwukf0AnfxEtsEG6Jmrare0RNUFXELANhxa8hL2
DVdxE/8P1zBlS20IorzvKV74AkqoZ2OU39pa8Q6aip9B9JZ86uFFUdFwttHXnVMz
YUgq5jpbyMtJ7+ri45tj6WdeHPKN5vQ6qKpXIENjjQcMkHiCDuCLo0b81kkOC67z
C3hDPmomthO75eCzRmZmQVgDaI4HLGN/vZlfmfDVbOX+WCIOT5/FNF5D7Wy4xynR
dZ2AmIjIHVSQMqp26V8VsFTgcn4U9iLkNXxcjQytXdi2LABbsm3oOdNMd95RIOC3
3q9neaXC0Mj4rIfKm2TS2vUl5ppfi8nLzLNVSWIK4eTSBIMVqTvS7rjORf0SybqI
R6qpiocNblztjD0bWuhH3j0+8xx5VTSrk2NvGHKWNexovln3agNwUu3UmcaSOe1w
alQaPg8DC3IrUYL1bKkDTIhZrgwpMdIJ61FQnOP7GsM2KHiZD9kLcXuEpAzXBX9T
au9/8P/ZxmC/mBevVMPzSmNzE7aMkqdo5+viEUPijurbQN7P4aFxnNGurjk2D2Y2
9kADK7uSY1JR4AD6lmhX2te18OQyaIpmglKiAhByBUlOa/PUI6M82vXbxy13nxiB
uVV3y7sBXKY3tZ8VNf7ziesz9nzKFtUnXmEEDEkWzQZlO72gvl4r1ibZU5MOYx+g
60OmMGTKfxwezZqirSmGd0b8RTJVhnlsx9Se1yK91ZvVfE3n75oKwad541ZUDOuh
OjMZh1WiEh1InDtXqwLX19KUiwLaBdORzndI9g6r7moY9PtsFiSrk43ZbyrwFFs5
LjWIzv63zq5QweGg0NC9BNQDUk1FbuAspLmogRRyaq7KsbfydhUV/R1FKZWGC1aU
ZtI5jnNdUF/LxHXPeGkYXTadO0crp5qOQdTIPjaa9bjJZGeIgbVisiuomhzjJUXt
beUvZJZ0BpKm9+K+9ef81yHMUJmCyLLI7MpjT2KfLDSEAzcj5Af4bJkFOaeSeMGm
3RkDbPoijiaxW/yWtv86JXnytsp+8TLLoommRqR2Gj1Dq/N1AIT/1/AYqSxBdHQ4
u/ICHneFQNKMRFz1NdWqV9coNjY/hWb/tWLhvaDqFhiPkMLquEGln3PfHXWyjBQl
qeX8XgksUbVs7U/KkYJJ3/QMSQSrhDrXzzwZopCiYrnJ7GjVnReFSyk0vjonbtA+
I0jAdeIJSYic6UOS2cPEL09dff+fIsEX2FQWBWQlt1GBjmMAs6owVTQtw/Kt7uD7
htN+gZnZm2i2cIzcU7eBls8TcYxGan1lahhfPPn6exLMvdQ8c+hN3mKMbmJ4vEtA
waLrCZaciPDWjTykWzcNQoX1Hj23vefHoA63rPa4O3okAz9Ot9nw9q+CpqGMnyHt
qlFA4al+1puDDDYu538Y8zApY5JSqOdseB7JLAobDa5uBPuSchltiLjZVHaYLKdv
neXqJKGyRV5FDAo4rym3NAwHsyaNqF2w+jMzgiQOYiqct8fQ7jKzIE3A/xYEtYt1
2joe1JvNtqm9t5BvNXXv6Qfpj4z1VevEtRrKvf/Uek6PdIgnSY63rhAFqMYId9d6
+OV7fBC0vZHTJ/BMWpKpKPUit1YWivLOgx7TIASoIoUwxXnig7iHHVccteuWcZlO
Wu8gMpv2GW7aqzUjZfxckRDoGQVePCMZfWExlngppNXFD+gynx017OrZu2UZq5C1
P4fYj09icyLLhi2cfjIJCAfQyGImoD4QIhzi191ynIBZJ/kVM4bPDl9BPY9gHoxn
6BoeLt2J+DF6sLe5kKdSHzB5LvxHZXb/g8v2ogE1md4ctq77XM6ADsK++Hk+TWyQ
WViLNkpVTIZUgv//iBzHmqrgXIF69AOh3JdMnKzBNbC/qOpLDN7x814twKN/M1JD
4qrv67j2OF3jZrikPOj33OyW7rSJIRfBwPjGgvdf7+eBY+SlcJaklL8yMYH0a7DA
4AgfQITYXWtZbWFI4POJABFwL/CblxXs7RUK32xkWE3vZiw2P3+CBlwTSv61HmJB
h9Nc2WquhFp5QcPTEs9Pd8JHa0u8l8/wKHoztsQIxLgVFdFICs8qYfEE+VxBf0bn
/Tb67pKR38CoFHgqggnMzcmoCBOw0K+D1mOaH8zbXjtjvOA/vbgw8+5oj7Sf8KEK
dJkOBWyOmVzbj0LlUDGIuFYlgu7gVLI5fMRNOAYtTwxFI3ZTrTpYLYjUHGnQJcmP
NHDgFRg8G9JrdmY10Xy0rTGb3ylTGDtyKnyuVp8mBNVu8cMY1g5of6moLvDnc3XO
zgYy/0TGXBxhODFQVa6cT7956rU3fWoBvyaq2tGrpFe8pPsLAJeH4YPpHTtCh8OQ
aKVzk8DVGubZOI1mDr2LQazalyTLt6xl9XKsxVBZ+AVNsJ3rhANR5iyDkDSf8a22
ci9Zli+1kimp3ypwFQPlnJLWo178jl3xLS3yvBfz8UfZXyDaOXVnDly6kqwYjv2W
itbrPLMYzFnNmAuzyJdZqbGUuDZKsiueCHZW+Uym4iUaSD14OaFnqQmK71bsl/D6
vvkWDbPV/EImIWs20n0VS+iytPxr/ocE6Jcpt1ARRUPl+j3Rd/tF43HCJh2W8Ad0
weCXly7RCk85Kesm1DK3Q63WymtNMhc0S4jvimRIjtntpRXmRwQ739WHu5QrOBkB
NGe9jZ2rLHvKm1a8plSdYBM5SwhNeGCg4tI3kN2JEhZjUfMfmyzlVX7UGFfgsQUb
Qgoif67t/KYZEv1F3yeoUXCCUAj1ymh4RCJdRduTAeCzlgee1cRN9pIaKLjSYFLv
r6rxBDzraV+qJf/lu5OGGn/5XfCCuD2D9GUaka/V7dPsJJgNEmsl/PHcep+qujwS
vQ1Hl5TFyoAr7XEwuXzj1ngW1m6SAldCrHZTN2sgJJ/OGuHZf0pv8DD+eb5DqN7+
B1ls+HpMTLQ7m8bn5dJORFFy4dacn7ZlEUax3yltoId/9XzAKkLzccmzb4pA7v0Y
ia49kC89vIYglC/zeBuIIxiil4n21FgvhG5Lfzc22XoAOD/rYpWeotomNVHm4axz
hvy2ee9eTmvzx4jEwUKe9fUdjvY64v/hQhx4IPTpO5yJmfBcGx7YnggSZyoty/AL
Uaf8qOhYXoapCmiPOI9d2vVpwxZlL4DnuJXbzRBn579q7qi0jfITMhKA4I2fmKrg
XplfzfAEvjF0T8gyvFOPj917uFIjcjFj2vOVIa+WenFczTp2jRV45vMCarAUL5Sd
Qn56O3eZkcEoJKkVfe1i2Y4DFwsu01pFVC7EPRVypvFuWVsdCeM6THPkQPjYqRBG
6PoEyDvVkRvvBrqBwpDPeRzs6BvayfChJK2iO+XeLNpjuCjzeGIOooMKfZ51eVRR
9mnV3pEeIz0RA/xRysBYJpXXJYZPPnppXAO3HQWEA/d7lYHQ8wY6hh9i+8EswLpY
KFIoUmD1xo9GhacW+BtdfiQPQPUMmTGVJaolHaFm+1H4UyLKRHo/3n2J6gzKtcMe
dJmVSoSrh3EGyCsYjOKF9Wh+l7vPGjlTwkZBZBPI2j66ofT1CORRGrbj4aiDsun9
co8AL7bs+fweKrHH997aHRoPt87s4qFRSXoEONV8QK/p/pSTsqr4SdoQoydz9y60
/Qpev71q6Wqe867pwWVAB7pDOVgfdQzlivsaQBSuVH5ibn5I0rfUrvnp+zdpte6E
iqziWlzIotxUHKKh40oMUvE7CJMAdazZoymH/EIFFm5fVoLPzuLTLIMFTAEWB+OZ
sftHuP3Z4PzG+am6Ypz+TgsmXa85CjjAi6K8jt9e5KT2VyDQDfrVim4gRhnBmQGf
XeYCCMCzMZloSzmQIDNjjXl59cVlneBgw2OftTR2rz8bbQehQUQVhggyi+brZHkR
TfUqepa+bXRdPGT3DR+6Q/saRb3bbJJimUuiGl+Sb/2oSPEKL2ep1H758bAJW7WH
2EwZdzemUA6X8dveKpt6AYdlX/sMxGucMSa7lcmXNoPSR5nwo8aovB9O/jWEku5r
ACgpZ/9w4aTEe1ib7Qz3u7Ab6FYCSVoPhhY9NOziLbKAk18UUD4r+eWsqoTAmJQl
2a0pxJPVU7rK7O7KwOhFbQw1gVtxDiTUbfndW2zUSh5sqw3keV1iyakzuA9U55MG
sEX6GJypvHoku61k/ROIPIcmgRvqr3ILUKty37ArZlAvhwk4gJUxCwxdRO8WaBiC
tg+/7jRe+5R+bUaHFTsC7rUYNYFp3ehWEt8BRy5bCcjtu2qT3owypMmYatkKoaLq
n3Pe1JAn8ze5fOFwxwSpJICkdQE9a+HLDBgL1SyYRg+CPCDFgzu1Fz1/O2ohBbJ2
EA0fedCrjKoXsKNNEhNsHXXXHSURJsHVdA98/mMbX11O6tSrQpNsg0LrKYO56uHj
1XEK2evb1QbN/xd+cHSnysVeirwelfurVupGR3s7g9bYY8LfUm9y3apXq0tRF0CS
Vxmzk6r2guZ05rUxkEE6YQ8edbsIC6rOPnvG3FNJsZvD8pEtHUzGc0x8nHKT5wFQ
Q0HjgAkGOmUAlEQK8Q85sNrLye2nMLAit2jf4WkFS4zu186jsSAVDG7c7LSOvXDg
CEZfc03lgsRf/YrZvUxHxtWSKSPXh2sLRGXUicgFjmO0tvoEpZSfzkuBWtlTjIn7
Z3DI28K3cqA6XBA7+G0QyUybbGnpsPnGx2/XZMDvE8aJzp/+fEKcRorUdzhdIM70
2X5YQPKuxTj9V4fp5paiFROslGJnTF1NkFdQE7ULnu+aa6KLn4jMP5OA006F6wfB
S+wZTUnV5b0Es9GQTIqglA8vuTeFzcMYYHXFWX/Ame5njfNboZB9tmk26C5tyqns
6He6H9b12Z3aKRWGcxMDa+UtJZQu9HkrNFowW+P7OlN6MHpNlaXAPpII6sKbNYwq
8JmPZa3uJ4S9MngGEboTUUoUXLB2mzrN679kQ4FdsrQm9TAnkrkhzONslHRp3EPR
q6YwSkgr79ZXpjXhVDpKG/K32WYfl85st40TEmkRKz56GHKAiKQHqTOcEu4hHFdL
yF3RHImYEuk13bwyxSnVh+OTtcQTyR30cVYIzHILdMXyJ+3KRnbRnpte1AE4R1qZ
TFvCQXd6PqXZofZ0OAT56Xe+1qfQONw71gJ1ciY6a982yp7vwMcQIRgd192v8VEe
6GwsDWrMuSDHqpdF9qfTzbFATBhQTZqMBnKKgifaMs9TnV6IKqLXNENmLVruzH7i
zdIyGH/w3iFIYTI0/Qns0C5CN5Ai7pjUCbJN1UvDZti4NmLJjlxY/FPdoZTdD14j
t1PE1cEuXidff6oWwR/uzeAsCSH6pClJYpZwau0k0TMoCF9ycq0Iq1aT5kFxZ1y9
DXpmluFPtbIH5ksVHhhXjMPy/ooVf6bgl8PHX3dAjG0rKskaBZn3VCopGFnShLjK
dGDXFUwe2kUM4D6HnTxQF/6846SsP9PHrfAbg8yDum4qXD940JBfBN86ECItHJdX
sHgB2C1ozLzJJp2q5cUp7oEVnW+qOxMsPl7W76VkSOvwxTmdfRvzHwmZQOs0/zL4
OJFGaGmHE48E3XnLHYr8XPb+Em8I4XbU8NAqNtVeWkLmkA5ktnUOt9jVZAm/FBmn
nBQ3VEcFuSl/WqcvhDmQQ3h/ZysTjWOFAITtGpibBAMtCXzMOJkeU4xhGc2UVLlZ
jmB3hueoL8dI3yIr91ZYflUPVgF2IbLDPCk5lm1id1rF7QWwyW5oqtabGy2WZ7x3
l2n3X7bK0LoiPmoiOwfJYDEeFlbIDQ4X7clCj8DSqtoshn8FppsfkERNyWYBwp1T
c0JBeciA5uF01KPxhtN2XH/TNi1jeimfw3HrOKXtNibJWkvT5VzY4mqhqxU4GR/C
zWLCA+wBFyTv+oxnRLBBkBqjoENh+X0UcJLeT5G4vXLcFWKNtAW5Kxqg3vAHMHZ4
jA1LoOJsOmdph6ddeJ75+cEvoPjgSOE6n3KWjEhaPmpt+U9XKQ7Y/etS1hQaAV9z
nIdof9H/uzkhYlIpz0Cs5HH25gOl+wodujimsNxjaoAtG55FvMjLl7nHiMJoikPf
K+ttnt/JBD+njjK8uEjyYGiDsG+FNrm5pDnH9lbQAu+gHzczGCvhmRdTBoRww4sF
PsNN7BbKFf35foCr1ezT2UFS2BtYZn5peUvs2v1MXpNktpPszGDUi3NXFnU1CcKw
om+Q8KiVO7NHikCd2LjlmkMqD63ULsGqPgE0+Znp0eLJpJrR7gB14w+Eu8sfTNP8
3go1wKDp5a+usr8CT8AINjgqXOlRei9g1AsOMuLicVv2TAGLNv0QagyVW78easF6
G1G4rDAiOaMtTLkJKPaiP+s3aXoziQKEJeJCMsV+UmpFgC+0VBJ09jtpidR3qnYb
EIx7+L7hhPW+xjwgSZuzZMW4SgCcNpJxwc8HyHZcRy7BZ6Ra5ph4gtguZGVZ8S3G
tXZQdr68kfoa5qeMJiawwJkIl134IYn3CBwkoXLImvZcXFDOeIYsl81HUuxZ8Q01
FpI47kImNgKlkNQK57GptuzBHHC/TDl+Oaxa1hbzAUPREOmSUxWJW0HVcqHfLjgI
pZkEmUS/VAwGUzd3vZHCgXAvDvm3UCQ4nM+ycx+gr64PAeVpmvjyLFZoy7ag9eN9
kTnLUDqfHQ4eKTXIFT/1emQBtdUIL5bmTXcbVQwOfn8o+28RrVfWZRPy9s+NBOWQ
3DQzVws4kjNpt4ANvIpl41/5meyt/qFqZRpeXhfx7rYE3pBczS0cD4PViHf1XRPX
hgjuRMvbT7WsFkRkLV2fI//uLNqa8OK5PRFkCWBA02BUSbWM+Fw9HYhJh5wuz9AJ
KfKEXWEAwmzfOSGSDyRonLwvSSnu94BA7L/Jv68seEGuX+1Z7V/5aENJDkYCufHE
u8ZZknnXrJUoUIvyckbVG1UR9KYSnWD2KL1wTpBvBpfSUzkfPNT7h64XnSzpDmvH
uBABwD3I5mfk+VYMXFc8BcWDUJR81s3m6/Cdq298x7/AlB4YCbwEOG70LjhtVShN
YJ4LWmjRjy7yZAgl8OhrFqpgAeVUb7fKgOLYhz0LV1Ruwf97lNQPlJJGQjX1Abns
RacRpA5prQkkzs+bJHh6PTL9uGbkvUyNh35fh45G2iwluhpvIe1vrwA10VDI7M/c
AJeZfX+sskObypTqI68h9MpQZpVxtMQl8sD8+DtTIcO0nliLtt2eUVfi7T5kwt42
f4BRVZJeA1APOkOB+iXyc7DBPE5FsAgV9PUR29bF1kh/3A+eU2uT/0W2IMQdPxrW
1Kifw+PLC/HvjDtUnmS5H1NM+ELFwpq2/gxfjpuUvaf/IMw5kT/X0kP9RzEZGNKP
X2Itarvd2+iCwmwohemujiJ3sCe5gdDQDP5mk5eMhNuwEK/qY6Te6qtnySKG1pRL
q6ilgP95qdNjnRseJGCSdnEsTpIVo7kS4v3W3oCL9F1dMOwTuU64DTbemhN32Axr
V30VaM87jU8Lw1Ry4rOrhJiMRSSJfDDY1c0xttjs0fm2AjAWYv4QEZybm6EcyRq7
19ARlG7P7dF3rFHLQpEyNHhshQ3mTW5fLOGRX0F0NdiTzuJjeF8i1sAND9NEi+cY
A+ONQlcn6fXreyBvqT+IDJH/fgOTrwC+QCKQJJthkTpo1umbIBg+3TUwUENf0OTT
2Ck2RHL6fpRyo8BcTtQ31w9ZoJZiZrYrwZfJrIeC8nL229Hpt5TvacmK4XphOkFv
l73ooi1VaY1pLzljs+pAjkvTj6B1tGrU78GsSSJE5x25V3GEOA+MBqXYAVU2hwr5
9oEcdWFcQ0jpzklgEsnLjHbQrvA7lqHBUNn4APeVFCZiqHEr0T9T4OAmwv4RqMeY
hCocuJ1UmfMrJVskZvQS1ZtFXSfVq9MfWmS3O3v7XX7sRZ0v+eOHaTWe9Q8nln3N
sAIPuVPP6L2LjFOo6ln1GCTPzyoJ/Jmk6hM+6+CSGx8cHJ8pJPlWK2shpDdA7QzY
LciRMsEGUajI09N72SmLiDZXhAd78s23/61IQKacd9XkEln8hRljfcdnbRNHn0/g
t44iKp3zn+sSRuTlQsrwRvLvyYZ96h5KdquGyd5AFVw/XTa+aevN2l3RB2FDsOvU
tPKcxk2ikPHjyUPE6dRItW8YocC93JmNyKu45uhrgxFySXZIPib2VYUJ20BWaRYQ
fLZhl1i2gvF2f7BFTkfFoNlY3m1uijo3l/Ronj1qRYPDNJJbgD7vx415Vw6xSkTK
6IEhI1WM3W1Qva8kATKF4lrgLwr7BLtmsuXCvl7mkbJ/OOlmUcYJcqJUSuiNFr9I
NVIOUyb/nm2z35ZMQ9BSLUVKWiFDjeQ+0UR4R4TfMFL8pJEnvcNXa3mV5+U+6wD4
RuYNiUYbbSpksGEpgaekrM7nPIHXdegQ5slNbANimruhj1zi73v714H/h1Mgx9Ao
ZmGHCW8kUHa0SEeJ+SmGknT94nThm0jVx56B6oP1Gv1gXPd6yhJ5/L4UlxxcFV6w
1cJyhW5dWYZIG+xcla0WoUmlVThFLLrANEr3AOicC13nWJDluiehF18hQmE1PyIe
BN4VpToRdiSh/HaGXwiruqO3X63SYzjZQVqYRFhV37iJnwJ5KChORceiuGEn1nr3
vHdk0dAvd61CzKeQ09sWRu4lO8d1p2uQOm6TB50vZlNNuD/TnWDufvg5VJtV47dA
GTOUHyyVzfJtKyFvlYgmDw==
`protect END_PROTECTED
