`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G2V5fZvCIprWI8ZiqagrU2MNkDvsIeEzlIOOXMcLi/WvHF5dPseHaj3XX3lD4q2Q
kvaPH7X8sa0MqznUiFuU1wDPlxUF4HDI95jvap0noGCooxE2F8ZoHwxDvnvtM646
JawpzRIy5/Yk811iSP851muvTO23sZxco+OuJ0s5jyLrSbvj8SG47VVVwo/UHMHv
eTKr94dJqmZts0xnPHVly9Sm3S1nL1bhHVK0hl5lAl9ABkWuCp5aCyqT6eaLh+Lu
O3FYG1Ov+Edb8fY9LYqg+TVS4iipKuuisIRcsJIFdF6xYpXHfGjZcCQwzBhZTgwZ
7f/wwUdaIdG2BKvfthquZllOJa59mhja0EvlkcwdDo0bnH77M5PZsDTwkcxdSYxh
tNyRfkkmvyI9xIy8n22PaIC3s8MnTQWqS4P/9QObQvWrwviZFPLjelzxAx2RRbQJ
p4yxmXfUfyymKzXvYDpEEbkgvZRaya+KfWZLsjB1lpXU7BGcTiOaKunGmZUht8xw
l8rxtciZmtFmMf5prkU7+1OC1MLZJOeBkvxYy8WCYq1jXQc1RYm0uzaPR7hDmHfq
Zq6HUxCigVZ0ytvIkTMDUPeF7IEXpc0Jc0x9xLbqtDw/SNZm1v8+FI1wmZTuJvw/
a8rlGIOf35bgmbRX7YLsVgnTQMAyhrC3pIIHhKucuBIlh2tQcWBdhrtQpS4txmm7
l3caWmJu4VTdGe18LafrsWmeM+hnHfbtHPpH1SHVetfy7ygo1WfDwoVHceRFpCmV
xGU4okwuebYAh16oeMNQHV801IQNFoeNWus6lkT7z4tHjovpua8MdqybYEEsElCn
scWSIUUuyE8ncI4z9YTDmilRaPtbDjv3Dells7aPq9w8MDhhSqVvCTm4MVKWNGl3
65CMIW6U1OCRfVGBiezE6EJycFUueCbqlg5Rx1SJI8qdjVcei+PUzq5iMt2VxAHs
QOF344pcAskeCuubtwW0yjzBFKrUVdhYmnCBBil0qC8ri1TFz71BuOoiPr7zmJQu
DsGqpBxKbgRepTumwF9OAqikZ8Werhv+7Y5zMCLjSiStoY/kvewy8WfOfAS/ZEhc
WwsDCL5pHVGAAgZdpspQQxZ6IYOIKDeNHHAsybewOEYt2ifTUbdG8eO8ZLaEpAiT
EC95n6ypBlCCbu/4FGaHbfi4LKZSWEl98E8bpCwNXzC0p/TfWCOCBTMnT/kgLuuP
rfM7W0KslSOQX8pfocl49ZyxyvdqUD7KMYcrX81OWBI6HAOS/tHM/3s//qCKOAro
eZW9qKy1o2b0qe7QklJHWROs9f4TAe/uiHPZZF75H1FyAMX8v0UTKezosW2vylou
6317T8Fww5Sb91zfDWad5DuNX+ldRAt8pfpK4kKzeQNcsXH4vKM2LdTcdjUOVYra
1mAAj5k3oJyj1iICc2QyjAC48VPhzG2mI8ep7S2bfNcaCpG9KJ+1SpMnmGXnghG3
kOiiQh3zH7XWR1hw/ml9Smg4bxMB2ohx7UZfXUYP6NMhOCenxlQd0jmr91/eIXbv
wuTj+0e4IP23M4BITvDEbkCiGVSZUGzt5pFyYaPT3dRF4vkoF0P9EA+svzfbP5pl
D6l7fncknnIA8tYBp2+CSAVqcKV1GtLib8HpnD0yI5AgN06nvfa+uhAgKRJHPxus
Xk4JpTLBXfNzfHl1KRTPhoHgFXiPhb+Uh/o0Q2dBy0qV/Ip79r9K+FgN6d6SUPGH
hLtr4y3X+HvaHG2BIwZQpt7ayyNz1YP9e8V4UTNYJmPQTpFnwLwx2Qp5Tl4Aq7rD
H5YDmmKs+2ySfBEuUlS+tO7JpsD3KgqVDeIR5ny7n/y44PqzY2PN91QxGkQnqW/c
tgMQRP3vKp96atJ6MwygDWVu9st5Rey12QPeiF5hZciUZb6TJltBub1lkdVTo2Iq
2ot3+54vaA+jbx1j8WlGEar4v1SkRoubXKvZxq4hiLwYJ9FHgSI2qVehYnVIV9HR
33Lc3WphP+kbeQi2g2vUrtts2ZJzEN3eforAfXRg5yN1cCrL1N11SlpvZ9JuCmJl
xubhVcbBj+wRXsXDfsK8zI615zyilImiEwWD0fLHCvBncbCilQJR6B36GvYNovA/
hAZq9/wApBOWoLzdMt5NuA==
`protect END_PROTECTED
