`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F7HgkfkJ1eNuhXt3PD61qETeuRQn7GD+Ny3hptTLcq6r2xgaMHUSNpIoiWO/c+qb
TbWGj3gYrg8oKzsZu4JNlJqLGcu5cV6Wvv35QVDMaEpaBWUGlCRAKTSuqOSCTyUs
59/8igIId8URl50wXX+mR5vpFZ9NT7P7Bvc6WHFwZGuhCWPXBC2MayN1JASNPrM3
pxIUf3CrseP3mq2pUWgmZ+Y1M+2UOH8RTqpk7dbM2aDgVQAWIV+f0dE7EbEE51AZ
Vo3mnueHxowxH7OdjOvtS8po5fq6tVxESwtCyQ2EQC65O8pU/69DtwCIo448NwBw
QVH6w/59E9AKfGAvdvz0bbcepneGc9m3fRAopspybhBAYAPr84TvgAMNQgCMiIM6
`protect END_PROTECTED
