`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C9qHideYPlrTTyyDIwlEEmSMCI/pzl9LDIsHJ9wHO92sqrpJQtMwH0W7zwWMdVkW
3x/lxBwJPk27X/lvmKck6op2A4/a2wGrWFAOedthjkuhATlz6zQp9SdPLPxQw6iw
QK2SUbAeSaoh8+xnE0h7OlPDgSUyiPsKnwJTYYcoQcZZ/rv2KfwC/M5Ma5iE96eb
yh/cs2eNAJCE+SHGP3grXalbnTer4WzJyR8qHnWsZVe/rlQOEVQt+k0DSS92FrRS
IfF2t9L8yoOXvR9DqYl13p9SOWcwaotyzjpGRYq0vsFsubTT+wxTSy6ByDunqdbm
Ygy7EgLsJjG0s+wXGfwlcw==
`protect END_PROTECTED
