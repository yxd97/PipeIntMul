`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AKlQGo76FKJVqX/9zvDmGqh8HZmZArYlfFUMMz/VKEmllb0I1LZEHkWEYJOfADK5
1bQYxbVQjOPjH6JENJsyl6aPbGfWFVwlVAijFLA8Vr8tlyPg0N0iu69bWSvSwBhU
UwkOf9fDU6744ek+96BBhyjo5GBzoHAXrbubeU0HDe5IE/xleXwVY1DSYVOOI3HS
4v7QbCoFSHMabD7mKolzFQVeVgjdUdiwBZJEJ9izIBNNv2mhlGSIa6qUwm/SmUQH
YFpMmNAx4qRxsZXv9QyenE58cVfZTg9ufa6gJKIAjs4Phpb1ijZ4dc9xIps1ow7C
c9DN8NUO9GMuCxbB2lPLqQcZkUaQYSY0I0zOqrEsoCuhkuGABDKdWpYh8mZXvFf+
0w5qPz7/pmGR9tC2EgWQoeha+N8kk4lh+U//JXhvqVQ8Rr8zAP8Vh7bs2OdTQx6J
UAzyVu9NRZwq54YM4FLdwXe04xr/Qm5kdjLDjUkv51t93ykIVk33qExoBdPJP08X
cr3uazh2vkGyA8396x3QgTpkw4SY0R0+7OdRgouuJ+c=
`protect END_PROTECTED
