`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NvovwDE2MOcJbV1vbDJYrYzfWt5I1d+1B8GTesY9/D8tOoLlDTW/Jz9zWbeYRrB3
GU79sH2BrWrlqWKY+vfEDhiJtafuTrhqHVbBY0blgeuTY8cZIIVbXFY9oO/+qaFG
g7nYIsI31Lx4O3l+OzkDhnBdzO0d+dINhLCwyTQlcKZFmYDzLX/I477E5QgthglB
1cvWZyaOyvZlRNYlGpLMhOwbfLZ6eA4dU2BHf+ywSV+qJnm2sddA3+PlZBHKcp2p
YuVCWC8f1C7WfQtNVZVM2Tqk77OWB4UECmR1ASmQmM0XkBralednHpVFhJcWXg5/
hdW6mTyNqmUZKq9Z5Au64NNz3rvkQNA7XgUXT9oyzDVvavIloaah6fGp4IFUB2RT
NFMZRB7LWSaoIupCgKc132DUzaIWbWF7ewSCWQFdvju/hwY1m9RQmntGHtQemVpf
V3aHUPPQ1YA57XkgTmaEPQKfCxZmSiZBDCqiq+wRU2ppdjhDy5PTlKlhXZeZu+2D
pIAbJYJnBRIfi2NVXaWSVTV0EGbysmR0E8xpUD0EET68/+tTBK8+bv2GLVCOqObr
kbZKxdmARhHXl7MYwk6IGg==
`protect END_PROTECTED
