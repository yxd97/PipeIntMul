`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjm4J015QPJTqVZI71TqlR4pA+7WEMsSo1eV2gvHiJGCkXLg4yGEw4k1LSRtshVM
bZs1QRKAFp+hUVacUUTVYZKQVJcUu7SIjOqkd2X9Mu1WlFmgiNXLV5ipJMU68SLl
iq3Zm4D+Yn2HG343vluuBvdA86jiuoDaizsYtjFs6EVDyOD7w2R0Pdt88dVfGK0f
HvxRcSQU1XWAdgNWRyYGTuKQnBfU5O/Fo9tged7zWrC/SxKLEhm97zKUHMQSzZIj
ZAsXhnu3spjMOxx9JUdOC5RQTA3fbmd7tVm186aP745WJ4RAZAatquwLuUCxktnS
`protect END_PROTECTED
