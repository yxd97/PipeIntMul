`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mma5A+49rIVZIGGFO4dmlPytvwoftUH5l+3T9yijgf6IEJZ4YvTl7rbrGczHPnzS
DviXfNDn1H4Ixw6R5nlKL2EEsgxn+eLE4LZVnXCnWlnKxiWEte68fYSEa5ZVFIUp
XMrGI7AFw1i2Ez4IO58equcjZ3IyITxLhDCD3p1RM04r2AZIjKxl6s6+eNIHfZfm
U1ES3lJu1sIjR7BpVOT4PmLvZyAqvSzFAuq3StESTH8sPgZN/kYW8ZpDNB7vGKqS
Z1CVz4H3o0edTeqr4pm7u4B/KtUwNFb2rY/z/UJ5HLH7lIXjTMjwgaMbPvPinJpV
9rT6riJMX3XLwTuAjxPbSjjRWmoGZYMKkgHNaSEBR22DFgaJU1dSIhVvmGAVbbcE
OrooUFUXVb1eS2EaNWjorHYAORsKckI/cOn81WTvAk1kicOSuHUO0hdDKQCONaa7
HPe/Lrb88K8jW1K2wrwdjcbEPLjmDDVbuzMnShjRB87RmQ+AUbkSkVTIcKR5y1FE
XAn8dW9Bt2TMthyMVoOIJHcW6CeR6rLJjZifz6/MMiAY+gcegWzuEuYi044o1Bf2
BpuK5sXKZZQJSEJUZwLHZQO2f3g6yADEVmiC4VOdCRLbjhL0gqWhjUt4EtW1DnMC
ngVRZc+xYb3VpC2UV6Ee1Mtlq68MXcvMDr9vJii4qGlrSkuyGW+tT/WfEGNRHJjq
K0nSRiHSlZHUK2jDLCAYLOU2QT9qagtBiQGywJtyBLJ/Ler9mnUhsi8IXQ0TYedw
1X9ekfuZE8ymPO6ZlBcsfg==
`protect END_PROTECTED
