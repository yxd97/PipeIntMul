`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fHYgRyzaeQCkhyA3Hs6CZHhe4IcEBPCS05Mc+LdhHbKUJvX4Te9u1KCaNofGOQH
PIoGT+CegbwlUO1U3MxrOKEZwdyKwTVx/r35Eq+8W8Smd3I8BvNtpJchLPH8zZg3
IoifAOF2fuVf3OualKBKv3VIaH3mqI66bgGRl3TVqFFdiMEIMKS3Ie2vk1Zevg10
z88mktuiU+DeUPxlr1CPl6pX2zGQI8+9euti+LkWw9mEXpExJVZuwyh5kg44Fefx
N1pd/23KBHdKxFm9I3Kzt3sjV8CQIsKMJkP1In0Xhs/YLOwE/SD+9qJ3WYKNLmSb
kbU73RemDhTGyRruhEKBlVGV2alAspcVzQk6tv7o0xnTRwUt7mDELyfHmJw+ROdq
tn4xSfKr8I/YG7OfpMcrIIEnxVuQyJu3y3JbpnsTag0AHsSaZal9D0zZ9sbuKALr
WFgloG/q/XZlthm+9n/Q3tvCZKB6MHQn68bJJZJsrzHjYw3e+0LfW915vJPQnvO2
42hNjQEi9oPyQDH2Ug1/cLUvgDg5YQPLZuHBPrRrEFp5gtfZFGCHhZh6sb+9oMq3
pGgoaZkzkaMp0ejDUIllMbLEYe2QIhp1EA3796kFgpbw7EWJNnJ9QIIB80w8OCPt
Uh5Nmy2z0eF2oWqdp3IhJAEGMv50DMFJOaqu3P7X9XbbniTwyjFNUq7b+7WuTIne
KMeurNZITNeGKqEzInboy6jECGvT975UpLt3SlEWQPOCMSnyng6FBMD10j6/klN7
ihR6ciX7mvvH1Mxpp8P13+LBqEehjnnC+Qt1HUe+VK6KNanfMw/ew7qSCZSq7L5y
jcRfJ/Ct6FLtGAqAONFpHLNSeiOgnUelwLoBu1/FEFK3VL0yFTnskLXmaQVG3yA1
WNFBCMUG/ubrDzAVya9fznJRV6/LFqPLwu/B37jCMgz5RvJMRaeJk+cljYDg5O9q
KkOumnciKeWjSmBzwDhHlj0MwnZWxMU4aAIrgE4XOgVIHVqDzy2VJ/jbgPZiLwQ6
gF3l6J0qYiCWPIXwkZ1mcyOGwr0TnrAvRucfnL7armgKONMlPndFrvyVVlpfVsq8
92bAUDXcLeBcdnUQeErOVMRlc6GtcjHtrGpk7uVmbrP/WRld/eDz1WyI5hm1/BAG
3npSTjWwUfxuOBLnNa8MIAn6LjlxH34LrHwbw18CzriTO+8nuvhmMJ6noJpzQRK/
WHbFlrnYr+ieiHZ7KW3MiGNZgIfQ+hv0VyF2qyJZDjU7qmyMx6U2XzYq+D0rFIwx
DW/+nCK6FKF1G03JJl8Po2sU9YrLYpX01IpZmiudkk9B5u8EUhEKa/Vu4WdafvtI
oFeJkos+bFq/BNXYU2cyvoSBNyb5F+W6BnYOhN9JvIDZn/suoLYXvlGM7mGBkF3S
N8wJ5SRJFz8zVzUuow4q6mOZEpDR9hDM6uGkkWrPl6acua7k/N7iITaTlJXyPLvw
Mb93pnL5RpRZ62hdczzExIzsPHafWJgGPmIkcQ8OoQahvGhcwf6BMl4SAUxihPqN
9koJi7NlDNNRPPeZ6l1/7u6AdmLsRdKpdanvNXV4XDDO2+0Z0hzEwByQcmpKFKK+
nvEUQEUCscMNbcnNBmyq/8FRY01ir+DnQBSBUZEyHOBvtrwWxKTFZa1EqFILIr64
ddE6Xoxau4yAK4bAWyjnOsfTjdKce0+DYqpKtmJvsfpeYa8oDJVgJcn+4g8U3mGf
xi6odNL1PycM5Q3o8ksvHIdA2fpzofkopG7Pi4D9JK2x1miejgNcRSlacMAuJ1qf
TdXm3ldMi8Ewkvhvf2r8n0cr4NSG7i+FCFpiH6nDCR8HIRHahY1YWmZEazmT4xC6
KXEyEMG4sTCT9LtSxyFyp3ACzUcGMFMqahPZfMz214prRCkFGn2usrEzuDS7hO4q
SjGuoGmTloDCnk4CSDE/WZBnJNX4AinFq/5dfngYdpBrsqJzBCZ5lYIGfobzECri
A6nSWXo4Szh53EaFPiwFloEmaFEeuQ1exrz3Z48EZ2OuaXKy9Wd50sH2pjW9pBKH
iYb8BNy3N3gjA0NPchAn767fOmk5zcMsILJZ4uz2XelczjUyKPx3v0VgKAw8rjTy
xmKm6gRaXJsnsra2xtRCt+/AZaXUSWEWMIj/ADR77fg8Ed1zVLV/DMGsboAZUfyv
ZxyiEWRLjLi5Xj3ZUl16q6/61jvW6ioV0FFlrqyPxH1Sq1AyatGLPeGN5AE1k+7s
0GyJnb+K+wcHCKHVSzUJ6JFEPC2jv6i1NnYAL3tnRY3nGbnFOZ4ECaGX7U//ySCi
NwGierPAJJqGg+qIXYGAEbkz9+BmhYH0wrtO2pOmpFi9zYhfYIzMkRFIACb4J0gr
GHPj/Hdu2PLlEPUqv8maz3Irfoo5HqFH9NGWhPAsBqBgNSEacioZBc5qP/MESQvB
Mi6eXISDvE/XqHttOAt0xpoTGlpOhof2pnu5+mRwB/PUmANpPifPfqihyuZqZGLo
iNXGfJvvbJclIbwysQL23y6QPEoO4qsB49rbYXU3wHb+lp/5fCOVdOGeItHtI1ez
GKowgFfyO+ARSZwP+YxxUey1AX+zWOlKUs0oaTaR6C0aGfuHEf0EGPT25FNnD2H8
WfXaSr9rhpz8xtKVqeufU/HNaarTt8ofRLE60Ewbjwt2coI0QvKxO4QwvAUZp2qU
qdgZ/RBrQ/+R0QDx1vBi0UqKja6oGa1EZOLic87XjnSinjwCLm9F9aRV81q+d9+A
RHtzFuv9xlE0oai5B7LwHYwOTpYUdRZ2Yjo2ieSKjd8zh1O35IS2RopDUy/ymgBD
Oi7m4lX/65BV6gqZrf85Zr95fwKAqqcWVmY+qznjbhBr5RETOec57V08fRqIHNh+
JmFjxdBIGMAIpQdo4rzorqFpZ57ic1KDpH3cPlYc7gRUinwt7+87i0el6r1qpsbn
s+Ifb3JNVSfZWa6+SQJYe1HF/AtM9H31hNNHSGT4hZNamtiReaYr5w7zR9cPFo0A
8aW+XOQTRaRfqeO0pVZA3GZTH2lKGKqJllSq5fZotJLZVjFULPOGsOoSq/qjl1+c
MmnLk7YmLIzcuxZ7Wzr/RAYyB1+z5SDu1zmaATdY4B0A2f/sQOymCj7WtJsi7QCt
GXqXOGplc6foDioX+X9irOJWCGQrUUfs1483B13XErZGHlhnVlrWUwchZN2jN8w2
UMBCcQ1pOoL/V+D6PwGaxz9VtEYJ4TweBXK0T6IuY97Wr98/6afQYzK498Yh4CID
b7SWvb92Rb9WVimtW+GETA+yvnLpa4AhJdBmSiI6onnuDyArE2ZLKnx31Xhvgo11
46AM89fiLrWm3tn0Ua5Rs6EGh9qcqQ8pLBcwt5i8sr4NSnbCsE9H1cI5bI88Q5xD
UaLgP3djnMyeh3JKvPsz9bB4sMgqcqVQ3vh1vUQ+mz+5Z1xP6OWkUtOyK6e/gdMn
oZMs+J6AB2L0UOpNAtk4vSnp0C2/n4jzFp7iieAG55I7i3gyFrcd+zaDowhGflDK
nL8dCbTLsJJnW8Q+y5ujziL5B7S8LP/y8jzPGYQ1VF4ELqJhzcFj6/6M0h/HKZxS
1EzaJuiogIWuTrcimTnWfHMqmTvcnq5LvVKtrmlAc5bw09m5+gotQWZ2owscQkAd
Pc3QGLL3maC/QMq8U5VYU/hFiAMWtUojfhlTUS1+f+vGi60rCI8OXt6s3FISP/16
Hia+NhEdN8DF6DMBohRAjcs9/YrcIm7iMSXkiQcEALsO2oiqiI1vnZnO5KtQj316
zaE97bMb7qTdxP6MxRvoYJ8jexZVaLykuErviHY8bsrgZL0Ix4UoewSsjGMgRLdU
GvwIM8ON/sIPbhA5vUREpRs1x8HoeTRzOENWOjltmBU2k+d4pQoc9f+zBNH2J3bf
q0qliDDTr3OXK7G3stwWWuDo0vy33PqRKfhAJ7Rr+4gyNfQc1+xJaAGCSnrDz5MO
MblxS2RuH4Ao02iHZ5Ilk5qxsqWqGRvwLP9bbPRu5mMvgteI3FIj3w7Ry+EDnLhz
gv2kku1TUdVWicImAQPOKHXbIVnPPBy+idPE2Wr+AbiIwhuOAj7JCDBR/9ToT4Fr
uygdhawDVbqzUJuo2J16US2+cKsUMRuy+GnHva9O07jhdFWLidVVnnMuNbRkasVJ
vf0PUX8IIgT4UvmDRpLRqyUK8P7xKQakBC08zs3esGhmDbt0oqp/ZzHZ2oq6ktwb
BUoq6VcRRE+94UlhYobgtrtSW+yHFfMf6s3eIlM4GbicRxJIFpn4pybK7Scrn5SY
9kUzWQtyit20PMOoSk9mNFV6GBqm2xWZiFRFPGI+H+Mf8/Vz6m4PJgtiON2KXyrD
79xn3TJhJrsv6E+uvdNqqO7VFij+0VJuUsa24el0xpMNhN6xKJI5Q1Roq0NNRue9
UxibeIBujp52adqdvLfTvJmRUyaYfPSJTraokXT1e5AZ0ltjbudht733n9mp9w/U
84RIVa5LpwWx1zbyH8GaEOPn95oCYSB1Vy1zKa/iRIES9Xo1/ffJ8iwegRkA7g7S
VCvl0+xzPMWEMrHV/UoIAKnEF3mCoi3lTeRUpD9SeXODl5hlH6/iBqGEiWIyQL9q
9ux2lHkWNX2Unc7uOrxVQEdood0PG3gRtGka2EKA4tpqNZUWPBs0gPymfjV+F5Na
jjU5GiQ3hWzBBx664Znnkt5Fs+2szv7dm02tM4MadUkI8REZoVsb6jxHHCPBoTsZ
1JO0ayZCD7mETBZqFBJGvATM7wt/PTanpMwtrYOx4dnw0Skli3yG9+ZaM6wKoVyd
WjYV7s19I2Gx/JLwDY9RZ+Cch+j/xNVw5SN5+HgCele1KOYrBO3LLk0IVjp2EgMw
nEq1N4owosFsqNauKlXF7/WH5nPBE2VEsdWC3gZA7+cIg6uHNuP3C2DxHk5eFpbs
8gObsm+7sDRny9TwafJogRJazM2Uozdk2LaD3Lnmov1SdqI0Q6R4IV13acY5E4zp
ld4gc/OVbI6QKI4QAEKfjamQwseUyAU+dpKKhr9jrzlaWpdPlGGOwv8TtCv/eTeu
Awg6g51Y+d8JG88xxi0MfCqvOA/HOWul23IhYaPIZDpXGI+zc2x0lfGWwaF8rc9c
BU7FGoD/WeoAwyhMjan/gx5jbx0sxK7P9jtzi1w8d5ldCnX0yHbUG+u+3Q9K4LQt
evX1Qu+3hFTqV8pyYXYlJlmAlH0EJZfWBnJf/weTBqhHSV/8/PXWNRV3/iCoHkgx
TWzBvUxwZURc8vactwd+A0dZOorLDpehnqXogiTLhEmZ44BC+K7cL3khhfk+P8Ud
GS8x/6xCUys1rklCaj5Ff8DKJmL80RoWZHiqgoq1Yp+tLosTGdsVVFhiBGW4zhWN
Fw0yCdKwYkjJGNGICL4xFdtZH+D5+2s3cdbsTCBHLMqCz+o/a/+SSSSbDxUeZkPr
QzSZCQNYfT5X81+rd+WHC47ivaXZ/pBTZje6oqpMdD0Dm9d1jw9OBbZOk+q9AasS
CdcngSFvASrtuGhVDN0bkGsTlRsH8XN2bTJ7s/1806cuyvRHRqrA7T3x8OjtYnki
QQfg+uCuV5Rr7G9w2vGpS8+OtLhMSj0SDSp1DuAJ7iVJVIH+zm9aIb1EwSu63RFK
x3e0o5uBaPgRMDT5yi1Laxaw0bBZVUQ75WMx93DG4HMQWrDSYFzPNh87oZY/uiZM
j5eCX/CXvcngukiXtJGxUhLvtaxk21YCQPyZTY1lW6g+61JVNVQu6d63OJVmYn0r
JeD1SD7zDg3Os9+xFCrQg+2rS41ER0kgA5zVfe0Og3Zk5p5TUdQERQ6gF4DdCooV
LlDkTY2Yr8S1kmVpJU2GEJZvSTx6KU7hoUXHpStG5/5//9sIjxlv89y2xk4JO0I+
5HVnDuI4a3Eyr7+VmC49GQKiv1mXSJdHmhDWfsrjo2XeWmwTrXjahDXRn6V8aRDL
yAXRP3Uf7XZz84dqOhiy+RYVTwMYlhamDfcF5DZplQdlb33HyIK7EIynMYT4phDX
WtaJ6LrjiZOarfcj0mdxd2gzwQRYPHY061G4/1Fts6yqb6CcuqCV9iMGz542ieUt
xMywmLz91DMhGQ1gkruOgTBgLVv8bFia9+Srk4RXTe+9uluCJv90llezMTptTtO3
xvuJwvGR7A2ecb3l+d3oUYzramrmWgGIv4yAxaNmB4EERd4vEQAmDqwA1zO94qvt
oj0FouV0bbFY6KEWHs15Yx0c8cSB0CyrQ5ejRxpTOK0M2ECIH23LIWwCSeh0QXMu
loka0m3LeMicF0vex8wCeQnS6AaiAm8t96Vz558tewbZOOcVFU+zSSjGRGCsm/Qf
cs/NmIpey2LtrXV8ooy1kJXdhaJkkjW5VLd/+2pQHNqENV4g2YB9CwJA3wyXw0rI
GL/Ve0uBOqnCs38AaQVx5FZpGk45leui6uD5sUQmGtUPmXNtI1Cm6nDzZK2BtAqp
DLVnapGCxv2qqbn/QtzHSleqyV3x+pnWR5DKRYCXxUbQBMb1P2du3BNyAa7ltNco
bL7hWffuf72u9Kh7AQ0+EUelK/ZP4yo3w6Xfru1kpRBmfSdx2q2k4pmZH8tfhKTj
kfTBK5ZpbA11G3bb4zhbJLlg7cw6G3r0dZYbEsGHhwEuRG9RU2stmmlci3WrZ017
51miWPk/L8mUGXgyJfMw7N08m+eIDSQ+DZHqjJMZIpd0PnrEgCVGACWiXkIvozbF
On+JUQBDwCKP5ZhjiLEM1cQmB3S0kTXZmHdCWPyy5j+6Cl4ZSr88zNx4KQajNu8e
z1wFM3Y+HFtL+0BRElnaq/Vk0qpK+x/+wj/BhMXVntQD/BMp9gyvPSlUb71/O8kC
ecpzdSXiD7LYCJOFx+sZEPGqqL70YlUn/udkpljcnB1ObgW2j43SMVVdlPCkXkOR
RLB5kiuqCR0ReEf1VaddjhMjVC0KAodOm+d3kSWDXPL2FM/gDY4FJbuL21I+JRxr
YUwYTzt3zJxeCuBLrOQ7BHowlqtYlrxuxrKSmdrIRz1dFhmfuySottGoZ7/apZFc
6RT4Wx+Ee9J9V2/X1j7kuVBLcAwVmk/3DzI3b1lsVffNg+F9KhDmlHYu12CB57yg
clwFjphUT8c58Z2e5dYqmjcGxLDkpBE/anZIKWlj2oX5Hj56xXEC2UT68laCdStu
KUvGT8EVX3x2ArMxWWaPz+tN70ozBjR0hkLM2WGdjSlDI6aKSqrlkoWgpjqszYnd
fZHeHmbn4dyOmHin49TBCAZ6N1vINu1ro8gkVl3rj5ZmOwnGcrc18GQ0Lw5oJqR5
EgAKk5rAljjwLx/H6fCVnhicCkPvm/GMU392tyAo/ndBTXFGkFIS0g0RBdexzRhJ
73N5rprQnJUglpjcOvXBkQq+aSWRWt6AZ63kxuKZsuvozFBxxGxV8urJvZn1YNWf
etPYLGmid7qAO/IAk7hrAlbx6CD9DXwVrxi9wdSHt8zYZEwCJxkFcOw+GISoOMbb
1HNKvLQqR4sXxMDPUs5HYDuLSlg74wR2TIyt6ZtPKfn5YzPIVXy6fnjBHiKgOWf9
1FtSahHou0EaJJ+rXKGK1AOF2SoHqvOgBMXnrMu7Om9+dGOK4ZadwdKMa7hx4wFP
/koTXQb5LYjW+DBGXEnfDR1zAxbAwXNm/r5ckyuAfySYAfQjnLP4kFd4QFeHoa31
QrnHM4KX4ccgu+akCrssvCuJfuZYCWYR9GTllnhk61TonlAK7k35nch5MmFd1pxV
AU8x9HuDO6bY7y7Vqx48R1Z4OXNFyBIeGOphH7P9lYlf8Dy9nV5V6Mg/xRMT6AXL
dwRkfuu4n+cUgxPI/Qo8387FAtBmnNDe93KuIFIVYP2S5M9njeoMOXvKSCIkJfhB
A1G60NPVFIvmrVyTIcZxIAHtJk1QLhCi4pi2enwROs158X/C2gZFYs743xc45O53
KafogoPXj2x/JfIyHTPd9DysNOtG0pZ7D6zjhm8JrEDZE0I4AkAfMMcfDl+Tq2Up
4JBaljCJkBVDTQFOE1YZV4W4m5ySdRutGtcsHPSnCyphU58MuraKtYRYVvz+W7Cp
JxKXEgUF4CjC2N7HlBwi2dSwtJleZkKY/qdYfxcOnHHBfquAtIQRblNEzVQnWMAO
hvGcGKPWtRy8Nlw0raeowJR5jZNpeXb0CCuHC20PVZx/y930Zs31BTxbkPSiTGkr
lYDZDmao0FmGP52O+vSeUgWTJPzp3bdJbzZuWiWi5s29nc19G7yopT7/uwCTMWv4
5efqbyEgm157vOtnne0307tZj0oWqDzVFDohQNM/OIZ9+wZABIiYp1YaoW4OcxH0
WU8IsyOuh/ykDhl5rpH1gNNufmYym0/3mftNHjvnQiOE1B2t8GvsKpNYfblCsu8L
8JC0jdAklaaDrIS8cbDIwNjy/yF0hMn4HurhcHCmKP1h3kBfhRmCt8er4rE9lu6A
GB94ppLGSwhod7kIbMbyHwujZYh8YE2zjvTrT+7U5SFhThjnF5xUbYSCQie5oCnM
FkklewQoEWdrOtRaDxJ+MFwON/mGCo62XhSYN0UhU/BLwJ+9Wwon9rChoVFYrMhF
+I6xqu51obMVtvyradRW3GTvAK2/Aehs8P7Uj9Ol1acdNMjdxVX/IV2WU8QT3nBu
HxxG8SVsE6gE2AHrAWYNLa7P3cmcULmdcdwwYpZr911s+1Uy5ftHtLlVTDQrVdmw
23HMbndcWAvXsI0xxiiu0iwz6BkuLWAzOqgj9hA4vtTGemhTtvSQkWQ9crlAcNmn
cTUEyEp1IWHunsHvKJCz234JSu9ks4C25qDlRY9ysr1RS8Yu9noCWt9MZDRPrBf6
voFXZ+ciAFunVkeNJq7BO2HE/TPnlURMK//rHGWkTXIN9pcuTPAOpHNNtPSm1JPR
I56VbG2r9770PpaigGdgMxU0BrOvHbCo2HOgskEAJlw6LfPex61aknKERNSxUB2f
VhDQ1yxoUaOU46XrrED+bWwOMzXUVBJO2zC7GkNQ7tKi1nI7qwJP1w3GeSSgfkBx
7UnRVnKp2nPSqN5jsfMxeBriYzdl9EduXGFI7ejG0iQYUWX9H+zuwkLra1eHib4D
76k/eIGfttrcGgMhnNGp1H8I0AtpCUke7DlF6MQ7YDXIb5gPuVHNA033ZHoXsKbS
bZKajSy2Gwtm2pZsbaC33D/YShOd89uZgIdt4DfbBgWOhoOAFXhweRwoVZD17q2s
Mjpqs+UqPyZxKxm04Hmme8UsxtNp75eidV2ejdz8eBqJlQP0ZepkUBZdl2M0zZ7C
0Yae7rew9s2u6aMNMoj600c83botcttBCW7mr6eyE1ynujggwjsNV20ryeQjKSo/
moeEKjqyLMN7joZIlujvngxbmyQbm3uo7a8K6rx+UPapVyAVgJLPDIHdqMs8pU81
zNrTbjlmCOKBRh+2qME4a/emEO3qRLJNbYhBOzTYPA4jKzUZCzK0g4XHWQhUnoFT
ja0yqntVFh1MUS8o0bQu9A9e55pe3jl75NZmkLfZcQKWWyy5D9aXm2TAZSgy3FeQ
aXmFGp2r5coBr258row+U7Ygp0AkFecXMApURwFch2ghByNBaRb3mku7nRmVdHKY
jCgUWGEnLG9TYmNZUErPU0cK59V12s5HPtPY09vc2nn4v/V5KjklZLckcvh35RUg
a+DTEJZgU3wT1rsm3hubWEwZP04GHIN/gLL4llHFPgj93tLuCdO/pOqFxqEVq4XK
LXWUTQWUmVuzuINTBQ/hcgRJEm0Uu/kNX/3MLrz5A5wU3PaFZb/0c+k6wNROt+WD
LP8w/C4FLHBC5dwgxidHfoEJgtjulI14FskQpwVUan0ZpYbo5Ka1tCYqOu+HDDCN
l03gWwPG7MCP7oLZI48pWTKzJtHO/W7IDJPn4JpIGEBKKPvreY2atNTNJ7Ux50YJ
tYBGJxPHe1k7QyXSSqLWdo0ZuhpyyvolqrGaKnpIEZrouiCgq0mos6iHSkmBcKym
u4n1ztZUJCTer7yMwiolwlFIaaxKtbGaE0uiCFpw+7TQtXxmyOlK1Z0Q3Mlq4krJ
d1PpRgAJSpPHit+r23pkwYhrEDtccC5bSHPw+mrxZHTReRjpv5Wqh4B7qhdNeA+j
jYWBKE2SLBt0DPRtTxVNsRnKOzN4MDmhF9DBaxhcU3Gfr4IRxbotR5mvC+Xot7HZ
5fQ1SAPSBhL8ZwWDX1NXlihArexb5XpqE4gQh+fMtZfCU0EcYBZk5JbCAsVrnUxP
BOmdiEU9pF1TMs/OXKDyPmZEUIInPXK//lSdTMWkF6psj4LVuMtJN27SE0QDhFVl
zaoRck0hk8N4jVFHgI1rmKwRqKCBa5fspfpkwa8CLrPWksDpwbgTuScncEDLvOc0
bFx32o9F7JSQAtFoRuduLLk8AAo7qZajoOggVJlaY70wFdi8ILtRsSDZuwvQIKci
2oLr69gROb3NtGcM4ARaE0c2yvVSjbjrEb4vKZNLLySIJ4r2BpJU1Oolo5BQxQBc
SXGn9jMQ0qfEe2wktHaSzqni6f/zPkTRHVYPE7G7Dyz/58cLlDWnVMcCh5fJEzpj
yP0OSYjqpjCMwyt/bP9TVW+H0H/UyM8jB4mX9+s6jT3chrlbCQ4QV5yszk9KdUcs
k4e8bVgq1PPrrbGEAgC2Ku7YdZ6CsB1C2sBwRvhYnsJQvwlTMHWTTgqYrnbw3eB6
qz1YUMpA9BJQ5uE6BozJu+B/UvfI/L6StmwKIoQfrQcXU0+OJHtE0O8JRwciT3e0
MjrF0XWc/XUiVYebLIfLayoHeCYtYB1S1OG6pm+E+sAS0xj4pMDHH3raT5mgDOxy
jZsqH93pSrLIc8KH7sJS4qv5EkolfY5bnI84f/5+51XUh2d85oflm9DWH10hysKO
nB9s+gwMSQE8PbeYMoI5dIRIGUtvce7vG3/1Ka3o1iBNio8qm7qcE86W8gIE3fhg
fjKJqQaaCR4POPvpIc2UrDsy/7Ou0hmsvLQrDdlUaneV/iLojDBrF9wwU9TuNoJr
znQ5EGrpWYXnUbwBqNIlIID2sGZphTbQgqfGksLZROMT7lkTdQV5xFDdRczLkelG
xQowlUD8taTZuUK0VZsSPrI8l07CUOTqxyRh8i5h1CDrZIdbOosn5ae51lU9YH0b
S0KPfu09XhOXvIvfstXOPOjyzYgkSofPgVL2+/EC9ieg4pImfd+p0U0YOHuDZdbZ
Hb6uLeqxiV3jFXzwpFlDtQ5TwBkmYFjyV3WmZ1OvZAmPf8bMxsnVbcUym2E+Pr9V
bn6ZCB9peaeGpINhyVko7BjcL/ToP0BRuHIu61i2IzcNGfOM4qZbdQ9tzY8ygmLS
JSAuLHK63lOBO+i8ArmwrNNiPHAhx6xNuycczS32fh7Kb71hnscw5L2R7/qFWqjO
Nh0ubbTjl5HWzYKalzjD3cv4iRDW1Li9isvBOk2GgfCZZG6vFAzO+KsFhzrdUDGA
aEvwRdkOzAk05bTqeIT2VMXRghVcgeUE5YQCW0tmS3AGlCP0vm+GMW6TfjnkE15x
d4rH939FY8yeUFMd5FAdBDThGJBkVxxkOBPB5gtu1y9V/pVZBPtFyvctgC/SciXd
VpTc1KNDUtCyMEziKgqYylG5FpPGIlWAJAS9tK1m1WHJ2UKc/jl0+Y9siL1xI2JZ
a5F9h1bVfOt9OxLqZl1J6/i4vdBgZUpAEp+9wWQMeCEZbYnA871bCNiUqtt4nyx6
hHOlZX/KXL3HxOkaYwsdjWql7WMBcy0kC+qXOsT43/Rmf5DmFNshvMeTfnCEclzF
9Cjqb9eMpot3vx9G5vqeXqZarR3Wh0VzXyaGXtBznYAoMuQvZKzkNO94GXrcmgSR
ZhpVEZaJ3sfkrNMvzqVWIACc3xwQk5lws9xYp9A4b1FZkA9dxkrD/mv8depcAlMP
vKPEmdJkuTiXNijUk/b5RxmA/SNQ7tJ23WtCJgnO67WmFHWf02XDYLS686cPKgST
wn6KUD2HTt5H33msapedC+RqVT+MVdGb88fK9VHE2yXbJmMWoHt+uVQJDSoT5m/V
L3sguiV4v2O2QLormZLRlkMa5vg4jftpaBNVp3K6F88tcibKV6YcFe/udNDFfnSB
PCYUHMV8jtRP24MZEc+pwQPi0dQmAnPA5rFp5ASlH0O6CvDFF/aipWyIxYfFtOIF
SvjmaiqNCVXNiJtHLlslrJ/4tTVN12SmpiqoAEgvfYMeO5ERQKIiAV3GhyyXGLI5
yzW10zvCG1+sQPJ6yW6sx1bpMziJZDkZcwSiqTSqMXLmZcdpNomOL6iGDJ4dSaZj
FSD8I4C1FHY/o5o+fg2MuMqh7WjzhG3LNmk2i8HQSiT6HuPONgAKT1q13U6YMwIM
sHymwqhvo9qpUlaGp7nMzL2QIvnklcX3jrOJV24Wk5R8YoS/mJ53s2R8AanapNAf
cgYn0PVdzgklpAkLlGpzE+FQOm1cgrbEs5hBdbjZyMrFgNSFix/XxrqAQ5j8EVGv
1MyYJg7scZN6b2zA+/oUNZhRY9HFhpW6eDOavUDukLFp07oxaJDUQytPrrYqNcWt
OLmpOtr3UlS6BUY0M6OGUZXvj2Ozl3h07rbzV5UrTuyoaAHKe/Sk94CC6KZgsnsL
LPBrDvy3Z9M5YDhsGT69MR/aUrjPsL8guYC7H/dqXl3A2WmA+0QiojE+PuGDkF27
6/2SEFIDIzzzjUf3hhUN+aFNLT0fMYQ5bOjSLmMkFmn3CfJCGtXxCgMDIvQQFwZk
`protect END_PROTECTED
