`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qolwM8yc3dOBw8Vv6u65GAwdpew5M+oydxZJEp2+NjJYSqE5eKSICLyfW7AGqmsn
XFVhxPZiXnpQoVXTer0FEOYagR6cr6MSHsk4YZtl+zJyfT48O8sywtoex0i51zQ0
mW0pAtoJ6W/4C5E25S9pvYU7+/Eq0q51kYB5DUf2yP7SNnsp4vhNnuUB2YXz1bPX
zabRPe1o3QT1yMhpJzZSSwDr3yd+KaF8dDQ4UHSIdg5s5knlFSP366NFP1B96fT1
QRFaF725UB9G91i1S9OZ34RhqNsUn72IGx1DZMYO6SjUX1rOI2DcJlx39xc93JoZ
q+qv3gKTfSIaWAjfcAFSZeKl138D1GPvkv3OeUWT+D/NMH2+pJj26+2h9dYsGa/1
YDVec/6HMtKzXWjUrbHLbFcnxQjRa+kdDnS1PXubDoF+jTFQTtiROxE+k6m6Zirk
`protect END_PROTECTED
