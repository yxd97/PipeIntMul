`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
57tQwYzCNcF9wDvNGg3NxLcNt4Zm6hJ6KfE2zVXyvHWLm7uq7q40S9cTyKxVqj3Z
Om2BwLK5BfzHn7WDNXLVt4HIZMfn6XhjXr/+1/SyfnRYaTi+2IaFv1U6psYLzGt8
h+oKsemoYu9ANNFFTgSD4MUmZZB9cSv1ZfBBrxBDzYMII6VgqP8qNpCAFhnBr03f
hry2US87sYqw4QGwzF60SADG6KmeFTY+kgPc7u9A1W6jrwyg4DxbAl4XtggVk2mQ
Phj+TwS14wpdQAfOKS40xL54As0l2y48OpYtptpBtlJh4CRn7XXdvymRd/A8OKU1
1n86NDr0locStIsfLzE5vg==
`protect END_PROTECTED
