`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xTd17o3musbi92gGmJixudbHrvgRArqIUU0o7SJdDY1CDRRZvf2fMCurV4uSeylJ
+wcuZTTxxH6p48nHEPCDpfU4N2FaIDSVUF2cwEKmiASc5nEi6bt9LcyIolGIop+s
KltUOfqiPszdYxTMUQ+qxbnreeuxILHSuROQJ8iySG/rqCkMTsaR69SMILX1TEbJ
fxfVyKsPcWfZLp0k2EgY4ecRChJhiLD6hOR4pIkCtH5CO2s/jLEijTyfSmzuV2Ug
l8PVtSmFP2aTEKCzUB7u9Nz1+muhOAYVA1R3Nf0+9gqqb4wX3yo3+0UU6SlNelPB
`protect END_PROTECTED
