`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
raDQMHkePtSknSxwlHERzjI1p2K26e3/Lu8KIfa71ABsy6tnMmuJiZbaNm3M6Hr5
HGsZm6094KaxC204ePA6M6mMPhdKYhxNOnKIDXbsNJL1v6CUwiliFl1bDBoUsaiZ
YGCHhqMa0wfZLsweol+M0zMeY9HKrgINBpdbpgQ7GEzKfQEwgIQDPGiwCrfVWkVm
HqswDMKh6Ib4QEo2lrsTN+F2zK6fBW5eiyPSROSQY7FuH+nCt1dfhYkpyjQAV0D+
2FFBiX6A6ZxyLeXyWCOfl1svsOZQKiBiT9cW4YjxlJ1FtgUOi4aUVvJ/hxTy1OxN
RFwDLlAFachTBTdzt3XyruoNEs/G5q6Js9NCFx0nB/tjaJLkaA2DijL8hnNLbYkq
lhlT/JKVku6fA/W/lhEe3g==
`protect END_PROTECTED
