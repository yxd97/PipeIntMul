`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MunQU4ewm/CoKtWy7mK4ec+yaz9UAIM/FSRT4eSB74pWzMaja7lhNE4AJ0pIA7Z/
VX5d9uyt4AV5IWCYQgd84jRUvO7Vf0a1kDQNpbNHKHrYhxSBrZaRgbihaG9y/9FR
oIMWonXnAafhfFq2luR5BKQ7TtoWpo/z/1JJZuGcTKncR0fvILo2Jw0brm9Z2dEA
ph5tbUafOlc3Fy1MMyUZ5I/i63YaO7UUxJ5FTdEG2QCzTm2Cf2XwQMdzqF7fpDDT
6Pi3+fgI2uWIvh1BNY6jFRe4GrsOYDeEPYHyCj9VfsGEYu5k8XQMQAw23wNDFHS4
927GeHAC29rhh9EHcaF2b1+y0i6bv+dFhjSUosj6WG8LKQ0Ef7klMeP7XgEG0jlf
O+tW9bVldBCNQmWua8eoxJ59Dg7i/reBjTFb/3GjInJ8BydiVu94S+ubTJ7Ue4zm
vki8Uol7XPfoTAcnqRSaRQ==
`protect END_PROTECTED
