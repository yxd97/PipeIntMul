`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LcLP17K6sXAyHLrzYoFYixidUUdRUIo75WU6tE8fWRsWVk8ULvGXEWNZ6HZyXpGY
4gfpqtOa1cpxY6p8JKrPxzySNMdebehMFpv936qYnWeR8SKRv8W+xRG/QymKpfps
AIDqhtYMgePXX3hgfshqSpUMgayTGcUswIWmydRg0BUw9G1/nRVxpD6z3hsuz7ix
7sWCGIl0yMMPCe7ttCVf/+eOL/TKDpzrnZ2lNmcLv+/Hyc48VHTsdQugVr99Hg1t
Arr7RV83Jfeab3vWVcGY3z2NaHTXuCFwyQNnS8gbz6vxnN9x3c1V0todmCkL5CPy
r7+yeFAeYzZWXj0jxRpcdQuyUEpx5JH5qm0gs2TVU2pi4gHLApAsiLM5b7kbgjP4
+o2Cf1Vm6utsj+0/9QfmU3oAWiptPCcUm6Jqb9YEltVewBGIDZdTyG8iBT3nUyZi
041lUbq/G5FpEFsALqfQDsuRwrfB58zgp07AJ4qfwHg=
`protect END_PROTECTED
