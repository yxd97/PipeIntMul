library verilog;
use verilog.vl_types.all;
entity CAPTURE_FPGACORE is
    generic(
        ONESHOT         : string  := "FALSE"
    );
    port(
        CAP             : in     vl_logic;
        CLK             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ONESHOT : constant is 1;
end CAPTURE_FPGACORE;
