`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XSuX/Kryd+jx+UEVQ6kCuWuywUZZh3/leutYDY3OHkX+bfONwZvw5N13nQRBUSX9
oxIUcsu9bmfKAatotU8jxnzgNIQ9X0avNMEUZ3I65HMPUpjqSnxn0HS11l+cJbAK
nEEVAzgupvcK7r7GPmZ0MiE02BuVAhP7AToViSvd28OR4B5zBnKi/YVsOHwL91tO
AuOVgjoeuwszNDXnPzuRMAYF2XNDZkPSjEdvUk/X7q5GCQd3ZRCzCet/ZyIXcI/E
/CW501sqpfehojf2iss6mpjnD+3fcZzynPTWlQ9TZjjdY8RtyAA5w4kDhzhWw9vk
6lk8nFUFN+jRifH0MIJQXzFqogHgzuZQ/rS2QQytFgA5lIzvGD5q1qNd63SqILNE
Dv2JgzXonitETaAtQ5zo1wglvgvSWIJnjvyiBW41Spaip/ISdFlqkQKgnzDmOOF1
hXrXnvAu+a+grcBoNBSV40dxnTOg2RS2ZbblIk35b/PtPlhJ9nICaFlV0dMr4NCo
`protect END_PROTECTED
