`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NAQwK8JWslxKmQROy9MflCr04uNzn+jgdUyxPMnV3cLG1Qgseal/sGEwU+KMDkos
wsqrnRKDEllDfqvDHyqTnAgb3qFvj1D0xPiJlWQIUKC1aDmEkiHgUIyuoq2X0Gzg
ktTUoe+aOpLJVgkX4QnzcW8T1vVj2aD4cg0d/0rL/0/wzaxtR+KevWnj1+06aeoa
UQHA0fpXkH974JDrhFSOeNFSQSXtk7V6e7EtP9bQ8rXiE0wwmsZk38K7ySi+AyUf
msD7zMofCMw+BsaWzKffDA==
`protect END_PROTECTED
