`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sPLqZ2pFgsEZY3P073MkJArt6w8+ILVMkY5ExNoRmJDfp20yTs/R/pX0YvSAt6QW
KOxpUjzSOnDs5/c2vI/TEvWjQX9ICGFSGxhDoiAVY27+klbXHlZfumdJFA8qT7+M
wELz8w45e77nNa0wANBGWp/w8jn6GIDySB+BxhyZxTkIw2uYLc05p05ErzRVKChu
97PaSVdz2MF8Jisy8u7RL3n5rlR3RNMqRkECmdyT/pqEMv6ovtkuGY6K/U7/b8SG
x18+ZTPRGTuzsvBhyvZM/esZjyf+BBoL1HsxHZTGE5XzU9JVIM5uYpOf2+waNrMk
bwOtPgHiQe5H5D1FKpUvQKFY/FmlNz6oEym8/Sp8EI3K/uZg5zfqf7H8TfX028Ur
O1c/55zT/hDYaxLgHboj8JoekxIavFmpwrH5Un1c9keFgBaZlGl1n5ZkhPfCskiG
c6VdVZFgAIIqToxVLWbn6uD0q1agQRzxcMGGu6F8cKjeE/dZowUlgKMJSHTDlFjm
`protect END_PROTECTED
