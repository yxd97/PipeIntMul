`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zx2U0oiGn/ddSguDt/Ib/3YR+uxpNmoLReALakygZV5M8E8FKVcI5TMgELfATbm3
Bo38Gqp53YAE/DX6H2bVnIR1oookqI42wUy2D46ru8e6aD58DQjYUMP3nUrgWcRb
NRMNyfvpP/u3Bddg/GUiU5i+oSPtc8SLC2DXQkcBZmqzhIqa7bT2zpZKKWNvUIzY
ircdRND+/8XGXEGaXeCeROKDj+z7/AV+OMjMZ51Fu85W2q8hzJffax0AkroyzLsF
wfCqBAsBWAtvwqQ9Vq6cHrYYzORBQG/JoO0QEPpNBjbi0u8ohvh/MBF2lO1LDN3F
Xn3UDtqIUuq6LwN4vh0DMSSl5MLKOps70/M6aIDCar+0xRWi/nr3bBUU2/7U8U9L
VKe7QCMz3pLI1KKLdlwkSjG76T4STuFFyyFqEw1fqjfW5gvtKBP5ylfe52+HKo3n
VnnUt/73CSFqeads1GjRCipVKZzOWsB6XTl4BCp9A0dLa5uCfS50YgyLyTzVLjVi
e8n0skIgmbW4C8Sfx28/mR2DUM5gsKwiiCyPJaMD5IVPMiKcFFYLfh/Hby1DVzmV
pO0PnjIhpQ1wMBeGom35Gg+3m+wFEcRxgkGszZk+wiiG4KSlHwLghNlg6CpT9tYF
3c5Uy6BHpGyaP58JuHjj1K8/q5WpMhtBxNiGX661J5USBTHS9PfVzZQ7ocTCgGxS
5bY8z1EbL0dN8xrzNlLNiPVTX+3+oDfn5pWusvrPF7hsmKSyfsKK9MQijrTkCPxU
VMZxlc7s8T+FENFSS0fQkH6PtALLHUU6l6QM/ROlzAeU9w7Dz0l9VbhDv8prK5nD
9ojpSauCNZYmnZ8Rv4f4PBiippNpjk9sMUNxwh+f5vCzQZmLupFuEVRlFwfdNV/a
0B8CPJlJS6Ukn0UW7F0lTvzM64PjTYGJ50inZZgZjKIjNVsRosjXp/wg+50VsQL1
6if2igiNYhsPDxMdj+gIw1CAvLRv2lG8o/Nbp4DmjQXJqXu82C+2jFXUQ/jNkPVk
zqX5P+QxpsSm7+uNgbOUzOrwJO/UvM842RKH4d2hr9l+9EaCyHjN/I3ARMrkwDVn
A8hvCBeoeYnf1n9FkFrXtkZjOPVvnIHJJZHwlWdAJg2psjMsSwcmiNpupmEugI1r
OjzRK+lHFSHZjv94IsrAgM5OgUnHHrUrjAoFVB1mGMBq/mvFVK0+FAe01+UYbvsF
7CPVOaSxAzrTZf52/phKyNrp7Uz1BuH48ETNh08Uc74vk3GL/VJKiqP0KwAmrtG/
RVSM+2CVo+tF+Fv0nuMXI1hAr6r8+QFNZOh/ZDRN4mLvvCe6rI9tUzIvl+0S2Q9X
uhYnP0/R3RagmStjBE9jsGeXMcuPKhNLJzag86+KgZdK0gB+/BaMvIz8SmLOJO1E
3H3aB+/6IQ+djU1wT8s+lO0RzQR1WY0ibG/ErzQcDuas0IrLZJ+LFXU19sA2xr2C
QGy+T6At0B79Lz/l/YFytisgAj0foNSnJK7+2bvSdl9sL/h8gQmA6gVo+OWO9s0n
lRS2P2inweGWgNvadwAaGMltdTxQs943xhJ0zrC1wHekAh0L/omX6OMUXiJcFg3J
TusvR6UeKSWM6uJu9xqebMK464wUsdNxibiTcQKYCsKqpr1SbS+PrPrb+9aHVNts
4obLBVCKShlqa8PySDEXZTbWB483uO34Owl1sGZI4+mWYqHSpSQ1diMczbcYhDrs
i3wawKvXitKkd3Bksq8Y5rg+3H1CH+zngA5audEWJPigPoBEl3uP6gUdovZzA5qn
sGiLsN/NMeKCTI2qOmyy7K3GScJ1f9gyD1peljgBmxx8wgo+GK/Co5WZRoTzKsal
bAB2WSx/HE3BJsqjsqw0JYO0CIblpa+LoAephO8NaHV1SpWsyileFxo+e9CFe4pq
1SsxKgofu0i0/pxlZfsMq/cIODSPFIq9AoYkjIpjaiN7PN3ckxxZwhSLc7sPBsxM
qqbdwM1bCjUSahGaEqaLBK+uMQirgStqlffhuPtCPTh6t2ZUwfS+ooyskTOcD5PO
PvKvpNkigiTLtDzXpVFzxReq0rEMVtwqHbXakfvjmLdnvVoJbF173K+Yptqh2Z/D
kGVtWg+xS20I4zsXNanKWHU6ytashr61MWaA1Fq63hlY6lYa1h73dtfALUJ8vxnQ
FqHtC2DX6xr5Dd0bIJjLxyUIFctcsUAOAog7dRbYva7i/8yBbcPMwFsY075YII3y
XYy+1wmYQ9DIAEpVOpWFalHbWkEQyUutbU4rCWafo5nIGmJ2zRVsxLL3k+BYBUXE
leDgYqh0m+vnc6O9T8JIDh1N4sjgNb+O5/uPWsgn9KQcBhC3NBCIEvF3jcpgzTya
E8e2uFAIj8L8qkc9qNIDx7Gw0XDlJ5YxLvxophL+K6QoCmr0K/7NfjYkbL+zDvYF
0EeUu0C5AovbUgKBwAKgfIG71p9Efe6stgv4Nkvu0293DtgXHymbER01I7O2Si1N
HUtZhAN5qxfLB4Xsy28CAcTe6Zk2OXgORsv2N9UK6RW6qwukjrL+GZE8BnmPa+AC
q9TlbsJ8r7D7ZFcZOBAqu9TXlhM0gCcJ9LkW3bUlAFYiN8Oa+nnV4YriwOv98cvK
fxoXf7FfyHF+r1KmgOf2rlcBEddJElxkx1cSXBZN99N1w6We1cMEcIYuW4a2rMn4
WCh2lBpuw6WJ4HWxN6IAZeJVfjSmmTsjvIWIouIssvfq5cuByezHM6HrZG0atW+4
IhMX8YRuw2gQLld2OCQKnBpj9SZiRu2DXRp+5GwpyMFdV3TL7suCFpPacifWT0JL
jnr4OiUHs/KYA3Wf0rI6iH/0SihmhPT6PPCoJqY1jM1l/xJ3HFrqs38QISoIR9kQ
BssEiNRvef0bD294LZYYdpv5l6UOq3gtsgSctm6LzElQLLpcW6Rk9T+ro1GuD3Vc
Q/YBRFQYjLEPYSsMV3jE+oZqqkb9UDT7G7F7V4qO9Sra6TO/FZSwTO7cEEndnCGu
qfmtQLiYOngNkr3CtZ4VgDoDs+KudIGVXaCZCX/dhzYQI2m2NZH6P59wuH2Bnkqn
UBFHod+VZmWrrF69nd1ldxGgbu2T2POD10ONDbttRQGILj2ExC7eFlr43u8Q8b+z
K6/NoV9yFSNazMTokBDJgADj6aPbL8GLyWxQjyAqMe0H4OGYaHE6eUH5NWbSMtNo
5m2Ad3vn8VKwghcLl9G6hnMy13xtJ8ZnJMH9NwqMmKdeJLQW6LfBDBEgVUcz82vd
WI814lCy4dEgDJA8jGWU1hYzcMRrcTRa8laXwZo3riClYlopvzPyjDuIs8PSLmrf
SoWdMRY7AuxT3chm4b1hie8S8e96G6pa6Jd653fLa33HKrYq4VumqruEfXj0Mk9/
VXkFV48NRhX88ig+rb9Tsy5uFA0hH0M0UHIXaOdV8qZEU9o01GMj9WYtjwSikx9P
zmWkAlx0iIlab5K39oFlBYMr+c9hZrEfcGeiAasaPUYEcKgfntP1CBIQ35PJhBXC
MQiXjJkEPsE2SPf0OB0TY2EW94APKEoBI0xUXX/c4wv7wma5A0pA+HUqZeT1lHJL
rFsK8LDVtj35XJ+beafMrMZOi8UzE2SmIo4E4sF2dgsLNBA8sRRfrYyP7Q629NnU
taylzzcmUkgxce/zzQMyHVt9Y6GSYVZrsFxtbUUZNSv7YalvSax0dMr6ucZDAAZD
0D7x3GZ+OGYR+IzAYHhQTqiKK0efkcPBdNyG1mTgJbiRGVNmRVz4+sm3/Jv1n04b
Gfrz2sR6m6VB6zh0tBS9WKkrCA9FtVa70tMrg4GkupXn/b7BixWBJkq/D//JLN9p
WGpk17CbSkLijPxY+zWu6gka1qHNpwGnRNRDj/3/mGE9ucLAbRYenyu4n0NmJIRv
ulyYBp27oEhZbpP6uWXiZb3TISbUko0HaVtoQ4fydGtBPcUYj/31ZwMDwNtVWV+Q
dxJg3ZOKI+O280Lo9G8OcOiUEKNf+fmfsl4euWGepp4/Xhcjk100VZ0CroH5WVUd
/wYCDbPPjYrpVro9rk8TN+CLLSKHnwm61SaVCq1FHEHm+RuMp6vWaeGgRDaFGnay
69c8EepIHEMck01UJKhcrOnKVNKnqzk1vW/dT7qb6Em7TyXIkNeJnQ0/zrIrpgSD
GAq2z1L5GGb11UovL6lcpXljmdqO84wXf1HKo++OcdXubJ86IYyLDQKmfQIAP2Vq
OIBNZ8EIFKtd279+8dGmpfOkGPxQPKiPEB/SJ8/FCiwArxJBDTkEVw7fT9hNxOyu
iqlCTXzufr0GOFvNllbtmmmjTPD3dT+dlmBGNiy7AhC49o3uKuwUx2UF12XkfYiK
XlW5DBfAu9DM40T2a7tbpjYE5CSdj1zXJGJY5/PBxvKwFzGWlRi2vBc4QccInpdB
HEXww5etEzYMIgwJ/LN2Mt81ltlAa0LFMyRHkcwcrzwckEmgAlXcUfJOZJZV5GRP
pdoR14Oq716QU0EbbIsYAi4hAk1RbwFbsFdA7jAAGR1w3ElFhue2wu+q1rt2vEp0
Trp1e36t5/lOB0M+dP2QYlFN04Seq4j7jSMq/9ONYF+Bt6xxeW6EMmUXydJ3Bv7P
VRxiMeicoj1OyimlPV9+C93tLrhoxFo4/5e91sYuR85tuz6dtGXpUrBwONq6+aE7
cMqTuxlXt2AULFeyuNcPhLRKjZ6oRi0/SpYsmoqSZA4ZNvqIxdVfA4XxGyw6Dz/D
oN1ppiAyOxb/b3wCFG6KczF6gisXS8Q3sxJYWwLRU2bbEnv9NoymYu/B71fhAXlf
KAelPdBIksKBLaJ9RcYMTQa2COXSff7q8D5vWZmMOz+juEYT1R8vesGAFSneWnhf
I6kdCuE+fI/Dyt0vv/oZnuiYGogPLoysHmLDejeOwOW6FzAvXDOSHPUZpdRO/dVR
dQ35uE2JlAQAozuq04LT424TT0p910mgYIw0AQ90srF2je5u9N3m0gv79E8yYXJX
n0fR/5pdmtPtRbRom+8cye9tYE+JTKUWHGf5Od9A99QeRwAx0UFxdndXIK/yNMad
fkBVkIo8etE7JrYGhWWtJHaeShA6k032E6nl50kzbkr+bRCVmLkFxZvaDlVEtRbE
7Aqr2nXIhcgXajO3hDzZv2VYn2Mb2NsukX4GxolzjpAbYdJ07VbskkX809Tkw1En
zwxvVdGMbwOjp0K/Oi2bklIDzlOI9wkQRGaBN6KtJ41MSr6MVcUBrNTewPR93iyF
02iGL5wV4QvErlRxMpOewO9xfwRjLgYBGmLWH0JInUReqtH+M426MSe6ZMjKmpOh
RghlQ10hLxXzV3AGR/W5BG264mYLr3/o3xHxAvrjQXIKPffS3N5h0Fn1PrI5Oaa1
Zee2GeHIzaoKE8Zp4WOenbpo7tYQlqV3ds358Db67/mjM/HHKXX84sRA56cPRfsT
KtqlH6DwM+g7/ImOKz6280WAteARoikhc9MCWXoWHW45dt9RUL2rYi/fW76LrmIL
U1W3q6AMboL50HhZicwX8FPwpuhMcwzsovM7Sq+76NmYrMQyfTqJjhueE2fyjnR8
6lswVhd2aQLBx8yAJZR1X7DCiSyaP5O6bL4tczFqAwBwgLoxnrUEU2/7wv/pDPb0
AHjCnOTGVaiSCe23kWmVVYPGCJ/VwTqQYOV8ZReFXSA44JuUpBvQPOpvGlN6ijsl
NTVGpQHI9AHWPh6kHCC4KbWG0RAA8OCCEaXwi5W8yhcD18+7H/DMgDjDzs8aYJtx
F3NAzb2QfkcmDXB1Yc51QXELKgcd4VecoifNkPrvQDXXLNyUJUXbVpXEW0DYC0sj
YSsqs8ysznKWJ9zbaJXih0Ydf3nBNjzbIRNObDkM1kjzGb2m9EtWiThuzKZ4gwN4
9B2dnrsDJlJDVB/fYy0Roj2WHB7fngsp4WYoXa2WfelEutco3C07zU0YtQqd/xZd
rEfeoFx6YY4ki+ksQ1hxF9pdQfy12UsnUbrOmFTvJygwLtWOR2qzUbqQQJQgXhul
kFCAosRfB6FcrGVNvrAAIiw4HsKIeRGokUAeeVuVHZLkumOUfUqAHDmom8kV0ydV
FA1vJV/o7Dv71uAR2xY48Q4pFupAm3hisghBNZBeKU1f/s0NJn/1jGmACBx/laXv
dYAuB6mn/JK9JywhAN5vH2490iyu6UUeypUaK/xZxYxVKKiBXnF6b+TdRPQvloBp
jfqFHCydNWBQ5ARQCodL0Dm5ZR85JDPQdZTK4kU+S+nJH66pSPaHJLfnWBgj0z4Z
OhjWeRvFDl9yaASMIvnBkq28X7t1i4kgGOFz+VdVtAE4makaeKFg82hXJO3iVOyX
XXsloWH7MtdbkVekuvWvpYbKKEHOg96veNWO6awxZ3V3cOzDSO5eJClAy8T9tQAR
h3R6/NswIar03b378cTYLJ8YP54sCt9dDMIsQRjHZJPsvksny9gdAlTJ+POYnpkk
JdwfSQ0BrdO49rx0vZ/E7exhSeLw/CjNigOmbaRjeGhDoS+GI8HPOIlrDX9ZVBpd
UxHFSwoKv3rmH507YxR0CZfyDaVAoGL/0p8tMdyZfmZhGkC9TAir3cl870iZICbA
a3jlI70fM0ChcrnJ6znvDr09VK6zQjduh4Tcc5tA1/gduiNQotTnWBTS5LtBvcBY
LIVbWX/1AmzeCoXsugA1bGZ+3K3tbUu2W+H5+E9Cjq7ejyLLKjNWTM5rpx8EB5yd
0nKgGOzQj7vbnUs7GAb/uXuRzymXH8Q/+rC3ueSLiXs0oKt1ad3HqZ0AuPs9OHne
gf+gjxy+tLz8qT7dDJKqWF1V3dj1h0zp00HJoi8RYmS2ESjmz18vVK6pztRzFalA
Q/Er6ZOw5KdH+JhEfPD+yUHxZ0Zs2OZTmmQxRRse7dFFrFCkNxassweHepU6jR2k
4OWLX5/nRDk8V6JRQkCkc/QKynIPz/S45VyrQwDj9WrUzFvA0V5II0gDCuIa2Lgg
vRaFFqmNLOxZF/8ONo9CbUM0rNTr9bIWqaQTThbRACrt/GzuFSFkuQEJOZGMSNew
rJz4onldsQ3d3VmAlOtNLw18onAMdzofgH18wDKrhPFohC4Lgt3V5duV9auD2T/A
RD164EtVYxAKcKcQR0p0Piz+PTTorHAtZxl+3pQf6kqRyzlaPWY+yTLma6pEpJ+H
EYJOuXSCgJ5wEa65UUY97B/CmyVVEG8UQdsF0zOvEzLmc/6v73TDjNq2z4odmiEg
5Ng33tUpdSVkclxOUme73k9tZwDJH2eh2tWabe5n2I3u4ba21plFEfKl/QoOybUT
Uexy8KaMl+bpxYdUr/weW6ouMIv+CzjPl0C+jkFB5FDZbojucv2QzuqCpcNw9NPK
P5Rg1YzZv8EWx9sFV5vbpG71u3eiP3r+Y66+qkpVxP/tiaYj5GWfFv+JSEHVqwY2
Lb4I4qEbwUKdt4SpmFFb+De0iwH00O4HPJENugFTKaBW/KqHZ9MizpRe0JGYHg+O
NuRCQrUFCs70X1C6/+w1tAPeBvKUXJoJ+59w8IiY6eI/Z7LEfCVn+2vMFRS7rcmD
yRSGhVm1YiHkp0R/P59ZCUMCep9+YlUp2WUnICOyEQacRUQj45oJduRXcnUFQd8B
4l1XL2674g4hWfjO3dTyMiL2TVZVq+DLBo9G6Yu0jlHw8ETKGo/XNHaPmmPUnOE6
5yFpbpsCQjG+kGNKpS007ZRebjJ54b2DlrmDPvUm4joDIuW+A84BxDT4UMC4+RwC
ih9gC/4jyb83sIZtlfup0fuUeiKfLBIupBCntuVGZzSm8rPOjEFwipY06dP0omtB
BPZy2KMeZR8hYA7k6fx01kj545keumMPMImC6OdZ9RLphPq7uyXhdvJ9d+Sh65Sb
3Xw3plt30nyjjd54NrUXhGa/Ytj18AiGMsv+20OZFvKciojjNFz1ZCULjZ5wELW7
q2aCAJHV+HUwclJTyYRsJfPGGdozo5pEkWAN8fKQwc7VPsrwGxYlmlr2pVR09xrQ
rVbUoWZtE50wKTw+uSahTTe1nMwNwwIrwxY8K3jebNBJzWSQv8GaSTRM7tZDbgND
e+CYLvi6VzYoHxe/pP1aQU9aISAa0qz1b2y/+/JWaXVN33+oPal2k2kx3+Cs1Yp2
v2pOpXHP80GyJTuZRH2aaxRfPDH9bEygtA1ZUomAtgFJHIrJWlef6KZFhYFZStGB
1epzrKz0/HjPPlGfZ2rkbMKr9oVcfV1nW7BKdBhZMaYrFROWb6+Sd6MHxaON0rNb
XBIeAvOgFNCO96LC4JusWuxXwz5nt9l/zwGOflu8h2VTcnaKq1bJzBIpTBhHPXNL
6u4m6IeWYcNsoRzUaj9SQxKiUI2di3iQr3tiEzWjR6r/y6kd7TAfRyW5mHQyQy6L
CvbjmUZoPWh5Qb1SB/fGT8rPfJRgzWaGoiWs4X2INNBDsQEFPagjb+7qxs3+omL1
ho+jZ2xFQ0W/2vExqZN/Buz6Z2axpejelIXO19KGGLiG3wsC8Ow+gu8xyneTr7hg
rKJ2YOQ2Sp4+LmgNVed6NE20ynQycdZjhmhlFWuPCGocvd1G1LesjmmxeM0R+cW2
8Nt/6qLxcxKQ1WeTEwl5l4tTYoeMyi+/X20istcbRKCT2klwnNBs2z23MzrI9/Vb
m5XEZSTkN2amCQGZS3SXT7QB+47yYQfOEj8Qyc43KB8tQTKrBj6M0InWWT8vxpRa
iUfIIaszCym73SYieCtoumRx0rGYxjodzbp3TuL8wz+Z3CpXCv6M4q0CMwcXlpGP
OqDADRxIVWwEqW4Dn9MZ60RacwiGPsX3rPMBaiBejxKb5co7zRIoDOxuIui0a1zP
ewpJ4cf44JsqfS/742+WPrYUR1c8MfwALg9bXR6TCWyATHVm2SMK5wkKGommjyJD
vAF6Bjz1BY9Z3Zbsm4QTOkTMKbRvYAP7RGqZjfwu0EkOcZCw/vZqG3SUtk+7Xwpr
eMy6w4tOkWgcd/qEVh9lwPpPWiMDJLTyQNbp+t1ztP3pW29j6jWWvZNRqHr3s5aQ
Y4gZauxg51gP08mUmZ3AwPQBQJmoMdVtkABFnAiwxkIcD06eqrl40GAb3XyM7Wnj
i3DeUQrk4ylIXA6GUcTyLcKzjp20RloaFstafT/6S+cDGX62iespnL7qlh9Fo0VE
3e5GDe7EoGsdBJhTwrJpmPsZPcq2weQeLm2WbLh7Vj8u+KfRUL9fHGMaOdNXiYyU
Z0jPoCKwi6DYoNNgUY+k+OTa9L15PZkuZXW82yT03idYcxFh91Aw5/Cg6vR0csGH
OL4Lzv2qEJ3jldKXA/fipwxE96vcpVmmm0xSm9Mpxgeh+k1TbUQ6ULuA2xiQ+g8u
434cp/4CcLCJE5i6R5zFbwciAGlQ/U5ZjCogcSrDXsHpozqRJ9OP4cj7b2OxYdiu
9wVhIKvEhTAjtg1h1AgYUrTArElmWUzNYOJqg3mnU7fe2qWTHaxhJNJBv2L9rp/+
FVoDG3zYSGogkVPK9CDDc3v6zWqOF3kDu3lgoIPppQp0JGyoHD4hJLdG8hOUFff6
gqNHsWoGO2M4AkOBwAwaj4S0lpoNINHlLm6p4aSzwOJzXL7BEdfqO2jhkX5tju+n
xwoXH/xR3YFKbuydbj2KzpQvv6bToHbY0DCWK0EF3Zq819wRXo7qTJLiQoDyH+xb
eiNWhfS5BowMSyWPQk/AXxf6u4Pc6CSJ+vgeYBfDskkZKTs6zUaO1GsHVgDYr0qP
8tFTZwEHch/3jSZ7j3yJlo+mmNOY4YQ3mNoFtbPCLoM+l6+M+yvF/Eah9FInjAqV
3Sy5MehyvoOCa3QqKK1MjcXNosQ9YyuCYHXZq9Qd5CNYIgCTUyOZTNG8iY1WpXdx
Xj7uJGvv2TGZ5wp/qNaCBTyFIILyimQ4DnNgAGGlXi7bCBurtWJDwkj4e1Et0sZW
tGTDxdlHmr3Y+8GTPifcrpa4VO9NFsnL7ZX4nkOQE4cwSWAG2Rw5vOKEJG0z38H5
X8wMTOpEQnZXQuDcAoaFiGupmRC1vklVGd+tPbGNwkjVtWLaXeAq4tq4yS1vbhNP
HTTu/dMV3QvHUSp4NICwfLDm1amqQqkAZvfAGePHY9BJ/O1EBHk58F8hLo1aUzQx
59GeqSaqOWka+X04PdRi4b1lFyfY0YN+gp84U7jq3VheCeX8i9MgPb0xo7mdcEnz
i7ePDbqLU9AAPxJY1Lq31cn2dDyMJQiaX73xoGjfBZGFHaInYtqrSVeKG6ixmrri
MGgWgVLyd/4eROh+J43HUW0IVcgTnqYyvpkkq99F8vFauacDdebw6b8rnyLbyB8M
dZ3lKkirIEXL7+F7mnHUUpXM4s1v9ph+WebdbhsqbqbVJyUx9tomxAivoWURPB0y
hWup2fa1DnsvcpGZZclM2yTwVMf2ybu3hQgYveZt/H1Fq+p0G7JOGzeEPioZFvBX
fKasmnmrxO8IQLjKIAN5QALl/XWzyrUISp6WFsVgXAKQCKr9DNKx7tD0ZrE1TO8R
8vJEnTo6+A5wCDtUuso2l54XFs+m1Pc8UnF3w8kDTq5YPvaW5+16EkaoTxG8WVWD
W4coOVnnOXEgNbwT0R+RF6oXBZzM4DyJ6XwKe9e1XfVh7Ddhx51h+XvflOT3c6a9
YXlQaXzEbUsF2Sei3dksdg5RadOzKuwwnHEAKc4knWtEe4gsb6WK4yF78oag/xtZ
HJ/Y+maR+x9vfRPfNfhyReqt95+OzA82mt5hFBXB7xVytteGeOiwgmu3StyNXX4O
IwfEnqC7YIXUfWj3JsEn9kv23RCqOebcY1fh2YyrgQYBr07umOoO2nJiW9NULNbk
KnNLEiCpO+0rz8OrzNMdqK2rjcsLLtC+Eiw3l9QUEVr5fAFrwXEnmwpHkgQ2O/xD
ntr8/aEl/JO+ROxVlW9qSOLviFoepc+bZPHeQh2ye2gdlJWfVzEdhg1DKABuuVed
QH96UQ6k6fhViTYEHulfwsy+QV9bo5FD+uBYPyhono2+syp2aRrOeLRAjuw7LD1p
sJDEB8c+EkizFa9cy4ry4hAixm5+6WB/1uKKBGbXA7vSxr4t/HDYcIKuMWmgnOer
9PZo19W1fhqxxwAgPH3mZNEiF2vfHyMJg6WruMheXKxd6eImnI6NIQtBLZs/CYc4
tKJWTA9MvlZi+SwLmNguoRhdBsZJBBN7EBqX/OPyHvkiSQco5xnD04TBO7/RLqaI
+hl6UHKu4l9WlDzB3T2zyMSCfj4+28b4lATR6Uq3rNPbozYGXJBexiLuPS08XUsP
p/wj2dIADeROwdvGAyMvkIdyVb2BzUHYM6Jyhw/xKQOrEd6yEKGG61s4FA7oDwgS
wVBB3AfqUonnrrrLPtVzcPNDWYXF2bArcgUBQey3M2OpAZKFL/GwK5l28A1Euji0
+M4QnNqBt0EqrvvQbgR090NPTVgNSdn2hmGHbOA7JotVtbYbtl1z1aUP4PRtskcc
GDH0Gsw1Xh4bwVbRfTalpVOMPxTwiclbXTBjCsPy3j8hgx3aTDvKVzt98zTPD2Rr
eH4turJcGeOxkLeReL5PNWhr8QpybBZaxR86PBVHJzvXwNP3FC5nG6YUVUsBRjHc
ZzofY3g9k/7vPKWdoW5KadDPa+L6xPXQkOtiWqBZOy3Jvog+hhEDAGu9qVd1JWsj
OqmLPpa2O72ff94LzfJPEJ61JvPLN6EEmaDp064y0aC7LkAxA0F+mPi6cXijydzR
87E2TIFLUMp1dRPBRyGSIHG5j4ih0td+v/0cU/qkIcXbgZlQRITsTr9omCqpHAYG
4LbeL2bF4suOf2ojMGz1GiuCyUyImOM/8oJbXNWh3/uuo4rW/o7kvBf+6WBQQPAP
StrmcLnqVLkjJ++KlIasw/w7ZBX1yWoGxHNfvPM4R6jWrYiqFJLOSZ3unMfZn9Ub
E17LI4+VqgvLAj2/uB1JQx6+omikRIjqyTJrjQQm7vNXtf6v9twkMZ/lAi51cNwk
JgnYdt96RFIBUk5O99WrgAFuNC/h7SrwzfT/orekfUbRRCx2jB9DspNaSsIoHF/N
2ASu3ORRcxTtkkF5H/IIZTzr4RDwYPm5xZgTlNNBGJp2IlPE6ZeuISAwcL1ui0Bq
W1o996mZixX4qcEJSJ5SxxXDfcv/6WeZVjfCf77a4FdD8E0Wrw+UILGuOP35POvF
kVGeduZCd/X3oJYG4MUWTamwh0lAoTYg5JBqhQtfrC3B4b341TAvs7LMDnMfBNFs
txzu3IQEM8TKX5geZnSwU4HbCI0vDiB4/3ZD+FGiplpWSXFwOhXH8rVQwWVP1WM7
RZr28sHFAgtecZOdPAEjq5+QCCgm8HA2KkutIRetlqvO0lKX4vVAY4O7XREJv0TI
UGkJk5F2PJ0TSHJFA8CLoJiRmDZFEruOJ0dGhtqasLGeDn9dFm/K7kv944NDBrA+
VZDzC7is0YoxgQw5r6f8MOFpUhL5H7E8CXe3P0F9YtW7v8DpPnoyZoCQXaTNnB8a
R0ynomikZ+Dr+X/Zt1M+GyJ6+MLxS9Rgr/b5bO8x7RU2XQ0qqw3meefFDPuY6fyu
bOx74WrorAS2jDnQQWgAE98/2IeV5/z9ZT9wBgTsNMHxukU2Dk+dVPVA64hjoZEW
NGIybv7QTIhQnFtsRaqyMktBFa4AwLY5Zdn6ZuJl7iu/JXalin5IBpR/OVJ6Lwt2
74wF/X6ne6/X/KBne0Sxh5TNNNoQzHhP/sWq5ngo8MF3qHub7vUoUyOdbXkbSZ2m
xPkccvwmDe8sKHwynZjr99Irz1FurWTAmvu4FDSX9AA4adJ4tgUaqmmsjEkf26b4
gdOqoOiIuAuoZxg9xV8MWULRbCzNUqoKWIiQffcWMRmL0nArJ1hw3NBCUqSwddom
6qXtah2bUus3tO8xTckTBNxl2dUqKvlbKb2gIx6oAHKonWk3mSfueCzgB4lKM+rP
COt/ACAsfjV5vHhBWbyqW1FXqSSAjeijvcBvDZez3yUMOD4C+QxGtKb2fJ1vxTLH
4wg+1wdICDBvk/6DuEId46wcDCu+MgDDPj4g/EfKEhceFUzjsCArdZQLB/cc4ZXo
uygYDawPta+7l3YQUTLX7PJEE1Ef6kT+uexMh4XD17VjX8ecrtU2A2IkUDQbx9q2
Pqsr4klMQC9CbSSwJopYMIcXjqU0fibNgJqdWyE7dx1cMd6RMDoob4+DQ8LEMNEC
U2gXZ7Nf7ZQZ4SmD2evuUJRK1EtjSjMmnBlRkemnIBcXgsvOq3ODEWa2F7FCepN9
Y91/hUoh8mQcYPYnNJvmYp43WkJrsrm8hqav8IWdtb8sG/zwR5Kc0/cFR9Q1/2wI
J8KB/0oXTLkZqrfC0ONvIx48d3qeiTRbTkz4zX1qFpyvOf1PTYgnpl3yd8H3htuA
d2Tqw1VZCERgs+DeK6JQQU14w/h/lZjXVWzSy9H5y31n6YCS5LMCmVrOFsKH7MrB
QgRgjLJm/tJCyvLkuD4iVN330BuwKIhDDEKXXoNIWq+uMEsoBb5fGL/doDu2v+Ky
9MZVsGlNbPSZ06et1axXa9SsFElSckb7vBecr+Y/f/fmAYousjAK99j8irVG6mpR
HR4A86Rhj/9PaZAgucEw8Y/uPg5ur35JTssUJYxIQuBac+Cd1fzIxFBgCWrebxDf
5GVLjIPQqB3QH/FU31YbLhkuyWFNGki6QsmbL2q2fARrnqd8R3wWw1eSvi7DkIgX
8iNjLt0QKhKb0EF9imtdhoDzH5y3VPrEP4W5F95tOi3EtpMJM4+dubhT0Y2gx4Zh
zDtEWaXMupb6EOI9O0WZ0tVtggToMwrjLBxYA/NhDm/S3u+p8X8QqdX/FkyNCfQt
KcjNk8xQ/UzeNnhsPbNaXuxTnJ/OKfD7QUstY9aKFJ4zUkRKhKDiOeeHWei3x+OC
6xZ/9kjMKW8Hc/1e5Qw0HghCnKQiRd6KXPVcRdNAF/M1tD8qSlJDu1nB0nw+KeOF
CoUNChBzRP+sQpLaAq/X8CynjRlSgvwAmPbYYweSf/7K9lY9WTNwto7b/qKmu4EF
Ebw1dI4wjN28g908BvGi2JnQf4gAIewCkOecKw7EtFCiRj3zVLQt8FCjS/vWiHGk
/czpgbUwBXjbySnXRCRNGbPdq6TlY4D2oVCZ709JfTRzJC2WYOdOWgMABS31a94G
6QhNsIxL/2pIO6kMAo+Dwha1XhhlV+A0qiTZO4HzRSodvOx0AXKnsSKs5PvJN1XA
1PWS/caZKZgV47etqjKgH6u1l2l91GEo9fS1GFgbdwnpGEORA/qnyUJMV+z5jlTq
K16ynGZ+lMEzzguf0vbcbfwhopUJuSx5wZjfWRMr2S2v9p9YP/HhVJAdl0ABQwF3
TX1Q0gQ612KJNLcgFYoA2m2p/tHC5xz6tEqGYOoBR8PIAuop1lkak8WSHWLDEKoB
1Ep5Zeo1jFIJ0XxOWSKCb0hQqgDL14cB1fmbycoIjLUBEOFW4cVVyCIo8JX+Gehs
O4t0qJ6YgEC8Rn7IV9qs3BH1ouNjVwrPyK3pF4pb6lJ9F7PcqBqH05cm6w7Uscv6
MwLnmW60pEzNMYB9fCJxzLfA3zbN4E3qbhfRDc6U+byhxVU4rLwXHoQWuSovIX0q
O89lc5mprSsIGCYaLIAhB8C5iF+X9A7vsnLvAeyP0fDdxM7Z6oVaeu6kVz9N84Fm
62lFcFwL309LIaNZphfEjEn+w0M516lf4zVtJ/x2QJit8ohKQeMwBC14ZjOos6Ba
S+Y4Dpyj/kDkTGmpcER9K7bQ4qstSx4HyG69ngYDdezy/cFzDMrcD1Aswli7AVQO
kGs0kIPDdXDWKij4E9/HEmvLb3ZdYJlVL3BwiTMq7KhW/ws+P+He+FEQo6aOe8eB
liS9FKFxvxq9d0GjMa8KeQXaRCZvaj6bwFMJkjlLGY+EfpF8Gx7ECNYcrUunR78l
eJd+Y6fpnSjroqSUSIKD45Cv+Mdr0peiEXoGcnimDyp9l2yVCBlz96OtdQ7esQqD
CqDx+vn/OIjRfIiviSnArXr9PbMIq62r/7DWBBXNVVTKOZOvMyVQSr5Thrm+5BFH
gjgws/+RDuistWrV7753wM45CM0DhGckGZ3ftxUt2gwruw9I8As7fxLHdZoBgxd5
sc+BJjFaLtsRTvA3mqkF5BUTLKxhhy1yN5boBqiFk3/Rcyww97tHgq64qTytPn6Y
WFgcq0SNS/hnJs5+WcCnkTlwae34ze2rT4xiEj3wsifEogMGk5rsEAiDeMTEnvL0
T5o6/xMbsgxeeZmFVT7/7etQ5XAV3EwPD9QC5v/Nr/vaD8eVW45+sVJldLVpHsgr
mSCLrbJo4+dQVWkHny9JcROOCeugP5myNAs1QbbqGqeikrEdcjTvyZENQLp3HP50
QRVZU6J+SekIWlRPew7Qzyc/xSLRvzr4Rq4+kOl9HamDaYo4Ms6+sibQsc3kHB8h
z6bHxBX4T+W2dYkRAf5UU9i+ScTqtSHCTNOdrtNPYyNqiP5MaK6Y/hhKv4643u1j
xnd4oi8OEy1Ex2nEkXV6PtpNSAFWwUvikAd8s1nu1sAkd0pZLA+ZB7iOy+UIPslA
3QV8m2LamLnqH3AFrUIz9cDPZ17tQEszlbaXCSB+KZWm26BdffxGXwDuXeyqrYMN
3opvoHZOvahi1R/Of9nQo0HDPw9KGABBT4WEyZmbEzn/rwc4CJEQ6TwMs8KKmnux
7uddy8qohqVV7HsLYQCXi0ftaYAnPM14q7/r1eT8XeXAtNPuBUX6WXs0sZTkhzD0
C6hSdchbtRkgnRCqGCjrbTGSoHh3A730tNC55BcIJmn37QyMNtF19NvsFoatJTan
+TeKZR46UDkTVspK/MHxbCU4NcXR888VeBhuctQmPUrKP4fHbVnnI4J30GrJyEIY
JZqd2J+6I2IfarsJ3+QfeeEV5y8YNl6Ht6kRIcWljDgG7jOnePtYW5XP/a5goITn
XiZ3p+7h83pXRWK5IzZS/dvT8KxFcVK89SYV86dZJ8appaAHxRW6mlJX39LJ5Sfa
0sXiHDSpFn+rYY0/3wTU/fkwQ6ucrKmHGCw2YK3Lt8z6Jh+5Qfv4hRqDizXGGVkF
m+TebVUU8UhJNpRsAoot/hVJQfDsGeBl3XWMYs7DsXLcv/BS8hD+tuXyPh2S8n5r
4tbjIxuDqbX2ptoO39sISosLYl4PoV1oSriwee1fm9ULoUR1qrjnRuWlJABfrqAM
7TOzsyNKMWshFhKuyL39QL8DYIiDo++N5KclZeKApyfpXZU8sI7QaDbx2fClaTSj
TmRu2Kv1WrkrX4baDXjIrJrO9BMS4obcj55UE4msvULORmA54KmdJTlV/7Vi/wxM
1Z5sYVVJ2rv0EZVHqulmD2QGnUwR1sNP9hOS8nuhgeZZe04jJc2pxvcVIxX3Lwdl
fPZLZHDtBt+Dm3Rm2sR0eVoSyY2tG8y2p+R/YJhc1gnU3LGn1xUKG6JFKjNNYblX
YWJ5zJDQUJNFzFNbZDNsN9idFalIr9GLzjddlvAeBa0mQ4LulY6gEehp7rFjoRjd
lqtCUdBRDKeo3q0las0D2dW0EtaRP0Wt5mGO55BsnxKZjaWsDP6zAkxI2SIfrVJA
nwj3dhiu8kxb9Ea/+peFIaTyri5IGbUo2S78/xwG4O/gf5COo4yr+YbgF6vBzpgY
IsGaTaReHuBIMgK9hPTC7s8HqOfWi5wME/PGa/HoXe+xZ8k7kDlOX+wY7ii7UWYT
zycrD6KKQfN30ldlxBnP3b+JsgouHkuzvXJKw8+ZRXvZvMArYiTVuLNbbybjVP3A
pIzba/w0mEQ3uOhXdLedL1YrWRuN4fvUhbGlKm8fruai3FpohYBIKCaSrgYmmTeH
4JEY1aBx29Gqf4LPhIvrWQpCwnb0lma1M5tSKqbDdebklPMV/1V2KeoVbKSIPPne
/N9mZqugyAUnL0khR+ckOjEPkbBl69AQ+m9hB7YvhCuxFwzxS3Y0K6VShD0l+jMM
/VlFxPWubRdgjJAwXlX2vX0UQgK74FOsVZF9gjMsBg1uXhaOuclJMg9HPqJi8J0e
niGdEeG7+NQJ2QM9THY7aWE2C4esV4m8FfHjlSRveEXEF0nOO+nfv4kwF3ns7wfs
jULd1qo464sQajE7/lg/x2hScDjEKUceS3rwZP49Revxzm8n61dn36k9zoIAD6Yw
K12GR1PkoB8OR2JQDQqj4eV9Lbkut17vw2sR/YxeeUiCTHwKKApn2m6Gf8b5VL1k
V6O24xnowKqxMh2ax8UJG5VUek5TXn1XysCVlaPNxuXfi0F7lIyreOo1xAaU9BmT
XfVDgDSWuua4XExU5SUE+ZTt5b9MTn0sbgSubDbT7IhsS19mHCbeBMfrLVPtaDEB
FIcaPZCdT/DXlurmXYw3lqZ0unhYK/rc/yVubiBtmx73bKuZACV0uQRTPJNVNMnN
K4o0+FM1W1MgYv1HHH0gYnLwjmdcQUg3dA9iwgttwk9ENuQffz+xmJTdmcSObvYk
VgUouYieTs+6CXwZMfmvlrLq/HHHORQzBW69jJB/da5jm9PShDk6hPMAZvfLPpsC
UAohSHwIirBaD3xGbmrbAtM5pjJr0e2biSDEJzbPEgzNBkg2NHZGn8Rw22evDMF6
gkpsDVmfTxLg9M5r/n51dPoyKeGUeY02S5P29cMH8FFJdFcUHEOqeuDBLFLW0LUw
SPTFijb7r/GPmsL4J5z7gH9sf1RXs7pl1cvqa2xhY6NTxC+gR8dYRTErMFdJRL7E
D8YOcc3L0RYVzSrysWfZKFbbn72wbMFR9E0XzK6Eu2dsbUXhage5QR/Lc8M1akPV
88xBTApbU6OtrvFXEGYQ+C+Ns+ksSs1TMQwmyb/zXi9kO/nQBZp8KerLbJBCluhy
ABQX7HIXTv3XA7CbBpRm3VzRGvfZKZdBnWDWWhe4Z3M/maULX49HYuIe1qcWf1Dw
FSz+EL7fIDx5DLtsKJ0Vqwqydb+PrdWxpLzQ668qPLabz/o3YnnJRA8kAHNLmayX
UFfoPBgwucAtDd/can6TNO2u9rWgK6Az3Zh5njbi3w5BRiaq7MxECQnfgU/pTtbz
cxBUE2VAsUHCT2fR6mVCUQ==
`protect END_PROTECTED
