library verilog;
use verilog.vl_types.all;
entity MULT_GEN_V6_0_NON_SEQ is
    generic(
        BRAM_ADDR_WIDTH : integer := 8;
        C_A_TYPE        : integer := 0;
        C_A_WIDTH       : integer := 16;
        C_BAAT          : integer := 2;
        C_B_CONSTANT    : integer := 0;
        C_B_TYPE        : integer := 0;
        C_B_VALUE       : string  := "0000000000000001";
        C_B_WIDTH       : integer := 16;
        C_ENABLE_RLOCS  : integer := 1;
        C_HAS_ACLR      : integer := 0;
        C_HAS_A_SIGNED  : integer := 0;
        C_HAS_B         : integer := 1;
        C_HAS_CE        : integer := 0;
        C_HAS_LOADB     : integer := 0;
        C_HAS_LOAD_DONE : integer := 0;
        C_HAS_ND        : integer := 0;
        C_HAS_O         : integer := 0;
        C_HAS_Q         : integer := 1;
        C_HAS_RDY       : integer := 0;
        C_HAS_RFD       : integer := 0;
        C_HAS_SCLR      : integer := 0;
        C_HAS_SWAPB     : integer := 0;
        C_MEM_INIT_PREFIX: string  := "mem";
        C_MEM_TYPE      : integer := 0;
        C_MULT_TYPE     : integer := 0;
        C_OUTPUT_HOLD   : integer := 0;
        C_OUT_WIDTH     : integer := 16;
        C_PIPELINE      : integer := 0;
        C_PRE_DELAY     : integer := 0;
        C_REG_A_B_INPUTS: integer := 1;
        C_SQM_TYPE      : integer := 0;
        C_STACK_ADDERS  : integer := 0;
        C_STANDALONE    : integer := 0;
        C_SYNC_ENABLE   : integer := 0;
        C_USE_LUTS      : integer := 1;
        incA            : vl_notype;
        incB            : vl_notype;
        inc             : vl_notype;
        dec             : vl_notype;
        inc_a_width     : vl_notype;
        decrement       : vl_notype;
        a_ext_width_par : vl_notype;
        a_ext_width_seq : vl_notype;
        a_ext_width     : vl_notype;
        a_t_2           : vl_notype;
        a_w             : vl_notype;
        a_t             : vl_notype;
        b_w             : vl_notype;
        b_t             : vl_notype;
        mult18          : vl_notype;
        a_prods         : vl_notype;
        b_prods         : vl_notype;
        a_count         : vl_notype;
        b_count         : vl_notype;
        parm_numAdders  : vl_notype;
        ignore_nd       : vl_notype;
        true_ce         : vl_notype;
        mult18s         : vl_notype;
        rom_addr_width  : vl_notype;
        sig_addr_bits   : vl_notype;
        effective_op_width: vl_notype;
        a_input_width   : vl_notype;
        \mod\           : vl_notype;
        op_width        : vl_notype;
        a_width         : vl_notype;
        need_addsub     : vl_notype;
        ccm_numAdders_1 : vl_notype;
        need_0_minus_pp : vl_notype;
        ccm_numAdders   : vl_notype;
        ccm_init1       : vl_notype;
        ccm_init2       : vl_notype;
        ccm_init3       : vl_notype;
        ccm_init4       : vl_notype;
        ccm_initial_latency: vl_notype;
        numAdders       : vl_notype;
        log             : vl_notype;
        C_LATENCY_sub   : vl_notype;
        C_LATENCY       : vl_notype;
        c_pipe          : vl_notype;
        multWidth       : vl_notype;
        rfd_stages      : integer := 1;
        no_aclr         : vl_notype;
        ncelab_inta_high: vl_notype
    );
    port(
        A               : in     vl_logic_vector;
        B               : in     vl_logic_vector;
        CLK             : in     vl_logic;
        A_SIGNED        : in     vl_logic;
        CE              : in     vl_logic;
        ACLR            : in     vl_logic;
        SCLR            : in     vl_logic;
        LOADB           : in     vl_logic;
        LOAD_DONE       : out    vl_logic;
        SWAPB           : in     vl_logic;
        RFD             : out    vl_logic;
        ND              : in     vl_logic;
        RDY             : out    vl_logic;
        O               : out    vl_logic_vector;
        Q               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BRAM_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_A_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_A_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_BAAT : constant is 1;
    attribute mti_svvh_generic_type of C_B_CONSTANT : constant is 1;
    attribute mti_svvh_generic_type of C_B_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_B_VALUE : constant is 1;
    attribute mti_svvh_generic_type of C_B_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_ENABLE_RLOCS : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ACLR : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_A_SIGNED : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_B : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_CE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_LOADB : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_LOAD_DONE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ND : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_O : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_Q : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RDY : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RFD : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SCLR : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SWAPB : constant is 1;
    attribute mti_svvh_generic_type of C_MEM_INIT_PREFIX : constant is 1;
    attribute mti_svvh_generic_type of C_MEM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_MULT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_OUTPUT_HOLD : constant is 1;
    attribute mti_svvh_generic_type of C_OUT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_PIPELINE : constant is 1;
    attribute mti_svvh_generic_type of C_PRE_DELAY : constant is 1;
    attribute mti_svvh_generic_type of C_REG_A_B_INPUTS : constant is 1;
    attribute mti_svvh_generic_type of C_SQM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_STACK_ADDERS : constant is 1;
    attribute mti_svvh_generic_type of C_STANDALONE : constant is 1;
    attribute mti_svvh_generic_type of C_SYNC_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of C_USE_LUTS : constant is 1;
    attribute mti_svvh_generic_type of incA : constant is 3;
    attribute mti_svvh_generic_type of incB : constant is 3;
    attribute mti_svvh_generic_type of inc : constant is 3;
    attribute mti_svvh_generic_type of dec : constant is 3;
    attribute mti_svvh_generic_type of inc_a_width : constant is 3;
    attribute mti_svvh_generic_type of decrement : constant is 3;
    attribute mti_svvh_generic_type of a_ext_width_par : constant is 3;
    attribute mti_svvh_generic_type of a_ext_width_seq : constant is 3;
    attribute mti_svvh_generic_type of a_ext_width : constant is 3;
    attribute mti_svvh_generic_type of a_t_2 : constant is 3;
    attribute mti_svvh_generic_type of a_w : constant is 3;
    attribute mti_svvh_generic_type of a_t : constant is 3;
    attribute mti_svvh_generic_type of b_w : constant is 3;
    attribute mti_svvh_generic_type of b_t : constant is 3;
    attribute mti_svvh_generic_type of mult18 : constant is 3;
    attribute mti_svvh_generic_type of a_prods : constant is 3;
    attribute mti_svvh_generic_type of b_prods : constant is 3;
    attribute mti_svvh_generic_type of a_count : constant is 3;
    attribute mti_svvh_generic_type of b_count : constant is 3;
    attribute mti_svvh_generic_type of parm_numAdders : constant is 3;
    attribute mti_svvh_generic_type of ignore_nd : constant is 3;
    attribute mti_svvh_generic_type of true_ce : constant is 3;
    attribute mti_svvh_generic_type of mult18s : constant is 3;
    attribute mti_svvh_generic_type of rom_addr_width : constant is 3;
    attribute mti_svvh_generic_type of sig_addr_bits : constant is 3;
    attribute mti_svvh_generic_type of effective_op_width : constant is 3;
    attribute mti_svvh_generic_type of a_input_width : constant is 3;
    attribute mti_svvh_generic_type of \mod\ : constant is 3;
    attribute mti_svvh_generic_type of op_width : constant is 3;
    attribute mti_svvh_generic_type of a_width : constant is 3;
    attribute mti_svvh_generic_type of need_addsub : constant is 3;
    attribute mti_svvh_generic_type of ccm_numAdders_1 : constant is 3;
    attribute mti_svvh_generic_type of need_0_minus_pp : constant is 3;
    attribute mti_svvh_generic_type of ccm_numAdders : constant is 3;
    attribute mti_svvh_generic_type of ccm_init1 : constant is 3;
    attribute mti_svvh_generic_type of ccm_init2 : constant is 3;
    attribute mti_svvh_generic_type of ccm_init3 : constant is 3;
    attribute mti_svvh_generic_type of ccm_init4 : constant is 3;
    attribute mti_svvh_generic_type of ccm_initial_latency : constant is 3;
    attribute mti_svvh_generic_type of numAdders : constant is 3;
    attribute mti_svvh_generic_type of log : constant is 3;
    attribute mti_svvh_generic_type of C_LATENCY_sub : constant is 3;
    attribute mti_svvh_generic_type of C_LATENCY : constant is 3;
    attribute mti_svvh_generic_type of c_pipe : constant is 3;
    attribute mti_svvh_generic_type of multWidth : constant is 3;
    attribute mti_svvh_generic_type of rfd_stages : constant is 1;
    attribute mti_svvh_generic_type of no_aclr : constant is 3;
    attribute mti_svvh_generic_type of ncelab_inta_high : constant is 3;
end MULT_GEN_V6_0_NON_SEQ;
