`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W0h9xobeMYpzFiZf3SpV1FncnhJ7tNa2Aj3ucv1XQqV1JIH1Z9lLeVFOgilDSMJf
//xXJVptFyiNtsbjtNkFOmwneOWBbTAHh3aXtFLSjw3ieGkqTZixbkGj/+0m/7TF
atvV5kWmXig8Eoto89DRTCBapzW4PxVe5ujOKj38eTx8oxbUMK7mnvwUWEjKPCFr
C5C7A+DhDcUDcItRHsJYgGW+vDiEsDvZDncbmOKs1l85sWq7ZA3w/dvdLjSO6iZP
09PuN2yBaCVcdvM1mvK0nroCdeeGOKBG8BXAqSu1n/ZIXPNn7d3/ysRYiDQ1yqXn
noiNvWh+mckEeRAazxCGKqYly6kZeev3t7H4ESAUa8bHpdpODn+TSsPLM2xRtDtX
7OZnLqhUXoEuAyYD3ZilpyRIJ/4w7Ut5lw15UICOgwoEJcxKMVFpWQlP2gTyrZXi
EfEMtrtj0nHm1ao0ANxlQiNlj+s39pk0aNrkG1KoU3GATLXn/OLzaAh/cnF+Dv1+
x0wURKbina9icj5ioJYgjYqxpe/uNm0LxeZiulzDI0YZ/piZ5H8lMRi55yBxYK01
MxExYAXqKAn2dVZeM65PWw==
`protect END_PROTECTED
