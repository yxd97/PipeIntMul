`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIE9bEWMPvc3PK9SIE2WPEk82D7V6zIHyvKn3hu2Zdll5eBYODEiLY2BVP+gyn2W
kclRiHLqHrLU0+nM7yZKYeVBHE6CLb6pfhD175UmhtcMf4pei46KO2ZYydC+u56+
zGb8mKalJJg5J06ljqKUxrJ3HShNp0NltbvftKodXIjCKx1lQKdQc9ngU67TThXp
x/oTWZ82PqyhR0fB+LcQGGjvqzvuXMd6MYmYBVtZr4Z9FLl/396SHXCWJXLYl99E
vDsaij4zbGRg2nbjcvVQsiQJyXbecEbowAJ0TWdR5RoqXD/xbWpiHXXKqXj1M4GC
6TGfsAnRjAAyZdzQM53xFBuIZ8Z02hY6k9XajQEJKQncX4gQbK+OaRaIzh1WPVT4
YewwtspHOyUCoWFgo5xfBt3xO/6tfnRomDflql5i1OZlkhVaQiN5ajtTAyzgABw7
OplaRg+ZFP8PlMCptOoAaNiDzDxarNFkXz4nR/9HfJYUl+p+HKIj6W2OaTcdlZT4
8McE7GBOzcTlJkAmwe/MOI5eR1ykfKrgiMdlUa0wfns7TpdNx2HWDvuXOeIxMPzM
OD9Jvqwax4O6nWp6+AYuTNXmL9MARaXkswTzsgrKrZ9G95glijsNyKTHHOOLcDQc
p663675XYWES5dTKeLdlo0ui4JFBgdivx+k2FooYNqh1A95vjHS9xP6R+vxK+522
xmgowu4v7I9HL7TXmBpXc9qKRM/kbMdYq/6a8kHz3VS07d98PUlOYpK0Xa7Uab70
/eatMpNbhrupWsPRuNGvuicalynmb2LO1DW69KjREaqE7InWGt/YEKDFeKUTXacO
8vd5gcnMVDjwC4SNl3a001PYJ0XE/4Hz3DKd8x9OECnL3x0ZD94JtOArzIPdnRMT
WKXveM3U2Qd9cCIv/ZCr1Rs1e1HztK3lZXY/ED9FOkja5m0Mg1EMmIUmJUYPcikD
72GXcDD7BlCS6fEgc0uYB3k3xpz5wy3t2H1YmqqgJBXxSQSIQwRz+v1TJ8D2rnAO
`protect END_PROTECTED
