`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4YcbT4J5aP5htFQ5RyI27WDQoNXDSnR2TGfFMzvZSxJ10qoHcPnBz1EHiWx/vbry
hqRGU9eP5KtUStU5L8nxB4VfknpwirKkLhGypL32MIi9xR0KJ+e5U6RH4hpeSjR3
Xd0aq4J2RGS2PIy3ZTUPLkM5AreT1VviGjRtzQhP9Rv6ZQE7dzt9WC9rXwqdNudr
djffT/ANmmuz7A6wiSKmZMeHYrita18mkxt1U4t6ZI4tHDRGPC8ly7izB20j5uX3
jyTAzZvBCDiv+lEMiD5L1/eYJ00GJCQz/981vYnCktVQ5K5hWkOQSS3ezy2jjcEQ
h4xI8qJNq52e4uaqALKGfg==
`protect END_PROTECTED
