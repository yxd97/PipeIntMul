`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2izcP4ZHWJEW8u8smZ1yKi+QAOZHA5am0MvAot127E0s7dwzXWwvGQ6Cxv1j8wx
xQ3FpDg9Z1KJctokiORPS4FcoYjpUgXSnOJpiZQkhHKQqpalqulKKiSid5CMtgjj
KszAHYGm3nMkmnYv5gCKbMIbg8Gfvfd5qj1LWIrlDqP847BHHJQ/yM/BWs9TXjbm
taJwsIh7D0VKK4zHP2/7+QuTFsWOrjtwxixMDvXT/gGNZx/uHjq5e05Rz0wiJLPu
xCLdBGCR2L0YaeqCkiJweeZ5fL7BJghzoRO6BaJQf9Ve8i0lgfv53QmC/i/EdM5G
LQkwkJoO0zs6I53SRL2dx0fKHklGebXBddd/KIhBfFDzw0af6TKoH3dbFS8VtKoR
FlPLsEBChWBIWDCvSZ2q0k1rjpbmwM2RHeVP2N/BGhSGVEZ6SE48FeddYsE5OfuR
DbOB2p4VLAswU1Od2z5flYtP82I+c5Dyt5GvROo1xJG4ADG7vf1zGc1mRZ8HRDsj
SpbZtnxRedZL//T+4hnKVCRdVfLTd4nHqx6Ymqura6m7G+hqD0li+V0p+AVk/Dap
zw3VGJ8MSE/Khv3myj1ZruyMM95ZFeY081dqtE8QdQQ9g4JstEcmFg6Msol/h8/D
pg2taEVmky1lic5aXuInpsMQ8oD7cFWrf0qhXgS2nDs+gIr7Px73fJnTxBxsu0NR
mxTqoEKR1z/pXUIE3tX3Yk2O/DxTNlvjwQ7GXoFVlSWqZ1PCsC9wNPcY8nziKQ6H
0bz7dlSECt1Tfzc9ZZ5MqEAhAwOuMdhM03pv+hiOhnyBdAOh/KnwLU76YuPZ+ZXG
loqZAKBI0KBluQB6RUygOm4ybTluvpGxgi6HGfbgfTwcYV54oKWlGQWG/aoLtIn7
uFKU2dv9qdjtMgXsAjJnr8dykOVG/M218lImaql1uz4gBBmKWP3R3F7c1w5UiKyI
3g759hOFTTymnY3hrYtK1SkWkxKWg1fhV8xjfkkn6qdfl1tvx4Y5zbe+F/Qt8dcO
amSAtqAaW5MvhJu5pFn97ifuWYffTcqYIZs4XCvbqFbi+JOYXPz6B7lqUS7VERvv
5eKSwvYu+Xn9MMhXkAfDBKKEHD5BEpNTLUobGUsCUYUHmYaY0pwAa/i7TcQ815Nk
iWEjr1gOpxfe9wtCT1mTEw3FIwS/5wo84Oag64UowwE+mx1gJXyLLvh9C3kO2htl
aDruEMa5t2HqM4trNgdLrqvGMwHtuwO6rRtkawHShI8Rb/n3dImQmCXKU9xi/aKq
7PBHp9UXA2kmkhDL1459RoVqgYmyCv7ECjVq//Eu24GOrmquYwiCAB16fJvewnX8
9EeTenHpLf0UeuUaA7ZPTLDuuhSNMW6791WBI0gBQz9eDDX7+y9fpSUOK+ITJb/Q
0HOtm5OIcSqWc8EHR6tKFcoUSzOJCyvXC8m3v+0LuCnHKqpLlfv8SkPvHXcem8MW
Qrnonk0uGkFfqPxtgEumIti0GAy3qtqHP/g83lkCxGUfL8Zvzw5q5lstmgq+KjvK
5cI35OMANF2qMn4hQ2OhjYQr04DcXvUYZjwES8IFiY7JQPp0OIhfAVFU66igCMtX
+C+8AQZFGI746/5AYdhkzg1w+uHYPJ0LhGkNzY//iWX0cau9D752EC4nXaud0KE2
qUFQFvD90Or3zP89hK/zUh85Eo87pl3i2tALI+9CachNcD4iCTmHaFn322AqZLlC
`protect END_PROTECTED
