`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlcVDG338nMGe3cYB+wxwaeq4OjMlu1bWvUDSMrc+MqBW5GW7syRi3q+8Ej3f3Gs
kcSpdKhs0f48ccTaBmm7l83T5UQSPzHgTty9hy5k0vaIXD/J6cWNjxE55RE0x7P3
zAUe/2tTSmEbFcj3hZYb303YS0Ms+iKs2gen2mgJ4xGgYxaNivX3qRhskCwbKTV+
lVLSV3maYNi6Aig17wo8jAWoRQyYkudHgnZilo5jMKTE9ej+4zLiRibtDNMMctKV
92D2ooJfrTawKMQaweyKRXulh+tK7YBh7AC3ZJkt7wDtMKRjzeG2ir8DsthQwjXt
dxdYFBtYjDC98KYwNGjQyDu4Us2oWh312lYw/bcMMaF66CInkCcwtmc2osJ1suHh
qVOb4bmW1O9oLHJqKbO+Of3ONcX4wUoucwrvwzZuWfOWkC74exljB7+U0UCLM0mR
7uWwLK9YY/7MtmfYl29ja/J74qXPAjM9Z8845Nw0ZzPTU8JykwfVg2ansa7PweA4
tDTAsGMIJtZW3o/iGvmiE6Bhdzuu+1sAs737h/blAeXj2+9p3Cm+WLG35Xdg/0r/
l6SqxCkeFKfkB9giX+MpsQh2yJ88J+e58+jG8YW7C5S/7HRdgjF5dO1sgWvziV32
NiKbqQejYwJKsxT181cIwkkm/rIK+gDZkTocsGtX4t50Txv6+CqwNbO1vriRPfPa
X+jR9MEyt2RI7FBC1ob8TeVXqLlAboRazAPWuDWof681I2bnZbROYFhT3u6AR4Qr
BY69SGaKsz3Jv7oHcqHAvyj1K6tpVrTDO7ugyVW6QYMptmjGn48ucMlbyXW8ECe8
0tEFdqKN0oyvODzSokCyMhVsP1YbKkv9Uh+1M58zR+foNo1Yfa0im48mE9fXxHRm
eJbEMrDyIYGKWe9Alb52Aw==
`protect END_PROTECTED
