`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7V/hvuY2733zCs26XwCmdxMAPRK1WGhwTCMHaUtEzGZ2pDxQqIWLyeIYnxcsSwy
aD3kdzDPG/46GUEJT/sS6Ypk8XP8+KlhhyIiPPiYmCc2rfGiNBQ9qBvg8gIIwn2e
F+9bi6AtLRz1PIlmcX292kKV9ZKs4RW3YafpUv4kF/FWpYuznd8GGcbZSVuT1a77
yxIpDlZOrqwsVTIaCoPSmIREmdFdYZZQKGMbD4CKJkOvzom/drR8flXLZRXN561g
7wJzZaQ8renTppjauOF6x4hxWoMVfE31OlTb6mnsgDKaHZL6MBxwoVx/84wYZQmH
79FPj75rtG66SQdXlkq7e1P7f8cIZsAwY5NN9tNaExV3JjHIM2i6oQlnN1OIPuYi
aUzeVd+9XUejXHg7lVOR7SNreC9oi9BZCy9fu6K6IV4=
`protect END_PROTECTED
