`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kEqEcr2AbPYsIoASkfsohDlHQ+imcy0nMhQ5jg9yup6jZGmx4Glh/fpuh2xcBjXt
PH5IKIKjn6ia+usnPlmZvAcXQ32jVo04LYFWa+sJPg/SRnXRia8AXP2ZmRXgyHk0
8CEnbfSW47XbgbNPQisGOnUuioguJ8NvZEiU7oj1T7RbRGtFYp3NX0evjc+mWaN9
r/bR7rfFZWRrGbGWkxrmMdVXGeF0So7QxwlzM8Sdfw09yAi/hXBoRRpah6qo3+t0
txyYSs8mSjXd6nIFmW8FI8C2oRaS9usDWRV77wUdhmcUUSapBbMtjlwKmtklxJDB
+XU4yX+sA4VOPTaU1nRX95ZneJfrIieKEcjqF/KUCa1X6IDsJytUipnDtcTvMsQh
sQ7HNGYVxV6oAuec49ndZudWipn2Pf8k4g08AuTze8bpuaQGxw1BWsxIE8NFIZ0J
20v2Fg8ksfm2jSiYqTVjw7o25hLugMbsifJK+G3Pfug=
`protect END_PROTECTED
