`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6beb1gC7Vx668kNaq/9wrZYF7W75A0gIxnan0JihFjhtCSC5JBNJZLddOFUkNb9
lTy8OQBDjGdL6qIOcjWVWHUbFe8RXZNWPTzap0rIfsLlJOK/5hvqIq2l6XUEQBfc
37rNU0GHmklSZVqc1/iFO1f8IlrOs8Qr3vtvLbDdms/v8G0mSbc8bQyWByG1hA9h
btAgpia5iOmCplVuFes2OVJ763lhKqvHYqz1dkWHNEVQR+eGI5AuWJivDvj9uOEb
kYeA0hZtflBd1ysFqSlKxgErhniJqr9CgIaPuqxC7L16gECUfbI/2BlBiiTh2Tmx
TtA9hhLney1/SfQP1alN12GktgauIygtTuej9IEH8zUddlMqGJhd5+yrKMpnn5VG
jIxd8mbmoQLv8wXT5NCnrgEueRITjkTveel9WbisZ9CdhPMi0tNaxHKsO2Ruvdro
u0dLPp0rLZ0nzQt8C5XCuY/2I9q+phvh85zgNqz4ohekrVy8a8Nz+L5UBbPWnai0
vBf0QSP8/folvHYWlKNt4NUO5vo4XV4ijLdF5KgWMdMx+35F9o/kptHl3ouWoICs
I8lpd1OEt9e/QitFXa9/ERqu/ze1FMjzfKkcwUkkkf8=
`protect END_PROTECTED
