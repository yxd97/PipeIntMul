`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZUzjedHjsjlpBdS5bylG40EVCG1GnxQ32aZ8yVJLTJaTTNWWyaVHoUiiZZcUama
gpgQRnWwnO1A1UR/t+N92ZQrd1Z+sOJgaa08Cdowtt9soQWh4nmSq9y49q5nL7I+
Tve1gQrcz9qKWZLODRiGK1JmBe+ufUrlMFwyattu2OcfSkjIByGQUlh7enWIT9+m
TvtTRjlU9sjTB1nHSUr3KO+2rVaWb9xH3kKFrS2doyuzEKkd76MlAEJ3w8OgL3x3
fIh0nRhj/oZF/A7C0bGZ5hmwN9FXWm1Z53cMYwgyOYvcIPJEqyf2BqmEfM/TXmij
CbgWkePdnKZiarSaW8LdzgoMEj48CBItumU3IwPDcF2NZNS6jNEU/7OSbleqEDZm
W21lqYjkWuHJsje4Vd0gM7Yyux/ED+bduqXEEV57QD4ObvA/UDua5eLUq5hr7jWz
1Js+lulBjEKaBT1LI83/4LG8xjHQ4+7mUvsgCRvSMDqU0uxruTmXQZWkNoyEVnYw
yDyWm+EyMyHQAU6jd47YBKPz94V3LZn/3CkZGbduz2mYiO/8584OgfrGwE2dHMPs
8gBX48FjV2rRyTKbMXhgXEHLFWR/1a7+07agcmPzbSxLs0taYxfIjstBR9MMifW8
W5ZDStZZ3r+J9Vw+8tOZ71kNoIlcNl+3vRkUkiAUknquv+7UM36UPFb4l1SXu1ui
QxuUA8t7ZrALBofOiafic6+vjVCczCY6+a3TSHasE7zl4TqufwJg+Ov8H2l1EmEQ
krcQEFHTf2SQJMeEMQpErukXvUHS06aI2Cx250AH2vYPbr7WweE1gLQv6o4JzwsW
/lDcpT9aqs5uNVmd3p0suw==
`protect END_PROTECTED
