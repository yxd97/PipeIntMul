`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YYunqVHlEK4UBf8iKBd+UNky1VQfxWLicSfORTVcdhdI2awEkaGnD5eqU+Nst/jC
UXHJzWOBS44XaTEcwLQSYPRzCFvrlkZTEa2nSU67kFml8TifUCODv0AdlDXAB67n
X46ttp7WJrCghOxGTJonIOT/UCEpExS/04lzDYxGL1Xty41x2R7kwadukm6n0R48
XxvFBeawk1QO7vZAj7F3p6BAgHJi7B1O8MtMM3Bb5IAcgjOlLbb2KUbOVxJjDi95
dxzgvuCxth1Br7GpHXLfNK9qvLddL7Uh3evBbDS8mrMYZeDMk7lnZ/nU/cXvKeT7
00y/lO25hqDBU/Ea0DryZKpkiHKELn35BZLN2jmI55dR+hwPtVqtzVOdezzWLaE2
PaKzx7Ag9lQvqotpCEjjl9J/OiHwcli21UVJGEGrQVfAF70Dutli2iuBXs5Tgn8K
mCqmSFkL8xJz4Wpt9c19sEHlrQ3JXBQD21fZ1UjMfiqB+WiAithcTD8Iid0rhcqT
`protect END_PROTECTED
