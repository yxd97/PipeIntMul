`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JM3Nhg5/FYM2JpTXiQ7byZW08j+Kb2jXHnJVB7hUQR8Y+tkPkrQm6dxMFl2yFlCw
0CI4cH2LR9/RVyw0OrgF2CMo9sZMOlrnghMuhtkwvCxCV+Hoicb8NLj8AdK8+EFP
XBI6k9xVV8g4BzJ1Zl3Th0fVHMBPl+QFhZNoN4pI0ElbcDZfwmKWPFEuuvWQETLl
EqqJ9P0kxG/sB52XO+9eb28XNfF8mjI0R3I3IVvwgp8/o4nib/gSCsVJINaOt04j
tcKTqo5BvVF4z2X0E5XD+bAbmQ+n9DRmzYvgyURzUWof87NAz03PS49kjXxGe9X2
JB5HK8H/NnqZ/8DA1yDzpYUnejX0JsYcIB93JvSJfO6YmUZm3HEXEKebqwCTjdZN
hZIe3A5tpPsG+FCgNmJ19YnNutHPjHa0j6JjtAc9usp8QFEGIlZnAUFYee949qAj
jQWjk9u1SMRM7qT8Y5rkyusdXQeYEtYOPES4Bzr/WG4I02og9FMJJI+rJBSYsVuQ
jvYeseDnG/r8IL5/jZcOOWpt41rLZthcfBjC0w7dPC1EBtMafjH4KmWyunGIneBG
XV8oLDVpiiYX2ua6taCIRsWrJtcE2YSCAKXb10HfvD1/QO+bIkZSLYcgs7haSkcv
739qFkiCpp6FZs3fMzNRtdFaQswOa3WpvuPVz1dLO0rLJhFoys+YQaneHGjOQygh
GQ5AY8hAqxng4YsdW5CpGGvmdoDEivk2IqSxKQa0pft0oYSkfN2NEXjnZjFN1HSb
3KoQVzB9CHmesOKvhwrG5X8UoIlMLcwowPO6HF6eJEgDu6uVBIAPrqq1o9yvJI2g
d/XBJvl45nSR7zz1mKX80D05IRN0sJPy/lBhsTpexUvPkqw2HpNElkFwDeyRNP01
7b+7Fu+1a4km7qT73KCMqp/bjCijVojI+/qqxZaMLPZjyDKogyFatt68iUiEovQP
KRZZs63daImvV3T55+HV3yXNkJekVM7rdJ3QBHEq4zW04O/U6+swGiaw+S1SJKQV
4zlnQ89/ChFz+vk7608GnXuCR1sqLjkVOToWW/9KquKdfpMGGtwHQFUhG0MOsss0
NT3l5D+myrCYTJv9ZSfa8To9ayw/jQEv9pPkiB1wq4k/6sTMhj3eqWYFqnR81oav
rRyL4h0GXPHcMaZ/pJ5q1uZgM15y/tG1EGMWFknKqBXB/CPzY/NdGtcpQSOPqRKs
Bweg2eLDVTQFx/dw79VU5sc5fDmlcgjTAHLm7v+qMpxxnzhE5vhrK1ejPOomSdyh
hob+ydaXsKZanFRgb1tyhbDBXVnzZei8bJW8MVZ49Wgn1jYMjvT6BCLCA3F5liCk
ELn+rSpc6fQcYOEszrTqB0otVUW+WLr6e1OVi+GqtwM=
`protect END_PROTECTED
