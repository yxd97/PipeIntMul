`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltAPbOVKHdVunmbjGqwBD2y8P8OwbiGflZ0zSXmRU0lfXNAbPjuBWNIKsqJJDEUm
5IEfhlRwbWJaA8/wHE3N1HNdstQxwRU48zQDONyQQdwedrVYmz+JjZSrZIQHtndX
sgNOEfKgCbx6wRYyDBvY74nzMXa2nD1Nisi7Rv4EtP75cgL8hHKFHdoG8o7cVzXx
pmayGnA+NvS0jY+W7AhsGA1gwkQDNf15QGu9dSv92V4zqxRLjKcQ1aAgLVYigJXS
A+f70hQgUKNQKIwpxrMnUufJqjw94yJ8Ub12lJTPqBx6YjofG/PYEznT2XMpuSWr
clQvZhlKA4cI5Y1XwwD7ZLT5XMDu9//Bmbbrp3PmJ0VMIaf7YJvzQ0+T9XSfgBZC
uNuCTujVw3n684FjF8MMlM8QsWsJmP7tRrc5XpX9UbhoS9BJ/x+9mjj6sPkMgU4j
`protect END_PROTECTED
