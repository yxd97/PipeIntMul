`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j1aSly54havH8OeDB7bNw1rQHgGdn9hkk/tt08WE7Hu9kODBLLKHBFAvYwCSpwCl
VkcsfdnVUA9QOgcwnIyEePXtKqZespIM6E5nHTZrYlyjcfLhFLb1B01PINotAY1C
w/n152HIlbH26XDspDLsDUYslW9mpiHdytWS/W+MR4MVAJPyIdu0rClrUugymyM3
ljER8wt7AQCoUp/vDhBc30Sqf/WlNqRhngtGY/y1auNPgEY3xfoBgds5VanyBODp
ZUnoudrKKtjpnAzT73X7zZ9uPuM16CxRVx3Dg5diBr9teesizM2SiYo+dnlMMwOy
31RiIo4FouIFYMUo5PeDffQehBnQkzdbhf8Xey2elGtNceXlaHPDYqdDkEoIoPM0
/lpycigCyEAiPd0fyYrt9jRGtiOS3DkX/7cj+1ulfBB3aXz5nr+om8giKqXgn9fE
xYz7PIs5k0wOf/vsnYRjo6+6O0f3N43ll4IKtdwgh/Ciw4vZuTHC/ofgAerjdBNa
t8wcDCPx0SHvUTNanwMADhGlG8aoWk7ZHiRTKtLUT6IhqKON6kjE1y0H8B8mPnKJ
W1WJWAQR0zBmCVoeafRTJw==
`protect END_PROTECTED
