`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IImxP9YKiIsgdHdvwXDXfMBZdSeE1L6oqNyxc8rpdhtCra0gjFOpywUSEwprZU0G
F3k/kaSLXVTEorbiVNZXLM7DmGrQURPbgWW1BQlGLE5JS+y5DiKPVX5MuGpwhBI+
UVeRyDHev2ikfGzpG0IIqu0TV7+w5bmp9lqRDdW06dnhJMdnu5IXnlDfRjrasNOJ
+mGU9yB5+t8jHgGbpDpOGkIzKmWoAeXBMTDKJLoboC7l4OPKeG2vVaxZqyA5QAfo
7MM4U6AsiHVsv1C522xdh0AyDv3iO2nPBxaFolBHtINHuLHKfIUKwYKjsJnyOdxE
0rPM5Z535qT5faCWZHTvDB4SmtnFYF9uKtG3OaZpU/YByKruV2gj135YQ9gtHGZN
unMB+TWjcDP4lkYXYlO2t9E7CDsewE2NdNU5Hu/sMuHbt93C4liPZSsNaYKdeMBq
kFt9eWy4njM0GjzSp3bGUg==
`protect END_PROTECTED
