`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/C00DroqVXBXYM4z2oNIeQj/nctBOBIezV5APF9pBblw0xJQ40rv9m7aJoN0iLCE
C2Jyp1qHzDEX6VfbBg8sPBtT0Fs3dk51ANhLu4DD7leLOpw6aXQSqNbW9LBgiSji
TiHQhxJeJ0sDXV72h5a1Y+NdJWM+pxrC+y4u07zYppU2VCQXAImP4bZgNCYQ1MVq
KdGd2dcqQxbud7O+UnpqJFKJ+p/6n7xPUJum7EDOJwBzAzB4145Pn5dNnhtTIhbi
MDiZY8GnVF5vqIkLnwPeEu4E3wEGruXbyYQWSRHi0XP9aGA4G7HMQBWQvxGqhCGX
UF9tGr5d+Xwo0azqzyNY2FMHyltCtId2C4Z4NycWkh/H6Ypnf/GBoPbvilvTNO//
XPN4K5mQe/Mvn8Fjtk+iiBRFykfPqL3R3Jeps0FeSzV3QvF/jOLzVf5dtYn3YO3H
unZ6fN5xQ4f+C+oROE4lRtc4FqyLrLFEkRbqi8i/uxK+LZCqfhsWVvmeDREcmavX
ps+8CqrfbAjv4GKuVCB4fEKOuAt426GLKkZ4I5FAecJ3SBG0Bid4Sxmt6IHUr+p5
INv10kDYPomgJHNm0ZqJyhxRUPL+Y/HzvkONY0KQ7E5EbY8qfKgqTD1IYH6OsFuK
KWdHV3xA3MwTcwDaqaXXKbaS6AovkkZAPS/buwQI49+rx1U6eCJLccLjsnViRfM+
d3aY9Esy7ltuZeO8JMRfs4hITAojG5ioGVfD2BwuxCNwtwxlElaPFjS40e7Coyzw
NuHFWmhysnFed6uAcqjEELYIAbUST4IDffPeI/5ZctxZHiYuogDKhC3EwLnovVny
xmYWmxXTytKYMnMiSW8Oe+OEOih09J9E2vYWG6Jz6XliJtskk3kEcI8DaOpex8/1
Dg3aInruxzlLkRnV2FmFO5g5oZbiolcFrFdlsIIY9Qs/YzOI4b5TRnNHVWMx7Cvr
k6YYOy5FyLXjjdNpK8OvqOpuqteUdnND8+zSstH5K3UbLaSA3kDgZXsoRnojxzkW
csrSlZoI2finRn4ccLylJp/0EPha8ZOYx/nqbQlikACwxDX9s8UBnkJl/aq9NKGo
qJksB/YpNmCyDDeeDvkcPKKABeFvMCOg1h+6TfzwVjQQbDeqQxP512KNO8JV324H
rZcoRdmp2qXXmZ+fpyvDUG136StH+0mNN0t1yaISumC++F+iBLkCq+rddhtC+Kty
F7ZwRpAIu/MaZSxK2bnsEbSO5lPVj4Pp0rHFJA3ZJxhoTpWANUvaf7qKppUEdjt9
2j60ieTysp4LEJFH8D4VnLMpshFxmzoRkeI/4cDMfihAFoY+FQUuBkfX2lrvZI34
GHW0VQ9/USLMPHAkx8WcZ3Njoteo/BcG77V+AyOvCPzoRUhG0nKWuzXPnneHmKrn
U4DLYYy8zBlDU+KIoqGL9UCLoen873ALeE9tLO6O5SXQFWoVjK3BL3VEQHvWWjtf
0tmhFpxGJwua4eXR2DYgvBDgoAcfD2CAFYBIQ5/erLSwXNeII4u/iyGeCQ3qfxH1
kBL2vfHCxIa8t6PnR1m8XoDinFpNeyETKGOo8jGo5cggzThLQtFO0XN/Q6aWH8uF
xsAwyxrs+UoMMxOHgL5UCcpQBWu7l0xBAyvcNGuF4/7HSmTGhJ2SZW28Rj2VInHE
EIuVoK4YGnLxv6kkxTJVFk/z99O1XknnvY/QlyqoBDTSzWh/CI8ADUC2Kk3X++oJ
asr8SbAahKt51efNnLT/AJ/FMAxywxHFobYT01h+pMadEj4YB8/gToj5RVTNaH20
lKnlNDqCZYxWe8DifsMXkqC0/QdkrooScF/vKYRiFPrKkNyD26YXwzO4JIC0V/Cv
iq4WU1xyLvvqlswmg8E/4o9udzD++i2WYonXYXW3KBUoh8J43Ti8r1Ano0isrkUv
E7shIjDrO2ufIYkVcGVN1Kw715/UqJP7lONDa7Pv3p7zafp841Rjz56Wzm+NC2Nw
+IqFq/dEItmU2ZrsX8ZgOw8U4+vF2orKHT6AGvYOWNqK4aNnzrEw3tid4AzDNJq7
BgoPP3pJ7taCwCQBYnvV+eEJMDtfS0QWD9FyC05NBadKIV2yG9RzstP7liOvNS1P
DYm7VaithT4f1x4+thg3Do8BuIEJyRNkYNwyBraC6AUyRGxmziJD871vnDQpAU6i
tOG3khSPeWg6ZGqchyG6KvTPIyHMhBwuEiPrJC1TPlrGTPOwcx2VnEDuk9loR3Qq
mdMnELrAa5P9xNz9Fr9Tej1MsLrQQvnNcfsy2WJ+J3cCQ7YZke1/SuWycYwP0xID
DMqjN/zDnSFw096SgRhrZ0qWJG4PFdf6CbgvHAis18cYyUV5IsoZ/TLf+PypG5NR
/l4PeTmNY/h4T0+xDODepspLX7g1UuJ8NDMp+0Z2ityXQZwUTyjbQPBj/bMifR03
cjz046yPivF99FVkkztycLdMpA9l0u0RajieqAPlcUbEYc8fK2vtUeuSwGz3AUjW
22OK30sFI2ZKUO5VpSqq8AjDNOgePlcgrM3JPfO2JG+1KV2J10rk2CMfptqUwwIU
DRexRxNYLIo21axUDoTtrw==
`protect END_PROTECTED
