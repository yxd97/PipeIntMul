`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/38ciuFnggSLzazil2K1KX85YhgaWS88vY0ExJnSiAFXHhQ76KBM3CG9WkNGMsqB
8Lt0nvQqbw8lPEJJAxt67YvnrmUK1BA/SBs/PCccGqEL6yPCfXc4/TDsONaSABzo
fAJCXkCegfHd37WbS8TmT7WcxQ/Br7IHHg9kNFMzkAkFkwONiMnmZQoAZFSqPqpS
jkujBrVdPagm6h+WZIC4sJGTgN5d/6Qe0g/mj4uL/+NJnRgNQbtoqVNQ5pg0bOWk
9IC8mhqT+3rdEkTA88eevM/RBQWPYZMskQXXRGMTfM6ySuaO0BtIe48t+m7dVBGp
t3I4aovE9qlTneE+hvyH2ak/89kSOfyu+CAIrKdDOhD9EnXF+b/KNz7jFYocr1bn
ywWu3BCQp4C9kZRL/aAFICA30nSXMqJzbe4q60pTJa5UkzfFKgY/0p2HqmWxMBLy
kDNfNgrG5CLh/xrZPYsa03Hy6Ejd971lAYEpZPMTkkc=
`protect END_PROTECTED
