`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1CShK+Bc4uTbgq+N+pYP018d0P5Celg5Q0NajxEuXpO22xxA1lBuFBEUtAJZBlS
Df3LewP9L0OxbyHS0ZzlzZmH5vFKEE8dsi7ffuo9W1X5Xat1ToqfKT65mW3V8pKY
YSMMf+NcE7wkoFeQpvsckqhfxTJWqkR8haSJ9pz6GchsLpTzJF7MxQMbBxvSKPYd
r+L72+EY509Q2gLqawaLKQMGiUkto1vGLf1w+TOhmoxGyzHMNRiR/l3IJdczoWJI
isQ+K1jkkaDaHsSdgMwNoIPw78ytZyOfrl4ZkN71cK0Rc2MvRpN85WxGTUMIJeRe
oHYNWBLBzSINnlbNmfntPXdgxl7x84NQWb+GhMkY/MoJ5vtTM4CCI12BxB93VXRg
W5GR6nCcJ/XmQ6X5pgOkP/R93qIpbsTssNjRwSVv297d0DQfBwkbSOzBdq3zWtp/
y4QaTbg5ye4dlY/qPPiMzT7ybgUGDY9850nGyk0DUMpC5tcCWRd+pRMdbH7mEkjv
C+48k/A9TLJxYV2mgKAfjmqTApisYB6FZWBLKAxwjVsar40W9psmgewAM2s+plLm
ZyMqQ1nPp47hYeKFByPm5vRw4lgONHro5ms6KmGjQYISOgEDte/h4oE6cfJSQ+ta
ZIPRrmihXSETKCYmPBIKaMMY5oyq9iqKz0zYfOJl3YKcaLoT2rg5p57wQjB2TwmG
L/pDXKzh/6p04/npqxUn717bTmjB2bHcqgh3ixFo8ByKp53YgYF17+7XKjXxOv5W
GDw3TMesbjhKsUpFLJ3W+IZdPHmGu2goDa5MM3lc8BFK6FC8Mf6G5aOIHQ+KGlw9
wzD8MMlGt7gH+S6gxFXMm25JknUgi1JdQemhbjsmG7Hn9qNIxpKCnhBrh1bKjxtI
jtn9FfmzXavw3o4hRA0IK3xePMBn5+K6emu8SmJlB6KYQSGOauX10jEjGgfqRRb4
mZmM42L260jRkC/48Uagi9S3ugTYcDp0ioujqPrS2jGUv1E1yfakCD127Ar5yAzn
o8kNvsGZDPAt5K+asV3YwJWT2sTyVKn6rNKKHAlezUmofoxrGQbrZnv2bjBh9tV2
SeoK7IUzFsOknaNTbRtKysdgNfbdaU2Dz1Hsz4+U4au9qMkgzNYD+AVCVi5H1af3
LvDWC8gCdiDGuZQW7hbfmaNVYnd9MLPHSuM2bfrz13fKWlSt7h0G2s2he2Mf7Aob
voPWj/NnYaI02b/J784xo0zvoEKgvGLrkVfaYIp8bVEpjIv/nqCVl0bNSVmpN8Ul
BtTmZRXaO5psPIbyzoy7pFR19UmBF4S5hOqIdbOWySJ7zOxOhHg9iPDaWu4Snlhg
zPLzVDa/kAqLaTrkH2c7Gs7DFoDgFVgzETeJrPyd3x+5pjGtakBGecgToDlWzM/y
/tSAZLJLKCtccaUul4QTGbLq0iwYT6DLLPg90ZU88IwJYL2mG1DHQquOv7NyRV6K
yJw060tTArnPe6xeeiSBuay/MZ7zUmqDkHmnIeVHIXGGFyBOGliQrTa/Yw+lyIls
MnRhCx3Wcx1oMx/qQWjBo9wB/NuC+Q7YikHLP+MBHknEZjkV7gs17GfrQNpL+bee
qwxdmg2OOvl7M/8fZlTQk/m7AwVR7vunUmZCm1ianeAxptwyRV+jwD1G6j284iGE
2wwKu27s7HPRCTmdNi3h8m61sDuXi3U3J/UK6qb2xT8k/aJ2NYrkiRGBYGz91WW/
1xKnBUbEKyJvvEJo8LfkZp2MJKGWsOmPPydJueUqHRsQYJxAb/IaQKkN/pubXw5Q
JnHDu01hs7L9wgCxQsnMA8zwpZP2qYVCFtbSv9tBWU2Cx2OY9nD7wJSU4MtS+bA5
g9iSmO//83kfCmM9utTPLsJgll+n1RoMAJpgFhlzTP8MI1M9mBn6Js69Q+TcKsMH
hnW+i/vSEKy1xu5zn2jq2BiWD9Qwz/1FYC/QUx8LPJ6QVkiMtK9HWCH7YOVzYNK5
gMTSbYNlC5ZsN6vnoHp05pJe/H9fTsCDiXEf86Rzw4reG3FE/W9odfDVQsGAYsmq
FSxCCAY4Rh5roVq5CTGCLMtgc48nzEiN8ntuDsacxkeadaVgytHS7w6/NNVYiulP
uiHty7QfMpm/Q8wmDjm+P+LWDiQA6VZDOd7XAUm7LIXwrnGjolnV3LMDJP7/uncW
+bInk7LONxOQtFcdIfueZIw+Cnlsvzy2kROa4CiCTMxA/A3Z1bQcxvDqErtU9gF0
IMyz7LSTFjgXBgUZc+t8BG+lv3iGIgIqQy8UA7h3Ha18YwyBEd2T0Y+Aw0PfaVIr
cR4CRAn8VQ5C4VyT5mzvyqTj/ZqPInckwGHc5jdScKCYT7nuWjP/qDARFGj1yg49
GKfw7Jw/ygxiwMJ0Uy0lGBrL3RO11kv3zvlk6Jp9Iyu7p3NDsvDBUb2l0+Nuuqj1
GloWtngkWo+LQx+K2eKx2A==
`protect END_PROTECTED
