`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zPidldAp/nE5sSQCmXqcCo/XJG5LVvJBstEjUuATIVuE7aY6H2MWM+ZRLB5BjrkM
6OLMF3zDtVSWDbt2kZSuh6a85/FcmKtF96TwocHbTq4OzAx+1KMimcqjjbcSe8iB
sO4oJBHXW1YWfiFEESPG8zsvtFGH9beh335/DEyB+vgFLQ2X722/NvTl1nzIU1Uu
n6C50VMDNF4/Qs5Dv7781LpVb4zNeCcD70/OJHcDhT4au52FofzdRZIDAZ83vEEg
CThckOX0cayIxBfrYC0liQ33vuXk1YDk+5YETVGrey94sNjWDBB5KV8uqjEzZj6x
TatpW8RQJeIvljtn6MrkyWsIMzVOlVVOwW06Fh2bXUDIPNhKRRXgNs/za15Rpyw1
zkDYe+3NfECudZT5q+6vabvy1jIWZFNTZ36K93rw7wA=
`protect END_PROTECTED
