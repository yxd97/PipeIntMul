`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSE9wSIW5xWV10X8DZNMpF+Rnzvrd9SVFjizytZ7ArSpiywfy/W999g4ERSjBjHW
Q07ouQsBJf59RM0qhr7f4byFwlU/5lWCgEjf/YrZiRf6W00hPOKstQ/DbVSolE4l
z6fUa+HMaC/GGcgYknL1kNa7WMqtQZ8d2vktHxLB83LvQWlkEeIPTsjVclRoggWn
xTFufBpn64PZNTzxhz/TgQRnN7hkTMwyDIRvJu6rbL7TvVSV7ci3uHssd0n4OwVj
UhGoYacJIwxxph3DI8+gfLGyScmnhlJPCcRjj+qVE/Xf+q4Ccz1GGyozknHKrOou
TEGINm0HnGdF6vUsb2HkI2K+r7Cb9nCvZmzf9xKuKyJezvnUa3ayiGY3ThuQlM2/
J7du5ysgWqtgx/79b/tagnEaKN7YMq6jsm8injoMnGJtGNCn/1vcMpvqslpXX6pq
pklNJw5brSUm/LzuT+U/L04UGHy3PoW0QQqX7s0p7FdJ8G6h4Zc+zpGA7IkRQ74k
+pRKXYRf+moVXVEmOUg0aIVIfw9M6uOLbNEh7ZQ4Tm1GR6a73EaRyKHrG8g5LFb9
VqxBQKRMYV4A7iNFpQnCirCDnGmjX6cYqLwkHBY0kGh/i69g14bL6gT0h/H9O6ss
cI8Bb1GnrhXB8xPQWweHeqytnBJdkBz8R0SlNMwMWTaox2ZhA3TKVgplj4J7lZ1y
tAVHG1eKPyENaib3I91Y5VYm/ZHqkmmIQr/W/7NoCNnXmjbG0eQYtyWeYCDLEyFn
vYeSjxYq274iweqN0+PxzKoPQ7Wc2k0U8PCRNV+GYkBpOgxy7UhUPHKv1nYOQjSF
pMh/8vnoHowLXjqFzybP/GWzj/foQNygKs8q204rVSM9duR+AfyGZseP2L22xmZ+
pjwu+Fd7ywK6+vNvl2PpmZvYiP/Jm6FA5/hFkXNTtLbFioIbFj/HczfPpLkUdza5
KnTipNUbhU4duLns0sevlfHQEWNN5F6QN3pWG8tZzHz3GNq/GDG51NMj+xuj3ODl
iioNpr+1dvFtVaPKpOiMF9wm9R227l3aH7W9twMrgrO5oDAtce9Ys1YLTJX+neTa
ZHpB2ngHus74fm/9a8iyiJbVet9iYJuAB0/gH/d1BZIMfrc8rFAcwDfDR0t2acMi
U4hlV06fQsnaDRALslfmSUh1+BRjrgRfFlDFrbj47/KbDj5He+H+aA0aeCUERxBu
cKZ8vINGmNc2xpxzg6+Fys+uZ0Mo03bqULs/xDEmB6f0RCypztXP9OcnDJqs69Pm
RI07uLOHOUABY62krT7j1C7EkVpfAa6+t/7ChNurVPAH3wt29spBFGg1DqvcWU1S
8bMNAuHq2t3Igzb9PqJR4gnZSy7imh6uoP1Zy6JmgA0jq5oSalKNsUwNLtbsGG/q
Bunwhlt3RtvUHPApMlUY/pvNoj1m/OTEGLUgrseMmF+JTsWmZReOGbWNohZ8bpvX
23ZKw23uKxh1FBy08sZCf7FE1sK8yjhs8UrfId6Qw+Wsk8WTOnBRz+8vRYKx8por
RsJsAEkkU5v1r7l+cm99dC5NxscXoRm0XdDtotmK60xz5ktTOSKKkvsY+fEcaOAi
94P+IxWlk2mVoVlQwliKWl4aMX5rzQarN4EYjyb84DsgkyRl2Wzw4xnBKjH4eve7
ytoVt0Mna9BM2Dd0FzhmZi1SIclBKcJ6d/n/IOTcZ2lJlnZzrAMQvpdYctl+NHaa
oLZCFP/VYsC0VOzYH1B5DViqhS9agsDspSbjVs7JVD5euA/ToOI44bnUU6rt1fsI
NQNrH1mAJy/cM9MqxP+V+Ztjr07+FkLemQnJSsCMVe2vZ8ElVx48BfRv3FE2qK3R
MrQmJuAEPKGO18h5xOZbQCyK4jk8Gmf5GSKXMZPbnSqok5thsDx5pVS9ytTLdtrW
nLi3okdR9kYC90xOPnKYXIXyp+EEwhZrM6eORwO5mK2UmCZp0mbcy0y284yJoJtf
1ZxDgn+GReBC245Bl36j0f8NBj7Nazmva640BBFx01osFy/9mSWurG/RM3rJR2r4
1rOzWTY8eRzV9yozHTVOCDYqLR+O5DQwBrwZmh+h9kZltz2WXz2IZy57az21LYig
VssqfjyVvbJ8F3WBtHkoCLuRFl8Tg24JzxWHcssYPdddl4WHxQK0KnOpFZGihE/J
fU4kBmkgKxNxav0Mtis8QQpQCxGt+oBw2Aq6ndXJ6Flomdb6disf33t5R7chUCor
u3vEfsPCTba4b3wPzos4fSND53I+S6Mzh1Biy7JOr4uIqhuuO8r6nmR31cIFzbjJ
JNfk5NquVuGM7PmshFmX2jj7ywAhEVGBn/Xh6/IIKI2HUDfSAdnRTsdE+W8Vm2eB
1BDyNR/iZj1555qAvYTKT8q5tmK/qb4IvzLs3stnUQHNhfd2C6KwVyRYcFUsttl/
q9aZFcXKNOBXTJqe6RUoDRQlHvJDtiJ087+FQKQilMlaEIznilYT3f4xiQGg5zqB
sf/bnJH6PvsKHQJngEySsucugO9OHYIsFLRsGY2//f9B63skmQWlVNOwDmeQpd+P
TfRLlWJIS2+etWkVSHQyqpFo309HHqG3DmQoANGX51L7CUQtOfJ7ka40A4ePz7vx
XLOrOIH/0MVb38ZQ8q642V4JWsamzbiJ7TWbeveP2OJCDxoluRZAbX2hjvK/qkz0
l67pknLcxXojj+XRbRcA1BHzywBQMgvlolbg13uJq3N+Drp8zy/ZKvbSE+TisNra
kYE6umnFNywaJGoA2OclWeIJ1bmW80Gxze5wTEzvsjxLqy93l0KdoOUuSOfaT6WP
eabe0QUC6ReAKKPqp+Jz+o09Tr2EKp+/w4ZWJeJcW7lspZsYC38h5hiMO1mmzvfi
czW7H+tTi0HdnPBa2tAOX1WhmOcwS88iHTELoZ/c/aiYOCq4Rs94BOFp6jm4fEA7
jXtvDTPHuWp9ODVnZuSkoY1K79ahGYde71s7FGkXE0x87Cqx6sEBP5zPqdVyb2fn
f9gpMk5NPD66SggjRgh5Mkm5WsL+uXjKt879sCj6hf4+DOZ8Hv2neeXGJ44izgO0
N1wY21UfqIv0+hHjYH6T3Mv8oLk/RZrK1ECvgsG6+TSj+qfDD3u0Ml4mBr2z74t7
3MVH52IdNl0/JRVB+KbETlHB8fqNQLFkGScRh42B1IZqEgrmsz+LV2KuTIbQZCV6
2NR1+OkJ16VTbuXePTC830ai0py7qHnrhhFPmrJFOimsVdBJ3BTq9f8EhU3RBd8T
am/5n8x2UV+hIKMhgXMEjqoPdsvuTO5mdMAY0uhACXkFHDMBjuL11LRudkOGYSyT
VxiBHIRb6dnI4T3AXjvr7XFfPNozB5/w5Mhrl0onKJKYSEJVDyD6oqoWZgribnrj
oKVap0Jsq9dXBPRxQCXCs0J46rqJXzrKcZkElHrNU9UBXuCMF9H/ZrlI1dmBHPoI
7FQz6FS/P8O2APlQdOx/kQrQ/+Q9szRObbwT9FWVK8BLlIXAZBxjD6AhCvGmPMdi
CMBEvOVtMY1yr9F03XzdXzXVqbjvJ0oLPZxg0yYIWncTyEmIDS6Dw/Z+MKuy0XyY
gMHok9LNSkX27W7HjYaV6fxnPUFUfNoQH2TryfeZQViDvod8jCX8KlKMgqmixUmV
HmjMpTvcf5UoPck4mxLCSIb3wAN+ElcBDROL+hY3cWXlrU6xFdRUMUrKYK4pJTOi
7gr2z7EvUJYf2EyZ4WZeGL892St2vJx9EXMAyBenIZ5uRvdyh9W9N9yJ8W2O5iPN
R3EUsCGB2xEcdlfbX1a6pwadE9OgaZO3eQnoymGFABCe83dU86AcSKaUMxtRAq6s
pj2wR4m43SNLX3AlnM/t/OUgQzE+Z+PM9a98BCpPFNw/w0Iifdf/CdV0X99vLf1+
ZL+YKpugKrzFrmo0zlR8muyHy4N1T7YB89eKCoaReoA3d7q5qmZeV74QVm3X+9um
UsmBVguMrrJOCujiRpZPY4GfZZfQ9tLhKlWqvlwllTs3MBnsmm1tRr39TQHAwQiY
4WPJy4Qol19hQgLDD5kXN6B+q+VDwUKiXvhA5XrrtiMBLYI86NxYBtXKLYX6jPyi
JH58AqB4oNv0M0QBJ2xwqg==
`protect END_PROTECTED
