`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
unhtvDngjekqNzv7iVBDFzq7y8Fe4OP1wO+ZoA2MTdhUMdiWQ+zH1Mj4bWJym1DW
S+umG7Zdg/KwAqHsqb4rw6oTokc4fK1Q/yIpcGd617oMiJHZbu7XVQVGcZ1v0bqy
Dbg1XM+J9ZL+7qbK2MKM6TJN27EejPmdBCZlrN1lwPnoSlYzeFWz/BzS67QEUvt+
JdzaUhFSzVGVAXKM0+0F8Ed3hT4dhDXb+/7p5MQcQUCi+Qqvif1RETkYktPubQvW
cDvk4XsmYdiyTykc+5RUsJbC8TrSrGvQ4lP3brLQWEFqKbnwGxE1Jk3a5JYJNvEl
2Tlyt8HpLRHuxxlYm7qoeuerQEJjoWPZtElVtI65KPbfcL94QX/9CRzWtomomsBP
/thgYHKY8jiyKnDF6OfVnLtY9CxEKhlQ1wphYz6gkgsmxQFGk0hSiaX+P96odf42
M6W75x8mrn8yrP839bwq6i3Ix5INcpmGS9AHhG6vkJmVPahX4byBdMD0ckJtDbEJ
K9HqCZZjuGcgrnzyv8xtRP6JR7gi0Ao12U8dmqoihTW79HF78N9t6rEDfvWH7Bzt
5QknfVI4nIFue0OiAA7dvBxv3qlssMr5hwoU2N4OHv/RB447Xjbfhg+wtgNCFSwt
aNH6pb86bMzi8oiKvUd6+A==
`protect END_PROTECTED
