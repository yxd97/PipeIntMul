`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTik7eodlIwBv++ZiCdSFoaoKqIBixvHCgT98KmdDD4urW9N2U9jV8VYAjFQlcrT
mABzPmBm4sOcWCF99C7jTgy1czP/rjqfWu5Up/AjL+9FCFrDcRRm6f69bCrYzmj+
pJqhlrUFcHzOq6epaeF8iyD4eTXgbj/3crZS9GBjUyzplrBsKCQ2WAZ3o2iSXyAP
j3NDUM4fTQHtY1XjAg/TpvGD7XZO7LJJbe9N06+VjM6ZgYA936ntNXeyjltRNESP
tgENlKjOAQH1xktBGuJEEc0Mvq0QAW2R/ebQpH+GzqIncD+SyiWrtwwMrJV3B1Cg
ev5puwxcZtn64tknRh0RaAoLDNCIk1N2NZK+Vm0UA98Bm/UPl/S6Pb0Xf+5YRCQ8
CZUBlneGVpStu6jtmT/YADSIOpKmH6AgRITRCHwhxzM=
`protect END_PROTECTED
