`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IVUjsPUhI3xNCOZgV+sFOUrvEo0wubvY+O+vGS5Nu3WzPB7ia/rloVzS7lMBSv0s
Ix+/n2Vfxj0BgyMEp5Z2tFjeUu8MXbqGT4tzyZa/5CYA3wvmCoxYMSZMlHCEp4u0
3/WDNWKqYVATl9sQHlUpdGVMOTRrVseMseo946FiT+EvWBN53wIyU+BnWITkEgUx
0vWBdVN/gjMht7PrML3tfqsRGpN5kSwqJMYx/pJGNefSwony9maQRadk53ZsQrQm
98c5BoaqWsfwoqzsGy1KqCNSZ3NCy1LgztIDfPqSL9NtDDL+efiY2OphCgMTwpAI
`protect END_PROTECTED
