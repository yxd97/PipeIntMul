`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkQD5HL0K7UuMsqn3a7NSC59Qj22VTXYUcYQTcj6wSgG7oxuwSg6eBxzSz13ms3/
+Vw3ZSDDYzd30iOtJXt3+XMoYxkMh8jQpuxyP70ejdMGMkDTWN2pFXHkYCeHTD04
mfE6s+B3ig7wb3KmUd9bS/pwr9EiL1KNMuiNVVDynFN/ggmoRWAnlDKEvvVGqvdL
x0nZnDQ3XgZ+k1aX0AAphZKJsEv53eelYKo3l0dwOHzloqzIsljsCXzawJM8ZAt7
4KKGFeRHc9L136oglOGg19eWhW4ZXnEClkZOOddczSn1HnfsEthe01lL4st00i4K
uII1Tz1FZidQrT4qUnYofRf+Msm3mzVw2IuNzS7XLssYBNo7dYNjW0C4norhXmVl
Ny9KIrwjnCGoAK65rlsXu8Q1tXs0tu1AeXJHx5N+YaC29XZUs3SXZB/KQItjCOsE
iJCQDY/nCOeIZlmb2IkaaMy13S725E7C79G064wWiJNBB4bMzJq1XX5uZj86B0jv
Okl3NAmbHOEeAx5fPYA3evVb1WUMufUlxvFACtKm5Y1BEiHoOn5qSnRQIj+JVvdR
tbtcBTmnUo9KUVG1jZSdmDxM2de5NFgQd4vsgd3c93gKEL0//sikXq5cgJtxjViC
H+Ie472rfvHuSG7rPR1vMwJ81NpKviajXu7jCSETNjH1dssakwIB19E4E1aODwZd
smt4hXoczwZacHkyyEjpNGkNCR5kvSfVUDx4mQssoUSvK1S0gW0Y+uSv5neoXA64
CXacGfdTywEkwY6iqprGjA==
`protect END_PROTECTED
