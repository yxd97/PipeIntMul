`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ByX+PQwv+UwWpLi05wUh9XOmC55ERhOCCuWUbiLck/rgte7QWvcmEy0xn1AZQAm3
qMCqC3y8NJqQJNyX+2J7Jr9q5D9a0nHynuIQJsXnMvZ1GJd1g1dlPXMwTW8YWEOM
tuY+RJozNnw4P+aCwlB3wVB7zLXiTDcTQSnkqpEZ4BCMWsWSTcuwT8OX0Bel3nKu
P21IZyT4mOm5X0mQqy0QKwNUwI6uYGCsKL/2Pk3GFousCu8LubUUvDweniIphIce
/7Ti3Hrt7Ptco+BLLHhwYLAutHja9hGtm/Gi52ZDNx3dJBHoieN06zCXI5XgkFWV
GqHjKtpZrzQLjVuPKxhnvl7VePDAMeC7uGdNIoNyTDbZBK+8/pchuna+JEV/PKfi
pB+u1CIQ+UIZX5a/1icAe/wFTi/l+Km+jSJGioonslDecgvXOBNdyfUO0Pfv0U1w
dgLQmrKuImXbmjJHwXkT+RQ7sD5jhdNXw25v76JBL2sV8fFpCI7ZsB4MNnc2SsaQ
JyB54fOAJ6YL6AKj6iJ9JDR06qJSz9xj903auv7eqCk=
`protect END_PROTECTED
