`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gRXW849s7Tri56KbgNy2TzIK1EE7oh4Fb7dH35hbwHOMDk+PNy2/MO2KpkR79LFL
AMHB6xEKeNQlKFYLOLc5vou2aN2+l6UtkGtuFO0Nz4k8eojoeH565Cn8INKBXgaU
K54W0D8kNHXfNtZRzf0U3jbhDeW/ZqRYEV4luJTOVKs22PRuMgjPOyWczFaUsU4j
d3JD3Jc7ySk1f/KpBQY9yVf13pXZVqmzmCj31NLFlEMZ7HIztVsYp2rCoFPSz2RD
`protect END_PROTECTED
