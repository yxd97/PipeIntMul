`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUuz3wM4nvV3KuNLW28FnoG/cco/778cnqPxGriTcJRQ6TI+febty2joctmzgZg6
NSUV9bFZfaGRI0gnTwl9Nt820gWw20el2aO1ECkVgCWgEANL6ns2yua4OB13WCX2
NdsnfGqdHu2ReZS/zBpoAwWmAr3bJPxwton9KSVpeixPB99GC4sBpK27fp3xtjY6
sgi4JIfjPjBuFvmOKlz661ZHA6z4CHEy4cXxHEx66NYOfAMQh3HDg2vt67JrV3rM
AL8KsNoSQwo0YQnPzOJMnV2PYGn9pR27G/8NxEOSA0FkyeoOoQjSbwR/yr1pWQdN
StZ6pMGMsVCHQKm9Z9ZGdj4pLSHs2GfmkUHPSMIUKCRWrzS/+nEQzORGm9TUyPtR
M0xHkWuSllWUqAEWpslQ8iSh/RwejpXIrapGZAadQPcMK+nulkfgw9fQm5a8koCS
lrOtmDGWOVa8/5Kcc8H9JQcJKYveIC5X0sCBmWR77HFs+b0lhtFUWeWQuJHQqmeq
SPd8OTPR3qqLgvHflFdvNngMxlfa5Jju0ZIHVaZIWGCyx7+SWeVTmH3HS2oeFXXd
LhRYzOBoJnZekUIJCr/Lb6sXIbEfXL1GZ+9xsx737iUZm7Mw2K7T4iHtKmtR+LGE
`protect END_PROTECTED
