`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+2hDmpXCX1FHRfaw/WIlIiaGGAXDA99aFjNmicFHss13Yf9Y7LPeI5/2acSUdgP
868qgSgL7hJmWnqrCGtk0D9OkJT1gLysxIEUIY52rVCT6m/lRpwsaChjxwS0J5b3
Ti6rIjG+lmfJ8w4UufMTB20es98aAYqtEDDAZ70FRF3ifSkmIlrfLgwskdoCmmd+
uIJKoYCSy7yMQKhYuhdCrg2aGLUtRwzw3bMaqkgMp8LWxnDNYVyqKmCAf8AF/S7s
83lYPeQNv5GN7ooYDBcatXkXFwkMl49tkdlmhjRuzjwEjTK7ag/C7ygx0JB17X7i
ZYKu8TPoYh4TUfnGG/cD7F29ar5efcm1HIolFYdlenxu6ml7pdCqRquXrYpDOc7A
mp6PDSx8YV03AmIG2zFlo1CJU0bragrYZuWsEgm2OumLhwOuz0dMzYwZ1dudi2/C
prgQexK02eX0AMqxd7maJ1TuGHV2D5boS6UTJPOD57vVCRixt3yJ2bahqcKq2qrH
7Cf+DyK8CM45DbvX9tqelE45MpvTkyNYTA9kjAlIsK/bOYFO4N+Yqs2U375+3lgZ
Z5XqwBfFaEpSS5RU3kj6D5Re5l4tvNnyBoBRGwEEvDdICJEbOzWOpRahqOJn4kvB
W8js17sfN181WbPcHYMhjRYdPxyMRZyIW+XVtyIV9zG3eMc5jY7GtckpYyC08oxE
`protect END_PROTECTED
