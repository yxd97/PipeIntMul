`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AcJ9KBwTu4Aus6hY5Xuht/WnLIHxKHOHnNsCXi2i5hsinIk64+gKRrYPtl5LaNkB
c/nkE8tkee8+sniG6Pfu/cMcoVCDLJ1ftbPLtyNFsCIacOYILv2Z9PbqmjjODhfS
Tu0iizxpW8HFFfDjbWSabimW7fmwh8JI+0VXosK11oy7i1AVvbCUtyr+zf5FCawx
LDBMY7bq4i1EMB1M1lg7QycJqoji46WI/tAfjFCOFedgn3T0bBAAfKLopq76NQsF
r5ACDEhh3gCV/LPlW6Mzi88KcFGkLMOAQ7Aj3GlBDZw+/M/y3w790UKokyXT5EGj
xKYcpVfun/HSzYMR4vz7q+BG4uYqX/XY0iCAo7JfSr+7LdnZHe6qWUG52NnKbOfJ
SEnI6tG/pH3yM66WtaVY9JtImGYXe8xihcKT5r9BHGT5HIT69hMjTQketZDz5zP3
z3PBDUFzm5UOdKuLGwV5ypFnBEEZCUmENPcQ7Jgsn2y6V0ZCNX9jdbIlnJH+NaNk
FyCxTUHki4Ox+uC8s3iock+DPmcyGJG8lw72nw2pQmnRhdhRwTXW3CviO+ThaaUZ
`protect END_PROTECTED
