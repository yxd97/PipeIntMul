`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PSI0pC2g0MzjA3zTVzBS7hztd9ivKGJLG75OD0NbzwHFWX4WDxK1+pJWVDLgM5Z0
2/C65GnEasVLvXl0NI50VEcOszcjA8av/0eFAlWIK9t/3DzCnAGe1Lf4kCH9jnWL
rXtEnFxJm3rHctdA8bzOsPhn0bBig/UEdEHTXyE2uaxUGGHq5znaXg4Cqm6FX9yb
/GCPitR8rTKscq0ogr/qi3BlSExMVuXhJBb65dDWzzRK4AsWKdgQxfc+NhRqUsts
A8j3lBBBnGFwgMY+h9dDeTPUN65wigQAv4QbQ8q/Hl9M+kuIHw2OY51yFzMJPZyq
CSkWIazo9Saq3Jq85GTeLtSrhPO3spqQrVZOjLBGwCO8apRSN/9nkLSh3wovW35h
ETG1v/E1Z5QirFICHngoiUEQ1urBJS1OxjQyW/+cGXSFjokrCZHvOa5qLewUe2U1
Ic+rf/RJYcUlA4eN0t08l9JjYYgMKQYog8Ha/zprDQo3ZOD3UMTwFAyry2P37tlx
CCytxIXTHQ7Em96CBNlLDvNYWnaKOBvA752pmsxgBxshKz9+MrxRH1k+k4KUhrnH
V87KAbzDj1fshKP9RXLodU2KWuM2+OHCkQIPAzC4Im+PcOfjcaoNc/4xwyAMFFII
+i84s9EWkD9yzPUBBymVguDs7KBLVrnaHeoRdfTTO64XoxMq4kbjjZ1Igy007wKK
NqGSYfeHmrW9DaIB2HY+YRf4GoQUvaDxS3ucfBhsJWHB2TPkPIlw3OMbjJYDwhHY
yNGjyq26/7hWx7TaA7PqjPq8kJ05G6nurUgJbwsZYcZc4V5Bs/eJOLrrl7QYDx1g
lTb/xnMW5lrwmuB9K9whkZvIw++0Mwp36wnKDHPmoz9A1SZTUUZkSriChrAVLeCG
soJOi6Ca4w4OSB6/nCPNQnIvRPNF2ffmgOQ2uoSqFoS7jXXs2eLS0OaJLJ4MsyD4
OBrxXYXlrDxMLN6lXQ9bnp22o7PSlJwrQL49Tk+7N5e9IsGjAxEM7NYkIqFfStBe
1qU269svQEMnfkAldv6qdN+aK7iOR6256AFPYNaxy0uB1A1kujHNlGRCG24JIm09
fUIMehEMJ0YYIuw0rpodssUN4n0qy3J9HNarEsbPd4N78JnD+MV4SAobPC3WghkW
Sd++hl93TWj/QcwY4CPd+S59cUDadHPNns5XHVnqhAV6o9AavQI7x/Dr1VemqdI5
SYK6mwMfm7Wp9S5F6OxAQMa9V2bzcqqZ72e8fO5bapiMI1vGaH6PDOkrpfUszWCo
YFlVaUHvmcqSNVZ9RHF5FTs+r2hbvkVLrXSi6DZKRd6jcbW6gV4MmvqQ8PadXdQZ
lz8K1uv0nvJ/U69y6FBORbkcdlCg7niFdgS/FIf0UGBX6zqpceKB43YlXG2dxzKS
TS6jPJXrOkJIZiY4vSy6XkSOsj5L2G2mH/9qmkAso+0qazOl/jHcGXxkfjCzq582
94dh2WO5lHKfxPX/arw+uLo1wKeJy8g8n9OYLNJSTCb8JgrAdy1FCckDhmyfFW/2
7o8kdS2nsG7T2uQMcvUcfpNXM6JVCF8bqmnHkiQbIqtyCCiAD4uMBQP1G2fJlHxf
aFBrwPqPnWYLG6E6agEbEnB1iJqYMYlz2r8r3hBYCvpLi1Yrnwz15Yjhw0rFS+Lr
OerpqJTHiqla2wRcb8rAD+P3L5uUQfryYJHt7KAiUN/SeDsXOIJLJSWmxDgk0KyK
Ph6LxiQmVVSRE/TrHGdKUx8qVyyKJs5YtbRM5/YY+vrHc8RVZ0u0zK7GI31/OfKz
JHYtjdR0fCi7aF0OtDKKhlRWnd75TXZe4J6Zn76+FwAiM5b1mVKIVEZKR1QXQVYw
1X8WARzjv4aK9/nqHxG4PFvcS4qHC2lm+tEKczoX9p9xBU122gYPr8f520/pRc2O
hAjaWfZe7d7A8sqylodZKcekqw0KnHGUGGFhidQpU+FZ2J2Ju2w4goCPCkoOHMVz
Skx8pNsAUzMfzvspF5MzGC/BwR2NgWMm0h0qafbguAu/gGfuY5sBXNxDGwMtg6mv
twLPvfVD9hUMu6eh9OK7ZcwFqTbFJLlxJK4odxMWOBr0pLoCTKK7r1FK4Wr6oQwB
Z596KHTb3CUYuAWhQNZ7LvgCgqDBYW54Niu+2yp+qmHhHtOCuW1+hcn5nNaIdZEX
uKNa4H2dH2pe8FhZhu5uAH9JMC/+b7TdvhSUUl1+rFHxGi/nq1dMhxH91jpnXz+k
txryaRx0v0p4HVxHcGp5vHRMrl+J6X2rU0epGL9jyKaIM4Ak7SroPWpNBHyzBpA+
EGO+rlxNga+g4vo/gRyH/EY4Afj+m5qH5PPgdeN1Ykm/JDW7dv7Cy/lgdffKqS7Z
Cr/hWBzj2/2k4ZAvyMHxbNgdBnE9vJcSgDx6gToMkZdYubD3Dcdqd50qPl/jfnZq
Id7DOXhmV7LznsJJzqMmxfVgsC3INUNorMx3qG+IhSJNSxv7Vxkx3rHi11xvegLD
ojiT0ZQ21Ia0GBa5iqxkC7pRsIvrAvBXWA0QsgJ16OiXKomb3qLRz2E0YcAadGol
RIZh3X4QqhtDKs1ryP26/+Zmd7Mhat24gBBaoyWNsqyCG4Ezgo791t5pyXWE8Vpo
kH0DMH9jevTQ1D2BGU1rnGgAbFOpHv5L5cYQblETuREiHq+ZkFs4imR77KWmegKb
pWfPdIeioSp7rfVZmhImbIKU5uUXo4+rOnIjhKqXx0w20TCuHO7FnhCbTaJahe84
MgkdRwE9S7MK8Jlndj0Bt2RluX3sy5ePiXx1tDWG9KWTwVujap0E8IYQvASAnIP2
67zW9Sa1uSZOPCF/cTVUx+DyVw45yd5W7jQu0JNOGKi5K5+tXi5FjsDGAvtcwFel
l8ik7ZZk1xSEQLh7q0ONAw9weMID6PXE/Gk3XzAUMwmEBR7vcBg8cAASRqshQ1Iy
kORpfkF8dfMmZXYpF0yOSOlZzC8kjYFDlePe6aqx3bzUWj3CcyUZWYuZ5poUeYxb
8Alcw4mfliBYJBp5oZCAT6pcn/k72LtxRb6qCQn6s4RpCtYIc734f3JU2nMFBqP8
sJx0ug4yCJ23rxqS0OgXbivO+Y6Ff+nniJd5H6fWmjDCcj6wssVxJ6bL3yCiEFWT
6/dtdMqPki4EQpUJr1nqqgrjSsf6NpR1xvBEvhZrI7WQ9b0ioOmSaZOazXSP8ovo
NXDsbw49JaX1EAs0gQAIiTeysbWq5rlRJbMomFOUIsT5Y6JpOCMe/8RhV0js6B/B
dQ4sJwDmtdY0Iz+NyBEtm2xZlt5FlMUU2MTOhEqo5EaaYw2habY2vByCEPajZBqY
QrKu2R3DdQqmWvvuMfX/oi3GmwuczvHEd0TwOOFozRI6RXFVs6obH0mfBV0javey
X3VCavtF2MF1nx5K2OrDf1JTNE2tjDaJOYOHhRZ9O64JQhVSmAtis7QmyIXQ0dGP
vQXGkaOQMC3PP1bgqJ0t0QaXRrRuYpHgM1X07IfBhdv7T+eFAOfGYn1h6jq8FR+P
/tY0bsKIXfST6LdaQ7M3CuENSBdLZkB1eI1qtL4exrMl8QZoaYJLyu1iIWHyplvE
h5VnFf624dEjUQhmV3IXlfpRzhFXhcLeLsRyzWjewFLKiY/VFk2JMSyFruLWqH5A
uY+yNjKYI577EAa0PLfkPwtaYpF2NQT6L/hRck+SMdMyXHyILUUwsZVoj8x8UeAG
dOur4KaVoFEb6Msu18dixnufVA2yotp1/gPL90ALGwiiJh5HyDH9p9apO7Gn3veY
hrR0Qo3Qd7UgB0rUqWTsLxjKA4flyS3y+XDkCf7pGh+0HZR3qBAN1yCw7LTRirD5
8fQNSFio8uStxQ1oAgK2YhH5BBDZZBbvHudU68p5KB9331brsXfwhDoG8Yok0J1Z
eaLw5/WhpPx51L8e4PHwAEORpRzFyWY7jaCdF8giOOaLRjYQLsm3tyeZEgIVcJJM
InFXiL58OL7bCffWct4NGvvIlBLQJOYY8+vWRP8s6Y13b5/KNII1GilZOueaZJzD
BGsdM4h7MTmcgKnNQmZOYVUqUEI2mtwgjhsLABwRxwNayhO08zj+qI+Dl0jObxx8
16S+jUzfZXIbGPpatJE40bHxd2z62p2itjTfYuo7cdqNZVwcNEidMeqkL90n+YCy
JxZhkLhOenJgjZZWU5hQCFsw6dZFUSyH1tYGaV1CZIeQxgVspSneQ0kv7kWdnons
T1cUFim1qGUMeHJJkwzY8HI1qTmxj+gXaxxn3HSGE+Gg/fJ/JQFaoPjH2TrCNH0a
tn9atiTcoNgkcTah3vJykrWwbcZ0spRWgo+1kt/eMwgD0THHTI6J6tCHqd3w2J3j
P42iZUem7qWjfQk9HFqWz8wsR4lhDe0CASmMzzbtGBRcTtxGqCMRciaH6XrmNkw/
h5K8QWf8LTJIXrwpxluTihdRmVkYdyd9jzfKHVzJcTHCMqlT8Nt7DX54kK/4uy9t
XLTKWHbAXjsHoyNJcO4fU/m9NyBwHK5CMwc5M9bj83oSG2wnpdXVB3pa6C3CXLR7
2hc9N/BRNVsAB1n0kaP2DYfHLyOuaMIpRp1jBQXyK+tQVzmjIJkKRyyjU2gqDxZF
dDxh7GjNURLnbE1SotwbkULizhKfIRVAcfsZPJo/J98wlbDbvDljtPU5seGxDGL4
ItXqulNv/cERWUDGEiwZ/4fyUnBkRIzx7rntsCqoJ7dLL0jNzJEUFanauV6NsVTI
sibUfc6A7K5PFKHgTGsphPdmDBcHlHBueViJ6+5Ejw2ZZpyqwWjucl0JRUVj1Y8f
bKWmLgyLfbNd0wbzdCFbWxvvbAI17Y4CXsUSbuxxk2K4EvyTAynfpy2AbmXgKLLq
+7E+noAFlD9A1EEbz3LfnucoDyZarwMkEv08+cm3MJnhbj7zZ2sMbyc+ipar/w7z
No4RIHPBksmqewyqxjHKw4WhczBp2TSSXyfayR5lQkGt8lWZIpqIOy5TD9vBhARu
xW2fpVzszvPFEBIpr46MDHs0BMyfK7eiGxqq3L/Fr4FpB3OpDuhANMX5EPcm8nF4
qK5zAvEZdjJg43Ia2lfolUnQ2Y2u/CwayN3MRWVem71lCH2TD9BHiyuyeFFIN7oe
OIY8gH5UBzKoJJajB20ifbDAbKxARXEiixku8Iff7ANVmuv7N/0nlTp39EodmlUd
a5/13b8SFfI4BQifqRRWVX/a+R3gV3YtMEHc9nsxEkvPKKZzllFltY0CtpU0zqLC
ZR8G6cJu1njVmNqBV50sZqdQNmQUVPH45APGF8gwiCv6BWCZrzDslU8nVbvTVXb2
8QYN19gopbmo9l7RXf77vICjK9tI4eOoSN5ELvjTINP4qbHSLk7/QrNtHrGOLURE
ncDZobCsWAq2Yyj+IimvH/LOhGq9TUbt5jJaREmNuQg+8OS5ym2+1Rj+UUnWgBYu
5KUgo8jDgm3VdOtIZPof5EyxyJDBvZ3NpkOPAEvo83BZCTLrQvx7izD6pakLSEUu
L3g2BzQG7xgsMvHrSOCqX1HEJUHmF+HnEGR5R5npxNWF9X4emFu1Fg7VDWv8dl3+
ET3sKAkQSzatIeI6F1zdhTqbC7n9MLLBxNaUXax+N9dzFQjfUXxvDCMdbhnwbnxA
V0tH2xKrt4PUlx56U/hj8F814PAqZ9Wp8LUR8qHMF1BZAG/HPWwbP+WBVD8wd6FO
MZIhLKVzgr+WwJ6z9xEsx+YsCwECtQrh+csNvW7v9nw11W3ZioSVsNYAmsQ4c9rS
C0OKpkU3oKSrTzqEzd338S5OnkicKu1H7xfX4HjolHRQIWU0yu1l8YoPclGLJtjv
+hvOfHaw7LhwxbrwuBTZuvvlkzvGkorVNiHpc+2BIns80k0mDE5vhpMiNwWECASc
e+lKKpszt9bX6Aj5SBaxykj4FnuQ0ZMDx4ZmtkT9v30tfJC62rM3ojqu8ws831DQ
4folYdFOHdP6kcwC4OH+95v1p1NSTgIEJkcnFG1oyRMHSbWwtLbG2e1vD0BWuPqx
wOtsE/vBfvkbvRi/bMHmeRUEHnUh6c9Qadv4xfkaRNST943QjJxYnmmdx1wyXuwo
A9HwIf7kNLsvfV4z7IJrR4PBI53ugsqJ5wm5/sw2srRJQoqpKucwAXsli4ZCQgbR
cLWOj825lcyInrqKr/pJizjaweeRfJpnXzU/CposP4p1mme8fug1mKVYagjxeIOg
AWOa3A7TDW8OiS2s0Rmr2HpchDA5uk4c0KGr85kI/L7XOcChPiSpd+7OB+fCfPKT
L0O5TcdGAQLQyRe6aAgBDgYF9Q3oSC5CpGGPpX4dlDYS+QyvS2t8useuZ3fkV5Fi
lS4XejkKs7avqWMdULQuUxgPjWy0qXQjG5Llif0LFxSpE1hfjUeLihOOYearGpNu
JYuEYpVGes+cexRSl2pCrvgboYelL3zWDKhvaiKatTYPAZy7nuYnXmCsOOeJU/Q4
IsteH1hW6JMb18W+b7LHn7/rDewJxl4LvMHf1IPhQJ3AVng6GHXZLVXUHF0NgnBJ
c0rcxVZaUyRjrJL4HouLyaN7Cvx9spYXniytAUY3WArIi6fqt5V4zf/sHM6T83Fa
TvBDwPphmfxBd7e0seUzJZPU9hj8/iuqPO1FTw1NvXfJmLbVXM2ptzE90pGtd8ZZ
QR+ChG7PyBGKkEAAPiZWbz6xQEq6LuKKytuz9U7kZnsVUWudey+++66KYUm0OIlj
xluEXZ0H4adANRpw6zHNl6bZXuCqez+x2HbiN9zCCXivt4KCYM0f3GoRbqYrEk76
ZvnC8l33G7eN1MzpIkpgWiMxG4RpxvMnGQMnuupfWIGN3bYQs1267JLxgubsObWb
ybbs9vAmN3wKtY0/smXASn8RkhUpxR6K7eE28WpsPuhDvE1WB3P3zvTOHqRWaxNc
I5i6j0aSgUEOQKTEu/Uhnd5IlZDXeocVUTlMYL9k5h5og84PQ1jgBLMSy/nn6zDV
VrYLxDGsVbwXIUlvVKiwvjrHAumAyBFJUFlXzleEoVZkmzB+tKiKWPEsfGH0QO4c
S1JHj5PjdSMKJFJjViYN8+ZJU52FQXEcGYQlvk6quT65x1IDSLx688Ap8TQWjQdJ
x8KmSlN+8CEXUw5EeUEyunYvJQYjBi8h8NP1un8y/bLmziYxO7yteHYshSKH7zM1
7WM4pcnvQ5tAbbCZa0Uqs/cqDOztTuJUYx//Ga6EtVHjL9dojI/jneXazk+cHVVW
66uH83roL07CCv71ShmY6nGYFf2VERawn2mBXFWWewSyq/KcBvIn6RksVtvPTbtg
eUL5aHL0r34hAsfn5c6/x80vKFTHLbfED+VE4rMPd5KCFHfUfW+eT2Z+xLmspb7a
6n3adMSW9Bnif4zv7nVOfE1SErr4S99zlle0DCuXmeqWCVOUjDrmoEGX6nRzCLkr
/xVoVmobgFd0wlcWzspCZaLyiN9YTzC/rLyk329taUOUMQtD41Sk6ohBk4zk6G3L
bqOUvhpOqwgw30pi7i6ImSk86ZNAeLsA1pIk8eZxt/amsTNWuSE60/GcWqKL3rAu
hhHVnFZHDBwTBYag1btLqNtbeAGEpRClcgorLshMozimM/whIwluIZAO8QNYnCXr
P3XF9kOYTJ/5EzR3/NSO8Y8oYSD9jGyn+uBMgsV1YMsVF7foOS3VkFaWkF45QDuh
i9YdPLR4QOn0irj1n8KQc0kjCOEJ0Lk2FRxi0c/EzhoegS5m0/XOnYtofcAxGYYm
ogpWo1EdBbhpiG0mL+c77e/Wy3vG8FG5eUSN1MgvdWllXBnP0ghJbmaMDfYi4gZ9
i2/QAJam9rlRlsv8mwTMiD+NNa1/QJwZUGQ+aEi+qLzUFo6hqSR6mieOPTypqPTA
bln5i3LCfczEO4Pmoc2Qfkje7srM//MBzXwbMg+JMM9KjiV5aKsG07EzZKPg0RK+
ccsgB+ZmRwqKi02mwfzkyfsiQO1RZJNp9Q9t/Rr/1l0r0JSy4tOhxB9YVnojA2TS
3CDyALSiFHFQIDzhAeFu91J7G225BEexYBnqGQRG6wAavCMeKXbnBGAb8+ANi4+d
s0ToZznjXOIfq4OrFi5ybJMFwxCyDOIPI34s9hp5PdynfdiwVREx6aNaxrKs4yyH
x3siEZmvrNi3I3pNVSxQxswLD1nkmWHXi6RWBtrUuF9Aa1ICSAhun9M1MDWkI4Ol
8hGRL954FGf8K7TBomViaX+RfZMrpOObPIRD5aaLCpQAmrWVP0ZdCdifMQSa+8ts
QCiiLFk5qhPHRai4ChxUN9925oSSOe8z33c/IqwVRf/pdZgGIRdp74iPD140OS0p
0ebYJcbFGCEjD51Myykz+HuTetgFOf4QJ+6xqAumFtWf9D3t7dMKy3ZmhocRsC7m
ntH6x0ueiKq6eUhBbjMUHstxI/fk+ufHR4l4b87Oz9727v80Cnie0C1vmXdOVo3X
s+UhEcMXKI+9ZqjwsENHXymgW7hRMQZbayuYzMgRQrVFnnu5JIGmg3gLIceQhS0u
GSXl/I5/EhvuKeB5JuNOKb88Uz9SR2CFuWOXNNQ9aUUG74TRURXGj1hHRh/f0CT7
KwXGUYubVZ1os6eJhQh3HDaUVgiW6m8kCLvS6Sq75JP1vlb3rbNzT6DrsuWUJX83
+MD4JQC8jzPe9d+xh5q4nzo/zinp1iSof5tuao8dEfigHNpXAsLtKbRXc8enC2xK
3QYKaFZ7SBTV5jyMbwCDms0OwQgGNjTitAPFU+6dUW87K3+2yeMspkPyB9aa8x39
sKxdQ+s8BbfPZJRHZmMV9H/lBRja6Igbc0aeIyR5odcaIQIPsDkJUSBg+Jtrxx/I
2fpKWucpoS2QcVK+49h8gqDFkDui49BrveeZJd7MSl0rRU6391v9dCBKkGMBjpzm
soac3qVMkmquXacZ1mQkpbWJ0vcq5kH3GrE5yKS2lyFSG3RZs1/tU9KGb7j8lx+5
eT3sHmzD+0FXSWfAzm9BtsVDbKd+qXr48Vc4D1312UjMleKVdcr9v7qpVSujOeLH
vQGGm4mWULSmVZs6BW6TupxOcJm1hdhWPippHc0nElgt3OcpIgTpxnB/zwzyvOWQ
RTZPkZnIC5rNtqP5OfyvaR4QEh9h1g1+CfZdc0YONw/qc2Ez744P/BlG4nnRcaXy
unJzbRebU4wHyuNOxd5Uj0IR0rU2EzgG7wtv3F3RSwrp4k5vmWP8WKTj5feAbko8
Mgx43HEKngqkllOQJt7jiLruIGivohS6q5yl1hb58K5FuDO+eOU+dxdluAFI8XCA
Mfr6bL4sCoaxeb0llq1UIER5I8zLwF8y9tsgvaK6fFVpLCWjbMTB0n2WLDIgdLaL
THWwfY5WOs9ovOoXWofHs8QxClwccgyMbB7O3ddxtrajSbDVsB5+WjpSZCZfeqrU
aQd9fpd/8RIDcqux66/Q1ultxp85H+uqW+xztlgeidPlmlVk2BjDVzoZcEqQr6Qd
P4mJaFM4cn6BiGmj+DhdBPBhbED6YySXxGo1lqdc0fm7B4jK4vUym9zo8UsQnIp1
LDRYrgtsSTpFOJJYCiOJxh4BEIcGjeK+mSP74RIX1GctAyvGAIPry1S+/2VhbASD
ylhYtnja/VmtWYn58olE0FYfNeTHFfRYAmjuCTOy6kWyMvHN+9MkYwuGPpSzLcnF
xUpyiQUKDIQQzAP+avoXWXrIBrqgrI07eKah9/bv308sw4QoEl3PzJ80Wzp6dzDv
twGyQJ7Pqsjvtf0phw6yjhhUuK43OJspOF/SVJ7N1oJB4fgbYNGWTwNGmQB6bmDR
J5dxhhHbV7z5EV9eTQexkfqiO2RcqrbJqoCwDd6sw6JJPJmePLImg9zpn5ILimxp
rB7KNdOYqIxf0kftkr0/FJrUgYCjTzsuyvxgMiK/ESg6HwpQaOzyRsIfh0MobOER
t5Ll4bhQPIxIVDN+jrhF5Cy9S4mrF018kY2LItQl3w0aQvXQ00HLPt0ktjkuwn/3
uSKb7wIKGM8g5ONvkFVsgSz5nnm5mXP507mzUoqIWns8heOB2Sbr7U3XUdRuoqaR
hVcwvUyvj2pBUaIpKMRH1l6CT4mY1UOVA7igeDFCzMj0n3aJfyBeJozh3DsjDnnU
DxrBCgN2ACJSuoFkVmgcoKL4IBxVSrhA8XbV9/CFyymsVH7OEw+kKSnKbQ6z4II1
PDifePunizV/ygDil0BlXP83U59cwGQYSZw0fgzhDSnVXZydh9qdI0x4uJ5krSob
TGX9NXY5e0GsgngTtYflaSSMbeC9+IuCwM3x7uW3kJnw218eK2/egxDgaVI/mbO8
1WWLcYLn96T6BpLW+c6mOO259mbI6ppASd61MfmSj8Y8oTAKzejq6bi/aqq0H1PK
vlrAizYqkMmVyS+Tv+YN3VLj59rXBxkf4pEr8qUYC+TG5gB/gQnX/vuLklyCsRzt
F5AfH7vJEyVRlcbm/T3jDXSaTGBRULEnNVuT7L6h6bKhyNHiRSHEqmfTFRVlrWmR
MSVrkdOU7Kwilt1vsc1+FfZpn7LMPnqVu1XZEL30xjw4YL+ym/xw+rJgy4UdV61n
djIdGQ07rXMH6B2d/MrWZDbxCB4060nuBQL2agvIbtfXabrepnUC9A9CdVf0zXhi
BO7iWszvwrpAwzu4US752tJcXM68rPyyFCLHXS5n7GrDjn5H87OFZsST8wvk6/s+
A+YmbHzf54eLf0rx6QeaopYqiSuFNOPZpQYvTnONoKrX0B6FULijWvJbHXVWv+Tp
SwTtAcrWBi8CoeEQRqG9/S4MGmAoOYnFJn7ZM9CYKwAYXSk9Y66qj3UivYh1Iyus
pOojs91+nMBnR0GIyDau/acOqoqN4NuqbybYY2LLvC08ipb8+i7lyqaTt/juRRA8
2BP127FSWtVW8zqfDAeNBrTwqZcPKU6c4oAkwNlVvfIUtT1OewbLnf556XFWvNfl
b9BGNp4fPGNyj0+xFZQufSWt60ga0+tHfjyrkX5zolAS7cGEHKtPv7KQnxzwkDmw
xl+KkSN8kFda5+0+PBbWgZu01VXcTdxUKrL1RTKLADdGAClwApPosgp8H9hl5ArU
XBe0ugZoT5saU0DvD7ZyWWc4kgGmJWJbaNsbzctD+53au+Qii6wIpZ/2dvLB1LNU
HYQ7xNIBfWd4eQ0C33F69nHITnEv4q1tuZcuIfGYq9bCTDYAdb9GZlx4JJ9PaRSc
C1SUFPP69wFo3Z/K0EqjYM61120NV1ObNU00omcwptvhnzRUZNcAo+OMDd5xnemq
kYcLzqLKU5TAjSjRDvqMNgQpz4rkCXMA/vnQmRFtEnTscDABGvXfKTpp8GIAsxu8
/7uk7ZsH2M69gcNXEKMyMqCnnyrNtPYfOqf5iMOgKnKACAlAVz0s+pXaFXNfEBol
wOojh14zXdEtyrR+boEnHKv33pmOAFuYbRhZrOO6XTUJYbReHJlH/d5hj1Wr7T+d
yzO/v8IZgttCYXbzTRFbwr26Di3wY9425AdRiERrNdSYtazjyW6vrKgLaYqAumb7
vDM/renJLiBRoFcfTpx1SaVqRqbvCcyYyuI9pudLfsWlAjMAF3cIxvoOsTo0vD9g
i62rCW5yRVmZtUtXFMN3Yo++R4PPVPin7/+4WxBifiWHSalFYaJPmxnkKn6l8LOx
+bXgIA5ACvRloM+CYqXst2i6jftIjQuYoUOOcQMHgVgtDMOVtp7BSxffRsERaT13
aPpUsnLHQyDu0Gb4A0qNs8A8wNW9qqCThUTIFiLlLVbvkIuBIKV/XC8yB/AzgU7T
ybk05OaOFlg9BC9ny0ZyX9z+bptbGH7iVaIS+6GXTMALJQEShJWQt/6AfMlJnGbh
vcDgT0CU64e8DLpEaXr+f+V7ZSb6dvPDbxNr77qorqMQ7cgmoXIK8GNaCUvAW0IJ
aACcuKNQzKmiCAzewpE0P3zEu0lxAWPeRh/iXZmkWXh1SVqKBoB6G0a1KvWPtXPG
hnPNoKuRB+ELh43U1o0tlIuDn2kFGKxAXAXRkJ+qsErtuG867/bNl1+GxRpYHkv9
55JDo+mZ8Pllzo07ZORLvQ/JlzFMASiHapC+HDKM1WdKZ9IcHnHuuvITb7BSIY3a
qOIpgjvULGECV5tVMHZ3FfjVIjRdOwgMJPXRKhsqW6ZGDsE7es7ocQmhVu74bZdh
t/rhiHhXXZeuAxzlzkSanbClLm12z5kmGX+R/lwxQFv1xrf7+yKZnjwW+MfddCqg
aTnDf9Sm/KeZL2p8fmZOykQ9s6K3wvoiapJDYtLusfea3y93AQEiuTfFGKr+dfQb
ouqkkMRGHruKg4FlQVtGszDGrWs1Nz8fkFn+0aBdPYSH1o74H0FC8FsTvzBW8Dfd
tuw+SNAkZdxXMixKLXTWN39tH5jrE6hBA5rdxcUH03Mwnh494CjKvLJLnfdw45r1
XOIzRryG409dC6ZN5GrY/LWX83TP47Dcx3dgE3P/GUOynbFh63N8WZ+ekani8dfa
Uf9gPIFFrKaSYYunyWR28k8fc6RvMvJCRhtH+RbkORvuYDSuE3hd+fO/2+Q+DagL
vhXweootfdCVwofrI0lC+WfGp1r/AL8ZXvFGrzi87GX1uiZCDXaAp0TleTlFZ0QG
uo+Tfq8Ljrv42xNE1cNdXn7GLtOTVT3J33Tg8ENilqkUyH3N+wFRTc02QrFAWWxg
SGCuF3OuEOb0LdMDV7vCGrDvgolO2j5hcH+Zt/qEzzCRv4RfL83G7uDu486GnJsx
cwfJv43sZLv3Z+XAimUglZBUPA28pWD6RjCiMXlHNIS0m+zMaJsmFs9lwrgTOPl6
ARBpgTYkwYMRzTfZ6rbqHt5Rv4VkEu0hkMTJ9oTlvhbC2EMptwv++Kw+pDTZIoEX
ON1XdnwqJwL6EJlDGFcJ03VSxTvEzOh3AxCZHpj2cGV/pz1R5YvSIylnE0PDQYYI
DXYIYa1w96Ey8oabLBZOMgnoCp83sI2uNOv1Ts0OvSDaRFE8uJ/rHAVzjd63sTJa
i5jxg1qvSCqAGqJmHBkstQd01BrLJATfScYyqljsQsLc02EsGWVkWt+GWAsNEvFY
7qKg10njYA+ujzAzvXepuZVHGWrrLkFxKeQVcf72+v6YTItH7GEYwCa7VuNhTnOS
pi6/KixYsJxKeI3E0oiIAecI/XC9mgjZlPjQnRcVUYaS3DYrrvL9HqzZz8nIAc8M
TnMWgc5/za+YQkRbyskUmcmHJ07eNJ9xeedfIubVl03AuJB9Ui5+zjNtIqtYg/is
Ex3fjPC0sBFrTmn839B/n2zeSDXfNvZxr36zHaIRAHKEbn+bgVnTldHmiJdawqf9
GYWI+QY9AxY6uue2oG+IKlJl9BBqzs/aWtMV75ORYwmXL8yiqhNxSlMpYMPnOnoO
V8ddPTqExvn5VhNP3mXF9D1wzLbxwEuL8ly0cF7Kmfe6yBI1AYDm35IY+agJ6zxz
wtlH53jAQnhFKnuLdtspZ5kAr8FAJrUDGhoBHOt7/+ioLnMrcrp4Nz5FJ5VYy82f
76z1urMQZw4t7g4TBnYZx37ooavTH2SOHJNJHyvwniDBdqWcPNXoIfDzqqF2x/Ve
rQrefWFoyue42xIjWUQ+95Ofcd4mlypITJi3CGFEB/vqE2I5QYoPKdvgfHQUJSbP
EaXnyCtsxf1urpM+MxWZBDeSQDo3CbbuJvlz8TM2tiCJvIqgvpaJWiNcM0LF30HH
SzJ+GVNom2gYM5ZHfJ5opjAEt4kuHNlEGvlMUpv/njYzPx/SPbSsH5QMO68tEjXr
3zxkykwKE/+SNpoRpgm9+UQA4HlfXaGa+yPyu6t+/J+K6AIy4wleq8BAn/gloG2J
SW8k8pSs5Rd9WUmsxbZsg2evMoEGjxXcTG73+HwQ8ioijlbAKc+NzYK0EqKi9PPM
CtCrrXx+X1YvBZ6emjtHSlmEztTzTUF/zWpkd0CVvnhCDlEUJe5SKdCJ9jRV6Pm8
vlpYU/tyEfVB+IlUCz/CN28LMnc1tYIngmYaAimI+6fYJFWbvFDCDxoq3NbYF6r/
4QdGK2pAAb/l/eZ7DyYfuWXk1DwK+h+AL344HlphqkDFc6OYavIEDocGwCR4UEQj
QenI0j/WXXlcbyLLJ8hWcZQ3pM6S4GGtHB0lhVsBKmdVD2dtgQaKN4NYqNN6KWcA
DbblgEjyECwPM6Nbki3oVoo0Oq5zV4LMtjaFtlGTw/p+9AURC8iIwktFmt8MxYzy
ihrvNdm1Dd2IFMVFIS31cg7WVajmAZ8TsFFnGmGqdQAtmhWj9LjPHHyWkVdyP/CE
ZEz+0grciViynhWN2QLd3wbxdvdzJw4X/VjCGtpxFnPbpWJQFjJcpUGVj96r7g1v
MHl1YLO2H5OVZ33POT+DEXdqJe4vCVTNO9z5djVhJPamXLblQtX3lKfBCFDKe7D7
rJ4gGn+X28S4NAt4iziXmBykec0XWJujuNR9MA5WnK8wQCNgYzlH0ZWQq2Mpnpco
DZxwrL64gOQg8Xsya5pQpp+cFBKQMyhGqeTJlFJ3lDk9B/u0ccoZ8iw+hszwFZ6p
w602jlh0C7l9NOSW3o+gSvugcgfElMl+4mBrJD5/NZdFEjblVIYGDDakUCL5tHbU
Gkf8Os5cdqGJrNShY5UEyJpFyuBQnPi2bG/YtAcIkFP2c/F0OY4QVD8bho6E3ptg
PczDqw/HxSxiKu/Ol6PNPEivye4c86QTjSd/Tf3qzkmxxNHwOW8M3vcYZXqqR1lE
+9T6yIsSBhDutiVDi2zZbD0JWRuiZyDgBOXE20hYtoH8NH3Y/M3WCjdgr3Ki33po
Oc2LxzmUAaQOW7h5M0QM5K3zzmxh+l7rUPAsrF+1Am50v0gDMGMf3vgvcNFuI+YR
AJmGOvGaXP1tIxxK4CH2qvGtIa7I0ehOgn4Fx6bHaSd4/g34OHcxr87CDBcu3x+g
jvPpOdxq9C8QRTU1UCUIRt0YTl837qeNjZRRPutNeomAYpzN+8ySef0Y5d2mH5YZ
D65CCwx2jtm17GZn1ecIU7VUi5JCrDDm3eIgTJvhvqKv1sMvQBtTz8kHCRf6SBgh
r2BfZ/CVByfytZZNcnEFJEWBuB4wFnrlaFMNGvqyn5bwQAdccDSx8j2xcxYjXvO+
iX/p34Qv5+NuqKcLczmoe8YKYue7QmQtOx4yNrL4c5JLJ0izzEXcQdARB95GvqtR
J5R9yVdP4WFw6L02CD3FymfhNawN4LH8NJPvEXuYpiOxrAeWjYohdPo/ZcbL/rRa
cFIDEo+MXZ7/aiYFSQRlRJ4pnRoxSGLx6pCrpmP4cnZXOnUI1nywqByjvSRI9XfS
cqw2KkX0XttoRN2oRHQh7gBLMF3DYoKnNt0kt3WZpYUspmPNjD+iDnxXwbBE2BcF
JMO37JR6oXCDlxSPdGxtFs+Gtw+PPY3IftBa5Pi2L2Gv2TfwHvNHemon/1SV/yeY
eyjur5/s8P6ceMJagQV23w61Qm2kWKtf2iMniePdcBjebCqNCFKd2qli3UAgd2Jj
LEz+aXWoBoT258ewXEfN3zR14WQwHdtibeVJzyobatMZWf2gZWgb/c9xz6eFIp20
12DbUzEBuGRsjuxJSkaPd4PtGdoIft0HLfCd5p5CHNLdaJUMpCFbXWtyIcjy2YvK
IylXBR/QNMWEN/Pi5AhGbqVp2HCMg4yrJZwBVj/NHKeCXCH8mT1sjyH0URbsw2oY
N9UdxL4KJ0/0PVcALj+H1MKmr4YqEwwA7xYRWAWgkK6XKLgMZQHv5w/rpsmhmhPw
uUSMM/sy40EVgTYx0mZnTqOieyvTV8Sgkh0GWlaSctIfNlvNLJ5Zk8EOCl1K3p/R
rdi96zPALw8IJ16Yjg4zZpdvk3eHx4KgpERD1MujOXHwLi/TQjuZYpdSEAywRu21
/lDoWsLkqHrD71zo3aMzS4vnNbysT9qglSw7Ik8mBzADEz9IdakiIxlFpY17NEgX
MMwbJw43PgUVkBtEB+4PGS5MJj52OvPmeSUavW93K/xFXR0ynpV4/ItPTJ53eTQs
3aXR1pgTLjBRlG+pJlgPa0q59tjR32zGup9D8AYAW9JUOsNjQB9PryIGHCa0ySSq
hKQdvgUh9bdsbwJhTtjJnSrd2fKguXIUP0SRxHPoaSa63oZ361x7lsIKDjKjAPCR
bgcUGwt4hkzvfOwN99LVg/C7F8dHbOTWB59hYVCv3pPNGtZEw0pPyZ3Aaok57D4z
mhpuUqVsXpLhEH40rhpE9gFo0EiPf0gvBsMhfTHrRKD3Sk8FdrgM6uQgN+MzZVlU
KkhGzCH6MPKuDduItHi+5rHbl+AEZFQ44LMveW1O7O4F3UYh8hj7/gVrUUq1w0NY
7KyGWUgirOhKsGcIWJs2etIptp5oOVZ+bJ49zJtvLNLAgUNNXe2wjz2INvaUAgQN
kshPE8+WFLAvZtfcPdLmCZvIXcWMLkgSUPX2hlDwB6EMGybrf3rK1n8DNkeZLZSW
1frBoRwhVgbNdEkUspy5bwmwolM+GPbTEDAdRv6PoD9wZA/peAF+/nY7qDeXmb4v
i3IxrD8Zo7Ehlpv1cCN+REGml2U+cPtukAqM2U3OCY7TKQzYss1p1oMsc2GiyPzw
gxqOL59Nc/YTra8Lm2QU+IkpI7cJreuY1Z/gA3gs6FtvuczipBpyNVe53/VPVIe5
UaB8CBXcRJ3UbzH20TBlgC4TLZgcC4qoENJbAwtTKSM4ei2OoYADB0Dfw+LiET+D
E9jdtmXpx8EGtXH/mWbYnO+G6DnI6t6gy5AZIPnFPhCdrX8R3iuzkY09NjvYVh0T
a0nnre375lQ+kqGOsV31mRejSZRgMAsMNP4M0qvsam22nMzzGD5CeY8On9NI036S
IX4g//4Awzaf+9jorKZm8Le0RM0Hlebha6rqnYk87O8QXSE8vebQv9Kf/e6qmoba
rFQoO+Un1ewGga83DcxQBzoy6zm0OkzsY3mzLht8bqYaTfOy0HU1ahm8IMmkH1uM
ZeFSFMo9gX+6L32jZpqU06LPQIidZ2enIUUOZgOJp9xEwbEG2c+S/OQQN4jpkRpQ
x8lrdgs0+i9oGy2xzNj4iswY6o0vt46x3ApOO5cOi1guBqklTLrEWFkILBzd0zr4
ny/mfmVUtOs3txL7z5UeEfO45oIjETYX9HmsfMZ/4q2bXl2sBUDe8Zkf5onjyk/3
5/n+t8JPs0pDZ5pYQDLziRqw3jOAZiqBpcW+HDXx+hv1qdyw7c2vbaF9xeOpVXjm
4IbV9e7iBalBYhPOR8hJP4nlfDuzmX/+DVobEJVK6FatX96rAPwfPyR3zrZ6anLj
eN0Vl5re62maUFFi9kUc08NUfxFLXFps4jdfPye4ct6OngkYbDP1V/h0e4KBr6ej
9PNbNO0jmynKUKCE5naDPD56EtNLF+tDT0qFRrYPetLvtluOzvbSokhDtjnB47d2
dshjTVfmHEwIM+z78KvlcFUOtOEZBIvOYrtKiIRoBrALBEgrZnJqTNb8ZNqEx0E2
U27NiTKm1V7CqMBea0BwXtUP3NGWIUc1rV5Ty1MvFlOctUREjeBCDP0/ddmWOdRx
+j9VbF3VhTTfo2Z/jTrFRuTP6GkdQkpBeQjDS9PGPbQW6zR9iclOaXVzCPRm4+Kq
njmbE1JqQxDQguRBy84ehh6ONgEFYxVp3Sr4amrbmkAg956IUd3chNbBNayoCmvv
F4tWpEnnW43WyZ4+7cs/89O/+DdkBeKINvJS8lYZtcCY0wiGzzCK2Ax2e7gxKi68
0Pz8MYQ/DXLY2BGzggHdsq9hX4MEzU/4RZIkbybdU4M6bB3ty8utBxVF8vvzB8Uh
SWYtZsRyveNT0dXibLRFFH/9Dtv7DyNwPNrzhj485GUQzCv9l6FbIs6yIndPrsaP
AW6Y8Sb09touiTER5ELT5Gq2UkH3G5SG5hb9uyvQfGohV/4Y0LyLi8wqWMS6YERq
Xkd7sePJlhzHRWwNturisg==
`protect END_PROTECTED
