`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gu3195z/UMHJXtH9Lai7A5pJXObyq2QROxofdgHUwYgA/Wn89uAPJN/Sv0Xgc6pr
e+wRnoGO02Esdc8yOAnDUakZLX/qbL+6EfinlFxrm/CfHg4CHFWjL9X85dJvyNs+
JBiTM/EcnzkK52M3tswRlEE3gej3izdbZ99Vg41AVWI1b1fsQciWpCILNb0XSEx0
RGWd7sHJmtiTaKlrDzrVy/G+LWRGJ0qKb/YUoqoOM1+r/FmRaSjHbKNm5/k11x4k
bSiKSXWFahqPfobaHxh3nsUv26MfrCswIx3+dsrDt7gWnQY2XVvkur4KV+DbobeL
gocRZCorAQdXKWtoXCq/zRSpG3a3MzS9tf6eKLNoM9UeSgdggWwVWzm7JlpM/+1S
isPih9NsGkw+wbGYfMg45HwJ7rejBo+rLycUHxb52uLN/zk2gP2Fe9o7phWBdLiC
4Xwr5utgYqvo3YOllIB+xWaDYFcuitWC3Ok8OmAfWCeTFJLgwKm3Cecai/B7vro2
KM4Tr6k3iDpv4+Jj5AUidx3P5ISuuAPiYDfVItfpTh2D958k6qoy/1qHCTSef+c7
t6gmZ+9IJqsn0sIT7cIuSH6sbb0tqSuPyOLqXD2V6ZIEAPxBv8BLeckNAAQ3uYh6
mDm8VgT2YlIuv7yF3s5G28vqkr9iHnQSO682/NychJL8jZUOyaB04rLu3j/GHEID
OOeXutKYOJgD3kbuIOA/vFazWoKOvGHuWCDmqALvHlt0BIpJzENMEFRTgIMCJNbx
NbL80wajdE5nUCYs457RisYxcXJhWF11zz+pHk8SNjAeA9wor3ZYOXkW8OKwMW3Y
mZ2IOCPqsLLYGn1Ziwx30R/g1UdDubNqKfh5nvV7Kq9edzWHT4ZTAXcRllkISPzC
jW0D9cUrA70JXjlfv1EQ2p8Tz6/H965eAXKizDPBDkHNdLfacBGCNlwYUTSvGa69
jWE3GwR88lP51bLGen9wROCVl8OoHEk+PRCB/LqprRNFqDGabTd8ez9JjDnyZGRB
JAx9IOO8iBefOeq8U4wv7upVFwYJ+FmiMn09owuD1x/O91ksqQe3bqNPIBGBTaQ8
DWRopHpE08TbTrUpj3GjN0S+S/+JuzOhwMNzm5CWbX1B5yOrFsLYnNiMHvh0cs3G
3J7jZus3jlzh//WV6P3y4HsaTXTdPpfxuyrK6mJKFxEoByIaUvgIkCgsLCd5ZsYM
Xj1+OTJkf3lLTjFdFENaUUDRWB3Rx6YjDaAGW/EqD5KpfKDOv35W8NadPegDPO9J
whFfwAa29lCD5jm6aid6tFPI9Y47/JAfeCH+/k32mv1K0DogzfKRs1o+5jWJMPj4
sU1/+bt/2VB2Siu/PqVqLFDZ2QwGEiOOtjMI1csELf59m3Swd4SEsgGfHAUZBiIL
l0Ovx6oTery44NxB57NCXja1ycOw7jKcI40t9eO0Hh1XHWB266DBs+QGajbjelfU
L7aG3USjGxKoaxGoAkhW7awf2sj4Ub8l1pyLi6y7ufGhXPHGmQD8h+0zSKjCuUMY
dOrK148rwl3VqXebwTKJs3UZ7jb/QT00R7z3hJglinEE6xOwLL5Z7lCxzIn8Va1s
xLES48w9fBaIeu4qXcPHOpui9rdzvfmYQ8/DqUS7t62+jLI2j+2vE4I5bmhjd2wr
lS8/rWHlaVRWWNZ49qlUXOcFTmn9i+x0ELmNWDv5I1HTJcHyWPhOslRtBAcXFqp0
7LLl8AuGwydteyv7qo7OFOArd/wFYIkWORa9VSEXpiPxGMLEKTQ18brx7KBAYqug
F7OYJai9Ima7gu3gGZ4cLm3JJHdDlIOltb7nYLeHHQqqooJs8xoZWzNQnSpajmbm
x4dsICeHyMneeJfbJhzhlNMPVAlrb3JgKA+y1nwJGV6dtbhn6EhzqvLq5kP2w1NC
UOw1ZSsvMRI7tYf7H0DDe2IZpp6x9yemaDDE02Y4cbFRrUzjMKXaZy1Y9yJBrcEd
w+XnqrWEpz/acTEUrwQgTLiBHErJ9ChHtDQT8iF02q03gUUcTXxOnka8E6R8QjDv
Dc1/qJan3bonrSDfeYBJ2v3cho5kOy0XUUeqVpyaevJKwhq/giaVPfuLl4Eyn7kE
xV6usTECbJm0lrHFomNUEjOfcUcrkMlDXk6iio8Stl4wZ17vNTtnxrE5O3iSeOdp
AGAlgL6YlZqDnI01DccHNuLkqq523YyTVqtlU8RTci+fyX58Vc/627M2neALrw8r
dJqu1/Da050jrULPkuiGWyf5iHpj/k6jCxT1bmQmSFNtzLdaN81IogC3ECenaEZJ
`protect END_PROTECTED
