`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihFj+st2vl4+SsnUxMUz0tmrHLUgmeAUIBzxy+dwMgb+rt5W5OdaHTeNYUyhkZQ3
jup8y5HsBzo2dRO6KQKoMuwxzxkdW8dEHNADIAsp1oXmxahu3qho3XD3w4vfBgui
DelIgXQFda8vtAkczcA9XFjN9DOHmEjOSAdmyKzEb2EMaT+BhN3rY8ul2Gxf/rEx
s/doJr1w7oxeoHeQhHg2trwYRJkyUnLk9153jXIRCIxFdjQv6V9cJAdAUVTIW1hn
5HDeHhUgmlw/qHcxsM65O4wJ/Z0clRttcN9gTju8EolUIQIZIx4CDzL96Meyghhj
kh+v2ArDqb37LixQy3zGOPLY4cMXy8nqZkSkVvlzqVylfomlrED55LPfxiiytm9C
bSZ2Nq+cToxQUYpV3Rj0SCkJj9tJGaSB7rlFO1+Degd5oMnzR+aNe6mzwP/b0VgZ
gOMAwvSqlXqo8TY6j9Bj4ayQXQW4wvpYY8u44jd7yCUVcXRakR4YiSEMxQgR7aVC
U4ekU0A/9b07i/8VSwDe2niD+xwPh5XgLmi3tlhp7mTiMHS7bfs/Ynu3AMolHlVB
R92eqAozkxO2j2MwvA4C5syWnfA9SZdr310O8UzUE8vU+iIMflA3/JB6s1rjlgNB
HzEQsOXUlN6xtlNYx8juW79eJmnvjy20MbPMpeLwoH6w4/tddFC1ImASyESNmtwa
0dgkVyBgcyXTfEaftSNEvw==
`protect END_PROTECTED
