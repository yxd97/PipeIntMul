`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sN92Pbbkguv5zff+nKnuJ0Q9dv49WRdvxGLpNYGGI52tmZt9IeJ80UutaMWPSz4a
JufkxYYUZlBziE8E3sZxVSEYhzzSNMvM9AdrnQ/jQeGZKVIS3S+p0zXt6u7Nr1Wl
bZxy7qbmBixMH3wR4g7z19HxiBn6xFJOCdl4oeQg1jPvHbWbKJXOHlGJ8Uo6a95I
yP/DrLPgrceaVUDpfeHjPKIXPaTwLQHtkcvtru4NnEZ7ESBQUzAveKrNX7EIWKGn
LoAV65QpRp/7kwk6BOcgW8jounIBRGQvQgFwA9GBkY1XMT9Q+6KaVwl92td82FVR
Jgn3pn3mgxxvLFFplb7H0V+lnRxBrHkWKJYyhq6ydtkXDsgtzgXnAQFki5Zwxz11
akJABSxuvJvDIP4bS7QsZSXUMTY6sDoZoXQ53K9193BHLem9J7QBqI0vJoAZfCrv
dSldbYedCSoyQtTOppnKDzkptEXM4T+i7YQ6akAM+9+pzOo0YffXFw0SrVghznDI
X1jKw1qsjEKbjZCHB5/e/cib43erxC6+d6vtTnL12UzYyzIC0IFyG10RfkZJ20kj
L+vRiBGlwRlk1qF2xmikELylxL7dCw6P8vGr4yT03AyVtrGzaFnEuxHnYh41Uv95
eAqsfO6dr1j7mL8jflcUy0HD3BlzyujJukm++JkxVdzv8YypTsqKJZwHbGcaJNsK
RQYBIXtP/whZFE2M/VXTL1z4WR68raP3XiAs6QsONdTppk8T2eF+Wj5kg4e5ujQx
PH07UDGQZU2YYNTeb3dsc+v8WisAx/WQ5qIxVs0zfdEsaZB4Ax1HHH5w2xMLWfFp
2Qw2uBT42O0KvXhzccRxxOu3pstQFltm1bbAQx70uYQ=
`protect END_PROTECTED
