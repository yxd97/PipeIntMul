`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSYCXx1Ive6p4yprqCK4jCQdgUC8vgtCebbATy4SbrrcqTJxGUF3tfzyKO9JgU50
07GKIiC5yeJEjb8WPFI1Rw8LvyM9b12O4wxiZj2V91iFxRFG2/v1T2H+s41dvGYa
3LrmQM4iSBMm2nrUXGcLRhyB9V6zsddu571Lf3GZc8FPhPh6V2TnxjhhN4NgIOcE
eYNAvGNQmRb+DcM7I8cD9aIcq4TM7CVA0txBE6fn6aJ0YXIHkoXaVcSEox38QDa4
SsgEkiPO5nH3uSZd/V/rwvu980vOBw/Vg4La8VptCW80GSGX0jANmVEwJVCp5iMD
nNRoSv93mYyb3AwhEbzbndVxBDIRXAEHuzGUF8a/laSh1hmUsS7Htw5daGiYolVr
z/my6PI/HXbKR6pH3G4jPG09MISvWBU5e8Qfi/lXqPtsYZDszL9DE5pAiWy9Twtg
fbFobDtSVN/E4W3NpbyZIh/0bDzNL7PAhBxtbCehZP9fpRXv3M6EFb+KzCnd0yI2
FUP0olPdxlF5Kxlvx6qCBNREbOr/41vcnxEDdeZj/cDRY8Ija57UQlnwzDkcXzJr
cecAEo38A6g24qfDnJP5+OTgclq3RGzyVNLbPYa1iAZayISs+A5nH8jC6H3R6+Rb
jD1PsrROkNUxOk3PPIghC6D1hBQmOCwMTDgVll7M2LqIzxG4yUiYxhRGyNIzglDd
gylN/5GI8FRX5qkT/ykzPhH+aXvdqxv9Qhr35j2jnXLtMz/ZvLThGL7voEi9txg3
mGOOX/T3KsBG7ZXMp1jvjV2EMZGhui8174ZCDIpf8PnYiksj4+cbNlaZ9VIequys
T/8Yy+qyeKtpyu3z3bnBj+tFfK7Prh4tuBWlJLYwSwWOrdEZVglc8mFWqJ2QcMLS
KJ/Q04l8i4lgi6sjcU7rzxwPCMO9Z6ZMPJmBBehCNAVnL0Go6GkQ6wxV0c4cGZM2
uxb0bHddN2znb6gJ602CPeSHVW8LaMoVXsw9SvJMx3KoimbhfOawX2PNocYcDO1Y
UOZgJ1a7yLQFsJeue8dT7heq8R9pM0+0WLNR0A3OYGMa1M9TR0NJ49E7EyB+mf17
z3M8qT7mrMbFHIrO7kVIn3Hrr4H9Hh+gvqby2rnb45cHZL9cI+dgpwqz1Rta/8Es
`protect END_PROTECTED
