`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3rJ6J22gpfGn/ERm6/arkBCgzluIsBC0/kh95EaLbHIooKWwPo3+umTFw0GGCjH
jlElQ0vatKMt6GO6zybRccOKLYrYZb3nd0+sX8sh6DntqqB9f/JoXKIEB1hpcTwr
LKoyw+xuga2DeavHf4JAN3S0XnuFkzYxIMbp/9pU/PdK9oD+hczvHocHqLEfUJce
l1cb81oAsnvfvKplxlh2qxJI/zt3c3KRtK8Z3+vTwW6HRGwQfNZlEILzBGL67frn
goLD3LI9lsvYiPATDrQBWbtcXvnYQIn2qJjAagmCwnQ2MFa4vxqnnnlhNvBjdwhA
Htx9AiPyS5exCUWb7qjpb1sfFYHKeDT2vcACH/+M0rR2UTAFuzWjU1eVV4Jjdwnv
TrnctryqU0mAMamtmdvQqpMqZ+Nn7C6bCaI3p8JOcUEGNJoLTgn7RxbA0aTBrcqR
MrBJkh3dqMa7Q0tM1OcdZqGtPG+bNNRrPk+szUElKPnvNAkylZkjBBEf9LSY+7d9
bOITGGeTf4iwPhsv8dCtqfNyAnMTSkfPDSoJeQeOgSQMrbJMWNBI5R00PU2TM/ji
5olN6kyen0EhAbbpvf02J8tNytc4ww05WLR6cVakLwKgiON+HxCF/zKEtYzT50Zn
WO57rwEcmEnFyabRi2wBjxlD2sSEbxCIImI2bja3tfzv/c//fzPhj0eQS9Cw+6d9
gt3R9pWRMEteRRtzD4gwV/wCUJPEbtE8GhZ6SeLy4Ct9itqzBbzj7mCF6xDt27Yu
qjNRGSaN5Hui8rqVsYhHKlHdT7zPVPN/7ixJexBtEBk=
`protect END_PROTECTED
