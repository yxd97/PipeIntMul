`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XPYawf/xDXevaabMXWF6ZAluh8UwDKi1EKdHp6BQbNLFzvJcvcKPpWAp9uoi0mjr
n0rwQo9kzeJ5cDgMS7BWqRSVa5UPHDEoDg5A9pkQgMhNihOFPFuaVGCgCUzqYw57
pF4uveHLKdTj0BvpvVzhjVmeO/JtrcN+e7nVWS5i2diTEYSmo0b+fjR49Xt2z1gA
c42sTkfKcJZ0ETPBT0PrPVp5nhMoTYYi/ztgadmX3WPYC2YBKdwKpRw+5ra8sVEq
Cb21PVhVMFtqNKR6ZdSMLwaAR2XSgNfGMqPxG4aVkQY7RNlU3SVGpluZfWIF06yd
4H4EVoFUQzh7wELfUDdvwZ4EFHrogxA2sVfn5pNyvXaKt/BOrjS0ynomqaC0ZgZp
CqyFGAWNHgjLmvi1cvZeCXfn9fF2Lc+TLzZhoAefr57zfg+IreyCSR40R9Ec7kFC
UJ17skSFb2wLoErri+NKkT+Db1aB+byDLx3yAr/HFbjZDXpVcWly0OqpAlaFayEM
kC4uCkuvaNaOxlgIjJ4JpmMJfHJWIG/AXng3dhSlYQhUOC35XC94AMNe/Gw21utv
9rO/vqfGspOGeSTKzjksT71vC6BWzQjEDN0xqtu48nrEGISrCKk2mLykofKOaAFl
`protect END_PROTECTED
