`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y88UXhV7rs+TzIYqZsbGJTGWat6KJmqc3Fi3JbS64DMDdM/YxDFS+OL0cCotgipE
faevtKxiJ0RcDIOm/mcdp2J7z6k6nv0uftQs0E5CM3e6eJQydwyW9ncp7mCGkMVD
swPn+znp37e+XfpOFkP9dZ/yi23WEgI92UnSPInGCwnHP2mP7crMIZpn42UDqI30
a9dqF5XazmQ8Eh1igNeptuWixBBtloLHJess9MrG5SCPlITafcMwgreDWShqYhWb
q8MGEUkp437Q0aUshV9zvy9egUvjYYCwRGZ1SqvMq13oft1GClUzmbXdtusWBhrx
lWc5lM5O8DdKoApPiUcMCFuSr5CJybGk0PofO66y/lnCHzJv6z0slSiPGoWcLtpp
qor57Yc/MgiKXWBKOmSuzCi3BYxRfYguEABhkWRIYUs7XAhSlpEEG9Oc7vGHhKUF
j2xS3z2KsSHz8oKyduDsbGIy40+6VSNb2xIqJfDT5cFQkeM5xx3e9EzpWB2GUQNP
owLWW/arZDnW5TfLe4DttkgoH6flOzdASmnr184SaJA=
`protect END_PROTECTED
