`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4ZFapukKavigK69H3ROlqEWEkYXI54QKyHFI0FdlPluUCxrXsxQiFN0fY0/nlhC
1a28UIgzV00YTV3sp4Md4LyEdsotjbExcLx3ihtX7edlWa5TqTUoqHrsI3mqaPyx
awk1qW46OR6AsqjiQTy243iRvdHr0UZeXYD+3amutdYi7OIbD5Mx8gxkek+hdH2Z
LuRdK0SZfNeD0FPPgQ8vowitWQg2fWhsXuIR4c9FYucpfcPmCDe/pNXWh1vPLvvW
AMh1w39cO6Id3PJNTwYLrptJ3vxelv1dt/adISh4oM7wnR0rmq08j/46Qn43q79N
B5xBScaR3pXztJNby2PnWM/Fyytz4F5Y+I6mApNjPMk5UHFQrK4iDL7zTDM2uWIl
uloNhJyRHbfMVRWd1M5aS+dubhI04JfGPmDlj9YRpj//i4gfJt3bnCB21P6wj79Y
XWcHSh1Wx9U7NF4C6dbSDWH/qunnGzLdnsBVkWR23Ne5nK6Rf2f3cDRhF3N2LkDf
CFf91fBpf5RUIxcFTmdaXU36exlK599HtgTN8DHVePHEyQK11UaEXzUIJxRB8WSX
ZvfM9oGfWULgUDEpbYwjue5hss0D+/7b5jEKbOj6DYIbVYaebjdpfwcmRC4NM9wH
kXuLwOw1vYBFK6WjOLGvN074/5EbY+j1NZ8aeCv1Sp0K13Pwys/cFrBepA/jZ6A9
H3HNAsY5QUZcvAmLsQ7mvIV6ShO999KGJmelfp/hsyZEjCHEWwKb/v0e8cgGPCkX
xxSnQmCMxL9koZs9M8xxFtZQGc0Sko/PrHehqnu/66CO/KflOaHFESluICnY2/Fz
LHrjtPd6iJ5pjPwTq9srOXJ7OYA1+Z4XyL10VRL0mL6309m6eWcXhkg++lGWB6aD
U9R9Nxf+kCQubTu2nmle96cmnlA/MWEwIjHpZdft7Q0=
`protect END_PROTECTED
