`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwBsXS9YupKzINa4bk0XybfYNRwCFCmxgLgGC7N6sx9Xxi5nlI/Xxi7DivrRXVKb
YhJ4uzFubpijn8GhGehJ6IOotmOxOCSWQ1/GTWikCCqN1djTIFBEyV3nzCLi2+Um
Mf4Rx5rkpPC3zt/i4/QAguhDuoWdJCLeOWa4lAm4eXVXRO49oIqHysQqkACNjDQd
fs8rZ2npHYu4YzdFDrGVs8QN01kNbnjGDV9Ghdz0Yqd47HsNv94tz9PhWUgSZDfL
aGndGgyFPzK4LJbyc78LAfwzD51x9SCAR5C1NVDDkgyzbn6WSjNbbJ66ZS/kvp63
M7xoS9kB9WmeXUU5t7C0RaCCoEMLZFMY0DvQDyIqpS4S9PNfgLlO9PoyxZnp5yhb
mset2yxnQgGlAxMmvczNUkROBxney0qcHb0xS9/3HIkzSEM1nbRe6z69QRCFq8+b
4Se0zUrwVEbSnXq+Drl+dqMGKt9oY1uXxa3s7EE8ONxTsKv+QH1m+dHQ6BE9I8nO
UAZdVV5wn2DpXAVJmX/oxC6VpBkrv7zJWGefY3zce3ktUqTEpoO+IxA+qI23s+38
xdcNL//DgPa/oeQGRv7lIzSremvL3NJCC65BAGhTMgWlyT5DnDoZXWqxJXvTcG02
/BcL07brNZqFYmGYvP1pRz/PaKBFE4yYG8n0+Lm5LOPV7ldOtvTW4pv6FINNJD+7
s9L+yfcA+xveZoViXFR7JuyMdtonx/3W5b1ArsjR1fD1bkuV3snsl5PKjItk9Xo2
6f0dkxuBaPvlBPvVrqhWKzobT8js2RidvWmNtpTLlNezvKdph3djMLOA5X67DR8o
xfmkOyxydcMc8P4EcJ90fSm7oZtJugK6768VBxHt74C1i6aYs+TuiGw6UUp3tK5H
JQ23YfarwZGIqMbO7zd2P4lt83qh+CCvKeD6fAWEQZSb3XPN9hRSKdBVzl21YlIo
`protect END_PROTECTED
