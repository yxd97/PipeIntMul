`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aTYPnDZCvmY5uWoyoHDsxTGnN3KpPVeNDuTptpMuFA3lipMq9WXvSeqy1kEtGA8X
bezTl8+hgVMWXiQOBRkzxDk93TzjM35q76KkzAsASLZH0tFQF6bBkCHKdlwOOMP/
f6fRESJy8IQ9rk15ZFQnjR4MF5Ln5B/4xqbr1U7/i8N7ivD26K10/2wKMZqAsEzr
7WeREPuAQTqtwJ6Mr6AlL41a2B76GDEvaHViMqtCQBozuXHbCeG9YwsDZYHBhuCM
ua4WN44bahrhtk7PhaRw7TT+TVy+Mt2M8BQvIhZlx6+JXIYXWP7M5ysBEFB16D/N
MZowgzm49IoklC0hIxDrd8ags48lgLaa/iPHD+3qLRdnp1WqxsEaBIgFA8wvLqDP
O3Ew0m0DwjBnR8DXvlTDp0AFLGInBAaXOLE43u7xPg/hd0i6CNr7UcJ/vu8qs5xO
3wKkmpfeLAEopVOv/wflOd8VhZ+EldciY0xFVRrvitljgaIWblII7xxjJ2a94Ud+
VrwDnsb8CY6FiQUm5o55LGCOgUxhhdDx4jf3+1U54AiOb9nfV1Gp0Upe1jlQiFAA
FdbLzWAQgCveMM52FR3h84ukgq+l+9rB1x3VvxVTQiXdKSLT5t/l1Qdr5U5n20Cq
7oqeBO9saODY4ztB4cx2Uex5MMUnxyBmOxr6E/42mRy44f2PGW+avBkSo7KvXC52
iweOFz8roo2twzT76GxDn/+hx8nh8kfgfVkHdB52sHX0QTzLplMj5nskrbjqP6MK
HyRJgSdtZ90L2vlz8o2XD30InhacnyrnAITQRJU9rSkBHPSeCc7I0Zj3WfUqF24I
bIYI1An5fTkBS6vrkX1XHoWveetJKs96CjgRV43rgUOk+3BQS1Ev/aRHDMhJDqQU
RbExnuUhSRZssTv4RJxMvECmZUwX89Z/tRpDN4//A87RlQ0JH01igp1cFHCk0xuN
NHnj7zCrhEDYDVwQXNIXNsnotWAoCsTDpaO40q4u/HGxr8FPfpSV5PEuavDOfmdc
jqJcmJ2XgPn3Gi7gACywwiW0+5MlBJv+46f0R2tXE8+rLA/CGFRQXDzetjCZm2fj
YSPOQLrDT6tjBsQ7/htYKqIY/E1OXEs9f8sgsisUeZAyYkFl6HPFM80VkkA3nPd7
bimZ1MkXFgVOl0qsSPwE32+Kwn3BULa9/PJkkwO4xQR4e04cHVu9L0srCixhtjml
dKAng3O3ejamX173m8uQrZHOZyE79G27OITLimMH2lMOtiM30pvHa2cbZAiJu9oF
q1bw9DJqb3m7UIMOtILsWjDDNC5X8/LzGmF7K+JN5lExZFZBB81AY/KYj0HWc7BZ
j9yDSHSyX21lYvW2Y0j4cjYx7behSqpcs3k+Ak86OEP4vLOUMgueRjCp3LhqXUx4
`protect END_PROTECTED
