`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIc++fAXRstu7m2M2oj6F6lgmZFFxwnpgfAHmplSqCiOZs4dJzQ6QRIe8ADAtSl8
IAES1H+Zi9T7ipmbhI/qS6/AanayF4BSAj9WhJfLoF6gTqGQwDar9JYfmqoVdeAV
DFN1KlTxlyMFhQtPcXXsaHMKiGT7ryBidLlvCCSPKsvln2n8RV3WDPV06IA6vIBn
NL6CbKtw7OzjVSQ1QESZ6BnFO5tpwSOOyhp/NLnFtgYOo7OJA2mAp27txsm69tSQ
3oyD1JO2TS5G3vAfmQQFoTHK+w6BxfJfzb7p4wRs658G3HbGVDMARrV/5vdtGSGO
NgjS84pu19YOEuWHUe0l29ecvmPxDW1Gi/FDHNa9DAjA/zVygncExxTLBbHedgeW
OnqX6gTbceigprNXvcsRtE4VSaHPI5TvE7RnCAHO9V3vAqfJvz4YznjYwnShQ/G2
uIAOqLkdZOzpn8tPznn144+qaW9DPh8EjdvfIlZm+Z8NuCJ7ObNarzpe1jVGfips
HmI7abU2FrkdBz4kj/ZabTsRmyAusWH6QovoIXRJRhEkm9EAjLpZaxHey5M9FWuS
LSViGrR7CVDfZClk4BiLz1W1BnXj+5xm1F5XQg1z1vEKBy3OpaL7f/YM5m8JHQO1
wWb0MUDZvK+BpkN+1y1tFaoJldj4LL2SBw3VIDtzltcHwMNGzoxNTQK2uIOn5rDX
jsKh5t8pqkPwjaSeB9nYKnT1/K++22j8cligI0/srJ0deNv/0rvGkDbIdR+Vtquc
gPudBzLHOQCeGwvkL8TuCeQ4IMbiot2ADMd+z6kWwhlnv8gfY2uwahhfGHFLq2w+
U6lOVSdsY8SW2CQnPDNQzDuRHM8fcuI7yB0YiXUDziCz+qWlm+uC9qLSrErdCYQw
l9M2cFVhlOwq6amGOpisUsKMV5YplGnSdH3kVszi3656f1/a3EozfnoS8374tXT3
TRDMSXH6w5JOf6q/ReOnbp+2bVTF5wfnt48HwytH4ep1DDDM5eqw+3vuzi8BJ3lg
bZ4CzdkRtqVU2zieb66eu0sdSuGS+niL3eBLC1jw15cNZR36E3QI9fzs2d7V5gHQ
3uxkdzNT6bH1m33w6RS+Z+iPIWCYtf4nQbWjj3KCbzaKigDDw/26g4iwejVF3BsB
9RYBr+XEzw1r4tcIiS8/tz3HDO8zh843PS9m+8kgBeZA8D0onQuZI0rDTM6i/KUM
2vsiL32AKT+OvKfRVmRMmyZrWKRczSznHstRtWsXotHmaaB5uqLGk5KfWftx74oO
+bbGqJT2J5jJFmU6PZf69Bn2w+f0RWIWNCzvZH2qsoOvcGBI3P/u3SDzOU3rgzuV
WSn7G7w+JUOFbxZFXMrcmATdqmEbWZMpX7bW1X+K1JnY5hwRjFo8jWjTEsKRMDdo
8sD20eRj0ESYm5S24+rBJgl0omyWWaijn9ClVKdys5AtaNv3u7M1SoTFdI+y5BY2
SfKINzJVFDZhZ1TfA8WYbwaHykasZrUZ9L23GGRn6ctmlUxK5XMPB/071ZEkLhgf
TneZxSgZGWwnXqciztMYwxKUQlN5SXQN15LQlg67SEDScXnBPjm+BqFEm0lTeByj
z1eg3bfIdRnAAz31XcXEfAEuPMNt9EV98mzNHqED3wxqyCGYF/ST3lrq5YkUrgcE
Wh6fQCuYQuAtZgz8AcMJRQ8yDgjfKtXqPHlyoVUNMvY+l61AK+ejyFEdCGHMzFXM
uHm2xtyAf6GjndjEklBscHRGftxL9bg6dp2yV0ao3RDUvOWiQSvFaZqiEvxCj4ku
6PMV3ZGKboaKm8Rc6VkjkoUKzAMCwImOHgOCbe8BIcvDaFe9oprHc0jot8eAGCAs
qBtisvtyBwXfqhsUFuwJ720OqKHNW3Owse3eGIYcoj596fJh5XsHe4jg8BAXgvA3
HcB9JdhiSNYFFBEtTe/q11FND05vom+te9HpLaatcT3zbsZvU2VEHU4mabC4yI21
g1HqVUfEV8dC6dPyMF/pe1vHrZ4wvfmJXmRQnP2QYM1niETPj5Upe6TG/fBWpdFd
saT4sKh/dWR0ILB0xz40k/Bj8kjajGiCZvf6xpBK5zzMr2kL5DZdglKd/0YOghaT
Mce4tpbUXCDjh/pvaU1LM04dPiwkbK2Cx0TFBMiUSgq1h7IrUYHQCHvJ+IifE/GR
e7BCSwBwQGnt7cG09FD+5jQsddm8Wn9U6OIZy7y7E0CzjEfSZLpDUPSeJFHvBCl2
b7QmaWifR3S9oB+PUXcE0RRM2ncm/GbOr3LUPS+pnuJ8JHi0JJlcpXH58XU9LDsW
alwypkozLJ0PNJHWNjNz1lL8xAy8QueLexYJkEbgXGhL7qo5UoggDNP5jbfcyCnx
MIvvxG2pNNRRC5PEvUdxnBdGp7XIEcjyQlWqiCznTZH6mlKsRuee4r2KHsJR74I8
4p1t69QNcChghqd5ZKQ2cTW390+TfYJz+pjihaFlXBed1WO6bmqiJUh6hDprtRNb
9BprsPvS2J8+iyEC3vmkg+TrEvk7lnH8liOQoypM95Xi5aLPSd18++lSdaeBYf2B
u0F65PsGPSYz9wzwF4ACz+TrDWl4Vn5e17HYSqAS5e7nviGY9WjEZkSvyl+vUOlc
LuOfFpUkLw9ng0QKpF3ceBaWBIlZhhGX7j4eDGv1iA8TAJ729jIkfzsi8iFzQNVJ
UOuUmTJPELRI6zzMyKzmnD9Fk0xKWF6iE4aXUsHATu4Ne3IVYG9b2D8endP+95zF
faus/i3XKrqq+sMZyB/yPfoInxWFE5Y85AwuYcaGTqFECFOuiQoCLc5jRjAAH8Yq
9pkxB4JPM+h3xqSnG6YjATI78ejKNvW3Uw+Cs9Qm3w9TaL11oNZdU3v1vVDlvYh8
6Gj1/3NlDPEruwZoZLBl6Nhsqvc/pMSYIMkzxNzS11hoBr4byalUh3nxBueDzwdp
8ETZFi1JxW0aAKT0rELlWe7skMRHucwdkms9kdCiEGrmTwfaYr2KAV8ZAZ+VjDuL
6mrA1RMv/VC7oX2BKn5mahsihgMA5fWYONID3sUt16Cno+FbRATTAnH0kof0Egve
tOd4xQVHm6OJUSvVl6ykeVgbuIBt+fNQYIxlJ7CGLAGbXI+e3VAOY7UnbHmVEtZ0
ngaJHZlpNyUHHalI6GXDyfvrlSYBv1U+AtkvuUnq62U9vzx2FBrPkRpZoee0rGgQ
6p1gjeAjg0APeEolU/1fUHZnxnXMutkw7wbg93h992q/9rood7HiSL9qUbRG5wWs
EF4uF0kEWRN7Wm0nEuLJzcxN4NVSOHN9gAo/iC9odAY0mMAfvcDmAISl7mlk9RLu
tGEFOj7sxfcvZ17eLSBBD2M0Jr2JHfWmiU262T4oxM6I0ThbfB7w6P0Midu22Gh3
mFNLkLrBIZZDvZAkrX/yqL2Noz8cNZPyAGtcAVBVlQ7oXsi2cvYZesncGCyRX0/3
AT0enNgDDjvHUULVPJz3Z+BqrNgazX9tGDnplMiAkhxKQyi2jvY9bExxz4D+vhf2
G1hujqnRQVHQoM53xEzQ2E33zBXSyK+JCPe6aeb2ixAY5vGDRVdWuwZK63/EnEer
PecuQzKRG7xWCqTiwsm5tnl72J5JRH0LGRt8kVtfqjEl9uS/yi5eJEb3ds93L3BA
u0bWE/0/70MYEdMPOnMEMwluh/FDzu3yo75CqlnzUBrauWWkAHXNJHLPrVKGayxW
fcscZSQNXVU2wMHwlrpOxs4ejCFNCvDT1q8kdBotDybtcWdnaIvFRtLt3x+k1BKz
99XldNRCa9a5W/7aDzt2yh5cS7bdrWYL5OthjfbHptvWAHkdiG4gig8+VEs7G2al
ST3SET1LYib6rmCtBwfTe4CYU9wEoDPEITsG3W/UCDSq1nn1RtNdb1raheBpZsBN
tZERlnU059niv/XGDDy/dP0rW96OLbbEegVfBvTfMNSz8K5aeRdMUZuW53QbXjWo
1KQW4o3Hww2R/Akiy49xDcGYOKB0SwOf2ynKn7xouhbpuikuZaCPgf676TTEwo9m
k/DMiFiLN8lxtncuel/iqCn2VWlha8BEcGDok4PcarpQWTM6/LLVEBdMG6ZfTdnB
aavzJkVjbwA0HWRQhdhSy2jsxQx/j1eUUxUAdtJdLMXg/eKLUSGcA8qb+EsQYad1
gOu2pz83xCEufg1d9EwQhWoWu1WwF5dseNIbemGakPL3/ShHOBeUgm/kwp1gr14c
9ybnLZ9V8D5mAGOQjD5OgUG0PE9CSa5V5GTV05lpZV7PyV+FsOmq3ZAtK4e0chmn
McLbsmqoq6KtvUhYFte1oc5ErBdnljHejfC6wwORK0zg6K6GJO7sIPap1gjUv1gh
SNIHDaFAzaMHLE+KgWLpC117CD4dO2t+M1oTpRSTVL+xfIInOZ/4tOOszAKqLXbF
8vfLvrv4gKK985YkJTFt8vmcieLQn+AJ9zryB5rp1y+kKn7+qN3mKu9fBuXwUESJ
uh3MgNLEr7BVrFjZohpLkpwJL01VR9xu3Nst0wCZGSLOnGATWXo50zhhPQTUSiMW
bHAqTbUGmXzZJ+LLCYCD2g/7WvPv45zTA9nWj9MUj3Rc5lWT/pQZl/U8K0AdvnVv
LJBQPTX+k66uUXTyFNKa1VMNhFUBRh44Tw/QaqXXadT3H5wc7n9VHsx+GRef4sTJ
4nBTh0u0YD/gG0bMH3S9lu9BVWUWKbArZErmBmQTeDbf9L5cM192woYyuzy5CIjp
iSfpStmvgcY4gD3v46h5oQa7Oh1kDlSfxjUBqv2ypxmX32Wcbcrsf6pJY9OulU/x
/G4ZbDn4+I5VmganfGnXS9W/ydFdFMDm1t4gqt1UcAI67vHuYmPedIWuNo25N29o
YNJizVN8afILjQlsIlRC//7xNDrxDpc5dEyCIFXoeLNf5VBSOUHkVxakgsK5jzjC
Dk65VBE/ZOOMsOET5qhVjcw6+j0Bp5A0QlI4i+bLZmcli8KxM2IkzBnKO5oQ63Yy
KP56kTnHLu7RyUWGzu+QY5trpXbBWLfhJkNDlgvz2k6YqOEmnAPLkfclGOpVplHn
SWPNAZMoOn5Ur9egvXp+TJywZDHPORjDek6m/GUdFF8qgXnxQIe4iQFvN7B2IHPS
LGBo386ZTVJOYeZPblsXYOgY47FrxB/nHsQ1iutxzvn/aivdC55iTd+aZKBBrHYH
JNuVMH0aiU33fXoBD0B3QiTt9dy1WayCnJNQ2xDOTBjdmZCZhxhouzFjuTXafpJV
E74NP6/wN0pWrgqd/JsQNYYEk2hNoVLSmEpRQnchNErzNgge/xWc8fw+KabiA1+S
+p4QOuXd20G4ZJuplE18oRcg9kCax4ZFTaJ9E1WpIEaxQQCOU2x2KD2QEmYJdRjd
PbtuXCb53XZMoTHOxTTa3I/OyEOai/u0O1rw8xv8PB/n2+qUvka6XZW3zBVNFUXt
ezuwLaGagJUOXetpJzydmVcY1N/1ED1vNVNNN6Qzcgw+PLl1SHg+8B6x/aTxG0Jb
wEMTOwmfz4ViB+/Dkxjtna8/ikcmBqNr+AFDM/ccJB3b2MmV8eb49DxDJJED8Qq6
L+O6LbvpqidktTnQNlkiTYw4qfUxi312Qw4doX6n9VYNBQXhrO1pKyOxBi6IFYn+
N7FjqrO9kt9yXqiDAJLdGoKe0zOp+wCgexfpea146xegNkTfXbl8HIw/sQuBcw+d
+uObLO4EP2yhJ8OEIGdPHG8zT0BVoaMfM8EpXiR7YxHlGaoRAW7Reslfl7+Eta0K
s2WLDaRMbXS5BH/ubFAEv98VINyRbSz7eV+hvTp1gCOecBCOrK2OmoVj27r0b57l
mIaGaoqtWGjjvmaokujMhddmZN/Lrm/rM1ihD9XemHEirfTqRh4jUdqbL8ByY69i
bJDljQrXI9q3ZAPzMi4WxJ6bvzgQ8IvgZm9TYn3yVjUb6NmEiu7pN6AsVn8S+dQs
3GzMH1zA9kImIjFwzVYrZ4nKQvH51750kFfX5FoUcMFCXlUerqjHDYHfqWB28Au1
ipuGU5tOpV3+PqrXs4AN2OuBOfsjvQjTiz18sMz6Vva1rjfEKSdk/nWNfZH/SNbq
ZlocwufbuaCbPqUL69RlsKjpGdx1NyyhGuX/ubag1+pkb1FAMcL5ZnimCbB6S9sR
HmOv6kcpl72BHZV47Bc/8fe/J0fqfwICc24Ekqf3vFcp0AbVkGdHU/DSj7r70Lo6
T1LnFzAtQVjTRKIzX+zbYGEoBuFdZQj7OgxEZeCeGd+50O6AYWp3lFPTRurE9xYG
CpQYeKIHpjt5dFk31Fq66MBaPdGryIv2zLjMhYM4FM1GPzZHpPFwZq1c07rlGfZ8
A3Tui5zWN9s5Eb0ktetCgfrgu6vXkyR6X5QUCOR8oZlgdUqBtH7VsOylsAvuASfg
CtrI5+CEHK7rIPyQvYVNSQPb3SgG8iHU/WJNdZoKkCzL1gaTfc4QQKBaCmOKM/Nh
l9Pz0U6Iby6mjHA0VLYb7C6SiRy5YtjKOODJSE8h+Fh5Lll+A+Ob/YPHcjw7z3zg
eCcY+kOrv4Z0thkvg8eWsm2BL52gOTpMJeh/vqmJbakL1BpQxWGy5Wk5tlk1Klcl
CtgCPuRAldgUS7rx0TAYmPSUclAj6mipv57ctVAhtcwgl4QZBXaePqKrvBPSypJF
C9KqubdQAcEA9wS7vT/LKJJjf5lfMe3tX/tr++z48oOKL4KUW+4JwD8tgLVhKcCQ
oYLgKHlYNUkNAc/PQFkvimJ5El8NCf7E+wYbXPhRsTtHrETIWmD5O1BcrYeetWsJ
eK5SOpYEuUwC1Hh81DIrAnutIRzaOwg2qrNKQEbfXQjWd2CYiWCMlPmn3j30Z3Qs
HHccE/ON2Wi540zk8ZXfzUjlsY2IPEI+dp+3vruQiA/VY4TQxt7jKzsbnASmn3uq
lTY5OMXG2hu00ZyO3JIPkm/NOIQh0e/o35Y6y45pGye8tEdfxenmm+d+BpBlwgI7
gjKlXJkFWuDwxfjVyra77o4E4xYkUnEKcsAOMRdWITS8QZq85ma0oUDmuUjdEGqP
iMndEPPj3AfVQEYpGAiFEPX1dIE3znI07LiqaB/Eq+yNZUo1o09Ntxzru8nyMJXC
p+3yrN4jnEgENUKzwxU/UvviuVVjfHpK4E3DWUQ/QT6u3mu/IN95PlghMXpK9Jv+
Gd63Y2lzB2MG/EFvKVGxvclP3mIBRRUM6LQa6ux6DSjS0S8emSjrfQYxj9pGByb4
EHvT/N9QFfrNV7EdDNo0On6t0LBff+vpBjBZsGsASkMRig0EMyHZaUnHDKkUhT59
EVNeH+nRw33q2KugTnF13Ve3q4q4Vb22a2Hvq5rL5tQIzMrd1F5k9pmJ4SCgwJWP
oo9moycVufIDfZy9y9iXEAUbVEyP+Ib7LxLosIjAduDIMbrUxOfmgk6MY6RSxSi/
CIuTpdDkd2FeovqgfjcHc5ICnOUvZ6KjV7nsdF+iAE+JEB1d/E7rOwR48rT85Wn0
U5KQcrmFs4A3uyw/rQCxWn3SKlQj/Iu3EUIZQP/XV+hQkAuKI4HtGtN77h5+1zTS
fypajnY/Uppa8OoqoSN+lXbzxc9kjExp2PXmZ0BMWiwpvKfUlEP4lJZsJbRGPjN/
Qq7Us5ANgULd/BmWRFjBbzLaW17W6PBR7oofD2Ka+ActYd5wHF/svvOvTkT7m8B8
wWtfZgtJMT8txHp9CuF+RFpdrqwHfPAk2L59CPdTFIWBYKOyIVktivDFuWH4LM3d
KiU8Q3tAmR+HKy2hlSGRcdBXrmTdTfZ+IYibWv1MUfC9hOEDyxcF/g1trAvhSrBk
/Wtp95vzVVEvuNsflkFcDlSU2tvnWuv2EpARWx8+hQK49tMgnN7oN/NsfnI+ae/A
K5iNA5kiSL6Kl2LS0dyrks7R/y1fSD7Gw1l1R4ViNh7WXjYfDBTcZe5cSNh9IXTo
w+2WVkM21ve2ZXbBBx4Pw5sFqIhk5MwQ5cg4YvUNvDWmyVNtFkJrN6HmsWP9PRYh
PgOFrgSBiSlO+jJ4V8Jg3vIS5vC3x6kAJ9NemidX5YZOXgWD+pfnKnMPDUQvGFgc
gdlGQKqQbTR8pYYadTx63YH4Ij8Fw3xjnjWQXTur5mOdfO2mcfSF/Ew5xaVKJpU3
GFamOcIvcdI2fPrdCNGfPSBwPmMRu3BrkwQbivshwhgc94X8wfrVqGhz7UlZNsl6
ACNBb+f/SX8EfRrHnHsJZp9+xTfpi08I/caS8Wil3ZoIVYmZa+aUtxFDS9NVNMSb
x80dh+upxhwCc3ZcL3fFk9x3Mhw9ot0m7IFEBqiKNcHCEsVr1Qd0yI/pe7BGtFNn
wFx+DYnwHiJevmGjt0VSOEb5Co1RB1IFZ0te12KzZvxxByf6P5fNSPzvSkCEaTPQ
LJ2mTj5taQyoKWo2l34Wrp/WBosgnSnFwImM/svG5RwJ9CFuVYlLjwsg0DuwFc4Q
pzYLTqx2dsOXGuBYT0lcPKjR5eocpZgXq6CdJTu/Y+aVCHrghZ0upweTosngKv6Z
WesgoR+ihLPe/xCb9XL9KXOPxbEOhPp5LRX9KFVnbvSeyFGa3S7gHrEjKCE0DdsF
5XPLzPfJZC1VEXXJ6Q1QkeNGfB/GhsJJMWkTBnFEO2j9va49ns/3+2e3g1Smekl0
WARzK7nQBMmJUdXLkv7ouKFXxHRtoW9u0muXedLiqvkobtdVVV45JSjUvMGa4kcm
9Y5KD80nwazlzX83gai/lgZb/tPl+pMd0S/FzXH48wkeyp41gR7CCXd+f5v4PYAf
ZPqrtgSe82Z1M/KR3WKM9AAlk3cBeP/J+OG3gyvTEX0n8hViZXja1RK+Ph92/3LD
z7N9U9WLlighQn/FPcnIIFFknVue7Jxx8SxVabyDOJzmZ6AgoSZIK3GILbeTggmz
77k7a+dYk8XWCLiH+GdrmYjUrWI46LRPeflxNYPDwMMReKOr7yaPmmqi2KDF+AT3
L3/6v1oHZsuB0q+mNwxH+d4/AtnLLYAYszn0P/ioVUbYtYJT/bedTfwXacAe26/i
Bw9oh3LLKWPK9kdtNXqhYbpM2JbHth6uahf2RDXaNZDZkbSy74RVlF0g7MDezBEN
5nha7TFzOBLl3lwJtE5VbmDm1eT3Qwpil4b8iRSpEuOt++gxTK5qW80SrAGEpCUZ
eIdx3Zg2CzqsxggqQHcLrBwxs4A5TPsSPnRKXPBuRXomaVfSm4M+Glfub48VT2ly
jY9P+fojL5GCEjl/g2rgaQQ+1owXpSdW0WUAwWv8KPEqiOHERQR2TUqMNi0NIdAU
p5v/iknmMjf39yl3WNDJeLiNpbbhZkd7pWmEjfOS35pt+eB5fFpXel7bTquxPBEU
Tz8KhFEbV5om6qM9RbLBXfDpFgYcQHCSx3gM0PWd9EW6o2mmGzEucR3gvta6U6j/
1gko3/kgdBbF7dT6AHThswrH/TrXckS3IjUVxzjau3JPZM1ziGr5WSsH3k00JNR9
WA8I863VYWxgyD3xspjcQGQRtlpRZM9AddjBnnVTuiErDaFOVEdMGbKxyQprU3ga
Neq9Zz5Opgl7uC29z6NkuPem9Uz1T54m64JZ26FFhVDoz5y4+eJ6SYb8Wrjgy3k1
/kDnIIU536R5GA/+iZTC6BPBkdnpIEsMhI7rMi3XtrbFc15APGPwXrFoHfHoD4II
x25M8clEKtf0zpbw/p/41Rlqy5gjGXEl7xZLpXGtT6Vmyx2d/5QGFGwIKFhAXRE9
3ZZuPUu2Z8sKrBeN3etEcr2aA3UGycQZ/jpUXI9a3rK69/w9B4pK8SfGgVLXpd8u
+fQ3xVG1s3lNjcXVq87sKDvMJHx1GrNPSVbsVl3qvLZ5dtZMSKw1Qy+iYXIhlBby
yFkIUz3/bTRO1oNZCG3UBxJ5hM4ClHQPTQN9J/c7r+H7LbxrbdvqGO/9BmW03SIK
2VgET9s57x8mjKhTksS24At0ZBXKtyMSq9eSlxx5thdK4wNU23F+2xLUa7IoRf/y
FlfTrFYS8Kr6ggz84A7W2PWWpmjTZb9mdwAcU94u4WOPaAObFhPrKBrKkAQVqS/t
jKCkXXg8J88JUya7OAa8w+dTYTsnbwQLROldB3HTSMrTaPf69Noww9HQbJZKcCfa
CD8ozulqUvGRSQiuKZP826uFMAGgk4IelM6ZaHQtIRzqwZffJCRjnRX5AyQDXK1v
FFFYxmiSmuyOSpb0bstU5ai0hukARQvO+f7VH53rknl4kbXjUbMCO/46JTYglqfs
UC9PHNBE1KOVxfzFg/s3SJTzL7QYB3j6uEzWT2YKUKg2SnIB/m28PmYWl3Xstzug
TJrEVdGEK1NEVNzr8VG9zkT91b8GMBtBdrSlmSwNXn/oW6S0snO5nrSYWOJvXZYV
GcM2PmTIl0+APpd3tr8yT709cFE0hCemU6jIfk+Fift33CVVRqEN8Fg1taYaoUcI
zXey3ORJR9M3Fge+20rdd2fmqUCfoClHOe1SFtovZ/JCKgeEqQiQFK8cMMYxiBmX
Wz2q0V2C5j7pO+CewsI+4SQPiupm0Tt+5jLic0qQcbGMte4VEcE0JqgvWRbBAo0h
Gdt5D9oKWA3p1y0xkySLO8PNp7qgVFh6e0fFf4oGfQSaii+8EI2lFbPz5tlBb6QB
Hj6y92E6p4BXnitaOBpw/F0CjKoY4NKPsE7vRB6J2ShnG/5aFx9cQ8N6NqGEAd01
aKDShGMveSuDXUQAgakvLiTqHO0ho8HsNDZq7FD/QyHI5GVoUfCMx/2FOIYATyE7
NyY6CILtSr3jxd5LzmrBXVIoZEiYI9JFpprXoLPMOaHyb8nLHxsxEPMwc0Yyvhpc
4E6QC9slXYWh2A/KVsj7fuV4LJds9tdyXr91+65wn7z7RZvOAlWpnsbzJbWSKruM
K0cULixYn37W5n6Jfkq+MDLPHSzTEwfmgG1P5knbS/CU1cM48tOXCzfXsRNqCYBk
w7WsuD6iRecEur7+UVHXbvAUB9EXw6KZXzVBfbop6DMFMzkNx6FFA1tn5JdYaqyH
qAmeEAYiSZftqgqjb1VO3x77Lwq7vnMKLMg1bvnv5KRCOapFUHdJ8cr3KECmXPdK
LrWzMzyOc9vzkirGjSTNuimlMAH8p0m6XoEGPbsvksx2Gmpt2aSB9CPbmjL8zuuu
YBr9iCsXCYWJNomGBUOU0qg0q9vbz3fAJWN5szg5CH3C1TxttYrCRduKCWtu8oJ6
+6au5WnIhtPcjdsh343au/jsGvi1rkCtzVgynuTqCqvGpYFQkgPf5NEXXln2Zfbb
C/+lejnq9knO4OjE5K/myxvZ2z3HIzqJ9j9B6HkHnvHRf++2SNePSaPul/Fb7+vK
ePHxi33GTJsA5nPWKMfWkf7qU19uhGy1Gta4v/n5uh1hIRITcymG1SijQ6Pd03y7
UtAtbQuO3xSy5y5sfylsAi5KrhuhROcv/OEk3Z+FQ2Mi84pqFRdixtY6dBmH4A4y
+UQIebVYBLt8xffEGgcUKLfBWHs7oO2sSUbTrz9xLmpYjB0MpbtEg2K+EZol9CHG
gaj9jM0xnxLWq6kRGErHMFle0IXdQGTsnqHQ4JAiXJB5QJWl0vXF8jt6W/uhvaRo
FvRtBKJ8EzN5dHFsA+5U1xS2+b1Fo3JMnIAnVTPFGv6G1uBwjc1m0uvJ0KDs6yrb
IWMVPHXrYnO1eqJaBg1ouFJjxnYWzwTMgTsNaVvsIDoXeZb31RLOm/2RyrEeXSMK
ZbEJN3uGF9owcxzJSQyeKmQD6sZhmzVk6xz603ELPF9I+gkCgJ68tedhBIUhuQpn
CqpWKcfI3f+sb1oBq8fFQmIOy7TKBupysHnH8fL4XhXn3XtoyBo0Y4DOPIxnE3G8
JNZjxLgT0BVOnmmhuzHUqL5asMgg+cspTjktB0riFK+5rzzdiBC8IEkrva52XEL1
Gg0zHp2PH/EZZZlAwh/CP+5SwUACad9Bz43xC+6f/heewRN7Rpcx9l/iqzeFlRB8
QiLDBbuPJF68fMGffV5HT8aJlA2t4AmQbmb8Ie1xqrE/aPxSBdESSEc3Bo/SN3Um
iuVgS0EPxEAFE2rW9VAJ9dkXh9eONCYWwJ/DNZn68qI83YEXZedu1yN+VRKGBCkD
ugWY7PJiIdopGBmlNoqA+lQ//gFQMsWYI4PUUcLyp6utxZjfhmVbewaUteyLhDeV
lSDhs6Bj8FkqndZ5cu8TYkjkTqOGRqNzCA2xTEFmSyr5FeNw39d/gdQPuy2u1YHd
zXVda2BCGOR3kipuSB4P1pQGulw+57+AT92akdLW+KUzLOplYyKvvJcYSD/zqN2Z
b2/y8EBRwBRddq3jaOFa0d8fWzOjMkYBGH/2bZot78/bMDog7ygjedEn1YlioZVC
ghZdcsx1nAHhOnojeZWdL9z8VWRmlBV6BMGeWH7ab+qrnRm6BTpK4Tq7rp7F5nIX
4MfBbx/mFIHKWLLKHqiAJB98eVcQ+f5fy7M0YrJRm3IqwzS4qvIyHYXa6rkluWvM
CwxS7mWU/znidS0C5LlfnqdV9P7vmbEQrf/nf4fThT15WVjVmqTW0zPh+ZjQWUvx
SzIrcX2XNSJ/Uk0u6glT4DYgUke5bEhlM6Qpk6CCn/Pw2VE2YFgR5B9d8Z55BkxU
imZpkQE3jKQTnQOpdIlgGV07op52Hn0S+QL4uLP3SVVGighfTCZh0puXQu8pjx10
dc63Rzy46ybD/NGa2dVX62st17l2ClkVXhmSyol6BhpxJ7YX72H84HebqccRZkSn
P6eVJ8hOKYjvUGpD+76grZtN/ANSoi9WlgysAKiZn0Ua11FOuKcIYTMNkDiAFJ09
7hcog0D3OXmRUqrzKYEFsONOBqwTaQvwuUZGPE99eD5eti1fBUaZS8ojikmTPRau
07PArr1OwRTFEiMhl745tNGjlVrGU7XBdUlOEmJgvPk6yMvWdwGQaak990k9rJUM
g+GTMaLwxrJCHmyTXb4cJGw4fAuFU0NWQCCKcweu/sJoNt6C56WiHrDZwG2Tte5I
xtZesgFRX1uYpypy+uVUTFAIf/jgd7U6Ebqqzn5B8CTzG7+I9Axxs6wVxqOMeXa5
F/zlO6ue1N/9atiXqP7ghnWkP+NULZDOc2PLbS/F8mr7fpZttSIub0SLdXtawiqi
tlkr69vQofnuhjiChyiVksKniu3ThoowF96S91C6nBO7P1hsfP+eFaS4+TIdi3Y+
zoVjykVuQe65Wg9xp88vvPLkWGdh38A0XOjVBT4anjNys+QQiH+sXs/xtkyxyRVz
ZRyP8BettOAfMDdVEebY8/KYZZ5kb4DxI75wz/7FHCFxpUnFc8cCSDh3RVBGzv34
HOdRXmNlSM+0/C/1vvUnomolOH/KI6xdFztSt9uL7fvlaSNE9BGySF8JnW/DEko1
klqNOkDpaq3VvHhGDy6zYTRdWepK+BGWFi28dlUebsOslyOmZvHI+ctWjhgDArcD
t3fksgz5suco2faytae2FwvzW5smcNbax6h0J4LDGXQWMfFHvEYW1pWT7G+DGBXm
R3A98o0QLD31NCTwb2nJpv44nqWBkQM6gvaxOAwEVYgXmDZhjuBPRuExcBtEW+tO
YjsVE23895os3oyGcxu1wC5sjaWFqYOSyv6NnKjO+3uOzv7aul7MvdQmOxkCmanO
mwWmI2pGGg6sq4/yLUwueHs+egUZoKDpChn6YbbxKatYNW/YtPGv3rsEpIU3aSIt
wrNcsTnDa2jBd/lN2/9m/I0xYelcdWqLmeWh0TvTfcaw402vMknMASg12PYv5gzl
VHF8v1tO1e2b8P+7HQAFeLB94uwIH2+HwPf6aRc/KwGzUM195uvq8VUcOIUaRql+
JASFZvesyx9aW6yRnTf9m1+kGWwGcrRyGM1r+Oa5CbeFtoG6RFZhSpckH94jNnUc
cLsmUWIKExZgPUQTCckMK/RzBFT2u65NtVPzwCNPeBSSBS6Tu4CJeSdCwfZOBn47
zulz6VOVvPCrTIeFGVd3I6gNAKM4MutbCZLl8Xoec21XKoODBWgr3JFxCqRme3+m
32Enu1FzHm0RfhHNV/lpeDvzDDPNnpf3QccjuxcbaHsYBholvhLlLc8yNCf0PyTc
k1rVKhUM0p5Ku4Py43OSk9GmgGeFtsLBIGv4tRwxi0zCG9AdcyY1Xs8g7X/pruL2
NObFT1SJk6ACJY1nBz3rRgibx4VWRXX6PooEn5NJYfvGdX2BmPZ3iq60Nm7sfOuo
y1M1WPK04+jf0hmy3jurZ4LYqs3Q4N9cDIfY/p4a2YJuQMhjzz/5ceIkzawFU2y+
8sPRyzgDhPQNc0oex8H6FB2mLyEa1egbYPX+GOc2tRnWvoRGwqk8MSKPlGjOIROT
h1nknxNb7sGmc6wEIdC39z8Z4UugZ+POLzArvsZBcB0VVRsbLNLioiaPnj0jZvqu
sfCK/8VkcuJnAz7URRlyGFw5UWdeCjxHcmZe67NOky6rAaLP6xBuXXorIdw1RNHq
vemkfY0nD9PMmumH85DlHamjvlBJ9mtZRi9i1UffZ7+dZFrWzIO9zckIf/kdR3eX
DwWs/hu+fJ96unN80EcW90riZ8FGeoLe/9R6RJuU8+d+mJcqdWhRqPrAW0DjF47l
mVI5jdUkqgCtcw7fzQF5JCEih/G4XU+p6jqVhdlaFZp6r70+ArVsKQ2U55Qa1+7i
8wa85Gt2n/fMHrXy/ouTqLbJLUpla2dKhliocwGkOonTw97+plwgkFhxfXDqUbVp
VSp5sAnqc+nknRJdkWNFVbO/CI8e5B0KnL/5VObgBb3B0uhzbylN6MAt1wxGRmV3
1eo7Z7LLRak7QTwVutyXGpfAk/ENPaqLBc8sR3EWPfE9MKan4ail94PAvXbxI0NS
lnsf39/SiGMS6UiBOov4hcF7ajlquoBG8MffP4V0jb2cp+8etrUBGYLd+FbjqHB4
E6zDZh39GyACHeM09GuiLjfsjkGwy8D0jbZOV/U6sBBTot5X8kmF2sgrM8w4rLs2
cyS6camGHJ07q23OZkHzk2lv16sQr17rMfLxZujYEGFRzqaeIxPvIjrGR8pMO4rv
Te/LZianb9nqvVanhbQNd6XxGbj4lbE2Mf9D3g5b3YHBSgyC9RIO5dOYxjED5PBV
9ckc/4m05f7DJAQ9/MBqCYFPgXME40S1kzWh3H37/Kfnd3HXzO8TUW0kcoAHeh5p
02OUJY0qOqrtKAjLYo1dxBaYJOf8yc4APwSmRz7GbGyJ/lnVnFaDoa/aeUuPqNar
umbmFlok72e3EArF14V/oek+31ggZEvrLeuHYlGfBy32k58BsLAPBfPzRrYqEwjY
M+BtSkarxFaixqeOLarmzICNX+Ab2uFpDFxNrmNbGVSyVxTPNYOBUjBjScM8oWi+
hRKY9RQasrKreQfB4CuEyHh76e9o7k0IlS+aIHCNS2UFlaUNR8UzzYpQT8Uwkv4z
zm+POjRRbxiVZPPZADu/V9q4Nkrxe0WjRRk1vSg0mLjTUARKyaaK7S1PZsr+hACL
2MWVZqQ6/7UMPjWXnqoEDwmWwNRqhYJO2GFoW0Nxe+h0ZDZF9fXnLLrs3Z6YBSXa
0yZARqBUtx55uHcX0MKtQCCgRtwSHBtovC1s/QVcIWGvitl65bvrUJzFRKMZyMcS
k4s2vVbJs/2X2Er0Te5Tj121dUezeIy3jjQkoygaJRIsxrPHDOgr377hIuZRkz6Z
w9hVV9HdilANIwIfTECD0/XlMg6EPOZYz0idrNrL4zTQjpq3Po4bvi7gYMf15Dma
x1fn0M8QTT6ZkceoR9MEVlurBeth7h2raOzCqP28Gl1sBG7Y9gndlrszFupGoZoG
k7FGybGDUQ7w8y8wP2zhz1dDL/97pmkmbXZlFXtLynKPlWnIowcqKRUTn2/ctM3E
QZfXb5eaWmWiWj4+KxBZVLCbPfSsPs9R93uetfo3JDwSS6kjy1eojLPca9tIryFV
PgCKzlaYmMUghx3Gl7WVDI2IBcOzJNaQ93zDSRxMo16vIDkXME9iV0cq30IWVwXY
70d4OveJRkoARVT2HF64kN+SUKIkS+A7M3DJTR68Gf/gcSd2/1rfm7r8OibhRX//
yJSDlNGxBu16sF6Bjge1EdUmCFB6ZdLJT/UMsd33Our56VGgO605588xw9xagPH0
8MANjVZj3xzHaeRyE/3ATMpRs5tOn/TWw5eoj79HINWSdpWCNhT6aUZ6bPub++jD
6PUENjBzq1Y48LgtsmyWCMibQb+FzXp58zrhnvBVgKQ11td8/se+TaLGXR9O/WZh
j3N84qSLnKow+rtuxlUz2pI8zNltuO0rvxUXOu0/NhLI2bdf4bGWaeQApNCpDa0U
GpEuJmplCjzfPH27JjUjhZQ3YJK3gkdC86cpbgGKc/x2R3UsR/D8Fg0zTF38DP+X
XjrMEHx4Hv39YnSrkmRMJ/vUEZjyQbl9NWlTs8kf9IIeUEJVw9Yx8413skBJCSJ3
QBOQOGTx3+ifEgY3RV1wqmxa7yYP5kLqQvCPV/qaRadpqgtnuyypSFtm3aWBSSJK
qETuLo5cDU12li3LkL9fx0iupQJEf0UB4j2lBKsRS3KrheE9Hz1xf5Tkjl6xE4Ni
DzqSpXyB21hwzHSlpTxVVgO48MfDnj7aCXd/0MoA7soJnwf/gRBeWhROf5pA0ez7
C8rnjVgLWHhQzw17FtyO3ZT2WLNUImHMh2SFUlzlN8l+5zeyoH1s7lVOwpYc8LZg
pCgyzvfK9t0nmhrsXogpuiQIspEdWWShFKrV9/UT3ymqU/9f2xMKZ7Y1WfRgLsvI
CdCSp4qOXcjiaanOgHkhaNXNhuhZeWRSd8rtMu2iaOeFZ4sFMeLRX6X1EigM74jR
BNzeQ+//E7sStghzyCA3iokNm4S8v+KJna1NISPQ9ZnaWnKZcchKyRzASJt4MsPH
KJ96SAdb/+cX7TEtsf3p7Q==
`protect END_PROTECTED
