`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oV2+q3txh3dvvzY13nUwK7676vDNV+fOJnsHrJckXUGeLOazXppyKhERH2poQ2bR
frqu5tKkON5gBWY4IfPp7SV3LHeOCOqCEmNYBygcNnWZiYy5Qv0VvZEN2t+NVcPB
KRJ/YJDVwjDU/RyMACsXvz0NuHUDY7zCN8Pr9QRu6TKxWh1FdU5qeqEwS5DvH7bn
xPO4TLQj6Jcov2JkkhiIeZV0oBEnlx9iGz9ErgD1S+GfaRHZa4xCgymjTdd/IYAT
4Qh7FJV3QaR0tSG489jgp9KIklsg3lfM4oiqdUNqPJFyqDVVDq2GaXg8+ph4+6Tt
HfLLCHWD3ilVRHoZdNuNcWBb5ASZLkAFbUUIWVy8qPVZ9PFYP/SAZU/W0ju0e0+H
0H01VmlYiBuL7XoCje31gQ==
`protect END_PROTECTED
