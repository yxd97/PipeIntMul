`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6JniVJARZLoinijOeIpfXOgTGEQZGYsh55lrtjfyDm4wNzR6gqFpyjeL8Y9ZnA4
UlssaSNQKNZbD3bobQurAFGB8bMDLNwY9EU7IAtSU8XmP4NYhkJEGxBaIfl++6Rz
5psIXXopUvnhG+J8sHyxymnInHjxLgEkiSQW9M+/Lsj34UvWRgAgLFdJ+Hzdfi/a
pY9dAZPMNTrvV3KOXeP1wcy3KWEl8rLw3WDsh9d7MchK3we7ecJ2zQwTreV2buoA
o7hSxJnyo9OBKYci326CXZIn9MG5usbOgt7AnRuZsZoBeVVsJsAR5WJIJiMGVQru
WidLpL+SiTiWWLE7cqcKu/ZmBRgsh+2MTeAAAqxq+9rW4luZgLhiigaEHI5rqUoU
vbIlkoo0TyF0diV37UqetI1k1vZDkZonEWKRzntWf/LccGZIic3GkDBr/qIyld9A
MqPi0llJC+8nbA7+oAPIocTps9PMkwtp2qdAGs817a45+YMydygjFZ3iF8JsYAyI
EGa5OUSnCeVAHFDqnTVbCXpuZ6JeMbDIa4XGm/04TM/cXHWl7usDzL1ts/D930NR
1vR00BNYphLCHMw66IW/AHlUahMhdh81PtEV2ROhAbED/OCuF+9wsFV6cRN10zuM
GEG4/L8Ui+zhSmYd+eV30K2RpcL+NiYwQBB/l/KjBmYV0yrAhFwTjRU2Ec9gdEWU
iPe77j3yATrIfAMC4quimyzvafpIgrmV+l10py9BOil3rY2i9jAwo7O6YVqbWbyF
sj1DoS4Oa5S9xCjN5LQMUGsBauvjkffHh9IF5ErIs+g2SXWCfO7S+iKVx6urpFfu
LyfTLZkkevvDyPuyZOXemH3z5nmYM3tcRHxhz1DgMmGUzUZoqfF+wD+QPeeoN9Zu
`protect END_PROTECTED
