`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o0RjMz1tBLYdXnRtk/o0PNz6GGwytotq+LANUjajvlr+QVIv7XOkvKlYOa+fh7Xv
pHdVv7l3KAAflTgjYwg2/CvBR+TQ0gg477c9M+ulHwN5YkqeXVOxQqFKhE+5PoY5
zAsfEWrug5/ewbOSm8LD2rK7pYIsMubTdPk2qDCPe2JgOiqFsYf5YLMhbY1cMQQm
vqJuSH7GXBkBZ50l0Cgi1juAOniA6JNKPeGizG2vaWTx+BfRt1vWH4UIcjXAHKJ3
wT4wHWlro4Ihoay0runX2RsKTYzSd4drf2aUkx+KkIhL27pQZJwP789GtbxuUq34
YSWE0wU0J6AGT2rY9tSf+tA5w0GFJyAPaX/Izk3rWPjrzhhElRfUJzbVxRehXCI5
OqvjXX9rKVHZv2R/zYauF+oTD4zMobw27lfWstiE50mqD/3HIfS3Q8znnabUVp7h
5MVhhA81PpyTaCs4RebnpY+tYiTH5wd5IbZKRQ29p1+j4DuveESaugJV952GGAtJ
8eg3+vf0UdshkLgTtzlcV5/5lf12ZAhenGiNrguctPIBAaqND2OxKMUZgBVbv6wi
viCUgRQeX3qAWBmtP5I5eox6af+m9YxCAfVIezOe5NmDPeb3hCjyNncmZsASySDD
YaIU2QQ0NgMB+82JOJizbjQcMaz4uaiZfFI4aXFvTTK26MaY7eaByxLNHerFjINd
J+l/+kHf4NOksXMK0GU0cnnhZAYdYFnKlh5M84QPh0TXAZqwcbR5xV9TI9VUG4wr
b+nDjiQvlFHL4ozx9a7TSPJ7nfW+Nc9eAA5wuRKKp5gK7+xx3wVDqAiTPd3BHszR
zy4e3qiBPWQEmYQVUQlPayRfylSyKQMahz+fgBREI3KpPQKF34sVEdYcLGbHGX2v
4WI9ZWQERIpPh+0RR4VQw1LE3R9TkLWMG/qHHM9CQgB93CbOWcm0Y+vpxVMObdlU
fS4WDwPBL0BHzw5jrQJ9oGqdyra+pa8/t4Fu0WebeX3q/Hwna5qlC5GLTWPRSQGl
MCDVy0sKMcHyT6bk5xDiPF/aRhGBbbBudvm/T12FUo5Pbz51nQhAHuhwZyMcKg5o
cWruo0aBtRPcGXFrNXqtVg==
`protect END_PROTECTED
