`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dgvYET+i7QLFylBAPgXcO3MU67nIdJlQzOwj6QCm51Bh1wwH3Q4jfg/EbnIWJWIn
IcedBsNq02FUaK/0HEUE4cFHqRXiXK5S/uGwrno+zCeiGoLRa5bdaLzz5/+lyfn/
xSzMHgPIHUuttMpNwlR/JPrGHCa4OolII/4jGZit4WnNKcHbXpTpQPD3grG4UzoR
DTNmFlqjw9tPeudLC4dImIHJrNz4uMLHx/g+js8isLwKHM6WPI96ofo/MFJR5WyS
5EnP6WUY8l7ge7JmlEWYmKdtuyS8Uwv/hzylNc5ltcBUZ89n2Flon/6LMAPQHddU
`protect END_PROTECTED
