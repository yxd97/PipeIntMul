`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1sFHa8rviUcos4aTTPlDPFYutfPxqs7XhGgfREjePbIINLUaXADfpz1D5dhR/6oS
v6sm4xQDaannpp7tSBFe6vMI7wWlIh4pq3nNW92cm8qaej88NXuWKQhWXb6lSwyu
DHMVReIPu/9wysYjlQNqm05xD5uRfDGHYQ4QLTJiLqXuIPJOiOhro0Gl685/hr5s
jZaQ5yW6aKqyUapi/OUwaubyKbGxtXu8alRJsZI8u6cckimjw4mUhzZYP33e+NOJ
pnMFkZZWb6K54udP9k5wFqMZhgfBdCAUsmxfZhQfiYGfth0l3wKffhw8iLf195Pa
7rRf592C56SBm1yqKlAg25HbTDpS1uF6UgHf/SJNnBKP/2/3RLyPilMNeelP2W64
ObGSj3eH7DA1vYD/am328oyN4eSfSut/uUjRmpOtf0P/XBO0svum3H7CUvnAAlCc
YZHL6H7MkzGuwJcOVZHrJwZ/j05R4S1KqpvmZGC99PwhT76580LsLM8bDXZsnSc2
mP8BztpUPbQbTgVO+UNLkLY1M2uTxEaiASBu9k5OLTcPhjnXtJ/SD3BpvvYG+q7m
8BlAV9a27JSQBokjQeJECarzyr9vneguKA38ZhCdN16i8emBy8EiceTxnEJl5AIU
1n/YzlHJycYbkHp1R+sCUryVwM+h9XPmmzPwr1VNN6cphl3B14H3ruUK81EbBygO
Z/TbKWZXFzN96SSEoGyE+Db2Jxkz9TKmsVcyKpW1mDtuylmMzVXZwKakB+GbIDpV
U4n17yUUMqOvQyvOOda9lPrUuCsJ5TioeyE682DevsL3qj6C/Y1XRPp7D0nDYqRl
73lx2FbNxlo/lc8RAzCRjmyHRQR9iOC21hWLv2VPzTGmBN+2/eEsP1jC21+uhlwt
P8QzPABTqEKGVWGxhrCmEytEYHSvOCiIEpTPSekwNkyCquMvW7/m7hK8+rXzY0j8
/UpCmbcWkFxLXruoZHGLZ/EmwyrLcqTJkdc3hEbagif+n4qs5CTiLXCrfsYXVbi4
TIaxCj2T3maiVM3hN7zwseBN88zaROVHCifOl/nL2gY0K9WB+jVUX02xslR6itf8
z66ggCeqircpl3kjBt9if03YWyVRYbFXxnEl/Sg/CiQlwD6cy49NaA51yaxT77VX
P80nvYwKAcHvR6ZJ6I1GdNePFJ09iUBEKkLS1eswhMZdlSdvb2F7D2S1VAgZwqNa
lMPCkGywUddWJPINsz4N729PKS6441P5tSwF2aO7VEjXlV9TZSJjeNQU+QDGlyjM
eRszoS84DLtlXDFr2ct4hZDmIuNNcTBLTUlBoyrgtwBbRAKEpn5qgIg9mss8P8Nj
te4+CaGK47ePLOW1OjlmH0oUrV+G6iNKXEuWSL05OD9XHvS6lIRNB7O35TDxSs3v
z6z2pPZ4EDDy+Ayym9d97eZnHLlAMFoAPhH/4l49+jfvlrVrwmzQQdsh3nIXhA2u
swRHUJeAGDcQBgZxW18M2gxufvTgOB/daasNbNOO9flk8Jd11QEebLeEUQRjhkkb
0yCsjNRO6ONKE/c3HHm3kH2nM+uZAzRK4FCdswgQpe2Asibc7nKWCgC+5IuiOfSq
Aj5sfC1nYkjIlaTfD5osRJxWRdbb1bMCbstBAZSr2qjrq5OVc/GfB1PUiTf2tIu5
ObFuhISayAHUxqgXosQlYdGiSzdIITSb/P+koo2IxR3UASZ7lkzqKJ+cZ9zRMJlk
JTMEURPUb6Hi0UK0uwkSQg+zGYONUA5Ixm7nGw48mtNMCWspDmselRsXHUqdLNWi
zZcjXLzJoyo1kKvKXSEeEdTAo5KeCXuCN/42xePBMaxSfs/S65MthM1jA43ahHEN
hZpRjLa8ysINVtsRCTEEKhyo0lItL4N5kkKAvPpVfdHdyiN58ff34xiJUzQ9te7c
H9VOetIaGWJmBGcvsGJ3ysaqkaOlCxiz5WJu3tsUSOH036Rg6MF8pU7kcnBp0JiV
sS4snmjxyQXIjbY6Zxjx5K/VUEEUFuTeCvjq7EQ1Hd2QlOnjkEuXyUZXabfC2Ws6
5surrvcXJzZUsWigwymCKClgCO48x+s0x5YT54OyYtT70PMDgZn+01bHpDsISNAD
t98D318OcgCR1YhQEtpaS2I0K8NYqBXbUAHOr4ngai0oGbsW+XetXJlrygWtEtnK
u0GCHpDqRbM/p88TMB+FMNqPqy2KNRs3lLgFmfU+4qNlqMd/ib8r5kGxoC8AdNsx
5ICiOcMti9sJrtMlHuGGI12mPPSLL/xNnBUVES6aR8wP7pj258VqnoqLM2yRLiAX
dg8wYOPMX7QdmzUjhkTgIWYgRtWJjvkvei7bD3K6mzn65qnFWnweQV8UOcrsTteR
`protect END_PROTECTED
