`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2HszT8TssL/r0l3iO/vR1vld2O7fkUWJFkWglVHtt4ps3dTmGJkj175Krpiz2POk
tm5Ikb47dW70t3wTytdNkizjv4euWwvMP7OyKtyvrGYgYpUkaRZG90rih9xBdACh
AdK2VeGr/gS+Im7PG1T19hDVFUThtVFiLfKB+baTrG3tY/hac84HdhkclTpG3coq
JrRMvV9kckyLNLHVLqV/N229/kIgazMagfA+YuhfOxdJNNXNsSOU4d1y59eEd3Pk
tkqPTxZHRJZHXMInPj8sb0w7UzNvZA/RglLa7RuI7q99q9VZR5dGHP4+K1tm45Yu
Lx9ofyB7IOfzBpIuW6YsO/acX00VxWk3zddiAw+CxGWWw/49hL4mx792wUQdK+8g
jhp42vuEZeQjOYbhCut+0pkMzchsLZ8mcGVfUFLs9ewWrxKeG6yi2xJdsA0Eo3eS
jszHDu2fEsj5Yo2JpKuLyQAdGeueul8WIQwKzg8ycHX8z0VF0S21yaqVQa/xeZEX
8MARuibzmMruIJJJXae1dN3sZQ5yjBItQTDmXvFyjpuBbcVXtF+BX6Jx2TX+U9cI
kmOCjeKBL8R09ES/0CRQqXm2X+2q9jiM/ofSXR0Z3+z17Lts9mNBX+qi5L25xgRn
WxVhKR+DsBlZvZmwz31bF8xIeGZ6a3sl5VLZVFToY4U=
`protect END_PROTECTED
