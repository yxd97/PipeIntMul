`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRhqKuWroItduE3VxQVGb1oTzJdFLaUgzKRWy9PfDyLPLVlcmQB9pDIibIgYMYyq
Low/SIkJjhf2Z0icfpHZr2qIy15HU7aD5A7j7CZfiLkQX+2ucxQ9/jz5pYr3Urqp
5aTaTfFrQzEjoH6QzjEJ+JvCvJ8/KS9av98396sOHqNqLFJSmLLVyn5edsJkcj+v
lMk4Es/dEkFOmya7YN+NvmEHugHUGQxaxVj0ocucGIGJB9Evk9yZWc7JF/V2Gjaz
RggVCoFvd3VGjdodPJffiss3U+CzL8BTsPRk04QOI3ABT3tcqO4R9kKQ8nClarnd
FnnT9F3Sjx+J4r5MQXYh842TcThRz37oODlEtnvvOKGygXFIq3FvoV+mojcvZnpF
vOQAhhu5xI+K5oHHSYLEig/mpr2A/42OmAg2RbPWId/u+fcD6s4QyHAnWQRIYuCG
wGx3ZohF2Q2KdwHkkNXXR3h+JKS7JY4MesriAXfZ3/bD/urPSU4/Bp1exhf9OA9u
FPm8USmwVpbYQtSn9W8lZBLh54rgb328dRD6h5XksSCYOLc5SCOy75X6JLBsR3Th
/vv64uPmT88nMZnwSbEPgExq74m+WvPaJOEbW+J0acEkAE7JHvfx6BcHhp6YEEBj
`protect END_PROTECTED
