`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDuCyS7pgWz/Mh87kPBLWR7/GsHsIU8h7FbPOUh7bMSirERd1hYqVP/uPDQPOBiU
sfkDvzu0x2ET7cXEypGddcVkrsEHveMWt8YNiOR1Hxq1cLOG8vgnz2hHwvrjksas
1fIj7zVGXWxeiy4PQZnZFTDHryo+4Z19YCrT4NIHNk8ov0PEK3tUVGuEK5X32crt
XTW9d/8/QnnZcq5ucD0lFnexaxRS2U7wztQ0gfmGVh+jGRK6vLM/ctMZvAJnzBf+
Jx/gml7nFHtCdkbNEclAs5ZEB8lBRZ/pF/2NstgLOfcmF8Y7AI9JiehTroC12Zc5
5BZU0ge1azseaIHPoJE1Dxg0Oqp75CaWxYVC9/VOYMHa6227IIoZGPc94wxtPQ3w
5qjfPS9RFOKGuvNh5VbT3t0YHz4waE0wmaXiTuJ55ObquFd1PEx8GeaQuSoqNhXu
Bav2hWXjVsG4Hbx21gs7On9I2KRFfKIkuRK5TiOkvwwD5C+BLRviZeo4fa2WRCh/
`protect END_PROTECTED
