`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
noi8dqY/9wGatFjtLV05hkArWX7LRnAjRDZUGgQ1mzNnQKyTa1K9IGjasGmngaXa
WPJArgqAXNRBs9C/LUin40k/Cac5zswNWVM+JuwrGjxPJXqe4impA2hRN8RvsCFR
nGSBmUdRNTIYhHdyqA2T2I0NE2lRoc1Myv/Kr7zZsOpi8LTXsea+25lh/I3XEBPK
QuallnRumz9T5dsf3v6XWtL+rFrOfnfFGUh1YCbIREUERTkDB+A5rRmlOU4wC2yb
XIJdcwXqOK4PjRLTf+cLn+5evfjOVBKtOzgFNOaY6dYO3uztBboW+iujvJJY9lWG
b4zTUbYbIdZ6dcegxscCwHKrtwN79BHhtu8aJSj0M9TDQbN1XW4F8saWeAzguDIz
MuvRCtxIdzc54BLz1XNtQ7DWmEVBZ+VNk0IkLzIZora0KmSbG8bvMHyz6iScK2SU
+1cLe0maDVaD6rJ7fcEBd4/xvm8JeO+lVzB/OjTJapdTgCKFjvNDsvAsrkVJ+nwG
`protect END_PROTECTED
