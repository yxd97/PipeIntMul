`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M5al3leBPF9fn4EPtLmPH91eJdc3qED2nahbvMextWhJETiISREMrfV+xYJlSqzM
8s37lLuxJZkwmVTH4uQUUccaUbaA6tUy+/0neTfkiJQDR0nlvH9mL8Cqh81lUhLL
JT6W9Wz88chdegJqAgFuw6n+JwGvwXGrVmJ08ldVvRhuQzAcDlHB1C1Xh41OlZ0t
3A7BoTi5g1b0/t2EGMxyokTxnTJTNyh7yzMkLT63Tx7NfpALtJG0Xp6LHfCU4awa
Ja9TVdOgNsUOCkm56WvECfcC7Yk9LO6TPxO4qLHGclIYzDG79epZt/rp55K05M3w
hliYQrHQ7D9zkKke2bOdW89Ry0k2Vxnej6DmWpNko6kRrH1sL7gLWeuc/vNi6U3l
mHXyeNKTGI63clPLNgK3cTx2nlTKDSP1g8W/GDu+asBxx+sJKK+ktIXGWQbV3pBg
D++jHK9QsI16vg0Ez13krrTpHtjHRk6HyrLn9wBFN5flXbU7WN5TSJPfqEiiBjSc
FRuyHJllG1osVV12twRjue4GePGVybAGK0mwc2QsZLVAXUB6qI3co+DOL997rt4L
VvRZR+gQfkA0X/Itghq7KK7hLJ3EQcXXXCPM5o3ogC+jvamvSy20EXs89riONSx1
rn68yol+rFZMoYYT7lfTyK7nrjZEgkqtGWrlfLrmI6p3Z8TUXWW18bytvP9weE+q
2F2JYr+bDYOiSnQ/PcNyICN0gNgheTrgsk+UIl4bRC0JICNuZ1oGXuWlezg4Eq74
vQhhGntbkRa1PtpPodQSgp5umBBn+ZSlMsJvkZGHXf1M911iRpNzmWmBpgmozzNL
oexaxtlRKG00vX7m3Vx+mnkl4yFkl3B241oY5lZLmqCJS+17/q3lcZfE1msWyb5p
U8tjzVod8QAqHJ40QojQUHns5s+g+VMFQ4iliGCkoExXtkJ1NHVpSKf0npg/+lSl
9FbiJU1wXeF7ahPwHIkldBm079URqJBDNMHYBQgZefyG6uuvbXmpuYO8n8xQzvTs
EF4y7MWhC2YUxOVXWT4vZOowRpcHwN5vusa0Er+Uh3TFG7KtB0Dk3v6LxGooWRK9
rXDUbjM7NbIjwoEZ9WNJwt+MRZA7dYuEqU/L43dnzr/oZzvXgkOkxMWD6fVO4R2b
ZMQfJQaJFi37UXjIJ6jVyTFPnAOcHb9/q9mg0g+QKCvlc2ZNotMdSXFBdp9C2Mvo
k/EhIV7S0iSZ1f8eRRzUWvthyaEF6/o6pgCQfooZqwWpSVb2I6ejsqf5iLhRU29p
zRZXdPcyooKgfa0JV2aAOtWS+QJP1kycTDD/KI70ROBJg31dJzXQSqt/uijNbqQ/
MbjVMNIkDpMhnV0q1eEPSkID6l+GSi++myJwI9lLSyzlRNsVdZDSyxwQyAaW2xtm
OURDMiiuDYzElH5GwJqyxpIqfC9H3wBnbRlTqArnNKSbbOHVO7F7zw7bpF/t85Q4
yi9XW020P3/5gRACZRnT+7T3SHMvJqtnouA4UnIzgVroqm0MMCqowZcK+7dWLpbR
4Q7WcjVyPDVcSqG5s7D4V47bIlOPcctTUvzfKLFFQF6vC44UTAqo/bOPWek6Q3NV
aFLokeLhEYSW8uB/qbyOnposcAXItRzJtw+iVjl00oWztmdXs/JI0V8OGj1uuzGx
M8xrymCJ1VEjrJogdBWHpi3GdEuA0tGw2U1L0nHnjHGyErFz4fKLlZCXb4Q1JKdA
ZuceTCD9dFFL1GuaOle+k7J45wH0eZpNhaLXd4dJm4/1cuOhJ/G4lGGvbLiiHacI
6uwSTjbqZnAcZcoQxHkF6Y0MBpWdhhOiDtK6afqb+2g0zH1p8vugILf4SmCUOqGP
jEs1ReHkByu6hkd9tXPVYvR/bhuytSS6Xbce+VGRfLuAQ9VAU6oLwN7z8vgIwvAa
s9uwTSXlnvr/ESzFUVl35hjdKzET8PV/z8nhdPY6WaAtL0ExrEY6P6QYKxTGfkqn
CE2PRY9nHEkvLCfCdJ9ml35dR9zy8Ao6g7FbCmjWPRbvud/tZ54tSCf26OmhwfkT
c+DvXORHrtUlOTVIfPef7YhH/sBvkgbqg+OnKJ+S13KFUOep2d2FK8dDbORasv/N
wVonF5Es7AKQ6AA6QNO/3atV03Rs4EfWc8HK1IbfCIDEpV8Zc6bRAXkXOHVtsxOr
7QVc14lkP0amrcm8JFkD+RPYypk7INXowKNLp/qNlsYuIZ3gBnK0xW4+frE2zMlm
rxhENh9TD5FweXuaOXyyMgf2dOY8blgaclymtL407nrE2Kgug6ASrGcl6oEt1rJ4
Mo0uXKC9clCsJNQL3Df4gv19T4k/3m+bVgGlhEpQ3D+EvHrO5zVwVCw3HgQdwhFi
lKpXzVaj/J+J9J79Rm9bhdvWa46CoeY8uEgeXFjR7Cn0P7rsZpcLHm8LIkY6mJY4
E/PndEkkr1J8OSjBkciW+QStBJUGXkQPWgcF3COmByuTDpsthVMeIdKBWlvMsoLE
gCyC26YjMSeXAyJZcLrWwrMFx5CHhwJFBxhDWGcbww0IAB3Wn52BDJxWYND0Xomm
o4fazcXQ5Vdz0hwtE0c9dHKOn7nEpWsDagXVK9Y0OFZp209JmPrw2zPvNxlBLTYA
QPkUkJiLW+gGPg3K95f7lWbkMe7BAcmFdmxP6JTDnNtmc0c2JZWg2NRif/fEkcUV
TAS5P0amseuGVK4+xdPjfe0C6JWVBc3qdd8INF5DyDCL/UeyyweJplczfp+Uw8qs
WoALC6CouxoS7vCP2aW/ntVbSj93t67pF2lkbe5O3D7ZKCvAtLO67RNqV5DA4KtG
dd7h3oFuZIG4ywv+YGgm0iJoDwh0XJcNGQkI8xoccjkF6P6QjkyX1Y8KYVAtkzUE
rjpqNG+4zCJskQRF2o7R38pAYpEeuV45O741JIdCWgg6JBuIFWY/9IQlQnBhEyKf
bD88JbdF0sILKAQmwY/wr+/VEZ7fmyKHXwXJfBuPh4jiUXG4yXCqSIvbI6Zi9HGS
WctEv2iNbic6D96HYo4N6Y1e3yuMiQnD1g7Okp9fKeKfvZkp4yuqSux0kXoH4A1G
OqNeTCiV1v0IfzY+Ih5lI2OLlqMqhXeLncQhMZfCMQGrNGa1cAgNnuIF8jHhCt9f
4stq/R/P+2MdcaMy2QcLB+yZgwkKhOUAnm4CculShmCvlcD01/M8FXcYW64MxFn8
Z3H94P5xxmfOvzZ/k137Rxl7MO7uejHwM/QBBNUMRc2rolmjmgCxHgePolvZv/Pe
dtchAZ8+QsOkuo2r03s7Vs7M9LWx1+vNSPeFhc8sKPn7hVr/qTAX0bmTGZOAQe6e
bizAk28Vkb+6y23PlbAVnLiTOkWfaZ6FcfDGmy7DI79IdUZ8WI6OnhodcdHQtiwv
hNKxoiQoiEmWufNNjidH4xK7i784cZj7gxhxQa8wuKeEi+tMKYdd3Idx3kgciF6N
hQhyj+zRG+ZS/i0nx4aFEk4e+PKQU0GOzaVRAGe3jsPNqUxDq+wWm9TQigEZIxHq
lI86BPKOadK6uBhxe5RbZRMwy63ForI3eLgVXiHf4OTIdeZL9BxPu6sZVzPjaANH
mg44Rm7KbSHEEXeqH1xiCsArStcLAcWKw9LXvJT7JXFKwVMJMjib+ec4uKDrcsj1
P6TwBserr6Efud0Y+4bC+uVgUUrfzVKH+senkgGVpwKjxxGtYiWX86UT74Fd49bN
Qq428qqLbvDF6F22cKAajrqmRCfJP5xcZCPMyWBqq69UfDiABIxnjRrfZd452hHN
a/s5T028SHviikQMaN2GsAQV1F0cLVgG8HUy9FT7z1VyhbiEk9jp18t0b2/RDLk0
riAuejqtNHCz8+ofb5ggeggchoQT9p/tammyZmFTBPVu3EevMn4VgT9XcfNARXIt
AtON/7DQEAoKz3v51kK+lxnuacpET2fzbqEVocREAue6STTWQ4+yV9iejpVlPER+
E6psprwofrq/KqZvrD+HfixOacYjEWAXjwO5tM0MsLuyc3uVJFfQelv0/4fMGg1e
k1hT4S0X/8wKivUPsn46TYEXdL4BCiX072JiPrN+0Rkr6FNR4UOwmu+M868ckywH
I6X7qQv62bscAkHA59MrMy73xE6Wi/VOp3MJNoY4isaq7ckhx8um8S9zBltKIwpY
U1O5/VpKFp8q33GZzafXpi2e8NFkWYSy7KMcaLwyBrXKeONb/nkelPDfJddvk7H7
IaS0uO8y3EGjtpp3G/fZgr2ALoKH5vlSVNF+kkUC+xGj0Q1HS89/CwPVzq3CpqDJ
W1Rrnsuil5nqMV8IXwwv8GwT7mcYM3P5gCXTbTUdiclaGEMjZUF7FJQGfU5QlDxN
fq4168w8lYPuTrJenuNMdVzL0Ed/ACPfIUvcEtTpN1Eka34hco7bEENASUMeZa5q
ROxTb4eveuKfZHzmJZMfJnFcJzrQkwEXOy1iQy+9RxL4hsrqgyr1IhyOhiHOgNnx
yuABfYEPOlCMvueTSTkWTT3pJImQedYUu6svA0JUrti8FTXZN7HGfER0aoXnjqCZ
4WW+RS1StpYxTVIxA+iYcXgrr2XoxFTZ1MaPz3SLxzlsJ3xP7nkw1KVyYfXfMw6E
15fp/0qRjUPiFdfu6kSU4R9bZLGGOZ5DIp7XL8vyh3PmNox5BBtAY5obX9jrVm9V
v8FOKYK/EbzY9NEKh0CMTW3wN9hQrB148f0Nt2Ig7DeTl5Qmd55paJ0Q97ASly6u
dWi/wCNDCypGidTZOr0Zs3akAeb/3TEHCmfo5tf2YllkYQ9ob6GhCXkDVWxQT8qR
aMzopjQegFYj9mzfus6qGzNmk51xGme4SRSQazoCHg791lydSb/2ab46mBqCqjcW
6OuuUnzNcXzvgqqNDbGMpl7jdZMBEN8p87Xv2fajV3awOOUKFOPfqtXJnqujwEz2
ATtsGhNRzR9o3jp8YO8rqjwiWjjg7fpwm+gSZvYD8DO4NwmMIwE9Bnm8AIziS/hq
xhChJS5fKSfhyNuc9Sf9j4CkFW2Y73NfuqxuoOq2vS/369vP00G7VjNRMxGhU207
HY0uhijYeeh4IKwuea7i3+NRRq2ChDM97U/OrsnnW5/jGI0ME019lo+li+pssJ3f
crvTM/4zcgOM9Y+3+3oMhK9ujXn/6UGmD5B10sez+a5uu5I8WlkpnfCKtcH/djjY
mdVaLtjHQ21CGSrACFer/nBPOoTmzpOrLpb3XdjzouwBPalEZ84jTfCxO2TXxioc
PKXvzj7NAqW7//bcRF3HfMIvANyxi/MSAfmJ90a5VXz3l9ei1nZ7gpz3VrhALiy2
sIjNe1eeTzP0vv8o4lg92Rv2WFmoNXyBTCdlh0d2nQghisbJgpu+ijuNDnvC+2CQ
fWdE5ZMzk+y4OpofrC+AH3GcCpOazT0JumDvmqJHP6zBIMn0cnxbZz4WDt/bg5F6
7Gf4YREELNPTbUx+SDlY4DZ9jmlzm/nP5bek8zue0XVDqxOW9sCEPzUtsGNmHDQI
QCm9YAkxK2EmT0723BsCuN1cE9cqAoPgVnAopFV7QStF7Ewajjl99EhU6zybYOHM
eHgOTCHx9OTbvx/C8vfqdVGJHP9+OC1HC8hluo6cyo2dRVKzA8QtuGecqah1bM/C
jqG6KzTAjHaoMdfuQx1eF6ysToN3eD+XiJT1o5dWfNBQzTJQBr6gKvfgE3mEAdux
BKzHnE2FiJYY24AW9TJL2Jdn6tHvoGoR1v+a+xPj9jDgfSZ3xNgnA/noiII+WUGQ
f9jt7iURoQCq+qFixuts0mwGGmKSVdStVst/VMMKbkHy3oeklbO7eYKLkbz4HSCR
z6wXHuzywyc4sT0MIYTroNL0/8qSMHmp3BGphAqsuJac3IrbqtusR1SX3ItwqWkG
IraZjoDrTOKsaHtz4FnS9j+GVFysZpPLLW27yLki3hpAWDBE01CvTWia+8yzVzNy
0BVfisMdKU8xbQdXaj0EqWHXdMMbEQt8KnunwAIpvdsdo+ujbJPJLU65QIZxU/UI
wfp7ARCMzSpVAURfIUoY2CJ3V4YRj3VNNM8TplcPW4TliDEutmxu2OFiJpMFEzpk
1cwwbi8b9RsnX4UWlBytunSbR9UR4VIaC+Lbe7mBdFof+8oSbx1Ylyy6urtwS5sE
pdQnU3RG9Q2JtpoYzMEWrMvP88W+TwaxLUQq5wk39Gh41LbFxyOc1e9nb7+gGuh1
mh2/K2CZdSX8zMe4F66sRf8cUGNCzd1veynPaGMEvg9Wu+6aXwg4mZXJrOHVAQm3
hfYRSYp8PeYQPd1S56S6qXYTEwp2QBd9uV6ObQsHkLc87nCcCjW2oOnzP06mBImF
bnsPPZ8pT6FgnjKPDxpT1xlB9kd0du02YIabOwq5nYnQWl1mPwBrXV0z3pxzUb37
nwBEq1A5CcAsRBhIToa2F1scn9j19myq5PuqZ6qzL9exHGgrWWbTgL7gv0I5JhaI
/et31e0OgfoyJlfndGijJUGCp83tFqzzIQqrVi0gTytU+uoIR8Wt9Ec80Rr4cFJw
rSBuaVBCM2mCZXm26wmcTSPci8WvzsRQMAAHVIBNVwSVWT0lWduL6/SUNFfV/k3i
4ItrHVerE/WBfn9t8jpU+OXyJ2SYvDIk7165MJVwYWToH0uclCzO3U+LM/xvhjn+
hPHUYTf0HdNeXWhArBeSM9sgUkRGfJdy/kyfYVxERzsDi5kqxq4bhUQcZABpHau3
/Bh5S+YxJwlv0Y69lXq1VuT+9uXD9s9upsWp6isiBxottGvVya+ACyf4/hNYKPoP
CyOTPZFUq4c4QGi9GYTKANBO12taTncDMVo9ojgAMRfxgqnABeF2RUaR/JppC96p
+B5L0WV5foiqddzY4OqfQIZ/TuYB6dpandbljWBqjc0tBcl1448CgyOa2u7OikO/
sDeekg/yZk4q3EyM3vORznXnZwwcqgCzKB/+Xy6pe0aM2B4tn8vbr8eKzZBTJX4y
0T7F5WlUicIbixhFkTM+uOCt3DsfslcQBTWiyOO7bXL7rxXrCEqkSnJ3lCBOqO9R
Aj1MHY6e+vU8uY0zgdoZeZFlq1lfr16TibKaUxk1lYWIqaYCbKeCU2NJnsh+pf6v
eUFGc9z2Yg0QV1KHrZhjSnRBuZteB6iAPVCMlJhWKXsH0SgxoYscRpzoCyLzwMbu
KXv/7hiha7FksawnU4cVSdGJUKYGDoEPCV2iJS7U7CpXndIHvkfh5h/hiuC2HsAw
qAjYhmHooOG9LkXTwZBCyHd2C8hfIHb+HVyGtBdm+0aEuwXVIRt3o+zoGBXLx4fk
KbtBu5n+J89XQ0BF2P6x6VotwyOa+j0GzWbzZb+K/1UenMg3wMCDB16PApZffzNL
/3c05Jqqay5JlZvZGO9FhwQygtH6V8X77tv3SiGTCCTr3azQHPJsVGEhWxN8pNBA
VZnJv7ooLy5ssKOAnxYh0U4uOEvolBMGI7sJd0Rz1XNU0Z04qyNXOetwib+hfv1P
RUPQQTF3xeRUCsTk/202r/9vdNlJJJvk09h+W1dzIeSYwtDQB2SzxsdgMuu5tpPg
hh0s+DCY5PjKsH6dnwMpJku3mrVDBoY9Y5dMfw6FsUvO0TAhC5NAw3v6mS/a5tx9
PCE32Hgag8yO7bIOxfY+PZSJHt8RxqcklLUa4RD2MggxFgKmGSQ/raC+GhCx2gQk
SEealFhrGXAzkRImGUfHlIisze2J+MPNJ6QDiChbq0uD3qN8+RJUGh2e7MrDXzKh
F53rKiri4+OHm+Wb8h5zSzfkHYkOpsemxbr0WDRi855Uq6NGU1Rw8RpBDCeK1dYh
t0rJeKksXheztL1BCh/AaO4RQLwOvOsJRYfjnSZff3HW0mtj5G7S2hrWbL+4wq0+
fUedkIOGMTEgSmRh5FjwciL+I325EChwnQ19/n6j2RAsPWt7jqaVgnmBSb+QHAUx
O4mQEg7D7acCQR5YaBhAMi9MGcA0YsziSvjjmPDnF8IMjQCSf5M/wEa1geOrgULA
foc+Oew04cemtq9iMCyySsWnhO/3qEy+FIeZEBoyoXf7jG631JnZqh5GNpebIWMa
uH3lAAeKZ2nHlZqshkkTtHkU083GUhs27pKgyVtITN6rOZD7cZjyEYBuVYnlJWqu
9tTOe/hHN+7i9jDMMvdOKwDMEtIm2J1mXr9jfX48SWys+7F8JcdAGsO/y3dJrmGw
bYqvJrD405YRxBklgacCx9c5txNJd0jyTJvfSfiEQCyBCOruzl4ZJavOCqtPz7sx
SPnCi/CTKOyXnwpfVBB9t5II8hcRD+n3h3giYAb5PNEOgeqzQe7shrBK1WwULrtN
v2ZMGXgTFkXY9p/q1RDk2SbR6EdDsG8afIjQRrkdTxzJJfzZkDm6KT64LWbFrdPm
/ILO7lAzGsYtX4iyllbEIicd58Mw7FyuoBZWqxpa74xviKYZQ6u1Y4bstfrOIemG
KSAgSiwd70hmpB05Y7KWcXcwWWBMzgxdVUDubcx6nSc0Rxqgbf3tSaxaX7isR86r
ufjZlbEwdjG64IvBOQTErvGrNbBh6ICXD2SLb2dr4MzElHE/766mhSX6a0Li2XPo
7RI1YYJGrWC9mxtURvSnhuasJ95X/yft2EPp/2ErSuLEllPUkDPjsjNp/SC1MePm
rM6gffiKNa8a7JupieB7f2pMlnYqjDT69TducoOR5rp/GTXj0lP/WdtFaI/eGXXi
bLPRI5e/vidnT34RsPBL5ISp6FlvZdKHsxctzK/9MYP1Ni0L/qkZ40FCBoCHx0+U
FubifZmgWQamUhsQ5EalF35B55Z6OPEimcQ9vYKq5Spny4OeLYZfQiF+nJuWsz5/
VXII3/AeN16M1zcZKzOtavYdQSC3v/AVliGGZS5M1N0bG0bkfbm2w4a1H7GZv9R5
QP+BbSDttv+8uV4Iei7s/Ajfnpb0ZhQegUc6Qo0hdCa09SqjfWR+y5xanbKvQ14H
OlPQ9rXxklzXF6XJxI7Q0E2tRPeG42acmaDvYUM8xODSNA6Mi9MJIQwNPcBYtAsf
YWfYn0DKBS1gAsVL00eVv0AhgPD3pCmXNQx2QcfdVCKWkXxxWWIRhImdGj1UJy3I
HkxNxuXgY4+EsUumf8V23vKYZUUlim9YqehYX0Ul4eWAIi2RNodm6QSfTppDk6iB
eyCf7PNjiRdSePEisreIQUEdoeP1nHAqj6kKASSkcFgWbr3dZT9N7i1gYc99LkX/
eIerrPgdmoIJGV1VPLRLmoz8XuermaI2c0yNbEZzkFQGqR0goRZCR/o6vuWv4LpF
gTRU6zvqCtwMl/e4SnzBw1DPpvk+6j+C1RxZDWVSWDsO3EF/OOJwF4j2fOoloTUN
5b4VT7p5FJby0XlYrI9iEdFyvzuhiEsz5LknqAxXMozoe3CDY7mtwrF/ZTpyTr5O
Yh4wKK7z0Ei5+MohSddfFSs/yffRP68HmJld49tIF2gp92kTWRqED7x1eMgUHafc
0I4XCe1PilpqqfHdWMLCzXXfkxXogomsODPzHAxV4CuKZn4KkELEm+Xi4djNRsJ4
EG5Nl/YdNw4Q1W/WlZK7os2DYqFC+NgoeqoS58KjhM4P1yUe/w96gxG9gQpkoYtO
mKWwgkZZ+CaW5arxtgooDNqVKR8AfKKDeZVdMmcDVaUn7mT6rQTcVVoeaixgnWsN
a9tXi4dwXJBkCLXk+5DygKSoR0x8e13EBNoUycHW9XU8agkt6JV88JwqsKagy/Du
4AC0DV3jF2yZoCmBdjZ1AWcKsyjoigVl4/gXZacRseDeYOZTIgf+xMuqLESiZYzQ
174aJJwWF3HR488oWIRGR5ovRWzGFqoOOmg41SknI3wEZgzymXX33kv+OGhiuHTF
H1HPSjuHYO1I3GdHADUNB11kduZ6ef91Gdg5G0BTgRDF0eb8e28NZE1/I3Zn5hlh
g713+rAppM/79prOBlzMY1NWRVYrH5eT/J/g+5yHvMqZ6ugCJBKSCv24+b/X0iFR
N1JiF1jhgxABV+ZC6wbeksWkykbplavXrw3FmVnrpLSNvy4B12qdzONxx1TrX/df
bW2khHvCi/HRHQ4qAuOVywJzZ5JxnwTCjTfSDy7KCyP5SrQ5wIl1CRj2nbrsxR92
FozX44ni1cnAUexb3MKVOaKxdJp6nK+hc45yxJh6dHXDz/U30+t0vOtxqjs+kQkc
9ipkeVBWKmeOfdDr8GvM6u5UqrYH0i+angy56pIPGC5drrRamY/qaf8U3nwvzIM1
fdonDcn0iS3EGSqztqaSevwK8RBQUZG6d+/g1AHzAVdh5itZ75nLEXp2/EXDe/SL
ztY87OJsebdGIaEQW3Mrbez2Jbvy3Gh26AldJhohDtdsONMi6HvRFXWKl4ipDYlx
voNd4l/XdAzsBlh6FJpIaWmQk0zGXro6rKCEaSNUeskOnpgQPvgdZDx7+eVYkCUR
hJKz3ZstxJNboyYC6MAL1T8WMnUlVF5sGNWWpWp/OttTWkNMQvkVckudjUj1EGS1
BKpCeoOVjWGRh7wkeuowxDOV5lohRHLJnl+6HAnfhZfKxyUDuZaykQ+FkTwx8Cri
phLddEPlGV+RYjY94VBWNMkb2MsOHsshQredxqgw5gFz6VNytc8MW8n6SvtAl+RC
sY/20bzmBylsiib8+bynboQOAo07xzAJPA9+QMswBUkQIDLuHsOd9KiVJmSJpM18
7HVKRLYOqxkJs4p1D6tF5OgeIMd73SFmxcHEsDFiQBhWiKGusG3da8143XinJvxb
7lUjBX0BYCEumqZDL1tkE6qN2IKQfPIwZLll9SJ1e1vfoK9MGfHuDea/XG6V8fqP
a5zFx9NR/u7i/Ot4Oy1hTwpGGVNWQRyke0H3DtjpAf090fzgM7lFRRoBINfXCJQV
C/rK8eNT5EHDGFvpxD/gvoeOLHHvMZPDLU3PReF8AO2BA1CbvnivtM8hHbNQyHJK
+U2MoLVd9c/xFcnZhWWnX7FBbiG4hRaI/pOlQ6hwMjG9OdQcZwucvCOTm4lNQNDe
U1sa12WpggpVjdAfuzcvSIn0L5RTJ3k7fTB7Sxb8SQe0y44WOS3KuhbhBbeR/U+Q
G0I3h1NoucJt5utAFx+mAsJRJt7ckaLMKpUZwZNdsH+xmGrkTlnw37UmZo+ki0Ym
+egQ6HI3oH6TrIzChOsL0BIIm0YzzWV4j+RBR/qxCyuP/DLT2UcezmHiWEVRp1AG
5inJnTkNhTwKNdGJCFPNl4fvdtv7MMCdZELPSJikQA7+U5q09MjpGEGKDR7+oi7N
zIYVX1F90dTmSQRStwgsVGeP+MghaXZfSgMrXi2VolTBpd3dw7GTc1F9WU6GUCyL
glUXZxKINMA6y2w8Yc840OTK5GkCt1A0xGXKmlyAorwMaIkYr4M7gu6jr6OhY7wV
k7aE48SSh+841yWbpxyUquofdL+1VXU1UCaPMS+bMlro1xjk1tHTTzzVRi8QUl33
KMKbO/WhjJqmC1b61Cua0P7Da4CTNF5z3NM010dfBepvxuLVPbCj5bQoCfuD0XSR
0j0/x+oJso4o3UHlCxRw7Ng38SSfb+Cq7Z2h7lZH4wfWfab6P3J5YN7Rhkza5EC7
Dmh/G9AZKzNKrSKsrZUj5MjtlqYMsAJ0KCILd4oLavFrLMWT1RDWCGbI7LtU88Nn
+qMG1o0N29k14MBaBlhk9d7xLhPQGuE4YZo/oyvY+V2PgNvGWjTirnll7h1aDXzb
84Txlilzb9buFVf7PAaVEgmEJ/ZV4RCw++q2a1Ah9ZSGbjuVWLa7jo50nk0vMcK2
kfOZny3PmMTra890h3LtKOLL4eXQ2F5H2XZakMmFb10YN7w304TtPceFqzg60AHx
YsO8OWvbOJu0kGjd/c/J32tJ4UT/421CER9RMzJnyN/8O9/DuFMOvi5Q/wIIu/G2
RsMtlYBCp/bslId0CQhr9Ls8xilovODmKHKV+6f83EZ3sW0RmeYDs5qB6icOe8NO
oooT+yMUaNBl2jQkGIa8+QbcECYcw/fcwX648mxcr+EKI3aGZW94MAEEfZ3h5Mbm
OjJraR+6Cy4I+JhRp8YeYaRkuOTkstvPNhVDREfZdEuvF+xUE3gstCDRSVXX0RQs
fYTHh03bi/0D2CfKSpee/ziL5IgCam7jhP3/RFwv/GvBHn0R+Bcbxs59V4QknCo4
l7Qw7TjcL4FphKDrs/g6RGwlrZJB5GB38RVQSSNVT3REUiVNJuquASz3co0v/ynf
gqbkfA0PO4vdB2eYYfXtUb8HPJt+mBp2wcel5M5lsgtHW4cWYO95awZiDmB6IpKR
n0D2Xyfbuamm2Cc/pcbanddH39H/d1NlgJm8ALiqFSlJXtuNooDRzEdOzTAFcWt9
vM1yjB7xAxnFu96xX+08F/epvioKrizvcZT0S5SXfJbb/Vs+0R421a1DZeganl1A
kdWHl/03eATYyV0+9SL6A5WKuE8K7kKc6pt/p9GsJEyoA52dxfISWK+yNWBaFoHB
vhgQhij9mYbiwbJyFWOaNiulGb1rPHoeTsNnsi4GqXnZAECWNqySUmpKiv9C3XWg
9ZHvqQUdDJpk9p2rwoVEtAp9BUx2r0Se8eX7YgDvcbGiSc/cx66wyNcN84EHC77z
8xm8/awITz8G2a/Hxx9JTcw8Jy3SxrWmoRsT/at7aCTLgtu02W/lOi0B2lMSnsx5
e16VALyUsRyLyAZPu5XjEhxvHkcY+HgGh9IR/2Kve5imPyVzVj5HqBp3ls9oACKQ
IDiveWyQXMriwpccy7O7PdlAi3/FK/jvr9GgK39/J3E1pTLheu6mfXRTKFJMXIBW
s2aJJD5/skW6ocS54raWmPkLdiLqTf9MmCmKpFT64NCat+hFhAlRgbLtNpjJsrsv
h+ZP0qikycJnivi13u5Fg58M4FJgI1GW75dVFaLnebH2clwK0M6sGGRnus7VDHAm
L6PcxWN9NjlN4ZAbtIrf++tvVxWp6S0xk0o2Hm1SzHnNQLg43texXqzL9DdC4N6v
I8eSDCaQPOAj2TYK3pMV7EFmHwgkNDlBbrBQfj25144ohGB9QwkIOahUa+1c4245
0Meq+Sm9pk0Zvt2oN9jpflTTAsglRsL9PKrTPlZewMkstZGz5DBYSIx6C24Yontt
MtuIY9yalllEgcanBiRg5N06e8GrXqtbLo2laM+XNSOWbzD+X0HLeY4MK2Qs/0MP
b2MwGJGn7LBn9hpD3dGhH6GzTlJ00cS/qQorw1j/7SA+Ogsnab5D6Fw1MoKXa0p3
L7JzVGmbMilxAcljEXxQdSURu6JVe/R9b0GbanGfLhglEp7cw4YYr5ss9OfamxHv
AgN0D3KZ7KhMWaU0G2UTecKtnlKsKdVreFFeWNqYWvb6et0eIvErFstAIVPhVHSZ
PojFxtfHLby2MYGONX7Sgdsc8AN+QM8MTP60xBuji7qM6DB1yAyz3JXsQQ3GbGu2
DULWK0Z8EwCxS7qxnHtt17XpI9duyFM77RDimBroDDuGuNZvFEUfebzwvzRXh9oS
CyorcJgQvRcjWka8hQD8OALv+NgCOQ9vt//a01AakRF7GXJtSZ6w17+aujB9LexI
Sd9Cv0YtC8hrf2ZiKn53i8XvPoELAP3+GsJLs9d5jBPaA524jEp0Zyz5qTHj8iyT
syAmEUoYu14N4DoVrtNTESeYy9VbKNUIkwCq4oA9njlomm8Gsw1LiKqKX+JHwH5i
DErdkVqPA9aELRisOozBT6ZCc9L6+dOpTI37vSaTVwUdUw6MEy5uRmNpkcLvOsN9
PHoeeVFdIh9pEG/8j0eaMXcjzDWTT7mKXc6DZVCNIaEfiVapJHYqisWDA6D4aw5d
coSEVVxYxzhg/8PqMyAJnYSHTTtDvJQVQc7/oKgJFDpFtRHxt5C5Iu6wfNKrdRP3
o9U/awolRqpOyVwM8zOO9w1bwzTZ0luRldVhVK7CzkQHh4zULki4jRQEelA0IJNI
AUnAuxE609p4FZcYjlRY4oMmxG6Z5B6uqtnWT+DEKbIp89l9NHsgh0rwfbBbnKht
Yu1cb/+rQbz7NYxSUE054WddCyFdbhzklLA9bStWF/uPa3MxmOQFUMYAq8gQtqLA
XfR/NDY19XPZ10Ovysnkb/sI1rw23eHAqk3TbOSciMvYqFol5zuWTF/82SbUiBK0
1NLvPaTzb8PHaHQP/w9pj+t+ixoC2cUi9lew+DpCgA2lhNaMbTy69DPIJdxVUFg1
KyncYgrVGzSOL9DqePRgb/DHtEJqrBY7kEmoKQyb8ahG9y2l4MT6O8+GmcZC9Thd
nh+nimv8f4ATb6xNOTdPKlc0OI1gRshZ/3GVpt6VkwuMrEQ4oLGSoA0DTcDXBmXc
a4THAtZXvKF4DS0usfdYC6xkJSutzIIM8tcY/7zPrXs/mO9ofrdilV7BABZ+PN9B
P0D4s/W9YxBBJ9ZACTG7fDHrshKqTm6sYTb24sdJ46seEZlnKb8cCwIN7xEykDUx
FqQ5UpLqJkRfk5RdgkY92jutW+yTAp3StlTd0KP38mufOK6madQX9mEwTv0LhZap
FvmT+eEfRk7ndnvtu6kkrbRl+lL9hB7uoaD8QopudRP2Oq29lapEAXIw4PSEX1Sv
LN1qBBW9RiApgAW0ETw10lknXz/Ty87bwj+2xA3L9/Ck3tNG8GR7iQdcnbsDyZot
/JJk7hUpFs6Hu840XdPwMkAii8IhOuCZ9prBuY0/IufSakSb6fSLQizdRXezQQTk
kxL/8wkcOLcs4eMLBtgt/8FvWYLLE/l4dUuGXv60zeRLbnWhnh0ZBMb11hltjPAJ
rZV0mWhCSHP3jWpBoUy8Xl8dYUFSIDei48QvaE+s7e9MmdzkT1dPK7CsELNG1/6R
bKWkjn+DcaETQNPcZwu2Gjwm5ciIzbwIidRXSMbakUioKaOTd7fky868sMWAtYrY
W2qOeDuKoAkz9ewYcWekNrDQcSQIXDeBvwh5d9ASWniObkKQZydgoFjlLj0LG3Sj
XPETkR5+J26nZ8fLeXWJbgtDQfZXng9jVBYjA55Ya5OrJofKk6f8dskKJNwi6ovg
XlsaGVZSvbziXW/MJF9kbTUe/gxj/1zPlntuPu6lLUHTPghRXkqCRBzzkAcKmG2D
`protect END_PROTECTED
