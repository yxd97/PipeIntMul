`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Z/gpg+G76GsdbtufrajIF17Cfa9niBtR8cIRVBXk5MudKxL8ndzxCzcp/AX03yi
hOhlCF2mANU/ob9WVYILxJsMkN/lWlW0zG1n6CxQOK4B/05Dhqf4BDFpgZihLZTY
1IVKvRBB6CsucjQLlzW+kre7p8elE1TcVb4DX/ERq20qdlc6iS9RlUhRUpD7DC/P
rFbcqV7up3MFFzN2m1qAGGx95oQIwXuNmeyq4yVwFoE0DWo8WZ+xMhMt4BqI4vHw
/9a+1LsioXR8iN88e1G1IjVp10sfNcuL5U7rfslSYq7QICEIvsGnPTW/RipDSbZL
HGu6haMtmQKZZKP8CyK3a3GXm4wzR8BmG4UiIa5NxZ4WAs+WqkcNye79fySmhWGs
uogQ6n2x4gHhb7PwhBcZz0ydrkiuKX/QBYx+rfnphHPgrXAue+WtaE9Nwyha0FB+
IgoxPA9HvPooguPrGd+v2gUdmBUgX/RnIZ4MJiWhNz5ofOF6VumI9nFK1MwcGiH3
bjHBsxgKSKiW9u4v6ju2AClG9OheiFdggrxEUm8DRtnneS+jV0CktD9CXPtWq2Tv
4oZmv2gsGHxHT2gD6qRd5zaIBF5En2LysWpkc5i2oEo=
`protect END_PROTECTED
