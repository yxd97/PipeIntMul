`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xr6fXt99AUcVm2C1rWxwfLofp9E9ZzH3odlASv5CFlC9yFDahEIbSPMnFgdc+g/F
Ogsf9skwyU+pnUvv2pwqTEWWqEaYuy/8IxA3b0JXNJDuP4u95VG1zj5iO6W70DY/
qa8ntwnXX6imODpF7Pei8U5x1BefrUQGQR52mdol7L/QMX6Cbnf8uhjTSnKCIUoa
V2T51KS+Uk8gcJMuTaSjFYH7FmDYepqjDRbUgayTZvPd85Czj3lySZ3mmr+wTo6i
lUOZsy9tM0M+aQxLcha3xGMcBWTZ2U3KLQfksC2egQjfUf8nGfExLQk7hVBoMnX1
G14OblQKNxyB/Y8SnYMmtVE5kdEOJlzkpVV9emwuD1lrcftqu9rDRQDX0wpMUxlb
b0O+4rVwgP8XminzJjV9qZ9avKrWSOQPxqvmZwDhOzQEoN8ivq8R/HoTYDpHirYx
ZzIWH4ByYCfSujF1fCxYf/lt/YkQ50X4GhnzwcKBaxQj9IlKMCrjkrt47UVILnmz
3WICzb2vzxDNHUWHnO8BNuJPdfzwW0mH8LiX5nRgfE94NBXldNaEUkkMJTER7BB1
i40aNren0LWyHD2R79zQY06xBQAV0mstboFYVflcn84Brwef/7OyuhpUgkQlxAuQ
p2o47bm8KYir3TeGGE8M2XIAhYZyeEb1UoLmpUr0Z8FlOumC5qlg3M0y8MKSiX9E
8P7/MLMdsTVnSMpvr54cKvQfSP6DzqSiyOM+NIj3bOU=
`protect END_PROTECTED
