`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KhMoTe+X/qokDv6rkL8VSDACw3/Xm63sU4bksD8NgPveBKyfjwn2BJrrNh7I5uMI
x5sxLc6TXs5FTTVeuEXEgJF24d8Ay5yrSyR2fds51Z/sNbkP6XSOK0NTWqNUYUqo
Rpw5bFezEGeCUsQwoF9FbfxgVSKnOCRsGxR7RC5XfFwXdQ0TkCrv2WoiRPHaC2M3
XtcbK3/Rj0m5PavzxMwlOs32w4YRM1e5obcdA3aOB4J/P24mzizqxl9ADfBCezsy
ZMBSCvI0e8WU5ZU8U29RtSj+PEccx/hIROmVZrKkzCHnTS351bQ3SAUXw9jItSwl
XOiabDAHwxxjlnF7MCXnIPWtH3Wz1KI6zEhhSrgKD47De9EPA5VMy4ycbt8nAZNn
RxY3Uu6CeaWAd/gMjUd1fOGpDdJpuPLahxESnlQg0S0K61AtjM5NBJUSNSkV1Vkf
iJa/4R/S0PVSmGrbwEcNtoVnO0m8WWBUxaKCDdFkDn3bVF1ghrBPawXIxHs5j3j6
FKlidSgxh/IBENrEkcXKD2ib62DXBvrZsSeqccD7l2zgOomSKOVPo3/6n6eYjkam
9sGYX46+PPWuyki1zrRwyDDm0oSuzusSQJ3inndr/hCQ34q8a35s7FC6epIdkdm9
Du8W+Swc8opMjc5zfvhB6JfKbVr6qKmFNODXAbRnjokTqa1RC9aKm0WMZybZKgGV
`protect END_PROTECTED
