`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ebek4186uHEVohMEOrfUuBPUyKtRljsMP4/WGlDGEwuWi0twx+B8c9CZlWaB1eO3
ft12tgR4yEM3b/Qq940yUzYBnDlZF8qNpmvFDErnb6o1jO4lgx0ksf1gg8iDkb/8
u7aV+ngVGUMDjgq/+NHpA+hIUs7GYvGdLU5C8NckudGIJv/7KjYQGA7iBizsMjI8
91oU/iv1ca24wtQyjC7pKC41KY0BJ7XYdUDw1P4GYsCTMTUqQX8fTbUyQp2a2+5A
0qwF33TFuZeViG0u84JlWeMeCWAKzcdXCWoP3xvGtqt6KQhthQubthYqgYJhW0VM
3rV6E0zd3zFK0+ufJd+Nj1uIWN54yv8kJ/EKv1xETPSZbvfg3bJr/Z6FapXxx4KN
iRpsHkmho3HCIZtHWmSOfEQXYBLyuAZa7gZqHCv9DpA=
`protect END_PROTECTED
