`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tZWEQJvrkHoSgF1gMwLdxZl6Ay1vtGQPiDwtWrfN02ZV5akzfpyfP6TFo5hvKlGD
ILbfj0FvOZamjVvrWrvkZupHqZmAcOADFDWk3sa9mXf2mtfpfsWZPnFOxKLAXmDQ
Uk3213O1g43Or6q3gsw67TaDANWyimarciNmk63J+pxs0saoS+cIt+jDqtbaRcKz
ho31uq1XUOFwhwdRPAuT7pD0/oamWgeoTRPLsBbEQqk=
`protect END_PROTECTED
