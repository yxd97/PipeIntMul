`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QrqbN+veuqjYEcDmU7jImSKdExshe3YMLdRo75zsr5WgsOmPO4nGPLj7lEI/c08r
e0hATaS/NBuaa0m69QXjls7ZqAMbjlC+vjorSdF0CobIAb9B79zTjVr1WUQWzpLI
0zkNXQwAMWY25rU/bmB0Bv1SaGxiCALeXWOmbWWxBm/384xzvv7ijljbk/UX5a/a
3DYQLrwx+f6+azOKr2PM5i5h7+OZ2JpzM1Q0bts9HR0AGFQ0qOu7oaMmjjIhBoLq
n1pm3zP6HqaX0jV6j0I9ZYhyYMbgjjsTrafQEdZERySeJOHZUnuqTSjjq3hd4HlW
LZYE272c+001Yhrqtz8OG3QTYNC4pOzkUNpxNg/7Fb5KBK2wiQL8GMsb76ChZneA
ND3lbs9jKnU45eQtVsmfkJmRhB/HotCv2EPKYmVgVylBOqxO5ATupu2HLEXnXLsr
8J9+QWtSw58/TldNCuAi1w==
`protect END_PROTECTED
