`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DtIyrdWOXFuMntnfsF8zZNKCIwGrwDYopMV6y72pIxw1cfVu1UpXyRWu0QA9+6tP
DflnPWgA9HSYzYdEh2R/ruCJaxAlSaoxM/NPcPQxl1JSKJ5rNQ8Fnkdk52tQdNm9
l9ryXo3eJUYvFyVNeWWqOHnWD0CXywowP+LloDWO743b1TDxOmWKG5nsd8MMgxm7
G1IktOkfGIfxlXZLuJMxKF6thoSgDV37UrdvdRbef0feQM8Ro5PofWQg3OQVaQZU
mndXj/ACWZed7qZ8z24r9wAnosD7igZ6yu8wXBCSvUECECj5G3RERNK4mhLVwGr4
jMOUnpoKAXqFdwDcE3LzJhE5WZdBpvkR/BcxU86hnwU4dDSKW7LKdxDE94Jmxq3D
QB+OslH8e48gzpHCa4RRCiVj/UhRYrf1U9uGkzNwSs+syyrrNn+DxXgP60rJNsPp
yIJly+lBxXiVeQKztxQTpf5MazYzOiAsptRl5jedX9dbdEsxy6SQnvTNd/hw4cV0
PJJfFniupbD4FpJNrEBT5OFgjl50s2Dh6HD9Rj+/b/DeeLGLUlhwAa7W+esM/sFq
/fxgYQj8SFgoGGCqIX+47HnHre+YL9rjev7CvVPTiYh+oRDJH67KZUgaumkNsmuZ
HWKyzYSacrwy4wiutwiXPUV3DnkOjJamanYw5Y8Es3LsHHdKNeaDeLDSjUCdhvJD
A92TtCvnq3oLoo/RkQhaDDPPLNhYadasDxzDNO72nZpWjnB1HbiSd5rYaWWIOTK1
qDas4vKHweI4WtJrZhE0Fg==
`protect END_PROTECTED
