`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZmPJ0uzeYZkNOxuys7fv//zKzFHwDbJxVw8sFf6qn+3JVUc2EQ9nMloJQ4bkmdVv
D9LlqpvvsntkUsyAlbUW9iKOIWkfQyMCDEctWt+/gy3LNbB7JMjKOoYQyH21oT5t
41mAnxAN1uFzX9eswabBwQN2WeStDKQAOQbsJZXWTL76X9/a6UzcngE4lzozaMKj
/H4CdGklzcx7OJUU650LnfS3Pw5RZThimhXnpK7FCgbdqsZASaIhAWpKi4jMUFGk
FTz38VM+zCypK0mb896b70h803A4ujYIq4IRHP/7tDqNRWrT6xb64LfuV6zYRGJq
r+P7Suf6sz5BwlBRtTGEYg==
`protect END_PROTECTED
