`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rg6kB9BG69hIJ5Ta82eq+EZtuDqkNgRszHb8SmJX4JDR3lkrzgM3Gaw1oV7pQEn
QiMuKEusCS1Bw8BREttw5b9OpxqAWfrxyeZVyfcrGTOcPvZRSC50rbdjWME+i3qF
6Dc7wUytq6LWIVKD7iNptGMG78Cxpx40iGxpkQ3lqokFxUuBWP8a1KvND+mPrsaq
QNJaVyh9hlE1LlYRS8ZwqG1x5fBbFyBaOXQG0qgRyQka6HgbyzG6tkRZBJFFDRYt
Xh03pnQ+uMlxV4Caq+35tXcpBtl1CXvRh2zzM3dMEdhES7ufsXzSTuIFs9s8Bl5E
sJPlHyWtWci7wZiHHAnfVTZPCxmjx8fN+TNvOdZsFPkaaDErPkfBauN5TlsMQngf
pKsjpSfWdefqw4nu72m6sI1rhmt3W/Gdi/bbmcNjivTwLOrGEKvgnKFDukPASqdt
P6DBBSyZ8/QeCWTKPLeUifnoOFn81tnbVNe9KCA/pWI0n2riQz2F10NpXafBuf2s
aV9lFHvOmH+EdG3jvKS1sMiFGRE0OEtnffo8qWZLNZN1puEjZgqwTEbqu59G9sh/
SGx/TYn00/KjJX9rJDGrQMmm4pyEHAtJ9koPznojhTfKaKwELv3JPrFaJKqQiqSD
sCXVSsmZNJMB2h2UocSU0ow7zYquw+JOK9bQ4yYoQMMEVeMPiWXsXA+sUmcqyiNj
+MYcIdd7/lvLtREwrpkez0uNVkx0IeE2p4wqJc1fuyowhhNxsqYYPYMMk7m4qx72
j6ULAwMmz2QrGnfnxQorgpJ7PMeY+0kyEpM551lwoWnsMfTvpirFGS14emXgnocP
YAoSenaduZqvqySna/UvDXC8qg6dnGX4BrALJMfUoOS3503BQGYzthA3/B7ps+KX
rvIu9Y23roaTjJKmYBY+x7zncRRug6CBeuW6a22deXvJGAxPwpc56DUz1BW0M189
sfAGRmzYbJws+P36/T5eDQ==
`protect END_PROTECTED
