`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ELwdsP4zw27z1E0lkM/Q4mY9+BYeziWfltSm7pTDHRMGw9G+Iu35JkO4TIWLcVOx
Fqqv2EYKmPgIkEliQUbQ6cmF76JesFQL7/rKzF1WrP0sGy9Q/dYqBWK0P/9Iy7Wk
LxL4QVl2ZzYTsqUKMuQn+1raJBihXRAvAT92xxZtlL13b5zJLsmNj5qh4KKwfFwf
94wNhm1vQYNm4yObnI0FOU+QM9XgZVnD72BCH8UyEawsZTTe73zH5hfMnd+QD77g
7vphtXhQhfRF+UOGQVq81UaVtH3iK04/B5QzY3mHTqu0qhkcLXT+5Npz5Au1LYbF
7UgyUvASO77GF6/IFIyPz6u4os5pTCAoNRc8JhJHNXRcezseu5WNbprk57jWcuBn
N9XnkkRvfMAVLC/6Tbl/CxG2elbaY28xrvsnmJZDafuDIdFdse1r6Ytl9/6+kHfi
MyL5pDV+Xt5A63ZpQGek0Tx6IlVLa13zfpqjtX20YIlybYmx5HQC7fAxoT7LfCTh
XETssPrEewdO5JQZH04psW8Z0GqsbVodKBwWPaBy477/txzzh9wbOEvyubsJy3lK
G9gMgwyjwSAI9pA47PWXFdEaIyz+rfG6IvXToGfWpJMTcXTEc9OYDYGrEUFDYfV6
CfeWnVXcdU/Ad09sHS401Cf5lWbP4/ETAhd8/M43Q0fUp3qnr30cvdrKQvx1DzKy
4JeS5eZ/cdZuUEY4ZBKya33wWrJdPr8Eo+CJPjk1IM0MorUFbiSlvruJ6IW0MP4z
Bgh1aM4WCSo9Iq5H9XbtBgkYxGKokeiQPI0Cy7W/0diewmplcoNrevbd4UPUJ/97
3l7hb4aTkbjF2oVvV+C8c5/I79OMjQu4ZQmvVBJw5dO+9hVosJtIysdmq9suShxD
Ruzn58ebwXDVHRRnNrE9TJ66o+rk1NRoSJsUBd3FaXhhE5EGNkJxGLTvJ8uKghPH
6YFt6Ht13awC0k7fcUA6THiBMaSWoI4xQ8QByZvKUKZH1TsnxN+ElYH7bmvAAykV
/3dILLlhxo9magwNvOqz44Waw/s/2qYMcYhjqZ9z1V76kwjpwLqe/BHBQ/z0UgQ8
vUgp6VdAR9mGfKylQqEa/QLgKoLIkComoZjrSHQ4XhgBLusWC2ud47wFl/CXBmA4
ER2L6i3fxgqyQycUjo6nOiyi3Y2G4JLSY1yvZC1/oMZQch3AwVKONIkvIk+/LbYo
qMcYxlnEsmlfvrICN7zzepP8CulqArJVrI+SfqXMt7MWscinFua3EElJmow4Rjbi
/I6BRmiLDTfKFK5yvJBoYFqgS8gKg0eDBl6LR83l2og3CbGIuBrBqNNBdkbmFRcr
sK5OGDjgK9DGgClj6pnPgRk02cUQIw9rRA9KxEd9cdCrFeTNjs/gX4eJPdZUMxPO
GoLsEngqiMXfksYlez+dDoMwNZySlmaw1w4ttSi/NKqbp/m1yi/B85Zo0Wy4blVj
XaGj0DM5LmwuU+0ISR3WhTQ2FvCJx+O8Aiat0IEKtIN43X54a/XU83CzGOyNN7jP
kPae9lD4N5bKVXSsw38e7T83838nMcvShB/PsgOKly2ah2hSX2qlkN/ry5ZCnRwi
7QdX0pXy9tnIiBe3AdY6IqADYmjyzXiJygxDgcFTMVt495WgXbz2oAaoikPrtmfA
X7QetqYryvwh4GrYybFJJ/Zq9vLJPGKXviqO+MHt/XhE5CqkA2iX9M+DUXB12wxr
AMoEoYKsiqYANolxnQdau29cWf8h2TdX7tYXUebT/HaNUADBAC1RiXmdzGTVjLMY
GTaj61qo8W5UG/qVurrtH3gFoIhO2yEWIR6HvMoodYUcT6pr91lRQOgbOO9Z6Gx1
yp0hLeDVAKEGDK0BqRLCcnHsLorvMi2Ze5jSVN95ZOxcRoLq3wt2YBoODuQDC11s
jl2wFfvqLlwvv3DC2rRyCpZ/Qt3gaUhEwUAWCoXIc+F/ynoKDCdf1foFi2gDqKjI
p5nJLi/jp+8+eGhLA9zn0Ry4GF7NzytbMgkODzCkrxgP+QHmMAUuQ1VdRyrdOqof
5w31RH3CuqxIGnMsaBPgGPXfSVO9vbsVnvuyWSyXObK59YGf8sHlpOnQqUYVmdWl
8zQ6GM4o3UKsv0uxZDENkjjoZfNG26xFQ/FSRL/uclninaLCjluqugZgBzg2Dp7X
SGc/x9RzcEHcAzhgLcHaRA8mtAghD1LghsTIQHP+VqNxm8D3FHJw+xGpN9As3Mhd
qP9G+TBXQ9nXI3tBsq6S2CtbzxFa+83kl1CS4M7yt7P6DRiGI7A+vEfcNOIl1qf6
OLS5+bByCEXweTBG1Hqe08oHepGuibpmpM0xyV4WZZ+IQfR1Dim06pEpES+x24Xz
mQJnubVTSjenJiqum/4H4KrpxlL76OvcP1Dnim4W8FxBP8uVciNkg4u24jd8IrN3
r6UKUAHlEnIZElTauVjqmD85ih/rEn69NSLZNj79I5Lk0iO8QkSDDfaRkZn1JoaO
bgfAEHR0UJijPaBJBjkQ5pGhOhnD9cBvr8ER8mXUOU2FmWOi9lqkOAnXGRaOtzn6
OqjbS/lxPQu6UF3kn1mnBjbTLTqEQLu9JR72UGsy0C0Wa2zNo/DttRV9NJh/yG0B
OxeVJc2WKw/cBhVjPLuGXMfinw1v8qVeSeBbIvz8zlSwvvsJYeC6lgKQj1ysZh8x
tRJdnAZGpjfaRPh1IeQrOuJ2V+JaGP4pp4WISCqn1TYqLYX9sPZPOi2pFw/IySRP
+X4mm7c+9dlafM+V/MLio4RdYll/TdZmvkgy/qiuRrajhgYtIz+Hgu8vJHFDkz5z
RbRHrIBesd5i4ShDG9W3dfCGL/Klsl1OlOUj5bl9yw0mzots9uFUjWwSHsPvuDnc
563k7q8oV37yPqWuCSIvr/Svi13GPpVi5SAFtFFPUtce/U80KPNzxq7zfjyFuxWE
YqOeVEj/3cP5NOv3+NfND5r3b5MpuucAPtY0ZVjWCKz/iNvVRDEQ+vT4ISAljUSR
LZZGr7drIU1EjSjr5H4CAw4yfvoXSHOoUpygt4A/2Ht2LfxdDmnptV8FmN1jzRWw
eUJj9l2sYZgFeBE8SYmi6S8ww1MhAIWx4JEaoguV1zTheKSDDF1kt+bP7VWunMNC
S6jCBP5/wbcB18Cazpa/T72+P1OB5tp000GnF0R6wWWJXX3k004M9uyrrzduzNVS
r/xvP/mbZycBRRRjaGQfo01lFx3iJ5bxlju6AM50VjBwvloC7HB1CH6OrM+ktFoh
wNvb6Zaf6eMHZEmBL08K6h9QHh+e5WOlOg9/iPRFRBKIkvnKnvjsxDtj4yJOqrZ2
UqhKPpJ0iRaZ0AmJxajzZFkjBZZ8wl+fsH1frLjz4EAyeFlBv+KD+LF5Q/Zw0lyo
hePJZ/kNqYDa+kyPcu6Z3NHOvr7wXbvcZ/gULvJMHQ5+RT2Y59PtI2qvAm4NzyCY
dM2zuMfjlRblUwOhyv1MSS+93dLJTPPeSrBsx/pAd1eASGaw/O0aYI8MB87hCm0v
OnZI8mlUVTq2HjL51KVLwRu64fLqTA/yRmeBEG4thz+P+U2q8TM+axCbbT9UHFmA
6eubDevDzQ9iFVrYsOH3QITdDyl/wmcbVmqTLY4PQImGWVOTjRZbEFH/ttsRZ9vA
FZmL0Ki5MB/OoN0uetPSdEbaNaLDMZscemDePSyxqBG6Sn4XWfD3PVjQtjgrS7Uu
GqkNEkg/85rFQm9qPMjfzu0RtyETauU1H33qXnyen4zY67y/tacsYeZDy4K10m9e
BUuSbEw8c+QM29XGA+iO8Td/8FaXIRvU/CHMR+qZ8IibMPuLsWNz3kbyC0O5tl/W
IDiLn0fguhzZdve0/leP8p59b6KVmFoJn2jerGufVs4naB/5r3nhB2jV5j0uBzoP
0nwuvZkYALyKMpaQPXpWPE+2PRbNCoYF7TOsr6g82vlkikXhxj0jYdIRwzyJ9u5p
9daft6sAoDNh7LxuOT2Wk4aYT90J2e/fAz/Jn2ijtHrYxXzAUexaBt2MQLVqXwnw
aVRJuPr8KT/i3gqXUhAGzROWX1Dag0D6LnbIuRg01WnfRXbuHkHmQrdirg/1ul7O
AIJDO1lRFT1vT/rr2JnEB+8o5inQKFuHDyoFE2fbPj4EpB2hf90vC4MmOk9YEocn
TGwhDB4Tba4bT4pCG76nLkfT6K8RV5JZZWJ0MVYIJSw=
`protect END_PROTECTED
