`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
np4CLpTzeCxQIf0IeHlVib+4i0ItQhb+dB46TKKvuTsyZ6AA1ouWrkpQ19RrLAQP
1VGBCwbzSeMHx9HNriWvB7GqT8qt5i1/oAEB2ANo5AyJweWQljJRsiF5f6e6mWuR
KAi0hV4CqUGxuiwJclsMf7WD63hbtEFY4ANUScyAZ+W/TYWcM3QD+wUGyqlQ7nMC
vERgARPFBStA03MbfuSCsAv0Vd8TVuXjlfSdsER2KYXAqHUeYU/XmtTRSvZYqN1Y
rve0w1MObArczS/paRSHBM4G++ZW9iSrH1NvdkEQhFYijNBle7UIA6awKfgIASc3
RpYjXtaR4rM63bExCozhIi78DsoBFUPU5WB+aHVcYAAVmKUDyY+X8uPsGsqAig0z
jnuIc6gR8JSaH+/a5rUH8VasijuyU1K7LZeCuumYhhvDXKIASV+1OUiBrrGVnmAD
steppisz5rWJVWGhF6dHea7A0xiREw8Wrv+HIqEIZ2N2E5pVY0CnadF093mei68j
pa/YbwcsAoCelDUtjy1LE6miRyZ2OgRlPPpRctZPRqswa92oQDA3LOG+I8iEzvCj
zqdUIlopJuebSRh+RR4zStOL6KyV23wX/Vtt7K6zTYJsxbZPvKVljlRNUUzqOGfF
zm8IUl4+WkMiydbVKNaTNKStzMnFHjuCy0by2TtVa+7fACKkOxiJil8aNUi0tJtw
rzqF76ns2K4j6pbkTzEyBJKTRMTOr4cpRZ4nxfecqJlY0hcxcBPdHpGVSwXrZonY
TxqCSDqun30jGBVMqms0lkZD9Lx2EsL7loZRlG2SqYU2UowslVn5gT3coaAg6bmV
TdytLOIXjo2omNuVi85Sr9dxQXSkbsvOsn9Z+rXhx5xOjwT6obLmw07vXPISsZ4x
7UqgL8cWerF3Z4fTTrswqFYOhF9kdfqws0XuWMOAJh7KKfbn+bC9V+xaJwvfe7U8
rYjrcaEhNzpX3a7RJp+3YyFexX3ZMsiGnYWzcOn33eZwBaOF31s7Q9owpTmbAYwk
9nZuigctD2C0c8c7Pv4gf222SmWf/HqHbfsr8UkrEgpvNWbHrtYQMu+RKFk42wfX
fssjgXwjjpsCCmA6lirilfD4IAxTszn37oNXbfXtDQEuWubpXUlvO2LIktFJNoHd
47lL33W9380jdJ7qRuHksvELyQVMI/P9cjiUalMUBsGKT1Si/DxAEZySmb3A316s
xWM8qfU3D5OWdH2+W07UegJMW1OXVVNQcv5holflO8W3g8zBREdRJtAvwBlXSGc4
Pp0nolINO7XUlCdhO4b85qKHqRVx561g01Q1AcDwpzdIOzqUWwN5VBFtwYJtfGwy
qw1fjPm57G6hXfHXOUUaJ52ssfuYsQ0U56AzeaxDmaFmc3BaoYi1Ep+zrNSUS0qJ
s13WZI+K/O2godBlwjN1+UhCZc8ooDg2VXi/tlo3/mZFDbfaeAQF7+IAatrHtDkH
waQk0VnLytPDB81GmIDpMAC242gOQ2IMInVqeHMpvv8=
`protect END_PROTECTED
