`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3+AmHic0SK3XX+qKA7HAUvyyqzBHMH/Oyf/XaXibD0GM+cxzG5XcjhsqiBGNOp3
jGM9xq+jpLSPa6+h7ryfi+8Xd/AGfzZV7l1nw7hgckvMXAOOfivZ5a8QtJu9k/j2
QQtU5zdIRcrHwe+qFVEIPU1mjuYZnOuT4DzCA+nh1xb6XkMT6pn4Onxc8iB4XROT
becHCF+cDAco+3Dc2r4LAzo7BwBm1Gw9IkSg0/iTV6XaHNoKyi9g9M16t75Vldfm
PBaHWBxMFFlEPkxA5kDC3fyjmvh5B6rJpu93i5BE7GV06mP0meS0Xh5pxbx6lZij
3xfW5AGjJ3Rm52XAWMeaFUwMUq1NA7MBJXFvYGaB40YrpfHZYsdk2khkRTRx4pFx
+Q2vKKq8C2J++9TsMc/bAdH/gm0uvYvZzp9uSbEZ3SFgiq7IQPI1ZycDjS428qWy
vJIqFRHvSzowlHubBQ7PGYMeqGxa+tmJz+XdqO1epLVDHjXSum64X/2EZGu3BjvR
LM/uLS+YwbcX2WqCodSqJ32QaSopyh5Zf0sXrMzQNaJ9M8sbSLf3E9uUQnVrsQw2
o0q6Fix0lZ6iCa7UTwOCcJMRMIpw1hOSsE0K09v7EjilKhp1HvgqW9qGkLvxOtW/
MSRJRYWHOGlsuy6VfEws/CCIvjxeO842tOF47NQZMbldq4XvfwUkiR923rWpnic+
le4l4TwjgYQg0C3Bca38BVJfpK2UNChDatDM96J8lV00/NoE6rPp9qkDvRbfyguL
tXmm/rPBfzS1jHwRdZ+kc7PMDdIXcnkjnchtze49vmmLrUlZxBH13FjdZG+vaeST
HWNiJFicoa/kjY/sJH9toEq6f82uw27Xv1n37TBlKhY1oxmoBSIqjcChWgQpzuLw
VaShH/ZAFQkf13N+yZqWPA==
`protect END_PROTECTED
