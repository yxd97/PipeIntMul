`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7sxXp5lqxGlV4U/6j/fYQOmAmJoSbAN5eOhdqElq8QU6/zCAMmwbKD/T4kEH96lN
NY9kYD/QPvqecaW9O6OxkgZbrrLIk8/3rytVjn5qFCMbQmFbdUomk/lAwRfUcmjt
iT6mu9n/sA57cVUqbLrwrUyaARes+loxONgbMwRjMWOhJN/0XmA5ffYoop2HA8Jg
U3rLAw1u6hOJ7ASK6RMqLuEwlIAeafVPnwejiTO+Upf4/0Y+XRN8uTMkNKxyMnt4
cLkO/CLzwTWBA5nJVtSJuH5CCJCDBfLlk0BHksXJd/whQN8oWBexmNhMp8vRrgmF
0Qu0PU11gxsDD2kPuB3KZDKsReMUWdGc4h/E9aN8Y4k6TbvzLgu3758U1K4bBb2Z
aQerChInn2nLQ3g5jJ6aKUzL7CP6DUL7UChmzuP62aNFRt12niUKYCnoKpgK05eZ
V6+z1churzdyY6sPlviYCQfEh9hgx7aURkXKs/Jeq39idLQ62dTaVtcxI97+Rs2S
pdSIGRBNXf1mKOZ0hpmFE6flp14FAafctqYWYjblxwkvsVSlVv7iKneOA6LTiCCG
vUUSBs6wCHPrDL3i68U7bZkcQDe7mjHqYNluUulbCpnOsHAwFOWmd3amdYbKIB5v
iBqwQW16opsARGHXdEXfgJa8e8G+Lh2ESIwnh+WpjOZ2aBST7RBJWIkkl52upmV9
wK4pOoZ5lRY7MkTJU7llelhio+WoGRvFNp+C276N/RRVnAX87e/1YR23JLoKMouM
+Fe2AdoOFejqjGVmOPlb9V95wR6i9CE7TPqh2Wy9NZgvdI268qvKYvPEj4V/VBZ1
/3SI9Gjoo8d8khcfsc7s/WATwfHAUZ/pxXoDMswVfMdaWwbR+pq0sn99o4ederjG
ovJee+5zgGtpmDy+wvF44/zuUvhmBASbS1cMe6jQw6I8LIwQwVLF3dnQNTVsVY01
rxFtiOFiFMNIU+pwKIJD+UQ15AqIyODWeqi5+nf8ldxNgqSEd8wS+GTvA0Ww8b5B
L3q8hyCqyDmyupnhVltN+Z6IodzGQDN66VdnqxiYqWyRe2Nh/kj4AunaKAt8FN7q
FiRJcaDbjBYTB7ShTi+m9QZHU66kslPXjCUXGHnUUFhqtlglQ2qvzvrR6C2Sxkjk
4gFT2ERVZPt2pxrNJFMkRCwKmdD6j36SRzp3wdsl+P361IMVy66L8Es87L9ZtMYK
Ofhd9f7KATO4ES5oJNr4uudPVzvLYlCwBVATQunTO3yMThg6ifAuY2Zhxb65z67+
0enkFv9rCedmKekeJFSi8A4mU2DPTBbJYOvB7gcOV9dvLvEFTliZYznAPINfj8SR
euzphha4zdKkmo+WKiusD8NLbUD6PheSgvgm+qvHvkQG8WxlhlGJqRvC5IuQMyIl
2I5YQ0Ta5cE8ciWCgXsJjXvnV74UKkgIb9jGID4kXuYCzHbDE2WM9AxpOon5Q1Ya
beVXScd+SKPq6akBr+e/G5POkv0jy5/ocpwBrZruom5T+JOmaTC7j2PIFNauexG5
euPpsqQiVVwwbOfua/aArcYMkPP7+SVtAb/w9Xj0pjP8xtcwRhlW2uif64MeWavq
GpAmIUEXIYP8szIs+T7pErXWypVpTtqv5ggDp3aXNWoSfnPQY4IMZhdrWl1crc8t
61vckX6m/wjVQ5baitAC4oRcErEyOI+kXOC5P4H5zbji7YaODT7LJl46Yrm2F78y
GWNZYdspRejbkWxzafpgKFhmObX1GDO+3rQXeIg1GdvEnDIt5/tR+itIEQ9JQWnQ
SpcVNDg+X8kItzCpmfRe+5Pjps7ueOL1h3HjiCAiefhDyMzE+06KgyoDAtE3ihGl
1nHXXozfnXGFOkP6ZHeD6kog0izz6w1sEKHDIMpoiKMxEEgapVA7xzuBV2R/PGey
yl5wjW/hd54tRe9eZym2+we/hzecGaSDT3L786LiYGe4RzAGxN+0my+cex1XuwQD
A/T/3ZFwI3xgG+3w/8qVWbHmDhmDdXCfLejb00xVjKa2ac2Qal+u6SFzUsiZSX6m
I927KODvAzeDnXVOhpd6D7GIIVo8SBcDsVt6AX9oKIQ0Nl6z8MCfEK6jnSig9rdU
AMvplTARg6zXivdxn8pahlMc5mdUWfIbbZ/bnej55CnlU7jJyhazdwG8hGW8cZJe
nNp/QsPVvngqEjEdBHQ233J5f8tHUe8mkTewdSLkLIEevFEG5NvxIMYkMrTWSibf
XT01q7n6y/ooKf0+tVUVi+gF88iKsNzj6XDHYkhvjdPVFo4VJKBGvzl6wIPLAwQs
SwR5r6+CnnltJLHskL2t07UIaHczlSFwecDCL5EYG7Zpvhtf/Qd9iIzLuUsODRBY
oo0erzc9ES9mRQnp3dvEoNdbxW/8oVOifs+spWjyk6yWF9ghFMnQDEg/MlJxW0wZ
FTC+TDx0CkQl0lG5HZBzkXcK4ye8ksQqoebyAM8NtCvCXhflqJfnC3SU1ggHiLd1
crUg6l27nOr/RiCmBkSDGILPbIzI0jK3kW8kOtkULgPX43p8NwXFbW/+snohJoJr
DqXzuR3iiNH63+e4EuAscwnEw3ABmqvDAq3W1vJaptmQNf+ikMltSwL9kF7sHB9M
nZVbGSUgObgorZ7hHwuk29ArEh3F/PK+Zs3DCEom8Z6AZQ1JBVyQIhH8eGmUQrgt
tsN4Mcn50SFLLfbsghUekDVfY+6iIfuhL0svkQzKRbQ28h+s6QDkATK38Ya6Y2AU
CMIgmyKRGxJRLnABynVww4tgG5nPnnz1Px3F3yuE8pnuUlKoRgmRAnSZaR0/RfN6
G4QSH0YlFEGiIQlOpYUUxb5LSd5CHYXAAuW8/lHFCz/PjxJ7w9+Rlv31O+VyDray
nm0AbtkgW3Edrwqpz6xHPRyelO803R4BD4YUxUKK0FeTyoTbt1CRMDZHlbA1sXIa
O6ym9x7hHeQnh2LY47QdJL8Fwg9ePjcUx02lTX8Lj//GTuNFxZzPbnr1pI5w2Zc0
+aFx7m3L7mQdzxJblTxo6cBO9fI9P7SVDagdz/Zq/iKgHdOfxDyiD37iTkVWgqVZ
Hd5y/0XELtipIWwB2wlQ89hQgOx+aN1Hht2szBJAcaysTvIxWH3T2gnm9EqzlSOh
DfzdKcW/ymmIe2R40GBNxDrlCeUD21i5HMVTFPvtmH4IWOarieKCd1zaAu1H+qs+
jIgAOEL7LTDeeyWX0JNDmwxA/4bURYkuQON3WazL212Q0hlFomV4MCXN9psD+x+W
fsxG70a8Nt7wutN5yEUHBALTb6ZgHW3C91KsCedCscWJO7nNv9Ss5mxymb0E2K0f
R9Uiu4VhIsjvGWIqka3uXtn78MEYpD5woVEOX/6fi4mJoPaLzXUAJ9KA4DcJvwaZ
8iG0vM7qTc569LI6mzVePgUu5J1L+c0jI2O5WabuIPBhCcVVFUC+EB/B0QozUgUb
Tdcg8IDdpPJY1R5iuzSRDbAYdqEH3sWKDW4lGqkB67MRvHA12ApFbZ8lWY+eoM4j
wr5xWg7uPguHzpLHk014oMRJ0ZTm2AAmdm8O3QURjmAAF4hBInobGzvzZNua90Dv
CzKs4UcagR0G5TyId8NSYzESmMzvv9dQzQkHwSV1yiAuFv0GSsk6ZZUBAOo8j5Lu
7elSoOZZHDGK5x9n+KYWvumW20EqCE3vhiXL+EJv8/enHsgLDOaziwYJF5myxVC8
uSf5ANb6lhJogyfRqvN1wcLSa2psIzNJLqs5RUzvVfnFN/gViGUxeIbJ0KKUGwM7
uuS1fS+txKNCCEbLRaPBooD2dHgdPlMrZ+ozmHclqfIywHjK1EK+8DM8omUR59hN
9ohdCppWJ9VSDi1QQpECcqXEcNvuXEixcdhGTRV3Mq6IXSMPDVaCYSB4V9u3QhLv
otCC17widgfpMlPxsMRWVXSLx3cuHtJyQEYKMwH1+ieXBrX6jEBwUpBMn2OdgynO
kgdAB2I1qg0VcQNvhdxlDHG4gGqBnljCgHqwmUr/o0g1JgSKxe9lbpV323azn2sr
P3Tg02GQzbZaFN22MuX+9vcCnbU5s87oWFGnVfJJElc2ksPG5ANdzj0yzGWLXvcH
AztJu01G8Fbx13cWr9E4PB5na29Gk1fg/vSsDz1m7GMRcxi5cHAouob9TGADtwQy
GzjQoF3X6tJ0ZTOUJv+p6xj/MOtbGSTwSrrjOsilT14pKg7Yv92HiywEiSLBL2tQ
MV23JTCc9aT8kQ1qsbPdC7OtZ9UhmwShT9pxlyVwSuPsOzl/GkL7O4Zcw/SfiVwO
73rg43sH47oh7S64r4Rob4qvcHILpDO8+ITldYiYSpTy2m4azz20lmma6VzEoeSE
lehAZt3KK5FqugOP5WfPwePjGZu6K6dGgA+2A1X8qLlUZWxCjusP/j79rlOYKD4W
Uj03XLBy32q71g8YIAeZhaZ7PNHx2FJG8UX0YxweyOQSZlq8b+N1il1zXHicODk2
34Eut7GKWSbZ6i8FFnqG6xUDazzgPBkUPGJS5A38F36yjA6aFzZ0egzsqEsa5V8F
UMn09dnXWwahnpW7EDSMXElyHrykNEZ2/qHjhhJGmq0mdxXOFRzZsH9F6myAPBCb
9hBS805V4f3W2kQrenaOAeA1PWfFw028ymyEsndlG56XYKnOeXo5XzkZEeTCc+WT
JnsDfDsmOwso7i96kTQopQ1kMOvkito/MYg6UXzRQLDAt8T4Gt7ssybINwX0F3Mj
psbNMxSufZDBBVkr0WR0XuU8ubKw7AOb2eLBBu67ViZ94jvPoovB3pD1/+S+3bHr
2MVswDA9MslFbNqlbSMz3qf6iv7NPU/B33tx9BFibvGqXfEw4RAesdt0higJvvde
8w8psg5qJPSo+BgHLGPXdjLwNoJZPmp6uBEOcfLubbgdCaIhcdv47LKo3vErf6B6
isRm4d/J+yOM5oJgDPmYNFhl2vC+gGyz2lg9Sbq0+DSbWVa1VgPo4yxkTxvtD2rC
A96ddt2gs/GdacX+Ef22PQOEriVA90wIfcBHvBthLGSTmmjtg8vDZGut4/lCt8S6
7Lmg5l6WR1V0YGb/VjOZpEYydPOhB47kZVU1hqhb05g=
`protect END_PROTECTED
