`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F0a7soBY1P/1jukGs+S3ZfIMB+zLYTBmq8kX7gRlWVgamQRminWTNM9cd+VrOJPl
qNQhWymSOr9Gtg9rmrTrp9SghmCYxsgkHFHwHpY3rlXlwXus9CVzCXpkYgC41wY6
ygd92enSfLj83CBhkIIYpfL7HM/lZpXu0TIFvWeDeTVk0kYZ8poaQpI9sQm3Jq2w
Y4BOpR4C3/zgK1Phcz3XC0zL8w1zz0lUZ62xz8OxT2KtQMhdAVK2b/ubOt4XpSqu
Kputgb7P1ARFk2ZlEKIAKUT2g9f1j0tlO2OZ+wsMnz+av0hTg4VBRdfbbQgREjOd
TkE36Zn4Jq/+aAkwMx7okNyeSCGkh9rt/UQohQ15ks0XQH6gSp/1NCuzB8fF3pSq
hiLsibcOd4x1mp7TaPii+g==
`protect END_PROTECTED
