`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1M5rTxsXEoKqmellBPkQOIwe/sPeHC4In3UfIH17ztSIO7VM3p2MOoyHzSsu/JWl
883oblzGZRi5qoEt60TAy1EtsXki2VcY2RG2qbzANvTGk0sonGw62pjnfSvyyHaH
KtprNASJCt/3zVx+lfEhCoSUDURIf3UY0ZZjGw6xhxbguWt1rlRommRlwRjoD5By
WyxuogQT7fWId79smBt7sHSYK/05ZltJ622sfuHmsnTZLsnYf9tX5Yh4KfNVC9F1
SIGmbxrE7neR4TjbOUhRniF5Uk7HPK9E1ewWmb89utGE4/kRvC7eS+qUe/pTE6ly
Ff0zN5TWnDzqX/RO6bAhG0aDIlvOpYoJAqb2zeSSia3o3/bSw8Oa75jC/tormhWC
55CSyWTvYJw2Fjx45E4hliPMu+m3oww/CTKOBB8b5Dt64tS5+BLCZ+NOV5Q0XZgu
J8lqwpkpkihdsSB6Oj3ANk8HrR3iHqR+9e+MbKt7JXelLeH+kOVcdyWfF7Mi+0+f
Idb+7+stUCpMteM5eNY98igAYn2HUc+bnqH/uTL0oxiki+ACDacWWXei//QGhZKf
lofPRiSTM2zP6jz1srN+0bdTJo++9tge13jmhnUiOO/a8x0CEdO2ZK0lP60VUlZP
YGsEP1PJbqz6tRBCiEogRMucy/0eBQEFjVSkljpM97McVJBko5XT1qQ5X2yLjvG1
PibCYE9PIlm8Pgyn1y/ujg==
`protect END_PROTECTED
