`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a17tqg1JKOUCz9/jIAUIazYBQUrS1ZWmUocGikqTkDwDExmqNz8FvE41aCuN1wOV
9fxPu6ifuA+Ka8A3LdCB1V1J8bcH5e6kW5YEiHDqDvvp8lkTIH1dqjlMp+RUkh9W
hrg5j+zOHwtQULfOfdtV0s9JQ7PdqIZ/vshvWiX/p77dzXRhEn5b580DbhMZjPFl
XrLlfIuVHDZMKBW3TFUzlrpgDQKKpkP85sGnI/tgDDy9WGW3XzEy/QxA9lH3Ki5w
xnizd/cTf7eoXnG8ZpEpn0nk5Srx7Stb8tWG6RFgxbiuG+yn2AGWbz4mFHJVZlvB
`protect END_PROTECTED
