`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILxkOO4Bq42EwZqskxbADOahdA0XtMB4WXmR1taLLymvAODQ5LtOtkNERV9dTWWQ
Mu+1q7N+oEgH9Hkl5RDM78na+RZkoIktY1EkqLZVUc56w0vID72qUCSVtY/TPOPD
5RtbEzv6Jwnrq6UOjBV/IXY+1Itq9pKcc0amc2kQtnXnUlSeZePqZDs5JqRr7mcs
XWvRtPbrbCaCZNzM0MKA3Tz7Q8b89xWUmjGuVkQtmwLmsbdK+iesPtQe/TNBHHog
E99gAmPWaHPJVu7gGYMXE9izmAM41uBwEwocL4EqHQxtMHTIFdu7r6NTkWYEOfFT
n/pAyfdWxgIGJEFQliiMFrBj8AptVLwsJlAI/7V0JEuVSnMrmTRbuG0PGx9okVqN
ZexBts6wmuIXdvfyE4tUzvhNW7fZdtwY0aldNVp6EPGGS7wuZE3WNAarz1/YTkAa
GlbaQiSeziC+M90tDwmlXAdWTr+gID/Tq4MRx7cP5iyrKNnD5/s19DG2VgeFIQte
Xbvy1JsCU8PP9RtsOLhMDiUHz0fE+tsAIQ5HtVqFh15ReDMsDnX42ipRPPtHz+ZL
huVGkcUqBXrevXyKFAaFZ8IvgKxTw67/mwf0+yrNQ3/zcNWiMQzT8fqdg2NWD59e
qffyvdniL7mMBzXJII8iEA03NOhnI7iT6Uk/pKunIDsrBa6J6VWvKwevSITrDHwF
dhVYlLn/b/RD+CGzWqRQvhDy9bv1gCtYxG3xmHIwGoMHudxd+gsMeVL6N/qwCfv2
TMGk+76l+ilNUSbignHGXb+uLLCqmVbHGAQDTvQi8CMQUPbb9qX7Fa6JbULw/2pJ
vxr0GJ2FzZpeWOmrZgonsAvQSUeRaUrB/ySBWPMCbTRSJXNNnPUL5iD1VGKL5UD9
4BXbtae/zoyfx2zC1hlfqJH5v/GP1923AbPrNsNt8lzcHW+9lpQ/+F3CebiT8uhU
TqDzKCxN3ojkO0roRHE6MJ2gXUG5V0wc9/+0rM/cc4YY5ySxh1hA+AvxDJzY88kl
rA3tlkC5KxG9kLXS+0yRnJ3o/upKey3gegO2rRMaW+Pv5ChLyn/mLPFcEnc66m5y
YzO8klcPpVNQMxop97hj0d14xYIcIZzwVAKMfwwhucInS7PM45G2pzOo6guxRGl9
5YBhiktCi+EEkLIECev3hXrybTi5xtPETnfuLRktmCuCVtLc4tpR70Cx5KFWThex
MjQDTi7HCi0ZpXE3taF0+1KSMOqXLu2FCOogqyZdZueUS9PYwKdV1B0JxHk8A5Pn
qlOuGU5o9WHQoGVcMloL2u9nSDKtl18zOlvtXnbpy93J3vW9EXB+zW8u4rg5OZXO
ENWK73eqOy2EKD3qoj6afG1vWlcS3XOwYuglp2iGvKhDklZ7H0tMC+VbsLxpc2Rj
KYvzQHcquKJlT4zSCThxnGxIdDHgrtHAbmUv7SlFeu1S51EL71KqSVHrkxLQb1q/
avbwDKFqBw643W+20LsVYB62VKvwJ4mxxbsTW7FjTBIEM7afz0imsQXwkWhxVMis
/Q50CkiKOOnCBJxCqvQ2RMNwXxPFNaogp4UW+L8Y4Srzq9zxnKYzk3a65DlDwrS5
voWPNuPR0mf2nOikv9xgNIZH4tftgQhzs5Wrc6Ged2SJBiqmgwntUi03NQai662Y
6p2oSPDD2JR6n6/vdHhl56q8I/+HwrDF9/wQsdYPuxyUI5v4wvJvKI+dQf222zht
ftDsvIO35VgAzcX1T8RIfkkVUUDDvqyp08mQ0qC3F1rU3YzGTSUhb4UEoUU5c/kz
2NQlpLds0z4RvQmzj+EbRwPIy4/DaFUKhKKJi8CZOxgnBzpvSGIz0FJABq/pYST0
ukxnNHkO8W1nvlN9PhvBe8/oog0oj49WFM8JLq4T8uWs8MXfE0Msr0dt4NJqdi6u
bVsu69WIBmcpE+S3pem3E2V/LDHsPRA0oD5h7vSERV7jK/Apih7+BYVWXXJsjfpp
pntavnhOQlLQWfrvd7Zws5yRLVkzc81qJOrIWflGf+Jx7fDF0EHXmil1ff0Fy/4L
4yZ/JXwZE4iQMpWVO/ZqEdCxv+d2FtqFTru5i9kHQDolkocEx/IIU7bFLopBb3TD
26n8d7NgJbLiDtcMShpmFoPoEGafVGBggdasmXCnMCg=
`protect END_PROTECTED
