`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9aLgnMw9Sj1ISnbj/0Z0HgNTKjR55wW4P9N3xNKWWPw6vxXeRLp9AU00os7Xvh1m
kXptxokzBdlGtLMY2ixBw5gSV6VvaejSWwLP1AwIuSrsYhS0b+GZ4O7MMJuQhiTc
6KMTdZoENyohsGoIFbnOjNC5MG/a7nTcyj5jUcm80aEaMiAyaeHxVhVpIhBjRhVJ
OyqBiw+71LvplApys6r2pIV6C97SG4ASUrJI9kRmrtcKAgaZfaSR/Pe7AOiYnFkw
2aZwg8jkJC+iBm0m1CjYKKckDAFpS3+mRcFUTF56fGJznfWel2YtTKdnO+ImxCe/
baPy1XWkWo4LLFL4MX/zHA==
`protect END_PROTECTED
