`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSHSsWisj23Ha09xexTL3BQJVJ5SEPLHRyvfQV4hlvxF1cqCwpHUC3nqWEgvPTBD
ulXjqxMfkZEvzJwjrEzVLYop54W5xw9p3BD3U4h8QEeXnd4C0EzHATsxvXA+CQZZ
VdIejvpwOtDhDaAqklWieQFALtQ6/4Vt3sJDdJO9YEx0wLHE6Y/VqsDx46/B0N9o
B7JMJ3dibbdpFRtmbUUhGNvK476ZsLSrJDgsEFnt8dm6lq8AX8sW5JYFmKoMoG64
o8OFONAlia7UdVR5SXyZoTjEBpYS/18TaBOQ3aVnbxco6KaEm/ge6qNrS4/GP8MJ
OHGllH4eq1xrWe+xGDizs4lTXxtAgsH/U6xH+Sh0uwzJfG7JfFtpvwMkFr1APpew
RVKADnkjX5wM2Dpefx0eTvKdjvznGzZt8f4WTH+X9mkOM+HpOzeMY0IvCBLalulR
dg3CPizLSimRs2xXUoT6T0o1r/48GQhW8j8iw1ST6jiA3nNOAnQWDJBhHzxif/I1
YcwlO9WpxMQUEhPIWzTAZg2uA4e3KRRuO6Kq7NSbE52ZCncyKhyCoQkVl3t/mft2
ysEHUHduMSxbXfH8Rsz8CmJmPa+9Mw6eGqeU6R9IR6zj5oIXcB1EPoWet8cuRvN1
PM9cRIKGdGHS/315hBIsuYks4l6TWBkok8X0rpuMlim2OdG3A62R1Q8QUmE2qSCZ
yHX1VTbYF2wi0GaQAFvtvpP1NkEurXLmemYp07po6QWC6SNFAKYezBXXE0wInBjG
h2mteselKpqs64mY3uszM8z3x6aWeOYkYj2y6Xxi/WmwNA/AQ+FA/QWeiedy4eVb
XmPY6Vq+Bp952YCX9j92RdIlW9qyziY+EE7cCpvuWsZCAV2Vq4RVQtcLoP9frYlr
ezD7U9V6xY9pq4prwX68mX3V1K/FW0fRAtURh/tEXYcSb/ffQVat71CuPBq0oLhI
2EEOatURDttPtNltgwk0N6eEMQurh3iSM/L3PFsiXJKwMB435kboGplTY9Qj7/1k
FTDSY7+9GaBD+4o8fzeGgfnrRLLr959h0P1IhL6zNBndwHKvphBBMF0T4t5DjAr6
GoBCjC09u2L3HD6Oe2jrg4kVpn9VjwsoXS4MZVter3qYvANTEoUBfQQv6ZDN9UqB
eaLF8RbgkR7pVuqNfD6OrVzZzyVO/pDvLjAhk/lVxIfbrSoTJVkZi2HZnsTcLENc
hI0gwMnIuc1fKc4PtuArBh1PPOaE6wDXsQSPBr7cdIZL2QSvcCuCncen+DcIaBlq
LmPsNH4CuHq7cFTrrv8K2Cg/zMf1Nz6c46N80OWwWyMPcDb11E9Khurj/zGp89Kr
kzVU6amj2MhfYlOvhD0wASQ+ET1bN7xldlYX4+Tgxgdfe/yHmcPvMDjqZyjg4On5
fX4i2B2MO6vJbPE5SpOX/3v59ixH2efiqwyz14jtxexDchoWE14IIGxRqGamiMdS
Xdv6Mk/9SYD7M0iBZGTLZWktECqJIb64dTfz5zAoCskxcE0bmYnGAUc5bVkJ6vE+
ht3NybuB/TbFycS1F/o0Tm8TlBynT4NjSDOkxmV6gqaQzJWLBCuzTomd1WaEHsBr
HV1eUSO1C5s5BmMq1kBd6Lf7zW3THTYfzZ6zxqNybRiY9QOkAKcGJ/Y/uRLtOk/3
t6n3iPmJGUjY1jWdqoB32kj8RF9DcBJ1uikfbkJYG3TBNJQ55ZVloPXdajX6B9CY
W9jUmShN6bmZYYMt6juXuRL9a3j1okl++6wIIqb0zcdEPIJQyDZu9PD9rQMAR1OE
q4yTi/eKcU49bYyH8lJTbd5yg2U37kCwAJX+mNC5FrbQ5O+Vr1mB7Rpq0iVm58B5
BKUBbIpVxvm77Rj3TbN6IukuHf0LDyCVIlBdb1gezDBxPLjQ/UjcvQMFN1/mVmUm
2gGk2OMBakO09UpRZ5BgIu1QyfxhA8brF10kJFrnulE2DOfsOLrzNNPn0RuHfSfe
Kps++3CsrfGCb2LCNZWBqh5FQXRTTY4/vpsLzfasCUjExCQj9tji1GRpPiitXuwd
1zwfjCEL9kXuRyrrKsfEfv2Y7hdF7K/sQ2yTtGB8q692Tu7oVXEyD4bAhsfYlrMt
VhmvKwQ2mSAb+HQ9NFj9ownKxIexa42owfikzTFuNwh00yrgA14DLxSiCCIT+xpn
P1VIiC9Uy3Ki47gFi4XLhQCfnNZhKhCGSpucaQlYfeBb7Q6qo1ibKWrBbRX+aew2
kgi1k5TVlGe39KLipC4Ezndayo2tJPKd7/AIyqEGgZOXC6m3t7oyTWpogKwJeA+E
F6Tq69ODSheXUlMM34JiBKj9NjattVS7O5LvDY5+dX704gh9FLhmxWMMzgCoVwNC
khy1Nghpv+xDgKTGy/vGZsEFPkxUhzH6x0vKMhUWrVrrOZbiCVNlDKeIVLFq2n5q
xlqncU1K+PVp09HdwdizdOAbATLlUnjUaziojp9RCdWwvVAoZ4sgdup+w6OYws8Q
SaO0lIWou2GYzY1XyoYfzaNRQazVusXCzZcRlMaAsf3jOQrMH2UA5GWm9gG7IQ9a
44ASRI9Nocp8iok3/eleYiyqePvylWm6Nu98zdGlMCMzr+AjPeScfbUukHTI0vSz
EmXE8yldlfmkHORjBKtFLiFdo1bW6ErwTidOCxEXF5LcJrKQWE5VlYc9dJJxSDnf
eehi7d2smz4w4CHgPVLoECsJzAislilLX588sp89EAm4d5F2fcs0rfn9r1ZxiaQj
K8+adtBw/DQBo4nKQwIjLdsXo5kLRGkfuZlpxOmVhGOKt1TzetIY5GFx2d+1Xeok
z9znpEaVsLD6pH8xPje7qNbOP0wWfrkr7kiX/MZ8Obs1oJB47ynJgE6R0ZDnGrtR
ZZFyGjhefZxLYUcuPS79UkyYLbtxENiRfPJo9RnrRqwpnWCHJ2Vkfsv67RmHgs+v
Ifm2sXEG3l6CAVd9qFwnQM7ubMplS2GD2qfxaLDn/MXGikvVq2rJyPhU4F0R8GlQ
hfjwxBqjOJ+30s9naXv0NqX3FMVYvR5VUhZnVzcjXSVczcvAYDZYoaIdvrladTuc
N+JMhjFiQffD4U4sQ/7vo5GOSz85+Ed9AeRzSOmoXB1fOOd3lyZVZv1hc6SHeIIZ
7HeekdOMJvqLmVifSjO4pOsRTOYsc7cpwBWbR5QD7LmqigIaz8akphXtQUcy0b0A
PsJOhdkqOaJljmKTu9zDe/ub+rUQmYZMAOeauoKxdDJGHxxyO34GpHXoWiAnVPFJ
ZMlSRsgtcTGEdJz8iJ0THvkzGHv+klfLGh+RKS4MEcgVk8IvzMW6nCoiDxCGTNgH
wHsE5wXnPkQHCQ34YijCsB+6TXMXJxCVlV5IHd4G5k7tMO4zrRMamOzKqXTWDlGi
JY2C3/OBp/qp2iEjLvkHHfIjfJGugheU05fwIg5LnZy3v2uZipyZ6LTjzpsK3fog
0LA26e0u8D8Pm5BM8xdtDtAPLsu6CLMRgah6tGPJ9e9bGPIPL3xV9ODg+bUvFG6o
NIN626x0TSi+fK9a4Q4Tuu4JDKJByb0Q+7xfJ6oX19mk3r+v7WQvpGps35EJ0O3C
W+I4BfDVXq1eqRlh5TrV5ZjMIVd+RiAKhNge9LfYdWJWraLS4WRC6dvKcphj6LD9
Afox/dir9KOpFoyOcYaF1LbmPJaSrOUJcuvzjr44HoWcJCZK8yxqr8OZ+Z/OQw4F
vupnyuMTAYRylDw6lfClHNd9VrDAwfo3pEFikT9D5hM85B4Y478uMTiAaS7plila
IQUK44olY368HnJmKxEqx30U07MGV2aiSbJeL2YGbpmf8wQCmBZjCrwizlVljIBJ
DX3BDhgClOwVE5EszA1vc/iKCSXXmp/8Cot0z4SBhX017gX/gk6TwJ/FuAvWwsTX
4uXRRIZERZizDI0HgFydjktzTpOboSfp4VZgomR8mvCKxntDZTESTiN7/lEcXX8s
RtOyZMI/7JdzaRRRuTQEGEANgmbJERfbVoj1hXcESDFDxD2x7AQjm3AAUp5OSFEu
hcVzzRmXDnuDV87OZHrevLIRsNmGMOGfdFyCXnxx8/HnZKyPxd3i75l49d5TFir3
WWvH8y5oMIQ02tXatge+aGF9jiWViza/l1nc0ZqGGCG8MfjQqkmtei2IQvXqv1zC
Cn8hF/DHojuArOfbtfJnSGYI192pJFk3ghcKnbQMSJorfjnfNosXxD2Pf19TTt0C
lq4RZFfZm4whufMIZm9zxbfgcCS6npjXDSV6s4dzd5XMu5VUmbW2H0iqwPTHtUq3
yRHRPE1Yejp1IuPvBglzZrc3Hl1rd2BqgfUXSG5pS5hfzjmNDt7BbAiIsxtdza1n
+TlWP4TS4HlUsTFxPzX1C+qeTnYAKwg0mryiCZDefrZlPHE2BzbZSuI2F9lko2Rh
/Pau8zJQjj+egBy+qUPuvm1AFAOVooUgrIJoSHD7l0Pjba/9n8xUhJIpDYmzq28F
T+TBAru8YgBa4G9xwnHo6OEJ+7vAG2ygMOE0CmFs8riLzHUmnlTvzoFO2hmb2hTk
+UodKH/CsLe5aIz1GUX2B8rOeDkJufM5/oK8UIXRydAxd9m9Q5hVSfQc7+9I0oA8
06vtTuNiWv4SkmVccNhMkiymmBi2NTJA8wl6bFsOi9bVKnA54f6lhOGAsnLEJFUU
HThRH5WpvUGS08vBtMODmHtKy4VQC5LlZlZpEpEl+p49FtljpOgmu2U7oqkvPgUZ
Sd/e8WE+m2D9rXkbq1EZ2VCMKIy3chABKG/NqpC94jDXa+7wXpH95aDPNDClZKpS
iBc0bFAx3vugr1NaCJkXFVnpsetIWy0QP8S90uN9BHsxINCfXt3BOS6ukpchwOhG
wiEghm+JA9mrgrkCup+c+ySaFiJstEdZccaf9yaaKkR/VencQuvpBRA4KEgIYvfJ
6/WANlyIqPAoze2Z3ds/6UAnq9xXUTdW7PRajcEHcfFj3bks6NAPKRLxs4X+bdYQ
ZxFyFltUb8b3dxnTj+nYx+VUrN6SAgTQaHg4ENSqKV6GxVedUqIhz/Xwu8dHL60k
27bXkYgmhBSVfQxEyN2hSck4Ml3aJ9mF7B3OFg7W9uaShtOlHt2cUk0+vxSt2U/L
K4TG8OhDsgNd2l9gxdWdz7OdTFs/Guwn+lPVxecQ+mxaWoY3cf6Xe73qty55eoa3
1InVdxSsyST5/D1LuiVxF/TTpFcme3LEv3ezhENedo+lcqxUupBGFQGTY6QL3Oso
sZpVNQZvMAKfAPlXiS9ewam3GNAMpDBnVpmjt9ziHmyQYca+z9vs0BjcZ7hZ9NNg
fr13bn97gSHkNBfdZNsQk3nIPjRE2KAnl6bVZtyBAbHcMqkdbVt1Gn8L2sb6aRz5
SumPYEnZ7FZ7AA++uHPFp33NrsHYhqVi9GbRtniLkul6Tkn47fFawn6isw57z5C8
Q7I3kig9gMqMdxQdah+hIMerDQz+hvRamWQB17mK0+m/yN9Ep43t075ZqZ0UyFFA
z7eR9luNAnUsvTJ9wWST8UoTd/4KHXkjVQ7rgnpxpDbfnShztWgANKoXqaUAAHB4
r249DHhmnXZpRa6PtXRdYjtnsneez6TDJdT9PRu2r72nC+0qO9fLe4UZQPj3mE8l
3gcMevdWUef2oAJYRbJjr5UmyuRbjAegn4csO3XM7BODDEQs6jKJ51mL8f9s8l2j
PKgPsROnLDELRQh2iH0w6BCcl2snyf2glapfZSuDXA4zEoiBTMnnO6xSzQLcr6J4
wyjyKOTVq7AeS86cYVM7tG4ID65tZzPdzenB2DmpQmqki0PtlNMtJWzJWAiAJUyB
TD5FJ8iNJHiGKk7W1gwX5HD/RmH/0sHCfEAd6dsgG3sLsS9ezQ5JCswofdtERTNy
TXlXzMOqiICcnYp+01TgvmA/eHW195ynOzZQdaAnqYeFQMLP1BP/RQyfkIKBCnGm
gx4F6/vZCK2FYiQumQYZnOrNnevsYqEybB9PPEKQ1xKIxjKp+rLjhpwQYn8CV/3V
PTufktK3MtglzlKyC2DPXRqmuz3m0SMEqYroVCsET6Gk0wOgLHlldEWslTfK0KhF
IVO3qSGXOHdWrG49ivmaus5uHRa0jHB9RM+zzgMNoTL+/J2F5Ps1LnTzMlQ4xbKd
LTOjHwUi/qWCohclLokFEVBkN26dHJEXu3K2nyuETQlX9MYI0wlxf0pPpRJWNMva
xmQFAFTSJfOsooKWKEDOZ1t02spKTCSuNHcyJrdJEjruuJ7ipSl29KWqV2LU9lFM
kdlJp/AQd2+08uaTmcSWBGFT4jCpre+2uUCg5buQNA6iWokfytZcPaaD82JbCYMV
eZtCZviCv0d3LMyyQ7fggOjeffi2ly21MtzXaKgxXtZxSxnJPO02SSYW3ShbqHP6
MjZ+LoKDxJ4MhNBf1FeF8SQ4+rAW/eUzYXF8Wsyl7TYwodbVCe43yHL0XsTAfywe
YZQiTrWM6u/oUOAeguACrDi9zS6WdxY/VhkGQw3BPqFDyixq5vfvVNM39ipVT3oH
xFClIkGsqyemWfEoFrOrydlAxOkx/03ny3HhROzUvN/GvIZEz+AYNFPOUv1gVPD0
sbiGmq7VMRmAeHDEIk27bnyYJXD9YGiyFzXOfz/SWBeqRYEdYTqBuMWSt/hfgEjQ
LFeA8WYjJyJfQHj7cmsqmjU7SobCZbfcw4R2KA3xiig/OnqZboQcgztWOK7Ij47y
+K7qcNExG4N6xzteAd6wAStPEj8UU3Ngcx0Yv0oYanZQyL/gNulgBDqhqbnnQ8ZY
sFBe1Ds7Ph3IAASlRbe0OMeErU7PLFZCvWJvxcOSkDKpTFv1ny3SIRv90kCPz5vG
fmFFTO7n1iPpIKVolFZQJe8yCh6vERuTXiGRqXvXgZUgWxGLe/aS+vAclYwDlcwy
PHRwkHyxI+jmovkDevsBygTqTC22vJopiSXugauuak92OXqZaarHjXhjv/KR3dUm
flwnVYJcpFcmapGiimfwwMLneLdik5x9++eIlxeC3JgvZCZTnBTPXHxTYRfS+49P
DpeXd6mkOIjttWxs/WqDOMX9apoJDchSIUeg9D3DgfAbtWfRx3+7HVsjcjnffKYq
pITYBjaI5fpdS2/vPL3odIOyaVQ1i/4ctqTto14qDrYseDH/iTaX8m3N5gE/2ess
LtWGpLiqgQOaDypZO9y0oaGJUKzth7sQ0oJRjaFLMDVaVC/tycJc3QvKQXIQ5AZw
8Mu9SKXMOsDTUf4wV+UFnnHYfGtdKj7a19n5izS2aqZ6qbXMaZMrbSMlQWf2bwQT
aXo+A7fLiACG9206HWjQKAEJeZumWrVyBFASBzOp1Bpu4hEu5UW2dQizRw9RprVT
VfTma2k6+1wZmkHz8elrgcVvaCKaiNEHJ2opFB4ZTZ4K0vCfVcoTUBFy0CGJmTxr
10Bg74zN00JjTt7vOgRRv5E2B5FdykE220wmENJECrgQdY1ScFPzFHfKdYPiDMw+
9G2J0Xqwd4fV7NNyqUdxRD3IS0t0A7q1xWOIApWNRNdJ+FTO0uNRP0AOjUS8exNh
qd+xg74jEbax1r5wbYfftf+3jByvskWHNuLs6NqMPgB+h/Lxeuyl2DiNJKLM5SIH
X31gMwSGKyCbZUKuraAANunH28Z3U6WrGHzxCLMOY1E/Hy2ALDDtLmrZ16ikYdcd
Q4tSxf8JbRSQrdPYvDDvCpCuPrdzsQGcw/ek0wHkLjHHN0hLScvP4GVyieN5V0A6
LKCHQwcEPMgdTQgrkM3K2FpfNvS6HoQN1rAWooAbX/FzezgVYeLyWkPEcwS2Lnk1
krcaTQooYrXwWY4F1H4QYpsE8zemXenu8Pz6PysPor50Ia4sr/F8Lti6D7vy/uLK
FejQsv0VSjXFbTA7mj26oA0g5sMc8iB/M4uqEgB8QwZ8UM89ozMAXlCyzMJZCXqv
dv3e8W6O/Eikfcyl1jy2CVseDX+DxT58IWW9NQczbPI/k0bO7F6n2M7fQRCHBYiX
XDNr50+JxztnjzkMyUzUm2WNM2XOXFzGsq5zH/6IekIVLNH33l1SG4Ok12CQ1Xgt
qonefpiBZ7G8onkb4MibnM5Tp9S0LBGTvl9w5Y4mfCihEpqXjeMY2Q117Qpqu9br
fJvCE0eHglNYkwAIEKX1pS+VIZTx7/BviVEmstabQLlCTUnJ5s39HeiIYcFIbsHC
9PXPJSvNMnE8NErKgmux6qKMVmrwmTPBbYrPH7CS0CMGuq6D74xDiUG1/iQlroyp
/B2r34gs5ckrjp6qCuqngQkEbL3XCLwGnqR/slUs44lI0RIZnQwN4RukkODuTxYH
wEz9dvSn8HKAFpU5HZcPX2sI93qSvlJg949jpaBhGjHs/A+5361c4wCrLZ09tH35
4TWybAo/ZuVWpmEbh/TwolRbu9V9/R5UXZ2XYe0tZrryCiyOkTXyQHPuF3uWWZ1U
qzXsZnLZriAUlsIz0Y1+AayaLRJeyf7HykvFlzEDmgiXkS0EbNuP05hC9mELbxww
BW9+AEN7O+nltwmqj3Pm6rngrAadqjFFwFVlDrNz6sAmGt9vX6hSZ9ZA+RoasVTN
BNLl1wpGQAZtW9xxccxnISjDVrjtealQz1fvgC0e5dWySy3/V23zYvg+V2+uc1PG
X8zg1+0RNiouqzaK3yY+Px6ssGrZ8rMunB4qcdE+R0a7aQnDVPZOEXaH4ffG3Y7W
KO5KR+DWEm8zjq1u8eBY9bi/jtkqVAshPsJ/SzRWltTIuv6DU/WvplKgxGlNr0t5
3u6fgo/pF2ECRJdBsLHXimOZAz7Y4J76VG4TTCh4+ecX47HXbrCvKYDi8yD6U+ux
5aHD0i53F1Mem0vJ7eSaHLJT9eGfXUuzRXlSVgEo2fF8dVgqURqOd/OUAxQIxlgS
JcqpBsjTDrzb4mN/nqLUqXFyZHmGZxWBVcINmOfJ4JdHWeW7rAcnDF+RkzgbidcZ
KCFh1gjGf+7MVq28YtWIxzKEBgQXqnLRiJ8CRtSCafniyVzwBh1O0p3w+YN4RYF0
cmDC4V+U1nTE65gfmoyqmLHvotcnW+s2OLGnXEk4WGza+aTXvaRf0bXBHLe/lfBI
Pqaq7Fv9bcUZRMD8N71aWw7lMVlPE2hlA+FwCbV9qFzG8tEIhitHSFNF16ioYuZu
t2bZn3pYhDgp4QrJ5rzxe5iVZTlzF1Mr7ryPu0rofwoKtMDD+2kU6BFxgzKrro4j
o31dALnJe3OyFFeLrbhULO08ztGiL+3bXrZmoAPKXpLoEEgARPW+xDiq7D4zlSS+
WhSCNIQOXMk9ppia4zeHea+3hn5hF7c/7K02oayvKMBvXXU9feov4k/h5N9ep+8u
id5rxnQTa+NFK19eeUo4zOaHXx+vo2FfQoapTlneObJdhlGZPWgZ974f7Hbv4Py9
/aQwGrLoz8QWbDNMT+tO13jXYRAa8nTg7J7nXUFljKwdfDw7+jJD0UzqngFcsh00
0lGRQ/9I6xG6eIn3RbVSqdNYhOkh1UBauNUsTrX2ag7y0PcXkaDoraawB3ChZxNv
gJbFQr8OpY/zfOylWoyXxbhvPnt4q0DEfkkJvUFL7ycdclLyKDLOdPOdHn8PbJpX
T+6Dps+t9KGPqvFL0ToYpw7r4ZSMjJVmc/vzBK9gu6gyWpC+t7DoJhI74+xWBceJ
FUANwjsfqcO4qwhPXhBVX3NZ+b3BKEtqAjBHrfha5tHEoXo4iEHL+S6XV78iGHE4
dwaPuZX1sOMX+/zkbRB2hA/9SoXEDD3XIsu1EOjzxr4/B0tsG+HvI2XhhO+24zhz
2eva5RXOk35XsmjHbGz1ijMOzUM2tPeYwF6n+tsxt2oy2Zw1eWJOag7Ay2JcULEH
Fa9gb/mAZ/pU4cDccwf8IIjGcEf8DqLiy4xwCNlJ8fzxAH7vEYfCl19RuEnv89wr
FaOkfm53A2quZoZIyiCtyAdMJD2c1HQO6gcZppzlKmRDjssbDKgNWwe8dxJ8Xs/0
y9drrTjQA54SRAfy7dCI+VY63kpQ+bt2oUrKyOGBO7x4tmzELNN9AcBMC0KQ87Ne
D1Lvhb9F4nEuOXaa3VPGJTtY/ndt/Ph0O4yYzIjD+2jeL4mdUgDFIVwsZF08jMcN
OzO0MFYnn1wYyAdCN3B3I7cgf3asj180Zig9jAWYQ8S3zBEDuSvfjCG6LU40H3at
aMqCVwKJH0E0M1Ya4+6R5OnGrjORYmB7zuhJekiQG99K8r+ceqEntXCK4bLZM8/A
TEID+btItfpkiCDNsjtia4cBoVxB9ECPWiC1hNZwopZXNTNICcfZxLoA62r+NV34
KpmjnckbLq+hyEsEZcdkyi7rxGBn+7X19mBuHn9nNXgW94I6Yk8wM1unghxitQY4
fIE6Anbxlim+73NzyuEV2MOwB+B3b/LTp6S+95HNgx9aVPN4LjZ2jKccT5SxeEYY
QdzmiuGAy3t5uDpq6s8G0x2EBLv7yiC0rKchiIOct7WBLsNjTESP3DoVQFO2730T
UxtVSZIaWGpSsUOrGrLiWBZancq06U3Lr6Tndzha0LPzB8JVN3onA/+aL9NsyYGr
gmaKhTTRs+/Z36V2hXPeDvX821P337CTKUOiXgvd8s0vfnUVoCjFPmLm6u6Xftg1
PRlD2NBVVkwLg06kt241CWuK6MCABs+z21QNjyn/MiXGZuY2pxKRZB71tN03ALPl
Ck5Vc08TLqMvtMnzQb1FD5RY3YoRfYz92i0+auzDK2/ykMKErig6U1a1io0wChIt
llP8L19LxlIAthBz/xuwZKv7ZKrjvnQJVMAR/Wpb4D1n6Li8E9kwVukvx7qwKA5T
RhfVgxiJNnTdGgpPgAV92h623wGQZRVFHov7qmc0tPBTew97MdMS1JfowapH/gC+
mdZTaeBkul8Ph1dpP8j5Wnulppwsjvfa3Wuj7ur309T1AVy4Da0YyR81BIMIkbqn
qilx+6OiQEwb9AHda3Vc/aXbkI9o7jJNcsorTu+CuRUYbrlZWx1J3y7CbMP4KsD3
UyufBF9bTieFUGczz3M7RhW3U0GjAqtKpnpfDpNce+teFRiG9fc/Pmz7zED2WMxK
9zjM8ubeYxVFuk90uPuKuTG4pij8mN4MOfB+YGPaXsaNkbfkxBMHtUcJFG7rmhfN
YNs92i+Xr4KgRwdFs35l/fvsiBuI5HKwVwBIw/vSYHE9ngmhig7foNHR1dizSFMN
JemDoDgJcQ2viPApYsj0X1WfrqtNgTN50qKmiWGfSV+Tg45orc+HZXq0pH8s0GaV
01lVRU0gNcBLtHveEm6gvmCQ0AE2kOKDA0ImMP+GSo+uadp6fXDqAdSgPGqOZC/8
ZE3J9UGpa17OwWfONMwQewoxIrRcO+EmDsG8un40uEdCYGs7UrAQA3eZOHen462d
i7sS5nW3zM5AKxPWuJqrXZKybzeKCYHuGVRdBiNqZy4tsXnNGb1WRjllMds0cd4U
r0wNHWQlnhqIzAhug6EEBUszUGvHUQUhEbyIcVmol5ml14ySWbY1gW2wTLVBcKMz
BwQR28OEKZruBEm+p1ZSVxi2+Tvh6XOeT5amoXGmS8TBpalWUMSim7zXXlcdmtHG
jCXE4Q+S3L8e9rAl1WvNjq5mbS9e/mIxpahahs/SAMn+KcUw/9QPujOIw++mDV/3
UlgzBny83aZborLi+27UlvlBq4YHy9yDGW3wbzsS8h5CAaZ/BqLeL2KmBm059Ojp
MTvm7UiWR0Kas4zYg3y0ABkvGJaWIskC8n9tbZx0UTcl8AStG1CL3c68zopaX3an
QtY91DKNhsY1os93jigMo8R+iNDQtYxxIgbuLIKp3pXZGJxSkzelfPNuUHU4dAsL
R5JVN9ySrQaL/hMSCP12GKSc9gmd4fCeMhTl3x2Xgdy+OkAAJNljJyppECUgGVSz
QPqbHCEqmClhTfBKWie/GUdGkJsEyU/8etg9voPuE6jojxFGJIwpn5lkSUh1Sv44
/fszFDQJFozTVFH67Cn6FP1QOj95epmRpxoVcBPfM3/uzVSjeu0qlPPtehoZKxgn
R1ARgoHUNNKNJJ+jqkacdGwuyf7JHUJsVa4T7UKtN2dYJpzy3CM8DXXqu8X6DV76
T8Oxef932q65voyhi+WqJuy3lPWkoLMGtldA74r7NgE8wUVZRARo0wOvS4OIOwUj
//k4TJZ+Xec6ZjFCg9IgBmu20ax8seQnsxO1RYtjNzn9KFDl8HBHBaOPiwyzNbUU
PA0ud1SsrEEh+5gFhv6yQ5Y92M3ihR1q6yz12zz72Zb8i6PnqfnnD1yZ2xzEXtRe
sGBhP8akmGbvhh4Ls7wYing0dKDmWyPHBYw3BJ2xPXogpwUCPXUPJ7LzjSqm6B9h
/9sQEGK5/r9DhGLo/qA6xLc4Vc+TGevxBj+3Gxt6mgv2HTD5p0XpxehXHHxbUwbH
5tbHfWwn3uj3a0bco/4oblNV8WRoZlL8YMm7PbTyXqvSSahz0Sq9Y0oBExxq06+8
gMKhG5Yt4enn6C4J9VvvJqt7YLlUTmw732x9tsaL9oYRsPQve/SyF8ZhQjiE/u4W
u05TSAybmvsoojIJzTILg6ySGgaAR5wvgdBLVXvbS5nvL1iucqi4NrNvtIy/mcnW
vUp/tpnvJbpASo6A4aTKUohHfeYLQhbnwC+Lb9y0Xnlm116BjtYjiDd65umu/tc8
GeF/1xkjV8QkBdvue3pFqmJofupS7mqUsHxXIKL7BNSLziA0mWBB0Ueah2IA2MRI
ngZpSbJgnid7HhDBpKvCduRleM4Vd233IWQpkiblA6Yj5CHECD/fUyK2HYY5FJuE
62Vl/yBb8PD3WrEZUi6rQ4wRK8IXmyiUNiSzxoKtOw0oORDK121xqEXnG/cTP395
2y2kVCCdAzn+H/Bor9nQP7TkPlAb1xldUcsXURVWN7bSGKGdmKczLX1wNux7jJ/f
G6DawCwIBVjMM5OPpMpNxIO/KjZBonBaFqTSzh9SBXpugl0LjSYdtIc+qbyrGG7J
fza9InDToAGAFouPmUUij51iUmLt9LsAQqszM62w/bSqTGcWQaV4foWqpl5Cyoxy
k2NO6GwaB+EqY48kuW8ANjUqiJbDeuEtNnOt2lbgnJxxr5dH8E9mJ6+qtB57IJar
XOdf5gYBStkJ1QLNwXky6bhCwlxuWZ9vFVXPD+WhOs8HVW8qTG5TKgZzlLHNhgFy
46IzhhccG1Te9+GZuNpW9MMbEC9LypKhO1cph0UXIeYEaD8hRBcmhdHEKcB264IH
/3MF/3/ph6oxCuBV5beYDiTmRelJee2DyJJx7WgpaMQk0f6L5noS/Y3opyTNdGoZ
0T4lZBTOe0b/3rEppMSLRS3dl6rUjRXmhHYnJo/LaJS3rF/DUTGYz833w+FgyjEn
srcPB5mT/hvz4wvPIbuZOAA5nxYiL49MkkSL9GeRE2yqCIosyE5WqBZECmmGF9z6
IN25jefOALsLzqVo2OQVj3Tp+ZN1vA1ZYG63PCKjO5buTLYpurvH4PvEbl5+QLLS
kkMI65/DyNn6n/POPX8fk4glGQU+MWBV/P6zqoktEBMHCFoLlTFFxm8bNqxLwuYt
H7k1LWVlvGaMUaVRQ02iUnaJb/Oo0z9X078+JgtxlJ3aT5+cgT2euBqNhXmrk7yx
ScUcrMGbgkRu3yuavIo3auf2tgPnjBiD7aXXkygOFu7xntb1lcZ93RQCIRxF6uFg
daUYq00IR2HBjPFRGkZlhR3zNydpbRefRjpWSRSRhscOHAUmfVwGzkEriLoapR+y
cLVjRdZlxoLToaC+zqmUD1j3pSs6qcAiA7TurlrTkHjdRpF2V3FbiE8zHmTAX5SS
DyZdbRJf6MjnwX/Ux94K8AqDVWI1o/LbmuK/1kfiafX8GsHT+hvTuKeZ9WYSvJGX
sdGJl3dkmY1E7u6fiV/Oswm2/SBnwPXBF0xEigCIFhfrpqrWnBne3+bAbq+WPDqV
8RdbiY+9dCKDV6UxAG5T20MX6UZcqSK76bgrKX7MOhI7xRKTK2WwxhhP5Ofyh5pC
zNMTrzx6EkTYe7joJIg4GicthpCIoqeY/vamkI6ILLKfFQU/JcMSFTfyTfpKUyaP
WKkc/wqweW4ii++JpNadqPhgXGj+52u8Erc1RJxhbS5JGFMoaJjM1dDC7E/y5jLJ
Yz4JtGdmQe1RQ4VclTFFXPNNUFQqJvePqt1t8AzLmrAYOWXRiWSiQsDP53Mw3R9b
bnk0E420nf88MJXz5N1uyM49cR+XIk1kgnzugiEnOZ667zKrugJHiZ+XIBqWXX5A
GwkbA5FT3E5MeORUQLSxleKVS6zGQPTX+yamh1AoVoTsk8UgCWLF19CTKeXNORWW
6d9Q07WS0zcykD7SEL/gec913PqF0ZyNpCkxN4MXsCpYRvTTjLZi7PaGvQTdn0ae
SfcKvkGOjd0N1wyd+6L2E72oS3KXMs5bZ6wUh29VXxDaq4YfhXE3VXvRsvCoYESW
8IKrPOdpsl26jl4lLQ+dX3Sipu5NdYdEy5vPxaJoeJ1bUvlf8q9yKiwSzIsX9ZWK
mbkMZ/rBfzBnJvd9lexAIrhFERb4JgeISdPJvDMTFDyNGgMiOVEVbaG+cRbVxrCw
kS9sJCrfvujU8orpbj98vetXEH6DS5eVPiJHVPp+RgO+ENw95mFOWnpI2twiuvBG
tsDDtjnwRQfrhAf2b3ga0sGepeGWSUUiyHwYLUXsIQk0NMGzNJSryqMzCWkkKJh0
7e6m5Gni1ASbMalTdRfT7dNEjId+e6offTU8xSeAeJfFpZb6FCLpmyjA/ULVbzp1
ieGeJJQDE4rVtsG3/v7SBLkRfcgfpC5d3Q8kzAl7Ty+pAL6EvkG15SMohAXVjP1y
M3oNJWNusFTNl16Lyas0pHBO5ePJ0IydmTYwYk9GK0AB80wfav8Vr2DjVOhyzRV2
0AJZLYzKsceWYKuZnABMfwMdDg1acrcFKASWoT6dMQL1dgjWJc89nbrc/IeV/O9E
E3to8C/YLNAmWV76ei/rt16ikeyW7poB/RfiIuT1QV9GuDRernk1MBCh8c6Qw2JW
giiSQQ7ZxF0fC9uG3PaoR9ZhkTHJfff1HTnyc5TJ34rnADkH8SgPvG84EU7/+w1+
1/4J/cTn3IOdZ8Mm46U85i3g/RZjg8n+4YYNivGbVPIrCpLmTm86y7F3tr+YtBwF
8wf+2q0dHrsRH6jE53nHqubLtrbegzVKVHMr4ng4KeIxW8/HQ13N2tTfxCLioPb9
3HBSkgI+TCE+r6lEQDmgV5FB0QzWGTxiJw1mjfEYbbJR5WqViUfs88qzhaRXl4pv
dRVylAsY4oU3H3KBCFuDJRfvJ6kfI0oklCGkXrGIDT3gaB5OTnXRsxeb2gnQazP+
Csuns8xNQxSRcwXdJ/U9I0VAvkW1sGEliqAo1f47V2nUlW0M6ZsQA56VGeY+WZbC
oezyUJ5XwfHs6JZmU5ZQTuyuCCkEFpQyCwkp97vZE/PTPWobEjfgfEvHaJnqu4to
8VpuMCXbJ4d5EkpSnDjPMlyRyXGEOiGb1yJm99V5/NITarIZSAJm0iP7k6u5FmKD
vDZl44I2mzvYWehBYVkHAzXuI/41gPKX5VpdYi01zpAy1SUwXhziuArFp5hKpEDQ
kRNTI/S52fNx6C7PPkheOqki8lST/vAz6sqxY9JRuD1Cs+8a9zt/fRGRnNf0syvu
7LrpWHJZeYJ4eHP7cleXzIGqKJBvQ5lh1YXWeFyupjSWS9WXfTQD0cvfQJNrHbg4
eqMBXQhNTgtajAe00vqyLqEbFjPdTie4C4NhB0EQX45PoQmdOn7zW/xa66WJIXtL
km0yVngGU+ALALq/MJzYTCtP5k/SPYEdQB4i8UWkd1wxDJXCCNGffNcJcGHKibsH
QLu8kqqAIkxp0Nc0uvbqRP+s7/jNzGsNaMkVHmiFssIzueZ63ATsSbwo53qThgup
WkBVRzUxygH56BeJrldB4JslZUi2xQ74uqlBZUxc5Hvx0m+tBSb7e6zaxGLZnCqa
knS2Hvd4R3sKGvDo3TWLOn0ZAdLcIyWAHYDxb4cTmLIdz428Pp0L12oFRWt/yqKr
Y0ZbvW3aeFk5uElIhF1Hi1RK5gcXNJdw6SM4PYhFf2VyFkrH7X+Yid26cZ1iDl/3
+AdTBwLabte1fG3Kc6uYg64U/ViGcL0TqbQrfDA1xX2f/OOF066qmdQln+6O2U3e
jAtn46umhrNjLmabBelwZYZw8WITKcILjQUiD1Vh6NZUX1P52jtq/e5FOxq9afKc
YN2YbC/2CtP9DWGRBK//hRQ7Iq/rPnakmesiJ3L6nqnVTYWavKI3NTeKp1OtYhps
MlCq8A8QHwq0dj+LdWGUczabJnVANUxsgPydSFkpanS16y+fqy9vfuy+ieKHM0+o
ziWBmFepMImPOT9Ydj7JmjlCSoEA7z4WK4fZRtegg6kzTwD8Fej2rQzuAiMRE5jc
xru2Mm77JEdyynFLiR+XMxjNMw46Z2uvDWCX1tkZPCoDyjXAn1BbwTs6owWGrrCW
aP0IRQ5kYka9AL87c0vUkLj5LqYNwjAEPnULQmIYvE0txHO71qh3QCCoc/rk7oQn
SEkdsaQCkgzvthk9S8otE3sWWk6uRAS3W3mlw1npRb8n2S74HPOrF9OCKmkO6GoA
e0mowxxSfj+CKTRQn0ZBaGve+4Smatx30uWdlhWWVWPayQvuZIORN871iSN1Cp/g
frJxfba6Vg8Yqqq7UERNG5fUOd2f6BzaZCQL2kHh9O0yrXWqVCSMIm1IRxjHN31E
GGN7wLhf7We7bBCD1tQ6llLBqSt6XB3eQLhT707Cbw3fu8omMy/r2Ztujo5BlejR
uTbZcDNi5R8Ga0veCYWXL1fxE2XtRls3RPBHTi0eutUnVuO37LIMDBh56zO4gJIg
mdbWZCcmMh6RGw2JB2Tf4AMZDrqcexDuTbqgdcgVUxcikklCumgJ5TIvWScgIxjd
LfJfyWu4SzU/P596lrjqN+vi3PuR7uCSOZAacqnADWkOaRUHQ+Tt0RADGqd6gmxW
KIjMUyJUtmGTS57oaPLdN7/iattjM5+pcqF50QInBjc+qH+60LxkLYKGc550Eajh
Va4uYcs4KBt9y3YGZyHodGF7LgPVf3efuudyWDAv6dk6TOCa9VHWRrWk9DjHyhMy
qFyFzjwa3DEZSUA6Ug4/0QJsyQ66mnCvaFcVXabWj8u2L+gcMz2aM44Q00oDFhtA
5i6quErjqPWGFQq+egM3eIh96lKdaW9BDEAWovKdmX3CL5SEmBrcpBx8tL4RZHlG
alezxWYxo3KaxqHs7nEoab/Ou2aerBWSTSXjRnkXkzdCrFXD60dUroUF7FoRjxSf
x2HUwA4YSHeI96r1PUani3Q0UZgyRiSSciESiBTIaky+K0tzsIq3f8F63tqocHiF
eANp8xiMy8N5q31Uo0r2r8kPPNA8PVamLdCtm1EPt71RGxLVQYdVxGTV7KxzetVH
rQZ7JZ+6c1sPQmk4p4RN5L+qkXTnHRI15gY8w/dB3mCVoWQPI78l8gl4xLoaftz0
CCHZxaDspNNCjJbPA16/64wugLmemJQE3xonCHOIaUjcr97HAyXRjnbRHxU2IZTc
d1eFpOYlEsnNq+YQ2W/RxTmqHPzx2CYIfMmG9MFKbQMHNLjNjR/BBSTlDgzRJgVG
/lz0/eSJPwsX/0Vjr1ovVYJ+z65hoFr6Yi7Z2ZiKDa6x1+pf9fSOI5Z0yiJcS4YV
vBlOJG7TP+bC1TYDLI5Zt5PrCDcZznUI/F4YctVRZ3PBEeBL4m3sUBjFtgSEvE48
rWj0IGHHyp81WNEJP+Mq6I+RvePdgObz+GXOz7/2Vyra+PYpCQWx86O9hcjQgw/7
gSphmDx4GjazUaLsHnr8yJ+C6FH6UrlNtpO6weCEqJRBvHZTNMNoIgiTea+tTOFZ
R5bXcHpZK0mPMVF/UbIy2xGkXKY5T2XcNqKiFBVbjtwu7wEa6MqWHFwGlN4dutiV
H8V3NBeuvRI+LB1wakDhLI/So/qgwZFCOEL5pJyrhRehjMQc0IYLLLacqS16WA2P
h4529XrKxSDXBy8QhkB+kp/lZgTJaMhst7Xc0AC2Lpa0Ujqdefxe+NDQfZ3VOZsb
sPRPMZ9Bk0Re5M+2WrOmIHkvpXjPYYpu5ejQyt1WvDzarwd84caNJJ9RvGBmfBPM
B78nt9Jcun6dEpvlZPDGm8tm48x8kxWSQbN7o+/i2RKe2s7nrQwF3w7uUx+gOwib
rm3G4SLQKYsI1AHnMp5+BQGw9+w2I3j+7AAUrqbMrsaVQHh27qiQzaBiULAJxAyu
EU5309IDQ+woGIB2ej8OKuc4WrN0gv9CDwuNHN5mvCyCthAPz/yAlEwiRCPMbR+v
m4NYsVrpgfVxntG+tm6jEMOHzJAe7vJ4Vm55Rg3oCkTB9ci8lIJgTpEvgOmPqDYx
Gz8CebItF/RDZpFbEiN0jycaGJByM7Od0We7eG9tRxryV2YMx9CCUqgxEs9jctws
goPVsypU2DCRA2WQibwjSA2jpmYY2Hh25Yvk2C7jm9bHviUjoSkyS69h/MotZQlb
Qd5eyldSDTxSkOql+uEpOSbUdN5gS59ZPs12hv5uKqNGBvh0F2M611FA7FMJhgb8
/g8f2K0DudMa9cjgLADJHwjBKn0IEnO3XaoJByn+NNuTmjzR6O+L0OAuKI7+WlQl
UXdorSuZW55zdod11F1dYtykflT/5Qo/sw3amEHV5+N1sv7EZvPZhRPxubahoy9N
GoDpREGMvLyLI0vXsrAgBh4/+NwHgXI3vgNIBRFWIJDaQt6dlUZgUfjNOB2U9vKa
+Qfd+GPBCDnOe6+trH5eC118tB43j75lmzAFUWQX9kss9vz4ro36zj4PGJ3Dzi+k
9FO7NHqjGa/fJ2Ze+s8w6YH/ykKtZRSHZ6WmQBWAdWmZeUJqJq9KfzdxIt/JQZ8f
95Tz4DSPk5WjgHO9xxzo6C317NBsxVbR6YSAeDz0UfHxm6FJ7QVSlRNbVnNyEQ9E
AfzcuADVRGOCH0qtTCvoPvZtLnUPvSFBhV3fMZ4hU7UkoiBmpCvNup9ikZSxyziy
g62LyWVqix2Zb+xDa23mMvOv+A8RYWemLnE5wLCOyf65r/XTB9rqOXFIFznLIpFc
hG9Z5IRC+ZuE6U+042mjCB7KA277yltbvmDMTr3UM7VjZEWgvR5jmGyKHqClLwug
Uw8Alkbfn5rspUUWzGeR4vbYP42qvfHppCXpOSYHwR6LwKdD3SX925ye15hiqL9R
g+WChRjd+FQzxRvwa7W3ME3pYMgb9GNhv1vLweTdAjJvTvw8fkWBDDIgG/vvQMY9
s6Rmvq09ozhk4lr98Y3uGOkffho1ZjrARQVjTqovCLJcqdP/9htBRTqaU2yX6W3A
LjjWdTICABHuTvjk9/TrytsFqIErjZWqr/8nDfpsrWbNrRNVpEaK15ZeXEVxTWQC
fXLmP837JK7K7xp/hS3tQjCwZOpNrWgIVHR3uw2d4XVfHC3kj8X6zqhzDd4XViqo
Mx/6MO2dqCfdX7z0VtBQQjYCwXIU8bZJt/IohQkje73MAFijnhCVZzNgSeZJpZ7B
ONLmczGamAxcF4+B/9KVAstvM48HbWd7ag3aZs40yzhJgTVWBJc4qA3hR+61S0fc
vhrcDJ+0KsumSYIxnHn/c0mWMUb6lcdS3Fm+uVX1tZwo/xcaRxHtYqYwGjWXh9+V
zxFTTKUyqTjVWPIt4QvxxmCklw1A7U5alCp+Ni7GxEepLsUAZQ2lQTxIhBmqGfkf
/Gt0amgTmqA++6N3YXJx0pMNbvTTM8v9iY+A0qVOmaw/xkCD91jK+Y1Y1Q+vGfdA
JABCXkYEufHaHeGswD/SM3SK5SXBhDoPKiu+16UsrfSQ3ss7R83RTc871CLSMzee
3QWY4kZ1lF6nyFrv9eO8ByLiaguOsFER+DM+cOM3ZjQjOxvIO/kRWc2wftoQ+Hs3
GSVrbJJSG+PSXs+b0MoobPQUiAKfaDSyyhhqmK8aus/Nle/UxE9y2ApQcGEKmeOC
mRTJLXcqU9v9VhvanRtOBjPsXnhMKjj1oEt/6F9RxEP9VwIRlAHU4NYvVOf8qZG+
zysQ6mkp5CZlSYnPhlW5bnRLiY4KWp5qUXLy2c62RvBxLnTyUDJ9WGBWHvYCg95W
xDN2S+Z6O8frWsETn2DmBsAJxPHUBtH26+VqUqIQSX7w974onJv0+811lPn93gwi
lkSd7dXajRxkAvbVfr3rzxGeINQkP3vrmQe5z0Z22Yr4Aaq9nsrIrXWk3NkibfMf
DX7674H4KzMN8/IFM/GFbvQR8xnkLhDNom0O+Qp0NAywdwqbjy16pA5975E7JCre
FD6DDjVkbxTUBxZ2aF2zC+XO8+xxsO9YDkLJFZPtQuroUla6Q2knz8094T6F4F4K
YXr55VdcbOIG+uwocw5RLYWPOnpyNmBc66G+85Z3wOvudzXukKkQF0yx14pVuHzS
+LWl/9hQfOa3OqS7iHFJyKtuAftZ+05L6eigwYWDSqf17BQpemCkjlIQhmVJhhnC
ijNGmVI7Ur6BMIAJvbWlHv4P0ObmsISDZq3St8xaYWO4ziwzZdyp9vqK2ilaJ/cW
wxfzydME/wW0XFYkfML13m0daWj5pRsVojSt04dDVXaCrcRtryh+okRAhBGsMq6j
G470rmeLypif2UBXxPwLOLhs/OP7KDwKXmBFT0aVlorwp+VRO/CnLug3YSXegYiN
bLgUAlHN+Sel6uTpliKbrzhvp6BslWqnFHaeX1p5HLbLF4UQQnEkMACgeJYhGUCy
tuGYYFDC7V6Ldg6yUHhiOlAQxJ3uRrGq70w2tQe/YixYXZ8sesM6Hm8gIMfnWeBi
wbxOciLRCX4WWKsrG0Um8HB5+YIR8TtWWH1NLHBr5tESqdvM2GyqrrzeV2MDIgf3
N04ZVSHUDUKNXUnIQe3zaUxPZa5MCgwNSXr++QxC96EGfTM2YM11NloMLKqq0dqp
KcZIi0YXrgWAiRZgkz0kgGd+1SzSnp0NYPIwCKgeyqWaPrAHTVk4l27tWQjPjAMc
H1iujUAIalA8JM7W4s5gemKsbqgVZwLVF72JjFj22iUWBMOd18FUr13M+tturNbS
tuEG2VHoBUYdVW6tG3zB9OjsbX8CPNhuZcf196KI7YYhClL2TFDUlBZxojnjf83s
IGdD0In66e8fL0PeqaIDyNHr7Eajh6DJlm+hjtS9KubVr+mgjg8wq/XQSiTnfVxR
hTYGrtHqPYLWzpe/sZVCYRhYpMT7Z6HA2hGc+SFAIRnvbRJLEllAdrawI9skzH6K
GFv2+H9Vt5RUsboXKTszPug6godJzxDoXlUWcsnUdmjXroU+4BraXK+Jevccx5DK
mMKblpRkIEAB9+1IXP0r61252DwjTmucdj1cnQiG1ltcHb276gD1vpdzMV2mBOzs
0j5aPgVnWYHmrwSm7fAr5Wp6om2O+BkxiGsQ3lph09XAsq/wvo9GlaBLa2WCvr5B
JlrGazJ9jHXieFHXj6Bdv0tvhjmVnCNKmzWy78q89f9E9XNN1/fLqi8/R5wDitvE
+DeG30ty/8MKwJonVDG0hXEBsSBgUk1qanRwGLTAskWJi2phAB32UyqI/FXBUmMK
o7sx+oSC4bdR/Y19zk5kD5dh6cKcRHQGnrI3CtRYKLdpOx4/bD9Tnw8ZQlHftWi9
siPWfBYdm6j6gs7OMllM3wKk9uYXhTgW9LqFO0WyDXQ0aZtjKxQu1Oatuj3g57/8
5BfR+zUYnum4V0GXBx81NVohTknbB5CVAZsxNg8QyYRCIhmEVmHV0ViET0Y5dOMm
Uccvxn3bhGcD6Vk4IPM7Dm1WWDu1FDcFg3fUUc0r89htiZOtAKJqFf3VxmwTBsKE
1kQa4biWAe9smDvv70akw6hVBx8cwYcUQe3c9OQPbRG8mrhIsxo0ct/mmjBmwl0f
8JTvMdiHPn5V3BNfHCICE+hb4ZjKpnc+XSABaRG2qqlkAnSNSfRA2AE5REdO88FL
BtPDQhlw8kigFdm8kY+M+Xo80tQjaCKEV8eOKLnwGi8n2YBeAdMbQ+N41UntmEzE
V0rL/Wu8U4XBXfutQUnZDu0c5pQM1HQrYHd3M80dArbd0etgsqUmWXlzKtA6BtG8
2E9dDliXQ8tY75I5JmhQL0ex3gbtG9WkxMahEVzVG4HVQr3YEmGvNzR2M7KowIsi
F6ZfyA41Ex8vR5HAT3NaRFYXZ68An7cAGo2mZFYw5pvrxVTXHEacbYotPHtArLvu
VdbRJBeBIgHnUny/OcYca6EhCgQatXqUp2i/JFvmXCI5c5R7rsuSEZTL7Hbkb+NU
9uqmjvhMChE2e4Ua2uiL6Ywrc096JjMZunYIa8Do5Qv6GY1hAmltMg5yvYMjmvPX
WLFyxkrdlnu6zZ93zDaYfs2U6a6mvtidOgR9csHMZmBNSrDH7eQbyZ1OGsYFEfJa
POmqUxIdR1QVH+nU1hL/XljySnn6m/MvJyW4q75bqMVg9wlKWtMF6JhznAWEXLER
vgv9tzNvt2ueUpdmaNrqCfDFVi8WxcSLC4HnD1KJrQPZIUp6XAik56RjF4s1s0T7
OaTQ+AuYXSilLLNlpZsy142uwWaLZqCA16bnmcAX6mautweuRGWA9j6gpD/SALVL
GFtE0Py/7ahBQcmJFn4XQybLmJC35Zev7RfDaPwJQOG64rWLmC7mbqYPm2/MSYUp
z5vRCt+yremThGmgOumwveCWCpyKiUFZIyKFbu57a9mlY5ZD8/qKUAWqp/oHcuvr
ie2oQAedy/bW8T1HQpnW/K7k7VC0ViSQCq1fDnK/2DmHTFIGnnPP6J7I1v+6alSz
Tiv/artiwvx0ocPG1h0cPPK0rEOWIleEBAQlIVitEqh0JXV7QgOxkrlV38Hh9A67
iFjSK/wt/GAPDkIkqPj2R8TAJOnRoJGZ9h4ebkaQeORF5hFTpJeeUjJpxaN8zXb9
5i/JT6G2YJaQK9HV3A4pYow+HMty9u7+Ef1T3eEnm0gBhTVBI4JGTfDVdEpeANXv
z3Bmzg21w938llkQ40q1t/3iLXcYm/zVrUv2hcMJ2vA0IUY2/Uz+jiP0NWEf5rM2
+3bxNWzHTMVxY12CSQvwkRPsD8lZ0wBz9VqAUPODBKH4Po2c36yme8J4OlcNv32t
T2Bi+tbbNE0tU8U1kyZU0gVcegsIF4yP7/D/9evwOltZ66aA5Bs9KaN8Wa0w7Rck
g1Zwhkjx3i6xhw6/BSTD9neIHufcEI55F1OzAzrQ4ruqX0x2lDuifTelErMaqWCM
oaEPcIYWsJVRfOFKuPQ3ZdGO7If94xHf3gxArLQMk/JRfC2SwWzL28kaMW8aZUDc
75SkB/QjPqobvoyfXnDcbu4NiO1uhojeqjtk9eKoR0KavInveS6SCz5pVnXdpBuA
kv09BotZ2unD6Y3snFUToYgzPkwXOP17HMM9ZuIjdkKmTka+3s052XIuh+5lU0V0
fyEy+ZGdQVxljWka4lKu6qfoHRuso13ph0kLzs43x4a9iqSaOp32mDYV5XFL0Em+
SWmVN+1wTPaxNpt06b5jGOlBiiCGd5f0Caw3vE0Bl1+MiW7pNvp4NOwP2Gz3LZ96
HTnzDozUlOaZHloXGJUjKNgXmBxLtntwGlZArbDdgM1tO5qeBeDx3rGCV0aZXQUU
TlKYM4YzIN7ww5bwkywzGhKhyXTOrn/mT2PvuDG1MAJv46uDYVnoXNb5oazujnkS
vZyWW9DSzrZX5wpCS6pofTLmmITeQk7KLEPStAkDbIQrESg2hpKnbwxLkamF3BcO
yRKpZE3gLS9uKRVor5krGXw3Dj54uumxq4eb/0LQegsnrNT/7QAKevGY8++yB7sw
Wdzlt1PDTnaa6DO1FfBPanAseyMLahHGmnFyIpcsgV+EszBDl8wQBylnjYtiAVeC
vetYaojruZN2ySA9TMLM3XHIU0MvbTa/eS+r8Rxlvp8dnPJ7vHuXZiYFk+hJWrGd
6EsAuhijV6eTXnjQuQcxJnIfuBfIg8QnknBJWhAxqj1nbgjYJvRUeSzcc11zgz6b
CiIFMBoFO7HIPDZ2tSc9Wvk7uUgm+Tf9ST62ZFp0C0SLbotDmUH/FrSR1BhSw0CI
XA30h9kWrIp411IXJz2lakZlwG6oj6d58lnKk2zcIpvIDrWj4NkNaSDJHqmTGrG1
iJpHhezC6FnofYApuj68D0/QTMCJboiYwOj6eAf0gFDHtJllkKFZI1fsdrzMqZhZ
f7mpwXN4QG05SXMJ9xJwhV8IP01Cbt9T7ogEW64Dt36iOMIBDs1gx5mhrCqPjkhK
LFjjQXwo5hIlDmlQO5XAcCcWZGeTAhnx63jvQDGwHoCSNd8ZrowIBMJK8fnMDI8T
5PPWm9GSGEscx5tNN8BiNPWpv0cNqBfDj9MMyVNasvMGtN3oHljkQyjQeKs/3EF9
PfMICGnFg0GFz3rks/YEyvYU1PGdZbX/tokiAkDV2/LR6hUbQMAVQSWEZVnrPt1p
qslVRExU3E67NAWF/pSlUwKO/8XjU+XPTNHtPhQSlz31RfrrZnxXE9QgpnIPlokX
OkPhF5lBxIKI3Wx8bS5Iu7b1UI9yX1MrZrn29zs58qCWTYOiY29gc4S9Mwai6DGl
d57oDKoHzmEZ2aFTJrK5hDEsua6NZ7pdknqlV5gmHtOs35l7cnT7poOaMomnB+pr
Oo+JjWa7Q8hbdy2dLErlsY1dSsRek9zQqXbowthublm7ApQGpw4sjMCIAiyG197X
5Mei/idJalt/WEWYkMhBOFt3ZU92Kkhm+1pTcDOLnF/9wHQumPaK7Fy9g6/BRcny
aBCebfI0E8fPLvcPqb2/18EeTmd11QxGnXPnzbN2Y+81KeL03D8w4R/Zs13jKKX0
j+TLqvRrsX5rCl2WIc0UzLIM7P6vMlGiO2nI5fmJnlMKJJntVbU9MhIqNofbhsn/
pPtq3z4GEuOimdb+dNTtrH3lvy/Sx7SHs4hh97ZgkexIhAAbpGgKHs6dH+vQcmBV
nX2Igp+U3nFRBkjsFHphtBVGGsQTvDptko0jHeRqOEBdbTk0A786uJpMWC0+j1ma
oqLqSPTJTauTgR93DA+ctlFZpz5p/6gRkqzYWiqumQQoWaX16+BoX0lr7kmGWZu6
HIRTgQNhkRV7zq10k0XMsi3WlU2hO/wIGHDvw4eN3bCUy7vAjim6kKLC8FCmCgML
GkK9k2K9b9gMgsBziP24Ndj4cDf1QYtfqA66nCG6GQUPUx0BxsIOo0B7ZJOcdcJM
m7LTJx/TSAyyUzjOzo0QTOwsxTqT99s4YRu6UeoPCLmAF89KAPWKMBhTUMmpqZ4L
4k84l5qUuwoXLdnZzbZ9NaY0WEFHTCwiZFkuBlE/XdEQVyWMTBIxVZY2asbK1Jt0
IN3thHPklkqfLvn3DR4+bhY15JBVRg6znMO3QDuGlT5cyJAUvs2rzDAUxTo9Q/9i
8MUNNubFJADlTJzMaupOtBpyNppGGX/Hkczcqz9vaCmq2uMCf/3VRNUYWaw5mwmx
CVZn4Vnm9eHgaC15lqRZkeOti580Yo6KYyDZUjfsjLeCEyKNwg+YrJ0Fi/B7GfAn
X+t/VjU/7Jy5B0IQ8yrn3FzRvr5zhJUOakpOKbIU8MHAgEggTO9A07syT/69OWZR
sYcc2Y2FzoaSNg6TaNOGNDSRDrzhte53HUncZK9IbpJKbFSDb9HSWwdxML4Ovp9c
8zjRbxrjfG+X4ag93k/wgiV5/s1tImFVsCK0qWYOL+/8wS79q3kem1RS5+btO7aa
dGPnVWg2tWECth4iOOfhwksEmqd5qmzwRY5WIMS+/b2rHnIrU55W7H0uzgB0v4ex
yxB0LQcAaTqh0QqVkOZ7x5Kw6a31Zyau6xNqRxGyjvE+VdD4aDs4zK/whM9nBDx1
iFBzk5kufugH77D+qULzyOn5ZgkbPfuCywLZ15TnjNjJus+xbgezCOgbZkiDOQgO
h1DQmw+xf3fsUAF9h409DnJnr9cAMe8FterJ4iGLaNWAhtqkuurTXc/XpaSNG9Wf
AXFyxguREGqsiwFKcwRoGO/cK6egSesQrVDe0/Qxzifq4dS08PrWpESmnucTivMZ
aDgbShIoRhl2KpxT1VDwBP/nXBe+r6OrQA3fHlo/0xL103bGwvm1Zw9dDYTo9AWu
dnGci/dNfCOYYSF83GHDziOUjJhPfK2Z1PtxKvQwtHeV92+oHQRFkVd7+yFCS/gd
UxVylYhuJ7ZhNkZU3eHmgYqg/+CTJFVvGfpZ5L/MfGhB8jHkj31oIlNbZnsVhuWe
Y3Vr3SP+5f/qnCKCuJ4X8KZbLPAQwyKGlFVc0pOyW2b0P2uAYu7+wvXq9h7bkjTJ
m50vi9cGrMyO2ML8p5ASzph6D/KENuJpwu1ichQQagmFkcNPC5Qe3Zz10RTmI5Xw
YoQS7UsFVL2gY4gWSJtC4iZVSSsga463GEC4D6XN8O5uFeKuxSF8slcpL7b4VLbz
yWUlGqDRQcirxBv0TSvprLrXKMPcfjhGcDfr3C8Vdtv6wgbuzrZ1cxWbj7yeQfiP
ucIJDF4d07nwMAfCNXRvXlMlQrNyb/KAUZFZQpCMbVQI651Ap7eGJh/Dhz/ebPOv
IRG/wrCdCMfIL8gNLug4S7BqTZVGfNqhSRpdyr5MsIXi2gndm6cvBDCYfyMywFyF
+OJzQDOV1hh8q4qNR4h3pVEIPqzM5Zi9AhGBtHEm0CNho10IS80TMO+hQGaNBkjU
vjbQv/HtbbTVrqdLsTNpfKdE70B9lEvZaGh0Y1a8zseHDtvHctvKPJNW9CrydAN+
IJp6TJ6psXbklOTygP62KShGI12Bftir9IlzOb22dMaow2wNxWMeHeQ0a7TdfEFW
0uenJfAX6rTd45UkL23U8WXcM9UE5+Mz0YcXXR4sHxTqE7oDK3DMfbFBxTm8CzLv
rtsBFEbn+gQ4oS9lT4+NS2IsDd7KzH9+ejoTj1TrU0NDWdu7mh/3lb44DAY3j2df
M6olKBrdIuAeC8GbbH9l+AIezt+5ZHR8C+ET3xn7T1iHRAlLH9YIsTSdKFY+b8C0
4frolI0xT8m4AJdGl50m826kTT5P14mN4U9t7wqTw6zy2kEfktw0S3O2gkG0sNO1
fyiL4Y6TrhGYwUGAcuF+oD201XQek+LyUnjx59nQXpzUPEWyFJyrf0PK4Bzp/swZ
cs1S0wsM7YFnPOMp3Fj8+binI4wSczPDtstDWIJrBTtQwg2OTn5R/8iKQM86dSdj
3T7nZ547XAsV5WVOuripevV0bd++SxSqSxlYwLXry+KFdHBtdFptxx/dHkpo/7YZ
Q3qb/CKrxVR1nGQ7v1R8oHE9eC39RD0VfeheMMM7fHOrhXzPPbSJTtqGrn+I+k0C
0XNheZMj9H8046Enpwqs76D/5AC8CyiChnzcE2Z7gKoh3qy8mG3hxAuqFnfPaubU
eAN8nflOcOJ07pezOa3ejGOUOzPKqz6VLsNmRkxSv5FMcW1WKsPa3tTOyiVHlaEi
wyvsLwKUpiFKfJNtYMlmVDMbU/1cmDnwwh/qCDUFvNBW0rwrGvvjSp9KcJmEkhJ8
jTqc3ShLDaWLoK+yr6QCAvK2Y0Q1G1Ndrz0KZNrc/Tiya8X4j2/ATKy3Uv4sboJp
4cgx9I4Van8vc78vXE+Iof+Xqo3kmXEb3q7voYMLenYslTJAOa7Pt6kd194mLxOS
E0e6U2NiXqWUcSyM1lm5Ax3Q5pBh2AEUVp1DbMr6xPs5DdS/+tLOs32pzjFTvfAN
LHDthZQ52LijWkh0Jv1RsQsrAX51M0ze7CMqCGlcdHhQipTT0rQtxOy+1QPGJFsp
td2uowvAIh9lcxix9mRYUBfAlVgVXoTqgFYi88DF/JD3YgbSL9dV9vH02lAwrENK
qUC9x7Mt0irt5a4BsHm9tllFmWD5ZUB1plRnpq+k/S2SVOgKWT94/Mzu4zG4x5TM
5J0SMpdIjU1QjgsfPZW90Ts0ZXgAnXghd8tU1GxYq3Hp0UZjpW3tH+rlYMD+TWjD
C1c3oUcx30Fl6NEgCNB8Of1d6gKsY5AMMSWuPs3FKDq+JnRsATKfC3RuxDARsbqR
uHu1xEwOy94XjlbCq/rsdRa13wOMoptGzmRSsGP2TJZb//+989LhvXeNwL1MPcE8
oU93uMN13XYza13uhjdDzKNo5aAGSRgDY7E+q4ot+0bayU4dFg0TjsQIyOEDqi08
N/3CMbdD/+LlxSoJwm5tonldSqaNydxArsuayFBwTP7c5iw2XwBheRnok0i52GLk
olCmqvFu3GsXHluW9tF2N9GGbKeb5QSxg9HRXSzTlOsmVH31UAswFNvT4kjq+PGq
I89ZTmINlhCIMyriJ/qwQTQHn58yafD1+PMxOULTNquVypkJvj0pf7PcMPZiCiGk
pklU4TJW/y+B5/B6PZt7upDGausN2HyCN+xMdBDBi4E5n7/7OYZd/JT5c5fIOtDS
Q7OutYt5MDZKnogaTLkSF0ppvGxFTOlJrylTWmFrm/7DoOnNpOkbYn02+lUxKK1n
`protect END_PROTECTED
