`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRWeHEh+tC+wxtX/xMGkk/DoAM/Yry+rxQ2qOCTBvzl/EFaH0NzOu3D1aAkvTggK
9kIce75r9XVe5quU8AaXuARMv/MI4VJeMDdqxIL5gJmAHNTtADPiIn0jGScGpmEU
PxWhn8f4NxcpojvMZicvEoveLEldOcUjIcbe5hIuZrHazhDJQAYQQ3jNpmHoLTJN
BxAnME8C8iKFBy/bm9L0Gd6nFqzq5zZU/bFDxnzqF1Zq9dO78nqliYpQv0SID3GX
I2//j2aA6GjDA/FDor8jXeeE2IDiaCygkpa4VzSF/t+pSKa3U/AYl5uoK8qhNhYM
WEyoSavZd2YuV3NefCKaFQ==
`protect END_PROTECTED
