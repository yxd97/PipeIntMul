`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7TScUF9Uuqg9KmWZ9G5Erlu5ZgBT0OH8QTBiCTCnXodUhNxUZO7Uj5FngmGPm/ko
ar+er37rGgE/b7DUtM9fgfzfhEl4gy43pSG5SM9hS1Alk6QGGSjkkVKTiYF3AwZH
s0Y79fZQiYiM0Ap5Y/A/PEYuS/8lAzu6SVi+zMCPLg8Bz2dTWTLJLcq0YPTMdYSR
TeQmLfAxR6QaxOOlUJpwJoYb1OV3LHu1c0uTB5Hn2PxH9JRsji7fwq4AiOyEfJbb
gOrhOEnM1KWwVE1/aiko3k83cro0hJBwWUUJR9PAjwRNge1uIFvn597CZYjmsnMc
oNEY2U/x+FXaJ+bf622fXe4WaT5gSGTWSAWt4bOaqX1xTgf+6fXQbjjWWHaCZTmm
q23BWFyqY+RNO1nDK6ZhvemwQY/L7KLnUXejrolgEk/jFVUJgM4WkNkFx8+2BStW
cCezaprs2PeLwh+cwMPCXxDcMmHpjy49TW4l3gGrBi22irAv8ADfj5q5qeUTezT3
YNTo+uOeCcC4W1NHazuCKT3lEtIzsDov8y2sL8tQ72EpkiRY3a+r/IMHhEf1Va9D
zb3hucU2M1bNNzgrM5b62h7YVhMEnueWwCXP0lvLQ/6MEY7fKVRjszQsIlRsiDNL
o3JzEPEI970EKnMO4O9yr8DwLLIQ9e+nXlIJY9YWe4j67T5EiXwseCpU3e34nG+8
KLpyuTLuBWOFeAZBQOC5ylA6o1AiUIhb18nXvDlqsCeqNR8EJ3Eo9kNcRE8WSyuW
2yhvefEGx71CJul/pxazHEeKpfnnCwZc9Nx0xVYEPLEIarPn++pgsI1qSi7FNJMX
U8xOE8xzeLITMrGiNbI2lJIFhUWiLpB/Z6D6KBncvaknknrgJMESUwe2PBkEUnLs
krRHySg7SjriDiILOTrrZ4T+bFWx0wfwCIkbK/2WJoO8OZHrjI3iIiaaBQ5a4/f4
+GUA3PwTrYnrC/0TC5EMsDu0/EayW68drNAoFEoj56E=
`protect END_PROTECTED
