`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMF5Kree5kr4LnAtvvGO5eWW7GjW9nuVJNqz6YeAnlWtO7A1g/TYzQ9WL2wMYWBn
Q0FOtqY2eAvN77Vp+rGFAzDs40QEDsf6aAoMfuVWrSv5S4PYsK4Ck+yEoElbcr8m
nzc3GOATjWZqaISRRFAax6A+eSYAJBif08jjP3C6OE07MxPSaPM0PTEG8HIhKGDP
r02A10DY9yjYyD+NCxMn0nwRcpTzzUZFG6279w5b01GRfKbMJWz4l3cJNwKO/Y6z
eu2cBr4MtuaHz5GkASKOAXjQfxWKEZmK001aHIVcF+4Z5R8Ix+mmtTl6Ieg1E4vi
UUAx53kXy5H0qBt0v3YTNnCQWJqhH7fk8FmmJFQHazgrXECXHPaYvBKnmhJsjmxd
/Y7geMn1NIxRL8u+jT7i2cG4wCdJNLZtm0OjF+HV3mnvZtsRaL7VSZda2iSxTD09
JyavAh4okiIM1ByrPe4fRjhKmnO8YdJiSMwYRJ6rPA3lLYiWc7Zk1Sjws2VUrR1i
eB6AbUfjkMn9vHvxIYcFw+AVFJtxzm5rfkCI8k/2ug+RYltwhXtrDflvW3VPngPN
D5ASHVw+CEWNreszbjBWXA==
`protect END_PROTECTED
