`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DQ+xLAkRHZdY7G5NLrFWO+Eg40gZPy25quC6TpZwQTNJ1bLf3sCaYCdvL8uJN7j7
SAZAxvOsBKafaniXdCkrkDhF3RddfPxmsgoc0yUl+cwQ41/U/mgiVFyZuGhKq3cH
Rv8Or1VUG14NZVRWf6M/yHHASeIWTnJVBdH/drYWSKJ4ZGMOXRgWRd8pIfgfiyoi
V7IaPWGyOBtCp+ua2BKoVYdCtR3o3sCiLUJIPQcTL6gds6Xu1BPDpgPvi+LCTIwG
IAt4B6GcetgnkUUnZ0xblRGsw02hF5omWfgii6yxRqx7WtJ2kH1mT+qSajc4z8om
QgBtQ21POv3Rq/zAmALYOJAL2WUaoxV2zjdI1oyZ0jE5FpN7jIiPSg+aA/JcOHnE
l9zn5b/uZwmr00qOXuoFDXfBaBK2Mw+4XA6mYU2zD8c=
`protect END_PROTECTED
