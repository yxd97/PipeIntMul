`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zOi82rvXZFfBPEI1fj59ZVuIihqCKbM43BTHnzjY+by3vpg72Gt5ZdQ9QWkRIng
SFiYlfUGX8buKQuXSaMh9sNoad5RHRAANBRyCl4BgZ5H5F8X9BJxCwuqGSUtHLNY
K7WYG0tQc/doUWow6eDGUJzqx7YLs7ahdHdyQjXjIXIXAMCTrFNcxsN8PgFd8N/I
MB5z+wVAM5c1AWo68XGEaBr7TR5qm5EyrLp8KYILCbmzFoxttpOUTVoG1qoufM7s
wdidBUR4vKUr+9KolH9j136D2hxKirGTICuAi+L6fWso472GVkSeuTS0JLbWAeTT
0pQShgpl0ySrfS5V5VIuU/7Dh7fhs5KJ+sVwlNjX3lOhhsoPd9hoVhc69HS4dcm6
lpF7sS6EFd8Zsl9CkWBOzogqHxx7kr951GHAX8fObmuT+JLLqSzalEVKErI2lhMo
zXuL6zv8WStsxr/nVc4JDcyh4eRk4ytzNST5jgjIKh+3BfLfq7dRRWSd2093/nN1
dtc6bM/RIuVZHDtQoGu+ZRoZXE/+DmQ4igI5LY9ntzpJPsW9TUAhzphFiIuK+mMf
vQhVp3Dmqr2m5PkGKNOTM/1Y3LPM0aPhcGbbuej0CpQ=
`protect END_PROTECTED
