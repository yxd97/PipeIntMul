`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMg0pmsuhQ9l0YtRkEZ7l/DbsLO+eoCsjmkSV6HPHOkm4blx9VSpCrIGwA9HHzjx
HbISa/OS3MbunYA2SjpSpW53DcBrmD9N9qne3axSeO5vSfDtediaNQFo0xRb8CXJ
LwbTQqtkL0fYwOYIE6RwaXQABrd5o5tpA38fKi5KaAFsbh7QTSAzZW/P21tDxPaR
kJDnjrlPDKbYPvUO05+EJWlN/jJNuieEpdH+Qddvov7iqMquygfo5jWnxGFBHkB/
FE2TCFxtK5c0qlpo4OwbKpNdD+i/YzUEOZAZEi8/Bexzf+ca2LqHOSUpa49rwRtm
B1f6INq4C5FpzbXQ5biINK/uWiD3TQbwyfwqmZGRX5UJha0dZUSPQOXtvIBSM8da
6vFKgTSFdrYNtNa/XgcW7+5DAIrcai83ueKL2oI+dqbkg/iy6FsN6uFNxkqh8SDZ
KygeKblLUGiOEX0cEWZReQ==
`protect END_PROTECTED
