`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5iiKuWxC5D41N8lHZvDCMHcuB9Yu7PfWuNLmNzboOH1iZnnV6UGjXYmnQkWqd+k
hSKbIHcD/Y1NZLPg8kAmpFFUyuqaO2zZ0mcYBkayW4QYVWPvVBWCsEdyj6BPbK+Q
UrMqGyAwXOZRYE9b4Ed/1zNfoxrltVgJYBc/uru5NOVvwWMQogDBOtKLL/nd7OvC
1a53WtMW5HQot9WY9od6fOvd9EnrOm1NDKWOOQVi8v1b+aIAAUFrCHNfouiojEfm
YP3bOUbuh+MxTps5RqaQBL3Nrpn3C3/zoQ7zx/u1gx6HKOGr6rv1DJOai81If54A
+ObtrPpJ8/51xVM7ttXvLA==
`protect END_PROTECTED
