`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xsM7Oluzqe/Dge/h39SB/eZFtToBP46rxcyBIEnS0JyP6mn73NyjORIvlbR+frQS
ykDkkO/2e9ORDIKlSVZGNDlX2kG3JBCKxJlEfIfWF7QiueN0ym7lRenbXqjzNA3e
noSDlsj/IyzsKd0XOLF1V5mCS6yfDDCJ1hL4uG0U1NDOnRxCiFIJbvODI/mMNMRt
KwJuLjvpej4L/+lr2VSLgMYNamJMDHiC8yX3at6dBcK8RO0lcqHz+ebEwIfH0pN8
00kL9dc72JP0z3/VcWecdnGwNM2fZmOOMEf0Q409hJcOIOUiB6dtCoRXVUoLszjM
oPXnq4wlS0aB8L5hL21WUBSPhwBlq062zpmMd9zCghw+rFJYWmBWrvOfmGbXXI/n
VtVwsYywTgduXBO/ZAVeD1qYoSnxzCMD4kVUDe8TPMQ3bDeWxwf5AaP8G+LCnqiR
ZQd92tUQLRs7lh0rusziUWccWiZvLpfX/f4FoypMoL8ybQFw+6o79umqneTfiMOX
YoH6/VEJ60urPAz/jjmBw2Im5Ub88LwFSebB/gXldbzCqCeYT4g1JNQehbAWpleD
hIrTypc2kGQPSvmmCHom5tFD5Ai3kn4vGnnmJ1QkI5Fnm0wLUDndeL6htqmWaIAU
YR+Z8aYEWBMJEqn0SWbsqULZkZh2z2DmiCe5VAUl15KaNj5h3CDcUbL4Qfqc5BHy
cWP3OqX4vbYsV1XA6wSxXYJu2C6YCZw1d4Mpb1aOG3cAMthkAXPPoliVC3POWbwz
rco/CiHYSRmoNMbUZEtcSobEr7hRZ1l+vubqrwytxzx6K0p0QkfbSfF/R1l+1kEo
WPE9YGtjy+adzXiipuL/QUeCldCWHuxvGy7cAirlLpcQFRAgQ75LNaSV3+/UtQG9
vEt+FOwdQyt5gWEE7S/4hsLMzSLhWa8sfKLr71oJ/FfQBMsJw/7m3QjEuTikv4Du
caX7sewz8NF0bt60dbXu0aY64UHHMe3IEqjGG2pGqhR4t13bCVPJ9zC8CT4DgEuJ
1pMuUb35kNqrySoGGx7F8GlSYvhl5HlDswfCevutH9nNm8zavyhVRmjrPNdh+XyO
Jd8vUCyRxlH5kVRZc5BDNuMemSrcEutXq6wwbP24k9y3Jv34/+QaUKp9HsxUEd6N
9N1WcLyJVs+f9Uxi78XI4PvwqiG6u8IofzxbxikGPvq9MLcaj1fcEVjOHpqvvIx4
wXodOLtSF2FC+O20NLT+03RZFTQjdebN94UR1bBXLP7QOKI2ggVmOmAH5r/ot8lT
iRBALgMTNURysGfIcJr/3IgQJ4eA5vvA6ZPAePxF6eoyxiqZa0mA3/8K86ysolUJ
U6P8aq+SK/iHWYQQ97XmzMClbIirinT9aVKHeMM1r1EQxnfisOZJ+FWAWUhnOCV3
qEsV8SiMqQPAdkqzy7h7NCKXuQ4WEA8gVKNK5sg4zSUEIcBPsVBsfMpx7Ll/Cqo7
zmxRjaIc04Pto90Jn7AAkqZjE4XlWv4tObwovWjdUJm6Rq+R0IrvH2vuzpCund4n
kGtXFqns95L0qahZh/tG8ibMLHfNP1vAkYwp5rJTRNZnUkFs+NbSUn2voDGHfhHP
pZSzuFitnm2a7avxrhEuUjuqafPNzUNaOzsmHyw/Yoh7urHCt4jkmBzrTxsGx9Q5
9bJcSv+dhE0JJtbJ8mhg5l9DQxkmYY8AUlVHUmhy7QV0lk5lyWb6q87RZIWqHOqF
D903RjsU9y4O5lUuETJ7UCROkqNmErVt+3hFtkxsRIpGqv4GCRayCl9wT29tV5Mw
NBKQVVvcSTwD/NXdABQiQdobPSi6NFQJgDVMrd9VuO+DEfxh6dTtcCsDycbpv3Pc
ovQg4lVOFdqgx1NEtvdKo1/2Af4TBXDqYLvdqgdrIEzUX5l2QgRfsts8O4mVgukc
pQ/jz8lTIMKxL2uEwl30INVQrrGTbLP6ONvA3aMhnC4fJ34XbetM+z8G1msV19TA
Wuwp10FR6CM4rudt1vhDdckVI/19iGQZURx5VZKdi2JT8gCFy4oJhCPPjeJgtrUU
83OydxMOsBtN5vTuhZlGvetcEJ3DyO12H2UC7MUxlAN2bIxgtsc4Notx45LRAiqZ
XwKMSIDsnTDtCYHU/cfST1bXQaP9OKc2Ex6hmkASOE4aizVXa41gH7+Zr5Vmh9n/
WJCo+NHleEiLqXht6eEhaa7w6o0sm8He+uA/FKgWqlADYfNOOAj5xp+PKmvkvvTz
phUT5VNKPKulVfA/rdExpUuHvKgVp+LNjq5vwZSrLQphHoTAkCA7eA2+Hb8327vR
e905QpzbdRPDol4PS6a1z4TxMBi9ua3B5+1j3BFL+nLTNHjzGq34c4B2Gsohxxj8
j1qqYqAxDkzJs5yh9uSVwqXOanf+JxgHBP+NgurJr9mE4bJpHcLLLo+M/8nweuTi
15ONBw7WhxacDZEh4wL+i2/xDC7ZscDdmDU01PJeTKEnxg6IuxB3c1ZBGcBc9C7q
C5p8FvL8/1hkNtl3g0vowsdKkw4ow7ZskzL5rgpZplgHxXRwCfykW8qQHyH+8Tiz
0xN1ww2znHAPMuV4BUZYSBPZHMEOOaSiShHJ9E1sd0jVwuLV7P3twpBAafPK1N95
lwBpCKdYAriHps3Lxl2cQTX0dIXKy9RfvLeFtVLxiVD2JzvyeYkApjm0LRqgeCop
gt1njspVlEyzVVPUoOOHC2T219q3PRswlMba7mkLKCvEpzUssx44fjwC9/EarFEO
x0CSsSNULK7LFq9CaCT5JDpLOx8QukC3w3G/OTUDMfEYZr6HSlcvzdFW+WK1LjBI
aqrLoy13BsX0SVLiAh650mhfHvjHB02tsPuEba1DL4foVxwkVyQtpi5zkok2QevT
1hTMb+2Pdsbipzk9z7AQfuQ6cMzl/qdzOMHWIKQg1Pfj+40Gpz+2n15NdvINlX6U
TKll3/8AQ8XspIkYdx1eaUiXLlEvKS8NpCF6x8QaJpW2GhKMtX56VKpGnJ8MFA45
9gpzg/GvvVFZyhnY/APcGtqAxAENtRY+VAPFoy9kXsH9C0FRr+/7/TvNwnT+HpPk
/ObF4+nA7rT2kYxjc+kJVZX6QAa1MaPvkkmIq1OA2eqhd1gU3gGwyfNZ3DJek1wh
MjuFJRBlS6RwoaLIaZrQkefo40p87Dsjb6txI04H4BFdHR2DYezKncAOGQQwHvYE
6cc1lKLL+2N3VPPlNZ+HnhYAVPc3i5L1DRcHsG0WmVvBgZjjbmSie6gMzpEDywvU
cCKmYI0TyduIbLTBDJJVtlQR0BZL50Rec+dc44xO8AITVJRvCULqmTN7d3F+IUT+
027fKyeoYeqzcPCWfJa/dmcxPeytc/FoP8jjkgE0UT0U9pqRqT13TchmdXp2+J5s
2MmLQT2PcHrrl3RnWVvZl+RbK1m3Wz4KU5qe1eCI+MyY43H0UDrMiPj6XIGSa0RI
3O0d65Z6WKbz3v948z3jF/HudIiBVjK1VBeFtYM/Eqk6MewIeqaWKHXa79xNHANc
L3eSt9h9f8y4Ygfwi1v4uT0y6JIiDaNVJ8EiaxGhrKYLOkEMLB8Bbqd75DUhH/0Z
+XI/dXZ+D6zWrNR24+wnZhaWkwwK+zaP+QHpcyKXTluXFlGGPIBuh3kaB70mdXg2
MzYPvQMs+oViQeOdYbPjkVfB6YN1G3sCA2L/UppwmF59HCHq1k6TW1OeuELf2hot
Yx4oI2ou/7plXzrshycUDk0kNA7DT9TV8T2tgyOshuHiCJvlZX5NuzcX0ji3IAjr
7RmxOuu7fDpNeeaCqKkRPsprNTIs12h3VVRXf1BSESG15f9KPTELxI+nFnzp7L/y
JEWsA2kxeF9sC1G/3gLTKyt3gibvQYEmxjQH2B4FDJNFrThU3k2npaFpINXNEQir
yt9gsKJwir5hxCMHsRNqDWRzQ9k4RH83HMBorC3J4p/xf9MJ5Nj6e9Vf+eLPy8b9
tY1xWkk7iFnskfmRHlFyB4Z1k+GD0kJKWY9tSNZxigwlK6cH4a/HVhWq/NAJBVPb
ziPJDSAZSWQerF6FFlEKzWfkqbZNjo89GrvzRExif1giselh2Z/tn6/Zrfndx4Zo
cJShYOc7ldjXLAvniPXRRdW22tJbhnJVLAKkOg7lYxsTchrMY4CBttbY8BbprHxp
0nNx1DV9MYs0eRmK7jbbZbhxORN1KcllSf9WO9hoEhvNe4jSmUMONHN9n3ftLnUu
QD0WyFRTSpmf1XvwgIAd2/mFkkBv0CDzJ6gT/R86pLAcPu2WSo6D9MOB+8kVSPgs
N60qEmt7QZycDPRtkbyCjMOg5oCWZKN+076aCS7IAGq0Zfrvc61JPxAB+UG7UTt+
fKYBEXmrQMbCUef6z5GszAalf8T2HaLtZbG38+SGLCHL2lCBF/3vlCkzaP8hY26U
OoP5NN7jFpnPVDdUwzRdKmRvQxvTcMPZ9PmJzBjBS7/aqwMjF9AclCvn9LdhJRBg
MnDK+QndGDp1K4pBVgJsMi1JTYEPHhY4RVsg+TuqVd9SNJgOZsp8qtXOaE0mBMMl
3hIHMQ/qxabrIRqmcFsugniPe8bNxLv9yGrZ3ogesAaD8Wy7petS6+isp6z7tZUm
kcNBWje7e60nq9PpOmB8hiq9mmC5349ZqmtddYc3qQzeJiQPXGq6sb8MADNpXby7
J+glVlsXxWHujwttyxstgyRbfNHI36obbpkxVn/Ft7KZ2yDFC0Dhl6AFgVUjb4WM
uYWLg0OjmIgESH6gVNKrrKAKHZ1bxLlSueYV7bq4wWq72vMFOxKvUJmwyKfsF64R
D7z5hpxiiT8k1y2ryNNE6wVtpP4o4Cd6aYjW0v3s56K09Q/ZLr5tYEU2rnhFCvWo
JJw9cr4hbXZDTkbkQ0Xl88ye9HtsO8Da9ea1xe6lZp3VMmkR2GY8LLAER+jMOLKK
+xaYK8ymmBO0tQkZiji5kJjmrLOkg7XE4aW+0Aqbb4S25CqgWPoWT9lAG42YP7k4
hdmDRyGvbbRDPgn/03i3EtfrbPBtQSfITpLhM14fN9H97OEHM/l3NlLLqHtj4JzG
ZT2AWH0cdcGTRXDPdTq8QOXNHRjjlHrO5PSFnzGuCmPBdRIoqrWlTVpv31GoUQUH
XnXIzutptHXNKAXtmyUY3AXt5Pg9CTxKhdKTLCjo0F+QiwUGcr9iOsXBhzYSTJXA
O8+eg3CSBfeX5sAtdD5U7wdB2du6H0xW9igQLTB2pccXXtA31OSShWp2CZe9aWyF
FpWYZSnon3+nKP6NZ9X9DvFujcOpMYGmtdG9ZW7Y1mjP81HCdETJsaD7MW0I5mAu
P1+WuMzHV6fIFDECB1/qyiFvXyZaSmY03HPUNf7lr6F9OC+21qK/Ux0jiAZ3Z8A+
6SzQPdiSJtla2BCxSo5pkqVdlREYVceIKprv/CcmI8eMR9MEH8btf4Gay+QvNJiv
t4OchRlu8IPCiufEuuZcD/I3cMRmsoquJYuMY1WYik5vCG7IZ04Qo+0GBMtrQubv
Wg4XVgawQT59P7MrcJFBT/val4ZaETD6l3NadjHpaFQ0cKRH8X4WLsUBbMuXcQQv
t1vVH5m9nW1w8TT4UX7SdkNCPUoVbZSXthozGIZLg3TTTtNobSfnhQCUii3j2R1X
7E8RasurI0mg6FdY4fEv2c2gcIPnA7Vpuf4w1IiztWhE5gOD2yhL4H3l8t58NKvw
Bval5WgtqKNd8FaB3cng6j1IaTVAb5dA0sfhWgcWuCTSI6gc3jGg+J5QXM/5z8n8
1U3SJPpSbUOQwsGTzdkzezu34kL1n8MHLZBw8UzZF2hGpYG1947Cz+VomfKK1YUn
9Ug6tL1niJw2lns+Qr1L17wxXOIlBigCQhbjELLgjxYtHr3uKQ0/OzjxDDm2gKc8
nOJAAuQ4o9ozojunGsShkIk1drcRQa8Cgy+1584RZrFcjosC9Q4eFZhe6nW3ehtb
yTzEvhx6z1BJBOP5o4+hkWfOQ/thEeEan21J+zhfdYJ1yozEEmPs/9ASUd64ieIm
RhNJqmBDr5jSEvp3qatQ7k+z3AFSF8pxPcmiskR5/O5RdDiw1KNLXGXzHXIf0P7l
Ra9PrfEEPJf22seZHhRrOT1JqXyGaydCdYea2ApzQSroWfuuet96iyRZ3wvslmEm
4OG+8xbVWzUphTQ+2CclZgto8XBhb9fPMR0Y8J5uOyChMCOtFbJq5QnuWCOXS8ry
nWihOyNN7buqJk4IN+r9SIvvKe8uNoQnnEaTa2GVqTxM90xnyGDuXlSplOSVPBCQ
CY5+rjnGUQMes7wIqNs6oGB79ggYEG3kpZ9D4IZ1d6dS/VVKxsutbsL1LG6DICXL
gJJxlg9nj8deDHmt1GnmA3Izq/tA56ld4si+EjrMqZLZw+ABTNADhfYJnRddYg9U
0HdaZTDYW+J/O16XcPgSHul+c8riVWrWFPWUdv/1770rT8mqks7cFeYhhlivOLZl
kYaW2fkY3ImsUDwTMqSBP5FFZdy/PsMekYhRDfpas+KU2LkzckOARYl/Wc+qGtfU
LEgJ2SQf78cyej5g00CWXEeSvcw8nAvH1SFYT6qIRBZqHHvZHx3fhKvbG9ORB/Q+
WWHN3WypIpJXlRmizm10AVUJnPy1OrdRd1vlmaNRLoxIJczCGS1sHP7zv/HXRMSk
OoqUGJzi7pE88KTfjil1QwfNOSqHZMQA2Ti0CYI+1hsX7l82Dm/KYjNYP+AK4qWp
vzL77PnyZh5gaxuhyzuPaqhw5pNFMwskdnDmSy1NTEWy1uY931InY8hI6qm9iJ0v
wGE90Ob0m20d4wl+nfGxtQFTDXTILOrYgW2LnMbPODnm9McF1hjppT2g44zkzHPF
KBm0IS6JYN359sTPf4qLh6B8pq1R8Rnu9ui4B7b9e9/wpw4ctgm09yusr+BjmsLE
bWlmrDFIYQ0Z4I3foZL0GLUyq2jV1S8NMmlpqZOa8vEHTbT5kLBCezu3jfK7PPbd
xsRGEPT9cTVyFsDt9g9HAnLT5fxiyDuDv29+/dFIbXyqeCZooGZidd2Pus2MNUJb
KsCZBeq0Enzw9nWfSsiK9Bz5Hoi2eAa+oX7Xy5G1QS0QsTe45sl0XnScY2gm11ji
MsLUxBbgyAdGVPGG3/dTxoPQoOqttrhFrIJafFqmS+ydSq8HlIEVhPHUW4FpP2Kn
TDKf+/4CqrF78AadjsbRNU8Svu3CsazlWhUWTqcoQCp2VR4zmj4kRTpESUZOBufZ
6Q8JND5seP0+brcI3Z5k/g+K1lArphJKX1Vk0NADM24E8THn/9hXuhkmIeoMkgp7
EreyQ0agxtpqJq8p1Pyw9EA9W4OZk7GFd3fiN1DsRtd3tX60AOJVbpl5HUCTyBP7
fakBNPkOG1GO3HaiWxstCJpWydZwIqlY9ZkKB/TX38c7Pj+dL48nZOhweGD2o7gx
nulQ2K2jFzapcT+PIYe4+U97ELBFOyGJSEmlevGGnQf4rt0VQzzDBvco7WJW3WHA
NxAejXXqqYuIBZV4Ga6Ry9vxbKP0yL47zMGU8bMde1CEZNEY1v/MA8rVJKfNGYx5
91ujy8rUZOOhzWfuTdm5QHEWBov+x1c3vsbGPqDNDewbzd5HEyCEgTEVmlgo3rJ6
t0uv5VJwvyD/ENt2QF+ugUSvJ46IbtsVX+efCMp62jjgPf34v3IMV2anPiaxAw5l
iQL2QNyB/M9VN5iIM6vIoHvGOfHPaE31AQ8CaCC0v3eZhe6PRISL1dyUbDWgsOaJ
Xb7WFezh/5rZHqA7paJEjL9i3Pdq2EmtHZxAwMX2fVy6ObNc6GlRX+y12L6Jj564
z3g+dFLaSy/OkiYbM05tfbny3AConXNyzsyE440EXg0Ta14WaLIpJC2rWlyb3miU
+3zqTUA3a3MrbRUB6GOJFhFrQxRFQm0dQaw0CB7L0q5ppgyeqj91wf7UqB5ctZqk
ke50ddY+DIi0N/Hq4D8V/UINszOFO5zW2i61FVgcyNOHG0e+GnhLcD/zD4OZLjAI
/AbDOWuaPL+UdznATz6MgNLr7y5WfPvcnuJD0PSjRiLAvouDD/DqhY324Bp81isX
EafNYs7u/DBrb1gudnsKPBzCPxxYulS7PfedpgAP/JsJ09X9rRb7flIF4izanhdM
6AFepDaQP0ENSoB9CrTSIrNYZCc4syT0VwEP2Y6VT4EzEZEmMKns0ySVnLq/Vl44
hy+tHX2NFw/kfHQI/gqOxGQEG0J1ntvog16i4OYScFbDgZZstekpC4xo1DbrtXeL
crVPgeRmBrjL8Imkd/Gz9YukWJWGvdyjUKZct/5BXWhMADEB2aLBUX+tsrGO/muk
w1yOnRMiFaVi3vOpjnyj9DhdDx24pEqedqOsEhvTh1NVPeSHMGqTz8cQMpU94g0Y
9chwlCyEcyOsKjdgB28/HQ5eOKzcAnxUffE7WMX2LWqtzg69GUieN6X0MQa1j1wE
ur2VAgcCABBixv8g2lJ2zzpblw91ICnEUyEvYkoLpcCs731GgRC1FgbA8BUzhgkZ
DDxua7XO8a0qeS3OwF2KVqKOiLUztfNyiqIzbVqINquxaC83/quAbWsekUnzAbfE
kh/VhXsafxKLqoXmjSIlHwrHGiQu9K4orhXgj8kCVOiHU8STq1NXvR0l2eRZpjT8
Dd6ueuEp9M8gFtOZ8uSA67Z7mwlS5Itnj1aZiNQB4Sq05RGjNGdcfW4anqRZ86nK
U0o9McBxzwXfejovTrPTVnEz5vCxlX7K8D+Lp9uB0rxucRMaoABKu1KDoeFVxBdZ
CqlR4H3I+YreXQtyBP7wc8pbmcrctg6LF+7QLkhzVggN9tufZOIsmptUBeuyjHIL
MbxIwN3BVc5b2Q7Ibt9S33EM+7ne2gXWIM6vH7Zh+KeQvhNPbEMtSA7Vdsko0H23
C6BxXN7W8Of/E6fkOwLHoOTrp6MNsFrFJsyOlwIGX+z+uES0UQD9Nf7m+hBSZ38m
XpPj6RKqara3XOgcERz9xFfTeDLPqA6DslBsMJx6x+2vQa6hysEWBCKSCWO7y/PB
Dnu31B+FKGr9xD+EgKq38tyx86hFWwFYw26G3XiENuNNl2kflixteNeC5rTK7mC7
LSn1C1qH+Yu4qUldDGa44xkYuWs1QgXFBWugVwNsMzSPft2En7ZZg1qhoEcX6GRe
7rXL+zjUetD6SN6x2EW1HGjv6IvqYCJfm6oAILQ6GYGy+OV6q87R//J/iiO/ArYP
OYkDjgr/5e4hcJqDkxFLN9/fRiW+muvQxHZFu+ApvCLqHuts2Q+iA6OB7DaKQ5FC
2+/1HgGNqCYH02G+Ktgcu00coS3Ur2aYyyLLnRK0v3fhzb/UNyUVVrbCDL4ncggY
I6i3Cf2tBDnKgnacFiLE/CAOlTMAhvW+ZFgaVeswJdw=
`protect END_PROTECTED
