`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6W7V5gpht/ZhH+vErrDoJCi7vR1Zf7/h/rF8L9bbJRnpel/+Yw8Kd7W2et2Qp4EE
GJsKA9P7lD5hczSS2eIKFVoOaDun1Yw0r5f+mEbINhP/kaH0gRlT0/35zZQGw8o/
DU2I0dHEpp0ep4I74Yaj353N271tSDWIZziUkQvCVLt6BOWnPo0DvJHdbS9d/hee
mjfGi6/yJtTwfZDdwdaT4zW5o8Yi9UVynLzUjQP8vCwnTB0iraAeWHakpRY0cwuc
7myIkpINsa/rNBVTN0R7QF0GIiZs8vh7aF5kBIYsMX+kgFpsEUolXAE6C4jMD88c
`protect END_PROTECTED
