`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FuUN9u3S0osCk2aQ/aXe7nlu+RMqv/Jlp0xLHbwUAweDucPHIO6ByqdmxH9vCw7z
wYqdK/ytCk7g/PYjre01KmkDa7epY/C6+eF5UH3FVYQp8I5o24iRZE2+Kjme70J9
2HwExP6XJCmXNpaAHkku1Hgti9Bq8eyGTLOBLih/HKCR7Im47zTIbf0bVqjpnTCa
UtvsjyuAJnsditVSOW5sYOlCiIgL7dHxA6Q/uu/DjcndvPJpQGCKQGUfy3igC0cJ
+T6jb0XZM2wbU4Hr1L2earc1dR3CBpzfWHbrNC0ybOCA27sdxKCWThVmLVQEVCoM
ULPnp3khnCy5K0Hr8HtLavVn9Ex03qmMOd6bs6ZHxh/Vjoai0l3UR+eKfkHYZlfA
+ZzvH+r1jw5RzI8nh+TtGA+m9EVFicD97IpztyV9SaQONIHESZniAYvDLpIKBvvx
`protect END_PROTECTED
