`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mT6KyUQ8hDNpTkOfT2mksjLUdpMQOuvh1EEy+Qmf3Hyqg8V0zl6d46qOc9a3BwJr
SlRcUUlpNL6J6ViOGQPU/ivjAxvVG40JcwWan+jDweHtIAROoW3Ra+pzRaSNm2Ot
5kn6NOfDJT4kSylK20sTYiJlfNHir43+Z+3JyfjnyW1vq1suFTwygTmqQGHhI8pj
bFwFJR5wJtl8T8PM0mEYMQAUqGhz1yBcz98dUx0w8VAID9GLg5Rn+zABzdA/LiAS
MjcEXU/WiZi017/x8BaDMinG7sv8ozXrjZyeKsT2E/+IymZlxFI5SanrShBY9tlg
wpGNK6qfyQWGXW7vWiLZ9b9MhA9fTfdL/YL3+jW9lbz6MFMVCAiqIyUdzgAXIrpO
urhNN0BX/AU4Ik+e4/E9plcBY0is50iPrxQ2C2Nu/E4O1U99daUgMLugW1iITIjI
`protect END_PROTECTED
