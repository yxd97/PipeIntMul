`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C82agirQHAZkGMovG9AZd6fpu8cIJDiy5llIeB1xg//YzCktBqNUH5Oop0Kakq/3
LQJ34+J+IiPsFO6psBkTpJm6SxWRNinP7uIHhTaV2uVX9plixK+WPw3l5MkgGOJ1
NF1FKp3abbFHGfipjQIt4S3zBSdAVzQ+ePw7FY+hBvx3qHkq/Km3mRmKWAxgYrzU
fobChwR3QM4CDygPKuRl0gby6AuvtexvqdWJf2MOE5i9yuKmxRPW13q9qQwszsJe
oAQ5bberJSlw/SVDm474hKDhPPu7Ly+P9QyJoAv8lBqCxI+VPB85uNThw9ukTiXa
9D2xbIuudEwsSgvQdP8Icg==
`protect END_PROTECTED
