`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQdA4Hz0Fg0rprbd0aIyYO3EL3iMCvrPSHJlBGk5gHbsOSLrzH8TE7WiCO1hS8d9
4CqTp5vXciI5K0SZP5zypgrQvgvlTAQvp/L9nvCqJvBXYpwA892qLJRViZNUUeOG
lDBiJYriateL8mc6BPTAlgnilt/43Cr5h9fJUEGjAUZiHPkbDY4YImov0ME6BOul
9WdJ9bMe+oNj0yq2vcTlwpD485ZGDCTMhug4jKIj7qnFeGnmfvOnKxO2A0dIS9v0
NICSl+6xrLbfD5p/rm5SeP4xf2JFDmGaLmEC7CulQiE=
`protect END_PROTECTED
