`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tOQDvcEjh/ct2qurcUpCq4X1zDJrUwiQzo7UI2TPet1c41nzIL2iHh47h8dYY3R
RNo6n7djkpblhcdvhbHtpuCTnbGDGpRLLAFRSiYFPHLVqeBsP9A9AMMxoqP9pIBB
36yoVKC8WuSbWPFBppywAuAsSYEvvSbaymm8FO7YWwe3sFhlqIJnuZOgRHtkIvji
TPYC5ce08NBW0O09r+iA9jLZOr+6bCm7stID+k2HVGbjuR5IPAt9GglQnY1BdDMq
qIdrCl3HslprY5vlKO/kNg==
`protect END_PROTECTED
