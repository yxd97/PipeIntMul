`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPXEoRwapMYP4/7MbdxHC8UTi8/5s5cFJAYBZTaRTYjntYv14iZtVdXS2HM+95k8
vHiAGAKAcOwent+mnHN2zsMHcKNQ/mNznJBj9CVqqP0Do29VN9tBeAWpaYypSCyj
9K2MNoWuH6m3z5RHeqB+36KybpcbfE3yipKQ5J24VC1wiffSs49j1o5WB/iyric0
cA7aNHsnfJVfavIicP+7YU80cHcjpFx53iyhYBoFEMXSO0jp5ez+9MykNkZ0R/SL
5IVckVCAq2IRQkFRa6JKiIs95t6w24VQoQgRuN/77XKn2UL01i6UDrAOboDhTg1O
AdNvV7ahuAmf1UF37FKm51aZ0gygPbJhDHHCVFGB7LbUk7VDUMhfHifytSLE26QW
UOgJEBfg343rMMspYOY5v/vl5OtUZK9UU6lndQZ6XqJQV7jxdyMbHA29s9bSytxO
Om90LBpsJ4ljcv0250boIPRZpMITMuO7XAiHSaI1zpj4xa/XFVqU7mYs/3qm7A9i
StRzLf84AJb4NObzk5YZ++nh0XMCEouE1+e/XQtn+kM8wME+NwAUhWU9B8cLhf9O
6e9KV0vBzWzpaMCGUtnGTrEZrak8BK2gwSvmU+5j7mPO7TYGOtYZCYCM36Km2Ign
NOG6Rv5Yq5+APmVFGk7kQMH47fRQ7CyXnVsj94lNRw7wEHx2gHmzoe7F6S4IbzUh
A82SEPn3uDv53JGnw2Qteg==
`protect END_PROTECTED
