`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkG0wUwThLeGuPV+PdnvZS9NdcNZCEp2yjOV2QjdI/WpWzONnkWDtJt0qDKn/Fwn
XxbIGGzJyezJsNNwnGFJOaAciAtohssukUCETYAOwl35085uem6eoAK07Zk1+etK
OQ7tWH0tdUtFh4D+8wDUxmd2OtNGoh7CZeIZ5Bz+WKhgxm/joOpTanOl5nvA+z1M
2qa/JPfCkLXYTFdxdCM2Y0aDO0HO2TCI5XeNHqLZZcwElhL3RMvllEpzAj0Sk9LB
5gG3gdXY0GFJ0kv7frNcF8KamxLsqGH7u2OSBI96ZIqilnxOFAI/7iz0UpGd5Dmk
nnxREvpK84WkkWj6VaZ7tA==
`protect END_PROTECTED
