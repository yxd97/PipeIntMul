`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1oTqK84JzTA4C1ArCO78pjZ4VpJ8NdsGambJAncJtbAWmPrsR4GVPwYNcsoLgvAc
ApAn3/YiBpZttSO3tRRAXeLiob3pUqor4eHxTpB2BHXJmNNSZ1HwAhZYzW/akYOO
VHX+2OVMg8/2lENBdMZPWTkYg6oMjoco11dvBi/lGWFa9r/qbhp9yqjklxPaxafE
B63+KUhOv+H5Y2p9JKVmdPcgle1KTWl+LrltODS5cvaILEc4zDQyeGh4tCUr8XRl
zuyupCRt1i6eSnFBh2+7IsfaiaLY2pX+gH2m53OR5NFBj3EFTX7pPY1u61azQ9Cw
7zxwJBcN6JdxOI/FzCsUTp6NCNWqUE9oZyOTTz1+jvZFpjHzeWobj540vN3Oj6st
oqa8yO4Y3lTqlp89SHy4mhzXDvpACZIX1i8ItKaNtFzB8BWwqkbLTwD64Eu/t24S
N0hsv/8mtypZbnlswPv5+7hXbW2dcvEremuT2OEkzNSJnr4KeVNtGuZqzqKtc6LJ
GGOo+aYTbhC1mgVTm/N9iIlmRKjLV+h0D45tOd4gKmBfCng7qqJyF7Pv1cjfrIaq
4XwDZKbeWD/Gy0EGhNtyPMjZOIQS8I2nVQ6hhrvcPZwvQtptoiz3ItELDuruBQbf
KdcAl5RpRPR4Otm79JmfqgerDjsp3zMqcEZKTtenFTtJWERiKbOU4PEJ21TY3NX9
ZOov7Wtgxl/uGIwfQ7Z0WDrhsQKUSgHpmReyNacJiO2B6RHG2Yeioz/KlB//g8SY
mvcSjuiMd2vASqf6+v0RMxtWBg2nbVIOOAPIwgIR+Ab6EkHaNGctiz2CXdV0n7w/
nrhr0cUnqslX3AV9MOa7LBv5u1EZJ1uNnMzjEfLpB4tbXlj+ReJ148ODC8CYRRRY
qzATghe9DBoBV1f8k90fEJJQwsIGQ0B7UVymli/Ml3m9an2OcYlyNdeE+2DtdwOl
U+MBfPfnULcmDtVf/AvJZIcVDhZuJm5EG2BBcMTT1eNLm5PAhPKW6sQL9GPJ6q6C
QSTicfhPQD9KwJubVoQcsPsZL02MzolcWDrmOinb/fwohq8CCp/OtkiQaPzOV+5P
7hR84xCUmUCmmwGVOH0hFN83DiiHx3AQjciAkSDwZCBcRinIXZsM16FaMP+xDDVv
8Eo3Ye/Oktrwky83W0HIBL+4qN2LBBcbCEBwCOo+CkxlIwej2txwSaEEwNR8QfqJ
4SG8/YCkGdVNmhbrQio7kwnt6l8PEfc/pCkQmPcCj03+MwuJlRHTvFLSPVwgKwVa
v/HkxHWPtUGBzITrTtSdxQjckurJTiwixnmjTNN/ZtmlpfuYqywqRedM5vTJLJWa
S5PYViwv+RaZFN2Jf2m6ojbRHuwn4xZo16xT95eFgijipakCv1+Utg/f7ZK3DUHl
PDEGbwjRY99cs6osdieicIdBu55bTtDcoC3wcOxSwSCrjz+fMNdoShQo/9F6JFAU
RNVd1qxP5QKc329/zZJg3q3KuPTLFTNeaWtJL/ib2MYPuT8R9cpyGmjtyM0ZtdU+
J3nXb7jNAFQsaK09qxyI/DYvNTi+bhV+sW7CYkBLXFlY8CVpxPnAEaHFM9sg8b14
gvNu2ZrkhwIYNAjXdWnLecaluQsgNqD6xpC+bhIEOj2CKx6oBKejS3nEsY8nv95N
SQIpj/AAhPefS4NbTjTggD0JQQDD1KYgq+McaOtqf3wfrmCLmIEVZiOKoRrn/ClJ
5Q5tKmdoj+KkvwFlYOLa1p9ydkFcCDkTdBHc0rXt4tEMF1hUewuXPkua1r/zeHPS
arKLSPvaqyjftPjrLnQ/LeHSvg7ACmzsp10jtUnXDeDMKnQzfBr5hUMsrQfCqOd1
rxOaVVQXssoZJYUfxMhjs5hYkyxHHJTmQYq1Y23P7WKR6ajmGSK7sosWhXEi/8Rp
GdYEVeeWzlOiCdS8R1PLbHvw5/jxK8yXjVHRbqoaCvcl7859XYifv8WlDD6NExef
kLuAQV3gWJXXP3ehqZcT3F/Z7TNCbhXI47DA01JCD/La4PcBezzC0LKentIAHKir
CsgEhDLfAndzPBVo2DwSRcUdWlHLZdxS/OX9G9lpVp2SDUbn6VeUFl6eLRnmMFio
GCJQ80yCw09ASeA1MTqatEgbboE1i50s+IvqKT/pNt8uKp+KViigzwYrH3BdqIZi
o0imPaNcDqjxXIz81OeSSLL4L8xsCgg990L1K+ZyVhCrIzZUVm9LMzkAS1woYzOq
b/HDvrFoiGzT/P1+U2oQCgLM0HIc10MAFZBQ7LIi0+RY1Pts/Ip+jBW/0LrQSiXa
/lqGSZL2cZtaKDgYz6jIHl2H4CKpm3Cbrfbgk5G0TAVszVcqX6X0aLsPPAlqOBkc
H8wgayUP0xiIqGPAlrGHtOT7NvY+IQJT+1Pj8NwAdmDeL7T7Zbz6DDlXOWkk73k3
CpWK7CjZWawAHB065ehhhkBmgaNFlJBz607dGbA/L3RB+osG+vGtiJogxJP8uaMy
r1oI8iVn7IF4mP2quWLBsCTtTICtZ2gsANSOGYlxvfKqLPGbNvmF8dqrO4bEvhTl
b+peGHETm7CtS+OqRBQ8QB9wy326OLpzmKomSm/Zy4jV5ctE3TfgRYovM2yjMYRC
kzWqNKUshamx122e3E2CbERxUMUSgyeUvOJ7kQ+ZTAApUnUVczSXpkyhD4SkbzGT
lvHhWX4EJof7pYQ/Enb/NgSlgLsm1YxnrWU5MsiKy2xN14dpRjW1JMLyrpUsrZFH
H/bztcI1MFDT2lsvjk5UDVMXXxDbw64TztvEo0H7KpCxNcDXtXg+H8LXfePdZbaD
BTPZmsl3KTt6xEEPoc2Vh/4o0Hai7wK8I/mAbxwLHUxakwWA1Jy9njini6VhOL0N
6J6o3PB8MikZLNugkhS4NplvohfJ+IJxGOf2eNq/wV76l59QcUl6ZlZST5mH3WGM
KqEM3KPU7wg9WVnTSYBxqGpKIiVS1dMpE0fzNjbT/c6FWPT/4ZW2YxaeO1n0d9I7
uhuXCMBDuvlDasfBf6HdfIGIHqpZM5iIeM3fiV4UVRgPuCrJVxZYQ9ToRPVr4/pZ
iKau69bE0M1kyHro0yB24H863lEBdB9fJnmFLAXWDTq6Nc/FrmFUvcVUUkKtAKQP
Wa6OWpQnyTrj4bkolt+fnCmZNeDs2Z/cIUKQoLodRhS02m96nU0QZAe8psD2Snf1
q99nVC8q4jnEImb5y5uK0ZeqRFnb8PdX9+8dGysois0wLEigd9ZjQs0wWZbqTAQc
t0LOd7s0MJPzWFHmy+i7CDCaNe1VUuVChHY6ovN4tfU0GEhrkMy7FDVd6IfK+W/o
P9zA4q3h0D1b08/j811DZy4QlgasPCEJtV207fF3H3L6Fn1v2btAImUxN+1Mm3wW
VIiWm9ksNPfje7oW7z7E7G/PiOTg5oabqQ5fsUSgfutCpo+Yutx0HVz8D7BVBR5o
+L4eBrJGOPOmv1UD0DMp9K5pW4p5CzVXxtCKITk5VWDPBHS2iqC1nAtRQiNmh68X
N9twghpnbouD9vTag4ZVx99bDSMmeXIIo1PuOn+shkgLyETeqlFo+K2OWiPGEb2C
yahen4+UsrYRxnb11YOuXyHgUWymr5FmPnU0Z0gVQqiY4r2VF8j8zPB05hfJdEmG
v2qg+bk1Xa38lEQcbQhSylbXNfzaJbL9Y9HCORB6BdiH9+DTHv1XOgKwZGKbuZfT
zCnKcHs30Tyh1oewDmlbIYgpRe9yChWjBAVjQdjtAN1WxOxBvj6EdbVmymXr9/WO
xgvwR+zVSw3Oq5LlaH6uWk7ie6pVKa7FIk/fAburRA5EkuO82Hyp7SugRcF4/bjd
UISnAwhJ8ts453ymCTjMvQyjFpEw0agV6krs7CEOhr9E+1eiIqosIEyALeMQjNUj
jgQCeB9vZvSB7zICiO6ybcHHRnG/FBQhzO1OwfFHezHe6hy2W/WKo5LIQS3Gg58k
0QJK6MF4XLKggampmIIQcbiSfkowDFwc8RTB5EmfMf6/H85GFO2lIPYfWxyI9C+l
4ErUfI57D9adi0Mt/HwAl/IzY6C2sd0b77Me3vOgQ0zL4wxRbp07aWkyWUA/vM3p
KIvCt+by5g+RSlgzs1Oq+UggwBCEqjA8qapAHwGg3ghfyfPdoZBfheZ5z0k3Czob
RyuzZA9M2J1wu27DJEyRQ1AK4PxcCzJN39+7CGeePNCeCId09uQDclfAMCi/bOPI
hvncxKRD4Cq1+4iJRWVqW58LBhqZB9m50gwJn+WwW+FrsApaqkUyFnv3EsEmY6Ye
7VEihtv8ViU195gcIeLAkGlXS4uvpuRp650I5hV8GpHhFsihrwH+bLGHVOms+cpw
yACH0FDMhrR/EwhBmSq8+9KlKlt3cx1QWlIlQcJOtCGLO2OkBkJkExNo0OQ1rE4v
Jt5a1U6WSKnKJWlGAtF2166hm60kaoZabdWVF5sN4Fi15DzD5gWeFx5x29RxnyZA
Q54p/qtc/HMWd9ohGNdtHLeoi8pQfeUyc4Opbup0SUEoon4uCL/gY9il9+v5k6LG
I6Bf11j3cpy+mUOaOxHZYVi7/uoPe/qf0Fx03mn2v+sLMAjFqU0ZmvUE5ipEzV+D
VNPIqzqgodYXIism5lWRvhNunTtLceE46vaKSy57Roi3otvsAiX62MZrV4JkqdnE
fUcPpLbIyAadk/0JcyrTXEhS5scOhWQLG9SKOXMJ0YsCGbrMO7EN9uPODBCNHj2q
Od7QGJC58bXqp8jdJsYb3+navVlQued8OVEjA+3kQylCpmmnwLR+D8RWWNo9PI26
Hldo89qdaV/4m4Mj83W2VbjrIxR5zrRtTSF6AHwzMJaGWHeNZygMuYbYwGSFyLuH
zAxeCtbMBXS7Nxi3jZB/H84cohM1v6YMSbXsGuHaM9ZNVqdea+DuecvAm54oYsTt
A4G/d5AHCleYhaAyQ3TMnmj1nwk2gs+k/R/lyRTgqrhuBglB9YYd9lCf2apPAOl0
hsEuFwbESrvw3w9YlMRW0FVHgidNw5cdNdPM0WbJsYwx5XjgYe4CvdtSs4cwSMk7
gv27+9D6okXbNA35KIbfeVNJJzxI5edU9NCUeCeThEG/0BOd3mGLxHapf2t94q34
HLsTafXQGwyazqk1ERDPmWYNHptB8dxdNPvaVwcCAjAfig9b3IAfMOVlhgwvhAKd
PpilH4WtOzo5Iid1GWL3cbnEWgy9A8cm2K8cwR9nOfAuj3NZgtj0phXg7olxztz5
xyECVoBQHtF0baJru5+QcEKIKiylKXPIhYh4eKznqoeF7znARn5krndKHP4Hf9LM
vqm1PapvMSibHIKa4JwJupzUfzDSxnN5Sd3x0Ifdr8ebYfADKjxnSvibf8BoX3K/
1D19KbniSbljBIwnfcxCWAcSr6zHs82cC4DSPade6gBm4oT6yTYbSV93lGe06oXB
y3HkM17tMCzcGnecSwCYxz9pnldHodCwYH1kPJgL2yprGreqPSxpc6hstVNq8MZJ
zFJDuAiohL1i8j60wJEKQ3CF5lhEtlgPBBxJrU71jtloAHDyht/uhJtNJqrBzPd0
Or/lm/f4NooVcQdFKWgJCu9n9s3E8VbmYQJzGqEZcQILW/tqmYbd1XpGLQG106IR
YaOfONX6AJPG3VLbychpR/TeCICVdV4wWzXUlZmQtE3P1mbV8XdP0ij1IhrIx8PU
b0ZoZx7iFpY9LScWmGbDz01P4e6UwW9fxP4sX7snwhHQZWZj50yed43FFUfaHTol
JsErZvRcRhzibbTARfVQTtN0WllY/d3gSf4/m48aBzc+WBH6FR6UICKuIR4QrAtO
O0CAY+q7cChlE2AiUDItjoFakIjYFxCGCwA2umH0aWxzfgVrxUqoE3UaFPlMwUSD
yS9cKlCOWxp09NVXBpf4SkPDJCIIzt/49+7c974ObDFhM8ky5ZUOOedHmnmFsKBH
i8BjXeSKpRstEE7YY6cQMjuH+cgyY0YAviVZV8+HMLW69SZEfbX1VYPyFEEg+i6n
fz+il7sN0vpGJccKY/T8JyvR1hVhbYqdyQGjbWqbIF2E/d4YZyVIQY4N/irh+qrG
JKl5BrQvNDiU3l/Lpgpnnty2NYNmoEfpOKG8NIFp2uy3WHBNBRP9RRUxJAQS6wq8
/VDnsI3wjYjrAAkvSEy6KK6AWn+j51OoeV+sKIKM7ANFOxeJRxJ+FApur9j8gdtN
dpcvcjO8AirD26eLSYoODUF0PlKIKRQxULwf9Kw4iU5ogOvP7owKebWSsunf5oA9
4zuOycUmEJic/OjNBVWQR3yswVhQI6Z7ZoJiL/B+LVBcJRKlg1SbftUF+/yHd1ah
JEdxCdmUNbCY0+txPl02XG8YPWhylU59oILvNMnTysZxGMbjoD77KW1+gUpdD09q
0XJ1HUwng76wNEvLDz2mT21K6BeAQ6abBLPLjeQJnBS1JMrfFsdq6IomZ2fO+whB
hbikt/2MLegkpI1RxgdC2uTjN+Hb0qYDNQm2EzFg8ThT7IyPE3W3VM8LtlrjMmH/
PDNySnflh51HRHXGOWgiNfZGEfMuaspjEMqxVz/4tGlPIexDCnG/NpB57vR4unxb
3bCUuYrcPvzlUEFmH43N2RBUHFSsplQ6wopAjjBlFv87/4zTIB2H7+zAZjtxa+g4
vCamSZca2XMTpWmYefCuWlR/oKAKlY5OqRvoAOcSN3tSUB0uYqXNZ8GapBC3E4Gq
hwZQpLwv+8+7L/H4FEu62K72Q/95aXzxAtsv7RbZVl/5FGZwqF8WB8xAzKgoqSpT
nHWHRO85MI2VcaN9aYO9qYSRznuvynra6eXYDhJP5K/7UGuU5cXaFIn9DGJc8CYE
J0Sr+2Isl/kGaBamkAD8TZKnCi3dQH7qLH9S+Io1bFdlO1Rp3idabtfePd2A2e01
BdSaPTugFQgt6m1F8rxPDJBFJaUNAbdHUw1ohOERjSIdsxRKXURgtDTvc0P/NnkZ
cq4qa4J/HT0jbM9ngs017oAICG4NcwQFwD82BhHezJqghFPdJb01n027n6el+OFJ
2CjGUvpAw9HlBwkgbTB+OTIH33RM1FfTJg6IPlQflH96MTHQOHwH9QTMg0hbDWAT
3GX4c9vwuBVNXtyAmF5bCMBdWUkQp8cNZrnAVHl/WWe23wl/3OcCy9OtsW0NLZWs
+vKlpY5dAPlaGr+K4Pgq4REQpFzcRwgfNvTZsa3Be3RiG5TNs6ydRyq24JbYuPaD
UylGgFAdvEL53BSJGoQqqFVu6Thadj1JgJkcaFR1/kSissw7Il7m6uhrITrkmcUN
8Ma0BlCK6Xo6b9EOKO+WrKtft5GxuaT4wlCjRlMwWSicTueldK22ahJpF4cx0Yph
mlupoBTSB7y2u9ZUnYm3wHOm44ZcJZAT+lI2Q23yYJOuu6IAt6FAsdAfKz0UAS/Q
apbue9ucJjkXbBCBMOUbODT1lQig8XcVbrEBqSHtA1DP0ZgyvvB/3iIoaQgZVEwI
d0mUPHNUMmKysvR3cOXQOrQWNVtKUgfiswr4oesHzeYLNmdYouxAdnbda/4jfHQj
uuQ5t+2YgA73DLWwN8Uf67/yW24NYwgVYf3TM+w8VpnnVtzIEeorTo/NGS2aZ/Lm
8GrD1vRcxEajvlnaF70UMTLpAWdOKPHnbwHtyHNPW1smK5dKp1zfWFmBPMeSFCP3
ZsWJPP/2Y2/YbrhBJkQBUB3e2SCG0yrKSLHV/BO+se3kEKlQtU5iLv84ULzzwY1r
1BztZTAFQTf48O5WwQ8UncFgu+iOg2JdFigVtdc6116zWRe1DS9X+HnrhKEnO00c
Dy/d2uCwnjFTWSqzz6IsaHJnkL/OUE2Bc7uAbso2RGude99oYGr6fJUhifYhYGlK
8A9eFrHxh9qX60folIqclkYl3hRpIBq8JYt4YEac9cSkSxv1vMqyVItELJiqoeXM
Ba77tPgvKa1N9Q/PUVxeWaBLn5nRcMu23KJoSkXqIRd0Zj58o0EbFsUZUwpoPhVC
eotShLj5LS3+Y0In1srqgwYIyOLcwYbF41RkKSW9XtsL7/AaVlyn/pthEPF4P8rV
bor4ttRXoJsSdyysF3HMBSkBiJ7y1VIugyshaFuYQXL+O0r+MYODNEGe5csWravR
p1l+ilLJ9gA2B0es5M6/boy82yYDZI9B9mKuzPFvaEkX1eIdWWii0YN3vn14KHQG
o/mgMu8Al2vfhFbUD4uQH9hXvPSYFBpkmK3tevSUe9bV6/zuCipIz+xikTmxWF2O
XsyXIyqRs1OZdFjKRe563vw/frCjq8KMvcaaCgkuecUelgGxar6KaJ8g2Qn149dz
tyjDI3qdO2rGPq25E5ro02npPhMk+q1qf5xA5Hr1vvhn7Tw9+X5G7hlhb4Z+1mpT
Ecz/nFmyVaXldGl6LyzonzjMiQdH6wSS1l08c/aC+mBv+Vy9nT9Igp5x0HaA3Vn/
1l7YzVGsAcMpVhZDdjSfXRyVByVxImi3uLz4pyC8Ca80KUrZ1sPWmggts57d3IVg
qCb++h8IHelpdXgzWLwvcMBc+9sNxzIDWMsfkDzqYlr48RSD36SQ5d4t4gVMvtAH
WueJG7ImdkFFRWMSflHFZFtLNfjIUAr+F3LQ8qcdvFrf36NEviNE/XdSvwzyGF6s
IUCmDWHDJw/oJD4qbHKW0XSOcLrVD/p6lXMJ85ZVXrj+OvOFvnHt8oM7K+J944lB
rYDkSO27F8XmfD4KJAI6uQszyGJ0HMYVg1V15/apP17PdtMv5sUP0aqwEVx0kUJS
6wCDfyy2a2LRMPuGEjc0mkgnQinvFpEPMBvVQ01nZDb5SX+D/qWgdnFYnCH4/rr5
G5gjEo9dIlffAjULG9zEqV2V74yG3vyHOXoHoA/kuK1XKVWijkN2KCQw1vJYIZ9M
Ub/wyzjl26namjIRbWhYzmLpmJqwaahQpIG0HHpjV9Tw/X5MpKx2gB/Hg6ahAUbM
GPx+dzuCIaHCFgrp3c+ECvf2Q1TcGljzI5EIlFwUqE0kKk0cOiM33t3HNVv55Z6U
dOQa8X2vmLGaivE52hjQIKtxj8y3sqS2Firk8Rcs0UdbZilN4Wh0gbPM7oHM1o5U
WXMbAm1ZgHYgFozah9jIn+aE2x+5zm69I848jA1qLpXsF56OHMAQw7Aiz1iHPB7E
YXdfMTt77lkvafBMHPsHiQ1bYqQGBeAcBTL6eyryl1XCNi4NNdm70sNiVKaCkLW+
KkHIyZB3OQDIKeLDRfz9nVnypGv9BeBZZxqWDZ+i7gnEFUCUWamj7x+R0E4wkxug
Y1Rt6D0KJptC/wTZe2pl3wM7F5cZ3MQc5DDt99AUKYsundZtZRQzuA89TbzVfSRU
uqHRpd+3+vcQqbMjuNBPjTlUfNcEDAR9/d+EFGLILgQii6NsHKkqlZzsssztsDNj
HZCJ8Mw1ePZ02JlF4supveLDaR5idUGP17UinzJuyi+90waB6ul43gosN91f/U2V
+zriHlSoJnFlyqjSOCfrFX4Qw9QhpB3WqjSUdzHNw6U8weQ2Uil7MJJQQFoQGux9
JxRpJp4EviJsdj7KT29TInRKrjDePE2z3Ra2/SGjEhIfiKR5scS3Fx3/ElPdO8rT
YW04CWJ9rVCqDLXv3hr3PiqXl5mdU/DZwLLlGkCp7POr4b8JH7SAFXUm1vz/BREe
nja1pwtBb2LgQPEnhuiTFGMHhG9ZPWyBhZGH1+U50rEJ84X3Fizgulnhoc3Gqtp/
bEOi6AOeIUTHnsYYh7admBCeT48WRMMOF1u1q7y7w0ZfqJiHYhejQFIdHqphUwuG
mitCHmTFNifC4NBbKA8yNM9HW6NH0VxWeztRAILQlTsSfmLTYdM0BtvxFvOCh4gk
OtWPMgFaMuS3DGdlO+PI1oO3Sd6sPsYNvlq4C4BbzFfuxDENT2kQLsc2EI5bZvFn
FmI4aW8WKWgLLeeFIgwdd7YBdEWRJfzzxiefWeYsZYCCiAIPR+M0vd3w3M3aStrQ
NprXswJLEg4tR1vfWq8ghYdjSos/A+5WtoMWyq6foQukVhIEEITRO5jGb+3YYE+M
pbAy0ux0U8X3BdxBWsL2yWnHC+XsineCPW6Jc9ZzoEsbRa0cHnBoB0Lf5a9QirJR
WQdRrnyq+hXuch3ZBmOq9Oeyovlxp+ljlc8PYPra/zuvPRuu6uQuUDZbqh/z7QKP
sOgBK1wX53c0f1l28n5sICrI3kU/wcc+EQU+4JJ9C3JLHry4lVLp0rx/S2ryRoZd
5NW7FUHvwnT91d5UpupMJ5rlqPgQrpDblkGutBNYJahN3S8VWLOBmy9bHiJH8sws
VbxDedlwWGwmMBbihh0EvdDv8Y9El1CBIq7CGoR1APUCm8BbeZ3sXrX+DnTtpy5d
t2n6RUzWbw6tQB+DQd4n6aiFzyxSRJ83ovHNjUc9DtgSfqL/JiQhUchpeqfS8fT+
GiLE3m0DsdOWJ9X09KXVG9uQzL3u9gZMEo3/9sM5wML/umvM3Fy2VSyS3e1pB0Ym
4e8Uu4KLt85jtphVvfHzQ1+pvBED5khokToHPQHfw6RcLHYDlgaXCCCmxgJ4rA4I
FBS92Sf5aHR/Prk2jLO0HeZzYQIQmnQGMhwF5589MBxf7GVb6BZDCfkB/APu9m3Z
AE+Sjjwi/a1wccC2SNMy/+SDVW8fLiW9M6vRnpczrDQXTWpPN+bdynHUgYnZ2hfT
3GZYQ5BamwvATUJt3w2cEx5nPhnIa+83NC2exv9G3cdMp6b0l53dHZE1n3wa+agV
Q8RCNb+a4QdGvguh7zAzSp2M93kPR55nfXO3c7ipzKYojMiceIoxKV7E7Xxv/UGA
ZWjRShD5URo1xWgz9j4QGwMmzP1Oh4rLGmclhIjwr6a+5vkJ4MNig/lCVkdLxyfu
apP8nOvY/zersPEy3EU+D7nUdlOF9ebRj4e0FLI8U6KmwatD50e8ga0j8BajocZV
VEA+rSXdngXnj2xjIUWzHsQGSeyu8abo9HSwos0Z94d/UwftFMpzTsixyySteuFx
PFzHpjvZvMjcmrHT/IzlJvjqkBIlx600iZg2zk/vaYMQR7OsDwPlPw8GeoQU/qdU
ziz3iQed0F4g5Tc9izOg+HoxejAzVcnjNaIcsK29koI=
`protect END_PROTECTED
