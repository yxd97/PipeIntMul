`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6ZS0YWigdVUL6QyENCs2/auo0voSCrwQNFcBZ+s2zCoeMEXQeVNhsUeCV1gUs5X
ffRnsaScux3SpBh06DchogmCVH8aBdsjb7fXQfK2MpBZwXosrU4tm4w06hhgpODk
pWb6ZthAZcRIxdS3FooGemxROt03q8BnI/cCt7TITnj2s2bO5cw/2FrTcSteQdg5
YFMcV0y2WDud4YcvW+iUE5AhoVmg2I6WizZZXEeYE8dVzCEiqbJ57wCc8OkB9MBM
W1RCQqIJ2hgHW/KVNNpQplUYFNQ+xj2WqL6sawkQ9WYyzBv/Jp+Ch30uCgRqD7qL
VjyjA61AMsvY29dKHhRgZpfOJ3GCmkx+v0EkI6EN+/SxQvn4PNHDi8IQfJL5VEDW
ePRLlY9om81S9jDUy43lElYKGNN9Yd25oV+CCJ5abDnx052IWTHx4OoGkS5ZYcPg
6J+cQbhShP3EycBNQCpeuXurbdbLWBMAa68ErR+IkCtgi9mFz0Uw81ByCjnGpJfg
smIWg8G/Nas4v955sydzvCW/goMjk4jrJio5fGwknxi0y1JNd5dxLGsUkTbOo7FL
JBYP7ZeiwK21PmwHxZDgzMPIi35Nrqh9rP8PFtaOv/FBUlA6wx4Vpg6siKL1Pgri
Dwre7b/3xgO5jv9YurFAH3GXUafsoeedhYRsSJLXSdkYy5A9MXf97Gxed2POiSEe
KxQA7Mdky0V1LMVzbAeJ3nndcMSR3bki9nvm3fP2BJxJCRJXqpWSnPULnVGQCQLy
cAjHX3Xk2uLA7OO3W8ued9QtA8Meq5k6kkpf0WCpG0K/eYG6y33dJ6dIf65GKQB2
e1PMgnBJqxoZu4jDR+osdKMcERcF0NOiNjqo/5K51ggB2pCymWrRtGnwN+OJa6Bh
run6ZhKEjfyKOYFjzgSGfalUc9sQ2iBJAAHqAuEc+SEXr7Zk0to5szrmVGXF6CsB
Pke6g1tpaaox4m/kL5MXjmUzaRv4TqkYcWN0SFEFYzZfunpWvLP113rQa84QHiQh
UsEY0Jg/K8UWw9vVyiYb03J9ELnRqJVHfPJeDpSUK0ldrQPmFKsTWhU549Zs7SyT
CfQAGAVl2WJFh7kFd/3kJXD9RwE3nSe9kh92FgABFOAgDHmO/LqP9S0O6kxdSfgN
maLp2dPYNOXFX97eUrckyoVVhCXiFq5mlFvO34WJyAu5YPnSyVilUh53wANFS+zC
cp7VEuVOiThifmHtiRn/nOXPkHjEgtxuX7Y9vELZZTHxcs8GyY6Dop7+LUjyIFyi
JU0FnMAgnKgr1uTnI1usBhNfUQ4siGFfGfBCpLQyDxQwBjh2wrsJrwWOVNyE2OEq
G9x8Otc+WKFT2CCJmD2b8hoRZC8CEnLfXLBdQM50YfM88BjTtOPOl5IlWwBXv1SS
AmfRvy5e2lnNITROYTxvvPG8XamFQw6am93CEzVZmakQbIwunfYmKbTZXz7bg3FO
ODAaPiRPEs5nxo2meG7LN1wLgfLzTTmu/xrpD9L4jHzDerVao/y5ZvD/YKeWzcOF
IXzjBXnSnUkufSqpf5Vdkr6agR5cZEkV1gqEC36AKHz2MACcTwgXaft+syGdkBvm
rYkYezMMyutyctpDFOMne/gdreFezjmK0w9Ip0a+64k1nXGEGxBwsRzIesnkiNe4
WroFbRjJZcOUFkZ/jTpHtXPrcQPpYQ4FG1YgqEysZsZtlx9JXZ8wDDN1iSLiR5wZ
E1WKk4b56LD3KcC3v2AIXYJ2hUWoDoScpJTwfyQrMgWEYJzKQpV3RSo8I8NcFk/q
vHTGfO/yx5Oi2gsbFCG2tiAQnpcE6+z7WZ9Rb803KXS9zSRpNa0BDg3WGiyTXcDc
ohXCFavlT2O5hORD3fRGfexQpxPd1EbJivKH5dVeeiY2GhLybPPqnBIIEGGXJdqQ
0t7m74g5C9ryJgXgoC5y5Lu/4WhjGUV4+D4p36FUrZM=
`protect END_PROTECTED
