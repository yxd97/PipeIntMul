`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsPCZIN/VvfJowKXhtqtSdneT7tZHfnH3SyR1utKhX5nR2eea0ism06RON1SfKWm
NogmgIqGrdWgXS+C0hAqZr+8EXc6dEj1qyUO7n0IDWN3RiVjCh3QKUF72R9UKE3J
5uJ4IlLMpndbNdgyJuDJ56V9zSsJk7jiW8TKu+TWp75Z6Igj18rC9fnoh+MMuDWg
M3XjqqiZJ9xX9zPHyCiOBjWO0c4TXJIsmlR4+SKls9qyHQW5ZD5Rrfq2rAMJS7TZ
irGJ8SvZLDJVbHh52Lft1ick7G0f6LKavVqfAB/69WVkWzD+hCdnI24Y3t1LTsDo
xTSOx74Self8PhR5aKTdq5ud+4se9TME2sFGdvFwb93syxmwUSnNr98BrPIwLAXw
`protect END_PROTECTED
