`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HOeVPklcSn15dcl4i5FnkF6/gAMemAVYzBxkp6smSbf6NGGYdfY5a//vauQeiPmu
NBTcwrgZ1ixkl2yPaZMpm0DEBuobIdX8vy4ISDt/4tMbwnY++sMdOGWc3TF9V9Db
tJEOdGx5ugikb7ey5rBQ6i32Wut2BDd3eawjaT0vHeOeGuRKyDNhuteCsH9KsZXN
cN3dHj/Ax/c+ckiM1PWvrhD0zgX/8kNa4e4orj4aGdn8ngoKLQ9AAeSMLTFBFfl5
9f/9vTIk7pMaunDHpvGgH+1ltzEcD3CdL1VffUiupjCaNGnyY5Xjpp5aT5wzT205
la4Csm4vV6IHVoiDvi7t0xVYTnmWFDtQtqLcmxj9zP4ydQ23pW3YW08k/2kLTEez
5EQWXyIe1QfJRh2/VHbs4RjWcWlEpyUwxh6Ot2Lx7zXoREvWkn7TSdibfCngCj65
yDV5hUkf4lnKG8inQaofxOm5Z4QUI7mmh1d6+NRqAUURvI+66tHkj1zI/iSZCYmc
YgwynYEPx9qtsIJGG9TbpbUtFbMU6IGOhiEEcuA3wzSkEqtbWWvApjv/MniwYL5H
t5B7ahMBeSISJxmzRpA1kFZzPdeEUxkPEGhfKgOobucCKH4NeDER1+8Ox+qd54xC
3rltL+PH1NrPO03EmiaXIA==
`protect END_PROTECTED
