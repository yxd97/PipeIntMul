`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M2FDAQX/VpTs5zE6lNBbBjvzzbWpxFOSOLCVeSsPVaFnBYBDAnlCOcg2Z8iNLs6o
f9l8qf0+JCe/gIAEnTNPzYZqERVfeSnTUOStUvPGpc534wHCSZwRzNhXZ3rntuk5
j/gtYT96rBBpXMcV4/lIHTzjuUUM7JxlBV4MBhEOP8dzBpZXpEZwyO0jXg+x9inv
heL8/gLEAiouDGPy2p414kSeC78Nl38h0didkUVBusZOhxc3HHQGXO2VVI1ANINQ
nOfKA3I8ugaLDqp5mrr/Kw==
`protect END_PROTECTED
