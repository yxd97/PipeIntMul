`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0p9KAkJWPhXJg03m+Ri8MHQ/92Rrk9EnN5RGkKvnudxkgdppIjGlUH8FOAMy0lmi
WpE0NdrOFweZnVHHMTND0ikJ/mRyxRltEXihMGzEqgDXS5QY8XDyx8pyRaWVBbQG
zi0lZQQWrJEi1kNWJHuaaN4seQuNcu6NeDukp+Hhx4qzI6Cj090zFzHRLu2IJo2I
eCnq2HIJ9l2E2fmMxS1B9aysEd/25Tru68q89SHUB4EzCwy1iNS9zz0mrHT2+Bo8
rToLZ8faRsQMYYZS690ZzqK1za/Jbv/3muRcRsv/DkMVdv00OqO+q2i6LDu3IRqf
T+0zIcNC8egMIC6CtK+p1xX64dGX2gK8qr7z/qp7KKgN+XW5L+nXWyQMI36Ue4qZ
2q7jfP20IeHpCeGj/guL4kdIr1nasqm5Wa4lCmxdX8nTz2NGyhRUS6AOfCZv1d1B
g7fLInBpQKYN/iuUGWSgXslQUSgdmFmRBPhBQnGxlaxmKvvt9UiPeVC7SOfthQ2E
8Xuz4Y0o0IeLXZQPOJM+pl9vulzmmv9jdbnDViLVoWm838DsYqzKvPpBHuRrTcWi
Ipyi/WNFweGM9l5xlR+2CDFnVL8HIPdEwA4jhOXriI+6HQGu1QojTcvK2+gmq9Fd
OqezksvE6PuARJw20c+i1Ti01BOJrDrxQBy4QEYI2xP/lUo3xA2ldGNErDoS0vAF
vXwj9PAbZ8+BEjJWUeUrzEV68/YitOJumNqp2t+qurJK6UosY4bif5sNd6mPmErC
MQL/UcJOsGsN8vVbkqEiaC9s7yaFItVhgQOtUz3MDmQNhRtHQenW8YNh0iqFZXwt
G2lwby1nc0yuW5QrqJzJYw==
`protect END_PROTECTED
