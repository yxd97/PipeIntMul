`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWtHRUaaEf16sqhM6XhlU9ybkEJGxwfEViDX8INDOm5vPFm7AoXsSkyjx+HBBphR
d2rd1vvXlo7yfhw9lmNkv/xWKZ/ZqlAFY7rcqTCA0FPcJtbBeMYK8A9Ji7/s8BBY
GexuJ0bQ4ooviG0Bw/XThg5NVHOhzqO0vRVWJTNH/w4E2yg6YaGK1graE5Q5nrkl
6ljmY5pkEmXPITA50RnmNI9EcC6RKh3t9WsiqOXwswGbtkaUYbhJAgRGZxvfjwT+
VPEoAI7piai0RsNlALsFYiTe6MpQe9VG2KcEn0pWj6e9lC+2GFUe/ajn2UvcYfcf
PhV7gFs7NcryJ1+zavH8fMYcwDlAKQV562sFwiEGOYZ+fE5e1xMLDHBQiFL5Jp3i
Xzz8bYN+gCblQKIF4x7LzFjJL6TO1GdUWmMPuxnGnEm4F2dbyLMF8oU1PoOZX3bA
VsaZSrhfhYHFIImE9sr5nknegfMYKOdokvG8QHDTu7MzTg8f5bAQoUwUojM/Obd6
zzPKPXO+cAEhqPUskn/KPQ==
`protect END_PROTECTED
