`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZztABKp0oWxSl31gxvUyVlijBFX0tnom6roFRf8zeptjYWRlPMBPZEMxIkUi/Jq2
h8zBxspyzrgwsO3Y41p5Z7bh5XPujmW6SH7swE0zAXtbGIIexllaFz2xsIDDIpat
wPwm6jUMLza8ix4n2uCaea1ZDkCg0XegzZL0+IrSLynmMvwuVlg7oVTIHYL7aGKA
0jJbDO36ZCK3G/QgZD6HXrFQui7HXCWU4cDjG3VBcU7eOs271bmxcCFHjcyUCRA4
5JwX4d6oUzO5DzvxnAM2gNnoquZTqMgIHKA/BDY4PRv9jZaBHT105b/NNbIzJseI
yu1xzDYdkgNF/InCuMYNhn9NHMbw4NN8eByiAlxjmiIBiuXUJa9PE6aIt8Qtnk5/
uG9ub6qmSK2tku/ErirymYmBsgKTYeMMT4mephXMRJxLqyRVF9YQCaInKnvLaapS
1iGmEqvukvf5wC6xFIlkKw==
`protect END_PROTECTED
