`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulOf5iDbJHlZPiC0Egz7YtCJ4wBXx2NEJdmT4cuMR1LxdsOTvCPXc4erCwX5pJi8
OamAcOP4ItMvOLPFbjtmn2466MWfOV5rA1YydGcKQGSa48TIrG9vALpyE4HzBwvW
XRFXM17QnvrHXqZRI2cwYVSu7rD2OsKyzvKRCG2LUpCf8aaXHWYNoMfnThZgUBKY
JTdMINOPaNqTvR2vOd+boMIAnaG2jl6l+Nl2d6mw6aJX4/rihP8xCiRdpq826KtU
4rRwgNPok0uzq5z3tJV+ztHJ7inRFr6n2TgEsBD0ODcZOWeIDDtDzA55PnTSdO0N
xo20ltJnBVJIZa6yLUm17g3UF6zNg3ISYMGMPo3MtparzHrakDoFMOP5WoxScBwk
e3AtWjCQV2wvahRfx166b/mLCOj3UEM/9pdxABvug/65nsrN62tLsUBfDpiI2lVz
7REUAVLjpypN3YY0pue01wtvuqSvV+vbVgCGvboIKGo=
`protect END_PROTECTED
