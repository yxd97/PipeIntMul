`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WF0b3Uw/xmLScxa7tB7ntvGPAH50nT1BUa/PMSSkwPq/9zox3jDCAB/5LPuRD2K2
O2vOkpqWVEM2r1G2KkpEQswO1qSpTlLHn2kxZeYsNBYB00PWutz5GNQeva4GeDY5
czBnUGv0eNsWmfBQUOvlEYX6MOGcm4JmpnSKlifYu4JvvNbTWxk1BOgPCNfU28wR
1TgjHxXWOkL24q2bCRkVlHgRv4FZGKMONtKUSCabDgYxkhlh6sir3yh8H9LjCGNY
DFrUKFCJ7jI4wnN70rtogb59h2wcaLdfbhC+F6+ZB7zICzrR4XkC53SagAfAsUgr
2UDOIZfhkqABCmVMR9lX1I4SbMYnxHjKgd+L0xS6RpxLW4zOtKv0po5R8rJY4BrC
o8vQie3WkUoxU2NRVj+rurKoHRCl5vKuOGBwRGfCgkFuZ1RoSoEcQep6zgAzf9a+
`protect END_PROTECTED
