`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGuUOuwbJdd5rw3vKTtjff20+Xfag3J0ShhffEgHh2GBWBzeeAwR8IKCSzwV5pyY
FulSJzCFtY1dvDYcbBHWn5RJTg4ozVL46QTBqUR7rpD2CVIyTNPxZLk/DICncc/8
lK3rxNM0rh70hLBEN21A+R3jggSO9opReE4jsngLpEz2OEJ9O+DY9tZvkkGMh/v+
sSiVv62bTSQF98DWy+G+Kdcsn5I36pYVBIgrr7kJBem3wSS8GZGe1EHyuRHkQNPV
JoxoRpc/Vs0hVV0Zpn38GGWgp6pDBtAgiCIvpvbJogPQvw1rS2xeMMm5TLeeRgoA
439JLevvzyZkopcE7bFClA==
`protect END_PROTECTED
