`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
adiEAPw966+OtKfQGu2DHJsaZT1M+Nn7Uf6bV92ipXEPhE4cEuxEHdj08Ugxt4C0
xBPA8vxHQQSBDQl0dBwVSMDyhflHpi0DeHK+DyG9gZZ6QiOqc3LTIr4UiCB1ZPyG
h5xGeqZqSoTEEj1PzcOnd0/MvujO+IuiiNe9X7Pdc/DD7Dh8Hj68oXQsMbktBNfO
FvNFZt7arxzG5aDQBxvTE/ZqPnRkU22W3eggCjdKZe+u53KtTDFVHmEfBxj40vns
qoK0nnGNgRTwX0R+3lpfaCSGJIRaxWSR9QTPuxB8n3Zq2Nx21hjSCnL54y4c7kO+
UVkjNZay+3fF+c+sfcvYQOtSGNxP0ajutC/BR8xLstWv2YIQypCnWHcrhrurFFZc
nnrMGmJ0quyq0mO9CYeBjtqb7Y8r3xfF71t9tWkUEPBflEML+mc4WZrgeQfCvQlm
hB1AfIO+/ldhbjd/7lhpJh1sVCZbcN2WUC2M+gsJnSMHFiF/Ix60ilHNoQGT6Sg2
KzG9yjy9fGV2ZSZO3Aw295xzas1BAjZ42b2HmjbIh83i2HJx/s0ZUOl2HukKHd6g
2ImFTQPbWLDdhPLBo3as5HrhoHbcjuOFxynQbkQ9N/bR+xscdK0ZkVmA+GM75Leb
4NJC6iDqZi/lng5yvd+AYsI1mBzUH3/Lz1Te23eoctU8K4N/Hv8t8z/zqnf+PRnG
JBsFmFCVrC+KGTAppUqrVHcN6dMeeT7CoZmcPXllBkJzy71OZ0MhJOmeQO72ypwT
KI84QO2/PkkMInFkFcyc4Npnqk81xCJY6u4TeOEvzLwJzmFfAQ/hWu+9B465B3gx
hdUcnWduWQ+7Rm//AYOlcjAFnw3ydtvezjgQ1z+ktrxSOusf5p+lDZcx4nNrlQxH
OpEjncWuP/5D33KMzGK/7w02HHI61mRGoSLgZyh3Um7k9vuTXgrSvquMse0pc2i1
7j50BsO6L/pp4+tJxB4yGu3FZHO7p6qy1S2bcDpvfIVU48F1Fec6C9i4afQarZje
gGWuHUsDoUtyeVpb7uCppHI9MJJNy3JuVGiVrSnZUMxBjk2l3XTIRFqMkLOAoO7e
Z3GaGA0jcV5CSzG6mywtNRbjepGEe6YozuANtYSK2YrT5m243MjSFp4sxQVyqkzk
eMUovyrFvuaJoma6kRzn5Ifp3wRWUluw9SwSyatYSnb8xwVS3vIcoPYHYKtpOGgv
j3Ie/LDCNyByW+cAb8p4odFMI8NzQte0qiaVN/BqdulK6fJ4qWyPTLEf2JAEtfEX
aBDjMfCP8qyVhBDJiYqf+R7fFTpMDAIekRO3E0W68GI+mqv+1pxMgrVWIcoqppQD
TyEO1lr/lLnYEJUEY6ZC0xLqKcE8qwaTnlatt2Y14db1nPdqpFZBQe+QgwV/EfOg
NS/FpXNPXI4iVKAkoQ8z9IuCmxCNdWmum/WAxNjRfx/kekcWPnn4NI5AWi7M4UqG
sUghzMMLVExfp6L8GVWUOGDKO/NFA5/aI1g27R6Co6JpTTZChyinWQTc2EeokH4V
4V4fnUGSohn+gKinm7ReOZy0pbVT80WucO2fTx/ppagOL5gY1Xbe3vj1HKIaJwsP
BjaG8BW31Bnsp6YGOp6OEVkPZqdQPzuev8T034RJbjBDQ+uRohTDkXvvugXlYAn1
4e5hhZg+LFGfD0rYpzOVSzhb7HovSRILlTeOtLIy5Nd2DGqIHVh0wzGRz14Ag4Tq
FtFbrpDD4ztSJztnLUFB5k1D/249GosT5RwKVlB90xD5YnzTmuT+o/p2UGvzJ9Qr
E6j7MXs+Ia1m9YoQUbvk0IZzt3E5sKibcvwAXghXmZYRAnJylYSZrnF0aHmufD4f
te7V9QHrfUBmo7wTuHqJcPzwLWf86obyNgz8yBYsi5fiOSH9GfsO7cf+0Yjik6SS
YOXM/nBeqcTtlNujaZ1CNUi5vWzsSvIt8K3uE9MfaY4bdvEb0Es6s9GTS8k1fkD2
QvrbJmNEZgSS3ddn2gvAbnh3QbeRpM7GhU7BMKXHyXI74h+8XXi2hecs4N2Pep9L
3QjRUr9fC+IYpZvVo9yyfOqdVDSgF4b1f07uNxiQ6Jq42zX3Bvk5Iyp5JTNnIIT+
A5/aIy1yR/kjFTbZJbKK1S5Yk2SsNCl65/hkVk8Ow/Og1RfG2PKe89/O0R+fnuNg
w+TkE9OPdxmnOkJCahVDiyrWtO01knoSTLv9FSaU/ZW/tQLZgSheSgqb6AnnLaE7
/mTuGeYZd7DGEHwUtCmdTNFDKDYfSPgq/NiyXWcMXAXfwGONEl5ttjn7UKjmCNJs
B6jv8WmTlwLP05hUxZhIh+x2EYmL0RhW+i+08IsCSPYa2Im4vARlMeNn9XmyhnZ2
uKigANWLQM3rFCKrYjmHot4RJsH58G/Uf8SOX8fd1ObHwtKetLGN9IP2gkaC6wxz
PQXdFLomkXrJfBEY1bvQC4iBFxsE2nI0OIJjlJZpZg918GshkSA1+iYHudJMGzem
ejUowJHX2zDCmFCidBDQKY9kYmAGCk+mgK9C+dMr21L1MGVXGWdgVqi7rm241+Qu
wuqTLC9pNmI6YfvYfHc+4a0CEpbdh/1wZe+0JBqUy7SHtnmxhDon5JhNkmLB4f/o
nCzoZxeYSDVdgu1M+ZWF5j56+L6AwNX788n3n7+GqkulHbc/gKk5q7EJugmVJvfd
ycVUgwEayobOtg0QCF9MaoY7abR3VGg60FL7Bsh2mDmtM/IVDs6z7Dhwr/3zdANL
KEGSdw2/9WFlGL92PUBAotfPDLTZhcG5SfgHRsS6/Unp/TfAGPQH+ncLS9DLYuHz
6kPlepFql2rUVYjIB7cXlvF+S4Eej3wzV+tXCpZBDDxvs0X77yUoxmFJIbbuagOr
KTdXTHr4AHlO4y1JS08vwgQ4c6wgjNIOyY1e1oGHpN90NAws2pboHd1yFtdUeqwb
8Ls2+JxiP8ieuQsa8YWR6RWtg+42p9ezehKeVX6hlP5tstyR2glqltTz//G6HOV+
Wy9EMn47VTO7kIAAN8ZlWJMzHySrzcu4ELrVwBqDnsUd7iTvCg+voAMXFEeTigtW
Ry3it2G0dtM813r3qE+WFHSLKUE/TeOId2w+4Es7VYDA4NPlP+wtOYxlxCLcPrcV
ktw2ZF1i1oTFcOsuXcG5c9m6cazmy3gJjcHhD3/HwpCxJ32YmvceuDJb2OLZmL5n
0FIwBv3+NyqwD/9a5aJZ9nIpqONSJMD47pHpPQOnMDS7qae7YwsxYFhVpSntv6QZ
tYN/OB04ivNEwoMGFCjlVR4MtRuycKIz50FuCKZr11pINPNxwJJof+fx6xD/aql2
ChHvQ90Hk47H3fU3J2GIPij6W2GrEklhW7DT4QqUgSLQoqRoyeaNb4Qv6EsBFHRK
eCjI2b/VqnGREkwQh9GYxgAB31dhhce3jNkfsLoG2HAaZpBhW1v/JHtkLgcsaLqz
8CPinfrmuVvrC+bMS2YA+BOZMr5czibULyGMhFsFBNbKSk0Agj+Ix9/By4OV7Us0
xfkRtATeuslfqkJ79GU7m1Y5azT0Vy79IZ02Mh8Oj9XKve0QcUiuSujp3TF2dglc
vZB/az3FFYl/+LyDwYgH1KORipPHFB7FxMvtT9n2INiDVqIiiCjRX2ENvoZ6Rxv7
21S6jR1FoV1/chGEbyX7RBlBAJBHNH7DZOsPHEIMu3IlATvXotITinlgVnyUXvSu
FhvPPsAtillAmf95nshsJhCSdFKg6Ggh3noYBzms/o5k/2sAkb70bRq4m583Nq6a
UXF0DyDg0EkQu0JCKt8mfH5RUTgPN2aTqbnfhOZ1pVEHRRKpZLCdN1BXbUvJuCna
hxtEZrGZtpIAI7u+lHqMRXTsH1AnzAoOYZkQ6UKM7Fg3N/aCGTt8J0drtU8JreaT
2z6YA+gPXquaUimjK8BR2XeuJbsw5GyzAD3CTUoBnfsPyVuwe0YTe8h8eVI9R/bQ
2dzHosL+fP4s5GVz3RyR6apv8ah2HP0a0cd3+0LldOVILWWbcrV+74J+HqWMoXxr
WgrpJtcvQ1Ofqi4+ad99Rp11yh/T4z7v20DLel3xrIFAHEPxULcFdN6aIL2NzQ5S
sMTz7Np7xPBvJOw1y0fOKI/KDOUuOXkvGyND59KsBBpe4c3h+gb3HOdP2uhdhIoM
5tj7Uz3Oyn9OYHEgoeDuhUNst6Y5dBB01tEppilZbRrhGmfeBtis04smrat8o7cO
2U2POAet1lWuFnDL/XuHqYI4isQrbbGunh3qBORwK2OWAufjXlKKdo918ahbm4V0
vrD0+IDlDGEDAYC9SQ5VFV3UHQlhHq4xKpUAoMV2Te9dnw2lPAbmSbBFanyGkLM6
9zmumCCb5J98buGEMOxzlgZdCLUD7elkbFvWTZMqCxOgac0mAjpkMgCLMbVjEJ74
sddtgP173TfZ3QBCBzNpglZcRj4UfISM28Nxdm+NbjqtoWXuyrZrw+/B6mWduXXw
rJiEpBtnxCbq0CM34VJCm/rocOfgr9tb9W7chA6FyCIfENV3kYLQcli2LxxP11pF
Lkid69z9ZEdDHkr5pjcuDMwmnL8FSAHYYVNghbolxAWXep5izRikY7Sawi/qv/p0
eLOK74Krtv4cjaySwy+/xrRkrIG1G60TI2MqGVrLwYURvFrHadHO/pe02dPRRRrg
cdWJx6S/mfLJObyaq0IoEAQuLtrI70XEC7Y/pK2WOfzvoydJ6VLa28I6lpPYUJ/q
gje86XKIJ7iBG1gtWRkZctC+Dw7B2olF8pvDpuEc9PE=
`protect END_PROTECTED
