`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DG7Rf9JncNhmqnVB+sDLvW7rb9N8O/KcPE9k1udEZi/50Oebw6dkou0IngYQljuw
0jEZs9WDEfsVaCy5VxJhnxlRpSQukRkyTH/XYQ9gfzKvakR828ChxIpSp1VHO1xz
Ck+xFsupLHJU8YlNxx3zarMFh8IVyWDNYqUbN1tUN8oq7KU0HdbQ/Iqe3PgQ1+9a
+MLYwhEMbG72Zq7jrMLLi+VKtQIizo5e01461gDhaU3OG2y7hLJgazMwxJGA+sR0
RoDyJ+nKn+jHFwqbNNI7+a6K6nvKCmPfzXEJQspSjk224vqPRRzNiGpvRe05HcRP
K0SGcym8d07EY4Ol+mSRjNEOI+irW8UVQ5C7yxY4LihTHmPP+b/FReXjh/VigwEx
bJNeI75hzmtxxAQmgFQcDMWj/fS9dfF1sU7b39nUPw5cRbgtjM4P2tTqJQQjFqjI
DvM5XAw0JSoi4VVuz3NBMNGgCXZf1XfjwLMpWmCfRDFa253JFlaK/xhAufcqXUGV
UlWcTTkFpx40TLoUgC2k2qELMA1Wtr5jeR4anjCbwMLA+tAf3+YcVStHveuHkvkQ
kgp3Kq+htgOOLKlJTXIanmGhaWGvk5tIfCCnCdaB+U4fJDN6AAlGKj4uW+VGW3P4
ft1T8yeIIB98+jaJdE1MMyRdSl2q1yTkLVV/ogQ1cARd3QhEV14d6gXOqn10WKtA
lgAEmj6SiDVO5YaXK0vYEeMWNXX8OxGNrTHp9ptBmm8U5SHtApGZpl2nk58gRKgz
1qj/GDJd3l98x4rLWmys0o3VHcsOMiq5UHGEIwUEQXAW7pQDG2/yvauGUW3SC3PA
0d5rcM1zivoNx2id/UGkzctxfuymw6R4WYaMYY7Gq0PZ/US1wW7IYMlhnCp1gN80
GjXrSB/XEBVnf30mf+XE2XL65+RpCWp/qjx6vGgjE//DwAD/NC0aN8WL0VigHHZ+
puq/PY4O8+O3b8cSC6HRBWi0ewgeuWkZQnS9rsl2hPGCXr9br3SZuureBEkTEv/i
pfsz5tDz+DADCFHtgpTWUT0n/Xz07w6wM8gBAHp0CH9PkMirIpy/L5T9ZeXFK6Xn
uV0jPsokyAmNTPipGGK/oDy/BVUugrJjIrbfFn+hk2E2z7GBtjdaveD2siq9WO8h
Qg+416fFQtpp0N/ibmBSD+mubD+nTByaNIKaai9WfP2ar7qCfPsQXQSEpEIjyaXL
2iD5CQ8DOX0DnorsdcrKBTV4hGoK1SajgLbbea8S/wBn4WDfkrKvZsS6BkhNB5js
n8Tr9dBsEyAdbMQwReSVjIMuUyxJ6A7TNGzAn1R0iC261/UquV2xhclUNkzAt66s
j4SkZ3aZKmkHipInEC2fli0rIwJOAWbk6O0DrvXTBTusCl4mfjL5+LfMz5hJ1X8G
OlJjtBjF0xpGJQPVCn6zO0CMhdTAXQ1AhX3kEkp0pnH93Po7MjkXj6lik80YPkbX
iyXE93pqmIlGGKnYfSYWD+kNI7BO6xzTEVKSFYvOx0PiTBCMJUpVaijA2xSdgbea
3UALsDECgPR9vNI7tObL5rhqUqKuG+K8+C3E4RAGwiHAkV+mByn1hZLoR92Nm7rh
EUih6i3fwhM/cs5RYioWlhNhXp4KJfxSciZS6dBrE+TfDaSFUaIqXyJvDjjHf9g7
s3999KfFqLikGOzi/wLAaW0c2r+i8GpHaiEccYQGivBfc63GzkUhZmVnc0VH1WUt
6qQnCUyo4y1kKAaW0l9SiCdvIs75NxEiogfuhlREnDINq/qJwWU5sFDdObTs1jNy
PnzVxiEJxukuMcL//4zqZ19vZ0CSJ/SI/Pn8gbGRk5HhwdLJqCpwvB4NW4hTe+ni
Iq+3H/MEQ/g6oyb9IR5lJitP2Ns6fXhsuaeSipFtvcIknYjpgSVpxAAL9/qPAFkH
eB7m71wIz4kauJyA8pG+oGfMNOaDQWFW1xSC77QeeagS1gOrOXZkvq8JTBj93GGA
vDtf0QDUuzWPww/UCacDXdsZajMOfvDDtLEykKdoXcuAmimk0cKOQG/9km1rnlHW
EzFX55iKNynlfrTNsglMKAkJkGdQEwNlOPrJkys8lqGjZa03ClLcL+Do4696qA08
5dVL+tYp1cy+ZYOh+XLjc+MrrUtb+aNY11d3Kc1wkC3BrTbuVWh28Sq8GkXSEv7w
LnaNtdHbjkEY017MuykGVzXuXW3pgJFxa6lUhD0VJyVBWT1H99EE9zbrJnfAJ8rB
/zU191rE/W9TrHPEcLrxIgVJlysypx0Uyt7V8ky7P6VbIg0rKwV4vdi+q8esQlJN
W/+rr8Y5+bh3IJXDmhMiyls0eQFk2/FDD+o9zrdpyb4H4Jyn68tpXMDtkeE/2h2T
iXn+5kiI6EUCv5kFZuuF5YQcZM58pL+KGQUby8gc4Amk7wmDJ59NcSk2SIXAxHim
xxtlRLXgj30c+vwrtF07+sT54RSCRFFMiyCQs/A/+ZDi/GNRHeRnzKxDGQuvvEli
ifEEQ3ztEeH1IjCFcKQY3kb6rW6CLk/VoReA3fSA6nG9JVtur2M8sdy7N+Y1K2N7
CuNrIkXAu6Iqk0wArbHWbW+XVCvQzYhbVlSA+SpwHFzf655Sbxqt5oHRG6Btb+v3
MASHN4ZrAHJWt5X2nUm1a2wfJfJ6HTcf4UFU5YKRa5GTF81DIYL0HTna9J7B+pQ0
srQcfjPbhAhx5P+JjhC1/ge+RZTDyhb9YrF/8rwTnxm/Cjb/LzN1aev27PfHK3UL
8y+QXGVrJEOFSY5J+XuBSKsxAehOYJaI2Rrbm/Hmvac/tSVklkcGyYkB6R7re7r6
87Yg0ky932Y1OSJyTK+QoKi/9AtC2WqQoEeecRbpA+hjdyC1DpUTrhrJYvLJdtwZ
2OWNRr/FZwr+SLnAyyzychVpSFfIgyErqAbrgq2whMx0i2P/xNPhiwERGKAC8DDH
TFN6LgfxJgn/B8VshLp1jIk57u+VKc2jjema+epAu1qTv11GIE4Cir6njHSBTxnL
jqyubo1FaSo04fU5CHyQKc8+NN2PpjKVFvDJMLeBmce7RUb6lVNC+ztzrDIr+SZJ
4AjQb59vf/WucO/mNFWJ1SDcYYBw5M/x5N75MWAgLmNMJUIj+9H6F+JDZOyinXFS
8uotTLoEOygKcaCv5Y5RKbA2UQWxIiKdFoKfUIsKuDSg9c6gLOCHiRDdXu2KBR50
0shn5sR1y2a5UDOcgVerb2ksQjFsRJS64FejmldHUxiy7Y6hFssq2MFcuQ09SCrc
eQHl+9YekzW6X/gAFefdDNS0bnqqnSywoBkhtQ2SBHK3PsDtZmVmwi6uu0CELWOV
T0mTFCKsuw2QSFsv6shv1XMlDPCgO84g9kSTkTucgn3a7OXVygVlKjP9dWeRl28X
u5fwECEFXtz8xY36xJaC4yRHLzKwWNDceN/h9ZkqJJCjWXHWUUlaF9DaHFDdCXvc
UpHCew+BCpgkvOE09EdsLGSvYLo47rn05oNW9c9VmhX0JuKY7+KY+elze3cBUm8Q
SLGVKWXUGsLk7UQbWjvOlZVi4X9yuEAQIBma3M6gr3bU/nnzbqEPnmaQ3Pev5VH1
jDBfDTv1/cRyZRj2wgIzdHGbnDgs9N9Zy28vRiv2iPD/1Itbh+XiKihyEeF2euuB
2xEpQoy6jLsqGc9mp9f41MxU8XL0w9up9auqTl0pRjN2XRS8AiO7EikepI3UGks+
Wa7yUALeHwi9wpX7twadLUF5jMUTo+XWkxaDcuhqRCuf3B33Mc8ODq4O4r1Ko9F+
kmFTDkxrKko0btTQxNh8AWK/8I8QK7ai8JQsCeqqbo57RuKuAcZFUKwnYxa6oY9X
vWwugjfOoX8juRSND1TdLsDD7o5YXIEKXa13hnNHljI+B5nDm7H5qqT2GSUCGqHA
Sn/fQ+0u3IWKAkDnN8teaIeBVbAVs5FA+CTQkBGexWBBmpw5kr2A5YpnVm4LCpj4
gta/QfELSkUtNe2Wxfz9hLOfi1gyBJ4GnHa8Jiwo9BKqx9TMtcxpsO8zya1aHXci
hfUe9Rd2vSeSCS82T0xBmvv6Siq3E5qit+UZiztj+HTk4tAr8zPVmCLlRcca7a6L
om35YRYIxilszcA5JYIxTDRHsDi5L2TIamBwZzMGjOMoBvIMtzBLxj7smg6G2Bnc
dJUlOcisIHl5ah789QfyvzXdDTNuUmWhX6n4lI4+2CmMuQYSSVo9dHePNwoNG1t8
byQU6IYg7OX+bYxo8GR9oGp0H5jlEXMam/sxqcLQr/cHXclM14KrSL577E4NcBVF
JbKW9pEMDRvIZVHguosRbb6BZzVH7A4Lvc4FkAeP3bPlVgaj3ombO1UfheiBc7kC
nu3S8kAPWmiu3cw+77wHkjfb6vxpJhG1hzTmrzmR3yxcB1EUKeBpTEmEMrTjo48x
5e9SeDSKik7Nb2RGr8vJvZiirkauSmSJTX9xFCUSjCjmVk4aWkR1/XpP/ezBDY9O
LNhqdlZoEYeXTUJt7fhdkmZhN2WdFKbmv4Fbu6FF3FI66tvQo/NEsXlPFbmxVu6X
xU/Gz76olQCCClJx9gSzjdw8P44/L5AynbkyvvwsmZGKcoBIVak/zUAKEKmhFhIa
7vv/+pnrG5cZ1AN92FvsvtsDbJJjCVEhVFH8z60BQQPEEg9r9YWE/gwbY/c4OYQL
9MfdFziIjOAlZRnLyR4rPg==
`protect END_PROTECTED
