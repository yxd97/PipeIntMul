`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xB+x0bMFfiCHXMHwaWuAdU5VOHEaX12DKN6ZUHsxK0OkvTUesdjwqRnzYlKzxLiS
2/XZ7PE/HgOtFmsA5q7Wf5pwCvvTzv8Q6H+At63sRNx+z5zugsc3GLWel/554LXS
Z9q+O4Y/U8NfI7IRamnRuMjnoQj7Pjh75uN8vsfrwuu8aGIJ/DlgeLHYPnAQ0Tt3
pmBb6jerTwbnaz+hYxH2B+pZGifP+bp+207upKe9aKh8oUd7sI8LH0vFYrvIhICx
2bQYOMj9ve+gvMzQvdm2+2hzHn2kMZVKM1iFM9J8t+WbKideVSCSgqiMECusO3dk
fkrdOhEfDKH5Vm6eWsYX7w==
`protect END_PROTECTED
