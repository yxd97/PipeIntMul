`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y9NQrqkfEJyC0SDS9YWzwg+AG0lL2RI5yJ+SogLEDvN+tkIxSE9K1PzmN15TUK1U
CApuKzDvnw6XLQq5ouw3y6graiBXIRyMNFUXi3P1xRWeMTnPrhG+qmszd+Us6iNw
5NhCcbUPeBpHPd7fABnDSgrGOG3nfMVcVvCicgKotzB3imqQNr99j+7EQ0ApzMAR
iwjmjlR/JDrX39Aiyi0rB2MpbDwJ6mssC6gLlms9cAlJo4B/zfNgHc8fUOs6JndQ
lTCtY3dv9kIw/girfmLmRE9tA7PuoUicEfJogQV0Rje74RhyohChPiAPMxFVCulu
qfrqsXWQRd+NaIHYlgqfCCktWgYtHDEMOwODnnLjnkrKl0E8fxaxJQBfExEGEAh1
un6QeUVk4p3C5H6vJxHIPn0xA35fXrH2ojenFJ8GYwG2PD+IwrIg3eX3LrsJqGp7
9dFqGM5kliAKgMVKeJpflMVPeMooZp8to5mO9Jn+HKQ=
`protect END_PROTECTED
