`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MQNmNpDJS0h49m5gJwrFd7yPhKqXdVwkWftRz47nwjEZOrSk2BRb8s58Kl7LwgH
1ycTbAYGm3A6hhfjyIIVywyaJUHswK0a9jsXmwo4So9xGoy8SEWKN9cKT+Py+Jfk
Of3IpCLhpsC2IQi+5b6OIaKAca4UauYluuMKJ7A8bLVPT208BFVKzCGmkkKOuu9X
azTeFgUQ76sMNHy5FonVbddYyEUmHGvk3X6l+VhZYIQscOv1VG7EiV7rixBBUTFg
XTlQQcC8gQjs0yC9VrLDdBr1lzfkD1SvaAlrqvFJD7TbP44xE75h/i2sCzD6WFRW
MO4TQ0Yw0GCz6i/IOkw0gypSIxbFW3toGf2PewQfYFCjirJjvonNH5JhsNjuxIsU
qxYnzwvTeIk7jovTXE+56EQxmd4VT/PrNh0L/VO4YPg0SGa4LEfVT2H/GJibE7+n
pPG2dEbLtsjzPBkE2r3VldKLnQlUs3FUDQERob9/OdyjCTkutzpulxvX2jMpPlA7
Ac983PV2w7NGTbFn+9DJwxqPvMvJT081bA9WyiwCZfhq+k93OlJhvYgCENR6ptb4
nyqqTCfYPENpZQ1gTROw4rDD/ApvNyTcnM02GVYhLyebVaUPqbgXvz6ZmtQEvIYr
2PvByIuVtI0HMnGIIYHB8fwLjl6IY96LBj9Zhvd4XzSySDwwW87Ehd4LDSDg97Pe
gbmc8iq6mH6v4j75x31RQjywitGtgqNnx67wovcZR/Cu9DyYb3iZo3QkMvcHotvZ
RugkDgGP/8zrTqthFfZsrSCe8nDBWMKfGEDZm6aNvwZ0ZW16/gGlO8jbgn/OIIQ/
i5pp0J622rUFLkBdFL9qYEgk96klklyUFNi7MpqG6vISs2sEsacJy5pE1aC5mh0U
+WQpNtpRJeMkQdfVYKOGORj0LNH/IKXq5fijnUEmqn7ABi6Wub0pEl3EcvQqwtpl
FXr0eFjCI+sXD9pojir9RWudlQvwakvjJOeBfzLdV9oZl2z9L/0tGrjBoqDeZpEJ
4EFmTDKejOkdc7UsZQMcBnXglGqxgVacwWwfUFYfyaeeAYowU1e4f7Ew6dXAq7c6
z4HC2xcceNxPJshcP9LAUtjSnD5EaNeKqe063/9ok9+pDRwm5fNavdxbC5B0hTFb
vzsQHEpmFnak/CpnQOOLxvWEeYTmnnyP0L0/7zv8dvKYis6E/mUDc8ZuYXXj08BV
8nvO7brK7poLWf/XUUJLO96a9sy+WQ4gx1bQtjTC1r57Q57HbGFgnR6TXHy8Miif
Who0nLqRkFWh4vkYFt9ZZsb4z99uVYHTYGIhg0puM5hXtx64tJFOGp4WVJR3DLcT
HjWEr37SulHZuECjD9XS+uRS5aCxthbHMxxBaGbo6dk=
`protect END_PROTECTED
