`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
odfwsgZAj81MoDnobTf9588SX4khSRiE4/i6F53akBaapXBEIXr4Fd0fx6RPMX7I
A6WB3wBrhc+6stDnzaIgCXP1rxb1kyt5/9zffIiH973xu3hl4uSHbi3JAwDSBC/g
yQjNFiS4PBD2zaXQeBBQ5dEjyefCLBxyCFYvEVn1djE=
`protect END_PROTECTED
