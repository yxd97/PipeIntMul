`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JJScetspsMrvHXC64MoY7lCtdtnuzbB3cTy9WYOtdTin9ZBYroMEJxFAvtf+RnD2
kxT8lrx76s5d/nFK0qVw4CcIW5MAELpN2bU+iOeBhOKyV32ExhjE6lejXmJzvAul
qiEz7H1fYaXMvsU0cKi962hgmO/t+y5wftceHZsICskElXQZ4C0QeIXZhWRYfsZB
NTGkndB8OpJAy8PWZrmIxWShPY7nDmXX1Todv4GsvLOOafIKcfT+pNKfU8BKIsfF
prZtz/tiXKOQY4Zami0FlyqE7bydLMPKs+OFPAUCdclvFsPuLYUmmXZnFolZS0E6
ys92Zqw1PlvFbh4FnLZomoU4ykeOjeKPWR2taIjgpKxfmuj7VvDpi9u9Ne+zxWhe
nJzarTkCPpp8S5hTvlUG1dgb/THk4PpiGaVx5OrUs66It+4xW+oCDOmpxG3k46iS
HJojEX2ybJlvloo5RR2Fam71dHSagaEf/PKNRvWWE1b+wfQoNSAVVtLYPBF2rn+A
ACzzh1gjlMjtMVtO7WiQ+NvCy4xhfgw3SFIp9b5kJ/tnKLdV8VESRx7d2OuCYJEZ
Yp7N3mr0Ufc9WUlxQtsxnsd8PpuHD1n8e0y+ZDOGyKodicTpSil5fuy8MKqM4Am6
tK0jXCCQ0s7Q/8kmilUCC/xhrEM9aIVX0zklpcs18p2gscbZedR+bkrWALVDKYTR
BDVO+aWcMb2uAQ+4H6Rb7f7meaBKMEQLhgUvwGZDJOr1oVUyhRFJ/yU9MO5ZYWhd
xP3WFl4GlkTKmMRRF+L+XQr4ztGoKPlkCvnA6CWZPIJ04sY9mDSf4bL1o52m4Ik/
kE3rx2cGUCgfSKbd996tjNvd6/iwWlJjoln1BycKhUG/Gz2s2fJkvLqU5+LX2Mbc
LKgE2BEH/+ouMgOLuIb1Jq1NFbEFjglv9aNn9GFsxtM=
`protect END_PROTECTED
