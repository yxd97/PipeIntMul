`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFMIcepRiq2WRtxBcl2xoHG9JKdTO1MO8JYCJgKkw5e3+kyRlZmpCjcbvwopC/MQ
Jd4kCNpVgSTX++69lE02XweoA8atetERta5fMK/19dTIe3JEC16WKWApvr+tk0v5
XQASOggT/PLzZiTnENjOJZz3+klwbMRzcLfTr36lQHBvByxzqHHrwEVYwvBUEzUR
WbSG/7IEhZM2gKwTdxqSnqbvGv8o3WTN+MTt9zYcBxy1J3mdYE7cZaOxSbziu041
80+gknetaJ0sfOc5K4cV6iMVXNgyQ+dKK5ewixX4922bq29KG0js3Ogiwb8SWbeq
pu/NsrAP7Rof/JVNeUYQPf+MduRjCC3vcScPimsR4UtXnDGAGiyNyujxvHvrywP2
GStE9wJ6HXfucC03WT/2URCAVJ9MtgcE2TXRlxREstEAIfQmzoYvwLZiSXLilJzW
dks2YVKOvuZCYEdsNgptuwAsj5aq79/7TVbTEyCorbx2JnAGD0oRY0E5LHVkeu77
3smbI/XXPn7mF7HsYEKSDYSB0tgd4B0MMY+2oSpq/ZT3erOZ3PXJUyvqcfKU3K77
P/svY73Nz7kKqQqA/I9img==
`protect END_PROTECTED
