`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
icW7F2jN03QX285JEjKSuWIzS5B5TqBDHOe7p/yWJwz1OapKvK+/llU+ajwUoYHu
BZzE3d8ZcxUjQKgACHP9Cr9AZg/yuTswXLTmVPT5BW87naq0SXBpFQThfvvdj8sk
6Z6kv99GJY5wEQmWZIS3dtdGY0JLSGjYzTkvrBVgK4yh3AvtofzZdi8nQScBGKJM
bAqPbN0bxZml0Ag6qe5kUIc7NuJrW9Z+QR7U2NPq0NKd02MmwwrtU+taJSQYm1Td
A2agzvtbqBOn98XXOJauTlJ9ULgiWAKfZKHR9I+xdf+63nrW3jN4Hn943/AcPpAm
sGTxjVwL8vDmzCE2btgiiw==
`protect END_PROTECTED
