`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6zN8evWV4Rl+sqVTQHIvrrNCKxkwJcI0VDMRgsqJt97Y1YuDX742PAyjsCWkbSuV
gQG++aCi1xIjQKtqbc9Pj6zLGxjfl633exAjSKOQBZA0h6S6N1BieONdXgLnRuIE
tlFMRRGXWKW6Z2byVPz2gJSxToS9XeFjHpbgeDZmo1QjBzg/HbOEo1cQEP+8HLWD
BNb/oh7UTccXOcx9F4Dk7JwFtkJVlzjWLfw8l/HcTSDgsdvyqxdQdV6jHNE6RRo2
dgb4FFnPDzX5PwQjTwG11Jf19IMda0K2yEr7JvJw6KALqFTvDvZCXL/iIepThiu7
67jotnmHGy3IW7lu/h3HLZuLQWeMUXIebihBZ+xaoX2rvqfdh/qNEenLL9QtZcoO
nJFHB0aLRIN18+o4UKMgtYfXXyGEptumJHQFm+Y3KnTHBttd0bCzNrio4SeQN523
b7v9jNxgVAZrDVzSODmXeTLK7b2QqPSJl4gLOEziVfdXwXocyWLuFTD3Ue62zZ8k
R6/f6KFA10rOAndd83+wNVvr0szexUlcwFe0reG6C/+Ht+wMXZ7/emqUo/ehUTxs
Ck5ygyplARLCYtM9+35v31MfRmCRunLEmUYGY7MZW0sF3OyHkzSEpYPA7LhvpwB+
5WsVCKwAULkUpZU3smHN7FZOtTEaESZkqgCKtjyJYSEX38fnqsLJV1VdnAby7vho
QTlbdEybivS+sV1EgpkLmPnFSl8ZNo7PNUiMno++unKZQ9b3ACLXGjPbLxR6Q0oI
qd9TCHERRYE+zEkkKjjAkfwn0bDYUA/WHuAj5LMsMo3XFmY3iBvCj8QxzIlayn2R
gOlsYl5+WVVadc8NXLh6OU9fvYpaW65zUCjzVQPcBTzB2iDaCbsSqo68lvcYdWiD
aWa5hh6XpxSi8zXqDCNCwILd5DSWD6DSwCT3cAs15LHl0UReOmhIgVxxZ6A4HXhG
sStt59GdLEf8LnbJ7/SSVXfLvVn0HJE41pf6h7OFQ9ZRmjO0RMeE8HQe/qdOEo/7
iV8pfHIdVOMiAPM+TLConqn2WaqfMXx+S63hbSxY84GbTEM+CF+SaOk1Aw72WLsE
O//d55wF7qzbanIzSexsn+LqBC0cDkM8551cTkzJX53zBZooJazOkISHEqfgkWvw
rOo+s64g+11oMOcjHXg9pwaKNcfHo91FQzygNLv2unzR+AmS4/uVtcOTLG63UhIX
uMri3iEtH6VuLDVYATvLzGakswi7Ccwgd4h6Kq506I5keKUjvMsUWBKVlGImoLvj
DAArl3zmiGwXSV52+0FtNJpjFLy/pR4CpYTMRw4BEfJJL/z+HuxJ13mGwFwSH0uO
tjzSQ3E6/xKuX4xpcgI3zEN6pClttxgKzZVL9yAUx+O6qiY+Mev34ndi0zb4U7tL
Oj+E6zGYkAla+qJmE9HwcMCsKPLVdOZ87sXPydOBSTkmJh7I0xlHlTkvWywvDKa7
OwFGsoKvLoz2+B4znpF7D5KpYk1NOeuxdA667GkHUtnqlBoEBa5x4iYiuiUNjaSZ
UdRr8UkMn0hxlq1dkwyfdH7N2utQb1LDffozlxUE05gryTpcOwiu4TP1+zHoCyhg
19LPL37DxuQCsKDwzgYDi/OWxGuevlNaesX0meEc6h9qCZ+GCYZKyM1RsKC/b6H4
s6MjsqC+j9pa2X2czuDRFeXzh00zd7GSwVuBsWpx6CkmoHlsT+2ciaRg/sn1gp1K
QtpD/v1g6+c6so8SBbplYtIMI+Jr3Ib5sEYwRfVzpfgST4Djgnz51FaJR4HmFDdl
w9xcHx3TP8q9vo/yhWyQqFpPhGT0y92h3lwV7q+OqWzfGthTWvrDDzzijpo2XbnK
KQlw2TKCDWY+zxQV1HH05AhEdpDgfYB17a2NMr8WVzSnzLSRM8XySgR5ycYipsp8
n7uqribZRmKLsZGnhFa8F4m3BJ90ss/bhW0rI+uUNoaLsyuowR13RpJBEKemWJOr
J3idnmf9/s8tZbwGCdgxaqpWnpLtMJL7b6ixq6tnRnLCXkThuOk4ICfrfzhLt7lO
E7o97I1s/bhXRmis9CPATd2tXTTWJnXicn2JZoDhoZTd36xoGZBRwnLlU6pGl6cJ
a3UirfrB8/gccfWB8HQ+zO5Cd6oqCX9/1ZjWOjF95g+ROeB9ozOIBw9kcl6ACh4R
ReXjtTjmK1EmL9ZWwkVCAqY9pvhbMqRYi8dCIF5eMW6sKKvcjtNJjf7aQbtTl6Ej
0bkDRjwyAaxUxFWWzPNKaTSfQaVqdbrG+BbPtUkm9+ncaPJ8WIznqx7tX8hOx5HW
ltAXQM1dkGH12ZQJ+zzx20uDeDYsaSnvNvxasxaoV/n0N/4s0kAQohEe3Qo6AV2P
zX2aAkRogmy0E59vkXZvt/bW/smKVY1+mGSln2xVJ5Zt53xEvJP5OFIjJiMmX6bQ
vAk0K18WAyQPbLdmAcYi725PixGF44XgTIgFOprDKOhjCxpIG9rTLxpFEJoBdJ5W
diymM4hmwaSc1RMc33OMxWu0nPNuWxL5oGzOcR4TuEvqyfU3W63f5PjYaVG0iDpr
GHS1jCUTTqocg3tU2UYH+YfWeeZhoPUifz9YZpNJ/XkYJVwj2EneOmz/kd2E9L+V
+/rkzOCRwOC6Nb3Clh+FFJm/sJqq8vOD/EdomDc1slgyW3RifI0gDwoJ2ygGwCy9
oV08D8KoTKyG0TmsxIKUpxOQqn0cPGwXL52rl/KSvjkFnxOkBFoOhyWSExPdYMSX
FWsju4JoHHqXg1cy8+lcFis8JduQuNgPM5kE/J71kQ0Y89UEv70U7GfUVrSBEXcQ
3oUJlGjewtfbIDKtpjmGXAA1etvUaz90ucxQ33fX/HePdlE+nAT8jR3DVY5QsM9V
mhxZbrJvHLz9m3rDZ9kr3uDBDQ4niIiD2W/eQDPlILY28teD7KixrpXakOCDL9xP
bfHgZ33u2DOo0remV1KpUlklGZ4xo726IXiLpqarCTz2IHcACZvJi7baQmOsE5jN
/jEqUvN7s5HY8YckXrYon8oZPcRtBmC2ziCqMiR7D+F0pE7v0Gfg6OkY2fHYM04C
qpkfEDiPF/vZWlkIXmVVM7Q3ljXHqPO4qnTO8pRD2Dztyv01H6bNzG2PqRpCW51o
vRF3KtJ0pTrdX6JC5MbFVjFyIiFYmvjSTjb3Zwn1TR9FE9+9/onxEcQbc+cqXsv+
KW4umDK9qDoyBeFranB2XCVWmZdAN9hz+YggBxYWyM1S3ZOLCFABN1p5MBpwO12f
ovW0bUV6Z4OR1aZhYIZaLLAxZCBE1u2cXMXVWGz+ZgybVMogVUPKv2DLPTradFRt
OwpQE9TQh2kZVK4aQpDh3YNi+oWgJMkWh5vGD8NgV7GLCL71NIvBUnxvlkYhJRQF
rLng3+GnSmWc6qm5BPXgN9VlnLJ1rvffYEhHM1f5JmqE6JYLPB5FK/+VUNWS6SaU
i41AF7NEKmC/k5n5InBamMzpBXCEB1pgiUx+FCcbUzfQt5ccS/rFmXU8oRBbR/xZ
IOXVi25/F8C6KuFxaD7uE1RydDE0l0FvFfol3UzZjat8My3JvLmFW6pcMt9cyf+L
SeVU3o6lB8KA6N4x3icryKUOU2kXfOnCZ0zIATlX8inaasj+FaNsULr7oAC1drZS
NEhdoasdJOolnwWzlveHwP6BFKYpgujQLSM/aTuFhPCfR+Tg+NriXCOAgtBwNMQU
vc7gmbQfVS+gWuEAP08zuVggeaYU2aklWWeFJgZnr/udUR/9fB+bk4B2No0jFst7
SGpmlLoycRXdDZiWe20JRw+z56e6jXjMPIeK6e0Le/+iogs5QVEfo/gOe0URvKsH
FHw/f6BR/OcK1afDsRVZy5IMDVfb1tPgh1UKjLV8ai7aVtLGLLsSVYVgebZIawco
oDQMxDVa2HIIdAQL13B9jptx/T2i6zSdEw+j/MoejfEggq1FZrNhZJa6HaAFenoF
T0pH3izqTzIQitH1EaWbzZZ0SMT+OZyZr7d4ZIBGEcgS+Acurf6E7HbneMUcYgg3
M8XytLn5QZkY7WstZMkY869xZ7PB3fWlyRkTl2odv4T1pojcamzz5Yd2cV95Fg42
wg3qeAKV/uZYQz6g2UpHGMM0sEKmfRs9BbPxItCsgW2XFHRMRZ+La7dwT9waW2hs
NnqkwYtzr8bvmOB1LPyUN0BFffkjYyLNCj37dT+5cNl3tJ91NiMAkXTZdoDanK/Q
6VQAXIdRMaVpVbeY716Q6le7RYTFfl3NEvIZB0x33dSFDqzjNX0J+HXsKi7n3bPq
D8n4ZMRl4MYmtoBkB4XUAst8kiqtJ4t23KBSabdCVf8+NHz06BYTwQkrQUPBo78J
ZPNKdXXybHu5xjRDKUzMRDvPSYREB6IKMALj9S/pYnRy8Q4ntek8n1v4mKHIWJf6
ui3daVouK1hcv+FCBiCpXICNapSjsGilFaCXwJFvF6U7nsI6DTDBinXrDlO0dK+J
TUkn+Po9SW20DgBAxNY4GIXNlPb5hZVSQAwuKvsU+beqs0uxOtDrm9H3EoeX94io
M0OXkklDYWO5cjAspA2WparaW1ljaNCmDakSiXi8/ez5GOPIfeKAVQg00Nc9VNy4
6vvjXRafUVDgowdY/kaPyCXaG9z+tb0StyA7+hg+ZpLfCEUUZKxJqClPJIIVgAfo
cMx5e7HQS2du2kL8IK4glqoUY+6uX5b0uEYMfS6/n4+mnt78BVoZj4gBX45/7S++
wlEIino7zwJgqYDLdc30n3sntWBS2FNW/oFM//8Eh2VPWwUdJxq0loc63raEptp1
xuFdcW5FPB+/PZrzRrsJ5tnI+jCtXZGYVo6XIyJIH1rb5gQYkmvYTfxa5900jtqA
yxJyIvvcJAecWTu7e4Bvsi+3W36uJnLuny3i5HFTHk4VtRmJqfLo0olne3f9Tbow
s8elmNUwPaCYWppX3+P7b6b8ySDtuCAQ94om5y80DuUnO6QplLpHMPFMwUNcxHQe
GVMS4neWzWLCjdS7e23NinD8k3TpKnoFdLHt9Ah7n1kxR6D477ObrUbMazX41WNz
YsNhVBaC7BESQfaUizu55MhvYU1AwbrVVPWIbpyrS89sTqXLiGbCnBueSj5XCAb1
VD35E38n7TU641VH2tSaPxQZdynyEcblw6cdHLR5YpsOTZb9N6j8yhgupRbcYc1T
Bv1uxdIPu002BvRGGk2Og7Z5o1VyfcqXuLGCP1nT3DCL09XMEnPqSUb5ubJYP8Px
60rdILGI/otT0PEk+L926SwWdJV2Zyy07j8qh9rV7w4CUbcxeZTG3tt8LEqD63N9
HASP1F93qDJuMEi924E8jJvMmqffaUHMwLQ1np7TqEPLMtcw6qeAEeoNIKsnO8kf
S0VNptqM4Wlp5gZc5efWllhHw6oIrE3Zg+9/u53AOxPH0siaNFUucVKKpi6Mez80
LNgADveVqYopDCGCYkVj8YT7HuI5xczPZj1uGvooYWnMkj93YOUCfPSNKnYoXEF2
ejxv84Al0bI2S8S5KM4bl+Dy/fIQp25JPJ1zxp9KXzkJaIC+VNEHjUpnE4PCTT2X
pcL+1rqULv9enS3efN9jedSRJAkcxucedUQ3fbjvjsRX7KAff1O0ctE5I5ITP+us
C5HgMJOnSa9Kv6pmPP/ghqQS8HpU1WWvmY1npQOwIJa/ywnSOmKVmKm06Ecz6Vyy
ZHbNuVqMjI37p5CV93T/D4I8JnnQEQTRX0IGhWqcXmWeDWAQcd6dmkkAFC+bv8iP
vUR3d2FPEsTQ3KOOsVj84xbGetV33PuA+ark8dFWboateKnxEZOD8eoXTdQ3xyGC
ycBU8efpDLd4zShd+ODD7HhFfdoYgzsk4DuwP0+bdVAROPLSAQPreFCjLjDrX/Wg
0NnqVssruHSXn/p8feTu230/Bfpw8xhuNmfSf5R92JwFCb7he4dfPvrrLzWpzdbm
gjWzMSROPARQDfegPJsETuSKgO8RxGndXtpkPxRHdAeW5ooXUgQlqKPlc26dM9nK
EemX6cFaFmuNjoNGkagB8ZZL5JZIjPahn4M9RNShHGW1jklG+SaKFXtLRmrPPQA+
HZP/CpuLRQiR6F8fugQVhsZjTQKQSodqoOpFRuDW5YYCoR7fX2FdpPBgMLA7oinL
qrqupFjDCeZAmlMp5zLnkD3X6yDNUqSIXAfqwteSyBcrcaoVngvI5dJyGMbmb05P
y+8MRSRvZMcqR5+0ZTaq4LF4/BCp3paVO6GhGQB5yTeEE/uoNOLPf/5Luddh4Yii
lVyPIpv2bOhUpHb/y4ZqFXS7I5+8QUTmVEB8BkJgLhqOQ2Yy3ZvG643b+V9U+8Z/
GX7qIkrEThx9AlIfnjHw2TZpIcG1LG++oeQTw+DCV+VU6aMzqEvI8IUm6+jjGDog
wpHn4DRqNc6VjpvQUjen4h5a/Op2q49LKRELiijHaFMTBaY+hJsqeK1ETiJLIaaL
KOa+/KR81rVeWQog2dVupwb4Ftjhq6wXBxoK3tWGzb+hl4V/FfiCKyrTMfbPZvVe
Z17zG+kvMM1GhLmwDSd9NwJ1WbH/bdinn+vV+fZWjR/5D9Ls8zDX2mEBkvdn6yZ+
pk345Yl5labompDHdQ4j+abCGJosTMbLI7Hf1o+dhsfkmbJ295d/Kr/aenn28UsP
G00mOBg2mtmsBFYWK9xYle60f3P9vzROMANkhxcLFufthw+XxhIawCIf8lci7gnB
o9+tISQ4KPWrWyCwWun8oLRgsgjLO1D7s2ZeLVOMFrRitzd6Z6isbEMy1s1jM6oH
uYETcsrLn6h5Xq8w6HE+xnlSKFRsuj+9m9Kz/ss8e4xEUDnYYoGnuJdb2UnEMtU+
0W/5DVg+FdG7AvDAyYa4sCwcF205nPAGpscXx66loxnVMuL6YqxYOiv9xcJ0SUV0
7iIwCJoa8ooRsI55Hurce6uNu9bq8QDq/D52WScuTtmRChDc/dlhTeYqTyKsm/Vv
DI5RG89fxk4t8tB61D3lQ5kh4E6jOAr2iSCwvGGnocTlAJDecLQAtDJAzgm1ctLg
jABUOqJ8hhd4Iv3X6FrSMij5GNW4dI84CAZsrJGn4puV/KQ47ofLfTt2PRHUyOaI
t/tE4MlR3LoCwoRB7G/1EbpLljlzCSB710uGlvL4ca+HzeGJ48ywKYF66TcxBPhh
eL1hOEgiWzZ9gzuOBamVXrZOURPEw8qtzPlG+HEkecbdna1vdJDIRiSYV04gSCTT
koAIgmhIV2nEtgJppN/Vns4O5acl+CXfT4xNzbl4aDXBvEJzcJYVdFx3J3yiib5o
WZkOt06XuobkKsjqR6A8fcuymOoKdfdd/EZoqtmkYG7FdYaCJKTnUR0/EANzFDr+
CXeDSoSwEDjl0EkX2ogJW9O6Av75++R6uUgYcIhThDI82pgS5NtE2j67md+A5ZhF
kl0QKFJ2oCyWY0rLHoEDuKAbpz8NNXh3F/7cnPD0NnLiZFe7yqu39/meWmIdQo47
54Dn8nnFf5HWREu1zIPLuuT7fJ6Ad6fogRiOk7A+EPkycoBNsQcoUO0ajnoyJEsx
tW4JB7HbqfSo+4XGCd78d0RoHxdOlv2aUZtXGRUe6eBK89SkjHAMsb8PJR/6U2ou
W9Grb1iXI7p4HDKzUuW2eGxFZJYUfx7BT+lmyXrkp67orMKOFFsb/Q9H6EUFxnAq
VjRbUD6n9B4I0JCE2JS5SWfJ0hIEYXHGZqt2ETuCqEfDf1vx7Fj2PLJmxO2QIyPS
z96GRX2PUCK8h2sSFak8zk2qAYg3Vf8ZC1vsh2YnLQ5IRVoH8KQ319WVY1CuJzX/
K90200I4hnJz+snlWvGbFLVNy2donrgpC3VVujGZLIdNTuIrdLGCo5TK3fZNYuFs
qvg03tghKZ7HWwcK8mfvkfuIdf89YMcgwDrZRVcmKkd34eDbkP2KHSlXm50IK352
p3GLtQgyVJqM5HFqjuilqCOFW6BJuOwheU/QRwh/Y18eMCvKaCeoqljxq5RHHWmz
RpNnc/NYLetTuZb6FeC+WQN8V2U9Z9ywQiQkxrMjBSwDRJdKmWkuWuaHWw1i+jJ/
ClOuHM/7QldXLboBPnBHaoBEQLek3UDN2PMNuiz5fEHew7VLtCmXOk9gNmN5Y34b
9XocF9pHLth7TAm89+hSJ6Y1CxliCWkfMEMenDlPzynl69Ibx07GsB98n8j0YPRo
xCmwXaEAeCIjiUaGL4kXD8aeobUKB1QaCd73wdMwi4Vn9LLG/FpL56h6W1TP4cr2
ChuZegtfSP1CE8M2jP+3Z5QBLNAZtwFZeQ1YYPVte2Vm74MWlIxz5SwiDsEuMfgN
RCW66Lm092+MMQX/5NsqDm/yQUWFbXPlfliJG3xLkAInoSdJt4fTUesjcwZicuel
oX9+6fFZCFRm1yzZAncsogPV67jzl0Q2h48DX32C92SyfNyqyDojrKujwNv6M6l5
a/I+FBofMBwwtBAFFr5wMDrlsWfsCYlI5gsTDks+NfV8slwp/K9oEukwqdFlQ3UL
TmjLeYneGJuOF6wKN5rZkk9uvrwd4njAOjKYcI4uerOKeO9LZHF7XAcLko68rJ0u
oiohvLff0Ss75UgbeMI3vq7JSf2PW3xS3E0X5BDTCWNONlJJsGMqf4FRqRjmvWOL
jWzExW2uI2gUwX2QEMt8NR7aPGVJ9g1/fQmnC0tVxGPK59lz9etouaTYd2hAlFYL
4S+XsciHa/QqwoqPABGH4igr2TlsDbeviVnbEwKej835P/sCBGwCu6kOWtPUTluz
74ICdk1CiPsHbjHEsy+/qzz/S56yuZ0iBbydoYsmcngMzJB3Uuaseg+AMptf6stV
EAibYhyhb1AUnZSTWJDubp+RXK7VfK7esIVtgssn3GRX2xZeRzW8UmDLUmebCKWO
TJ2zw2dYUtMHY31Xwgk58LwZEZCBnmuEU+JgRqY3c03BTFAmpFkLEefTqaZDpRBE
kjU1alj3Kpyo0oM4Wz2GDMuexpDN4nVLzrqjV2uN0AKr8A03VLcH8wgZLritknXX
Di6Z/6H72rxEMTK/dcDagDZB7XXYNvPqLivsxv7mD9sJM8cocJ5FM7MLAypXa9s4
hn2lrh7J9ESHO9QHTusFzRKwtBh6TN6Y8VRh0g+kIlbNEkK9AFx3EMCDkynU8/V0
DhyahJHE8pnVHTJDGWYT7Ss4U3MnsSH7RaFJx0MPB1aEEegh2DMQOrG5+b1YCNAQ
fZ0GvAYugZnlgnl3i5o1M3VS/Qc+7+/ZLD/NHSRSwDS4ARhoNugT7i+wMSEk4VeL
Gm+kotV6Bvs/HU/ZmcGUngytT18FDyqjXEyFqo3fjK1Wt+42Xgy3yKZUdqhhogHt
WBYfWr29n9fkmqMBWspInQafMAsz0n2thtNe6AfW4kNOOVlxCM7LMF177O3nJkri
uezgrSYtCAIh9DqIhRU+aMl2wld0P/1wWiYE61PYcw6BjGr9lK0DHg2LDjlif5Rh
xygLHocys2ZcUPSTlg8UWnMfAmJZA1c/dZNm4nVJRNHE9ohJF3QH5ZaFxe86QlMY
OcriFUiio3x+MTXi+Rh9MGI+q2UGY37zdOah/NsV1zBnAa6rKndrxtlFYJnffC5X
bKqC7GyFQSsTsLX76chJbtkTDaBhtomQCZG80KPsff9UqWqDSuGZ4lzoq9LBY7OU
AkCShkaBtbsnhML7vCBki1dsaF8ZJ5w9XRMnY5pqoCt4wi7HOg4Z0O9D3ivXPCFb
8ww4Xcaf4SMuWIgQlmqGm3D7EvOX/K0f8cNrNuGZ42yiJtMZ7ifoGJzgk7GlURAa
4PjUwFXEBUjbCvy82SgGmCRe8y+cLOVlnCn1iLd6P9VNFmD2LGslNRIIMKwsboXi
+7HUDGFNxM/bSe2U+7/2CA6EPpXbGZss7Y1p6kQce80J/nJzA6QwKl23UtEpw/94
fwPtK04Wk9C6o243jP+vua11xsMhvsCTgk6FPXEGane9whIwq/Icv5d7vGtxMZ8l
A6d2YnOnk02fNppl+nU3AJP85jekjgrDX1x/C8WuBaAF0PN7R1bwGOO/UWpczX+y
+C03slVEC1+43w5QCWrXprBv11WMfQA8hmzS+p+vS/z1VfEOnrwZhgEJ4bL0AsN9
2aFp8aYg+hTwbRSWF7fXltu3t/kIOym0l3PcZeVFWqsBmxRzYc4cflUkjwT/qm0Z
V+abs+C4IeBu3ejITYODrlO1vKUEAG9KtRs7LXT3yBIEt6hKXYZMRcWwqwD2KUY+
RMnMPylpaRnpRMwPQyMRX/rWObiwPifktz1u2fiDvPQ558c9anHYscXH8E2Rthgf
F3jfJDFInq+h0YHg0/5bu6OW380QxmZBZ67OPKBtO6rTJUK1PbpEDsbI/qj4iGRb
TRWRf18ywN9VWQmEy0M/M6QxZZh4ThcjqC7kO5GqGyXEK+Y9RB7AXjsIOgEvd5fe
7iswgzYup99zdoKUYieYT0V8O8rwNAZ8CiW9Ccpz0KMNqihWlNIHeT9iv42Hv/TD
M7jN0UybgkOcTEeulN3DsBqFwzKyysvYfR0EScOzUgmjI86eufJ1t1JVFG38wrUV
aGpCidG1oUZLfcYQPqkA13eASvqeStycQIUc+g6efYbJ/a5jXwwVJso2VbRCw3hK
Hrsuar+UInLExqUMwEHkwEdWtC/2HCLkU24WZip7jDg2ffJB4CQC/GhWCGeBrDLW
PFo6tLEbCWcGgIWeAYLV6DA7aeOo7zbVn2jLVZoMeiVKdZqAnBmFHaiPvum8qJzp
omS3VydeNaIWrMfNZ5+FnG6XXgAy7TXuMtVCjogy6V2UVfepak95hEk3z0gTwuGn
Y1B1LjItaAvQucr4bZzqQWAXxb3Xq45znESHIsF7lVpZ+6wsRTnpXWtv3KIiCjLP
2AmU6pBJLj1cVTbWzn7HS/yjI92LJ8fDdki38u6dyhCM/8+oGCWCaXaxndlpshZY
WIqrfp8HjhXLBnJ25J9UGsE+NVJn8ya0fV8MhZlKx55iwhDrf04WW5efKUUHg1re
hvEebLjMSHaEV7cgLQzXp6SNzZaCQodzx0L4R6BEWNXBWLrm9dPKG4vhmeIg7nYY
Me1/sMhPpA8WdOXVrYHu2QxmO5CifaWIF3+njaT/Sic15S3skzRf3RWbceAGFjxv
0UYbc6UCrBDFWHVCFQU1KppObykSWV+9gIrhDeeKiImBHeTCxPrb79m8KXoKGjcN
4TsQ5D8EwhhAzXcpGnaVaQ23voz7gnIwuzyrCm1EqSuQKJui3+YqkxQPa58DDo4C
xASjktKuqo0bjWa7Io4mE7BuuS+tkmYrpqk77HOZAlYrAUmMzoBvE9zu6jvJV6na
0DMdlW6dyHGEnyLpiASs+7rLT+5WdVd024u5A4PV9ozb2Sw1IOIsi7OlwlyL/olr
7L6C7rmTn1Xi3PahGKgBetctJJ6viZlXhImHWt5lUkEMKJQ2ehB0YtbGLmo1ZVPB
fJMOonrbteU8f5BpWMxnT+IH8GhWGJZrud0NX/ssi/U6Id/uarGHu+TITqn6dzuS
xrsiySnfcADKp/mZoXV1kudrkBVNcmEOr+oYHy/PV2DTKUtb+WIkds/7RS+tpDID
9GPkblnD/dfupmq5mtCodOd3GX2Mn00RLKplSQRQCs3mrwwQ64YxXFlaTQXYuaZo
Ry3rkDeqT01nTiZa5kbNkUlvjCbEbp+6YQqvBRentAKZaPkX7HtFj9ipBu22aHvC
sXnFab2KgY7FT5XiECTUfv7LkqJGe1U9PJwB5rzTeXuuljK2/pc3iiOLC2qLoWKs
US8c7iYH/LfUPmst2b2Qt1DHkcGUILNyG3e5yBDHCnvJom0sRv8T4fkLC1PRJZ9C
XnE9W4323IIFKHIKL4hMqX4qVboZbyKEPQzbXQLh5jzSmiDev0glG+Kr5wBaA4VZ
EPbNxX/LOWMHr2vJBF60rDQZcESN3ksMtAel9L158dz0GMpCF6dsKugO86VRLhfX
YGg/52+ibF8gszxX8QEz/UvrvQ0Q4F/qfJ/T84g0VKHfQ+D0Rm+FICOq/gBTWL39
HBybM7vr6XKeRq0o8yGJ85L+prNmSUbMF/ddG+mVrYpYQSn3w2GllsswhuuUpFI7
JmHiT0bD15Z7p8qOZIwv8XpyqBt743LVFb5OFxTC7FVyxE0AuqDxIhjz1alp7gu1
xiJwZkS0/OWyzYO6+hoLyYCFhXoy2wSplX0pQBetVFbueRHS098AAkCDMwuyK7yB
W+/cJDv7c1ny0MULLTvUa8G4mnB02y2Iw4XsTriyw1W5BcyY7mwjrl081ZzF9Ua3
`protect END_PROTECTED
