`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nc+9Vv6MKtOrNxdLxwsAH+/qrDuf2Ym+zBZHYy3zVjSr4XHrcCoYRuWBXd0brXSA
RwFjIA8Is/p0osC/r4vybFtTkPFuy09tNAooFB9YTxNDbcDxhOG/+YJrds1GoS1F
5IdRLkm/tFiGEsteZaukUxtF09Q94N8mpB6/TDo53mCoXyxO4jCmftNJjh0HTY7Z
E9uT7qv/J6vQTyMdO69e3kSgSrzvzR2CPEZUnHELLY/iCjerMgxT61tOY1j5MpJJ
vpl8qOGjsCGBNKviEvY7WtnCeFQp3JTBjkfit4QYvnky8RAU4xKhldKieIddXaDN
OgmneSCARrVQ3FthZVaIjMNXYHOFyP8yoT71VA8ElpmACCQFo/wl3PAgV8rwbPxj
GL5PDr2tLXve7SwIHwc9N3K0MbquCL98CaQ+yizfbtHzHnlPiU+R6AOUFwZty1O7
UHBIG3VCiFrrO31S16p6W9cpa+jPtEvYAXuRDmwJtGHgj84Ek2fmt9pbI4fv+wbn
`protect END_PROTECTED
