`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J664pcgyJwsSfip93Z6hvuTj8WAlligMSNCyT2L8fs6Z3JxQErnnLYrUPG386390
MjMtWf+uMHhYmvg6RHSTXmI+EoSR72bOh3i3qp6mHFyCJb/u+fZ2ePKCuR7V8Xq5
AmstFBNnB1/RE4xHNcEpoS8Tiiu/J2mTAtzeuVQandQZAXnOpVj7Ftjxg5UrzY8V
xs1X5/u0R46keBRYCSM1979LZvoh1w+2YrW4DCZ2+omM2bJE97oKeJKfcn3c5WGq
PUredDwNx55bWFAoxzh7nbT4t278h+SFFM26TGmN9KXYomCvM/MgKBmETou+9QuW
5OgTdjGVRfdLho/i9PAsu03y4AGST1PhuL/5uKZsZZwBlWAx0zulifl7jfdO0UME
zP84bnjlGopy7x7zx10BLZmzu5N6mbUkkH/3c1PePCo09CrE/mEOflMiWHTMZFq8
`protect END_PROTECTED
