`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNEcU9j0IJch815XauSK75ly2E97ZAZkfLr+zokJp39vf5Lvg+iCzreSuVZJxuHP
53VwJKxeoSy+R3/7YqU/nYGF6Fg+QUlRAE54JyydKfSjPCLHT6Gt3jmY5Z7acqL5
vfyUAHjJR9lnqCKfJbX5arp6nZz95+E2d+MYpbZkE8Casn4GIng/jn2QutyEyf7P
OawKsgEYJF+UKavKSq0Tn2GXsPKuojhmFmZyvvWrJODpSD+W84MNy35U4kiodeoQ
tD9QbV270fZ3HhZvGRaFQFjQOnqgDJ3beNUh9qZozpaYaMmzlhKjpn4rAtcODfqx
8m73VSQq3cv+w1karX9yhRhw4GTht/zREOIEu9ExzX1ok0ue+6qpVNqaKbemafns
LSrAr+9u20g0Nao5A7xPvP3mYzIPu6EfL38g593Z3TD4ab+qWUgIc9QjvibuoYHu
Qxaa6HT+zd8nfECI9Etk6Q0V3zxseCIt5pKaSlXpkbvfjhSDj6fr8dpODM5qCVRH
2NaWB4hzK9irNyh75ix1PDJciJnSsywCZv5NIckG/iGTc+rSe1Ssxl+TPP6U6t0b
xy6cJpGzoPKzKkyJlcpbPEmFd4px0ux5JeRVdJ+qQidoCOxLKsUj0Uli+YVOvaNM
OA0HZIQz3oCO/8dm9IaMFd+WR1gtzquERTSUMfRArAS9eo96YhlnPv7w7Gsa3a7b
qIkQx+RhwUDxHNgcxtdecoJrzimvZ4hV56hQVTTg62btabVlljMZTLJMH99sM7o4
Edhoo7/zRoGtaLdPKqYuPC/5RNxRvo/ebgPrYaiEEdFjFRRZkmTOqhGKPGqqE2q4
q78i2PfecbVuIBtHV/Jdrw==
`protect END_PROTECTED
