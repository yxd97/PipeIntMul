`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2fIHnq5FjPxZTfzDJWBwOYRPJ8lDaPYtmhQx0eC4XGbyekU1+K+PnoLaQT8naYk
NzLSkwtoq+aDfTnJgz2yg1oAQfn4Sg/jlSlGc99k/y0Esh7glQVPskrMacS16EC8
I+MZXLd5QllMOIEXXPtcEHKML4bAOb3kOTjxwr+ui31DLfE3caBFVw3i5I2N8yW2
AVOThSCQrK+8pSqUGL3OlEmexm288IJIUwVg2xFbqt5pFK2PI9cGtV7pw1jLO860
5SJFUnIuYQWiReCtkbNQLQ==
`protect END_PROTECTED
