`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BoBiYcwSiUfKoo5f0kClZym4p/3aT1pVgwXU4hbpLBe3PnG27a5sAd7X+z5GfZLb
4DaJuzd4WnI9vYqVUnQlVnxjbKpvxbedsq4st2ISrAblyse6sT0vWQaxfG3taB/N
Fl2W/8AX2fdogmL46tDRuUl6UtsmrysvfqdNuCDi7Yi+C6SdDO4L3pxBAGKIHQ/A
zbLI0tWCXwR5F3IrCgxKYd5pMcojymxHRWGVvu8nrY/sDFtpR6jg7DLFh4uyYcLY
0uGhMJQbxpmBXA2t59cRNIrd1A072+yJk8ArI/mlrWAmAZOhhTqCgfOf1nR8RA69
8gkn3UoIvCIOwk0iH0h9abWNErxR5k03uaqGqfORgGiHzeKA4UykaBtVxUpWhgyR
o6hLxTYckmdOtnw807MZrvQvMiQH3OjuedZ8Tx14UKsh7ci5/+KxRyJ/6GfHPDRS
yvpulceEnRKfkrAblvlv6H9lxUNun7KRlN8haQpjnjQeP5hmscI3gQKz7245+C6B
AaaV8UIZYh3y1fL1l6pK3LPllzhA2p0ouovs+5DUf37G9/1ZVJle/BTPb1EkUunV
3SRAQn096UPLx+tH/WCtw0YXTSM35Dy/HkzfxQ7huUQ1iyecurco7h0WM2abGvN0
`protect END_PROTECTED
