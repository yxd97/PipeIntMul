`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qV4cwm5Fd4x/JioUbI++4SYylaTUTh8MvqBW8/WxW+6ujcScPPSMRxJjHDnUbotm
ZVoPAqJOT1gW46EODOLZQDI/U8flN7G+cbl1FaGj0LUSL8qrpawBQE7KSB59R2X+
OwZPqp3txzYIbV+6/sQfatCzPsVpnrvpT0njambqRT3Skan0K43lmtyxbhTdAEFH
QByUoyJcKIh0ZcrNL7Y09qBZfNKGYw5e0Tdgf3Syw5hHrTAaJXX7ojiyUKnGy8jk
`protect END_PROTECTED
