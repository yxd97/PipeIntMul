`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qG5UDMtpz6PfKJaduWFO7ubqtz0TadMqA/5gbxhE2hWaZ0FQqHNpSjlCw3McXq5o
1QTJ/VnCXaYTD6/eeziv8JuZ6eW3nUmML4f/eKGN2kNXLqSpCJ7bGmyofIBWibri
6NRKK35ac3O6Yf89rnorM5IEUm9RgJwMaMvkLmkhS+cyt3LuD5HfQBs0NoQZ0f/w
xNeydh+4qjJiv9lz8tAuHY7dC/MwBFOsL8ak9FEt2LHWuPdbyBlrJZ74pY4nOa6E
Me7HHkmO6uovoxSm2w/w9ud2kj7PfK7vSVqO8p0nAFlLFmpKaIV6ikrfDDp2Crj1
odTDcMI56S9NnreAiG38kj1zhKaTdzNpl9O/Hn5IBsiSN0m/9BzdS+LeEbpzyAAz
PUC1PTPzicoV60/pXDIngKIJ1x5Il77lVugVGB2c1JyaOuEe4++DowxRPoF/c4YF
zrQv94jqdfY+faQCpf9nc6LXDJwoQ/wGLdk9pS6WDNY=
`protect END_PROTECTED
