`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
skZo3koXqh/aPvJH6NLHh7vSZaakTtM1/F9Kh0trVm8kKjYpBcgyOHBGxIR1B/h+
hMh3ex/yN56QFTym1VhfiNn4ZlbPYe2M+SgitPhwZuNZmN3Yiljb+jOSDuLUQmSc
O8BdTzOtT9fj4blqRqF3TSaE1LbrLNxbdULaRWoB5Bn0Ffu46p2LkU1ZGIaGNPtx
7Hau9pQvCqad3L7OmVU3oXXTkVGcu4r1lIuxAQd4MVtQLnS4i0eEHX2NNCYR0GKN
7hMpi5phnyYMHaQUO2Ml3oMQ0lfmMV0M0l3x39xZorOTOLGrOdPU8ktD1Crc1LL2
frcWDbP8GtwRmnl0N1diJ5IQz+nMdbnasznRW+PUVxb7dk361Zuc6BT2FnIIn0vq
hmJH1mq3wZjaY4vab5MZMPulLI0kOLW2I0pMsQvPvEghhoVEvvDeK3rCnWUy5NGX
bmxlbYXxnCHyf3wnEHceZx6YpcRjmql2CiJLLsxd20c9l2U7viMSMzZq7xfs7wCI
sX/vwwDDJBt+DD4D+KXukMeI0wxCjb73uAtBcoQBqml0KnAUyRBPvxeE+7inDQ+L
6putDj2r/iCrUw2ysJjE9+AVf7Jcl10N9rZhcKkrfXlgaNEieL46jjwyRmkkBLVd
VBJj79YObry8yQt4SvOVpMNWvqCNaNu4Zp4bbPxmJioTHxdTTkuZ8UDhlewNQSdi
6d11Y+N8a/t+idrBuPWHKOBu6QVmiOt1yQi43Uh0SnIVwa58QGN7kkjeM1YA3IRo
JL9SgCx1q9XjdWCVJNAf/v/XVVqQUwHFMFNN9HR7ITP9sNoEXNWu+UPRH2oDPWlT
ifgl0S2Ub4dLnb0OjWtTnhRbyx2vDZAlLA1/Nk2Pbf8N0XrivfSvbnNoTBFzMVUw
lIfSNUkwCrSsPOCLzB1qE6L9HioVIeJGkKaYOF3bWFWKRH9pRwnP7/FAe/a5aHF+
ZONRKRfL82ngzUNX/wevqg2v2uPNkMXFrsXdDaKPZkFG5yhJziGuBb5AQXCyvNCn
x3PrC7PVr4kBuHjTtQe32C6P6qAORn4EzHfa3g6feVidY1OE18jAQw6bgQgB1XuJ
FJdxfk8XuR9VKY6/uQjgSpoSb1sR0oABK9Zx1zqDQVSMJOOabIeKQ206eHwbfGHk
tsAIiL0GLOqTuOF8DEzxdJEA5PrRHXdmIuEvMMti421JDCU4tbSKz+jWWvtrdeSn
7OAcd9cze5DaM+fBSCiwbm7eDbCbAFv3zpa7LE/pj4bxZDBL08msmLvyt9fBkezQ
Gf4sY7hi1k3ARe9DpzzCXpJtSt2hdqMnUeEy7eX2oyFDUhhHfxc7ktJZNCsyXAHv
Z/NWKy9/JqPBShsroV3Z9AlfcXEFuAXCdD3mNdyYtnUKgALzzo4phDb3XVhyLAFd
AjdEsq5c29GflI9a2Sl/l8zf9N2Xt6J05dHpbeY6U4EnJHdmFJ06fw1J8khT0nHz
F2rDWqMPVgTaZYRwxXo/jtNDHFhatvLOU1x/jQe5N/xf6g774NiXqC2cYGIubirG
g7+5zAbrr5lsdY2+BlkmbB3+9NrEY+qFxVZaqyMAWsXPllxS2cBj4OUAp1N5E46s
FKcww4zR79f+rAb721/s4VdrOXXKLZI032FROoYj9XuyfC/GRl7U2DkUj4aVOSyk
own0tCGtz0jIeh98+cXicftBQyR8vMX4h04psMnnCYdnCO32VUm6Q1dihH4ksDdu
7r4FbVdAi8pf3eFLwHA67DYbhf7oqO4EeZk4gU/hG1VFrlJGrN0RXCKRJbub7sVi
DRaMbxQ4XoceoIKyN2nCuwd+st5uCmRfigoAZdkKt9SAUNv3HbqA9L3evuwzOPs6
hfiX71cIMM7KETGTZdnEnuYuXAVTPtJDz2Bt1pr5oJq254BxT8p9kxGwXDzqCKFd
ooI8MkDV16hSryWai31ZZusZLGKQSS61VlbMrMlvNH7ihR7I2TPWG2aooxssTmGr
IEw0u7bu/0RsePJmu5Avt2sEaG41e8YN0UhvvDeTAlhpNWP9EVaIEgkxoPj1XUrj
xP7Pr46MbYhr6J4lD6EV0FVL0Lsi2mIwn/7BDNn24CBHq0gpMI39XhbYVDHMjtkq
R9DZUQizHVoKG8sZ8axt3V0jUnvp1oXaMQ36oD45RTXU+wkkYFscX3Ki9XyTzDOA
WPSPoFpbVb8kM/NvJbbTaItY3HvUZAX89z/dfRxCq4sMwEAIKKXnDBUNiSY20Ryo
BBO0JBxpmmC9VhR6kmnhGRh5RFHWJaEE18N5/2gxa70VTTvkzZAKQWSiRkAFhoKn
fWgxX8srgfHGp1S1m+kM6N5A9l9ouYiov5WHMavWwxdIhPzg+LFmI0+arBgmAXAt
inWupoT+E7gUPbKlAlkGIkmC9+OsrNKHIbyxSAwSyNhW5opf+2oT7frdO0out9oD
Acd88FtdBA1zFprkASR8GBpRKuhQmxkip705mg3MQ+prJ+NHUXEy09dstuoFtX2b
CaCADjoWZM+BoNhIHvFoSgLgIap1L+ChGVMYLuUe9AyJDNOaoTIqpIjpAgang1wX
jg7Un2W6zj0zIGglv/AeCVTKcPPzLigfBYBQ2RDK5GH18qMdLsTJglq42yTov+Nu
ya6uoANKEH66FcgTm8ns7NXarYr2LF+tKNVyifnmH9XMorr9zNxT7O4CEVoFEsA5
Fm9iLpjIWrZMEnik5gYBGdlm4T/B5WjsZXLXIOXS18X6wsfmAEwDjaTHAz1DOOXv
8bo6V5cBytKbUwi9aV9r8BsaIZ2oV7ZNOMZzaZfurjUHVA80rFWh0I6F9yvdHg1b
MpQ/0K90aSoVdNTxBIFNXMk6TXi4y3Ha/+BWnmx++kGsn1tEPlCk7ZUmRbKY9wdN
i1kdliMqNudv0LBRFsRgeNCt0oBcdBz+cigF4JCSx/BEVserr3MldpFEcW9mHyAe
knFHQrPFf3fugOq6PBWt5U5GbofeWFnvnwHmJn2hsMTZfkUjD7iYppCt9fj/Xr9+
QWKhqdF954wOrD54/D2GMek+Vl4BLFYVooLUBHbGiDu5ZjE55eI+3I9TVkgxwbxe
xoXXzZMuvy7ITnBZxigF/K26znCckISde95TVFyAW9FCDoB/s6ftbh33AdYVufWD
tolcLdMkbtzSt53pVVAjI/j3Vb3Wn7ImGaESDznAKDgmjUXOzegc5NVCD2ClN/pN
jXZz2r/FR5zpR8wNtvqgZdC1T3MhzlmKVTqhfhlAyI8LiIw1d8AgljVW2j/rO7/O
Y6sIv1YJ5criypNg8877/PhwY5LvgIEDz2YKueHWisIqQ401bJ8IVeFWDprni6uv
CFKorLwbQZKuCdRFbDRGwU+7dKFAL9eTDtt4Oh8rh+yKBg+vhCUwMgxE09e8JSnL
b7vi3QjnJC5YFWHbsZj0DGRfZT4bCnCHUtdMbnyXK/po++DofzVL+aS9dGUKf3ew
dDI2cfiw1GHCbcXSaIsmA3Qz+aAW6JUNs1713E/GlmeiLeCzkXdYG+hRyimuLUCR
jxTHqbgEL5DxZQiyhAqPtBm/6xvUnwUOtpoluzS0HTBN6pGk8O4LOxPOFzfHmBRJ
ngfWWjYe3g7vt1OxU0EcS8520MPRNU7a9OdDbPnb72DAQ1cP4AgopTwB19h/NEQi
WxWZ0ljDBdiZVNMin4VgTzM2yvGMaxC+CBePNN3rU2sLuSLObg+hylMOOYMkHA8+
ojGIFLNXB7f/xatu0h5mlL/m5eQqOphWjOzUFTaqd7Hp20BVxfkpo6EwRpecjpNm
pjlGKeWd6WimxFP/HM4dvfmWipjKnwvwJJqETgVcMlgQySlsiizeu7ZxcrmlhlWc
BrY11nLSHxCbrwrzjd8hPesjKDDc92me+oWyPqBGP0SWjQ6IG4ivkKr2LaUGRI/U
ypYsn9BbpVjeqHczoumtr/bmMwsBJ8P6ZRkRKzWa0nycdfKLM4pnAey6T8Zy21qP
LsRbo6PgenuOxtT2wmgyu2BlOZ5YiRyRi3CWbdkPP286Vuu0GUkRtBNoV+bnTUcw
P/skJBGjYBnchJrtCsZtUT7zNP+A8bly/GJZm6X+9fvs7CkGeVuDwLG6/CP8Ucll
MW4E2NM3cVYngNFCwYT3n8nIHMlkOU5GIwfNdw/wXpl0hz13zN+N+vGQ3Jzvqmdv
FCKEQfoKvDZCxIswd8lnrdDZlpQfmIHQQp+kDV8o5cV4H8qtVIJ3HTQeKcmjWVOo
Oe7nweUbnheS+4ZJRjmzeeekkvxWyw08dW4FwU15Kscarfq151ZDIblHoOhtABmW
OAq3PdY3KO2W6oJkOB3UvA==
`protect END_PROTECTED
