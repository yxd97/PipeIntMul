`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQ2ib1gwSe6z3gmSDh0Itu3tAtDxPJvZ/umBDS3030/KXbuDRRcIch5IRDPbFUNx
4yo2eEnU+v8PxHQyfBA022CmcJwxbwrstlrRaRoiKPNUbnUlT7Z1zHOZuge32XRd
3iawtoTPwykS30R7Etbz4xnaxpejLPGzdmzJ4/bb6AT3kCv0EEVgUtiN4wxoiqRz
2D6IjdbOe2FwuvwNoBvb6Ugjcw9Ar6TPRHN5zCrtPJcj4K0xZWW3ka012fOXSlJB
cB/PkCndclmRFPc3VgYAOo5vkycnx/xpiTAQKn7EMLwFRBdt0zqx+VfRjMlCiKX7
lOxY9Fsm6hZwY7hsbRLYu98C+k53lFNmVwqugF++QgN4Oc52ZMN5weI1sA5azyLq
bzBMc4JHSfr42RiS3iyvpbKLGM4GEbsMmeftNUZgjA6i0pmKfu/uW8JnmHI4D1Xc
HxgPsIjhC/o4FZTqh3wtm9ROa+G5Nbdt2NExOsi0iCLfq2T50FTKjsYNwC+Ct3XM
s7ScTruhRLUR69XayvVEt3YxqdzGqB9b1Yb+GIoN6oJlpZxwXMFT2zXQXi77KucT
obU/9PpF4Llv3tGSK7NaYA==
`protect END_PROTECTED
