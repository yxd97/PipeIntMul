`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hDmlDwhSXcbqWa2RiXqHJdMYfkdyl5v8BWaW8Fn6wbVZIh/bqAbscUE8fiwVTtJd
2XJ0jGJKSHGYKc54zWSeI2zmhvRbPd8EQzvpFtdlUJsl5GTN2qouob0a9UFpAuzW
NkQlN1SwbhaZAqd1VrIdmuWNTgtw4hvsacPJmvnkJ+LvyxeBwOUaKtFfnQRJUsrw
MjV1yLjANBia0Fqm0VGMBP9h6Ocy5nvxEGQYBIOxNoJ9x0iaBiYLPD57qiMSdBmR
s/2nKKwyBzwksv4E+WVdNlOnz5KM5Zf9Yuhe/Rxnmrze+AyPQKeprh+BaczsdPB7
uqBRid6JZq49NKM3qgo4+3398t2HXomWQ1/JN4qStl/XFw5Ih2pLUj45oGTBG4zz
/qZP2VWXljphHH4yAGWjolFDtoIUwdXAMof9TawUzbajcXcvCUGU6EMS1n1Tij5F
Y/1YGTF1mwksIdcV9hMNFs365vVhPtcqK1lmx2w6GOU6gBmYeInt43HJftF1kJ51
hV0jihXXH9gA40Fet61NkWjNdbplEJa+66ICR2Hw5fwqJJT9g3ALI83XwBHuDgMm
lJL9QinRKpebS5jvugwWIABfNaiKbm+4XbO169K8xt8UlfAChBNzmVWxyCLQ/wQs
8mz4ryaOevc/Kyrs9KLNTrZnBHzjM5LuKQ7nlLSzEFolwb7fV/jGmVgtD1mSgkO7
jUW2z1HJVKNSnsFrU0ZKZXFbE6s1ctDoNShzv3G4+CbeSZpj8dtvN12UuKo/n8Ph
NxsJbBX5TlPM6Xve7LFmnBCoQxTnkyB71OuHnXRRIVYKE0vPgNtKNjJ5wUpNK8qu
2LCyR1Ts2HtxPfsuV/d3h9tIi0sK3lTFSaqjt91QLswCekOrSc1kZsepzdzXXvT4
7oXLjlCpR037UeDSzEMO2D38apUy/7NZswEL6Eru5D7fe3mCjzkwFXL45rBQIpoq
nft6tl6Z36kvOBiiOUcJyBGIwYVGfoq72DALbvyL1kLoFo5ejnHvxdGvuFjJbd9j
2Bg8h57UglcU1YaZ8Uw6EoUHEECZ3b2N6Cypz5y5dYnOaPEmZTea/yZH2BPk8jGx
/urpzCeEBUZgWhri+Nc5Rye9i1a23ucQKZS80tUt0+AacFXatZRq1x+xDL8Sr5eX
HFxpmS8sghtU2mmxKmEkHx2uXDWmaGQbOiv6XXVHWsY21UkRI9fifcolfbthFEl2
`protect END_PROTECTED
