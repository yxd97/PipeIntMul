`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkpEDQDdszzN2SI+mrnRmQJBynRx5HqEYmSxSG6NFX94zOOmznNf6RVl+ovV5WRH
YTb8tJR9d/Os2BTDAPFmUmaYzfTzOvzGZi/CqFwSuGGWepNteIfTgZyAJOCyoHtX
x+omHYYhkFYlO4XaVdB5nSyGqpNU4HGcmgAylm7GOUHDHhSEneSnkr2ZeFcEY6C9
WHBU+0qrRArUYiWQCf1IrwhoWLwKfxnSqcgc1zsQPCZ/xqGxzVjnS6RXyZAHD0Xj
u0Kxd/hJeWBSr1i+YVGpvetUiwKUxct9GridVwcF4eX/qv6NN3I37OEenypsW21b
d8dp2fczqyZJe9hb/gy/lmu04DkBue1lw/ZacB1iMtJf80zCZTs+pARt2CbtRE9W
cAOVmytLbSNlwd1qR897a5WgMjYB6ETMlUhvzhkh7P0K9g2h7Q4urJq3mfeeHdF6
RtOW8uryTtgAlS4TtB0Z5DFD/7cJ9fJxq392ZgHecTU=
`protect END_PROTECTED
