`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jU3UISrcncQ97S+PEH2nNbJ1YQ8feKaFhdxiWFpcqsZ13kI2yzz+WSxNUtKjndGo
fwqGAtR9JUqz43wWskkeTVH1/T5j4eRAu0aNcC/2zK99u176s/pR0/FOE/VG+mAC
XPOBdOSWVoyUhfpVsa1vBB5LnWT7VeFoO9pApnUlA/mS47f49r00kQs/XxW86NU4
kk91YADWLLinJhe8n5bySFtTy8pIRZuMVaMU0k3MzwhpEbozwQEtUrpfvXJdNMki
C60kZlau7+y8i7I2ZQAV7aYjKkFPT/JirZD5xwxnwo1VXj7pEVVPQx3YwQqkKvx2
CaPKh1ldfFUxgpb1o4CTIsCKD2eeOvo4hh8/i3ZSGmNQfDcRbSCqX8EkTVcjbpid
JFy0Hy5+BVvleY8qx8qDNV2QEr6qZA1VEoU67NkA9EAyWFTasnhuTw2dl3JsEXEl
mXIOvmK74nlhLRjCivy5mItiBraFcd0LMVCAIa0J1ZU43zTmbbMuZ+tGsbqLfi0V
PE/5bope3J/WLWbBvEtHNKErTox8Ku1pXnlJUVXjz1zAiSNPhhcWoNsiDbMKMmKW
1vQHPXVA0naPcioDdqn8rFsUODz3bWfPy0DEg922jgJfHU5+d2tyBwyjQQY8feWR
a9hxiG+hczDoiR0dPAWDGR7ICUF+4CzRbYnwlgvJfHVt5E6g9vt1dXt/iIU0+U4N
Mj4hCCDfe1/GPqKAdb1SvHw9sCtJTlxvhBcI+GP3a7ryuv0tF74R9SbJKf0SwT/8
T1xfLSl9A+oP6XrGpppncC+LDHLzdsUIpopa7IazHmLG6gE7n85DIAn6qcVqwXKa
QlyonehsBdIsUfuQb2R7aQ==
`protect END_PROTECTED
