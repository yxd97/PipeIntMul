`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HPxePObbl0tgl6W6pf68mElS0tmZk+tpFIMDnVd4cVjIOH4yle7vQlACApVFJly8
1IDEoIkrrQMDvo+Bd+hKptAeb315bvDwHebMK8yWmQdEVI4lG3NCAhzgrX1HirY3
Ddih0c4omj7JFsfdvq6SxWsFBWm7jKHH6Kyzqk1kDQ3PcQs+g6RCsQ6QHX8RcdhT
ICULvk3WAO2BJxQJX2V07YBKAkitVSL4mtzzdjrLY5+q3EeDTSXuYCHCPrzUjClV
bjA4ln9bMHwp/CEdF0/a2bHgmQhDPP2rP7lCsIT+aBbwTe0azICPyUrrVBulxxXQ
9nwBKbxTzwtnteOr4vWzOmeksK1HedegTijv9qxV6/ap81bq0By9EXpk1eywDoTH
PTdxT6rh4gNEXcnWwBZ0SV70Y3UfkcXbeqeJRhpv5z4UFqVYGhcWhvmd8QUrcOfz
4Hu/uXUyQXCYYhoNAAzbjruPpMsbSArXOhU13RpxmJEUSALckggs6QvCOa9NFEEW
eM4fnKtZAa7EHJvgH04DYQHQVmHeDfGSwXQ5b5s2tbZ8HCEpRSDXKuQbyL6lUZog
D9SpZSuK5NrOrfpHu5hxKqOM9KpaP3IYgWrJJhtHb99+bVcRPSi5BF0HLFmH2PL6
g6D+9IrIvoDHJRWpzQWyUc4rTfqBqiYOAAZULtuKG5wauilzDjp7sThS+QaD2dsi
FDtIwWHajOX+6WHRw8i/laaNeOUGuCpMXOCDjF/ibvdoyG2YlbLeBhkukkslagRB
EXb6M3RhyrXy8vuZF3T5UxgysbZ3q/VGLsh8xpXymRQ4U7+X2Cfg83NgXorXLW8i
k40jk9pvs2IGEKmDoaaTMb53xmRsXBhtbq/gEDfowhgMjwAoI3u/A3ssMnr33iWV
+eWfJrdTWYfpJajUq5OqXAl/D2U3QlWWpIaLo38rXGXrqH9wBJRBmkONK2JLZf6H
dMnCUid92k3YnF6dd1NQo3AjLmZOi/U+32Mel6r03qcU0D+ubRg7fmAqfhTwY2Qd
M8oURLieWaTOz1TBLL7YfffROaQNclErO+r1ycsCzl9+dycJ0xYBklP/r+PIVSLW
d8IYxm/9QlSx2PyMXwIEhCLfEN4Xb3emhDXT+Ksjg/TrR1p8XThmYI/jyTkD+5/2
mEg9rvk0CizWJ0EtQgo228ZHimLF9J/NLT/sS86fl+XXBSZ2HTxnEx3ZUuz930Vr
MzBg5QPy0nOhAwIkswBNysw6rw7oU/ekce2LctdS6lVgEtgFoWvoh1WIwwlXnb7h
4NPXWu2fUIv55rCex+AwYCjxznK0L5DaAZhmois6GmULGVUILLVv23Yt/aiHIfIY
yCJZmwf9/EaEAGAmK2HAStO+b/AuSt/x0j160V4xpM4ekgBAyonv2nuMx1p0uAjA
QJQrYFbilGdo+KvHRNlvdHHz6RIQoNvBk3lmrjVKOLUOr4jG8pOJTBk3vgtCLjMl
eh7wB9hOoxxh+9E920XTosQlLUapnInVfzwk48sEaSLJp+Bv3KqGoqxNR5ePOyZq
afWj6hScAO4oYUbO6RQpd2yNmUz1HO2a9IGgExb5kruXqouNwSdRQ63y6aSrJLIZ
4RZIW+h6ir4E6ZJGNosgoIOiqjkGnz6G5WoQ5FibrPvrQP0BNtaJ2b3CFN8m5Vq9
ADwC3dCjWKDpn6VJ6gL+TtHFYwiNLJ+xe1zyVhiS+DvKKRdJeT1EPQygF8q+LGqS
jWqoxTtmWrD2SBv15e4CjtQfKm0GUncwPRm58g56JmeKrz7ysMSfUvpbRovO6Cef
B5f1z6efs25A+BnZNzHEh/PZoPE17boeqHz3RNMDp7A55V/jpzhZzpKHiC0k03P1
Sgz8Zj4XyVrGE1OLmo2KHFtL+arZTbGKZQXSNNpXEdBq7yz9NqUUATSIgh+JqH1p
06719ewrLIxiDKLmllUXDi5RpzC1Jw0F/He2gsiDgRgZQWdOOH0pjQAOotAP/BEC
NXxDe0XWgn2gwHC7tMoJ19MQDsCcaLGwb/IuX3h01obtstRVGM56dTcLRewZdOQI
NmPNUJM4qNaXjKUyr/GnNXar628zXefiyHJ9HO6tcNPLNI1IZSzoi6q/Rld2uO6B
/a/vud5oNETCutxTRbzLWs+nMy7cjcA071aQ0z2JyI8uJ08vcKFnhBHPSt/VZVY0
qd0S9cbKcB4ExDmODR1i9xIAzEAj2kTAh3g8VZZCgxvzOAcli1EDjxhSEOVFFnAM
m7o33zPvHTeBwFc2YgMKuLjinjegzb46Kbz3vkm7kT14bfcKIr68mbLIQE6pqipi
lUe6EWgS1UIU9fWtDf8ia6Bwrcoy7Y8RvOJ/dZDSzP7v5NFrZxsFNDN0ldLO+YC8
UDZYdh8xXqO0o2gCa8TU6qLJaEuRyrRcVzXu9DerKkYDVZm6tfwVN0/Hv4TRBJ4H
mKuu1zMByERYRECFd7EikeLK4c+o5fQ65myLnVlciMIm2K+p5rOInsH30sH041qF
AyJ2NuOQCXjcvdghLGXQt/k8bnhlEniYtuXA2wgKON4onkhYlVYZf297bAC0Qgke
1n/ePN+zFp52c1tRSCL4fVbN1mlp/8KrolaWKbBTuzir+gA6f+HhLnL0R4oPZ1b+
xMizsCozCKRwOKnQGEnapgsm/DY1EoUri/O2QE7Ai12/EmE5m61FeZGBeqy+aHxj
8k5WT53+ZW8lbWtEmRxtS6WggcctX/5xlxwD8pU612UHwjHlMgUx8TD4p7gZ2OUl
W6ngyw14jOzi/E/iPbThuTd+FEg8lMWlvBwerHouHXfPM9z/2rrJmm1opd88pyWa
8tFcgNW73L33MA9frOxSZ3CwLFnh/UzfAst/lbr1O0ftczGIYaMPeQ23UsB0Esdg
bo1FADTATO5t3Q68hJy1IW5uJb8voRVcdn7NC8nQ152Jw0Q4HQmjfX+DBD2CLZA1
m8pgif8v0KIv6kH0fNqWxm0dF7S/tXMfsgRpUK78Et4vdY7TWh8LczNbIULmJlj1
TiXb8mGKdG81EI45VUX5Wm49/FfTUwMKA3+r3HXWntxOMt1RLtVfQr2KGjkXURnZ
NUHyRk8l6HgO3dWSmknKdbld3emyqNZUHkOA6mLQXStbRURD82B6GzRFYwYAnOrN
A75KXYSC9iLO5LbhdYNUb2DloyPiEZ7wrRICeHFSQc9zS0lCa1pK9k9AKkceoKX0
FKIqsaJ4svvq3DBQXbNr7bMCtn9G4W75ajob+f9onr4REM8irOAdjM1fRosppptB
G9B/4QZE/QkKX8Z8j84siH8tS0F8ki5vAIidK4nvsHMuucz6AXDX+0EKV+1rCyed
I9Gq1Mp8VIwKllw+ULe5QnV6VGq4V+MSq/Q7m/drXueurHVjBenmvTUeqU9hUXRR
0DCFkKNcdhF9aBlJQIHjIQ==
`protect END_PROTECTED
