`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/P0iWFCQUCYFF/hJVMeS+0/z2YE44JXDZUljak7+XaEHegm62FUdV9i4FoGDYTg
XJ3o11EEQa9RMPceSSvi5VqJ5thmQ+uHorkwU4/pRAgT0OcU7r5HrqzdpO4pZ/pV
6xqjl/aSHgsHmlSG6bBFNjPCqNHLkPX/fQq9/nNsl4SdAYuwKhgA0A21c0wZ5pMP
FWMpBgHx/7bOAhjcZEgX27laIl/K/GbLbkX5Qoq3yQuN/gx1OVJ95kE2FM4OkDsZ
FldivSLlP4Op04SwBQeo4qhl965fBIZRHfCY8IsIZzPRD5SC5fodiWJob4dAl/kK
S3VkLROZIGMGnm5QLqaz4zxdFvN1Y+t3rdKTk+NVVeHAbl5k7XOqINJd+Jmdk+Ae
H3q+P5EacXFvSzwwnCfHRaR8DMJrxqcDiLmNYdvG3TT/SvCxbf2c6HPYqff3Oqds
`protect END_PROTECTED
