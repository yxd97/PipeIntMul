`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yTiusJr04boDpKF87OefwD51n70fJOk2d3eGun5jcocH/1MzH6ZkxIwnhQvxpZ/
d3xbUHaWfky7p7du/PLb2RYhra5uu0RI/JQY4zT/68ikDJvMf3aoeKpRAyhfnkvG
RKW2FTYGTt39YGIqFGpnME2Ej+1KfUV5O0jTY9VJr8NYq1L5K9ZMU4b1eaWpT8lj
KhR70oc9JOUHEB5QUD1PbUA7wMXOCytLwBUVZv8uT+xzr57Annm8tURMUzxPG2d6
6JZwmlnKXMR0cm2TLafQAwQXwRXSl085H0Fj2dZrSIPN5qzYq8M+6TlWXb+vxW0b
`protect END_PROTECTED
