`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mg3J9OR8Xz9PnDIJiX6snbzy7u+w+qbMNyM05EJPEW0jkY2/Vv8JudbznfmAv1yb
A9qBdSonMA4pYnC4JqT5p7iJxS633l4UA2qLwoQRMdlkm8K4+1qNNeDqdPSzTzaG
+Mp47U/M7Sq8+mqFZUIJNPwRI1dAgMZ0becKx/3h/U1aSTolGkkVkFWqaZ52/mri
nzlE80eHIYEt8LOhlSBgpU5axIFjywS1AG2RcnYAysUMwbM1zzBt5FprlxiCru+2
jRuZzjLKN4Ib1X0M/HYeKu/Q0Ljg/dzbIsnlVumIH1acfGeFaMKiz//MNTfiyhLw
8odV8Sr5VonHYSX5sjoYmMRO73PQdREGzx23E8q+5puyT/AdOFWWOdKu2lQuhl7a
230sA/uKG1DyJboXew185K/WJbmVZnNTSfvHN3tbRfyKgI5sln6lslwL2rC7xryw
jJhWHOqQH7W6exSlXVdvrGJwVGS3hhq9GKyWwKsaLZUwehU8Hj5ywhG6Lvk9b+F3
WYcYbSrCu6rUaoJc5VYFk7Q6rYtCE7aM9NgQF/G6IxfJKfSLLF3TUNjya1Cjws02
xVASvvlwDm3pHITeHHew5lrFalFilCuXCbJvIYbVJNG3PyFd0Nl2w31y2RBhjLrv
4/9mAiyZ5nPPoxwxv54Ue0l23sW/32M+euPWgksgjI0bF65gSzqsyYAOE+syo2v8
c06o/ryLG2hryhAzZwyk8NXO06HTBki5ZP1iTOf8TWzBJHeHXFM5PqMpTZYcSGbt
QSngG2+6rqXbaJltTumzLH+Lcp7xq7Xo87fl6X7HaOeDb64eP1trR7Y880fbfwtj
eFQdvvfcHZsND1ERX3Bb2sRdXZj1aqJs/MM0ieq/C4132ZjXhyOzPP0H6TG3sVn7
AHpH9luWUTpEne+3IjLZK7PiL0IRBz3olCqcOyt0cyjvl8zUyqdoWtCTlCUydZ6L
`protect END_PROTECTED
