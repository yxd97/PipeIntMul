`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Hok1Lq1HX+eByDJ9JxaZYLko/dbkUxrChatnipIrNQuhkTTt6GKLclqVbqYCabl
IR90Vys3OcHochmWkwtwmrj+WZN3noSz/vH7DBHQSEoGJ1luMcwOcSl0Vk7ssPYT
ykPUxvafHLfoIsvncdaFI0oNhDyzMFLWJGcB4cRWhCrjf3RBvwaDOqNnmV4NwDpk
w3ptLoksxp2MI5z6DJC8idarSYlYybggTUQvWF7qr7PiLwTV4KSaABXUTwlAUCFc
yqD1ZZo5+sfMHUZ5eGyhXsyKn84BPOlYFmwzHrsKVLqzLlLT1NNIFyUc5maj71s+
5AjAUx6VT5t01xP7iRy7I53HMObS7Ahg3NlX71pt1mG7Tf7+LEFjuVwMbc9DrIAL
LVchTNcszFcBBmzVZH2Z5GkgJKuRa2A2zlD5TZ4DbrNSt9waQ5FgqOEKlHeuMpOP
3yXTiU9IG/BzFXK98LCqxvjXzM0sMBl4H7MuoQHEnX7GqmQs429xLf/5vQqECke2
ACcDqW5wRhvu//ZgXKHjVLSzD/H3/7LBTI8obfWDgXiXRkElnGb2g1m9+JOidNfv
Fop481NLgBjlqwAaeysfdemge5vTN0d51nXTaMFF5z7wLrOyAOqEquyv6V/icWzB
TNItm6eKUMjy0EOmQ29os7IdqJ6kia/G6PbuYKIDjESCRUVbiyR6F7eS+JYMDCj9
3Yp3TQYK1bTEVXpoLVX1GUpUs3Tyg5gZ0HK7f+uuDeK6QLrBcP6N9cPHB1pWQYg8
uf/EXUsBz+KNOh8gavRr6xl1mhU27f7njwCrJO6atGohkbgmvnYXlWXHHKQE9nMk
1m+K6aHYmmfESHVPYTXC2lVlByGlXqmQbzJM6TIsjojdc3GJ0JWfdNv+VcVnaXrK
PDS/mIAMXl8z2a7h+4ERp00MNKipBpqsGRMGetS7jYab4+sgKMyQWJMESYpLlDHC
`protect END_PROTECTED
