`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2Xb4fJudfdTJn8Y9Q9iUnbAA0Eo4BmObu7TapBcKw0pJBNNALNkhZ2uFLzLYx2r
uz482LiwKODDnnBgSFffEy48sDMlNavNe7pMiHMCXCr9TmAaFpFCC8dLrRLAmub2
T6Rt3dRNjvbBhjTOiiB66VGgzv2fc6PY7nEyUDBBPDBUqdgtWXsYJufsrrduoQjV
iAKojwrPaK9iTiieLTMi+BU6Ms2qPnuPbeAAbVl5j2b1oMyXD+BTeqhv9Scp5ufw
0jFUTxqEdpejHkkEZ30mttKFucdoLVkG3fueo7cqcm9SYwyXK9Ni1MrkwRFRn6Wy
4MnglDQrYBC9HdVTncZsE4V5rIKEovWAiH37ZoJmQNk7OgUqshvu93z3i5SnY3cL
GAqxEIhdjuMXaNirBfdBCHrGF/jWidxLL92xDIxP3h1uh8NuaGldwCyK0SbdW/Jj
PZkoZNV54TuXQePOutrCb2fFl9PPj7BxyGJ1jm1DKhTpUKRrD15j4Pa352xVCxup
`protect END_PROTECTED
