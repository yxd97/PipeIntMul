`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QTOsEy3DtdZNBQ7/rHp5xhiU0KDGxMIBhUO258OX8ADgUGoD5PA0wuqjYGZYuXuc
e/DMe8DA8GVHz3p8cATFXqRlU+7bNJ43u0Yo0fFPk5MbnRrYgRAdsA+zgQ6bgBOx
uTwigL5G8e/1lyRi3Mr2ht5aCR/tnOf3ISnVU8IZ4csJc5Du2NRuvUqc7s6aQUDU
8USCLtQe4cBjGlwt+RPKRe7geQ3sqf7OUyoTm6F4DEL6OpwUaiW1oaoRrTRIwbms
a+irNs8woJC19CVVCT7WXt7P/D4A+mMNgvfi2UHkZY/gaHqrIOH0x/lok+brkWxw
XL7lqDMGW/YK4/LbygYSHlqASpsCcNcmwaT7ShUY6EHXkVPIpZroTh/yAcjWxG70
rmTgE5OscNKh63JVXHhtNDKsdqPAbJ+4BP+5ZT6HQ28KcFYq12kmz8KJaIJO68Ze
bVfop5nlBO63/4Q2AecHFE7EZgk9eEx5/D07pS4QM980Q0eGNasggci6fzF4F6/F
LbQaiGcTngLHQ/emIsb+7IDj9gvCD7e9SaNPUCJWYDjabofIVHSXTyXmEWeoN//z
xsqDsMs0QVzKBM3p+h4eGOIP6LreBIvAxU31yX0Y6Uq3xltegibb0dNu6Mi6Jtwr
kQe25X7jxMcNoX9U5UJ9y+aM1/m+rjHOXt1Tmk9OldhDySJmBNp9I0ZShjWt20k/
L+rRG4L8ZLb6Xo8ETyuEI+Fxh1xI9jkumvr6Fmr55zeZwszYplWWpkOixm0k8+tb
/JlESoKLzVbcBdYf+NT4xQlBlvLi3iBtq2YptelnEPUPrIGTfjufW7XJfZrDhMvV
H031+N6UIDqTbQLgCM/TeNumOxyZ3QY93EQMixeWP5w3G8pMhHrL/C8u+LHyoevI
iSk1lh41Bn+aMCXRQFZ50Xwys9iyVqiDG0Gdci0fbo9d1JBdydWqjBngfyQw2jsu
3c++s3mLGyVd5E8mwuRT2LrNRd6x1pBPaua8WAAtY2FZUDRlz35+nQLmgtnm8WZZ
5Bs37nE22o/77qBz8STnPA==
`protect END_PROTECTED
