`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzURhmS2wTsoYmb//cQe0AWE2/WIfuLk1vYI3Xd6GkkFpwxPPQXNMr/bv3+7WuRT
lukM5e62GgnKBNAWZaJ7tTcJ0EAJgO9hUex5AyVeWidtsfAPKmy7ciWSU93lNCgb
cuK0WowLfgl1bgBzJsjGfIRQyYEnrkNeWcQFQYquGLX2tHDtNpFJFBksiUpi7NV9
daOa+rYi831ArjrPMB08gd+5S6XASHorPxnjySTdsXTrUrRfwsJ0Eb1YeI1RE66A
kNaA6ydb1UyAZEr6hN/SKHm3+cu4qOWSQ2njjqbvd+pChfsoP2xPVlrOg0b13eyD
tT7fwoMeKkdd/rSb4lbeU0pWDolGtx72renZ5+A8P7affv2nzSexfKxhlbNbDH7M
UOw5wL0wJpmQfNdhAuETuZ6+59ojZqmHyWRQYxP8KTFSPHhTy8sTXZyha0vTNsac
AU+jiflOavPXaBK/QARguxWqtXqsHiWyiu8X0ueWuHIfsEEtsF97f3FqCsJ4OFNY
`protect END_PROTECTED
