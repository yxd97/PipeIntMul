`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2QwebOBLvIcL0EWWNK4Q7lJzw0nzR/srjmTZMR1iw2k6L3RllG+LXGEASmZZH4xa
nyIBlJzA6rGgzj+Qj+Po20MlMkxTlFzSneHO03zvOfTHcz3Cp/cCqh8NJaLcEhOT
ZY1fGnz3Bk9hHuMinepqZkmsD/whclVLB1/gmCuYzN4FWf4JwB/ZIFWpsJ5hI9Rl
AGWuhCzle2OgbnvYazUIaYQ/47suo5BbYQuU0m1SwFBtJ1C/o1mMF/tAIHQ1yhsN
O/dodrv9maw/ns/9JGe4I+KQt3mS1TiNIPyh0K7U+7pSKMBkBhOLM5svCS+MVQSW
00NTCISQUNv9t9YVyAn81W8bR1E08VnypG5BRxhXeumzTeZaWhSw1cNTfKJOe1ab
H1VTnPPau2jDI33BqBEM6qlVbjmWIZXgEg/d+7blHy2NZGroxJYSYvN0Ujjllz3k
aJQjP31othfe07kRv8EM/HKMJVcO3FtzwHf7+MYGYUpOq+dp1jDecqF9E/ajyL9V
Vl508BY5Iiet6LAIvec98A==
`protect END_PROTECTED
