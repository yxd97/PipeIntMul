`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jUSCRLszBLc+dsWHBW0Qhn1LGDUhZ7BI3AKBPRLZ4qD9sAjX8ZbZR3ROoJxJFI5h
t8NwIiYKKcmQnhTac2y4rMCRTxYtQzRjFrDKt0/OiK8j+RdPH8SkZmCjH1k+yQKv
lIeVfnSWzbtQ073uRjWLjSGtjjoJ4X2HxpTBru51e9eQGvmql4ZB26zyi+TeCZqC
lpKM1zPWC81xoLxqQmBy4DUJw2ttspHe0ibcEVZ+qJD7/Yhhwu4TFbgN83+XgcQh
GLs7vARwFPlYnTW29vDz+3Grb+mloMaqnI3L/bVUQ4l9h6z2aYV4F6yD2ifOZYrs
+W7v8GoB5ittj1WjkPaeavWDU3K6Ip1H/38YfqgZlAyeCMRtWdhstEPp6S1UCHFF
oXmto+qcGCjOi6i6nA2r4i0J5o2+HJXspkfjjQkl1ILxNXG/SWaFC3wGv4sOzlLU
cg0hhCvpjpvZHMr6pDK936Rk26rWadRmwuMUpHWIC9osNJ5DCSV8gw+DVdU29u+g
J9TiJDSmQvkfUu0h4lQ34W7M/pCfNQXQ2alIwq3oRzZUAW2ElELvdTaXPXyWniID
Q1xvNIL1dQVSxDNZSK9+FGNQciXvKkrJ4i38pxfCEgY1LokRUuqMKrx3M4JmurLz
dtwEkvbikKi8iW1EjHxiQCZiKjSEadHXsoESCLqQzE/gpj2ZD8PD3sGkQ3ntTyGH
aKxqZniOdfg7q9QocZ33iAHLtRE/6xTmte92zZOB1QojtAiFmQC4vwxJSE1wABZv
e3YkfV9qKWexL0giTX7R1A==
`protect END_PROTECTED
