`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hi7tQ1Fou+XUaTtAX7BNI7sgMzussA3LeljMAC/R7OEH4zBdp9gZiaQ+JBJFdOiD
ThdOlcetvyLcNVL4/mJTmobfrawkrKUxbndxRFR3ortwUuF02kSvUTz/085WKkL3
UjVGtwWR30aieAjbrYlOW1BmReKH/RG1k+yIB/uPrOtVoc3fi7mY9lqkXLZYTj0f
eA4o2H1VZ8Zxw9QTvqmMqySYo4j9zIWaBdzKWovXSWFnmTpGZRiGsIDLXZ43ka2Q
2GhlJoonm/L2j6llwTccWg==
`protect END_PROTECTED
