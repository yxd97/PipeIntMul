`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6IEbvyb1BWgiB0UfKl23Ep+SI39exf4ccr7SjeqUbUaS6DWisWm2zfwqqTbZ3gT
17so7eTQOtoe6J44X70X+rfw6sUxxvJHovbm7Kms/FkXZQ6s9o4AUYb7Ge1a3bbX
pvnb8oIef67D2/baB7cktNFJnN6WwdJ5v0nzSLZOdeB7/ICAyOZufS2XabcXYIvj
iD0VPOdK9UQOr9P2vSnRKWJPnhfe2l4xbv+Gq0HRP144aheZStVgg+7RtGgG161c
CLzdRvWM1Yp58kKTohKt2L/YReYrSI+Gwe51nLSCat+p8qdN4EE69zlsYZzGBq8o
FW1x7EnEiJQx3TsNOD5hQo2v7JJt2ncGhko4sHolWaM=
`protect END_PROTECTED
