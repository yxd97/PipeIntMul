`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POHneZiqULISwWSU5yiAat+1IIdg6tR/7KBd/J+tl2joTdf/bMlEY6oOlGC4GSVT
dNRTtFoo8xNCjYF6olwgs9lsH6wKKNyZXPGEbECr0WpBPZ0gPz4JKVEk4y25YooK
8BZ66uOZqyaWRXbrc8QALsRwKT1ZXTpMaF+BnmrceAWg/yBghMZhUnKB/ZwBf3qA
A2epVDvecEQsLHf1zStZT15BArRJEBrBltXmc2l++m0Rh47NRomkn7AslocW/AJL
/z2O4Oh3gC50M2KrmIWMZL9J3mpVDQPK2CCjUrWkTWZdeQP+ntVmP7eQ0Dj7or35
MN/0/wLdJ1OdqKRiaoQj8XArsKdNvim9zsohw33/xqtHqFWXi611Ba4vAJIcfGGQ
fQPzGJl+9iaSimkGWb+eOFtsEOAsiDsQTxtnvxYsVV8Fm90IKNPKAC10iumLpZoJ
I39YwbBccpKn1sZIM+6FaQR9LOOPY2kfT3hfh+/nu7vxGyocZB/QAhJt6VoKMDk/
NPCkNpUE+P7Y6CWtfjeYdvq2o9Nnjq2AolYwTf5dbjhMwmRQ1VLR4am6PQuIKpPR
kQk1GtI2ttKC+5Fxdv03VxRR4tCIyZPGiuUE2hSBriU76VNysHOMLa1zf7vrpJOM
ipUcEHv1BMjSmAjfxQ6JaQ==
`protect END_PROTECTED
