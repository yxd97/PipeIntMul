`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f5+XhpfeOvpcXfBI/iar+slhxJCUkfqhUOpW6ojS2qMvEmO4IiB3P0WVD0EKDlPI
jYPu49GE689fDRd7NxDYGJb0VKSbDH3oX+0fwDvClvrZHR87XD35Rj088VzBrXJu
5YtkBckj83KQICSRib2a2kuNCLqOXH50Rpx6uzBsaro07j5+M0Djrhd+U82JgE+A
GcqlBqy3FlQ5lfFMDN7jPXPRSI+aVeYcI8bn89/OcGO2DlYL8p9+PM5eXhy0ePF2
w9ho0lJw4usqYEMJ1/Q7sC7M27C61dIugjc6k32Zxe6kSpw4QASThwrv8Xz6IfjF
I/DZjMGVR4fdKMBW7scb+5EJAhb67nZaYWjFj6uiA0x/+oFj7/QAUfd9C8e6HeDG
ezhMu/59In935NUDOnFZ60ijFmaWhdWArBG1oxQXlxs=
`protect END_PROTECTED
