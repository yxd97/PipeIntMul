`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rQ00bT1DeHYkvjTSDwCvlnFbtTLbaw1YB/v8EBeQE9HTlBCdKvV1OUTtlL/MO5CS
EzymgtjdQTJRHenCY1NC089aqieGjxnI8+RFlMlTXc8qWv8LfoUGyGrz/CD1kMr8
hmOnVLYcFlrjW1K0yKlNZFfmfWtIpfKludnUoTcu3/Np9dAF/UYmx/54CgcjJ5uP
b2CwTa99q4/t46P8I/wliPik+p60U8Um6SknfW+5MoN8xYUK3zwV9GAkmGzDlqKb
NMjoljpZmTRXwwX3HEs6uSC0x/tZROEIVDQY0O/7JZdnJfNFiaUwk++M9rGSsJ0R
37+N5LK0QoG/88gMBsY/392Y/SiL3gTtjuJf41PSodsAAUo//WprVAU+V16zMyaW
CPRfGjUyz500O/K0+nkj9zwQ0Jz81BZYv9LwIKLKMoadrctofwWDM2ILcWbANc5m
oJ+EDtLSpaTDaT8hbroanZwLnOlYh5VAjGXAfoVhycy6yMuTEnA7RazdLV8x8kYM
HCJoQIr8sOamdJ76qmjWYxKZSLUvEujc1IGAzMYNLbFTbMKzhB3WUjH5MFfa5mA+
zgsh5gbaQMpwSJQKoxTzYzhnmQt42aESOICbL1LREeNojttMsFZITtLC5feR7ZgQ
BIejIQapyGbgyvcGwWhlzw==
`protect END_PROTECTED
