`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0/32iDvFEzn3aZSuDtUcBp4skmgfrw1ZiLKT7Yu7pYa9+s9yr07S2pN3NzJlisJP
UXKdieCAZXqBMJNWdGWCNy/2pdEnIuLRvDf0/5489c6odvCbDDZw1PlLDFVV6aCC
CpdIWmszPBGk/rpqi7CCT8I/TS+RzoVt4RDlZCPJeOaksGCoEjevp4US+80ihhuw
NNcfBuhRqFFQFwdti6Rm3xV1Qct6y9BQkndlhmH+WewV0Xe0Q88eW2+f0jVmQ3ja
Oz+r1PPTiIFOQ7mMN1rJR0wlFwGc3HeIXqinGymFvMsQIgi/EDGsvxu9QXHYkSPK
PMe7JCAiSCyEcgeAqpFY0Q==
`protect END_PROTECTED
