`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iriSTve6uzM/PA4aLXQ5YVfirdXU5cnlMqcMAmoDSnInsBUQRta4EIP/LptifDRr
2mOE5nXpk5zzrLGMm0U/sV5p5oZtNhwPpKP9Ar6123Qwdc//x4asI8OxBb/nhu4F
Mw2TL+yGyFUFWLxDgkdPUe6CqEfc+swV1fLBVUPMergB3RzrObzVA2ekPnogPO6N
nN74Ql2Au/cS7ff0BSN75nuqY64MPkAoydFH7ED2bak4BQm75gGIv8h5BECNxUT1
cE5J6iiC35mScPDl3unk/noYPnbLN/N91HorkT6R00LzIy9wUcNKKdcLTbXg99fn
5nJNdiTZWTcqdZzbGLruD1nIYpwk2gJyng4oCyUh2uS0Skfb+/F527RGp360827f
rO8opcZyZtIX+DMIl+s+wHzNzbFBOtUa0TRWxDAJ8HsMU6P3MgevoZOkqELpc7X3
4JEJuZY58cyR6WFj8TDtSr8x6z97t8VHgF4LiMHKncxIlsKPe1IJkEfaOa+bRgEf
3N3KXKQQKg//CvL8g+MlNYXWadikc5NKwwm4u8gXBGPa7dZqqMMaLKpkTuc602rd
ftsqS39pFg02TC2Drl9Ze937fV4CFq8sZ8hu2hxCA4T/QPuAn9oss/T7paHm55Gn
syx2L3W03noH/wLk5a1I399iZMoF9Nv+vhHIhPj6y+P4duq9Qs6PowlrGPIiEXrl
l0v8GeErmmWSzj5578UEIV3liGfiLYcPmZd6NBIXLLBw3PZxdsHccBxU4wlFQjAD
EeotJr+O5hSQF7Y0jufNoiHHsfxhlxJjt1if4npZsinlCjyEJ7MFSMBNdgT7qZX3
kiYNQUxSQHMsp5VOFSOBTKYPilF608eSsddC/1D8xXttuq9RL56liypZCPcuUzy3
H1dCBPKyrxLeKAzqVBkcR4L0XwOB1xZTr2JCowy5B6CiBvtYpJcaYk2papyUQ35g
7mdafva2WW911HurRLmdL1tiFHZWRACBVxh1+ZEnCts5MLi2dYAeJ8IgbBLbrw13
5Zp3cOBNdYKuQ9CDS+4Fs88Z+II6161/aJFtPBTpxqvKlZ79jHXicFsOAuBXy6zC
9mQ5bVP7wHQfSos/7ySFza9x4W49ZJX/SH+HD28mQNVeEcD+Su32qZWOwxD4oFZB
G6U+tDlEkBLSGVf7P5oNvghHadoCchcGon/+lldULKraPRyb/IMPCOCBwWSSlk+d
tlrF67if5gXHlrLcEs98jtGlHxFkMCvveD+VaaNTQd04amQS6PCklY2+23geS1Aj
ZPBY9sbqrotMQBHplXP86fhnkM6VAIF0QCPGQPxXdGMDnH46bJ4Nkxbp9fdkrTUj
/WvdXlHzyMtiAqDpqgpI5ND78l0RRQE0kf1+OIowFylxBjEDqhpxjMTD0dj7VRDT
7t1wQuBhdm2nZwbrZuP/b9OEuIAQ0kCXgKRZ/peE7FmNM5uNS+SmWNMoH4CA9l/8
MxW/+x/7FsWpPwCtNEZbGkfA09EhF5vbcX3acxATGhA/qx0PedC5cVYyh5flvLfd
NbvioGVOE9QDyVZDN79sfdEHUkmm4TxOCz4BFLsg72MfnUj0+hvxhpU4mOWk175B
T6wWkmFbv0biwMx7m187nFuVfDekeXdul0JGo4l37itv+2HNHKKterqpYQCag6fI
30AMRaBIDTbt3Lc515eCxkkPjKlNLaeQJ7WAImfImJz3Id5Uet5MX2/7/uKvWpBS
ZzSO9U+M+2sJOnkfIcRDYTO/cn802FQB3B1NaAnmHVUJTwQyq+JKiEAddC2pK1As
Xm39OMzoWKZ/Hr/KNKKPWfocwgw7Iv2skTjDoxZx5o0Thd7YSX5IX3DippIRTNjh
iBM9eKTxa/SIGN/qSvbYV32/lGfNr5dhkBt4+9N66nuFK9EbsZ+bXpehudu8KmFi
dX2A+FtVihrb8zWOva/cTA/AOd67c8zgCYT1ejXUGNoRdvd4yW0X/rtEug+zvQbO
H9Okn9aTYMrXYJg30K8F6lXsrFmQnYH0KjTGZjTOAtGiAt7NVNxjICZ5x0v0h3SK
1Cpm/a0jOEozp6UP7PwfA/n7SGigRlHatrK4y+UZwcdJCmreX2JITVU2yMzwDKFS
2kM5FLDWdmkQL7+PaprztXK3cFEl2ZKifVAWC9Kesmr/fmUIOCDax7shUnvLNWvE
OJq1j+TXDhhz+S/eLKVukObJrl6NdqCH9Ujz6Xk1wZAQt2utaeV3SKFSNesZEXpR
x7vF1MwZpq1yviQ3siM8hFTmxs8NOdj0pJvAHAz2n5PvhnYmhWrxcNrRLT5fDrEy
flcWQKQs6zsJYxWos9/75vHlK+1oDwt8+C6mCfLcFTb7dLUAz2Lm5sf7UQ2jkcGS
oTxS63tQi3c8mvObaXPUF2ICpDmX/FS2MuKVC04piPId79vj4Spy/YvxQZZA5MJI
OnN8zUPsS51I2u0gBbhLpRgP2OPBnAnmd4HL8oO2sBg0f1n4X6itj8ThdAr7GyHU
k2yzV2aIbbzaekvYvCz4sFHMd5lneOJjhMUfF8s0dd55c9yl3Ikh8XdESZl1sG2Q
FBOpEuSLROWJLfYujQ+UZNQw4rjwJ6cdMBioQCQgYzdPA+/z5JDGTTfqYRIOlvbm
4XU1rgpwrN5JeA6gzJp4RYwLSH81fwa3jwpuAmL6woFMjNpFLHs6gui+IniqyWTw
IIRkd1JwMv5Vuce8DVxteQWSdOqaj+9DwQ8BNW9UYGOS6kRNAbcSRUhKEFJQqfub
+yqVJkzoDcO+44Lx1HksIa3LEZ17qDzMHE2zgYarQR80ExrXaCTHrMzFd7ZS6414
HKHbQsVMzGzCrhUs/Okjxzu1fG7fVtE8CF3hjjDG6cJQGxj1x1lw0vbn6c+EqDvO
TSvl/NjpmLmbb46hiwAnbGWkGydkopuUCga8QNXvP62wTH6aeHm16Fvju4ZKOGy3
wPMi5Z3alcgsXdz0asbiYQjRq5VL3gRspcBpPA5RrtH7XagipZwBNoTwZv1/yFOY
RpyHvaqnOqVjENXx4jlxqrmfaAnOZe4EGEvjTopxoMAAOnNgkSUiVuYOqqTYO3K+
GHzYZPaMfauQPbZqIH/ZVDhLTTWU88ECHpqrqW2wlu1OuQ15uf44CInSIZIwKl9r
URKg7PteA9K1udMo4JR6LMmusUjUEL24ZxOtoQYe+A6TNBWeMT+xOBDhFlN8IzQ5
r4EosVlobniQGKLwWWjnvB3tKOI9RssmlpVCXgb4Tt8H2JdAdTXmx8L/cRsNc/bl
lM9h0lwOdkRjl/CEXLf/EFd8EcmuAUHDo7f8qGbSPmWbNXjBhGYNS6oBc+T8Xmml
Y5RWB3/RJO+0FdTyWok3UnfFtajb/+3o7x1vCMW0n2fRTmQfiO5oqHxpz5ejin2Z
2Xoc8JVij+zUV2B8OtJzXc+E1fcFnymJh5gE43Nedl4lWfKrcKvRdB4Z+Aa0aBdD
nt+vNK/xAEBWJMRpMPEdzm65moeYBGPh0ta1ECzHJFIhlubG8QBKGXs79o5Uwmyn
ZYBUCTFziIP1SYzXSc2F4bKekK0djesyiQOk9/BsZaXTYhw1C6DhTpXfja081sAj
H3WzWyMC9ziHnSEAXOAsz3VqtkHk97wstRaFmaGLLpmLVjRAuhI2SFCY0e0LuJ0P
wUhyYhkHBHpZEUtW3UwMNMEYxdfjgHYLhn85vBD/XJ0Ve5QNkrcVteMkAkjLJbhX
sHYA0xn4LPDh3VV99BjZdKL5nsaocH6zh+ukvwQN+xFwhrxpTH3yRTnlfz8gnMmF
hNaiihO0rZ6gpJWh38juwPG+SpZifzgH7UQXVw6Iwx7ZjjJk8Osxk64HcCRD9SuB
QLLz2QYWoq5or32jlkvCT4M4evAwTjfmntHyY4PEQ5ff7mAPpo+tKivBEfjd9axG
HiuwGibi9qLF3wAM7Cu6R0mez59VP075+mVwd55Xg6aZptGMp6msovelt090kDj4
NxeAKsFYvAaG7s4E1e+qcjlPtCtrti2NILoFTOp28OUcMyDo8L0uI1UPaNrNj4CM
G6JwGfRazOZY6XUSTy3AwPTatJ/0ywdXd3OJeDn9fChBgwsQsC4pYoH5K6S4XRzx
gSNED1eBvKkV5LwYPoDwApax7KgWscOMxTLe05bckXQ6Ya/cOmYFxnkX/lZd1GFW
ORNbZMlKqBCvmssK+fWbnmFJnv9vcrqJyRY2cMpwWcUzIX6KC9zKnEfpNLQx1494
diDorzkvJTLMEdRiUlsWMsYFBHJrDGkEtyowBfh2ldXGyqUZRodzIzD9JVvg6t7a
/5PkMa20qoDU5ynAEozGd3dHT0FRrNpl0e2nuCcsoAnBEr9aGqxGSTVzVl3c3XsC
KC4Ik37eFmFljHQl1G3EO3HS/3wdUeKMOXzNAzhTUyPtBlyHRvwPairy+vFQlaGT
2sBGCDmwpImE8aHp6gPGl94KfSNaJdUH4Pew2dQxACE3yW3Ck6XLT/PTe5FYZ4XA
L0mle4TDlU3gn1CsLJJwrmYiw69TAvKdYiq94gZOkzfH4U9f4Il7rP6Xj0mUMqHj
dgYuRxxhyG0Io7hFEjrfjGs5GZ+eyq5nzHkJZ2HqRoLAYCJXnKEY7lRJcjJdVEEB
iyl57Wx1cHLWahuYPHhfwieJwZBWxqhBJw/gokJrTNYoyfCPJ2gsYbbj/K5VSAa4
O+LGb5+mY5FguLsPAXmXbzyhhI6JMVYLryrIe3vMdMZ9e3EQFWq8S6t5djnCAF9A
2CgQIm/1dGSmCfq2lhNNrnUPsNoRqgrFMVCiY+zLlxdpksdFGcYebZPcN85rDpBP
WwSyiJB7yqW4zpZOez1RNEVxd/xoBJFofrMjZwhtTxicbQhfO/uM3kvqotecs4al
GatZgi5thZ7FuNh447XjwpnknUNPNLLfpCZBx9qoepka8GhPrFX1+ioIdiDzFHES
l2J2/3ARm86emD6U9qAQJwGtOtdNWbZi3Hcn8k2iGnunFSjRLN7rdfTpLxynHJpq
d77yOPbnQKupmKlZrrDmIWWZs1PvMGiPXAzTgagwP9fLQO6qFjG9pGfECl3OA1hA
QZFZ5O316XQr3XNmAsxEvGPDgXISUPuybAYIEMBrPeRNq3OkCU4mfkIoDV7kKWo8
5sxMolBxRu4zremmA9ucN7utZe125+jOk1wyYnr7Iow2nCJqa7CR+QwYVydSv+A6
1qXJgtB8GPaoV+IwJk20AMf9LMYigdZZ+Ql11/zr7GFnA4eqNk97nQWHMOo4h5by
121y0IkOxntgNvDFKpW+hkAVcbaaI+nczA7H0XZTZ1Q8K+Y7Lskpi+4X/qFucjqf
C1RVt9r8TXtnWf+GP99MamyR3dzOCDtR7OmmGXBD3ND/AfDPqRYz1R+S9g1UO8J1
7AL5wSrno2oceIAd17u3Vo18pEona2jopJxOurmnCjye3JFaMaIvqOGFlv98kyIT
ZWoAPUWZ+fH6+g/NET7p5LN7Z8tPRDNJGCM4NeWk2xvDfOP/tqVIRpIj/LqTjiOt
xhTFkn1koOUZLfk087nCehjVmAc1BE/Y25Aap5ve93yhJUlbb0wjq4m/2FSO/dLo
PAFnUuib+T1kcht2h1LxmUnc1pdgzHkQHhmokWaOAAI2lYjTNJ4U3xsVZweeQNdn
IpX8zicNRSphtODDs8gr4lMfchZjQOhyDZHlSSOvumYwVQYxV08vcZ8EiE4n2UlJ
fASfbAfXqbCICctVcC443C9d4ShM6yekDPtcXgNrnziJlaST1cKyjAfTkuqASyYr
Ma+pb1s604FVwc9WACs1xs4t1hRX7ISj/3M1oe0cv50yPecWxOyZK5TScENZB0NG
82NfLCnI1opDchrEJ3wboSQ24QJnPtxdBEGfxafGyYZLmhEVFoNCavYaRYVbNrkX
JJozQgqIft5lKCpfY2iVyjKvHCJ6gwADVnOhs2AVaH7gyoR9Geqv5kUChYnMeoeq
pKRefFxKmBt4L227j4KozMznfTgfJraLcByylaf+uOKJ4NCiAfYrCTDXZo+k9Iza
DetCYCyjFmwxhlccKNshb8wY6tKncxn+bKoAVwvXb2ldoN89CXx9khtQX/jqW5uO
6rXIPP6rck/J5uEYEyGOw4A6/udGMhw+8EJnZV4scZUm6khwRwhYTWSlydMkBLNd
OQG8tIdmPc9MW3p/pCRyJf/W1vVTY5OrDt+POxs1NIwjI0L3FoVvsocIkvFOIj8q
Hd79Yo3dATpe3aaalpNWR8aAS4XpqheC8fMceYxM6yitxumGygGl5+wtuqXy+0EC
vZta823fSSmPoaHZYYStP2B6QPr78EPe4Q7EIsfgvpFgoFvgym5aW8Kbuw43hptG
a51G7BYR1+FG+M971kvYHH4TmVL+BSy8H+Y40NuTFoYTmB+mHTb6EBMZB47WeOl5
1tfjoxlh5HdZhFSkw1UbxjNOMHg8CA69hhLjsrj63RhAKmOkTYE1b+dCPbhDkiJ8
czdkpXkj999VE11rV34CuuVoB6F6WIphp8jncZ3guiQUa9T6ft9rVsDsfQttUHjk
Eu8OiO/+znI5LPb0qWLK0ZI23auSjerG1uPnvjC+vFvYmgyJmxG/qFvklhUxLq+3
sp9xwRC80VykqPFsattZJAUX5G7Z9gtBJL0dSAYokHDG7OAoc+s192kZz7dyrJbT
P+Dh7o3bpCGjIfdWZlWBs7LKHB7t7biZLJNk68CXiWQm5u27YdsDKyaASrIT1uJa
eKYW9uiILJsce/RXJ8fgdfDAq+YnBNnT8Fr1qhGbzsutwlVLM2jJmjA8FM9bXaJV
4YXK5hBEliGxneCjvkA24RFYsUyAUe6mku7WBqkDUXgMTR3TdB+7cI3w3FpGvIA3
aGGu2h2WmP3x3J4EImMo4u+HnbhUCBOPZ7pRX+KGn4ReHR7oiDEpIWn3Vs6VytwZ
6PexBF9if/+QQ6RGpfMd4U9P9y2ZPuW/O7wMHikV9tJuTU70ghI2LnJwyglPvxJ/
ZRLMN70Q5NPkmiJLcSzkhQ19FGwZhQPTPAM9pq5ShjwgoizP9z3wXlc45PkMg4B0
SuYe5j+ejM4IXrl6mTfh0o+dvELkQNoyTWzzR0S30pAqs/irwTnBw/C89ZzGzByY
jPbb2wVWqyG68j4CE/Te756GyyntzgygUQbgcY54zKymJe033FZOx5bCwTPQQMtp
ChYxRnd3I8qFIq3O1MlDE7HTaWzOrzv93Vpk9+QR7QrffDA/MGjwBV2jz42aa6Nt
7IJOaOCd6vvTjexhahxUWuBKs20fdrKOMVqgPlYRUYb0F2BXMi6dmykY3tkwhqQA
KBgYE6vIKca7uLQcc1G6C+Q6E3XaplP6XG7mwp18l42wTIQLOMwQ0VsL81dkgvQd
yUXb3vLYslIDsZSK1Wg+eVbl3MGoNvncSF+DEVLU1U0Sl1UvbEESi8lvrJgQ0uZr
9VRCTw8Gqw2wk/lw/lBS5Xodjg0sG/UbGFN9/m4/kzhhGrSMnvqzb0dUzXF9webz
+1PdIRa6tphFFfDpV7pzPhuei86P58XSJ/cc6dz/HFp4ZDKr727X5qB3zJ3IOuP+
ot0Bpnl2WHLVcWBrEoF1l/pU6yR4RIC+33mxJ9mntlcWWiTGtYT1ouDgQK32fxWX
YAi20gqtUsW+xFerwkORyhcprU+Qhya6t6YPDc69/vgLcL3QPb+vlJJUY9QaT/Hj
DeUTuiUScUZPfdwKYjpKO0SKv1ffQmdWBmi2gcJ+zMa7FUyqciP+CWH+aGsobH0i
ZcwlPWs4XexcLJO6arJ+nvQxdrpl98G448VptNhDjuFm8Fvkn+sykQIxekFbRFtV
/Tu1j/DeUZiGeTSEVzCOtBwdu4FpGPKj+FBdPwC7RWz6O1syj8wUzRrJABfFv3Fn
qSf6KdlBHkHCxwyBP2+TztOz4BWRYG5Zbqto/ZWNsj3M1vbHH5ZZmvqvlelnCWue
YfuESlt+3vTvaLCBkwOPRMNcqF8bVZGx8LbJGcP2TbOWQINlkgxD3dCyWVlj8HBh
Zditx+t45B5Gg8l7rBvWH83zPcpn9tK56CVknmT07ME4PBLyHXIoWLJ8QJbxbfr8
FZ/iUhJ88pEJkFrWK7y+NbIWnQ7g4M1/GPEfekJs1iOsW/axT3XGnA1qwk4B1+Gh
O9q7LeuMZaTrrFL5xbGwMTBmnVv5yo2ltLyVceNKEkUXafL/HnFFWSriS/QnYYoR
xSPwJwxR1d0YdaR0NQe9lcfHrbtXrD4whQt9am43aP1ABbZCgArv+9Z/dhDncL8T
Z+tYhjN0sgZcGCggeIwL3gmSKxAfIXn2UQYWR74wUt6rMUuJfzO8k5L+bf0qttQS
/rEobhBtyElLsWRhI0VGUb/vPEUuwtBHHM/qCfIvk2C4l8UWA/JBcRvab/yDHBoT
JQtiT9gYhqBIsccvSJbMFnCjadSApaDzQSVHRmSR+Lypb6KQtcEBDP5Hr3fyvHHr
3uONDVt6lJP3CvQX9+ubKJ2qXnF/tFJw0uFHAUOjhE6GJF+pAtRHiIDyv3kbn4mj
3yIadk9R7gnZB0AqswxueWhvlXV5iMRfiaMLqgWzLy7Zm6OPj/0hX8nHYaiBHmIO
LqI7Rzrpg2r5doYiBXhq4QP8mKxRGfp+wS3N1kBDMhlHQo78Hv6+aKJ8yGuImwAp
RaXv/a2tcMb++MvUi+43rmCSELGTrtvznGmBbzGVTUHA3CmG1XUhqgynt0vrEPE4
TrkeDan0jrig1xo5pHWVg8jLFvBrGHSyD+EsKxpZ0ZYyf041aeNXhVBfOlWfrv7U
HwMdRTay91LBXeYY9Yv0IMrdVaVGOmSii3AjvrBGIz/S/IFOapv1EKyLJoHnBqEq
Wg+jhXSfObXAyZqFES2J8rDOZLr3sni/HMhQQYUgqDutZk2OtdY+h7mrLCox+4ZI
k+svgT3IV+P1wTztGBFfhPfflQTwb6Uh/jjsAFUZADyiGbuKkISC7nlA+en8Ozni
8pUAJGympBRwJMmsRwTxdcPEOdrlDHJ/PBdbAq5R2LoymBuMfavEzfm3YZxQFZYb
B891JkBHrJ5BZ2L5yaplQw==
`protect END_PROTECTED
