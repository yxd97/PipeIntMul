`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRSljtjahgGDTnwdLABYnSPIoePu8pxEb4lxpBPNwCdW4iSnj2fK8aZIZmzD+pHP
HpcWbzOa4Oeu0x96AmQYI4TRvJs/KJr7pTyuN/55aAiswaarw9SAzaHH0ka9iRHp
/Q3vPAaFNFG0SdxBz/xksIdt7xwwxmHsbk9gfO3UYjsvhKj1xYBMQmD9S0/NbKxK
izSD9RX0oPEjcNqGCORICYClANadkgzyg3qaC5lWyDbKJsDXpw/4mHJz7/D4A6oJ
Q1Zn7BNKMAjmZV9NnpMaa/eia2qtMjOJcddYO4pFP4T9mOnZO9RFYzALpHIpFfEd
4++k9+BfPyqVuahTx/JzJHsZZwEabzYIyZ9OpsF7t50qLH4IEA4XoYRF3QkhtB38
MkUlSHrfg2YKvFJEX5sqx2JMVoFpSlwdLvVkFTQ7y223kcpzCoIFD7QcIeaITb5p
NcaIvqZVhBZ84Bz62B9zO5TpGCA5eu0Dv81QdgJXQ17Psto5Q7p2qTwbhdLYqqFL
Xr6e80pookVa1J1IgVkd23rlHN6KvG7iq5H4M5zwyOc=
`protect END_PROTECTED
