`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIEJTjZGyVcF6dXBcj+HBkLliKSSFJbjpbrHhTwkG0YaDqMRv+8UGfbOlDR+a1t+
sFD4JnLw6i3yHaIJso6otb9cSGG3ZsDhnyM+eHKem4dI0GaVbk9Mr/hxNUhnfIYR
ET5S/EnCrWmhDI4Gkkegq9lHLV8+ep5uPWs9nQmOExbAZvpEk/Y808coZRUv96aF
tP02DOOwDceUqWahWYYjbSXfIhJErjhqfyv6p8P6tUg0vhrami9KmCVOkP/bHjav
+BK7D9g2gGnEmUpEdZtKAEwg5P7+/cyFS0ZCHQ3PCRSbIXTWLEGD5Zx4NUFt6Vop
ScDcomVSRKTKEHKuz0FN/gCoq+RAVKBDdGiGiuyQw770PB0+TIz9lWy9WUYRyGcU
9+7qWBlHjKkPn9dYqAfwBulHN+iHzkgs1VVDpquFyhbKl39vhFlNdy3Thxztzycb
uWEZH+2mDi772cmsHsXJMA==
`protect END_PROTECTED
