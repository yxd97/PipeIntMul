`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WAQ9spL6pZYJPWO8TEgJBzeLR9CqEYgWz95FEOVlvVL7B0h47vO5JIcV6aLCpaDi
FkZ0O7Uo9ii5aiLcU2kxn1sRqOq5cWqj8zzn04j7PenP4bhp417hZcrUdznyf0C9
6cOhCNF/otkx2HtgKDVxnXWfL1dfFC5lbbnFbt+ZLsXSb9RIOPmoHXS4R/LRNo1N
/kFU2oQ5KgbrX1e4pFls8pj/3D+ayQLeMAN8sQyzdvJ9Ca4Bnub/DvGxH4Y/CsPq
cFPV1RRiQheU3g7TlWfDmjuicZscZ5mQz17NXvZ02YWl/gCu/Jwsk3c0o5o8p9XG
wZPyGnqgSIi6O/kcDzezhJKcMf1GiVaE6I9qeP0E6Y7da4gnbE0zxw2mPtxuxIPz
gxFhvpBrGfJiJRkXU8mUvqPNFG+GyUpWf7w+/n3MWsIN7otl61wfuiKWVElCnrfw
PWsyz5/ScY4Y2NiVUKU1tg==
`protect END_PROTECTED
