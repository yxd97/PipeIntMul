`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tOWSfGn6iJiW1synBH9qHk8Mh1IsUxyXZCo1H3KRkKEOiDJjAkL37V5ARLbj93yU
6wTROf7Qt4XCjETSJDtN6ibYU4KlxYdyhO4YOEUQZIXcnoYKfx9RK1/NVFySbLdm
U2ltHrHVyL9QeDnjf8WKWRsuQ/jGzUQRF9CjQJP6e0IBX7OIOrEHFMruriWWT71g
s80tN4M+1qdkhKYQY9u19uSFFFh6cMsBGJWW3AbXI7oMRQRQQ+XI4Xtv8M1NHL5c
UxoMUJWW0WvHUabAQfDW9WSvgPc675hwTtDVAhWjbKLvbgVpFXLD7JdCkR8ZKVk5
9GuWMRJ3zTWmMJPXknFwrIV+47v1xSNSM2HR7DmcHZ29yvKm0HQzqDXiU8vhFGho
LS50v8ouKMJlO34JGEIgddQJ2f+5hrGLQqvOI/7awpwlqUHzc3BTXAm2UT0CKbYI
h6hMsEfl9gf2Ksi7bLu1WaIIGOStIcpW+7dCgWNRb/lz+z4qcnQ1G1POBKkJCRxS
NcqUIP0WKA29yQB2DLmdsmP7gjXr16eJCyyMZsPdHX9twlFBl4c9l81pop8+NoiP
wQgrjbAyJSCJoalKTWx8TpVnm6nT5MKmUOCQ4aGljxsNZ/SXt95sWZDh7Qpj+nOv
tCFu1IQ3ETXi8SDABuyNFIc2Eruf+W9Q7kG6Gb6+MVCXrmYW5yGbwTw70+IkVT+m
SpvlQpPRUcLjPfwOvCAs4s2gc5uokDe1U5iDSkvuVPaS0CAUMZjAYKerhkTJ3Piz
QEhjVCcV1jx6aYlD5x7dQCrbMBLz+tO8qaYiRxfcrabuVtFmnnCqoL/FTp5DYHta
RkVnSoMn279xT3hbWsQc/zZ6o+NdSFQnMRi7ttvAGon2mN7lrBlhaRv2mRnx9JYw
qGEho4WEZAM2zWbT9e1XxAQx6KF2oaI+NpWgVPWxdrb7A0O48WXoints0Ai/Ye+m
FhWAACDeqXo/SM3JXIoJZr9FDD4N9G+hdU64LnIVqRTnFs+Ix42WaBzpBJEPh9ay
`protect END_PROTECTED
