`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
egQbn3ErA54q8WEF6uNxr60VUYwGVg1eQjj3dQf1QdGGjaFOcBtj9/JJU6GgOtTH
BQKogpzdsbQypDbZT91xuBtVL4nDFYF6Pe/hBkArMDjUrT5W39BsM1EQJPi/8wwX
q6jgS7sk85ZAhc4/4U+KLZRX9tc6Vq7/eDcjcHbDMcS9+K7qPktbhBB2m5HYaSF2
2NjHIShXfkM+bwfLE/ZDptorC7nIRlhJZLi4LfGc8HZH/R3dFX2xejtNI3GbDgRT
2+rshctvqhd4JBGAiW6e0hhniYbpW2wp+Pwlh7T5w4hlRWKMBmIjYxYS2YFYINkZ
EMcjRI+7hPeXuWRXhBSjmPH+TjT2o0r0EXDSAxHcclNDB0jIShaI4O6dszvsMu8B
BFYHwHS6iA2J21bDL5um3bsua4RW0vJUG7mc4CJY/l2Vd3zCCvQV8wGfAxr/2dLx
QwXpwKAoeU4q6ktWpdWtNuRx9IeSAsfZ3DKNR/xAyhhEO/4PxV8x5PFiMRwlgF1I
Zh+HJ/JtrLeLAUIqsmq16nMqoHMZiRJmHcd4ReWLn3yvEMgrxw5WmkA7lFyD8Xu7
nsswb965t8sjx4mYxg16kRneq2+5gzhWCjQV4UeKWnPlA7UXoZi8tMpqY7XsGwPA
L0WXe2t98W3UZ3/RS0F3jw==
`protect END_PROTECTED
