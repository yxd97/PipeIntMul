`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6QEL5oaM8Pw3qUmXQ7hYIdz539NLdKntdkxMJYXfEmIP+szKgm09UuF6z4xoWfvk
Hz/0krRIS1OdPMU79nKkpc7vdjptD4mOGbtZhL8B5m2jPTDnot8em8MtOs9CSdru
xJEecn6xwFhZN3QLFYD4quwBpKhv+FYS97Kw9qxhXdm8J0Un6Ia05hvK0LUih098
bb+13ZYkxN0IVmLgkHZ/C9iJQhTh259jvWJ6+PGRYi0KlDqzheQyTFPDaUG5KtMo
5+0bO6sdUZEz+gtjkpe6JWRMkZ5dXnqVrBy40/spUUr1HwR9keaqfs0TK0ZRHhJw
nJj0/b4QL2N6OQBYj7xo5j52v1mF3tbT/f9dp+o+3gNMNsJg+yMwDsUDQRMQ3Sha
rNUWHx0Qi9frSBoyCjOVVcp3c77BJ8qTJjWfYsNvoPYF9i/LW9UpTbt5K9sgr2mc
fU+iSx14PdX/lA4OGJ83+w==
`protect END_PROTECTED
