`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VN/KGOluINNv4zrzDg7oWYEUQabVxwRjNK6BAjg3U9OXe0DD9qm6HThxSNnk+LsN
AKCBKtN41DMJKwsaPe03+qKLczoedtfi+E9h0fX4pRtsd1Hds7DO9S4DSKyRLYdm
n6QHlcJxrH2xG59y5jkz6nSizFKbnAMrkhtbODDPzZfAz63zup8NzMCgbvYApvMW
hhO7tBkYixxzqMyi0gon+NBk9USIF7x3MyA6wOWzlslfF7jOp0F812mWgGvsWTdm
8kDeiHyZFCoyMJtOMAx/B2exDoK3tJADasq9clwedQ3jWp48YI0QW1RQXztxu7nV
8ouTEKTjoDDFauvfczSXb4kA+Mgtkz+N2RnHwnFk/coIY/yfRchSX2eVqVZHQId6
5dCNz+LqsEEWXQelwvCuGdVrYN5W1qwqfA5vmvwHtMTQ/Ab/9wDPvPV+SEmpmXmz
8j6zxEvjlRDjnJa9kVxzZCb1joUL7mKf6P4vqUQ4Vpondkt7VYGWNmJOdrob0upA
GyAfkrFWTwK6Ujf9B4N1ZJcmx2baBoSJgJ9+8AXiQyE9Bg+TVBb2/Snh8NNggQp/
prEt9E14Shu0d4Xvdwjq2hFMNq7D62momyBjd+AQY9/pJMYdOj+AtxCkChAopsHJ
/DE6llnPCCyuwh6u30rXvFPJqXlZCa7w9vSHsJN7hIQdVefd6WeE+Sb8Ozw7C8Dp
Ab57dRYlhHo7OuBz7d6jan2+DbwiXE4jsFcxplw3YXuhjTe0NGSeh4in30qJNWS8
0sVphM4EdVOGCsMLFJr4luWIgiB+Hs6IE2ME5xaIVILWOE1ab1ehXF+MAYWVJ5t0
DI9W9qvK2yNv2Dg12QJ/R/W0Z+rf20DQXKebf4+NQ9284wGHNb198AIuJK/EQ6Up
WLfRKsRhNfCS07GL8jxw5Fg7x7d9/FkLm8e5GV4EXiCeCYytYSMtmiPWToKqLwfN
NJLgKy+EqrQ8ZSwWkS7c8x4w1r+g/wdN+0dunyWRL+U6cRhv00IaaMUM9B05eWTm
ARoUBK978hPvgPCGwlBz3eLR2dTVBgGOYdQHZRhX7KvHi0FaB6kDhDjokDVCaDRk
DeoGfa7iAiKgaRNa6XgCDxYurgmtDSgrsd1bY8gKBGxfyVfDXqowh6D8xAp9vwP5
6RktDKCK83E16imK2DGDNvq3S4YTTZrCYg8jU/f1PFCp3DsZUFULhYFNpdbfV47r
3e3LcN+K7WDyJrU4/e+dcCwNxliHnehKteyXE7z6D2M4Fvn7YUrYJkGfi9NuyJvl
qoF2Ib1tcmfjJKjvAFYqXk8CQ3At/OpGDqP7LGuoC/CtxYzhJ/c9OUHGRaWZoXqm
IXfbU6QFKtXZdT1PiBBNjglMt/ijo5jaEe/r6C4cA/7pcx2/E2wwbSsX311D21zO
JBsy6EkIWXnATZRwCp6sa1fPeKDGfoYD30i4+QZs+8J80Nc+9Q7GSG6lF1heR5v3
FTBmjFl+KDUMI3hYTWzs3vlb7mcPup8YR4PKXlNmcs0oLpyFuPCiglm4fJvosOjB
3P2YncdpP8jrOw+RaTMueQvyVxdPyYjggDrOjlQuAhfvnq+DgretFMVq1YHgDcpt
mWvzFjz3VdHnnt+wrNHMJasovKsrkcOlvMec05Yg+80eIGBc9GSAMLRNM0EFjB6v
aXyj/VGXEzJCGq5DNZi/63vtOrCusHjJ5VLnx2I4h7TwdSBf/jCkXBJFJkN7/W1a
RadYL6qrIfJTE6f+Ck3JN/c/u0ppuWinHuobnK5Xiq6k4triGa0/niMP8gu0C473
JGSkX7A93oUwgPMNusJO7x5LSE467cLTTaCPqEmXaS6XT4ME8bJ4n9eDk3pJnlCb
wQqGxWE+pjjh50AnVQ43diJb4JQwj6fobho7v9bE4Amhp825YOEC4X6eJsM85Zau
wah1lUNoZByxCpSfuUBfm5hbeqT6ataQmU3A7jDOwf/AAXzyTOgW2Fz9xjO114xs
+sot79Gto1WpG92fDtuHcsf6UqmP2fiuekZDp2fJns+o3G1i1EmoJujf6VE5WsVP
JM8WWOXmFRj2PS1Qg+Q2R4Vh4290gHuEtabMh+RArWBFxm607tLTn3xlWS5fRQS4
uyW6EtxGpP2gJHo9l/X8qF2UyfapHo9nL0scLpmpbaEuB+o2Fo13GF+oCmoXZ44c
TiPpteVHV6qgNgRzV6sXYq0eMHsu3odcfmO6IMJEPkPVYzSU6LojPv/wgZ3qjCnX
sVT321ZikweLAlh3OPZfB284dqIJaBqpNTkUk/yaDerEnxbT0YtBwy8XDeDSSdPG
CoKbTRiEebB7W67Fxo1loG0pWrQ+M8yI34cUuzUpZ85GydPNIVD3VA1PvfGoLqd3
kZhPGk8SBRTd+Si/sPPGrW8maSMWp2C9u+eURyuNi2uwqNwkfV5K85X1aZev2rAE
SJhy/LoEolamACgvjeK65YGDTh5hDR/frBI4/RAoxRhOY4FE6ucxRbzDWTyCX8ke
`protect END_PROTECTED
