`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBO5uStbUoKdFoCbA2Q5XPT6H08YSXcmcX1Pgc7S7EWdRGMEv+YnPF5IxS1aBEUU
bqvjPuQvyrsApWW3/qIes8TR4rtFsY0u3rlwr5SZyGyRwd9/VysJd8Bux4rrfS4K
p6MwaC/K2gt0aUzbtdek3fItqsPTeeAIKkPUJcR0l4m1F0xabHyA++h6QfnZrDQ1
dtO+MlVyKqx/gzB0xOi6hcqiPfKbZK6jUC/r7wmY8PPTa7yWYRcPf3Iwvwq1Pfz2
D7X2qbH/U7ykDqOefAb2uhhFwqnxYfL9yA1NpYe1qU2LQub8muipgXpRM5g05usE
jZV7LwGwuFBW4WSZRFSJyrSVb4o0g/KTpiA7Hy2AfhutR9faFH5uX2ZilVIhOZlr
HmPNnrNU66DlKKRAO/4zK+ixEMana5VXTj3Cm6MPZavCfWg+T68PNXbWXkNww25z
`protect END_PROTECTED
