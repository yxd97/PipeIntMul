`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I8Q4Cvh1CqNHARIFUaPN9L4SKgkZ59RmiDdlhj/QqADKMeLBIQl/4iwHAoNaoFuF
9ZCNbSWBuzs0FvZUfKg+AKDVeZp8cCjeKM8R1+USTKiR8v7VXhkuvhIoCPNtPIG7
MVTnfIWehCJ42kLemk+kUOns20pTxteRv2G/xsIzZi6w3zFHcldGKWaoVQQBGsQr
Ei/raRMTHYNYDH36KaYMA8EQWvTB+ig23GKvs4mdgflj9rcJMXK7ZbIpXkx0H7+B
q+Zx5GmsPArjVQCfBluZX8SSbN8ylCRi55UcrbzfI0tpHFqr3yxbaXZA8QlkK64Q
WhHtAHjdh1ON51CPCucb24PDXN7RZE7GYphakBoQ8WtqjrSHe+54F3yUtZ/LzKGQ
GYkE27PosrlR0HSZPJi/LPsuK6cZ1NrWq4wwuivawjmlEgxffG6tdIMtMwJqHh6v
joP7VVVPC293L5F1Mn0tf0h6yl/vTeZ/fI4kq6n6yvUuQGb9VYMkf3tlu2TMT2Zq
`protect END_PROTECTED
