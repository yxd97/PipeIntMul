`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+noPZiczuDVxlXey29fl3BOQL8JWy/jdxq6FSKKPXVGDPvSWO5vIeAakGMk+Gh8s
AxObHXWAmGJ9dNe+Yx/Vq2QUkvVyH69Ai71Md+9KG9H9XQ2CZJ+Xm6lrcJ15WPkt
DUKJhoVdldg1DcBomWrSJUx6fa2JHhm4m/evbk+lwposWSksXge9rJOE0Tj5d6cQ
HFekVbxRZC0BRb/BigjlDTmSv2NWEBVpGhuy4Q9RWffxXb84vpLm6xhmTs0I8vHu
/Mfu3N3LdMUkJYQ7voc9MaNX+NvwyWDvsLQzQGinc/Ge5Lcq118fPZFnK+gPTjwX
3XcDZA3h1F5xdsiXjUjr9FAZzBaM0t/sy2aBGtPax0SM6K0b6l2IIwThqrttYQpn
TFBjsjX3mXP2MU9wSxCrHQ9TNrBe9nON5M2mrLwv1PTU8KfAmlhpci7ds7k1prf4
/BMeLjB7V9f93zGNvNZnCqfs/nVVWmCygema49VNPmcWRc3i9O3il9xMzLCMrbyK
Z7mTyXnl/J4pGT/H/wuq9mjc6eVI34Sy1z3chT3nYPwbNMwPsIaj4korvuWl36ES
yv27ClDMGGIsPk581X/3KT+lZpqxbzfSKydkOZNLSxzv7YVyo0bZjkuZBtxRwya+
yZznYl2e9s+jxoLIn6whr1pEYGGxdYNyapaMok0d4kX8xwsLhNQ4UXNDlE6YPR6m
CTHXnwrZjFo+Le9cKsgAohvy752JBbSvgh77oZIHWPY=
`protect END_PROTECTED
