`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzzAzMw36GnaPcPbw0nq5pCYMNPDzMEKawKI+cLQNy3SOuQd6l8v8qIM7UdM3clu
rTAHMgKq+Z8AZl26WbmeND5k+lSNeJBE9Y6QT/dNm1zJTo5+tFphqbpVGeeO+K/0
kxLreL45yyCfs3rRbUd838M0lBt+hG0bnD9Qph9DYebgLNnO60ulv9u/amvF0Fiq
S8ojQbJ2O0ziNvsWRkJH8mLgDxUBcbis1g9msf+vpqqsj29WpVLaOY4sm78sZ79I
erQF+eRLcdX7iimlOUaQwDkA9TzR2HgUDQwd5jXPzfolDwok9wkb5Cz9Mhm0ZvAT
UnikfEy3dMBfUfbtDqVkL1y07gewE8EnbtVB/RSVCt6514TQZ1xjQV4p5W3eAofG
pqzWht/x6oE0wb5U6+94YVkkAngaFu9XKl731sewvLC5z5mWzQKmbP1B1yTj40iB
shfHry9QgsR4Nuc4XqWJIX3ZVA4JaUQevwlwSZT0sThHc6731IfNyv3HTmvqXhFv
HGgYN+ovbCf5lypf9DokhbAjtA67DqSvd2x63Jt60TExx75ntZhfXJApnNOWHk7J
Ym8T/G/V2JnE4vwNdtDzyFao4PpcQs9Sfg8hKb7B85mLY/8sPhkSY+xxw38mt55f
Fd0W4NtpW6SQ+NP3xtF61Xx1cWtpdw8FEQiofsmNdcrw1OJ35aC9tH9UXOw9Nik1
N7Z0RDLiB0lgIt/58uuGpiid+IvJMDMDGnFVJQ/UEMm3vxbxsm4q464rlnesYqAJ
Q6ThHtUcd96vCPKQDctmBH/9G7YXvxauTqropibWO+oH+iJP6YUT8W8Pn0gtSAPD
aeut97DjqzXmMOjPk4p8iqtT4enjEe2vQK1W5alxRcRSfZtjEueuU1dWjfRbdo3m
7IFo6u5d6D5U58kMz0tGp8SArnWaSmEc0kIIBo6xnKeyOpaDHYVxeqh9x7W/t3lr
7jHkrMsFCmOQ+jJZZiYCRA==
`protect END_PROTECTED
