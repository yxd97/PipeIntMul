`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f0u6TOO2D2QMK5zGAyX4gX7y/g/fyJ8pF33hTsjtcLJrVyDQp2cTDYWFLE1jh8zf
KMohhmm/Yk9l9xdsXPR0Fd2Pyo6uMpioidz2nuTVwIroUk8LF0PB4K2y0tuttb/B
AX0XtjyPDmm3/OgwkjIUXESBF2R9teks9CIpaq6ehkYwUvvmaMCKdrAnhCx+qHC3
fID7SViGd1397cY9B//T2xan4ZJNJhX1zUPsCsvxb9TNsTVSrGCqV7mnhtmgfXLR
`protect END_PROTECTED
