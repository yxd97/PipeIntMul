`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTb+En8QSYTHqmU4sFr65Jt+0RCzlZNeWP8iqYiHMPPoqc6gfzOzjREonjcgCjUb
nRKoGd1QGwCVpEZe12GxMrYmLmxazdF1e7tienRqKhRBM/yuQNPtwTVnfDP5o1CF
P3ziNz3DUVjVM6AKZiWLJH1seQRuzF7wL2IdsUhqzwHuYcWTjfZXsEWkozuoNn7T
9p9GeXuvhH1yXHtXDXc5u3kVboHbAKzoe5IkAVBYfHwNYtHWcfqE+2Z8zWFbw76m
QoJzHJtYAC8qz/XtsXlF8Ok2kHUhGK7C0YXip+OMlCvGC12m0SMKsMHfelGacfWM
XOaPhRVAOyKPOuNphE/yPw==
`protect END_PROTECTED
