`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
elGhd5EjVIAs70DCps/R55CQgvPCOhvqH7U0BZJ/kebh58U2DjtaQofTh+8BW4bx
Y+65wHLbkOP+4I2mi5h1gYEDVcmjItrk+E7tGeFjqGbAjTGPRrWOnTB4+DsYuHpo
JmOxM60jStVqzQj3foCO08PyMz0KZSG20oes+N7F4PiKnuq3DFerGwWLq6aSiknh
uKXsYbVKWVRTQW8x3y7pUsMtArW186O536nJAKkDHXu6Wr7r3QEUsQyBTG+pMODE
/LSvTGRM956a0mhlsGkuzHXKZYbLvflQEnTRW5zx8UNd4PrkywxkB+s4KXsgrW3B
sJIbcpsGHLml82zrhax+XZ9yZ2vs/+5HQXbpT2fhD/LTCkUzgNnFaZiNLqMml2op
ro5mwvUVWYk/i1GQUofZ0L5nRX57ZnAy+HZxwR1dIb0RyXVtkLBekwXqoq+geV95
ATIftFvTEulfuq8NSipfAC/af5HnlrJarBh43DbyaPe0czGr7veLLV+TJvdaIc8Y
R/E79P9uo6cCJRolwvkSuZo+hfvM1ZqwBBZnkUrvo1xv7zbBTvVZ80g2PAKDCpk9
Me2JpoxFtQ4YV6stLa1lf3NfGsqTfQHbZaxCLCGIqRIKzu5vLuulT/IqjoJRkQmL
Fdqgy2Bpozu1OCotRByVyg==
`protect END_PROTECTED
