`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xiomakFDzU9AKKHax3prPDD0xcJOp3LlvyLAjRkuB8j68IhMQ8jZRlX+W874AoVS
s7nVNA8cblWfEdHqSoLw7XO4Q3o0UJeN4OSpLBDp+2io0CgLkeEQUFuBV9Xwuhdg
jh3yz0U/dhQfBzvJbW41J35XQJhmxG1aPTC4Fxvd81ikW9qMjCJ5B6O5GgLPzN1v
1++mxGm/EHlcBqgdz+ZCMPwJlMXQ/xPT+NCe+F9MPjFhhAS3RTDnbkUgnPJFlGvA
mQj9Ut+8ieLBWm84wg/fxD6lzoOFYBOdwMdmeHdPV0llAPhNIG3p4gI0OUS7GWJi
gxtuFNDCIOsUQTbV0ZTTx4fzVdWKJ4+/xES3VUgikkILIg+3Th6dkm8kr9VcPYft
57dHYhNx5cHVCjjSS0sfeQE7+9JYOH7Go2pNF2g5Pakcfw76jvBfXxzqN+RkOKGp
YL167VsQQc5cDUtRYfUHvfDjnWddFVY7nUVmzfWj+7Y4tBpJocRQy0b9zv9rd85H
8NNprEP3GhMQCoHeTCs++MAFr5T1socnRWGZZA6VvUM4BRuPLkqWsMTIhXkGMykt
yHq5cizATCv7RpFojzFMGga0XvqLYuWn9sJMloxHqFJN2PquaXqcmAuDj+8RV6ZS
d4gH0MfvIuNI6IsibxZZdnHo5p/UpFIn87XmCZEwU4/AP9e6kaTC77CBQLi8CBda
2goqteAhvG363akXHrCur+5IkvWunX1/RQdjxsbOzyGwoZh0Y7YyvcvuoDSLIdcK
Kx2/maSL8oQCzhzd80eHKigfZbWhNbi7Ft/ELt4iU8yFeKV3NG2+Wk3ueBsUT9B0
h34a73bvjUcvaeo4n2VBgu5/GjicvU5T4BYLSqnjymKFC34BpPO41DYIMJbxD6+9
5DxcUkSK0v6UQ3Dn67BetX/12kq/yBKsunvarhxlRbA29gZQRjcZwGrFK4rHADMT
U4WOi1afQaEGXN9cqVDMTe+hbVeJFRFzEeamMpq1QpTUshH0+VOpliAgBf+yAj3a
IaDK7AEsjP9wE77NAE+prpTJhaRBznguuDxTQPIDCgZT3iWEVKb3Qm0XDxk9ZPvd
RCJVs3S0IDnM3YMuJwklX3QyUxHhpd8zv8kWrGYgUst4jDZqJLPTE5tsFeiOmY5U
NHcF/zNqFHrHAc2e6xRxVXx1bL4hJzxMWXGoYTuDVzEQ0vA29ipsUwpuYxW3A8Zb
3pymn9giqJ8UDoDDx2WJA3OixPFdbfJwUJIDSg5aYy/pYRqrguSKje8SIFc7rWOC
a6C6ctMYMOCA1mYrkTjH+HXODp7FmV9y19HjYhsVWywH9JYmtRmmtyDsLoFy73HD
AF9QxSjafay2iBevQMiK9pqxycW/FFV15mTu/MoVRYkk3Jy5sbgiW5cP/a7nfVDj
lsHAVFek3KXJe4VJAuKP/DEvUcdMdAwa07dY5xRXPgxkR9EGH47Er67yJbv3oRJz
uz97Cg5qKjwmmasrsqMVLDuPEduXrI2dArIQHbCQkP42uXN3WOxreVR1rsckUhfB
U/lp/0BdpfTrkFdTe1bE5FhiTT611kI0B+3un6dlX+G4bJK/fz4f98Ey6rAEbOKU
DeepxXXunSCSBo+kfX5fe1RFOe4+2L3+RMySSyNgMC30ZMUpOsh8b/OPUu5W23ts
wq3Oa1syd1fj+aMtZwy8lKQJ3T1YuRWNO0x681dJGhPLbuis/phRbStZAu7np9HK
9BlxQdItCbPR4Rj4kzQQy1QHnU1PclNJOOz68z5xmtePV9hBE45ZzXu2Bv1HwqUe
0aAHLxgTyIakRu0/Cw9e0ARooYdPObRQBi5LmtOzrBt9ejUFEPB9xhbW8HAQlpLQ
+ONPxVSZNznDJLV9PrC4KESc+Wrmd9/ofdSx7YdpdcWsQXclxQAEH1BFwNquDYjw
s0DVFliCyXLFnMTp+Wk+fiXF49Q6jIC56VxGZt53ae3Y41InAk3iNYYf5Bhv7QIY
b6j+Zn4VYciFvNkIFlUkMlItPwEyg+jLbhAuUg6UYcMiF1WebAEBwxs1BpheUcvT
FGeWHDp8QdUMDUSjKNFGK6ZBo2B+1Da4F1ouqHJisPs7AZj+TIwLrRu7zAaCpAoT
nUAclSbEWwKemjM2o9jOMyuNTojZcbXMJolznW2/DsUz1YdjxGGElfJWXl4U5uO5
RQ6jbX4EzR5+1lgAPfo8EVNWwRwOBZzVlT/HhC8aTwJZoBClz5SbGImlvb2ilEy+
96LDyqQlo2PUavRQ3GnEzap8/UHXCyNjgD3Xv00Okj5NQrvZpt32AK9z1A1tq3DZ
KApWkYd2sRl/KsYOfHJeSnsgoqI92R5MXyGEKC7pNOGh2f3gZvn51B/ft5JUTuR9
WV6NLTdWUO0KmbQG9daNw+1d6K7R4DMTD0h7z52epHMvs+i2NFJoWtnAKmDvyDZZ
6hxM32ZMfOXVqlHv21/9vfwjiWC9Ei2ty03ZBTfpX/ZqMirGhKmp7d2Kca8ckSO1
Paq9Wd7hoMSFBEGlJaaTzq0K/+9VDDLxqCcACCIIq1c=
`protect END_PROTECTED
