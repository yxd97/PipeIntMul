`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dU6914mL/mYzhSBofs8wBwqB5xmgRgUblTGRmVg/sudF1BxMznSd5mISX4D/ypY6
St4Nu+OMaLlqXKmAmgf7jxBM8oKyTS4eGWKucEg1bwluVSvzoA1Nt3wbIQNeGXPw
2ddtgXvD1Wf3tKN0RUvEIY/ffuK6y0PXifF+MiPMQNcs6FhrXL6s8eKqaXSlFFZA
km8v8WsKlNShSAx+1jPQDz901cTRYl5qXDdhIs4W+SOM4vgKc0worQ5lgg1NXfX4
s8NxAEjYpyTt4fUTVj91N/RenD4fRoT/OOmo7jRLqH2KjuRD19JS8Kui1+GnbxeW
pLJy0qpCSiLyBl33MW28dCdCOQaoQEGlyYASBP/mDUKveFYhJiAhWtZT4Ym8iWST
ahLG7CRlLgp9quCVdTngEeNKd6qJeH0tDr9xFmnBSzJs2CWilofNWzEm4JnXjZpB
QN5TCk1DNmpd233Drhdv9vSzgbfSMUN/5Mr2i0r2kdP3HPV9wC3qjGBgQqMRsh7c
a69F3Me+P+88bDeDCIqRjprevdmmB9dtRl3OInGP/3qJvwQwS2GtZQnFMYbOYMY3
jckAqjx3xgEiKnmuF9s6Toxk3n5WyQ+PMjz/LkXdJpNrbfhWMdO6Wo4hLfQPJUL8
sZbaa/XZ7AlsN6qYlQdSJPfCn8KRNDzx8s25jYrMQaENWgGR6K3qk7nM8KVsK7wv
E4DpYDMTEEBxcmkzK91eQSdAI/+KQnFKNI3kHs6rKzg1yXqcGxs4IGhFxWbyODa1
uDqpJeIBGdPHLBU0aE8xUA==
`protect END_PROTECTED
