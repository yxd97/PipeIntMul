`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TrQBjzQyin8yqmgzOa7IHu/3M9C4DXsS/1VCyljVbnNiwIFeHKn91kc7eWyFj6at
ZH/VE0o2/YiafcF2RPoU+7tFKdnrCqEIxmXi1NlGEsMZ8lH749HCDD9105wiAfPe
S5OtCx3eP7QXOI0cSRTb69SR9SfX7jdm3Twk40TjnS0T2CI7xgiYf1KYQADhSrnq
v41kvzkXMoZ6YI7M3ETlWN6hZVPSqKASywS8yLzNvTUu14fvFlu/bigkbwXuQL+E
+8B8HcX3/OuFQYvxexizQ8+Q1tcCzoSPSaHLnKiIW87Zb7WW0m6YG6ch63sqywfs
pE43XLdSI55hfM+sSOovJyWDSbPJrMo0CPC+7t52qclagnjWAAiEI65LUwUDs6qu
usHvJ8gLFqdVerxx4amsY3j5VItcOolrTBjWT4b5lUFPTx4vCW5Y/mM0XWqHYXiI
LbD5qBW4YyGFqJUOr0uORVEA0nm4QOp6FFnXVS2RkbnKFqWqjahy4Vpcqa7H9k5d
6gj57/xdy9OFjhH91Nr6uKRHJEMOum3OJ+5MQMQTUmxMAlLq0ZR6rtr39vB16rJc
QAON272A8q+99vN7U9uFrc0JvlJ5PLux3lxozypYX/zSUKec/IHGiBgcvhO0Jizr
7t9cbcEmeow1z1MYQSplwCa6W6WiLIOre3LK5Hfqb8A=
`protect END_PROTECTED
