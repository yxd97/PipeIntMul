`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pkr4ZobiW/mK/ffFeeR5oHZn45lGDDF+HVmGgteKeg/WeUF0zAByT0I2Gu0/IKVa
1R4YaRAWd/QWIRUb22GzTBdufsLNIX3nHKNShMe+mua3ByJhnz6zjY1aWB8zcK9S
QCV90/7vZ/go0Yte2ZG5ris4p7jrB4Jr1UxgZ3gCxWBVco4logRe+U0aPPasb2s6
+MIspOniAMTFiG9Ve/ETEtT8/8IXWPhsRjd805Dl0FhwJ3ZjQpsYiFPKWDR5fdCn
6Kg6xgH27qfSOWhDjupLpD98kQHIXnaEh9koFUnqIJ5tBFaFOWOpy/hrYvZGHqb4
GzwCUJI/o9DD4Ch755MF06wwIi+70GFycsAe5eQQ/DTHxQL2P1YKTlfbWL/o99W/
NPdTAx7xCsyznsq9RA0qlcrMq5N/jbGao2cmDXkCZfyIKXamr9RgFAEbaNPmeHy7
`protect END_PROTECTED
