`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BKnKhPUA7YLfVMNIbd6CojtlAXHLaIPm9dFxZcZGhycIzrFMQFIKYs8ujIYoDKBR
sGukO1X5tUIfu24QTC6Fk4KZrJfSupjoTNH9kE1JW6PXeKON9T328hU8M+fnxhc+
j8Y6Ekz25gpp0wdTjkW+3MdomEFCdQZsGpkDiDth9f+OaEAaxHu6enb3TJmU0D6X
cSD01SCncCHRaDuG4QgKBQn+0l8gRPl+AWsSD9b6f5495jc81p9s7aOtP/WdCqUF
SavFKKN+7CFlA05bVrKjtmdeCjcQ32EEHltnMAtQqVDHJjnJyB2u9/6r24FwFScA
+o8fqMiv4PmnyDqPM4XWBDvRB57BiCj7W8kwx+ku5eWRESQRt43i8dgzxDRSgLFf
5WoX+Ks+K45grbIbcIXEWsN8CDsPJB1vA/ODYbIfkv4+tJZ9Ew9cAlFq6V5hfvYV
WMW29PbYlSkRVw1xGUDJvoUSvCmkhzZx1xtntNAJHQEZ37xmzBfa/bUlM4eq77UP
D0fUZ2Z+qlULn3IEPf/Hc3LTa7eGrQ32uzPDRs977mwxQjTc29WQ9zXfvmm5v0x2
+fb1b8OLuOSftKZLAl9rdkRwgsvvvd1pRt/3FW8jQ9SOaUt+yDe7zZ591ZIW2k1C
sKIYJuzqFuArEo69zMuwLhU+OPpStXySLQfysReNLc/imW9sO8Rjz5B+BVlwZMQK
QH12AhTGLHg+mNRCCFkXA9MYd1sPwPr2oQD8Qb9UgNSZEhI2C1YqpWqzf71vONE+
/ZhqSqmvHhnY780xTC3eCEozdaxX4G0gbhihPOTqgbLb1Xgs4HT1qcNTx5RYABdr
oFWysxGNsK6YT4PeIwqGIkwecX9n9eKTpfnlBtRei7y2ByVS6271M6BKtcDwJGCk
n/DZzGzyKbhIRRO+jQ5PT1qRn0fFqAp1GYMjFYcFPu6FlTXjbZQ46BcvROQZHygf
/S+sX92brM1w/ir09A/6GR1YJkUsps8ksEhNY6ZCPxbS1HPQ26Irjh+BUuTP4Ejc
KzwHtR1Vakl+Xz1EbHien/6qSmO1d/i0B0VLRbCK7j8D3AXjhHGeY4Z0pYh8CIq7
1pkBO7sJRorOc73hTgZDu1umtA4/kGM3z4ySBqLAKL/+40l5N/qqMIDRA8sI/YXg
ldX+rd4v+pUYxa4R8HI9YxrfLim+a0g1sz4FS67fuTkrBsxVG/MTRBByja6TVThO
WbayOlnOnKWI+GbKDkq0lMBgH4yfUumveVDM9+2YGTyaFbRRYcoKMiwXtSgUWFXd
5kCsJJ4zsNE7NfZDybG2/isgZGEU7H4T0dFrG6a8rbU5MGc5eI8M7vq4rc+3Wil8
VylNkUG4N62j4DiiA2YLNN4tViNA5ow+Laak5TGADaOnJqFHcDla9yXLsyXtHvuK
cJ+uDksgclusB1BDAsvERCycYvgjy5OpxvUZPLGic8Q7tfaTs4MbAxWDR6A1VQ7h
I85MgQrNi0+tky6DMBYLOyh6BNAD1Rh5SWpaqqc/q6qXbcVWgrfDzIGtyvrIsCet
sq31B+JMGVd3dXo2hk9qSMLcvpSRclEPthB/Z2DHq/TP7Vd3RolrhukDrs/hlrVY
8yHTryvzZ2fl6K/Y+UMgY4vblqjnNxKHzjeXpoVJZcCIJSvXSDT7U5IJxqGjYe8X
SnINbUgst3tQmIJ7RB6/wxynJw+KSo9Y/1f+b4t29FL6FxYAN+IAd5XDngMbgQNb
z8zgTuS6Gh8QJUunT4oQIzW7lIVmU9QaohIJq/6E5vrSnPC9En1NmLTqLNgIYtDr
NGRTQk74rHb7hTuOI5W5I0y+3cLYve5vGjqOs9i4ccwhPcYYyDT9s+hbDjWZcSIM
ggUvlGXpGhPCd801/L9XpY4i4aJOEosiCN3JzQHUNYdjNY+fojkMUUgtJjcvChWC
qwPdi2ANqyvnWblgQng2O229V+4XSorq/YMA99ItgnNF7Y9t7Y32k+J5z2NWRSKf
kVKnZ1+02LnfsLc0HLnr2YN6InJM+asHebKzMzOwTpvk3PNiB9Y6rA2yuzKjVWRF
kALjfe2vc12iA8p+GDLPAAugZOf5VZrqG16ZIqJqOTHjUBTSbnTfFtmh442TFo5W
++Q3bQpsQWl9FgCMHFGRWN2XhmtqbDk0RSTPD0ZXlhzzWKnhnwDb8gwWgs/wreM8
0Ao9RGvNRO9qnQqZI4TlULkA43yjL0zGggWFASAe5dQlpIpkAO1kiZ2WdvgD38Ec
i7tXwEWQJHoXL30qBbbaSrzbIcwzZEVVv+8RNW6zO++YGC/NuRmQ2S5GP/d49nm+
wr8oIdqQGwRYAdQp2I2ZTbZa/br4RQkFGxXB9CFAd023fX4kRCfL1D9gbllCwrnf
oAlWQrDTDngnd1cv8/7JbPXD+gZc3ClEhMY1yINujbSMCQLHLRoAi+Bfu3DVyhEk
NBVYYrDS3mCWD60ik8+iK4IGLocJ2jWRlwsJaTcgBwCwmdau4oXa8yps0mWqaIuK
WBdEym/SG6CHMhDldV9YjG6cLWxGDpoV8Nr5GYHIp9fAoWi2xDSSxO21oLyCE/gX
rVgCSNP/7CGmv38wVZVikRKIRyODytw+b4d/hQC5FN2qcYjUJJ3SqGWZEaS9QjXl
8xMctnHY9lqe/PYs+Qox+9pTYUqlDmG8PP18IiXhxX2WS2dCY0pCp7OfN+5WUAy3
xcde/iO7QkYf44lWRhlbgHheqsHQ3lM1gn69bRw05f/gJ+lRuH7m9yuqD9rBN2Hr
ukWjWJQADLi4ep6oHy2wfB39TPpI1uW9tjEAJsZizgz8Mn6GKMsujyj3uxMPeMN3
OLhKP0HGBliewitO0FhuahEk25txQJuEgqkTgByfohW9S9geq/FiqaFH/w4A8m90
o10QrntI7e4UEziHHmKKYQmzdxeu4D2BzHTAh1t8DRf8qEE6ZG84Gr3/vu8R8F3R
d4HnOrheCJSNZzKAk8wzgj6T6hw8LcgsT7RfRH4b0F6sEMlh8gDwFlFRx4SJmSh9
jpX9XNGMDo9loaFzppVvPFl/vy3wu0dzUj9UzrD2w06OX5o1r5YDvFl8V12s4rYQ
4q0FfiNUGp5V9xegts1ofDPFWLU6eMsCimYbNcN/tM8wfSLq8FiQoLWs0r0A24r2
sJbWjRy2kur5AL1oyokqCPRBH2mNo6Ewhjuynen/ZgR8riTw4edxq0TDxVxdH5o9
InF/lHNZ0DlG6QWuZyIGidGYs8/yxWJD8ProeQUSKuM8h1okZNr7gWtcehcHuwES
AoEDXZJZC9WH3XDhEUFoNOCVTDcIQgGo/NYr5F2VdmlllppIf5CdgiRwWYy26ATd
4Cwc4m3tCzy0Q55VYmhe4yrKNSOChzi5xI9TZ4kpZkm7YsPvefXjO3nVRqM4Za5R
/IrJhKRHHB5TE2NRfxbYzkN2RASayKUnPiBb3TytMiyEKEg7bQWT6z+Dtgop1Yi1
azsvemrN/2BC1ix5KZ3DyGo2AgTCdewZG8ygXBECA7PjAa2oSCvThrium519sv7K
1J3q6BAn7NDsoA93kiZnpPQDk31l0I4w5agLYn/oKY0KgcgLxjXsODclT2q1YMNm
/j1zgMwWhY8EvczWT3hFqtTLilo31aY4UCjLzfjkqiD4PidQxfivGqWBztT0PiO0
Oi2XWzCefiFXxL3S3glyL6r4AnUmUe80t9JahhJGI0Q4XhxB1s5FC71uAJ75k7mS
W4t2jrmmV/hno0mptrXMcyHv+jpGy7imyoy7xPowzRZ2JHlQoxB6t3e1VF1tgE5E
RUJkpYYAHhRQeVkCOWWD3DUSy9hBt8XWWlwZKT7qXJBfRfEKBSL/fbJCCbOb+ADo
CE2UCPJRV8rRfGHHoqklb/9Z4XYmSLnzDf4W9Lmvr4VobbLo2mSZecZt1ms3PoDq
ojIPVwlo+HhppsH450wTQO/SXIvQVw2dg3caVBGWrs/gYNVonQoQVC+Ev/AXwRlV
DAnd0TL8oW1Z3ImAY2WMT5cvVGXoCSIUBkc5H9alnwAbIXO59JTaqW3XSX32O0Io
a6lHrhkusDoIRle32FmWIEmoXvuHsx1dn0golF6+mxeS5tp+MMc+So1AigwdoebW
3m8G+6rzZQRsdjiCN5tH27t5deA/IrWXBvKHoEmrOopmXvYEDJcoiZS9lv6cvS1i
g9wQwJmERTWfccBoa7lJvLYlCa6DiDWeFECvruD94fxtIMwMcBFV6O/2/0FYnWRW
XG3IYpDL5MpLgAcB8LfwhwmtZD2fXIf1D66BsoVmBbNHGV4nr6GxVF1Wsl8n3ZGd
RZQFRKiyobhDHFrJorO/eZT4MEv+dOL1WZsg/cOHw4cfSx97xHdxgIbkD3wUnmge
Rzu7mNSQUorWDaNYZuBGJ1Du+dcPt+jYaqFnJ3aSYVOvm3JjYxbE6XdE0XF/O5X6
76WJHLuPxIcg7Kxafk69QI5VRqg3T/XEnD1HUbdj11H5I45QGCj7tffilBviStCo
KxjLWD0KAKR9QkOk/Xzq2Gr8cGWiVtL18vxaAGxZNMopZTSGEr3yHseiTFwrTsK1
/Fbt/DkI8CSeWwkn35n3HTHA87NeynhcTE8XJery+Cra8XfiJFV6WLaKPIwsG/ur
osaE487yOOISuUKuBALQgX1EpK6Tzw5RqldB67vsAVwlCVrBT45g6z3Trn3OsATL
/Uun4gALOZd09O75/Xi7PlrlGC98Brgpr9nPQscjFy5tWt029hzErJCIvvC1+yje
4ahOdnfwmYKoI7JFz9U6bqrCic/Odn1kFY9QmkkfpxXsXMNfxLgYBXuoGD6FS8tt
bEDmrc/2QZEJIlenClaefhRtqUoJeZqL4zUTR5AM92kzR8UQJ1y6R5G9wsB+KLHF
BC56JAQn0X47S/K7pZEAeN+F31LkKqa2m4bRYlWyPY1YnxDZBLZXyM2Tjbl6uQF5
1YpupS5egyOmOJkW6QLf9aLigd8rUSJoSlAo7tbOQyWnw6QW4ZC2mpIypv7JE7jD
V/KDkyMWDmnvqPTIKWdpFLtjM3sSp0uNjCEmm/QonWsFiG+5uNTWQcYImBN1sGcb
7DFitqy7+Mw02ZsPfdDFpg/xChSXAYo6IbgddPcZafj0LqIqcSgHRjlKrw+6helc
Q5Z/Xe23oNZLrVnCtG9dkJ6yYvPdqH8Qx22fTeU4cAsQ1ib7IueXCaVRn9wHuEi6
vS51y/3OBZSx/BklWE/sxSX+Lx2waRtt+TPWE9GxaBFALM7zxNzJzc/rhQukvdFa
1eg43N40W4VkAnLrZ/mmCP9zd7L94Toh3wZjsINP4LBCDZKHzEY93VKEuXZOuac6
81v8vXRSWhqdeCcdCaYAwvwmSo3Cnim5Tokg/JBXQ3iKO7jWnJ9wTAveLeEa2kNK
Sz+bL4vX31KqadmBW1mYnELEJJlxYACw96EIO2A5XgYoaiR0NM87bKJlLiw2vm0D
nt9bHKeC4YuYfY+G079+rUrvNZky9eqlQrIssTCwJk2KVaiamPQDll8DHn42NgYc
ZD4vfuDaSYrqOMh+0hSLw/1cbdylpvWZteP40qhpB8Q8E9eFhIUhl3/bUQHBdcSn
Wp9MZw18ZQDPILEnBmMQ5zQZmVqu+PCBCqxqYkIZ8pRS5jv8UebZyXdXXcTnlRvu
c/6G4LXenUboxrvfy0dt6t6GsqbPJ5qGRnTT/mNBoz2y97kMYYltpOFFUpIKVOMt
r/mFUU9Dx2jNAXLNwMXWqDx1C/XiIOEQWEe8KTQoeisKCOeam6QXl6zyCb8tDFcg
WkcMji5hIpFMhn5Eqw8tkQCwciBRbe30DeZ+K6u91aNfCEGk9426XO/wahCmSUOp
vfSqAy4ZHnrB+VLOH+9eR1lCG/RgeRPE8vIrV3W5ZDrkpZrAqXwmLHxl+lyY6so1
u04jFDAVfSeigvcShclgnUoHBbXc5W99gMj9MmaI893zrR3rqBb28JA4YK7mmISS
K+QafxLMXtke3ik6IoJgdq4ZOHIjMgUct+8ym3oIQNXb2P4eC5xmxbcQq82QZ4Uj
cUh37HdiRrhWOZAxE0MQ0uUi4jHc01gyYb/vVEgIPTkTbj/xv32A0m3yaNf3JcZA
zXEfHNgu4i2xSES/ACGzJFDeRzwKUfPpHxxqXEUYtJbeG9LXBfPh5gmtjSlToOOc
kmlKd1NRp4zvx3//6aBpf6JpGSnb+PlMJ4tuNTlqnIaFL2DciXAogIRBaWMd0T2z
YKI2gggCf/CKCTCbK5u3J0FkFRVgJ7drpFEgZBm1wgyzqdeMC5MDMQ2GU21l3J61
Nyppv93oKGdK2Jc8OWsNrvcBknBjrUTmMTPJuZUYufj3yiSNyruhjWPOS1+uVTHl
Qqc6F5YBchQgXMhSrpVaWZoU4F4monAmP36lgLan0S2fp2Zs0RHVk6zdWHVSKDc5
33u0BH3QR09dd8eE2OMMQS5Tnm06ljUvj2raneZjAUq2vXMjD2aN+3vGrYKoN2lS
ZhV/y13JWxxaNrDx0/y1Qory4Wgo1ZE2wBK1Ih6+S3S2T3lBPqkiV0WTM0Oh2g8M
BojGfE6svvSKfkHMXyLcJezsnreyLtUo8iXu8Ex+CUfa3+Y5D4yUSIA7kHSV2ujV
TRccqi51hiPvkcexUqYjiQUVLRp2xTPKC/dMENBLcBlZhVkNUGPfxpndcz1ga0le
WVyzJLoeJB1XVOaBgkHX4j/Uzug4b2i9L09mKWxYeLvMvA/GByclIdeEn+hd//HO
FEPsX+OHAI//UyTC8sNgC4nswFoOGz3f42hqHwQjXfvDYXDiIrC6adO3VDecoP2F
ajlgX2icNn/khCLQ2uEo0Fq2nMz3f6EDCMnH0QBvgv/952UHgui3Ta4w6EixRhH2
GmSrwgiP8gKFaBXqWbMOpJ/hvMR7aTvE/SByDsBH81Lxq+My9OzQxb8h9gJEH2aa
N0uT2IgosOgdmPg+IAIX69w1v8w3iwVcxwM5+UfrB66wEnoz+TMis/3wZVg3//Hc
4zQip59fm4zNbMk1HqGwLKtBpp6PVC6lst6kUMAXtDT6aUCscjoojELP0TOm8i+T
xIMKvJC/p/m6erboIoM10aTdrICYX3awklW2BxzIPxgOBaAT3n570DhvUoQ8aqWa
H3D67omPZUlZr5ppMlZyAukWVT+o/DXky0CdyLMrD1WO4mb2DWJjnXY1lfLzhB1+
VJGoFBHRuohrghNc0WrXZ1zg0uso7PVgwSifEXZtvwLS3JA+hkPfPUxqMkPo4RKN
TpaamA94eCmorM0xRy4QuPC7VuA3VaEp1QU8eErZjLn0G53lxZ+yw+EH7f2E72T7
`protect END_PROTECTED
