`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IF0pOIoCvlnKybWr9r+Zkxs1KfmHIK92nsztC1hm/jw4de4hxgTZfVy1oZoRYkG9
7GnQSElHFIGZMj7Dy745qEcOQrfPqFhqAgnkLOYgyLolFeBuIGmaFgkdIfRARKez
YfWuLWT/sqYh5qPPij3M0rZ53mJ3nXL3pxXnhsHYPMVe3cU1LQjBSCbUhGgy64Xv
0xbF/MTdOfSUBGMoTT+FF20W2k+oyJPRrFmqwAc73T5gROV2ul+PYMYhce5NE7pE
FubUn3QBfkFazVc9tYyLCmi0LJ+BweMDfMYtBQYRpWDdA5kBHbygzvYCtSupEWzC
PK2ZCiXDVMi/Z6alLVuz/HC1tv+WZAnU+E6aLa2UV2+NGJmCDsCZURf+c58uUgSW
cvyIR6CA3y8RDEzfaKrklQ==
`protect END_PROTECTED
