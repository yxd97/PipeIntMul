`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CxyCqEiW+pJlVoUz2Bj/Edr/AxBSEkOr9Qa7TvLVw4ajN5/G9oBMchTRl0pT6VOo
sq3UzGDZSkP135TINPciTaEcmZI4vtOIBvqyqbOqk+guGy9XgD8KUMrx+ziErdkj
frEpTq0k5SrWWEVoi9TYwgIzHmdBeztVPT22wGLnL564hj9nzuO2aG57lm5bkbD8
DYZqk74BE5rbO5oblltMzV/+TyR0MYo+3uUGObYH6+q46jnebrHfxaDtR0lMseN2
/zUxTfsvRueOa7Sfe4QoYy9kidGjauXXuT1G8JzkZWdbMZFl3pPjzcstcQH2Newv
eywPX7gH3toOwPAFEKs3AKAwliRUmIK/ep1hHIXr4k/tLZk6n9eIuRI5f/X3VUn2
YqIee8vdBggyXAf9mqWRqSDXfs82K46RFeXhzBJ6UrBZLczmT5azxlcvEi/oX/b8
bfti3BJQ/kTpc7ixYf5gg6bPetK9roXtOI91VFVZxv8m8fdBMkRcIQEj83Cpktdx
Yyjq2RwuJb8/oxTpHs8m0ROIFA4U5BcwQMMor3r1ZrFYOz4Fd8ooKRfqQ0u52pAY
gbPnGKgt2RJ0XYNQWjd3AIJzdGuArQCX+l/iQoys4xzaQQA/enLgMN/UFWzl6F7N
NWjcx86M8OPRWSx2mmv3aFfIfInp4rNbFMV7N75p/w2+MZ4vbtvxcp7Og36wCsgi
8Gdm83Dr/lZl8dR2mGLWvvPrb+1APCEnqjSUIFlU+uVaOUQ7e/o0i1GwwqdlzOem
Rxu5dJWLbcEXlF/Tsa1n5Sf/CGVdfWxCu+Xo2zYqT6H0+A6cuDO9pbGq3OVXLBhu
`protect END_PROTECTED
