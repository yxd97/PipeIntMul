`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PAX8OHYz6p3QRA3quqPXY9RqI7nt+Y1GethLFQk8YX0d/IPzIvpSgPgIsm/0A8r4
+OPVUkg1NQJWXQSm+KqwHXstJL7osyXfpfX3Z9txA4lZUD1j4J7XsHaHpvfIUkHX
KN1EqPadePJKDFVOs3vwdedacAzG953Nh6dEPHpHCaNuYVkg2FkrPCXWOom4cI6u
rdvcZ0GD5kwnrApOte0t3p5HkQpjU27fQ7abw/Vz5EVOjbXnk4LwGClX8lo7b46p
WbAXGpiZymQgph3/RRfK4waBJU7P8XoBxibEwb1sAcBl749NankLCZjAQm/5FBCL
Ez7Me/JBgV/YCDMZOuksC0mEjKzsGQXNUGee1dl+CCUM6ssrzXbkBBu6JKGKURZK
2NgkF0gRRRgJ0L7SKOYYgSdwsx4Or89EC48sSPTuUpGd1Ln82RqLIapsy1x7a8v1
iJB2zhmm09kpUl7y8PY4C56zH7mbrcYyfVkdlh4QzKKLcN2fyp7GparLnLtRKjXq
7krd/pVofhvOns13X3aDkg==
`protect END_PROTECTED
