`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VG9yPgsMdC7pytCT2Yr3AhM1yqeyZhfqDKsKWxlJcmBTKbB6EsdbLejzRiM1Mim8
+5Ep37/AUMW8oWyfNviPGeVzJARad06Cr+YpYsUr2+SAPLrrPR5PMD+FxiE9Zs7Z
XMsmQglvfC+Qch0RjwHwMMiRUYsx8OR66UMwYzlUlhfSmDxam/c7AXv5khMIC+Q5
rTf+UqbbErQMhabCqE5FhMScDtbgXDKCjy1BCuluM3M7dmG04k8O6ILGNUMuGwFr
ehUYSJ8rZ2KfGbT+MoBvZ9qrLR/ea8O+RLD1e1fj3SugCHpmVKadGN0boibKvAip
QlDdjnHU4UnqOeC56p6nVNhhbNib7KOJDriTVGel9+MXy/FkOK5q7mROs4GquSdl
50pFvERkbvCCKHaRS++5aISNkCUccLv2opQrF7LaDBnR+WIzvPkui1bktGtIGVT2
H+ph2VOF3AwDusJspld/Lf3aNwgirlZVBg0rn0g8oCSR1EOFQ2DIotH4HP8QAagN
tDAPAXalNZzczh5N8zJ/3jHT2x1JZfsmsKkufd6kbtFU0oCCNmOjobV7eDVcoM5W
r1PbHfXR09j6dccYSNlaFKTnPHVZC1PqndHRixbRaB5GD3Kl6A5KLMoC7fW4FYoJ
DyhALBodNWNLJO0ADwgwVHhR3rH2r8gQODED/Xrdv5CXBAjIXxAvWQD1rWBdOas+
6zro10XnomKWZwgnhkQwrDs6o8DZAXVxZ5nmjJ8MB1PyxXh6eZul9AGEk42jlnNs
6CEXN/BouQyKb9yg/UNjJntiMAayNdZYnvMaEsIJVpJxCa6l5v0zIYClyXmPiwXv
H0nVTLeXwQ/lV5V9sYuvbJexvmaq42Of3a75xl9SVhDmVAGqi6WfLWjpNbrjlnCf
96pdJZH7n5MPVIM5n/RFoEHpWGzXnjEXWGq57E4MKEKixTIHQe52JLoEEXXf2lRO
SxD3Q8wFx7ZbF7UmiD2HzEGjBdgJ/bf5WOITyhkrE8+Qzcpiwx0TBKlox5Ts80a1
UNwbxsSwIoyBeEmAvz6PIr1hKZOK2UEDZFq8Ei/xZzDA71n/1WxfDqNa2brcIsTj
B+Px40utISbW5Jnh0zQh9dLVOiyxrIRmrCnvpdqzPoCMfrTOqqpngp87Vl2fam27
mw8xX3KT8wk3jnp2ipvNA6xDvVtxB2097EkXkKHS8L8=
`protect END_PROTECTED
