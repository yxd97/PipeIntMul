`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ZAFkIMTkl6pyUzdoXis0NIzoaTSiwlr3SP14cF+rRrKom7FqjH2K5FUginVcrK/
zmMkpFEtQR0eBYP2R0TKFzOnEF3+TfDXSxz452oSW5Tifa9EuBMMc5H+c2l7m6Kg
oj+szogXNKXKzSxl7JFmRRQeBhCR1dtBzZ3hoa0/8hDqRDdEELgQzvoBiyLqVVT6
pF2tAfSU72k6nPJSyvQqLLE7aDHTVTHyujDxtIx+4ZMirmhX+7MB9IXoi8GkAYdy
ygGJS00IlsMXSZQ40CSSV/A34BNcbRWzit1v/WSilFRtesFTC5tJ/ZhdEVC5/XkL
dCU7gqw6zRp4wzHXFeA5ovDQ1au4herK9UIRqVJ2rK081vJ+z4UgP2fHvVmrWJIK
ozP5VXxKdbI+r/WSzaoop7W6xko7VV13QYg1Hd3aiepVR3JYORXYF6T7pIGeho9e
I02VfeGja/YdLs9n4G59NGa09fI44L80YNhCIVb+C++J5llcGUHrdbewEsCeEWq1
cisc2gELs9v+YEjAEAgNcIqjM4mLEa8ZcSdgYn2c4q8+WBitsUHVNtJuUZ4EfKuS
CfbcfeNSfudvehpx5kvH44pznqpLTbDRI94Uprfa/LuNXe7NNLoxfRPaajnlWYjf
g4JnFcB3RzWRscREVXCQ20vcXs8IJdeYSfudaJdymgFQn9lfWTsxWcWAenDJnIbS
`protect END_PROTECTED
