`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MRZnSj8xTXKNN3jwIvRjBJm5RiQFm6yAJVttNpd6nHYzjLdl2ZalkAM0wq8dRXuD
MYyXNF0JWPDiJi+v/XR6DNtlSUvZx/ieEcQ9LotpZ0y96fxWlbF7khxIw4PWSm8Y
lPoLgnY8qCsZE1L3pjXxPkOfPqqdA1Vp3H+Mk9LyDKB/OF4/JfiRdZENyANYmHS1
eFHIm6RCKADUFr/vU9H8LvrxLgA7pUPCpla3AE9IN37+gkm0mmht4t7JBO+5a7yr
VlboQtYfQAM4lNq3t5yVh9uFI8kiqw3pxlO7t6qZE/1MCdpdpfSq30W308H8/f4i
wkD+goHb3vqZsowd0KVpkNnF0X5qcUOd8Vd8g0cBkQeEFkelIEBw4KTO1uc3MfUi
Iwfc1FhEbCc9vHcYAUhsCA==
`protect END_PROTECTED
