`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dsJ3910Y73Qd+4qXu/v5czwXMMJOS6pNEwzUSzQs+w1Hm+OKl6butrybVkhVrYWa
rDDwCzvlco9un1/v7BjwFbk7duSNumTChN+Be8zsRnYiYg45YbXsA/Fpyrpkn2Jb
c2WKN0qp8MGphN6bBqTDRCDj3khlgF0TXTiMaEcaWuV19CpUt54gZbi0Zee/b/BL
YMe3yT6d5hCUhmPm5SxPCKUc3x9Ji4KV/ZSYwCbsEL+uoXO8vIlIfg+hSD5S3loB
V7z8XJgA4QIVeKV7ydQ/Nkpkp3R9aH+vWs8PtoTgInGSG2JTII5FLMrJnPao+usu
OO7B/RK6HoIHwEIZ3TIn+hVlaxSUN46rG6aCUAAU3W88epR5f7fl37CnzeMJMQhS
gnt7FMsdSzOjw0nE/mYHTS7yYejFizYMsX6gAGFcwkGxFTjMdrRsp2T4JOezpaSN
HINQSrh3UXax1GCZWCLycI9oHfMHCgJD1djuMr0GOPihULHZLhZo0nNUrtQnmo/4
guMxny+apXRv+5+uQOeV36ZiRFQwbi/ls6jnm1tLjgVmCu8FpXRlTW/nn/qF7rKo
JMiceF80jSnTARp43a2hCKdFiZhbovBLWh6vKEKKgIefCdf3m/4xGCxtn9UsM9GQ
tdUaGkkg7K9kPvDK0k5BR3lcqoAmqlqUyb/U0UxmP6h2r02ro3ioHk7C0E3GS20W
AjRyJSem5+aO6ZR3Qb7YdL9w5kI64epeT1g1nqlZKrXr+Hvqu5ZjReB/Ty4HyIKG
IN4rKM5JFaMlPxCBwGKNp3un8l4ipoRXqjFSL4QqjUmH+gRzqc4rnZ9jA7mPI3ep
qlG5Npa9UG1j7cUV15KsCdms3iZkDz+3hI6XPcLBCPL4Kz6x5h7j8y2cMZb3lou5
40xtXuN7z4m0lY0kFp30ZKnI4AQAfmYA42XTo73/RdruAOQH1/q8v7Abzs+M1TR6
nXUm3Lr6GTtWayKQ0ACO/RkYdD5xOzL0K0OLqUgeYr+2AoOYX5wvOzj221atuj2x
wXAZNi0CWLWnApjQddF1sLkhLLuJMMM9f19t2X4C+DcYZ2YaER404GC69pBoyR9K
/EyrdcjGkbbQW4Tw8j01CRW5pEa/ngKiRnow6+7dpa0tRxC/G6lT7CyDSRd8K3NM
sLpGRFY95NWZXd5c+zSoBOB6UrDIOtj3ao2ZVoR/tVX2W/N+zGM5Eo2z8Sh7x1e9
81qFBzuHgGEXcSWpdFrTNrGp2EwcfAZ5e6KDKDjUg0u5+eUKlQhMYUqqaeeHykMX
Mxuu5EjrRqo81EshRfGv9jXQ/l6ky+pJwFvt38L79Wirt3CUFyjfTvwoaCshLWIX
aFGodXr8e5eYrizG+2414PB7RL6thh6Xfi5UFYeNf7aa0RgrrzZ0C6So1s7dT91J
UpQlaEoBdcXAWp8MFYVB+VOSCp+fcj3NozmPCgm52ZmEuhWlclnE2vU4/+BZ4Toq
N2dlvvTm18wTppvZScIZYtzycHChTles6a9iPU516PZOBPGh3EbhtMI3ApmMAAN9
zs3lwzCnVJ+GFtUt4c+hofElhcr+gKgbultZWyRi29IEK6iWWpBEtOQSMHV5Ip6Q
DD5a//PNNJaIXn7UDe+byNJcasdat4zw1dsb1qLHFEXNOR1GjSeEs+kFNKzLEPi4
kwTnziouz/PJLDvRBKIvhsSb3R7yiXVKdXo3x0rmKAoYDoNwLe98PjANXeXo5+Dd
6AojZQ0D1wuAzi2BQgB9SIYhiLyYsNW/f7yFuN0Hzj3pKBJwDegy8/EAijA9yTkr
JpCxJ25cTIMBPfq8aqeXVafNTJA0ooRhgSL3afrkuvPy5Cy1IbsYLVD/unGUnXhp
qPW7R51ChBzWEOq63ctNdO8siTWiwcuyanWIBv7lKrOgOsY/PKfSs+QQQqpgt3OM
tSqyW3FyqaZcfhet6gf5tFlC3el+m1rUGuDRvc64h1jWFnx5ghyybEOjRpX27oxY
SAvDIkGBd2Svo4AUXTSrJObf458wVzaKqcMDVYdtE3CFiWaEdSb8ZLCK4oygsWAI
SfEULRkgZNgdIuhq+NRUt+QGI0NgjBSbEvES/2AxlOPY4csrIL5/ywrVdnQZuYlC
etXiCUd913BnMhgyRMT+5WNvmfi2zl2nSA+M5CQXGtp+02UKkmfRqujQdYCc+b/9
me2B74wiDRBPQYnY+iWi2+RPPm3QXUwokvQrWMx5Rlx7QHcY/+aLz79xHTWTxNOU
HA7BysXaMfsED/WZ9ILDjLh2bO9NTvoe1ItzQR2FQsenoX3uE/eiBc6A+xwy+bE7
dZjl92G29g/C9sgRPsIhwEnDuLdV9DhRArbgrnFNrUxBJVAlkMUv4dZs0QRkoBLE
/jz7PFSgT+KwWuB5iA49qRw//bXB1/bxLkGPRvUrYjKJQoRRwPvVyJp0ejCTiv1k
osisN5oQIwazlrvEgGQeXtemPDnPRDe1/J7cuHZybv2+PRdh1sPbcgeaUoPJOBM6
SFUizdzSCxuuV84fMDhBgv5yxKaRWwCs+PXC3+8GMIXK2ARyxpDT5LShArcmbbG+
XxWbaC9/gNEiaQQh5i/c5kmDm6+lplNC/u8BX2rA06h3kmaJymhKfjOi9vC3GqgL
1KXGiDnAAFhuKqr2L232149V9bT8KCvAbrsZ/46qVRDZQ6b8J65QFvIj9RZclnsE
3PEpzcFfGLswaFYJ0FOvYPFc9HMNSwR2IqiRCSDTw5PLGhkqX0wFVmABz14qw1Mu
9a5fwcsivMDeuLxUZIx/liy/n6VYZh0+VqG0X0kcTIRYFxF72tIoZ5NrUcPBw2VN
IDH0wBMPZDFTtP0EO+UfFYsQ/10vPrBmIIfGCF7BpwsfuwKG86zPUl46DVuw+75C
8kX+rNg0epN6RQWuDLTpy77fnHs7YXRtR9iLz1j2seoI9Un7ItTHwa2Gu7yaOq2v
wnU5cavwIrSTgSJP4uoiSdGsrm3bY1FINCLcCxSJE+RqVpxcGemDBmLbSYzy2PkH
7DEPdytoiNzIcxXbPNb7SfQKoR+3HSGA6nt5y3I1EFV14ovFANxPO5Fm/n383VXF
rRRGQGJ8y7GR5j3q0MuE+v3A3Dws0T6iIQ1/xb7p4lBGqb0w0UPxMIb83HgMnpXX
O1MHpfg1/oTfwDVHa/2n910pTZ3fy6ZxCh7Rp+4ZYJNVMhJg3ETlBapeG28UPh4y
ngJOUj3HGmiz9s9WIH+IhjhFzaEh7egj1o5QQDd4665chygBuaaWhxMrKVKZOXJc
SJKk/NepFiB6gs8OgczP1+lPdV5On4Q4tu1oKyg/JZ50LK+9MwmdwZksws0nVpjW
FiU5R9AQAkWr8nZ11jVeChxrdeYzH8q5mIJMEoIFl5SBmwP8T13gk1hH5RIZAosP
TgoymkUFsLDqfwKEez5x8biyZ8uhJlQXxO8NYMkb8oyNBOxBIYHBsBu6GmdYcS3Z
6EC5t7/ASmA4go+sPIh/cI39epzIkI656lYczVYCMi587mfhewJYx4dmfzsVcWaj
zg9c3AdflRrGJnhAAB2HlctZrmxUWANhJgpu2pei9XlQO4a6+b+TgEc4THUSR/fq
AJe9vrXVsf+VKyt3xySZZbMycgc9nh0f+qH6Q7679L8YsZkofwziig9UaP+JHT25
rTAsiH9ANYwATl4lc/sBCzFMV4DwO90mFD7OInyZ0Vqv18cagH+HrTObFhjdr/Nz
r6Px80lqHyAOFZwq3HjM0dHfOGXUiA6mgrCUuEW4z1JWyTM2zDc1d9cWnigpUdz4
8nMb54PTRybId4MfQt5pqL1XaOztf+f1yxckLna+SwrIQMESphPY/eIadBczVh4t
56+IE9WAXiKzFWu/V973agJYtjyPg+20bFrQ/HQ1RlIWtAOk4R2IVCBM+xLdkx3N
DhqDeUqlCZqBQ4e5EbiwBpCLP9COt4HO/3sS+ahqwwSozrVjjYyJVaR8BHpGTfT9
ltp9k//s6f3eYqv0CAS5TNgy4K8Xyvi1AHS/Edct1aaxUdPLpvjkSsSa2SDoe7Sb
uCss3HT9hYRsT7rnp7H+oc+wMJ1WaQSXz/v/Z3zdcbMNpRLOaqJTUEvyjJ/Rz5uM
wiqcH7aQ3JAtdT1CoBOuLM22Cu3bRHfrL43ndMPVWoQHka+ZKj11iwrH0oICKA7k
LBqa58nmGz0QJDZ7i4PpMdEv5h5OF8Izz4WdVJSR2TR5gb/OYDEFjLHx1gtzsXjf
5cJf6J8uBjKrwg88bT8tskrxl4PlfQe5v/BmxMJV+tnFiLXYxDzvwxZjJ3X6JQaU
itR37kBVKEI8aHJCMLj7iJVQ/7TOMJrplA/J+7ZcDt14ZQt0hIrQKjLj8IYu1cWQ
6MSBcdey+vDLZuYf/UqttvdxOytWOLUFRL2PZOt/AIwWPfNIjLrmpncrlybMRb9q
RffXRB7+bdOcnsRLR2g5zwvOk0e8l+jgNnK2v8/SRDEvkBIvb7DUaZqPxNnSjVtn
RE3u7j5PlGI5VqBaWisBOv3FAWmgy/Ll5k7y1Qq9uuUdeWlF3UZwnshWLoGTuEAJ
93UgJjnuSQ9XfTGgKLrjBWghr22Qp+yU8JjaHl2xW0lUBH5Yq9SZ4fs8accjOsL4
/MWac/rSqfpKMq9P3BDnKAr6YcvHCAq+9Rf6BIuWmSYQ8poc6DULtvpWBpg7t/he
CuVJ2Jaf26GZxd/+9+T6ckp3n5P9meD321luuMrSoKLVbe2B277E0OrA3UCj1TG9
Da8cT5HJgGrs08CdaoK0zs6soSrhrOlsg3z2OMIjSBGNudZtEdzSO9quKOo4aNPs
xvG9sQCvJxUpEIvmDMMxYFNyMZWpKsqHyaZ6JahXa5zSWYwJToJXzPR9NMZfheML
3BJOM0w6gAn7gj3hRF0O2Id6p0Udxq8U9/jnw8DD9+JoGSlO5ZLkaQ1c5b9UrBqM
i8vHOiKgdZ7XsglPhDK9260tsu3HUlsIAhyUMHuEKMb7cQUZk3FWyya1oJdreC6P
5eI4vpBAhD8WqiJabNWMoj9h7SerFehc6BV+YOa2Rk30P795lLpEzbNY9ciqTCnu
pzH/Du1Nxn2CwCnxXis9gN4B8S0uGO11aXj7CfUcuBwSTuLaLzpB/B26GWWHXL5j
2+o0Idg+j0CSRJGf6JEpo63vw5Oq8kHOwcjMDeipdVZipwZg8R42rbIYw3DJFR+F
qFVknE3Mg2/IxGg3jbMaJjdxHebsF0HxcZX48yrAnGCvz5odU79FILpcU3AVXzDd
ilRKEEvWQKV82wZFj07F491wqUOUrJAV4dmMp4gcVzZ55zexUzpAPisd0hBOWLC7
PtjDL14XShrXqurqny6OU3GIfTDq7VB4/rX1ziFzRHYmaKtbWCTHhxN2kG191rTw
J7Jbzwk9V4LeIEHvtSle4YjupiNYpVwupKOB0Fl/N7z22C/uB8dEeJKc6Qi7d7gr
Aapz9RzuQgZkvMYkU90JpabVXqAMetM/qoZzHdUaJXaCCwZusaPHfD6dUdiWxxbB
kxady5SZ9+AkIqGPtZC92hLhBn078YWgo3GhFWnvvpBggEQ27AXk3xWma63rn3Xx
lQInQ3NWwribfO3bnPA5FGyissKvWNAVajvVdBhmPUdInuDyOCJKrvCECSmUOQr5
mokuX9yH5rwrwW86j5yFSs60yBB2XxxtDxRMqAarNHPHlDEOSL+godd4MbeoivQO
`protect END_PROTECTED
