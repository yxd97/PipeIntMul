`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AZhQEbF/3w1eq/aTryov6YUmjOinxe1GZ/znG1WZSorciEwxOqphPT3y7sQe5opg
GBZjFpxse2XiJHKrSXHKn1GE3tCGIf1NIGK4d4kYeynUFR5zWLAY/CdrlyciiTeH
mrhvqq9BeIMy9fdfVxGAOmPHoD+gxu012Xb39ZUH/DdXcP6Wh/heV/XO6DRjdcHU
dDNShAAK5pNPgKqvES2R3xDw00+HuL/43LnOpfd/Pzin/j79gQsxdpPz3fjMG/eO
TYVuIQ90SbJGbhc+m+TLarQFwi9OvA7u0eez7v2rLiRxGkXNz2BIQb0XSF4tuDDO
SmjD5ZaNTc/G292g53SI7Az4lydDTcl+fpSRT55hAYp1H4aezA8IQ7Zg6OACYu1q
sHSyYULdcDJHB3Mvt5mzuSfo8s7sv/X5UCwU713kGvjT8ULEvlPpDrUa6Z8QdVez
cUHlDaeZP5ZxtFLG/B4nvGa44Jg190fndxojS1I1IxkfuAn37XZNkis8gtkCQHQ5
PCMzGDBDAJPSiA0Mux4yAYP5fxPzH9iXU1TL3guob911I+1/KneYGg7go5hHlwFg
TZUXm4I9Xc2qF8i3HPllF0LggLj6Ru+HKrX2ooC3J35NUtxON1IZADZCnE7KDUbG
05lBr3FIimIoxoK1j9glSKf7GFU4L/7Qxv7KzryPnfSVLq7uCFEug1AtMo9khwTf
6W4isXCJro1NbwIzR/U05M2hQyDhUIe5ZzEsu86UzMbK37DH6ShX1M+u/5DzQvF6
temGqm0y4smyp18yAJ5I7C/xyJFHHWBuVCjwUBkYZBconIurl2mUUGbndYrMTLpW
NsO/suOtCpCnUeONC30BXbxkKHBMvbBd6wgO8CggVNT8L0TEZzf/urZvpn+Xgp46
AaFZHj/8K3DJtl8fGGsnmHQX+8Jpuu1zB1bic3XbXhQkQKLyWSWZ1ah+PxoCQIme
`protect END_PROTECTED
