`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5ntAFRwvN8ly1sPejv85Fe7ddj3m13m0h63mhcT7OW87fkdVta49XgYBYsIYiyI
nasOkUgMlOLSvijZIQwMMRFsSZrvTyAMaIWyM7TGLeRdg2R6GRS37Yd3o+7N1ILP
/oQL8UxODVuGuE0slIj86dw4yx0UiLEJypZtQMZs0Yuj+TWoew46abtko0jGZsEU
39TnVx5lAxvTc9Q7T356rBIMefGBXWes9+XeLZhT1UsnMjs5M8d+RvzAGd1w3hTJ
DxfrWrZ5yIVATNSyvJHhDP34tCuako4XGvjXzOVjp5FnNa17hd8eLov6HLFwy72P
sk5xilGIf+xyoZNJtcKx2sevRJQ2wuIXw99+X5pwV6aMVWOGi9bpwHvOHqSVLz90
jbcQCJ/FZI7d2TcF7zoRy5rrrUTJdxt81wl8kU5Fp9ib8OPaBz46ubVQr2JkrALS
eSZpIHE78oGL3I34go727Ueog2xBa0iL+XiADOI/xjfxU6QI+mZ/i+hj7gqmfHfW
t/bFapjhDb9LwefTe9P6tgFfDlzlOojrmxgkUZFM/qwESmWbYfII4jkEIOtd5iNI
ZM9XynFcg6UP/LrhBgW3KdUXQ1IELkA/TXof5ZWXvNoHlcd0PV/9IEUkNzd7OCq+
VGPXVjUDY656oHIZdTbZZ+K23afmRdEGqIG4abd1tAKcoUTcI/CSSLwWRepmuCYn
uO5rH0Wl3hkszQou8qGY/LQ6w49iBLjMw+mhWiuVyncHBxwKD3W1r9Fh8vsBCRcr
OQwkjBGMSF21BFEJbwkQd8zt4wbnqrm8mE+nBQuV6sx9H0poA/cljAwUK/Dee2CH
KDLiyAjsR0rhlcBkr/yxV15URoBuV8plxcXEvzC/kJfxqupF3KTasxDLG1pcqX2t
PNosM7Hjh7qqw4goiDlQK1oqY85/1HPHBeYGP38Vg2GAOxawjCEqXVD8Br7pEiwE
FXxPrRP+LND8/Sb83/jmQTvN4PC4VnUP+xXoWH05aBtKsUw6rd9fV6rRFKZ7cnQa
`protect END_PROTECTED
