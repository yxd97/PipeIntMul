`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiWQ8LpQ/rv1hgMBACGka/Zde8HI48ibWuJXHYarBcisYp3oIdt7VRVybf/Iuhsf
0udthVhP60IVn4G3rVuVu8AITH91F/gKwSDV/G63JcC4utkwCFG/rr1yv0qlChaM
WvAr8PwP4fJX9Jc+3G+LQromVizeyBtujlErDWY7JxnTdW1adXPXBB8AUrcXpeaG
69vAQXloYLmQOmPf5bnR+tfHBy13ZxnY77/U68jBcav3fnx2dR3o18atzAuTfuDd
MB3jZuku5+OOu540K3pcFhP1sq2tcJm9yZIGR7MwJcUSE8Bay8p0GM2niRyqnv1z
Bpa0r5/6k5dLsDLmghrduRMHOrHT25UM4GIuBmU7ngOeiBZOQ6gahXfzKkhIh+Wg
8A5g1gavh15NmKKdyFYzqPpxWkmlkQHfDqfdA4Z2tkVbt1xbUYhsHoxejGa2nkJA
9C3U4EiU6CF0AAt1m0OZ8GCqW3BfhG2fKy0stuEGn6rvbn/kwR21JWIIl0VCRgzC
NdARsx7TPa3b12fJoOZm9DMGODmUHbt4Lty/HC0ioSASetymiXKrfNhfVidIVoae
gX+1QgJOVhE5ZMUUaNpOaBhK6UQqoftSTUMJAWltIXLoNrZ0l7+ZRmYr4/akeiMw
647pwBdSOvI2zT0plkHAkAKN/UiGtglaUMdhTkTcFPd/ZW9edpsqiT0K/8hhbOmz
NSHt3d2sePml2Xt5Y1yY4kMT+6qWN0i9HbigiBaifZu+98K8W/2ZopGk2y2gwib3
mYGIHrO0eYhgOiu6J1LMYCIXsassSDHmC3AJullR/RLwS/2drKvmB0tTNYYtoj4V
DT8eqLPPknV84hbJclmTBhy+o9cgMI5QIPELl2hSpjKU0TCVIeoytFc0K/je1kva
ubfMU7PuIFbDgyYvONegdVuojT9avqOp17VUE4AcpqnYKtIKCD5ns126skPXFzdp
jR9cJOVSr+gsm45keUFskV93AKJ1Anke/G9Sw6Fl0g0unW/UG26AOUAeRKHz4vnJ
hoLlqQh/3QpDfpG/SPX5euV4Grsnt+/7jlU4D+0L73mR10vTP6pFAZSYzCQWs2bs
WlW85gt3aWIAE5moyqNsuLLQxqvHfHfafpn3jJZIwvpxARQweWW+GjTrzXl3ov0x
KiOqPMn2+921g8O5odE6NO2B0ovIPKtJaih6S/ZsYtGi2K0NBoflcEiak9k8Xdr3
zzHhCZzROHj83jtk1KQM4wcOqnIKNyh9PCO7uucNJ+3MjJIve04NPcqEq27cynpJ
bmQgJOSxV/XcFy4Z4zAEsV+tRVnGIl1IUvDsTdWrB6McQgZW7LwqtiBS8Mskpuzu
rWRgphuMcNd5pk1rgSj4p40Dc2LOpsnv0FNHYSoL9ZfzSSqjfLaJ0V0limeVnn2n
torD+CckpKcNUGJXZC7PfqScRyixoLdlHUav3QsHusEPFExrPOzyaee6I9Yce81J
5TcCFAyBJGRfM3jWC6lmiqiNFRpgS4jguYlyWvfHlY+Jpr53/y/Jm97WHo+28Q87
ZQ8Cwz+ufzg1Er1I72NUTGNAVGpvwQYRq/Jdu7ppZ6EOHFsCOyPLPkKJo0ZRnmlT
aXaHCCxJP/swRl4JXj5r+p/KGJbg7VE3bDLok3/oedZcNc21jWFi8Xu653TLdWoo
pH3vIH1Z3Ae+nonYJUcItLRPLYgrAjeq35bHR2dlRLddkyBN7sv/D6J1AVcJi5/t
8yOrjItxfvnMZ6lTAyw8YOuYeLZVyYsDfVslwFauTJohvied2Dumj93tpSMwEjby
UW39uQY6fEU9kp+jHyptQruIlyppms5ma4qRq+hJw4VpkXzKCljfKv6YiG5Z5VO4
Bd8cOnppKmm6Ynix7IOPuiRK626wdpmWGyI0lsDUnOohIf1HCW8Ih/xhDsbh+9aD
ESM/sUJqhdMwgHsqQktjgA2rDBouB2ah6xQxKYuwwiKcCgunQfM2xH8KexLX8LhD
/rJfYP/Y3VZOje/2dWNKjEpEpSK90ZtpTHn6NDzaUSP4Cv272MIl6gndhcr2K6D8
kcg3O5XgqffiZwSx3ZeIVB+SbxwnOSSI7Z3bHxreLkUoTutKav60j9FAUD6GF/Cp
i1reWwzE8y9rY6/0CxYAGxC6GPVQsh1GiArc9USlzjoWv08l8GahDBmqJ2cctsuP
7TA36CjXwha5to83CxyL9bL6zOrwtGpq1wvgDKVN6dN6OE2L69xbhm5MxKXPLjgC
0EoAf2H7+mTeSAZGDZKo4O71WLlYWe6tRF2jkMKZJT9PmqZ0tATT16aMfmoHE2aK
opY8t9DMWY9CHkmNhPD8Qw==
`protect END_PROTECTED
