`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DkQfkxcZYx5yNq5aKoLAhQZKzHKKO9cn5GxKucg4jSQw9ivT0MwR0eYu2JyuNLy
WsDpRdKdy07Cbyv7zMeXhNQxc4N0rCKeQaKTe9lfCkjoxMRM7uRJwsO+ExvUzZs/
fPlkMM4eeEpgWp0hZLuQmf2dZfkSsyGRKi/51rH3Zp4n4bM54tCGz55ooCvJQuKv
BWTDPz7hAG9a1g4cYezA/SiT2XmgPlIY8N7wZ1Zislyn9mCd4fifTi6PY2ELUr5D
SpHdwS9za54B9jEo/2cg9jpzUqCKavUhPhYTOa7/+4ckUdvlAG7B5azCrJCe7eZY
FrOdlFGPVlJ3lzUZV30UKqmblJltqbTWg7aPvwd7V+hhLvy+h1JJ97ro6JIDhsFq
TzgbuuHy+tOK3j1kWe2esSrPMIu+P+0xwQIJh2ucuGgFAcv6zL0K6e5JruJx8xiP
RNUOn/D63Fh0wI7BXCAvZ89UtKUQ6qWmMkeSZ++zy0Br9WnjFUVGjoKQ5sUIrezU
dh0TsDQ3Bk1kovJO6L+vxK3KI9K0VL4yrHCgacxqObXYYgV13WKd6p+b3yVU/vc2
`protect END_PROTECTED
