`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WE63JJoXZCwa8xuy0JKY9TfTT3XJKlXLYZVIJ8sxwaIIsVuzWkyBFyzA8LFUMEry
t6oxJ6wLsnGx36yDor3TGkfxZUAv52DPjWK40LnYHNmatkRNdyRhXybFi89h8aJN
ckj65FmBFZDm+VUL1xB09N0uTwC9sTx5GYhqrALHpAA3kFWPxfQtsszNuGTfMXgD
adcLi+QP6/8ryZZunwJjxla2ANl2OfSQ+/PU9S1nF9AA+lrc/rtCeRaZrruAkTY0
4cc3cKjUt8cRJEA8YtA9VG9DCYc5nNM1aIuUMMPdaT/Kvmw/ZHQf9s+HbwS2MtN0
8JPFRSD/Wrv5f9rVc3wqrPByjHbr6gjOGjbCZAtEZPZfR2UGRYReFSqKos8cEdbD
RRkkKVA9/Unx6NPtQ66ZEoxKfSjhi+u7RwQ2nx1oboA7eFNRykBGPotTcd+jlfwY
Sd1MFFfFAakL0c+fCMXEzRg2WYDqKLfz7CQTDBvAFk+X3cv8I3fGqbRlEd1TC77t
m+KY77gQSOC3F6n2BhY74i2jIIZxKh94xYuYHDJsZwEgWuhR+rbUBiyyZzTZvrBn
w/6iMshTB0iudlSPBuYDriTqJegKFSIzqEtBNSXDHmA5WCBRetgdrJkdDeQHxZ3M
yE3F/rGTDBqW5oQfaXC6IjuFA3GfAyWhXZ8SI1sKofdHOkgYqISaBRe535XP7MuJ
gd49lxggj+hqwmG01ris84JCFz2UKZTEjoffM25veLdwsE7VcdPcIssKG4QFOC6K
Ce9rrta2mubab2aHxlLurlyuM2qmC6NlBzVa40Ue/YJaIIR7FB9q47IpUmjimDLs
sBjBAatMPgNxIj/MTH76xhyeixIa2z+b/C/No6AwMzcFoG4QK1zja1TeGTb0CXQK
Mkb5ODJS+YtGEviLCjUJFuIOqgsHzQThfnXk+Yq4O/NuAX6dD8e6TQkt7t5oIS4T
0crfHQ9HQComFyLLfLYgIuFXxTxkEPuQQbNpDuHobYbjsU+gWz7fMQMU63fds37g
Hk7GJBbZpFuMFN/wbDaT3mRb7ft1g5b220TXpaQUHgAEscesVmzwbgCQlcCXZFex
dGL+FTGlMm91N1uAHcGYoOp+ZNPKM8Pe/NHNA+uZt029gdZDtMQVVRZEFFl0zd/G
auwJI1MD+s8JzjZxn0Z16Q==
`protect END_PROTECTED
