`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6WtRzxL0M8AAWDLhVTvN9BvSC5kvh2cKnj78sR7QGbG8yuk1PWe+IgSHBAWtKXWy
WrYprC81nyq1+9/vK/htBhCW6N9mwWWmvq6/DjYykS8z9j2h+IcJa8XUnbRTzHoP
h9HaFHgxbLATcdLnO2oEwwmfznK1uA58yA6rmqlq08wVVVfgmmXNPaUmMywNECIb
dIzHHO0zkm/rs9fA7ccwQ7D7JGiJFkX1xDZJmK/fPMAF5mrCshys/dzoIn3WOXWx
lKGfGlvFi0ov6MAEoKDDwfFbPlo5QRDVg6Dxze/KhS+JtOnqVCX0nvQFzXE5kWJ4
un6SFyb44ctrJecQV1zn0QoXEjvUqHkeyVrtqkhWaFVHfSegQRjo1ykT6wMBlxDS
YGurDdIHL3CwaQU/PjYcHsF0jwpweIiUgHC1i5IUdE16/m0dPpYLQO+oE/tyjm/F
jWj3+GELmfeLRpuFz0KDRtYx5cjdP5uZ4ahlD+T6iDAtl5Pn8Zlq9m9m9X6SQ6D/
i48xF0y770xRM2+SYMjgnVc6yoxatT7X0z0oyWeIYDuEDFb60tHOSJrlLuhM4oaT
ig0CBmC3yyVZy0ckVANErefZD9a9B4VCmpI2QGXD2XP8EOl4IriusayWHJ5lAcp5
7+X28PWB5bd00n4TL1gwpBu1/idH7gjw4t8OxgogeVk=
`protect END_PROTECTED
