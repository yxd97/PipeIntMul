`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nPxl7mwNKjPgeGd5xMiWZ6DPFzp/UvunWS8kLcpYc0OdL2sv6D+c1UObMV9HNJeN
ikbHHhuee81cR22FUwRCtiKo1OdcQ5PY2WR0EJwZ3tkvmBviMizxzLais9966hZS
9/JEP/YenjAn1l5xxFF6fQ8Y1vZRVBfbEdbgKJxR3FGFKDnUJCt6oIvFDZpGQOOi
hg+2066HXyla/mfocMpAGI7inwYbPAB8u6hjrtjxM4SD8kmPAbz2CXC3+b4TO5bY
`protect END_PROTECTED
