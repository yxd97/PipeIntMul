`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WfU4/ndZThZxq+Rv+IfDNVIJ2OgbKkw6/lYS9/+2+1wwRXPO39THlfKEl84pTAbU
xpupyTZe97jjQq0ELP1c1yZFdqniLEnR/YmzQZ0cT5VTTCtL1CM1pTSFDaQFlSJC
DmakRwISV0wNDEPkbg11e6Igtsr4/sZ/fl8ih1RqYVSQZuHNedEtUG5I5vdbhkbS
0kTkCilaw0dGaGO/0xzonOgTE7jrU9AFY1+ESRea66sznAgqmerjwNAtj+xG86d+
Vcfo/SwS4Aj4DBfJ9uZE+25xkDn1Pa9CGV3wZ/GI6/OvhVrmu8LF/hEtfld8Wsl6
c1bvyLBhuoTTgrAw81lyQFl7JA8AU8yoi9Djr6/hbBQg1eCXsR06CPZR+QECt7cx
FUQSlXH+KYSqI1OCgBVD6u5eHNHIN+ip18b8TUCRxK1LlWJ6a5zNxxfjJ89sYfwO
bXPiqRJRkLOE9Fyjlr6ly5IQtPSzSApNTK5/pr+ug5+qtjguRNxl/sOlBOfcXz0l
rMOEtj9FqfDezMiOZMh+TXIYgNiloXbFHhSmuXc3/dukuaO/uhFYKHN4s9oiVYHz
72YZ3IZ1VjLUZjQOz1iGZ7qfgef/owgJScmdqAgt19nV2W+16oIVtNpmb7krCOUt
K1lI6Tv+yJ1P6kE1ueA0Ja7Ag/3k88mq5VT9jxPfIyRmxUTpndvEuxw0qb9LwNM7
kISDUKy19EsVhOC06qWktLd2dPkG75yg8yGwlWMO+QqB71YUsn70f0KFTtN50ZL+
oOyhjF3BSJ/WIE68yUL19mPQHilSwUb18wW7Nb/m0SI+TVKROVsLg9dE/hfNWH+b
VuBLcloMXc20bsWQ1P/kESv6atpaCZzN8Cqjq6OWD5bXhVvQxOkz83Tkk/y3WSFd
sv78DApCSDrxSTGlqevRhZMNY+vwDh0t/sR7cZ0OS477HVc73Tfte2HPOViGqPCY
4u3W2CeqzohDKxhkrdb4IeQrDd6gBbUTZdefmZoIaImSHmi/OrPcabC3nBbZs0Hw
WAfi6gil6LQrhqMQ6EoIrMe+gZ26OwBnVSnWkvfn69ZVmvrboRx25c2wR3MEjItU
EoJwLspLVrW1jQh2YjAGwETqPwCB8WilOKI0R5jAtqzFW4VodaEGxpZBWF1hhTuU
2XcOGaL3Zz6JJRpLpLmXbi4wsTeUuhT78cjV3C8R8bAaffObooP9ebzyXWAkde45
ZiVEJCgu+2PEcj6qMuQIvpvlwVOoEXewLkLg+cgoU0jTx+GQUquQCYzwRfHZ/S1n
XtscNz6AXV1UEXQpn/7vAIlMYXe8vt0oWbbbHhn/6eN2pGVZJoqICEKcEsxAsnrm
nmHZTz6BI+gO/KCqVwIP9LA7hpkTxFKySSqnqWVHOJY=
`protect END_PROTECTED
