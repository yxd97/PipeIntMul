`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70gpfMAG66/N92hoMG9UGaLsVPjoS55VVadMj+lKpVoeaJCef5rDxaMvYlFHNd6R
/KkgHyTOzy42U3krwPrHGp3tMQ+piVaqpYULkmdnus/I+hx6jphCa0u3FHs0tDQN
rd16A0I29Fujau/YOsTNJDaXzWAO1/FyXrm2D3mNJNK7KL/XgzuktrOhPBPoP6eW
NLQg9FCpCkd+wIeJR4DvbH1W52pjcuwPaKlpXp+1fjhHaI6m4hVUomy6aGAy9w0G
6/n0UsW/LGgskuk1M6yI2k8+FH8gUco8uexL109uPLlSX3fVQ+7ajNVVtwyOoqma
W6n7c3AnPNsPxziPG3b5tg==
`protect END_PROTECTED
