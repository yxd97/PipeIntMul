`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7A+Z55ZK2k/OXIsbqG3HLUASPT0KHlTJs6iZdAF34P7qgCGDpYrPGUreK/86LWJ
PrF+6eUn6kFuQsaNx4o4Ebgeh599a0G/wVypeirl1daVfNo/0SdSS9wzgPWo6v2J
T1hsJI2cM02yLWwYehxt5VtutwXLpBAQsn18cCmKp+zg5NB7OlaCRBRa5wXXRxrZ
lwwcAv1kvEzU4msICfVH0lZQtmY8KNxNn5jfmsqQ9Sxxme30pkeUcN2+V8bu6dGL
L1aK1Sc8Aw6ymVBrgku0k24cgORikKGED5dhKdtpPk6obu4mgs6QdxFgGeZoV8Mr
+18dJD9E2t7Z1ThX5J+Rk1Dftv2dwsUgdXNV3R4AW/ERy6BLZd1EMUVuhIQq8GU9
`protect END_PROTECTED
