`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DNXIaRNq0ZCQ+XnV1cd6H8Lrxwm1Z8ZT0FndVKgqweifqD7iuBgsGT//M+2piABl
fzQtKjAt1qXzoHnP9NVPOuippKX1jS+JvZvNVCxATec3h3EHOm+gD+l6DY9ZdMXj
bIEHETAhOQafgpjtR6hO/O8zwZyT9xxYkK30EAd3cYp40dHjFRmMNxIUzvSngisE
u1+NH0zj04CRGJJfebKvBPlXAxVfFRTzOXMMqfHEJP4jDYJ4sJJeoJNQkBKmrQdv
sgiRql/31NdciKSjIzdr9vMtPXzHK4UFOCkuX5qZOy4=
`protect END_PROTECTED
