`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+vn7PmEZspgwpQaxAWJ67rDg1pqH0syFhZZixM7uY7GvqFaACdjXq+dSEDQAqK/
ZIeOWw3h9k7WeOqUldpzam4gMc3UzgTTI5Xo1/lf8eiw49tBBKSBrpstdKLhNYCK
WIwL30pAImpmiq7asaFYaG4Un0hJeGDSsL7Vor85sCFjYJyRJaZe7NmUjKGPThnR
+h6gYsAL8aECW9rMeEm2B9UFhSuVCQ5xtyxsB2MVQLgxsylKNb5O4TMiZiE7Q7+T
XKwBSfBGqCXZJAkYC2tJMaDlKfUnfaBh7v13EptUSLnCEaPo7F1mipXb89MQG48H
DxhZSubUaahp4a8OzhZsp8MrCMEd2psDhtjbGx+iIR12z2OhL7hSdNJg1ScljknV
xOF4srnOpRu2eymKOZSEm186IRTGNu7oH7qForzm6QJc4wqb2U1vtFmcFwWgH/ZO
BX+Qk+1kwsJryzBk5B6prEKmnWK45S6D0sUs4tOtkaDCryjEGoIvxjj4I2O8UqTP
q/0B665LueZANFxDMjyU68/T8NhCEttlvmDMKXLaWNMew+XvxafoTgfze3F2bNjM
/N4NJ9HhtOE9STryxwEu/MzguIumKTvA11tOg+1kxTR0wz1YQUogl1s0dB1CEslW
DUq0u2IRA753JXkAWEhe7QifbIqsxywojQQnZrTjz+TLWcnVFt6F99lEcXJH52CH
oJPMZN1RuugIPY8VYrB1Oqorx2RcK7HVkajTzQeW9cndw0OFj+txPVcAkbbY8Rg0
U8R14SX0gmQnMcKGGr/8VtOll6JeU2yXG8cQwFAE4lTF0OsEaNd+w0gfHHF+kV6d
eRhfwzWQg0BvdTBeit2Oq0Ihv2tVNfJSwC7tQDOfOn9VJPfOoTpDRlzENr4omoOa
/6KCMtcRGgNjc1Wdlw/xpa2TW+oxsboIDjibyc5HzGU01u6202FxWOeNmBLN2QlJ
ecKY9RkOF98wLh9Ol8EWDwKWeq2MPBxIrCZ/9Hao5eruElavCILspu8k5qTzTWqQ
G4COB1CWqd8xhEdUyKMwB803VNlmloMT3iDd8JV7ioF49rS+4Qqq7csfpDAcBM6r
taXf2e3R4y33KWlCxlXnvmIzIrqqDiI+l+D2EC0mMieDEcKh+CcmI5Ty43cdiPWz
wrAvEd2ZPsnoH7Vwslp67kfqA4X8Q+yz8ceneX3mCOXJGSR1I1aOYEd2T27kSm2a
PLlE8gJbqqPVxwUHAB8XMXTiRi7QlOC/HhXGrNKtpjs2PIESLdRf8N2poB9rJLpX
f2gktc7yGljoI8P8vLlD4RPDwrPuqD2xp3PoviHTYpRwZIaZ+pH47dgiybmS7Zm/
I71EIKkZICDyadnhXZjJU2X7X+knU0Rqkwe9nMU172/uHcJSrEKoN79IUmW7atYm
SIyObk6+Ys0nNmhXtBxBwnT06Qeaeq3j3Po4Klzn/hL8drbt3zb2IJB2G6IMBYtc
/5jipfvjS8/CA5MLf3/djs40tyPKQwO8CEhmfDkh5SlDQdsSzP4s8mP4cxCBt47G
0PDPLVTPqnNbvXUB9rFiw7Ra5CjIv6+0fjCJuxfrb87bej5Y6LyMeh8P5cQ/tnwx
YbrHTGA8S44+ZmPgGv/7NcaPnfc4m9kRk3gODjJcE/gKYYGjLXlCxLSaFly3aJ4c
aZjGCPeXYIln7QV+w28sb5clq3vF7cTY5GlduLwMwSdRPSOJLVeUykx2Pml60rck
fncys/Vs98DeS4W/3FTFVjLJUS0D00/cyPjBcXHnZGhfiJ/dIPfcDLo1U4LH6tR/
ijxb+rSs97xo9enNwnrUZGz2Gvhq2wCufzEjeCQjq/xU+KPJ/FxiVv1HJEsk7tcG
TmKsqRAfUyOOWoQ3wpcnqHkBsIriIQqJjUpPtaWOsk7KQz6YvFRe1nB5nDXgyYBa
/IgUP905yM6pCBZ2cMCWYIgifSQulL399osvIUsPqDFvFkfvu1SoIAY0U3Uvq6+Y
0H4J9cjCwL0qXB6MJA1UAT7Ea8n5b86dr07aJykz5I8lls7vHTsyspd5yuyMNuXu
Mc68pi5fx5QEXCtXByx/8JrC28MMMsZSKwKXC4ovlwZzgv66KGzbfK5A1DMINXtp
CLi9L5rBdEeA5rThHHEhwa+RgiFSsaMrET47votK85Y4YaRHoOyt9T+t02DAbGki
9kPeHf95xU3kkOhOPwYTScO5gqW+ozxNSlEzDbLEG09btBHNvVMlAEu6lCqxog4H
gP3pXdYyGtCridN55ze+sMSErBB9fil8BR2/dsk49sN5FJDgMk/lBRxBzzAC/sAe
iZGgAPkNnOFcjd2Cm8ZdAACmdsRuWOuXkpLPA80U98YngobpwR3wDWX2jJy7yDJI
CeaYmlw6hc8lvht/jvhvpXuX0c2ihTnZzKLKYQMJTUyZdePogpWJS6xdlcNTsQyX
r3AocB4NOHM+dCXFVA4mvM6lYUxl30PFDULn/KnVslKKl7HFLU+YJpmov2juySZm
WSLc6dSpi4Y81QdqesyJO79px7oaulFmkGN0Bw0nfYq6el7bl11fLnHV60IlT2wy
8GbmoVppsg5zTcx1bwDVq8kuToLq0i74qtC5dFoSUQB5lqFcu2T7/KQR7aaLwfWu
ZO9emXTfRVRxOT0xmqothZuuSJbdI4Vqn5dAdLpUuEJp8kWGkgMfg9FR/3Mm76xi
IuFCuaO7wBi/PKBcaBue09E+5GH2NeJAxIJ1zBnX7skzzV9msa6kR538D1dHOE0C
UTOApmuYbi5aUHtg7FX247Ha/K7adxLlF+SCilmSx4DcingBrFE4SXB6ZRz6EdvV
hVyVYeWwW2EIuoxvLmEHKYBeC3rQeKC491PrP5VSZOfLKsN8dUBmx6ZzRywE9Bpb
rbkavzERqM/gzmLV5DV3ljAMrM0vrx3ofqGPGaZIdSxtKbk2SDXua9bUh2EvxXfV
BwOUuRRkXSZxigXwIEq14sEf0JmbdgRGpP2tZnljdfVQMJ2YlFYlDWrvidRuZES4
dgpYTNj46osUaEPmqN7xHM47poTX9OBsBHfYnLzzwUlE4sirGUyEvoR0OpM2MMUO
ymkyEoCG6+yUmry7++WF19mciywm8vQedZvfIdzIsD1L0+GkzQZixhsgHkXXBax3
3ypEGcehphVMjdTJa1kWXi79dXkfNlN/5fO9lsVuBw26uEXwVlE5Pahvyz/QVPt8
JRc+RbX9gDTFLvp17VbucZwP5myz8CBZ5MYeZqfEU3daUN3Hxi2J2aG/d9BdBq/v
o2d7xe3RxvOsd45I9+Twy9TOLwkgOOGwplOLfkOgGllopICT4lqgJtWFv0k6ywSL
DMAo+pLjuygQtg/lxpNxnYWJj/h4QCKMPistnRs8uQFI1zFaHCnq88l0spjjZ3G+
eRYNC51QUwF1/LnmJXqWR7fy3Ub7UQgc51aK5V3zZoFlM76MyBsfkpCeiZqMMTo2
5qC9Kc8QzoLkTp6W4NMhxyNe6jiBTlwCFwWr+09Pko6WD+K92giPwrPV7wSTYy3n
ccLSkQ4fBKPvzDDQZwcAwVeB4v+KWJUVUmbxymx9IMJps+9LSF9pziyTkuakSyVz
/LXEN4HkhX8PVntw3TPChXKKkptPKQ2MZq+o+86n/HK/nd9i+wI6GyblnI8RpF2n
e+Te4ZiOAngifsfaGInmtEzcEI/3E0kKp+w3cJuG4jJ6Rho2JFSXuQILuIbM06h8
RyccCdxU5aDcYxUKwOmgubvuLoFFG3A0jqAjverPdhZtQb74C3/na7OHejSCrSyr
j8WKsc+XV6d3cnkOyx4K4PcTXWidJ5WkR089vO6gpG8ktEOZ4oJ9baUT5znz87YF
y7fVGa4ZcJBgzT3XpaQQNuULTv+txSD4CuzZ3FmMYuAnKIQAqaY8tAg3LJ5RZ4Na
uIcHTIGhLh7+lsuKo+TEveKtJgCABdwGgVsiKO9HecNdH6y1b1bfRxgyfiUEmYVN
FZhnEa9eHSGJfmYcmYV/uyuvU6++lEEotSesWbzbSa9ECXK9IB37m9Dd6+IMRCwX
jtZIxCa7/ZVoj5rmZSR3Jh21RSWyVD8H4ISsuiYYIGyigEhJKcy+Udw3YumC/NHH
QwEiXqpOfimBvcsAq+XZI4vdi43TOC2LVTt/W0jQO0xpY961N1FtsJTh6EVSBamL
Cm3vTAx+2Rq5J8aTsGImrMXss5DplBINGyTEOR9W7l2JA9g8y0RWot3qj0+yPOH+
WfqnWqYymcJhTv7Bx93PVCStuGNNGI1XgGh8uKhJh9M6tqXhdGFTOwr7jV0kWGqk
DPvkOOV22O/LGs6e1MgN8mnGIO6VJWKTOAy4oLIEw6tz7kx7DPJGepDre8uwt/Zw
7qFCtHRtZNJCNICw7SQDRNEy/APT9kAa4Fvxga7jTXwCzMmoM19wDTvYZcmZHuf4
uT8tCs02BjrFJD7S4ynLLmNOZDdCltH3pYetu6gwM78yUjraI8xZEFCTWFGYRZ7O
F9fQce2WWJrt5VrtyIrDDmVmlmYLNjwn8pzgnzFFK1KpG3b5/y2Wmf8QrXFkA0OX
PKOfFAgsKMffoooNkne0HEBSXTKetfzMgfTN/++coXPZnIBK9e9WY94K3JSbT4Mj
8xGaluJUBHTYqrwks7TjfjOUW0QPRuL3xSub7Vaji3gTPH71K5Wu3z0pWTukJQF5
HV2eKKbJRBa0Ojyod6B17Jal+PvPi+nMHQDIhxMVrf652IbmH8Vb5Pqh6kDQ/XY5
4pRtQzNNq/zTLlO/MpBenuDaJIIdICkVHa16LlyPcbcv/A+n9xsRrzRTz1QRxM0b
OK7h+lSXDyM8zhyvZ4PQAi2vL5WZ61QwZQXOE6MdgroiyuPcCIU21DmK0yRLECby
wlOeKaVvYrZqF1cI4PKc554irIcYkbBdaPBu4ygE0tUdmOp6qJLaX2KUDyLkcKuY
FWoBL5wgerCuKVrgnIpcKpPdVFinQqlP9oAuGFXa6xg0DkaonZ+gCR9S+G73gfjS
Pn1ekslkNfDB3lA9HpUCzrlgjNPjQ/37OhFcfA8sYe+x2+v36RN25PKPKOJwQhEp
Te+Xomv5mRjaM8rySHM0wSl29LypJZU/j/6Xz5nuyzFawXFxGxfM6+/zOywR/NRc
yD7StvIzxu0bN5oKI/3qWbbwn5PmevD7Sa64xr7LEtMqekSo5I6Rj9J1H9O05hrJ
ESOVgH3HFiuhJKbod4AUuSKG7gfY5KK7FkqD15u64Iprg/m52Nyf5zkM2nBj8iMY
csoaYqK5Vn3Y/cJA6EmOitZCtRs+00bJBRYz+WsnrYcLB2LTKUIDgpPIl4NOttdd
BiJ0SyhYk9lsonOsCfowbghen/fWoY6aueIdvHeV10/HOXqjfVZMqaZUhFUFS8eQ
bFVC29JtVUi9RaIZHN2rQdJdig1ap2b+WWzSBTQyzDvnc2Y4adlBzrD/wVOeiYVc
/N+3bMKgauy1IP5kjkI4WTv7Hw6hvQzaR8ct4NFZJ7D5FNS1PhxSIgNBbyFtFv3F
UuN1t5m0of4qtnw76m72spmUpdLamQRd60tS4gEpA80vjazje9WAQo4nbXoRzHHs
l2UExRO+WlasOEfVMfHZyt0PGpNxQoeSNP1cXv1loT6Y9JiGDT6u2D08MQRvJ0Y2
gMXFqWt+fWNNbRnXdhyouK7JyVnduM8HswCJIBLeAXX+gSKgFKEXlQx2eVbbjQ+a
1cXbNM6OTRlo1tHj3VLiKwUMj9N8wG2u/xrQl63dg323D8K/56nEfem9oHm0kCp6
vYvksWUteIctU2LS7xKwHs1iC7SRB0/jViF3/LhRHujQWrfdeJxNyMiMq2tUtHI/
3kNeYFLfnOxE4pgdiFLhYD+jE1ctu3UYv7/fECZc7OjwRISQiM/NjRBuf+AMH0DF
Hy1+m7Zwq/eEl30ADBdOYA1UHdJptn3uWXcE4LcA+kbm9iWak71JCgQA6MKS7cI3
2HC5sQXo5PoVZUuwoKwwgpVIpnM6ChLOIP25NmxFm2fDvme6iYwyd/RT8ejwWiXM
VSxjdVDNc10Ber5U0QWz+sTWTnjJsv2SUUFwkaPSfrw3+edIDJ/x961GexnGQTan
NnSK26pyE1FYkFIYvqMKbD2kXxT4C7BQkp2IXWjN1Y7CvIEpzfR6aRq7Zz0nlqDy
bRrDjeYYSKHojn+mOF6DjIhEcYqMCQhyP7Affgt8I5tN5M462j2SSjyYa43+7Sct
1oaM5Wyl93LDoh0m5byuCxRMKf6LZC65Evc8gOrLthUlFoNwum9/r4mK5zVA4Woy
21mzWa2p2qQrpXWHYWdhfaiSkizBZjCX/Hj7lMyDVRZXloLEXyZNI/aJmCZnkfUR
MKwco8/yYovh5a3ZtUXeOxAR1QdyFLE28SpJLFxbqUu9RfoTuPUsezwRiD5PzmQc
tHvX0D3DUu+cklerMwXI72BXj+1dK5zm5FUMwEIlJ5lBAJnwO5aVYeSVXztAh+TI
M7E9JYOJwqVvvIKuzczpT1Vnq2+Quj5mP+Q0jcBsI6z5TCz2sux30rF67x1Bl18w
PaO9YYo/bEI2XPsdTWKMGNo9JJklbn2NpaQg1id0IYQHgiDgnhG4py3a/4yGh4RQ
8jsXxIhN7BSlkgl50uUokJ8kGt1bXieFEbs6VMtzg411fTzr/utQGiEE5U9ElmSz
NRw+CxmcL+um4iW/w0RL4JIVUluVQEqSICOyHKtm8xgxu7cCfhVRbGa3uT1Dwe3u
5az3eia+iA6Lslabi4wwjvWI4Dw9gFJfCslXJKUBOZBfQVkPHLJzKjQi1EEm9huY
fBYrgr8eO1qembHM2SG1P+OYvUi70l0mptFvtPpDTeNMkyUebV+np6zTWW4l8FHs
U2IuuhTIStuk8Ic2eSWJWok/CNg3MaSZ+8gB+cLaeHWe0j0la+MP7oU1cwMwcbcf
WS1wtuqe1FTNp00oGXXIgxrWwGIBVbUlbQAnhst71Ihnc27kSFA2yhXG+S55y3RA
CPaL9bu7zyEjpTaRV1T+hrx/YhFdKDmmh5A9f7G9n7erWIkj+D7vAig0RwaRC+tH
vWHYJKIM1HRj9tVNY/gGOPHQ9kQmfBsuhtu6Ol3HNDnYiUmXufWEhvs0BJuJkrMf
DdS90mzjrSwqJ8KYk4Url7C0dDPQM2iIN8KPMsSAaK+HGfttHgoQkZsX029ljFND
ygp3I7r0x40yI5k8mCURn9rBMtccU8cDwIoLfu5lua2E9em9+ziaAaHv2kuA3bpK
9MQL1bmBU7MiJBym+YFVwLa2XcDkb6wwBevNH/RUVKPk4wdcILDgdvBlzAkw2MNp
XBK8Aud6mRRv2ZG0mCDjly6Cof38x4ImVUPpW5GI+z7XpIWdWsE69Di0yZ6OKMDN
CqmAve2F689FGn8hm0QpytSD+G/JO2sQkoQ1M3XZHIfX3gWpFCbMGQ3QIBofBAR1
wjeWudpuQYtdwyp6oIfQxuDTANTUIFW3NccPzKq+nnbdlhLP00UfcYGXLUk1DtLr
2fjGg4VIAQIT57homcjjN0LU4WoKg8aggytnbaIQ9xUoRp+RUMBooQ7MMLg8fO9y
NEg4EcKDC2mz1qFT8J1fPD0W7I4VgdAV+MKmV0LNX3KYOy/uH608/PA8TyCNxpvC
EU2c9g1nY5oWdaa94wAz0KDy5yycqAatAUt2niIYdHV3aEEhTIgqwLq9NKgfIatT
SyRCwWr9NAn2n3EIl7b8x3bvma4q8ZOGitQ60bj+hVFfiEq8XqKBy2RgIfyfaOoC
FqUt0MZ6YcLqyPCxxmynLpMXRO83M97zpu9c2LWJX5108JQosknk3t6gxgtC7q18
Hn68Ggn3uNvrVKFjTAe3yRjD9vF0fagAyRLwVIf3zt33i56ZK4FIFcnUbio/c/Dt
59j2A0H7EhVZB5JzAALsxIFE4SB5vvA2Nl22xSSdAapII0cuXEk9ahSpMx2M+VAC
yAnfginfI+DPKSbefYowLZP8Kkxga2iRTkFEmJq54UfJlzHXPea0bpHVt3MR8WYa
5gLo33+pxL3DAnZzdU4KE2jEbK1+Z8VvBgZSAk1fVjyQKVfDRcUGFPZBfLmI0nX0
AJxJoFyYur7LX9kC/VoM5dV3HQBBNjU5QwxYvxDtt109KCjYXHgQHEQrf2kh4UGb
oCkZwhZXvzTI+YY8jiF4dDt7B+V4EgpK5/3+eCHJgV9ix8ZJoKrhyZYAXvTKU1q4
Oiu8/D8+YrXhFRt3qM61Ib+tGZ2VuHxIGiq9dgs0LZtK+hYCYf2N36ZJEK/J0+MK
MQ4mMxN7TMsHqcbfQgLEZ6mTUfgqKGMGVowSncxDYjVl9Ur500pYooSfIhVRO+F6
WiK3JErKJRg8xnCHcpy+sTpomXbetVMpK7gMbB7U7pRiwbYM0J5nKKD8fZ2yvliq
ar+vaGE2LROGpN20fGTr3s7Vtv1uVVWhr9/ZS/FReKGuw0yMj4Lg2aXRf4q4T7+G
ZRYHaX4XVNJK9+/2RJzdmjyiCF7WWJDmRwL2hGVxgzom16ASpaYQssoTD+uExa7S
EPAYdiD2z7jlE7Ah6zdhZJxTj9to1y3/5UgW7VcMVdV4ViMNWv8nLkMPKPsDen9/
vGTzemiUqptlsHEd1MZj48FxEvxIPHMi8ZHdbqRHOUvmH17ecjY5QcnLmthdklkM
uQd75pogYxH859JL6fM992BBflJdVe3V2acQr/r8sIZLPSUiSt+rTp+2SCtZiC1w
TiI8enX39NLXLnRdys3BZQpgUMB/c/t6c/2sRWCbkUhUTGQc8ROwz0mQH+AbmJbE
9KTjTgFVr9zaPIBXtmxp1XPxap7tz72QFrFoFzod+lJkdpkju13HZlDbKzjyvVBI
1SEx0qkdbK9yxJeTn4S6SXeOkrGLbMiBlj0pwzVKsXNgpTOxuvS5VeDtr5F3DBT9
e0OogfUEDkaG/1krM9uW+zdDgaTGPNay73+g473XaumZI3kRM8d1DgWqpNJzNN6F
lsq/4s2Nso2hV6RMclrpsUHy6tatnzxL/uBOTeXiswOn38/esOaZu2RkqHOBLrbq
G92lDDvt4ir4gDJGXJj2gS1ScvdzJ2JwgfaUkTHaQE72bFfmuxuBFk0iHlWznnFj
OP5SHL73l7jA7CVqftaKduNMKK5pScc0MRdSoYR6gQW56WZFedvDPcPeEwllFza/
SJBcksDPiDh+MqdG2YtWb5Kr72NunTWJu1Q7rLzbV0acHOgXbeLll/w3yEp6Rr/D
z0DnsFllkK6Z1wcS6e+Rb8NOCGQ97uC+IHcg/1JBShaYkfBfQYUdQgZzW9ELdW7I
ZSfIpuAkGcyGfwKyXJkqgrMofyMpO2z9oX003pB6utFaXvQ/6q094lTfJU1PlUwM
OFfwSZ0zzVhqJ7LNEVOwDNLeWbsWCMgOcKDBT81Vo89BxR7XR6oAbyJFNHc62Nxz
umfFfV8YcTwCZMmh+yBPKfLY2Twg9qy+XBBMtLl1MGjBctDdvivEuCP+lPogKItn
+4rarFPAMgBcAhAUsSpwAPc5Qa7m3+iGTmsEvXE7Yi5U3WPR3j/VLRN7Ab1mqC/D
4kn2Ow94RQZqhvWVfmG8f6shDYkH2BLXI6v8yC39DK3NNQ0MMe0jq9/0sJ6KRR2p
yR/DafdkjRwVo5Hzl9ahVOorjd/EhbreXCHpaLqYsxsu2Ddhtp0IVo8MgI2DUKKd
O4WbdoFJW7rRgCG64dU38bhTjbU6MbYXSQkWkbsnR8F+/EQBwUCj3tVFr2Jbc3D7
T9kMKd4X1tJBS744KUsgcyDzARVwx/m4pZXhjEtx2DVAkdNF8PRmqPy70MzS7XC4
HkQq/qvQNcKCyRchYhWdRnUS2wWdcLqtEx7Hi2F29w64WST5YRrGBVgxWAfT3xG9
3kSOqAzlin4gKQ4bvSq/qWqWJ0G9PbGcgOEP9vjEyUSN1bdNtEfr661Wzunud5JJ
HVlq4wsXGhUnP559XRzL6xcqSykf52fOaRIqSTJInCjwQIZQ/e5DieCu/4Qtgqqf
rcXen+ntHwQbDK/ZaYPQJ0miXDSJWgLQ+qABKiKZ1OaP/TLLj1FDsa+M8oGGkg45
llmXx3RNgPnz9fFbKoQIwIfXzI6KgTCRSM9FeJcNx3/R5hcYYsg1wvau5zm7RFUV
bQOEugNBWkTpOfNFIRiDGNVYXBV3WI76XvlBlZT27+w3Aa6bJdMClo0iFESYgTb2
UmBao07ILpXpdEEj1/VsYjrqtwfhEMRQEZCGMaUE4acvII4CmkImVyfpovuTpKTa
leFWrfAWoa+EsZxOQD9No3ojVScldCGH51pRJkS/xPDBFDTOKb+U51nYOsTYra0M
eaJUoD2GBeWQSlX3HGTjAtLWBA84R9DEQS178p4DGvnnUymJWJ7Ls54+xK6u9IA4
7MjVebBHPQtUn8/UTDZze2IdBpHVBFiy/riZMtzqSRrhxHwC80265pVMv3kT0Elp
ilJ6zsrbYk5opXjFqaJhNcxDWuIHHKJ70drEeWOZr5Hc4duV9KmEM3Qj7WJCotpI
8V2LUOeo6IGdtITh4liABmw5VdWs8qJdkYJXN/giyqVWalqHAreQ3cG2g/a6PgI1
e8zl6cxjpyc5XjK9+j3PPjkqo7KZ7jHlsxMB249kwqThq3+RYymfzVNWJ2KYkFgk
9di3soFb/QQU0Y+c/oyTnSVUT7I6E0PUahDZO1aR1bYZhozFfY9UHsAUMo7Egy1p
YtNooubV3SVdzzCvwhnVmSMVh1BojjDrUAXrKspGW3D9Dt8iL6yT4RUqNSRW9lXF
gAMw3K12A3tDMAy/bkgzC1SE6qs/DEN1IITfVAF7kEZD+wfow9WrIlBjGY9y9s2a
jMHCmjiqwFaAhq97Isaa0Shx8qpgzEPGrdQ3LRqd/UO7HCIDh60Ihg1UK/jzGO4U
su0lkoj4PwNA+EurOpOedW6LYZJEB5zoaM7/T498oTBL+i+Oz4uE6rZY6nAS5LqR
VqnjHiySUxi0wP8xoD/JvaJIltxbf9NEod1R7GxkDbfjsfR+hgNAd0QO6HauDgjv
tTj+wnzSiQynEngPXsFs5vutZ4H61yFb0VY6I4mxxKnIYHv1u/Tz2wHmc1NpNWGi
pftGW8nXpx+FZeggiefW2AOBYrMxyEx5UOLSTvB3GLfZR7DVOD8bscE3X0IgCthB
TdQNvCvpvbcucNHZEkf+eBF6cfz7EN+4foE5FSMA9ZP3fdpQM63TAtvniUItX9Rc
lEJdLvYVorcWNRK+4PGfZJQQFQMAncBphr8wPmbg52NWLRjvStcqZECPuiF2TOJF
cb/9PNZ/u5xw6ebKNUGRlUDPIXXoVKVH5OqLKT2yI0J2qgg0E+iH7VRYK6GgqJbM
E6yaBp84cSTjTfk8MbwW+ZKuE3zUij9HPQkmU0h3ftn/wVpTE/Srtc0sTMeUwGyj
WbUVBMSDL4qBN/qSy6Jx69Xydn7nPYBYj+jYlma0E8jSBKE+mOMI1comag6Cw+VJ
jVBDPWgjlBHB+EaVsoTN4tF4bthHoYcR9gFuaGSb7LfeFIxB/8TBbnUEtBryu/Ua
rBmqjzQEefgaTb9KC4EgIE8WD3UOXFRd+HH/Y2vIZOqNWAEwx8Mp0zM0y77OAd6j
k+7vGl/kayugpWgsFThfSB3+caKhmbG+xzEYhc7ZN3ZkWDiPoA2bIferimiI9Rc3
u3dIIf7orGTTmaOLjejkKRPw0WMrAwsymVjndAbqusAcb0ddrTc/DdkCNrFhTcsX
YAMb82XSK3mg75MojLNuis1TPwRMmiAz0fqKT93UMCQl1E/w2KzCfjacQfzPwu2z
M/HBKG9awKLXv7OJrCbnAPErFOjoEpxdooCzIj5cRIXlkm8Tpna/U5GOTic4z8NJ
GfmTODv8G89+lyvcKW+NgFS/6kSp2+vhC7FzzGlYWgW6Kxk+QWoNPbEsYfoBVsLm
QyPKVFupUypJ0gMfODQXL+EA65nxXmJjELFdP2nJd7iqMxDPx2wPpSYD8gODOEwB
uBRdFICS4qRiANfWTjiwh4i/FwIfEENOjRTnfsPQz0hD5UDbXAfJzyCFNKeXaPfO
/VHZVoqfK6lUC05iLfsOalMlF39qPtOBDVVxlie5NUgOMBVehv/sUVw6VIjesSp8
BFG84Q1icnKkcv87pOpmiXoNHGkjKRJMaNC4p24znmTz0GqR0G06maPAmLThC+gW
rd5/uN0lFJn6bEt90GSIr4dOgkQYfiVL5gJFwkAn3zotvtV6PYFbrlp89e2XZkq5
8Q3MDC7EcOM6Q62sBEJVnsJ4APx+JuJ0QgQOrzxOaN4m7L5nlCWIdh4CX8sVApu8
aiKysgWVemQqJ0MWHUyBj4uOuyd+d2yffwcXv/bqY553DAa003MZTziilWkOeWAj
VKniuJqRKCKKABVot1T+csLk5nU50EDx3t58SVputGzEhHI1uBjuz8YakazMrF3K
cXKXCy6kSjNuDXMEw4JGVr1ZlcEEPVAdJaBjYc4Ux4j6r1uV0rx6GXisoF1xRzwu
gW+XYgnGHp4JJzNE1ReFtoaZLbbGhQkQhPMsSIl1G4MaydRTfOBNL29HOanBP4AT
Jb7CC/SwbAoX3SfJTBw/qTbL7L9CSFDN9465blXu33DwsCcURRPZoekKdT7b43qQ
p3zq0vjWV4nOJU/qi17fta9eLxWA0wTpMlfJ6y734CMXRZH4wzu+XVmPnWDo68+8
Hu3y5iFD2NVWFg1FNs7K56H6evILKdcxlhfBbm0UjemZm5r61+sCxfe5pkRxVqHe
iZ0BszAbfkb/dQ90nwGhBPD8f1oLtzOrNRfxMdgz8Al43Y8IL/J5pulOW7Cy3yzw
uxGOt6+A2t/zu7H44t4EEPpqnvoeSr1xvtGKZ1fv4Sxd2e74+tkdhsa0RgNdX9Y0
IxMxXDvTb9oE+WKQR+M78Pdr3nmEMJqsOOsbQgV7mWC9L5l2H0a5AzU5DX4GwR6D
xKdYJzkBdUUj1jhKFbhjkYSuEpDeTkbH1JZrmHlRls97L1Kqwq/38+xO9yE2Mii2
dn1nEh4OhbtvUn7NKuo3ZSqCUY/IPUAQA9R+meWfVYfcJgnQyxOuE1zwXcXB/Oad
Ol+HMJWvPnti3al0KoOgTUuaSJGNf/WXhfeHv5/sENfjAOAwqqzVlgKh9rwZD4W/
5OjuxprihznLnpvDsTJHeWWqqkf7oPrVi6YG0C/Lmx+ZKuiDolB66/b06ihpzYMr
BvDGVnDqE4IEtlY1jBxehmtIEFQPcwOZG10P1OuEt5cJwSyO1hBYPMG9sDuhoQW3
8Omz68wvnGMHOgG2oOXk7GTVa7GZBSiqhgEl1YTRBrjSADmbZDjKur2YL75OlyRw
FiamoVs0d9BhTFLi70do84sqzr9zS9hOrxHMeO1CM5t3XuEEcUtA9rNTt+mwGM/Q
A9GkA8lytK3S96Xh3zrE6tWzitYPJ2uaA+LgNPbAoS56cKD7FJZdVkdX8wIb8FBz
x1YXwtQyNycLKXbWCQ4QA1fqtbXnc/vh3I44+byc6voMD6E4/3C98KFRYwvrrxQB
QSZJQQ+WcqvUO8EdBzM98/Hs1Pi8bNHGWhghJ5xFBSDpIR6a2zd7Ps0qAfLBkRNf
9fN1tiMM6vOsKDO7krOjXyQvOdAbQSIqPIo62Z/d0sUVKU7xuNosl0qzKv9dB7SU
Zb2WQBeu+r/TV+v5ceLOXgtRzln/oBM0117woEJzZ3Ngy5VABMXcXDkQld2ETXz9
5qsOc8ejml8lmjjkpcelsd9PvgOtv4tR9YuzsE0wTOG0hORdAJa/ox24qzHneLe1
7dcz9j6lcUhGOGWT1SKdC7knDPmrTwGAr2o0R3pkA5zosGCqZj6u01J9pDG+LAZM
VfzhEdaFpeJ2ZEajtSX4vs5DpIWMdoIkIzBB1NGj/V4t2gn40+aHbUf0UCL1CMUZ
XRtyxHXP/iJad8hPRvgYJmQX+snxDnYlsQXNfXpXqnrh6WjED++n4rVVmpHrNhb3
+e4oCrM6oNerwNsLEB0tvPUzXkVHdMeIMbsMzaQ88hixhtalxrwaCCfRHm/AwGBR
g9ZxWXciD6OoXqQjB6gpsxrxnrovLf2fRgZUkOqnR799ZmalvTdTd5QVbA3D1PRA
GBdg835L3pQGLyTCtfZrSaEL/Q1I5maxE+PrrSQT2xiw+2swmxBh2dETvqTgmdKq
Y09ZCgJ1EpwEhHsSMBLsifvkz8xjbFoY9tArpld2pHMirighIT8YICvIp7QA3abz
vNeogQCTFqwzjqqVPkmu7fxQXVG6+do2WQl43ZqzughpCzlfOcAUnWVcyQGbiITB
Oj3+P/oJLhbTPSswlOU/Zu3dc+obb2hklRWj1tPvimfICj+a8zs6ZGsUVI/v6cly
zPaiajfGic9lp22JK/W/Xvux5Ouv39md13qC0grxmVWb+aYWaSWVK6DLPVyPOMG5
MgahgGPM4Kz+gr6FAzKPlAy6WH8OX84cJ4RP0PthqD8cMS0J5y60aoNDqtNibIod
y4uzmSdlzctBjvHZpyte5+hEyVHke6XQLGyGvl/QH+TsmE7nIQN+zfidV79vmqTj
3/Iv/LCwpzCbb+LofGnZPOxNK3d3uNR4yGx3dmzzSk/wGGH/484324QdUJwKlueL
BSvYyZbjE1DsFgwmJ5crTwylU90R9LCGdsr8xLrtxAcaPDSnY1sZvfwk0shcqTpT
k9VBiuNm7uaIQbV3N14FKDfrvbEJQnU/oiPfgsm0KZxwbsS2NDhCP1XheEYnDOlb
eXDEwcvB+4ZDwlFX7kaVLmmZ9hXrMmd5k8Do3VX8luQrxxD+KyVLQTLxISablLHU
O2+ZLwOZaq+kl8MCGoG6IlPgJDXj6hoILxO7grEFlPSH2CfTfDKlMO8Ih57+OYXO
Y9RgJMHMh3cAl66tQnvDHP5vFmDt/pVZzzAPBTmZ1oStVz9otu9/1IevPJo6TjRN
r5Ur8qAMfw359flJvOXfAkIm44vxaXycxRLNc2nlJlIY+c/ahu1TZxXoESPCmlrJ
FHOY8UatdshP1KE4GEwcDjjnWwpeOnMYT62LvLEdePgUAhqGSbuEPw6DPEliEtyp
oLXZAbTm9491/uGI+vg1QmUb3hc2kI8IjGQVhLRWaUWYu6YSUBAr25R1QxpuGkEb
WnBTcJC+AUXcQO0EkH3jCU43h+mvbBjKHArxJ2ks+Y397DgL7QSZXGFQq6hEkKkX
UeY3K2VZItZ4m+NEunPPS761erakWVELd0/nqeXvhfI107IpPLprF/enXvFFYVbR
zRvdFZOUXVE/fizRN4IsohXfCldYzKeIIyRlQjr+6EKcSCSXh88Ry9xxxaf/TzVM
LM/YbmZ4B6C6IhNsd4yjloD8lEkt8SkBFA7k5fvz6yq2Vm8rY30YWIDxtdyqdrNn
w3BY/quJ6cYo5qYrBqpQVMAkhqAXJKIe9VsFaGZSpCxoY+dyhmbakhwUaY5WKqIO
2V6wAe/UlnvrLFOu6Cgd3oCUR+53EydrKZCoOENaNUfrhu7XdADNOj/MaLeqDW5Q
T3FMqIei8/lvxkmoBwO0xx59m41Dl2gKAvzUz9fhLiVQgmRtIQPKvuasxN+LFvUz
0rcY75C/yFQ0YL6894HlH9/6n0nRtp5hW5mrOzbSaBIPiMeKK4oKudpmFnZMf6AH
8VAwGeI1GnlBa5tVTAlPZLy7wkBEfq1CJo36r1Pa2lMKccRKGbbmlRAO3YBug3dH
4SC4htZ4AHEFiPGaEbvYE222Wl1uVe9LzB9obpRHv4ZBpCfOyWk2UFXkHRkZv/I4
hT13gKbMlHdx5uLV52FS283T4bDkrQXQHkviGUUSYG+Lc2RyImirwfacjZisIW5W
HGsKx+1iu7/nvtzjBcO/gZvZ2J93J81kB/k/qqtanLWYOp3sQHN78/Hv611YeXny
jyVDeH2LxscjekEYaBqw1ooKRLyk+hfNsCXj3HkkektqU03Yck2zKNBbffKzcNWH
ptLtHsAW7AN7fxKGKyFGwE0L2ImGQCkSeWIEzBnWOYZTXpdATFflGaOy66dmdatZ
CJZ60UgEOFnV1XitiC3aMW38kCJFbBMVtjYu5zwpSNM8A/jKfDrVDb0XuCCKkPcY
Xjt+d2vsVZbPq9zH1tos4T6ILIkoJ7h/J+H8WDHLzlQy+o8/+mvaES65o3Lf9DzE
RSnfPiuEiKKDeKbBofdUrfxrlK9DTdTnmh2LAu8d9i+Z2ncFGhsEOWThOz4rKb7u
DXwE5R85eO0DPacG6mPsq3wi0SuQCghgMStTkLIopegjk3FpDIzQ8VEza0whtDhw
6sHCx87W2qVGju34OiwL3ul7MI8ozrSTVkJ49PaoXP6twNPwx5KfTCcZ9gJ8yEqY
4DIYwPXlGl8a62j1VsTuv/LFfyLlqZQLI97UpCCQEEOlMk+CzQYn6+PZfLXf+Sw8
DC1+4yHqSwK9cv36cRiSxS4fqrAOO7XpKcqA/hLCaHmb4in3nFW3g6uaSFvrVGl2
7sy/hldbu6/9GNoRIcf1m6IyPJCqjNWD9cfQQp2oUj6GOqCusMAT08or4FN84FZ8
i8tPt9qsj4tYxd/PWO/TvKl3iRTxY22Vapv9nsLZR/Z974W/D22Mr1lftrxZmrfW
nug4uWpzpC+pLeLF/hSguoBueDI3R6ZFu/0sPdnrYx9L9A2JfEiaMKLuJ+1rEDqr
zZbcfim14dmFAonqR0S9UseRF2mWv1Abno5AhqxzFjziKDNoF+IAywQFHmNuUqdb
acKm2Qs7U0fpu8bjBi//Ld+PD19MZXfLkC9+l05PucXu+0OPu2CyJvn+WeVD5HaP
vBTBBCXvA4bq/3Be9c6bFU5YhgzBzEFMadYB1hHLpbpnDbb75Lu9pGfh99WZirmv
8A4xjsldZnvKJ18HaquSpSsHDQWXOV051UDD7Sz9ltrrZpXxTPbNc2jAB3SR3RK0
N2cZ8u7XMNZFCwCQT8OlTv98Gud1O/9ALaUBzbVqJTuObE9UuqBKiFMOjfO8GQVu
aFBcwpOothkkP0OnXB8eJyF8r5I0oBPMghnO9MPj5b6mESIlfyIH9gNjw7v0QGWG
pdkbwX9FEakL8IvoJn47jPMU44vfKgLpFoSLotSwcIpgwNQPMNeZIbLzveoSAhQ1
tqp4jOcUjKBc1hmwoC7sCFgVXpxV7ITOrByovEosNOURQIGXjcvoCfc7Puzyd+g0
y3m+BfX+gRCpHJ+GnfZ1cS77NmvmiK0xj9BGI+dhF/Xh/th5jPh6beIMnw9tWeF2
seq8l7r0SDTCLrr/6x2esVjL4KFPe4cXpTvDyP70lutt7gVu4B5+BhV3hrA2AADJ
uFjBsKGGE7JroUHldo/7xoLX5ASghopsCMMsP4+bG3Ka1mNoirms0JTFerJoyUNF
tYOH4HPcp+3ISdVA8k6p5OAtQVAGQB4WJUfo3DAGESe3IABkF7N5O3pPUuwTd6dG
D/iTFpI2xHKcvNj4x4l3snsSxwjG8dcV6OQOLgnv9nzvlbuEX6EhWMGcvfVFrrSB
l9u+lyefMjf2McrX6fqFZbUpYJ3Q9CAsLW46PShmnh9LGf5y5nasA+mbTnPnucD/
Ya0to0mJ3sGCG1kQ7ltrN7QXvJwkSLmEYtKOAxcjqJOr307UelFESJ2ug+qWFlEp
sTMC/r5C4dOAgV0xTywveZTjZlBAGgGuG9/aLH1Z+BOS92FadaK7GUjqlpf/lwjF
GMAIJhejTVHQ7MVL9cMAxJGdI7v+wnOZzInusUYiA0cnFI2MTLUEXXZa7T/fMO42
5bf3iNsmmoFq1C6/X4GbOhnONZr+qd/iYnrpPoCMb7NmQQY5HdWPuVlaHIcc2aEm
du5Vzy3m4WK5E7Ir1D6Jaol1iSTjuF21nYBxXuYb4VWtLg0rdEg0+UQJPzgkaypE
O33LGDbq7LNT+UAP819+5rxFLxBv/b3zIvn7TZyYWAfeYdWzdKFam6gRrrOL0UZA
ZRG3yIzJM/UX7NAO0GEresfFbQsEjs57DizBLkAnW6FdpkfwZej/sqmf0A0iMklH
42z3PEa42wbWA+R0PeM1RLhN0/Xcd43YyfiUQ85tby79hXYu39mCJqnoMKWAnWAL
//j4acpCZwAmFsN5P+RbCJ9ILN6+w2ae2I13xhdTsTqG/ErUVO+YOHPWPSAom9+L
9QL6tV8G0rUARwZb7EYwsS4atk8g0xljuNht1S26JOIgSUKj6jm6ZeMqsMonG1BG
mkolf+MasYsyGlk+q4FoZGSG3cJuU7yEVFfqt5sCVaFWfVPccMOw0daYcvy+yO17
gQgaFLRQGTkMhWucukjbUlaCvZkIpwiWZ+1c7ZEmQT63bWBWsZmAVVXe8RbB0sLf
J92zVv73XVKiNQ22UdwAS5IWCd1IR17kRr0lnMq2VHCaf9qE60bIVxgN90c1nW2m
cOae9gqmgc90X6qH5hFUBao6muT6Rt4bonIKj7DmZ8mXCBuJzYlMjNL/1WFHlbJo
9EhvGmqKs2tURBeYYtsgfGKhHW4zLDkese7Xx0C2v/9YNi+XJOWgUNKnaA0mwy3y
7sliecTetYlvou3A4wfw0dy3cBmJXRDuRnZhdnEh4WMAThOQKVF75eSgpe+xxaJz
E55Z5OiPUrABMapRVnDPuSKHAq7IHiT5kvqGFLe46GL+4uqGdlyPz18vwjSle7w5
QSDWsUzUsxxp/+nUiT76Py5w+N0G2DAHgJBsb1StsK2ArXMndhvv6+vi4bHAemm5
lkkt8jlNsL+X/JNqCwnHwFs1ThvVBuDv8c5bCq+kovV6MRCAzqiijcnfc5vr9gUQ
du+b4skqgg4cvVBLO6WYwCqx1Fgm0DaijiiQUchFl6idSY0yI9mdaJtU3sIwJocX
PP8XxoGDfk0AZZBhI/uNLp2XHSIE/SdMuZmRa0b2e+EZ1SMvQ+JtOf4gMttvTGIi
oBPUbNqetD9QxTWhLF3MybQg+DWsNHpnEWdfplEDQ8XVqcQq3dey79Dfjy5GfLHG
sP4SOwosfKSU5N6DFkWwWOpUIGbqa58Ilz5Vot1iYwxIA7REML9gngK1EjwdRcnx
04Js8wh1lm5T4D1/+Y5tnY8Qh81W6Xm7D2gi/tIX41S2vLxplaVhmhIVZDVKRKr6
2Vcu2w7+3ki8bgSNsbO4tzHuk0u2PyV7zZpw7ngHGYGgWevFsw6NpqBMZQNnwTHg
vHDgGlIVRiiJLNL0SWUp5UMMpju2Pu0mTZrPz8iOL8zTH4egRjP4gXSqklHnZ7hV
AObZ+7/0q6E3+gEdC/w88PFXiVgbhtGKkrdQAJRLxN/rw15IBqAZWVAb1hF7H4j5
RKczjB+aKjO9Paldc+vtPhItKs9Eg0OkRsby1rSULIygZ3g6GnnRnMBTaLb+hH7y
TgnkjLtJptIGL5hfIR+PKixjvU/VgLs5JNIvqrS+nepwEiiPToiMy3wOFoyQgLF7
tNT/3UKZTQi02vV4Eo2NCc6GLFcRTcztUe4NyEOgG+9bk3Z0FKvDaFJniidkZ8ac
harz20n47ossPT9DwsWUFgUNn35Z/VwqaKRpXSmpzHYlkKTFdM685EPZY7J6uG+k
JDZOQsjgDZxp4utJGqPgu3BIqAl4pPzVR68D0cLGmI/25g+ImmCo36JHGFHPE2WM
1geHRV26AAgq0rJuGEAllLfWlWYUZaWzZKE/7R2Lj4Hx5TD182ufAGHPb3E/0MTA
vkdysEfJpyBSrAWAqPMqETdCseCJgXn1SjL/B5fNnsavab/nPHHCSvkQKfNiBphR
MpBkVe4MkIaS0pf0Dg/T2JvwG9ULISN7WvaeCZZIfuVUDRIBahTpcV0czLoWCckp
h318G9RUjqTlZ+LAXHuEpyJ4YE/SGzkkNjVVtPdd6PV419HFdwnzzYxoTf5iF0M/
4Tdh7pEE7sx9cE9ksBZv5YACLgqO/i/gAec6Mz1HAjLz3YQdCIoaVBorHt4Z4uxg
bm7xWztbhbY+9FVE6WericyREkWzEzw0EPUv67LhetaSznxi+Pr9DJk1CuwzERNG
N6zM64fxTApTPSrZcAV8mCqP7sBZdxAAjbm1VT/14i3unCqqJ4gwx+SNWogvzYZ0
Z7OUk784hov9ykF7sILi76OJg2pW0mUidITh2Yyn1hovF1DZZ9FWtE4G2ZiXmAg0
aLqjQjX9rdvSE0/yn2ztMCDmA3nkCUv7MAaqrnC/baeVF+cVc4GLUuF4u8MV/YhN
YEFuPowTYZMNqc7JaEP9g1kwbg/B6AHflHNgsDIEEq4IIBQnB4cjYSew+BaXihGw
ilEiDvq4uUnYkNZc04UNBL1AKNUpEr6yepyLneBLwNs1xYgNMB5weAfXsBkoRqoH
eLD9q2V5+NUux84KfHWU4imXjIDDfeDT0t6mpK31sbeWf12A2aQn/yvqfoeSFg2Y
1QRwjhbhf5vxxhU1Q0/ugRXANbg7WEW1QygCKPklDfpKFoQqphO8KMq+1eaYwAhx
5UBePO43K87HmbIWMsb6kOW00KzQ2hsfF2CoF7TQ3UEP/YMR6/Wy+0EOBRBRLe2x
OxoGIeAhoDuN05ZSNoj24tknBe+OAEUrgiiePMZ/7TJlYhHLqwf6myXWAtN2PqKb
AsaPFCJYaSVJQOa+4/zM5eNYSa3QRuqv2usBWlF6Gv04sA60OA/KsEMdNwpN3CUG
CH/Y8yiU8+dGaW/tNFEr6xN/ICfumvRcNzMejAlFQYjhc5E+znMReKOWSs/SV+MS
OW4eq1N0S8UH7d5suPIA9wg7kQKKbETTQPUMH2xNcCeB46NJeXWKtOnH1q/O7bDc
g+fFRgN5pVUMwJ2clvzK0xtLam5y8t4phQIp6Vq44FaWJjhqxAzd+5NRBzSlrS+9
foW+GLCy/t0M8Vh77LjDv3EF8i/PCgq1io4eXdSyjkH9dyQWU3S1A/GPHFsHJAov
RQkpofv/vNT+0EfeWi0OXgLxtf8OwC+c2G6oKEZizNmAsAOrTXQqkSdEK7F9gkDO
2bGFfon9dELUv50JECYeqzqSTCi6W+9V0Rgwlcd4c0Wf9QtuE9BFoiHeBkM3awET
WPklWC144lFcNcq4cnTs2KOxPbOXYKi1xGPfVPrKVWlw8p+2N0kZBwliseExd+k4
qCni2wfQLxJ0pvPKc+OChGMKJ4/yRbflFrvxZ6Si/700/2ifQuRvRvKim4qpsiZM
X4gB11Lus2oWREQx/KE2fM+95O1FIMytIQ3k0KeL8Qf1luctN2fEVZx0PYjxM64m
wIp5YBit7LuxLWW3b5V/s24adOWNpW7LWKJYGfIDQkyScFnQT42hlHE5FPE6u2Yk
hGS/Pd8vaLqrGkYNorHPe54P7P/Fjq2kcn5ezK3RU+AsGjkDYeZAXBWzSlyLHySs
+j7+1CWRc+w7t4hVtfkUo5B1r7e4734g40QgfFegHrwL7mYkNwrNwHCzpq29gjuG
GHAPxzqenOnbjsK2GH95cE+T0x35qtEO12we6bdDbsCQksil1W2YLxTfthE5jsPs
Hf6KzwVg24+06fVaI6pMEmUGblyuRK+SJTchY3IbEBwa94Gyci13dOY4gx9pBbqu
tFKbmBnJ/Jg0HKyqL/MNuWMiX0EWo0+SY97p5vlFHT/KmePwU8SrKl4qbwTfBHgc
pXXRF4FTjNXiuP5DpiSEu91XGNOBHOUMiDTWJcA+Uxu8XbfDNOPxEWAUGNg55Cjs
jlQdTTxsODzBDXXG0gMj+1O0+Y8Ce+PHVjQqi0kmmd4Vj9/Y5T094OmULFhckVEe
ViMwyLq9WiwLPWvhcEie/DR5PgeUbe1eFmRMSr7GV1q5IW7+f4mqUP44sc6WlKiq
Wbc+sxco5koicNyKHek8xauukoF8CA3HXuxdEQOo8miti6wZ2SDnRtWEuViIoRAJ
2YwjryB1fDRcuyJUea1wWO4nak3N/q/4YqSGDyvBYanlOeXSy3xqiInfNOS+uVhe
S++ZYYNBukesNautLrGZQ5CwHTrJO6Ljcn5/AJSnKBhKJt3NyAFVL5uoJw8Lc/92
DTGTqCY6fTk/oyHRypj0+IAiM61vLY5fHbRonOfFU7Zd7mqjS1B/NsZbzZTQPvbE
C63FRvaMYC5ljqw8zPD732JNW3gnFMm0ZAn2iGbDtVJrG188DXM39cEvy0TSa6sd
JG9bizp3U7xMuy2fWI+xDR6o5dFZ9BtiW6fgNHJQAiEMBwdYl4ijg4h4r+FoAtQd
gLH+/2/sNHx56Q0Dy4w1o3UJuOv5zMJuztajmeg5/STi7nBBiF60IjWdrVbOjQMr
AY5tw2m2BdCpMHH7OoU62ISYiqvHa1Y4oDlnm8DO+N20Lm060pL3jK3fQ60AC5R6
0iRX35lX1mbd2JhBIHbcjDdFvypihfWpZvgkXnmv9nVo7fI7HZ2TF5Pmnt+pD1qs
J3+0vHT7CdDPqYqRV34/ibJWbHFitQJYtDO8u4u+zLo9squtBJkNypM0KTQZw53W
Mbi2mTuoZ+JO2JydQXdK0GCchcnF8bjhhmjwbxRyMu8hbJk3x9kluEB7ClrkVhCK
UYMOQ65x8hOqP7wcuJudL8/JSRY3s9P/Ad2S9ujeKAoZMZmqN+X90SXYh43qi1J+
zy5zTBGhXFp57H8LIn3Vy97XuFq6bhoIakWPA/D1lB6s1NAU6Xi5XRqTeajWUbWU
4z8ZeTz/Lr2KyLTuVqXMRGo1pXOITbcZ0u6SDK66o2zyfZwVYkzWMEXawOvZNXxp
tye5ENy/29zgBdVFx2XfJLNw1ZJO0O82oNT4YjeCMjfFJ9zbi+DYXvr58mTlGNp1
0j6mKJgBL921XfGFrw3fk0B0IkC7XGGqAO91/iQbqHFNbvZVDA1G9skKnGOc7PaP
qhfirWmIQMgje6qkmQLCwuRf6CKyqGS1kw/bB3OVxu3vDhgQGZXH4K/kyOU2E+th
fcqPffQAz00gwlnZ/RPFGUXwr4pXBj9mKaqlFgHEHY3pz3TjKi1xnpDUqMOtXKOO
v7kvTMV0jSwCw2KM1s7JiVKU1Y6oFj6Jxes3eT7OAL7msODovZE6RV7N75umjfvl
QOpaNOK1PnjBZxYIXQDyrg9GnELf9WfziR+oajYJFCQ/6N/bA9Z57ObTCWFggd3R
VTQG5g44wsrfJlcIOQmQZ9QMWo+gx41e+DTeio2sikWBeCyRNbO52z2WnX+3iEmY
GbuANeBnTA71B96XJ7U/pvJiQszBGkDObG+yBam3QTIDRmBkhjFjiSDO9GzEIaNb
nhNYOhP0uE2T/NklJhuDm0d1fu49S8R2fWC5yhoIB2XTsQhdnqlKcYbd/G5Ej/Ns
yFz2ZmVZB226o8tLdbOOHXQSuOSqkYqfkACSsOIlUrfAYOn2AuBq3DfqCx4vDLU5
AdMdkj9alGU8lF/0qlOKjdqUgqeeFQjzsiQAa2sKsO7Nnexe1P+PmyoZbeMnWzl7
WJ7SFFHUNONSZjSgiB1lDpGMoKnPbacCZHisVWY3rzf8YYhV1eU7Yzye5e8ItyQo
nooW/1FTrDvDKeh4lOZ47ObBFWp56Qz6pKc9VfHiEOeuda8fqUwWr1orTIdtmJpj
FfH192cf6RM2WcLmxOE4N7SlR7wObKVQCOzGC9E5l5KYYjVYuhifhnqqwjzdbfZ/
390V51Hxm/SKoNKSWSdyhOWKRJGXvY5OVogB/pA+TbHjGoDLwsTJYvNQcQWbEqI1
BHQPSIQOEiDKN1QJhfMq7dKw+OR3lI8/vpElqHG1pnKEdi4og8AlS2PtP1wAftdk
lh9RIXftgMTc7vsFFyvT8h+lVVWXcUX/t60cfPZ68TPPmajJJEzhvbjKAU+VVr8P
hvL89LEGJbohvL+tvhYAREZpfBlp8DhtKz0bjrqIjVAnbXuBaOq92oafAdhdZdbX
nIDvUgQZQElkjGKIqhR+MpicRT8O8WzhFbGkbLgJZqa3q7cSDkwLJkEUx4eD863w
WLvcula/lKTE8z3GGd2gjIiEZSozYx8OkKXdf0uu9KxAdYu1oBrT7RMpImi0rK/W
+DRLOgBdCmqwbDyWVAGQpZ/TO/CrlBoh9thi07midfNk/KXyhHrA1TjcN8Ejka8g
RmYCchjigaZQlM3ukPsA6DuPP+IpTtIebuP6bDAvPp4/H8ZCaQGjMUgT3aG5S5Sm
wJ7WLrE6/2jjqZTbKe6yIKpP83jRvTAf2qlxpvfxBjwSYVvHjAjXylpekqVT3tea
qyaWr2/Jfobmul7leI8DjD9jcmZV+gXd5d/+WC5g2EBLi6RPJuj8i4QTGSu+h8XX
yWG52V67zTkQ4OqmiHAxNX7wV4oEJ8pnk1aSmpevKmGcpQNxCHcaLW0IIOVm8zOb
Yso6tRivORBzm0ARRV1xTVy0Q9910KwhnPbcRoFIQpnUVX4J2agDLfBn3g9va0zw
qG3EUQaQcT+G6x8/Pantjmh6wqpAkQErFjfPFCeY8yN2U7rQz37BWObssUcYP1Ji
CnKwY/r0Ahdwtwuz2YF6e83V3XFy0XRVIpn/LOGfAbFSu+a4wR8KJnDLF6rD1872
e7Ka8ecE63D7/JQ1/4ecM6TPBM7/G7xNOTC2KChWLfCKffdB4lauDu5aGHH6GtAf
zlBkWUF5uZjviv9KETMC3wxf3hlr+RzACSIjPPIZpnGvlaJPTu4kc7KoYIcgEs2i
B6xPeHNXD3xtin1CwgaajDaWjcIMTsrquMWg/vhsEzQxQ92OGma+A2OOd4jyS7KS
BV3cUgUbqIIhVNW/acqjlO7VybIu42Oxj8/Vzz+i1WC6vs2WTMIfBxKya0I+hIGl
XU2CITGr852OpUctQQIhHbXdHxNwsVycqVJ0sK0vV5YU7g+rWkSWw2pnoGCtxleZ
TC8f/Cdt5bQ6tBR2HyFu7ap9GQN2EmH2F607pHut7OBrf7HbYHOJ+t4Ho/9pYe72
HcOOXd3KZNG01flKAnP75zmNLNE++C+SarfY4d4u6RMBdPDpSqqvEKBxVV+Ha33R
ZFVur+PU11M3TcULNIisx5sc4vNcVWIRheAqUHZP5eylFPadvif/wqDHg43ywjry
O+2VY+74tcD83MDLROqts6sorIMF6sMxuSQyOeQ9mSco3/vtkNy/OD8/7HfN5EdE
RA9Ux1nQtzyuAHp/8GfcFIYNSqzOZFELRkDjllwxUUL7+jBad5fI5Dfd1hj3NWcf
Q4zGImKbiXCog40OMO6Uv0u89Ptc2P5WNzFNRzj0jjrYdOB9oX7t6xLtkKKg9ARa
9EiJAzNiPF3DnFSQVYBZYlkpb/g0hrMhdLIYj85nJII3fH9+miWM7R5C+MkENnay
MGhPrfi0kVUY1oNrJPvltytcUlXBv6DvBpmrh1v37A9qYeutmhcV3MhyZUbDmQs8
sEXxQB+efv+/YdQTiuFKePXYepNVzYWLUZGCIETBWXtT2U2vLEihnl+ZN0ZRGcBs
li6c0lYGfJP8gO5i8/Bdc5HFPEP+eXgIlLy8AOdzxx+HcRnwnktgIc/C/0zLPu+c
BGmYwb8eMy+HnuopYljjquYvcCNvpRCKd36juw0CCqwUYhlb9amI+dqldIgRdOiK
gS3uvN3n9yqvrzXBDmCjCNtF61AdEbtjlBdzzEITVjhYNlAvIv8u94DN8owMn8Ng
8DN+YSXsW9XrtBsPXemH7ZIoBljwT+WTYGOekKrN9vaccCzRhJMdn0Faq/8oQFTp
acQ10NewjPEn1iXsKJLjyHqlCVALXo9XVE1GoGkLVpjQA1kX5sLMyTvSM0QsOYa3
2sqJ7a0drtWZoIEtL+M6EOYoAtnBMXd4wWozIF15GtIjemmz5xyB2kDwOwHchwkj
y3wRUzgyzN4OG5IPhDUMTSQtTV6tNdEyzGR6nELk2cTv2RBJBNYTzRTjh12uMK2u
SkKXYIx0mV9nSMCXgZ1IDlujdmd13cC/qtrUI06sVbFh8kVfixS7Gk3L+Xh9KZm3
/xSyvMiQQx6jf1dYb+wuGsWnt4bwNqFrPgEZkB77eF7CiWNybtVf88z89kmGbpGG
XWcGM+iFpgxJQYjg+sMZ1jGOdgE5mQidKFq77J2wCZtRyO1es4weYvDCTxonBhDy
Cyv+PCrKDT2KJtj40Rz0PP4+hE9v1f/+hU1vF8uakniyvYaoPh3W+bTf9o0oBCMV
YnYhcY8p1bOboQ46nyO8TyK0aW+7KmUAZtB05Ds8wifB9pBJBub9V0/Mq8wUrKWI
kAR3xccxqtqcUZIXYH59Ywu6Gb7bBLT+OR2CD14RcGL0YazNIgvjp9VBSCIg3ip/
iw89V67UyeUwaIIzJ0B5hKFLlS59lyrKKsUlKcvLGqEfWuhTXzNfFcMShX4Nef21
N6jgB6+dzKEdrKvITF3lWHcjJrx43pA849xruRIPbfEio2LCR6pxc99RgnNhHMv5
e4zH83ezWi+ZsaBMy4uqMp7NNT9pXmRPwlmmkD11cJhGV8Cjxvu8sbRHkaEEbwbN
i6YOl+xq3O/5+6euMwxlVtu0uE/c5C6Y1AlSocOKpEDjYwEE+77HDjko16TcDXBI
FG938em8b1c20Qo7wWnWh4coaF8cbHibPBsJ806Uh9V8NEk/zCBf92277EtoyGup
uJtgyDf7Eyy6TJVLW96iV3q78IrlysVynOQEQsTJr2FcVG52Ttv10WHy1XhcBXPW
Jdpl8bwiktiQpv721CDAiZouCH1hGoGP8IWf6sdFQ1jrEn4+9W6CV0Dv1FT+ha4h
k7gARAFReR5AhuNSYY3WCI+fwTrSUY90r9bONVRLF07Ck4vPVFZ34PO0cIVW4UCk
aZIVw77xEhxC1Xn28xVSPaTStJcqXpSVTvPg/CVpnwX+37qC+/PHpnkJF18cwPnN
qsAzBNgDunu/94w/zTGl4qztCaQo74yD1vb2KMx93o8mcvHlqqOJsJY7VeucHGrI
eTihAogNQRUSKet2KmHtgG8nDYLuKxFDLdhzLCrn+hFBCzpnVphme84NgipeupRa
Uvr4EuLU8ygb1AQOj+GHYWKC2A4ymIq5NFGEF8J870iZqiv8gf5yk7wLNp8wfxGX
oLDjVd1qqOfvah9o6SipUyB6OeedipHjE2OvNh+rUee3XFO9B4orNfE3ixqlNh1x
CsZ6xct/efMFmrf6gr7boeB6mQf4FuaHasDAxrufOOI9Ow0/MJa1cGQ08zoFkI9r
vwl+jwf6DJyjYV0ICUL+582g2r79P1Evi4roX8pdRiSkCo455PX5KwKdMgYcpva/
CE4fCzg1ebHK7/JlIH546gJEX7rslNbKfLtsWkL3tvUlWlnQVK7/x1u1c0PUQ8nW
dWy1bMrXCLnr8A70tgATnecnamdJh8taE7B0V8XmGBllbsA+vY8j+sintZuPd9+P
e5kx3K9XWUtSeSN01MMIzm3ifseCrx6lDY0Ys6KXsEqkz2LhW0H1ghDz1YP/P3gb
bhlTaQmKzOgKGILKUwpDyJykmrFma29oat96YbOVv8/wewWH+V5hzAisR9CT7uAb
Oa45rGEdySHW6BsjnEzDbIC5+wZ+DOk4hd8ksIJ2no92RzlZWDgPIwQYzANbf/w3
hEzOL4c9lnfe9DQPlxQ8IFqAehoLTF0/yhyuHHvZI1HS7/Tg+bTbBtKL7ldzG+x3
l8D96K6GalRtCaH12DeV2aW+wt+CJdzBWCk9aefpTsYMTGTV5235RtTHVe7o8Jlo
Ia4XCDzNXmemcae0AfYlf4eEAwpRnfg/1LPrfAAWoTM9/Qv0JYQSKG4bIG+PBQBR
sP0LBQtiwWqLETYGe/xoZiU4InDD76IFf7pBOhMdahzj/ul8cWX0Bc7/rRiG3P1E
XNtcqGvXHXiw+UkMNMcc/vHtJFfzw8IMjiCKBmoOMYZgA3U1z+HdRdTdU+Kepe/C
ce/omEApacF0szhPOwA5x5WolyCX8cy5sfXRoDr/r/TCtMZ8cob6EZVhKQWgW2CW
fNye4mnJTM7u9ZK3TGNyfxYjUbVbWVsxRnyLv1Rgl0zwaKYWUEkqP+acFn2Mvo3k
m4qBYSqOHPhpLNnxd1orEV3eGbkyLpOT8J/g41paNKx6izRor7JiMn6dx0ZnM+At
GW8AFGf4izH0tz1Ydvur3A74X0G1oz/LpjlElv4sBbgiUFvGB3C/fPRvjxke6u+B
ZSG+CzvK5BwEHnxnxuJmw1G1V9D6EDpUGoN/X9kZsp9En4aTr1SX/UKynDGII9LD
KpdScESsS3puYMF5S1Nw8tQlTEgeOGrx/PWJGmvegJ51GvxyTeFq2qb23+pbZLAI
d4sBqYdWxsXrss2+1mpG3pXUwJxmeft0oWgl/w2u6EZ2PDKtQs9CSAomObiY5ieY
c6wANFFOweG1uTg4kFm5z7MTFNh2SAGEXuONrkUPf4DsvuIGjyk03Q8jxYcQjWMa
xG9ejoyHMGeadWGqwm2SRHmGVHMBNqYHwAQpbrOrKqBNjGR3jXRJhsYFw7dEWJDZ
ncekcg9m5XqHopKJqILmbMOFkDFfZ8j1CK0wRKAWPzAqhJf2Ss6mCHP1x6LTuHNF
r198moDCVLn1MkamSvyIc10wscRzKAiHRHDnVHgFG6NKkuVzduF4SiFxonJAvcdS
uDIYYAK1hXgi1NoLJbks/wvYszyzo/fkyI1S3Ryk+9Lhxl8AiBcvJ3uo81AA4AiG
4fa/G+hJmKVXbid0tvrEyko7iMvyZ5pj8ySObekZcXc4H2gT0J6CxoADKXArSwsc
rN8KY8f7of2RpqWnPebf+9/bk3Efqk6MvQZYSkRD0HFYBoj+UjWxBgau3Cw7PG8u
PW/5Tom6BUjcyYnZEEiCCh89x1pfdoNIMMIzIYr1cjoXCTNFstbObneBIReJVCh+
Xh5rqTLIu8INJ0MQ9xC6D3zjgpndTuFE9j2l2LYeeqjiTiaHpdysiS6aAR3MFqkh
FN9jLp3pWSN2gxZCoPULCGXl+RNpC05w3+Z2g5L3HNmcNo6nk9uPEH8jmyYNbGUo
nfp3mYknVVwSQw6uVQvDuicXy/qCNjMJdZJWAzzWxaG/uaKZ3EFTmV46mQOmmOK0
et/HtmlgkvukwMl9dBQ3FHsFytNYrmAZ5GZJFxLdimV8YG6VQWTTYX551CHejVmi
oBGm0UYn4A5yVgJ3uM9jiF4nwfGpVoeAL+UobuYGUrQpurh8L1sTNCtChdeK6/I0
NkT+1PRSlKU/kCmNQCOjWOYGswjO/eWEuu+igF3/qjgCr80b+sHTFJBOJ1tRFnWV
CXdkkAK0twppDQudWJ0vOl08j97g0SXILXb5VkSKVL33Il7twOp/QZ+bwT3BDS0S
VCts706mMarQ1H8pkLi049eDn1HplCa+mRFZS8XrX5pFD4FC8uT/nxAjigoifLFB
llsQAeDc918iH6UMPbeOMw+4w2hShH0QZkmrqLUx+lJHO+U3a23DxoJC3iNLBWLt
RzTx64psd9ViLCZT/NfYY4iiDVV/GkNG9HLplNP8GbIlH4i/aqQm4rDLStGQlRck
0SYcMfgw3woCV8fX3LfV4tHM5H0gc+iEqg1Rt4IAc9Km0l5YS9gf3Bzjw5MgPHNk
31nIys0o2VUE9+RfR7QmApjoD32mXG39kAzSInKTNSPhFOJuzgDgc8opmRkateD2
Oe4UIo4QkVCggSuc/rMsFRe6EDIF1wcEPtFujeE169PoQy8ed+XP77dC42u3fWF9
lfFIlAd95rA7lxaqyWF00SzyiY7D8i5dWofY27dMFwnfEhawNCZz9F5GcMrNmFYL
flXpxbRCIDADIcXZdKHKvMxV4X26iwWkTOEYPkP1J6OH5sbf4fiag2w/tFjYBpzE
Ceo6DaiZXY9IXEK9QA3PIraUAhAujvfwPnLFDSW1gMrJk6uqbWb+OIj1lhyPKl9z
x/VZJKkkmGPoQT+73pgwSlFUBv9xUJW31h8ouPGfq/uJ4sxLvSzeSRMO6fZM6Exu
dMfgOlgawytUSE2XOfzEqbgJsNzFtoz5vqZIJkduzcAGN2nlTT1H8desx9ZeJPF9
6m1XH9R94CGgbfeyC99HCPdUBZArkDU3ameRvIi6eZXfJ8xAWiX081OPxLDvHUt0
ZnPs5gAfhaXVykrGxkf2NJtR4fSS/krDe05DPjtGd6hwO6GhQXsgzyKckifHCfwr
3qq6Ah1jo0iPUPxISuyX/1SDaGBvRXm2o0SJG2rSTLqPoINq+2txVYLDT/Dymouv
eHFhqGDcOzbR83ZM1W7V0Nmo157TetyRaLnWU4MjcdsYEHECAf5oup3V4FJhhGIP
eVClC9vS575rqgDJF+OFLTyNVvvI13jw4wsD6j3hVK8YcpIr1q5PnKuV0O+kpTgW
rpxHbaklzr3/CBP01BXt8zZEYh4Xo7WBn6CyZn5NT1q3vNCzOF5qMv/Psm1+S5Ob
PmuQadCl6rVX0tmrN4MsoNxpksIOUSt5YATrC8+ICQGkMZMYudnbnIFYVzposYvn
n4lqqRgeIUZtgExb3TOJX9xmTzefNqUTt8HuwnXOWH4sOoZ/dTFRAD89nm0UmarW
+mq9m6ppleKZuovBUbh+wzMqlLrJv6k5+Uk+SY0pmsZc5xC4P7dI+BnaYOFiW3ML
K9vblspycn58NafNRNeaaKrbe53PoYoFJiOJZH4UQsyxRrB4YVCE7FbqJAbHk8Ve
jI9yvEMwD30RQ1N5PuEXQEeE2rhovgNE+brGhS4wBS79vYBiob2fsag20k2mikCv
w6feQI2jN1XSbQH4W7U6hKXRFG/oFGbrad9rWIdDmmZFoRuJZfCH41rca8bnwHOi
hyA36E/SfnAdcl977r8/JsAKTCX/RYvKMvpumPARscKTI8LL2Ac9RvJgbxl4yHoI
JRbup5kz2QnSPm9r1/cRVtgzgU7hdv14ADIVgfKKDQJprN4HQuKTrQdkTRi+J3bu
1LaGxdjhLRRZezqQnfFCX8g9apqRPdxGNq0S657Ne9/T1zNZB7v1NRmCTqhjJ6KR
mU1fZQ9WuCzgew05/cn54HS/s1SKL4XZ6eP/xJAWBsoZ5hsjCC7nF+ftmgFi9im1
WUo51zFl2FKh7OacPIvxaYoCgI61NxLukp5v/+j+QUHEefqkbVLAZisLuq/7/YG2
UtE7lWuTdQkRCCz+l0YZ0B+85TNjKizVMB0N63YU+H0rF6i8/q/2EKNewbS+5f22
7VqTBdBk9C4ACwGfp2lKkesWxfzrXNHfoxK34hu/t+Dkfll/LB83lSwkXAIqnXcn
KG762ntImO9kxZvkpKP/FxlWhlwKkkarvOLo123zzEPW2KtM8KAHMbB/vIbaEXnY
0rqBY7w+DFmSXi+AEjJ2REnKfsJ4eNwCOiW9oYnzyTRxch0vjBwQ3+TRU3DEyBwp
H+OuRhpI/NhGLgkR++4SzW4rf+kqgrEGvNpQfbIPi/VkRsH+4duVggzcZFZDZvap
5iY5vnd1DAcKp2NfoKg3ZPfrlsMm5z6GdZh1IOhzMULNUdvHfxnMrwZOczeCAlgZ
NFtpcXxq+KEtYxuXYv15c6XQhtiO8tuM7mGeG/y0wIq4dVemuw8fI3CjqTM4gUXT
aX3FdBO1BCjMICAmGXYYbi3qZTuVvL8JfaYV+fRCw2ImXpXd4O06E2VAS4bWi7Ll
0i9a+8NZnQFUdcIwHi/eTrl4AmqxJ5RInjBEsnapt/AxRyaQ2JEcXDoThinrJCPD
dlex7dgo1G0CTCe6iCs8C0ihde0NGzAX+Kt6x5t5280hVcjA+35RZe3Ep9gOG9AQ
jvGt2zaXybmusANI93TLXXIL/YEjX63WfO1S6+zzqd8WQGERLEc4Z4XIubSN5Pil
14gw4OHagC31HzU2qGKPa/XElCCLUILnmtWBgD6hzjbG0YIlPI6AA7US4fCqd+un
IfDEXfhZKM3XfWKYHc+ZsYqlRy6rxrBv41LCM/9xnvGMs/B/dOJnIzs2I2zY0C2G
pA9O6rVMmIKjvOSNtTnU2XHYfMqaunkFDogXxhj9pkm93O1kFtuJ/8i+5eVSDgoK
4ibuqVhKZpTT7DsJIgY8NTEXxZdpVY6r69Tzi8m5QgEmXOIJzJx7NwueOQpjsgiA
lXDsSAVP5FAHr4UZQqLS1N49yw7jLEyS5yx+9ocRQ4jJHWxpIMdxeNhF5IsZBCgO
QsRD5v+inHUQgXvGhqiUIe1sAaO0VrV1uJNl9+pr0QaOgu3gQTpHyUoO2bI4RNgI
IHhwJazO3bNuoTD3F3c5nIja63BtAtKj62NDLfa1qrGv0CsOIJejpbodWTbboRXV
kSwDe9zRe6pl2cU4Tm/C/3LJ+0pmBD6mvMMPIZyMd7e1aLDFGUXHox54TN6RzGT1
6nAcRGb1ZgJumO1wGsAPw0rjg2TEUbghMlCJVN0lop3O2MbbbGYikewfTcApwvWX
CIRm2+iGudSpZ+GibAlx/o7gtZTgJtnuAvnYTndWhfPFL3FVda9+/NcDSOuqE3X6
eHtVyZYR3s2Hjt2vtb5P33FWPR5UpoWbK5iFrlFrfghUdI6X6Z/784gXySutPwUX
elZhfTfl12ZBdWDSCYEIPmQLzXnCIWREZiyDK0xN/DmAk7SpodrCwYn0IoyPLfJg
xEyo6tmUF1qFTnCHoqJX17lFibUHgIPg7w0YFzNt6tlwj6l4mq7lWrtZqw7e2g4o
Pm+pwplsujUNXI8bnvQwzcqASTSS4PGnn2Y4/BhCtW0c5YvFXLDL6JK+E00giI4E
EPt5WzWBcFQ8M8esil73dF2aaFE9c9+IW++OPt7uVbrXZFLMPpR8UEOdV0Ibo398
1UoP1LXNv2EvfctMS2+JF4+Pl8Q+c3EFD7waNImTMLN3bZROXCLYxef4vTjWlwDV
zW/LxNaXM4J+zUmDuBOUlS8D1YFPZ2TW8Cl5JpGkpzS2MagEPBrOMYRolbLJGsfP
G5qQ3h00kDoaFSsVzMQvfJpgoZSi4de4aeT08mTcOX2BlluXRhG1C/Ggz2bQFTyh
f39yx9/2z7l11hgMLb2sMyrsdXnHB2IAmdVUmrWtR0HnTzK6poWpXU1KeQMJXC/v
V5eqe6UYMe9jiWTVbyXNMICshlWDBCUWcUJygROKOy5Ah55w801a6jRpv2BdA8G/
ogI6UwDtaJBkwG78XhcmAIFruikN0jKIVKCu6bMzeZBEfaItE7/raXI/xGjoxAQ1
GeCfDXYlWxGBBasr78AaU2ynMq5y1gwNeLMBSq4+XLmIbkfCm//gCoh99N9TAEGn
E5bwHhx7n5mbyFvrnKX/WUHIrO0dqDfJ+1b0mcadrkDPrkETKXrM8C/YpRvKOKSP
pxZTYe5F3JRxPd7sAki7nMuZ9TObi+WGuvuTmrwiIHsPZokzS7y/0EEOZp0WOcn2
saA6ke84UDyxbqbA4Nz6xlLhp+xPSQ0OI+chOnmMehs44noGARBqR+VpbtCJBtv0
ZLJCGFWBd9nG50iBozH3f2w3QZx760wJCLSSUaQIDnbl8I3Qra+aW4NLKWD4uAkK
01nUCeEqr+xk3gFjhxRtAq/JDYurmQyK7HHnJgkRWKeaBTVKDwtI7zXQgejjO9bc
ik/rHwjOlAo5Jz0bPUWyXlu2NMRYRCOLZnxDsAzhrpdB/cjkJGt7RiSqr4aRGBTv
fh3lr43j/7S/STTxfVB4pSlZRPDxQX39roiedcGtDBmV01RAyXZZSj20w/+u8fg/
mpfth3CvwbJfgFPz5ta7IxhhT+eX8eUkzZUfJmVZtUGKzpD9hHw3s/imwWK9xOfc
jDo+dBMsh51xsuPn0OG6iobWs5RAe6xc5/BwN7xXSVElHXh3QTJC51sqxJaX76Oj
QQp4ysy2X6VOeyEP3Q2//5VINC1iXonBowz0xHIOnA0hRANqUPpzTKZ6m6fyDVmh
U6CxQ/JaqyPVv4+MlZlNHPqmpQU/AsIyxtrCH4mmo9lMyZACqvn60aqAa3bwldNo
eD0VPmTX1uWPTYxT8eDVwAh4+AGmVdk0N+JcbhD0U9h0aycROSrEfdqC+FkXVtUt
J/9ZxpsrQlWY1ecHpjEjD6Wcc6ofjyAOMqyi06/9P3LVDPEUGnZctBdv/wGhKDYj
eGrgmvgJKJZRyNPn/MFMWzkBd4ZK+bC5FYi4ReNytSSdjEN5r0UuzKq8hOGefiBw
VnysOHqNKDG42tIZsSpZWFGu4PUOTeX6jsZx+i+fGpDofOExNmQnsKMBqthfEK9w
1Z4XTXca6OZ43U1fRW4s+PULxu4bgpdlstWB6f/WQ8Cs2ptsMGnr2kt3fGO6xoG7
riawjCrozkoJJlz5RFn1FSVqTffP7Wh/0AODJNBlMYA1BAmoUuLp84G5OURO2T1d
LOkN6CA26e7w6dN79erhwELEJ135/U8p+CeoOA4o9JDNKUlgtTMWgOtDSQhFiKPa
Mb9b6T3cMa0uCQeuoPbzv8R+hGUyZcFGBzA5m9sL8Sm3QhT1yH6OGTRNE6g3Q+EF
5MZHjcouglK7dIaeySJsuDMCuYEttqAuQTrDQo30+RFb8nfwKxSkJpURYxL53DxC
y7pllQTG30Fl6K6iSNPHOkSFu1ddr+NA/5xmsBx1fSx2yxh81PZ7+LHPtoF4LYK0
eyb2d4g4KUCkJkKIw0nOL2VkVM+nxHftHrp692pscGIgd26TTOkat60mMW9OMX0l
7gYmRLYXD27lWdIS2OqnWJnzkbA0+By6Jj8cZ9OQYK4qfSQAtlNatFxf/Gy8wn95
RT0OrilssWIuWazIkDNLHSfhmXYEPodzp87ZSz+iVo9lLvHXTsOK9yQ/fq4forLR
4Ht8z0mAINj38nHgB5gS/UeH1tslkjDzxAXnbaqZaWWz28K8uU/nbUFiUj1gyF07
dB/dIqL/FY+R2wud99TamByIRuYKB57ykkXfvJ8/bpV1NBAvthrMa3daBOOCsh5H
eIXzC9vS8sYzTKYak7fLJHDenG4syJfMbfpxWx6Eosj+SNaaqhNtn4fK9VV6176o
MZHzTnRA5DG66ozxXPfgiVCEuK3wuiGfAiIeRMeoYEFL65Basfiswhpu3ianaRdb
Jk0af3nxVkLWBHy/g8UlQbXYWeW55tmnvCE5ls6/p6pMbD5tT7BKAC3DIaWJeUCx
Si4KH6BLt3/pbpghZfzAcPNm3TbQBV5j3e1EDwmZla+n1rLXdlrocXY7ubcrSNWQ
ZUYtMgqiXu06knLgEDz34o+f+lflzDRDYNhfPbs0XA5USmisB07HOHJsDdjgyZgd
3e51utbtNoMVUaF17zmp0mSfOx2SyyjaHQhEN8HvEG15584pWNHI+9s0PMtboLV8
KNdyYihcRdO6wZPDSdgNGKZ1y3kvPd5ayFpvS2mx7xWoHs4uDlvYA53cBlNQtTv+
1rJi+2kLTHTsYz7Yt06xT3ktRfr7XyuZcs9ngH5aqaYRITp4olIULW0Ls9ITehEI
s20Fyi1sJOK6voS/VXgge/wqKAtKIuw867fCvnBx8KTV3i/IvrpAnRsC8c//mE2+
+w6mrGOmIIIR+bESjeV/QUCqS7Gm8UrvvWjXXTssGtMCZOlPjfxvNO0gC8TjFIXc
b3pSl8Xk98NF0E1sHs8oGaMfaKS3aUjHcuzFXtcJHDjwRPBfzlY708FI0rA6XwNE
HpYsZ0qt8YcJYRX6Whm9kn50X+MN4ZGq13eyXH0ES5f7jHTZIBr8fn3K4SdvqYTH
1VapxURNismJ9g1+FijhLjSnT2nGYJNREy9TI1o9q0MruxuVmyA7x9YylqGJxXei
s15nj3rbfrdOZN79N0K2aJG7pUw5qkpY7LF6MXIy1crALHc1+pzk6l7/vXIS4vAo
zwOg8+nimwo5znKLkkgdxD2xF4fwq0aoXbZAoi4z4uHNbLLvGYi/9JxMrTqsTGMs
HDM8NReag0orKzqmaUmcXeyn/vYj+ra+x5cl+/YFXukwYNhZxfINV1jVxNMmljfw
Ts0RLzFCXhj1UImNUxzMSQGKBwn8lxTH2zvcsfhjt8Oxu5vPuMk65j6V8ZELJHqm
qIe9EN1v+iBVHbch6yKfUMPqCSJad8NUZ6sZEMrF0k237JkeIMMK0pNaeIB6u8Zp
DxfkVPndibYQC3ZljUqxJw8XQSWWECqZBaQ7+cTwqEX/NwuPBYEwJ05D/vqG4LWy
km58pZ0vCH+uwu6U5FRbpLDrCGMhccShuVjf2Wvp5SUwjAq2wZSq15lJBs5M1pnM
o0ZtWWE+43pvRJbcwJDyrOa4c9WlDt1GLm6GUuzwqe61ApLEhi2cippfhO/LgEQ9
jTjmPoKpqyfU452igSIwJf5eCptKW75/CK5hnvObdAHDCvQZSW8ppdIWLJ6oYS9C
8jd56NuQtYr6XNyu2/lUuOLRkF9YWiEDZro96HWI+4LdzYsocMcUwC0m8Tz9IlGe
uhQt7UsconRhFS1OAHWpXwJRb1BZIRUCT5hFvZCXUhCm1C4fC+IkCQtAtQAgzyMC
USbxVafPD2AjZBDmb997Gq3T/vFyq0frD2JWE+AJKmCpooRjSn5aM3OuSbDKMmQV
fYHrqreb4HTQ0NQKd/5e69qQhlBQ8QxpVOceL2L6UKRr6LxSAukDi3ul3GJqWsy/
YDHvXy3XGzjXSPE+ukikSUHj5gmF1kXxPPeu8/+PyCjsvF4PmbvIOigEe6MPJhhS
5uguCqsVrcLWTvDyEAMlYsM4nZEMXJUVBHSIVWoqqBrPTkMkUt02RL/QWxLepqAb
Na2+sA9idVaH5HYMQSwSW57cViNBxqhR8TxFdK92RJB4oMthfBIhAmDY2f1W3tRR
ITGBpsIRFWfiSbFCQr07tTfvOxqYi4AuvQVUFI9zNKfupLjKb5/eLS3Ya8DUepi9
fNNs6Rv2M2QrGeCwXpd6URvUgI4A36tCOBywuF96yLphk2AfMb8FKcCB3CofPeu0
a6MEnjteb6Qq69ZM71KseJznyH5Mfno+TSkz8+l+0TAvQQMG7Tm3tHSMKfzo+kDl
eyY5GNGpFJ5xyT2M92xxweRA54SDP4lzEykbQlvXaq2a5sz4n6TmcKMCkJeMFv3j
XscHpKBuApl/z7IPd+2kNVQegsNN0V6Oh+vZoaBnf9pgrB1U1azBYS2O0jkngk1a
nSHz+f1UJsJaletDUZwEz4E2k+YRummWgAAsVlqCGwW702Mxtv9yrdtToKhTY+M0
b0gt8zJLrimnfgarsFh+CfrxbjikCWSyNcOn98KJq7gf/Kcp+Qjc08dM7oDY7ZpC
LZd6SvXVkgqPnI61DEvx+x+O083sROKiQ21xDH1ZruR0GshjMTqkVu5Ry5BSdLb1
6Jakrr/zmAZ9aiio6vo4x29wkAE9Nps6do8swIe7SX7HL8Z3ymOZUjNrKDKgFsG/
k777MhtXnzD+Czsf9XFD5AZCFrddcjIdxo0kCHRbQ5XvC5VAsLUyMnOWpXmHURtA
xdlTxto0/iMbzuw24p7E8f+HT9qJJGYWIvdi6InlXKQbcC0HPAQyEgRz7FTX6YnE
CC+xkaJHKFPh1p5Xe4FNLCRUoXtFlqxOg5uQtMoD6Mu3N2ekmIaWCGXxDWRl4sDZ
m+VTKwdBI1f78nSxiDk2BFUSOxIy/SfPyRfdrZ69S71wLVEOSbDZ75TIEQ/OsFjF
BQsmIPaO/E8hFdQ3AopJbDNRPDcYe1ABBL/Lc63nYOyFJ+AjVWyLAYXC1ezY29FV
KDgYRxiCSgCx/Nz30PYS9+bBm4U6yn8My9NyQVn2p+qEefVuppSx0kb/i0tc8noy
GJCxOdToEpFvppQ5eA9A993GhfPgDPVlbYRmwWya4fWjYdWPGPdcM8bC6sLx1e4k
fz0yFBFcPZsnm3gSscNzuVsIRo/PvNCAFlbpdASqysBwxaIWRduLKzeR+8jp3+GT
u26TIYUA2lIbXfMpk5mpIhBAwqIp4qFwN0DKiXoc7VPqh3OWEmagbUPuCgTE8YvK
xsfsehsUyLK3DfH4ae0n5Iwv+5cFhdTwWwVb0Ypr8EndQHEgrSBgMya/BFEIa/Fh
hcuaS5EREsbk7mnCWy8i+AAZ7EzhNP42G2DOphpzALAQxfxNj5YwlaLDpIry0JS0
xh8Kxyl6ovIgy0X609I6i1yxD9+wpY9PZqZ/Sa0UYzLkD8YcVICUQkIBiB419IJ2
BniQ8Qzra8KvLk4jgxE5xgLUkzRn2BftYHpHVWNUQqzhyVc37x/dCPqzpugPm5CQ
RbvrKePE7kNDGu7GGMTF2YQEes2/XW8KIqy5phf/XZKV9RYunjmIQV16T6rYhehL
hvyvBfWg5PLdSh4QORI4H4OdeFYfFfEjRZn+pUg3Z6FHndhGF0Q6PSu9hBulen5b
l5SjW9IP6TwBsbZkKWe/JLOBarZLaoVvZ50Rg+apAHDx3xwwbeOBP8erePObpYzM
nk+7Cq6ZSfTROBqnfGIKl4xAYj7X+URs0sfQWoZzbTV6/RtfHdsxSP5Nmyfk+HJU
blQSdwn4kusAVT0wr36aC4dvDe5ccjUG8DDntq4BykEvhIl2PSrfW0wE5Zgo3gN+
Muc0wHBqRcHCAogj6+kKplPE87fyZzBapAJT3H2PsiT6btq0+hvJzI50Rp3bFUgb
3sRTf7U17OoMfjteL5C1Se2P1QFvcTccCj5GFa2Adpv++hfnziMPOUTCOcJj8BcG
lZQttEQejvTHGvBwrLEVwchR7n+DqHgBn5gdbEIwHxtEKz8IUafnTFo3t2aArk3k
IWzQcLRV0WBNU3iC9DFzwLxjI+m5mn98ptSXlw4fX4TeZSgaKrdSuk+ucKsIpLXf
iY4yZPYWqsLdJzg3NMXKsSyZUhf/BtfhXlsWfFk6RE8F7x3iORZ1qubruKp9uXNx
68MmQvGC9mCug8EE3q8iWZXPdOhVTRCP7urkvcqOT10KKZGSbN2G2JCRbduv6Q5D
aaptjlF8Q9rZNeqr7WQycDNFLZmIDIfSQg2KOk3uCSE1+YsIowb5pwfNIekdJefu
UFXzM3jW3HkHjCBXbApYMSlFUv4gGWDnZc7XEKXvR3rRFeN0+hLaBeKBVqcfDiGK
JgQz4uzoOKSyPNDBD9G6/5b5ZUmJg7wvbP8Fy9mhgDrL65fXeCKORV0urTy46Ryq
HbS7BIqWSf6d5/LQMMO+mx74cMTIwGs/zQlOnaPX4k7u8rmd2FYoJ5nEODccqQGC
43F0PiAK4anmQvoEOg2HOfKAZK+obVJwjS/tUUW/e0TWB7CAvFXetA4X4ClBYs65
HXCQtJKtLt7+ZzXTmaO9RSaY94s53PDb3j8vcn5uo+jWEssRwmKEEjVTu3Qbrcv0
VdoZJtgORrvkbxRofiYYENaSI7prEmYE8IeRT//gN6hK3jWmSD9BI4d6CxN1YXIo
LD6Chcj2OuAft2Sv8of0Dn+KiElfCLb3FhtoKtl6ofumZhayGurydCB2NoP4ltrw
H7tqBm0CASIw2GvxEaLFBQMU5Y9xIFvkI98sr4RMCUjESvERx4CqnAmgY3LLFrkT
8lBsBmWG9PDXv+HASNvbRVWXBpZfJdwqAQY7bTyBA3AOBJo9/i74Q4j5pECvaI3R
zBIeWPi4xgEGfBRulmQFhM5C0hcoNsvmYBirOCHlmENshkYg6TDHbQxudwcvYCZg
8RyEfmq1M80bB8//ytnaFHsgmRFMTRDDGUWvtrwMtKodU8JX5GQb3VhPbm4Dx9Bc
aEqy1gwDnmVLi8YDsOF6livCRviqCciT8jAFschJ8nbUG0aIngRYv5+9HM5OlDgJ
XDRz18YgqED0UpzwdYP5XOGYCmFkYDh3KUyMQCGSHOhkgVbGfhGjpDtqmc9/7hzg
orGueYT5495x7Zi9KVnVGq0UUjK8rPDwfj7pTNtpCUKcvPDXa0qx0cw4Chj5G0Vh
S+VAYbBYEOlRaUHMXfwPx6Lg/VTNndrsee4XmUY2ANYovriTX+EU8xIJJRDL17G7
rhAGWsr3s+9syttmIfrsGmSS673DGgo2pW5LDQ3pNakF0kLD4zAERxB+k4AmmgxW
mHu2Kfmj9hskwnHhsgdqt22ixaanT38MII9IxUwh1DIAN1UsdZ1hpvt76zNZv/Yi
WKZLBkJslXpA2HBQwRmSWJ2p9n+vU7kr3njqxkJCH8gE7H2gNWgoZx+waKMwuhDw
BVLCvHMR8lRfriI6pghizZbzi6FeumWLEOi5cF5gWp8TgHvwJoZ53FMRUEkFLUjv
cEsOFTJeV63puKY8MdBcJRyVVSRK0mM3KQoeP0wkNZrFAQAsw5cYseSat94NNF8R
ydAJOcNJX/tmiJWU4zwL0Wr5T9agBcAbLyzoqtgxPOb5ObJp0ceO5r4oQS2pazvT
MLZLqRaMjw93Yft+cPKbhrTQvDFT30oMkv5Wqq29WAbTo7bgyo4Px+8j0+zFE/tZ
AD2TubByU+Adzr0eXy2vaqgMX2M0tDNXjKvn/CgIc4VLySLZ9LBDeAeelNhRg4iT
Oud5wBdaYEv5MOPU1oQehZan30tC4jbIxyk4s1WjHVFuq/7/CifXMvOSrrE31CRQ
pdbGnpxbac+ZJZgdhRTUsF71PHwyblHMGOCkfQ5H5pam9ZQaUfofRw8sTjFgHSKa
85WbwTKCrMs6HiWBFQ2y3XhLeGySyKp3mQ0Up7kOV9G+2N7Za+kEOuIXh71hC6x7
/2mgxM+zJMQDszNOO8G1XINcoPNK+fvbFW/M2taU2M7pHstdzPrUzMEotIME5dNB
TA7NO+dq6DkP8fxCm/dbpBR4jzq1gynqibaQqyxBQgFmy3Tr1iyBSYStDftS0Kj8
svHzsmwvc2F2AZksVKSennP8CQTz/FSl5tkRPpp1c8vKrLaL+Ac0jwlvxM6e6ypO
tQRWt/QOlwWkqLBV1rGWMew5A4LG5okYUsH1Wdu8K5Z2ulAiqAtGRJT3GCUx8b3d
Rn6EC5k5BiE9HegR+FlGQ7U2gz2bypVuZGsOfwnzLJg137bqPH3hEYUBk0uDCnVM
qwDXCRWXXnh/xu134JH1nDb7ZfTf6cLVxIIo2Y3jr2r8P/TxJaomDIlphsUtPf3/
OgtjrMorUgplZgmMZdVa64w7CcJmCg/Lg2w6PdoxvdcZeDm8DJAwe09ZGsoETpc2
AubceIxZAIlnwCzilXseF1u91GA5GS29MtCgqhKbB9dsmbMnC/JSrrZNjJ61vlmS
zW8pwtpPWmJBspmUnGcBSVV5jvrrkJvuV5BWRGYoh3QwMsLnGckyCbkL6zgFyRYR
saZ9xT37wncUBYpSPY1zyVGB8vtGgL+MQ+FiBK42cHYE3J8RlIYBrDT3fu3mYNEH
FuSRBv6d3VEVm6F2Vb0+NmSUTATLAv4q/C/9E3HuHGTQ0t2lDVQwFWmA1NYurYtc
S9ZIrRJEoUcUDTPepSAtGGAU0jOCh4OH3mCn6M2j/8T/YPFxwfWHTwnBmcSh65y6
ZxeJUsaZMZ0I96BClT0YZowh/7xpGBHUwjKq2v5cCdkuTun7Zy4AH1XeqjZcJk7h
oyRwgEYYrI/1hE35nxjDrpSJ1X5BiwbA/9lpLRUAl8wPxFnP1mF5laoMJ8z7q+72
7DAcujr440aGIvaWd+C+h9f3/Ac4OclwMQaK2caI4HOMO9k4QA+ecz1hhiJrFN5i
bCaLh29BV0P4FfA75n/nYKY8F678RYee8iEXQQMcO4NC9ey3ZzKBUNtZZmpzTUrk
HEnVFnxSGiHctZMWXiak6iyM9gJ8LGtq54+/WI8PLF3C3XODR2cF8FM7BhNuFH7h
Xj99Dh8GE+3lL29blFM8c6Uix3MSyteG6XSoOsH/TKfOnBnWtS/cveoKwmlB3OwU
/8gSKSIkaeVn1XoUV+nMsvXda8T4SFBVhhQ50s6MizZbdAVJy3ua9CFDF/M//+GK
rGhJKq08bdQ25TMnpoBrrzIysGy+rqqqSX1S6+HaptxRWrbdnhD55Wa/dKyDDJhj
uK48JpGKEaEr9GueYKgJLZXq+t83q3W3Hn0ZxcHHwTq5UTWQzsxAn6NCIl6JKUnp
xn+XpNiHUzxmRWl0mrjPlAEcNnU7uTQWDWklcaPRwHsm1rzhVuLkFUUSvQWUdGLn
KUulf8rlod7UMEbv6NBnsq/4RmMeAJK6lcE9Wkx2MGtMsMmslCBSMPs8dxfFspjE
i5/XwigvLmAjLS3YYwkWpkGVb8YA42XpUQQRIj9ko/QGNg75F/r30P2Rg6fA4q3j
057Q4/4uGoN/pQABwNqBiguNMJGOD/ySwbok8FvbcA0BJt+wh4YgO0POAk+KVU+D
llBYZm9RZNnizHfP4hLaBMoueKfCbTcczroQAMntJf0xtwdQ8PEKu0vPD8gS5yK1
bjAE7SUs0SnBAi5ZmUUC8KRKlPNeSBpuACOhgijuB2cmcFgLZU4Ng5S2iynXJSj9
97gEHnsZdVcnFZsZnGjY3+y+QU75pBGYznm+0z5JjKU=
`protect END_PROTECTED
