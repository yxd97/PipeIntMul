`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uSKYj7DpBYFaTzKxE+R/AkiC5vIBRtcXmCC8y7mGvwPZugaZdvZxJDOsc58oG0nN
Z4spmN9r7TWuQ4qtrQ/TWZPAIaUP/3fxEFMFV6vkv1lO5KB8nVDoBrICousyePka
p/DRJjKjl+6v4O9OZUsPHkj133x1AH58I4chh6jl8PjQNCihkMSL7eQBbjFock3H
TbAWmDrO0jYUf3ix3H37v2Et2+lApmlipJ3ixRTQpbvk97T6u4L+ov/UfZ5pdDjE
2ncBuAH08tVpa8u2wUdXFzOJDFwB7cR7a17e+MdNKDeNJdxeJeGKCp+b1zD1sQsU
`protect END_PROTECTED
