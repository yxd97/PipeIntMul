`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twxPxFu3+uEQtQbfUAGEAE7PGH683tX3kxEI403OJR+7fQoIbAIkFjjcioL4bqJF
9BWB8IDugWyCdxN61mGSFLlbzZCY0FNnZHhdC15XmZzzWjDc/aV+eiWb61fvx7Nd
neJSpcFtRS/4mfqfpxU3jPhc+9xj96vCuc83g2sjHBnLCiKAz6paiphhHOesqqUn
TcWaZB7ZmkgAudooIEcH7/Z01TiKHAlHMSwVzLIDqs0i5N613O6D2/+LwIwJKXDw
y07Yf6Mb50Y6RH3xRv1i7VIPQPn7+byGoRwYNGc5S1j6hBR0JQ3EN7jltumrRLdc
eDbACn1qcIN2uf3NRW4kuEp4G/bQGYFDcFy8JbCHVZj+0bp2AUlUK3UgXCNBIZ+e
`protect END_PROTECTED
