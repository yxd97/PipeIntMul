`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88fzTRu/RjsQ0xjsBWFOhy17dAkxKPtdXabChQKGPZ/pePt4gYLlPs/Fqq492UpA
0TdiYSWrUlI84SIEMcr99Wl3Yuh+hjV921fV0lEQTU51qYQOCs2FS2EkSY9PBT3t
wCT11uNJlpKS2npOFGnK1BUC4z6ECdtSse2ycYYxOy8kbprnNPdWQnvyjgxQJ852
5uB+2F4eUJLyCd8BZbUp0CyibTrXI/pvnUy5ya+VhkUM3cZ3fy6/1HQf0tZg6JQZ
bQp5NijqF6DqCu5ntYoRiFr/G1tJRzX+TpRFzA5tHd+tWoqEkOBwtXeN9Ld7lsZ7
YBsllgWF8SuptUB2iV9nFEqqfwEiEL3tc84FbXCeNrBqgIM8xrDZ5MweBdjys5eg
DvWv8+I9QzvtF5m4bonnaTpksneZ5qdrrgVEeVnMXyY=
`protect END_PROTECTED
