`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rES1xtNWG2GcEb3BhMNlRSdOxlVZMFZQejIW0cUWiLHbPpAI3ZDYXKRdgVBsl4zf
DaoGnmfoG0I1wVHNnSX8bjHdU9My3nXJRHfE1H8RWGQbVSs2TxZ2EYA8SrpsQo8Z
0H3TVbhHiozi+XgDZvuQfFyOEXYXyf/aHk6IyFEfRTFxzz08nRs3DDyoOdGFc4yJ
xSunbkiXHfmu+l1e4ULp6KRrcypM9xCUt/xVBzDVrR5dsF6bRH1vxkAurT+WuheC
RkRSsBQe0xYh7VUK2HkwFLJtMVJxOYr1aqStBsJGQqc7RR1Vh7+XTkhkdSA3jE8a
YFZzpICT4+mr3urotzLYErj+MPy6nXO+sWuVyK0kPUFxvdmfhwGOkO8Brw2WNaq6
4PgiM7vaO9t1o6nuWROhzs5mi1KrGMa37KHWhSarT+k2lDEO2LWkh5JQORL2aKT+
cm9U/ch1tms+OcJEFFMTeVujCpdEv/C0iXLzqNIR2YPYD9tjWeyvPQC/rLUSSuZ8
DR4q5CHnbui6WeXudC037TkqrElPj8d4FyvSSFqfK1SNOG/MuDGn8PQI0xKDjD81
0vcXxln2iwbi+0PEKFmj+mOPK0S91wga2ZysW6+VjbDuXLf2O8GLjvapzsvHFeU+
coZuyGhOSrcllctb+L69Zwfrk5HQhxrbx76Kipjddi+gJtH6Q2ALy+XzbRI+ctld
V1x1/zRF2njdujZ8JturDw==
`protect END_PROTECTED
