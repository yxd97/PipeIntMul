`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YZqWLEIIk7/FiQyJd3yVY/q+WYQGaNVG+kpusUjoISmE38HcbSDh2cW6PZN1NIQ2
CGNlnGr/2oVbdZEDfwW/J3xlvrdopeODY6+VUcgatdIfmWPbKEq4rf4h6eXmdoVy
SwGdNbYIVSU+H8SQt1UADxt6LAZykvAXPCCZeiYw7ZMLUfSe0tojQ3kBeWGuh1B1
/pNJQigpFXAzjQBN675w57ryNY5lU1N6DG8MJQtxAKQS6oYvhzIFqknVTVYnBc+t
kd6cyArH6d3JEZQQ/HfhSKf13nPAP/RQroyOR282i7uTDcW9umPlp8/PBGVkh+oK
2zc/gwBmK+IUmPgo2d+gE8AuK9YzswU0b/zblxjzvodRfY8kbOLMWKjQrSLsqeOB
fdJAPOJlAg6inkNRKnJpXY+1VhmMEixxFbNosOHGETBwXPeQgXiXcmg8TlCZygl/
vO3XvyHIV1mHGDLHcpH3Xk/2nuzFaPrMWRSR4mpY544=
`protect END_PROTECTED
