`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7kzuq+p9gOJEyoqNTVhVaoyGJemqo8ZnuBxos+9uUZngqWQHikyv9CMUNqqLB2fY
NGGNSg3jGvJqWeZNwOVcfe/1jc7aV3CJihvIxbPgWB6LVnyEoaLia6+mfnfXleBM
PpiZp6/DTkYlZ1Rt4MsEQMO+IT2qPdRdsS9b/DIRXlR6ATpy2r5MN2cQZbhT24rj
IqryyL+Q5lNBskIt46qi8zugsMqB9Ci9oiC+YvfKuc+TtLl4MDM6WbXnV6fZGwuM
Gn5Z6uiVLdT6E2XpoDxtyd/E0sa7jSa6jD8oaSYy85Ju2hMh2OCf1GUxPva5LX22
LG1XPbKAE5AwZZm5RILEJw==
`protect END_PROTECTED
