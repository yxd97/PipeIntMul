`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QKVzvsps+bQE1utUJviww4WtXJnssEEcQfbqNTx5CrpyfofCtjGHz04rW5gFR6y3
+N5Y1PPXc5LbWt1N0VGlfsPV9FRv3jxXhIPLZ3eugwXdzmA90qmQIdIQ7LVi0O+r
SG6nXyO4VRuayoBch0FWgPDkSrZ6566CpzxtcVkoGg/QyGPrqBaPB5IhXJs6049Q
ErbMKoq1WnYcYwpydQ95kKVFEgmnBenhEExsysSonv7ewrtI+dLsfeBBw7Y37RHV
fdJjIQvuUhMJwsqwQpc3uDijOhcvuO/xGs9MFUdnjsYbN41exDu2U/WdvP0PwrLz
dRgvKr9f32uqtE4HJE3BTzIXjDNwXfapnG7YbHo9iRtRWONRuzsB1zKnAnmS99h5
a4Grkw45etUhML3ZYhGSk4/n414fDT9+KGoSgnKTc9TgZa2SYR6fHhhwMlfergg5
4t1GwdTraOJIv0vJPCy6ATIRMK3+KoKld7Wx+C6Jy/ks6Bzr6gyQPj76t1f+Otzs
nVc/jo7UtTrKvIqb0sfB/hAirh7zvU6avljyLiTFXw5l0XutEpp81uJB5bsewLy4
g9ds1pVFcZzmX1JPNkNGN29B1QgaNGvNQr9gmVo/Jtj3j1DJr5c8LNTg+y4VT1QC
EWeKyqqXkYJviZ88TWauNDcaXrisnwytDQ82Rzqznbm4AB6rEp3uZG2fjYpcO9I/
ien5jIiJctJBUp1fWoJWh1XY1t1yAXAGdxG0QLIYKEC8jRT95ulGh+qAAV0aem7t
rSDviCkGuX/AcLzn4fet9sGuhwVy119HvIMchsqe84RMHPKYNs2GP49hH5RE+5F6
iktWHRdIbD9m2Gg5MjGkri4SMiMdrSwEQmM0Z8Qt+saaMCVkv5q2bnvuisf8btbv
P7GecaCvdpo3ZUSTDY069vZxwkpgzUUxsaEPUDoZCKiZdkYKALA3S6iAmUidmhUv
kSUO8BkTaED0xjBAeQnGt2BwgMc8nZoL3V53ucbpzF9cSC4DWBTF010m8eZcrb4s
RudRnwT645b/XOskVQ1b5YBv7uMF0CzfpNfWoXLixX7wnwyAXQl2aJ1lrMjGgSQJ
O0t6fyCjGAUb2YgFNwnHUrmxpK+5psAAhIfyQ9VP5PDGF7q72IJaAwzFBnJ9OoQV
LEOKPz006ZzK90p5a767++8jMmyYCapxRs2T5Jto1Lh8+E73iIBRYp80wE3RIbsE
TbMsAr3Ais+5QW72KGd7uoEFkQYCSfreZiIBt44q2fK5XCynPXNic5O371wiBjjG
cnwqtAcbTJDeEWm2IFzxQZV5BZcs56fINGEZJSNa6pbZoTu6pgtWLXpwxw6eX2GE
N1pkj3zPJuMU3FH+05NLBHtD7xEJvcwJybQpIf8pfbtAK2WAi7p/Lv8Msfl8QYTB
4wXt1m9AdRDolLHKE9zdCtGmGQvSRwe/3wfX3b2VwpjpeByInav6n8Xqi4iNb7AH
AbTx+Rspr3P083Ijz4RBCTvBZoKRz6tp7EkzCOLNMr1fef8yN1hMc4Lxd/+vat/A
0qfLtNjrGn4p3X6f0GVC1hf8xYxBJgORqw4KoRl2HO/HZuU/effpWPjt9NN4J/CE
2PTpWtth1ICl6RgpxX9MIamezfSqRrwFdF+m41AH04eB69OMV32RXfxaKIAQmJF9
hJ8RJL6kQgmZLfi5dTb3mTeS25HwL+7scT+yZhSuN2qFBKISkfjFG9rJuErR9SHL
yhlyeB1xJONUTm01gmBzIfzj5/ZmjsUnhyOj8sE8mRx4J91gwOfOjciO4opU+yEP
tY7eNw8RUhc0Ge+n6V3z8tGPF57PR9k8AHqC28v5MSLK1fTvastscSa4SXo19png
a6sxg568oKUwzFNVlBcKydhskPQG2W1jhtYNC+Y15OnW2dFtacCm25k3dBFmpxuH
PWi0sP/JXvhk0mhTOWLMdIl38KdT0XHZFc281gq09rG11vanu+q6qaSOeMX2KY+8
tcogqM0EQxWohcM2QMbgbpjS8VFa/vW9D0jvug7YQo4EMjcZnbrcGoX/0qqOyD26
MgpSuWMKuFuYmsPKc7NR6TAlOMCX5YppuWqGPBoGpzHcuVyWoupxhSxHqg1+Jxfp
kfNd0n7/OSF/CeEP0a3KBkT4G4SKOulnnXlYb0jfff5EO8Eg14okTsqRG60ZI8HH
ltnF/dpRSYU7n2eC8TtJr9f6h5pHtNefd6SX+iBO1X6xsRs2M2fUR0Yr8ldGy49V
kOPxhxQPeEMHN+HIWguq5j9Zhe4o2LCDNyEy63WPBrNVXSnxD1vXBPUz4gxoIKva
kT3LRXZzpcsGtaktcvs42Jmy0w9B3nTqDKKHRAPOUo5VDJ0sseJCze5cUlDAbI/u
PB0TE/5NKtS6BLj/eEr46pB+d80QsZhcKovY24AIhbjHlkxAaI8L5gIq4mMdAHtl
V6dLKalnLTJQ0tCGZKlHZ3ykdnv5vTmZTmJYR58P2C5j1kujeP1Zu+2OJSbt/2mT
o79/w4ey9iefa8ePzOPFq4osYMP+CA81NGzx+KCsPZyQNN4aC8hhXBna/4kM4+8D
zo0BD/cish0zO8rIOBxpWa121JJSxq8wewDqZoXJaZdctQD2MU5MFMm+91iUR0hW
5ouIxL4B38KAbp4nAn07gyFQJ5A32AyyreTUPRgsms52mH4OpY7FsI4XvwwQjE7J
P9LeHEyAOzU7le2E1SGVnjgIxfRov9dOVdRRwXp3kVBr6BeCdtEo5cck4/F7xWOr
RvKd4qOywBHVwU5pWJQW0c9L4WtylWJPk+FcZo48tZzBftQfyJw/WVvbTEL3puCR
RSKiZU/hXdIVs+mv5jhiVbA2g0hxUzpAF6tfzQdLFqA4JnUl6hiay47a3GO15AvE
0aaWe48Yu/uU3JUEqcMoGOdr9BXq3/eoBR0wfgbzuqNUGZH3LGrk9NXZpQe5n2/M
lhDpi2ljXP4/k4HWF5qhBHnjTeYY8e6u0ekxubzdoH+M1YiXfW7f/jujWGcV+vxf
faoGMiZhul9U7pRFDACNvnBV2ySGfAaxLqSBr010aLwxy3mVVaZMtT6eccbTPRSk
MehzL2GgJuOHMvExO8r9R9VzU15ddHXNP+Hfvd0XglF9l6NPRE2vgc+D1RTJyrtN
VnhoYKdvCYyK8pCoGdkXzflXD94LexPQK2Kg+Q29N3Tbp9+jGSFLBsc6GdK+GNls
eiKMQdxjbCLMQhgGibugkjxbEMbEu/lO/RB+C+rrn5nyvBL2Vj0h9+goCFaMIXd9
h6THXoyILZ7SlEIyEuzXZRl1OQ2UGfWqbUlUGl0c/DvWvawJaA542N4r67EZaW6e
Jr4iF7SQZH+0ywTgvGmnXFFr6lFM5TQsCToVXVVs7r9USIMMF6MZPeOtbduojdbC
q2feQIYSU9PG30zKJDzz0bf4FP9XZAJSPFr9cBRNzSG4K/B2ipcfEpb+0t6P38G/
Ewctvjfe6Z2SaKJJOME4cd5MutWewthXEd2IwKFrUtYJw3jKpiAnCbWR9iFNjimc
HPbFvw0Sh7osMRHdMDQUKIYzQslecDjyTOtJ3mIdXlnqvtRNXUsmc6sgn7lsRE/d
p0iCsN8GXoJS171QBjxUGOtVLwU/gdp7N40fs3x4yPPS5GuRR9tQ8vIA3CcfzbG0
qc/cn08WDnf8AzK8+P9zymP8I2YZunpRtEdJ8k4uoCsch6mXG9DoH3kYd4ilLgy/
9hfl6a+ecrgWIQd466Wo/YrRTEUCCw28STuNOtQF9aXXObooByIaEXdoy/yUl3p6
vR3mWifqZM4UTyy3EWjMBNGzJy+5s/HQMPxf+Opt0J58xmiRveZ4nwetEP8qGRnt
PKSpBz1Hsj+qqpbvdiuec38w/72PvKJ7shNajrQ0+UX3ktPiKItO+IOculnYwIYx
MLsof+wu6VyMU2AVWiCWDDvjfYk1/TcdcAflkTYFzvJFc2xtuutb+p1rJaC6EAXu
2wBfqegM7kS6qLYLSTfcOTEWQrj9xF276CN9dAVCygWfvcQvBezmJu6qEWUJm3Rf
VbSd28TMxQJ/Y/sienzvNBe+pcO20wNtWBDybLIw6m9XyAV94mOF8Jc9gPPFDJo/
rvsHZqYb7zkgyVwNUFGci02M51qcHVPPdC9e4MoNySO/2i/qWGQ61VqsLFi6GmvR
n9DbyaaXptf0pwa8KLLPN41tPgBQvfqQGDGFCTvOz7a3IES99WUslsmgfCyK+rO+
08JF+u6Bl7p4tIuSZKlXBxYgri+gJmCZ6hiukdbJU+zKZLDoGUkrfzoaOZl+3QqI
D4RNp4vI3pWlWYMFxLGiJ3qDCBhyrwoAAmH9lX6YS/LaltSFjrWHkLR75qCGZwJp
OyOulYjYa0Wlf3i/4SS25UA6gAHvOuFnrIAaI8TPynBt2t9Mc4oA9C0dWlXmGKV3
Kug5WT61QM9kTZoi1zia5ZIivstrfHESiTr+aHbvHwfU6xNIMcQSNenWwAWdWFNm
b1Pu3xRwHw9MvDkg3Eh11lYSK0lIueE7NTskSa2qBpyJCbc8Q/oXhaJVqXQGrC1p
+XYamAAgwrImMmhlsxWcJqQClBt+F31igf2Le6rURE/eE8o3OW3RLzVZTyWEumjg
kn6OG54h5TnMdt6Mw3ujmlnDh1yRxMRHZ7f4QSQOlxT663TbQ+gYmAixrVkQt2EG
qjEfzWW0nB3kQipNIDewg9OYxfqDgcBIE3LF7Qk/mutlF/lPplT5vVnXTuVEb7aO
ZGR/Fatu0oVmnYGUnrmJUgBEI4Jmfhd3z6JGkgJX4NYs9zMrVZq5kd8Lh3jf91Yr
n7ciJVcT538bfAz2a0P9lOytSyxOtKgxqxRp2pM0YongkPtDIc40Im/pAqOu6oaI
1TANXAuJ0htoi/MkbbzZvV5zMjHRzFecLjZIGtTM5gd+ZBhBIcbg9dFk+StTJ7aY
AFUUzCC7iqeCIN6R9TplP5e1UNlSBxfBptu0mjfwAu7aFgcEOvUiJ3QAlWf2Wzwu
e8Yu9WV99jtikdVtfWD+gJRDb6DgE7m3K5Y/Mc65ZpDktpC6ieMrOSfei8sWoe+9
yA1CoqJVnBmmgR2Z3LTK1Qy8dOn8S6UCQuG9BvDPCwKIaax2kXEkBzRX1X36cPdR
Rq8nC4GWOXDNA75ByBcq5wMHYxXfT8nYiKWDLgBCgpvm1KT9qNbpv+VA11qn+F2L
n6uTurIxmbFPj3hcBDpHN2l5HrjUN6+WIg6U03yJOkxJ+qtYlOmlmXm3IySmQB3q
HzZ/znYqpstxiv+VQhVsXeuDHUylp70GcvPVnCL6fc4Qb9noGIOEO/FMGXm1eyug
D1jvagyxrBqz19j7CP9nSV2V41v5iEGsrVMsHd8ITPqydvlxFJPodOPQCIepdwAr
mmNs25M5O7b7vxMEthB0BHbiRMKOl+s9+iiN+QpQ/5a10dwjPs5rgVwobmhfRWFW
+WHn9i2tsGwdE7QPVtjbmxdzsDR2UFYWdmyCcDsLtQizNgseIpI/KFMObTELKF0J
ZcCiXPwH7tASFl1xRM6JdB7FhL3ocm/8xruPiyevxak=
`protect END_PROTECTED
