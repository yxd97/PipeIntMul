`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3wPgifWRl20bK+/eRxOslpWsFXAzVdiyIlyo11d3queXaJApnfnwWhkXA6ZkS5s
bKpBzZSGjrZdca70Lh05IogR3qh8R0B0icfcRT/q8XXUVOE1popg7Vn70zwtE3L1
vKr8NiclnLWb7fO/uouq57Sul2UjIqJ21jO00wrhX6M3a0pC0iiclM+ownmqUuBy
QNMRVFdpYuVHI7IynDM0By48RdtWkzCXlINiSaA57sTbTybLP5jlPZ3F+KNMibaO
5J0Oe+ggkfa5imo794ihU2kIiaoOpAW7SFN7uyVhDXsLrskFxeu3mLgxPcfydmBo
EyF3HLTWBTwfpG9QWixWhRuzgajIND6rjQTsckuyzhNhNYOcDaPlTTG6gZWEKGD9
OVnpSii2Yz+Blv3cDCQEYQufbUaYeDwHx+ocSVH8QOs=
`protect END_PROTECTED
