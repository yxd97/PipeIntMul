`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99zDyPNxd24KfWW0MP4Lxh6X287qm+ZUiSfXfKrM/KNCq4tinZCMenQ0oQgGiFrN
wjzcehUDpv9PpFDJ8EwMmoiLrYOD3w3g80VjU3dsb6kr2bmgHi+QCRZdvXxexQYL
wZJp6JTYWTbb2IbP8/vD5+EmPgOUW4CmmKWVDWmXVyWVh6/ykomjmL+DL/HNVO3b
+yjBFfNWhNOyWN7JEwsVrsMDMz6oexdByFU1Ep/LNiy/9ty4kTGyI7PAf6NV98xf
dOlQyrEWKqxPU5hafNPZ6A==
`protect END_PROTECTED
