`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmskL0EawDPVEQU8Gy91oSKuLOjHEJkmSr+CS2M5tPMzkKJI9RE4xoH2lwXadwIo
AFVRYPGEsM+6v5TeZUnaIU4biA1XMWyyYBZv1BeIWjiHG1HPEHbmVNuAz1TgPdHl
g1iFgtvOxTLEgQkVfHmsE4DEbmJEbcd1bSXzPacKNevoBsdPWeYqpUvquo0BVHNF
YrtUXI+qbqq9Hv31KU6D+FVn77Ezbx2CkVwGhzrgj+SzFhbLM+sjcV/Ep2py5vTm
wyD6aNPspky+RrH6VY7gAMeaB/ezm7M/cNOzqcH6PERlhOsQyNREaURVxtsVGrpd
5zob/vN3Mu0wek7XdT4496BOj3x3UEo1s5F0HIpjTsI3A3RCHzJURigOutkAlFIw
`protect END_PROTECTED
