`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkNswyFsfq5HRGxi6yoqfjxOIKVpRtaku1SM/U/kePJ/1VveiCgTWb1udl/bXMzf
smdcu7JQ7neX6d/eIyGplz+YHdQJpGMg95wk/UeGskjbqwFQ2lMTY6bWjwrk/lv5
v0L0w7If+Wk6xKR/5gVrxyUi05vJGMvMFyMbuHfxus3SAaBp3Orkn1kbHb4zSqqq
h3UI66dm1DdtMjgqlFmTDm6SBD7GuZ4iP0lvSSAyhAMK7FyX8nU8SeOGvyZK/Izu
9lG6nfu2W/sI/9j3K4jDQTMlAVeD24918QAV5QQk+Lq2djczogpRmatqscrZH3T4
WUrt06X3quZshkjuysoGK2E9s5QM1MbQCLN/UxK/Q19Qj6BPJYFpJbAJdivr1eeE
mAFTvr8Kh39fYLP6+mJ87GdXJPhSKgCvGtATBCu4VEffteNFAfvLxZeki9i06aoJ
KrhyQxXzO3j9QYPgx4pPfipxQk/Mft0AP9HKv0lkNSRl/D/gRaUcV9pCvDHdnBNE
1jwxgix8FDgTrryzHLRDd7h0IlVaU23s6aE3QF4Hr2Zb0xiR4HpPF2pCUA+0aD92
hRhdOgtWo3H0GjL5hCUxq4SEcFn0Vz/rdWB7bk/4wGLJwnaa+Kra4vnbegDMpqCN
S/WCm8SaRJz+xn45xKslz7ej6ZiHY/rTL6GB/rwbO07LMxj9jWDne/v94NvoHDyt
QuF40UAbHAl3eltv0x4iWddmWCeRxGhvmHtcEYQli9ss0LiJr5N2k7TV5aLv8XLB
If26IvkRRNkiefyWUpo+oJDSFuMRg3YRHA5kMVbx1J569Z+gQfX2JJ6c8kFSU31T
06vHE7NMODslicNHhEkWYVEydMLLc60IgX9pxQpEOkEZ46vBJjIiHCYeVKgtGysz
wSDCToIBHzjAJ47L8SJIpQ9voEpPpyv9h3eHs4dGkd4lz6fW2tFtqzwfEDbys737
HIwWWX/PBRQ1P8UjvRv9SsFnn2w+yKJoqL2CB5GHdqg=
`protect END_PROTECTED
