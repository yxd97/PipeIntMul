`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
879lSCvLcmwWlM7aLnMgxIT2/hDN35lNfQB1aDNVKczkMwFAovNUr4YoMkQbatsC
fVfAm2hwKq/KeFufdZwvhCw9C8y5xmVUpge7+9Omr/kjB0L18jSc82UEsmAqCrTx
/K8w+LGUdF2i0cIzInxrmSGonh+amlIzv0IwK+yvMR+RYJ2+r909y2v2ZHzB7LaK
SRA7MgYXCWR/cKqV00uj60d15Snw5UwlPOIAWYZZduAy6DrBp11VKDWxR77BNPXw
`protect END_PROTECTED
