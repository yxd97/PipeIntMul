`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNcintPQMY3lO04jUT/ROzl5RvOXCWdMAM+y9F+1ZpKJMsndfYyDOajFnXbbF1n4
FNABqrKf5ux7rrR3kxtC8Wv2DS+PMKLCl53loOik4Uv+wI9RyEkSBLAycqiHIS6K
aRtycV8RLBAN/lVLC+JmzFq126uNJhnIHy+WXuZVij4rdCjEWwo5QLboKNle/dLU
A7/BJwa7CnzDyxekjLUquvyDY6sF7ZwaREhau1ZSSkG9DIoGG5x3FtjHbkz3YV7p
dJ+c8sfjcumbAAffeft7tVsyo3LjzdfFkZSrUde7wAIe3uhEbsPVrMuxgccosNM2
W7PeT2pqFVlyUEusnZR6Cl72Kq0BZhMlQJoXaJGfRSC3jm99RyNHPqjivEVWPIp5
oAKQQe3+IAyaMcSc/V0TWYxw+WwPTf3QJJCpZjjcmH5/dCodCmqgcxkMC+T+jxcl
gFCumXTz98PACcBx+lZxPBjugY/mEOhYcQARdDsgLmWleQCiBF9CtWl/uyd++BKH
Hf9eN4XvDC+sjNFOZpsVyCL6fMitKRZlUx3uv9HSkJoIAJeAqIeOxBYy8Ib5ZmD4
KMQOan8HfPyLPlBBnr2uQQAGVyGRjl+BUTvRk4TtH7n33PLBwNYnrGbYV/jPZMym
LnEvzlYDatiblzpJ0GAo5MKqf/Pf0bmnbBcu3FbiTZmiiVWzUJh/eGiaeSbfbEj1
gvRJ3kwMdi9EY6dr6cvc9+g/BshheAETocraS6xIaS8yPTG1cpxQEqAuQXhKV4+r
oruXRPpWIAzVA2yg8PdbMJgrcdxRhzISbSUBbwNIrF62vh1XRmgeOvSs0rMfQ0hp
cG5JjJJ66CFZ5B+3w+rbcXFyWNQhwmdrb3w/h5NjlVgZtn8PTB5Dt7Q490kDymhV
mfPNPqzLpugLKqOTEq24YimuJuqMs+XXjQch2iqFoALcSh1FZ9tlgX8FC7bkP7MN
xy5bF+w8RZTAeYi2E0YUbRmlUOortA2cLiCDXZi5heU=
`protect END_PROTECTED
