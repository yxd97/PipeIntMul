`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
plMFYtQCPOXBdXDyUkkWm8T++ww8hCQUyGZoMA5saaKlA9CrPo4+w0cbTBqfInL7
5Cqr0W8c2yRK0MyX1mymV+BpEwXZQVN2zBT909GXD1XFOiIyUl1+LZ/3luXJMtgm
0Cjmga9NT0eyGNjv6K853U4BlMxHynYoXAYAQ+JEZ9uoBcQV+RA+M0TRDC7RX3BQ
DSzyHjXH8vAXzKvqJd8lX6HQWDSiUhVwDBJgAIV+Fi6JPyzZd5Snv0EENlwp2oBP
4UmdBXIaFhv60Am0Zj+inRHxKvvsjZuRI2jldWsVVoGJwigItDypeimP+PP7MrU7
048RY0MMWx+ZXtzVcyWh/BkisFbL492DPWILG2rnQFYC4ryARH0Hb1OsXWNUisE0
nSNU6It9tjZlbki12wRqLv74qUww5g7UtV6t33mBTjJgCWGkUXwbD+9MeP1bnrgU
fc/HiJen4+NQXo2c/GrCb3FwKmbGGRHqfaF6M01BLJ1b4EmpAxQghDDAJaCs32so
FoVEE5W6J6yqfUA+8EsYq6x5Cd2XA4zbS+2FL4cc/StfLJMkZHFDWrl6JgKvfSCJ
i32S5MC6RGCegCSt55UpBpxds1R0Vk92S4RvPZBe/mg=
`protect END_PROTECTED
