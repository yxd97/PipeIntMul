`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5lecsKbb9xFGoTVSow2kh2cVWs690Knj2fnn+FsJ3sZUN/uM0yScYtuJ+rad31/
e1UWaiqECImofRa1v/h9tPWoNLdHM5oxRTQQ0fVtuM2u44I4aj16NcNmMj5N5Vkb
RT8EpuZ6Vmj+5fYph+cpmXmmpynUWePG8zrU1hJiWO0QLHdB5nFkOSa6eaf0pvUS
tHV/7AOXAZ88DdXMk+wE+L6iW090yeSvwuI2UxLoi6G3g1Y3MDLLOoHwNix8zLd3
QIOyoL3adbwZmSoP16sTYOoE7+Z9MMdWtlIgNrr9NWZtURRNi0vZxSPLiQ9csvO0
LmMg8VXlN3goyCXOJXog3wWVyV8KJVT17gC+4Cyhh5d6+NYBs9ESrpP9FI0+J5s3
UO1ai48RVu3v3apPETZonSS5PoNNKbH7rJXHkXiLPxXffrCQq1L7s1X3gnF9p4Dc
t3VWQziEco8FrPsUXuHZVNmIaTMXdV1C/LsTcE+lt+y4CFnM4dAASSNjoUit2r4o
xKfdpZp7IMQM1cTwcpr7f1lbGyxIB+Rdj4koPbDqZrFy5TB7elvtt6IO7FAQMvLR
48KhCuyboZid88Lr1bj8YgfDbwhbhEOE4TDRRTSc/OmBfY3NUT+Qu32RfQ3mqi41
xrMxjoWN5IxUCswhK270hFmrNy/skbu4EjpEa5zAC9CbrLVGNifuPdiGFVoXy0ag
w7Bqvw3bgGw1U0odl45Hajjjcospjo9bUuNXUtc+M6YXD99MwSse0AHhconlwY2S
lUhCm+BryvvEyVrKFF2G/A==
`protect END_PROTECTED
