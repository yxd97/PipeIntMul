`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oLZJnnCTVpnwOGYz50p5zNYLx5lcvyKhn4uBcFZG4uvlRwe0WJLzVImyugQTgmbf
1lQLfaZy83ln4P+Ijie+iLZmA26gKu48zjyyZc3mSBaEpnEkNgKL4MMuCsnRpJny
4na9vBxKyvBLSqFhMPFyKC5K4k5jwz8li4fhy4Y1YKb+ipePblRMkhOlmmhchKr5
0rPD+iCRhc9qudK3NLqBQVClv2hsAaHVWWIGfglG50UQ0ZvEiCYl+XifLyQ37Fgt
oMJre2QABPvABwf8JAv0Jn4pusnfPdJFl1PF90ST9KmR/xW8iCb6/3BRGuSyOJ/j
8RTmABzyeS1068rgnOIEY/OEgW/0cvHd/vsodNKrmSF0dGVtEVWUGe3fue+V79Ey
TfeXYuHMqyAq3jUiyRVNAapBkB4IPlwxV6AwTMhbx0pF52ARtlUH/6tJGka31yXj
iMujaVHqeY9V/J0LHRsMgHWoZcuwxbjBD04QL9xCIIvrkQxxaV+1akSW7tf8GUxF
CG/MfsN/TxU9Jyn3rkbOwazL/XTb+Tq1MRSw6q3cwc6P0xeK2cEwH2W547c5eVMd
AsB0ilMQOve66I+5K2jkF5/H5DKVraWavpA9LyYXNq83a/V/Gu1TUaTNfk1k24cB
71Eq5BrTnHl/B494lXMkb1tL9Xz4I25M6TbzoGIdozEBcGc60SW+1IzSNe3jcaQw
mCsEJiL4do0phYvsxpMWeMoRNBPKznCK/0yueCVeRRftS4t0MQjN0MUMu5L4h+s4
20PHYBtZwPr+Mev3ihxSVLGxtdT4uwMkTgzlVSWFiT/t4LVbuef8+DJQA0a9vGLh
+Ri92EWWlQPXcSdakpqI/egF8ufUrIO4v8cF8X18dmuSC/aYfs4lUjZYmQC/uENO
Cu1oijfQrUkf4SD9FtJaFq1o08nu85X5bbxBjM7YGIbaU0I5rJfVbczv2j/1MHCf
9k2j5xsdgqd8DwYsUR5vnd1bYIeggsJ813r3VPu2HvB2FZnsXdDtTL9pZEn8WFUt
trnuarWTriMezGFJ0OKiHyoRloSDfL16npLwu0XIHIH2qaOpEnpkvbeZOna4JgkW
FLnq1qQ8JqGs7/6DP2DPhDWpuInkltqr9DUmQSE3tItxdxbJQveP0MRN4EmQM0/t
m9GKzf6g6aH8ldFYBSgKWwxSjQiXfNL7TWXlyCNwg6pxzx9axt4QQ1qO7rOBtO4O
4rGrbRjhEJiKp61YNxqqVfJ0UZhyZzShgqtGN6HviZc3iPYDJnXXTaAMqA8oKJbk
AkeeVd1Fs2KysT4OWbdQqZe323rozZea4GFzBBs7hKX1AKhChArFcgMgrwlXCwtH
ZyLnILkL0CCP6KOu9TjsefBDSc+qm0kCej1+mTTUKYitRPNqNrhiOeb58n0qyP3t
BU3Y0DZ/JvNxv1QVGBJTNL1/GxzWAEe7lsSsC+KhNihs1crYA7BMTRiL//o+QUUk
YNW1zbKRZxLYEIi6GdFpjgTGQoXVRFmySlHKwuPDOrwx6N0TaZdDzqXSFee3Ygxz
E3QNwIgSrVIsqPLRShEQJb7uJYRzcrhHl8Elt30wRg8vHg0mVT0tdIk1QLEbGGmo
tNyVowfuVsQkhJELqrSO1MQK1l+e8VVdgutdQ3D8nNYz61AVhwl5GauKYcgYyLIJ
KOiPTESE9lAVtw1P/4v5HSCIPO/ZQbWcZV1dFuouUvF4HYpKaSGbFTlQkd2Y0e8+
`protect END_PROTECTED
