`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrNVJLIzkOPd/XzcFoVxFM7bUIELkxsNcB4UzokukZGMK+EIX4pO3u4SpQ9N2MjC
PzvDRQPvP0hdPxt8qP9dOSt3tMhes9qjVlx0ba3uCS7OQPYAvPGVKJ+flpFuiUOO
sQSrd8mnw6JC6JnunJ7PwlyBd98Wz7t178JnoAFMlfTfo6b4M9thakzC19C8fP+V
0sRX2NcuUoTIkFgCW9U2bY4fzBQDHJ4jK2bnpVYYzr5p02QGvJOVEMrNkcigroQH
x3pFSSCm+4V4tuYZ9usmhvtCxwfWJjz0H6dx2p1CYQEcBztvDQ8j5CBmPTC9lnaw
9a7grGMVa06meIqItQi5+6fcWq7ld5BdcFKL6ta4CL5AxfvSBCo2OSsIuqkM5M/a
qiYX/KKNN23ehEIQXaSE9eWmpIMONa0jM/95oOmu7iXEAOZGELfxnpPzW/rXGtxv
z3xQclwgeHyPVD4o6SHuGo97QlUa9blat+XiXc7XK4vaORyaGmDygHXb6FhuAusx
vqHaQdUE8hw0NarzZRVDDIQ/a25AkA24HGgeRKV5RqAOP03zwlvpAwbKWVxSiVyR
Nrku17EH63/D8f4L0E1eDPecohJPJS+sGQgngl3DHsy6KT6yEPu3RjeL4bmXTzEl
1f+TSAe4Moz36qFxsOgaP5Tvj0aIPpvXmF1E3DjCg8ta17qOnrGm+Lg1mHS7p+fH
nXm6hzZ+XzKTREwGaH7lTXLrbqsbFN6zja01+M/fA8frZ9r0ovIoR8E6Nerk25lK
tMRlwACC7rGVIaIGkETJItV3WmWmlNKlC762YAVdrWIvy7DozHgh6pHf3Bht+kz8
B8cG/6jEnWi2ktx+8adBMdjXF+6fsi8G7ib0Z+9UXVr4sEaXfUjjeuRWMFu640cr
Dzln0wjLPEz75FQMONVxlhDK+tm5E7pAHai08QmmTdhC7W0L/7bdGKSYdBDqM0NZ
uMVP0+98YBhXC27wi2BrCicdEKxJBahmK8o6XB/HXkdfv1kkkBjvUCy2mcSAUo0L
k/+xwlONXUjMTgoSvcNRjQB5YxVw1R8QNgskNxK69ULTxtUWgN3xMzWUWqsI6mWp
PXGzciJJodRIw0wEfjso+w==
`protect END_PROTECTED
