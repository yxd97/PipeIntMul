`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SbBxhjBQNEeD7nzn9l60Ml97W0pKc09Et3BTvQS8AJlQA228aBvqEALyRCZMa60U
sZXdIywsIdgMeq/FO1VTuE2wSgTu8CV3mZuo2sNcfH+dVyqQhUZcgtwKWImf44aM
IGL+kxqhMgvTw09/8HXE4ZeTQGVGVqCJaHPg2ijMSPcOi5WZ22vDn8We5DSgOjzZ
QOcTgOEZHD+AHYyi9yHF4CObJ+Vp4GtW1L27R7+TwTD6CWAYn+nlE3cnTza4WYfu
H8mMg0M9dZyCmz4Z6o3ACN1G2NOeoe0ysGg5TMhhim+1FLLuGFgM/346cMw/7Ko6
BK7JvJh8FHVhdSOi4dZxMqmS/nNgN5Ha/3j4wNzqytXy4Ay9JQkc5x+xQCTM7mPB
zZN7nC9rI+l5rmcMZVQyuTYe3AK0ZXOcdnWKe+YCKsr6zum4V0HFXDcAPCiw6gQc
PFWXOAxwDNhtsni+ohopR6yr47r+hTI827Q7wPIL1RvfI8NLi++O1jYsFKKnX43I
gUwKPkatekzMJaOxP03inE78+jwmolfPND1RRPH5VIlM4sccx8qTAxD2SccURozg
jB+Yq8Oq/t1FzC1zT4NdOpZG0cEU7tRheZtPfLi8+EpsYmdPaA9CWMaJQO0Z1tYg
O+j1SALxVQP8Hngn+HKiCOBrId9qDBXLx31Hah7SOhd/GZ1WXK9Jifo1VaFA5Gap
FF8Xa2Kl2Pp/TnuM6Nkng2FjrbPcME9KA5sAa1YpyYc=
`protect END_PROTECTED
