`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWBjLv2QMxUg7d0jkflwG59/tQbCqZUkU6TLG4g1uEkwrZLegS5d7ZITupwEPNOI
+lsef92L2j7onQueWk1nzJKifix1qJMASNJjyjbLY/BvJvB+9jFfj1fwXiJKZZY3
KdMk7632MUFO3z1Cu00tqf8X7W0J1EfghXLPC1y2xdpKcTx/tTbvortsbFAG2Zoi
WSlpVRaQujcrg3z8If2gepHF0jexxo00ZV2uuU+isR7CBb23PQYy3CDc2wMVzN93
OqShr30gJM9NPtIRbpbKkOIoGs7ZF220whI1dMmmGETxKI6FEXvK5ofwB80tUFLA
5z6XvvOuwB0UdKu8vVhZDu/rYewFLg+9dSmzEhFHSvrXQkR4W7aPsx1sOKTbMwiu
jZBKa4EIvLhKFvhyRQV1u9jXI9FYEsj63UHaarxMbaUH8icSbjTvSPkMvg2Y9vQ1
5USdsCibVJnQlx2NqLUKBoeQgbaWYLBzoFeaAww+nmLU4pHI9VkFYs6QVUIooX6R
t6DDGvBoevIqb4VP/Kmp71yHmwAe8JYfcKCe7+BUJmPJ+5tI+E8My/IJoN531I+H
NdNfmkG47X4VjEgGuXp1F3N3reopQJqPz4x9sUbxCIMiynv3kmQIBc4k6sMuHhrb
WocmG6F5RHMhsvcbPjuc4iSSagyDcKMDi0x+r2rMQOMvv3pHwJruql3uUg0AdHXg
PQ+G4ddp6quhFkR4tGr+NfNyCfwPCy0awt4E0vv3iP8lUjGw7Vw0N0heHw91j3d+
trdZ/2HVr61kRgofh88ocXeedumdbYT7uahcbHuOs0p39aaT/IBe6tdiyMl1vtXO
izBBjChgrdtod6pYQzHBq8ck556v2KlndoS5V5RUcsheqnW4DskyvdIAq0DFDLhx
EZUNllNnpwDW+6BJrdrkjQdeEuwk/Q5sK/Fz1OmoaW9NOCX8DeZU635eN9gqL/ou
IO1cCVz3wqjmW31l6w+CVXa4KtwZXIKf5JtRvHAgvg4x71GXMncmXFnIQ8/lVcdO
`protect END_PROTECTED
