`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/1bS8QQC+l5/vR2mexZBfnUmyZSLnLbIME9XVGBpQcuIovezJsZqZgMhOBPlyfaC
S7NVWpf01hhiUD8VjtnMXEOyu04HbBghzB6v/LDIiqENhM4SfkXF3PJxv4r/nxs8
tzDvxsyQaVJIm7+5WBsbCXLCHg9sBsgtWUaP3OpVNfAcYo+Z2bXcXqjckbkV5W0J
okG04/gbC0+WaLmQzVnpvPxHRLuR2zusHhJF1GcRz2DVRnGmT9GXu7HRgqroevnK
YG2W5+ObTsI1MhRXX8dkmM5Y7LTarJElqAhzTnJjBmkjUgzw3j3aYSKj9j8AaGK7
1JuNOQkuA2p3jurHUDDUJhG9kwCv9PfhhSQr1oOaFYooDctiS6Ws3HlFZlBRsOVM
+2wZJhcrfsfj/caHi0n7wQ==
`protect END_PROTECTED
