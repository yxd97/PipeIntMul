`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQHU9puBlQefnmoVr6NyLINStuLCuimnb1Uyh9XqpbOeGoJikqncr61hugynMuc/
y3VRLhRF03noI4emziskLPTvN1hrnzrKvNTef1s3y7IXxPCOrOzkf3HvF2tHTpTM
JmUayIy4ICNXYNvO/X+QNn7VBSxIv6NM1P8nTlQJdpauB5fi+4Z7KZJuyTHELeSV
6jf0UZB5yrdjX23zpDyaKpsuVfWDRINr0i0s6SHZgF6Xbxhg6asIjwWEI8++lVMk
tiRorJIN6T2Usdc/vEM47mTVH9h+qjzRL5kxuMV7k5j3dQhcVAXFzFjG7qXEPl/F
Y5Ojf1efir5Z9L0q7UddfA2t80HEVRj4fiDCvrqns9hLNLOZoFuBBzpnNO2r40lN
VyZWvMJMuFUf4LPJYedBwcOcEfljn3yh9eEpDGI+DsZfP2p9OpGfhHUcHuIC3A7g
/l9GoIHkm70mVCfsMpJ51p3mh+Emnpv9i6Z11Fc1QmIcNPh199A08B/HYZdEDB5A
1XDDuIwgfkxedg6zcP/eGi1Bb4LvvN4vbM5SSBPunOCX+MM9iMoei+CyITBslzPg
ukTpWH780mi5NmiQh0LK/W4qD260jgG5zR/Q7+lqu2WOuOo5b0h4Q7cjiD8Dx4lr
PhyuetGbS7Ilp5/LZMLO8pavy4DlEjp3SY2sYtltv0ityodhBylcjJ+2fIl/eEIe
8usaV/Vx1o3T3WWUwo6dxFnfkFfSBuuO0covjNCnl/XQ8TXAqrjbGu1Y+iYMp2C6
eqitHdr6wDA6O9LqdNUv5qfGSrlhRJReCfYsiCv8p2zj1WYCXGYtZ9bXuv6SJVDk
MLsxz5EPUdYCPqwiQPVpM57kKJoM1oO2JHQMLt0PuV+qrwhlblCu2gxfC60rMWpv
1xYFlKj72eC57vem0R9+Xwy/UBe23XLTwRa07dc8cdaI2N3aakCXvMt5IgcQQXwN
/KRpSQAk5AqaLeNSz3ZniiTAQqZdkHpfxsoNyOVRddHzO+KwUvkk5AQtq7AHCud2
OJZLcBVHZIiWebnNti6HZtSJuMTTbS0avgA75AJOxV8T7m75MGBri4Teg9VhITlC
ECV5le6F6qK+VNxwEFog6l5MIR82Y7HYCtvO3nm+3W7MhjZ02lR8Ls+4Siok4v8l
4GPGkt9nDP4OCFnuswCZZcfs9P34tl3L/WG+u1HuzXLZ6K6uPmVyXkP81hEYKJtz
TJU1JLwIhGUJAjfqbLAcXYLQzZXtTJ+ajlWNaO7QvoOgBzPm35lDDo/IQ14ssM/N
QB8VU76SgLmfFBB0iBQFx/LHWiOt+naniwM4zCLZz43e4iFq+DJ0YXgWHuvW3QCm
vuib8rTSCUsqKYWdF7F+86CsEC0kfwSjiqIWyKO/yIxBH19pbTtZz1FAHavvR0if
Sr4hEvu+UWhbuu4SS/q9PuPmKdtcGzBHr//zp+GjUDXmy37F9UzaQn3ML2puX4m8
idgVgE/QOEBNj6EqlJe185WsMcA/JSdO20RdTviUfoIAReWu2+T56bMbBQc3Ymbx
XY1YJAAXtAGbWKVkUdEu/SUKNv/xKDjZRB14SqeA82jReDkygo3IygKhJo/FTuwI
wgej6G85N/SBFGRj8AmWD5HovHRS1qEaNefp5P4ZVAf9qTiFJPS6+To2NOAAPo6a
nKCewuWfFI4le7sEpHdB08UFG5Ikhg9fC1TkbnC1JhLMgSnliM3LvnAXhue/GyWo
LQfbbomXWs9pBwGuH+UEfAnsEIDqw9tq9E3OgfXgN/IHwRIjOSVNTdUQvY0ulTb0
9RBvKFFeumm2UqF0oCyxANb3TMto8/lkqNP8XiaHJDbdPEvzeEs5yJRNJM1llX85
l6QNwJb2u9OfQzv6QeWO7ErYQb8ufdloANEkDNE7Ztpym4rYQ1jinszhwD9rTbpC
qaRd0hQieFHqMQWHUSzQbenncAXMzyMiorRaTI+dV98YTjC1ujUBiBQEN+Fmc8Nq
9xPr5pkHqBX2bLc2nVT8sK8iKhUOCge+ymmx98IbTqnMSVo1yZeWJtvzjuvl08Pp
flrj2M+oVRwAN6D6k/AcRgH3GyJCVNy9Key3HqnKH/aqqPrrSS20bU3CSwvxSghD
T9j3wrfknu8CcwqqevJloMWHPzx29+LQr6YX1pUVuRBPu8wCF0LcejcCAL6lwHx8
rwpsrVEYB5pxJst9Gg6sX4NotjLrbgBHLrfJEAeLOvUU7uw9p9/fJoP9db66vIUN
nZ7/Vm4+51hGYCVHInOygHO3S8oDBSmp8hD4HEHhOzUlnzlXD/fzILgldnjJDL45
QUn7tKX07g8AG5uZIz/qkq/4j9qi8AqetKhN9dhoyncjzdIIlFfaAgHQqYbLSy42
LdR8ATAExxd7CP6ovNQwzxO7gM6Sle3Hx4y25WcNND7eAwNZd6uQQi7M3RcDLybS
laGWf613wm1262RUgLHFNFoxleyGjFGqRphjLvrPNbemcykmdRoeiU71cPFVULx/
q22786EUElijg5fIpOtF0AVC3/qkMqcvWFnqwFI5y99+eCrbiujsJOyA7ive27pv
07s03W6snsilhKefWbRmJ8uC6TOvm5O2uZ+kefuWpetNlQt8vpeh2k5NiGWphUE4
10ka4/dafEU80nw5bvtyDwsz4BRd4uYinCiWU6dw3sInNABBwEPODNYaUs3gLDlG
ALvwcv6XBD3GVOWB1O9HDHd4SPzOrINN5GO70qoYseRQKxO1vzDm5NioVh8rD6lV
c9jhB6QUKfx90Bqv2xpAVC8O6c6fl5Du+BXYFkIgtc4YFZnZVjB0qQqRqa6fsMNl
7mxnFNbETLqgXvPWtCknPKopAg8VhK4brmcyZXgw4L6Q8sY3F+KeJTP8ar580pO2
bq/8zVSyrlfTqLjTevr4wPqBNDeQrJJynSEyD+Lpuoh/rW1742Fe2GiFzoesLzsV
LnhZgjUFpz3cGxGHWSTWc51atcRDy1aFGz93MYhGNwaZWIQomn7s70uvgw8poVy/
3MxZCLkbHqpjw7U2q3yRxqO0TEmuMhvI3gxj6vg0Phj5aXPtEliV8hUsKZ6U8RAc
xUfPo3k2L94heLITNp/gOl7ufso2Ph8NZg/bMT+snLycLs2RsxqHHjVVCBSZtuRi
iLe79GjuiM4V0UY892RledW9AFX9v9OhdDytJfhDZ4fuvfRszimdEdm23ki+FkNj
xbbJnUrqzD0Z7TKZSIXofxDCBY+aFUOQXk6e36bboFCZUvDk8OFMUFvu6ZEb+zez
0DgixDvfwbaVTLG/GH1J5d079iIPxYqVn5xpvIrbxB9y3JLeWJ2qe51DbHhRXiAH
HkGfaxEo+4PrgG091LoytXYusQuJBZw1eKwJ9EHuZEB8Cc1aglQqviUaeRoHDt3O
EAWOTG5MxPyIZfdWrdvRMyH6dupkMHgk4dTz6y94oVgZroot3NngsTkid1ILINWB
MEZIPkORVu29djGKXj1+bJ0z1zomMxrmMoXjMnu9hH5vXLXbxuEsK/mA61b7bzFp
NxlK06kxDXgr8gICUxDsd5lXeiz+mR0MdrH5xUpNpNp5j0EFNzHHyZcD+gQG93Lo
IOzJ198BvyiPwcvEMWQrowrDQvLf3SIdDvep/9DzaFlSOAc5rzG4DpKunAJyzPRw
rS5MLTw0RK9O/aIBWeINApqjDkX372S84PNMBth9+PgS27gM66wFKI4L3asmEv0v
vfa3OcsMIsgZrfYaSrvxpltogOW2KUE9B0gs1LljmMSyLqjxcMcStjHL3ezmrPst
GL95gD7gbZHkTSIta6SI7lS7Zt73RY1E+zKeqp/TIkI+HJdlCSyrIsUg3sReJipr
VZmHI4DyRPSpbsJjiQFLh759/sFEY/vdQSGZ1iu2HfbxngSXRLSDIUyg2iKRrQdh
70hkJqjyxTwYoJe3amddy0RHobu6FXNAWbRRVvpKEjrPgc756RKs9ElNdOPQAmEL
WubTplcjeMjs23O6gJSL5F/fc7YoAIwLQOocWqxhvVER6jlYMcOZCUqCKctZFyma
MY5f2rkL5TtgFsx56PY03NYFcsC9lFj/YseGgSnWuB8TSubALDMMcMhEBenn5am5
eInmBKxsl0jYC5GslqcyGcwarazPoKDjxzcwsIYO/RPgLuWZhNjk8tQPfS1KLL9P
spo8kFjH3aUIBZR0wE3WNXmZrWWTHjife+0gfhSOiV5+BhdvJvA6W2Znsl3HYWd4
PJRz54NQkCbS8Gl6PraTQ1o/e+oIrSc4sGAuha3fLjmQ8hm9WYlCy3MM2Dv+xexQ
dEziZ+C1KhWboVVm44H8SJ0HClmkHlgjxfuWh748Os15jarcQtU2B4k5JNr3ln6M
lHF6OF6+OyHxwEoz614d/tnzaMyK2a2zJrRvWPu15jTLPBujkQzYZTJaaE1vv5kW
kq6milgc52kcaP1vRSkST1Njo1P3rlGfKARH9V8xwFQ+vZBXVYGpScB6nCwUfcsK
62BLJIpT+NqDDjd9b5VL7X65iAcpNmJyMBdhdFOI5MlKujYs9Wrz5gDnhfExiMhf
GSIhUtHEFIhj6UDewLlRPA5Ic5yXIdRmIsK9OdsNZ5/mbSfE4XzISu4KYCpqS07a
rvJX05hOmQsR70VLARg2sDJZqDDKJ/rxvMP5DYVUauGSTU4Z7pwpDEFn5Br4B5Tc
lQKPNXcsYCd++GbqB76RfpX4x99KlLcaMYt68CKDq3V8dFfHfHHvu7C4lvZK3mwL
DwhJixEMmHlYNkKBW4xANw==
`protect END_PROTECTED
