library verilog;
use verilog.vl_types.all;
entity IBUF_PCI33_5 is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUF_PCI33_5;
