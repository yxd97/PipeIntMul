`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p2HCfku4mA/r3Vvazp62dni8UdsXeNUdgnyUlo5CQHfjzRx0chgdToAnFa05s/5r
kk6SaHBiv26BPxALlzFuU/VIjJwOMtx7BbJ9NcNLeE4CkVA1GV3u+6scm1OLsA0+
3dpXXAfMh0EKymdf1Xgopynx5t5t29rlwazmZdVmrOlPdiBd4xYeLybm4RmdeuIl
rdcQtsWSpMoR4qMq2WS+FS8bn4dHENgjHzgPqJ0LQaV4k052HDDQTtrZL0ZmtxCx
oYKhW7HcBEFv/oLZeAs5bw5QyIkT0Bp5mvZ8875JuWUD2Hn15YSaetS67YvNkh1i
uAJFHbesEOJr+NfqyOIkMw4FGvZS7LZ/N8A7v8TQvW0x3zo9UP8NmWmX5B+5vdie
+/DeJm5cx03a8GnSOCyohhgci6pXCaJP1MAS4gX6AQvoycbr0FJmsCRcHG3qRug8
Twmh7LQGH9KLQNhfwEV2C65dyjorUNkfyKs0PXpvGg6SSJdbZuXwOOFNNRKQDS+J
taNqb1oJDtGz8VCLpWmh8YK3tGMCEQKATmOrD7GhXQ2wq7w1BcTJtZaNUa10+QBv
H7JimXoeWuiul8/SzvNHkw==
`protect END_PROTECTED
