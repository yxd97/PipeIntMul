`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMDz7l/J+vL8wqVdX1Zhtfy2Qe2RiA5g1Iaqm69tNzO5hlOaA//NueR2+rSqdEJ0
jad0ZYdWdfLGeRHq6oRK+PinL+IQJQSCyN/CuSx/cnjA0XabweV0vaOrVfhxdsxs
at6GXq6i1yAh/HCdAB96vPyDs59WNqBl+D/BJreqnqJIzdbEn8vtsBWl6YOWCboG
XwVZ9DQCsbgTcoMOhKhZUtu6MQ6GrpVInvVXV7eSDuTwFw6mUD0lrKDwj0dzd4cp
E9BVJ9grW+GZD947t8RpxFWMwK7OsmU+V7sKXnL/d09BOjX9uSsh59tnaY/PG9Ld
IcKPlee+sB8s1EOMuLOa0Q==
`protect END_PROTECTED
