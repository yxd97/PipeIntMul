`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
us1PBRjCyr6VWVnetpVXqyowJQx8/GG1Osj6FCq5kBtu/72g4eni5ianhFVBU+0f
jyhpXa0xt7knzZrvPyqYQKUO9nD0rChUWoK6TH5W+RidWdxyLR+uLag+SeVGywbE
q5S9JfWCBAW49xYkyXVvNBncaB9nELbx6N4LGCCmKe3TrPnOeIXAvTFny7ogEnhl
fglGOzlB+40A2ogDVsSH2dXgBQUvYJMvyr2LZ7t1AW70FvbTf0zwy+UMeqUjdNZS
2tMwP3wfdkE35rBb+mPQK1zjWvntYuhBQWFUMWO0/VOoL6lOuoP+E4qSIiROIma8
N5HrQ+/TPDHVzFkrpw9EyVUPtmRM6XpOylfwh2484T5sv5t5AJ3uTZ+658Adwcfm
`protect END_PROTECTED
