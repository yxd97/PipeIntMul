`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZOnVUvVZ5ylQV+Vkg06SJ5cZmt1CRnYNCdHJ/50Yh5zEyZJFXZcBpYRfWzjtBox
Hbvy0sSD/hZZDJhrq2rNHvLj5h/j/sFa5L59jDgadXK0kmPmaKV9jfcfJPkaqwdc
iM7w8hux508VBB48TOVPtDR0unZYW/4ReMB/2l32oOas6qKYZs4C6qvMZ7RwI5kz
aDSvcgfKuM3GXKqTCvzM8BfaXrzaH/Qv1is4+ii1Qh9Av9kIwnZKqenjtd5tQhkv
PC67dcVcOg+ykNANoe8ZTI8sLHanfUO505E6wDceVWmXvQAzyVcP/r9Zix5dIkFK
oZgZjbRE1kGqtgGJbLoiNIYWzi28Wg21Bl4L11CjGYuq5sV+6G+QaXDrhRrE7l7+
KliKHZLFq58CrLUtLXxwqYwA9OfJPzcYZ5Z2P3K1PKz6zyP0yc7lx6LFIa8SYnuz
vINOy4np2rU2OpMiMuomdBd6qRMK+Jh1g+g56OUYBqTW2NGIXJfMWWlOLr/6cgFj
sfqgxzlJnwPpFAtE0q6ETNoH+dp3m7Og5anGyYXQAS2ZJcLVkQ8Qho8vF2yBeYlD
x+1Xxo+FQy6aJFfbwWJL4qQ7WvKNY01Gg59kqJ/D7g4qojFrooPcSgLORlEP72wQ
K1DBsYO9Yods1Wmn85kAp+fzks2yH6Zp0RMQ/j7EP9fOn9vmxaLEURYry9ASJq8v
qUPqEvJzFv818j1uBA1Saiv9aRNS+jEvZBjv0pz4Wry8GfJh9zdBXLnTseB33iUp
VpsMBl4La+DqTcLItzdYf5lh2YmB85s2FzwPclQNswxb9hsNDpqWa8OAeceBRAIv
q+vbD+hmQM7CTfT5L14aBV1g9umDwjS8UARfWejIDNxD62Lw6lmfPfaI+fiKzUeh
L9+5kx4rlBbgwg2WGbuMegZHtCZizH8fcLO36c9kY18hnaVhEjWKTb4vWwfMwXug
`protect END_PROTECTED
