`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KrWzKO7FM/0mtpojRBH+EixwsdNgceW8w6YRLFtPyCQTNGRMLFaiutGrh06ZrJ/h
xZpf3DA+v/AHLXEYbhC2JEPSHcGcntIAaMCot9UYs3djaPPrqUMa3W4dwduwfBWM
qJuqPs9quDo/i3iFjHgT/Tg3zK4r32ythAaz6NxHiWHoAMJ5Qpwi16NnLm16ZBvC
xSDYmyOd0lFO+2CVuEtIPvaI6lZhW2bTKo67tfVfCJNOg3HfTV/50mGrUEN/Ti83
RJJTCZtK+YFdqma3G+2VsfgAdoJUasOwGQ0CDChGgVw=
`protect END_PROTECTED
