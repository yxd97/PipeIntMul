`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+DHpq8tvk6SMzNrjZ3AlSHJns4RssmCAeYd3dL9wKi6Wd/rww9hyom7/HBwSFrhQ
IYv0hyUPCx6Ryz3/wpAPUzpDlSpgzBzYCAQEfxUSGBW0ETKZPlrRMkRk+h/cIw1l
28lP6qdBwB5x75XhhZx6Bx3qgEihFklgVH1RaEYDe1r9fvY2fyRCIHH+Uu74QXYL
3q9aH0u9XvegfIRgtqBb6wg/DCK7UHEp9+nYfCqE1Jf3UfeA7ngzgN/z5RAXUrEy
0v4DNwOnCh00vWKmcQj0mjeILeDLyb3OHhKfURv0mxhOwLlZp2h6HRXDXh8ptXea
l9pgYJA7nkW+FnOIDp5VJ3tItrLfaWkU0nflZu5Uwk7OjovbSdQ3H2RTzqDhfaOK
kM86Xxc7oYxBXvbr5EYIGPYBuL3ekvUjg1pOO8k14GF6Jo6Rkjmpr6IyC0BWqz1U
ow9Av5lA8L4vKF0wWwn955g/BpPp6Jo5j3bQA6HKtnjrcn157muX8vvZeddNls5W
`protect END_PROTECTED
