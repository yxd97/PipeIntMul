`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9TJDEnGPh/e2czKJVoEvTluLMKo4jFrgZf8npM37O4X2k3lf7NYm0mNlwcPej+r
PF4eaUaIoYsqw1VdzqGm3h2kpyH4cLqEQwXfEZOCJGPXd5c8rk7L+Rd7czwCA4I3
gAre0ndFiPxhieY15wZ5t1wjN1xuIya4A0R3rnzSsGbSAosSgXlTjR1Nn3/h+lkz
4Szl3jQ9QbO83qqk7WjcGq6hZFfYhaAT7gBBL5D0G98uB0muvtO6eJfN9nj9/sCh
2YAcIIupHilNeQ6tHsXnuOH2P4kWGTKICIcqv0kO8U9W2m6QDtbbHkRmCAQ4Jwq/
dEFLXel8yJ4fRV3gGO6xRdergqSnq62TmBG3QyVwGoqtdijP6lhNH6OxN1FkvS2z
D3X+zDcWAdFbmmShbcajSacEgSEnbPE7UUnMhcQ48IbRY5/G+oHNUClOrLPX470g
7Xt+dijKvMn0va60EoyVvSdt99Q4cy9L6BTGMSdwCkM9DEGIJZA3gF+KT6Hg+iZy
CK055rNEvjtI2qyyi1HoIhnO4wdiMX8MTuBKfjkAFJJBnh+5ZbKlYW1Gw3emXsjE
9I3LpPfmaUMVeUtR4vHCPg==
`protect END_PROTECTED
