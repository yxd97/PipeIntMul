`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UhRYzYYyJQfkht8RZRatkkL0GA0jbFJzaOJ9cNKfc8wyEpVbFBOBVUqLXwHYyj3G
DWyS8GuhMn2rXte2zGYRY+Us02V2QZeb6GgELJSUd0kCKX5ZXA/Qow6vC7KLCGMq
lNCe51S21hCs1ysrkG21f3R74/PnoVXOelax2ZBQkjZTQSX/mpCS7o4gNABgltN6
sbiSEmZuvOoJOk/wtAS7EqxRTS1GuYMR2zD53nVAL52ZZ4mMLQqVXBUwnjzQAV7+
xasT5i5rukGCDNBAwki7mhRbzQlS3790f+C0DywKSZX2awmEKq5x2h7mBd3PyEFg
JA+5iCPzTaEO46wtKuJ5WbsH/YAPsGmVJmXVVHieNGZ1sRdhi8BXQc50MInS1cye
OlL5KGQKp5FIHrrZFcU1Aq4VJyBGjAXTXy9XwQKEUdFV409WtVZYlEvF7q4B3naW
49EuNj47NpbZ4xyrttcbW24UUPkj5/OXM4x2220hUNz9+T+LFKlyWWIGJPDKcJqr
KKuwI4ihV7qxeu8uwYwCXowxNepjQSw0o+0NLaeAXF6NRMMoEOw07/skcs0gGQPM
m1fJkio+Ia+9iLe5LcTAHiFfchQKQ28jmP15ft/498VoDaXvsv+Ny1qro5Yo6sl0
XEwaeobY58P5R1PQyJKnYHoPIhgScI93DiTNG8KrQm6q0LBylAMGfxaCnLap7qQw
g6IFeJaQt9MB9H5JumFshPa3a56GzVmnmQ/4CJyuHrQKuyKzmXV8dUNzNGblgCrB
F5Ydnc+bDpvJ2KktXteeT1ByDThpUXk+KsQrybKhExbXPzL4NXv++OtPnv6Bd+W4
6k7t2Ba1DTZdEPh3IxKPwpkTiENqGDrMbbLWc8JhkZJZidUhnfUmLZ3w2B6MYnV5
o4KuZny9zrq8DyfXTnpM2wC5qtV78Jt64s3K1GpTBvi2d4GrA9ebKfAxXLSfenN3
0v+YNtxI3jZPWVlmGIrgfPc6Z4TyImY5exR/Zqp0SOTK0/oBLolpCH1K342foIhn
UbL9L82G8XImz1wfVFKHE2H9+B8W9C62SgAUeDD0mS0faWpehyLLCDnRb379HfsS
y9oBBajKbw7mltPScjn0HhNjTsL8CiGbcGxhSJiXwerwNJAIYW+07vbtUm4XCfAz
TqG7wHgNvDNvWo25+YX3WMD93HNRDFk/sd//QMAUrdCN96Z5rc3Ba9BFIisA5pAM
hKbtl78rkMPKIJWIAvxcDOvpwsgiOPj4PMvm0N3bOykQPwsa6sl4/qZsHtKpIwJ9
U88/HTo+Yi4fvXtTqQXyjBBxwvD8MBVVvWuZf/9e4/Obys88JsS8WkhuI4rl2thw
inQ0P/evj2b1a1GQMTo0nVTtoyR0EMyFpVW6Nt8MsrJNbn+tb+4zNGGEfIEsri3h
Q/GeWyzBtfCTWQMdYRr2Enu9KxgI5iCCy7JOUUz5LDJOxI+03XSmpc1vgnkAWk+/
rPid9ixCEV4nPQwcP7N5DnP9ZMnNnLZzI3hVfdqIMooG0ouTEb5fOZA7mkK/N8HG
r4DnUQ8QneJQK5Ws6R5+BaCG5nkn6dq3n1PwFds0/f1xJgZORNYYvGirg2ZN8Jgq
KsSHujP+gqnUx9EtTt+iZHL+LFq9ZAQw1OatDxHGdE6ycrfFEzbzSCb5/EcaKUpH
vKvp2Vv5mAxra2gRcqVCq4gK8dkezbpozmpSmbTTTLyA1y6M6OxlG6Q95ZMQhq6f
mMEp688Ck3ZUMw2pSbFS9TDEHE8WkOYqZVfhcjZEd1Yca+roPQz1QdZldPIjIwmA
8JU7CPFpPT+RdjEcscXeL7okAlcrryIkiKLD27DK3uanoy9kXby27xQzwxl0NoWs
BzkLQjBQxfPjlWpHI+5i0VHFwXGSbHcFAfqOakMFDdj/4Uk4vP4WM76EGmhshWrz
u+WsxmLzDispWU97NUoDyjzT4l6v+joC5xPZnWVvCwNOiBxFv9Mj3xRvehxJbTHz
hAZPh17nv02sqe+e8CZ2lnoCK/O1hHaW9ynqhRyFILV07AbAOlsxTPxZWWyvK8sF
O7mdp+NUnGpbcSbJRDqOj8dEdgI8Oiu+kda/IRtBYk9DarbL9I1VLXDpz7/7AlcL
KqmdGiFtXenMzkf15yQ6DsPLnhaqJVnsaMXrPxQh0x0trq4HAQ+0XISPtq2BPBJi
hhIqfd8tSb80BQlCUAs1DkUXZXRBw/qnyKi/BkCTIBYM6MPTUgeY2KE1dVDT1VD6
gnz5kODlxbRfb6wwoRXdjFg8LnbVW6r68qlvxeNCQPajPQF6WYsKNlC1u5RB8Nlf
6zis9eiFks5rMmUtWOzWSY05f1eTXlA4sNUnaMvyolHsZ5btCtP+I7GqpFtNF7cJ
dNIcebUqmQN0HSoOk4oJPUivH4TWit3vLJuRKKNWASkZXl1UrtY5X0DWMs1EDVxn
1y2GaQorTOfa73Ny5uCUG4WBpKBVe/1tADccexbGzpFtzYXjDrcdNcLmeyIUposG
Tjv23VMKBFaE5436+XRTuN3pD26ami5XDsS/8oKDzs3L46b/qfMh4tIvd3m2aUoT
brMNUzyMikZ/ti14Cp6189WSGfftS/bzFDrKpgkakJwOuJfmC325egThTcX7veAw
kG0zJZXrhfYZOM5kN4wQOqMSLvoEpJpK5ApKsZmhedJFtX1XzNm40KO8+4hvGpq0
`protect END_PROTECTED
