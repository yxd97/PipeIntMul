`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqJSXqrNisHJYt0BKEb6qKaNL8U29asO3ub0QBk+OibmbrUfU7D0dmidtPctL1iC
3F0ZSYZ5VyWhBYPqyhsgxhkLUgQRmvCnx7ybApIwWeYqA858GtWRCqYDqpEba5BL
UoEynN/LPOgVnfNAFThj5qGsj6ZRalAeeLrQVaTWyRE3NYN8aJyqRqIFzJ0az3JQ
B2utLNsk4Uic3GLrEg5opiMrqAsX2nxLAHZ7OxZBP5Ne3f4KBe60JyK2zpHl3aaI
owoGIm57hknm/XnDU7Y2uQ==
`protect END_PROTECTED
