`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mUZkIZOSmTdF9yjgnHHfPZWQmtcvXaT1roPzpaFRTe7xP4ms7J8xm3dXHX5i6DFt
Vr4bZa2WA2vb2txOYyF3QKvLp+gxlv50AlW+SCxnu8vYREp6dFPjWexkR8rRk6HX
SQaKGRH/Hek7ayts1entd8JuWd7WAkReQiPasCHvspgWps6wugiNSHs4He8N84vm
QZyrrFhlzltxfLKJdcW+1IMH6xPWQK0HOYmaRjIPYekKHj99zmp3zpa3FwqgdOl5
/bPAA8IAmzegZ6upmbb7hPOBVyLhQQqCK+g328QYS8s=
`protect END_PROTECTED
