`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+KFyO+rIVN8nQ3SRBjB09EoZz5NHUnJByfIB6HMlO7RHAkW4JZEWVpOW6Q25xAps
sWQtNMi3D9Dt7qJHN107IPFxgA1/X2quvrQ8K1G+2PnU/2ZabhdSot3OH7UA+HFr
aAN1nJjpWIIz9fNn4y0PqZCIoo7f8UZSLDI41OzhAQ5U9N8DYjGq0zX87KBUBtoj
4K7I6xDh/g+lB25+4bKy2iULPLqOtCzrb4OzrjAhwGb632FqdP1NR7ew8tmeHPRM
TqaVlQrhAX97Nn62bhXxnw==
`protect END_PROTECTED
