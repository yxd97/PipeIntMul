`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aY8AU6JoyQlZEIoQsZdVxT/ePlghEWQuKKgC7yKh2XpmpsqRfs2tSovrsLz57ZGN
ZGvZL+q+YxAT2a2dAyPpB2lmW//CX6HRLQo6ho45K0rrwbme14USDlGVbiWSKrvx
F/oz9+2NGxHaVTqNxTGqeMdbxT/qnl9L4G5c/F8uqQKPEwQnEKt96bJOFwN228vH
gwGlYYiwB3TFKiubC3Y1+yEIQcOBCXtb2BGN9uuQRQwUqzX9ORhfRSsn+PEIsRV3
pdbId9UQxvDlYbnnaFQe7zQCR0FOltWKy7omikLMkwCd5oDn5vUD0qv9BQUYL8T6
FIAOdxYNWLPSBkyMm81p7F8SsbsvZpe2Mx2lMM1Hk2vykdtRfWeH+Er0i/JyrzTm
9Ao2smnLC6u9qXW6lAWBXMPrg0U+DGbyzzLTYFCWbfr0kA55RnQ5Izx+FNyn7ytQ
MoN3E95xKgvncCHk/zdjHxwrvnBQK92qWUuAFCY22zX8F7mXQYFk9L41qjOA8H+S
ZwS6bcqZpzbIyJ/qMlh0t7FUxMzqK85g6rkNqp2VBxqTin7qzOu4VHHmWftdRY6m
PJp/UyymASA0/wI04Y+ujf9eWgs8RRenuA/1KOFfBeQvFNKsfCXr97T9IKDQ5udO
5kPdPmAAvktemmo6KmDkviLnjgoOtHBfH+rIxfJMa9p524dAOWn/uuxND1zntzTW
y4kYERl5ScckzREGalwLnOOGPmCwcl/10oG50LygcRzng06Hejo+VYAp4xYGioao
CUkpt12yiWcw0Vg/wrqILhPayA4yis/n9a3C5PYCTAw1WqkxV9/oZSMl4CsjqEZv
kk5wrOH7KD4JV9XjnvHlFC3EKpueNUchgSPsQoWFqodjzt0AvX1IRaYKL2Kpl3Rb
i32Isv6Dn9NOzofuTIxTk/lvFvFXL+TyzdqrxxnuVi3EfV8ZfK30BsATQp29Fn+b
7vsqDnvhsywy7AE5iH6IEH1MHcZoZlOjZdbi2k9HbdOa3LTC0mcjOuSJG3Q+uXaE
J+Jt59bI+TmJnrBnHQ++WP/8/0X2D1S54/FCk9s7deHMhdAq9RwB1WZSdkAvCP8M
CUuwgrkHkwxDW1ovWt9j6emadag4XVpAbkepk/mXe8soi9LA49tYymFClyzmihm4
X/BlQP/A4jsvRxTJ2X5MYPzM7Gp9IPdCOM4TWK8VU8mIgjzJOlse+VKGFd3aOtm+
apFHTDQBS+mwf2ZF+xFEGsFMX8H1DjhlmUNuRoc0vNEsULgedG4la2611fhxQFp0
MHh86XCvbPpY8p+qTLZAraOSkzkA8d8U9d5mghd4mvcTrN80A9owCS/N6QS7RUkk
JRkH2DOgjU4Yz9YqAjd1BIZVrKcBJGEeWaoUz9LsVNpwVXFLf0a8/vXMJyCtgyIj
Gs3L32+FaWqNuZzeWpWLKzYDEFTpaoIduEPDqZckn36EnQLtF2TbIfO00LZ0xw7E
X83lHIOK0OCV6rcepvW2589s5bMmZTwRf4U6kUcxb/DLAp3YGzcbHVwHca4kco7b
hREHygn+3aEKZfMbJSi8ZC2oodzvGdfa27NLlE6H9NhN9ApeTXLcHYmd3etusM0O
TagMKfMlqXpxnQBe2b0aDmgslr5Dtg+d+YTEDiILuYTGm/4Bg3fRR15BG0EjI5Jo
URvcRjyNn0K60+6av4/UlQYGM85PEytjKSAPCuUBVR+4EgjTR59+n/GdI4pl6LeX
7GYL9Rj+7JFBY6EDloFCZKzQIc7hEh8xE70/Wsv+h3DbDeqkI2VWQIO3VsEeHosO
yNqcI2kBPRz69rIGzsFArg0gxhz3IKkEooJ5rCjBuskhpR50x62BzCYJdjjCfkfS
a2hSnp9ljJog/lLj9P85JGztqH+6JMsS+b1zz3zGHSks8AtsS1Y/GezyJsDmyXe0
P219B+jFt7+MH12dgaoa2OxXUp8YUAnuTEMSpM6fdfboPoFd23RLiV6ZrZGcdqrm
hVTkzEdxY6LCMtV0h0swM4ClglN7tetc9by28Ceb+6mBRUX677GKyGBBGgJdTYn6
/1B+0JcVF2SU1sM5j0XECzDsI8EICjAwi28L+Yn60jfsYQxiL+nTUL3pRBJ2kp0M
P/cC/IGBabtRiu+aKGQas1INFB4cE/34F64jwNwEnNJbXNXzQ8ruZofrpqAXymi7
eOJalFBodsxhlK4bxj0eUKWxp4LEvbQkDaqjcB8jwIe3R8ucSqMaDzsKSnLfMpJj
7+WLFRn5NpWVujuDiFjMST9NPC8pMgXfX00gVxs3c/+4LCiPMzfpqMn65QYX1SnY
r3ruLPUwjPQGMs49WjQHZcY4Up2eCRNLG2viRdmffbf7KQU/d44FUMeHx3RTY8bN
5KM34XbOoZpDzTV8f/otl6ktCAtQA/4ttLkZHPGhCysXi5imSpSPwTMO+AxTzQQQ
yVru8j/aaZaYGpZLzTCZBtas7Y+wc+aPBchT/feC8CdMe/O2uZxaylOLazHkeZZ2
TT3NlJhsDwm7HG9uz6O0oX8TJS8iXIzMVQORG9zlm9gHtx1pE9u2+Ivaoo9nsuGW
XcWtHmg+k01M+OADnfZeChiM78l03SRvtov8zZbM214ffVvPA7ZBc1JrO7RhYIOj
Sqr3AdoHzCRrHq0+iyYrZikqx2uG7bl+iOnEZVCfo0TkVDwvSZ7lyTovcX1C3GSZ
ukUtex4B52K0OlKRNUAiXQz5YsX2NKNTr3XSpoB9qF4TEvJzGtW4BdsPJbXChgWT
O5ALMqh7lG01RlH8aHvMBUIlobheX73/I2FzCDSho3Ks0SarHkKHFA4FwXNY8c9a
hAozSHeZGu1gLvtnb86qGq2fLvXSfEi82QfY9ZiK9AicCSYoZFNADRW+vN9N5UsK
SPIzB3J1CalycJ9XKBmDI2ga1k6QNicydsKDZG59J0qrJjbPUrl7b6oDym1fihvs
tJ0M19uwzJkEqVTkeGC76mu5y/aZiFQg1dnquVg4NJVh0TJPGpHWlRt7orC0H6QP
jCoXtk9uP4Okls2NJvYPUHsne9MURV3SomNI/C9a2d+faISW8ZCVUJxSqOxsVDdB
tb1qXlWklRXrO0shddJYOyGegli/Ms5DDqbBD5mbFcew5/zQHYWLnuoChjG3RCZ4
Hx7PR8Z2CG0UFtTRwvG2sbOyvUgJi+TD5wjp1+S7gmAlue2SP747+yyrPtiZcPBv
8OrAkCqYAPJVHHI75iWWBjUWvkbFNmnxFeR1h91tYkrcTZIBMfGQAg2XPEM/OQ23
hAmX6RTyDXkZxfBNt1yNjiTlYiiZHpHNgRxhTDQ9QqbcD4sE54/68CyVwaXauJQL
6/VFwCJizM5hRmruV9Z5nGw+hYveVTFN7Ayd74eKGJLYWtqdfbAg9BdH77yo12OR
fXiiKnL4jyD2uqqewzXY5Fje+xWcFLez1LE1K5xEKapHZeZoQJqbJV7b1pePNc31
FZ8HzuJfuF0vXo7nL44oue73oWp1+kwP+xa8n2026p9C4cdR5rNdo+qti/u7CT04
5OGkAxUpG7kpPjaL0E6pzztvPhAC8d7uE3jWgWlIwZ/gnNeYtoOAjab1g4yUYKX0
yYxNa6tC6QDDXiVE+2a4kcMYtk7lRwmzz6PCc3cdM1kpR8amTj+mhDnZkLVEtDDi
SP5kgWmIn/TH3OqAcBZpNTGYjuQEsq8tob6/ociSXReM8ZlM1Pr34SiAFG71vvom
/ZBW2nDRcSQvLsqDDMZLNS+yOSTy+Yr+fcMA687M9p8XoHpqNKnWdYFiCXd/LSl/
N1Gsqn9/HFlfg3uZptyZkFuvkikW0TAkIPsdOsIZA2NNimlfKJxXmKrd/Pn5AdlE
cZWuUORicWBkZhXxJSeMTHeq6bApp5U0ghrZoSO6jBb3KksQuwqO7oRIYngZARw9
TQ1ILuRAb0486SwlY6YDwwLaR3iA6zfQPkHk7kknrEk9RtsZurvFPzpT2VSNq6dn
AEIQbYWo14pzrHynzpCEWfWCR/VN6IW6S02Z0mqBZ9n+dcZi9Qkw0chFY8WSToBS
7/3QapVPH4rxfdcZe9BielOcD+TlUnuEKGeX2G3zEl+x1sJTDDO7ssMrxmT3cR7X
nbDTAUA+qsddXZA5BkCAQmiuE3yRGRbRhBTrV9/zEfzLsns+bpRT4Z9uXDRUoNJl
`protect END_PROTECTED
