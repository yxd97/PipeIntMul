`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSmmlJ+ROPLL8XbsKrWwuFLwbMe+oXNXPa9pgeYRbsaSm9N/BYqCOQKK83UXZY/5
4nG7Bn2x1E5KjjylJk6tCQo9fnj4VShiOKLdRiF++7dr0RGyiRwSZISsnMAHQ4mG
CpYgVEE7fSwp0H3KUHTr3CHi2WdWl211NSHYmhlTTdFXXNTlw39YuNTlpCk5JcHZ
zppWTwv7QlJfq8zw9y+19+WclF4YJB2h2UISp8wgNdgh7BCtkNYcKKaEJUBTqRxA
qBAZoo4eqC7dtVFlnYzHFLuFtKt4p21ske6FfYK9AbziquLVg7hFXxC2sQYYoIv6
ShQb/cgWXQ2GgbVTW+b64T9TBqTErsrkmjnIBsCnYND6wjuZj2YEOh7XtpBey3I6
zgZIgpvoPNksEFfaBczCsCsWd+sHFBv9Mcu+Rjn7B7TtVBaU8k4HO/jps0NoEVlH
`protect END_PROTECTED
