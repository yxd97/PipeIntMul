`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lzSvsAyM+ADvXIAGUQ6CdaXoEz9ecgSB1RhRewVGuHTkvtnPobvJmJJLF6Cjwjus
ZlvspOMudFtybIpkLwKo221OToygg0SBH5D8glvCvjUg3GBg8qP44pp9QTFs9LTq
9Fvm/0Rkx/R+SbE+zqlQLnVAxGUDjNTlrgayf3n/l2yGRwRG5hKQsXlwpmzeFA7T
tQs4Fjpe3bO6BLlEo2ZkAViLPqInXYNKW/h4aPhAfeUlsJCa80bsF1qVneygzg6c
lCfy5+qmxvwAKy3/vDkQsjthnwsHGRfRogLc8Ft/lRbn16OJ3ZpzndkKbtewnc1i
Mq2eYRZGC6dbXb8DXki9xSC/rpz9L8JvgsIXZ/ko5KOARjz1CGWFShw6hFtlHu9r
bRiQsRMW9k0kshtGsw8qvRTV16DaNxtH7sFkWdLytYNxUJYJYZjOMO0/7P7m4DF7
u7FxYxjYapkig6AK85sTJd236ulNz0BSzyIcxda4aPxFXnQoeQ5UovIioJyU8m9j
tl6eeSdj/8mPpOcdS66O8aJ5nwmvYahUr6MkHtZLN5vhoJO8dOKhzIbsbRkukCKn
TlfptKZo1Avm3dDLTPh0dmIr/vfjhp8rHYkEeSzKXA0=
`protect END_PROTECTED
