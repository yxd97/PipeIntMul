`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzMWlYRV/ANprtvB68lkBsXZ8CTCAP81QhcQaMuZaSzp0NXgzKOaWloaPdOo76w1
UBaNZn6mhtkl3BHJE721mblYSBXv8s7QFT17SFH9W4C7Wq4yc9C30l8ttjBto75g
6H+bqbOF9jBt+N2GMaJXXuI/2zG7G3UpzNm8Xe1N/dnsYzrdo8OjP7T1XQUyXtnp
UDQ6OhevOGdeIKDpn29skRjv+ircZMlg9HcByyKvNZ833pGhIPDvs3E4D818QqXO
dQrAmemlYjHKOxbJCxVXUALj9BwLkkRr6Bm1bTlyLxv4i9MHO1oOvOlz2d8CLSt/
4NreoGaqIE/QIqgVzz9/ueN79pHTep449LT7cACfheqsruDnqtcTUfx5cHRmkWuK
XypimFYFq0+jKkBldsBWnXX1IKHDrmrN9PxiG2ph7GiNwf8av/VmIKW2e+fSa308
`protect END_PROTECTED
