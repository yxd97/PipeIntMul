`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uwKDFqeLAAx+T4NOIPrYPyNZoJQDYYPOlbDAQy4Q8UXHCUKBAfNnB4XUBdn/QxFR
WLjm5njeY3rI7ZgDWtqCqWM1C3JOkBHCI5wRzrYCZ+sMOuGKgyNHxVz9JhHM27yt
aAfo53YzEH20IcN8XBEVJhQ57Im2kuW9UaAmnJ5c2nm8rb/6mavlQ+RRQuNQxC0U
Z4CpWvegW/7oEAfIhpBBwhYjeTnMmI6dfqaSTTq4n1mDBd3Wm9Ne2AQOtHMJFIxZ
6XBFZ+SyNzCH8VRoCbMdmxfsjUwvfK7fwx7eAQABhBOlQRj/YpfwFmGHeNF+sKY/
aLeXqjFz6bWyw/GNt+dE6d+DmE+b504rWwdd2kfQlVI1xfYWVVc8klwd+oJ7jNrW
JW6BfBBryz9uGO/FpQDQI7+DOKyJ9Qwk27nfbuDBaAqXKkG6WKNGi1bjlHg5Y0qr
nA5dZ9E0z0+r3fnkLlzzCXEkQYFID/kul6bXyn8EyTncBQy7A7Kbx/s0PxtL2+nJ
bgQlQ4bW73H1zhdYV7QBqfeei7GDWNXqLq7rYjAsHP9xASP9tZ0RrC69eyQIUIPT
0/e8fSWciYxAJTRIE9GFqo0GFKXaVuOSMVDA+ifcIBRSEgI1d+uHNvWLexWxVWIn
Sfji3aUj20xOCZQyfK45LcDfZX9mDakKRvnnJHU+4s2xpqVMBtA5/snapb/QxuNc
b6ythe3NSL6HDAcY9TEx35eMs5OG5DGnU/7zx6KMEoY5dwbqk9Q7sIHuHljNh2bb
K4IKWf088wxw/M7Pcp9UjUBwTYlfBEY7MEghafSU75qHiQN6SFrgOeeSn2Spsq18
lDxjJMPmMDskp+86usau7/q9hLCT5jIosMpYHn/Hil6TvRYtiXgUvyYCdObE22PT
/oDi8I/SndkmvpdlumRTCzKQzkPqjBMxUrNAeiIp09N5OR3cDOARjkTN9eWi8KOp
NQmOS1ICVPy6UR2QtHmBtmacKbEIC6fAqBx8kk+bfhgX/EJ6S9tlBdb781SzwyLb
N7hZlF43r+l1LOd55QiU1jS42kl1m3OihuVCsK75loNSm0lGMZnqVmsAhURv+/Sd
pw+l9eBAZ1kUCnZZm6D4GS1WQ5ctJbWGksfgLTBo4U2W4NQyJ2wV7W0xlcwaApnt
Yfx5szgQ/NVQEofS8LN4pS2owW58LA4FcR2S13Jq3gUt2nKSZPBei8TrhLro7ELm
Leqlt8TIqMbqdzcjFxWkq2pSMlmH+shD/dh3mIR0YkWoxHa0Ms+FfwXMvKyjlCPN
wcNDKVnTvaeCh40Qq/G9lXjOULtXRXfi8DMj2rmRoLAmd28oZZxffes4UPPjx/Ne
Ret1AHDu4XWS4VcPRS3qAtprSpKzGspBxh+8uiR5qUg6fU3pBr2kFJ3cpgNfh651
FilUkaPDbvMYv4WY1I2OKe2oLw+AdrTmbFOu2gZTAprqXNoCa80flVlE/24H0lIR
1ahZSubGYHq+lPJB8nJt/B1MK4rOAbu+w1N/dkFJKj8aprULk+3qNxteS6CpnRmG
pH0fQvu3bbFcKgwQJ9dMa+pLu8/w8dxxWD7eAGdcRk8siyDbV6tu7n23BNmSvaei
54lPB5fiKGo8klBRgE2MhNxHe2XeRghrbzx/SnaSYjODkAKqzDYbwtCDZJOohAsq
MRJPpaibOvXxIaQ7gJReTT3+jFeNCJZwEvVVVg+RCpxNVdrRc7wUhQD8dO/TbB48
8rMaWj+21Nlap2btyD4dAnNRGBEnGAOE5Z1yr1dn7eQNmZz0fy8K7vZFIwQuU3vZ
071CnVMc/7aC/yHW4JZ9Vhtlwn+VJnoWFV4uY2z4WtaEao/wQeLxDau2+ljQCXHK
xADM7qrv2t4Ke5IAPUNd1+68FRseiPvjulpjs1hLEDvLrVGl9ERObCj3nolwoTkV
fd8RFnax46b/d7+eydF+fL5YxrD0XCINhJQa1kyE0O8t0K3WAdmpzltO/+g8oocq
`protect END_PROTECTED
