`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eAPg6SiObfO+da6Bh+qg6qqkstQ3V5svmCQs+S1b7DYAJIZImGB/m75PyA0L7jTw
8J0Ci4w9+V92c24jyLsU2ZT52ik2G7zFzFxsXdVvBoonrgW33mZ+QcNYhZMYmG0P
s+H+ogHHAPieIqQIAgSsjKW9Y9PM/EDBDYH2JoWKG2QTxS0XyQImzE3ZNjqZkeWj
2Cha4ehPKTnLX8d7jWMKxOo0gqyuQdLFX9Pr5DtN5PSRcuyCHlEpNmz4J8cbCM8I
lHy3YfiOAXm7XJqr78m77PQGn0LuYwreGpdTIvre0INwIfpK4j7Cy0+yt1boAVQM
P1tdBsznhRy4LYIHckRb9hLRGceEsTgEkBWkcXD1N/Qhj69aRUAcmhRH/G0lgO1X
BAWGW6GUFXC25dQGqLlIzH5iv2GMmWXD+CVZ0CioyovCkxbcRZlSNkpMfNYllXjz
KXeItAkmNDoCEU25t2XM0hDj0Nta8bVCtuMgWcmyuXLeAMn3fBWg6MRI7IZdT5q5
lojoKEFrCc4s0g6tsUaUpbN4nh1fAUwfNlImGidWkTUBF8QYWBMEjQ6G0YtGa2iv
y6ovq8/3q0VhlGZK4mRbraXBPhv1q/IsrV0gXETH7Uiidaq4mvknsqZ6ihlQVrRL
zL5tqGn5gjKIJoSDKV8SBWEBUMKxoH75Vs81DXusX0Sk23RM4YjlnQ817Kg9Ssv7
UwaOl7+iC77MSznd8x321lRT105U+jCM20fDaPh4XIxfTHryVw5pcc2phMdZDHt6
1h0CFV1sKt/rWvClp3XuIWGa4nIO825L1z4bkSW4P1wq7D+EMrgO8EYEaCExPxWL
+ibOOl94RSUqn+zm53/TXu/uKdiDH3rLT37aO/0D/PjRCoajRkmWApFLEwKD0IDB
Ogj5XSIhKBDtoeu+VynAhgDKbz8bR0f85Dgx69pYzqOMrUXTLqVgCqRJJaPb9p64
5qI3pBeOeYtlTWvrFe9XQa9mhORByzP8k6ZT+8cd0UruXZwPdXWja9e/uqZsWQqt
xitfWuvKc8kZaKS2f0YiSNRUVNYyM00KtUrEN+E7eD6XJpmaeI6hGtNNB7VQ/msG
njtZrBOxX9pOf9S+hpzQRusVRh3PGevqYtzCMBa9X1pPtQ6NeSSDScUUTd44AUPF
syDka6LQAlnguwM/URcL3pTxAILq6lSKimKnfmAo7od9nHyOQXH1jNGZRrkLqAZa
AVFeGqmMY2aO+KzjMIYDreQk5V1NTByRXiqJIOIBo2FxOz4ltXrBatWKcDf4lja7
RqEvzK+6ebXMFjK4VBV20G6UeYpue4fksE335VUNSYIEwzbZ9M6YYxGQGUMl9BFR
A7osOjjaz/RUKUQrKkhLZcdr3XuFMITtGcXHuB5iav8cZ4JjTeSyZxKqj/ZIirl1
/kvsj/WZUc9D0avcAw00GiUoDxf9OB7pi1cfuQgyHaFEIHF5qcCghZYT580sRuGK
Q/EP58s5LYW7rynRkxxBmm+zwTl1WqBv/uAO88Ba+p6OqFfWOo1NxssaViW3Se5O
35HdzdUb2oDtCqrmCe0HGg==
`protect END_PROTECTED
