`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BIZ6QTbEvUsMzhlTdQv+ddLBaQnrPs93vJnjD2fnTAxvDgWd9Jku8eZO4bjyWvW
DabcmS7/0QBB8O/mhj3iSadv47wqkkfRoblJWXbmMWJgYb0fgFgdJSsgfirjjybc
Gge9aIYI1YIOzMhCy/sWCEG0d+ZqF6g4akO/lWaddI71GTpkgCg70EEDxU+iqPP4
PHGB4bbGz2OxcvFfBfcJsrFB2sDN1iA51HC9mttecYSzc0JyApRwyECFe5VON6kd
sKZmp9HY5vyvH4M8/tq6nB33xZqzrooD4VTVzUV72U9P3y1/zp4XSORyeFhj2oz3
fuCSsU01CNXKGU1qJ1O7cPkiLjfvsi1qD3M/3gq7D2WzRzQx1u7+kr7mC+EXRs+f
+7H7AFJqndq4voT07bjRKPTf12Ne9IBhuX+l1ytT/2VsWN6fLqf4mfAHCHEQRovc
X26P3W7n9u5uzhZHy4mg3MpPumaCvptuzWKpsXknupOpOAl1DiWfvl0lwK5/VfEV
gCf96ZyFU0IV6ux8Q919b0UjWphBf6YooOQ6IVV2eO2uxxviYukIGYsfo4B4qj7W
wwY/TzmQEx06XRFDyYEtEVPvsL4y5R2JuO6GSQR9cyV/j+Vt6RNeMVsgR/hi2Jfc
YUVN30ZMKf4ktaNiPeiwvnMD7M807be1/dyoCpgijGomIibiPRbvloCly2ZMZzo+
ynHErZnFbfs0ue7AnOySKvfOF3mImc/c7b3qIs8eBpUpKN0WzNtrCuOMqjiFjnPM
oenZh7wEvO1pfYmuzRKV1Z8v3zGLIwHwekbsufBMWex+Z5jJzkG6X/otFlNTpZpM
h/RfGUgIT5GvPx5HNCjUNrD/7r/PhgHlXiUWBn9cwpUMwYh4E0N23n6IWMjyVbuG
KYp0ou7+x+QdWGG9UUrNhbbXCqyVQIxiH8kmwQqjg2Ibvx+ehdgPZ1f6O659kZ1k
8Zc3/neRKJRcia1mKduaWH/cgHOkvoFP7KnLhNKmZisL5xwz42CkWARS2cNKlvNP
3IUADw18mY2RXZ7fMK2+nJCnRgZQZy8IaxsokPFCfgfWFOIHYork+3exgjTqFJnT
MHJCXGbQBuANo0Rmw/EcMg2RcDJHaEpu5jw6vWETIh01KYgiBUt4o03FeulpeKGR
4aSzEPgvY051YNWrIsvAXUUxesJQCm5xJcgSQrNF95FZdp0l4JW/nntwL+tKWEYH
ZbO+z3eJ4HHa6/kPzAes40UpWLBegHQL+I2eImvmUtqOYY2QKAMQDMH6SdRWJG7W
FaaKV6mjMPrPEMqBDjlFnJIS/V0xRZQPC2ozfr1iZdWyIXnlUd1XDyQmx3/ZSS9k
P5XqQMLTrHsn+JpES0PDzjPT95K2BKMhwdBEIMLXcnPL5M1bAi2FmF9anqxxb9hT
THMQcJxD1K2SuqZ75jjuUJ5/jZqYBKb/NjTVx6DWF1kWCyPbrkEIDPAkhqUX4K9I
eWzjFzlrG9yayF8RSbGwbd256p0EBVaK9RsFGRbP5aXjOTyDuiaqRTE0qep2+DH3
k/wVS2fL9HHfyhYLZ+dVHOK1Dve7fTNFunxSSx3O484rlQ8mXMvtFT31yMHEuZr3
onoPgZra8BcKTSLMNnPnUaVKPz5WwggWPhKi6aknfm+5N3vno4wdMYcXB5SaSjU0
ZeTTPtY7W90Cf9qJMM7sjkE7YALCOtDzIppe88m7bBhpVnGyjDqtY1N4tkiC7twI
PeKCq+9nKDPwiJVpIGeQffIW2wzjeFdT1y0+Wz90C9U8EXM9RiiaiA3gRFhtWZSS
orhmfq/fBM0PPpQolvFSifcG4JUafbNYKLa8DAdT/vuUtEYa2I/Za8WvVROBjTvn
CRHpD8R2mEylsP/6zlTj8UIKGYsget9zuKak6o7BwWuEsnpbLRFkrPAxWJVIqHju
OQnwjZ2Tvd5/N2JmYJ/zLsuFVzr6T7gKYhonZQdxtkI0NlhiOEREs9ltTOM3t8Bb
fMMN8YbjqQ2veroEySGDBykzPK3XIruvangoNyBttoKrCBOGVXBaF9RnD7fmSVnF
uODwoRXO7sr29UKjFas+Gi0FWmGP2lx5xFpXzViPp1CslHIE95/C9chP9XS5GXXr
Ss9IV48fMQA7jjhCCaErVYjftDmqFfJUPooo95gy0acnL13fYLbRSuotwo9Tr8Yx
7Z/oiQHwZ+AMHj0bsVELudaj2gvwGl2WejRQsU+XinWDuNjgtzwhr4G76AJSzKdz
8vO0tJxaLysub/B2WoBmKiwlAiLXz0Em3rJOypLtlNY3PlHDu6dgZ5s788rFs0o7
Ms1EHFaaqYfx+5iji6TwIDYQJB3UQAvP1mFQTgRxAXAWDsYcYQLd8+pqQpW9FmtJ
3ULEZwPXRSCwRgfYZa0cRc5EF+caPH+Ho3Ip67o/gjLiXyG5lMBIY0BFZyhaVuvR
DhIvhE6DMl53PQFgxA0cQZyNrYXeb7qZ0cc1pa6Pp6nKqOKkzasuUA/zA5MuB11i
FJ4Zix8RE5BTvHSBU7r0iAXD2KjrocwZ5+Q5OFdnsMm6dl112rwBaNVo4jMo+i33
81tv3X3XCnR0eyTDc7iCbC0dVwKsl4PIzXPPXpB/DhNezLYkOkBf+2OCxGraQ9FP
IU6iALtdG2pkdmVazoDeWC12jZTZo5vqpY1zdFhS/BtmT3QH7JQ2rds/04/BwhtC
Sr2W3ijZEB0EJnw1ff4ILFrd1beylmzR9IIAoVTwC6vya9+kBSEjfBYM0MGUDBqE
RGAHLj9LbWqGGynvXsHp21QgRwshkTYcEG7JJfuKcCHdYg+4uoN4aLEs5HhSvIs/
WvMZMjMog9igMkVWXVD3wmbECZ8Be5tYsg1uxyP2YYG/TkgTcuU1cKCRHsc+THGi
SqGeVvUAzVra23X3Nbk4DaJM05uaZbSojim1cReqfj/BhHxCB+T02eKT7LsRmre2
BEMFtshYtOXcXoBJ8qFx9cU4ojAD2f7GNpCqc+PfQHWiXcBtjQ7f9e3rnE+lK3g9
regTOhUrnNKoQxaNS+E06LvsSdjxKvQzTpGIC2xgF+8pOZZCG6vYVvCXApRy2S0u
sNY0+IucNL6OQiNrpiHBqjrQcmMBwwzrB1DQpJo/lpNaGd/S7pCy4I3rHpyShl7t
R2UqHjBVTKWZt3GJMbcssym7h1FFuU5NT++3tQv8UAsKn8MvDL1YnfWD4xKVP9Lv
g3IvIF5WNIb+3zzWZoCgbbhBRlLifD/nC8dM5us9mZ4sZAuwVkvdsupPEYsydzBF
2rD+DMgiPJ6o/67Gt/BBy0+36wSA277dtOcSo0JVWButp0I3RY5u0YQe7uc2t/e7
qc6EE3avnQwa5GWblNyB5gfVfi1RhiqC0IY1UUNJMpA709b6cH65CyHhTRPMs0Gn
S1AV5CPQSIrGwyDRmxKuE9ZVTEzNn5Tyrpj1nFvf/Wd/b1fH4ilL8jWhnhmaaGDO
KSLe5DWBCkC2q+UHetMWB278cd/Xmw6bImm9rMEsIYc9m0BZLSgmf3STKMJQTcip
+d0U4xiqWueBktpACIbXdGRpEOQij9BH0+3gaBMCY3Bh7nm5A28xhqVXkM3JxQAR
mKvXrsGXd/L635s1HlIbNF7GWUcjz6XUuxeGb4O8nurflj47aWwGxnqrgQuPYVtL
ZmxtOktkyTxOVNOIFGBanKKRiYWKYRZ1Yp3t9dVD7LwKGR+qyEwtpMH69xF6cTea
eE61tYfNAoPMdqQvmYJlSsmWA0Ybd/Wn3NZtcnQxWVeXJCnWEiMyR3vJsmBp8sP0
yItYVKa0DGYYsTS1abZR7OQb1nYKHkNaeMyi1fl0rYUa+CwtH64/i+9D5lGDVa2C
qDFnpkHzpJ2Mo8hJkH8dlZcLcJqq4ukwvB2Ihjb38F4wP0wO0LQkIVRB5+PwWCI2
hsgAJFP9Yd/OS3JK9DzGZi20fidkVHdJgLyE5p+zowzPsKRZynzH2UG9clbUXrC6
fcBAi9taWI8KrKi37DAKHMN+6L4KPCnV24z4db2WUbiHNW/8dwwZ1eeptf7QeQai
i3CoVOsHdyKekouc/IIfpkJt1KVXq2VPc+dClMXm4PGTbD52boXqHT2C7d6ONNSK
M1F7O9rzAkNAC5jfQ/e1wzFn6Xb2OY1xinzIbylNy6ujMFQvJiyA0J5ZZ1rWrmLX
lV1XFNNfAuW7l8ZwB8WVFP1Z+KOIMEQQSTPENSfrVx9Wv9yoH8DrBDH4/deNkgeG
XyXXMqxHeUXlQil2tR5KK4K4CrMS19KmAgRXlaqLzUxnCrXZOMdaFavf5ScfOalV
6VtQIZwJ6YEbxlZpf0JU+3nDJce6qDkEa3UGH1dnkaT4cT+FecwpwMl0d7uSWRNv
83RoyNkvQPQzU7BfaBNsbDOa2ke26DmyQ8LxYFVNZhyhP7gaRt3hYYUpM3GXvnD4
1G6RggFHRuJWPw0M/sss6TtZZYg0X7QGmJ20v64bipg=
`protect END_PROTECTED
