`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RM0MyLAhOdOmUqlK6JS0Miz3FFiLEZyw6vPbPIdV8jRdudtk0vSYdGd7mZw4x59c
nDUYvZgFbCwF89ddgpJxkH8yqAAWGPfPTsgMERDbtucanj5XuupZvCImfMckOblb
lLBQ7Dc1z/tmrrqtc/Ds8OI16xbIU+f4ognk7QjMMqUOeBWiwJt7gk9zxvMtfK4C
HC106Zn+KPQKbyD1BpGr1qg33ctRyLYCtNCq+dZVsyv0/UDQWWS18SEx1FQJBw3h
QZu8EjCL1W0gyuQ4GTquOtx+p9gTiwppNdPTvmrS4Lk8n/Mw40nB24r22LAKMyaW
KPzbvviM5rlo8ClB3Rhrc4DtH/kx9SgyMyG6M2RqmGIwtoNyXhjZWf227gYClRLN
mjg8VImfzY7rJWY3R32zXXxuLHQ7RzwH5sS/rJYikvf9CWxt4yNfh9nwHtEwxt91
S50ZCTIJ3GuAS/zbvVQ+Mm7b9hQvMoXnZuTixryw30QlaNyy+/NIz3Z2agsFgBH1
Pyms0fq91pMdRvJK5XH9jku/z2pO2d4aHdOlJFxb/ic=
`protect END_PROTECTED
