`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DT6sYtym7SoCg/KEDiNyWQyetEu+PLNF6vfGvCYu1WvGxydQeJvCgF9Z2BZCO1EN
gMv019O/G8I5LKoag3i1m86A9vJ+uEbBDPss25QegetTCtDOSaJyURRs1iaq++jS
Iv1oRYmqRl+2FMXSBAsdRQan7NzESmbbCG4kniREWkfJlrges2rw/Ne43wQXnMGQ
9jsDX+HhCsXo7o8loGWxfFaCJNE8/Qwqlux6i861vuV9v2+MgbuLsETwUUmaIhVk
MWuJSWCnrLmukmCZ0qzvDzMUzIgJc0qIJNNqbev6/ugurYkExs79OHzbyj5FnQfB
EL7RIVZIvStyjzg9wjkyFf0FHlIEEA8z8jh3XErm1FyGYTFZk4Sq+xwOfGHVmbrA
6ky06IDW5UFOWX0Q3+2gYIviQ+0jAGCBxZFxnFm/Jrs=
`protect END_PROTECTED
