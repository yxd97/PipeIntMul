`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DG0fGasbH3PKMCFOxEyEqU3CrbpZdSASqNUMAUHzQWh1fEHLYJe/d+FvZa4n8uRc
YlLHjsG4kH+693UwF1Nb3J2by3vnCBoMAXrdlAr+0gQsg9PjtC+eVomm8xfTSV1R
YEnV1LvaiXyEvvHlU1KkJRPmYDanVUB/N1vBQQTbcfr6r8oStB1c4bE0l3ZIWFWC
GcUyP5/ruBCCUdJvi0JU1uSu5ySqSn3mWpLPJ034OUBpS6qgIkosn5yDNMgPi64V
vV53LLYZAcG5cfbawT9JnE+RrjT1s9oBpkvlUWPNAVE1hyd8MOzJI+7/9eRbb1zt
rInsbRzAH0Tkn5Hm9Rdm52qF7d42V0ziiuHHJmcp19/Bu3rUDx9jTanD29EMvg7a
8apklpoE93TjUpAujCF2sHe/uODbBNUjGQKh06a/nll/QY7BHUaHuyNMnvxJke+z
ai5xfS6OMMsoHgpZYdnZl/qKjFRIAt+Dx5a0L2iZYbHtGXgWcW8O+iIPE5IMHyf/
oTc0UP1hnlkH60zEw+dlr/Y8j4fAXZ/pg4i002AsUZ5AWTo+c9S6msiSsq5v46sR
LpEXEmQCS6KftVGBKRBcRg==
`protect END_PROTECTED
