`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BaJkXFbuhmXWF1qjlGL1wtqlzW/fu2MjDhgZzd8t2Xm6fjrqmKPqPyz9q5H4wW6
rJqScnW2RpA78s7zOWJ6fuAeHhvjUx8XAsL9uX5+zvxMvGt6DMpVagE1Yz8t3jGv
ohhx0ypY/JxWGZhSHb0mDUdHcwtoVokC8ejmS70AImSSrMszwLYf0fibFjC8Nnam
zYKfYXehTHAU/s+X2i75TfpTCRmhWAvRJQ1o3MEGJuiIgUZzVbhTD8loVotIaJor
tXXAizJwEh9Nsp51rOAChe3K6vd7XBSIs6P8EAFR4rHBJSZOnjb5WFKHLoCKi+nC
Zhsk7681mzvV9Az27yve/PupOM/fL87wMaWyWXf/zJw3Z6qDD+E2mbAgqyEWmsxu
`protect END_PROTECTED
