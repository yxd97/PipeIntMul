`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mqCruHzSEabflageCdtvrq3jlLaAUa+5B47cIwfnQbjA131rtquF4pRr0muB49ds
+BpgT+6e+kcwIB68ZBy01kYvqV/DiYajucpmz1x8T8GssBoHNNeW7g68BYxvSQTt
YNbt8B544herQA9YbFDpjv9sKLwsGWD+kXnYGvxpZKXlebkHgR92jBkiJx6XfEWv
ZbfdiTGSKkQwl2acZnuYKe/ixvpb95x/nbY+N4Uovbf7hLBWId7PfTWQiJ5cl1Yz
PUWwMdvn3uTXdInw4Ipd2kuillS5hV/0ccQm/o/l5dlK8En0VSmXezJ/Tz+CvFDO
Pvxe91+YaXjRbekOPEWsP3pYeTqgHKUPZlP5cPfNTlxKJdfJJQIq1k2dqcbRXzFp
tiOHtdvQAokKLDpdXL58HCQOAQT3q0u+JYENI9O05hZL7i/QzX27lTihH5RDW43u
6KtD6ccZgzt/d7dvDBuf0FDVSLvz5TS1MzwjM4Z/nYT04n49mglxMzCrPbZ6UsZB
hug8/nZaGZnuOfrD4Iz1YJRgwb1cg7LNAJzonONdG9A30Uwh/P5xccw34xtSSlhv
Qh+mifZruD69CzZMWO5+qsO+w1+5rLL6VBsd75pjziWZSson5gjkLO+Hlv14Yvq8
ogEMyFY6u+GJGnaCtdbIvw==
`protect END_PROTECTED
