`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yaiUZ1z0WEVKWetDd3DYqyzcXiaRu0/8Zk9dNYD1v1sd6Z9Xxl8sZH7fpbGTofud
CMiKDJcwIm1fnGm8kIDDSh+5Fenvjvs6YHfVCqHZFo5ksQOvS34mSuKbxbJjIIWh
mUCHeNeBfaolxL4gMlpieDHHw0LCRZLpssXPLg3exOORVU7lfvKWs5ggdTP96npv
baJG9WiCiF5cQk0y6YgwXH4n9Qp0lyiT+3GM9FxSgOxCQ0vPfvbunCE00kl4ELAO
te2z+KBm2/oQxj5BleQRcj6becCDdWr230tg9fnkOIh5sI3Vc3FNXP9PAiY3hOiU
nRRi66oEGeTzpO30ReoOJcageSwKXCdlCgFYUpb+0JgjKRgy5zLTbZn55bZqdbQq
FKtfv6WyebOauBuuUrGfsyDE/oCQLDRaLwBRuBXuVpjFY2B/welE/C/clqSxOKEB
l2IL2xqTQNAu/UH8htHGWGoKY9ofrd02Y/n1307qzPZGXk9FcCgm8h5CMOWh5HT+
2BJUKjWxGxpZKZVGu3YnZ/p9ws1rGOhjwWjlNhWBGCCji1ajrjIDW/kOU5SLNxU4
SjJJ4Sj5RkNyPmgdeqB/NIO1vwR+fiq/ajp6uo/Ag4QLUhA11D/5M+GMxQ2Z71aR
d6CGK0hRrWikjm/Jktp74+IcOTDpW6GPfaU4XoYjbWTKhNSEJsBkeh2KD9gw1vz/
LqfKxoKJDTUkhphXkwH3Ghhq9XTVlRrAOV+PNWFNsKmtWHr9X8jq0x56Uc3IJz99
vaaL+quEzPu4yN67D7aCEIIFQa6wzl5Cdnly0ywZG0x3au5EepboPOEpBHJ3Keuw
Sax08Cn20rb7WHlTUkrIUmQha8v/dUJ/2c49+wX66dKJNQ/8BoF8m57HCrnJvPbB
tGkEhVs5pdChtxXYylXKH5Fi9cVDt6NnrWnwUH4COzyNlBh9dFnJxYA3WgFWimBT
K8dHkEzOvydTemIwpjguuSjnRgMcxaeE6TOWCqwykqEbUYadNC4tL5MiqmmB+a3N
fyZlKqTvOI4UfpGL+lW/T/2QJdGhdDOjDvEzVYqrW5z1FQTXTgdtbUBv/PnOFyxO
hVkmO3XtJrZ958bqv0SsPh/9ZWbMXBZuSa3dnoSBiRXsxecIoue/PCS/dGE2VRQm
JmQ6yTYuIPbPjn6jwzMC3ViCAaJvWs58HtSinigkj0/P25yeJ6BBJJW6uRd+BtWz
ce1nJJZcZyov0tT2+RxYoZsmZGeQNSfwZXk8np6QXZFSWl6km2FOo/F51lMyvO0e
9S7MbvvfxazSQFUj0hUxKYhWoPsz9utTOqDi9uE/JQoN96yVGfbYP9UcIIZr7DaM
rSwnqBqXkU7gE1CIsiRzDUaMAco46ZoGr4BwETHQk90kS+8JZRVavl4nyyWTHNAU
kncNLjs+7IJBJfDGibAOx4eGOAicTM6YcNZcyu1TZe+y7JJYY09umZxQaVkElJRR
G48l2/OfC8BS3GwczpHKV1q8PMoF/PTEj0rK6rhYGNMXHgKrxr5j1naQJ0iV2GYw
tErbTRCCXqpkzQy51yU/8xmIktIJFbXGNiXUtoHfO9BzPQNcQVRr/a8VHb8U2uL7
keo+dVkcajLfZy5rVEEGbybKKwEAcyMjex2NhTMYahfU8XcmtQtv62lo80U4E8pj
UpKXU2IaDhYYy+LA6TBUdsXmWn/eADKJNNn7wZZzPoWf2cJ6uZg1MBNBlufw1WDU
RBYM2Ybur+zvUnQcBF51euKh63P/g4BfQnMWa282QtLQbXLgHXBBu+MSkZ1j4hAE
+wNabmKc2LnkVnufkO+pzeNh4Di0rnqhcF25QFQwGex6NPRYIy3EnAiuXOD2E+CQ
m2lOj5yLSXK3x3b0mk+ymHDROm25cDXz7a9T5k+p+dwBA0Eidtu/qsm6wo0wSERK
gpCG0Vz6u5nJn75/JeSwF9IrBdelWDMgemz+nE0gj1gMDdl5BgqbsLUnoZZ20z09
ss7fByjbIVns7HR2roBJm/OPIhfD3k9z2ILVJNm2an6Hl2VSJ5ArL0VEVq8KoKwP
r8Eg4gJ2MM4vWJUHMp0TT63pWJ19R6rtqKdqdJ2l62byrLm4mTBNXBJ95BzPAVVb
URddQunJNWe3reVQi+NYkSAwDC8yg+Zf6q2+cKQtNRl8d8+PJIvfhN/t1Rjmo2XD
SmcA4VJekN6T7J81OSg3Bp3yLHt+X3hssTGHrMEuqIWg5NSubJxuFuuaYPRnkoBY
WhSc/ZpwKWywb+jbeEIMQZdeuMaYHyD6sazt30VuGtqbXREmnWP6AV/JNAALXzda
Mqgv3NAIuflM5sIAagc9hcwCEMDA+vtahJhhrt+2As74dgJ015j+pJXx+nygAysr
KBGxm/hsfNl2kr76ed3FCy8OGNb4UuIjbR0dMD+y8880qPaXaTFW5fKweQl7EdPG
gm0PFsRe95xQLOWe3IWBOk/pnO4Q7K1nE83vjY/0bCZLrYLJpjgeNbEd6xfNwEvc
rxIX9GqxF/8CqmDpTv815HziuWMrzzVQOgjTtRonEynTfHWX2zv7AkC96CYMN3C7
//4mQKsh2MDl+UZ/zWmmGU2u8KQcoLjBx6e0r3m4gd0q9h6DGnYT4w7CQq084QUA
4TbF9qC3xGdVbYfltH3BNbjpeYY4IQ4kOJKBlepJEAfv7iMGQ1cBebBpptbWHImQ
p99eDl9UxcLVRKXIs7fmU3CSqIU1q1xPA4eeL0uhJR6k+Phjf9e9TMJtoIIPupZ1
H6s7VcH7L6ULrbqgi2s8Y9VPl+UwiLikmYeFFVnf21hMoOC35Jcx3PS4YllhAxMH
y34X6DNc8Miu56hw88HIVbpM/AvA/tlBQQlVrYktsMpOoA9ka3QLYroCpklbMC8J
r9ZwsPgtPOgHGaE4+ayOawABLUuZpgJLzkPZGJR4eXyTv+JrVIhTpFt7QHgd6bc7
`protect END_PROTECTED
