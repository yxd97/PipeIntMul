`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6efymILiljZ8Fc02lS8vVTyTBmMwHBdOfDAXDWucL7Mh2Y6hO/zb95d/c2HuqQJE
k9rWL2uB/5wGxyg7ojHLFVoe8nK5HohyDiB84F/xCoXek/7mh5MykUIkm63ewx53
9vcFqzpTiQLOqDXfLpjLRFRsSHMWiJz2+uIejGDZObbGep2WHnvBCveFbM28Dp1J
fb5koR5koNgTAKgza32/QtJ8b/Q7q7rEllMsHbxIvF4p8FOS9M2r6dFP8FlnjZYu
9Il2LI+ZoMZJOTbS5f7avIX426syTXpN4V3EW6oM95pZJwwB+zImvWN356jy/Bf1
coeV1Alf+hPbsgR2e9MAgCOUHr1yO9E8/Fl1zExTUTpYECUUXgeGyRD+y+kTXufQ
V1LnfCbG2s86mREzcpuagWSW6SMvxxqRIV6Il/+wCgk=
`protect END_PROTECTED
