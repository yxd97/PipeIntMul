`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GMs4xzk7CRb9IcsQn9B05qx4WFIChrUhX1NVOyRhI2T4i7c8ncyTv2e/JrehHQtT
lJiPM0n4P91DOk6kAeha3JlGQbImAy0YkKGgdy3YtZNefRqaTBBr6zYiSfizixx7
e2clCKbkcuK9+xE2Q3IC3lzIKyJhl2xEvHhpCldba5LXiVV9KMnH2SiKUdVrZ1sW
Wcj3JKWN+ZPKmukojwhabFU1xwVwHIqh9eH+1xgjiLlOhs33E6jjwl3i+b5Y/Y6M
QsidTlfwOE+20OFT3EvRQA==
`protect END_PROTECTED
