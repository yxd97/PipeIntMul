`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HmcFfRnI/0RPFNTr4ubYSQuqo5tFLqAgD/HUY1ByuwtHOhSENEhAsSeOBYIldGBA
rusrP8AjxVMpaBRyRlBfUue1tcICdAiD6YD9qMz2EXR4HoMbFTqhQb0V83Fyzrht
1QnoRvEAgRtOpVk8R0kcx6JeVTbbhgGdA0x+zbshCsCO+0/3w2jspfPw2SZhglMG
4sB+uTTbraBi1mlGjtxOJN2aoLrj083bcpkbG1dBcSfshnXdalfuUAnTHCME9yiz
9wPZckuJf+5JUzlOxmCTKw==
`protect END_PROTECTED
