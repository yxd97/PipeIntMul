`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
54YQQcWSVGqIRilUvH5h9To2yVNW/ULVlFHLSkDQV3XB1eTJaX5ptgl6vR3gHRVM
4qddEjUufZ4MI3oor17/hcmsyyJhJGbxY6jt+45Ucpt6P1X+VZ6uwm3zPgYmXoYY
5J/SeNRuxSmgT3wkhKOhlpsGudj2VztyJo4HtlIt5sDJcGC8ogE2cOfX0GmmAIev
lKWKHJZciKGFGdxg08vk11bBHeMCue70DIOROtDDelZhCOpvJ6wph7tE/fGiddHq
IZ+ho1HA1v0hTDa4UZe4DIg3aaxABcfGUfrrcC+0T5icdh66cgTHbc7kbP/nx390
APncrD+JJuP2z11VB0OJt4zWMfnFCPvWaKSXpKCUMGVbWVUaTeNfjS7Ok21ZQX1l
8xp4IfHBp0Me2zJAUmDQOw==
`protect END_PROTECTED
