`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sgQ6PFoGalZwD3BoovqRfhJ9kynQJMc4m7M51XbpamcC2Fc2qr3gABaEUNHFTWow
6bLXSrQ5+GsuVxGgmGXv4Q6sh6ujOf1XJuBZl39lKkcNG+CoxfvX17cF+3V5bzMk
496d06VK9VOVrzjSpceUELZHythYIM1ynIWxSItbts9/LqFW+KaESL4fOOBf2cJj
MdAtgxjcH0EoG+bWyiqdoxmms+fMJKp4bMBIEyMK916i8Eun5fcUXQ10oZhZOoLb
4uI4wtts/mFRIf53ESp+kY7SEm56xR/6JMedSbUziV0mHuvVZPGOTPZNPcWjl6Rx
EkiQR5vL9A223hrphdtZ2L+yKza42n2I7Blx9HHqhNWyTuilhNglR4ldliym8Aug
kMMhOuh1kxFtBd22lpu0RnQ2vXKnYEh71TJlt9ynQ3yqT2EZS0LQgXcitz0CkT4N
7bAH3zPAx8uXJAhkS5hdp7wtnoemRs8K2nkVcCQYjXoLxpt80wm1ie9duahKGVB1
T0ml1OXb4E1bROEPhdt2tTS642QDmQL2b1fPUoF6JvdYdfBJ7T2gynPjSRHg/ikV
r51LmGuQYk7OwhFyP5NJq4M45K+VXvzGhQfPrrVjAYwO1SkJit7k5YHTKoR6rjkq
104INIsaNGzV1rno7EbeGFKc8+5xvXKmFnXnY5xkNhIlFVEG2Ejejp87e0s6gqfs
IYBWcXAnEe8C0RYUSML9MZT2bqWFa4Evy+8UfIyD9MROnWXa/QYHnTQp9V0Tb/IJ
`protect END_PROTECTED
