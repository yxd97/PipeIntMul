`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzPpx+WESMn2I/DWKlxFYSivuWo6DrAGdIl/P90j81hcC/DuukrgOJsJ7flFa6d/
ogTbYgZCXHuHMxnN7v5IuR2kW96dj4OfDdaB7M8wsigoGELhvGDB/H6D1heILLFJ
YJPQimIqbJGxb7cNiTefpEVmk3BG+Gct9+GeNBZH6qEEdYVmjX5nWhyc9/6hkBHq
rDEnES1MbnrOL+YaI6hmTqf4JNf7xZU+32Pf1DgNgvsKjXaf3sluKGJ8xWqxmGrg
68PQ8m2odqlU71GbCQu4YA==
`protect END_PROTECTED
