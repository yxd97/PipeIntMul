`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvANQXm72De4aVPSJr4hQ61zsSOJuONb2J32sbFXBe5U6WVBWot8GCxN1UBwHB59
BJAPz/02KH4tLqVjxWtUyNMApZfDgIDumy0V9zaIpg4iLk0KoSB6D2dkwUtGqjmZ
rZRWTW1sAKeKsqPLIHy475lndl/ZnN0v76T98wGl1Hol+YdApXYlUTeYwp+ld04D
am7nc/7cCzKLa4ZU0piUourulEARyAy4XcEsKvT12ONaUTBSKrZv5DCI42nlCKL7
VUHwafh3rZgGvTUrqUUBSvG2d1G6ptdoBzP9elaHD/tWWIrLBYuH7irDmIQ7+tZl
HkLP7FA6aCj64HGuPgSH8bAx4HtMXnvEKIO/6BAtPxuUACrhhDe+uanRlCcGLBD+
kjXNU0XNwqjrA1lKhwxTXrV2Ues31bEirs5Ta3nI+hJvikiaJEqZHRKQ0o0lih33
`protect END_PROTECTED
