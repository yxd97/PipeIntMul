`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S44zSY8BAS29E9VkunZFPZQjnT8O5KEHxyB574snXmXuwnYYmPLUx6VawUEfeaUe
MSpvJV7GI0//xUphASAUkRV/Tv+9esXBssY32ZnIOE+ltwPZ4n6wGb0hbfthq3No
PrboaS48wZMqrp/p3Y/wcfHGHOh/lo7FVs9ZJzNAz8bwcOLPDxTx0q5/gCKlm4mc
xx05W+BxcyzVPKJAQ1pPyZ46SYFheEfBPHLJIcnOFl0B7oSO/5RQgbP7o0wc2kHw
dTQUNhe+i9H0MLClmqK7MoqPYAgTIbXuyOaI4Y/2Pji/47g6uX9Wm0gWQHPp4oUR
EKO8pqTFx8dir2/QxGuMJwOZzXC3njYmSBVjJjXSTxmyQlNbP+x5kfzWeXkrpKW2
QrdEnPzCPCojfZRl5X6I/6/Z/npL63hyFJ8hDFjPFI1+LY1KtfI8LRw2+RfIOYWj
j/E2fyDKD+a6moO84ugTvCnL7mMOWr1jRJVgbhNRf80=
`protect END_PROTECTED
