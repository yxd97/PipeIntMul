`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KirbWHPYeo5L0EXvgJnP3UqtyPsU8yqMzTgyggOG30a/MXl9Z0cD2W1OtB9ieBNE
+xgBAhauHV7OHC9FBBhmrw3hQrCF8YuFTNlbB4XCBbMJT6WqR8MZtFko8wo+JLAK
RZJAXMlF6rgubIIxRzWcVLgMP8TkZBU0ie7Z66XojBZqYGY6wuxQzvZQbUKG+y4o
wod49BsiSnjlTuh8sT2GHJUyt0ZDsYuX1HVVBgWWjMS+vQBLoexhKAr+dvBpPQiw
A10uK4pRUUUb0fVukzDWasZd/TIzZOe0gyDtMdM+W8hlDAAUTHAKj96Mz5E9EGF5
KuoMA2WZLCgoFJrD1RtUP0acP4mjM7w3agrguMkDA5bgR1m7BoyZmjvPyuS9dKDZ
B6rfKhYyAmDVPl6zIzL0FB7AMPU7xBg84ddH7lR+9FHkelAQNxQQ90FH1lAv0CoD
ErMsspGj5kwyRDGZft1FXIUUlEmgI0foRjLMY4qzNojcOcjusSikzDH3gl5iMTQ9
r5cUWEizFASIOxqbGOuVK5brHD1tHvjShyOjVsKXWXNKEumaXaZAEsL10WVfGtyY
UAU60Wqdh92vBlUVbeF3TG5Oi6Cd9sQbwrN0Qpz59aqXKNHxy5XuxGGV5qXWD4zX
N9XeFlcSe5kV+yGriDbCBX4uDmM2ztBkpQAoUEDSeBNVafqqod67iwyBvbn9O1iS
ssF717Gb731ao9ryaHIpMJdMepIqRxZymZgkr+cq4ybLwQh/xxvswJOWetQag9Tt
Gzsrn5vChpvLF+Pzq5F0jdHZxwlvet1JseA2961AUqWmQ12XKgoArfeMDPeA9mZj
PuD11iANAq0NNhP3+wfGpKbGlT3IsTNJlyXkJ+3XFz08uBfDfrbDicsNgtknJzMs
oVW2o6MoyEscLvlpN4oarmy0IcwHHicEZgm8wzJP+QUL4S+sDxgAwRZ8jaF8YtEv
u0XVSAKHTlt2JDVQxVs4a3Uo+t7+/EVS6M+1kmcL1N3Tst/y01+aEhatGeZPbG/A
CiV+Px+DroBeyJjJEC9JjWjLLkyJgy1daFZAwx4DsBE1fTzAQH7zdMP74My5zCXw
PVK2RWuargQg6HczpDzm5DqMyzJqrCPLPPSsFftrnucLO+IT96AnNv4SEyrquaXC
nkycOiRaBkZeUkHZTfAi79LGYzBe1iRysGEEB3eHak3LjEGYBBO7IvmfZs76nPPq
`protect END_PROTECTED
