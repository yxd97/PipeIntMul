`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WIeEIbbqvE992L+n8FLFZvDytDARshOsKh/kxGJE3fO3DBRu/Uo/qpFjhmCVe9j4
sZaOjTR9MLcl7zmgQM0mCm0HchUlLD2EYbdap/PGO4ZE+mh7OdDe87jyueRbwy9h
SZ7o7PORosWK4mYGp5IC8CijIr8FTjsvP7ilJRBSNfQsOzI2VqUrrf8fCJG1ItWK
vnHyKFpeiLmSLBIrbChxI5GGchLLtwlRRVX0MqMmJpM3ycweOOEGr5A55fPlZH2V
0N2dZJtmsPkU+S2IOKocrhsJ9w3H4HDeqWvBpX7T28C4oAcnTZ5+clFOVyal/iqk
e0ThP4fW4KPVP8jmn2q7cut/gbFSLhhBngIsLKuJHQGtOnitReEfZtdhE9LZvktg
8JQPfp6+kIRuUY2yX6jJGvKkcnyeLaGm/om6rhCrzJCiCYtIlX/kn5sF2oa4iCAp
jd9kulAxYBkwBjaM3UZ2X0x/b9Kt/aHJkvusBOVNU9fFsoTZUUOqEKLZRBMj32JZ
5wFfWGKGvKn9fFOPwHSgSnYLa6kqxa5haEugVXYCShVKA0m8ODw5buOWpiUypvrO
WgH0Emig3moX0lbglVAovbDRlHU6KpomxaD5LiyYwAd1GMKpp9MetpltaqVdVNaj
8gRnMxipefJw9SR2XsSmUuj3g26N/9Gnc9jHi3nPxENrm0rIbm/2d6A8DLBLMdyR
BZjrMLN2PdsZ3UkTEEwsC/uLy9/VbgZ6YpYtc3Be5J78+CcYipatV9ciL1wmxwov
etKBLqK/+8rz5+sUyu252GFadJOtH2CmTwAz8L9LJTqrRkqqnxr73MJ9lpUQT2nJ
qlM4eV+eV2ytNDP7IcEC6oHsoNJFY/vIWl0KBu9Kxrx4p+L/Nt5B+RJTV9O6LZH2
sn8Nv7xrsyC1i8kn4TrNE6enVHo59cU+bFb7Ymr3P7qAyanhMF724br+kA+cDkX6
GzyujFMQ9OPNcEm46bDY71oLZ/YA+KJFgl/AfvWbiOnZeS1d+TFiwYNIqMUu/Fyg
sCE+lypToFckJz3ejPydvuo1eM9aTvzwkZFm4HKrEvig5dBuflpP5ObMLX96DV4P
gxUehnEvwDgfYPhJPhtUodAH3pclFLrXA/gmaLyR0jDILZhgPxUim6M4mVyD2zJr
uSHowPrbuzsw+c4OuZYP/wBQyeUajyKdElMr2ulBg7VN5XwZrpQmo8BbE118OY/a
O2xmiiFqCuZpboy/i38B93Fq3v2b8OMU4PG61Oq400z+YchaWef5nyE+1jYvfBGz
mcJVI56PFgUcsWWGjBi34faZDFS0LZp/ZieiXXVedpLaN7rgQwAstPRCk1XfS7u2
dUlfejXiryZS9RQ4kb5qIYkvVK8JdME/+QASP2gROJ81WM0sad4gNxNHBdyK7g5j
jDGFx54XE48ZY3Q5HtXxtda/tXk/3yLiTvQGB1w0czGezFqhXBjl7k2kcl1IX0mP
oyQRipt7N8rxfy6SWD4elMUEm9fFQwA3JBTqrbxiO7hvmzm41NvLbViPBxy3xtfR
jgfBd1ykazO7Q30kVtJjmccTdPLQ9ua7DYu5jYMrh0Jl/clettaF4ETgFRasIg9z
tYf3P4hBf0ZvrKyeHIn867diZrgH3vjdCkfgjkTHqebgqMfJqGJAj9zfL7509pcF
BeDSxapciyo1HpsnYhLBQRCGT4tQWgo2LPgvmCNcylnQx1LrS9p/NJS6KPBjceW4
2B9XXZPDFdF0AQwXLwx2AU+v+djGV/LXsuKHtXYx1XP7GYy7aE3Wg7xqp85LmTcf
2iVx6N7RNm+pmctKr1X1bDRf7CTvbbtKbCoQ/jaiGRYwtagXbuOGm59twCCrjGTR
N0xk5QXZXa2L+/+HdYZtkoB/6aIDASF0vENve27ldJjhj6E79UQRwYP2t1gmYBwm
0DtI1jZyi7bebhZCDwpYNCh7GTKs2jH5+R9epSIjkUrj7THkXN0NIGoXUrY+3ioq
jmqUVnKmSRXBdEeU19oqqAtqQ8fIRnw+t8Dj+rlckUlgxohxKhGMEeIRH/4+sYob
uP5gftKsv0NkRIuCfa3lHUQ6tOY1Ldt3XA2TFn8Q+21RFLyVq8jupGNK2wQ49j7w
tIhXnMCZhtzpOnlYNoomAlTYjfgVXE/bmqyVRu6gPcN4okN9aFWTrk9V/1pLCgDV
b/PqWS+ONPRfHRpG3mRZ4RfM+k8iP4cJg1CiczAEZr5cHeXv60nv3d3E6KxwR99s
uQTXs1Ly+ZpNDaXxglnsq8WjhG5WYEc2XI33w+vRO5gUhXZrQzBWpF05sesgPU5w
jJK1/r0x42Qaw+PwOY/aTX2AwwV9D8Ks8QhN27B+u77fwuh3LpOD7AzGQgD1dR7W
NyiX0wRJw2wngrczjLS1tmmSu50yOGR6lNF3bhlqURknFpyq6nJf6qSLkrJfTTJ9
+jRfgMSz+VKrTpO/EzbfTzavoH+06cEbqP3behHUWhNxr2iBMa6tVRlct18Evs+G
BEjOfKmyb9MpjcyhsXk1sZmr7FU0Jvtv1LhVbk+bzmpj1gQeteDdGM1fK/AG1Vjk
JvES1DVxA+TSNE7x/nx2T59CcwyW7IGvttjPCW5k6SZ5RkITo9pgq0X6ogABZWLs
cGnVvEsVt0EzHIYIBlVQbX3NuYUeSbvPvTbJCN+zw0pjKNId9CXNt8ucOCMPDDMd
jPfoDMwP6yyMhqf0MMTTyLHp2ekYoVeOzqwOmWloFZwNIhxjPAvo51jAVLRFN8ux
+ttCfjwn3axJWukShQEZRU6clkQvani7So7QF0YHL6b7qfTAIo7VXPm76J7JOj/4
0VDgHir2RoqzaayFHsWiiDGls43nD20OPsp66IPUgp3tm89M5diJeRmWWtobFWqe
zSIHeREV26AvDhqxqj8YMxG7ouf/5lFzheGewfQnm0DbfyuChr0qd8SWkPtYK8e1
EwchLMO0vCUyyavRviYzkAAN4uKRR0NBSSzlC4YE8/Vjg/kgGJL4rXfSKrDzv/wT
n4OXN/aw7KE6ojGE5sdISP059ESP+AWZhn1+cxa2xJ9OqlWzKwjDmvvOdi+SLUS+
QkhK/Ml96n05lah1xFg57KxKH+MDR+OVKRuSxw+6hqq09Q6P8RVLamoFSdt6/rsJ
GIV21+XRqxuB3lXztkuzAPLqTxTl8pKCuQe0jwuu6IfXRtRuI02CjcUfMELI9GfR
zRE3pCt7SoJkCy13R/OfwWSGwbnUYZUp7joTvivPrcFZQWywI9F0MwX0Gck2ipPe
y87BjrjPhh0qmMeHVc9M236WUXt2EiOVJ9MERrbh2SXsEFKMA/53y36PRsP/5JLt
UBBvRNK8g7ELRa9I05Beenn7NoXs0AgxqFRUj5Qa2PCqyTuXqPrZo/SXjAbvpt23
LeTajBEf3QiqZigAYNEQNn5/0nUj6uvMfdy7Ua1ELx0jSBSrqG+HTyL1kxPVZ9mX
tS3vZMPcTter6fI0p32ibJr1NY2Op0abIUrL/YM8O3t+RhcsYv6EUjh/myUmevRL
IvyD54gJt1anb7vW+b+/Nkqg86UQZ57fdyfWCpHnyC68bTWfSE4VXR1QP3g37VZA
jyR3r2nDADUFrzmbnEr6k+zgJnV8+4ZQH6nhbinWAkTohFGUXCNZuvVbVqPREPyH
un46GIJOD2UmqiV2ZV8ExgJMsFDy2bmkh702LEn8+VinyeueIqOON0ulBB04WgW9
ElvvzBs207nA7YueqXxN7/8kVvV7TQ0lmmlq2nR7UoxQlh5jmth86JftTX0iNd4w
dy6tYv1zJY7Pa+rM96B0geW6sC4FqfuJqXIGtd7uF0JeyDnNdlDsIb04SoA0LKgy
VSSTErNLKxt3ayevo14Yt77hCyGA3EEmDNhu7QBl78UW+KvFOHzVw/N+zPXPu+9D
a6qLbqPjR+M+Gg5irJb/Lo3Ow1/FSSLwLIzLGIYKcPiPi47RRR8V2c8qz95Yx48n
yEsaWpW34OC+NzctHRJTL5gE/WWwR6MGnjop/cc06NrkSHUtj8qH/lm7ZTORQeWX
V79Eo/83wEp+wO5WaWStks+6O6sXmSePvAJyT2WIOki/jgjCtNpddU4t/qrS9MnF
GDnS3cEQbahb0veoUBVQ3uHpZQr+wnVw5pcJFXdHB01spNkN7gfpwSJGLAHnZfIP
x+wknYZr3x/tkQpx8eIi41FaBuYnTinwqzkA14+FfGOXKfQE4oJP16wXiSiTgIle
Csw9kivPym/5vZkm0UTE3vXb6Jtgr6mB0ZBC31JyPT+0eTb20Q3M2Wog0xuC6cmw
lZWsj39AnbynSKP/PkSClLjYfPNIz9Vno4Z9zCgID0+67V2Mi+WablK+xk5OsAtx
KnKVlklSSKq9q+5AM0Sq1KKI+8hpedld36+6+Zmw/qfB8pJh8zw+hmIupDeVDxdg
4dE4PT/aUpMh9cplrrbPnxg3uE0hScvtqZRxRW2C66WSLKu7C9Qy5O6leVfC9krh
5yDK3W6Sp/nI8vzMKf2/VNXMy85zV4hFEJwAq4Du1RyYWo78Uh9bYBHCEib0j2b/
3YZn6Rat/m6srcWuoMQPM25IQFNspFIn5DydEbAxZxBAgQvTCB+7J9Mg4iD/cwke
UZjQuSd+ebI5oCFzRlkZB7Z2KUnZ4ioPrDPAyMoPU0PsHORFi0NHDnWFFSPp2Bl/
JTuckxvLEOe6uJ5RYlRli+YEivOPircaW7bgpzM5ZyEQSOhJeBTN6vC8G01AkwXi
ng9ON4t+vHnlstvwcS+V3H+P8mjE2FPNetGDEglWizTiTSeRehdBmPQPFfbndFd/
vHm2+9/SsfP1I4ZsNrEByBLiSo36kD+p7614X5U40rPBOdjxhJFxgT8KTLAXMKcT
Yknl/kgvnmloHkn0FD/NnrXvo10UFkCuJLL4ksofa4/oEgFWsDxaf6ohG6U1biyp
iJSm/sFLpbDynfJyhr6trzzUksDs97FLgcs0dJhETP8POeI32zPmL3tBk4ke5EZt
NeVyNIM/SJUpSCN4alq4psg/NtuYvvq1eNWzTGdcdaa2dclquAPh1JbF5MX0VJil
z0gIXr0TG/8uHaA36ublFnM8muRoz1IELt+8EhfX9cE3uH7lMZHcOJcxhlvR5Eh/
VXD0GCsrz2AfQOieVh1ObIv9ofP4ad0j3xaTau2272aY7oTT9LkoLOzY7BXqDTCL
tc6e1z6NlMqTw1HoRgWGErHwYV8HbWxYT/vATk9//6EmB0+Vp/Jjp/LNv+l4Drh+
QFvfGqfnx9Q4ORA4996PkS46VkvrtbApyuQApPJi+4mp835LMkGhQ8MUccimYuWY
vBUWWIEFgulAJ7FBOJ/jlJl9sdkImoHWKr5/MxF9NY5u6ad4sDpOPsW4jZaMBFv0
fN4P79CY6IQ+IpbnugDZC4i6sMGww2BO2vWb3koQmlVdsD1ONZ1ijERkrgznWJwD
zsodqhj8UwcPjsleU+XgJuI7Lcdf7epueCF2iOJf0FlML7tl/3/SLgrwA3f1V08A
PY8Xie0TAGFNlh545VY+LbOi2mJ1lroZFjcO+L9HPSf5qiyTK30vLiYspJh7tYo7
WBHwkgVgPNFIXWfSGiDiP2rDS59c9ycbwM7wIVe0rTtE1vXlOVvln+8ECarRLKeB
z2pm5QxT0kzAGzgD+mkH3aODMYsHlQHVg44rUv8eMLKo2ITiAUmfKXJfE5EoY8Ax
pyJwwM0ZRoa3tL7udL8soQpuP2jwr8IoEn4X/JsK60HiOJKmqKSZH+ItVq8ORZmv
p6KJ5mp6HX+zC4bx+kTkrAvttMuh1xYqaheGCbR+XTG2xO0Lufrk3voEZwAmvRTu
RLY9LS9k7Lv2a/a+G+FFsDBKjS7VI1kppckYoBJTpROUBhQ38/sty7sk7XccCX/3
wePkjeROFHbC5mVx8oj/LtThujF3KhFGwnwwZ0OVzn94z0O09qZ27cfIgwGhCHZ7
4FTcWL9TVAR6RKwNpP5g0tiqDrJOGZDvnLaNBgRvdqxo3/q8quk9SMO9tMKubLkR
omuct1FKM0PpB0ZVV8/DPTI2Zkyn9eqQf2p6EPwvZDXsxJhKElh34IIPSFkb+Ee0
d7qiwfewg7biLkGcZxHeM+hxEVZM833bJ1XujW6Erftlo/33159Y02MsUkIPpyPe
gurZ2AMNhc1m4Tc5qV2VDQJUsVR9SVSvQqr4jAw4BoS6LnvQcAr+wNqTjD2pIr/5
HAyGfqCS1DO4y6g8T2JF9Ac3dUV5XCnV/0h9hgc7wPvfDMByahukslKXqXGeN127
HtrhC0Hyv9hwVVbLcN2S8GdZiBVGUpJfFf6rx7Ob5gWVTlYmbLUZZd9OcA6ak9zQ
Ubq7bSvfvnCukPJXI1ttOo/eWAtwfZmXeobXRAg/svaWp3+Hf9LymxOmTIPwRz2n
ULmutghFUJVCXvbuGYVahyX1LbQdxyPsuyW/t/Mm8Mil1GUMXZAgwi+nWkw39s+N
ImVsIENrVbZAB8+XpzsJFMDANLlmV8jkVHEp2dgpw41wxZLBuQKad7QjhmZ7X2Fj
TBAKguOrPq/lYGomfOEAB2b7kWdl9cwKdhovOTcfA0rFPL/2gJupXg7laD9Z0XFT
VLf3iOBM3gV4IC4FvVcAPfiP1rvwsoPRYPchWjiZDHHRR2QUPaVXbqOmUDzC/+4Y
RXgYOjkE+Tr7AecVAzj0nSc6NNzJkaUsVX6V5hzy8UzZI9IC7k+p5DreYpw7Sb4Y
xAGEE1OPzUDfmI3in08iIxe8XXxBlm+tnCe3aEbYtMU1tL4+BitqKfqMVCqreVbQ
JQ97zjORIF2wVkFETscfWh5yK+8TR0mw/eYPtguSroj/IHVovDUZnsQFx4d8YTMP
X/SvXJmdliWkHoj7YpVwWPG+NmJLSerrNE+TfaHvbCWihUcImcNMy8QPLt3htytO
G4XUSFe5Zl19EadrzeRGqGNaHhCXjmLNPTLg30X09Dy68LiTTmV2jFy0Sp/bybD0
f0P09aNOlciiaWoAN7VKR07yv0enSTdQTdgPTBVxtIyqkMjI8zgwpOCIgi3Ax+Id
y/Rnpz0sqh1O1ILt/pNpMssTJLIHXN/02I5kT8yU02sJBZ3t4cfBGvawwVGP46Mi
tPgZ7whiA0xzYAz8RIWbMRNK8Pp2HKUx8xPw+GPqRy3xogZ58WiQsZlODGq+xPxo
o1p5ZIwV0YmHkVU9+7YLlF0ImgB685TcHc9LloH4FYGB0Ze6SN2WvbdNXpR21gTQ
mHTZBEiXJ6Fnih6kGgwqLeCa0zibXBu8FSiQ0ARWJsvrEQhZElUoMLLQxGTK1uZ9
kA6r1mo56+IFc54OyyQTjgPTp1fhcsbDJmP3VrY11Z17gUT6UvS0Wi/0GNZyZHNd
+cqPEkD4rvsBglfOpSeR3OPfG4gUdBwZclY+wML2GuTvhJ89dvbJjQ3feiGvbBL2
DBp+9UFs/k2/uymk74Dgwx+mS7xtqBrdOIwo/VCR2O20Il1z5Shlhja8NXKbtBdw
r3z/oIJ0JH41Z0dXjZLt1GPMQ8ab23d1WXh+4l4k2x8BXVfE4C5D7NXuIlIr2DQP
Bu0Iy00JFcc+GQgVNmT25804fD+2pbbainbPPxtAnDb7sFNntj/GKH5yM0exrp5E
rZMN9zJ534n3GizgTEH+N38Js4mzECRlOO2+f3qqpSNq1yedtN6kW6I1J3ggN/y+
hiXp/tUBBeAyS+H5z9YXGjkVGfj3pcU/JN3BgEpWthzmXvI6jHqCrFtaSrH0Hb2b
nbsQCR1bCNRfYH6GaEpYsDf9C6z6jbdJA2EXIbzkrumtWIVghge5KtAm699UsPse
4pJbGBQy18joHqDWyqwn9JydUBkkrUUbO6cUjbafQ3AhIH8Q53m9EMAuJBv5HkMu
dI99Z6/6WHM0R4BcZZIWWA4SWbJ9SqKqcALNerbJgVJS15WjT/eP90cQi1B5uMXA
mzsgzOJqQwRWUrALypStpPtIVc+pTAVdGF62F6fNdJZQ2qWjvzeAiWvzoxqpqQ9q
CbNJRfXKab+yHbipjByzfgAsFOQm+FLroDic70Pp7N1BOmM77zVrrcNlgOkzj1yF
uaeLrc8YB6++1Slqb3MkF3gQ5IvbjwK+rP0OdYlXTElKx+eOYTs4pTe+f/iUCrNa
gMGyhcCkhjiYrLct2kgBioT7rz3krIn6JZv9whNhS5CoTztm4Nwv58lE39XDD6+6
CDGzEfOr0tqUxj40/4aWP0jc/rKGW9lXKDD8FMgx93i3/lfWbhYFYa4IOaqgySj5
T3R7aVC3EAWfsrycQNIkZ598B/qhis8rlX+0wWzy/eG+aE7z1i4QM1PZ7/ZVC432
dyxknldGQwBnZ//sEN0/aBsBQ6Q8kBTIkHgCjXMTtMhuQ2C/xmY01dUx1Wp80lwE
fbBnNTC9V+D1r1hEHyroLhEDCcjW21eGKqkzJy5WK62XnXcEJC8cEeg5QU+KWNb0
87bOh5nxfE/zH9SJy4XO3z/2txAgqzcCxKKyw+8aK43VNESYsbng03lJbqQvQqZl
6pDTvkD28m3T2uXZDAnlOSt/XI6k2bt0fSf130lhv/bt8W7m6W48rIKF660upLm3
DYLEerFhOszDbAimRCm04A5c5h+pZ5d0AHcgcMFjejV/8+nJhTj3x14B/Dfh3GLp
VP/K9NiHY0S23Vo0Pws0iAUfUE6XMdls71q1bSZKALBjmx6y4IL9EZX91lbMBHjz
NeAWRhlZOYbL8Yy8ttPzKFkX0iYRATa45c9tvH4eWjKGIWE3UiHmAMBiuqwc7ARt
41/7uHDr7T5CmX7L6ErZljjorPVFJ6iugPNkdaJs/1MvzssI7h1J2Cj5UAktLWs1
fF7ij6b593p6QmHn2cehFbFot9BjR5eUtwl5GJ1rsg7S/bl9Nvc7KiCu7XSd28JB
SKZv93+ak2155ZtkSi9j2SpWT+JKYTE5sQzRqEMVn9PCZzCnHgbxm0u5J1V5Lzi1
DJZrG5a6USh0vnzQnxW1CajFpLCZv82bCAh/Oo8aj6WIbn3mqF7a7ewFjqk/hTZf
AG+nKTew2lD+YU8Q3mVOad7oXo1iVs3FAQh1hP5GEFYmAKdp0xbP49CaA7DeNvnj
oG1T8P6jnz9/t5j5v+S+t/MADOcL0cHNOVsESCh1Kf8Wz9vVgO44uK6quWm0x62N
ubUuOaxUqVKjpzNzI5w4TtIxOgG2EIAqOizyX9fMni+Hpks9b1cK3jQeSbvEDSHC
FT8u+y8SgLpxbz/7XSAmAZtdyhWVvD+w7SsyQBgLZgLMUbvXWV8lTwCKlx7ZyMVt
AOhnd2IxXEgBsNYk/u+ADel0IM/igwrRqYI1ptXZzoRA9bmTMG6i7fne3J00axR7
8TI1yVVRU0Hqus4Z7yVQYT5sRwuScGbRxFCmn7WAt/U/dnKKp+csnZfufYA2G7Zv
dJ0QPtLIawjARo+i0F+/7D45YORCIztpoIKpLI9iOqJz73QznMwQO2zU13dyiXfC
7GcXerVpadGDbd8MeRYsOJQ8kBqPof+qZNngoAka4kq4jwVEBmmMhL3XxUDAz0wu
j7bQ2tSxZCwbL0LbokJvCZwwAjNN6FNMFibhKppRYUncAgZgRjctJEL+MXAD/yZW
ToNM9tLpbcTYalXsJKfGWeMKb9hj0ref/s8QECKLn8WOk8xoMUt5EkL9LLvdtc8U
94yTgYMSnMTLb4OPnj9Dp5v5AoxCsVcovtCXX9bEP5+gTkBa1x440jLP0zMEesLs
Wfl8e59+7sXkh9QzKwHG25Ibbcmu8UnpHP4+ibwBIRYmQFYkOtLAesdjpGYyV2y+
xo1zzN3VywBFGX/uUw+lsTdzYRgokWJVT9X7guY7Qb1lWSo/ThpNB407pV6xw//U
FO04R+62zgASad3bgFSVCCJ0JWTrY8DjgyuqbY1jsAQmhgG43fzPHXKt9n5sFt8V
Heopw+uSU7kEeuWuY12fM2wKeLn/rEiG0MhAoAJOuE1tyjTTtrEvQt6r02kQXy2N
FzgMzS5/6GyM+uHP7fB2XhAcQ/eZs5qVehNPz8hq4sr1Igcp/0h+9hVTWOvSjDzz
0lDgpvXfoKKRt3oO3CLGZrKVywWH2v2c/U9lwbXEXj10M//QQa5FgxWqaqdYz7Pn
e/NFqHEnOY3HD8TxFaO/nUSuk0ArvmLL52pD4s3Dy37NR5Uq5siq4UD0lTaedSsf
tIGlGLPHNF2hhnwC0ZtFetgr5vG3q0Glgco+uLbmy753hUUmjMpt7VnyHqNA+SG0
NW7F0vDCbMtII4Gqg+FLa8FKCPPAMyAeU+RifvtD+MPI6Qx67BolbuZn1b8ZK6AK
Fd3UIRMHiO2Z4dM/o9BBDUyUhpamKJqN3y1YlDQwRBLRHbZ67txrVTIIplBLWSCS
IF/Ws4al6cpNvyOGvqH5gsgwfDBaRW/HpJnIszj6oIJjAgnvHCk5gd7IBKuhCrp6
LGoeTJomKIzVM8W4+SZtH5AUvE6Lr37WXWwJKCFBVafVI7CrmeOxstUkCy9+Tib3
6oww9DwJRYuy5ur4qs1hMSCofs7gxntxvahIy6W5RfyvUkZ6zta/r5ExssRmVSAB
ga8N4ssazdq6qL8r4hYGMwT5B+PmX/GCvKKgHSgYNJTC4v42UVuO3ysetfdiP+nZ
ezibWIRyHgmLeVoyd8CEdWxEFjI6GuCEcrjoIRn6J934lyj+s12eOzF+mmow5ptK
VyCAx5yfTpX0gE4pnRgPfvLP6rlHp186ouVhkLasEZ55jKYY4IIQwKsGPJvxZtOB
6XVG5a5vy9fYBaAT7gKGaE4Yf6lGXVt0BlLweS76H1ZDPL4eFTC9tb8CcqP0tfjT
lB0rtjD/cyl0BIxUlixwgKraIic6/UPiCmCvc0mpH81wLef+fsAR/nkPVTrrQv/5
2SOTzj0EzyqUY8OGP8aufWH9If6QyI02WAyT15tQnwil9+3mWPlk4pDRi+xjeHn0
KETsk0OjFv0TSYbSx7/kckTww4kY0Wn/4HLM8EPFqR2v2QZ4Q8YLGYE/Tt8tC/xo
sCK8PESPFDpxJ8ZXHcWTGsRNpPUoHv8iw9XznhUin9bgkweSxpAFyy39zAJy8S9X
otnN2GGVENOagsmtJ3V5D2GF0TKjWySadxvggjgj6gViZtop4UBQO+tfTIHJj2Lh
mz2gO5+ANw1ln652/IwhfXJuYq0frGmo1BjKluIGlmDbm/E4apS641XkNFuh3smO
yypXcn90ma/R3xhk0ZoHApkPdsQ3utc5Y2uaZKP75HbzreGkTpDCT2UqcqtHTd3+
u67k3NHd/YGnCJDaVOgAB9cmKnkZW0qdtFxgscSaV6yp09pQeuxGGMwnkOn/DG27
dekJhOB5aYg+jwgCy0ULFPv6kviuaVzv1I2+luuby8eR8bcE5Ob6rAjdwhmuykXY
2oD0dc6pvsQ8+E6MPIOh8TJ3YyCcOVFGe7c0ORrjC3nmCIm+KrHDaUuBg7xyjrGn
jH/1jK+NVAGAV0bdUZBQ5ZWAIMvrDv0bg6TFUmXfsOoy4g9OAXfRL6m+aa4Cv09Y
ceRkFUDWdVmuJoQhpaeJ+VprWCOsI0nCMzI+B3Q7HUz2vXPyNGS+4hkddMd80EvF
qNqLydGlQE4N9H+/l3lBwWiAOECKm/olVzEVGBqK7VCm9bwPztudJEoYMv6RIQ7O
14ycskAdGlYkO4zmB7q+B8SrGeobzD6QvIfBg2MOrI/rj8J+9OfgAsq3wHXc02y+
uUZxcigC8OpGOC4yM0NPW9mZBjCDZT5xP9pDjHFE9C0AFTuQXC1evTbDVZs02FjC
x+A3zeSXUneU2w7fhKiT3QqXqrXqhIMwRpiC5so1c7v4PYqIWkq1kocY9yEDE2lw
taVJZgrEEi1tka/aklGBIcNvQ8qsQgwWcMV2MdtUMIZZwYy71ZWZxPFnCMBPXo/Z
P5Bf38jjpUIeX0/r68GHL+j317lWybS5aqVAHC1BbnH4EjAPPCJdz3CO1IVgDXEh
lZ0TzBmHTy/IURuXaKCISnEieNwSPqh9TqNEqUCxXWqtEi9V7C/USaKaFZ3Y+c0U
nlqFUY+/DGqP2xE1PBCzmEaMhu3S56cNHgJ86yseczKZlKs2teeXapo65JzIv0XW
l7hEPAg4bFjzryYDEsM1kI3+0K2TK7uNw3rgwfThX8bFL0Q5m6mvfu5hHy+KbVFQ
zremczXG1+eK/nQP3Rpsdcu011TvbiHZ9x7yIcLx1fEZBN5QMOSHArGmGi5sSKc2
KS7eWMO82avKlKpxgaqAS/Rd86vnkhtLkoIxNJc0sSM8b+VpWcoHfoi1HMBXa0nm
kBccMHf4l0jkt3hqnxYpq/2ekG8Yzc4HgkS4z/f/6cto9ZetZxe97Pct7BCdik9k
WqN4qUG4F09cs8Hryk2IQlarjg9Il4CXFVncpSpYNv5Anm/W5JE8eym+oXrkVpvo
17fS/LD4s/mDMohrmDi7BdIV8VKSjRktCJ+/tyL1Dz1OOUZIN+oiCtZyQg8WwWJd
jNsjoYkjhLih8rUVoQLNzT5Bch97gI6OX8ECHBDGkDQANsHHffwujgonWpTCfmf6
vJlWTIyzh/mfnWFYV4iWyVr0XcEWfs8BlO5vUO0zjGrwmvTU6u1e2OgsJnzoeidV
P+R9+kGhivxNewFe4COgPQqBT4coGpdkmAuFrjfTkACjSpsxG2j3NzCQcIZ6RXka
o0jB2JYZKGXWqvNDSAyfFFo2jV1aTo8c9TRtO7r+sYNH1ihP+EiAVD3ZaXa/aDag
QHg1o6I0bsFymGRen5d2QRBwlCnmySoPurvLq8CJX0yLQzHmg7S1tfBbRG9tcHLp
vuHXuEoSzEuuUm/m/oXDgkku8m7woIV8XWx46KmuFp3nS4RPSC4lBlvKcpdQjVyf
X/dfl5UeiNadRyMudQKKuymIIAGyx/3KQ4afYI6qhkpTpzi5tlumsH2socAb5jyx
O0RST2sCtQWDj4dv0RsPHKatJtWtGn/8lVs9faRDEHV1c48UcmLyp58kj/ewWveV
VozorqzhE5DW3VzFMI7G76TDEMTWmgoWsdXOyJHm/ue1zFbkyU2keKBoQsdSl85i
ATL5Z6BJUGvkz1Z8FOFFb0SJCA/rXzkIO/m0li4jQAIMypVcYihdOeJ/yOCq13E4
vSdTr2g2ATUSkdl7J24jsHGsoQFa9M2JhQN1I0m26MUujbjieBvAw78CKMOnYF3s
QIVOyQZ7DuYbAl9YVwcFrh81mCrl3lp7GfG36wVPb8Qup7GLFE52bVFjXI04Nclm
gCKCqzpZqUfWjWi09f5JG9UbSkTbDfPb68I84FpIhUZYPQVTBiTFpr9eNAJ7mRAd
8smNHnUGD3SfWwBjTMoWtUkCbUEAomKd8+O3zBb9fXXwucf/r4VV8qVjzUPedrp6
kaJNU1OdXTyNojbiGWlglIb4YjES2kp1DBF3BlQ/ilsRkOWpM194apfs8QDoA46O
uAh2NoS3IUH3DbIIhT8+tO8gHeEVRsdeKKXCUSRbAIpjonaj5zXfNhJkj3elSiN2
+XiQ9l4VnZmaNOerYnmiC4Mi//7AqzydwimqeQ4BisYEOGse3rjyuVf/fGNZN4n7
lIHAV9s20sVXGI6dMwm5tZxb49JyYcBGOv4o5V3ZhcvU9Cm0JYYWRkmO0khVziTH
DU3hAWO9WjN0iQOAcsd5XhOzrBmlGSFgzln25lSrD9I8KAFu5bB5+7CMDNN7yis4
/iZEOId1nmXblMLgzpd8oheAy92/foXey2vaAePxVShtD6V6oP5AY39PtWaS3ZZJ
4Nuozr6i58bwnBwQGaJSsK7nXHzbFO5gQtNT6ad/XHqxWbU8Ju82p1GzHLK3YZwA
Ex5Cyf00QboKgHVWBZU2OXBq1efOYXAVnZ/GECeKuPDRfBNCnM3EWkgn/1xvTUu3
gsaDPb0cs9tvBzD9dlKNgAIX6/WuoHxV3O3KxGwZyGfGfyFKFBxcJQZx+hKuCAcZ
UWeoKHLBmJpGe2oDQ/Puf4gbPWUltXEI2egDLsa20a7W1UTv/LyW5oQI9mTBojiv
o0QJvnK97H8wHbN7AgvwvAiBXU3bnDQvLAIokiTH7cUxTPkVmRMbg8CnnN/OTN6S
4FBdhDAXAzMJoOyQfRY+iLWOnDwLTbyMutwG37bwHh9G/V4YhAUgWCtIGTnXvoH2
d8enfe9IS9TX054kWicAWyIPDEVfYfh8drtw2j2wm7smrBTln7+okTAMHHPt9uMk
Fb1GzOc0etgIbVTvIBj69RwxjZ+yL66QV3inhLeq8oS/veHzkbnHHZYqXp2qIud3
AVJc3h9flTVHo+/rjg1GKP5LnYurk86dXmzOgGuDqJgEcY6dAQqh9/PQJOl3Q0xt
BZVr6eoP9w9W36I6zHecHmWWhxFC+QAMO/Zb5NVzATr1vyuhTGcdwV0RBcBhIhwp
gK2MxoeDBBExwcX7JSeqH75pXlCiI1UVE+k2Ko/imNqSWIHZ0hvDIbcrkxC5vaFl
LitrmWV7nJ5W5jej9WgIXMg+Xbf8QEfzEqJavLXbr4O5Zcs+Mj/I8RBG7O3Sc+79
fF/ndsdd1zjY6Nu2OHwRBL58dSBbVyQyhWbZfa5B+zvP8BYfqCEirHj8IewylfVB
W2IGA/11Txy7cx3VkT1I7Bg6Ml56eEOHDF1mYXSKo+gyVT+q1fA9Bje8pYYHer8z
lu0Ubt7aE1kOv4N5RWXKdNpkHL0898fSYSoqeZQR9hyXizfOZZfPXuL7AUQx8AYm
XM6RA1HM/3o4yhh1zOSS0pI6du/VTavKydB/d6pEFnxsxmOCxX6iruhzvJ/9ZyAK
1DJAEBg9SfDqaL1zkMhL2Rvm91aveHImwtlZU0FwkiFWqJCI7WFTq5767V+KwLyg
L+XDYhDVLz3XOdkppDQ5emZhChuac3lt6Er63MRiGcTUbDRtciwt/o8+iLtR6PwP
rkBglXNjRUcL60gbehphFNEIbtgd74KtTtyJ5DavONHdy9Un2VTAO6Efl7xF2TZ4
/6kGc0xoyUKJ2vBb8rtJfa7X6ydoX8WXLRC3fKnzZcbMwz1nnRFoH301p426gJVa
cN+iVeOUCV3y92Qbkl0zM9QuyhBUvt/HrpGpLrP/XdPuv+hllZVTxJcJw4uOy7DK
EaUhr6Y+qj+QzWtuflivjVJAEVO2autyaorGK+C79yc/jRLvEj9AUFgfidWlHQU5
xUpyRO6qkgebcUNaWz8XbKlDy75jsZRIOvfs8V9TqhzWVTKi0YjXx+aRyzhUiycA
XXzY1VBc3WVvy4wBL9D65uKpfvCoQ7Fl4DOItRSH4qOGTt7VQ3z03GqTLheiRUV2
EZLsPAh7uPqZ/hYSEYVw8X++PI13UGL9GS29AKitHCzDFS79wLmi0AQtPxKmLv8Y
kz9wkScib4Kog8QuSY6j8V1+p7u8wf1wYj8T9a0dWAR1JQzFzJygUt+XZz5xFsEg
UlRzwb6zMJq2ETW/PQE8ngUhaFlpvnJNqcK7vp+ldL9rGqxy6CD+H73GkDYpU5Qz
byQmhn4zyh02B3LzCIUNIMVuyyyapkvWwwiSW+VQ74BFB3r3dF6v9BQtarNj1G/u
tOHV9uGVuoGgUKw5OoRtx2SjK18Ez15AZQma6JrgBNeHB6+6IPJfeR3Q5v6rVRey
Vu0NSBqY1ZHiVRMCvWwMU1VnL0eC9pzjaA3zAOAtPJnNNaUFVxQrCcYQhE1NAs/2
fXMvg/F4itNsjopJlDe7k0/lNdSfGPDf15y9uec48b4syuSQahdtwotCDzuDQvJh
wL13wYA40/uLBVtaTo3oz7Aydr7a5Kw2E7CYP5bw543sBKz86qmgNM64EhMWRwtZ
h6dv+jaFBVCGVti8ZrTcNIRW4bIyKC4ojDK9XPoWXqceX+Xiwl+K20WLEUOxCQ7p
SHrhC2ce6X2VuTiQ5Gujdulw7FNn6xRCLfV7MF30Ahr5MCTHrjpTRhVveKIdUSvI
zV8lIQPpxAN8N6HS2rQtiwJcTRv3PGL/P0iIZAk3zkwJ5LOb5RH7rhXWQjsGar1b
snS6FCFw6I+RLL3xuv7dpr7Y8d76YVnFNxKMH6ocdTeozk+UQzXvxETQ5A67qbfy
g9iWan4m5QTPhUbQDvHdxSC6+qjNvOsObPd7/efpYbvNIe9t2GqGh4/AlH6+bLNv
pWMIAqL0PvpuTGds2zxwmAORg00I/oJ1BChMGQ+ldB/VPBAcj2fGNbmgCI0/VOrM
iLgy4WNO8Gn73+o6R8a86sFFDPpMzhf+jon4emf5wfzQXPaYM3U7atmIKyFmkoGd
6am67B/l3rnNtXr/d6qTGa6gpsL8ZsmDkJhWMq8UcL8CuCecE8ZbJ5u5qJgp0t2d
BcDq0lGNXEExLyQf0/XEcuGdrXM7zPZV5v/2GlJIDNq/jxFGpz9vgyUR6FTxExzs
ouhs/xL0yxOnJPcroz4GypkwV6m5+YJR/PF3f5m9EbISorNyWaVTA3UDv7pxjFIg
ZU+tvH4snHiXzcX2hsObl3vfWiemOI4DRuPFdUcVmSbmtpARDyYdTesmz1QaOp/0
t78O/duq8FfcdXAP/WpV61zVZkFpHdmqyR3LV2+vEYwOVvLs4yHv+f2QbjXStXB0
9KudypWodvliwvenlYCH2Y2smyCaRFsGaCzoDM4McirUQM1UN2t20kabQhfkarl2
I5OYtXp9NU6D9inSqi22T5Iu3bLgatXxdyu0URxQ4P9aPSd0gTVP7newxAcbh+Jr
gk5J/2XYDxvebN/ROzTS8VjstvtaVI9MqdFjjrAxUOv92x5jVYTEj2HVsg4bcRPc
6L7XYukObZpYnoYdcaTY5MzifOJ+T9nlAJgiII9EcOyNT3OVQt7lqd0ok8QtthbA
fIj4GTkqmG9CGy0/igkFLKKtC42Zcg9Syxm+bnO9yDFZ/dOY0NbH8tDfLRRa6Ktv
Bj2jgZys99bLwDxjglrZYh5uy8vIfRx+GGuyK3ZkER54C7aa21/AF0wTu0j/s2gj
roWogYV9DWD5Fw+fL+EC3CCt35WxvpwzIF/f5pVb03LLR8UdTzVl9GB19wWkm6Gq
3pG8CfpoQ2UUJXRv9fuYmqcEwVmcLZ1nIat34rK4ArD/Pm/g9re/0jCqI+x+uUcJ
Txd6ou3Hx9+GvfldulrEbYF52oVjK21w6Qq+831SDoxYeLcJ/CQKOCwKfTM3Ldz0
MKm1CXIx/2gXjTsQFBU9ehAHhSH81/hd8K+wTUyLmXjex3GM2J6K3MKVwBbcRmYc
CE7R+J0c1vn5VR1QOYZLfSqyk5FkrX+bcFB8vCf7FsPXxHKGTVZmuYn0ogCxbk9+
+T+PuA0G97mv2Mv0nh0QWqGsg3s+3aVJUXp8IoaYdBuQQzXP16qxCkCSgY4SQPsg
fwGPQM0MrDXUE5DdMtHpYISwfHUCRyXNjGcUbcAOVHUHP5Vp9pqmzOBJTWgQ5RTj
1VgR74eNV9Dyp5T9BzUzIIguF7jGAUWcLzqYa0tyDh4Ou8tJPJpCItHiBdnCrzVX
lopGBGnFP+DqtXKcF9wMVo85RkG12XLx/GsJ4f6dJATVWQQspOCqn6oDbmlCRBHF
eArq/nceoEBgzekeZZvrLZ03pwiu/muBX83GV5j6Sx5febZlw3/SXFhYSYp0t7de
nQYnCirB2TPhKSPFsYraaCielAnnAL7bcYVbe22vEadVNkqRme2IFrKrliiXkwWX
tlPld9NyWqs+WkC25KtYp0x/E3XDiOU3w8P1x1QWFsUIFtIZxN2pauoiJIfjPItY
45tRN1ivaF5Hh5z6+LAHwoDnOVLoo4Ub37hlUAB/WUswT0QJLthuTm8liXWCKNxY
9gCwDdYCG5S9lQqHcLlvWFiaaIkbu9mz7IscFncKDj4eZ5qAZG3t114nv0iNDVlT
7k3cmeh+kRu6SMlEJ1JzFhTb7FAhznYY3gSmkhF+nqxkaJZOcXmh/hXI8euzGtl9
2h/ImIqcFMKKrcPbCYmiWKp7GmkAT1BNurAL/aFqer2jV+qpl/upfLY4VZy0pDp/
o46SweOdqyxAhyUi6iSY9GAa2pjXmhgNg/vTfDpi/PB/2lpmDJPTopKUHdWjM6n9
wpTET8e5wzj6tzSFd1vJOvoK42uisjvHUQT0YVLzmwBz9GR2YVb3OaanOGo6WsRE
WO8U9/dSY3MQJSH8TKAp53t3c56/Piw2Vw8AFa+G1WaNzpCl6nEAJgdbzSQgjAF0
JPTUEA4QAWmrt1EtWP39I+dJKkOhqFLvcA/y+1JPZRH/yBKwgLpnq5v7q8m8bfem
`protect END_PROTECTED
