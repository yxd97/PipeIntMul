`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dg09A9YW63vkS6LBx/uECXe+1h+pLQ5QVydAqG+ALBvqVrHmdUZ4lhjkXurZoZkE
07U0ofd6B7UsyVJPyNJMM4hjdmWXunfUh29uI76BCncvYST6BxOUbljuug1rudoM
1KAcyJ2bhHigrD8YtNW8VvDAIvUolJA92TvzztL+0ocMVhhBnbiME1jeXfSxac6D
Jt+rI2Q+lK79BaSi+vv1bZoN1VhJ4kXR+gcF/qG9qr70N+2gLox8r4pXqbIjfgSf
nt9i13vLD2I3mxevNIKhM5raoG1iSTlWvw1J6Z+80QjXxIM/Ua8gYJtLdXnUct+K
ZUK/tk1AEtFnMDfDgS+KmZCqkw/IVn5j6sOJaSonznsaA7/OWkewhSp4u5/GYjhQ
`protect END_PROTECTED
