`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ZS9P+Rel0YRnZnUmF0w12AlTXPYRFNShc3Z0K4YV8dLaC5uIPuUWeXUKuPpS/Jb
CuEp011ir6JXxvOoAhjBhD1dqtyf+g/9FKakuaEaKdJTaPRdrJnibEUhBYa24gIE
OueCxTL61EptlzzT4KmFswd3FeSWbhNBaBB86q4kRs5xoGU5x8wH0tAjSWm8xEtk
YzZh8qpTw8OK+yhc1T4nMj2O4agNrW9Oe+1gxe6tqugjRz8sIn6/dYg4zoca/fJe
ujO9ycbFBw2sn+qIMBGbq2kFASg9ejdELTqNYGGnA0gX0ixbHnYRfNsn8kCz8g8A
veKQA4Iz8aoHZUlhluMVG0BTjacJxY2YaYGd7hbEDIz2weMjoRMYGX16HNKOE6z/
OS5IPfikG0DjYMC9y43zHzTp1vbBcEQoyY6tvzl7m+5h4ZJkoB4R6JbpJSVSlPWR
02mlGeIisNYsLI7I8ZkmBT/bVUofchiYvMeBaDEWGmqD8hUYEWjQ0JraQXuJnNtv
xxRJfmoJdOq7LmfP8clhtVgvcamqAz7vGdnGFFljkscvaiMmYE7+p7enJsf/GjdA
UlB0ki0B4k5CV7CJU2efc2GCfHkob5x2fv0QsovHiqvUxUmPv74Fbtn5zjIRRg9X
gAqQ7RqPP01UlKrKW4Dr7fVr+KM6HZn4YCgF995Q3RBWZX8doltS3JZegPoUarob
z6bwmiHPBs5C18df95O2otsMLphwbrDWYOoQpDqmpmqQ1C6SOh7MNwhcEnks93RP
5S9J34y9UI+NnihFYPLTRNK+Z6NnIwm99N525KUA1L59xE0keFB3F4hWBXU+oGpp
g7Hoqtdn0y3s/k5MK5E2JcpyNqZXE9RanB+EK2XBx/2BZRteeHVmR+ZDvrvDb+2s
OABlfc9BSn9/EKZYGIhUNZH+DkCv8b/85s/sTvuCTOH/6gOkOUeL4tukrzdMzrcm
RhY8PQfShEB2LV3ApSeBbhunzfxVw83W2xu3Gm5+pqDWAD9JwQ8FDXdXnijt8t0c
MWmV2rk3nsEx5ghnLbSktohNBr+KUvM2DldCgNcpJIj/xhyS7gsrb2MvPxrQsjWY
6SPX2PBRr2rh6CUn6CwE8MZ+kCb6n/FCBzu6uCZWA+P/iTw8xk0SNLja531jvo0O
7V1kv6qswiZ5ViH7PNHFSpw6ektNx6uvi4MFsV/OmpDOuMpZpGzv0T6VzIQ6UyQS
kMLrMTngEk4qFsw8ykD1SlojKvYkpBxfhNppELDF6Z1QYjrGR++JFiNcjlXsjoNW
hnF27IluackTsfo4S6lvTlTcvxEhvzyPklT7fWJ2J8EQMQK9ctFO+IO0BlvpvykV
Jp57ELT7rH1PgrZ+iXl4JGrlG1syzSXSG7NhsYI8oQjzy3UYHlnXvIWQC2D5sg7Q
i5j1S7+f5Y7nbtRtKj9VNb6hJxA0orRp0ShHPZtmIVud8dznmpYBsnN5wU/Ot/8s
80TdbnrWrcHPkhbyM3i2wVwrgzGhFZpoAwv7WtIYhsvJGkhoj2lnRxoS+pN/D8l9
FpVkPAgiBczU+8zn8K16pdtngNAQ7C3X5VsSTt6gMZR1RA0t+9Wmxt7zYGN2RCOT
HaapzhKCCDW72pK/Y8p+e0leAq4DEkUqvok4amP1/vSNUdSVtuXTdDR6IQW0smcE
Bedb75q52U9K68go+jqgqEvlOGKKuPoCdGy/vBCck8+yC7gE0F+A03ZoXL04yIyx
DonQVSv2QPzL9GBzwSxuiRqOLIhI6mEH0S92MZoMpwmat+US7iFjEXPPMdc/2oyQ
N98D10NS1z+z+NGIr+PleR3tHqrbBWbn6H91YXnbyOCOSxUtbvREFqAgthFwFe2m
xM6CmlXUuB2pZurBb+yiKzVr/vlz2qsV+YQnrfVcxwhZyqRjT6wGnffnPJ6NQQiV
aYXwIVeOQNcELJn9BkgNUjEHanIFh6bjBLkXJzBXRapNHQftI0HHcfa0o29eYff9
BcAlsqONLNKHRUnpDTAEF3AaNIRdmSVRatXH6IUmcS6V2l1YGHVNq3zL8UtruEKu
p+3gFeZ6l9z/lE30G4MehYbpb0EdYgeRKu0ovetcE1yYPn5Gw7DMsK9OeRrYPaia
mVjEYgU20CPVuXBL9kfagjfQVvRGhdEQJon4IwfUzS1xfiJdMT1nWMbJIWfdV+jK
TTUTDz7FE0AkKZAqXXl6vPdScoQMjMKbyWIR/Y+RmDNch8KnGJ83IaDBIX86+HCK
4v26Z7i8x3pj4CQx8iD+5N5RAC1KKeS2ZQfRWeAkF0uSLDeV9B/6e4h3Ul0fZ9CE
iarDsASiujPjg/dU1sVil5LUJJe/2wYTq43+ji/GDvAmUQU8aRmKCuW0eBcBhsBT
idT+43UvgpZm525moEMkh5hWesMOod0wcxunQhSkK3smrpw6+bE6QZ+BAZNbs0FX
Dw+Osccu915lDYxM7NmW/+s1/he3I6EvtQ2cBcB8KiwbAgppQIuxZB8Uei5Q1lxh
6h10iwCw4pb7GdkjMHlFKzU8hMmfdG8uONEmOJGe7Gg=
`protect END_PROTECTED
