`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FXlxXlCxSDNGRWnqZ7ZspLRQSqjaLXu9GCvlZQi/c+5eLPd6xwQBfOeYU4D49NxU
eQqu3Vf0STvHepAlD7SY/OwR5BknpX1jxTAgMekPHyU5xx35SAgVuxX5LtieosYV
vNOusYfZD+yS5gAyOsNmOuS5sQ1JSEwjON4Egw7kWyoFqFz/NBXT741FhC2SQGuQ
+2neoYZ29t7H9c7nz9bIaUHhgtKFJY1Cr3ML8Fgy626MnJpLqljPF02FTA67lr5t
EWSg+i5+QVJxAFTGlgIWVsdfhiIESacqiwCqMi3LvvNzI73uqCEOOEGkTw22+LQO
Amni//YKO3GNKiZzgRAQT5oxeeP1zqI3RDFj7+HEaJ9SIaIZiw1ZmFz7xixjKtWV
ERg1HC9nLq4NveIKdApth5LrnSZZ/dFu9t3qn1+OufD3DhiB0r+/oBmkYfrTi2C/
RS4s8v00HkE+TvegF1yvXsHE5yfHF7fioZZ+qTy9OKyAdqlC9mzgcE+nKxQOk/qY
GDwJXQ2JdesTDbDfJYma6XzCRt3+2N0loZQq1xisylKpy3b1P/80r6vVZDGZzv2a
GqBcv7DV1Vy5tuD3epQ8L4Xb27acEFi/2CaBfd5nHUZYWzCyI9gn1QXGWVpmgBpE
bKVb+7KHLky2jPslslNJgCU3fAAukw0Gj7trHXVgZT+J9W2rlzXnI3ko6H8O/MHX
OsDce2UczpOw8t45e60ZUKkUnuwM3GOjLFBJfbZ1Ussia/p1KeGQXPH9mmKZVOUa
ivIp0goh3Y1FIAoXd1EYNfcqdeQ0YYGTNswID7l9aE3NkVmiZZ2lExu/yWC30cMe
lLrU5hDg4jqJ2E+0q/Zx/Vz6t2exy9zW8LyhDKD7+F9giIcbfr2q+27UmYNj/AHI
4amI6Xv9lASfk8kd+iqqZT6o+HRY8w4gxMM7WqhOR3ZieaQrgdSQ+AXRVfKhW/61
p6sF0snhD5dBJfWjo0HlrDKXgy7NZItMOk+0sGAWnbpHkwFf0GR2t6F3UxayCXXw
iI1DX+qf5Ee87Rz7Ip4orBW6Y3h0NBT67Pn24mENKUX1CFW2xgq7KIqVQbMz1Zom
n5UTqqVcN8I5H70tN2+XcFEBno8MvQEpNUlW/c5Coc5raIcyplfvwbqKoMuVMYHT
ZTevVc8YgGma5IKb8Cvvfap4wgup4U4vzHY+9bxzvhYfSpi3Mw4ZTjLckkdegpYx
QGPySoauliwwKC/W3G2hzzbmUUE09VyDV+J3jCiwRdelm/OLkbB3xudvlsGy91Vw
aUKS44cApvrhlaT3PJxpfd3UDrk/fgXrUJfCSBfKznbFHgmBvzOvxpD+0QHwIt4J
6a5fvhL1B64voV5IOybFCmQyz36oMtBMxChTPx6cfpYlIZJvJHcggdM4dmH7q/8u
UOAzK+z+nCRO9OG+9NWlvtLKq0rRNo3JK2bUO5wNtU1hD4n/C6A+ZC31AmeJlsI0
R4TSFBsP5Ht2jAx2RDKIUc0FJpp8/WHQkdBpQSYftXu+L7bpNK7vMOIuv7DUqYPw
EVcyhTgjHDjENzq55XOFSdayvu22K2Rnhv5twzbSZg5xSmBS0vbyuGfr0cEnvUf3
X8YGMSYyK78UiSUxRwYsJemjPcOBHPxxhAEedorbd17gqSYKYNjeZZm4OdmcgZML
`protect END_PROTECTED
