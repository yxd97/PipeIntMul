`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n4Vz81SBm+6OUKdZZRowDD8/Ldj1kvEEZED0NMQIvxloeaPUAqBwhJtb0gBOogcJ
ZzipCeTqJ3jfw/RCFJCBFafRygiyb2wWIE/yUOFxCoH99I1ioSbVjbylieAIbHqt
VYkMgB4HbawQJ0l0fkazcgqi95MJ9VxDgAIuXJdtyQhoXqjHblTn8AJ1qM+Y3n9T
NOSoMURQ3C2le1+QOlvQ4W4Gowr2WsVxp/s1FucRV2d0oe/63oCDpjlIxIuS7XD4
cmYnIQL4982p/HOr2Jl8g17y8pBDV9zRbpIc9dT+vZHNtsHugyNJQgHRpSpdW1Ab
I9pxEsxaZeZ7egbX4aoU9GV+yxZpDdkt2PGEDuyUhu+aNqcV4aAb1EZ5DS5KcUvS
WvS2dGL8avHoKIfSORKpVk4tTJg4HvwnFVTIpZiJE5RoqhPnDYhFoEQu6wXaUpmB
NUZ5J8UPogT4c1SrN0ZTG99pXEXfILmIGDzCeA/0YvzP1meXZBQzNotuTUTNpkMt
yRlzEVo4s95OKd/OBrRBBLYJGHtypsGfk09sO3/XSFYYh8Vpr9L7YSFcbeIC0H1S
5shI7TSCWxHoYVDdrGAVC18fLWP+J9HjP18dzPqETRX46NyfTIzu1X9M/B8NU5S2
oRzYdgAnaFAae6Ti/BwyJL3Lud+WL+4w4GIc2jeb/Zr3vlwMSzShqI9okJOd1iOG
IEb3gyc1wd2U0sRgl2Xa9eRmE1nOp/xcKrzyjUqcPUttmFzqtRJuC+BuVEFzz5g3
xLBkt2PjTZDAfLIKXIQX2fZPyj7bt2RnwT6Ztd02C0pevJSaHRgc+1jN5UUuQmhY
XTxf+NLyObMUVS2CMjoDAZIJmoaslYOOUJOq+U5YCEWMNmCGaIRmJW5O/XTMxDuX
Y71G/l2rOu9fEbBHXZb/XwVi5k9PFZpHSEg/wJGleYecpsXWdl991HdQGOZvjG0S
QAQQ1UjURReI0UDKzQprz8Ua7xy7NudrJV5C7IYibe0=
`protect END_PROTECTED
