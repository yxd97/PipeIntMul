`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFBgMv0alziOLlGoEFl79iW+VL7ukrb/w7icqLmA9MQE//jNZKabi3/wqUqNFcVg
lI3pngzXD7fMF/NFYKqExSG28jFKahQoQt4iAUhKE5gGUTutJvOzD8PoQACwlF+X
4Dd/LtZPfXrtaK9rzLRgl8myynVEx6eHu9tIY4mGt31TDUsUFgSqv6gptUDOtMdR
Jau3oUUDNV3ZSpK9XCQNSX8v5zAjfZ3yrJ9BfK4LHFt321WBha+vE/fYqwMK0FOw
LYSs00ABPD05tcPJuT3rnpAxkj7Gsm9QslHsv/VAlk73ZOPaZAnJvR8GDLonL9KI
CSc4WwXZuIN9SkAunvOlRlWCGkC7pzSUmSucYlg0BAl+Vu13tkTF6971TEgqPlJH
DXoimaJMARtnyvbhzOEeEkKjXU9vqIrh48tTnYQ1C+OsebxTOM8gkusp+TbRNar/
OaZuG+YHMgps+qs59EAhySI7axOXeRU+pzi9YISJuAJ6Xld7yLHdUDZU0QTv3TtG
IEi9poIiyjOTm+FYEyWDMErxy/4QA+27Xr71wlf/JkT1pQzPgEggfNLnks/CCKum
aB5DE2PasoTpyVRvzykfRjUycUtVYVtOd6BcZw1kLg5w6dOa1hrLVAzO7wI17a8V
e+958PVEV632e0Cy5xppf+yZpXoHKPof6FYy0WCZSzgmPH0AgjeC1HlLAR3qZaUx
3sj3++2AlulWDb5RBB60cKZgO/7I124KGPXdd+EwssMuWtbCOxfeS4CEBv1YCc6x
h3SLScKiZvzD0TLAUAaL3QVWyaPaZ4GpzDTBEWXbbAanHJHVSmuSqEo9jSV5BHH5
ZZcENDqAhEBfpAkZ9+foXOU3AISWMZS7j8573nblH29XFsZ0p82thoEzsigtQ8iy
36lSBKF975e8aoZz7ZK/8wEZaInsGTdkFH4wbwmUGFWtYvcAv0ifCvzk00fC1sh2
DAEGGJnOGyeuMRYa+DdWZ5PdOKI5F4qJTjgm8d9tt3wq8yFJINPRYk4XqZRB/gMr
9vU6rwOnA+Iark8OGvNr+c2dxUhcGKTPOD0Mp4BgpPTnV6knUKSO1wURGXJq9dUu
qgvo+qJoIHZMFwCHHcCk8dna3t8n+qMs6v2JduOQ+GKwV0EDD8FGiG0gBiQQGOW+
rpLTfPN7xOSBKZSqHXi9aR+BI97AGrGA+p8gQWXrCGgCvo96swXJQuBn+RDhMv3R
Ln6IyV91TF6UZqOL32Plzes6zkj6VYKJ/DIQaBBHzS4W/Pgzk+Kj0cr12qj+4bUz
2xakDqQjYALnNuvYEyDoqbGWZpGLwF6hD5b2bulwcNv8sbUewQ1TWVJ3aVuNV9dV
lAgzzt/CHQCKh4K5p/zDzxFMGJkA2+t/EhXYHnhAY4iH+q+NIbOjUXR7X/261iib
/HX1Y8CM2q0POi2fYvyevKuHHZFIjN2FbWjVLbF3b1cs6pxj4kzf37QUvAPwmGbj
EcgbYl0d+bBeRnHbkJRofX96XI39vHOxU7rH5DKjOS7zmdB5AHkhWDELThFL8Gmk
8oZu5NrrfnrkOeMfoyk2FKZ/nC+CbGqczI0/rGtg9BcdrhkYGndb1hI7P6Vktf79
36Z30VoIgODup4KFGVPbK7LFTY2RXNWtMjSxov38bsufWIlj7T5TQTBR9wAOEzVK
EZtXgLPTdaWQl5aprzXepBcOPxaUiIcE1kERCxnzyZNYxxdC/GpQ5MmcZlSF528G
KDblL40V3fLApC41LDWD2eQWPt0uZGDRDrUjlpALtg3TbKoCEGVmulWvUX2ZGK/2
IwxZfCvs8A+VrJWARbxoRiPgypTI4dll3dB7Z8Hpy+d4DYeLDghOiFEuU1Ny0yhe
maRoo/O52bMFqqaVZB1nJ27CuXsCoUFa/rOblh+b2ac=
`protect END_PROTECTED
