`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oq0/+st19ZRkQHy5p7lQmHwk8xlhihp4L6iFv1GY1oirpZS+m3RgTkLS2gbDZSxp
TK85q6G7lq0PnLGIMiGlpI+yqvuX1l1d/4lG90RTgJhC27nRgqKuRBixnY3rbJe4
ZsFjA3fsBkoj4NTkpTrc6oQsROuqS68Xi31bHldR2tLPjk9x4+9U19lM3xt5zEbD
y+f9/Bf6u43Z1kBS4dFOv+ZYQWIY6rUeDECsw7DX0DTtGGowlHMJ2kY7NUb5+dI9
G0aVeB0PezTSsAoZwYcsgSDG2y7VsoV5lx+cZnV0yGQSWHrTEPkCLQfNIqBWrY2B
CzD/dRGbMG3RkvVtpRwyP9QfJrWrDgnW5mVorPux4R0hjR5bGKRH6ON99CK9TlFx
QzkeFPYK1HbR8KyWZ1ACYjsLqhK12M22nsN3iK2/NVuV10zy3IFWQBiJ0Tve4ssL
wNOFIf3KayPzeEB2Uf2wfQ==
`protect END_PROTECTED
