`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zyRprZviLqrUwggEL8YpMKLY67DIt9T/D6/A2HmlL91fJZL4IIQaJAUT1uBYCKuH
fZfRRNSTZiLMlUU4MHC4lNl3/dtMJzSjSftMmWhgPdynDxrVgC4eZUSTRYazHsfT
xQx/KqiVamBvpD915c340fHoZ+qKdR6Us+ajjAMiEGWpUadTsfjD6NGsiT7qAr9U
on3Dm2lwAxT2D/7GfjKURlJJkr0w9rINoAFCXGrKDD70IG1OO1n4+v9qj/oAWcu2
g94lpzf+5wzehokOUA2+DEs9EyDoh9wTM9qC97a5At0ade1xf4FpPstj+6tvxm52
JTT+Z1JgFQWKC2u1gO0gCQ==
`protect END_PROTECTED
