`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iL1kM+KOx1wGi9hQl26R0YtDZJdOUTGW4xLRyMAdm1h1fR4sAiTdNqkBYpCdHy0v
QDzMRYmfujkDazCZAKOeoEEsqP11hAA/lm5/Wi5D8cLa1POpuF3v/ZDTA1eKX34W
P6VQKn/M3dseMtlbnPZQgNeUJQmhMTP1DRQvalFXqqB31pup2O39gxpz9jjEocRy
cBxQJ1IFOn4TJA7oe2JsbFcdKbn5u4Ox9kt75dV72N3hoAksoFtduJRHW+BIesbZ
QsIM0LJ3mqV9ZmC/KdDYMpKhkOkhsD5+OlXxCnSDpZdAGy/Ww/R38gOAjfJFVfOU
nOisKIRSp+/JQAdnwTEcSruZzgttn6wjAyctZKVtPG82TfHBf5vU9IhTHMKYbU8S
iC9GEMWEd26ayY5QmRZNHd7lkdTUPu6/C5pEnGnc0DZ7lD+EROVxp5kWrze3wE5Z
ujMqjg410/qcwrkJJ4x+pQTlY1vvzq8GcPsQ0B6D8MDeClIg8yxaGI6vHCPMcXCo
rLNAZ3ls043SfPlmuvDm7lAIK2M6lfMf4+Dn8B73LfVtKeG47yHRtEVx3XwoY9Ct
ZzFSr62JNqRK0BDK78D79bCK+H56B6qb9IZrmYxRfEzUrzfBKvqVLB7Ve2SuOcPI
+2mdd4+e38pdBx088t32uZjBumAVZCN0GPAy2FbA5mNkoDW34Dgo+AK5Jz+cYcUc
t0AxOSisTZdYy9zx8HODRQ7lCQzvQlX3PJEISvovE2onJCyssV90tTzZ1+LLIv20
tbDrD1s8Jsm530IpWjl4pAUg9SgC67sjsKrwpWGU/bZyJsVv2uiilRHCG/sfGZv8
O5HSbjhLh4zaKFSWQKgddXzdPNDSAVVWpGzlUkFb0HNAImMzru/4eLdd5zFZYXoI
ziVv7KRDiUtEibN8oWxQ76ZLPhE3e1bSf/AXkre5eE8TfPlJo5r1Ij2Px8x2N+hJ
x4UPgLrDBuKrG2/1kpBxN4P9v9juHRQKB3NR1BcW2mMHoMyL9pgRbfk83BPyGay/
S6hntwar3cTA1AN2KYAchKQxRLAIx5ksf1gdUU7q1UGXlre5Zi9hd6gg8jSOWzcI
tyaR/n/G2yLMukaZ7SrVFQ8BNblhS0++66gaoW8sD5ycI6ng8CsVRigbG5NlJN01
DrgTlfNKh49Womiaz1QKlPmbqleTnggMh3LSWLZnzJD/Y7T2ENIe9iKzPCmrTngx
jiZPUlMwE/dKI6aypGlo5k3cwTAbCIGB9Iyva7eA5eGWQrGMHgMq9JshloFlndlL
h6IbZ4HOsmHbNZcyiP4cH+TuqJe3h09dR9EaLpgb+GsKKk80rtrpJMfHClcrL/ip
s4vPIULJ+vKIVcErVWWULx6Wnr1OBTlzELSLYqjqE65m3edyG1GEv6zftfJKqq5S
NuZaqxPsInR/xY3eIUNs10ZBlBhNmQHMDu/+28U4NRLhVKct7c6SP9bMiNsDc5uy
Bt48yLb3rxoPrSCQ4LYzlA==
`protect END_PROTECTED
