`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hYHMoj1Dk2VRUpS7pFA6kyN87wXynyx+ukVRZxaZQeIjLJqRodPLlXer9bKhCeSW
7x/IpUq/pvs3/C/bxZtsy+c0j0fS4AR1aP2M8I5wQnAEiS0jk2LHq2uDTALD7uJz
nQOf9InkhkseZJT1oiE8wx5Ou4iRPJtkDbm4xH/4YmMRjFZtimblq6b632CWnv17
CqlbOs/HeYGdx++qUAu3QcB9HCgxvoZYjCbx8x/57tt92GeQ3u10wTdPH4/nE+4F
OjfFrvChmuZOvxID/eDI/95wm67MvBmI/ZXEI5fdD65sVs/d82PqFdR0Xx4gVUDf
iexVO3CbjsXbt35qUOvS8J2vpLDrSKMH7uuL8etBpp87QwAW8V3kQuM60CyLoF6A
rvZMP/vOqU/og/dKMx1G0UF1g8lyx5bn4uzeZEgn/uD2NhBmiQEMcGFylNZ6Y8j8
q9opOFk/vl/ex5LAGZrCQ9qHQhXQ+qd4d9NwkW4+/Oy1HSTDQtj82reVhlXHlMMq
`protect END_PROTECTED
