`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qY5aneVQHFj6AE4H15EgJssKi+zNouGetTNsUBe8UEffPQvqM2yyDmWVVGSXrNsL
gXJ6AbpC7f4vy+B7k5pZEL0eRDGFRuz6vxxRTE1Ytt7ZhonqgKb9/fN+30IfRwOB
pAO/Anf7qMsQdZVON4w9shm+SeOl0guJvldvhmZpO+c8ADsr2styz9YOes7mS4zP
0G84ojMK5B9a0ChaheJvGRPtDV/k1HoPuTrYNukzHr1ivPHLWTucuYrxF92vXvfy
aHTsHL//AFdQhRe38J0vEpLdxV42KX6KS1IgbL/tG9yjs89+yTMQa7UzALgDSw+n
yXz5DMQvBPIWXYNAjTWDv/NmEoZW114u4YukqVd04KjXvQt/kcBFH72ptyFOBiZv
Xhbn0GHkaRrcrqTkcnzF0g==
`protect END_PROTECTED
