`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8h5OGwuCdqU3qQ6jbp5f6wZlcQSjr7AjmCUUoir9PMDlVFUnE5SERwBLbIX3ZTlj
Aq3IsfZpxIEJGkKbBprJw4LvuAtHx1B9l3SC4y3/hk/Q9hPb3VmzHaL6ImNU6YdH
koXGEUJZ4PXdBQrcEvwXOBm25Y5Gr3vs5ELp96vmTH0iy2EK2qEibSSiq4BDgECW
b/ivUNOwSWduZWFdjHgnggBZe6V4l2BdZiGJUgGym81HhdP8HQyn8pRO7A8gRM+E
`protect END_PROTECTED
