`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BnIDgq20GCFndeM7W57DVoFcL/ekWjLFSZyZZrSxUNB3MyFCDcGAJX7Drx+J42Wz
ks8eR2wxbm4buwJobYqxDT/jWx6PCQAJ094DSqVrCCURiDc4okte4id1QMASvHvX
8JNqiuOylxwedsp6jFD739VZ1K3HVH9F1wkTecvW0oOwon1OIxJ0c6vEDbxdKuR2
Z0BQO6ooqfCdGb3Q3h4pRih89xpR+EFMwqEK/WJMfn0QM8i351e6PUiPbrrAxVrz
1P+iHIASpLtBif+6ukHufkpya2a/JbHtUKmyBKIs1DYUrOXjAK/TZI0DUWvQ+2FD
1uV0qYGWMKbY0Hbxz5UexIdPj9GQrbqRxxO5TUAqiIQ4pVBn6OiU8tP+27LuTfdh
j8RGQA94lODq4LleFZfyu0u6gmK0KD8tmt35t67KzeWIn2GflBbSArx1J0zFUYZn
lluh4KkCBM2U+EfNiaK6UCZu9iPJnJuz9aExb7zIWoq1J7/qkwFx4UW8a2km2RMf
hyYtpiOdXDnvK6Dr/3lqSyIjHl4/oQFvK4VP+s+ANjp8xtxwi2y0V/h+e86JIrQI
ca5Z8oTR3arS9XIZpHZHuQ==
`protect END_PROTECTED
