`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOpshCNwH5dkmY/lvau6+A3l7bLfoKK90B5xf09Rw9ZLQGFbeigOYRYbd+lHLDHD
BrI4vfAM12sWO6Ea+BOnmWhyVirV29/GTRQUmbGMtvoFbwVumJHw4ELoO/Bl9/mc
S4PdM9lo2n2BhW4MZ8BPT14wqB4OlyUl/Szg8Q2iADkOxDK+AIiz31PB5bjdMYPC
NHKvwojtn5MaD7Iu/WDeoZERYl4XhyycUdIbadt52eCh51/U7On/y9KxB60n/fyz
pG9fvFn7kSi3ZtaNUW23uyONvXK8K64SpIi+A7KofSGi6XleBHswqEVgRb0yqAd3
/NqjeNsPSljoFqIE0czBE3EZmuFDltEaE9SSVtO5dNUgbGZKVkg/4UwOZch1asqV
pt+I6OpiW9gLZNZ1u4XalZCXvT/kAuPcLNBGoGBY6HoDb+lk+TsSCouQBzo8Eem/
h5KDM/uWgUQ33qkM4VBxVMyPDSfOfDvVEFoiZha/ZNwn58aWm1r+mfoJdX/oEBWa
MaBRxoFfoIkS1Q5tVPyTN3D1Pnq2mlqPcPTPqXSwjiJMiwigDuXFEtKm61FmwHOi
BKUkGOIQ8Q+VKueXuELOM/zNopXE/Fa+sEBtfjPckOEEGRyqPBGx013P34ntvI7r
OWvWSaU2ZmFQaBthv4scsoHade/lboF3JphCnplgJKeTZXI6rGVZAx3EXzD/urUS
N6tCRSP4oWAvc/nuD7J/p3HS4SaYr1Qx+ZKgMc1S5eU5e4JL4V/lxijBDD1zwCai
Xd/b8RkaOmGYtmlWv6fZUGBeCJoo5lGaJz/QW1nWkiiMMRtGwyoGwYeB3wy+O1F2
LsEJ/kYKd1ZNUU+sv9T1hgIAgXR6R8fLDHRNlPfCvSKPHluOaXSP6NwWBOI7Dcsc
VNc0XajfBMxnW+I8TWtCqDpvz4uWqNbwu6ll9pAAn+Q=
`protect END_PROTECTED
