`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpZOW0AQsrrvy59nLF2/LzAl+vCx15DOGGzEUrFpVi1l5Czf9ty7ukok/R1q1J5i
X8sNQ6TmsubfT6QwPtDbogg+8zHThvMb2ee/nM6ktdgk4Y7w7e9idqAeZIu1+jZc
9+zm0H18s/MMtAXTkx2DfBDc+Eb/+DVPbzJEKZ9BaKSn0F6ZpMLGxaLtCJjLkgsy
02TaDsiAtKEYU+OwCkxLlQaWaSzMcYso4m3nU6GN7JB9/ThoT3p8txwowERgk4cg
P+rY40MhCIMSwH4zQAOEnepo/Degnm9csY/meSoTYFaqd64VXE2NxVMhXaBMwW9E
8U7rOemyvksXiaKMMKABgWMTYR4s5xZOU2zPKTgSVU1Znm1dfMWDfdl1CmKjekc1
whb/x+cMYkznXgZUrkuGJ6q+HTeOTmzwberhb1XZ9GDtULomggS0yovUke7YC9rM
AyJepltvna0RuWz2UXIPpzyCF5RggRMj2WqxIy4AdRMwyyCMIBLhr8AmPXfJUTrU
WDzCHEsRlKPePdyntgMoEyHyoQXPtqWOObTo9TxWZl/WzRmZv9pkAkuqgS1oKbps
eZ8qGRF5JLXyjCtE8E9n2+I/yIoEbcthH8nBLMAV2t7bs7pq6oGYrf7vTkT6XQSf
lXUA4loDL/irbXfzXv5aRAn6bHe3JL78iH4aN4LNhdQ6J0KkaNFQ6VfAxclL69m1
kPHBruyLvmqA0VrC2XK5QgXpdr5Ze7UM0q0qZTI89tw=
`protect END_PROTECTED
