`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rXzkx1AGkrc2/REpCw4lqv1OSkQPo96Zx44cLWvBkaUcGnL3/uJXNDZMzvAuY80G
8dWn5UZyQktKp8IMo0aZuchkMa67ZQDq00My3lXeD9nirCbr2PvhPe+pq2p5u1SY
nA4oJhuJVhA8HZyFtNk4KSwKaXo9ugt9yLruxZPy5Om3xoJ0Z6WNClDJTYYlc9Fw
S/xi3d8wCTYpiNnrrVK29h6Ee9puyCWCUKyvz2GkMAAKoaXNKnjT6CLBkPrV7kr7
klASYeEgFaaft7uB3DwRDN4m6i7ZwiISoBSOdunA+0qJ9suu0YquPg6dIuWSO3qX
ZSYkWiz0HwVjdwfdEZnX+lJuWiMtPF7SfgMDQJama6Uhrnqe7JjHhg2W89xZ6fib
jXhtZc7hGELCY8ugxwnF1nM9r9H9Pnv9nJo2xnAJ4vmnXDL0xhM0vCamNdRNQiRT
VVVcn5hxgfNX20J9m4jvM5dEVWf6KvhW7dl05PsmlSzD2TrMJIcGN2TKXL0aiGpR
aXOQ9jvH85oBGVZj0U/0rF9zSclWr+6iLo+Hrqh7+Xj1NWg64WmGXs+1hjAOGopw
27bBSPtflr+2Nc6rhvuxGzurHSNC7WWNi6VlG3PgVSR6C4wUXOVkLajpazvdcnH5
EvNdGMJCnqOaxl1+P4+VRgREiIUknzRp7AFI2VmJlA6XopIK/uBstj/Ra0VfbKOp
6d/X1cTSjHl3VgjCh9Fjv15UwGPDBA+nk4TykIh2brlZtjbOBxjVVFSXlBsyMd/V
VX6dqFoq9tVPEJZmfmSzOr2Iyrax5+rLX6A2xkBkbjvBeHqi6OZY+Lcr3b9u9N9A
GiChqXTwKfa4S7pDnZ9ncwUOfRM4JVijYOBZbzdEhaHos7Md1LEu2jxIQWOZDXeY
dbNZ5pxuvLf1KP+AWmEN1ObfON4I1OQZTYyYz+bhk5op1iYnl7GAA/GH1+Gl5yjV
8zXrU8vxGIfHExgV7Ry1t6yrPYz9s/uTef61+mbYmNNb2ulnomSOzmT71Qc8oozW
8ftMhd2Mlcbc4y6cH4oMJg7qEKWGybBZyXy75MhCQmIxAofdrJXlnpMhm8fzCPk/
99my9oyo4kbTNYuKz6z3MNr74Wtl37DGIbHPS822T52JIgF3L1BY/oy2Rl6V0IE6
h+dT4e7JMLafqhEKBnQM6dZgHGUL1TP4qWXmnOyRkMUkjiXJaAEbf0d69sZPlJBE
IFLC4233SgpBfirq7vTI4fI7GnYirg4suVL8oL1iPmrelyg4P+Mmi2FygIQjxz0D
4VmZzWkfB/pCdn2yXNzs/Bl9tsc0RWTvGH1kB6lLkalk1chp6OD9Ledyvg9RuWKz
CEedS6byL9+f9EWCEqow1q/7mKgM13RYfnuKAuMyA9JeWVSBxWkzeksSHv18c5Ne
PN8vyo6VxqH75AR1M4fAMH3VllsbmhVkb4h7kUJzRZdEYMTAxc3wCqJOY8E58fe6
/e3QW81HnTs5ofdnpJl9xzb7mVVfM/1G1/59MjGbmx6YX3klg7jOXrWXlih0TXGz
5UEhyCmEC6lBcU1v3iISdpBxsQJWgptQS8OKlZF01NQlv85NeS8gWXuctfeWRc07
NA4JlItyUddKMCKLgKhyAkoIq8kJBMVF1ZFMGTU1iiXlpJg1QJjZMBMZUj/PaEZD
vZFQddMie+FWyvPeTsoQdS0QynJ/+jJnMhK58o0SHpG4jRu0WCET0/m8IpPC0Zqe
pzKROJY8N0ktE7M8EG9wjW7qkmy/qdYulJH3mb6uCuVC5jT+0qlY3mEmuKqv2kLs
zCq06XQK9C2f2xuIbDvq5J54ej+Y3KyK+BCQDgmi7B+2/V4g/JWF2wv8qLGAkb5G
ZOjoGmoKq4WWxy/ys50Kiw4QL05uSl93hEZ4BDq9zgSE0Y+oUxuZduAqzbt/rxnT
ALRZe+UIb7I3AATVfVdfKQ04dQSMZbNWrNZ3DT8S+37tFD2TdB2Xwx77aCB4qV7V
asM/vGd+X0xzVUPmtW1o9/ddNbkHCtAEEw5r/PvHeMiNEQE02IYkTJry4hpK+gwr
X4Gw+cg5L0cFVGBYDPVxweBV7SmuDOtWbVbqVzprlnri/cx26dDPujYv1abiMhSm
nPXzFXXFoOOZux1f4k1AoxO6+RYR/NzR2YXOatZFAIhGbdeD8ExB/ugUkKZOG16i
SrZnTiDmocj/8iRq9akwWcjEfk6kFbZbhKnrxt579F4RJBezJRM/KPMXMP80m33/
ZduTxjTMys+MKvrsLEK6eyFY/H6LkwFC+UxSVu+4HrsxSkxgnfcOKaFu8YmZpMFL
fIeLuJgkoepFpZxZZWUf1ynutVjAA+Vu/SHB/MjF/6bXvn+BNve7mcZbrGI6Lwky
BhN9+CrZWlFYeAY9LPcBaKq2PcdODL3/6pk6hvqPNZs89o1UrSm51NrUDMaJmaqK
yyZa1u6t/s87vDRihV58GggQpiXJoMVfJpImU2ZU4nGvFb2G8ziKzmrRCaXQ5Uwd
zfaU+q4C709giM0alu5yfNFsNdH0+Ubq9Vq97UuvH2XvIIscvNJLVFKB1w9z8Nl9
nWy49ZiVsws4FP9co6R1DQaDSWZ+wDwt1JNS6mFZDp+5zhzTIkJ0IagV++F7kaRO
20DHhSYTZ6YIuLchsFI9pFsXt/QV6KXbAeUZ3+OJnJs2T6iCKRcm/3vYllxw6ssl
1Th8xma406K8sOxCBwpzNJl2TJVBhCxW50QQt0106NklalDUtj2/rVceKNHGElyj
bmJA5YJ+GJK39WZLZlV6Gbp2nS+kNEeoMYQFKOzlpcM+VgKNk7PaSJp2miRUNoqB
/hxj/FY/w7flHTm8zw+jH3538hIlWmUdOjdLsGow7Tbim8MspRD1dme/M3oVvBB/
4gs0LuVB4uX5EkNqfuxLtqV3OjsjATl6Z8HDKUcgqMleU+CXpCa/X1qF3tfNvQqI
/it8fznATWtwXlDrm9+WZheoME1jZq40D75BcMn9pjaCFT82ZD1QC7KPBQPNXhL0
Omu9jel6PyBXxiL9unB6ZlNUPmoIV8iMlwskrtrQKYMXH9qMPxmoUoWslT8y+6v6
/o5MwT6cjd1+gcwYSB61p3bVLKmXBOAjWICZG2ibXQx+fCRRvgn68SgJkYgUwmea
zJA+agddwvonMcBOyyl7NWzqspFS0tDF8smy9/lfmyh5JbZpKiyCBo0gr0ZaFuym
`protect END_PROTECTED
