`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISGw5+oPpJNRqBXyFqJtFsgZNGtjKGKacnOi9/gP0aIgRowhfqguxRcsDV6pJLrd
611rqSorQfU0o82mwiFtMZvCxTEN/f6RjN+fg1rmStKjA40wiaQlGKR8b8z0nFsE
P5Q+SLLoFwKQcdZCBk5jeVExU9N9U0+XuCXDv6a3GUD30Q0oH1yckmgtfL5F3suh
Qe33XptRTXCAf+ypesTly30ns4Rdlbl5VHeJG314dpTmORouA09M2cmQOMTx66Nb
Nj6u5VGMvaSMDsF1yUZfzCg81/pcfULJjp6k/oPxqY620uV4f+3AubaSxTDPG/X2
GcSBS/EQFyER1Gd1FQhR2g==
`protect END_PROTECTED
