`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLdoWN3ULdA2ScMAHZcK8ZYfx5EqJJ/lvr+/zM+WTKwa63XJH3jhQHhmGJTr4x4p
A2KRG0rTGGZKYrUdGVI6vB2yTvY7D3bna18NIRhk5QGmFLVFWdsh7goarCU9lmus
YRqUgD/8rqI1LmNgZWqv/bHeX3Oy7p2OMphDf4hNZD6yjCuFkgQx2HW2WEH7Ws7P
AZCFkaJGbX5RsPux+KzkqFv2g5aCosyfZ/7HpTMeDCR4ipIN7iVF/hLhv8B5lMMt
G0rv+JnyKI5Q63sIqEBzfMzGflFPNZ8Lld4SxefrPJ2SsYL7vuE8vozqjWGWUQf7
SQkrW+cZrGz2CGWFjjtaZFDAquSEF1UW50F9RTxl4tWzxGUgqI/AbR1w+RTsnf2W
G+QPxHncEXvWBLyPxf6TVFbYphvcW9J4uPhmXp9OYjqe7rm12AgX9WiDNSNHwYd9
amDvF0XkJ2d3F7Mvz3uJHHn3sgm/FxjS1Zv14fWAhH4xWQfFR+G94Rt9UzOnubTD
MP3Lgspdb1pps92cZg18DzVJ31vyvRnNyt62yZOC3gI4ikUsdXre3rjDAwUgZMJk
vYpCjWGkJeV5CWuAQ18bPnurrHkMvZBun3fJqYC1HIB+ov8lceTN43E+a2EdqJjf
DfE5Ft2IvuokMJvpp78NkBtVKauUHdImvTbekSos9wxxQ/Cy+GG5ulVQpyTzU+wI
tjb5yRhfmeIDRQaoiM6ups0qygfq7xhgwIMMacw7IzWiQ494IiPoQVtzzLquYmNc
f5JxCy9xXb1cID73EfGXScqWurMW/fBP4z1L64rOfL0/ODgfST771bNfdJwgFSd1
ASq3bZY78AISHNx9rX2eSItFVo4ZFyq+6me0W9ny3DDO2dTLi551vLiYS4M6Mn0C
KAkklTzwNXdxwNRBjH5RIzyI287LjyGIAXwqAnjXPUbK+6cmlkTLQAwFMHCrUXgU
0BNBhld9cnjfY8ow0fLxjf9YhwGEt6pK1vxzvwvnqiHgSH1z/oUKxunddFBW2gX5
oaxB1isiRv/VWVxQ3AnrQmNQA+v8Ti0XfAQA+dG/oY4=
`protect END_PROTECTED
