`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMRaiLngVEvCVmSir9bATYfKALHeXJ/crnKJde11bwWt8lCbiNS5WFR1jpQX/JbC
ZAYYV8aeDJzOEsCQ+DJx5+ZVlgZVBrmflMeQ3ukv65sHkcoyOFObUb4bZMnmO3hO
w+0bza9S+xATeMW6/9097N7tQnY6sXgDqc18wSfwe15C8PQ2F92ez1ShtxxHj3No
3HhJLbhqzgAE4xL+nCePWYomt+IbBqMINXSqWEl2kooqIDccRyRpKST8qnk0XAtu
uYB0DFYPrHkp0wojGUzLhU9E0HrvsGGkIcYOJQwpf6s=
`protect END_PROTECTED
