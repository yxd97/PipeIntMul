`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eG/s0i6O+d7QcMZsA9Ez5K9Ohee1+O6TdcxvCauuPCHKD00nV4637uFv864BvHTb
ejPBpjzkDnqAuGuXWGZJlbqEVxjAxTfL02pkTF27yX+bEWqxOuRfNIXTw57FulDA
0NyVXSmVCoQ3LGGw6TSL21w3r2KTO6v4C+gByzX472IKN6ewvjKrxi0aOcDy6I86
CvnrhIAR74g6G0VOmcty6gmyZ/j/ZPRmcCVp8iACEZgcglETGtSkswC2CMy0uyjp
ju0hXKunja2ecbXAxjdLW437DCswvKcA/KJAYljsG4i/i+wPpOQ5tn3J8jtYJYpw
ppwo2s1/9uyUZ2ArfBiNAZMZGxI7l1ls2RuCvzNl2I0Qtljdt878vn91cyio1gEO
kTCxSo0N/iZrFCtP2pfGemmYiiK+IOUxHr8FSerhGtMagkwtikS+LYKqzbVnlgKa
lmRbbRnrC2Hzo2X2XvGhD12tYH5PMLDdh59DYpB1iLhaW2exS/bcjePHBL2sBLy9
vuh8ZnHAi7E4kXULAMNeS2QH0eyLu3OZ8/nrxxrBo5W2khO4+B9gKbDQqHcrtfat
9UX3UlmG35Eu//ED0JCc1E34bUUd1ACg6fG1U14JyieJF12zXnPaLBrfvWeR23zq
bwgJ1djtuAYv7+iBrdxS0jeJOVi9iu2IlCn9LjSyhQuMs9jhEY6I2qoJJRWTBs2n
HaOqneXYiBHm+9xp2ZfsCvHdN6P775swUnhXF3g+Ygr7lZE/nMnWd2vP/O+tncYz
qOFqhnGOztWyqnlAFyEfZ2oxjXVSoSnUlxrGIaB6dvzDClcwvngmPUxnEdzYYjhK
w/wC0+Y4fav4gMBeQnjikD/Byjh2MObe2wKibzolIi4oOYv4iCNojqsYORftE1KX
8w3vGenkk5xtQ3lsJAoiIiWk5RUuTltTIlluhKk0AX0/2jF/niBiZI6isWezQlg9
6tf/jSTfjIfRvMTjlQmQ7aliJpvsaofKl3l5tfollcBDbq6IotdQhDLoVsLUQsEM
IIQbGmVlKMIqL5EJ2+grRwSFOXNl2hQI8Lf8cX+6pHcePgsR+iR+QL3LK2uhWf57
lo2vh3dFrxqW6p/JMh0ZdelHK6F76ukM2F8P3l4YV2LnpWU6/Z5PUfl13N0Pxw0z
ioSdi/VbD037XpapDV4jHLtSYBxvMlJUlKH68qlo5/V+aSJ2IZqu3Z4anPfSXzPg
e3rmlrZH0/nT0roh/bwzuB63/XfZYTd30bffB6OXZtwFZ8I59bA17NsEbHLfcD8x
`protect END_PROTECTED
