`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7hpkk5Lk975YDd5HCyZpaL5noLumQIZ0+PdSU2q5fWazRSOjoT/nO7gOPeAAt8b4
9BDmuMZz8fODzxWIhc48ULXAofryd1zF2nLu/2KnJf8/sASDByKZKeFT9EowD4i1
Ltt/yrEXEkdUTLqIDBus/3Mms+AjPxDIa2tlkh1D8t42mrMkjzK2nEcwX2uVdoyz
9C7RaAUN3V57ZvCgAjLpTP6blzoUEiVCM1Wl5A1YESSvAqgYbKcm96hZbPfM6Jzv
0Fj17r4InBfwvPLdc9JF9UJwsVt1LdWX0GHQIOpApwkifxaU/oiHMGcOfeUe5wte
IkFbKazWsmB1RTm6faDrNNwXODcVctu1Huiu799/sYYycTjzseBx1jw2AHpnJ7qk
H6RdWpWFV2mOQ061KdV2s5Y6XyOcCskZP6rRBFCGxX4=
`protect END_PROTECTED
