`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uft+QdSxL1At2aI0VgAbAoAolOMpRCDUCZfQU37OULGytaFYnPwqCIhdCuyF9xrS
tzccGvh0hoZKfffS+cBTr9HolmAGzzAFC0FLiZJ2V47x9f1LST1LYxqXTiZ/lPQg
X+0U1qZBDaZpEodcw4e1pTOh9b4gMm3GKUATd/ohYc0q3yNFYuZinGcAajSHQw+F
HgxdyTk56D5zU8Kzd6rLQCgsl5vd8A/0lO+QuSvm1KhIdht9wtM45GxpZxFmLlEK
py98PBxTX4kt26okATzp9JkBQqNblHrKfUOlOwu+IkGq4hmOqXU10beElX2uIM0d
dj4JlkAQmP3zSdnu7eE2aqX50ARP3H3qdpI1s+YZtGoV4xoG5FhXoliTRgOBb0iW
tVR/UKz3B8vCMcfhDtjHds9xFG7ZIzyN7sEOQJPH1qAPISoPavhyeBfWC8IdpKfh
xdVFErdA6yEsW7I+ypimJcE6JOKBhGt0tU31t2ci1b0k5mAXDk23ThBB/m/7O19H
bw+/fBzS0KTdOHvlAJQdvjfeXPo/H8fBgnBIaho99bIOCriztS0vNH8Hg3pzkh8v
yklP4ycZp8/hl4izWE08BO/c95K0wFOrBMp8zvhKiG/kxs3SYALX4v42HUwt9ktl
YZ727i+9GRAdtbl0wBsWKw==
`protect END_PROTECTED
