`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eb2Z6XD5fbYGqaruEKO0c6mvKRDGacD6kk28/O1vrB7uzyBf10JuMUL9/3tL9YuR
zXkroZ3Mdv04kM/VuBqIYVbWLV++JD0jIhcA3ovHUTybYlxEWujNMOXqIi/UiSJV
5769HIyedr5yiA/VQZxLje1QaBizX1V75+b7qooGsXAjC0ku2xqjtngU6kNOKW02
s3IgzC5vU9tlRc5do0ns9RkK5Ggri7/3w10buIpQ8uJku1ITZb7YO1lBSP5Yej63
IVsHcK59E5tw3umDIBh0Riknb+VXmqKSyPMYucq+mXHnWt/opgq8mfavGd3QU5xe
DYXeHwcBjvorY1JgxsR4KRi8okUDVcsWn0FxGFYjw5+QjFDQEvl0Az2YhDcRKtDE
FTAf18XUEJfJBtb6dUzBfdAxD/7M9KWalpO0CCmEmkGCG3Caliya5Xex8pzZ18go
b7gHVi5oOMTuUxCJZIcN27uPMBeQoNsyjLF3xoDYCWDrQl/nOPgKWxEZhfhByiz3
2NOQtVB/dVBWw8Sw8IWBFc3CpFP3mqVr6Rp3EDct8X/BqU0L9G9sdNImqNEVN69F
37boK6ftVJbuq0p3/GTXWVUct044IsGeWQFO5xlPaliK173AZ5fBxSqCCz/NuzlK
hmdep8NvLlMcRuneJvKDdsqXKEpP01t+0pje5r9D97FaMSnw9+SV+PCVXn0cSCTu
Q2C4ypMdkP/RXupHbca1i+zzij/GqybM+FByEe2Mrbk7Jg7YPvSz4K3uStGYgvti
B9PJkcIV2+hoUE+Hfh2eByo5sGjFhKv+vGV4hghOTIuoLunAGbtDVqsKWraXTN3K
WguRKBZiJuOyfQF8GoI924z7GYyef2DidpVZbqB3eZfriFWwuvOmdMG5k1bg1mrD
3PdiMMtUemm5hwDzspB9ZH3RuSqlkTEfMMWM+oqHlEeUi0tah44aL08/ZKQUq+Mh
707XgtSIXEHF0u43M64McI8+hw7oqBza7yTZYebGLUX2eDX0ARdqB4d6fP6rIuGp
4NhD2vnSqKo99XyFdSXYUitD90wAphYVPJAn/4NpHfblREn8MvEObKMlCpez+UrW
iNgGOcz99gVkhuHtpsAzmksL/KIUY08AO4XYBZPYvyiBypN6/ErKhEtMj3Nm67Sh
vX7BvpIphu4Aagg/JRex/DSBHvQMenWAleBE0PqVp10WBWBiI2zScvRUlnisZTpd
y+Ra5IfWopZMWAVXK4J2AiXPo5cCZZ7FQeCimAp1ThrWF+O+WDOJDJCOi5xKYncI
grs4ClLbVWj+zvOqf5GQkyQik7Rxqoo7MOefB/EQ4nocO5UzXR8Sjl1Rllaih5fn
L2HqAFKmyR3bQ6JLFWuL9E7rIxoHoypbaoBah0vqoSt/yMUDttqZq5GmGf8g/zO/
8uueOmWTWYJ52YAmuad5bJ81RCl0DLhTQ4Dr7g1syZqrRs3KyIU4DR9D/QSQbM5u
rRFFu0qkvUw0nfnBKHvkKETjb+qf9tyqq4UNjzoOx0jAempZWHzyj4fu3CJ0snjm
1S8m/nVU7Novntv3k6HiHYQgiSK6m98ZhI9ZCQHD5lpzbdMxQgZdPeB44ue8syon
GgcVquR3vx3VxlMX4EOI7tivsiJPu1qyF2qgDTIuVXmP9VcQiSRWPNBujubZkU8B
4h4JhPpMf4mgmGKL3KmOWMFAh7h5LCUGrPJyvliXXg1UB2kFT9CRLi2dEH79p3ZM
oe7d2G6jmYTbwMlBDiM+FtYtzaSXCZL63OqNJvaLKaOlc7Or6jkkSBujUAFmStTe
btQKKByKUhxqhbVN6RPk1B97O4feBhNDAow5UAGqqxaGqNlUndrjMf8VAKNFxV6m
PdGlW5fH0OM9F9EMDenThWYCiuSidy/q2A185Xay+9Trc7l2VPcXC12obgiDjyl2
RDFngETIaVevT2QwJGqKYDI6OdUwykJDr1uRRH64pgO0BY4sRR9U7oZNzWNgOyqr
e8POeckkqsDmuV3BFFEpuovo3VPL1NUTt2K3jC1zuUjEND6/V3hNDakcMf3MVdbN
WIXCZW8+6xuHQ7nqa4uGFkA4yw5fE15F68oj2EHCPDsGKJFmHgtSoD4rSG1xQ1Wj
pe1M8wd+z/3LpN6LmjZr8wnvUn+/Ytndk4uVCX+NkGdm8YGw2M5BHtc78K9eIVuC
hZKn6dGi5Gg/5NI6OQofAA6kyNXtCd3Wsk4fly1mbqM3oYX8rXL7S0ugwFrg9246
JOIdQ5T+PZAJE7mjOfMd1SeuQD18hBYTNuK5T9/ALf3KxKFCxaaWqB0QUoMXxpj4
hLiwlcXP91+P0kyFC+yHD9yjcWeF3ag4BBFi5HkN5wEkrfZo1mO1m1Ri73E++eQR
k4XYQh8FqO27jOA/gdXfG4fCuaHTtCUf744YBPOOIMLyQik1+50d33/nIV75HWs6
XCPAyrZGS1UgJTU0JhXnqY6as2Py2ph3YIK0JfC6vcs8tk/CvdSO5XSMtbpM9qoL
LXsNpuAe27ufLjhdeXp1ZQMPiLwnJ4EhiQu068Toc1fbbZXI0ZmoYp+QK8o7EIOb
K28jOyM97N1UwM70/EvnZv2qU/Ys1ZYKK4506ZU9p/DRbTF+/KlF3WIDw4Dpcxj4
ZPepDTE3T4komx1NV88EbXR/FTwcg81caP1TLsa8uQ6mLsv6tPYUleXRaLZwbzmR
eyvzKC2faBiHjVyuS+SpRnT1utVGWBbU1EWQ/YAcw0OAOiqvYscOgLW0W/q83QJ1
HtDUSuS5TC2N7H4BibhNP1Z+rIQNUImnNBB/LmAMW1gH/jnFSBY8JmtCzz1JoQiJ
OoX82ZD3v0pR623NVFe5lEKc26HnW43DZQFVQm4LGcwzBiBPLb0gAe73aiPGTL64
0juSj41WtGYtaGEQrozKkqFmNmQoX12lvzXRcas8zidxmACGN/TvOFWpCgY+NJVb
nuGuTOlapf3O+vYDZZjdz9yeBq71G6FqKBIZhSJGoTCw7KMQ4RqhsSS2lel9r3jB
cN2rDQwQhPUqez7NVpTRh1hmxa/qYzMTS0hohogJnWWqGBi9l1PkLoQNoRo+xTOj
bry/gTrjPuXEGvYtDFV3NCIvkCe9kSaCGacGsLdVyvo7TXIJ6UpOWXqFtv9ZYzCT
PQqDvbA7cxaKm6z2ZuAL1iz8kAI6k+xBfh8rrKe5s09q4wChimHpREfpLFE/9lap
XiYtQSf8hSno90Q70NiVagyWSkWdkrqAKlilJE3PtO+EYsYstRVHxDUog9Qt9oKd
WNxUZWog1H+GdHOuahh+1VTBvLgREGTnSG5bxwh5IMWJdvO4MfYiq/gca30cDWm3
T34e+2QfDm2m/jQuX9llvUHJ7MycELMp50TaQJnftkcEctN0/5v7BXacADmQ07dw
`protect END_PROTECTED
