`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AGF4qduNM1qv2IhA5pUaB18SKTAdaswEd74k5Nys5eb/TB5uX0q8IU7yooQx+Grw
0aFb4r/PHJhbSv9QG2KaFz9rm0q1wEXCln5dcplgyhsfy/CoZ9lYBnnXFO3GKSNb
pIg0lgL/wK9D9yVRI98Ot8LO4nPPF75WMsbiVD1ux2ZKRJpipufwGwv73q5DVbNi
69ykXsIRN6nOxvu/KpX0Yj2H8QZOxrz0IEecYH/jPPg/PfZmI2NfxXKEzqZQDiRS
8y3DX7B1auJY9J5wmq9aDeCJFwIfudIw2oE7TzfmGeOw0sYIVa8Mp0eBBngIqZ3M
OiVVX00beRQ+2Zvdd0YtmUJAzd9SC7Rph6IZVcTR/hZSOqLTVKZ7xnLVF3REpCTw
cT+0yogFrFZx2uNu3Y6RFptxC29BCV4e8pyCh3vXnjPHOyqK1Y8kiW4MUpeoUlxI
xpqSAh5jBQCsVn8bwySsft2kN+v7KbLMT8Kb8FsXirftnjpnMrULYvVmH2GcKlj7
X0h5MouT+5GDEmWxvNdZbc/WyheTWDuKqb540+5Gr1cDUTcGwX8Oude6dgnZBER1
5Vnq19BChkF7JJtgxDDltdHbHiZjP56+q4J+RLX/YaHHuO4jDmvgcUmvcQ7FW5CK
Qmk+DlJEDxBfDFLuTU45Ovd8UYZRDuiWGBKxnFvodtohVIak9QyK8MLlNAdpbZeo
InbNsGDPWtzG1XAWNgJGXZZ4cs4liCgjLAXV1ghf8w23uJw7w2eZCMM4UyrkLTyd
aDEXkmo3C9tqsgUGvNlhX/i7v3tMsqf/GS7MaxizNFWTJR8NG9Xs70N/8pJrekh/
ndiqEIwGQNIWUbZed7XAGqb4anKVXnZsZWoEn4z9rvSbcB9HPKU860D34gSlhL6A
mkeVcX5g+Ub23GOl4g0H03d+U9gTh5ZlMqL4r0AKipGznTYso8Njoh6SS86Cxln6
BMjRpY+Z9K6EntwtMWWavrAeRzxX1AkAYC+tE68zn4b77hXy6fx4N5c78zs4DM+W
S45LqkFamwFJ7MEiKxvsZ8BvJXmSFyJICIJ9Pzf1Vs5ige5yW5X6N1ViFhySyPLh
V1Se6/bVrr2jsKcVEe0ev2alJlnS7Nrix3hcehrUDuyYjodpjrEKM1dgJyMAKngU
`protect END_PROTECTED
