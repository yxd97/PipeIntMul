`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MVBk+NcEg0QyGXd+Owjtr9ULe6G5MswxBEOG3CI4v7Zjc020RmYob9BqJobqzC2J
AEaAlol10VTXO3F6LTCYqXaQrJW2s/SBqQIzboISycA6iVaLq9yyuVANlT32k1IV
53w1niJ2R391psyzrJyZXBDArgz5g9yAn1ukpO/89tVPdDZBRMClwpGYT760MyAg
wXp0C2I2vmqG3mlf/fOrIAvZB0mvwK267gSf4Q2pDfFypidN2CNmOJPrN/ATtUyY
3d5mFfjBPFi5JfMJ33sEjRa1V72CSYHqm7woLyX72ocuxCex8sLu2+m/UBaMSTKU
ljnzRYjXFhlF363n4DRdrkV0VrKh8WJcG/DDDtnPbe8L8pzvBt3wYbueTbXPqTsu
yRj+fkJmTLXJWHYegWCWoySg4lKpdeqh9uFRMd+/q2psxEGP7rX9tW5XOpZpQusO
MvF6M5hFJXTHPIBssNKXFYkIY6QkeZn5OUScYjIAbBJVt2xH7S3PFY/HUaMiQbxT
8MUAa2QM+3SC676Q86XZ0GaP903870zF24VgFFMA6xlm7QsYNWkwZWSu1jft2PtH
IqkEcylGM9q6xP1L2SAAWYdcE9sIB7QJ4v8LlQx+PHmzYe1Bgk36yFn5OkssTV6r
dLhEzHxkUneek3msdpBeTR31oAA5fwMMbqzaJ2a0vOYy1kH3CVTI1LAutoZSTxqA
JeC8ozWayl+Lp+WNTzBQLPTVyaFGMiIgoyR3UniC+83VDlv1PxWwCsCzvMXFtXc+
y7dD5iySooAMbCJd9GQk14G5vaSYAyiVU5Z6w51SzHdAiu6JrEnL2uPrgggOsQtK
K/KRvvekmoAqZIidyjzwVxmm6mbVZkHJvfvCC2I1XtMGcDrrDpI4BL3fqj1k+vYl
GbRNJj0kRdCwrMvR0NqacQ==
`protect END_PROTECTED
