`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+8ZP7p+LKCajNExOjak1EtQE/d0j5NlvlY8ZaaAc9JplDhIQRzPcwnBR+sFeeDD
5Mgqy5tZIMMCMm0Y2rcGwgigRq7LA9MUjU4VTW1oOyD4nmIdgexKfb1TzSxY50Si
tLk+RpkblOm4WV8sdszRquamUMHgEyR4R1W01yGOZDrqPoeY/bWBw3peSNT9+wkE
0NwBZYIFCW22FFo5/iYc5hvsrEn74Sz90PMP6ckLiyDK8cIKr8DkNaCrfG12PanY
G3XJNcDAJXTjOlIJz35JDNQky0brH1R5RYSXKhy7+UX9wnBr6p49SKNipyoa+99P
BCUbzbI7isxWCvLZ7tW/sxghyPJ6PfgdGuv9ZCDbRVGjIVa2g0lAjH+sA7loaIIG
KpkgwESmBBX2XP6He7EC1DJYirkx8pTmnz7Cqz3fl5ohXRlnCFmrQwY+EvGTeelt
A6fIEeK7FBlUEqgsz+MLyVXc9e4Mbw1Ixnq9O9z0Io2AOmCpg1h7VA/ImfkKqyW+
0KXbIMkmZtVhVF6LKxhtNFkBjrI1rkgfcRzW/KzMLMnLkRXY8+HwA1on4GvNKKNr
4gK+gfg/UEBW64jg7hQVXgKsCcPznyyXY5OLQUxfftHlm416MbOivZgywtmcKfF6
0VFiZV2ttqw3RwNNpocFqQ==
`protect END_PROTECTED
