`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bPdUuHDgr2HCzzH30F7C1J8JWYC86RyedvMD4p84l0OGXHaS9iuqjtmJ+2enId9
3R4WVorQuIxgMz+VdkJM3riKrAVH+JqJ5tx7av5cIIk5nD4bHqsWWrViKVWlQx5o
FdcUWgf+1EXi7DZ7JukR79eTih+Cf6kpdoT9uvEosqrJWdj+HHmzHulsxjQ/1dKi
FKsRJ3lhRvfeSR9r9s5iIc1M/GjDDSq0qN0mfa2oftepoiwPs+nv8qdqnUaveLm2
xvsr8S2krzvGJxQM8jPdGStxwgsFM111bUizu9LOaBc4+PG82G6RKpJxI/3/Ai6v
tlprn/keKpuXvh0COJIz5JRJCEQO+M4k6ZO3xIYu1UmMaW45PMT9Auqw7OEk2d3o
7Rkn6a6R9MgDpGl0Fz3m8UPq/nlMDMEKHtVKQeXE5JeRkmCZn8U0EnNloAUU4L1L
yi87lI7uEPQ+/kkGSG90scfN1tqxw6gdYn1uLjjl/ZH+xEQWXUtXQrvTj1bj9Ul3
OUpcUFhBAVRU/DemsRF1zUeFQd5QySLCAv1LaStOIS1UmpDoRf3CGctGOPDYbMtg
deuWP6SC9ndYkIVI1RDSbg==
`protect END_PROTECTED
