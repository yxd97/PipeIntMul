`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kf3QUKwLLdKeaUjHyLc474CmNio8hIIKsEzqFRLOjmIsT58ftRbTgbPu5dz6j2gX
mNiDJ385YnrAPhIUyMeJpUnABg3URlXHsvdrZSLqY91Zrqc0crv542G2C0jwv3xU
CZ7TuJ2iGKIEpzWhmPJgLDYPNJos6OStfy0m+KEpT7rvqvgrSvj+Lrhd68KmsCnX
iRV/93YYw4RquEwDs4R9Ivtgw5ckiU6olIZEl35uxPf4uk2LbcuK6SYXTDpsJunW
wdyoQr79/fhq6plbhO6xGTeJoMLYI6C42V6Jb5q3QSaSlT0Xw9vos3F8We/a6uHr
`protect END_PROTECTED
