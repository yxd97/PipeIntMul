`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
llTRhzKnfTYZ3UOpl8i4jhUEpS29G0ObcZwsZ48/Hl9cy3TNsw9DDJfpCFf/lysI
mTsENFVeyyCdBGJbSQwWM11uhKW9Mo+qQU0QMiuJF8XoY+X8F9bQDUYyN4drKE8b
GxhqHj15TaVXjs+FUYFwvX0k3LZREiyBNCOuBBUXrQejiFE2bRuKmW344BrHhX6p
fk3MK0eqVai2GLwiq/9OR4lYtKvBydqYUXDjxvxjWCUJa7yQnKrkfDHJedTApAwe
M9WMndJLeALVMxmoW7Y3Qg/Y6YIs6I36C3GOlvBKpByWYkF0x+1Or7I6r440P8jh
gYZdR57Y+01By519AK/GYx45KAktN1dxK3OQpyR1CNeulKmAohZynJ+267/9zR7s
iXAknFmB4z29xuzGnpQtkFMIuIBseBtOJWZtW4HkScQOGViLi5MDHmVkoYuDNET8
69kZAqM0wHZcPVVNUgtInPj8BMJfp3BE0ukrraU1C424kG58NffRGxQK0JoWS07l
2lpQemtVKvIYLhUW+1vgcLrEl1OyvjiTlYhipPCTxv+fq7m4ZZcWnpT7xGzuqKGb
+IvJae02UvSU7knglb/Yg73D5dXSfqU43HEe2McpSihlJkiLL/LowwEcTNiTw1Kq
FBFy9y8h16DnvxxH4+QQkkNw88PMSazLp7BhXQZi0ynpVvBfo5iGF12+QCIcBogL
pmdoP81okc9Lg3nbBRrR2olyMXQLVeKv9Qh1P29MtcLgTQxy5mhna6Dy9GcNmdoR
J2A8Zbp1RH9eqe5YlNIqUA==
`protect END_PROTECTED
