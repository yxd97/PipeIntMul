`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
etT2D6JckyvvhB/PHo13iW/qiT5WPCQcnfyReZghUZzXFQ3GuKnLCpRTukej/gWW
C6/4/u6xSD5dMujh8XQqObsq+TZBxSzmLHVc8C/ZGHdvHNTCzTwtQvNona9lvy0S
D0gIV+V1EB10irsSbmot+w78uqxeNDuikN4n+Jtu1CAM33gUX/iHBs44O9LsXWGY
uaw9jBMH6xF1d/L868Ifnq9koJZnuuOslr91wQdRhRdPhjE1moTOTUyRL1TrkyHV
6qTNFsWR8gzEqmAlCY+69qEzrlVSwOXlRmHyNX6omFBBueEoxvi0aqBBtPHk9e12
exFdb3+e2rlV6xrZJIFC8uE8cdk7tup1tZXUntpgDD9ayS2SQEbOidSzBaCEf0+H
mhsWs0kpLlmvAPMpARa/CQ8t4HvTovI/L7AYgg0sEP/GNp8gP+JuygYdBoUq0wI1
N0E9hG/zs2zhQTHhijyAJtFqpdcYl14f7AHAgmSKLizyR/AhPXYWvFTxp+WfDVFi
9WUQNVgtiX/Nbd5y8yFtI3gi+02x0Xf/cCSAontFb/YHlfs9BEETaCL8C5kQraTx
iqxidpgOj//d8dokMsGldLrJSESRSfZNds1w4JQHccn0d/g2/HQ9ld2ELrbu/ZWK
JmrF2MOYT57LAwvhPUx7/BNAArJe+e23ge9LazwDp22OKleHa2mgzV86p7gEI8RT
IT2wPXgdwG5G9cDxPplTgUb6KV8DaS93oFi6GjUrbCt1MuBA8Ea8uOhWt6ytToB3
MCLbSvEvdFNeLjTvZH/cMY8Za9/DEvtCNzNbjxrDWO3LyTb0ij916GlBYVhvYZ8a
jw9JaVgOzer45zNnzkA/SGy7/BAjZyM6OgMwfH1XvanHJXAcMKsZJL2oe0RG+bcy
XL88NH4AtmHUyWDME1sAMr3BTbSm19eXDq1ZhfR/heF1nOg0bqmBRj+1W08BtIfD
rr4LhIDowyWcxM/7kdovvSdk5cSGjRJqyz0atSFUxesRSt9f9ea/EaTE3zZjluml
9aLAqu7nDIEG3Z0t3oYMoA6LAKM1Zte/mTFM/kzuWIKuetozA2dshCbrZrEeTZtX
+k5C61lcN7ZvblLya8/Bh6JS4miRdKdXYBsjhQury9MYF8c0fixmRJZDqfYNwGrQ
74VhhGIjLBrumN3grsG14Iln+TRCH5l9NmEnPbCWAGzN9IF54M6d2D+aBXQ/buqK
iRFEGB/xZ5JBLppirv/LA0dhDgA8XjTfRmcUK05TPxK3Dg8hqC72Pd8ruEsh9tno
LfugfnOdTwoLwILjQGNJ3NYiEeyZcfzdLdyLkC4eqgHUn6bez3yEeT/LkufMZWOS
`protect END_PROTECTED
