`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3FFSina0dZvgMnp0lutW2+TT7W+qmNTEiuWoTiD6d5eU/Dl/Hnz9u3OGQG31Uv2
StoJp95jdY4tSLYl2SEZbVp0o8Guu1qrN6qy3d3j9F9n/4wlYZg0QYUXjVYztd7B
JRQYrFyn9ujTOmnFeIP1Wrk9vbO6x3jWTV16Yl392P7bMLDOIdaCUlDXgrgiyPJp
jP6ks5etAwBLrI1RHlovxVCm3CO4JlJOXlUnmraYaUvlns/UcDX9yVZ6YEyZFmUO
PcOHRNOI2ucmk+ZY8i4wkyaJELbxqljIveNjCaxnGkdpp9fHxA0ioYmLO03csHTG
wpJOWO3UxosKHEzOkftL3QYJx320mH/815D+H5NPv97cTdiLr/v+0tpdiFEXTFdw
woSm/gZ5yzxu54R3ckutLvxcwYu7miYTrXwWwqsVsPuIixmICLOrrSCywD7N6r14
xszK53puWFggKDkomb5JVym+Nm3mHQd0wqjXhhjJzIE=
`protect END_PROTECTED
