`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7u4xBaasX1ehpDP12uoNWvWqY/7FVEaPbX5POzbJxjeKQwj3JxpFz/f9PTbdXBT
k+G5OamSfgk3F+WitMGV2LaXOM9s5NfX3luFJgwZW3K8i7tSsOTR0k0VZDaY+iSV
7/asVleeHA/JnmEdzobCZa8yJ5iLJGBK7t0rWTEGey0yFgtQeFnZ8l0W+WslIdz/
gV8f1F5jItyqbAI2GHJFJjgDrkwc42FFfPbf3SeGbaI+tkU/cuRvlbMe9HXuNE52
HJlMKPU2ywsljmCyR0jzZUkympdvYX2FClJ9Oc4Mlt5QRMvECfBnWwyDefsMUUe4
UAs9u14iWU6/hYac1Oehq5doh398AH+NkWo/THu+MJxFxO2Pma8SpnJ55vZwO9GU
vvcG3JRebyXCONuJQl19ZsVZ4nDlxFGmDmzlq5X3yUxufMpdajpXqkdiqIr44wou
OWIRQFwoswaBb2R4mC750qBu6vKt96Edi4A86X6wuLsvonPwMlDAQyTSuTDXLH0W
5GaEfeRI13H5aN3ZHoc7YoZbP3wGqm/OMD4CtBc36fkmvsgHJ9YsOrh/B817q0/C
YWbpwT9tnwLLB7TZ6Zaw+NsAF87g+PpF1wwJ0NYVUiIbQVhazEySD8eub1UhZK0W
a0ZWg5icBP+6qVzbmPca16CeIlFiUfvVLFH0S2LljYOMSIjefKvYusQp388p/WiX
FfnbfOBBRhstkefkGn/qfFCGhbbEZjrMgugEXIK4veUENb3gkIJGXJy9yBAhuJcn
yYHn7cBQhJVFtQ6QeunV7ra0PPfFzbvp7ms+1YiwQyeSYbcIxjD9iiSN/SANQoWs
OApKg+lmbZeJzN+aV9AB7AaNkKXFDkFURoNzDxb/Q/td+DgxfEsXyoAPylPehW72
EPkemK3qsJAyIvao9FjfRUgzNBOBhJsZiUjLf3y+IWqCYR+OS4fWagfkc23qR7N0
dinBJg1ePHIvGMdcTeUk8dXEMCJAJ0jlDlRJ5YPlRgc6a8FHIpSp82ec5Bdg7+gj
DjhySBYgfgbhpjNh+RRlkWuAKD8f28O7dynZgqTen22e5QmohRHWdiexKrKOmcpw
gIwFaRIL8XMdCVz6LPU5HiRvQSynVHTapYAPw0gscafDr7N7UXRTDxGy0YowYy+Z
YyYzK4/ZZ35YQbV0KwfoEiWzJ5R0SvJ6FV1BaL0b5/U3ycqyBSSSUrz1a4lEMvsB
cyjAi2HdCbPu0yzZCgDN+gI0DlVTEnDtpOHS4erz10aUSCsnQQhftE0+ihYR6tyk
+zoutphTfegtPZY33a+7JEzbKIc0ybjJWC/TJ3k1QxZ6M/2PZjQ1huHLxX5DKy2N
nKFGbvZQ+XeuslKckgJljSrbiqyoErSZs/OX55VWW0NxETjzL5RxgMCWpkDjrTbV
Lz0td3aymmmnq+2NvD9iljGLOX/vBfnmt5pmKKZUfNSkY7WcXaUZQoOPL8XLodup
RrrhS+8sDKAyey6Fl/nH6r1dzNFH2eDb+puul9JhEF3R+0i7cPA+mtNBEFcX6Zrb
YKplgWkYYCHOGpVZsZvU54ih8/FCuOqIzF0bM5xFAqLQN3geL1x/INGaurtJJkEy
l1E1a1eDUF+oQGCM4HEiCzH18ttkMJ2naNIkCgSFVkp+eWIXOSfu1i/+EEWuIkYm
LGCecKkWyws2/KVaUGoJ0Q3d1hgsefXUMZs5H4xOoHTRGSPnT58nDkUbfOUJaBxf
9N/yFrGw75Xahn4UroAU5R2nZGl/bWZp/XFdKd/ODUaj6W8y8WE7ei4HR8KwZ7uF
X5Ye/HRXJ/4i4CgAPW1cw2fx/hK00EN/9BPuLTHN4OLZhwHLIh7mKs3+QaUmb7B2
FnthBRq8Ji0g8Syfpp2Ze6qYZM2hr3Ked+UfVa+OwF12IxxesX99AtZv9/acK64d
i81fp0kmtSkcOfooGW2tIah6WG7lGG/5tC9U6bcYptjbjZctHwHdGZEsoCqM9D8O
RMdgTC102JCnXYTFK0SWBqQWSG53PUfRE1EGTHx1pOxlSea6FCW7R13uZM844YhJ
+1Ue3Hnn8vDul+/Yx1JALZmkErTHVVVdC2e38+cubMwOa23LCOblxOud98G9PGHd
kb7u1KNpdDct1XCCw/hw76SsDNSLi89tXHZ9DYnydRf1+0Dz/hhctFd/HzqOCrL1
P9jGH2SBLbYqvhTGIuRXOiXw8zOTrInUuJvaWxfaw+nciyaGlcjEQXt7HnZaTMDW
Bp7Tr0iOuCs3yTwWFKhwEXDVnrMTtBtZIZIhk3AwCd74d8JVU8VdTVAjHQVysq2w
lBNhqTWasI+AcbI68i8zFcUUSW3Hk2Fpoalt8I6SKuOvSs+Zf0clf/bevXxgycXp
aXosyNH4fI8XWO7wLG2oT1Vf/lGODvNf220UMFkjRJRrGrlgWe8PhRJVeccaOR+X
X543O5Gw6IL5OjvQPE5DHg+YRlAGBGxK0WtbNA+2zicflQW2lhQhicA3Leoon5u7
kU4ORGdb+cUOEoIw02c7UMSKfEBA69QH0d8kxXvrC8DOqhx4LaWUwZBQLRjxQQoY
JmGVdUM0rtxY1ZNFfi79ugn0njlscnKa9aBTxe0CudKZa8TUnEvQ2G7KDjE/T0cD
FiIENyaV/6r9vnVPG+05K0SaTkPsJUUx+cpLppN9F4gya6sglxdcBhaabtNx/3qk
U+4OAEtx1WvuDMhxHKtEA3RHlBgPUhbcboye7qGFAQpzw5tTtf/L+w8oG+YEnP5z
JIIT6GMTSkytM9xPmFdQG0gfn5YItIRUDJ0lmJV3TrSQN2BtauE2OdCg1bRa4EPq
hnyVnqcbobBjN4XjOvwPKitR0HLXZFKJ3iXpdHK1E/9jRWMf0I2Xt8TQ5PTohGLm
2VDd98EC8yjFqo0BOMijRsw1exqZuwjP3dN4eIc/aBmdEcGVG7pvATQelx6HPIYy
brj13yaaMujw0PtsZnlzj3jafRymCfuaKoaUgWkQvvXkOUaOLFFHP6u1obkhVPiB
Ote7+sty/rKnacuObS6Zc+ofampoVNyFB3aKqXk0xHJ7ml8QYikmrMnJJg6cWjvP
ZLpDEPJ/l2VCxCyUtuGeLh5qhzDJ1MStVkWCRin1M2z/vg5I0ZiGbLp7O3w7aGuJ
Gngru3A03+lB1pt7OiNLTwXMGiWPGETncz0JUDhHXO1OHA9umxJ99yP1Q60HVEp/
Br+aTlWntgv/E9dwQ2/j83HvWE78GtEJBaIAHIHpV4HKvbIt1IeBIIl8w+0XLUHj
27hz6+mg97VWcqU1/KtjZy4A3ho0gOwtO7VmjUA+cKUbyMBD0VSJ1saKFm9w9PjP
UAPpOOd420g+Z+0chAX19GouAAJh2aILWjo2cJGw5TqjA4E28coOiAf9ZTkPjYdk
3X+LDCbWbj+CJQf8Pxbh3er/wT3qSTfdyPyvJ+jjokAQoCgit4ZVt9iVc0vyCofb
nB7qUQuNLfQe/F/q4cye97YkXgXjARDLj6haVWjX9hcWPljDVy1EeT4ZXObp85lr
VOAU3YSM8hOXgoQcCAruf5rhT64zxp60FamXAEDYISpJcgJMfnbvBDQKjjF/f4og
+lSFmHyraTrkMjCXExnGVVJ1EER2XfU+Vbypr/p/L9EFGcAPEg5NOyTe1PpwzPQM
J0bdjILepIQgcdWMr19DcRByxH6m6XCv/nEZnrlqy3P+3vOmI+zJYp/MgzCgqjpF
nXmn39kqTcl7bt4sb7qIS7FiclHYdqyWnMmobyLdSQAG5aPszGaKC/iUqYb2IRK/
vAh4GRw71dE2ITHkPpAQyysY0Vx9/78OzwDVlEofzPPD7MoS6QJR2CWZAA/CeHRa
4qf45wYjgNNRU8jOzZS9IG3bt8vlo+9Bqx+tkGNxdYZ3XrlDcF1JNrXYoz9BXptz
jB6odfARK1abZVpgtDOnZ/31F6r/Re3GUIsf8HeeThLS2YrWCYwS6xiQpN/ujqbl
Twc1bsgCuZVv+KEdfZ6zZtO1HIMWfzxosFjhIFO/Pe3MYqldhcQg5jCuMmMkiYPi
H7mWJnnf8APv4OD0liHvIjiie/12GRjIz68SATvl5dXd2fih3ayihP70VWMNMiI7
mnMl0cb0MP+9rYlZmsZfROlb9fW59lovIDiPdvzg0S61ecVPJ6em52n7elV+eiw7
0KMS7oS0khRoM/70y2gpCKyWSd/Iq6sibIF7PDSChomLtaLIEYAiXQ0hmMBaZkcK
tn7Oi69SKX/o/Db3ggNvd2scVvC52nfD6SOy7o3n9yKO1cowNlKlS9cLMKM0/StE
5iF/5kYdEtMVMB3F4kgBvWIRrmcZfS9srSYjmMdgPPdlcqi7UMpib9jHPOF2vb1R
VUWJwh4VX0EciCtLKUWJD1zbxYzd/4VvEPbT17P8/AwLkOtDCqC6MxeS4x7PG7IN
apq3zgvNC7Rh1rH4RQ/X22W5RSUM/tzl/3Gi/8hnq/D3cNmGQnBA1Z5YPu/cuq/J
cIywFSOJZGTBh99ZMCKAgWpptM3O9LCx974uqZRTJpLgquG8RB/3b71sUSJCfC8z
/dRGZ8F2FnRKq+t/7kO5idNNyxbu9gLKqK43cTbtJfQ+m7gaTKCX8ai/0MC31Wto
94h0WMlUP1rbjdOYPp+ZtKEUYnaTI+VLTU8vJMPX/uQy90lBs2S43xbqXTdUebgh
toBfy7No9uZ4+KlWODeXnE6MZbycu5MIRSXWd67Z8K0KEd1En+pJyExbnz3vuan+
1VP+uRZNSm5qeblViWyBFM1fvXlhBwYCdXCmN78RH575aWdFRxSpRyurf62JObXg
OjnYEd3PFUQJ/pAavt0IPB8H3uuILwGbsLZQYg3SytWVt8nroGGOZbM5K/DtF1yn
2HjFHft+ef4YzhQ80uh2/DGnHq+Mlgbuccf11k6ygd6xQUHrUv64gQFter/PhsIk
77TU0Bxv3peFxydajrGg/GZVdUt5PL40Gin/vhnOYBNHc+AB+wG/P8K0V1sZeKL2
TovFk7m23EL9/6NR7AqcPYKL4c1skJEyM5mkQO0x0EsUkLykm8QlPy9d/QbdcZ4f
odBfmOEd2WpYFaQNuo/Z+3jNzWCRXMEBXn31l7rdm39QETzyx8c6LT6MlN2gtE64
jn7CoxXG9M0Evkxn1Qx/7WLRCW4Db/ENuWmt6mLjy5BFFSC2GybOLy5xoUz1e4a2
0ZyLBcTfrGQpA8YyZrowvkRAEDjTUkz8ld8Z5W5HPvnlp9LcT/sVCtT0wT75rZmF
B2ANnC+vmx4XV/p0yWGZeDv2FQuXxtkv8NO6Ed0K0ifQusNJ9jou6zsdXw36/oeI
S7ONteb7f1cVGlvHdLmke3MXKMgaRIKjVhv/FREpEcIgW8Y1YLtRzerthIeLwC/P
iSPNcMeGLCFeLrtvumsAN6qxfM5bHqIC4HmvyJM+9soQA3O2u7E36gSZcdFoCL9U
VJprGsfZWooFY2TZMVTnaBmt+gtVny1PZ0cQydtO6WKPf6EA07VeU9uwVxjAvo0T
uIKdFttiqBu93T2I0xJIrKqKCkpHsyX9XmxrkK77VhK+AFNclhYcQQOc+E5T5CW+
PM6/hPAxlXmYUc+8NRMxxU5HAH4C1OJzc4L9dSr8FmX1ybNqSDkSLCHaOovOPD15
zp6cDfc2AJ/luh70GB+lcLTCC3CFHILLp2QDhmUKqp7VoNZRczDpQdTxHfn2I0nP
L4pavSB/PM9fYtIVH4cmiKgebM14G56ExFsdSj03GtJxRvrtseYhlt5OVZCBRvGp
zR2KUPUpvf6V9ImfPNP9LeC/OXebti61n4BXxuGFmGDYrzc9PRLxRbzRZ2KMxjVA
Mkci83DF9E+ZI/0r4I0eyT/pQT0tzh+LX1h3GQlfc1YbF6LvSM/BOKNOtqIJPR3x
jfMktzOd8yQxo/x/A+8eNLdrtNGGk+2PBX5mUuEfRy22djGlhNXmEBRH4NaG5VPy
wJRjiii3XrxSHp3auUcHWXtYCqLdAq+KpETnd4lbWLVRK1xtxXaO5b33RWwhNpVy
pFYuPzBguVnn0CBlBq3ECyc00uFpKmW2bsh0Aqro2kNd9N3NdhM8+/mjytrOhzec
CLF9WH2lnCRB0eBnWQuhQmSHwBPBK09+eW9+kL2QJn5ol8Vqo8Tttc5zw42jzUXn
Ay7xfFg/YXKVG8DvYVKv/O1FLjDVDNYQqKpwsUY37k9hYZj65ZPAFNgPl7x4ltaG
1nDM0tbuQyuMbTCnldxH71pQKsUGAi0WK+INGWqhFE0fSKc877rhItVUdeDzhlM1
9lYK49OpM7WG6iKEi5FEiJO1RO0Qjkp7vGSJBWcHV7iY9YE4ix9advBlfjI8Bjf1
W59MmHnZRkPzEcsiMq/dUuPs9SxuxYIzLJm9+aV8czSGW2ZdLmWHj3XPHOSJ4p/K
yg8lbtm+lxVcrMQ5PSC19fi/S9E5UfzvAAeCZHgfqas8OiEoFVTILW3tw+qDSj6L
D3fPfmFwtWlRSbr/aot5UOAhO485HaxXGy9L4aUua7RCZQEhtgC18vmdcsgY8GVC
50nrCT3Y9xS4DoVRYXP3sn7ZAzxMNdWLzH055qzQglZOKqNQr/BwDIRJacF+fhxK
RyXZp6cy2LRXkVQpX3CEBwsUGHrcdtGzgaRIaMt8xFlSoPbmBP01Hzv9tI91Hwyf
Qr2XOVvvJLVng67Y9P27fWTKSEursyVt7PS62d9d36vU128O8YqosLT8sIJx8xPY
PC8J4ZrHcl0U+g2sVRr7F9vc1TO5WrhUNMP8rT0QqceNrDhQPZfzMpdUvdu/J4v7
lTDfly3nQdg9cRHFwJOL6xU7RAsrkRKZONxul48FOemxC7Py55Um42Dv6T+nHe7Y
R+rqrD5pCEtyRRNSFWf4H1p4mVUjFmBM1/4+23JR3IYm1GemC02iwVajoXckzrh9
f57LFW/zpQuwQ4ycnlxwYREUlPQGd2+aRlV52nP69a8CV6nEkfEN0HsDcLEOcfAK
fF2fDFcWGs4BSTFCoxei3IOlPbwrcITX8TUDn8MoczHqCiue55FDbDHR6WfD6Nq+
oZ0GdqzJ6Zr60+4wrruYASmnQ/XY+5gTkjaGBmmrLlVWXzqTX5tU3lGqX/ifY3wV
dfhR27B3sPIt3LiWxNYRkM2wwfLVXmnIqJ4y+U5eEcuiETKUOmyRvrcpVYl4sq34
LiSsEzdZBwhnY2WCbiZs27hEWhaOek6xi/hzLVQ3EoNMU63PMHCjFyNqx2QxoB5h
GoKFO0HZYgUijLCeTdb+jywSgHE477ziVd4A2bNsHNlwVOuRAUQZbp2XJbL1rui6
4sU/KwSCtHWx9AHqXj4NDaDOlbrYX8LKG2z0CKDmU6Cqox2+LihD2d748rRBy+hK
QjhnnAzQUXG9X/x4869aGAVMTbuzwrngFmJi35kTvY8JkHX/KyuyiLviiqdSV1v7
+gEpJq3TZ4daRHmw/cKXpaQ2T2H/VSB4o3bNfmldyJaM1G4faOxmXeU7sPj3oKIJ
B/3SPxHb9AdWZ9JWjp17XdKpeUoaIY8726g5zsVfw3m+3/66/BJ9GoelzSnpBptp
TQVtPvPBFI7IEk45+qwUYNV3v8xL3n/AS3+hs7vmiIkGT0JUvBvj0x+IB2+t+VBz
YkgumWVNiRGSPOpZ4pD0QNNSiapFjV5+9NyBtkb5Bji5RQe9eMwqVxMJZQNJ4hFP
t18f9Ho3wiiRtFvMrMbXMcr/L/a3rbL3G0NSjzDgw3QyFJCN/z/WKTbegTEEAQZo
EifeO9Wjuv8qEl1VSQvtXOLj/ubuZ8Ue+d9i0zywbV0Ki0DqssCHGtsh0gZWrqv+
KemK5J4VuFZgFMWkZQIQjg==
`protect END_PROTECTED
