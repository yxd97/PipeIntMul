`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdONAsqFoT2K97MQTgtdoavIgSEuJavZe+iM2bV2fBkkcUwBMjl4G1JZG5sdLnYX
82NAYBHXLhvSkHJ4egW6L2x30TzJIGWJnOH+KkFUtnXELQ6DqlVVz0Biwjj3TKLn
xdPKMnpzkzS0MuRDmkaNI+gg/6JUwUAcP6zfNjkf/doChrSoGlUEILRjm5z55V6G
QUlhFY/6jxZrv9YpzI2wwCgHQEFkvF2KrVjp5kXrH5w0B8teYjZLPEzi76a9t10S
gQUBajkbU+O9KsalIcRZAPwgm6v+5JUAp5rqIBlBDqG/bpNuGdrzb2yvgAR3nEkl
TMm59TVl2q20FHQrsIxu3ejuUL41g5sMC8PQoqAJTd/5DEUZ1dNU4XCNdVtPJSZP
zbAr0L3sPApvK9mNKGLOWr2Wk1PkfSo3tFpMCdAjfoY=
`protect END_PROTECTED
