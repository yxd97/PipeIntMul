`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGpMOHlbkowiE4o9ulDU+fWFiuTQpP7ipoIMJHVTJ/D+eHxT0aaexdTmZgeuFOie
l/kWbyixqMWZ7VU2RJzAmrfePv8LEGxvNu4SvPPK+rhaefn8YYrTIHEeoESqALka
h6FivStNNQvCEgAIng0E6Z+sx+IojXnffW3v2nsme3DdNYWwI1cfsGnC8LXBDm0o
tDv+EYSaVl3c4N8s25xyZ5+C9voiePowFi0WNRPhgId1MHheaBEU3FznJ0+Wc0A7
0F6XVQbMQvCXVrFr7Ci9lOHcnThIWk6ME8U06xLW7w9nrY1owlKaxvaHpBROOTo5
erBMQu+0EMg6Dlx1IvgVVuTFF+jMdZk3W+eepo5Pwdey/qcVOlvUeiJsBFZLPCMs
eZMNokwxlHVCzgj9yqjB3w==
`protect END_PROTECTED
