`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NMkCWItUfYfsBCbb6UzjqiMbHsyPUn4ne4iC0cKnsvXokrXyPlLTnS6TRowukixu
A+RYyjTUpGGTA/LdEuF6Y1eBQHWYYh6gjz3M4HEROO7N/ZiB5H+4kolw0bAp043/
XDoWAFYtP4Y/46fHdc8i1loFmQKncDsadkxNA1Zx5gd4xJ+fqxKXLoiuTvzCGJq6
kpuhw2Ybj2oDYT7PnHmIgLKlLVPHNxDkXgvCwSu/XS+G83H49VbEmZHJktVHuEFp
I7uk4AjWUWOwsI1ErcqJwvfjTLrqBq6z5t+hreN238yWu/y3WWVH5FLacBXsu4fF
rVcDuuVtYHkJ7qetQexQBDZhYCFIZbaKJqIpLbd+77cUqE6TiYS2FN/jbr11oGD5
v00Ht+UuyZMrkWJcn1xmQmLFSA0p0TT8JnyIpusr+mt/1f+TGD33Y5tkj7nSkT7y
1GV/7Dsn9yDIwePnD3dtH4WK6PkvYRgQTtsC+zysCdnGWou3LcoG+/IaXSkt8+WR
hCdsw2pkBWDZ9IiyWMTray9tnVi6116ncpJGXWrLOQlq/cxo+0v0/8T4+1kxOmw1
pi4fukpbCtSapE/YtRuG3PxkaKB8tsHucRd38tPiMd48JS8MaU7+W97XDsGsx7/L
n2ScTPpujoz1+JQFjuec9kt3QUKOkdQ+Hr7ZDasCL8cVDNegVOXA5yVs9UxbR7E1
0NJYdgb7qtR/n3OnXM6If3CNW8ACtvzitIwrNzvKMEhuBufRne3QL/gojN2eY9VO
C2jGFNQp7vVLj4xeNBYOdhy1x3cfGocHpyJoBxXrXXNRgS2f9FXsPkz1DPfWMMod
ElCmYqgm1EN7VJr6uhdIiysWuGKxIYz30vNdcUurBWMw7uePrHGU+rQtXyqdv0Fl
WvQDYi8Qtvo4jsqzY81k+Q==
`protect END_PROTECTED
