`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkkRk3it8Qq/Fob8Vs2ulAsnsDV+yfBc2gKYH6xg0r9nQwrllFrRHYgiR0vMASr0
Q5+tuznkP/yeWQyARh+7BAypU1O7Hv5vqZIparL7JbRo7HV6mWe9q4TGzhIF9T66
vRkkLx72MJzkTXnpodAQQqxwfOHBd3Mcf30+4zuGEP0Z03BVPopzVSUmxHo9eKzO
LPckKnMC0M7EyMbd+TiNPPiInM0cy8TK2Y1FgzpBRjB/Vj9w/O3KJdLwIbt67W63
UDOHflYGjYQqvLs7zhXgbqwFt0iy8XRuL8ydNWYLB4h5N+SxUiRE+r3j//1vQoHL
w9F7a153xskYq+HFdXZgF3Q0HLv6sLzE5w4afhtt9hzzn0qWuC1lUneAVvTLGOSq
hleAlwequlyjs0FEAmBoEQ==
`protect END_PROTECTED
