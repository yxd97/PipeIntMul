`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67nefprvc6cVZj9iYbAjCcF1a7pc4w9PeVTfe45VzlzApaF27G5BvBQXOCznGkUn
TsaKHi1dmkYr6r/toAMPZhI6doUMJIVge3P/ZJyfeb30FDWmVH8HreDSp4UxN61k
ATXH2jSq0Fwrrlw7YOJFQbiDx4j0KYwHL2I44X2OJWTDBIQitoOacfqJPr3xQfon
UD6mKAwICAurLsQB38Ge0QAqZxzAgr7kbuSj0xTRbFD8+a5VrFOFt7uZ/5lF7+D4
LuE/FHLRZQzV2pQ88oDgSXugxXxOgpL84ZK6CR2rmnNIve5eHpgphkLTY/fqMU8e
Fyt0lFyG3hCM1C2Bb9KchEO4NW5ngM30C7kUmV2bIKI+oGBetFyX4Vv3mb8PNbBE
nmKpHp1KpI7FV7qObFgrZB0pyuMQRBuVEyDa/MQmcr0TuVTA0fmKRD9E3549otKt
6a8gG49s0YAthv739TyzKU8SE5mHsLUe/YVZdcfni1vzECTDfr8Nd39RB0Ys00Pt
`protect END_PROTECTED
