`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p2JfOfK3GLPl9yX76jacpUxggsb/5t56N5z7cTSZh0Ft/oyJdQWzXDxY0cFS1ng4
iPY8KHiz4MALlR9fmDgKPaCbDe9p4HJkZHR6ndYJ/QOB19ghkAyQJDBPGcyERBj/
IGNL+Pu4rIulnXILSKR08MoHLBE/5zUe0o7MmAQUkN8JeHdMDINEzCw6/qgoKLo8
SrjUJ8oMbG/gcEEzvJJeqJvAtw5APRiogYfLw1aaOhQr8zh8aYO+KGYyYk2FpZ2k
KKyDT+TAUTcNDjLF2gqqxmkzz6/btjZdNGeI/M05q94PJR8QxmuOWvLriQ1ao2y8
N3dSkDajqmqICvX6a2g4ZH8XJrqwxrVWuRa1hPhJp40brL4djMerTjOICM55cZID
rj63b7esk22RKqHXstjNyw==
`protect END_PROTECTED
