`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VufqRnNslHnSPd9V4PMBn/GaUj1GCpjm8Np+P3LJhIlFNiiSQuMMwo1zZ05KfvYP
e1NEpWDQlTjfJmUziGOnUxWVqi3hCFwURGrm6CuPtz7aQhd2W0drtAH10tLYqGip
Rb5jedzq2U2XvKtOCBLpmXCD/IFRY1J8iP4leMmxixAxdoXhptQ9oep9ItGr1mOB
FmNTa/BMXicBoEs01lTQZmiYvwJPBcg+f9V4Xn6pcXfNxIvOi81uTUDZFXzegjoZ
KOsAUxzSTtUzQN05OnBY/jY5UBNDSElLHG3Qbbt1rTYeivNC4yIJWtCUaf6rNguh
N0XROTaPERoq/tmKuIRpZei9bQKozvi53yxlFBQcgOlu5YDmhS88dVPn3kf10IeY
Xlkzd7i8FZTW7ueXMZG0767OpEHsVmDYqocEBouA417JCz9kI5zhp0Wilihyioct
zFquS2IrZEngjqTVbCWnGM0896Cjiq+43B6e25GHMAMzXOYyy/f+v6j4WbcW4iRQ
FMpuA3E32A/VnDGr8rzRkA==
`protect END_PROTECTED
