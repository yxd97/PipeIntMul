`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NUJSAvwSvnyS+qkUL0Sh1mug7TKHYxFzjxRpsOOMEihIU7+7E1UkAw/6hJDu4UoF
9F8Sx8NQMLsCN9KEBr1D7VF/w8s48SzghDUI3zGoVjyJxqV73Dgu2HhwQwIPOj1O
ZxX6/Z9beNo5gQP0KPO074YC+fyO26E4fvNIlP2SQdhNvuEQBrbdhkgsseYJ3ji5
nIInpk6b3Epqv5dFB/HXPX+2tAPeoy6J99P995v9FGPF9Yxgwl7CsEEgUWXvzmgN
kovXRA+3Joq7vtoWkqYExEreko5GOkYlhM1Xo/cUzXDMkbAsf1y2u99Kpwb+kf5o
WOdraLWJxRZkeDZCG1aWIwYsHIaMzxOHMEpX/gh6Z9esipaqnwigUivA/MgvTp+u
ptFntiMvxqlVXdiM1xs69b3q46eqWkCgnDiIfGrsCBscv2YU0GfXii8tqow6gO9S
39s2f8JDb8u2JRB0paH9LbQb7poftBXWzRkhls8vqpM=
`protect END_PROTECTED
