`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+EgMHo41YJfa7ws0AWfYdg8oaHQnV7yrjs6tsgn47geLqxJH38TOJswf7KsYIb+x
1MNd7DyZnNYJ8+kLGT3YgFoicyQuYmcng1w+VStOHNrVkpcmBEs2aQPn9B3AEIyP
T3D44xqoWdzk0u3oPccbHVqBYZCISA4OX/kXoqfqgtB+aVgUjHzL6DJQXbwWKHSh
NvTMc7gwH0WmQKk9+5h5GmgFBAqyXhUzBZoF5kGlRYHX3N1s+YIPmcUC7cQaZTe9
Z4jp+OLz2pkdQSsA8kUOnAtP4DTlCxXMe2hMjxFguibWCM1px2k/VWBm4KZGTSVE
o3rg98f6aetFXcntHHkctMW0eBLp2Qlju61slgRC2qlqEYwnnwuRVFW8x5DIkLrt
3cvokwRZ1s+Dxxejq8W1gwjA05jRHNbZMO/+y9HkZYeg/pEaPmQjmMCsZSKE7xZx
dmg84KDuvwr3VMDQbAQKar12yDJgYcPZ+BwvqSTPLemyvSvef8bcXhG1MbWnZsre
bgPK5tXVUE5Qy9WjHCPwdr+mjVhyPDJOQ7jSHuvk8K8AlldlB+STB9y+elQo3AqN
57eFCK7pglL87k4V6eBpHqlYm87gqo/QT11Ru7jrotFjiU4NfW+myUchOtYYzr05
m/fCp7yQ6yVOPfXgwvhAFauRMRKBoBDo5NEEW+0/sQ4cLpcZhpHxkUvQIbRhzWRf
230NLvKaCBbRwpre1GqHxiE/gyyGEVNW2twx3TUKWotAoJTOHu6t9qJdBK9wnSar
+af5ip7l0p1pj3FW7wbGRQ==
`protect END_PROTECTED
