`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kf4HLhvPeFgftj6mtzdP8kiyj8oJFgfT29z0QDKct5uWgiczbQLu2mlSOLTBcc/0
5FNqUylW4q2KK7TwDxr/xOgQkD1wnOG2FPuXyRu1aZor0p6b6ET724/r5W1TdGAA
oo/MGllT3W+9ijioMPi9tFJbvgp5orK8Re+5awqfur/Ny+klIMFzZqcBTFg56S28
JsRVGgaAIvRbAiHWLnkqZ3mEONydJvW65BtT1qjpyAM5Z9xxiGxL2rtH92IJjR+g
g11O6CyubJb5kkgCspp72eA1x9i8eqVgZJvzU+dtVHApwdBs4sNqotwVnmFkp/1q
npbOja2/s/UvaQGcb7pKjENx/tV/oNixha2dhZQZuc6Lo6GMERRCcggHRlRcBCy1
MQYf9vmJn4CMrbM6bhJ8veOT8R762ivVLMsGi2ITk/E=
`protect END_PROTECTED
