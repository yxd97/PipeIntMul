`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GuVeXal3oVEG6FiVIE94/VSsX6W4EWTqNH5rtx99enuMvwpPt5uw0rKAO1su4E8T
SstFXoXU2JN1IOTlQvqdkJax05SJgDos/h9CDeERdHwLNuWnaEN6c5ETsENjspLl
7Ov5E3jA4T0ZT/5+y5fo1IWmgGY6LMC9TbzV3VALTEVSaOdOV6mRI7uH5lKCqmkw
hFctINClxx2mle8RHe5kFPEZNLXBgIy0QWs6MyMe6DEDfhVUJKTKynbQ0ixwMkBM
ZT9e58ZH0RRaq2iXhMLzaPT17Hht3zH4IswKCJuIknd5UXhK0/1GSzMwjmqYJLoI
TBaI2ZU9TnVbu7BKb1xQdeH+Jf/HNkvSKQfgqrc1BVvpFAtE1HZkipiwdmvxTcq0
LxoqyMiC6YAcR3VYV83bHA==
`protect END_PROTECTED
