`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VfoUNipvulncQgIhVmtLVBoHN/k3WiyxpzpgEiyR01a1yqufpVz8hGncX9flc0mB
gfNd4UFJ2TSEqteyYSm0QEpkh7ZIbbFcASEgKJ+AEIxhJ+rgayk/ipcGHFEah5W5
oFOSEKqOpJooaDQZFdjkPZ90mF+WdbAQnZBz+WBQO1F/oFK9Dp/UkdFpiToucDYO
ebLW9+pZz6OidLSMJ3m2DTHB3moTYtEBC9L4uCqAUp/fuI918VPDxysDcFzEfeEv
DaPedSK6x2DAkpPgHz26GcgCuDfIl7pyLq633VpqgXl0WpMq8bja1k0WTjxKho0b
3vjzXy24oipKNqNKtSt/36esmNiLvfDc9il9SY7As5Cm3Vmbp6PLW8TttwWFwsCH
qkSxMZPhArwkJtFTo0mTGLYOJuFGgs9wh4fsR8M95uXoz7yrg7hqoNsoAkNwsDsX
/83YKyaXEuCizJ4NYt1LW5gTun9S+p65vYUh0hqj8BcuX2z9mmT6U0cWk3hxSnvG
0ObfALow5GJ7oI4wqsN21/jpLjtMtW2cpWoS+F0JkrzpGSG8L9sByNmfrlJ1Kb5h
WoNd3QnKQaigo7WgbTQ4kzUD2AyHqQkramS8MBUJ/WjN5NLqRedKG08bTdq3ED4P
jumAFQ4q6rfZhLVSQmH4YS8C9toD1Wb+v85R8LxJ70LErVeRqmOHUrlDbNNJavIc
nLu/Z15iWvz33Huj15rDIQvLSQhkEWFfaPfRToWdHkVxPyil03MVKepoil3MkRsu
gAyEiltpLX8a/VzRbbINX6Uame0K6n99KG9+4QgH+q8XLnjOKMWIvlgMiy7ujc5F
8ZYPIGIm1gN+dBr26UbKnYMzqmHPfZVxDLBkL1wvBGFVrOoHBxc+Tlag9QPcR3ZW
BYXcayU/GVXM7o6IeYHCJt2obXk5UDTGTc+Zu8Vy+b+JFskjQcr3RqGsYbPj5cDM
`protect END_PROTECTED
