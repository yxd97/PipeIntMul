`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
903rXii85b/72HfTiqgfJCrHAW8B0h0nTnimYNifkkm+LWQ6OWnuqTPFEBHvwsm+
HDOTu9qovaJSM8CMfLqPNf/4CIol5uMUbTWfEggzAYS2El+E49PKr03Stn1T3XoG
Z7optWO8KZ+ERhU0DxM+oClz1/v4bxPAWzKRAaOf9GTQHdsWDNS68GsRCPSRvDsL
uVRbwz3sosqABLCAFEEm6KKn0NMeuWYqRQGZm4090zpRK6ecyllo64OCg2DrR0wj
zeL5RClfBzfqzV9/HHksWrIow02gLvIbeN8KT17U1ltmxv0yk3q1WniPccJF68NP
f/KFt8a/vbjC+wPCcUnjxkT/daveiX/RSTpPGm+zwJxGefwDss9HxBtKQOmb+0tM
4ubI1/QxaksO6NkMuGszp+5YtYFXnHOxFSWFQuGlBn8A0sJc8n8rPsTYYdL6OUrJ
9P9cdGLY+7UseDW+Dc8nVhE3EwgFYbRaHlr43P+DS/MMx3JJHn5n8SfNT16xCqx/
yoJD43Co2w7V+YH5GVKM63icTukR12FSolaqvFLoOJmcjNjXmsy33GHuzTjaEU1r
Sz4sYyGXApwccwEZ9EB8tuEeO23fWyk4PwUUVucrYTBokWA1DtK4yMi2k2IBLMKS
VcMJomZC1fatQrXVWeNfNsqunk4a5bRMusAnkzlz2cv5XIVU95TOcs5mr5YJu6EZ
FUrVnKVe2AtNWu3EnGks63BkYt9dHAXiPS77NSynTJ2WBnQURMcARHKX0g8Uv8iX
Li6uUcOvxzeWz170sDcwuC1LxESnFR2zu8QhRuz9H5f/ckF7rFRW+xaIPZMEvGw5
Rm3qXMsyf6DTGMVOW7f/nVxrqcEjqCvfQtAvG8a59/J9bXhMgfSx8lzhNEHlrugL
E246+1n2wrVu8mhGH71ICEACYUA2m35QRX7CCkdnwV2Fj769vOgQ3qotOBw3sNNe
`protect END_PROTECTED
