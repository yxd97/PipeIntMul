`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OxEXnvKfU98BDtYIYknzE8QkzBkdEqG8mLATLuPs5wMASn9ZrZQ7rI9GEkapHt4m
usnMSQjYKc9JzkfxVsN75GXEgSEGugFkh7+kbYkdFjPg1jU7MY8vE0/GkfVwNVeV
xIcPVWe92dB4E/Hm3loLyTtJBicBWBnik89jzaHBUcye8W5kcO5sLIuw2bYD0RQI
uEmJR5GUuMBZSQNRMCc9xd5I6fcj0T8Ao3V8M5RMW1nbwMXxWHnP67xlSIlklmqd
YEd43ZiaJ3hjfQShtvM8Qhczw0W97IhCXYxP4b7QGitIcsmvAC9ggWk/1yZnbziT
5wF4pPj6dzWQwYpd51Ap58XAMoUQTCTLQwdocxAk9AqdJIu42ha3Ox2udFY/jJiJ
WqsM98LRDYDlCPBuWy2tVYLUhsSzkhQ7Q7lceeWYhLI=
`protect END_PROTECTED
