`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ub1l82jbRrwQapGBXMZBmti6qw/3qKlC139B5LW/iUgtYx88Nqala78kONAyx0EH
gbezwLfNowI2zee+zhiI+5RW2JRdifFhEog+bqUPCbiMTCK2QbJeOxSxhNtBQ4wt
VLSQEW1OiVuq4Gbx/1N/ZKTgJD2oPQuEFwd4H+/kY0/CcszBivALfaIUjj30T++m
faF5wO93oKYjXuRymIzpfIeSGhrJ9UJ8QUryyasonQCng7JJeFoB35xMSlMKO/NA
dSScuO7thIflibjbQ25vhPk4txAGIeTg6dGweIu04l6uVbZbxNlY8bLUBglgFPEP
zbGPu58xSeMv32Bbndwl0HQ6dWukjVw2OkElEI9BP/+/nIH6n9Zl65hKXh6M3v3z
X5lBgVpoFvdl4I0Mf1NQJQ1IWdyRAnHG8meE+bk26egGf128TuO+oB8JotfBulCf
5h5uWtoqOnW1+o92vJSyzDLm3ed5vLJLeubhf7Ia6wqJW0nHV18QXqhrTZKlv5Q0
qQnIKTgdmq15LG+fvYtw0C78QnB46Yebc85Ld14P1BJXg+EMbeJzOJDbw/GSbOrH
SbdQz4+bQRSZw9RtwHj9p32W57vwCztC6w2vmttNHhN5NHxsrZOGkB/w+CWPRrju
Mu1MyqLeFHpji6gWnkeQPF1AP2yZVVou9XdQAlbkt9TU2yE+KyUMQQm2KPJNvOCn
/Zisi+bUFITVAKQFb3mGBvgtSUwJ+l5AS5et9s6T1VJ6Mjeuv9qxw0sEfpTvHW0X
En9Gco5PUWVf9jtIwbwGjhOmbzacXBMeVVFiPZbAwipNSbWCGwRBIvn4KbCWhU4v
0vvYg169QUMDhzlfSRkHw2mWuvgomT2ccuRs+LhE5gwxkkXuIaFpFI0P5qKMp4qa
VVP2wCtFx5KvVPWVatNTW3+HJj1EjoiI6QLrrdIcQLDn6BpCCjupC3VpHALSx/KU
N8jnphITtwVK7Y0SzdhWKllhJUo0VL9X4bs/QJNoVfZGFYFCoFPPhOKFeHBAeu8m
/ZlWCDl2ENaFdKE9/bZQ8Vab+QT4wrMGLctnY03wcQjxD9sE5wPqF2TvffWHJZla
VKVXx+g6g7yPC+P09S6G9Su4gAwZEhdKaQzaMmHvr6iXYBw0GAgzSEix0ecUI50h
u4NHTRWqoXnsuBQSmieOpGargqyHpb4jZRIrK+WpJRF8Ub02Ag8Ob8dH5AlRg1Nd
N453/8YhdPy7hwgOc6rh0vlURSwTdbUAYRPXfwKEKeup5wvjqi80FLFUVCBq1P5u
WIklAO6TZVXOxU7IEl0ohdTjyL95gC41IcYLXDBlnp0sYDNZv9y4xNPgyHQpeYap
km7NSdXqGNJgLRI9HDkEht8uBNWPh+OPo00phCWi1P3Ctt8ziKHF2ZLZ8LGVbEeS
Z5BwyI5FSBK8hiEOz32+uA9WJDseIW9EsMzp3jFxP4qM7W/vFEV2JqHd3qFeucZt
rY5zwE1beIDQR6XB/6fRXtPyYHmUeAAKN145PZWwXf+7PWgvdPwugw7ktzciZ+9/
PpJUUaXnAGmrEesMO02Toaib5OpDVpzAuOd9gI6jFgKiCtajVKitO+uLKMwcjKw5
cJ7Mg9thy6h3UQ/WDGOfKtwP8VHcjd1LRUgreXEPsSEA/MZVADkAfsj1V0cJhUkX
LIKDWM37wUoo/RsVM6UlgL7zjzDg3GAdYUC1/AcgwZRVS14roNg3eYXPHvi8oLh/
6QF32+wTOmSIeY4DNWtWn9/ds8oAudbYSPYlwzmP+BSSrge3KlK9gsAASa6i3Vky
2ky3R/c/7iFSQK21dygui96R8Aung6TaQk9Y7fzuDTGmia1SG54T5A/E+L0YSHx9
px281hgIacwiN/AXvPTsvpVlNAGozwv/lR74Ux0mnWYCu3rYBS/yRm+tbI6S2g+l
8frZYrjoi7sQUJfua+/amQEGuVB+25s/ZXqc/AoK6nCYIGxMrY0Tw4SpiPeERr2O
lPPdRnUpGbGyBRjRJu/R640rp5JVeOv1I9U6c9y9/cBf4nH/8wczd7YFSlKxD+DR
WsPv6PpLpizIOLotYUl5j+8gwyxHj0qBjLOVgYGhKQD7+UVcfSZrQ6NnDKSmJcbQ
fFBLs0TaFoc0jc/oTEclTwn9xJTXKKWa2ESc/AGWR3Sk30llPqQ1yVQ9rgxQErKh
hgKRKLo1dv+h2wEzmCo0rvKGVGhFIQdzO0kjF52TJYUurBFEv++cbWzAlaeb32Nq
kWsBWEvN55J9Pfg74GllM4DJDaMromf9imsFtioYRnwehE36NQLIqW/0PD71AZ4c
2YwcwZxVhBsdbnnQr14fv672HuvsXg44X2kFXzzWpZhxH39J8PPT86Y9p6W5i4PI
HoYzcFgK1yK9961IesVMF3zqrILn7W2xPEDjWlvP24WgXR+/tOXInVMn25T81rHu
AT4rdLtl+auJo3quAi2i6N153v7REj+yt9dOVQJKVroYwAnddwXqLgPGM604OXFE
h+DnObkcjOvGdlx7PhXbuvuX8Nz86/KLeDrWtdYquSJlYAs8WNed54O7VsIUALeF
agQ1cw/t/aRbdFFI10vT4yl4IT85o42l7FcH/T5rtHk+/YhhmdhDfxVhWD++qd+3
J3IaZ0hTXPpeGSN0yRi2P+vT6LC6voTstgjHbhu8gXEwHnooNiQDARRsgbU5xyti
JBM9623A6ySq1xqE5YR8eBELp8ma9tQqjaPwk+cSMpwboarkPCspP1zSKRvYA1Tt
Jy1PDVX0GyIzxJLjZoiN9mRnHlVDupzTWvckrz4F3j9yE66jvQova75LIDcWx6qW
Dnj/EUxw1wcCLbTNzDx+mKJ/4+RmbpfuHCROFndgqZw4b0u0SbOfDQq7TEKdv2Oh
Xfm2vnkvpTJlf9WaT3n87PdP1LlOQdwagbNRHEiVyE0iZMPPabbsF7aBMr0hwUAg
ta1buR2eB2GtmUIyGE0WDO/K3C9P5pNFcUQExV6H4ArGNEj2TYXowjGc3qNkZcNi
qzEpg5jDuahAJ6R4XBaHfWF1so6Q2a4TGJrHH1BsbBPlp5IQWdlf2YAQ1JC/X1KA
zK4O0sILP/JOFGwEx+mAVA/vl3DG8TnxmHBFI8Qapc2yUcsLjCXsnJFTNxhRXLUY
T/476GS+BfJnyTX1kJeZCkjm8JSXwzSPVrxuwUbbjkiE4nbN5qlYslYBM2LFqaza
E5D+vZ2nWjN363/OsM8rsxG6q9PgORPOn2Chg6W51jChJpaq6IqB/f652Zawvu5u
T2Ukw3H5TXUz8wE5HRNlzJjrj2XLOwku5Y0Yb6zrSKCgmy8BWb8ssw4cazX2mfKG
ZmrtyGcQVgbsIcy313RHCVYLuVVI5cQmAC6lELm2PsCwYau2nMMasDRtar2hzGrI
H/tyRR7LHfHOC5VtpM4uol1S0Bg5hcNvLs4CN8Y2Ik+n9tRSga8fybQphOmqFxzz
Gir4U6nppQZjN3SnFIHcsFTiyWVq/30RMILMLNxZZu2J6X+pIJtQcK6DEvtUp7f+
SZp1yHfWXaKuSeCgj0GvJ8GmlYYTi9TDjJzThA13O4pzWBWUvdhNzCqlvUSnG675
xfkHIkJas1EASYw3EIqYMvvalrVKxfCDN8LQDPEBN4/ZE5sXyxP0XM0l9Hp1gXqm
yIqGwk62TXurql4R5UxRbzyn+b+ApP7wLRrfxQzzUduynv7T2AHIZlHyoGoveiig
`protect END_PROTECTED
