`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bWdCkGhBuSmpKaVapuQQUQcqxPtHsjGKPx2Jevr0LZ0jRENCJ8aXr9qt8l7lwWGU
Q2z9qGBg2ZeC4EThq1CfuH47+WSIJKGVyoedKh95vfkNW9y3y1fFAOe2RMPDeDSZ
6SEgDZ7Y3K1CzaWWXnusKMSvTFudPcmnzmqoQd4vBC+wCbW5l4PIG/Z1LmDywPdL
stdivqC7PdLLCjJZqg+UekyKIUq9Afp2M1Afo/h+9g0ukweUVeNI6ILd/PRwBhOW
tDP6wXsVwRx1mfOhU35HuA==
`protect END_PROTECTED
