`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3xpVK8t7UQQR3MayF/wFHGDoZLnYaxlberivljCDnn3BBCCl6J0HJACU8X5fjui
PRUMl5m2JzJ/P3geW6IDqrX6siHpYA4+Ci26LSTia824Z0Pk6pyZmZBhiX2+WX/i
6mbiP1SKZhAS9oLZbM9kgOlJozEZU6LY/39LUUr3zMHhuD8/kOjNIMOrYty5IAZQ
ajLx6/RUJnGuxxMreSiLUrukLPCsPLRu4q+RBGmfCQrS3oD7n6m63TGp1GQl7Rct
uspAeEkL215eYMGj6QTxk7UGiJBA8Dc7qvFIiMGyyL8TvVtnPOpajhuyKNtr5vdv
LbWCIX64hoQlrJEG0OQIM47ZS5HKvrNkhnKLFSEu996QBN0RYoSnLlQmlcS2EubF
Ai+h6sPps3K4yJG1Bo+TWuK7mpN7m9NaCR/mcN+e/7qfLvqU3btGjcYhc2yEKjVn
bqDy3UcsN+cpLLQDrL4nurSY+vT5x5Cq4Nme0K6dN6qruIcLVRKIJOgh2ygW7owG
`protect END_PROTECTED
