`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJNAfjo0XlfQ9lkL0xEfupGWi5HlZib+FIByEzTknD3CIPLuOK0o06BUmzgEH+2a
ZPTkmH2m4PUpQUl8ca83j8T41W74AJanLj+9UeVgULOJ5cQULLPufUHKsmOGBl1K
xsRgKg2fXEa5n/twOXNJSKKmliLpAf/WQTOp/Hr6Eb+uMHIdsqikJA3jalhA1hs4
8AN11SA6pRXN5thTiAXDPve2MJXEEKk3/cd27RL/fctB5VW+O/ok8ycPb7uh+gIg
Puq7aEZRMHao5c6r5It2YAPeuExBS20rWcsaMfmgtOaht7fHosi/9gj+Q69iiaHg
TJfpgM5EcBYaYbqNXlRaQsgzs8tm93HLwHWajr5hgic7TLrjlO5pDg4FbRPkvTum
PE7sm+bMJiS/d6MA8+TBQFhaoSRNok+LaEr2VDQyp6Kgn23xmbrcDL27aV4E9RzZ
lcAA4sw6CQ5puaefp8bC5vcFCjIZzqV7X32decyDtN+r2avWdNFRSta/LEFdM2pl
Ovk8NUpL+NYq5CHXsxkpmRJbJ0vIKuobx3Y6OgR3RjQDP3mV0DwN8PIqdkGNa0Op
hPJvqiX6r1Y2c0E/yACHTYcKmMBFEKAraah9wa/bCmXDHwXh2n0e5dJGvLRQjU8Y
yq8j5x45DQU/JmQMMmQBEnCNzLKVh7gnnuWJw5Lcm1dxJJSykF34Sf72cWPucIq1
MK4S54xuurxbm2G6IPMWKMyRsxvFkZ1S1QiEtqLBEWDLc2+XmTnisJIvoNq9lzVy
HgdrgdLA/gDlOidBBDGTrWmbfKqrYb4ED7lp26im+xlsnteO/5tB6zqFnMSruJXK
XjmddX4gWa8k9RKX6+agqQAdl1XZ0H4ehsWQfCHA5G0=
`protect END_PROTECTED
