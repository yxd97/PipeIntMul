`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3c2NcxGFPMYCe1MZjowGqHMS8/TkckZPKEKjFPXDEH4EK6Gsy5TLmR2wQzGDQJn
6aMvxlvGRgiRSfy6gwbvgWTN0wQmcCrMZeJhK9NeJl3saY1zMYQ0I3y2/GNhacZZ
zb+OMjixRz5Bel77G8dVUDz02R+QPTVumgzrhUJEbshOhVqpccjNDeKSrj5ahoNH
xCnC8W/pomdXiYWMTERXhFYEXUIz9crJGFJ1SM3kZHPQ0C4r+qbFq+b+CWh9DfvR
vhNLBsOnYyHyahs6aisRpOkfLaoeXzg02SdmjO1bMR7Pl66bAnJEJ+1danheVC7D
GI6bD3inTA1YTCNFEI93JdMDH87pndM0AuoqZWTz8u1PZSZOjb7AkFoqVC9JVj5B
PC2eRRx4Koe9Uzup0cOkHNzr+XKWmXPCzxyhxyoO1ZCtBR8O/OzRBryryamX59rq
67arTra84ORz84NMnpTn4TXRZJ3n4fVrcqc9lAOyUl60m5QueeUE8OT+Y35kUN+x
UWqJg90D+3QCHhGKS6lI1boYZeEWzG7giv5WZK91fvwiKDV7fsk9VZKkQq6qLSav
TdJuvFfqIif7FyHpuVWpbPs3zcxa0adrvZeKdG2mfMgDfWXP2U5MXL4uMQbvnJZJ
oNoRBenP8isGQO6JXqnjxACWfee8lJ0p/noARfwDia1ANoBJiubPpYpaTBf0t1yT
mCUkz0zLA0cWV6MwquF/VMtoBfz9SJFoUYauy3XWYosEffs7XviNPvw1pV2axWot
+T+GN0hZKBo7pY3KAdvnCg==
`protect END_PROTECTED
