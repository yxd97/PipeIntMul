`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJNqpn7dJbRmuiOKTq/2raCVchV8fYN9nn1eVz20eKonQzECIdDJlXsd7lfGn8r2
f3H3RJCqkkbPB9CD0u91CxSbjgb79WE9WgaKt4fGD0tWb8zs2KeV6xJKS3kl9g2c
g2rFQ9KVJUSlvw850ZVEqCIFWtICEt5Yn7Sj3XrPfb6PKnQUbfx77kzz1IblWETe
pJTkWQHWCGbca1ORJzvwGGE0tkf80PeQQlaRlZ7vfgXzo9axuw1A0Esvf9ka2OiE
abEUiogSw8GnZLdaNpQeGiYDIuX7VJq0NH+CcYhKzq9YUhjFlqEva63PXYoUNWqN
01cYpHTBVRBbcAKx1Ww7D//qzNOJyVN+nehW6ZNxEuVjT2Vdkcd4aUDCfUuokQVT
z13Y155Y0wXY2/ABocbFb+Dav4W2nde0bf9LbXdTbGbU1GTXOet5u4bh8pqX6yWj
UzhSPPYPylAo2/sWFCDp2dnAGq85TEJlc+6EX/0xNI69QA2YlNCdQ6hSo7TIRMv8
`protect END_PROTECTED
