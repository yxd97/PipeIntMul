`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7clYYf+HfYI+2borOeZl6v6qpKz3yaAoZzz6Q28HbuEVu3QO/3Rf5YoUpsaT6Na
Z0yyr7oXk+VpfGsbWJysBZoeDxWhcy0IoHMUY4H0NXWRdYTnXvJv0JPSu183vx8A
6+I3Kr+YnrV5nJ4pu/zkiKTMmjW4dMkBtTuyT6fivPwMi3OBK3AKZclvMYkCnhPB
+IBcidxudjeRWHVvloTT7i2PuEHxe4k+u2GP5yRdhWbHKR4ZU5NRgzvZqGY/+UqN
qZ6vLj+Eyc/qfEgDtFHXXWFfetf2QeEORwRJQhPv7sI/2j/FTnqIk5t4e9M/CxdK
G3ysKfVM2iRui2uLHnjOgXnieOhZMQpAMgYSA16VbxAjdRKUyHa9dl2rEwxtcHPw
+csUfppAI/KQj0AYnCWGdh88+0Dtzv/myF7VwTy29jgAZcYZkNHQLrKn5eY1KbQl
oRg/FjPpnORN0MpW//4vmEiHiFqc1fhUlTh7sVVNIutWm/8TGeXWCLiUAeVCOMZa
E2JRhnUk/mQAeI+CglkUsuMF4chhpjz5IcDhXarzdxxdoQuOJesAyAvzpt/qKdYr
hT5O7gp9Fz4jAqy2bwly4hJbkjSoNwbS+sEW0Uh0xJnE8QPMwoN2jfK9T2dPURHh
08Ycow1pGHaVBt3OPwIJ6rm7zvJx6rqF/OMmiFpKzTUo8njETePsL1/zQmMWSvkA
UFZ+qWN29SqODzNDHDti1V902tCXPvbNOcBGM+srsgtiPk2iMcMSBVYHBYODQGdO
sPjiCO15Q9cuSZ/WMcIXzN5MLdH6A9sr4AgMusLXBc5HDAWm7EsJ0C1eAlh9BtAR
vG0s3Q8419beYadn3H6a9Rkg9Qa8GgzgDtBCkyfmkA0yuMgdNOw7OU+GZFqz1i6Q
/usItUjyAeGDmojbja/oFPddL+0Ynl790lrPFJSpn2A=
`protect END_PROTECTED
