`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QderpZRNzeakC8tIuixpJtIOrP3ypjFD+hVoLaSV2176jKZgKQXGSLkTb8Al1efE
ntu/Kzy++ZcOOmYWPniZdQMX2eJjPzHadVbE9oo5tUuIN9Ehz+pAECps/lqhlHBA
ZdbiaX9APKYMAwixAzEzYt4OY1uTmT4m6A/cjskIXJ9b7XaBlMndDcJHbnlbiDRP
jCu3PBKjyWhJjrsdI/QM5DdyP4pQw5seMrlXXK5TQ9Vu70Wj/WayIfXH8ffZVu/r
zJvWQrlgMqlpJBiGOm52LQ==
`protect END_PROTECTED
