`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+1qbFWiF5eHgbeOJyiO82KsCh+OD9wo10w6S+IppDBfeXG3f6ToWdI5/HK14Uyc
OJHJtKvQ4TGc48Bz5EYVE57YmwwyztmQCKVzqDYV1nZuP1ouXqjWgHyDQWvrBTF3
ga9KrIZuYfkj+2UpdQHZUj3jeCg+h3rXx3hnborcwV4b8Z+OHbsW6jlcNW/yd4KT
xo5WpzgWHSv2VMqpKGE37G9VEV11nbe6RnOSQlF5ELKizwzqySEiiqS9kuFel0gh
QpWpkANetVA9CI0cowWIHL+ofh+ybOoGmvVUNrFEb+iEINSF1rl4Sf1pyTBfT3uR
6kX8aQHnmnyqb9ZtEzBl3sGmODLwKSqUk2AOrlQ36f7IdZGD0uQBU90YGzQc4fNa
KkT6Plxs7SNKHugT0RkvL22W/nt/OBYhMpraK0YWej1bYOjkEs/oiewpfCaDpABL
v6sxwnGpoxPOCdpkaHOUSbGBFL47CG0OKWq3M24jUxIZaSPIAMp4XYiJwithOk1j
HSWEkLad3UC7vzPlJdbdL1ZA4iYEtkWjCNA4gXf1053tST0rBMWiKZj/ODc/ueYV
MdskCmTw5QGj9V3WLi6XUghEBty16ZvoZjKeCgbEODA=
`protect END_PROTECTED
