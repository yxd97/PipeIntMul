`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukBN8dsYbW5kO2zao2QREFV3B2FAUkAJTZTHqwd3vLyTsXwaPuHg7b7hMpdpESr2
LY0lwL1GGqcHZnWxi76UyNoxoQY2FPk52XK7clBHmO1Ql+svJSmrK2lEh/ajxpjZ
fX7do0KyI9xAVbvEsY/qbUXZRFEoVPFm+6x94JE/3niWoHJV7xi0NtXB3R6LEsnT
BvNw1rmSYSoCZet/+EZigHvxQkW5+csHRVDNF7F9JuX6oLldxNLx69gEov57DAZq
m//2/EbIonlyE3Jrv1d/TPzK2F3OqOMR4dgqG5jS4d7GJnUoNzF2Ggcqg0mhNWp9
krtvDS0BQW0e9ENOIN7KIIA3vrXuwA+G4f4fNGNv7O8hkVnNUyRvAN3zuBrPWyjc
Ml30+6Gw9Vjc4/yVtcKW5UP53wRX7oJLkyNaSxjqJCBRN7w6PyAL2JCyXaP6bBIb
h9nYs8889FDXEhxnh056weiGUKJ+NHxfcvtk+a/N0t74TTU6Wle77Inuz14aRaes
nlFxhaTEvYQ04AsNWJ6v/WVsLphF6i9L2cDjaSQy6v+mZepnpsW2GLFX2dV25afc
7zRiZA4h93lfDdlpzcolNFD0ZH36HmQcssa3E6PQKMSX+bAPKdAzXyVS9jX9R2lQ
`protect END_PROTECTED
