`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zYSTcb++GsX+9Gm+C6KLyipSxQXB0CjBN/VAaR7uLdiUeXIz+mAhQJWoMcNS0eMV
jZQXHN95U2zOLOqO1hdMJQfamcuDPjqAvxe+tBU5GzFGBfUwQvkTi+GzGucw0VTT
ats9s4BNhmRB2SOYB/7RL0AXmb0A4xBSJwTdnYEKnF+FomDmAzt91h9MIeYBJ888
QDu9pm4kvubDrTyOwDywGTrQB83IX/cvdO7YtvHvOUflJxs3UIy0Hai4gVxWA0KW
FC9rTmvBqp7j8Hju01ps2sJWGgXn92Ai3Y5/nSEtD8VraeuaOVZKUkB1pL9DOYZq
vIzTVrPcy5hydWX/pPmcnTdUN3YKjsrShfYV3nKOw/ZqvAjpRvH9vhR1bHRq5zlc
jGj2m4exganEXbESthUym8BC5oV3w6GMoWfD/jmJGoACpuUQCumjBGY2ZV/cP3u8
dKSss1UVU0L+EezwVAd2i21QwMwJoYQbpLkBEr8PxAf3kTcS/eiqafEnj/UDBcfy
jyCKms7ZL61K9AlNTxbSKpJUSDTdFfUJqPLHvHE6HmFz5NTcsjwb9Cg824mcw4XG
fyiiO8RDZCmpFIGg72Gg4M2GyGN1XJPeNaHp+qAmpgq4n6Ljcvnf6UE/cKth7CIN
JGJubiOl79NDu3pm9XZuFq5tk0r0W3TrekADGGVFh6+diYmToXz0A2cPuwiK+D58
Mf4sAwGxLuQs0m0b3PY6GgUydKLNZ0yNTgz4glHG6J64h9S+95b3/ggPL/i9b498
sIQJb6Vr/8j7mKqczI3kzarXHqYrDmJlyZH1hGx94JFJyAH7VAXR1iAgY28RaFlR
qAEJZptsrkVuKJxwuCGK4lS2w9lt5S4crQn2Sa+utlcUIypf8k3SElmw5ZIgd9x2
v477vjc65gQh/FQnNRtmGfcCDBBQqosTDNnNad5b+Yo5A45X1HDN3QKkn1Mpiwz5
94OjWJamvmjdcklGanpGt0O4MI0rDNoFjJ3WbHGLaGXS2Wbfd5MnCBmiPWmds9pC
m/Bz/gxeCrpAeqZQiLgYHR1Vml5kWylHMuHp4bxuB8W7NJDi9QcHsovt58eGhHqh
PzV6BUvE9IKX4PMFQaHUEHFzwNVh+GrGk334RlwGRBHv2cB8LmQuQGzraG7GRFOC
sMR2oBG5CxAsWW9gWDPRTR9LCkfBGuJLUkWXxn6nrYyyCpwz5RlQbS03TKru/Apa
lHz/ltpgEZYdG9xI26pJJ9MOAyU+aGN080D0b7RGpWGyQWy54rNVBJEYqiDwJqvh
zv50UV4DOxLskXmVgiyvKiI1Nkx2PJaE5WiR3pnsWW9L6JfMVdVgYYv/cDsz2UPS
TqvVAl1zyVkXGYXdJ9udag7wh6pc150cUi49yWMT4wZ7RphE0IJF6itaz4i3wXPT
Kz/nRCKLT2n7Jtemsur+ZS7He/oHJ3gei/7y53fwFiYWuXOybqdeAa4Kr1K/FlSu
vPwLQ03Go0opaw3/GUoq5hfFLBoRMXEzFXdvNO2qUhYx5vzM3IEg5q+g0sR3XiFM
50RiYEuhINm4cIZlnqSXVP3uufR5Z+PZlPcUfRclID74vfM/YbAMmsgViQx2Q4qK
3slru/kJpUh55LsQ1Ch5VaPK2448AUVdRx+do1u3iTaJrVFwWCBK/J5WJZUItoCa
w/kxrag/Qw7OQcbOOXGlH/5w/islbBtOM0RtdL7/bAUcAx4PPeiuuuOwQt8gj+gN
btcdMnrXtzqjupajaUiQHVgIemnbQiqUzLtG4yapYsTZu2ALIkjAG7wGsemdKCDZ
eoA2X27fuBtfgOhkqXGV6XzWtImUkmGfjUCm+fht0vwaQdwjQV98pXJZWtWq8No0
UCfJTdZt7CT16EQSjlV9VoLs5VC062a04hcgiGBcbObA22Dx7/0BA5bAll1wTvvS
0Jr0ZgTpu+p/tVFsgjz4teHcnX/4Yghx1iDdAQpbYuaNCeEj9jLw6uzXpR0F0Xpz
hx/ELPUnqF8I1JHUqaw+Y/NGKWBlAwG409E3c8mEFZYUHqqbu6TYrKhziXLRfvM/
QlYJO9V5rd/w7iWJa6pua23u/PNVEJCtmQkAGqMpjm8zPjuJPxwr4SS2y0eJGnlL
s1VIN5x+1AAkCotuoSseLvVaPPekWCUKrtRqQPJdaLKM6yg/JDiady30w6fAAhSt
XImIn8iKQa63R2NR6Zlq8/0gm0z5qoQwuj4aFybtZSXAfj7zyjddf+xpuW1zbn72
YytNv4MyMaF973/nOJ6Vahaxe18vfdXG4V+RHADn2M6WY/V8c/NI/1ar9IhXJt2G
sH86Rf5qGw07T/DvyS0ZVYC/f65hAJUz0oQIpqhp/24qnIwF+tmnuLmHjXi++S0+
ICJkXDFjrU5CLVK9ehyEoOnzj849bFy7yD5puu0ghkV3J+olo263AtgqOSR35wP5
dFfik0im0x/7gv3DZqYN1F0cOhwbi41q4Q7ZFvW251b9aVYlZDL5qGnj5WYLw0cv
CQ7AoCRozTPmF2PyYIw4WOlPQRJWtQzW4YVAss5sUTdzzGEplnaCo3l6hiTP8ZWD
BI9jQfk01alLSCJ5ZLC8I3tKlOD4lkMlfxiL4N+Mlod75X481Twvu4q19wluPvWR
sAvDC8fwRyGWZ7CnyUwwNE+syO7LWWukJHEJq6rW2w+PaQnwJLwP//lV+kZrj+27
Z2qs91NhSW3d6JxyhcAA4Bkn9xUw4T4Ft/KyzPtbe8SBXRjNObzLMmG0OeZSsvrN
Q+uD1Mz3xRJggROBu3QfShYc/9CJbbtLdVhDVD3wg7j1EYVlTic6gW/6cnLchPhr
68AwxE5Wnb+IbO1i4sssTL9l777hJUxi7Vz8GAEWPzM/SQ0R9k1hhXAbfPH1MKPO
2rXbIivcnRZezdNQKdARGNVga5njvVtGUtzWFXHGlbZofwi8UEiuQKZMEriCsHeW
cSlLxz1+HalXg+IDd5xisSm6KhDHvtULZsVIwl3mHlq5eG+SNcBFjXiAhhypTY87
smog0HhuYN9vskydcqFqopp9wSwaBRJZKyWGWgg53CCMgkiwzvujhouRIQLqEibz
0j75CWgvFOTomSN6K5Nf/peR7RJ87Ed3xifLqiCl9es0cWmhUL2YBqGs0JmlojLg
fl7ScujDJOxL8RrBsFYF+6YcFNNm1YFnfKSpBaH+IGcSIFh/iXIhgUI0rsOP1TE7
Crwq32XPIe5fKvtrQBk1/Oxba8btdjfINC/Mm9C2SSWa+KEYgrB4uFV1797VyKUF
LwMgWvv3Vee9jzneCOViEmc1iJoybTYrVN1kSupSY2+Vjjvd0zDtErLSp1BfvlAr
qDoeh4XZeFxZvc36WgZPQ+H3/sdxTL2aQQRr7GPb7fHE47yYjs6XZlwnvoq/feMY
FT4z9A3/q2xHthULp5RFJc1gVg9fv/UezFhLLrQ/w8Nlt2mLgQGo/sEs9g4me9Fc
LaToRUkGfAZzkEqYb/zephpz1mqrTw99WN03eyA8dl6aEPDL1420p8l+xchaQt8S
f9i/KeoyCbTtwzkfj3rr6MG0/FWBhtnpuQ21GY9eHSvng2EV823ot0h58b3scc51
5I5MCK4wnX1fo9/WZghfufMFhJxbaxSGhODVH3rbHXuf7styP2HT3IE2pgr4ueAF
caqj0UljPiRNQPG+8FncxKJ/mV1vv+Al5EA2mJ88Slm0Cq5L70VEqc8ty8dscVVc
Wot80mY07/RvH5+1Ph5yw9dpDkB9nw+tV18HGYeXJrYBfMfkcqp0ZjUS/tbB7sT1
BJed/7qa33sUBJxWfK0u16+U1Pr8YBGmS/rQ1Hi/powQkKAqtGlO6AXIODeYF00/
PlBC81289sQ8Kvlq5okPyDmZ3+nf05uU3ZUpyxi00rCuGJ4lApGV6+l1IRPxKAKv
vUgCsLyxzcEP3rRU4z6drcWU7epCZqxR49Ri8p/nsXLoY8LmUU/Ua6wvISf9gb8l
jVIp9MQGaHnjCTa+eg5nbAizVN8h2V+Bax2p8+OzdVEumMcK5BPzUsiilH+PjF1e
pJtKGDkPk3+8QaoKjdWcRiBvviCg+n+oyqzRz+B9Unf41qXTBlm426jAT4OGL7Pz
CdzVSF7zWD8SDIYjQwxb+ImeO5/ugOz8QI0e4U7ZCMTodtHgn4znpbkFZr1VxmSv
9nFBm0zKepZtAIJGgQ+Db2C+dE4K7+6efpRPkjDu1KKjVwn1ImWo97tq0XiYLMrh
Oerx23dQ8H/+cSsRNp1oA0HciDRN1gux/3CIaBkiI9E37chXCVcj/NXFKlzebIDE
W8tPfVmZEM7CxrE607lWdrQQl5zunLNSBNJEtXoNjSaPgZiHiWPtvNn5WlEUb4f+
HpXqpJWqPmhsokx355BuSuj0kxt9KQPCVslrU2lA6fVeS8HlXqNhWkNeUSQz1J0a
D4/ELFieGFLmoSdLNd/asFEb2EFCC4UfXEYEkcGSjk3j22EfsWO+/pBSdlbUIW+d
sP7ggbTCn5WBY/Yj8NwdR2h9Tmx7m7g+zvWUqKodhGJ9ffNcx+oueAThsVg4W16s
K5mATK+M54YEliuLzDUJkoSK0kOqc7dDELBulb98dNEXgWwi5zfQNlIH3DyGNWuU
Zjr/bX6i510/BI0Rj+6G7T45ZKtwuBPx07ZJ6fquqAnF0pusEgZ1cgmQuLYSkATt
TSn2AHcYX1vrZNSsHvy5+TvytqSdGk14UORoT+wB+KUXWvZK6utFvFYmV4YU3TgK
k38Wf+MuncfAMUeHXmCw7T7p62ICppfmUc4h8fGCHsqk+BRPeAkF4zheM4AMNVJ2
zBODfRsp065HZ2uKRqPMvkda3IEbaj8vaz53/aT3X3zd0WD+6581oYIpjlhNW4Qn
Ff7svFYwlYF2vHovDgkmPbX7tvONGAdPBkCekgLGkhsF+gBqYm86PXKrIF5CHCJS
6eT9q0Dup8ZBlBOBONlaeE84eYTC37AH5xiHXxwreTTYXEIifc8kauXWjitdFxdh
ybH2uDE4sTouRE67UNhqjmOnkLgJ98IKRWtOwoNZEB/9KrP4h5WWEkve42mAuxdU
irV40WF8Vk3XUSgTFy9Mu8WfSb/mcG2PlrTCoZMyEibSPqRmQJhLT4aOWK7d3s7K
ZLbQZw5WNsiBccz1d3K0sqwd0FP5cp3KLqLS0MZaKBvN8N9uiqNHqjTQeQG91hJ6
+jH32K93/6A7JrGFs15szQsbFMDarSBlY4boQeO8+p7p9norm37TvcHcIBHfsWyw
NHmH/KB4VffSMG1EDnBlLKNaryKxeBcCZstET6OPSRu1Aa8uGR1aCkBzszLc1gMX
ZB+Mbl/St4rf1rx+ffx3JGbhufm4oe6ASWwyONlOORRqqJ1BvEaemmFXwcvb4bdi
SssH5V9vVDxfNkXSlYLsRbcxZ5A4O6Ce1DF4N8UXsDNjLCrBVkXDlJmy9oaa/xEw
Jjl3mWgDxQRa9ND+CgrXEYVQZDIX5hoJvzJfxYYSoLj33cv/YlJ5EALwh5F6hZCw
Ur5hVwU03jxaWfEKITFCEBugTBZOGZrIAtP+Gl5tqam3++kIjlzHSGa7Ey346HaZ
aQiCzMepvdwR6cHdi7Fo2b6i37jANz3BQMs3vMEbSSfayPs+qZYLd/M6uCCK3Gj+
N6/dSR08toaQuXSP2hZ6UUUUPg3zmS6TV9Twc1Y+JmdCFGr3kPzSrZ3t9AnlzhHY
6iW5bk+UrnSpZRy4E3IeoQbu1Bj2bDFQpU5e8+0kH9FfPjDz1sPPuGl3Cpb846Dv
uceOQXQMLkn3tc90DRT/Vm++nsjYGjqfF7SB7mB4KECLNYuNMTuoHVviEnvj1waJ
DhWhisdzMVHnLQbLrwGyh/mwXil4h20k77tXnTouJpa2Myrmw+SVQmJiVepf/Nxv
3cvQgDdBLDZY0prSDCEwvt64lld2nED6FnzEH8OK4T6WZ0FW3cyAYvwYcHgXHuM7
mGF4t7Hi+4qGoQENfheiZp2l66VWt8G3zbSnt0DgssJaKDdZmrS1YIehQgM80CCV
xsDP1cAShDKjiqrWhTeQ6fM2EyiMl4BqRBsVzgqaa9n2qpdA9SP2h69HdZhZ1OMK
RdWJ2fGb9GZqSW63HBVaKWOTNU0PWPMYI4J95DnVUgQoofb+c/uvDa7oqde4w4pv
ulsFFFiKWGNUYjXAFilAbpNw+p8A1bpdoJo20Rr/5iBlgPH9+gyW6LZ4jHIvOegn
eomsAaKkdg4Y55lsbzkbSvOevmdof7dcnPVWFFM10gMqfRiMTW3H5YO3dxdD0IoH
13MrYDDZ649ybcHuB3pZ4YHHY6Jp09zjsRmSrQpY2xzgLfvpL0n21Jwta4cgjf9C
boJUNdOtyS7w+bGCuXm4oJuZ/NeMboNxY8XhAhUh81IopA2dv1wqCWIyM1k80oJG
NsEZ1Q66IemkjBT+wFg4sWqtqr5szmOJTB/Ny/i3YaZ+PSpOjR9/wKE19S6IqTdh
K8GWJqzhjoc3zLEAgBsgKunejhXurJofzVfgPaN2kzdPBMN3by/uwPo9StCCTDTh
BqScj+FJJvAcqpcPkXf/4FGWohVDavB2XNOTrI/DI0t2j9dzhIkM99XmqhaXtAKr
B6w/qXcm3iktWrQtz657bKExLLyhdmdfiq7jfZhIrbQ2LjFy6Af6c4f08wGBmMow
+XPmkmcTquCoFXgiTan61x3Kf9buBW5CqTockHWgpokZqrYLT6w8Z4OX6VO2bOoc
3ximFD6EUzhptrlJDfMI1GHRD9bZg9x9tvtnmrVAdNUdYHZD0xLCNVwtBXQQMBpF
xtlQ2ghKKefcagGoj2UdpBQ+pRU9Y3llERdvzvQt6zpcjeVtzHQzEXmoInBjI5pv
TCFmWRcyRmvcz/FQ/XS6HYaiL5gC9dtXaTxGs4xmbmNwh39e4tJEfb9MyI6VM6zq
LhHv+f05jct00f9zgJ+8X6bgfrdE2uf7XH5qCORykv3F1nknk9fUE5YqORACsK8R
WdpK04AFJa4s9kyUGQiuAOgare0puSNSiiKjPfBrv/TmAVUYg/tlAZfhiIpFfnak
UdL7h1tyYcRzhqPQB+9KR0OyLPHa5eMOgfyOtfx/IoNksYOCkf2QUwW+vEzNQ06u
xmoMDVE+AmjOgeMSCzZyGAwyjO/oETAYypw7XXlK5UYDX0675yf7z6Pt6hLGhgJO
eOJyEPSO8jnyU5Rd/r/2mTcD6mDyzvyapdVSPHUHikd6RyK7PN0ygUa+V+q2XOyX
w+w6sWLLchIHAodYA6ZmwDr8JvOuKEmaQUlPCjpq4z9BVWCHQNJdN2p3XHng9NgS
St/9dYruu1mmwfSOZXh2+OXjcYXtFboATomtHalXXsaFsgR721Ppm7qLae9qMaVW
THAhzE88YEg75HYwpGHdLpoF/kyLUj4ZSjDdVVM/YkvBX5GTXcMLQ3PnpsGT0xjA
+hWiRLQvFipco4cIlTFi9uNpze37bITk0xqBRiC89ITHRxWypgaH3uwUaVqSsbF2
g6Mm26K0HmMniKFUYfdJR+pQCRCSpDUKNbUbxggrlcQvfqVPAo4/bBn+t/YCz3lU
blxOUr2iyL3rshch180KGU6fcWvdbanPH9cmOiNfec/P3l4X877POit9z8vmSmjz
CJU1+KQBGJzAPYGc1yP7cW17j7My7AV21LWELOFZqdCFR63KmtokqQTfBOreV1lS
u2EoJ3DJH/dcQn0ThgdLfwilqQrvEAYByjUl1oEymIxQSLutSFoCXBTy3D2N7Uq5
mS88LSh7cKycALfbrxrnTbmn0ITkp0E0C1NXPm/d0rgQ8aoVrQLQODAw+XnkrcE8
GfTXIaeRJIbdY6ivdKioTVVBeqDhhZFTwoYelFMeubCZ1+UobHVCrayjfq8mMOVT
Y1H+p1E0PKyxwEDkLVr7JenDuwldeU2xSXMNs66Nblyg43AW/TJqHY5PYF3JUOdF
JZZhfRPDLqNqLq0ntXIn++Tmx732N44y4o586Gq5BUJ69JIaA8FJpLiTGNY4Pq89
ZXB6VjWoT9j/06OKyl9OU43b8sW5xvvKcEF9aT4yomI3FQPyydtrKZuefFSGxfQT
Bi9tPfOsC0AjaLKrbCIMg04WCCfjBh0qF80ZYMiNiZULt4y02T/2iOaGtLtltf/+
SEOQghwWhwk3i15DAQvg6bgMpDuhj9ckXF5w5Xk5SeWOYu5SDCV+Mb4nGOO/QmzE
Ha8Y1UFu8+V52KZJkeuXbMcL6YzfPLDGWJSZ15et3hShuAh7Lz+PaQwSCNiyGWYB
fT77rvSMSUQMBOkfgz5MqOKTsY3UC0VwdK+e6PQb+sVU595pftxykcrMRBJZxshS
8wJYyEqHzBMNGaBUKcdCMwkAEOoVe3l4WgtyYvvXAnIdky1cerx9LQcYEmnNJCTx
qw6cg2VYzs2KiKbXFjJeZkiEJMb8bHYcM1d1i6fWC87dkxHiOsokXc5aXDD+RRPR
3HBmsD/5SGGbxVCHTowTTdDda+/oRELVVFKk/x9e3q2DboEygSlrjZYI8yXU1d63
8/3zKpM90DNPzhKYxBdrJI4sDH4YiV6JVDybsO0V3ZM5pU/oIJp8V/oDybjq2/kU
mjD3WivZhzqgMw5+b0mMy7k0hDRRsfjvoS0hpAAYPAlVn3+ImygpZU/bYjm3nz0b
6h1ycZ4iRWT0Yo6yhptOwVO0Fj6PkNaylvyoDaP+BA+IRiA3NxtWBH92ujYM8jqH
k8D0ADAPY8x+NWbQfT0CfG1TFLFehJizm1FKFfurQMtYMMjr9f3vX8KbdmGdK0Ez
PaJzwKNd8DDRebN/02lTHXE3F2dugyeQ1CJ1b/cBiJ63FvSfo+93f3CXATCpq+rW
DWL5vWP5IgK6AjQVI+q2hfDjiOQipNRuq1mWG5dGqlolxvcWkjQ68TSeJTrtU4rX
EkUhvOMLUTWP4EUhlnZ9lGdxzTh1Uag7W5ID22VO5rHzngQ634DPnqIMHuIaobyg
SrHVztfHdK0qQ+d76DANYe5XPChv5iFTI8ZXW8FW3BuCYjClnQGlfKAvLb5HiUP9
BUOqa87FGUrBWCZQLqiWog4BBouwzWFSjLZ3cLOs/7HS4jI8OBcvV9B+ueGhmlbJ
KTons2sNbLEqA3LwBuTqgCTBuN9STNYy7X58Ze9KX9MdiN1WaT+kY9jrztNwvByv
IYCX49WXEpAy10Iv8Ho+dcmpEsnxiral6KL+CwRAEoVFgzRIVFnpjcWqM5NmZTVL
DSDhVj/n/yfkHA95tmE+OedHOkPUKfpNlolk2kk94kvhacfgk4mrw8Z/DrTDjZVq
6y+jQ7NFxaqmFSogynRvq5mq5DTDQmisevRNCXlbMdgNa9JWFdSzy2lTQtK2atol
++C0edxLx/9hLGoHJJNlAIs8ddOHyiaqUf8uucXsFQ4Athk9ASTzf8shbT0b9qEz
X6+FsEPJhH7nWTt8MB/v35GRSbErfJf60gPNZPNY6zQwAJtcbnSle/qzBcgnQsfF
vODXjWB7hkZvBgMUXSmbejkRukJOinPN0spraGabzHAmNZeD4pHh5m8d2RWhKwDX
8ei0PWeIr7OAfTGoerwuli930Jlqnu3V2lsVsKS8wImw49MZn5ODTDzcwJrBqSFD
EJbJklOLjL4Ie7/QFvtfaAtSHFXoN8aLg3EcP99l7VrtzfzDcQf1n8tHxvf/kMGB
LkZ8TyA8PiwmC73JLDteQXSAol9NHf0OxqmsefRt5tHNMpWbrBiUWcWhiXW5N8Bg
jcvcGXFD9KQQkaRfA9Li/emPg1UfBaZgsyO+ZpwuhWUKtw/2p1o18ihdTQ7oFC1y
+WeLa00WuoLFnzYGxsU5hfOy9HbZY86eXENV7DkRc5RPZ87xlCG4MTL8HcIzvQBb
i4uiZ6ZJ7jjYsmjvB3Mj4/o5dgrhI3RGNunCRf2ePOYt7//M0xHhEyg2SkLBoS1L
e8YUWK4NjT7UHsUBRoHgRs+nE1QYDPuR+BISXVdzeywiKrthyssS/lGi0/Vya8y7
xngKwo8sUO+Fm91UXNf+uwuVEu3d6xSDyrOJkHKMrC1fVmpK6z08tmabl4aFWCdR
q19ZEZwQBYKRpkGnLB4ZnbdoFduUkqCyTGS53LGgzKfbvO9fQr8UG5vLnjXUnTnQ
hQFL+Tk3Ye01Om2tVincg2QqAOM5oimNyYSgrAqylcp5IkBkZBhgrK1LRx8etBw2
JyEqwXvLo1EHroBXUvcCZuHg/Wy+zuKIr7YdsVAJEYwGwZdECTDdsXSOAaUOJpW7
/x+jkqmgpyfWlkjeSYpIgvwMJpfnkdI+jvmh+Se90V3n7pQpyoEsuwR2+6cfkyCR
muMt8wnAkEs7NKzYxy8/r3U9BOREddvoo9siMeTGRhyZpOs+QL3KaYhxvU3519HI
xPDHIwBShyY2cJYTaTUhQpMxMzBWP7nbLf6QcF0UheZEv78jWiO8N2whzFj0SYbM
GNTBgS7tQJt70T3ZCsg4x/ILtye68SdE1T3j5B8rDRIXNjloWAnIj2zS/AcAEIYA
Swi6wU5q9w6oGzFPbp1scQGddKiBc32Hzw911u2rBDDoINB0RmJOItwGFNyl8FqP
hMnokvEm0EAl866qYzIaAKNbyS94mYPEy8hNJzhg9qN3WN08WKtOoOrw6ikLLIJL
YRkjncWnAiWJfQvRb2Vj9jiFPax0VM2cA38mh80zAuclnzDxp8n8vZ/ctR1Z0NuI
iDlNmRD+ul8uEBkxzI7PBGhJoHL/nHw6uCS+YkRD7CyX5NcOxF1AJH3Ks9bR+P+C
fZqmKWE59qX/0lneUWkcZDcrcJceXYl86z0pQWKSwqzJPN5rz8GMYRbdslkFZeOa
CKFAcK85yX9uWfP+NX5mQMIDJv9lHM4oWD7kxWMdKFmHdiQcZ6rnWM2bY2MAcQ5D
kNno4DJEWHu9AYO0QikQd0WwAn44zfB526pBxot7sDRBB7r/QIlhYl1hxjRprMCN
0CLzRHP1uzVuImyoip4xJRofuBnnR+9auQlgZhxlU5u+nldxjHX4JAOK/cFnoWyf
ybGL4I4ob2lTjBel9Lk2RcYXyaS/daCjmiKkKaV1O6pXYOy2bH2VWZn1AqdMFy7w
5Jx6mf1dig7mziSyTqjo8msEWn85wh5KhrAPiH26NL7B4pWdsC+Z2Z1S5Su5xkB9
6O/1VnTcT0Um0u35cNu0FNbABzlEoRmbtTnv/f8yjOIdFZc0YXGNP47L4JPUDLaO
OD6B4NBUprGB2PZf+/zpQFQvFTH31j2QtT2xjV5+mh8tiBmv76xhftq0dy5FOy8q
ljftFhKyB/wtmfHrji8qmkWSr2Qq2tDn8meM8nksbony8saFL/7JW4Rhgxv5eXDT
3vgrQwkGhHEdFuRQyNY2BkvGnkQvBqppTQQOWmt2U/DaIdxH+fID0IbxoTLO6TkB
mgLCe4TNafHnafeslXGafrLxg43J8TWFBBqq/nI0jSZkdENutJKxwMCFsfpfjjcO
8lCBWAfZkgzgURToWjQrHrTObIWBGouFUBloXJvV7olYcBWmNbMM5/Q7ArepTQ2k
NX+vG8axZqeQeP0KRvFS7trU0julapl290RIMxszaawMKsiSi5dPP54sI8EpT4yA
dwRfXP58rkyKoy1H8p9wt7emf9rXUHjpWAHFOvCg5XG//PQ5mTJJd7ebSfSqZe6n
9VFpJVHJaess8cR572kZ4X/YqFhFMO07a0B1hecmIQP8UcyM/Mh2QFF+xkDLLMIJ
syc3Hj/ndxWqyYZBqXsoupruj2qZR4dUnxXbjZmwwn1Hgr4rkhqSdFvjzG6R1gC3
v7Ud2+YXOhPdr9FIKTcK5FIM/qLdR3fPcqg8MS2LXwOxOaYrgIUsTSWXv4W8n7xX
IiGluyf8cVvGc0CZyvFYcWTrbEVdfkgFfqS7jBPaPLjlYM1akHwcINrAQaJGAo4f
EBTF97CHQbi4X+MNYB20UUYS3rzj9Y5nJQnmbYANNF100jqsreqW9RwVkQQcAPC6
1RcMCXL7jsStOTmnWUNpOoLnhGG5bGgz1SShpAWFGrwfGmsbjPRQYrM1LpqCvKcm
ieGMtNSh1rNsW3Z+jrffDTMb6H+QNJAKB2/oF6AbCOi5tCzwpjNAj+3OuN3sxxIX
FpkRy6eScOjo3hC+/Z7NG6YjO9F26MJdGNQP/1m6b8hJechjUjpzTS6Wp696WiMQ
96Nn1nepYT+1DPkLniLGSQKA3aAUS1KoDwauB0Pg09+tejNLH4d666Pyn104ITUX
WVBdAxYHdf6dGBMZkwiAzGy06lR7oXPMgVajIm5WH/zo2HLc9s7oj772heb++7PI
bodTr0P+qoAYNwgnS1mn8QtHD9AAf57hXYN1FDwOMAW5twfhaEgjpc+eakXuDiKp
XnFO+XtgMEk1RRpXDDwj8KXZtnfSibSriWjX4q9S/H0Gqr4C4Dx+CdIHPMwXlT2q
9ONmipgzH6Vo7QYiQNLT9Sn7Pthm66eexbAXHflpk/x/uQxGCOYq5LNg0wEerLq+
RhZdyXiJuFE5r7lsXzxBagoywJ5XhmTsATqo4O5fmqLxDiqNzCCiz7iAu4iWYQ0S
Ovg3Tcdp786cBik819Is/RpcfEydBIJM8P4+KCyTXf29Uzfq3bP7kAQLFOMMdJp5
60ICVy/s7w+nFqOKRB3iVTiJMgAIf9r2iOmxKKJ2tjCrbMmsQYu7AdyS4XRGrIeL
42EtRNfitvQjHeZUnSn0NpzwfQm6BrsLjMMiRJ4OkTJH2utcj5XdtZAXxrGvT0AH
/ISNLbATtNqgLDjgsgvgIyPth+Rd24bVKs137L1x/VQMuqTuWegbo9MBREBH/mvi
ziBUlWIrUvL6APJFiUMZdjye/vL0oP6gSnuyCPrNr6sv5GdTdQk7sJHSVRpjK/Na
r14CMItE2ITRCdg2XavbqOT607TXgJtfVlbNrthfjBrZUd4DP/BtKc64o8hZl0w1
bZe4PlS/35utTlX+0U5G+SknEhYR048YcG4eNDoRWy0UQKOsL2yT2pkCKgi5oGTR
tvv/L+pU5Sq9hG3V5CsCKvGSDeIDdudfPZ13jP+VgbZLe7ACgDcPquc3gtxQZ272
gqHLf0WIk9IAlQY4rC/Ax41owYhUvTAEVcmAwG7TBNimo+EkIDcVF29fx7jeiIU5
YR5zbg8pRbyCFmm0i4v1nS4YG0cbyjEIZQhbx0FtCIoqI3L9q23TJDvRnXqMwNxg
9Poi7DA13pt/yN/XX9sZH8CyN8oLNaSciCJu+gKab9SzS5S++ebIQessy6w+AM8U
/UledE7ThAPXfoQoEQ7qUwMRO09VAxyB3VP2Vyol6x1GflWCP/odV3vCBy8ipmVZ
6Mr7BqZclz9Ty3jmNX4kOAyqT32keu5Xns8b+q18OuNAfTjwTZaPt2CWgOo2nEKF
rkNGx07VWooiX8U408ddo6QHeHe+6BMIXru+MohCQ5HeERzc6enbU0Jja0xwzVuR
SvAgACIwiDhrpf5BGJUvvW8i9ZD2q5v5SoFOWtuL+mRQCTAVDy+hVvSQ9On2RNqI
Z0G6Ou0nMzyFJVBFWVn/lanxxzuTS10zZs7/uHuQDRi/sPVbf4leZUuGepc1xhw5
ZNmoM7tMcYz8/wRMbekk7a0RxFJ0Jd6IgwlWCJpEli2VEO0CJ5bWBaJudlIKsJ6x
6ADk1FDnOsdvLxeoKUNuxcD/w7GWuXESZKdVC8cyr8vzQsE/mhaRoev40SBlI9vD
7fBewnPwAESnFc3R5J14/Xlzgbs29r4wWZHEceisG4CmZ243zeUP7gsTWVMYH+UW
fLOfW2YKjjZ+FoslO3PXg1onbtlg2OwXkSKVjUSMsp3e29Oqo+0vTC1yAImsE6aO
MTmEHrAdvs7qV58gzC6MpxCG9LH29+myhOxI0MeKZPtjbJV/iKSkGUQY5mhuUpKB
abw6E7fqVaTuvcZFjKLyBLBEBGFw79KHCcLCRg27fN6i0ypsJfW9x3gPCzIvmA8B
dkSlE88W6A5elJ2vBPcrmfYMKlj26KiOIWXjZax8WoMccOOKaQbxffY8rrzY3pI7
wiyYkm5EgtOlvnhlwkuQaSIP3QcSQYPHh6wFEasZ76wX3rmfdECfntxeYxYhyYZd
OTwCYRGyOY1FU9zCXlxj5KDH1yA3R1Se+GW6dQ7Fl3HGbJ23Nvp8v8wZ/9cnqXYt
OKMokNFLOE3XbWW9GFvVv6+u4zq1bPXRP/sDeozNEZdjplWQAw0OydHSvpI3UsSU
WkCSNShiZm1Mcgqxdlj0pDwZiUi7hXp9pvo4AzyGoZSStLcT1Ox7YAAlPbABoZZ4
yIOVFnoQerJgoCi74zM7qZp8wCFrvg7Zyi/gpgylBG0YoKFEzHfsatrSjZLdvRu9
1x+mNSXFEOfgslttp1HqrOSd7z3FXnveQI45txBcRqBAeXbnRNpUOiURQBvtON9J
3z+W9OstOEMBTN4BjhxpyVPw6wAWGzGuBmfZ2KKdeNofFgVscfY55RVdGi01Z3Ok
144oQt+K7aUQWU34Lml+PwpjLeY2SpT6/WSRYJtsCq4XoklpT19rA948w+U5SzoQ
yGnPPB5BrVQhC3PDo5vK+72JK46yRaBd3T335CyDIwOxWejJoJxZVoZU0t1Pv4BJ
5bHwWQNc2uo0To0jPbveHxUoEY78umNE8/0rC3kbbvH/IAx3rO59OtDL2wzmulu6
LBUMVKvIMnNVqBp7mqY7Ke7DrCi60NS5+1SHs4gg+K7tQZEGlbOktbZAr+WlpeUH
11vZpjo6j8dBpMziD9WqBOg+ftitbNO4q2W4O57PlP+RJnEooCmsE3HtuV/cJeFn
cEO9cRhVpomvYZwH2cif1cMi6YHVZTH85wZNHNaIZe+4IyOdpm8qbd88DcMeSgbl
wrj2gW/tq5vtFlHmwx5GQBeZKg1Fb9Yf+gjl/YGWPDgBQfzPQjB0Gvz55mAeltJF
1oYkWdD15jUOQxjDVouqFpRAgdr8XDB1XdnPlP0xWFAlRnlmvVb7qGKIlrAXHwF6
hd2azNbWIitVsJTH7uYEqqh+idRYDXf3Dqq3ZOKYOikWpjbXs/wYDn4B2Ni+F3eu
Ek+OPgFXKUUX7vV0M9kdu77k7LOp+m7aOp+pIw+A+X6tdc75RULwl/krqAJ2tQfL
Xiy+fCxRgvhr0SZuqJZLqpt8lEUA2+l93pp5/YxoL4bCK9DcJZgCBnpuSfm3XKun
ZweR6wMasOQS+BxRacU424SueMRVjq8fU+HMPQS5hwLw8UHh5TaoBJleMvrfN/NN
9LQltRLoi67pstRvpp3ATjnei8WihQoj4GTghaUz1UiiJi5ZB3hebRAB0beh9RLO
JWcHq/1+DBnKdsxmu+5V2oZ1XpdMgOaWPK7sOGPnP28satnqY4Bt8J8ccJFkYYvZ
2YAsShfY8S/m4lTLSExV/CACRES8zhOjIuQIdu7upnTty7jZjzgmft8rvWn+Jd+5
z0Ve+ic+FypzD5v+81PjPpSUK10aQpJOPvdqUnLgYDmSNNR7DHsRjx93RtvL3n6h
a0RyZp6aMwACeMtdsVBwkqMfe/lSVjrQMmyw5f6PWa/yN0q/v8RLCuIIVd41ifMH
Y54XuDIlFf+Sm2ZFso0AVCK1qIB3E/Qqoh1EWKHs8bqR+9c622JU6iYaVREYy1aw
/8UTGaSmty+PbhKU1s9uHyluRg2cOycSXb9bNIgL39YzVoEVtgxGP2TiH6vqPpPB
tkvx0+99d8J67eBq+TJXDJRHjDwiWXek1gNQ9tRcmYa7YiIK7H2WA5Wtku41CcIy
ygNiF3QDmte1TlPg+lA33TyZHpieyYIeOjZxprE2MP7UBQevlnWfqZya+wPRsJtc
xfuQyAnOEmHY1uGZZ/+6bE8X99HnnCIrx6tE2becNrSWBEUjvnOO5sKMP59GI12f
7bcWj+RxxyIUyZqpnU3jGsvw5ICNBxFyWzgPEi0SWyQS/V3BHFCntrAIj/LKYBQw
Nj0Id+9Rvk6Ondpy2ZkxcXQV14dm9obUac2YY9HoRJ/tnRa7reMF+uzyrD5EWTQC
5IO8/RqLj7LVV1AkCpnZGKXhhn4pDs475G7pKancOLw0W8UyDSXP6GC1hTnZ2qxo
xgQ5gS+/onPy+K+lKIql65G/xShjEggm7vIQXR2hIit1HtDzwMMkMsk8baMVE2kO
jPKJqwT+C8vVleyv64yaI0QITERJbv9LgxWnB32/vx1gfvXWEToux/gWMmclYAfS
aHk7bEr1E17On64jxECQcITMjAcZrbfbCiVjOvM7soAjTfnsgu2HACODr5l3mQVF
qojE5706LIanQq7TiSgcFPHGyKza6q9EW43tWeRprOLujOhz2dcdA1QZttHncBoX
LqoQzNFC9JcVYFL46fk/wWQmnoNP1EpHgnX3Kgj6yLdR3dABHuZCYGZp/lKZiHFA
qrx+QYFCuNqKNsangymBLtLuTmc7rhiXu+V+yDMJ8KPYZ/JgH92r6XDFmKYmNGzf
H1n2eCmlNa5TBGIpG8b4TmDSza2E87z6c1jX0BkMhe5IbwJiiGk2ARxGiByUYtL9
9t3N28oXWx6QMY8TgcW+W+CP1VYEet/4v0Vg0kg4erP6w7C0PIrcuju9LowiS+hY
kEsyHLAZx04O3ZZMvP5WMNsBx/NJFlibguZeEKrb4iTAeKKG16zmI+EhBKxGPytZ
58/HFFaCufcWB8ODG/2A+VtbEGVCGa746mpNj9xGXqBrv/+7CSojuqVAxnnzqgSG
cSzPfViw0/mmUXkLQDBdKSNMK5QB8p2bgzLc7AuUMZcSiFVrGpUILs9uyLgZgRHy
7hsAZQb9b/frBTng89NjPSvhn7zJZm+lddMa+NLpdxB+GByRKi1YtWXcJFr8I3Gx
M+v5YLp836fb2a6muzwLtFOwfpRUzM36Mov8LUFqi7PU0FRQbfXj+FwYCM+3xPNA
Gk1iicjXq2VwRs/zYEgaVD6MSIAtrvXA8CLeWYqJkt3CIqHHNTQGWGHkXclZ8KT4
aSSfliwMewDlU64EcOc1+T+wEOKv43+KImFuCoZnj5Bb9BcBznOthS1zEwM24OG1
r5wpyWSpYkprs6No2B2ua7uGHmMsehXt8oHyvOvxtP0Gg9MxhfOrlPhDEq//+qYk
lPz7yvVZ7EKE5osqzW6HbOwuypxOPQN4oD4WlV5KZ3uBhdeCwRyBDvNSA2ggdJ13
W+0akJUjWwUr4HYHqiCMZKmN9g8drF+vnCMlWWN4y0NvzakMiB1o63tgN0LMhXmE
Kg8CfYxURoEDuwkrYq2ARNpVdn4R6X6k4JrYclYitbnesceckKI+O8VeLWlimafI
n5BwmpE6TVg5JNLKEXZ81YwBi7aqeAaeDs401AzpWLqsJFDO2l/wchk7JAk+0Wl7
hPLQdu8P9Zy6lCqC5yxEadmXR6x7DnzWr2sUpB4LbcQ6gXvON/2DRl0jEQVmKQad
3HzleOkYxKm8ZPRlrvFz6VmAqR1gS524PcXA2h9+yzCM7sKyvp6RWUHtVAL4uoTb
KTMIm7D9VKoFUZGnE1+KbO2xTMdY1b9D4weQRVPuO55wEUREv5a2osPWxbnO3SWi
hJAc+k3KFFr4oW5AbXr0Js/SpsSmAnQgdtIdK9bNrpk9DPcARJ9JLGgmqz5+0Oa8
fQhDixE/faSM3u1PEfiI37ZrXKPW2godXGjvInU0u4917N9zYG3x1jXD6uAKs4+A
Z8eTUkB2T36wI0gnc0foUAGoKBsTilK0Vj1Zw48b96bMOPSLqRHFFM8pbPe0Pqaz
MIVQpIDd2e8LLy2ohiNQqJ4vRtH51OmYQrF+zZUvx+C/O2XpYb5C4o+NQXfIrDhJ
dW6whAKJ+GTXYI+kJXWwOlNU2Z/5MSDfonJbHQNzjQiR22YCse4rZ25qMpRKCA1T
KXvzm9u0Ug71aguVyO+VuUyey9akTqijfqJTeE3j1SoKUg9GnzMLapfca0Dlfm+V
KtKCs1THmONRxxLMdDlRuOC/L3OuTAGEstoWGvjgHL8K8zjvHhAf7O8E4ivIuAcV
GRPhrb0KX9GITb35NamRoHAwnp03FJj0udUGZHt1pMckY4Koto1ez4EPvkibw6jm
VgvI8SlHW33ISF9Ye6zmXMzifgz2zN9DgTjPFYmIe4R3HDNRJkHLh2Wx/UOVwhN4
KNbUzbuLX8O6WWYDoJoC9cdpua7V8jGm3KUVJg4uVouEzSu0sk83mI9Ort8KjfpQ
7eZrd5gAJV5RtZ4Ou1NOTnLI1ekVFSW/lfTRaDRzeAV9Y/GVx3sLnJCeZUzIK/ID
UBYzM/hpJWQMfkuOxVIGLUkKoJwDccuNNMCjKfvKU0GKZF4V9Cktr72vn9zlLAI6
4W0cfQSCPbY3i4KeWolNaW1WA/b4+9Kp4dLxx0fdhBLgl8UERveqq2pCRS+WiOX0
vhJOqIdYOTXkvuoAtuRC7FYjV1SZx17Y+cMMihVWvM6+jKLCjje6p/umunsTtdei
uWbTvlERp8RpRpXuJsKhvc0aSTeFVEpM05N9ugjUzSKCH/3f0d8mDz6DXgu76LBb
w78rsQN3O3lmXlu/tJr0bbi6LuqbVtrpWuiqmFhr5OecaNwQWh0cWZdZkQm8PCam
S7CYsRJzi3F4pseJWiWQkGhcxFAt2IyHjGfkwa0sfjtKwgeMVi+filNYEOK8ZhqR
jw6PmCNTSCeo1OKmr7uOy0sH8GsHXrJUwEZtfxHy68pvE9eFjaiowqoVU6oDbhRP
vDVeUFwa7X+IDAFI31y5YRONCgr4HUPIFutDbRYy6CSE3G84yTIx+OcEQqmBQ4G9
rWtpC8kj05wF+2AEe+dnW/O1TYD72Ef+NwgEQcb9aThlmeWOMagONXEwVRzCcqoN
K7DTk2YkqFvSpwL+HtloB4Vh3F+05dd4UGy/AnI67Tb+VmaIvkXgq4hcfkdAsTz3
C7bbtDTIP8l/3Q3pNBuOEKCVxTi5uJtmfxak4Tbs2iRtoZgeKpt3wz4qAHj3lHPb
GXiJRBZ/20EHv/LElPP53HYJn6C6DN7IE1+KDmLBxuIDSN6N0rGu7fBA3RcOw2yf
FXA4fXKS/YSsrkyJOeYya5mu6we5T142ZEZ4IEVKDB9d9MnDxqnF1MLA0mDTWEIp
Cletw0IApIWBh+4OE4Xa3TnEp95EpTDHrdIAOw4z8iFKBMV34i/Q5xNpFbY/o4z7
eIN+SSDglKynQzuns7K8TGisDyGNCh14enNCiceL2X5a3A5ZLVpn7hpO+CFGKNDx
YgEo2t3/8Q3BN5dWXWrnQlMw/Eg4wXa0Aw8UReSV2NxtFe863M9fuWLrtCpNlFwJ
9GyR4MrqiKvk9k/tvbYNwk3F/kWSuOPEdoZoSYmBE16ZthEfKQ0wcdN0MSwN/I1x
9fGkX7nUhzrbZMof14wKzcG3T0QE5ZM24Rm4yLCW+GToSA5aM7mP00qggXA+6XD1
0CyAT6cdDzM30wE2rwH4g4CRMLqGqGp5uwlYwQQFH2iecadircPmfWFc+lyChVD4
s+93wn3TRB3es+hvrNKs5OcXrbIqbdlr2JfoQNszu5fvzGAhISNek6opxtYzFvab
VxGadbd3M0V98S1TFzD4nN1WMl6sPSKe2awMVBqPPSY1Idi/jQRPKn0N+AnbQgmv
NyhpmYLJ53CjAaLEjP1FEXBXO20QmkjCKJUh9PN+97MvmwP00dF5XQQ5HO7uYbum
/Ky7loRG2nfAVsq9sXnhWbxXT+5XW86fj187kJWIfWvi936dNSFw2tF5B1qKx41b
tCahHmWx32ApabIhfqpaABSS9ICvJy66B8QCPioX+DkUF6QZ9RDV5lTYCg2ADLFV
s5MSpkWRAxdzT3Q7cF+MBi0ZqBGHppzKlC3n/YxrqZNIA0FDXSnb5qa+9GFMb8iI
fkR/c4pmGF1maPnySPzrM0yccn6FZJuqeQPVzkUaixvi3aQ5G/an8tcHohrequuV
qPFRh0HKbuB6EbDJ1timp+HefYYY2mO5T7Y/o19QT5En5IhsqqBBu78FabOLoJAd
RjNMHjX1EQEptByXog7W08IIBm9JB/ISADzTmHE4HmCyM0GtWZlQWjrQ4HYVDjCe
8aWk2qFgmXq+XDrn2tglgbF3ss9X765/1ZM+QShd9pifnA3t8VDxSkrylUKuPbza
z9FhybQVSWrY+vWnWCHC+fiU0D4z7Jux0LvgpJ0Jmm/CRhNMPBxshX89s+jnk14M
fzfKYlVBMkQ5SsDvcsx0brq/n3mK5HC8Pg0caNV40Tx3adVhjNtOiV8rgDrj0w8F
sAyw7+WbQhgrjYetd48xH6ZUITAK45dQevY4eeOFTf9TkHUdBEbhJiksQ7n83Vqh
gyv6CSXdK0TBoAbiTNSF3LmD5gxOj5lKea7bjj4i5tEVajkLKDucG/RfkfOfhJGD
I49hduIW5INrXEgZMmHlPfArOoh7J6JKIcigG+KgSyRPmmg+yqBfqsjXYsLvVfDJ
H4bjsDFCmUYMpLjvRnfxWrCoEosdC/Z2eeWYaVT3fBXxI8nEzPGZzJsgBS8U3OEe
liS9KUQ9N6yGHwO5XqBMAvPiKKIqxEygnmYnBcQCiwtex96chcjFkdykdCGg2jYB
kNElx6bDsVFisNY+b9e/61ZPqldxyXUR3AHiR0v8PrAMoAVOR3gcInWu3Bz2t9Fr
PVjWR6nZlk7f3hQaW44vOw4NSGb1aHSUMRm/8yjvWEcYjLzXCzdjX8J9bcbRdG69
N0fE/nCcO4atOOllrwXDYIITDOuKWVYAAMtwO4xyZzdAHTLzx20+o2o+Nuem4oWV
BtV3SZepCREy+29U2jNhtXpdu8AvBsNb0ou403lldOIZNtwZENDcLKQTSr1NzqJL
n/ycTdQMLHMNoWIBOoD5qnx8Wv/WaVJ5rmeyoU3VsMhHHMYCNulPLW+EvduAmnOG
CvFi6MS/EN6qNqgjCz7xJ7VrkROy+KxKDCagtseSF31vNk+T66LlG8HnjutRzb3s
bpmBq0nqvK0Pgq7+8gm4D88csPxm73az6sefi3p2d91+0AetW22EiNcwl+pzUUDh
dm1sEuNL/6tstK1dOmRcKo1q7fmhdS6O1GQU7M+pCoQC6vRQtFJfjiEZ6N8R128b
l8/P+oPgy82NEHoBOUgkdF0ZcfASyZiaWvJkX1k29hUZDin45mKzD0XI0m3wp9sS
GvKM0jPVfQeHBfGHuNbi3Sq3Tuuf7cuk9/0LahF4LSEL0YQ2t628/o+VVyoUB/+g
4YmOZL1iU3pKaDBxBhSKY7eVTgtaBt49Dffuo4ykscRq/4pLpc+06QbwKfnJ3DOr
uwC5YVwswsKmQuR19p7IxkxHcXhnt2bTOdgae7MsWjWaNFsj/KlJikETTbDzeM8t
se7QKhgS7gYNTAhE7BW18yeqyLjsg91bo77VMf8V4hsqaj+gAuRsy69g1iEj4zvL
M6bWrocNrbKRhBfuUgEByfcCDhgZXBtrYMwRBpCXc533Vhhtcga5e3rL6XCH+Tbl
WTpkFl7LynsvbUtMeFHA5rmB8Ba5bvtNOwbXB88O4IblxUrfxLwZ/m93G9ZT4+eL
jaCggFQGy4Clzz3JaCTH4DxlHOExX+VWElcSu0ATBXHHHAUilgP20Ub3Gra1gUz4
NHBFkHrnaLGdTVhxqiwfXgdUmELf2nMV2if2Ne+24duCJzQCgMdrgPQtrHJ1QNOE
0GF+P3jCicV789xSYzlzerzWKZnuvZj5JV0IrhP7ywlOiEWvZcT2IDbPT4h6QW6+
v6rOVi4zZcTLCt133VwkCBH44NjdgpJ+i2Ghj578Oljax/w9GUq7IRpPoNBOzaGd
Vr4gXrMKfZ5opD5AqNOMjaWF2FfpgDONZUd+0KgWQshtqO9ygbH6cRzTRC7/L4tK
dW1VITDjCIVuB2f1k8heAydProMZowFp8Va38tMnj9zHMIRngaDOQ7YiqOgIOEL0
19LPwnDzPVu6sE3DdwOa313etEaTvQ80QVLc8fp9FHsTFen1XoaYy9eRD2PhwKvF
t8uCAZJaTJS8PDazmopi3MCtCN/zU7DhHvzjzIA714MWsRZG6k4NMqq9nbk+Ru8h
hrTdOHxd7GOEnZ1NwxGpP2j8o1EtaeSFJBgaBByQ7JJY/IRSDzaNK3fcEPo01jb1
NEelKFX/PrYokNTW5ZmIxwnx6h905EHP3yoIc1bUirsPmI1GwMBv70+DEErW4aJb
EhLn9j7cmkF5J372K0P4EaIxmniE+OQthzdKQTuzozRHhC0WLcT5B1F+FW/2VZVM
rqG8sPd1opISSCpq3+HnyvGKUoVvNeTkOXUThy4J5q/fJvBiFA4Eumn+8DPMsGu4
EeSvC4+j46vWwIesjFKOqeOSrVY/U3GML7JFZpk4z4HYijgEBae4+zvwN78ur1iY
FVhu04/uGIz/mAYlx4It0+X5k6iDfvzfekTxF5+HxmpOjbHgkiKfYil4x9aYsGxC
1v2bLfKfNTdg2KnE5xjsttdJFWEJGQmydX59J/M51APYGGhv9IGvR1NvB28xPUiK
zYbOPI5J45y7kCkc7Q/7rPiUtV9DwKYg1ZlSJ7HeePtkBEjwa1+bPMV/OvE62NEl
GLBij0fYic2bbpAcnUdNipXbrnM6YC5eUnVrxu1G1VzZCtsjDifqfrHTnwtc2nUl
L+S9xrVxKqpLzTTiVm4WFddN0nKdBunLFiiSSisujGxPq6kSdwmzddnfCGk4G8S9
qNW/WUncwp8/l8U+N4eQ59kiVA4ZLQvHMuhZRSWjQLBBmM48/Er3G/JtJ+mfeI2U
1/x8aO6eRHk7y1/4QVT3wwIP9ESIXY5w277U3p0P3qaU8UqF+TfcjqYDasEhXb0D
s+2OTGdNyCQUmsaYBDehRbfJdPRyxA2eSFP83Ub95KxiEZsw/d6gUJjbBEb3obfI
K98ZcGBWuAX1hAyTG91WbIW5P9F+zq5200hKconOXHrmpCpZuAwALjCNu+6I4bA0
o5qBcLDe+nNJ3FwarVj+uJqyo7Q88f157W4ZZMlXKudHdWxD2/HxRsdcT4DumeJt
9UgpBi/b8SE1rN5GXMkDDNLejZvevyfScdoihuXf5y6E0rvjE+ubiPJRpwaXI1+/
aFGXzifpt08ck9hg4yph8Kc/Tkxqp5m1MNybIS8Ssi0LmBX5DiRG8s5Z2wrs5uz4
ljUuN1UqLgvvT5Qs4XQthcYrOOpSOGbSTokVX6/tv0wS6ouDnemg4U67j3bdDkJG
AGIRf81VnpczLA/F24bWFCDpeoUvSMmxyDETZJaQOHevltMy0pBI4eR6jX/Ewy+N
Gf40iGzm2hoGwfNsCIZoW5GrHt3mrKKQIdUwOlN/S5n6SBb73jEQzdAVnkIVE7jH
jy2CBnQ2IeBDGIVg5EEcou+r5CeGb2zdkDkU0mFTlkyBK256EkngP3bwsjPG1qei
oTjQy3/9hTBEMQ863ePlxIf7lwC5FKSYJBR94nGOztZ3SHQycg40L7OGNs/bJU/g
cQw2bIIr1LrMsK+/HjPfb6z2Rm4Nrlew8RNuXD+4iPorUTbm0+D0Q/7lFs5oVdXh
FTQ+6vAho26Y2bIlFpdsoBthj23ut2sP51dL18gZ8fYAFichKHocCJ4YpEeCdRJX
ZBAsOSg7VmpazH1Ex6vTJ6vnwSsMwBu7UgjX5PqBCDhoE23B/w9QvSFne25cf/WF
8PiK/FtEtSMvTgQr/ZHj/iuc9/noLsRGtt8qoaobzDR5xMnXFmSfYxpIWBRvIYuw
D0gmXE1iPx6Y2TIZRf2TQv4WqJhSjy7/TEBHgWNljYc+Jn9mIjjFuaWV5gyES9wV
LG9+vRB8ZnVuJ7NRClFI5Igr2LiX59bFO8vQAR4IFrskCyJnlK2S+ppY9G5npLqx
eHXfzSCxhXvucUyeQMjKEI3JJNaL3Gd75jI/qCRo8jYUtS/MAG1Kil2pTLOqNyoT
NpkAM5fIxsgMnhnn3wly99clcXtrHsXLkeCxJaxbpJlkGcQU+MCQrkhVMeTabJ9h
B+E/1JG+bz/jO1vOS3NnMpfFgP6XjbZRrLP9ekg+mk8gHzfjNrm628bod7kenusk
fXj+hYzzldbqAKqRLnuh5Q5LG3mMRGMbtZtxgitFVOrFz2m1J9F18UU5cyZLONgt
BKAulCPcUT/oAKhXQA0i9IRoW6MYEKAU+ghoqrmKEm4FTJ26mZDyZMttDNqrXzCn
Tl0CBjRVDe8FaX2p5vKOCyZgf1KSLMGMJ/G3KORqOWJl5+oh3Z1FkVyeKEpk5RPA
ks2YYTM0ywjVa1z0cOLN5D88ByyP1Ol7CEgSuEMiAY++YoJf+NpmThRHqLWze2Ba
ZkU0VDtLpR/CBZOFIju3XTUJbfG9Cn+ebREqdcNDoUFqKqrDVISW/ftWFVEh627i
efantK0SWEHvihUCfXM0qBH2p3Q8WOUfx2vrzt6BNVVndtsdY+Fxy+NkEXxUvdK8
4Yxoa78MS1VukwPPgft8eTB4Fw1fJT3KF2FDDHDauQYC+4XE109CUOSMAoWHOxE2
TAQuay8UZS08q23Oo/XnNOV06mEHKbsvJwvHGkXGppy6mLR0F03b8pNZaQ6GtDwZ
s9upqKo8VdN3Ro5ysbgqiFxd7I3/j8HQyX7mJlNADvvR4bIceKkr8lpWm5xmGSRF
AOCj2Db9dLU96wIyowEry4H6Yw24FkoJK64wRAy5QOe1AipntFxTRhQST7MLKx8T
TgGvMkYttkebsrQCAOFzX4PApnIJW8Xsfkp3GSdKEuBXM/HSeX0t5keHBUp9lPfh
r+PU1NlWCPeegtwARCk5TBNA7/31oQ5i+kXSHti8r6h/S7zpHlugZptCxrflWQUb
2mwZqqy5QPJAd2mCbuzZTMgCxEUGctXItzXtdWghtINoq1qvharKaMUtZa/+f95R
SKZ1eIp1JmHzsHuhkj/sL3C9EUyJBOTJo3xe6W3kBDyb2zOG++nsrwAFEEpiEZEl
mzxHyEJvaKY/W/K2ymMchNIdDgIrlJwf3HmJGC+rfL+5cd0ebAUhzjSOGAjL2wXP
AHUsXhizl8+4Qq1rZe6tzNwE5M1nG0Uvd1EpdPCtRm1g7ATxlwyyqzT4a9Zl45Pj
UYF+1ZjvcP75SH/WE7d5rlRA3Rb4z5OeKLWQHu2HLN0YIKG3i4jP6WFaBgr2XtiL
qvy25ZIpyDeMr1NXj8drLDl0gViphXfcw+RpKGp5YPLVAv7zqCGCKwNdWxWsnvws
kU5CzhNnKwgeaN9tOZ2z7pLogTLKxEeDtLBuv5JP2sMI7juAmhRYh31Q4T3f09J2
QgstBjYehm1tmbuRrcUPxxbRbXxwe24W7vUDMrRPuR72lLIapvGbHAmlKFV8kGZA
78fML2LDegd7Xt4EJocxtgcXSgqO+Dnavn1K+IOIQBJZU9wEGhRe9Yv4lexBZ+tv
gITtS2qhxBwVeWtx6dzaEz1d5k60MddSBvXpaCJHawSg/EHcAJLnUP/UvlqWT79F
hl2SYgptVjC3huS9RBoDalN6v6Pi7jwRiXpSsY2UjGVcFYP/S2Li4OdmD8QZ2xAw
6hTJUkU2vzhjLRRo5xZriHtnaaOircM4qbHPwyNfk1umzQqed0zcbkjLqVT9q2hr
CNa5VQWXUB4IXl+8bGZSYIZuMVF3vonuIuG1aX3h7LQOk3J2/UL2LMelCYIXjVd3
8D2rsNDcbxzg5NAPJon4h+qK7vmBSvpVmhSc+1Vy7HFmTXyIgusGdXiADnp7PGc5
8E0PNfsm+fFNO2U+xs58RGv+3UjLgRWHg8fwSD9ZQf71CSYU6JH8AJFHmuz+NO3D
U2yLhZJE1yKbO3sxKbpdobI9ywfhFizqAVd+VENcuVpByEn+GF6GIHKKWvDKXvnd
Os6uV5Qsm6Nw00ZZvobJntJ8AqPHeIhpHthuz3gfNqbpbcHpohan70KgI7AyYC+F
zpvCUz3dptRZUidImCVunYJywwE+Yq7ZwhPSndeT9NglrouGSOGxcNTtD76xbCVb
RnXtYw/xaMlwJDP1c0QESprSg8MGaWTjBKvbLLMJ137kTzVvxY4Cn6bPVIVekduX
OEUFZtSEIKgI+TQC5ovLCiV+hZHzdrSroFhKYQrtQkgqZzdT0CPN8rXd8fvKh62H
FwBNUIcwxRcd4YgKUUoADMZnd2f4xkMc9TCx0yYoS/39fK0oJEd9t00s9uIw7BEB
q3BSiZj4PAKWQKseSrKn/LzMGG8Bn140UMAZ2dSxBQTUnOZD70DeUQq9hPwECyBk
WsKzUoJRlCNgRZRgpP8j/cozeS8CkH9bCWu5TO8j5SXk0di4uSRLAacb6Pm2aKfv
bMnt6inXzh6bTmjWdw4oF+QRYz2Rg1oM24d5ypUsDQw92R6Xw+Soz9hElEY0gSfa
75draSjXg5//GtNi3J6JRrr6IAB9rUMBCJs2QILj2ynSPpmRfO/Cfz8Y/8j3GLhD
0uUgM6FEMZtcmy06YYuVYGjp0cTg4z8GrEeIIJwrcpxBQ/9AdgIQTWPtZJi0AA6+
Cl3FpbqkwqDFyoRqxIWUFHfIVizf6A7RbFX4Tgrh7hhS0PIHb75MXT/qQILVKSFe
wTsLCXmVeatvFGwbxgV39TebOKxLbaeT5QZ03fhm6esQiAMq4eZXs7Fu4tlR4jy2
uAdMoad9ktHj/Hsm08WwfIf2XN6Eti7HFyYu/oz/VX5NAgA462YjVxDEpCzCWnB0
ruYxR/BDjxDb2/y/TPn5axtcKAVWh+urNXCjGiaNK2FMHvY4q76eSnYrSVU2iiQP
uNOdB9fKlR29mU8xlZzb29Jj0hF0eqrQYgM5lgyttEquRTxW25rYAvKlxu9/t//i
10M7SYceSNSKhjt1tqoexRFqv5DbOFhTPOY5E1zu8km7kfZwf2gKEe1HzK3c5Tjm
kw1Xjwpe7J3TJFi72M9GEOoi7192us+oeZ73zvy43B4/PDjhA9+H1e2b3Dq2Gd5C
oIs/IAG5NckUuah0CnBA2YqgVMljzWjHRIYUeI6Pdy3p6hizMlku9rvDyQoJafiX
+ghyFtiauWoKywq5Hq0L/tq/hxpkgGhgkT4m9EoLmsYD6MJND00i+Y5UfiyyowcT
GPfy6F+pWsnDh4xq4dRrDEsR88sqvs+Sy1wPGjnGOP4TRHfHg/t1+zDYRUCaiVrZ
Q+jsPt5OK1NnOvmG8kgKKDEskdNOPc4oJLdq6wOBA1FDS7k6q9tLlhSUdLBNQ8d4
K7nRATtGrr9xbA1J7VGhBFsdNdsI5F9H4BQERJgMbaRvtfo6Ryi2+T4KaPex2dW2
H/rIT+jnd2l+1pynRs5xFQF7xWmFy29ZP7h5ddAFm8UE+IEQAXiX2AETE6Ej9R//
88frT8nRTNJPUdBTJvAGofnk9gT6GzQCsdsdvxrH6F4qk9rSnc4ukRP+usZJ9xN3
CjlgUhJRnfpwgvyKYYieYeuGe93JfBMsi9sswzvHYrgmAiuQF4kren9l7f1/NQOn
skxaA/96noUXT8Ia+NB3hRLJq7kf0h0NQEmzX0ZTKRc7Oui9Jc31u+tBTfL9KZ9d
f4nIxC20qhApCPcr+l/IEPTbAZ1DCpzUzvn3qJmnsqN+7pF5wpzsaBwC3pdj/NAc
sRBGIxEY5MiSSZCYYvRqAfppR6L71c+/mWKIfzdz0g/4u8Sx9C/1ZqIG9XuxhZJn
x9+OIi+sU5fWDPsgfhW+WIS6W8A8fPW0It8fIsXOUBaCgZHOTY8jBt8q6BxVDM2j
GvBIkZ/3V43SnhHilL9/QbNrmd+DBsOA5laHawwDSEgkn56A4GIxh7/c0gxWf8ZK
UOWIOFrDJl8f0q0bZJFZ/ABHvoyUsryMUGZYDVYKvKIvuUSlcURa8taLYS8XOGaN
O5cqwDPbc6GaZqvllsY9ZlMzpxgImJ8xxAJJ1o1JvUIG4tYdCTVVfTrZpuupO0DD
tEexgkh9FfZE17x+n8+iYKT0AgoVxwlEurpsa5iWEkdv7WLKAu1KfO6HjH/toEuh
H4jTeGq9KznWy2k1rm1AfMOI5JtdGc3yYxbe2JVOC6teZLaAcADmLsPD+lovu2pI
d1ITck2XMS8LMyITh98sMfBuXtxX/TPXtD+csrP0Y/eL58JP6tgiqgiq3MobnjR1
9JCHvtzs/ZrF7VcfBEzPb1UC3Xi5FKUxxpr/pzLOtL5+WhK/FfRQL8MnOg7f0yR9
RmdGB8cHx/lnrtZTfLj8yY8LI17Lwf0RkPGUkDO1G99mrcoI5EAccEfmx9hzNwu4
eiIjnBsMG4HczZlO4q22jPYO8njuHteUkso4Rk8PDA3HJAkaaFVTjSreUbjjrxrc
7l1Nt6utgXUs1NcepLqnMaLh0yZm3h4i/dPTqxPf2tu0SBBb10xMoEERtT9S4V6e
G0lKaMgi23onemyNdxMUDAQouPo9juYe9EwhPRdv+s+TLCI/BoOSmgJeM21KSPns
/u6GHThYkKQoctjRnoiCSTZs0YNZMLpZpfbqeBDFxPfEu4aOcHV4ag9cd3BxI3XA
UITvC0UPDonlnCVu1my0NsfT0RJl6P5223QwsIhC9Mu9I0pr7F3i0YA5Lk1LSyCX
I6CJjG3efIw982iwikdhhIMabWfG/2UL6xuV9DaoAWBisrYkFk4BYUzZUBZiGw+i
4yi6EaOMYwTQspkxGLyprzMd8DQNWYiLrCUsD8wNWzTmYgD7Gqnc4awNdLnBHlJL
QTyH1BCyO6LfYWtOiGvu+ENqsXdAciVcx2k7IOzB2v+oumsBt1Tszrlfyk4zsSTF
Ai51R10NGf+/XD7kEI0uekMS2AIPTpk6NRR1/HsNFyzzAt3pORkmslzeFCzQP7jZ
pgoQc9ncyvb9QqeqMhZFaBeKOdV0j/VIY9qraPendWdDV5N4labZwuopdpPRC+eR
fbBTimTmHDNd1P0iPJagHseteRQpTjOeCxbx847/blUFxP0OViQs30NPwrR9jCuH
4pyGVDiwzEe4fITORcS9JutqtuPVU+RvTPTgd8Vwue/x18ZHu1UR4HwkLvcihLRk
6LQe0VNgMMe3cldwqDGRrIt29sj7PBOsiqIYKody9zJoaQtkQkFMNO7iNlzm6Rm1
Px3tHaUlBlz69nw2ip9xZG0hMH/Pkc8HbEig4qFyiblLuG8ZWxhv1Iqhwg3476X+
0o/5NZ0T7Y70U9Nea6k7KOzgLf5JV2PbyShSyqj0jYU1c+eLTlamylg6HuTu/6u+
t8RFML0xn9/Mbnx6JYo63aC1rgEQPOqAisLw3FRwV+Z9UB+VfHi4AiIplY/Cr4ft
hk0jLISKEI4pP2A2PltKR+2MgWtx3xyPLLaDKsr/9/5ZJaz2cON+Ig49xn35gQTe
0W60dKkUxsWtbRbvhODdbdulmvdrBao9oYyHmml9BgP2OFSHsG7VkVHL5j+TeKBM
19W8RndvDQOZT94OqhicxgiRGr8ooEhCPmy97SLjebdfj+xgpI72yHJF/dOBx8f+
PXaNavO38VC7k97NTk8zahMtuCl3TCGXmhFb9HyGRuKp8gKeCYn4LmIZhKCfWKGA
zcoePcvvparqBbJ+sF9NzmvwxWC6wiZTcf0QMTMDZMyuH6BSwDqCSMA/Lx2QZDT3
28YueQ3FPUjQOMEQ2fjE0P7VRXBbPvYcBcNcAarw+0pyVCxXReI5naAK0v9+CKTz
R09+3AcAprkkdmmN/2GRtNIjgB/mF78XDXjrUK8aEBrrji4syiytRPXUHBW//OVh
C+1hoxqhX3G9HD9/SNad4emJLV3pWjqtGlYI4kreKIMMEvH0CnafU/RxcfEVAUnT
Glk+dmZ7Hzqw+mhiByON9ZUGc2FNBSC86tEwSG/ykDwDpr0iFEApRJLN6nGO+q0T
Tq/J9UN9JZlr0wg5JgvVpkve27d1M/u1NqFbzFEArngJzkanlNAMQMYFgRFLFlbK
YockynevsZncEK/Pk84qx+tfvia7XB6GpeI3EZucm2Wk4RW1Q7DTP08kRSMwnzTn
7FWIEoIlp/r1ny0AGLG4lq1W/L+4bkKqC173w2S2iDi4No1Rljo1MXoVVfiJradn
1Mpodd+u/zlfDfxUSC74FR8RQUCEvYLAiOEgyDaE0B6/0YK07qo3nLJvTvntfCTp
hyc+oqAcfvSp8hmm1UhW0pcAylVfgv+75Jur52iSUSWVf35nsio24x19qzA8017/
x8ZWPYciExsGXWlWyzg2JWyXmyEb5LOULADPA5gJW3vKtZg+sROMj1qwLY+IoXxM
bRhLrXsDkVkx649eh9Gepp9dEkdhHsvFOMjFCZIsT7ZOq3d/wi5yRBkQHgbSJVK/
tBEjkIUS91ka/uB7dBmzC7VHePtMifioN91AqXHjuemv4c2RM4xVZd6ErXIXxO/a
ZRSGmIqP4tXBFOlRuSmAOrAohOrTW1e1Z+wC2CJ9DjDx41r4MfXAqajRmrlJoV1U
PkfHkWOTfR4CLtKv2wtGknQmvSchkv3rkLRPNfFs0Xe2LWQJd+mAtmhUBuh0PXVv
+5Hqn81mducSnzlwJtSG+ChFWAJO+24zSRlsxgjSS/8J44RjlkbfrOyKBVCXLvPA
Utc/pdHTgGLolRP6EL/xzU5AYHw+risc73xjpy+iJVPIT5CKh5kMBRTJc97WcGx2
iEpOmwe5ln7PFuiFZO3y+F0vfNwUq0sClH2SOiMFj8STtSWDl69OxrE5Q/m0Yrxr
hkcZWmv6qJYEsj2jzW+m3G0VbEF8t0f3jQDC0T/jjxM658l2woorrw6LuFxPH9es
ykO5iv3Ye/6P3u17+Oo+qcJI7wSA9ExQIFYjgicfwTAF8MM399UMj71TWr6lNj0l
x1g9CI5ldr21vkI4zzDL3FgLM5NTHpE+Fxth29V/67XqBUSrvSAJq43YlRK8lLqc
YVCzE371xKvkHT60Hd2WGzkkWLPniwuSNuawnmlyqMOQZdyRKU8Ivw4vAkIJtb2m
y4jwm8H2NBNw68LAX0+rTW/3njPIGoTHI+nKcBN8DvXqSK3FNYUKlI9zJcKJcsTg
wHAMNVEMYIpjsGxQj3xH1Cb7xunX5bFWvEUmcu478A2PZHazzI7uOLfbHvu2m18O
tZ/S45+hw6cxk5HxXQ+bvXczwp99UgjCP88eWA0JdQu4vDGLmH0Qec0z/B+lEcuV
w8Pi6tl5p9n81HfSJonPFY0t1DzvMskNZRoB/u9toA+N3TgZFpsu6GmUu15JyaXV
7jU2TjedjTGs+fdOknEbDKPsYXWvSkDOvJElTlFpcD10An8ZH4DiWy63AOg/vGJj
upSFzNP8esNBOYnUa7eqzgMqJ9rEiuQ2UCt7S7DGrNa4J07jRbT5vaXVnD+X9Uk3
dZrqH3j0scd47MFr+NO9PLitNLrRm2sTqZBunNeUHuyycUA8bu63f7cB5lEmwjdj
HK/KBZVG6l+87BqBvP1FdirmRxPvofx28I+gNX20L1mHqfyIlDLPad5UJirtGabX
9Zqwayfw/ac8/reNIHaYbg9lwYbDDTid2n5ekNcsZaW9UgxgrSG72zHxIGfm1QSZ
rcCTz2QsbZClgMvsn3lUCOeptIROL6gG9nEyep1T9LH8Yjo38FtzeirzesFlk6qv
OXQ+vdlCSVOMNXEC8SHUghPMVce7CYD2GL/JEB2ft+PfI/0dwLTEsrLSPFdj9iQE
wkFiCEHnnI2fdQ3UpKJoNoYFepeqXpdVmSyfPs0NR+Sqy40ec2wUhArfgkFYrk6H
7+DQ42xwRq7db/Q35Y65JENkT0HGHob0dRa+PzTVgemm9hbQSnb8AWHCmtQ5/kxR
3wQGWHdzQGJUc3jkvrbM6N8K6J3zfSFr5xZ4bgSd++fVas3mJCVr+s5oBnP2CuqL
reRA2QVOX1xVMdcoVO5hcQMUXvNkRyJ1r+5mrN9veAea8hgPEVbAi88XorEM+isS
Qjlvt0jeh/UfjC2r8r8pKhxYQGjrLlwWW2shmOWpDPeaUCgnHTb5HD/MqGu5OKZd
hgXpLj68NDIo0OFr70JWQshTRnnPykxJcG8biYbMaD7pxzMhg6q297dV5ztKrpGL
ZLPPSM4FF9axaNjB0y8umYTjycLObo70UV476wagw5LDbtqFYjJfGmXgz0CDdGOP
BgY1DLZv36YC+Y3PBBY5BLRXaGNw4gopE4G9/4CcNAzgYFDRT+r6nD+1t8cLkp3r
D5xQxjHkBb1yuE8FL+Q1Z/rRempWD8aK6Jt4wqLTW/8YJKutbyuE/UsDjiLSbVFB
M+d0n8CuIydRYGKgPlnEH408kME9p6frRYP0X5GuTjfKet+Y+vTKfc5KaDWnnxnH
iJOTi05kD8RWIAcL/vd2DFyQhysympHTzKCOiXQtO6jH8OqW3X7J2uYUT8O3DGJW
bDFzZkV9IyYVqWxQiIZ3luPqRgru4aB0H2IntYqUK1qJLk4/a+0sTOOf2kjzetsx
WXh3D9mHkwd2iV4yKdDpSEg39uWwTw+UtaTFvuYjWDQjHR+bHk5APeIiiubbDSub
qniP0pCyox1VL6RuiG/OkdrCLl0sDv47Kv3oEzzzaxr4K6qYyNRkooSYkmz+676L
hEHFUAKXWgi4SjOJaWsR4z0Wax+7hXZT5B8p3f/BnuYL2cMbbGPookGhkNPfEPz3
YvANkRp3hK4KSbu/CoUTgHGiy/VyfNXJGziI/NOGHWcgQS3C2aZskfU0MiMX9z8p
kctYRdyRY/+k+lkcnxS0w12PvqUyxkoPJfGbrHe5FJHjItbXNQfz8Y2GBpFrQlT1
pLlcMMiyWwEq4Nei6yHQIcnfSE5MD+3cjcRu+d8yOAN+JkcurcMESQIPNkOJ6ElP
pVUSuXTzvMswFyaZikGFUuJdEXptKfliDNUGsQ6acfuBEvhcOm1u20e955btpVur
razAvO138hDEdXjspx+vSXub+m0iB7Nwlp9b73p3BtifIiQWe51eeEaDpYcPnMwc
2EU8KR/v1Zr6WWAVYeFDjY4ZBqtSZxg5mEt0uzu4HKWtCTxyvEXTZewmNN9sEJ/L
0sBKNE10Ydx12VwgnB7ATLDfoJD5X30N0baQ6AN7tz4qjkL8w6I2WMBsXAJALSUI
GfRqhqC9D02RbBwFHeKMgldJqBE9+1Jz/gxJdHIqgb/H5D3LwIGUf0Fz3e6UlCov
a+69j6yTcRlwgMfCLhkDUZyNbngzQ8/Oy97YpKR89kVpGJL++dHVfdodCQx2SUnz
k4BqI7zkGXFlfBuJndLJtWvG8vQkh02wIE7eWINjjoGp7n+9CmEz8918SCRgWsw7
R9s4Bm5sAFIF8i2MzKY6EhQpDSv7g0z/t5/7uU3IiZ6Dr1iW83bQr+jnUy4+bN+g
95OLtfT7U8m6TQf9+szbDFxolMfHqJszEdoSzsS+oz3MH3c57VPU+k6k7Adu8fNJ
Nl7yjfKdrZlNf7MuHjWQp9K3uVkXLprhIB3gMI6A9ixNLz4azFHU8zqD5lD5U4M8
xBMP4vG0FttQSSSpugxuCuVnX6MgbN/IeqU1y0T5Y+DVYOxz6lz0O02HeINi32pC
SW+a61amg+1ZRIWxHIRYCwidj4A/lY4xBsc5QXe/RAFbK5Xh8BIwk0lNtJEDRVs+
l7m0uAuxuAbB6Tweu2ZsD2VdobBMwzOQkBBOX/SVvnPYuZ32x2mIr+SYe2t0uul+
DSmzd12WxByckgpBkxzFrzjD2/NvxBrL5SDsdjMSq3woTlrhVCVRd6B5eSs6ug+T
1VsWWfktVLxtTPkvl2fTZ6PJ24WLJkp8p7m66lUIwGy1cAbb6NYPxd4ue3sh1lEl
oC5vdl2Wk4nOHMUIOdKWK9maZBdMk5xCvzJTWxdgZMEQEY0Mygnww0wGSOJUOscO
PUAjVNHudobnsNoKsLNanWfh7cAQEwx7ovJdfI5HeELb8Eu9zjylX1P5pzm2H0h0
f6YsLJmKicnw5zvMFzxOaW9f4RYgYItNl52XvnuVFYP3uBGNU7aQQ2Wb9PxSh4fS
2rrdaO6mA8st85mYufSbmuFV+kupdIguWl+cvjJ4NOrGkE87apA8Q6r1HYShv51h
YSCnOwkHvmBxfb2ohFHsWNmcXHiSj21bti/0IAZ1dqK06ZhYSiVTgh/7GvmFWA2q
wbzY4MKeRlOmb4ZthwoTqqYDl9pEB0Xnwsp66Kq9Odv//0KiIp+foH8MtjPADVvE
lirwiCWXR1no+Qbpl1eXm5jWqDTiUZzTSx3aCkAbSqCkIHoxS6kJTNsgt9P4cq+G
lOG/+JTR+qalmzZn9E7sNE+ZfvFM7eGLKgef2c9gMIjtNH1ixJ2lhI+cCdj4aEja
80kANtAwKExE7p/rv/Z0c0rFabysyd5aKHO+fRkywpEnVVQWnj9nuA2ysnz+iFNN
ToMvFKEetGMvG2zdAZH9oD47OmOwo5kNFDnB0v8zpDm6eMMRWWX6gS9yN+P7wyAy
s735olLlJzVcN6jL1LCWvl9Qm1jOKC7T25elf/4hkTSp3QwVFJ4CB2pDsLN0pSnz
C/2RPPDjNHRPmjFp0Mtn5j07Ba0biQGT5Zv5znK0Qah1F7uKiqppc31GITmUH8V2
by6kCghnmKRdvCplxcmVJKrzdRz3jiBKyDNAjZQpayHtbWbuLxzuXN0wPIGyRnAR
ABIWa21r1RcWqq/0WmbiMZUHRGLf1Ja/1dy4XoJTA59w08q+CVbEKRvXYklShSCw
4ZvxL1iTQc6oKd+u+BotaXLXgtBzSnJDspMsZuVJ2gmdfXowcl5mXHk9aDL0GaeO
tbn/nc+EmQvuHp5k3cdTrG5nV2KtEtb4x5XvjdC2gy4vP0dEWQS82Gj/7mxnUf/u
ZpNxd/yRCDubbBkG5cxdfzOveLzGuY0pAjl5TW09Ysko8QEQPHJxojruLdDKenN8
x8Ho3aC/h8bBgK+00JT7MSEde1pdRyqKSLyGUJqa0x64AXqjrDx/XzPrnuQsvi8m
bTLYrdTJSrDDbIeERsmCd2YVveLeqptK0liUngS3wND8pUSWMB947SOvnilZKnzo
lQOll6+lASLkenj3juCc7499wwXCYm8no71t/JqXSFz6MlcbkrwmwNT2kZGXHBce
4uinM0NiPtXBufZKVLUoKwbi3Y47LP3/bgHVesnDHjGJDBR5B7+IXdfNidx9JUH5
Uvb++K4PorYK4lHVnPiCT4fxeT+J8r7/veNK6qdjQ7kym7LaibmvQ/cN7mmC7GF7
bdmzU+/amMDWPhov+kpgIVQ6EIl2vDmz5Bw2jRqTvIvkXNH/YtMjsvXeMAbBKyaK
gO0O1ld1N4tKHAmygbIGIrWZlYOne0Bh/BO6OK1kOmwQ/16BVqC+zykErX/89Z7G
F8TZ5Ntu6zuTixK0t6SyZfQdP58DGLxuhlKQtRCjNSSSEgaXmlgLp3ugs6u+qDIx
t/7OwzC9H9isUadoXTuRI7kx66RjjdUqCqlTwW4cYhEXNEn/5ypm+hageXhwnofW
ZehA3Sc8XF5f1PXNx2VsyEqJzMPOccKpiKd9HXZpw3KYw4v5Efu7KV1AjdDpp78d
mZ4U8qMXW2aoQOGwMjDV10ai4wJ4U8P9A55kbCf1peeMsHyJ1DBTP5uK2/lu8PIS
pyC3E/vQYLuCy2bcMUSxV+TugrP1lBy7CSkJuG9DMPAeBDpoRne2EEhkgAYW/T7l
SgWBcmgg/p7k0wu9hHhkmctJYoqsaYrd4iH4lhLuFvH0SJ95bZlfYxEduRyqqE7d
wAfyrb994Ns2qK4HHBk+CjZYdhZAbNe0dAWITaKBRZRbE6a9sLdltaHPxXkwFR7I
ijqC/hGrHI3V41H6QmjplBvMo4knjX3zT3QDjsDjl4wabAss0iO/Cghd7T7q4Ki1
2yvfI6hGObJ88MvlbxRPeelYZvXAPs5eFbdH58/vXBfEQ9hOgzf6j/ArHew/jy0e
2zFUPNMWaAt0tJ6AEuye8jAKfh7mJsCxEemDFzICG5RwIqxys3ZIryGRmztNK0nZ
oZm4eIjCPqYhXZ/tS2NZIVEiZq2TV+4UGU8PButZT8vnss+sVZiFXY8DnoNh5Fcp
X9Zl6H/2niTZmWODzOHgWFB8FlZcg9gcn9JJd0EN9J/582zL1cjBHVYjsnCoDM43
pM1axU+rzQIkmkidzUQInL3PIPY4cy7d4qF7hm550trQwpwyk/2rMnQKm4jJJIrx
2+OrZbXx/oQRRRuciq2d+Vccylh27SpVVuUOBpVH737I34p0/vxVv527bF2iYmw8
x20tMgGI/sE50z0uznZ0FvcyQOI31HiTzIFdFsvrCMUOjVBH8TdP872wfsFDXgjm
S4/JByYEBLIFJ3ah9syOFXyT/crAFDg/5zuSSz24ex4cyDpV3Kpwubh+jrpHKaQB
Rm4yycszo9Wpk/gKIEk4QyMRmf3ckUzu7PMMNGAyiHKL1SMOaXlTuLcPuXFsV+AM
z5g02vkvB1mNHAeJ140ZsFf9w/HOY8SZMHgnV9gDumwdiwiYZcj0fjOGYQ2X8E6L
svnxbtZ32F5a7SjP5OJ9FbhdCsfVf6T1GBc+zAM45ubk2mJSDSFJLMIm/OEQaSzH
oDakGvojwzMXjmPBMFamIjq1ZRWQRzuqMrhpdC0ouksfQUu1I0r3ACNPcRNNOlvs
M3+IcX5esY4+b5bFcC+qdPQeSoFLTO0H25gUtL/OdcDBytDXHZVC8uRxK5fDgrUw
hgIWrFww20qOSxC+2sIiz2a/lTo4GPPj5268mz1v19bXLWKhLd8K/agxmJV+pR4b
kzj1ParyoxHClA7krqouSE0WNdg5IoHDGkLBq/Z3k9bzIT4QgHKaJ6c81/FPbCw2
+DSvbj+3TewTrVBrIfRtZ6FA343gSVdh6rY0u3+zqgR4zceIwdWW8nyzktz0ieV1
xn8ifedVhqKDJ/Q/TeVmAMC+LgdaYIlds2jQUr1iokI7cZZqc8hniI9pBM++8hfm
nbrLl8DgURGuL1pZ0nFeo+Guv3mZVRQtNV3OGVqDXzCzHKpTCyC7zkyarJcjyRaK
Z6CrX+JNTZZ7cFmV+Z1KqrbzF3a9BU/lwfEYAUBZ3qRenR+QwXaBAgMctw4SgsRn
rWOj7Ra1IViT6vnB6gt4/d+llKsP7xGch6wNrbAQNoG6revYKrMKoAU3jt7nODze
h5jEmIf5TsMnVOTzHnOGLue6eleIoIwCplZrL/DQ0s1SDWo5ztW5zGX8nDCaDJ59
0Lmbr92VuAY0bksdloIehItBbf00AAMBOvrS9KrntRf78uuPJGuFxdqgIsSBXyH4
JXLxNQEGZ3AoS2yt6YQlvu8Yi/5V0dj7KiyBbDuDPUBO/xQWY4YWQMOnYplaJqDF
frGHZV3GcicCk6je9B3TGeoWGhG6LCWxJRyUVeQaL6WpHUtVjxM5X7Nlg97NL2+U
SDz2oVzDTc7rObVI+mBtBulDlLg3ili9uHvp0vjuv8/ri7tzT+pklAGJ6L9zjE5l
nj0X3qnT9E4DoUr9W7kAnwjijy+IL7EdZ3MWTSmGRtuX5u5EQU+s2HuUjlfBTMQd
y1mQIMhANoNlO99poE8BHpr6yw2B+/Dkk3r+pLLoIMUlCd71Y5IKCxU15b+wzZUQ
bUt3TTjA+gYHrOdCeP0d+I6HkHrrWcFvJECXNw8BAvwfhTlkAv84x1Ql7oR+N9zg
d0ZvKeOrIYjiH7U77HsY6Zb3CsZRtCmTE+LXYqQRTa7l1gktFFNrFFR7piiYWvpj
bKSbr3koK/xFWUzlgJGcjdzuhwdjzhYE/bcd1W4mgYeVE8cC1SqIQHlh1MJj5fQM
5B+AFNHOAVpjGx4sK2addq4yixEOf9kCm9zXsAHhWLQ8/BFtAw9+z41VftcGHI7u
aQD51dsq7lPfOrRh/riSw48ddXmYegZMkRLTcpCRKqw0CJoln/oCTMgAkYylMxCd
e0SaSFr27rGqfuYXSiDcupadCj6YVuYpBoD+qVLYMdQ=
`protect END_PROTECTED
