`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGg5q+/183WRg2U5Wv4X7IhI89Zgkf/Vm9woZQdLWco62rBtXy47kymXqiPj1uL5
ipbYqEym0qEgBm+oWCrZS+/ImgPvmq3kQv5A5gAi6J9N/o509+RLJJ7KT7pc3pVR
1ktSERqvs9c2f1725EqpaiU4aW4epnkWyyQ+GIozvIsr1egwx7a4OV8mVD7cDLae
pceGQqgEp4Gq15N8TnrnO0EzqnmWI7yndW29D+rYh3FIYatB6t+5PHOwAWCt8tsc
GHLsMorUT9U47wKuoMPcsV5XZF8NuvGgdl9eGe7gQ0IK0pdV1sAig9U/Fw18RNrX
NfEBCp7pqH2mLYjDu/HnEhWAN1err2eqHKSGoqyWhfNxvg91RdzRXXbptt9vAXZX
zg7fh6mAkQRIF/C5yc+CMQ==
`protect END_PROTECTED
