`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLXDCAdU6dHoXHmSgQwhENaTLkJwQ3NkeM4+OZ3dyzlS+T+HH/8/RJ/pzqaLa+RS
PfsoVs70Ln8UD0k8mdnW0Z2EdLrvul9yX9q27gmgs33AsFf2pZq9ITpFCMq9WAWd
JVjO8+gjHAU+1DlBEf+BP5AN62bAzwwDqD5gkSrT1A55OmT8BkgJKrNrY4KEusaZ
ecz/ro1zpBVLMi5cOiI+89PY2odOMrLU86pT9/kiWsTU5leWxgxJ+ePO6DspU9rR
EhMAfc5vk0z8iSQFOOA6q4/MWpBqChW9M87GQVOIHzprji0mdFI6ehAB6pXzu0y2
DGWlTxp/WxaIbX0Zr/ONMZQgJeeMOqULWacyNN6ACBwekzJ2L5mV6lFA0q0fDSzp
Mb1af2w5mYmzG+QmRDby0nYQgBUsSdAYRP33nVpa2o5grMoTLvW4oY8bqXMxl0aZ
`protect END_PROTECTED
