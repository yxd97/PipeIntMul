`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jYmROBqSORgPQhZ8VP77zVmL5sG433H5MD5jzOsvFBXlsQ637/I8Zt0sGsDklaD6
GOG+JOvWctCLGDX1Y+GmzEDK9xFDB3xfEAZSoTppsB0TSF3hjRniQGaeeARZC8ZP
6v6bFGH/V9G9zyMgDtxffMKb5oug1lYDi/ivlwpy/Ko3GibBcZS6TD5q/GtloqP4
EQM2nEjieY7R4WZF1EGAEDqtJR3OtGY4PYYXqzdXdcPDzA2ffv1mydrxFsFo2IO/
IaerwHjSsJbOySlRiXhyF1SdgyGAN2Q1g8WMIKli0zJXIAEMijKebZPme6eUr7mJ
1sG1UX5VczvJ+niLtTeTSJhiSWkkC0cQ8XHp0Ii1TqCJNMkQ2QLZ5Rs5S2CKX59x
CTfs3tJelm9saF2zQepM+lK+V6AadCp/7+hfKQq5FtA8Xks3iPstzBiTwaItS9FZ
CR5bpZ2C+qxPNDTNsREWC5yrHDoz3MIbfQe8TG31bMZ0IQkmCsf2axjJPTHff3iH
r5JuDc6TUBeyVjHQ+9bxgLHXLo2utvGEhgcPbG15E1PmH0fb5JH4mxmYwI3GR1hz
oecluWNzFM/uFbP+zK6j4oL4HtpCY13/ZqDH/8ylew0osPk+Lhxi9o9diK8LrZXP
rLCELqio0FV4qq8zgOD+52T7bHTiwvt6sl8tJ9YjFSw=
`protect END_PROTECTED
