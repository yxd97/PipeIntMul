`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xiLxtrQSGgRQAJ6ooYRhrbFLr3PZ2I4QdynezN4kc9FJBbPVotipGwPp0lDuKiW
3F0JOdzbhELCkeBk3hiDXOm4zSkVg9NVp5BXJsaH1N2ih213ZOEXy3spIAi6ut7P
vfwtc+74uEdSKOczUwVWxB0M9yTRN2/wRN0WYUFzspcIcObS658Q3OTKoG3HFCv8
w5RzvjWi527V7JbuQf9fbNYg8Kv+FRfoVoIXSru4KnYyhKqYJeJUBIHOITkDXiTr
W6iY3fjZP/nTXKOYqu2/lbRIuOgLTrBYIHwob/EGbkKZkzuSRDip1isa1xdxwYSd
J/rADX/4h8tEGLbAgOXUfnaqu/FCKCc5KK5R+ARVRsKyox9pNdJrIaIc2In7HHUH
Mc0uB1BGu11Dwq/dYxr6cFCBoq7EEMM3htazPgbORcpwo5n/KJzVtOp15CzYzO1o
i8geUF8NEiNEDJ9ZrMCphKtFC8yjyT/IO4SL5dT1pNomi/pXSyt80qYZzq4Nd/Ll
Uodi8LgfN4nR720m7+6yF3wA+TqegMFLhHEsnVq3gaMbgrQxM+y/N5qofQRGAfME
jFfSSG60PboifWa8tuVHyRY4/KBuICqE5bmvl86x5I1birM8dkMWP52+PaXysLFy
uAoG18RjKEvrutzlo3iM5AULoy0dTI1Jr6D0TzH5ChojjE+UP4oWDoNsK3TvtAwe
/fd3cpjz4OvbcwipBIRVEyFnmMltzpwSDtlcwqvjvok=
`protect END_PROTECTED
