`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HlAR+BzSmGrY7BgSx9jDKEqTlfO7uPTbEvvmvKqinkfZwTl92mEHNR3Qz2KZK4n
U/xBLtF/KfH1gYOvSsE7KLLS8cYP0WTs4K2W3Czjap5DqRco4KHNXMAQIZ8eMYiz
0jkgdNEV+S3q6kNdPOH94ZE/rKKs4SnHaVdr/sVS813p4ZH61RsSc3iUG5Cadvdr
+j+ETmWEnmcH8CBzC7nflwvaFkNFM6RRsix7p8KO6YElnb6jB/M0QXdVTJINNNdk
44KeRqUizFyjoY2Nt8MZFzQ3Q0l+L0FLus1qV3J0d8a4HU3UmzPo1Z0bPHJdVylY
57FbHYF6QInGNtuDWzRcMkR7r/ttVHiB7WlLP2zLu7kiRtWZPPE+E4NEJvUNrOm1
DOlXPwdgal/vYyxjg+O5WzfeU7MEaihUwhcW2ThF0sDH8cWOQJu3xO3iI522YyXF
PMEDBe1wHuRYakQTEyPGIFFges07yGa23hEvYAdSgUofNHZuL7EsuTEua5s4y19z
mOFiH3G/vaRnAUvbqzRAmzH++SVm26oBaCI0G4mTuraT8LWXPeBHXaPt488SnFcU
xqZ7beCVRJv47aYI0m2ere5Vv+NaBEXIrFNRAR9gP+qp/RQntUFwOoJ2b0a2f3uT
QPNqClvDJmKI0AnMCljTcmA5kzn7E9X8ZRPgddYwmELqasO7/OgMD28PqV58xY12
YF2/lZhRq5W2CKkDBaHTcbvnpuHfo6CaG1XWC1ib2mh2Av+HBhPyW1waG+qduUpQ
KusSqsXwmJ3dajfuJ95IIw5qBBvqjTxcLVCIHsmmEcg17FrSAGJrkFi9d3joGGfw
mzWAz/FA2B1EUNCbc9LYSQ9rKGUghkb92bj68v+l5zG5wkUw2W/z/hmpresmUxRJ
klb4+pFAo+r41itA7sYqOGQvIOayW4cg8GZ6r8gR6ObUnHeCvHdKCZuBTbMiTMLv
pJe24xP3lNDQ6hMup77weKSGVEriR2w01Q9PAMlQcoX2qYqugT3iKVMtyYTEO7c0
B/WpGUOiIBPBkuUAoxEHWXY2h0q3FeZXRii/XQlDcdmxQQXV81phqI16kiN9o+ZF
kAZksDbzrF41OHxFf6B90F75XNubpPgtDMlgmWceAQ79/aQmZ5hzouxMqeWTy5na
Ize9Ith4KwjzjcCNW1t2Wb5db/eobXkWLePD5xeVtKGyh2Ru7TrX9lRgcqIa/u0q
HLbXFIK3UhqVATXSHwpEnY40zacbXrz5TfBWyEIBkW4wFBHBMOlxLLmGJg7R5l3l
F10zWerG8yQATBZg+7Jd3gjxa/R16NZuSTwBhqV8UWiO2NTgHr8jqkE7oCGDluSy
dR0JuTBXexyLTzVEKaSRWiSyyBiOoEGCAN/LeuqJ+xcrUmbWt1jsuhVGRVo5gfQI
joyDpU0UVWMPnnsCSNgYsji9KfnP9UCO9lJyDmHiwdVAqpmO0j3Awp1IOK5nlURY
YsJuBCXVdPUr/7DwnW5sxWFAO2yNVd/TcKUrE8Wbb2TAuoAD45wR9qWTwnT6r9CS
+6C3q5rfFAkAPHbpeCgDgN70pAOnUJWEGVpaM9DhyAt+VjPOE9aS/A9cmMudPwb5
08qtHIeYoHJpU1YyxZV/9eL71BlVpji055YKn2bGhdnYKHW5RavNhKG2C5HYhsn/
Prh/6iWfA4MBbOGl6bAie53bHg+JGx5zz8ZlN3GcbksQrM2TgJ4CvpOk3buSLSRs
u23+l0gs89OaKSfGCMSQi/rVnrib3ZiUmBCOCyHUcv73NIUOmGOFF/sDonfEpeGd
pDg6BK4vNyb2zmIo/xwSfCN9DEJ+Efda2KD8lEhB0gxZ3bSHCe8Tk0vGxXVAnu6D
YBhAGHd/yNvHrCy8Stgncz00XntoSdvnEWVQL5nNPQ46UE4zyohfAenr99PbD7/R
8pWbCkXrtlxsKVmwiQBA+5KUwzpid2gpvdiF5+8g1jcm/6wt7zcaryu9GPPkdMwS
Vf2p5EdhIHE1WTzoxEb07CGTB+AAiwXX58UYdROSNNs21/oSAhhe4AhwE/+NRpmd
zTEhfDvYsSgGASJb1uDpTAsC+utniowPUvOkgDijIkuUr3Hizs4thdMwPSkLcoXz
oqas+UX0Z/OjUHFSGdRcDAZNkHN0kN4JhUmtvNkgKEL/3zVnwzvWRhQMW7nKIws6
Gy6lHEG9xcaZYsv4sII/POeKIcsIYSM9LG+vveA7rlgjuFIQZjF8lZSJH5vbNuyi
45ja8muR15MTiFsdP8/qf6bYwFKAJxRfvjrfd6SihYgFglHd4GaezLPseQlWI3p8
4m97K2vewvnwhqcV34dLv0SGLZUjY0LphdSkiHaNL3pYDnbMuUh1w0fbcLYfAPWs
PmY0HhaZmE0IahSqiZC1FQSZAqc7AfansJKALY2Ahh13LQLAn1pX8zT79OSEtjio
p48TItURBX/5Lb0o1rxZaUWjf6qy6JrFbyBRMMvPakLW4gToFyKYN/iLYIcprPVa
u7H6eKrK/d7hdcQzv0QEpA==
`protect END_PROTECTED
