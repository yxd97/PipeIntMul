`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HiW+Mp/tlfpBwTYPOuGDrU758sLD+/zjehbbfSnZYCBXcJZpn9iSjxlA+uWWrR4N
f2x9pJScqHdqTUgfaFvpjRAnKs3lcUP9LINFosXfeHDMlY+9STi4w8o0EQuxhJHK
JVN/lltiGQyPbSfCMRjcqW/FO/D36BWkccyvcK3DWCyYwIbgU7kgY7IHQlaIe3VO
Sjtwph/ARQurE/rtFNsQ2gVP6ap7KYkQd4/6lDnF1dfyoOR7jyNl26N9DNFB4AT9
1oX6tHKlVO/w83tdmZYXrvPfmF9Kj9uQ4qGA/sHeT2KGdG8Q0i34aR+T1U8gDUrI
B84tf3vg3RJxP9sFn2RPg5xg9qtuzhI/h2EYmKiee+78bl23heiQw0+o9xvdw0nW
c35hHkvBeow9mevIGfHKpqbie1/dzWvBuuhoD/gr9KaUZYPZbL+qe89vlzc/G/sC
kqa04KDkpeUSRGQo8QqQRH33hyJlhm0twTahTeOelLo/5ANP68Svlr9tdGtJs3ZZ
IUjvoPf/YvWXPEpHMrFa3kXwR3b4tqbKCvztDWRrF3py2gzOHYsVwesL7LEP1m+2
bFYyDFjS9MVPAlFXsI2xMdeCJo2GpsWn8fz5O7WDBuftLX6dRzlKS7hWCLzr4XTN
zT1eKPtUZjPKjrxnMxL+1dP9kKi7LCAQt6isr7F4IzV9dOPB3idQFanYITcbzsJ7
iGtNz+qqMnK55i6rz8cOWJ8DqxDmJLsfNzRXflCqptVET0I/1W4XW7JfsE4P931V
GKNkPwHblc/61FoZHrKu6h3aNbzZSZ1oZSsgoDyEGWZPtPoY4H9aHIqO6/p2I7Ma
WT9Lpq8rNuxwPSb35ffsjREYgjBjXsYs+6gvqiLG2gHxrdo+U3ZgSYWZplzobjl8
DeKie5Cm6OphHatbQPPtZR0ZMX9Yl0XIy78OTRZPJDq6XxKyd+kD2402C5+egnSU
7IQhDcPqIWlGJqOLgZEUo/2qfv1r5r+iWjzQVHRKxIFtXtUuCSDcYVdDEfMG297W
22wYvTLPhxkZUyE6I9oLDVJM/UAhhJtbjjHltJxIJ82DK5dAcI2lYIqIlOUP1x4a
Armr7DOkPoMqv2pOjmC/SqkqgYWP4SsjKzduErGK7xABS3tAQS2/2NdEj2Gi3q4f
eOraeqaBVeLddJQfj8fkFbg8GwIhXAht1l4gZEhECFskyqtPo+eBYPZc8Ak7rMr7
69ZjE92UUnaHgnQfrmAokhsu+dOydUNIQsocy00X0mc6hTt9FPYxyuhztXE15YxB
q03sB1n4/HjkRYC/N4/ptnY+2TaYDMyue3XVxXrBevsD8e4VfGftjr6uA8sQnYaM
RhluqooRk5RiDEQthOkw4LocyJ+86CO1/t82iNWeWc9TgARocYhZukW8OC7Lif8w
aeC0OaYBbzwZrdDenI3zwVAaRIqAHl9xwZnFutL12EU6FwnHYX1Y6qkvycrBynub
6yyN8Iuy8ji0KQhlFxtHW+qaeHVTpab2aALdK2Uzl7orp3SoRDOmE9j3zpuNs42p
+gXMfgCbCPdEZ0Fx6a1ze0HVuZaEAizGcKs/vo0imb24T1nPeQECHiZOiDiM31rb
KBmnIXw4V4GIrlDmEYpU+YG4RFI7UULbZmfjoEK4jaG55g1DC7t93a41z+U56r58
LfmjowjxWBIDhtz4KEdR0TEtahj8F/6ku5VWrRg+9d/2ZvzBAJ0pdOdyGWzWXvS1
5LkgkTpkS1eUb+xeN7/Ss/tzKr9JMhxi//JRAa9/qbLpCCK812NLr7NdrsoGtptA
+lRr83siJAHIfnGvt6GgLwg4P+nbHEKsErn/7Gk6f4Y+kAcJLzJfry+sovB8R9eT
wYwIQDDxtLIT65QTCkL8R6iti+ZgFNK0JpVOebR4aRoRErIjkU+7Rkb3K+jAMH4j
C+n2Iow5/1tsS06NR0jttGfqsymP3fspHJEI8orAl5i4CPSMjhEAPa4GHQamqnqJ
382BPKUU9yi+OYBmQNECceGytEMgUIpP5rpaFvonqX951/FywRPXUj63XR3CNuCk
mqaumIfXZIfmzsHgy9gpOirjd5zx6tVHd4Our1rMOGe6upbfG0a1vygZDXFxmYPe
JibSnPe1XE7X0tSWbvLPfGPLT8bVfQKMVj0Sp1Qk3j5uZtz3VHJS4bMEBiaTmkGO
sXEaT/m+GiMx6NUsOmUB6lyvyioPcTd2u+NRKPfnJeVDqhBk8c1MApyHfYEgQAfH
O9YDOAwHXs4SZUcFSxgrae962wRh4rONZPUphIPf7faF8GDyD6apkc51xmMacB2E
mKOjujiNfIuaeD69776+xtzU46kBtVmMTEX6zdWQW+yqJp7s0RZVtN0VWpaOsFab
MS7fphef6LCVzXWClpVL39pISeTlUBXeW3Sl1oI4hDAJcHwoY3ZBC1HT8Er9y2KQ
LOQkTWQp50gUczo6grOKaW2dowkWzB623jMq8D3P1vyKVOifz/s45+8pWRTiqrmx
8CjfqciFoce/r09oTL4rkagSNkB5vR22rnDpU2NOdb6AiG/txG8CbNyHBFXG3hHN
hHnHA8vBUbmXQJQNWOHksnm2tNhk7cm9o19m563cclvYGqmfznqRTSA0k5OKrf+9
9jilhB2biG9+Uk8dm9QUAo2LFZr0y4pBghEBnpNQXYJDDE4C2SY6/0/GLOmgANu6
+nq/AIfxKNIfzSzadIKksdOKtSIQ/k/v0Q7rbtexJjknXZp0QYPqwy+X9ViJUhL6
NrJ7oDy2m0T804pvzRi9QGUXgu8hljfywAuYyNFSO3JSs6I/ZzLCR/3FtTYTgNKm
+dQGfroDkVt6+qg1iumvanaVylSejsZB18rDmA54+zvK5zMZiuXKoeUW8vKyc2qf
SPY0W9nv4u2wX+6P0viRr5enaJ71++Bt6E+RiO0DuaP8hR2ZrrTiyoVJRyeSGeLu
xriKkTi1cz/LNvMtPAIyTQ==
`protect END_PROTECTED
