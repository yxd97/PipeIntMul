`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhB8p9/TdaVKZ+CsbYiGy+rf8dQWzq/2lUUxLNX3XwUWPgDYXia/aAylPXVnrjOH
MYQ7e0wcj6XmAoGBAP1CG3hm++6pn4BYRosW6Mgt8o4w0QRUx01YbjxZck4Hn4nC
RXoVqgKF61Ekteb8N5Nax5id9ErANRzKXbLEI3/XIzrj0kAffZNJqhwHAtt/+Duy
iviigeNkKFZlvKJaKWcdbg==
`protect END_PROTECTED
