`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0fpU9DpEM2H26qrTYVL290BP9dUi+DTLFqkAQ3TAFy8f0teWcW6sI6lhoafjA3Y7
f3tdpHMOvJap1vmOKERL2xTZm/uZBeozbBmldHvA+Fg9Pqrvxyg3e3nEQ8sb9bib
8a/4KvSlHMVFBj/PS1iZXEq69Gni+SBjr/4LFfq/n5WIu2jJ/5ZsLDbi2r6p4CJR
YRYyJGLHHJMZEhD1WzNk6/YaaHTZlCZhyl40fDDME6U0+28Wp4y8XI5ybzh29p1A
Ag1JcOm/084wEYmYnKJ7BsMKNn7m8VvO6LK4/Juw0/MXwf1Kqhm0mMsfsb9XdWb6
FgpxjhXu4wEaeAbu7+DarQ+SpzhOMcrIK+rQz9nOY3sRM8JmqQFHA55oDQCRh+Js
7/gIYJEM2Ii2Yd/UeH/k6a53RtIjuTD+br+42H94ZZ27o5LJgW3+aBjn3BmJdywM
XuITG1veuv6fSOI4E7v2zmD6qliqO6BYkg8BH8bbVmzzjL5yD7zVKjfZNABCKs7b
n4hIFismVnaOl8VX4VXHi5MdWcSrv0raQpbFzzpkQHT5p2KOh54Fo0CwmV1zdex5
`protect END_PROTECTED
