`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QcQwO1t+S9mbvNyaVMsx6fTupbKuCuAyNtA93B6VqhLcCIMmfZspGpjHYLDhlMy
Yw9fh/1GVjHtgPK3AQ7ct731SnyKUhouaAQo/X2cnLwULRg9AGKt/e93/jdu7v/R
Z5QAj9snVDLSSbqJHADSNrP3x//FWG1gamoAuYn8w26uauGCzJDDD3lWhtkNb/eh
HZjJEoGJuFLQw7V88y1+ewo8IYbWkiYzNq2CjxnlggV3VRIYnTsVOe0VPc+0ndD5
ix06oRPggTMEEB9WYIFR+/Fe9oC+KZygdBxQVVO2nsjHYk9iBa4GOH9VqheitpLE
rS7mPlPkWTahn1Bwnubq7R6qeFqy1/WnwmyZsL83mhqhTRp8psI7V/bACUNyVsTZ
aNSaxnX5XkDU/IfNzN4xrOrnkf5qadWuVEYsIrJF1LNA4UWonk9OFkS+fAi3B7jx
VyEyesBkqHzPCqcP/MQJkfeLRKepL9MBjaGh1hbZgojgKStw937uyoEdCtw/aVUL
HRa1u65UxgPZjwbiDP1b4c1z03Ag399ZMZhTpJyBiCSoapqTrSquPY+URG/hXonK
`protect END_PROTECTED
