`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dqa0vcAzbbLRP5g4NHYoNqMv9rPEJOtpCBlWUO3grqMWgkdTdKoCot7C721k8CnE
GIx1faXsLNyMzXWHlPTi+DG79KvQxH0zY+A+7v1OW+skHTUsT3a8ntfVgJ86Nj7/
6WfegoGGqjiJJPuBzI38KRF0XmHTeOGi7Ut0UJIedMHeSWLqxvWO3UOifqIUmO5Z
gd9Si6g2y5JUcfBhRC2v4Nn8PeKBC4qW0LlZM7lqYeVErryLSq2Zph6jJfV6r3Wo
E6BfdM3KAvL1IQFcExj3DOwPo5q+1K5vP5xdUOIXlfhDYKauzTHtyGaMeSgNytl/
2vcAZll0/Cms/oJYIfU59YZDkzKQI+u9qfDH0+eFe2Rw7VKusJb7SfSonCjP27kd
57HmV4C3FFivor0/AKAq11cjQ2m42uatIGAWs9ITmXvqf0sI1GakpObcBJXJnqPC
T/pl+/Wtj+/7vAm6mAiut4XS79YI4UJzK7swmiu6BKbTyYGqoQJ8ixuuOqL8sgT6
9DOXWGI2CAz9rCzMO7xw659Ub+hWtzofeHJ6ONPY164BKnAwWjLkR11Z8doKhS/V
2WvNlZArx62sdmnu8aQLMJ+CAIHc/I95CR1W+Nh2Y3A=
`protect END_PROTECTED
