`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rh+7k51lh4bhxPX9qQ3M9NFDpcnNT6BsKS6ZAjJiesyBbuLQzhSAq05aA04yhTt
yBbtGXkmHMAGwCLen0Sn9+4qRgMNt2j1aKrUuYiAx/1ggOUJvQhYRWxMDxzGiSxM
WtN5GgQrcYg33fAxEFVkvDXnydZdDx4B8+/weEerzTVso03ygoim1MpksuNjZlOQ
InBcF+vTBNyyfwoOz38lQfVR/Q9+xWh+/m8j8siv3R55FzQln0rdTqYPZUdRNJQh
5gxIUPAsOTUxpb1LB6dTwuscKyInytJQBJF+nSo/Be58WSqIQR8+qI3sjaH/vPIv
s2Gb05WGZnRqo3PO3v7iRIDGB5cRL8iTv8UJa/La+YuAmcm2B3/mguGm8wsnQpXq
xewyvvLgxeQaRnfJlbQztTSSSOnTx6J7eza6z2k3tCAd0ONXTiYSP3h7GMRx5T5C
tnt+/jNBVQN33/2enBEQ+wEzFJ/yrViAJTQURfVTKtRCQaGyK4JyjGhmuo6O147v
`protect END_PROTECTED
