`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zp9HQaRsNJqEF0GmPyL0G5QzWN2LjN7tILI3nT2BBBWHPFobT53ZR6uNj8/l4vyg
413U1pImHFHSo63AdIQAn0Ac3/l3IW/jZWHpp80Y8i16bBJF1Fv4ZHbhnhO7BXMP
7tBLt+SbkKScP32+f22LukxlWSg/RfEX5uwx5PKRp4//8Y96Mj6N/EG0/AK+1Py4
1UhINY4nVRq/Vl9m2BOCMub+grJMagFmI2GreR6UwmFA5sqSuOY3zctK8RYDARB/
hPwx9y3YhQ7tSqyddX5zU8vXK637gooBrzA45ys7ZNeo7g4NKZ+4iiCWP60qQ7uV
qdDZy0MO9W5Q9X4d1kT/JvUCSNotVQ5WDbEu6ROHKEkNsMpNxxQjilOvG4PYoddW
xEeT3xv66mMfyDmKxdJAMaHYxy1KOU405Z1d6j7ij/jUhe7QBNjo/7HMDz2E3brq
`protect END_PROTECTED
