`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XspOERF3chRfYFYiEkLL5DhVK3itZJjplc3SJ74WM5w6OREX95iJLGHZ0pnKpl1m
0SugCkbQ9ZZDKQBUcnV2jz6ToonCs/nPnAUj2vWL+ZzqDbUWksEdmDERTu3nQSWh
fHX7Lai1vwuRrGhZGl7LtAHVcJlGomVq2z0n/FkZ2UhR8JXdynC/kk7UI0FeKxjS
KMMX+yebkyjRS8lko8AHxedrBnXRdmjTZGTR2h4g9i5/rdqaVIJg/IIWd3OVgp5Z
GWMlYVQ4UmHq8QOqvaJ9n8lS5dVbjGKWe/sG9ACKglkJetr1wzWYs1fQZ2ll31No
D9iKOArhT6zOX+UEf/Jdvne2I2KMWU8AWuMlpkMUuBo=
`protect END_PROTECTED
