`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SSAsz0fxkrAInp5Ei6QVPCyFSrXmyMjBfG6a23im+75xgq26wr9V4/a5qoj77eoI
k/nGALjc/HqBDN/q3DUJNSiN6STD4HlYaqsY1eDacC4xNhmwrVnPJDiFJAwC0DrE
vFHFhBJW0B7b8WsUkZsLuz9Y00GrdU9A4KnM6KRMGQWdG5cidufSSriKanir4UmV
8rf7WI1eCMR3YlSQg54ZolNYg+xjZjLea2kPI4kxWX4hJ5hVnByFuczPb3qdE7Tq
Kxx49pUc6ogjOUUjBK5Mhqi4NXxL8TT2C8ps7wkAXEaBNi2BMk58s3pWYXSOXFYO
xp1dgUU0NXP/XW5S3q7UN8qwnybedu+bhmV9HpRjLABx4LmDpyfq+kaf9XIuJxVH
hA9PWV7Q1eASuLgfsTeIAla++zP9vx/jvSWvXqxhNbOax+fdynzLakOkxiwjkjs3
iuJhOXWqTWaybIvxapbnFZlimmXcJCMZWWlb0VBYSgT79vonzQwgBu6cpkbHqJk0
ybPXnaar8kd4l+G5DMu+VQ==
`protect END_PROTECTED
