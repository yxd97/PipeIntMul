`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mpjhg1lbi8AWIzAGtVeQJmFXT/aJsNwcwne77U+K8YN9A4QLkN+Vd/tOuU0VC2P/
2bgryMN+dKNecEswqeUkYyn5vaCSU+s5YgLv4NQYMoDfwR59YQXuNGsDb5HIFT+F
OZK5+7XXHCuc1PTsBkXBZYUzg4XarSoeEQGT9c17h+avax3+C9aFkqL6SVvW4uJX
9BTgNGjXRMQHdc+cbMkyl6RU9FuLd2bj4YDNTiy7PfhLy9KYUgmrNST/Yvxp41jv
yQpz9s4vB/GzSo2RN3m542T7NYkz+IV4FHiGRvsDHS2BTCvzxgMbEWiYc+gyHYLX
tkf75SgIpIDdD9lqVwwBL66pIkYEZseHcUMFzt/dhHPUg+ZYTTVfi1rD/GSx6l6Z
YsR8b7QQfCYDZbrDly0KqR87S7yNrzGuIQMPnLfC508Lu4lfXGDqsnIjP95UVcyU
os7LLNdGOKzsXKDyJA+P74m+QRM3SyXIcZx+VRbbPbcYP+uoyrrfkVPw9fn2AloX
`protect END_PROTECTED
