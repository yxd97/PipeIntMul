`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FbNxaTfXt7S31TC9JsCJOF2hnRY3NZKNi+u8HgOd7KcclYDdTzzhy8K6nVwLQg7x
za5NvowcqYwb00zuwdyHhBZoVZzC/GQ/gcFxCCe+QoITmZaaGJ9SrdIL9CLw8GUC
KoHeQfyx1DE4WbarUoPKbAOEg9nUVGqWmn0lSDR6+1PutkHiGgCQgySqGqfL0jT3
dGnTp27Qr1ru3tDHYS/26urnjuvkYHcDYind6FHQ0HzyQA9uIFn/JuqNAGpjhkGN
Vv/agzFpEo1ZCULs2s9mYl1OJGZb5B1Nj364aK36Fn/HJR2kDa3ue23Gwm2RcF24
Ur2rnyd8vNDcuFh6ICPckOQWMj+Lp8wBG7NzQpakcy5vcKseYeGZ21RbZSWGvxzc
`protect END_PROTECTED
