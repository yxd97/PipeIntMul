`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c2MeLfIz7ovLyMhHZfgB/S087ZamzTdOSjXKt/30aLZUaLjEBhMHMLJyShRlF7GQ
jjitVpk085Ec8c8ryO2RtTO+M1THanweX/PJ/xW/Q1UIk3apqewXBIq1upjl2qQK
DFCLJP12tfC0OOPyM1reZKtKFzuFdZeEVwqW6h+6ln6WwEbfE2Xx9YmBy+SZCOqV
5RqJ5w0ZM+65fmCl/NKfn3UyNg2Tket4G7iMMCuOAOqLHCvl0HegjSjFqexm/Ofo
ed0nc/bV6IHzrjVZju+V6CQ9cYmEHLHcAioRriUxJRmgIevXc0kFQJfjod1jGeKf
CTPHucENj2hkXwfHYCNxhv4IXojaS+Ik5uQvkFbdz6dRckqZDKZyCF5MREHkw/Yu
k5dCLEp/YQWytfONjokeAOcBzaOE7JXVyZESdWB72UU=
`protect END_PROTECTED
