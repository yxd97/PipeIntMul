`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rlykur1dZ4HnWhHZDtlWFOerFmiR61J5gHk/UvRwqircDqTDCnrHCEYIYSt2V60T
/NjjRDfAGqS0QUPRM284GLh71dG7LlO7oRf8Q5snggxPVy82XMS7f1nC2UfbnzPI
eZ/4TtEJHOypX3cDBcQgI6K8xaOhhLQzfKdhuSvYmwmOCUUs/0JPcDRjUz+Xpe0K
I6nHrtsyswZI/ThCAcMfLnNDNH/XyNYQeRLiDn64EpcvIzxhHUS0SfA+11Nnjbdk
PNraGxunrSLelz9goGSaXvfSHBcyoLYMp9SFRkEy8BCYXt1k6DSsny1wUJgVjhi1
4EC1lYzydS3N9I1xopOg6VKy9KDv+Qpt7jphDdfdWw847pD6q0Uit5BIPewueCvB
i6lUFUJhJBYMuukoj6ckgCLbIBWfXPi/3M1iTpHIbIE=
`protect END_PROTECTED
