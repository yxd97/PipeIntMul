`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0nqd9xvbqywPHO4PZo1MyA5COdwu9b2oeXvqCB0y7S5BAU7YbUVkflNk7uwUxVD6
gfAbc12j/nB8gl4pL6pBxmOJURnshd6IhmcLwNm7tmRlLS0WlU4O3z6WMSZ/g7Ud
dM1e0uX1xNMyXzu1w8BLttuOor96glXdUVn9d3FBwThAeXjvswkJLqcdL/C11Mbx
+IBs+KozgOMV174ga2BwPc8cJ1Z95uLgdvpMlSj5qqvltgrEE+umwoBq+lo53q1Z
bNrfQy59dorGJs0SXDHf9UqMrvvfYMbp0l4wiB0iMx2tIQVL1C28YaGn9/Kt1Sj3
2xvQDM0SL26Sc4wX1b1OGN+pSC+XnD45O4CcT9I7hoik931Y+m4loaNY8eM0EOCW
tCW0DFW5F7DS+ZGcUMWMVFr4ac4njmX6UeHVEZ8S8crKYCvacU5KzW+CCS4s+lAF
N7ZMKqQ1PhvihURMBrMGx8hK6emgznucZx+zuwrX2ZcgbTb9Ntcx9pdAji6iazdF
GqFYwmc7m/pdjmRYJE3e9IuhMDqvcY44jr+b9q36RbxISgEGFuUUEjJNiOWmxBfZ
U21gh94uyGmUQLJUQG2aeEj5QL2w1xWtM2EMdyS3vZ4kNBpjQeSG23rygzWU3DTZ
ITtKV4lb85l8VEfLfWR94A==
`protect END_PROTECTED
