`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NuBGYTPkq0dYMj+lASMkkYqLZ0DcVwR+CV7XStJsMV2rzn2kFOPsrRLQxhsPRLWs
f1kRaIDRztb/TmdfzbOOCp28sJT1vLLC1PwWi2RhRln9JMSju07ULBm3ZoKOCMuN
JjSpgJxOe6EsdAmy7kSJCmnIu9ciqhE/HoaWjgfx0xBp6BcitAIfoHU0F9u/sJ3q
YKfbmhJMNMq1defmXkvr89cZ4e8C5KGo8UvbP6iaUphls24H+oXiTQrAV6/fHRdY
QRFHG/HFYoGjM1AN3rjI2dRXkznYXyz38INpmXpWnC3Qv1WStXppbptCGXpzhUAB
hy8ZMwv02M3xpMCJtGWO3P8vH+D0gu9PISvh2ylKRoyMx0BafvW/3gZypKPHsggz
VSvs6SrjqhOn3RnjFkBg1q5V2us4JuKhrRDvqOO8oY0JIM69Bod3Ebj9ZIS+Astd
cleieajoZVEzigvnBpzDcAensqfCebjbSpT2uQCLfzuGynWQ7Y7SWck4sT0yc8Ag
oUqECTMWTHzz+0jvEuy1XUcMO6ijVqGJZ1iSfMuZbuGqAykKfFLy76Ff71pmo5ey
p9imD23l7pRRy11+UNe6yDdBb6QeTMN/fqh440IgoM7IjvLOuyPSdoL6hA6i3LgB
Nsy+ZKDs29hQqopYXcujIzpYnjsr4HoRGLTkYPVKkpGTYNiklcz1wLgbc9jd0Cua
`protect END_PROTECTED
