`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lSko7/B9Ppjxgrbw1zCCaTi7vQkfXmkN1lBGpwipfhUAFih1emHWiGgvb7fSY/5
ZlT5HhD8cIsDAgzOy+RQ+SwAfGkOYXFRXB8XB0sCEO3IWePGENAQaTeCaabPlWvL
Qn1y6EQmcCxAH1ihCTqyEB26Lx0kLUAXq39s7D6M8L9DoNrBtwpxYnqShSHyhmx5
sIKslNesbGHFmeREfODvhKImHuuBt9Rt9GTHHxASL8UidToI7aSRDziEVCcsOSP7
k8SkIygWBF5wg0qdySGjAOQnIroECcSq7ArFrLbLiyxIXE2GI5iQpEVA5++VoUcM
f26T1LK1Yks0yikTlv30W5TVu+WnG0r6x6TeVkuArOV08wpKssbRZNcb6im69Yqm
bbm8PNsQzOnzFtFXx+ueuF6KuaW3O5Ui/map58tmTKgQcGUjAf6oIEhboE1H35eg
rp4+s+vSpfdJkcjGATl2Ay6avi7EjlL2ME6URwKPInpIKqVPJexvakenmzFWZaj2
eDX4xY6uVlv+9bQvgR/1uruEGBQUII1mw7Zc9OclL0QMCU0fINHZBOORO2Utw7tY
WwDwRr29jDiX0yDs7OOMklOJ3Ai3qJMLmd7cyGyuELk=
`protect END_PROTECTED
