`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1OmNK+7ebyM/Nqkrg1Ak1mxAnOUIzFOrm3byKhgGCGhJn8ZRB5yQWGyPhDrCDOL
M3htkEdM9d5IypKtgaL2h8QyrnLeF0ECsBA0asJWYZNgAzeDIVk4VmanCfls/Ygy
vshlvYR3nzLszluSPhS5wOPd/voKLKXHEG2LIhPVdX18SmYtpe4AEJBmwgeVhZ3t
0GRAEMZOvvbhjo4ygdYdWEpoCMpdhreahs54lYTA97XunRG24YU3zuWP5+f206Ff
`protect END_PROTECTED
