`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKiLsNOp2t6Gj67PSiXpzGZgS5gm3GtKzoB4FuJzl9E03+DT7Jv81P6V2I0cBjQF
uRwo1erhjAK2Q83nX7qiQhiGdKHANH5O+B+cvhMZcmm36LUK0dniyAn/VxdL/MGf
IoZB4eWfOrliUOns7Nn0vGCs0EXFipcC5GOy1B7X4JdmycLtWnK5heJ0ZWTNGxpE
21Zke36V9Ms0z0+zrMo9FTmyzxR7sYgTKC1aGKiKCGKss+n6Yl6vYZWdLwczy2F/
otm2oLqsEYvZF8P6AY5lWh7J5i3yhNfMzIIYjIDgMXRphyuRIVyjGqrxhZEXvhap
OA+WK5cis8+RfXzdN4LYazVaXvnUkZ9k4dYHK8xqbqlPyxcG5eTOs4I5hi2613vV
knpA4VUt9oRRE1ixkMYXAg==
`protect END_PROTECTED
