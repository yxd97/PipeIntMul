`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZN5bcWHPdarcWfo5bszWCyfNN/tm4893iE7ritRv0JwVCCbHCdEhjKsBAaUEedCK
+Je3MvJ+d6rh0YvKy07zuzZf8SsGXoyXSTHvGBm/yK6kmxqqRqugddvjC5N3sqxB
O7HO3B9zyMDfVAs9cCEThtlyKEuRFQlHrXKiAWdi1BwEQcBnK5riEAOgl3mYtw2h
KTSeKsdL4A/pEhItYGQvVwrhEJlmYE9Q1yKNPtO6FRcJNYCWAgHI4OaD8/UIP8vV
x+X5dXhoBHeM+6koWO9HswatSqQxwOsAzmy469QZTnw6v5YUTQJ4uwCulceOtvfL
+cLSgDxwfVmY6a2aI8mnHZy9MP5dFkq6GR74a6lxloVPjHk/tG9/HgNmzWWqSRyG
ZHEjSzfXfejhXL461kV2MKI+5rfERqyXSzxrBRfY6tvle2JOZctVuWMTxSpzUkxM
RHjR0BHMUZuxuWw3BV7JRMNp56eCHWj7lZKNHaKpzJJqMaUYD5lPgB8VDjYuqnb1
lLohSlnlf6c7LOHKLGzjlH+fnTPEwnJz7Jn4cSqAwFeyxWX/V9wxTOvvg9yUA+Ae
7w908mLilWUrSSKIP7Y//C7Iv2yoc8y5nTRFGqhahxFQHdasgDzsgZJ++4bXA/04
u84eCADx066w6F4WhzNpdXXUcrk/lW7/2LBvXndtMf88dM3zKPWZ9zIkZ4dsrzIu
FhuGJDytCnmtbP4tcL7AL3eyq+PN/z099bkmy/c3hJ0/MbUzKJ6QyRiGDZ6P2pk2
xJB5vgTiAnd4KmKg9y1FbwoTtWGSWBj2yXhcW65gc1TfbXf/NQtPha038mYePLSX
YyLGez4MvGDrm03c2hCP3f3vBviDLbeMbgaXpHO7bDvMFw0PQrmLEqZhWxynggxx
eaRqQ0wVAFw4ufnBpTSIhkQMbhoZa4tXrDRmj/nR1gTYTaV/0DOF4/1GtQnY3oDe
VhxqCJI7//8Fj818WsMmNWJZ1OSQQZ0MVvcDfnxx6rLw3moaCJcrbRLdARQ7NKBK
1iLFUcHtYxnb2VTKGeUaUan1UAhEtXSukkUjzfpbVuDlvWChP/uGIu3MR0wRpr9R
8QWs/O2eCDFmYT212+YM2E8O39z1FkFYDaJBsfbsaJeykTTH8ra/zNrmO73oGpvk
b0k1U0R9/1P8zVbwduOeZpbvs8t4KmjcdyQJAgEnYCUe4PQ7Srgtn+AKHNteQXL8
LqiJQanhoTzF9qRAMtJIzmD9U7kSC+TJuNxquI+c8iqccYuWMfU8SZFf7fguWWv0
1h4+6bHwu1YegSlsFEd6s7R1D+Dvkr/UTWrGhVJ6wSwPQHcgqwRiPWEmEpAmSAnA
pXFWlNNSaklnjlj4DEby8xTtSisgoU4SX/rEhmeB0/DPmC5utLYXxBpMEcIL596C
k46bfX5jUoppEDibMkz5vanHk6mGk90Bh0EmgP1afKaBsWDzZ2mls+uTt/02Z5I6
Cyu/4JQl7HSLhEK+VBRFHooE7Rq4Zz0sfDuoVRAu6OWwo4Ty5yQgwgIwe38oB0UJ
aDUKhUhq5NIlndnTBIdawcCir0zMAlwjpG30d05rz1zqbdwukUvqUBPyhKO1h4Ic
mt/No9Mugn7BZbVLbew5eQ83ZGtaUh3vN8KU/T1+9EYFfm3BjzLKdLLeuPpuI5jO
qvyDyQshLI3iyo34VYZg/Smeh+ZS3h4Z+YAOBPK26/dxYjC0z83yEt8J+UoTlohX
srRaGQ9djC4XLnCJosDurbvYfT0E2gfyHPsQF/ndK6bWY/JGHxDdaLYPK5w+sB86
speHzGnDIkFOt4V0ABopKqs1ALs3ujAHqotC8eTyEzSJ5QKhkef3MJX4LvvI8rkg
MIjUjD9CBA1M1Ue8+UJk7ujUzKELXYtm7z9+3gxpzmi3Q+ont4/uHLZNOKdRmLZj
z5y1TxmoVSWMwNdVRMFQXH0KaT3vDGQ1hOw/yYK+yvxHY6uM9gtceosiwNNNw1t6
04SNRUnh0Uf9tIETzYuWMsNgfgN4z/noesFL4KHpfk9tgyRnq4qMnF6fr2uHdVn9
WSMXDDS8BTjx4utiqGt/RAD74LVSb7mmGO3IdYJRzNa1W5hy05vdTy3FyZMi3+XW
kQvzKLVzlGQNPKRwYtj4VV/T6l9HXW0AZ1krhpSJrDbX152MM4H+xrTTyWGR8ZAA
Q0S0MCLYpHP7TN6ALff+12ucRrUI9+ciEQjBVve4Jg+mVohg34KSylaP6plp25t1
66KTv7xaiLfwZ/lI/DyABYd/LawDDbnWFx+nF9yAWOQeKU5kAHp7OXwTwuT7gDi2
mgHH+DUSH8rfSg+MqnVVhz7NT4+Rmi4qHsey6iQoR3AQwmLt0I2NDnqd4jxyGfyH
uV+5SkRkLyTYpySIkrTscUxyHu/vVQlO+Qe3nL26/iv1Gwp7pcW1/A5L8TRmpusm
/8hu2eEtqXTcjMMz2tRtiBCtMHhx82eR57JU4y0BKcbY91F73SYBCW5+L0HHePeu
qxKuTmuRB0rsOmv821HkJ0KAW4NhfC4R2VFr7Csxp8kvEASfPOl+p+pCkWQliKE6
6V65zCJgGiHIimACbqEH7wQ1SQy5m3nG9V//xDBdJewbd27sOGsCW3Y7DWvpnwmg
iFHN7C16TXRfeuaz3UpM6/0CbMHeFb1EZIpz6Cq840RJnqSpUMeNtJlVc+2HWM3u
wsOJOdrFeW4rxzDbX2RaIavZHqY8EfHgm4QW1cTh8IgdtirlGg1adsPIb2E1GyIV
`protect END_PROTECTED
