`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsR3PYkH68MoLREmQkk0QuZjO74abYwoYDj0TcV9TAlPj4CeXYNYei3iGnntaJre
CqjpCdYX7SncWFjilMbePAIxWtTOQLBBeeM677h9Ml3NLteG0MZeP1xqmUbPz74S
slza6V2tGHDluCvpNBXXqpGVrMhszLJ7R5siGkB08TsszUi0yPI3hsyZeU8w1QPb
Rm+c/7fnMeGq7KOehjwZDe10cIqE6rrfn6Hvw6VnU1rgrNXvhTX+JkW/kMIhwdBo
rsCC86ZxPweKwlFxA4slz0cGmuLaz908mBmy8KwmfPdxIFKOxFcgmXBbjv/QQ6sx
WBy9Q4r0wGeJiHOkXGsPaqux6g8EizdztefhADj7d9BdHe/MmAFT9KYGLPVjaPW9
36YPPuO85axf29e6xfI/PRGcw/TRRVn79ANK5Ry8Oizf8BaaPaz96CJ16vV9Ltlv
ALtAxjNqxaeFPVU8fna4Uw0gde9k5TV5/WZ1gfSi1sp7aa6dPiPb8kh8uY6j7gCE
aKZ5GvL9zskMfi2TjAFZ2zlxp9x+/U+2YcQs3PY7LHf4+MN+iJ3tmJNDuL8tsB/z
yD/HJAbcQc0Ov6QF9JWZ/W9banrNYY+39M1Sv744kgwr1iCKDRDBetRm9lYLKHTw
BTFF8o0DBXKFc9szJzanjBb/+9+GAvdsvu/rBiew0yVwLbEVfcwfDNv8IyZr/uhl
r5pktO9OjEwfu5edM42cHSqVf/tRnTNgc7ze7bMxYkI=
`protect END_PROTECTED
