`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbcKhzETiK/XGPvqcDRLquk2E6imJ3Wz1Ofum8woayqVbmWbcL7+vSiXqweveEUc
30ZeOy04ck+9rJy5f3o8tssn2CfpBrrRHXw3w1b6MHQBHsWkFlxsu7PL2YpsVUzz
E0ZrYOKVVr4cs0kIvBZxXTVAS7BGx15IoP+/r2Z03ZoEKdIdCRunInWlT6EOXxp+
qOatq5Z2GnI3i96/1+zloQDdMipk4Act2sm9+fH+WdtyRFAp/L3fn+sozUV2MyMu
ZktFXi9NHb/VzcI0Fb4GPrVaCpHZMwCfQuHj3YjNbcE2PcUK+NE0rYHA7UsFzqz1
hvEEoAqrDFqR6G09gavixddkZsPK7gWWe8TAEDpoIo4qBd30Y/yqNr+FneV/p1wx
+D8FQKfam/XhPsrFaOIJgcuxfXHo/ADtRgAJ9FCoBUYdLZye/eiJfsRAZS0aXpTj
hgGA0QMtkBsD1PL1Tcoilix7Jn+LFWNU2UHZGE9hFvlFCPcvlCiHrN5q/kZkgatV
qNWteTonCnyE0l/b3JKYYqogLlKF7ONihpTGucIe8rCE8UMuZE12T/e6YzdZ4Zqs
ndI0gEeslAclJKPgz34/FP4b1+2yDu69GffpIluvNz5Nxkob5BGC1aKkXxbweDHI
k5NXWJAhHhn0ewtHEgvC1sUTYXVzgnxOXijzkTZymgXa97A4DfViYWupABal6flR
NyGCq66qsJu1dwV1sSfM3V3vBZewIUuSt6eeE/t2RDqIZXDTGzozm7xFl3Kh60bl
zpVsz3ZQ/gl7CohBf8xeHsv+VOE0adk06qHwpd+woa9Vu0qsIDNfC5WGtMepGKpS
n9dH3o4CWuNjlxj+as9RxEER2cd/CuGos9FHgWmzJkoIR5qfVgbXPbJReG8CAwAM
6RXNjhpJ/kJ6vKyDDlxdQYg5kRtyl5Xg80lBDQqnbZuHoinVVZLJv4VAohB02uzS
YlVs+ZcDoZT6K39hz1PlAnt+J2Gj7cuaPWISs1RD+ONlA7UaFZXOdmliFaYr955N
nw4HWdCMRLmhhuFB7SZReg0roGv2D3Wr5zpr42K13L3UIUSaKZ4MxSXPjmlwdIMh
OSRLTyxA/N2u4JWg1Et2rg==
`protect END_PROTECTED
