`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PFPsiKjGYvlMEEekd6e7ubyXcmW0pHh+QtHsZdmylwlAh+HRo7bij9AP8IS93dsM
sRdqT9ZxiB1way7OLLc6vjsBQd6ZtjX6pXARO+jHssAXRKUfdBDqllPdE4wl4+xj
TAA6g71G7vWsYQflFK6aDFeQXoasIn07oiUX79QS6i/UG6XnBjuJ4qp4AHxGcl8t
I7jGQDzi296HKgpqPVIitVTJ+0kAGrY5WZ0Wt9PwUnLkO4TYxgAOGaldC56Nqk6d
g4hYBoTgDstdggjCM1h8cstNxZ4c4vGXHwKATzBUrYcFca3m/Ml9jNAuCWAncz8i
biigqm45LUgcV8qGnXKia0M4vgNU/zYGtTaNdOgf2VqcobouHBgTdTxi54MRrn1P
Lh+f9HDG/W2qFX7LrvL+plyCOITXeJpQV+7lQQgwjRU=
`protect END_PROTECTED
