`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bFsf49Qg7pK1gkjtACFMaSOncZOEC4UEOnwNaqOMQ2fK3VjVVjX1VcUz5d0QOcoo
//Fi4DmKCDOAVIMKtsoKwQTibmbAACllOtnz8fzb8bfRb8KLErpDEq9LKAfNBkPI
EtNPLSLaBZXvny7DhZuODp2qW8P+jF6yJH12+JcCh5dtq7RXCjRgj4UiZyVUtU1F
ifVtpKMzFlz+HgmjfU00GGQ2Nu9L2Zlsla88FtkvU1rKr2tDV6Tc6u2+DMa5W/8Y
D0KFGwRwGsEa28bPtgB645aygMs5vn75DwxPh0K/el49C2hUdFDFgOwHZjff/H3J
NMcjWu2PHMSYfcU1cWKm+RqHWQjugvqY7Uw1OISB8D6fEnwVS4sNYzkt0K5s2Hrs
5RQwPXnKx830f9S7NXfJow==
`protect END_PROTECTED
