`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P5g9m+crAlmMH1SOLR/7tWyqcxpoohseBwPgd5CyGQ2GHFhPA8qSE6532G/BQA8O
RRbrKzQQ2FdjjC3YSNbxjd0X9gt3S5sfz2bTmzeEjDuh1hGqQSR1L5ldyKjMX2VS
e+Y9umMNKt1I7fWIURBAPYa0/NqNoXhaDuClf//wffvVGY+OCwiq0LoEFoywoyXG
Rvjwh9hQDeh+YiC3jZTSV++hYjLzkq3lxZ378gOllXVGHxgOLksG+aUzxKICXYLm
VY5LmfWxsPJ/1Xp5XBkcQG+/wskYj16uda+OiGydpVOvkine9UFIs50Zvo3rc7my
u+h4wfR4+Gf/ShaxrZa81EAdpXql+7Q0TdM+n2TXuiz4j6hkisweOwRDnbGF2s49
wnlwuju7qcWFzLQYei5cOlqhHycYpvOb9vpCmFsM7HWH6TCne2TtlBZq3X1UYIgv
xNr/GD4JJm49O7lFPlxeAbgxGQbPvrjWDJ2Jb9DKW+2CDLDw5vSz++wzwAn5pr7p
`protect END_PROTECTED
