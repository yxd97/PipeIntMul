`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hBwNQ+Vwv5fFMnQQWWiXNgV4N9uqx4iAjP3qv8RU230D/wXhcerE0xMAE6qYrFOx
hupw4B0Vn2DJn/4azVhfZ3TEm1qGRRktYLXht88EVLTRLhJGIj5aA9Ymc0kkHPPc
yNN/JJhETrxgOdX94ieBQpd5M0d/0/ffvuumDMkhtxs9AjC9U1PlnY5kmtzYA2ao
0pC7LJ19S9kwq1hZopSSvAU+uyObQ2otCntRKQ1OcT5nf58r0DCXecx1q7dw0212
tnSdThY7+KOuQRam9qsf9slPSaDxWsYIsPU7cjcr/sjUj1u0wktSy5N5N0fxIMGO
q1mTk0e+6bCfxKCPJbGhNj5+H6Xtw7ZrsJ/DkGzUHFTFlPCJN9CIfpbO93XNb8kM
oK1a2Tr+CURaNhzQlqEMVJsY5+B5lHTQ8bPPk/tjRryUgrJCRxbSwo1D37Sb1fic
eE2ZYwaCzHp2I4+S+DBL7M+1G0mlTmnQOll4Yfd+qG2uwLsTW3lK4obwBsnv/RWy
vdpxgxiW/+vtdWYQwBKWnp6m8mo2XuJZgA/GaBcYNpXadXr9Qjc25BX+UQkESOQa
g7v+EXJt4Cde5IJqGSELPuXWVHtR4zD5skwcEtQ7d6+Y3UzQvGjQvHn+h1EDwRbp
kkO/7fu5tJ1lV4BO/WwC66wGhbScjMOpvzgscmHaX0+zbfKxoLYnBY699fSe4Za+
7pvdKcGlcIijfrdKi9Sw3kTKPfgE7s0dBT3r+QfjgdIs9higHlQrqx2UUXuq53A8
FtyQOgyA4AwICDYUDPpcMAvwsGWvIkGYHyheCGdbw4aGrYUD8o/yK8YoPBh/p1JX
PNSXCFPhe4HiijDcEFFdmCY4YHPqprfSOIp+zapB3xSpDixISl/37MMLkYjJqo0U
dAZmDx97wY/yQvtOp+VSIeAmAm1pS6EkMpQUSXSE/YKLo4DJUvvkpjML8GIIeQH3
yNGI+7A5hBIttNb6DfsDF2Z80hN+4bxBHYsiRzreDPuA/LOHNlH0OZOStxmFs0du
l37L3DnPjEqSKqyx67Zh0gcYxM58NfB+0sRlg/Mo0ZpnrVraw45bLmksJuOd9DLD
J6WDeNLclKjPVv4ibyvhoKdfrX3Zxt+t4RltH0jS64wEbqy0HgI7rA3dLp2VqgV9
Iw474EfBWy5zl2JYPKiGdhxQrOhaE471C7gUvVYHOFWclBudnxcSlTQXdi+KcmEs
7pHy/XYiOyNyC6XRtiW9qFJVQ8L/AX5jj2JJnnnfyZQkFtUIvrnDA6JxCrblO464
vgy+vREKHszSMFd8ld90rXOlWmBnxXUkRuUmuY/s+sFOvYvmlOtgVvIZa4R/exOX
WQlWHmLqS22a5unohAP4FQePIe5eUsTN8+Oc/co3J1GyGt4244U5ZKDU0rSEdpOd
klaD/u6pQAIP8tqR9LWUJpu2o43H25jHdLWz5ES6TlJAI7AhrMeuhjt2o2BPz9jx
82jFtvWAphsSX5iU55KP8f7+AuMbVBCQJKdr2xzxmfbkFFKHaEckVpIT8xn6YJwI
qhbeZsPqiYdYMKI+ESB81h/jDU1kdOaIqw6sv3vCtfE+OxvI2L0f7ID3ypfC5/47
4KD4mG1w3dasQewo5SjI6T2Pmz6UVDUiJlgmmKBsQ+IXYufQjXnhe+f9tLpcok3L
efD6zYv2C0HX+v2/WtTn1maq1Mi89Ll0dZj+iHp87I3v32Jg8HWDCXw1Yqerj/ts
3ox2Bd5HQlKH8y25yLrMaDLbRjDCIAFbTd56rq40CQnKpih/0u91RTztTLm82lZ/
ysbsK1I103PUIhWfKyz6E2PoO0IecJfdkwrNfAoe008OHMA52d+WSrYOLtbamQyl
EFIyq+zVZPlEe6RFlQxD1xb928wwQUc4v2iKCeJ2mhb/sHTDCxfzavV6NfGruOhU
JkGKSF/8LbXlmOo7x2WSWOxor7tLwm+ZrCO0l7euwur8dS3qD/fJAAaJgnCY2xAa
SO+JJJQyXLkqR6RPgbNLTeGjAYwlkKpJn7xSPHa5oQwlQQKBJISQQAZ+gESh+nuJ
B7Uz1KzAlDhnABe2sy+LcKokLpDz3MaOfkyFUwhDeXZ6p/298RFBomWcq9/6hqQu
Su4RM/cR5nwyhhuV/J6ZZ0mm3IyVV97wTbk4oYLsHGQrVwNot5pdlHpc7lOJnila
X+Qwf/vWd7FgLpIUIiLLK2lo2QUs/eecQkH0q16yNLafJUmk7iuA3W20hCj4Qg7e
CRRKobrFoWeo8iJLmoSU05KviyIcna8TpGDHgB3SbdtE2lOsgAOClHk13alwuemb
AwTLv3F0VC5OYRwv63W3lYmzM5gBwIOTynn3RbyWDiD3HzUE9LU27H0CcgXl5z0V
fAz0FSkQZtyZ+MXhxK+z5HVfbLSXvKcV8ZwqOuNN49yZXY4A6TG3QorN7IdvKd1u
9TTqug9wN8cj2ry5KKMOrGZ5jzGFTeu2a3Gw/MH5Dfhbxz+VgKYtkF1/oKst5AAl
S/27SnLhrrF9qXuAQitse0ezJjX4J/p2UsvWQhkfoIuHtFjdYHLaZf7/2XkHGnqZ
WZGHywBLxMVhSo4BYqegYCpdRzLjib7MWXI4RJ5yKEvWHy7r9T5gFnFFuf9LZO9j
jNt+MA6bxuwg2K7b/k0/R1JQg3diT+hkeolIzZD2Y0T73qbx0Ir0ZnhY8EMAyjbk
ds79E9y7s+iLw2H21aNu7P3G9kvgKwACt6ITZXTGGkalM8lh1NEanLkcTDvvKhW3
8/eZMS9SWIO3HVnGSV0pbfea8Z+5Htnrlbdj0JK3pJfhrj29jOoN00Iimc7DQUDv
9r3XqByKsj3Z7/OXC2e7oX7Xblz9rxOb+M71IL19FfJVBmpHchFGR4179MqzAIdu
PKvj63vzVmDAcFvrvqCl/Okx30EZyJHJFFFWNKeWAXKnEUpuGykfbn1US18fT3E3
2TujomZ1AvsiEx+zHpXBWG0sbOzvVIXYoSpHKRe5noigywCD2UYBHvlInTWwM7F+
ia6deFiEHqHabRbgrEdTo5+FwHUeSaDZsN71XIm5Ct2D1rkjeHVuDHuz/Dl7Zase
kfTIyh6mhf3WeOrgeTo1upkUunEz/pmg0du8l5lzXVySz1iDZ6O2iiBtTmTUjkK7
UyWeGGtFvYtERvQWaykH7TEsEJ+akh0Bk4+mNqCd5htwX2DpJhMcrzmOGuLnHOvz
QRsuYfqtCPprvRws5rfYx3TSaxSVcjl5mDmlEWxij/GdVidjG2r9+t0U0BDL0Z3S
zn/YpdQIzsWS6YlKH/TsAd+uN4tsgyqeIyEHZNqXWof5F3JSoworjl8mEfRo/pf7
C6bXqs4lYzxC9vxpHn9k0vk+hfzZSUBq5RK9jmVfbyQMFewL8H4qdhSkk0rpf1mM
wBYwHHcWgVGu062w9q4e5KWEr2niCc46Ozhfn9wNr1WufZwpbNdFiWNWiw0JUyWl
LO8pzgYYYzL7Yvbd4urlT70HmwIHSFJqsNKzWG2y6BY=
`protect END_PROTECTED
