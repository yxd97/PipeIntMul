`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KNVCkNOi46szswvIMT7XE7dA3rJ8AzoV7sj591UuS1XBBlFJf8rCfJ7kmbrv9nV4
gQFhslsd+G9aTDCRTJ1xbEcZIVMUERaugN+vnxJpwr0dTW0XV6QTfmXPkVE1j2Xh
bwwNWulNKzOE8w46JjraUGEJ42QrHG1oatFNh3mSAU9E/vWFbgW4VOdyW2glVvcd
mzbxmDCcIP3KVUArUsJYc+esQB3ms2PQ6E6Ey0SX4qWJroDeHP2CyzJhDP6fY2zQ
p708cusNWhcqPp1wm33ACtj48E9cw+lj2WRITCdPcfhj1a3szJnMeVhmpR/fAHO7
RIMvJykedWQPpvZb3bXOmz6qnDQQ5knHzReCIVoYf1Af2xTTWLW6t0BH0RIMDU9A
XNZmMzMy4DA0kBinlbw5QopJdHIo5KJlwy9Hu6SuujvZbHhtnhRsZe5NXoCDVfNb
6RtdPqIv6lPx5YxRyCGDdjmsdQ0Emhw+y5GKQkJCtaNne1/DETpmCAHL8dl4ViC3
KCrLiG4eTYt6dDfv+kxEBDvin8ym/lo8qcChWmHL4XoUMKxD9QomRJM/GrWQrQEN
Radi0YHif/VwVH6mwXXA+FBh32jSCiUQoIYItuCEMld4X6hPENqDXaqIdyzY3YSL
+o41c9hQVV+qq/yvdVeodaDhB8JrAa+SPqurUW5kFk8j7yWfrHmrwQRn51sMbZS+
`protect END_PROTECTED
