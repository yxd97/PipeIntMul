`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9CoWcxV2vNy4E27w7DaEBQanns10B4s6duzPYcV5+Xx5tEb7dOCPMOxW0kogwrUL
4WQ36HQ0TRPij6+985PUWWExHBws1lsIoH6f7F9HiVRwJkcedA0RTIBjLpSZrZb+
A3jZ2hHqpKa1jh7Iewq5XLKaXjYMhx7ySerZGpvTyMw05hXNz1SZk4EKrZarCGIU
CwsW3SPerKq2iWCN1l7I3nwudtiT8z0oxxS9TrNDGHV8dy1YQo3zd9SsvCKDk8Ni
EfZkmlP2ChMraDvSYZrNejXYw6Q/fCditsQUoNcVL7VTMKumR5nRSZXQxf+7dHIV
+ovI4n+B1rqASq3PEeNQJHhfwaetndhtISLXo7jO0DBwu/h1ZL+w2aGyfn/SCfxf
UtEHK0FOlXFGDRawX03R4R2rECBVjXI8S2yH2wP2NL0o2LETxDTBV8we/HiaRyyQ
hvI7rryPt/4PHVk/GgsQzRuFLlZK3WQVEMRnFvCaZ6g=
`protect END_PROTECTED
