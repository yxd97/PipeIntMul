`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wL1SMyKQ8cfE03dBiFR8FB+WIa7l4tbss5ceN9zHD67tQFSOHelnto20vn8Z1g22
1fNPSlCaQpT2J3p06Xsg93twoXLq7kRQuni8GSQlCMNv8tCYTYsm8SI1RaE5Y3M2
OZOn9ustCvsDm3Z4rkuXFQiykKfv3URmEeh5KSv0Pd84gL7Y6qsKZ/lT26HzIbO6
4x36RIwQu+kAdqhz5Uz9mJukdZQcmw3RVtu3yM60/7sjLSXdEpLCgm5Rp0HsyMSP
tzflwT5ODpn5fC7UovC30tvJJHsgpfTd+dc26mE5/Z/L9qO4kirxIlKvVDYZNvYk
BCN1xFNJ1+JVYQ+D4fy1SRrg2TH8Qw2fv3pFzMfQL4fHnML+xok5fSIqsCrL3CNc
MOWoLRf+V0pYIvD3HjdSBQ==
`protect END_PROTECTED
