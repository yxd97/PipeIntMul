`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swcyxCMVYL0MZL8KSUFrSIoNUqiQGgy3gcQAtRFGBE090YBAxm438qxAZDKOErEV
gb0k/HQ/e0Tw4Dwi+tRDRFu8EhwWGv5ymKeciu3zLJQU8htZ6S/T3He5dwKi0VUI
QRdEOviCHJSJ/P54HqCLuzX8sUoDZq3vucR1RPPpt2unDrL2M85NkDAIu5jH4mm0
pt0FCrjJkEFirmjBM2xUtBuSorkzXhVtVDZw4XJFA13EWSO9bZCr6soPnO9zxrIU
eY8rmdvLdBsTHKMQuwegwGhGvKdK/vk3i+IUWll3z72sNtvFmqTVRoYyt3JAtMMY
`protect END_PROTECTED
