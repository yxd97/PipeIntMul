`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+qXT196WBTwfJnEyxSsMygAlDpaiRTfnXf4X4K+W9Utu8GMCXqsmelRgjJBnX2Bz
C4aGOqggyh9whxZLi9HoxtJmdHwzl0qyp0/buzt80nXW3VBWDyizr3SuQFwR26Bc
6hJsKLV4FqMNRDt4is92Y72dnWnzAuFcg+ckScWq6fAbVX+Zcdff/8jj6tQcENgC
i9W8GcyhUl2BI8tcr9HgFCo1i8pahtFQ/bYvrqXQ6MWoxWqUtVA6HTUsVISb0Lsl
e3wr3Hyfi+ziMxKQpa+27/q4HuKV4mdp0HYQowtBNPFE8T2SpglDcL7jUEzKY6tC
0SBDuuUwWm/+K9b5woJVeoAJp5VEYTd/bgYthsIG9irqAdOFetztMa9spjVJmx15
hXYHkElzsO1OJKiRJ6LUQN8IRXCJsKrrQG9d9/c0iabQRy0RCV6dsvn9/7UyB1bl
veqnqe4AfnbhpOvPhdDlLMy361fqoSO50WKs11ZgsUzlUTPqnaiPdtuwYdNaO/Gb
ALLlKk0sAdTWxit+2+toRiyWsA8kAS3K72RXwUUf/RjVbBpIukW56T1T011CaRBD
`protect END_PROTECTED
