`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3SkonB5R4w//J361nSqxDTURBlY9jAHcIcTjAY7VSkE69Wqr9oiZTmwCNQYfUxv
bD+bgpzJ1r5K8qIBMyLO73m/3+FH7s+Rioq/4p9Wb2Il74jIaiQEfHRZ3AHqFl3p
hY27miXm8n7qh5e5oU2ge4Nprty9VIu/Nwr4x90E8ksrcATW8MovJVWisU8+kI6F
4RR1fWgSddELZkN3MI3UTpr7omX6ITfRhg6nRO2avBeNQ6g+sh2QssxD75aX3jgC
qGnqiqjDiCQKKFSILDPDWgz+5lfugwc8Hes4Ks9jr3dvqulKYfrctnasBh00WCxe
LZOTs0CI+SffRYx2b3pdnILtZi+iqgJKQuGbZJO/XUW8Te1u1NVXuzHGwNUNrpkP
UzMa9wsv0aFO+8OkM5LgomZuPte78sD2KQZNDVWbCJ8F70cliDNuc1FWzP+aZ24N
iMAet6uxmHQVBytmkV/ukEAv9O76xijhNt3r/u+rsVE=
`protect END_PROTECTED
