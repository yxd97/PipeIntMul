`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gq0wQdcwSMC9H7PxxwSxM3x+9T3wL/iiuJDBz3o9mSHlE7Cm61+qgM/++rkyqB9K
LzaroGjudg9b1+9HVqf3lA5rM2laclHD5kzOUSSnSMgqCHs3oc2M4NR5XWOTCWbB
tF4iJN0LiORARu62KdKCGrspVyEv0Nx4DS0vak3NOok8DV5kiUKfnwbofjlkNXTg
YbEgHxBZ7indDAOEBisWnXE8KTpp0WnlXUY54iVdnPKW675Eoe7GtQM+M9pSAUFe
AwhL36lh/1YOE4ncoQWquuSH9WkOzNaQn8OJxubb5kHV1fB68qZ5Um+H6zmEGSz8
9hSdlxtpPQa46nvqzpp+ZGEs8gJaWUtrdsjUoL3kdNBe0JSIyFD+hcl/pvQAzjSD
Q1VteeT8FMwSBM8kJbW68Rbq010bUTUspR3gZhElA8UMSH5apGai3XcsnpvTIUAg
FFAEPNrtOjufDZo+E1QN6yU9lO2CxHz0BV5MZScIXqqtwuGtW/uFmzmxGxoXmGjk
dnn/TV7377g18E6Btj7+qVgGmnZyqNcPKmUo1own/pgmk+CYO4CAzv3GaUfH7Ftu
/4JMhcoxQFWGAyAATkn6SA==
`protect END_PROTECTED
