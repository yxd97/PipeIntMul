`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jovTZISlAIGBwhp72l3SPrDApGZwX08HS+w5jkQAtQ5mCf5rJEQofRDhg7fz1jMw
YI7b6D5UUEGvgCnRhwwPY0brAV1/EIY6rPQ3+REwOH3gXUhbsAu/O2gr/+heLwuO
ctVVAsLtlSX8On2tjxIN6e4tDvRpMBN1BAWiEzH3W5H7yIMSbbG8cyKpgz1/9nAP
fICLRUgOKEWpFCDoE9w1PlOvAxI6U9EwQrjWRTx2GqMKAD5KGkwZkkDnzWDaoHRa
QIqll2DYw56ufCIGd+jP7EVV8mxOvCbLbO+T+NrP5+8L9q04y9UqNIqPjoBVZG6d
E+qduHRO8dpmU0EiRuTSvzrVNAOJem7qyg2qw3U6hVHaLdlXXagosmklAOfiAKy1
9Z56OS8lKZfHiXe2zdceO7DKaA4JrrsrqBJobO7MrqhIfp3+A3QDMWBsqY/fVC+u
W8ri2HjXJ/NlY1/UHXLa7MGRkqNAYmKY3nQnjZYrmZPOJaXZ3aoiT5Gezhe6NNav
BXpDvRdEP3i0bhWqTWAi40EWqiGeGJiHR6hMKI0N4tIv2nGSR1vxy7/GKlhFk/H8
MdpCb3XFZaL/jigzdaa0bUzLRrJYT/6Qt8RMxNTXYqQwe0W74ZuyZGJEofTx177+
MJEWf0uMHpbZZHbnFjxT+WQXCVd/Tm1XUQEW2dzLl9Prdk1hPSbPNwMdrPTWnGS0
Jn9R8VtQLr5cjk2+cy8MEgZB6HlOdnOtE/f9kV3BEhl+7B5sKCC5yTtZx0xNqReR
`protect END_PROTECTED
