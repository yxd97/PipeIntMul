`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4oLJjwfbW9NQh6IaXMnkFsUh/CaLBdwGqXri8u5krPm5zVad615GPAMA5ADabxay
wwQrWlB1DPtHh5bkwnWLM4xppFvPfSIZMIm4WeSZ6OYgBe53mBy4NKyW/xh2i2QI
eJ15JwQhQz6ygXeA06NSK2F1sukwz1AITRMKiW3/ENYZoT9vzLk+V5mzc0taVTq4
EpArYGi4pdmNWbZlhIi4PLLqKPD1M8cbFomr9CC3SnGHyfX7aSARYVVVRko3spbk
XEHOW0CUksXLdxeFMv1fbywr7P+JKi+ImPD5hZ7vk9uX6Buz6O22sjXI+bqdBB9V
cCQybNXrlWHULR2+eVdYODgXdZdvmiE2bFcDKjZe5xdMo+HVDEyn4qTewgif1tGc
2ZdJ8pBSOsqGr91zNWIKuNyHoh0BZd31LJr4RAEXlIwhXiCNyURfF3bblXNoVHXx
Vjz74gfeS1vWFOSfNNhaYa1vQWkNgHtMs8KbbGrsnX/SRIqSr4GxBgEnzK1QcHOI
Hlpp+vGPdTo5gy/Q3vZ5PIqpaREJBjirOj8OG0/pWPJp5LxMYaq6+0cyaTShZF8S
7IkYx2jb7fiBntm2FhITyQ==
`protect END_PROTECTED
