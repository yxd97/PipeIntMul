`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
okAoEApj38W2xWQ2W3tRYx3kmValNRTJNgVOIqqAAQBnBF1o0HWWXFe2Ax3ud9GA
Ay6azbO++im+KuJPAaRFPk2ZgEqdIoX5KVNwYyi0SatZwFFJIAI95NKWcRiVuhyP
eNhsNAO/JvHLx77+0gWwnAvqnkdVNpD8stTX6wzSQZka1/8sXGRAykpgv5Lu6LUK
eH5Ew0HW18A7DjBsD9+tGCiNpOR/o8arw9fI5JnWf37bSq5/nDTKSKhLFOdfqIkU
oNVPheVh/ZXSFeU8NC9GUWmszT0SzCz5Xka81t7Ax8SqKDU83RYbnraQLdukUA4F
t6TfjKETOeNy+t5Fu5+KwX4rI/PGEHxn4Hq8tLQDTcdDSjDzW9siPuPXaByyehKu
Q4CQWXlXABIfsgATioWs1GPxdkhI0LaTNaa+NqqM9v7HkeCtjQ/5RNZJhQzx8gb/
+OVTskRyE+jk9zV6eNdldGftF/3dp4EE+GDRX8CzmqRLAV7e2jhYeZB7OrcxmFgc
`protect END_PROTECTED
