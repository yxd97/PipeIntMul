`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3q0+nuIC8RVz23KqSwqSDOSNZ54MoNokhaDpE2ndcVgEaVBzmq4NR2B9oecHOZn
2ZPvBsI3FgsWWJJQc/OoWQ6EKFIUJYPPi/1HUj7krHrmrfl05NoJII1HlWl6CYb5
oVF0SSB3g+eMfoO/f8PQx/s1OYOk4VHgWKIb2CQzPueHbVAdquYYRSyaokJVgREY
aeKOsITqmGeb4seUlz/OjFXn4e47gnV14+r263QnY+s+IiqLdcIEHuWmXksAG9C8
atus70z+6Pjv1WLMBOQTucvUysyfk/lvkfpGQMTG8PtB+cUlIiJIpYUYblUqiUvi
KirwQ5hTin10Qd/hOkISVQ==
`protect END_PROTECTED
