`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rei4fN6oyu9Y2/hz/71WhQZxWYGo4WjnjJj9FyWSN7CSxRjHk0b4gsK2PU4/7+v5
KufnFgCZYrb/gwZqlTfFZmwX3fw9bFGRRxZPoPYmC1tPEpfmAyAN0tINy6dLnzk+
HD9O/NqllpRbuG9UTKAq2T+z3VNkYHGUTb7bA35FwO79pQMy+hMhurf+289UoMXY
U8JCujCDKTbpD5KQE4pbaYQjwyTdkgx4Q+N5spWyJaAwAl2OCDJbU0Bnxu+prwTg
AJKW2DFdBeEgH6Y03p2Hq2kLjeNhXrtaU+OxXbnOvMMqlHA8ljBUF+9KVDC7jPqZ
E2NzEcPcwDTRtS6HCUTSIoGSWkmrmn7bIWFCPMbzhl5/uwSAoEoZohQ9kjy9uvCm
DMauAPpsK+oAtnpEwXwX9g==
`protect END_PROTECTED
