`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrt1IY6DrDHJc/Ny73Lsa1rGgcsmunAYQVVIdmKxQZ0IsA4H3qusG4ISyxI0SBES
vNdhIkBs5vRQQ9qJujgwIaw29MajrLOSycrBkl30bbjuPWsHYOaszZ5cyP5TDzab
VoiojJ48q8/KoSUvKjb7RQuddMlDqOPp09hduok9nZLA2g7+wNumFH6OPsOPphSn
knypNQbcClMmNCYAn/Lz2vDivmcG/RkZBFQHDGo82sEhji/Vmka821aNbHngafNm
53Ob14pjYIyoj1f9+wEmNO4Y1lgEtvS+tNeXpnzclNzc4ty56lKI+wywPxMr5IIK
TPkY8VIT8TAyvLuXhI8NLyDfDRCge6vN/JvPA198wVcXRk4uJNw76AcfrD7/x+GE
kUHUGYP00A5K7YATK7JW86+7UJnwM7E/8OgmWn/zM5TM2jF98u3z+Ol0lY4MBSwL
0L7aPk2W94h/qQD+wDZZW4JiU7XhWiuV1yrKqH7lqqPEyymmB5klNTJmyLmdjoO4
uYR8Xullpt4Jz+kpcv/+MlhFdemBge1scc1Etdus39z9GkGob462AKK9KIeoLPPp
hI8RjP+wf7+MTnNzNSS7qY1MFvi2s1IMb3h1WYrSgJ4=
`protect END_PROTECTED
