`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
252gUteWn+okesxDX57ghZWrwWQCBFD5ykhCCQt38E5LI8VsRG5JNl1r/Jmv+4Rb
fuB/QyjKKVy5tpQSxUaWPcznk4/MW3eTkzKWQPSiYA3k5aaF2301F01Lif0ajZ2L
1CQvhI3fxCbiRJJMeaTqpAEfYh8cn5BvNYagXfaoC7gExN3PcnsoZ1WAyLclAKu7
jqZIYeRKvT/SAW4blqwybiQLcsCC3uYEUAjbYL2ZvCQnwF4hebXVMs+5KxSCYT3G
8f346PEtAA0JyHkSIb14xByZfyJUur5ErQX3R+KrcZpMIUsQsfREgcj7E7oTZqUt
JpY1BDRfpbeDDhXR1kYX6lTwKhCvHhHy3myhZ3iQTNVPOYkAXi7PR71zBBaP1GTM
9ZjnNAHvkRcTdVKj/Y593IjhsJ0hi8nHBwQEgSpSa4G+ACL5KKhzWex6awhsPUcK
lTlGIG4VjFLj4wYP6UY65FqVx9s979c0nFFvpRNcbTU=
`protect END_PROTECTED
