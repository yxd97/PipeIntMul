`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sVmJ8sKu4K1/agYCC9tclu8bn7/NpCaHhqWCAlcmQJ2uDq7YNRWqXQLgZ5w5WoEB
MwPshAGbRt22xUzcfhKKQrFLXpzYtbSkh5ipiW075Zzq5JSi3jGOuW8HQYEIgOPz
Z1IDfD8SudCb4tKBZOQgUdNKU6hzAYB/RF+IaqqiKqZBpYIsUdT0Esdyin+tvQk7
rTeYlmuPogIFtLtdtbwjFaF/gE6fBjV0HxSYDlRQ1NA7HU+qXbdBp1HSYO0Rt1iw
9yu4m4jOjOqs9o2wcZFh3iknufl3slVjNcQqpcZHWHaysWGQ3utPhChNwEYDBEUx
ZOYvwWHlvrhfgy6z/8rnT9iswC/2UtcXMKb8LPG1qRV9crxZWk0f5yK+4SjA1Odi
5d+BZxA0ar4g8dMaZEetZSRh4jfbm7r6MGN6q5SIKpowRlo+huPfOxO2uZFhJVHx
OcP/JF0dbLVjuFiswMMXCjBzNTzAHD7A1szPs2+N/cwwDhSq9y7HvnreGsMYdh5q
ZwT5jwdixDbZk7FeB/uTcYI0R0BNRoXnHWmHojf3v3tMvMENeIuKxolPdCKTVwmz
kArqMyrMaQoHhImqXOU7QRIWT7is4406vZF+Tr4EdUwAMtvE/rGwKBKdyEKdiMpm
TYGyBJNFGirTjca+EwQkDvXMXc48Nfuk4MIKHOQpbb6QNxaHRoN8PtVJ6mgtWhIx
QChxGEOvz+QGrDLix8LP0bRYe+yGXATa9OfLUvTUyKxUeCgQlmDOzbkB6YGZ0SJo
1pemZr3vR5i6iHGKToPO47VpwzA+yzlFPFfVdrX0F8EFbGrln7dJSlexNlt40JUM
u6+VoBnZeg+RPmZC6aNZigD5IBJePZVf8EzyUTrkNGScdBjFNa/Z5epEBy1j9qjD
xp2NdXzSEwcxa5rdoyRPzfOFbtU9x6Y6l/n9rL/H6pPS9YEuJkQVN+WtnIXbeEo+
EvvPnqKgp2k1VvNg84uLa2f9vXqsG4ywIrnSnAECUzR9kyQdG7WRNChXBzxHZose
DwdxxWL8mhysNfM7Sq616eGcpcu0PhlVPyQFnvCPgTDAbNE6dHv53d44d/17FDDL
hiLdLdAecqN+Zs6aDHHCJI95+0axV3PZxLwT1WmqEXw1d00/UfqeK45N/dLU4/30
JaLSGHQk8LXMjvXtVklUbzJK2p4XflhG7flEqyKywBDf2Vbj52+x3uNibTO/Sw1f
EjrRdZbVj+3/tDge7lD9KFESTCSkST0492Ex10reRUJmF14rcHmy+evof1oOQ3X8
WGc5+ovLxal1XbWSFTYa+B8GUOrDu0ZgqqiV6tDoCjQ=
`protect END_PROTECTED
