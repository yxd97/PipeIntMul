`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OpVEDb1AwknA1qarIH8qtp75JfKizc43+1zx5TVln4ZK6c/MJLeBKEB+xTaB4WEd
Shu1IRVq7I4raFFkuhw86OSfGRNX7HrVYF5PbuAjjURRtOaMZUTC3OG9UdZMVH7p
ug5FG0W+Q5tvim2ZF4v/VGL902WD7WegyEvjoZ4gY/zf8s6zCvogUzlZjbkYAMVb
BGEsee867rHO1QF2jP7Ljof4qIlBOsUr6w2rcLp5hFNHu0W8vcS3J8oV1/MTMoa6
wedf2ZuRWo1xAkSpM08wgoSrEAx6aD4bDkvkTjIDKndE7+mxWgaqhIxSDGxZYIyc
zbotslzB11QcF8ogP1mHpJl93l8nzYsKmtfPsNUtasWKlDuU3ahQuE1IhglLhk61
l7p42Z0ZTyNtrPNoao4AR4Ik/jDsxETGgxpGMluMvpFckwNxozKhijQnuGzuP/gp
ja3SeBuUL9CxqsvoW9sEK9mUGf4mNYSm6Fo0F+l+Mm76iQStIH/ZzlbLBhI8+H/p
OY1h9REkOW2Kl9eEpOLs6sD5htosDTnRr3Tf1l7xOBU/SYIXNS6xjns+sqlIiSGq
PfjDy4AbOkkj+kNi2NGDe+IYEMpNweUwY/xEciL5fpcj2f2w4Vm9TkXswbkA6I2R
Yopgpq8CZA/nxIjrR4Pb8IH8f6lIeLquYVSWAava6VSr07v3PYkryZpuVISoQl07
r9PpGUufGI7oU1g863bCtvtSBCWP6egDTS6iLIZ0HkmynAKLu8wlciPK3yK667nc
UZwLK8Y3EhMU33jKkNiD4F8tGX89t5fpS85HqI96ysTrBtPTZ1zm55KCzEptgI7s
7WgzVkUywClEDbx6e4LepZ6CYkaKTDEillveEGdH55jgRI62G5v9kvqg8djpT+Lf
b283+M8RtbC2WVYLpHzF3B6wArp6ZKCbadftBoXOW79y7+AI5o/zSuhaAWPfFaC2
FVR2CCydn0KUYfNWzzyiconSmOvU0nTeiUNlCntKeUqYc/itYdBKoBiPfDsK+sTw
AVyNT7TquX6X2Wm3+r5VQzjWtFcYfGLG5Vydy+1AxWeLoTHeH5pV3XisaB19Pp2u
+CtXBZ70XalXTWWfDCYxS4KhZuCqoEW1NYQlTgS1qa+/Def00FIa6P+bFPKqSnyf
39j+UbGrucWBMBcZ4SrqQhvRiRRZ/LIqRcJcV4GCJjjsDWoLaDMPr/K2+tBBFyOO
TFkldsLCErlLfzsmgKAdXVAg22ewy+n24VznCFMZM9d2/fp0XSe28jzMjGDftzEC
QH1WhIle+GpgH7yuo2hOPuAUSoKLJMJ0a33nAIWvjDr138BHHn/S7gK6N2tQf7+2
gun1mxW8D/gFIAyeKKstK+lgaT3qais80ChqzpNSREil592M7AUI1bocjiMVSzn/
i6eKVEXV7jzlhJ2LUf6AMVjMxmvhzlz8eR+oeLVtYwsqrO2+K5RhI/XHXq2wWqYJ
Db4e/EnjsCnEomRM03r8uk32Da2MHbsE+Ob5N07+dkXzABAOoHHEtw3WmMGLk8Uu
5R7NAKy6rlkeUL1XNcrmahIVMzX2hEPDu7/eoeGyBrfW5/L/WKM256x/Gg7FnGo/
htQj5j0oreciBCoRVhFXxWosLhlnuEW1GVa8pRv7h9RoBpINNYtuL+47uUTdLs3r
xiXiGYIEZslriUzxPFeK044K9T4Siyc32PnikzfVTbBerES1bFmAC6mE5qk/vtjg
APJ7yl6nrZvTTV4/q2YBIh2gDF9lUtif2OZqHceJvjmE2RN21EQqXlySmjlY4HZN
hkQKRw8v3RNvrjXSZ2u3sjndsXrjInYRhw7zEQVJmqqxAAZpF8aQdwmln8t8xjsM
p7d1cSk6uvye1pbBfXGzYSAUTm4+NzAvGe8PcWgM72i9u54CmrQV17VQG40gApXC
QsPxanwK98n0ygNmSjjFBam5Omv2Lh8+qE3OvttwpMkSQ6IjH27kFgOQ/RM67XSm
+YHFcGsbFaCc1C0UM/zHFXacfTXNt7Z3XsipvmZUGNshXkYckBvHVjZn3OHBzo0B
FV2akKGlBV3UFVP7X2v3oJf6R6HeV5juqar6VbYykjh02t/0A06KzI8vgqn6v1e2
7F5kLv2lXwX3cS/BGa99uHdwTwYHlta1+nxsv8lWNTHxLQJSYrcleJajIac34PUj
67e04qoZKrAc6afzZM29W1jecMkQXGCzNUkcyGPhjrBr379rMviZxiQk7AEB7OyN
V9jg0xCwNnXQS9l0XBjiPVuJkGZXYAAQBOTtkR+SUu9nuQ2AY2/L1i/AZH5jhcDb
aBUWOZu4VFjL0xgIYLknMPs8B2cke+tJwtQmBkV9HwY+0MPPjHda4nbcblvIcsQP
tQKvpgBjk4x4Na+LfB7w4RCu8y1dV4OURsZJZym+VwIK3SzQm77vjlH4LgqdbA92
vXmcL/eHt3HGQpLKZQo5foZrgGTO/pOZ+kufMJpyIbRJhuSITDuVm+BC5lHR/1HX
YkdNhgzSkzLocVyJpyP/O6q9nEWvgJpW1JnszCATInB7wRq1wHgBzmO/zs+Ssn5E
v9VnfaGYX/ZVo2QhgkjTVx7Tr+vVXlGGW1ukLQqZjHc=
`protect END_PROTECTED
