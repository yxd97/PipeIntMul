`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWqQIFCdoNgrVK7XAiAl928j1Hqd+cCLgyyUmZ+IWutGjF/HHeuPpKPvi6PLEHlA
HOhAwg2tbtPX33ULStUZfDNVbq1ttbv1Gt2ux6VDP5RfQtXEokBRTbJyh6zOlG0K
Bt0PHfvBrfcCnUo0H0vFeoSLMFOtixFOVmYZUpxNn2fu67urU3xXndgawICjmaek
VUSxIOLheNaMX1OkFYELraAFoxo4JIdYAC7S0c844rRmG/RQpIjS1wFtY+5FUYNX
C8rU2eBjzM3o85/uHpzSpdGoV/dGwhws1W4QjKwQqLwz6HTxcbeZ52HftrfgZWUv
fh/RIPwkqS3Sq+YZtB1Oyw==
`protect END_PROTECTED
