`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fx+xViUk21JyCpgubS593TJ8sGcyO3Dvy1U2pZgHXy1Uwtq/Z06kF4hbW3D9BhHI
mIpjMjErKSumi+Cng8ThPWZaxHORM89auZci3QyepfAeE5MbeJkOwZrHn2E0ZZSI
ua0l5UIEySKxdiOW1P5s7mfM13q/+5es58/MQYR0N/dns7MEePrDpfACizzohAML
fPgIpAb1ldlln4uO0GKiSCj8g533o3OMrHn/OEVzE9ryHJAYgzKkpODCnNVBMNdM
F+PxgAIGMH9VabqNzHsQkzAdJTyXBGU75cdHKIL7dypHdnvE9MKBhDvNI1X/hYZT
Vs/cayM3h2ztThNgyTUwcf7qSHRtgwiv8v7g4x01G7g6209G+n7lYVmD05Xq9tQY
Xk9iG/zCLCYoiLTBm0EzRl8m905YA4K7wKRUds8InNFSbicsTANE0jVXZOQ276Oz
Pw9X9yP2fMD+P1sXLJvovY5rRrYCGXD4Zm5nXM83Y0/yeZHEg6KiZMHPXGwmIQ1Z
aBOqTXcSK2nyo9v+Azh/aSSeEMN/6q3KAQfbw+JwIs1EWOSgRvglccbKf9kvVaOH
ywAJOI6lh54dRuySFzW7qE2brNzV9cE1APl4vr4FGjiFcwvi9nsj6wLj2AK+l+SM
tNLbzfRd0A8dRCvOprcUmqmXcpmetGOVy/cIdkrq/rq64iwwTd3TLgyBoDynCcH2
HN0RC6HKgq8rst/7xjjIZT+bExvYJyFvGpHEU84cE1ZJ/KOOdrix2cqI3q/gF3AT
JP1/j8OyLsw48uDgyosvQY/xn1oyZlM5rSxjKQLM8EemufH4Mer3UEvW6/PrkkMy
C4gWykYKuwaVGE1j83dh0AzVYCw32IDAud+wg61rIqSqDJw0dT45V1ZGmfNRxEyI
1kgUHEKwN/gc/HQFmDpD6zjeWwp3bwvDJPEOhw7Y1aT3hIlPv7yN1Wj9ohqD9mrj
kRlxd1uf0YXtjcCZc6aXaB87ZG7ZRm8acTWgqbjvwKXWW5B0PP24kBwXS2Mim2bI
2yn+nRHkJjIYViUL10FLPVNKaZn1w/NZtrecpTYp7/Bdrovz6+jSrktTfwvREgsZ
ZsEzhfFX2aQAdSLZV387fq7+vRJYvuID74LjqLq1Ks3O3nrahlSscrST/Sdxl0yR
jYa2/IW6tscEvb8UTVwqiTyWchsneiILawHTyaTi/yL1lSmYE678tngIa4o+D748
Bhtg7Y0IQ1JpduPBTgiHTwE+Zo1YknSxJKiqBC/Igp+xKbAQpaYOx/VM2MwaqKl+
eo8Gd0wK9w1BWE1NovpYJlkpRlxnb1k9i9M8abFVp1sc55B94oslLjhEmjVeP+xb
NZ5ja9TbmCm7pYnACY2y5oePBQF5OXTj/RMTlZZjuFfMUQs5nMZ3rwyaoKCx91cD
0HyFFJYrPVv1nhMWc2hBIByZfCaxW1kasgi4s2FvfYsL/kI+uWGg7POrOMMNxM/F
6cvvLmclM9it+ps3G+MG3Bd5N/5lrRz1R8VZ6uDmQsYMxlNjcYkGh4Gmfd8xnLa1
MF2BJ6uIiE6iQx2YbWV0JMrepqExCXhdu2sJ85gN0fGmV9NTnHFzOxvqiKGVukm+
w+safBotpc777V8fkO/IdIkEu+nd+duXjnZAjZ8qUsOTP95ZzhAn+nddEwfJyKpO
y7xJ/RrIueBRSQy8+wIwkoy2lTjBYvGrhfGcZDKRlh4rSuzopEejXQugocvu1o8q
4apimqlcF+xhzPVxWQGaZj/DOCasr1FZ2P/bKVqEnawtoRNsecLiFLyBSwoIqGWw
zyehvzE0ithwtwJ/eKXw+faI57HV9yimvKZSRoMfmtWnv4Y7PzGDFdE8U3qP5Py4
d/lD9IlMmbLW6Rz1sZqmKLUKV5bNYrO7VAd3U4X/IZ87Qaa6BW7QAx6RaSaeJT2w
+Mzgr8V6Yjg1g4PhvtTK/yEIORNDwxIJfleaxuaMDrwcY5+8H0QJFTgmDMilsn67
YL99beUCPCD/PLyrVCk8vXVWEKQ2+Drvr7n6VjqOQyDwLTwhDUz2LA9L7GETA1uM
fM7nsewAMZc6dNt/UMdfvKPEgawDmCfq6pmPax0CTnzOt0nq3DrEzv/NA5kZAg3E
T5n0eevQDPZEHHxDXRccQU22PAU/I+p7hdeG7QPDPa+HXfv52q4gFEp+j7UMsx27
Mtw5+m2t64ekX2Hbp+GyAzubqMJE5TN4Hu6mGlReRKTNe1Zy0zBhA8X+V/8M8XTF
O3bpNB/LGYtD8fwvjCKinsAdCPyyWSvMQNv9TizPgg4CSmZyj/OlgpMS8WlrMKgC
zxth45ihzykFtPVJwi5/6kn6tUV7no1q3kv4fJ3xioWqQbxerdyXFfL06Yb6ZGkv
fuHGQ3zr1HZS2vDtHEsmjX5wbEaxDnvK4yj9ZwnJtHy/UavwgNXd4PClw24gmIKD
Jd8pilGEZvBqzLbEDDYcc6Gug9fw8T1Q6rfu9cBxp0ib9+f9fg6WjiAKy7t1I7RD
OMdLI1S+uIERTW/KZr/wdMY7XjozXyb9WkT1+EXD4KuGwxtQgKeDyU5qb7VyaRow
M0MxftTjQJQmTdlhW/q6TJSIjX/Gjcp9haWaHYBizkXhCFTe44oKRM1/Qg9IsfwD
LC4iAWDtIqYCf+FTsaTczgT54xyfHMKltImFeiID8KvGb09LJbv9YydDGVuShwdR
T4Hr+Z1pmUF1Fw43MpeyK1Rw951hhZVjudYnyhaI7hr7PfsNZ8MLwqWRvm97/DWe
wyhXAsKBYZdG9mmsD5aDCqAEoZwFb30ZLvMGD5AgjD0a371JTGpEwFf+Ur0iSjuy
dLiIWt1OcP0pNAfyX+8JCL1vfQLyLRI+QTdXyAqn854ya7ivjxhraFnJyUL4J10R
0KZ6jeCgZiLYJHIJSubyURrpPZznlNrh3hpItYRj8Bu+pAAn2v1/2RNRvPYyS42e
bs+AHOt09ZdN8I45nvb78C80pdKtcBmGrKn7JkW8x3Sb6FSmeqVW9lNO2nkZm26a
jNFueaEnN1KRnVb5wObv2CP7CNYJqJQ4YgL8N5VnAFSZKi5d2pqY6DQ1iakKbUZu
Lyrg4g1D5Ic4TQXJ1I9d2PlEGq8EhIIs4bJTU5S6xJoA20modtZuPczgps8LolgH
vzkg3grHMM3vFxXGf2yDyUWC17YWTyG9PNdAM2ESCFMKI5Q9iMbc2bunaikN6ijY
E+BoQaz2wjZ1Kgytic0+7Hxsvq0k/Cv/PzyIkdAp/yx17eQMmiV6YFG7d9qNVGK+
D/VORuEpSUkGrgsuYDeZ04kuwlxsOrzMhPz3LLnq0sHOvmhSgNmXoEkqNcB1XDCV
opoOfA1OpVyn5gseMDOtCniBk/ql/WxPDcKSR/HdfnzOmZ2biDaezpoQVgopYfgk
as2Q5y2yqSwrFF9NdnMV26lnb2QbH2aAcSHej7h3FyMlVNXe3wltk86JeJukFPeI
D904XRVdsFbCVJCo9AGE/jmdFueEgAba7js00VCW6W54hRhnqbq0DNCBN3rbmkWd
UTNn+Ei7aNglSXt1EwcNc4PDXRnCjfLCwmWb3XEfke/hQh5KqSoEt2+jVRZVYCT1
UU15mK19AbtCa5wRVHN0W1QRQX1X6jdpO20OQDroTV70rBDOf8olr9O77S+LKTGM
g0XTwS1UNBtwmI/1pU9h8jbP+UqRv40NVCZIfWJUQPhJnj9B7C7Aeta0kVhwF6Fr
GWLkEQvlGaUu0WlRejvxCvYKeUdzt0RZF2XUr4G1bE2ENFAKJDm+xDJHjiefHFD4
MuZq/mtFrAbYO82rgPIUxV8h7/mk07Y1EPh9TQ1mLpHbs7hrf3knrw3a9x7R86B7
cli7NRM2PI9HP3a/EEQA14GvQrdvg5uYu3skZ/8WWhxCUIYECeIFZvWZTAUrOatz
KuoFxt+/Wb3jCLc9V8t5+lf1WlfQRD0/iLcQLcwGbr0+8BycSXWjZXfwruMAMsP0
vBq/Ef0eGyT05ntTjatpg+HzWhI9m6Z2MMUx9apPc9SqOch7sDphCOAWnVnRaMtA
Gqz2lIutYqVU627SEp6VFloTdsANTsdG+l9toIWWwXhhNe/ZCVelY7VuPASiYVne
okjh8cgF4rgkHxhhgSrNGe3m+hNFyBIicn+FaHusRHeHJvd+2rsKzaVAhXkIBZRr
TYcm9uUXltYmftT4mrPiGhOWLUqF9tA20OBGnFBKkp1ZCcU9q/4exn++2zcM3pUD
9rtraWyWa8zcT4WiHyFWLFidrKfllhKanPrUAztsBIuOXM7TAqlvodaFNXJrQd02
5gRTfal+0YNa4oEMWFjKrHQtVwrrxn6rzNDr2gwUNVko1pp8PiG4clc1YHp2OfuD
25gWNOdr1OUH5IgEEDPUTd7HteTnNqgxDZm3pAPdfGRG30TrBuYQFMNypkzIck6A
4ueYM2snMNlQcw7nOh+ecvymYc2G2uSh9GVNm1wfeHaFx9PMi/FQANR2Zb0qkGdh
7kscTeanhJNvcwsO5wUHarrP06WvQYtnBzURWkxdYmyTmlSc0hZBLBJJ9XVo4BMh
y9gOIFjXHZ5S/E7Zqhdzqf/E8Siug/vA/w1tX/uZ711216F49+uHGQFdrUV3sHPL
P4pMo/hneZSMtAuWih5dHBDhNWBuo8btneREBBGqA9nA7jj1Wr0qJ1PgNIrX98do
4IxdsEVgZ17jQfZeFS3gIRJpbs8yQLwxS2fKlyuhHa8FMJ6ZvW1dO42gaas8eylB
JFNxyDVr5lE36d19rHMPYQ==
`protect END_PROTECTED
