`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N73t6X4zhfdKGSPh4v6wegVHn8xnAyocYJGCn2nG1r0s9x1XIqp9H5TfXUBh9VcL
Oj7MXrKKlWhgyHPPrv/76qCxT+n1HKgOIZ0WdW+aN8bna1jlgFPQBB1cGS1jxWIS
xfb70F2H8tHXQ2auOq7sknaMHWZVxNjg4GOx8zQZHraoW5jLPEHdoij5QjY63O8q
bVQE+3JOezDsDWAj0qMZPQrLYLB2sU0bk+Z5SmUMjgGrRuEE/wBxDIfPKiWgs4XU
3pn4cf3Y0q+5IV7BDRtH6Kw6VAXVwUrv4KmF3sYKQWDQUr0aAWbr1KYqmfSpHA55
iQVhugXK173AOBzB/A6Jat/AP71N5OHZtuabYgQtvb65gKHRgg2Ers1ZXUtCxlPr
ytRi+EovEVLRzMd4RxVTWH2RDlletZFDptbGOAVRG3EmXPO8RNM+T0yWcXhEbV5i
JglS+JHXH+MgEbUV8OpXIw==
`protect END_PROTECTED
