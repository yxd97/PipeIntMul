`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tLb7KGiQGspstTuNuJ9J6N4XFKlwju+KMfnXzJJ/UbisQ+RFo/TLfhkmE1fbmlr7
eXRRI4XGGdnXdrcPy3HRC64aFv9EDlPZEkM6DYeJDSqSpBAPbMUEekg1u8P2biWv
2AnLyh3vRptVFv4k7zwsq2Jhh/kicIXf6+f864qLsd1aaJegMrd7YPRW8Hksqq9E
l4LpBb4i3YKIOoPep0TIgOikAwfR9AepDtAXbb4fefuh0A6xXrNcYTH2prbqtGti
HJC28a/h+bmcRuiOufb/7I7Iol+LUU+G/Za5hh0KEYx6NtagHpXwNZYqALeAEnkj
6+LDrwMbJXaAtFGi6yDx4tBI4atFwGxdi0Poexa0dm1kCtJTNPH1S9dSsCCL3S+0
ZJWksJ6BTeC4xBhcwPg9mcUCjmUYmXkgX7Hd3MZ55KQuaLbt7uOrLigCR/Ho33se
7ZJgtfsZM/TXm4SSu3C51XUd3klO4sv0HJxqeMM/KWHtuLJQVCnRf1GmbktiWBDw
FqGymQhkpRWy4/FGU9lb0VFV//kSNXd5uZFZkX9lV+2hlIJruo4BuvXSuXz8BT4r
gVf2dpQ49fylNT+zSuwjVf2ldf3IjSOd41qpLhf+h9uC1wtoyp6grfDmdUEe7gc3
smyvzoOb2OLqotk/i1Z0Bl9m/ePGN1+4F1OK4Ib0+pAYidt5w5U4ZMdxqROr7tj0
G6hIvXPOVeHhtKJj1EH1zhxhWfKiY/aXeUg14E++UqidMbrLbbS2spPP8zvkDOzJ
T9uuN0erwG2uHU2LXniG+NWuwFXF28NXdRQuAshoLTgcCB1tC4vwZU0le65flMSM
i4RUkWc1Ej+/6cM9sXWYfDFLMGR0tDTc1/BKoXQhx1N6ZZqqcAJ0SQR/4HOa/hvH
8G4oibuT7803A7Mykt5yAE6NHZ7CiF26xFxpUMvxMthPuNHG4+nyzHIkcQ/IVdGD
wmFcEoTqDQ6UpgmprPwXjPlKUbM4dGQQvjLTZ8DkyF5MfyxW+NL/cnp75aFDl9dC
`protect END_PROTECTED
