`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NW68NWSYu1wh1gmKnEGeYJO8pX9kO5LWPkEWbCnjzQklDZetDGW4qRotnkNWQjq8
rkQ/jJjDq6M5ztn2WVHSdm22CIqXtroTWrQ7YSI2CoG0ACI3v5CnACCjJ4tvNEAY
Vpx4yOAf4MmtJJ7DMtApUN0Wv9+BCIzjuL5ZTtiFNyOGwWMoDYsUu5WgQfo8CPog
wIT9V2lTUdGU/c6NEO4Jeh0+pht8rRa73oYUQxjnscIO0gd4wDeS5gauwM8M01BA
zmn+XND7Zp7UmZWbXFLLmzh9HRPVdzFiiJp5nt4/y5cmVPiVaUZ3Z+FsseisGC6v
8I0Ai/vA+aG5ktrF34sWAA==
`protect END_PROTECTED
