`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hl+onr+6a4zK7L6OVKKzVP/3iV5uEep4vZ4a4f+jEyGJYtaJF62cNRBOdstbFAfu
XALmZsa6o5+31Oo5fTJUL7yBc9FuMLbDqzk3fKf45RjEfTTcgsML2QYXerAGIJ0u
hjgj7r+7J8OVkmIGJWCaAs50uj1QgJKSvlk2OSrUwn2MrlAKSs3cJHdFPEr84Ucs
r/wCuuhiNVvnImFL/r3mo8JcbdyhNNL9OhDBA771Xi38j+EEXQqdrbnrdcOdOsdg
60jX8h4LtXaRrS+nlXfrrvf9AxlK4yF9rIwCognK+N6xsXxFzQwyfxlbdY33zyjk
AVLUaRsHh6KK4nHBYC+JDBdTvcYJhYB10TXEadFCkFko+sBZ6DkCkNIbUfR2isPE
H0scBo4ksaCgGlo+W4OdRGudwvK5ZJpCK84f14sX59vg+rJKa6pOZuYtJLF2atHD
JrdsJfO3mdSU32YylI9E8VdHa7/M29DHoqIV9J61Wj0ECKoTYTk7NWc0fCTcULZx
Wu+EZTSXcB/UVRvSF5aQ+hU9GAs5Lu9vKKxZAUW0RT1dJgf0GE7lz/UGhG7YbcPN
8MDLu5J+7DURTiiaZa9hCjsVG2nXlYkU2aT0M/pYZuo=
`protect END_PROTECTED
