`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/5gVB+GNc4ayXFTr/p9HcCBcy5+YAsr10e3wHai3EB9GPMtFLzUd8X5GceC5d0zx
SXIPGXIU9FKpraPm2wZ2lb0lmyK37+ghId6A9+4Wk6muafb3Uh27wWrwGBez/cOy
HJ11G013xN6Fxk9apN4bOuN5R6Lb0E8Tc3cONzXqmcxCwRpmVRMdaQeq31uGsu82
j7Hnb8Bt/UDunhirOE4XM5xyJ+MKeYhZ2UkTWMFi1PE0dtLGv6UmEDNhHdq2qPca
BPlKHpv96+3OcthaJzjpfNJ2FTam2mWgy5w0DPtRXUIIOOZYx6Ma3DVJn7vE/GuM
KPajaP7pDojhftzNpJG2r6SXpdChHJazSPJZ1+50FlLW6Yx8Lcs/sGAW039UgN/Y
X8VPIU5g+SVb47Xh7SdOPg2cWF5na+D/679WmL22VM7+ouk+Y5c7BdtpEOe7UY5Z
vcQdtd0TVz60BEWnGg/IXtcpxxQof9ZzFQcer0gBs9Yj++22B1mCGldsMP29uMAZ
7LG9/ZR+U+4BCrfrkOXx76VnTYMJ2ixg3kFTY9BlQe6tX0ahFRvKeXgUznlaKlic
7oxyVOfe7axN52Q57lwMwjbRyX5GZ6sFYxCqSLogGcoINg/IP4DnX1KQEIQB6hEW
Vva/6wgBaorcwalkTMM3CynRAEEsJQJxtcqwMBBU1gHEEm3nmWnHLNHaSxVYCzV3
4kp7GaelSXSVOBjVNhaGMRnqIsvvOPQJJAX8sJ2pSQXHWxJSSBTi9pnvW9NQrXlv
geb5njCUAW8GiNAgM5cGQhaWs0tJcatcQln7kUc35jYnimrJTWZxEgzUnJOmbgyz
lpYCVhMwTx1XTIJLfnbhd2UP0ZOOSeqUiuZL2J1TaUsVconQsnUsz3bfLi9i9c5Z
Ej8MNeKUh2fRJbsXVVCUecLrB+Zrt5GYUNyCEFWgkvHlI1UJIEwdbIU8CNXbQR4c
`protect END_PROTECTED
