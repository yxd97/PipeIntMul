`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ZpNQxMTYdQI8/tz11P0M0xluNxRXoFdGB+LgVYA9/6/cUavJldGUveCCk0bj7bn
CYA97pHMl2sGiljlYJsyi16WvYLeIVKhF0th+mhO1bWA5hiXnUUisBxzkTiKgXe2
RIg7C3xChoIH2y/i2MpAydXqYpBq+ka2WEiOZnXMlgCSrKJ0tKKuwqYSmIICI6y2
3JkCtK98ctl6qWfCceclYoUXIbM8r6B8937g++63fLnaz1Kl4Bs0ObEtCT6cH5sN
t96jOKPEw7WCN+6FDjC7/cak3507xwECUSuRJJY0vBp6tZAbkCRN0yjyKWfXF2U3
XnXOgZcig12iJq1oMfe0s/aQnn8TVdRO74DDys1ONzBtI/9lF/pVImf8SS6UgGTd
QL96IyfLb4qvn9juYFeaGbdI8y2mmB6njeFlP3NxJrxDfkCdtmbRGBE122y4ocvO
O2/cZSVQyyATAH0EqsbThA==
`protect END_PROTECTED
