`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pB2yVtZpsPBkJKoXGdyhsUS0HD6kJaHNtMxPrZL4k3Kg3uxyrU0KXk+gJhskTpi
Q56zU/4flngiUlFnPuUE16PlZlANz7gR+W+ClEdzbek+qoEDktGHZPKa20uHxJuJ
jGGEth8RIK+bhk13XwkcaoRSFka6+uXh4Nv9ZtfkrNDEjKv04CFRMrKlD6benoe9
xFjUAgE5eCye/QMrtxUhltcpkJwy5c/5A+4XHlJEkjpw8omFPK9Zuh3vqnb3qDuH
QGShS7ku7g+svhXXsEI09cYHy+Cc0Aa+md9JcQTwuwq3BAT7n4bE2tOV0khY32Ty
Nxuh3JMR1HQh6xan3ZEctTs6KXRsCrBWffTR8Da6jQmmbvbUs/AVvpIGe8O/iUmO
HqTxUtWI7UY0/4NJZrYDBKbu7L//8kpxjoXvItkYaKuZtxWWX16+2hA/WrhbD/1F
eQICeh091ydHjlTacsCK9xn2TQ2lTV2fqlN3JUdOnwnj0x46kgMYI+rSkoU4kW3a
suRAncwfEibYiCujd4iTvHCiuFl3jRrhFgWEazvlk8WTd84oHF/9xCjVBhQAsMmK
cckFiB/romsxSm3+ceL1biQalBI+1bkdGvaPzIt0P6V9622Z22P+x5f3F6IBMMhH
FbtMUSwQxh6GnszXkmEI5FjizOoA2iv2u2SyudgJ2vs8n3W9ezVHFbjSHSfxyIJC
STPviI+Uk4JhAocCyEQ6DmZ+741YlMgRbEDEBgk/w1ljiB+JyB1Fiw9iKwEdjUkJ
gZ08KfQIVpBmY69ZrvLT9KxAeImWKy5CZsR12xnNuPPMRLbuDKyySd4P2fwTm1KI
hwsF/GP3KBsMDID9Wq525FeqdqBAzAfh9RjopseAS8WONA6XfFcdD6L7YyijOE41
hfpojX9MFpQUDdTsbHj9eKQ+yllj/PGyaIDOvNTDSrEeH/kovEhnx2ZKDKv/92ph
1Ngq6OguRfHKyzh/WwhLhKDbiHl3fYJyaOempjc3meFk1mwkX8rzy/ozI+Mp1DGl
sCP9UejG6b/n2BoKR6jK8V3vWr9qIfZPmSRq8kQluoNrZILRVxSOve8hxCz42Eru
FoM0tenu5OCNtNK37o1cAtsY/OCxWfyoF5hujQoqtK9N1LSLFMXAuCPr3k0o4HLA
lX9pJd2tI529ugMZyruxrnLGk68CnlV/7Q/8TmgMti6a3wZoqS8pwt33ixipHWt7
d4mhYHREK+pA0GdhTGBoBHYpoG4XaYODyaJpMVVIt5S0ZRiDV4cc8SAiyPeN466o
84QABHohwxve2BUppz+GzmNzJ7o7cknXUpx5qGvbKlw4P+V2cLxHX2SAs2/WI2ja
h+j8giAR4VFzBwvfYn0FhdHZ/LdZ3em9fcyvIPf3IER9Fk9lxdwuWWEKIhA6azMf
5sMDIj5WNftGCK2HWoNhfCqrAYrBh/r7XPTcOT64umFiMkq7HcK9aTljIQ4a2WW+
a6WlUAOVtkJfZgAvc2InNT57uNwjbeB8rTeEAADmJYOHZhTR0QS26LvlZMF4Lvbk
VxVZ/dulEZufGvFxQJPpwu76G62+4+hLCZvGjTSqIyvXp+OmoGlmwdHP3wqQzKHe
nJlgH5N2Mviskxx9Nx98XBvwumysujQWRLlzpSghu/SeDgCsKZ3JFGmulJ3hjkez
Cf37o/kyX0DTlOLVN72QrJCN2kkcZrkmPeq0UeCK+2TCZEEPHxd6cy3K0+4BKoez
yKcMIwZ7AVX9oHgEvpXIa6PZ+wHMBpoFGg0cn79vGOMJjWFYMa1LQuJgnVDBH20r
5iZp3avZHuD2toMlRkMWZEwiRzvcind1I+cubekqxTzgKnr5we8bPqdK+qIMgj+x
g8reB3SXVMrUPWkYJK5NuyRZE/tSCLeXSKq8JRAK4PpGFhPUqHF/ZcpIN/TfiKy1
`protect END_PROTECTED
