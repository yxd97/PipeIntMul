`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hU1cnsrqSzNTSHwz6eKrxQsTa2AqSe+QFp3wf6O+Xy6sd6pd3AG0mM6InCEk6Cma
uTRWfp8PAR6yUoCQ3J7yS59TZIOx5kF8a9CipI17EXvpf4mVDL2+tehaqt/UyH0o
X/p0hLZ663R73grkDOfoGRzz9Kv68ZmLnpg11fcy5IyfVOHlxV/BvKCfU3slmihE
mieE7ennaelZqjGOiZTvX6QAk2jfOgX6DeeLwS5fdiVo1lLqNm780VJyIM4gtiWy
eMpcKyGHfQHu+mr3VCqXqW48OyzzJ4J9SkHYHvK1mAhd+eRpJbrV/dfLkUX+tX3e
0ceiod8JnK2tRLEW9wKfLgnT4cOBsWJK+ucFyNgruLLGCSrjAZKDlRtUJXUnefLl
B7/kfv0o7eKmdlCoiKzUnfeDkyOc53o+DZMFSNYMpqSxM4lePh2AgMNWpGZL7mp9
OYqx11jQnmpm2u8huG1tSC95JgSvjqdH6lJPoOnFZgoWl1R54BBPWIMDGTxWlhdF
6LQg5x1VSZzU2G/+VYblzlEyfLf+fi/8i2yfqmZfT3hg0+VlwSsgBJ9ui2tOlj8j
MnWK9EXX3fTCBBRDpooPrCDiZuYTksv+13FaJL04T0k=
`protect END_PROTECTED
