`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+vpEkPCxkOjJ1NNoTks3T2pg06F3RIuh8nlU2xL2m/UlNk2ohY9brn7YL4mE/l1k
8FDVfbmNb58+bqQMeguyE+OBewA+Bnry9WkmRTu+K10DsL6utGJoV2jWLp8zVGaz
2oNOy1s5Hf5sTi/92otC2Et8PfKJ7Pqlfh3qy6gDxuhMZ7XKVM2FIaLPw0bLfTsm
EbYdUbn8rdS4IboV7ptJsjUWgjRvAYlmjqDAvbW0LYJ341GQXIk0O1YTkCdqfa7y
+mRxjCuD9Iwdu6L7WT6yyAQ+K6oADFPZy7acO2ENr7sV7iwOoJjKfhxLLJjoGjSZ
21b+7rmiLJAs5vqNI8pW1ogNKDwTEm3b915GdNNBB3UP54HBEmuOkjP2UO1Ov5VM
QBsjVIV1wlSE/xL1+jXgOfFJgfHk+bh/M8LduJhSwc3iQ1ZPJ/XzPYHVITzgyoJu
4mctyNCzU4zbbyEn2IB3Krl8O8BQR/Ee7nK1b8NGkFg=
`protect END_PROTECTED
