`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehgu5ls4b1KlAmrJBEE3DwE0Fa0sEgeSK0lWLnBfDHiwcRf4PENuuApLJw/50scX
OHNNt0SCZUxo0B7Kg0AmHQwLkq933cX/h3q70TiT5+p3uY2m5axJDUHIllIXnLUQ
hwWjVprufIlj89qFiPPFAzIfIrFHrNqtI+1LusbplzDms4XV7/acAUEIQTHq33GL
LZ+jvAljbD3558hWn2/OyU9EP5aMGRiH/xIxaMtix86oGnwwNnPf8mG44dUF12hu
PuFjjMkgaRm5X41gQgPjKHuILNR9OEuMhubiAC19NltKmHwS9cUsXCA4eEhQkSZz
q3hG1C9MKhUO97lnc7grc085sEHF6oj+TIQ0P5/noA8q7O82RlH47HewF1v6n2VG
2kpNQH05Z14e7FZoF9AzJSE5O3NPiDVi2iVFGjDxK6zdrauuXVoiBH2R97pV+02i
kmLDZaLpkg/gxPHdSD3UeDtYyHOLW0fAtikVtwq2C9UHbGu3x4wOVzykKByXc/Qn
7L5aFuL3PhkMTZvEyYfy9Q==
`protect END_PROTECTED
