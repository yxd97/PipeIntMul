`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LBSybOu9iFHFIed4EIWlZV2mKafLVSIm87JzJO2FqBQg2xRnx+CxUPndqCKgN1pb
XMWsJrwl7n3he612aD9zMsH3w0JJjH0YjfKtks2fXgADQDBbys9qLWp3porjSfv3
jTljytz34px72cu1pW8kfWqQjHjL9nAMgWNbgXEyBWZf3lqXzAWdY2YzucbLJvFb
ZrCboK1wJZkZ2WBT3zifwo9Qvh+UeaOHPSil5kowPCHJn33aKOiw9VsS/pjUEw/d
VylT9yz1fpzUOCqg+3EAMzS1DsKpHmwb1MU9acyN9gifO3mBBE7KQaGDl/wEmD+L
Ggu89ais4gW0mFEl0uunWDutD9tjoHDAU+0K5/04VOsW7g9xukz2gVBfSHTPSQAj
MYkz2UI5LUQPqwk4CNHKzyvmMKG0fOREttnXZgGYXjnWsiR2NiAgOxle7V2+53kQ
EGx12SftiZppDqyTVZ86CJBo33Lbf/IFd9nCJXUnPObr/z3/L8AUKQeiccCS3YPg
zUdp90n4coOTwLQa3OVHMH4JUIVFkTgjxas8wRs+zlOp9SAQxzg+4MX/xj5Qssv2
2XCJ9ZhwPXkGn4qdR4d4K9sjMWFM15RHdKwi2l/Kg0N+s2h0wsoGFg/q2cjoCcyk
+JmZHyqxe9kpmOzdYx6s0DUX8pBhRGfFGK88pN1JKKa35JhZBDtEhVgLCnDk9+dd
`protect END_PROTECTED
