`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFNaYo/mtuVfi9fA72ZYCt7aGKy/KwPXF86hwpcAzMVn5VSI2iZWnRRAyZSmQWgJ
LcUY1APWkQkBRfpSF1rmfuJqjtz8MGkrZu41yaiPBnhsAnohEsjDoFpMkkaGtPou
sZVHg0T4FnhGxwHWc+h+byJDzMaH74RqzG7tGaJ5DdAiKQ1HtA1yNVafuP9itLiY
OThSEH1kudvkaQkQEfK30PDPzePHkczHHBMM2bHCg3LJNqPbkQT8QbOr6qzUhPN8
fCF8xwoFOJ2SFfXcc3XCaWiEOSbiOr0wnRh7JbxsBgiSwPvEJYZpdoBzJPzHWQre
ehPpdWaA3oe62kOwhtec8/eJeSWZrNPRjy1lMSj/KfDWHAKtPzbaP4rpQrmYTm6E
5RgWj1Z2BjlkEKnybo7SC7sDe21OxfzEfIZkxL+S8K1VeVQUutWj8ucsCIOff8le
uR/WzzeLnDn1or6xrwMZ56xHscJpmfSuceFogmo21e/wCPUkhH4jpJGbuq53IPuj
ueYV1OV9h9VJSWzobqDuNCbCAk9z7gatQ7H53+gcLGGNTZFZbEwL1cspMqpdggTE
ZxeYhq5fkclM22Nxq35Nbkm9Wr/OhgW+e1ZIu4p1GnAA9fwX4WS3mXunM7F+iVtV
QmXO4u8vTf+xnFbVE5/Zlv2hfsCS3xUy09T/Po1NRRplye2t01Sj0eZQdHZxCgfM
L+YsM8hdj6uUVeU1twtwbx08/M0BKtq/XaHUTnajN+CMqTYk32u/TVXHUC6EXq45
s3N92b7aD+VvAgJamLD/jpeA4T0ABOy/SLgfe7hLBR29z5PJjE98cBK/ChmL9Frd
Jtqg6coHI6HHL1vGO40x0N8EXSHSe25iUe+7IZPYr+0j3PKdHyyfnLi3XJV0OaYg
g1/4ghVWDF+G2nRUuZZCoBhUYn7V1kz6/BlrVZi8LUrNp472wPivhZ2fnPyHGq7u
VRKYAgmLX1QWndULFAiQgZkME4n+D/+YwkWs2IqxMGl2TeWx2MwHJtqltsrRSO9w
mTCqU8D+aUeVncp2W9SQ272nel9i1oYwi4WJuBYW+VKbtYz10jCXkUTpPh7bLg3c
Wlaa5MqaCaGgzFB7UiBjR+UxTkOS7a3fHbZMAFjjvi2MzRZxBoMGwk5oFmv08Z0B
XDwyPukCo50Fl/+B5KCoropscgtuQt43q+AbxdkBrSYNpGH20Ax77ct9VwwZu7aI
xMU4jpQ0WfeJi0k/KX09zxA27Kb7sVbs31Rf/p8/d9SZpbwLO8oAC374kP+jp2yX
DxrbMhTAB1MwtTKiD26vZiP8UBJLmc98Yem7q+idW/F19RaoMK2eTA+53kjFtd1+
LtOtA48T+Cm2xya1hx2FZ/yVZz7D4fBBaVHPlhd9HCpKKs9Wc0hSFvRG6oq6pgHg
kkyvb++NInsKo9VUBb8e/sAb99CScSyfEMMM7U/ickJwxvoiD0nwv0acJrzAd5/r
`protect END_PROTECTED
