`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNDz8E79vv2ogsAwbd27Dwuz/xlfYriJi/42e1aZenllMblnDTlM4w+cs95dER34
7+Owd03dz77f6bTkAdGhAb4YnjG/P3r14VcnisBk/Hg678D6g4SIeVl0ohIycLE0
8vhvwfaUnhdsk+cKTbw7RZmh5WR1K1dUTNN3XneuBR1oXxX88v9nggtsvc3zBi0b
csqecj22Qte4c+xUEYwPMW4HDTizJFkd+L32oNQMF1UI8+C6uKtR3nsjHXceGkC7
bpKnEmx3hm/xV0bzjlcxgRITEMAj3CUb9g92hfIbJXdbPQ3J12/lx7KTuHcuWXz0
aOAgKwunsVubUOd8b5YKqf4i6Nm3QCK35H+RPHNul6UErtK4LVVtdh/aFd9sp68Z
X7M2OX9AE3hPKKo71GMP9Ex3Y7y+hgqHAdRzAmUGLiSoraom3fXsCEcvUuUN29r6
PAAHhrBy8P2DbAp3HbrC+3n0AP4gv4V7yxLvgfgxViqylSd6zATBarfC42f0APho
Aegkg4hxSGsh5YAUJkGPWhl0zt9yQYeWetHmvIbhl9nTExhzJIcC4iQtVfN1V+Eq
DGDOi+HEduqzoqM7CUoxS90l1qYhMHVIUEOy18bWcxhd0mc2TVPYGQSBi+I4OsDj
rhydgiI8WBq+YeM1hkAO6bMYvL5taYgZP8YGxNs67NS4dnNoKxd88w+qdqAAczHl
`protect END_PROTECTED
