`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jrTukunS+YKrj2bW0eEjHU4tbQruDkaKqRsNzF+3CPd3gdKvngpJ2MelGH/9pPT
+92+35mxLpLg19xi/4GAFZZt5Zr9bmnh0aDCYnnw342AuzhScXjCmGyXR9byC4Jt
0UnvZyZFXyC+7HS83/0aJ5xVRB36+jAry7sxFnN2gWiITxpSUismnfASljslCdE/
rViRabgwARO0warOgMmdQGtgS2f5NuUrmuKYUJ7/Rv6ldSmLqKCPLeEHYtACymIo
xO+OfpOm4NVUDTMMXsTisxsVU2vcA7F/BCtQ4NWeDDQvoUF/u1hbzWZ1urNiO1Si
T6D0MTgRmycC4bDfjg1ViqJ1Tcn8kbSNSy+md0R8hkBlZygRJOOBVYxg1ZoeAu0+
zh57bmqwb3vnxC0n78J6bTDvh7Pj1rCBL9KVTcf/XdI=
`protect END_PROTECTED
