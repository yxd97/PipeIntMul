`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGA30+BdchQ2RGOS4MGHKkM/Grkg2yOo78m27dpAtj1+S1Ga07MsmsQd0AdgVkqx
WBEfsF0Eqe23y1IrvQk6+dymfNeIZF/yRMy0lWiSk1eJcMi6UFEXhsRzJ/VWI20H
YcbPh6lbtLNLlPYegQp18kQSsYTHYw8UbLxckmUjXB0MbrbtxkBQJ49qdpKAmoEN
65nWs1e8xzn4LdhhpnqpWjBWzCh11WwLR0yfL4BrhK1HKs+uaX2hhwmlffGTcscE
ig+eR4hQbCGr2uK4pIGTnmeFXJEA1gFqXwGcGvTUE9byWC6AHF6Stc7NA0yOpJE3
HZjOOuz8ERVh2mG4urBP4/7JOve0fTlt5T5Ei7VWRVy4x49wkvRK5FLFbm1CJy9Q
qlZ+HXIUuhCBtzyGgYml/FdDsSSZBOM7IZ5XOC2wZ8XsvwJEBcz5kxMs4hB28H5m
mUHJFR6jCQjHnwpgX3uSl5Q/cnAZj8Ee53T5Du5kzdbDAEbJG190N9eAcRkSz+fX
NBZxpxNGBtwmXBO/f4casmmSxuVSIcbMeLThXqEAVhUmVxWGkTcp55HxTwC3gZ0M
ubmGFR47WNfNmgSJfZuqy83XAqvA/jlvThXhMFG/t7q1nJI+i3RVty8gudIkJZai
EF7Z8fUAfiG7xakHFKx4Swyyb3wMaPQDBJu/zrhF0kLvzBPm8pP2LxrHtk/45HvJ
l1cxoZB7DWEdn2B4xDT3nGjOBbOUUQkGo7zBLG6N2jniYU8wA3HVR88JedBZ80ZZ
augX9CMTMR05SflvEzFSgrwfy2mBrd+a8hEnutZm9KGhZYqAlmvw6tNb3r508TCU
aLQcIBbEpwxdRuHDIv9VpOygbFGELgPIL7+h4djLIe4POiujSi0VYD3ofU8WkJ1F
EEDdAD8Hsgntrury+E/zKS4W7peLVPYnpWW9lQ7SjPf5N/ZlxTxo2XCoq6qRH0az
5v+c1MYOvzDcsCmJEOZxP7xdvJviHEwBfp3I4NDtliPW467n5K7LkYpRqXtAtz0M
z0ezKI7Tbc4UTGHN6/ApghZ0++U5B1yS/eCia3aLdPJYBUK0PampejPwYAApyqAD
KhMoSmxpYju1PwGJZkxAraR4NsjefLuXKOMJjZEbh68tN8adw1U0p1vRS9peLem9
HfItNJXOj/oomkMrM6Ahzdg/FEnODJom/UxSg0kH49Z5MyRfLSfzz++punknC/Uh
/YUDnuQ4tzUvTQMNNITJyi5V89kAFh3mxFRNwTf/YkBKdyw5741MILpgA+M7WV5/
avuNWmraewCtl5uMGG75AuF0AWUNOO3Bw22WdPf2830ngjur27CqRQlprdBeDK9i
3Rv+3OoxhfxEe45Z1tC13RcfRBuJIzXWmzBrksJ1m/uXKuq/8iA3WYbexv3MiG8k
JaxR4wCvY71LPcEeMzIEKV5+UQcfTflrPOo0O+ONe8P3kPNAmNsXiGlbtul+QxdY
`protect END_PROTECTED
