`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Es7xO8IPNUnRCbNZxEWMNW2qLlrnajPp2cvfEt67W7mf5+dRNYxgir+raF84mDDJ
elXTcH299MN+Mg9SyHHLjVbH4SRMAjAC2KhpjN5PB6nSky7/G0glGyaiEIGHaApx
zmDkfsXxYzxQRipCcBjmvJf/dYZUrXGx2nOr1EtglO3WI4QszWXvZnvw3a4wcwqQ
Sy1rOdIo7awFamlWuri8EcRHkG/I1DPOuhIV98vpiQ42oRwBq11kqzEYiwxK0Zfz
zu0MCA2w9YKTZroIHFq8aYCHt/zCZBhcWSEcyBGrANIKUpMSG7SgWF0h6oLR5TdS
sA59R4s/JyL6aiMHTC1q8blw6aBBxItGQpT+EFeqcr6X59fCISyw0R4SXYUA3Vr0
2dRMiJIBucCHkkXJaAuQlg==
`protect END_PROTECTED
