`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D2FjkUET73w1LlQZJapG34/ffnOaAuxeStelvei19aw8xNGas3sTed50sxVK/QEb
D5CeiMdmZ6Ec8Gfii1uMqE/IVxJZrncctD5bu1Qf8YlthoQSIlYSLhOcUwteiN93
mmhrrD9DIXI8Kn1XqPT530I0o3qw2lbSpW4+4Jpmhp7hCbUa4kGosTECX7RrR/xC
x+aGxSFtkRiD1oB7a5H54DCyZLPJBkplVDD1/gBdDn7QGD6phtvXg2aGMAp1fCDb
3dKtzD3JFECqpkxkTrMQvaKpTMpP3JvfS0grpQgYncrzITTTBOu+gLre9d1s7/DP
QG2Da2Q1YkPxyiUwhXHcSURYxb7pLi9FSMmQBvIwuN4KCCF5aYbXhyoRb6EtHP31
0jFAPmbzfBXwpze0XFdxCC6XMT/bV2mwmD5or3O0eYtZdZxlqkbBsEjc/seLefZo
No76z6vmR9YQ3TOgjva+Mit6xSNzu8JURj7GxpwGjF0hOGtFI3YGQtDPHSbX4KAY
I7W7EDv7EZJjoZ/uWdi0pdTIW5noOc4WVXqwqTEZCPRlpU18f+nCZpq50EyyeHtZ
/ZD9S0x6YZmJrwy31Ev8jG/FWTSLcYYBNj8RLUEVcncsUHtOrgCArsIDLIp8/4V/
SLX7k/P4EMjpGoSjoUKLKt7EhhVrxUxaKRAybXRrOFdS1aWdC3vDw5qtVMJlCESa
ZCI4IutU5J1krmBtFuTACvNodKm40yAJ5KAS5/PXrk0gfDdu+n/d2rsBXLKbIP94
kQaBUWtjQMo4QaXIMs8RqNk6VXtCdTfqx8HB5V0X3QYItVg7L7u7okBwr0lMqO+J
u4ZYwFzCw+E38qYXqZxC0UCTQjD1PClrTfa4ZJcV44+OMxIEJ9vODtoTfv4putH7
xxDHHjYpHPLDQqjW8z3kVIkLRsm9dhh6HnqOMuqwg9oy4xooEKhfV1JCzy7n3r1b
mtltvtVr3+pZ/w0IHFFI824/rjIKKq71yKIhl4y8gK3d0nE6cE+ZGlfpAS8/idUA
ijUj+aC9N5ChKE7Ky67+dX2WyYeKVQ4GO9CDlLBzBffUJLWrUpn2uVPL5d6iGVGd
u0q7P0UBp0swDDr681llnHbBEjJWDJRVdccAd93kM0S+pvD0A57j/V0q5V67qETW
n310xlZUL6NEuIxnDhLwaW5IUbU3st0fJ3nGtIrXxz0Tgpg3IyQZoX1ZT52KwYPY
bZDN/4GmjOZitbB9IWGDIhI+63XeFU9Km3tgxt0ZJZ2j2WqOy00S85cD3TCNNQ1d
wUTo9Z6YRn22938MM6o9/TI/qKd1+/VAfZxdW/gDMtKLWGgU42JsnNOid0+9LONd
zuab5/wAfyaStLmediuWkJ4LwOxOzt+dOtoIcBWpS0UL+0jDxhOmhHzpmlvBO3rQ
jGzqp8FfWDJvDFgqp1HFSnrbTxTBa1WnEO0Az0fMnFPfz2b5EjNzyhyjBzu6fjGm
m3bQhS0dx/3Tvjen0e3UL15avhOXyXuXIPYgvNGtB5pasOWumqU+tCUFJd9sfxba
yw7wyDYxk+vnmdjHRn7qQRyRCUrliyhTVm2hkJUoAzlB7mQ1skuUbBWbfcmmBqTn
Xt7aEbtx9hNSqtGndVjIk/6MY0kPenzuCSz9lIg71Eu9hF6Cw+RUtu58kznGP1nI
xhccK1LXEWF2GLGLqhzghUTKF9gnWPNs4aKmIcsGvdPJHXKBikGYo8+3fogmjitw
IrFoIf/XLBi3LwsIBFkrZg+hMy6JtOUNQfFx//S5Q0w8sbzgnPh9tJoBarnYcq5e
nW7BHRHHW8as9laZm3hsUUP+hF3Y4WuTtDGjWI+YDjzVZw5OiaQKVTsyV0KFUZNz
ZZ/JTLjd/yx3N74l/X4qf4KouiZWRHrr6XwaKeJmz+wTtThZ6gXmS2a50SbWtgpN
A7WZP9aKc4Ao6Q94tWFr0uspQ5ylWxyFk/vGkyx072MN0QytFD74M3y6BQcRgoBR
z2MslGP1TNFF4wpImBtKI2Pubr07ONgJ8nHW24RfY7UC10fIiGXTaN/RIv3ksbEX
hyePl0m2bWDXVAWvUaAG9w==
`protect END_PROTECTED
