`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLaAKsjTjdRxyvpfX04x/2tapyYl7Lot1Nh7dmMU3U1oiRG0j4P0N1zdo+zqPpmO
Y7lC9vq67PYzWBxBdwAIWCNzEs6tJGNjRoRr+RuVlBB4aMWHZ3kpzYx0gKusYgJO
pbjl352X7hTTHmaLvofGGTnM9CGhLKq82nlszE55/GciN5D66p8JdtxMw+aUqDvo
lThFDFn2h4rUjHj/KAhTj1lo7ExuB4Bd0/rzT0c+0buxSJoihBcmd26U6U8BFSUg
EL1KCDQcwYbOE4jAPZPBtAt/4osO2p8GZ9NJBi/oALkW2Dv/LnskU8Ugo5kfG5ed
E/enRDjdvxFU6NryJWnflrQDCCjD0zin5uIJhLKJhd68V4BzznzxDR/oV1S9w6yF
FBjRKagL9DJAynwPf6dccJsm5n01icjHuv41ZSU+AQpwFQtWXhqy5fDoJnQHTdRe
ruyQUrQgp7m2lZvaSUrOlmzdb7wpVOgbfZki4Kz5mTjlLP3OPl7xa+anUEC1sc+q
RmAzuquOagYhYQ6Jsu4XYC67EtG3w+tIWQTkAJuQjyM=
`protect END_PROTECTED
