`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5A9t1MnFLVaY7l3Ve+LYPR4tGlsOH4eNUkJFlhpL/lUYIAwZpiEM3fyTyPq2tE5B
7WCCJ52nz6Lxw4dLh3yzjXNDgiFXpEV0iTxI5MzbWFq2h5Rxs6QJ+37QQSUS4//C
iBKR6a0MKYcUwl5BAl1p7xjgXB2jtPApiIi5hUIoEUCxj7nQsY2dwo7fu6aq8u/E
nFEgNhqM8toO/a48KJt45hlJ9gy7A3rLoYwjy3UFX+L2kdHgVBvy7nzinLwcpwHi
For2gUxUqZwCKpNh3cPtDfnTVNwKCWy+RNSo3LWTavDDQptHLPg5kCRyl4X/NIU3
xEd3qzqlw56QnzATmOcXtk/xvpj5qyMeNXWx64sWS2oWiMsnQX6j8j70vt4nnE4S
poSONloBKAU+HgVl3YBkZ6xUvVrx3G4edmzAiZITmrb1ZDGMUW6L4GKgAXnOD3oM
lhpg2k6tMrX4yNd2t5sGsHKAogtbJFR5lhJoTTtv1DJ0MZW0pJgMfZTRtU9JeGmD
KiKGBYMPATi3RYLUFklulfga7r+qeSrlHQNleEXekQiTxPl3p5PtDVfRSXHrRfUA
gcRA2XaCf7Xi2HL89Evqnr+qYokGZf1sVV1NXHMfhDk=
`protect END_PROTECTED
