`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4NggRvUVVz5y9rcxF1SV1Ek5CIMr/PU7XrxRdyKjRg+2bgh2wqb4RY+A5IZPHhAO
lj8Pz/ZRN4Z/IJOSX0pQ2alNZUO2aErUOG0QKWkX9APJnAynIuqg6x8N62kiM+6V
RRMlRRw9H5Pp7Va/vt3JZxxZ1F1D0iXgT4t7XDMs8tQbKxPXbmw8W+uLqRi9T6sO
OJH+kd+XH1vJ00JzSgXyWwToMdonV/7+KuGswTvotksjfp8e2O7ZSbG35wnj16lh
AHfBI0kZ7zonm8CPBTdf+w==
`protect END_PROTECTED
