`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/x9u/8qJBI7IvTZxlEbn4Vi65p0DmikS6krUjHeo9xMzt8dQkXrIfPP9pRztsasE
1YN4dKtvuPFvvrz0OLF+bFMAnF4EHAxlVkEPtABwZOHLkuimh8BvLKmR53+We87I
Qp0QVH5wUjNOIFxZlkjxpUwczQPUh1iM57srKEQTYG/FKN7A748nexoaUh6f5TAW
UvSPl7PcsUn4QIJOMP4gmrafwCVPCS1dMDfzlFRFb7zVpG2GrYDQDYecH4AJgsNf
EIltwj02w8FBofCBG+c5HHPnNxEketpr2zcAW410bmohNdElqiQDvIPmJncU9gnQ
NrObMgn1XOvhTCCt/hZYS6JLFLojfc4pJ9nJCZhH+85PH6aE3AjT78TtDYtt3anj
WlSB4npggU6qqP40um8AyPuJO5e79RgmJ/RI3dFFjGzqXSrimZ90pOU066eRxb4c
TK9xe6TT118JT2pgv6/E/7ZqIEtfYPAgiazUQlwfkx2frmAkRgOKGwHxVniWQblz
c5slszc6GrGwI2UpdVC/l9/V1RbBcKFF7DUeigsywNzviV5BEVo6IA8MqrSQ81V5
7CcMeBkDPRiQqBDBoI893p5+gx6sh2+UEgM9a6o7iV2Ip9DC4rvniyYri/bECuQa
+paoT8m3QrQuH1mQ16HxtoquhksHYBkqmoea71qQz0E3C4ogQamHjxSZKjpAXB4/
zOo9Qw2xGjs2MAxlvYWI9lXFzZ4RmdirQ25ecw6UM5/d5ASocLhAcwkZThLPZVI/
mqxG1d1xlyu9aHdgiVM0cfDqD/XMlyMR342nzM8yaIbLsXqKkA396TX0v5ymhsSe
rxWqlqVuZgwL/MlL7TGmeaDToC+TPyItcKNlgk4Mr1kgkSaQ4wy7Inx4EIDIRMg8
o2LAtUcvGw8mUK0xaeuQS//tzMZUbkGlP6AaO9EMdjmPP7Bb6YIuLL/IJEPmUfdO
U9ge/0CVFX9mzBN8k02aSPu5gpaq+nckGiiZWeZjT352j9b9DscSRClwj1GDw2Hl
gSJOEb6UwBZI4PsI2M0x5l/PkwZu11T+4oREKqwrb3zgvviFrwg+7celMy+qvSiq
9q2TX80M6LUbP/uh+aRsJzm+zKXQgsECf7jtFIAfygql4Sz3kXC9UqJmTrKWDvAr
+z3GQM+kY8+WeGCz54KyfRoGQUirROxW9wwHWNKUfrs7E0RLU0UM5Y6GsN40TCjF
2pFGRYH0haVwKY4OQF/HJW+Yw4xwl4payR6pH56ts82kp4eh1+gK+cYj7L4yLE1p
haeUU0FZXydykc2bUuN9ZNwvdyBKzYRvvDQ7WtoPBq/Iws4dUUzalbuWiRnzAigs
dlJ6zhVUYREFc3dtoMixljKkFxNtFfydFATiNsaWb/i1WcaL5OeO23SydtNH1io+
`protect END_PROTECTED
