`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XknKaV9cQRZwt+tBXsD5qUkv1xG44ZDc3kDPfgpJuIXHyPS2jm7NoVuvMWAmj7dC
ZZrBYdDj1IHpgtk47ome93cBaGOyjUQ+/L1HU1h4lKa98gKvXqOl7BiZwca8HCQ7
ycegyf0A59WWV1qd8oD78gn1wQcfGHjMgHwlxYWCSJX87yS+Xy0HodKIgrV3tOUT
dGydCu7A1/QT079IRx4ZtRqvREb2i/jPHljtFLJdMFk/ikUD7dtmpwqYXi49RAni
kJUoul7pWWRfT0kmBa5QCma3UtnGlfxsYZHZqEx68KQH2QpPeCPmREAHZt5MmbAX
9XJx4/dnrPwuLdEaXtmesOXg6BKtGxPBn3oZpckaHmd1vFSbwQBa4onkZqGU2Gvv
nzZIxDF+PpiEKB5Afdsd5xousSfchlHlJVVqVbMgyKstK5Goe4hD6XPNS5V2dIjd
eQnf6rfUl4xhzWG9nY9Xaj/Xr8pOV8K/OV3EWhkVeEQ+TPKNKdIFIP9WCCUME5Gt
W8c4oe3+4alEBq6WLWyZy1/uIZCqyvSgu/ZfmDv3BZP3cnuj6e2T3wFz1/8iViuO
0qUt1oRINZvpuZBPBHxi5dm1pkw1Hg/MYMRucTGjVAssO9ni1SRnEETnzmtjP9KQ
pIgFvYYehoy0dUFi6rEak4+fSPtVd4n+XZkoB5NJ6CEfAzM3ELXh+GXXjj1n0CVK
hyCheP+FX4v/7lpvnPrC8GgyBcCH1TyvliZLru5GMdMNjzYZL5+jTTp+XQWNP5Tu
mPtbxRfpN+tOiAXtNFQY5Y42TmVZg7cWCWIhv+Sd4VTNZhC8CQLnm99h5SPUpjLN
dJaMIBD+Bs0B7rmmWgPXhCRzsKduNoZ7OZZCYzIsVPY8ICVj3R6rfjbqsLk0DNmV
sO3LLxim837Ngu+WGgAOKZWM0G4wZQ+a+4VUMkOGYMsGOSau+pRQ2QOvjMmd00m7
7VCaVIl/9wcaWGA8zVqCUwPTR9JB05CvdiM7RO745Ep0iuSXyHCmTnfJxONd7FWf
mTafeEeNvMWKVaQw9tODHtWvvyERkLhJakrmo2X9lcE4i1O0pVJCojHl6f7nbWys
d/SDpBLR0Lf3eAH0y+eUF+oOMkk4Dmc/jIjZkopZx62cv30ut5W1zxYlCF1DryXr
cWV5TllX3mfrS9j+LGrZgomAG1vw5XF2e5Cc0VsM860rd/e8SHsSgg2g2QMVIEoK
NIBX5e23T+bVHTJovCWi+O3eIegZH8EMT+Dwlh0Ij7NRx8Hfsrr6RBVdTv6Jh+Ld
wbI2wFBB70O+ZT++wI6FHVi5V78H4Z95lHODtDDxylNsooMJPlr+w9WmW441ecTB
4R3qyv0G9RdQKrZr6zZDAh+ji4l4PnG3xtaAJvLx1Ve5FTPECvMBfIZjQ5oxYFdK
VKryTPPbggmO1GdTr9F0Wc3w+SsY3g2fP1CB6SKouiLKMtX/gM/41+Pw3DPxy+lU
H/rUcmY99RpB4paRZm3iqMiAXJ2jWwpPg6A6rWp2xMDflF5FCc4nGbfaTSHcAYSN
s5yTQ6qAhjl7nLr1wnXDBUXQ2kQk2hpDrhySLdlC8Mli8x4qeeSAmB1VGpkWbdGN
Hbt/flfHfiQ1zNJC/RUJzqMFuMpS7U89FdOIzzbRAtRFDF5x3LT2eXsrrJw/b7M3
fXRgEbA76I+Noc/XhEfWhPp+wY6AMb8vtRO1mB5YiqQaTnBKR1udzifZ3GidDcRx
t2/9PIT/K88/1IC7IohllT2HL+FmEMwi6vv8m4zlgkPQ8/OSK59ETll02RMKW2Ry
8qGpzdwD2t5aY2XTePygLf9Z5KiiM3wLsLfqBAVGk8P5gqkTvw3RCDKpksAoPfCA
ZtK785DjtBfR3Lw7WM/dg6d9G0lD9Tnr5EPiuy7UCqI=
`protect END_PROTECTED
