`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Od3c7dxtkEvlMenBcOub3iprkQkgHZgvrqyim4GnKmUzPUGWdj9Jvx5jXHqUD5zp
4S9V51PFeo1ER7EXHwx2+QpXC2GIyYOwBo8ZBoRjHt8iCRkDuNoc+aBCs6OTvJnP
AdN6diiXMnH+XpoFgfgwvKH6nGMnS7kODE+RqOMnjrdgMTtvEsPNVlVsHUofKkkv
nAU1h6hwg/pZfg4BToKCbPh3ruXe3WEdNtr9DbQZeYQjXTld2svZfoPodxnW8nTB
RzKlbVFAOW7ZGMs8rQdYIqEmhD0i131bdF3e14sdvbTkGGOvMBj/NlYoTMgPNP/Q
P45TZ8E5W1r6+/Hf+WS57g==
`protect END_PROTECTED
