`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FSBDqpdpKfUmy7gTU0FLV5c4WbBXO2oImmQfVNkjy+Vj72lYumKpcbPQsQN/xxoC
KPB4+g1KP/3E+wPDUopuh0VGb+GV6WYX3oa0L2dKgtkZwizoTJ0lwcGU7FagMhgK
yutpw829/MoPbzgXxReDkHnT8jW6mRp+ARqFNNZg/DxMh5iaNJ+wJeWQTRGvty29
acpg0Azt6HSD86ZScGudh6rf1mgwu3lp7PEX6zCaZ6x3I14PP2uWoU8fRDSBTYTk
t4yql5gW5MJHlpz5EMvPrCrXSnxEHW+5I6bfJh0Y5+NjrwmegPH1vtVY2nY+Tgad
dw6ZMmZbDxYJ35tBvu2tIU1+vIVTcm4DoNSy41PrNBqXvnE6BWq1CFJDkSvtg3Cw
2k3DrD2kmdUozzUllj10Sgut2UQo8wCtjkHAIgnLXeMUnzp4MB05vsJ4azUFgtxF
XyAAhtpKMEw3ZSqAyEan+9NcKCt/mRwNswpUlPVts4MI9gmVprLWGp5WTDNhDR3b
UX4kqBXagjp5vBibV7R6y6UNhs/N4kownP9l1Ix2Bq15SSf9+JoCQIMOjLQDs4Oa
qIa08chwLFTtLj5KMKw1idKMgZ+urAD1C2xnBZ17wA+9POz5foiL70InX5IfqTmS
6v1XtY/rYfT+RegeEzIZ9QeM0D+VNcZZUinxsLTDVYUOxRICNFrNGUPI00jGuUGW
Rib6p9/hF2dTzVBnx12PNA==
`protect END_PROTECTED
