`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eXrEnlxcpANy6EzLl469FvINnHztbUMtonCHZ0rQsDnHq1JIagCH/WTtlmmZV3tb
AEKqQ33YSuETrzjohqaLkQLRjeyk//Apulfl4cPHaU3uwPIBc2lOSA5BD47JIv1s
O7MqPXmI4mO4l6NjWG8cFPW06EjzXIYpYUxGIttXInwquhgSgQMVFJMmiY0tGNAu
u8vGaNwvdpyHKuB6U7F6Zge1mthjDvfVqc/1gSTxnzrmd9BaQX8WMyR2QpK5L5vg
tMT2TFh/IuO96PcyamFwjIgM/SvlsXOC3Kb73RBQdb7oa6NOEp9EyydjZm8amuSm
A5AdrMuI096fHffQb1w4SQ6DeyUOnul5HzKUTmJUTf6LAIJ12QLVcFlMI8rYqzJS
outTnjREqjOuAxP7LWxU5EOzI/9IkzCCR+4yIocdS/DV565/6Z0LIWkSd42gd0/j
BMZYfikMEsfGmNyi9wXipgEqaH5PjjU89Sf6KrnX/yXjgNdewVWayyTO8Lrd9IBl
poHTyCuylRPWkbn94XDMt4KRZI5KamgzMdGqU7loWZIuQI8zDR8ObW7gI2RXZLtq
UAXKR3h7S8Z/m0p1EHAmlCVdmzSBKXUGsYOrM9XfSz4+5Mpg3rM/XWAn6OUN0lpg
f+s3KTMsgn2Fs99pScrCX2qhvEIf8rbM3c2dxbpPrOvtjdiIR0QOXAK6HJCElHQA
`protect END_PROTECTED
