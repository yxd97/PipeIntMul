`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8T7PG+v0VwRDM79WbPYtDBdcnGYYKikzrmurLyv4sZrny6zh1dljuDBIKTbwO/i1
6dIEZ1mzGnjCjueHDGOiT5BCDKlaQZWJw8YfOKKXOSpYXjMIuMQRJPTfDfvvbKZW
cWCb8D5kt+pYM2DQHlWlzhd9o8WDLFEShG5ZuSwlbYUm1MDtSvsFKvBHm0Vnj2P4
pXtyfhhzpdcQXCFNHiiPsk0hkaKhvTgu5y5nFHwpW7AOSpa17ay1KGVL/uG0GjjK
19jAxG8xgM3nHGww3/4CCmYY/AkkcxLWEvhWfN/3PoOrIhwvQrzknDUnlzpPZ4Zh
cu4vhYCf9gvSjiqrPVab1JHw79PWoNVa1wmcqpy2NQDXR+tAaYytjdhk096ZA3ob
4aWPVbP0KIwWbkkXc3RfzIoelA7AoldUmxRAZsoySSF+Bh0+7DZzPrExJI+/P1la
Oy8z8DMsd/B0PeBshftLVwlMr5UzxM3B7J7wfPgsUkEB4aL3sSekrgrF19scOMZy
XgHZ1ABfFMcyxRk9pwjnsHR72pNntknAoFAQYXAcw0nwOCUHU/VpL9EGKw11ltuv
kXdOf8FObNfESCLrQ67WBWIdvnGc2wzNY6fcKpygtcD7aP4Mdmo8n1qjn7j81j4L
7rgk1MFhiNcUvRxPTdn9A5T71+kDRJCxYiGI5DGhqQ5OMKq6H89gNsDNCqyehAse
SHe6h3w1uvcZ37qcawIPwT9uFwyqsH5/iZGF18ItJPZdPpWRYb+agRHnhLcZ1E50
neze/X1ygKhk46yI9sC/IBRDvGJ3OlK8IiSKxHUElshUHSrF7D28M0RTUAV+pRCX
w4UU4kv3qq9KYjTSYb4gIYSfW1zc5CVNLoqzlWFRdlJ3pS+MnXgxbVrmqSjc0rCX
rehMDAf/AkkYy6vkOGI8e5xnq3z1QdS/LaX9IM4WenLUjdbNrc+1aeMQ1qjTf0eC
Vo3G+/3i4NE7H5DYZ5egmibMTMcgEWsc12doE+LcPjIKyVUcRApy29IQDjvnq3x7
CJnF804WOUrwK9Q4yhzHtCnMJkiWqkXqyT+TOz8EO/fyCCXWtRonf8qG1quKsBBG
2a+QtkmPkn53c6MYiIKrMcvgSPMDGoS01+tX8U65wPoJ6jB3G0LTiaqB5M55DzQe
cc0RmamMB4KPk8U2860WGyGZxFGp+vqQwqLDOXaBigjtw1aEaq1q6OnkKo1cilfU
5OcdSiqdGZUZ/YBOVI0iVnkeFEv45qMtSjyMbLn4ZSKKiJr8nN3D/upIxbVCo7+H
iCE8TsTjydvjfx2sAQ+SpxIC+PjyPX+uRlSqkqqsh9S7ub6FTzt58DDsoteZyGMP
XcVemU47LbiIfacJQqwevfpTRf6JFpvre+pN9GX0Ga+QAxheJGmbhttf65TJHpBF
PtRFyqCxoOfXjWTks8WQT+OzpHoBwuT2B98V3r8K9zqam2pbw0xatWErWjmE/Tda
Voqst/V5zan/z40x2aiMEghjs5n3SbdYqYpnjOt31zapxqrE5cdxb74IW4J9xk2j
UtkNVSk1c9ACyouD+iXeexPYp4JzuuJR5YyOtpYZe4qiDB78T3hUgqZul3qpV1jW
fS0SRBGoVSc4xFgnoAX0zq+2nBjFWFatVhATpqkBmjZujI3X3BEMrwGuJRVotXYN
nwACerg5Uo1feZQGgWaW5g2IhSkhBmWuhLOHv+bQOW5H6W60G0FyvFfhWHsfL8BM
emZJoYGO//VOiPt6WurLcxSWtE92PJr78PFEI4w+mZ3P3paMfPFK4Oobwwo9qd2K
rRj/a9eFRkxrzhvputhZQfAFwqDA8OHFNj5fUksQyCdbd1t6pIRrdU9hExlgvH88
eDX90Wbecg7zQsh2Q/pnAT7Nb3VabM44XZ3CdxGUUxTnxjOhozku3lUDF/XpUDmy
onsvgc/YOwywkqLXVeRq3hYYhfsNSKCA5JB9XHc/bOi3vC9gh/Xnzb6/ZZFrGpBS
uoho6gRWqTpPZvGUNniuf0Dv7MeKqtUZTX8QLAnd9MdoDEfBE/90rwKHTbUz6g2P
I/lIa+04sR3TvDqqfj+bDWHIXxLS+99vI5J9PJwwp1lb5drMM1vMsuGeWikdSHVr
SM6ALHHjer9xthj8U5vhn/rJ/mGIoB0yq5mp98t/yv63GlJ0moT0Pmpcwtx1EANP
UkwAsrpCijbyoARceBt4owZD621yykwjLNC6UJaPrT24DYC0rI9xOFbTg8vbN3cG
dJ4o+NZ3dySVYjCwBZBIo6iRnPLkbRhLF6687H6+2vjN3LSpj5QqqAER8B+pxOWR
Xmz7TYbEz/36gtOKFa5Bpc0OWIMEyf8rIWPoZV4uhQc=
`protect END_PROTECTED
