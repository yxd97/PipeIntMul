`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yglHLuICybXpjreMZ2IfmLX/1pk3CGrhlCRpAg+n9oiNsD/ILGden/YKREgt+2Ka
dgd+SEMHvHRGCrjb/7GdvkCwkvk99z9plUxwQ3BbZv7CnLkmAUzQz+3N5bbdSbES
rIp+o9bt/vMbXCzR9d9z2lJge+4ThfCc1ssiFqJTn6viOK7TdpGDvX8kTEPsqVyJ
ww5lAoXPSVuzjuANHt6ry6N1IivzaP/KxTJvoPSjh9PyGsEzdS/hzY5enbbBY4YA
hJRDTOyCBoGdmfsSRjnNfXVwP/oK+n4CowAVpSHJRxHygiEgqpKXDhFT9sZuQAk8
Do9YNk2u4252l9AJQGbpXu/GTW8r0Sp9YwrY/3gkVM5DoCA/G8bqk58blAdUjKZ0
8/+7s4ehOsLBnNTywr4MYsFg+auih+h173rloUSstiU9ZqJryjC2zJmyhtqA+mPn
TZthJf6kfHy8Hz0eBX4WT52sSWvCjyUksYK3W8hOP2Q9MGQHp3Q7iLj3az4Ixr5z
`protect END_PROTECTED
