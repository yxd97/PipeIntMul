`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/Vd+vQULxcDIHjnF+xpHxO0cc6JZpUbLPb+Zn5DkCSuJyZojolLBu65wJwXj8fm
YjYZx5ui1k7U7lOnGb2lRKXOMXDASoYUnyoglWUPZ2Iz87ZC9JL5TPXp7CJxBgmD
60XmQqB8ZjWQGepu6oHBDrgumM2Ts9Rg+cnOk+qWxszs1ZsJ6U8OHSw55ZEhXfnb
VlR5y7SHpUpdGhu7qM4Tlv+rjXMK6I7Lqb+kTGUq3PhXsCjV1dJKON3LAIXdwnyh
jzNDoa6DitfK/b4qX/YhrfIcCkAbXkA10tW4d9Foe1u9+k8R2U3GwoxuSP4aglLj
CXaPxg3CmAaJAEeEuuoSRYDJOiu/1UIrLoqz8SpfhwG0vFmuwypQDCUuyzchhFqY
EJUsI81jkzdoktzlFnIADtJ4odrH7Qi+tXutH5AUAPn8pURYaomQiLkrGZZsvFoa
ZGLF0kYtH2lfhGwnGASbryEM/1/c4/Wkri6ZZ0P9NF+GyBXEQohR0IGWJ3hHed7b
`protect END_PROTECTED
