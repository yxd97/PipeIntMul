`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3E4Zb0ZXh3XZYlYXjd9zXgX7c1e9kStY+9Cy/8oa4JoIGkvYP8l9WFAEPVq1qHV/
d/b+TUJ+zulXI+tWZTJJ8kXvH34VGhrqf3i+TLsAXfkzjYlLToYq2TsvGtAEcHm4
92Yy0g2XN+zfRFarWHF9NzKBq2U3UkNhzv5xRCEt2SdtyefRML4Gb6o9/Wckz9/5
E5Y1oWS/OJ9HOEX3fQlmK+7CGRzyVdGvTE5l7+cudmJxuyJquRbShgN6Ynzyn1Gq
gDmhZK0+cRXK/+IXSMiwh2RVU9EFX0mVh6YrWlKxeh+Mej/f/3fNBqUPQNe+TiDE
LCTHKRwOmd3yKCdetcZQwqo/crDwQ2HkTooIswRah32X6u+NJnoxh7j61NgqWDsC
ghtRRcQ6sUZB6tgcql0odr/sze7ZLm10Zi48yxGmg6tyLrhoY/onnXEHsJMIr7Fx
uH5VRI0rXBzPxkW/LnFrf2mOC5ilcOdeJjjwQVkbUzGiq7Nuu7oFaGlg9uevTgkO
TcU+nFTIgY9pf4uVICfV08/QGa+ckqX0HHd/VtRgZLXuv1o2tksY8N66uzCHONSD
ilm9N+01kK4XAlo9KSGP0SJIZaFBtiwIsHr10NObeIS/yTVpKY/Cr5yb418wtBYQ
skGbeoEL1NVA4YBQsD4S2l57/8Dk4V+EhtOShIp3LLYbiqSTd9AyDajoQOpxWKlJ
dwsXD0BzqFkzZahu1Iaf5g==
`protect END_PROTECTED
