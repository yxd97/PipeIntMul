`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVTGs0Xgl/YGMQJ9ljC0sb9PNcSNg2KU7ZwgizkpSwjt7Kjjgc08baASF5Ty6NV2
jNIe+/VH9D8oNtSceryP4e20U/xbYXPDnqYOA3j/XVqkPlh9+he+SPx/5nTJ9cGg
0heWzVB4NuiUsRQikB3wujDNg1AqYxdVql4kmiHihI+DyMbg5I/gBQYvPE6Ss+tC
Z9inl5vvfJnpqhrVBYVsO66Yjr+Y7QBYr6LOsWoX5APtUClKKNmTRX+Dx+vnONSJ
zlnGBpt4oBPkHjEs5Q3suCx5IZI1V6rBg67pBq07c+1RH+D2A6cqKs/hGUERvrQi
cnzAanu7zDdUxZ+TFVsxYUflZ2inbKb7JLP+uVEcrLNDYF1sSSzGGkgUlo0vhclQ
iE350gqWGkbY089wdOp+mWRcjaubQOdm5oOPhtlAkj4=
`protect END_PROTECTED
