`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gSR7mbkLy91B59piSwPwyJ6H0cgpMnCOqK7tQKZ+cLX1xVEBIxPajkdRY3IofEML
5QLZZZdsM+UsXwzAMq+sptNBWJfU7ViIyB5Bt5CqCrjBxh+u4gSIpyp6C6eBYG+b
7b8bw92+yKVyNN/8CvW36t2rt11fqGTGJ6sgH4oo6OUQb9fqZG9/nwkqaI689ttB
Tn33RsUn9ONd0i9SHK3gXm4xllEd9wup6tbqoHeivU8smbv9ksy3cmA43fePwBv1
ZcsMe+HxFaiRJY8LdD7lHbY5FgdAhm0+wCNynK9vUHKOwJENBf48I4LX+Ne/8iho
BrRjIl+zqQRS+RU2BZOLezUr+ioZNQ8c3104G0v+y2T9IfiBAM+9zfRnlZJ1aqeU
ZoKKvMuwuFXqBIa6PUJy1W2hi40hj+f3wFUr1/UB85UB+0Oc03+9RQF9AmprwGHg
n9RKs58BP3R9HPPrBxVZrFDTGL7668YmuJMiVpRR9PovPzlB/02E7+4V9NsYa7LH
`protect END_PROTECTED
