`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rBqnlDWbzTpmwTpL6CsO+7maeQtp1IGSzsT3QMtLg9xtoUflynrM60PY1WjISgH
014cBqL1uOt/lCy92JV/wBFhz5o0C4dJERfEJ8PZzXD/wp2G7BLuzKhoIS3h8DCQ
hAVo8m7bRK09gtStN0akS+FrcqkcVpS1piKxV34nSlnLyXhr3r2bd57FjyyNnncE
GJAaOluxewx3ka7bH381ZuMGnxvdIIU3Eq5yuGZAm0hk8j0gZM8HxrRGp/MpJMHz
qiTuxSaB1LFAqDKyxwffAbaYqHTKS3FkB9BV1YdwSCYkCmP69HQh7hfc2aw/c551
1Ukhjn0mqfMuoGDfFGjgUSXauas1TXI6RIWI2IwPj9QIuQgculDy+AxvERAaALRO
WHE9JJbLqUk2NmiNEo6mbDfXR6emmvrWFgIrWAJ8sGJBh6GO8H8nUh1o0SV3gHRk
hvTiL3HgSlUbKCUlz0vzxfZxSLs1FbwzYZn7g+/A2KJNEvCAp5+e3Xj7g8tL+psj
foqSMpQYUX+/NFw5EOx/aZHOZH4/8y7xHBpCr7/AmJHBWR4pdHoHBE0wRSJtnQzH
dmLRLO6/h/I50hTfaS+vhw==
`protect END_PROTECTED
