`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iaaAxHDtOqk9r99ngKMJOGEWAccgaak+NElP4oJXNAVA7RpozGXB2l2tmJSS9T2H
AcVq5/cbS0MjHzbbU6HzhjMJoU9Whyz6g9nAcCBTs+BHFdKG+E5qz+QEclEzCgxr
ht7zDKF5orcvY+7I2Zy/64pz0x0F/jn3ViRa7LUL12EB1vDKfMHMowa3yfag8YBK
DlCBMjj5z6U+tEZgn7lr/Q7oxjnlSI6bvhpgCqvwup28eVeZgdISbwRagN06DHCV
cW/jtm8A+aqH3gBy/QTokzpslSINNRnOiSRmRjpvUuYO71IZpz6qe7bGCkKadj3H
1RtfPoBgeRvTzbW1qLLxjK6Vzutzcg6TGY7o1WzycQ5SJRd5pcx8pna3gatUflez
bXyVHeqTUnmYsI3wpG9li+lrIzklnxtcAw+zCmmPopJXlkqEG/nATW833zjxNeiB
J0mgjZH2SeskOKot6uHR6ZLYCkYQFtDFJkYPu0ywv5mej4XG/q7dIDkrOXHbtuUO
oEILCjPO4EWZdkSxhIWD+DizBINwvVVrI2ZE0F2q6YUs/rhx3I1YXz4L5fW+IA1M
vn0lgmYILejfkWlKBaye5jIvJHCl7jPmDWmhro+H/NhW5GWMjD74YVVshXe6kxgY
rr3+gXDA2yMSshlngEdhHKH3mBV80ITBDCguZBnzNX6sxiGo/vHGJQDy+OZBccwb
ydtI4hK2XFtFNdIfjBNG7scWF6xIZC4DANk1h9YKab1mDopwezUHKMus//Bp/pby
5w8AITTV0EzlnMhkSniVM91kiBumqgOoZDwXLxIU48+/5Cg9NNPScW3z4I8gxLi7
/3rQ9s1d4HbCfppqimpU7C38kWTRDDWAEQBi6exWCwy6YRQpAkGMFTCJXNzEMEsH
wpYIX8pLpbMlxU3I1/OGvkHU7nmLbdsRYYCnOLgWh0AP/oq9R99CnBQJB23tzjG3
`protect END_PROTECTED
