`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rx4P4LRNlGhjtSPDhbfZ/hqlOoD9YUEZBqf7tEQe4A21Ag0VB37o9keZZhB1u7xP
/leY7PwzMTVRi9HLS3XYit57ZfLNVzao1mabXKelJRIIZdnvDd0OsHaqwxL9iv3S
clXabht6rZCebAvp6iqtBEulDMnSm4k1WdfG75PcMaKMiUrw3EqiG5vDFjoL18Lh
2LxTfAKU2zIjLq6/LAbiIQvEEJRP7q2OMj7fBcw+Nup/hKbhrMz8PCihgi450Fxr
h16YelBEi/Dcp6oGqoEU3FHTOdgoRyD6CwARJCvqINrEtu4dEhSjdLpPebxkPLcd
YAcmEiNf81WAXbmvhlnDUAxOY/Kg+r07n5UmO+Nfid3knkkUBdx0GPsKLX7R5tUT
ouvNOsm/9qaJm4VavNlCC04WAD41VMOJsle9BvbpWU3Er5kPNjZRsPAq8tc0GMD6
4RzzDvoL+r1byHnP+VfT9qu4D25g00mn5/2wpoDoJ5r8+Ud0sDPV0KvOHUzGFZ0t
SROWV0OLxIrWgbXw2C2UAeCqlwIa7CnHn/ZdzEOzvTuMTHdRmz8tdpeXNV1QtEia
9LzHIcpe4ACHFyUNbOfU5aJpS/5mCcursTpOns6r11Ek+JZAh1NqFUjbArbx2jSl
1LM3asWD5j6sKIdPTg92xsz6ixnFD1hreFwa/NZwwf8T7bdsufpFiqp7oWeM4t1P
IdsR3TOWSyl7KWic9XGo5uDHEVjSASuNRtIcz3fs1KCIzRXELjoiegS0UDNP0Z/j
eqfR3IDcNpQ/ys93tLWIXA==
`protect END_PROTECTED
