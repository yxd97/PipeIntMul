`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/SBx81MaeHB0NXVAxI27JrObcf9/HRFvwmxD0OI4+btxSAogKK2klXMZGY5hgx3
bFZfvnvSjdaLWehtasAAAom0Mulz5AN/uqVWg8tha2T775PSji9HLzhgmdiB6511
S/cJHU7VUzUCDbex1PphAn1IrQ1cj0YmxU/rHAHb44QGq5n54BA7vONcp34MfzmK
r9sOtHzceR75XSuw+GSKbjznqZPcr5w7DJHnZ+OEkdK5wUIB2dz8RuENqDRiiQjA
5zQcu+ZPrkpPtrQhs02Oi6Cvbo5D93pFuiR2ZOpPjx2H/4PMAxJh1LZLKWD3CTJx
56+iJsn7qPNNYyhCYV2iCWgp+0fx/awwO9GF42dWWdlVCgYyptoorR23Am5v1ZHR
sGMxbthtsevsryOQn9h5DBzQX7FS3JynLyiRk9uUCIrHLx1M3gz3RtrRxF6hYf37
j9GliY1EJOcK1UhkE+Wt7aMhVNK+W8KlIbT3rftWAt+9r3+IVfSWl0qY1PbMktIU
`protect END_PROTECTED
