`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29K0oeBnSv1Jt/DrPKi7tJ+OqqxuUQwF2elwSLjRo1hWQGKeTVLeFw5YIAfHJagF
PfdS7jugBxZz0Gv/UZxssuoPe/HspNTUdZ3YHcxaPHpLK8vhiOAtDrGc+tCPz4Nc
tImEQmsdejZaxaYIURrYzw36NC3jPLvXqjoPDzDZsyFdzTKdo5gdClxPSwM+fDs/
KZMjv4OOFNfSUSMOqKb5y5Oecw2GXUrDpADtE0ngZXpNKIvQnVA9yOD3ddp2/rKw
WBy/bt9p4hhcXcCQpJcBoc4MnEW0LlEX6QoLMpzLK8c2thopE7LUdu4vGIw2U0St
8J9oT9TqI4RHCTmxGbOO6ixojk947wmwFv+prSx9mvA=
`protect END_PROTECTED
