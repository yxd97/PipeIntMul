`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4KFPFnI7VFXGpnoaJf3WmdHcasxJeVapvM067ogJ+XGXsVhw8A3TccODG+e/LZDg
5qcbcSk9sj2C3clXDaEWDi4/b4ccgbmBpu7wbaY23HU4rVTjwAHWUz6lA0FPg6O9
6htfb8Vu8w99oJzr9vVNkkfDxCougRqxINbDUi354Lxr9410aKvxpNtBxtl6fr9J
ZAYxeFXzY84X8eXLmKt3ee9Yi4CwpxDe2VKe6sH8dnI8nxhlWxyE2gDDnIdzMn2E
VebZWnlKRKgldHpDjsliYE1gsiVA6kPqqDqgOVNBcf52+h8b+8uKYM3bQQ+uHxG4
YQJL9yONzi1yGMPW5UfugFR6nR2PYvuqmyWJcXRC0PHJBiYgOUgaVLdghiRl0Hgl
O3H2G2xb10/eAbcc0wENXlj7E/1suenBL4Y9LyBaPz8/RJnro6V23Xo6dXJ22oGd
J3y3jLZl2haV2w21MP2/MKpGa/6iphZ3NbPUFIQxRotYdxQwUpzZdjI2DbCm3zOS
71CEbaBjcwc928aEUZa61IJbd5ILU25qN+F+Vif5LniB/zyE1PBQlKcmTOpo5fwW
+wO54KKlYVbTJOBkU/KU2Eb3udnxyAyH5P4E39L5YPepbD89zFirrqhRV2hjiq+G
p/PBRzpIJ4Vjply7VlA1Fc+1CRN0ySy4DhvbD4mqnD6fRBeTsFKoWgQ/0XaeQaT2
cJpKi3W4MZ3aDKuKRJxL7E14z1K5Uo93hf2PBbnRIESOdaRy9DeIMoYkzWzO905S
3OAxOxMxcYW3ZTd837WXC04odzlfrYZKNMSrx/fKp4YKcw8vuApExEgwEj1092Ef
HqfxBFI+LAZxc2DLwNRM9JyEZeEO8EOVv1pwz3Wbx3QZHTSUIzfa5NhdI+7mNv1I
5xGV4mAHcTRCC57C1JDeoO5ABXpSrnQD/8A9LajCKQFMTHVn58nhDl7LWPAabq0q
lVipYjqLxqes3c1i0uktTHyeH8R6uuC53VYu1wvMPXR5IolyULYeB1DaCeF1nZzU
TesmNxUZBDOPg1kE0WFaqHi958b2Fqn1ryLWD9pLqwnhTQyIpEAzJnXUxcdzrr7v
xrvs51TlYAjRZwzj5KUil7IbvTNYQP8PJlZw1JK9l/vmoyr4LSPBKuKU3UUUo0rT
yZRo97ZSo2hGoigSkuRFrUWBm7K9m5uukbJA5qpuatD4CNByCJ7Wp6GLwq/LYePw
Vy4IBKicLKVPzikoJUMTcdFQtTKX2e6HtpCXa3OKWyTqwZPsEjSX0yZ9BJK4K5m+
GbNGYVQhi043p2Oh8XTxgEKDX/a3SZ9or2tWBZKl+UY=
`protect END_PROTECTED
