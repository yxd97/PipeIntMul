`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lgz2Uc2XUmi5zSL5gbyRmZVuceGQk3QGzs5O567gFPulHOkaUW3wWAx43xRH5fN/
0G6xUlAYUIAQ9ZQxa+eBao36Koi+UMR58DLFqG3ngRickwS4poczvGi93zvPQLTa
E8uvSGh3DpvRM5M3LFzMB5QZDwmcqvccbFlXnjRgg5+0VEikwDZKYqAlAo7pXhLn
dIPuiEUrMjJoANBVgadAD01+umM9QGLBwCosP7HBlSqTp+EKglIhszapJpbqZxMH
vR+Uki5HqmFNGwkwRcBrCXn2umgo9rJI6WtCj5EcSVOOegPLOUS+aPsSdo0eJ4Cg
RwIL9vD+3eylCI04n8LiCdt+mpu+9ylUCbFeO8lXFh4sn2P8cKieYKUCNzjRYnG9
qkrxtXmPKnHKR7SUA/edYcMHijYClJlYKwNLbcCcPH3uTppxahGU3bHxlV2LklzI
w0WXxxLku2UObQOW7ecx4eGhDCi1oGtK54W+kbTVmaGAjJ3Nuo9UZIvpYFas5tzR
sl0x0uI+QhrlPemGFxZfF8mxGm/sRER8tXmyMWhTTJBX8Cq30LfcirA9W6RkHIZW
fF4x7R+dvhDcUAK5j6u8UssJ9r2eBrqMhOItIhg/IXANA7Rd7Dz/uu0cVK1k7Tq4
ulBVWgDkXLU1YpL6hiwVtz08cajAf8NomFjKyWLJfSIXZ7HtovdpZgcHO7xNLEqw
8pyik1HlqlT1vkS5MIeOJz7+hBFLPEGPz4rO9t7nR9nN2CqlTqTMJG2TIgyThP2f
wbufmqkUruunK9WkuktEiAsfHR52l49+sdr08kfPOdUiQ/zMpq2Qk7n4FhM7rT6q
CO2Ngja+t8D4iPZQ8QL+qNw0x0kqXCU5LZprK3JunhWly3K6TVOYYYm/CNJ+RWzH
OQZFPUWCVSnz66ospqaivlwOshbJEr1D9Vsqmu2sBISy9no8rvsIpMOUEzRFgpcm
YzRKtRrQW1sNF64MuKRfoOSAh971ME/G1RHGtnhJjZbPhHpD5WvXJskQON7+8oyA
HwhRhU9eW587wkngoxsAsOWGHGf7aj+YWZ5GeMOi8WP9Y4tUHEVWlaLzqNnx1t30
t1Q3bUly0dW9TJk0bXfo8q5Ae8dNs2B3+2cA1F6S42Qy4WyMab8KbFj4UHE0xx4c
T6+AHNMHIIe+pUHEhWZfBqW3iH1SD1/PYGnGpHUMDiPcMm4ryx+oQwf2SoR848G4
jPBkcAY5HRA5aokSncVsuCXzhmeUL507T41kSbIRTBnnRIsgruNGhcnb4hOup9Tm
EvWWHLb1M5WHrD5O8nowu7gCZqPLKVVMkTDm6B7aBNIZw/6d3WPJLAdiMWCdVSJA
bVrFWW8sGCpEDczk5y3HND1WlAuW3ZDbnobIgaonPjTmbyE43LqwRS5FsxgVBtOw
655/iFqRG7IAKWpSFOovBeUEejwlOwfsRhgRGqiix/bCmVMEnivn0kddKcszixwx
M0BXwnPMY2atLQ1PJ1IOGuWCI/+yXm0fxEnc9PfcOZUVMF9QWBGbz29dwutgdRkX
K3lV4/IEMMfop/TGr+c5scLvkh87a5s7X+HG1MOdkGIW9geP+BdYh+r3bdKJ6h1m
k2icOf0J3WF71s8GT6erCpLhpRKMeUtN9mFxUnie3VE11Mv+xFHFyJYA4/46Lske
KkgF8N/5kLbTu3zBudQhDO10gtJrEDE82b8WLorfLPcW3aLcBRNOXTJCseIxzlOc
6uHEL2TqHKKdLVPX0ohIkGKWabyfGbVyb+GTE9tgvJBWJNtT1BJBbwfqWQeTrtd9
W9HBNnCBy2axN+vrqSbBGSTf/5uPNOpeXiEngoTmaKNLdGDMadQAqrgD3coa9n/Z
I7rPxIuCaipM8do45+9rOyAOTeU32r9watyl8wi9eLvpfm8XN02+mLruouHvZjZT
VakaFvplrt9GHnGlQ3rQ4xfHI8J4jMk8CQIYmIgEQXhTQzQ9bX/0qCTrj4BuEAiI
Mr0mfIytvL3/HN6skhjz0oSFnoARVTQaWWfiD9ED+zCeSQbw9nZzGgHQVU8i5D+L
zeK8tPVW90NX9r0ONz5cYqVJKG28ATP6cN2usqFpWac/vxGT0kHsMWlcBhF9JYhk
6l/UTq6YF9H7c47sPgBuqR3vNliHJx/BuLMZmNOzs/oh45u7nEitq5ieltPK0PqH
MMX7iRWi0u5RGKFyiVGmJxIc7TZhLGmsai0rIk9tdiYjx0ktPxztBm2NIzqeleRs
C3DSmrKCjRVwhAwtLxrSOIlFTmylvTpkscklfMHH6ryXgsPYm7ZZ+caqfkrR1gQF
Ss/NK9NaQyy3FbTivJzG9DUdPmI2qI3N91DAyg3ebpFYZDRAS7BPMJ8xW6nddXJ7
lPbiOVplukSAlPijzOvmYlQyjvpit5lSyZ69bF5BrSSnn9Izw8w4K6EGpGLG7lEk
0fagoi/ehAmFM6TIU/5zLRDnvZfAcS4KG3lWRJgbBNHGnO3C5bNH32RJ/5mcda4U
1quKEPqEquCTBe0QRAiW7QbCcWb7wjjUelYYzrmMDf2IYqr/EsSeAQe1qPMyOsS2
zCze/P2HRy/ZWCvy55Uh0v22HCukUa17GOX9JdZ+cs4gGbk6PkbgdRcJVmbUtqk0
5S2QVj2d85edRhNqNTUtiIl+yhSNjWjpzSp4mlSOSLyGnahWP78HqANP1lGH3ISD
r/gjycAz243LmubwYJwqNI65iaJRJlAj/lxp4MhutF7CXQ2AQzxnC4CQFVUCYeu5
8S372Mm36rJQ01MSitjnrYrn0DrrAzJYVXwOybCJ9NfraaHIFjhIBEEX4imKlr7V
tDyD4hMq+UVg8lMpTqDEKTHqcQIqmPDUkMEFRGBwDPNS9EphDKJ8znnCQBepAkfL
HL4ix2D668fdtpej2ta/kUClCgC2WSfvSIOXVmx/x4Msmby+vW65WBX2PkbDWbfV
MI6VNUzZ96Z3UYMsDfivkXMr8sKPW4vCVhzwM6FOucyMaIYx0ogKYZUG/kcJ6tFE
ZlxKt8MAf3iseN0pveHiX2xO4nnK3pA1gbMORcjSpGnQwMDhm+N3HsnL/sEFGQv0
R8RbHEOI2e1095vsyhLIAOhO8fMcrDvpWUGWt97P0NTSWAZ1sKOIRwgPSIveaWKl
hpOZIOYrr1xfwAyHo65CXD23gDH9ZdalCIn/FUQfOGZnR1q0FYnMB2bNP1SC789D
IM6As2imnDIV224olsEpi9FzcJE1Q3EJVGEZ+esQ4cZJveVvu28hJJ44nzecYAEx
N5BHVCnY2OhWs7dr9UdSjOV0vlmjCEvIut3zlDVSrc7dvtIyenbx+JAs4/5pzhV0
9jR41H/mci/we9JzCDBRDkDV8EmczOtaUKk8WBMPJgK9Y8IWlX4vIHquoiRJQm+L
9jtWxPo1Rk21u0Tu6+PTmtGJczNhy/Bb/75ITlU1YcIaZLzIJZYXuAm83hBR1N1N
vF+piRA+PudZ+v2DeBpT/ti44jU4SH4jAJnmD7BFw83ProbbIttG3YR0/b89jnKK
Pq1jr0Xg6LNHPh85Q2Hpygv4xEhXifhavtc6S+BImQJAHKGd6tAV30d8wqAjFjX3
c0CjyQClVafCzygvzW++K2lgfqy7hItzMkI6d3NgpLmO5Hob9Uq+dER2eQT7R2cB
wFEgRhHpEox7f7HxFzl6KqE1uP5u7mdnK3u8dudoq5bDne/KfUdvJlGpFfEfZQpC
Or1+MXnQvGR3M374Z7QByyrvyY+Jsb17LK3Zb/YmADtw/Q4BShxTpQSlLAeyJD2S
N8My2+ciSHQHK+qbtuuAqE8FlnzTNwYJjWoDT2ZkA1MCMLjI0n3Vc8l4rPUUdBbB
6dqe2OjGEC6HgaqjaaeMu+3hja8Fsgf/oqnXZuhw79JWat3JEmgpKyrJljKOlIjd
6v6K/YzuxsZQeRi2q/IaG8cnHK96uT1ZrRw/QitpDZRaSMsbHrBB9naqRIflEzaJ
RL2fzwL2vVqljLnyawTj0t+cmGzDVGcu4doToKwBmDvzYz1CGPpVVljJ0tV55vcn
NEgKVdW3Pz/KtZ5ONBA3gDqHn74SJpSyA9AH1Gpw3x7KJhFkk1K6/iJq0K/tPtFQ
OiRqk6cX0DgugAPShdszpw4yKHVTAf/s38jfECZi5xTtpFETUTPqM/kEDeTrRj2b
Ym6lPVUI6Ti8kC0FSGvuOhof1SYy71+AwEbHZlV6jdME8dgRLAtOXbyGhbLR/jDq
O+ik3aRvTwSOhxQL9ZSi38qOwjc4GFbgRCLxnFuW+r+3vwWNhVs8il0dWv0vfbw9
w0E/NYyzvo+lTY2agYk4t7zQ4gqjTCLTJB80U2eMRst8vb8+NTYye6vCyITdI8RV
9zdbVlZcpSPuOMGHBh6Gx1G0gO10zfiwFozWh+QEC4kOJ5bm5nQV2y4H+aKzxeIw
8g/UmSRmgf6Z7BA8V1eYGSs2iZ3l1fh8IpnquZyBpV5HEyZYbrZWPGNS2641pCci
pu4AySLyGGfF+QW9xLYwIFxvjA0Lt3saHYey/1gZssyBST/ffbp1Rcs2Mb/wh9rK
DkRcfh1Vz/7BflEjYdvCaPZbrShrmADNMIqMdIM+mBfS249JgoTT8qqU3uxvfuEY
obUeSuOdjwNqcoMFJQWLirzvy6zHcHX4jq6Yd6HIekuYtIvRovQXwDaZglFGJXen
TB08PZrqSk1TSNCt0uaSGrf15VfznUufwkjooHYBme9IgVBKp7rbinPlgPaAwINz
1ig1l3TiehK3vIbcPDLZLrEb7LjVR/0CfuIC3MgbQO0M74vYjMYAoQHjfEdHZCgu
ATh1sCoiC2I1Nfx63XAeKfPhQmiBHbR2bjKa4z9Um4DgeqOtMsVRSlni2ooJ8RTg
txPrcQNzczTMclz1Jsz9y2nQyE5LX8La7dzPEHaUjLfqH5/oykHGkNwGcQKTq6dw
sZbM0Jmra5DbUsnKxOzhuXkVOupG9vJMy4W+unkkg/lxGJaQnMGTCS7Nkzsj8M+n
9ivrGLUhC14g5x920HC577oPCIDBg/Eoj4Px6f0XZhey+x4ll+Qx8GaNWYNpBvz0
3VeEkJhuHC7uBdysouhTZPMuY6MdxtyU7X0v8D9xbJEnrZa86YXF/t2wzcv/sOQW
h2ITYkXochBTfvPblUajy8Q1Dr6p3w9cAyfm2NfV2JL/OjFjur9rEH+xYwqOW37q
5Use4hGTuHYTELCf7qgq/f2iXWOTtO6Pi7HUfIPA27pA2gyNQBZBofSBqrZX5xqm
fGwZPSeeDbusyXAr8c8ZZiFRwMrFfFCKTQVgoHCZopBBLDRoRzJdlSGjIoR8FgjK
ylMPnHYW/KkLxLDp6WjUrwSMEwRd/wENQDqr1iVLVbd6nrjys6E6zsaJyzz32jj6
TbyCXaBitVG0IEKlbjnOJKFpb/5CbswnZFHEO6lFnyhNMcCiXkM5jjYtiqqNFkIr
peXRe8loBXKpfDA9qhAn/UGZEAwivrRqpDNhcffx+yCk3t5+YFF7HTES/EfvH7Qq
glExUy4v6tH4Cjhr8Us7XN3WVvcCjHNbrYBLOQqcR4ENBzoVJfn4q5FStP6uDX8m
g0NFWBTtJdmfb0Vjv+dhNeKASzobkWg65Wo1N2s5t6CFlh30/vCEFk3rnpx1pclF
QJLLcs4Y20CuVIm4YsXfilMENF2Lll30ZDcFPvSNAST/Gom17SOthDKGb2NwK/RU
sil4rJaChMgAGpp4Pk53/pCOKeVGKbqVjk35ehDsfdmoDywb2aP3SQIaNEUOcto3
no8ZekBORGHwuDfxLv4gGt7CgbnyAyX/cA077KViNOAOi0dIK2kmhQHlOCaGIc5L
f/d0s4y2oI0zRq2LXf5Dqdbb6hdN6MSXer3gfpe8pbg9Cw8u4AD00u+cdwFkAIp3
dsnahTlYH6WE8Pv8XkXR8Pv+o64r0QN1rVj0rsMINkgqG5pMJ0yX+QxCneKwwUOk
MG7869ZscWBk+fqyvZMog5hi9bL9XANDSP/pqI40FWHlRjdnNrfw7EcnjEXDvrqN
CUHg3htLNgYw64+5KmTZrD8RmoW47Zffvv9L+kWsK1uKaktg9Hikpy8o6Jb8Qnto
z+O99XtysRvEVS4bDjFz1YUJ7CSYsU+a7xjy1Rx++5KYApEvxU2RQ2Wu80Q8lnXM
KNaVUz/ft5KVHjTTUHsk+WN/dAgFdNPLnR0HqFGFmvjqxmzRYfjWnPqTvkXk1isP
T4urAJU12uFnUnH9ExIXX3CwhRgDr+CTxDbrGyjagaG+1bvzneHen05QGLhPwppH
iLT6BCgysyySXOr703shFO1+BUrTNgKXYLd2qN52fumxBPM1/WrqcUCCcLsUna+v
Sj8uwtYArsM0ri3ty08eRQE84/eK7A66yJZA4qir5OY6jnczPMCcDnnWWItzVVCE
7Ejv06/8hSZ97ImNsWZel7+ke4GBfZEn+83gGqcG9J+6QKe7zuI8+r+emyqCYQak
N7TvteJTMEZirolzFJRLJSEEguBS/tqHhfEDIhM0o1tm6E2pCz8UezejhvlfqIt3
bzWhHPSmW9vfPXWgTd9H77iReh4B7nQA57pkf07pFkIDZnlv2qq6F6phZ9gaSJ4D
FVRR6jmx1RTVIL/UpZoxpibXZJDAhWWyYqZj09hV+tW2ZEvT6aKNpDrRi78J03c0
r5/k9Jh8hWiFQJztdAJUWEsl73MZBhZfSIJYJz4DVCYteo0JQkajx0QIczNlICbO
cl397MLcIBIIXztzS0GdXFE+YSkM09GgUXJhJlAoaHSG5vAFvMh24SQ1fSJ0qynn
soTt7XDZI80wcetkl+I8MkIkx5J845Mq4m/t4QndRqfLAAarix7O7L6DdYupdqse
7NiHzCOnae4TuGupI/x2V0zGeCrGLppNC+07bjH0tFhUZlh56cIzSBC5vt17tqRo
fKVIMgws/mQG6HWne6uuHzY8nAErdZFN9/UC6FmXVyNE4NGfjRUXbzqGRBKKdWOZ
pJTNOqR2q/uV6+J5F5OaUuKrb+k4pbFeaWMI/JJiYaZTQsRNwFdNewhp6xULo/Al
qmmpDZcEutrLImKBV04jbOLNyIehcGf9ELlBGQGbhCMFNL6LX0fOGwPu+ccWWRWF
INP55siDOWjaoVyQJq1Ov3jXXa0q3DswbegWLQUhYnUzicCbeZHlzKNli3Fwv/ve
7DDSOeCrUnvdyJwKqrFzYDAj+KiyWqxQW0JZcGATC/jlzlllGZ7XbSLjw3iL5FaU
tQT9cvh1gcnZk0PI5VFm0Mi4VH2dFEsM7CBhsa4w8mDz4EtZVyE47CWhTI2YynHs
WagyolBUPw4oCUcwH5k/+pZz4No/MYDZv9aek7QM/iIL7fkCiw0yUEiohDKMdwAy
oa27O1tKtw8SQ4j8jYRhSWGT6Y8+PYdjBBw/UkvUE8vcZHSJrghrLESa1aanaX2F
KxV71UHTreuz6U4S4WoKz6VGy82j1u/kvXwczSZ8oaQx1Tqn04tL/1pWfDy3T/A3
If2DshmQ9bIhbWE6myPbBV0bObAXx+uGja4xLCX9PqZ7fIxpj9E7J9APyuscSD0J
bOn08zJaSiJrb6HYrPRhOARB4s7sFI4IayR/pYLwPvbc/pNaSfhtUTsRaykfpXWL
P9+wYQB3/Ou0lbvuYzFG/Rf2MZs4SkzE1vq6sRqjjI4qm2iAC5++Uz5y4oOtOA2V
fWq2A7wy7fBXan96bdI7E+wln19tLKdX9pDKy2tvn15MaHvD9RWaZXpv+gBFqTZK
cSCriPSFimJqxGANGdpiZRct9wfjTQZ1uJJ7dKQGB2NCnFZaSth8Mp4w6cJzYRvB
pKd72WWXaZGFIv9buoTB6jynu6IXInNtazpZJinu2OmOs5xggQOsyfNc9bCSoJqI
zOusXK8WPgPXSTrCYX12ksd9/L6/soM/nmW/TqcssFfaGiA3B5n8UkAhM9n+UwxW
W0tdT6V6qizr6qJX1FKMVqerLZms+NaxoGebCt5DaHqxDwY2TQiseVHBaMLgEZhi
UH7bZyNYbe5TBDDoof6VToNs5InrudJlhuw/jUvHPUWYSjDMtU95lVbOZiA9J1pF
fjjz5eDTkwkNGKR6v0ptoKwr3Mzmk019MjDbHoQR9P1DEZLbyD4lYWSApH3AVopU
Gs1c99RARFaRmWQHahLdIdQ7SoyzgnjfFaQVTjmjs5x2W86Iwr+TP6LhCsWhpDWV
eoPcXPYiqEknu479OLdqm7yE7+yiAyYD3f8RtDgK5Xh26gy4qrEePkIrlP3FoewQ
UjNMnWmh6iZqF1qVF7TEGLncYTvUoaiK2CciUQPauz6ShcqrIP6tAdPNgdc+aqIM
97vg6DaUoo3lK/ZnBLKMWAJ1qdUD5tDZwm+i0tj0Zy+RDEmmifTSzmGwKVBkyPaA
ZsoVDzFqgv14z/mYBuRGfhpKmnnsxRDjb16/jJdyGnA03FlqrcbZ7ayUipbMrW7p
5rPAhjTZHkBia1GiirEn19e1TwvD+cMEddq+wY8ReD790tic3vAD4vtCaMeVnXWY
3p59UchZv4fC9GekfcGRO5GwgGWt5KyqX7AQwEcBC4yANGs+mYLGDRKOrRTWFG+g
IoASeV/W4n4hfygx0yNYsgPLxFSjfQedCj6JSACB31DxzclIs72CISS/V3b/95dj
87Uy5b48baQf62TWDpqNOiIpUIOCTxVJOwPx2gHi/vpZKgPp8aTDDPCS0e8X2JP9
KOqnXPYnmfnDKOKmXDaXv62cH5DJOr6WracI70X0QNLbcKsEVjamxRQdkTFEijYZ
oa1OLw5od5/CaGO11KmXInh/fgGIcPJcTOimpsNQFwX+hSaASpoofwcj5lRbn/Ho
ktiKdsGlLFAEVYJlTYiG72tqDP8zZZMXDF4Hf8Uza9SW/7UA44GsM4f4O+wZqjjf
gyDVOvmgXHZnv4EA5R6bhVi2QidMpMcyljoFY6GzOnUqNxf5WOhUgRqYqfRV28/T
NHUZzBGt3S5qx9tgkVAYCdY5s5oiIbCrUcqeebSCkLnne+AKP2smSITeTDk7vzk6
HtP1Hq7qeFZeEaxh5zFlq7POWKi665iZAqbJ5cNMuQBSzntJgn4+GiJVXxk30DGs
M0nhANotO41GAn0azS/6Wqjl73aEyXThVeOGaQvvyrtUkjQ9A55qu4E29M901MMQ
`protect END_PROTECTED
