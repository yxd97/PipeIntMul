`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nw2nDQkNzqmo5xYa6xX3rwsuOMKmAA9Lv3aGx3Q3S5HtsgE+8lbsDYB28yc9KOLd
fdo7QLVp6IOgUnwoDnCfZ8uVt+Dg9YuY6pEXu/GqlSMB3Km7FwRKVxEANBy9b06B
vF5+GJg5wVaaws/XyeE+WvBuJS/glHO7GC4VKfaQYXYZdyITioAoaJ1044qV1jeD
njxD87jZnx79y+tC9/SD1RpEbm5VtGRsdGAoeWErIuyLlqjJmr0eauea2jNFA1tg
FEcopi5qWVD0Y44Zf5LXyogtwldLD/KlSl5A+U/+V4D2ZlJzSLuqp6zT3f+7NpZZ
s/IIqi5+WYjavT+T5EXfxhgPMJWxtjf9CeFmqniaRPz46lro2rRS68oAKv5TgBZy
9SFCV4cWQA16xNKGi0WIU4k6D01S7th3u++VwF0loLWXUhzqjC5w1eS4YJu4K6Vh
1hZuBd4ZeBqn74f7N5Y/eNK+WCD0/f9RIezYzYKmJ7Ykkoxy0xyspWzspBA78exs
8XbfpAt5le4phTHxnZEqhV+h9/NoTa9hJqEeowsiKYYSLyy4pQsiSFz4i4ZnCCx4
VlErlCpUfSzhIdm76iVbhSTZK61ssiwNqlAKZyK2ljaZ2SDFu3QxFQmgkdOHiyio
dDBJTgjA/UJQwLKyh6hPMsV2QI+ggO+aiCKj8OK3kUC9TkKJAc6YvZ5k//eygIN0
T77jYjTEeSQ1zl5jjnxuKg1JdM++Fzi/g4JBaHOv2wuKUWqdn48WMDpi37oCtoNU
MC5HP5LAdtoY1F0Bz7Fvgx5lA1Ei08q75yT48WiWB3Z+CDQHZ5FiJIv626WTBiK7
E5F2S6KYbcOE3pCCVQe16FaEQ+YcUkSYqfEx45DRb5t7koOTQq9YJndM871H6Jrc
zea+C59oeGTzpv9UA13BcfnlEyi7uiatDOUH9puKaZTQ1bZpg6bGgXbpgbLRxTak
pFXuxoj5edl9uF63K/ooXHbSAr4w37Gehr2fprHiW6FJJ1uvx3BXHpdCPoPlZr6E
MjmIWWtnjp1zlIc6qrRsEzqeuCq+KFrFa/wg5zaJHOU8Dz2h3m1XYfSOBysWQHHb
101Ri4b3Gn+Do/6YBs3Qr3PdSBw+JdXtNRgFaDxcdV8fD7XzKfOz6Wg/U5BVax8O
zA+xKNkt/Abn6VvrmleczU5IHfb5TlqcQnvfHkvBqS7d/RqR0mNTmqJqV0eS6SH2
4p5E0aCLzLeV9yLUrNSChfgckfYn6SKkkugTk5CGs8WYP8+k38LLxa04vHT7b2/q
rdOp3IUD0i3z8v0etXuod7Z2qeY9f2uNYNK3Apo0rzbAaGA6xKuQUDg/C4FxzJon
mwqTQUf0PxJrdyQyJ0/GHSX/OcMg13Wzh8F0OhYywzqb6Tv/m+t35p6ivpLWG8pF
0CP+K7VKTxxC6fWnz5jiMs6PKtJKQ9cI8l7mnhLRLp1k6XmsSjOAXeeTnPehP0bl
qQFXGBw0MZx8X6Oa2veMWD8mjPDzP++3WroyE5HaNBuorgX3H7O3pcu1AuNmsvUb
JZ4aNFfpH2lfjcEhtZTNlU+SE4NIFHMXKS5WppV+0BP+AedMoWUDcAqWQZm/n4LD
j75FyPnXodmnStwWS13ugjk+bJ5rEVnBp5S9GJ9NxM0bloll0BosjQ1wNS1kctX5
8kYP+c05iaqdnLrWHcJZ/aToX2ykNK/2M8rqIk9foRIObEODnpTpVwU9xLImqzC3
sDQE3iCYV0BT1H0qFnGnzmYfa8fJG71JCaoq0JHzBUY8Q+WXCkt12lqPge+ET4Nm
/9QTpzOcu7nsfUjyrYcJogIjcVJj107aYdbVlrSNp8POEgf3zz97YHMwXIXFj++c
7fTpiRXUD3hDbAAJHr4MKLVJrsovrfaAqXyma8Syu/ieoz8YFYHZHrKw2XZbNisn
k1z2I4X1vL+kM0xvxh6lnGRxbnSfhYX5puajV+HfiZavLywo2PvyToyC2Qygf1Xr
BAAnb1CnTBUnw/d7HvASQVbk7iJi32rymPGSvAcHfXaM4LZX8vBdrn5rIkQ1UVkA
zD1ZLkZo8NPpzMpPLMVySacJ4DouooWphJsNqk/w3yQkoiW+Engs7PJAVZ5bBXtJ
sqg02E5skWCh214yPkrWxIkO0M//DRUXHpBMVysk6uFWG9tTaHWt8xTMYkpmRzmg
k5EoUI20i43tOovzR1Y6htzENwN6hP7JbrUG1nz9WusL64usaRtAE815YZwHqEaE
cSmLGaTs0S6TUKaEGSijj9WbnulE/i+gvnPNxDdV3/OX9mF76ATJQme9uqVXp4hW
YDlrbD1FKk8f1EhUJ7eDni9jyZjCvJLatbcneOti5Fg5euuIsOnscT26d+eEwVmS
kuGFxNzcifcnEPR66qF96hbm6kcXXRfVwkiBxG/56EPP98MJLdVgIbJtKtmGcRwV
ve7wn4YwrKKVioJT5BYC/ccy4dsesFaSK7vSLB7gYai8jSa9BzJwZas2GIqmZ+tu
Ua2x1mxdV/TG0V1VtZSSRxOWo9lpgGKoup0xfoH/zUxTy2nckpR+ugS45l2XKiZf
5fjMsgZAttxHdFLJx6ye1IYGrR5ktvusX0oxWG/8/8NOmxW9szYHs9QL5dU1Yyvn
92PoVbELe/rcV12xeOpekj5uFYjxdhPuHAVlzXg9JWTJpP9vt4JEzfRCS8rVSCvb
Os/sh6M5jK33jjA1zXOf7Rud4VrSfASFABaSQRue8y1VDZXytKyjS4q1Zf3amVbN
YCmXGS+8m4HKYdZSP6g+Zyx5n61lZj4IURH9ibSdEkjKuqNXMxSNw8F5nG9rWKoS
QgINjz5B0HG4c3uoUTPkclyOLn8cWnSw/btnWRty5zUkspHqGZ0eqXhuKmJUrg1x
oN92TktX9kkE/T7o+gxZxBVp1BXKKdnzMZ1A4+ZLxzbwdSEqeGDiM9DSNtu1Q+eB
gDCs/ue6yMof7dUnySeueI39KtjspsMRjS+dpql+C3lb0AHdDk/nSdYSOzPr1CEC
5oLWPJ0NYfSGgsIbCuzae6SODzQK5dOp4ii6TCAglnCFSmF84xWThH7PPXg+ldfN
tKmZxUDgTBVrWJLX124zvsephsObyWIoKYgBLiVQbRO3uSQtd7frwjTqORso5PNV
cU5/MtALliqUgdFq6CxFQqtsppV8iZxgz9TmiMo4Tbkl182CSdPCNhRVySXBGA7M
7gORqtY8YC3movwtiWlTl3+Jxati9Y8qMrwTqqJxnWkimacE9KJb6unXLCMz2nWx
L5Ux/9L4CCtNrYt0SHfCR2MSGf/ao41Lj04RQzxPX5CABIK8DNMtRS1wju3cbssV
OrPTEroPsNSck3tSn8K1wfY7SfHM7+wJjzNxC8ufJiePF2Xh1dfR37C3WrDJgWre
n12I9A8ZqKyckvdhVEZEwTy3C9VPAlp3g6DlGqpGEKikqF7Q3sWK5xHOoYtnjkS7
FbYJ23j3sf4fq35r3E7IL0hLqYHJaykEtUdSnF7r3tuTiZbLc5lETi9lsHVSTNSU
347Zo7tnLzWccBZcSKkb6r19CoPT8XNPTigJspIzY2/tkpS0cNIFrSA+BijvAJDv
cvVlCNz/YY0QeGM0LVrltiroad7fQtNPw0cFKNOU5vSeoy97v/4ODuuaOmceFFxN
`protect END_PROTECTED
