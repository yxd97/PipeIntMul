`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r067n1YZHb44Co255CXOxyR+a5OtGqn+z57CVGkmd8/Fdpj4Xk3LcLw6j8NoG5bF
AtwaW5J2BX6uGSdbnVfUUKpR4qLS6zrq3cBPwRu5+onCsTjU+hsfHFfzr9GAplZO
gwRqDrawnx9An6aj3TUqdNzOmEiFQRdVAfn8XLW+w3zTdIPNwSh9lle6WFSypH2C
osciKQ4jX6XuQkQPgyKnWUjSfhnjVcWTrr1ZC+ZR8H1/0N+yFh7wb7ykifyhvK79
NyQhFaSVXUhYbUOSf/nn2Pbct3Y8Tc5wfwDyZzS8k+ywDEfGfOCG6hrbpCwXizJ2
+TLJgRasjn06YiYaPAPs5Q==
`protect END_PROTECTED
