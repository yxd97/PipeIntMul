`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/up03ngoiKE3SrcjliLyL3G2TLbH94cy7mJAWFJ6aPzhNrSEnejqkBYZvYC+ukL5
47JECXtSWWCB6dFSh1knRYAu7F7Rnc/JYbh2yf6GLkRaCuG1g1Zk1r8tOyNXl27T
y04DX/oyYsn2MHA+0NMFKETfRkiq0kudAG51v4ufp+DHYs5cyByv6gf8EnVugM/E
QY+IYPF2hgZje5yur97+O4Y5dibPJ+NyRRe3hFy8MC9tvZG/7AU6YyIHMO+Bmeh0
dvflY75FKL89GYlVTHoUXA==
`protect END_PROTECTED
