`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBC5FnRn+Lb2YcTOXfW5Lft/ZeOsEeSM8BNOjicGmgnkBVnok/jfk//tmXjiHMiJ
A/6wiWtn6Zbn2+mcgaooHVBPePvRoH4d6ByT5c1NOhRdDUqbhCouWD7gOpQaAz7m
u10MzNYjYxM1AJztlvZOrEY9dE/50piletlmxH79oSYlTRtZinQRU771fU1p5hQJ
jez7tL6KjbqQY7NMBvfAujZt6wZkvgu4kjbEOi0PNsGGMzTzzENnhR1KhRNnpkE7
y6eV35NSMfNV+8EP5GRTPzCQmiuN0nxi6tuF5I6mbMdzAdfLxn2bptrlMD+TLPuU
AHIbNea0n3Xy+mIRiTul+nxS6x6J33z0yxAUg/nvL5JVKnHJ3j+cLwfTRZXlFeXO
XtwccJhHuZPrLk7R/TBa5ccmDLB/RQpZ+5xGYQYVn4ggJW0uALlEpd+txKHwVOjM
ER5KwNQysWWv+qtI3jdcQI/N3/DVN+vRNQj1RiF6J3Xie5SJV697NO58EwqMsEgB
S52gcqHuuIXEzqn8+mYxQXyLshQQIehDYjApgwuTfzXCXI355sWxPpzyUMJZC6HT
FVK10BHofbj9jacUPQW+tBr3J1cQV4G1MZV4/XjP/2aicxJDKIkFKPKNwk4umLpH
EDivPXSUvAP1VDQhzaBTR3mYHTuIMFbYQbGXZlwQ2Fq/teuqX4TXejc6Zo0u1V6y
wlyt+Xwqo07A2VgWvcMGa9m76wMxSAObJ64pbyg0liqHD2AjX7DMYjSGBXS1O3wa
6UXu0zTU60ztpezbkLBhG1WUuJk4lbKYI/uwpyblmuNgJNhUN4Wn+nHH9DVL58jc
PTPmsgTeHh6BA0TS3WKJ5qCNIf6L3kHePjW3b3ELsZFILQPfx/iBuz/p37bC9WWi
hpRx0oxaMFVWVfVanwiOULok4PzZKEJepovqZx+hPxTWxMeTf2O7KYk0zOfcXHK+
le9lnBBpUKQ10FG7TcNYNTzHAC0B3Xw+U1yKH95xjmbCEOjpDqnv0sjGzqUqJZ5q
Hl4O6QViF956kdsfw9yvw8EPTq1bsZjqxCoKrttnp4OiHhq4bzmkXhBx83KP6X3S
g6gRzTZYlRr13+iRb+tqgTbZ2gMfl5zklshAOGdSeLOU+GnZ2k9JZFdzAAJyRny3
/XmRAmJS+6DTAepXRruBbN0r9LXdjspLSFVZletAzVUvlRl2qaMyUs7/+vXtuABV
HubOFxrUqGjffFMKQXq13hxb9hvCN1XBSo4NeE1tcEniZRMYTcvwA4zoMHebBcD7
eQ/PIVNZrOAn0qETh+hthpjKxoPx3ASaI1dHF7K8mtfSp7bkQcnTcYU/355sb/tM
K9dA5laYZDSrxlD82VMpl6G2jw+aLLWuYbi6c+Kxgv6Z9ZgSQiiMoXJEnNu6a6zI
TSMSsvUoNwwMoC+JrY8J0PWj/lHfHDHU5mF2SHlLmoEcK5CePEmCR95axbcGBKh+
Mu2anCdaR2UiPtNj9P3tFdWhE9BJQZoLNaIY8/7aGn07Xl7lzBU7qmHg7S2o1zD1
O1gCMO+kJ8QnQVX4McFVKYMckM2Z5qAlHrzN72revj4=
`protect END_PROTECTED
