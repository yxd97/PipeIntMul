`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h78ZHDGwpHcd6eKLQ9ChFFSgs4KwrSWhM7y4Ommt1DsJxb92mEJo/JvESRzCDLSN
6ZHhgu5XojjgvCYM5DWFahVppEkIcuyawu8PYHrxiZ1a1n4UeAXjwwdU66CWe3in
B/hJElTCF/7QKniYlGbCvmAMwKms2fJKPeBYwK7GUDxErfX8mAICJhtRlkTzg2WC
0IhFyhVFfs2qwOgpVe8DsFweI2PV9Fosc3Zr81tj4b/jfMGjEDGVbUXul5y3w6fU
tYVaA9CH3GaIM66WNf2q4az42ZPpQ9hoIqYR8ZbwQj+TGjO6bvUKYJQJb9UuqOrN
3TYJocVoeko7P3EJf5NeckoBolYPD9Gq8m2vpRLoqGmve59eeZXaEnMnCV52Zm5C
UffLiuiQ26Y7zebEK2QnlOoEe1FvRVpH5HujQrHvmMiRvY+HAqyur6y4kSQ2N3HJ
Sf6NTTZ00RvSN4IhW4nQf85riS8BvMeYl1mG8S1TZfthT8MLD94djmA9CVKh+hd8
yrNs13ULPe8nywoqFQg6d7+OsLM8CR6oahTnGaX87PppzCudUpKT1ajWl2+QMpf9
JSvYOIyEMM2V6D2MdwrATppwOZaMA3oJYVfe6vDeI1KecujGj5CCzRBSwLhRnQrO
8victF5yvuCbWUE4bSgAMFHzaoxfSGldSIiKhINIx0aupXhoqka3FupRXzZraP6L
FWyh4eRpWNbS1xVVKUe0OoC4ebPEL6Mv64bOD8gGWnnZ7DtFAbMDNaCl3JIBN5oX
FAoMiz7g1p7uAF6nJRxUVVQeagsfXEGe6wXEIOACOwYKgcYkQOhrGqz2TxwHmrbq
aqTnEmuHl9LGEQ6Vj4+kJuxxl1vljbTFue0H1ay7XFSRRWxiK7l2vIHqpydKASgU
ilQIRN76crpFUxQwLBq66AkoHfkFyYpGCilj93f4h/T40st1X1PLaRdP1xwL6D4T
8FwUW08+h83XjuVB/cBcX3XK+XbL7NRuYoYawKcqmd0WHS9jOeuHAkN7SZRKDdtM
YbnGrO/Ffllz3Wq1gXbYCCnCWdhlr7MRQFcRU6IhiH5G5QZAT634wXbIFAm1uFqn
IF3v4fwajcn31B2o8QTKBXiiHeA0hZcji7Fp058giXFivG0YgW66QUsUksY6A5uJ
j0QGKg4EONmMLOFI6OGGqeZCIn6ij5wLsLH/5chXrfDIxhau8ZeNzfjjUi6U6qQP
lk/R2l0h/oQD86Qx244WX+0YN1YlxG22q5BUQMvTjKht6jzEXCv6JmjJJIUHBqhI
`protect END_PROTECTED
