`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zm8soURiE+KKZvtQf7I1XfSq2LLOAMf+tg87xQ6M7n1WAn8XRQsbT14gcv6IUnNr
B+5Z7q3jm/8ERy/MDMp6cex5NYmTceO6JnUOBQpl3TuI9YxaCauFprqxkWwr6bUE
7l/2M7UVhzGMUrbRrtIBS5EeZbOIcxG4q8PPS0bI/YAXv7Gd7lVpBiA+0ASkddtZ
eE2jH8uyI/VhfGLVgmHLbAxPOIiJc+IPwKnC+T2Nv1AJy8Wx5pfVqEZR81xYTXfi
uNAc37Emg/vvNbhyoLFR4rqQoV6gOPVtlWaPkYnYrKzSMe+Hec2b7ElWSB03sS5B
74JTGSXIZTzj+7jkymo7KI79WfkHs/uz1w6S4QIXoyXfddH54js1iKUP/9YfRSDr
+4yRKp53A31jCWda9dYHmuVBToCGQnHMiSEt7eCCaWpt5/YzWx2d4u07Xxt+z+lO
yWQJ9mWgf2bzCa/0yxbGGA727pQJ2o8nOnfgRSMSQoTB+djAf57ctiUbR4AClkqc
NiQOJP/fuOkJ/9iVUgQA9znZzcl/dJFwGCXWb+fu7Ijcv7tq1X616KjsTKBrM0VP
1Hi5Va+exshrbd/SiHfteDnxcK1GszOZZQ6XFhAxd7Xm4ArR2sgvTyN8quENleiO
2MYNlrMvN63i7G8PWPCkn4x/tec75DRIMbDl3VAORuW4GeJiAenIQasAXbnWv8Iv
pqIx+jGo8FW6vWzJG+jRRtQP47W1GTRZiELvX8qz4a+AH35qWQOMgtdihp3xg8+t
RAs1sRzfQKRhW6cZbiqCHikxjMdYHGf7XfN3nkJQlwZ1R8SQvWT4SSe+iMf3WfqC
abL2LEvETg5t/m7K8pDtLJIr90g2WaZP4+JFYMPM5X/9SL4/xS2XZ7RnJ9QV8gvI
PKNzhwNPvxcdqyGylG3JDJTKEo5XagTdaKtPikcZ0W49L8go7OLXZMhUTfvR9FUE
2XL6E2xOUKSlMPcLKDEz3Hrpf2NunJtD3SHeaVxYzshF7AUs4+u4tZbuhHb/0szJ
s4PQ/9t0SlhZyz3dqWN6tBb+nloLLDO/fUHac/PCxfaLNsng+dhUHuZ1qdDB5s4O
ZeQX6V7hC7MTRvCfGc2z1nSo8M4+y9L/Slmd4As+YbcnwUsNasd+oCctIBRLdJGR
MKpmlnWKBpj+74/87oX8/FFZ93Ah/OEGczPM/3LAaeQSr4ET1uP5tegFSqNAvZ+l
Bp3NFAaC4s4QrmAv6v3Vwp+Qnk8ObKxZhA8+0Wy0iTC6hXSGY86BO6UpOfNpcYrE
WO/c9nOpVBw95yx/MNjfeRGIUaI9r8TK7ENfJvYIAvodTlq+MesQkt1Ko1V6Kbqq
DX+ONG7xFazQdjWfr/flkdltllmkUN3ZHqenwEdXZfUAZhEwv0AxnUcyhrPU5Awg
OT7SIgTga869Cl4fyqWlVb4jnDi5pBonSjR5ty0fJvzYUwAqf0/gDPEFpHoE6Pzs
hzXvI9uFKnVm6mxt9LjyM579W4g5oR12goCyu90a/1GP0fVBtgAWityskaJL3PAt
4Sx5qLJPBj0Mx19mFHdueVDhiqrlPR12nhH0eHvp8MiKofmjbw7KrYRCg1rAFPkB
4I3Ume/2FyKCtERrwZXlcXVBLvNfFh3qt8SlUgqEokbxUrRCUeUAzxRDQerFewcQ
Mm4SUI8Zu5loLgRmFUl9tgoW+yIWr0friAMs/6zfJ0DMyygBo0A8TgCCkfFmqAsm
ZCxJxwOLWwR8ClfxH8vTfi8olN7BMrkATtQNcA0IsTytdfXizV3ns1W1KnIy7drI
11ylFFCI8O6dfhSjzQU27WvbUzypjdBHCC1J4i2dg4JOlyy6kvVo42VNLLK8Y6Q6
IA/E4M/DWJ6DL/7hraedNrRWjUekiaVpbCw9VjwWjvStSBwF26YzxzvR8GjjkhsB
u0NsZl6JFjcwMiAdromggdNF8yc9/8zbXcOIqe3AS2FSAB4Q+TyyYZZwZrZ9X+0i
PSE7UD9i3dHXmeA8J7xvt6RE3rE29zhULdPhM3Fg/6Mt+P7/EnLJuIWxACbByoU9
bV+ezxbc8CjbvH5CNc552qwpiNxPP7hLTYD0PaTn/DA1kCqumQ2D0Pi+hRBKvKPb
RzeUBoB3kCTscHf7rgx2ixNTz1XC8cVo/rYkaQMF/GwJh3UbqQIJkACeIZxdGwKO
4vSElLS+TUQ/bAc2QfIEl+BHBG4hYv6ZLAcVrLrmpK6orGxpDGQAhFl1Z+7FFNim
eI9Jiw06Z8eVJUV6fmrHTm2cyPvtmjBBoMYayCguFvG4aOlXPic3X8nU1gZ+1uEU
v2ewYaOjs46KoN5Nt/9e6LQhjf9TvfC7Gv+jpSrZCVsC8G4G7UunnUAsGCIn5HyJ
/3Gn7u0pkRF/3D9ejqRDCp7m9Rq/K+MCyEAueAoOdcUcfZEPCvcqkzIQ/pr76t+D
NiWAQJemITQBNCAZUwi4jaksDu884ihGPFISj0St+d7epVJfM7oMxO6tbfE/j8Rk
ew6zghNziP/EJmq6UR9X6KwVnvSGWIPGVQ9Qfz4CVJPmRspYP4QQ+Hp+AAWA8vqA
t/LhV78OE1evIT3YvRCNW2ZVXqmzqns0w/ez31BPek3YyfYCD7pWNda1Bf71qq5H
hYQuvqsEGLrCcAhBvw3NS3XD4UIKP24mTwOSKm1VIF0xtUpsA7Al46+0WAyX7X4o
9PAtrL1LZ2XMLDtyDjO+3UjsoSNx563BNWKTxWKFzlPX/mWMlR0WNY+Fp3VKdnIr
8kXK0UPZk2ZRfKqFhhgM4wdVNJeed8HozTiLbkPU9UGZb25j5QvOQne4mpFyvebT
Sgn94FEkcESeoVVGoCQwLq+oCGVxICcqGyPDEt1JuwXCcGKIEbCRkhE01bNllutc
RbUoZ8ycGO3wpv/eg3aqJ60ATSXdL9kuKcMP9/yo9lOAoE3RXxBBb0i4sAbn02S8
c2Yjfi1zErScQB439CeqYgxXUz/ZzYIh+dRThokHyB4=
`protect END_PROTECTED
