`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ImoGS/Qmp2DJAjB++x5KpV9AzEZ7ykOv2VUR+6GpEZJYmfT+GmJEsPmDm/fb4Qb0
FUrlSBTEEeHgxRzPd5kG7iOInMu8Xgd6VakuNljkeU7A08oDikIV1vt2zOVIwJ4u
v5UtDnkt9mp81xPIlub0i/72+QYPTS+bLZHNQoOpWGheNjK88B/m3pp6QoPw456q
1+/PQHZ4hIIKT+k3OqcnoL6rTCT+qAv9/GBo0IXuyLCSa352sDE2lf8639oinEmS
XKbLim4rDVHQQlyd+O3nYv86GSkHS71gkhyWm+6Ilpl8C2VNvfr/Yf1wptC20A83
EaFXHavOUqmhSg6ueHQHM6I/pP0WaSTp6ks2CD4P8SxS17vKyVsvkSuHXwvmF8V7
NKkCeL7uvSuRdyKjPP+gmpJz9u5icvBrc0vuppb9wmQne26SXQGYmuL3qY5+hlTQ
9eaz496dQFhwsmbra2xDDtD6p2JjFSdBpzkThOB+RGs1obL5889MjQAP6FcL0gvG
NT2fv6xvUAjd2cp9i9uU43NnDvERl/B86VIO7m5WBwnAYfmzDvFi5VvpcGG2HnER
dgKwDeKCedDFcAv/09Q5kqXS9z6uo3WEOOiQexj0EjE45xW7OLgmo2ZNzAQPwFW+
SwDdekY9mZksehXUHpAYZY2QruPjiWK5iyyJiVAHaPaBdlelvkqVlLUnwY0pAxkU
Jj/EMnjDeriCP/GuuQsUGcxB2Vl0a9+6hplJPjWflqwVgRItDgm1AW6HnnIusAt3
qjrUNh/icB1J6Q45oanbHubc+wpxY0/xpC4AUYfzaK34c2h92pAb8TqWo2k2/kds
rJRpmsQbjdO5VQ0VPMH+kgKzDTrJU+hpVfjZSvrA1+MR0XoEiWldySIP9/KT2DY3
NVOJkF/lO6gj3/LKjmDoWzHaWlBQDI6SEY+8j7cYSK08PbtbevfbolMXdCTgI9eB
DhriUuCwwM5BzCYz+vT41GI41CTZ748f/DVa7WQZMJSZ0d+39bu4iUYZPDxmbBlg
lOFTnUX8c3f44356cOOCw/2CG7xYU6kxA2B9rNBDzcws4CNkv7xNsuvf8yW3ppP8
/S4q6KyVsqEZIcPsCuyd6AryJbrIoumeQxd+4/HxVE0mm4tPVUmnWLSelOtbW7x/
Gcw6jacNXJAKVivy5d4QRJ7xd5wF7exIPshA36tmMg/kFfzakArAOYzKlwfm72cd
jqqDPzMzzYVE2+Im7Eov22hBsn6oFRP0djxog+uU150dKw0AFfAvsHZZp+hsr97h
TpIClT1etOJbg4ccgj51OWeeT6nls38m0Yfcushh36//oUNVbwYxRcwM8kLXaY17
koy8FFp7pR9BhgeOzuWoY4MygIbCndAZoDzSm7DEAFHvUbjDeqvWL6eUZiZ7U+1A
oalHU3nCH3VnsabRUW/jDCxg/nCsxZmUzlGNii+jfhbMKfkuR5xci1WGZWQsmJ6e
ouU75/l40b2rA6MGHQrY3+99aK+H7ki2ABbqljEKrKLry1UiLANEOS48bNL1vIN4
eyDEMjyTq0omMz+WnUWX5ST/Z8RyT6RT0S3ZnVWieOlkcLizZV1A4pGDwLuXTv23
ycyhL6m5Yeeq0nYeIcPFJFn0OC6FMJQYTy87iUwG0ixSYngM8d8j+HLsq8iWDB6Q
j3i2Y+9zronjVxLCDQxYyyqcUpvT6o909SfMDyTBEyornAzYERF8eWhd1kqDZHZr
iDqtJ/hOPtSnVkMZzhxy7Ek6gvwPgsA0qhLpasSQ4t3xPylD2lEpteaQf/+JLyw0
9/xlRPwf5AQPgLdtE6kjT+RUT2QMa3yGwl5wMMZ+yi3gphBOBKdOGRjXWS6WA9Z4
lD8LjRXbvAlg4Yd34JQpKt4S4nUvufAMmXnFkQP7eO2dUOKIsLHdRWPonmSfBy7C
aAO9UQ86rNHwvL9V6kqLnLZefRwWfp+LIoGXUL7AU17QQyFYH9hujtgBEbx4yHuN
i+nyZvJgtH1D6h85vqmvD0JLrIyMZO+DLWfBVvTGRl1eNhS6GAw6DOGAf+oyLmhK
3oNpUGDEdtlmTjmAd0N+9Yq6IA4cZxG1JN0FoH1VCPG49y4EVQgFmp5NLzl6Fhq5
geEcm0VQenrOFjg6lc8O6+hPupa3JmlziUB2BGBLcDVIzxt/Zcb0rtIpA6yuq7st
O/34Ekb4ZWAnr0Y1Wkt/+7DVOaA56KHDRGm5Jq2g+vJvUYrLzPihifdndfHszPVS
dRiCk6Qp/mTtLUyCjA9WN7reE3Y1QUOdgCrTjg+26CR2YDwmNbhGVugRhnYmQtiZ
uwzo91X6PVk9xX6i33XkzefBCJoZnsJhXbX5PGwnuRnq65cBZFUYzqDUJECvCBuN
xw3++lpe+YFUt3ryJNephKidFIXSSLruCuQoi7mxccw=
`protect END_PROTECTED
