`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+uDDLffn6W3dllU5vKu/AUGmLEDsTrx5yM5McLb14mYMLCqt/BGb34UC9u5mjjE
/7lvy7JgIYYxkvz+FBT0gY+j1j6JSFidWr/rVaQH2CyTJYWwtDr2CpzjD+LLeVPy
25QGLxgdkuhWYC+I6GGtdmNCDZ9+8JLnGXOTEUtHTxkoGkxGgyTPjq0iw+B5+Hjj
y/MkfCBCQaieyvG6zMB9eIog31G9FCvQ4GUr/Qxs53eP+qsWrzSTf0UfGhUqb/Id
t9a7GSu2wGqNTsvxFba5aAuMgOfTS4ek+S0iAheY4rqtlxW2FRxyBxLLM+m76RTD
VV5Mh4SdrcqSfHat8jP+pecsNqrFnX5Nt9ZOhsVITQtvxFd6QXkyy93xIrJFQ//Z
CkBze9mxUKEJNyOE7tY2vVneLwwtFNI1UiQzY8JwNFkzlO1ilspctXJM/CN8Xl6m
6pnpRfOjWCB5yQOlFNWIoS42ijSg0Evakg1/NSUEpwM=
`protect END_PROTECTED
