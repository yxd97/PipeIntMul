`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3a5PhKiLix1ybkV/MpVtZs4LJ0Nbf3I9f3dzTH6T3NbQB1mpzgD5GXS9a1ixc/aX
yu0RxnIVaBw2UAYGBWNNTv5xE+qDP/RY8cOu8Bep7AzslV6cRJS0NskcjO7bM97w
DV1bkK2nsk7CuL87mW8DG22g60426R67u6WuJ2uqBIyc8gCpO+2uN2MHdId3ldyX
rT/2K2A2LfdbcRoREDbXph39BfBv/Nk1OYfejQYWIePWRyG/AJeNkoVtlxolEs59
IhS/fCMckPRaMj8DRLoUbcQvFN34qg9l7Yhyh10+AmnEa1Qd4Pk31wPHOJi7Jpwn
a5kXJw+a7cNTqj2tgXZ16Kh/ypWh4zSqDStxxekarN0oh20bOj4XaUnsKTzAUNg0
U8DTg/rTaxpo0myKyp76BRXRSUWxSIIrsDGQcEP2weiS+rQA3aCsW9ypD59JX+Fn
ZMqnIvFraksKbK96NpsyIiB150Fh4jzLRSTUZLbdO0H8t2AxyHS8N/ObL+dtLkIw
v+bChrBvwW1lLUsBzm9OzATNGtYzTbRDteTAcTSXgiR4xdFejOcOEhj/GKRkrIhF
DWL8Ee9HBBquRr+646uJJbpcIHhW816vX9hzl1bpksJLk3mfW3UVxFf1KYcZi08p
VMPxujCyvHgX8+s/nrBEoshG8m1dq64nRA3NiQmCQFqjc+OXMN65RR5vYNOlB4DX
Dyj1Zv2kYDAfAvhmQsnurD0NCG8Y3rN8zR5n31EHZ5+y/trsMSDKWdNYDZ9Ftx66
km22r1tTjxyiIQE9tVvT+OnhYQ9lXSoj4kbCi2k/WoEsDUf9FjaBV9664oZc8Vo5
Esff1JKIoGa8i4MtSvMQBWRzLkgHig6Wiu4iz+t5FheXrxb8GxI5yM5hI2rU6Q7U
/7QWx5x4q26MZ/eB4R341w==
`protect END_PROTECTED
