`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fV3EX+IdFeUaursR206OBsVEzoOFlf8VV9XqMOHlwik8K4uxW7QrragW08LUlDED
yz5VDG2JFZSIQ9GC39GPpRm/jL4nbaL9znhIDmOT6BAGwmfX2GAxIQJdYPF8qQCs
Eft7D5xKmfVNVHkX6QDP4/Qs3ZuaBRzKEON1HGhcBBNNM+t70+Q3JbfREcPBo1rq
+oNN265zEsK/2Fu1cs6sOgCeQd4FiWGCplNP6vpdT+J2Q7Xq8o3e6hQjZ5Dc3ls3
0gN8glMD7JZK7nGW4vYmI+Z7A+x13tN1NykbPRVkdqzM1WLk93GGgLxwXSDVLilc
58wir8DMrIoertJvVKoREhN2xUeMgTp3FMOhUJJc1QdqRYnEubt4uJR9Cs8tsxXa
fhnJPV9ktBywpdI2HROXntSLugGlp87izbdI1rkqGuFrwgJFfqLG3NQuLVpVFD3B
B4Xt/bfIYljHPhPxVDto4narlFrDgw3tRroZDbAJG22jQc0GoE8ioGB6gYpuUNOh
Sx2ZVZLUQspZfY2g5/MpDanurtZ75wJsrCKn9g+TgwpCNYJ1A/P3DyMvgSYwpj/2
PFSRcBSD2HOw8p/+X55uNssBzDgd8BKOrGSKAN+yvsd4a2N3FLwT1sPQD3nZCNc4
mwgTqVn4vk5/4WWjNU0KK567RM8+ZMBzV4/Mk2NIUjnXKcrHWmDv/ypQkB5HXsov
6qdf6HmwK2TQYHEjD5GU51XYgJSVpqiDtG7qjda69tLVo8cEhOo8kaAdEmWZPYli
8/TRB05SM/9qdywwSnLU73oYTUIlKhOnXxHcdZn1R3vP5PVFVaczJ3EY9gFnHJhM
O6+w4/KEyNi+0DcPH6uHnthXN6JUqxI02UC26dWeCcV1HwpYOiSQi8HQyUNoi+FT
tl1GfS/hswzXSF0Sod1QV2/qLTF1G0To3UhgA3wDR7vNlayzOPSctDCO6yFah9Tb
T/+5Kza6E1D+XU2FJXVSSim4/xS9zymmCteJTtj17XWE7NDFG5fk222qqp/UeX8C
sbqQzlseIwmbwfohIABSzgA6LhLhp0w4wUPD4EuuwAW98bxlyeVngqBSJpgiCGls
PoT6lv1a2O6WZ8eh7Do9NAqAHwo4Gdj591+a8BwdPEWCejl7g9gmqHun4tOwvamQ
ErYT0qc7ti7WAxlxskf/svnUaw0R2oIODp5ZkmJcUsDqnbigJPlWRnYTJ+LzuYAY
2Bph3j4W71KgyfL7JeGXI8mJVZ/6M1Ovs/YfeJQ5IIKZpyh2fi9muWQuMjvvrcZk
wHlqPRn/ZZY1zVG1qVLhAF7oYdel4jRL0mn57fFNZs+yd47C5SoYUJVHyoRFEX7S
OO0dkTwqrFnHlSNIMlf6K81hiE5HSYEDE16wWJ0O5/pQlkMIQmlBPRziO7EZVcKI
oRO9SH1KcmeVzLibhky8m8uV6P6RW7B2f7A5aNExvxoJjiciwtCJiLbpINJsmiDn
uo43Hi+G1b8oRDIFPeUwMCOFzP4xV2RxfGgnGhhxs/2it0A6YhEdCtFGSP8YBmAm
kez8+tV7Fac9ZN76J70wCt+qvbEQhV1k6vQYfE/E2r6wsgwPSFIo+rar9oVIFjK7
8eE8BNBUrAgrki/JsmXqKGxTgxI7yFzZtwOV2b60mNJSH0aubEx/2ufw+P5bTDu7
TSlnTs+1dhUMsQB2ToTKIgCw9HCqtdsQc/y58QL4lVcDpAK19SBi91/LDNQoHMZk
GC9v+8lIeeBTtysH1xmlsYaWig9ypmal2Z3LdvrKd9wyrQ4tjCoSbWKVv3//R4Yd
zZFI0haL2/lYvqBZp7YFAjkbM2bv6EZvfiAGVEB79jTWovR+Z2FDR3XGTqaU8vgu
quDfpsVNxrQNc9v9vQiWE69aYXr1pTjsGpx6D2iTjYJfQAFtV2eKD+NJMg55V+iy
F8CiiYERxwhMUQ6d1OauRnHoY5tyNzgklRWAjPR5G1DB5Ws8VIzQ66lhxNPDZF/t
08YpsleTE8jD3S3sQlFyNYQWjtfAIr215OzMVqHEe0h9M93NTj6/DQJNTWHyaUj3
hE2qhYGSh4i5eWS5EWzYGh94cNCV71f4znmSE0NXPgE4/2wuJERknYJsbb7oZv2w
tOzQWoitPX/rBZtIJhdOZxDeOlUP0Zp4ebnttjmPQJwjfrMWJQ6VLnvTaGkPxqjf
GjPcP7tL3fpX27rqiIA7hY7zbaMKjeGdyrYORqWXnuR8bNO+TsG2m6cQ+vqP07Ou
yj2VeAz7Eppysq/MHIprwQ0rknbYcTchMReeOdpNsxtwYhHMXrVMpcBNwI3tAcAy
IFgIwqT4i2t5TO44elfj4BLHsGMu42KbQ6TVwrartAtFGsfhCw2oDFaXK+xq6YBM
pFa8PX0zCFm5c8SB9Tvvx9f67ANnxZVCt0kXpJ93oxMh4UGG8nRUjHR/c8oK0gt3
U1TbsL+nNRKtmef9cVgGh3wr1FylV7BEJ4y6qgd3dQdb6pyw6dURGfBSjzn/xmK6
qExmDJBXT6+oqqQ5ZN7t/pfiGfk81KD2YLpG9fZUXZFxOrgXsgwVR7pEOCILHJeo
DR0m4pVgI6giO5LG4sh5RKXYESXMUQf0ZbUVBsQa5k9khQH7Ll77bCpPIFqcD1S7
UEOD/Gv+XvlwLjBG/W4Ydpz+5nM/CFoz9XF1NMk5Vt5bVJa9TOYq4Ka+8QfKzqec
kiRNpKwKwFHSddiWgqlztEVYOb/W6xWbquqCjDXH7duV+Hzfl9CpEEb0LDE91B+g
hj+DaVLw35LcclWq8mcEWbMDJT0mrV2DNvKoif23SCb5iCfedW8zanJ9Zf36+HmE
Z8LA+NuIDUQ+wIOGfkKilE7apMUGaYecOSxWlHn/XaWju6Jal/UIlUoYff+2eGri
OTUvEFN/grwLtGcydC04uBBF69ThTgyOvTZxvn4doSWgsIs3IuH/3sdTuuDjmQyu
GiOT5wOPmTNBv+LQZV+zO2u1JyR1PlLgEizfIIUxhL+2bq87O0tTyB/QhaCmNkq2
088tDXXAj1CQAPW7c2+tMfqRL3yq2eksEUq9myfv9JtOtce1vRN9fHC/z2y2TMCg
iMZmMAiaFD2HYEEj7wyMkIwT1XD/m5mWzcmxhoQJQfSnnQUhjIsn/vKOSa7iK0Kk
nmEPW5MjdsCgXCrfRIqmji7ib5vcZTjKR17QmaAGYkVNTHr54CNm8y59MK52HlJ/
AqlsW6GOtClukBNygzJFyGvmm5AdhnjVcFWpveHRveQGtcfGWsMZ/FVQuhhQaWwZ
TT3K+DWu5Ru/MJwONgjdx5A9hARlQvwsbQM+3h3qgQPm+NunaST/8eKZk/p5AJ8O
74k6+HoSQdk1bVG8sAnnykz0gzYKyRNHAeoXk02P17kRcaWkBDhJGdFB2V5VUoUQ
FfUQuoVrBU3pj/mJAwTKhqzt5Jn4tDEtDpAtCslUnpVvZtx9R9f2KHBNTfnu9iGY
tBe+4OkA8uMpqzvWR/Jn9qdO08FFkDR+EmdxVj03kmQNml3wgx2Oquf/q1vgGo1J
Ug8AF3V2Dfilr64KxPDxDp61tl0e98QvNaMfMOR7b8A9fffzwJQr2V8/SJCTTnsw
BA9r+atjZ98L1hS+H7vZLI/DRoyL+xUTMFLW/nF95NRG1L35c0nKNi747Q0tYMNv
B+FIQ/Xas1fc0QC2MdukOrXgDzF6ZAaZpHqM/2wI3Fk3fCBqDkNqPliFlCZ8PSA3
5dNTz0PW7ygNgo1oLJeOYbeZlUL7TQYHTCGZgceGSVd3KYcaeoI5pWN/66bbi0g7
KBqZ6UQms3llGS2LaT+4GCG0QBBbzYkU9y2Zt+Gr0xtPVkO1ucVL7p4cGsgcizy/
w0wsxWixOyNRVSddbS7d+t3NZjM5Y4zZLoP4Hm1l97/0CVIMnk0r8mIEzevTLqBa
7ydQOCXpo0sYuu7EbU/8bcMCKnI8etTr3Hu6RUL1wuDtl2f+CG15BTDfwHWC8wEo
+zsepn7oMAI3Tlots6+mChOe+zhyfZMw10FItlas+wf0UU3fx6WKMnz+nDTYh2xu
5AUrKAg6DQO7VVtbemkiwrkeGG/YI6dMy5IyBYL+FfGhu6bzv3i0Jnkk5+klDY+w
cXWu5JgJVExgLl0opIwM+KVdM6ces+N3Zvr70hODpspFNswZ81vg+P6GL9KxBLyk
j2d2E7TCFe8EqiLbW61OmlpRYB0aiFFgS1Yjk2PsXExw1BSM1WFILPB2s6X8zywk
yIcAKZq4PxRjxAUokRP3CGLPLSLkSP2N7tBv8bezoHgZYy9haRSjOK6NbmXCrMhw
3mrcpfphew73VgTO2hl91RMWomoijBzXCdcS8mu7QqhXrBu4+EqO5R9UjZMveNHD
ISWZF/oY+N+yXwXRvJ4Qh8/c6T32J5zp4+mddt+gbbycZr5faXB7PJsjEeJgOKu/
3KtPe2zVASp8htTOXi0pZmy+7I3B/BvYwmW78XEB4RZMMkZ8LQ6HeeV6HFups5IS
Kb8YGYnnOHj1FTGpIKDJW016pkpeSKZTDTDIPzT6QAZAmHIupny6b/p2fkoxwSto
/j6F3fJnsulUFkRba0UbK7wrRURttw+wBoazoAW02439QlC/Lfaw06K1RgNtgK8r
6hxO6ZUJjf6h4gSIzRqlByza0BZByLNg7k3kZZ7SJ0hZiG0Fpz+dklg+iXSS0aEl
RkrzRL1W840F6kD/W0YEbI/H3KFg1RIyXqtydqZCBPkLGBN4O8rV7zEpenVFVdKL
hJQFKLaByh818s6vpjxVbMvbEQ4T82UD7T0ESKbIMrrCUn/yOzL2qqgn8Hpa74SL
dpD44bM+6di825rOogfgihiEZf3UtyPu1YRjJFrea/wTRLY/pPXJnxAb11MNv+Jj
XhRwcRHBxRnXQWlfZtFfVzfDTQ9B0bEe+c5ESWwGkoeEEBpZpu7SmHjhlyMFXxlK
+6GZ5CP3q5zebWrdzLQhi0/tJ8cJLYzid9btse76ejRdwJ3GRk0ZZEyEG55h9gQ+
a9au4L0p4I5+RBgXKrjjS+RT9PeWFVHSIY4xI1jc+WEKDbKrDzl3XIgHUw+fvqiV
2FLN3JYXQK0UoRGRwQg7jgof4B3oQENkwlhhh588zDxiIPsJJA1LaozOZwTsRi4j
LE3/Lkm6YvD477RSO6V7vB0Q/RDnvnGwINPG0dr+kOV5x+xNl25UKpzDwgg3fLMM
jWKYs6KJrTBP8XLvZdpBaO+0vs/mB+oGq400+kLHoGYUZIRzo4mwD0dllwt9pIqH
oD/VaB54RiXKRDCS4/e84roCxBNPtvTKdRPRRpKD+A8=
`protect END_PROTECTED
