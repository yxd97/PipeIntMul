`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OyUDv0sLXzNEbi4RjVei4BpxbFs+2/4Z+oJ0D0Rh5vKJnbYPG+RM83MgSLKVhUWM
N0cMpgpKuUyEjBEdciwKe7t28v1wlXRyX1e5UzzA12pEGD0DQWhE+e6GgBcBmVw3
sKj39wd2/Ghb9OYg8PS4HHidH+TcoHp0vRMNPDUzmhirZut9Q9bsKmPmSDbrQpNr
tLuFjOYyMyjmq0zWrivGxdY/PGgO0zqniiOYprDhTVzpWwHaPUgx96Wfl5gCy1z1
tD4vQdxEtz7XqrR/ZnIwusfsHE4O+GW3n0qoET1GdmQ=
`protect END_PROTECTED
