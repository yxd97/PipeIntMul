`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLpjQl0ZdsJITY02cm+fDxgY3x4zfvE17gM7el+C06lbnSzkW9kyKOM5N8RaSYlZ
An82Hy93fbSp0OaUQXu+6NK/rM0OViZ0DpzOk7I0rkfvWy461R72CzSdNibVMLqx
/bvin9pvp/lqCIwAyT+CCaLZCPJSeJuUyOKT7ds7Zqp+VEb12qzBlPwCEoELg8Ji
ZBef9mxHSFUXDb2yzc0/xTFDaVPhDuWMtESX2hKTZaKBGTn4RWtx1mn3DuV23n4P
Z++bCCPurLI5O9i38RC8CI8UNFLZn524EBFIeC8wdkUSq8Q2DotGgiSjILCI+RlI
x0P5v11lUbxVJQeOR8Z2VGtpho1H96kTsZjDdmWkgKB8qTyrqfXzL1RkjGRq/zsp
smYy9jSbgMoB6YKylAWW7ybwHOZ6ZShRL5+DMAsaNxeh1Zdya7JtM5dkk1clH5dI
bC/McLTVUC/jy3kuYKOmiw==
`protect END_PROTECTED
