`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7/gq8JHbGCtVvC8/MS3NuRVxEyLY5ueaClaaNdUd9pUUFmTgE5P4GRCFSFflJNO
sLycw7k335XS6ip2vnO2qiL/4iJ2eOnBlYICSRYfg13Ztn8uQcvJToz6DVq+4IXT
GCbglSsgj0rKGmu5WN/H4inTNXW2owp0tuo0be9p6eXJrDWPXeNnBQoIyby530ko
tSlFu6D5Q5FM9mvIDapx9RDMMVulYPlGwpPNbni6FnuY8/R2RvX71H9muH9Bwo8H
`protect END_PROTECTED
