`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aCbCp4BW+5xZIyq+gqwdREZYKE7w9rM+6i4HYF9vCm7uxVJ/Afq8CdKaOe6b8c4B
fkwRpkcFOYmPFJLW7WgtstkH+Ha1CenGL/Fa72PRPtio2XEtHsLWWAcjiqizpOnL
Vt3HBqCGYlAhb7Ity44vkeUq+XYCX8OiMYnGE/4UXgJ0Ibora8y6lZTMBg2jY7DN
qFzbZZwT8AVyqiK0OTwqnzvI9bdWWNeK2TeBhK6LtkaGiqLG8M2+4jy10Kx7QiHv
DZ5IetXwYpeWQt2PppAHdyuvmTWdlkkgru1E4MwKFPbcA12L4uR0d7ctQMsdtdID
qwKWFkEkUc1F7oYSoZ8uX911QB31lwh97aIviRzvcFI=
`protect END_PROTECTED
