`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q63gFz7mzrBIsVUSTRt/WSnMhTU5vhgfDoQ4lPP49sFiAbW4irZpW+GGwKXNpVr6
T2Rp6kYHrnJ9j8QPeT9e6J83d3fLd/9wUiPAuNisZq9NXrUcq/mDdFrgyYxUkUMh
BsjAO3rEYaEoGzNxcub/Z17Dfncv+7yppZiqtttdS8CQHgtwhmxKPdwQtTj1xKFP
YBuDoN1Eyyya2cBOeosv492RMOGQSAO6m4aLFixAKcfJjJ8JTTflXW/Z0WSw+wMy
xKyFw4WaH29kEtSn5pfbgkxtjO6hg9QNmZv8MBXAWoYCsn8TCO7jQYylCh8Jg0m9
ib39MsWcGwj/HTpwLWe1wEzmkmXRUqZCeXfbHEJCSI/Idyh0XahIRrASlMu1uEHm
QPVcTIuBFygmTeHfATaQXu+Fwct0p4vbOjsNfbRhBuh0/yKOWvqQTQb4GfsXh66C
ntNVdZyn+ac1EHMoUlqP86MFUQY31/cA+QGvchiKoWkIEJ0JYlcovn7q1hDdahPE
6NhAbNCocEqVHKTmf2zI5aerExv62poNty4SUSDNDgcod2qacQjul7zM2xDNbcqV
R5zFQsZFKDZjwe0qNTqhYAG5Vv+/0ImcUHprsPM4VAdIInk7tWywyonyRm7QW6d8
sVJJa061Wl1fqOSqRAYNp1blsOjj20hFsaGb43H6hCQsujle3TBU0DmUxb2TrTi+
xkSGWTIXbcH3cjzKC2CSIHtjC5NM1I9vWP+MyqX5RJbFZXzmFyBP1+W/RonSlP/K
SLdK+qiC2sdNToGpdPQpIPLRYf35HRe3tmdxNf7lBzJuOCbYnHGVVv4YTjCIUZ0J
nNC4io76XHhk4z7hr8bzTX3HQg3EIzoZHdoGRtpJCOozipjCnYYkfeya7FRz3b8g
kNUJVlyAx2bxd3+9wmsOAm1B4vfeilIrv2EyJjiW8M7fpmUxIgwGZ55WBMwqs5U7
`protect END_PROTECTED
