`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z0BcoE0/RRZg0LGvOVMRgUtKxJRhRK1Mvyszp0XHz0NgFKgHwmScF8r1gNlYFH2u
iyIdPPSwvZxymLWoRAXUcuyB2czr4CUNPWNYsNSZInwY1vtXx1TL0KXHYzCwL/LC
I8NXRueyaANRzr2HjKgnwvHgGHjsjmBwUqgr4JIX4QJJkxpJhOcwfikmSBcG+0qj
LUQ1Buow7ENFOr84RqNR5QmgT9VgUDtKOEFhBm1GeimEgq6fuxzpuDLbNAcaSAAe
uGJ5ADEkoZzX3dEgsL32WEXZRx6LotzzVxNMKuFknnwLWDFFNAeAImAeLfDWpfP2
0QAyEC3T5J7j9oauHnHNj0wUPtnsKFwf9fDep4Dov7N4Tyb1VRLXGUTiJrJxuLTy
80pQ39wkxqEEufMQ7IdhOJnDCCtPG8HNsQbPTKZB3uY=
`protect END_PROTECTED
