`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VUh7i5cfH7ClKlYH12oUF3eIWGf6n488tnoOuAqQvstwUE3ca1IAItDciluTCpJI
evAnVMO92hO57+fmaVpmO7TAYH74wVTHQIBoWcJb812gSJwAsE57mnR55HknHijk
qJnK9u3HucqNhccfqOex3LgBXFuj5B3Uyh+unX3TMfPF3kXTF9NLNQAF3PqdfKr9
LPDhKGD8o4ukC7J1znyIMA9D7VzUDFLUVwmj64enjeJZ2PELQ87Nydp5ESJhZN8d
gjj2v8bcPkQUkBR5n28ZrN9vcU3pY5Jz+Huh57xO4UmufAgk2X4eQI1UNHtWKxpF
Lb8sXfRa8/sBB6AtzQdQoefTDJqidRmeqG3XzAnGzCEFzYKjy40nsXc5BFwBSbGy
rg5ErxTd/gRLSw67dnY25fm0AMVB5nxNhvm4epy1rcyRgALjxbf7I8f7i+kGs5q2
KFykz5GLbwBVgHDNe93dT9uRnTwoGdkFHHz48Nh8DpAcsHUf8a6IKQ9luraC7x0L
wwZ74k2ei/HlpDOF1eRizWE28RPLjwwlvhSAVs6FKFMYYVxgh2uRamoeZfIogJcf
pt1RF4CJxVymwKHNZ8HEXsjYZTshISGWzXYrvyoZ31a/xsRPvkqQc+XcDOlhsjce
H0D1f/PeTADxYhIoM611as8HCKyjBJiw6UG7Y3fIVkY7KxwewWjn8fMgkwhT/VdO
ZFMJuETQniuA7J4npL6R2fRq55518RYYZW537RooF5VXrViyapmi/e59jYpPdj0o
zcC7UMmeKdIOQ3Ka0keIbciFAmi+gYqADBgGhsk9J4veikmGJEO2Z53UsvJB1/wA
+t8h/QKn4pLm2fP/5AYNCZK8qYRsFl8JXlVgYoO/65ZipFcpp5K2XvFjqCAPr6AG
HIruCqfTTArvLT9Nczf7AV/R/sOxxW/U5+WEAyWzIzMHL3pbIHIaT+JMAslzULxu
YEVQDtcD0/zYr3dLaR4yL8aTtmqAMBnBvSghMTDiwlyswleVSLMyY3cHeomfR3Zg
URc1F6ekaLXIxCk575u3qEWKmw3Kh06wT7K8QYF0BSXvcxm2TUIpxag06eQ3VVQG
e+bTiBdNgD9etsBjU63rQYI0yYLVw1kuqJWW2uNUWS0=
`protect END_PROTECTED
