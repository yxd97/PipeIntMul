`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LX7gfMGJmgQdJfG5TOPQ/aB+0cusWqQ0IPgXRNDVPz9ARGxIHt7+o2C8dgFdwZaR
+TxBn81mNMrX/w6G3AN4cJtb89GhyFXjuMmVa5Dg50YJYHVneJ6FTdlbvoitfmtj
A2bEJFueoAoxPoRJBlrFVurMS4N/L4k1oBo0ouew8eqO+Xqz13yv8tuYpcpXqUGQ
3mpn0VGCJgwqSLzKYWJQxVFZua/EwcBV4V9hfJfaQomEF39T0VL11Mlk7ZxDf4q5
K/U3ApI5EtcPzG3u8kuJgQImgWfhEcEViaSqC3iu56Y=
`protect END_PROTECTED
