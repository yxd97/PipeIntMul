`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ipnDSCKQrBL56Bja4l5sC8JOWH0tS7uC3KgZpFQAGnEx/jw4fVa0CXnWeWy05e8
eI7jMSlNU8lC8I+Az6JuPim/UTU7HzuOWl+sUXcq+6FsWPGHiYIvxHycPBx98eMV
623+6bkKPxuzSyKf6/L6XOzYzHIvmgrIsHzHtdlONxik0T/wwSLy3fJy95Tnli8l
YUepxfEMgXVL7e8OQBkLDV9/g7kq7WVRPvN+g2fhWxzAkJhCfssKiNAVgu3wYaPX
i/Ztj/Kdml3KpYgkusqJ7aynRnT19zGwdDRkhyiqJV26UAxb7H0HQid2V0TQwZAM
8ZxzHzsf27iMyXTAZvzy04aqtGa650kOsBaOVPQaLrXSy5Hy4lyYzFe5vdMecIJ7
MzOMlT4Wh8N8HlJNYh2lCg0lXWJw7oGUKipvmZSzdjL0T1iGpYUM3RlRaTsdgQwv
fFm09ROTOn+bQR/ZCRxZmfI7H5kn+rr8WJCaAnFLU5+ncocuDYu3DXz6ZCeUc7Yp
09XfO929ocdo46zWurCh4WCaLzXt4cVht3f/VasrWj4luRUiX+P8j9FdH8Pe5uLK
2byipdcQwSAANg9eZsTwxfleJlXfNxNWvihr6/V0GTwAyRUEJ5ODyhfUk9sNeuq8
mUD67agTd8SQYhq3CjJRbEbatLDMFqoyZn9KX3519GWkiJhTJWPWfu/wjdsmF6gG
CTzKFypEMEPoVkrJUF/qjHe0/lfXPyL3W3qmmgX4oVkJ6jhNHr5KDdWMqYZfAm0b
VHl/bBQmNTm4/ayxOnod6Hs/WyNCM+u2oDNeqhJPOXY=
`protect END_PROTECTED
