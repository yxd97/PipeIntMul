`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o6uaNtb2nQE+dEDMvgzpDsMoyZs7xVtGTBVAguAsQihkc2FQhzRR9Lva3xTfJDfb
uhxdY3aJ1PwQ9PjCbqkEJ7FIGjfvKp879UjdmIwwx7bghlPUACGv9+Y9SQMGasW0
9jHJBtrQuePj4qcdnm9RZvn+j/BghkCOk++bSregZDphWS6lyR44BhbSto3eDzD6
GU76SDYRwWAOCyAfGO6+iRLnPoPWam40hZ1iJz9Idv0m2zj/38DMTdBdNmtG7uPH
sQBxKUCnVup5y4rQBgmtcxCGQnx5Wzm4pfEpANswdJEEyuPt1xhYWo0GjY2pH/Iv
1RiJA4M6KfqBgH8gISRWlLqHayFJ3uh/TxlMBZbcNiPIzO8a5MMD5QbRqbFVIhe6
XXTEEM3H+92dCWhfO4xMdgCfTbIkE3V/BsbL0Hs4Qh4IfTJWLlFpaldRtV326Z3Y
O/vz7CSNbDQcavrmV8iLrQ9v65fLrj3lYXwRPZB/0P4PiyZ/ltSpeDlmj5BfKmhz
cZfhE6n/ZEkyXsrWxmOfM4dk8ilKoKmken6v1RtDX+hi9uO0Kaa3UWCWKkPDxhL1
/6gMGta5wWXC6TX7LAQxvdCdogyBLPH9ts6Bck5bIsfUsY8C9pxWGav4pGByaxUR
DP8/CQmgbeTD5HAxpPo/fS/G8UYLyjtan7iam3odxMKss1yCna1wyM6kzZc1xKER
KECxV2qhzFKf/hfASHUQCtxtAjqOLSkGIGhFNjYQY9XrCAumRyZ4Py4UOuc83UkH
PyubRu4liRmP0LU4HKvoMhbOfhRR0BHIJrjGJjR11J9J4O2PtVHbjuFy/wsK8G3k
OHzJRRTGNitR5a73KqqJyAF/wn9R7rXDXPq9X/TF+MMXyC4EwiOVjqGtSmRjG9vD
oLhbBkSZ9JxdMSQnwNciPlPFA8Y+TUnJnQ/zqZr79N5IsAMS73AfWJ4n9dR3bHhN
ud6K8qc2071mCOHZVH6QfkN9kpYVAm6GUJ8mrgrb1bdCGXVCfekB7OVmP0hiLXUq
jH2akTuP8zATqY7c9TGzSg/XmDf40F9ppiFH/085fmj3iTVfnrtGx7RJ8Q7s87bt
Vzb3CBhavqDC1XQ5sspNE+MI+zzEz3ALDlG9jO43tB7d+5sNjyOWqfyizurXKxod
4f7LUuiW5Tyl3hoXp+Ug0Ys6FjMSsFavmSlqkx1nLqqMhs5IIDFAk2NpNkDO/9Yc
0tJmW/eI/eHtxF5CDu0nYL+2VO6abEDrrbaGsW4fos4xWSXFFJutOlqxe9LMwYHc
XfQO++ZGNI/T297+lVunkZ2xUCVYn993Ju7pRsmTRzMDV7sIc8EwJKGXxXUj5iFR
B4knoJDZ+Yt6K7VOWBtfZnTaESE5a+Ieve9mjPWIA7ePBIXfN/COPVbeRJRoX+F6
0pmDe6iwPgRSEwp2m10PrwCWaay9lcZF0EKt3Lfum8N7d5fA7aH5Rh3PDR76Dkup
dJx3dawwDYahbrvxFnaTvp6msa9dL1XNrW4fw9BGCpjhWC9jPbJCbYtKkpP3kM87
frRGF01ePJ2u4pm1x6g1zI5AaWQO20EagFBFyD0cRslaOGMxjPzxOIADTptox870
S1fq3HDHLmBkCymJ/8FaV8PjRgNUlkkjn+V0FoWW63fu0y8koIIX5yk5aCbIRA80
aPiUjRayLzO/rZBdCCcoEw==
`protect END_PROTECTED
