`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1hPP/xNkbTYpcE8qpi5hXbo2hAUawo6wAo6e3sewsjNIJ7mmeRU1cONm7mo/dwr
LMBiC8gcC+uU8DXFhLS4hDrIunKYsUJPDKvw1aelEfs1cfTl2yC4VX9J4l0R/VC5
wpAIS2KAXIvhXOic76ibcrQZ8wFzOqD+8NtwnS9pM3azMUXfQ2Hd+SKkaQNFVl44
hbcavTDdB6Yf0NYzyPApgwQGFpuwxDpcGiVSPgBTGQwvkCnqOnDq+1y04v+WEt9s
w4a0G5RN3jNr04AtDc7mBpnYG9cC4Jy0NSy5fPzGUaFvUcJDkoU2JFtvAkh952w9
3y5jplPD2yXy4wlgeX5qfkFyTxc3N4Uu5Kn15XaNur+uomQ528ww2r+Hu3t+ERt9
SRQrnhmgBfoCZIljERsiVFZW1ZfFev5THyitRBTqZ6rYRzZjT4QaOFOit2qnL3tv
uuqhj/FkRv8ZGY9y/6mlfwSSF/DzfnwEcqwODwcofYmL0pdz67NIOjNTDl8e5ovu
5Y0ckbnCH0ZSHN65KmAy0lJEBqOrGlCF/rpeS4muaP/ABHsw6OPToHSBo9MiWjiH
MxvlPmOYQ8m0dOc3Tc2jL+1mbZbeeGjrl417qRVHoGVv+9gju/07CV9WgFJV7c7F
7/5Ego5O8X4x1EmQjLtZuxaI89FcrDmX0UrTauih2zrde7+Jtx8ioJNr136J1grY
BUiZjrmxHlpX/b5VAb2Bjb6F5LUI4iwwZ5cEuAFfAp8=
`protect END_PROTECTED
