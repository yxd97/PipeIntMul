`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mskoJO7pLn+sRecR1crf0OzHFTzfk4kkbJ04oonURr/OOXo+Kpb+fi+NLm5Eo/MK
USJONHI4yjj1pymhi9TjQpW2gk5qq1bDQIf+peazvHFPRYuq6+EsQQcXvOaFSdbC
dWWP1FKSrkuRPOx8pq6RzB4tW20YP5OIDv1WSvjJUAWzYkL79hkgPY2tA3b7WRZO
bxs5IhruZs4CHyETSLojdSv+WgkQy2Y5MQEFzEU4/uYQWiZ2h7ip03s1hEICnz8E
w/5HCfNPjhKjJlnSiiXxqIswDtnOzczK0yIeBpni731q5Qijs+/jEjic2Gtq7SAu
YPdziFmwTcAqTsRN7rMH7UTxUhBO8N+q6WBlUe2J64Y6QnzqgqB59f5ybLhG7ayN
LrXNZikeBZUqRS6fTEfB/+ZUn1HSeXkJM+NgPJ6X6qdyVasNuC7qznm1pdkQBHaW
dmk6fQVBOjIuY5gVIOQMdKXOwGhKvEjOdaqFEnZ8ZuEDhc77yW2esbNfQiLvuuMq
cI+h5wchuhOJVS2NVsE2zUwr1NbUgQyStdOlvdu28FqyEr8AgxWsxU611ARBAxXo
COAiHirjv+DHN6MfhlT1tOBbyyuZnmf4J+gLh7hRoT06pqZ6fE+XmwdBnHoAKNuJ
CYagmbzCHvAKgps+naal5SUJ03Ro7aFW/cyb9C7Xgk1jdZuAS4hzIRkSFvWhcUBK
3IeS8Kb7/fS49LhhiDXTjjmqkyk3g7jZF+3WHDHMDuXIJQoRWicyAnIx6CVomQvi
RHoM5og+PVdBHFTeyB9XB4ubN5y3UT14BEvHZsEsBhWHS7fIt1Pwv4gAegpwd0pu
ESLUvWOZr0/zbqpHzKz00IyDbymvBthc39HVSJ2bjdHlgiZh4dsOX1yhaAvSkth9
L4woBhK/UzEUiKr4b4g6786R0lz1egn8CibvhEnMlfL+FmIaCa2v3veP4YlHI7+0
RT9SVJjbpjou9r5tkdezAbustNFeacB5NP6x+j8KP8tdBmsjGCzHD1eOI6+vmlzi
6fluAJhgfY0yzX3BgVTgZo9L3HvcrbMRWQOPdrjxvmU/wnM9RLlMuj3Xf252OvgA
btIhXfqKQ4c0/fwF0iydJKUeCzbvPu5Bpdd+CmldVQzAjkSJrhQcl5t0r98wCgTy
dWjX1+rOG3ImhC4AY3qS7mvr3GL749sZ603JHVC4HzQJsOK6QkKmWeRuPq8pRynY
jvsUjo2IERiqru1Qx0023hP8s31PV9va6CAyrbQ8Tru+dgUVGWxZUasgmSlimIir
mhm/bUOzZ18ET1eAqIb8ZRbanVZQ7HHsqLGhkIPiZdDNtQ+M1UAEM6Fyl/dN16ff
NrLbapyRmlrNh7w9E1PaoM+L8jCBsP0lIt3CBpvaj2wB0N2+YiXPS2hpU3kNb4dl
+vSIBntNyILLsWvV9d/sliDRlulQHecLfX0UZbQFrTW0ZoeibcIiq7nUo5XUOZB+
b+O8/0eqrZFm7TB+kV/9qJEQsMpUKl9ccTYimrYEaz3QU9CbcJWHlIN1cMk8w5Zj
5/lO1ALsmKXA9on9+QJZOjDrCtFj+QThCVkp2M95GSSEuUInFlqgJyhRy4fmEbcs
LWkb+rm3/47bCY5eG3Bks7/pCCpKEKcxniXr/+9LjcH88UVvuK2GhDwF80LP4VgV
GR+YgSjD4fcZJkOz4vIxTFaVyVldf/7JhHM+t3m6WiQqXgLD4baORXH5WIE7fnY0
UyIl5+emP+ZxY/nipIKyyyWLcXBMMmmwjyCTOmZ2jcWIoPlN6JEuP55k6ieZZ1dj
N9VccMC0Qt/QxfFTBjpNnMwwXavjOZ0xQNpGfDIodDApv+XbmgrLwRelQPwxzKRS
PXp3Fl74SSy2bOGguvzaIIupAhQhhQQmWGelGkrKiq3yPGHg7otRqU5BxCHZ99bA
18Ed7pBO9R9VTVyCW+tob0qb/xcZN7B4w35/EQRtXVczOa/g3er6SGsf0UXYbkPa
GFcRVIalqaxc/DFV4p7PEhHwbujFu0Qi9BeqfJsqYafD2MmZz60ywEwXzR8oNXE+
/mobTKKhlCyrG2UiamPclOJYwyUC4vaaj4i5/a/bGXez6vzspKRSLg3FnGXtTlms
t0Tqnq8cU0ZGm5qWFTkUfO+jpTMfXW/N9Rzyoj1TPL9aj2CCx0L2xDLTiD24X5pv
RToJEA59jwLL928VWLFAd6XKOMRU7oCo9S4bQ9o3rJkB68KYqpr4kabQOKKCdmxa
LV/0+tUW8gtStAEghhkj7zYi3FYiW3mHPFCgUKE0XQ865kjVzlBDSVIrnGT83AaE
B2yFi0rIDx1ek12ENabTxNxSeHnr9lQPCj5QPBJP0c1Q2rA32BWfvldjxq0nbaAQ
5Jha3Ns+9/wKTVfYoJ/wKmObdzPdmyfK7GamYF2+MoK1TmCbyQRTIoA+jWABT8eT
hbnL/NyIBLfV0eTSqWcZTMf6Bc8gDxEVYZnXzyemLbbMqTUS7L9dqRcmiCQ4GFDT
ZF9kIHFRUoBepXlZ2h3uaPAUJH7W5anGfPapmclm3K26cEqUqpPP5kLUDTTWj4Jw
J4ylfj/zDw8QScw1Ek+dJCCzlk7TDML/Dkqedbt11VgPtQ9NKeQUzZEjPrEa2v7i
pY0tzD+Hoo8J8fN3JabzoZQ48Nq+CLxu/9DXxjAM7Jw=
`protect END_PROTECTED
