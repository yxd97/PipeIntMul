`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vppCUjWoAGJ5Ho846exVOrbwO0m1iaUsOOzgvQvTiYEtcIvo2uy5aDvYQdNA3WUU
eNjHnn2kOs3X8FLn1F0UO++PVFrHtqX/QtS/Pf2+neWhgracZpMZiNKQF5HGif4h
32LCCUWvLIPzC7xksS7oOUzt5FMcxjgqFTM066w9Ny1jRzEa4oiC2sjQYbcMUnA+
HjHm5axSQxAhI+cUWhvfnPT1L1f1O1EFLFlyg2CZ6k/XxKtejBvLTquVBf+w1i1l
D1wTLJuhFOKAKhYlAmL3B7rQTIhFvKRtAGDZCZUys0bkCAq12/uAS9SLQXuQiCKr
u4G8H7Ueq+TCYW2c5b8SwHUaBvsrh9t9wiUd1X4KG6+e6mB8Uy20vYjn4TMeBUOF
gvod/cGOBdkAoljwSjjcfpprDpAsep2PkQ9/0/Tx6pn7lZl/LwfFCyfCr+lJ+ru0
eivPjx/fhEnmJQ20AT9FmrJafeXI5KcbulCTihrjSrehnNb/D8Czv4hTHEUKKm+O
0qkFq56EEPugQEv+7p2ZAy6i7TAvj8chCiRu8B3rllQtoXqyACEOWGeujX25Hrrj
gx4pN81c+Hm0AIv9AmJdlUuBSVN/qM1JdSD0JhGepXd7c6Xf8ehlNJ2u3P+kLH66
WiL1vSIQ5dvYtDaCy2D8/A==
`protect END_PROTECTED
