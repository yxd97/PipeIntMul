`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yiGYvPY9zQCdP1qDzIgEdmVBw7Gzz7ScXZLxlDkkAHSQAQWGJowWYZ9sJDkc92Sp
rxGJhUUNnyUyh/7+KD22Bb9Xym4v0UJG2JjEOPW8jNpUwCFIYaOsoHXY21fABMc8
YIlHWSPUHVI5245hlDHmuY7gl6s0uEgq/CM28CeNjxRD8/2acM0qqemc5XWXAlsR
eBLaOpmyM1NsEUBe2XLm+146J27lHTT2zopPUlWUe4d8faclOzpe/AJb9rDdaxhJ
czWoSmKwFMq/ObKKj4UjQhg7VEPPKucU5AaK6jAQc+IxVgdYirWXmlJe0RcdmGlm
lM320Q9TYv8cVcdHMtKywA==
`protect END_PROTECTED
