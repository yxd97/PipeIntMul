`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ob8RIJA15yPyfgdlqyLWNx1VVxtx8dntlc+PFmqaXTVYnShrBAipKY7zMxZSbmcl
dpEl9NRk7BKO0IJb4fKXo6i+vTd8n1XgfcQCTPRZllH7mIr7Jthqdhu/ouWKUdj4
Hr9exlzpZjLnqRzHUYYcwxmuKmV5ylPJHwAeG4Z1UR49ygzLGybtFlOtqYK1iBGq
zahjAzX7TOs85Q2e6Q3SaiSbS0BzxcdGkXAhN7ACs6ctoaxZrAX+VgPxypB/gQpt
S7/d+7/JIytlrJj8lhVo8xR1EFhHyOkRbs1S1XsdxvZFi4KImvp6c3hvyBd5dQcS
eE5DD45Dz/FpeYgWHw2b6OzFVc0kck6LL46bhlKH+BWhkItIW2586tK5NDahZ7+q
shxLmkZGXex8vaH5A4qtINsHSgTSTpMviGNzyCdD7/YWTXQCH/0gk/5/BfHra1lx
h01VXK/GN4pGUfBHUNGQdG1WkvMr+EZWLxCwAfjkeHMzlANb714g2wJPTS7GlPai
dfN+xV5mkl+0NyM5mDkJHC3twUVusWzV1qvkl/lmeYA2inhTgvIJn2IP3Y5BdU6o
bHHwY4zrDpnma4ciElps4oHL/vTla+55R14/vnRPHDzMJmJ+B6gRgU0w5rjOWhCe
iezBEQg16Vtq/fn/K83THmzZHhI9q9E2UUWZKx9WsN4/E6euqlNfsirQ07wOHp4p
1rztfbpFdki2WpqZ+5R+skYx/EPi4wbx1G82kLRzzItZvfKItDdLZNO8EVlAstw0
wfO5UL/NNQnyVzQgXym67/ap4x+zTGDQpfJ4UH8MK4s//jU49OH+aDwTFBcoIf9j
X6o5dfB0c3dMcDN+BHDrgAmIhE6wJRohkrBmx9qj+/UZG2+DxQdXi+aEqwmeeg0U
7B4eRE+1eY5oJ9jLH8zpBe/sNjIx747UfhV9/JocO8+4uuKQE08bheRgJdd56xAf
`protect END_PROTECTED
