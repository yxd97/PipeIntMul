`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HnBO8+6Y40JcnEIyeijVpCXMerD5ng7zNtrOdtF2BMOgy9mGni/YElwN76d5HXMo
zOEepBmK8JPdglga6Ww75sen5PXKhYYZ2qTlJF8DYA3cfCPnHKda7okRCoSyGq7R
8E3tey6TcRdt9DCXIDmNXSuDM/TuzQJzFxtCwxgYuAIdkL+vq4fZSoUIvRwOEIWZ
Idycelr0cmN1c6s956ZZNm3McsL7mVwE1rHyLMbgyCGBnb3YXcwKzGlfX/tzHzJS
cLiOp7Y+oarZ56f+2QcwbCrZcRLxXwVmoQGK/SBqvi/aAP7c0kqM/npZimzSRhSb
TRTet4vdpUEX04xygwxvHw==
`protect END_PROTECTED
