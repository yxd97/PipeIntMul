`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IfGAiLiJm4w15ZkfUF8UMSG2bTBK/rYUDDPcGMNlMQe6ZN3zgmcBQW5ccnpuNA4N
zgnFruURsIGABpV8A1ujHlW6lg62siufX9GId3dofHGdybgtP7vvW0w7lJvmzp5o
33tTinWDV2HUenAiAmz2vE/IjaNls8l4f0EJZUQMsTT+7h9qBn2HejIDhD1CBrpr
8bPwV8TguAAkDZto+rQX6W6iMVWr4g2mz+etTiw+SHTkhuQbz0TFHSHnPsMYz7iI
PAVAR26JDkej66IBPDKOVwbvq8NA9IUE1xf6Q3AZ9KhHlbBnpPIByhhUYOLKGSNd
qb+yJJhNFa/hKCpyrMplWg==
`protect END_PROTECTED
