`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ip0M7PvVKt0XjIdcIaXLahrpEg1FPBTzABi6qwPcO4MXnHMHeiVLWgY6UQQfshkb
Z4jNmiL4kVyFCZvYeEZ7CpktQ7E5v3R6c1vUBmFecPWI33P0n60CXpb2sfQ2mxzY
yN2HjTLYDWHzbggzekBt0lfBdel3Jyu5Mc1um45U/eHEmevA58UsRH/4B6G3uT+s
mV8BHmoZ9IYh2Wt0isTCHkegRM0vT6yideqff+4BfciCzDONazKo8TaKoafyFSlS
a/upOZ5H0Q3bOeXwUpwoy0gqWJF3JXHpwYSUU5cghiehRIW2AFMjzbsNZ2Ei4NuF
qiqGy5ByPqvF5+PMgvXkEpJpdzvaEdofis8nYsyrlHVyytj2dpjdO4yuUrgznq64
RNEbR6V9W1NofYiDy4otFMEVedKCccIKOvbdAhncbR3CWUAPulDEYNnqvato8s+e
mCy3kEFCHtyDUtsmmw/Nt0SpLJVIXUsDm3G418/lSGFD3guNLJKLWOTjF3P/brMb
VoXA95vzdUYbvOHl597cdt5iF1CVGanTKYkXWCQTYzMJWJzSY1Y2LE53k7uVHoH3
`protect END_PROTECTED
