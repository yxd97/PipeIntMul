`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlctM0NeRCIYg4qqocOl/Ues2G7LqIj2FG6iNmP8y1MP6n+PHVhhDljSEsS/PhSn
rvCmzsJ7zaWJLo+GaGAXLvvMQb9T7Vzbb8b07fJLm/wcOAWvXnhxZwqKjCieH+lI
a5cF+G3MSa+Rhiok2TjYWLHNkM8K9hRGUrotYL7FQiK3rZ/PV0aQ5NBc20/af3xN
7E0S32H5g42bN+kw6rgUtUvFs+UcNX+l5zWWijhiyFIlF39vczZ2CzfJv251qOSY
AmLmjLOZcraFwAfN6Xf9eFGD2/idKCG5tDqCW65bn3an3s8Ylj7cd3ypJ4zwhO3g
s3Mn+li+fK1V62P7jCR8pydLLJxaPs4ZQVoUuZCbBA+mC+fP0D8OCniAiCNUQKAu
gM7DpGIrWDYm6cpcBUrcLse46XF9ZTX9VzO54G85C6R2fFo6kXWikMutpxhPGiYb
lFViwTVIBjuocSYGmT+9WECgJAwWszTmKh8Va+w/dTo=
`protect END_PROTECTED
