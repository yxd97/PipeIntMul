`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RqhdmJunvAy3rBi590UvmYvlfy/I5Dpu/g4mcEPOKUOUSil7/A5EdvbTneKxhmcW
lBW7zvPKMSlzDW2kqburZxHAvfY7ZciyAMAsE5gff+BGC57wxYryuwG6vRC2LQ9Y
J5xWq+iLNfKrKGUVDGBjvY9KMcMQMBYgWu3zDTYULfF5W4CBIgskXCNPqNogafXc
2jxZDmIiJEzxDAEbs6MxARP4EyO8TpbZziUusl9wF91JloiHN3/ADDa1AqbOWATb
iW05YrkdOiL6scyyC+qckKnKOPbzRwCCCm2zFGSsw55iKaewDT17UvktXYOjFS9s
O6eaOY82ZB4oE1S5OgZxnacyWOXofXGAGY5JtqPG55EvU8b6PiQlKbUo1xDilUNG
NJFcEog/bEBGyUAVN5+m0Ztl4p641S6R3+rf6b9N+7g=
`protect END_PROTECTED
