`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q4gTrTj/lM2XHf01bMx9zNSGCnNPSgtskbc3KGlnaFJdBNCiCJR2bdDiXjZynQyr
SlttBkdI5Ze6DkEBhWwzA/SPO7tRCG40yZfqq216gQuP1gGV+AIMIJudnmQ+0Pfs
LNnJnftlO2dP2xmHhsL9eXWPBxyOuYJJi9vesmSER+7wvKl1tZI5qOxCigQYa/EM
gp9cWHTi0uwZuMG8k3mo6X8QW1CLNLs6CXVoMdQebHu0s+xXgEpYTa1QLzAYjdh/
bARDceHW0tjgtZRTMcEyQBeZsbtRsofdMkiIAp4naY9iZmX70c+B1rkAoXzmObZt
lD1aYbC5huqjru2CnuGPrISkBcrRx/eb1WlcODazIFJugC23Gn5tn0ptClXMr+dT
`protect END_PROTECTED
