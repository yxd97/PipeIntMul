`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iZuXXWYRVRkbptvssH5QdSTiHwDhFdIDKG1zizCjpjP8o+477cpGM5RjYwSBbnWT
uqBT6hlHr04alm0JVh2X37zseUT/hX5g7ynk82lZ8JpuKxm55lT8VcgYdCetSf94
0JPM1lk7AdTQt9VLTgXreulFPRzwRIuiWCB79RCuAhcJM4sbb9JEYzksNv8M6QeJ
toTB5HOdDA/JBEEyrtt0CwkIIK1TQwa2yHewyUoNReTkg9ktxr37jnEPf5BatpMl
NPT5XQBboyq8c1aYctWLvBi2V49uqegnTUJn28Lp5AitZOhdL/krogFj1ZLNRTp7
wsoo76+196kr2fDJ5cykg3riJpWCO7wzkQxRQ/9O5eFbc5wW2m5wrXCkX31GmSTk
G/gb/DDxv6wRA5jNVH4hUihv/QdRitmulKMU5SjMXyfJqejhvlZJfk6w/I6djGgT
MdOaJOKefzRMZ+RRqn48Xwx9+WPwGyyGf75JkN/3irE2ZfmMkO8mdEgTFyVCJty5
4Li0RZMkCJHlg+Cdc329/1lYBlWaXO3OTmCPjo47nly2yAs/nKwAq6JjXAFdr4pc
sN76aEFBHWMo0Gi0EAkRmhBS2v0+rdyrwQaZkVMOGkuQWexYHP3uwrry6CMpbEsJ
CO1xyBwCZOJykJ1UFOWhBYnGBjDiktlcviN1c7Mk7sr/VKEjLOdUglsNiF0AaU7E
TBTNVb7g8Klio6GTx54aogL4T7/GkjFYwPdrAgu67LSJAYVWhhfYVp4P7hDW+hIr
K/J4QPvJvoMS88jb7NcfMkmc+vbe3vKoLlQJklwY6+grUtSk0B6wtfpRj4UGmEt7
LdE1wpmgxD9I9jo2Q2aX0h6e4TfELW6ByIZb1pMoPFdM+V4DoIJHpFOai58ivI1d
cILiLVYawYnweUOwTaV4S/881rH2tfR0wuHoAbqke54CEX862KjMILff50jpjph4
k9Ph1CKNjtnY6kNJ2PxFKPn6VqGxL+eiE8a9liSMBjpDmDo6qVss9BiKJwMJsB11
uLsvZPoABTqYv3uqC9ZaQWus72d5GPxHrDs/QLrl+3LlcKZTY4udpYeHBBbOUsNd
uKnh4oD0q3VmPo0ygX2yGZedKaBXOKEnvZAdD7Ile/3QbawvaskbuFi1rC6ZyKBB
`protect END_PROTECTED
