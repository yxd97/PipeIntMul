`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ruut/fACEZEK3Q2PPoXn+50pHws7INtqK1C0u13UF+q3dnhSK/8+SalqZ22xUP4l
M2yoKGFouW3wX/OrPNSHS2esj4YK4uU7i+P/jNhwlgi0GBDURsFLucDweKm+gHYN
5AoQrgSs0/TtePrmwqi+BAaAQXU4qlZA3afDSNd6fbBanjw9LIu9qVQXmJOa5Vmi
lR7tXcs1GEtBG8h+dGY530NuxzPaHn2vXniygdCPYgETc9Fg/m/RFUHg3m0l+gso
jS4W7Qpar/NFpkNZTALMkZS9+kZoQNyItca+ELlmQ3rZRopOFycPAVKhfVX1qJmY
xziBaOj0NwKzp0KRTTZ8uEt3triMdAJEpm1S1bC091Eromu7TDCiOmKFp9lu1ooj
LQQYD6SUKotoBuhYP6oNFzdpjAPFB9325c3lKBUCcNw3rq41mtaWRl4Vv2iYFOyY
ShY7+1ElGFExGVc0aa8/FlBjHNlIc4aOJ9Tc+yr/wzEuFwSCarjUeArIM1LX3JmO
`protect END_PROTECTED
