`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQsWHCtgtId672hsFzxWcgAXDkeCGx2wShOhD7djaxctIcdj3Hny8Eviiygor4hN
uYweAZvOZAZ8ewnSAQgzz7hZGkJ22+XJ3sNUUCP7Do++NB1iACDz9jV0qZZmOzpZ
lUrNtP3oaG4F2vTBh/dN8+Gz5vHZmgMTh1tWHBUu+qBmLEApvXj41v1E0pDIVlW/
m4Gh/kQi1alpG3KJzbiRUgVwZMqmDU0IfZL8MPBhag7xM5/1tn1trdmDalw7xogG
nXQfu1xvMio7d8pnTNrT9RMWePb3ay/fglZYBg8R3AjaOtzKeydTIvnPpwSjR7Z5
qRQ7XAzCCqyJlGfvPKYnFA==
`protect END_PROTECTED
