`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B5LnYaS3Gs+PB4pXCHhj1F1rYaTz7oSypixMsgY771VN6rU2dUf6v3LGwNPUuc3u
rrXgtX8aC/shshBjsZsBFSAqZJcnnLoQtF7OgWLtKNiUDqvQqAt4eY3rtOyjrDYD
pCZkCz52yQFy5HozUNeX6qiWBOeUhIxc34byjXLYIUfrXUKfSAIeAGxJgykxca1N
CmxJBxH1IkyvUDXnLIpBcs+72KV+4vs11MOTFc2no1BwOV3AvQFDVf1QmQeLrf+A
9q+25syhMekTc8SEnCVw8bjQ2xbJUwjUU0aJdQwOGfXqyc8R5tY6FlFbG3y0tx5w
wVxO/PUxcg7bN4mFo+616WOeJmc13trzhpdKy9wMUUaodwnTYkA0bzRqy9Oe2U82
zRSmQHuRZeARPK7W/ntHtw+sW+54EDf94i206oZgtlUw6Xs10IOfXIadpN4/2hoL
oM+Fpddba54c7J5qHYWdUsvfo7oMS28Fls8ZkvldeZzmhpSyeLc6mnJWLWQOS8VB
c7ZEYtbxklusEo2M0R16muwlnhJ5Fu7TfsvdeCcQ2kL60AxhEDvJMeDruFMYE0Qy
NjH3IRF+cstZfKSp8txiqDRG6QxybOxG+GG9OFsxE8jLWq68NT03uq1iBztSACF8
Fgbft/u7ObZIcfghwvxi246+dTDCOzBDAUEWLTX/zE424wGix9ZYlfthd+cFqAPl
bMxCoZ7GYoPXO8YduVEF5M6FpTvLL9I4dlThx1hqhRPA5cHiCSqu8EWvV1yC1wZv
RCDRIo35ZrYWQ7db6QFc6yPF4UXvwf1xeHrKE7jfwTcmUIWBk/9DPFz3kwoZ0mq1
/VU/m7QsXyb0qH/kalPau9py0oEiS6oDY9FAIQAR2fmz79Yxu1QgybTdwI55wCK1
SMyxcZkxrVp+/nlWbkR5kYFT3Cd80bnxpig7Fuo1PoIO4uvxLp1AC+KrO2Jaj6Hv
`protect END_PROTECTED
