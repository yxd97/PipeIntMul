`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5u/Nabw3TKIfdh7E6WcjQ27Z/B+7Nhhz2tjMX3LBilklqZMhA+J64J5qBqWZbEAb
q7HSwRGYjg62ktpGy6DkVnH/wBFNfBKA4sOJyWwfu/VG95FgShZgqaUxY65zQy+t
qR86DvaAxAj1k0CA6S5SgrT9kHDE7FLIi76HLUkFOtGfAabqQgKv5J/fOTDWtdZG
jAzM8/e0dlqJs5Yxw8dNyXXhzWv2jWqaFGS8NyTxKED/mfmR/IiuTFsDvnZL+b6m
aNUBwinJIDX0zYyxlYZp6MFysZ1P8tm2gMZzewUzHmF90BzziaflzHI3ezxXRAyD
JTvaC0Re+zoqIqiw6zfOh3zQHeB+ng/l/ePFxo23gY34YdCUXPO1D2SH2Vhahwpn
HBNBATZG43cVJAkvP2z7zJFsspc5YZJmYkHMXYj2a9rKjbWQk7nZUzD3RWmEXwOr
XJHQS2fVGkhcljFSq6iQ0YKwov3AcB/C7mu5TD62+KCU3esxX7xnw2VT+/3OURkm
0HIDPqNuGyzOuC7ARlXKD/MYJPqrEhpHpYY95YejCfIPSD1yxd1PBUVju7a4wVQc
n/VKGIys0s8DNw0Gk3W6wXI5/5Rnped47HMvLjr0+qljF12BPT7AetkEo2ufOArs
ppo9VsYI+Ok+0A57kf4PgdqQv3PNHL5/XR4eLlfgwFEG6gAngPfS3QpBQFHHlK08
yxnTiyjHwxJm5lYYI+2cH/HGAM69CinTXPNkXhNrjzVfUqKSJj1yuLcO06s+7zjj
XhID5FZPS2HL0nq/VYx/CPxxXfy97cfBwojkOgR29S+Quig8PMZQgS4iMxj2WfXG
MF+77R6XvFUQGGtB6k1ZWLReC7GvyJhZEAHqMvzj+HxKxB1kCP4kjfHPx833pQE8
Q965aYaDetPdtaPNOnqE/ii8TZm7lySsk0MZDqyLRd0qyQMsdx5Bq2YEVOrqX7yM
o5C5jmRUE4XCC5NL2nB93qGm+Ng2V3Kd4SAPe4iRxtkr3ckR9/n+7je3Li/rNB7d
c0xm3pwQsGxxpxovqBoqAsUhbKdMtzHFu7PkuRMvpQMG22ObVDnWXLdjTDlDi0IN
2dCaUA/blMOIp0Ly/qR1xathjfaeHsCJBtWpmjwS7/xXHRYJPrPnsWizn6iicnbI
u3U0hwYfi0HajR/uV1aF3gq0Gi2dSFLuAXUrK/eng2CCK4VxjZaCDEKyx+vKfCQh
`protect END_PROTECTED
