`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdR8fG7DhWNl5s2fpvJATCaDxVlWecmHt0Jg/p9WzieWOCOR57MaBzsx3yT7A28/
74OIkiZrpbrGDIPnZt4Q5xVEURbaLeMFBwL/ijNbDM6EkeNFMRywcS/TcUjKoSuP
K1s02ofMsiTh1LgrWQeO5d1BbpN6RLz8ILMbRP9MuLSpXHY4sqtHrOikpcKW5jl5
01aPbQvVdZIHRvGoev6iYmHSH7NDc+7g58p6gkpPepeQEOZs8BI1c2SFm+dG+6eJ
yU4UeCjtRN7nnUrFyRoHXpKe68Nn3eJOysgEyPq/RMfzS4dVgu8JagsqgUuhTHOk
roz+zNBD5FVKQwEHjyVR204eUVz9SlkVGHWJ963ZIvubxCVXtNV7Y8/2VbbhNOOh
m0l8lwUF9Mis4qAmvq6aFdNRLTObN6p2fYt+O7OuEIc=
`protect END_PROTECTED
