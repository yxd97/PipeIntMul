`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqcVeMgR9TMd8adX4DuwJtERYXJeW9nCjSZ79iBCrXoednYtlxq58/J/aSAiS8yN
qbuh5pEgJ5TRo4pqR/0MIV8ImgwNYEzg4svjkzWKQKOSd8UuFybedDqKEVHDEwLU
NyQzagcutYWBQgiEiU8cyIum+DM6k3JY3zZYfwwsHq63vqHzKHAC+QeAz5bl0E9L
rjaOVIMqY7vRfpjmNaK14GWWwrPTmfeH61XIfeHZAyxEiQFaEfWO4RUfO95J9sMb
wmN8cjqHpNi/INMUmMnbF9ZzGaFsX8/ynwhB2ZdZL7YrZF+0mj95rzvKFm3iUoP1
u9hTGB7cB+x4skru39NYwpS+J4JXMPfeh4quPtCXH5Gur+PnYCElwSPVS7tdRToc
zI0FOo1HBYXivHY4Z7wCMw==
`protect END_PROTECTED
