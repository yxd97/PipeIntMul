`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0wIL1874XYyZPmzGzJtacfwzoHWoKYsSQtAxVXR7A0Lg0Pz7FzzZhlMkl73uOLA/
GOkpSp4G226AvIY1HBF4tinOaJsMrLyWJfezLXAdXjY0RmgwKJB+mlsXWLplzZN2
ecqX7BEYd23BRVaCebBcb8niXn9A0GW/d2rzbTsfCUA6sq5IVcQLr8yGLqJgJgnk
xJ8L9uVEDZqbNNkiPHYtSjM0L6LlJa7UoZ2a7/y2HRf3xTEu4P+Q32VhVeHxO88i
+jSvytIz5Y9S42E2BD0nKszR9JmgMhYuZN01JKAuMsRr2qDlxFwbj3O4TFAvW9Cx
EPmovoMGrTAVR8E8RQiD6qu8m1V8/fsZhsK+Zg2Cz6rH5i5i6km0H34pURHR/8kQ
hU5psH8htnPF3J6dpUBD6E0PFNjhkisHjLVziU7cvD8Qcs5mPaOQP62c1jaccP8j
sX/E29pPluaVMWnjwjaizOhRR9Tm9XXscK38Y/hxERVtjnwLM9lcbdGugdi2pYMY
nQEYpXF+J2RGNOChjtLR8vLB1uRbtTI7/hXhyueX7Bfp0Hn5Hb+4y4l11lhsq1I5
jDwq1I26WYExf88gDdkcSkISqKNVNPDASe/lzX6A/KE4f6Y/At6PdYyP3uPnlqg/
9HPxav0Jkwz/nQAJ9jy/ZKzvSxRFrVnPEtzreYItLCLZP3BfrP4KhzMdMy2UIf9w
u1VeeM4YbVLuoF9cq2UbpQ==
`protect END_PROTECTED
