`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yy9FwsI32NvrIjz3TesUKTS/Gd2hB7zrJuRu0rlKzwb2hNN3WvYC5G9pqCHv7YJ
IJv5egTBYx53blDaz6sccDBMoNkmwkeH7BAaonxvNiY0NGjcD5M52p6DOAPYRt1g
dmnza4pSPovnXRZsjfyMLQ/a7sjUu3l/R3iRrAh2yFZ+xwbh9Ug/fMywfiR7izB1
Xk20flK0fhAlFVNOVEqVDlUS5FQf0ehsZvOBg6K+Hh/wxSYjZ/H8/hO6hStGdvNx
h1U7GICa1NOvhpPiLebXIVSASauT7K7qi2KZn3dD3IJ5oTUjk2mWSUSO8PJmx5BN
E7LPE6BWVliTKxPWQIfFWa9QQ1b2w7eaCgTj81+We+0=
`protect END_PROTECTED
