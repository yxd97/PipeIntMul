`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2sMsy9lt9ozgnaAjTKTI9tc2LmMmxQDcKCEOMgi++TONeavaelKu92tiwwjBzDC6
5Qc6JsOGFW4GrSWuGSZE/3rKJxd6z2Wyskgy77P7HPRzP7P7joIBHb8sCLansoNP
MvWg/uokZRXZxPNYiWZN1k+AkLRswFOyEd2S2EA91ZO0i+WSr/FWSFFI5tIFsAMC
9ehErqD9ARwi7TlLWUSQdicelNLbR2pIxPwgbhvrAj8SCE3YlflijV+J392UTN4D
M5dxcoOK17DXy8qMjk6/kfRCCMnD0hs6AAtW2ZIPQeouD78Ff+AgbUZcOqKOi3FY
qPwtxwmgsgFhYM6Pnqi0FJGpMKuTwFA/d4pqEHpqPC7HdUrHP8BIiiWGG0PS1pM6
4eDdnPEBF+jhs4LDACllcQ==
`protect END_PROTECTED
