`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkxJeu2xRCaH4yVOFi8/jv7g4vHUbn5rxYua6JXnpBJoAThY1rR+aOyLl5rimfoF
QC1gu9BcgCF4QHR7d0skEZpC8Z+6I+Wy+z14GPHA7Mtv/nAPFnBLsQUCC6y5wh9g
QCpIZkALlOQLDNrBz9D/DS1URBUAdpcai/iWCRXQfDRyCfw0oJ2nAwWc198ApAIZ
N+5dCUcG52Xv8WWnP/aBWPBThs0GyHMe68ad7j4Au2E2YmIFNt8pSTxioxb7swHd
Bdft7wr+D3QsTfwr+rdACUT6rElQ82a+7Y4oqoO9W2pHL3xl/nmmOl96g5ukXLAf
TOrFN1z0wiBPs2URZtHEMNNsa0cDT1A7ArshyNa0dDVXxq58Iwrdp+YFw6CVkGTB
GjHwMhIdzdTLG5rFNwVLbzKw7wnij6TXYZ3YKH1R+jr6eJLPIhswMq8W1X0z6JJy
1VK5tcvrImN+XgY25dSMXmaMernxY3ac9K7qfOZICOyMQ0M3qemxJ1Gpir449IWH
9nrlxXGzQrKO++vcEUDozjnoUKCmEUr5bKaDZFqcu0hgtFWIoPnF//uq1QZmc51B
XOvyDHzHqrIoPFO/oVG7ekQ+qmHylFs2KJl4QAmfi/1ro1vQdigJ6lpJRcXX008T
AiuDNbQR0T/O0DBOwdy+7SNWp/41Ssfepfq2YkPuI9bBAiqNbaxEIWTv2w9sF/aU
YnaUKpHSCQMs3bOF/K3vSfNnh1MzjkKHU8gg2GM+GK8LT/EFyW20agy7xdnX8ktI
CDQBVP/gaYlfuDFiV9t7rDzoFt/mRlbazpH5d4VclAJxdCFm3ORrcHNp29GTM1Op
Y5rNp1atqzruXr72ERkDyQl2mKuf1sZP9tQASa7pkZD/w/v50NHxhp3DJW1cnue2
ueIiwzOpntDRIu+CnBdddCGVkDv2sFdbMQRuc9i+acswi34zKnaG4InJlF3OmdLN
K3fvHQC8/+noV0lw/7BAHPbZGHKygOfeEE4+RgsEZ32X678pd/Djs+jam7O7jHYa
6xRSM1hHkvgw7yKzaHcd8TfAlSER5H8A6RWNr5dtwEp7zZ9Suh1DdulNyxLbwQy3
M8CiEQT4BX0Ka4JU+IxfZ0pOO00879P5uo+zxV9Jax7YJdfy8jt16eNb1EpbGmF7
SJPpGZHftUutQ5rekx3KUrUHZbIpF/EoDFmaudpEskTr/Vif+B9VvonRAUoewxbm
JgtDKwpfjnyKQabqvmCKaa/mGo9Y5QJODbz+dFpipW84TtnwHMrKcxYbPSlc0dOX
8kv1ikJNN4vMid+eyCXbCkTs2CO55pb672BO/jREZeWeU7QWgCp7NbZhuWw8b4Uv
`protect END_PROTECTED
