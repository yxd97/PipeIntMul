`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6jIQ6Z9hwK2Ub5Ra/8tlra33ghOmXc62wvnEx2jETfSZtQEH1txy0+D9yagT5Bn
h0URWLXVtZVszAOn0hUOxzhhM8nOOwoWOc0BREC6dAu+ddIA92dojbDb//hOrGp/
Lp6u9qMej0aIExeZ6NzaplAvcQdt3QcFSw7qQ3+id1VBV6GARoS0OeTFT8G2E07q
FGYpsMbQEmv6tpyVv87GJZH8VGpU0KcLkKX+zxsHwjpX2U+LjGrves2YCN8aWiri
Ikh/4oNIU+a2lT0o5rKB3EmfdDnX61tCHHg13p+sc5OHjn3od32drIbO/5BdwYSL
GEFWKfaKwzuSw2PS1kOwYp9VMq3moMHGR5RhQuTlsJDvd53//XV74RRIVTBYbqB5
ndwIuuqNqt8hsY0/79W7vqL7JoYimaEUalhmbidK/+UTxpgyq6IIYHr7I9aQ39Lc
dkoSiUr5tnyr5KefkbZcJA/shD8OGtyvOsOs+8yPafh+o7v3DyY/1jD9ogUozrea
GuJFn1DJ6YZdmB3hoSI2Avub/u/1cKOgjZKCS29vy7IEmyipzE1xTQI2Q/mF6wJQ
0rBpbl5xWjNxfPdpjUDrTtcey0Hhw3axlYzoVdlg1vFktjmQOB1TSMHVOIPJGxhz
q62Pl9IUDNU0FZusdymDwIdPn1ur//rK+Sr7Uqkumbq7BfLiIMk/KpgeAdLsuE58
/AwkE8Ya+ZZlB8ByrOMEQaSLw0WC1Cqsd4H04HjQGvuOVQu9Yrww1usbmiVuwsKW
RO0lQ2WwGuyOiS/aTS3E7u9dJ//7r1w1V/L9gMrKe8FNOekaSfZBG4l+1RP7/J9X
BYFJULbyb9znozutnuFueaLDs9CWkHJEvAGfWMJxV+LqGGb7+AnNcyHqkuswv8lZ
2YwFubJfqQI1r4ayqK1NBQUueVwWhdRPNYw2syF4lEQn0aQM+Srh28K81uf4potU
Lqr01rBiUhPwEmnCuhLOq++/fm45oEiYA9Bvq90YPvIiTx8BPbi8gGgzC1/5Uv6n
FOjFPBDnugqt74ezqBUyRpY97j1hH4nQsmUSoMOMPgUZ6JJ0w5ryceGzjinv5bzS
QT0U+2j70XJHVK7X4ZHMpCtse1np8YwbFFDn/yJAZnQ8qaJt7P5ulEojpHTIug8Z
3lx5qnlyTj1SYllUzObyJ33v42uQhgK0zztwIvsn8lkIZxCFDqt2iBFCs0NjsIFa
lqaVEiS5STQQBSejBd1FM/Tgs2jykebS9qYLF9qJ5V1ZiJwe5u0y3d9203D/yEG0
TzPqTzwbmGcWyaEczdY2UKnD6bqe3sH4tXwXOaryqAGmCvVbvOmY7uOdpMQbrgq0
hcyJhT9NYwgAMptBDiZMEfqz/s0qgEv9kcQ0xuW7SGGcs3QpIOMFl7/7KdcZHxJK
+2+YaA3gV+Derf+LtaiV62kG10F5TYK4v+rXQZLUoQiLUBmYzUZz2PYKRDmFzxEN
V/XzQ6b15oR+cYrseENcMyWWbuAlvk4hadCwUuD0MXNnDXt3ZXeGcPhNRBEE5nYV
Uvsv5eh1389EN1k5DdoF5o8U4gcLo+82hoj7AHtNmbatzirZm3HQt65rG9IhRA64
oWgu40jv95XPlVRjVCmzwkStgV6n3pNMdJvFKgA44QUACUr2+dCHuea4ua7/JOEV
tlZkn8sbayqOLBtOVvq2nY7lzAx+mVVevg/EwD9DvJI24pJL0hIQwB6MHOlKsXba
xyzYt+ZJefQILo8RSMffKl+ooJwLI4D3fCg1JZ/0kpF/Mb7ca8LlWe13jonuCvcP
+99HvNm6y9MiHJPlGeZsNiTtcOyU9hChCwaLosCUIpVUFY/Hex2e3hV5auDUxF0E
vEVWDYD+gWr9w/c3+eDWJwkYunHQ9qITigN74XRxe+Hs0NIZZOk59G/zxnOjnEzW
yxyGRi3f66HlGVkOV1yo3vg6EsOZxTBnYji/OPlxiXTy2YNOMnl7MMzGbiGcaKjF
jJQ71HoEUnlFhZ85/vr1Q0/ZFuz3q7ls/SHodiOsvY/fGxLqH+q6/JqkJRkzI/g/
yEjIOpYeNSwe/BtJj9JSKH1oM7tiOV8EYcwajijgGPpUXmsxCZSGcuV4gZAxAKkN
t5UouLH3TV80PlTOjfcLfcMaQvD7obJy2EcX2/ZT+1dGiICAMMr9rqbQh14WhHA8
lc8SZIRn/vgfhqz7RmY1GuYfq5yM6rCIg0URxmiPoHhIpayHMgW/WpzasO3klBrg
vzfyL69MXSPYbAT5ul6oi+iff7YxokrKbDb8f867CsJHFGp/1oVEPG4398ou6tx1
Q+BZx0q4Z1JmHJ/jGvNHhKMQ9P/n2F74SoZCRxkwg9EwGX3sO0Er8/tA5Ly+eQrh
rKnF4gNKHoPxAP5F/aY8MUGsG6i+vyV9Hh5+l5vS43iVdU0ATxiNd0rua4ZzRBck
F83q4WoqEPAzCsGQMdVdWE10wThaEG2w6a373ZUD76BmG8shr1SydbLflfYAX3Zd
RVum+KkGWYFOITS/19YascFVc4kZEQYw1phmCU7HzDBqot2oT7CgGzco2o1Sofmz
KGYAZAAtjSPkv9+QzuSqACNG/r9KpsIXbWlRzbXhSmHpNS6IWqKGEa9zqVofufoU
LuFBdJQ28VIDhwHnJR13oLo6AG3iSykSjSVsESCb/bkSh3LXqwecdILQfAc6tH8m
98xKUpHx+ItxQaPbGSjkrZTv4abWLlE8qpaqrdlTylLOm+a3TP7XVEiXtzDSXCmL
aHUfLb0QIxZVNpn1f+/+k+NzJ2ITyXXRGKOkH9xnDQvyo758AtNyiFAPy9BNw7Y3
b+tq8Wm1miMtGcwEjPAsiuDhmoxpea9gdDcWYZUJPuRfXMWOvtRAHOktzGeGT3Ag
+XUONeGW6BRmQKQL/2kFs2MtQTO4G1qS2WP+bYOFWTf0hBYCWnR6Vo3hJobMWBPp
DUuQUOroGAcRwQjVas1T/BknI8EO6dHjY/OwhzU+O7ZP67QZsTo0PC6yx80wxOzM
7lKn2GD8nYZNiNZl4QjZXDQY192loyQld9rCxpu9202SdZa1W8R1ur/8QExqg91Y
3I+eKA9pm2bGOv0S0ByvXe4kDyOSIq1rKgx1U41PUixf38ZSeJVrXr5P9MnUsLEM
UQ0BhUYK0XZNk+XYxK5GNjpxg624HD7QT0NK/IPmC8LVCVLgEpJkvHAapa9aJsUp
AGlMtSqS6dzUqyFrRpyQBJK8R1KPavSRKXC7nwYWv4qGHDQwl6Znkxty7X89gb/c
gkITNhkM4HJ/Fpk8J+UlR5Vc3dtf4BeXiWk9FR12J+lzvs+Hm2PQNoOA4APRh62t
1CBOeQRWx53bm6qHKoz2y7gENuMT1VGPsPpDU/TdZhDcBPw3Sy6i1l3ZFTBPdV6M
390TIQdb1ovQYkHOGTbnkuppCioGLpvx0P/gIdndtg9SxF/d1PmshyVBI6RvZaxj
+H9QIBVl0tqv5t3uMzwPyU0lCQ6oRUy/s3wCmOMJHOrZN2ZiodSBb3HX4XaDk+W2
0/rmBf6f/p90k5Hh/2kW+Gg2yott26DUk2PXOSn0kASSTAOrWS/mQu0W/J8F7R+g
wZncWGIdQhh703YW16tFSSKktVOIDusJRa6Fj3GonL0bZ4nUUZOe4XSHEttRZCx9
eom81BxNa5snLWP4b2iefBjqQ2S6dtKMTv6NfwG23i8Mi8fsNrs18F8PDoTSmWcy
sz5NYHYUX2rEoTbRCNJZhP4HVkJgzo8joh858cUkq24o8bUpNjMt3r6OxJuJ4HG2
9HgdPUmeWUes5phFvRi7x7YnRxS7e1Ja6TE7wz5IvCypic9T5pVPa2qZm9wCh9Hf
kZJB/0B3TRdd47XtvF2wGJH1Xn1JPhk5+fnjgpnBODAI+3fdHYUtTfuGrDGxGinE
isRqvLVSJMReSppnQ94+dnWGGumAVBsT5RLLtSo+j6JRqzjCzIvx0BQJsK4T0usa
qBIVQr9lhb/dMH40axHwbJiRMF5nOc5FCkrLkXzFbOg7asXpH2VlI8XGh/bXBcyG
C4kNxJPogo0go56iaziW2snZScX8qlw52A8tHbxukvoWzcygcKyYiGNLonpdKFHu
28MOyAWgEAAsB34LfDYKrYpg9ezoFZ7Wh06ecXr2u/kyTs0WY5Al7bj2CBcG4WsN
ZIwIdjDofcQYrKm89rNB1WRKkheAOJH0OmSl/zpTD/llF7pR9zl4aFCRh7JSdO1/
5X2Fo8JCyqg/7vIZjfwm9CWojUeco1VsrycIERA0EDrksyj+4aP+Yg/m9LPGkDgQ
ZQssmiSE+HBlFvl7DiTIv7RpISYv30LgtzksJsL1nH7+OL6RCmCNtAYiRbCNMStQ
fF4saQkZpFUb1JIhJ5toge86KQdMh3HM+B612c5BildOolofRchN23W8d+Ms9nS1
Rt79NhJTjMUyDWlJYyJpGOxz6Ll/+v1SMNLIu829mm3tDWHdpkguODcG8jTdxHoG
80/2dsXOltVgaWXMfE8RgbLcDn4SzaiZyC/TVFPHD2Sdmd+h1gLgF11AGSCS8asM
y6bYHl5/FLM7qEcOUxhVA88bu4R7AGAGvABEsgxOD3I+QuJPH/CZ5jf0syUNSt5l
S2CqFUZ3bZG/eCA+3fF6ZkY28b3MjZyVPd9KMRJKq9Mc+YBG8uhPIhgaIm7JMRY4
H5Di6hHLOh3KWMSbiFmDdrqEloh1bmgtNn7ssq3YIyuAbV/yW3NIwolxD+PeFqx0
W6W2m+UfjHvU13Qt+s4ZzaOiBbkDWV0F6wULkIJpI72XNQbOeZW6aO8NliQcndbj
FTlq8frPi4Xytq7UWAdtEISaVVzGec317X8iJd9y7oQ4SknFOk0+64HRtsA/iM1B
nE4CsCD0umMVfgVs2Tk7f/VnGdD3398LE222ecZSgIJLQBwImY+/qHkl6T6pDkcU
24O2E/+cCDOIhjqLhUPFMXEzOGUUJN8Ru2C+SsIhYsWdepQi8yDjNp2E0H7HSTCF
ewF4b+F/q4NEmfoQLIViPH5iZTTvcs9Uko8RlaSWSkb8HKksI0ghfeX7NDFIgniN
zmCOpvr7NiWDGEm7F0VjIMXl/R123AqsO30MLcINGW5pHy3CgphipnILh/sNYF0L
UmoiV7alhFCwTbSgL/Kiq2p5ewSYbb+FGgLwNc0Ul33rTpxKgRmDF7SzzaUxMpJ6
m6jQUnhr/ROpZf5C6v+0JZBXfBr0tbiI/71mvFSEcAjL6I04zpsOSXlmmEvlZgFg
C7CSKFbn0rjvHrHWMusfqQ68nKDCPXcly/hwJlFmGAq7SFH9CpPrbTqAvYtJfnqt
NuaNt5GCMsKSFgZ3Ry4PfFM1vZBUrGs1/ajq/Ql5mkOnY9MzaGXsW+Zi9YKOjqQr
83/sghR4UEeZ0HL9y9sVv34IaoAXhde8h1l6ueZHPc/6ejGGTx7UiQJx2OkdPpiu
TYRQ8lvW//Ouj0d9O6wfkebAeSLURNDvGoONfZTLqIr4IHRLy1b0mFEIWTQ3NphB
nIbenpJLGe0sGsqS6QwimbmyGCIAnrPRAFgW0X4IjZPtQcVnZC1VjTjjHz7fssi6
P11FSXY/R/rPKrA03jv8GiXHim/OZDQiQ5L6BXQoA+HNmqQ0A6GHCFlFQquvuZ5/
f/3mI6YWgVNp0i+0pEEugrr4JIWspNNmxcTXToJiao+Smy2FSQLaP2Xr1qSnugfW
cgo39183H0E7cF6667LlSzr0BELxVMAp2+7ZZx4772ndhEW+BFiFc+gPoV8nXk/t
ZEJ5ejJ1usbJMhnxEfCvqcMaBreF1MTmgL/l8MSjiMJD3uwIEOWGbqnK+kfMlCwl
USz16/oeMeynOiLNzPqgXkLaIi9KPRFJC8t5Brtcz4XdSzgpvoJgUSsXdfPU/MkL
t7hgPn5bGmDQa4DBO3rNq/ox6GB1Pvl8zH103y6wED9xIWhTE7t63msYYePCMfjD
dimN7fCUde+HmFtM9c9UpSo9uYTcDL/J+Zb4aLopog2ZWo8mm5T2KsPIQkcWWVvd
mZD3hDbwl1PEEHhoj0+PhyeOXW3LAzGA3eqy/tI1pIVvIQQ3j4+pWBcpoRbCRqgS
72ragtPOM2mTEOXJvpzbx+hfqMlXTsWBKAk1m9Xp2UMHhD94wpoH1JIIEN7wVlFQ
YweyrIftNGx3VSJCbCy031MEmLA9hRMaTKTicNIpORHPWxMn+eA8xm+CoOemRlto
NMHfiQPfqiIxDfbKe1eMfmkfftIfGwhDxcnzPpjs2QhuJRYHYdCBPsLVC2bg7ygz
On6XQmh1TBzcPJPib8Uku+maot7WY51eTL9QNcGCw94yIrTUbRSUkt6sydqcwtmU
4bCDwK8CTTh9qWQHSOjUWfjf9aG5GJPXmGWYO3INfOPFT6UoI8Qe/qbzyck0B7hx
bO9U81aTfh75mxvJT/LaMXJ51gPE3WxugsHZh1UC982BF8WDgijiMyoyOYakwisp
fGA4wlwEn9tcp7n4sBSsB0aVJJopTtOx7HXTScbbfmRh4m8K605JX+9BL3AQJedy
4LzMI+SY5Os5TFr1ivYXsHJMdLLcGBRg2yEoo4lUyg4S4VKPKeX5OUyywlVAuAWw
Orf+9rQNv1GaT92f10vuNier+e8zgMzmb0gQXdBKqn12ubX52K4TxkP6vzwfO29d
faYvdM2ScPoDJKwQn36eW17Vq5eWHLaBFz5f3xmQ0cUlm6Fk5Tpm61J5M9RXT9qf
fI3R82lUKWIfGN/iC4AwdlIcBinQnXakrItAn7q/XkLgVdrU+fFZRGbUjNhKAAYP
Ew9WSjFY5ZuvBGkin6QidzxZ4WfvSTpmM57Xw8E6jPnVR8bQju1m2fO30hdn2eQg
9OoY0cWhvnH55lcYJYeRLaCWuawZja3+BbaszGgPdk5r+XTpGxk0+luGprjPYqc4
MHT1/vKeGYvWoiqm+UJgveNmS+V1rD7znpbAcLWXdfc7SU+/P8tkhiogt7ybjyN/
LXKH495G2t1+eevP4YeOUE8+E4FdBxwAV1wIHtnvFRfModFSQLRUCb36rS3E1rki
6JRKZeXMXNODcJM5RO/T2NTmDhwdiPDcasHnuEhphyUgwQH36mwawgLN4u5jVbPm
h6Phed+mDfpJJuhENRe2j6I6TkZBPXT/zlA9tOfE9Ff+xxlcFhnI6ogYRNLkonx8
VhrzKHxF9DfSJenigCEWIUVRdqDEOoUgHfVlCdDWiuz2qTWQ0WbZEhQ4WrOYTwCC
4eauAmchDqqSGV/nEX7UbTSoxE6BvP1UvNBvsol3IztGmbTW6saBpXgikxKVtFHl
hVKa1KRd3C4zfAN01LKnh13O+DZ88uc/sXz5bvLcbyFM40/0PYInm6DJsVnY98le
Vb/dW4jD6oaMBzGdOc41d8dCGa5Fzb5U0of6NsS9k/t2pbg0rXwhKVBEboF5jigk
X++dOouo65DXp+0BWu1zel4iDcVsRkspDfbA5iJNwva9YdsrClTPK/p35YCVrrP4
JjHTvEzYn312mK4xY/DnlUxGCegeFzRm3F1hW/ehSUB0Q55WKKggBbbUmG1orpp0
JcE5o1OfNvR6jo3ug32FSfjmXO0ch6aRa2WHTKPiJpAOMy5dsMITWj6wGO/zK7yM
9UtYIE4FDg7Z51Ph3vBHCBuC4vgW6E8s1AN1St6Av+T1aJ13+X+qv9CET872lMnM
t/9TLhLCKKJS/xQYGt2wRQgjKL/wJy7kr6srInc5sx8JfCZ+b9mkfKRGx1gd5IgL
ZCSF8JvhPZOZ5jbDH05+xIMatFPWfT5wTTM4cf/Y8B44yQd8ewYdnrwaAWcGoKOT
MWaKLgF+arhDm/AxXcbe9LVSBf8v0qE2NhhwbJaBcnqvgNXsBnXDrL0SDdy6jN0t
Bbk0pjQS1adUVYf7ci88Oe2y52oRkpvAX9S0PnRAzg1bE8WzLi4oVep8+xP5hvpN
PmTh1WW/239/us65IkCVZk9hBnXHdlzwcvNop57M5Xg/mRj4zn7JhT3lOA8/5jzL
LCbwGMRdeHzo48wWO3A0kBs3V7BTs0Q0nbQH0rrpdkvE0xGPsVi2JZBIpnk/TJxW
x8glG0VpvWR1kHCiZsFGGroS4DiFUwa6wTquYRt7csQJBCpsVC/HHz4Xf4NzZHIn
EEtCBRO7Qw2TjxWVCzfB1+tKhFmBljKzcrPa02OIgWHpVN98hAlzFHJyy15Z9eYx
3l1mXae8FS3Ji1230qu0ag4ugi5pTD12hEYXkfxjjlBro27HZvaUxO2xfnAFIVFl
5pZVuWH7wquaDiVKC9vHlU3XIqSi/OuoPcCToWTXPzw3Ltz3fqFBgQ+wHEvy9o9k
Z8Tx/hoDJA5kItyYU4sH9XRkojwXEXYFkk6Hu2zNpIwX3/sa9pJCwQQLt6B1MBEQ
UvJtBWx4jMvV1PPsaIT95jSoj8QsK9QYe+ShNoODO4eB7s+Dxwvq4N0s6f3VyeuV
tmgdqJ1zC1gWiaCuC8Ws/ijNSrqkcQ3UOEc+EpJcsaO7jGzk7nDUvgo7ntFwM/tX
hJx/OWePe7oQJGwvSHYEORIQJdP+SAQ9vcBnX3BqQ0QUQOYla/TrSF7F++lY1Eyd
5L8ZOLO1EwVsB9mLtbOZwijySdgO07ZNVV1M3D7ZNubHPV75l6O9h4l2DRGetmqS
jm1+NJyZi/u/ClhIqwtx7HG/d59uAAS1wZgb8Nq+LuBmMHHt1kN/kcmff2t8ZHux
1A60iN4UNjeROaiAeQ8DazkQ1nyRl7lzAY3dTqiEyG1mJzZtvOJQm8sakSZG2/jk
FwBbS9vc54peZOLuKHBz3SKTdN6bcyNS/IVUhe7vkoK5PRQJxw8UpdlRbb7lXfZS
1foZbnOQ/Ei1NBdZGzYKrXVJzrfNjvlaoVOr4TGDcoI8Kgn0yFPlBwIuQd6UVkvd
PzCvn2IFjxw3kV/wbwp62avo1WnmPPLU6b1W6p2iJ4gFAe8W5a6umJVLeVn415lF
huqSm0b9+jpNCUvsSgLbJOo0lr5kX+WU6xtA+Nfbb8KFQls74CF68CupCtkuZWEz
upWehcnh9r8+1wBnlyTsobSoqgeSqFbkI4KHgn11Kdhc+FHOMnRfAuUkyPEcL7Tk
1LJXPvarVLKL3AzROEuRHbjow0gIoW93GJy/WH0Am1nAa4whua151hAPKmVLrop+
/wdz/lj6ZLcL+vgRoBg6U/qdWN8ZqtHT+rDpb4s9qzoQBSw9y0KID+aKescKXc8f
mtNDUHnQiLBrC9/TW1Qwzq8myL5zMVEokzxFzdKWiK4Ie5HsPQPM85HlzAArZk+t
MsvK0PnbbXrJaNbLkb8tC2gK+xJ4ATjKTPD6LJarQ4Z4QRVWBmBLV43V+phTrOn7
hSIfPl/083AWnkGf8kXU8OlFZEqGjCFlBGOD43GXLcpfB4rySJEwF+iJ5BGbSm2y
M4I3A9jGqAOXKr/vDkoVjHFl+LVRYJATlXH1gCnPNYpvWN7dcb8WxooAgWR1vGS9
Ckd3qbLqu7voWCkoAsw2BDMDrc9470xBftAFOafBNsu59mRzPw2rjCv8RlzWtK0s
8Tgv1sozfnGR2QTgoVDbngyd+jR0cjPl8cK8ZjluWmsmKIWPLfGXlnR1XftpBiYA
CxpiKNhdV6r2TdUDRb5dsXupQZ6V77NFQixuvfPq8dPrIIFQ/1jmzAgLQGqjxRYy
SwLpOnttklx7xkSZLpG0wIRTjBsqPw0/A508SFPQKtiMa3XZ0ALKwHfIvmyPX2PW
tnWsTJgJsu5yA4ob2kHcoSz1NPDOj1rNYe2FErWoB1dxgGsuK/D18f7WiGwIMbXI
Uaz3qorm5miuvWbGx6Icqh/E+2SqgL5UBYaY68l2qfXXAqtLV7O2FEO36nyvfTKy
udGYX+wZ/uyIEV9/0vk1nM2xMdc4dtKIdjZyxlhWFmJgaAAhdtmqzNcJTtSMMl95
k+GCBT/0gtynrHh180/UfmwuDlF9SSYLxo0m+ZJxt6BIjz51THeJnnwNF0XGflq9
yYwWkh1B8VQ+7766zo661DG8UpoTdfD4UdK8FB/xywkDGGn9iuLTAXLX2LslSu1F
oz3ld7NB1Em+fU7g8ptjLTYo4PYveSnSgh4/Go2CdxFnhUuzCThsutBgyJ+O1V3t
gVftO44Bc+JrYd1A2kOYoGdG4MzzKAnPjvOw+Q7zwceVt7hQ4LjmJPRbEgODFzj+
kw+AOQ3pbVG8Ljtiknuyd7lbu5lQnRuu8hy9sjnRZ8TIK+oLc0KKbrSN6q0l1l3I
fJYvxJ/rRcBDNC8g2o48Mrc+lCiO/EvPAKGsmhVbsfWn03u3gcoHi2RFWNT6hNVF
Oknj+Xdx7zFgFn+os+0aD5QafzI4herNwhbIGJnkdRCmSKIMtHFQ3ibWMug8EU4D
yjJPrV3SXqwZw0/Tnsblq21oulYMiJqc+M0Scq4dBQSt07imOiePobkcgq7ExeIo
4uKPPUA0Rt5BtgZ7fiOiZa3/XeTqmGKO+eGT81BlXuClPgxh646Di62rTG98Gwit
2l4edvau0Hc8lUboHveFDzgFAde+nToUlDmwvGxJH3ZRJ7By+BO8rdFB6oHvEMKr
IxEpXwbXzkcCB12XHiy8JSMa3hBaIWUvATmNi3n0jlCW9Rj94o7+Clzw2R9MYGRn
ZkSzTsRIIK4nn16hh38dCSoe65RJEgS+QdhOAbjiNpL/xNeXJEz4AZ+yIMbbXuP5
YKOThY3f1mWUx60ezYpdi/MkU/+eZUlmd/IQP0f/PH2lMdjFyDVfklT1t249FP1e
YGZE2CYCXjdMF8z/llHLyq0A0St8JwPMvCaTItpz1c3sGsSmN/1QtgXEJ7ZAmIGP
E4JTQ/3M6OgLaxOsPt9HIBw9peDdIfNeuBLT+WBdSfhDAVdSMGnG1K5geMfyxC7q
6E7OPGGuUDvq2DFUQUVj+iHjKdyoFD95Mb248dywqA4Fwo4thgsgveV23Lm2lE1o
vEN0UFM5+MiiVuahFh5J4tKWBLb2V6+bzLJtR61wa9AAVKVI00KTSFg7wFma31Im
kgeNSzM2mdGPCk4vZFEDC6JtXc6JthnzVHA5SlocEcFTD9bVhEaRqs/n1lrWIBJ5
89U4pee6Hr3iwvQN1Ye2OgysFFQGsoZX0eT16qzA3APDp1fPCCXiCrpepivRxmmq
lmQxqMowsUttfu63MHaAW3ADOvmjbXP0i5j63arYdfCYANsj2EQxmo9luAkiSiTN
SfewRcBxq3ILRQ1qJy89JcONQO5eY/o69+Og+1tiJctcoJScbhoPz318a4qL/DyX
HT4kRsq3tT41FwzOF1YhXSuK7W4/xtrMTbvXTgBwdBOEAchySVJlzoXWkNj0fLW9
uytbgD6i88kIP9zK4uL5IOTeaMYjV5uZvtb7iXCzV55n/D5iSvMPLM0g64EndrRu
i3wB4IVjZBtC9Fr/LseC5W7P4u7pDNZELjG8JHvlpvrMwQNdNWEEn1aNThzu4/Tg
KfdQyQu93UDWzZd6ytbZjpxABXhsKgLniHcCuI79VBPI/R2Z41c13QNN93dnvC2o
sl27JyYxTzhNEx9HTlVyQxriygjD03LJ+NtUm5gU0LyJQVShf7xtyPmYlmzPXJ8z
g7qHUjG6tLQ4zlDkkkHGUFmQH+7MEep3+R3TVHKqD0+s3LEmD0zcppmeURqr5Ocy
1bf9BgaXfXCoHzFDBT5fj7JiECJijfR1TCCdDvzkt2JeK8rW7wKd4Tyx/PWybTcR
dxWcR0Gbew4IwMmHpzATILMXyZF9awja7TAwjFLZmu01jQAj2uu6FtjJ2hbIVmss
+yiYhg35jJUOh6CNt0gAhY/GJ5hAlpgEecVO1FbmwbhSU2kRLFidvbYtL+xUFzXW
ERMOrfL0A/fa4zzPtfndE7sfncs3ENglySnmEgN7wQPuqam3uVfZm1iuBTaGcfPM
d7oEuMVzwF9nSaGiYzyoooEsDzh8nITK+w8Q5pNIBe2Je7cV4lehTL32/RyT0OUg
XAjtfXzAcfe6pADWETKYHOTMfaf3F8O62YvoN4xMpADVLPs468MCd8ep+deor1Es
sLNJpbIhHLGAFCorAfkiaqlI8gTmNwbgzqdFXwvcd85xzQcANwtXfvSHLPEWTZbB
0bbwLwSRcQFgAVnsDzgxx6Y/+w2Wy5+dx65yX0+eIQmxvNc9BTmkvia/nwbAIBMl
nx45avkOCsGv7Pvz3lP83fxXGw+LWjGRhM2IhYkEMolb78GuarZu8U00lbmDJLNI
ylkIUMqdy8hjYisur5L8s26OxVoIvgqTLTC12MTIw05kpS8g7VfZVwvfspzgCz24
fTZvRmYKDSx6B3VFKGsZ0LSrTgolX1HzJjruj3hWJsFhZm+IpnbWCg7WYqfAiyd8
Ma2guakQFxfWoQWwQq4R4Wr9xza4L20Dt21UdvNADomB8eqzmmEa+ak74aa2v7iI
h2nm4jD9Oa8ODNG2PMZLjHlNdy9/2HH+qFZn9AWz/EogvGEot547V7FpeILKJ3bL
j9HdKDDzsLOI9/R4wgmekCahRoeDSAp6keeYTi/Ab7NaEe8VaRZ7jleVHPkeWMkO
kecbhdtMByPnXm59VKz37fErWdKF8Qehjx7vi9OkhtUGDitWRz9NWfKTUXYrlfg7
aACdsq+KqILDv9gIKy1zbStr+gnLYYCeGK1Jv1pFlMYQllnUZERI+H5R0wltN32d
1ot3Uqqr5Va9avfb0B5NmBmftHUmyNNlFmiQKa9McJY6r65ZygeEs8Rl+AfN/4Fc
5G3Tpr9ZkF1JxxmIx8aDTaz8vQF2EK0eNQ5YQhxsBoit/+CE1MNPoOaPl74mBqDl
8ER6T+Lv2aJlHLS+bRQj9cG2kA71+S8JmpkZvdTxCkyAnwklycQXh2ZaT+JjfivB
K44I6osW4aflss6dN+9+1ZIkF/geRWQ500aAbA3tFECdjTHXa2s2mhasOdm9x/8I
bWgXmTQjCITeiTPlrcjat9T3N+wo5JMz5tE/ZNctj8XQtazhS3LpjjZMa433RfQm
R8HSE3qg/LZYio/Tgq9XStirPIHSDbfNS4Q0U/VlUSXhYUzL2FQF/cnVranwLJg3
+iYuaJHiYJt7DFDwcNZHjkYAqd2WWFaNZEV/MmsrFNc3kif4ynGPLH0mf4Ssdn/+
gtK4lZI1y8vMtCXpfkO467ci3jhE+8daBOzuSxj2uxK1BbLYCvQ8um++VgjuPjHO
ROjZhV9SPTwkapER3O7FKpc5L+8HZq0jqyS/wpUKROVAs7FXW71UKnTTF403fBge
r7x7ykJcZl/ut56PZ+V5MXtrHTNu7y23CD+i0Qzq9wAaNKnGeeVPolEkIewSX9i0
U2bfFNoOzXOBDKpzKrwL71thXGnbiHtSYcmppc7D58qFB3QgNmiPO5P/EH9gvjen
KoRVTZjLiYHMPbMfDmgsInZ4wBuaT0KqcZyNvBO+vAVv8T0bFPNHYkcc0+LrVgQn
biPZy0/lU3WnNsxFvKHB2wZJrOAY4AhpUzgaDGXIpg9Tn5bu0IKllMiJ+VJhaRXC
9U7RcxomSg3UDOT+fQgD77vwkHEMPMkApmTGTVkQ02XpBJmTaRBL8cMme344sSz9
caLtHWd3E3tkyBMrDEtnYCaGiYbx18LeazWHbBI0dHzZgp16tBRWlMiy87NjBX6J
e23yiKz/ZG4m0DARQSbZI2rKW/8R4ewsnTNWfj60N7bDJ+5qjcF4ZIpyP2zkgvgX
6yF895BpK2wjsrjM4jEqC33MaecCMWIvW8GfK+bb7PnJRyaaIr5HCd6R8WVbIh9p
Vyzap8KUWNlGCF6hkrQ0pvt1UpOi1BYE41VL5GdEgxVk0gv+zDrclQ9ZhjZQojXr
OLWi3Q3tdxDDCLmiDgXhnicWgWEOfW4P9/W/N5d1rkueW3yPzdxcAno0O5vvRcNh
lPRR6CDQR5yz7JUByyQULCqZSSNVFMpNyhD5M9qG7iHCQzOalzWrPehawN6vaAX6
BcEAO4tDOYfziGtg/MfErHvOogJ/X4UiYo1v8EpXQktVmQ2LYzp+AtNKN3n4/W4Z
ng39fs/Aw5Lf2uBtwQ2NLKPfxYtbEEoWjtcXa+PLo/X3Cu6Hx+0ER/WBmweKJYZE
rZXK9b68DAGyXU5DyhlAQ1wlj0snMqctZL9b8hgtWI09Gh5PfFES8dqwus9DVEe6
9CrV74zq64s5/2mr5VS/Rhsb1x0gvrWGEcLUZC1H9mVRqQyV978BRwfM3VIcU0Vc
JWpLvhqQpfVnnVczEtFI5XAiLLJYRMaOXUlA9VhO947N9K3rg5rzrY29fYFTWxTe
4OIoamk/DXortVmivyjAEfvXORKpBcmhdyMC/N9h3QAclXZ5HOD9QqE0YfSwkOnd
wXL6scMRSlp9yI8rBXLOLr19SwDBDxZSILzXnb0W2ycZM60NX33iSaxNs31SXT5z
1gK9xIcbF3OOnh0Mz+ITTr9ImduIYv3Ku4D/wFmM6/S9qJLjP5Gts+hYP9BXTmWY
CyQvhe/WKTcBaFsc2s/Trw6wpfUPMR8FYtVVrn4Eo6mSzckAWrs1ZkCYa6IGhRTs
5fWHVa0STy/Eot4tVFJwIqDZxT3cTzsOEfh7U7ws2vF3z1r8BZ6wOhAd1dglZ3y8
x+r6Q2r2dZZoMiMLRUUnw9jagXnsmlFtuIun1CJNgUFWU2owd2/gWlD61tvltHOa
Z2qpezMdFSR6/c62vZO4LlOIYfx0zpskrcJIaoK9GrT7qaDmUJg9YTZFxkbk1Ohp
rwuhF2sjMPIWR79/aIGJSEf0s/2iMLbPNTpx5BgK9bgxr8F+3LOW6TQ6AIBe0Dx6
VJ+MxXhETrAS05EjlVe9MCtgvv0hBzpR1+3I/2VJOVm4V8xFy+24pJMnpGe7B96/
EFbfxTbVhGMMkLfjh46t85dEeB9YDkKo/wuCweaolqk3FfYPhqFmPZhpgsdKJjjs
foOw1qgOIo3nYshpgFc8QXDVtAE73m5RJBJ+rby0d9YSjHalKOfT6TFcbxUI9yWn
G+g5QYBF4A53IcsT2TX7DRhT/sHdIplUnMWgYqY5I4TN0exm4zqEdQY9r9t6MPq7
f96omWqEU7hL3F1xrhubN1IoM7agKRczJIMy71+zJMt/NrzKZaBjjlgdZtN5FdQ7
HMqLYdQIZlxyeP5JepfRq7FcCy1joZJr8l/hRqBZKpAHwaMkgeEMWdVExosZ8Bzc
CEO1lKDZzcqY/O4K/SlA/9mqQ52/kyPpX5DeUqTbtMAXTYq5KfWUMuThv7gFTD/U
zGDSutFIxaOp0NxkhFUtDR8lImod3BCkNJnNHsTOQ5/HREnJReGWi1Zbjo+dv7+C
GMWOnc4kGsN3hNrQWx9cCrVbyAOoFerziwko712xv+mzeIvnw9fGYAsCFgnxKOmO
FVmvrzo3aQwSgM0nnCRydikXeEkqa2of/FtJ9TxgjdF8CGt9nANg8t60sBof6Ska
84azTzaIMuJsCRUdK1X887yh7JQXxe3D5h9LhdbChLI6UY1iOb0PLDJs+IjDK1hR
QJaA6TKDLJjhjvbJhsAiB+8h3KBawSch4dOfzhUED06ToqhnPtmnkgdIc8cWoZMS
OxFRI3kLNpA4x8XHi4hasK6sRRNu4P+fq9z/DRfVplzhDg1IQ9UL3fZL6RBtOg9h
ALl8HMqIT7gUgV67Nel5jjX7OLbRF9v7LNQnpmtKdnqojaYW36eSoWoxwveNOiAy
SVRFTFkSVNvGdMZ7VrztHwwxEkyqNw/6PxIyJ+GMLXmKy6OM4WrsihanZutsiiy5
PHVu5hc5Bd4MI8P1Q75TGOxy4mV7EXO4yFq3vPsduU4PPyrHmr75fiTgyjZVP4SQ
BHh2Ct+q4Awvvd7lmfacvbUpsGEVAMnKPKmGzaN40/VmbFt1qmM++YT194AaLHs+
mc5VLrlkxOmMAsLdSt4wLIynLzui5XrbE6PZufYDneq2nyHJzwHDXsH+/nX+/qaK
PT28ayC0srht6hXew0RTKMcByPuP6yuHNuOOWC6+XCckNrVGgCVBEGMgR7ATRTsO
rzO9//MNMGRAdfWycN2x4KLh+uPGp8lSDRlfT3pCJK8Uk2GGmf4xwlCUiFr85q59
XffkZ4lM2sPajPZ5q081+hk3vKXsPY0SwDCuH+VJGQYtMgx1N2lIq1d99ANEWmkd
GVbCHImhYhXoJ4M6KxuLM63GMatFfNWTemMl3VkS0ld91bYbZwtmRSMClf/j/sHR
2KProqodFRSRkGevhW+OvYHhpDdfK7SWi1j/szfEm1G/rq+zZ/uZ9PGhH1Zn5kzW
KikPVfYnYGYzBOlKwvtwaqAzxECG1VozA6AoquLkHcyuoedSdMDNvyT8sa3HZnPn
8t74N62YNMZ1g+e+Y0DYf6KnFSMJvlDkUB3OCk28TyhbeRzKskkqe3NJ6PvMlbGr
lo35jB3abWNUeNMfjNhykpF5WHSmECfF7EQUZ25OHv9igC+AABl1nayj2NSRsptu
9+9momPrzHDfAaJArn2qzHVOL017RZjjgJC3ZCS0tRxXAgrBTBvEBVIJVG1wR6od
gwTpRANH2CfjIu3QcL+hV2ygYG77E7lNFMnvrNpLNwjQKReVX9HJXvExSNsJ7TCy
SBLa1x3Q+h4FBec8c/+y8a03ynxDQtCXKmbndzNoMNr4iu+kZldN2CiYmGanaT7H
yh3c8DwYKnBMp1UWmLEQwEmug5f8w4Rhu1t0C7s/NZx/XzWKhI8bs4iIxkvQDG1y
CdAN46UeCf0aZ/YAt7EEYR+Vre7m/d/LRo871L8MKryHmfm4LtFXX8PuCnBgAlkv
UZ9REYqaPgnYyTrqDtGcQ7l+9qxSAx2xNs7oBInpFiNEq7t9/fRyx3hZAdB3XWNB
/7FNpQIQBXN/wcx9ck/bpDr0swaPPAIxNp/2u8UzxppD+FGYh9yLPRwwhDdNCSXR
2yazaZVohhTkobGj3x7f4WYr5YAnEo3k0zTAp4j81ZgPYpy3iV4hXNCjCfF/tet0
aDIRetq/ioGe1+6Zm5gSkMUJnc8Sk03WgW0HROX+pARebTueOLxpIp2rrF/UMGkk
h6Kyh/QTYERAAUMfq4wkh+WwazU6muKbV5y8rpKPQzb0JL2TZSwPSX+PVlkWZMDi
gdsy/3vWOHQSoGFUtTD6esrB1Xm/h/u2NOamyFmetNs67L1bAGlY5fFz+coPMlHZ
NRzTQCjqdQ88VIQ3F/XDOXZJ4frMjjdH8WsX1DfWICELxA6GbqQOVguXdGoCp3/9
gKytlbmZbrMZAoYK4///m2PCRizZeaBFrQW4h02V81WkIilvodR2+qRUcwQKL8XZ
GfSsiPTJiMQEX6WKakMWA12n+GDWZvR39MAyyYs7ghG3R9dFwS3SAChYG4cC6ZQr
KL1/uF2Qew4kdwY/FIdBetIikJYRbjKiWYmoW8gUH+/S+mNL/ZSOL3umk6fJQUWm
GV4YsBw9y/wKNZ5Em+7OSX/Xp8cPrNBWJlXGZMRQjutKhe6mO0KzB6rfX2kzIsRz
4IW1aXeeKJhPh0Jl+vkjwKJiMNEInaEvIC3xkfNFhgqv4pVs9Av4ggl3nSjWbP6J
GAUJMVEcyc91LKLFuvzERbx2xjlRiueA84nAi0OMqORexpyO91Pa9HU3mbyf4DlZ
Eja0PzRac4PUXbgRYpBgFOIHs/qJvLq0Dm7+HNY8YDEaJgKhe+42xUaFcVez7wNz
w3Ts69iOrFnEzcpgIC0PSG1eDdo3vlUC5c95eLcb133jmkm4nUk5bTDC4lVDxmYx
cEartO6SVnJF/YIdlV7NlbQxUGZW0SKwqXwhBY7Xq2zFTR07zDCyNOce3EJfI88C
C97SsnVfbCVA9zMg+0wI/70Ml5ZuYvHvi+TSrKkJmwVVOBi1AXQ5yJkR9T3cR6hu
l7/X7eIdrrvMr+3nSHa/wQYbM670EYnWE7VcBIp20LHRPTB33tJXO5o+lvHUazoX
xlWpmF8o+p0y3fxIRnIGDUy1AEWFVmWwLy8G7T3bMgnJJsEsyv9VxwOIxmi6jzvw
oApTYLfGdeBo3DuCG6Em0FrGcNNW7wH4thsfjk+OLuSvlVNLbhwvpOEFpTc8YO3E
cLAnXp3OSfjEvFTZB3p8OvqyuWGtVLxQuwXcBORaSNDnQ0W8CMfr/4p+JVNI4/E3
IhX3qMHsYjr7eQkgYPrvWIqgDbNPlHieT5yUsw1UyQBy6jACtLC/MOyTexgO7qxd
ea7+OtmWubiPLnQf1Rcqdt1YrR6PrTD3fSdqrCAyYAwNWHoo2sU7FP2b/NeipJFt
0btTCkPK7KbxVS/dnf1rT0W3TBIOZ029mptTDfqK3PLybI+I5UFicixV/lcBk3Cw
UON6EiFecVegqjFRxNa47P6zoynbgsajSZ2qkpVLbE1xxilQHVsNSuNu+VLO0IOF
Mjs3I6kQ0IMzcxMXzTl13rot+wApAr2CfiKClrYGp3OfgSLYkYCtfJ4SLGFt+1x1
exdz9n1fNcivvLfRQO/X0D7kw4gXmfF8FgxGQwKEGxeNj1sk7oh78+A+X941W+JA
pHFW+eYk1+semCmstzhTHNk0LZT3lL/EFTph9BsPLkjox3/PXMTu6pw2+mEqIW5p
6PqCVfOWiFPPCZTnVVzdWTY2L37gwECu9A932ELKLtb/EyLRppJhkoXyAR9OyxXu
by+UgcbX8JQS/EEnDxHYQ5V2Rozx65LE4orIXS4fBXOrlxADmFUxUQ6qCFqWsJpn
axlzZQaDlbtNeYEHQYdrM4oBUyPpWurv20sLBl61dZrFA/osVrBe3xP4MQChQnwS
go2vkHGx3bE+0kUejhBE2/qx5EstUjEW5CKh7n3BzaD9B+Tg/e0+zen2jbETYU91
Bs/owkJG0eHm2Yda2+JNIlq2QBnIWGTES3G499dgiWxKdrjlVa7epXPKk8tNJdYv
OSGRYfMs5ddnu83AazTM3Z3GKYvYBVcDw2xsy+fRL1bvk8zeb2aUj1aq3/aeaFNh
UudHOfBd+wmpDu09SgQsyCBeZU9SyvreumcY0nC6Id7uz6XrQmbwfz2LcXvQxphf
4/XGnqohTpsziJQ3LzX6txREcHLRXa9gtNxqyhKttEWJm8Ad+Gru4u902KAM8Q97
uTOVXDhuJsfTcaYECcfAz6MYnq0idjumvFaRIMZZMD7P3Q5MuZvZVtV++xz32mEx
pG+MDEN34EQ7aIFSf5XjHKEFS/TwpZzhcItxdg45ZfDuxXGB1SvJ1RgLHBjggBA3
VL1t7Q4g9LKUm7+tRDDCsXIudTkBQVeEqeIrEhd3xM2kvMvEr/UDIcOSLHcpj06P
591rPftBYL3bwPG3/f/tv3ybj7khh4ntyECJ1IfVgfUZZuhGx1MkREizw4opdgiZ
IyitOVL6Lpn6Sz1Sui9VzO99zKKVwFwWLqNMWx3rh+/A5iqK2ywNfUD4wlx04AmB
QQulXI8eWSmDq4jEADcAxkCWUmFwDsrpoAfxA4LO8IBQjHdzFVZyOOU0ca7phyAY
EDklkG5PCmZ5gtX+py6WO+J2QhAeXeyRXm+12ozLBlmsIe25xUhbaPwnBI46qgsT
KDrsi3UJWrLGKNEzo8XPuUz/anhuuCLVuyBnTcxPJ7hWqJQA2UBbAsS5WUxIM+Td
qt2hm1Z2DlvNGoP0hgkIQNZYOX4eqydkiCeLlpYKZXPt/3B8tgFADqYeUPx1sazP
E00qbAeJPLpmzo0207HowKzZP4xl+7Cq0kwKc42eRm+HJxIPAszNFANnf5m/vr8A
cCNweKuX8TZwO68GQq36JtUMjUO1kKoYytaVwI8zfzlAQbvTAGLXBhtpiurH5nLY
454lc+CvwOQ2OroC9ixD04yTtRx300D8cfOjWNCiYNC52NSd9WqHyZSRcCXS60WK
Bkc53quloLbZNA5iXdSavdg+Px97rc71rSIZBATFLEnlB4eMdD84Fep5iUgxSHjf
+iUC0kmFqYZFc1uWZ1hLvv/RcRaQcfhSH8EmZNSiKf4U0zbBd2Iojc4kNuptbmhc
bBVUbqjWbiWIf7CGBbxYUjuOuA1qb5TBYPXCFc7b2y3k++KiEcMdKYFJX++QRWrS
E2O/gphAxBx7JmZ2rTYYGl/YcxFPO0NLjZsxBpaogeuwWtQa/LKbA0UM/IGrIdhz
+ExaTk4dNlcwo9Cckj2eRgLkrXi3mLAB5PLoBnXZA+Q7hO9cAMhvDkcTFPVDL2p3
Dl6wTWTtuZj9br/a2FlBAoCdQ714+wM51vHgpHBHh6DNfD8ctJh/UhuKhjbD5krB
ZmU5rhZzaqox8EV5R80n4X0S/ceE9+ZrJjY6hqZWRo72fw+6k3Js0OV+SAfZseYQ
KxtkQPI4sW7JyERECixp/yTVKCOpusfppM97xZCz/I7P3hGN3gefWGR3FaybfL8f
iZFSF/dbWxo/4frqVqwAdVB67DKyhbsmCkELB1UOvG0qns2fvksEdLqmf3bTMzit
q1q4pdbCUBA9HtAK1AjsH3r+g1L9FSv9Xu1ULCItQNHTdvtQH5bmdiCNIJclyGpF
0oDiwp4fnKpLWqLIOcM53a+j1UuLgkCTlhyag8TbXB5uEXv+dgHBxfKxxb/vo10d
60wHNLH7sgWQIeCftIyhrJ2dc/lseTsd/VZSKycaQlhJCZ1jIEF0LTmh8gxQkH9S
nf/rH73VBZbvEW4abetR1nG9IX1sMOusml/jjktBL5WMRU9iDglhPsTKzcXpAhow
83ldKH0xsaTxWYjL7vuT4CyyxVO6JhvnL03NdgWbQjjDvyu1d/oD8wg70A5gwoTr
CXBTVHa+QWJl5KlyOoH1Co/7arQXbrvROfoNW2jjnYwIMYI4aEjUMXKJwBjb2Ftj
XTsPX360S9e5HIvsiIpMsrn9JOVVlI7dgeESpY5uPVa7jwbDg88Bn/pNjsR4n3g5
8jx9K3ZUqvZmK6bB03R57VA+go4unuf4AHl6Qy+UZ4baMDZZCTxLypvWze/pEdQI
iSVr6yE1NUgLZ6E0wB/n7QfQYQRWKLcMkrxNhDSzx8lrM8rxGZVzrTM4XKN6rj4D
NTSTf5gNB5g+wyNRTWuAwVNrhObRhalBBV6MGGa3xNJjxMJHJGHDT4jbMMB68oKd
YurNDDf6eV4cCfL0H1hH1gCwoqkI2oYnZ8f/47d1zj4gyTlJl/YdoTNcR8fH0T0f
Sb3vgjwYKRF8AfDhZmWm9VcFfAup2N92NCRKL8v7HEWT1uAtDNcwVDIrXy7LLlrf
o02P+m+RZrj8ZfoV8iCN9exGRjpxxX34/El172fZDibQgs75ytZXuGBDFQRccItX
zdbcn2tq5dF38I/pD7M3Xw4ZPpB00yJyd/4ss1bIR7OTwPk5FFYvvpwTTt642j3+
A70YT+Ofgeb1goHlOgBJP9tllsaZSCzzzqGhsJ6tQypu+82pWwFmvtiPrwgLu5PF
i8LzKCCi5CdGHQSKP5dUpUhr8hAjeA+uWBEPxF1jT/2cP989ynG8/xrCKfupwYSW
zbgBb4ilvy2vmkdol46wb7yP/07N/la4ia5ffeqQLl8SOQlkNUXSyQvwChNIapxF
F/7w5hWE00ld6CBpFOGnFPuzvytz1qB8hQjhe5QnrV/zZEbx4ZZceHLBN0Lm+iCR
Wb6ZByCsLSzag1AOeO15hSvAo6PbSRVrkgG48yYoGiPWP9JCMeXvuhKOCB749PET
0FU6BP6KeSOYuptLwRNY92IcS3dfwV1WLvtPeDzwn2rZC9gRDhtNUtQLe3x5crxi
eQfkq0zZXNVw9rMSZc3ovpjUJuoBKY/7dnFlSQwKhAFXhHb9151BkoAKf/IKi09g
j3U4GqX+RWehh8bjRU+FTH/BIyBE3kdUlxFUQLBQNLM5D2Kcfwpc6MoMAEGIb3qV
EmCybU3iWNVRQapgp4Tmz8VbJeiXPsC85gVdNpLJ4tFfrcruJuqAVYyNgWWZ3X3U
y515PibPHcA8NEPKWEOhWs99r9F+Eq6RzAVAgN7hX/DrPJch9cjn1Qs6lSuqb9Lo
98VfyKzuKHU42CV/cNiymEufN9qJJkpfiZ1s3qGZ1vAaoCdI6lCiPP2zyBaQNNzY
LO7OCjM0KE3oQGD6MiGPPBuIeDZxvdHSsqMaaLWRZPpjeC6hG4VNxceIqC/IQAbs
yJDuj0GvLVkV4vci5WGuJw3RpeyFW8tQL2zTLSRuUi1nCqkmZ5+kmJJwjVVcCLvA
PEoiy4zS+CsVyZ0NibIyeNep/U6JW1pIkG3MiXAXfK5O8tmrbnCiY/6y4sw9UC8C
824Cdwh+BeJmb1cVFfGqwNvf72rUP1lx5ax1nqStzimXURcazfFiMBpKtg1j7hZl
OdFrTBMp74RbeRNyJlbGbebByZc4kZYASA7C78LqbPyORTAi00DPchaEwld4Iykc
gi0Uo7TsqsDmLetLOwo4tCXyO0kpbXF06ED/L4DtXHO2AtNAswUX/N9NlYbKgR2O
MZ3e00pdaRWdapSSix/SGBtjhutU29KMOgp8GlcRo+e8ZAw4CE8FJEStr3iFupgS
qkQy6XtahXeFltdZ5FoYCquhB8Tdvvi6CzFwocShj5FXQGD9W9e+zBy9t68BTXaL
Kdrex1KrKWT13yVseoUqqC14IF23+fHOstj7Gm/zLCxvyOC95X8yn04yjBNcKjBY
GWat+X/7QdeoyBexmBeePAL+dPvKBxr4FitWovR7lpiPFn+RxOI8UHH68/bF7Jyj
dUppW0S28BsXqtL89FNPYpSV9AdxP5Ucu6PVvHzUQxsoSweaYHgcp41We74SbC1m
U+VJpmJ5BmeIsQ5E5TZrg/JRveWKZuAVolQJLNjuj92V5BY6C6RDDiUKnknsQT2B
PohAf9N3MoejYfz55M/+KgL7ujXQHcSUIjPdyFjdqi/hqOqz9qspOLhovaojoTN9
TnNPaDpkNVJmyK2vuxf4/M5Bjr+HTO/UNei2CiJOnGnam1HLkEK5Kkuc2czTxueQ
qQox6kgyHn/2nwYN911BYwSbll6IbCukWo//PBFamW41HyYka3b2GDyRPKpeh999
H1O/17oqxCtKc3MNJ6KVfm03IW7exahxBA5FpCehOXNPVUcevdGDmYP6gEvpMtyj
qGivGclTfM9ZKvRYj8RXFCP1E5pVUTCrtu+BuNxMAbEzxYR2+AViZDNJGwFgN9hY
mgPfE8jmN7biehEQgd4tMjnf6va+kyT4Wht0eP8nMDCnvZxKOsGy8vdAhMahzhXB
AE1btCS1A46OKsrI8PzkgLDKVMY88Wvgn47xUvXUsLutcsbwEMsqWIC6Jk21hWxS
NvvY/HwiFZtQGgFTw96ENMVF9XblzEsrZLVQ3Y8MFL+pPoD9cHfCcU/fZ3JBuDRo
uwYFIOex1RPES+cCdm/ZYEbkKDsqQ842EAdW0DzcDikXkmNFSVUl55+FMb/qvpta
T4UpRzPHCShtGHqvf1MgWumLb9VuPioJMnJE046lvDTCc1mO+qggJFXKIDtTTfsx
cPqIMZ7mtMbL0ItnbT5YHyWccGRaJnv3O/ZmRnrkZDbqyrqR6IHdxUStQETXZ2vh
cSBLoUr/+0PPOeVWD2WPIaWWMkkaFyaC9kY2bU0IyUlvd6rHa/jWEPbRIyiwlKrd
/OHL5IfB7V5yUco7zLdi6IrvCczDYMRHxhzL7850KmGN9AmtV6C8E6Qv02+lKKd3
1n1t/6xoxu7MRxHAfuVh6vneMvha+qWvL9H34R2NBFMME/oUG/jaXbg6z9LDgqw5
p0x/6frRlE6QhLBY6lmjddrVypYPOlqUm4On35Fm04aDLaFDjpVStpORGCKQyiue
jxQOIOewyBAP1aXsWaml1fNsdudwrAqX9JgY8fq9esUo2lRs8OxlVr66am5wsCon
TsveCXJhb1Jfkd8p4wWvRZNzXuyDdjoMkQfF3vauHk/A1YKfiInKo1wDgxcBq4UT
ey6TR90JUgl26cwo6KvtGXQZMAVAYtuDPYVN8Zy/8lsy4FL/A8aoYZEQvU/Q7xkf
h9HTfTfO6wkj7IprLr50gtFrbY3tdyNdIVe3OZAGaAmzOWXXp1l7FGL1d68bewu8
O5i2dE7dMDI+1PV3OzUjAUiSLuHS8gqbZ2+VSh9mOmAiWHiEa9+qgHmyEfRlKnSj
T+HioM+We7dujLqQ1ujGWOXfk+f4Dctdx2yATu0380UPZjxab6byiqKXklikYGff
dTZ+Nb2wsWrbrUTaZyoeCOZPIZhLPmD+XCn6xs5STdRSSmeTm+Y/v6n7Ctu9/H1A
pagm2brOvwbtTkaqoBpQc/yHnsQKlJcM9gS3WI36tW3NpxLSKvixP1cFs71Hk4Dl
v0hx8FyIAhnKBAeIv1aRxLfUSgEy1LLq2c2T9w91na6Gdq73AJOcZMWlhHOP7UyW
oKylblW/o8LAPECCUTOSbKBjJSklS/PAnmRs/pqE4nWIUH1H4gZ4xrD4eePe6nED
6lggQG1nInz7a8SAx5rH1oSKg1E1D0CvugQoeKUYJxnjp4n6QCoAVuPpmGksJ1bM
ZnA/ke7eYJrUyBundZo3c9UMFx3jx4Scw1NpqvJkFKnG9nfewULO3WvPk0K6A2hU
tZiRYFKJfq0XpXn/kk/JU12N8RNURJi1qmkIG2PlvDOM6Ie4SBeJ3pniFKdq4F2v
3+JZQLdvWel/8x3I9VWGwlcIuep/ApWZYRujrWpYfZUTxrEJ1v31ct94ePHlhN6l
pGY4xeFxoQ/zE9yFunPVSxDcECUW2ppxvZTaU44uk0XSJ2NGVq+p/gQ0UNc1xG3l
V1iUbzil8JDDX/T39X+JF4QZuatDx3fWRAp++PmSxolOQj6qlruqmMZnXktilmlz
kyeA920xqEdYEZe+tQUGyYNCO/G5lR0EwyweXC/4j+ocEJ+2Nnmk6DPmqxYVAKWG
npzrp/urI97Ao7qzX/bQ3G7rx/m/uuTWYjbnEwMynMqs74MbybIVGU1JKl4hKuHv
xAB2Eaz2q5M67wzGgw3uD8sCg6WVtS73ogG/M59dIL7HsiHtPavpytdEqJZWDuHL
lmVZuiFxwJk0OfxrhqVw9S/6/RN523wUBZYibCv996Ab5br6VRAOy6GeEvlYWpk8
N+QICg3TNMUyE40hOJUki+Dy/OXgRcHlVTAmYbTeEmDnjPNo2GpXeqOiLLR7wMky
09QxbKBoBy7sJrz278ktAiyABOYkht0pH8tC5UNcXF+aO5+EgcxZg+rLNkej5K65
y+DW9lAKE84I6JaYteCrXolZ6xIYDt++1LourtughgxaODIty/CtjMPUwcQ8NHXh
7AUPRTS3TyxKykic4jxjgy8R6QNRZJKIQWImWV++gF5n0+YjEqhjKpGYfHciQ8jZ
0yKiLumV9ozTvEFhuq0PBOufdfG+3g5pyjpv0kV6XY3Zym0p5sa1DSi452+fzG39
4jXXHcsCF2OqyPelq+r7IGUz7WlwFVL8uZapG4t3DKi1E/SRWeqFGn6bUwVPT6l/
W8UlFieL9ZU2Hwds+OBJrAge1ppz/q9A/fkqt3sQVU/n1AtlgwHZALDDdROxRN72
DXLo2Jf8/NAMZW7z+LTbc9uMrA2lEkNQeY0V2jy8uYGVn0g8fMtF6rG6LTnSO+3u
knA1irf6M11kYBXQ1333jalO49+GCHArCYa9br0pGEEF8wbnJ6ANda4K4vxksnrJ
V7e2EkUIuPvIbsVYXmljSAqEcSFzYjEVxAlzFjhwXwbMDTl8RuFMqcdfgJUZIcne
RcJjOCzA4dOVj1Hij1fJSP1CffE6Q1YOqSj5MjHyG/iYBdPLF9MbXDBEiECfGNA+
oyaIlxgCg1F7yLKJEQUwiI+v/WNITyYfRaS2FfuXrV5JB8CMF7J2cnpVaYeySS1I
vYfaatdSiHj4PDCSpI0pSkvGaWjMpsWpgBAM0umxPjQ3IlqwIdDAr5hdbk9+zczV
0RAuY31Y+ss+MSIEH7efzjtsyiiXq/gQFI24Kw2sQRMp1QRZzwlvHLUEwV+siUDN
1+sk01A9nCAlimaOKmrXpDLbK9R6tPknn2Fz947DP50UGG6+Chb6dgvaLUqiPXUR
9dsnKPoOjxjLO9CUJ3y0vVg1GAW4ykgEsAPAuwTYmkdAL09nDyBP57Vt3ZU6Jd36
/5S7nGL+FPsIniCPVf3gzwJle3V7Y81Ge+dLHcM2z1JbEF0iWrDqFmTfTTpx92rH
d8U6G5eNtYt+aQ9qvgufrQiuz/bJ8jd1bBGzJEcF45xSzpB/AIctm7AdJb+UmJmO
JCMeNOZtxdIyF6OU2vrC0L7HJV+oY3jcVAzHdSToA+vHcUZ2Hf9xcyXthWndmhE3
BaQcaO+jMpsLUgTAjSfL9zGZthEdJU7Vg/lzJGWeO6j3Q3RuygRBTVzVuFGYPzRp
+scziQJ+qipEuakWo4oQDAGXIzfe2bd16GkNvvhEU6T3Dn2ImMjFvCTaYFcK7kdz
zr3FWBq9OD8rZl5EIg9ttFlnaYxQXHLbeeKA4PVA664ul6TvdtJg19T3yoA2x19D
PljzwojRqaStj9sVFWx9j06KLutRIMOPGydzMCnQ8Dnk3TzYZmb9ecQ6ofeueZ0G
1QSGHclodcpZhIKuvG8gS/eMShQyfLnmVRYu+IjEBCur2UF/TKmgD/aePOrWbwJb
2rQGqOXKYoLoAIQ+c6CrkysFfq0AfdgsmHPKpymitgQGPQckx9QGrYiWFVz2P4Ai
2XPlni5mLJENSZp8OB6yhae6MtnksJvqErcWcgqbxEn5iFxN2kf73B7dvqiYU5j4
Ozgb9aArlhczmvKhgVndRPK8SevE6KSnRv2GH5H02DVOxKoMD8M7kD1xaZwGFDQb
71fcGhf7XmHQ+HNMDbVXBTalawQGAEl2YHfymVBcyCiUFGnPpJzHTGFqxVq+AVQe
ndl+467MnFEWfO880DMCGU1bbgmM+slvtyhZ5Yh3AJBwPCzWg780CpALDuVeM+/o
NIYOiFXQ35we43lw/cuzR3UGIWM6JWWEOobwGkNPzZp2i9ouoGy8gn7EEx2OroTr
Dox/fcJL+LlidW9EvIPdw3Y3hv4jPadQ/UU3xsh5/Ra8xk24r77oGg/Znk1/Q2NA
q4Yj3c5PCo8cLXxCSXH6WcyvhzvOjeX4nxiSyWkWirlsuRXHrUvIejomAKMrAQjx
GF3sWfq6epFMbri0KF9je/qqnMKT6h8gAFldG3WAKzb00p/fn6bDf7YCoDUEvuV8
eXZ5IUKWlcfWqvYJOBG+FLQPn3Xd+ALraNf6M7GSyUowGwxb3xiHgooko80ngV1W
A3yYZl/SrnmrzPBNLhFbuQvdxZ4gR/cUcYZonuGLWc4lNJ0x5x5a/p/KIfZjNFYe
36vdrio/XNo8SvmReK4XvNWjkRoXu5Nmkw2WLaZJF3jjpOlqYnzkN71QmAhELrSZ
DMpiW5YdhBfw2L9cKjHtUZZv4cWZGxA9TPswEOnKj5O1v+zVCSPbPYfTnnGgzeNk
5iH6Q2eq43lGZYasGCntqZBjpx9xpbsXe3H6MOtEs4RCVgkTIgtzKRD/7QUlF2us
/OvVxVkxM439ivSZd2bd617wHJbRiWYInMq0f/FVwoNj1tR1bWFfkMteTKVkwd5d
ovVjcaHn6ooql/ZmcpSJiTH4sQcbvEx5HNj7bQH4yXXIH6E+1oGpwKXx1RoPWt9b
f4NOlSvZjefkZBr+do4ewQ8HyjaUFoV+0ORUT3rytgzfQaSsnLy3t+gUw1Jak8NZ
DzPmaQabgUTrLovXGf3Tp4QT9z8BOlZ6ckVRMfmHkAL5sKSQS87LvA2FVeUp+79v
SRf2GMOLrmUKNm8aJ033BjyBsHUtLR9Bddjjd+0DgIogN+qdVDmaf5YjIE7dQNPc
/EouOQQwYlOBS2zym2L6jDLTs8XddRPXkzpJNUH6sbYJcA/dDgicXexaUeWY66JK
/4mJMBIparDxGvbrcPI204CO94woUpy2JN5ew53PCRuaUPVmiSr3JyBDGieBtj6V
WGV68i6IVR8p+ptxQCRz4RdUnKy+kN3B/qL8iVqy+WXGlSgTFfcnNy2cJQ0vQfJJ
pb+RR5YbZQDko+q2OhxTrnhRPNx4dvg9wAFvx5cUnYDUgRwcNEuSxFhHma7l21Rm
1O6iS8yvu75Ht3Wf+b1kWB66odFsthcRgU1tHnsFGErqItgRrX9uVB7FzxgIXwku
0Qbm7PRkfk8/9DSFpw2WHpDEVpRaZLEqfzu1/S3IVROIt1hrlHi6n1+dU79GgSfk
Kuptvb2o19tkPp/02PDVlHWdMReiMI2Nmpdh9Wd49M8hvqUB1CasElML9rJq5Pl2
4H8Wbqu67mFMUtZN0nFLouU27qNfnRkS29k+7p598TVan8pqdNpHsFfapRkOskSk
8b67wuXYeNsFpgJGzhBxC8XujV3O/UijITIQBzTn8Xr28fbBntQsrPRqfszAvaCh
SVKPFuFvctk2wYPkbzWXsGZXT9Lp2VtND5t7/P4NmWClGjHcgxtoemgEmGeqiaqC
ofZJdpn03vobc/fws44X6Ngb+/Ds2DX1nyEDLD7hVvs7TlAxXaK2ZamiCX9lTpNI
dqH8ljIyP4VqmJTgxQThVYkzV3/RqxImBgAkgbi3qZ1bALOD7Sqc6ywck4YiiT0b
K7Q4KHvqquNeSRsp/1UA9lJY/BlNjCkBFUkrOC1E4J/8i/043Rl99VFdvg61Kxb8
xKLwCppPkheXAyDhMlhsFUGcG4Yo51iJy3VvuivpYrwXUOU41Jo0wq+hgmo7vAHd
iasuxsVjcTXQ/9bs/pzuovX3QOUFCckyG9ypOZz9D7UWrZXxAmYS+KF79qryn7g5
gBriA71GhoNR3Awon0xGpUTCPHbZCzUT/0EHvpAApW7JxP2G3QwLpeuScvfb89F7
uvRvGmocbCyHzpjdQTBG50dLx/07wlcj/ZcDssH3ukae84BdFZ5R7QoYFedSo6T3
ohazWFYCLe0d61kffiIhXET9lo2iqZAZqjZqP8b7VPKk3uNWOV/QZMPlyHGvs0fZ
duI+CYrPli5Cm1jlxU9HDutwUe6LSMgajoLN/WVewWW2An39vDV4d/Al7yKa7iJM
FlkP+FpOpeVxoF65WmsRKCSnafGl6xQO6Seah5N5+J9bJsK8xEsyu9YZX7oVbQg0
oXceAbmxD0O8faC6G5LypIMy/0cZwEk4zfImonCR2g55xE8usIH27yGnqGKALIDp
e0P7TG5oK1UC6O/XP5aCXRV87bdrPUTeIwOAs5w216E2d/5qQo8KSnW3G4oKKbx7
FoxxMKoSTCq8bhbJyPF+24D0KdPtOx1uied9qpN+h9Bg2w/rgFQW2zf6nxhBPIOX
geiM+FeBK4Y4/iWh4lI3ebHHZ517HDiNiT6j6YRg/ADD83KxTYT2xKmbnlPKhbIF
BiEmKZpz67Y9uJF2g80fcUNuqScZrGvslacyNiFKsyNiF9KC1M4djvnKFOQsqTCj
nUwIvrr+bLK9R6EsF/sDFFzaI8zGBakbLDdEfBet+/5oyn0o8qhFUQOMd6GN4NZr
+JqpvB8AzPnTBDEdqDQwJOH98lLsdHxnCotzpEXklAAJM6An1Cj0St0X67WXoAey
6PcytzDEQ/Aoha6RpNUvRSY4Xpaglxh6lBkdwhMh1pcsJeoKrbInStlDoFO2ViDi
YIqN9dlegOlBMdz1q/iyTdKQKobEV98mPqvwJrnaHaq/TcX5CCr+26k2TjwudH1x
pU8JNdjVLBOMEKztzkmiM+9kE9m1Xn+vf2y6DaVzQN3mDR7r/4bN6NxHBa3LJVFD
DGXkYdzXWppI6ETEuCoUkzDebSJ/p/q4V4vxEY2lxh9GChm+OC2veU9P1Z43okNt
o40PAIAaXG+76vFm5nVbGxj3mnoDNi8JvjFegVQ99QVHINbBwvqJPwKTx6jPLWwI
MD/zIB3aS+YxfyoWZSlE+Z1yjPKfZqM7Ny4lSrhfIG/5qsS3gNKEsLZxHJ/sknaw
CkKeOxF91Wqual8e8ZSZzFr1pk3mZ4Ia7CPTWLvP8zBK9+5funh19155ebZx895G
vxzijkCwadF1vvugN1e+RHgR6ZaM/jgF9ftUTZhkxmi4cEw7dqh8YZvhlehVDUsI
s3JrQRwXiaw9wG9V+AungakmBDmPpmWUkkLCwSl4C/5rmlearLSX/ukBJ9N7qJHx
MDHdA3KP8Nxa8/fy9gwRt5byvPAgVuTf0Is9CdA7nItkjvUkxo/TF6quCoMjgn39
hFPC3pdmGR6qDSgoLIojOzaUE0Y3+aqZy8wQkL8e23HybisPlI+brkLo05D0JR8Y
Zh+/T8MZZ19NYRJ62UEmL9lEDlsh+ViaTQop3j8mStmY7m7H7SSur/frkFhYZEhm
pfoTNe8CdFgYLrA3Met+jFL0HHK/g0tr3rQXSXd96m+qL6t8d0xQu107YfPz3lBR
i0QL99r6kzI60AvJ6hgZQd2xH/2ElT0DpN0T/rwym4T0Q8OeREHMybhsjkss5TEU
1A2+k0aLi9wEGkStz7RV8jK2UrV1+0AI1KeIEfj505RHjXxT8LOIM20svUexzTb0
9Io6lvjcDOjx0hiPHEssL0vNwi+FEtTUuSfkJ6xv28oIxva9fuuRUs9/+UJYXDjz
kginWmsUygbrRghardjuHzFqd7j7JPPNmTLW/dtKTKxrS55RWvXVFqdm5Z0sIDmq
NodTuqtZWJ38Hgqm29l1iLmkAePgK7r6uT+61pLvrje0+A/WoweSWhg0IjwhedAp
gZg9lswbSRLXLAL79r0CY9ywoxS2THVbqtmvZ/vXu6PPo7UNeFm2LFfbrvgGwDuZ
Nz1f5PnswzdM8abEbvDSAOi1ZSXoTHeb8jASoobuqliyqYpcmFZUc0DlJbo+7fxG
pKxVbelwxbGMSK6LhkEglJyMDnAfpTjs2rpBv4Q6x0XbjwXDGA/VNiBJGvEOTLkK
es2ybc3RpnhhBDDnh7xKddhIVSE7IRhGVf7OhLJqrXNjkCoLczigOTmxGl8J1A7C
7mEaa9+eQAkTk88Iuw0x1hfTcVlGDzQueeMVH2QiRY1XtOO2rzeSS5K79TUCafoL
NRktBQOhFwndH0o5x/mdQi6u8kCFKTqsniBABU+fshiBJK7dxp2XzKBaM6gUpfpL
RbUGaf3LEKmXT4ETOM2xWIrOCUseZe1DJ6csfgPkk4JGJ+4ZUmR9QI0IE3jvooCv
MtZAGeQVRkU7Lekegq4uTi0/HZp1+W32qWafCwBGNK0+dLJcXwGKsCZz2VxztoSX
bq8XO43+gQ8Lemwbchj1jv46J6FtJukuqZ7wn8hcAot/sbHVnMGY4v3uo9czvVIn
kDayCwYI3VGieSxj2iPn+BukNjzwgk4L7dV/o5z41/lWSbJWJExjnAu9KL/SyvU7
ZyMJOl0zTHq1sDE1qd85sR6gxv7b1qg0c/ymmsfP5ak6/M1yO3Wvkv4a3uysUJJW
shBfVvzwDPsRsGXt8cSM4jboIlqT5Wg8oYVuHdnGNTfDjoLGznArZr3kNSkKmsgI
VJzwU0NmBAgQUXAY0sYT9iCYSyMlJQO5CH7nyc8/qtsyNknyWPYX+xlKE6msdVw5
AlRjA0s8WKtlEOMfPjs01V6k/vaOY9aJTIxiWg7CRSlZigCDrQf7XSu4T8fRXWJ7
T5kiwliyCyJZaQigGG/Wh4U9KgfcXPcXUftW4sO5Mv837AADe/RJaqg7nkgVrqM+
7MSHijq9YwZrBwG18eQvJj/0+KJOybuliXB/jtBg70ggHdCn2SleeGQTFcw94t7n
tq1AT3SwUSWH22cdP4Pa3Wimu5WieajdYGH1ArU82jyMpCwrQjVqTE8pJo63o/EN
pDqsQ+ZRhD5bc4rhnNWJc0CIGqJuzyxJGWrO77W7sgI3avgLNNSWspLuDGtjG7HT
C9AI15tE1fLSSJZUcw9Lh1vPAwhK2yteja433o27LQfunCxDRvUak2+z30se8Iix
gi9mb3MRsMlVPAuiNJg7AyLB3IEB/puowj6CuNQxFS9orvsWdLw0+EhJjpUWo/9U
p45xMsA/npS+6hFjV1efzEiJ4246xCU7xGCZDwj2UhDJ+ywuOIRH45RcgCHXJYWm
GCAAdF+QoYNUmRA5aaKrp1dfIA54p/qAbz3JrDpe2bYM5lN/TalxhjE8j1MF23Xf
tJop3QAdRwC5M0mURAzeDeWPyR7RvmjVTnN+VLQT+L4nEX6FpcM6NEDfa2o1xwSE
No4EQF3/EwOmTZd4aBedrwmEF7LzYSxqCH4PD4e4hrogtURl437046oia91ZEGom
lQYNxF0p1lfvljts5dRtXBnJCgYAzVesGwk1fg6ciww1tjGBeJRjVLPdyrsMFvO2
RWdhOgp0eA6aYPUSGeEjYlm80STmhsCWJnSp6FTGLQRjCptpa/+foaXH3pXykLam
yIsN2YJtsvTPeSb1qLnEaO917lloB9QQGuI4Odi/+qvf2/k+WOsoWwJcV8v6E5EY
E44DzV5D1sZawa4NxAKb1UkIGF72hQ94C4TBnz4RDRajpF8cO4VWvnBC83KKe8vz
hw537lJpjVDZLXQzREBFe7Y/l1Iaosq6FZ1Q6pfMaNOcV37cdkysBRll+SZtUDCN
0M+DNrtriXRDYCA3VokaSUXOCgwYTdGYosQL8dfnspNvbenJ+10Su19EPIzHiu+f
FBWHDVZrm1mDAQwtrjSb4JIpEo/ic3jNbhXTtvL1Yoc+QLVdJiM4veBXBqAmfko2
qznGwGa3sHldbFouEYbQKZIRd89qd6Q2FABLeTLw6kLOCQhgNAMcH84wQHUzLWGq
jnRkS24KOtGdDAkyuJ777FLgNZUELULPyDiD77XmyjF25wDT5TNQdJV8tklOZJvN
Rrn0v52N2oy4eawlBAN2SYlI7/m+yi8Q1T8fTWcS5ghOs8DmvUK03OmF3PkW00e2
nETzw4bPr75f5fBlMYq692JBiRdIOhSsbfs2DyNqgjnkt9JufO8i4H71SAyD4z5D
+ZLbIWytVd4Nwup1IVmdwa+8uvQKYe6owjGbBKcws9D6yKGfDsn7P04ZBPG1Ct+F
vWkj1VYIO+0EfUC+MguoE1ybPcOXRZH+5zNGl58YEwCo0K8NIjf0vhD7w1iWYCRS
K6aRWWaS9DuIPMIcXn17cNCpj9XT+V4n2831zaAqKg8gVQuL5Q3Rmj+TEa4hqUbD
qV6M996DBzYiXMc/1qO9Q6Pv5+THlR3MZDcoDxg4HBSuZ5eZ18d0/wYB1IHMt6K1
6/Yz8RRGo1pHEjO0/M1yeOgBDbQ1W/FN0CiJBXPpgPS46xMkjevVhs2qL8hASP/Z
8lf78E0KMlBZE/jIVWX7EWASJPwYoP198GijKNQhA+fW6y1sXd8u/hMSY+Ua8Dxi
/z302vzCcuELyQoBsTWJfYDnZqzTeecCgpR1+H/i0nPzsC5AH+KX8J1FWisg5QXJ
TZg+8fZ645dkzMUA7arCpfh60QyuuMH4P6wfdGGhW2HJc78cpBGVrfb1hZNdQGgt
qd9JM2rlsigY2Rz5KjzMNdsrdifWNMhWJpIGZgQKHcp9vS8+jdWgsYPcnpGzu48O
RPslvOtXPipg2rDTXcnhtGJHrZXozpzO/yzNuhX+myUTtKlo+6TNXEbwN606WqIP
Y27nsjfONdMwwbZOqGR34p5t6jG1/ylanD61aRFyETa8BmToJiaLFhgSDztf6TaO
GzP+amGpW/hFrgWe3ugwwlldRrseiR3n4jBvGdmgYfGukr8w5ly3Piwone4qgbcz
Buw+mE0SaXSFp6x3HdXraLS/M5FCy+n6GeIGGHL7+0RtFpqHMCVohavKjkqHpZh2
SVukFRFNWvHWokAzPFmQm7ZfnSRsu68+PU3jKxYG07VnOVtXOwfNcKTYT9mJKJ8Q
+NixiFMO0wGXEUhx0+TbNQHqwimwzIFlrZ1DhfE7XEEUvsx3b+i8Wx2qwnRLKDNq
BxsxX8NYAMWDeunF+TBUKyVwtC0CTfRwfuBRtcNSTUQ3EE415MFR7o2BQ6TV90vA
ESRUr+OQQQ96PDiyi88/cmNWxLnrh1JEOe63kOw4+3IZ/HFJJ14GVUFYc6IWjrqC
AmWUpzppFY0dziNYFSRW2kkvNZdzyAiEHkSEs3RK/2NFzV5HEefMbRQ3d3mCT+PO
JrXXLZGSHR888yqWjsOsjmDkdz1ACyGQIwjbN+GAOzDX+nTJPX30/wss4pbHfa1u
AV4swCQ7WdulKRT3skcHl3rTR2vpWBsA2lB2z/NYE0WPLV1K/bZJGcKmaEySSUzI
QincVxSdk34lkwtYCwnAovJPGYqBG4shfsfuuxgufyXvkB1evELne51jsxavssgK
6uvM8FirSd+48/Pz+Uv3PCnEZ402qmYRC8aGr+zALxAznvkOtRnqoLGuUQi7ZrvT
nDFU7wXuKaxEkiWuY75vSnRbv3CDnflYfkU/bWNosIWju17Rlv1ZE4LAfbDAINLx
M/2G6PCH/KFxbYKA3fKqfIdanjPz7S6azTQsGg0rx03ImzoA/tcZ68TT+XYUgOU5
izMm9qTCLALcmUrL46OcXCNyEFEwXBXGO82Fh0Vo5DkIxXNut86FUXvICzU2yK7v
JPpt6kKpdLkEywRhRI4Ylsr0ytNOW6k1hITGtDWjuYsGD03oeB1iSgQtMMCcQMqU
PJ8rkwT4ob8/agN7F6BphbJzJlbEZENrth7crNXv3u74+9/fhZXKX4ETF8RrJfpq
JUE6vJ31YoZf4gu2l1xXwZnKl+a8S9mDeVJi8PsXUKkaDd+OA9bGD0ZpHm1AS1lH
H12DqsoakS3UG5ArdqlxL33Z/AXhV1gu4TtEYW1/10CGEP5jYlpVthHofXUWxjR2
Q14PpMgeE2dwepi6qekFOVwACuMNGG4TfO3EHKqyY/rIAB1r6fy2MI/gLVC1uEWI
JgRk3VqAj1ZJMxMgYm5os+eiuYDezCpWqUqIlxIPIM1JjWmyg0UDNV4fpN0/qhI3
lPMPZ79YpDpvn2bdxPfyCZnIW79pGXs2OlDFQRWED2a9EqHX6SRpf76i/kxUa6BR
EAOAbtNC0jezV+nS6QtmJ/MEOHsx0UjWVzMmokfZm1GqVkcSQenETBXeLLB072nQ
fnovn5LDSDZRRnQEyk3LX8Q7TJ1oIu1FDy0lPSse5tY6GxhOmLI2GpOZYUJ9iho2
peOdLfhJSNuAuKn/w5dgIKgw3lBlc4tg/aQESfpkr+tfVOQIPEQHi7TbC1ubUDI5
QrWQcn95+oF5gvl5qOeVLPoMae46J3TAH8TCcJRGfKE/iOHnG+ZYJt7ud43Iy+Wx
hByxK3Jz7pQSwgd8IrDXmV7skYn617XP3RBkffPJZN/PYIqWs57+W6Aa/oRrg+m+
q1zrhkA2hnIv8Bu7XUQ60/eKR9oaGHq7AEbIpyosNjXDSt1cSGRE1NjLAUjnw3i2
p65JVIhG9oSDnn7T0MQEvbOSEFGSEhd1hDeEzUU41jdXa6ItaDDJFf2kwI2NJxyP
CPv99s/v7n2xcQwPbkfxpmQozudw+HZta0ykx3lnCGcRcImmmu8AH4CVslHRkuGx
VlNo9zIiNJ4O14EoaLXdX/4hm5zY8ggsEa0Cr+FRditfPY30nVijLeTbH6hJ/tXW
bL9AYnOalJLjBwsrU6IgFdp2KOgRLE4WQbjFGNUuijyHZ5b4H52hL87eijpxKVxH
lDP7bb7XMffj3KbN6QRwR3rWCKnPjoAKYG0vxGH7xPV5EjAIo6vXot80SVnqrJ9Y
9EmFghyPdE9dbWb+euJlCE33XAffKjv9TteRywRPsLwM4kOKxo56l40XX0FjZU5e
HL2gQItYlMUPssDexptahRrnmnM/XjwNBXov73i975/je76AbdUQXbjRHzG6qt8N
E88igebz/FPanDkkwkJ2Lt/VAEEzrD5f6ipLA2FFDpHIgTePUsytPeuBTxp05pz0
UjCyq6r4ev4THY0ZVxDzt3UGxstaCA7lAjt4alwRVt6qib6lbZZtT7ilpcd8cj2u
O4k0n+gaNLLKPElWQ+dkjUhIB1g7SropzPHU6a9VkYzr+TfF8LNaMt31RsQcSoqu
agdpSg7ggfRWC1d4hFkMa7ywtiSn2l+Rmd0lpTxFpcw1BtrApjrkgRc7sjnDIdQB
tMS9jc+pILoIimD7pLFYhOhcaIjRzQOU9vROBF4N29P0mCvnqegGYXaAyN2NncmC
3elBAjeEp5r1uAZpkNHluYil0+Vb02SyrP6Xb6l+g4aNsV9EOEN03KPyfs81iMiT
i6UAsU3a4HwRqLTqR8YtqaII791pVgUxvhAYpJJZ5FXkkNceYIMUSwl8ORdQx94V
+MzVhZDcw3jiN+0p0OPygn/D8LtVhbNuCFREc9Lb+EOS600cCdK0MH7237f5uuv9
5rf8sRcDuQP2KJi8UxydJPoCgNKhv7tBWaPnzxETLfc9PVU/Be4VACgH7zx2ZYF9
bhHYAw0WiZJKoaBWBPwhggRT6qu56EgkBZ3ZRIo50rhT7R73QpFHR59pVsTrhis9
wfEMe8TyMxf+maUKKuSON5/cv0zWa+IDUaIIsgY2DIHQoOoKG8Vig2sl1sO2yzDJ
jsDAz+6a/CXNocuHMKufTtREnGLbr47jpGgvC1wEHkFB8fiytlEbDISUljbDSwg6
D2Nu8QcatdxGELutMtdohrUxSJSpvvnM+7Y4lyiiOGeD+2d9oeC3PkLhC7EJF4jU
IAzonSLxOTN3VQJq03uPdTVLxh9zVbdQtjBZYU40USJo/ypqH87n90N4QnaYc+Ae
CBZJw+rU43JEmeK1uc81SESxmeXnddF823O7jKUW1rxGqsItM7QfnLb4ihXflWrG
TJOMFwMmL8nIJkZLnfv5442SqPUgfpV99yLa+hSYBuoh9v2K4JtwDY5TkzmTwke0
E+CzVNjK59BFvPk0h4OwVFPonWKf4naKXCfc/xcksVnm+41jJIG6Gn7aI3tgN4rZ
oCIBLcDjOTjnWnkDz8uIYQgUbcQWCqh9MMVHCASq/rHchuoitZj3omD46IVr06hQ
MkkIn/UCMsuWCwxBxS9OnmmUb6WIYJFuEYWllFkEb1u+D7uOVhMwFLwReSFn7VvW
ltUI5o9iFZCEcBcOoOzqseRPR7Xd1klPifSYpyqIwZH5JiXh+wQWAHS6o1ySyFFO
wMbdlBaRVZf4eqCGERlQwAkJOEWum+uhKb+Z6ne08xnxctoxd3XEj/+FilOZJiP9
CFsaGCO8+eTKoljUv/xcP/Vo8G+AAOL+mrTB6GfSbdvnNtNczsRap5++sBxHL42R
vGiEInCLv+lpfUZDqBPp4AgqGJU6t59pJoo4JLSvoPKmwyFo3u4Kg7qtcyd9FxKP
jTYV5ENaDKvWHLkoaoNz8RX16DHwD98hBUnIk+KKQij+BSjcT3yUsJW0Gg4nWy/N
znNxCTpdhOnCby+2g5KzSfa9FsBGhiQD1yIcUvYc5hvQvqTggHyiNLCma6XbR75K
JK+KtyV4AxNSxsa+Q7YuvE6z3YI0Mv9mTnOUqjLrDXAB4m4EIypINaW0c+LnsxRP
SxfMM5pMjTawfYF52N4gyvKSS2JJntL0fJnQIa2iBo6YzUYhni9m/3nmY2ePoqNl
8FlRSOr/n/FOjhc2mn/7wT5LJ4T4aJAsL6x3LADwQnYJJYauS3bf3w70KuBG3NIU
98Lwkyg/ssb9MFJYF2cg7BumgupbnrhGUBM4od3JFs+GVMJTH4fDXBLCDct+Vj3V
fk4emb57Ysnfcc5iwECBCFUvlVbrsFyts8G0jYmvvpRAJDavLY8kXSd0u9OmVYHz
nDVpIAL7jP6x3tfSTHbP0gxQIcondIlbWXD4r1wMsIWLlvn8hDRBhuYFqTbaDtJL
NGFffcqPm6HZwO/skLJ5OZfclYKuH34Lu8d1Prwus5BR2yR9xgXmDvcJVpZdEV7a
V92MEHz1ojMVR6E82TEtYOTltndMToNlUD4QfOBu2pcAxPQ8+1xLvLdoK+YY0o4e
sgkfnSwwvOJBjeCcmbOH1hiBEeyunuK1YvCWCq0OdjoG7bohQeH29JjGAzeYWLvz
klydJM2Z+CPyASac8cftXv38jzmZRMlMJPHZ5wImCGh9OWBHGHwp3VozqKwemLzh
1td/P9unBtlJaG6NDDLs+49h03GYEg2o4yB+rekhC3dIExtbFGvzbbPw+osnhlnG
vHBeCCp+eBNfngELo4pF2LvrMwwEIJ7V/OAL7ud1pwfn1rK3nsuHPyXcogWZzJqG
GA6dVIRUj34v+ncRtrRThw9be/T2vyv5bc2W5p6q7wlXTFFWB9/b9JiX2ohi7IVz
FnIQrmelqITTP5Q2/LYHH4rAuKfFRWZWcLjTVrSGK+OY0/gUpRvPPDJXJWWwbLnw
jy5lj3xCcznjfCzg7RbFmfBQ5BW8e3yvDMB8/NuORMe4VPSgWZNI9nh+XqHy6KSU
nVgih0pkGeBJDke24tF44Z/PSkNjfEvls4xGeFXzvUSSGZvunjFFN1Ij2apLWQR2
/ZFVxkM4fewKVv/13LUqEQ8Kl+4dSVRT6X343++o/0HaSwl164wgjJvvYZ/A4EE8
BDQdIP8IPH+8/zKlmv+uLLV/tXX474YQ7xuwr5PHObDQSJDG2zi/MxBmWfkV17N+
uDnCU/t7eA9yThiKbfV8O8ml2hjLqHN/CmQ5neMRIJe8uD9icoDJ/x80OJXLoAJA
SPXfbt4TRq0mZogINLlEQcEkey5LWHuaCH2iKzrH0p9DxTR+/7NwqErUeTog913W
b9ULL6e2wLLBUxGatjN08RfJcHscaa+5rsO7ujq2t6xaWsyEBk3/a43mUOTqkJgX
yK/SXCmkidVxiJ3OBA36lU5PcbqF7YZ1Vt0Vw4FIOK3Yp6U2bCQi+VzoMPbaQ7ci
xXGzV8z+Yq7SRoxFLkvi2aB9PRbEx0wOWgV8ahHlx02zuubUlTjtXBDeKMx5KcOe
FnmXl+69yjhDLzbTIpnaPUDj5UPdUz9RIuiljDIwQUKVVJ0CLCmP95KTkLjq8JMs
wMNcs/00Pjii4QyB1t/NBq5frl8xQzXDkkpSU2CJZ0fGBYky2QBuvTfbFw6ZtLRB
oc5o35GxcLCniU1Auz0bNcGkSm1vd4zKX5RKe5SobLnYjPI0htmdA+lCnaF6HbiK
gteSZ756o7Bk9Oj+fPQNETyLSTKKgDKF3RAXHy/ICH8TNsYq77Wcij3Y2e0Sg6S4
HOde8d1SOi09MlAavXiH+Ryfjt0KROFApVT0c0PDkFAVgW5vJou8Og8K1irAIwcx
0t7NB6hOpdOxDzqzqg22E8j3gdYQGrdm+j1+lqDSbnGNI2sPUhgjhdoPi6qdelkV
C2SvOMuP4mVMd1bcxiEOpKw6XSPQR+EvxyJ+KJgYS0bQQDpdm+YheAwdgjXDhl9y
ovF2p3DmrmKrGwajsHhweACPmn4fWy7guq3A8RlGkOWxs6oY5sqOCsZX8P/OKXo1
30wWCCYL/lE4jzdlZOTSydHv88gg2vVJieBKpMWl1fDZZjGUFKcTMVmFu0+l4Y4j
9oJuMHY1vKcDudzvXIX8gPd1+1nOPAoiP2D3Ua0NNnBxYrv8sQYAZG6p9ws08meL
q6dcGW+L9OzTi3tO2gQNsHsFi0n/XqgD4jT0yaMYde1EM+SMZ9DG4lK1cANc6fSC
KP2w1OKxn5KCFAvzeKT9M4zbxIaupaqQA6MCHPvAdHVOrHLZorGw546TKI7LJazi
qH03FhXgGaE6AUdwCPX/YmfivDrJTuAtPpZNGGY36q/CX7AYlIqw5YHQau1XPPZi
i1ff8AeNkSqL3arZt1nt5MaS35LXTBdV2Fxzwbkhsev1aMHedfMy8erNJeGtIGDM
ZPhHOUwg63IpJEjgEds3QX+RqFGL2WY2WrN0/8GL8HkXzymbPWbwHmV9g36oaA+M
u91Qx0cgeOlxDVG0kJ4ZsBySYxsQuxMeKWwsPZDQ/6ILpoDIMRjdp2h8nK2sWTJT
Qlc2YV7F6kTqBQPfjr+CKQC+rJjIgGXyROIfaU/rbEIsCEkXIsZAey0domi6sJV/
3CFwG5nZsf2BvU1Z6VJO2DICbnoQjeAs2ZrMLwKB4OZu2OeAmjQ4wITP/+Xk9XWD
MhAFja9fqlkNEzq4d3xO2m8CUlM3at++lfJycIBP31LiyWG6hq1IeSF/D6MWx5iO
iLkw2rq0mTwf5PMB5Vyt9jXbRyXJ6HKC5mXUXqAo9DPIUyz9V0ZG6bqmKRlGtJsN
Fr29smpBMsrhqbCELK+yAltNn6Jm4HQEnOp4IKWnWWJuCreEiLIN4JzyQ6RoK/kI
C1lodQfgFxMBobFozMXyKk+9ZJN0QbFo8S9im1URQaB7mvQINiJHOJ/VwvObaCwy
coa/TBVUB6N1rHGLJKxIuAKpNI0IzURCo5+Hu42UtkXHLS8rIOxhpRKnvXCYWq3R
mrBmoHGbQ4rPHfkaGJl3ohn1h3bV/KnDHudLd5+NfqsPtyFRYZcejAn9EcQfXxNY
i5BPXlZl+c4yKSKv1CmDVjW+PefptDtSxASniVy0Ix9hv3cHDI2d+iqUVY0zxz3x
8WEKkT0BHm9DUWPqPZZPMaGoojEYtkNkDdFSccOqs3hD7tNF2nigEc+0CZm5fSYN
I2VGECHZAdYXKdgiZtL3lI5v3JY6ym3Su1/rdXJuzOBrCx8IaLxJ3diDO7v7R301
PrdvSRRj1zUVYcBKi2w/Q1e2x2e2PqkpnwbivD5/CrE3Wl0iTORpgYdnjGftZCzP
h+rjUor3GlH76E0Dyl/3775J1ocZEZu+EMoJQ9DupYj1ZPVc4m3DzM6My8Im1tDb
ofcTf+2msWvrFyoaFW8u5vmG/k4KJaQrGU37NO9mvUloMDSdouO4am1K0t8PUb28
AamaItV0Nf6+nGY7lbYJnwtZy00A01mtVtQiuWrwlnW7TsAdQjNa31FIOhpIGEf8
FUjcf9iQH1qfVY/9TuwlX7OZf5m3rXfdJxaP0gKjr5wAgsR+UxzqMHs1rV3JWjj8
MZsDJcSTXNbVwUSD40Dg8hRcGoIITFxxCldvfrXVYFU4wytImHpD6VpH6gxlSrGo
Q74c1Z0jA+4toizUhz0pkHVDAUNNbP1ULOtSbME5894eInsHsd9tR0Xj0AX/c0bX
aX9jJ+XxltAuRQvTWLVRY5dIqouDoE0KRzisH0RHqiIFMwm8Ve/sX4rlusPJwK/M
KgaVuEZpbe/mofvLxNyhCQXx0/jrWiafGyZQ0sPls9ManY/YB18YDXAk8Y6yhDjV
/WMb58/0/D2kHJJAwXK3adYkNdo+i4jgyoOpNfEt349otu3LvjtMc136SiitVna8
A7mIGM/7RHlooF4WVN6vRmYoqxQ78dSTY6DmCNp17bDPgOA941uRRLJEiqF36Rf8
EVRoqMK1gfWSUN4YydYEDxsBaSXSKDZYKyjyLSvy+15XCDJoAaAB/Asy7KxVVr7v
Jzy6LbqzX6rosqykjNq+IkliXLmZ3GG/l+/iqa4YoxR5ivW9rCdXo0P3XRpS/gT+
0Jn9qaGKIGiT1vqowGXe8xe5UaNjoqUmM2bBQR1/KX/8T9afigVW9CI1lHJ0m29l
DBUyMkGxyIW8b7MM7ZIU/H3PNKpYytgiQqUEJov1sMPYOUMkqZCKGZRBnW2icnYO
D/9imRj5sbsq73EQCEZBKmVJuk4OVAZwAN/IBukDOm5aMWQf3HHb9hnvC/E5w06i
BXZgtW/wSludPr9q959jq7rinSngvYsqO977kGIhGQiKyBaOsdqgkWZnOh5Yr7IN
aYqAvC0YYZ29V7+2VrOEZ2T2xW9fFsosqUBL1s7qg6kCC0IMn2cxh054qirbenr3
Hm7d7+w0GHG+VLM9ZKwGBt12ZlfFE54No2SctfXu5RgFklMIS81fb6pdoZFMuYg7
HkClZIqzSzpZklqYYvrUx7HVKRpmeSiaBcjmLZcpKrYUE1fr8OuGxO6frUtgKIKo
uk4Or2TzgqtkhyK9Diu9TH2eNofmbjKBv8VDo8h3pPp1TAkxxlprg4txvJ2lmum8
ox/Vqes/DegpcPEbtkWUS3sgUIlTZotYraQxyVhFp2IuZ5jd4QW0gQnDMhs2ypAB
MpU6xCA/PG1hIyeLdO+l6hWkRUmKWZK83TulhGMhc20A/74Oz3CpePAws62KETRb
7bo/pGC3WiCLYYHJ9hFQ1AtmMRIORM1NocbadnjkUZCsH7/OE5eKKER1Xi6El1tA
rpNnWOh/MLfXxXF0uyl2wlN+Y3G1dhOImy+dL7cjUBJUsA3IUH6vr72KJNAihbg1
j+k1NXIlJMs3BPjk7z/fIS2I4hh92hkefpiA1N/ljIRHy7PK/wkWczH+tZo5ro3g
pYuZFnypkr00tnYOhoErytpcm/8Yj2unPtPSJoiAWnfKb4soEZQOSwUgXV0cdknT
Bivtv1pymt97caZihlvk23G8zKf6v/0gx8e3SOpuzh6mPmSzq+aptcRfkWj0a7e0
syqpsRrQck0ggpRIQeU8iAOIEdBBUA7bcwGyvud9dEbzkBKRzfIBt92x5A/DBT8P
sLQdsi0dWC+FcWR/bWtjRFl6GzdazQ5O0j1ipoFgd+Kxg9seDufCh10gbyXhkL4z
+nZl0fzwdVjADYDu0UcaunDOqxRQfyVq9tYrNvmGJw9Xs4Y38VeKpKQ47sALYPaN
R6GsWhOjlVhnEls3mVjECnyaGyW4SwPOeOKOSH1H0FrJuvpdL+kY3Eqdf1NZnMNs
QIK6Bv1GP72aNdSCAmZte0cmETcgX7Dgoba09kyhi2dxfc5pWOQQB3/Yqvxt1YU9
NJI0RQa0WA6gjDb9TeO3zTU2BbvkGg4OVQ4nWtI8GQ/HRCvfuSyAywCmlWnf+J8O
7+6pGzXHlRAyItHaWeU3OxQFIC5ozLyVV0EDK/m/tveUl62/9CcNL4BphgUdzfx9
4RegwwGVd2/kGaFPt2RECB68DBvCFuME/hjYB3NczRcjudZ0Xh1CVqdPmpgTzRme
TayAR8M0rZN+XrtNo1u7vUWFjDaT2+av5dTgL2S4snaKZld+9ZmXiNQgmTnAHNBB
foPbM8yZSaXwpdoogMqhQwAsosxQGf9fvSFf4LpnulD6LNvNgv21lUUsvFoQd66V
m8M6kod4TjiSKt6C9ib758whi42WdtnpxAKDDVz7BS/zaWAFD5gH49HYBU/de8IO
dV88zB1MUmFiaHnu3pXwFgBihFduCSPnvWu6qMLvBgc310nh07apsdJI/H9FBoSK
w1IZdXO2Z4Fpfl9+nS4ri90Nkt3WBtLU6x1a2SvhkbOeZgmklNyf82sU3mwaS5pH
NE5unlrUKjDRGNEatO1gseC5BtdVKxPs+EAPZMgEHfbwSAqs7q6r7gjMx3EqgfgW
npPQJJwPQyyKm6GWI62nUgv38R/ztiK6k6YIAqBOWKN3AWyEoUUkRjg5+7ZL2v1C
8AqDyjVQEqJh+xym3qlNxGq3cBAx4Fzz9pbgjeTfLYh3QpOqNbT5EqQeAmUhwl7C
Ezmk75qVdCZWDa5oLdXA9MkJH/KwvSCvgk0MX4/+GnTY3HOn51YHVxhUbOhQI2Rf
AxxOJypONVUwsHgJ3x0gHYLn72BVEWB6pF391KqC1mJwemZPkDR42vQuq15t5RMD
EJUEzGNAsfmEfyCpdaagzm9R0dWAtSUXo5REvxJ7OHhlR5TMimcqeuU3S/TWKNTE
PMAcMRFWMEyMiTwO3/khCLY96wSihHljtdepsQauqKY3ztvUnKXocjqMhf16cUDr
o853zf+sKR4cLFjc+vjTsB29dx3v5NRzoKeeFN8t3qtIldfgVUOAVB5CXEuSWvh+
aQnCJRHuJ3ChQA+9IaCxex66Q4jYre3pznBQjjPfGfE2oZoS+d6UAuxP2bizZZH9
qlj2huKSA/Zs1s+OgTlzTt9Tu5/DLDtcUcdOjC7lCER2MwYiy/5vG6scCMHLPC3Y
EiHqdFBMHXX/Jru5rHlXBfhwkLUZmYeZWh0OC0P0MCuRPM1C9oKRd4xW0IE+ze+j
GY1gTJeznpJW13flw6hwpdwqEimgFYkwlNidttCWaqrW+KOikSuIlFHMxb9IBYke
wm0rsAp8Z/l9bDAszK1tXtV2r3B9+niqJScF28KucWGOpp8QE1QhHHCcDwtON5KB
7B0Agp1SXJ8JIiaGTj3wKoOocWmiASDy5/Dpqms8zGI/1WhVZjsi3eS6mIXfP9zW
3terCu7Bif9VDNvj2uYVkMnIPXuhEOh0kklcOgqYH572LlViD98W9dQhxDN96Jf0
+f+wIpj4mfw1rht4LQPo4NOdX4HiqI+p4z71Ppzpig2U4vEplFItLZyhWh6htkMH
XyCj3H0dFXu0b69UHPefkvJox9VGlv63YPl0bPK5Qw43on6sKROfiw1UUt5QUtgR
mttJYyDDWE5bnWZvjDYe+EGVQ7Bf8pSz+gTy2kezcFQMSnWlhCB7GtZpmsATcLdJ
xbx5iwnAaom0kVNDqx6UhnXOxxLWYOO6s5S4laCIAPw+SabWlmIxe0WPLdTBpilC
QWvIcbT/v6S+2NnsZL131UBymaOW4a6BzJ9zllEzWpa85WLLCpB4dZgRRkLJLdlv
052zzkZFyfDdcAxiTnLupPGiqk9cou2I6fz6pGNu6WxDnMkYr+tJfpqlNraXJnO+
e6Ygv1J/BDLKvs1+N1U4DJfzpoPWAv8tNIlQsoBRfsHiW5w8WN75uIL00LFkK6I+
k5puFEOW8fa9GQ4Up7SUnF211jqHa73j6S+1kC9d5Z9NJcrR99ZIg8fnsayWupv9
eZ35qN+i7GN2a0PWknuBJSV7hVLrsdHYPO0tz4eat7BBgHDDsKjEaLz3iI+B9obH
h7dFq1WOWRhzCSUBYwAFDOrWTosF50gMUP/umWYuh7+jgrY8UUnGRg8vk0GcARd2
9gideVxjjbBEd1Irzi9SnMeOihNQEpCf2ezODUtPvwLK9Op+iFOQ9EFHlU8K9SEq
rAnUJx5t2Utq2SmET9AjkkmSt2Cb3AbG3fbg/J48ImjD0Q9U5Q01z5sD7a9KD0xP
ComUqdeazghZAuDraCIwtI9x8ZHkL+GXecG4yhX3YR/0URVM8BagGOZiRGBLsc2M
bGzUyOF9xq73S6npEpyZEp0tg4JCu9u/Mjbhg1optOxhZgLHKbUoGwAIh2jLdxNX
y7hkQHQdXPuCyRduj8F1gZ/zO7SCwdKK7n4+k8+FYxuJr8sdZZ8vhX43Znku74Mt
kDZ+p9q/e8ok001ouaA05W92aYhxyg2G7QZIOiBM52B32xFit3T1GJjUXxWLmTRY
esPT1ffjpPNEO0vX4lF2sCt+VPEg++03Nk3/XxN/d4w7H01zqkFkuEoFHnTR/aRj
BPSGj0fUaIZ6w/7OXe/q+uJ2MuKn3uamcL1lSnsYYzl9ZqduyVa69fyW79gZoOWF
fJXllDKGmsGsHfnNBU/YFQOFf3uEoLty/ZoMtgm9Chry1DqjiCGk8RiipMtKvmrE
mMS4ibsRDZGWZeVEMQWylc0pW5SMgL/BgHNfGINYtTTA+68FpHNcOPBMSGb1PssJ
mRg/mcp6MNFZ/h5UMngVfkYJd2zBbqPmn/GOGn1ScPVQdgQo+tLRPWmOaaQxNlmo
67C/bvWkw5Gi+lAnSgLptsXgwpnYuDbj5iLraA6bfy8EBysnSxCftnDE3so9LgIy
D8XcV3IZz/p8mjSbfcAbbIrWhtOPJS8wjqja1I5UAdeWymxoD/r5YeMWygMm9HHx
MYg4O7CBKWgVsuIktHJlzxsIr5QTA5jzjiu+nFthbCp+JxOlVBG//SrArp0OmDC2
ny8qlKwEwP6XkvW39GFkFF5sP8TaNWxdl1xMQ5pTGb0kdcAq+BIh5/xBeJvN1Nqh
GXpgr5/+rCqbyxG68nQEkGydIc1BlkY9MZwmAGjQjPyB95s1GBXKli5x4BqAvZ1Y
0MmpVk2VgX7Tbq9E8c8VdDBQXaV6EfxT85dFAI5cOUB7Uxzc8F1cm7ewd8WdmVli
absJeGcd38eukpdgQJV5gRikK2e5uhAdWBc8yHPEv2X7oKsYs1+Hbga4hJq72OKW
Xg+2aXgh3mPKRrPPBLkJJ4aMnCV3V/tenfHfUFG1CtTTJMw/2T/H30G/3mckGUds
tzxNvwwP6gskbwzkIcpB+9eOYY26N6KBJ/ibxsbwpZCMqsQkg+K5l641sBlhlWNN
0A4o8T0qlISWx5UMhUMVKTGT9Nkst+Zv88qCVK6C7dn0KQTCFHKavcMr8OypLpov
Qu1rTDdaFNDiGGMHj31vlUXhus5cRIFsRAsWH52Ub1rnG7mcs7FvPw9HfjGu3Gtf
jnu4tJFxj9Klw7/AYY+93yLUux84MF1nLcR/CLf6mkmck9Uik05F5subAKkfO9eM
BcO5oZIVsGUiOiH9QhNLNtuyQqAMvEokWeMWdNnPjKI3s3oU8kQZQaFwF1aYhdZX
+1t1NfPoGi6hETTnWoMSYwUvxug/vp3XKFTpG635USVcktNHfzdEgk7gF0j0PYQz
MUxzqhEvOSbsxwlzO7kn0OHQfpQn6BXduzyPgDMMwmHeD6IuLXlPwtfS09QiJQSL
hCyszytPjsuODR8jHxgjgtoDx6fsYEo0F7nddWLYN4o4VAn27+xD+bOB54MCkS1L
W27w4WJkcYAqlJ71iLW4H1AhK+k5LJdzAI9QCE+mcoZDl1Ok3pt6SaipHxX5qQ4z
hG+Vmo4a5F5rMKZRP72xsQ2ywIOOXSv+NPd4QIjzLBO7dynoXg9ok1mFXkhHAzBW
MdFjKPcicJzPRomZ9m6CMxJVRcX35oAsxRd1yELn8O1R873dKDkhTdRrRIe6z9Uz
uXanc0mwv7iliv8oNtVW6XhL3ViE5X7AmeDKXNmL3geixiZpk1Kn55Wn3M1yPUvT
HeRYnf4F23W7a1Iy+g5UJEoYnpe1n/rHu9/B9z9xBIHp18G4kKMnkGktaGicYtLk
kGl0Bno/vNCQ+beyP+tX2TOkxuK3vP2e2gOueM8finYactvui50LwMswhb7MhLHW
wCP5uhDNCCksdEsEwzxvuOZyktmsIXCetFimQ635psXkw0d6J1o3iSMVPzLgrS5g
qJzp+fsmPhYYI2Z4uehidbJUYxYoRrOfUHlEVS2yA6WL1O4NMgbFUc5j/llnn7US
MmkUe5lby4a80BPHtoFQUEjWZsPFCNpwVVMDXlLOmgnYjnfMXVamcigack/OQX6N
2yK4njc3lXh7UBYTRMLspVd/hoxGIbaS91lKvQxqzChHrwYf7CY2zB1+ICegjFxP
P+C6ZcWwmyCQyF1gMOys3+QXRL7ZyM5egYIvEiSjglpNv2sZT382fjYBhW+WMU/7
mh2kuQlgKKzPnW6qWIzJ2p4667eH1IU7eZxwW8s3YKOsYEuBnupsX8UOfg0n+diY
oDyU4jKjlzEGBFp/rgESiqfKeETL2XMFMHN33wdWf3Pz1s5f2avUkHe83HGdpfbW
vsB89dNMMBn+l5t4YRdK/DcFGyM2jw1C7poH6JGSTLFrSsYUQhW5YepJdvUWqOjW
iVBPqEc1f4Swii56vtnbwXUWeyWjOqH3IS2qsrhi57mGpsqhI4DO8dUhQ1cbkRwf
Jh2F9qZpTm9HPnN0AWv9JikcOoqPhg9vxgfh5fL2RQ9H/K9um3pxyim8f1TRZoqS
rm/BQyt0RTUB61iYdANo34RGZb+RlZXJwPN0amAOlBng0sOzXRenNLnaosbijrdt
2NSYQolsXkG3IzuRwUctJMJjZH4fWq4LbfyZPTA/ugTcHLBUVvRnxEVw1zvgqhra
CTKQWdLqsxM8qwnGO/CPEmQ/GCs1nClo5+TdTayBk3FExvilTectLwH8+goTFf9f
Mkw/3fk3ad1btkSM0LxJrxnLUZrtsjqVAqbvhT71KOnZbcm1vJhMpAk9ZtE4qZMd
47vvAJopZY1z5EAgJvyhtroaDEyPxP0r+7e5V5AhXgi6rzItSpDpPmoxrRMRFFbb
zk++HLn5f6qRuhSeaqlNhoo+caw8iXDpJKtjjOISPbkhcL0HbqJp4O9pcv23kco+
D4k/ZhXagyHC3jBzY8zEGgIn6V3PSvvQFs9M4tbeBNSfauNoGjYrQ6PBGQ2+LVD/
VjQJP+zDNQDb6WgTu+00j23StKcz/2+4sxt7PsyExPl86/qIIYNf+szV9NR6tEI2
H/OyPlTuwrafjrUe4TDgvy5UBtOCHL12N5ZzEKVdMPL1OOYetX+cCkm/QVVOPIUu
7GHkgSPWKAUNQ6elaKIY+E/CueBUF5JzjkF9MoCAeVpHyb0w0K04qqZykSZjfzEc
VIxYD8SQLftFZp2HZjUeA/YASQaZYCb+0dJiyZ2LjmCIhLxPs9/WhGdHy++GQMux
F75AYDOAh5LEK4TN+qzZvW8tRua96HqlDdXopVHxu9A1MIgmYaLirccIF7ZToycu
wNryOFDUNoobXChQZ0oBwgNrkagtvXPqQPR8MpuxDLgVfkMSOaL8mQwbtG0JchFq
LrPwzVAbcZAERvNTx2NvtTZplA2Tw1wK7/gF4SGx4+7llstDFPgq1FZepvY7SpkW
R2HIEhqrKTIsx4HdwysfcyWOgIxPu/XXDC+60fM87f7ZmqPO5S3jgtX7adh62szB
b3bmwk/qfgx4mnjyHi7r5tic3AHyneKGzR8yq/XrPCJjdiM8ZtKGdOSJzL40YhbZ
D4Mb1rLYooclWk+G5UcYoQigBVNGiv4zovjHWGOJrl6Ep6vhSsV5MWgdcshvWvFV
KCv6VLeO8Wzc3qt+7pptRgsXjKHFQJhY1R81rs6S/YhybiNG25IOwuywzPIqC2Rt
VHjRS/UpPVFTtjtswQJVQDqV2uECYxUQvBWKeb1Xh2HmiJE7c1h/pEj9QFcyFgnG
vawIh1sV18knDtj6zQIaEJDUjYmGiGv3yCnk0xDIX0RJaZRKcPlUWh8Wa5X6MZrm
n33RERZeO2HiKBV1bQg4PLpPGZKD1ksr9KC6Rj+IhkKBT+9eCWuBh7b/mPtVc9FC
jIujvkVqcCccdNUyPpdVuJ2SzVX0Q2qIcmxoK+UzlKMEJL1ZOtR8V7cwAtVskS/x
qAaxbQ9Q2XQiCMqOW+vr141ph5MDiCMnOGPXGUVUu+k4TINroFnTCxQKpM2d9kfz
m+ngyVns4Fqxuss3uMz/ZyDMDeKf0QX8erkPARz8SMN3BMLUlvNWt83vwhLGVKDQ
GHWG62kuM5eN8qtc4Heel/1HxKHvLx2q8ft2jU7ip2mG4t+Kw6KJ4u5Fq8wsjbur
TrGt7moTFo+xfdtuu/RMuGlD6VzNSMfjqce3AIQGXDaN1UqPS263CcnyPd+1wsi2
vNto5O5Sd82SoWU+WteVwPcYuoRCWArLyizm5FTYY14HbU/+BcJNXakYQzW8wGyi
6lRF6M3x6bVv0B2+h1SbzMMJRCT580OScJF/8VGwofW3Vkv0cvyaWN2ji9sR3Jzg
8U4D4+2WZrVCiX+AWnXc5pz6akGVe2jShjdWkxcjZkvd099owrplyk3ww4VPAu/H
JX5Phdqbc41Znc9YpWJ8n9tPQO5c+S/wWmAJmLEQk9a+kavJQPJUrVN5aZb6HbDc
UwGGYp5bX9NhxHQpR8wim3/wXsFMIDgrP9Ww+b3csXdPMqUyAn5JNjzrZXAvc0oo
nHe2Dpfw2ACkvNyPEajT8g+KQSzF/qoJhffAMw/i49r36fyd/coToiv8qy0wAs9Q
wYSkffeqxq1fZZSIjqesbBJiGAm2tn+UCWINSQH+1lLmCX7OxTzE4/Hvmn0mpjnQ
TI6uyE44E+QPdrK8Xln1P+k/4vejSYhLeC3pMnQVoX1cPVfcBp/AcJc14ly7eGvU
ixHJOXCDf7wZ9VS1bh3o8RGUSpjlqnPwaH+xxepY9640hWB9M+HyNl3PJwSUat/h
Z69+0NfkkgVWfOdy5K92w/Yg6NyQx3AIdFbvAv5eMMbr9vuWwRVp6oFCwzyxuSGg
4WC5Ig431gWnkygaZPTPB+r/ukg54qqrwccn4WeZmYWF7IFkigYmvY1JE3iDI6wc
z/L0niTG8Tz5RrauYXBD2Tzj3DA+iJ7pIvc1ITR9QjiNQxnycpmb8J0G8UZZpaQC
RjNv91vRnDNkkqpqFxywHof4Frf8VyKOztKCegtfvzlPdAyUWxDE4wi2A8FoRwBk
+Ju3R5kBP1C03wmp2TE0dj9GcwBsXD1gBCR1F4kfpjSJTOWunIqjZx44CXeyIflv
3eLu+IQE4paMjoz6ZpmxemonisBKFkukACvFlhMHCCpoLOEPYfiM4IcBBVb17pCv
uPvtkOTAP20yVFls3dtsVZqTEGjB3ezu6gCkBPuAaB1+b3o3rMZds9zcbYX0T33p
Ns95WWfAL/MSBR3LQlsL7G4Q9aCaIARY8kziHlJux+xjmV+DbmnN/E6lJ5YEGN1I
RbYW7HlkU178w0xcqQoA04To8VcPi2nmaMgtiK2XatNKxGTRZyTfT6863g9DDKPY
mjsKKqP/obnkMS4T6MOPK5JEcuhen13G3WYUEOAfHbilQYPN0we6OjMU5f9EFhBk
SDrm+gE8zSmllNbjxd2qW8Rh06wzCDNoRm4wiGyZeJj4ZIiR9xqZUTxziTBO/qY2
OeNDaRl2YTth8s89vCxNKq7sk1mtC1+rOtAQlY+dG3ptegsCLVl8fepar4raAD+e
UWy8+6VI0LHtqZnbHYGBOKAqz6W6SLqzstxKWKM/wXT8MtB4ARqstDOo5mE9AJ6N
8Pw0VMQE3zOiMH4PKc23e4KNybiPe/MBlOADTA/BLBDl9cVWo6yoiCeUq9W/6lVS
Gk0IBH8xosi39CJOd8WLoTx3SX7jzetRskFkmosobedYRmlKvHOs1zv1zZ2rhzou
iQI/nl71PUFwDF+WxNF9hXTi3HHXDgroZi3dU0AjvIw6YyNn3XCaXMVEkvMQPVjQ
3IjYS246MZdwnuSZyO+pfYXDrZpTkd3/xq0sbsEwhhGGbIJ8HryDeszncOegdAhV
ofiyFpmLNaJv92zRes+pSsL7dnaaMjESk8TOOrDQQ2ODI8Ls+ErvcnzNhftGTdr7
3o/YerbBAb37XpTc/1ZTUNG9X+WvZMsgbENnL1WWv651GXXFMTMS+Yq38smDEfxB
ZVqv/5HGc8fg+En/iqUAu4EEIP0t5fcCBwbcdWJZ8jC8eXiyiYZtg3HD/+PIx5f6
VmdRoFPDX08+F+EDMBMBHYRCns5th8pFGlfPezQpWDTTntEYZpHDIrQQBvmBSDf+
FuUWW2tqu/eU6mq17k7Mo4j/RcP/shEBTq0g3GaQSKnebgW6P6CsJd2+6hkAsuxy
UDMUJpodAqjQu4cOoiAtFRgVs1uM25E+TAll626dzsqIyzxnwrhWBBaPCgc+ywu9
f6/twZ+MazyOHKWH0ndHdmEdeU9IP6hgTWQ2kRDvYvyuPdiHVDQt1NmlZySBxxwb
49CCasAUX5IbHaUQ/kQc9jJhFhniMTCoe6gvQgW4OupFesMEKTOXzjP75WKmREBL
+6fZyHTtwj25NAP2LvrGaFRmkgSsedyUmVExTngmP1dw4sjy2JhHq3WYBPWDxl4S
SjSiqHn0y53gYOpdVxRqgJaxh56Bmm+s1VqLQdrN6duzT3BOR2G5CDDy/sPWjuoF
wHZa7MPLeaQ0uVfH0ZTex4EDqpK/Mv4zQkgvw7Jww3Y20eokUwe1LZ+G8LeVIW//
wzzx++vqwRcvz2S0lR5pR+ZFzrWO2K5HT4jw+XNYwamhqXpV3vL00GE+c6xrophG
yxvVP9aJ01Rp96uM1rhlumhvhg2lWOSWXglaihmNHJWgM3qs4lRHOH0WslAglnEu
nIlJHYG8KXgfR1v2I2XSMp+Mu20fgxfR7qBXg6MvTA2Vj5IMhksjufoGrj1dnCb4
zzXr7rALNJ+BI5K0pFofSVvgcloaoUzMlJ+hdmW5WYSre79I/Fp5/PvwS/yNJ3fT
jDUWZJfKLLyCygn3+CDCuupzuUN3s3DbwWfb90rnhOj5oux+LHqZRKc08PHHzjab
+aktxpgMAKbJWdKeEneuOTVUApgCTLc1Aq15Li+/q48Ba7KHL0BV8MD/lEABuSpB
UEpcaa8WjeGjoG8CpBWkqbOUOyxvNTLptcvQPi/5TjsJ9i/1njbGgjUVCOaQco9A
wsd8xg3LsH4iVwmY3Hf8J/RoE/J5u61mtkoZm7SaHy0OunACDPdXj4R8L7gsrUjV
RxiXeo/HSR28XopHQHFNYT8sTEVSv/Q9NQ2Ni4hPowEH8zDMfC8r1MaEzLGyj+gk
cAFhBH9Av1ELVq8IH9fbu+9dGPBOOJQPhHVOV5CC0d45Sd5DwSjX7z6Yi6oLadzx
eYFfs6lwCx0qBtQP26/rONL5AT5SbTlvohgW4xG6hnbcAaUrPGu4+l9C+JIdhNNR
nCddA3XPcLU6wnU5D/kzYHk2b/wE8xFpgu6NfNVghrDx3AIrgvedt47WV/wZEqmF
P5iRNQTSriMxFrt9rnPsLOeG0HOHO9yTmMPk0ysXkSb0dPYniXg7QPJQ9+npUOXa
McZeg3JVDv2BmF7dTKaS4TvqH0ODbK3Yl8bAaHiZj+5XEHjrtRZppQdnT0D5tc3x
fxhS2/AK1RsX3BRARM/vlkrKWUgjY0qYF7uxER1Gj9pi8KdK4Dsq+nh+ifk+gNIz
Qt7Dhri5hwONSUFrr4YtB9Kr2aZrttwMP+49DwV9idocm56xrLacnZKVBeGUs9gA
x+5fmquwp2tLT8CVmYXU3MHJOMsjyRkNi1fR+GUpkIl+5um/pUyleJsdPZ0Y7MXi
w+iRsuhUDd2JmWYagi0dQXkN5UowQP0hldU+zFv2FCUyfSxmZwdrV+iCQUriKae/
pzUFy9G31DteVS3PzvIl0T8qo5h3iJje58lNJU40Uc2r9qdnAtkFCol7No5NHQEv
4+yp1zZcI+D3t/VdKimN2MRJQYDIYETmjvoEC0xiSuU+AZY918TiUS4PIw45zF+K
yaGWt0RNzjsVlFrwdrLPYRe9S1mzHAkmGUfhOMGmKmPhjgvPN5Ha+24ui9GQfGrj
+bCRitUHVy1R1IwlY7+RLn8PezsEhxaJbfnexPqXitu3JC31PZ6Dq6VJ0BVmqOgT
Yz33WFcUNedf3AXgE8FxPwaYGkPV4St3oYttClZ1bl5kmcvGerB5RpkDWT5UA6de
dBjgiYvvVcH9UEOrnhuUW5h7+Dv7toWJHQxyk2hbRrWBTb4PJ3eTsJfkd0z2153R
8a+asgz+BO3Z1vOmD83w004OKhav95DxmxUSvnWgJI/lGZM0SmK/2I27J++1AVmy
I6Z6iqop77hKWuJpv+ILgtbjGvCWnFEtehDgD7eeqB+KAulTktSFa5Nft0JqlaPv
CoISalx1x3Wwa6W3feoqW3YeILgP/HTRNTooTkhX4TuCUoFm4xFuvsIk4LoTxc8V
1pBm//glxn6ZCTYjSrlgxHrU7h6r8sxKrpCte+8eJIEB8ccmmTlmx1DTo3ZAoWdL
me2PcOsbfdJpYMQGoQoEXtDq43kIZcJhmGcl2akUQNeLBTrmTKQuiO6fTF7Vesb7
E5avYPHlMvgxm3/aYrQV1h0bMA1TgWtncW4GmIpTuFkxI7Hq/gFP5hXtbtjR5y4e
p25FRCrbRDNTgB3VgCJ746sqnjBKKRxyabeuNUpoNSeo2oqKRBQ/2amp4l/x4JXk
/ddnLiCHOgvjLdZnfMPywl1yyjpYstnD87M2lcpt18CKU2+jxVCMIICzVO2eXR8c
/cgc6g23OWgEFNA/i+YQU3+RLp4BJhZSpwV5ZqhS/cYgFXaJ+hhi9lqPO5JMrpLv
bIoiwG+qnkoCl0QG9vUQpIOIWJlstVc8oDiJ40qTsPheXsud8bbsT5Ei6I2ysIvl
lJ+CKrD1iOK7TT7UXRC/UeISZbdLwRChrBfmcDvudLUVzGZxPLsywBpP1aC2V2nx
uox1qNVWviUgcU9slbT1DFG1VwVC9LbnKDN2qikUyyf6TNXGnPjBB6SsItdenuJt
dGuyEImoTbWTOk3X6nE3IvH2mCblbkT2mYMNFW4hM0wpVeMrc50IhQXk/OkUU4iE
ByBNx1RXOJ4oEEnI4R/ee+26YyXCkGtJgczbHOjTcWkXNKx/bqEecc8ddDtlmLkz
S46xIB+fMnsBKQV9xjJvfxN7gpItUXiTYvFcEg/HyWXX3HRGoK3uMuvCUA28tuX/
5l0MW/EZ2xbPgtPgVi4964PF+M6dts9KTKblgbCcLOYUXM+3OKFxUe2ALc7tOw1e
WZeaQltvGwIf8jQzLR2u3vF3ZrOx3oX2jFMMLAkQknUbCCgX7OuyyQ/ldWzoF1P7
a8uiLJknJelRcqP2gBVcqAl7h9R7zENgGERVmAcVizrruJeW2purhubl/fprx3VL
8+vlkN5SZrjyne4lkEunArzfEIUAJQ5bWcBkAmXOGyM1tCOsCtVvMROVnhO20KdU
/ZbzwvYTu/ZRU2HuwafoCCv6VFKozl1IBEMxStCdMRRe1j30bOJ6u7dntdfIO3cX
fUUZy5GsEHbLqNBYBrH9lNxSVoQNepMclivnRSuqjWBXoXkDOt5jyYDO6/gyt4Jh
dyZ+mUxH+6heWuV8f5c87dJ4VrWzNZz6nSxXplED4TtFFGzkwByyDCM7WRz4sIDg
mF3jGCOdl6uQAPNKuxneFiuIvbCNnie2QzZDU4WaBEz1Kly1uPoAAReaA6AeTfQA
DeDwk3yqjBYxU4TY58goLOqQMD4QaFXuYOqGudCFwfgpGXQNpIIhyWY+GdoX4gq8
WcuGl68pdqIctWUyROWR+xRsHO9hKihcIzxfLr9xqzHmWTA1h+SVElUjoJ4lyrKb
lYDMM5AuFqbSDwvwQouyk7kLbzDCg+slFybgNeBUrXdEDxXavdAw/E0GMY3yN/Ba
UAIcPSdwns3mq9IFMy7D1pjlU57hQ1DLksbBd0xcgjfAPuuMBoxyRnl+zzn/87ba
/Rz/f+LNQ/iT6O/jPB56PFtubB6wZ36dzmj+jeyaBL5D7fdWAxbUjS28v/WlAxGa
ue+Hyb/4b8qj2+5mOucWJdProfWbedcLvBg+Mmkp9RcEmDPyeLSSpIFK1s1lmnNh
CCfoxntc7tRhXaxt6toSbxn3EvycfxxdGbZM+RcgJuEvH7Jr/s990RekjbxcPRBv
/H+nV5v4pMSnHIa4QBNUKndTEwyeb+gG7YhRlS0Dhxml6hl3AObuq9bglQa4THBP
EJkzZGK9KAPQDZICaW/URB/WFwJeSjRaJZAxwmL1HeeCmEEvZiC6rPeRtHjL/e53
HUU6GXmtR0bAW1usYJg/M7YGEMieVK1BC/UuKavshXGSLMidiw0gEcFl9qbfNE24
Gk8bzf27gj3Z0BVUJsQKrYtIYHzwK0LZKkjkNZuip6HleZRb7rreKq9+917/yY9Y
C8BnfjDzhveVX3dCCTgb8KttErK2ZP/rfjktvAYZxMFDn2EDT+tND67HQRr4gmUZ
9D20mDogTm5MMQxclIwrhL/MqXtaY3xHE7qVgbHjLsTzHNLv/0e/E1skkai9y3kN
nFIXYNPW5hC5O1TNlEr5/Bp1zdVFV88fNjrDRwI3MK0ItKQXfd8Jsz7sjEJMTqqX
lGBRMPmQ/4366oKq46xRPHnd5ryWFF8eH4UFjT7mkHyPTuqN1YcjIU6/cRP/Go1B
IUiKgJ0g4NVVcedsuGiESDIHLhrrfDNr0BMxkSk9WcS+31Q2NMg+wJAx+lyRGtM6
5IqDRRE3u1DSPHnjiGglOsp4gdvQrWJ+St+Rxg/tvVAO6k0DXUkMMfrV27t65iIU
xFCpYbhVG8S5v60VRNmifryBjwWYvmPmk3Uf3wThYiPa32gAt5ls7axrjNKMIQZs
fEM1ira0hYSSlIa36FSsQjm0fYGVNGv0vkoxHCADWepOJzsPydsO3VZE8tHQHjnz
qYeCRJkzBxs1wV6r+Q4TUihDfhu5QmY5E2g16VCoswCvEuj+hIgh3JmzbYgnvnEy
AkR9vSbe3SPWIaXrQvXrp8xzV5AAi1QuAAJcx24+YKd7NLL9eTzHOzIJpSJ6mTaq
QOtAPnlLaLxiaVvvRSq4PtJUyZYSdMrJJ/E4Bex8lkDToMqC/SSB4oaxufcggxXM
GatcunNxTSezPtz+g25WeZFXRbkjtzJLfa0kcJMuTQV/vXCaPFJVwbb9dk3Zq5Gn
PdKCB3izwMpnE/GwirOklvCxUguF8ozFnkCfYLmXiNM7YhU1ltF5BP5cdId4A04u
/r4gQJPWar3mbxvc2NjhxhHmWdX0wrZKvx6/GfECPUQSqRzmehD9a6jI2ec+nbZ0
c/1Z2U14TtJDZko7x/7EMdxOPjYPdEbmto/WGvYmro3WzgiNQ7KVHWbpjdHu6vCD
b4Mw2GrImJDS/mOP0P+IvDgQv+fZORr7UGPIQdyWig5M40KXq3iSnOaLkmqMDr+p
QvabpNgXm77sGYMTloTpNKpDbgIz/f7kWqqgpa2kHUhxqct8wNgoKwS+yhoHoU8u
xHS5hJrExAjdSswBsF9//xqgVCMsMmV6mtL8gB9k58+hl3YVmnmLsLq8XPqo3cs2
wnsR087SpqDghbVB4VpopSd5MfTz4xY8U9wTvFGxzW6JTIIaI1yngU2MoOCiBgtu
Sti7PYwnNgRfDxKfAt2tCvr7TA7vgXpSNoBc4+T5sU+BxIUwgXIBQ3qtTe0wpYKE
+sFg1TMqpVwnN3jmhQoVGOI9sFW91/5Nyq8cPw7pmRmg5K8xXmmxyo023iFSMb2S
o8DlJzE0H1n/sAwkEpxNU31v+olkF+0LY9hFmTSQ1F5NhXfKVELmODZxd/wa2+8n
6kWsPdc9/7wN4kKnfUUnws6y8O7J/sKGovML0d9y8XJOycdZL+uZNwhsV70Gg3Nm
+QkKUhU2kk7kR34dEmDwxaeo5u8H6TlGsyEFFIAFbZqTbvW1nEK8JPoZU5Xk1/uC
x8fohq8yJKekKYb3O2QkIbYJivYPWbnnaMOXLRv02Gkw7Jhkf0EnHahN22M/7Fv8
jHYOM/9WsQxGpydGAYaj093joSWHyg/QRuN1x7Pjeg2Gg4Y9Y4rNWx781BoxP6Kj
rXqBNN5MO6mHKddJmNeH+CsTRfsNTJIw7+oHtucYEPMcs7+RKbiZdNTt0FfTULvY
EAhZcuM9Gm3WPRsb24oFJLb2DYy8DrczqzFiKc/fttkC7gjdTA4L9iXtkL9qKyo4
Wkhin0CzASTMmkD1uDrQtYBRXRrMoMTHk/yEP+kUrHS4pCd7hh9csqqRN+U9hooj
vrgQEIfedMnOfP3DzsHxnJzUX/VS3JDFTs9/yIF4goRnzEEC9CRIQ6pAFJ0Gz1ER
/EQ1hkk/wmsub+1t/gg7kjqF3wlgJkpoG7Dmeu6PLzXMH8nOov+QLi9RT27A0+RT
OYwZ5jAHhSmczn0xZC4oRUWHQO5P+w2MynIk8meT5I/NrbkHiaUCbZBl9voTTf4p
EI35QmeZz6AUy+uDOkJhPA/odJKRn3viC6nKpKwKoI+AukGKiqC6DlwXfNvWtCW2
ozU9CEBfCh6WvjowQyhOY8JqHs56MgNDJqz3oUIUrwrwlEaY8RCVU0JQyqOy0zmi
mehiDl7AtbZNyPqZjfzqCPMWaywfNUDuP34gKp5c5DGIvhZk30/LcN8TYsQ52Z94
eBK9PdBettyPaSBg/QKxNjZ1I9Bedo4SASPeXZflbsrWrwvS4A9Ihz+UlRK/dM0r
+VzEcGJijthlsTJV5DB1AmqP0MVz+eNEeLTcOowzNA1bG2xnBebyH0HtT2MWItZT
sNfLnc1e10bIaffDv15l6q190iU8tgQCpMUsaV0081x1V5T47IcP1rGOFss1BMiG
1BQiobgg93hVKoemv6uWj1OU1TT8KvRMulQJugx/zSvjpqa/hOXh0+moN/S2xFLE
9ZksV2ds0J9AmTAKKcGZS6Mi/YGow+CCaTGiXbnl4nSxa+Od8c5jZY+uRShbjeIk
C37x9tkivwejJVR2b73G4T7+zwyJP+WHZOzYUMZqkvVj471S6s/LWrhrVNb7wPZd
F1fv8iGbeOszOGy9ShpqXT3oTiZFq2RUY93RfXEAfXghrEhblR17DARzGUb3KNTL
t1NNpia6PcJwUcjMWF6SuoZJyLuTB/qarj4tw+eGANt1bsTd5omkLGtW7NWtdrnU
pDtgq7tgNY6miv4ySBtEAqJ9PqLjG+5kVNkahp/Kz1V4gZUGSdkWEfZDTT8B64S9
0I0jHqyEI7yyMmmz2Fu8Vc7LhI7jwXbV9ic6CV/0YnT/DeNjKqzgH2riq12IXYzU
MA0QCNu7RY241AOY0OovW9HGCPUVDWNR+BSRwenYk2YJwuMFAXL+rEr/5jKqqzyO
qVmRd8CyI3IOL8+cEtjXs+vwAtq6sx4gNDQsg1XOP4UQBVMvP64HI4Qngh1OWU1I
Kf5EqX+ou1CES3Yy1EUw36Efo9jx0uiESB0CARIFCtem/dqHDN0NVClLAu5z+9DA
sRB8+w4NQuuZ+3af847AG8L2z/TeIaoZmNG9Lbs6DPjy7xZZro2IlGn1+lfhf9rW
neE1pMqNz0vE5IqyDEVRfqG199faaFqII9+Zo/v5gsuklVyJN9XrDue/X2w4Q7+p
PMAq+XGueA2md8aTsa42JX/0rAO+lN6u8G0FGMsW7RxRqdGCpnwIB7XjrS72C4U5
IpivVOyrNlcbL8xGbvS4/wGqdoXCrLvTgINtaUTdokXp4P56CUjvToC2H7H41P0j
YoRRvidLqyIVqsvn0muGP3M0mhwjtLseMpNFOsu/ylLNbOaSKb8YtBqw1Fr83V8I
zMrUbpDkK6sYI50uF5JIzKHwNAxReKNUQb+gQvJzhJitgqU454pTJe1wEEzVctim
wUpxgTr/lqAoOqQGHCGOFc7PZ1zAh8xhMcIorh1d9uH/2+DFq4o6kCEQQWDQa/yJ
2cIMxar8CX9ZXjkTkZId0vLY/wX82AIARfKk4jemeR/9xAEiBi0EMky00S8NErCN
Is+zf9W4Q4B26iu/Sxv39VKzizYPO6YOLSyPj8hbJFNQUhgYWceOBgGdCM6UPj+c
JwMusmhbbImWbCiHaoL4HxMWDCFDxQ0Q0Zm5fkCDu62Byomwzv3/A97w6An63GuT
kNXpo56bo8Pc1Qw6bZ9GDsMMyB+B7l2a62OznKjGZs6mAL+N89Dzab9/ZkkIwMtN
83KRPPdw1sLQ5MV5WxrbAvKuBRfJBz4ksz8cY7ZMujxX7URU/nFM32N+Ixvv2FrF
uPZ3ZOUKMepSEgsC5VFRBA2hnMl2at2XOkrV3EiY959Bg+PpuOaA6Ps0I1Rg9I4Z
fLfPAbQo5eGTem8hgAfkKAN4wWUvPAJmhTRpzGEBjH7xefanKy16kY8IgEZSly51
5wHt9wyob8vOJIEXYxQ4TDaCIUv+c+AfyS1UBZqHviEBUn5yC1P5dOguQBt4GDc9
U+L6yw3pkAozQCYKhzPFoP8Irm+I+f5QCq9jO0V5yM8VaiJ9DP6707pGEI8Oc5+6
bsQC5Wfg5IjG/y17Fu0D8We/qvX87pLU9LjJqbj7SMZK0zlS2GDZCfkh1h8NRtoD
/kfv0CHZXPLboK5e8j7ecuu+Ka2zmXVIBdAiJnuBKTP1znkny6hZ+9c2Sr5dZ0i2
CnunXA2mATs0JTrtDo5/oQrJ4MuH8ITjWSVwMllBXIYuR36AANhiK4xgvh80mNyt
gnSXhRi04Slu+Eve8xzdF0V2MCyZG0g5crwQsUI85JQnDszOCTYYzzokhwyjKanX
QDOn4O8sqYk5TmoQhBp+k2U2JE0xETRtk/NTDvWtZpo7WzTzAid4KScfrQE7vlmM
W5A3t2VSAXujJ5doyk5lfBoOLcfODRrLBQHCr/gQjSvzEDltJq2i+qwU3nh3zmGB
aXp+brS2pZEzxNgd/BWzo0A9DAnf6MACXKAvH4Y5LrhK10REMIPBprB+gzBPSNg3
XHsqak0n+0xZQ5w0a715GBsuckjdc+xhD5dzduNWEBrQrdFRcmg63Xm1sMSasfnr
ZO6aG19qKVM2yLg8bQiGBEZq9cIpev4YPxuAoRWcHSphg+ab6v3+qQd9+4IxjHgl
nXPHPATXxtjlh8jyir+rIw0jhzI1LVfED5EOznyxOZUQyDc7IrGaf/5T+LiNOcIR
pkAkgHR066xDnmI/vVu191ApvjCY4/aFXbMIWSXulYv3KEYjJxxjShAo8R8ysBTp
Ez70XkD0txA99zqRxAM1HovCHWymi2FkELbEGGMFJ3zFrvJgXzvpYNDJ5rwEzmG4
4ELAmY2yfkOaL3PRtH8OYaOmeIPYfeOSXLQqGji+r0Th19UhYCfql/makcSM/xoB
jze3FSGfHQZqiPHMqD6xhWKxI8MbecQoCZ3hdLJFog8wBGoPlIc2kU8Cm/IB3H27
czSwp3P4+rWQOn4cLX+bdyDUl9JlF4AClK9Cou75ZlLNEozdeuDz97MSfDpnPCMj
rxJuyoPbRH1D8gY05jeN3I6CKW0fuOD499qVZN13NfKiptYPP/Wx0Qa5PXhG+1Ye
vZ3/Z0CY8Mm1wtvx2nplstLu7Sz7ON70beDixwjSrmD2jkOAH8t3nqFYWxrggKay
YlGZjZWoD+kSLhbuLDIHEd30sKFWQ0pTnVfrA58DUlanjsX2eOJnpcnRujOaZdIK
21CNFCueUTAGfp7qHsnOkj150k543/h8ZuW9vq3N6eFNvBn2dub+9LLe3KTFn1bv
nhn/xZLKoLVPwjGLLwvowglpfDlrO7R/22R92NuuD3Xxh+HZkilNOLMeNr+dC2SD
pGeV05M4qRlSqynXCi0TzqsitYkBzvH0++qkuMZ1y9qlXaWoi2OE/fggJYk1tLSj
zZ52b3RwJZ3oxkjDsG1GGzeJK9fOWhmZ8nHAq5hRIpYV4kmpWZaI0aUFo/4IeEI+
n/HG8enz83cSCntHFxPKgE/eUTKhKmZdCU0M2z3flJgxFGseVhFAOjhAmWXyETNb
enVHSXNyKIjjRGIOr0azehpg0SR9nlCZLoxb7q4S69zxUaAOcDNjvejl3Wbe2eLn
eWBT9GgtIJvyDQ+DIpyRl+Sbb5YtLPyN+ZlVz3Qma1f7ZD13p4w1RwGn+PrH+Yku
45A4JYYiPqTe8vYKf6W6lkfEu5AtLboPfRquPUuhiLXBjZM8JuLNJf3KXTyoDngF
KnXncquJFoLEeMBnA0+tYwuo8D18VTHZCYcc2M5AcNN0e4PcJUggiGoW52lzXe/E
e3K9P51edrWBaHos9gBssdlQabprttVoXUqyLlxuB2Tj3U0hRq+dMkEughcJWwim
Hmam+k1TrCGXTnkEBFimyoQkaAqXLx2ULfmJPlvOflV9MamkFn3fsEvtEetuZwAy
Mvs9T/S42TzMuD73kfMHkbdTUPL0Owbzuwja6W8ey8LXJdz/U/JWRY4EdcPhb666
vgYjZH6zG6iuhd6KqqPLMd9QbGSPA7UCXuAIQMmgFEnMq+vD5eNhkeJURL8z+wQr
LA9BnpQFX8iFrgFHLYiGHBoCJpreQMY8hoMW/ET+vUj36/XkesAW4QgwV4mpMq+r
Fjt0Zw0w7wfQLZ6k6IdlmVkbXzwJwuHx++ioy5IteRbGoP3t69METmREEO2JVJNT
SQ6Jp+4XZzreipjgk7MBNwoxUbVmvD9D+tttImCFMyhp3C6B8khCluDEzCHC7Ddq
JO3Vy4fTrvHilzykOlONBUXH5PR54dKDny1UkM2P85oSyun7GsjJ6Ov96hZuvpP0
58wZF/zHfwGb2fi2g/Su31Ks+WLKGUJI3DWwDt7wS+vzSObjs4fBSey1skW18Buf
pABZUs+tWESp+hHw5rsM/OOYmANOeGmZY5ky4PkRfbWbMSINLvxCIHCdbU2uVlek
SZI2NDCKNI5LaXyFyX1BCVHuVo844WAGgtoaWCz6Qz2IduQ8iQVn8v8i+eGQbn8S
w0FWJmkWi20BtaCN89atmvIPVsbuklCbHDjTTgQTP/GEnuPp9Wt5HZmCce0UiO8X
pf7Ue9y1DFGp9iy/ZHyMnsbRYHifWecr2jlnvEu1iKr0vWd0kTRike3XoaG4Unt2
1+Gx/lNBZTgODuPf8EMiwewCeZWvzRfpHDONyMGEjEZAGjdJ02j4LmAcZldOieqa
kyoZDX+LCGHocFdrXZYsKGLuAGhskCw6FCs+mDH4DQsZmVEA/O8oBmSgTKmsP6rf
nASD1Yu/UvUw/0M678ct7vC62EEAtEqQAIvV+D2NZNdh21pNa9sMGDqWqru2eIY2
91Pb4xGXc9w6SX2bc9WQxrK1brbvJFN2RulfDYb3ebME/L34v3QxhIKYQddlSwXC
MnYLI31KLz//NqzV7P6dPIkNSehFGCSG8zUNodMgb+Ni3/r1V06CgIXu7dXSsAWK
s6ixCV7FK3AIU+X7I/WJxwNSFGyJ361V0r5EY4cZrDEA6eFqEIeIShxKHTA//9m2
sbfcdccsP3AKUsN/N21qlgkXvv+l3PYpIPbKubVCxIKS2AeOdxaiaApGfxa5cSiU
PUQnZADTBSX9wDKqLh9AWSSiPSZHEf5zouY0J4awA1NkoieQkwzVAHnL5sLUzA4H
trygZOchQOWD3A8ZYmmqOt3HCK4KmiTNuTFZmBjObJEgtZvpKchAUAWr46ikqZ7I
a91W2vuA0ZPeWlw7CIhUJX+ve6OFNY8lHpxbLTI59fmJjjv+nfloIe7/srLdsJUS
+vH5w6Cvpq4dAKEvVSdUOaYtXSK+UEKGhuys8zSGBhiAnyAtvCgLBUkoATWQwhhW
xc9e6x55Rs60GQ4uOybrw8tEW0MuHLKvmySS+FhTcmMuf44M2uvU68z+Zm7/bms0
D4vnCZ3r6fBovB89L+FjxblS5abtmxvXZmri6jg6RXb6Fu/WQByuR9t2cmegRo+6
a3m7yG677QybNwtdhreEjw8tUSGBztMBIJ/ICT+fJGYKP1yGcp7DD2nXvgZQFmzC
h1VH89eXTAjuZXWvwaM0e2PaewriRf0Xfubl6tkLgFFU/sJSoa+aD4MpvBn0pFjw
euVdpuWOqGuyCYhhdzkOSdXo4m/4JVWdFz+qb1PJ8ZfWNjXqZFL/N0h4SqtuNZT6
Sv3IqHEXqKhTXOnRoIu3rp6cZc8T3yQXN9KX0xL8oMFgCrkc9Ok7thb+u79oVwM9
LQtjCVGhQboUrvAG+snj1/uI1gRfFRH63c6VhAFu/iKBE5U6RoRKx4r2jhzNv9eW
UA8sVlIjKNGky0qK9iUeuC7sJmTv0RWIsjYYZwD4/LPfcMMfwjGnA3c1ARYrW02P
mySz+wVQ2j22WqF1pWapimIyq59UZbGwQTvxSQzUjLfkP8Muwvk+HOgGGDrHcMZ9
2S6e//Tr7ZJzwrqrISaGhBEUFziY8WdGkakPsgw7fexbcbrrfVk5oysFdvaqpTL6
Dfss/F5a2MVjzRhi/DrPpbIkaAr2LRqNYBS0f7XKGeWcpGkS1JJDoLqOjYb++NtT
XifxUJ75jypdxvYVzYFrAbyvaewuIDO7BxECn4BwJd29PiNDYehpyvFx33bTlQJx
PIrXEBJSYjQjJQ5nzXBtaRxWAGlo3yfsvpv6GkbBGHaSip6OTl7yEA7cGLVczMbk
I5Sm+/niwgpcD5GumN/i1bCFMUEcSE8XHYlKNqWvr4zftbXeyYJmxuPufgeIBh/H
1I4io5eMKVF9HUm5VgJ5gJdRicOmen+cNT9VtzA5PSZcg6Tt8gniMkGSORtuND+6
iSeLKmsE75jMBhK3KNiTzHLT2FcxuzH9yPN5vGoTzZfoPjrb+YXOfPReB3vfOYtN
N32USQ5A87IRiv3eewDFH+9VO3MSs1/l52JpwqFLi82+R1gzR0zwkihy7LPo+asC
sm5kgk/qXRCT2/lHiQHGwHDMj70WTMZS0iCOWliYCH8UM/1Fc1mBhmfZ15MlI0Rb
YLVzljegWSTdlC+628kiRzVDgHt4O4H8KGpNh5ZCFoH2qhaeMXx9kA96G4M1uT3R
UOz7b6lufMJomJKk6K0/wqqUXMqY/bcZWVW79sNuBjtMsWm/Ml47r1O3fgExfD1H
k9OWfOMbbXVy1O9X9A2U3zSQJ5T8hlRrPMKOUrFnRaChRVsvI2J314fHAu9QRhZZ
YIFYrWPCMdzr5bG4Kn9FqJpqcxRycOG80Cnkh/K2mjURyDFOXLYCI1zeV3D5RoMS
T0VNUbjXrABE1qeW23SXg5zX1C6gPrTVn123xTmRc0qtYFGYdpMc8y2fLfEGtJJ+
vFZbiBsKYbTDENMFufyHau1KDfuipi0nAcfxGg7YToTdwSt4sxsiq4poXhe6bkIl
/28Gd6KyAsmiRkgfTlVJbkbw8Xo457ZBGCFmBW2O4vnQO9pWYXxhBDgA/3fUNP7P
drPVppqwCbGq+VJgXp+Nrlp21r1rPu2j4B/h3vuUZGUrZVRkXFb9EC1jLuympMv7
FL0L7H75CDkOTsFAE5IdyjZPkOmrNMh0Li6ZEo3NV6IsaciFY0Ak9zHS4ZYdASzO
8xCiN1jUZ/5bFjjUnECWkIfF8+J3me7EdfPpn8xcymqempA3DZ3cdYwxrHP3mC/L
5gcy3VOaSrfsX/VQhKFrynbWxQn0xWTNCNRijLUvTSaXB0oEdqa4EdsqpcEF34Ak
Q7dqoCMYA+6C3VCr4yaX530fwtANV6BaDXJPQdDswr4b1hIMVPfz2F5d/sLROVDm
elOj2pcflGj67nZGalYzOy41eLoqVa24T07eRTcysrUI9vwod6r+6yu/KUxZpGc5
klnsW3nzwxj5rPWpvrmzATxee6AXOswvmgKDj6JbNU0URshfCM6GJK7ENYbsy1OK
6iI4MS+Y5YihPguIVXZ7xIphUlMjdaWlBffmwfky2WEcWFi/d9LCWpcWHXG+Q7FP
rm1YVjSEHJrxgjkV57GNoyWEKZzHNzCuVCSsGhAtVNWAnVZMgsfx/M/1/XSSO0tL
RHlqdeA0qS6wv6GEISI7PM76Yqv9kfXD2b/OmoQaBSvXRaJqjlTzy8RHpqZHyXle
+118/nxecCn9SxoON34+rzSjvr9sq9iULA3XXmh5KoP6afdZS8Su73cpdFup/3aX
L2dz2UGCa4y2ecTLZKpIHgsPPRnzXnvb8rLKBJdeFhpgEbIVpZVOvtjowF+pNTye
HjRPQLiBjEyC0EbRjzbL/88C0+6q8j80JQxUgQCfVEKt+7rM4eJQo6QLxtJcuILk
hIOTH6hDz24yoZufL1lfWBBjvCkhFkxpbbZyrUMQ0eBoqB4bV+ilpRil1ZwVFTVN
pggtMA/6dDxb0uifV5yrIU3t1r205gsW8Bu1uX3zN/OIlp/wP1BNHlKUFW+qYUXw
TxNbMhRAlo9bR79XHGV5iVzSsoLKL7/n1piD1x4HaQeUhInYLAYjMd8710BHagNl
oqvQEQI+M+FhNt3H+p5JWlCRV2gRvCAHrwlRVtAhIr1v3OfhV813dZNGqFkQoBl3
wbc6QbAhuwWcuMK0+HsZfbFTNJXFx6FcjeH2Kez19yFk6D9SI+w5WossVWrFggkI
CWsQPn5v40k/zzKatUHZmPF3Vt+IT4u3u+BlUHbgGcBEJaIlI4v3uSKGZmRANgEh
2PgJCz0GdvJlW+Pzqwri3b8vDbyNz6/W2PKfyMhUJrQ1N9mN6GHfSskRd+dPMUCu
W0ClgoP2g0amhK7hn1azW8gVBcJF//nWIW3i1sW9lEE6oEcml7pU1Uam03x3RidL
DHv42xWKGxcKXl4xLKD8mxuBvoSGFEC4xC6IBNnDetbiGTRTv9FKrtDiRjtR4k5u
d/X/6bBdlqwqXWBhKCKK6B3hbzDAiYHPCbInSQf42XgaIWoDxbBx1+coFymduh9H
df8npmL/XLvtDnOHtSQYX0eNH7QFZrKZkh67hn66lomlpDFeaQiYJ3UY2/0oG9QU
MqU9o3iRH6wqC9wqZjholFpfFpoDcHQiiLc7aCj24A8xnMrJssOdMOKLqAewkK6o
Xy9SX5wB+m10ELrOq0KMnoyvFhr6FVBbzWko1Eq5rxLPazPRibSjkDaNuXrsxwNm
h1SbtbZNwqlsteEZZHqIyKspccVUOCGA4hzpn2f2E1jiVlTk+P9clsNLw2N6GWFt
jQ7/ytcrwrKe8m63wZ2MyVkeh0m/t9GSUkK3Ggg/gb3B7KWf6yK5fMA8vh17JgPd
faJQZYQOcuyqMRk6rjFI6O7NflWs/YoPymE/fZhAH12dbDbD6R4LY6wOSYK3p16r
yztFiGWmN4IeYoMaDPjWiwrQ6LRBFsDwXQamjJVxb0Dn5yxBsEWiRo2NVMdhfcxt
MatM1Bc4/1sofXhwn3n72qX4PJn0pMZ+mIRzBPfWJ8ziChGq9KpXvuAdAL5BLR3h
snmPzhZsVWyfP7Ebw5OgmHNpymWdkNRcLTmuF8VdJTDx+/OQ2pcIL/+UJ/kxMxzT
2HhuGdSjx/5tvZuozBhJ346/s/NU+ylKp+LRk+1jEXHXBGtvn3zB9cgtP3c/5gXO
HmewiZXqznle36Ltf2Lvt4Nv6wixaLx0YkENa/2Jn8eaIjzicQtDpt0rax/ro0H4
Qm7VqrlDdb62JR+gLavoEoQELBKMg39qx3pnmww9nxVkuO1uPO3hSeEQif1OpItr
LZJ/pzzXAE+cZYZ8fw5DHXifUSxPUBU4lLMPTR5fTLvemVSbBXo7KLmNoh9CgkBH
zI831uVpx3r3Jixlun3uLuYuWZVPkbgwghu9zn/iYkxjNSw95FlwvGQZUoUXQ6Rs
NGvsr6InTH2kqyeTM/jo1xGY406RZk4kdbb6+VPLJyGJoAB8DbF6Vc8p8a6pawym
vwoZAiK+QSdre/qL98SoXhAnz9r5zCjhFmXBKCOGbpc4l4wPPXx4lLwlCckVSoPR
1/mNbizw2bU0Ro2OzJXFHWKGkaZa1SWH32ARTQnkp8SfbYO0jUtBhu2uva0Jri1b
fs3+PHmSnqU5sLcM0GYBqI8lxLFfI5fkgHFbHAvEAFgMr1etqi7qRMOoVKOcMTev
WGuHoO4QmIjD2t05+bZBFcnVTHOi795E4yYdX8S7nxSGnRwvLtCG1m4Vn2WoqXLv
nw3+AAewY0q9w2wlyHTUdrt8t2N6jXxP1UGvT/h6LD6HMIzvnMK8HnssyV1kZzZX
2V49OTPQVQxvgDH52qWQoQh0FTxoaVGPL3sXKDjVDc0q+tU05KCUFhdUS1lpKUyw
UjxP8OeEbtmVdt9kRU2eilDHTGwuHShod6RD5aOsIvAWyHKYRyqtLIDI8OaDtOfw
t4O4bztJYXau0QIsFHwtlUL05CLF8i+qkiawcmdb1LIX28dpvQqsvJFE33RlcsFE
noFWxQtkiziDUcFI8hdXy/PQSt1AvzTMXYg8Jcamz6Le/Cgn79k1FqPgrwxi1Rwo
q2vaxU5XNneSuwp/DyYJvCxEdXgWMfSi1PGRz/uJhWnSWg2Wu70sE7/dvlMVe5aJ
vtyu+3SwGWd8KoosdcJGQlVKu/GbzZCAqD1OhKYGWL42dgnGElQfDfTnw1Jg7law
hhN6/4jlmOEHxN4K+wMu0aMr7eV832/+Nc/0Gc6A2J5tMU3UZZ4som1PzEhtZMn7
RR4NwWs6VHOnYTB1B3t3WL2xVXtF+b/Ktt4nkK81Ii9Afm6ot4e4oseDQKNXgFVs
wDC9KEG7ghY9shZ3RrkvEwFrpCanAtLZ3LhujTu/78zr2G8Rpd5h+9bziKyAK+kT
y01GySZf+pM+G6DpHBZxqAiUTTkFlE+1fIFwj5u5ER8f0hhU88fAae84AcLuoJl5
IBCDAkDI3Fdgypw9uLOld4fngtKLRy+rm5jEcRPY/fRwPt1AdVD8AhrC0WnmK6mt
sgHnbk19sicHDRfQglhotTqf3DwHqARDJnvIxJPDbUIUZ+rytHLifG2FqIZf+M1v
M4I6A35VO2nd+mB/jKO8YLQEYPE5NMaIomumOnwwJKJyNnYTakwOaoogjXu77v5N
aG9SStiJKR6y0YLpzoIyPFIj6e0/HB5O7X9QX0GwJLNtwKUkmw2X9ur2OWTXGfwI
WPKyTItRW+uoj8s+E3tVciY44bUR1He0Jcvg0nnjZ0OpPc2cf0i3moiy5fw1PQ/2
VThPazWMlSCLk2YFovL+IgZZgEGuXTrDM/c5ZW6PfA+IVlZWeaP53i/SC++ngrjU
35BkD6EQLC3zS5Nshfu5NC4HQg5uL8kT3q0YdXoCeBjt8/z0+OmzPzKHZvYq7fQO
obTLC43sZdEjanEdzklP08oZpeEw25lvXK1AwJ3ZYtkK5SwUqcgyui8IPmXAgA+d
39MtceYj4SFqaSn5D0LKCM8qDy987p7eiY0BewNi2EwZr1F3ksXWu0+65PcoV4mP
q8ChJ7tkYH21mr709VtQ0EYiEGzh9ZyBFxK7g18UUnhE5F2WFXSkAlfNNc+v8QDg
6dUeQjD8jrI2eG6JZUol6EJFaBqOPZ4Sz84+2Z0oYDNu505KxTTZRNaIO+3/sb0m
jmYcfzy0r53VU7xHzFV396xXhWdUCNCExEb003jXFHDn8gSznJoZvyvzTsS3tsQE
eOg64FUWAiIR9MEjdL7Npw7zDOB2UxTdkBTCGOGagCS7qsBHNiukRJCKxC4SgGm3
vnmbej508yxcw2scc+T71c7vZFjGrDHfsPGTV11rQQajucI4muaWBUEq5daQozP7
EAgTQF6ztjgPDWrlkatux6NkDeG66jbFseYmAS79fNc6JWpTThlAxkbQZaYdNS21
3CK1P7CiouOk5yA2tipYL2CrzWokWVF6z4Zgns0kx42feaLPdFTKXcH6+rcL+uH7
GcZ0eIdGUVwTsJVJdkbKBiYCwQLw7HoPIZ7LKbcDPNlC6kEQJLaIS9aY3Bb/I9GV
5qCC055RiRut5qgZoAHiVLo3Gar0KyH+bdp+mrf4M8fEvSMT4ZSaRmrTtNzXXYZ3
T0Dvv8sHdPhMeN05PKAac53aZ9c8Hqhx2lkQd0jbczDy8UnUrLYvVVsJFvwdWASk
C9kI7AK2EGjfs6vDALX89RLoy55+8NGUVHTVjtq0Wp9M/ILItYWAOLwu9DXj5oEo
DS780dTxBtVz4b45NP4vdEP3xw4+0Ty8bIN8ZCBmUWiT4MS+DY7+7Z4182Zzt/Lq
JJvRSeEeQnZMp0ODAb6kzjymTVPfdFks6QFwTBcJAQWkvdOw41mA5GMRr6f5bmDy
5xNymoYOuhjGfFeZOWzMxLp9XAZh6Qb9lpZSRDfrCUu7zQ+cSWNXfPZ6ggQVBvHP
0JYnqTkaeMXyWhqhkntsiIXrVZ7bpTRzE10mReWJQbdReepep2kbUdqriqmpFUyL
VEM/saIsimhpVJhLtQnTNXT/mJuGoQjurbJAMo9kof5P/GDsUzGOhfFkYT3CZ6FV
D0eGo7vybPXEts5T1bqYWXYP/CucHTG/FMyKDdlsKusLCcMMu/SIfxVoA5weuOcH
ZPYBNy5BORLa0qcIiK/H359lYdMxWU5hRLvJMpv6JYNLJ9cNnYSXvGpsttaakvJF
eOIvyEAV5mbUY/1ZjBoFmfjy1nZ3Ev09SPX4puzwIKETgGQImLKb76Xz8WCQHWKj
5Ep1o6wx2q/A9dItkiXzpLGMkk1b0B9UJcLW0gh7704k7DWWnDhlyHi6GbeKIy2O
s2+FyS/51pyJWKMnQaQvsEfiMThOQU42RQD5SbBgdOW1jNyi2mWRhfXev1reyKr1
hvGVXeYHVZNvKR9DSL46Ml3uLPiw/Te+zziwPLPHX+Via7/1sfUUmpnXYkrvrv6/
JSSbLEWEkd1c9OMVh0Ds58r/lBu8Hpldi2IsMwE9jqG7itwEdGcIpcGfPL4nG+jb
vHKqq1tb8ybOreqY7aNRoHfG4lnr5dNCAyfnTCLQ8G+sXSqp4Fe/Ypx9Vlc734J1
IfB2qEvHgz8L7k0eB+eMLtMcUNA3d3b9pvQm5y6XkvJx+1VOf9tf65hQnnThCrwT
xCM93OijB6KDhEt7Ju6kFCYo477k02/z1WS0hkkOFrF0GEpxd3STMep4rX7eQZDU
kWBOdlGM5SaQ733HQmIsPtfHFHtnpll71mp34ZTz3d4ZLx/c4lJuihcGEgU0cZer
91VclMEAYXPEx56KGD244OuGg31ECvZoyGFYPDysu6zOJ6yZXiE7MmMi9FNB4NmR
ZxCqURczhB7wUMf72lfaDn+ebZcMOKb5ziO18CWCEpxatnc0yCF+4vprOUk4w0R9
iEpHf/gV+UXo9IZAuQiak5CK7yfhN8DJ3y6txkusMewI7P2rkK8AOUsDweBthMNj
DMvo3ctKnYQ+19oxcHiBRnMO+rVcB4udqGbxNK84RJNafLXRaNLNd3GGeVDcconN
Zqv9CfB8fPPzletLwV7MWgdp3CJWDh/AY7bs6MYNqZe4gEz7vL3T+1i9R948cPa2
ej8voS7rxUA1wJjKC/o4GV3aLL9D9KFH393096FCF21NbwDp/qWSr8vGNk3bSstG
MLQx8KCYr7yl/m9K7hhqC+EAfwJ4RHJyG1fmDQW0dl+iYpRK0AssStmS5IdNZc4V
PRz9F3mgwYh8fhq7r3l6pAVRSzBLg47ZmN+hn/NsFBSuZZiVkpzm6GY1vKrB5pI8
Viuw9lRwhiy7C/GKCDyFT0Cks171OQuZ8b+kl5dsm9hUIlkmOTAQhpsHj5ZCZXjO
DF5ZIa7nMd9vyfOP97o0EKF5k6l8dh4nubY0EPHKh4dF+SIVvMEfJv0hnJnCdTFm
5zS5kfZdlWx4FwIXAcdQayfyhRDfxXaMPuqJzWRRyztKcFyi2kfYEiQrqgTcEJyg
k/IXtcg5NnwX3SzQkYp9LnbH1r4uuwR0B9xVECfHk1mKquySghoJWQLzmFOXm3Kp
4l9pyfF4ejiQ0IJsmk9Cfl6zeL/J6mJFBOSOR8tqHuxPcDmKt+lrHHPmAzOSySjr
b1v0YrGvNYRKKc/WDfsgJlhKR58+XFq8XNX7LZSh0tiAzAhxhoMB+NaJ1PSiQ8iE
/mpXNLKgPuJ01FW64NuYvPvicUnJ12Kgtr1zxzTrNcntiWoFEuqtd/kXIptEcm4V
zaj1v0Hb61Tz2bo7ZOs87g6d7Il59IetrXWQxmHwe1/0m0pczgM9O4OJpapBsZii
FUOCEWDjyKwiLzNQS5dwkwyZfxaVodkk4fJt5AIEaksF1L61kBG8l2nz8xoEPR4w
7ofsPEGsLOklkSS0tdqe9/TxV0HkXosVJUMpZBBvtZbdWsJYF/JwQOZw4zz3/Bc6
hMJCQ17DMjjUGE6cX0r/5KDNTLVuEBMmHR7EYpZ9WySGl6kYsRpiP2fAPnYaRcNh
BWrYD+VpojLx1VyqWoBuiMosfT5Hf5HAf1KACUwja6YDgCTrNy/AU8Vf6FpprbW0
iOd++nuBFnjtWPpNuyL9V2saoPdCb6xVWlTi1NXjC+Hs7gDnKh26Aa9XJHoHXCTP
X7SY2hgdRNBptgqCVQxyeE+8MNGPXIZUJYEwLp11P6+FGdcDaLaAFT+W2TvlZOuv
79K6taSBiRJvwt7lDOEwbyV2FKHE370I4MiF8gFNMfAQc845fo7A0f3W2e8tyJmr
1rP/BlVLoh5Xomh+nM9HhcVq9cdOsvaQRoPxt0XuE7m/5c5UpiuxvV88LJMntoZb
oqFuiRmmuQ7wKPfCUktSOWP8gvN7cs47aYmb6lkb0QtvpAT8hUcNZ+/Nbap7GquZ
6oYWZvAQbNJ+TyDffBVg7OuOXkA+igJGHAmkcFQ+iZ/EoHDuw/AHalUB5pZce8/e
ZCq0opHgjrmfJnyBasLCwwGk/tGNpjcSdHt2Ayxxs5GljdQJ5GOhxTgXEE2WT0IL
KYJ6641qSlUEwvbMJVMrKvupq5imHCboUj1CVCSk7cE8V18CFzceGLonJ5xg0o7W
kySQBa9gv/1Kzeo9Vl15gFwurKXsiKnHTJKWZHRthw57TFToKkmJ6u/oevS3Dnge
Xh6AGRsmsmCkHTHfjRQrMusa6BSvKYv/CKeWrG8s7cABt0dhODtUA9RrIU/CEK1H
+QzyW1R8IM0QFSQnFkMaLRUqMDbE0/pHylns+G0qvz9S/ty1krDLASsZehVeEd9z
bUXFtHy+YC4kRUdq/a2DVtgGJ1gs9y204uFwb8Ww2pYcsVqAhlcUkCPNcLIZrDND
sjcXkx9pyNESEBTIsrLVxx7tCG9fZodUi56iqATpgDM8zCWyqXy3WiUlC6K0aFSi
HJhIp1L5N7QY3yx/0chwUyv5BQLznrDqIGrHTcM8NBNCE5dL/64zcCf/pY4rYSW+
jOrnXMeHKJPFhBvfnd82JrBUrekVg78jVNdbiIK7X8pRaOhZ3Y01N8XxLVm4ddhl
lN8IxcZms8/CfNpqpcI6A7idnATvyB4Al/TJiogU1rblmKUrLBNUce35wXCdRAoM
eVifDSz6Rv6Rkte/r2pCr6kMj2yI5zalswdK0vhswSh1jJeVE7fc9WSkTiGWPPnN
6IvjgrN82utCJ6tyDtiQvHoq96RbHi00RLcFeSTuZYqjmn0GXHDfIRh6XVW/R098
1TXwBPo5qZhX3YEyjmvPdukS2W/zyzCId43dc0Yexdk+NeCNP+sphxQGnGu2+LBE
6p/7gCpZVEeVgyjiHDNyU6oNeNuteS/QP36YtYBwsQnQlyLDYcA/tBwlnXA11toP
SFKE8B8i+acgtQkRJZro8s3fKXNYlGf2PqfiBjHcgT+P2Ybo5NdqPHxLTo6YY4Hg
EmaF8EuuPrjYjIypFG4Soo9gZ+ZFeHPefyA7qNq3P0OJR5NCyVpVP4L96tcd/7KE
qhkv9+bjUEP58XiBj2ebthe84GAda8+zdkd8FiXq+uccUa2c7HHeCK/ulXQYB9hS
gKSfjz6lYOnjPb+kb2UUGE7f1OHLptfxsfk+FLSd/IbxTUn0Tn0IxkSOm9oRyQFU
HiD3qCH1NbdKnUFsG4Q29Jb0HO7Hp+Iw3/SC9kqAkcx7ybVptZMr7Jv7+LxbAVHr
fND86Cbn3jmwBZFsl91NwmjGnvqF5k6PrLPPJzEtSBXOtX6N+1wsgCLMGc1qpsU+
2vsFg+TkUlF7G4xGfrHNJPE2NZaBOeWfVxRsfLb9ZtbWzl6UxB6IVPPSgxggPlcY
FE6CZ7HXNxVPLMKXc3pEhA0f7NjdJ8y3nkpc/ev0vBGAHE5Z4X/ioVB/nhRmLeS+
aU5u01d5GlXnM2UxWdAXQUG5VHXyii0+6RdX8XZVicGI52dyVEN5Mp4aGGp9iNdA
UbyTZOTObm+jHcwV0XwlkDuIe85aCUHeXFWN0XrxpNlaGS/SS/poVAHtGRwiAF6T
rmTc1n8wx+ImWTv47LIGrBVC8EcWk510kH2fiODF8TDKJouzzwbBNEwVZvA0boI4
j6yiaJHjETn+dRN9ljAuWap2tQ6zybpJMnfg2/drWnRbBLrtAmGhyS4IxVuSGoCM
qP7uVhpBQLaFOiuZQjWffyHmweKsmz5HXUSrNoXccNouswiabDK3dE/uD5K719z/
2+aNi7r5MGZCS/2jQPlLF2PdECKzc5oC2qj3GJTuHH8xb2wxrHhoXBrMlfipE1Wb
gh9ffv5SBlN/8APiPdNIbmLemgu/Wden8X4GsTH61cGbfWSwC5Il9S/OvjYO/4NH
N5zgu9mOjSRTBRZMYbTj9/P5UaLezturdptz7abtxuIKBRo+0rhE2G687OFX43Nb
eos+LMRN1bkW+Zef/Yy9/9awha0kdH6ObrNQmRUfaNwbrHFNIwkYmh/huPP+vGRD
FMUPwzFDNd4DlRoaQcHWolqKpJn0ECz4udY2t8qRLYT/WQPG+TMTVNPZ2TYNQpU3
xBEBqY5zMwqL7L9JKafjyd1/33/YnVWOOZLC7MzuwGfAOZr60uuW7U7mQakomsxj
KnU1/iymEi/SRDr29RccaZGEnrKH74BKOY3RTQ6csA/QRvu+GGCvag3B1n2bEEMt
die/TCyXhTv5HhFrnddLlCC/AzEhShw3f+0s8tsG4vYkJP2W6brbyE86xFpSUcAo
VbE2R4pDfo08qilyxFXYR1YFhMVrpyIreedXQNKo0Ob74VLwG0QMUMsd6eBGM+gz
Q6021ai/qbQgf4m2WlV2/vUu4YnclohznKbkdp58DIR3twrD0h5lN52ZRI6r7pcK
EkSSH2QyiDwb81pajC8vs0QVPhBjef8qYOxgID8Oycyj4upayBbuCTPVoiqm900a
RzKvSRyx4We/yFK26+1SitihjM5134CvkTLxPKJwwoU=
`protect END_PROTECTED
