`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OVyfDdYsgr++XTJnF6OYZ9ObX3LmDDZHeqnLpc8w96KqvQXpU6olJXSfzixj1Bcz
jsib81GV/hpQOaz3riiDF99BdJztl/p7BycDSZzSmrJZNogoMoAxVHkRfg5b6pUc
ElNCRpM6ar6ufUKauGloTYOuNyfHpRSNJKjkp/EvH5FRiDFB5xr6rkJwmRasZR4S
lNi/cSESyP1Op6h9qklnhB96186y6vgINy0vSqJ62jAIvzx6vYK0neCJCclhw1aH
z1aDRUMhcRpf0mW43WuOT4UefrJ3IHMauOM+pX61Vm+iQC6XJdnVMK9L1mn+lmsc
sz0Ut/n+lgZCJVnWlJsdXuCUKUhwGG9+ZyT4ysMvIjOQ8A07VkCyh1EUlJyeNPEw
1f77vaDwyFQdwnscJlD9A+aQzqRF3VNqwSOlm93UwerRHegv/66sPfiDQmkRbKok
`protect END_PROTECTED
