`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4oEMF3Vhut3B+Q0ooJBQroLCCvVUgamBdGZwNEr0aF6lGLiydhdMMvxQgVdm+RYx
hhs7qtp3WR4BssGNwWURmBwACeg35rkKkrjEi0cimYQR+E3AzhLBdFGgO65Gmr0J
AAGpEyDfR92/STiAGReCedjERAEn0PFRA8sMxfaGSmBRYm8FEGb0zfsauESiFcU7
Xd6txodXHKslui48s6SS3zwmqDTFC+g/DvWatyc3BL9H/iMCPnhft4iOiM9qMKUO
pptFFP7ZHuJD0AZ5MJHWonZ65EwPxqnRWgOu3vHqD6FgU9LS6mfzN0L6W/C1N4CW
1f9HJgBMvBWp/v6yCgSkMQ==
`protect END_PROTECTED
