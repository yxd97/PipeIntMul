`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDExjHoLeObGST2sZkYmSXmLSgv8kPKzNrJ8RplXedkl8FrHcRj9MkfLXL4yo92o
3BnTkLD4c2q9AsLskaPh5vYt/PbMR1M7vRto3wkqwL+/UHrkZOy0KKgEseQ/CFIH
vBsNDNTI7GT9cipcL4ZuBw3K4Hq1olzUkDlgVRpgqThbPRUqv7WeWOiELxhe8QGw
3Gq0f6ZWLdIdPa4HA81Y3OfKQ/npwYxhl9KLeV15rQxJfjwSyNCxe98oCqE8Vyrk
OdQ1c0lTdoRqHdIlS9VNc10hsPRn8o7ug+VCCTDA0QCsKpq1cZMG2UAkjhJgBQIE
U1dofh8Wj3zcbmqCbI15wg==
`protect END_PROTECTED
