`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2w91iFoNFFQ6jVKKRgoxtjUpsG2SC0l5e6G8Uswr0HwsaxF8xwsuwwIBcSChubZa
PT1LYEEhY1iDTHB3fZ0KWHiN5Tv2QjFHI8SloZK8nWGIlq7/11cF32GdqUicXMid
tAg013j2jP2vs2NLtt/AQOJAOQKXH+X/39NMhZo8VQgzvvDgdkDG9c4TiD+FGTCJ
dYYKOZby3Ek6ie618XQcN43slrrSlwZfnT4CJLwp6pdQGndFVEiPclOT0paRPOAy
dLu5t6V4hgAGwQgiH82umq/R5OCh2cOlTVZkiU0UJ1fh1N1DqnzOpfa+QEGF8tXA
ArH5ewPemKFefH7P0lI2fDqsprkS6NLR4zF+fIzY1ZMO9OFC0/75gYwBHhg6EoIT
W0bejoTW6cWThfEyxxZK1Wg/5tYH6Z5SreEoyo8D5AViKPQ/PS4F+gQn9aQe0yp/
ZNlwCT+leyf336cPQSUZYrMgDipkZYSGS/tm5BhOdjByZ/7vxVpBdENbkHfyXqZM
7yu9aIvoVoxZrl0itbFClg==
`protect END_PROTECTED
