`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMf0OXvRCu+YAJ8qQUh6WZX36drvdjX6T8c8eNisQFVS7rnz6CFNA0GdhtB+rz1P
fdLt8dyEf4P79+0kqlpqJBgiKuPptPqs/GfKtrHDBIK/km0jNMzF8nsG3wVRFeJf
HfaPwzIVWkfb5KvqYS3A1tW+d8FM/OTsPYeyylfAGpl3h9qs+7ctPECx9/VR6/AD
fc1nwHrtLYUyl6xTNxxgo8PowpQSBqhhesg7hjIVopJN6uJXjFvc7yxHCWbjy+wj
kAmchPFYZYyGoSw2L4a8u4HLAE4H0UueyuxpoQCCKXSjwYhfV/Hoixx1e0TJ1DnR
b9VDgOsv0ly3FUJOiMZHsKbgfHCg/9xHoNCa/kCg8IlHJ3v5Q4MVjRF8w/50ZQ39
3pT9pLyVrUB6/Y9PidFJjw==
`protect END_PROTECTED
