`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ompRlpNJt9+ViqS5ayo5lkbH/f7m/S4MpkCglQfWoGKPBRCzOfk+I6wsmX0b2DE9
hhTEHZK1Zu3b78IqLM1RqJnUOYAB7piJTNkq1+wRigG/FUxmgrrY9t9kf6defiq6
PaKwrbZR4qhu57JBPcom1xvClug9yewQY+iodl/PVSqXa3lnq2JLqhnP1HCfxlnM
QoFWbn4xu1dXPoq2Rhq8wzcqJSeZJXoWNScUA6N/XTljdWEfX+RBS9GMKBHghIbB
LsOQhSX8Ph/IfbgzNsNRGx/sYDQbQRuTJnauKT4pe2nthwdKNDWMTBmZrfuMWDz/
JtDJgnzVwHlPFuKRhBdp9j0SPAgFn9y2GggDbxW8mIwsLnyl0D/AqHFzeOkU8nOd
TRTbMymmftzW2mTNBafJeIWfIxi6NbltG6e73LkiQuJF3awMAAWG6G90pq1pL4qv
1g+tO6K4B5LDB+txpUlAv9TI3mHE4hUc56GB4l8sLOhcopr0Inh7dKNo5yDKLMu/
DhgMtblrjQ1nZFmhw1nvwjc/HENwfO808hRZ3GnNunomc8RRxOp1NFvZRgyej6JO
T5JvDmg45/HZcA8FS9X8qRguotpfgrbXrLqTHYa0lviPyVJwIdowbaumcOChPEno
tuf9YWaRPa0qntE+329E+hJn5RGyQibntH6hCSZv8/JLVT//eWpTBGRF2erAQAsF
2AC/E4IboKGfCta1bAFExPTJiVMZR699xyf7EPuVOcXL3kI5/ifTYDsMVoTgyGpY
2Qvpfd4AR1rntb/3wg/FzPaHnufP8b6RoqzF0xMmPj9I25j1Fvl3ijKkn6wUMHkV
c6IKhqiG0eGElq5NUzD1GLPmSujDvrZtYRjFWLc8ZtgH7hDcPwlQXKRwr6LgkXZx
qYtQyicIv+tj3X/9j7nxdXq+K/rfpu7eH5aM+mHjviZleFmqlMzYrsav32iEuYPb
sCxYvpvCTKuJ5WZxkqjtTV7Gg99EWUPMuxfZiEzNXATQt3DlYW7UWzKbqouXrTd3
ruNj3BgZgC5fRubJiTJB+89IxJbqIa48H1ExGEUrI1FcLm3PFsqJy4KpNmHdl524
xai1rWZ1svFt4T0g4LdPIRvD2vA65bbKMI6j+Wx06R71vDoC99wpFB2nEZ4DmdNd
zMFetOgs66bcpzbGM8dfp8J+vCMCnKbMf8ZQOqzisN4=
`protect END_PROTECTED
