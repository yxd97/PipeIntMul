`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HA01rnE3uixsF/WX7RzTAy8fNoP2RYX13nPzobeQUxu4OhYEpeJV4C8PADY9SNkM
ugx+d+Lb6qfuOo6V05hM0EmzUbs+aClJp6sZ3xYtvNEJ87c1lStPi+zKCY3Is+XV
EIHKhPqMZSBH2aWH2m6wZaN4ACM+FDd+Z7sckPxSu7qXHI3yyjPhV0XKC5BVl9RR
hX0vi5uzqm4n+89ws5KWw+gyfmGn/15P5p8Ib5QZv706ya72ESwv83Ncz2LA/Uy0
pedvvFcZLZ+fDAYWdnH2+fLRpdOVuHW/hYtPV0jgcy1tjF52L1wczhkDDeVI9Qt9
CsoPUyN0uAtyy/cP6IcG/HxPXCLALdM9KCpqGmt9mSLgiT2MuvO9KwAE706XMiDL
FWYgwzMXznEWHIqjRalyvpSJ/krp0n01ZLWLOIqKvItt2q7xorRHQ3Ieb9GOPPMn
o3mQ4XOotURhUXiCO7F+pwEHB4M5GZkQhDxeRJ/LwOG6r23dVUFb8dvDhYpeyRI7
S0gAkPinDMvC7nhbwjmrqH3M31RfDq9NIeSoLB6CpxRy8OpI0JWfBLi/rbMavjnp
gUgaQ1a+wFzHEz9oiQpdUNNsFXYBF9t5ufTN/zO9t5huuH+7ZFGUTajTFmo3HlQk
6+brLgUev8KZZBV4J41vQvKgKrBUSoexToE35zJ2phezL9LOZktMroWQjX0KeC8q
w/18mNdte8oaSg2YchbuQ8V+X/YyZo7AjyKm620EKOndSbRSNyfvTYUJMkPVRcjW
QVV7AIELNsCEfTU3STtLfhL6ljOcB43Kt1WgM6bs82X/wbe4mdMv2D8eO+w/nlVR
f+PgapxY/WN+ohiSMiZRUNFbSig3vipoh8SLu6yggDnmbwQGQUAhpIX9LJCsQsad
vvZt1Hw81CAX39jDil6h0O34ByCN8SRrZqw4M0D73xpV86KxYt+GieG5mZT6bvMZ
LV6BoV5JIwJfATgFI3iNacpootGCaFctTmvAIKhGYotRAzZgYaEM6wtWiZD/73Ms
/oRFG1G6DQipwA9RvNBEv0TVnOYJar9YbMvjJUKWz8xFWaEgLp4/WSxhNQh08/++
EEi3z4jJgHEY49TIp6Dz4yCVnjIbPj8piyhfsgJVHbIzytnERbg5CLRdjZ9q3PhK
haRiPMfDp9bhtcgHWrt9K5zbrQOdh1poHvAS6DAXwZYFK16nzG1rOw1C0vf8A1uf
qGUaSAr8kcRj7J2G2ssnBsr8lFngVaxV2mEZqzXyPk8BgUX3GI1/RaOvzGJjZZPg
+30vkKS1EpD81bRcNpAikA2cVvgn9VzQR5eXmxVOJcnLIXAeuX5FQhJi6mVD2AUS
tckcrGXfmkdt5m2CBQQYEvHHyYcl9wlTETaWt5deYbTlJSncQZ6tZ35ZAZUUkbUl
owitwCINevrCcanOOySR8g53SRAzqKz3wruv3KV5NCMSf6/R8Y/fssGD2EJxTLXs
05f90BlQv57nhl3ccCAgioFsVeytoiHnZhL+XuaWolOalQ95SaYOB0BEzWutkoUk
vVhIkfmZkrjU47E3nuSLkf3lWDvY0NYT5Tb7fAR8PEbcCwHetEJHmIuS4A0K6qzv
lEuiSMGwpgnjShZ659BXKpobuIsLmwy9XSt+FgFxjdcdX5z83ghfNgdM8uqpfN4U
ZAlMV2Q5av6bPmF4cb/LA8uHYn6ANgfIrQo/ZYORfjd3o52FdkybhiHet9/Q56nf
fvqRu3BYoTNNfJkRKxZ2NKPoBUiN9BmT/wo/RArwYVgECTCCp1QuS8gu4XQ8eGJn
M+kUKJhgbQ4u6er8WV3+dnPQsCgYycgQv0dA4CnsoaH/2yvHrj0OKzZdgRD2Ukkm
pJcFR6U5EE5nL3UsHUBE4bJeBsPBkungiBBR6xU7iYavDGDLcPpITjHgrkcjdudH
1edwelVDQsdwLHtQReYAUvMKHrP/WHg2r5wySFTo3n5PR8GNHsGNTyDNjvNHsrFq
FQ5qpz7CSjQ4iPJuSU7kWz6EwnshLsnJR4GFIAQWvkg0wn8c6TlxD1msxoagb7h5
02fgwE4vO+xDsTInq6rqcg2tnUkS0EGZFZSVM2CsBBhZ2V7wGNUy3eo0JxZIg36+
pQqDthFbI7lx/LXJJOZEuB42NB13L6Gla58Bua1YsPuybEQFUfHP3D5XzRVX0k3K
F+P4ODg5qSR0K89FrneL1NwGFqscNBDZVqAb6W8SsJF9zEQD4eChUYyvJ8hWAfAB
w8UbwnsFbC132LlDLhRrwcYumjFQCHLnyicMs/w3cyWBYnjiRVGf+olueTtDZfQe
VqZXWeNv/F1mEtwYQEzfrDSE0QmA1mr1Ui5lrRS6tVKG+lGor2rrH5fVxileADSQ
cQFTTot5yL9tpc3tRYQNax6+DUjglUNuZipWjvHWXVOm6e/nkUiRVegx2PC+scEi
E8fWumDVYCg513GpHUMg0cv6U9wSwr/5Z99La6wKi5UgCWedIctnPWHtNm1rvrXW
iDL3d++iXg2SPSGhI2EGY+Tjlbt9iNj59Xu+tUqm2Hz9My+kT+TZNBEfr+am13pZ
g4kuohVj4BTXy9kXS56e03rsoHfEkRbPSF5trSu9/D94zmi3tBycwt7vpGqgD3SB
5ZoUHkvEKJDNcL3ayfrFDavjOyXRi4qtFLf5stZkDEkEDAOmcpkz+f61N0EQuIlF
Eke7aobbdV/OTRr7rt7RyVeLj1Ei6pBU8gp35qEts3m/i9jVPCVW4yaCXgiRrzzn
9VzoOuIu2IY3yUyNLiyly6a6/cjd4HWz51N9i/e0+L6/Qo9y7/+Yu1YOBQ2r54b9
X67U3/NfXdjY2w6Kd9CcDdfURm/5ddUajQhLWFqybn3PjbUgZKM8OB/2oWnIx6mQ
D5UT1uUwiD92KNw8+RGjO15oRPtw/xmsoauuH2XoWZtPYm3z0QLvRPjXbZUQMFSt
MY4g4L1hcNoYoZ8q8KZS2I95RdMdLd/H/8OwFpyRi9GlF8TNpnC1BSY/vHiBFlvU
ud5z1MHVi+liZsOZVytKzhpCCCzYfGJ5R+iVlHlrNjQ2lRXtINXMGd3EGI8/Yh62
2YCcy2fc9bcxwccaoQNT7BHrVb086E+7vKk71HbfrPoMD3sl13guMJREXolmPFtL
WWF4BXjUTvt6qoQwjup96PbRvoz+WkwUT2DV7AWZisMjLdTRRMXTxsvkhI54aICD
2pTjm9GJ69qY+YgZ6nwn0OWH2VxN55wH0GI3/WUa7vHCnBpYriqLcH8y3+WFwdFs
0+0DbAD6yh22RLva4t/CxIiFWUZTrqWpFfqvobNg0GHbW2jIKcni/+nqPVnK3LM4
4svuc/is/71K+iX3p0/ITT10gKuaeGJHsrMutcqL2eIN/YP+N2LBOocGuilsMrNy
O2aFWJEGz1TeutTtLXVo1G7Vlj36Gdheu0IGoSIrB800pEPa7FVPeMENrn1SWiMV
sOimAIlc8vHOO9LRXWg3Zcp8+5HF6ZFrJ79LLU8jU3zUnRnkWj+kHbP7lmSklDhf
5WZ3ii2i+PIcoEVNae5XyHW/0pMdqK/HxiFsEzbZMXqZj9j79nM/hZoTfqnZgbbq
HMM5rk5pmMuqTD4xyacaStx5qsER2g/J4fErG7Lt9aAfBBCHyOgk3UG5H0OmP+/P
v23VCvcdT0dSCAbVhSr/C6mtuvTblO35BbsrWUQqU5T2eZyjAdsw2VvnSAmac+QM
15JBfF/BuvMhPgT56TRrgBrCybj4YCoNYfo+aWHd2yOkZBmJeYttk3dMvQrU7GDd
RRhdV9qE2ijCmfgXR1TxaL24Z3X2iWfJECqJx20rVogIWnaIaD81OUNpvI7b9Y/B
dgEX3uEk8ohcIbjjneJgvjAyXi92NH6xKC+sm4IgoWmq/Xm1MxDVUJXtlg4s3pbl
f5oFMgY2MxwrNpeI+XAIHeaEMn00Fbt2yMXRi0q5puz/x2LPl0IbSPJy+GS+xqHl
tU94XD/f0X29oItJJncBsT5MsjVN8ENvLu+dMSqAR2PO47PidfTBp8SyO/nmOa73
iKxjZux4lS8+ISTVjPpXUvxJitnxpML0SYcZbFpR0iE9rbvw2XaGKrXUo7sSKpba
WBXd8nsL7VwRzRBVWtHKIaBz7kQEO2mt3tJUoYyJ9Ksse+NBJifnR3BlRogBF4/l
faMB5DqojzzdQ2BiVsSgnv9x1wqmwHc/4uWy1X7q5H1y/3qgM9Z8gdQPIZDBF7Eb
SNM4I4iHU7worFtXsx4W/zJaTR7ZezSQZkcaheTBlOjg+pDXau7qCPqlevhAvk7Q
y4HOHjIcnej0eOjXrWnBLVinsRjCXsHN+icm/13WJsq9UMLrUORDneAACJeY29oC
e1yjGg+23WrXhmUCqvPFzGISGhw6/+BV1vhox6ShZhYOj4sYQ/hGI0Y6A+AYurTA
vPbGSjH7nWgoS+CHqCSf+4qeSZLM+0/g1jXxE5N20UXzEHqN34E4yXmZ6UKBu+mn
+bG9GwGh9zOGCOCtU8NoihBF4HqKOfnnt8H/bIK9K9Q=
`protect END_PROTECTED
