`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VNgDM3S9qJom5Ce3EGhcrvlPnk0TgshpO5sk6bUavxWuKisNCIvA/gRa6qVdvQFV
bSnSVvyXcK3DHpHEBf+WdQHKECKh13JQiIRo0Yp7w80lBnPWTRj0EOlntCntZ1IF
SPqHm6UoCDBxVnRZXp5lbLCzFIlVsFNaQdo/iGj3L29/+gbsKCqIbGfR49u38H4m
xCN++IYEmzTJENrTRQs5rONngK2h9pctYT1QMzyPUQekUKSayHzAWeopOX0wFaFn
zVt1sGoRORkeqEPo/nM5dd/5IWGRZwlpLwf2m0nb8XaG+N1AFUNpOtps6XdyKCFE
yNCd+QX7Qyqk71HIGGyzMd8ZvOfH26gdZ/9GXzzCD00hHxRRvLz5ZZXgQfoNW1MX
RcQJZSTTwK8UG4KDLQzaL6VJGm/jyifQDfpZpYkN7qG+vlpBWh4TL40bTlJALHdl
`protect END_PROTECTED
