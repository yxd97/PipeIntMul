`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RSRORQWUqtTCYEHlJxkhwshTbSS1ho4LZr+Ay5NMZiUY6wg7bubrTsiDR/Gulx03
uzz2cR1rDVnMyT535zdkOY4hxVDBY72YMGNw6/bfUfMD/rOGzboBi1GzK2PE2iQ5
FbzeUF1pMsSlXGkY7TCxbDea+Lc/zNXFjNfV4X5b6eYisM4+c1YOO1dOVZqpqiT8
aX0hhhSDSoQecvygippRqUq10E1L9Ok3+p2/hMx9oNK+dRnp0b/V8jeXBpTSDX91
PtLtmxNUzR+qJRdSpkTWuOCXd8HHF3yEnuURgWszyPFDxyJACDdsZyYHsolhF0rY
U60zo5s4DS0GjnVMEwXWpQ==
`protect END_PROTECTED
