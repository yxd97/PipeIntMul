`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nSBjwFS3G/ByTm0g18xAqMtcxeZW1aTtjEUguuiuZPl65BBf/upnT65gPT8ffd2v
Xq3RRbSm+wD73WggwtPwQehadJKFTUFcqDoc4oKcpvDCmOctJ9KM9f0Ateg3X+cg
QdvYjE+d3UMCXfN6mRJX1FSUvOKNzKYF0R7rfaxpFSzvdXm9ahkksy3D0r53jAd2
IsmMpW8LP3eNj7+eMSFsiOTQfvT0luYIvr68PXD/FPH8DNBnbWrwzKXESNiMmRMe
ZDPnXQElAPELC8X6xBKm+6N7kRKXJ4qR9g4/CUtZDyiVOd9YzPqSmZHwF/KGFzOR
`protect END_PROTECTED
