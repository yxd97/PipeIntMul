`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
siI5fcvogq4no7dSzQDLx8gkuaiwzjHmmoQ86DN2lt7UIW7Wpg9wWW9H4otGb5b2
SHrOIHX9FpxtDBpSEmIF97QDcN75RCrMC2NMkpzTVyXPaqPqihaGwna4b3q/lVMY
1E2/e9EpqQsCEu6+sJ31tlUgqrGDKSEvZLhFIelB5afa/hzVOx/+KRL8u07OfIBu
mjHzIhz0644CvJLMMZ1bGfl5UNoDh5o6o1njQaOtpbEpMz6WRyhoofzE87fmLLmx
P1QdMYyTxw8I3yPgkKLWWPQxUbwalyX4Mu9S1DcmPIJUMNrmev9OyUS88KHoykD7
q+euVIhyHUZw0lnuVO0VY542qz5IdwEYIr8Cz6BmEtDa15YjGkHImAZSQM4qJJux
OMj7LmWrI988b71wmaR70Sn3Ms4EP2KmA7KW0O9xlUx8JQ2bNnLszm6XbfnJFMpj
0MQkS01Bd8+D6U1BhVUjI76mBoBXko3BHhcskBbgwplj5SntGZvgDSX/29owkd1s
`protect END_PROTECTED
