`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hu2VwAQxtaNi8gQkdUTCUG+OYYCpg31fg5FCfBmfOFQeCYFoIKC6g1EWoIwu9Lhq
zzMwuruu4iyw9cPAaSwRrUhJkk6pnKjpdQCkez+OETUT0J4Gkay3qJS9V3uVHPKC
yEe+ixC/vHGLFH1kIGYnTQlz4P2HaVtsMpg7iS17+EQDVB4LSrhdU91MX/XcpcLb
lg/1yDY8J/gxpat+LYSm42dtF3UYjpgiugQRcGK/p/V4PFnNpSsyF7b7y+X+0+qo
mIBIcXIpdsvBPlCSVJ/OlRb2I1s3NurVNtEi6tt9wClLChPS2BvKBRVvD5VH87DY
F3j9pLGCCTGHZBD6ioeQNVgA565elN2kyCgEHsXhnOzcapX/LXeBWwWUJVLMJIfH
rdWKjbYmpsSZ+t2MdNQmDGSn+uBVMgn5CkvyXX3/qUzJmzai1sIDJjwDjY3UW6k5
gBohQkv6nWsqhJxH7ypCyUEGimhFDpHZPx34ga4GfDSuJNypOBdKHIVV16caffDY
CqWr5sgUkR1JVgFcGUZil5f1QPhcpLgRzJTU9r0DZOPWBg9SNMZ9arUmcsRRqQwh
QkiXbagYUidIpkxxqDWNXCVJPfuiAZXl+ALUEmi0SPxWvxRb6rpB5TBNKY9CQsBe
XjAxJdXayCQBHGcb3WVY0uNzait4rCp6hh4jBW+iQKkf03rvUsRPy6HmvU8DLLpm
3QQqQGOGdLNxw5h4MRobi6jCLkUe6/RnFV1B9gld243OBNYQdjndM4RwOdBCTEZa
jQnfYanCNGumpy62qjaxxCDsHQs3ueaewQCBNVE/km/y9uZl/DhQXtkVxzP6/uwG
2y1JqArvUosvuhVEMpeP4gdpnNiEJeFFsE5+/tOqgfiw0hnEGjdGp7jbW2Kxo7Fs
H614n/kGunLecyHTikTDUxKIXMF3tVtX6wBcVk85UOzjvkh/d3JPCBq5/NaS9Bc0
Wd3hH7KQDVwjHYiCVZCyK0y26yJbMbc7yKJilaJJVSlnwWhDzcKeX414gXohLGHP
cN1DYhe7Y/skxEvR0Yd5rrGzkObWl83xyrL+WzlACGNoMu1I7rHvXaL4wfI1+ixo
3rBoeSxMwtd+BzgW0AmejGSqbHA1oJaDRL9uq0oSTDWkJa3X3eh4rvZCO5fbnwSx
jkKYhpGintWiyZeHTKgc3A2PeboAPC8PE+q4tFH1QhCfPJ5WJJNiBb5nGQhJDizs
77aiIlHxxG1Pw56Oc/2HY0HtZJztuEevuvnnYtTfOXI3N3JxTL2p+E2aCHTs84Xb
wtWYtoITJhPUz5ixODWPLd6BrMvPcaR+ssrqETrVJNYzZGR4UVzLuAYBehjGCsBc
BV2r47juEA6Fzu7zA88lqAZzBqB0jb9XsdE2Nevya2yv1A+v8B835d4m0Zzqjz0k
TFh9kMM6Sc9lwiu2i4ixR/Q+v6JaVBl1H76xc7wSdjJVFzCvYF4G1mI+quyTGEDL
OG1ChXxyR7cWZSzc2m8Trvv/ZmZlhf0moNLibxA2vPZLlR9rJZtVTrN74ggfo/AP
IcUC0qqIpCamhOkbf+XgUPVyTCal/iRUbB5tIksiYJqAFNHTmxSYKu209/PtSykA
jCK82KHcGAxCPke1Mnhong6MacvmjMhJQI0HLL4Jgwp9Kk4Muc2HR/zFASkanISG
xoxEb2wCrgpv9hPlDX75cswEKl4owOl5YpVSLqAggikgWklgg0WrDewkzHWKHW87
6FxcvjsJrzk5vJ1x9EbTSmu9483Z+YTVQe7faNnZdh4vJIEGsr+BdlDvtF+h0X0R
l0SYFdZ0nT9fberWkqbc1ijKzIoUnfAtlaprIxNVqcnEKclCvfrkF4PgB9vY0MST
th4X/U3sk2VJsc9sPUkCEqErv0XB358+BvG2gzM1felrwSCyHSAP/mtmJ2NTuPfa
v6xTu65dI8YvQGWESMHcRS9F+E9FqQUb8l97sLvM+EHltb788xUAlVLcEeWr9eg/
nx/lzYnmGHlEkk++6u8gvDwD+rNMQp4ourI5uwqBlDkyifWoQ2fxf+vCvVqECp0j
B8ecLaz8u4b7xTjIiTq0kEf3DbisASISLTkFooSLnoLrLsbCHh5kICxSPo1MXBZj
iA9U9zPr7AAO3F+wScouq0OoKIzZIrFHyVrV8tCGn5qSfPFj6tnD7Zxj5eMXmJSf
f//EGkTBgWc6FYwulTKsiBy7ZXrgRN7RRiCGddMiiWrOPbCTv9McR593eAKBkalR
paGQY5i6XC40K+IRdmiZXU/dNEOgR8whuYvt4u3wvBeSF0fPH7CRx01h5ZDh+d58
a9OjZPuE1+AcB1P7K2BgKUybVSDOdpPe7RrJXd7XrOM=
`protect END_PROTECTED
