`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IAUo2630JNPfMy8WQi/B0ohJmvu6er8dJDC2yauQDUEVL8tMcjSpu37hpOmsSnZo
QzyJbnLSjLmvH1XcLuFbIP1ykogiuhj6an6SdPUYIXCLPCe+doaid4TaPf81hQ8N
ffbKNm2nD5GmN7RBrAP7u5hkVZefIMaUwpxZU+6xykb/lD6k96fdO2HHKJ4QJg2O
ZdEvFY2igS7VqP5/Izw+9jHu6jNvv00ZZajAirAOjCCty2Who7PS0zYV7+Z5zXh0
rynHnysIVGPwS5HDpQzCfwB4YVGN1hOcal0dUD7AYzBPZoLhOBHRh79KFFxBYVKX
5D7NocgtYVT+YVz1kaI5uPbMpMqs/UYCtF3B34+gpHlAa+OIznES2b0tXShcmFjj
`protect END_PROTECTED
