`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0rz5CK06VFsRVTnunBA/qP/ICvoFONYiLEsHzTs5tJS7IPEMDF9v6/Ki9X1LcBW
BXc05kdloYSPzKDPT51bMHi/ytO2I4IC+sNULnHyxwDkL2dmgA6oek/JUuQ/ctX7
2RrNO0ohJ9KblL9Bt4hcgJsDOl+xv4jWSaZVKZ0wGccWdHDprDm8KpcrjU9jKc3f
nlPAKR7SxJVq6orZl8f85BajKezg5plGxwS6a2VUpOeZZLtGCESpthUu/WRtb+PB
ECmzIVxsIpc5t+6Loa6bKtY17m7h+mErM2F44ci96gURFKCNuA5KNrsdylTMdHN0
G6gO/XsB566Y8of6V8clob1BY8nL7fZqXVgtXE8G+AkL3oPS8mipkAOXay2JLnMC
W5rGgwreY4jbf4xxHBDpIIyZrfrSKgbGOoD4djRKXkZphWPlLkIDy+YzT72i+j1Z
tQKpvHqHULiGtgvtlvB3TuxeeZK4ApADkbvHIT6ZKIxaV0vx3TejLJevZkDbUEEY
4GYPQqgPSh01izdCvsWDdg3bYgCciRH6zE94hbnpmmIfsSG40bz67vNsEp0WAiqY
vjGQqKY/oE59q2yRm7exndhO0xrXQXUXinpjyJjpwvuhMerOIZYbIbN9A1OL8olQ
ru2hcIuoBYwCqqUaCobPkf8fW+V0WI96gv0EpoejgeY=
`protect END_PROTECTED
