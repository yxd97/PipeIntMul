`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5ei4Y3Oq8XVFiTyu9wfDDLtSG1IoMBnrMj10BQyMs6GDeydxCkz8rSk1O2neQq2
/INnUl6fQuyFwx+PtOBydGGzi2dR6DzI1hqpzP1jh9KfdoN6bRPQxpOOCFLFbghc
3qloo8dayc4TYVHH8+Wu+bOxRcA5h4DzrSpIOXqFk0kN6GUs8QQsplpO98RKm16x
Zj1L+enjP6GIkeyZbieF4hXJkI2DQCo3MRTjEbgdqaMG6Yk2lAKQHOUdT3vVQjkI
VuETd2XQSiyNVVSA73pHf1+mItDczpPpPkSoumTBM7Rqi94SZrb9EFqYPJbpU0Op
CceHzuDYQ4FpTbUE9j8dSWKxVVQf0QW6NVB02mwQfuAtG2skKiwBgEwzkjVlQ+nG
TfLr2yfCPuiCnPoV2T4fXbkp4OZf0C/K8OLApqUYuNlD7tbQFqcTVAb2vJVyruxu
PIQvvcdcwhhIUwkPVjO6itpFT9tEzxLI733iEH/hFC+bZ/AsW+jv3XI6SRJNbjCi
TQciz/wNAlkNSchhhsiNrWr/ZDuBxS+q+kUiV1CqAL7svPgeg27VGYv11Kc/yIF+
`protect END_PROTECTED
