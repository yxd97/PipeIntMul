`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxaIX2ZPz2PtJ/GtiVqjh9S+GkdO1bq/N90z8lQQDZNxytYwNtHhr9TxLh5ESoUi
hjP8sc4APp/pGh0tFM34/ADfEHSkgOE4IyJMQlRf1XiGcguYdCsRf+M95254E0me
6qhi399I+d21gsJZl7ndBR2DFvApwX9cWS1KJan1hSYmnEfYcpET5JqX+YqT8Rep
WvLwIkXH/h0VXHbk581ZDg+BbMdMJqkJj8LhELHHDoNU0hFGwENCyqcQ4ByWvC0j
6/sD4Ka3o53tGEVqXbwtx7hlCZCASIJKg+PcGXZCsdyDp9jr0pm1cIw8KR2o8qSr
VYCAZz0KlKXpQql+v8G4JxVcT79JHVMQQCwAdyR6cCBhWEbkhFniauzArP0Wgxju
DaPuTLwZtDAvgJ1xdZvh6fTi4omTKNxi1B4X17D7V5fjKoKIYyrPpnUIktswaNyl
`protect END_PROTECTED
