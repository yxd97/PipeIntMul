`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IgT6Ek0rOzt2RIEaHaX8NF/3kMG1xrQe+e0ioD5QirGPfhbIE4uFDJ5WLYqoHv47
Lz1wUVIOkeYPB4a8O0Sme3Rf6y6vxH2OqPQMJ2Wg5O+y9pqBI3RFj4gYQcJyJu+K
a7hr5p1gC+MvOGwnnuSKqZZtn+FH+I60pGaCULoJpCK7VduVZS36Cb+PBjhqGr7T
U2LcipYwcfCKbCCnkkB0J+JVnK4yfiVqOtFOnFwXJlcvailP1gJkhH74Y7drhISL
SHE5I6tbfwG/Fk4SRSOSOr3905hqeXk6sOfAjss+IS07a/OjbFlzz1wR0JLPeo9d
cKaoH4TIeiugipLt3SrSFFOrfjOUpxJDtXShcm8LO6dLW6hmhR8q/YXWFVaLQQlk
FCKU0Kg5tcNVC53DrServCVKtGiZcGnK8S+i3CutRjgZ3Xfy1viSNYnhGgSZWsbp
vI9AteCibFxXn2eSk+GsUcIPEHqOJjdYkRqw8dvH/zXulp8YqCp7Gy4sCneveeuw
JNCQ/BL8itxGNM6HjwUvRfi+122ArLiPWBCr1QXJFtckbwNY5h/MzC2FG64iiOQO
u/Ct9cYTmdvIZKBTdRr0T7JPnZF/WsIWDjZnTaY7PI6PONnnIZ8h101BiIfWJThJ
/ORFNTqJ422tpNUuI1/wsfLTVPFPKIkx/xqUAW7g34NYv4ZRgc3XB0T5C29bHG1C
7/euArD3IMv+QTtW6ihfN/tD2jutKCjkarufwZiARwPGJtQqvi0/Lh2zTErdlUDy
3Cl8FzQwM757c8Pyp2jcuEiksuKhWYSi1kzX2tyN9qC7lsYO2TzuQJBDy7+aS15C
p+NvvVYi5G9fkna+g7qqfDpPXpbL7uMkjbeH6WQ69gcaLiUxrlLxzNArzxez4kLg
0zPfn2o2YFHjPzcfYOawhoNhCKszv8LSRnf8GQvaTTdKlsrMW5wAlknfXYeOW/Ub
ozA+b+J8F/1Het8d4XqK/JYgjse4z1104xjyNN50iZPLWrHqwgDVQHSRIORcT29/
bGWV4UG1KinPh58jLNgO00PlYJErBPgXJhtV/t6JaUpCJ6aGJvvZTdTJGb/wVd8a
ZYd0scNcIKdBuCUUHCM3eCgdXDJN/rdZPvsAN5m27CNIMo97Dg5/hMhDPyYTCpcA
Bw//gy/ALKahx1lgXnpVxI1aNt3NVjr+n2FWVKIzGntv89tUOaX5Mt4sXBROIem3
csxoSE8ZRWJpoPxaEcqY/KW+uMezg8fSpzm3DY5G84wBD2Qj8hXERYn1gYmpRmHB
qf0BHbDGNlG/0fVMDgXuiLHjg2f8Ihp/3sif0kt25rYetYvEM08o+SkUAqKnGeTF
ABvz1FiT5/OxqtMlI+bky6PQ0PfFn/1S0NhRnQuZQNKxbsQ4RVpaW0H3UjLRO0NL
pckTP4NyTIAXRbniUSpuJ8fBUYII73GsCPb9SKTB9N2KiOiNX40ZSDJFdHtYuPwW
SABjyPkcYoeS77bPCFD9P7M5VFmkxmxyn6dA10GkOtZL6e/buk6YR/+HnZjq2OPY
xxE7jSA73933m12k1ufXZz3w8YkNZWUjfTEp7bV7ebMKCeHOZAXkZUZIEARMMc8i
oljO3ZoUGVsMQkjqgPDhdf8yQr3ilGkwus7C6mymhWI6bOaQ5HlIMS3Opw2WIeDu
ERAwFZZ10YPiSWK7sKrC8EQDHsKcVCCz8bUZJn8jy385FzYXhOPvmE0DtYXW53Ke
B3bdZf9tyRyhUSc1oMMv5uwF6DDcfiIB7/9vpqwZEIDj9rXdTU9dvhTmZZotJIr8
YXkq3ijVnWW5cBgQzP+hBHvEKkNyxI4FUlXj7C/XxwAzRLd8rVCfpPiQOtI5+9fK
MIubPKVe3q+LyINroCA+Y+86UhDMc2d4QSTTVdLxT9H4VCHw7i2XbmFTqN3xRqIo
4wVvjl5qX6Ms+jhHSr7+mB09IIub6aHkA9tVWEYEguH3QWJI1vzySLzd9iPS7SUc
EjU9oUgFkVR+HEhDd9d2kVmNR1YybZsfHfq4D2oX4QCDo72ze15CUMBhrd8zKqt6
9OFNnjIiA3kWd/6jVxL97R2r6Nrtr2R6GiYf2zO1K+5TgDVmRIjLB6iDrzQkYVmP
TFC9bSkqGpclXoGDYdoPGUmZLBW2JoynONo3utdZliJ2KAlE362wwT9/xqu/U3sa
3Mu0yOvmsbOgDqwAX9Y+tSoW+5uMmpzekl+lcQt2PuoZCQg8HHw42jLRTPDmWu3Z
C5EL+5ogVztthlxqdy9GzO6uZkdazsk8SPsfHaYsGPLkAQQyiT2ipCgn5c8qIkKA
RRAfDfQu1sdDqVzpewXL2T+3DGoYgLDLLRTMhGfOF1A5fV2tlhj5/yrllTr4hLPV
/ifFuvHPMkII75LVGCqnRLQxYfayWa+W+q5QPq7MPdBFVdn9qoLrbpzbD+2NqvdU
MdlxfRlENtZ/9YNJmaHxWmEI2T4kph9bnjZTC5dmygOzsU8Z0i+cLYXAdi5aXtOc
k7ALXzEre0SAprbjD6Xz6Cddn11uCo5XSc8oQFKJcyUAbd9oyvTY+Pr0rW/Vf9mG
3/4gbzSm92eaLMVWDO2El6Mu/+juFTQx+SA3z3OFdQJzTEWr/DaMspccrjTCAxJh
ehyjBLLQFhAVG9+RUuD21UFkgk7gsxUz73ZQ8yWOxOW0KPig3/oyFSrXi5/vESZJ
ysEVHhbpinuJZ4DYfsqzdl4ozlHpDHJ7PLydlFFiyOm6KNIIWJPpc3kFUs9i4SfC
dKp8iIXJ79rMzX5SgwquF9gSMh1ZcklLl1Aff2+Vcy02PtoFkNHc7gOWBmDnH8q7
396fEeRGGXPcxaHeK/Jq1oqd4n4iAMQH52MSTfjaF6qhsfsUUVhHuGyBldGoKbwB
TtlmBVZDcIKys9ATIvhzCQ8OhilwVbU7n5iFElReiOyzupAYsHd8Wk3pNkexZJZp
BSeJgTlSmKS5h2hhOeMQ866z5LoDDFutPtR3znAt//A5LWV2JFfbWUfZQkHQ9nzm
+Q/av+ApmMlGVJ8k4BWYEvDuBsbKXrZOSX8/IcrwiDlz+ldDkayJRF8K8jcerKyA
T9iOel7HFPOC8rnhqLgBxDNjEZLOJAkpjmHri6UR/ClhYFVAeuTRf/CLZklv7Qxw
Wt/XnGaUbCugJ8neMkNEyxUzMz80AWsaASMdZv7mkXqG8mSu+jMiM27VDmxVLNyB
QFjLeu7N34UlfT2sjYQQi7gOgn888+QN6aCJJC8OCqcvF+mfj/CeoYirGyT5zTdV
yEKOuSWiRRlnUdaweWaRJJl0qIJlBcjHPwiEoUq9TcHFCdgEjZGD+qKDdKS2FjF7
slFu0DACRY5qWITsAVcuGYLsZmNdH3E04TYNXTiAWnyHIGh9OJia5Z4EsoMrW2c4
auFbOy5w5nkD4eQKNR13PELQGWssn2y6EVGcVrjhnWyPKOIV2KXUdjGU8tfc43TL
8m+AiT/BLmE5QgOwtcqgcfbfgk+pHvuU0Bm1eRC/tTYzUEKQpfWTRscCoCWA2aEQ
fuA6loH5STGcsKHzgqIqG9SpEFhiuRlNOWVKjC8LdHnpGMnBdBP43MSsDzA9nHoe
c/XahlKuWff9OtFEaQrWliTk9ptRBOY7IO6YXUIvQIfFzJv7hckTe+gamNCgqKpm
vrSHtVLsQ17PowsMlS2DZkGZJ31sUf37inxKr/J9tLRWgnLSzSYKF6aXxU1P/k0s
JPagso/yuX6bNZwxu5OebHsxfOzq8JaByAFdh8fxFS39WBesKiBKmeHNWulVUd+Y
g3vhhcnn64jB4Z/ssYmY/cZQJBVP8kqoG+YP3T6Lr4cdJ3ZrzbM1kmYttLzEVfvw
k+B3BVg+hV/bacP0Z9iPBAavfsIKcAb73Pvf18EMnXcBhrVte+OFucMGs85vglsS
XrnulZ+pdRmnMtTEu/cEcSUtjmrq/NYsaTHV9wLRnKSHI2UydvJzOCGDk4uvisAB
BKPOesFeuzmQWABn9NzEO0zdtGQt+STNcuoTOoMFY0P5szUsIbqigcu5d7ufCmz+
ustGPe3GuV0m3ndgSd+doE7PDiHZHzXyeBveUyVKB/Bnt5DIeutUem7D+euOqLCf
nWG7UBrZnQX03Kqp36qkahQvqv1bPTxJGI4Ymh9YIhmCMuEG/l356Ctqt0duTG8l
PZwVo+0JazpN5X21hZSxWvG5z5f9sXcPh6N7WF5w56rXUYh512zdbCsf8eI4LCFS
jeGFevxvHnBy+GpvfE/AS0wBk6BJoKXuvoXnS4vGe6kemRtiNZg1yeAUlpNocQnN
N04vuem9njLokOfLEGDjK9AyuPBUlImkSBVj/uIo1stOnfvGPf4QkD9DwlLw7sq5
D/g3tn8pReGAozwnuvW2Bn6erFcoKzV215TR1wbeF/zWbGuLOqWQqxuPUHUnzKQJ
BuIDwNyo+iS5GUnawsaDSE/FnzsJqK8wmjEuk+QWdhN1k21USYVl810aGRwxv2ze
dITpadu4ElzyGZlErbz8OGR17gbVm1x/hZTBfRHOavPxts3Yy6zj8lQg6K6cogSg
NgKra7cFXtjl+j7WvlMjRIe7PwTb56U3l6zFFq8/Ye/Q7hbcD0zTo+XDNDzxiP45
QJtYZCfqeEm7tqyJxb04xPlBwHbjNm2twxuOGKvOmV0RU2z/H1m1VfR1eaV/Z/9W
cl6g277lpdQdOxx3tM1kR3F4tkcJL3OIpOuxo0uq4loaRM3XcIdJskjSI1ef+pf+
HQuZcwcwDX1Obmte2Kuwak4ZSGszskLvP3PILRcw148wb07t9gb3Ii+xEoA/sOJt
1AVBr0YrOoQZOchztNi2+mIa1eiFPCfCGH+sePglUB7DMvlDCJNzhz2iszQv7f4d
dmx8Q9wF1wi5DsHaE7EMi52C3lNVOZT58gZ86oB3yaRCrVx6mRwTtiK6ssc6o7Vt
+NOkzSfCH87MY2nMRCy0i2P7QKzhE9BgoRV4XKcXy71KXexFuqUCbJ8bSOweSqzo
ANgAEX9i7w6BLKH9P9oRke/Y0bSygfDKlRLfMykVIZZWOTTzFmo36MJ6nwedW9zh
23wpdEU4Kj6DVPl0+IdaUpLEmtO877U6IfF1t2gnFM4XVoVar6MnrNbDdZLUMjwA
NGIfdk0Mnup1NX73OB/6K/5yY16RcIiY6QpX/kZLxCz6+9DvOAHjaXag0ohzocCD
A4xgplZp/1OC1vtFrNK6FwVTEU3+h15vk2UGNteQ9bYp8PnPqk61ZORDxVrOxG+9
dUvVOI5Jhhj+7TaOaTokhCudJW0aNHI3TMMSROF+ERkSyV5tgdJTgwKr5cBMW6nY
1vIXf42YyU4pTsS7ppl86oseG3rim+Yr7DIsg9MPlvbbzzyQJhGy7ER/Jdqc/RmA
Su34awfsWdnSpnt4aq2wDyTVXsMapyHsZYv8Hl/C1HXLWszQql/a32yXuhjhs/rM
iMAb82a5w3uJVnZmWbFOfjZzYSlBF4b/Gr0uPfaEqiotHWGEtNHJI+JqAK0y4ceA
V3quGRD1yCnE91Uzogn58eMfYwWRYMFMLdK+MMdWGZnCw1H/oQu7gHpEZJTteF/L
RrPq97q+48SSFtDIBnh2sxuva/6cVImeeI609psd5P81/6t5zEaYXZgqBXLIUNDX
bV8fURA8ZtMOfYgbt8yWSXoxIZgRMfbhSy1Z6Fil3Kng+YybAnL4wVnhlKLPfF89
LSdWFSNaSDoe81aGWlZT1RgjE1U3yJeWck4PKe9rTPI94P87LswRY9hvxrGv9ZnV
cRyj2MWuLp36yDO2+nHw/Me1SmxE87eMMHZ+YsR+CsXg0A+UVjLlI4+Zp6bx1a+V
Phk4QFjiLwGHpmh52fdz4b0ymE6A521C5X+7z4SWP+rh0x49hARo84gtKrdfR8Er
sNuIJaPpZdVc0w3gfbzjDqW7PIbUxZRxfoT/AZQaxSgtwch3TrpntbtBdkwf7oHm
09x1idA7R/drcJsWxmsEYueCAc45/G+vhGUjkEtRv9QxD+1wDRs5bp9k3kHxRbuY
e9rXnVBE0630ajcCIil9AY5RCpJjALIjRcgHs1CpRbFamP7RELgZbJbAa/+aGQDE
uhWtZHYdAa72OjXS+c7o2DTGkzl59wlZKD4j8aBbihoKURPTr1rDSfw/gaCSp7Px
sNbMZr1N2itXQZPMsGQDWBtJxGual5LpOufVI1zHXNPEKbT3lJ6Zat42rGxEIJx/
CBKwcI1nTOX0TuOwK5vbq8wIZSxsRQdkb1U1B1+7ne0tDLIEscIiAtamU6txQ2bv
OvSEEwhwKGokecknNqJTmBZhOc4EIXLmlJuktZS4v6PyCzJGkIc1F9iJFuLvszJU
jhIIOc7Rj6+7HGM4pgPjflZ0tUdFGp29NbdHyiQdiEvaR51Wv4m5h5cn8s5x8M6s
mqe7PQ31XEu4hjUm8W1jlxL8xs0m79Q6x2y3uTpWlxGV5zDPcP4VkGCeXYu/o8ds
2NXold1+PNtBsM0YuiPXI0Uplp+Sx5FG9xlhGZdv9rO7sKijwvqY4Ddi2Cs3xzSk
QMfHVUBQeYnbpeozPf3eQQGH2ODd/FzjYfB9pmXL8Ka1HI85H5nbvyk4LOHM2QpN
SgVOvBXm4GV9AepPxiIlCnlttpISx6cwAASjsY9lQtiM0thPQqnKzfZuWk7R/K0Y
8hFJ88l3gxzK3oYQ9xczR8JBEQF2rpp/+WLTw+HrrWB/tignM0zPO2vgcehiHC32
/Nkoz/saYUs56r7u+GG0KFr6zLqNTG4si26mF8vxHjBdGsrPwyIKSvARbJA8DlWM
Cw4RSIJ/d7qH+3F4uSEIxL3pdNyU/WKrWQCTC6EiVntXP5bWO3kiHHMklf4m0MvS
YJ+dK+MZoiIITlJEfIz7pgMb8bnHo2CvKr5Z4rEltfDtDgKsJ5aD+8Mj6qMoy7iZ
atYBRsnihkz1d2R7RRKYBBWIKLXY2gw5ansQihd5OZxUlqCxlAkoVij1laYlxZ/7
5bbJI99VWbjVCCBXN/e4HpgXK5PbC2mUu9Nqsl3OHPcdWLGBGI4Yzcly5ukULxB1
8iubCbtbB95e8qthtyL3n5cJ64bvVbiyhvx7eYbvipBwM7Ei4aoqYP84rWnWtbF+
Mq+810Kj+cRjenuPF4vEGehb96BL5Nw+1PqaKMnnzXdnnLnSVMBwByGiRVI4FRC8
i2Q+eszxMuo5PsRq0VP/VJmAk7ta+YeP+iHQxi5vgR8tUOGU7D1u4gSpS2FPw87G
F9k+zR+9lzJI0+j021THjeYBykrjgf91x5l8dngA7XtSdbCQ8XkGaXmRWABgVeL2
uIaelgXwK2tySeX4lgPpbgH7f1Dkz4JlhI6Xu87ub9OXUZslwxehbbH6m9ij9ww+
n3VWALtHVi8Ul19WOz+z7diZMoazsoqPPPjcp1lWpjVzX0/UHGRTCFVfRFuWmdzT
+IK7JTewyy/EtCuWLeI5lroce0JrIbdCHWVY1fcZrsGWbXTy1QoGi0ZOE1opBFyS
WYeA9/3UkSKzvLR+uUEWHSJWaRjst0x8xwElb9N/0n087nhdf1UzB96Lmjpu9MNA
MchdGo7TUS529pkh2Dciy+gf0xYP5TVW9yQCq1u/DtP7uQs/Y4KdApu8+FD/bf40
gUm3RjJjH5lN5jBFzFbs4f/rWKFTBXOyChIZNcuj2vfgGaY6WLZ+DwFKqNEanZwt
pLwlI2vShO5nqEF1/1zaM5RNUslLLQrNa3xNSzex39kgsqpGcUC9ZbRi7KwTPuH2
2C++aTBWyBsXhgTjrYese/1RIH86dxc9figb+uda2S6qCAuT4hBLlrXKHXKEZSfu
PKt+LxMi6vvdQe5DheT9sIshqImbBtXFDiVw+TeYD4FvSMGoqDKLa3PXDnfntthg
r3yRlkQROA547Zf51xBNl2Nv747jfeT4jiAmRGVEHlL2gSJ7abtwvHMygxQCg+UA
weMeljma8jHL69ieoZhn1icDy5QiA87UjtoPj+Swtz8FxouxQp3MJb3xOgMla+sX
T84hwVOZ88i92qkAPWw5CIzlFZqqSCmaFkVI+JXPzd45sshfRZMxzYZc0/9bqCQ+
9tNBt16e5zHL0Ag3pxV7GL0iKTbiMhipPZ+55NsO40KJiRdsq7vuJB/84VKDnmae
55bqbviEzchuYD0yxcSlSv8jww/c1iPFymBwyu1qsMzlWaikCOALEIG4f6i59DpU
yDgOs4pfgKYzvmrGxBwMc5yvWnCGhrYf70PJpg3OMqgaQ3TPlhqQS5U1rTyXb59X
srcu7rocEnpML6gDWfvCnh4VQucQZsqhH86lSnQRl1HEaVQEtb5JyitWIH+lIk/h
WGvlkwkI7VIpDWCsIFE8zytkYY835lc58v+ucFtLCxwU59cO9hPMwtWWT+2KxH6p
ZWRb+YQH6yh5vw4ury/JIwBbOUosblfayUd7Dcco3VlH8J2KLBuHUClNvwWxiqV7
z/sbZyM/rQOaB/R6pMBairOV/rW/Aj7SXG6T2M9Ns4ZpDaae6P1GT94x+MIai3iC
up7hZoFqp0fzp62KYMDEZwtztioO33BoCSzqxgG+HWNO6nS75vmZfv0/f83iHpfP
n/o7xGHSvxj9SJtu725/PN5CmP0R8PArsEg1XJZhJf3PrSgscaWdpeizGkk0mq6V
4Gl/Xdm6wCKGyHXVdUlJPfdYfpB/jExxVuM9RhP54l+dx3FIBdMQsNxFTzCzmKAy
w2blFvmy9Z/Bre2nuiRnLX8bv7+VNvSyVWUbK7wjZGIOTeE8kYHOQPM3++CvgJkp
8DHbNcrC5jLb+w6Z8i8B33vMjIIXdzww6alphowAd6KPsSMYWek0KC07wFa3nlUE
x0czUOHp+qiboGhnYjj1zyyThcVITDHWlp/spHucn9BLmSn001AycvLPIggBlfAp
HdsxT8lmKYPpJtWtPhQz9lxWJKUtW6+jSh5rUh82pyYATlWiqbaW1GIkLD7jAXgO
BS3oloprHCWzKk7trXPgJlg7vSl36dDfuT6uC20jcsAnikMG9kL1CUBPRZFSGCG6
S5jFMoI+MvMKV9oWLmIdl6Z6nIytIHO/Qf53ECTKY60Ts+NJSezNS+A9FL5dh1xf
K+ZiyRHzyx7Terltpp8oEyY0eDyYY2n41FFxcIw8mLfaxpu6YfQ9rEQDEzqRDN/F
YGNrHu4nP4ZJCWdhrSbNBpw15r2de/1GhZHV9C43vuv3m041juUI24s2aq9mDH5t
5xq9Q3W4xeU2hXq411PfuLqLHqxEv9O+pwEaKWprCysUNNgSEXVCiKbc4BIsFeWd
3avPSVFZA7R0iIiXj60VB+wrpEd/kPblk9xdsVNNwL7EAAmt2DTObmLdLptzfjtR
53TLcqSe2WqCszijIIUrGoPD6nAU1pojZtScLt7HxgbBJVA0IzgM6Ajvzw342h/i
sbA/CT+o4kWA8G6BBS24Q3fz0OvLam5kKJ7gnvZzakBJ/lEdd065XU3/9NNs26zU
6hFVmL8nXD1rROXWYd1OgGxSNSoGPM9pbEXKCuV7oUcxDqzqulwbNiGnxZhcuQpq
k2CPmjousHJ4SpwSF8Q5bi65VEoIz9CpjGFjQq3y0V5av9x3KonGFlFOsim4bkts
HlWJ/aUSMUY3Tkq2IQTGF/lNQENEezI4ETD6WdwiU673AmX5khfbP+giAPri+x7G
ErtWEQXq0AkJBAt5Joz04aYVcSacRTDiHrH3lpREvB38rZh7kTJ9qWpGl2/EBcyi
6bGYw2L0AMFGBCN+y2uF1pzku7YzErUKS1SI2SE4YreRru8gryIYDj2KuZVH/qPw
Cmt7Jh1ROUN3dK4YskEFkGj4rOc0auO7eLwmMZr7k9CWE3GfjpykzuE9LEoagmvs
uQpKXjNn91DaGBtUGnI8/9dOY7Oed1doF0g9PZ3Ks+7MNLdPEBXwJIdr1zRAwfAv
sXZdUfHqt+Ku2CKMD7DP6ixNfIM0/anRNKWc+42i51oolDDtdIZ4rRXBOa0CEAFp
TZ6Gq5W/yFD0vIJ8KXNmjJTYQ94nc2Z6L4FTMxAPGvDTJy4lpnlnOp+e0E0eTASW
doIP4N8RAdEBkKBVu/PONBIgnV6W5+VVwClLw2vusyeiJeiDoKBV85oY2dHADv+2
9cLG/ShSwnhv8u4Aeko1GSK2WaMkXVRcgj2ixcvpOAx9N+IoF9OJbA8O9CvxH+kH
/Z0ceVZO5pHFTbg2Dk8hLh6KjG5vyCE6mB4rmEBFe68schTjld3msIaGJP150taG
p2gtBkYdT+ylp47a3lDvXEs1RlgGdmn1xvZn2swLjLV3hHit8uPZI6Ge8Z2QGLeY
qB1GMHredQbSizM3jgVXsW6MKk8sNO4RrP1SddDA1PvCuSzfjVyb79nW6a1gbWzC
Zsd5uJxltzBL2ltaJ9QUvdBFzfNbvwOtNhgEojgVI390YiwVglgj26QaoM0eTgFw
xG1W4XPnXf7mhAfOeHiRcNlA4Vu4+nIkn9/Xyd5XlL4WNX8LvH+wuj7hpGKRbwxV
1tso9WetmKS11LSVMDHPwx8L0jEw3Mr7IJjZPmlaM8tgVk3mB2ui3HifWeUENxuD
Uhs3D8OGEk+GR5+2Nlu8rwwOtMqAECX0Ell3gOr4Qn7wan4iBVNuVdU4PscSHIcN
2NRRG+Lzg4aJ71acmm36Q1prpnq7AF0LVmqfVECTldn36iSmv23iwvSlPueId8n/
rq8GYuiOFjrWX5y8v8SCE5nM6B9XE/QyiwuEvH96CnF34uiabSfWSFssbBlyPFAU
fnWYMKOYHfU/ES7tNu1qHa8SH7S8MmHM/KTrIiPREIYldav4c5Nx5rV0HY4wGbRk
Cir3YfT0vhztzt3puPzm3I7M06kjErvXMilQbp81CE+jLwNAaf2ihsuoozLb1L49
b5b5AZzF54NPec5J5+Ml0+PnEDb3bGHy6vNehSL+yXK5RhBAvSxnh+I1M5RIsLqg
JCvs87lU8R8Bt04ALGy7q39uBSPpNzyUJIvFMnRz1k7FITO0nmMme41V2SyDwcUM
r4SETxMi9JNxvhsEuzZxzywawPZ07RJF7YuiI/VCYfF+XvVGUfvOcJUpyeUAYaNy
iQofIIKSDd2x8bi6yYkNYoufrq8DTXbiInd2vqx1d4jdYbY1dsydUm966YKC/gl+
LdhFmYismNOLVjJ78EXorCX9eWuGkGdcu/U9yjnjrDRK6ArooZGY9hLWcT59ipaM
yGSKjJUlo7SeD+xoRpN6oDaqtWmUKAZ2rwrs+7nVXzgzFdYfHVIo3ct1tnkkwuPl
Z3nu2NX1IYsmO1Kzh2pIp6gzTJOUKNmoGxj+XSMgns4TtL8F7wik2/OF9Dg4SB0P
Ak1m75PVVHAkoJ3pK0+erIg7iVQGayYgxVkK/9e1VGZcg1xzqlIfTCVwr4Ih81c+
geo15vl+9Y9cVQIu3l3K+25OvsrLhVlaPUdVB1i8epgOWb7g/5ffgrrUAsuRBPI+
N+8LL/9vQQJBesujb4xT37xWnenFs6qlR9J+6pdnsLfkCn+oW+RJKZht597RQHEG
e9re+J2uHm+MkWgIlHCXbkv/2Sz5OJVA+XstaZrr3tCmv6UZGjC8K7mZAvC11UIP
7MzawLZH2SwwJZrNjLZXwCNV0HSDDzYAPusMhfmH0b1VXkhdLfPRVf/uALGZao2o
LIAhqq41DIylOO2eoO4gnNYNj8x7LrHgYt14m+cEXA+PjOrPkFBZmz2yvQf88KoU
uJBTsHGS6reTlaL7JwHVnTIA+0pLGip4ooO0T5bMNuuLy2NlNbt6TCbU/y2r5w3f
mJMWEt0NxG7rYxDuvJsrICqlCb1FE8oyLFb456R3WHSLWx/kRLwkdl8XQUWpwV0B
6TBiu+WC2rAESfxxvgJuigNj+6ldcl7ctzompqAleU4cXfnjaOYyyBmyvyQ0bVay
TEz2qV7plyySEJQn84r698zGju7VZVfWt9r2vP4ZyjWpku40QNSOkAE6XOGGBztr
biih/DTOFIWPJc3riYt0u7QIX6va6g2di7eOcGqOtQqnTkDVx+yw2cb9zZoeZkrR
uQBm7yMmkolh73A0ePnkXDQ34SKZqlX3GW5BtgSDJ4Y6Kkix5ZUj87Ous9hnYq08
wdePOr1mQCAMtY38MZbwSry9eUatFGVUQAIUMKW3K5vP0mLXNYkPX1mrwwPeuao1
kIun9rliQNn8sbq/cN0XNQdP3azQrXKD6U8o3K7CkcA6iD9SEU/F6ByTwT5jLUnG
S8aU0MVDzcle9MtaYZvU7B5Gj/fC0hj+w56BaZc5HclxzKpWg04mkQa1U4hiJ1EF
c2qBIp1qlGxdOZGmxQnPZPNH9tUd9zhtc7mvNzEEKdg0UreiHF0XEklk5WSMy2er
DNukOY2YQldNDN3sPd6B1E4zJu8Uqw8j7pIkbt3fE3vMffoHEoJS4kew98Zt7Q9Z
zds59qoMSCatNPS/39wH0U/KPPI3Hv4C+sWK31dqGXRG7cVtO4ZbWFRU7DQoHnOh
DOoosOEcCZ1f8xTOTjWp30zeceotwl8VT5H4ut8BWO/cQcblAGyZaQus1JgQrmQu
ht+G0558BD+2L/wGOrCLrv5/0iEW5qS/8kQrKOjy2Dwe0sSRuqBB5jTAWqiQT4XL
kVd7mHPpUymFOCwwvSYOeHknYss8KEhSJtOi3VhD70TvF4ljFqdK5yFc9bcgFj8w
RUn68ar3NlHlA9r8OMhBqImbr8PtslJoLZKTjQTvUQqNf37uePBt6SeLZ5tP2cqB
PNFrWFxsXY/b8knbpFmODu1tupSX49ZwghbmvJsxbwXwFPiwIwCou/DVGqQiKI5G
lTIcqVeGgLDTc1sGHQyZhg3FcqA+wNd0sn89KcYReKyCqerLnRlikAxw7oJBBfK4
tNjKPSpotwZs9uWFjbNmVFa0/l9lUg/x6cQpqER90Geqk7bG4gG0TSrXjlcVQolg
Qi/Yk6drHHiVr38ap/CdAaR/PviymYSDPs4WcwPDm5+mPl9OzmWambxcjpJ++XCh
8aAX+MWSY3zxVBl8UsnM9orZWugewYeddrNYEi808GbQaSErmhG7CLKRG6uAev90
SPC/O5Wx4hguXxzqnlKxYFJho3YQsfrir5z0FkTjQUMNkjeWC4inmU2OxnrFGM8b
wt0XWe3hWPq1S20euz6l6tByueeKLdRo3DooCgYjcoPRrX2L8uZtGGqmNLdGqwPs
0xUdeZbkQxFvcJgLsWE8irI5dpOdrIJEipz39W964VwfmVz2/QzoZRZUa5CqdIas
aqvbeV9V8WXj//z1tPTdcoqOX3c0dm4oG7OaksJltXvjNbNVTllsFXZ25VkbuyJ3
Er4ijN0qaX8xrBVosYKbAQ==
`protect END_PROTECTED
