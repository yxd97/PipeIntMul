`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ip2IWIU1ErUUGLc8oJZIzbQb8MgNw3OrYSJ5PMA+RavfVe0lVRm5D+cLIzfe5Fdl
wC5VPG7hm2UNDGxqI2ykY57ERlVJGPX//ab875pxTFG0pn/naomL1FMhLRNwNlGc
PjC1oD9Y+U0QRzsqGdbmoIsEq/zF+yh+fnftVerlJZtZ/0tvljF/m2E8JmPirc3U
OFmBaevwdpRP9Cp64ATqM5nBqlUye/XDZkmJ9Si7jVReDsOuJyvCOMbUHTHG7szm
q9ePH3ct6Kc+wdDu62hvuwhoDSujZ3Q5+uhMGrPxc4gtMjqIrEA5uD1roVe6ZyhW
hzbJ1PIjBPik7Kt4H4xLhB8TgzS1VgLotey2VFB4+wN4DeqyVRw5Yw+NOhCYI2HZ
ZId7bWzgAnXHFo5bvEonzY/DwlFZkPxx7zhejDH7msexo8ocYeeiy6ker8E2+die
`protect END_PROTECTED
