`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jIeIwoJMpU3YahK5jkoEvQz641r/ZdaRZhmHotjgC5AMuDe0J72nVTp9fgmtdGXM
MCwWXDNDfdBW0ydCKS5UB0eAZXz76BQp3ldMVAgiRXbj2VZmHAZ7lquXO+wcNC+C
+LBOwDWFF0qqSA+pdnQlqKojPwvoY1zj3VLA7N+a7hM9z6STRdgRWJtn7QYUsoaf
MlTo6oJipXFQaWMLtZqOq70eh1/gSqjpoWJ+LxCDxQLAIxuSkOUSh+Ruyh/Qsg5Q
1fyQ2bRFd5KwP61rhTwGOy0joaeqQZDYGQfNcsFOYQxwTH/2uEn5YWDYQ/91m2xK
WkC1yYIidgohhhF6AA55ZRpSOi2+fDW6dJgzyA3XEuGpePc8XOmIER6RON0+rUeC
Tcjk4VawqOiysI62dQWZRVvmTVoDhQyI/yXfjElQWmMyGy11bsnGMFB2smri1WIT
y7JQhsgN2ouOJE5LYv20EhLqLBZ/6iAza9p8WkgMXtAZOpB+5e6zbgf4jq6tc+NY
3VDuCIMCo3xFEBvzoPPo1MKGCkuY2x8k/kImE2xBlYsXLnkp0t/ts9EtYtPVv2Ge
VrrE2vxTh1zOpVhLKjdh25cqpWmLu/aP9dw7s/UY+HadKREn53K5cG1Y38Poucxm
JV1pkYsMWiDpgxwzogKmm66j11YH9CwEQ32mdp9tGsA/p8vna5JQX5GLC6kokaKS
Pp2ugrd2JemTctbrJitrONRtDK/RkolsLfinZ9MrjopQGB/m+C4GukjfvJ+/XSpI
6tUIux5+w4dQy9uW9K1Y7lWcEc8EHlF3YXUGyRN+l6QLWHA50S0vmn4gLWxaYNmT
7LJUP4j3GVh6pvBTSXtXvA34KIiVERqabTo/w5qRtvKPVOGjMVg9RCH6+RXnNnV4
AKZewtm+Xcj0alL+AhXRu1cHm4HtgiaDgr2LAO5p2yoIHgEYThwYErbgQQ3o5FLO
ENZTGrDWzjXGPX3yYhYIEzBhflFd1x2eEdf9z3+6JIKpVP49JhhStJhPOLGJ10ke
N5GhuXfoNTnHvh4c6TBkVBpVw3XNdNcyFNgkOI0zOKMG0/YVhLIgvMgueDGcemhY
p8GF/L9KMbJJo1iz0LWyfqIBH6MI3X4tamGIR3s9Fd5q7axVlsERw96GTMybVgV+
hlVIYs+KsUWkqUC6t14qe5Bj7572bnDHHnvpVW/GFCz2cjYLfOtQGkofM4ki4TJA
kUl9xZdLQkRb9mT8cj8beA5ET/OBek6/O3xKRck2Xw+qxqvNx0ZdjJWW2Z/JIL9M
nH1rA93PvaA9dV/jrBcKnMTNA/9oPYkQND/NO0/PRb59Ug2g9j67twFS7z9h6Chm
gS0+M/TTgIClY7RprT+y9el7k9AcGFlzmjk4zfONtyWLiyBl3MqoyJceVQmhJDpf
CKLn6VYlyPbS58ZRTpz3X3XEGclV9yPPnRP/mmaE9dOxlVsIzNJtFMgdB8Ub1Inx
Kod17xSvQJvIWXBlgs0Pq7YQ6WNfcJ+w2FnBCQd6nNn/EaS+UL56vasMhDViqxXc
b6E7nBNruqC4XQFsd5UBD4dS1N7j3pjXQeAsqXWn3ZTF8lvG1rTgZJGofqpkoNqm
p63VQSiyYlcPDvWMxdiNpedmGV+J4INbxRefFmlWbMy1gPCdG2lltW2AmXWT+kQI
jiXmYvvCH5gUrR8QK8rNTwsVHXReeSXC1gS7k0DxJ+Uoz3LklQ+oxP07yTkGZZfD
L9vbK2R9lWigTnu4/DheonKWdT90xSv4bVoH+4QS/m3uNf0SQj6nY/0Z5slMIeoa
pEqks9IXSMw5zxX05eiZ1FCVHA6tueyMF5U7+375yZsRfTy5dPrcqZHpGbC3xpv/
SZ71Bo2XnUi/535EZss323+HlZAnarLu6KqKPzZdEx+eqNAV1QMegtQwGlpu+WYh
OLpOnf6l+FCwZ/PNdPNSpr8UuqoawPelqfPuqkH4FMBcFvyGoDakRD8GNMl47X6l
FzahwQVrHRj3yXi2WjUrF91GzTPHQHKdu5EacDOs+4MUQKdX0klJymh8a9M5JQF/
Ovtuh544sl6mGBFSwsiUcS2W7tWU8mEgWnNTn6+pan4s4QPmxYYY0mui/QVY3yMR
jQkx3ZYgRXFLArf7X3ShLRVHweFFdYiy5ZV7JWWcmLGh+WU4wsIjmjVVuNn6Hw3E
UzH2CLA2DsB7gjZJvv3KVUBqNlvAMiPaVt8OLs9EyEu3RL56vATcLqfOv+0q/4n7
3BzPOblq5W/lOrK1p/6Z0swxJ5U4glEwe5miNB3TVxgJ0S8Jkq8a6eAVQqWP4yds
8txNBljMWt0Phw3jWd5jdKTh0bnqRNTqvQb3J7vrOnPr0XF5SWFxkynZNbxOhRwn
/xHL+xvSSaQOoDPX1osRAvLTrOu5AeWtzahT1NGdyjzPI9Ax3g0hKo3gLfw1n7qs
+oj0EMVh5LFbZhqHR7QbZBMVTzoPYF5Zb9An84QYKwD+lHbJ6lDlj661cZ9Sd6mO
jGuvk3C3Gy4rVUEHcg1ndUr9Zk7kjkzSz92fXsM3lG6j82Rvmlh/2PuBGcxE+lpL
JJYi/LdXz+lx/T1t32GLqDm9jmOtNcZRgPsLpVnh928dFyAgR/JjNkef0cH+a6JC
4FkkS0Jw8RD1GxXmJ09q5plU4XZnkGS4351f2n3D3zPfjE6Xyhux2es7Cc5ty8VS
EU2W+tTOB+r13iOVdMWETKgrDqWnjsAESjl4mD3Ebl4UCyPKHLBQfns+wsstll/L
pwAF+t4LEWGifl9a6CiM6ly+MhYkoKZ4fhRzQTBbzD6c4QKzRFRl2Jri1wLfsXMF
zP/8NlSziZi894XihoN7+rrZ4lP1ZiKIzdycRGlEE5dEVMnXtzpHietgyzQD3Raa
fJQ4puHf58zbaFlRIdlOcPfmXi0116QdnCpC7R8gQ2y1Z8NVZ/MLke18WNR++w/y
qT/ECTXD09kc9Hj4+gZgpvE5FTXt7g/VsTCwnqBgaStue5paibTSa/EJiO+bZqlh
9Yzhj0MRkp9xKEHFFD9jRn1TuFpIqCrW+ufew1vkFUYcZRBu6O4JOdNAMLisU7JR
MQzm/nKInv8D3XklD0zLX/TrKyHx8vPdZ95OSYK4nix5ihHcpDktCAy353qIYupG
4R0VgVHmlIvKER4OEQVdIlrIDVGEFU/RyzObTxePMljILdRicJ5N+hFZh+2njYDl
ZutkuZYabzcjj9HEkTsqpn3j4u7w6Kyi0H6VWyewgCrVwwSEiPt+OYstbNe0ZF8r
0QV2QJe2d0SDbK/Fbd5j8dgUqF+iRXLgv8nHVXd7ppFx5zz8TngXHAZfk92fxIDZ
NMWyqU+mV2r5j53w924HN+qP8n/xJEzwqs0QQZ15JcWYTMbBvWijev7iEZ6ldwGZ
038bs7oGLmO9M7xlVKCC7HhR6pQJPQa0S8iZv42/0GMXq9iad5plu3QtkOWsRJ9v
8hYk+Yr+2jR1fIrAXsS/FzzYng4ed+xFfvxOszPjs4T/x/i0/PnIcS3nIaIFlPRs
lHl9cKih+MwRdRICofza7cIxLNZxHXVMnzEXRsVnYws8XEre4lM0IB1Bgb/abRIb
Zavr0ERoCSNk2+Voj+P6W0e+dl8HoK7jj3jPM8Z/BvwC0FpIJJc8FgCUGg3o8GjG
RL3cuvCrhY1XMxfz2nudfDyVs6o46qXRhEEmEjyaBnvzUg7uJmwjU+X/pzi5zzLg
WvAfr79yKgvqcYb1VW+UE3JPeUcTxQPkZApZoF/WTNwangGX75qj2vzSAV3vs27J
IVl7o5QGJEYHXJBb7qEo4d38mainlVnKZx7qG8/Kz6ZaVaSukK7WXSR2mXzywy6v
VtTAnIlqO2tyIhpvOYzdEJHLefVyUTVKORKZl3nKSljcRUvq1gOOlMEu5DjLJGCy
DgyeRvhyPDYFE7XcOtw9Qp7MRS7xF3FYT6+Uk5YoHjxutLMlkyQhWkVkf7i5eMRa
swdQw022it+uZA3OoK/JFsmFwB1GM1GTW+uIiCyippawzAeAuMbyQ2FGVFW58g3/
QSdwUTNWaMhLHW+fEDW28fuXIvQuMRyW/dLhmYaLLvEdbMz7iBSpQdHz+vZ7kpOR
joCOudeiRHPcF5kdijO4aMTYK1lgTmmg7FJoHCoWzR+SlWhoyvyfH5tUEgPTUyyf
rjatgg6O1Gzw+/imZ9aysmFnVjzD50klR2dlhDv4t3YCyLnOTxIt9uB3coXT64zl
n9wvFzOVk9kguyP9GVlX0sWj9U52wXfsZu12YQIruUnrjDfHqBaRdrqwTnjd0yFo
j8sSkFD+5R+aG1loC3cDFS1n8yoeH52xsmscqOAMobgK+pfnwg51BxzJFiStEkO2
Nuq/WQyNDxmVMQovt6Os7iHz61/yCtTRdlaciLkuq6l9EqdTn/Xl8vbe6UYSexbZ
MoaWDErdT8PXGQZi6zGcyQ3bM/79/uPvbAPl76GhWtGttOv0RHFcTH8YIjnudu+Q
CZu/tmkJjTUrItSOuFUg4Blu2Gek5M/iIOl66CHJSD4kg9owm5kmMirE+TfCMDQD
5nYw6OAAMLrKx6QzAup2Ku9OKmeciRFRo4ATQ0grPDEOUSNeqnXciuFP7qZqnZWf
iOLA2e2d2J+RJ7ZLlz1IJVdvBSX/PEsdaY3BG8U5q2/CnOnmdArrIGtMsqo9WaQN
2sk34xTZdDqZKyIY+iW4y6pKfQ3N6VpvcfMaMZvhBhjMTde6H9VvEJlvXuaye/xt
CQbWB1Xovd4Tm1DAWbs3U9v25LOwL71/ruiizC3fsNl52XwJ4c/QPYpWwLdLlMl3
w0E8T2pKXOhh+ArMJkeYrmnhPvoUfxswsU5VFoFMtAzzzFAEYWTI9/k/3H7jJUk3
WK0G1lX12LQBd7SjH/0V+vCZuI4ZiHjvCUDVHj1X5SVbb8rzAzRLvzudNto1HAG+
`protect END_PROTECTED
