`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cc4whyY8PbiteETndsr/Z9aS0slGjRHo7NWxjPQHVKXMnnBLVGHfBRkwtD7/+Wj/
gUV2iIxjaKBg6+45ZNxbhjuWoiAFkmi4YWlV0wh0eUuooKMbOEeZk5C82kT864U8
WcMwQjv6sYwdRBNRoB9j+dtAVLWdAaoKH/GQqaWrGSbe1mHZPjIlEFw7VTC7qpNJ
A1F7xWAbu0o17V5km30yCyGUUK+aL3arr8XYMAYc3LkJT/RPV1bsD54Q2LqAwKCc
VsfZtKXIM3wqMs5EPGpxE2Ly23CCSYfhx3rHHi34mn9MSF9yR7h0PbZH9Yv+alWD
yYEZJZlBYGbtfXTE+S7kEI8mG5o1eOswZD5lqKVJt0Tdp1Sl7/94aBiAAtX4tC1A
9UUg7AoJuDT27uz/xnxzaW73iuPlAayljPkxrDlT4HQ=
`protect END_PROTECTED
