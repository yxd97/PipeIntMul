`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/bRjGPs97i6eRzLVmjYzFA/OmOA0xQUUY/xD3/305DZE294g+d9E5wl/V6RQuAT
HZjpEtTzwSm+WkOetumgECIIFh753uQ3rFJV8yCKd+hLVPWVBk+lNYVah3yuygRU
/qMZMHIF11d1XCSaIAt+wgjluWVWeg6wyG1yxxXZb+lUuXK36qWch+IXmXMiVqPL
tj0j00UB1l1KaowRNSjaIWTT64WWLznrpBIqdHeQI0vjDnfF8CotnAHPV7xXa6ON
K9tXykesXmnlR8LfCfT4G8bZnZNvw4pE1423ylp/mQqibvDE/btDgDOOC7WFr83I
lZWj1iOAW1hJKwcGxHDBbksytAbRpgKTexvVZoslJJHjETL/GCLnvmZTK0HU61ph
VX89aXspsEGnTp5VLDwNmJC485o6eLkBWWIZQdMe10L1A+oMNaRvagqLaT7noR/O
wx0ttRL8DDHFuGWQ0HMkTyoGGYwdgys1KOwFi4j841zpBCABVysN9ZtAlzcRljDW
mTwwuuFHIW37iOTdzvUJRv7Q4RQRSr8ya6SyRvcYgKb7ybiTWpjLT0S4rePg+FRj
h5xp/n9+wYg/y94+6VL8NWfQF96cKVQLc6k6W3YtgRiZjLZjN9vmKvd/fuTCV2Jd
5OBZADux5X6iV6Z0bB9WZOTm49Hf4w3Watso8GtU5KpOocokMasrPQ5eWtr53wpz
YETSRqepVtyFSRoVqtoYDhZI0HzEbMcdLgyGJvHgDBQCkR6cpaixR10x7V/n2I/K
zw4W24uH+v//dZM7MnpsrvBLlS3T0rJmzfRk3skJKTA/WKtHidGrk/vUsvmtzGBA
2Ft9tW2d/s/+j1ad4jt0tQCqv+Vd/5TlDWQOS2V6Vwe0arWGdOLBFj+CnjOZQ6k9
8UsYzM4tZeiFmdiRCmzmvDAhJEwrQ/7WNCcjHJQVio0cH38gWMekF76KPZ7YGxog
IR7x3FhyS7afPAYxE7dDBsz9TNMlZZQ7Bd2sWPfk8ednisw8XK/oQaaNr4xaJ9zj
o/n8LviVm0b8y3hIDyncGbz1+HUkwhlsPYvYgf11GZ849v7d68g7zC/nTS6IGlxe
W22/n549cqiFbXbYkwf56hPaXMl+XBbzpTKr9QlxcM1+hafiniw34KRHCTtOrFtW
AUiW/QImXnr1O2caexTbIpYIx25UwpkeM4Vn52bNvO/pFJ89MSrWR32EIQGkaKum
EG8lK+MNnAW6DN8N7CLUdNPVVqL9yKzxpdPr9bI0gJ9kHyAeCbtvYZiYoFiE+9ZR
J89lY7Jnnhf7WObSCp0bRbLxkyMv+0JWke618mfSGa6CPFlT/RMfNbb8GYG3tYl+
fZJ0JfoofRLrZWP2Jr/Ubm4VlJF2Gn8N9sRspRI8lubpSe4xpx3sHPKN7iuAuyPs
N7M7PCZfrTZOC3N3T8ghDqG7n40GN9RHw+tWqfKq+q86tJGH0wKAzMvyW+e4wY+J
GqCFUX4vzE6jePh4a60m5+oC0hW50TAcrxhrGNAlkl7yA4kKxjy+umvHBbr6ENau
OJcKTXxs94b+QWMKf1miBSx55JqZsWLyxmmJ4ik4rgFDDyZYupPSRL+LuwifS5aI
CiAwLw9PDRfTmiUrD/nChAvr1fC0E3YHBpoxhYjgYkt8Gp1eeooD55j44f3CxYfi
X8aGJgVrKDKG6KH170Hibcw1UEe3aY3SYKt4EZT68ZASrIdWR5McurECrV9AtG+V
vNLyXwk4W+V+98uSRNhpKEJmDkwx0UIANaYDhcSpHHN+G69fPxhDowezVmlIeE2M
w+1pHibL1pPpPAjKTsjU0DJQKwskPIspyntr09T9Yl6MZl4BTtSTnr+U7a8IszzU
vQYzcXkJX9RUVIiK2+S/vVxQTjvYZTeab2YeHoHORta39xlIyAbJOh/Z1EZ6Qy/q
4wDH3bHIXV/N5EAep6HKYoExsb76bmlO6tt8AW/5dvjn1fMIQOStSNY6UMueXkR9
6hb8X+hajqa+bNL6qAIYyROj04nJudLFRGuiRV1Q3Rm3ZbrqKpPO5J3YID7gsvsf
PO210dI/CnrRjcAztK2wvPybI6ZTyj/njMsJ949FIYQbrtKyPW0nw5aoXfYdkwmg
Eir7lJW1ulRlcMKg6aUiV178QO8nD7Eix+xrsPWI6S+mDr+muDmKY6YISMsWoASx
sIl+kNyR1jlfdil4/XiLtDkoSe4A3Au3o+BECTxgvyY2dmqQIrsRo2WNStVwxIPZ
VP08+dXeQoR9pDTvn4Vrwt3qfZ6RR31fGuYirAlyo+lgsn8D/8SsDiae3pmNfAr6
KnQxWrdBr2v7cDSkZUzYdQA8UUvyhGmS4fGc2dss/obIKFGEUYcd7t/kCAZ5jFfi
sY0B9deO4xSIYRRGmat/yx0GB3oJDCix/Jc0I6Q+8hBt/T0e3NJSoGAduuF6uaiw
TI/r+e1bVwcc5iBf3gZ37urBzLE1atersD4XuFn9bkqvRL79jWr7GxLyxBvWibj9
GgUUCFaoLxOwjjiONnfoYsDPBFngFBaU1u+Oj76XM2f9ZsCsIITOCCELdQ5jDhLU
yIHnmS/+XyLF63TM6mgojP3JSWlFxww1mAIPL+jFpHQUdHw99sEtojC0/a+a5wkZ
Qy5CCQ0Phba/bcBAN0iaTZLGwBPKjFgyoxDbmuuW1ie4gDIFUgRA2MrbZ4mH2pki
I8TuZyyI2OJ4KlN3YZd4gP5N4b9cTMsOgoW3w0TJPcR5KneIY8HmLKnLhuwyiRHu
oFFUUYpWKuXE6LjJiPdlO/kZYGmVczUrydsLPLnL99R8yP2nkctep4K9e3axjPq+
f8CVVr2Nx+0GCKb1A/PR7hJEgc7qAwuI72gbbd4lL3G0gbh+TqiRf11MuPTOff3/
7jniuE+fewMiGdzF1JKg9a9r96KsQQ/L9/wmierdvauQ1KXRinT01eR53vowLlre
IYF2q4d0scROBR8pSP9kTpqfG6hgRCAEV8G16z5HDOVt8uFn5e8CmlVlXZtwQEPP
PBEfSdAQR0UooCHIarG6wuFO5t9IB4nFeV7DsROtJ4yy9ed+STl8EhBBynWl+WmY
5zpE7aOiXv6lX4pj+1sq0sxTWTiOes/rGyAS4T+aeDIFQtmk8Jb3TxgLOZ+bMaoi
N6xwxzRCWyLNIaLfGbMXTlo4zhPRSuKbq4BSPuAc69SwZ8nGXRqp7frSqKXPpgFM
FzkfYwEsQx3rzH5k5uaQ8uu84CRyxoBDN1WeepkETw849KQKv6KYPRIgbpXS7fZQ
uVJGa7rogzPcyf9OfdtHjbzGvTQ5D+VogigYsmKnhOuBbx9FiU9tZNDr41YWOW34
qXUddn2wfSCmh/bFQjjIl9jE94v72asda8pCmc90aYfG/2e4bvxe/rGVv2QkubG1
dKI+pR5/6b/YZSVJMoXAXNKi8FXp2O/IBPAem2Za3OQ+iR1ahYV9Eis7r8ji7aJP
MsPB6ndhfUFuW4jJZzlRfpsjRb5eB0eUEspQ44M0PuJcSKatCMzh7GcpzxNsSpBa
BXiZyjvp+RhJbEXCkAw3JkFM1Ze/kgSiuWwBmDoDSB6XwOjQ8fOynZ8D6ZsCSZDZ
9PdRomQndkPVqSu3KyNUrZ1v8TjC3TR7KCnkgUXbqpcvBwGSJBQ6/30CwoILgxN0
0JMOKTucDv+9/37F4en0b1EQDmbZB0ZUARqMmgt4gx8/44qH2UcUZMrMlVtikPKK
0LR5N9na3gHz1vPZ3VBgAt175qB4HnwJ4CJy+vmU9Uhk0Z1yaZGZVX40KMJXzJ6P
L+UrA9qvFTZa1sxeGV4YgaLxkl4dovkASs7q0QcqLtaoEiBxOFf6TUrsKfcishZ/
0NNTqqaJY7eZA3OIGHbS/4qXs9vwtDAJ/TrBUb9UwKVACTK3WOp6bJjDvcehdhkl
zUA5e/ZKlwmeqyCwqZoaNPixrK4yjZjRKm7/nD2ErZala+4GFQSO4ND808KktoTv
doZlbw01T1ug7x7xrvY7zrh6SRMVUm2jNK/MWEJQXEVW99YGlMGTpin5vNMYNaYI
VBbGFaIif5fmT3Ggy3Of1GWFfpNEygJX6YC8Cwz4JSWOqyYNNAq+A2KvXK8prXOX
oLFwhdjiOJ8I5DXc1MmQ/t7Epo4xBp+nebWNWd7+aL2kXIlSKgvgMIyQ5oUIE+ah
I7D3ci6qOhmiTAJX/1rr4l7sj3nAKM/WSW8VhnvR2343Cnt8rVurA6YxxFXGvyUL
o3VsSWTWLyUIhZ5nyzzcZ7Njf46pLqRer9wfMgR4ySOK4HjVLwar/JS4p4+BkUeL
AonfoM1eoSNZ5sLaEJ4qjrR5cQLpWm3im4J5crDJXFAAAQtFRbXuxTFsir4j51fS
cAd/HlOAn29WiJMzg1zRtaMNNHeJKuqFPQ83hRfMMSQiNWtDL4FAhzAfmew8snpZ
SCemyyTjZ0lHFXzi7h2t5/bOYB78GcTgAovroMjCaRsYoaBbfjaK/uUX1vIQctDD
S14YSLJcdKCLKHBFFQF9OhvUkwS/8JIEyQ8IvLg+0ZQRnB9ZdhSnOYh9gmWQD7R7
1OqlnFQ7lAMAZMqFdxFdC5ivIojFiE2bmQLeV9HIePyCgpbMJZbJccStP1Uqc0V3
RwYJFcZXyjBrc0SLRBS5KMZE+ajhoM+eKXEsb0BHeLy7vYe+pF3koNYLUWDGhY42
PyKFkk3QNv3AsP56BXBfSU/v4O1CtaSW2D1yMO0nLWQdetvqjn+gmiyDq27s8JLx
VdPTVPw6StJM2SlSZuCNvmNPF7iaCo8g/iTp6yQMtJgqB2NHUfAMWOJAsLl7anX4
n0RcAjWJngy3KGH8RXM7oCof4GhyKm+32IOPO2YOXagNJdAZdFSAdhloKnleM1La
B8G22NBYKIGJAnS/93bMlHDtB1sTGuklB7c8iA31+NoKSb5fFr7IjnNyN4O+JFOT
Uy5OSwVz6xoohrtAc4S83SMxtYcGDjQb/OU/uJLMSxeww6Q2TUqcqcwEXzs1uP04
7haCKoHLyQf0JSsPNnmSDmeYSECPnX7gzRlKLvuZtNXmfbPyi8InEpIYHCiKnPjQ
y0H5g1tRyMOAb3BgCwPGsojSgsITwdAtsMT4LqPUF0vhqcEpQatEKFwXj2zBe2K4
dWeWm39n0l8HT8CJHataMfl0Gj69XpbWFCQS5Q7YWtaoBRhit/Jl4siayXWjdhk0
bvaBHvbelcjnrm4BqfFF6MkE6dfKHGDka/PewZjFfUbTfPr3UELU2nc6I6I6zCVk
LDyFQhVBAhNDg0MRfg3m1jXwaLkzSd1SsKoyJxtMxlxIzRkGbS4S0lviRPyZfhHb
QlVYdGqdui6MAoSZOlxm5qUfLGmCx7sGfe8Y8eFrOPVMCelQVQ2lxx3UoJD9/dru
SUWpUVNQBAL76gcRenwhZGGiAg1Vmz3m+3gJhqmBRficoljuUddDiZjpSJfktn6b
pwK5GUOhQUv/Sc2Dps4MnBFnUOi9W2A/LSGSkS3AzRD8ZKeyScGI+MIYqFhLW/7u
S/ijfxo4n7b0FORzoVJzc5q7tytghjy4iytTnGr/h5rVDUXAF5LUkDyYgIioLWqW
a6fhAI+NZzt162WIlQjbc+uhk2v3eRPwBMcygQVHKaBaEXY9hKBPmOzn23mIagki
76GoyY5k+ppbw3AEDFdoIX8mW33yBE5DJV17Dqg9YsSAtOrlHsAMBYYVVN2AVq3t
1NKdbjiOozGy9Y79ht4GKSsjaR4lG/zg9rSTivgnsnJ4Shlf/jhRu4GI0XTfgEHK
GkMIvJG/RUIkag5Qer5DXGp3y3GoftLpnrAUDBNAJe90dAbj6Dqyp1bTPgKoRXMW
c+cxTXIzweYf2mncJkNOBiHZis/PuHjcUOxWow7Bqi+4WtVqut+CHyt8dLDiRumq
ESFrzclE5kpFORjmF1dQisLtVVP/KtxpKhb/MkXB+GnJ6qigZhOc/wILZhwGmiTB
3fPZEDFato2LQlkbFAYF40CokTw3cZBoJ/014P7MBPcqVuXcqBdZip0yr50fecDu
OUCNjyFJzMD1tLhGqJnaIFIPwhJAv8k2yqOi3nsLL6UmrTXnDmEL+hHTYv5+9Rh5
1K5HBGV7NbI7YmCCyGHMasimGW8UQZy+Mp5vhQuTJSRxKHaiyZqUCfhyXXK+q1dB
0xueF/cN0+d1A6baBuET+0gmZet9hMnGL0aVwk9vZreC3YW9zN/l9xhq/KBLbxyn
YehAYSP5EmJDjBL5efdt7fBwxEKBWBs4RkZ9CsejJMVnCYVUenDHi/7FLWz5h2Tn
15mbNTd/HuYInsutN3NHRn5hou61po9I+lQdVkBkI40cvIdgXHOucXQmP7NflsG8
C+mnuY1D2SplvBcy8QbsdyDYUukJx3+kWdlAIeZyeZivyqAtMmckP0457ZZKgeTL
y8vwiVuGivuFOZ8JkT9qizLY6OXeMCYic0rGqkL5V/WoMTNViBXqgcqXGXFSM85l
3qj4/1bZrClDBaJ7e1o0alWAWn+8PgZDrZjOGqQ5d9oxPoY0D6oHVZztGR7uQ6pK
IHV+BT70MOSk/ju+N3TzX7w++4BfEyER9aikIVMIsPyA9WYQORMSQGaGvvbh14P5
OG284LFh9Dk+kkAwD6l983T6f4mgmUFaXPT3C77sZgc1T1VWovGi1pRwVqjgmiHM
uLG/ba0gPtfE4Uh2rT2ZO8Pqj/IwJcwKTfFeQLThkcqMWKL8QDs3I72ZzqOrlAty
EOYHImlPZKkGGBgWRgqTbQJ2OHzb/J3a0dLNy8JA7alN710CYWgBuudV7oiVXNXE
DGwakv6uctLlMdEFrm6HtRCoAwbMcGeqxolOeJ6EPAroHsY3w8I3vdmZPVoJgrZZ
q7Qq7JwQ5AqlMVUGxqFbbPK8vvjZsKa9k0kb+ZTYAASbHAzPJEI/IguPERr4zARc
EyJT7AXLSLdevFQA7auLuvV6LPm9TjauTMs3GUuOmvVYTFByQ6660xRFC1N9/grp
qu0azi3PAnm4aZf66yOEyu7mz+vVYQIyJr2hNTOyf8HXeQoJ1qIg6usdP8Rox033
WPOeF3xTU3/jjCQP52vc9l56Hm2MGnHG6NqGYXun3bnMiypO39XK8s6s3NH+RnhC
vjWUPFxlovoNXG4gXlk9vsNeyCCUFC/gOnNGFo2n5A1xrHdGCRPl8YrF1az8DlXv
epK+l7HzCiVIFNtd2G1k81G3B86hsxjAH+SF8ru1OIloHjc/Z7FUq9+Bhdtbad6V
slZgWudQaluLUf78H8v775YkN5yiARA/2BM8PsExa1pbiD0W0ugu2A8U+HLBty5X
P5i/g/GUshd4hMabTblXOD66xN1Wea/5jFuyNeHWgc+NRO8Y69mMOAm/7PbcAAI7
OXr1YzC7CTxssHcNDMmS3avuYnGV30qzYZxmiJIL/Dun+d5K6sBrVmJP1aZ+PRoa
CxhvylOGCAfQiwCgEj780QIPkLsCqwcqSDD6b9mobJ0NvwlMysdsdeadt8nY8YrN
fCJIRHRAQ27bweUvdt03kbphAZN2pSsTJIGbv9tvLGWlcBOIZdBgSgyk1KXTCXCC
I+gofkbafvBciGrZeus9H63RD+ybaXfelGcefy1hl0TvX7nq17TkeuDy8s+LpuQS
imJJjcBHBvLEni2BsaukGargZ77OJfNybgZsjIa7SS64B2mmjR3dFblNor1UJxLO
g0oWg806h6M2hSCLe3doaKCvazD4hAZ+3PCE02uum1LPEPIE/y/NcH7ATB1VrRls
xiOUIHef+KQjS3CL0E2skjTKnF/2Sa25s4DScmmRyDgQtWYWFlKmUh6tguFk4mGW
P2Dajr0jBtpnx0YpappF3ZJQh/h8Z4wyu9r2tYg9ii6Rs2yfLePgU7hQYd4VeVvl
VQasgLu1+X04MLdRpoK6HWx/buqObWeFz4fzr71lvSJXOkSEab37Vf/NqIpHzRHC
xC+C31Obhe2apI25ehUVAvp/kkwAUQxmXWOyvuANAPlRmVuI/JprE+CdDtkG7A2B
PR8enYxeai/q+L/M5QeY+shYGckaNl3EPXtl1UYH4uvycaVfmZTccYioa72D6wlb
Hcyp7JEFiukQbpeMFfuiXIJFFHrVOECW1QwoRPqUXb2QNJwdd3huwpodoMgXa9zZ
DWCg4FeTPsRjQFU1OrJ3O10vce18VGx1KkaUPfR1Blx7qGSfHQWC7Vj0GqSkB0aY
UpPgHKDD0IxFz9dnbQo96N45E22VZVN8m0xItyLHnZ0CbYEHUE9ip2W+4spTWJ4Z
xiIrm1hpJI46/Q8ThFOahncOAf99TQVYDNKHtBac2iV3CwThlx1GoJh3kE42OnLf
mmgCLLtZlfn6YECsLBexX9nSHpH99/MWn84rhZdakcegO/4jHtGh4Z9JkFAg4Bw6
CU9O+QxJEFEOwxQZKPC0Qbr0Agi7j3fbFiVhshaqNCB9Al3DoHYEf81zVXPUPgTX
exXC/HSj6zWV4Jzn4RyXFOJPyff2Kc1jH58ZwiD76nG2lr94W9pHy4g+Mp265Uil
suUqkymujPG+107hwVjU/RI+PrqYRqi9Fgf7nfura58eYSbkA7uQ8euegm/36r7D
FvbKYVrrfVKCMTTn5LdwvAwY6rnpFhvw61F8sHQX5CVPlHGjQyK3I06csDjNFaNJ
0BL+Tphi9AZ0tR92KM/hg1F8WIA5ILE4cDpW9ygh34kJLeRtElA3MLAWshfppJFn
3yzX9wv1cj+eOmNjK/mv3jopzMwN3Md/OEPDCKXQorgaVumuHH0AZzDH3/6LB+qi
7oOgHp+R2TRytJi8LgR6UKZSL0A/TBbGn3vO0XMP6ptyv3C+RbHX3QA0SJ8CIwgd
hbxOfpo07lN1fEG7IlZvfZ0F9cdgnIXud2NPKo5uziAKZudvaa7vLQ3ONXfPkVEU
J9YFy2h8kFK3S2jA9vHIt/p/GvagMkSbWfDZYfnzHNJ21gn6h9GOtK8+E2YwgRpe
8jhlKh0C+ibG3Bkbj8vnfbdzl0UGFGb9xXkC7R06+luxY1aWWNxX497FdwNUX57L
83tgYkd2N1JaEJEg/HrlwmftjP9GO7pmG9F7NQhCZFRHOp7ws/r62oQ4+8EI6+Y8
YzlKdhhkPMcnSOOjZGIB9iWIX68vCNyQDGo3aQlj9+CIh7Vka/bolVfTw3ORjwJT
Xed9h1HrlPow1xZXcDWaczEqcsw9KwxiEv3oMXy9iSX/MCXQrhHJAJ++r4RwHJId
QzV4mRrYrGjd9Ej6LUSUMw3azLHBx3e416kqNYMGaa1sQH6vNcWBT6xieWK6pxdl
zEPe3yRveTCB8aaLyaWs/79phWC0ozRcXWh7rGVDOTvJCuwTf5ug5CtObq8lEQU5
3wEMlfC+3VW0IX3JPdxQ6q22xGcqCV4+bNWVsGDkZ52k9KCvbTy2Z80u6pQ6DAru
8HJ1c5ys9xFprY2aP6MwO76gsD9BydMeylM3XUVJjelsdd60tgYZk6mBq5/cQAM5
BrjwQa4ryJ5bxelD0hAFwied7q6LirDbej8FCOEu9TGGuk4bLXjeZF40PsAcSEjL
D9kSC5STXlJgJ6RG5QPRHNZFK+IbnoIORgv9aNrIgwnDFNmUC1QZP6S32fM98Luu
lQ3hUhllFUaD3B9a+G+TTK/3MLcw46TeiKbF0V7/9UD2tELLCnhDkBhu9Ciq6dS6
xs9xb+qLUZyRS8a4Cq1wBcMa6JZEU+L1/EvPcyXB6ZUm3bORE7J2mhPplnO3Svf9
+zJaGYgE/ltgH0JDYeFA3pf/T9azoPlPKoKL0d+urLUsdk/VJuGfHrEmMZC96lfo
v4yBjzlVToiCuUQd+7YX2DAr8Sxj+2CchD0FqTXps2ehzzEqXmBzduWy+xCUPIot
40xZaT87x6hbcAfXc1efk95zDMERl9S5tebbY1kgY1A2A6e1u700lE/Z8DoKZtvq
tMRSvPzPeJHL6d9lNgudJRB//f0ffy04cyWnqopHsZOqKLj14ODERwQxknULE+QT
3DS51iRuVX5OVgHqXemElvEUyLPX481ywNzAfgjs9GS8UIO0PA5FEBGxOkg+qem8
mZaLmOftEE4YuQsosLzhJ2Gqwiuc7H3c6rMFDydvZ4qqh0XFeycIe2TtPGa7V3K4
zR7PedK3FpNMnzFTLHsEl301ZgtXkzzQmhVCf1dBCg9QxaG0552xjIKey881riW/
sGIS9tIh25kfMJeORis+NzrtXxY7ccdT4ZzzW5wFcIscOSJSyzvrC+hcXccIMl7q
rWnKWq7sQHH1/0qftwSuMlkzFmAc8MEZT+tFPGO3RITL4ddFKiuxhDfE2W51UvpV
T3gCLjHJYcH+QgilbRMIdh9+eY5LL68XaOuNhzQCMHmoV1UyqpUkphpfT0brURxT
+ePf/lTbSB0qbmKbdnR6SMx03w6D3r8enB3uYUogC4M50PuLKjgovDo344XVdKit
lniC0Tdb/tiEwysJVJfA9yE9ItmitIueVw8AQN6pjH5jefZ0qqsGIWUNnzkT04LB
UFflJ2QbY/JtHq64DOQ50+lkE68uR0Q0L8bwkm2Zrc6b7O7hMyDywY03OgtDBT1O
O7IdsSGD1vxzNE23kwGpmyDU4MXTPYnr9cVLLrGy58E5zHmDQtCfXSns4Cd4UMaO
hWmhmSWBMJ18lY7voj5x+WK00UveZE1eaY9JbzOeuHVIBoQFRzK+rQQIiJaDSWp2
snR/KWiw4IcOG8cXon5YWmaWPWPfbq1mkgaPgZq5+9q17sIhVp13m8Dp41u0u/pn
gk6CvlyvkOkzO3ZvfJKxsOwyYDLv5WyTsdn+h6jmbFMCqfQ3Qajjvd9+/HMRfWUl
ct/GfzIYik9d72SsnHsMBkWjfT5C+St4JfzW75nPXRkBe48IeMDc+QoU0UsIhVA1
TZASa47k8+doPFJ0mkhOSam6hxyAdmegA2ShBtcftawexUWxkMLxdIMyJbmrcCEL
/cdGR+of+70wrEQC22u7LioOmTBek3O9X2rT1bavieLwEn/ulLXFiXlKpoe/IL0u
Q/h1IGnf+CWgiPakoIB8v0NUAn4u8izCsLJ+qro0E5+3pZeobtiD5l8LJ9aSbZrW
JLim2O9T7gsMZC2ZPe5VVClwDNacvnaeYxJoA7AqcSSWHARDWB+vz0x4JpRX/5i0
PvhAH5Eh7uIgpksIoBPdXGSvHx7KtJWvgMkY6JkPYRbSbCdkjd/uryNr7gsKbEQS
SDyb6djMYwAYqS/nDIu5ZwvGJyAEZd1r1rzNrcUC+DHuZ2qABZfhxIz1/GzbAfQu
42FsIeYbeIGXCgI1Z7kKO+RkANZCRpmFZVIu9AbjMKwkNXt/WSCWZxfmvct73JbW
JXzLVsnlohKrSXxqn6lL6GPTYIZQ9eD+88CG16O89lQTlFo/uW6vjuhYcBAegTSz
1LKwJQAaa9qewjy5NHe64Txa87F42c/N+19Rqv1GYQgYA3z97pk7p5esnRFwM46z
w45HhDROELrc/MhGZ8rX/xhb2DNMytAfoPAivuFjuKgf3acP/B6gMO0oIJNYTsAJ
kPVUsFgGDYsa04YP7a6ChIHnk6PatG4kFDkSc9CuDH8opX5D5sxh9+dTHpDPYgY3
Y4ce0XtcqCjnWYmgpJOOuPhQ4seiL6/RDqSiQdZWvE4cTyWi73tZLWKtJ5XCyYem
7S5wSPOjE1RygM/UUT6SB30DJTMAAv03pSMc5ofDJy8owIt/Y+h5opXBx7eFDZPG
8pGmcr7UNpWQ1xTfhUAzcHWz1nsXm/FjIvnYfSE52NZeFkmJD5QvqXbU6xBZFWsB
7FKNbVBQP6NkTAYnlQWLwVO+sw6Qewyrvv/FFMAFV0nLbfELssC1GOQYdq7tiVj1
5Jfi33c+SLoEQMk57INjFW2+4KjTVG2Z1P8h3JERVytntmAult48j37SyWuE6Q+2
1eWOiZhKvGT7WQ/57Tb4u88NPWfPUHWQ1a86WNvJP97WHfeJB1Qz4Bp4CzXrZ815
B1xgzb8v+YF0BN0ky9Lk+zg71LJ8HXs3C5ffDBg58vRQbiqBZOb3PvuLzOLm/7Bx
4PWK1b6iArElGUJRtPjXLso5XXXInAtPQ28W4sxqvbiquFa0A8W+OfNh2/92nYsZ
4dIeHTK9aiLgV5zYXKFj0rioluBfNi6qL284b4/pyMj46J4PMhU94kME9VTt78+q
x8Ch6ekd4a1vamP8+lXSOdJ5PCGRM8tnVrK1/cpNkDcyyL1CNOvfP5FGycRx/2bk
CuXVk/cS7B6VJs+MfbjkEr/eOfP+tJX8c9zqysPLB3qAHdF5aAUrQv69OsEpDHS3
1I+f3Y1kl1RhDLpUU5xjlUw5Li4K3MVzh7+wljhQGt7xyfkB9W+NemFgq9z4zHQ9
EaS/e4lETa/q5mUqGwnKQLzb6fipacYUDrVopD8ueDMX1bCmX/OrfE7RsVPy2BA9
g4VADS1uUY2HhuXZFSGVG5NlJYIhr1xFZUUSbzUpq937Sa3BAJE6xe1vse9hMP+2
0AxwYvU0FLTXBV6jQxrSw+DCnhtL8B1/bPc7btfzaDV3GmIw7O9/2cuOPby0u4oH
Y8xgIco3n9+DHx5KDoLKZ5zh7L9vy9yazpViByG3Us6b4McWXDDCUCGo41xKg671
zYmK7MON/ztOIYbyMwjbeLexXjFt0TC8spotxLajbsi682QqX5foL3C42t5li1Tz
mDrD3MpxRkrLBZ4grmMSi1vV0g9FUpcgfdqlpXgDQ9l2ZpxNck84YLrkMVl7gmh7
pknTQhY4EPzZZWmhak9H9UUOJZNXCd38KInJ0gsw8cD8AcBrcdPZ+jBcdMUGTMJ3
LfoSnf1A+SLIEFagZ/7zaEgOvwm0fr6VyeioI4CMmdkO/m80MTx3dbl9Llp+6t+L
3OC1SLbt9xEKOh5ob/iq+t8AqEYd6jMF2LjMGrPuVdd+wCyQkxpXoclgVK+nsCxk
JT2GMSd/C9pFAk4NYiiHuLugUltnbvAka35hWqLvzITqygVSv/UGkenrwQjehLU+
RvHJIcjt4wQfw7uiwgXqBcA5Qxsq/Z2HcusIqetx6QTYOQE2m9GyVjEmZmR39HLx
2sCDUEgztCeQbCz3YjhgcBKb/La6EUbnkNYxmWsSkRflpR4SJAhcjFlZylXTZ/mS
Ka0jBiWLmdxVSaYLryGiktgrQUnp2cHfCf0m6yf2hoiMP7YZMvBHB/8Ed2Veb5p8
nAIcRIesQeRJx7hoV/SLv96YZSws7Z1QnVQqhHrKAspApkeuZi3K+KxMK2YNZyJP
S3xEm/H237qC+JFbCMQBLEPaezZQkkk3j3NjDZXxx5mhqAX2WJnvXEWCZ/6pRv3p
ORTC6ZP6+gU8Of1C8+l6essbcZZp20XGNnlLQVSgl/KDEOgw8uRAuRo9CCh94LOC
NLaulEDCra3KGdBBZ5cKe4bxLt+MeiRrFKsVlRtQtch2DIG2g9wuAjJocqIuJe95
hmUrUNnCQ/QkG5I1KxdbOA3ZE948QlGDMFG6J+OKiLrZ+9XBaH0/Zf1pE+fVYTIX
dFS5O+DqgobXkuqFdnIdEA4zbbTXYhhegabq6dYWnWPI2pixFToN1iOTkQvti6e8
lCjHwy9K0y6Rxet06J+L4dJdXcXb2jG2ZTQBDKR3unenpue36KFl+3QFGA6mwFy+
4k0mFQozAdKJ5qRzjnbLAonz6RHPE7ggewr+WpPF0mlIdF+vXgAjYXR6OhX56bO8
qb+MAyacSWm6IioM94P1dTcjCu7vFq55Vl8FaRCrYcj5LKeWVPkNhVm1rloplEzD
QJmAMEc5OYiNGOW2sHZ7aQfepiuDT8rLXwESXWwmoogabURgro9joldg6WBeTcpI
u6Ztmg4K1gPzdvQh1KPw6FDHJcC+KYEROnqtIwdBmgDff/kall4Qd2EzErgv1L/D
E1q54Fcn2MuHdbu//xoXpy/VhPRzJOWvpvIkosn8vXsuk2U1W/VtPt98gnLIGcTB
Prjc7vOP/uzNvhMhbS6M8ZSotcS+FCIeYTyTUxjtGXPhDfzO3fGef9geV63nQPOu
Rjr9Bmv6JoNMmYZe5XV41Jdl3kiGM7RvdDM2lzEWvNrYo0BhsVqXqd5WpPtQ84L6
2egBB6OCe7RsTEveBqhg8OwCPt89beIhS53B+9MOlSK9R0KsOl8o8FCc48S049N5
tP72REWRw+/Xt7E7oKCAqkQ8pWKkB0f5thD3Rdk/eRMywDDUVTuksY/obdYH1aTa
CmRpEfkZJK4KAdbWVLM56NuJ0799WFgbytJDaQNAbQNOanMb4eVBwAd2KULMKMUD
UcxiE6kPBQmpKTPOUVtSsAuYZA8GtPUKYj6uSFXTlIcAbpcm9ES90LT5jiYdacZv
aH3QI626V9Aeoj3UlkoxPXjUZNZNb7c0ccXJ5E8I/fDJmfj09GW2hhXlCACQArcl
R7uii4jQVUxjVr+I9ID2ne1CWQrOxoPXb/8bKRHig/WkDUvHJ4ItgMNW0fu9lhfR
e5QPe3lJbwAb0x0wavKhsEP3FDs8SJq5geujHIOxUbYX1Ai+Pma4OLKvRXT6wwgR
kg8J2TIJMEoeztuwi+TtymqhdnKGRr3zgTWAn25tvd/C9293XVak/rcNmR6zWzvu
LxPprmZTP9KI1xSXc4Eeu6TY5by4A/nW9dVM10BIE140ykpc1OyjLWvWu9TNiBET
z8opqszEG0w9plhOBE5mTPhwl86XmEGt8pvoP94G91SM54RvcaITf7FmaIsWX3ZY
Mc7CILDchEweEXlMTfGl0Bg0K/sw02ljDKBmT9lwttNsWt5yLDPdmIBzMF1jj25y
Kl+q960t27Kgh7IL7TxMvgfuhBBXimSvUrkw039lJgoyRaqmxxWKMsT1nsR7CvRD
K4jjszT3uyf+LO7RSZHl8D8O2nEHJoN0PZp4pnh1QTPJ5yQHmpEFZvy3IiT08jxY
rS9cGi7yndzMyy/8mQFjeieEG+SuevudDYA5AyKewFPG36blHQ2dU5hHXhP4L1/X
ovjCQyTPi79oMq4ckikPORQSYi1fHufaBDh5oE4CIsNEEJuLq+jnqovRrP6xrZFi
0sO/VwhVlMmlM/GW8W0ir4sNR8xgvuUDPkw5Zh7vB9IfLWc/696ctuKVJD898xzr
i2xvYjwm938jZ0iCUHieQFXwuqRnxjwefIjTK0iNvZIjUVhYJ/CuWN/+aNl3Oj5X
g69XnQSDOBM9eUNcQ8xPX/Ki7Cu9K5r/vDV7p7hxKew+YZfXe6WvtObquNsjV1to
hSGY7XxqV3Db//3pKYmE3RGCbKLizJ82evFWqRSFUjshNP0qSIEpHeCA1PhE+kFB
yCAW8+kKkzTxBLXN3iZoccuVlnsEtznek+4VxyOcu/mnCBzjNKsM7yzqY0EjHolp
AbhcPGZXyhxH6PN+yP4KLPyCKuv61zYJEBIbTcy1KIjD7Dj5kFSv0ykQEUpR9KWj
qxNrk1m53qQqAiVuiezxtos+JK+EwhhhcbbxIMHsiBCCaZcyUIClXGMwTqFNHVLH
NmsMvr5XWVCTE8MCfJJHlZdhGtO6Nyty3GnnYmOHrdPReAvQPeY+lPBXvCsjSW/1
g6uNU7LIMEetDZvL1TFoskmkVuV1tv1kr9BEE5BvQ94q5jkD6M7pFehcgm7i0Ryi
hMHTlyRS/1KY62R5PlCTfL9K+8sKTKNxrJZUBu4kP7PZAYsE1CBmHg7lp7rVZ/DN
+oT/pRjRSl8wcYQobn1OlybBbJPxSpCv9TcgIyyrz7wL7lVGjaokAvILdZ/JwMe0
SNKK1c/r/kcoM3AGfx84e+Zpnq4gj2q2fHkpE7AkJcFvJU0dMU3z0A5kDXZY7B4I
qu/LU1JdeLMTPv40VJ9tsFTZPLDH5vWBvn2e2LyTt7gI/ow4R4ZsbSBx3bFhwKPX
lmqxdjyxttpdLp3e4NpEcLAOxFXiaWBmyYgnURPcWyUwSH2Bcnk82qjzbtkRMlqa
6jxqyqdxBBdsAnmvYC+8IEQ8C7hWI4NnWyzReX0aPbTwgkdqV2InK4tA0ARp7yvn
2a7WnNFXSADxktL3UmwJJ7E9ne6XSziZRvgdIz8EPZAt3yltTJCV/g0U+3UFkeb4
L+85JI0LUyAmknvWJQxOkcmNn2yrMhg2x4o9f09golrDLlAGxbaHXsja93BjOQii
n/CF9X+leXWqFSsyXEpHtq56FsYcG8tMxSzWUL65/zD+tnOlSWy4zjTkIfkvoQPX
HXGFCyLbqHu3p1A/oBajs8QsEQDZ84nx9Njem2EeC3I/0oaaT3NJvNWqaG4qSjWs
4jxy7bqpmT1x8Rj1X79N9gwjzA8roME5Kbk1aN4EUiIuSnpNH7CZzegThcFeHQeA
P5hs8MyZ901lRbdZ0KPBpfQRNvZmxmVdwwEKaaLjNBRpoU21QgwskvWj0D26vBRv
xrzBAZXIaZQ5IMLwS5IlczlpkcT/lx6pPBsQpSotpkdDwhW5jKHjE0RwSHdznBDQ
5Wl1hwa7Hw+bHvEGAn7dH/cNeJswOxxpoRM8EtmGhCFStQ/PdvpA4hFcJQmLDIqR
gMHZ0PtdSoF5R9KAipkq7Vjyu15EbRi82HV0ZMydoikq0gjCuoZIwE1h6ey/dP/A
hdyYcRadthlQhZqNWGPx917kZmUUPDJDtpeOkSj7bP4oTHnv1ey8N0/O50pOWZ36
Eb4zi/lFWVL0iLCsNg/jnI4GvLmUj064pMQHuYb7MfBGEDZcsIdT7rs4P2pw3THm
xFoiJzJi7KI0wXJTyOLWSUrDADA2MnenaWHC6uePXd3WTu82jmhlpJBr13dxh5la
bDYPWMrRr2VfVgVR2wlibLhSXo2S3aaNYgyoe8xNYc//LRICQDGYhhATpj1kb962
wXdGLa9PZjzZmHpWsrfmxdORByKm7Xi4rU6b2tAF9OQA0zCT1pgNWVuGWE7QyOB4
Y9XatpuTKBjkpzXWFV9Ba8jH2OaXkL4JTlQqqcNXNSEi0hkEFh+J7hIwc4Z1DsJi
4qz04XtdiAex2tseOvwoMzKR4jZwPcUVKYCgZvJS47lEnwkxzp89TSsfeJJH5qiW
hl3Do/9b9NDSb9TuAfiWCPcwMNzrTtiL80M62hsqypVMWumwe0l9YGqnTjqr10HY
uMfMMJ0GeRbNGsFNPTH9m0GKOH5PWtJzst6xH5fQ1CtFiS8s9faPxD/dh32DSyKt
7v+LE56LhC3jFdD2/+PfZQIwxA3VJsxvjF3UXqpyidxHCG9dFWb2BXy+esc68tgl
RVaYOH8hEOlUJoPyehwYDUOeFzAS7jC+Mjfgdw76J0QlPxsgTbg9o5nH4nHEDnZS
mgmkvwPA+fFPOlRdBvLhXpNiAZDuI2laWxefqZYEKE85MyLtZ55htDPbM6z+pIf+
3+JQ9OL9ekiSKYk8TkyBHn9DfibXgS/yU97fm9dPCWXBM9P+JiueuSFZP16mU3vq
fIvLp0FrtzLsCh+rqrBWrGm6yF5nEK1bDqI4xKmjUdmwD2AHbToRODprTb1EZx16
vmapMqSm1+b6iP3Ns5ww+XLJINLfNbglbaEIlX+2x54cflxboyy7JARwztVrC4Bp
eOL3wcRmF3Owrx09bykCTbhbosrBvUEQTzbubxV8eJFQlvb/Tl42dqwOA1xIRhf6
sfJGXVWwa1IfZOY6wtiZ+ijqu/Kgrq1mJA1ou+e1hv6ibeLTxD6UK+T3PaA/eAbf
+gzhP8ELMFYzbTK69Alyk8RdUYVapS01vWRDrnqaxvOFR9N71NMl9uLKyqyes6WB
CxIlpAYncp2rzssP+zc36/2DGveq7hBSvXlfc1zSbd87ZB/q1BHiDBLntWuX3MXt
cHwM8bjPjw7d3Vc/CwxUEUpGI2lgQgAMKGb2MfgZK/OMuD84URUCtB7i4Uo9KA9H
cdFiu3Fv+LqS+HPK5FQzEes/Wa0D16M1T3j0m8kNLT7zVJQO2B4JdrH0d9TwcXES
I3l086Ks//hbpcPciOJYgenYIKrGQ9Xj8ISHBprp4cP+AYfHJMXXTWjy3q+3ihyX
H79Q8yi0EhxzAPUuwLVSPZ8KcN+4SA19Ypy1bCBqbTGJAekFnsxkmZuOQw8p+xxa
JDsrVH5G4iOvO46kLymo+SyiVdw9XDfs7gOC+RfasuxJe7jMde2YMn5g+w7Z0R1/
TQRayFo4Nw9VpmUFffBd12DZy2aPmu9dKwCpltQOTpRxL/Uz8K1QhZSELXt4Pnj7
GumGWftG2rHctSISvIOwAHWP3E1D/ik6t8at6jRiL1Wicr5sWcT3ZEsSQAFPR8u+
HZXT/tfBKKDKsZPPIsiuWToSNVVoWvjGmLpsW1oHPvqyWpP3yBgXS1TlIC7yK/Pp
fbW2Lm2TjyeYT6F6zxDyWittHbqDwD4q3HWz2m1jlH2drpCqNV9VtHD6OySTyRxA
j0QP/xnZzRH288n6MyPgF1LzMF0uLWd6TsCCNZMXl5yBAen+NSeomHSf3eXLZD3/
TJaS90uAy3Chsz7sBrUvAntnPY1mkjzIHaCLA7x/35YP4LoVl5eF45IXcS7uHSOg
UeDmKf5/48gZK454u8PW/mw5OQFIVGESqB3OKFWrNAVjKTNORZOmZzOu7SBRFqbn
LvUIkt38YSJSEOqxROFi9n+sPGthh+AbNEj3+BNmS/8MvTQiRaUIzDHiHpiuAVIH
N67v6e5FLqzOHzhY8JwtFwy5U68Tdz5COlJQQYQwp7UpRAZ/5nAkl2Y1JtDAiO28
veY7l3Ht7nU+CLIk3nnmoyC4G8oqdq0nlzLKMT8k9ug0plRGUdwhU1wY0vV3NzTy
ABs6PVi6QGTEZr1oly2ANwsVSFEuB1HN7eM2JviE9oxOK1RoN41L+9+UmT76EUFF
KbBOWP+mRVQCKKYBUN4ao1tG0pf+RnnIil22Fmfz5CnA17R7cYd5yAP9ugYqx+5X
6RpjEdOFCh+oIj8MGdVUV9LH4ODpqDAIPFm6Zx9pZruuRKW2Oe7l4d70k0kTn5eJ
eIpZGXZGnTDn0Gl+u9hTIFaAy/bNOf+HPxv0ZqxrdskmnDjcdW3yDIcKukaa+QdH
n5V9Hgppf0+AiHmznSixUlRYf4cRj+4v/SjfDsrjJRK0vbK6wjI0AwzKYJ4nWjhL
0CFRmNLaVEUCtdSTZr54BMbeTdAws1N0osDES1FdxJXdeb9RuQ5bJDHGjxICOgVy
XOcY1wQJXhin5Y9iUEdV+GRwohM7vwrJ4Eof+jXgxAGaLDzFpQRxjq3GMyRHSbXe
5pnrSYQ1MFBNYbjKRafNVcdeeTEFbahC9Ox419V2Uc5UMaGnAzJmCNfbnS2PMr7O
I3W4DgUP6zWAQJVNAIidevQ8uemFVccCgEp6E8GtiP1a5FTXhskpO2z6uU4m444N
ROO25zuj3wXuEZ1fnfrHxptd83PVUASVvCPk/Mezq4SdXgLQbB8VbAm275MEvAv4
jeVDYPFpW03YBMeUpSMId5mUXP88zg/K/nafqIRnKr7MNgE6mBgK7Mco6RGKEumv
qX50sE3w3amlc4EKdkfNzuNRdbaIeVbnHCydq38B7YM6w4mS9d2QaBdCWfosHq4W
ZXywSWj1qok/eH9kPNGODzhzGnQ6QCZQQJBBSEaHb+TwUYlkG0nDkXfrWiPl6riF
HI1/DsaEHbF87jLBYFQmWW4L16P1v+7P5qmGT6qwhK8ecnECJ62S2B3bLdKD9j43
jhDJYXF7ENqZ2mw6KeLkFrsMc5pWybOifjB+P4UNQ3L5uEBb16gSoiMmHaHwmHzl
qF2+sbdMjzaulgEXsVpzliSOtuw7akUkbjEi2uG3guPlsQVdWm6R+imtvphzZSSF
RbNZsxbI5weeX4/Rm0zj/bHVQVou4g46FeZMnRBXJhI8JP3+ZMRnElAzPWA42sgY
iPCok5b3SFUs2mIPSrOjTlsl4Zaa2G5L0D9NmEvHBKTF0LXNh0oDXczwOtli0Hlm
5iGQ+UnMA7uSghl72gWgiO/90dwUodr1KZF07dDrncQRMoxVVI7uZYAk9KpcZZrh
rCgs/5EgvXA1Lbs5LaP/deN1Nn3dDkQq+jkcdbAwBnMk3TC/QEYSplRQLSlXCKhG
MTdtNmdxyUK4+SZMVrM8bEw9JRmycPYvbe3Ce7AaOHdLuglbUTg1VkVpI0DwCC6L
hPLCHoPjdnbwZgjn42P1kI+CfEdPufzipAKj/bnV+yrDp7R5kgL6qCRyLpgwC4jo
Ofugi3+WZgWBZVM8Uj3K/rMB10tQPMTJ6/gQUthkeDeX3r2BtIEooCk/d+qLrGqo
55GHZm5T+9XhFOyOV3p3iyP3EnXktLv1uRGLfbEvFen3KJ4UFJgmOqvk9LbhoZZW
pA+fU2CScKjF46oaU5Xv2GdAx5q0PszuG4gLQlRjuB+gT2AfMx/EMcIsiykdqm4W
fzT9xUHEOdA13rSwaiUi0nHWs0EvOz27eoAvUoE4uqh6mujSBj70fcK9RAM2l/5O
A8bO5GqF2HzmQiaCQCvdIPNrt0Y3QeJvWfnh04zb1g5h8b/+Ys6bodwZDzsEsvht
4wTlPePY2o7PG2/z0E/xMXJTu1QmRy8re4j0PF7sCL8dQMJlJAP/XXxFy++5O4oK
5t8XRYNwexk8AV/Nt2mARR+oPM5/MtpQrpW7cY3lE0Vm4+Ivv+xgQChuo7dTC6If
mXJN5vZZu/n1AJRHYgRjMqS7QccRcHGG6zTtdWiA09lPtxM6sbBzMLJ0UV0nqHiD
HA01LYZHrCynvq4dvZHjoDexyuZOpMgrz6J/jaKHACPqGPZ+VH7UCUa2AYGG0sid
ESy9kH9TpzVMpuarrtd38XD3C+uh6oCxp5SFXXvNviqxVrG8uEVLHUxxlBDArzfG
HGvn6JghhmOP/CKVTMyP6BGz6TElj5zsukL8WtuKrNXsnVbGGdfe0OaCJk5BvKz/
ZRcmI3k9Xw/C88TYVuYC9xK3Fi/m1aNtNdXtKj43xFPvd+npABawBolAG2PPL4KC
8EABNeBU8dosk/+XxZRdxzbUx7GImq9+UMJc11TexPeAYUZbwl6dtU1MdrRpFsuY
qbbhY7+MtRd8UKFOGRP69BJd+1DYT7hLqqVrv7Vq0/bfDDLSXEGhsi7jMbxnsoL/
mX4+W3um+NkyRSKU5XwnNhAHbj3rEjV1uDsFb4vs2FC1/y2umd/dzny2QqbvTeYH
q9OIBFJWsSaXWWuijKVcnR6liU0QGTwuTy4ld0dgDLLIN6NYFtJlgwfYVogq+cO8
yAxrsqGRA98YZn3jTFLvU5IOQhicjrMJRLDLwO7d2SsigDewJwU6WOdCXacpig8U
9wKpvQpkWJfZZqakqwwyXrxt/LrNbZv1SsA3wM9PnTQMW5LrjjD9USNKXQEICDxW
cnxzskSSfoMqo2jO/0RkG5SePLHAbPFZ8RVrvR3aRlrtkHGMck4gk7dD66MGgQmW
PUgXvItPHDUqMO3fG+bbWink2ZZ0CMJ9T52qiOtKrEvDZvxVn3Cb+EeYRVkfPJ4b
hQTGBKlzmfIFkXRUB53VONiy5CuNbeljK8ZvcgM46cv/fAUdmM31xvyVNGboKptq
XDDmQmg0j0+dHDeRMJNWRAHaGwq+g7Ydyafpbk3I7F5l0d8+FejfHUECVGBQBJb0
pS8s0Wr0DJq+fh2n8Zo4pSYx3tEExiDOJ7YfRrB/n44N8orpTRdIJSenSDOT2XMa
thRd8QTjUlQO+29UOrV0wlOpruKXgSuCNfzkjqUSLrT4h7WCf9X9vcWPVbLZYxoL
Ao4hsCDyMkoPFu97HDZAhDFP17jnBJprvqa8vzwh5vy2ucakuXGVWUZsn7yMY7CJ
QgdY2R7ZGYVuPnrzrkO42VeFH2JU4if9kt5SID/N7bYZiPec6oTyvDHQwT69nmU0
9a5FH2U5h3TZOmHxkF0hUjkt5511gyDeSzikpRJVpWAiT3riLoiT5P5disP6CkeG
uamtkx11t0nk5XpcsEARssqPVtTMTG5yvcGXvBYVbmFILSfxFpcFM/1prLA52oij
WsMmQeLUu88pQ6zlv0AhO+82OuakO2OTHJrDqtT7F1M2OkwLpdlYTKLhDvoc4JJt
kepLFSoxFaMC/oDi9cQdVg2xlYxGmLxlpFzr4WAW8hbUMWxKhHQcqAcwIAdnDXBL
HSnJcuG6k5b0JH06uOVVcL4EcZ3guQ62+1BwZFK6qz+laKQKJkTxt8aflAPG+tB8
IgQKwWRyWcVghEBxM2uVw9ofjbSGWuBvhszwBAgeoIGjrSM+I55caLr7GC8APx+f
kuhn84m0KeD8qAkiMRriwlQEA6ewIEmbjZjCGtlsTQdAjC45/8wl/WR6HOY6AqLo
7B1NgENVd4Hy/yZyQpBtZePXuUNHKU/WfCzSEDfQEWhQ8glVLc7367Cbgltu1ocM
Rkw76GvztjTSwRR+e09yQIT8+B1vZ7e+F3X3d9FW9yZcC2cj9vzY1PkGZ4l+HXQm
CHGGNOpty+6EZzsJGTViB+oiATeUNS5kRxObM1IcvPgt5CxwA2u1xPyt4ru3mza4
x4tMprqP67ctFC0nantZQxNgDU+SJ32r8ybbnQGv70pfqPpwO95hj7IULrFIf4uP
uEX/usLvjQOtTTRuqqFzI89EExe+VhNiJW3otPyTXxkSx0iGoui3vJ6eaGZHBOb6
GMiU1yDdHTOVI0C/K68/oe7Fft2ebVT0jFxil6J6bJmrh+4ONbKxqB7rG07IzaP8
B2zvtYVVxFQGkCp5LLj5rBWQt/eyViTVOmHMAop+nn4tyG5Df1gJNe5lTV7wXNHA
+vS8CJx9RwTTT1q9gFXA9ce7UdS4RplfMyMjBthrpMnc+0i69PuoytTJRbtvhZPD
gEYLlh/nF4esWTgKj/tpYQcLwAjPqqg5JmKFNmrHLi14QRPv4jRqXvsvcOCaZB2E
3gJ7BoIjmkm0XkOibglYtN80MsLrAGNVafnwh+TdIOYCE/o30eIV9x81dB1+rlEX
iC0Ywp+xkuWTLbc9moT5/Bsp6bfkycgNSq6u1POsNq5etqDT4EwyMt0KXCKmt/El
Z7uDN4tMbEZB2Ybc85PZmImVg1iNVTmXiQipEx/5F6Ga+IaozQNdc5YNEdS7r34v
9CWTS/fU33RoImLq/tB3/rC1zSEW0vWs8F0tKvvMWtc8Ig+vpNMIWUgBzh1xynaW
XfbzexlQfVaLmMUiVMSRBlHKzQ72pFCbZap2Fw8wwlZrNl+8vp5hpDciJEChcptu
HFLWuwU9olDk+tEm7ibW7sHrfp+R0uhzrUhh7HXhmoERZrwjr6uIt2D+X9NfptDd
zeNvxFkFOkMj9+Awy+j/JOU56FUTrX8zXQtJ2skbsdMwUEDUFjiB8s/ZnBqM5vsq
eauS9PaU9rzk2UHrr5scI3SLNz4OugAyiDXbAY5mGmIGSylB2FT0VBtyR8PdjssW
3MvvF+q7O3ABeelpL7TaA6cfkFkKwsGe53VYQf3ZfnFCuYMzdnCYkDKeY3F6O2p6
prHZToAFyCFpDZuQQEW1Uhgiju3FarwdvKkgOHS8RTDwBD/gbdrc/MOZHqJezZ0F
Lpg/RwW7kgfO160b7aFFmi08tnR/8+ErrK22vjejG8l6LkfvVuByFl2EiDru9irH
0K0q09jw4EwzwnZiaVJKqi4OY3bG2yR7V3bk8+NHHMe8IBR/ZjqD6gqSQ7ILhLSB
LmoLEnY1WQSpzHIg7YNyk0uPJlTQIQD7b+W/lSUhyHuQWKfyiCEaf7Iy61qeLXfK
8KBr+R0KUZ3dLdSblYLR6mo6GM/ngcY8XpBi7qQcQkTXiuIwQ8EJSY9xA7HWurmq
b9S0qO/HXxPB7WfKXhVrnirgfRDw8k0dNvFP2rznxiEg1gwwIwuJiue89KtPJZWt
UuqhK7bRs54xuIMMyPe6ceIH9ErSN0HQqFbuwzGzMIHtOZ82+xGrZRY3YYIa1Qll
ixveQHuPDWUAKg3a4/AZLRIbbHCq5qJmclhzlj7DAeFiTO09Q9eMW5edFWy5qWgf
73u+J9xk8QgMhuPwVP0qBtd/HD9nWTkvqHE7dk9UMByyANLmLYh74qzRhCQITOYt
+XXYLS5vNQIGSgMSvZeMhtwMPqRloucYijmVhup4Qrg4cfoF3cl0/nAI7RmL73FH
CWy1aV31Dq6qz0GnmiaLg1IkZX9kl8tqi8tcIZQARy2ZT0yLro/+W0b/KlM3MB0P
berZhiFqJDge3qukzgi1CL0AwH3KY12oSvG7JFVM/TuZHifUmLRTlC5rQJFV1Htt
kDk9gwv3km8Xx8cNbpzMYIByb566nFoQ1NXC3EbbmlM5Jpa3smFIfrbN2HQJaZfq
wDlkhiuiUP0lSAkD10SCUaUW2LhdW0LpGvnb2KetSQB2bUlhSgI2BLMDPM6aDP2R
LdXK8jfePNg7oGIbFauDGWtoZrcWanhMAkvBHptqQ43oNEm2WQ8B/Rl4iXTF+fxP
GUikvEt0FtpKNWxd10i51WmtKhzE8yWDM1uWYW8ok//S6m5TId4/q4qt8mgar+Fm
GI7hkW1rOAEUmReNlyms2jf4kLTz2LF5zqJdmGYqXbEwf2kShJPC+qiN8ttPijmG
J+YuR4IAbB//OWezgOOOm31UKdNWWzWe2TSOY6P7IQA2c6Z+Mirj14gpOqp/+Z1r
XIKCLc4cJnbm9IPHKfWG1CvX4UoHKxfupr7n7sVT4EpARik35YO0bTkNQBtSD+wQ
1k3z5fO2TtzN+19/QRpjfFICblHufXUExs+FIxRaPvGdgklIiIcUN+vXHbT4aPBy
tOEr0B3b72ZGjuj0ybzEIMj0KRSmq14JluuvCJ/GMmUoHGdaY/PSY5uB/nmdTIJB
xOrD8fHZfQEQ4WFiH+tBvPIwcstfmLwT6EEF/oxvI3eXu4uoySrzd9ydUgmwC6Sh
88n6ZnvCiLRoz8h4EPkwi9xItClD4Z66swiTKsxfAkls0+KN4HGVUDUyaVjExwFO
q4pxwHgzLJKSXMW5mLDJT4AEWNPs1yWGtN0BouwPwhgGlGnokIPkwPwR4rUMMaTs
FglK6DyKrRxrcQfqPphUCewHVSthqCFIQjlUkzSfQaTW5XqnTW/j7BbZOFXSytRc
GF2TmCyAc0fgDqLVecoVVJ7LA+s3TEWLGoI9ocnbTBYtE66++eODM+nPVaGfFUUb
7qXnbgrUGI+9rbDlXVElbP39FAU9yN3OPc/ALNu51nMz+bqMan4LpLEeACIKrdea
5deJSQcgv3olBozhF5TRjko54idWibju8nj7AKpd9KvedVSe7UqjoCnOQ/ADUJdR
FAH6++63z+dRAlsjV4QkuQ2qWGJ0RE63+UjF+WmlgP3+mWwlHOZu4m1/nnf8Qrbp
W8syx/Omc9FaCKWmUiWZDGo5Q14ZKvYIB6W2LypcIpXx5NAJBi3NnOiHE5WhwCjX
G06bpMV6d1OwIFYNJEi5Sd80ZLexaEQf0wAVRkWhrpWuP24KN07kUCesmeAY2sGj
GqnRkp8qXLnxUZucPI08wrKXsNkjqZ3W9RlmGqIeMWCdk9q6Tz9AmWvY0AEfNJtw
/4SwUKSLiJMMTsFd+m0oWLoPitUHw4z6AZB3pvN8blcsRxLW/VzITlrKcpC8eo4g
mq4QkqMTVH7gj9GyJLX4GlHKbt11w/HPcIsU+0lajmDC+OzLLxR7R+RjPXyHpD1y
GsjH6N/JmB6uqMrM5znCBHW+PMBi25E8urNBFaCbYNsK+0yI4z+mdV2lhLnUpYdd
ZVKX9drlH4Q5XWYUc8To3AAhtIZm20w5lbCASoks1zrwHq63Zm/10PoCCuLKmUpk
GQAQnkwjhs83sVVyVp50sWQooj0Mz1u6m8IFQghWS/Drgu5rWt1j3vhOm6zob+sY
p6BjAhIiieEOJzo3IEZTnLuIPo310/3mEsccakODPoIdJJ9ZXiu5jXrfqQ4sxgmy
o//d2QTiDpSD4exuR0vgXalzQT/prUvqqMKOq+SnzVxxHuouo+fQzCw7Eiky77t1
Iv2PGptl4ReT7DwlWMhGgsbg1BCiBsXiWlXPh/sg0Yj3DahJqXZKuzb7zWVw/G3W
bZRpK1cr1oqfm+b9EaE9IdAd7Ow4+6OiIg0pjPrhAQBtx/aCOVvLRLxBpWFPSfAz
BxnoKa9eEEQzhDxfKlQWS7mxsQVGmhxKXzgDAZRlIrydRJ6TU+fP2QTW3Rl4hT+S
PKtVeef8MUyMea7j7SW70EMtHzzzRwbMFJMjrQV/Ohdncf1Vd2xMGsfnRexaCiro
2euOBtRvRVkMjaC6nStDHjnAI5mF+WcQ4nbZWKkK+N1mzY9chzKUiFbH86OFWc0j
eWmyT2nXj/RBZF92tQw0fgHlgxkAXvQZsR2YDEg9mmGCqx2bLZlGNybBPNyoyzhK
HkX5TdgPkd8dkEu2uhiQfMPvwIvNyrxeDiSlKg8bnVeSxLVD0mOgLhDeyG9gQ6mM
ByhoXpa5hntl+JM0R3hRQVRnwuA8XEhWPEoVYpsUBQKv149ycQEp2xsYujDNxY/5
Jt1gq9NxSyfB792O6U8WfGomW/prouJA317TPgoI5qV85gmzcbcUcGbLj1hq0Ooe
rL6Wjrr5SzxmIp6Dy5MfKxK4XrVnImGxKAAv+h2fncYdvdDxaGOF5lKo4eBWdB+n
jJz5PU2rNunYUgOD9hhqqneT0vWlVv4SRGLy5gGrjytce+nlCWBR+zh+7O/RH1gT
khaniFcFX+6WEvcYldP7Q+TRRj1ewECmomC0bew/SJL2RFtof/jH0G24068E8iiT
X47Iwn+dU7ig72nX8Y3SOZbIl1oler7/LWlKTdYU++pa4ut4ppR1zK9AbWbHbrdf
WbxLIObOwrh9uJ4e4GiyUUZ7RgidnRgXPjBHjfnIRq7yqDb0Rz7MxuDL+2xQ9zYo
03NpXRJG6fUfH7pJZ9uuci7vBwswziBkMu3u8Iy4dIbKgv6ZeY5J93Rz7ZSHoIYv
mb9e+f0GFSAPMZ1amGmsRZUhH9joH185UZfujbtxV2fxF1vZXBobbFJgBfxAJO1t
/ADeOEr8qJeBBfW6nmNVnBDHkUyK25HmLd0WeRAldlxAbkdIvOuqYIoHlQguuxh/
dipUFlGdzf7JMcv5jjCx8rwxup2157y5T6sF3XpP2ZPCj0mTBltzkST/OyYgf/K/
JU0/Gz3dzH0zHa4svnB3RQxuEaoA5CocTfXXgV5noghjd3H8bLf646e7ZxvwhIGc
JNP801q41L8eUKGtxuLrfxDnxl6CZzyWiiU4j0d7sQg6Bcfr+WeXml91+JM2HQ2p
S6aaSDy/b/azJdeAmYRguDlYgUrZhUEPVOLi1une1YRRqSITpn0Mk51+Eq77isaL
xY0PBwf+5sVJ/SwTXCEIVZXRPKtqql73h8v4HPXuOMfV0eBiUpIBMf0HxtATXZwr
XTr6ezGYvlOPoWEuOgPKb2WyCP7kNsfUPDp5tJV2IuCpWgJ4ikD10nqnnZ/LJhQE
jXU8rE9kk4TNUTONI/73BNPvT/XZf8RvgzasHEeToDnll8cH7sPjboJXfjtyHMJP
E5nFDccieMmVFNCsz2NsP079GpoVxMvB4s8uqon2TdvQV4s/qFrDQbvpJs0rk7YT
HBrzf3JBumoBIgyFZBOekp2UrdJDC/ox/Og0IeSV5peoLa8Rzn2segGzElQWMdl8
1j72BzFERqRsDlgzhxlMBIq8IfNVMbOVC02TZS1jBHUBnwSiOSFEKfYxBOSuPIks
qwUaKpMgwXwZMEUxC9mW031MkdWAa1hcrRWr/xkGzSvoCQzsIP+uMY+EI65RB7ZN
3oxpcdXrC2uBmJ6DgQBEau2yI8KuHl24yNi1XmLKtVcIizVHkDonCQ5dpGdj4CzP
WDsiyLUgCrBKkXdCSIQS4QIsNjXBq0khem74UkBYM512P5m8p7j2nZ9XcgL7FEPP
vYlNnuj1Mw4FzUwqG18jZYX35mJwh2nW3dUP/GpJFxB5jl3XcMs2+fRVTRC/kqbu
Xx9/QZ6tHPqJoB2j+l3O0iptFDEpnmrfBFQYf+T5DX4+jcjeGtSdTr9rAaGGxSrp
qXFzbfahibCuHK31W4AyFBdjNeDLQ5Ghi12ehPnURue/qMn9k2tUCairFcXF8lrl
v/On1Pn+MbQERdEdflVpRNms+AN6RkTQ2EPyBjAS2VI0BzkPn+HJJhnIYQQKYAoV
0Ej9F+Jem0e0UBtaQAnojny+obSHkf8IZy/N+mKSK9vl5u7ZupaQd1CwDBHYlGXb
WsUGzStzSy3nnTS4mOoZHaJ0qc/BuSfmt1XMNXRZm21r+Z7eyPzAf7NCTp3qo8WH
EyzvDKIauDwv7MrNnyJbBgtapc+lzfJgTHSvzO0A9pzAsSR9mENCHKmWE3AdzbpB
+8ec0DRf6Rmd6gzgcwUC7yylOmp5ZNefNKsX/vynqWVOidYzLw0VG+XGEBfH4RPx
4egmpRociVL9tOnOMmr8//gh9iEZEmySPIBJaLWZzT7D0kjGWt4d0mzhQjjtvSKm
CbLzsU8xNpbWIbXMZuCEE2ES4O1vhobVvJzWBg6l6CSg8wDwQbrHPJsp/+udySX8
oruWmxuGUuLHOrhe/JDLn0gqfLuUFuWEUpr1sitBtERuo+YvT+YP3Di6/ZoI1Msb
fpMzaQ0OBn8fWD0NCMAJstXiE5fkA0biBaoH8v7cIYyl4Fa9R1Vr31l5mSNgUWPR
6POmXpum1ISdZJFpjBrrYNgt/EVGYfDT9YlV3uYHLIaba+eVFriCkHbSqedtO1gB
TwPymbMfr63AkgRAtnDotdEg4fNMtIC+Lh7EdKYysTVNOXgO3g8QgbPflqYonn14
B66jb5b2PGCCD+ALhnA4SiymPgBX7qJXuaZEsc9acu7ESoDxlKD/CB1YF7Mzy7Ep
FCkctm7Ntoxx9zvFbwBRVCoZcAjapjh3pDmFEzOC5Hp0cIonYNcE7Vp0iq+5kkSG
tN9BndslccaXIET7t7gMjMtmSyNQsL5nZFtm17QJbdYKSXOV3El+yWGPhtLEgkSK
I3qiS0nf8x11jWiPex+a4mZB0CyXzKuAalgdIaMTY+equrnzNEe+udfaXYjSV0i5
7co4zdPIrx0ssQgolS14K2HkOF4XHkpxbV3+tUT4Je5z8exbMrXmqQVeX67mUfRU
S4vks4+lJ756cVm5Ll84V+Dr3h5Nh55InqpejyCTgT3LBSOd9oi6sEy2CO3ub6oA
u6uiZyjDXEgu/Y3Frbmd9mb1qdy5NUi7CaJDAEfBFsoznc2mDlEP4WCoI7Mre//S
+j32M4MlTLIAgpZifrFhGFFLOwhbGpokV9FcI4ysf80NjB8qpC3pmxfjva1lGsfY
sC5yG5s4Pa18uYltuQhaUGXGd10Kg9YKySF82AulTAQfiSWqZntF9s83Ty4jHRYQ
9dYD/Td91vcoq4GtGfw16by/XiHQzg+TKToyhkUmFr/sASiw9jubPs9Ra+P4JD8G
2U432+/GbwRKeENpkNMl6Q1uSk45413tR9VK0in6ixz9Av1amKMGfxoC7utfWwdo
gnGfeoM1JRW8fEEZ8PP4RuWn78ovGQ1Yfb2pNO9dn9EvIwqXZo+E6wRIFoEZPy7g
3PDp6OUWqwQ9wFWPJ5wOph3NhGIBZZ4gamb0+OxYdDjMO9Fwdnt63TnMrUZ/+ieQ
Yvdpg60DiOQazUBFr7hAfazwqSwbutu0U9cFBIfGBTIp4dT6bSRa6haycNMYcsfA
bWS1fpm+Z5l2FAlJQx/7HMCPZXoz8kyaCSP0FTbXRt6a56lEa2n4ZrbvY03Pg/fU
qsWTK53k69mPIMfSw1VnItR7bIRSDekTs5Aa+KuUR6/E4NCes7TvvLWAchwrjhFM
keM+TF0Rnx64sBqttOdkqSISWzPinfN7EMufacewEkUusoBsJmRX/iPzLrnYncd7
lMhtY7kX+2rIrJMFalI7C9F/FLIMIiN8pdbWGnILSqiutdocu1ycsHvH50UyDVtG
wgYzZ71mKf3TKhThae2tirrLojNJVbduEuTEe3Ha+K35BqHlobX1TbNWvZ1AuCNO
jt2O7mm0nQe6Xltnrmz7EnQInrIuEo85xVhM5MRGpZ13SKnfBBE+XkL2P6ZWxBkB
Cp1OTX55aSOOHKHQuCD12Azrbr8r8rKvElae82lkIbFST42GoxnURGDvK4Bt1DrQ
ymYgxv9KQm71ZESk53WsrDoXcWKV9wkpx78LEXR5p7i1e6i9ynySt6nfNnBQTixl
U9lMqqP9PcfGQu6I605E9DwKrJxd3k+qzJ8XGhj2bvPnoaHiDNjKo7YwlISWnheA
rG93dT5OAVcSTFjt9BCPUJ7t/XG5DAqZPYHHVk7Cwu/QIpgD3XN8oNv0x6YunFhC
+1ofo2/+qV8nSseQTGQNHR210aklMXOrh8Qwzop1r/olt+9MwilATZ5iWDj/NMpN
ndt1I3KNqisPHyXwAMU93xV302hXONmb8PP52gJVyXLfbltR626rQQyXD+H8Q/XU
I3W/wzmGAyJkXa4hY9kONCpBtBCH7RbJFtORocD9R3OhPYZncdI7pRpHkKD1Q9Cy
/FVQkRz+qtLgjmv7T4zXqig0Owu7r3ngE6f/zFzpZHib0igiEsr7KvyEpeZ0No3e
W6dvSVAJcHTkBnuwETKAAWoF+hk+GDFYhp7kBmYs2cx9jWpobhQ6dFiCPlLBaMMt
438RERj0pSMeK5StL5ag9Hlvo5DvHQmC2UhMZc3uu2NGxPAfIz946+bYdvaSTTMZ
+UoTd2pVXolfs3fjMRc4r1al1OGQPdDeBN+6FeJkPMxHd9bDpZqNA3md8KdPplpy
GNggSRBGqCCCZaeGt2iP+jAez/fxbPTTSf8JIo1WXUEHbD1gDV5P/eILD9WsVmaa
RGNSirq7AGKFsNiFjX0LX2WvOCZC18V5ol0iyif6dKw2ZHqRBaP9FrTQrwYkyo+G
llaSMvOnycNEr0WDsN4EDJQxkqtfz9xO9SL/pn7E0LX7Ds2y3mN5iuCOaSc0ygnQ
DOPv5CTXV8o68U+q2ZUMaG9JKXP2+I+1O8irVYkvgKGCEj6s9FFb6fsctE8Mh5Nh
QwBIK7OXPWLhJ0PLqUu9KcGskRp1YE2/L62FkNemmnmlbo4nYw/9LZtmyPeOyBq9
IVlVbIqRpBgpYBCaotb7w0I7A+0OEckbBo6Zrwl4sCoRSoIKM4ywhi1iaka1AodC
S+IYTS++aht6+c69vnU4qlxO8BSVLSvBtiXci+anEXyh/MWiOX/2Qck2eqM0a9LG
tnXwjX4uQ1Y6A+PVd020FfQ81CQlheOEN6236NZWn4W2tmJ10BNe7iiNzrW9v98I
NMjwYWQzOJwPCjPFy3iedhOTvJsmU5Bsunw2+EFMSJFCJLF3txYJqJtgdkn/jL9i
TQvnoAq36HooLE+AZgT4D2oB7zJU6Dhxv3TtIQNEianaw3ayI38OnUWOaC+5rsjb
IOFnYUIUMcBaqfjFTA+BrF8nmqEyIssFUbVC3nQ/sNE3k+S74LYXuoh/uVrLxoXY
MicIQSycQqQFgOaFIxi1y2dlbC7Er6qZq2giTPj8hNM9QT4Xy3ZDxMAT+L624ToU
HlxHprsbFotvkUPEECa9KPU8CTa830lNSC7qWdWJFnrciL46kY3o/JhwLMZ5B7hL
eMdYZcv5Iwh1gOlrTVQPqlUkNCBJmF4OgPHYJUPz/nRfpAxknoBDPhO7RPdAZo9q
a39oP3CQFJpxYzDXgeMwzegGzQ2z1wmVnQ0S2cnXcGiHj1Uln0Mzv1luo6o4dJkV
JS/Fq0xeoBjXEj+6Xxds03+Diw07c40bOmTte2MQJy1YrIOtj1LLa6HdGyzNS+Bx
8xCpEcOIfoxOl+q04WzPe2JviQ3eBncocn3DLizuvuyWvyZFfo+MSTJ8DgIKdull
1qCTOuYLLlzC64crpU+twpMiz/DfaUnKf7nSvDglYEjCNFEB1G15Y/NGO8fsv4bv
wk52/Tgmqw0pWrBvb3GOgemi6K3uTqgzz8a+qAu/kgLanKeetPEXzTk9QZMRFmg7
OcNwHPXhiMERu5URBBE4o5VfOm3uAfiC10BwebamE/ikyG59F+TZjdzHxQm+PIWn
sm453ufvX+O3ZBKHZ5dKzbTn/P86gLbctDV7JnPjCWn2MNLMx+M+sLZxgu41X00N
EM1S7oAFjrON0uQVMBKbNlYp4fYke3tixcTjeVoWZD7zhA1ABGHEEhRGmTI8HR2f
`protect END_PROTECTED
