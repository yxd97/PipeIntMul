`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qbZ31ffbgOb3zZcQy4rLY8neSF/8MGH9mPBziTZUwdPN44S/yngW+0DhaovzDEx
PAHg1YPtmSV55omiDRk0950wwSVcV+RyGP4/dgBcSSOPb4LE7SDQvbQG5TGPMQou
JY0wtMmyPVZrJZPWwtOz/fodNREZoVZr+Hak0XOaZy+KPTruAjY8Sbdi/8/DsNfW
lLdilkoJPC7WJ4eCALAkafvWPsTQuls0ump6KnA1pb+nrIBXGgQVSfdwnWfvmPZ1
7RvJqg4NMUfUSQfuSZrGIXhY4EbIyjrTaOmTj/jd5pU6qVbFD/TCs+P4hVRDd4pG
VkcIm+nnFLfnBcOwhUWMYcBKpMK38PaUeNeEPIBD2OuuoMPKvCRn3ujgZToKlyMo
CF7H8xHF8NJK00mhGTuXi858/zVTLuQNLbWDsAsngCoPsj7X36q3c/zO99V/i5yR
kTcXhwgosqAstk0J5KTh8XBUzIDGI/xIEWQcwbFLqhaszBLd56NTJEhWfgBunxGp
vdubw7AG6TbitpzV5lTiGwDdzINupVV8u4q8NEizcG0EWWyIGnOFI7jkA7VPna+0
RDJ6cjJjESZZ6bT9A0+BYO88Pm4KO3YNv5x58iFaCKX78K1Go7an5+uoycvABaUp
MvbX1yz6jTtXJA92aoG3pZfcET9amkMSeNasryT1AKlFDz9c54HQBjeInbzTOpop
wyrUjpKVqESuJKCHvDf74Q==
`protect END_PROTECTED
