`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yS7QZWcUmOXEJcEShNnx2J4d+G74ZoqfFb09rkFTJ70IDH3VdG/uj9LWtFN5pKDw
/CBrLg2YGOdTaMZvuKV7bvtu0zCjfk48cmKE19BUMEd3r8B5OwzcI8BWLW4Xnax4
mzihZ804KM2pbTnle+Iw+IvxpxtLa7hFE/jWVtZwiXBbG6cX2G0IKBB5lmKNj96/
omLsq731hBjMGKU2q9FLNQlrPsxXsQdGZcnw1HEAVMNLKYh0JP06tTKB2jBNo0Tu
SePe1TemXn2qjZm0QVo5tlK62dDKHess2j9RXZ3mIz8lesFRiGbmwZtjv2+GvqKd
mE+X/VuuQvjQSCJ7nMNgM7HjDJz6ddSmHwmD9eFLYUs19fMf8LwlhFIEcv1h5Dg9
1WUPlLCz9fAPpAIvFz62QQIBYrAum0MwzKxc24a2CMZe8khZUzauCDrhkz7uJYJb
tEoaMGiEgLkZ1sJ8lvX4HCvEvr+/jyYFLv3aGfYUZv8q2gF2EbEDP8FXp9UKfd8l
gdysyLwE4FMcgel0yAXqClk/cR3OnmvqGYlZ/WoO0SyCihFlOSp1XT9UJGwn01sw
S2XjPvj+ZfjWvfUQHoQCyUnYl1Z/kPkrM002Kcpxjrqpl3rj4UvLtpNTQMxIZyhm
HcW+0M6twsJ8gzqE4LM5uLQQ+rXXbgH6nzCoFzEF8iUTJ+tCqbMdTz1ILlAEmTPQ
327gtCubXhYMxmUPEQkYNsAd7hnz63drHDDa/mstuGRJOkzOFdxLHO2mxg/W+TNS
4PU0vR+1HaQDr9gg4B8oenxGOuSACLjvDrdLANSD5p/zeZRUTXqiLc1lAdBKfsHI
UQO0R3hS2lJSP1ivFiYTEUsgTig95ehNzEWLzeG5QIPqTIgB0W/36o3gxrrI6nbP
X4uMT6yM0aX8l8PtkmLUF14gyS1aPW2hC5CgrLNUMBVDDMO609Dul3aZLqj+mWQZ
d+2Eo5Kra/plA/h/Yn2TCaYRD3df+ygp3SQ6G8UdNhx1IxPyaI35Qi6SUAfTSpf5
muiqRlh2sCrXjHsA5xdFRWmvhtrCeF9QphXTJXcJhjreoQiKHITDrRb7ivwjMBfU
OM25i2gptUXGlyiJRfkXJiWYKZsMEg8MFjxCpaVeiocTap6nQbCDVOud4let3n3+
8jm31RRLYUC/nylTmbGZCPnCBS6xDK7bgLfvFjvFNRN7isJggU74xN5t1vDLAR61
K1U7qEhI89hD+PstKvc/LqX4NljFP3COFwPv8a7q4WfhB/j31wnAoUNSeNcGULxG
tN5JeqXm+5sDKQ5TkvTAZrGCYNSpdm2oc/O+KokLspeFCKwmHS1LJnqcXLlvndHN
nfHA0LRRszzgHdbWTFtohnPtqSkGwMxsfsvbTV8JIX4+M+Ue6DvctxFN4WOJe6Zj
AYA83PAF4DAjcjhRl0JmMcR6eqt3b7UQxFtV95hnxajbjVQCjbJZBqjiyZTlnNNJ
PO0d0VEHNJCXrxcrwaeYB6JQzFPpcS0Onc63FplIqnDYeLjP84aOK4yZNp2FpmOx
`protect END_PROTECTED
