`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s19nvw1NIUqkGYPZmuKm3QFJtVEwC3HonIVhEPFj1dZHxYlb+rzqLLZ7wchNg+AT
1IYRRfvCc0MEo7UtnWjy7hBwUZHIE4EoQTFMRLdpjvBL5WxRM0EkwYiPMH4LwvY6
Zgea50Acmxv3sw7sFGQFK0PWLHwZuvVAd+D5pRMURZddoi3VL3XUVehj4cxdEcjU
t7sH75mqSAFp2kA9H9wuivba3fmN84YGrqhNuaL20RU3T7gl5k+FefvtcnIy6XsV
6yEESJTqGvXETombReasb4O8sQPmrOB/B6T415b5iVxpynMzKzy/Hxc602313RPG
9fuK6XLoYZlDpePN2fxfle/KSO/X9hgy2oAoMlYWqH5tmw+NQxtWX3b1rY4virh/
HwvF3E8wDYi7Pvod4WeSZ7LjAF5031DTqul2cfo/BgcyephZ5QZ0g7TM66VWltaA
leZzUgf8oy3fEDKLpxxIXCtx81jgR5fYJJwlsmmei36pers7ySidbu3MZPDauPOJ
CTIk0yUQBZWikCNZHSnxjQ==
`protect END_PROTECTED
