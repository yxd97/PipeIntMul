`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehFwaupvcRJDWXYf0g/Sf/+yF0PLikHfPEhnX2jVUWL+BkwPU0Y8Biev8jnDNZro
mAfPJvuapMRZw9bSZdKYvlFas9U2GtfyOLKKhR3LuGyhLxmGZ+f90HMKTJeloyBc
35aQpjpTIY9hoyVwXZavARNpwhA7CbsBZFkSUPVnaDCyJ8K2vBE2rm/CF9abrC2Q
lH0+nEkgT5UxutiFRCxjA5hlgUUm+nAEUg4uqjtHq8NGE2H3WBGWWEBvgq085tlc
WvaTbKJebGmbKGztyOxp9PCnpp71Z4YzuJt/tF3BOl3qXWTH6iVWNF7M7LugiL9k
gCimLQhvmh2a8cmkJHTIlwYnb0t+mOVwoOzp90wbWbk6TcZeIkcgPzPDr0tLY7rF
+V8k1/B6nrPmAo86EryYQxrX5Ww7/3kdmhrD3VKP87VFWTYB1lWWooLrY7GCK9FB
UbrggkeYseF7SBdWmRQr7RZzs9wz0n2CPBTXNIhTYC6vEyF2+CwowH5aFTlfqy1u
z/gv9BHnog2exLAWix8WycauO0AmZwRPOfz/ztyrM4x2UQi5xSedEfZ2bn/lAKDN
QdY2huB9koeymCRg1ZR4GzpSX8KBbKKiFSpx4hdYuWDwWn98ymcQJHwyBnPNJjhN
e+5UsCmZYewpaW4uPbXuLWOU7/j8V1P5fuS1ZybBXvivb3mZ/nIN40DV+TmSlawo
Ct0FLjXdcvRWyEvvzLosSm8ICjgDGHfrvG9COKicfdLe5sH8j42YJKd8arzgiZB6
w+oD9BapqEA2Di83TqvNp9ugPmj9Wo+xqf6oncnGauEyL7zQ0wwXBY3Ss95f1uAA
Mzcg9rCkkFoLNOpWY1Z1HldFevAYNudGLfLk5RW3jFXEWC41DcUORLQHweztKeNp
k77OJxNR6eXwWaDTt9YUmB6EzEZV0k2uPY9gqDJcqk/iDnHRHc+AK/rCovVaVdkc
QK1NDLRrgJ8S4Xpgg+SdAkDnLWSci3yzYd6xdnN0/5QbediFX7LrRLGYMhNpbK+W
/tPkinU72bZp+vLzAviGt7wULwX6v8dWZqu8K4lsiqbISIQ+oVvIeLVDHJ5cdgzu
0tu+doitQ5fL6axpQUojwVD77Dho445OL+2O1JSDsDWM1oL3ysVOXZkNRq5HTTM8
7a9t0Q18C1DzYXL8gHjsKSkAOc9wDEBOai9N7o9NdU/YhwysU3lBHfFyDDQb8mbO
LyIlv5hBzarwf2TKGZXI75PNU4Qd7ry9+oHoVI9F/7fST3ZQdFQuapZkowtL8MKq
GAa+MII4OFtRTqvJPHJxDw6cPFj1aN59SBan8A6UuP14P+tDmRJbn6erKOKmwQQb
1hdrPeDT410wf/yslz/Kcg==
`protect END_PROTECTED
