`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wo7+YogYPgZ2ZctUjaOKxu0iaKYwAmynLFVquPX9AEGPe5vAUYx++IYtrfiVq3ZN
NDKJ86BDSug9dyT0hMFcXvHJwpxC3Jw5oDekx1EeGZWbg5wXpWJnva+x5rlemX/m
BiMK6oCuhhtfsYT/L3gYKFpv33+FxhnYM6/LlonUudf8VsJVxpNNRzzcKeTbDNyS
0aqird3CX8Aoeo10KSG4ZauuH0FFZMKyPN+PXRJwdAPtCQLWCGoE9OmKnwkxe6Cq
P+GU1mDIB2PhMHM5BwAO5QQJgQmJWFVxB8ehTGtj3Yo=
`protect END_PROTECTED
