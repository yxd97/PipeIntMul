`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ipmoHFlJc5tEp6fWmmYM9qjrKiA1oVpl9ImsogrvI/TSiXOls+r/vZBAiobrDIDU
eR9Mlw5+jK5G0nv3iGB7MpvSXkSu9C/E6JuKYAA+VTQVl6uXzRw6e0CthL1msUOY
RpRCXzB5l0TUoULpIdgw0FMNp4eTceUyQoUj9DOJZPrvTp2dDD95IIAH+EVQOuqn
kw7YhhsmH3H0ltLnBm0EgozU4FCPWpjfELZZUU6qHEtBZNza4UI+j/U3pvjggmDq
5VNHnBoIAtfaaK6MX8/Y+Xh1PWXeaqNprNF8Ndt5H0wbHitlaJ6ZAJBFJSh0EyhH
bo33FyMOjcEZB65w5QCCl/rZWPQHvab922WOrUO6oFo98PPYHZrqrKXhjV3IBMDR
J1lx3ttF/jk4s005J06Xr3B6Gk/yXt+3Bi7Ul6Za4Yw=
`protect END_PROTECTED
