`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PmGj9/cSaRH0zrPqGKbXsnKMLx+5wQHu0s967OAeCwPNquolRg4QmddajYis9+PI
4l+eFOUxoilB2QjOwDw4soWjVAW3UhqEjVZ0QbKOZzvkPUJOPMM6joC2Td2MjOrr
/ipHbLb862ivMzW73ZrGXuAHu5xkcrXuttwyNeeZ9n6e+rGM5eYBNs/8wzV1+Vs3
oaQC97LxiH+GNohZjlUXp+8w+RRM9taO7hsAOgDXUzAoGh9m0qUSecoUZlxrtiW/
2OA+7UtDrYjeBXW6Z1Rj6Qs4F3t6dJXl5i/4+1R0McF013bYsPNCOKVq+G83seNv
YsmmerkO9Hgw3dltssJyLjRKy6tDluUuVH+HzF8p5ecWd/XhBorCd45ozhi0yCDI
8MXGe7ilukDvzhZIZuG3a5r/BvDEhhV5gof57Tl5BiM6UoKWLzaarT5PfloCX8/X
uzVdH1d1KF6RuVN6uPZmpiieXi5Rg6kgoWR4VDo0sU+T2f0EiOpll3za6pcsONKi
`protect END_PROTECTED
