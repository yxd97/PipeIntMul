`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+sFCBZGQnryyvqLIQo7e/G6P77UpBIazcxAxYTbk79KfT7u4++N9S9WjPAiUOgZX
+G98R3DcEv7KMiALwPdX1yFrvVfYyPmtBXabGNjCvqn9h34zFzIp2I7Qqt+lld9N
jhYQBtwMry4kNt/prlyVG02AFnD4ki28D8MOYmyQP3EBeSQ7I0wIlwAqXJA/KXgl
zOydwFMooA2JNoA6oqoHQxUMmPIW6U6XGtxvA9raQOQq4un8qWAC7eSK6bTtlQrQ
nw/9vIiKgQ/CQzUWEGrO5p5ol5r8Ho6zIbj6Hcl6hxVDuj0WNWGNwx36CUB9QXSj
TJ5sUE24d6b2m+nFIlBTXtkxZUQ1GF4eLi9fHkv7K30o5vj1eTbivdZ9GPuhRqns
uPWRpg6B9BcRH9tA+/EWmG0nBUzGOXvqHumbZTysennpKl0SaesnN9OFAsl130AK
2L8R6r7YUtjiDkLKajbLJueG0ZeMahfXShArpByTMRmGhdgCGkBPYduULYXI/7RP
0iRqMCf1NTb/Is0o+fx4uSC8q1NSDwFA6ze0QeALOe/6gJA4kc4C/I9BZvNDcJb8
`protect END_PROTECTED
