`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXmhEXLpphGYyjqTRaJN6UM3NsqzE5ZXon7Ux/ODCmCdDAKPBYI3plRdBklsP0X9
pBzC/dTwOQWPNtQ+D3XYVbwId8oj1hx/WWdUqoG2w3O5SqanL/fyYYlNtCVMsOMN
g03s4cHY7JtWFRclj0w8CUlhJfF8MGeROHXPTfNCvjJOFzPzbyFZAPry8BFHIRnk
lVkn46/A2cHRxeLB5jkx6HpcHs3+X/F8VHP8KqdhCxizM73cLFIcaqB/CrISypjV
KGrmoHqswYEMcno1WSHiavxIzuIKhXTYrGZYppyVHNoUPxWHwXvpShaKCegIeU/6
TROP1ioTQ6j9QW/Hh6zyQ6QHF4bpAzM0G1M7ar33c04TperJQOhOO2h3slUSQcWk
hpaDpCNB3cGBB9v3bpDz/oV9qPjOhm7FJMJIDcFgjnR5B5gQc1xM0HY326RD5hpc
`protect END_PROTECTED
