`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZJ9sl1yI1oOOHTyEjc1katQ6jMMxbzMa0CPTjEOc31wyTjlt/49763DJWRpN54Q
QFMniwOMnWK0A5tWwLh7zA+UmQx3Ms+Cxp0ywECAntnmYQw0D5tjbLcwxYhf0tfg
3A1Bi9QW0bSn79TicE29Dtvbu8h0c1h1fL/+TQxHlkfrABUXRWX1su6LC4UtNE3V
9Z+IlYpEvPWqSfNAP7EKZ6mNWYN2OBzJ0w7UJHVb4QEt2rc+dVtK/bpuUN7ACaU7
OGCdHal6QSc9dnPSV2fSwMrz3dboCkZO92XJwd3opMcmfdEY4hEFWcRbtwCJGKTI
T7i8sqDK4noIsMkmPW0UpcJ9UQfas0HU0Dv3tJZjssv7dBoRvLcgV5jFt9wWaYuM
ZjsnQ6WeafqJHddOGDtI5eaQIu9fderIGysgblsR6XNT2M88SHvY15Wso6nvxBj3
dc2WhXvovgKOMS+PtAJZpBlvUa3g/5mZSY/jnN+tkJmOxZtwxecr/B3aKUPdgoar
gWzokJnpCXtRw7oInAC/COe13pxox6qTLHR5jBCRDhz8XzSxSpqZjxxZykf9/nv1
xkeqisozmLgkjwJT/FYY9TiESV/xCEokODjEd1gpcN/RuQ8loevkqIbIe14NjFaY
WcvKD82Y7YZHrvtEuPOiqNy18JBy3yIbR4YMLgyxg+/FhcOGysMjAVROOxhiAEAH
yhK5IEG7SgxUi20axphKuBk+P2P3WDMlSq62EcE7KJ9MVkn/jgYkR//NIf5Wprd7
vEuomxV1fajyg45UNZwcCNiiVTXYtf8mwhvq8nzGkJgPfeifXOIPfpmKQ077FIwg
VwrLquEPKDmBpmigRJW49NJycxO+3nFnsbaUSMBLYCW7rjXYz22KZJni8S/PlE4y
fY+5bCfhBuvwHb6qsfDwtri8hEDj1qF14V8/jSSbn+l6xT8E5OVLGLqoZHbSL/50
pqglRmHdIgfWF5+Oue0dcnX49JpyR3xTB1hzqdBWVoqzLr0B4jGjDMic0Y+OkHXA
zx4IRFlCRcOrztvpm4yfEMSL4lRU0zxRsUMuzN2ZpZujOLiSpskr+vSVh6+ffFgk
a+LBzPdtfOXAI+w7+Lr38qRcstx6Fao0XfXJZZRNcOPVs/Ho74nyjnA7zFmOvG6A
HyrpJXhTRisNy/khXg08kyFrxT0HKiOWCZHEqTUU/eeHSuDd55CqluVxfDHHs9qx
5LY2aNov34jQ29bV4hsklK6koGGh401OZMj8oezIn/KylmunvXxZcsdXJZbTkZPX
fPB803ekDR9A/FhhtjU8+pKr23/OiHUTR9XEByN/XHwyqnmuECRvGmJP6Spv/76K
2yvYWOoPkef99uH6RBBQkAqWZSqNLXJqMmlONNaKt5OfLzIagaoQ3avXRq30Stve
bayuiN4yCXC5JGWCF2udg2WgomNTLavmCbRzwtx0MtFrkiFB31TC3ANbOd51y+Zg
xVZ+HopNVLjQNi4xrwDwUlQQrGy2nJfwQ5zF7cq9LCdAyf0YEah42o+cEI4TjnnI
zgDj71OVxfs9AgFxjsC2q1ckB6OvptxMpMdfzCQuw8BYoyrBXGvsMcRSG/AAjnrO
nB72B9cegrtw+sliZah+c9fXo9ETYajXV02adLsDCAHWp4pQPXB5k+Hs5N9FfvW+
dkj1f3eri986nVc5B3l94kQbY6X2r3Tj2bCsNT6pfSu1S6BZn1ojvmdE/9D+D/5b
Okrb8heFHvF1IBV1dKgzQXIr8WyzMQVZRqbkip1g89mXBh+eL1Aa8oE6EQx9Armi
M+o0NHX+CSWuTGorLYcB1ZcEfFD8Z5JzSaU9K03jloOHUKb468ui5HIN6mT5Gy7z
M0K6mk2376UnXpAZNCvcx2Waxyv7oFSfOWmueIBXv9bCLC5LrQKa32woCWH95q0W
+TlOefpEJER1RogTiPDVFApd5qweep2GiTdagM9yHK6AKV68VU9LSt3d8c66bA3U
TGMLK/Hr5AJNKzyhgQR2sqyNLq/12DREAw7/CI+5UwP3S6h5ijWQbe7fq1NCl21m
7I+3BUlN7Lb18frDikXpCtYrDKtOeBc8vaBS6vgnD2pdHSS0SlEBztsTJXMFEKWt
9kQ9zGIG/SSUsWF/RwGukSwbQgTzKt4QEBDzhFCoD0EQ+e5jC0yA5OSSyzQ2jaAK
qi+YpoiAsarGKy99wkFTNiepQkN709FpCY1CxNCWeeC7jhIDtD/EU/9GYmsJBHt2
BzTFM6xYTC2Y/+wz8fpPh9SxQ9NV1b7j5oju4vQVyf83MgqeE0986i4C5nneA8nF
xCfeVfHdAh2piRvg4IUfPgmm57cWF7GXY3C9pAzLgX4hWbnYRrMLagUjv2mz/Qem
Yo86+dVr6ElnqOFEO0fEOp72Iw1bstpgtvv5NofhE/TojC3E/aBMUREOtcvme3/Q
TarPzZWyNIGztnWQWr0SRFF8g0n+aEXYmAKQfhNhlVRCF3nf2X5CKUNUnfe7Cilj
/TgOUgJUqFAcaIgqt4Uc+LH/iycIMy9+rE8zZdO+XKdEDtB5AarEIss1LuOrIRo4
fWi077xJVaOVKB2kXlPyfcgBCOKxmXeqmVBKWbbQrDyyjrxeHSNa1jbHJFqduuQw
McjrPqTK0bcsJKgXZbyF+OeogHIonfXwsLweRHHwfgdJtvPsohGMwGYThkefUDTv
j8PCUQBj/dOT1JHuWx5dQR6KhwU3c2n6HjRctFLuNdAGd26fXUNfiKHHibClfbLt
RrPubwB2bEA2qozvmOaYQMKs2ReMm6y/n0DR1o5Nfw+zcVb+zt9kV4ryTJQb1zcZ
WYCSIvcLRMIIdD89fzc9Nz4oEYRGHA9fe+P6hxL1zbfLWMThQFzKcFdwTtfQzxuZ
WRaWpsRNssYj6RlePSp2haTOTHJ03vkzQUB1eHfB8EqJ5aZRHQudWlFjIbtMajtC
2699z+nWqIq8caqKpv1N/xvfrURw5uzA0jNoPRmoga8xrQKHqBhpUuaLiq3bNFP4
/bETosJwdpAAgVWl1gnnu9QXuLdJpmFskJfX/gAY9V89CYxj/cErQx8DnVQ2ZQLh
Zd6sh2fyT3B5KwjR0GUnj4Y/+4ON64otWoKyOr5KgVMty8nPEKQEYXVF0O6KRuM/
CjqDY4IPG7ZFsUOeY1Kjn8DYE2PORISbfqyDUUhJK5Us/IfbhBDNoJjs4wkYrwHw
pLIgIGIen1qCI7J0d4qOT4qrKPCgyPS7DFApqZMXgxTTpM6C2BLqyB0rMPkuGjXL
HZtrU9ydplK73MnXm+CjaWiADXFLB76RWFznjG1TQeVyqCGLvnpRPRre/P6RERsI
eOYnaHQ0ZsK4+qrCfYlcllHeS0asiYwddjIUBgFxzXmt+0PFPts4okobG1XI2oMK
BtqDA3YsDOqKm7nkHtWjw/4LOu0JNppzXG3zkJKL9iHlJ8W7+fPx/4mS9Y1D9zho
+YBKb8r6rcGTNLyq7PjoYMq1qg+V3Fj1+I6EzQhpvMf8Ir2Y6Cd/TbDC788m6PUG
V78Mlw4p3i7YC1DFcDTIwAro1q7EbnHcMLTMeVY42AxtL/jycSOLllCLlzi9dFx2
MlipxUyjEIepYiI+nKIjaGSSi5TsUlXilJ5Nw5ZnTOth3TqUuCo1qf30Iof+hBlk
kZaK6e9FxYszhklLeVHMlEfDA/371WTrGS1/JkByT/h0VX5ILMYn7hZ1Ms5DZ3k9
XzJ29uA264zEmV8dIyCSMJdMbcbBDmC3dNOklzjixuxJdFAJE4ndKEIi03vCJk4j
LoUszArrzHD6MUkHAecpZRbtnsMYvLrxnr8TAhrDbca4UsuTe9CZohVMPg5lVPLq
rVy8QXOUmVpVi2MyG8Dy1RwL+AgylRElyyiRIBv2Vfk2gWxvjKkV+BI2h/lFYlXZ
eZ4hV/Zgh39KFrAF7UunRmgCDBD+JdNYiTXQ2tSXw7mDrP1MTipolrOADTNS2JgB
SV9We/TITzTtYGX9+Pf/VhF0tyQXTZ1b/qy7ClT3VV3VzO6jHI6L5gIWhULA65OQ
3M3I4fLvTBzn2m0dumO9uENqnS5pmg/+tSUihyXmGOZL/MvbUjPXPL0GTAdLaRhj
A3VkjhpCNya7kipCUW0j1yRI7UaKJDpM3qszW4Yr69j4hC+CuBkOPKxeBJisaFp8
97zT7b8z/RvUvN4NQ1jrRmGpNiJD0S/zuzikiFpqSehbTYsr94Q39LhKkgqrU0tY
dsK59HObnKMg7PaRW57bVmfR3A9RYSxy7QeoiDthTKcB+1F4sFy/OWWEo+l0AXVX
TCp9tnD80O78EtnIlhDQtMGQXE8MQnW+lQ0DYNZp2UJh5hXxrHFii0Im+LdNFMfF
8upiqNQkwnxN+0wNX62QJ3LPMqn8xQaPYy1WdJwev+aGAV2vvnFhbS1gqfykIyBA
1gbwYgS9YfTLrac7G4xffXjl5tFgU/17tjFwSl32bGaJWamVJvqyJ39PCwt8LoFH
LzPvx4eZmy/np3VR/8KYie51O77SQ49bDkOanSExNjoeJvju9sn/EZil21jjCPis
ej5n6jIJyz668ewnbBYppr7R5EW76xe68m4hDB9jpZqyXHiDKxIIddcBrHCmJdHJ
5SBT8I04flpgR8O//Rl+RnzUmDA19fEds33XAVsPZ8SmYFevPq6Ex8k6J8rwOnpZ
XI1S5sp9O3OWwa/87VfyXSwRf+cyoEvIt2U8O094Z6ESeOid9rwoMH0Ps19LuUZV
MJMsrQ7sQR0tqs5U/6vFBv2JYNTMXZ/79sTIRdVkQrHG83m6VvOCT+QJBrJhiCyI
FAVYZd/8hAZXYoPx3sxUL8CeoUA474EwNmpDxh1d6C2ce0pyuvwSjt8iSGaiKRAY
Er3AejXN1E5UnAVmzwxj4ylCC6IXFjh9rb67FZAUZBtCh1Os76MOt8G23NbTcpHG
LTlyymO6Op2fXbqiU5BQRPMT9SKUvSYBIqDd9A1D7S3LgcF1YTF30Me3KIZf5S3P
4G/WZM94zsw0V1aMlVtwdDPMFIRgzTIy1Ag82CqiHNUb1w3dCa3pLffFcYh4MkHQ
t8603IMAgAmeMNjedkqHGaLKE5x4d6Js1wRHmDRsAYJZxAOxbVHatUc2drHugvza
N57NR91l6L2sIwcTjjbh8rXYYF2f8MmGm5+AGDqdEOSkZknMjxrBdAe9xQZxOXRA
Q9gWok+Jf2gjzG9noo0joY7DmmiIvkxj4u/pqrThrCGXjGujyWSDUW35hhHu5rNG
ekyqqr7MY3np2ILJrajwdO78ISLTbM4MPs1AVqoIgbiOtwSywuvVulpvh3/ZRV4c
qr5as1JPFqNqstElWx85MjxOeO9zQHWiW19ibepA3l2/ZG6pN9rwzfTMlAr7NYJp
F068IW5olAfNGMwVoPgCNuFNu4WtlkekDwCYx4c3q4J15qVGIA2FCfeiEcbD0mTe
rnUk2HmGfYCrNN4lmzrLagaMCN6NBBDoNzaci7cj6HOfK7bNn/dhz68k1il8n1aS
lODMkTxUTTtf/RKb6WUwi9DTnL3S0ePuoGhXZQuZq7f6AyTsFpEE4a9UikloH7RB
uxNeVn/fJ1JwkKXyk1w0ElWU32D6icPhJrUa33XWtINR/ckinobiGwub58QoDaWb
wPie9hQ4MTscukqRbb27C3dOs9a+Nta72ECvYPGRpEz79pZ/pKofvsAbIPxU3MBF
I4HnGvVlReoFycQ82gJuxj4vkfHcv2zFujCLX8g3sLX1S2xzFji1GfBRLrE4lRZ3
CqQBchdXtvOUdqGoBSp2lnwRpapAvL6Yl/Zuz4Hj0bKDOfoHbG/pzftWV7UoUzJp
H2gmUZ7X+qgfNQFwPUf1e4SfhZms5KZrAT6iTsw91e9bbv0dWZv1qEuN59yuDHzB
xZg7MfVozkXkMXQ//qZ4LgAVrhP6C/KMzsb+QMmPFVzqzG1uFmz5wzXrajCskoMu
Blk61n9qDpj0P8+qzEMEGxOjUbxd5QZX3KRlOJ56lkC/2cPNuNwJnbYvSzZXtUc3
60kJYu8brmcDb5h1hP8uyoVhKJtlxGagmrt0rfLq67aKWdHXrsUsJ0WnXJZNoAVT
UcPF8oOrSsgoie4koZmDU185yBLSnOATd2VOHCrcgSyf/QUui760/6qdTQnIS40/
h8YOxh3qCSJkDORk/FJPlRzzbdkkmOd7LzGM+AL8iJogE5428d5aST+5Q/Ke4ZzL
kVNEBvgytxZ+5Tl0y5fi7EjFbVnT+whRclBW5NkBs7QRN8ZUtJ1okVtOt0aaNcXh
GFeA8grYj2kQ+qkPOTqsnfwu+r6/vmbfABRS3WiC6qRy5LYUOf64C1srAVC0TWhe
eVhErqfZ87yD43X43savCbcdjzfiK5+ewjCROCmnwZsuT2H7lPNvHmlVRevKsUst
oJ0dvq9nrPulwLV2GHKSmD2yMfFlvJZxEKe/+rh68oK+f+svsxN4RDaG2wgJOxib
kVcE9QVArQbAtsFKG2Lak4aOqfZfkHjdoyxn/sqErDqNSPDOZMxnVNh9w/qf+5Xt
20ZQTEz/xREfTRUPvGwCCZg14njIj4DyXdyqPHxEXfsDxBCKC6sNOKx4xtBDUzsu
Yu/qdiq3W2eDFTQ69JH0Ty5/rdr1u0GxxORLtGoB6Aaa0uAXdBMRIsR9VV8G/VTV
MV4ELIel8i6YDQiwhWUrqD2kJ+YGCuDRN6oy+PoMRJdKkQOMIZm7+ErP7ANFT735
ik9mmhfyzvUey09d0b8wnJFRKwcmyrl1SDfChVq7G+A0hLtBH6LJ+R6bUZNVm67F
UPQRl8wbNwGz40PIC+wsoWsDRydqMjo+XBFJC97paK1MAtHBjjoN1HtWPGXki/Nn
6Y8HnoUB2tIB6XZEBj4VE8Mt1CSbtXrJCOBZgklIT6JDEXStpcWTLZS32Od072UV
EtaAqSxE4DdmliKBtD+NEUgls9hZsvUOrCF7tiYcnIeTmMK5z2ggqlwWH8p8Je4A
VsB/Z0ko4iTHpNdamfoepL2nAyLZr1SIrA6E9NqP1TvgMHotoMmY3/apebmdBTmq
RHTSILgPev5R8ZTQRV9Kai378iw7jhZsYWwQSyYbd34RDN2fT9YrAMPNe37Vk5sx
38t7dviC3fr4zkVxFDdaF7TYmLIr1YbM8h7fIS1Jx3zCK51vQthN2J0O4lYmuwxl
21mC8Xb9hMhtefXKXk2oV1hxwCFqD3d/CK8lwqSpL/Cf5nVk/rhI7IWxkWl7b1Z7
wgv0QbJTy5/Kl+NKAQhkAjy1YqMNGcw5m3B5mTmVjA7VaH4yI4YRQTozoWm6OxnP
RjrPUq/0jJ2J//Jq6nmXXqB37n9qql3XasXFp9vSn8BhJuvCbUQBlBTDzmXJjgAf
yeglfsKuM3k41C1XiYA1h5oBpIMUgT2qMciYs7CkWqHyn6c6jpEufF/Es7nyw4UO
fXxB5mdE3wt41KM1W2sdOUcCyBqx4L+RTxY6NGqgNX0cWVHgjXN/2He6abGoCg5N
Kt3COcXjy0ZvZXeEvTp04jpjfIPL8scPjqHz578bPp/Qt7agSoqHrj4XWnnmCCDO
tK7u1g5n+CRdeyFe6NfHoo5YeALSvEn4GM0TgMPE039sJ5YJeTSnD5z/ezf5jH0P
h6CQf6xbsFQEIxGrDynL0apVcDqAJNFUcSkDecYwpUZgRKSQcOTVu3mm/WytBMc/
4sEoePa35G5F0N6CZWDITarP7VBlGv/MVSzGvCI8oALYtqB6KIzS2/uhIfvgPQBN
BwE6+lPJvkt0876jFJ+pe7Wf0hxQtnTnUXSTLqtMoxrtVnUMP3ChGrNzMpAdE57o
pR6WSnQaVJ4+U3P5LMgvBAToyvPAzrFlxs+s66y188GuS39t+s3J/ktB9cUVJp8x
s2M0rjnDttP1yrmDusbuT3U0w/0fS8f8tA8HdcygBwIQBoWL5eDswy0to0cmfjju
Vawojctk/3uRR/6WiezuowWg0JcXe86pke7L+XuPs/NMNpDtQz/NHzveHjarg7xc
WmZFzvEm0ttYJgAEqHnvdt5EIyJToCfV+T+JqboE1tMwyRMG0QlbQSKsHehBBIo0
x2RQeumtarIcmOJ0tJlpE1GZvaIxvs/2ZNMOTuD7GhgBQeoS1wNy4kU4UUmja2U0
EsdhTs7l7HNG15+mone+VIGe+xllRhrH01AUDyMfXNVlJv2lz8hLA8oglJ5XcSKx
p9/ccEqpfwMAHQCQ5wQ2OoRQX11uEmU7d7+sf8eTH3dvRnXcJGcniZUuUL6rjUw9
DkDAFdw7GUMhVK3Jc09KXrgd5vQzk40mhw1QIo0VTj8YBO1ijZ1VCEJrFC+Pm1uV
iPWXN/J/6z0MJJccAwwhXyWWVLmzsA0VUgIAck9iKcGI8GZr4w/NRq7tMarSvfdZ
wEyUZcs3ykCjHH0vgz8tH2COd337nTBpnMJoP2UF28NFwlUVpHvalbI5dZNHmIsd
gdDqdnitdPH6gVd4KahZUYLuyejcQVZCL9ucbvueLlfKjNUrGsgEIbaT28fVODIw
/aQ8MoNn/emi80+W7l4nVEvY3ugOorFBh8Zg2v1toeHoTj3IbFb7E3I8NjoByKRd
j7+wVPCklK2oqgbrFZVB/G1BZ7fMjBufeyE9VRM/hNyt3zmnRp4nLtKjHvLX0bCX
vDotUTt9vK5uw8IH4B5oywyPTcX2YgC2m9K1KH9QfzrXArvQH8slwt/g6CpbltEH
LyYPYxduqvYlq72ESUg+p+0R5x57LGIjpTaX80v3Cnptg78lJ5xZoCNcfjhpqO8Y
qvn9h+ZK0IbF1czPzU2tg4URSp4xAEzpQQv5opd8qwoZ2FiZPQ1ZIUg4xmAx764q
rbbZ3ODxOg2URnZ6vDFL6NCFf9Z3bCu4ly1tZc/ZBAMjNK0yKI9y6F3HSp+BYXEP
Ed7hrG5UqRBtVPsBDkTRP1u7qC76Hguv66o084NfgBIFmeS1hIWDcMKVWtn+AH8i
qZkY/EPX+FpOQuRYjB/VJMmL0eF6ibhxdIUscl+vo/fTnp7XAAyaWF6pGGv2Yzi3
9Lj3INmHjY/G7XsMv6cVYm6hRouuWtbZPKD1k2FNNeHMQhhh4JQkwhGXPdvRIu1+
3xYh+JIFeUaWcmTGnjMTzmbVjQhHh8HKG+egr30neBKM5IYCVK9jKLi0+Ef2PvOJ
UcAMr1ujgPduLQlXYcqcBKEWq1uHYkg7NA85E53ydYc7wYa+H1TwaGhs35b56Zla
BV3tZohpDrp69G27PiOoOy7zhQaGQxebFvQgMCuQ7AXZoItpiZFxDaB1ylA60emt
1Sj23tPg20CZVD5tCXa8/LGp1wFpHsv9iBKe2REbrs4CUaRZzb9plVBepO5sFqyJ
TNT1C4PN4M7bQ635Sa6gQ+usCiGP4XVG/seweUDppff7fqGmhVSDA8Wn3cfSixkD
a3Ub7Dmlc+NiY4xXsL1gJMHowSP7c0d+A4/1IkPV+dkoYALvWZtOoeGmN2YcnkF9
kgVO7tdiCSG5qBxlOXjo4qvV6hUJ1XQzwidCyMel5m7mOThvBzU5KIIomdOh9nVi
n8mZS2W6rP/6nEQTCDduuRAU0KXZS78eDHyn4XcI9w8uUiiOOhL9vMBfLSaOp9yC
iLpE7T0zTkv72d5e27nTtgN6ePhZhEtGi+HKi+HMT0qKpyzIcsZzWz7VGtHJ8yCP
F6vA+b0C7YjVzuD/DPtcKBOunDb+v56ojZIl6NgVjhbv+Sxb63FMHTaycFjtaXVz
0+aTAv+2vXOFQDb4A1ucH0/opU+x6v5CraXFwcpVH6fRjjl/UjEsYJ8vT5hXwLDR
VtoKCz3TIqtL3JMG3XDLspOixxSJkaUPiiq7Mov2OqcpQSp0RQgk137Jg7cJ5ecB
bJPHt96yQ7+e8R7+OQPxMadVEfaQEXHzZO6PMbqMRTz5OhlH+3Nv/laQa6EgShdv
7rF0EIeYFFCalfwhwid31VwDA0AaedT4I/5KZ1oKa+RX4k+gkABVOcPySpwcv/JW
eMJxRuah/7hCMkNTPLHCzA+HOjmWdhlUaoZq1QQWhLMqS388irpgDXw6p5MbsAdM
PT7pONja7waurDgSjUtF06vgO7EK991jyRUyrxaUn+U3GRaPofWkqqe1bMYJbxp2
sXcKhyLJGJ2KKsex4/ybvyzfkgq2Bvov8wA/bVd1Scv3EDRJKjFqhDtraz0vs/kD
BNBXYoPRQ3nFjQLiqST4eAxwxSjv0k1MR+BJitwSAzOzIf+9AheyieuDuRweITP+
dK/7juUaGxVsFpYkxbQMP0NiNW3g8ccXfbAyR9EHyUsHDNUX7zcW2c6ITTuwnnRy
JW+uYsgCaAFWc0StggZFGLQRk46knjGMmB2zY8LMvCCBqnpo4khG09eM+xQATVRN
0hBHoJWIt1Q3ptkMhr8uFNBkmpvY6U8r/o1YxHRKL1nSc5q7sXv+XHhqHFWF4Edb
v3dv9fPN/bYGoc9lBwHUEeCgXnpV3kHO3eajTcfVqsxOR+eQH6UENzKO1YTCEhvz
AvAu16qKo800eUnRQUZKyKGdI6vdqr7Lvv/vhz9c9KrNQLgT7wFNCNFLBbGB91Rh
sl1kENN2wtp8m1GOFLOZXoItRWJsKcxswe/V4HPxyGLnOaupJUBHZEoRoGdxLeBS
ATG55qm3wPQ67uep7iccTqWfLm5NOLQeSD/MBsEfP0v0MsNgBxkJ6xig0VUpHUlk
g65I/Xr9bi9ldQNCyTVZP9X5YolI07Tks9lWzJH/MedJcBLwdIydPCbxyBZBl0U9
PMbdraDIsbftPpVtgqLB8uHtX35WiAKbDAfXJbKIQ+0XNb+gLtFWcBY1qgi68TLv
kZo75kVXDYSnO0mu11a6q3uUc83L6K5fxaxdRZl8Eox7RjrpqdXeXh0E/9H1IDBc
OJg8QoaS4MXrvmYx+GY9O9AFowYKUQAZfI/yQNsiA+UK2B/EcdNkf/jfGREaD/Cz
0xQ82UuJOHnjUw/e5zKZxQndBAGhBrFq3Hh7F3IIVkDGkqCmQiRFQok/Ng1XKbRQ
vK0zmzWHIrVuQcBMDXg8RRGdbfCuO0NQpO/3h2E9Km4wO4IgbL0O8j5yb/fUHQ5b
Lyrm+PFqbaG6SOKoG2Vl2EFgv0Ko/Hs9SOuaGkuLRgTq5o+6TtHk7C206hbLDCix
fSB1bKTd4R+nViZVbRfCDLSekYLGoBC3Uit5GF8h2TD24lCuSGUxckfvEbbTXEH4
Di5+6+Nq3AFz+RCY0FABO7m8IjmkYzG2HrZLt/KWMW9VuRVY4UPTYDVZZ7LVaKkK
YrowepWvznGiJ/FJ+ZLwCTsYd+wAvhf1ZFiyB5kNHnDvj3cZAHX82Y+gk+nbEj+P
gfQHYQhALk5M+k4d7geBgO+k1Ox7SoVPbFhFbL7SwUQWDFP7xK8B1YDLug5FJ0Zg
sqIa2w2PrI4/ncUUDfr9BPMTLmKGWsWAlORnJvSGdHgv2vsqfCIJKHRtz/aArQuZ
QRWce4ImYAFl+3nBJ+giVlbmHx4l7QbYRWavhKzZS2X6LhxghqdXAu7neUYNroU9
imx8+vJoAys549mqbGKsSv8j/eneP48ihJdWSwpGQ4b21Pj7IQWI98O8IarhRcgM
+WMumiqVttJrUQqH5J1SrKI57a3dXdhUGinEJbnPvtBrn2oIVZiJ+o7BvVrmj4cY
pShYE5bF0z1dhylC3H2cnNyYQ4f2qrCMmeIlHthOC57hMZi26KF0lDRLQaXbqmwK
/XMZ4eoE4MM88GWA+FpkYmxUonqRPVkzmuO1jQAMxzWrCMOKRM1EiiA4bcT+8s1R
uU0FmZhsvRjiIuOjMm2Rxlpgia6qyJQ74/8DbrJGKDrmQ67ut7e/xYSPOLLlZsI1
AjUxpWWrh8y93mrZPRQ6f3rljUNjoIVaP/0Er88WqAvwl63PUG0pgH5dzN8aNv8q
eTF3pjU/ZjK4+jnQqwTX661VG8xlRCwTcQT0laAnGNBbNAhc3cztNPblljr0fGFd
wrmKoJhK7sIZ5GOtXDwIkutyyZ1bJPJBoGQpEkoCBWhlY+Msl6ETF3iVOZnbH062
vLvfy4vRW9A8kwOipIk1F1laLqCRSeKcIhQJdOVDuzTTdn/frmaqjvD6bGYl+2XX
ySXzZG4gervV/TNeJsyMKEF6MzajaoOmf+w+TS/ns0aezYyo3TlzCm6s+Zq2CFXo
dKq1lgyhV2gjog+Bc2da3Hu1FkO/qMwrEqK/6bZosyBQzE6wimslFKWJoopSZ4t5
JwRu5UAWJaGs8dA5EZF7XBd2QLvz71q+E5ID4bna7h7EJDZAALWM2/Cb1KHJU30R
XdII7efeu8r1dDRwKiW3wnQ3sKuMJcdr3je8blp2M7WqpDxF7F767J4iuxm8wKSI
y6LeqDJgRkiTEdfbJ+HcZHGj2SvYXIN7yrdwMucc3f0vN+iZ1AuGMiF67he1kYwU
BduPtbMbIFe2RSzmDwT+fzIrwbdTXqSuSxbtVCxjZCAtYLG0BVfegnZeYT4rJ24V
SSry4QgO0kkZ2O3eGZF8nncIw/Rk+zzqELehRQs2lYsc8PsZn/f8zviV0jxWsKlZ
F0zWcDdPLupScrivTirba7VnQtpLX/PPaHeo8b3AifS6CE3wK2oHCTDd0mw0Fl39
SoitZRUuwp4+x7bMdcpFu5pijIo6eWAK/fU695/WwUuKaIYXRrFYDUsEkMON0yNE
j4S+fkaMb8rC2Hrixxt6BapUIy5DDGFeIzTc1vXsbVpSZEiRRXy4TDeITFYumVDA
FFdfj7wZEYmRdMuVKbG2KSP8Ktz2qfKlP1Rs8PBe7Opsca0HsjPHhicV3BJPSYcq
Kqmdx2hVuq3yonVHLzb5MyJMlzm5mn5igZevj6qCVMhMPrkoMA8bCOiiy9VkSNFc
rMeHugTwtbGh2HSpoehqwTfRC7ET3JZXVUjvy+y7AOpdJFMlnLSSqU08sIE+5atZ
gmJrpIjC2Ti1RLpgB/FHJFyz0V8UwPKMw2PMa/QLKDLU1vG2zN4mC/u5VZqJkpoZ
Wrfme8H1priwNKtd3QBBDMNdcZc6t0/KxzeG5EPHUJo5fJ0rjG7uWB5fpGPpAroC
jO5zTZvjzeAYziAV22NY9sslDiywLIavhF+NWkzFwhyrLW88KEfqgnd6Cza/8PAR
BEnJQSEc0agdWzObTBLsqH+6Yggdz3qkMxPIfeO3mEwIqgl+YJEb1QZDPXBSmhVF
b5bcRKgQjkYlCzkzxWnrCHv1uYW27XXVJFufxJ9FuzPyQe9NMP2vlQKfVhNJYLuN
9hoQNHVljHBpSvwEsxsAMWnSDMYX0glFldVTdEiBHeEe0gSOK/dK9Q85nonQoUgO
xhm2KrkS5KNJ2ExrOdKqlBJTaMnpFuYQUqia5y1k1mReZYZmTwcQRy538Ju7t7ZU
a87J/8bnKYCxrc1tOktOGyYGNddd6JWLCWOv86+sJbALgFrK6QwcWRiie4abzpIo
w/3hrFBey0Fz+MlTi5uE3nwwJBbkvpMKbt62yN+VtrKsgpvj+FtQh5vW7E6XTaHK
Cy47joZ/CfU3aoviVe/y7jqz5qZtZL6DnN1ZTM7O4lVZ+gtKNL69PXcZaYqz6v5A
QOLkFMz66D5ynqCX9BEQZDP20QLVVvgae6nU0uK5cPIjV1xkR/J/Y9Yvx7/uNyzN
RchMakuOQ5dCR/VUu0h99oPfLQcLy7PMAJFOjTzmwCgekohBJbA8A4waUdNoTg9h
7QYEq+/t8TBKa+m/bnlIFBEu6nV7nGBsKEuSVE/bfdNWVAcvW0pkKldVCMAmRo+h
EXe8N9aAvG4r55zx2917vzpmJri3dEU2wXMzIq+mHxftC1YghiP9r58g82ric4Db
2Sspc5+zwwW7MWbx45SnQt6Tj3B4XUw+bNHvfAClOHhDsdfBKpYlMq7IOcCs3wVJ
iuq2lVn2y3+CMgexu0tcMKJEDTIVxMBfhQAYg1GfNzKpDv/jq7MXTvi3CUUh4GbW
TJtw4qGYSBvj2tzxNvJ+1yD0lAYwv7K1n5BVUg8RJa8mFFGNIwlDqaxQ4skAz89P
T3/5OmievbTgYfe0yKoHMrMy/ej1oMlSVAuuzy0fVABjfiCVWFNu1eN3fc4wlJ9a
6SlM3JxVAuncek5plTlOlspvLD7xx7iZX2r3r7jjxZ83CtFqA0wR1YCTDYDYD8gU
/CZKfTSugSr167A51jjy/wijSSD56minJlfFvsMZf5RQ+FCCXoF4+BTh2IACfySo
XjEoCyzVW7XWgo+VCWk5+fPnDQddfxWSYEZ9Frvhfde2sEVVmHkOvGEQdz9OSIyz
EXjpWsQ3rRpuGkJ4GcKvL1jqaQE8BCsH0s9scD+w4yMWx7X0bTYuv+iqZu6qTN4S
4BqBNvV7bLxyhtxW+gL4sRtQD7/IDmj0CZw4mOQvq0ZBctvPAYbquSXzEPYOEShd
hJlSBIwCNW4GbewA+IQaqqBrW+3EbT3+588st0rdbEsV5SsHT07NKrrhfs1cVDSg
caSNRpWOzLsWMx40MTetHO/dju3MpHEM1dZnZ0/X17HOFSdQBNQ7okQqRMPaamgQ
ZAOv2J9OeteFQ9u+W3QYIIBloYyb/tuUdnjD5Ne0vhenvUO7b0kYyZ2HIBJIuLlU
kuTVly5lKE4qtMFGBoFpI3vsVH8LEK/eEhO3E4Sd35ZRTeG+Pto2Fwrhw3IfYEG9
Qfw3XXdVr8KYPlPmlA4inUiJPgFQzsj4fBFqe/fUxvj434VqxnflephDqtIhJ1C8
bfT6vXwDfifSZlwlYEGZfugL9uzF+VrB5fnCBWEsv7F/cxwLEHdei8m+S+H/IwG8
/AEPUOnGypYq9Vujs1pS5UO2oC+LqqdmZ/5RSOyK4NXQXOaQfmRGykdF80F8EgRS
Q2aaMFnNklg23q4GBivnGrXAcGa16jiWEI1ZBGwd1T174E35YPss5kiTR930W5CS
A4jxjESAJIGhKc6JAiD6q0LGhTC+ZJptbX7uqCihIIverfscwCjHEb0WHcYl9tZx
m9dBxP/yJCqoqU8wUXJb+UUiEjee/INOS45gE8PwySjkxfeRRTE/61vW0FPb6o4s
51kMvf4UsrAAQY10uEb+DpiL1ky9tNM3XLKEbjHR3yDN4C1Rl9yz2R2A8IhiXYrS
NsivA92mbFId/Gzgvz7JZPvWmC4y5PwdbeJbjNeBB6Oagrq5YABazs7sXJBlhC5h
H+31hiM/euPrgxPCCQduHxfmE7Cxf1aiVr/ZZ2Q8O/fyFhsQcn8gIRfeE64XAwUp
xmuXUir9eyq72nk24JPzgdGFc6eIUTupaujIPQgo9Vv1/NbQHpN12Fjkz5YBgyzV
vKDRoM1g8BU1ig5AOuAVU/oVB+Yth8WgrVg0oo9vUVQivAIJfv3QmkkGOajlAWDx
5MNF8hl70mVZNgaYPPHZ4jdsl5gefoR/JXsvxwh1zrBZsSw9IHAoAdfUFJnTEZEw
mkOlLPGWKVtt1vZuyYvOeiJmkcaX4yEsf52q1g+OPaydjnvriuWp7aV3gtannjg+
csWexb7g3Ji8T4ovWA6u5k4NutE/wopTcXu3SQyOyKmeYFhsIQvAHKZtRlXwSO5e
6JIpYSo0FJiFSZHg30bDOngxX692a5JBtcfKCdYzdLjQ/Rtk12PjUDuLN8Y1BCHD
VDUbzdT84FPuTFUoPjl1aLxqCCeF0eM7Es1r1O4T7UGJ5yVsDa6+VuCm5O06qV6E
3JWcIub2NBEOxy0g3bxn+lBaVNRa6MfXhZFw61ED+oQlQze72YiXdr84OboSQ1KK
LVhTqXp3QNg3yRpKR/WHuGVfQTcb4tS4++JFTI3SVpJJ2C5oVmbfg4b6NTqkCMcb
6F6npjoO8RxIe0NDFXq+6hbL8HSi23GacG/OEfdXMSAjKGugnicQrMa1vmh0vjvO
SETq/0YN90mv2niC/e2ryDZcBYJaA3Ba4yPF50X9/KDYC3aAodv48sWBSfux2KGQ
vtnn1XmE4gzEkbmK+L9kgtUhlGGO5jchEa9xBBqYIY9aJcYZ53wfmUxYVqyTxPDH
MdIFQ8o32kcu6PdZnxmcmRB3By5ojr3Wv3zh0DSSmBqOcvUjPp+d9ead8u/rld2J
4Ap1ucsugp74MaZH9TRzYO9l/BZiLVLNM64qBm0iOQSV1gsETTWJLDcVtxlgOj8e
a7lCkR06E+E+MwRDyhX2SpOi8aRaJM3i3GMT66lklh8gXuRN5En6fQ8T8ZGFehHO
ouZcUS6k7KW3tXElL+hDw4jxJfAf+nzqTrh8ADFiHAc/SokBxMaVsZ51XuhOAqjU
9xtHG3yMvyem0pmNFLH+ZaMIlkeDpj+xNtwUthxzeHu+QawaTfEz2Xn8mPWI8RBu
78q+OC1lOK8BpD0Uf57czlZEmhVtEhaCjo8/i9nOvojgTRg+STZ6DCyl7SEieg0X
NTV5m2XzjxaQjk+n65Kn3kbl3mMXRZIDKdvEJlOzbIHycQroRby54l/CU5kicYIV
uAJ6yEcghM9nJl0Lp1GjpXfQ3/CwDfD1LnzpwvnbuqS2uyO1lWgE89JmoDKAJ8Mz
pycUnvQsyUyUZIkOT0g6lhEXaEpKFX84PTPfRuZfVgl1HxQEykA2mHMbvWYU4mA2
CJxq5r1r4qpUAhcBFqT7D0ylXA7JGd1XLUXOjogykkqgtyRjPHBx+xPA0laDb06P
CI/q8KMYG78rZObSOZPHr/VYqlEP7UH0fyt58k6447+VKHVVAMF+eJmSIl6sLxQj
PzdlaBc8jR2b8J5bH5nh2U38g2xXdyNS03lSI5W7x/kXXACZ/F+xvaD3WQO3Q67G
xmVnHcsQ+nXHCOLm3tg47TRhn8/FMM9ydZ4BvohPd3jIe2ip9jS0BgePz4SKhyEu
o46bWdKHreXnsFumBofTW2orF2m4vjWc/efRb6MZB4SZM/ttiS4qx8L79LA1kfJa
p2jTiiXFT97Hki7TIW1XStMyOuInLobJI0/hoLR05c4TjbO8h+qjVlswQ4BdO9p2
9jjx7pdJsrC35OyX0u9GR9zjHvN0LdyV/g5b706NoaGWcVebfJ0RvzOG/nNnEGHs
sUlvDtmF7nhH3Bo3UUKhpJqTUNBwLnFjCb2/Qbp8I5NRFC1HpSRGOJlKKzPflF9I
Jcb0Bs+mmxu0rj26stXfygy/yBLa6mkY+9KrRDAcrFJ4LIhP0SHQnDYBeIVe58iv
AWmGHVnV4N5X28liMoRZiLLAqoyb6P4rl7ZfEJV9b7U8EiwmiSsqAljB5Wpsym3l
KTrKhxlsmydnk+MCcamN6yHB3LOEehg7CyP/QyKPpaWv7f5lMhWRUQRNzIKgQt+R
49cuJxdWkU2loCSmM74GBBEWvJgLkV6i9eyYWvQvXf+pKc2Bc0dBYJjUgY2bzOqs
TZ2gT7grRhHPnKqxoSzxvO0qJKzr/9M8B5ZHkfySx112bK3i5PbWbzJsCm0uzq3k
roaN11iFNmEEJGqiA0fe3oGEofrP24/jynMYplq8phdAa2qNgqigGge8/DDX2j+M
XeTxFH98x9S1TZ0Jr0JXV/pw3CmzifaF83J58D3JgUripw3u24sc67MYsxUgXqHh
enpPhTgVZqEN3Kj1Jsi0+eY4WsSxT6HXr7xutqOxjkkv6Ov9bQVChfiWaJF+NWF+
mlLk63lMT7C1JAhSY8ihdzfdJNTDV9Q4z30uG94x5SZNLQb9qAbcGrnZ+4efb60S
LaYYzdNsfW4vM7q1bRlglV+rialLFONBINQ6RWj1bxtdgZ5S3VmwDzOLzHDxYrmc
8JGOi58lJwRiO3dXgRMQPqoJh7vMPU9QgoTjkFUBFI76w4ZsnthEdQ/MiqqBuX+f
0usAaqDXvF14a09HzSSKACYR/qocCi1CsT5EJaGDJ1nhfEZj4ionqEZrDY+UT/ej
E/IyefO+H3iis4dRaRa5DNKl1maKlz/2EG2JlsnEZu6E6kEebo8us7wwtnoGlXY4
yqcS+1cn/IfIBhCL1UWtJx0cwg3oQcKL2x+bU/4+0G3qwIfKXBwZz0gr2Zin8CRL
IHXbeH7YmAvotG0GoqpKCrMIjdF/2MWQB2uYnC0SUdOfjqrUfAyUnrpoHcaROMK7
+hPBSiiRNNWmbfikD5LT3UPEL2ToyY1vsz315FMCDmaDpnu19UbJzKFCkhseQ0Mp
yOZARYnVKx97Y6RuMnfC8Zo37pfTSMV421rXU8/ktQCUZFQ8yuvsCzHxGsY7soNJ
rTJITDzq3GnRIJiIrfSg5EVJMXRA/SmtH+2WOIgzd9s3KcYh7FnYtpJb4zRaUXOG
vQWmxSto5tGnteEWwy12UxvJRDzjpET9gd6YpE00BrH9ckT19LyAowErbxkc2llt
/dg3fB8i7c/G4BhE0c3zjZW414ISVOy9vTB/ccZgXGdIfkZojyw58BScKKgWjBHW
y+iP1VHOJbLTpkPiJz9DNSelkkqtxBFl3r9YKb/fFsu5MMid12/Y0hsxcX45hpQp
/lSbn5vN7XAfUpz828etJueG3PRN1nFuXk+ohA2i8qDvzY6n4LM1sGPUhqGlO4Dr
QaRNXPJlhttglbGtIZqNDlWftk7TdFfPXyE3AY1WQf5Sdu5g+iZLvXsI7LDkoI7V
Si94XFclVSCI78XYuMm+vDoXmSnDauucWAy0mtF32J1Rgu1F37phUPVWHSD62+zv
N5YLwZAqRwpaNdOXSmBk1JFYmrkaCy/ePQiQmrL/i9iPu/DPEIa8bykC3u/A49Tw
JfkoS1s+epRqoa80QL/y3Q33ryQ1IEds3bodbY/0YpU0Ihw30ROZOwl7oQ8H9nWT
1ulFJOikbiAjQAL/IRgzQKMKDe4xaWVP0NrwF5TbIudssUdtiMQOOb1f4mjBqcbZ
+1TUvF0RvH9DUGValy7cbeKOIwVOB2qFaOFYr/l8Zo5P6ZpOs3T87rXRF7yHK4a+
4M+X2TlnD0AnFOfhWGeDRk05K8661M5UXc6oYgpVHO869CklcQBl9Wm5PekicCYA
8tsi4O0XAcg4o4ORi1jAmIV4r0OJYlCQu8GLVf2KsMXg2F4eCfYy/qvIUNMK1KA5
PNzpFVZV4th+Bpx1ARX59XE4pz10uprbfD+2/fUJ6RlpPQgt+5HgqeocFt4Fhwsf
6/zDDWlJfjz+WoVp3k/mcFazqrUWawwou0GTWlXjLopfM6DWyCablcA736+gT4nE
qyzijHBiMd0C/cJz1QfAF/3rIccYi1vrW5KHMv1SjAjYnaOCgiQUkQkKaTg6llY9
obwmbFR9zwZdCOGgimGYvKfqs7K+cG4tJf/5tVedXBE8hCbddrb6SOYswlwO8BaB
imXdZ4sJ0krbsqZTZI0ZbXDaqzihZLcyLSPgBkUp/uTa+vm+SaTgBlmJ7ab2iDPN
QG9PnsjqfuIaRKe6SMFSEJ/4zr8MS7xR2Pmc1lI5TqIr4Ecy1BUCtMk/D++ShSz/
qMvf3GJCQrxRRTZhzg5hm0NLUaYX/G6iwyIP+MlAcb0Oh0jPe3bRB8rUFiihxKoY
uAoWbwKOqMrsY1jFSPc2AjJWEbAsKCFlP4gRBsQpjwH+NtiP+UveJtgnkBw5gU25
2nAHOW4e8dE+HRH9QKgSGFheGg+L+dShsVXLwaD5h9NrthAQmI9gTmJkyNv1e+C9
q65CHGLkO4TQOOr7MN1USQN8fL2FiNBqf66ICtYaFLOJNwY1MOHRMAW2RIfIRthj
vPPDHG2v3GfnSvJp67TOcr3eQxsSXASPyJGC2VaaItrC8RA87kn4ZHS8B9Kfr+8/
bawPu15R8I11XzI+idxjceJWbHUY+5KKenSa2DxyGrm3IOjnYUVPe4Qq08SjRRS4
cn03ZwD8C1Ryajl5uqSENOYiIVeGtNjYk/cWVFVzSwnc7uxua4kOycHN/zJ/5lYK
Vo+YU3FXSboTA6axGx8z09RV52Ywfy8tRpk/XOf0jTW0VKxPlVMam9zocUB+Ho9d
g874jljfdHyF2bQgTLgpIh8mJtN81yXdpaQbyqRbezhJT8lzeNarLL/iuKN4e29n
FbHM2VnwrS+K7G1/69GhlvHm6m1Tkyau6iuHwyvLtELmQamhO4Qb5tH5p9PCre3u
uuYbSRwAxCwed1H2P01BZZ+az4jEK+G80FljDteu1Ys9UTAVK7kr0ajcaMn+jbUz
jmyART4OH1VefUjKmVxY32EyXgldMDhvGZvjkI64Y63nxapllmOwzI78krkNzO9x
B3VdF+Cu9m4enWoO8cCPEMsGGjYT177McEGEGC8YaFNdzF7uyHxm0HqQUakjVgpn
nKBUJzg6iwukT4HTOru6Bmim+dvNwV/FzLkSKcbQKf1hOn+KQVoeW366efmZ/zrv
efpo2paJBTGtd+vM+80YYbipwKrucj6DrN1tWfdjT/eytBXr1rPAhesH2UqD7OMI
rWuQ4UduSnyd5HMfdlk1KYJMy5m7PipDs3WWoADiKW2Hfv4aRcV6qT+W2wC6r2Xb
99zxiioZ2wuoSBn3So87qzx8bKcCUFsr3qb17WKatH44XfleF7Me49KzgfeLCGUX
K+qyI811HsnqQvTYwObGPbfO4iwXmlDJlGCuN5v7bul9rUKk/tjBECrCkQ4JXwUb
8owHCYG+K90mq5aNTC6SlJRoMpCsssjkMEZSOeFzwX809dXxQaO66na6b+HYqDvC
D5w+m4Kw8kQd7694HQLzZoVDlIQw82lr4Fx/cJ1yOqE5w2+dhpEhVXPSlY5O8B3E
k74KEQjDHpy/Kj5Q2PY/DLxqc30DyvS2QbMRLRfJkWS6cbag0VHv4n/zrx/fiVPV
eq84e9NuYsOrg9uk+Bjw1cJCKY6bP1irXOa21OdU3HMn+fMEAOujECM6DZyBRKtH
EtrRNUjDtYZqZQXZyFySjz1fwRvPYavDZ3cUBmSXE2pS3Sibf0YGgEuTuXtNL1Ro
5yR+64WL05hlVStPoIyj2joz4DEUrgVqP5xvAL5ZOTvUHmnEI4yodUjBYk3fHeGV
ety3Q6EHafSV3WhKe6VeFaJGf3+qqTR4Jam0ZiL7ojH0jHoVemhfPWGwT/nh0hZV
dAdn1wvG5lypEhxfqwPE5JuQBCKGg45/FX0sNWcfup2tYfTrB0aOdqqOM4aG6ecP
QuzWYyuDuTA8c6daJYKxG6cSxD3e39uWiAtoOoT8IQhHxHsv+jrnNbB8jt00RetB
JZVRXrbIStspH9uaJKt0+uHvyXkw138xWJoCi9ifqi6Ci2Um1uCbTMZfw8IAFY/r
TZCsXUXokM6VTm9eWD+U0cjzj+bZ3XhmzNXFzA6BMJL1XhnawB/2Di5cUCgLpzoP
w9V4l7ngptMhovkgzK/rnjlnLeJUuI083GvrX2mqtp6zO/F7VWUDeavav2e06O0O
wtyJdNyXrg9/bMmZBt639KLF5TNrU3hFE5lqHPGnCm/oA28V3298xdEVeaVukE+P
R+1SJLWPJNpvRUfkSyh5poD9QyS84Sk20V6qwKxekyENPXyjdP+dk6R8N3G7zjUm
98kr7HMTtQWp+HRe82K3IErXslS50sxiAEcbybJL5/pv1DcuHvE17N51JxOYVonh
q8549tmsTX1sia2fuFYZMfxIy8EC4Q3Xplht8eKwQf2U4/Hu1CA5StkhhI8Iwv2o
djzT0oqTa5XK/eZG4a2rT7rAJ8QyxEfdnfAeDgtuP+TC7kel0clBHsZoYeC/k9gG
PW/yUMzD61qgyt/9a/3Gq70GHM42ZGevbCiDYo58qHqlZngOII7dYwAeIkbZ3pf2
3BTYB3F8RwhJTghhBA198EvgKYm2McjZnp7zFfTcih4s6f+jZVSpQqrpsTN5xn7z
RlfiZDeixYqo4oOSLkJNzYGebL7mBNG7ntrYZMysAzuEG6Gf+/MZz2kHUT916BQ6
C9nRym1Q8QF/tZRa7GLplXH+9hX4SAk3dQrYavwGtGSEu2LMBEeT7kn1PXry8jEc
p1znWgyQf5EZpwsDmgXPY4iCvYwjfRJKaTBpVtlYCUz/MQE2Zj7vbxjxNRxTwG89
yw1Liljv16JzD+Z6Kx22fzYy36R5ruKKkPvMfdjAWrTiYH72GCzxJjlEmAVKYVZb
FlMJm2yyOm30OdsrLjMvBxTruHbyHynbv0RBerA1kPrAs6DO1XG/08kdqlXbo0kE
GO9IDL5mLsAQ0yq7fHbsVTplLljxB/xaL5S22ERyb397YMYwam6N/K10NJeWBmTl
4DvmDlOnhC/U8XrtsuybDYLb/kg89mV3/3RUWGd7u7xPwCF8Ha0V9kjldD564A07
g/HFBe+Ish84hj0p+K1igUrK8etDafcV69wTR8xZeGWw/CNKr4QEIanT1u9iqKnU
moERAXEhHdzhm4W6uH5IlHUqZQlOpY9aUby0fHZQujlCu6t+muFObDJ/zM3LO4du
V2zYApKt/pmtl3CNh7LGjD8bHiEyqbgziRWo+bZcTPuNFsyFOJVOdZNaN3nkHgi5
YFnQ5gBlLEj+6qgCrS9KvGnzOM2pDwsxpj5J1NuzVGLlHcykgMDlJThjZlRkIHAR
RZS1yQs2AkhvcPBSgSumHerTOwH2KHp91UyU7MP/YVke0vnMzLaJ81Her7YrwO0V
4Uai5Kk0UHdu61JeTAK4wkbNgqQoIOx8XCGceqA6b7ScWP0wpZGKnvysCkeS3wKu
3t6SGOqvqJFgiPpltMuC/08ctBlV4A5nqBcYVDlx0vJVXFbIJ4VRLT99PTv1RUmq
LJqAIk6eIF5vpLW9YW4c6T7pEQ4adS8JsRtGZx8qtX+fAMKdaWoTdAcAZMhJDZTH
k1V/+3EgKF1JtO1lE0gci0Ca2JlyryKzYnhCgDjUQkD9eU3iuHjZMYQGqkmxaQqA
qabMddOj+Jl5iWfwAMK2E14vQHN5tW1fWUFsUJxic8NHkij/S7I79XfWb96K4biL
utSLFA078f9kaJkvqgMJHlfxr2c+PAyLpoQDg/F4JpJOG722KplBetsMgq2+3EmN
tKOwN+a/OArQrBfBq88ZXI3OLhEYJ0d4DsebPSObxfKgUJxa5ZtJnVW4B7goYmFZ
eq1/CXWJ0mM3hokM11ZoLIcHICccw4v/y1Zzc6AeoS6dyFzbWVYMMbpeIIw2ULr4
+QlVoReDne7mp+aUXKg4smuXIx7aTQ/6iDMc8edElVil2Mx/Tj3WRf6E/HjKevSc
nWJvQpxj5otKVcujcboPk5rGUqqXnycPyUJK2Tnf7jTlerZDdyrpdqM0ZviFbOMm
XY7ewp/U4aW5BE8XQQg6thIIgecuHioOGusQoeaHQzKKfJqmM+KgLULI2omqwHBI
IfYViy7Vjg7m14x47MKBNN/bxwbIj/+qQh4dHlwXX71vQUpEKHth+1Tj5uh5tJQI
Q3ojH9Dghh7ffIRQJtb769PWU3rVAGeYNtAWZmXCFEKP9+kQs13L6qqssoQhGr2a
79NsKr7AUneJAsEnkxiJJTg95nYCJRILq4hWb3qFYEL272a4VjRe9dJqfIKijW1F
o+sEenLukdyoLwGG2ZHGIp9+vdwUyocra8Twi4NM+Hy7ychGraYuR2EsD5AYoCDw
L3AwF5SyTfOUn+vkP+jSOL2l3X4shrkftp/HVoTgOjLpKSYBxc0ePT6SB4Cy9nXO
Hife4gArLwVSWuJ7cH00ULMQGjWUClvHYJUwEokS6pHoi0YMnEl66GQq+GlMO1Ne
SjAofiZRc9/o0c8AmsDs9QXyTJ6tpp6vINBiaOq6oUOTk11azgMf0fijLzM85ZW7
mvpV1ns+JiQi0rfbvtRd6Xj+jY0xTnueSAx7j+l8JMVOlWSeAFW0I/q4JiG0uiM6
XP60leOQB/ZjaOmNPARI4m2WjkaPfX33tccFjJlY6dhE1W7njiQx5EGLRi8aK3j3
f7B0mh2EI85XM3a37GViwvBhjfiooVapkfz8S61oHOL7ksvXtOthfvGsAxDUGcJd
2kq2eLUCsCbE5sALt3mFsZIU6wDPr9AoJvddOsBY+OUkv/3hrA3rOIFkpm1AhZ3a
p/N9F/MTvM3MrareM081rzTpAME8t0RuNtfk1vRFlEGMIqdfIz7IuxBU/AKoMnjH
fvD8uPd8r7QhkA1QJoteDETBwP27wjejduAcov0is5AiM/VJ60AM5Z38V1xLGR8h
jZIuUtOcK/GDiWIXcytpB2AxXD4MkyWa8P/mwE4iFrIrq0hAZ0h03ToKV+e+TngJ
RRinxZ5iEmwcXaHGslARa+rN8uRFLBCzMD2aSmNAKlWcst92Lc+kE9RmH13fHIAC
vsm6xZrRCgDOcnrrTpmr5pieNgfnVEX8+dx1hBlx3dLsxq1XXVIRHdyG49GFedLO
9Ua789rw2TrGGkKBA5w2X1e/612IkyvGLPJqga3xCXA/LHLJWiVrOLf0huRmPMIh
mg4iCEK7je13ngl/p+eOqUSSpWS0VVBQtC3VcfXtKg84zq6mAfsQqZACeUozG8Gm
OYQ0k1SAG5Qh8DjwGPUyCbqcixJ5r+jui0pmQ2Kxg1VJ5L3XPLBrB9SDxHRyCG7X
d/6eNqIZB1RT8n4tNexKyhMzIjuOhv7waJTz1ElVJD62NCxK6n5kSxsp6s0x69MA
YznfeWEu2Ig23xJyVac1t6Fw6USZTWCoZYVwI4JorHTdMVtdombaecL6d7QLrF+D
DwhxZz8lvmqz5rJyQ6Z506psDq16ioP2rCbZky+np3lcFpiQoIYHoYdNUt0HQSJW
feK79LgLvRiotcq+/yVTeneenA6vFWgt4GG2IakNktnR6m57ke3II8qmp7doOFUR
0x6Ms1y0vlEiGt5HSk82tH4ctA6mSnWdU5a2oJYTzKMHMhJK1jqkaLZi8oR/Wka7
aHxQ8rr/bXVahh8MXeUgiAC/PmjpOWqE44AlMWwOGhM8Es1DHaXU/atHCSj8eyQT
doRGWIu5pS0KBYltRHApNaplFaj8209bbCidUHuWB7VX/xDtdEpnylR1y9znTcLV
K/aXsO+jsqabA8ucOJaaykn5AwH9DNZv+zrc+jKmhXbBGCmChT4PWk6UJdQns4VJ
JnYfDPgVeYTTzfV/sEOZfyJol8qgIyxrVdYFSRaQOlkALth78rrl321odLNXXpK2
oOF8BNVKzQjsuTaXK/6ZgpvImRvkui9wdg7496Ej5IpQpfn0fh/58FmIzq1IJ25g
f5EixoEJOe/AlyOEYU+TsWmuFeteufpLg86imwX0aDhHQv0Tfu0X+iGN1GHUJ1uw
ZucfUagzd6fM6/K4CV7E7fvEO2xZ204tfDh9NA00DZDh3BETjnGIr0NNo7Eq4umQ
Sd/qC1vlv6IsAj1fBhreh9q2OL5h3+wdLtL0yFTIwd9t/MhszYP6JGi7TBngrj5F
qMUtiLWr2bNweMlsFBCFqCJauwRRuNuy30mg/x/pAqNvfkfDsnF+hJTvEKm9MJKM
AHqOf9ZKzuJAbfXEyrgLWXSNzgG9E4AItLVIKqnKeYxy0LcUxrepJlGfXMSF5f/o
FZ4ZCgSXJcriUS1KOmE6hl+DHnx2DKf6wpNIEvOW69gpdGkO6yqydQflLBXywJ9h
a3LT3HyP/w1b/nThVbIIm6iMUKGest69hQos4lOicFk9i3+wk0iR4TuJg07/JJlr
s9DFxTbh23SyP2sM/gIdHEpIv8NZdSwHwjjuzs+6klyocexiZrnXL8o1jyamH8Hq
yEwdDoyTWyT9jXZpYmlAIufDRs556J1GjJZR/CKmnxeg+Et0WuYAe8LnYop07XO9
M1WquMg73UUQZRDgpzOrwZFRiQCM0pdjWc6NtrP1CaM2BIoSVU3JtnZH0SPS1zIi
VcxnOmMuA311et3R0Pff0jCJNaMSZCYY3EZGF7JTdVcO2dyr6MufIDYzhr+/fr6W
GkCK8GBR/kpv8U4dQH42cP5HnaXKV6v0p9RMxp0E/P1Tzp5koAiUbpsHoprzzFLK
NsYXhzGFcCMNpHHCCKX0No9HL550QliJophahqsOKjlhPiD6QPLcVD5KL+6gu58i
q1p0OQCxVWbGRZ256Ia7IckoEJAmL6HwhIrGDhIxCASjo5tisx9F+XFrTFSMGiv4
jnpWHivHUsHo3qxxkYnctHJeMD3OlfBTaMtq4BvJ45/xPAvrmQfU8gjt2x8XuQ+e
AtdArG0magHDhOuWAdO/yuj4HZhJ47SbUG/wewksQ5P4XAdfRblskF8jnXDLfqye
tpC49dbqqbiyUZDPzp/rQGy9MDYa+voHuN05tknL83hsqRybepNbCNyiDCu1ZO6K
DpPgYTN0FHUwOmQjbhBpXFBemrBE5l2V0Lx5ZYNFsGdoI35yThuGLqao680RHQAe
mc0/J3H3WCtUwqTcXqzhNnT9pZ/0/um71PEOmYmiXA3XWwePRqb3/y1+t8VOvQqp
On7FOoG7aODbtf6qNLPvsPeNvCL+qle5vtAr4TW7fMHqEsk+b4MGqgkHoa7ABaJH
oR/U3Kr5NF9/+m/VwgDWNwZmIgLwtdy3FbyDVd63QGXdm/R3b8HVaycX22Jrku2L
ahliMLZo5ZkHHe4QqnyI3mdEUu2v6Nvn9IXrFBCdttRpi4Dz8PNcSVoZ+q7TjoME
1dhl2pFFMsgX7iWUNIqdI8TLrLscMPIuuHEi8+qJC27xMyeVyKr3PkQjxujg2xND
ND/Ox4wzerK+ck/ffSI9z1S9xN1WZOQTP+CX6NxJwPk3GdrbXiYgf4tH/L5zJ70q
s8yKGiaMQ6jwAj4QbRRC+v2k19Tt2Oec8hGncuyMr3v2eP0Zta1+WXJFPz7ZL8fQ
oRqu4t5fElmVDhPFr8h2FlPYJbjp7EH+PhH4/zAc424TJJPiDEOwsYujNQQdiZsq
hLvJvOBlydOlvZwAHOBb6TIm8nsGO4woIcs2KjtHZi0O6EedQrHD5ufqJR927l4k
kCBgCkdUbOoqjCufCvN8H6LVQK8d8VU/u2uuVSHDi4omHFedtJpqa8ehSJXZp9y/
6cmAkCNgeRRK5VJ9BBdemwx1hTy+Pl0iHE11IQg6x9msFPEQAUnqtqy+gTF1BNuv
tE8CtHoNCL9ljDLpGYUUpKW1ILch/BDPrmFocofqTrG9Hm1hGGd9P2ed0O4c8M9D
2p962jgbF+37tfltJRe+7/n2VAOUchdS2X/8qhEwMPJ3YfEN5t5fANchLiPbU/wz
Ox1KShH4DFJdeD761DK4T+kGYGf7jve7kasKlC/E9Pqsh/hh6sE8mGWQYyWnV5t8
G/Mded8JUIDI3LkutPijCf2cNPN+FaCBvEJbSZGpXToxzI4bnX9BkJEGWTaIg32u
dcorEvNt8v3Zi3CAIy8zu6DhHmwh+1qlawwiblYQXNXZ4ILkWodybGVuU4XwXyHA
E3V/5F0HITZfABeoYj+IGlkb3v7vzvxn6puPxd47erEoVB68ES4Pe8ELNNTn++KF
4to1H24fsTWMVO+xaLAMeTnCG6tJr6CDujKwMfEi9Q/oJnLZfkcBNX0RFc8R14E6
vvlNWnw3gkxGP+Ji4meqkgl0WAv2a/SWJxpZpF5Irc09Azb/ZDag7EJAVCXWL+CE
XbtH3X0lN/KSIFDjtmNKw0Wq/gWIvlZPwyYvU/4JxbjCgm/Wq5RWO67iwMYAH2no
RZtXO//wM8SOsbxpkElfGhyfvtIvcZzqG4sHvcE5zjS168VaSMPGZ6cg3+LUC+Bb
u8d7hUhKzg1VHrrL/uAgGROeFjwKOZstuYevTPxqNi8EdciHeqcT/JpB78V1b10E
Me5yqVUKiC99IIhzfjau0OoKrrD+e/wlLm2Pxz6ZUVvhte4yMieksFw9BsSHryFm
T+7x8bF/72TC7JTWmR/YzfxYYMDzplKwFmS8Fc6Edvx6dBLs1nvO0OUyDY95AOUP
s4rVHfjViN2Bs0KjPJO0Pr9Owz5odQYx2cmHxUF46jlaMXXE7CwbL9SFju1hKuWT
C84I0FsyCDSFZ4Ll2zlw+bYQt6xSTga2mKfyq0aZCx8im3QPzooh44JP2keYwBP7
bLFUgMzZJuhePFFXfSZQU8H9X1tSMVBN3seiGV+MqaGE/wLMh2FI0qVFqQylR3A3
cq1DDTetq/qKmHqaJk02HNqqosHap6UAPvVenox84ZBohUHV9U5iULAk509z309y
qUMg+MeKdqDPGM49ggn+euvNAn8e5Tjnk40oPHQmruTolv4OWE0e64rbW7E/fxgA
ctoPyajYepCSAMJlvNb4kctZsL7Nk0uJRoGL6Pe5n93ieqr3CGDT9xVvS14umvKe
FgL5UAyEi+JRjl5kdMR4nJfqRuSKmgEFcShBXja4ZG3a/KKNr1ACWQLOHw/hcemZ
G5Up3ktdoYuCTI6w5fN2aeczvLCXhJqM0CHxHnv3gzIR+kfdEJEfTi6HnTQoPnkR
8un+ka1fx7juMTL7Djrr9KEwOQuXtFUOkgmdJalF8QiCc/YBAnpQl1rB6jJSZcWI
a++RxA3dOQtbmwvxYfxkyACqzLix1VdtgPZtt/Swwgdggu68w1HYGLIZNa77qmIq
x2ZTgw4oiPREJktASfNqdzra311pZfl2WLD3ypLLBhXhOrtw0LglHOgXOmAgEjgy
oT53zkRKrJQ7vA9Yr/mmmQL4Rr4084zHhxXA7lLt/wYiILBI/l54tYblTHKCz1bo
f3mFPfQMMGdQ9WcZa++qYD4gUGdiIfxun5YVq7nb2xaXnmNq+trIjX2BnpArw8m4
ImZr9epoXvst37g+YUIL7y+yUK5czmWoAzSQiHICgAowR4GJds6buzP5m+xBUGz/
KgqvDe+lGidoB8aDQUb/9dhc3leoqJMoipUH2cQF1vVFiI8U7o2EunEVTp6IvLCB
yFqX3GcthRqR+gSzKtT6R69559XGaSCgYDAPBqwvSgKZ6fvDSWMNei9/8rRTyzAn
TSm2C8et/AVUBZ2KS7eC9Cyw6anW+YNX4vOPmM0MgPaEhpFN4nN2C2nsvPuk7rtg
Q5vxI+FkxZWcQ/cr2heHIHhmXpX0ZWZ+jvNDvHLjgqlCqQmtfTNif3OaR5VDddJE
XioQySyhOqMaTTuyiKOAzJ1Yb/vaGWWqyeovrDisnwCG81+Odn2APYmYzC8laRDe
4b80VVU3/B+DEyksqr7NhbdOX0ZS/Wu6RFifSKEmjhngNR0Y6q6TvoJwwYBWXJdX
sSBm6k4ZWwtdNiwSs30JCNwPxr1x2ml6jrGLY4iPVBkMImN/N3TBN8K0FziCusNM
0bbOABtza+xYfCyHF4J9Z3PVwoFwUBthnHK3oXrN3oYNbUf2A7D8yefG2zDfx7mD
XN7e8bvKcHqi0fgj2oJDUyz7RPiDTCb98BK1DH3+KxEwpEL66LslBTw7QC35wfeY
OKfsZ8rXZiMN1pNViUi0cG9D1rRHmeH10Hd11tXGoJHZduifa/byMXby0NiAVUwB
5J6T+pJAsyhbhGnFr37gt26jFNMWXfiPQh7TNVLM2l5zphN4B1/RcZ/IgaeusiSO
2Rxw067UuhJLyJU/vtAHX1E2FQ0XHLlT4kWeL4Mdp6Y1qUYCmh0tesnY3h0e52Nk
k4zUIZ+Z1k1lhp/UOpxEVtaWlMHDsPQhT12QCsK9fkr9xr1+zBZizAZ3UpO1ooeE
FzXSyUnLftSndQN1HtR8tgfEcwSNnc3sjsf8yWBPqFds+EGHKYYWWZHd4C3Tf1DK
UA1xy249pctjF8zpki8nJ45CeN8XErFdLqM0+mPlOT4tGMyo+WvZXT7Ap2rKZRaq
Pm5enA0nVCMUBFJr3Cmt150cGLzJ7/oMNXRZEaR4pVBstZAx1S15susHzN0vjr8N
K927BHdX9NntTTPF4exARK7Tb50TLpB90BOMeGXVV95KcjuNplvgao6iXutRjG75
ZyY6NLLjs7PZaD58Nb3rNZarhzb8z1dwU9b65SS9A+2/GK+ntlFo1vluMk9V1Ing
bD7qy3SZ/qVBQ17lKguFKeEAZ1g0ZJXwQ3kHW9z3dgGwFADKOluYxxvgfi6NGwbg
Xu/ApAfGYITYrDOYeqG8HeDz+RqqPr0a6IQOZpLwnW2OnPSAikufXKoc0mz0DhTa
sT5h7NEQzq4gXr8eguFH3gc0md98zpzPuDlo7Y1FJ+pyJw/dAzUZ/bcTAWZnD/pG
RWPbrpLKONa8nvwxBUK5MJaq14RHKfW+ri3OSbmIy/Kq65dtT9cjewN0OCQDDmJO
L7xcIOu62MWecpA923o0XYt0lKovSzA5cZwqzRuLgV93DLWDqyo7A7hc0S8Z6zch
Oeo5fwzJSgalTSv8+kzA2xVmMX4zasJ3GwCkb3fpbPiLptCEGJy7G2gdIReyzGcc
1nmPu5fYzQEFWzunitytvk7/RnfBeDgNAZci5y4Za0QXYoL6GPum+ZEMblBGHTrc
CMA6dYJwmsJfh4PX+dZikIlcGwtbuVob31QvCf+afpsxS9dYq3CTGP7+DvuMkeey
DebTGbhMVXwd8OH3wAVoG+rIp/evB6TlSuHkTgp89YQ5FdPVfHXewZHo1mBh7vKq
fEquMIXsEcsjqIWnjGMNCyxgzn9722NOuwTgENrytBm5nYAtPpGnalLIsnrrd1/M
gIg9cuoN2UIj0MWJPgc2rWzmnRSOB4slb+nKT2fosNGutEkn8HnTSyRzptV9C0S5
1zkQ9fUUCpC9RHdEqZ1Hc3T/5X5BUlCTZ3H3I4dTHpUzBGBfXFJ792FNohL3dsux
4YqByoZYtk4iDTe8TmKEvsPi/URe1uSFLU/7eDgQZkyC15Y332wp1oXLcq1n+aH8
K+X+4YdNdfWFRd/EJxcPM0gaD7elgTbUtMsvT6bnAD4sN5506jtcjSwrkMs2zceT
yHccHmW8QJVIWa/cd2VoErl/+90k8zpG3W2WotgOnqokYBmiMqq4Np66CP23MhYi
ujqMbIrijZG+pOStov2bBko4OEdkIxTnlxcf0FaA82S9FSWkSpRnRXDfV4cIbtGN
6yk0c4HdgudZuciCWT7sNMyIhWcZU3HH8q+3AekSStfnYUjXXDjRiuCERQFfmKY2
ieDJJIvg5NTRoBxGT/lhPRIFFQp+dhqVpRaeuUcyNWsKR/oq/GfTTfGo9uH9WHH1
2ndFjqUbp/tV6/Dij9XCXscCyoGok+mKgpLmca6Qn877G17QCOdJBP/RbYOx6m5O
p8yswf/OPcX4W+h6TZvmhE8nGMimLExXaXpvDmGu09w0MPwcRMDzMWpVKPSxk4tp
asbC73Yj1WvcKju+4n7/X9GNq7JX5+MIfHMDmyD9yOvZYlz7nebFCT2MKiM9xoCg
fIkNIBswXkOdBTyIAkFxDI+/oJ39pzN/Yg+KUuriezjgr9QUgV1F7ZJTYP19G1zj
rQOQy5LCPLxmPCCEEyG94s9DGIPMxEk+bTaIzi/xNpBilodMpiwEwJtyXo0PvFxO
dujoDsvwUXXgKjBPgDyTQIVHKXk5pQZ1gOyVoDQhoaKelwrYo8t5N4zy0YAdZvYP
N1REMIe5zrkm6WK3usV07Ei2i9yC3o5aRKjVAU3aKFbS4pPC6VIsX05s5FFHjx0D
YwsLU+97s3fxKF3JH4Qk5vV8jAgYeUG+ggqPT8tzYnXO9Q+23K701IloXBp56BBG
F0Y4MHMTUaqGc0PPdziLxFhg4p+jeQ/yf3UhJExjmC68/J88bDzWmVsGXBcAMVkb
1QbqHucgi1kPk5lAI3WtyCqfdHZtokf0hZUtQTSvqcxyFdQXi1dTFQosGK3OgX3W
aEWz0X4gsktF6AKOb7t048mDKN4aNcA5qqkRNuDbNE2/pzdlWpKNNCvVekZTdjSt
wgC9guxFz1D347qGTFaKgwFn8uiBLdlEnS1AE+0NCganTDztEByou1Ise2tZEeMR
ogNJjKT2aGsnQFHWgzVgioW975ZUCYiGbI5MNb5kSAEYblNUspOFil3SvshhPKK7
Wdx5DnZa9VP0zA+v7bAYsMpDyYtGCXEDgO3Uph6t9UNbst1QAGbcNd745eVtB838
MRkINL0Kzn1qZ3IhlwZ7MaKYMW9oDMEyYJOV0CvgH+N6I1vxQIWR6TGQ0z8XjgX9
NwpEgq7LwgcwgkjmlZMdPz1rHJRxVEpQgy7oAXl8x1MSnAhGIIBGVN2aVO3LP18G
2B/3Hw3D6puaUKB5fBqwM2oCO0zg2uhcPTf60DfSXMLp6BIEuzzYlV56aGRwoBKM
wAIfn7eOiwXyktKMBU2B57UoQAkARuTVLHveSs3Lj2pWBkPpQfZBv7Dh6zuGpORj
ADH7OzzIwlwJtikRVLpC7igbqMIo3PR9UuVsKac0a4cmU8I9tPJkN3rddu3QYP9x
zIc09PqPds/wQOSc+Vj9Zc8agnBnpE4rxvDM42udZG3L/9An75EMi2MclFg5RhC9
mAc2+4hA1+1oAIT0L0iWUOivhdSEPWUpbSwx76r8u7EHoOEO2YMqC8Ni40eOujNI
EQRjyrPM5bBmyUcfiB/ERHjid7hn6aR7keJ6ZuLTRZmdyY5C7+QvpEGyMPHY4NTf
XrIHPifKt/lw/If7iLnmp/uP4YTLDhpy01hPX8eKiykFAjcA6u3KTT4k6HbBgVT1
0uzKbjmL0zj/zlITx8OUKjpa397ntv/vOoIUflzYTN41zMdG1KFSW2Z1LqkaL22L
B+S3n/nrxIK/USW/H/kldBUjUD0Lnt7HRes4+XeFRohWA9CFGM0O8bWernB9W3Js
YB5ErQLNu8eJWMCb2w8u6RDOMQK1RVdW+uYg0ue/98Ty/uucFQTFGCwem8RhErA1
5y30LTwr7AT1jDnrU6v1sn6mcYAHXmf2yocce2kGkWaaf0WgRZZIGYE1EGPXtXE8
Q7LUt2SeNGtpi0q54AdU9/m9xlPq6N61EFGrLQ5bCYTf40SParI9EaUzbIir4+Bu
HydPxwyHA6rZMIJzE5W/X4pA/fZcpa/e2fs4DGs4x3e0cUCVVVmwW7xwo/V1nrij
vtxQJB03TdNOOWkblFFy/OTJUVEn115+0hfy3O+RZ9GztLLIzI/Au9nUFvPbdGBK
Xom1MsLmSCH6fb5tsCLqy4OhiAjiYagBcUAn6WIt2RsV19RAaqpwaiLNG6meLa+B
S/jqGOb3W5SiGE05Oim7M/59CDZyYsja9lFeJupqjFMxBkQgeGyYT/Ki+bgig2Xi
Od6rHtWhLsktJxmBsiFMrvlxDwI1xtSaf5Y+WpKQPFH2X04oDFKw0PWFrKPgzo1Q
CTlJ0HveWufs1vZJwQW+tj1UtYeMYMH43SjKlOnlH0asY7SNzR181dfGhEVPYo7P
NZ9AKaYXimC0c9+GcfRj6fgLdjvxU1qG3t72pcisOwGPPVTumk0fM+likhCdu2E6
8rmeoMjkVWo21K8u1aETxtyrEJsqXNseosPayBihh3Ox8iZn+fVMdlkgf44WjSWk
/jBVoReGRPX9w/6uUrwm5cdN72ELu3T2E/B+1l6i/KIvFpEa0QFkacxCgZK/ECXb
mQE8n0qMH9+/oMVLscPuVEVk/dspnLZUbVPg+oiP26lbLOBp7Sr6ls9WygcgfWR9
8057yHOd8v2dCJXgXjI+qc2y9FkTXL7Gc7IxnoTUK1jRcjrnf4VScPDe/EMjV+M8
NDG7mSqGN0pC4mw5ajD5lD04tPaRQyr8NNxlNjILP355WUWIePotqqRdxYWs+jyV
D/Q7oUh50zQRLzKDUAbNXUH6OXMcrIDpJEwvvmZh8v68WNhdnydPm6SpX13aKcqz
aqpEkc2oypn0j5t8BGV0I2JusYJmRq9SJQ/JqwCKiEUBEF6CO7a/kFzd2vj2+0l2
PwJFta1pjulVltiT92jLT5J++pJlZpNJGpGWmx8AnG5nKqkjmOdvTUzI8MJC/+Jm
LsHVzcRSGEOCNh5jM8H769NkW5suxb3j15+mZwOz5nK4Lrf3IAgt6ZK/ykkk4E6d
TwvZFfnUd/OC1ODbDAGnuG/Y864thh+YmnfwWSEf/+CdD5t5uJckNLWdE1NfXIS1
7JI4NRai9TsYf3ICLy2MQmoRewi//FmpbWzF12jMLZb2Zi6ISpabAWnqhxMGrc2f
ieGPOAB0UgoJxuF69BUtfeFK7jQTpWOftbEObuz8TKXozMNY3LZC1EfDFXS/GyDV
T1RgazaJdwTZbEKpZegrXKtZzlj6VJX+dYwC50hJzJ56DvBzCMdULAJ/k8iW58EM
mW9TNpMZMBCSAiOf/qhEAwbCSDtECPN4/VvOpcUDL3FBsA7TJhpZbw8z7mQl0cew
YVBU/XlUntfxErSD3s9HRe/x352keMMR1ghaamOfdwnLuK0UkThL0AI4Z6pvmA9D
1NZlZv1jXFV5aHIUDKWe8Siv0KKCMDR25WNesiE/Ot7q3ITl4G8zHYuv7Wl2vowq
AHcKQ/hfZkLy+bz+zli+NRcxixGF4gpmKMXKrUngKDlxTc8zODHI9t7Oo2Xr4rHL
idcwwrR+/sCagjtz0+PFwxsc+b6BufMl3/2pR5u4BQyX5kzLQB7ptiVueRsOOZkB
zbyZ8I1xpDmZSZBidGmdz6r8sepOT7VNs7++2EgqfuPjd4zreBWfUsFkD+ZKmPEZ
mn6Vg8mOo/qJbYl82Q/0Orz0YCZRW32Kf21JG0L+pwpLfhpJGq5/g3oPEIt2nQFt
NGPN0nZvEmSvf757WH2z+OuM2amuTPvoC0YyYVv4XatLqTD6DGlXRFNmsiAjWBE8
88TRLUS51lBrZeie/OgA7pJamScB7OjTVuX8bH2jWMDc94JDPQblQAQFFOLkP1Zl
6D/1hqbXK9AIlenJXwoA6PF5T6EqA1oue0ZRPRGIs4kzCC64Gvo8duPWAeCdEeRg
awSxfgkTYmxVhhAR7KicsiJzNc3ZWbSRBoD2Y+gLvDj1iPigVPGjgHnFPLU6FC5v
9ZRCV6HGDCowsnqowxFK7p6oIn+HhFiZA3PDKN2v3b7+hP5Mh9cKdUILZChyvHCW
2EmI1oBj909Ncht4E5CSrUGwv8LIIu2EJJarRCrZliPLRDenAD6seYd4iF2eoSGj
t2xY1cj3rdxE9FRHSzR+pUjxdHL61JHFdqhSXLWfuyfkAL0oGYeCWdtJbCquLRbV
3ueU/xZgHo9M9rCzb+eDVzRYNLV0SFrjQj9o6uCnBBIqNz5W0c7wW7St3FEOx8qY
5clBwRY224UGvPL+CDMlgf44fLA2veLmeT5IbEw0+fiNhXU4D99Ue4i8APn51lxY
nxR3RgpNLXcvDJvPhCnd4bvcpcQWKO/wAKR1lCW0YLnmdSVarMvQ2uut1YgKIyM3
R4DzNs355X838pvmFn9J4Dzlmd5h1SIFKXK+8lBv3Lvgb98DxN/ml9jX0BiFAIyp
ORWXJ6Q12bPXuVoEm8vwxI2F8+mzKMV7w28DjVqIy8j35suNHB8GtH8D/g/+v+OL
hPrs/XgcgKvxnNWyxdpeWhg0H0qozRe/LgF/TulWwibqrUEfURnnQRqjkjePFLgk
WaOvaFZJRM2WjXEVV28bI4wIrx15LeTEg4UZ56kho4mrAXL1JRAtX80B5naY2OU3
ghczH6S4dQn+gh/CC0Zp9FV8eAZwFYjgq+766WnKk991pmgHw2orkg/YW7rYyjkR
hA4WKi/jLOo70dsJmEoKSF3YVKXyT8/Us1PmewUilPvAVkElHlgcpcxDS+wB7XbP
00BZMtQi+hOhGkjP2SUBfCb1tKhsfYtzp6yPU+JQSg4KTYarp5i8zEsxfP5HhwOw
ML91J6i1rCPkxgJ32LeKTRPAiUI7gu3lLntiGLfKp1bF6TKQVC7tu78CNaSsKL60
JwE8eC9cIuzJLkhg21l5eGIBB+40pyRjjpWYyRq509Pc8Te6mZQEkTXYcK+Dsm7G
5IMW2E2qJjFPi8RycQ67H7kGwPMUe3C6qeLSYGfw0CFX3WXO07mFIQuH4NfQjq9H
G3IHpLcBWz+2Gd1FKQIGiMeuKzqdE6S+L4pRALq4V+Pc4Y0psKtjh206gAgeU528
Eh4A6QAcK8YTa0pYioSKq4v26/ihlZEHEMzFtQKiAVLT8fp3wnegf/kQB2b3puGE
7b7YRXr5wJMDWCnFGHXx0VhvLqnXFenesYwHivuBhG+WJB4Cqr4P0TjP6YZOFQXT
kKUjwrLswmZgBYs5d/Ogr1DNXyoSi59tXiJuzLF27jfLFjMCnrTm+9YEQvhAvT7o
CREwNRvbA1k7+JYt/rTsLktu6HjPbCgEaYV/mJajGMNeLBwpB40ODi5T78RN7jrz
wRkYU8FyMAiWYo2dypXZ7JF13XJbORsiIQTFZA1k/GpU1kd3e/rI3zHs9lNLgsHJ
1u2w8NyZ0C8vW7ShBij26XdzjCnNz3tBlQp6b+9SjyJI5Lys75t2j4VY6tJ6b449
3Pldt9l2aaoH6R1TzMxmJmdeYAQdFij7Q9KFk6RwCkAbSfANnZvUhrDig93OijEN
evZ7ncHMD513ki/pMZXgqsC2RJl5RNXNi3bir0Y0dbV7rafbYwhWzmXeDeg+D1ft
d9VaGxMWRSqeLwaZ/iPL4ZO+LD1icah5inbtAChlU9SYj21HfZV2vARFr3ZzrKrZ
rjseGZ3yZ0EmLFSPCrlBSwpDFivxFG+/Wo2MT2hEL5eb5kU/kXGJMHfT7vFiRkou
hJuEDCGlMACFHR9PTO57cOKnt44zFz7KiiGgsfJPKRB0oi4MlSl+5btNhxR3DBeo
xwD4PEXKO3AOEe17V1QhZ7Va9YyKaZTmEAk9sZDbd7nmvMGEDHkr1QmtLKzc7plf
D7qNgWx7PzNhk/i4dMyyULg9inm94P+pBwtCAM0FSD/oeateSOhH6wyCzFyd9uKF
FVu1aSyTYj3/9CsGsS0uOTSPewTYPVL6pUsPOKIBntTHmzum4VTpZ/hG6FNhO2Tn
qaenlPeHhAgAwzpzl1NxKmOiIvuqAFgghpuEzRHCtQCpJ2QkHJbXg/msdPMXQ7ss
cEHKoSIXjkU0eIIL9OZn+9VeyL08AC5bMuEmZANF1p1VGQPUV4Gp3NwOVYT6u+5C
sEnb6uCC/pzRbaoQiEt/EYrxxJHyt2tsJ50dw7hjsfPlt9gV4BvsqqEmzC4mMfXN
dbJj9OCIat7M6vv4V6hrDtUaMB/0rlSlS39gnrKcnnscG/tYcJAxeNcFlivlVqIH
zDFcY/8WDJbiULItRozG1LjJG4iofxYRAXYRDxj/hV6jNCAQ02geuElrYGQRY6zh
+5l8oEGbJBH90GoDZX52WfZcsYNLswW2nTqSlpdm5LySHscJ+/G2MnfeWrHSYXJ2
6Mt/LK2QeHm4ZUInDuxZ3k7wci0AVhuvUBOGxihImmhuCPS3p94BhEM5/+j/cvYz
ejBEljmw0b+NBZhBK8GMsA0ybo67i8S8uHqm4HotSVhDyptyWDDEkPMn48bl2Llj
m6qz8UbmjvEBi8bg7yV/eU1v1kUQp/4RsiCaDISAg08uDfEilmh/3CxxXgqmxacl
eY0894K8J9m5lTFdog1iaQ/umt5omSaG3SEcrVpUeY0Z/24opNVxzOX13pwG4Kqs
WTXU0ad7pcDHK5WHMZgbjwx6MDQ1JrsgxNjqddQNF1IdFdxH0Mq1CYZEdu1PL1dh
r3nhgERhl7Bj3wDBr/1cSjIBzKw8VywkfKlriprDOwdMkTUdHlPZKS7Znq5ydQs1
ot3i/AGIeZrCGbOeb4gH1ulYfeTVJomYXEdwDjl3aW9yFddaORuKXvmWBPyfa4eJ
1LzGH8hwfw6sIaNHu4m0vGhcwXIn2VEMee8TVrnKDrBLSOg0w9R8xlfmW7kW+gfP
eEQgvpOPKRMr/tEOTNwn5JDOFSzAKexbObSQTr/Ll9cOYzmFgDhN6XF6peljJESd
vxCroYP5m7jNryUoUvXn1DlZIf56pQtz1y9nyCpxL4W1Bp197/607v9KCsI1g07P
ynGGtXdZYfbMeSsnAmod2HhDywLe/DC+yDxQ3K1/nIb1Svy0c/UAJzUdKM54dxpW
GRJWyfcVZwVyCB+SRiVatCzoduOEh92ivclZr1UoyEVF6q2un4nesmemcrSSCTSt
TzMz2fTtUjCI7bJeixyA4ltn5OiCWBfejMzeddanOD9xwC8fGAS28lA3PECgOPpo
EpF8xhV9m2rHa67s4Ubbm02IAHxx15R9Uq4uFftbTZb/s6FmHsARfnDJZm5OwHqq
lMbMwEv32fUtqUYbP92kSZ/WqXLi7Qc3oldW+5ZPWNaUyoHqdyHBL7BBuNtpDj3o
2NtkCKG4S4GUI29McrOtu8vnYzViAYyrpCNQktCAXl18depeFOm2CnvxEwpnBIQS
h0ZeX1kpMipxvnDRKOJ3MAr4FVui0xLHiegQwKvaYXbrzocv4B0FhQN5ndXp+/qb
GKwbIzhYLr340NHFsuZkdeT+P/GiFu1k/YrQgaAqyGkHbi8Nr6dM5rjWNa14yMJ7
i1Ek1ssxUujJaJdkQOJBIKXPj26jQ6i82YWL3BRt2ZKFWFqUK4R3S+mkbWlNKQ7Q
SVLYbXw1na9286A5KFNz/ntcnWrfrGFCCyRJfyA/nLXqtprsKeNHuwdf5TpGYANf
VgQRIPeli4o58XxGJnNLAlhanOSirnQt8yFoCrza/QPcwrd+UX+jTqYarQ2HLS2n
4jm94EjbUdhm/X65ZOg5DIcXHWTTZ4kE1hVLgoH8M6eHfKva0mR0jMnKpU3+/xEk
RfXqKjiSiQ2xvqfrJHx1s+vRj7he25mwCsp9XEF+ePWiP/HinuYWETk05JmrZq4M
2QwZBEi2mosYQN8zmLx9ZUxCwmN2CvNwO6FbcFj7c8f37ZAeWYMZ7W5wo940TZJd
OksbyVke7EUWyW8enS6SXXL8M4hBua2hLR6Ba9AVUHHULBbvXPMB0pVx75yFJIRD
oCQaPGYiHH9BBzs3LT/acsvcnQ760f65VpFuD3BphcVtYwPhsd0Z6jsmktlKywUR
QQRNkH6HZyBJ3N+/kkNNQi9Ho/tPcVPqJfgbyA+Rs0B8GJrou0w2XLWo2bKjsdYW
V9YlW+z4hjo41hWBKA9MEgMnC8QrJ3bab9G9e6b2BYrzUSod4J0L4tuU3/cuyQA8
92FgNo7Ua2lAK3GQstd4J5QMADsIJgFK7D8iC39Kp486pUwJC+Cz87L5IlcVUJYy
f+4QSegaCtonK574Q0sg3+4CZoN43E41msIEOovzUaLHw+Zey1CXj+Ei4j3TDEet
yZ7qB6aBrGOZMMIxBES8tCgIW0u+53ID5YNMB/hSY9xHX+YsaB2rjGpgjXfqMrJo
VhxL24M0Kpvm+OKrDD8qvIe0T6Yx7GTHLFhzehHF2wgvdhw19gDYrrs2vwKf0/xB
JKLa3APYkZOobSsvBofxLbRbrczEK0NGp2XjWrYziwybcCZBv/CDPRJYsyNqZgow
n60y+zzSLbi2e6nVnfTR/eop7PO8yzJB4lNwLZnmFPZjsPQZw8w+Wz2d7G+D/xKn
6FE5VJjjydUvPajaqjr4AOWIyZJx5KjtH5zr2FjPTixI0qCH0SRuouLJ3fF4sPVz
dArzlffeq4eLFCmTDLnBJhk2mLEXI9soAug3OymcqYQV/ZRhsRb5wRPuraXq6hzw
ynMRK7n3otlOBA7IYXVX9AOJop5lYF/wVU9CXKzdWHZ1ZKGOVLEWSDXUSC0pIy+J
Chblhj3xm7KqDT7Ce6cve5VNm7tnNDHZ7ZgVUY8VcdjmSPctRgK01Y86JmWn6w+5
Eq0T5YZpynJfNS/pWJXIt6DG/9uSkQSTv+T0cPs0du4jrvUkJACma6YxZvtBoc/E
RXxfhEN3XrbpYPY/tiiygimfmbuQyfCC4vyATuvSZ5neY7wL9ZZLrGrAFSYJCMKS
6muC3KEWDpqSqPGUENfcA/7j6ZvkY3T7W0OgJMXLMy2kwdHAbOX9FRwxsm3lnj8i
AErc4MVyzZuplnr4B0hCav9sBkM/HFs1MWEqILTiWi4iAxJ9AJTtg/DDjt72capJ
13UCoyl0YiOjvkAdyIQoO72+wycgpZE9w8f/4pEQIjZk+XVq3+3ojrd+Cnqe3CGQ
1a+VU64NtOxDz5QlaTMNTNrmfPL/T+a/OwyYGYIP891yesORj5IAnPFwv5IEuBrb
55ZD4qPi9MmNqRZhWn22ngxlqHO28NmJfYpVJwd6f6PG35eyMg7V5d2zAKlkssLA
lc0wuX61EIBMlWKvQGX0MUzZSw9K2JfBIMEnOMIA5Ow5cL0F2ih1LKeLmK2QWgpV
63+yVWBtXC9oGF0AXIdmq/jYqPboVYDfkfdFSBCfmObqH6FBUbmg7jO2McCg99y4
FOZuEk6+DQxgGkVa1N7jImEWIQTgASfb+g59O0eTvY488fA0znJqTJeJGZ2KWMGQ
/5Vvtwxw14GxvEBYtPilpHuN8HicoHeXRZbfD53xpdtYWdcD4x/HKLShJA929cUV
/tacd8t+81Qt6RYVjABlGCI5MFJGaKtp1uLAxkARpqc8JbDZpx65x0QBgOkBRzRq
mRiRXWFTijDlJ7zRwpyeim1lN9JH9mBBSsVHT6lt9qc2igD6Dtg9yGoOsp4B8Eh3
CNCYnTI7rCGphlhQKq9/ssdf8G+czAqjchrLYqXyPmtmiuHBQOzTdlOYDsztpCne
xNlV89LokunxjL3hu+CjbL5ilFdiB1GZgvDPQ8dh/3C7Z6Xkzg/e44cL4JTKFxEY
KsJlt/8k5kr2zyUHIRQggwLtBS34s8p4gwnTjbuRghZX1DcPCOAbOXG7LLXuEwRA
ZSje2B4sR+WFdzyhF2yZbggr0MHpJqAYkxbAUlx9F78Kx1hjHMGnMzxjlazXNpG2
K4KECIexPU4caqtc2AHZ7t7QmnpGfqzcbO8qPNoWR0lJG0Qf13PRIFOIhtvi2rl2
FtDSNEzuyVdWd+wV4sWBWLIv2QGzww34zvvecujRSMdEOksIJSLQ1MIYguq1ZZUQ
CkFs/1hZdSs24JzhLDTbSEsmeIc7S44loxGYpjVmoneDXOCcx4fz8CyAHRa9n2+d
RAx8gsPtvZTojq3mugT1C404/i28x8rgxoLqt0vkvm1eDgWiZ1NMq8r7t5VDgy4K
9dBbA8LQvSUDDrq4BQDn9kPe6vtRPTr8WvsyPHro0FQIsXJamvpXNTbwwy6EeWoW
fXR52+MloNU32IVhpZamyZ+wYUk4Jq+qzO/EIhRzmrw8LHzUSJcUXtQIxY1GF4yI
PAEJf+Hkvon/N9FYh/W4oXKJRIW/DuBURocV+caOA7E0NZPpguVz/UAqefHQfI7N
j0wsjEqpZUz7suHu2MG//3Z5SZUIBdRnTfxzfNdWl0AgRQaM4l2M8VLRgpTavOto
EbvWO9w0atNHYVxdxJRfHVGkkIGwwEKD38uQdDhVWAhBOD1csfup7W4DcYfnTmke
GVXQ5t0blZiLeavhRM10niibkbzG482J65fID/m//f/cuXl3OG77v84HtGHwy/DA
8Fpq7lMvLRN3UPjiis+QyB1+0DHUBbxf8z9cpvI70aA3lqXaBOyof7Xmb3c5vm6f
dU857WuTvQ2OnrsmksAIqSau9cTmJfojO1IKW42lVgtLIcBf+HkQUTjj1bjPP1HJ
5fSSWyfM7MSabHkFMkBlBeaMhMWCO6AL0qjW1HJ0naMldmpeOWmzU59c/kyeH1Hh
SvbM95Ke7n3T7fVxrP+NtGO+bjjVoZZ1BzlyotIOybIlDj3TgFcDergg4iZwti+v
3s+MkdBXQ1VgX0kuzkEx7D3dCDVvkGGG8pzZw8E2Z4Yt68AZU9+4FwNDGP/utPZ/
seU+JZsPQPDrgw5eGbSCM34hsiVpnvRe7bWBL91gegD2cozOeqeUgF+ed42jgUc8
p602cYUeQYJSTYuk75K7TdR1FGvk7JB4h0SnbwcVWjTnz0XEDBsq+raYxV3PtMNU
kY8y14JTF3h7YBOpOlohcN9iDARKR+Vtd8oCFSKBRNRKTi8o/MDoONY1CBR4PLTJ
swzdSg1mKQfG7rS5LhS9NloexLJ2RVny9d0aXZAjkCgQsOgfrhc8/2xeayiSP4Ro
0hBUdsNnbT7NIWLdLZq/Dv5OCQoqe89eIjSIQKY/trFUGAqqqZMXpZV3bXR5bWpi
K1YFxKRU54fE7mWyc9JUPq/S1rnUNNnFA3iPihTERulnG7lFg9OsEpF+9WbOpz4C
vld522VmSUw+aYF3WT+UtDjsiWTFgj6SHSkg1QlZF2zFIGcejLTPaqgIMBt46k+U
LSS9dxd8i99jmNPxVBwzeAgTZkoFDL8Ef9LAoTSSmiYRnFycbYbE5PAEkR1m3Slm
d2kX2YvUHUSji/MvMLcBuspxyj2KOz+nD1v+VnwhvFZuwD5evqK+p6L6i1nORBm3
1kRmfewOnLsHWiq3HyxEgw/ovqi+yD080mP8i5NqffQ9o6W3DACUG7JWpqp3/0H/
7jGiSMOvcDVl6CXJwTmT4SDDGML5crJLduBZwYMUAjaBkBDigW/y6D26xtL/UBUj
uxR3ZR2EEuF4jFH5eh5IqywCbjsGZzEIL9QA35skmDd83qrWYeoz6fCLazDIEJC5
vWGqfOw2/8aRC0P8/HpsIlvLKVV/PT6vOVLIMm+9oJPMobZ7TjAg6JZubbgsqQ7F
qqeePCrYZQa62H9LS930IRgiOl7JcUjt01vmw4wz8KVBg08Yrcp1QQzTNO4WyyjA
Svu5jMep+JEhca7AogWh213a0d+3/8i0TJOm5F7+MnqQxBYozDUVigUbI1U9Wk3F
TFvZ9qUvfPQbdPjExeBdvSTPcdnKUAH33rRUSSyGzme8IaqPkxOlpwt0BkjaXELB
06AsVYkIerWPaoPglAqFrBwqbqtr5kw3rlqxYPtW5U0AOy/S0ioxAVBCP1MqGRfO
1V3RR1H6vxVmJKudfCDD3UYDIovov0TkOk7ScbX/juifnKBgsu10qp3vP2O+w9dQ
zkkxgUKjaHY2JIkab62yig9QYQuS5xHA+WhvY4L3AKIwy5bGM8s2n9OQXN8Zi0SZ
U2AvHJc1lCEWjlhUT9bRIXzJtyaaRP0eluheJ0m0GILdvFlg2x/zHwXxBzGMr3mT
2WYNnDIxbWeDGc972xE7TAw+4f7+NgUSnh8xSGTTn8Td4DfTXFRrAWyre622Eoh0
E7C95SpvabPCFgZRtntE/OtRyKmBl4c7NPfhWwMeLmg2/K1OC8RJK6iVKJIA+p16
hfEMnjyUtnh8zYukakkAI5VdzZSn4DQM2xdgCZcMrUXlSSUjNyH3NL4xcqveuHSG
GVOQo9E0+Vu3P3BPhysc0OgpzEBcPWL+pMBXmxtJYRCqTVwFmTAb/1DUug7o0FLS
j9BmQHrEctvKfLHWhHe1/7roS5uEoiqT7mWHKb9wjF2e5TZmn1RQaFj8aMT6E7JG
J7KDe2GxN+Rg0t2A9fCf58KIXesjuD/m2GPskxDXuoUKvAyhk2Xgceyj7Om2+4kS
QaqZO+gOLcmepSUg0+Y+C3UnKl972F8u1uudm7DKrSBye8Nhw2YwjKDL+3CQy6u7
wXtrrh4+YkF24wgM7UTTtvLsjk4hsudge9oo3BleWB7mnfyu26CQQl1CdCaqU3r1
hfig0AuhlaIPoUhhun8S7u5JpiN3MMSiGUWt7hRiJAzCnZxpmW7rGCZOg8aTMFNB
Oa2IXWLroYMz4bfj6lohgROncGQkaPvfwCkaDhRkuKE/lq5nQQ4JHvEorGwNOlhV
SUeCQ2/B7PpmjAuUmYGwZo3uXmDSqZbQPr3CIzySxw728fC2v0N5Uutz2iRjVIfo
eQU++djIKNKVaqGfhzrll4oRua6biiJfXNbSmV2keuAheDadQux+tPZAWtUC0txj
sKN/5g64dBbzeGQXXkE7yPhbqYjJXWKMCfwONow6wGJ+jgSoXipAm720XfX8U9Eb
tCiw51drHkIOhe/qEa8V/+90zHUYYeuSO8GKNzs6XhxSDseiA4qlOtEZTNxf5F9I
4EcFIB/byd49cu60rL5YTMIWJo0CqNjmkj90jIXsXHkacGRGg/hrWqJ144IgjmXg
XssocKe2TawHETbP38Nly2sDkMmmPA6Isq8Ijp5KsrLwNK9XhmUOHYoSshCiSZzj
RMRbqaSzJUPTeyHZfv6ofrbkLZPUrF/IT1wg2oe/XD6jk2judLjCVlzpOJ+OiE22
xhgoglepO5vkZlbxw0BC49fUDAhYoF5a03d4ExKRXfWO/LOr+wJ0Kwov8ierT85g
ZJN+KA1jEe+LSRuz1+xrHG5gIX7QqzJSFVf4o3RYKln8HDYZ24pxhE6ktqJwhQke
bl5BT0/1Pik6S8nCcMYXx3W5NNQg1fmfC6nTIO/zesPii84t1vxEBqhPEBc3tHGz
FJw149kIb/J77QhsyBMn9oeApZRe0B/uu04Q8PozYGb7OiBPO+/wC8m+qlrhrUgl
PlPwUhFr0i1kwko2qP2zjoZ7uzQX0ttA4Fpkynqu5pw/4M81IhGbThlQbmy5VL77
z+526nrBiD2b17SM3NQujHt7XHQaP0AsVWrN+F2mW98i6C2ow0vbbDT2NvESy8/q
cM591v1iZHq2oepI5q2JQfCUg3Mmk7vGd6qRS4adJ+r9QxwGfRrNGUX7HN0B2QRg
ka3PuZHuIrYenFL3NR+NkZU3g6M/TZBkPlY69o5as+My+CuVLyhibmPDnhfAEuiu
9RpmqmbcJJYhhcGSNAzY5YcCv68ONGGGtgBWbQ5caZKA7tT3mf2iA7RsKh36I28V
AmQE7WaI4+O8hiaAtv0VvcreDzPSz0yJ+a5QYKUZ1Vbg/xWX7oYRSn31F+LHNN4E
xEd1wiyTw9mD1IM1JoR/XExscpT0mvbc/Pf43lLLzd76KnKMhtQLQRm6ttaEyg6T
7q329o/hgqhcPU6Qyov9tTppwG9YrBJSNeGz0wi7ALRXw10ilPESJ6G8cRbHyDHQ
L7eHYjC4zBRvj/QJbmVH64dsEfzC871CgZuk93sGY4DDZQcMfjX+x7nq41i4Zocd
gp6Lq2czVBwl18t09j5rnwgcKAKrrCKtC3L2nXK8nQOs16wS0+Y5lLgmoK5K14zN
V7oFWJGkjq1cNQq4/Hl+JJQChM6ezHAvHOYpsNkkmQUsJMrjV5+key0x0Qgl19Ui
1SNj5eUjjp5tAq/mGdbzVL1NSCWA/B7h3OdffdfF327UyvF6F0sS4NHV9sB78d58
JNfuO6OvQXFE/kf0PCGcEda7ShWWC+Sw4FOYPV5G/TcEP+/tNSLP3BOm1pAdL9DY
MQ51eR4LIWFbQo8vXjlRylYGxI9QkaufEZovE1UD/1ZhBYOpqUUKyrBTerx43pQt
8BQe+IIJGh+A47WzyAfVXKxYKAJ1SBF30BTqUt7C8JHFHt1KZwQI7K+35aiD/HsO
g5IMQTwDWfriJ8MVIGqgt6xZgtoNjOBLbZW9guEa2fcHIEG34/sAcFTZYrGkaypj
d4ox2dY4x/hyCqsF5gXlQFWUxSRx5IkOjCe1lLsMcImBgXBYVibVc8T32kvjChSr
zAFElyg/AniuV+jBdOLSsVE6PcamGe0KCkPqyjjlcF3eiQMv5SuK/jS4SwqfxmKA
PdrXEvEK22qz9lwo9AuiYNv6L7ETfRvAwnzOclsR+E+p/7Q8lpgyWJyKXRkPq0pr
co+2krAYQqejLR8HEEBMMwESFvGDaIfJNmuNjkxcRoQ0WeCq0183MLp7sirofIjF
q26hpd/QSQlqFm5kkvGa1dbEKkzFTa+thlEztr0Df+0hjTYZma+w5LCocCu/Yat1
cd5fzWV9D4mZgRnbpBzIw6n2rMiRBPEJcU6AJplThyoWpb1S/mUXjVZPQFUdVi9E
PS6Tlk7dk+VnUTzfMF+lZMsg0L3e0vAaDgFf1HHotXUYMOdneAqvz1WE5x0L9UkK
GztdRz3OfC49vrF/o9EiKRaoEok7lIllyZ6PxiMzK4lZ84k06fmK5oxg/6m8j8cr
Eu31Aqtjaj42PIESb64a9u381YZn1oA6BVaX0DN00+t8uUT8ICScgC6B+dou38KY
iIOUpZR5ZycYNiZdPtO3Atrj6vDCv+t96a4RJ8Fk0OM9vrJ5kIyNrEhJu4M3aWy7
mLBU4WHJN46caz+74kbgScoRNgN+n/r1IZH9OTRJrmIwKS/1nTtMHoqq/pMVZJEu
DGjV+86Yqc6jn687QbfszHUayGqF7wkU0LWghyMMSmSMrJOiZ0vfX7FJTTicGZqs
/Yg4q0GcC8KQKLf0+8IQ3q4PuUnwwCmLmLHUiVeoScukkrLFbCq3Kn8UQxRyiIN+
Di/pt40As8P5e+Yjq/cRJqN/xMUzaD4wVG3dFu7IQyfRU8sJ9mUAMta1UqYsdjfI
NlKeFDCIenB3QZK1+PKL6b5Lx7k0mlkhSQ1v3m15zBbCmdNJ98zD0LLvQelozS+b
usz8mFjk7+VV2LpuNXVkajJyG/DSjFX3pp6lqo1kXiEmIcrgdlnw1Si3NdN39dpB
Gz1iaDHPyIVplylagv73SfuzcD3e28o6vBJGkaCqMZCJoHrr0zEp/gA7nN25vCoT
5RbVB8O7FIjle63S+D9u0FdIwqOGmyIW5i8/xjz5fWg0ZaCxRMaSr3VITZDw2klF
ScqEJzsTzYhNT2T4eszLxmLA3oremrtAwUKchB8Fo7hiM2OfTrx+vUptVPn0+MnU
ac3D26/iudh0gMnSpvFjKfumgzoB9TDn+nJMP8uXzbR9PHnuM+mvp83JJT8hE13h
VxaxUMPKInx6RVGpFGSAR8qJ/D/FoAm/y4P3bFp/t/7qWocRs0pUGv1l5Yh5rZ7z
Jx0u5WaogNLK3BYZiipeizonLXdczYVr5xitmJ1w8v8c4B0gBtNs0nZCBJ37q2sc
owQKqKIjlEgP2JpgBN/Bieb6w3YkdtdPK0KvHdZoSqPtUsfq8+n3DCcP05wUKNUx
JpH2NfWhJ8IM/cP2MReuKHpxgYX4jNr63V2lWe/jan3A+eY7/fLW5/VS4M6zG+Or
EcGhptw8W9R7EfjZsujtMT2yMDPH522IO8oOdHWOjqAjmPx5V51pa9z+p2RkXS+P
RFJLH222K4MB6sMNv3c9v+ljNSvjG9VX+7xELdIAn7hFvNwIbJ5Ruxno/fgq3BnP
0/rqPlTCl0t1LjpHoPa3C3m0JChRVfmHZp2VqsSZaw7MqFrounK38oo+lbUfhFoc
i88WoDmWcsVDXnhkZiiKUndxOmceH+uz8DeZ8skcg7XeXeliPFiOIhAe57naLHhf
sYteYUap+oYETUA2S2olGVdFX95HKtC5Q5jkCzVg9f78H35iyucHdKexHPmex8l5
hPS1WWPxkU4JMVuKUAeeWsKOgMrADjZUGmTqBwKfzTL4DZtd35V3smBxw1KNT/T5
ix0nKvR8zeoc/fgZFuiP0CgkACgu0nBjHd9wNRsh21R25G8/wc5EWm9lP2Gs9UiK
C4/XH4QUZ2DmOSU/XX6AjPm/q6T9ujQ1Ydru4/bicU1LbmHzzB11cwIVCHX0HbNE
zmi4Mn48PqROzGIoNTr8VuJVCqkzPu1hX0n8EXdm/a+uJE/JcJby4proYo4rPYNl
ag6F2JMSxT0kO6RzlNbywG7yzQqpcDJ0EOORe1E+8DsCea4/LEJxP+jZ+l3gBld7
Z8BUSaz6BfTSJXVAKMubSbPkPHsWxefF217gOHDLHrxKenDg1h7Ql1qA9MBAfK8e
pE7ApivEKEkIob/TEcqjQ3DCKc+16/ySzrPfrcCvU2h9VskNNcAN6TkSvB2hZsuF
17NGkUA3e+nI+9xrSLVP3tPa6iGJDad5ltgPgrCbIFsx9SK8aCxkZE74xHfnkSTI
Ud6nsnMnaeCrRQf7MDdnmhH/s9um1LRz5k1YFceDXzIlfAYd1p2a7wf5/Verd6zX
LCqytUXa1tt0YWKS0fAuDtlQ5btTVWRGFCsnZiAsoFEnkZygx+4GBWpzJ5kLeYyo
v4tRRthFcHDra+hBesHiR5CYsADPN+nb34zvtcp6BIsTkDvRji1jM0AYuY+O/oTJ
8oXHLWFO3gfsi5M9+/VyKp7hYCZp9HLw0SFWgJarkXeRXXlyprts095Aq/BU6KDU
4ulMNeDwgtAHwFROKgeQ9tb61NdSBql2HqWMNS6wvdSliyocPctP+3TycpsEDGh5
A5sZqHXbtwSP0I9aDfw99wCURlG+j+88Pty+Q58UZ+D2NkOSrzqIgG66POhStgfQ
lVR4qNN2c3CkFULh5ysmkE5Oc8JBDL6dPoqORhy2alHGej0rTqHTvZj4ctRFwqa2
DQjp8OmoUJ9vTUl6skIyWFE+Qchzg9i47n3iADOyB7XyxjOQ7QhEdupm9ucKH7/9
/i47V/l3KmWlOnEAaYYia2NhPnvdL5djHYX09Z4tlWA3fAFvyNQ9tI6v2d89a+D8
yM21RzfWDFHMrG1vToHR6ruCvPOKf7Dx2fHPwVIEurln8GlA9jz6jtby30KqqJYA
fu2bkBnvJWK2o9TPpzZiQmuTmvvDcamw2Uc7FIaJpdQaJvLEMUWqjVa9sLiDKjjj
Xu89dd07NYKRcyDrv1Hz36UXMHKEas+f4DJwTKPp3BtRGJ3gSCKL32qXC2dtS78Z
V4Y4aBnY06ywN3uU5Ake5vXZDoB/QD3KvtR1T90QkNUqDktFGYAEWRsiri5zd43s
q/FF5BtvephfY23BQxqvlTzPAq/pi3wptzkzDjRVzbyTI/VuiYmtdU+C3WsjBSfB
GcR5UPJvn2UYrB688MhNB+yhpZ7/4CMv8AS2QE4iKcr34YUDgsl7Y2KKJzLlvWvu
6udnzolYEhDJX+u41b6JCVts9hr4UB7rF7CORY0yqhUNTnk5/v04SkESqyexMhO+
bOr33+NmqWRTyvJR+4xlFwIoETbpOi85i/Li9i8WhWFIFqglBzRYwLpx17/xyFr0
jz9/1ccxSqtGX/rTo+CXqZ2lZsGbBouirvm2OGp/0wvFCmabEoiMZLJtKRmzKYRR
P9LYal/o1kvtejgQ/2gFAOGloq9Lzh7iOFAA/Ss/pDsUGxW4TQ4X4qrJ4SyTtx/5
UQpxcYFddZXKoc6G6mhbBzlJwkMZoPce0roT9+y55jwFhIX6PgUvTHjU4BQ4C15i
ePWnNjz/caXxpoqM82/8mqcUoFvqLmK/gnC+RV9EIMWxnBGMD58tpZ5y48ZZ7Hdz
2QJb3s2WjrOKTxUf4MlpSqLt93frGF8L2D9rwnQrfO2u45xxy9GF0cUSuxyj+Af/
5CfSDqM4p53jgdBH59/4kM7EsGC6e1lrFKOVO0bwzxOl+rKazqvKP5sqixptbecW
Lxtfsvux3DcGrH98cCtyszHxEtxVph+LK64r50fsimeJu7p5J90a44Uy0QwNTlQI
duvq6F5NSnGxlItWrjkw0L+elB+9jmNTLftDcPMhByaEjgWEALC/7K38rWw7Y9iF
Kn4ynhT+oWyd7VXqCumUjlhXAVCXywyihH5qhcRx9J/kCccDfDbGzOUdw65zB3a6
LfyIT9WxSiRIMaXDlJmeffmu7PEyKzjp9xhni270LeKZZAf1SvitdkBAr9YcaJe2
poUWn8/H0FCD6OESrVrmHhJYmrOn1bfQ/brDn4+/THsNKo847EyrRHHbsHvxyFcl
Nwtwnsesh/lxCZTTeLL0CRBMAJCas7kvJSSoM9ix88E+fscA+iOXfUe50ehgwR4Z
OdZfRNUUuQLT4g8fGgPbVf18bBTAbWn7WOMzjUs2cmLUJygnGGANpmKlcNCJsZrR
FmVlTdDbLRQdblaRhxJox+1eW6HM5RtDLvdrSeINECJ5bEraGKG+Gl7siFWnGyoE
2k3tPTJCIl29TWj+CLtKouKEB3UFJMAOdicZmJwOeYlyJSUPELQV+D6um5On8M3g
dBV/zdPmfqxxoIGbxGKmTIkrZYypkvpfaKEbbo0Wsyqrgxw/3tE4UQZj1+suHfIR
clG7WOXb2WmY/ARuRTIswzcv/q2qJH/wqmysybMXS7kbQHnD/CvzMOZ0A0E7HyYj
r02F9ar5/tivExdCZAUstFME1IaYYkhXbYfgyPmBtY76giX/U3FltluMKlvwJUtE
wabm2+RuYWNMqPHW4upJmkiY2/YnrSHe/qMZhUUAhatqcquYCdNyRrqe9cEMoWim
xyUpKP5/ohFby51pIMdo9PzL8+VvBh4ClH3dpMNHvPcUDWNlnoz2tyz1im3o2niA
1lOAw54h7CKqhDzqeyszyIuEX0kfeRRxA0SK7RMGOTUbA46mPxunfk0iPFQCsBk1
wNaVtDBTanThfjW3ec6sxzJMvOAtJuWhlcfgjbKe+XyqW3nRkOAPFoAaPNeU02OA
aJTgDHmoJvWmYXkuNLSgbDqUAZCNgMk3G88Txjwa7UZcltWQHTX8zBvphWJ6xswW
M4XkGaPSuJpzVcv+ClguUna0PssgoUnnkGX/Hq48x+ufWBfapsr50i/HHodgaH12
FORolsIXLcaesnHF3P59Z8yDXEcwPNg9d3s+J8gPY7jd2veicF3DLDjUOdd2A2Y3
NAretxcU83xPDe+Q3GvL/BSjObvNzgioNW/6sCEmryMeeHu+CX14gJ8M1ndhCWLe
9lRgdLqVxt/62ArBYHUPKZWxZEq+IU+3nGWIgsexlx4esxjFDeeL+CqNdlQCjICH
XUHJhvo9Xj7/DuZDbKdDvf2z2tQFW1dD4T9Ac3my/nlHhbNLpgrGgxKxlp+PEj2n
uwK6zX763WwUYpCRakAOfJxNJSBPxAXxwOrLS9ass5qyiuZrP5+zETNNvPLwFHij
SVz+F1QJh0aEckaYuDYN7DULbX0dmtg8lQ6wFrUqf4qSI8zEPR55qtDhM4Vqt8Fu
pRhluqlz3J7+xrwrRkEUikaR7V1h9uxg5pE0ZTVb+7bDFW+2krjQEzMsroMBBrRh
3pxVvSNrxwourJgTCs1eesAS0JWmMPg2hstNUNy7Puju6XhUV9l+5kV83lO5XFl0
ff9BuWEyzgjx5ODym0g6UCMm1NDCl+LTZlz2HfqbqTec4AsW1MzF4tMsWFYsOWv6
gYa/ONWGQgQAxGmGAakPkPoWlWVeIWSBTuGGPUZIyAawNkrRceI6u4AubXgc051N
UTuVjw/kZN9TSGUF/zLys2oX/4IHvIReH3N6NVVsLINyplcYXruVeyuy+gqxesPn
VFCRoDmM/oegTe7b3BAzEiw4esFo0bd7KH2oAob70BevPsqyBAUqifS4acC798mG
YXYYnEe8chYVFHGo4g9wYN4Q5Tpi5J3V+ORmxTEHHRTcTpnUkTj0wmue6AL8WKA4
qJ/wFK1V76q5SdwGrVTsoxsMIiOhg9zGG3VfsgPN6wEMMDZk1gS9NLKBDLWcqgv5
hSQnbErVhAL70PhWdfTo+29ySDvkpQEzW/iC7qrX5tyWA1Zz3ZIc3qF/fz2cUuZe
uW66XOdHu8WryF4vQM5ZaHZf05MM9qDorviBRcwXJQiHiT7FUx3AEC3wDr2D+MvH
YcMZMFaavfXFHCOCI5U1miiAV1zX3IRGChJbcyysk4HI9NJF/8wdFovX3j6DlVcp
RLLQl8iTop4p9P5jlG+RB2QULCy3BNhKWeCxfVOY4ehPZa+6g8SDA8tkjrryanEi
aXIlG+Uk73w8XTbTfshSg+47X1GUTkNSPsyBqmrSJ0k2tXKxN5iRptHTMitu0nnt
Sa7VQkXEReqJxdqJBZNGxE9TxaezJvDxd5HM5yUUXL8+NRplNtCM2AtXEhlezUGX
LLdVhohp8rPGjAL5U4fsu9sZiFg9FVMZIgF92+DWqbZnRklaO5pRhtwi0pODnNr8
FIgHLKEq07zx7uS8PbVGHBflwU/NAHgnd+TmbW8b3ISKSe09Q9vAKXB73zQkFW0w
+wgdVwOZA8MiSDsfPpbType9PM2VYIKHjnbdllYBx9BMvP8t209heG8y5Ei/sSAr
VsNaf9nz/diO3nh7ns4np1z+vOnBis+Vvx/CLJa3J3ldSs6lDZT309l04VRQ4WEE
5EDrAoyGY28d9HSWK7eXlOTatVcNeVgFLf/QgZfBXi5MbwAbtfaMpB1WxyTbZK9a
Y6u0x8S76Ef/bpCvQu4zbHQ0jZIZcP9BiPHnd2+Jx40IYi9phitqQi9v+k+lln9n
VL1kstF27rZz8StIuxVjNXO3gTzE1tYn1lpmfdh8XNfa3dQVsSme4HxtZD0EafI5
QXL2Rky+z5Ch3e5scSOZGz5jCgzEZaajLzPcDA5APoYUhDAZQ73ELFvOl7fYXsN4
9ac6RTephLxugQ/3y2EF8UOSaaAGC7YdGs2TLwU5wm299qE3hlQXhCwx/bYNyUKb
FPb0exryMOoANxQ/a03MM7KLRt3vJaEi3h7r9EO8sdmrxW0FOW4PpjjgNQbhbvJG
qQ6ZM2/pwQcorFQQlZ67RqhHLRXxAydQ48El0DtLW5/1YlWW4Pa7fciEjFqKyqmN
6VHmtBei/xaSKW+wdupI6/DA89C0lJ854HlWYSYvBTNBIt/L1EXT8UNo9chB8Yo3
1j1liMs5tKZoe4xV0dGYfMaTreLvpQLcQEPJulTzQxwlxTS+SFa/akB5uJzJrnRS
WKkEOx0B3aLCsWhJnFLu2zSXZcFOxfGmSx5zNfX5W+hKZbqEsSl3h3v6PEh69bvt
uj6BXR6GZi5T7kV+yQFiwvowmstWB929aDU6Jcjzyz5/tV8BTMQnrtXK+yLN5uKO
qeXVZhjm6BklSomsRORPvAwvgWQEl+sQlYTk4lIZtwnR4dJgh+IlyM9nt0Z/BWsW
L1BXG243l8OqOKOAbLDsEQNglNap3sD0xBqKcagW7px2g44HHrVVBDqGOLMuhJeq
sJIrDUwT/iJU8aZfk2jSc7AtPdhOVx4piIYRPhkzGdyI9F8LBkFTAk6qiVyCPjEX
uQ8tAZ+fHoa/YYBmpo/geq8Y12dYDf0ICHAV6KU7m517J9GuS0enBLRq6b7tvDf2
ABRtgNFAx49EAyuyLT4h0faqmoTru2IGA7+1kxH7zXA/pAEHLTJ5+GgNAc+z4ZSd
jTxyXMDcxCp2crzX3XEppmxuf/hP+UUuFvO+oUa+kQu3jsLLqGD0lyCTItb3QayZ
ehpjwdL014iKATrwXITIKJOpRAdo/CDwE920P5VubRzKxZYomcNfJ/qmutk7Insv
dfN5Uf8vrONFwrXThnRZXQDx0Y9U2leBTLLLziO/YjR76KqgTderG+e5ShZTvPU5
tOewZcVnnVxw4Gzw7xxJNLSyWHJgvgVO7fhlHGQQFSoNheQpsNaWoLEeL8OmTtP4
AJCnPSTGSvSmv2Bg0CUpqMhHXwvIsc+yRmbsKPOZGfuqoEo3EsRSz194E6UArgfp
y//oogg06bHfz1P5+72bfTqKvuh/a78LTsaejKZWKis14kzMw4H/gHkjIbT6Uv7o
QwwSnGKH5DcOp9a/bRYtiklUqFxWbcnxwx/9r15+AqTlo2NI9bUSHxnk775e+fxH
zTHtLrDmi9ArZuX3fduxMQYo0KOO+QPYKjOO/d04/S3i8AlsYKFiG8QKoqdgSjkI
YJcn3ET+KMySYnhqe5ejrKnDtbrEDRWlGRXAPwpGGuf+L5VJxH+XYWmDW6vX62cB
9m/XYyaVNt7G+QcsHt4qBMsk7vDG/fR+pMdRRvxHa3lwDZynokB9Uxk3iqfsjiXL
aw0Jesgx21ClebhyQkRS+1FUJ2ZEac4j1cWoilHC4X9ma2lTJ5amdktd/+ntpump
3li3nLn0t/nTSDaBQ3kKWkSksqSJNvgk0WQynRJBoCi86jA9WCXCu+aXj4uS3cRq
IrSdaAMaS+3frwV5xCc7nv2NnzhXj2WUautzBk3pY5BiHXItU35c5I3W1JfCWtMr
gyvGor4P050yrT5M6cXhwEF65B14LpzouEruIWbTndTU4qpQsRt0Citul+UvBs8N
Spdq6gPA4DSiV2PC39Sniwicp3b2ImQ7531Bz7cdWiyBoPCEUC9YtBYZvjfRv+Pk
HFcSypMezFv30DSxYc8hDhY30qlykJlQna/FGpAJymK6gXx6s2wecbKKRkauIykn
+/87ngb6pOz14YTeucN7WHmYvxWlspnei8WV9LTOIQqufZK9szJU3lKwnQ+dmRH1
5vXxkIjDaZbOeOLnlN+fbkgjifoG1/VdNbXd/f+OYauWWtBHkkNcmi4v1lQOvCRj
loP40T6iPezys/CTvX5DzlkJM5IAbKGaE0L/9yEIrM9fDIKAA5/7jIIgLxD/Uu3s
9RU6OA/74HauQTfgwMJCKPPcQ8XlqS9LK9t95ynk4MZqfskjJFaW3IW6kkLUBfCK
veaw3998P/mqehMHzXIWpXsMTnjqlKImtNuoRwjclufE5XY9RNV0q4zx0w88NyMx
xvz4ApyPbCyo4NaBTUIejrB7dSF3rzcAYVoyD+JJVMkVKZTRvi4/B0Co1EL1hglc
P1Nqdgd92V2WNkOnOPuwfyBQ63Tlj3CGns18hZ/cx+gfi87JH+4Yt/mMKmX/QZqp
Bf/ey6uRGGgSmLhFD8WMifKiny/Ifn+uGqQMmk6EIV2vrZ2Msg0JtJWXGkM6VZY3
BsP1hM2cyBP9ZBZBxLpHiA6rMhdJFrO9yVSn9uqP0J32aY16jfceaD0dTp0yZYn9
UvfDMhD7NeCtuMtY4WFUZ2Lawo/jQ4evdAOcmebXyLqun2eZGbw8pmqq65QD/vMa
XmmG724r/J3eEDYmTDcDSFWi2kMgRq+lR3HE4ifwVxZfw/peTM0mcU0YzuNj3AQF
70iYKkRnE86I0zuuZyIBjlxUUyU2ZN/V99mhY6iyXi30aMoH0bOq0vFoojPXgUMj
h03FWzyxBW7LD+kOE/GrSDKoUUudd9lpB6/EFpbHIoi0Ekse/1T4AczoTn2Y31hI
BAmc7wihtHy2Ah/JdW4iALwS+pUVzBBSJsynPMujHnaDbQL3dq7AM76T9SRjgYcH
ltOy0OucDzjasySYnS4UvJeRmAcjKeyk7QcuEzQmzv1NpgikYajQbrTZ6/tOqti+
3E51Pl/UeY7sIBvcqZydBEI2Q6iL+kzHIzazLlPISwVrkTygVOy10w7WGzqBuQ8K
f77Firff/g63VzB3ZyO8GhShR60W5gpOikIsFUgxW8wjGFHSk7aIWC/0pnWToXZH
5CqeQbf8ff9Q+sQgKdUoT8KkVrAPJ/mUSwMdiduhUDrP7vbLXp8kit87t3hzO8Th
M5Jgaj61awF465YqMuht3I2ZabyDK1zO1ZHrnlpeN368rjCs3EnWxuXMBwOT6Xc9
XmmVUjx8DuKiYIQkN4LxXUOX99Y4TG/ey8u2gweFh6SYiDmp6sislHu2V0zTBfCe
vb3UULepwiscQ6NIrGKn10lHos+g0TMSLER90frYyYDHtvP8ZRkp6YQez/HL4++T
i3FmClbWq+kItsrcXAdoQRs8g6W0FpRlYCPgnDMd9ArM6FhwzwCzRIpDNyGDM13i
xzM5JoJwlQXjK1xkvK+8BPIKMr4ktomWx7+UF2+WB905UizHscSYfS3/VTnYJ6qf
lI6Z3mDfATSqyrghZ0At3vYI1TlHtuZJ9tdnVmkznklVPkUgulYzIjfOBgoCGzWn
sbIKuQKfACvBBHSuUXaekw0MWasiTNyVm2lTpZuYPzUXA2wUDJdaj27SHy3kjNnr
A12vRdIw47EIvnUS3idvJ19f6EGWdyIG1ELeip4LHshxskmbSSqotn6IM4Etl+QJ
5Yxl7oGsRNSLliVL/SuVjpOVqMcEdng4StGFgATuR/fRCNHd/wKO/5/V6WatQtKZ
+5QGbnVpDYtgec2NWwhwRLQWKTbiYAZoYWxV/HZovNY7NiVA52YoP9xnL+4zWAWB
3aFHSf4Zwh3yhr3/+YWnfJrEYHBTdC1DnF6biOvcLMHIDLbNUcQC7ca5dvNfGIw/
NLCjqwi+ndpNhKzqdhGqxy8LZEd6p4CTvkpPsKVRYbdLvDfUpt2ATLLPrQqxXa2L
wDIT+Bo4y9EZ8ZnOZfIIaWg2eiNm94dtEtXhK93WAdhpO92gnSDLd83wdyJP95Sn
Ok6STQcPf+Ci7iPdeAatcUi7DmE7e5BNxyGm34JzZfwj9oqjqpJiQ7/S2rJMu+ep
7IaaKMkatwyv3m/wRd3kiQyKKS8fYxQg6+3Ix52rDJcbrZQA3f2pfBVqG1P8oco9
hyZ969PBGF58tfwtlVQCufyKGzYmBrUbPgl40QGd/+NQVo/2YKdNc5lfSmuLT0YR
NLdozVbsNEUzZJv/Qhohnias7JgK+YKnfgYW186AYPkraj2xVhbEOvBFnETXSYT3
CEV/N8LV+mrSLNpDolqP6knXApVvnVV6VZj64/yJnPYo669dEpxzSbQrFnSxG9D1
btfdlmW4sQednZRMPwvArIoHGZYRDxISE0f0djjSowgv6X9ZPY4MSLvNi6mDxsC9
M9Wxhz0rBPeqVI9UNuNgMffVbcMF4t3ikv83U3Qb6aushgQCiTvHIldMWfWUASdx
hVeob9qRQfKj3W+G8mKX/UkGMwxKgjLSdnXKQi8tCCDoMLtQUIhAPCCqECcIgPe7
1szyqgQP9YAp7nBrqowAwRzshvq9vUhILS+czHTvOlVFgsElpnFhxmHTmj8ZeQb4
w17+1dxLm3XU6iUVu/Aun/lziHkWc10P9xUcVNDdcQNvyIQKsFI1jcfcGZYwU7Ji
S/G5mR9BDr9DgtOfwoO/8nFx+n0qglPJBeps3BRAl0jsPQta2drMYAOW0sbtEcw8
Ioq+xqhWPLB9FCDnWbjvZ365mZp6iYToncrqyo24dfyAUtIuUPxfJA36jHqZ/MjJ
uODsxGiYz2NUD9kaKliYnl8DF7vkrlo5xMTl1FcWzRjLiW7iwbOtHK0nLIqL6Fga
W2mjIOUjddkPMMxtEttYHnoIEOr2KRzli9APtjqLGv623bUnJmkp5P2HDiPfj4JW
+u9G3rJRzuo1m+Dd6shiIhKADVgkp8Zy56LHk5DyxAqPD6oSHj3PFv0RdNrNQ8Nl
TnHwDFGKNypkQb7exv+H/CIuQl9f4T0B6wSst1SZWniCc+B9+VtksdhAwQfT9dXf
MtJoSh5Zrl2/sR/sNzqCcThEN1B/ZykJYtzcjwyY5aIWJb2/efxT8culKAjCtBgj
vRMUiXpgI8qFI4WS6hfVf3nYC60GZuxRIx9G2LJZdxezL6X7ydY74RdFyLC4o9B5
lzWFWWgLHwikIph7Xh5MEjGnym5mnJgCAqd85dv126rgzk3mULdtiHq+JvV33RFH
u0JSStaV9+DL9vbIAeaeJHitEXKNQ+cnIr7ixib1t+ttcA/lkHnWcjjIG3aHKYzP
9yIx1BZ9j35qTH6EJrXmwRBtbTB1KJMS21UOvQ07G4DCBOjDKDVppBTVlLVFBgKK
DkgRJqTm5/pfZipOq50BiIwtPaCiF0HlEhUHOvbTFlW7HkkK0HSADHE8XMQIVRno
iMynO86NzNmFhsfSq821fP088fIlaUGyAHoEZdMkhu/N6fCdhFoIexHZM2JUK+nC
trNholKv7Zm3D+4nkMtFy3grCdRQcIIcMuXyAP2NM/XYa0QWA8pBmbDGlecMrCM/
sZ8ZhD98/Msp/WIiZYSIGj4BuaeUthQBguXbmDC8HPl9qFtxTTrZv6jrK/3Sz8Es
aqtgp41AT8kOqdAVadk9OLA15JK7EelnG7qLDcFMxWUwhwUJuH7dtGawloBXPpXD
sRo/Ehn7UvxFzM4tmzvJwt4wFnK1rFKYw50NlMxZ9YjXG+wE1GHoolm+ee4DkAOP
idO040+Cy1RntZTsZUABCJkWxOsiHFgMweLyGfoJQmuex9TwSub0fbQminLYhSUF
qftKYpvFit4G84jq6a3fLWkx8vfY19hJa3GxmGnwdEmhb+4jQs3U1ew9WN+kGRf9
1TO7Nb3BnQEEJBvWXfPtGbfj2hZKZRzT1xANqZ9tuvOPqyh2iit5rYo32rh4wB97
DTCB9DlqUW7VinyJDvxiDBIoDsXF9RkABssLrI36zlxkqykCDoNvxJoE3JOHuWJr
1O+5Mky9oBdkQST907/Wax02BuFX5aoEApkCmZLz1oLmGApH0L2Y66kCXErZEliX
E7rcPXbjGv5qWQrTLsoq2/0ZTNNCj9EKkzGzFyBrLEzYVoJPJOqBI6m8ZTkGxysF
jfFf1HxVUCpC8YkmK0/9vyzrQ2odLMegqXxOMwLv/9Gd62MXtTA8FpEJpGO7F7AB
I9T3sGJpe6C/+ipNvJTHqlpQJHaKvWwk/0oY1TMSMYbN/afnsFtsRJSzjs2c8Uhs
eHd2yYiA0bPGtzA93wbglKSkgsu2d3G1CgTR18EtRhfK0VoWLTbQF+24vK+vUyBS
JbamSY9JpQS0dtfemQ7ernPctpDMqqUhBHA6u5LiRM7R5km1rQ+43zhmfIb5vdpH
Q7F06RKneWkmVXzL9L7MwwbSDiELKDAixqvIMmnw11cmgIqndwZZN45ETKuKlXro
wUh/TUzr/87iqCmzaGGIryrkIHxnVSyDRSB0w9Es9bv2NQ29tFuiEve1BPViLcPo
p7fCP1tvdvBmVzmWkAp54PS0iZmdH5ax5eqd4nGFpyuy0uI8N3cTnS0LTIZVq/XM
hNOEwM/95KbzpmV4zcJqqOVFrFuMJ5nKgVY0B2ykHgFAVgLsWtqQYMe534xqhccM
XjrP2LsDy4x/QK+ejRW3cTdWfYNzmsZ24IaVPpHsLgDg1cx3ocvJBDy0PYdhJrkr
XhikOVspmWxH5l9gHQ35oL6nK0fvTzEl3CRLM/JDI/bK0URv0aQjZvNa6VWsy44y
D4X2yQPXx0Vyw+Mkh4ytrNaVePIepqPHO9DgssLHNLmL0u/744S3PkNFgfREXuAo
EpDlW4M65PRzIBeFcqeWLKnkya7xhdW/QdNg2f8UZPFsy8g8Oe8lv89ceDo6NyNU
3Wxilv2FosXjnYYk77fRbJXdtGoateE5O+YIibqD7WuB50Eky0IpC/noCy4D3CQb
oFOoMBZc54TZS2fUXbUeqggXgauZW0ZFk/5pUr4Gc0yE2ecxTVud/acFYloCbVGa
YAs1/HsW0zxHBaDJb/8H8Pia3S6HpkXu2mM55CHnwBzBuFh3+D9RALaSt/nFmW4A
oWzT+2w2fkALcyAxcNjkFZCCT+9zvKTtmfEzrtKINnCYuszwq3WdFOvuFJrgLL8y
V6Wn5KvOjWZpe0eQKS4AnMSgH+GhgdDLrCV+1K1nKyzc5BJQIU3Nx6P1xTMHZT9S
7UUGQP0mLn3Q6A9zuJsL/mxjTxFyrkgzjPeE+zZpUQCvBOzlrAOzPETKlhVKZ/6C
EDZdgn93iny6EjbdDA7ykWw5bhgsALJWQk3CLqRh6fYOKbCGeVWFskWa3Tzysu1K
q8QDihf8asDf13XoVpV6NwszY/exYbGaLmPE/qJmCtJaCf7lf4y0NBJYhfqADv32
KwZmBSCWK84CDTUQ72J5R4JWnjkk7nItcY43wY7AovsNRRi0IkCRJg/3AQi5kZ4i
KAPWRNlAD4EEix7eoPNHWIp62EevB0GmzZGRnw2z4UVYdrH5eLnxDmfE1nsEv0wh
X5b7N+Da9iq4ThBaUWb4arEVEsjvDaHdDalp+xpV/hhIkMFgO/U4Xzrn1vy6mLH/
GrvphVTzgM1dw05mpaWxTimlvkxJH9aY3N4dtAcPjBQk+v9bjvPa8kIB3j+dP/vS
fhXMsNa94rCKI22qrtJMwGRp5LVi7RkLlld1/4IQSs2JhcEGl4rrh4057Q27uxii
YRZYzIoXfEqpxiKSoDZQ7w1OSS3Wu3vWeWhxWivw7S3SszGwZFpNLHKVbvCz1nER
E0uVy8q8EXqNWyhSPd/+dCgw+mZkPXjLudZUjL2zg7HcMaEgXxeZhSgCQv/xd9/c
vHYKtRfpov//UmXms/22IPYbd+eui6Tq/o+nDzBQSsRCwCyifNgnheDL165UQRat
j79sDfkEp4ot6pF/bOKWG77cqy5Ac9PV18wO416HpeK5wbKMMjwEBnudUqA1YEde
4lxzL36VTXnYOZA4pd6gcPI5P//Yt+PK5xKdbAaqtvxxFTjKGvlvQCamCQtUmGvJ
EuIYorOfhVKcsVFUMJS7qNq9X3Z+4kPSp/9BbYX9d1aLrQ4oQtkA/iYAC34AYDZL
5jl+bEYHr0dC8qphLYT6x+P4uuQVqcFuiGk51LBJOL/KPBGCXBGSmcHSdooEMTyY
RZBCLgAYgMwDyjnHgrzN1Kpcnw6zW1oltBRIIYC3cYvXVlZpvGXza0yXffV6jX3h
EUqXoH2b3x1aIVFFNdijojMSbaE3P1n+1LwtyHfj739pgu+jogTXn0AZg3rQicto
pUKiULYeTKMeKHPoToDaCHYXWFz5zsnzG5pvCy5fNQdxDmTSmlG+nXj/4jHj9Q8o
rRNQej2VajARyEiC/dkkiNvOPtcn7p6kQ8bR9kprW4lmcK3UvJElzo+0/Um3h6kX
NVDepO1rINyLodlLQ/de7yvMSee8686OmllQiFrahFfx3+IeR8DdIJF8+UUFqB0R
rbHSTNx19n7hkxS7QkLkIENI8Ee/NC/pfONbSfZRsyBPSp0XDUesoVfiYnbkxIYA
oGv+43QsWQHvGI5zKn21+9sAAvxcCEQwRXMOOXcSEykuxNBc/38u8gKg6J2S0r7W
OPoQii435x6S1vF7ClHqwkjL+xjJPIe0YFpRPfRONTZMgM1z++BMCkBauCPePJa1
NdNPZubrPLcCA/L8KGirKSuURxsYXQyckZZHEdqT4odgoapVgCnDxBE33PssNpjQ
vB6nH7riHjQ9EbaZ1i8lCT77VSd2TjEgvWh2wYWhXFbTrfrz/PI2QP0y8DkzSrKz
XY30OMvnTE6nqdXeWkRVQVtqokci3Dnk2B2MxkQ7t579JuZIU1vnszOpR/Kc9jf7
YjEFdbt6Uh7cKskyOaA7yGbNAyOO+UnZgo86bv6odK+hJLZEcNj6n9xUh3ZBCmZ0
nCfoQLMUnaDBRjnzt/flcqJ57EKXJmeoWuFJtjgCn3QnSNR7oF/D9vQGtSEsT8IG
iiFA3ACHt3NgmvDbofGDmIOf3kQUIUh3MtTIZCNI67PRNE/d/PQaaG/gxGELFE9d
yUFmdAnpdU5dQXwvc37WAHDrJWrnfYmiVOGA20QvPi0t7vZyOECYkf/swJhRwD3c
mETx3uNn+BkEIyeSecy62JEEDRIMpY3xP3utqqyrevVDjpjzBwSE0Xv41NwOxJR1
LVeJMiYl424ZFZvWhovw/ZtzYVFJS+sFxz4HPe3FsmyTzytt+MEYfOrMpY0j+gHo
VGEmLl4/cAP0IGjMsdmVUodQLpm1SOjp/iFbwrei97yUcYx7cXD7mTbPc81Q9hJX
w1D8kDpW80Axe03t6SP+wFnGw0yBeKFVxb05KfiNcSd1GaaN9JyLnhG5j7Z7CGah
avo2gHpywz0q+Fwdv/bXExu4MKlEKOZFdXL+pqjjf36KL0l3/2LhLClMC4KLpgOi
JE3NbMeFrt1IdQXFBqJD4PEuZMyM9Xl2AQIy38fYKO/CGPswpZhmNXrW0nKOvuAW
QV6SUNg69vccycbepwMS6y5ecalwotWFtoKyRGVjww7xwEQDyuMR+WuTgx9LmHA6
94qIh+P50nRjK0JqbWr9nn9h9CRmNCRm/njj8KfRgntGk1KYVVJvE8HwTtGGd4yv
8YR3f1fesdq6xmpO/y2ePw+jiJf0XNIZ+q4fRsghrY6pYbMyvGI4tYGzr+4xJdor
wevIhbn+3LTbO9ap9KPSWgYCYOYQ+rk7loRB7TB8ms2MwtMGdHiFg6Ihr8JuyNbd
QtiBb8CJiaPK9LFDg4mlnIrZsvidJoz+Iy7nQSS7RNQoVaR3H5h4v+awwV1anWRD
LNgSlai/oxw8KTNthduPP/31rmUtOKr87mQoRgU8piWTIjzSq8Ah+xkmNSZovmMX
IPpDB0fNJ8w9C9S5jwBdujI6peDG+fDQA0mG+UdqO41au1HpNDqJrgUSrqp5sKEe
bJ7Bar94b2E0vWj3fKBJLCmjuxGJeLX68PU36+ipKNDCWOaYFmR3Ay0bfRiosmX4
XB0pgg+W2I5d2UyBpgyYOLqCXOYPuDoXwO6Uy8Ia9Ckfrma76ZLY6gRhxl8xTsY5
V0ZqWsHsDMuIm2Qp7Hkqo9eS1RuOtD/Fy4RCvZ59ZTnEwQVIgRaWUWebJo+Xmx/d
zNmm0biDfAR+sozreT3Sj7ih1DTYoliN4WoPblSIl+0oIwootwuekRV2C27BAyfx
TcnQT/2Y2omD3RAPXwqBAq3vq6M0ATgcdgqk1S2+74HlG024+iM+L87YUAKfS/QN
h+WN9beOgMd9yyy/cryAhUBvSHlLMhs+ht+RC4A4MY7HSAwQO/FHeAy5/Up/yD9t
DT7XFxsC1uV/Fy908WF7S3+aCzMSn9zdiIvvlISKSlNQsQzynvh9lhoNirR34Yg6
OAHgcVe+zNHuRA4x9b+rvbNlw4izeCaTq0GDTmzEQSJcaT/1/DI6HEscJocxL+AA
IJ+4TZheEwaqePpDOPhn5V54jYsSj9nbkWjCTNQaf4R8v8DRzNoJp7A+0wZi8zU0
ilIKI8JYZm0yAsi06Cs2mHsmssl82YL5J+3FzG8/VHBi+iiXPm3emZwGY2QyEruK
eIQL61wXq4KTOmTJ3kjIVVvTgpgVU0HXZkL7Sm0kNWj+RNeARuaoXxFLWl8F7udN
hplHVM1FfnwcZ+lM8jg6uFYdRpYrCFCuByGomLs2ha6iXkik51PG6OI1kydGw0+b
SpPL3qUZGOdnnBRyGe00lASCuZfoFOcZsO/yB9HSRag5h3QsT8VDk3B5Bl5rFTL9
ZLkmklyysnS7kpBiPWZwjrLcXEh3vuOL2/tHjxjWgHypimsrmOyaqwjWJJv+5gfI
CE13m0dK8yMcsBOa7Xu/nB5dHSnbaiJM6hwOgzOqunTE/fR6I2mANqxNO9Fwb+/R
klxNerfopj/n9/qH2FxJhmTaYdBRgxwazT3/baAMNV6XDblLgWPttYdMqeJUrYnJ
jDRGZhLBK9+L5QmKyoaAGZInnPXuAaTx6I+pWj4vTNWcCR319P5L/oEBKKIUtwlO
XBP8YGiQaDLZYVJj8AOq9PPunVGkYjZCuWbzbAWGE36azKtvK4NWWpzJtUKYG0Ov
bJm8L55nfoiKfGAiLq975Bfavi+BE0Gp1DKSlxOFIT2pgKbhanh5g76fBJZa7fev
LRLzTcEVZ1kgA5JYZiO5slWG8XI3SqiIrC7eFB2cBW1q25IachroUt/j2SOoVrcD
DKOe1NS9b3Ahp1Y662i01AbOeyA0PimS6t/zwdprSNQANBMjzeW561+vkXvpFRg0
B9GarCI8Sl1I+RqxiaJTBfLsdGQqiRf+hzEo1+li9NHY1rGeW/R2Ys0cyd7K8rCW
wOoch/R4lHPQZ030U7IkX+n2XCCRQZFk/aSaQhfjmipqckjljU+hBi+h9TTvZJ2E
SPS0sFvw7P4aZcodArICLgV/CiDTClFc9tGsOnBMl77qrBMTC1IZjGDUQsVCp6H+
6rX8LUtP3c9eKcpmDRrLLSUTZfDjuc0Y6JoOqQXIQoIdJCoRbBKNJugzizQw/r78
Wq+UmTbw4tpKNpa+y34K2NIMbHy/AaxTrl4W4xR1e3+3NU2rp3kOR/QR3yo5FRl1
56RAk/ZDFjcjS8HVRe6RXm70/8sNCQGTnk5HZUuIylOh9qHbGLt6bgKz+cT2sQHm
AGl814haOc8JuN6mANTDpKZIjNUwn/X6ywpDD/NGBwvP5IK5mtRmL+5S2ADtxhwT
LPaO/b4OK0BRzGDM0x1EdoIXitGKlXwS0aUyyERDFoXzRlcFdg0+pfmh/m+Gvzu8
RIQpmMsA+AWAnPxUrJAFh+fskP3B/H7sBSgp4+kKqXn17GQawQsJJVWbS6rC7TVP
d2huiK4v5Jvzm5QUYzTKx2LIdPd1D+8Jk/60xKq207hIUQU11TNAH4IRMWHZHphx
5vPflmD8m45JjG+vGv8o1krQ+uM5kpOVj2A8rPuCqPX4BZg1W4dntJTl6M0R5W2p
b0aglko8fO8erSJCuWJrsTxDIlaSnCQof7CRetL24aW2GUC5rvl1awaX7T76WXsa
jV4IR7Lskxm5VQOdgeXupC14ISxgoqcc6PPEtnXqDUmw4LbZcauNMhOnqMZbJPO4
iqMHrs3LwTn9bAEORpFvrt2SpXpxC8CPU7ZDr6m6b7kNLDP14OWd1irTa09cksOg
kzed5EdNDEC59+AGqms0+ToeanW9W/p13ol6u6D5N8Vroip4VaMcKTJGckgmQcYD
JgzQgI6J56d9b70eKVDNH77vRbY6fiSpaGxRtK1U6hvSHroaM9o9s3vkWqc51NLH
3Opnip/ua7u/wiqH929NRrOBTlu41uo/ugFZXQY4mTolPNFB3XmA2VrvfnDGPPxQ
7jnEAKkJAGWJeqvdUwXnDRLJUlmf/X+VwJaRaqzZBnt912A5Qtg73PVwspwOnW8z
88YUxz4DIzeo8ymJAZ5D7vqTRVpqqnF3bCWN5oxLGv2ZqmHDU0GQnDKGCt8MSyYN
nsrBoEuCDTljlIEn1hi9hdzBTMGdjp5hD3rPGmpcgW4lXxBW7YgnHKPFX/JUmBjs
BfnuwENvzNgjAEEQcPtL8nuTmO5x3VmlxwmXGL51RcPaF5NQelIRKMlroksMcnXG
YOvgFUINNr7hbMEMfz0Avdr8TwVosIZOF0fyiJYvqNJcSO+OHs7B+sTDPLxfjkfG
4xhM+AwYBdZlaxllcjdrgTKTKTf8sgyN0FOlVizqf93LcreovqINFZebNt6rj+Qz
5ArPbHLKd8w48AMrxJ5cRQP9rsA/oQ04A/lFGOeiP3BaPOkw+ZMisRFHGFJ97FRu
0oM9FvWBlaUF+iMPsdSphEuOjxFeoljxF33enYk7JhRkD6a7kZ4IMEaBTQb5wgxD
H1GewwJ75Z0zNy0PoRQoptb8UFjCDDr46f15zSRlXb4LG+RHnRuhjWGKUlLHx7Lv
yCVuWODxdTbYRk+/HKweW1z4YjwDp0QqQPrjLyVXYhZXp7YFRfWPAvXvMw8YjX6o
crYF18YLtUMeAEtGgHxqmNGGlMflefXndkB+lkUsHVmqBvzdLgAY/9GrrfqgZUI8
pvYY5M3UIl0liOC7SHlz/KKcX4iqhspKimNtgAzM+6SR7RYTTtId4AK9h5CAJZ+B
mJtyp/B/2W+hU0VxmhlAYJZ+edRPPA3Znnq8RbI7Pz87yOLkzP1gdBrpp/FPZc4P
fFRRmWaIZvNSHjlXcDEL0Kwh+voNtewfK3n3Ov5Eq3/eCN6aQo5TI9jiqjLLxtNq
J/3INKE+NNetjuQ91pv1gBQrouJDuqJt7srJwXCO4l7DP6m82zBYJeWK2FCM1eNR
1WqiLSPETSkVKG/cxSisV1aOjMocqO9JHGQRlldBWM01iDFUimDI4voURZPHVsMH
2QgUSCdL4S3+EdpGQLzMutc8yfkx43geGhm99aqS7Lg5C9y4Bitnpow4XqWG5dFG
zg6y6+UuX35/K/tu3nsVf+u1qdGxnRhuV8/hJHxdFKS52OFvmO1tr3gfNQQl1Spr
5LcT9b2Q03IPxUr2bxdg/znjBKs/KYQK8I2Y93k89rdwU3shlN8tx5nmWV00GYHt
hSkVT5NXjUbaLC3AixV6hk0r/AFibGIAE3HPpJiImcs8eirBO4fXUZidgNctd1lO
ZLq6Yo6pKd6qU08Zx/37R8XOCOUWvTQhcS0VFV1gqYB4Oh0roY2V+0knf1Ozq+Uv
VF6tWgV8LJl75d7IiAZCTrWyOd8FQPwreoDgWCt5DNJ4GmCwSLJJk0RJnTQV3h9h
xQZFql2ERDOub4anbklVnZ6t0Gag4FintiOfsVr4ool8nQv7i5BVcrTruaK04wKr
FFHD4MINVBk3/a0y8lwSHCgcbXnTfhD9Mo29wCQBaLl7UuEwC0i6zvcpO+GCotfq
WVxz3V2MSvaHgL9vbFhMvMB587VE9dF/GtKDxmfv6P+xnsLxl1x55QPdhjd5z0o5
RUNOXTU3OSyeRy1i4SURnBf7VHwE+X+S9mHZAYdlTQnYbDtuulH/1fI/iqzbaw2J
cOvwOPtrp+GmmusU2cPSme6pen1P3gK1wI9LKIeRcJfQ7nnkWjm3CFL6Q4IBpmf2
llcR2OT3z+AWy9bhJPoFV+x0dh1pqrXCUw8NHfRO8X7KT4RTXpbczSIGXDB2z2Zh
G93eLcqMchp5w2gcf48codrWh9uNot6s9gAGNf9ajudjwh2DXwmEC+snvsqEWpSa
dBAStDD3DdMScW94FlMaFu9L5bhZ6AWV55uVWf9KKYMkjkTacNOftrsEX0GicI2a
ZbIUTGng/CFynGYiW+R0PSwkzjOOHhBZNTy0203avBDf6XSTdsgn11fPDKWPyefa
bkyO31QI9wOgKuUzPAIHuNtGHqMCItys6bnDqIXJDSWaKowxSRWnhB+brfykv5Yv
zsq53wmVbi1jz01KwOYpqhUOAcqwn7MB2ofycJMPSWiKyo2tpgETIOgs4RzwlMHm
y12dN+opU0elT4VJiUutcRh6YmGExpe10uS19O+0IBf6QOK3iwOZexetqjIFQMrX
IQOM8P6H6SsJ4JdYJuPHaZjfpb6qfHUHFLchgpQVD1uREwLcRAiY2LkN4QXCD8te
CteEEPoKYK8WlPelUKOWGcWLkHBexEvfnHzIU/UVjcg8ndS9+wqOUNoy/rt3BS/n
W6sMOlI03JqAt58kLi9gwZtpNCoP164nl8yY2kVvTGIurgzVleoE4ijK9Er9BR6d
gxHp6m8DfEtJsab0760F8E4HmcrMAioHPioM2Qw3tcmpyxqu4tX57JO3w+lfg63S
L4jCSOtqDyhfZJRsH07iFM+OC7QWxeQs3IQwtTCHMmMTqg/FGQ/etO3oXpXtETEK
iaBlqS9S95pdOp9RHSeAqkwPlvDlRmNL0uNW317rjZBjH9/2Kmjt0wopnPf+Pyjl
4KCCo6C3y/x3zWzloHkcVVqkPmZno3Txz8HUMY/gPUFLQ4hF5iURjebuS6GVu1Wi
4E/K+v6lqeS9rAMeBX14hfMEp4M8ml+76wE9o03zj2Mv6f429T4kcfAxusp7HJTo
AmjgMnSKgGFJ23JluWf8pEVfMIOPw+mHYXxf7mUhYmqiMxzDaDJ+buZgm8+SxgmY
uF9DdMjQLmKoRkC+NvKSk8WYIidNtWifFQjKrb9/bGQorB4HKdEtktUcKrBF5Bst
yfKjb2S+7Iw1bPPD9OK7hDC/Jn4rglD9oPKaD+pc9Af9i+RGlH/cKisOy9zWN3AM
KIrnMcUAE96+u9vc6F3aWFkRedyajuB3x3kF6rCAAfkN79OsX0g/6H57agiSeQJh
4sKYmo7gvM635pv1sN01CpfqKUXX7WYbMFsElUx7M9MSy+a0q2YvYRxn3zKBiQqB
+Jm03Ng4sC1QPSbIgS8uTHCo+TgK69fQlWMU1fMFviv+2xZDOVF7iBfkswf1XPlA
w76CjjtFtjUmFr7DUatnPN0SN+j9vk0Jr3rmJ7u1eE3TVRpJ2PpFMUctEFHSzLdA
K7y84sg8w/HNVa76PNCfBxZW6shUrkNKxiCo3pAMCCF46gItjm5NCet6YUzYpuNN
Ae5gD+qCu+yhPUYpgUJ+xXiYcLtgcd01AclfpviG/BYfMP6JQvghkmQB6EONm9YJ
icn9KCABVSasKiFkq/X73lIevN4G/TKZ7P/Zjrf6a9caaKSclfCJFI02AEYwum+3
cmTpbun/mYhHi4iipQEqplWjzke2wVRZ8EeKQtZHk4BYlBEpMK+SGQidpXJdDXse
4w3ONK7DReSiesPtrp4A8wbhhohIHE8+5DO3NQhClGnQLtkvKYgDWENnIUsH8bBU
UGb9WdbeuyUZz4YFXIUc5sP+raFYl9jV8OqTWWjZzDiDC+edebir0zVG3laeFWhf
sk4fMhmGWyOim2PkEm3Fy5QMXKrxiHZJPyRYKlcv72aNwgZ/MIc0ITYV6risnfHe
3FblLQo0JGF7aWiDWQFX04VmzJtmPOO4CAsdGJdqOrj/P4EahH6b3Gg2YGyHDVCO
tMkQVh4OxLzmWg3rscAylIkR2n5N8qVzJSwtFqvR8uKNhaQ9cGBvDzLWL/NUMl3V
2b2MYRqfua9HvqD2MbdkPaD7P7lcUaG0iEhd0sp5/eVY5GX81NPmD5wE81R1NQwo
R+xe+SqAI5kNf6Fupe3dj81IvzY3SJ36YKshQpW7JG1PvXAJRIoQwW7GZQHdq+Lb
ONfs6khjUqZxegwiL4rwOICLDPI40Ub88uupJSQMNFy/4+GUWutu1VeU2QYX+8vd
2XDuOrEeyC9xD/a1ME0+Mgqiu4gvZ1KQvUxB2B+ISGxoNcT/HlFeYN7xs+60wmQB
fttR4OQOB8c94IAnXBS4R71G2ULN+bFrK/E6gN1YRYSUxhgieGk9ReJvvYhDtdpH
5I1JvBBYMoPzbLHtL/jEBgpBJVfZK0beSTPye9HAgbxhLI+jBGsP++L2czYDcYBp
mCJpU4RTkaieqVpJTfr5EjYBZgkyLYxaHRT93/m2mGUvZtZ7f7/kEM4qtymCDGo4
OBxG19RI2OA9i2bqoPeYctySGSsCGPOzzM7GjQzSkw4n4TR4akC37KAkF7YLnOdp
3pArUv8ZtYIQtUeZunrWjRSKFhdNN3uWtcq25GDGZFu2dEeaYRtoKsUj9OJD7ZI+
zLtusyHB5+BO+maN4BuHk1LMlKGuLkMwKCfo3Hw5a1Y=
`protect END_PROTECTED
