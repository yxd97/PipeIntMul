`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/3jH4zs3KcXEFY7shG4hapvaeMnNcY3rfjRRtdzke3VAXMvnVkBHSMYcn1w0cQaL
3VHr5cXJMz+gdAup6Q+FtT5Q137Dml4OHopNfbZV/VHfKX1sPXNN3G6H2WfD6DUd
1w5e3Qa8i7qRiU6FWdSIkYN8qdS5vymsLSCmlEhAgqyq3Cx7x6BNTz/q3lgn3sFI
cnvATplIhPzhqyhPdvpotK66vOSbmQgHJe7AjxTOKIxC2O7qc4vEGwinHIHRctM+
QJ1bTplG07Jb9K+jJwHaxvKQKMqmN82Dfwb0v+R/Dqkmus7THpis0c7F7eUb79c4
Yq7nxS8ML3YeqHJKVTccvawZpuh1wCijtV2vlUYTI0DXmYWmJMbNAUc1JAlTtT2+
+JSHWmaH1axwBOoq8zoCHGLTnS6n15yVgnWXNWMVHwOydS6oa0gOuTv24krZgFCb
/cZz6MtR6Jm6AvCzWWBDl83iUNav6g06NQi23GTQi7+M99EYuhYIY1zh57ZZAU1s
+FxBc2LqEdZ9vvYs/5QPplqtcAP4anJpLGlRuFmg0pR2nipQj7Db5sD+hquIMBg8
C5+Y7rPCXXd+rIVHRFDhbwrIHMMYaRXicQ99pWNCVp8CTMjHCvABldAebOJQndSu
Q4DzcsWla18bYoQMEEG12P1/CJTbLPTu6hvMge1lHSG6lBPaSLrv89S4fyz/kRb7
6Lluezmlfha1QbKhVTpRsZlc001JHEgeczs8xvT9azSULr0GxM+pQam7zNJdZ8FE
GxbLf4iTsiPQ4WT2MIzjjhMFhh7t18B7XxFzR+voFetx0muxxtOLSXaqXWe5/97J
VSS1Ux0H9WfihDNPuB9wosABl+yHKeEpVjAO0HD2Ku9I2rI42lqn354C/LYBq9Cc
/Nb4j5uqWl/sW86pQE5F2w==
`protect END_PROTECTED
