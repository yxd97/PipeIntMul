`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LY3NFA1uub4sRXl0nPoHphippXEZjXgU+rY8hzRllIoad0jmWNBCmUMhxgh1bqdi
ui67wvRPN+vXr0cjTV6wW8qrskHM3ig0nf7B6tK+Jv4zGxfeR3vZEPUZTLrNkzOf
mF6q/S30fz5zcEebYNYa4Nf5Mdr0/QOqa4g5KDyU1t5O6zA9gzdq8PdvSulErV5g
usanBq63Hh+3ds1cM+ldfYDcVVO9KvJsZGRQV6OIyiKvHpJUqXz5HaunThJChrcr
QTgtf/hJLLtiIwdo0vUllsv7HlnUCSXZvY5BSq0Jj7KfMCOPWcM+0deKq/xWdrmj
QHIbj4nKEhafrndOciP4XHuU53S92xsfOLTTh7pKflqUz2GWuus6/O8sXQXACinQ
zYJ5L2ezR/03bXqqqimJxdWHGKgIeRGUMuPhB/8xtDsWvVTrtnie1AOQvyixS1+d
Vzk3X30u3U8QNWg+1CoGdgCg5BX0JQK3nPuKnNvomYUiTMgXd7gNKVQ7KdWDiamE
Ddr7Lczsi377a3O+dS3bXvViHI7KI/R43b9zEVmOVA7p0ysnnm2//f7ebW6QUTUE
PTHeW4uefpf/ZLorlv0n+jtsiHmS4K8m4eGY4aJb5JB5aCDjJkK73DRiJspY9iar
dGTCcmjU0onuBiRhQoD+3DbC3Q2RKZzqpb/VEqWEKd9o1O9IvykyItQ+Xx+uU42g
dobboHf4nJ5N0h85fHjcCi+D6+n5pMcfq8Eof3O2DrzSqOlpuCGRe2ddjbGSQUl4
ekSXLeSq8LVxjSKe8U9uZphMSi5fNY9goXyjcLW7M+mdhpIsyCAC+EGeezcelHrA
BBpMewJfqHzPlysvf3Fyn7XMBmjyL+7sbWU8NIesP5kZrtWKAB0hnvjfs46yLvie
KZnCbsKveYP7F1ga4NNztZ45nUJEnX7pG40M4czGTxz19flReQ9tUy5cxB9UYx+3
kiSTotC9RnXcQSREp1qFdEMwTZPcn4PADYz87vzHO9L04WfyPBRIkRxUbQ5qPx5Y
l3rT1VuRaPmsOHHzZJgfgmneB3QqokJ3SXYNqk1VqN5aDzP2uqqZ1fNrA7Ro7o+7
SOx9ufcGC/nK0y8Tzf+0zClqDnVnd0FJTrS3027ixn1MOZeEStpLMXBxmhFZY5hd
G9RJZn/xiN4QuKOXXblngdRAixlzbqi4+Waea9jsD6Q0hcSc4HnruLylN4lFfQ5B
baWpaNhmjH3/fMOIFOEZq5CPUCv3dN2zlk/d4f/snFeCENrHdMwIk37IqwgDtVe+
mpYWec7djrOlYP8Ev2nNuWgyCcDCohB45QPEPz+WbFFjIH8Po5+0kPb7OadywM78
KDpPic2QsxA/E0k8YsB+gpXn3jPe8IZMkDrBGJW5koH0Y9+XKaGodXOMQNQhyInj
zKCgo7BbEI/veGX8Vwo7gj/aUSCtNAljPSW7VR/5MThEkGxgY8IAgyPotK1imXOQ
iNM4McYsIq37f5L5FtyM7vz47D5GuCkl4X6kIUYkiQ76B9t1+OFppcwIOvFSZYdz
o4Z57pJfpmRdbwio99Et1fzBSSWbcCESlz3JAl7nLpJV9QNAcWBtJsW254D0rg9g
zf9p5+1wpf6snKm2d3m+W1UlnNHdDWCiFUoSCLaAqjb9xoUGcFkQcB3TRARVcEul
tiTsZN15ptaJVd5TY7w2nfHYBtHI/jGk3QvX9IJVmhMHuvrORMXKP/1ZDQL5DpKV
2YM5B4mYD4KfQ9GWOfuoKMyIKt80/FxW/bn8l0P5gGAF78YYruObst+S71IOONc0
bhOMmz0Cfb0S75Z4kM/R4vEBiz398dzxf0kPN4ITVovEO/6EjjQBiQRfKH5dtTNO
+tydz/SAjYdWXTC8G/jdEhqSvi9JZiymObJSo2LQ02JYso1UJs3KvgWqK6aDnfeI
LAQbTW8K4Fdl8kTDnCG+Qq+PvCK0A8HCyTH9Avvo9RAYbiBu+QA43tLNlCjHHaNC
E8XvobZydehr2KuPxjyBxVeIj/qUaYAQHt2NHrkARkHUq3A6ePzTuzVQELJhLQm/
FVGvJ++7hZf1Dj+dIn9AI/mVI3SIdcrGt2pXBx8CCGKITcxG9oh7QCQwn+G8f5xq
M5EqTRf2fNXqmN9U1oXvwBLySUzzzkqS4A8mi8CxbVXh6kFbdB9Q4yVSpjC+C8+M
3eewFg2zWQx7kKZSq/aEg9URi7bLJkxgkafEeDASNvk=
`protect END_PROTECTED
