`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/Lnw9DbCpMZmwaWtn6G9XnYpxit0kBPLc/FgPpH+HgCs6SHeR8dWX+ZvWakJW4P
UXOj1WtfnJ7CU7gsvyqUTzYt1ghx1SQgdx1rOs+q0iyHpfD2TICCvSoHANC2ABtw
X7a9mVIY/PIDXByXwxxStibs5ND8K4g5yfV4wAKNB9AmvZIjS2VOS2Ol/NLFKYJa
ySq1jUrmUlPKA/5xjGCFqcnmW5loGFA82PqVcKzou4qutYOsF7sVsNqpPfA8JIj0
WWxaVeUVmYoatOI8bQ4GXJkK99Zj4tLCbZI/+MFwaO0aOQUAau3epiHPjkZfUnAY
nHriq56wi52eKty+1ER03ZyBheKHpd2URDNyd99LiqeWLDjNgIGocgPVYNRfE9Ke
iu1CJj23Am88nl7quN1nSA2T7UiY7EVT4qRKU+skhGiTChFVpMzi3YKoqL8FXDnO
4HUDFDXZLZE4R5YV97xhf9lGwHPq2cxg8KSHB/U6vr/i850cHAety5to79ADXujo
zRetv3SuZakhpBv7vb9A5YN8GylT24y+Xs+hWslduV+Aleh0sa74tOcJtLlpXUfL
D/x8Q2mPUFjWqAM9hyspGICbQSyug3XUzm+CTV6vuoB6yuurwUL14gZ05JXKA7Z3
daMNDagdRS9Fm+Ka6uBYDBVOWj8Nciis4EpyaapFQEcncbhTbaarIc+sY3ytRFeU
6+38m17Y4/6EOe+9uolNH1O3miIJNnsCu/+Q5psuVHkzRbXOT7yfcQPRYhlC+n7r
v5KnKRLv90+PN5+xgV8ZYj8rMPJmdeeVqJh6wTAuNog5hSumFa+QlR8kilX3RCoz
+M/17Us8XstdXAuykYB0uw==
`protect END_PROTECTED
