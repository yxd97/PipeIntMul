`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5wIXNYE9YgkS0k0wwUjjW7wBq4fr8PFwUEjXXskOI0okxLMGilHmfC7c4pyih1AU
OlTvTijUcIqenlNJTT5yOXDcQTVWPn/W10OB5rFcAA8heq6daR1cqCtXmWYlKnb1
26aUZt7MNbVPuWl6IUbtWsyPxbEvlJxKvBD+9TlezomhtUyV8lMOQVhiPzVP22m1
KaXVzncva42GoyoN7h7r0g8a8XLUBw2b+6Tp371QsVeNe/xXO1ucmlxxhmLGrcVf
vzJKc6pgQTI+6guKcp5MaylYLVJUo+qmWsl3bTVKYd289VRvdgVOROVTxWj0z1kx
lAQr70EWllIHmH8P0ncj6A==
`protect END_PROTECTED
