`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7b7IgQDoD39DqPo6jHN4JSQjdLL+wOIbsHdwnvWof/ee2QfcZgTj8ApJJIfdZ9o
XRTOsIOHlE4gWxHZT4u10pTnTZ6NJWmTsZCNZdDzn6xBhh8bPPdIScTjK0+BqiKF
+AvjlEpRjQwKfwuG7Qn8YP5MOAaWyPXcrbDfaG5S784gL74AHZpAG0noKproBm6v
NLY/0OsIjLXIqr49+nL1ZOXpEl7fx3Lh8gnGjeaHZgci/l9ibbZU9gCaVYNc++/d
KrmIcNhTC91hGjtDq+2bmnw1lcxBrvUJHLfQ7Sy1P8FPRqbq5axECYvsYbiPr6QF
E4wcTaU7vOkcVuwlnLf5eOIODhuCR6vz/e4KOabPDK7P3k4DhzWvCVknDCgtE/gp
7LS1T83IbbQ3eimK6xfbXSRDEnUzNoYQ+yJ8uKhs8sp9B7X9Wdry398FSAY5r46P
eQFKdIkBB4FJtwBgysq0RmpWyOYk4O5GOPNEntHZDt0YhmtMJ9KeCW0604O0Yxdr
`protect END_PROTECTED
