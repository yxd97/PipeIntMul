`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bulw/P9oeJvLsRGBQ+GK6z1+3TTRDeuMCe03wOITL4z7HnCN/Tg2mI4RSgMAAB8K
bGI2OJUxLG8xivLiPG0hJD+Gkgc7DNmYF7K+zaAdBMm8np335hfR/lSBN8rs+Fu5
LOyYlQim7R9phC0Uv8ONIDj16U3vQ0y+bYUjdQYqCJiGzhpbdOvHGGdxDmizFo2P
XSAev+aQpSxfGj54vJgVu3C2Js8fffWywpTeABGZxzMiO7+SYTUnsVNiluTJoxae
Fpeyfk+Vj7FE5EhPvJXY+xolYv28GioC6NhagynOcZrayfkrgJfMlvPoZVBW5TpA
cpcjltZLH0iud6Dx80DdrYwmOJXaAntqgzCEn8Dd8TZV1xepa/ASG5qktumR2uvo
4fOHcFDbfggr+2E5clusmbtgdKdXac1qqOHW42ESpiQuIr/Nw+GuWoL/ON13G+Ea
dy26cHRcID4tKMWnxyT76x3WHPEwqXKEOgWPRtWDuYRUtVzQEWt1tQZVHny+P/K0
OtNSdnDh+x1KFhEXV7WTe+ttzGbvnZvzzJR0I2uYE5SVq6mjK6Q7OtTvWLx/lDrc
C4PWzHwrTl16ezdCt8G6rH1p3EMvLiXvJcWefyDOhXZikdN+uh6WROZ6raLXuuoj
dXoMb9KvBpiuk3hzNDgy4o3BGVGfyKCf7ml1FAeHdyU=
`protect END_PROTECTED
