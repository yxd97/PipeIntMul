`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+JEHZnzRl1Jfx8e0dlXRACAGsGggPLrGQd8B5+NXux/aTAzTpF6FQqyWvZDlhw6
/T32yrH9fRI8O3gL9HK5wnjXaLBVPRi7RXGsIGCez54Ula3V4yVoN+EQBpFC41l/
xklB+J5g+mxioor5hChX1njPKBx6eDwzXJMQxnGGuQzGY67kPI+mLiBpqZMnq++4
QbhKHYha5AD1DHhJUI3KzYUAyXKdei+TvevSqYbyw0lev4lVOTEZMyyozzikIYCO
GIOl20QfPgCf5s+l8JSmob1UDUSHoc1kRwG2q3aU3sPe6fsVERBHKF+5moXmww9a
IV3Yy11Ktyg086W0wi3ZYNLzb+rl00u0eceqa8l1OtQSD6sSq88IFgFhGcDwsWYe
r/AkGjxntwtOy7hrcZbpnelhcs7rB9TaUaiILbdCkIRsuWzUPhnDxqzWLixwpP0C
mGz5c6Ru1KwWEctQ8YJdP786KW/ah7zvgnYv7No+AsbPZnP1Vcq4mpph5UKsfTWi
Q0j96RK87m5OsZndXUDysz8CDhl8CDepU47nh/0iTR34hCsfh2wDCupdbYlyJ1IE
`protect END_PROTECTED
