`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hf7xqOcpjvEQCu/kaOQ4uj5iO5YDKeB1MH1SjHcLeJ4FWJ8yvb3hg0NMW/5Mb8yT
ariAyDZMWPe7EqGwlzK8lBO7cmi1gUVrcBo3gmhpTUv3N9gE6LyZM7y1U0n2WHmS
lb6p8UbgT+3mly8rvIMzb9QQ+QVvtmfJ0Qiuk1ErzjcO6vTHHJ9Q0vW1ncAJ61XB
D1KsYSJXGXlJ1CcpQHuT9lHEa5MALLptoyTcsXBG+IclFLx9EJ8VrG24JvDlEqa6
qPZ3F0e46eZQag1napHvuG4DN7w8Zi9PsPS5LwlrYLPnYXA24wzWHPzfLB54HWRE
YIDYxsz22byMeBdp9GaT7vnDv1Lr7dM5UML4nf9EJe1Qbq7jzFqz/AxsZRhxK71i
o/au3aTPAhN7INfMCy3uzK5t8mpuwsNQIj7AMgoEq4tA+7JAXrh7WofKxrHGFg/v
xKthx71nATGRXLYDwYs/cmWRtm0ukwd0nWQ95yX74jEgDDXolr/2c/hRZ5isd4db
JpUeqpFXVxP8nwf6LTvMv4rmPD88ceEqDuwsmHmhFFnk4lvoVf01r9xs5/k9j4cQ
OIWdT+r8ksql1xXeBinGwFLGUtReuvIrfLMfJLXSargxNujIQFrhBXlDvypvYEOu
cj5bR6Rj7mKYpUFabllMxKPR/cgZS3EMVMd9G3XNVM0A8F0hb/UK/jVMjRJS6j+3
di31Cf4rIlb34hM9F2cD5HqQYquL9a9zIf9wqV67mFmg2p+JEJIVSOBWLULWWCvY
AaYs9YUJy3lS6W0VHI73RoAYSv4q5DtgpIbH7pOn1ZYiEZeuXxvK4DYUUIXetbW/
4QADJtY/3/czGum8xf99Lo8QTspkyvYySuzr/Y2LudT9gT165OBTFz7n7oxN8axM
pI1IHCs6FrLX6+7kQ/PamnriF9PKCppQdYuy3D5oNqCAtETpYyvw26q9OqMwak4m
W0sIsc7+n/KSI0Q0ECwLk3mG4hW53G+TEXo6yM4pyB4F8W0YL1DimsWwP3oDOAlv
cuJuEBafnjIUeruhRLPGYL2kjIdT95oLwrpTVG/gshZ5OczbL2d8RTcxwWPW5PvW
0Toa4HsK/8aFtek5h9Qrgg==
`protect END_PROTECTED
