`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oml+rwVA7hy8mHxVoflx6RcpDKSta3I8gIE564Y0smkMTmyiNevtRe/tNVtwcFBv
MTwJT371bbYEnCdPAEpSElXQT/34B8RCYu354c9DktAxBelmKndywC480AK1N+5Q
HyPGhed8meL2sXGG11bYKRKJRgkSGzqgslnuMOI+THfCQT2lsrYzhtl5owJ3v2wR
Kx5RtZpbGK6CaFLNtFqvvbhfL5ILzQGxMI0WfMa4GKs1VdXMorgnrTi8zGnbHm2+
ekLka34uKi+2yQtG8dvCQB0HrYkiHbEQSEJQi9zbsIi0tl7MtIY+p0xYsto0vkg2
3yI7Fwh0eWmPENWSj4Mdko4bY+K7ZtQPr1PZ2svrJxD0D/LH4VQ8C+TkX9cNeV8A
WDHjbfO+FajNL034EfIjSjswme/xzYda9SuhMzLkuYQ=
`protect END_PROTECTED
