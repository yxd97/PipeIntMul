`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlxwwHayLRJlBGpskxZXYMfQ2z56X9Q06oJlYfaMS0QZspeqtDy+NrkuPfcRWk/K
u+z37UBFP1rK8r5X8rEfd+gW0Wp3gYi5pVGCD0K55dvTIfD45rfdpmWpb3PCpQur
eoPXG0xbEle+BipkT8ODz/EZLM5ucmi24eE12v99JIf0NdaboLFXfP/hn4xuElAu
jHeGBQoC8jvEG9OMtc9/xt1zVqM62oRy5wFLo2b9C5IU8xSBbqm+WcXwfKevnm1U
QcZimlAtDPeBOj7o9aMKy5EvjgG2MDCcgnLVWZ5Mgi8jUspqNt0o92O6nD5ChOdJ
nig5aJJs+NLRpHzbV6AWYnXw7ow2QCOtolTnvwxgsvjwcZUpEF2XFQpqFswp7n6m
XBhUOIH4MxKxSHWDFozi9XfalZ5z3bFRqwzGregvXV89WAFUntV2dyU7tVlj+Rob
puRYYfazTk+aYBF9ZBGkAg==
`protect END_PROTECTED
