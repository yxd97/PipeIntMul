`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vv7ASNmEWe/zji2802lTYmKbX1p959HqrxNK1H1C5eADACGcY7Z/eFujanDeneJ+
Yly67pe68+2GAU2jqkTHEpi/YJbWFf9oLh1trAvKPdg0/VLxl5YfVUD7NDV6chpP
Hp516nTdIZOtzbIuG3cMK05M4EwSnRp5oiYpV2SUNsY6lgINFtAMUu1tVLtvaEfc
EjR0yM5I/zuIG3pGxnGRJ9GfHMIW7qhE9BbJYj9WaV2hxZsSg7fOqiKtHYNcs15j
NDXeltcr9nsH/hDNemlkw5OmwxP5Sdl0zqaqTgqaOfxGSyjazvdeT/NuxRRU43+m
vw8CnPmfL0tvwUnRgBcnI2x0xt1xbemIwpYgROhWn3vbvNgj42dPViGTWN1Ymtmd
ENlDvqAsEc+sipPW1FCfnnCOwkVvV7ffgBWspXRTUuwIkRarfaVjEE9rjT1rV5qi
7i+/QRPKgqrcwcVQ3X9P1mdy/qs4ZMAyqHspHyiumAleU1ahhcKejV890GGyRq4+
KIlkSBlKN2hI0R7+HYrekUmdDnCqKP/fsaYwTeCw7u6raIfG6FuMvcuAxyIIuEAq
xrIdu5f7rIr5v8oNUfDQEjojvwrq44uVHvNL2v4cGXyXvdKSgRYd1OwESXrrGAR+
99+iH6l64gEO3iYwXY3RvW9xRBjeAUpqedBKyih33m1O6izDBE3g9tmDd5bN0K5y
lsoU7PNzREJTlUlu6MmrPQvzGGtgq7mtHCJX2dOoZxBpl13aGPCMbas0qsLRFDlD
GdLwGvHsK116M/+xSRfn3K/7F2laNQsLNnlpAXr6Qzj1tfXkKRYc/v/Dg4pvABbg
Cofvn2IaD5NXxwmBqg1h5PFaN2Do4MexmatFupqCwgJGX0i7qtvqBwdYt2q349oh
hIXOrNLGHNDbBnrNt0XEhoF4xBR7/n/XrBLxxMLWwtwAPVN7b6oG9zhsPea/ATjv
LUjYIQ9/wQd4tTR2wNibAK5YK21elmNomAXq+oPoWrSTQ7jnUnhyuBIaigf069K3
E7zDNE5ofE9dDKszENQNkLclRfcmdi6PEiacEdfbNkh/ORFEyu938+TVQmyrh1rf
dutDYmMj46V1Y7AlfPHW37jUCQoxlP06whea2VAwfgvciPxp0prq/RYb1Vlihj4v
EMOrG3Ic2TJgb4id8t8Jjsk2ipPjUhfHhkvfzGlqmwQXeOoVkIeTBXnpsKSkNctb
0qi49NY18bDl82zi/REgO/Y42HNd5YCzIH3gE3S8S1EMZ5oo3faQlkWsYz3XmbfI
byPf4Hjb0tWgG187z+YFcjGS7aR2o4h8+lxtVBRlV1yay297ichewAe/lqPxnptt
pjvn0m9yiOoN7xZTQ2pTe5ys51mt0iwgm0vZ9v8Zs4C9M4MYzXTnm3+tZNxuzRVy
cIBEIlZM2WPHZD9iinzUmGXXS6oeaXDfhf+BqSiJgqvTMGqtEolJ85eqmgn//4eK
`protect END_PROTECTED
