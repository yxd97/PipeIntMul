`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3CrdvIBaTbqouseVMiESgybo8ZaaG2PMKgnxAj2JCmmODW6nYCFuFVs7P9mQ87IV
9bKnNLQkIkmJ1Ss6AUt1Np4sfU3SKLId8amfmQzsJjvvKu7bngJqxiBIr8pKhoeG
/Owycdw7WkojRQkDB/TZFA/7SzNx7SpSd5NzoQBzsoD7D3pdupLiBEsBO0+JJ3Ok
WS4EbTm+u0RUl525UMAvswjcPg+x15OYXbEhaS84eB39lOoq2/PSZK8k5U9jaDs1
LQqC2zPRQtCWX4qCwhH5AYfqhBNDX2jVHZO4vhoq3DER4os60d65uLwulODt03k3
R/gXVSFTQGYDUtliaot6VG17qD01an82+EB2/Xp7Tsytl3CximTGU5CqsMQQY15t
M4OupW2pCV8Dp2ZPdzriHf/BqLV2Par6wmIbwdDsOZiW8Oz8SpBq5c0HiL0/fcAf
mk5ghSGbtatPasuPLDlLtV0EIqTNM5Oaeu8VfRdiJ5E=
`protect END_PROTECTED
