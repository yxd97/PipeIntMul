`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCJIwiPD9S5AfxhU9RYgm+unxbaLqQIcUrPouRtMMDbNvdPPMvqo8MaSUsunhxjQ
gGO7kptUmIzienHeaKGPa8rEY6/gfSuhUvzBgS++AQMa76Hb3Zw7alVvTHLBm+iT
htxh0iwqAmw/4WjvDBYmUwG2PI3QQKZpfbgc9tXIV7XvltKqiKeYeopR310TCZQ2
KQXtm55z31ERoxjx7CcwPPUNVhu80X0jm4stbiZxkSUbxf/yroNV0h/hzpQ1lyAa
zn2rFGum8Vr1RqVsy0DOelJqINCQQtlL8Wulv5wJyTGWxqa68ppsIZ59K1ZRXazq
Z/MrrUr672MnIdiEKMMj6w==
`protect END_PROTECTED
