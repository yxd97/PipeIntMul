`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Eerf96GAvQFHFfbqcgdxZw8QZn1BPon8dGS+Dr97M6L4itn1X0HFJSsITzfapzu
NjTiCHscb7CqY5LkjUxEDbTxNj/6AvjDRe6TnAgtRuu2O6D8JKm3jhpfC8wkAnZN
QokXegnJ4g4adp3WyyAJC3PbTkVQ8qElTd1n3rbQkRMw+P2XxDxGBXEqHn9ZMj/1
7vWH1ltcC2GXfph+0ZcFmpE4OPhlpn/rUb+wWp2PvIXcgr/jUAs+2y0fJAXj+e7n
DY/+NKlJS5XXmr0hTTdq9hSubU+b32n65c/bem1hwqVHx/82yEc4QvKZCfjRh5/K
yuDY74euQZjcbEhP3s8WMoz15lNi+CMgLxfUqQKnhpSXhfWV+7Su+6cTEDtAj+7K
cRNri+o70UHgDX9f8sU5IS66lQFqb5XSJOvWXGdHp7Y9JpbAFU7u0OwCGsklo3nv
eQsQQUz5bnvpmMAnLQJ3cRXkyBxtrvpJBtFAnHy1CEs=
`protect END_PROTECTED
