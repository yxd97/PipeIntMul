`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V20rWIrrEDLZXkZ1z9sW6usgpoFE9YU8FNd+zcJ9uFgRp5ok2J1m56sd4LmbTI1H
f8sls37ylvPO7DzEgs45k5NWrgV2fzIfxsUajRn6NcGNPnpN3LaLIhBNbFHLYW4T
TjRwO2YCPOvhDeoZUoIug/Hzqw4F6L2n3VhHxsEflS0rCE2uij3fpin91W5rSAkn
sYcVe1//yXRq8guqHg+CA45bZcYbILMaGtB2oGrLDtRJgM3LuS91sMlieq+bw5FY
VuYoWnmUn+c8UOqUjHw54AGH/jN3f3fLOSaGj/uXVT30Ugg9v0yPitRy8CackNNr
nJKIDgNvWiXmf0SPiPhi8nmxSg1eLC0ZcpN5AhMZNMEHYM24bPxn/Wwd6l6S+2Wb
E/cLAk2W9pbfpC0E19yZn48GjwkZdze9AGFiyRg3W2Xc2Qf1AeN60x9pRmw3wmKF
D3TwQ+TLezFmqFRdVRNpGh9GzplcQ2DtAHoAV7IO7O13EJ6PrCdNCDI0YTZ/9l9t
LXpywM/IPWCZ8kbKBzImsMeC7IcckO6PgUBSeFWXHz1Ks0SMx1S8wKe9C7sbYkjQ
`protect END_PROTECTED
