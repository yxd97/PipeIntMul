`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0L+SD6pwtfhbPgTIoRnJAN5kryl9Ig3VKAuh/ralpw/27cixUzGyQu1u8KCEgF9F
5IX374dorC4PDvRe82gO1xzmuke6WYHuaelWrZnuQ8UD90h6LqQtT8E9pknqJ7M1
gP7m6mY9xi7BViVzK76ifTedei7qgd82Ux6DHDB/hkPv2nnjk+m8ogltIYbpZEf1
Ldm6STie3Xww/rtkaTSmMsGfVW6oQSwvK7zAWdUVTVSqymc/hf4NzWz/UT+RUArf
MsWr2g4M24SgytK3u5JFWQUyyq/L0hS1t33FJ/QFQToYUiHj4BvIhVknQkrd6Y+a
`protect END_PROTECTED
