library verilog;
use verilog.vl_types.all;
entity x_dcm_sp_clock_lost is
    port(
        clock           : in     vl_logic;
        enable          : in     vl_logic;
        lost            : out    vl_logic;
        rst             : in     vl_logic
    );
end x_dcm_sp_clock_lost;
