`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bn+MB+F5PEkla9WJljv0lBmWzkvatrhh9GVAp2rayIUfXIi8tpYEW8RpF3LG6czc
IKf8ybMwU2zQ2eE/2Err/6bPc4+j7Get16bdS4XKFP31rbEm+Dcurs35ia+jwLnq
byVyb1GIf4hehi0iecLaTZAmC8TE9y4Dih3jh2yp+tpCEXcgYBs3/XxxRdTbPmYE
NjVX/aYtN/kKvLtQgkSFNx80fWqNUjSYQJPJLZn65uAMy03SCAEbodCzGbVI9O+N
bcLMzX6ZcLpOgQBsCqYmoq5YqdT5AOXqPuyRgJrP59kGBXPP+W0jl/l+bTBQ9g53
p4X/yfO4rcY3ZSr/T9uidZYj2qw9Qipz8u3XuiHKeROxK2/ye608gS5oBOfM6dVk
MjkncRbi7zbqz+Uk0GCZ4ML7cjXKQSJpf9Y0P7Lacs0=
`protect END_PROTECTED
