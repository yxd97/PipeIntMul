`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3Qzu5sSvNmiZ+z1C8nHIIWLDyUw8SoWX9FOY4mtWBQ721jEvGeu9hzrYwnTYef9
4q54ptykAWCON+OtKg84tuZL1XdMyx+CniLGsEMtZu+uujk5g6ZcaQhkBHSUExK1
SLTN68v4209ciofq2OmKQtiuJIw0+HwpXLNqtzlC+Uk5CUkL9JNV8nOgzr6t1BRA
MXpOETu9mfsXTNzEK5CputZ+XT4tZtLFiSZgwLxZZ8yfmneTgyBqF+Q2/qkt1U+e
7y9mHRewyhOWGO22nCRrLHRACXK5ckdjJyUEFMQhD6sg/uFtXlbnn0vmujaFeqqH
KWsvbFVMZb/DvGo/rnuhk3LPgTR59rQEIcQGnIKLgpXCkZtoCoyhKR6XbQEGyY+1
1JIctojKrY/xrBTVi14ERhnnbzQbCuDWA8pUxIclKQwhR+TJkMh/qufMLRBBlchE
KnSIPeUNIvOekqGlxEKqoWiCo7pxLzvl1ZkV31OdwwDMpDSn3Z+k+Wxitxif6kdy
Jljt+nRd6NlRgCA1T8uHLM0gu/dX4Rb+s7mXLal+RABkGUBfa7krYzjKns23LTu3
5ONZ2gegBPt/Slf+MSWQz/+tNiSw90uQYIJE/XCD0N78M50StVmmicURTOCCpS7V
9nLxSRZoiks9EVtF1LfvbgACWag7y2zrg+0sMy7dEVcjQTqOV+uMqI/15YzqeoSB
pZRi9NXg7B+QhWvyuWWWxt45S4bwO2sxahNJhh+r/J3oyyMbXK7x/MlaU/JQDZ4S
oYdP+MHXQG1wiGqdwG6vcgyl1PLc5A8KoDpSDXykPlQbgxMgWZMbnybW3P95jT5C
mnsOQq+78kRwc6hwQKmY8aaiiSJk4o40tyYp3gM9d60alrg3/4mKozD7JFksB5LU
iipxj4GB79zqdvCAhWcORI+BDiSp0t3Y3qc0nR685WfTzNL77ePFX/vXvbcFK/JX
6zjcEw6ulcwbQ3Hdwd2u6c/0VPGJGniakbG5T44iwOJ8+Jcty7qEvaERgRR6zqF2
vIjPdPwSDmClLbuy0d9JuSTpkNERimH0BNg/aerHs6x8U9vjoFKXAvDoFkN/89H7
zJfMSwJLNQPVNLJcdR2XcjXKNi5NyvyYzsQJPmyV+hS8MSQlIr14SchEhU948IMp
ZSYvQxvWwiAR8lOxRTL4YrwAENcjelrybg/dDvNguTq+90OsmYYyy5lTYocfGzO2
1lHojNjeiRc/pH/DvfjhwhxYm0thTuzJ7qpRf5aG7U7asZPwZJB4b/5WxmbBp0kL
hjcqSN/HEFKgGaG8XSYoZQceVJNfZhIcs+Hx22cqonCwDiWQAUND/9Q3KW77piA9
Hm9CB9lnMg9YQY9RMRkx7Q23Y608X2VlffaRRbOrhnvc2Y0+b3QiZZmI10CLjQmx
/YupCDc0Objs0zCHvD5PmDLmjwcFUXoTAMRdl8DE7yMfgJsZD+VVfyL4QrvU96Sp
rOeYkpVwmNKJCvMJ18PcmmpeHVZk8FsTB9KxMbrCOkRAQuYME8Vb6NqbWlQD6T11
d+36lxB28Ka2bdJgnK5SXIGdIQD2PeTV66OSsXKvWoNYnxTVpl7FypPcCjak9/QB
r+TwU6RBGNhWAc+KbYfbYBbjocYkk7tBsxhACfbjWqy3IslDu2/TnFiqYdOPO2Pz
ofC0FKUGqTH9vn/nYWZrM9BMOc6VCQChY4A6Ve4IKJDDOhnx13NFLHKTG7MVjk0b
/Yz/jJohiDzAIEXy1tlBZ0ZI422lxmXRDrfVoy4gmTCPHyupO3SbLXcZJGEJv2V8
E/zPw9WuTv3ZhtK9jfhpJ8k2B1x2ERHDVuDT36NIuzp5BN3K97BjVlH+d4Rwh6ck
FLu1oGFlkNZtPHbyviodYiumIE6D7IA+D0xS+y1dZvV80p6gJFcEjQlgh57Adv7m
gwYxKl/MqBpR+IxtxuRdQAe5cl7cuUONjXwwzTMzH37A0ThsLv37NxP9OfC4YgOr
OAy1gP9/zzouptv4azajvpwI3SCsXrWfsviFewUBad33exjulQZwF+EbdDj/ODsn
V1xytYVCB+7d+kFiCvn02g==
`protect END_PROTECTED
