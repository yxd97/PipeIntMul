`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70ny3MZDgpBHDV3zmBOYT3CCChB/Ql9Yz1bSacCzUaZf5hNg6TIrciGo6UqNmXQV
rxkitZ+8z6LMhAcedFvdY2hhL4lTvK/LB3nI0tlts2ZFGBSlOOXhT5rR9pkSFbVr
3AZdX4Wnf7CvIqg91NZi4MtnPFGxDUfJaavGxNoGGnru8vMy4MFo2cYriJBNtUrX
lCS8Qau3IZGueylA8e/Mli8DRCsokxpK+vvxoPsbQDpE5of9zqRwdHS0m1E+sYhx
Y6n7tAUfGBM4W3PdjToMv3JU4Mb4oaRNl58WeTF4Fmiv4LWY1/17VvjyNCUjlQXa
hcNwEdXl6IWtT8pmG4sw950PLC0Tnnz9L8rENYNhhrzHFqkQNmb4XuoYLVzi/tZR
WPVFDjpnJSlWFInGSgCFRNqnZCaoHV2FpyVu2xEwHn1oz99+IXUfGl7MndFXy4WF
FQr4si4ey5aT/FCro++bz3K9Mqxy1tz6RGlDa/qvOBVfexnFiB/bjPaopTHAP2t1
nx8oB99CGzlLLL1RePbFSF+IM75ww5eLiDxxzU07pRwLOQwo9tVakjwuYbvRUUly
B3+JJ3jO+A43wYisU0MfjYyjbX0RM6j2B3YOLUxDU6y4jeIpXhcXo59sIEioxzW0
ZkhqWJB0BX4L2j9H2yCyZ29SUn8kLrHbeg+IG3ONEPHaPv7z5UHsg52hVHSY+Tum
bS77V8ErO3CPOgHKRoT2JY8jTIkRTrVyofzxsqxX96i8Y6e4xvZFQaYLFZsZbE1p
ov9O/Nto5nL9AQkVMePMws8p7CMSGkoHzQ/EBts/P/jcWpUBipD80+4O53GQ0n5k
IQlzZtvY8BeXsExoRjLrRre6/HnEKRVIt9BeFhzcoMoCh3PthT+Cy7VIlGcc4L9t
yly11ITYQ183mmuDh4a7O4+snA+uxSAF1yPvWnghZuylOfGguAUmPjnpZVCVKSym
yGnhP4MWBxXt73Mg+llypmfyI0Ztu0eTeKZhnSTGKw47IMrADFkodz7aICbYf2qt
7IwJMSHitEZqmX83DbTrsjzF1SEhmcKhvtMgCDjayHmF7OaI3iFpF8yuuBe7hqRa
WVMbU/CjN7SA0g6bJVdGPxQnE0rcNIqCnvBt+99MscXNMH0/KlBaUHvErK19NhuR
OCH65cyVlDrntMVJ4kBC0lywSyov2T6bGGgp7aEUvM0TiqSa0STpXDo/NFBtC68X
dl9PSVvl8axqFFQaYA5WYVM7gcoxXP1nm00jck5aGDwOdhcQqdKzFfxyBkgcNcv1
/LKJA6QQnIrEvIXba4tP8WnU7L+2LA6go0yUo+yzNh0CsVxcapCvQqR5LZJNC5BG
MqZ/4OkOEnEr95/NHsNypcA/gfPIBxfAE4mi008e++rVbL0tdHpudspIrFiOEcKV
1L90+PBOoSdU4+0i7cVFOqTosFVoqUNy+/tmLhztQVgiVlS2XV/KaWLENc9xKpu/
O29xZYHo4Z1kqWD/9MSwxFZpD9XaJeYOTOB7UOpj6PZUhFVbvtr5NpWutC1c0mlP
j63dtILJVOiZxl2uYzM2pAEZ1ns2QNvrjTELtJz85dMW2w7o0bIQuh/qTAzhY57L
qUIQqb1AJYsEBdRWVYn1V7X2n666Ys0HUmQoo+/rA7MLPYFh3RYAapUJSYpYjIsu
eIceKd57MDKWXhU61o3pFC9WFexdqfVo298rDSnVpnpfsFcqS/pKo2XkwwPDRGdZ
JMdmTmni4SsE92VS0TliG2/PQUc+b8DjTRy6vUZ2900iryJhaWyfbl3poeHmg3JK
xrpf04xFkkzYYuRgniXB4wx6/gnNrC0l9FDPFWGciVcCpAbAoayO6jUeJplpTyLJ
Msw0TKkRXmjnG6CR6dZA44xIqXpWOGQtawuSY/jjFvvX6mJO4UhBFhlSLqx3dILT
FU5v9psulE4RkFuZY9Q3/gbEzRplHU0pdH6+p//5aQfluEWU1sXXI51Hr9NmUJgI
9oMshiKRgVdBVoS9WrtrBI8RD+XI/EqkjNVPbKJqIBwWVRjmps7mkm7tPRjcp9HY
PZepU5Sr8XVr8vlg1F32BnblNixF0FZvlw+BCMDLQLcvzma6u+Lc2xBPiZl1p15k
JHOV8fgJk1fd1v8hT4/tCXFBNjc46BubRyNnVN2YfufgaE3gt2vPho7rKJZeQsfR
oKBXr0TaQF4AzA1l3N2m/EEtizFn2CKAqp7UE5ltXtvzl8fwWKaHg/e2VOoXPfkV
98ChXgi4Y3iG4Igo9xKK92IuSebeRimTCBpaHL4TiTSsYcMrVwyxjAG/p5nOu+aN
dzc89FtxFpmHxZMe09fMuk8/LOuexGeEfc8trZb1NqKUSH3R30rERYH+87zynKW5
KJwWzyGBMArBUFDsPn//OXdxOMWhx0XRTtyuCQRvIcnsBWkLe01HoybXE5KkrmUe
MM6tQniAtab63D5OwAItcb+OcAYZRwCaWONPx4T5klEQ9Ieg63zC1WkJmbAX57bo
uC/MQwJVzVpuII9Ye0WL3wXHTE2oZ6EOtLXXRhq2aCntSNhrFx/m5RpdLrhqfjmQ
HdqnjU+v6nF+5vUOTbAJN8icC8FDFQIpY1eCKffIMK3pqwjH91/aIQ66B95HynCV
FQuy15mDoEDYeuwsQfD+0uPt41LjhrWjry+9LFsG3BdAQIB1J+FIjm5oHYV4d+rc
iJ3B1Eo3NqwfL1A6BaZH+1arQIPUpX2C0doFQFExLwl0qA8QkQoRHOnuR4Jgtb3t
KYCk5576ieTjc3LE2VrOLl1A2LV3UEaoRgUakD2djvx0yIV7L6h46rc/q48LFyMO
EcyZcXhr7irWzj32Nrxwv9mXPnmcMg2vO/5j4FuPQt9nRGU6S7jQGFyonf9QarVm
l6HF8U3x12DG8VuL+TUaxEdDCuYdakVG+Zx3xgdd0g/+scZIBxebtg3Js7A/Y4lN
P1V8mNnNPkqdxVeILbxF71V7xnolzhhwGJmJ2mw3B7RFkeQnrdOzkAThGR40Xh9f
u7s86qKIb8VNRSR8mbxIuteYaT6f4pZ/NlDkKOEf2SUNmo2tyDevqooViBVyHM5o
EtVa0aw+rAcq1O8j1LfQvO4boL4pjKgr4JWxk6Lf2V5K+W8Bi6hFw57BtjUSNmxV
D5+CFxXKQfgBza5VrzCvwS6JruTtRg4Z7X/1PhNN8xaKPsy0eqY8Iy5oGL+gNHc7
hP5y8TGhf3jRcHWz2S7gXBaIDMgzaQrdQPOMFQNMAEr1UnHe9HlnUUCjSuXV3DZa
zpoWswmUMOkgo0F3LQgVlxPVRTGwbab8hc1kryVu4irR2XD0c6fQgw+Nuk4ksktX
wHIO0oSzwUA7iFMCQwfcucr723fiwIq7A5lSIgl59KpOqhFwmBnQThKmXOL4pMhY
IoZ/tVIUpj2lKJ+3itplsfCGUIi+0w4Bqq+g3PSiaCjl/YjinfOkiYRZK1r2SNve
SYl/erguqxnJ1SqRu4jSlq0VJfLzgqEUkrTUklgwGJoFUhvelAPOJ4q4rZaYU5CY
AGSeKrU++NV7FygXUGPFrtLgVdBIQktH40zOESJarPaVrQylbgP4yIARX/h+QDpT
Tpn0FUX60yTYjwYQejaHuzbVtyV8nEDaVkymrdZsyTygWBVeIZNSy5y9HI9tVGTX
HuJezYU9Fg6ONTaeP6I9Le4DnPwHX5kS9Cwodo6NjdO9iVZMr7GuKiP9UqM9ZNj5
RztAN83BFeh7eeOHeq7znDhNsvHqzC4rqDjHhPP1xmbinfI0PNsDA+kta4gK3BZM
XenuqOPZT0c6YMreI3Ri2gkPqJbyQaVrj8cOiJ/B2Ll/Y03xWj9EJirTdvvto4Z6
l/7JjMoePhXih0yFEXnE8jNl4Yan8zFkm8Wa+0UnIBqYaz3UAWhyQuxi+vX+KsSm
a8vVk2gGEZYJax7EdRQvH7PynZw+LM+GZgnt3dsJPTr1Tqz6j5WPJWh4qDY7dS2/
Q1BozLT/NMl3+TooRe0fFfh9Uz7vd6V6qaJzdnB/FH1P7Kyfhu5Y4jX8BWjflNQK
Xthftn1bchBTqpTizIC4Dc/j14Pmhxad7Z8cBdlOxjx+HP0SHe3B5y2AIN47Ru/l
d6xC2zG/lcmihmP4VLr/bV0Bh3Z/PTusw8w+6hYhu9+F+FvVohXIZHJWODIuK43J
+ljmExgzYgdV/+IjUmTQz1/Z60beLcXnDAJVIsUUlkC6cz5CdHt4O77o+AxgS2iQ
eT5GrTP7loV004p3Bjmn0cA+rh6C4JIA2il69jfvAyYrrqIgEa9gritVmlQO7QiL
TkPbcZBZ1ZKrkZARiTqXveFR8MdMs3c3S7Byfi2HSXKYl3L+cOSkxBllDhioyrQ8
MXv8ath1TnmQbLu2IipIAcyCa1RYs44XnIemZ5ypPOcY4ETV+8jrp4vpxQZ+LHqS
Wd4gBkSWN8Pq3AT6ie9UmaNfzOOfKx4ssVZlYaz5Sk2qRnqAOyT32x8g7xgQ7Hyw
UglutEMj113cgDviZzUw9ukuF3HcllmZ9fyjwdnTqfuvtjG1Vgh0NzftYtYj7nck
mageW9WhPre/oPYfSnlgmiu9b4Nxp+mNC/DpbMo+Ipumz3Q7YfMqWih6hEW+WqSC
KiGO/bn7b7dYLDjNbGHS1xWm3muR6/OvHgVm8KqN/O6CvCX0VdqP1oVNhrf9J2nT
1HVoGG2L9wmrntYFNBxzGcnk99Rcq3OZRY2Yl1twp4LYA5itQweSsXuDbwa/X55g
usgkFG6nucIelWQrqxiwVAY4wd5xaJdk+ztikCtpVZGUntleMyzlrW3aVOM0bRyO
MlJAbAWVJQJaykXcEsj8480yrk6kEYX3Vv4zlpw2bJMBo40FUitIiE9ufeUEszyW
nwb+6woWnP67huSR6flpylGi+g2yIYpW4iRjenPkn/i+GGaQJT3EuZIRD4Jto1OG
dqtWrPQym9YE9wElh/V2W9NS5V3tg3NcnngDddo+IKkdJh96Q0Y4O2euapwt8wFG
KSiP4I3LpLIx3nrt6HDfkh13o9JMCdx+cfrO9UOsSSjPozkAB7AcnXdpOwWIXr/9
Pd5Ixglo3EAAz5MGeVRQ8NLfF4GjITLFuwGaIag5wCn9K91tvf+xN3jC5joaBOGf
EF4o3W4u6eCBgVG2n550Mxu9dFKJYt8llHOKQaOCLFsqPIpeB4D3sbbblOVM8g2b
BoMpmrivq2hgQnQ286NQp6jrK0CC/nsl7hRYMEj9UxhYbWfxAdSY0RG/Hull7n02
B/SVGvwNttjAAGI5Ps+cW2YK+wsELmca4AmoPL3eQTwj79MdZyyhhy/w94rxw1ke
7sdh09bN/x6DG/lUJjG2DXzxwT2hDpIShr7tJsoXpFjCodnRjXcE+K7aPamL0JQ8
2gymetbvWN2rv9xRToh8joEB4H5I2Ge20vtbbBo7WVWYEfYc/LCxEJ9N1+g34P5p
iinGl8wqFTSxm3JhNUHq9ZETpxxdwEJ/6zaEs4HIG1TE908pI4noMPtDOHHWkvFA
BLKQbtQqRqxNXZ8xmlGWMx17sBAcT+Ttb8lqaOw8S1i+lghFEU4LebRwzrjVmn04
xLAQ4+8e2qodoSidYTBuXxrCkVXr8Y6sgdu9VTfEneRfqUIdbsAQeSb2SgORIrAY
sFxejYvyA/wmcuh8Tk8u32Y+YgPHFy7Wg5oq73yvbv1AxlYRVFzoBVw3l8mZqBqm
k+I6x+Ejfz53NvRQKzTeZlQfG1r+qqxSUVwLq7xQ5DCMPs5G66fq7z8hp2PzM5hb
UUslWvaGm/e1zf8Ep54O/oXDONBX6O33L+AvcMN/p50ZWgeVpJ9XRgZE9/FlHeae
3FkqxlBHl7aGzhsYnK+seEQSwmvUQAKZSDKYPPlbcwxaf48OWpQkdLFQhCrPO55u
gVXuwQ0thf8I9OGHGOuyCZL+xWJcsWnmZDIuaorUl4hCPj099t/G7iv2HwWNMOnL
0TtVxOxDNiwvz3xqyCFM1rQnPucLFLdVsq3TBtyMqaiSIEUrHzFGMoH0EZKkRrmj
+fUF7IH7+9jzrEu4q136ocTW/rWQwO0QFrg0OainTyaLUnMm1Ny66Kf2rSHQaUIG
kHzx3i2v3qR5ixKdurta3bIkG2gR5x4PO/kyxluTDO9+w0GwJxM4d/uQJcrm9Acs
AKDvcm3Bef4aI78yaAacXZNeFnC9k8nmbMNfAfYC6cfpKPqPjyCfc1v8YoX85iW/
W/41aashk6i2DNsWhrmewQlEZnerNxU1YTHP4V0xswwK3rdAIrC68oO9J5wYmTBx
Fg4l3fxLQMYKVQjV38t2IWvwuJ//NkOon2yLyMt85pl3/KF2p4RMZuI1rHutoZQG
THxkwAzNKVK3Q+ElXergWS68uYGstG0QoSVURFtBVnuqxdy0OYabDNvvsvWAlzWB
nriU5mkDV48Lx/D9NWfWocBVK2p469pKtdNat/zU101Pa6CIpE47SBHQgXhIZlB9
gipgLrvoTB27kgomwAJc46qXJtFHQK1sT5RvatyMTwB5hY5+Yjz9NQVsDivOEyS9
IQPf8I4b86NNPhD8cUNHLz7tsY1HNIhOD4Xrr0tyKgc7kAFuME1MxtyHKEDYzfzD
plcy+JDYhBDEhynofJ+T/AnZqvbl9gdhYC8+LZKeQTdQzNvVS1UBDcesLHx0hSYk
hWgfbL3B4sfmpG2DOcxgHc30FE/XVEDNTfJz7QHKX1NpOazvsSivpCxiB1A/CNUJ
PUhIO3Dtgq9VRQDcVYSHIufUJ/Hr1ITYK7by1oPUAVqcgpLwKKzwZJMO2AzQIiji
sTkZeq5tadHKr0zTS/nBX6Ez809lMXpsddR+r2GauFV36dAL09pmWZyS0Aagj9Uy
k+7hkmHjTo1r/pv+s9YuDIc2TOc9OpaGT5Dy8kWQU2gHsyHDdERVijHYIK9eZ/S7
EV1gl3GqO/pz04kicixdlPG+4buz51a0hlweD2G7jhjxpiSWegq5/TCDFoNV2a54
SHSoI/H70gL0oMY2hKF8JhZPm+psQRP1D79Zc+1d+P6DOZ2QRarB2p+XT4BMLuAV
Fdt+0dUxyXlHvgOydi9xi/HVHv/mI05BJLrFtyL5A/WnHuQxymk2aaj2WLP0An1C
mJ1TecD6BxaG8T5fmvg1591FZYtjOvsTbxDtUuOd4BgIoEB7ElOdg/mOswkfM1Kn
HBQlNlCkQ+QAyXYN/VPxVtqtaJcimJnivPapysZpG+AGRmyqBYaiiQwR2wJxumRl
DgP1+CmlDugewFrbWbHo5x9V9B+t1EUy1X3G5290G/YDijO9Vvv9NWMgofqKQ0f0
XcwTvyuwfvxO44Ryj7nFBeTGpX2Q+rL8RorHH0I1+30xQEorpdM9OGn7UFOApdfC
95hmAovaEtQrg2GvUK0ro0KgYxGxX+QlYkB+0wUDilwQX7vnLJsWXwgzwvkIgrTl
WRAPYvsOMtaSyzlvXOmanPvHzewUAL7a691J5z2Qixc/Rr2oQ2dGcLuWLFDQIEOM
FyP9hrLX8uZA4AK67N+uOWMATxMYH9Cdex/IsJpMCJM4b+20sZKP07kBzRYn7KnV
pOQ7QX0UufrIPEgY8qfCXR01G8XZHk5kChfnW2Mz6K4aKMIJF1PkP0o9ZUj3xkf+
IO1yKwZugqsKnoV1fkSTUplk+/rVxI7p+FPtA9mn+4uoIW6QrOxCjxA0Di5chguS
+AdhRJqIindsy/gdPABgOh/VLOzPBIkBkq9IUqys/JRsbJY9LP+dFOXYcv0miALb
ByJyyTis8Fpw8B4vkvxP7MMjXr3eqnC0Rcyntq7IpCFDutpptZ185Bq9gGlQv9Lh
Bv0SOp60oqu4SwS25cYiKJIDFgla7Ni0mt9IjUuBR3DVIvu2dDNSBTDDlHLviOU8
7UqcykbqCmaW63DlZ3j4mFuwezrq/6pgO8Q14OYeTe1xcXACOppPWfwKvbrpHfeZ
Ov76zpezXUQg+joPETKUBiwKhNwo/WaqTRmv/9kvZSjbWDKeXm0ogDcpKEUMaNF0
oR9epR2cu7+TMXPujASYVcNIugjJmnbduOLjUNvIRWapSUNuku5/65AH3If1QeVX
xlDbN8+WjYEp7o9FqtOKqtFfcLpOe0c7NaWvxx0feO8LCR7oj6v1jtShz50GqwLi
xqugieWORXJu/4FTfK1V/+rd+lrVd1xA7x/ePw/ElhKUpfXBX/rzqYpiMBNxn3BH
0Rl86UBd5kg1D3aogQ8iRyR88M/+dl7ngGgZCQ3lo3/I7bgrew9JuTEzzPnZKUKL
3Hro43NlAJYs9PQzlqdXNqyeUV5cT1ri7tULVJVapMpx7nPw9pXdLV8DdrL3G1Ce
j3oI30DOTC4EACk2SqT/a5owNL7r3rCBgMS/Z+pVfvOq4MI1oNv9K892ZH2kvkO/
WdQJNhwjWeQs7ZCAbjCIzJxdpfsnkHdKXtnngSdhmLt/AChG0Ijcr8JRCux7SRah
o7MFT3P3jT5fcBGc3eXs2Y30GcrvJ+/wfajuyLkyfNdBDJ0qcGW/WvTMj79cjKkt
STQ2Wz+UAZ7sav8twGBHnpxkuiivntnMTZEmLnldRT4YtO4A8K/V0ILxc/eDmcnQ
SSErjGzjevNMvKU3ERkHZoZpvCpquyO3C9pIhvN7ukEVFt9ipX8T+/oZRidLbHky
DugijI98B+yh/xrTG5aJOPJyI38ZJoGmzmbN6jKgG1DTvJWydrxJKLpMgi6rCO0G
DgggLnwn9MMb4mtUjdb4lKwUqcMxna8J57RyMISy3xWD3/7+paMd8puV3wR28fjc
0RfZK5saaW5u3ZBf2HWou9qYG/fLV86rans5/rdFDwtUKR+c1T96xhRaYfCK0i+9
4pJ6NZIZ9a8VX+3/b3a8xswFCKBJ4GMabe402QaR/gmY4swHWXflCEjzufDp9g3I
TQQ88+nxfx4yrL5yo0enehnGGYqkGzmJ6xoRiFUl0f1hoabFHs6o9/7zWcX1CeBT
WkmQSm0ECOY3ODCx6+61hODXehF+5j2v36G19t8gMRMKURIdydSUJJ4tfB0IMF7/
uP1u6hdhltOgIBJOaYp2i0KpYmRJiyaHUisH9sFCjpn32ozgkAYD/uAnBm7LHX+t
JbUIejClxQE/KTtf6Zjfcafmek8ycJP+N3XjHoiOJxPz0X8VmlOXUcrzbzPDpdTB
k+GfBZMVeRqUf6yDu6OsJRtzwUK4YD6DxMIr48FeaDpFefzfiyQE9PO7gBAGAZRu
MoHXKMoPiT7kby7I5RfS4/lyIPPPErZ4dS/armOMX3ZoIB1YYWURBigKDC2Tg+e2
owjmtK33b/4LF/vklyi0KOchBehi2DeYdOyMCkafiO1QE4j8W9J5WAg2YLvKLNpV
t9u0DmnByk9Ku+JQeSempvurIRKVIZNzx+PMXVE0KK8K3TD0TA/YezVhjoyBGWk1
skcZ4DY9xPWTpPQP5i3u8ClpmMSKF9qO0C+s5RzIImInzvBuUYsIZptRk8FlzOma
s344XjjpXK4dWrVfre1z0YZxCvKfaWG+YIdmS6ffmLQ40srRK3EurxXPGxXZeNiJ
H+gtytl4IG2U8l2/0p0nKozRzjgvmH2PcKfcLrWZrsmmCPuurrlTUN4LQ9kfivl7
YbEo6BDCBD0E2zCkC99b/lDDCV6a1+Z1nC7Nh1HJMwcUKg52Sr40PfzNwt5Rbvax
G9l+08P58evGk82mPz1xVAe0QGN+d4iQ4daZgO2urN5RC1Cu3tGYIxLhQWcAId9u
iP5LymZaNaObBCsntr+8Z9WOZknFUdaDQX60S92sPfO1HESPEXecMVQMLKsVEo2O
oUnPfzqgu8N0Aks7tWolVu7CfqJdhd9aaET2qlyJcHynUkCvxfvdGQ+C6ZJAHJzn
HqLP+bvYcIlab5PNTEbAiN75JGGD58Ak3iCflq4MQmMIXKJFqjaPEfxCG5wrwr98
MlF4DiPJI0f0H63b2g5lAuHD2seB+JmcKkQFHyf7HXYGj9MhhndYJSOOIJLAH1L2
jf5TVTE7hm2b5PfBpSJLL/vfRFhAJyqpls37mpxv9PcmTba90dmwaP+m6+Ks5qyK
Hb2a6tLQbNIupNCz+5JTuQ/M7Z6JzHJ7fQc+NYvzJozGc3SCSvXrv4wwzMqfSQjn
1oNpVkxoEtA7p5sJawcqqdauAs2Qcc4dzSI2/bvbHWUMGpIvk+TR+kkVA+0r61ic
86sr2VyK6UzlvCiecvPVHnOqiln4Vu0N001oajLgyu/txCqp1rPlMS5SPwSeTTF1
Ty3rpVetwnTcNDsGltlGvzEk36ik99UQzq/y44bPnQYK5A8UcW1Z/jsXN/1x8Fwl
Z425C+7k/eyYvmvGwgAmYW3BCbKMinMORpDSFzViJDl0usMezu3KWGjZnRELS5lQ
MS+98wzdiB6PMTASHaKWmPBKVBOm2tvTLmsa1hmE+Q0N6I8FP+Qcfah7WfPDxYsc
58tLGgX5eNgnuhbIMR23nqJL9aNfRDeHaNPQMFHtPOeSn5l0bfQgkcoBN9l7pOli
V/ncKgctCdlk3KtO4vQBFMQpiPfPj0M3RUcC6drLA56V5tz6wGrBnf+G/GtiAew+
RlBJEQ4Q9mSUSxZis11YzHVd8TrTGBWli/KLYat5Hiqgc3gHi2vwyqmkNgSBDrl5
h2u2bqm1y6IFeEiz2t37PRbzZYvD68PAMEOHujXk6gHA6IMr+afj1smD00eCJO/K
DWHCVpHAFsaU8Gbr6vXktPYvVjifmw+wXSQuoXPd1uwWa2PN2bEq9mdmJ5WmZjC9
8hWr6iPiJwkYCqX4KSlWFb7DMmUl3HXC6B2uqYYKJla478zkpIjCP4ZuIVmKe83d
6/lAmgSMIuJjvM9Or0LxIqcDVQznkEo6vWuh3l6iMohcjOouIltx4egtL4ksNjSj
vg2vV0OzDGOYKQrNhPCcougysZ/UzUvMq8TZ/kftIDf7LDyzt+JnuvtFOk1SSSj0
jkqKj2tTyj4Mq9ZAnqPTHNhH9letdIoCG81NZXYN0u0RP6h5xRq1mqQ5BdSDbaT8
XhL04GNJTzHcq2VT1R/Gq0iNChUjg2MM0uhrJgG8Y3xA2f2ym06CRFKw9ukxOy8n
9fqbQBAj8dt7y/2wbQxx6WzG2AVDGMFizf8cRms6J8jNPSTVedj93gjmpOa4Kl+K
3/IZTddlkywDTTczAyuap3czEvb0oozK7eVFFmlo3bzOZmiblapII2Unc8pLKWEM
qMPZntoSfRpyZe0oFp/+7ILKAz+HBPp+oVvPdFHO0qFJEggajuZFf3hYSqwUdQj8
SFansd6VL7O5wzg2YeeaBTUv7X3kpu7+bZ9sMoWgJayiG9V+oZ2AbWUhxxv7EZzM
Zw8TALNqcsrWicTi+a+13Qdqc1xuqCpybbCgPOw1nFdPSD8nHMQ5xrgur0iSYLiR
MoVwARijf14hPSNwy/7LCW2WmV1Q257bbGBVb8gKfjVJ34wN6ONSGzKVsF6xZiN7
8LA0Ifq+D2yGmvFHwXIBExkF6HoWjCwUVIBk/KryIuGvYFmTc39keQyDbII432m+
K1LU5VMK4KRVLw71G0SflxEmnuVeExH1XKszhzl/Z6SjSNiTPA1rLMwDDtIDfwdU
rFwz7mAEkPafJvw3XILgToAFTo81rSOfHGivNFiTri5GCDOxja2gz3ZLAIGA3pJx
uQFQbvi6DP+Z1CT035k4BL+3gqX3s/CftnitIuX42hfkIQ4cmdZ3hSGzNvYNQnCm
PJPcmG7V2yu/N/zLUNI6rZ5EeG7jn80Erw8Cu36q+Mk/YRQKYSZ8wNMRWikutigh
TjJjfZUq8O93nGHLuvRq3uxbg2EPYs2fFrmUWtwpPFtGr2SUd+SvCTZ8yoB1It5K
VMOlXH3knZvm0knEryOmw01jilsoSP6pCa6Fclm32Fagf/MK9WuAFkqDJYfPaewy
5VUcNu4ns1vrh/12tpzCCDAyAAiOhgvhXJ2dL1XilelsI0XkygS6fruMu7QV88hK
sv+X1uzscFANgdGFQauvPl7CSpubtO0PvRLyIfyOnuaRNn90oB/KkTy2/kBh3RrQ
pohd+bhqFGWHX2NH2d1XzGVAZhOCcDgXx+t/aZdEbX85W49RuFbbL80AdfQYi3m5
9WDg9Ou52+2d/SZcNnrjRLZvK/4abU352/kH1+JWAW7aoftDeWVlxMosWaZY7saO
03JcrLW8EhI5/wtJfPKv8t/XYGGfadkGiwGRSYczOzyRT52yMkYH8o/A1XNAE0+A
BYN1NF3FFXVXGxaGmNJQrUyRlu1oCysFnKKnc4l6cXIijBQZTsQ7q7RR4RRz1pia
bLNL6Qd6ovkpJ8G202x0zX19BfXhbfYiblAwY5I8vFQnQXu9xmol5bnMSUEfM+p0
qrfOygYbDY+3h4ESPYVv8LfaIistz06PzEOqFM8mb50WY1HIkrW3zzj0Z0f+hNgI
M2pOrYEgMeHgZZp+Kis+7r8KgqWCrEnsYu0arUS6zfWgDtdVJPYVWt7mHIyOtSgP
uMq3kaJTTteKZdOfwF1ppdhYueLzeSgP8SZRILLyaW8EFgoGx4QO/1XDDXwKBbcH
yjRC1daBSAx8prD9HmsWufex8Tmwaa/QxuPUyHTmIQzkgySfeteaq8sL/a+894q9
mRzUTUMzlNUY5BfCQtWGdYT3rnj9pKzZFLcOC+hUA1qKScAGp3FcEdEFFBooGCIs
9/Nv+i2uKUNmdniKWQWG4Fo9XaeAd2RzrJdDdgVhPnwr5cT9xJrdP0BxXnzHAuni
wnvD+Q4wz3dwRxrbSrzAFbEfBhSZGMmA8as43WQ2GtoZx6mRllAhkMyxwbjHukLN
aONFvp4qTIvAexJumvh+7yJLRiJm+7h8IP+Vfv6I8+T7Oin3zjFdd6WFQ0fE3Thv
rZQHYIk1dCxwMh2L3cV8KDkeA6+TN5g5EeftYMdmSfM3NS4TeA7H56noX3zyDsyu
2H81wRQyyc5oNPyNnybk0mF+ybEup4cPchYLlnTeBOabe21yT6/n2hojN9ZC2q9J
UY2nJkNrA7LNM2dTlGevuLsVa42M7JT/dtyx431sguzdwBhBJPKeKU2QrZrFghwU
mtdbn25URJ1E9X8Hx2zG22Lf6naoUPpLmQddmNLpzwtwszhmvzaTM/bMX7qs+s+i
X126d62qE1u+KsZ9zIq7kM7mCJLynea3Z8zlSs5mS76u1+dTi6AQ3vV4/Cngxl8G
IK6MIpDaxTu9J0YquJKPE9DwBBGN6F3FSv0PR9AITufd98tN/1ZMnJV5P54wW6ZM
+ye0E3fH+Kv/P3ZDe9w/zQyxC1MquHDp6Miqj+Z53oRETiV7jM+WxoB55rWYB6rh
j7Lpl7MwodWDfzMaJWs3BUe10og69g4tayDPnZmrmxSkA1YC9r8bdGG3CGuIKur1
ty4ujgGTRILxhrwJ11WeuboVKbz4nzW2fBnctdNn0YFwIQ/7kkf46a7M4nK0ZFka
FL+EEw0klOgDXFkIlLMydjGssKGuEfbnYRhrw2xYDXkfuJ2VQUfdUMdqoy7Pribk
sX/t5ua1opHBLjnSOJcruGPDa8/S+CptWhkvEuK2ARQyCF2PmuvUNpxAi/0h0624
hwnX36nAw1WO12O4MaULTkv9WHd5McRBvC1IPy6jfk3z8yJfOtqMInSrDwjQ4/dJ
qU+HQ329Z0tFZYyl3mrvckl043E3VLqAXrhqrOyq+d54UcxNi+oF7fVyLzXGybeJ
8P/SuO8+o/kpCE7jF0aTNRaAeuLLRVoyhhiRmGgZ30dxm0Zl1hHNw0WrXyf82PVQ
iPV1kDbVWBHRXO0R6yQefDGrFDCJRz6OpX+Nxb8SKqLbBEjlzTCkMvU5Hv7+kl18
1AahH1UTcfYFke9Utz1hUQae5WoOP0r7137p/lY+lUNabIXmQWC5udckeONpzcBy
JLOQpHnPHIigCsxwemNb+Jyi2b68OZ8j1KMWMLCcOQlRg4cH4wQgut2maN6sS2yo
paayRpA6rKJcSZ4RRs/WIxBAiREVTuDWYScshIvHGGRKAbQc3nnn8rWAgGgPg6i/
souJonT1qO7/xT765XmDhkK8KR1U5eCvxOuIL6DhAmxbqDPvBsgTrPTk9LKaEm8V
DdVkKpXTKABBBY+GajhNa71D8gj/MV4znzno/IJSkhGnA7v946tRlUoUjnxAeV0n
QYw862d8cUZOGGBeoL6nZDBAfdKXjjqXJzMQBwNMMSzL9D8+znOXsa2UXRYbY2YG
tsbZNz+4Ke2XoidukUCaMVSlo5+9g0QxUw3gtBVAVPlh074HVhsNrc594Swfcnfv
iCEPKFyjU4PP0Zr6/HsVuQELsX3QIYFg/ec1C53HkrEsiOl1Pj/CZtfCFrUAHpY7
vIzI0YlhMsKjZEcN2wlSTtNDrxXSD5i1nDQ+k9SHwL8L9hvw80BNHp4+r3/D8l1P
ujZYSf9O/jZ5GNQjp5Ho33AxW8c/VIJJXP2rUwG0rKjG7p70g1TBzw8Uz+Ghz+gE
uCc41V4Vei3L48KuxJFjraEYuadGBy5GrHipvoyie21Ykkw+SHI6G1pSspPqGygl
x1dQN+mHe8GKPVzZmWNTyV/COgg9PFHEpr1BMuMRYBp1pME0e/4WhZGsuGIk/6yA
n8t+TNzYpnzeJ/nP8wrg9ILeDItJC+uX5dUlPzWu/vLkWsQJGsQOxA7WlwjkANCv
7gUV0W9u39WboqaGMdiFrsf067H0ac9Gmbf0BQxpA1BqQeS4jZIAHg3roDIV7q3i
BPq3UWqCjYUKeHEUegEWh7lrKGlOUPScc7ZFj72Jjtv2go/cggl1BEQ5vjbrD6em
mIjXtx+Iryss7rM7Z2shgQAhDj0yyDLBuApCj4zPFKohKUyt83zOOolFXLsp9dik
Vy9wzJ92FHZCrJ3c3MXUGdWbcBD7//idjkaCnWcunhFLVbp/QmmDOmLdhaS1y157
hIj5YyYANb8ClWH6o+TmtBsfvuuwZ+bAF5sWKa08hV8Igy0BP+pr35GuFkHrYVCK
7H5wjAH02nf0rCfivi/VXIlxDKL6G3Ek6aYDlcHEob8pxBOoOZbsQZJs9jKx+elX
Yjs9d7EuFpoObOB1fPGRR79kgrE7iFiOi0Yepiz9DQG86IxRvs9o9hYNbIwJLMc0
qtWPD/8UVp4uWqcbrQg3PjsLxH3HTVvJjzp4FvKSM5aIVd2BgieDxPvHy+ez6W0U
MA2lk2ZthzdAOH/ZOTiN6YDY7srvKy9hWXorkOEa22AnHLi+sE8NOUrUksvxFHpZ
YyIRj31tl1Gxc3vplQU6eIVpVz+FO896oud6FrjN6+0rMgNVaKG4GRhYTGdz2y7z
dh3n/CkxxzN4t1EnCpF4wYetjhhuaEj9VRyLuy1C3k9CLsTWfu2S7/ILRPA2UWFJ
Y98410PDZbtFm7g+1yl5Cd9+cK1/DdWoHlC5BDS69AOajUqS9Xzt8pgeFnnEpKYh
HIwRcD4qMQIuYm6rwki0atUYu+dFJ4W/F5+B810wZzzUyATcQ0Ts8k3Lj4/65uwY
pZFQV7Z4MQUHym46WPh9IT4Vl+7ZPfUXj43csHEmDsv7HCAbrrnhCqhyZKCV5TuQ
0RnMo4EooGR9k+nUUJtssWMOEQVTtfnRmPRT98ioVv2E99HheD1DOVYYX3kyOg1v
vJqLjeN5NH6lgrn6IW/UGrDlQ0wxcWlwbZ1YAHkXwLXnmNj9YhjVFTTa9HAdznYa
/Sv67RKkTp7sJQr5j4PTRw1j37qaxhRIo+sA6i9SpqftjrVyW4HowEK7yD1yudSF
v0wtAU5SKOeA0Fi6SnDMnAtePcNhcJeZYlS8BYsX7lm6FRCAiSKZ6sBkpXpXNjB7
HCAcN7ikQkiO+woSNyVn9PR19nrXtkrrleC+4RCF7OxPFlF/BdB6DIeutJbQgJ0r
iK6bk2TWRLDJNKossHw4rGAAJN3dcXr3UjACBelY07PuTy68R+qFP+4oPOk4GAVZ
FANdlufs9esIAmAqL7qAJiYZL40OCv3gB64gizab1qHcO1RGmqdha8WsjeDenaAO
f/YWbIHv5yeObEWGR5kt7wCwgj6Wcp0qlBfFIQrVWZsxsWm5SyrPw+sZTbySzufL
DeEjOMZ3V3Kpi0T+F2UraO8W86iAZPk1xiUkwn6KIFiv5AMbpGdixH3NtvLAHUfx
mUyxUUoIrk8ToTPdAnoWA+F6Bq3kMmblf6qxmEycIoDS4cqCvXPgmGg0azEVUnfr
l0X7sd8/+SO647o0JNfKOnkSjPMdhBy0ra5UDPJkFncmGEV1NFgAvtjo3IeJseYQ
g7ciMgWqoA9KDq4+sF0fyJ8KWRZZaK5VM/UfKoBs3/BkMwqX7HRbpsLgTAPPjYYO
nqObb/s7JNd3Ek56rpLI689mJS+uiei1HCKnwQS9ZuuUCH36XquDfhW6G37cF0Fs
mYfZSZvEd/Nb2UqeJjYy5r6cXUuB8LXHlm+XwKSTQqaZVPp4Vkxc6MlVw48+nVur
YKXCcZTUJTa2sNcD3xylfUD0g3xcZWTltts9PplGQsquJ4+vPuk4Y/yEHGHZE0h+
vu8oDOpsGNzTV6dVxPp9zvnAGsmYe8J3k2GrgDwdrKW1sxZb0OMMaMGDnn2kqpNZ
IMohm5vOkxZ6tUeKVi8s2mDcrL/Wo/RMMJaw+c4MYFRroQseWqfoK3eNrKyIGp/H
kQcxzcx6xOzf2g5HB4rQaTqBtIIf2x42MDxxMTCCvLHFJAinvY89Y1imVS6V0I/1
+x8tI4pxasAkPznlUMhPUHrVN64mmwRhMg1WN4xX54aONLkDQdQTtMVlo4CmP9vm
5SIqDHxn45/7UQ9Z0l9opJhLQCjxpSdBb6M5NbJcPUeoSahaXW83auTR0BDtS4ss
HXhQc5nMjIwJvsqh0OmZK9vIiQqqr4Obp6XOKDLNAgG2c0J07j0YI1dk/UhWE6cw
DakTAF4WLcpSyvZLG1IcUEfkl3ll11XRNZ0h2s0ubFNREaKW/r/EIU/W2OK00vlz
w6bFqNoNZofFM99vD75GWhgIeAM3x7AFD+iKal9kpK5mckURLe0NdCwe0E+MHeH2
8XNYoAtmVZA5SLZOeeIPLKlrazbP4RkJZ6RBKLlANs9gIZebidd2M5ky/OGGvo+Y
OaRs9PLLGx6e9t86AiDVWpirnLVUWyn0111nrne/39D4ha2slvvQwUYoLnlkVAK2
zqK+lK4mk4LAz1uAVHsn0RiijNvlgtyxR3j5NkY+nQ9yFLeHg4j3Gb2BiN7U8SC4
8tWOr6xvVXmyXHeMJOeE53ugUNOj0XUwOhD5LQa3h32wxZB9aGCp9CR5Fl2YwW5Z
uV+K4VtW1MGCel31uQZDaaPrlGUdiydohTc4dJ+7wJdIm/tJVBC0PRtmkNnJ/Vb4
Usi6i+6a2zgYKMYcbuHaWEW3ZHxdl6XkZ7b1oGm6zRah70upNgC51odkSWLLqr3b
xPkInnKNtCqfOiR7JqKPytDugf9JF0ijJtxX3/IZAHfc/AEp79hr0/oOIWLC6e0I
Z2nLMVtnx0539QlUnw2RcCOsJ7xog1+DkL/3Va5NDRsI0leG53l4hTJNXCEZpmu9
iF0fEw1M3LQZa1Y9L+3CKEz1xAmQ7fDlIAOf5OmX5wwX7VPV5dx76XX36XDPlFp+
9MSlYLeKIdAcNHDGpiUvqCPJfC8IcneTXHQSzMki/f09rEaDoTkCd4AVY+Njq+FI
F81o1tXmz8zGpHqLeVZqhQv9gvgLcmWy1gP/Mb8Pj2yIWhfGBKTMFIt2UmNYkLg2
U7tWo6OZCbG7POBN/5WEgO5DxRB5NcWNGPXiAz+eL60s6RIl9T2dfWkWJcVVZS/l
82/UJwx++oepCMPmHpiFKvPq4tgkBybUFGoCZqejyd0P5/q/71/PDEcR1xSAmOkN
cfyS7TaWGTRZdcFSKO/Ja3rGRGeu/sj9vo3KjH+FFt4hk76RTReFVUdueTvV/YJC
nyAE+PKLt5BSw8z47ngGdkYG3v+m9BhDCM4gk15PculjKcSbxTbSjdvf4z7qdcpm
EbGpACeOoDcKnwl1J9m3rZ7bn7ysLRYcxhhtFWUbLfjpr8C/AoX6veayHI10g/MI
XhNfwFvearukx36TIdZDjcd84vkgnlW7yk1g5ntUKDZtcdHuIF65+Ljmg9jqLu+F
3y5A1t3arVuAf7lgPiMOjhAqM1a6Gg3p2fQy7zAng7Qj821Q4b22A8hpS57oAQe9
XtuK1VH6BGK3QOq8yR8tYUjOA6h6FeOwI0lEcP3MNO7YNpahVeGjepsDMhYKwAVV
eZphLaJws9EQH20zlzGAiA==
`protect END_PROTECTED
