`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oXrNDMZIltqzcj3cnqbPUOcws3gV6sLrxm1XHOS2i04WS0yUgFuqCUPgyQrUJQWK
yjwJ+lnMgSv+XQsyFWzoBPp4s1YZ1/cmKuBHSL/othdxgD3NYx6CGVkMR0IqupAg
Xi9kuprDpHEEJJyGqhd2MUT4MF9rrjE9BtrrJZgFTBKMlnN9GdOfoxXjaQEH4d+w
+A13ZSGzH6crndfGU/5ZaMe3ATrn4q4HeP27j+FBoDX1uBTCIEeDVQYob1TTH0Ym
UC+W/wFHusMmYNPOezo06s0IqL4V3vD7rumhVtnkUAN0R2nyUK+X69HcWTQ23o1x
EwkU6d7b1tP1ZestfDTZdL5Tbze8RgpDMibEXzZ5FTQKnk2meqJ63vqY5hpkmHLe
9ULHMAtiTF8FikQc1XnvAwF0o8OmHgqHvTUb08eQMu9MtdsX5Ko87oXYyZirjt+v
7zEn3/wKIP2IKY8evkzniZu/VlClRJVjEvCf9UUX2hWlpNDfb1zv7+E5sybSv3EG
UXj6QM0BphckkbZ+VCWeDI8VYstet2TXx3/ZisBs9fuzcLXDF9AopdkdGnlM4TXD
`protect END_PROTECTED
