library verilog;
use verilog.vl_types.all;
entity TEMAC_SINGLE is
    generic(
        EMAC_1000BASEX_ENABLE: string  := "FALSE";
        EMAC_ADDRFILTER_ENABLE: string  := "FALSE";
        EMAC_BYTEPHY    : string  := "FALSE";
        EMAC_CTRLLENCHECK_DISABLE: string  := "FALSE";
        EMAC_DCRBASEADDR: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EMAC_GTLOOPBACK : string  := "FALSE";
        EMAC_HOST_ENABLE: string  := "FALSE";
        EMAC_LINKTIMERVAL: vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EMAC_LTCHECK_DISABLE: string  := "FALSE";
        EMAC_MDIO_ENABLE: string  := "FALSE";
        EMAC_MDIO_IGNORE_PHYADZERO: string  := "FALSE";
        EMAC_PAUSEADDR  : vl_logic_vector(47 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EMAC_PHYINITAUTONEG_ENABLE: string  := "FALSE";
        EMAC_PHYISOLATE : string  := "FALSE";
        EMAC_PHYLOOPBACKMSB: string  := "FALSE";
        EMAC_PHYPOWERDOWN: string  := "FALSE";
        EMAC_PHYRESET   : string  := "FALSE";
        EMAC_RGMII_ENABLE: string  := "FALSE";
        EMAC_RX16BITCLIENT_ENABLE: string  := "FALSE";
        EMAC_RXFLOWCTRL_ENABLE: string  := "FALSE";
        EMAC_RXHALFDUPLEX: string  := "FALSE";
        EMAC_RXINBANDFCS_ENABLE: string  := "FALSE";
        EMAC_RXJUMBOFRAME_ENABLE: string  := "FALSE";
        EMAC_RXRESET    : string  := "FALSE";
        EMAC_RXVLAN_ENABLE: string  := "FALSE";
        EMAC_RX_ENABLE  : string  := "TRUE";
        EMAC_SGMII_ENABLE: string  := "FALSE";
        EMAC_SPEED_LSB  : string  := "FALSE";
        EMAC_SPEED_MSB  : string  := "FALSE";
        EMAC_TX16BITCLIENT_ENABLE: string  := "FALSE";
        EMAC_TXFLOWCTRL_ENABLE: string  := "FALSE";
        EMAC_TXHALFDUPLEX: string  := "FALSE";
        EMAC_TXIFGADJUST_ENABLE: string  := "FALSE";
        EMAC_TXINBANDFCS_ENABLE: string  := "FALSE";
        EMAC_TXJUMBOFRAME_ENABLE: string  := "FALSE";
        EMAC_TXRESET    : string  := "FALSE";
        EMAC_TXVLAN_ENABLE: string  := "FALSE";
        EMAC_TX_ENABLE  : string  := "TRUE";
        EMAC_UNICASTADDR: vl_logic_vector(47 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EMAC_UNIDIRECTION_ENABLE: string  := "FALSE";
        EMAC_USECLKEN   : string  := "FALSE";
        SIM_VERSION     : string  := "1.0"
    );
    port(
        DCRHOSTDONEIR   : out    vl_logic;
        EMACCLIENTANINTERRUPT: out    vl_logic;
        EMACCLIENTRXBADFRAME: out    vl_logic;
        EMACCLIENTRXCLIENTCLKOUT: out    vl_logic;
        EMACCLIENTRXD   : out    vl_logic_vector(15 downto 0);
        EMACCLIENTRXDVLD: out    vl_logic;
        EMACCLIENTRXDVLDMSW: out    vl_logic;
        EMACCLIENTRXFRAMEDROP: out    vl_logic;
        EMACCLIENTRXGOODFRAME: out    vl_logic;
        EMACCLIENTRXSTATS: out    vl_logic_vector(6 downto 0);
        EMACCLIENTRXSTATSBYTEVLD: out    vl_logic;
        EMACCLIENTRXSTATSVLD: out    vl_logic;
        EMACCLIENTTXACK : out    vl_logic;
        EMACCLIENTTXCLIENTCLKOUT: out    vl_logic;
        EMACCLIENTTXCOLLISION: out    vl_logic;
        EMACCLIENTTXRETRANSMIT: out    vl_logic;
        EMACCLIENTTXSTATS: out    vl_logic;
        EMACCLIENTTXSTATSBYTEVLD: out    vl_logic;
        EMACCLIENTTXSTATSVLD: out    vl_logic;
        EMACDCRACK      : out    vl_logic;
        EMACDCRDBUS     : out    vl_logic_vector(0 to 31);
        EMACPHYENCOMMAALIGN: out    vl_logic;
        EMACPHYLOOPBACKMSB: out    vl_logic;
        EMACPHYMCLKOUT  : out    vl_logic;
        EMACPHYMDOUT    : out    vl_logic;
        EMACPHYMDTRI    : out    vl_logic;
        EMACPHYMGTRXRESET: out    vl_logic;
        EMACPHYMGTTXRESET: out    vl_logic;
        EMACPHYPOWERDOWN: out    vl_logic;
        EMACPHYSYNCACQSTATUS: out    vl_logic;
        EMACPHYTXCHARDISPMODE: out    vl_logic;
        EMACPHYTXCHARDISPVAL: out    vl_logic;
        EMACPHYTXCHARISK: out    vl_logic;
        EMACPHYTXCLK    : out    vl_logic;
        EMACPHYTXD      : out    vl_logic_vector(7 downto 0);
        EMACPHYTXEN     : out    vl_logic;
        EMACPHYTXER     : out    vl_logic;
        EMACPHYTXGMIIMIICLKOUT: out    vl_logic;
        EMACSPEEDIS10100: out    vl_logic;
        HOSTMIIMRDY     : out    vl_logic;
        HOSTRDDATA      : out    vl_logic_vector(31 downto 0);
        CLIENTEMACDCMLOCKED: in     vl_logic;
        CLIENTEMACPAUSEREQ: in     vl_logic;
        CLIENTEMACPAUSEVAL: in     vl_logic_vector(15 downto 0);
        CLIENTEMACRXCLIENTCLKIN: in     vl_logic;
        CLIENTEMACTXCLIENTCLKIN: in     vl_logic;
        CLIENTEMACTXD   : in     vl_logic_vector(15 downto 0);
        CLIENTEMACTXDVLD: in     vl_logic;
        CLIENTEMACTXDVLDMSW: in     vl_logic;
        CLIENTEMACTXFIRSTBYTE: in     vl_logic;
        CLIENTEMACTXIFGDELAY: in     vl_logic_vector(7 downto 0);
        CLIENTEMACTXUNDERRUN: in     vl_logic;
        DCREMACABUS     : in     vl_logic_vector(0 to 9);
        DCREMACCLK      : in     vl_logic;
        DCREMACDBUS     : in     vl_logic_vector(0 to 31);
        DCREMACENABLE   : in     vl_logic;
        DCREMACREAD     : in     vl_logic;
        DCREMACWRITE    : in     vl_logic;
        HOSTADDR        : in     vl_logic_vector(9 downto 0);
        HOSTCLK         : in     vl_logic;
        HOSTMIIMSEL     : in     vl_logic;
        HOSTOPCODE      : in     vl_logic_vector(1 downto 0);
        HOSTREQ         : in     vl_logic;
        HOSTWRDATA      : in     vl_logic_vector(31 downto 0);
        PHYEMACCOL      : in     vl_logic;
        PHYEMACCRS      : in     vl_logic;
        PHYEMACGTXCLK   : in     vl_logic;
        PHYEMACMCLKIN   : in     vl_logic;
        PHYEMACMDIN     : in     vl_logic;
        PHYEMACMIITXCLK : in     vl_logic;
        PHYEMACPHYAD    : in     vl_logic_vector(4 downto 0);
        PHYEMACRXBUFSTATUS: in     vl_logic_vector(1 downto 0);
        PHYEMACRXCHARISCOMMA: in     vl_logic;
        PHYEMACRXCHARISK: in     vl_logic;
        PHYEMACRXCLK    : in     vl_logic;
        PHYEMACRXCLKCORCNT: in     vl_logic_vector(2 downto 0);
        PHYEMACRXD      : in     vl_logic_vector(7 downto 0);
        PHYEMACRXDISPERR: in     vl_logic;
        PHYEMACRXDV     : in     vl_logic;
        PHYEMACRXER     : in     vl_logic;
        PHYEMACRXNOTINTABLE: in     vl_logic;
        PHYEMACRXRUNDISP: in     vl_logic;
        PHYEMACSIGNALDET: in     vl_logic;
        PHYEMACTXBUFERR : in     vl_logic;
        PHYEMACTXGMIIMIICLKIN: in     vl_logic;
        RESET           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of EMAC_1000BASEX_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_ADDRFILTER_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_BYTEPHY : constant is 1;
    attribute mti_svvh_generic_type of EMAC_CTRLLENCHECK_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_DCRBASEADDR : constant is 2;
    attribute mti_svvh_generic_type of EMAC_GTLOOPBACK : constant is 1;
    attribute mti_svvh_generic_type of EMAC_HOST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_LINKTIMERVAL : constant is 2;
    attribute mti_svvh_generic_type of EMAC_LTCHECK_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_MDIO_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_MDIO_IGNORE_PHYADZERO : constant is 1;
    attribute mti_svvh_generic_type of EMAC_PAUSEADDR : constant is 2;
    attribute mti_svvh_generic_type of EMAC_PHYINITAUTONEG_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_PHYISOLATE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_PHYLOOPBACKMSB : constant is 1;
    attribute mti_svvh_generic_type of EMAC_PHYPOWERDOWN : constant is 1;
    attribute mti_svvh_generic_type of EMAC_PHYRESET : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RGMII_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RX16BITCLIENT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RXFLOWCTRL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RXHALFDUPLEX : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RXINBANDFCS_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RXJUMBOFRAME_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RXRESET : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RXVLAN_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_RX_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_SGMII_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_SPEED_LSB : constant is 1;
    attribute mti_svvh_generic_type of EMAC_SPEED_MSB : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TX16BITCLIENT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TXFLOWCTRL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TXHALFDUPLEX : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TXIFGADJUST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TXINBANDFCS_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TXJUMBOFRAME_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TXRESET : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TXVLAN_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_TX_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_UNICASTADDR : constant is 2;
    attribute mti_svvh_generic_type of EMAC_UNIDIRECTION_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of EMAC_USECLKEN : constant is 1;
    attribute mti_svvh_generic_type of SIM_VERSION : constant is 1;
end TEMAC_SINGLE;
