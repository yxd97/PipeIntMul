`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2pr+J6yHJf9Q22yf/LFMHA27H1zktak8PWXDludumqVc7DykxFfIEQ5C7WJdUrS1
EGiIltZPUgKNo0VpRJXucWZfBaMEmkM0SgUbG3lFvmbw05IUPomkq9HfppXq7x8j
2Se+ofdqr9mFm90d4EwS6aAUFVdp8wu3M8cIi9hJvPgz1nb4qJgsgrFfHBQFNLqA
8X2vJ6mnAMTUI1CjVc4+rx256NvvrS/KiDGcL2bXjwQ0HgBJw7WoLvdUg4tbMKCJ
Z9qmYx7QgwqizGVVHfYoZKRmGtzPXUEMwhNZRDUZuUp+vQKoRYKGoG82jfEuGRu3
brqzipW5TCLqzIHa3aRbT60r+26zSEL+ha9UTOdy+Tu4DBZTcu1RE/NEfaxJddBX
kvYitmdwwimedb3dKn6T4+WmwLud+tYcaCTOdhBXJDGbr/BjgKo3KwcqA9+UgUCu
zTxqyuBseFiqVXQIgvLPRcG85oyOrGdFKzAaO7bAVTSnv6KafL5HY+i9VuUaMDgj
kGAKjk+yJiuzKax/dlDGarfrYTtAdP4cO/VCoVXd6vedUo4CvYosO1h0K3NH0sbT
4b+CJcjQbnDXk+BxshmEoWS0LfnXB2WT2AHwiXz4sFvl7Je10nSAqR13dIKQPUKx
J8mgfXoov1TH2I5oJNw3BRFw7Z3Mq2x4dCzbEbRrsu/3yjAp34u/7gPheu7TENSn
nYbjxmMicB19tq7sj7zLOb2gYzD1vpPTw4stUyr7ErsuPVLADtGOYZvxdsZcv+Qj
6TWLxil7fbv5SZyQ+5EnIwnPB2RKDyziRsc9DwqHkef5PMYK+1NTIYVv9hWS1ijY
XApEwW6ZttgIfKy0fMx0+V4f6+wcQOEUj78ZoLc8FF4r+KwZVikE46D4ggLN3kza
5TQEQ6fhEKEVOrM6z7QAgNh+te/xhkB7R0vD13sUOfbzP7bkcVOuWjxYOj5Zxi6X
CP12C4Ks8ng0N3aWdXhAAtIehbZbii4tD7QRK0PPmjT5g/qennb6p+8EnGg3d39Q
7HPUhxYWm01IHaaEBTWflRSvc3LQqfabb57sM+fMK+vKqRmKjYECb455ODlED3Up
8KNbhGR6Am10FD+ywtZKvjBPgHp0TiCsGjO2k6IZ9bNS8xptDuzP2urz3MusDK68
O1daP2MtyVAOBavZTuFAewFpviAcIEvgjLIMS1VXThKSKbiLUxONxzQ8KD06cQKZ
jdoXIV3yVasHwpxrKfLROkat65hqf3NUeJ2Dli7qWiQgQex8DuWunuK6Nb+TI1ZU
U8MPg2uVU8NtJj2eEPTNVXLGeZzmp5DeqlrX8SCsxSpI/lKmzwvSpBbVtRvHJscm
qW16A0jiJg5eDBslscEfx5oqOL+nHYhZnVtd5aGIZPYyhqbEW25ChCeaYtfnion/
3gMd07wI5k+++hYy78PBFgn0yu/gMMboD/Hywcgf2u9B1VmljwWcKRkIL6ZU/n+4
3k+9usiHfHBR/9WJd/rugoqo0IFuqMJDeg1XZEpA3Pgna/HBDpvaKACJAIiAvDJt
1X55J/Oh8KlcqIiKnocx6PxU1MjC6h9ZeBBNUvZ43gnw2Zsx9BvUVZkR7Xzq2ZK1
`protect END_PROTECTED
