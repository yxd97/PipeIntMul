`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YO0avegFW+YHEur5ixhhQVKCPAY6Dckd870C44w6dOMgsJJm1qCWsqvZrdoTCMdW
f3NM9ecOmeRqxKFnT+Sv1mfkMRFkbN5CSjG62Wn/GRN9jPBmTPxFslxNtDL6rLqh
/VqNU16zJZyzRbM4kFwyI+e+BFRoetgOgUXnUY/C86Rl6Z/eh/lFgxupFPyjyXph
rGEG5JZO9mR5I+0AoO5ESHVEaqs2VP5+/9KXVPx3qz0Pr7E2B/wAROywVKlRxbHw
wVkRXL4ofiRb53QeOWKVP/gqPURGzkqGEg+mbRqyZOlPQqx6mxhmtnTlU2aj9Q7F
foQ0qJJIo0NIGet3kFy/vTO0/I5tbZ+W26W3uiB7crbJ7qFwKoar3c9tVQb08HS3
zHVqLFZk107CcFBjgkDa2Q==
`protect END_PROTECTED
