`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4H4IS+BmVvvo6na006gCv+P9WZEUuLOJag7WCfM9aiw2DqpEgogGv+ppm8nFQlS
3tGNqQPXkoVBdpEjPRFvMibGrrLCbbu7b1Xa0PolQqftX/tAr27NH2ScTe26+xA7
LYFKvuU/jNLj4egl78kfZQ8zunlfycSbNU48lyPgQ6whjhAoeUq9QEwGwPiOLq2+
CyJ3GQtgW+TEa6ZxEuvK/LiKL9rFtzOWrdxnMUetma7M+hvPlycyVsg2Y9uBi/CP
6MXvAJEWHlh+XCcRtv6dvP/Y1fcJzC11BYhInN3VkirO9JBWHNHhQKi1R6owgo0U
x7wdsVlwbd5TYTNZks3O97nzr31p/2eTq2q3RrSbz/ObKoNmaBIb2AcscQ6+l4au
6FQOzWPOg2iHu+DjScQQRDZkzjgnShRTGbAo3yfPjGWFVw1gsWUzU6Sfe9fDmW4b
wvUm466HHRQ0qFSNMBjVTdPhT8zLp7oI/hF2Px78uHBw6qha4LJODGfIRP0eOXtf
u9JbvIPd0unQ9RI5/b5WFAB0kb1F+noWSIppiU2tHp0wtEFDE9TUgxMwv2JroceO
cOrV2BLjtdsv2yybhchxkrCYsETOR5mkDpPMNjbHUj2+k0dnoxeR1j+se7x16Kqx
Ss6I+at45DV+ZiOVRB/U4MNLPtuDki1YcY83Iasg42HRurY3gYZ6U2832fhy1nDX
gt+JN7UphtJFFkbsX4V5g5xTFCgtTE78UhoNpcDwrz0LkOLFu1jU5jNLQ4tcvx7r
7wd54LybYTL3v1P2p1hHWQ==
`protect END_PROTECTED
