`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67fdru54hS4ra8V0R6v+VKZqJeg0NiCaSxVy7I52hL3io0PjX5cDauJ/Wn1bKndl
4cE6J0u62SZGudnn6UHWt8ACT/n/WgdT/sdQbkxx7SzicBAcCCN1x2sFZjcdfZ+N
e/useFTemDJEWIHTsRVoBKJ9MDd4RiKEXiugv5t5kyod88Zhs2989E3UA5k/KlzJ
43m+ZC8UJA3Tk8ryGPQYs7dic70JRuPNRrPerWZ0fj3rxiXVsYrl55rWxo7Soedy
ZR+7y+DB8agqmZ1hpbhFt95FUNf2L1PDdOMPF72nFf7GL4SeY8rjFA4V8cOrZ1pp
cMo+1sqMFHMQywLsQLrUohPktA8EvHFualj8zxe+xQz/U/I6QK77ovJ7OxqNr3Dj
4Z+BTYbYA6G6YvkyWcM29QSCbt92/RYZstSfRMFAKEbnUci6/HywSUwEEJXy2Bbj
b6HMJTuF8LVI8U0deUfuV8nmk1NFdBc93ZQFDq777KW8tYDnkhqwTTthluU/0OtA
xnT0Rnx/bI5DXrr0PSWilw==
`protect END_PROTECTED
