`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epIkU8LGfcpl6L0PINPrCQO06MafVQny+Tfk0cJOQeGQqvAse2/z79h1NE/reuSM
cDPPgkIrslczjfcjt3tQ3FVWxAfBqnoRIunWXXM8ulrevAB7GZeZHF5euIskt4Ez
vMS11FXdTPi/Xv5K7xpvs3P7utwiwpcO2c58FM8ej0pN1wfH66X8hRu5Pk01NZFM
VabKffScxHO36I4Mx+oHEZ3TBYM4p0w6vp2ahGchzCyLulHmC0VPXr95OhzB8Jjb
1YKIzwRmE9Q2p8RJRMwdq6NkK9f6USAuPMCAfkylyjbTxD8hh3KxLtmBnm8svVRM
n+sZJJYvTwqMG7nXCuIJxuD1qotafezJztVpMHx9abtM8OxWRDPv7Vrqh7KbRUCn
JcHOfAiSh5yatdmONhSEYBfFsb6yzJ3zpo5Gj64BfEpGQ8Zj/4iI4Vd8QwoQ4VTW
0jooZpynAAn4e9ldynjRCawhww2E/LiWYEdO2/SUiNVFCyQgDU9tDhfaUfTpbQWI
3Tteg8Cs5zG89AgqM7ohNRAlabjBX1SxuDNucc+cvLAU+/wWrnxvDEnEIb5qysCG
sYh4/MlLB+0iVZkdUPjRAgxKhoI8Rme3JjJfUJ5ztZ2JUzAUh2emNOsf0/jbW/of
`protect END_PROTECTED
