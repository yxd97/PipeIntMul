`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B6pAnq+bw7o3yL2N1IPrj0u9usqv97hRiOmsw3zHlf/UfkJ8FngX/5cxsuDq3AQM
ww6BcBEhjhxWC+d8/p3cyizHRtg5p+pTiMZecDukKZ2qhWZpkP85IlVTK5PxSF9B
bsNAER2CC56fl1S3bxOikW0016OTR4mrnJ+CRdmLKLVv29t+0eet4g+bJoAXfzOQ
KIyGCRcI67yDKppI3dXw9KKQ95dFZgy0DByRxekP9rA0YLJswF8Zy6fn0TlGCPG2
92AAJXzpAoJJ5DF906ik+idbg+A9cLAtvbld0ICtPkgdumLzEIH+FzkObPm/tW+Y
ZdImHNtdZywMNa2TFprwrg==
`protect END_PROTECTED
