`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONkSNVZ7Okph+5LRVx3UVoFmfPYDgO7/SQJfozA6e011q+hUv3wDhsUQenVoDNL7
LGn1QMLtPeL1VOMmuQbZhR0iVSXzGSvc/sajZVPO6JKGAbZ64CW7KQr/4urVgZNn
6+5+P/aQ5+uldVXChnMiX59GziSrwBopTQ++9m5GzuRJ0TSlxBVWXQk+rWH8dLGW
jrSftG8SsIya6ZUUOyZuteX74eVM8UF/Ziz3G1TWYzDc8pBQZ7dMvHbpr5pnu2X9
q6IzhvitxPPlCpzgEZQAA3XdqTvP+1pkzDGs/zNhplqEArkKDMd2KhAU30Kpp9MG
RAdXAgvaApXRbk1kAd88YgOol8djyJbXlkk/dV4BV4eAiFTtx9uWwCKB83qcfcPR
CwNZr2zy/oqqexat5B7KFQ==
`protect END_PROTECTED
