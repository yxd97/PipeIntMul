`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
icit1vHOJ9Sw/qfynmkwdxJsnGT2RJN6hzLJX1D+zbvZOHFY2GibohBuQw9/7SnI
ZWJPrQrFfCKbDBr0wzrCcNq6n5d4QrifIPipNfUxSA8aySDqjZ3aeDI0C/YKs5UN
5L7ud1Ru2pOmp2fMTDerWQ2iH1VyioqwzNKYz3A+w4dPS640dVKo8vzPGwcE8200
4jTAWex+PoqWpBkpre/Li6Fz6G+8Sex3KlmXYVyw+fXxmoZtSrpeyi2R3g8vcSnT
qOzWPNmRojcd/oo9RwI5DUxD5ojE6F4gRKCTrd0v564PfT8HQ/h87+mujoyVz7o2
flOZQQiiUUwKRZ/+zBxRChdUrdX+SXxOU9xnfwod9gRHULVG/gcnEwIA1g/s53TW
L0TK3O3TduPQ7HGirBOLv4Pa3I7DDcgxG1etJRKDcMRAAzp0jHL7SKFUWo6wXeFM
qBuQlyBbTI5Uc9limSWVPxytJx74ZTF4YH23317kaLctYis41huq/6nsz/AG4DwC
Bq0Yrv7bpO6p3LLwer1uFOrnZzeP+YoYWDM8l2majyO4xiV6pgapjR9fS4rchYA1
+x+8xmvIlJU+k6ha8wcdjFl2Ib5wiMN654ByGOq2U7pAM+lhvCDkHA6tf7xrnuKC
DEzcEeMiJLVfOY0sMB7rYufwNsfDGm/q6YpQdS6+BfD0m2qlsxos7oI2eRlQbccV
xBnFYADDTeYT5BbTVp/DYW/XOMCzXzPnvV9lCbZBPvzPIDEUFo6D5tPVRx9lSRUF
mfilTlgvwxQk4IFEegnYCG2VHoSIvBP1VOWIzCLDqbb3caz5bS9akfJCli29vKtB
AiMmU8Ihb+3beT3ZgziexWw/mCqPBQUoITbCUG7BlAVnCIWy8mlHGStkVsBzCCuu
Ua3syNO0B+0q+LXNkJVIiut8RycCf4f1iq2xMgzrnBgudJEC5wjNHINXYDrHQH9I
j711GMrhavWUfJY9Fy1rXyZKF+DN3g40T+7ElxEKqGhk81pWaVcMB0of1fU79Jrc
/LwRIAC/NcHT5XqxsY9fOlmx1QQ/wLwLzvBB0PLfWcoDCj4EnzzxS5FhSHhdNG7D
IPg7URPUVEmCRPDwUAJeIBcLsmqipVtlzVI9erz3DxWy/6IaVendQnwnwTxV6+0v
mTa5S8OXmrfz7vjtcdVQ69A30eowzKQBikLJTFm/haUnqhtZgWGN/iW1aUXxYMpV
ylzkIGvDG9AAGOtOKxQV2gKJO3nJthaOoPqCgF/CHrxJCwHHNBdN8nRHBqsfvJ1T
UW1evDViJL9PRPTf8CP87sFlwABM3jzwq2ha8kJt9P8Xu2Dh4iCmVZXte0oTRYyI
hfqBpJVZyLLGQxygMGF3CJDmcafHbJOWWXxQ8usl8/z7gP+ez/tBDT94g8HXcO1h
yFOFUP82MDzttgCioPYgffJVm1pA0OokVFs/Qaus6emGVUe7yK6SxG6Jv3lR7Dus
JQue0vTm32OdzyA9Zzp2o0qarJ4JjtIdtY5tuP075CanZnN32FUSdy5w2N48fP0L
HTX/kX4T37xZdZ7YajuCC+M+E9iRJOnAKRcLCcAjgyG/B5MtULh+k8wF3Soz3V3t
VSQbWu6ntVwEaKiJI/Ew1kfR1KgP4r1nFhrcIy15hqJ198V45YIqMFw5K2YTkFxU
OKTfW6TWGqTD1KMDNIM3uJMHNN8RmqBpdqhJO/4YUkihQLjodCuurOlheLiAC7KO
OwomMXIxe8vgdSKCP3I0F0LE6w01DyUxQ/6us7F+x4Dnobhx0weFIFL20eVZ4REO
qW+BJQSWfhLtPLDAzju5PCmB/XWWO0wT1n9NOOIqeNmVXOvNfH/g/gaVHlq9xYp2
vtHTj2y7NmwdmbX/2fi9G/mv0SGajtvolDYF4k5riJXReQ33MzfwE9Xq5ENhw5LE
uJbqIdaaJ36i/WprWPNaFrK0q3X+zFMDEjKNkoylDQ5LDHC/Qtoud913A7veFyEi
6uDgUx8hsxvbj2wPcDIqzvQLV3T+r8q/2oKkbS/V+MjW3Lzc9AbhWGcoIC1j+698
IaDXCtsySRL6W14zGk8Id7Afm6F2B9JvQXgt/4JW9CFNgM4vAfYaKuyyJVGp6Xay
rB14RSqjcQ3xW93FVzZI0k/n4s+ZrQhfCaT+XbIHn9H2qU5ONVWfUI82QGme0y4J
vEzb2xjcm7+WDtjah/M6LtinqdGqGC55BUvpFXrTDyq/X9KP3uss9VzXmx0IvwTw
RENhvoIDEdxkuk2/pkXo6kUW2qW2fFeu+gfDSAouU7bT24vCVlnjT3deka0kvFVH
qbQrWD80hyAjBBYpERuJlOUHSqhY+YVsb+XOAoBQVGBuXmJ1IjnaTGQdLYb11oWx
CGIA85Hy6u3wL/9i/kRj2zrF7RpST1KwLd+KK9acg4xBK+JFyrtvB4FqOQgW5pHN
bsCpX6WUhoSSTPWnbkxko7C3XI9mG1O29xHPfaAHraZcqRqC8j9GWnKMGFMCkVx8
UbAsMdq9QXNW1JOX1qqGOJqWP7pW2Iqra+PNEcSTqc4aw+pxVZDIOfG0d9h60DCG
o6dWdrqT1QZdAnYKwoRcLeLVRhtK2QBu84cOkZPAiwruFRzi7Iv5DnsvOfplkIDz
8gnUP0wqEDm6PLeIKwXmYDtTHYQR3OF8S853z6t2dXwoOpI35o8Czz6r+jPG+6SE
GwxEboikdmDgMVIvMGhGZ3POkVHvAm5u67XPlt4CAxktJIzNYE0uRQaEp1KJXpNd
Aa1pNjkEc5hgGLRy5NUcG4ctCdDjNPCZNOQO/mHSi0vd0J1BIkf+jPS+FXBus15K
7XLvCsr8J+SqXB+kTmuKaZ8BkKV6njhtQTAGOvFxshmugy7ESgz8thn35Gq77OGt
iqy/EEd603dATGEDrms6eTyU6KIOMN8qP7jkTXmxtwGSQ0dxGNMlDW+xSDC8NXdz
7cBvkUVbALpbxguxP+u/hgKKISkSiPOLplt/t6oQ8u9pkj+5UfI/E+/VRsQR9pW2
rEk5NjTgJYMpOMN4d+W/ucYPpkbh9jjbslY4HAQYkDzo7Nq6sABvSUm2GblGT5S6
Yb2Xo4wBz+qiMVGwDnOm+7LCwso+KKXrSv9UlpbUQoWca2ry0ShqGDUXuZjuWEu8
0JupTa65XizcKpdZZh04edtL8XKuszecpZVl1Xtq4B97JUebhVuobLBBIsOJzlzw
PDY5qEVSiD8ofC30oqA++oFGBJB+s+pGg25kC84MIHVxUBbD83mLzY7g44MOGIPP
MFSa5I+w1E+UaCgBiE67OdfN/yuPLtxFMvf/v7ghlnMfRiaZiYA0QJShORrNxq9D
oltRE1y8S639FRMJHhtL3mAog5a8elAARuIk4P+DXci9tMUfLmRpSCQbd7dAxq4h
TnXp3Ak7u7rS8xNJFe/RN2PmrrlpxZFx+gpqD5nu5KgeTye8sXzB813CehZZznEM
gC1i7TTkmigKw2RsuxOZr1IVqzweCRQ9qd/nQbWg6XOn21IkgjPTbCc7b6H9sgB/
zotr6tcYQzJg4w3NAJBrLu0sPrQiWhUNla4LzoCt/LvynFTHtoD7FdBtpACaVxFj
+jMzpu/fDD7nSaK3HVwFwOYxg9FGJQvXUJK3rHPTKHqsTWOvhG7bMISSGIzWnZpT
4wA9A8JzEmvuXBRHPscWun32LcKLsJkEq69iJVuC16hg/6OmI5MTSDVN12OHBzbw
HoNeRAeSuPLDQcfMmGBbX5DGt/3663aRpRtTOiJwlJbK19FKmd8oLSBM7OMc7Rip
Cl53aO+JOJ78cM+1+ogBPYIeNQypDEE09GBn62NGD2pCswwK8RUR2Z9w4kH9VuhF
xm3aNEjLpS94d9W/X7S4pn/rkIADxDF3aq2QRB1EYJEWJDOSh0MJOuSGm9HeQyVy
sB7Qwyr3xvnP+pmHZzZAgoPgOnorZexnBnB1EzfNYT+HTLXnU4ZL+DxNPRkE2uo+
hrqYZj3vKfeieXr9YoKeTmGmT7tePQTbH3L3qYLA9zfyr1GJLuGeG9av+PgqGpDG
p8JzVs+5INbAxZ81WI07PsZwcdxtXdLTXQ3PkFKwmUrloE4C3GIoCgAH5+dIGkHe
5S2vIjx6je3t0mYCL53xCmNBsQ5xXNgzEDfKckyLVZyRXJo5Ri+/9oRPLSOZr1OF
NnLNikx98DUbbonbgJFRjdZCGkm4TuP0cNyM6CnpDS/XEVXoh4zh7a02JPZmDQiD
xL6TtAVHk15PyBxZQ0kbIptGZ5ceGtNi16gaOxBavfG54PFKlEcQJgUe4L7Gluvt
E/wnPWDBloKxi7oX3+SlS/uHnTuyO8bgTKa3iY9vBlr5zX71T2KYbviLuewgEzKw
xRK88u47x2oyqETCu++Yd/wOCsbz6TYk3RI95Fvscn3tjlUWgEG/26EP/QDzeZLB
u3+PbTesAfVcIPLr1MhYVZRxlwWIXbWaZTb8GpMa5FUSiQkojwPKFHghFuNpsaUU
Uf5Rk22fhIblLuuVQ4xHqe5KLzcT1CFl1EbzYacPLIOFScwvcy76qFWQYmfH1RmT
x7Pudw1yGG65u98ew5eMG8irHHvzg8kzAbqMSy2Bkd00wzSN3mwSfgMZVXZ3KW1G
WUJwe6Pr/0fuu5Wj/6qk9ZUap+SyCnExlyOK75E6OJOF6lJZ+5xbLoduVAP+iSj2
Yr7vmUe3LK7xIqu/nnJ5iJ4Pa9gVjAXWedrhPTLt9xOJMr5+XtT5SwIIu8bIIfQN
zFr0KfmgvozUTxhk05beRmJYeY/YV9DT/tFbV2R5EvmImPG9IoLehoFKhSBvQcGJ
YOxjrNOiRVEiFASJplfpmBia3LYS4H2MLOytfGpTOjntllPuf0y+BpohCJzaEBWp
rl2E6iuh+E0FiPFYFSAd5nHHhXaFIk6Dmmsh5avyTRMBSI4PoSS9YMSaTg17kW7B
Kex9SdfaCy52E6I5c5IZ+1tB8YqJbzrDWwvEHBbBcijW1X0U+6+NcaWRVNyylCnS
pVSHmjYf+oDbpjGrQrFbpQLxkoxb8dc9Z7F4e0dS2yERmBHOlgTpsVCcKqqLn5IP
vqTv6avxyXICWnJZHVtuoGKlYDmxSZSPsyzAGRlUP9YOpdzjlbZ9jZKkrGwsxSm0
/J+awI8XbpvUqaM+GDJF+8PBDSPS+qTojwiCuzFUTILYipD0Z38Tsf1nsOziZxuS
kmr5lpWCRj2GauB6YXtPryeOj9saEXtgrYw5t+dZzpKSosWWRA8biNOePU9x6TvK
ENJVk1bXKrjpvKPTks8QSn1MJ0bwYMjHCLl7xAsZtirRKQxxE0UbvyxZUpqNBLdJ
+s6Zr/6/tOi+Xt+MQNAb1D3XhTnm0BNXvuFldZZEAtoWXHyf9IJHlrD/oxXreAqd
Ef3YWfiZPWGd8v+B3Jd6GgiOAzsKyNac8EyVgbjTP7ee5sydcJx3b8Uc6deFci4q
9UU1X+aiZc8SMo9qhXrElbdsPLr94C0REyL+vmT621GQaQfE9seSYXuWY85sk7P+
XR4P/guSzd+ZDl8mrwXj2Ao4dW/qqtL59upyHQHmagN6QGDukL79FRMpnjyMMgZY
VKIUtqg2CbVCslBdak7fnIaKGyhVUHeDw63/a/+JnPns5bDDAUkrvEsq0Wcgma6G
3uEu/WMbowEUDuHL0x6wDlKOIfhUxo/aWPaUO/oaoYpEBCsPUNpArPMqmlDZAD3z
9Sze/ioJy6sooNVfpR7ISmaoqNef6M7ALuyBhWq5MDs9LgwBxO810HY/4mmtTKeO
3I6w/xz9sWg7OBtckqyDgjjLbqu/MwIBxFZE4WV/uulzAQMOsb/MGomadw8VAb49
ETwZdcoMpdh6jp376GnYP99BlEKNrGshBvsYEc/gJi6YUxXeLp/Bozz307KSfV6U
eK685jEdTqAwL4IRc/QFY7ktk8FsgmBX8uuyx50PM9d1p2SoizqnItEq0ULj0r2t
rYhCfh9OY+nnbURf0hv+ZNE/EZCLFKuaae3h0a5LXUh+xWvuhJm/Mne1An0gtYAN
2wJa/hlYTr/Wnjjy2yxGuawi1iuo2KG+6DOHUi7S6t+sJLVtazMszipyN0aQeZHY
DIvvAZT/09Y7RqkGrGgavTJaNd/SYD/mWhcpN0ldK6fzT+E+ZfYYRahitS0FnDkm
g+0DTTihDAHFNAeSfjkIDY+FdRqY/QUnqC7JIL+THtRUmvDQDchz3IjKi3TAqbC7
ocLRcgDOGz8MHdX9HG3KmIvj5OE573ODlzo/x2RhuSah0eZyya/vIaSUizZ/qcNb
AA+i5670frZqoMxm56XJKxHdRWVmIHs4pyzts42It+5B3G0AQtqwK5iN34+poSN2
afF5CG9TH3yO2mw2fHvqfu0IMtKfsKaVCxBsjqHYgPw981xwCo4wbNcEoe3/gkxh
3sUlvSEUY0h39ffqQcS6R/AqcpZxBE7Mu2pMyOekkFpchlTeCXLXkwunmnk05N+c
/UzOSWn5iKDaSetCnYm9HBQ+PUGH4lDR20pWaMZRsSMUn4WyV+juKGoC2IxQalN6
q8rvzFOo9w33ftYpfockM6HzR3fV7sMIluYzs+OTf6bcHIUzdtbmH8ynTiCqNSek
DerOHOWVS1uanQMfAQ7DfEo30pfrH7yuYfuVmRxGlQyOo1oOqHPNC2NYSzPHvkt5
DrF8mTpfvJaX6NsIp8PI5l2jkMJTqoBY+VwDt5/tJYsftD9H7W0B0n26/259OcAa
79to2/e9r/Qr6tLgYw+fCVpqdDzNZMiogfBq8JulScjB7o3r2X+WNV9DSRNPjg6E
Jn9jLJtXta1gzl15+xd7s613RRAblVWq8u36UiWR/rOfuuNIbwa5+zSI3Xk76bY3
qNKpFOzclBOKohci5wrVjOUlt1feadv4uqU7fpV9KJeZ7MLS+wuHv7KZwsvClsaQ
kRJFtWcvgX4rkzlm6+UmN4qtsvhDtmicuXWCpjsEvrCu/bWHLJQkoNe+PGQlgmea
SjSueZIO3Ml1Ae9L1BVwnGqJfz77bw/glRHh3/IpjI3hK6AZ8xRS/ETM8HPZA/jk
6gvMsBHtxnR4QS2lMXq950L+76JZlcRd2n8d5q5iog2Btf1vsnxOeXPWcYRM1FgT
/36qPkfgnIiaCdZeqiykKvsjvYBpmHTaWTC4dACMJc1y+pOJZsdUWZ4/NCbfPIqQ
B6DeV+3/fw+K6lOHQyeo0+BdY8IRboPJrSziB10/u6O/99tOBNrzqhnavl6T/u0j
hm/PU/94a0mDtc3P8NygPuxIhXngXuppArdEJwiHYpuxbiN0wQK7ljncjmibM0en
FvzkfI1i3NvKeSZ39Wfs0OGKMGXngC9Zkz8emIE0N0DVu85rKdBWklBTRQu5M9xs
vRP2f3GT/K8/WecmW7KTUoowLsOIRytvmCwVIca7vBPSFL1IJg5BSsnIBY4+Dvrx
6svptBFzlKQJ+n3r5KuGdIlN4Q6YYgapvIeBmMrfr1ei0ThcRmOhdC2ddjjpvyTD
Ma9FMFZf75fXGvlyh8RVbMrUnR+Yl1XhEswKWNl97qLTWrNbge9Ll8O8H7UfjPGS
k/LVb4Ev/xn/dRfwZc3sYeH5AWnSCintIpguPsIKfiAChfG3FrLBvT272VK6zUV6
q8OgtbJ6mM1B/I87ujqtmvK9SRv24SPKBqYkNLSCD5zUDaUwlsPJQ1aPPbbXdWzv
pQpmFlw3VDVDhOrrV2kuTXMpcO97EAv3JHpb75CebcZUHa4unrcHob482sZouozY
Or1OJtQYVU50ss9onotyVwkPetvLQ0u0Dm70K8EzFlTCXlAMG6S9nefw4A8xmeSD
uR4lxLcwDHRkUBW4ZgNQyFdbmdFCbXYAbuM8a0LP6eLtjR63B2jJS37XLC4qCcAl
rfSwxPsxRv48j2CGk/znsWyOMhXLBSbrdT6tbQzGFDibZ5d2dDhU3QZctpDy1IrW
JyhZDyct/CnXkp/74HzqenS1L/APfE3JtwADGFNx/+EWlTX0hw19glkxRcgx1hjO
lh7KDR+MBfMOOhhe+0Ebv5TZIOh6MSgIYpE51ZM3WPpyeLZ2F4WXhmy296hheUMW
+WAPVFZY/Tr1TlXT1gKewGaAFJ8jZ5sHRGYd6/wJzK75sq8rxYgZ5t4LyA6xhDxa
hYbmvQY4+mv/vw8G/LSZiktS6YZDjD9fUn3ipbUoPQnXVj/nrYRkXyaHEprXr58A
5wwKmIvxOYJ2QXMp8vUN15KAM2Q0RJZkBYsBsO1N0bUSRJadBtKvJ+KkAw6pfY5r
aVqXp/3Kov/Jh+i00vlRdq27qpJMurQ8/uaBhJmw2NqxaJ77Nby+JQ/v+T8gc9nM
Hqw8XUqgToEFX8Uio7Vumnr4iN6mhEpAUlpOoqA+pEfxx6lPOZqAQSxGVcBMNQrZ
1wtusTF7siuzK9Adt3Vo6D0u9FXmZt4UwlKgX7A7Gkw5qZ2g0Hc6H7C86lc+P+2U
QlsSy6NdenLo+4tqDmpn5RuZ/qkp+E6kpy/2JmMVjmIu/1tS5nBxOWFZ+iEvjQdr
7n6uEMdLBiGFL1vnKH0fPIe/wr+i7+ohDl6Iap1vFBlt9uWYm41cZ5cQ83pmjmKC
bafDH1tAXmUWxwHzij6wjCWcS52aC5amdzeRWCprCLSixVobGyUoQ80YaieSTPIa
vVok9EOvq33426Lv5q7XtS+xoHOG8H4f9DUEIo2y+HJSHyPVlXwZMEZQV2iptfiX
VXVmB4cSis4gJFgG0IxhRnGlgXSK0SJIPJ3k6nCKZpGUvp4Us3zrPgvZg+AnoUsO
n4RgOR6stDxgtC3BkC6G61bCYw3/aiCtBY4d+gnuru00f8IMFTnwyfHCbDHZfDWI
6sV6BR/HoeK0QPpnzT5VEGCU2e17PStPgDe8R8PtR4PxQZTKBgieg7TgN79IRnPa
tunopzQhvQ19krczV/gtVfMBiFOrbPliK+dFBcZHb9oeGDyGLWhyg9R9sz7Bgmpg
apwl9pFJVSK+JNML9T3tJHew05z0UiDWdsVkSmuoaHAK2aUUWUZR8aGPkMnRWGv7
n71D6DQxVKd384gewyDSmt9B6fPjvBZNCIjfPne6Kg/xt1qqIarHy51ySKhqcx/+
55vHyHKDMFnA+s6MtDeLJrmcNYtqX1J/zJDYgdxCYsAVNL2GtouaC30F/1AZoqH8
dKbvlHmZ6PmkqdrjU2Ey6lF8Mv89wiDcYiYYJ3AmwtiuO36xF8bInoWX1xXz+ghs
Y2mMNinREnSFf1QfS+g3dpRIIWCsB/KSQcpVVafi9EoZcs8va9VwTh9BhTQV+fm7
X3t4jrXIm1g72GVcOSRLLFIxrTn/vMQhwmxJB8QrTF1WBn6OV2+TWnftvwyO1ptt
RfWFdUaPlD51bEvVCHNu4TmoFSXXplusTZftsta4GioRg2U6FjFty+P68qtbbc+y
n+UaBlm7ldRTMpfrjmdAg1/vvfCcv9VJONIHcEVGhZyQq/QQBa9ek+KcUVTgzJHZ
99ccOtxaqMtQh7V+QZJAtIjcC94DzEOuLbCyQFCVtLQcWmT6yRNmsd+69+bY0vgI
o0TiH5KWgwBStVwG3+yVrIRI4AQJx5bPsCU4w7pa+qsYff3BCvRxsP+AR0Bp9J2Q
PCAlMzx79WPdzysLwgiaUrNjflDSgzC8qIoS3kPDUbDvU5R1zsn4ua+tou7VpjH9
ua4UXJ7k/+VY8bGbkG38al27dCaGVNRCU45wc4DYm/V3djZm5k/JL0m9m1tJudIe
XATX7d1mX1L7MXYw+Ff+9gY1K06K7ZGRSgHi+029rmbS6fMrrP1665TEg8poPOWb
hGZR2mIlMfCysMPZBVKPLkxUT3cZTolZ/8/3XR5JbJoOVnYa1RO5/ze6YTqYVeZY
3xtnwp41nbthR1fiy2LqEI56dkhltNxfwelOnUHPPT1024Kj1GduE7oYSV3LQ7i6
0Mw1dRPmBIxgMT0fcjb8tgkQ0Lxf966uMxxUMg4vZZ0CJmHfc14esFyij8/guOrp
qhgYRo7Gn9N2bpBlSUqcH6sq0vON4ti8FBD6GtvPsoZjlj5NqRfr8W2ITNUdP5o2
GrMjU83Ph4iMuWUMc6wRkiwEQHOJEVPfciF3uDKf+oLAJqiThcSx7K/S7f+K1Ynp
rr6x7X10CIucnopxy7xt20M/+ZezkYRULLiwHJrEsWA1v0FtD7DIKdQI9eX9tl02
Fi4QSUr5LFHy0Z6H6tKt6AtJSeEmY2Zht7qWIZGki9OdAr7mL51c+rgzlF1Zpo8/
cfq8Yum1T4t4+wrHjaq/QGgXTJPlLnUVPqqIDWa+qLPkelLuO20vHpbRHHyH+UZA
XjridjKrS4EGJyswDexKdDxSZ14M6R2cbo5Ad/PVB1Loc9XLElfTZ6dOjFY5oSg6
pzEPR+MSwVWhBCzf4yySJCVIY6+ergMXwKxuQz8LG8KI5qqg9XAMnwdJo4kIQ6md
PS6asr8ZFc0umKd8QET0AmpEHLdLY+RzY27FO85GIJ2Ew31HTY4anQ4HTRNpVE3z
7pn8vv/gSKVya+L3W9acPeXIOQy9ZkgujLmvVL1gSyKpK9lijmefj2g1I1SuzJHh
OI2en/gHxVlTFJJRSqQeB/CYBzQjq9dc/jW8ubPqYt0RmQtJk0qsefEbPjZWUaKO
wrJC6/kVLpq9XKZYI+QdW55PiZnrjIKaineKn/FuGkA6FJuumNo52W/bTpZyD/bM
+S1Cx8TDjuVOqQPBXQ+NJ9M17E0cBvnz+0gajlTBhiRJN2M9jHXjOf8iFVYnMvQN
nHLf+xabJlKY02vY7dP3UqPUdxgwZtDzud8UJn63ywnOdbHCi1mdX7a9CpDT5WzF
ym1wa4tRNwegal6sWhxFw3XIEH5iHgQ3vPUqgKYE1Z6OyDMiWRfVlUMbWTe0btN+
h0zzdlOMF+mCswDgmG8B+BJo8zKnVdM7mPgHZtRaBiDt1GtWKV+Z0qSyaGtXfBLT
O3WAgGo5kkQEjwc9uGQPGoaN+9TUXrR9GYcQvi3b1nOQG0ggiPjY2l6mqz1H2FOa
q5eJcFbLK9gpckhlIccHWZUOKnl7jV2d8tjI/HBdYezky42pS6Uk7FWgsYwXJVyN
/azdnhKqTeUBlCg103uOznnPanmsoS+mT9UixeiA9uJeHFMAFCwirjucRW57p5d+
o8k2/sldxc6W2p7OD1drVhITsRb7mGHm7YIbBAQzIPSG13RdRov1VOeOWN3RFHJQ
zet1GWn/0YoaCjVePucEr+dqHr8O0jri8enekAgxG3NmXq2ebPskwtNCiD+4PYG/
uPoJb4c3jLsjBGWns+7fe3UHEr9tdQ1AuAI8CpwbExituvI1LCFmOfOckFyFh9CB
XMsLyOlzCYRxLTkdAIHgRkJzojtbduMuq9c+wIiolJlS890KFoB+OSK22UBGKnmv
/vFKDL82LMpuqODCppu4MYQbrYuwiZxcEbifPAUFgG64niA0Y9nhQQGHFdg+FN4/
m7Vk8nALkmb9KBDumCuy1ROljjvA7nQ2j7hkoB0ua2xb2Jt/zHVXffOcQQzXP/C7
h6YbVw8AlFjOnfRlXLIdTC/ZGTsWgeA8mMf+9WhR/iDt+EFLdud+ytEDVD94IIwi
pTz54K1GJXeoLojNoeop1F+17K/FVlLfILfOHVEElYQhkOs0jokkQptkGOcX5LWr
0ceLTzKliVQucCcCjN6NefEKc+eKyQ5PU3iPdVEwlGP21ZyQPkWL9eocJaur0HxF
1GyvkJOk5VKxL9jSu8quZttlXvjWnlFmLzdjDPpJ8bvvTt/+UtdKycV78mjZ27jt
KGBAwSPgClnrtRUalMtSPIc91frAXew1IWQvo1dCq1Aug3nN/1OsbAtkmbXqGfFw
vIMSTE+xPKPHi6iSMFqGXBcj3r9yAbk5cv2rwnEl+mV5fcYvO9goilMuCM6NZzMS
N+Kr88YEaWx3aGEW/0oubNlonJpCeNrxXmPlxeUGX1lMpHeRSSQ/jekHxQ2X6rDS
UNjUizbLTkoMLkZu1x9dLwnzSZl8Ffn2gB6ZKFd25FuNB10OoyQUJJMBz2IcaeA3
CBZ85b1Vo2p10YhcL/un/EjNJwYXapFUFZiU1alwPBIgZh/1OJmVwNsHbX0SHnOP
deDxlSwctS0U0x6Gzs5kpGqeHa381jhUBrnoynh3MF5kdIY3TdDpXUcFKqpPVzlP
EU8I40Cpd3qy04j4SQ6fr/evOOwJC4jgfYVdSHrU7RkuZxOfqx8/jZHsbrK6PSjh
oSCZq1xZYIlUt+KCmSi75fQwhttKaQUJSm5TJaA9e+vX0o8jiUhTE5qQ8xUbFETp
wB4oguMwck+bub2KrSHiDI7it/sTrkI1sQFCRusmqVJP1oMLmMmUQkwKJ82mwQgx
4mvn7sINNTeTb8RzBoiu9zOFoWDgyTOX8LX7A27qb7VEYhGiNBRwQYvtUpWihyCv
CPldUb8apVL05bnpODssNeLUbS7PAtnYaxUqUik6uujdQMvVGaGubJNMKGClzuJ8
KgJQZVfCRYuq5DN9qgpeqmjOyllSuXE38yLYfV2dbv4EjIItBBsYYwkz1yyjatTE
AVvV0yk12ZWcjbreVub/OaFx0LQCkz1o2akx6TMeTNKWped9TuqHmjvnHldov3Tr
CzMvy/08FhRTJUjlpZPe5CNyL9nR6LAdOmDFiZj1DdH1JwXvq0//8i+wO3f2p3aj
U6LIo8ebAWecbwtdjOl4GRZK1Wbi+kQiFP4luPoAUSrb2tn1Fe+H1vHyWXQrk+NQ
mKbZvo9uwMOGuUvEXE6UbsQZEL5smGEmSbF1Oj0El72z6zSVMnGYM4rmcqPrQHHW
A/pURioj1JjeN2BVz23UDx2tua4hV+SMXTNrdrE0W4nwiTwz2z0oUrCDoJrVjqul
A/VBGruqoq3JgJVhntG6gwKz7w3pRfSbM4OzAFWY2ysHBwG/TX4AH6LbN8FvtqoO
hJMIZelEg7Ll7WfBNdvm1dMuWjR/67x2/n37eadIYeMNS7xsZFJ8T9KdEe1YrjHE
i96inO077k+cqvuMq6HBQWAmyi7sSF9dXMmIaxLIEtQ2BOoOUfn98OJlvYAcIEX1
hGlY3xLgxT+YEdLcT+ATv7bjS9+ZzQg0MbQaQvyBRUJ2zVOmbtqju8rAoPVKEEa2
1pPo2JXyOJcQPdDJv+x6O7QqBisdGior8nEybQk9Fiiw07iVtyhyqSpWD6qPsTvC
FvurS0XFL1/d3QlA0FOcIzEs7+9QBJ19ub0w/6P/7/WZQ/Zvnzp06slQLE4xUws/
K2yaqOHEXuIOycoQcqb3EInYWsTlc8zb2DK5XviAHTVS0d2VwOBMr14jGgZEPDKn
aXN9mKfAdMCXCTskSBoQ15DDflYceClNzrJdRyyimOIwONlZvKgfpt7Yadxvbwar
C3qdHZTB3PXDC9xb5p3v8YnoVzoXAs828SxoySz5W5J2zlp1k9DnZY9SES3bCven
SFcL784WfvGfPzxJEf66sVccoDtEbsgkoYDQJ4QwLZXtyqrO/vxFA7t9WcfvvvHH
0DPE/AiSGo9R3VGSzBxjc1nG7xpZzOcInNZ5Clj7CxbYFZmG4NnpNcT236jSxfww
7/JvfwsTT2Qf3HTZYq4I8WBvlXru/2vpsiuYk50IpIuRdoDD6tQbuYXTMJlx3R5k
0Kv52DbHo75jM7VUf1c3hMRrDg+GTbBIxelitCpmpCZhapNy7IcYGfd3j+7+ylah
TKMttUlCxmuCJs5yJZjQ/L23YSm5wlaNwJz1YXW21xbaFMtHEMxijmNxS14iVfdU
rzbLp9CBKl2feaP0vvNPxIQfZXrS1hxrfrvXyzTuM9UCd5UEfM1946u5kJzTi8eX
S5nuP1vl1cQcLF3DnoSYkZXin8ACZxboigXalPsy/jMFF1yD1lv1Ih30eGvu7jc8
S3cQcFdVme/MCHTbJsOyZgSXfcSmWBmC3/mAhH4SMNnsuL9pMmp5raCkwLdwdiGc
MBz/kZmwvEDAl2+AvR+YsuFhvyxjQQBgEXtKm5TsdA+dLFX/gtm6n5oUPLPgiS2x
t+j/Vw+51A476x2SNzo0UDKMrjj69tNErdjDRUrpA40hoRc0Z3G43HU5tdRbYNf4
J1KegAW2NoRxtdQndui7GgDzSRPY+p9z2/dWPGHPBA5W39ujunf4P1mT6ik+0zIK
lzh6fR0CY+cz4gd7wK9XVjaBoqa1XjSuvsuOdoU4JBKWKBzuCswlhV/riUpVVPXO
XfnwGopch0NpiUUTMIsRcrhmQ7FtCctYy9jjhQBoqViPbqLSO4yOr0Ugra+kmpLp
R+6mh1tUtH/hHHiPUWtS2F0wbF1mpfX0CsdhW8FHQF4RM8nDPjxwhi+ZZpXhqTJR
133ROC/4LYfxFLz8wFdEZHePHbbUCfIrxgg+nK+qJhAodPuxZ3RaxZRtQ0WzrbCO
/ThlV5DzrXG30FXTNWzY3XqudHG+5g4aFz2yZDM6n+tWfdbeY2iTbKHHCL6019LY
HbN/aDgKSeOwZFOkRTsvGDJPhM9ZOh3ln5iO2buXcB1ib52yGXhcA2y+YHxSgZTG
VQ/bwJFtWksZEnq21/BsILvX0kpBtB8APYpYzufadlTsb+n/ZgGM/AZSguokJven
HRBVc+XfeyttBPUG3VTHs+uFd0SNbC3fYQZFC+bwcdADlKW4dliyz0GBCGAL61XO
fQmb/MHnKrxMyQcqhCa/vX8SW/LtQr51KpmKe15SQKHppB1gZFW/bcfgVdtrl2OR
um3lbRQWiWZk1cFRPZb2SiGJlT2eImNeDY32BvRnKN6WCGsuAl9o6eq5NqNnRPbu
S6pmkYMkfjh3C/Nq8zgu8+4hAA8ZrJgPKjEaoXzmwb53UyKOVVyr6X1p01Po9FsD
LMaB7IUD0eBT95BpJJPG+wNhZFDGL5Uk/szxzhh0C2g8ZaDZPNGGGn6bdEt8s/t+
L0kEmBsLnkUoCuPCchyXUhv/ZcZdhu4/NnRZRJmPLYQeHTg+bw4BVBUBmCwtRMxA
V3BHxTYXj5dSSFc/lv9desqBoFTiTQeh95cT3sHCc6NuAy2OU00kPXSV1XMG9R3u
cB5BMjjLbb34YUzWG7oz+swUJHM0q1R2bqrQtnxVulM69mydKUtQ3zYHB+EGPhAM
+29t9/sFq1DyhIdNoz99v+aN0D/h77/gqIPKT+kCh1mfjfUOltVxzlQE+LdxgN20
ExxIhtBxXyoG6VJx4tX+vxycmy6Oqqa4M92dqGzXMAz7mXoaMeb53k+l1I/7jqAu
Y9XVUWD6+fysd1SQgSn04k7nC0UB3cm419bPrtQavBUv2eahHI9OMGdHjqtYo6XI
QcrgMPMDGnFPo7UIDQQLd1yn9IsbDFk0JneXmGFwyhtTjgEeqzBS5WDOcexoVTx2
wCsCPK2QW63jfOYiYXeCF56u9ScvN/rnK5+V4rQj2dRoNAOdMMBp18QNdHnPEK1v
Tmz7v2pOEGLS1VrTNOzLEEXF32eKbbjyNC415vfDvSRAr5OMSAcBfNjc1iBRCRUk
bX8zVnG7Ntf32aoxwbHmCoXbLiy3+D4X8dnElB9PAlFnF0UPLL9eUe7Cw0F4nnNj
xRwGi70nQ33EBwN6EImh5hgfRc99O4yLKK08hO+qsyGQTFrb6bickQi+w8mGMJo3
yw0GI/2B01hohfHKwt1HWF/IP2MNBm345nTsuk6Yq6pcvemJiJSblmwmYXiCYnuE
8e3HVN5Y7Q47f8jF7ZgXAbOFLnA7oRBfyBLowBHuJKBlg63De4Aij4aC2IhOgsn/
E56DDN9r/p6GWhulO8NHOe/nIiKaRkxjCaqRkG9bA3klcSbdBClxem4ZyaRcfKYa
9kwgkNXIYNZLre+RVAztJ7g9OH2OP562j4NdN9F/siWo2THCErP/W3R5Qg2LKyCb
Pj+4Mq+zcfQK7PK/SS4vCJc6qWKCSN88FwVxP93zYnhK2yOZ+Onbl7+y/eSytA1y
LimK/0NHFLweEbMUE8nwlnewyiShq06pqm1gaWzTXusgEUCVbWhv0vwnQzKcqUmk
ZFEO/0p2wVNXQYIKtv1GPBSxCwiv6bo/odpudU+VKVJigIKNwDtPfpjuppASsvtB
SHRniRMPFPtw1ruZZpahOQ8y+s8Xj8GEZb4lCHBwuBMNfoPrssLokwW/WO8Gj8R2
RqY+ZdplSyC9yQ+kn2sGSePewaBThzFMimx73hQik6xr7XdhIr+eJ0fXLMlXUPcm
v/+2MiRZtDU92MKgIhrVotC2ckgAEKVT9qCl+FAsTYsH7fBJf21IflvAVdfUZPev
gfHQiyfHOnkuZVye2I5O6aeIPknPSdkRkn5V7YB3bUC+V1oJ9EFxA1+KeG1S+DVf
JkCX7kZqY3wnnd2p9j4hzsXzk2orvPoouJPBxy2sXunZRWQJG0F0guBkA/sfHkbN
WBBou6HR0XGT/oYeDbsAUQ==
`protect END_PROTECTED
