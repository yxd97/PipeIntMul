`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7gnxGXdXD6JtEPB8EhKV/cYB84QbPH3oVmXE9YtBg3Pp5oOM5Yeor0fNLYO5GZjL
kMJndNuu9oDUkyz4xaa0RdP9VL4Uj0esr+tcNcdsZ7dhtR36kt/ZN0gK2HHr1zwa
uqE/jPGvqplp1sJJUwY+sUGrYzjittZg5QEsUPfdejIm+nMbBpJy3NaMuMGOivpJ
Lrg818XuypWcXVWzhunEljxIM6thSd1rwQXBDTmm/g5UWiBqSx2tmNKQareUsdGx
Bi6+F/tyiJRtGz19EkZatt4v6F1fGvCJcPOGTPecNEl4YSI2ghMAPXkCOkGOnb6d
vCQost4bfmNwRY/FIroh7inO8IBcQGzf8JQpWovUSyyfJrFjxgqkejG0JOEgzZgx
sdBe9fKiE+ebOxVvBhSlxQ9TRaFH2Ra6rYOtyRTV8TM=
`protect END_PROTECTED
