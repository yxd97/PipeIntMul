`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6zNiKb2E9Zr/iQ8tOhgdIzKjrraNfHkNak5rtJxbeTAZy0TxDw1NdkJxofSLzNG
ykH1dN+EEol19wQzed5kfYygPBIfLxpF9FhFJm9gIfg6CvxzDiaySO/HqxFinLUN
XwMlPau+nNoFR5p46LWJHOaEZdylPusIuPHE6oYDzLVyDJMrOqqvN2pmZhGTYV3I
1s29NHQvqlXPdQQp22+QZgwK16u6Ld09WRmj8nW+sCX0gzhuczDDH05q7Vdiu9eB
H8qp4tTuwxePA+eNtAvs8YmDnemD7XM0czN986RAPqQtzlMB50PKyWyJOt3FZ4Bo
9uYRzGCBR3wrFEPiVQF3lQXzj6cyRktTtWbT20FnUQMB3QspY2Vn7BIYcDf5uNFJ
NHaJkUyvH6hAJfrvWUrw2qGvn3jg/Sk0SsOgr0l6plf3sleJq1jN9h49okYE2fKN
lzdWgx0I70sxGHqHEG6JH8rqg1uujw04bPMNp+TIPZwhTCRj69p4+WXzO8eweuO3
MnS/we0sgKVeL/9WZvtgzn/iEHE8EIAquaQn+AIQOdyM4DzEpQBAfUBGf1Wp/+um
mxHmGKo4jQ3YYADNPa+c3phefV/Ijze9x+n+MuX9qRyaKQ46UT7T42faBFEKoOze
plCSodw/5cC50VD/+ZIHBL9Sn/UurdO4ZWNsNEukL1sP87XLYfOsP+zrcD4HER5W
vq2tLubmLuPK33cXZrARa+5kBXiAriXjp7HNywtKWpNiVKnkOlTU1IKMU8RIG9gP
3lT7xinNJCr7opzbY7jufBDDyPs6RK7FmCTOFA04aV+baALwSaN/ZG1KmpIDKMhI
qio0Z0VZ4a/eDk/GIUQUaiY0OFeIzb38BWNPVGq/0EFdigiG4xoL7OmS26GOZHjw
cguz8L1lrXp61PwJU/qouHQxEWtURYdG5D0x24CSE8kpFoOkypw3F1YvEHKgStUj
vRLuWBNJIr8dPhdW+n7Do/O8wBTAY4BQQzy/MtIm0Wy8Ghkfw7B5lSW5HSlSL3+C
Fq3Nkx3Kt0cXVUHtHmYk4xavPj2eMVFb+ae2gf/ZQAKSI4u4nWW4GjmxFZgD6x79
ORZqWzvuTINyCvilDo7Euk0OJThvZuS6QSzdnlHKYixS4XuuBMMZ2qoO66AFk7FR
x/hvVtt4EBP+BfByjz0J56DbkIxKPhQwIuztJ7y5eDEkLHKa3EY/NX3JT29R1Q1m
kRGPs1BBUh07ku9oeCW2v1lC2CcJ+2TvSda5EaWModonLiGNtWigIQVshLN+mhr/
esmDg2nE7NZECo79t4SDvubVyH3GvP/1wOVouNONi94RYKLh0XqXIsWNpN+ujR6c
vJM4008zsrCLHLyDW4RicxpBXUWuVFPmCjEQwPu9qTgP/xtbVYNzraaA4eTRzvnB
zFlcNAg0/k0UlWnmr7BUkAKe0VyXimri4PxQxhLJTPYK80S4S53HokUZ7Exv+lId
benYIoamH1UKA7U5MyJ/uOer3aIRJJSBZtZQ7wZkSKqs8FsVWNjCGyuNr1WVd9OA
BO+ACXoz59bIYXQLLEpISfwx76QhsrH1gTzcVV0SrY3JM/N6qnMxRGKFmjKIcq8k
AfNQKtb9w/39QLVCTV/y9aTTThIgKoGXgDRPfowBBBQjXTXI0gyIH2La2VavSfHh
3dHWSg5B/EL6QZEsqYoofVaOJ0XYWBVZBMDmYhANf4sxcT6XAvq5/qznfDFctN00
JolEFX5794cA/l7RtDy5rA==
`protect END_PROTECTED
