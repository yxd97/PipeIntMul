`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZSXRd10UosQbBOqJNh6VPmZDXgXBaN7GHZSklyb+23AjpXRSiEN2cMgYfVqP8Qy
pQLvFrUF9B6wSAMT0hloHjVlZ3bnA7zmXXunEjKf2yAa2By32epkLGOHN3myokwM
4FnUAfY5cDlqvNUt/fVftGUB1H9Xfr2MIF8QYzw6mbaHMvMzwOaw2E5QEgbp8J/f
iXQiQsYptF/0BvkDdVXhJCrskhWeVFys+dzHymglaGjN4MlK4h9xDjSbpfroNBSb
fRw0gpNoSOehCkkvL9cL35rHHkAD7OMqK4rYs7L4xH904UDOtcA3ZlZESUg18Efc
1+qaFm9ZGixF1vKPyZJE87fXkVgEJkYHaINtPcgnjLsNossJ5Jg8D9XRXadN285R
W2okxBzpuKpmSD/IBQH+Mpsvb+VcRfFMz+NbBmQJ5dbyRKcLsWDPPYxKsvjdyj/9
mBJUMAYncHPK0s3uoP7enS1/lcCLtpqMSS4EKOx1Cc2ubWTGuGVLZLV9z9xgCTBw
C82oLjzBugfZ/9e93R0/meM1xqymek1VHH9wV1eG6/ugMsBpMn+KirentiyVxad0
vNDZJNAFIWMUrFzsG7ZbZyWTGvK+oezvD9zEbvBgcEi9WF3nwxy+obgqWl2ewtUk
ZnQJVg5UqfRdzXRSdafbm0L4XWeKuKQq+VMASa6z6yJ7F9bS+E95e1ze//W87Wy5
TVYPAAutMEeghbY6TqGZo5HSoEK5YnPG6XDs3y3ohaY4An0cHGOayEcaGoJ74iYX
VM8s133ktvDfb9kq6f880Og9IuosmePOlfq8kOED7KQCryOdwvmopAVpQIzFSIt3
3ocP8ELtfdaCGKv2lj/sfBVMTg6SBjr03g/Lld5h9uHf/DqMVo9kGFa8NzceWkoG
Lpv5Yl/jDZ65orYKUX/rHohpqf/Q3UNv8bo+hWRYuwmm9rS96v4Zjez+MLWfgt/d
cDklYetwHG9LqH3di7AcK+WG9ywKul9oJIA885UJc3CulTloIkZNmRuXs3LyTU/k
qRaAuQzIUxP8FQCCrLcIMVCVJ70ZybpYAEqK+FoWAVRNc/zE/fvKCRN5S89+RIzQ
qKj2gDA07BnHXGD26w7jBNHyUyvbLKfI7oF3O7mT73X+8t839B3tRHXoiYEJgKLP
IMz8n1NK5oCJblNu6Qf7V0AJuzrNs8IWTM/MtKjW8L3cIh32CdK1BBKxE9MbCWG3
a6YcaoCWPnfG/XP5OT7T0oXaAMuMem97wlP4gLyQkA3ubzzYKM115IV6MTovhOdm
W/BFbOf6bkt7C8O/UExgPJrDEg/b40OxmZ5WW49Ukekh9g7Lv0ivw+07iE3QiUlJ
pYfURL4oKDdscFzAUOisTeK7+X7NhTcj+pW3wEwFP+IHINgGcwNvFSTNgSAn0OKZ
Liuk3k8UASdiMcNx3fgwev5Y+TJ/6sR2joTX7kDXW95Kk48BwK00SknN7elfce6l
`protect END_PROTECTED
