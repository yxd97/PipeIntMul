`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2T3V4ZGWLMyEsCUcn8fCHpdJOB9cg3pbRSEDiWcWWmexr+xajvQuHiOjXhIB+Pu
woHoE6P0OfwcT/DB7t0CSAepw+bC7QsOqwrXr6T9HsOZ0nt4UVSpkouV1+M8AH1q
5Qos9l2+kb2cM0Jbc4VuH/aZ31vMV5KNHSF7sZm7PeyoLY35xmoW0jEc4nso8JGO
jIzhS7dcNaWZpDwwpbEM+kdles9ILqiQwp9qybRo0PMwGD++tMLjcAWk9WNz3N4K
t9xXXDdruRkJe67cC2X/SGPEq3z9lJ9ZxPhRjIUvwd1lnXNIQiTjLXZJhpAmbl4C
VT5q2oPn5/w4s4zlz8I5A8IalkNMP81SzigeKNW5WXk07uu/uNOQEc2d/Y0ag+Nf
8xo1k3jap/EkDT5RRRonyO4ktFRt5eJ/4aVwlxZLA6+FTuvUm8NWpzydZOsXpNM6
6eZmwXm0wY7AVSw4WSH48JL/cF/rW6j/oGcy4EnE4MDTlLP2tcMAvYSpC5ru9InR
utYmXf9YhaP0Ua/uVHKVbfU1SUbRJeNx19UV2MC+T1l+rQ/R/C8gbt9LRS/6Q5go
WEgUoGO6d9DcoMs8ny26V7aZLvKbHD+HAJusqZf4EywfoOVZ3oENnuQGJ7oRbvVc
jOP8MNWOVdBKM2ofLZ1jFcePWyysNm+aNbLF83Y1HHBksBqAMMs7nkmTlLQtCA7t
FkkWz7LUGWxmKW8HcK4VNgwwHuhG9PvDeCywzPmB/sgKMMBO7meu9C+ax8U/TCNV
ihwdxfUNNfkNi7wmrpEx25+Z9zGThqJquJ5951/JyYsR6bTp32+0l7MhrJkWlooG
/UDJGfJqTBVQxPLHYepBQFsU9pgLMjNEjsXmaYkS4IMO+lkVwpSFYqh4qO3a9nzn
lMsUfrhulntC5E+c0o0VoIGSF6R6Aj5y8SNrAUeIlraf7L33I46JvbK7kp1cRWss
vUTEDq3IWrK2R33C6c8hyP5K5gNrMC2xMh1fx91977/TdGTXauVtKags26iTAxdh
23iNO5Ba9EpXRQPjG7T/W2lgERNd4HXOEtBb+SZc9Tqo2+77kn26aWwYrSSJWPUA
lWsfHBc7bWzUV1FGPr9u0NYaZt84gEe72Gb7tVMwm1Llybi/wtVAjzykhIvsxu30
rCq8tCTHkQomcwyBh8Fo9DnwMwniOPArylCVduHNX+qYmpxCTtxN5QW1kEfkYJ+d
wwrU7GsJxGMPqqD0P2g7H2vd0b/XJOY7uKpZxcF1ytQ701v4yxQyFZn0GmhTkqd8
`protect END_PROTECTED
