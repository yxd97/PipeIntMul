`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FbzPv42j3gF/uz+NEmhlcGV43gJFSUEW8dp99+Mw2oig+L5BPT8pGy1YY5bdRrSO
1JhjZWzGtbIp9PsdXAumOAqHyt869qi/GuoSqEo01mv20COfhx/+FG9mX/Df4Hxs
1qdEsKVosDhm3sX9r3YLzd66wzKdF6E8HFcLwEKR1PS5b3KBVuDtKfesCLQt7nmu
MkiMgcYMPZdJe/R8awe31VkLfN2VBf1GsAFHZ/qHZNKFd1dsce9tN8DcDC/ncYTO
fEL1EYvvRuInS/lrt0UJpIpA81MnGWv4/cjOwkmGPQiofIpinw51klUMiE6MmrVp
GIgce4a07ihIoHPj0Jr5phJWj+bWGCtXcxu5AtoJsWLOeE8diULyg0fL/2R7aE+p
/xGHhHnShqjVLMVBQV5iaXotwliBN5Yx2OwWRkXrPgxtXYg3UA7fqec3sxoz7hEc
TB/Cd6LcyIyJaJTIw4Kyc9Oo050mWwU16TMt/GMfYpraYO7ss3t6KdExGm/kDAMU
/lsr/BS0VdKeFHsOfGg1XRkDmcVT/HCchPUmrawPsQqYSHaALAFh1AzghbRqc0va
/+SAd++8jqXShZzUpG33m9olGnp5iIteAX8ssZGWvqg0VP7GLtHoLBGMQzEJ7iry
IklIyJv8hJ2iMzet8l0AgV/DV3r5/adaGt7nzebKEl/hPHePWpmkrRY8uXGrrFyt
QA8fPaqv6aK+8Vrg3wmynBhX3994t+L8ZUN6gzno6P05qI9SB+JoLnZFqocPIhLI
zDrIgGFTxTxtvB5UP6xcJIC02GLD+/sZUwx0fuUMmneuMofkRIgOJmsq19OYkIU9
G+uaVXdd+xwohpAUgpJ0iXzLDIaUB4uMwVBoDMkM9Xa2lLXAdZO7UMp5kEX/nwer
f6c5t3o3rZ2o5MCtxG3p6fVq6hTlUaXeC/PL2Hsa52Q9nV0GYvWhF0PgOUGbUO82
DbcpvIKW5pzAZAE7zRq/vU2VWPpjhD0sE/zJ5uGL8duhhRxjs9TqTM+4dkUCHBa3
6LOD4PM1acu6GwMVzBGFmPkCiYellVwkddQ5lPZJg368vYOmhDbwhoFR14WKTynA
x0jOerIXZN4yMEOFBl0+JTqZOvxe8U4JsU7eljVEx0jOCqsTd2mv2uHOPuLuRFNI
yf6GhaAljCIvAnRknEfu9I9T6O4yr4uX5UQn6HMeKku386k71R15zEowj5wW2niP
V73Zc3U7S4kWoCe7vnAWu7gma4NuLCvGO2CollvNebcphRqfV3LZRY1X4NgbmYON
w4tTybmDBD3DyMCRvDXzQ/arCDRk8YDySdUJv6SrQtdtrUSdwLQoPxY36YdCIwfp
iw9L7UkpMblYVa/IqeQWUkRPLiwsFvEinc1KO3foTBmmbo6Ertxi3ztQzzmZP7VI
heuNlXJmiXLU5LUoMobILBP8HWNSnCKnqdXGGRNvoDl6WNONs0jjvcTbcJJam7Z5
ZXLPXWX7EC5akP6+GD8cVbCBoTk4vcl38q2Lsq9X+t5EFjG0Lh7n71yD0XeG44PV
a0ddPL0uNz3xhrHCjYRyK+G8jaXcXeo1MrfB8ZI7U7sserIZLdXAgaLsggzQJQth
SlCF8iah7cgBce9Xn5+SYjuC1YHqSElPvOdLH7mV4Ui8k0XzLK1Sgt5+QD4dgtkW
6ppxeOsUfuFFAZGPTFYMfrBKcQBpVTeudy1zmNSpvmM7ePkh+sT7hMRAQPYgbM43
Z26+WlJ7CoMmP1MoKfZjjV+Ri8ZK8tvD0Ab+dqd1pAHoGg+dtXSqJnXNhMTV5/Dy
jIAzRQPn1CcfLEm7lmYhBJmRyELvqDx0rNdI8unNTRo1k/3jxnkaY1K7x6m8du8g
quxdKg65mh5C0kU26RNyaTOJ9S5Mi8MtlObxBsz0KxBTcdPcJI7+OmxlnD0YFjI8
P5mzEB5hEUa9STvNNjm/Wt6cbmug2rpQMBt0NMHbOA9au3aprWsgi+OaBAUKwZVE
Bs+XqBevtYbpFZRflyICYPHIVm4z+RSw5CgOzSBXTZzF8RP4vSgmFgztqBf2Uxqy
VyrL8CyAJPl8LSV0dyo/ZxUjjWZ9dBlEFnmkuyp/38HJEYyaBhL6vMLg+DOEywIa
PyNV31jVMasRnLKpo6NgGIaN8dVuBc0CAkuAOi26o15gEVyn2QsMzFa9eyagO18n
gC0Vj34Wm6T8hclE916eOaKrBE/AOEboaEITOCZD5EOj4RjxeUztRhzmnsDvpyLt
wzVotFIXRpNr1w0j00WcYJdAwuJS7Rn8LMHfXDzIzb2t7tkqrC/jp6MNgULXE+W3
ozfcyqwbt3a59ry04UKD7UQm9QqzFwE70i7obH+RxhtCffErMqjVAxH7dpTrhCOS
txR8LPAc1Ze4syxvpK6aEJ7EptHzuJ4SsVohW1lQnfTJVIHcufhwfWJ1SrdcDJ7+
qD3jmhvhcLLr1VllGBOhWADLHUrbowRDCnN1yBrB9Mhu8p5msGgPDTL12xZwRzsZ
ZGCAYIsFv3B1dssjTVygAyK77EjPXX+k+12zYC+iJPK7wBZwaN4L6YTEYH5bd4gU
`protect END_PROTECTED
