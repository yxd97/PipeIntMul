`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6LQciaXnv1wZwfurRWU9s56p5+ceDz+XQxG52GzMGwiOE3FIzrMZ7DPvXvGrCBAO
WhrPMDB1tKPrD62PDPmldFy7cGEcOIy3R1c5XhxuxHVWVLgi08QLduBlv86m5S4L
ujhANtOcRXu9P3df9QWuVOJ+eOMFSDBEnlcTZS6hOkQru6vqGVLq83Gk+uqeQFxB
2YsdpSXICYUHViz8kpZz6EPTACcNSXi5w3R8n+9exPHCFTi7NVQEPb8JdZwYWoM6
cfGc4QwQ1vdJ3LJO9C7PmTHDBUD3JqeUXonaSVo03MkvClXCeIujetGAhjWiEWM/
5Trayy7esM5tz12318qGMixPwHSk3qR0l14lmWUrlYOdUaGv84E+6DFV6GSQfNu5
9QayBCuzyiVsD1PeWywBnlQgjeGmvNNIySlxDQeUaK8sNM2RkBUr9KuuEkJfL4Qx
zN9pCRrb7XIl+0BKiag+OFRZcrtoHAjVlPuvsgnytQKB9o3aXESjeitk8YVauDSO
j2zkC8+h/L7rjV2Oe1vTsPzrlTxZn8CoxgTOXb3qnIs87wYXpZjZhgfzc+On2VXD
CkPYIU8IVQhcYzxNibW3lpiad76UfvysaakxVpJW8XhaCn7VvUpUQawrro5lefnk
RkswEBNdy8d8MmaLNX5gKg==
`protect END_PROTECTED
