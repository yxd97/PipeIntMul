`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TuEpVdRRHipSYMeQMnZ2y/k97M/HJRwv31pbZn4xwzjTHxNVWQHQo/S/wqhy5UGe
C9ggmXau5PmAqB+zYG61cpOUXjYurwqAe9wwFTgic6vMG2TRRbsm45WNyDl6yMkK
EDx30C3ju06ccIXCbqaS4jZLaLJVl2dQo0FcOGVmVXY5DXTaf7fuFrmRq4ySQiFX
WT4OKpTiPHynUmCPLU/1LJB8qukVaH4FqWtGcPUab7CGHEs3uxB7UBTgXgCD6318
5iQPLZYbKVl+nKeEm62r5MgNoI/iNbuBFKyTa/LCHpMnMOWbrFEt8yp39E8tD114
0OJZAwL/72RVcywLAqBm7RI2zsOvCRNnx4dVyx72cWgOC7n2xvbBbcSktIBt5tzy
frue8cu0eYp7ny/U+cimdGmWkWxSzok3oxnS3/XsGg66y8iowOO8da/u8svGNXJX
BH43DM9X+Al0duDOP4GlMisCcI+m748hWawjVa9dhh9ZPSoo8jxxgRPVQLRh2RNZ
jjhi9gKP/zm+cDHQKxZdCJb5bdq8S2aLZY6z5yKBbLBYGKuI0u85mKfcLUhw1viT
q8Ss8Yqiek6WI3np5846Sp9DFBBBYbvgq1U4115Le2cI9tbkCIbQsaztCC6r8LhE
lgnKxMYBbaZtQJL01yfESoYmTdektI63TgZWdqQYjzVbKg6czNEn7i6XHHlWzRV3
JSY0vj+h3lyPy15m7MmcIbBxzfUEOgyxcTvkYrS3O+wmih6X2afz96na9QExF8nJ
yvbDHuBzm5PZAC+ZFLm5XglqaohlY/IjY12IzVCKHNmVOYjmYc5O9OctCMeYEDA6
5efEvVPXO30M461UBE7UcXrKu/mO0NjlPyd5udAZUo1QUCwSDbjQxF+FKzdZfSLX
2KPhu7l6TDvIc7CSr9TENyppyWhdJM5JSv3AW41aK6yPvIbeRLxoIcmkzqv/nIwG
oUlMqEa1FwV5sXYb40yTkirh95OehArUqmW9ln2rzerP+uXXIj3M4tTaUostzalB
W+B6XB14Ia6H9TqG78Gpmg==
`protect END_PROTECTED
