`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
reJAh7jih2xe6ezPQI/U+1+olGRvdXutOkkf5XbOfyqhvFIsu0AbyacmEOP/SRxV
J3tmpCN7HRsAJzz0eBG1tsaMORgoG0DeYnJxlHwi0WtuTxjlPuX4zxvc5dlZI+Th
+wVzJcTSjTwAaUXHdVoxeHAs3vASj8m3QfyqMTddoO2K4Zv2VvszPZjSpC/uBwUQ
BjVFXiSVU3QCU6bz7FMF6zHeCEN20kk6/Vv/+2AoIV/ERiL/LL7KHK+H/ieii2ZO
12OCFVy6S5CKT7DktZLzB3aWrDx7U8z+3CkY+cyOb+rTSZDiU4boyTgQxTQrqx6W
6yXly7Po1BbvrwNbRHCgxU6Hx+ZEbOKL4K+bAx9Wu9jbAM4mc/TTy8K6+mICPlkF
TxUoHj+yYH51YaFn0l/Ogp5a3s+dG6mjcHHNQU0O924jZFntEWsza62y+2PvwZi+
jsqptOuFdhQDNIDoEzx3UI+/0Et7CU4ZF4C61gRI4zDX0Z/rBRkpSIZ9J1HW7bFn
KMMUSDoctvzUfdv+Iv7+v3rjQa3VJnD4YMRopDt55/6y2vHTbpYk2ssrgre6Xqdh
ibu8wAkp50R6PO/FC3r1G5sOm0RVUQlzGJLLZpEOUKS1ip3Ecfq9cBOFHRUn7tXt
fYTO8oUbz8s6DO7n69ZAwa1Jo1IpGplX9ma2f/DFxJFtq9RKq5k6WtV9jxS04Szh
K86Ovd2DkYMl6umGE4aDYkkGsv87nx2arJrNWe5Li2ceI3yL9RBwhJGydfrJaOHe
bDpX4ciVak3pzL0UBomPNXXSwulYC4GzNzRNdUgQ1iq8CmF3ix23tuyapY1+CHXt
laBWYaGfx9aZDHomPdzfCzoZQ/wsYmJ4BluaR1ALBYOeK5Gur1brTwIpcHowUxc1
VUNwCqEdvOPkux+TTIOYb1DT2MhnHv0GL+fdbnUf4JJ148Zp4fIwM87xpv+sV+s3
0Qb1uw2GqYVygnXYnQxa9w==
`protect END_PROTECTED
