`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1zbseOVxirrckrbnblypJAVTjZ7TTJ7g7jMwSuXTUWsC43alA1IFkCVAB/DNZIe
SMo+L5H99jlYffzuUtwI1TBrpQwCWmDaSfHfYZdQtAx0468GyM8HgZIFaOIBr4so
54fyuHaDV1LDipKrh+1CVECIvEzRezbQMckoVBCOAladjZPum42qooZV45iAj2l3
KpAUaT3OYDCHbFVqJRvcdKZ/m0AnFAidPp1XMcxjBaRCpfcrUku7BoEfxefplIn2
fmP8L1Dr30TvhSCeb/qukuh3t8b6Sk0ciXQ0lHmwukyglEoUYDPAz1Lk6qq8JX/M
+Zii5xEum3ntJ1/p6Spj0pAgAmyVc4CZe64EauVlqL3gUyoZ5ZzLqibOiT2JJq9X
oLxyTkiXhJYyLiWXgZEssLVhSnktLn/UMJhDTTGfYWBHHdmXhkW+Ku+4jX5wcXmo
uc9b0J3elnkT1GUfwNxRgoK1ebtLMdeNOzLnFRucRO8fzQrdvjFxI1wCb8gkmdor
GpyNuDJBJ+NgjPrpv9xpkfrrtAQaWAyXbuIiRneoMQXvocQ4gjNLhniM6bUBJq35
4+q7bn5LaI7IbFQ8u75pPXgqRnzbfi/uCVCLzx5Co4Y6rXkne1EvFn1oQDJYTYNo
ijejFQuLqANGTDVNHqespkt0g74Xw2ndK1kvgV94urAYrjcAYkIKLEG/ASA5Ze9g
36Pdqg4g90xNK0Gmhr5xIE+JcmXptnG8qnAxg4n0So3MY9VWAAKYicTYwky1g8BL
EaI1oyJ6Z+9duRO50GEAYlXJ260+v66qok4RAF3p4jYtvSUfruR2NXAIRwWhuGC1
ADnQS5w9ppKQp+llMIdmIFOhIh08/pOASRIcc0B+LlzkUxIL+CK0EqhFGx8drmEo
cjOL6kqFxII6QWPXicWKjWgfOMSJwj1sA6rDvB8vpo2RjeyOmcCb0He1HdWdFl96
goGfnUiOdPBN0CPrzPdV4EuL2EwUWaRemYa2YIp02N+t5oWkLVHUr0gIZ55VfnqC
aiZcGDyOs4rpXNFK0ZTUcnTDvawbCoQN3DOMup+TMymVD5jmmCp8vVvH2LD3jji6
8jto7S/dwHpq7rpYWK47prjEwYyxqNpeGpV0d1o1cQ+3jEo/dPK2cPGUU07ywTYt
8vULyr1juBLQlp/zYKglN2fvA54f+QPhd6GY/g9uXIpkcRML13325mY4GzwHt+tk
eIIfdaccHl52xFetONERHqcl9jWrQiHY9kXeWHNVtamNnTaFULJ3rB5AjIuH7YRT
2x8v5wDa1WCnEsbk3FuM1GICfNUFKUM0e0qkqJIkdHg/ADdZpJi3syhtkGjM+p8i
o/NppfpE7UP3T0bKlMP9t0VUecfllw2+I555ibqTeHDkNhotbEfv6emjIaUISzZF
hqkvm7fyCrZGjLscqAOsuBW3pGJa0UvQxIsE8aUvdZHmFNgjkG6EtL8Lv3U6RfQE
LVMm1VHWE5kfdnBxlcqOAGSUaJwmrHlDhytqll68kjuOriIZsGZOrEaccGaKH4/0
5cUpTzalXRKLq/b4lHM00qF2n4CQZt7svVvnGnHsnSano4q7/Y5q2z4m6d0I9KyX
9v4kx13E3cnakQguJK9hrCvgMlOo7D/UZLaybi5xyBK7nzJ08lSHac+iD0+h1rKP
9PaSPJaYjHRcshfy0dVrV4v9kfTrXGPvF9uOt9A186lwcT3tnpJIM/Kf4UE4gshH
me64gS1IrzXSnKNNERN3P7L399yNR9WbLZOuMB+bj0DgK7HQlUZuJEmWu1S+r08A
OyGzbSzkUxdiI/5+0sKb6rmaZbU0zPmTTBDCFBpAiVKIh+odcNedH+DqC/i4LSOh
1xzuuv2fkJyMoohweVG43Mh6OiB/pb7658PS1ZfQhlAMb6WvJRE/SK2gFVZ6z0z+
1sP5s3SnI9ypn2XNY6w1/Pu49zGoNSSc4H4dpYa/FBRojNnAeK/x/TiUq4vev71J
ukf4F5A8GQfLcvpVnPs2bTGbO3rdgpAiPrMvXAo52ddr6y+GjlJRJO4YaaNTS13g
wVBXOFsZEL5SmUbMaFsntVl6E6ULMYS5QS0uxlh3KNJ+BcJDoe6kLEPWN3rbFAqL
v8tz7SsUjvbUE5ke0O5vO2YvLFKxeAUWmx6ejLWsxiycT8CvEW2is8fubnGHWaqI
yyUjX9MChokek/Esn5FHIAHUMLX9YB6vEJzNu24+VLKDTwZdJWyxANcag9/nKsOS
5eNY/HDJVecsBIVs9qmc/i3AiXKF2M8d0LfkJQQw2660F9jFu/NOYYCOgwar27hM
FXmUUwGufkQ79weu5MMjBDxM8H62NW5CskpHByig0jjfUHtoh68NZtLth+W3A6hV
PSn98FNkRJeQfDKiynDCz3b+indFnklEEFyL0wMxpo9rM4lXIfgF4cTR2vv0D5wc
1Jd+VfX1zfEb5EKkJPlr9yGS96y3utq/o2FUSbeCmsdEHuXr/KiHva/QIeDAXajR
WhamMW8gAX7NOhhqGtfMOxMivJezl+aWfwHFOX/DVIL1uP+R4m1oJHWEh87d0X3n
ndUVeSjVs4lkcIQ3tWp0XaQzz2IYk5WtcnnyLz32xuKU/QCt6oa98Mv/o+iQgz1Z
gYhDfVYmJh2E0k/tE9mhzn8RUm847yqZVgmatCAdgiteyi4iG5UDb0PkzaMC6LB+
D9xK0Edc6mxtXRApSDbggs2ImL7KCOUCYyAS3InORUJvf2hh0UX5f5KVfU9bmKDy
8WVpsSMjqRKvnwiD/wlP81D0cfZhSIKT/nJSAnpA4YAQtMkXDNwPg3weL9sLzWae
OHA/HEFjMoGWRGdkCBHjNBktrs6U8CzVDKfEB+oVAfRRrwsl4CHt3COhvyQcg3iH
Kd87sqpM9Ey+88rmYisiSonPB5O7oJ8yQtWR5M0jjXYjzohKcn0sUn+J5eHntIwT
EZjtgp0V0mviyF7a4nkdav7b+LqMk/2AAkMgIvmvw/RM5L9C4ZyFaQrhtXZo+qc1
`protect END_PROTECTED
