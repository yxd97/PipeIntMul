`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kYSCzIKwOxr6RjIcvSVjo3BwuGLmVP0iOuea43RzWsCn7kVO0jXVQl3I4ap0LMTI
WoWA5Cn+xkVBSkF3nnMjuVBWCLri7VIIC2m7VwpbP7UcOLxQ1QamXvx7q0/2n0/T
V1kFPjHm9IcvbI2QA+Go3bjojQL4ZJosRiN6V/eAr98++kYUHqu/eWjZ3jOH0gbP
GfhRCB1vkRvezCWN67ztjGMw+s4Fe4HdNzD2VIhgBViG0CrhlvXtUW+FqAJvubSb
2EC347Yvvejk2Pd8wLTrWlnB3PG7IPIdNN5zsSSRM/nZWWNKm8pPco7wJ4TUbuNd
nJ3cz909+UvDvjsXa0f1nQMuiixvjtGwRtsHzHyrVfX+MvLGRtiROLj2+lbRWlzF
qvflE+GbEgH6xsQvZZGreYZ60Gqdb/A+jcc7ex1hKcceHPlu/Gdkcj/sEzKr99RI
7w1ZUPxCQeNnqy/VrEmDFa5M5y7DMyUS/jIjDhMrvqVBC0zY0BLZwPABBgwXwZDf
lwUq5QDjGkpXZ+W0GadGEg==
`protect END_PROTECTED
