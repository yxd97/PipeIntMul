`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VD69lwAVczRUJ6XNFRaeaOcgF7KsenBaQ0vanYLQ36wMOXJrGGKFeNqdEHQNg4lD
kysMr407Na0p8RJhjQbJpnF5zB7tKeMZQ8eSyP53l8czvYvBGfj1LOcTd6JjRFVm
izxAlhbO9DGAV2EgI2YM9eC6d8E4QKsLAvlNgb/IovjtNMLYZiwT/ljRrAZd6hVa
m5I7LbKZ9WfjL7jgMrld+WrSS9mY1CY/lfseEpcAEUMzbttEmTUL6scdUGBtM2t0
/5kKabbsBjb6YUWBFQf+dHrHGd70uGMgE0zDZc4QpWORkfnOeibidf9yeQ5GG+9/
e8B/ZrU2A7bjGdqJAvF6/UP15X95F/aMillVX1mGJUAlBKWLx6gSbcJMcunn6tei
DO8aj+7nmIcZnjR55XysMjqjQp4zR1fAGG7yWy2wNZW7Q/EDtfxRXccL/bkpOmoy
WMU6Pr5g3px+wC+9pTf+s02jtxbObPxtCviyiG0ctaiOBO3MjkGRNUQS1gXztJ3U
j0V3hH4M4hF409FdyyhPoBY2d+j+uj4Oz8vlP/fWoc+TTVt3ILSlnDBMozVk4ruZ
DB+di4ECcEKWiMT1RF8cmG3SDPH5S1sRIvE0aF3HinDdguEbSUb9L/44hhZIUGqB
hQkfUOuuXOoDYCD6T6YKn3/mK/d53AdopOnVjMXMmqPuHda6F+SQ3CbhaiKc7Z2p
AR9YxAiQfIc5Bm34tMh1r6RRhzeLxiUE6FEj1v5iAZLsbWulFhRzS0v6GyfJAb/O
unqzs6qo0xNKOY5EIywH7OXdF1VDkYQpZh4LN3qILNtrdGeK0LhrowUBcK4sh9sY
CUHUOVeBflUE8zYhn1tC6ljUCHIJ84+mWW4fFY+JQNzRbqtbrIl/jryx8wNG0+Bc
KUWn8i0w1QfLRTZVRlHMZgdDVWiBIbzcsbzttowurjoLKYuypIfdw7NAOkSGkVtx
HbajxRiLHaQZaOPYp/B7AId/pMMcT1supFY6LdseP36rrkIDHk/XBoC0cOt74XSz
x/6inrz1ARakpHu9jkd41YPx63eEpffNmN2fbNVcxtuB5CUzg7wbK/OWjtlqWuJH
3EKfsgysNzH3j7Jn5qqhPbvM00Wgxu5+In9fz5Pc3JhiSnO/JyajSRRRygfd+7s3
j4AFQ7g8juX2n+K+bZPMtnTLoNUR5aHqUT6SKscs7YQHYdW1qqdEIfH/6BGlm+Sv
8+VpZovl6Ws68cEQjVZ5WDPq/Huw3YnC3sFNeBaLbOlmPy/3t1jqT365JHn5Pi3f
Xip5+Semjv/Vr4oKt3gnmMWZAvMXP3nu/Gq1DCzl6YfwOGux9zjmodALhMkuN1Zt
354LZXsMErGbRQ/SfogXStR7xtxf4nHSr4AGRdKubIhF0Soi5w/kF41LvoLdDNXL
6vNr+iIojSi5AHvMSrbpinRJa+Ket+D5sK6lHJp7w6C/lCsF3cBT5M/vJsT+cKjz
xFQZZ/5dGxd46/wex/+2aGvkldncfbuLsKM37R8akm9Bm/mNgl1YBjJUDgueHfkU
czkO4QtflFX680hmaeKLWCTMysrvUZitNc4u+ic3syQMjqqV7YASXloPvlr8ybgv
FHOnJGUMpH/HWuKs4156wllprvWF/nj4Mfj7SegY02kmtlQBxQiQgYJ2wi/qR21q
q9KsZblYqcbZXboGSKi2okRAq38fq5RGt/SmI0XzODA=
`protect END_PROTECTED
