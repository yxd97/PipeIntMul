`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kuq6xRbL7vEC7jd0/ikCkXcTj3RoupLl/7dmwylMCKwsKPkM1Jlcm58WsB+HaVlz
BpwqqyYpZGTySMdqyPfuc/ENdIVaLByY9vH4fTbNaQmVdSoMAatgrSR8PnWcuT9Y
CQMZeZetLg9uXAncFuIAUHetj2Q2PaEUKuNASWC6fyzHav4Ah2SBNWxjabKa2i3u
/+TJjzmBOTqofVKpC5T2NIELblHF2eTecFVWmM9d4mztaoxCmM4fHK0xNVq0xxk5
nzoCxCUhB6IeQRt3bU0GI7cysh78kP84leydjv8Pi7ypNy01HOFIhjiJQu1GQLnY
EZXCV9zyJ1oZrWZhxhApAhjq/7yFiRRudFUSVkpcIUyqB348Rc2Ps6+EdG2ItDoE
S28vLos/dJK0Y6iDFJYOsV3GtzSPA4svRiOGXPdTUgCJPsFZIu4r5Y+8Kutntzux
U50cPKyHeJj1j6Mv7PFaKaQdC64+D24leeeTgPdLp1U=
`protect END_PROTECTED
