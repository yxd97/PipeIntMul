`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DoBPFtRExs2y1x1TjYo+qyMgD6NR0Sm2oIrHPGcG+SDXAxO5OF/szv2LxRuGfG8k
t7uFng7huOR8LfkHIM0lE2QKkp+3ULNXFvEDgrgzS2bO7Q9FspcIXMuIh5TdkrfJ
LgNI5toa3udqKCCIaGyhJHyVSnXOuY5CnuTBAltwIeFDK3aX6rDUxarEEAPw1RTZ
70w3fIphUeH6KRe9rKyfuU9ZG3BVSfbvCSCTR+SXEoLNgfPyVclrmKoqAMm1CUCh
a5tA/S/K8dy5j4zcEiWqxCthFgPjdhA/Bfho11ClbCgC7xZT+9CHq/nnwv+EvlVm
EmdzocPh0QDFO4NtCYU+OGCp6vEkvKC/pLquy5OHitYkVNVaR4kmrJ1TcyNYHqkM
oWeIPPftLnfFtXESb3z/v0VC824g7B9/nPmPrnURuSfk3fv9xFBY8TA5+JHR8YWM
K8zBwWbOvjLlUM+SJjQGyfJ9qpqJ9OOghNYi9TRBeKq1xnPcp0knnZkSTcGsFX7o
FwWIm01GNFIz1d2lqq3VoICwhXB+9zCc4HASLq4YexaI3FCZ/iZRL8IRnM/OTMuI
+hJu01lvH4T95RvSZ4tRCjON8Dz81ht9sr11nSuq5KWo+h1iDtsFuN6t90DMrWGk
wcc92m3wT7MCoaCCo2CDMg==
`protect END_PROTECTED
