`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+XiiFNOhBhWvq/3P2YYFiDv1T6+CxSCvq7v9H9Hp0KyM9wGhZan9V/NlKJeu0X1s
SLMAy3Hu2kMNQPlxe37327nLXXUxiJWna1sJSbTOpg5vphePD4ISdhXto2KMI7nF
TaYuS/0s/VWp2jhmSX0O73XhIdntipQseqFVKg5OCcz2PoSs+FI/Xlmdscrv+Xks
BXx14Cz+I5Szy39EBSqkbYmAP0MGTiMJCcMP6ZGtrK5r+1N+jZBpA1SouJh6QYWD
OzNyp4Mjk6YT/xcmJi73MA==
`protect END_PROTECTED
