`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7udqVXLxRbaKcukeFRj78a+ctGL3qWBfsXTbpkbawy1+IQNgQam8PSLNAXEZaMi
QzfO0WlfjE24vkSGn8OCQW60nwl/o4zQVdnTC6F5/IjFhD9VeA2mgtJ2HrTSP52a
hOx0tXHP3ItCLA1Jj2qmYo4e9wQVV8RXE99MauDQLUmB82qaob6cEjEerybZUG86
JfbGV943F3L95TlsoelKc26YJdtVQAvaFVAlt9GIyeJ9Xm7KiinUi17FftXg7wJ1
sbagf8hSpJs4DT4OfHSL7YEOiuiv0l/nB7OtAjEl8dWomJvNecKo1ZM0HKqF4YnG
I/gU3z7698L77LMOVbAsBwNFUeN8IMiXta7odsroUtxu7NE5GPsvKtpbXLnWWSOt
zppA9R5AWo2acsA9VqpbkSOjpnkyNVZ4sjtf6GZVW8zr6m4IuW9rXfypJFhXHbyM
sfU76eN0v4C5W+IIV33+ONpPTiz3KaYIDC5hTDf440HwwCCLVOEYrkblcpmGSX1s
g5Mn5tYr/TaZA/YEKfjnTZF2PvtsbyhjJaMMwqdeUKKEIzbZLLfVE+Bw6zXUSd1I
`protect END_PROTECTED
