`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TUgIw5ISiLiAgrbYjDp5t67sTiVNyc+nbp/MLWg7Mf47h9brb8hzAio7n/8JaRQN
nPbOaS0cNO454a4hB7UujMaAiGacbCoAcfdTGIHPl2Ej3yUIhmVh0Y106vaPUOES
DJNw/owirsPkV/bULThbUp66qn7VZPQtb9sF+/uKUIl3GNckXF24oz3UBH8otapK
7TEVSiPnpWhhD+PDNsq8qkEqW52eoq1gp6CoX0dLjO3uz/TmWGdhrjmeW7GjvnO1
WxHsPcAEI/oThnpZdiuu+F1JrAwAsYxPtrrrXJ5GzjyokpzQoSSUp+waZXdQao9U
z0pHn+2VQexfU5rX+9EzAkyFWTHRmtIfG+3z5WDO0H5swhOgARpvbpjV12Vdf6tt
`protect END_PROTECTED
