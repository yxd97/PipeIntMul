`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUwF7pSIfzmsUP0MTWQmTnTGG7eSxIQHPHgdq9fpiMCqwLgWEnRziUcmc/20okN1
o0ROGJ0/Xxk+77pqjJkbVmllr1/PVsxy+8enVqBD9Dt3x929G63OC5wN0C61ho4p
Efrat5tQMlNb/QPvnupl81snY+MBlzBahEBWzMmKPmltrObCOHuaR+VLorwaM+yt
4TU2wglLsaV/phOQ0/lJGn0uwhp/1XUXtl482TyxknIlOGKivyWXKu+vRNr9V4LC
XAMIOLWEsryzZIVqT3Yv1Bd5w6BoFSmZXJAJMltGkyuRm5/KQ1yhVjf8gytNygW5
RFGrspeQg9gfUPGk94u3KYYA8nQHecwQMyMjpTS0wcmqMQWoI0xPKWEmBT3mlMea
iukthe7uk7/U0KS20aRE0lo2l71Lro1uKo1u1IxohRTzVZg+e+2cQOafDJHGLA5g
hvaXtxLkSNyLOD7fh3jV5M2vOm/lHZmzCaJslgQxvWj6yaX6iptKnCU0EH2w+3cO
oakC6wM8vr0tPhg0slWASmpOTOv1DKjr+uBg8M7X5ej3KgleSlXCpBxD9YIn8Z2I
FEK8SPS1fGdTyCfcPfDQ/ZqYPE/uleBaRMRokvU8sDe2OKp/Gi502hQhjzVZP2G0
cUoQ3R1+jIVDapLSEdplDBmBsGBELZLP7GrFcfWd9T3F3mhbwUvxqb04dzq/E9tn
CHjc+DBe1QyaKpmKBpZRK45iq9Z9/3i19K3chpUMsTiZMF+34T+szbM8xZEsGdUV
SNDdl5lNhERLPMSyo4EIgQ==
`protect END_PROTECTED
