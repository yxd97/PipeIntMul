`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zkqcWUOC4mU3nsYJIiU5mBNQTZ8UrPPnfY5Aff+EVB1HDTnCUYLkNS5hjqL5f1Uq
8PK/+kluqgZhy6l+fOCG5xY+SGfgCkM8aMax57HHjsIr3x+NwMaO4ZjweMFmLf8i
FEgGh8UekMKdq9fcrlpHznkcDYJxtFbA2v9WP8tRerEgWCxc5Qwx5oencHRiXYfE
ajoFyUkMpsU0cojp/oRtA1YjKDFRREgWlHzoNN/ZRpI8iMEe7wBU2kuL82hFEj1n
SRHU/OpltwpOgyvAMJyjh6TcBKMEO4uFL0QgSQwe+xaPCLBeS+kDdkAsJC6XuFas
yj0X4wJx9Ki7PXr2RGHgeRKKK1Pd4mTsGmk9fh3xJFjkCtMD8cWx/t6tj2ezxRtY
xGed2VGWSfDSWq1dAx65gBiOUkQzCQq7IDmAtcRHvT6FFa3vwvI24knS6ckmSSdH
/4dt1EONOomR/fPx0VKHpJLUa2kbje6lAXBuG4xLROPDDlKe0OZndXvAHqAnp9P3
WbyzpjnIFx8jyjqFmu9iCK/UrH5HY3OjvBaT4nVXC1aUmXVe+CaF6RVmvqzuiiIU
`protect END_PROTECTED
