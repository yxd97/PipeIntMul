`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wpyzKJ1pvKmrzmRL46FqBRO7Ij1QGTkLyXmTfFf0T9VAr+4mgk5KUKsuyoipIki7
HxVGB3sYNBc1YaFzbCOn11kycgy/PWMXJzgW7L4xkz4yXfoyIOA25AxdlPvvm02/
f6Y2ZMkdqB/0DeiTeWGn9EFowjCVVLLuGYb4PPMFu+QLOdayn7H/0CdQd3/ROcF/
HAb2Gt/Fr9C1LtzAnYXTkdwMIeVqJA/Fe6Hz+JmWVNr3U1UpX5l69N/x+b/WS9nZ
ecPOvZFWVe7zGui0qa9L88KltlJLlyvqrQONlpZ03458F6BoAgbGTq5sBv+nFrEA
gBKFY25E/mPGzSn4+xlR5+3MLLix0GIwmXmcNSb0FpI=
`protect END_PROTECTED
