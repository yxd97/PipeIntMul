`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wsylF1+VspZTQJoAP65RXf58hs1d9veIIv6wyZva1QOr0vxt9RTav7u1MINKH8zj
ARkvlD/EuU4WmkNS19lFDExDAIHCsWPRQVIw3OIS07W8J8a6Ja+JA8ZjWU4nPn5y
mD9f4ggf5Bt2ejIb5vXbAtCKiRhaHm15wBZZhFzc2jLsCit/sl+xjJsTFvVnjMTT
ospzhb4TmliApqBjBnHOHxqdiEqbf4BZledXpOQa8kdVAvReIaYiFwqqwjswuXPA
js76PzIz80GwsAqt6f8+ZuOzIHcVS35UxjiM9oydv25CAGhJYbwlGDUlcJSl73+5
o0kJqMh+GBIXy4XSGxsKluVsqUKKv1vbueXM5h/ZSOj1B/q3ihesO0sMJlZGlqsL
v0+aTKrfmQVHMSMJ7ALd8RLVrHRaUc8IJ3QEs3lM/cseLwIesDgTWhUbFADLWnfa
`protect END_PROTECTED
