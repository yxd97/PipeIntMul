`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vw4HaipHMkceA7Fyxz5D78K0Ct+IaDuWf25+ce57Ze9oaIPtfIN8eoiCQhb79vCc
LYKmTGQzyQpYJiJ2X3lCWN1tgcJlCPxTEopKsDhW7emTDtPX//JOmBOLF5NO/9Ei
uUskck2E8O8UOsw1UVqsDHLDES98kiUriDhYHMAG9N5c4JAd8KOUZ6CpkfNRCabX
FqUWR3IdgXPOPjz73mIQtj2a9AYQrqU/ic+zkDm+pwPkYx7V2GP6Q57qJYxoCR/z
oO0GPFbG5kiWPz058DjE/3Q6OQTX5XjIAllhq3p7dzW07UlnUkftYy+thmg1+lMu
LWu4wxdBOffWEcpf1Rmbj3KUCg7euz/Tw8dVCYfIp7/zwQrRUpvGCuikGpNkJdkj
iGcmF5SzwVjf8SP9SgpcVaPAGDI1bhvovvH6ZKXsdYn+M/HOec9eM2C54LQw3vsE
lZVYKlcwOyk1HMSuKLB0f7t45cCUheTE4ll/RNadW106h4Ef/iiPWKbFQ4JYjMm1
FHVcYitg5kFwu/GptIxSpwbvzR7Qoz68b425wT6s9Kfg5LH5DS1SvM0kT9cXyzS9
oV/Y2oY/busnDJT3nUOzd4CN7ByrtZsbtHs/Aq+KS195jvvL7kcuqdFx0FOHm24z
E9iepHsS+S540YcHQGwp8Y9IdKqCx/VgZlR+Dvab8v7rTanPVn1M9B26eggWkXwZ
GtpCoHQBY1F5vrU6VYvMXfzv4X+m1XFR+MYeQdivpPUWaxiKrjdBBG/fXiYL6hFR
ZfVr3S5XqBZ7snIH2ddsvWRZ5VdJ7H0ggLkgcd1Mhj7zinRyaLAafckC6fR0zBqg
oJPG6fs9Oqpb8rScxh36F0XieuRp7+n+IxxPxDyCt8b7obK8LUgzOYjwy9lKQMLF
`protect END_PROTECTED
