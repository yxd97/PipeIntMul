`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vfgT/Iu4F+M4wEkTZmFFj+ZeOZLTnnitdfxOO1mnC4OlePGoGmaQlOyIjSRUWLYT
xgh11N/ZXqTvTRwrYHJ4Rpr4K+yvyuo3kQtI4aFr8eHRp+5klXDY6Yzlw048vXl8
UQArRNlL3hQ2WwwBYbd+qy3Zr/X3c8SjeCfuRlj+TvHbUFof/qs96CcF4un3TIf1
qXKBhealgLwlClQ0JONvW/r9cc2fQ2KnBrypgCgoy0pQQ30mzagEYwuYmSmoi9gS
q6hnXnmWbkzBrOLFdYMlagizxQChlYCe6wqTQXAE7bfRsY9Xmx0lhw6UYavyS7rn
3QfKI6iK9hGtW+sE92v2Vr7VXfXqoZqODx8azBL/fMgDmcg/mPrqX5fwD7ENJp/R
p3C5HyxsPWWOdnh8IwOswNBhWbmhaPQpH4rs9T52zgSsJpHPEiPP9KFOz/CtQeiD
U9BYp95yuL0YrQExku/hNsYYqEKbXGolKEhuZ2x9QRhE16x58HSBCsqGKbtrO4MW
vYSzAQU9QGMFlUwA5giVFwzcPnYlqZeO2i4RGO4u8mT2tSXwvEBmuj0FkLMeV972
zuK0ThKuhImT74p+uJAc89osqN1toOFeIJWU65adt7TjQJvRDg/SyHDcZAq1Wl0Y
x69+360lhNgBzO6d/RcImKxWP5V67uior0q0UL914GYRiA1zunb4H9YasTZ/yRK0
cmf2aRh445EQk41Hn2JexL0WH28DdRo1PiU6O0t5Fz7BjofxxNJrU9Nf/XQVE5zz
lIvjju5BI82c7eyYeDiP3lQmBfELnYfShJWXhyp89747hqxMTohwD1fUU5NZDI4G
ggsAUHH7m1HqaWhf73vh7KRvYXRMVT4naSG/dGqr8LxrDYQ8yMPDlkSqaOlNhoGV
57R7PB5d4Dq2D5KEFessVMOOBWEtgxRzVuOOX5uv5XDfAa+VLsTMpyCobgTjCv6D
Q3fndy6doJhR25obehXnN1RbS2caDmchMdLE4OdSzyNtpXJgQM6mxAei5alh2904
qI6XeXvW+k3MsJMu21PPVw7r51UZpmQh+fObdG01fNoxNEWuwBx26BeQaRqhrTvN
LzykYPYA16bNj3PmRGJUXzNbPOo8eL8qFxw4ETojJayJrIp1Pgj1WRa8TFB5ejlG
42WwJs5NI/mthE3eWyJYaRJxiEhEBdkNdEl9d1VoULOtt84hPRGC1VqAM6mvONpK
nAW4xCq4fa5Nmm2+fsIxhRyFYZlfFuznnuudrmexkemZ0AUBpEKjdOX85mrFTYWU
VxBmR2Gv/NqXc5aU+Q8SPks3sBq4461DKPjSAOa1wamYcajk/iesyxWR6TPxpGkj
rS8dpSt6PYPgCLbC43ZZvaIU3reSCXV5ja7TkYIztx3jUmL4HhotIXBYxRdYLFYy
YbBAdM0245ROOLDp2k13wXI5wDr8TbOqtjivtKt5XpjmU93nHy2mgLQR8KjwaqDU
69rNygy6UKOztTyd+3iajodve4zzlCQ4RFdtgfgEQNPYIMfJK+xUnS8oSRzoaFW5
GI3hgObWbWWxcsDoE7Cn9UCNC4iU8HNsfrdo4/8WOHwREm5pQN1DLUbBSX2hBzf4
zo3eBpVTH69n0V8mL4gLJc2Xub9vbBx0wM0lorVQblS0CBOai1Rin+pGo5SfRrkD
ZT3J2OSv7l5jzZyBTIk+eE40Ax4TrJbvplhL24f6Sm40ys8mE8X8xIiln6nmCjdJ
8j0jQB+tPOcb/YngZ6PcrdD31iSEiLT784bKyPAdJs6TdDNPjSdgiTaHpHHQfy3w
BdAq8A62m3yYhqpAVqIG9lS5LN0TwdahEr3SDRWlwjBLM+gAUJLjEdBEXaLSmXPk
AaW9MA/qseswZCeDIHUFb+IEhFo1JCAdcp7Nyu3r2yRMmlsKhQYTG3/hqOb5/OdU
f90YgM/XjhQvF9Wz4XdYjM2hIFRkkssUQ9rNz0C2UVBYtA+dFmkr9WBgwS/ILM/G
RaqcHPdE1k5jAzDfzTI92dzD29yFq759IJdKEZgZaUXkH7R3H/CPZLf9Lntby13Q
O1voi1HvK5iNdcb//RZh0hOpUnEw648xgXKYTxSbw2w9AtbkxwXGsAeTVAY0YnDa
XiI9zmPx40Wq5fhEdJTAsvuN9oPWXjzZbM9wyuMg1AMf+X3cuYNGp/EyIUVwEswf
ENWPQ92gBnd3uocYmjhcd0DCH3UtYW8JCVyWaivQtwdsrlaxCnvJE1moXWYf4qTI
gu5uLaqi0UgKaT2czqMhtXgMi+eUzTLMKvfIMuw7J8j8HNdgu3nBZFydO+php0+W
AsgpE39cBD9ukl1ysTZFygbl2wfwRI0NvS02HGoCtvn7iH8SftkWA+MaVj5ezI8X
67QJ6jecU/F3kBh4NdFuWI0afqQdzpzvZYzHf6LBetq/n2+Md2miVRGjtBwMkVcd
RMC0R9FJNya14AysMkGz69g7oQQLiiFKcLPJF3XKPgMqXuNLaYKfiSkgMd9c1Z7Z
+MqfhkURBN783MeRqz8XdzLk9H3NfEv0IwsqN6jH9QGdBuW8kfizhqjznFgXIIz/
DaXulkhnRW6zCfdsaorU36RPKxVgNbR59yrABOc5Wdt7Z5fnhH7KbvPoh4icyXi1
JcbKFyATTYIQJFd6/grnvhlbaDDtCNTGq++XireXQigLaiZIAK+buYQXOYzQLwZo
Saj02HzFLq8/QZl+I6j2zbWhiAO7VJFdrIKWpk375JZi53Ydc84wF2Jsc1f+WbdF
kc2/UTG46nQ/F2uQDeGbu+p0CcMZXqsbdkL+d8pVz9uXugP4EmgU8pb3MPp7Z4ax
lm+t9ISPfmuO9HZRtEs4f1KBHmh7dbgGfcfUiXihAB4SsrlPMRWjzFi6G1n6kOjy
sSHYrQorq/vYH0bXTKJr6MJCcOwkgEQltRkgea2u6/RL9/l0k6RuV/87W84Pamme
mlZKfkoopW3ZguQ1m/1JnEInoE/Y7DWafIcgk4HJilwWbgZrplbFLjX3iqMg/FOK
yD5kI62JK8KG3/F9YwwNEVO2tAuGYnAgEhHR2Fe5AaP8LT1nIvmXfnOZghvvf4wd
3ES4YXPJB1BcTahRUPBQ38+wC+RN3AfE9YiHJ1oI1kulaFLyUjrU43kULyCbGtpS
nbgKawIiZZBYm+J7jUi69BEfk2gE8LFH9y9HZGGTsLCGeDqTBqkoRueQh+aJHq0I
/DgNyvz8YjWtmkt17ee408HNM1NcLKxkUXkYT8KJlEkTgiBXOKB/X62i13oedF7g
Q5WvwMGD8mnjBPJftoaWN+2CaohJjVrfB06tTjazq+3Vgfur9jtNNiMYs+EH1g1j
GnHUZyOrgX83dzasz9Fg+nTZX60cQOYLL/RMZ5u5nuJ7C0BKH7DMvMPCt/+TFENG
FPcR5yQs0wwjJnyzfvwSqPUCzZGCIbYoWlJ4Gq348rRKXR6Wp01WtuYe0EcfLXBP
3R51ubTzYLOoT2frHAiC2ozw8rPDfm/YTXHEu31y2OZzVT15IabAtWmCFNC4VrYW
t6psoFPL1RhPFMhFWqHwd4qIgedYpNjypUwSsp9kEm6e6wHz7Yd9LMrOfPXRj67z
ULfXWUdGd5vARZThTPOafQYL3+kfHcp7x9nCWQ7tO2fdWV379bjUwiD6OhN5rgpE
92VE47E3YoFxEXWHU0TfdY/e9VNHQctj12ofBN9fe+H2t1N5Hm8uUdYaWKZQXQ2D
bQl+BDTsO14frE0lT1EHrOs/Kk4Ss54THEnZUoIvM0vjOgLF0K6nFvVgob1M7IQR
WH15igHAQAdjQWJvUKi8mdS6aWPcz4MPlzcaUu31VuJwPuw2S7sQo7fWa4+2RbdJ
a0o+JQ+b0G6pwiOuvpB5MFXaxirAySRH90j7WJ/3xd44hwqRBHv6RjAHcGVXBJye
fDhLZRSRsTIkIvrXgNEelCOpNgTQZA7e57ebBxF8Bq3fZyTmnsiiLGpg+BnkyD8E
9lDN2+X74qp3+2BbYoamZAGzjT7uxlkShqTdRjjszRe9qBzjkYq93pXDXFDJ/PlS
fjuyLDDx2KJr04S6BewR5hdRSjbiahhgmSr3QW403HbUUhjoNp2wDhIuEcOXQy7B
GpacX2sRrmQcA/uDO9ERBdyOAI7BryDN4DK4wd6Y0K212XbedKCCpyFU3OO13Qi9
+Hw4G8mUqQaZHk8KXKLxbVdor6JlaqDdiVwdaYXtgE/jW0fQDfqVflOz+A2PlWUi
KkPqLyCqwfgRpudFH23ecipXRK22K4j2Ui8NPF2KYPnkqzgyniEWcYr/h7wej64W
/Ij6lTL7gCrkueZKO9zPzF5CvQJ7o5T4Dviko2lKzI3aa81HFbIv199pnpOUgZBr
gH0i/0zlliW2Rx5E83Qrq9o9k5NFS5PhZ10QZTNbHFZDQzHrQlDPnpw91I4AoNlP
XKtXxgd75x+Htg91vaqaM2hm0k75SAgAOYOzW/JzG1BZP/arapkrftdUXeQKaNYh
zU/esgpsZ7PusRrUrJzWV3B20mMGjul97xKg+y/SQPl2StKaLp/ZJF14Vu+j5X3Z
YJXd3PwcrL8eFYk/eMZMdrvicswlRjRYKk8TfWBGSbPbKfLl03tSQ5ERYRWC6Vxw
+sQEodWfv8IKsVpgqPb45WjfeZDNTnVt6PJPjDOiuI0LFaM9z9Mo0UVnwxUtgb3G
Hz5sj2y+TPOmYEOZ86hdYvwRTRN+JZWWf0EU+L3IgKekLbaD7OTGhKPNMYJ2vsbJ
al8VQZIQV7G0qSz1Q4wCMj8pCqZOgy4uQ2LC13nEh+AeRuNiYG8BOb0vGAuWlOCq
rOeUDgYcc6YuuhEfzQ7vKe2gmiE42WAgdwplIUTMkwgyBfV5JnU5sN7TQBJvB7Cs
+4W28eqwAuNe+lqFDu6PoQHMUGpFjNNlbwq3mChBqguafL+PN/++SXs9vLy5xGCm
O53WbuayPIEt3DgGivgbu+f0SYRQT7qS1ettakLRupWmf4WRcbPx3ULpb+Tjw89S
Qzu6qDjLFf5MD+wgFZkj/CJvbSYAmj1v6m+9enTGT4xk2Ujinah0+6bXE7oT+KlM
Pk5AzKtq7XEbo8CG3/NzWJ2NkCrZ9URefo5Fc7vkAILZZynJeNZLnnlBSE34qyUF
/VAo31LJPBO0MU2xQ4t+gyvGvChkCxlDL3miVsjwu8EUarvTTWlJK9Rf7dbwnN+O
KoNqZnBWXETjLoccEGyCI5Bc44S8cmgzImZKEPySkdG6WY59z6PH9pwCh/JRoqVH
Pq1ykDN74BlHnjbQD+OlnIlmr8hOCLGWtSgwZx5DlJvW1s21wXMAqcsFd28A0Kkw
acjcy6yjBu2KTvrP/MV+rLRYddZr+60oTXhMEPUbz7zySIXGadxUKKLzeJVaF15u
/VTN0+ZchISUMK0zK4Rkdvk0l7tgmjkCRofFUOXni5puzMfIfkrUi2SzrLgb/MOI
Z2uJzmzZ6hNBW3AT+fVw6MTzMtGJjn6nB0WF2a++HwBNCsoToDx6Ym46VOGQCd0K
ULo7IDPJI4LAjp3Bu4HNjIPPyIDSOSHUWkBOSaPGVgAVTbHltvMGNMuUTxWO4LmA
zPycX4B5z2PNzXy3VVzmWkUx0tfDtAU4C/xnaGp+b6A0W54CcUPaHKnpzMqsAjHU
Mks0p9pTTTr0HQEz6GWlj42n2z3WrmsswUvI9rj3eAfscusk0LUEUA+7V+FFhlSV
DbsRMhZS4aOCtEU3J/CXksZDhmn23yFPKu6IVwOi44TJxoZNS9k/SjKYhIewzizG
IKUYjyHRg+IUewUhxboF89NKZnHubdVwtQmDQGi8J67x+48ge1YM/Qyn8gt+ycpK
BSy0hfuNXQTvLhtjbOngsqeAu1gP3V4rtLcHkn46nu6masp0pvJAxMBcCfSU0occ
PbQf/cG+iFpXe2n5UP0SVZjcnS9AnnFvF+0xvO/vuXrEa3Vny+ILLf6z/mdwDQ3K
r059Qtv5AZEd/TTDT+v64yNOIlJk8ZTmcg9UCI0iLVkmCKPyEInFqeCHsI0dy6VX
pE2IoL1yWejDp8AECw8CfvN4CyPT04sku3j/pOYEzYtpvCa1uh/NUIA8gDROA8sb
/uvtkXdYCTkXK8cZpoohq0p2QObqlND6mzN7NbNX0G+VFTEhvDZ8OiMc/YtpuIl1
n1rswpHYsf6OjvWKO1gDQLBF9znYrj2qEo7jWEi6V3cwLfTolDL+2Zcpourqayf4
k6w087vQv3VUhOpcL8ZOJ6gwPY7mkYWqRPwlJxjA+E1y3HXUVX66nIqzxsGn9R8z
srZJUtfriErXCYfk7ayxdGt/scMi97ES3w5uS7sbFcqrwau6yhmo9uWs+XMQcMyF
0yEEDyUrDbepQuUodruVdVsuE1vin8pEeUiV5BokRPH0a6T/J7wR4hvyugKW/jzP
/kBm2JD5GMB1wf8Hlz69Vk6TnFc1f233PcI6TVLh8jAO1wtf9a6SH23a9j0EDmn5
8WT5lRklpfg6U+TJrdjgM4/R4zN9H7NDOIDR4wTVWr18iFNrNE2/2/et/nE05oq5
wfalNWqWHsCYvazLNRbTeT/VlYIQnGo41xE3qa6LzuTI9McX7u6jIGVkXnE+9JN/
krF6BWMEDBe8cBpYIHrWAV6G9OVWnqWdMPY0sBxmJeSDFYhpe4oPrmV45Ffqz/AM
Fn5UJx2jQJOL/qZE+oMlsMk3CSax7QInDRylCRe7/sMPsUpd/1Sv1j6yXQOoGzTF
+YZMiN7Ds3iL9AGQ8DwgLRGY46ygc2QRDl/JP0xPldS/XSQS23vJSQLl8xAKrEhJ
R+qk7NYs8mCSMj5+FbLQWtFFcayrvvoivixNxqsc1EdWT7iqosrwrtKMMcBXalS9
A9/Cxdb9ALoPkr20qCx30PrCX+wPXir0hutxwB6sGcLLD5h0DtrOB+LLlW9ROjiq
wnaT7g9wuozGY2U29LO5zcCk2yDWOkSQ2aHQgg9KD0V2MZ4ox1c1sM1V19uFuny8
8rWH/ag9VsOkYSx8JBQIqKar+Mb5HA2T1nMKuoQ30/lrQDwpmntev/7OIKsv0Nmd
6I834iEVsYCkJtcTnO3pXAugPh1zZ1Sdc+dMaSEisy/EGOkHiTn/deYbgbTMNqaj
9ZyXFIo7d327z4h3kDanGYbgoQFd8HrvKQLA/5HCfZ3f0s4/yHvCeyj9UmFuUPg6
2M9OS3S5fEAH8jsImbPvg95QN2nXM3U9DoPEV9e+7dfhRan0oowRd9fuj9rKXV2T
4vI299IuBJmnIxRqiWOBzlvFMPkIiyXHYZDV61n1i2nls/U9TQFnyhmsOlZVhN7c
rr0X647UUR9zRCQL9t0XZhyQjZYEXkwrn3vvM4p4S0e6qgDzIEl+G6aKfL8f75Tw
gbCS6bf83EEFlGbZ0MXtwHGZa+aQZE8z9XrzLsq4w/t6xFnzVTu7v6Nu0GVPkNxP
tbaash6wxLj7NuoK5SOiOqHPDP/s1/Ym5tkSSAHNL0m+nzEPOTtyEbc8Q+no4Gh6
rtSyFgKBrBw9hHRHODEfJVQ4porSQukPKLJ/DsiT6uoH50n7MwpP3ERqh6KXvtKz
iyVt5i9h7KMmyV1bcmlbHXSF76hxpQwIBQQ//9roSg+mMLHYVflZXH1r5W5I0DFp
qZCsC9LbUBlmsf4mBfZ+UMfP22n+o6HM6Z4u6+cb34fCjsv3L50ARBepXlYobkKY
XiavbYspNt0umDSQYDj4J4in1/ZYc/hzfPPtvwLcUKQ024ybSk3SFloO9eH98psF
yKvokm9GVL90ya5IhkJ6GIPZQpe5YQaSAYGgmGIIbv++CYbhT5j1yV7XaVndSuKN
Xn7F+Cv2ebNo6r6ash1hdENaxigtRCO3ffoVwVF/KBpsxi3mB+hCZMZQSC9nTjOH
JjAOYEjFt80dkZ1Lv9MU7DyzzrU9YErtB5Cz41T/yYG9BQ1Ehc8rw0jbRHP+rxH1
vbYiOeDItFMNYjprB1ExDid0LzRTSmVdYqJ60YTHrfEyOmayk9s51IqhXMm/XHz0
/uUjHyveoRy+weTsge7BgIsHaGOXAJGRcHlYTKw+QrbkgSpn/VWNHfsUbmAdwtkK
WCH+vR6BmM1TAx9qwkGnBv2SGDbWDpjtt+HnknNuKisph+lya5dEUZVtNvgjz4m1
XFs+XOsse9xolYrZbdwFUL7JAhSgLCBxpguqF4gGq7zrgVjHB5PawuN4RRgCUB5C
kEn/xAnpB2dVagELAbKXqnUCHwO9ou08oTLOhhOhE5x4YfJ7CcNv3U4/0lce2kY4
Vugqxcg4p7ifCsZZ1pmGZ+2Rbi+TDGKmqMeiyzoGsMibkowC/PiEZeaxN/xLVWzB
IvozcCxBRIaBTQ4AovgQMeUX6tQN0JsWBFd8kdELerNbE6bBsWWoE7JapersbpTw
wX/3hym3yGuy34G+aI6a5omrvSwPAPMO92/fHA2nGRxHn5x1RGvvigmkpJN5MIyW
sNUxBHVx3/OTT+BSNv0VV3Nc7ZsX6AWhYODaahTymVyketNupSntwX3cO87NG6lS
9GzmH4O56oQhKJ7oE9DeNg1/rHxQz7gV70V5Hud5AhwEig4vJJyrJMgkm1hkdJVL
UND5rKzbBVk/f5P5xqAS4dNklyF/147IBBAmsZJvHqP4I5Hm8AmYMv0fggCAiv92
F2Jto6yxs3Ao+ngCbwcwDWir7v9AqKlhVudxg5GYxIBccWg66IH2fnST/9XkSdMQ
hOrVgTB3VZYlmPbstpmKgmqpCa1or963weGqZ2RkgeQIpIKhzazEjjzgZHfM43pI
hDClOfPb+TK5KVF5k7CetMk1bmerWEACkgp1N4GdleaNaU99gaGYhoczWBqjVJhs
+vqMv0rfAHFd+d1DbqBO0/bVR5jiHOYscEr8adbO6r9cDrYzXv+Zn95UxZB4pPVf
wOIjUn3Y31Ai8TUbRmUstCOBM4Y7T40KJ14LMzsXJqYCe+kVnUdZzzRk5/LD2o3u
+/zWCFj9pLlHGJfrjTUwt7lkWBULfu3mMtWsjaunVZBftLWCvajs5X2RW8/baRWE
/BmiR52sGZlEqw9nzjGxeWapQcpKdkcHYQ9iCop+FXBiF7FdB5TWyNcK0QcRk8b/
1X2ComeLwSgu35oGdJP5jgUyytEcPp8MkymcHe3TwgYmeqm2U5C3sosbwqvgSSOJ
6Q9sj2DnmLN5xS56mvB+N3oV2W+c64f4+yukQ8V4Z6WSKDLDKMwECF0sULvwu8uJ
YcGuJa0OgA4zwRqbpACXdLEmg7SEZA+vkICKmAZSHVCsaevRrdF6ctqbMBTqGdhq
tZmGk9EsgB2WtoZz2BpM7Fw+6zpHfauz0st8CllKz+svj7kNoQ2xgOsyhzmXTs3D
pmozwi8QT+CR85pnroxYQ0oEjQg8EIaGmDQrUyPtg3WoWFSiEKNt9XB8+GvcbVvb
8G3kC5i4RQXXQVriVr9R752xWUFXuFHz/bXF76gc0s8ArGzsuznUylD1RVBu0vq1
cKZ+AKM6u7sNAnaZUfZHgKuqfrOUz6S+HlEYBrTaAiRmOwQjfb60Ua+gbJKSVu0/
7IPug4X/dLnLuy4+c7fgRpinDeT9dwFqHa22s3LvckO6ZRPRZDHtntyYVGGqWWeo
7xykkmcw84RaOEEDhXUgBBXAq1NXDF1pI98eWxM0y7qC2yFK/NRhvfpLA2uoA+kL
AUSUw4xpDVyJ/alV1rJCa0vIlhwcDMEvmFbItMFO1AdWodXj3gonWY5TkXmFRktB
lNEdzZu48GrIm9Ox4gyVLQc+GhoW5ke66WwO6Kb6RvPdUJgjd1VciB21dU/gDumq
YaI11X744qrYnl9pZRYgqs3f6I+RNy1DhPJGjXoP6pPdJVgFG9NrFGQja4r8xpmT
FQleuIZBI8/TvA5gEu6sSzU8AxCTT9b2EtF48luNLQPWzjU0O2cbnFQxpVbsDSe1
iKx2H8A9dN4N3n/gKTGBmMdds4hXdxNz7hzqYDqjU8wcluOQEdgar7HlxNVroyZ+
e6H+kcKoEYxSxp4uujcuL8WDFnot8ibYnAFDwvjfKs86XE9JdEtdj9z780zmNPRq
pn9FcK/D/YnSU4cn39bOK8gL3Zm2i3W5QCG9jHIR10Tngdmrm4OTlPnZibkogA1T
UlJNma0t8NzKwwRFlxetvRaZuJUeEtcqI8n/KfvrzRCCBKdIEWCtaIiEuIT5IE+p
mAJLlRw84KZgVoEDowjouMIySdXlRp/+yTykn4VTa8ZL2Q2By4r3rLeCtdVYjuMU
yaTXHRaidMGQCMJTn7cHGtwGYiEHUaUVuS5tiRlOrOppHDAOAr8iNTuShnHO6yMA
TynEZLducE25EJDagVf78j+PSKIzIBuW1e9MuCRmcTQ468bi3i3JaxU5eL0bGcct
P+z18ggvdJgliUvNQSXPgC0YEv16C41r+aGJx9qyhLdFrAIVDomjPQE9Np9ounQp
8fDIwmyuvljRkJJ+UeKa1b+ZAvSaOPOtPh3PEPxdLD1Olu+ljG9aMp3HEEPlSXPZ
3BvvvaJiE00lt9kpYyuaS83rwuq4E2rsrlDEzphvByIiXthwd40RtnDyVh0nX2qL
hPp+aO1+CUdQxamLo+mNlsDctZn/OidO4ViUsjw5JNe2ojp/5OWCGPgBumR21x8Z
tCqTTsjjycYibb81yGvAf67uRYEOgpVDS4CO3N3iitm8F88OqLaSRu7cEYsAk4OT
QijrW6BorwXYuVsao/7cwBTVemwyroi06B9OEbPlaguKSFSFQm1Tln7TYysY8ze+
KlMxqcWjbpf4ZQur/xOjBE0CSqViU8CtFJcHj6lleK3U34vVpBWJgd6zyY5PY66T
AENEsuidjoW3A5N8Vl+u8/k/mLe+RpEWSJtEHR4v1pPGgbzpiiUIElqutS4nMqmd
yDF1Junp637quX3anmT97FjfSIMqdFAtfUcbBJCOoB9wqKDpTrU0cse0sTu7cCBg
hHyWOU8NTdGARa861aIqvw9uQOMUfyZXiNLqtaXAsP0apHn7/R0ElqAZy4Rpvsc0
WYw/fc3yOLBCBDlJejFjiVEmQ6ktFCPx1pcM5lnh6XH3XE4ZkZXlHpSLUHL6XEG7
MNS2UmzxyTjluOGGRjCNJRPzBNKI4Frz6/hVPGusF/kDbvI6GLVwFkseF8yfxMSk
rlz2qLIoFtXeEtkiuE0GTy8eAT4v+XNQtpvo8gtNKz0h4YFT8ucJD6KhpCuc+/6B
gRrdUNtC5/tUQExlrlulvQkjg9cmq8/+AZzpxTBo6LMTrDNpm3p4ukOJExfNmZrp
PpTZmZtKC+UARBT3PFC1y+X8uLt0U3UAIgxyAZgKXCbCoa9WAmOU7doXSCARclq+
9uLz5pqIrsdTY6SvKnO8bGAwY2cyjpaCF+lxBm1ocbb8wmMhMGUYzBtvkJzmiKVc
Gxvp36cVCuLk9R4a/4mV/sz1PzhhUxyltyQOVm8BBYEoSfogVWDHu08kKWxoF9mo
QnKJzgnKjq15Bi5TjN2Gnikw7TIkTY5Xd5ZRkA/y2vv3VGTh7l21ozPO9OzCmCME
QFsXsV0wXr9IJoYhFg018vA+89/2o0wPicETE4Q+00ppYqpul4PvftdROzPIi5cX
0PStgR5iXpKPzragTUdya2A3+QQLJH6LBUqkLJbdIUSj4TQWgaE315FOTpvfTeD1
2CAFmUmtr2ibU4/XrsCThMU5WEWiIdu8QQi9c70bM1v9FfXa5yQhvl8BAzwUivKg
rV9/ph6bjgdidDQSGUqfCy+si5kdn1+N47RSmun4yqsxefKFyBOUcw4udKms+BD+
G6YDH9Ik2hWRX5+evZakHwH7CLTcojsuQN1pB/1bhIKRCvNvPDdxQAwsgCMizy8v
m25BzHjyUpa6i9mVhsotexEVqGKbxQvFSl1W94Y8Yd1bcOrTy2KUxOoX+JFnuIpX
XvDbei1Gakcb4F2kUtPunJ86AQE6IUK9rKnybhkWM6OJkwGQ3B3WrEfKaBPTJhUj
sTiHGb4Jw1nAQc62yAgIIlum7UJo6vt5tfnmAQGPNr7sAUDeA9z1QZGXLoCdz5Da
TIFUYxU+HteAdkpWF0KkgCfg0xiDeXyXUqgsWeVAtLKaa5eRJ5AtUBhuuEQ3Httv
x9CraK0Wyp0rCtIujwlqrLcKWtAyyZsBAvx8bwDmFGxXL1uZvwRzNaS/IsjGxTrS
dbLzoUg2eZdf+ycY6Fyp2gAJ5l+18LIroSXC7Dip/2lG8mr67YppkM5N0NV3ouU1
CGIZjf4vnlSi+BUCz0ot6xmSC5bFdvNQaFnr0RDdTc+aYiRZCEDXmg9XcdVVPL4U
kva7J8nn77SvVaT+iaAmw1hlJyuJf33u80ZyFplZGuI5pSA/rjtxeEpeaEoVsJYe
C8fSG/jiH+98MaC2GwQBF1ZcBvrH9uZk09zcK7JSn6VP4w6b2QQEYe1FXecBqEzs
l+a4L4Ac0OSg7vSBfJqft7XVHYBhBYvK/0JOMeqKgw3vBu2ejt0V7Gz4vLVZn3ul
hVbo7fTF1YwK6jVWW3nmJCs/8wTnruv4YRsk70V+vKYFZcKiZ0pE6MVAHw4XjtIW
9Go0CwdSBfiHP2+cEDKoBj+qg/8KHUZZLPuU3m2xNB/yno/rh6qBY7iWfJIl73Pb
xfx7/DN9i2E9mumGTKucU+LUXxMgGAcWEKBq/oVptZbRWUCd9NR4+M1NQ5GfjZ4O
OCNjX2WWX2k80djd3d0ineVETufRt4i6v9hyK+ccK0Nmy4eaTF83mRQ7AsDrJTtf
lTUOdGOwEtg7h+Oh4TkRncr0N5lTPFuRQP3eX85qNzygi3gRv7PXlzshFhtrXn46
y4j0M0BVz1d48a50Ue5igknB2lWq97IiRrCHkLn3JMVBsvjA4+UcBL43KSBUjtXG
/Eq4w9i1R8TUGyhiPZAeRvLlHD80nAutXOsSNf6ClQDm2upkjKp9lXGZL1zjdhgd
hbKKVqwWzhZW7ZnO3dD2dIki+VHW6XVyDQI/8Nc85oK7lt7DzJMhDlQbZc78QlAC
+QT4HHZXgImPvQCrYpU/uYAev34mmYgRD6XbQylbApDZIT0GKhgPmNZy+jD5l3RR
HN4zl+LnHmSb82zafEc3GvAoRdQWUGgJFPYXLPk+VeB/HoUMXD1FWDGGRrMW4kU2
H2eVhnYfGiEKPxH5RBNfawsFiIZ4WxwGv+LeSX1i7DythGe+Q29wsunDh7Bwv56Z
qugpVCEtXDSfucUpnRtm6V9NqRapGHspxeX2dgghJI3ZCjP3Ttlgs/DFbr3HLh5j
lfIj6xHtQCS/BoEJk2Y/5S7kgF2lgxrKy5FRXpzb+iFAjhJSdYKXfE3mbewyuVBB
iL4fEJqsHTgIximQjJUO96+B1AqScoTsY4RxbiwcG6ufJGo9nW3xh4oHm0w/pS2F
AA3/WPiwimmaCnfio3nLZmzAI39TcwGHOBrA6fTJT+QrTisiwuBTEckOMXXmon2a
0IaDJ19tms3Y+Jbo9yXynMEbrDTBIjiO0C4KU3QpLVcPFS1kDN5K1OGTINLe2njU
fJbgYreu45n1LuuxFJUQIEEfQxH9G6suR7ZoahxxP6+9/Y1VDvWrj8r3yofoT6hc
6WpEPrguCVsgBm/uSkHWvrSoYFuVzEbQCnxj94fkHiPtNhOfv1aXlJVEhQMHfOfP
v5fuPMPwExK+kSQQrsSlT0ljBFhbOfCaxqyI3GpVNgqbrisKjkSEcmg3DHjHsnHB
4/hFisiOcocL7sFlUv4m0qIyIybRnSPCFLgNONG3CxU0HESsn8eF02SjejYkF97c
AlOyDrLZmDB+d2FIp4WxyTqiRDUMY3LCzeJB1xaT3gzwn8zSq2hi32uID/cocNuz
MZ/Qv5ZGKinzKLcBNOTbTUSpaK+g2KrUbeNP3HomMxUC1NNnx3obRZawmsFjnd8c
PsmwHo6R5bJ0hTwNahTAdI++DbziDxQ1/XZHxvSo2wVUZvjhOtvdViG/Sv5x18jB
/JhyOD7+BpxF/r2m258lPDp7coTtc8bCe63bn0l5cgNoO40ZE0tMCXgE2ZEpYX5P
AqsTxGJJ5cnCF5Rk5ClawUCCKZWcHoJptRFWQh1/uNzZSy7yW1WDIQ+EQNrF+eLD
WPJn15bnPuK1VlUHiqjuREIbwhkXkDTw6Ex5hLA5usH26xFxcdZ9osO1OYWbc9c8
L7tsK8vo0LPhgj9o5kNML50tIa8KD2vSOiJH4Mdhe+JbrF6bNhwDRN4UOWNDozqB
QIZBl8DzHN/I895vFx0JCKIVtiVaJhJmM1zguSvaqvCVxitUc2tNmDM6ctNYwP/O
HC6tXciw7ZU4Cd0jtRbOa15znxNvhdL5LcHcHFNYVB/aaW55woE8Li02iS47yeRQ
yjlMa7An7pYI9EkynaFkDD33/LeQkZnRsDsEV6DQsajbwAplPndl0nKduh4mSjV0
wbNctDzme3i0MfbgkZJhKkpYbCDddhnwOk/Cq/02rU9g7ktqLJ0x2nfgdV9kCFQl
djQhzjtRY+bkkKVh20wdD0+fMOlLba0+S+hGd1PuUtGFEMG06A0FFKGY4MZsMeex
x2nsNgLWu70D04RCPjUKZ9xf58mSZWnA/B/jiICJ4IIvt7jyrllNnOBQKHn8crce
0zOUefJnu5iR/YG5DepizdQInbPlMjys0ht3uBuJxDyHJniZOOg0w3WCVHsQcK8t
NVbdFcKF83Dg0LkNdKUJpa5UMxFhIpTdME0TormFcW7UgNv3IDNo/299fc0EaDkz
HTgHGalBLFBc1yQJL7dGHwaTwN9lv/AGIfm62EEQ0QK0qKQO7QsnXPLD6kbuckmC
CK+S8PUIano27UhC28f46oqha8uam0+xv+x51WW3sMXTqosRYmEdrMopgofWvN8i
+Ev8pb7twTk6DZ0SFSQyrIs12xoe8X8UJVZ4Vk8zdTtfz0/NO63SlI+VO68Rp0R5
s88cuXsvP2PvaPijZlzhpPEQ2PQdLkyUdbSiVKHQC2aRZHB7CRgZOL+829FcylqC
IiOSN/MN1tcYF0kOVNUWUaY1RQ+PJ8iSRiGWCU2qhU/1J/+tNO+q3ZIeCv9FiiMu
lBtiJtfF8QfCcGZjLge3iBfYMunXq/LMak3EV7zt7hL41WVLtLa3B8H9KxfqTZ2a
LMZ43a9UdTCbLSaDWaPKkeIJvtfY6mOKIT8zTdZ4lkKEJAYEnFSnktu0onzjbEdf
ZbfZ7qE++iyAC/9SCnMndXbUl6/ZgjSCT6u4D4age5LpJonJjfaRLDMZ6QI7yg1m
ztKtGts044EGxzYPwm3eijSQytMciFJ6PUs35dreL8PrCjyCeLz+VlrFW5BiDEaH
HvtylXXp4QtWE3i6VjhJOiEVjLACbOTykeLQQ9Zx5LimvYa+9p+KFp2x3VedInrV
2sbRLExNPHyAOUB5OEsM1snKtIpWQvBKT57r25cOwlzXkFdOKagwfbZ2Xd2qwHFQ
BSLD1mEzTKRDx5ADe/iJEM95nhoCbkfNeuCU1FnzcifKFo5KLMy3wlndBXFa1aGm
zuA2hO9ADaEJ1vy7Kyf1Cb33q8w8OoSNydbL4o1mUmtsKoZsk2uVnxs4KVFT6USI
b2wBVFXjwSz/F6pA9qM2OuFD/5LBXoXqgVL2oX3HGetWfC+/J04zhpI/s1+ofnV+
iLaYv1DyUkOPzClbOYWMavEaz3GqTXf7WaWsH/X35qobQNPuq7JFmDWsL4emJMqZ
ZKbhyYXbHDNHZfxHBrkK+X5lOBLnjq1dWzza+GByFW6DuBlOuTdQzqpjpiK+h8Ue
n+BHxK2wnahzq80QrclT5m1Q6hx8nE39u5iaYkvVXDF7SXyazKSRcgoSUsY9EijG
Upo8JG3IKsVIeQebnWcxZQlf44xXiCAUwDiyQu3X+kFB3v9hYpsbuvdD6j4FeXkX
vZmP2dpIgsUhyvzGWTe6E/uUBUZnfb250exDydfWFHqH7LkXwAqvAdKuiLOAx8RC
W/Cz6YgLuXsxWmxRnqTIRh7HHRltKnkJlDCQMk8R9a5hZr8AqdtpLbBzwO9kAZ77
vLpbN2Trs15MTey96TJPYTinB+6ouAn35Jf/w8AOQGeGFCYjY8QYG2/ApapK6gzj
tFQgz6+5qiBDNkgWtWF8x2ynfIyReKlW7Kgqe4Rx3yRO18j5clhroZ+wX/ZV9/Vm
AyQI18jZY4vz1PfjaGR55uqg82oytBiOsSJSFPXq3UVncaR7zufoyjzxO+RfnaH3
UeH7e528cBC4Cgm7UhxHuKB6uzOYlEwDJ0XHrbSWEUvKTT7unva608MQ5vFxKybw
f7wwbtLHOsokP6+POS0wlPnPH8Ch4C6atGdzf9/P/0pY8iq1pIdS1RYtzkPZGlvd
n4Y3LwCayhXx6aindz6rWdKDMP9ehuTl2ro6kp8s2vKHqLwHCBkIW7/YU45Ei1sn
mCdAWtpfW6M3LwO5Dtfd1t3WyzSHvvl04T+p6Q25HviVUYa4TneUc23sZwpDJ1uy
N+dwFy7ncPR6Vx6/vrvuVTUg2KsolBVMw7sknlD0E8zoiCEf+Fgl2KD/HL4Cuc/L
qoETQ3pjCUfVcAw//e65bhhup9LJf8d4wTistQEJXrnnE8hF33Np7cSHuEFjGiIT
BrQx+IbYsvDnVRsymqykY+tY7xeNNAun3AA34DauxtuarpKjFjbAFvUMAH+tu8b9
AJsWPVL4pWxyp84/0/QksPr6CDe+ukY0LxRLAwaMjMhoKdcOqt1JwSWI8VuE5WYD
wMloX7iWCJSE/za8d4Jb+yqUvsgSgIY/Om5eoGINtxInirJtY1E3uKdFEqbtQrTe
gN3+Y0d6gXB3ez7o4u9oCKR7iFswbUfhZXD1bugeXI+/aMaz/EXBNYpK/mwveSwX
xJ9aBMk1TnSg7KxcfS7D1iV/PH/TAsjOlZ8LfoEZnW+DJ4cwvWqxVmWKxRl3jodg
XFdHJ8fbN19jfQFlz3GrH30gQR8okKqSY7RxV+PP4KM66DlNEDvCoMOxUPcD+PwF
lAM0+yihMYVb4mqHzFb+vI/rbCRi8VG5OZTKY+6ISQ+CcKumpHDSpgLINfVtRQ1s
qSlHo1d8i05SUuCVuB8vKrDGzG8AkL6D0ZdmLtBNJJWXTkCaSrW//KtR02riwYMh
jTJu24swp8tbDAWoZXoaIjxiooLhvNj+e2lFq0P4xxHfFwYFNQufEa5fgyeXPAsp
ar4xQIWOZ6RJ54PEqyfK/7apeOovwZcZB0Xiw/Hyve6Q+VHv0k6H/JH3ex5Y8Fvp
Y2BXV10rF9MNUBgOTkez9uI2EFlj3dtKEgo49qMkLyOkhMnezc6pDwSZLlUFi0a8
RsSZm+e3x+jN5NIftmYb7yS8N15At1mY0f99gZxsYAy0NviBUl1uWVud94FVW9XX
s9ZTUp1dBFCWryuM5+RuH4ysmluQGJS7rtEkWBUZMAaQHjKr4GnE8eAWPR/KKLm8
telnx5fVBLbCsdHiMtiWa2+VfaLgIbr6YeIh4iC0OqcTKo8XpFeBEgx2s/Pl8B1b
JtYdou9QTEM6UezhVvQLmptFr7n03c62+A0gp8TYVZURjX71uKSiILJfV3rLICnp
/Pa2CnYJva3FqsDIgd9IzjLdQA9XsiasgWdAvvsmFtFoOPHR1h2D6k6EmN5eTEeF
yrp0q5Q7G/97/KBEHhGs9sO0tMJcfX4hTpYSwuul2n/Od8L/t7oJ37k0FnPUVVtS
nmoDsm0lGicwy61BWHtu51ccj0yj8yT3ZHgdYi93xUb6gpoo/UcKuemyA5kYolCk
HGIejOPVzl63Wricxqg/OCiUHfxBEWO/eGzdI9JoIaBiRuRYAtIG7wwv4uer0Nee
ef3X7MT/3/LhQBiY9DYEEqPmfB6S0C/MXqTJMPJn4Ju9WNQKEZ7w3XZEFVz1dmCN
BIH3ZqEIEKOKR/DlyDwI/acKjM3SEW1EVAkRwJaTUefOrr/rrN0I5wP6sDMaj9xT
yKWL/K8J3xsxNcqYLJ5DH1RbC6lGVsLTwRh645pcmSw+zimd+O9DU34wSHLg5sOX
0u/cL78KTjY5wT1UIdRTssZGzULGF4iWDU8qe7kTaRqNk5ohnGgZbqn93J7PFlVy
/aSJuwbmPmXufb7b3uVu+WLREACfGaIDi4bDA3HeNE7TZgp4bKtX6582awg5HFMG
mHE74SbGGcUIRMkZYcoUuxuM0ie2rPHmOqpThGBouN0MFGyiluqqZOpzojDyMNk5
dSXnw1WogHpOuiP6vdgIMSIGRpdmO3Lzidjs0lmCoKPUcLKl6P1R4AGQLAHmvMs8
N69ThBnJdAO76i0XzKHXRbzguOCq4kSZkUU41ZhWQO2lBISIPf/LnpkQpls0jZjW
GCBKzI1mSOZ0PS8hJUwO8OaI+AaTDCFks8vZYSv/+VtWZMTcaQ4WTFKLIYMYNnw6
nGOK0LG1tJCioSPYY1dwuSJHfZsSh4aFPtfRCqm1aP8lP8wVH4IlmPiLzATmGdoC
QE/0O6t8qqZrP+G3ddp1lnPAR42mYmSISPRzw5f9V5+D2Dy2LKHs2ngaMvdSO0Jt
21d/yQHWgPL2RtG7TA+PlE2wdiy/LN9QFmNp53slDBhWWXA4BsydcXCI3Rvpi8iy
Lm4TIGbezjPu/zQgn+N94iJdcYeDks1RDZK/JHvBltjhkNcJG821GhuiQLRTdyDw
Rss3t+q4GgcKes/vsPWYjCQ2s9OlXN4+ATOKabIgmHJu8HTVpcW89+sSkRkDIeJb
JXc5geouoYDcyNFresoSUUV8Ibc5HRFdTTb/qz6e7bCN35rv1+tbFZiWuXsj3vnR
PmjCl4rATbdtTCgpmKmzLIH9EVibFFjNi8NOnZORd1b2l9s5HxZCzd9Q+OMRA78t
qSTZ73UxI25RGSJGd56UmTL5uV6wtpkSkTGWykxTSKLJ7hgUHkxVTAn0GkM34/I6
wVNGX1R9LnSVntzLVW37DTKvUHz+lyZMWD4apQqOJjPX/4k97gKPr3ihcgfQFtyl
RsqEciyY8l7YWEOKLJKBnfM8KXf4/P01CL0aJ12qEKluhmaT1+euLdeRGzvOki1J
/slQc5dDKRi45vk/FQGjznnrmvXll4Z4ExR/4sGaSLanCYLCCAYKpa4YgPNxxmfI
iuWyiw0sAwwv4TIxbp4GQjYOF4bI79cIVNMXAb4O7+Nfb6Wzsz5zU7of63H3R7sn
Gj7yjRnFz+snVcUYpD1eGIEURi0thFyYkYu7CPfiLw5cQwW+HJRoG31TeMI8FZ03
nXwAAAPyar0dISc31xOsR6i7kS+mTNcSPQUrKzm2jobCdtAGN1ErrdGgzFsCzlx5
PpW0wUXK1hwB93sr/+7nF7kP/zynrQ2kkzyQ8ArCm5a9Qu5WActxConCIUn/bLj7
+U5N48oTlCvh8WKpU3tq0Za38EI42ue3MW+22qDqm47AkWa+OgUjTmVvjHdwfeJz
DxDMAoyNDA5hdqcTjb4JYg8RAO7HNCVHf9zsseduBJ08y/AmtzAhs0FFXOEznMvg
QFwdgPvVo8l1chSNBeABHDoFVdYS0TTpCsPg2yTsDS3uo9xvtLipEBuhoVyqbBxf
bzp6zjEV0u8hkUy4WcVxptTUHq+YngC0HXWE5Dn0CvLmFAjUZKyBlQNp5402vlCw
7MRwECoDrITOKBRKC6YVQi8ycLrrRkj5x94GIkeVtAODH9+faRDEyJmWxm24W71b
G2z7mJXq5gW+dCDquGDwBXmY60Ks3VuAr/DAFjULKeIRecF3l9/2jPRuuLcvk8nc
JbHUjlhteVZcnCj51iMOEWI7BpOzDSJuZJeqMJrWdowgVLNYRzzh1OEDfRtF/j0E
iOOwklFN0KaIDWjJ/M4COQeMopyW9OKQf5uoZOi6osgzgZL2eGGZaRQxRKGp3h/x
ec6i5l+30MvPrZ7uk7vOBrxDn23P/+FJmnn3t7u9wAkzIX6WCQEuyespswoY89HS
YA1lP+sPpIdl+9SEFDXgHlmjld7es/epXt2TR90x2hOKb7ATk3Cfo7zm1cHrIqgf
UNVzwH+wQGmxbSKVNjaoq2A5qkkEs+HUai9EwJTIxIrTa14jlaHtUrhI0Hcs+WHk
VeJk21kt0UhaX+IMeiHd2A3SrqKMgAvEWSlBAo5KJbT+Hs1WVQ2L+FcyQ51ZVR7j
0L/8GpgEBnfQvOgqFVjmg7+tjAfxvHuFoOrqv9+3scq/v2KTHY9+0zXhA3iu8HOt
a9mhsp69aT6scn40ynQq5BiSly5zM0ii1c2cBo0iQWJ9ENRRcqIH+3TSXjd3Ozn8
j51c/0As5pR2+YN55HWdf1cYit7ZiQH1bYRMGZuVv6n12pGOMryu+HMjj6RGSBYn
wHS7UiwBjae0CvimLOhU0FZ3c9V+sdrWPj8La1ke9EmmMX5iGUxOzmIQZAPQofTb
0qG+VRDVQN9orQ3z1vtjxqP1y/k+iYqdXCnwcz2FIJ52vxRxTKqNgsADByf5V/W3
289YIJum8uI47J/iITDAtqMHdsV7s+f0g5xISsbmVKlJ4Fn1W0rW9XDLUs7YQz5N
XUIoTghCb/+PbvFPPDDwWOtohKihr4gCUWwm70eWI6h2Wt0e96R4kBoGPuw7xPRG
JP0AJrKz/bug2m5ns+0d0ITF6861gy4dNuM08LtorSYSspQZ76nLOushGMe3SC+t
tkmsQ4mMzZmWfW+AtQVGKuhTPaTJ7peF4oElNnVkORQPlazs13Q/Fv3/iQvhXtSU
pJ6frfadVOWgw6lQi6LQIVpe9TE7V1KDQiGLWcrUkaSn9jbIFbVRFrdozUAD2G79
m2Kns3nKJUZFm1qAu9eWtYY2boZuZXXkcOWUq0/8EjFZACG00jOigk+pcg50WL88
RpDWEMdr15kN8UdOmc4G7P+xxcpiCAXOUP1gmDTLxNexTEYY94td5hLh3cq9IVMF
yO+h2q5tfY80TyN/NBs+VSOgWNMdQD7Ybhx9nNeAvFevfy2SPNLGMBUdENNXuLDh
eourd1oMSn16FA1F8ULn8CxiaqAL00+EDoxndftG8QSZCGTAgRt2Y5LMPPzlrwAi
3oc+ev5OEvSiVVDvCgMvGtlHoBtmbk5GDRjyfm5WtEMJhC/5ZReZOdm2joEFtSEI
gxaYcbeRfNLFP+lhQXSVdg8AUT3MafgsHNmgLFoorWXfF7zWqru7cjI0hxKbnpI1
Sah9sQRYNlPc4ehgFEDKLMOgo1DRIurKv1+Byk9y9ElXYsXop5mK3Ee7hJ8mNazu
EpheELM6a3TLvffawHMzplZDVChFkb4eW0FJ10KqQ7rQpC54LD+uYFLrMGTmFgZO
RXmd89Cw+bfnohElDdi3ZFPA4rFj+H0SwYG3P+CQzUGHTWYqO+arAuJ0jij1wZ4t
AEDHeiBJu5YuDieC3Cf6gy0gupl+rTvsSPjdo63oTCxqJpxfrTrLPr5R7u902BK9
uPdhqy+1Z1qwlSLwYkwrT9hDE6bOneIGk6MdpjW8cpmh6YhIo1/tROxw90TSukgZ
9M52+MnD8X3MRlMNU0k/T6Odq9xvDGoCYdSRPPJ5j+hvUvbiCvBCTUlIFEQE1v0e
t/d0rIYfKM/rlm1q1YUoq81CPQkmXxstGltyOO8OEcTVNh+5V/uAmXvpncgHCgws
zksleoWDZLnpBR9T/+jMoRhAhVZDohTC3zfngNxCUTROwX1rerG1kMMSIqpr5ba/
XCyLHLSckswAikY2cBH27JxKrbblHDBvVejRvHt1wOMJlDNr0ZjDJJ3eTvODQNGg
AlsE1UScvkdBNt39cIW2sZfWR79Ty+IJ+V+v0WG0RLHhfYJuNnbJ7P+WPddqHaqb
JeZJ3OBwdyWpu4T+ju6aW1SZD2oyHUOZeAlj4iYvASq3uH+ewhngvJu/Yh1hRl+5
o7Pk34q4+l7LSaTvnIZ52bbcGbnlcuIuX/u2P8rqVDnajoIaOv+8P8vWWUmuyUqA
xhWhQXJ6nc0DRgpw90QantF5SP0Jbph3CUm3LhmVWPCOkIpsu4Vz8kPj6B3yOKyc
WtMoBqhqTUx80CtZqETrP6bM9j+d7RjSpS0SLzD/GpRQfceI6wdtYdY9NfNKlJY4
72UB+XM5T0dTGNPTseUiKnYXWboA9T1qU5xugGuwTOQMSqXzYARLrtPPNpObvsu6
klfpLjmiah/Vy5PnN5IMW2mZAa9gDXzrZLU3lTU3UtRP32kWHhVA394vhzifRbsz
F87NbQePf/vnj+p89xdscZSI8QgNvYkL82qoNrZA/mUJsqvCv/wrT7YyxhOGKpyO
S6PIw3HJN/DdbUowQd7qVR2l4hMBYjpP/Ln7JoLFhxCDkmEX8w8BVTpS2IrlXZuz
h/jiOXJIR+PYLQYaZaw/PjJSuSs0GwqbodwxDWuS2uQN/CBEHC0KTDLj5hppV/PW
ghObr7eMaOidYDxv/8F9Hc+W9vLBXaWWthjcUyFv8oNLFOE8uaw5OXMt4T9ljZ6t
DzzG9HLioZ1A+kYJIEhgkVZm0fwNxOFxI22E9zCgTznTzDK3as12hIVgb5p4UNMJ
VZEGbhovO2OKH4tKLawOfwSeUANHffBeDveEVAo7gozfOp98irpWXJf3dokq1l/m
gsUHEIEHQtqZleXSZfEcftAu2pGmL253uzw1hJJSpKF5H9SQhMfRYL9qTSBfEnL0
N+u1F88WRyseys+WIrno9uPIm0R7WfjIdsmdDNl4oYvbwU8CDVhYUlBtrRukghwG
c56QLidR2Uid1NOULVY/4c/phyu0ngKCru4m3o9N6OjCg7n7kDAhQyTIGsvD9MqC
JsiKMKvr21a4ElxNBuqcyepPqXG36/53jJLng2GSmSHEYTWOtlPRz59ASWixI3Gs
pz64RtMfuJ1B1AsLv+aR751UlP1VTvBo/DAtuivFMFjvcoUP9ErwoWwdSEEeJD9f
N7VD6b+VDNZZD+Rd9W6d1BCfxsqpIgJX2F1vvMwm1pogSTFmwWf64BWEsItju7sJ
lUZMr6FDrnX/rfYeMEKuGma80/IFgTy+4fTlDI1vWguyhH4W4xexyCGpag6eWVh6
4JLvBC68iIRvrZnRNAgQ5l38nA49pbH3GxDiXPZ3hGbn18d3Js8gJ1m+1Pjlxn4u
M2TZKuxSaGRwhYaJIb5PRbNQjeJZmvkSw5zda+ApdeqeNesNrR17/ogl/QKvLoEy
rUDVkWDcFNXwez8FbNIyNkqkXuoyR5UnTOcqcjj64M/UYordJ+guxUL8J56o5NnV
T5xg1ZDuO7Q6nkmqXj83VaF2zQw6HisyMwqpLiDG40H2QynUz4vyUSFb7HlMOEzW
7vwPAqyTSRRw9eOkLeDQutvyvGIcaOx8bZ1ELf45BhS+XdJJggZMQSrOD4SPnyxI
KQsJgb+BW3qIUevoc6+0eLsEUtFCzbQkm5KzfZIxxkSNw0s+5CPEzFDxU2f5apWR
Qs/MmFuGXMuaY5D4+bchfnr9KwUFSahF52ptoqDWcyvHnClwXn/Sq6mwZa3T6jH7
vnsG92ORQDhFDDuJfJMdKCG/S/j2b/mGBP7NDkc4rbB4FgNhKaogyJ7ojU0CFavK
UQywd25NpYJMAO4ohZbxMTHFkCrW7FFG/QLZjW7phbTA4lxhGzsMRserevbNKTiT
8AbtBMxBgBM/DgyOGCiLNStwCRNOMYfpyFLISdshmt0NgRxTQowAM4vgIWBlWy19
/0u2/vTrUTLVk4oILlhKFi0rTBm9qrT1A/Q2ATfzxKgVbeocCwm9SKeuIHQULk8/
qwzqbHOwnTqcGtqpfXE9ePcEW38OP20Ob45IGahFKdy8lVrq4kcNdZe7q0swDjla
/aeL0WYZQhZG49CPCJ2fpFuupxkGCZEYIhL4sg+FgO5C7ROVGt8dEoqBMeStW4Uv
FVMkYt9ABCIaOo2fQg8e+Nfkl4Tj+Oab6MzmvQofjhtL7chFrnsAkeZ3BzbX8q83
AJQCj6m7sE7LGwct286HC8kgN+Xwvjvij4bwhz6SDfttMk0sOB0HTc+GpczTVs5a
KOZQpGSH0ydWqQ90aFilTkXfriGoLpjzBMmGZnmHE5skoRX3fx5wGuX/VR5o0d26
hq3Gbp9D8W3qh2915wPV+bv7sZNtH0LjHmvHfiBwentFDA8sjXkUcBbfWctyslW5
59GCor6Y7jRqY5gf0GVBz3Y++6Npsbhmpj9m+il8wcNleopdGM1TOhxOhsOlkaeA
tlmtKz0G4nNi08JniB/mdPa/nxJAubE9uOG/+LN678lcNqrJwstGu8kjQ5/w5Jb4
Skt3Ddfw9v06PAfQaxE9TVkTbSUF0bGhMv1dp1km5uMXaV/BHXVSDM9YwBG+ukO0
k1NnmRWPtzaLXQWAOu6T5rGQ54s3FqztlRlmzvi8vlf1kLd+ap/bGCxg2vvWbPIa
G9t9eKC4q5DyPREs+AUHYk0ESYKMysTzMGRhu3r8u+Qn73lvKqWGcCiUxbQbnj2I
nKq7T0/EDB/ZzecWISoC3kDV4OL36MtEbUlfRuwf418etu8SFBn0ToyQBRtHLYsi
M563A46jgWPBIeu18zUAAL+EYUpSPxK/lUVrjuOKl9OAzsVl8Ny8g814n5vWY5mi
34kWdzsuiCSEUJ0g1dzfDwbKuTgQgTBnxFZxbqDA/Qsj1xHPUKwBP94uUH1GGalb
fdu6G+m1f4TKPPNF9i0A5Fd4+GCAGTfMJs18eaFPMF2VXGd7Tq0nEam7Mf5lOJPV
7j6Ng/zaAU88rdih1upBLal+9SkaMDQr/6pjtisMSUdro/itzbTTQGrjR5hMB8yj
EbCMe0XqQiBt447vArepmC0+vklNiep/R5D1ZivH7/0AqrVsoPKPuDZcQ6RUF+mw
wJJf1apg91Muje3gnDw2ZcrCxEmg7o763GyeqGU8IuS7W6WDK4zBOo6u3w+ax+z1
KJMr9rpAWzIP4Yq/gIPvUXNqYGsuif+hFxHOUNZTs4U3ZqP3WmG8+IX+pv7ycDzY
r6O9V71cioEJ8yD4D4NWOwfCGo3TRCnCc69VfL915jDDt2B7T3zBYbQbF/MPb/IK
nWlEQQskpF7MrM87f3Wco7CUKwOGIHFOY22TDVx5sFMROHdcG03Fieg41fTGcJ59
eflIMGFGZ6WKbKy3Qhz4f2v+DNn9wOS+au1IIp5GfpmbpTSbLzfMx1XYMIOeS/VE
gX68RYTki1sgqHOVxxSauwpuflfw6NW3xmsrvok4smbBZu/8mW3vq+2HuBC+69FA
oOD4dnL+CGLbZcyPSOAblCwdFm+Jndn5FSOK7dTeP+USDDNLKqaPoLG72MD659g4
/jmlJhnlvRGJmniaZwd2PTNjNCtLKIOIajXJ7CxREfdV6/+KiUN3khYn0a/m5rsW
vdmAkAM8x9JyQRTjQDZM3DlDAyW3lltQBy9LBWjFrWuKn1GlsEQGORuuOUpCjRHC
QV+q46YtSvvLb8kRniYeH9/ACZekfaY1AyyOWhUSHOuLJiI44cr2ZnIyVtyM2suB
mMUPs9N5I5SGYJWooFS3O+pwtr/6bCiRW0oKSGVMzDG1FVKeiG7zkf4+ZXX/AAzn
hDpk1826dlnMi80jvKOrxKi2k0wwj5MSy269CcqPZP6tq4yF5QhaEeEC+lKOWIpH
vPWv7Q0lVzoIgxZLm/NM6u19WpyWjyN+y26IXLK0GZ0Sv8w+SsphW09UtUXpdSKr
+Ki48CkyIAa8mHWvrSzyXZEOWdRKwAQPAF0dt0xWPKonKeOKhAQNfOe/uDpRcJFx
jkcstqTuvzxj3REZHVEQncZ47dHA/78yHbrDpdsFPv8dGb+pEkgM9C1PRr5IcHCN
vMRc2LZR7m/ZBvScfFOmuTxp51gL6sK8L4RPnmzpVIWdYb0w1wEr69PD0c0NW0LK
jeVWO1hbbjgBhizf4SNlJuvcvsIJj6XxKI/oNF8N8TiYMnYe5BoaEQrsynHVZHfQ
ERAzX6LrGUFvVp8zFJxjTenmmRVxbAjys+Z4Q9lfqLWJBLzz7T74Pj8mRjsIyjTc
1+sNmrRWwAKM8itT+UJ2tPGJ5uxoePb1nQunS9LpHope5BWkMvngRDpMWpzBv34D
7j1gcRe3LWCbvNnQhZYZozvehSXyRbrIvpYNb4x5HIet/wJ1GNvWlQezI039MH2J
WPzjLZD+j7lz2ocZML0x9WIwVJ7j7RbfVFmknsUzyJTNWWE8IhSU2XxFCRjn0d1M
sONljTkLc1v5apkUL+WJa7+Td0fgRQMjTnzom9KdKJPV9K4ack4CAHu98D4KYNu3
bhAH3vPnBJ83JBNJB1GcyCN0usbpBkbuZDuxY11YP8HjrQYPtpPp7z2rd/6txQaN
sM0AbNkId0hYMm2OHFArL4aQOCgHYL34j2BBVkhuPSAdperyrgZQFm64oNssbRnj
sH92hk2+3+TYpA9fLCUYsMkmPHGMLuuD4t8hvoHkApmh/zY4KldQf+fJr5nMyg4D
J/3hzUy0y9D2L8YtH39hEyNFS/pwlmj80/BPfW4bvdaqmxBibzk7Gjv4bkKdxxRD
0ukt7vFr3gCsgmWyxNAAGAahlIscgXj6kqbkQShjD0U7RF7Tu2XUuZJ45U4HzyCx
hk2FndZKemaXWh1/uN8TPAAF1TJt1fc8PTIxuMBoQXlVfgA+BhgyiehH37qG7AVQ
3HOuUbe3IS9FCiRD3QcTEvNR/9Y95dpAamkWeHi+9K39KA4tUaeovHUnsIU9vruI
esbV6xx7jBI5IpYorW7ikJUXwlG3cWWv1MN4NDJI4+WcY8xu+IEw9/kZw6/PnnBr
O6Wbjy118703qfnz+qSxSvRu3aaB9mIW/bM4+YUwiMZmlUjJq3OMK9G7kh+Nr4B/
Sa2r5vi9jA8JDyCsqEwVid8SwcBQsft+dULJ4YnciSvGH2xISnB82T43zC7QcA74
QZP5EUkrbDOYEGTcpxGs2kBbmUNzWSxvUHn8zNzSZ9koH/lE4T7aHJdP4xQYzRcZ
RKTJ66b/jDGhBTMbrjGVmnynd0SPEhHw4akh1mkTh2KDLS6EYf6malP4RvuLFMMn
eyyE4uKnHFT1OcShQ3EwK8wZYcLs7Wn2K69ikSCTXBcyJ2VD9t6kivfBL0NQhzAR
LlDt9wi1/KwlawI5oWRkDEEYUtLvAwUZIZdYtaWPlfT3RlzTwtfWv8pUsYQeWGtE
Mo2sK+cCxq0NrPI/5B9CfdtNsiAFfBCNbmCYCp8mLaG64Fm5OxxeJknx3Z+k1Kbz
xhaQSBHFuqUEPAfxR33euaDcv7ZcSrUwwX7ZW8dTeAa2NVOwHlAFJGCHI59WpZaN
8DftPv68znByksp0wqzTcGrsTuJxbuoLf0+7cQn9MV2XUPAa3EhMBreWhFT7kHAf
6Lwg6Wy/wefXnR+gS93S/JTA6TWk/vbgiEZBgUAoG1TmWJ9uS1vt1rkp24HymB7H
7JTYk/Sg17rdY6JXB+sz/XkiEcEBvcsra3kd0rUOTM6RZROTsIisIIfZGmVpyti5
qnZqsPhmXAtmSlvP35YATqFEXK93TDIRMk7InPcw8J8k6k22EoZy8pAkhBHtj2fW
LcNFg7OnmZVhhkKNftVA6d5tbkhnkzH9ZmS7JzSahUz+SJoCuGQeXlYwyjAisKQz
qxwVF7WXGPKRQaA2aYHgbwGQwp+myFVW0/Fu+9LKD6foV4umk03O5+yGDQYmPpHk
bGtg3vt452z8063iePhLsDhUcxE3J7q0UlbjJwuksM6x9kD+pxs6nJIC9/JKVhwk
gu+jLFBK3mmUwyIWkm4r6PRTMXUnte8S3m+ij4FXVDUgMjW78DsVjCuYgSuGmGWF
B9vRcroBq2R05PQOz12OksIG/0fbZQaAKOKkaaiY4cc6A3DKauOGoRIZaMgDkasz
JosnE7/EkFeFGauQiilScgn1XxKG3v0PStp9NSL6Fz5eIJ+3BCNVrhme5go7EV2e
aRDppcDhfZRzKqaMjMLVAqR8R0g/ewZ/yq7j3LJU+yF451PvWeB/cdteGhmj93UJ
XvsZMAAcuXOUxexPfnQJ8gz3oW+rgmkyDSB6kr8d4LV0PekVEKA2SeQwSXpLnYJ8
M0b7qyPVHyHkMPs0F4rXnjVDRSnY0AGCUy6LOEc9vQZ4kkbal0YWDYYZHwoSbw6N
26Rz3NDkFZ43+JJJ5wtxxisnaf2mpM3JyHD+E8vfM+K2vIvmDzO6fSfW1FwtXCLd
8xdPK3HPXdTnfnXjhHUi+p7gJDwMdMS9z9FTJLrhDxO4kw6YSgMmHgr0EdbFf9t0
UwUX9cwEeDzPs6LczHAnxSQwj/mvcT1VK8YNKMc2ZWPalVZMZIq4mvQQCq/Jj9qH
nOhpR8OijsnMSRLxzcejkR8BWE3sWe+H9FCrUjhErvfGxmgNt1YCpcrw0/9/7uHo
f+3Fk9o5l3MVS7qPNeIpa2knkhqQo5GreNXLtl30VAui1NSciVzi83w49d38xZQ4
sMSFCvNX/7djRZC+5741fym64oz9PNflVALWcXtLKsmG3+ha79Bi1CpReEL8xj6R
pzUNYgxnA+GCbP5sryUo9T6/flUIAnGJ3KxHXPmmUM7QvKrEFvMkADNlMl2ykRcY
MzEkDDQJ/fHRBrvmgU7e8nUJciE/UG4k/Mz2PvnqIWmFqADu2ouRc4VTAhOOnCM/
PqwkQwcFrrCmXm8brvUSRrhBvbTBup5FBZ9W5ez8Qdrt39cdQieyJAuYVJZ6fx2n
4dfMSH0KzXj3k1NG64abexk0L7AtMTYXiSAsVkPecSRY+NBKIpwjYq3jW0bOdmXi
31mjfEBegzrsgur3yyIFTsWpw/9au5wz4WBa7sLJ5nIWougJCAWSe2/b1UhzKWs/
WvHbF5mb0MZOt9CesdKhlKgPijax8gvtYmAq+3cq0Rhr05p0mUaU3+U2DxtL1Vhk
5oBwXCqQWTTxgmF5m4xKU4hyYcyX0TzuDKSBwgPzgDTTsmgzARZLTGn+LncLDtYP
BOK8e+ioDxtrpxMiMqHRRAfmeL3uFfj08gBjmkaTe1tMg7I7PDDvbONGcwKWDIyI
/uuXv1UKc3mmkzaYh9N+wDJi6XzYrL+JctZqmUcTOk8JPkOqpjxTOZ/EVk3mZqmH
aMcTHmyisIPlY5gb2ZTDGPA9uJ42j39HUxTqrOx1DvVQ6YyFtKuYpylf4ta/y5xJ
ek3fRM5hWr5qhQ78zKJAJE4sO3M6lRpLznILJpFzZQ6lmDEUSH1FXsN43U0X6NMX
ctqAQlnCgYyaIkJbvXX3PC0DJxGrGpm76uLHJz6MoKcvdIy6EUXBTpSH8+vRoU5g
D68r6ozhUucEweJ3UOc6QFipP0VEe6pn9vXAnESUjILeiKzAwcJgvxbRGjFBrEO0
8pX5Fifi3GF0qDiZreDeNkIvZvfr64Z9CDrmWZi9gOFsYA8qGNR/yEL160uK53BZ
lMc2IQXCpihmAlvFbW0kY+4PihQh/arDJHmTltRSqOZ5IRan+4GNM3PU8yPfe51U
fIoSnGlaW4gEn2N12nxFHH8dMZ1XkbOR9/6sgg2m4AwRDJRZYr4FXp/h1Q/Fffrm
iHICl9Dao1fEdS4nSWWqChq4EvbyDLvgS9EOKAzQng/18puA0FEjDO9tCap/WYku
wWf2pg2Dc0ogKlwBeeFp7apsx83O6OujZTRFWAzBCi3J9NmtEzAuCAc/+F7dfBl4
rU5jPN3JxKkN5EbDbYJ1RZ2Tzjk3e2iSULwMOLwyPShTQujjB2JpqrY0a/xRFtjf
agjxJaANP8kxTUf17Wy2lXzP+CBCLGDFD6zbm3Fzq9Npq5ig8QaAnQ/gU5b05Wt5
8olpLGn6Swt7i358IhMyPhxoE32BBAqGOAWBy3nL2HSRmYFtVlCfbiiYtqJ+B+y0
j8Mnzc5XlOXgZe6CDU0CmjfUG6Y91lf3HdVc8jGfwrjQ+RmyLBY/U8DmpGyLBLtX
rBExpvD06/j6Y3bM0Y9Wfn3JfSGnGHg34R64upMS+Jm/IISy/ElrH6Yd9770Zi1B
dPfIchHvHeOcSVb1e1Qexl27UIV1yozkAfdfE484/hxyHKu/cIiTqDTI2sUQcv5v
IFLcXUWlPWRHxqjMzrn96nMfApx2CH3ZViRbGwPYZnF6POsnctR20qzoU/GN0PWx
Hrw0JluN8LMEi0sYHPElda6uo8IGZfXsYS0uzfXWEXPVlzrvg1vZ+br/5gipFf39
ew8Pf9Rf9kMdffo35p6vtsKGthkSgwkOGdsNSsYRFJOj72jJjoMx60TBT5inIbqQ
qphwd9R2n3qRAT7Sp7kpXTzvA7k+1U9v5KoSjwMFJTbGa7K91VVpuaD/yPefyzL1
dvrhYhorp3lbBPm+mQUNi88tP+2a88HWRCECS8u5QnWMXaI+QxWTFFiA28eBmKDx
q6cV2emCbnPD8UjlN31Ajg7scgYGq3l+ieKHTc4slmBH3ahxXcyHaZfLBrXq/j4g
2yoQOM/W+QzYw6AW476c2RYfZpomFRXKfplqHGyJEgJuZpzRalBvLnjGPBxDHaFy
pNrjBFPlRfA7P0KtlerDxPD+hwdjsge4VXo6JRpDSBQ0xtpM+REL5UXUu20lPeXW
tEBaih94NDresiy43yH6qYZYgORP72Arh+qtcFr52y68yBi/DJM2HRFjtcs8y4pT
Wb+lsn2DXp5jQi0ZVv4Gq37pNUFNUaXmMA1RKSzPeLuHy8PNMf9akLj0qoPqkmHb
O5589fGORA3F5ATzg/CaweYwOVktR+WkS6TzeDT5dGAHzp18Kj1TlzWFhHxuHnRz
hVTUvqrSgSyhCNvrat3lmr1mwXoYsrk4V5TwPpkfYUJCw/HITpsRDVhwm1ZL4y37
lmK87UXAe+KAizRMjZt0cVI26+L6b09RnXfTJYIolLmd+VFiXj1P9oQz956AyY8e
xTPa0Obf9VUraEqTXS2B25Zc6gSCWXIJYreVDeyfVGYh5A6f6MSJadtiIhXI5VhF
y7LMgd4Q+Rgdw7gJDk7U5Sc/x8hCvVRErqNyXEjhK8jmtK3IIwxZbSDC+KfVTjyr
ACJtczsj0/BDk6srqGiHnrDB+oPQb3Z6M73LcxwjLVcoEphxwFUhqd20SL6m9SvH
2f3ZbWt/wAv+elROCYDThCLoJs5zVsOaxXjGrNf/KLfyFMsrygPOgeaZLkEbLS21
H38T5wuQc9WulGskvAYKRrLhWYa+nXCCPcvyepd6MonzHm7KIjnAAW94DSdnKfI2
17sa0gkpotqDn5+hsybc5clm//rCp+1gJn6T4dapkFsjwO6IfwPJcEjIWoUesKEL
63pO+ltH+iAyTlN0Cu9ltuGJrCCN0Kts4WcegJEEtbRULH6r1OKXMgVUB4EXe8AK
0V8MRj5BKR4J6mkn8lcJcjsq4Vh70b7ywf+C8wIh+eRq4BbnfjG2OqNWyrmnXoOl
emGJO6s/fQLAxUrR+FifnJcaL7zySvPIYbepzrxL9uxFj2U0qtW2ca9+6hx+R5iV
LA0DpLYHOHljOcLbxj4aWbbvuSZXCK47GsKgXx42w1MxMeLUYLjPsVIDhPkUIqjc
qD5QPbm78sAXuQmc/O8WLMlTnNROC0mHMt36BlduLMJrNDro+poOPXHel4HTLx14
gwahgWb6gyuonSjJgXsazx4EL4ODjdaVz+IFoSYxTEoXwY7kT4an03D+Jen0b+e6
dl/aPg8vnglf6LS4eTvuWjIhmjkCDJ7Sh2LHIX1her5p3ICKMKwmW2GyouXziLDf
L8Td9ZO8zijRdHBon0Cb2VPgFZ7+ASMLZ2+mgcfFUoM6r1q47wGjbajDO9uN4cNb
Y4hdb9O2vzOMyOA4F79GzYVunPpRh4ZGlh9eTNkgsQwgWb1iZ8eXsPqFr2Du5X13
2vagK++JbI5P1zE5tmbveepBMgmDHG5G42TV5OwsrO1CGCRwOph7FU+2Ym7+oFvX
UMiMRFaxPauOEthhQ+WkZ1m+b0GUi+K5dJe45riw7zXqoOER1RMFIxtlSi2SrNN8
sAMDcFEKWfM0TaAw4z8zX4sRt0IIxTl6poD8wpHGcQ7C5GhzYTMIe/x6ZOtv2UOc
kLAxuwaT/39dI0ByuxKs8XaJ4D0kRQt6JsNnzp0//u0+nQiTPtd3DjQlP3Xpc/LJ
SEVjUa8UhMNdqKqaZ4iByxDuv+SaHT4xS0NkNGxqi9G2Gn6Kp+ntqW08zQbScvHJ
MFOUXwMadl5EFdssSyD2FKrtoTxBPlPy/GNaUJ4ygyqlttUAHjlfXtx6XIe8oL9W
SEc96ikRUPBPZD7togPwsuwcdSEsXgA5Bebc2oFDZ1IR2syEbg89wadyc35b89K6
ld2mieCNtC4Lmato1QflfJu6fHxzZ9Px4vNInVSsmSS3T0R4xz3e72bOqRwEFCe7
aqmXrrsoJMNeIy0TuFRtC8P03I9KAFMB4nFx2ArjPmQt9xPp6N7wW1MurGevcZo2
tSfiz9JLW+UUr0ADY3QkdzUzoq+Jk9+QU/g2gKWBceAVBUfYyv78UvoU7k7Ff//P
irycgLjOMt+yEwix9axHIBYKuviSDh4hd92R3UdmR37+flzGGc6qtaNSzwDJaDBn
xM5EzluOY8sQy+LTCLhS6LBFGENJnIFud2kBKz/3K1LZF2cFmcZmxG8XswRYqNcV
G1WkWQiRj1EHtY6AMq0o83HkIxKsCu8cARad/n83Fcdh5/Xtieji3M8e++mrHJvF
vioFwvDhkJM9eeyq4ZI4QpVsnVgNnTajgRTKvKbTzZx2Zq07le8h1uMk//+dkBGC
pnmmP0fYHJva73BQ72kQH576A23AKfxg4NOqVBYap5aRv0oeyPWqmU0oIPp+6x2t
cC1szzcV55xywRZ1a42HIUZ2yn9XdEAlZPJjZUroFoqmp5314osznLVFZOvPsqrH
bXaHFNPllNLMmoM6m0dHvCe/ZFOCaD0LyNiCH+hEalOhiqzvX7bRqiDP1OWMRRRD
zYUcSYpMJl0PIyK2RedkqCJWpeL++Ne7Tt5Q/RALnMjgFbM8Ge89mFw1jgip+26p
LK9BnWDNVJRlD0wP0qwl9UrNd6nak58D3kv6aZMzFJ+eEbX7Kr1SrSHR+yy0Pqt+
oygiyroG6E8D0yyKY6QnVYW7/YI6jVKCLPm2F8f8son4TOvnWpPa95l7TAhsv+e0
j4E2wWTkqk0/UH1revbVx39Yq+50Xlh3CSoJgxKz7alJVAx2zhdYr2h8lbJPRsS/
NTiiSYBAWcj2cugCeodgAMPcHmz0Bc+7dbgvj4kuJuCbcLxD/MKZP39mphxCJac0
1L+IESmOfCNOT+uB+o6DcFKIdkBRe8a7hvLVv6cN7YaccewU5y71jnxQF6iHaeWt
vDw5aYYWdndV+WJEGlXbD50iYSWw7NB0kvaq0d5qlp7wipUQFndKLu2i9wSbod0o
To6TL8yUubYbxg4uyGS2ZJRjivZP3/lwGw0Q9KEb1MQx35zeaoLeRonREcVl6RPf
+neJgFXfv8sXfyMEPTHM4dqZRmlAEUuPvtp+EutnoOlJ3j55P005h84VvGGKkE7o
jP+0mPmS417nlZiP0u44QmbkK1vkv0SSpNrX8RcfRRSUOfL4emBXxOOpokJH9cZ6
Cmywokfq0c14mLz2b7xDG//HEBLEe0VQKJTzLM4T/AyBpi4JTIO7O3XIUpgvhDnr
340oXB2O/PlGiDHNT6TM2vuQFHoLp8jstwCnR2XBljzBk7UcUgeHN+sxEncFNvKh
QCjscoPyqLyYJU/wbd/UsX9SXGkcgxFtT3IouB3aFof8JDN6qQzX2aRvFiMuZDXL
/bLVI1uUejbW7mw15JXkmHpgzAB9CeoXLKQcKXiBw5Bz5q+Lo3AUOgPKfPbEK3LO
Fs477pD7R4LHL+SxUmiBQzlWEorDUaaif8aSVcz4RllfXwUneXnNuEw4OsVNt0I/
WAA0WUM9hgJTj7jWk56+FZhXUJ+yITFNXY72aRGgSmWD4Cfzb0P23dSyNCVYU9vv
bSFLbq8x9dipYzakJCWUjOHxAUcPTbTBGUYlW1DWpcMFmmQU9OFzrPc2Ed9dWUlX
WMKtOqYvjSdOas7sk7Z+5tB8zBdiPVyTQEJhHmCzjLbMzgEVVgpFipO469+rcwxt
mutLnM4757FZ/lhotnzob5jY1c0YDyC5MR9zo7lMs7mjH698MRop6Nn84KF58YCF
1nNr7148o0Gqagcr9uoT8A5yedIsi/8uFiC8R38gxkd4dhrsAgXZTKtPr8QuRXkD
qY8/xBpAh/1B17ePBhy9hpZnse04gLfs9OBuOB7ZZLSdVjKICkxeu2ayzgfIXuAe
Fa7RtJWYPUYCnPnCKN0ntg/zrC0daNRbcwqiHvht4/nOj6SEn7gruTcEB887DYFq
xakOzQxiyJfgJtN6SPUv8d1yi0tyyHzjPWVdwXJYoSXX1b/MKeaiyFrf3LCwNnoY
B6oXWJ29hXjjDKLyVp1Lj3ci2LXfoS2P7A4OlhJyAtkqP+xi9Gzgq/KeYe9Hboo0
amajoc+zJ+fpAlRiLl4ttdEzM9J1+s6qMuoTkmDDEtF7KuN9Zd4VAmRLBLIUWw/Q
+0Ms7Uy+mk6vHxAiTEkaThFv6Kd8lPQtJZpjOEEfmJk/45eOTpqFdCvZfxRs/r93
sccGLx+qdPgajgx1aIUJ2G9gYJCM3THgnclnIC17u7vBmFSthIcL+tqAvQUB1412
v6+uO6KCuLQYYHF2mtycg6MmW0F1Dcxj7GhGPzYSotE66Lv92T/ApyT2xdsVsy9U
zBddc2/yvzJ4/rjWnafxthgctbuHQm7R5lVTb/4QXkhgG9oIF2zfhUiwCNVZ/EjF
joadYA9VpD62M2Dvy+L7XffdlGtmXiCNLehYKjI4WkdRnQrcGqeVBj3AX4KBweri
TZwsGm6F7u2C9iMMQkZFGiBArMqMHAkTdiG3SSID1L5vbDZRLldFou+ZsLnS1bNk
NnKXl8IiGR5HQ+8sN9bagTZPmeacDl4XwoZldGDEQgGQJMEmLDSv7C8cKmpNjbLS
ESWirUcNXjtqDt5yEKXnUp1slq8qM6ae0PlUY1GXMnw5ysadmb/oFQKwe/Cwjwcu
XNQNvXm/DMsue0egfl0NUoSsXhbJqfq8wbP4gt9MyMDnxQbOCQU4yMKsTNkS/pWd
cxyhq8X8q4qWgecIx+S5qa5jCNQFLf9rl4H9NHu60WVOd4PeLfZwxZqwwi/9ZKHV
bNQgAlVNqfPHnXNICAM/L/M9uEPCa9g954I0RKhtMO9Yyg3U7uWQHD3hfjRKpgOv
adLikFXhkt67sQjU+5ITMXEdyO+5cfseHn21D8qLlpcIdFP65/ZirQqATAk6FCAp
5Uses7jI6kdO3bvoQDXkMVo2VD9ykamJnoXedbHjMzfStXhYHHad3+AtBdyf9Obg
t1S2SBsPN7Y19KcN06AHm7ik+l7h1cB1C7ce5JG32mkBcg5/Ctn9laJ1vx9d4rpA
4mN+RV0iKk3o+xdK+um9ANOMsJRk9Mokf/Z1e/YdKfggxVx612EH3nDN/D1h/w+e
SbUOt8uErGh1LT90e5dc0gqSgBeu8+R6pn3zbKHf9WBi91sHNjvn61O2Y613NbLD
uYGLcNMRo6LINoVB7JD925XQXMIDRy7uczkX+4kmig5gFGs9QTRFWKGQIGjYFNap
SlYeFbfQH2qeEZwIiNQqy70Gh5dJVwKy3SqsIKWMwHg78pJFHt5IcJOwb+e95dso
8Rc7p5nTz5Z0WjlX5HDcOlJKhWgYkAFdQ6kNvs9ApLfvE0cTo5H8IIpZBRsor7Cw
s3fQkFY0leD0M0fO5w3L53dGaL7e2Yls5kwmtyrIMA2Z+noIYAaToEQarAnv1Mo1
3OM3dcrTZFa1s4ChwdipmXt3nlZarMhvRIBRbR/zIVz/CgSVWvZ0UGc2s2HA91L5
H3ir/wvDzhA+kjkABTnDqaPmRgecnvEsmxlzz2oDSOJVB5I+F+HywfsBcT+hPBuR
Cw9yqNeegD7jZydjZFa2eAgjSad74XBC6DOkO4jKU6Kp8YzoAS2qfKqyNkvlvpzH
dozpGzKdDYGQvv1Xg1TruHILT8Fy71kGa8wVI6TA+8rJCW/SicE7FYg1vZ79f1fA
EjS9GoOyN4QbGNn611+P/frFpIbOvWFggy5zAAJToHzelFral73shQy1r/e9yE/L
I9MVJgP5LuqP4jlVyqImwaCHNWZzBn9vr/c1CT7k2I58VG33SGnd1mSnn9ET50s0
KRJJ6YYBt3jt+PzCnC+ln/+jvhRzshcgiS0NFHsdBKhakY5k3HiQr3+yAcGEXhx/
bVLonNEJNISzfJxYeETeTXQpIGNEOMWdcZbSeVXYn5lM+xOrTOrMV9zT7aZ6CBdF
LF+JEIPLu5GRVSO9gw97iuJ8MeUAwYfwz+WEuJr9fgn5FzkVaqdxX4INu0M9SI+I
7l8XTEuxI4asfzxO40I50fwb/XvvZXKZywjKTWw6zcm79vNxVX85P0oIyq4Rd9eW
jCvSRf/dZTglxaBFa7PiZH78kxG1tXs3eXcAihEbJpXtgL6mgEoUv3xW++EOUiY7
rzUyqg0eaViGvYW3IAZpz/6nvaXI+kbJN+uinEu3lr4Bt8uXqhemnEpef5td+EYI
cZuUJW6kx56Fe2v7nhjc304sp2FEXrUOAD1j7XJNgE8alSRWhseb54a3Om57qNY0
tV6W5fhmgzQzd0dz1RA8Qm4H01cGwpRrxZSr2gyGq3UOEmAaJKNWY1G5p7ZOlqi5
b7EOQFsy3R6Ri0+lslmU3Pcoma3uWkYKJNLmTjzJ3+siRPDGkemIXEHqEXIEllxb
g6AnKByU/Kzp3YkHtSt29QLWFwgqbZcslCWP1VG+PjszqlFLzKUNsNnYGINixASQ
XYprO4V0YvHv1C6NcQCR84Zx6wXTULLV7eCERDKwX9QtkSWg7wEj7izcigSUEIQ8
jZQVW/pxRPme7jqIBf+nni4hVHEEsLj/8nWtKfuNKJr7ZyrqhozAacwebhC1849j
v2noS+tPx/J4b07H8jLvkeASppwrNzEc0TIlJFnSXoHJNn/aoRvFFdAsKid09V4T
fn5u1IvS0LGHlw5vUIIwnZ+/2zFjmbdz3TlcdKvqb14fSk33K0RPUL3qDfAj9qUO
lI8/4lqvBgEWLHs9xMsx7DDpk4FCG0SmvF0qrCX3sJQ8kUiP6XEJwRDYJ9nk8QD5
4NdVKN5VL1xKHPrJJT9B+LvY3EQ+uqBYv+5jhh6IZfWHCsG+G8As4iMrL8/pzPBZ
HYwzW0iVlCHre29DRBHt9qCbXjg8ESz+2Wk/riUQ2SlrAJWnscbO5cxJlGyfhamV
jBPbdpJGoh2kM1u6WNRtM3t1zT2ePJmV2sJOeQCx1jNPn4dbexuZGLUwoitzpDdL
h3qBCw6V2SoMP2QYWWL4RFM2v1ylXMmk+rMiY2IRmUL0qR1ggV3KTG/KYDaUtyqy
a0uqPPDVZ4Cttk1idtUMD5E62y6u1WhzF4naMWccQZnStbL3w17/t5dKVkxo+/vL
efTr8Y1RFz7wtmAYmRA4JZ7g3XDf5/NmAhk1/vPo2jsv3AE+QZGUCiUaOSHGX7kE
YOHLYefeKB6XKWAO/FI0LUCZCBFNyo2L++EVO3lRCqelZW1C3bKvm50GT5bljjia
mo85vTjbVIMXm1coVhJE11efoVwZxDUstj2WoW9aawsAITB0n0XzNggYemlPT587
iHU7SvAfXFe9sG5FAnTNlatnTEinX0Cs4cXwTbJJzN2GztQJoFkdU9eAWuITE4GE
jd2XchdMdwOD5U62Ver5L0kibrb/Q8QADSBghgV04vPhXlEw5S7M/L+hJtQBJa3q
UpF0XHv62b7eBpSFtnnxZumlcjk2bvNvZaA6TJOwgnwhb/Z34j9FUW7T9rEzw1F2
jQiMZI4iedpFZPF6ys+aHPirdmNS81/pPQc0/4x+MkWJAYwa08KzmvaLDPv5d/mT
oC/OEO09U+AefdkNAvaYqzeFrF0sFr9GG1w0NvQsxFmRU8yWI7X7HPED0ejf7l+g
ARgazNk9WFw3Mc4XKQXFNnOfCS+u8Wo0Ieg8+qNX0Oq2KjHgRYxs5S9DbIWp8Z4z
8AKpL43lWz/u3gtqcoJODraiolhKlY3CtWJDDIdClHVD5JA/3iiv4Qz0VCiM23NP
/qyGFmnHowCAJuvM+txv612JZmglIZBGxfCcjjHYdH9No4rHDWOjRLfkIyYwAJss
L0DEonXunS9ITHS0ULLlLZVy3dnfimAFyGAP3NlH/okYSfrHi3oxKAFvCz+1drTz
A/gSXU8a1Y1kA7TmWlNelqsCUHofiLMiMNd3/KvMJN1JC8CQcLiMcVvf0vPAkE6W
L1KFzhRjnDvEkKCXcRGxx5XKV131uNJ8mvDnJ2XQt0ak5F0tIaBNiFmxMqA+kmhW
MjqZidRviSwsLB6Z00qBOjxfcnEDKoLZlnipS3YBtX7JC4iFblb1O3nAk1FlJA6u
VMUTjZNkMJYttvkVrsiczX4loN2yFk1n9y1HwnStRdOEp1GvcZIlJ7e6CgKBkJKI
OhZVXHszWuhK3nyUAD3S4kcJHL1/XrTjz7fRul3KuR4Btb8b+UFXGF2lWQCyxaWe
PzqzSKKy7LETZTXqat+fSc240wsv6aB96uf447lLEtXA5IzVdxw1+mEWnOCYDrrQ
0mrjq2bkKsrGrlT2n+jdHRZZCuhYfEAleabP4ePhreXtoVjTDBV6vde7aEjNCZPX
DEQuSnJe8U0qKBzO5WV6dMRhuOlZ2r7kyz+z3/1YymG+wkNlYHeIyviHAYXFC8Gr
5Nh3pIT6nd/CmXWnq+zA8mKlTgZnV64SGI4Nkuw3umnBtCg4sXfQMZ3zsnzmzREN
nNs1X97J8uu7zr7sjbc9hod4P2gJ9u1b5JAfA6QYdAJZJSuRf1R/JwQ51NUUdBVF
4yLn+C2twRobx02BIBTSyUdbunDaVRx0A4Y9iJamfPuBXzEY26ynMLRCK9LH7Ffz
sRLT6RjmObGGoR/cjeiB439R6+4Zbd5XpycPu6OrlzlnHtIvbUdUTYMKvLw9wHnd
nVJ8KXcyoQvsWeplXhFRnpz4EpuIP4C82BaHsuX/4QXaGJWvBja/vqg6k1Va2iG3
j51tD6AbIa1tjuo7crWy/WSqz/ugc2UUIe1J9ou/eqklV+AVzMZNRbf5DI2EmCuD
66L1lEzSEQPaqgpvBT7DjjMHBqZIauqWH562wfv+YcwrvBhMFZyS1mLLQ9pYtjbN
wswl5fo3iBzixbQy3o/mgwaNhswJJZKJvOOkVQBbu6ikB9cGpUpUzFeUkm7+9hT1
zb1wapvJS7nY8c6i/0qlwe+jpEaR1fFEPMuKhqp9IuUWDnvMca59EecAe5WsaCcU
XgbNneJUvi/6XLlC64JdLTctRIUZ/Dup+LYSnIWBiKb4qeq64mEpUATjJCaIyOlc
g89Kj0L3TNRtZgiqBXipG/PkuRiRz6ph82WYDPOGAuRTshCANDnB+OkgB4ZIeIPp
qsMIE9IyKyJG+uI6RTdpw/arFWSpLJkdLDsN3XzSXsJV8htOgjV+zwVal7t5y3Dp
KYEypNir9E07BHq82QX/dCkv7ZFCHPh1AORlDEeK6ddAjqTf4UHIKLfFJOmI9FPb
Aq8Ek0Ka29YjjLaFSGR8Vi+Dd4DLQe+FZiFVPRHgXWMW9gaNzuz7rbg0TThvwIsg
CZQMyMjBzsvKAY4006G0hJ6tTLAyyNU+BwZkwjl0C2DpPH0CRk6Y4IBmzcoDiXYi
miqKgEyqbOqd9JsnWyF8R0mVG2BkV6AumBY0Gs6l/kneyUpJsNK5al2qk3cFyUY2
EHz0Lx2skowsn1br7hSr1C8eGTQRlG4N/fMIfx0Yb4CKZ438swqOT6+KOq9x0qO2
f3jeCZzMQDRhdnfs93ZF47zWqGCHJB2XVGARZ8WP5pd+4d7TDwGDfPBrowhZ88n8
1SWEPc4QwTu/sJDkH1e6ESlZ7MXb6eEMVwsBbFU9Pxyw6IorIWYX6Oyl95pyRLHm
X2n4PH0dsruzPzOW7rQpiJI6VUpJDfv47iNrry+EKNzcYfAUXZZzhDxYcLmgV1b0
JmmvUA+1+fCk99NXAvevEswQtumHNppBJa5hXhl7noMjbyBlUDBj67PJkrRi4Yll
UNKRPhusGAWT5qIhXsevDyyfIxCAr4Ldhf8SlnC+qxW6QuGwBLu20UEhUp0xa+Vx
TdiXgHW2JEalv9l0K6vTq+y35qWmSZb1UbmM10JxqQ0JsDlDuKI2GTfNadWqmuYj
8LapGUW83/c1Et+2CMRqEXmmiIDJ/x9nulsvKTFi5/ehbWlH+AobgPmCYeZjpvvK
U8QyZl0rVIqwf/FjOt0+HxVAxqCKZhGSMGNH1RPzs2872Tlfn/vCI4Df4by6TaxJ
AmhPHE5J6YQiaysn/pDYnZTrao+KpI7d6crs+r7s8wDwrE9bIltMeBreiQ2hWoLO
Hcxglnzpp8NGnU1a4uQJL7xj1kGa0Ko/fq9PcfeeYzuY+tJOQ0TK0POLbeAzXYh2
EzzSQxrJQ92QjMu3QEEgcMWdT7v8Tg8knUeeSBzlgNw/59L0Mu3KMMBYPqsgTVEz
MHSfqFnnoMgTjjDcZSDRwM8ii/uIvGwKDAJicIZIHtU+pWjbu1mvLY0p4vAg5Yjs
cbypikof/ftr1+cumVAuhjdWw70spBgYeIGw4sB5Q+fQyR3b2mmKMJ2p42amZmDa
9iZiEi8TC0zgmZBx1/2cRcZW8T0jP02zSHVIB/YsfVjj97cgmcI6L0lAE57nYpfC
HQ3XJlazHwkWqkj7luLIBYrCAFtbB04HlOUp+s7NvfeZsq27CMRzPC0penTyF0+c
rQKLTVRhjt4kevirwHkuCBn+blR0OMP/heVRIKwrRp7Wa7HIseQsSZJIExbZ2OwH
KXUyMgesIvVtJ5XeJAoPlXTLr+w/3yEzq6SqygHGP3vPlVIfev3hxZ9wHfO8SEiR
gJ7NhesUiSDS5raeVdzqYwlBfrsTaLEwnU2jwht9hGMUx+QFjNd8O47rDyE+SW5O
RC6K1CyNQ9hQRG+d2cdM1guWArmK8jKg+iev6DaL10n7wSndgg7bJYrRhwagICSH
jW/CutMzhYsQC4NXnr960aEJHmY/LgMGsJByFIZnT+i42HMl2f3YsjFvm8FgGWtI
Faz0JXoJ29goz6YIWnXKy1sjcBNtxB/l7wCJrEC8Yd3AsP0W3rbAix61tDGZc17p
kZnVffengmkhPXHMFkiwmKS9mIjVVcI+9Bac9n0dSvlGSEBKeQ3ODVfbgpN2iBPb
XoSPcusYbO2+k4rDvN36Lhr5B4Aygdt2JjOctQ8I9yKslHNZgByFTu0xUZqSPM0W
ctVJCcuc+h9bmW+VbZY3/TwjriaKEzbD+M6E9Am3CQxtOl3cXeYWNgnMw6+P0GrC
HRiD4P5UZ8Dx1IwH6E5BTIiivDEQX8PhCtWLTvlPsdjVQuezK09CCYR/Cpyi88ps
d1dph7jsHxl2aEjigzqukeHKxPN9uguky7GeLtkUFSw09y4TBbJBpQNKVPT/y9Jo
PejRqwbgUeNes6rI9PUnRQHXdwog073aWSILlM5AmVtDQix0LbSQLY3Sw8KV28Sb
DGr65Xzspin5vsZqc2CK9kOG+/ndlaIbATid4KUJQI7CQVr454Mqi/cdfAKrsLzS
FifVM4f71ewWyHvOXquiwJ0WSg8fFltFLjGZJja9U+5HLRGhIfm0f0AeV1P3hiQ8
xmB0GH8iiaHKo8Q/0nQAzpHG+pgTHzi9Dsgtac1EFEuavuTxParM2ghpdlibirq/
Je3L5JKZOvSZuuhYOxEjSepwT3wAo4omxK5S6+W47Kaky7QTaVU3lNDyRrb/6JY2
UkkiJEEy/YRLywZ5ASMLJrNu2GQoqD8LjV31q0BwN1Thr7rqMSvJ1RfT78knE+uK
hqigVrUGvXmROFDwAwEpaizQ0Hw5RPrn6j3q1TjxpfK5QICTRNJ7eFnRSj8k0EN1
iP0Qdw2I7OjZ7tunQ9/LbkGv9ic6XCjBYASl0MzH3ckIlxvIuRvfYfqeLmPZqDDv
3O9gCXz/EcboZSNPdRX7avZgDaP8gOCvCJyZctA5FknHwehI8xkfDLNrYOJEluRH
Ph2vUKVVROixAeSGQLM9g0doiinu+NkVpE0yJ+K63+Uq+b+ShLsjmdJ0Q/OFPTS4
Hm3CHDP0cHEEBd9VZBRc69FB7DHaNG0NZYYmuK7oTs6rxsPyVz8FldnTj4QsS0/d
+P0emB9SdDnCdBZCMYqAIrDX4+LJgjKDbLio/+PSuPEHxN30PlfomARQltEqRLtT
qEJwvO5qixmfktn0eLg+1+oZjeECV2GUrBz6+arCPjAI9PqJXbY9cSs2oqpifci+
fnGNQr6IBOxHcMPU//Kn4m2DlDH0xyybkvxS5KsVUqXhCo1t0xiTQT02jROp3Te7
FGgSZF3gMwr34y6KI1EMLHXKct3taEYGhmWlzi3AOi1dtqr8JcBe5wyot/X2SijG
bKx7O77OiG9SWC4ST2fVgvVxoigTHPesKVcQY/Z0Nu28V+wmlTVOzUclf4f3l5df
Qnz/bl0HGx4fsqwbjON8Wsql75ffZPmo8JGUoSLHDMW6Vifiz8Prl0Ra/KV2vLqy
/7dwcRK7L4GQxH5AlCjM+SLBBd1jEpx/NaJHP3bxTbfG4FwJZkJFVnAlr/v90zxK
6ZuHIlrx8TWiWc5p7yXscvbfKvUS+7P/x8hnYsTTOU+0q/hYTlz31Kn3t60D1NNW
mx+vvqpeuT6P9BKyH2kOVaP4GK3BwiVJ6Ch9Ze+hbOsFnw/26Q33ovihxmbXIAZq
yg0QXsJwfHk1XoRcFrFDB1K+DqVqnTluT7DxZWdrFoFch3AKHB1aLlQ5HtHZnSjT
EgQ5PT/lCLV1H9JRfJnDRxmZYlcAhG+Jv4+jT3EURFzn5NefTBuZIlzJjeB3ejkE
K8wSFnocy/b1JfJJLs0MbeEIWBZgeghMUDk7HOut9F8Qnq1TxEQXeuDpSE7hNp8O
RfT8yiaCpfOJCkW5oQMfOqTwZeQGFEQm6saPVEZefRQH+ciSWGrYTIHJB85ZrPV3
g1EvmKPV1dzCL28pcfZd6oyMB7LtaM1ij4XOrMDnbTIKUbcayUWwO5qG6HZXG6mi
lbf0Xn6sGtvkltkbpiV5ZoEcARM9s+kXW/AxnzOLmz9T2qWeh4ZoZ16w7y/PznRH
FalO43/McWTOA1sWuAUmCzTzjL3e+8RWJSAcTCb51uMrY1I/Kz53MXXm5JDP13ra
cqkmW3jyVk+gueYPZ3qc1/Goxbk1KZLr/tWwRkrN3KDu5GhRwiXxlRbRaul3FfSc
avcvMcpN/n0E9kIXOMOVzPK0IXzgR4jukq3Ay9Qnmmfp1+lA4mOcBa9kRGyiv3OD
Vj4Kvu6jRoD8NhcghyUHtO0TPEyplX+U1/yz7llbCfYu57HPAJ/9G2FrpJdPxuX/
3yKOC6LbIUg83v9tZpDU7pKAQpTbIMmwFfHgpt9siBbjTrHFknSZq1v9g78y/rCP
8bidtJ5/jDlK/ezwPmzS+SC1Lpmf2YuMjr513lTkw1lXcJZWYZ2TWwPWzNK8ZL0u
SeTqOXuceWoC6hkFJvOtDET/yiIkC0eVUNp4Hz5GaX7bBfw/Yf+ZN/ImmbZlF426
7676i8JbkXm5l0FPLoi4wEsZyzoUmft8pviPFKI6Zd97nwR+FdaGHJHaN2pHc41i
h5o+PUC7I76IMeCNANOuDlFyTBzfPa3Hiocq0k59+fQTqIfnEkMmiuW0jmRl9095
17yrvx/frySe1Owy3Cqh0tcFqCzyAXIUwtyYdQlcUhLeo1IIL3Hdz8cicOBd0oXf
qA3G4WBygwEXNJ4gT0Fu8SNn7ESVRcONesEN7GL+6KqsbENUCXgyJiE4m0a0+Kqg
lLOqjT/K2AYAb0Y8koGyc7BgmTCWRu+KwtMrR4H3HpJ1QGjAntcRmdLdx775Loi7
uvY3NTbhYdmd/anoryOZ+QCn/d/SNEDLR16Z+FyhKMVuWm4q2dajD9jtUxXOgSCr
XG13rQlesqBRfXsXhEsDV4wCE6Jzm5EaX5qA8CTG1vWuxZ01wJCx/f7d3ur6Jq4l
SlwxSXBlZqHMQhHd6DLcbUlVN91r8LxLjbAmgjqGrmSEqwc5aWIUsBNebrPuzz89
lgqamRyvDYhBNe97EfubG2yu9lIgeWo3zmHPkh1JayUHFCW0NUphR1lKkLXj3X1u
+19FkQqDcG7iHE3WgVnJWzun3op5XBMce1cY0fFqbwc9UaPLtvNchMFT2MeaQNKz
5h8cLsvOZ9RUiWbUZFdBhhu4zGRI1PiZPGKRZhE93utxzIWE3EHasXNoqSQLkCmo
PK7hm11s9BjNezHyTVVuUre1NhLnCXL473gxcNqsHu3xJ827ydyrIo72jzJTaEpZ
57Vh503QoP0QBwtm4f0Bct1EEmbLeJNcdp00SeCWg8QE2BulG1jnd9gXf+MIfah8
EYyvtZVfA3JHS1MCfgNYJ2/RhTv/oxJ7ymRK+ElcS2La2K4jwexk3B8/XUEL2x5c
Qhn+e936I/JF2O/amR8SXxQzPHBt69mv4zoNV8UF6HkfZ/54m/M6+5un6mTkhYDN
OumeLaPfvbqdW7+unFA+Lmgmoepv8o5hmrvCJXiQe38tP3DUx9yLBiAKRW2MZ1u0
GONPm3sqLEvXxcAmPbdRHySGxdHAOvYsmqBFjWa8qsWPi3Gb6JZar8YaiGsx7ATE
BZ4Rx6p57Im+3zVhSIyuOKnosBYdn9IqRfPgNLec05iq94ImTAFvxiAMlRLJlTSo
fSISi/g3zytyfjVOKXoZbDDV3xpT8IXF13prCsV9FnD6T76CXkVkriEPw7uc5E2a
5h5IX8pyH/BWyE4ooyhfxosTrBlDdjaIpZg9BLMqWfpDvIeaMyCeghFtfy6P5hLJ
M1TFfFs4Ggcauuhb4O5Jn8rOMhHLFVuK7n+FkNiMwe+SJd5MaTvJPw4fFxBT0OeO
Q2gyK8YLSnh4DAHHKHqBJGgsUAFHbN+e7dC5cl36xbPanKGiB8gXPIfFPfarEl72
bpeNFEMVydR8Z5IDoBH3SbyqfXyGplBRCjS52lMeneZblI5GMGVhropGS2KU9N0f
dLAeOFtV1vAHnwt9Y7CjCfcH8E5NekjdTWsSNZBg0NFfS89IWM1Ei5+CMlEkl/wY
LVf3T5Bh3aXuBjaRR6l+xeRH8xaXfvrpTIsoxFKulqUqqYzFHGd8fWR75hSAZq2T
mcQV3zwmT6BTDPrWgvv/O4uax+3fpbmhVJkkv+SS65TtfAXBNdcRS/y0cV8YkbND
nFJV7GVJRqp7iDhI8NyvlaiCcG2YuyO8NX7eietfogujdmVTxUiv3fCuxVYxN9DI
PANZPHjfbjDOox0q0wL4Vz02tMaaKjDuqmpDMGKvPhFY8LiPUlcK7TvRLakoxSe7
bJ6dCfwMKUzMLvxASnCa2AV5yE3+RweyiFxv2ZP7ZtLfVA0UtNl31k63B3FDSNiR
2/lJG58rCswMV8AI5iUws/pQbDJA803djQdLe/E49hxwVC2byj40UzWH3WCr5Po6
rHiDUf7CxAW6jG1U3eHqDFEIGeEM0ecVlC7UT60miSd5Ndvj42aNOCl5jXA9eYdz
TD1TyMvaN899PxhJIkugKj5JgJ1w0YrsDry9a7IPvdYCH5AGoMN7M9jr0KXQHgGc
YQA7VeQSdJ5Vq8qAbe3fBIFxlLedwdv+iOQ/3iQhoP+/La8EsoTJbCVHYA303Qh5
J7nGAg12wHBofSxW1mfqTTb0R4UrCPrOAnGqZykLZNdg1u9qZ9xYhza4wH3mKEuj
0+97tMOS4tpbVxLmYsuLNj3M1b/5kF7ds1NEQ+QuTYiJY0edYUOYxV+vZslyCcJd
ND/EwKAFZ8W8z4+5naykaGM6bgduE19zbdH0dbd3qWi30WfIn7wXbHJgOJDeyVKX
7hFPKxvRG/pEASHRPKmtj8F3gvPe070Yh6tAp3TRihv8NSAz0kuAKG/ISO6cRygv
/ajTj47tEDD3CFa6rZnWocPmL8xW2ZCrz1L4xuEd8rudD0e+WImGPS5a80iqRviH
3ZJsG/5TBT5gqDBmruLdzJQkrAr3iMpK5+/ne8wVB0vSc/6+i1CYgHa7kKu8gGiQ
Norzw0MfuWZyzqGjQw++nEjcGvkFMfFJ6VKdukx31yY7I7HoTp8kHXwg396ojXFA
PKR6CDIf3kbvBayGk/10zbEIm4LdHfCdBVfVcTYVC1AA6/JaJF96FMRmRLnYg8sg
aRPpvJm/suqjiubqt3JSYJSQ88K3+OQ1bhKBcS38TndvrQSMxQPnugMlSARynapM
IXk0a+J5jrs/QbKhcmBerGuOj5gEEw7fcPs+LH0jtJY5IrrHwmR/A/KgPoUCyBVK
7hwUEuuzbOyu01yGWU6vx/P82Hwkaa19LgTawuX/rMPl1JENgc/l1APGMYSyh+gm
WMUtNH/7YMVUyqDdpGvbuL3+j5MwmykNFgRSMxVxx9I+Z9GTrWOC4/vYjdvUSfWA
LC0orDWF2kjXEFitu4kF7EnU9ivWAwpwqlqZziqYw6+fF3KaPWGcQtUW4muRVYUE
Fn87bSnj8qVnUwedT4vD9tBULzg20wEVZCw0TG2HNVqh4Xf0seiyJGNEMZCuk96g
5x+SpScSgU588VRJ7v7gdwyeCdA508NoQtp4Hp4u5dGtZcbwKtCpvhP0jrZWQtRu
MseVMWLYHWXXfxcyAflvx1lkr+XqqzVBG8EynrNh38A6SMtSlVkI+v9OtiD0N2ir
4SB340wyccBURRWSjAWagbB2E6T408AikC8rTwy6Ix+1p4ErTS0oq+QW5wy9GRWs
VhO4SJ0MiANh5+bVDi8NJAGG+p/2FG3fWDRxYfAZmjqo2+GR8swZGnNoGcL+Hral
vGTVYn1pCPotAQwyNxn2tldzi3SkLdHUSBE/ttBqEfuhl9Z7KDH/2p89O3Bcazn7
O9OjjHWMfmeTuRnrOUf2ZmRcwxs/meY1LFdGHc8+2PCcj+sBrZEmK4mv/pOdhpi3
zaU1FWS3vlZW4l7Srgs3PpI0pum7yGlf8NF9FwtuyjCVZfoeKCBDdrMyVHJvymt6
rrQ1Kcy3qPAOV0VelL5F5Ck5FugrVdoBg51Xmq/9E3H7u6wU9eavRWqvbbid5J2j
4nLF5mhGWoeRIvVRmt48oRdqYWIGniSxy4PV5NDLewdWz1NNvC6XVoT2ARXWUF/6
DNCyEIeYDNLs32V8Or71mY1BsWAXhvFxFOdqtb+8Ikoqc6m01NbaN2hY3FswTkvt
koGLLTqQe1xRQuUmCT5WyiZuVfdBFUxWxa25WUF7kLchEAAlsxZ8xzR0ouKedx0L
591qwI+EEOeqxkvl799ccdjb8pH7hdahVpwHI1ivjs8OrGdaD9EjOO90ZD/ta+8n
kHsAWbwju8rrbC9ig3JGsRdGjIxpvRxjbbiKjkFePRvA1XwOuoYdJpBrQ43zIQh2
R/lB3TxP8l9ttRdjOmu4jEAxTpbUc/HZBpWOUCXc6kD1ej47PUzUCAYnd5BF5BXP
Ws0l9c0ceu9ihoefYepG5qwUIFS6wdqEXUFIWZKdus2QlySCQ5GX04xJpcwArwKp
p/jHcvmWkvmPxLjNUyHmz8SiwIjFrKUd2pX62noVyHfO/AK4vy1RYEqku0fg9OD2
vRRDJpOEnPJ1K5xlvgJlkUjqzkGhPuA15621JpsoMAcZCwAPhWOUoNDvhVg3G+sC
0dg6uzcyuWG3AJ+qBCE4yW2Mrr3CYRnVCa/gT8MvoVDWJz46ha3dESXN+9NAg8zb
mV8aTznA8glgSiGn24n+ey+gjh84Of2Q14Z+kLUcWe30/qihwTyoyNOE+POQxoQJ
yTbF/HIZYjKiYKzgE5hgkm3XNaYxt54wE/l6X+9S5tMfrmDK+Yygf5arYbkiL6zD
1Ws8utMkHVuZA+DesBl+wCg7gIDz8lEfmSGuAjtGQrgv/+fergeQ5VB9X0gtB6l8
AMFKs1xa1UVhnevUkqcr7EzyTnIZCLoaxn4I9pqgPW8z9lmbpSenKBFYy9e7cjmi
pK6ztfNOgYKAkLUqvOuqd1yYeldBzZgczCK2S1I1FUg0nW79Ou5OrJnq/dRTNmE5
g3F914S9NCI9W34hWPQcFdjvTxLeociJPrdBRp/JEGpwasSJK2HegZYUjyzzZjm1
SqgUUZoTijL4bRQVNPe1klTlKzaftO6hT0gGcUREYllMBZFuw1rkEa/jkDr8pful
riWoh5isABAYoHtLU/qNsIXAnXh/tUmonhibwCzwj1JCQDCzfK85euFLNSCMaApW
RM4W7eQC/9xaHIjx+UAJbdPC+ted07NKSPCRT6OOzmmZiNQ+0MyRuYL9n0sp3Fkz
T6XLLjB8SMEu7sgcViq6mLFeGQkx3RTK2fDPhHYKxIvwqSaR7q4gwmLD0+Bpg9WT
zwbmYYgOF/fKuqxgUujlTUhngBo16bwIW9udPzB0kBe0jxVwxIOSv1yjJIqFyQRL
Ptfhru88FGeoioEczDvEG/bsNjYXr/UI+aAKbn/w+9sPm5ukkbT9WDYsd27v3b0a
LIAZI+MnqPO4ibv0SIOYuh6SOE6h1rxTVvHs9BWHttH8P+P8Cf3JOpdUcfWhvYXm
uk69PuCAPgOJHFSUygUbfAnOzYhbU40pcgwfAtLn2Q2v/ElEiT0bZXC8FXHPZhLH
8+jEo/vpSFvbQgwC1IoockhvcsqHF7/TuiVFIKZdsNLta+beVn/8ev0foe5y1O+F
/u34pL80bSjNsXXnRbotAEz1/1WLXcxNidL7mgrjitfMVhnFwr5Mb0XTEc0mPv8D
YMoCbpBLB8kN0NKTZtEzaYGXAb1ziuSuDifu9wctX5i7Zc+V57xrjibap+O3FFO5
TOso1s2rgSNdr9iYxSOwyjsnmkUgToW56ZpbvN+IgJOPgN7SGI35RCQa49ilM8k/
4VuC7soFrMtkMhiLAETV93D0x7eS8YbpZcRIETsZU5SpVgIFWnsWOUEqfbTBkMCW
8/7xz5VO00oOgDrgpVIeOFNe1NuQLXjfPQND6uii9Xv32orSuldHCAGNJPzRCRzx
PaDXpR97eqaF4ZEykmmgqZzqOh5izfEtb8A99qV9DNolY4zb3mjZ4sK8wg5ZiSmK
nVVQMNuN+6DQ72falw/1xTD2/cGNzZk7Gnnayvef/dVB+iw/HKw3lv+6CDuTqgXi
Keb2Zj2Mzo8artmIfd4B4E9vsWpTN4epCg/HvqrRYW1Qq9SqBQioKVZ+da+TB8Kh
TOql6xFIat0ea3XS29MS7x0bJ9PLW3s2j3X3B8dhlzVk4Mr03G7U7cyhDY2TR59T
R7kaTm6Lh+ux69Os+ESiGFd9lotn5OLuU+z3uuzrTmbs4YTjDi0ANviUrGmJRYLf
+ssc9pdcFbUxI9WSlgIUDbjRBc2EnKd8l9Y6Xt3F3LMYqgjsj/cI9awurugD22w5
yAHv3SUlKvlw3eUyxk6O+moxMsGkouotCIlIu630j4ykvwIMpXLf4cp6eeLw00M8
7fYLuqhdSwyZjXiFO1fG6e1HReFC/OCvwXNFyCYGhULN5c0ejMr/jPJGHCLP/i4O
0FaKNBCeyv+Uu5/ifY8jWh4AFN28/HSA+8kWIkeVEYemDg/YzBjHy1NEuru0LrpI
MtTxLPGTHNJSxOjEyDS+uFtaHF6vQtRIXvVJf6fASoqzNOBd7gS5+Do8tecwvYBj
QpCQ6mwQGD+KSjCM8b8BehYYY3pYxumLwd/HxUkmtRWKBCXQ0m6j/ySH7/xX/cwl
Sk+J3EZYXRR5iv572c1sOWrZgkPHqNc2mADDdQO/rUzB4P6Mm7lsRNuQPq+hW6oK
QLCRIN3z3w4AtPtCY+qPptG+/AxhxZzYnqseXLzEqTDMk2NzUBYQsCSZXGT0WOTM
hoWAE2ZBQtjsBj8cQaMsuamObHDqOWVc/gt/cDMJX0framNQvgwAu4kKNlS9lh1J
63/AmwiH9tAjVHW4vOP/6+sIWQ8K4HWXOT1XQRZ4Sh63KEDOr2+mmwgXh6UPNK/M
PebFkvLu/Ih8+vB6TO37pIWH5FXkQX84rfkhf0ogn/83xc7cHL5I2wnyjKWBhw9F
OEyXPBSmtZaaQwauyA9juksy3Rk791ep0jXH3EswNEB1GndWiFiPs8QC3P6AZSoh
notlnLK5hF9QaDv8G09S0jip+fBnVfTtjVUG1zKQUpTcpBFh24e8u1mX5TCzkVIb
vOo0W5hZvUezQQ4MKjz4hIgTM/zWDPz6j6T2VpSvUT73vqQ3tqr8FTIe7F9a7iKr
7vQDk4Y6HopsxAyKvvT8FPYMKYcovdKbHrmgY+7XGEdPaqDR5eyPOEKnRZ6xySW3
bwkHdcZ/U4E9GUsPufMgkP3xNgXzTkByg8bt6FGPDKNTR9HdWH9BoF1rSMmt7pfS
AmpVqFPgIS2tMMXv+u4I31X3vktrexc4su/riqMMUQn2Iuu0DQF59Gi3ZFXRrhWP
MofHCIkSR+k/g5kdhz2cK4GniOD0bJVmKXNfBob4YGMcDxIA3X4nNM6MpnucXtuH
0rrzoCr43AXlptpt1hF4DJATsxAkoXYH5Ylbw32D8iB59nqux+MvMjhuIulL9/6C
7xFODpjuOMfI2hmYWM8wydfrNGZe1ma2tQV/ZL7MYsMbazJ5Ot0e6cDyD9cxCtBH
EVI5PuvySJW0uwVM2yEXhrcIo7l02NJeJ5hMaJj4trfSUTGkz2pOPC5JU5avvzQB
arj8wPrTFTB4zEAvXPvBrVr3+a8bzJqUvvqRy0ycl5tu4nD5ppW88qfC6+5+iY1z
3ljlDTPy+grpv3jlOJHeeDRB2xROdOKjNSRQsTNZYvID5ONaaiRNCtLyIl7Q7VOx
1f1wcs1gYBpoFOINnOMc1FkoX+Od7zGdBYb/jWGfwH2KUxvH9Sm5mAhSq6PDlAjK
FSLI0rVSzc1EJ9GJcez1Q1TULYrItiJ/KIaRGvLnhDDLpIUfy9I/2aKBvKcUEEjp
mA8AlI3E0oDb3i4CNGO5V7OxK+s4BRpEwEe+L8Hw4f986F+tDO/bcyE8kUY3znrW
SpWGycjAY/SSffGCoAmyc4ZUF4uQ4BXZ6wpNnloFzjTis/2cZ9LXUhNSfrR2eHtM
CitU9I+euNeelgNZ+oydFJoFbFXu+niPoxi6/FZ3l9tXLUpc6eP/fSLxp3bh/x9q
xd406vi/U6FlUfM4NcuufC3DUgs5h3s0ZM3taPmvFHybmy87nEaXcTgFOXxEHd7f
CUUOtQ3G3JeHzgS7dvQhyVqLUzFSR+5Ku3UYez8WF6KCOrag/2VTmF3znUkQMzBt
WTgKOQaWuX6aZRSACSHQv7V+E0TUpDgGrERe4F5bBBvA1S0NVtXwqKoy9RSxVk4i
AoP4s+MX0MsdOOXq+BXiosckK3JKcAn6t/Gne1kVrwqoElzwVVmApIlxsa60Q9pk
IukW1WPRWEX+th34VSbGMk36n9nEL5sol+2glDeW6zdrn7/bC+/J/IGmoV9gHfIB
XLjDYSj/MzZrg0/qazF7X5eh0X48x5cAcIIBfUtaloQC5/YTMRxOmZoNm0rpnwd6
IkO96NVLnJve9RWvFoNtU/THRL75ZOI+Ts0J1aPRHs8gafO1t1hWuUeLBucJHSU7
+p1qYmQR9is+8565rQhSDm5X0lV/hcjs+lV/hCoB7DFADZvo8QZGugNSi3cVkOLi
67wwpVahfxrqcPZKTaOV7ckBknnCFhGz5hAp7ibio55rrdvqMDHOsHw9KA4rQLBO
6kSpOUcPcBtk3FsKO7zTczgsUckqK4CEhO+aAddjhATV/IzHGbvCrJbALyqZ5tec
zQzTCjNQ456CP24nPTP/6xN1wnPwPhDSUeb4/nsiK38wMR6uvr5i70KDvJQeQAKF
ZsPoBPPUL581l3y5+4RSsPVjk4+Wtl7qQNcsp1yvbEzQTsCtqa13aE6o6ELEtH9n
29tZr81HgTFeDgkszIzyZH/d+BrdtvUXo7iuMoJB8gneyaHFqlxt+uBL1VgFzKrv
G4jKMgkX3Nd8F78N6QZMzvhQSymFWmrSAF64WFGestSKTzKedVPUcxko6UCrAZH8
D9rsJt/V8Cgya4Z73xsqZGvj3Olp8D5H8kblUDadZELQj4uJVwiReJrYx869A/qP
i3x/RaLksG6OWLV0JNNv9kylyTZTRJptRJ4l6GK4G+kifZpOZ4sdSohaRMRaVMzj
fQIxpa5J7gW5ZnuNG8xqsyMlX5XQKtmsB5Fcx27El3wa1wH8pz5YAH95J8IAI8I1
4RpJUq0mKkXcAVkQpQZB5pRtpNNZ2cC4uOeuODSeF2pB0617p4oc6TG6hfCYrWlJ
u9psuvWeH2nwT57xGYzV0aJZ72Uc/Dr+3LhIXpZtvdQmRdy+nkUSft8I06rCcjvz
PIfkL+uwInHfBlATjUSnjaoMOx0n6gXCNA/nV/PAyLL+NptcGomCPx6ZAKniZ8L4
rRl09SL0MscsspZr45eaXGAeHsAYx/KEvYiP42YAEL2knibyr/xEEC3ubQFdjNrJ
wt0IZe3wBMHLuNmqVI073I4fSh+QnIlHd6gId+nI61+rqjQkZxyFNTQ/UyAg5A7g
S0m9pr1B47zzDOSKGrZxJ8aEvtHei5OYxYM450RgzsTD0i8c5ZeG0qKldWrPd9AP
fSo9JYImyGj+UbCwMXZOCpLSUq91L5dQRcvp8jOrTrcwC5yOLumBak2KnlOlOywe
+tjArLY4+d7OWeXU5/gfbs2AWzxRU+PdWLmSXuZGJ4v5OXhnCoToUt+xdkUZ/cLR
j6OidnQk0EfEdNSzYmkGoMir0TGz685cDIsICpOqev4qTFLWqQ7p6ZE8bN0P3C8Y
aN0u4J49EvZMwyaidykdJYHkhByoVKoMHC/9VGl1fsdTWIHAXDvtJeMJVbTAvToL
8dl5PxWWt1OoDilkHZo0q7jErqsgE6iR1EWGvnB/oanQgiJ55qyTWLgxzML/DVL7
hXxbXFz/3YL2e9ZaeCzwIupDej9OuiIq1chlV2WRslsR6fsJ8ccvssJm+m/pINYi
6u5bvUVOyd6X0fzQTGvJ7NXz8GVViHZbVJHGMWX62mgFl5btESxTgyV/PAKDdqp4
6gSPjJse7dpxVlVXv5L2TBnisgenPexvUrrsV/LtX1RlSdyKRTcaS+heOseNdran
XC9hPXKYboKoT2tmng3EiqmOFWmwmQKVSBiryWVBsgUazWF5lTdEiCAnji9xVf0I
LUveL7a8g9876sdGf6IBmFsL944DtxW6daomuVSvLijjLgBmcFIqY/4zmCqZLaft
jnV6xGIu6eRiS9hHfEsoK2GWAkjNNhiffDZI6SwVYS178B5EwwNAurCQGurax7Af
LeNQezf9Iyy5j9tN3+kn2IuwWigkzsWkC+GsmSlmgF9n0bZyrZ+boc5MM6EplW5f
4bCjArWDqwHpw3ArBnr1Ldo0WS2IPuX+KAO2eAZ1Ex95/du9snl45neTZCwJ3n7I
6UzY4GGUnaWcVCZqRO/4BsSNsyqRoukONP9JANQtQkE7TWg/jf/viX5ADWJgABEP
Y3wpjQcY9CwrSgSGF1xto7XHTaWWiMzVtNblk1tycKZ7Ni1EyVnq7utVi9rz+lqd
qMQW2tcDGvTqrH22WEnYVfMkhTKxs9b5ZybHhLjZIkcRSkniFKYCG5Ja3AUWqvnZ
XKXH+bfT3xDpTDnM3KK438rgyIM3gT6Ax4baByUoGwillZh7aDaeC7xEYOApTzR9
oVqDfnRNiStD+gCaWrCCfgzgGhmgXbGcn1oCcM4h9OP/zxwfUoyN6R/zLIhRz3cL
7dmObyWSZmmqqs4ux7pFQWAOTNibScD0giwfJ/L+ir8ytyAiRuVpxqO91NTZiKwD
BU6UZz44RDvwj1dflEcroNk+krn09Gk/kEKeRYI78kTevh2jn2CjE1+kRXmFJqiy
jOFkEthz40e/LBrBqmZ+H1oHHvJkLE4MKoCSXz1jWvkWbaIueYp3B+4gsy826GWU
1ynt/QBvP6zupBEVNdtk+QvwBxDH8W15c36LsN844GuO1+kxwcgznK864MWnLotu
6psi3eHvaK8DXxZyQRb8djWUvq47Vcg83xuEcJKhVZwxf8N6JrhzRERMRIO9dicL
Cu6CJlgyVyFmDX7ZmI8OscrzWiMRMdyzYsuc1zuUn/ZuFfxTTWN5P6gsZEkY8LfE
xTkEhw+FyMkFmZ6otuywTxuym/KP4sn7FhHx7fP0al2tRAr4iEAQzN0xbaUxXGCQ
UZSXiE3s+yCvHkrpW9tlnFqK67bAIyutFbYWey884Ea6fSexEcakGTViELiAcKhx
aCfzeDIrsNfxqP7fK2SqDvOXN+Ul0eAAKnacqHJcYZnsJMry8jepP2WFlnjfBkCS
UlxsilpvnPiEBhVHqfvJYWRydZn3Yz5ZXNc5bEYAJN9nGkJyXS6oIu5GfI5V4vTF
KmurRxH/cHVVPqNKly0tqtLODUYIpBKfkKmCUDEsW2RHN8ziRiGkD8S9Nj9sm7zz
k0FeZAF2J9WDUhU7o61vUWjpqFdm/DZhJ9/MXi/7TK/qDsqpNB2BeiVMZIfx5jSJ
QuEh/P2igFlon2g2UVGuawEspd3E7XY4/Xe7Qm/tNQZT43kUYwebFSizot8NR6Bk
CB0hVYoBpmkBWWQBkhDhcFzMVRU2iB4JVIeP1eeJdrK3kIle7WrYLbVScl60PpRG
TsHDxs5k8weSAgjzqYsUxU+lPDqXSR5Vaw+hTrmDqNwT1OZNoLyU43dmMz7BbUYU
0lbUoqbjW5F/2yNEdfzwDau85peniMkJPtcTAHQlDMUbG01GjX3CxGx2lLq9qRH4
a8yxxsAV716hOK/nlZ8/NHHeBdPaEYyJIcF49rUlEhI+C+3EwOiW2d9Fq9z/eDfY
zpxnR8MixjPHPh0I6O4I3MaH8aiqdJVnma6YWvmziXTK51/0rySX3dUNZ1r3NLb+
iMddyk10YxlMI/cSVwrsZBN0ejcyNNQXZN0ujnUEGTmSqJ9CybRVW4FqibZ7k8vU
J7/zn9lic9tN08Lbz3l05L3FclyZuAHRhPg3jpr2JzsuEiqCKcIpv9KQk/2Ld7RR
CSAAnz1YmIetuRalHataVSVBJPmUekoJi/EG9sUnsc1dpNq0MWGZ756KufLlSPbC
EJif5ioAkyjNusfaDrzaf9+89ePL3F4RfyDcME5Sem62Fp+qPtZCoGp2eM5l7nSa
xULd4I5Vhe+vSs2OoTcIp/FhXc6ELTdTRmvyodgmCGL0/vFHnhJ6RApLYTogx9Rk
OKz+4Zn+LZ9+fmD4NDfS1CZLVka966MPvpnJg5jAhJ8cQ3lm99xg35FHB/G0YzAw
KMqeM/SgfbzPwomphYkWb64nopfRy8kEv4yZQ14Rco+NBI6tCGrxCeEKCPEjPs/C
iznd1JQUkcUfXrgrUn0ybMwMcuskLlqykLqPNWlAwxl/ar3idO8LaKsz3Lu9k5oD
4W0AMFpTxjDlA3/+VvolT3nPjyhpMDZyedu69GxIjFyrmnNYUHsWqc/VIjdyn/31
ec1pr9bP2gz9sfdMttbdo7cfJOouDw7R8fGb+kYu9oaCb+zUle8TR8bDG1vFHjTb
NU7JfLX/3FN0PX1WQLz0kQCLmbjxq5m0j5+NrBSZmI8GAzthtHWhFjAf8vuQka4q
/gi77tbrcC/16sqT6v7yq1uLkv6gXViuP73Log+r+UzKPCuIWILZ5Ua7LHvBeEsn
80EIq3C+Kqh19b7CUEbbKQPUq9kJYPqJOzrwIhJAa1ubYfXiGhd8sYhX9hjF9aZP
KmnGwrZT5UqRVN+dJlIJ2brdaUjJg/mCMm08a7Zp0lbxa48Aj6+2S7LO0TIZGIA1
0/ykaG5BhvDA0AB+xCR5+XWtd8EMWlppQPynDG4gn7SaxSEy4WgdKIkaBMVmb7MU
4dLatz78r0cUQ0SEoIbTHznpd7bpajA+mV/o1cAjVF0yGlpOEV4XysN5Ikco18rd
a9LucoevOFlAHXKAWKs/t0FlEvD/YWJXI5pm3yNsqnuRJIFPixjWF1TZgGDQAjJI
/ulXEoeLkHUBCQQTs+ddvh9q5Ia4oVmxvKd8KK6XgJNIhETLvok3qaLT0nXwZ43W
GTzzUpe/tE/85pngerNgrlPxQ+1DnXrYKlwope33Lblvv5FmhemlUbN8oTAfBI4U
Y75uazqq8Hr5/zjaEUOFHwG3+xl4yVr0UeWc8yr2jxZjVywQ3tS1dPac+UC9/hTR
HA4SCPodlZ6Fxk5jJPcRUgO797SgrUk/HBpeQLdFCKd1zFIEFK6OJp8GWk1USdYO
yhOUJtnwCNoQZPz+YQyv/1NlSu/loore1NC7MPYoMsP+m8f532wYJCPsOx6YTF9u
4pfnjH76GWRxQZWBgolXY7K6kzmocLAhDV8xEFga3ResK/7GgcQ0hWD8RF9V/XAj
uQ4xwG5o6SnoZwVoj1wJd1hdBgOZA4Md1fOH6GFwulCgPJruERm/hqe0R8508gQt
P9A9ymhUcxAaPpfVgfWZ7AesHzeqVd2pm4ibVJmMubwx0K0gV9lVa65hOLNpgQJ3
QQ/1yKmVeiVyMwRuweGlCGQeifHXuFiMOZ30ONQbAfo1LNUnA1fyL6pfAC9/axbA
E0aknn2Q7TzHeAqhe79HHFdaqzGiMF67WODlQyGBcN0GHWALaA9ApkCYH9F5FxZm
h786+HA+Sabys6Nbr4kcFiVkTZrZmWDCuO1L5rTbNsibDCbDuot1mgBOdW62dy9/
S2OInntdWqKMgiIFGS/K3AnznCgTANcEWCzEfHlCedmNPWIL/u+C3M28S+vHFvXP
Sb1PDEGS2KtMdVumACtPL4f8hmvTsygSA7CRPmrkErnTC4ekfrtEbJDyanNdtuth
1yqlsBoj1/e45ehSN+xlhgtFOsiUs0rSJuF+WFW/H3586bs6X6/65y9mr7HjpVbO
3CMJI2pFCGWHdsqx+HOwjxi37wVMlcU4Qo1u77DnDASrdD37+lnFJk1txHUM6TiL
ejQi+JfUIvYgU9c3iZLkJ0EyyCuZFwm7LzjdK/8bxtEXrxDJtWqnodMYb6NHRDzb
3tq6btmq93/FwKdEaY31bk2urjcowdqyZMRmeZNzrU6FiIPDxKLw64WGoryCwDNT
cGLdXeLXfywZxYp4DiqWdBVUb09yo/e8CzMEhaGupeNN1ei/lXPOQ67M1BTsXnsY
T/YRpDH7W9UzsmzFUNX2WUJfWy6EfswsG3V+Jlu9meg8FGT8yQEEewQ7YdvCkI/K
PVYDdz/WWekBbnQKLOSxXTQ0m/BiiKF1jPAznUVIDBMqnOrRNMM/wz0UyxMjiWJZ
dmfVImFxCX2eNJei8BQX5ZUrzHldvzh0tRDy0RXPQ9Z0EBFDlJTBE/4DU+aGqNKT
Cd/ffFPmRPgB4GvdlHcvoPn5ssu8Z7ThNEEuS5+RhkI7Lka+MB9chsUD3vG9gt91
u/rt7z83KC64PbSHgLmTU+GvJhI2WAC5hSD1LO0BP7HDcBWjTRbLT5ixseWp1kbi
T8QXYvyTvDosId9nFCdqKjkj7aJtCx4fYWOBkgxqpbqacXKGkNcUMaKf5oJ8+rbh
6JaMW9nZoy35u9Ob4g5ZPYj38f1nNvYNHI0I5LCBPA5lQs9+/xCPRawG1s61u02+
Vy//C8KHT7PadVPnAaCd8WTs+9VLOg0YeJVnWgaDKMza2d/0FApuPMuRZgvQn+r1
0IOerEoX507paqo5t0ArYee/K8x8MP2RMf/OEjnS37yLLM1VS76836w8q4zVlO3C
ZvkN/UJZyouIaCMDBnv2DPxY59QYtysHttXjycQMMZS/yaSuJ6RcSRlYl8S8ZIBe
jfCLmDCFXc3dStqEvZAbaQIsaBGbIB97JgX2e2vymF/7LRlFkZgG3muV8m5QhHGh
A5W4AVu48Z28yDvvveH7cAajCqI3fPcNiDzd7KOSlbgzw58SC1tKackYf3q9PDrb
+iFjlx4HOzXCSLJIPaRFVRrpCSHkEAJcRXHqouFHUykMOK/rihk9/Fv5ogRuH5SP
utW0ATZRIP4o0tBAzzwAtjdGvdtA1cL/i8deDbludIPWhUo7s1p+M9sKZasMnqIz
MpHCil7FSo/3cQRO3ExP8dxTvB7RydV8MzVGdS4PklwaiO2ojYu8p3Wdh0FKqycM
5IDQ3TscyfuxQEHRbzCgFb/mZFZWglNLE1sI91fsVLfi2nFaaP+N3xga9H2UAhls
CLIFRLdZcbzbOWH6F7vu5wvJVXCm1ci+5FhMaJ/MxI36Z38fHbuYagAlfVY8vk/n
CR+Kwq9AclCrhYDl8yUfLU/WfNQI9g7QhSXXEue3xNreymzopa+PSagHxsEp5GDQ
NzGIJqaJn2ypoTOgoKfc4PaGZaWqm0CNMA+VoZyvGyoLTTfT1XY6pVE22w4KKx2r
nA6SgiM362yrBWPskSrkf7oit02+FR5TpDHXZVMM7zVM2l0WIOrte9dFPx/eNShw
NTkM83+5Nj3JX2rTx7uNAJZRpdcfeQFGRwwHWOFDwXjyAdL99ZxYeKmylAajKTr2
yqinRdY/B0Rm1/6ITdDkRJEo4Psf/dbQKxEYYJcEMxGNuUn6Y0plGT7Ke2AAwfIl
z9F8ua3qWtHXnzlp6MyHozh8nnqWH3V2tvItqmJFG4FcNb0lydZudVDF63JdXvCT
X3pO351PBGH8+TbB/AGKURa5nVTVlIlLXtQi7LMPA0PEDTesQxldU9tI8nxLaAkW
bQDje0Elw/VyKs2ByULFV7FdmUGLSXtVaDZzoeXRdcFtDEU9sgtWQLpacBFNt/OE
r3z7l1guiItfuI5s9k/nS2yw3ARnnCOBD3yEVlzPTmBrEJyjCI4pVq7l6CQ50KD2
heRLGytD67cpS7myX1rc/SbEbLamhXxoz/68CBbsJWeUyCDoIzPRaOs5GLTFwOto
cuLHWyxYicLuiwB38OS4xsh4Px2hdCrftenfFgciODm8EezX23mRaz2R08+E1OWe
pjiSclGtmGFytV5mSXNE6+H3fGnELzjnmbc8+p1nU6+3QMHP3azLWSXxzaofz2NB
PYZSY0xzhrLCYGSi8BWWyso8T8GgR7nn573OKDIQmCDsh+LcRO2uuW46kqLEk5Fw
i0KpNinKEqcFQ8cRl7paX+suB7e+AC9rgnDVg8iWYrYP0HHh63mWD+LnOZNYmrK/
LiRIVMuWpzT1K1B2DaptwP+NztJ1QKpE+4TrOOsjJaU8X2z6d28LZ7lIpaftxB0G
/AeQP58IxX//TWAA5ZsrKxn4d8Ft13qq/sVL/HvOOvSKPzS8/I0SF+cPiww2kpca
RIoxuGLGSjMC4YzzpJ6mnwZfmyXNrF45uzLnH9aYj7D1j6U06KeBD76YNUj7/hl8
5HtjxcDse/HQgikJe0elkVCKSe4aMrffH0bpW8xMUmzEK7xf68+gYSNdMhfnVJEd
cv8MDYGbXuMyXpRCVnLtxgnZtkd89GfdLwkYGGrZGhPHfQkQWzFEw4VMOGOjZp2x
bf+Dl4NVe37FLz7JGgu5ud+AhmFnDb7hwj1uRhNr3JaCeE3ZmTwDTOQfgB5ihNq8
n14SVdqGtx/OlzqBl9E27B1Ep8rz39UdYPB4iyLNVAK6pLEeCQ3CJk0fDsBhqaMS
X8oIK/pkn2in9n7zilRdc1dPsE4yeHUw2W8YPS41EGnXkqFXyX0c9mLwEw4UJmDJ
zZ8UmazedI8yWtX+/RaogoMuTeFXfWnDgQ8T8br2OdNKF+wgfbmFFKk1sxfEzK8N
gdJmAnZqCXEvcBxg3vKTntvdGCufxez8N28C0NrgtVnw8FAN4gpE2upwUCcgfigd
zdAOxqohitf15foO6JjvdvMxS9aW11VS2QLGTHZyDGUx+6TQpfI0rS8HanhQIwty
eaGNSgKIty7EMPoEu/ApuuNnXQqdtu8z8mZqgOAmDUiNH189ZP/8dq1pLQQTrA19
Vgi1lc4qV25ezQGT4/lz7zMnBmGx7KzWxthkHVIXz83K44LbWwm1z9U+ur1a6GA4
O4RMe7+wz0RXaNZqTm9Zfsh3ygNUXS2s7mkXCzoj2As7u90HnJx6/Xubrtfunxq5
sUbtDC2LFTsNuoW9sy328AS0aQYRoNuwXaFFmmYjVB9cKO297GLSU/KXzssbeOD8
mtHtEMhL3ed5B8tcyQkBkSNRAaQPsn405HeoTboQifEvddclriADudJDEBNHs3hz
9CDfbiP9th2ODJXp9aNkFyKh8ZxqJqn35AMElvDHTiGEbEbCffTn7/suOVpKaFul
NHyEVEMjfZopXvuPdBTjcBS2HBJhkIZWRJ/yEozwwFkOtbg5FjJVeRTwjkcmoDCr
tWFf0CSQFIRlqy3XkhwRyts+aJIL9vW0L7mWsqQMVTlKN2r2bvxkacpob8aDsqjG
JMMIw8TxZAS1+VJlHJFfncLU5Lm89hklMZ62xWCUTSFKvBNP9lIhzts3bxKD/Ll7
WhJLHHmJMw2a+nfnDdpqiDysSyaw+yMDOuMCKmtLrdqU8T72CFfsbGQmvZc43iun
nX+8V4/Bl3G2sRcdaiKKwdLg9/x0GhOWshusCwPu2z0UuONxvfLi4pATRxBQim6S
Mv2iBLaI9ynapFufPZm939sm8KPBuEkb6Qu9bqBfXdZPmYGj6UhBe8TNRB9AS/gG
bBrUsD8WZE1dI58ONKfzq7AOzMQksXW+D/JTVBVcJpp+6rujOhJP54xzXE1KfilG
2cXoXngOyXQl/347rIrFOstuZKi/UL2Pwzm/e1nL6CpPIatTGAtVlv1/gJkUc50X
EqvHqlxKmhEVtEGdqnDpSGJmjbbh7YJVpyfCuAVQNA7pAEO0dV1ymbPq/z1hvUiE
f4zQB62kFpU6wZv9rVN6J06iZHaEEQDalVx+RROCXbAdXgkcMjMtD1klTsAUVScP
nLmhVudludwRtQHKQ7yolDtD/ko/ogFkjL+mbTUbHRTI1RijxsHaYd5Iat/t23tN
3WnYusZ7Qtk01io23NXZkN/5QMw5nwGGlOmq6Ro4/Ojn8GdRLFQfOnB7dPguG8LK
mVfu/GLYO/BavCEndKVw0pL9KgkTi1GWra6arpzRsUqAb7klUsx6kSkAkXZordpu
cZqWcE1x5+6cIxMO9hZpNUz8/6DmoyoEMrZ1sonco8gguqFzZ+eQRnrG9LrsuZei
TkHq9dLXU0q0y8tpstiDyTtFziwW7Jh3py9JAO5AFtLTY+v/mLjdZxQSKkpATiok
TbWMH819wekXtMe3LkX7bwe8H28GlkQOP+Kc5dFWft/ucqmI6s5Z/yKhjlZ9a6Sd
4cWG7RLqI39Ju4A3cirvD9KsbN/WWSHnoBU5ihzfouzBBkzfGY3xMaQgfgqWbxWG
qcMRQIeRFUMzI0/8H9x1R0/zeZSw7EnsD9mEXR3tq/lwqo/x4Kw+xEYOZIOESui+
yIolLtNKIFRLIMe0IR5rtbxKqaXY77153twR7Ck/z6fHI9RpG2pZAXyti71aUTo2
MY/B6RiOluxjkdOx1q0C8gRoFTPRgNGYT6NybRdx0ZdQ7dzuKHj+jOz28eg0YEDd
aaKmuI03DYGKvrh28dtofqqlPA/9wLV5HzxOLOhbc7EK/GqdCPCud6kVAnEXPWe+
vKB9xPOUWdz2L8DBhU1Th7fGTZppDum3z/eXYTab7H/9mFmZArYYlo1PnvqbedsN
X/43tc9AY8bkR++7ZW6xQ6gtTjJ24VVGsgXls9Vlad6cz2o7RvlphRAQvA0RYmXa
W73MTLWA6yMgoOXGSS7V6VuHYJ/zzUxg0Wuqky6Sk1/Ol5qKMys7MJO6doQJeCzu
xzUPPhnWVO63+OzPBlAywnAoZE2YpfoHnG2QtitonFyXMSDnEIBGIsY2F0MD+SpV
LcJ8+cV7mKNG0Eld/8QOt3sEZJJVqwUraFBoyLsI4QKHd+WoydvEddwODvJRyw3h
zuiDW4UnOz44UFyMePilN9V23wKIe+eU0kbv4NscBHdLApIHM2+0PlfdKZnwjMBP
jSnH46Gmoans2Vr2LkihYMT08aMXZOJ+jnJnBIuMkbB+OPXbRC/n1EjXv4pZTQkS
w8StAK6jxC0qwkVh85cUOGdIz6vRugF7/c+Lxq0+c0I8gZz/RJcCAkV6X0Mn+sg6
Q/fsSvWuJtWnJHwrO/Em4tAnYF58pO9/E8SYdQQYzQlPD0PzlJfpqPOeB6QPUDlb
D98fXjWFtPIWfLW0dT51BDQwkoI69if9XZHCq591wdl9ciDROvM0tOYsfvKl8Tmq
lw6/Hk7uNVbHiTyFgbc6v+7HAkb0aQhpxLugS40OtnHJzR4upwoWGPX6wEcGqItp
1+NMDdKqGAZw2JH0lXVkgmJjfZqEOTjMVbUyD15xpXcbk5+VAvCjNXy+bKUctxKF
79cv2P76JrqJHMoVyUfFQVssGzFeXQR0xg+sNhuRCf+002wjhMwoRzSi2Q5p38j5
xR2qUJeX3bb/cV22Z7V9Pol7EhWZ92b2J+brh/aqLhHqvsBpZVVhByPUJ7MhDXjS
OgK4WQ79gcVEoBb9p/saApUhq1F+BgMQGczqm9oEWsGUVS/Z+elQ0dbaAVqS9KHr
49UpRKmeN0O/q5VGu5yIrOHP2c4ZOgC2WmZ94Z0dATEVjB1FVNHpCPX75da5kaBK
WiXe+ZNGRU2J9X5dpAqj0PACwsbMOGUtzNWx5yu/xLlypuTlIKzeQs9OsZFWFmEp
NlyDH8eZMGR9FfPoOiHUcOMJ3/lCWS/Dsfaz1G3CBfLKKcvlbl2HhXKumEGVvQHG
iEbzLfHNKimUpL1rJdEJNNl4v8f4rG4jI+Wg6TLRZtDfbJ8BUp3GZeLOjyArOvqV
jIsTWlmMEWIFp4U6ClDfmGCNsaALNzLrDHD6daP2NOSuE1iElmIkvhJ8MwOmGGOH
4qwu+qQ4Ud8gksJZEPMOcG345DA4sOVTAOoz+xQUuaKx6GyytJfbdH0dUwEU3B9y
MhBWpVtlBknw9yDcVmkh8Y/RPDW8hgokgWYVGOIiynpt/BFSmDq8BhVZuawta0Gq
1AMwnRQBS1PgnpFWNtaTyVGGeNB49tq4DUJS+EejaQ7nmhIsUxGgFVj/0AN10xEm
7dGZoD/TXZKjFHyfNsbgb1iC2jDvYYpaqy9ZK/qEbg1BCkNEam/hbdDM8EsPST6A
95yCyAxKCan//BATDcyqtSkBl+7RFQT87wcQRVmm9HlKjKSLbctmmdfCvmxKgjQL
V/Nld/WBMPTA81WLmZNgP+DAKV+h+kRQVaMpIhOV3xIVpEFq0Zv1xrvPOJOLZXKY
eRBRlZc3OC0SiKpmQNf1fsv4TygeEhoAiJnp0znZ+YNFahVzF+f9lN8vjxn6iXzG
KlvSE+v8+Q7GjNqriXAIUl6NXteGVtVhFAA311OT43Cgn8UVWFCZa1UPvRiHsoTv
w5aVoEXTCLX+bu8d3HJIyACZrlhsVd1e/rt2itZ2SHgOXVH5RZhULNz5PGCskUde
wGqiNUMFcqWCka6aidvKjzext3F7ujsjIDdmfnKA/ESuN9G7j9/Sd0KWUYs29hhl
Fub8sl1YkEpG+gtJGHX+jwiQ+jrDmyKbHAkDFsfTZeXmt2GYARER5JFvHVWgsi/c
jL3nlXM+mIUzHBI0pXL4qNodgfeAsGZn4t6ynZzcAxuYid5RWn72qZ5my3YNPDvQ
6Y1fHcFnFFZNcRi5/wdtyMCKM/eAG722NZ1HIXEwLx9l/2Uit+SoSnS4MZVYGANE
qbkJyDY8zRfmwVL8TOzrrqjgOGqhDK+3pxbPMk0PLD5RFUr2dfdLFEqRjHQVaedT
9UFVDKPVEC1BmKvdxIFA4NcOR8K0GMeC8NoIm6uiXEkYSE8XGXUEizFDCBKCUhkc
M4ELn9CEUJSmKMVNxhzT8rLjTN3uGUqooX3GBvO6t0D5ujy/XWmdP36lVv/ksCXW
6Ne0Pj2RgVeAGTfgHZRFAysQfIJlsD1H1JazLKhpa0XLMCXzC7gYBMDjeRy4RZkC
k/eM7q5MFkCoSUCwCJ+zxLQkQICQV5Rj7DkJPKYnRRvpMMUnLxq1+a0BcypRGOut
qsjM51EIuQyz6UFHBeghILVGcL0aa+tDvwu5XK8R0O8RkCD92yatGeNfGLOki7So
4H45nTcGJUQM630PkUcfUbU+oxfw810dqTj5/ZVVmGc3X+e7qzonmpJ4NduP8ACC
4iI0BVBKzs7kTzoSQNiHRE8bHbHKVux97lSc3ViNxHo3qTgRJOaBFc+sVWCEpl/h
pAskG2kKkYcp1sCIlucZkLrXkueMvUw7x9F67OpszRz0KqHCFt1XTvZBHzAGUe5X
pc/GOvPcpe1BWrxVwouM/ZobyETf8gLJngju6w8tHWU0GmeXdd0vuFKX8YwFquOs
SaKqfqeBzteTYeBBeXFslIs31p/KVPDz2JbxaSjfXV8ykn3BarGZjNtOAv980I04
MxMijL8PFmeHJMSmJ9bZhehQssYypqsNTIcLPTHgIRHt1UOVgR0PegnDXo4O3w7A
nhWsBbo0KZ9mnCRBvxOHDCYhYeLUdexCIAU33IgSulrfukkkBkAB+NDGPSBKgV6r
+zORuG13ad/eECb6gjqoGirAGiNzHpY/z/IxUGJSd7Z/XzhZ+FJjFc0AsUCXN7s0
dg2F/JFLpIxRxQlJk13akqd7Aapso0B65X7CwtGZCP1NjE0Frgv2ZGsp/VL0Q9hq
WvDDYToP4kehxMvDkNywxv1cgpyXTEylBb4rE+o9k1L6I52c9KXI84BwJp2mBdjG
K4lW6Sz/aWQRX26bbcbDkBUI9gWfLHbcl+EKLRo2/tyDLwOE0ZwapPKpePKV71z2
C1/0uz8Aw/ub5wbqfDE+eP9F4TvbPI6HzNRrvir1LD3Wm7RhL5+tZNYuU4yBnCJd
sBSoe2OKRbGJXOI+riy0D3/Ix181dsF5xkOU+lRETjzyEltXOgXyh04Y29AYvuRb
fnnYXb2pzVCFiDyXSADnMjiODVtP0u990kAYKP8kUn7hLyvMlj9EUUQMyVcKQg8P
EhskwOMkpqfsDYCiPBhQkyVMMvY43VT/ODQ6toLXNmrld9ULve9zbYoZDyy1khk4
RfM9gAF7cGcQqD1aHrBpvgm0rsD8tMPwPQiVmadOZeUPyItBhjlqfH3FrfKfqkq1
aqyC4eyJSmlHoYfgzOKZ4ZypGqM6Ghcoyl9kye8ukrzjkCbVdQ8TSpxm8tHJTm6/
6eOuJniRSeKDIFcIzBzZdHiFY4q/Y9I1PXGnVUf2/EZXLN2m7xeQtjpW8RMlZCRy
zwFtuf+fFI/Fuc5gyTWVT8O+wZzlT9QYThPq3EyWnYDLLedyx+x/MRKP/ezTehmx
MRw5YZ3tbkRAx1WnAuKQL/rHkSP5185gVvFqw9XnCu5Wy2hUww0QjC0hvsTp1jSD
+wh06mFHsc5tSFGK/prVbwaIw53RYPe1KASUT6nOEhioew6EjLZg9YH2a26+qg3m
CU3K9M9K8Fn+8xa0WqhG1cxNjqsb/vXy1VJyMws9PjMcLbpxsxLd8MgboR7oxLar
Iz1n8GIQjSkZi36xxnXA32QckT0nj0YtswzM8UISs2WxwQ9Q7OLl4idvy5oY5yox
ElfA0K16wcstXMfe8yusZWZJj8m7Qr+4zwTEI9xfuKA7ENhnhp8qBjaXC5t8NBcF
ml1rV/wxWmhO050gzzoU3Rfem+KYX14obXxiWO8p0z1QlcxC5zuOHZg9A2RJk0w9
m2eOhGnJ8SZSPjR5uNmdxT+BbLF/1ahyRf5Jggo2SGtFGnbmANGqwQAMFAxyDkfv
xrkWxvRKIvd1e7lRwgzOwfpjKMmWdgc5/uM/vGWg1Ou5XsAiphWVmNID9148HuIt
gTUhwa6aPBLvo3+JC21xB6nVf2DmIA+y6a7W292uTNFFnyXDHTUZUb+Ykp2eiGDd
gYRwkxWJ2yOwI48oQ9KotYmHAHWipfiuhZ3ZK3O9z1phCOcPeIa2e/bCT38mN7Pf
7hC+/aXTu5HVCCJGghF516HsTRDjAW3izt19Ns1yw5A8sAlSlxP6uP3Xbr8GkGl0
WuQ/yG24p0bc6mNS21ByQ4XDWZdT0G/0AA5sBejzBE2sm4EIwx9t4eDnm0l/oBtG
n4VIl6bcBpijFYi1HDs8siGoEkZp+9wiu/4cXpUGz3ExeE910KKPleNuTDkwM0C9
9hYOzdRsImsmB/hoKqKav6vkrVYCW2sWdaM7gD9KxWLUJvjJlsM5ezuN3yUzR4/8
fTsD8DEzmO1ywxloTlmK+BjVi+DLpBKqEQ3/2mcYAZkXB16jrFiNart0URreRuQ4
uiP2qxk5n+V6ePlN1zNxBoDAiAMXpt30S8axfMCL8V4LEdv4FcqHkkWcFSmbDR0g
sHB7+7ZSflZmliggUXp8P5A3EQrjsXptp6c4dNs+WaY+gpMxsZUIWhENkDPYJfzI
n0bbEaeLS0ZME/iqYSpy5SIAv9t1vlcKLIKumj8VcRFU5mBc2Zu/ywQuzqXZYJZ6
JTrQ4JHh6xGPOtLWQivocOmUukW21WbKVkizkTFH8Y7xghQT/DQ1QR7tdQvvopJX
wLNZnOrNLnKWoV4JHL0a9B/A4FciD6RKKg+FHwiEXmxfXxHXBNpCLybRrnBiANVi
qNYUYNVlm/r2nIt1EASroJ4Dkl91Zg2PD7MGj5lPgXJ+d68Kp77ANtETADYgqZu4
+fWPeBZZ4YG3T9zEYHYksxVphUPF+y5M7IfKgL2mx7tnoxqkFNDuoH0IQ4MreUUf
bmv97KHFsi/ljvHxq51IB6wsjRyi75wduIdya3spFoMkZCsBcwt4hIPoD0PfWouB
rQZ6DZCHgFXaXRHtiRamSM4tz281niwNZnRRe3LgNM+HAbdS1RIS6dgaxDygZ0h0
9tXP6QQbKA4RTuPPzcTyLWNy8EXy+wDxXSKY5P82jAhPKtGdI1c4n5FMZ8dE9HSS
FJZFLKVVXvMMkwz0MFNwsYzTXGE+fH+XxBCvL4xA014MtHT4fbHCIdb52JLvLylb
erHXmSVe/Z5zBjB0DiG0Eo/qtR1kD6b/E9Yf3mg9O1W9kK/eZbfw1uvPjIjNAQ7r
NqnYMt56b+FN1GwocfYcsI+OoxSY+bXjeo/9gK+mp0OVj9Q3Pezb6efaKaDzbR84
OWjJ9kfwAC+Jtsml22BirWFEANow/FSHrXTly0OnNA6eutgFZ90JT5+ceWT/sjFS
zbwaOCKAVTRJxV6Rc+xU39+bX1FcM5g1K01BBVoOIBAXxchFLUSyMwoc20FM+t64
eWlpM3LH8HeaEkm1FCKKzZlDGkBISdDzOl2FNPmFOXOdJ819HkT6YFKJdVmV6eHT
4N7kTly/Hik24gj78yatIKFgjEJJ7N+icX2jqeParIwd/Re8l2mUq2g9V6FuThqr
9iobWnMEDTFyz+RQzN5tLww4Tb0ywlauoS/q8heKu4XcNxK0DkDoDj1nKTZxQDOs
ryOXfw0wglOtelsNJBM0ccW7HX3BjtmBGOx5ZJBaKzeYDhlnBPjdd0mK5l+eu9zF
9wPxP/ht7DoUYZbeySFTJ8Z9fu2MSny/KzSJ6dKWYEgT+rswXWuTY6zU3hyQKJ2E
g0wq5wJdv/Zjz6hMNo5TjWMzSOylvP6gPc0JQYWlHEMAA5BbbyM30k7i+MnI5WwZ
h1GPmV6CA0SdRGPtTOwmD1RsM32gyiGcaoSpiDUgqrBirgyoLkaz20qBEoq4m25q
fLLYNKT/Leue5aCYrvXvKFTEn/jfabZLusfGr00pzSefR7GcTooova4AJIWDg1Lm
BBxrgeE2SVP6SJako+wjKoKzuFRG37gctKQLEYYGgJYH8leyd4WgK3POEXeZbDSs
V1cebbvGliQlwFPZXw2hniWkHazobQliyqzyWi9N1hb6+G61/c68srSphkCnOdpF
Ulr4KWRG5/m9Ci5NA40id2VrMw8JxvV6uuM2fc6APMQl/6XWXVtzLQi5GKBcwGPt
0Mn4J9V5PHxdhn7zVn52LmY3R5RQr9VK1iCFDC94qm5rnzqF9Zzxc7ZmY6ONZOb9
CU9z4Yz3Iii13scPmz1KAsg7jTVr+VAoz96vB45nAHxiol4PAKd9rcDo3x4uGbo9
xfhFJB20OkXw9jCEQiG+XHoUcrClBcFOAZYteY0eUqpLXqwa5RN/BdOWfIzGXrCT
ONihckgH1pXEWKLGKcNSIFKVcaje0QCC84j8Zucfg02eKk/8WId2ZpcLUuXYbH6t
00rNAz6x451YrCQWR6z+7VOlw1Et00IQQY+GS3+Ij8QYUqB/cUN/ymEOIbbC19Nx
dz/RsJTfYZLWakv2ghuktMToRUFgGJiRBVLWaQpp1z2wHrOrwMeL+4dGFaVMvHFE
4plyAR+hiBxljg7wi8zC+ojXjV16+WLnk4/nBpqVoI3jlDLi1hq2dQMODXSJossf
BiPiSzBNSu6WS1DulUOf+QKDBmxCjsWmt2gn6N4CXDdM/d+t8BIBWCO+Uc1SWXc0
QtVkjxzIZJgQvgn6GW4hzBrYY4oFhDWmKrHuuXUUME6Owbwz417R67N9NJ0Ct9E9
+RLGDrW2c4hNCrAy4CzkGWYihO2Uq4ofR9/uBAW62XqpDRS7gka5g5EKr1tr0wGn
OA/6CACujpFRETSa/bLs7BkUa827XAo2oXaa+Ae65ASFif2ixu9ciCy85IQoAkhd
krtgJUkfCU9CcMFB+Xi5/6MKctHQRVoMIw3+/sV1X/xJds6A6L+XUr4exGOenCzU
lZ9K5ouWLnp8j4Xtd+7iGcRmNwCfFF2S/L0IN6oq1ghCRNHW1tIhBgQyCpfJzcyw
QqY3pD/w8eSPW+R0GzuRNBgaHMki1YP9g1AfkiMEo5mrxyHiflwtT6uZeTYhZAVw
ZlEf2S+7XrxdeQ0wvfhQBfNkdQ6Is/08Enrtlg8/cWRA47avyzwuLkGFABm8i2uI
pIS5fnMX/MfFQk8wX6xwKHUmJ2rmQYxpGrzE0LV2o/BEBARu7z6lgezFU+3b6M/y
HTFZP/QhmqnFJobRSJAmPt1AmVJjeMdmnfqbOaBYFvgKZFzX2q6XcG2cFVB9lSnm
j8XQjhTF/xGSzQxFH52IbOidx0m7C5u8fmvhyTJbFPvLSMNLalpwWrtYPSQF+4Er
1SU4vUaNl0z14dz+MePSwyaIiERXmWsxYDsf/l/D9gsSaGb6zxA8vlTmv2q9frlj
fypIKhh6ZGuYhgstQPIjrifuckZRktISSadQhQ69kKvQb5kI9u7jg4OQCSozDe1Q
+QU/Abjlza2tJ8+1XXIsZt9vXUWlhnPeKC19akLEC4Pidm9OGUDB3dUjkj0sAUN8
SPTeTfomFT3JiNPYWhyy8NEDALTbGe45niVdGuxW4uPi1iZjTNGHOCgb6YzUsXaP
ak5FJHlMZaOgP2RktWKHtxhaX/rP6rkqX9htcC17Bt7JFCCGH7nEsVuHnGIF344i
Dnltj1b8eUy18pB5dP5OPDrCL4m6m25Ud8z9p5FQUsiYNPa/Lk2JtReciEzCYfkI
xxR+Os/aAplq8jwcq01L/2SHcVHKzJHYV7kOC9t8detqYRaha/ETEQxlvsbNwxSt
b4TMlXb+TMc4Ygynm0zTOEpYvVgdKEWCc5wGQJa0LRi/1w755KjOXPCH57VkdhIQ
dZaps8NdrsWDRBJuUY6G/DEb9J7V5afHXFka36SMmS/2GgHCjxf5uJZIAOJ3gEYm
rcWFKLYFmFC9WphwtbJ3/QCQyp7wXRu6imWVAZgsX4MKTG6QzFN9NXSnIh8qDlqQ
G0ewqoOaAhn+nmgiNUi9FwEfIWUiCWJ+Kwtu3Cv4jZzMPaAIvdEoaaP4d4K8kmEx
V2DszuWS8t/hc/M85pu6BIdK6uWidDXQ5CYlKz4tzwkpg8jAF4ux3HgMe3SI+Hgn
l9uc+kGcKcJux11X9tN1/AWfxMWMCG8sGex8myyIZfDL6FAJEY8FI63xccTK29dA
DhRoQsEyhUfbJO+S0z8fy+nsg9TvPhdIEBluP99l9WCMBV56ltw8QpcjiHKD8hpD
zysCFh2nhQo1YAvgkKri479jS5i7mepAuQiLfNP8ZXFcQyCr9WTeKf08lP8yR88H
lN/tSfFdgu50TffiQpAZ9FERNaOWJOrvek7fqJVgvNxf/bUapCD9REHi/CsOCeC5
Qi/i3ZQ7RkA4BuvVBVgj8tSZqGW/TAgSF6J+91Hg0h4vkEM75b0qE1CYNRzr99id
bJ0bdRHSoX8UriSI5QRMxJyp5eE4ItvD2Ss7h7UBaXETfXy405vuDsMhsufCguco
f+9b16Mv590Er2NchnkkJW0o7tmW7PcCquct7FQBXyJtNZpd5AhCceCMEYQTtO/e
kIK5y2oapoRFy2c9gGfV6lKO4AcZ7ou5olaquAFwMAYrOcfC+KCyci+lq4z7SPZ2
f51qhNOPE0p3IdjW1nATPJSa9lwcueG7k2UWSFX/L8hMzWk6/TyHvQX0CaCDwqEF
TBp2G51KNxFVOuRs6RdFSb4SdBSDB4q87wma0LCyGRepQl5WDKnGPuMIro1m9nc/
N8/Wj25QC+Y6UmUj6U5ihtiZPDCQYlHel0vdUfUfvDxLk44zd8v3nj/+fccow+UL
tkoLMKoem1LeO9bjMeFga+jRkCVDkXJARdfoazIwNon1DvNVhWENfl6AMMjo5Ne7
+4V16iL/bpbT9iN9f4utKL2ZyuKKxHvKO2/cb3B0R7LHErAmuLJmj34RgZJq2csa
NJ4HYBPiOy5bnse6KD90cpiTWo4fPhJidqEpV4YsqfuqbeLMQ1DEmuofrZ74aPnc
U1eaJBW3KsMbskXR4ikeHeGLmnSLRav5fVbUBT/WeV7P2u3DvNU20HaCVGClsstY
gaCrUJ6VsldwmUDhiTflYUSsq59fT0zlPW32G3rLewO3zcew/b173b9W1ithWlw1
H63pbtEWJX8P/jBGBxk0/+pNFTXCXSSGqTS4wXMoZDJfe+vxvm5EieawqiBcuc7Y
Rw2bsd1OEP9fMszoc8eX5C84BcB2k32BKmSPq2KapU+sQ7xGeEGjFUp7viJUPl7G
CCthjQ3UPHT6kcChLbrywROJyvNVuFFUimaTRn547MkmX41ssE1qRNjVnkam8hY3
b/z7vvDrQLv7hu2Av9fiYnMYcUhls2TQxR3W+IjscimT+fjZyBaWKQAVM8u+gJqt
Zs46Cd9nmV3pf8tmtXbrQpGnHdxh5mzib3EFBTEj/IWBosLziDviRGgbw94EBRHN
viKKL8d2vOaltJzpNpL8ZcPtPPAkv/48bfbQ28VXvZa6vsdGdR2t9Fi5B0zeD7+1
Y4rTX1PrQnW9WLX7ykiMN1tAlzXye1R4W2RrObGEhKsaKwO+CgznYjX3WuNjk0cE
poAb9LT+WNxeyxPm1n77Z966ktjqS/gkKUSCSHKHYQu27zwndtCCws6hkma9mkZw
q7lQXlPWbPpoym7/c8A/wHRu7Bt8SeM8mNTfo9UYPwwvpGEi8fu2u2dZBDedBhaH
j42N+uQjiFPjPZRoXul+zdWBCHX0LwRA9i394/p/kN4jWD3dwSaQf1CkvBPgSHaw
CwlLYKXTifRldFp7LBnIu0IK3AkVgQxkruzDaMfW0ZECe6lU5BZPSUQ74u6PhPFZ
ArWoD7VJGtJiJ1mF5d6yDL3qPNRrrKGz3NFd2sHxCU7E26D2PBjHXZ3sb27zDXan
xJuIBAraDL/ROcyq9c1/qkU6h35dfhvUrLiKlaGMfe7LFo1Iw4H1+yapkrfOsv7x
v7HqlyHrStt7o6AeRXL0vGBX4+0wxAgHyJ+6OLPTZOLfCTy0B7B+TZSH+byATS0H
KbWCYn9jINd4xuf84MoHWTF7Sicbpfqz6bW720zKEJtNFk/fd5Qgl6aif3ds6+gr
cuQIts3dtjmqNwmMHaRXDywh11MQizYML5+kIQRHWU9Fbv4IA1OHSqsjRPeoFVP2
7LogSi1/ta5XanpViMKdUZL4yC6knD0qdB9DBEkMJ7nM/MZshUYZjoT0HBSKqhJI
9BNWi9u9qcuytml/NEnVBxVbz3jDzXRFQ/VK7QAb5d0WiAx123g+uGwY25cH9b88
hPva9oNTboMvhwFf63JFlyavzDN1E1/4vNUdhaMIsKKjD7A7EATzQBAoUzM4SKoK
wou5Ua/HYbg/YwkRMDvhtox69IxB4axysecZj2mQN3lOiuwDtOpactKW4J1L0whT
sDQ+JuY/ZzY/h2P09GKJZABGLXS9SY3qr0GntxipumeAUzBUiATCCHcBtrYtFTgI
wZNA4Cw3U3fpVegCQT7o9u7Caaha9hBqMM2Bt+nJfUFOZG/wwCOtVz6DnEN2bTYw
EDy3JHcjhH1dba0pfIiecv3/438z4wY5IZ8NfnaZTF9jbAOdkj5w0sDfxfJaKMQI
iwdgGtwY7vGOfS2nCLgoXSoV5meS1VPSvLK/V3RB2Dafvturt+0/8e5pausmG5+O
175KUC5Lnc/Ue/dvdH++K/oO7CW28rOozBJd2vBm+QBw5o+3HB7asEMr0cjurpN2
C1kvsIUTI7TVKCYOEfSwAsLGoymC0bFAf7jHnPlNpzcmPy/+Ln27Zx8d86AozKQG
J8iLAZpvpkssh5TbIwuZHtPZUN9MA0P/rbONbXsHpo5355cGT1WCXueZM95GPCed
bkM07m911TAWTqv8pXTevlSyY+k825IcJRy4eItosixj58/VvCQQLguHaV+jN0DG
u6nesYraAyxe3A4cYicgqfh68WbfOyhe9IkWvzFsVcQF62JhnYe5nWq5GPRtabx5
NouHib1mJesW4y1pwRuNXZa3taMFatnsgaF94BJf679Qn0pYKMcsrC9MhkmVxHtJ
PAIzJpY0n2Riv431cd56fsdOjNY7ARveK73j4Fb+BqJdGUNkH2XYRMN8ovDuX8yx
KpHav/8n/TmVLLf+d8h7kpzbMn42ClIDAobTvz1/Khexx6K3QOaavrAd935iPp/u
Rapoa2kT8kNw2AstFIYkr56RZeyRZrYa5cjOoCPdwB+ZSwub0Dx0aMWSi3ULDGff
H60QKC+w1MXLMuDisy1vo+HW2WT5gbvwnM5juih6GtLw3iHfhQmRt9TfyO8NFIx8
Wn8jNCF9FyRHyw1QhGrngNS5zuuevfklgjLEJ1NWAZGe2qCyyYCdZAdtWVARlTrX
QYVc8lilUedgfkA3jjxDAXWHHVH2xugxK3h91DEEv+gXIi27C/eD9DCqLsHeHJ0z
L9xeG3sN/wo7aPLal2LGSirffX5lEw9Tro7/YRB1FYgjaq/ZNeZrkMbwchBOzJdt
t4IOGMxdGg/7+6CJNGqBWaJvQgZFlBk3Q5UNQ8ezx2sy3/Y1mUg3OVlkZfWho/eV
fycEGOSzLkd8kgbvU3pIL4n4Yx/IagncexaOenH2a2sTQpXqVNJgwwYtvaIQxQ5q
aGFqmrkUEBmzeVPc44/aFbTIz4UVjlGqQxerLwewfB/aFfLi3onOyZPdbLzzz6MF
eSWbPWUxu6mjyMaTSfIcRT3Two2wG3t6wIjSZMKVJEeb7kzEBcStG/ocykc5WEJF
eXugvhEljz1jIHlANzbybJD+M85QIXbBEG5qDv/bmCTjqjxH7DYozl1QWkSIDe7K
gKVwTku4WZV09R4OupgLthksFLzIIcvySH48vu0XM3M2cIPe9mLl5Tbf+K+/rtG2
hhhOQdGBmo5Cb5a3H6RLJyj1E9V/vM2FV8Y8wHgBt1OBtbMHZ4YIyx049L/Ixn78
/tHxk3kcEairJEOqfpaAuv3dwL0vxut1ROmrpEqkZpRjK3PJDt4sDo3wM4YKXXOj
AUb/TKiaemgPojnHkdYJhZhCs810TBPoPUzBFJSjxTwm5ICdo5EGvArf0diDkKcV
T20OlH1qQk3QgAN+PmxYjEM+5tLFrojAkaXWb9u/C/lAjM553CfeBWj5Y6Y1jitc
azQIUHFZK4M+mxz/rZXSkbRJlLMzukLk/ibKDQJ7L8pOXwoi3vK28/L/rf4PSB3/
CeUlcfkHr8q9tzjxIZ+LQA41LMmYWM56U0KaBc+qOHoxj+W2Q6jBNtDByT2gRfk9
aLLJ6B+85PtqIFT8nmTm6O5VoinX/mPgE4wWONPHzh3Lh3+GW5GEo3f+9L1Dr0zK
6mJobJncRverWPAj7RECULBtl2YoIJ0jQCoIomLuzuI6aLuWvpRbFCjb8qs94Hxq
X2Gp/IhI/+Y5CBTXHHPoWEIt3ZdDlrEos+kL+VuECv/xE71iH7Zcr/o5uK3PkPZF
wKb0rKsvhUYT1fZ5TiO8uuW689b8QOCZwe99P161fPX6Yz5cQHUJtZxOTERDf+bj
ubnIRgSeHi1948P50oM16EmsNFKRcwKfTL8JKm1lRoS9fcoPmQ37PkF/nY688gMK
lhqtht/lsVdeVahBZ9mTsXE/6wSvev3sy/YXMufO4oNP7v2vop+XJKSlBN5zj3VO
W+oy+z0Ls0KfI7Rrf2Dkq0bQm5Zsvf7WrQ4Xtw1M54Xqui0y7RkejF5dLrgtOhmg
cjAN9pWpLvcuOgvPdKXllWy8v6wDNoS/W2pfGeT0PmTg020osoRmrmspcYV5dvNg
wFJuOHvgw3/CbS4VwVPvizhqQ4dyy+KPbBnvbiVaeReZe4LMOtXohLe9mtsneZuE
OVCIumnSC4jjb5YnfXncMvNv0jL47PFjRGMmGR3l5vOnhdlG53XjNQpjmHOWhsrD
Z4cLJJHoKkq0tYl9X3bDQQLLt87Mh9bICH4fd+/ulCer0ZT9p3Kdu4t2If+VHRo3
QnFaIMTPgEnZL9ibllJG4cSR/q3P1vMkI6Q6dtsmIrVjwlSIhpd5phcn6rsZ/YxM
jNWP7kk599qTNdIXMGTSJGJlUBo31CiJK/Tgf8vb9p8GG6/nlHa0y/ZjE0OUG/FJ
kb+OdvrFX4irj/nU0fMvBGqtO7aviTzV0EoC40tZJDHqCTaF9Uvrv0kPmRwc569N
Agxk4rf8W1OWize5YQfKqssTUYGHfISZ9YwbbKB2AWDdpr1w89YNj/ykRG4Om/Cb
4znEbSssR9/n/F0KG2f8sPUsaLNqfGFJcelHyL+3WdppoYFhO4CMejPRLTCeeNmq
seEnH/3xCVVX0kLyZl8Hf79RxFi/HEY7IbjcAGYL5FTtZnW5DT23GXWxSCC4nC4r
YRMC9wb5vp2wO3vQ586qIQVkoQ1yXLHF/XKWURtFQ6VPjZOhxfi0hSB9v2IvkLYV
QOkS+n+WyY/iWKhzffSJ28ot2iC/UzfDLXz9PvkvL4M+h/bpu7uw72owaG477q7A
O37TG3+57m9OFyhQ9J7lJ2m5MrIIdgqUMuMYl7lI8xdZ2RepdKcDBx6lMxNOjc84
/R6jXQSBg6+R+mIJ/f+qcVezb6fn+vE/e0UKvPCjXkDSC4wVMKGiMky8FpIvbwGn
YQOUDtfvqWecruQ1NyR4sBjYBXIQr9Wh5YbBquAsc4tkA3WyPaEG4ZlhjUrSbpx+
NFVp65aqYylJvFRji6WYqd/QpiArC8n2zSTZDiCGnBaJ38Zk0kK1F+ZlNxceAmxX
xVpY1ba3Saq7Wt8y5aHKHCJzTtTCfCoFbuhS7p1bFuwC0wCjJbiS4xLPrE/Fan/W
+E1uk97nPYF2JLyT+nPEAU7TgSsCcGGfQAaQ2cIPQNlj0SfOXAEJK8Hqtcf04xxZ
ax7BsIW5yPlA8WhpaFuHoEstkkc4LhDskV62pBFce4LxGUdtLW8KgYKmySYnbDT5
/uaCvBhyMn17OinGSo5eonEo9j/dZVUqzqpwQtbSMoSZwgc9ciXu92cNKO4jTbyW
IpmlyGyysPwgqjNjyavjphx0B7kGAaT8LE/pObSxEGOCC53p0oEjLjpQvEqipiWV
78BBTr0QFjYag+mJ8Ui8WdOwoLwZ8qLc2jdqEJWCl11lmwBqJJzZy8eYQoehBJ5n
Q+pR8uaKyPSxt0D1MxHH/ktSYdvpXcI9IEliLXEU6JWZw6S/Yqmtuy9iEaeCJgww
LC+1qaecfXW3aWmk2hJUyGfk0UzoWapgY/ZYmIBR0rYCTpQWfH9lJG/aKo3pnbJ4
uZxBztpzktoZY2qi6OLlFsYTs0c3lrov+N+NSj9wm8YpaKdb2Twsfayd22DypWRI
YOh1AU3Q5TaUe9LAX1+BdSc3fknmKLV/796RP21KX9Be8sBBl3D0Hrxp546ogRGV
ANsGYZY6FsKXtv6KXjlXkbjM54STvT2ubGnwDjWYWwzPG7/TQ+FDKmXJFsFyquDN
fQp8wC71DLUhZToi3HQ9gk0BW7Fn7A7NneboeDSymNdmIKbPrv8ppQ6senFM3YTS
rBqHJ3JunR8gU60Wbz7SCn9vWxYtk5Dl9zHSKvbZT2kFrfQt0TbzBNPeIJFlbnXn
UJ1hrQrHCESu7juO0kh87TUJe0/rAae0n6aaGEKKGN6xOyqCZljnTGDNeFBs87SW
fYGYCqr3mY2apYNRd+kDbmeMtORLDC+GF5dXo5SCB+BvvRLQ5wTQdt3nIVe2BBxP
1FTdw/cvf6+xBUwq2QdHhNqUZ2x0EecY2WAFBZ+gmbITVhNMLpCNAlLdUBjitieG
gDcMc8oyLqJWb2RNyy/DeGGbVNNWjn2wrzpTm35u9UAo3JpuhNweo+w4ceR/8o9N
QlXXOiXsAEQvd00GP/oOFuWzU/Y7qQk9ZjyTuHVhXTRBZS4YkW/J7uJNxFmYTBgM
GRNDnEB8/rebwwcY5pHo82GmXat9dULwQYEubNabQS1Cd3zBpXuHVI11GIrpCpBS
M6jH0/F84wLNh8x61lNlPX35mTDxjVWW68Qj3O2Lpdqi7An9i2z+ZoXXsDBOuRxr
IVDr2gG70C39+Xhq4M9HbRN2HEDIqxh1AN/TRSRrKTXAGniVRHbIPCok152XUEjF
gs3F6Xqcw1KmpkOZp8yQJcb/hS4OD0B9qhm/XdK1ysxx/qH5jFmXxaJiHWghhGll
K7iC7Oq/PuifkkvC8r6NUDCzLjhSYrnqhi2VNMe8XGb0bfctLC7bTNDhpaPsqHcn
jj7Zp+Ir3XQTBZ0KnmzA41pj2yE/sZ4KmNeBp6kQ1bOhz2LZj931xB6DkfYbDUFr
ujQMcMu7x05xPwgKlweZ2OnYTGRY8eJKgwBWFb7SW/Qyns35pCpya5zT/2ifodKP
MVZyd1sjwE0jz8m8fDFnkwLd4q6mljdbDrWfdWBZz5/Z2DxweGjjWVHn9bQElA53
+HuOZk6k86VA/dTOqtFG2VICOKr6fuC3rLHvpDMlf5u43WTOnf85YhAcBKmlgJ8Q
yM1JBAuBpnDg+5Y78iFqvoR4OFW8x8tq6VoN5BYb9p1v/mGvUXzNbe3ZNW+wtJT3
SAW1y0Xoq6mq8fZQGRfSNdWLgAf5CnUH41zHkyhHsDg6W7k9Azmcc7Jy4rmWmnkG
R7pkbJubhGhP5T5fz0wx439LztSKNYYT7rgmceQ2h4atCf01RyFYTQQy66Dyzydo
OZzsAdwea5niqQ9BDn3L27cxy99m9hjoqh92e3Sfk0vYyf9XAXCHjWbSOCFVxi0k
9pfsYHzquM/422xqthTJfhprm68Ud9sXJq5eeSoQTezFZYaHidccyKoZlYBb/9My
f1YRrvoY+mpaHRjmUY/vS/TZMiGs/V47FrLMo+oSZtJ/20pYaRk51XqCgaijI9Kj
UdQEfNJhFgtA2mrbH/QpS5bcGItYsRnPAzzM7ckhlcLa5JfXkPJQ8fqPFkI5r8Cn
q+gejbMEFaMXdDnCcTcE8MOLSffmvlqZi6FqxiU6up/RWVuEWt2DpZ/AX7aIrHbI
h3CB2/IjZd3veJ/8SU/6jkWwIaBEMx5Fdlla824QHQeLcZKw1Ze7Bx2r//pCrouY
+jWD5U59lKyl6t2vJfvwdtLqIMpgDWH9vTvUJVWXEpzyCh+7kXey4zVmhvoDjeM1
0S9OGcRZ59SvP8ckpYP8jKceITqUkuKErB4AJuN0Ip2iupDJK2DQXBXDKCltdYaY
St9QMr5TItJInG6QsMkQFJwG3AV/Q2lDjRDvt6Z6ADJKlJZ84952tMbBdFSZnmOb
s9uKwP+1ILhejAMB3wM8F/cNKXYDF3s79A/bthfVgltVtqmQUFCJhfdyTc9ZYlHp
vIxu7R9/21btPI+3+kwszZ46Jqyxc3z/JQTyKrHm5Rx2g4zYUxO+B1mSQOEpX4lv
R2nJVLg7W9tMfrnhwMV7WxnOg//vRwSq96qwxzEG9P4huQL2HLnbqWCcQ8MWOiAS
OHFyvK9ZiZv1TQJIUFCUNtmqWT65u2oT24xrTt9srEuRJGZAuEzAuvFuFZp17sb+
D0sGy43CfPKaf8bTr5NoA+/wV23yVztxunBc4BbT+DkZmpFgAkSnKbfwHizOleSa
1l/o0v2FDe85+O93+ZH58wRIfkhGlaXKcv8wHNA6IClgZpwfNWgnKQN3wm/aEA7J
BeFtr5UlNsEnFdmyewdg+JS26te+LWpGFhORcVmp4vtR5kJa2miU18lekbZWfiZJ
SF4v1qH5Ay5XIflqIL6k4UEpWpj52YGzKazbXIsJg2qEGds0y9UYKpGzO+uhBKle
niKdF2UTD1c+jui/N5iCX63tuPtuK4wPnTyKINe6jeaY/EJkQCpXx4JZBQouPls1
o2QSJHB0kAM1zgoDHqFDTqSaqqN6D1xGjItN/XGeYNKsaTAETDzmUWwtVuUukBIi
F4CbW9yJIDMwx7l0XrkYMR4rEcv1GYKxlG4szZo9PkVMfqxWys8eC8zVrdD3hjx1
akVdGuG7L9yGbQvnPmnbk6pZoPjxBCK8YNQ7oECxuEUPoSikBERfRFsTfFzYnD21
1BhtSwe2NTH5oSScf9MxBJ8JVPUqQMbzNZgWBegL3Wr6/MyhQOQMsKHP/mxN9Yqv
ySKOlf/tKgZjByg5w1iomhqF8ee1hEnegFGCUqQC4pl0nARAwxJM7lbeaNyT4KKE
R9jUJAFGSknh/kg07yPp1+sxVYVKhTAiKHjaA0m6AkIUPszBOU23UBRiwhkPS4/q
EOxWsp+ZZ4ZaJg0MfaxgZqK8nihLo8SxQhrPDT80TncbwO/hsy9DP8OyYON+4xNK
D7t51H35qjZk6+0VG3ijRppVQ8xpa5wg6LWdSW27dZoXqzf7JQBAcfQA7+GON8Ze
3dlejl6G1tQ0cA9vTFM4DLdgrW/yUtJ82XzDpDzF5XxzypNhi78X389IVp5eWS3p
usr5nCDee9FKEX4Wf4vmXA0XCSiU5cf7kOjzAPBcKvLsndfhg0q5ueoSfZOmp4db
bXxef6GRpfQeZ9p4/+2tpVWFRL8FFKECNNQnym4AJz4/urP3iWIQMcV98+DNjTos
EGhvKc1WdrCHrpoj94GD5FxffH8RrdLzwh9Eo6PW4oSoChqiTl6ITGnDwo6Vy0Kb
Ui8e+2e+lPiM/bkcNKwx1etjv3L1frYQrI+btBEufLN9J436S1bREIv0pmz7gRQA
nTs9D0VjtTQpreYyMjliRZpW5i3b9V94jRDLgoEA22hVnFzs4JN0D49uj87NQyeg
088EsicMOJW/xbCDamg3eydR6D/fOAirt4r7RYkpFafeXTCQEWn2W7wJIP+z6OYT
V2ZAZ1d2LJs0mR71LeRoyNNIJyTTbb9kw33NYXGhHNVxdTexzVa6N2d/yXPWshSs
a1ULTA0F3Pza+b8n8mYgN8A39XtWjFKUPRvgZjeM/XKZ59cu+23ulCkqQS9hqZuo
gLcEii8wPGF8WCbbJN7tlmqmRxm15UXY+a7+rLmkua8UFOeD3hOJIwj0N7EzHhVl
06KzorkMvp9viigQO2K5/9OjUAF/gsrdUGQLgkfK34fMIwZw59oDEq2bWjZ/gYSq
1g6KUpVeaExRXuh4B4y5lYUuG3Z3o3KbyyCSptepwc8TmTljdmq6iy4usowsf3Lj
4R4xNclHhDriO1tDAD6zhe6k8u1Aa5CGuOyNz+UnCo23fdI/pmPeRfsUameniOjg
V9jCvWbknD8pKU52R0ceecaOkEPXJY7sTAI7wfirYLTcXcKIPvurxnQUs/v6VMiz
Fu0OP7/smY3JxpBKygY0Q4pKV/d+tdUCIoxv+/dFzGHSP5raTZwX8Ji6R13RitJu
hPDKGNnuT4u0yoPxoxNJ6Fm+UHR+se0nmmAsI1fxyVyJTdptfjoDbx0XEI0cElAu
P3zwqQJqH20NKbT0U3rYs9xemQcVkgLs0zAWd0Ex6+hIYD3qvbZwpNkvwE/8wosh
/u+8b1FgiLKJ/KdS6nZ5Bp2LaKMoOE2qIRcQz0sSJFTIe7fbW4w2gpeJ0tde8UHU
dudh6wUV9VgRnNPmcmQnJwK3U7iI+LPhzlIBg5kt5ed9y6lvh/AOdR3Usae6kN0y
9pC2NLg+K1bH4BkBWNTxOUlLB1Jl9VvAciuCx5gCvgY7iIdaWE/ffofZ6C8dzhS3
B+xK5my5sHz0RVrVY1obj18BHvcUxXCfC1yYdRda07eDwL7xg91wwnAg6F6eg+kl
aEdMLZz8esmTPhhKnf/DsCETyyqAjHhXAu+13hszj5Qz6dLU9c3pmnOhGF5ljf23
Og2sLm1cU6wJxcGPYkIKcNqqP6ru+7ML6jU82q0KVSButF2KhyFBeezuBtCctIU1
C0YNOXYnRIlaZxiV9NY7c0akN5TomuHP2EIo80O9gloyHHo5iQgs3qxXMA2CyCDV
olzQDD7RsNm2xpJKt3SzDNF6RuPdt9WSyJ0sQ6rXEvp9sOd2MD0zvm7TeXlxqEoj
FVv+NnH2rzmCdN7WxoL5zip558yDxktCCgyjcs3b6uLlBrhnuSldUeKEKLaba0J6
SLG4wxJrgUS9/cFGiGIapwLEojM1JW0KG8h3IhhteGa34DLR1og63D8gnUlbFUim
RzuP5XC1L5/4JEGMlSlJrwdTJhodB+20YUrOFb+RYXlHJf+dlayzbM8Fl9dzBLmP
W6RiagoWmuCIHRZn9RFcJZZ+w4dPnE1iDt717K83inzsDrAeVA0+ZyNI/dNY5Cel
PTOEXC1W/izzugk5E7DT9oO4/arxBWyRd/3HuLZV3TPUPq57vCJVlxNFkq3c/Ub7
JW+lhXmevjVDI/UJ7K8IBTMYD+fRBpxf4Xojq8qKI3t714qZzEGwNLVGzFoXbGte
Cz3/dfKboj4TOmntgrqA+NUtxKRkGSVmglN758k2LSkpQMp9WGw7+xVBb/BLFEif
Dqc95N8tgM3HlZg4NSrwGY7CuX/hETafWFdCseTSfWb+SQAXdOi07IYwHaqcpBWr
QmikibgqHaPl8QSF28XS7oZWQTwVHWGYifJme3y5DIn7Lh7TrU9LdSJMgsWntabU
Xue4E9+zL3GFB7712Cw/OTCKej2IPRyOPI3/AMPI6Nu8vWYbYRH6l+N94axS6lwB
kYtk4kQ3d54Wa89l1vcCrJ5Peie6JEqlMj2SykCaPF6uNGseFpfzBRz8TbbUZu16
jXZDgFMtjpRSxYmD53u0T93jA+k4cSNePkYhS4R0KDlHYiJ/LBLtDC8IDdSRTr+X
GxDPlNQN5J914vSV6yQ5e0HMd+G6d/Kr403khxMX532GI1DSGwUlc/0uxlGcFV56
xS559Njx1la3oS8/dA9CubthkM1Y/8oQfAoPllteapDn+6Yd5hke24m15dsIdCEl
CLNsM5t9GwwG/1QKBQEWTOCUChpaJJvoBhDgLOVMpOOoFLWudBQmIubtwPh9v91F
57ZqaKZDR7Ca2ToXWLSi5IyTaZOr9j/2CBNm9PrGoIHNZRNVpXcPiWQGDZP7iquo
sgWgqKxU7Sfy2zILdLOI3uNviQsWhM7YXHeKAm2Oz7NrcQtfinq18lc7g5jCsTsg
VtflICkTfZ6fLhf8YMDKPl0Fhr0mWJJayXhdkv8SOCQwXzL9Oo1v3rvL8cn2GT9k
QIYZp6rsGsKQZWDPBU9DRQF+mwSphz19jdL7UJL5qpeJOdJYvepTCr8re+QjbB5J
jeo+zqxkAoL0oMI5DSdmLqoCzKiCedZsOh1Udh5BvaMWHP+vgpuM0JFu5v+vTy48
jsKhZDo1AKmn32YNt3BU+qKCr9otbI9bvOHDFuoRrcsb4mAj0o3YlmSdexFHIr9C
T4WJX1mIqfhZXotsx08sQx/GwvBKZ9CaGC97WxGTzidz5UFbZu78iFX6G9hS5ucu
CEEUZcpATuXgIYo85Q+oEZ/T8VFQ+Gii8znXxsXEG/GhpKvV1ebhRQmEI/uKKDR2
RvWV8mnDQeoDWtQdFaLosl6CIkJE/4qTC2nJe+6wFTrITCbtuc+81QrOr4lz/Gzq
XQdql2zOQXYf5vFHbl9KVg==
`protect END_PROTECTED
