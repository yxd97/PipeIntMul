`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1N2RLQmUSBFjvXbS227f1bAmtanGPf994XxxcKgif7/KIvZknXTJj54fQg7+rw9
b4sPpIeAzWRWdWPuPRW0NHVZpWX6cSl+fyZK9fInY03i/G93TJ4/4NMCuKki695o
298EK7QeXbA0UQNZEXiZcA19hagYYvt3usKfGVBnoqBcqiM9k37tO6WZAsu4g0ov
o/tmQstVTp9a02u6u8cG6h4ZNaUrrp71Qd0Vs+aAy9OHI0PEfooztu9tGy8u4MGD
zsbRmMyuasaxpccxZc1105GLI2Xgipt+NNr5HGiTVgxbduhodJXhVbmyayPicoz7
aPOJdzh8IwVmrhMOSUXZqlWc+IjqdefhaWXN6PRzIE3NKZZyuKhy7Qz33jHc+lfL
Qb8KBBLfOVI5QOCFGwo+7g==
`protect END_PROTECTED
