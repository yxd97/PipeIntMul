`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4X1R8NqZE+JRKcgWcZlbMgbJViiD1XfZkzc072RqSq4uYqOnUeT7QriELM27lNR
x+VOLwCApDqxJb72GdsuztX10bMU5l2xkk+GLGG10yayPy2Vj8wkV/y9UvxQ+sna
y9gfbVm+J4jUVt3djZs8d233WdrWX5COY2VplGIEb7SSqjuxFg0LzeVoTwhHTRow
W3S3WrjRp+sm/kRTvTzP/O22GpJzm62KuiaY+bH5DbNjTdEv/EHb2OJJEI/Gj7ox
QsOTcwTw7FapdXx4tWmqdX33fqLYE57EmSOjefSQZoTScyxUIEuFKhnTcf2N9Dh6
p3m+64YRkEeUPNNFoDwXhvYOZsrCu//dbBpQ3hFYYkUd52U0RLb8t1Godu8tLsa7
`protect END_PROTECTED
