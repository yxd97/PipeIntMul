`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DacSNB424j70wHIATTTYSj7XyjaRRP0pvvQr/9S8jxfHwXwc3S4MVDtPobd2gnoF
LfSVK7HTCN2gNGemKOn5LDHrkeut2ieZAEg0E4/WizmTtx6yhAPzpEkt3/2zfJID
oz8fNNyqV9BZ48rAYpzsFAo4irX4BiNS1lZrs2zjAnP6eAix9kkSbgq3SEtDuMxk
2d8SoC9prlkw3bZSHgjI2F2NqJfIotbKKQK2SLDsyt2nfDXw5cJwcTE7CMwjmUjN
EO8Fbvrk2Dng+1T++YY9XGmtX9B+slPAwsxQB/cH/41J3DsdD8op7SoIl8irqsiS
alpd+B+Kgllalh/veAPzfobGCG6wNaOsovufiaZJm4BD6guQ+JmSUvk5o0GGW/+k
ozWgvlKlgZJNPr0XlztxLsr2xRShcd/VbCKLRsM7Jqh97N5pyloNiHeoSASKKjI8
xP02trmajmz25/ZdHBjo5VfkMHLrAIh59cyQyGrDJeGO7Sia+N3LWbX0SlhRc8sY
co2QLxammy5JSj3H3ufbfW41oJL1tQv4GSD1jVT0J8Jc2gp52OpfusR5eN5Mg44N
RBEVIt5rxZGRd6vszSTHjxhREdtm9FPTp0fmZoZ16I2TbUT4VThKPG97okyLfGs2
mr4Eo+T9RBj769nvZqknwB6bu7qavi5autWCSEP+JoypjzJ0X6TxgqX+05YCvqrh
omVrwL9ELFahbaby5FEFARxkWojiTHjIyCnopz5XicB5cDYICh4W59HOATWk4uCg
sdY2S0Kq60jw1/+SNAw49OuRE3t/Oox5Njs3LQ69eXl8FJjnAcof058AAysxQYrX
Ky4BqbYwRCKkrj/YWWsAOYmOj4cgQsgjCvVqHf9rYLZFNCH72BbPTHj3iBqinSAF
eZcyXZCC1R/OoBwQ0UiLiYyxIuM/ah0qipTbi28P6kmPnTfwcQ5iWK1N7SwIDk1O
38VhMlLx4/sUdGygc6sQz0Sau17vNMn7d1ySQaU/6AMZAVH7YlOrehFlTcshNUsx
eDiDlRpeYmwXb3LTtKQhVdHWnZDzi2k8RFByDhV7fKptSL5t6VMNbe+/942NeIjq
BkVQStrlgyPdUbrag0kj9kwIsnnZWK8oknbJWcoXekk=
`protect END_PROTECTED
