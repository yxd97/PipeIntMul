`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/QZN0gliE3+gETDf+1UFWbiov+foZXwX2EtC/WnP1V6lAcHiWh/UxXSu4GHmEiB
YAJM7Pa78QMIWk0ddEg+cETJupnWzUcqEa/pYsMILpitN9qQ93kpu/9OxAWRwdX1
VGxGMM8jJDNquwvuFJCRWGN8hHpv7Mx1RGHz1RaxHxi37XmmR+lHe+MWGurTYsa7
SZp/7SoeN601HrVYwuD4+0lERtNzFDnkbdrRqZsfDMzRfPactA5h551or4ALpa3A
PjM2qyy9a1kxwXdt4zcF+GK/G9651cCzWXYRJ9RJDz0bCHhUQ9FmuxCOEr2YRn/g
veAyN1aX9H1N6y9YHarLhQ==
`protect END_PROTECTED
