`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cKqUotgCIJJ3TxRTikyfAS2cx5mC2IenlBpAb+5v3iV7v8Xw5TOAJ8AxeOymIKXN
V6EyMpkULCeTYKQlE6onIIQy1iEZoaBRjyj2h11XCHjc0+onbi/5hLFaZuJi6DSQ
9xGeTw0I9kEVGwTeZvyYTUYkQb7xzQPGAWtw3ftgM7lbTdrGc6jAnJrawYv742D9
tbdi3Cq2+TTiCuLyvz7DnfgFEEgY4+6ghuN/XheQ0slAyS3jc79DjGIuOwy9kEsL
XY5SgqqdKmMP3iqMBpwyjPdnYh246xMEoi2LA2a3t4gVIj8oRYx+92Lm3a6MtvR8
iiUN127rROyL5+Vd6O1i2/1GTZlVgAFkfsEM6nDRlFC2JKQxUIsBCb72pwvZkn54
OOawhdA+EEBtEm5Ay8sQJf3L1svftViMo5cCQB8pAWs=
`protect END_PROTECTED
