`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Be99zVf7Bx6TqVniH+Jw+jImTyXz63uw9v1h+ROIwF+2uoJA6UgOwwAgtgZLA3/E
JLlCynWa73gXeJajNvIzyPaplOTNSq4h5bqvqh7mxdkMH8ma/jhEr3MSzSMmWth7
3xEhO7h4YSRkGkwK9betxR8jb8da5dZi05lo7mkPqsp2aEx0i8VlzdvtGlbPb0sG
WSTsCSNfPm4Ze9l5zEUk3zg4MmzgkWYYdLx5pB8BRLtUz7RlXlW/Vix8D9IxnWB4
PfX9sK0lJpTbhB1ruvVeiG7g0e6wPQu8FNwF9DD0SX2G2soJI5Q45yEF5fnq2c/y
Ty8MvaRbmFVbMcjIUyEUPr/CNTPuw8AVfBza6PejqpX2DfgXSVQJrf9QbkjHFxj/
dvt+/X+Slv8joJKWswHCWihr+PwOR2+27vPbZcWN5OEr6c0g3fLvrhRQvXFayXFF
tKXRteJ87FITdFtwoLV3zQBlS8gLAuxBLUlOLgHlXiQ=
`protect END_PROTECTED
