`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PcHMrQdgYZ0bFKXElH4rgkkahpsEJUE913UozotfrsC6Yvntj4+ZA7llOq6cvDgc
QI1DArVZxygrewj/yi8+j3XZiCvUhwyNYN+b39sV+abpP5XfE+B57XuJuvhyYnT2
SEx0G2FzJN6/Y9PFqVqljxUtvyaBlFwgx3gSEM/keuItaNAP7PMTGf3IRagO/EWP
GwJ3IhN21y8hOWBl1in2/THJ8n4nEuazcTNMbwrGXi3M590b5VgoM6j047zXRnBk
92Xv7Rmh3iBs7kv12ZD3M97daX9rN7YTvtBVwwopK/LMR/xMtdDzePySrss+ddoF
aufwKqMkqlY1NY0qdUsKmw==
`protect END_PROTECTED
