`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qQ12JklFwnOZNs0bC5BHOoNzCk4WTvkIZLjL5Rsjuy0ntcAUYwTZMMTlvuAM33J
J+LaebduSoOJ8reQqqw3ZW/wrDEcaedTXxuXacLmPx8drzZxocxkrbLsZ+I3QpwE
CicVI2xsVYU4/NFVfufIutSdhmYrZyKFy3cP0qaNvINfhREqtKRZbhhjF9EXBQz2
Z6rkr/DgUf3TAR3oqTdAd6PdaOr3pjGAG5Dp3KPwlMh5jxo6LqVIfggd3jl3iYpH
0/x08MWNmhTxurOqYy2XS4OL4gRbfgE7H7jlNvoB5T0pqw/P4qEpIrFxmvOYoFnm
SLWsKoYnEXzgXe7WVLLItvPlybA1wbfcBG7dsVG7PeYJPcCUHUrBafCRRXPNFxh2
ttLgW/OC7xY/quB7xhW6cub2v8YOOQ2exHHnR2UFAspXPkeFsssdEG3BhMp2LM10
mpWPgiteBiEu34qHP/ge1GNPX68yUjK+6+/tIYMxFt4VivFK9RkxGuXhY8uwluv/
tGgA9dqgrQUSmadtxDj4wg==
`protect END_PROTECTED
