`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQf5Q27QosUwUMsvRhejtYe0+tvbrWdfxY9dLll8++tWL7zsFeAIvPCqQTgVBX00
LTHVeeS5UZLXG02vVHdWb8ASMjIzOhZEDxFBJBHNdInbO/xzwuu22dtDdgS/tu3/
gt0n6rhMo3CKKYLfarLvg3gcUxKxBXAFEe4iwcLP8VSHbWTqd5sFhmTSHWbZz7y+
3szTl8PDciEYLtl53ZPlKZf71PPgJrpK6rCCKrROeh4JiWkeI70dgjx668paOB8/
w0I1+dvoNzBX4W9a986DpN2nt48q8QOvUYA/IsLRCMrv4E9Xg0bjUb6pNL7uqftl
4nS9789S9d44PuZayXDPv7sc/excVWQeLvSeZfdZbrlazbJaLZBYFAqY4JNsOEAR
1Ztykkx/0mY8tsYq9R+No9HsPXeZA8ddQjl4yo3rRNh7D6p0cx6S//q5ezW08QxQ
wUTKgBaeUJyLkgw9iOV8E/qBlbc2/iB67SeavnnOhSbkikMeCBjWXI1g4pZh8XE/
XUWxK0RHV4jh+yhqR7jQZk0DYr7yjGPFukD4QQMrncCQ4DiBP3zFl7Yz4BcB+DJ8
1nirbRKJNmUMfOR7RHYhYSM+Rl6oHe5+G8V0an/AdZcj8CHrrdxGwhrkfCCR/F7v
tss2884XcOVBOp4BoRDcsY+s5g7eivDyxLDli6qmA7fA1obSTFPpExaYOl2r3vKV
EW6rhaghcsUgTjXjlQOX+3+FhZU7D7Puzsz+faTGkmQ6Akagcruglv0SBeXCC7p4
Ac4o+3i8KSF/g2Cua9DiqC82EDa0RlDhZ/Zu85ccPLqFl2u0Qg5wyBtqVZFXBvwh
4iKWIXiAYOVliV/8L6O+CFcKwtFHQQpvsVe7fu68GTKtUKTWQf7uEAQaIAaCzcV0
dFeEA4c4e48OGBLzJKKSphfLRCMeQNnoh04gtWAJl3FpLibpkgmCXTowJT6RZTJh
ALt8/afKAVZHISZfCSv+UK78u13mwPbNvEEvnoRpZuzIhDViamVAjI+pGF1Gmvo8
jnOSSyIOyOmhai82XJjRwZ+zBl2VwvJ6anHKjFuIRVQBBdB0zrS2jaNvTlz9xlBv
wS3M4BJ/I6ei0zFM0r1yjVT8himGlwiwbRiag5iMHRVnQsFdYJIfMOmBity43Ci3
`protect END_PROTECTED
