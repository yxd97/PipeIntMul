`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2SV9EA6XEJhhvvL3Wlgb+JNn+YfggNLia1dCry8ElLcvuANrsFUpWMog5+rBrda
yCODfW+SkOi9gdoYN7MTc6kNOL94zWMKTu96nK2xmbyPuxh79FI8oVffFhZjHlf+
6MJj3AkqheEH7Jddq88PNxxwjuQpMyf89VKlX99KHC+28dSllr1fQVQYIyvLXIVs
VDkvWBekjuH3b228a7xUujDPPvH0aNj8ZAwjZspnq85wUS4gZExEsBMXDX2H7SGK
ZGUbymceABJk6LdHtuUrgCGcES+OgxFc6y3keqX+EEsJjZ+MQMS1abHzjtTH4MGc
NSV4+gGMHNVnFhN4bJcrCgSsySR6wI3yrDyyzhW1TqUyP0T8GafcHEIXShq7eGrh
eMScIllQFi/DQB+P0W9z//+/ACEoutA5LlKILe8HJVtETE64FgsCqB3M5fDp7P5m
2hyfRJ7XMGKt6F34/5LFMxsIzV/+88QqtpkHKjp7lYI/5yYpQfpWa++QStZxpsGH
dBA+hs8Lx96oS7sfU6/7DiZpz5vHtPlvd6VsNyMuDjD4I4FQG871Hk8WSfgyVgpm
u1O40yfdzukP9f/mBkR1LRcMjizsGB5RncgDnQvmTvK59rPQdjzFEqmdCUGiIHb/
wUal9lVxNKXDcwsVwV4rRFF35mJdrU5FbeBbleCKXdT4tigcVqLI+dF/RIQ1+F5e
zD8gZz1RyIMH0XIvAFnFo1cssSM/rGkFz7ESVJMKQhvn13oSIyejaIIGc2cmgW5T
kbQYZV4Dka2a5mOjdy/igJw7YTyl1837QMH9/qZvDKYxZVB4PFrbDgtpczs2qgvq
r1tT1GexEIo94FuQ/OsCDpm0enOnu2JmOkgGBvlQtrT18dULUFgbazt/DHY3Tr83
a3KHtHgEhdkITTEdtd91nOGU4kcPet3pQ1kv2XNMpaDUNepSn5N/XoTIybdRWxdK
X1USzJcKBZmbKPtjilKsHxhhFIhIJqVaaJ0krmjG9lUvwbq7nURzXlFEsG7Ch+fy
vbTsb8Q3Ye0hfU4GXKZQiuotwAsmyhQLF9/OWeGCit89k0iOTavosh8nqy6fXzZk
VeO7zYi/EpJZG3o11WLgwg==
`protect END_PROTECTED
