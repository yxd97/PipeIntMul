`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7VdXmvfJLreaOeCea6dOPDDRCl3E/wdK+HQYop7f1Xjzfy+1ySs6wLAVIxiDRVi
o/p4q4GsQR3iAUJiYpBjDviNZZinXr0d/wjvL263tXDrnhHj3V+Q6iYvh+8Qe+0n
GS9JSXJv4PW321ZCdVA1rbXMjm5xHyVgdb8TNNggDhMO6Q4JjVZMr7KfTHqhtgwo
XHwwdyK8BJtsONeDoazJVwOSErAOAgLak/m7UZuzQ0/RhtQ8XDCWdxaczzP38kEe
BFLAYHzAQ2W0avvuxaDYiaQk+LD0ypBxsa1KH+X/1Mx6X2LMXrIvr/V2ULAwZNJD
j3sKlxkv+huNX8raH+i4UEtzqa8moxUi2F9FV0iENABR6hR1YFIUR6wQ4WrWjrON
o1zvisfKjWUrcUZIdbBUmF6zwDMwWCpUsxZnRwpb22/oi06+smIYo5i5BcE9STCO
`protect END_PROTECTED
