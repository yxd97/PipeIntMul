`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/hokJnevLYFHcQWmTUscQzGYtSdML/g8wVYK55VeIneVejnp6NM266M11qQHKjs
7KvjKnQFsW/JpLRv4nBCgzhksiuad/TrX8Dt09fiv5T8fWJM/oAhryR0TgK7J8aG
m3kOrLiOLLmcGBtwg7AqZhstPoOHUhJKoV0aEwR+jE4Mjhfb5nQCe1UBLdeC5XUM
z9PmSKZuoNpWQ8oelKplI9iEYdjJjmyChlF0tgVMUihu8yYLKouxclV7lYHdYNUV
rE6xU4k7hA2xxoCBFm3M4ZqIDziJtsLGOCobNorQGnxXhNeZfhTDlFvhNUmLRpcM
kwTPHE+HYgDsc0fGdOe2LTNkkz5Oe3ubcprQymbn9EnxxDy2I9kluNS+LWWma4Ll
ddyB8wfuoy0bv76qCgQ7JoDdy0YH5FdrJOeDnfEib69YsuO6xOsYBZpnFs+FvKRm
rIvdlhJYeVRrjeCnQFEcVjG+N18seQKlgSTGCvnwSIpzUoTOUZGBFy4YaK7lhyJY
`protect END_PROTECTED
