`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9RWqeZuPw2XI3njchHWQ+LbJeB2pbW0WcxEuGC1HPVswAaPBOqL4fp00onnymur
oDfJgHHpsqU3cYgk1Juxj76p5CClwLxJZfBDhhHzvFPU9Sfa4HCaHifqBndMN2YF
cCVoUXjsOjjxVL3xYi0gTZ+S2srwl7jHp2Y/fujGgpz05F8Vvg8eeySxM6m9c9xI
cB8z7gqsoKHRggK+tNmxBnMUYQfl79Muk/pgY++0wpfE0CrTXwMtp3aptQfHtw74
oaBQ9wdCHNnybG89cbIz2kyJX6RxJi0nHhTQ8+YOZ2eJaPQE/j1CbJFKm6akCtNl
lqv4fb5G0tS0zpotRZpg6g7AfohsJ1pXkQAjjc2VgjAiv+FkO4/FGEAardl3dDMs
JTOzy8vXO53pYH9i6gjHI4JUZc6fecnukLT0OGZKkuv9w8Qjf91O4FP4PrzMjrao
JeeLD1IILr1Xy6fFf4tj5+wKID1bT1TMsa7s8dx29IMZHyZ8Nt9JgeXgEiOX5cZS
rcxXSYSb0V9XFbbbA64zBfLsd555uHT6bzQgBrv6irvxd2tYwzFzhFaxnhkFsGUR
WPoVZ2rW/s0UX0udl8UXBZiIKmA1w9wfX2cLaV0SdiZhMiSvBtGfqGNc2IOKt4Qq
GC3PjAzGQzdeyRfQrcPuw3ij+ImyocVbj4Nj+A0wiBBpnXZPllup81hL5CmUyxlB
1DAFDz5+gLyv2m9yEqu2Rm/X/eCMpOG3B+CVKgU0/cc=
`protect END_PROTECTED
