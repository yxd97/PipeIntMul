`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LXOT/VQG7AsLu0SXkoFSII5hL0UfZmJYPpybP/DvQtgKvDK84z5iOwgdCFwOsNaV
Bg8lLxpq35CdGJ6Lffpn4o4pjjkBhQt7xcFSt7+ftVnLbrffMJyY7neVV9tuwbDQ
a3G/p1N/lun7CGGS8udRESpNPsA7Gd6Fw9dKTJnzIy9ksdZ9hMJTBKphXBcDNvb2
/qWhLLg/qqv81LcU4V9BJ6zneMMWectIEOiSrQ+gpjL61FyO1H1JFnL6xh1elcsg
pPsMVgdjbInJh/9gY7gtgMn7aI99SPMMV0qdBRVYVQlIe9PfR7+2DEzSQQWK86PN
ig7e8egLXUGxznZowYHnM5QR+K7DisthyoieAVeSDCzeiRF5diMwEOo21m7bHMHp
IXgM9bXCFC0gIzN8A8MREQ==
`protect END_PROTECTED
