`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfVYEEdqWPpvdCL3deAgxht7eAOlinfgX5e32EEBZp34myeyZiyAX7WNrpbR7Gdq
JonJQmY7ZBOdf56Wmq6DdMf1DkuOxuMRPyjo4OprkDHAkxEeOb+VKmiK2vd7Q9BG
YXLMqlXYxy1kLI6OavIWrD0KJSJ/klIPMjnUIjrx0pX9mOESRQ+ubA/0iHYu+njR
rq2QzvK6lY/h/WAMwUwqwZQurmTd+G5iyK3Uur9a2rboaLc6QPmvfiEEx37hCosV
FOZRMSTaBe+uyaNrIvcw6bWXhfr99h6fAOWuX7x0U38Og/9fCH2rN7KI/OB/e8LK
+sUS65L/DK9sbSJ/pUFZ+NZDZIVXgy4gy9AsKK0SF7wMILLCGw5JIXsQdcQrDB2l
ZHQqOQ+DHQSeKcgWDNwSQw8ov2aCx816Q+ZosC7TRyjPrAsKKPJ0Aws6CCPCSRaN
`protect END_PROTECTED
