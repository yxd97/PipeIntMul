`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbBDgnxj5M8HeFYS/IbgFSlKJdIo3fKsz6xkAUw7de67len0ZL6un8rnJtb0F4Sa
aEOKkz9LywNuMTJKGQhPfNcp6WVpWs6uReMLM3mp5KBlvxWkOjHSgDYxR0M8IbCX
iSmB/TqLhxjbnOn1zcED3/agh0IRuTiOdOZUj8EK7EQI2fLe3g65bjRvvKEdrxkc
kOiI3GgcyQrW+0C9FPp+oTrl++m6FwgJ1BV02d2W9NxDEn6AagRawofaBJv4TU1V
CYDvQSPWJYpBYK/DLzf8vEPXoM2b+tyYS8qXx1kzZVHClfiuAKeYB7mLcNxW5nxv
QStXrGpiLpLUpROfowVT0qFgu7K3jIcLMP+paaZEVk2dijYPRYic5XlGsU7/YHhO
mtwn7eNh7GEdt1Pec418Hg==
`protect END_PROTECTED
