`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0AQdDyNrY/UW2AS2aWMpE/Tv9Cx3FHkt2/nziimtYleHVp+viq2wRthudSY7sjtm
DA9gkhZpkHChpnOjEGRC1q/YtXV/XFQOR/H+QwkeJ2F27Iece55Fe2o+n8DSAJKM
8hDN08QbsyK67Re3ZzM1LoXZ0DmoJ3fLc+IWBfMQdkMBKeXrDcZ08fOQ4+cr0y6Y
0O2XbqaTtKpl+kD7lhfEHfm5M7aGcyy2VvRALbi89mf4JRZX1R84OqBMPQYhaE+N
NCsR6YSHdzqFyhOlZICKddfOUUnDWr9y8iKG7yshf00MKEPON3gX94NYlcb5x6te
tH5Y3+lwZV6CLVtOZb0+rNpAzWEkkapwItSCtlTb/sgeVXILiMJ3wT3F22ImQduA
sxTFS541xtzriRAkpF9er85/KanXgbsHBHoheQO/WS/+xg1gw3zRypockS3zYj5S
ITL03WfhhLJYgLMJpFMaJWg7FaWarb6XgI9RqC/X+qfUcW98EWyOpCfkpQEYhfBb
rWcO5NsbfniPOKFleRLM6tSKXCTHDqpGnZWM2tJ/+3t8/kiIw1+ie1wtQ6oez8Q5
C3AaN/9vxgEew6aGpwFNIBujSc5sAF0DX71lgIrv61NBjamELypOv1oWLdkhW08Y
6D2TbViPmtyPZDMiYBS4W5a591TG3zJKmpEiT+J/CjunLCtadm0Swj6sqfTHu6dW
axU6jgTOB5Q/bD51c+qibg==
`protect END_PROTECTED
