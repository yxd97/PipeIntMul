`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w15wa6LC/fAIwd/9kA6erBu8gsY+NG/v4wAJMdkY8YFwrx8IJv9x44pa8+6WoRx7
wIu94hHwouZMkV0uPjhVg7lLUFTtUt6sCOlOiFE9mobobI0Y2XzPo7AnL5PsX0FK
CpgeMa5UH+EQ/9OquAI4ZVmrMQNbEzM/JrdTDVAC+rI8m9Ri0L5lwAPGRSLJW2Xb
qbEis3lWeuJsUzBb9RQx/xVV9GxYZb/+w1O7fe0h/nEe7QTg9E05vlWH64ppT34s
BHTUSWM6U1sgRXCGpZOdr5axKwUMoFr/DmlrpsqGt1tR8t1ge3cgJ88j4/LqrWT2
dyzMOwQg2ybabA300926oxqEp8WR9qUHh/F9eXhecAfG89JDlieiwASx6GCgVAkW
IUvWNZcrfIlVhgZzRBP4OZvUMwyY4b9rzu9mUXrW2Mec+rvefOjYW0319blaiVMu
Fqzv02jCBCi43an2SmTMWJIEoKFm9qZbMdMOduz2TiCx+MRjJIcDC4oySjfEPSci
zyigZX9+w3YMFZMfbQBYRLjJGkJdhQIvhebNQGuXzy+5uBLHdTv5AsE8eWOchyIt
veHgcFvymx9IHEYQHArjRq2AYY7mSTjNeopejXjBfvmMtTzUncIMVn1QUXnSo7k+
InuEpRtX5DLahtl1bcUVfbVf0Fc+SwaXfKL06UnPOutMoCerWoLea2FoR0pJI6/r
nC6vIDJyHZ6SqRcheBSMR9+iwcRM78yFsGFb9QH3NIItqlmo4qNAykBd3z7pET7m
WtV3jHe8TcSo/ZYv3nzofvuetutRTv4/33ivvkResdkyB/JacL7wUzIZLs6Qeucg
sv3ezFckT++ZRy7KGW2Hmdd476FO7fjtn5OAgpysDhlVgnszA9Z6X3mZHVAar065
`protect END_PROTECTED
