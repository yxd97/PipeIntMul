`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rGJVpFuU+eDsbfXWFXvE8UwaqsNbZuIUHk46CmZMUL7jSuqSDLRhGkbyACoAnINN
V5Sj8Yjw8MdrlfEHc2b5QcruKrURJb0IwuCnqloV6Fx+eVi5iisDJUVucpOf0uP+
FG1AjJSv5kw38PxVfJ++yufePcKbRVLtV9KR/cc/wDs2GWfjs8a2uYB4fvOtNmUp
OcJGsTquWQm+q1VadxFEBkDk0ab3NH2vzZxEH8L5zvNBrnN8z9yzuhYPP8jzvF8A
A558L5tAJJ22m8OkSDkX99iuIg83DLJz6qT5PrSm0Clii/DYXhRvE4ymLliySQAQ
bSQRAUR1Bb8N0ERLTaGn5lBJEWbYPL2Vw4rAovSHHrT1Q+/Ndrz+W7w//6h+TrSt
6MGQE7dR4l/g/Ds52415vKkgNgbAGjQ4mwUMDocyOcC2GVT0uEJYVUAam3OZTQGz
jfqrZLUcCJbe2JH+b2K23Y+9yrE386MKH9A8zlIOvxbYUaP5cPgJY5J0/HG4fXtE
e/4tR31HOXayt8kO8kLtOLPikKntfZzvXmVHALchXaB8T6mugIfDOCWdLWeE3uID
a2p2YqBBIoyK6asvuFPdSB7QMVBfPP+UJkweCT9QTfztl2ZoZx9BPvkHp3P047As
rLFlZA1tbuL4hEpEctYHvlhIe4eBl44GjEagvVXr5EvWuuhnNJT4UBGlwEf2eXQP
kyV9AnrVBNj2NQhwwsNps+pQ6YNkA1GLG5WapaNi5QWdiWknu4HJFCCP8OGkG1HF
o6Toqr+lymlYXhAoRZCjsxiDb0imvONH8sr6DCIPFfTkgyNkNbfv7D1iz+R1f1LZ
UEkC3fD4MNnjcZfSb9GlNpMhK2aMmtgpIMaiqHwI09SJnZuJeECehL7mDWIY/cyE
M+lWDNVYWxUJfDPZGVEhDKP2pHGjjPDbe53t3vfOv8ma2/FUTuql1gZxCUnpqwIY
+lINiKWqM/h3IPRJYtarh2pnBegFMdXCRjdmi4rkW0P4yk8imezryiPA5sc8hWMF
Mo2O7BP4/ubKa0/fPxB/zJSgXlEfMYa36Gip7v6rDfoJNJ37yjvAbJFs8/0Yxkcw
fLBVPk6Ybd2Y1JDeA4m6cq9W7JecJdeXRmzSpjny9URupMfR8TPRKgsIeQZ8lk4d
gz66BSYvai1icpaBH9ROdCnqI3toOl3qxTuh1E9Bs2ypygRJ54xC5yJSZGp8Ml7l
SswUyO8QDSGdF/tEHeTHtjB7Kh9VY+1olGmY9B9UfCxlaX3Nd2059vyiokJHTFyV
jJlb3qr/ROM8i+nmP/ZVzb1pYP1/hneWy3Q3KGQG5ibKbNnwVb3vPWRgrgd01yNS
7eknTOpx2UgXuX85fgSemXTeatqTmU8DcFF8TE46EVuwCzq0glhx0yQFSJVOkyDX
s2gk9oykU/SWWcR0TVEOd0vjkyy/7EQitPhSahWFjWPGWEl5NzMWSSMO8bHYuZ4j
VKb9/d1cHdJiDav3zeHgiC6DSrQbfnYMYvCx/pHk9lo=
`protect END_PROTECTED
