`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sd9luc2MX/NDfVt0jN1lazM6oH5Ud67OfwWotPEyjyqKmDp3RTirmurljer05msr
M+ruPFtOXUVssMr9xBmEh0sddgi63sFDo0h6YujD30GUkJO7Yb4Rvqy4gFJ9gtSr
u3nVao4gXTz8yDOKho+dLTmHz76LVHx+E5PNJmz234l2zNO6VdPuQ3cHaAsByuhG
AY3czv7HAKMMGAtt+rc38gT74F8SUq3PXCFm/Mj8AYDpTsMeCEIIgW5Mx7oRkVoj
U3OU9Y5Hv/mysso9beCn+6LEVZgKkKBPQukaWGnR2i/zz02lu9NO1vwkp3HidAUu
56JrRIAWa+2ZDbbP4vBXzHTD/3KVqiPYt/WCvTlr5iumXEAtZUDCY/6H+fAfOB6H
2E+mFaPx0IBuSAv210fnLtXFJWjxrpEkQs1hxvz4rZ/6nCRBaNTHoePGtXZaJLUg
ilJG47PERYdcfBOgaSjphKceTYWplii4JmAj1zKllufZ3Y2xbs/xC0YrhW5ISYNX
BOauvdXn4kumROTd5p9+OhlgLBF4NEKpRkckKSKXXFYSykE799QkTsLnIdUZkxFN
EdwX2t3KB80w5mlXQ9I8j4E9DPROAdC9jlbDeVmqwsoPmBQ7kwH1AQGO1HxAlkOx
smnwE+EX0vdwv6vYrRguC/cKekZzDA7wlhM/bxubX7OflPmLxZmud18Yf+M2/bTT
e9j12b1aTee7q9Ek+f5iHbGY5uzah/8LL4zyauBfAdFbhcfBbpdipVilp9vH4XD6
qpA5lefRjGWXp0bwlr762f+buoWg6ECJhWNCVU4mvfzwkc01XQ0EtRR2FpbPfTRi
zLztifVkC9r78x0xuhDCQWa5jtl1F9EwfmUSnJGGRQCKte40k1vA+I1tjW04usKw
06JzefKM3BBZfPtzABvZTTDVwypMx8ji7wK+g9OTezw///6S4+FF0l3y+rwxusIS
Sd+Ro6lhQJ+AWQ5ECxMovN2sNO0f12ouKSMwwa+zdDjEHGcNtI4T7eZIAlgMZi+K
wocmezZzTZT8EF9LJp1yNcHL98V1EsSnuOvs+FWbi5TuHN3BLUXzwm8LlX0Qzs7U
KYDQlpP43yZDtLLHeBiu0HiqHXntxmj+B82nRVg5vKTuzFrgNw1m5+JQ1//6sBj0
AnRXhQauc6X91IQaXmSklLrP0XNEgxcZZYcGZ3DWaB733VPN3cMCRchU8oueppBe
kEnDyD5b3kmh/fi2z1nqAV2xc7UQvdm5U7Zja3JmfaYqEDSYQqlOZPQWHPBokyLA
NBtRXVkOp6WPkIEamFPz7MpEhdYOMvBoTY9TSMjDcKUfMND5T4Jh73OOIrHDUoRy
OPPoS6FrFoTh1bgF6hDtqbPjGBN1Y9CgSS11vHkK5AZz3qUw0mUk7ztgWBMW1clc
`protect END_PROTECTED
