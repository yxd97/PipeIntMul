`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDydJHo9SMtYHCdnjDJt1VDzkrOMGgvXeZk4OuvwnfyPn0+Or4AEZQhuK6FUnaaL
3Rjk3P8FtZuYzjFHeJsIwuvahTHMi04fN3Iye3lBZ7PZzeQIJW2ddrHYdWzk1dzD
JSNJjDp1MQuhFaj4xyteEt5S1a39WseUWnD0gzl78S1fx8wD2vC4H2BPzaPfB1jW
6Mf6fjmz248XM+NULb54PibdMILXT48BlCf2TXefgbCupRO3PJ1rdk4bCuVoclDI
5ldXBiEAk15NRunFxWX+ggQpiAgZuI6ske9kTwdKEvh4qUUavv1KmQ4b+JP3aV7E
WISnHIpdeVMsX42GA/njGUBUIpW2fB+3f2Kz3L3af/7Uit7ehj0ygx57QiWGgssz
hVpOi+/aZhPQLHh7vGiI6WUtjEQAQM+ho1b5wvSNJ5SKvi8SSUHE/7TudwP824AS
xQenBBxM4rLNBMAfwysdHGH/IfGUaMUlhGWa9+li5RZKm3mmpacA9oGLwOC80byH
FhwhsHjDkZa4J3wFmeMv1jW5hR7SDecxVVHl4LDLTvVgRO3i+1TBKVKtLIWqoCv5
BDt2Ok42yizgfj6d57wTY3xjVR8xnUdE9ccNGzyG901YY7+X0bmgrKnykzZ8lrIu
/lJnx9HecnDYmSCR6Y+8zw==
`protect END_PROTECTED
