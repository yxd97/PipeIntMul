`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pi1XJSVaOZmX7rlyamu549lzNXufWDRtFpEcnOjJOaQgCKvoSlxgv7DHiu6M2/eu
3xsenWNiu0bfdpGu9eEWpNMLmP20kY0XYSSSvXKGeJUYYAIX5g9qzs512+2gSQfg
sv6cdCNXHglxx8wShBBWaGeagKBv44CTNqp5Md5z0+2+BFmQegKthETROsmFaZTx
5vgLHDRLZTCDTLxfFo/Rf92gY6MTRCCArXs83Th4U9ODN/xu3as6oI2yVy4NidET
skBkMd07ADAgfVuP4xS+A8ksTWqE99JfcarjjQEL3g8Vjue101UWGomCS5CtcLvC
GtnV48wGC65IuWK6P0/EyLGiGE8QiBHT509GPeSoKvV+vo9Zxs7kPW38z4ok1sT+
jK0vvAkPs+dFx6dT9aYqNQ==
`protect END_PROTECTED
