`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmNRvY6KdWdMeoP30ClsE5IBDrNGD95mPh+QUk6xXl+zDDXT1mFMFO5ZZXGX3kvP
/sQFi8lvP7HnBajPmQVxP/pYCnyc+oZNqlaf2JIju09DRGLPOr63L5oqqucBdFEV
0vLI3ZLAkhOp0tBU9TmRMD+Cr1oAz0k/zBBIOTKi4Eqzg6T6fVaiZqTy3Dkb5BU1
Oo9SHy8e91Y6tkH2k+M+/UFl9doJTVYd+WMe5qxEYhj669yi0dMk224vo6fG+4oM
aq6NBXVSKSxOclxWhFVVFvYzcsjtYwdPl23CofySH2ECmGFnpaMLJKQp/W/b6brG
JdC6sVhTmuoWxAO2U5oN02P6MbARHlGFMxHCkFUMWMgLTLg50mZ7U1ZIsP+uzq4V
gMd2kuGJTY5PxX64KV0PfvvPqQOPbgY9iuXW2lcblTaFWiuO5Y8ju3ioLWQw4IjE
4iy8kmUZtgJ1uvq13xjry2G4zYKIszkjWbO5z4vhwCCJX3VEPgSRyXXlpK6vIFmD
LAf3+C5WOttSB17Xh0+v1Wh+mn8qUStkUG063m2TOh4t7QK15AI55HsNMIDJVgPu
P+RE8TD3QI6aUT/qX6a9lLcWUMd/2O3dX3n6ZJaG7Y1ZDBjfhwddHo7Lle5IZBpE
YrVgt258Fdk1SBdHbtgduw==
`protect END_PROTECTED
