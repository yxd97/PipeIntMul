`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHaiPbO4/tN98cxLnRoT0BSYTJ4mgibbfwm5Fb87VVJCvILC/LM0ZXwn9lPb+x0B
OnYnu/Bol5raE47ejZcnMz4476WV7SuNyBN+sam3Sr05SBcV3zlYrkv1XBLHdMCZ
84bifymHcYyjeJCkcKe1D/zw1GtEzBjnegSW4iOt4AvVABLSm51l5qNgdDeljvPK
WEyHCOfUWeGwUhrXivVQRvd4QVQM5/e3UuQ9g7HiWKWAN5Bs4A6rd3Sn45N/CuYy
y4nr0HXyEJYDScMBOOipnEXAQG5R82V/6j86mFysY4+2aAxaq89A+X1t2OH+HbZ6
zEMpLciSFhp81RS6eNYZx7DlWUBYG0kBsjzdN24k8bLRgocqCqD2yhmNnjR7AISX
RFcJNPdfXp4q6Ftpbj1YSLKkalRGSsxZ+cZ2zDs1msPZiwA/gyBed0m3IFVeaTdJ
qZNLP3/4H5PvYd8XkcSgPU/sXF30ZTD6B4MJp7WJAsh/WglxdUHvLF5x/Jx2Eg5G
`protect END_PROTECTED
