`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sLB789NaEKGaEGiNkyhrHRp6bvIEOR9fgA7UF50yVCI1vagCHoEGzCJ8unftoRnv
PuZV69p1alD6CDvT0ZtEzkysUfZ09j8Izh+1rRh3EMw/fQviRrsu+1YPdcNBlf4z
Qfv0WO8myAFSYW7OKBJ8qI9m0234uDVXyS0B6XEMl8JlCM5igcfg/C2kb5WQS7Jv
g5kPM/EVndi0BIbi+JPFAB8323UpRJG5PCNwAxvKfMWcGEjVmLsQlzWDNipdPMzW
W9Az963Ry2qhl4TNgrOqBm00vBcSerKYb6gsfOhm6APA7ZLe48hesUpyZZrHLkVM
AJNFDWZiou4bl2y7NWXv4TF2fqssPPZps2kLqmXXfOngQRCfW8VZE99M0CJsvC+M
Cl/lDSb/PE1HhphTgtVo/QNiWhDw8pBbCSMW9gmJ3dk=
`protect END_PROTECTED
