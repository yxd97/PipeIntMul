`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ydxf3zu+OnDDpW850CrkJlEyWK5pnkgUT9/s1tbfJBdny9MA9YvpF+/dkXm7DxYC
XwFJchDKs2KtVFonwWQjMEdOwnWZv3IQJ41NEx4qbkGZ8/U4N+kc4N+3wxEVWzaj
WF3mYbHU3nm2F0r47oZxdnsOpnWcBd5h24aWEBgIYbMFuYUVRivdxs8qFdsHaJqA
KLthc8UTW/BdoesuCaIF7HzlmwtAt5YtrItmBupbBC0J7rveN4F9H/v5gGsG/sTN
Gx/2G79mxf5q/VNFkpPbWKnw+i0sLBYTz8gV70gS0X3FyhAs1SXALT6rZSiGiAgo
`protect END_PROTECTED
