`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHznP95PpWCqIHv6b78sxBpiHsRAB3FJ1ZvY45l8j2ylxfyBr9lMis4fvjsSzfF0
vy8ydjWnotjQNDChblyIa3ICSgtOc5qvY8O75lLTJybN4hv3VTTh1ieB2nrdm4ad
8Q7uSu0UiRzf4ZvQTpNnW7GrXXErIw7Q46D4yNHtz8+ymxK0A5gLf6susdmawWUN
7KJ18LMsoWLscyaPqT0OvFTof1xN6qJ0aXdyx/sZX0ODgD77AAPdTdIBFMBVhJC0
vdLgz3TU1zfs8Av7kjtjNLc+55d54U05YTgXEKoht982NVosHi5P8nDqBGHeoS1A
syhrs2FUafSLSC6oioZ0jA==
`protect END_PROTECTED
