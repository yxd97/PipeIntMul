`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Whas99x+jb4iga4Zgy5Rx8nTm2pM2/YP3DJEAlm2D7ltekDwaKc0YN4hJZ8SR9M
SjqPKIz8drektGThaPDB8GdXJLLcgrxeWXwN7iFsjAtlodLFuQ/yfsFX3yB5JxYm
rtlQQjW1y7HqUohTt/n1xhmhhJr27bmigc0zwpCFtB+ZLPa4qFwR4F+zLYCQbjlq
zxC1AtQkOcBZdr9mV94qTZvbUAzlMBU1eLhIn0o995wu/08c0kjjBuULe7XJgan4
AJrt7ksqraGlXFTbxWbGnTZk2/ZLbsZyMPVwsSIwu40=
`protect END_PROTECTED
