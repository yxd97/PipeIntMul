`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Mmv7hN9JIKM1hKibodF1f9QEQwovWbCqj9vJLh9dQek/FD3J2BswmqY0ap4+o8S
dP+2mLbvMFhN0oKvAOC2loIFICPOV6Pyu0c7z3pSMdJjM+k1/VQimZS5coCsGFIt
rmYUlUoy1mxufYfjiA2/q2kfmZQJfrXIJCB3YDWM/1RYdky7S3jYg2OqrOQRkKNf
QEU4GBlufg+DTEF+C5GkDQoxIxULnp8OBGWb+d4dxl6StMiUWp9d5kSlFMG1lKwt
wXEXgi/Rl9KYvOLiA/aAI0nCaMHaF0f7xG6HiwpuJC3VhsACp9uiMV8pcwzVita2
mgHdfdZxHCkltStHjTPJvQ+w825mHS6C5LzqFcVlCd8MzPCfZRXcO4WWiBnlNTFA
o0m0wsIZzyrjDhWAJhL8vn+c1sHqzNhcikpWHav2Dn8vxZgNe75ugUa8LajXxDw3
8/Jli4M7dvweT2Q4JwiNOp+cDvPJKeMp0sdrhCvIcyx/ghud6W5666pqPqrMyFkr
KfwcVriw0U6HfQWQ+S7QMoXRnmQ6BDOWFcQVykhiXjbdGzlbSd7eD1w06ZBNSWHj
Re5U2nJitpQye1NeLBJ0O81VHC5rPSOFFzQ116Nzx0UygFgeGONM3RNZIlc+7a1M
feCBhmfFuqJ6osDXyt79T6ZWdH+OC+L2OpWg0aRf/k0=
`protect END_PROTECTED
