`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JnmfcPwYBpdilAhE8fs/SkqtyVdcWXL6Rs1mzb2PwsHlRc/765KmF4F2hwBJudvL
93B8RGmgptFD4WjF69UCtYeEiYDDGSVJ5uL6WKPg+5CPSMw4muh939DyUTufWFjg
8BZScMmM3QN5hCEzd/gLeO/n4zEqHkLVEADMB+hL5fA66SHJmIK8OJdScII8Fuak
wLLCR/5kEzpJti4fKYSugD3mCV3MWJuZtQNijn9AAlEBue0bTnUACce0RaRRHPSI
lIcYi8/6DBxe12uqNEJ4nfVGp1jdEcBt4QfmcBust/GTLKSwzUgoUC6eE5Q2OtXv
hXxKKTj5gz5ZkUr1VrO3vZmQzEh2Q+lLEqCh10yjNeAruTOC5QSDEV6QrAU3FQcI
jGm+ItPnOPGaY25vSOf6jRz5mICpChOzx19kVUufAvcfspQUVBfuB3rpT4RTquqC
MB/pFcUcKZVswL87OHemUYh+c/n8ykBmtaY5KqxsZAjT/A9QsN2JHrzIf6I/mGme
FyE6IjdVodhRsBPzhXMnmIrvABw4nuYzPT28hN+PAtviNWOqgWkgqcuvdNccBNIn
/8JK01KA39zAzUJ6XOq9jimsX95ykgtYYP8CXBwxxeCye52yxSS0C85chiKXhDFk
gHlRY78sA8tGu5oGArPzj49j2Kw5/VwZmE654PY6KyowtiHT+a6NGK4ibdv9YqP+
qxlnO4cHZeK1av+40lEzsUZnpwZay8x9aZ3K5iFEx4b7JV/TFU8hU5aZuLGy2vL/
ddktZ8nRVgS7k8vfzYpAW6BGyDoqiWOYGfEnJ7mfSGHEaPUR8Ic88YpKorCkQ+3h
ICYxkqN8HHJgx7NsQJS4TwtG60LpQid5qtEZXjeruixjZPdqVXO+GJGhyUuS9vRI
YydCdsfZD/5lWPGqPqy79Q==
`protect END_PROTECTED
