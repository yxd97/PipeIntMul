`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LP6ryqmpnggOhkWetd9dbjarag29vF4v/KzCTlSHcSwi25WzWZqBr2bM/wfxyx1e
j+xOJwW6S551BOEtpy2326XuuDpMjBPS3CWHf5exfRgSAD8U8OtZWP3WzLxbr1IU
pWpoazGZ+UlR9AZCH5gOeTgBPiaN0DdAPCeO0Zu63QMUOmY63ezHK5GNqKoGPysl
cfObzblL/qSuyD3dQmYFt/G+z6YhqccJ6QHFjapweuWuOhmLwOCv7s7p3/rwJIZs
ARHFgCatRLil9VWCB7zQbIrYVpkGc1jpMqymRe62HOaa0HLymqFLSCay2CZrGGKu
YqSKhxECyXUDjR5E2MCd5wzw0fgnbnMJf0wuLsWT3n7PWXU6+ZsuJL8+AxhrddkZ
1jIbQr1DUHqMHZgwtp3UioSZ07R8XPogEaMxZqHKu03t0XTk9+ol+v7zrWU9Q3x5
QOEG2AyOMGDNlcrCe8AzpA3KQQmXSgJ2TwsV41xOugMgZtsXJrvpojOnpkDRbYDB
0E4Il1P6xaq4VEW7lUS8NMCIsXdMkH4PKduUkQGhXNe5HeBbaupByvJAbtRJehD0
JFxPJUQxKOnEMr1XA4hK7aR+mD1/DF2YkZci7HuAI9NUEjz+C0F4KjvmPnLmkuc4
KxzB6gXBSsKsSRqOCU6f4nXVsIAKOcnpjdzPl1dNhQXpZMwZFU/2ZrFfqdCJOKU9
yMnEJtxwbbQR0T0Jdn/KvMNzCX2WE9W6JKPAxio0YOTn68tLNDr2zM6YKr7ZouP8
aBd329mHqtCXuX2izdIlqwgZNSsWLfn9Ix9gfmA3r6t7qLvSrAKQ+i+z9L9YCEBN
5SEeLGLKdQO9OSc3GZ22nohsgWeVKHMVHUqQR+kB9enn6S4/W4CtffNUzmeH1Wqw
DuVkTL17VqGJb6mi74wEHr9YKmeDajLwlNLjc3/meaM+JcBBBXucLOV8oFoLCuby
jHUVyRkm5MToX/PXMij0t4mk7yRhvs8XXlptlrKwgQU=
`protect END_PROTECTED
