`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dO7WOrGKQy26ttG1nJ0V2ss4IA5x41vXg9Jqp1Pz5CjBJNdZhXQIDidwVcgR1yby
EIOsGBEUdzdBRlZuc5mGGfmV5mcxadjcVzQ6OijnKkjHDBFb599pPdu8iqoPOdhg
tBxmhmKEtcp+KNlFPVJOzHuwB7P+p5BDt/NBuvmlB0fl7x79CGnQeY5JO2FFSvJG
MeGRHridqRQ+J/SIeNciI9RMZmlXwof4CSrWZQ2VcWXAHaIYF1aSEzhavKeGj8P6
Buft9dUK0c2r+CfIFVLzkg==
`protect END_PROTECTED
