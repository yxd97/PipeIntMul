`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nX8h3jww1hzZJHRP5FSemOTRr/zIUdWr9s066fKt4Y+9Dw6f1lOPpb9Y2r24SvpI
B8LsWXjhBI20kLLtg/eSNZpIUqcn//tsKuT93mOABr8EuXymL19kX255Zj+pHIJv
0ALAeT9Vee3XW9qORZOAy2RUAoIP1IQgaynlWp9Y5MmSeYjHDgOPZCZHSdSpXszy
ZifIhvpRxHnezus02Vw2QIwUCubJ+C268lEhSXS0M+zSjKMjFopHlRMs8zJCPs1u
bYowS2ayJMHoC7qJY4zTExlX5Z0qp0voH5OzfOsSFuyUKc0Cy2TIFXoMdbNmPoOD
GBBuKByDYnsJW9RjLS2CUK6gCw8Dr3R/vdsubXGt2rZrrs+acPfiWQH2NNU3JwrF
2TVM8+oZ/eBmppNQLZnndVQ0HrBGTbf0fySc6K7xEsU=
`protect END_PROTECTED
