`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXDPZ+E1bufFbbBbtxOnP7IxNh/54isJlEwNkblsKHfzhVI3JLZgotYvklEVFX1j
Ma04xdSzkHoyZ4pryeyp3npbzwI4YUcSb0ppdvTcuMVixN3AW8qwMjrgVtWMeyd6
BIILZ13f9G/bAkqhPrLZ71d/0C5GoMI8YQEpDXErnxk4CWiSRKNQ1CglV+d+DwNl
VNgIfWFXMXnfYcIsxGR018er9GdyZzR+ToZ5iHf2XqTxfyUL4UjkM+Cmx+N+Pmpc
cJW38IRDhla5rZl1LIV5sb6XPaNP6VASqCNk7yyHJ848CE7EGmokkWqb6gUP4kAB
gbFG1u5NL8/yARlVD/251eP9Dfr21NZ0Da4Nuvrp1dslfhmj0wOXdSrohILSrHDY
`protect END_PROTECTED
