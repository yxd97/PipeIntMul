`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VI5mTa0Z4Vo+JmbFoAsD5VXGJetWmMtiQlMjnr15VigeW/UwQWoVb2ArHJzPcv+Y
jHsLesgZoGTkr8FwgtNjyojyTUZXhEYTDDtw/RgSuGi6dS/3R7bHSdv7yOu25B01
7VmDIFcF7GUy7rcT9VCwvvarM0LiJNOqOXCJCpr5K52+sWx0Yj3hZHD+gu3VTMNe
QQfAfUGXD6zzLiuzb57ys0Bq1I3LmCQKu5kfoFGU6+iWmUfSz4EY2PR0Mi16qX9l
l/+7RZzcYbmHLGBHlTs7KKAJwVpAoJSsjDOA3EqjIlW1ZgWd7LatQ58MY9ggkC+B
KehOsD+c8qbJamy72WCRhJ+3ypwhElARYPLjzf4nCBoOzuoiiL4uD1p4qpES8+ZA
uzhWFCvKfy2yJVRj6buc2ohKxRKbx9hwaGsziMe/9LV797ue+J3VjngBTBz6uhFL
i0VRMPhMLf1bvrwIcONPzHdCy1HbEATZ6qRIBvoiRijCMUxwug8dUmT/uHXlfgJF
JPuS0ynzg2bLA3TtA8NGBOeYkL8yhKIcxKmd2KB1YCXuWUyX5jyMcwoLuHbBXOd4
3nUrmA4BQZu58j9TU/YQfBNr0s8CauXEXaOvgVfRNci4X30TMd7OWHqYqkK5o/kb
0e0ajdgzDDqVPEn9x6gCpw==
`protect END_PROTECTED
