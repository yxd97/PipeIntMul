`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYwEM2dnf4D/1/MZzEkcPiE/49zXg5+6hq/sZHe2Az+D4p7Z3EYbHmWy59oHSaCF
ZDZYbEOuVBBUFQBiwn1xSrpiwLcUyU2uHRXjPqDOTVRhgS4mrDXyHH5dAxVjB2qP
iPzOPeF3NmbjiFKDUe3PBIgGeSKuDiml194SIe7xeevvkfZSfqL2lXjFowlQK6cN
GnmxDsex3oM0XUs/XQJ3XJtLOz4KmJXCoSFwjiHWfHhQ6w7c4q1HCzR6xeHgofnU
DfC4mtUS1/0YCxy1HkuQUTLc0uamPF0vzdeCAEqAZvjx8SYtktbI+wDIyAj9bDd7
IgzvWgAZaKHaQgoxH/2pTLLJI4ZsxPl76AiXtuZufyqmDkqT3KCm1qjidAiGl+Vi
XbWqjcakVi38h8yyotj7ALYZf/SyOCLAxVGZK4iPVs61eB1IDROwZVks6JoYgk9l
l2dbLAWNicUBbLDHlU4EJq361sKLHDjRsFJprgw5mvnC5SFjLtPbmtTMpug7plo0
mcntKZG06mRsFT7iTuohCagv1k9zqY28yO1KnMjziL0TOJ7fIGaLohzxmGcoHDD7
2J05qKJLMLeXTe9z+HcS+6xDLezXgrBBfC1GGsM+NeLnlpoqYJwDCwdZAxnjS+SW
xykjYkRyTnyhwGioej0O98XzYUPJKTHa368UBTLNkPryGOdPEU6TMWgNNg3uisPi
v79MtXVSlUBJLcK76N2sAs1EOze/4JxEz17FKMnAmYIkZF+uUwfMnXrJF/F1keKv
WiHGeFYkJqE+vWBNB5ABy7gg1J5qWxgKeiKNhbPFE6VAxO6eDaW8uJ9SBcarv7yQ
wL3YDlLxNZDX1+jxuce+KUntPe4pQoKhkZ8j98g/GDZyKtiu73JM3rtaRDZMN7s1
NOSMpPs5hetkMCE6g5ihZdgHSVsKKUyhnMF2cRq01gwgPXDe6HqCjcXmwmnfqkGF
oJQ5sTcLOe0uz8kr06WKTp7DeSx3EijHPH0PiE74ARzfFP9fpLHtUwy8Bp1Tbzcr
110RAXxYhH3SZUe8AYeHNC+iCZ20fHC4jROoN0Rz/RZpVd0Z59v7EPf75ik1eGvK
8hVBfX7XltKUo20baFjCJtgmW3vLq7nRc8EqU8/s1ZKy45rW0Bd8zxWP9Ffi+5la
etVGRp4QVmOLhIrNfV+IMqxwMw7/E5/5N3QpxyvnxUWOOG795hfSrnsa5yV06sL8
POX9r9TQQDUJdCoFGqIa1g0M9mVjrab1Ci1T4F0SaSwbw5pTW3lEN6CBbUNQne5l
PbHDIax7/8RL9S59bD+NgKUZqngeahFAFyuEhP+heQbtqXkyFv4dwgVtTn13BQwr
H1kiEO1TuPrudjfFD9+tHNjOZcvnFBoItBBgZJTEgt+64vHGS4DN4R/TEM7+RKdP
Gx8EpjUczxGZtMY/i557j+VInsa/dEVtYSq1V1VlCJQ=
`protect END_PROTECTED
