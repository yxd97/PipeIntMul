`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1B1hWmF1ucf70D0zESw9YhWW6HPCDsgFUgK5d5d0Bua5c9up0KzKYZzI04WJQT6q
Hftw6+nqLqIQq7u0OLjhk64gmPsoXlxysM3QWS9r9u9gVZc35fj13nJ0wOfriqcG
GMykxJQLH/IHRWX43CxkTphy6Al89tqeKGB56u1UWfYZ1u3dseWdJyHucGsATOQX
jeRlIEwIpSIV0ZuTfWqhbOsuOu7hPpqWchNFSKaGBeSU04uzWbRZXM+x1eiKEXGS
wxXx7bzFvoHpUf2aI4flZMDxKRz+SDiHFaiwz54f3avznPyBOPftpPyAD0ymXV8i
2+msBfABKN36vjlGTVkgZUtSOCzpfXNNOxkMSplWz7axnC1vR60rNe0APP4K4tZP
dPgKkqkOP8oLd7HozoKK5DoCuWuwsIvI6eCZ0YMabxxx3PE0kmZvMdBohVL3PXT5
kOcOM5Cf0/JUFn3wB9i1ONugoHpo+dHhupk1whNz7+aX74Ws/Hjb4cbAcar5F5NZ
H88orw5jlP9SyPog8BkqmioifXasrjby1E8i2Qr3R+Sa+TCz2S7Hd5OHnaQstC42
l2kuGIE6Owem03Nm0iSpGFKk8sxS/7o3kfLwe10rxC/BY/y22lVmyr5vhsmISJ6Z
ottlMYGFY8d8Pll+6Axyhwrt56gxub7VKolLxg4izq4OgjA6xIkOcDlcQX/JbITy
69jIo2GkboqS0maBa6OlqVmH3KiQ6l4aCIeHLKxF4Jm4iJeRakCYqEtGZKLEVZlL
v3WAiG5ftPLvME1937+O8z1cbmZ9XKRcpe+laMRPvFgPu8E7HB1NP0gDQ0Z0k7fD
Q+tDh0epuYY1Gm/ARZDS4UX3Oqgx+Uj6fgogEFNpghlFO4UfgHpFhbwBV0w7bjd/
2KsItAHKZ2EDAm/EB/E4BNW9UZ2eloJsflrfT5MZKgrhbFtdzS7Y17uPFd3IDViz
bFqUJvgK9TLcurYoss8CaL5E/aoW3JcHf6V+Lh/BYBNWiFLUYDtgADh1CI8YkXC3
UiZBoirft6yN1fBDlYSFmStCFGk8oDQ2MwKnKD5yKXJNSCU5psr/Mc1K2gL+9m2J
33L77509araCkeso2TM02dweEiZ5BXdc3MSRoGG5gXP2CJHQrnaj2eE6RiPlafm/
kyUsMzue/hOHZYO043eyKqdZeAZeaovz1lyue67KQjqLIMs8RaDSHpa/g07Mgt0i
DqSOCwN59asMYPDomJMmd5OJfxJ95qiwBIWSzTm7wfzPRu92Y9QQjjhWATnWLxbN
W46QjOh9EBchTgvxCwY0pVC+iTlkp1eNWd5OASSRiG02d1vmE4SjU9lwSURUMEtP
BatwyUBV86hbru/XRrNSBc76f1uFdNo1vk36Tv4p2pYRWJgAABFAFdTD8YLQCA9i
nD/CCZJFHunBPQhZAwx6TdD4+A3WbJR80uz3H0TcIvoK5/kCxS+NkScKIWPqb0u6
LOalxSQtKLVBMrUXr93id0BoclsuXjVkxXn+sc71xEwdajbwJFLAdgNHtj2Iliwg
S/hP40O9UqHMcDpmjASQ5u7Rua+gRp04p02AUoHgYiB5soGwfFojQr0SyfMJUhOc
buXHbWJ1lreCL8tky941wRUrcV5g0ihg0/h+nxmgfpLpZYLqHXWc8FdCr1+uf6aL
4YNTzPs3fEm6+8cWmSUKiJPr3vDHk2vECdw8iTxZWsNCtsKU0gS2RUZOevl5etMH
9HnhBW2SaxYlrVwCySKS8iOY8xYdav1Y1gmNNQZjb93ptuyq+d6g6eEZGMVZuQcm
JmpqV84ab5B0X7iAAEfyIY1XanSx50nocxngyQo2jGjt72WiX/twbsHhMGnuoTBW
O/DqotUkacNX4q7lnQEneDv1rxgeSgV0pk9BV9te4G0CIkYSIRHwFN29Qk4ANBUF
Ph+Ma5qrYFSI96T9xW8sz2+lC0znZyzjsXtvvWyUwL92s0FExAZYsqVWgb7ew/Hg
WiwxAd9bp62i3NKAW8mA+CHUw8LthTn4zrTpwM4M8E4hdwC/68Eqrvk7fJb0BjZg
TBkcGgLYhXw1RdI+DBOWqX6+uMP21h1lRH8ke/epzVRJvU3m2DN3d6i8uqa58TzB
WPiCy15bGF/FiUsVkwIi8PMVOfBko/73bi+3/UXsDIhSvmEybjj3gOcy6cbhGHwR
ujg+WwgcOrl/hgpOhZcwTxKWpdEzq/rUBuhRzKn+QqzipKrVun9iEpcHhfvdRi69
Fl9BxMRT2hgtSuDcDZApbCwvewC36ClB7CQzQ3JUFM2rZlB4nTWPORSFpmu56G7i
hF0sScsp6owCp5QvGex8lEwb0PXWfbawZN3r4sULJRj7yjvMo7b7Giu1ospPVkvR
VRY/gVewa8n6NAMER5uX2Fa4zo4smuPSqbuozTRkFbYBK1NoJwHljbkW1kgRj/pm
edE21/KIusro6ETyk8RsLaNR8CJXdFJKAZ9Aez4CzkUcgFjPHLraBIE8pLiqU4po
TdFN2raJYKIVDgtADNmw24YKMIDQ34FBUCDlj4aQXeBBn5aacxoX+Z2u21BxmeAu
0JU4hscpk1x87T6I8gGQxial3Kl0tNZN5no6SZudLlKNAmt+cWGNNbFHmIbXvbKS
0vp7WMZYVdDU63ZQBxqEit6qTX7SLM5+ih7ER/xnUzb6A2qBN3NXdVQt6nQhuNnb
iSmOMsnW7iVRC/63VXYC0YBP9UAGp7VLH635InSmUl9EyNCl/9qQPv2jLVNSgDdT
56xUJsyghtlrl2CgrdhaDA5aJku0Z217SU+tv2sL4wQMM4ZHbg12Uyym0fjd9SJc
oeplU0anl7WNC3FJoardUfrGUZMt9ERbvYcm5Rp9geERmEa+dhinzzi+qOL9ZYcp
Z+AuyeehwKTl1NZkSs4Zj1zzMUYj3/wvzEC+EcaKwm1Z1VfB18lHtsIlM7Gn8+Kk
dHGNBoO0ZsGkwuaHGQwCqHPnoHi23uZLzX0m4T8FnrVwzqNLwdIAZ1oaBL9fhHHF
7HUi9K7Cz+y2YQIskMj74y6awWu4++C/ybCCyIWexYdqYcUD6NiSR8KHN0cB8vAl
r60eI1qgFgxjDHCRP5Of4kfKUEsf2yQs8DVFPcHukYyN2zjwY84plFlw4EbkR00v
NmVIRWF8HDbL3S92v8U9TcI/tT9vYlCl7Kh7gck7YfkZmGP8cZdaONnnX8xBHeZy
u0po3cMef3nLYoUP3rvgy+W0UamEMet7WCWPoA8EJnC3kBKLeRGw27UelvipCAy+
d0Jf1XKmdfUqyMH927Kq+4OcNofNNacAcSxE00rnxpDBLo2/1Nc9yBO8v+PIbqgv
Ko1EYGiRb7Or+RnKFKfEKFwHAjYvfFyVtCMY/CmR1bWa3M0f5vyr84kYN9zEAdNk
sRAP5tkBZfNr89EmLI8fLITklLiNO7Nly9mgiXrg6DhkOWBiqZkObu16R2FNfwrN
1AgqUw472KaSId3eQDoxw5X0wgzEdqmOcV5RgRm099kwHUPUJzwJ29idgr4K5XgF
ukoEfhenR1zhdjNDTmup5R+V5H+1ZKzyBxUjqR6sk8g1DBmhm1uo+kctDerTsIcn
TbgKa2/E4/6EloxNyNVKKE116H6tdoc5VTU00ZdR9P62x5XKXPAmR091KW4Io7hI
ibHm0KR/008D/rsnKpVRJ+vvCKUdE3ADSYwomeLPvWguTNkOXov26NVq/HrN1JDU
wF4ZwHXsg/gmuIbRE3zsbmsA5vJHemBnm0rXpcr9jLzPsVYJx4CsawHuBBN4manz
e7huurCekRqPNqoMumKY9/SMHGthOGz0m6Dr7I4wpBJ1PJTnLFZsROiPcQx8yXTB
neMRJxSf79ZKCrq2ko0oczq3oPL8kSZQYW+RThRKi9jM1kwrj3rUj1WR5RQXPui7
ppY4TLfBaaARb+HLNgoHrfRJKmYXGM8y3Q8ykfW1tmOpB8rG/8oK5npHhnDOkaMH
jWsc1mlMpGvLOTlN/9sgPXt3BWeC/sIoGk2YTyzJM2A=
`protect END_PROTECTED
