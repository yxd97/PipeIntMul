`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4J04x8FVllCll/4dEBYgw7O+MGNyJ/Lt1wbG6jotOsmzbJTwWZyY2tqvWvFQ4+H
B7+LCpXMcuZ554gZsgG7jMYfmTE7oqGEUGUPv4r+VgHg53Aj3zphMr+ACTuxUAHf
ZV82T4J1GleZIjpA3Z9WoJaJwAWYdRBER0IDX/v2hGzTkmFLe+vjCd/y1Du+dtNy
8LI6H3yihq3Qb6JyWxIueGHEGQru4LOa8nihVZRaIcUf/4E7xTa1ub42d2NdumPT
escDC0I4d8vCAgopXQx6EFNLEPIKjKQF6DRGCyaDmiqccW5CXxqxDSduRgF20glH
XZ7cWghG3IeFL4s11v7dnIyUBApW+lEFQWo1YZX7GCNA0xJ3GEYItHKgNVO700U3
Mp3X48ODL4P9EZ5oEfsjOJno1V97TK8Cbn1/KGaqqR8BM0qHJIv9J7ZVIn0/OKZe
VSZUNI62Xcso5m44x9lTcQjGwF2rp+2GdS/HBoRRJQ3+ubxPrlsDNIHkzi3nG78G
7HKq8L7PwqcEjJT+TSCJnGTaGu06GoySEY0SFgHGPK5XpAL/MwACcDQ/z5t4je27
dLLqw0JHKBp5V6UCuJN+3puGRB2b8rj0ajdpIsv72rZEXbuSrxp/Tb0CfnTb8awW
Sw7x2AoeIIzu65CibOBsKR5xUJTUQdrpbVj3aBYybjsfM02UZWmbAukKnpsf2aHa
weub8vDcJewfNQFgh9sKHW6xzjz4AbWWFOqNNQ2ssdfxOtf8h4sYNGWPh4Kv+JJe
Z24Ee09aJj/IJxxz/b9bvW2w3c45KE/VYiCUahIWAME5GTznM89WYnms2nKuCi58
pkK23C1F0a23iPoWFRdhmgti9WmArYHvClVLUAEgjpn4O2+VFv0EGCsNiSUGw+0Y
6MYfXEBA3oVEh9kmAdeYQsY34X99zYQz3SebbygXilY48kmpQovtXdhgPCSVyEyT
c8SeLGcOGjfpkBcG6O3Z2W6xQp34dNL6LEYbIx/SyyApUs+aX+PqtNCIlIvEc5QE
aInekEh59lBJFeuv4xA06jwSItLOjoBZ5juPpsvuDX+zQNWoK+AQhRapeyXL4+3Y
pgijlhkw9QTcagPdyP+RdZjHT/+7tABcV00OOrkfDRnml+NQriLk0UdHtiiryNuC
RKmyR/dsEG1FqR5tKT9ucuNdlxEjQpO9F7Lxz+PbDtcXHK3E/5EIFw8txUZ3FcKc
l3YOHnCaQ8ybqWVb6fIItlwyTf5pMHNN2mXIEjgUwphj4PwgudKlCO6RUw5BbJQt
R7jldkjSke8IuYz+gu82EMa4fS5PpfJmFJj/qgru0SSEm3sDP9md8AGZQKZlXTZ1
pfyn6SsCO9DmHQSqAEgmXALfTJtEpudf+RvQj1k0BBfm+8uURSAcN2a3ePUQxdLb
D3FShMfd49lzYlUBUitfzHyLNjeZ8rpJal4tl29oTRces7YuwAfN7mkj2ADVj+kK
WAGbooxuIcrmPfz8Syjbd1nCMru5y1pM1EWW7S2bScNlP2xDeKl5MyG2yTPyhe46
yavftLjXNf+JEm/BQyqQbDOlhN2a85KoLcb16TZU3IgQZqYJpT3gzL2BPILBefTi
m/Uhw7uGGldofTq32kSiDt8QyTRKc7lGuh58wbMrpcUsJkX9YYWBXK8/WUmlLLpz
sr5/cQExVdFQVNqWJmroJvd+MxV9Ib4IzmYRREtAcugGWVQ2Usz6po54e0fj6K2V
359IxXhyUA+uC6fqlLCjdU/+jsCFe5a/7o6ZB5K5olgpxM2Ecm7HNR6aEJ8mR4nT
gyxTGuvB4Midzozi88IDvS/1L5jl1RU4TuH57G/UEnIW2WTzKxZlUiq5D3vIb9VS
/bQ+o0W2S8VVO2WUWspsxg49zZqth6o+bP3elUs6JEQAhEWlydNHjfErRUZzNh41
yU1UEswFP3Q6KNm42liAe9oV1Uij/bAOp3oSNYg128jWYoE3Y5OlG3hK6D6NJx+1
JKVvJ4iQAPAoa9IOLp0WzmD12zEoRGI+TqsdhUMBWA7R1AkFFXdxSNXOZj+Cz/am
WsZ+TKCTCsQ1p4GAnlIgVig5mUpLuNLfjPDymSEcdauuLK02VZq7EfK4prnxdqw0
XxvVio+Gl5+/mpPCUq2AhNxiz/S7N1+MDJ8gz4Cnlt8=
`protect END_PROTECTED
