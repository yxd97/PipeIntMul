`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RfAJfs9C+Cg3F/0LLPvLmmhms/auf13ivEkfkm7Cr1YGeHBCzrF8RnfEen/Qg1wU
bhd7CarN7I02QLwO8O3rrHhYzQXuaVlPs2WG3UoArI3wQzvSvEDEboGDIcgpPPAC
9w96nwydVJqCrpQfJYO5XZ2JSJeqANhopSSGBhm82DZqy30e0JSua0veBtlo6FSL
seIfyM90EKt6EASFcYNDlMj0ln7AWMtMbiGzTbdDXJmvBsr1hIPRKwQa+q4Rtpwj
P+RV56IhEZ50DaTsIHjRMg==
`protect END_PROTECTED
