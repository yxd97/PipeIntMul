`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
autgTMmTg68aj7d3/x48LqQvzDI35Y/2/n5ZWR721OcSHFdAmDwNqCFzsJKGzfRr
ncT40G2/8gBLxRFgvGkfWk0QG+GkiMNfw+gus8xhzNbScW5NnNFee9tKAhhKiWsH
9DRBAeXtMppLXYRd63/e4uTkrDSkIeN+XreT7NV0rP4kKcxhHnsa9OAe766bF8iF
5FBtOWqIjE+jQOTSR3iVk9oopb6Tgz6Rvmame7w+aRLEir5ctzZGIeWe7iAV8AfF
hpTeEdXxxDkb2GAa4dZxERSv89eNpmmgWKxipggBqOt/skclwTnIpztkQ1QkfOXH
7rLiRDPbBfTrmulQLkDZ/hurUH+vqC/mAOe3ZtvgVOXe0vtO3VRLkeshbANGmHUC
Y6lu0Oa/YxmL2Du+PZKI6vZhEhyV08gSnQnfcR38zQrRQOWmSA6NZeJm4rHJbkq9
ZPP5cu2A4WanZiXIjjmazShrpYuuoMaou+s0jMzveY8z0mubiageS1bZYDyd3VlM
G/t/Qoojhdm8ecjnhojiSY3nAjXmyqkVAFpCDlmwkH/f5KGKws97Zh9mCH+66kF3
zNTWfEkGBUSWHyLc3PU2HJD5nBj9Ijtm+eWBqHOm/1QW2ywmB9CfKtMS9kWZnyHX
aJ4kpgVuf+aP0qAVLTZwoDgsqlxWolkLECGKKxt3ulB1A4FWXXwtmrYWXAtFXwtn
KiDtV2BW9h2D//C2kDjA9YS4RC+UoucC4v1RmHTbg4D76Nz+r+YGA3CVJqg28909
sbY54T2iTBOmxvOOu8NBeemsHy4g4PMo9Qbq/AB3sGBOrBbQ3IRjJLasSbYaG7sq
y89IzOUcxe6pHK2HnnhmcujA9eyUhg/pPqJxK9bqmrU1BrTllnLIiQ7cR5pPkneC
2jJSJAn2EKptX+hev1y61B1wD4NjwXxLRr1rM39hD+3rfAbiYbiCRNCj+LfmLdDY
LGHGoBhnu5O9ccdTxrqW3nduVBQaPh0WjPeAs4U1JuI6pUrvstbmE+fiKAC+9WI8
KqcIxNCTrq50sHoguvPW2LDypKbk78gWikf1wUAkcEWhEpUannD/uE37Uqju/v/G
SYlPbXMdZV4aouyzbXDWkm3ny+b4BQ+pezPo7IP1LMTxDSFcg+43k+c5m+mYAcN0
jxLHDjqIUwR2swgJAM+dWT8QQ3wCX6EO/LvkZ2Y/wJ0F2u1efIxOxz/aFRHuuGJn
jHNoxXIIhehSsGyj+Aj0x3EUn/kMS7JeQgmqv99i9D6X4dRksj0dhzFpCQcGbpx0
GPecufQfMTZOEykJJzgX6mRLC2txroa+nRjt9mwWN0VLhx1EPZacoSXWrwqxvyrH
8fjWHRcKkVqe93UD+P7eiRFuxZ0aUGqcK1DerNjvKqYTwch4NdTPJdKWA0vLo79z
xKDFQ2JraG3kJkkYGEPZ0jB/OJggYID7iV5rdsuw0Pet0waKwu+pXDq+sUpivcZl
AKs7BwDWKfdoQaopmzIegw==
`protect END_PROTECTED
