`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YMt1Ns/Bnq38Yr0asogjroNBp0EfYCcMBDya8U564c8E66KiAtUMsyrxeWQir8UN
h4ZlfrdNLzAygCh4g/ojQGGGb40do+yG2RU1I9x862WQBimsVXaLbC6n+/Cras/e
tvQqF4XPXztcULgwK/9vpSBxZUxRMb4yTOInbblb+7Y6UK6lKrcUQp16hRDZdfrk
hL7s4Q5+DjzB3fMMdzOp7gK2rTjzLLBWKzj63xj5jl8bYpbIF1tKSCtcy+PcHoDv
M+qD3TZYtkZEbATKksLnsA==
`protect END_PROTECTED
