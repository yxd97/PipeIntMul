`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JILbuqRjdM3gVj4Fus/lqRCosWCG8zTPhDy89kCnz3nLoaJ35AFuj40AiVJw0rtA
O0s/PPh/nNblXB4BxnzRWAkKH76GrRRirswsqhRHcJng/yJV0j+poEbsYb6ggedY
z5pGAH5ZRyvfmctVuXyhKPK3JSCdc/etnHKK/9yc3k31APmuTqgA8z6oABZe/LJB
2/Lv5dshKt4OboAhPEK9ei8znIuSjz1PWTK5NkHR5aTdF0/A711Dq+9jehqwpmvw
Qw6BOAb2xjZ4kzXQueLRw81HODKK1GSdNEdMmyPuQ/pONTkH+jxrHdstksze/Abl
rQg1h1xFBAFvNUXBLIyOwi6gcrS4AZvqblMW/bP8f3LX5HkUJU9lf7dZTcO5YHeh
UR/cWjR9L/Ubhikm2oCdvXbEE3GvF8MJ4Ot6qBXLVKhBQx9R3bljXdbPSQwK+1aO
jC/ZaIFv3izZKdsLgpYRneoAVaXTo4ur2o7Sgjub1MOf6Pu4jAl+1SH25ZOe+DBK
1XMVFpJ+pVaGTFeIxgmQZPk5iVCqAJ/Uwi+fVBHIGDfTO/upXtOdTHg4Tm48Ex6d
/dYCed91IK71pACcyPcym4rMBNDM7GmNStwcZN5WSS+govBVGxdt24+PWPweHJf9
I3PE3Z8R93qQFn4wxzn6OdFsKV6Qx8sVtdeTutkVW14XlyDsVZjGFsfy2dkZXWI7
7944WdJXtv+a5b0SvzxXq+ESfqt/Zf+sipA9QxLJt0hbIEu9yhKtwpOZMdKdqny2
UlesjglaMwpSJFPWIKPwqUGG3UwTeHVjBnqxt+ysPJNtO2mSb0LZomPFKb26rJWa
VD9GzB26SN6NJ3gBJ1d8FLSTw3I6BbIHEY1clAIG4Yh9y8hMqgjJWo+yzs981X15
3owm9qXF4ZyRTn+NpFi1YaxmJjO/1loZRioTSdwZshE=
`protect END_PROTECTED
