`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Viz3v3kpVMiO8QkV64IHscjUX7tSp0rxmQM9pOlFnXQs+pDbUmwoxYJlnuGtgVYf
N8+xxjbbGri9K4voujxUfV2HEGLUmeOYs9fiN6sLpW5KpG5WNpuDYALtstsTAYrV
1BAUG7lxJmaNUVeJtZur4MC9YZyYqDYc6dJoQFwVQF3u8E8toyKhM0Q52+2nJmVp
C4+OilCOHeaYvQulV7bSO1ywiuC2SMYn1iaoWjKgdV/Unr+KHerBV5YmxM5LYSg6
yzlyFXwUb5DUMQk5q0qf55I0Ywx525lEaJ7VO4FReizdDiS9LHhJTfA9FAU4SHHn
LHiLpR4d00494YcgifQovxsZba+k+psCEkLojhPk8J+gg1a0+pqC0U/uMY254wlS
hljehgDBVA1Gv7zNOrgW8wnoc/dXV2/TVXHPJQAMGB+1xR/isldEN947o0iEk3Rf
eebYro2q6wmsF/3a9Q707xV4SH+3cZKgcaW5fE06kjEerSDPMfX8973Sr79kb2qg
RByilMkprwYea+pDU01YYXTIQZoPI5uzV4GxpOB+tlAi5HZiq1+GxBRC6zm+zxRV
ibxkBLD2uD9a7ZUQ9RwevERpt1DazfgHDIU+YeNsEPhXOcyhAt+5b7hqK+BNIAMv
IDVC/Xy6CrUR27imUznAO/z/dro8ZnC0efO0saJF4vND6VlvlIv20+tqnh6tCqw1
eG3Bk1w71+phHc0PRc2qwbdRcJ2+lOTG1kdaL7XV/CEd1ydBDO0W1D4CfAUIM7xB
rQGa1/Dl9ivpSTKEdGCFHjJluwRD/GZdu/FqisMo0DshufQhl9gNT/9YJq43dqL8
QTLpBNkpZMjmAkBLB/JkgnkckUh+ZZfJ5HsQzdoXRRPYOhAh/CdB+LlZbRBCVfE7
TEPGIrQdQLtou9x2+znQZQ==
`protect END_PROTECTED
