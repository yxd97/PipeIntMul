`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X9fB5X2UUxzlren8/AxdUVbIT8tiPuY4He7XhWCgwTkHZsCHCRHoL3cYa6Qj6D+m
mzUTjxDJXnzwMLlkzW/Ohc8RonGPECYuMZUtpjnRzV1jlvkpShqUPW2mZrUZiEfR
leJStfN195T+MJyBDYepQLL1U1RyiPfP/AjM2jLlMD72C3V1iZuGtV7XgK2K+r0w
qctwwRXyQBlWm9g7CvBBzA9/4L5jNG6IEWqnnMksTsb7WSc33LJG3PsdnxCOgqeX
1jOIDPWn73alvaDRA0N8uWd7zGXAPy4nGsBwVh49f4zsSNoKD7tEU01MQ72GtMod
Irun0MJnY5nP1+PzlWN5u2O9s5cqwTdt7EYkZry5BxRQDUk01hr7EiqyWEGCTeEu
vMZlvXNcejxaWLTScgT6JXl48z7K5Gpj37FjYLRwDWC7mtBAviVHac3+iPF/5jPm
gDDYCnRWTktTAKmn85U4NOlpF/wK/22DUsPHFMWu9ClRPBh63ds4wpHvNRv3RhYA
MkoVOyos30UerA09jia55xL0otqy79skkFIil9YKChv1+/SsNBjV8LgN7/ee8hIR
+lomXIOQGzbsVGsE2eF4nsobkY3M15sKmWovHSfVxThPSJJAmu5+prIwqBKX6VYF
Kyh26zxBHsEtAFAveGTkcJLzGfyp7exddXEO+Z0Q5Jv0EW1ryoBQaoSAXZa2eW8t
3dOHr6zoH3asKxefzqv24yv73x0ThMmF9wUu1BvjVneYmRHAvqu5uCMVlU8RZWht
GNAapPWYXiBcun7Ok4OJSmumKl7hBZkll4j6vJlwT3I7wnNzrYouITCCoYM9ZFlN
RQzl9TPHYFRJN7JpnZmxucHrR/BGlkq8jYl3m7/eiNowznHyOlBQ+KDWnW6IKZx0
h5XzY8SNzzZ8CC/5WbaS2D6sLJPEc5GK9+GTqqh+Wng8f/j1UpGa7sV2bV7RSpvg
FI9RMTmgVFYUV4i/+p0Ipuc18Q+Iap/Nhiub1n5DOQExjXcHIsOjORIRD+hDVADn
YXitGIpxV2KpNuaeMqKLdFkIo0rDpuCh89m+et5mmMsnjrYZWk+p5gg/IoKRn9P1
eGiQyEmNIXotdSS3gL9ZfjKd+8VP5xhpyZQLFec1XeiA0KJESjuYUNIOgaZldL2X
Km9NjC3IpdTYiQfTtEXGCw==
`protect END_PROTECTED
