`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dS1yDaixPrPzJ+/8LKyVLfl9gFOuq59pvNyfoBgYRNxEdZ8Wwo+nkbcBjQuoxqhb
CGhXQTbJRzFRzHIDzmRpOoSo+pYxgLd5XNEt0qta+Scd96f+mZVgxKoFUq4u5D27
Kz7/mtU8F3ZaqlC+IjDJTbUSNuMAOi5Pz2fCt1QEjfKE9yGdvuLHM3OtSVLUjSN6
PxOxqnFBzEZSG6nASEKLUR7STlK4Nw+5Zbiiqh2KAAE046jyQ4srTjzLd4j9ZPZf
zX9dPJLwsMIwVe3es0kxtUpErHsINCr1LvJAA6p4JhFjt8x/0gfpLHkIi7Y6ByBS
9iIgdtKenkiI1KkAotc00L9tY22yXSlX1RdMGLLqR06FUDKv3my3DiwqqOaTLc1m
nFJmxobMukTaMemusTwRSWBojEbwDZO7z7GBYommbsr8DPemHGdNxeS5dspCDRpk
jsQ+XBSiig4v7ygji0xoWklH06v7UdOl/KC1rOrPVXP+di9hKW/J38Fcvll6vG7q
TrVcB3QP0Jfog9jJiixRet80s/FX+muXjji/9+YVwjv5ch3Ia60IfpiHnDAzOIUo
g5R6wLZC0TkNC12WlJsSc6Q7VgT90/l2RcwmFQgdBRy5Cn40DJnrDowVd+w66eAC
+fzd8p3gJtDQT6k1BYn+hRhO2qQnHZ+MAKcMQdFD8hzaHbLwpsgoIZ0dcUjm5wbG
myz4qsdM0LjtHBwquY11ViCeEq0/QfkiZcEeWXPmhU01jS948L/X38scGv55EQBa
Nz+Xi0esWHVgDQxJJvCQB5gFbUg68Nixo4jTtRS5jL5CFR6vRzrB4XB8zKOwjr9u
byl/ufi2P4SPJ5UOkHW6Wp5UWgL1LU55n3g+2+hbsT4=
`protect END_PROTECTED
