`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pfbfNhxAWd9WciZUaA/ratUMiTsU0k4AnmpS10FLTX7/Q6N+V+OvCytLuOAgn/sx
PzU+YIjZJr9hYCNvCJrpvAxWuArU1paWyeTq3sPGCa0IZlSY44rwbNfZgq28D6vZ
itGiL5EESlius/esM/Mi+wnFnXOYOOH5xQBDBBRlM35f3SXIXS6+wignvmWfnYLt
5CVEAZzIaUdyKavQvXLIiOgQhKeZRrjYCNxaE0UUpRBZBfw9QPgFaWtbMJ8q5M2i
8rtLhFCOWY1xc81QUa3JsBN503Wn1ylO24OLpcMWrTIvOkUIPZIX92OIpE9v42lx
JGg63yLwd0/1xun9gx3ww9t4S0bGEFZz1xytpqNokx3A9gy5ZI5UvTtMmr8ANXDx
/4tv4kQrWZ3FfW9QblhIEy2uGThRqfFJwSn2+llDo78JHv4OEVdGYo7Hmj1JR+jQ
tjATY0Lz94fTkdDyKK0F3d9dbrgrVrtMrCHJABVLE5U=
`protect END_PROTECTED
