`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dnIE7NS9acseOHMJgQZ8IF0J9q3tb+TRH9h1VcfEi2CRNCwI1Tr1D8yQG4XFls3C
ZPx/Pw/dl7yjFBM3H/qrRobOjs6JUD75KA5MymJD7/rCPaSLLVaqIFPjeJBF3oi6
1aFZfoWET05FUq56nEIjDV151kKVXravU5qcTurKLKOvfPUxStROzQea4+peGSaA
epAup5f9SD2oSfRQcUdAeSoAzKGDMFm9mRxHHzjZNm5vszLL4HwjJXC0VMcq5r2C
YKRHSGfN9zsCF/K4g3vfdiEgN3DY+Zu5iwU72QeXg9e4ZRjgRc1XqhKMTJzVCqlF
Yn2Pp/gWuwvA16mtzAXk6MOJ8pXkWDu5Ap5NzbLsRaj99OkAQIw+RAZzCqNZtN+0
7zYArx44WGvAPMHQaBuCBs0naOw2fvoT+OaE1FXGBd8fOa4BGl8ccHZY5MTqs8fX
56bwzkmJlwRe/aNOxdNem42LFF9MttwXxRT7fqg5Vh2cU4OL3kkXUgChFjc3lWN8
`protect END_PROTECTED
