`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ERsfsxgMx0EptQF04nci1vzvObWH4RUS3C1nyCTOCiR39y24eIxxASR5+m1M0NQ
uBQmQxO91FFR1R1u/IYhzHnsJMToNcOaOKzXekbsUKDr9fBW7+M7R0DvoQ2iAV6X
QfAl466gidnfRthXZCD4hNbRHmmwhQLl2aaih3vrAGo1Wvf9Y8FAT7Fs8mWIZ+tk
ihtYM+EP7ZzWigfOSWw7ZoO4LVP2CACDEE7l3hcdty9frM49WfFSi61GaSj1FFOH
lKeLQvrEpL8aihG1Gs/WMsXe7evWdGtHyvTASR29U4aVyBUgbyBeGCiwp0qxUVxl
SvMam0VRX8Xv8z0oaMyPqHqFAizcR3IBMiRRVzuAenP6EyWBXpndA4EiuRIw9sHp
pFVt+c11AXxA+P82rw/1z9QelFsIKseIy45oy754jRlcuBaZtVyqXlexNuTMgZUX
h8sc0eKpJ/lRjwITdc8XWOhd8f2bcA1NpQVCurlInHeepyC98O2UhFDRJy3OXcFS
DSPWAjcORoCowbS7i++rJVPybMeck2ACLTHXtwNdJmHqWZ9NNDe8bSoWPUh30n6j
FcJJ5X/XnmtlqIjF49MKwwfpXTulQuTbe2ZJL6VGL4iIJZVpjrqx7Q/hjQOX2Lbx
xYcPI5xet20d5lZ5vO9NksTqaZNegurGyOF6u3Rnvj+aBVPtXjuFwBLFJAgTYyFz
Iks6TcHJHKHNduQSE2OwPw==
`protect END_PROTECTED
