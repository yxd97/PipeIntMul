`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OH32iahIyxyNwaZs7KCk8Ywj0xjTswoSgcYMB8RWyfDNPXe4euFmGuwM/Th7cC5f
aXrf/4PFj2NZQmnrLa/xUnxY3i5nPymFDiqS/HNcpJvTq3tsjowvgZDiTM8V1ZWE
8mWVVYvChZGWCb16TxuPYuRh46vQixupYwK6sUzD3T3Bb6OKI+dOEdZ6iUUBd0wy
sg5t7iNkL2PA4nHvLC//VTtRJx3Q5T4K7n612xFvMxJ3EaH6KGEvniXDqgXw56xl
Cc83GAMRepqvxRQKVPz2xM6JFPbWJBdN2+/OMlM3k2ATChprpVaGsRosjBgrJgPM
gp9Y0QxLs2R/Dljqj0RmlUZm7dCEJXsN9fb+jMOoxnQg/fEccddt7RekC4Z4KPZq
9sx+2zqBF9w0m+x6HHT3Dn7b8DCAipyddFi4jjuRaiDfJjMOjpoPzdZplSHuWBmQ
SdFYcxldysvs/zSoNWDTqm666UWd5h8K2mrQxtvZ20JzwpqJYuqIAiLgHc6NEw3X
xbTtm1ERF/jN5dNtACwrS3zC96bJDEXWGUkyIQQIYcjRczE5AMi8rWqZZwDQ4QTG
gRJ9Ph+nZ+uKUk6fjeTZ6xYDqAOsXtFt8M8JbiSiFqGCo+lNyG8BqJF9U28Ss/SY
j5+Lu7W0+YkYY7bqDap70HH7nY3P/+kXUH+PnXlChnD5EAB7Gj/heYLdbcC0fso/
DeCd3RKApQBkaT4BcOw8ZZ8OKj+cKHR6vCvbLxZ9y8DgG9Ygh1yrkFX7EPFpw6YC
tv4iZG4ArX+uBqNHAv49vXR6+SYOI0zirsc3jZsj04Jix0ifXI907xzaDwbwdxqy
aIt0ax7NyMzRbWgaDiEC8Gk42qPJ/cCQ3clfctYZQwAITqkAp2zDznnVPxppBArJ
khdh8bafgxihp2XopNZ3S2Grj9/p8WjAwBQe500uxB5YgPrQwehcqJ1xemeN81bf
elbBspfd+0TXy96aBWrOJw==
`protect END_PROTECTED
