`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EASIyDXOk11saoiaYa0ZGQU+x37bR3SKofTC2z7VvNrYPdXz1aOJYZ+pjIPNJYcv
gbYzqYW5Ol7IOGOU+TMYSIiUYpPiAyWuNd2hHuGCrB24S8W8Nd6QO8ZajwbeiUjA
aPKzoRZMsDb6ucY26LpH5LybQYtYWf7paTrfbeIFHVSlrOBfqnGSzHivfQzfEp4Q
8FlaYDhZynJZ9iLJ5Kseqedg6OSFyBr0w4zo31AxukQ7AXFXCHcn1gkemLmIzdVD
jtg6OJYzFWE+0lVToBIweDNOcgBkpNdR29f5L6l4THEwwTc3tE6zHHkrgsPp/lV7
2NtbLaDnA5gACsX2WURMpgkYXlSjZb5yFmD9GBLK5ZU60onwo7woapvJRwzeN3D7
xRSrDhwGVnKWsvXxVV4lTaa+C6BfKb8k7MRkcVOp19pLtKynjlz5tzQxdm1mYCe5
8a3oia3FFuHOT6zJ3DPzT/G/w/Px+IiX0mqtgt4Uhyi0c3DGFqCBnF8iEBYExID/
f+Y4oP2WZ9j9DUoGwp+Da+dMt6bf9UJRyt9/hl39xIplQvYUgmOgFRazYs5bYQI1
JAD8BLMncnHpWTNH6MOJB2EAEZ6aQgkKDZjT081Faa6mGmJpplx7yP6I0o2rzbLD
dpOkzoTTq70b4SDGI7hFbVMDl4ynmsOr1vV3LBU2qbk5CZT3RHivgkrKUX8lnNQ9
y68cInM4b8W1hQ5cBhTQ2mcEnAbpAv2BpXHYZnTZC2NtnNW4nCfOUP95ESUTI+5a
Mc1992n3S1nGK5RRNaKYgxHiyw6IPWa8eo0FDKzkzKSwTcJxfgCUr1RgHKy3bVJX
Ei/v5njvPCso8ERMMcJJd6EjkDLW11oT6swUgezJKQvc2/PIAGV4XARJiM8ajSVh
c97a+ImQFzhl0otb+DB1d9WD/45YT1lpVkyNGlED6Gq5P10K1GJXh5le8AS+NHAX
YLIa77DntQ4AyqTOSV2II7q72rALv8Q2iCreQmmq63KEHjnbTIlQ1lE+GeIcjNvu
nmGFPXagku3OgLPql1YlFmGJ1Ws9DcsUHNbTODAW/kqE3tiGyhBPO2exS0KjHUSR
CxfJaqn98V8gRYXL3HgRPRXA7dofYQicp3v9zDWWdwjMTt811UtVkXfJCo9IV9QI
/7FO0JL99thQXbQRpXUALXqR1+n5Sq0dx3AN5bD6X5j1LPnfGq8DuyFiN692yHKr
i6Q3efdJAgvem36ix7twIxrnL4nWktSpRKjzVe+nkckqqgKJpSgk/RLVchl97n9a
Bu/mD/ssvtc4gYO3OvAskpwT41e84qX+/vBwGkdIFDwX/+AV4JmU33Cv9pbbhKiv
coDO+pfIs9Xkp+h16tLiHauQlx5TzmTZhxMOjYmZf4/7jzYaVIDSo7y/q6fjSeTJ
3t/DHlAXCvbn/JYl+ztCreiZa8uxy7UeIyHfp4mBnsVR7/ZzzImHFbCpu3sBixM1
7tm0yFOSogH1SVKvnKtsyC8SiTzxqIYonienX7bwawK/sVQ2VeKEErsz9kLYG2iC
Ujh3YefbHcYJmA8Q0wzvBW3Bc5GunE87FbUgDZN/R3O4YuH5k0EsG+3egufLy/M+
UG6kg25GiUnVVSaVuCC8H2WB3ibE6xVklNv0i54iejNzwPhc9m0lP3EaQSKZEU9c
reNFNhxtrSsoshiDABcUjY2AollEv5rEnSoIKgIeNma1l9WBvR4dXkBHSAg4z+Eu
62ZgxigVmRn+GjRSbytWruvTfhWCRfzVEG0UGp1KRLqRLZS+2W6th3xni0GWYMSh
J6MQcZMNZtNwf8klj7si4tJR5dbFjY2t25DZiOFrTt3Q6WooS2qub9189SjQvieg
GazUtW0tJmCcvfARnVGVzEffT7bca3OhguLmLh2qBwcRxYoKI05bpbAgumEqnhZ9
1uNXeXJpnemvtTE7MLvYOEl+hl10NAk99z7bViI2coQrttgr5JbmaJyJNM8TTPes
h6XhoHtr5rH3DdaAKoK6Htpi1meI9n1y0z0N+mkY9JTo08tSJ62H3GVN5iLukKZd
0tL1ABhpFCLeDYiNznoxvCAUASP3DKFvGCQiB8rCuxeoJLcZh94LVx+blsUDo3By
Sh8XQiOFPDRMA2YXbeOrCtBAtOqzT5zwW/wADj5dxg7iUdgkxc6yBZluU3sOW1Yc
29SNOeALEVkYtN8vtYezcm58p0rrgZYFtzwsnx6aOH6XN0QkB3b4MmHtqtUsr82k
Mz3ut0g03odMSCU9bckqC/WhskqyWzfc51ZTC8RNWVlVKjnpnqwsI94TkLYa0i1X
WmSTcmXoU8vvwjMjXhxogoXYo51MflgMuUrsb9IGSFPvTqsUrDEOSQKa7HLeQGz2
OW2uVxOaVGTthZTL/hPhfbdkv8WDcGGMHpBiU93TAGPehhkAV+NtJT7c99N7zN41
SIj0RrC1FQGB7of+uWB81laBEOezpCDowLanG4lTJxCBUMv03+RpI51oXmpa99G5
MwCSH1Z2C5iRWumtvT4g5c590tst8ZXAotzv4tRAH8mTdYF5xlLb1avbVXVBgwsB
N5/Lsw1WCOAVAks7V329I/NlM9lqFX7ih7tGCTl8oqUMCjSSNKY0AxNlg4qkAxOB
J1hT8N4VtrkHJAX8W1dvs1PTLy8sRpogp/byVMPWnyuesBVpctZa8TM9E/Esz+XH
70+nve45sI6JfPzFGGZfkwViorhyELMohorKVAfLATXMYynpMA6P8tL/S3Khj8Gp
ND2xs4pQP3Fsa/7iZLB8fnqSilMRPcOVG4CUGr/EnIhSz9oRaIbL9h4EQEQrQJyY
axKOqFONtfq1mOr+ElckbbQwvPhRvgiz3QwRwprrMoV7UTYdK1X4juXjMNe/FzRZ
h8ivqyHG+T/F3n0e3H05fmwDXQuP3/I5yUAAR2FBKGCkJbpY1vSJTkPvbLprFwjv
4Hbxpd42wjhTFJtY2zbDK0nJEAvUfci7sFBce89AFE4Dtq31ky0ga33LJ+drChcM
0Q22uOA3zopDHo6C/Kdkrt1kN3ZdZayZUiMgvN10OPg41qVvdGtQCa7jbZL2hvtc
l3rjFfaqN2BNVnhiJ7Ch4O0NceEGnM7zUXIPsjpxKk5CmLCJOVNlqteLsw9ze/fg
fyQvbhQd9k2XxL6UiLY+9T+sNhCfoovQvhcz8G7ws5I20Dh8xMQspJvdJdJaidcg
IuCaYJxVQUocPCQPffptBdF1lVqwFUjZ5z3Yd04S+Oia6SThKpuDLF1hq1G5IWAD
9xKsuqHLTVmBZnkVJU6Jk/5ssM+bQNdqNFJSh5o90xuuSpfTagqQW2kS6Mif+0E1
Y0lxWr5i/a0KLmSfNsgFx4WKAJbgMi+Qh1SnDzfMPq/meAPSuHuLY96t3MyCa7uS
xAruBgEsMjDjzrjWVFtwcEf7QmrcnsTSuv/lVdaoGqZPUJVvSx4J6nG5tCBJ3Tn7
SvJyC7mJ3Mg0GguUWf3XQRqoJ+E64msIYOz4de1SwruAkduO/kqJuYz4JjjvObWY
/wMNGGmkwhuctpleI5vcvR0xHI4rMzGt94dikZnUJ9eQr8YSl14+OyYYBJ03w6fZ
rN1QLrur7MowWx/LqNZa5bZbRfxCCYdmUKmIpYefNx2Fk+/bwBkcIxRXxQG5SY9e
POxEh8RmaEinlV/ctoj7FsZpqpSmjiBfJBKccDaTllQIpgrs7qGsFPZOvG4sbG42
cEOYnMYqDrS5zxtCahXuZWfRWvCgT2KlUd+NUw2cY+NOvX6W3w9QEENvjWw8ABbM
loWO9H/lHNMUgyuH04xw56kd0cpF6MR4SxKtAHgdJ6E73v3d4iHn/AJ+ILv4MZ9b
e5/F3rRY7RMRwB+hlgnb+M8djMrYmJjhXq5KNt+2p+hc9K2PqcFHSlDv+up5/tFf
uyju6EiM+4XNpG/MIzNTew==
`protect END_PROTECTED
