`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/c6ySDyiq48ENqz48/RwcjeatkSodBt1KRZUOFqPnEyGe8XWrFsukMmVz3zgic7O
t2mLUs+UO64ysqmr2z9fgGtXsfbCmELrn9H/b7ZFmyQDB8JtANhviWXAXd/QEdHy
pX6DxT892ySgsD4P6KnXXDIIsRejLGJZ6fHZvv0ReiebT1h3Yk3Y0CgbwlsMJQtn
kiuj3rRVsxhw/Ww/2kEDGU1Fq7p05Q+5e/+XXtgWeSuzwKBeqsT8w44e8P1wvUuB
b1AKr6sKJEnxNj8syXwkbOGzGfDg4Fi07TAzqVMQIcUJEgKN5y1QWWjZ9/pCbwbV
O7PFwlfV6wl1fFybbS4K/0e//PVK+j9G5ZtyZ4Retli0lwh3Rg6nREZkz3RqT13c
H9+w3LuH02vmquphjwhbRI2q9Qml7TWbeGSWmO05hcKyKZjs2UBOUS/8EnlYmvlV
Lhh2Qlg7VRYEORmaUqbylGDIf7B1WB3qK45muKx9tBnDKlWVmtbO8Lv2OgHrJgFm
HNdy5dvjkF2H47drAoHQP1WLNmbIxdfbk//yK+0fkEVgvORIQjjikhk9y2vS8qus
iEAULNsCRceWB6qyZzhglQ==
`protect END_PROTECTED
