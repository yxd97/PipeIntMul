`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJvK8+hv4qmQ+LSbCcpiRjNJpQUKJQx/hm+21ccxR17GnbmlQkDlxYfqNfFw2/Py
L4t0UJRxDm8afT7E6Rt6/wURsfHdtsKrsOHkDjBZaxGY2Skfy5ZN+ITagH4Neinl
dbmSR8AjUn7gmjvXtBIzttb3LKKmhZAR7hFQG6OJzJsNbPMj6EInxLdfV8tdUdsZ
5OLE5xC3AuykmmE8hAmyqj/DRRhWesYUoTmicnB//04p7WjtNg9ROKrdEZNePBXf
GPYP0k+IP4CaWTKh7IfI7K72MEdbF/qUV3uZ7yTdbAgzZlgr1oR2j9ofo29z83Rf
wRfOmcA2ImpSNXp4xHTVfN8VC8jCuE+g4H22Hdl4mCW17J6TyszqP2QDviMN4nNm
wQomsi1WLuktu/df9jcMKvimeefwdBRNhpV/dmpLNafy5ODbE6w7qJ2Bd+X0+VjL
cqbJCgslKJGYSB7GrYQPuHTGqQ2AUH9TXme2uaQn22MPMiEst0skfnqzb/B7oMqJ
U0CwWNdOXlbG8YTNfCgKl/3V6duJOgmYHHgGOh097I3mUX8VDUQigb/mpxtrhozg
w3wE9aIPOaz45nfk5HumgCsDMW1Fv26LlQncAQ0PHMaeeyBCfF4EOo4iQQb5OFxJ
`protect END_PROTECTED
