`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jeRENrHLiLXeQcTlhH2pk3UiAxqHgjkcxcISwpAFMblYeuheSG7XnM4PLFSyWYZN
Jvi7ACaqEIek2hE/fLgDCeBFe22rjTkHoqHeRGblF1O+lSP3TcYNM/qZ5XLydsFs
ZBF8Izl0uy0vEB2QxivQJlQ9vvZfQqDgbp4kQEEOhUVyCzzPbhpebHm7S0lMOkWz
KKOUCAgEOMCRAB/qH6Lq92FxQ8FxY/6CcQbKruaoD50+J/aX3zglfSueBBTfR2jB
vwE17DWm61Zygnp0EbePvELn1j3wQGJgHb3Buql9wAMFaJxLO1NdtKYQ3NrUy4nG
QdkmMJJ45LC4x/gYRtHhqa0vHDxH5Dk3uZiNB+GbgN2aDN/o8DktOt+kEMawlmCw
dpZK5RWO4nqgwVuQZdjxTqdRO/gjQelEE3QG+NAsCHrTOMN4NegNWEJubk2U7Xug
rU+o9q+ZPwUfu+PKuqUN3a6QD4Pv+MQ8QoAMYTSkVsx6gk15icotM4gL5T1wXBMM
K+qQtrXVrFSbA39kYir4LkY5FZUOwLO4UMyDEeH2jqIgmOqTs5ErCxBRn1ZXCs78
XH5cHMSj4XJxsjj9lEHzyg==
`protect END_PROTECTED
