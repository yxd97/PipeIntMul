`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ecGnPblyujmwce2XDs7u2Ev7p3naKJP8ntfHvUUBktNdOnI+ceBBhD/Oy4KCnEaU
GC0E27mCqbZmPl+fuC7bb9bYgdGskoGUPNMzHChCWbZXCRkBWsw+MJCvjiaWa2z+
CzuaMT7mcVKryCTziMyZF60Qozx8s0F+aN2BAq1HJtCgIDNRqK1hm8duz1RRFBFx
/obax3Rp6xU7+As/lRBsFAlmUnV/+t00ukuRkiWv/M2qaPvim4IdBI16OGhUAWgT
cJ+4P535jk0BmldE6B/KBhuqo9E2szzzX5JCIZ6s1lxI+Uzre1g+ZAkYSl79hFx6
7DqXjxjSKiEger5XzBJw0A==
`protect END_PROTECTED
