`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mhGiYyK2DnixE6kWSVXjSJx6Z8Apczhqhy+Fpv4k+HTcG5nevmoeawEY5Jt56r9E
q0kR4wsnBVyyZyjx3R4EELPLYna1uR/3u4fOiCDDweY/+yjLTyi3PBnwCLBgHdqN
GtF3WBUp5vStTEjPaohZKoWJ1wr4ZFDgZv+2AWzKT6VBYv6bwBZOgwUYo6anZfmY
tRRdF21LUiNvLwgWXX6coUFNpN3Ki7nlOAMZvmDcORm/5WvwMgNXukmRJJV+kpHf
FOJD1sCyG0bTSjcNbTB/iLLX1aS6aeDQXNqADZ+cPyA7YEFqcdATlTQgC32qOERR
p1swqgWGb0JWes9fzQSgxt2GytKDp2xt4HjGCpUwx76wXN6fJXUvOROfwYsP3yuA
qn5qvB5pmBQQq+bEKRR/c7PCj+RVgjjJTJwmCZ6RB4c+sQ5TVaSxSM5Xh1/nZJxP
GhYBw3aVvwqZfPP2vhgLfXLLhofRA/9uJgQIOpe5BxyR5xCD3a2URC2bnXrFV3iz
Noy78VsvL+3HAA7Dc+orahhL2oW6vUDIrtFDB4GUBwCLO0Bxc/msrMHLsgo3LYGj
PySIk/U67eeDBUHGJNuVTxPWekqnXAgRmNDTx3i4uQ4zt55zo9TnEF1tl6Mf/UpF
krdZO8a+pkUyaZldshVQ3F59lkFXar8IYKlW2XVhNuv8X8OEGJTVK/Xx/P+Rc1Hm
ktpgHC8AnGendTXfZshh7ddDdy3ullUilegY0Cud8ftzCXnSYOmbqVoutQkM/M+9
WFCBpKcWDLHrbRxuOqme0HmPQN9dPpKz3YYAZFlbtUleJKQ9+D0Q1oTi369KrPBG
crlCKUPsT+2V3BJk449n0PKWp6w0rpfSUKY4IF9dvidSmTikMn37PgMP3PmSnR6J
ScQMFvceFwFzOUgLvSNXrEoaSKrjj1ZcA0rHrYQfkXIb/l7uVRMSchDQZAhDnPbt
WfVbDMlSGKZRbqFAmEukx6CGxuJ2H3zq1V/3xjWCWoaOXVK+7M+LtiFSPyudsjy0
zP9vn9bOU7QxdLG6qe4Ig0mE8HHEynxpK2WPjVoa5N5LJwbJpZdCUc6cSao552oA
ZAQ0P7JBqWJ+emfYQsIDX3yVE1A3R1fh0FXeQ8jB7Kz2a9fVa1M2EDDEKHDJ5PWN
QHr8ZFuvjEqyNTFGgY/5FKE8sGh71ZC0xwa+fcDUU9ZGa5NYx+b2usbm+v9XddDt
vLJhDiVJPyeLC7oUIl8NWgLs+DnUK5rG84LNfKkdXRRwywnXN85bpUefYCu2+dmy
7C47CdcEd1pK76lncBpUyVeFVHQZaHcnu1QhPHyc58qsSJipReh/FIMCeTcnjo0d
02lmdwBPUfTeSSFHXFCsXjNpEDqkxZ+f/QSybMaP4SWYS0swtBhb8Lc5kfOdjtPU
oET8apVVJbITyebQomZyNcVvjxfyHKnfBAhD/tL/FcgAhmEZJPc9X7NJ02/xze1B
kZHLNFeeFr3QMZWZk5LhGBCFujLKRiRG0rGOqGLWpRopxrVg3ShC0VqPgUnfIj9x
oPX1F4XQ+3SFvLwVWdj4fsUcFaKT6Kxc87N0elTG+gEu/kka33aIwqjQFiSaQqv4
`protect END_PROTECTED
