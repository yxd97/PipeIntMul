`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KAAzIQaPuCr2uA+tOOQiqOWxEnIWFeWINmlRauQl5KrO3DTSJvnhTPcxOM0G37Zz
p8D7McOADqZWWwxm2wykiDm2XyywF05wOGK2vu3uLAOCVTn7Yoti8Qz6R22zSoWj
X+21wLQUmwWXxo6XnZGFnP+LLVU1Gg1scjM33RG2FOqvpnWdg83p+HLfuLWOdiKl
nKFj8m/AsE8bUErSrHPrxyC9S/Ot4GwucE6a/QVpUkJmLPi/miNFBK0h9C7tXhGG
NALqCbAwKlbUHUKtrhkWebM1xxA1xgfjhdcSTltYtcaAx0Q/oT6YK1QllCGBzXAP
2yxvCkSYHPWqfS9MHV+3J27TToV2bNpgCElpuxp3XE9DdqJHsfwTtLsH5kjGWodE
LK01PYOIiPo0TOZvNs4TTx79y5qd8PqGeKZT6pOEju+dIj3qT9sXw5y2YQiKSPnH
M+rvO0pdWuAiBurG7FJ3f3RrIg2TwnVNKq9BhxpDhK1b0SFVI+4hB3njpFAMD41t
nAM9jzJHqY5TORql1R9xDp71oV1Ntq9Ijgqtccf8M37DAM2DEuofmk+rbloL8xkN
fgXJSZZ062Iek59rx3jx5E1EfApESECSobFS1BuneHHRHLt9DxuB4UeIVMrkFfkO
IFsRIjzj/PNvNDi7BR+YIxkGlxDjghQ/GZKza+lILDIu2EJGT/Oyo7hyp0OIT3wB
0B5b4e65zx50amepbSKbU4zTEdWQw2gph1JmBiaoEqqhuaF+NRW2ejAq5HSftgyU
HDpYuaHihIvOfVrhd+QUEw==
`protect END_PROTECTED
