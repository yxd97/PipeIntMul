`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahW6/xce9pmry5d81Pm3YBaf9Oc433g7ufrF9x/s3lyyq0aK1pzdxS+d+GFpjxDD
f/BHzycVAR8DaebzUYcLPonYurxl+TNtfeMGVSHWGr6esgZbVfbByZBaoPrPllW3
2IrhCJs7TESLKKTIrFYbeXJPbOP2LgTRNlQiYdd4uIVYPJPKLNoZ9T5pU7JI0lMg
7Cp6oNcZv7B0nhqNGQga9woH1DNHPIyip244cokn/XEBqTLtKM0Ui8RS5vzXlDIQ
H2Bna2yq0OLEZq+E4/wULCh4sjo9hanEAU0v2DlbydYDckw64eqmSTC7tSswamZK
6Loybt/OFBAg6/ZkghCyPItTuxVtEkP5xmziTgvCp7dVj1Jq8RtTZ+z7TLZkRhfN
SoL/kk1M7pqEKXdDp09UMTg0GPM+S05RzEmCvbaVNDRXuv1PHmy3AUaSenDQ6uCq
F4soqMNODz1Dwp8wE5k0vYUVth6HK5QEpuPWCXbGECRkhYbEvtfLKga2DY4Wf+EU
ger11jzd54K3wMsje7LUoZUjLu1Jv5zjtXHhoMFsAqhAbBZW13pccIgOEztlY2C6
2mdOUIqBJKwrmUxlt49BY0IrAg5Hdst7HTZvoIp2CP2vPPsgIrCrXPCdveUwa3xa
A6UB50/GAm/r698z38EXiYg/vpwz3ksWtxJwURHs564wO1i5x3uwWOCe1pO8/J4C
9aL53RR3J7/3M8uMeNjoSaJqvDMooGiYrS78Mt6m2xIH6IgD1n9B4zJFahU1DKVT
BG/m5faXUFDfoYCxDUVNnAPmPY2cG00AuKqoCg1+0e09+o0vdHIWCwLcLt9/9vwe
uUedPS1rlhimkRELZAWZN82SGTjGLL3g5i+EgT9CERXDdURoWks2rIsQEo9pVsxO
MmGvbjvMxuerjUn9abKIQNy3arYPToltFzg3YdXG+MH25psp/YQNKwmCg17HbvZe
xqdh6jjcpwZx7151RE7aOX5SLB0sJG2no/iq0x5QFYBIF23Ck6J8AVrLMTEcaBm6
414OUTmQcsB+hfVXZ8X2oJC3hKNhL0Y3h32paOCg0MvfPnouIN8q6OJbOOlIXh26
aXWqiZPnjesUBm/p2t6LJw==
`protect END_PROTECTED
