`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmO71Bhn9U+ilbmW61/4OrJshkfzsRt17CQAUdiY3vl/HC7ABt8UeT5aRw8uj9g0
bGEokwSaN12BSxwthtOZBHrnzo5urL4farVOJrU22EKf23GVaZWEuCHxiF2E7tXo
TqqktvLa5CMiQ130cDliOW1quWJGE1u7OMy2T3im9avADniQhqfpTT352emrhSEU
/uzFQDLApooiGV06dQuc6Z7Le3WDGXYx/ybBKjK9u+p5DDNtqGSH4KECy0FGWScn
9DC93rZp3tw2EQGeaa59uLRZ1Nm8YIjr3ouZVZg2LeR8dQc5PMDKa64cLI6N3IWg
v0m0BwC5PYrliGoypLG+hPzthU9WChq7aZa9Ib/e830TlQ+hiBtptDl+5FguK8PY
+seoKtU30lmStdMz0m2YrQYDvpMkaWNIJ+yrCDNOd9jAuXS8WbpOG7ySWX+ayLau
fbtnqpSF7UuhxTtVJFfsVHpQPSk02HFU6nj8hDu2UGJJ1iLsTzUPdMO8kDz35ufm
QSXf5VzJ6MwKISPaW9yTatqxr6XBhZkiwWnWNTHgMlkrCkEC0komdHOhaSDyeDHd
orB8Zs0hHnXYaMmGkfemL9UwyNZoaZEd29JfrNg7J8h/Ek+LXhdGb9IChVA39zx1
srtsCYoSKhIa1D7GUn4GPze65ywtc/f6xvHISyTm4nRaOaRUJakLMesKZOeJVkLb
U5Ibhk0HkQpyY1zPPC+7f21NXG+TIv+LoUGVaqSpeKvhymXbpTC6xljflQ5NVRCU
urYyB2iREgYSY3jb1pyH/V4XSBiukAaTXnrSjUfbsBpBuz0oJy1gA1JPcOjE4jb1
/L6zKIFrIGjPi98ngvowk3Ukp4nyCIqTWUeEpN8fLz10wSreowULJLVF2I/DBKzO
5bF1r2DFaVxtYIrkRaYYehV25QyJdMUdEHJ18SF8XGi5kTVbgVHmaQ9wpX2r44Wc
EZm7nun3tVt/iEF9AHvDbYtAzgfwxX8Ge/phzmUoTYPaM0NIWoH9B23jLBxS8fnN
3z5tATBLb3BcGKPibKjlg8z/7jL0rBehCmYgD5id2f83eZnuLPpWjuC3KmQgrRMr
dAhmLQs8WEArDe7AkItVF4Bu9LqdmLeg/zPJyVKEBKWXEvhx43nF9fPz879rQB+G
KVy0ZYRG7Ec8cTBXqhrgzoomIWMQYYJkSvP+/5EwW+3g4usPkTjshFGtK4alpDAJ
UebYUcaaYYbZyZfcj+KBHOyO/p3bNv21HtTKmjs5pSZvx9PN7Ht2loV9mPvMY8zM
H82czT33BTrMVHCK5f3OlLhb5wA37NzMBshLnrvLYoMjX52EObv9occ9/T0KOqn2
LcAvlZrtIUCNq26oA0j4/fIkJsW7fEdiIRDmDbQ4jJgXRaDcNKy31VBcIMcCh/l4
qQ6l/vvkgXeBzs7Ux9j1cbN9Yr0Gm7GzJe+KuXImTLiOH/xg03T8CMpLaUkHGO5Q
Km4HiKZirPTuEEoabBMfATEPSOmG+QvSVYtm+qjvIjpG6pooTJ6rIag0JpSAwYcp
qWcM5j9Y2ijiyYxqWyrHbZsPAC5z8ah/sdlWCXuTOTAaxi4UQthkHye88k5DBpm4
sdarBKh28mmlrgbyvvBg/Vd+5QWJvMFrpWPP+lpaB4OX1ocBz+CgP6bWwg0fQRKB
hBPrzx7r7xb311mW58hkLZFVKYXx/PCrEPdaUZAI7pAMKokuJz2MG75hW4J/LsdT
PWw7lXnRJOtFfwMDCp6PrfolMJEs1TrbXujQ8/6+wZpWoqoWCA+5vTamRhOcdUsW
ByR/fRb0PCHagBqkgs4qrtFrlyx80mxAv2CG8K3s7DfBKg9sK1Ani7EH5qGcALKB
LPXsejfTZnmkrbWmv2pHzSlEMXpHyFQfqTXF3rGXos31j4jPU2/+EX/1N6VpnC/p
Ys1PatkEcKxBkBm24tWJ3zo6Ma2oFlpBd5HbDVXCj2LpLBB+9XqCb6s2pXU6IemZ
fP5MxsFN6KmisUL/2KgLPbEgwtza0zfSbK+qOGGMSxozorul/e/71J9QB9jAN5c3
tS/06AzpcYhX9kiIpCQZRenFKZMt4oNUdK58ogk2xqzh2BjPS4OiQRxpcHHnhDRO
6E9EG+3HaFGFMzpyMORIE8o30mIKgD50nhiPHblcWg03a4i21ABjY/49rH51gyIg
wjnC9G+KJqm76RQX0vyQ4d7TpvpMHdHOOTfUTyhxoN/aWBLqtu7XHsYF7Lc/Ts8p
nBsS0dBJ9+vdUuVvkKcdLYxZHG7ychLvf3hh3BbBs6LJjVAhsaSuTANtzo/q1pfU
Ph1n5nXs1oqlFlT7JeUlbw==
`protect END_PROTECTED
