`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0EZAtBK2C1+2Q/huXhCIaSIWQw/2ZYRlx2cxSarZOIACFbxrsWOPOB+ohMG/zi5b
j1rcT/xURLN4zY8tz6QLlsTE6SSkPwVjgLKbnZiTDnjwNPnDFLZ5kFRu/oldj33i
kEu3jRbX9/7yxNHNREloass36/bovO33AgU6JHQZo6oPmxPVB3eNDVH/frpvKH5A
n186fISy4/sDxfIUKnvforcIWKhxmTBmgYhI1rKGixSsKcFmgDwrlqk4r5C+aDVx
aBfaLb4a/fd8Qd40w56rwwbMUAi5oVVNztfux7PK/0o8bbi9maAWJk1uJTk3E2h8
YQu4Jb5vnTemq/8NXJmiQfXjEUhCYBARaycU0hUdrAEHN+SnLOdRdrUfqD8PHar1
J0gk2VvR0C62dkHgGrvYopHID249e3z+wOyrkjJmXk8=
`protect END_PROTECTED
