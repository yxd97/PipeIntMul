`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TI56IMQQhsfkD2kMKELEzGgmflhmEftvsnXhn0EZwBdYuokKoHsWycacDNGSmRCr
M7YUfR7sPJFeRdMrUxNap0OzpYB0iKIDdyAAlcqoQq4xpVonWjfHjH5+bWxl05Ql
YO5alpQfGIbbu2lg9HPJjU/Kv/dP45zcqBuErpEooTIPg2C4WhHvbH44+v2AlWaV
TSpw8Gd8K9XrYKuBH8Tfp4YC1ofUdhQsraIt+zjuEgGbgdwWzKn/gFBdTHb8Mxxo
4Xb8VW9QuagvACGpX//Rj6Syt31vY6xJ+A1yJxLAQu/8eBDolOOWnG/bK2fsnDTP
LK3ogAoCHPbufofeQTGOVrAJvrFVhs4zCs2WWE6fc94XB5c7FKjcHj2MsV4YvcRU
1hd7CFxuZ4OUcBmQqsGpvgw63sjWwdoL1aaUr3ufl+md1sOU702BYSAHco7GwUt4
tLWIt+2n+1qxK/o325NLcSgWMwGgEaMH8xBa5Rm0X6dQ5FMYY2tUHgpos9dhJZQl
S5QAPvzSmapNmB8SMLyvFRdn/rJkBIh1Nzyms5R4CQzI4i5Z8Vg+YXDcmRl+9San
upKO4BFVYUbR1p2NbJH5nLJuEDb8yMZ87e5Szfj74pMTZ9WKFDntqAFcylO9PXCj
UzZVqLDtzQ9HeDUEl8JvkIYVZohiDP6Xyuu8qd18rxI3Ay+N1E5JXLd22PBUbxSy
cKZGg+L75CTMct9RACwPNg==
`protect END_PROTECTED
