`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aykWoTsdxWs24NDjpXUeGjqYuvzELeX8y0Czbr09UVgrvBKwo8DCd+p34QnHcB6z
eMUCfdnyivt0VwMtkLWI9Lccl2Agsb0JSmXbX8SJq3HHVtapJz0ZeGB47t09aGFv
OK5vOcDb8jFsN3AgRrLViyg1zU06ybPE70gCgNoAMndiI1mwY8d740pvg5YrknK+
VNn7gNZLWnZ5noUS2f+cu+TvInS/kyUDfAcNzoCBwcEEsZy/RQAYL1cZY9/eYZvA
oO80XlqfW/d6hArI540OO6n2rmeM5pEdbHW2K9XiTH/vlIkurKpoydsC/kU+21OB
0As6VsGg4kImhPysAkyVpBMYVzu30NnXuvI86xRPwaTMCXVkZXP68TNFJp9J6UCB
Rx2WnlU8rtFHPNMj3VVvh5YznoVi2BZoH6BL6fZIu34=
`protect END_PROTECTED
