`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ueQ0LRcUUXgVnttt3HHMl8PbESd89E/KMYLnVVE4wuK4SyBRsSgNRUUcgRlhfKMA
Hk1/lX4ZBW2AixaGx9HJNxUjEFnzfLrrRvNLEs+FCs26rjMP7Do1Cs9xBrsLrca+
UsUkjrBHPXfS7/kuE5kwlMEIDzRc2KZw1NZ4cSAe2wbTirqYpmqn/UZrUDTSoqv4
D9rth1rSkxLIa/UFAs+fzEqChbjiKyOKUCt3VhXfAthPC9DNwaabv1Hmyry4C4zk
8/gbhCTY+nVXU4ioYvyIC3+W6TsIpHNWxER54PzXgjBQW2uVZCBMqmsmhM+lY5sM
n+sScup2hwoOXNzAbEeOXhd7FDifTCYb1eiQesuY0HQ=
`protect END_PROTECTED
