`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exS7+ACUr43JYDC8NBV9wMRUDIKeiS9ie++D8e9l4h8OaVEkVijR3269/pZsypr2
T2HLD54RkAR3mnUafuL4NkcwpoumtXC0lmjGt7/HdkH5JE8Vep1VcWYGzbALlpDz
ImMrXYlz0ogxaCCfQHkgyt7Yq5kYc79ApMbZtnl4OQuSDoW6JJy1rIWUS9UmoFDF
kcw2knscz8TpRcv+x1HGgJm0mQI6o8gEfRQfzxe+74FUNpsiS0WG5pDtpj8D1doq
JqaH/mFF8ea0Sl7uExghXtRx9YyX+OJjCfQuVmPhe6o=
`protect END_PROTECTED
