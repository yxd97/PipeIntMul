`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9LYzS/gLzXSL5+SCK3Fwd2ybtBPdq6k/xAezz6XFL87J/QIqBFkokJx6/2hJwb/7
82LCL/yudm1SDymEyHiordN9i8VZtTwapiXHiSry26wJC4nuB6d86xpqLpdkkJE3
1u80XYJ1M5wijJo9AMVZVIHUVGkoPO/G7+GlRHhN1/vmsTQr6dPJC5MrbFA+tYtd
TJPZX2outDw7P4CtBwImH6GbNNNcHAeVY1oJQ9bU97DpiFbfEvsCacfk0eWdo7+g
lUhucYGASz02HynX4Dvp7fiokp84EMGMzWcN9zFK+VId+bGrQB9B2XxaIqd+DvEp
feOzsCwdllDY7SwUC30vMXCNuqIs7T4hcytJvLD/BXoPt5jV02tgDCQ7OsViHUPc
y/5FRN2lDm/gkEx6kaxwxfrmJU48Pm4234dCxIYUijgWMe8iZg1FvVar6kOb99lm
pxwW+DbJc/irjWH5xnmKkbnr5I+7gp5Jkcp+KIfUFBjvgRxlk9v1U8A/7OkvLQ0W
JV6MNolq+Fs1AmC52/a1lIUye/jRm0thNsLGpZG0rmu2Pu58VDdwEKiaIBnRZmeV
f2RlT1nofVm9VboCY+0Out7F1au2e/0XSEMmoGo91wNsCDGBj6y30U2QxwFD/qcE
xQMu+gePwd+Hzc7lCKhz2Q==
`protect END_PROTECTED
