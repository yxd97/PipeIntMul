`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WhQPpvfxgxp13VG8Jp/ADrI2pN9vOndSV07MscBcWFJGr2RVkIDeu4vKVJZ+IoP+
rL7fBbjAHoJBe0oVmBjZMhRDhahAamOFdbm+2FI5XxI8fc/Lg3vW8kam3rG+Bp+9
DkER2r2qf8db8UThR95aj2YqCyriMMcvhuPv04NQ0nCjUZIuEDpP4bYalst7tcR7
Dj2ZHmHlaOkFuMIlCHA0qt6hI7joXTQ2onAaP0fu52eK/K3psxN0FthC5NReHyI3
JjZEvjPMZf+BjKSgNLJXqlzyGy0Va6KfEtTFirIscIZlEwFRGyt4CMs/D5bQjM/o
NWT/6XmCrwhH11BSvJ+EoUtscYF+TVoqfUzsVngUDsB8tY+eUnTudasikoJlJ99h
ppAOC0VjnyoYX13wmCGtzJM24heQWJvCQvKTt2LUitnVg4mrCp35vP0wS2aM707N
6RPVAoCkcoF5rBn9yb3LjSOCVusrq0ypFR6Db/pKoZoUo3BSwjr3rZb7/OGhpVeE
WnOH5CfJeztP3pCI09NdE5h4p4fhRL8YNNz1oZgsagNRDoQlXOJhCQ5lC3aEODVB
QJQ2gqAg2uhFfGGGDf8Lfrjdwpq9M1W5cM3eXlYQ7qCjFW4cy4JCTiBPSnHBE/W0
bVNjGeBDUypPuGK6ATPDVt/ng9BOUAVqY7KR/hXiNYV0uX+vb16XktUWKkiC5IeI
H9QnwfkAHbyIjIjnsWm8dKMZ2c+IB00LgrHDJ17aLbU=
`protect END_PROTECTED
