`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4jQRnas8p+496/GnzJ1XVK1Pwo6/Xvz9NpVNooXlrotIubO6UPr/5SwjkvPuw5oc
P//bCIqEKytm4sdokejI9a0ozjgABJRlv05alye5ttLtCqPOIh5VqG3GnkQqFKWs
fzszM3cysZKEV3+M0RJus8NxxK5zvtnrKtp5CrklROjLwxffN+eXrjEC+uOkm6Rr
4vJxcs4wWsNoAtJ9B/t4vYu+5pVpaoNfKOM8BHakFd2+X9YSNrkNxAQqhvriTDB0
ImJlLBx1wz7qeC0KC+S2uGaK03u5VlZsGz0CLFjKI4GNOc3CEuMw+a9iYZ9jzhzu
tBo2bLyrpy+x4pAy4whPRjsGDWGR7InxFG9lCdd8gvH1RepJoaCFLE36cUPrhn2W
HCtcW3D3yMxACE4Gxi9ki1N3IEn/ZQKLp1xY94LrInZlvqcYkwvKQV4+Msg0YesU
VQ/8hSupl3XM14oZ3xDQlkfw5Qn0q+MmzEvM8KAgXw6JsBBjx7Qwgw0B2PPHVPF3
89KoxJgfSwM/EYp86OVCjDL+UxBMENQoob1aFw2BSKoCRDiIKE2c/cpSpEOBiMbH
gYcsbFjN6mCM8fKCNhW2FsmFaXl8rNRIkFJ5ef8x6+j9iSov0Yz95PhgeWA8ofxt
op+zj8Gvg5xV+ZqEfmvW4vOrrvZvfNp2f4wxRR89WuvtFWTUhf4cGnrQzKE1m+h7
5QjikDBpT0Mqnc8xlYM4JQ0IiKAcm3u1tFc5cl/XUrH4bbCdkmH4xcGKIwgP2qle
TKm8vyjUEpd8wmV9dd7pcgPzPxV0LM6jnBE5jeV9ghYws5c+zsUuK1OUmjVm1EBd
hE2eNlG2xErCuTvhUHCLXPyzSD5boQiI+Efri5RWCNurEdYg2D3gChgnye7Pl0P+
4FOpUGjXzBwcrj4J3YlEtaIeoOQF2DswphBRTTLCV04wPUXt9SZ2PGQkdfm8oq1z
QQLWqVmjo4I5H5ejib+BgNggZo0Ci1N5wVwwCR+LHlq2KySECZ7QAEu1eDhfI8lG
EQeRZCNU7KdwsGM2+qEgBJxZfK2Hahxhfn7itkr9ssGEjyrnsiXgt5adBZIoW8J2
KekBtgncuQxt38usvLBh4ZCuBEJ++zka+JupYtjJGJWAOaaReEk55mYgN0s8i7yy
`protect END_PROTECTED
