`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6xTzEDH67W/FA488a5IY63w/lMPiR2FRO0Pg/xtLUKha8QqcvuszQEM96CwhmR1Q
f5wZcu9uBR7FrZn9+p2CNeujvpx8WfXXwvHqZU5oyrWv5gDHk/Jlb68aJt/DDUBp
Ckv90qencASPx8TRbdjWqahx2rlYXEGy/HZ2v6vpBGyvU0I7MzajX6vrZ5uCDYUf
X6osgHaoLftn+7nVHo9/acyBcxpk+WO0+A5mvKtFHygvevrRGKucDuQQ5gGJX+zl
jJfxOzLq/cylfJf3ApABl7V0OLwkz++BazP0POzTw20NRP+T3EefBZkbwRADMeua
+RBDZCABAnS1iI5MS6tnekkRTQbECP9ZThuKXNxzmTJ7+WNevbPcLqzUxYa87vw7
8940IE5ghcJ0Zpsi2uw78Baos4EGpwiRrQG5XoeoRdHpjW6rjfJejBMupY7yS0PI
`protect END_PROTECTED
