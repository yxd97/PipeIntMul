`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvC1JFS+gS0GbzNMN0S/hXP/4HsJ4bhKbUjV7QfJVzRuqjQQuicohZi0vAShxAhJ
nlrRh5BOkVAunSViikbTDq0Doo0+7WLgAHJrr3CTE0+AtyE58ngIoLKWRXnjHa+w
9CKzeiqvfmjjEzrcI8DG47uPKt7KQGZdpYXCge0Y7XCdZ+vbjN1++zmWhpJYlssL
tYHA4vCl85k3tVJgBI50+01+BcBjOyGAn0nvmHlPlrVs8j6DiqW8g3brAl38q2eb
o2MvaQwFs0tU7mks9i96tgsQMgiyoCnDB6deymyjQd8a3cN+G9RHYYUTW+50FBCz
1F2gNnb7+B8cG5JNHaBFIJwCdeBVji56cdSJZ5vSErEnvzHOmGq6jJili3DcuO86
G/IomcY2lqZ57qEnK/hiQhMcoMzkJl9JjwKci4UT4vzi3fNqdvZxC+zrBhDViqAo
JHzu6b2M/NHC4Zln/SZzf7h+nv9LDAKiLROIx/QLYsmrY2xZ2UKjL4M6DJVIALVl
`protect END_PROTECTED
