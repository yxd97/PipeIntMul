`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iS/9Ps4vc68sHj7pTP3uXm53pN/zIXhzTRZYSjhvUskKo6YqxVeF2vP+LR0/I8CA
Ot/JMDNiJGzQcjG813pwOTvwh35gzhoSzneUe89VuxIcXu38VPU7V61LbH4tnjNI
8lDaasYRdIetFaqCNy7NcAAA3SALTfhzd4wvUL9VTIkjR1LQVEv3NCmIW/9nyvBR
BnAcl+iZZOD926LfX5K9Fh01vVmXfPzDuetTbb5CfnIjn4PUsgQwcI59yl9/YKo7
3zZOHIlVQXbIludTP/LxjHH0PwJzKFJoSukv400w8qPo124eJMZpsI4E8SUsDtUD
mw0+DUF+CCijUIQ9S+qmrJrIlHNAQD8FqjU1LPrxTUxaBP0xwuJM9+W8j5Aa+JBY
CLA0pCicq9/Hy4rThXNa3KFAm5Fcno5vVipCl8IzRmjYsPosHa2PazA27DLBIx7l
47hPNK+WTDqiJhhKiE6AtppadIWzeBiTLPJ/3W0x0Ds=
`protect END_PROTECTED
