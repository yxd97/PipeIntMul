`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlwPsIqb2azkwH8tdvMty6j77A4vVvW/h3vUrvFcTNM7RLclodlajLxTdsnVgCb7
dQAoMxk251u5srQ3JCn2XDXhiB23Urdoxu5IHeb7iiiyjwRoXv5GVnLMMYFLS42k
8sU+lxc6+LnPym4lQwzhLvHqEITmJDTDojAIpCSM0kYov97cWIiUYg509dZhXqZr
FSbK9Q7QgQGEACGHyLrWJ+X/j8dgs3hB7v2F8T8aTwje24VygnusjT0keG1TfT9f
00Pc/15+u1pE9PGF9DAua8zgQR8nhj0lhS/EJuya3Ji83rS1AvJ0Q7pn61JSPbug
tymRwvJJ9FCUyODll9Lfs5xw11jSGgbsg6chZ6uZPxXq3eTV0BtBxJZu/+JZlggS
RPCylKxMQuRQ48yygtkf9W19LjPh2czk1FzN7qWWm99teVGs2Kl9QXfcEZN5dAYb
`protect END_PROTECTED
