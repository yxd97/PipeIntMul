`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jzSAGhOv59guSAONrq19a1fl8ragdQpAs+WX3bmmIzfDE/wFOW/OWw1G9HkdWbRo
0V/ckOh0n3JEXbx7iEIhiVwus1jqYEDn7W2o53Emvk+1SnIs77zxwlLQoyadHiVv
n0Z3r6xKds8PxpF75z3GTRpzwgWLfb/+ny2OHD8srDmeiyi71I9s62QT2Ls03gjs
zYlqXgU+T5sVqRYSTpDl+djXLoUhBH6PhxHLONviwiFPTOMT8baBfAZjmCD2WbLj
am4mq4HmcL1ooQjmUrybcmKiN1nPqdxYAsl05HumVHqyLN4OVNhgo758jL0lTDye
PByFYvQgwmbuOn/DFUCuanmEF0bwhVAacDxmxJNg2pMThS2PHk+ergup2JscXGzW
fjwZl6tOFEVtC0XmG7RdBPpSW/9mIla/qLceT/go2ihnVSS9vbyww/McAiT5NtGf
RBJM8dpv/BSTZpu3dmmdO0RAv7zzcxHc9qvCfClFoIudB8gNq7L76CEjPK31+1TZ
6ZdVTOXkxRtb8LZaFime1xsdtqvq/390GSV4TjZE+Sg=
`protect END_PROTECTED
