`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/5El6sGlx5mdIIyr9nHeIxP0aE2vdOQSNKYfEUE+aXUDzSMOgjuQmxBWTxEXNIZx
4CRin1fvYjVmjOM0LKxSTXTJFb/JimZQzh9UoemVk8U9J5VU0ClBe3iW5O3R94VE
BvUTPQJO08lysEhxKwcAOiH5k6PJUCz4XT/Q+zNOTYy7F/XBZsfTaHfG1Psbhxir
vB7nfZqkqWh05TcHxAVHLra8ACQ9VxrIJt4zmP61PsyQXEL8nl25OrZNzwc6lwow
6G58mWOqd5Vr7D+2SSLSWP2vgw64tE5DVL3r8gNzDvfxylTNu/tgtV1yabfTNp44
2CmtbG1F1pblEfvwkDwMCA==
`protect END_PROTECTED
