`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0lY4W3YoxdFQNZRC+WyyAnlbK9simQCzsqJLaxW0hYDA+rDpZU9FTet6MMZnQTy
xz9WJkuI7QFoeGyf+GQFH7QJjHTDxPBCnflrr+KckwanqR5brUfVpO5VDETXttPO
BQBItOvWlEWgKt0DHLkZcxiitgtEUo8Jracsu7CukQ3sBqr9gp3nYORsygpx8iiZ
pYeqLXOF2U+MiMnXutIVE+jgxytDp7GZaXw7Jtpt3HQuswTqnT6kQ/J4C85BgQm6
iyUI63zaj6wNy8Unv34APQ5eJ0bQjwJl8FDfqfXWeHost9l0C85RA/LszW/CBgMo
hkwE+wJI+RvInGX9vmnk/vCwxxRlAUBaQVU80fmdwb45Zyfrur384piqwhhIrRMW
TJXEOmsLAh1ZjznPTNEbZWDEpMeyIb99hX7r57MiRUxasJrkh59uj5ZC4Jt+wWh3
jN/AewTr6CWJAWyZ1CYT5YJQQLpeIHbYtclmFoPUvZo5T3g9cMAtFJl5enjrOkMm
+yA9tvDDQTHbdtRtm33vAgBH3kCjsg7wztg0e/nElpaV9BRf0wwEQ8PFGVRA7YLb
QRctg9oTnWnfypMn/w66gJBGoSqLx5ekJte+0U0pfpsw3sFSq6cFe82RIhjbPdQa
EEo+SrCrIo/42rVDhjdR2yxjPbO2QmwGDIJeoCoVc8obMAhggB9R9QrGd+icY6Pl
exDh/y3a2Dg90ZnHuSU4BNCHeMTzbSVzE1G/uPswhue9u+IsOfugrNLMh+da8rkF
cmlGYVJ2ycce/L+v+InAVLFR0NWVLJOQXsYdocd1o80EwOAcKcHiGhEwcWMprEAU
vCuN3a7vdwVLNhGFz8g+VEaXeHf7HPxnEnraxs4v5xmDhr9EgD9zJgsRJ9tH8gYp
BcWyJWVt9YfThhV8rG6iKoG9/LjjJVE1Up5f0P8UC7HKm7NX7cj+GDeaOqTo7lx6
1pIBgv7Zi6CkKPn3OGuIdOqSSiiVqckQRR/SYvkSs2JTsx2FIL85tq9AKNsPWT20
vMQp6VfR1QlFuKiM8opCLD2NuZeDJNe+I6PK1EXa6nDuonjEVR2MmsTIvxr7YqVb
ICqa1diUjimZ2i2+8LJZ38/l00lz8Ro2TdEqJRfWU870edTDIRbPPWj+zB6EM/in
5pnQ2Uw5FZRnJ2YXPEVcOJebR5wF8sihPYZgwVwjnAwmxfjY78TTRsyi1nRVDj1x
XrbfHv14q20f0VNWjD1+yuGGu7wOq2j6jDWr0XYJIs1kJMZ4EklaF+vJk/MdZxzJ
KQwvyQ74SiQiZ83r2lfYLAI9aQGRftBbWCZdN0i4SPD7godsoIqx0ZAo+80hiiHl
mzZ4dKzXmZ7jpMNIsbflOEkWnFBd9i6ta2JFLu3/MhRS641bQVfTZEkGXuOmGEmF
4+tQXAvzLGYm39TUSPIjqAoo4SiArXA59hyk0nzS0dYysfNUJ3NzrxLYsGR8MsgN
YfQlES7EZ92x9/uTY3iNF5P+u03AvLU42d+y47wDdcOu0me9wNPQ6yETf20u3G9U
6LIpgTcrrQtTpi6+ThTNEuZJFwCp9BxtwbZ4iXUz0ohaOnmegOk/NABQDfVou3qF
3Ata9RuP/8LDVbXTTFsql2DCspUyDAS37qh8rKCuJOoziBz3qz3d2JUYCs6Ts6MQ
YcY5nrEMaWGFdQrbb6xu9vK9fLqZkS44eZi1tDaS7Qe3icTfxS78Hz/QS6i2MYDx
ysD3D9ScXT0k9EL3lsoSWhrh2IGlqFiM9+k9zUZ/5SuYpmAdkDzXs3xXi3BgpnLQ
9jguP/plvScD9tuu0/kKnH+iHP5BlMPXpsgAFZd4ckIQWuoIcp7VV18bolvZC+Mo
`protect END_PROTECTED
