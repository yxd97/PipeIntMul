`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c64yun6+sLfmqKy8JryM4SrVaGoUyJIyESTLxLOcrhDOM2UqHBiGB0rC8jEyS/GY
hauHabyq33NnHgz0cN35NZXKp8RnesTBxBe+DZWSQDqDgymCGRplFIlYrM4XOXm2
zzzpx+ppQ5+6uOuCKhIPaleIQDj9kKVMnm6TQnl09W8djRzKMs45tjCcQFLpS3wO
vtxFqC3iRrMZxDUb6Y/iqqsH+ZuU18DGEAXy+qeD2/LkaMEOen2g30ve2LfvZwnz
PFMe+gE87aKxKCpYf8zpxrSjyzSlMLuWJLvKmxgFykp6CpDDUGlfz+q7F5om6z97
YjAfvotZCVyiHykhUbU1OvSp+i9APaN2dHjLg+VUQCEvnL8Z9nQA2eayGwN4lh24
`protect END_PROTECTED
