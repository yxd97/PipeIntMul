`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FXhMKiFV97tJK8RE6SNxBbMbfa2lJy9Tp/UwD58Y4JwPMffMzlw7M3/XVPTKAi9S
CdQ1DkZ67TFUA25sDy8QlKnzNP6nDs/kdeAaEHiQoLsb0ePnW+4fxxSmIzyCOC7n
CNiUIkrTVLH30fteq5bge6hmpkZjjJ49zkpQL4WL4kboro4izDjB/bVZl17ExXwD
nr9o6UFVpIRhdC724/xjfcukknbFm8GxwAhzTh0j9p+OytMB1QECAbkTDH7thvaS
cv7iVK7fh5g+nDNmWKXPRe4xDZTXYuryJLLMGsnea6tN/t9DRJpX3uX7Hz5WgZuV
7XSQ2kMfGXN1CWLdLYtU9bm49GiPQZwHZJH8UnWgiFmXNtE1ZfhNxPdpE2V6aEY6
84wk9ujp4HjYQHtA3voaoPnBJtAMqAUq0YJsQuTErDKWJSjh9cinGQ16KPDyBu4V
ruVSS7UPj8J3/6JJMMupaLH8FFde3xPgRK7HGfjIaBzReYewgUyAGnJXeUfmqQwE
Qu+kzmLvxcewY7KcRuLRFluNLL9WEODlCgf2sTqtCWfFUfd5hoz1pL3uOtBnfKLM
RCyZ8BxiJ/s08EPgIeG8akUvslItgawWCqRXwmNG76J7Dp2DWnYejpbSYIgKfolI
djy41uVRHnS6vWarNEJQuLlQigRcBI/4yA2LlYoU1GrinjClXiSWJ21irRGPdMY4
sy58RKPtsBEV6CXbf1RZvSqpx+Ea1UdTW4I8iiUgyWB0aA4SFRHJS2oUalBsJxzV
pIM3N+nML3JWsvmzUyXURD4bEBiIg0YBt2XKvF9g4VPZ6ETQ0eWJQtn/0HLUFLY4
tyhrnPcRm38XNvoXBzJkX3KGWnguNSKn2XSDfMP7CV6kGuni8k8OeFiZIuD8t0hE
ggTchpjThB6oHMe7AbHiM7aI2iQpPG////ZZm0tkztNjVnsBp20csF9kWtazeDJB
HTpNkmL8BCXAApVWbwzUjNMsU/uJM7JgV3GKiZnOISuiNK83E+n3aLUTj94CQd2V
/ZWWndmjnohCSPd+8wxJPkZh+Qj/SaxIcg/Whn/9FXpsb1Zul2DKteN02TZqy7Wr
gwIE2JHuXlRjUunV/wxq5vNyk6E84j1GCIdeAK45wu8EtVaPmSFDDAfOwmIMjLdl
3bpdlKsYhkZmEE6UN9HV9N4XgHbrKrrWX1WiA3k4z820aQQQHgyk7gKv9yUt3qUJ
Ap4MnkE5qGgBgSRNetMQbb/NxNTX7eT5OrXbZIsXngYQiI4tOfLMcFmi3YRhIK1B
y4X4ChcdYPotCG/H7UmMbVhCu/yd0wFnnrKjzwxCB/Q2jI0Po21i7q4zwxmKH6S1
Ruu4wb2SnmmTvGkbvFBQAP2Zi0HQp36/JdDYHEWfLx344oFjK9T6xelrjLt+bbc8
czzwDvtugcEbFg83d+q8PuRkvP9QSUueNtyozw0r0noUXfaPk3XyJ0JlXBABTuPE
gXUjRqHKbleJeRXvKkpuQ+OFgEh/4wOWhVYJ4e9tX9m8s70JsQljhkAevqfZgPtT
Bpwoyku8rIIpgXhrwTiaFjTpYLjUS1WREUNhjbFBZsC4Oj/c+MnyzzwUyc4yb8w4
0Sgn5vL7CqsyLTo0Mrl2wmh2ox+Bmeyur52xXiAhVratJrQDBf5tDeAdCJ76rdf4
vhcvJkdfJm+rbnDZldZpD28xSOlkFQ08cVaoz3l2R0xi54fuugHwwNHu9p911d37
AipdWQucCWbTC7U6RhaRW124BmMha6tMBfyBdExKOTeKOZsZUUNmZPUkaSjGff+O
JU92YKm/XhH7cT3q1gfvDTvI4KFXdzHHufHU6rH+ELT22WeOpflodlw1POg1qqW7
wdjVMDbquIM9J+xfcQb2Ma37p1gpquvNh47nz67YgclrEvQZ3J0MCFtd/yISwKFF
6g2lH9FNSIQdElM/6y/1KuJYm1UVqC2ijn+1co9zMyc=
`protect END_PROTECTED
