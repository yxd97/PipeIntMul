`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vZMN+TIMZVODw6170YEvkJOCeCtU0Jczk12cwsv0sAr3qH0uLze88+2itpaCX2ac
I65m6XF2Ck2jSOJzGooYgEGMTNFx2XsyZvF7PIRVdUsI5PL8M4u4LLjgEGbDvRaC
8Yv/qlIa/dj+c2PUGnHycE80NOQSmrAPv/nXpzVooGRo6Cxu2OCsqENVbaS+u3/6
DG8fU9cTfwzW82iq/WLvt9jGg6PkRaqWeyXswIxdGihAi5H9/niMeWaBUZRIfnYU
xcRgIJIeQVEtxlqQXB5603Lv8o4THex2CuD271C9Oeoc6O73fEM8yWieiSAKFzB5
ZU9H8817Q/qfqrhlaCNERc28FNI8acDdOAZOiKKnLsQKyur0Nrr6rInlMEgDi8a7
CITWqZ/74CTjyf/kEjWd1nbuQPLfMkQN2BGdfJzxOArV1nQx9b2EkOgWAmY28+Pr
PnDt1ZOVhEd3TDrZFIv/nQlCqGe63Gp8M7iG8QHJgfbRWdw1Y2K8zOnYUFB+KMxQ
M5HqzRctBRuZoKe90hm3scYTRIi6ntaMnFtypfGuGUKUwfIyMvdXaQZBD0ZSuUgT
Xw7PlUPYrSUjZyMfDSRaIZAM9k7sTZZEk9F27BNWRfkQ4QXye43e//Mc62tJXd28
tk+UwkpHnmnbTDqwzNqGKaCYipasKC6Dm1UVwFg6bIK/vrB5ia15jiGoNAAEA+0p
VPRw/bF1fLAI/N+09Kz9J3wh2VeX6HSHOE40DiQRJBQoIGiQJfxauidcnMuoT60l
5BfiK2K9o0hEAvdsNAoI+CN+puynjvhr3OpEYJ0HfBQ=
`protect END_PROTECTED
