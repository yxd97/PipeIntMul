`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NFG3vYYrBf/ldLxCJT9qCCS2OC3hgFpkW1YsF1qxc26yycfMv5V7mtMWsp5bnSR
lD8dQY1ZGnd6+weArnXD+Vf5syXI9dY1KGZjsyu8bpJXhL8nPFbWoqX49O6EMPi8
2GDk1+9wju/U//wI2/ozUJqiEfpLFpx5devYI9k/HkI+KzIBgpEDo4QjHU5kDkIb
h4ds2Hj5YiFYfl8aaoPNUQEZhBVTnJASyE+TjfWcbFlaZL+YEABYEg5A/HDuKFJF
prO7zsjTHR7cEST0rfgucyzmxt457NXlA9l8arrcYuW+5+jN8nDP6aGRZLl7Q19U
FuMDoGofVGrO0WtTk18Az6zxwtoAsIkLf+uvlSUHlumwN9EQHKt/24Ssytd5Zgsu
Un/30FR/3wNSmdHmDR+v8VZwFNbdHmvMfyARWoR+Luo=
`protect END_PROTECTED
