`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JYZhZk1skSavUESgZvx3gSKvojsNjhijNuZ/OQBSIVtQhhQDEBAVLQr9j9URZfi2
DhNr/KXhrO1n3glsGMhFU6JET2AxvVrRC2XKP8EXsdoZrG3enoATEID6UxK5eOr7
Xd+98KX/nHt3RYiyHSJGZsraD+Nm47QW99NNplvF0XB8g7cf/PVp397sgE16n812
CpUhoZcM6JqNkM2+nl1liJseu8SfuN2IIpT82bivu4oZXolwprcKMX+8uta7FZj2
YeP2CzJufU/e+zd84M23uxsK1h+GiFIgcQXaYaKjX8SIcM0GcuMnaZ+wyBzdqT+v
rcNTFHMu/tH3W3oXTJHLJHv06rCtq4OS1gcXMizU0JRv8whjOKHrDECB5e+QU6lD
VJoRIIVTvt4WaCUnzvwqUpL5j8+5qm0kKogtcKP4bhusc5JGDVUjFSncRO6CJ805
eaCXFoe+lvAI0vYtRalANppdjWEPiTiL3lRukZdy6jC4ok123KWdm8Vg/zc5Cz+k
0+QZIXHQplGU/PXoA6d0kqWWnteAo9BhdfRhVlG5gaBRhfBai228bl1E4JuRFHLW
oeHc73cKcvGnSk2feVrtOJ8rn4ymlWJx3TwguggbcJaDQTt2Q2ee3qbuPwOgFh4M
433QfHV7v3wW8fju3njHWXUgD43PsZBwbUbDmvOcy2oA3UrK8qWk9LES71P+XgbR
inSHEtLrIe3U8i7kbwFbnLXgPZmRGwaBul9moHmkoFI3eBnfVlyS22OcRgclMc8v
hTialu6LAXKjw9QNOdbSbMVYuJCFJB/eca1kRwdlujhkOzkcKG93rqBJA7CmXIhj
otS6jQuSkgs3rAfOytnkz8TNtz3UeE7hD5aCGcIVbRDxd95juUPAjgY8jo/c48SV
Kb7eqIsH9VOP2C8i7jNELviGrcgBy8qPMYGYMVve6DstEp7yjqpZiQfbveYx+IhQ
XGrJTj50HE81XAmba800eUZt/zLVOQLu5k6jBzWa91cvuinXF0aFPLawVT7E8Z+l
Ws2D8eLnZJscdHdCUgB1VfJAzuUoIxLxfiTvDztQjDdERMFJ18SZYbIEQ3wu8utF
HP84xkAHTcaGFc0GnJixPs3I1tt7WWiA+95JCCgDnZnOtUZIbQ/KMYTUNF88FPxA
2KqMvxK8ysIRu2tZKISlqQzJyf8uZM/vCXqoEYkJcXh+FYCiLckJXFlVqKk3VyfR
GqwFXlPrf66GAJjUc4rsVdJXju54TbF/vJG6P8lxWkotjS7vK6tUqKop0IH3F+k7
QEeSuGS2gQ2V97EU0i4LGzZJYMUU2LfFKJ2/pmfOPDroxBJ/r7mgTKc3el8dkWuA
3bJ9HqICJnB0Ir9sZzqh4A8PKyBzGKYxtvga33BrmSobXXAL8vR5qXRLrRg87pqB
5C3qPffy6UT1ealhl0AgXJzL0EPEQbKlbX80KduVoRfiW0FO7Jp9yZ1v+nYXS0Ok
hWztOxbtlRSucva/TNCVyv7X4Q9O5reMAV9xdDBXPKmvyrhYZN2NQ0KgXsDI0ayk
D1CmGMo7zx7kGxhlxVKwhFayFN/Jyh48x4znESmAm/hOcqhoWKCxvPbVs3C5iaej
2HPkFnEDpdtLbIzrFJP9Arw1na4A3ujhTzfFm3j+eB/joOfwJoKFDYl09whEQefY
O5f26qub7hgV/VyETVQTKBx0Y46oDzB40cG+KkCqwo9kNTx5cezU2dDw3yykGdBT
Osbj/9iHFxGUxuK5SYfT+Nn8DrXqcWaOZq3K1Q/u9dAclJPf34gkPMRs4fcnd21U
14cGfn+PHTP243OxoZC/xl2tws+G4wYOLHTAEValM1wLVwoy6Q2e61K1/jKr7Ahj
9PQlk0f19xJwEX67CPpSfE/hklEvVHrZv2hZHmhoF5k8GBTGuj1b3EP3Xc+0bA6o
5DfcDnJvGKtMG67v5k+l9nlV8P9qN6HgnSN/efa7StvN2E1p1dshCzrzJErvtQff
cr7jNbSGl2l7Dm282Y09zyxgAd+2IAjR9cgCTNp+uwiepqS8xNm7K0NIUliGKzPI
TPjdIq+xFSb5DY3QVZ1CxJUjDdPmV8GYQPuoasGJBo2HAsm45PJq92GVP/4ljI7m
jNffZNJ69Ee3Nsmr++v/EOLdULxdX/TWxFsN0mgx4SIX6MQ7Qhc6uPKQWdd8l5qd
9Chu+veJHstY8hJ4dqxZd6Ct4mYFriHAe6faB/SF47DkpDO0vFtyllQZJaHYKU6F
EaKnn1QBeBFPQCpLH7tkfXZBhlUNN8Iz4jOVcc/NCUBJHB/r+VUhtQfJqq5cjKHx
SWQ6X5tTFLMIrHVAGlLfz5JrJSoM9okEUu1hxD+pVmhxsRH14pD3D0NRLczVOx+W
BfrFfWWrEdTx4c+zo+KHCyNy6wDv91xdzNwJkL/ti+GbEGLV+l47Iz5NQoa4GEaY
u457glD/haK52nHdi88o40UOftaPFkRW9u77zOfe44yAETEt5+QHlFLmBMpmQ7E3
6e+tRbHPeeg0ZghwAm/n/1QCSP1RpIJGzFUADjxN6Q2GhcGHGojo+MAGTUKg0d6U
HAM6pcw7MuLmkY9LPqlUeVvZoawHMW2s5s2so0ATWL5KxWMP2T8ir7OpN7LSiKA8
1eba5N6GvdevTMPLpHitwhC5yaERTwODSo76Xj9wHjECvslXkUOaIjzYxv38OVC7
LqGEfI23GI31HycmHM/BvstbfcS5SRfQ53AUT2vz2wCyTYDy3rvRbdgmgCbu3upp
oEBGY4+oeh2BkS5Sa0r3VNnCv5g67I6No9lcPtxHcoXdTskHr47pUaOXcmtrGeCO
TbUT9P3pH6nnqB8HyvAGdjz54XILuCOHgmcqJMqOFWPySyxVQp3NGlDXJkczsyLD
xIN0jbxE3R49VkudaE+qn7AYw4YMpS9027sADJtjO5o4YzSzYqMYu3upOEKmGZWY
94xB15O9oMLkaDTrqijyYSSbpbOc6b4GnygrLAgPALnNKWFkNX4umhOt0w5Mo34H
PTcd9JBBK1APtvk1vHSKfnXHuGvJJ/uraNU7y8glH1qSKJ9hr/z9xfJ8vDb1sXO2
K6dMN3Ugki/e9IwRph4M/gL6KAHhguwSHNx0S/uh2Vo5zGVemiFfTs93pEcOjAZA
dNgoUJ4qUwtZD+0wG2pS1LWkEqFUpzprlIqU9HEVIqEZEvU1uXzvDtcylox0eJbx
dOBEJw3UPlAl1R58iCBlph5QGITBuIfU3fPlBRAJ7Z3BvdJwj6iahLrnrkwFaBS0
JTtreUB1OTYT3W/KwQzuzu5PfXIF4KI2rk0ZdvliiCBBP2c+HExcrhBJKVwLJx69
FSezQ6B4lD1tpq0BpHYQwM7zs93tsZNFwkSBFgIxWJD83hASfHCTDx8Xzv9ShNhs
bneQITI21UlKbiWBjxN9FKzccPRMdKsYjCOq4sK0cfdBBrtbAiy0pxaBZ7A5WB4P
zRgncRdYOm7EKGpYp2Jhoedm978n4R3RFjH0BOYRPSOvnHoeRla3RxhEi/rzVW+v
+JYu6yvhtFtp4As6R2maQoF7Fd73je36NGVIXEhKVMvkYg+UKmjN85jXX2YaDGH0
1Gv1nTHY6qpQ3MacrbuBtMDwGRIJItiuFbs1ndXnp+m5t38pPnpOuZ0ntvaGYLSb
Dgp6TPL9+C+FlNbAockwLPQgSdVxICWpQb6XpwtHQeQfxHS4kmJgMpUufL+tA1Hk
rnFpLtxDXphyP7ZFPZUEBwbSGB0R+ikzgo3jEkBj2mH7CK0DpGENPrGnFrHvpet1
0l70PZjgAI0+QYltHO0YUDxkanz6zH7Dt3dIN5UwA4gccDZlnATeuLmVlfKrY+l9
lydxL+m5MoC1EXIJ9xzrH1g+mFzbpcry2nWNkzIiSQghvZlGkrpLUa6TMfNEx7V4
jcp4Slt/apWeeLqRF1Q0xnVnhTEntpRQhS4TTXJhSRuOFzppTq2/1b+Uwz5jw+iK
SEFEOlUuFU2AOyXgfyQZ7suAnBf94wuxmQ5w3Soqju4D5bBUtCv2uqTvUAFk7aJi
VdwJeCkDto3jPpYW14yAMTT8oRTGHKn/ipIHz26GTDfgGTe94DFSy6K4Qb/Dkdyq
nvSNfwKStoYANBy8P4aZAe2FwaztVS6rPk5GQKwOedeMIPXAPuee3rBuR34j68L7
djMQKRAjeH7PSFSSrH45ckv7MPdIUjKquFIN77pW2yT+m2bRmknfPLA6Pxfd+Hj9
d3vdafrbnXx8/KNmduVKAjw2ztQlAvgEpHuWrj+AtQr1ua0c4uXyWAI6hCXYK/Ys
gC9TjBX9ZM7WzY4yhAL8eA3MC+41vChfVLyRzBhczybbmsdjQ615g/8cG8vICx1Q
O+NKcQqiQWKE7uOAdpKHimyG8MjJW828Zph32MDOYTpz+DiVDjKft0bn1techx/0
NDjCe02r2/jlFSpSm17uGvxqA8DD0yvf48Bz+5M2s0JvFxJCdvhaFpjwJqA4xA4N
+I0wudlxG0ra56xHo+llbZfEoIw4i9yGY5NhOs4/z7GH6eA/c+klh43GPdDuv/Py
7i5CrTfBnIdNGmtlpD94QiNBO9ulQAyrovqhTQagjfIzLjZWCfmpadWDBFRpvbvk
2pqIAV4eSfYpZC0l4HUq6nf0sIFSZf5mUM3CUCpohmZ57Y8Lyd0N+qyZOV+ifXEw
XND6BGv5DVVss65uoYE+XSv2tiSvZRYklce6QP7hJP1BHsgz+UwHQy+DbX1KIwp3
FoGmJ5YTs8dDWYYhL9mD+YdymSPJXVBae/+HVIvECCEOr4cTqY164Dh0E/Vs9tdd
7MX/nzfmfOxEQ/xMnEUpTZYozwpjerNh+VVs+fYzX1kwxwkUyyLtfe2SBsgBqKgN
EKaPUdG1JfydpdujmGv7Q7UaXy6tvMgQrRtVRNECgdGMM1C7NeA8l6q4VEpDWJoc
Nmzl8Sm6C69X+hHtsaCnlqoLDVMNbBWg1XM7DDnreHC7BO7JJ5PX9Xa5AtAgrBDN
l8OS09lKH6jlPKUq93rgjH2qUdti8zFQ2uDdjlxGMQErjI/1EZ5x5v7Cx5+VXui6
eDlYnINpvOl5JP4v5kIfKGFFqGxVM+eDSq14+I0dOGtduy7VrmYLU3S+mRdOdos/
9zq6R/ZXhugWJSHJYbEt79RysxVjcrFsMXZN9MjypQWJmIKBq9GexstIFIw7bVdL
m4y1WZPpDO3t3oZKzNg5+ZbQOdzw9uWg5G36PStQW02jycUhhEmgimVcdt20POE8
boruonlLhmdN/Ck0lTE6UgiyKQGPCxRiR6UnBFcHF6UgnSScws71CWfLDqFNFCNn
hPhUthCEGYR7J1IiNgZ1UDic4qO+OcAsT2ZjkNnVr2kJxrdQbY8WHbL3w49cTwyF
SCd/hf4in2TmqHALHt5zKeEkgb+aSvXagb6Vy1M+fzGPx01Cx2vepTcX0/KleTjH
CWcJIqh0DXdKRtU8Gm3dgmHpcwyAo4h+dC0GujCQt6gbMhkiTxtmwUZKt5qPzK7w
l8KdN14Q3AXyC/fGvxQUhfm47fUzrW794FjsepF/WJiAgk1R93ZClZeqvN3a9kT5
2dX16cjRs23vBdgmuLWYS14cxltnWVl+1LFpN/QuwtKE0XKMunUncwbRRxb+x17r
lykFzNpGCfa2GCBaQCPLaHAPpwPTIBauZOeZlX3oZqrZhYk58YYiXO9h/fof07hR
OWMlErXlbxsRWPcnRPLl8T/YCuMkDYNYz1VbAEXRFG2Y3b1SE5fWH/nM35ZOy4w1
PM6u+eTUvCXL6WRny012LIADs6iO8KwdBfQf8I0pbCuX2sE3B4LHjcC/RcKsr5oK
SJKhXNmASM5c6DNY4oHO74NqRKfppJ29zTOByBAIW+ZOyWofgUWWsK3a5I/9rU34
XiRsnO9wA3UGAZPDl7PE3MEbLQiZk4hcnffWul1D0fBjkCnNBoCAsXvydvN4VuAf
4FWQK7iAUnDUeg285JHjzp1miibi/WQ0VwOSLvL6Iu5aIjWwMJCRAn3OJP8L6E5u
CXn4YYm41/DYaZnU89OMpp9eiSTeHbKX8rH/1vNgERhbsKGX58Z/Fl2Uj4xiehka
SoaR3T3mtuckfKvoYs4CPfZfQYkiEpAmdZf68ADlUmK5ptFVkvap12OBSXoTllkC
Tif9xnx1IH1JKkd5c+AaZytcWPtQANeCUV38hIEcKxXCig2M6d5AiklEH3l+xmUI
ZrXo/xRqOMhedxStWGRbiht84lun5pNI3dxDh4ymgvT8lmIZMXGyDJVscVFht+s+
b8/YV8WiMA4KrUAJAfyhJkkf9uuxl+KZDWh4YfI1iudHtKW5oDX7QDluTWeXPX8A
B42SlJptevYvGbZv5GS0y+/XC6mSXWfK2ialbTl0NqhekXNHBYlnVBdmW//RQUWr
UPasu4Wl2vfkBucNOKWesp9F8NTkQCAaZuBdwESqUc9BJ5EFhna/B5e4tD/lAwAn
xv7C9LrRnzu5N1sjuwtdw73cCJZqO3aSE2WxaUy/eOxdOkxJKQRyF/Ry00BleJSQ
jCOwhM9k5pyd5ls0Qqg2CrD9sSQWmPUoQ6h3Zv7s6q1ptacYzj72/Z5NSzN99byJ
rccEOOfvvf/96n362/b3kjBsWyQxJayvBw0dY+gPLtEOwmVFgeSeeiQxre+M9WlB
r2PHUQvl0CS2EnIJCOU8AJMOyNBGVoK08uumyxAd84ju/Ge/ODTguYs6+eHhR48R
vfIERwCpcTr5+Gd5OTyPoNiueZLDt8L74zS2sTjf0kLzDRI8OL1c/EhK4rGM11zp
ZLOopMZ8YzK8RZOdbMiopdMzTLnZ1s7Dkmo8MYJ9RdtoIzScmhAxfBPjF7uxIUgP
OfI8S9PorWgOxEvRxLmLQ4TDO2PAci/EHcjzRpG9COVtNa9z+jMZkCNzNfiqADLu
2RECDOAuq0ceDLU9UQO4QgZWA+3ku9+nJs6Q3wIVlsHffn3NMLivj/Gc8/Z7K8Nk
RvlmEln4ko7SVqspKOdtphZ5AIYzSZuarsI2Rd4dzCxEIWOUz+xkT1rU6Woxb4Xa
Do5v+54hCE7awhOIp0aYL69kMbfpd3RNXt48Offe8X52sGoKOAMnrMfg/XYVaoZa
KLBKT3UZZqSFFjx/byH/FCvBuh75D6cYN2vceenvXoeDTqgOJ2ZpaMJftBlNUyGs
KU54EK/G8vSDmtw8sUimOO5a3KfvTp7CKMFO3SuCuBv6tybRhNgClrYQF97umeTx
2aj0H1Ns8ikHJL8RWflsw1fzg1czPgPr+sH48bsQ7RhsbB5DBc35PFVtt/8zh9AJ
543mTSdSqAWggivpb+LUr85+dHRKTyRgdoio4snK+m+Rv59iRS/h1buCmN7CT3xV
R6bVN4bFijFd4eHtbKzm858NJbddrGZTFwF2n3xskENRh6Vxj23WptgK538ZRybe
zvUcrBHLdrrgV6Qnw02RObG8ki7QGbrrN6Ga9d7i+DrTnR+9w8oQ94uLiJlw4o2z
aXw57MOAnZQhjKRETuKtG7ioAX0CYhQWi/7T2cmEtZn0/IO2BLjSovKZTeNAfjqK
d89u0oGhLEqhZeAbVMSbDSJygpIK9aihQh/5AjpFr7ZUz2v4S/pUR3sPc59E3+5n
xFIPRqrsvnvejqJjIEO1ebPREjxjQCZ+u/ooTuABgreWqqd4vd/WX3I8zlWpN2HA
2G/3151Z0FDBoUS41FbX3Wa+Ioy8YxZBNFImRpMV7DGnw1kZ1pNeZZ0kGu2AAP0J
DVStaZ0fYbdzsg2CGvNh/YsSTlhVTYRqno134qi21Fhka/edSxriqnyCILilgUrg
XzLz2a9a3WNDnRste4jhj7Bh9LHwB5fIECamTArsOavW1hzUyKUMMeGb6aLFjF+J
GQs+jjLR3AxfiovQWEi8xQ76YhAbDo6SVizKWgewd0QpZgF+/P18HSdQM2t+BGQy
bMOIAVuLIS8b8bwleYmvNl+LIVWr2o+QHmxLsCNsywihtAq4CG10+xVoZOFvbgYo
X+6IZfFYpY4nXueFBf1Q9gzEFj03/08Kj/yUWoKQ3CncTp5qb5DdIFETuAH7WXZ7
SXIW2toxq3yHS04uRtQzMm1/+0KIOpvlBeOrRa+bv8irpcxUChQkClW0h7uK3GKL
ySS4i7KDISSTk1CFJF0cu1ktEdpvMtN06oElvBcR8TNUeHCydjOX3PlR0lXf9lS+
+bXx5l+JEa9itu+NgK7hNEIDZIuit5fiTOizG2nqxszf44MQHls54xlFWddNht6N
5OO9PlouE96Zj/NIPyPa9B5/xP+XwG0aa9n4xs4BUSrAVc0VwhNUCYGvsqJi7Tud
xb/avrg2jpGD1KFGuYYtCZvS4KMYf2MZ9UvsNSD4aQhchB5XbfelWvNEzlpwHl1n
qMOWbtqaS9dHmitLLoWN2IIf0tqvXw+ldcRloBNpfEL1jM6C6dkc3AwONMVOdACN
Ooj15iqvOKH3H4/cfACUtooQiXSFQnlAGwevfaQ1Qe16zmNVj2AKxbBaP7ufywT5
CMElyjmddmHpYVe6H2mR0ChtTmOBpos8WNHOwwfts+3/OEkaPJmwHfwj1KA9oKpo
cusWx+qJo23grdtIy9+BYrVdu0Cis1NX2JfahENuWU1jwGxQ4nuTX/eOZK6bMrXW
AuJbeltzs4l0OO2dLNrmGU9J3VYt1TLFEPGHvTpJaLSM4DxeFudjctAd/udx9CFI
idTC+y4HaipjFO13Tcm9bhpLohocJ+9PQB1wHgzH9XMK3TlKZ1Yh4ATvmGqhW7w9
YHigjblPx1ca7I84ffehIKTSeWIgiGN4PE4MBm2aCNX6bst8NoGh21kCEe1FTv/u
kY/oD1BHiMOdwHiW5vG6/fHtehle9Vmx9MckI7xR/vs4ChwaXm8N0BXJHHIH20bW
rNQxhsZR+SwXl2g3bkB43Oh1k2UMCePTB5dGgHnY/+h5borqpl4Gs/gO0uIeZ+SW
7Ju8IAAkfgWdhQaUdXzPguhhOdS0jqv8kJOR3GrbTkt2nzsBTtY+rIr9i1Liudo1
WvfIThIyO0Tz92vyp5z77ZaI1EMGpAMc2/Y0E4O2TWRDvtyX8GERheIQir5oX3zt
q1iszSs9y/SWKmGgThawmKOXack/RDnnWKDPk7p5Bw9pgeYBtj7kez3ByymO0uKi
0iev+kRTDJC9ZDv92u50jAMZtI/2i1qeg8uhgoYET9NEqBNih4yTqFnvD4sB07i+
aDHtwkyr9tvmB+zZ+GDBMA0WVwCkbIrqbas6ysHi3s8NedNsWA0BZDbfI92VwmwI
PDGOJHDFhVtM6rAhv93a9AWv3KjDt1OoCzGuYz0J8Ajz69GlGTnV17wvJVgiO7jU
eyAysvfHOflAopyWDj+fUj/NnwQ9sn/R0QswGtG8Jhss3VLpr5YBz7OCljNPYLPR
i+jivNiLvlTd5sstWDW20frlAzS5rproV/UP1v+pXgGxRbSZibUy3f8fZyc9miMB
U60htsqtedALGxzCEj6dzc7QQzdF5l0GgaCRoQ7xP6iTP3uHLU0kGlR2RPnM6Bq2
G9G8Dsx/Tvl2WrSmpGgzAfIt50eaddjidJTmJr6baV2v2V1QqiYwoPM1mTbI5Uby
DEAp6CNEZsTGmWdhpj+kWa0YrmaDZUWFrbGY3IMyLuTCQQZWaSZ1x2SVMBvUlTLB
y7rL7nYlprpIK0ry7xCospfGGQD3LNzUod6LkRo3dAdPvqNaT4zOrE+DP/WcFBAq
+3zzec07Ni+vJNvTFVWR0y91GADJG1zD4b/V3aepDQWqw6xeCaydJaVlrvrXL1h1
DCwLVaptnaJ2JIV7h5qQSYVsV5a41t8p1nCjtMjJWLMKo7p88n6OTVjzAJLEzWWP
u5oD1AEX2LJqvBNK3Y2+59Vw14MgfaBytosCWI1EgeUgRcO5mqB/xvGgAVVtM7tE
ui9h84D2ggRXlQrB7zLY+yiuB8B6bUzUEwms0DHH2LzUUePviNj5HEW9dOmImVFt
Xe4VOisMQYDl42YPUlpuw7yj8S8ChkgZ3UYizsnTZwUrfv2VHL3Bns0ASN1z8GgB
1HKnO8J6gF3SzDspecWl8XjVVHxQhnWDqT523KbcuuKHga8Sv/dc2+mMin9zF+ly
KyTbdrfoVGoJSNgEhkHFBK+IZW54X8DN4VG0Go2DSUlf9H5+6P65UJ55PhitE1HC
G6/mXTn1HnP7d4OCcQXiixLL/jda8etOrOQf7jH05mh5U6nQ5C4iOkZ0wpp71+86
A3uqwU/S7fp28kBoOvx/bLMBGqkug7JxBOll/IOyQ8i88O4/saMvRXwZSM3jsC8G
34iac3D3ghnKPcfTSaZeWvPN1dBOoc5+xX2GsQHFZKP+ot0fg1wnAjRHZnK/8TNN
QAYFIAVHg4TF268v5CbS7g5FK3hcwinJIjX/aQqZ4wf/kBDBZP4wCx2gjwotJtp8
bDjkJ3C2X4B7hrUR2GZWj9Zs7EBq23gvj2cqAjinDPnI95iaxVM3mOkM0Xwd2ZOj
UqcN05muxcFZfB3VtjGgAzb9blEyL0idGdgsfmYbGrXfg4FhOiSKlcgPfMuH4jbK
YcGEl48QKivh7PE8Z4Yc0u1M2YJS9D+qWjq3H3wtNE42Fzb3cAOz/7dnlWbpnGj9
dR6M08uFWDFbLefckTjsk7eFeu2z2wPVQBc7ao8THwqVeP/4Ir5JIqb5ymXGth3e
ZcgM88D49v0XHdQ6yH8oXE84pmyX1pDzF4O4nei26uLv1FYqVR3o8TjaWsMtSXLg
zgdxHi6xs/xVblP7ACM3L5CwJ+rJuKQgqvYdc9A6Q4Xoxy4kSOfryXBZehzXrR7M
OLUXhIQoiVLwpyhuhG1ZMgsvnCHn1fE8gXbKy0qTwFsM/aJ8KQupFpauEpcdHtlL
cyo2B5te4yYfj/LQcvvEDmu3sj0S8xUX19Eqq9F1y8saNDviRjbDc4sGHx//7511
g8wWdyfK8lWAmnb8u4onCXmeNna3NHiFaJ8vb9JaHIZ3KgX/aA/gZEfJyYO1WVcl
wQRNAv/uw511uc+8bwHUU9Wc9xkoS7lUx7ux+p7r9DxCYtA+jQZwaFNKpQXre1a9
g210bdYcGak3S5QvNPOYqAMVBAQwjdWAkDDCXlpHX20Aus2jV9Rigg1u7DY/ESwT
UQsgg09DSz8TCtGJj0XKA3C20HgnfThElo68kH2niE8sQRPDWR8vBfb+BwTaiSpn
wP0bNKMpJ02DKUjZ8TyW5f7PaclFbo3kmyctK4EniKghKR7zaeqEcS9hjkKaNEXJ
BoA2u2QeYoN8X9q2tEiZxUoUmv7oAOYxyVCCajt69GfWQub2PCD22y6bDV+Y3lC3
5DgY3XgCBso6QI+avTclhTCaknvoiaWTS5ERFkqNigJaLPS7KfWuoeDq3UQ7E5mt
yy/4FOpYQ2aESN0MoOyoFNsm/jD/b3lW49+HLon3qX/VoLG4101/csWSMOisLilB
Lbtq3xPxy5PfHDcqA5ECnty9gdOjk6bvUOrJn4pMwMkq12hLqNGNCg4aHBI+PCrZ
D1snXOna662gYOz1YIFt830FsgDRnH0n6EPMPikTHd3a0jB2ecqW8fvtbLRTuXik
Pw0SKyCv3NPgziV1WkmORfdrVW6B8yBrx2bn/VtZNWS0HkGtEj5p3Xykt6I7IJNk
0sL+gJ8t/OUNd77jvk2eCWQFMoZAukH8LN215dInWiYURhDmTp1gKlQQ232276Pt
/78dmkBxOuYgR4Xejt3UZL6uruVW+X+NqIZBFyUp/QNUi1ulfbTyIg9nOQjnJrRr
Houv+p+IVmonBsY7KFmwZA5QUYli8fT2KTW2SLaClYq1USxHG5klzzcEve+go5KO
ijb2HFBCe/+LEAhiPYlrFpPfM8cVV98a7jdoe9ATGR1/EgjzfrEIrrpxxAdSvdG0
0Tr0GQArNvtOBsfcsj/XZWX2rpEasvY0ydNTsvPL63yy9wh+AvyuJKPe+kcp5Vm1
a8bib9FNtvZFZF2yJ+EyVQy/0lnvGcSbJtYKR2TuOgX4oGYtr+4PGcvtuOqgC8ei
60b60kbw5Cs7y9ru3Ro9ZqtLCoyDBK7o+PbZDOOiv6ONtL74NUCrTTd3OSgvTsMh
9q9pUOLkShmHXvsQCOisCjfDbm/dN23O8fquGQA6dQXxJ9cIrmDp5gjlL5hjcffW
yzytk1hcRMHwNvT3zf2NIkrdOZ3ZYYSRCF87fOocLpqNt7PnvWpCZChQz/hw3zmP
elZoW242xpLQ4kbNTMM/rpbS1790Qkdkg3Uen9Wt6w0mNIPaUeqCFo3kTnhcjCgd
O8BFWT/ZdpmJJP/FGVczxNTzjduBhs4WL9hPU52BfGGEebqnluzGKbvddn/cBiXu
1e9/dFjBIns8u95TV7a8ktF/UeM5qzYibG9NzaPqbZdWzonWP+Ekb94lffGXCp2W
qkmGGm++nCuWEsSCKx0m5ldKGUltS8bqKFN3SGnWgwCZYWcM80viGyNFU+VorEr8
gxSna76bhai9fy3/nWNxkJKXzAHwaHemnHtuuMYR7a6H2JNX/2fiGq38/F0afwY4
Frnx7WAiDZwpHJ6vMvevMAqty4+A6iv5HrFWdrSPMXB0s1WIW5TBs2lBlzK8UVLg
YdGo6C3L6tGkhN2p7QRsM6ZSXidypKeqDpTGSBVabbIAvQ+J9pIaJcD5ddqsEc6q
4SgPTiBvVchThhT+Otu6vV+jZZ709MJUFRyAzZhbyodWy4T6sIoX4RYRi/kgZhYt
0FDLC7zYrXJZy0R48uuWJ+sjeFBsL265mBfo2xqKjAwLs4o5eDl1yTE/G+6YABt8
x9goj4RUYvjIidPDGGQ1xNvbmt/r712nFj5aSw7N64BwOa/RKY2qJxMrMk7Gx/8F
w7yiD6tonbjfEaHdXJ1L2LYvhNEiS8dXw56lkip1VuJ9ZsYJKrv9xzz7llguVzo2
m2+P0KrHD9JeKaa8eVPD4HEm+t1PVC6+O8Oecju2M5RtZ9bw/pBgJEHBofWOX4II
owCH//qlDKqr6mlnbjaHk+HAh/zrkYdMRwubZK7Uh/qu0aGjBR81qA5UEX2PcISD
/GEz7/Xbxxy0d9MRcAvJRrmJj8Ct9z4K/+2cmddFnQInr1OfK3nBz0R+J5z2evO5
9vcM41sitDM6VBk/lNAMYBTvQDyttttzFm1l67swWTTQU6IQKLqY/knaPtVNElQ4
FavFFCUO9GnGLGAqs000ScZLHBmYjYegVJY42MH5P0WXj4tt4d7r9OEfO5UnnSHc
V1tgVvPxBBJQxQqHMtoDFTUtz24ia5Iw6ewU12rqJXeRYtGg9Nd8M8Dk3pkLEAJE
4ullpj7KJrgrSALImxUx98RgeL8daj3HVxfKr9C13xWRkkJ/kz6TQ6PFYjxOBLUJ
Bbw7LIykJgdFHI+wdsYSzD58vOoTH0tRa2pec5jCjqRw9wTWWtsDsfHpj5zplMQP
3qmPIsUG68/2svI9LsM1JhQ4b8djoyqgo24kKrlpNly+ndFD6G8+W4hyaYTyRVpC
S8nvE4sqhoLQIv0qE00o08ndue/3JyRDz8w04UypQDnFzCwZuvdM8WxQ2Ic4T/9b
MWlKCiFmibuV2lgOESUVEC3teW99sqA/3iAD06vCVwBg+Rp9s0jF2cYthS9nRZEe
tG4rPwjmPqpC3XadDUB8mJlKeM0TraVDjX3y+zjMYjWpJ9Zg35w7NnBeHQELXhE6
XN93RDEvLQoNq2SESx31CQjdezh5YwRxiu8kNkBvxzc5s7RvODOtxOhHJOdus8Xg
sV1LOiGj7iW/HSoKnuLjozrv4X/Vx9Wu6uxUTbx4bRYRYNikfJBtwuEOaY5Nh3eX
OF3lhB/QFKIDi6i+ftrk2uqsLnFIgQKszoFRFMPGv5K8fIH2pf2IhBDYpmb5NWeB
Q4omFi8JMMG83iKyWWIgOlekyxVMCAFS+FwrilJG92mBKZFQNPRqvr7sOQPWvayk
Bz+TawXAsvHIsb0k3U06rZqz5mPGjPGsHJeZjCUXeTJ7XCP053Gagg4cwA52m0XL
NJ3r/l7FJ1ZZfDPr5mK+bOT1LNegGkXb8jLoKvoF0egQhvn/arH9I+MWEVdQHXNh
pKHJGKuF59jfZnYCKeGVsoqq221T0QSbnKTr4rt2sEfxBE9wshlgXZv1wfpfpPSI
aKmf4S8H6r1e7V4YlDiia25091cQws7KE20ou3NQopO70keuZNH4Vl6qK4eFxAEt
J6HTVDDvEL4vYQCQ/+xkySqiK1skvtYWyjfNkcJG/b0yzSHcx04fIoi0P9+QdlT4
KLZ07ROQ45QWRgHHP1SUSjzVcydr4Vr8Cusuf39heMykSko8WSA2cYy7ipCIZuZS
JDla78laOqESjuxsQP4CmuhGhXoq4DO18Ep53vM5IacGazJub9n8S8r0iTyn4xAZ
pK+G0RkVXoc92m80buPehzUYQdmcW8X/asdGalCn1A3hX9WupoziHzZoRehjMpWF
L59vQJattf82QIW9SvUDKYRBpSfHuEDkmLvBF2bfcb13KCZmrHyml7KDbDAMi13W
S8Z4fYq5reZOp3Fir7N3YbN7N4jBHjkFax6LEhPFxvFVPI72A5toOj+ndaoy9izr
P+xUzf3zeEezn0GWXBeqBGGnmDc93n3Ji+MNf0f2sNc9YO4kUoKo8URqh1AM00Pz
oXkwphq9X8+FbQ3VqnyngXUy8UwiOoKb1vHrgZwYhRzuiCHfExJxUTOMxzgCq2rB
3RfGrPkDHiPMxr9L6xuoqe+i+6v9IGklYkZXBh7FFq9GyJMCmDjJcnxRtnCezlWE
UvvLptMXDm1bCjLde6YeSWRnsoAPYJUa1qPKcRdjIeNEkcdwa8AqdDEccfe+a075
JpqgizF9Rrb+v8rwd8smpa3JL4Glymhs+L2LheNRDYJDNezvu5JiYNrIvVkEsi5U
HfClKMOg48oHNiCFLqubiQCPZUz7+BtzbFw1JSkcY469aQ4/eRY+BQVquJ+eY+I+
MDshavB6/B07fztPQOzVJ3UFUrs4DowFwWK4gvyo9uFXFkCUP1MXnCpqBsf81S9o
5HPG99iGvRbmM27XOVUGHqX/MXKji4O4PxD9AN3ByiDXlFqQranTxpIiGbyGaHKH
dKMNR2omshNzqeHw29BXWolhZYvUSTGcAMgDd491aGn0tzz9RmJgb0z9r7CpJpuw
D2OZR6ZMjee4z4Q+bYxdIuQf7t7q1Sw0Lu5O2ksNktcv/+mBvTK9qROCwx+V4ZKt
CRDJ4s3aLCvZhHneBwTewq2qOnU+9akiLKca3ab8kGuUsxVkv7rcpyJiESyRgWGz
Nj30dUaCofK7iWuifaO/f/2ny+XcvUEJ91MXlqbmEiDIpjHk8qq7ZVHcnjbjNKjJ
Md47D/mUy5w79TFpb8T/IUyZe0ioPUgMNBEaLO0XarBUjzF6in5NSd/EMEbLGrxV
HD1xgPeCGzkW7qbRE59uCKgstiPuXC0RAs4ATLdyjRH6VMFty8Ec1vQCuF9RKKbd
FRG+H1EhClG6usJgeCiv8bDmrbzRMUP62ZPIZbNWqBlWocbgHR3pO+qxyPF1EOT9
PAcXijfxZsLLHqC3d64iAu1i6L27+HXeAy+d7eWu+gMk1+vYD0r9fLWbRrgz72Kt
xldADvFPiSqdGAq+FMmut/6xdB3xjtl8Peq7Pp1Gni+WfapNWgrXxkfFOcfMfwNg
i6gQCbnQxPusyf3EaxcZ4zdprtG0Q31wuQt8DxH41PHee/KkSjmlTFDV3vCyG3bU
iAzTt4O+Hyu2XaJoJ+8TJR6ofkJ/sqsTIcebHycSundcriL3/uoxIwWZA7KNXrIr
vfBUxD6IvTgY45bXlIYa3YHtTgFocrmcA+7gUNMhV3VCDCe9IyOWOyO9p0eoFnNj
Ts0JdCMUJw8FQLT2K1DuJX0rVPtZpnl+iVrBZRy7LmdjByLp/5KqdBE/IZ8mnot9
wNKdzKgQ+e6ka1T4wnMWj3S3xCx8pxgFMRl0wc6hfCbMjqmKGv0fGiLLQ343F9lA
bc1DkFbsp95YVzcZMvDHEZmqp5ilwFkiG+ml+cGC1jGWvljKeViACFbX0Iww358b
7CsQtTQkWVp4lV0Uwf+4ijYvu956Dif1s8DRJYaid8KQbY6OzqWpCf9Zqno3wlJu
7QI7384N61tLdi8W4sDzNPXkwHrIt3WOw4VZz4ylUDwmfTcm83fFm74rpAcawO0o
bWKsYItw3l4omN1HPsWwHH9GKn/9FoNuM31rTJHNMkcVOpnw2g8Yu94feydb98fc
eyBe9dK4OXGjrD8e18H3zdJBUpg0rweZY0busOmJwcJ77faGe6QKJA83Ocz4pAoU
rEQKE3oasEs/LOkL8faOIPof5PdojUGMS7XslN1EyQ0jpsh4kSHpLZwdC7axEufC
Xmpovq8vcSEHn93wmGtba+64xqtFfvRWtyLnMXxLR2DXtiD8WUDPs8DnHs9Fq/e5
8KMq/UVn50sk5jMnPsXLVY0G65TK6fV62jfz42JvtK2+MSZRM5nlTb70eNAxrrK9
1xcOCq4YSYDOqk9AsUoV/ryeEQnJ8yKelbDObgt3tl5ZJDi2IR9si6REFkkxD0Mu
V0kzfZo10QJFE7Z7VFlSxXywvMAaD0wGKcL20XEkVdNamOlKub/DqYh+syi5Y2/1
Zgnn8UmaPsUF2csey3Q6ZeA2hwN+mTeEffgqkNcEStf9G0+yxNSGESJKDew7BEUk
EPezn/i3QwTri2R+ERjSEGB5sdas8GZfqQLpnl1vs4pPGAq1bZG762vDmMSOa0y4
60/9VCtBgPfg0UbgUD38IDlb88sNI5VGFdCKQFovGNckF5ZJLzfQawERn2JJfDdD
El1tnFLIw7sLd3+/CKnNBmL0Zy2kYEwnJy+ku8TD5Y5fNPpCiMDy9CeJbnPPKNmK
P/OvKkCxz91nIws+1T6dK5NxgAijOwuHlthLEGthf4vTHgHr0eALBMi2B/Ml/H9A
Cwmm5fNktVmQL/LJUAisBzxz0yHvL/QsdmjNxg5s4dx0aAuWdpqYz8z7W7Tdu+Xt
R5+9hi3jq/UOhbRijUBr3LAlm03pkWhmSR8cucsvd4yO1t6wQQZORiWOTSj40PZb
y+NGj32yGCBjdRFkv5cidBQcIzTiVVTGRnA3/rvPQdcjKu5O++XU5q28qdxXlc0C
BmuMLw3HOgOq2G8CzCPTdR1PkAI+sFV703BMbj95Z4RsoF12B5mle2QuHm6rYEwh
0WIIt+wNbU5GLGf++8Xzb50BQIU2RHbrorBZ8p+8P2l+CY1Adia060HSzvpkfE45
xJzS9M0ZbbqyzZRo4NKJWqNomB/IaCq+uncB5EKsmHNrLgn+6SU8lVclnezVwqZz
hfZF+euvGeUHG0kzckPW054C3Vw6qrsTyQ/glas3V6M3UltQhGz/FTXkOqwWgDV+
cFuoBw16E4gGSpBAmr1byqj7LqXaXIQjigrzmizF0OQaas1pcLrK9+wBvbhT8+r8
5582EtZazUNrMIhQbyNN5R/eHeZlR2NDRelbzRH3x3WvS+lsZgl14APoqlmAwuhl
pmMroV7KW3G5141s8wtx3OoV32uZdW6s9lEFr8MJuReZlOw4nVNB6ul4rFZQoBzd
GjExodvVdfgpvxXvHifMpv6ULi8P3TAfFxK8bu1me/wuqIzcuYE/l6ZFOHL/WMOY
8ctjps+t2s5YXrjAJYw/iXSRRzB1JJWqmqU1armNos8Q60TUxsb1OUfHNQBeDfVd
plVzbbDGHnz+EiHQv6a8whiDf7NEflRhezwudGmbsnRzsuI/uwbsgGh6SpYIJOnH
xqPi3RDnTI+axMUJ1Ug+xdo4h9VC784WNov1lCbjejNhVgl3ItzzfewjJzHQvGEb
ZjF9ko1O2EI+j3KHNgq6RoJtVkx3n/sq4troaQHijPU3TaS/4BSvBmf3+OIn9BMb
zG2MtO8iOj/roCUcMGgzlKBNh4D1+ueFLiCLw2kjmLhUgCzy4Uddo1m9V90tyakx
kjSiULxBmAKBAIQQ8qm3DAqzbup4qeXGxDE2jo6ApPhf+mTnt/Dh4JbJKGnGRlPB
OhRtQYzOSt2eWgolDN3UZE/uaQ1XfImpl8vc69GQ7XyKXTJaLNmfBKdP7EucGikR
U58ALhlTw44IPS8Wp1S2XAnt2+bK0rfSGPMNx5Djrf7uFIEpV1NNiEjKNFb2Z6Gp
72tQrJ3ehbLntUnSY9epRzwVVVy9Yx8L1EyoNneIxX8XXuFP4xlPmkJBRgtWwWWT
liP2yNN8fxg/2V2HNrO5TwtWNBmQys1hcQcI+1ROxZ9SVex8ZrL4/GTpT3W1PY2d
DoIo1CeFtStO+nobmbvUUTG2yNX9FdiiEaE1l1gDUZWJXAMDylwtOewjEctwgbR5
4My/8STDm6DMb3vmHxl+0Nc8m1QEaprOXfrMqQQNLG2HVKpIzue5tOkzQitG8lPy
Q+05Wbk8qMtrqfz9StDm2s8bz1L4XePh8Pi3xYFYjdHhGIOV2YyJelOF1J0NllBP
NUsReuTdStwtQFg8nE6O4Dz3Jqpt5w4+dOMNO1ZfzrfhUKtfFHngkKk6qvbw1mPs
hnEBlnAwgBhdbSQ3AeYLzJTBYgPQzE7+EHGeY8d6S/iINwjs7pHk64n0MBwkuK7O
msBLCdCEp8pMMJOYuRzBlygoAi3eHvTL6JwYs6ac2z+Z7N/vNWXGWCfyX0q+hKRs
tKO7OF1z5L2Wljv+IS6WHQ==
`protect END_PROTECTED
