`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VH1UTuM7WFwwRsCJgdrlv/NlxdT9VxPAjW8J+wQnFj2yt68TQVvN6OHqo/0AnXV9
Nw+qIjqenm1uo8sHwnU3fiqETTPm3ckH0cAIdy+QLIoxrHsaVHpBr8/GDCz72J69
xNXurrLxucDFRUbXAKrmYzXXETGY48ghxCxWC62wlTXFDM6Pej/jK58wKZBB+uwd
ibeyOGA1REYa13FBtpjdGlzD3EISmgYGLSsnTEUH9CPVpZnxjxK8HuW++4Y6cdkm
01dSDL5wVM0Iunwn4LgYm65heUacYuw58FAsflGAyl6EKwNkA3AamrDRhdYCJ5eO
/nWnyF/nhXEc0WZSaLA8wGXzVUP3+UJDm2QOVmRO7oSyh1q9EbPB7nkCKIRLaEZY
jBFLbNvlYPoB1QzheFdLSzTfFTGWjRWR5YfIkU1yVK6EZQXU00uYReqdob7Xrxlb
mcANR1LqgEWL+WvqrEXkIE/sS1mBk8Uw+xMdKGgv0CGrjLYtrGGuy6E2FHkeqnMa
Xi6fO0dGpvq5o6W2pIxVOxefoN7RAbmYNSVM/udoGBc8p7/BMAa+3N4kjK5TkuZT
ewb+JeeOlZ0Ug2Qjr/TQKnFwpyn5EnBjNrSvr0D3tiIu2nOti3vpGOh+UIxw8AH9
7SN5FZIetEwDvtNgryqsOrRmVihSrQCcWQSdlcmXf2VTxVTqje41ilpL0Gb5HcN/
bovrdYSqAufKBtR4vrDqxMI/boeTZzqIOOqe5vmzT+7qIn/+DXgTLKqPY+4gpZJ4
iwQa7eLS0eVN+KYBpZD4+u9+m/qiSjSqWQRuvOXa5dJ7zzeRDTyVGqPYSQJLTuf7
XeVBtArU5valwNAtrf99Lvhska1O0LDeX5lbvJbW4bXI+gr3Bh5yq3N5DRdseUCh
ekWm0wgARlmwWNzQrvCC3w94hlPypRNj/yaIB2qDKrII6SkD4pVm2B77/XU1caoG
O/Oc/vtCBD2KULJgxju1p1w6VyDU6BmVSxPILEEpC48aiiw6p/qNss1qULznO3kZ
121vkFMJOPDEe4re2at+DPNFfbgTJRgXbauw0iId3nE=
`protect END_PROTECTED
