`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t0oxLwGWU2n0jbCrSiD9ULKVhYYP7AYLeVjy+dNEiUrbDg+Ey4cEFmeiGmI7LlLQ
vcZ/PhO2VRwG18wisErllCuhC91inn/34xSKftv/X+IJ3O+Wg47t3vUGEDm9CRwN
kNeUfX/mu2azPTx2m4nvhFH6Fr/VLPWPJ4U0oGBZ0zazO9VSDoFP4hZkCPKWcE1j
pgIJ1C0N3ElBLxbSFUoddXO7LXNhAgPRiKH+RcN5jbMbZovBzgXbGNOVv+PvOedY
jBbU9J0sIVohwwVR6VCPixLfsVTFkILKQnFz/LbS5OGoLAkczkQJoN81YYgPsG9z
659Fgb4MYfj1GBP3+7kIaGk31Zd5o/sBPbDoHEfF2eIl7GpHj+bG+6/gN0AQCrTI
alPnyRDJ/WTdUEBdRQPqM3W15CCZj5PG2EYei5wswmVXmASsIhNzQl4EVjjLoz73
`protect END_PROTECTED
