`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lqRxQO6d84z8e/dtI1AAmQRid++WI2/u1+CPCgujaeYvGzTuDzouq8RPLve05SAj
jxeJXowxt2keL4oRJxpK+wu5oAyVHjQ4zaU5vqP3gwKuPIUhnopuqxrPorkak44e
MgHcHWEI/tjX6n/8wgRzxxc4QJ5pRkauq5bP3sQflV+z8vA7tXDVIkjyvRakOctS
1EPQmsS5k28QdtBkHbG7zQhWr3n6YN7BF1LNPL/ZelVPzDpROIWUlnZEzWi+SS6n
YmVxT0CTeQsZW+ifNPkETXDyZe5o+WBwLrlHhVO5aTl0MLO7CTU8zG5mnqrkxiuF
xsrPNAAdVtU8t6me4qCwF0Vx9EqAbppTBeJcZEL4TQxrucxyheUgfQ2x8+o96k6M
VwEznDxCWZG6hT19g1ulhGcVKs41M+KorFaaMCjOl//Mh3KiN4xECZhTNhCeTSui
aw8WsbEZc/S49rk7lLZj/Q7W0DsQbTR6mq2IpMgU4WVTtmmq9a99qCi79fhiW5X9
yumNyr3pnApgz+QDHdaCrW1UjfZonwK0JBRTxTC3leM7tE4ZSvntib8P0bYzkuWB
Yv+/eK3rfx+GTsk/vd51DecuzIAXNuwZS3AZ/3Mcomxf1WqLwdyETW6igXvngGNg
tGg7kUAuUBG6v1tFP3yILw==
`protect END_PROTECTED
