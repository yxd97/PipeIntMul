`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6k2hkHHSJVuf3uRU5gL+yIMDL0DjN+txlOZNAerxBXut2f5a6oMMTnJmz6UHz7z
ESZwoabhQb86xXY7rJDJ+IzNzWq8PZ9KMptHaw1kPovktowOQf+cLMLyk8cvGjhw
a2LG2yAx/ZFpJr0k49KtFahbllrNI6j2doPRXG6xyzkN81Ef/JW/lWJ0ueF1oxvL
VB2UnNdToHNEsadSmaC/Fbccv7tCC1h95sAUAQJuakCcK4OOPlD2YIiWCxT9VxS0
BO6esssUDD9c1Vis90aWZD8epXpfAPzgt+ruuJIZbuBWCeXaew50kwEOxL1OKRrC
n3kf4qhqgnKYcyJrgTKgTBGh77OOu2KFFYMt8k8btk5qiC6I4fJBU7Ns8fSC5WP4
stgFL2yESjfYIdWLuycevCa1j7YBhmZ3ht/6HfMSQwr57HvzdnJzGRWaBM4+sAPc
g+Jpn7eW6YEBceQM2nfuAQ==
`protect END_PROTECTED
