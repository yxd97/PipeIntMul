`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hadSsmHdvTdEtf3RdN3yzij7QlFW/GzmDlkt/AQBI6He/+SpC9J/colLdOqWFVhx
OXjFnT2hWZUejLCMMk0VzdxHY5WEtdL0ni37u3l+9ZdeEq6GopSmde9vo9qZ4kHv
NuVtN9nHDdjq4PyQ6KMjVuUSMwqKhalo8GckRtgAKlLjAin0G589uRbPSqcB09iu
AsEevahz2ymg2NPYTLJ3KMbUo47wFrJE06L2x7gfj6nsM+LzlAQq/tehs8izqD/o
RD6Pfmm4zDqf73pFPM7n+Iw5fDKqhLxbJ3Gly4E76UHkqHK3a0Zaexn80DZDzzLY
NKmDkFaf1s39WMDUHuN8zlbLDfxfHebdrZlDcZ9tyKpd+PpRo38IgoTmCUJlHJlh
o2L5YuC0Gum2KZmUpcAXIrttwli5Ng1NMyOHCgX15G1eFSPjbdVQ0yGeoaTjexar
OShgOfcSYub0N/dZd+tkOfONRzvjDwghud1gQDx+oTmvi9dFtukSEt3YHJ+RZq8j
rHhmsCexITZA/sBRwm94XnMIPoz0JPCtit34F5J/Yflh6ZQOUa1WKpnMInFoBNIQ
X0T993KnDBCYu/U5GtL6pSx0NFAaX2IRd8Gsy2a4q4E/SwQm374rBTaF2XFaJnfo
cK8qR/ynt5Kg6CUh+wVm6my6tyBZC0BNpNiDRtJgxx7c9cxWYsaMfqK56LlvpkQX
c63g+0ryTgW0zy27R8GkLynA5VgfU0o5NlFh/YdmPeIl21sStRjxIFyXtGHcj9NP
Xpmg+fulHlEdYY97SrCkyp1orFbpNfe9kT26+TOzz/RqBPtmRHNAKwZaRmV+eXSl
XHnUhc4odz1ztg3Xc9IiJ9dOYL25+GE07oeYQgxq90rgGXFqNrpQsAHAuH9wbNrn
J77Y4PIBDbPblkaD+EqCCSliIRGthA9mnNWgGi9HpHum64RGccWuw4f5IWnczSq6
dgeE52+Csl/CMfB7Oblns2A3QSZHalbsIxmoJEyr7oKBRzN68SMNRf52EE8nWxt5
5nkAFvsfAe4ulB3c5zdHZim2xEqwUFo7Kb7wu6Y8NHIyclxfNMRAsm/FUogDYjhd
ikXfc9u42r7l07bhpq7nOBprrySLxaAroeAmcwt2Evp63F+zpRfrJdSofz7NIzky
7SMMfP2EAJ5d3lhR/WPdTNLPRHvgp3g9euGvPDPg9de1pSHREgqyzFyb8nXeu6Au
yI0bQNAHnfEBfL6ehOyi3KdsfIUlR8GmclJGFKY6NSRJYU+58IcV+FFEZUUDsZqx
anPmchU3BSlh5x/vL2cc0m3Rl1SrHmQixygaCNnvZRuC8XnFM3AFjhjqBtEQgQfQ
DUKUVtJzoxwluUjp9yEV5FUbycMKFS2fIvE8LQIPDdPB+3sZW5qZSrAOKTXRv7WF
uJv4+wmhLh8YjMbl7HZUuFLrqIGe4U03Onbg+YdIs2Cy6ngcl0VrzlzxC5kwx8KB
01WyIGjShgF17qEZVVgw3+gnx/ofytcma20RZS7OfX/zBW56cMliAqrVGTLKOTqU
aqCFyXEpXzLB3xCPUR2M5v2qEAUFZYpfJsIw7FtAZtH1LNeTxEcl1q5wcnHTPDVt
SVG+4RSzVdTaj00q3fsxz4S0hILwlqYElWDEQsJIPSyqamJ7ZUM03/x4wdYoLIjZ
zqt35yYaTKfVyuezLxi2DY20sz+/eq1i3LDgvcpU4tQjBigf88G+FwyaFtD6BJEd
CYZqMHL0ys0wLB4lpde1sIPoQpgcewEIn1TGxFJOK6E=
`protect END_PROTECTED
