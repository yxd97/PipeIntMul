`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x3mVT9rV2Zud53COTYvnKlvGDZocRHkTAmlULDvznHSDu7R1+XFHbFvmyVMOBLJP
vkVVKAYvQsgPeYB03WFFfZUUeJzXD+YbyHGPScPSP6qLeUqMCcp1EzwfKkkPaIZH
4gYhZaz8rIReDZZiv0Z3W6jvGSjg5KnsskFGDUOfcD8Inttim0PmtJTPqSPnWeZd
2Kw0Nf6jTd+BiHLAFw14iC+uR4JjHPc6NKUMo7VJ53qSSCcS6g3BvvqQ07PCpnwX
K2k6fGmDGxinW+JeDvjVSQ0wxg5ApQZxuurEsmpYtSBT5373IENsfGFjFaMU9NVL
xW56wfSzN7Y/uZdr/6WasV3B9ESVm9KF2FJe5ejvcLhlfn/ctMRPkHw8mebKOLGs
8tEUJQQ5znY/0BmoIP4DBDJXUQZ8t12Iu5vsKssK/suldKWaZb8UxVlhjrMBPyH8
Vaa+pJkTTEvaZH+9/fPRqkcFIVRU7kT9VZ7RFmjRPDdsPxhJHgaBRmxhgyiz+Zfs
3uLhIeP3GRGvERzXpcKixnF1WhTjHdhfl0hK4Ds7kIZUApSpj36wiuRXKj8SjdnM
x06Ko9CQUP9SBg+JhpxSCvEgMyjIwuZe0klHl1RtVLlxZYlnq7G0QNPvwxegL+5M
oE+vcJRzjwMaThGzfW2wp3c2K6Z8Tx/Lp1x6zRtc/d5fBqiFTIrzV/89NAtkWjP2
kCq1tO0B2o2M0PTXKb0r7mKFyAUb1FVvT3RMWZOm5Z7H9tPDtMU40oTQQRpVaFwO
7c9uN0eFe8HZGfIzMWmgQpfzV7ofR1BitFlAqe+fDoFDxd4iaJMQEv0GPabCz5Y2
aMl+El5igegokXCoCvMQM2/bf9clbQBS2TZ4d7FuL7M0N9Ylmd+YbCYMiDobvjCs
H4adDiua2/n3+Y4Ez1P37IYmCaYMv4KcxXu42IIzEfRIFEdxxDXrIryUiXrHahIE
n38ALRB2K9aAeu27qVEYUofk9S4GjXbi6xigu/M0TQEWv44uW94s+5PUGvdO8DlL
jbz+Fsb1NIsIJVHL2hMcKbJkwPNRO0nEpO/p8YMvF0Pv0B8zUZ5iZG7UbxxEVnvU
9nBR6NovkayJzgBztWjuejALYX2BAhTj4shoLYc/htH9oozEqKBOpdKS7Q+JUoA7
gdVaJuwbz8UyjpG3qpCcrGmd5BDWqEuvllpBF/+EdObzJcLmXXjvWyOfKmADlJaJ
56UT3d5AHZ6C8M/2XNJAmi+0zC/u6O8IdX584sg07ZZR8yxEtnxN2ye2hhLWc4Tb
O9F4Yi3ACHzZLqJHKdUMQx5NhWuqOWMkSFKAf2zNnflDJEXOdKIOtF1ASJRc3oOu
91RMvlyvQrLbr8pH9rnnII0cYAHk1TusMwcu+oLClbAH2zCwekkBoTN3RU4fGT2m
b07gen4gwMIFgXOYE22H2XTa+4he90MWUza+AIEscbGV97t4ISk1ajvIANnkwzBl
RyrAWGRSKj+rOnN+374CujMFLAyuBNt4iQxN55idy1c41QC9zUbztes3GLUEXMiH
Ie3CpAe+6FDzNMo7Azi+btM/VjrjScahu+gtWLxOGHO21xtS9e4iYjrkeKXlhtYV
lQWkqCZ/1BeqqjAthRZAs80v+wfEmm9BzV4HmperAHVStoANm1HFMdhksn2bfhVf
RW2YUHdFawirya/mzABtWuItp3rgSjeZcCTY+v4dbcxIneURp+DzIbdPEUtCxdkN
dfhqQzbV3VaDphgRriQC1xXoIvRXqBapRQatdfR0OYwfi8YlYQYaWPpZUfrW1Urg
dSVnBJHzwI/MWMX6PsYm72/GgU9M6t9PxQWECqSdwA1a69RDYEkd9TzGf7HDHSRe
U3/p0dDakTdIp4NeRWyKR0AAKcDazqS9lxoAbZ1ZlbclvThUyIEDjqh7JDk/hwH/
cf5ArGXBjNQ1jVGJv8MyLTqG7BNZSYlPB+S5rXhUl2Y2pgQ+KQSDLKAnxcqCssjd
qZzX7ad8yM/EVIeiLF0/6rHnT8feBaGFWi+T3qgB3qM0nQ2ULF7YIc7SmSBwbPG9
jZkULOjK2cIIlytLlD7DUEybziubdmAuLZEsLy+hrJA=
`protect END_PROTECTED
