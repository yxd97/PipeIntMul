`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6eckATvKX18g6V7hzBZXu+QdyAW24MqcVViGiWq0z28+pXn8CHTnNyNcAcLu/vG
s+shRFf5j6EYzzQxihna2OJtX2cP8TIo3pokAfW54DQfjdC2AXDjsdUuGh0WjNjs
nUOMKP6hSkzyGVD1HtXDnifhtpzoCRYV/rViGjiPveHH2aHpluVckQ8olRts4w4i
/ygUkQ3ecVBGZAH/7MkkGFfPvinj6KSQQrfPcQpV5xSdqGOIEbKEec/bEkjRPiVR
KTsINXkgWbL2ckKtb2HWhFin768jJQvo5mm37QswSLM8EPvZd67H2FINb64XtZ7Q
lec7XPuu5SUbKkw9vjCT4DmljCo334myc8HY39sY+zu8rlYJrD7neDbLcvWaZNfB
HIM1RsYFiPIGqW/NKFnJg761t/Or0J8WsbTVjxoCzMuyZnnvphYzGuLe2QsV0JBc
3DIFtGhY3KBuVNr84/QvIEyK2E4FIXs0GvWDQYZMJdt57917cgXbvD/XGNNeJMv9
yrLNswiu6ny8G6BXvjGRWsMrIkPx4mRRYwIF8S2yvTM1+OefXEVzqpOCMxDV7fX8
XFd5M97YpQhrXJg2vjjkQtd92AeGGcKYwPj7xZWkLdmR3+WS1tUQh/1RnHWy/ece
5h5cF2C9vvsG/QIYt1vbE7ErYjs+zUDIrDmAJ9JLfcQF7Iyji5IYNIMHTHJUg2UT
pJA73D8XR4zJoNF+t2VW39RZVaP7XzWJ726jnmrwlATLi4JmKecRosrrIQEQZKiQ
pe4FfLajU+hmid6rb9XPTwWQR5yzdI1D4+zFx271p83wFL6NYpumg0zJqBW2VVdY
0wjtWFVrfoiVuM7nKwel2sy5sLdhWAiSyl8O8mVAqiVfLSNmoRnLqbZlzzEb1YKW
KLH1+rtMK3qSoz621MCS90168jcI968sqGI13QaRSuOchHNuM9XsHlV1q1MIACRG
449ka90L/pMS3Rj6vI3rj13pu6ZIlH4W5Y+YDFg941q/7BUvvfS2TepyHHfLcQHj
6O28GkSbmLJOGWTDa4bRx0Gfx4UAEMRFhk9ieOUqYT9eNvBKTuJpn8ygfgz8Vv5Z
x4nyOOQfDauKHbOAB8n9JgfvU5zu8pXfmEqYlV8S43BxVVIGU48iFVLSJ0UYSBun
G7KI+LX6YIsqMouPbWYOelkKMjlefPwIuHSeH25vX/mfwmMGVJYvITnT49e/RmbQ
nbBpnyX8brUhc2RkGIWcwBJB7+lJIwgzFXQeBXgaD8Bmprvmv41ZOrJeiG1VosRp
xAYKDAKHZrht2bCNH5mlmWvN2QGPT4hxYXaiYanOgNGU2qi3xDLllll+saWx+vRG
lznKIx4JqwvQ8Dc9/nv3OLx46N0jZEdfQpms4zG9ZynIC+KOWGpfJVxE26B07/BF
VJYkkWC/C4I+donNuYMwj6h3sS4Ri/Gh5LeGkML4QWFJHjmCqnAA800u/3D029lI
cDPIvYU19nIXbbTIA1cOEg+pchAY0THQ9yt1+vtv1WrKJa0ivj1BvRroH6K2kdrc
LV1TTEHOkNv7EUYFUD9WOk2nu0RAokv35u3hhlYf2MKL7wl91HqEa9WDVpeE3v0n
RTLk6qCZZLinAfrju3xHttZG3mQ9O4WhN5wHK0qVPXGhb0k1P7Lw6nSITEzDBxXQ
OCRCPcTbN6uo1tNSKAwOfrmAKotrkKZ0jC3FDH8mNvaSt9ki+PYWZp+3TXU02OTc
dqoOYu7vJSbwsNZvJpJXmOdfL++emsCZrlA9sZZO5mfK1qIY+Hq5GaKOdQKblHbZ
B1i0fZP1LNEKZODlP89JdYkCepun1w76u7OIbEzSW+EJy13Ex3gZpWXnUi4VJzOU
4OVi0maIFc+ehILxp0AWESc6BPfCHHJH3B3cMhtFRr090XTAiKa/D4VkEYBYoyXv
qejtM6IokCLqX40l0x4iBVyBgwjLqLHSkGt2qlEHToF+9OZgLOajr26tFFGKgXeB
EtSe3jDkCBjFVhOm3tDGajJBcyRawXT5uIjK6Mz/s2ucnhcoNzqu7y2AwzfmTXVZ
CM6RpnFDLa38PSsRve51Ss3sKmlb+eA4ze7Fqd7pJc+mF7q1Sl55Qro/ZasS5NVU
`protect END_PROTECTED
