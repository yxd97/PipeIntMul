`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxIR/lQqm9MO0g2lZT0Fq94MAUc91+62nQIdLaBlwpfWyQbJK08MH4LdfF9HH3OR
PSg5pwvLJwWJpLrdhdlvlsipqdMmR5PvyLRjNxf1yzL2rqj+JCnOgs/WxjK1ZJL8
tyOIs3AAjdEiMt4Mg0eCnjFuwwX3Lu4yMFxhlgm5nOyL3CRczkO9rzgby1mhdZAE
2ic/K1BQvXZE9rC+GYGkyxGyqu8D0+zri8OdqoD6Kcf1Domo8GuORX3Cgp4i6igD
dT5P6eeeBi5osfhTt0b+QrkjDaq7zLpNVK25D3rnCFpZx/N+L3bmK+zJ0mm9v7r5
HX1tB7JK14llwRb/qDMTw/KRPAWb13D+2nO+/nVfMdp4o98up7tWBHAKrN7d8pKK
GUYyfh9W781HL7qfGRK01kGsIcLU7aLA8J+p8WFQ3/ZHtXqdX5WeojEOm8eEBNqI
YQJkOUPHqG9leDGS6zyd8A==
`protect END_PROTECTED
