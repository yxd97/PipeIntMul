`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y8XGOfrpH70Rxti3RQ5jypqNJBqLd/b2oaMtPC/pz2Omq1LVcw3F3/RMggUTRV76
1zHFxWfl7p5FgyZrR98jywrUG/J9d8nLwooQYKVpsbU2sUiizzP1QltjJ9hjl15f
++2GGsDIAKpVwQhqZZFakr0XCYjiuZbRGLPjDCFoaBOtG9GQ+8AWNT25ZoQ/13As
r5Ilw2pu4CqNa3yLMnW4MrTbfdv+Rmb/LiZhYGXesRXlYUZ/qYLo7AYhbHdxLkiT
zvyUYZE0LK1r/lkBzLF1zU4zqs6OIuYvVM4frJuM5zMPVDt6ZtFLcOQkpvQ//U9j
BIXr0MFScPNPHdTrop3as9L5Qzz1bbgE+Kzxwy41K9IGpg48KOUfBD6kdN4BQsRb
ngaHgdqOrIeE4qjEvi2hVpspgA0xCXCPUNEECioqSftBdsZdlgWHohTAqxeAa4EE
p8DQRGDyw8h/PxiNV7G11w==
`protect END_PROTECTED
