`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EtnkxdPpdBC1U163lOe6kipLN7sLDrgIvCTCuuLoZRscUl6kvzq3wbmq0MKo4egJ
B1WEvfG4hQ6q23Wp57d/s871McrkPvvqh8FUUvtlnLZ2xm3CCtYLBg16bhZhKy/G
RaFBUMUyb3iYVStKjAaKmhOzmlEz5q9P7ucjfG7PO+OJB0y1f7KaLtfEZxOiIgc9
AyjJyffUqCev1KYcyzoZUHU/w0zpPYHgg9Ahv9U/rhlJ/RCm926MC8iFraG6mi5T
EfyFAyMV0VKr3vGkdwCTpBgPBdQ/9lLaqGkfTjEd3XQUyPZ/KDYGJUSWPqa8P8VS
i39akV+8fDNbFblFbcLcXTcX/y4IIpWL4iP6zR+5kFNubZii4TubdGuzXYGeGuds
oKzlyn/l718WgYTI0rDymubhrXQo8E+DPBoG6h6NRwrnsC1ncnfCfWgCs0pAfMez
d0QrFg8nCPUQ01SCfz4oT/Lx4ZzN+4c7kcE9JdY/dYIXPCCJWKfcEDHIHceh9jhy
iUYr8qetV62TQuX7jahFqAsQA7YX7jYOIkMsBvADxG7SYHUWPmV+LweOZbcThku1
eqSIM/Zb1ibUcLX47mqBzigQPXZHy9F/o2CuYFKPfLXRe3sXTQoBHSJ0Tq7H4nVv
2G6xznGB2Taq6KYKaH4UjWTVGF/cTK2VQmkJ/5Wj3dI9GdbTQAi4xPeClYHKDRAu
wv+NKyWe0i6mIaOIjiwmDwT2lFzwu/blUABkI8faS+ogK1ZlN26TFu5cuSWbNQ7x
iGZ0jy8+APgvGw4n3YKRTSx8aFc7+3mO1fu2GbEnwq/ssYSWgASkL3qlDsOPZ8bV
HjCOZSloNPXo4S/V552kZZI4SriD/q9doB3LO9znR/M=
`protect END_PROTECTED
