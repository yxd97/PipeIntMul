`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X9PIk6vLkBhAqp28vtNs5TyU+d9pvYy946+ovV6c5PkyuTiOvoj0RCDudLk4GP5k
v3aJMi5rNCIf07jmrleEIrXaSKmwR7TNDj9OZakqbflSY7jjc6PU7wPISx8dHQAA
F7QY5QIXH/5FRiePUF569z4iOcmhk6+BhuKPtL4xlWc4T77H7Hvs7uFoKLmhfBZh
lOiTvNaN/PX97/rUOfr7Pp0aky1ok8zfPfvqd4HLvedFnuoNvIL9VWYEVbGh5PzT
QIWpcldjSk6R6/6hu/aSsgtDN80hi5Vu0gjTrwWC5AK84bmpaciVtmBDi5ONFusB
oWnA7iNGhp1fVfKke3cUhHo0GAoYFjGLT3Gew34TEv7uZgBtMGnFAqICUIeDVfqj
UkeOk+b3l6i+r1jpimaQzEAzyI6/egff9G/CbpoRHt374EOvYX35eDGs3Gw3x61o
R3lRqOlJaJqRhh7INd3sHmWndFXsEKlZc0DSPcfjlqtKOrRy7Steq7RambgMDSmG
`protect END_PROTECTED
