`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7uRE5kUzVPjxuk6zuBhQbeuov2/yFJuVsFJ0tF4mTclAjvFpSNqYegYi32jpbqh
l9O8XPpdwh/ggFwSmt9axVuambrBPSQWgCZuDjh62se44R3vxvHWG5rWI+P270xK
4MhPrMhe1acxyI/mM4z6JbuEtNtycS6P8O6t+pwOY63Xiho85BHxiMyiTYjI+Y9D
ilk53Wf1uNaxgOQ3XEdfH66CYnNrGnBk0XS2X8y4Qa8QI0oZMYa1t5nxI/uF2Yn9
jhrGyvgbEKKvfgFUpVScbjnzKNOQCY4jeKmRA+ePNXDKXry7zAJYDE+ZNFsw0bKs
UiMT0KBNrCmwXvgyIssAz1lPd38btYV9eGO86nDB0In9KSwcUSXTj3z4aTDVd+vr
FbGHi4dsczuZur8gWcOV5UoCYkeIyGX1xb/orBmddfyPCZaJCpT83y2PFp5YFn0R
i/otNK/jkNjYS+dtdH0Qbho1Qzd5Q1nItqw2qe/UJHnB1RoNd9g+8NkNLKtTiQOl
5ZVAGXAV5QcF76+TCOYiy4VZs8lkif4RHiPB2CXtilHLAUPlesSKrrA+wSGHRQ71
uwjte2w/+38EzLBj4Hj/qYgFRlvYwzx1fIWxNxeq+Vz6qO6iDoqgG7krIDDoYkTE
wTHfjnRiRdmoSEcPZgcUOQ==
`protect END_PROTECTED
