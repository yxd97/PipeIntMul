`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pTzxMHUegKEQJxc1urUa7UQeb/O/jGBITf7ZIMktihhzu268g7gJH+SG+v/RipXu
H1jAUypg60VWZ3JimE2FImm+XzcPne/zoFGqxgoQF+pMhPIU5044Xuelz599DAL5
rOdtlrQhiO6LMakIsrZZcGUume5xV4w+B/kidNFcdMBJpctu9FbKIo097n3Emaem
FcbXbcNEg6svfYjwYpFzrrof2ZmUi/kUtYCtFGJAVliSHRwcunSc5yPEEmE4oL8u
a6pACXodcAFvvp5P0lCIjQZkp9qVXLc40JP/OyVhX8C297qtn5x27QG3OG1RlJ84
26DEOiKb0E7EExQdiDNmd0vwKCaGKJK9SXrWNHazLfrl+OJ8ge1Si3xaQHumGbGn
YKpRmVpn5frsu7cT65/zSNLU2tu3IbMLmmPlKVVMViBRIPFcgZ3OVJuEEoPaNpwZ
`protect END_PROTECTED
