`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n9u7j57Ov2Gn+9sH3+IFZtWkKAmxBT1cLtifGfQkiI/otz218GbZAqB8dBsgoy6N
9wCeH9fyFBecse4dh26rXVi9f26kHGUBXTp32DMv0ETrEs5NS0RTzv1z3fLdR42g
666827RJoRMnhJ/505/tFuhnBYwUJFrsqwTUh/bzwt2XdcYVqfgzo6fSN6oq+g4i
HlCRFbTtQW5y7juWlfU/S5gU7mXP28EtYTTqwSNebKktdV+618oL7yBcwZ46IbKJ
+ATY9MmVnHHVTtC6T7+yOspMO1zr9krZK0SLpI05QShOJoCb8Rl9uFlRB6cpQTjE
Wf1HSBwm5HuSMjiDDV3rI4NQgW/sGNIYebxTxsxwr5ww6vwpYEyq0P1QttH623n2
`protect END_PROTECTED
