`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBO1aSIPKoefda/+7YtDRxpVCJoj/CUPyfcp50cYFKvFS7D/wxu0AMcs/Usi8VOK
Tla1iOZs2QbtON6Tx7l2z6LlUMHZvA56kpeFYch6HksmQu+1ZvQ5JdFGk4mE+aa7
LPeHnnWnH2flWRco/YedaHbvJFenvNk1l+Z6lNQl9eEyc19rzlHOmqTnsGd5mDRJ
SZ51uN0CMfDtZ5fd6ByMMZIeHUG6DexSJcn6Q6nsh6nTtljnhpR9fCDV+8QxNG3A
jEFxvMc6fczvRhXlXDeuDOCeM62ik9MGgFdqCS86w8cxmvGz7CyrfWd/FEJmlhRV
ifVr1B+Ccn6+AG9+Wxzm23j5VY33GcH82/59Zc3IPNUueiZ7j3wAXOEeg9HTvsx/
YDT0epZ8MVPiW5Pqv/sBh1ZmmrGJUcAs5+2BUw/87GbsUAYrtvKhU7TQUalnnCNN
HKtCMMTl0lrxptZ4ztZRWHQQ14CmD/dDlOpSlsOVQx6DeIL3V4kQJLXOwcbY1hzI
WxVDqRg/mLJnZKKE1WkfEMltAQoLXXPe6XVGJIE9p/NTXoNm1+H99uRgyDRklZKQ
7k9Gi5Gs7O31BjnyKel0UBZYIYGSFVMglEiyUnLNWz+qPWDDwB4lWX4H2wyIzLyp
`protect END_PROTECTED
