`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjX4tSOKOKtCaL8RBgjXQF3CiVfVL5XzTt2ZKBFvezv35vlU25RQcuEQvMBkJQSQ
D1yeWtGbtW/Xk0SDce9b5x4jdn4J3M+TUVhhMeJObzmj3Qir1HvdS6XMHKLusFPe
D+mta0/pq185CuwZOq3+TYGITWwXkM3zsaATu5ZDLlol36rE78CzvJ/LqCbHrLSc
hhBsgPuD2jQHs5XFPmJ9Yn9ZSWSMoDc5BsRLRBazNsxttL7b4leRvFsszeC8//08
`protect END_PROTECTED
