`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
crz6UUumxyHesjKOxU3vLcuZXw36lnio1NeS48tZYc4XvwO6v9KwAF9CbDJjl+n4
JFUtZ/UsYoQZ1qnN4I+2ob87zbvZWQBYzUcY9aib/aFmjoPpW/ETWeGXYH9ARI0H
3vGq9e+W0W+Haw9D/bu6lzNqbc+tiQ/4QqT3euxhGB+/G+7nooKc5U2uR3ETDrrG
/4qcLdv7xBDqonhy6clxPBOiLKPDQru9ag0qBqRNujkPEPQDkBzJpVYqSL6Pt+bS
M1UHOSt1e63oMiBREt9mTR6NPE5pnthfbBhugvTJra2ZFUZK6sGTxdK0oVzvEEX5
VuMbHkGt2cLmdEXYeRtZ77gO/phzQTj949TiDBQIkSx60m6GeFXz9rIWiHmRuNoW
+E+UdA3enOkkkaWEJDEQ01fiTy7je76dKVJhDFHpYX437+NiHAxqP2IOYFgEnAc9
Ajcns2tyAY2mJMR+BlsH+SfxG0ilYAsJzNRg4s3h97TORJImybIHg7z98Fr6yqlB
g/0rdsBH+aoKq+wF5iYtdaXclX0ZJOk46OhWgRs/SQkHuzTGAThhCxxVl529xVJk
mJ23NsisRlOuYg3sFqXC2mboO7WVqCuCyfhdlTc4e3eNc6J+23v0SRXc9moIybJ8
Q3cIsuLpQ3P0pVVSI+v/BJ+8n93t4mfROnerTwJfClYs7Fzq25FuzKYtCetM2yhH
mAwnxpQZrLWxc7R8nhm9jMyUoEzZlJ9Q6Ubx0WBAA5v0LTxLNvKArzgJ5VHy4YpP
dC0cc+TxDep8H053ulF9Cxj4vtYhAKLhog7lJuXdcaNwkQypl8EWTMZlBAVaKbOm
q3/PGUrVOk7G/VOVeICmjybvixgWyxvovWaU5wQ9N6NDNKaGZNep4XT2MweTWqyY
VxSkve7qi+cERiG8EnMiAqg9Y50dE9krv0RGiMPyeRq6e0e8cpomVhTvIjgnaTdI
5Cd9KsNjJMHrggq5kEbhU3ldrki25RVi342tS1VuR2+IjvKraOg8UqC95ujtVcwT
VUcEuM2t1AVEDzYSLQLuGtephH8ZbFZ+v7Dl/PVIG910ftK1FCv5y593lgev23m/
SPEQ6NiNPGZQpiKv95tnceVkbVdXQuuyK1envC8AxdCZMh3xl/Hwueeo2NCvFlbZ
xMvcZSsUbe5n0qbgSZ0iY7tESuSNt0mJduv8WGJbWL0TUKH4XjQV6A1cNKUp6KGK
oHAR0glORj0MDeOLa35SP1hmGcpwtryAAMbuFNPnXIWzHvNywSN9ug+nDA3trlo/
76Yhdjk6JOncdfqsYhjY987quN7VLeAAcONJmDUtpA/cR5m+WmKF0/bJRt1rVlmH
Wi/7MwniAryNQzoNIfZq5HTif+aXLXce+6EOfTCFJ2VVevb0RM+mLAuKxu5r57dr
RCcfagbxy6N7yXODcy/m8BqKtsvEvVXVx1EWbTuA1U1MPbtmORs+/2TAt8xMu5Fz
NucDQLxMlYhr82prMCxj+XMx6Z9U5e141lDwDcFHFYKDR7zrL3VexkVtdBfjyDOt
AUvGetRPCBAX+knVBznX7zYWiMkYyZz1k5POlNtwwtTA1mQJ5GNyj326Vq2LNblc
yHTuWX9pHgoY8E3TMc68vkTro1VXYLIOCzYYtQafgyC04H+zpjOIh9S5IeC463gJ
wHqeEAJtySLFixs7n3qak27N+noDeoWJazdLdb8E5TUjqfcyu/edoDdFx5LLZG8c
n59u3XdU6g6YTbGalev/mrMXYgcntOSlldJxSbAQS/EXM8iKKXjIQsR7SBivPZmR
MuhG1wwu6M8AaXhs7EJGKOhueoLWvMu3HQJD2h+wb1srJdUVFdtX3AX9m9XqCbJA
S77AgolJvgHhxLGXgLp3zo3uYTDKAysNez5ND9jf4AxxA8Ur/YXlt1KuBOFfrbcj
JAkA2O0K9A9jfvMRgBIZmLI8qeJVMPNKZf1AlMSGKiarHK7m02w9DwF0E58TS+4I
xnS1An8hMOwqAMIO/WSwE8ITDOas5DZgQgUsuCWEZ29lDD7+S8e2TkdQwPs9efK2
44BRLkEZG6/QwG7gG6X9fbhXI8Gv7W56U9z4L07tP23Y6rEmC69aLUzU80ULBbl9
O2o9fwhzAgudRvwnLb6dIq4LS6kPEXwsreYZddD4e5FX4iF/21h3Y5X8/ncxU2ab
jPShaHSYGslwI2xctxzXDOpeXUvmqU9FeCRgtV88x5IJJQ4G6acMdJyfCwmzpMCs
TvZ1aU8PNiNkYjsSeE/zz3zv6UZy5XNpljY0P+muFp6Q4uxvTDcQnjvcxUktOjDc
kDxENECB/vfgqMfHdqeUWNk4KFUiBFRUDixsM6VWaG1eAs/wQjEwlSQFAik8oFrW
5OPSCdBQ+K6pwm6ALJyvP/2QtKBF/HSG7EtfByrLEKErehUqGQXWDWtM+Uwsgvbc
svNrFa20i8ai4AfPpBVdLtOtHC0S/q0e1Ekhw5ZYimzzUPJDdV9XhRhltFMLRZSW
4hdnWWVFvfaK/F5ri7XZ0L3i1qDnwWG3DSrzNc6VspRgjiaX7l9BqJ2LnXrMhgpI
aNpEP6vAUEOr0/1agGbPxFmwEYh0Uv/AAfMw/0Rg7jNorPzZabSY7FLRDT7OmLc/
xcIf68PXZtIa3Wx/g+EKOC40Yr8lLsW8DZU58/k4r+W3fgYDc1iUjxJOZZJeJjWo
dB0qx1dG0Dgk5gMFFPYGnwIlPvJlLDhOb/9hJXmY3AZEryNIAbZUdbTZP/LYjxmj
xSyp/zfHmjzYXHLvf8w9EQe8qlmtgi2nEMdktdIDjO7xKsyCiSk7W78Ju0/VgfcE
XzbM/vBeMenq5X2e11/DDOYZePBCt0y2RDQnC/pcuMtVZF0djOWH8gVyrBXMvEiE
sMDlvfxsTSaLO0QVliIEpPNzyuQz2F+GCtAV1rDQkHHrxCdRqI/BgGFECPS+fqi7
bTQlTJceLxPWq85f+vbsnR4ts7Bk0JEhEwPGy904/RpYSqqMPkENSNGupj6Y0DiK
xo9JgV163I4CySURa3Zyi8A9DOd6rTcrIhvVFlMp1mbremY7Not7o6UT/zRrsdaQ
/1Zxt3XuAPpahYk+19JLklzvLSj77ELiJM9ZykKMaspIjzyH+iehnXJmiDocgVgF
uGJ1IrBwNX5OHIsC8dspRk64fejwLSiQ3nmcmKQ7jY75PCEx72m/w8tgT7+GK9Ni
I1MYnw0xdi9uN8K1TMn7I6SLifkQCjKtjeIC1is7W7Qr007H5uxalJNhTjqHHm4s
rfonREUWKVEI7MDKv8ZmhfqGNpgkSwun4q8fDYdiVTdAhrxdn6p8uURd8lMPkxnj
yYpXuS4WosDUzFcu3aJeKBdKXLCbuWeLH+oLp5FXiGh1WX3SAGSdQrppvHdllTY5
bQeBKIGcBKoOq9fWTeSFrQ==
`protect END_PROTECTED
