`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6EOLE2SExaAJj627CpnFS1N76tz2Y74u3LUf/qz550DE/vnHWmJS5V87dBxngxYb
NLs/T48v4Ym+0/9Vl4mRX9SFFCPrUhkPd/iEgdLj7QJk0TdWYHxTa4eVDOwS70E2
zDtqetCdzgy5gvW0DiFpy97rho6io7ndlHA7a3O0QVYYFtznN6pQg5azLKKBwP+Q
NnG2OD6VB5yZSl5XGbqb/daHRWXX6Jgi0yr7676EUy49azugDC2d4cvzBhDE8M64
d4t/QP3YgdwT7adbKIv9Cgi6MozEiVCoraoNPk4ECkrxjR2O/XOUl+BdwoVgcFgW
jsh7C0E6JXoNFr6w1BdHiRDT+YGp0D/jEG2grx6Y+eBHUQ6RIdAyf7HpgjjP4qwi
2aSa52QoryS8CbwuWdJLX9GobUCyLVh6NezhxszkfFXUAyicuSha6559X39jBQ1+
7nquod5LGj3bsJJzRHJUqh6rEAsrJ2vyDfW+OpEEscU9a5D6+FbE7TMZmm7FmIqQ
VJnggqUndjBUCZHq5Dk76gqa4PGc/tRoqwVhBlqcEPjoFHpR55VRMQoOC9J1hBD+
a/sbZ75eCWlyAdth1TH7p4aK0B9GS1Psib+Der7JJhUCz87cQqsP3/vABBuGDQ01
My2Nh4kjU6vdrvdG2JvY6xLxz8Bg6kSt3ze9JCdj6f27wu7hgnAiNbytLbJcqRqV
NmDa9DPBLwRJqH/A+p1mdJONQOxXOUS/YlB9nkvDfqtE+3d+u/gNC9weqPrugNn9
0bxhFjKcU5w7scEo9TLhEJFa973QN3ZzDgXRq4oZ21PxCOh6mrXjjCwcYnBXmmYQ
T/1nWtNeAtF0f2G7Xfrb1ubtXJ8PiNs+MryUDexSDoQVrkcm5vz87/RY8bpvMdLF
4UmZsxmn5ppOzFtjqMhTRGYcooiMtTULqvmUX0KOjTgrlip59ROMoS1IpfcdCc6B
CScMnnMOQyoT88cDSeu7yE9pdi3WotH8UXZ0ediQMDIvhJWWgok6mYjdSVAMrofo
riliNBy4XL+4oWUZJ4kkT7CdF2PFI/G7/Kqy8SoZXLtYNQUYFtQwVCX4wvwfoAY9
cabs8HP6GQe764aY8DtbWRrXxfnYY2T2mYrEb+Jy9vJ9bZDQ65pUVxH9QF3QCvRQ
XLELOh4hF3/Elsv8seBcNkQGaFIsIlkwlM5IMIr74rzKkX3GrpAEObQC0Cm1e10y
9+G+/Ech4IBYt1XW6ceT9kz7JqaJ5hTlsryRjDw06aIojqFMkQcXsMKVMQm/4nya
Px6VjVOHPXYeAhaU5iEnZFZw0mw/m1CdwM+kQCm4uIuT/yge2arC9w9NK+ySCyZ3
pC7F4HNzKsZj6a7mBDAaF+DEHYNgZvjMH31Efqq/V8Znye2X3uJfzuP9ejWLkqVy
UrSbWkjllTAQiO1ceZvgcXyg+E17p4bEiGgDCnjknENboXTSF0TBfq7F0AK1/3zS
2rd2anIWpMg+Wk/OJHK/4TPbz68gwuCDkIvvNDRBSRLpODq0Uxg7tmBERX7Bf0VX
XoIVxlbLiJGG8XTLgnWcXCYOCVCMn2n3hhBRGfG4TRvDOWk52Nw6p3Slq8ZPRGMZ
AC5PtQXMn4kn3atvphFmtxgipVyngnyYCAGeTnnaV2U4BMs940/eV4YMo7dmpmdX
QZ9ReW9WwOLM/2EaAZ0YgoQ+g1uiRrrte3qiLHHt8wIaNaPj/mmvbMS9j1sNUhPd
aLtbKiqKE/fQ6viozxv0MU7vvIQezHlMJDkYeWlAwNnRK55gZeB81ab8DovnoiZt
vgmcTUlw5GZgMzGjICBZIJIKvA6de+XOoYGGbMdD6Tov1Ig9RdGWdPlXKxvnl59G
vry/e/bosBe3yqzUVDHPkzwxm9c+EOjE4wvKIRu40LqcTCNwybMgN87HGp8eI6Y5
VoCUmAvWrazlxkT5aNnhuHwPNzre+PvcF+EL3+rRzuSUIjKdDLn90wbaDc3FgLxk
smnGdxCexL9wRf1Up9L6GnMyr9v321BTRdjhxB+82wM+CnIKCp15JPahwSd2/wjo
O8Vh4WhA/YeR2JFwVvDJHCW0fIzKH4cm1V76g4Ht3zmLG0tALO7Q6O1Xm+5MHHII
PtvSLzmQ3qT/QYadYD+z/jaGscTpy1pnp3pnf38xcOKSL/gomPDJhy7t5S924HBV
AiJlfHFQF7cz1ACAObSSrPbGCAR5g6vSrfhNRH/ibcuLfcq6szl+jB9/UFxDtp2M
ZJOw+o32TW0cM6pF1xTdd3rhDLjK5WlwstHlYBkzAY3FurnSVLTjbzgz7HcO3T/X
byDqQWRPFrWwzIo+/O+DGP5pDCc2MMwNaLEmffOZRk0xg6BBdLbLtwNOViSke4iA
sn/B+IDlEYmDX5MG7d27RD5Roa42Mw9LU2bb1ydxO04408T/z5di4JkhrJdwIWDl
hpf5+xiceyaA7gOxyfkzNKNeMDAkD+B/EU+m/ILloJRk5jNSlJf4AKIG86h0ikcN
U8H791bUabbhKxuUy7ffW8W97pARiRB9xE1lPbY8XyCO3c8msJ/bGsgKaR9NnZI+
p4MDhr8NOwLVSVSF9UJkGAm4wVWBB2b8v1Y4d6bc/ADIozSIp4+Loxd0+XimfNHY
LHDVI9AJXAP+PPDnwjau9HRGsAmwjTS0BllOegJXcLVSFgRrfD/LvPRvNQ4njsCL
Ba6TaSRO4DyDa97laacvWdtmNn3hw69mL4Zt0ZxWgVj5cVNInKdSvpygHHkFbwL1
A/jDFYRbzR55EuJt+pN7Van3XuptBQCHo5ZPZ7Hm9X1dTP8JT8jwtwPw5VNwreK8
j1b3EDhWQ/geP+9vnUhb76n+O6G6nIFRwA034wHYfZUWppxOMqy0bheI9PGkk/FG
EVCVZgFN49xXx6RaV5RgCKRH+4SuW35Lvg9UNBIVNHNG30JeC6D7KB7/DQu/apa+
31vOaTsXkvd6Nq3jCs2dxvIkikESLAmnuz0KW1vmCaE7UgAjtGsLXvapj0t8hMUr
mq42A2T9mLVXRTIgimEWbzHUwcK3mLsNj8WixBa8hWFDmR2/yHDIeR2tANmPwjRU
wciFZp48HSD/2+yS4+B91KqJyW+lid1tXGBlhrJcfET3HoPyDCumu33bK+9dtNcg
OAvTBmzvJKsuLivTuMWXSBHcQaaheIBXNPN+AKw7EHyXt/wQfBfhj9DMAjFnWy9c
SB9/z6PX8wDI3sQM4ylhfQhQK5dZiNENWeThtsT/5lsP9Lv5Ur3yCX2pV439MsxF
QMhytu9b91jrowZx+puec136T1M2xs9W9DMue7K8WaE+pz7q+eEthnQKYbH/YQLe
m7iz/8X5ifdN0RmOWGzqO++jjMVnvm5dk9xcJIQ6chs35NKtMzpf2/xjjYEMmNuZ
c9JhzUFGMZTALtbl+xG4BTDoar8CoYOdCXP9z7HdRdH/ZeEj/spHhry6y0oa6ewI
bocVhE2VVSgqlAQ/thTijUP2tJDbIT1/WIvqHRu3hmFgOP5E+Lhmknp8SgNasYyC
JDsYXkPwpBKI5kicXKcz/EKeOMhnk/6qMDdlixBiWII3f1PWA50ehkHbzxyXUaXl
6iKgIBHzbyb/1liMcrgcJ3lDb+wL2niGmiQvdPGgwvoI6KC2hcCmhIq2AITlkykt
Pxm39cRsdqV6II1jMBXPM8Rm82gdTLMtFgCf+Cp3twaFksxR5t5bEiLEQQdjRbfE
M2cneLlPIkVqDvoXYl5mIRyiR5K3N0iW5ixfKRGWOseFXRnwCmdhxff5TcsuZPGG
LbslS/WrStFuBM8UMVMAOpxB81Ff2ZA1uWIxsQ73BvdF/WR+o/CVJ1JtZqvE2NVt
k9ShIYyYjEnnVf3zJzLMS/8tDE4QI4lYUfogXifM09nI1+gqsqZpmiT0HamgWuwr
jK5nVtnOYO9JRrbBXvqGp9bHv3SOty3/AAB2GzSKx7NXPcBuWoOtH0HxaFg/dyrm
2tqNK2vdmyjniHavlQxYn2kGCE0npo13EPB6Mk0urNL38vEI9MHoHAdAvNsi8GnJ
Rn+BTvps+QKfLh6N7xvDRcgWlaf2USSDODdv+ex7WWAsEJJBLZYQ3fde+cnbIcRi
jMKo6ISGnZcE7FSHDGc6iTMZ+8sGlscL9IfZqnKJEs5NO+sXwX9jhUVKletc3GFT
KD2amRfszmDyzBOXb5jK82WFeKhSf+sJEOODfNCI8yK/EeGAX93wVLAEO7Z5dgyH
0E24Ci/i1DXN7bt9xEjNu/We8i+xEY+QiijGjx94dlWffF8v0CvcZbFfkxwzjP0/
/hw1ujsUMy/docUKWK7vDtYxfPEePxRdo9bg0YMgVSPl8+TmuFwUy9jO83z1Qc3p
aECsPqDVBB+9KTa60fz57phIWqabD/R4QzIC+nj0ESrn4IysT3JZKMKUry/4Cscm
hw/auG++gfv965NDSy6wmeXReKTTRWNFaHFTy63Io+NkYQPaiiqjZ1zPCbUsFem8
+Yd3mVW50RHqtLCftFxMvstMkRNt6UfKcBxhHSxylST5OWyMe75uCbN7hv+M3G9f
A7xo+iaHsB6d3zG5E2o/2s3THKdUKeEqEATFh5S0xs+j1r/5QY7Avyx0WJRVGc/X
s2zj8vAyAWe2DkGBrV1zQBjlKceRhgXaRBSlhSHzBtYOcSk3D02gPjWPAevE7Q2n
5+q0YgO9MWoMh7lFo6wiK8iOCWE5oGogPb6+J4aN0YEnlUYOIBVJ+hAwdjqFBqCD
lrGQ0iqBv9FI7wGzU/t9TMy3+BCFh+KUA0Dn4zBujx+ZVAcfHfYRI3rJG3kvot8h
Ft9NMWmFnNsAQ5wctmzYT5YS9LIOC3GaODrsJwR/GAgXPza8wjxpa1qU524S/OgS
DEM6BqcTwcfybsqOUNIDIrghJ5zmIRblF1R+DsEzna9okmmwSKkONflXY4mi+gFK
GBzUOBlWcyJKveGJUqzcUWTgky+qT5G2ZPlBI7aVdiovX+klT9ywLdtBX9GbcHdd
wumdw+oLys5lmSZMxS/V+keaNAo4qAewjHDROzD6kGgUaknnGcfgd6OMMzslrwHV
i70hYLrmSGx4RB6T8ZGAYWvVkBPFO1xE+2lBAJOYVatHqqr87Mb5Vy76+GJQcuTS
/KBukVjSttJvMloLhGRk4xFpQBa0o7lD31dID8a9YkvjxGGGBn4eqdV68ADoE8e1
19OLIps9x/DDwNRcVIZE7M9iXkH/OtAx+1yO2qKHVjqwaQNhgfupqvKZGC2xnCjh
1i6EO3UOnhY6KgdDhQfe4CHUkNKeDggD+QHC+JJiVToBVVWGYsZIG4iP2z9aZ6jR
6dp9FR1w2qWg4lG/1Pfw7m45anTQZytVMvbYZsyRQAWO/PyH5NscImCR+hktj53y
nIHMbR70Gh+kycJr1xolsyXi3feCOLKTPjstiQT6nt3SuezwxU7U3S4u97u4TG3C
+FfFsdJEmk6OoVNm2hwAY0B8IV/6z2LHgJHL0uasvfjn4yjJCP6xA+529X+/HWPt
6M4vw9k4O+XzxAKmH5E6gGlKQzP9l6MaYZWLpDiSZAxlCqYV0AIz3pkey0k9gmYs
wZtVybUM0WIHnHFqBy5rj6VSWxqHKp6RxvZT5SGD0kb20cxPELhMKBgsbNeTEMC6
dy2Ex0WHoy5X6YoxAy9nctoHO8ZtbBjwxwfVp7sTWm3MSiemf8qR3xcrfdO4G1sG
v0fpVveq44tGvm+C+Wfsw2N4nN1RK7FQUxVYqekacTwNH9ugT3LPaA9dmu0weyPc
+GlVPoyCbI5KChAeVZY0qyss1hGQjanomqQO8LgIiXk3WKBc/Y0lX51Hm0BnhyCV
CfdrZCwLoOKdRSN4Mg2i6VzPvzxF2FdRvV+hhX7PvBCwNnlgMZP13jJ3cYZ/diMP
GEQlQtDzdwDDICbQpGL1RpUru8p4V+uHKj3b5zmA7bOFowdl9iFQlRFvX/jqNpXX
ruPr9Y6IrydeZbiZ+cnyErT0+TOdeuoTQXUPuTg1kHoSU85idaSSMkOw2j2P9J/3
wfV30tEiSlrLWSO74MQDEskc9+rLVuZGESAOmhX/iaittDQZIlipY2aYku+9tkj/
pzcHcNlM72RsUsrCK6AHLwhzteqIAzKHHujsAERwKlpGX4qcHvvQEoN70hiKzT/X
bAQaGvrGl8n5ZnpkjmM4Ik8mDx9QfSbqYkiz2IKgsTAiTVMSKOSAZwXHDxxCgqfd
AK19je3GO+B4Xalrdd0r05zw16Xsqqjd7OOW1DpMYOu3wCZQnGtnpTWRvnw1XiPc
ECpif+MkAlYv/tn6VTNrDcZQyP7qH5steod+Bke8NJJ6+P+Q7F1OW20olPC8xz83
hhAqDs0Yteyo9LHpA2Jh8KeBZM8VpQ6DuhEWueLIzf5lzpVneqGN8zC5AGLtLK9u
AIQs7cRK7OdSyb+cUBVy2mCYH1QIbrtf870EA4OfqpPeSt3ONVOsU7+fdAT9dETD
pIuxUuZAZu6Ca45KURyF3ZY+G40ppZxtoFHy6g9fC5s=
`protect END_PROTECTED
