`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/T3Eyc33h+ku52WkMy0dx6uEQYyDiRx3S9M1oS/CQCiu4ErJBi0xq/HcFaNzWSoP
uHl1PXcptv/WYvNkNT+zv0wYl63d9db90sr9DFJrVp+WuQoWSNRcUb1EoJynnqMA
vEz0X/NIEwLFQ4/ixTFZp9cVAIsWdF6RuhvWAyzBLcRAqgiOgr4V/5dzX78GAW39
D98KE7Vd5HqfJw9vFFBbvxjZJlCAW1FmwTTIdtdQ2ZWc7K23r7toodtfP7IGtLmJ
2uDg0GPrzy7mo5PPJEN53SzcOO9z/WfXO9fbLlbWWOY9uooWGPTBvwkpQWz9carW
9eOR9udjVgD2bGTZUQYo3A==
`protect END_PROTECTED
