`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TijFWdt/mY0lwGa/Aug9QrGdj7SiCxqrLQtpBMMpD/HVJ6awYMKi/XdGSKgsVjA4
+rpgx8yrItRJN/CrIOHn2UYRZJZdN4oSb9o9oYcami/S5W/ZtQSyF8QWdaSaVMNd
ayhe7AItFetPTKJZMH1hVIVBqAV6fkpDlr+2sVDnpEWRQ3sdeamA+berpWQW0q1i
M2q/LkbtSpXqLn4iYG7a2ZUdpPQX1ry5t3QrNroUd/ZdIGQSqy7/JoV3RRlW8Oyh
uqsFUFTChFhkhFipsOc3IcGtP+fPh2NTXTkslXyMZ2bXfmEYZ6vJRsVW1Yb/3YzB
F5NWHePBQ5Bm8+OK58Bk+nLj4EASphDYybw5VEbf8yHSM2696F9LVVw+xG1GvLZj
Vo957Uhqj5fNhTMGjjfQAZiacyMhmlXzQ4A2NaHkoKCfFXVJUi7cYDSdObNfhJ60
MxRtJ50AlrSmr5TyGULCEejqA0bCnZQUEu2JvVGio/w=
`protect END_PROTECTED
