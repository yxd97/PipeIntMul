`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2I0q3WurYcaSTuc224chok53WZS9ExBncTBIEQfLSfEt6SxAppopH7chIBDqwU2P
ewK7TJ4sY9SC5TvxBLcal+kYJOXRcQtfmF39JxJPAY5J4+tUmBarrImC5mESrxuK
m2IKwddL6lCcmZgC+IEtH9Ev0tEfE0hJnFBahkqSxN51ru82mwCi3q8piV5T9d08
V8HlmP0DJP9bsi1AqWjDGCoxhwFHNlVQsO/8OglTZzI15BhQim+6kk3WX2MOA8Cg
6+1MRRssozx39KcVncyzog==
`protect END_PROTECTED
