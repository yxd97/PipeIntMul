`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgn1ri8Yj2PBPFQP98Hv1l/a69XvrHpHr157xOe4lbcAjUii3VWOMrZ1lIJNpJGl
fY0DU1m/x803RUAIV6MjwR3k0bTPL9hPXBLEvYZd5BPL9MYPEAV/m6VyLDV/1vWc
ZzW+VywRnhgd7VmgeJYoz25MTF1KB+IGiH/aEYTRchtL4l20r0O7GYQbtopSTvUP
vFj6CpXbMGdIDS5NZuCHK98erZlswL06hClC7+8mzLShXC9qKJaj/3Qgay2j6MnN
VQgy/TJDobl5urXSGd9EqLUqc7W8GnOqdNFn3hvEn09k612eUc/QWiUQHaRBZFkd
`protect END_PROTECTED
