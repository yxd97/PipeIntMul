`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3kw8dyK44/CMB61DflT6qu+lk2XvCvSS6TXVQJPnb6AkG7iek+7pFX5dtSfnDpU
dAY0HYOFQFCUoBNG7RXYsSEUU/g6Pr0odMk4jnXGjKOUtYL/yIZRi6qnBDil5aKO
6fBlOdJ/CboN8prktIBZfIVKrDXGbS8UGK08u27wdSi6Gdf7B3vXJfZdhIzoFiwv
Tp2+1bFw+7bREX3iCLWqbDLdzEBE5Efr6F9mYnHbOoIUVTexv75q2UINCvgD78EO
yxv0ieKRIZzYLefVii6Q39jLp4ijWQGb4SLqBPxsiLOr6WUrbz3RbsK8T3rqICfM
dVFGget08rU/vl7eOJVXOD5vutA/6jY41K2tFhv9uHnnRIVC6Kdse0a7+w2gzQDd
M9w70kFHUSMisrM9ZLD7nBk6TJTILGc2d/ZUMbQw86Zpku/646tKeU/z3BWJU3n8
dwDr7Mi2OtMhfpKksKL/Lubohe/9LUqp9qMqnk5B3OGNrhAv3Kr5dni5VbfR9lsi
vq5b6U+lk10Yl6PKA/VabSW110z7uqApslqQZz4KTJpuEpOqF1B9KpNPi1YluoNL
khHXFGOdGmMWaC9SMd0EXWIW8Xv/bZ/fqy6KQcewLqM=
`protect END_PROTECTED
