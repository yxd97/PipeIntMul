`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s556a8y4Odsa1WNq0divNkM3tsP10eKORTxPhq1UkZcML04imMcG0QJfTRUEykDw
B6f1HLmOJuIrPadU5+J4H8LoD3SdyBvWy6nuNkYzwNf435BisUvdCs1M/yq05naf
KKWuKkMjJFbPkh8ddekgHWXbfEG8VJhjSW2edqHnttYezZN3gpmHR1pnyMs02ynK
GLkjiCakw23ITFQDOE4paIyJUkLwhwTl9RhTrOVrEFH0l7JQQfgwkQPHlR3MH0DH
L3ynGQrAl4stDA7iPEX4K2gCNKo9uGQL9Zal+XJtjEF1LR70mbxkTMcHaqVZe0H/
VR1qTT5Fvf/vkY63RThuMhcru8kAjqbvgSNWXN368trymDtxcWMEyIU1Ts+ZhXxJ
A4jJ4t/M4vcAL6z5cqCCoAme3y7AqVhwKrwa7M6e5OKk5LC7m7iDmBS+9m2IEem7
aGFz1u760fAomwIygYhm2jN5t26m4LAp/0umgUCfibUY7oKpw1aBWY1LuADDZzSO
RcIfdBgLCVPLGP+GLtMBeLNUKpF9ZY2eP16dvpBSPDLCyO2zCn3YWO+8txpEF4J4
7jJp85m0cGpiGB6pfE/NXSVrT6tv4ioWr72KmUfFTRCTwxJjpAyLB+8OUmMHo0CI
mgOZAfGqOIt4SKI67lT45oFvnKx6EsbVUeS36aiZjPS8IFIGh8KvM/1TOIMO0HPE
qIA8joo28QgTJ8f1dATEr0/G7K9BLVlkMdh3po0IFK6dxaoQiyZXow39YVgRZip2
hhefZ8rbDtrs6VC7n4YWBCNBaYPMyym3PGhuYhUcB06GWWY/Rcr4XqXHeOmqb4C2
qNHPQOgxIWb1UhdAnHeVINePUw4JBiUSp6I3c90iq1ODB2wYK+Rn8me92luAb/IC
geS7MBy3h2lkuN30lk6rbOpfGtKDCuLTMszuki1IZ0a4uRvbPcsVb+fs+GYcHYco
if68b3pgCgcmdRGxt3oz9A==
`protect END_PROTECTED
