`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BROms4kj4FBvwyxDpvQs/P1R7DKh4avzp5GhSVFaKdfZsFzgFoMPd4HXS1M5zYEI
xvKF5jhCgiKqkvy4vLV/dYZ5f3VvjPZDTFue7ZMMrnS/CzTkyAWNJ4TZEO+mmoLA
VWIzdHtfXB82m3MM4Rn1e9X9176hdbTeuc/hEdrttwIjzc1HAUgbWFIU2/o/XAo6
dyHhMkOpe9JYbJjg0F7eLEP0t7Tm4eK0llFJEbln2E+5GdtBxhejYDOVJOg0M9kR
UlQfmN1rXLo+eAjODrU00Wi6qRoh5WP5oOEgbuKHfG6FGHZngXIY/3FdQguih4ev
+3O651iO0tw7X51eenv63RCuH9g4Zm8TZiLsHYRcuHVPHrX3w7ygTUeotZg3n0DW
yOiiy92C3FG0QmFPdNdcII5EweXT5pJBMWVZQFJw7bgfSbGPwfqG2LoRjZ5hRgMi
+C6wbz8MWZcBDlsNbeklr7bxNTVthPgMNpW+y30VTU54u07hQ/PErIS3zFPD350M
015QmbdFIUYj3XjzBqUk3Qrhpbo/YKRAgWaJ/SyT79a48Tv7jkA/ZYMerF7lQTbS
sToZfIAIzrQZXigU9s52wA==
`protect END_PROTECTED
