`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQDdtT1ek5EAwEYwQeYHkt1KfzKNMCHzp0hLi9Osp0agJdiEtzUCxF/JzF5OvwOr
yBpmLJCSb8AW1fOGzIiSiSW9pg5hAdWZ87jvlrFoPnagceCSFLnkVSg8Ib9CC3it
M07Ok/8JiuCxlw8pgC/0GrqQO5XWU2fkCgOuNWB8MRsP4NesH8sKiPFjXA8gB8vG
61PhOo9hgE/QVHx6hkzndvwV5r1sZAq5/01EzETvu8Uim1g49etUXEo8oZMs9TZI
U3qfU53vsws9oRkLui26SKJlLQSg5r5n5fKVJRBuIsiGCeQkOcUpCFeRczUVgrb6
9I8Y52cc9W/ho5iamaCApg==
`protect END_PROTECTED
