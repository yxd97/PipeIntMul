`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
639FMtyCkJSbNPFYmJuyCOILgRmS8m/AQLyLhyIp0Bfvxx7XAN0v2AWmtPusCAvS
C+mllGBB/149FqBV5Mj5R44KjJc50JEUEypUvefn8Sc2fELDjS5nY5EpmIShtyUf
nqDIFCsFIyE2odbY7pj4zGVjJ9w5uWzAZR5hw3XlaPzehB/H9tlA7xqaeFupIZR4
+cuVcL3WcAV0riMa2Rzs6AfbHya3VJZX9k47Mbri7wuz7/yHYtE2lZ19UX+4SJ6z
m2TN8uIUaOkKGGa6xxPJoTHPmyL+gRUkhMao46kCLixNBTxpbGBuctXw7IzAsrEW
eLEA2DJz8506yX8Y6hhNP/9uhdaQrKHKB0UQ2ePiYOxP6iuDrkY2Dq/FGNdCs8V1
`protect END_PROTECTED
