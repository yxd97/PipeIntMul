`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
trJlzXW7fsuUvcgetwR5Hr95WcGx38XPYHTKZ9x+jH3Ek49jtfnEzDUOEypm73zL
Jdre2AXuYU5204v4KxiFhCZW65FOKJH1LlHZ6ohvzhwnCPm1THG7VRCc7wAjnTCy
hX52U/OFY/3Hcu3wrlq1Cd5cV5gVRV00jz22FKoLpqUG+688dH2F/AMUAhL8VA0x
1a6SLWaPIKWjzOU/O7mYVpvTIt/KVMOMKbNkbm7Omurmlu1VsyhQuUH8cxQqDJa+
QCNr3BLLPLXWQyEiUHdtsBPWP8mRpjmTu7fxfqv65wONHosvrBhpeCaJfyqA5Js4
Us/BepaqNDSecIE1kP7YmNg5abWoVBljkH9//RQagRCQ4kXDI8740NY65Ki6f+ru
BeujKJb+zLURG+5MXXVVzTpi1oZeGdAFfQuhDM3hyB/hhh34QEwxxmoT75dMK7nM
mtYoAE9uh6fQD1VpG7oGUWyDZp0nmDgEbHjxMa+wQSWWxfGvFR2JEnwE2VKIbx3w
we4fzUIB52ePtwVvz2fFK4kgZCPO0+fBqs8MvWlTPaxcaEOd7nT+IB0TtOczBXqy
ONd2Qi16bizm+70+WlRoRJZrUjioEslujnrzM0nwzJQsgAZ5a6iHEN1ayt+LQe8Z
WWx4Dz26jFY6QW13cYZz/f/dNWpDxH4ra2akGCQrsmUbmYkG5WRJJcfoHWqZJ+v8
9iqoasvY/1T28JeraIbEURZHBc1fAOliNIEUgd3MVAX+fabUXvcUyV8kpLbCCZAc
2KpB85KFU8hVWIXcwUSOPAChsq17qAbQ5RPmvqiZqMT6TT7fJ/m5lywkgooO2JBb
x63qEeOdIsaAs3reNt+ZRoMZ/KvypXNbeBcDKdsiiEFniRZHF+NZSqikchiyl04J
FsMCer/0qjiu/Y4T8cxjd/mcUOMMH2oPTFYmliN6e5x6GKrnIXJZiRBzX/KFN28j
y3TTjKDlB12JwxPoT2cedcrG4DWpGzAVg+Z5Dzwk8Q3VsQu8MaFG0l3OfFhRzTJU
g2kXafHcNuxsYh2w4iKRx6B0k+4hwLw+1YsPO9MvZxsKmCuGI3ANAwRIwUvDcZVn
FWnnmn7TXQXItm0tjiPhYMs7eFCMbNpTD+mNsNILfTzi9TTkPkSfIzz3xaDmXeuB
CN1vKrbdgeqtWnEFUR4hb1xNwbjrVVlj3BUpRsHuE5pbXwUkP6xd1Dj+qKoghc4N
VHjQOqMkXj5chM/UMX+ZGDKNwACnLN7JQ87loj3x917pAJUlRYfwrzudRr+X2usZ
VcCxDeBP1Mu901y0dfeLFZ0XhzgZhRk6zw2+ujguEFjMLREMUHHLHXeL0BFEmJKD
mOqKbU0YtW7F1mZIXoZOSibnFK724VhugrTrcmFUhAqpCawlwZnv/4gmOajTNngI
zTrShorroH+Pkc3TbAm13pDcsbJhdZ7p277bfKpyifqYJ0Bw0Y2+vEiGxkrRGDV9
4i5aBpal5/CniArJB1ezHi9YPUS5K4EKryF9Fp4LilSeKi3gH2F4GU/cMAniwpMI
pCbOhQAgny9naM4o/DkAGaaIkgIScIGLAQzPLpSsZ0HsP4gMcKs5pjtvYEtiT6P0
CmGwA38aqhIioxYjqr5dgof8/pM8m0Tviu/HTWRDr7fFyYLhCfv0GHsEQ4rkrKnt
ziSGEms+9pIP3bekwtbNCJvAapq728SRrymReMx9mRQ3L0opU1nm92SFdBkK55Df
TCaLfrO1xQnQR2T/LK8TKnBsSxAgqgZhmA/dFFdGA6ZMezynyjF72iHjUg0R+vkA
RygPpKXepxu0p10dme0g1cQEF8xpHuSNvAikXY19QSv6zi5l0RTZLdFSgf06SZ/4
yDvw8L6HgkoCQpmGKSkbtFv3QxkuCav4i4TvPe+tKXWLNGQ5QPCOYKlCAkTlE1Jy
ufZXsGFBkCrhIbEjCHCh819jqyedmchYUBp65JMPj4VcNrUHQ+pGi5ThmNtJj7rm
6OBn1Dy34bfAMKliZy8FmIguMEBV8C7atAR7GPfKZgi8PHcN/TvoRhiN4Kag0K2v
0LqvwDvjgwj4oysLjD4ZkgBh1gL+qeh5DxXWX1PenwEfKOWUcZMOykGr3SwCHy1b
vTT6b48Vj08BQxDnPjJ+jluYPHTCl1SbIvsAJz8JdG5R+HPVYa0Ukq4JtY3avOD/
3WIVOVPQ0z0js3Jo0C7Q/ta5EPV1YpIAIsP3l7xP0taOPrQM1LHSa8XE4xiXQw/5
pLyFyy3YSZ8W/0MeZvoYvsvirWiStXa+N7Nd2nDqeWSNe1gaW5HB/hSe5KkFjL9S
kOCP8IWIaJG7zvAAsqdAsjGWArHywPggXfZQqP3Hf2Y6fzCWZqMrtc99suPnNiuf
F1hvZ+zEzSaYEFDtcLVAo5i7/KknUXMnwBKRM+XR7J3pHYYV+bSfrFWxuAw+TyHF
CSEK20WunlUe0BQc9bWUNoKWB6vv5UOj7AIUlg86JPq7ViTuE5boQzbWxTPgmp+8
sKPZbN8FHp+7F0oFYpo9uFxndEl4V4D80IaT289o0fUL/o12ObCE4jTBINnK0Eyz
hfZhVPy7qaH4cQALJHKCA8ulio0jrLONBpGeW7LCYclQMvmbHTFXLstrCfF1ldM9
QBw0EkiW5iMDUlUH7Vak0j1v6tb/9jyk2zpo+0G/KCv08y2MDwbQ0/O7+l7+i88V
64sIWu11uE2eYQoW033oxGXmk0IvJKfAZ3qDYoNvn08Kl/ykwvACA40/ZTrc/z7u
CDyS5RFJyd7DZugLjy2YMn29Nn9i3WnQwPL3HGzJXHfMiojwxwkGMg2ipAg6Lq+G
91UbwpF5Hp/0mDlHCombfhrsAEBPBofG3VNCkorKTyT35pOUaOC+R+S2cDsKXhmO
rPykcv0LuYoc6vRmGxx+0qL7GclQCR9/hG4cHX8vwKa3wn8ZBlI2ZSlSStzePFP4
n7qG9xu68iNodlq6VrJUkwJK3BwzsrcXymQ4/wNE4lx/322Hue6FFCxm7PpDDFym
3E0PnwhP31GkZQ9U3LJdKBotqFc633rf1bdBanZ77FmW291EhkUMx2nimV1v+IOA
/c1YYsZT3l2eCYlirmgdTkSIVjZW6wLCg8IuBTWqexutgemrsfGqyFI+bcSwOl9z
EykFUt8dQLey/G+RhT4H1qI1jx/ufzHFl5ZwNm5gvQiIV2MtptrNYJKWx6i8Qq5O
8sSn1blv/l/Y9WUxw2JCDX+dR5tDGL7jcribhvPlxInYxZihRxWhhSOTCnuDmYGs
UfkKxFBLFpEg1nbls5Fp04d3+DmgTO6UFrcqL4QnJM4PmNV8iCqdEjOtd78se2E5
yWm9LANAJRBHgOlhHTolBasiY/K6U/1cxN8UHJHyM8pH+HSvNtoOuAPblkg61knp
y1IZrapuy1SNQ0+xLnQFQRX0Zm3waFCwSK6M+s2TsFv+ZLL5YjojxVuUbRiRo+Db
l0ErBSs1tT1KtYPHX9S/puAYfn3ViK29zYqZPJ4+U72uvTT+rDKYcPkrb1pI0O39
crBnMfdF6oXvPr207qCMwA04atTMK/RpawagRfFHKdsWSyvUhEJr78D53Lx23IwM
8z6mVqC3v8CRfEeXRt+QwSIbcsPxzb9MgORhkj6iiGs=
`protect END_PROTECTED
