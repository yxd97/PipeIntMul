`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ew/d9AJ17zsCLW6bplNZdXkl8MAyxYCTneLCI5Q+RpOa3jzZXykblcc4MmTmR+Q
PlcUtxYycAf8BZrBtCJy+MXloaoCkCAOcxwTJeGUGBT22cZTLxEMvd3z9+iGC1cf
sIvLd22DHCRa1gxNbsUC+ywJfUKfVD4fLg1CsLt4Q4XyeCAW5XG+zTqsxHxwqo1P
+/UJ5NQ3sUzGNL2bRn2PIx2qgfyk/xYgNkyQGIngRlwXIh/29/Ya9ulKmzKHEhFv
NJXw365MCWoVNVkqJZHX3eZLHQri3tiID82apVKcN6dmxB51WFyWphXlSY3wx+0z
x/O2BBtelnuOiYOG/fXzB/VkuhT0dgYi5RbSlvzW/5ThIE8nZOX/UZA3QamwR0lv
h5OKFluQIeu0EKiD6XdS/J5L68JqC5/y0/vz4oaN6kSm+DOo5tp28+ecz67v7N1d
mQhgCgUo4nskMYYo2qOwdn5JKbebbSjHSCkY/FfITPcBpG8Dbq202wbgTC91NQR9
mcK408UFj8fBi4pNd0RG5E/8FaCJMYlySgFD1/IazelOoOSN8o7ppuVqDrMdW9Ek
TxnZ99+ibG+/yyBoNV+jU/N9v/NXSJIN3PIB3I8tnggv6HDlE++D04kRuzThahzA
ScCh2/tihcz828hSe7va26RMqEyV+t9sNYfb9BeOW8gv+bPlxTtJBGbWWqk8xrGG
XD1ScZ11Y7MsbJAGh2Gc5AFM6PumRcnqrxS1fEbNxxfNT8II+itkxKrj5TKNiHlX
PfkeC0UpoicbGxCulCqWsg2ZJL21eaEvvitRMMu6rVEh6a9Dat6v/fKEInpGc/D7
f5NJtaTfQA1kdxjBfsSz1+hW7UC1xRDFVNAbIr+954tOBtN5OUXwhHAtTGILo7IA
bfCHIMGTZqYaoYWl4HPDUsNgZhGskmboNpHc87GpJCJhVgKLWKJdeSgSVSDobbfx
zZyZ1kYhWnPZd++exuMoe6CWgOTO6XzSL9rhBfF7uY0i9ue4oEP6NFWHYcprNRWE
yA9qUGztqRjnEZ4mgE2LW6IlRSZyQqlCLME5X15fQdeWdGuKR/OmFxEnZ9DV2k1g
hXjSq4x65tenRE6s21BxU601MXHdkzA0w3OUsZsXNQ208Ku5rftlUcuT0std8+yu
+8uemr4M2dW4moniblmPyz9KmG9sH3urxKiPoVQ9geCPTGbtspxdbhR+wGd/Uaou
0WdfAbLAWsUUSXCGlLjSXBlhxFi5CCnlllXkc4SdakKls9JPR1+jeq8FgXfCd9dN
rCWF+gAtMXRs/pALqAPTaMkK/UGlju19AOV0Aq+XPHKNQZTxlsZx95AfFGq0UzEa
j4AJqbnhDvTRYxE2lBEFnV4enPIm+gSqdDeFLNHKGarXmSpXukxVYzjG0nP6L7CX
d1sLxqj5slEWwt+YZmeOnetEFOeP8vTGyi9piX+T5AiBK+CMJa013Nn5iSYXzCkQ
B+n4FXfXXrZLv08YS96J8OeIkrgIx/6elKwSnxnL1gwUViJA6idcLH9fIFHik8IS
oO5vpn68eg+H4RP9DntvUgyCqgtPbTdbmy/Muw7XuDi5G5ftkyVb43UBTME3tvHE
+HCrpoJ35pB/UM1OIgNKd3O7MGQAHujti+wFwwxCBeEAU+Uo5oIpVd56n7Oq0pC1
ABV+nSFK5/Lm6dtPnWPcwKmU144//tSDC+ar5bd+G76ZAvAnwj/+1F3OHPdrDMVk
3QeFfMzlwPDmx9UQjhAu/R437RGxxQ2iNyLa7S2c8ERkjsjKXmnpHmEne+h7ygB4
xR+3OTxEQCkVUHFrU4ehtw41fUlo3eVXc7OsusYSo9n8MjVj23t00afXigDgRJTj
rDDqo1uwuvJXKWQK+6Dua7WSzdG/AT8Lz+Mbagy/eHiXT2Tz0NCBeJWKNpab5oam
gH9v4r3wjkOoad9cIwQGU1ILgkWiu+V8U/n8qITlRoFW0GksomxQIwKpQHdLtEg8
T9NR9CiEvOZHpsvkH+xW+1Jobc3oiGXVU15osOhTkFNwhE6E423wWao0qEuRLwf6
lq49U5RQYaDjDbIvSF5VsYS84BiWjMLVipnNBDfusqTuvktRHYmXLiyElDQIGhFF
3Lqp6kxaN5YpUCfBYUK782Q0iqITpSWQON/FY1wmCrR/Vo7vsuz9CqctYpFWMZgR
PiPvHAxLSehUjQu8wZ36m1ngD6DauGlmixOpZY+Q9sutq47HBnRIzflO9L25Mx1t
M3nuxR3SE0L1xCwwhWFlPRi7Eho9qPpUZTrsFGd0x1+n/FpM8wrftWsiCOqDTdtz
AwvI17F+CQEuzfvUE4ZtqOqWOrPyfqMeRM2/zl0I+TpnGG4q9lzR361D+eFUq+9H
WuPfL8n2EVvibfC0GJAGnc4HYqkLLvDedYkyriZMmKQvjBPkecSZmaSzEEL9nHqF
nq/IQU+vK+3Do+mhfNI+gNrJtFfMMRP2WXLoSj2DnZev58Z3oRbGKywDP96fhoQ/
x9rU6vtGR2qkq4tPmyI53pnrYMwj6AmGY82SXA5N2XbcS2bBJvG6tno4DzFPNBk2
5qyGTkLEHpZhlCTpASYsKNTAfpxY1jduwLUCTsIOJj9UT+dURlWD6el2Ehdhvr42
sg9KyGATi85VR838biyBvsz5+JrE/V9lzwKMzwWDVW0=
`protect END_PROTECTED
