`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/6tJKYn+20HRDujl+58qMtGZlQpziv/TxhfIMG2vJAbqViBAMkgAOspNji1+jOz
xlUArgWizUZJ+6aCUCrDvfzpMY+V1ISNy+t4R40qrqVXCRzMCPFDIa48Ig3exsnE
QoV6t+woGHBwdwFqHLkJk3Mj2FTUAx6Nlc309sPb6losTzuouA4EcSsTyTpj2J8m
Wy98zuCVUEe75gzWlJzuru3VZfVHrHyLkDAeWnHKbBfivIFstkZu/MTjun3mzIiM
7yaRQDFwV7KC1SFc4OBtnc63XYkrEILPwAX7A1xSoCdLk5wD/GQVu89bkPAbhKm7
5zJp2a/rWnnKTUW9NMbtC9hyLAdLN/fyyyn6KjeHOHRlGRatDYdSqJfA9MH4G20l
J/fL522O3fDCfuxQOYjUWB5FcH/Wsc8huTbsLqSJql5Rdh10Vt12gUQu7F75xi+u
2o5E24O5n7Wo1CIVNjZ4p1zsjkh6frY7UHBr6tSKlLAjBsabvyGfwhzLTpeLsAU+
hzVWq5l6Y8L/J1bP4VMfYSogL2bwdM61CXw/Axbb4S/4OF73jK/4SW383MDIPKdZ
U5mtRpSG97Ppe7nKEfascB71T4V4A9riU0Vr5Q7O0o8ENUn8McDWU5HMrHbc14i7
vb3QwEnnvM3z+WKvHDUeOw==
`protect END_PROTECTED
