`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0sIly5TQ/UO5s4d1jFp+pxUeb+YcEnIe7mFJo1/qFi8EvfMzBCn9xU1jewiWVd+
oQIacvcR0gy2dDWe34e39hC6DJOJAUpoBI0pKKZmCYiEHJ1jHXE/3O+F4kjAJ2mh
da6VKfwUz+jIIc9qhGxB5Sct1WXShddTqAkUDL2ETo3EjXq+FdRHWn1fD2y5O3Wh
hra5/RawQsmMthiRq6pnn/CzJpYrHDVXt/uDQVQXGHC3Epq3Vpj61iUuZT8x7P+C
K1bPqZFIjqrZNbvUv1Ozt3yOYLF1BjhozOTgZ+zilh0wtWgm1DsC9tsvztuPwfJh
i9Qv1um1fYyHwS8r22K2Aefwv/kBLMHvJsmidvkKiAp1fm9OuIH23SjgXMkX/Rkh
qQo78ArOAIxrHO2l+49j2Aifgp339+I2D6aRB+hpXWz3K7KdoIAKPMFDTI9Ojk+X
nlUGYp7+pHnr5+F2S+3ptWm8bAdP8rKrI/RO+EQoHAU=
`protect END_PROTECTED
