`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4nmXu4GScjg3Px4KCPw73NhnZKCxuZuG00LFtenxhYWJBG0aOOxkOg3dnPFGXuWK
cBJlgPlvRQW41+LcV15AH0Ei4CcCDWfHEwI6koDO6yLsNGBxou3aX/KwP9tKFjwA
JQXvvdNYXA3Us5umMmKUfJB7SQuTHddZ/efN8JKeVwC6FJ+VbFC3jiyjzEVXRnl+
SZoFqJjJ1jaCn7WoWNCO+vjwIek1TA5vX7IqM7ewOd/Rvle7ClGvrs3qxYKnzn5L
dShLgiSw2H6/5oUu2JXg8yLU+hgQtSQjowpLSzIrMpJnxBxXNvPgGIOIrf0WHLZ7
60SPiNKR6a8AKn9uUwAY3zK9dkGog4fJpJJfVBJmARpySmyXN8SwEguJdMCrc0on
UBifT/g1vUB5wzUOx+dufkVaYwEP1VZHccwA3I54ZDpauxkgwUYZZw5mdzwq2rAU
qTRPthxiwj+OyK/G0EyBDSGfBJKRRf7uwyoo1VnDn6RHUyLRuiGnaIR/i6QVTF3V
Xby5XsgCZNEok4vYuiGvDEDqdIKkOJYS6inalG2qUgJ7cT5NTHKLhDLTn7a3bNje
eSsBVarZnaQw9h6NWv7VkveC4cNXeKd6pC0fjmkt5CDO0vGtIXEXaPhoNN84B+gX
eblQfRTXBhOKeYMuY6lPHBeAqMVv8Y0/DTlYrtcpNSFeQgToA0Wi8PjRafKgWiYU
zBSGPE74rqXEycQ/NrLqjDiFLtHZcdsZDuwCb4s39laiaoQr5KkaSYyJL40Hye2s
wysSfmO2FkuBhD9Ojw/IJ/XKlwoQryo9vk0TmnGaMxNKPLa5J4jVDSko07+JkYHl
SueckvhmVv7XSCnfl7iAV2WMmzjSyW/t/+FbSo7k3fUjB5qlItzVMA0Blzcz7B0U
hcGmRce4yYglzNFGviCGq12Yd8wkvWKxOpZiZIeZquHbUaA++A8lcAiXmMw6jlrT
kRW4v/bQZFpVDlWNZA4c1HZ2KCdolyKDkqKKyfVWKr+D9hHHsr9WpGypbkLwj+Nr
jljT4Y8lVOGxHXLEm1jBxxExW5sYHl3hlHmiujWzHivu9VcH4CQHToGhy6bbLkBe
fYVF16O1XpXKd5telKVWpxmHNGBrCsmdOd2EZPQzF9X6SimogZtf4n80SExxCudo
GQgRAjREK95z9QDQ4ElwSSfQ7kX7IV4MMJH+lEhpumaSKmQfbfiJF7SEGy7/zxPI
TdK79IK06ImAXtm3gU+EsPttZV0H4tCLv4MggfFST/sYh4iCZ+68VdSYXHyyFvry
LO25sjWX2zk4HiZyRUEnfZnUznlMi/5Oz9Kg44Un8910Fh369bfwlo5ptC09T9SR
9zHA4l8rN9nodjT4AXodPNpmWa9J2PoOyETbNUnruNfxz6BulMepxd0FKMrbfFEn
auX4AJ8rKY4Qgo2UVmOHV096G5yQwRnrcb08R98/TbBIreoRoTdf0pH25Gj3YF9g
UCsgh3uyY7cJcuy3MhFK9SBCq9VsxJgz00YfBf5q2bu4h6rk3wznGjlShUxg83p7
Y37r3htf+tgnugD+Str3dEzoBoUcznP5J+Nt99E+IspF86Jq7sfEDobPzgu4RswL
vfb9pBsrTHfc3JuiuutLQByZSfCPHrz0jubtcFlg8znjTVLJfQGqyUglCCiGGUXr
IUmsAbxnbRovX4alSRSYsGfD9UBUSDSTGQSQWlUOJUJrDngU5hlujFiV9Q8sDYYw
jIXAi+IL28XS7qQUdO3DDl8pmeudF3/S+6VX23d+NLQMxeto8AFnYwAQV4mikZC5
0Yhqshjw+6+FKipZIBT9YlpTY+1om0TawXwN4AiSxpbeHORT7qETngosk2D7q+yY
OrqI+DtgtjqpfbDvWJjfY8XMIPuHZEArFVjuC+TeKjA6ivuhRIcQWmPzLIPZD84a
UyMdjCBzu9Rho7J7Dhoi+X6uwWghRN6cyihVSIQyddWPBQKjMXn9qom7hSmYSbXI
LcRilMIOxuYBVhn0crlN+ysCBCZpVmSqoAOs3vMofuBww9wkJ2iHvvuMDdD7zQ/j
lj+bcjR9PiHYCCP2AY44UoZRZb9cUzKtlVLRb1xUQu1k0RB3F0Fwdyya44ayMLKt
yTl8JvMCpqiFILl4R6u5TIbAObQj41ELN6CJ6L2DBqgrGoL18RXqhiPuNnKHx01N
on93fgDOqqruuydEJzVFoGnTaMe20ntkZhB0rnsiRHtCtkf58AeVtHT5pEUACEzy
St7zoMIBQf/+uw6sool4qRnQ0d9rPFQ4o2rOxYigS+s8dzVvML8EUqW/PX5zgTla
sNe+E+SNBB/YnYHbQWa3VkBy4tl6CdeGrTpciUt2LGZ7xgpYfrITOawpbOV8tXRH
L4LCadOcnOxM0wGrf3vt8GqYtBQAge7qY+oRnxx1LcBa7vNu+FhRz+1dmGaDz2HO
ZaNwBwReuVyXsYq7PtCCPg/UAC+m8opETzfs3nQeNTjohOhf8BaawTVyGqoWK2Gj
3U60Rk7/usqxCPpJZe9cMKI2HfzkAZ0m4gLPJVCxAQIED6EC2nvWyoIG/T3LFbx1
1JklPx8qX8JkMSBAOIzIoaoju0mDcNNfYGbFPJvd2XF6Phu9FhYtEAbEcKjpDdeu
GsApXLIkdVhv5ijWCNFjheNQcXDuPShc2LYQ3MXWykUjAwbSysTcmTqN7ZCcQDWh
jcpNyhJHaonCp15z2+ZaDxuxBf1Fnso8YCM7H+N+R44RaadhyArcvDx5MO+VFc7a
EVjzVBEERMPUKY8OJFKpddicIz1KuzeYrLeoZviMzNfk+ZFvg7DYrzyUHa6zM1yw
c6gMhneeOQZsbkV2SbjV4ZkTXhwapKSZ3nxtE1acsrV3KH8GSYg/2/PmfF/iRs7I
qKYVJwmu+jGl5FvU3jp+8Tepj5b14S2QT4RgSKUphbCcGsNbbmnFHxGagTP+O4VN
11IxIz4Z5ZBCp+MSci55oI62otRumVrSMGeCXNwskhB5+qPIojBmttZJNJA0ke1r
xhDjXHv/ieA53c6MZbVSySxVXPUqThfZP4LGsIwNgeBeSQi/b8rzeGrrUo/uZWOG
3ul8aaRu1v0D2KXKQj84Qbuv7vhMg80dsDgNhygjpa6y4V/fwVupxANo1yYn4vGz
D27WpXj+cfkJt7MHm9qOqLEMTHnBx/GUR7MMwoO6hnXh6vH0RvCMVdFlfAz7fFGR
qqjH3UJ+uJMNoCWO0HlTLTatlCsYecCkGPEEm5JA3V97FCKtslUtO3UyUUuY4j1d
k6OZ1ScZ2cHaruklgO7Z10OccGTC5moaQvtERZGaZnGnthxB26UhVgN3GqWibRvD
RNirRsjsM5kmeztHA4JSJipcmRgcdZSi10/8er4N7y/qZxGlc8Cok74y3jMsASk/
kwIV/06NjKbFlhfFaBeg8MIVyyLCm/TnkOT6OpRGO0v/kGqM4Chqh6ANR/al6+OH
uUm3M6pOmYfr5d26IjvnQP6M9+JKRfaADkzoWFNR9TLX4oGNEUMU+UZajK1cMmBx
gzwp3tQuet80lmZUBUl7Y36XgkETGsQ9vhUs0IztmSy0Pe/Y7qs/cXkiFJgrXZy9
OlNfvefxuEwWW5u7uFl6x2beQzZMxc9TjlM8138I6HgUXrqqr+n3CKqxCBRqGlnO
bwcqRM6BV0YrNlnrVzMpSPPKFBG/jBE/T9xtJ7b0P4SbZ9RLBjXEZ89setVTIAMq
8wf2P61pdm72wSBU8LcKrJ65M/tA6Bw/LIEz7ht05sj4saoz+v20rOS6jN7Y3Ebq
6gtpi9/fRUox49cf+CiG2j5GkNsRQDH1/JY9nU43tNKQ0LBGsuPMS8BupoJjL6vu
7aQIvEKOmqgbsWQI2OZ2h+8i0F2DhxEuevo9q9VuUIWaTp0LEBtTwigKn/S4Be+c
hI1rBXN4Ldl7cy+WQp3BORR8Lotp7PuH1cDstf7u1pDlG5SD7MDAlyVGQbpcGP1m
i5lOLSeqxoHq45/YFvcQRFiR2ihIP05VD5oFiEGeyHK4Bn0uiShNOQfaT4MUJ9Ul
`protect END_PROTECTED
