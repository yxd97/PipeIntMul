`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNq8J95ULKSAQS9m5bFc5OYDBY74PNDDxSmKWanFoR+1ORFF5FTL9nkeLZqwRgE0
vPmHdLT9tj4o5ZItjMoK/7g+FavDwLOXMbparM3HxWaMmiO4eS9QGdgKc4ouXaeQ
qvBJhuR7nu0idhLWKk+aT1NmEreKRwvAgvU8sn4lxRGE4T0F4IGSWMTTUNHh7tZp
48KNERUNodLRIPraa7p/3GhNaKRVPYBWH4URm4H5tFPnjjvtPp/HAbOUbjAhlCs4
94Tf4zu7uIRRiLoSigHUdMGFEZJBLhdq7xuGGfh4xRWi+eWaq+BTu1ujMZeINQVf
`protect END_PROTECTED
