library verilog;
use verilog.vl_types.all;
entity PULLUP is
    port(
        O               : out    vl_logic
    );
end PULLUP;
