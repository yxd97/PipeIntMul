`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SzVGOAGcnmM5Ngal7jPPgjy4jAw2UlxTcgAK1yfclV8/e5dwqGnH199IskzzmEXp
AOOMllzfO4CZPAVTYl6c3kqRsbRBIfsG+qysjB2ThJIcssNIdV06dP4p+EuYfYwJ
eYXRE8hf+Frg0HmFEO3AtKYQcJFA/STjCr6+F0gNasxCvL5HrQUuwIiuPHPBJttx
5+B1gUv2Q0gWNBw5smPrgTmm9SvE0Zdwl6mojIARNi+nT1zyABvOR0XvCMPoBOTd
`protect END_PROTECTED
