`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JeGLgNvWbRftbS0o+57Q5ubJfJrdyvljgK8KlQhjjUSnw+cKmQd47qx1bn8kbdRb
wxZX3Z87T4Njp4ii9s8haCETanzlpoJjjCbXENpfxi4G4YxrX9liRrZt7aDgQ6X6
sgdMkCj5ODWlWg1bv2fspOhWbQ2jXjoeOif71xfJMhJA4X/zqpJqtm9L279euO1V
Jw2+eO+MOrRmpddZN6qNUzh3e/4pIaW196iO96SRxl1mWKMMqcLn8/aucNIsu3RM
9FK3jW8vEZFK57FArxRG/jXFphpGwusguXKoWZogpxgrzbGIqvfOWzAf8Utj6sQA
h4JSz0VQvtSd8miqygMVShIA8S6JwUNsvib4BOQBAe30b2CqAnMdYjIF48lpO+iz
3x2Tb4ES0mScG6gLwht6+YwQTSM5y4w9ygmhfG52uFuKBVl3NlxZyKS/Ww+COSBG
dZgFvIGPYXnrBj4sfV2tywfe6Dlr5u4kW4KTEiVCReZs5K4UVJbeizW5zQxKVVcD
64VitpRh/wIei7CEOt7NXwYvmxmNTAJSGXN2SjFBJ1UK1A9ZQVAPEc+bRG2OIASH
ovOHNnLMIqfS1HVh2/tdLX8TXmtymo35SkgSwHZ3mc0Os/SELsiqnjWswzKfxlJj
NnJkIAdrwEtvgGPD9fypzUYg9So856CuKhZ9OT+6580oJiqVwpR5eHsBWTnTERVr
S47uVTJu3YrVZul+ZwaTVYaurPOdwuyXTFMVDP68RFzmB31aVB9eicxXLymUQxTf
ck9TpDllD/lQJbVzcDaat0YPrq2AAnaJ0pIh8Pl0KUvH5iwocC1DD6V8LIi4S49O
ymXjyIxyb7WterBOMdBEmvm4Cr6sb28GKS2yTRT4ifFq7XuTS5Ubx4sHneWFeKHs
Y2i7O+HlvMOss5/ThAUFZqvsha2OwJIcDAGAf5knYR2rmBzs2oyigCZYC/z1KyM2
BAwGfFNKLj/DDSmkjQegf8vYBLr9FHnHAq6r0rFLwe+ZWa9B+EY4oBTtdakHycWo
AnJsLWWwfq/m0Hc32Gwku0UBzOlyOuAEe8Nj1ZjwesPU946SFvUZuMAvXgUvYAqO
7YXh48e/+X+WJ3GJ+z/S9JjxrXIoJdYEZNJ8AHXw2sq6NpsF8Pl0Dpcxsf+iEP9/
02878x/BFVmO+zhdmkdpAg+Ed4c34e7d1gZN4yWr4Pod0itdkQDrzzS/QViVPZ64
MJEBaEn7dISoJMvBbhBLAKtvnlEQqzvt6JSeFh/3AdjOUf1+r4mCgwDUnlk9sXLs
XgddbsUxCAjNMXaL/vlJSh+aFtkbKt9Rkr4GohsClGpi6EuVj/3k5YCywvXSd1Tc
siuIr8D1rXnKASF1VPNXguneUxS/KW+aziRc8r2A2X9LpLx8YgWSlqDNVt5ISZ7E
X3QzQB3SBSDooEo0ZI3Q1LfuL0FyqHTebSJvyJ3Id3igJU9vLmmeAaAfPrPW2MQH
i0JRaCfi5X8ut3zUt2KgyAq3GUEqEzGo82zrOEb0gHups6W0Ygxp0oxBIkCl5TBh
Se45uFxDu+U6Sn3K1gtdIJ99Kd6944uovN5LXxV/LPHSivNK8l4QamAi+6lGcRfT
phwj2JlwSTdutah2jusm6WJIqaxWwd3GRYDeJNRsPY4KwfunYa0kxia8LmyR2EAd
xpX8NiawYLPRU/jWCWociKm7gJ7UKspM63K3t3MPlFgYiZ50VlILUECUZUWWSP2M
NbM7G+eogYMZTeieccKqsDeRrzNp7NPQv3k8/tpYdR62r2nNWTxzDHNiSk9/76Bs
wADE0zCTE5Z6/94p75evcxOkfKhD2VNMmfbar3gWffv8SGwGqLt6Z3qX8vkxxfra
adrYM3vbefDacrEE5UVcZX4qeLW5g6ssFxzFta6upeNJWykzx1I8h0nas+LY1K8W
SUA/RQV3BTm8NtczlP2LwPud1uKUW0KaW9TAMoXQeQcOBdSIcdFUOimJITNkS2zB
o9TXwgGU1f+kiO6zdZ2K5gKG+NCf6YP6dy6MErlH89oV7UScu+bF+RzlXEvLlHP9
NLKw77TLVTaehDcR3mtF1UfTVwm2NXX0d52bgywvbWpa/sxdsGCXI/pHbceZ77ef
SN5FWfF4B7Wcu1ZYnGLHev8/Fs9xsiqmN8NPpbpjEXZW2Fg/TEsCIEFWsjKyYHq7
7AGeDWYziVNKF4hUtqu1Vmo7It5dM6prs8LEE2/RyN1XledRntELbvfXSAnT2asr
IQXlslyi2fn2GzbULp5Ri3i+EbP+07d5NV1qgLEVcutl8n0iPQ2fZqGifV0CTx7/
PesYo3k115ZfAWWUKcSu1EGfa+l+/zwvTj3koHeS3C5FX13qCxs+vbGaBgynj/s6
UCt13L7sp/VSMyYnQo57GtLlXZvDt6tOoxDgJozst1PNT69aXVm45CdLbfcyZ2n/
c+Xvph6Q8zlHN4isMmtvihsYAzauzwDCUbP6ILElG2DPDjnzxEWksTwoFaqXeVe3
xMnSYSetijy0zcM90hNI61vdvv+2yNz7GKCg/2H6tlVWbke8bLz2Wuo3OImAXg/I
Ue0HtYXG7HEq0HkiE3fjAhvOdQufA9DEH5sOZDs9bfb+vfsbUoKRR3km6qd+zneo
JhWGsOBks+wi3Wbi+O5I6gS6+W0RKdR1G3TYuhueQ/F+GpvibKwMs9XNZ0qY0gyT
d7T7L1Sx7sHAzT4nXvtqKqbHnRusuRxIr7jIFcn9s4/+e/1k0I9aBRpMRmvRHADo
jKq9L0itMWhrp/RO3adcx9Kak0uKwCi9lqGBgWi3+6bIsOI2j85SBXo5eyzRcNbe
TkXApAf01NQzIoJV2Je5VN300Izm5Lg0mfLrx3GPyHQ8IezMx+NI4yKlka456SUB
uXfx3qi/Ybu/el13laHY1oUNnzEgGEescwyfa+cFXL/46Co/oxVYjC4DAeu0irs6
ETQq9wvtzr9kpGa1NXgLYKiQCZY7r7eEC+bkBfubXEvUL1p6WyOXjofWJCiS0rAe
ZEUtkNR7ZvfqinZuZW1X07NzNLCYVJYTLBFfe+owmhrZlzxEnVkLoobcpILoGYRN
eaXffrjGw1SlMB9qpImWxl5L4N3NCEaoT+6rHIh73raGrVOpzTvxURHTLIaedOrX
SVnDZ2RbkNWuauqt9lPzgpkUmcH1vnWIPqi9jY4ET4pzWrkeNop4zNoPJzSNgIEX
hzVFgglbAPSoheGDTmBtPW7uGbQLZTxvd63CcX/EytxD6MGOb/96Zjat1IdlLq1p
IpdXCa5h9NUJI3z0Wxd6wA+BurNQJ1hF6VzMxLoLxnblk+0H1gqyVOyOmXEfK/KO
0GuMX6ktjBnhLoJ1fpfSPQmyDqbhveCOHDmyLVSgUcx5RmtqNRRHHtDbA2tovZFc
9PQzfkVgFO+zWYFGlVcXb9qCOCuk3UJeJcEt5Bd1p0/hz7VLAXzjt3DD3hOQBs32
lg9JmeL9mIaE4b2/Z1BVm5KqtsNM2JgUizxAjNQK1KniKTFSllh/i8tkdOkrPVC6
gXAKThvSJhLtcB6KkqxqfpuwUyOtEmWE6FZzQtTniTju/mlJvuvMaCjmfKPG5SG8
297Aq1eg+JkEXsclesZtt7fGnmJx2mG2vdiZ6KI9ROsAtIB/6/sSAPDX/vEifhzW
eWvxS7honI2uGxKKUPrRpB8qIFtI+51gIlAJ3op1SaaQVX4uEYE3w9RvJXYbTzpo
TJ3xeBhrKKSAodj+Mmpm9h9/t4uW+/BBISW6tAN1hrZqJqVKiNLNnL1JYLP0KGkX
dh/HToIYLPUP9WFCZkWuwq6JHtU5voOPa8cModB4nlyrhEJ78VzH9p/4PYADRLal
4mLj86/8DdlJ8T4QyGl8tVb+JTMXm+rsT+2d7NLOrUTFPI6DPyD8NZ1UBUXOORf/
7/TVGxvhqdYaCcS10/2XxdcGjBaNCOtqGSDxXvfqL+/FHG8Vc6aogdv1O3j9CD+X
1K83Sq3XOXm7/1MmBHf58Gq7Zyv+xaygGZsF5TqQDQU8JdWz1W4f4pTY7h1z9KB3
f5Tl7zTyhuY2gFttuSDX6T5LkcgutxItVSVgIpL2o2oosj1O0zvNNNJ4ow72jGQ/
l97cxaHcvy6xUuulHssLXJrgl1gI7EoRlV3rYbGcNMps0S1U07USHA6Gy4xGHSFf
jrlsSUBrzIjgfoIaFpZQh4F8CkUlcZl0F5Ca0nSJGtmkSUtXFNJdRk6EbVMftN6d
YzKx1V7xJ+rSQM8zAko+MTDs6QNUPXMtdd0u0tJ1+TcFuJCYiDEX42QxWF5G7ux+
qo+OCRhw/ssKfCSItyG8XPqmUdtAGxBzXuAoNsw907pzHps8mxRUPG9WL6dm0lm0
rn572q8C2gz/TxT7Ogx+ZHU9FtSnb+RKYDCb6pkVshjCIr/XN6yjUXTUuMAyrT6S
XSBTpnoAz8HYMt6kY/K2fE18BEREP9ufwHwbw4s+0DdbQdz0Q9WUC82ExfmaAdTc
G4DuTtvxYdW9VXXFRsDK+XkXkAHAVhW/HGUebrfW4e0ym4pvvMF+eSOoJb+nsoK0
9jdpxmw9R8aUX6xjASdSyaaLlBEcVHMYcfBXZSzVryNf5TrIuegRmIPnekrmUOww
D7sSFKTurGqCJtEDoLwIMOQgCty12RqOUi9G1MZ+AjH7pLz3JVlQZESlSwYXjcHz
dkAFc1eQwwkgcmMQ2dgRHfnm/boRiX724WaMRuddgLHSczfPAdbwrM6Ph8fkh9U7
wbWdyG1mpCSiMOsJI83h7i6vxUyOd1OVhZ9kiaS4YSJGzPr/ZtWnAVoBOj50Rf17
6UlCielzIr87RD4yLN3FnRKIbnK+8WXRdqqEeEHujHFZYxLKUWmkZf6J28PCDrip
UYClqLXJt0H3GgYjoG486znotkEkBRI0RGTYI5668t8PmQIFGwxVs7/+7B53ivcI
FHxa2OndjE3Yp6eg9Zkz2aYZOk+uJ7+rPxmeEOVZW3wMigMjHan0+qrAftnW9RQH
G9ykNsA2HNa5ZQvQ+GmuSKKnPjTYhDo/5ET/ir4j1RGzHDeSWAiwHBObgsBaIsOV
UmCHYUFqXN3OUrhulUADQEF1NSZmF2zwRfST5UfOjBmiZdl0JzKlViFhrjaC3uBv
eEtgpbILBHe/rlVqBK50GEyLqORtZXT+25DtLy6cYUSgf4LHag+87/fGGC68g2ls
hNkos1RO4x5EZMDj4sfKdio2Yn4xzNfculFoDgkRWB8n3ysCAx1x7CbzPl8CSPnK
4T8bC4Pnyyd4aTzWUSb8q3ro1a7SvQwuvhM3traqk7ewSe+sRK6liDTgdDBKAUDj
CYd4IVFju8YyBXcZdrs8Ud9SGMB1VHMChwjc5n/Su+KJdPaP0AOYY/1ySuRWBO5+
eeWFigq3hqxOoJ6CCXcQBmxvg4hlX32ltcD7YUNEWBpB3CHTbiMi38y4tCTNc+z2
T/H2oOIOsMlg1kr2Aa5QyUSUKI1Gs3xSmB2iH5D0qYOHrZun6Dc8lg5UpcMGbeR7
mgKKG9dWAQ7eVAzmm0w2M0xMlQ873gI5yQlk4N7ZfWyqo+GHyGu5glhX0oSkIOJ8
I9NvvwHwrfqlUScdowgV7HtIQNpDEOdeEqC4xl8toAD1i+UcI0c0twQN/mwwRmXe
52lkMUSrz1kzcNE7jQq+dD0TUxmPk70dt6VNEUz1raypHGS+AC/bURZ4UJUwdRFj
BgD7oiRl8uuQz/t7VO6P6E6Hi8W4ss5yNr95N2ucddkgNb5XIKXlgdWztLfnMecC
Fh7lXSwLe+bBHf0/11WsxKxyFT75f0/dzt/WuhrJf+4EbHRvuRcHhu/KzDUJiNT9
9izD/gdpqq63PXr+ekqVTBXlbjtVxk4TYP9VQcJawqClIB5iyvjlqsL4umYhGHfo
y2wZtC96FSFWcoS3xumUEc1NKE/ptu/7H0M+aWWB6Uij/FoPi0fNrAXAWubN2kh8
RDhWDvYZvo7vQmR9a2fBtK2wWtgOYJegSV46LzCebak3GCtuAb6Y4USCohk5qcz2
Dc6vLKQOm0xhBhiWRmwFoO+YBoPeUAixXC6jZNUqNAULZvVdh0Xs36mKzaR9MxRR
s1Vm4pbrtySD4e/u8x43LExBnGlWAWw+WHVGEOMKcb8sbbLE+7+maMD95kJHNiD9
FtcriZqi76jqJ47O1YhvyzRme5txqdC92peRhIs+B2/XGtfX+hz7UnHw/SL2X+K6
uXKwos4vrjtH0Ch2XEMwqfU9RTnu+5ht9W70QxNo1RZcLqV/MENCThOzJNXqsI3M
61evbiDywkwZ3nDlEU9d5Kim136cN2VxDK9rYeEm/wJoqiawcS3PdEGZV8bmXIKM
g/3BA0+UpZ7aov1gq3Cj0kA0OBYVwbZmBVzlNKqiqm1EqLFIYxYSoYc1n/adZWDQ
zJJ7Um65qjPsWclIGEf1/iw3b2GMXZGppLSsGOoJpvV9rPLPgIcV0mJp+G+NDqGA
+lg9slxQOJl6bI779vSWtI53w+we4VqXjJslzRBmSGknzd1xcPglzrUeYL5CvV4F
xPw2V0HYY2wg2lMvb7Hm954DXfzaxXm9mDpFfTCUJjW8uukl+YGZOuTdLrqNBXTH
VUvEF69DIqORlM6YFrAX5jY48toKYT+krXIr76cHoi3LRCW9838vHtkX2I+E3Umr
Qn4eOmdJKeYnYqWkqtpr8kG6WWbRcY5hApC9LfIdQ//h/O8JI7BT84lo0SIcBFoV
mQcV0hgupK6WuWuna6bKAqub9MZFa+AIo5BQ2+ylxtpPWG2OBYNblerH5tnoczJ5
+tSKNDMH58obYWwYgYTMm1dI9ehECH+F8HGHbsH1ROxEiXr8lnVUWmoQV8d+Jbgt
+86n9i7P0tU/2pdzR+VzHYpKIr6xGSVkTsPjynyIqX3xKX5gYTusWRGXBxw4W+qE
fUCLTB/zKTcNbZM8H43HT9jAJN15q4ODAVF+sutSadlNHBl4L3a/MVZs5QrPa44M
Lqp9W8wO1r2gqKJyW+xTdTSQ1PX1Kog3ek0YO5tKy51iQQv0NWrD1+x9XiUBEQ4g
D0XTjLf6vypmohrxwjuLzlqc4I3/Vd+djaQpRP8pVpnlXseZFNh6qcXyii8bQ3sd
10gVqJHfoP4/5IkT2J5tFEcnrLHYUibojJFi527e9Vjo69xYyxEfN53+S7rT0H59
gswTpvVw2R455y63ZQjw4pbTZAxUUcQcI8mVsNeLxa6vZUK7IdKlzkUqvbIEEXol
DRjKIMlaUV/yrqdvhSL7Y6yFMNjVU7BvUczSd5qtuEwGYorKcAIWTEUvyLnzhJmw
9ul5SA/rqxgTkoZoIxVU9twdCBw1lhVSJwdVDFyW3bmldsO+ovouvwAEy3IN/Rac
QDpbuP3XjI3kBIJnH1a67BwN3XoivAdzvU/YtBSLiO2ftyTVFFiq3CkuU4qt89Cz
K0WkrNiICR8/J3kEqsq+7Kuqm71MDWpwG8dE23pyDV/sIVU3yYkqNdwJJ9nW+JxV
zqqyQriEJWZyLFmfeGGuY0WpwZ2tr3cdIcjCAxZwWAQYTvfp3yxNw3yUzfm1U812
/XJR9X6/O2WdA6TjnIQ/KvD8V8lmGUDPTt2TEIho9jxAUlC7b8ecglGNTzNG4IDk
1BAQiHJglDbIa05Bw6nKLBxb/afJibzNUFRPgEIps7tXv8J0W/pdbEkrTdmKDhsE
TS+4f4J1Vj7w4wyI4FS6ae3cFi/E/U7vWsMkAuYL165IL3TOtw/bD4LdVVPKCrjg
51BhaSY1+FRQdJ7XM0tRFAl/Xh7McOLxOj+DGD5HYM7EciSad9AYPdZj9+3ZwOUd
PNWAUVFbzQfuZO8CYpjwhmCcvGZUluHp5x6ltH/MWoQi/VVDFOYMKUZ5tzMxWuwr
vQaZGYa/VZoDWtlNFPW4pVIT/YtauxO+AwThuNTD2hFS6GOxGwQNUm5sL8N3GCux
jLEmAJqh3IHgkxLMSed6U8ffoozfPh6TAorcrQm9qOShXu5yMBmhSYhAk4GafkFn
PCEpyVcJzkt8UdBijgQ6R06WbCckfavE4bcevdheo46vwaFUT8y0ilKqp6JrgRTZ
HN4XaiI1RW3fJokC4lCow7AHYWEoKvur+j4Bl/AzSUJs7MA9kATvYF39aus7UPEq
QXUj3yaaFbGZy9Xlt4O3k0ZYeTMabsNZwQ4BlbthOOz2JiZ3QN9S87O6MPh2sEfX
65NNnWec8xfqg3kyOx54PhVYHRB4wHF85MMTbfcNJQx/HOjbbDOICWg6MG1adXkm
IKJmQR/xCXYBc9ngxHZBpDbMCiNsC/ecR0BgFLuqdx8YUhZzDj0PVfF7OIHw0Elk
HyyzGWIhBhxbYW1fCGPKh2Zs78wG/rc0lrgyFNtI8hcvPiyB6HcFOaQPC4oH8NWl
u9sveZ/fpWqxYccozrynvuDBzLMekScnY+kMaBI2Qf8+HIq4kkXlH01lbJ+k2bYh
jB9pmW57ew0ydAACvkUFu1YG/F8hRiyROpUSBnQqcHSYB6mPapFGUoFqs+7QVkRa
+jXH/wPxqGbERDFKnRycHdHV9zehan7iStE+UoTR6TOdecZCrmZdJDnCAbe4GotT
t6wxZUZ+ttaOIkqCOTutVs3oBkH0yTMe/r8m9F9MAPUp3TROCfqfO/kStwcWgBue
L7Jann8wxBXlSF6gsX4ZAQmZ8xCM6Q51AULsLnUAzokLZwNeqzW8/ORKVma3uKYW
ozJxJd2M46m/GPypqyxfXg5NUxY0IkYr/zy0kfEIFwglJqVPpIrSTRoA/I4IX0cY
d6SRHSxXcVKE1FW127tV26tptffaGdcO2UbX/v2+DHHZf5ajPQJyekYLtmucx52Y
s2m9hLoBYzRGXDVXUKeQCePNFqPhUX9hEk6uGHvbO+RY/zGnnyfjvOL438YXkHOi
jAFfDKOgRZvA3q54//CwmjidFkLS3ZB8r4mWeFI4VD9hApF3sQW7HmPBkTSPlczA
l75x1uxckdLzbJHlEPXwHoXUW4ngMOZVTx5wm1cgUhFtKpDrzmjD9nmzY/EorGF9
UZGrd57UCakDiyF2b07n8k5hWDVbOb2bewtGuEZjGD1FBbBCxpqXjFk6r2RccHqo
T3Lw4kOVWspUGindx47EFRNpnpgvym4Qi0cxyph8nYNma0XSFvwdu+x+xFA4ayo0
0oqtrck4yx4yFSAe/vEDfgpCF15yPfq6VLKGNoCJG7D1OSBAvjXMHqVFKG7zewZG
G8/QDfPGakwp3DwSwuwRXRi9zpu4U+p25t5kcs7gLp2PYmnMXc0E/YXApuG/YbcO
UPt8OtVUb762/c4PB/d7hNCmgF7Pz+yNQYLj0ZltztxISVvCh2O5wm4qvNf6LddE
GkaeEZCTQLYedsQm4P4In6bHVJe+FsjksWR9ug2x/FMBwhd74+KwryPa8Wsd5QBB
dX6BxGdDDzPLBj0pDzGrboXLFQLx1s3c73EksnsKe0zJY/+zrgPynmTp1+Ijv+I5
Dftcgt8V6Aqt6NE38Wnqx4Bu+oj7HFBXypjmy+wc5RboQlzaRBajk5P0i7Ing7/d
HT5wDiS6lrpdLgHuhITYox/Ypgy/I47Zer8ClsjytzLrfXxKkJD+DXX738SLrTe+
rHRwPvt/gsS4yVkIY6+MgEO6UhbBXijWFsaSh683c1PGNY+QEit9n1u6YxUJB6sf
YMFws+MD9p77oTJ6iKItDZeIjIcQMHet1m5x11P5U/VmHyIiTlzncrJ0r5JHf1BB
uZhtB1ed8cuClBurPEtBML4qE3720YoS8rFpYrMU6bKgR4Xg+jxGXEFx0G/m2Cyr
DhjKE/AImo8Sr7hhULcDh4ygbZDlS8fXt8IbRbFeieH5QlpOh02uaGI+dNlkBSo9
R90TyvCttLVa2PoROlgfV9RbVPMiqP/IGJO8c7A4V6QL6Dsb3T8rNSglcIigI2ct
6gfyrR0cuOSwVCBtfbq6OYEXoxuaVcdA4zTlg8p3zTMyAJTKZI+k3wuxDaBFGs3p
IjfRr4Tg6kIjdMy9hN9e6CO/f3HIwzaZYq6eqSznpumhbDtohbqgPAune3tvrOMN
IS1Hs6pca1nYAKjoSls2KCgPEThb+JOYlsPgKMXE9orcstc7NcYUx3u6GUBXslbh
l4/J3d5Ih31+iNfDsrVg/kHZ7su5Ltoc1L35Z5aQY7PgjfEHE5S92IzA4T/Nxuah
52QyrgHrZEsg+XkmJfnOio+ogYqoj5GlqttRV5oeUPP+aKD5+gmgB6/M8CHifuNl
y5MPbOUbgc0wFfplVX5agsISCxnRDw3OcwGtk8ofkTmNH7ch61y5dq6huuyiLs3D
nlzGDBf245kHIMF6hpcmTfKuxBLQJU7FMQz13X43GjGpz2MZgJ3fvfwhvlCo2wdL
QZ4b2x7bvarPGcb2jS76YIYg/DjsxDMOw7eULFLOKG+L4I3tLdmeUANRdtwEqaex
M9fNcATLSE1pw88Dd+tUBrYVOv2aqtQ2QB9BC83YeDNGqm15oWSsIHgxo5Man8qv
0B2QP7qsyUXepIcqeIBpHacpaHqu+8iaRuJxN00rfl03tvP/GiSgHs7oPb5biXSa
tg9o0UCnBql4dPjTCDoH6onNxAJ1wdAjrnL/wN9ODq4hgxbrS39TxEzZKeZJAZtD
m9lA5blwIUWr9AlCJHGO18lb0lMdz3z4ndGpsbBzAvAjJVZqL/oM3Exq3fiDPVqU
4qKdmho7GvEzG7dnSGnkTy+1XlXgqJQfL0OiFbwITR0hC77bSk0HrAi0IAEALYrd
mUbZLNwOOerroIQYLNzhJhT9CpsHWxz+oJ/Evprom7LD4fqY05K7wulHO5BHzuIE
qFwEq6We6jgNKjqSvmHzkkDfowCj4WADKN8lk+jMiq6j4k9Uds0V7MQmRyizfCIz
dbyrtN9ZiB6iULG531PwX4NtWTnat4XEwLiIcRcv3M+PiaLpV3x+z5pGKLrx0ehA
GkgHuhyaMuaZFNkbNoCPKVyA32ES5Cb4xKe3XvkOi6Xl6GcgjgFD7c6LGIrK8ckI
BUI/ZHnoiT7dksm4ivsC3e2L9jeThFz36GUMU/wydEhzV/OL1A/s/JyJvbpgTssV
cAkTQETHARq3Zjw/nEKTB6YmNIxKNFL8+TEkCie22LYY9iVZg+TzRw1DQhgXzmyc
KRUK4zAanZf43GH4LTDKO3lGw4AG+uDicZQrSyUoiIDzjwFTFSawLcmwLYZRPhvQ
8qZlacMbkwFeDRa4XyabU51oQapY0Op6Wp/hTObXwZUzT7iW3phcktusHo1wwni2
QWgauCtO10WXxJVRnAoF39gEmsIb/hb1Axu4INGINCF1vSRCYij3m/GUIrL5t1pn
Evu7wNDr47SpsvGqIpWPAlntka/biOrHEfrnCm/jkAgsYuEbk+XRFDxKGyJVRWCT
Nmd0r6kOsXmygHDPBuPgplGRQkg4IJJM8sZh1011dOOs+ZCyRJ2KZc989sD9pQyq
nZghlI/KnNXJ/4wv6llxVQ30YPKeqYVZlvvBzddlqnJyP2oAKTYNXkgtiQ83dBX+
KQqfMP2cTWKdK5tArNHelHowllYNqCD7IMIz1nw40frdWXpuQAPIW5pVz1AIY4N6
sdBVL6YhBssXtsIQZPqz+bS/CpMGvxjbLsS7ueDXCufEPTZsnigbzRmUMsqHY01N
qMmleVENum+ergnTKvnFXShudJHPCVDYXaB865v3uKjJ/tE8NRJ9mGsnAOwUNK5k
Ob00C56EWTCDoxv/NFzU6ngZQ07VMKDDWFhBDCPbE0rRYrRJgIRINGc/hX8QQTNb
uKpS6gIE9iy8U4s52iIm+KMSVwNu5JQrMtR6wineH+612CdpsOuYvlgjbSZ7TC7d
ZT5GUNeajLt1iiGwVn9CP6pY2PB2VbPw5ZHvFc1UHH1N9rIzCEN4aWmtmNt2eRxB
4ZX0q4ZlZHhNzjxGUpOq7y4DEl1WsJv0UaXWMqmdFuRbJkI6vmvwVvs+n4JF9M5C
6OuzCY7WG341FBLaUkwLC7UAGYGvQHDCwuIUqD1EOTTKZcva1LxJOY9dbmw4b3mj
NSrn0ZDDu8kCkJSWULOl53udf7Wfmboiu1TQAN/w/nmHrukncwZWYWJ1F23AhX/+
AFJThq9MAGfQ56mQIwU6g3PYPp7GdrphdAesHO14nqnt91cWjKI5O9edHjpC8pqD
SbpV28YB348WaKSuZ8tGfLkCfJ+PqohhAMV5b5PqHtNFo6/6oh7zToGAnQLc0tzQ
bdWqD24lYIXnpqQF2VCOmaHKh6jG0gbc9OsXZnguCucnoK80dIFJBakea88cV+Dg
Hs4hv5UHw+hDcsau9HfeB3ttBRTF6APDLgCTA92sdNJqEPIhV41UITMeg/96nfXH
ngSnz0opgYJznDChJ157s88Enkvt9lrcEOXadXvB92coBa/tmdi1oCtlZRoyekDs
6HSeTUKgD80/WedD8cLQvtojQH3nqp1K4PXIHELwKiXffatm/1dnQQbIKDjm1fLq
HmLAOh1+Fnzy0p5GlnnzuNg6U2DT17UD5xUkRvAz0jiOBha8W78L3aLhflL8606U
I3FmI4LE+ecXunevB0RnkBugignXYtlVrGOV/iZZELd6koY+5Rl2ye7MF9kibeLq
`protect END_PROTECTED
