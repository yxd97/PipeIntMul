`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2k98XrWLt5haPjfUFeYZef7JcH3PRGsj8xdfGDqdRk1e1gyNQjfyDppqcub+Kh1P
5usdA+/I4Tet2IgE4hqo9fo5PWBhOAqEvJtRYpuU7euv/uFr/9DH9wZyp4jv4abk
s+CBzXzhpuNDbGQOtdikPzOhVgbYLLGWOmu2QaRfA4TIhgzXx2ss7dIvrMfu2ys6
RFKtyxJV4uCuBJ9caDPPIOG1k3nAJv267m2MvjhF2BW1u50KBbJYp8ge247VW4vm
b/mcjKlZXFjDFTKifBj/xORV4WvcV8YhFFyreI6txUJMV2Z5xQRQI2/+ljgeDYF1
2NdkNHp5CBy4sALHDQWBaGtvn8Npqm/BWJcIUYBGd2/oyX1/rOIl5HrFUV2ay2jS
+avHCyvLP9BVxj+RTMCEHnZmSUoedi6I3HYng71Qa6o=
`protect END_PROTECTED
