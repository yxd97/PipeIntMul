`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVJ19ZXRdefNMKwMc9CmF1JlyC6kMm+nVe9ZmLm/dBV4eENKO2Ktf7ZCBvmwi1lb
iQQGbtUbzbMFr3PHliJ4FOplUMJTOWGBAnb5xYR+21Ia8Z2U+h/RI7iPY5mmOF+h
bGx7BJmNAS0hfE2AU+ncvMQHYO3fb8KOvvh7jS8Ct4lp+1mk1GDs/b0hhtUVoY1V
rmZAhMRmH26DjVnOj1IYzClYfgI3GcFDi71wAuHCUmqDPqDoXQb4fWiWS6g2IM1Z
DdAHBRykifoC94yxPsUQQt17wQ2WXl8FPTJHli7l2IVRg7uoa/3hkFe2GdIb0C8L
Gu0Ctk/VHs2uYOCe0sMZgQ==
`protect END_PROTECTED
