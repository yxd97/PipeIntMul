`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ACtj8ReFLrRE7BO/zpQBaMJHg69arNRqUHEoY4/439nNC7vRgD1Eh5evdigruhhU
OwX1U9OUz/QlUiUHHtMbbIuH/4ULb/AFzz/8nWXo6R4fnBJcAohneBD3jyKRna2Z
XAt0DzkRUbkb14GbwXGjph8cXW64oFNtFL1H90Fb+a4R+ZsT48s+KV3atIeRo72I
XIXQmkfW1LNYxOkm+osszQ/Gl7KQXW2yEf+Nw9avhp8HQ/FSmLfzKuCYsmvG1L3a
`protect END_PROTECTED
