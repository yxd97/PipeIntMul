`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3o5Q6ADTrj6vpzOudUH4IWMJbWyTxjFse92UtpIP9Pk1W7gBkrk2qmPiZ+Iv+Gu
R2hl2qf/AIPm3+QcTqLdqqSxzefJuH+KB+QP3OV4YhwWEgIytHUA0vfkJ7hbb4N1
VKZUh1TqfN4yzNe76GjXK1B5VkgrX8SZjna2ZPEmTegh7jKIQ+6LxwvvvzKSw6fX
20LNL6v3h0haNvrAy8SVNUaR3Mw4dcglSDtikxfkCXugIlDEqnxdgc/pq/gZzXBC
cBHUCgtDCkYN3+HFWeQCCpBQ0b4sWE1DUb7GXFaGJRAHyoSBr9a2Bly9fLO+E2BF
aRhxFjtKe07PS2ZhpRz9h74wmOyEv03FFMeiVHQp65tdraY6KpQi18CNjXauPfJw
AivMoE8wSzPOZhx0rD+xIUcngdPgpZnHyxSCGpRtvItWdxTtaKR+M8vwg2NJGxlN
7+NIxLJcMIdFkDKV14rjxxdtqvDeE88ZMMWu0HC8F2JRNDMJPLryoQe6Holyte9E
YorGrL89xAOzY7zIbTr5XQtRw5RjE/g0t7PunQVfrziMEqhab4xfDVq72js8vy0x
wqRSCW36fBOx+cSAPGEwHEPbt3NY3qqMamr6XzU9Lmg=
`protect END_PROTECTED
