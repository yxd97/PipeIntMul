`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ijLaUhReyIMfeD5hC8hR93LPSfwYXhJRXdQui7AlozorAADi98RpYN4dbJHviNl6
u9YhCa555RXImRmZEjyex0yGpygmzauWsYpxkQZ7z4IAUVCKAaIsgvXN3sMrXeuA
KNw0+Om1ZpQoqWP1Ho5DCLsn9yLUb4gdd9So/iK644riyt1aojucDy/4Q/MDwp9T
CfwmMJ7Svu9ZcnOnTnak3cnonnbnxqgyaFFUsZR5BBk9Y8nmfHOR0DB7Ok/AF4MF
zKaxKMo2s8byHEammrdp3SCKREmDII0TVn1y07A+5UpVzh0OkIZlDuQh3s0WXKsW
6/5vK4MsD4lEhxabysCbvjkZmgYdm8GXocRutrowBMZBQVTxzIjaxE+DsNSTL9Mq
PAwHPUJI5XW6CWF0SA8eNIA36EB9iXYoCOfLIGEM3oFtFD5qjpRX/krydvvVzWoD
MJvUIwu2RZ8B/cQOx7TOF6rNOHlN2LH3yoYrKcJDSujTfLW0BHdH4OxzzlfIhkaE
7eIWEPRufHgDv+6smQpRX+wMPmN4REQdN/u3/bQYXJ6qrQ8gmO7gRWmvjKMXo6Fk
GF+EkhUeNMH8PtcjZG6vhbQiymAPxLXoBF7Eu7LJ+DHG633za+iUGXTlzfaCAMEe
toDSrXSxgSGxLMOaXak4ahha7hzm33bto/KHaxaaE6FceYlytgdqlwDADjOJ8VAv
C/Scw+pQUfTldXkyeWObmrsCDoR9K8LT2U9ILxvqoOxnF7diXVcl51te6+j7Pn8Y
Dqw5UhJSXcnOVUV/MSiM5+BxhX9+NP1g2Jb0/Y9ySei71mVSPL+/2Legk519Cmr7
nmwmXyZ8hK8t8ywAaz4VVYuv/dt3ezQ5J931W+6YtZYNDkiNUpb8kbT4dww6KH1S
3lMvJ6F40dbBv/OYGxaWz5MnkwCOt4pkCXVWeM736ErbFSke6ZDSFlCKPlFtbfzn
ULBAwaeMCFTOSH7aZi2cp1CSpGFdk4vsIpQBHgJMhaNddEafn8hYUT2hv6ZK3q0k
yKkqf4jBBR63xWN6o0TGvkUA+tX/bt2E3nF8TpKghn9ptAXpMzcNbPxYQr61bz0V
NvEh6KH9viS6yGOj+hbw11NHQTYys3e3XvWn7zB/RYmVPFK279+/Tu1jdRFrFlK9
HpkNGeBFAxv+ukIPWyebLVydyE/P+chKkfGhny23FfwKqvXwdHPYtdYzkb3ZJM78
qTa5wefUr46pccnF+zi5ldBxqxmPE91HmVm+FI8iMB0M1X3WcDRaGwTXv1R1gFs3
SvQW62K0978XQJg9Oar7h8oLtKdzUove+1UthKPWRoWge42yv/ZdNMj0UxUnSc+y
hG/V04OfJ/4LbeEdSpIfHd9ixjolCigP+HJpk4wklOpG3iAtYLrlS06Hukl2KzN+
YSshb2AoiVIfNaNP1aV3nimlfMoFi9e3wdUjGO5VOob6fdT2meikicWt+aH3Fpsa
8DOpTvPO8wnUHeXU7tXcMTszXBIk7a6BTQwojlOVjMF9aQqWLmoGESFpCM/6JPWR
ft2WBPot6YxCQs52fY2o7ixScmNRWsKdpK+HXgH1eD/ARNcE+7TYeGeo21UZYBo/
CC9vFMiCNAdEpvmk4HK9KT4eh3j/4ZVz1jDuEPVB9L4MG4uNYF+WDupMIgp4qst9
dj8T0OwhBhQQDOsZgKW4su70FtHH5MbLdSmtvi/qwWn28kyAoBdIEzTYCPvmCjqp
IK5a3OrpLmRiwSi4/4Po+uf+uY9Q5A6N6u8+KmhFeKFipSwmKmXg9hhNr915eJsb
Dpq3aGpP/SpnxgCGF5p0mzxkJ6YYVS/hKmWCP3RCoS6tY7i0fT5fJ/uwN9CH+OW3
8lRyTd0tCycrAKRzigJU4X1acAKD+81oHESwFn8mjV4BXhPIp6xWXBYNTsXtDwuw
UH8qzsa5wqtVIV0x2wXhStaBZtX6XzOgBsFBoTJD7s3gFIKQbo5XuhfiFdEJuL+b
E3Ap18ene1hpiQT6TeXeLq4B1l5p+pIwt60jgFtgR8C+3i+AWt0Vs8b6Rve1rBN9
9QVkjFeoh55mjaRtqmSVog==
`protect END_PROTECTED
