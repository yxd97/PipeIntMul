`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64+cIFzH5RNAaKS4RopDP5fiIh3uYvEgWanQoV/Ojc7YOhHZQDXwHih5TTZDmWnh
iSsE1kSsLyNGTq+5HBdXyi5x4moUh6L/T1cTCXeEAhRtiFMwQzWHjd0FMd8wpoGM
slvaejAxW7NbohNX9WpF/cNRET33h6t1An8QExdkHfOBHiyy7LKqKCmRqli9Zz8L
UP4eSyluJvUKD1SY0e8Ku1RpwYVXXp/Z9ogFut88asxzyK2Qz0z3m/kaQiFq2jHv
zV7W0IZ983PldlfeWDn9cw==
`protect END_PROTECTED
