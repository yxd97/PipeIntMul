`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EPxxQ/RRSU9VbaDbX5B2QkdudJY8HasImfeXK1CT75Js7SR/YEPyP1wUUpUXgL1s
pYTI906GH7AVgeMeS41FDd88OQG7OWcTVbf51/bqJTEJHiCkgto5BFwCYd30dSzG
ZLdidpvwlTBAFVObTAeSzjWmfq4P5/4VrZZp36pd1ufgAOVRu4h5GivIkXJlxf78
/mh1eNtgebFm6bblma/njQoWXrYtBeS9odLTdVDvx7qeXbICqEX7Oao89RJ9dPrg
4An3yQX2HXfwBjZefwRqKDOyBKxgOlEsopGDu4w+1VQzP05jcRGYx8uM0vKM2x3k
VuKw4bxWp85dubpoUZFdbnfAZoDtt3vH6c8OOSjERR3Wumq/zihZZEm2vLDVIedX
zcXIccJURbtucTYcC5M8NB6cWJmAk8+8hmGzepO4cLFY4zMoaig1scALcPlyMR1P
R6MVU9eFeu5CR/ekwAgmtiaqENvzY8JOkuWvHiYjbE2U4E9f6kAojCRcLhnW50yD
cXOSuwSsapENEdVsNHf0Z/iaP0vI0o5bqQJ+orPt4UtiFZo/EG8cFujvKMU01raI
wV3gLN/+tNr22urTNET5qg8T5ai4Ir40aXGqBGaGpaUMu8+lOheS6tqSJxd10M92
Z9QI58+IfePEDog5MtB9NUK4kM/iFXhenpcngsUa6pUStlXZHLQkMYf5BfZ0h+E9
XQUJT1g80T8wFtn/Ibzp8j7YPs4VWH5QkjoQWEChrW1JssHATdbYgKsLaD2pbWkl
4X0BYi7C3chsSk8UXi8ocdBXsGfExaRYRJ+Z5n5UoCS/Bel2HLILaWaN9KDj08fF
VaNnec4i7laUQdHQs/RL9XEzTzLnxVbYS0ma3vZGtlL9oliGVw2Sks9fRu0WghH+
Oybh8luJ4BmXPnMFTroT22YTB8MAumUCoOo8h4BWhCXSe2PBogytpQJPcRRdeKqQ
ur2nAUCzaDZDpJALVElMWh7fghU1IqNQWKat9wn+FTbqz0NBuW9+xXyq9z5VpaZM
7uAAsI/KaySjHGU1YGKoL59WO0tbaJ7UyyWS112pBOuBIiB7Uoo+WbAaU2JU95vI
zfVyOJPh9xqjb4pW7DnqE7ffXtYjKcZdeMuqonUPejrT5BHpBvoE+VeUaJTYttlR
PpI2IFw1Vex5aqVrkkVKNKAlIZFXCQYwfluX/k1OKGMCR//kpC6QSzm2ka3365ca
T1kuN7pL7VKvEq7yJPkCPWP7tqWgQg7HeFgEb1qoK5UJxVAbVIyC9Fh4wxvfvj/N
4TqrwttConk5x/5GQPe7tuEGFSv4FKJPNcfwhXUUuo2BX24gYdMpoL8e7kV+cTtK
LdV0QgN1I+aX8IkBSC5qs+5dK2jFxL34Q9g10uG1ocOiB8+lCEOISRGpYLsQ1zC0
ootiQ6U5vHU4FrQ9rMkdISWWPEirJF2KAmyo/YRT5/mlnhjUuzCUur1Ay9l2B9Q4
Qo6Ifj+yyUQlca1PfnpSdbIYigP64E3iJowRCVgwQVl+s7AkLJiGPJceX6KDfdAP
4YgHCODASYOtsFvfufm0Im+etL6grlo3UNdgNSoRaG9wa1M96nC+EDYxWO8//Yj8
v4E1YndDvVbZ6WLRE9vOecxa3JmOQsoXhzzlGVLSDkN2W9VDMwjwXAu9LqdiHPEP
kcOQoaD33jXK9m/GqMEgxGObJa8JzJ7yhJkGCr06g4rX5i0SrgVYBjFVNG8CavdX
fTZTDUx1VNnCyDkgtn4btuvfZ3oVWNbelYprsCZTMOiS1b90W6eKJv8A6DDELvE3
+J1V6KlKsPsq4/j96H9HpqIRFT0MEL4yFAXT3BArnEvkNB0TKGDuNDUL//qtuOfc
c+vHpvaHrrFMTpRfegg5UuHKThcxO7ziZVYakyVtME11S+5jw5DEH5GNawFkJ3xM
JCDNbQc4pTPsf7lcLLDCRanLAUVIRfrQVsz1ySlO0m7kytrJfpKDdhNq/MW3UQZ3
lUznDQ/k515CD46bAAXv3+3zFjxg/KMzLL+RN0yWlD7vYfGy4KPibHD75Mlft0av
UqZZBu2ay0mefiu35fJLSFKeWasHP8FBMk7TLc8J2V2FTdo0vu9e/HZd4udkoFW7
UuJBzN5I1mSYmBqJkLU2XsX41hzGuAH5hRIu9nQhi9gAdbTLNwxXkmsgYBjHNk1O
QgFwPBJclhXWLovM+Ro2xgQtN1Z6p7So6uoapf+vyV9pknNfkowJDFCRVS3LYRYz
sJlGrKE5j9J6yNjA/XgJYVzuBnvcaoxV/3LEn4h+HFqGWefYdHvbKfQfXwQfYoqB
43X+iyjv7mRT2kEBL3rqauwX/SW5VwwWL61x+NJ9alXcyvr5rCb7Qfzkr03s4ry3
ykyZ+tu3bojEeR2J8XAWFmr0g5tyO46oJM/OWyh+uAnKHRBNm+yRmCC0yi/iQPDQ
5HcbWwI9oAnNkja5MS0yGIVaHk5lqzq+qYcsnMs41SnU+QkeT6Pq+KnDpGeBYt5c
q1hACyn/vIRJmKHoaEZf/ct0uV6IRWrpzZJowIfikGt+qu7pRlL8so++KWdYBmDh
u6cLNXiRJYLdOFnKF2VdxPVZirRmmvft9PJdtNSBRypEw5ns2aMQE83b/KXlfUpA
0TaXGn74wiPFG6vDDAIDWwXi4sl/u0l/HqV80/ytVdOFyqXqG0z9jUqXtdJCAMed
TbtwSLeBLzlVhA/FwlYACnsPiwsMoNrRdl56R84o90GD16TX8S1pl+1LMAhewm+E
n1rInTLdDOa32lGKGctmp5VGrKTpZnCjzShKMeXK6eajQ1rljVbAtDTMkGZQ6khr
y3gFqKr/LgWlSGntBiCKzwbyWGnVprMjocVdnmOycjyh7l1uFOWSa0GrDs7YJcsO
Ox2joaTfti9F40nXi9GBZ9dUNvqEKnUMS4SZfxYY6IDarLKJ/mTMFObpoawyD6nX
bkTlocOsUhPkquLiOn3Ykdk18Jvu/WlfmccSvb2y6zozdCIajPJNCeC1n1CDMhdh
8PgeRE9LxVB3T+6Cbm6TQQs8bRSKfB5q2sPrfX0tqcD7jHkS5askrahyCb3HoJql
6xmkylpZFvLngIO3y79kVi+zlgocaplMezKlXngMz2gv6mWWhyMT8gvkFeUwcnvs
16t3HepLS6GoCUsBLET78x1j8WCjTeAyxqleyVmtyRxMK1328fFHKgzkro6HTZp4
APmpEmk4huaN5S60MGY5wdlOHgRUZ9S3RUsqiwvKJclKbHtkpvIWbMmOVNyWXQpF
mvoHNOAW3xrEOnkKanUUc3FfDcSiz6LI+VA/50YmWNnP0k5oHxb6uIXwoY8UIeBE
7DJpFljd6h2Rgy06ihrqvmJEPFp3XLDNKkYiv5LOKu5eJbI3Bk8+mUc4As8roI1C
npkn81hP5dpNWKMULN3y42opuG3L7MDuw07OAMbaaBBWRtrXcnWZ6aAOOVKfNIl/
v0ZpQq5s5uaqRjshuWLFDzo8L4qNiFaHdiy2ZOv4ugbkth2nYgFLXl5sNbCQC9w7
DpJZ6uqbLfPJ+fonnWPAWTdssHdjDrmFqDx/drzqWJSbhwRyV79V7wWMrbZ4ZdnR
8rC0WZgpAuafA5G1AiLKeDqCqu/gkf1XaqIFs1kGVkENjAURisvJPqyfKDVsNXgL
S0rRBBIOyrt0EHwRhShqMhwjEoMHbhGKBGlUPBGJT977NYWRWc4aaE3fuwUdFj/Q
U92KYuwsDEc6D+8JOHJ3DCUnpYItDURf+VDfVFl9lhxV2LhlgOYZtzTvi4eVSTml
q/+ihLKgBbRTx1o+5ORICuVUZNG371n5pQ6pPDqKMaqOob/mYTbw/bKyZr7RAC4A
ZQTbGQGsskTPA7auuAw4o4uazDgwqm6aYuepYfmWdsZy0z5zc/hA6qKr1LZoetnD
qbDmSODowvP7Jnai/leFHlK+293tuM4KOewS7vPYH8BPoVn6+jG6iu7+nlglkGY+
SHxKVvVdcXiEfivABrzdFG0Q0pfUbE6UkZCNjgaprLy7y6tlpUmSGEw84rUgQP5Y
d/8ajFuqKDh4BoZAn/R2crsrEbd048fshDvySUlHLL5GPj8kuhd4iq3NAhleVKYX
8eQx9toqHetwLCIsP03lnVACAhWdGzpkL4ieqpkwEEcEHTuOyA4Xpikc0zpFVs+r
tgqH0LINtfe8mD8gZIEwq06R9VK+uvBOWeKDajDd1PF6igaN2W3e8TMwhpun1d+6
6X0rUlnEDtFoTmk9MMn8MnCbI9ikxlLg5o/XO995BJTI0uG4INRn5iOEhAlhnTjo
16gVp6+IAxk5PeR7pFGULKotVsw0ITeuaazZdZxb0rhy67mKIGLwmeXlDrK34QST
MlJeS+aR6KCuct8qImVLeTRJXJzHMK9s0oSploSUjBbjkF+PGDQZMdAi+NNo9rpl
OwjxHA4nO04rJ2B1M11i1B1EWgM7A/+0lJFZrqVsvSwfYX5YZFJnWj3fQL/r+AzS
ADCN49AqbU6WawgNErRtTVedh1T0AMRjPhvLP4zZvw3sMnNxyAKfYbYWereQQIxY
vaXU2T4PSXjKDgi8p3g6x1Jc+uSfd8Un5OQ2yUFf3yQO5mCzZvRAPqz1ftk640wE
f3P4fbJNFHcvkbBWskG8Nh8ajNHpXc92qHuUHe3bJnydF+Fs9MKmBn4w5IeSzebq
c3PRjpv8PVHWsU2mF0N/VqyKHV0JzPFOptfN1RekmpPmlfhvrYYKdUK3IKCgbWI3
otAp3qzos/wYwSbKSQAtneeeGHzTxQW+iMXaXrU5JwTL+flCGhHUlYPiIoAHN/oU
EXVsqw/aqChOKgSdIcIE6S70OizXZgnYEzVZM/BcI9k9fTXuMsMe04WdhJ/qGyGV
4J89zcjrevfyfuwKoTYYFPR0hHjjKRjEX3F6pHn8aO8+qOWOtmNya0egq/C/1LSW
wu5qearZFgnppqJ6MaeUe48pxsPVIDEGcPBBsIkqS/3SHqjx+YST6OZIKlmb0zly
/Kkrpox3WCWvPVt6R2nvEGUYr6AuGKYO/vTeHmaTsPbw7iLgqSNnQFDuj/pc3ZmY
/cu3m4kmfAMi5sLhRMPnZSSOveNpiNg68e6HIAkQcfOFwZY1EPQUkLh6B+Bxc+ZW
kqdv2Ea0tSmlFom7SU08JOneTiciCtaohMw0ZkJGMJzm+WjZFDzDZ1T9WOsymd/x
QkWlDLxgot3E1oeOhu0PfnPjaAG9Hf6BaQaEiL/1iaUuNm4dr5YoAtTUhM9QWn8M
81uZpC8KNKV1LwszX/PgMyIyftcZC64W5S6daAm2+KMwxo8QgDcfGEqk6I+WYc0v
5abRaR4cRhFPpTOGO3fAHZ2/Sxh4c3fetv4opwxCO1/B2zH8rOprpFz4UqyqjELr
zIyxvsaBlAcLeFbgk0EqB+RsfLBKxiu4Hkh0mzLhfZIYkllDq5nMIaxGOeUQEinZ
j4wPiyEH1SYmP9TstY/Vxiu4fjCiE3fClx+FiPAsZEER1+xyuiFF4zJP13KaKXYR
srXbomR8xHfn+eQIE82ZgkOdSAV7gmlFOqoFJRF4f/y3um5p2pN8rIE0qLkRaFyh
wV9w5NK7jVfiTLTn4IwVzKjtDhVYf2RxL/k4Ch2G007gcN2Isblc69p3bzSK/xP/
cG89b0Fw1omR6P4yx/c4nRZnf7rNNB3gYamkUMlLKEcmx5HWuTXMD+dLnUidI7K5
Uac1vEnvAe1u+e9iKd1IMHcrf0/bX0cp7l4yFI7mGAMZs6ZZ9hVIDYgShgUiG9x6
kCN7lD8UdNx+3pnUApeePrgOcFiQAncIgkhK4VlO7BOoCexZuQg3IShSLXAR2WdM
Ok85AIeK/f9q6kNgl2ieCqJ8jTKV+frm26uPs2rGt8zJERwOrYcKyP+p+5EvX4l3
2i3qil/6k4GiTxXLWsQA9tDuSK6IS5gtDoVS6b1zK7YukLrVN9hQz1n/NlyUr1PI
IgeR/lP0Ys4vLv+/XYEFqrS2UGgL05RnAJEhLXSxa5EovF/kGdBndVymY+b627mB
OVZre3SjjaDfilFAjtXEjOGscXGcbV/z9DtXVuWSRHnzwpZC//gKtuCGBJkVG6Sb
5dgvILpGYToyCGPnJkK9LmTB/L+vh4XDSKHURHMTx3ikvUf8DG7MkA7HcBm9Gohg
X2PG/12fNF3AqwKExqnrVEVOXhSCmGBSJnewwEz8ohnp87Biy9G9w+0wuBPzErou
ZfHJunOWA08Fd9Jy/CJjfAIjbHyd549q5HhFOBgQYTRmF8rX2yIRuNzX+lLltuvG
2gYWU9xaoTSpYzls+R+vIBjFYlWdWdK1FvomsbPbI/Y4iKzMlNwOSS4rnzLVDzUz
dkKKuK2Au+hpRtGmoFooSFh5TwJ6lVMRz2lixEeBHg/80wMnwhOYFrW8uistadoQ
gJ2Fs7DchOW7ptpxQinfnk4ke5Y4OtRpogyN+a6OtOJiD6zsRfEiafo84nrCfT97
sUAA7hW2P693W7KU+PyaSMemP/UnXbSiYblUY45l33qMpQCYmfzqzuSNmzFx5/8T
QBUVIK7SEi1QflR0r7vRmUB6RiZoUGpT5P6c4F4OYv6ZGP7pjpfc7xF340yAAQOK
8rrqDtEa3rrvPkz47wDQXUBMTF7PtMd239G+zhmqTWr8Y2MhujdldAp7GXv7+q1q
sHREUZUBZWUxuUXaJcTQuR32O86YlE7/5j1AxD0h6VywdEOfNo4kykgQU3ebTeWR
gYDQtw/LblLJqXkBWCrfom0OUbP5vXH68D9jyZu9s0V7ig4mBHnqcHB1vT1XWW9v
YgkxEkVUWtYIpTk6Fp92Wr1zEjDyyAfKuqShF4kXwjaZE462gelsjJ8/NIaW6DV2
4mMkoLyu4ZOEp/zQ3/QhkJqej+pjOJnK7tVG99BBPIra+v9aDfNSDmkWhWanCaye
ND6M4+e1gp6D8jNN9KcH8DZl2l67PQgrCplWk4yknRP7rkz8k+1ekLzZWugZAQ68
VOEqnYn6sOW/+n5f1JBl7mqRKk63QoGF0FX+agLf4uqKr7YMPWae+sIdV3kuLijP
iLKizLGWjOGmnfN2PuYyYQ652DrSbLSW5T+d0wWjUrAlALgWemsk7oBruMeoLcbV
BoKnFytLftZRXo7EFl5pKVEcrS22VDT/7Ldzx8c3dz4PIoyQRgUd9HyDMirbniH+
THOvqjki72SKfF9SG/IHQjWjxtV3bkvGqqLzSfhZE1ioa18M3RqhpXm+vG/Jxf9x
cddQzaSm6nj91I9dWd3pDyxw2IHJlSRNQe+Zjll9n6UZ93pjaq4oqTDyyKagdzK4
UVnaz+GEr02wOiSVr9buc6UHPTs69OTVtqjpAxnZXsM3UWKI/Pn36yR41X2XT82N
QElxlegdkkgm+TFzEyH3WVDfY09CjrP5qwnv/mArROshekhhkwTen8xBqjjJ+Hif
hJX24CWVvvMdeF1894HrgTdSEHyPB0nTWYWMZZ8BoH+IuhujYjDwg0EAM4lvUFUU
LhdWr04SdpO4zN9Nh2my+7Ra9VjFxHwGP3AVLpw+NPPKOyUhHMrYbZaNIqikncxX
d7xWigJHANUGQOAhmO5MmKuLtTieujv/nt7KdfTRqRkpmkyEu943Bsgskju2tGNP
2ghxo5rq2Lcu6gljSxb952cdqiK+hMgaPpG2gqcj1PkZj0o1dpFjCk4Eu8uLeUuy
BbcJQi4dHfL3WV+LJiBWrFypphdcvdaThxXAWEHxI5nn4fe3M9QpK8u+J+pDpQqL
t7+It6cR78YHqqgNzLA0tH/cX0j8W9m7iIAt8ksIQL/J901/9GwLYslsvH0EcGw0
YqtzQU+69CpZCrpW8Opxknw9C36fnDKIEpQjKqRSmY9ohuZ8p8AITuNp3A7Ojyx3
sCdU70nPJrcSP0/Snx0dfd6xwqxou37SGkCpTwk5/Ak1BKpdq1g1GqTKz/B6t6WU
/WpdvjEil2fV2zOo1eUTk2bz/bg0C56BIRUTNfe4gyLqKhQD1VfPdAjFyrp1Y8uP
UKfwaxBjnqM8bGVh4WA60tBvOmTQ5KC1gMmFohH/fRzB8OqD1lFXnps3E1H6E568
UnXIdCSVubL1aS4zdMwNg0Z1JQVKASje+HyqKvJLv1DRWizRRMoguGGPxnmAea8p
8FqNmPrAWOCZA6pNzO+tR5iyLEaXMoJAvQQvMDoHxv5F4RSU7wE6ISWhiTASekCe
XmTJaNZZC9vqZ3kXN/AtvIUCnHDTRwXezHTIsoh11xHXY90xF3v7kn0dLquwdKqW
2crKwSR8h0DjbLReTZeuSGxHpcL/bo6EDzPnbP2NqDgAa9gSRa41WmOySctnBWSg
vW+/Z8sjXI6nfdcR56rnME/tJlPdJLSUAnB+abK5L3FCnKE1RsISxpEw0AH8F7Pn
7gyuHYEriz+FPd8h20wjT2SeK8cm7jQB4gnrMOz/4X9ON3QtNYf1DLNTOWjPWK+g
2oOBV5M8FnJs3m6n4m8UN5EWDtpoHZC7/Azr5jW7dCX/ghso+hR3PJ4yKixghyiq
q6nzuP2QXF/phKIxkYbNpRQb1vrMFHoVyFwbtSFZs8MyD2yir3ltA5uZIuXe7w2y
urcV2s1+jox2PkzBZ+ZNRsFv8xjJCgSzAo5JLmv8xdaVF0xHwLuue4NsRS3TiYfR
eXWJg/kPjatAZlxoN2litVfYxoPZ8JIRYvpgMn4BcRKC5a7C/vk1P9Ru10AQooN6
tFikTa3PAUjqKQN1GuRZcpyveuvaaySkDDQiM7dD2DgEbnRpdtphnMhsR914aF8P
as9j2qHioQqe9oTwNw6Qq7QhETMesX+WNwjkq7JDeeSTYUV06IvS1UIbyWDDjgdD
v3RYcxBh11S+By8+plpr++2yhgJJlftwTYqXnc/p1LzeGPUltIwQtBjKWQgxhJJi
5llHYHAh/ZcIVRcSK9nYKJQI/hz5bQz3rnkgN1PQRPfff8DzlFZVeL4WvUPD/zft
SnxhjGyah5aGGonSWJ65+a5zdj8q4WQDhwmiFePFy4pUpjjG9aGnAi2kdFxaP3b3
RPAIsOVVhs3E5Y0r0Pm6siucs9pOMT9eWUkgocfQTAMOwkNV4sxXZbShD2piS3Oz
qMRwBRw8DMi7BVzdBv2s801LUbMR+BnW9ILDCRj8wQRDxs/PmeEsMA31l2riGm/K
/OTazogHbmTR+dXDdU6buTwlRSIT414zjZkjfIwU2alu0Htc4Z8ypAyLnC12l0EF
+cTn7Gj7+l3dHaUcTDKZ4775OpAadWfq4BPDnfDsmq+qmj5M0PvA/AW7/pSDP+K1
h1OrMzKSzHNLuNfptV6OtdkrunbHjaXpQ22yvLZ/8ogMdiIC1DSFX6YLfPMFKyoy
pOx+v+RgqaXeYSZ4pDRy1MJf1rIGdsLNx/T7wv0x319NTksmxCTC/RvHJHt8JAb7
3yvZ6ck/t9njzuVux7zMzSvFECev7HYsshPyg7kKkrXtm+XBju2EN09OyNviZ8rZ
BGsQs8ePwW87sV7ZFvpHVEKiwUUWalTcqjpK7q/fc3lb6pGCRfAE1r9BN/IYx1gZ
U2FmaJBma1VBKvlXBuycdoOpqPicKMXJIpF82aYs9amC48zlc3R90pwl+FIBNjnQ
I78t/VfAZPtVCIKrggtbyTAkFSQGJbY2V/nYzRXHgeCLoA2VG1p6R8+p6q1UGR6R
q/BPEJ5RA/Z6kV8MFjzKV5ze9CQW51e0JHRJvjtv1OdrdP7XLeBMdcy9/OH8i5o8
UmwidLrxmVlUtKZHal8fhk9SQxAhlksOQnpP+SimVlrNy6j9rCqOWjNLvPlILX38
Em32Hzshya9PhUe+cCWzFDREVVn+VPk4kRysmtnOnc7ihaM6kJurWzfcN31Zzumw
rS6zw6lsIwDd3EDLvbzu9/4HC3IuiXAJHszE74kRxciMeiCLjRkGeYglueMQ8YP3
+MECnXVpOxrgQvpTWcMTyjEWGgWALiaaulWIX8p6co5Vo4XbmeaG3WMpmRF4KUmw
BglbmlIwbWqwl30U5EiMETBu1PVHvoKwEBYYZWhPPYB8Um0tEbf5DbuJn53iG6fc
r7/wM+RAAfBfFYWHv4c+4RZ3k9jyiHgvHlX4e4cZy4NSwfZUpvV6VAQ7W27WO75g
9y6aPpuBkm1jeIyjP6eyoxzOfV+fugjidnkHnvjZtOs9s5yo9jyJZRa99LjK8wA2
od1OV4v9KneC+tvgoqdloYcTkQz5upqdJty93mtiMTnrCYEE9u8IvUlb97kgzaEL
KoSF8PukdIl9DSE84fe8jqAi1hY6/QVxgvcj+tY3Jp5dAwacs/sJElOfCPhVz1HF
yHUAa6OWXpU7loZ93F/OqFoFolTNLrTrnY115hP9yPKTXgyIun03eL0I9YpIrPnY
Gx+ZnWiWhxq6X6qtMpFPmWlRnRQ7rnBA5OheFGc4ny5JTcLtr7h49OxHbV0JcHhv
Cau4uAl+aoXXLIeZ+z/zAyIOJIe1jXu3GHvSTGaAhM8tVaTgwIqPQd/03nImOtFX
8+JfYIMXVYXSqxBXt8pfDPmlpy75TYRx/jSXCS3yvxNB+0THszhaMoimcoqHQe9Z
/TrhjjrUQ6qqRBj4yGFo89lxXBm+qWuY3ZO1oIVbiNQ/b0kDMJnLWbw8BbDUJpIx
lJqBjiscNI9EbWvWIpYn1qzAuGvO9oVfpp6KF6RuYiakzqxUt3YUlDgf4/mtk71b
DixmLJsVOZZKTukh2L/eK/blDOsrhoi7S1lAe2LOUGP56uUCEDT2xhHAddM6/Om+
EqXA7/Crd7V6LSTtpLb20qiNhmInMgRKgUzHku8U/Q8PbJmRT4fprcEubxtcGoyB
IXs+17yNWfoPn3PdTBJVx3p9mVC/lYxS1+pQ8Qu4kvN/kq34q8zP7vKCyga/HKaj
SQ0wyKGNfTfVOi4b7SF7zpo36sWYmxONtototCynWznlcSVF8EwHB6FNUhHAm23q
jVA9yltAHv0ZAQFeZsHXX0VhbFv4cmG6hqAphOpEA7AtEolUTxOvV5DtDlCHXzjA
fwLAyMdJFusUeoZShViYzKsa5AgWzHVoRlQBtBAwMmJDEJG/4UmwFwTldjquMRn4
inOZIs7zSamQ7N3p4I+2W/Zn894n0cX5aBosj1Ij66GbufUb7RsVcPwiEW/Eu31L
lZZzz3tdW+fisy/2FGmXWTPivcwLIs2YRUyWDpvtDsdZCKIVuEGIK0NwXhdlefQc
R1tZthDyA5pVQwKNtBggSKaCLJsCCzEF5C+j+2QjRGQhJ4S/6r+D5XN3uHWBE2ZF
GLuUwJEJwAE+PxxV64Xo6Y4kbGusZMKS1G/DRiEWTadMRtwnS3WDPmgaBkdq8Esm
eecQW6zGcvj9gzlC0RtkAjFm9fyDOQy98gyqEWtk18iV1NKLkU2kzmygcHf+yabS
M2DX+dGtnbcAGONEkQULa3oYFTRI2h+9lbU3nupxPMo4ogogIwlLmfl70HSAzR1J
Ov0uXyYkePQXdhhiqbjdyVwLj2405vHu2XCATP9sBQvBmcmXzh19ll76tRKggKoI
riQK4k3eHW17HQq5y829qDKjtN7sl1pGeI73pLHvdf5YYROkJsW9qURQCD6NWI+7
Tw4PFnd73KuXQV56Aj1BZ48cBNZPJhzsppkP51O8yxDD8PD9hxgYNBavNyQ/9WLh
z2BhqAWFjq3vrqlln18Fwdy6ndKLesNUNXAV/BWsMdw/cGs3Fhu3MqAfo9FTbeMV
DU0weA0365EEGAlRrXwe3PCjqtddjuJyL92S7W9z0q4kX2YlKIqVV/hQd1sakJQe
7eSYxAy2QoZtFl/jZGehJ87U90/zrOPFYkgJkXsLQfSj2Ju8yb5bMs//mx/QF6kG
Xp7nfT9KK7dzBqFhtGluX2e+QW7YPvwNNCYsDVJGy/s5WMg/FcIohPBmDoNn6bim
2K/eSuex3Vrg/KSy66ny8BoWM1PaiMj/cMHCqCAwWy3HYWqBWv0W6/hp54NozmXR
/rmWuJP08xcyIcpn1lL0ULbbHLGJW0bOp90j9OL5Eq2QQtz+RDCx/RymLtm9uOe6
Y906TZpSic0DS7tYvVzXE97v6XT0AOUBU4X36g+nDapiExVp2ydbTECYg+un8HIv
8HWkHdFH6+wEnspP7cx8Ei0ZyQ7fIHjnWobMmsNskU25tJjS50i6olMCq/H2g1Xt
AeNqPNUs+8Njkq9Kbx6rS67kLDUhILc+HHSxa7TcrcchcqoaD8e1/gyDSnHnzmLn
UT3yoTJDdaG9zeS4hU4Om/ZVkK4Z9HCpRsxkem4Wei2oxSpl6wLnevAfF1h23Q/G
vp4QMc2HqpzdxmTZXoOQkiKqwYPEyFPqm6q9vtEUa51Gm+zTFQNQYTZwkXnQvq5f
YYgFmI/2YN1WOwfJLomuNGvFEzpdR2OPFx5WfpP8gwdzYIF+AFsrzTfDNuuWqEmr
bjXWc+V0veJARF2SkSP14H/7z3T9qz/1wd50hfpV6OMFf9ZDG49cZ61bjdL4v5yR
0nJfXmlI9CPdwRfuwnv2AUpoMZQQReVyImEtis1z2kmHka5sr+EAmTaimlWdf2Ne
Q91P3Rk+G8OKT0siGM3kJKvAnHMz52P30nbLIEHtYRNmkAWLl2oUN5E2MCh+XBCM
fwNuo2ACwIBNGngjfO95rKA7CXUj/17YW2PrmIRK5rjYikFKckTF+EvbxZY0kuyR
SES9mpw1MPIvwnazeBb6CHeXxhX7Ibutre17lq7DYJlGZdijVJRXoXBL4f8Zi2mR
IY9wdLeCcpNYmUeA6bXKIdAAtUqP/Dxa6pB0kdX/HTE2cNmlucc3NsBJlMARU9pX
HRbkpsU3xcfGc7PeE7xka4Cy4c9n6lBfSheAtRXe+FJUrdOQQUW0snK/Ge+Kqa0P
BACKIE0Mw5cER4TOE0pGrw7ddM5ZSIqW/JT64gcgPZySirRuuej/toSfdfJ+vZsF
VT9bJ9FQVFa19yHV9jgKXxDNhtIxe5MCvR5SbQc9yuAhw5/d/4G4x2yXdd/wFNhX
IU1oSJH9xrPuSJTEHq9V+Mm/xOxuMpvy5IzdMnTWevtozI8C/b3pVkyyorCowz3a
/cwJgtVSJd1OnURTja9EPzYOwUDnnNzvzJyGU0kAL1CwFATg/a9ynck3a4pYOZVx
J3mxom3JhmAu/bzCSxANDu/UI4S+T9fRoXsXdlWshm+WmQLZqv0wpCZJ/Ry+Y9lx
AmACG1jOUqVjDpKQIRBYpAL96PvkSGX0r5Wj9nqXgCTSt/TeYGwCn6tlJ3jXUQVK
mnOcF50MdUCEhJ387t4fKWPNUN2LoBaBbaND1dUMZLFdSuSO4ly9pI5dVY81l+BL
iSltnPy+gjYTRWAobrt7/ZhzEihbVyvEXh6r5a67rx4CeVGbM0tq6XWCPKQKwOrW
`protect END_PROTECTED
