`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgqF26iu35Nv82jj7O50HuF6gLyp+jxsectGjRMnGa1uUMgZPPyC41NTLBv3yA2W
DIROl9BfuCZyBJ6Yq3OBSPb6OIuMPpmzuWZQGNhHB070liYtXUTOcMzsO8z3TY7X
6AVJp620AXSUIE7pBzDqvQ1lLFiVpueWB4isFeXNsb2yWk2NKFj9MoQ7cxmCDqrq
jsfy0Btp1aCV0c+/JkRwre6Z1d4XZ8vGIVbtAICgCHFywApBao7bPGVzmjOs0039
xKFPTTYn9zCxRToeJgxJB05qPaCICZgPCnMldiyee2THhAhTtr2VyJDJvO700QNb
4iuzJYN0tyXO42xzBlmRiYVgcf171j0OHIcs9vIK+fAqs28Kkb1yXCdeefPJhxO1
iMU3J12U4hWu/qUdx/EufbNYWP/RMSZ8a/woAkCTwzw=
`protect END_PROTECTED
