`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXgwwmQNYdfA7KLmnkXIS5S3og/In5a4te0KuWzW/UuqXG/wVRAJpbCy9lLBQIQF
GyS699hR7mVlLAF0eZ89NSdVlh+d/yH1kOXdKGClbXf6sg4+DOQZoMg4NGKtqEF0
5SHYvScNPIc9lfbBQ6UwYNsP6F6azrPw9SSvhCRv97lFtYYIygUVsHVid5p7JV9l
h5vea0F1omhN7R8RHUAJQjE7Fem1iyMMudsMO4kLXCubkPcQGgyb22puxN8nKdIr
14FyEkvaa7ZrQRHzKDNKHyNG6CeApMtjxXo9xXVg48PVRADlc0Y2wrQI/FE48W+0
UN4P7uql3N6v8mPOTQFVnDcWzrNItysNuUC2nB1/yKvgSfilh3z5hztBA8rhT9Gz
yy8CbtrsCxm8PbRzd2v2Gw==
`protect END_PROTECTED
