`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26icUYSDEM1/qBo+BI1fCCwW5C8DmfHkR0XQWQzb7jFDXzZ5zy4qQTDq/tVQtaLv
AT3MKy7OxZmK9XmESW+uUGnAB63d90XliAEy17JOpLfcfAZ3oBa0KI/35KctG1et
xE2H8zTvIZi2dwWb7YCvbSMAaiSV0qznSFg0HfknfIg7h/Rb4yuQ2Ll0cPrPvS2t
vd+6hBinTb4aP6QUyLMahoTK+G5nfHAGsPRtnvnVZafjmYjUQOC4mwMml7jO++gF
/1y42S9UZN4PcWga7NZrwGUyK5YSZKYSbfmqlkaUeCMmtqc+MJE9z9lcU4XToFKk
wPYWXOyD0IA3YSfPgYMAnEhrKuwsPZZPIaGmjsUtgOsAmyK+dkoEaxpuueSJnb3b
DsFQJEXyQecMYFCx9cpNT7xso6SQKaTITpx7VI+nIfZzgn0IJj/UlrYtmAlBtKtl
y0u+CvzUcDG/jzhN3kQAMfrqErXfMJak2ZNh/mkh2s2+RAYRBXq9fYlSyn/hrPOR
lgJEOmqoq080o0zUIazjgXWWTg/J++CWEl1QS0U6JO6rZWsnJqinEqwVzBx9SQ8f
GOUuUShmXv82E7elyxd4gCvlcZER5M6PgLuGMT4hSvl/6AX0SJVHZ1F6G5FUwoqS
AuPlyzmi55R2dUqvP9WDAQ==
`protect END_PROTECTED
