`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kxok3QtpdD7ZW8ke3UQy2Oih9hn9mAYT9sEDlCYNZy08arf85HWP755VzKapxjKr
HehN6EsiOSySwU/oSL6MtJmAYpDy0lE16dFOtenUbTtcrpZnXnvLeCE1RTwNOxg5
FA1LXjCFnZ9p6+2s6JJdW1CSpwIxldHVuLu37yhwVyWtMU+QvybJSUUm35KvSBLv
8y0D2SqTBEKuW0q3ZYtvUUohIIJmGNsJXL7xZ6mQ0YBqdEfK4WRbqMotchJlWLoM
1fw6Kj7SI4E+FJdzaiH871sOsQYYrtAlvQ22U5GM2dIhFpKbwTDhEPNyobH5/Cs6
4VeNmWa88EuhzPP43PcIOw==
`protect END_PROTECTED
