`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1q+bHRp3N+ZsvswY4wWfvy67G8/moPAqo7u81KrNtOkgnc/TfnMBaRsVEdrmI/oH
mCyHmj/mt9kLKmg1eaNc+KtNTkvAZdKmjOIkEgh48t+b+L09mg3wixkccDb74YvE
b4czPduEBlPI1GIFZd7+oKqOwAdDxXT2Z7EMQ026Ai3KD6ycSKnuJ7xSdlnnPrmL
zkwq2tduGDXA6xUIJNjBE9YWA+OnPp/YyWm4CpF7CHppSrHS+vMPZF9EjJRbdlFL
16nE3c7J1edxxa8GI1pC3OjqoaUw1g5IPAR2JmjTQRieTdNGppBntz51BzV7X3jb
PDxpbKSdH8xr0O18dKHEP3ndzvaV6zhi7nWG7MRYz8pWVsjNR923nMsR9K1iCwpp
7HgYIO2kzgeyOMXDEsvGxTYg94ChOcoKkGTvPVBzoMVc1loaAXILsw61nwZE7Hox
fcHIgL5HGn5Q3TBbzSvzRoAj1LzxKKyCu5cHNXxlO5qgR/fmDSInG4dO+6bc1XLR
OzsDn3T7HMU6nDue4ao/l4rP5Ia1DmBHHeFq129hrPh/12b6EUvt2IvgUG35B1ZW
Oqnp9T6lpUZ692VNdjaWb87ETISC8VncLXpzWl1WSkp09ViZdl8JIDAbjZsBvm2/
AlbE+iBPogPBu9kREKcJdBynnhHhmZI3FtQJn/gNXFxuBw1He2ZiLV9vPYxatyKB
fKNi1gz0rsUUnp3dZT64FiAv7NlY9pT1rlzh8/LOtnLYzNjYFN4gNG5Q7co7w0ZQ
uzRCBHT7Xn3pTS8jc5wM8VMph0CnNIuEKSk6e2VS2DkqqYQoJO9hA10I3rQFnZt2
DtN5wqw/pQ3CT9gebV1mUKu8pfvYXz+IMDhpIguCx0M9yhB6ZUPoJM7Avj+o3paD
aazXrZHvWRxvMYSMWsa1jjdqMgR/b/PDvvr4hAPGbmhN1qtmJejgz8pHJGA/V8SY
iluaOOc6Htt2K3GoKa6k64aJhiS5fIG5kZG2GIinaadqne5/GIAiAe8+igHkRMmh
hG4QGKeIAy8ruU6meEvZD09IPvuKqbdYtQhB+uW0lvXC6u8JRfnrtRjG7VFOiB6n
/h56WdRHQrRP9kgK7JBiRZeTYjHjjPbz0r+YXkU9nD2+jSaBsKs7uVUn+0ZbXddt
yb9MRgdhVk9tVJ2iynrANNI33Gy9iINIX2MggKELxH3wZLvlwGWAvIiL9PO4Fdd8
qiRGcFl0PZXZ+7LeWSWM9T8bjRhs5F68qWfaEVXMmyEOgmChvgCsNw6ZlryhGX9+
O1AVQTrGAjJoE4Kquk2pvC7xDAwc65Babyw7AHDHHacQNXjfubD2Zzc9MLoxBYAP
u1BuPMhizYdkBNRYyHMv+D4xePjemBn3NQ/Da1XuL50=
`protect END_PROTECTED
