`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EK35UEpcQHAWMOUg+4Va8LRtyeUvtlZcjrZUB31Mje2fcnH6q5cWUVhMJtPLLmht
MxAROcnfzc6n2Nc5gonRJudylgfL6nbtFTfeP8LQpvjZ69QwTDmTSPIWkquacg5z
zzbQ0oUXIHRrG0K6PwMW3CroCbUI4yKJU2z69C4MEzpxyApzluH2YyiPr7LtOY6c
o4KlrjqA5wDodVMkyp5OBVcN3ehWRcp2LXvidIE9y2/KVXtaY4C9nc8r4ZQ5MSJ8
Ae7FyRdqtm91SJlGXYk6u4IyFjaj33YNzYhaazlyJYZf2jqkwLjt4HqEsFcmHzgw
80+NzCcf+/poyKeVBuo6qawBJbcT7SNkR1mM1wKTj2R9ONRtHhhdPqVyQJbmO7mZ
oL69pMHRqW/9GbPJdQQ73972o9Z/e2oQkP68mJhlGlysipLi7M8R5r2XzsPe5P7p
vtmg1rAV7rYA2NB5HFIselbpKYfCpagCBocHikuK6pJ1FYB+spr8KuAj+a0cQWRQ
JYyNFex0pcn+IM8gA2FubLc5RC2zSohHr6U18KTAIZce4XaIVr/bBP4PWZ6uc2g8
S9fDoSidnrf4FxFsuFRoZA==
`protect END_PROTECTED
