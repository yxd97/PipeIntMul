`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzGs7oU6TZL1EjjnB51mJt6glw/Th0FTa+8r1EL2P2QZvg/IGNPNIbYCICkL3NhQ
WWKgfx7MfS0cvOoxIHsAeExjCW6cvOzpxTlgibQlQ4es+NRDvsCKZKWuAG4T4Qzw
fKwl+y8ANWBuzgqPiU7tXkXtlf+B+On/sW1t0WoMD4AJGfBgTnaF4u48hAzCx0MY
4EExPztYtUgEqb6l9Y04y6RT8JCV2Z67Y4baf/ukcuR15NI0+fr8mohNjyw4HS0h
PGkk/Si5vCSW8rs0AsFLjoobaMDfnum1/Ep+oywNQnUOv8LY6uK6AQDqOuetFx+p
ylKLVHSeprvo/Fl8KAlgLshlSvO0rxYPNExqW0JMqgumeEgPUNKMDXnKqVeTSZTF
oa88oiudemkVrQMgmXqy8n/R1ssB4Sk1TijEpvC1mlRFWMkKDA0wiCV+Z/gy4o9V
3OoeESIvgOZePj6idJgIA0/4X8j/uFYxucKJE1iSC7YlZl+/X9XSvWJQ6AdRYUwY
xqk4mpQqVyrISfqcALm2pfEG1AqrKb0VN12hFTf8DdEM0VjXVxhuCemBTbsXbtsB
W3dvvt/3QAtMmK98OPdydId/66iqXlu6A2jcvxLVS7g=
`protect END_PROTECTED
