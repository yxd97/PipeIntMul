`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DHQ7UJ7PcAMMEStLe06L98yVczDZLletq1bnq/0PvXtOZHiavu60VlNSLLHJ0KZT
WWLw+sT6fFdGIlio0vi8YBc//0WtQ8b5v7p+V/gX6BVVl05RA1YxArx1PFB61aBC
Z6Ej4wxugPDxFdM+sb1JLU0C0K1JL+tKM7Yg+36MwaFrPGUiHGbLx9Shdlbaf4kW
YFRjj4ljsuFq5evqvvGGYXp+pmexefYVvptbZsYEuMn98OwFDxEIkFfuvYJUF1jL
j4XaBszuj4iwOFAWcO+UmQiieWcLaZHMUdKUsG9YEk4=
`protect END_PROTECTED
