`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HB1vG7ONn+Lj2zwV8yjx43DrdrrZQ8q8EdigNijquh2h8+59qgGbBQz8anHoc1TC
P1KQMgxwEfLZK8CxUjccItRQT07pvBvp379W19gp/R6llmDbZLvRGcuJNFX6n4s/
hR2ut8hZ8I1ZorxIwM49u37BamH6fht/7pfQFIqWM4YC0Sgic/TMvwfS5kYmnm3H
0L18SFqm3UaP457SPJToKf2XZ9aJL6Yw7BlbrHpCzrxxTNMJNZoppGe+PRTmAiyU
988YMRMecFp8sf1JMq/OCThH+G/tqnv0CofDIQuE2wWCoryb3Q5Yd4W2CmaLF/1Y
ezGQNAnr22/scgG47eRfFgWVEyHZM4z8O/YZJnV2Il+9p7armyB/Gtb2W7rRYZNJ
FhWMLUXZUF3kKZrm4JCe5kEVeW0t4vMvxx2ZaerUOIxtllmOEtEc+Ee10JfPveGM
3D8zH1K/eDJ0ztyx+5TS0WZh9U6TeVKQcvTgfE/WSs6wxVymTGJwb78LEIMTCslN
VYJIjivEZJvuudZ5EhiUFRYRTl9E1fTqUfYCBIbllN6jLqIweHCUuGnha3HJ70EW
4cByJ+bfrYKNYJlYoCqmDsZUc1zbQBiO99VNAhuxhkLq8a/GIIYtaHVms2t4YVGS
HP2zkxTG/T9AytSJJyX2Utso3e2+7JJ3g3UgX0UWByfDEkhos3A6mZC1DxNgFBbn
UfyBqo61fhx3tKzDVTPcs2yhv3h8DYVk6M2Dscp7Cvf/rOultTwJA4VcApeQCFQD
EbgLhfqrJ2JrtYtPl5RGOIg+UwFx+8I9bKCl1N3iR1LDE9EusAZ3rFH0pQ/X+r8y
sFJ9JVSNsL4NerxdoNA7sFwDF2YlwvUxmp/c1d9oxKVrat30yE9yKHoRqoZDbeFx
wSmy17l1mWZTpE8zzc+P5+PzQxRqv8VYc8il0haROYhhaprxxTrzveGSYSz6MVkV
JCLGolvqbC7B84RdcgZifv9/qrsIi4V+EBwnaSGdTus9un4Y89AOgdhdt2aHxIY8
C8O0D+nIxXl1LBu2/iycf5qQ4M0wRd2paaRchlZ2TbaDPwonuhgI5PAR005HIkOU
16ZG+dkYFUZl+gOyQE7OicxYXNrcXAAkibENlt6iJEhQFzYgOyG11w2eiWG0ieFf
fWz7H5ZYzqMbNwa+2zPU8oMpBypMKw3oXfAWaeb2kuoeVcYngByIVHq22oX1RMqc
XFHutyeje7+1snTlTWeA3snW7cBDYANsdT00mbv/8NtKUBWF8Obg2Zd0HBRbzon3
ilX0Ez0zliVyFG2M375eZ1f1Y8enFp/8up0Wg/5lYqoe2UIi7dkYQu7z2dnv5pyf
VSo6K8nPYM/Ta3mrrLI85dVs4SuaJWcSGwwbxbDDssoJmIRDdQuh0AO86oRP0x39
hRw+bj0itp+emgNlEfWQIULpKlOenSYJBDy49XHgA7ugmSio5G4zCB9bYUF9o++P
jFk8mVghZQPOZBllbEKHglYPtz464y+NhfPtDan0u2Q10aBfOxFMSWYSsFIryoVz
AbPs/PqNgPeAJiqzWPW/aVIVcumuH+MWOBLcnC6wcw5ORAMpcn3a67Fc4XxQXivB
75EbuFFp+oYoTI7OTUcNXqAYGkJ5HVgMtcn133VVPWvToK0Tp7u6qeLXqa1WuHuW
xI5sl85HHKEcyROiSKHqg/tf0N64XT2cxmf+Shh6ginGuKqk1cQO6UtzxdxMacBr
z0HH+JTBfn37oLdjJvmM+KYPLqli5TgExGh5ceA7w3H426ZjldyB1j37/O65wlYz
OwB+U53RMtlwGbAxSULd9GSErFwqsauKKbI1hOJbB8zMviUJ6GDinOGuQ4JpFALz
Ak9KDxSV+6m8iqey2xbwFbooO2ulUI6n3lySAsNNB+BE0VjMTrxSGRbOptnNnNWc
j78G3DUCwR+Stei28SfwXLTq5vqRZeH3rGibT0AOAC8CuKGJEpCREszmzg+Xv/tF
7sVBe2NkvHns3d8M6PS+7YmN/sQUZoHpKhAAW9W/6CYKZy5d/AzVNbA9gUK8O6gx
HW+ZlmIEEsxxcDier1GczCeazl3daIXmAZWxEX5/iyGOpSmDKDo3WbushuE5isIB
MOZUVOX/tq3RvQ9yNXQ8ba24IGjIisOOtqE/IlDOc5xmSVbw0rZ/FbmwB1YAPKAY
abM9ZRz3M7+kbHYaqWjrPkYLv29821ydf0oFZoJMz6jQuskbDxbbSIqfYUZ3ko5I
y52KuKFMpzn1NoKEDDUMGSa0uiRRDORWZmcduM+YwTdJqWgn62VKApNch7FrLnnx
DsUKvLUa/TvSLLuPpgjtfKknrjrjAPr2fkCGgm57GxkNY+Ulh1Ei6ySqY/wPEdU1
UkS2tUGG3LDQ1a249iv4Ke7KhFGoz4AzhsHbA+FWcJUerCaWtX70PUrDvvLh5ieH
PLOj+qPhOJbs8ffyYXwngDADi9T3Dxz9RZywQstrvSy8kQ8jOOppgDKaki8BLECV
3LHVooEi7OC9uZ/FxdEtUp4UBDKKcF0EH+kASmsGeWz6OBZMJ5ZWPuM6OmN9EVOd
IIirUquvJZ6qIB7U/t7uT/rEaHPXb1AxVfsezJlMj7VgoqbR4ZCncpmU7wyBQqHC
Qm9LrfdOQfd9y7zJjRsXBSgu6eK5HouqgKEUt7yFRSDCpVfAKrxhIh43TaLrV1hK
nZezLwun38tn7JAbxi+RaXHvtCXgxuCmYWhjflYRCVT8cqyJ/vQZxiTuZHXDGCAz
Z7Vg8ol2gL1GNO8Qmj/EFSzD3sjjshCafEPGbhCEo4d2zQewQEP6PeZFO5zgkF1H
jOWQJvkA+vM9PJJhY9te+xAZnfnZgmWmpg7DEUhbb4ZWE/uM3irt0USi3xpCnq8p
+t2h90R3WBGs6WNo9fiwDZOzy5NYKcC8kr9luzJZGkBozQmWOqDjxyrjcMeX1HGV
jPiBtFcKBg/Ej8n0mQ2mgXjZ1obeQoQ9zcoSEu9uyt6BTUtXeonNfbVN8MbgHxV8
9HybMCV8ciYnjS5hgww+0rHfrpRwzWp2JRnnHIWZnrLjrU0rl2jemyt/G2b0aIfj
7rOqzT2Ow/h8V1pA0o+b6QPTJtFeEbGPldBhTvUwpTB4cIsVd8cJffv1scrbVRJx
SUToRnawkYemCLgPN4a6YPKlzUBohvydjxEQoySTgx5WhHpemVnlZ+UsjQMwkcPG
XtRsJLECdNiDEnZPMohPMZoyCsXiu4aHud6HmjWcE7vNRQo6yY2gIwkr4dSSDuPz
QmIDjSc1GLcdZQUl07bcks2fmwjr+aM44+LHR5c/du2x74HvJAhCEsmNqsHAGtmt
HmGWjjM073XgyseRUr7HzWQeJGwyKTOSvcXj0NYNIxX3h2ZUU6DoCPuD/3ze4jjc
dS+9XFUemiZq6SVKINSSf4Opgt1BL9oH+kgMM7mXKtfyznC+QwfqFmM2X4Whxlql
j4bOO2a0zKLcQ4TLXrlUXxiOxJH/s+V51+NFPdJm8tCoSz+vFthxiwNDqOHFsqLE
1EPsmgH1QzgSQqJbCspU9hTuaaacgXAouXEpTUMBw/Pmn2ntQ2QiirUEDYU+drFY
elxdyBKMmgHoZYoViT94FdnmnuJCPi+xi0OVRZP90UNA1SdD9iVRHy5yP9DFONv3
`protect END_PROTECTED
