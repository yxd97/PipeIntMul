`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4FOdMcjcHxfW75TQipJkCxILqSGwKO7BYaD6LZjYdr5r2ngdNFqX8bLl0GkV2QcT
Cp7VQEzKFiRPHR2TTM1zqVcqxeFZ0JcrszOk7FTxFzrn8xjH1A0ERrUwt2ppXtUn
1VAbgcjc8gwRVCw0347sXXI6aTPRr5NTE565Ge98fCXQNTw4R5a+TPGDp9rP9Wak
tU70ERcBK5UJhNzt4UOVp7DKatlJdAezoQpDA1OvsUeD6c22IpqUiz7/kqO9vabo
twbkxco4AFCDFs0p0xEnBkZwGniOl2M/dSQHyqORN7BH46ZXWkpbkJUMmBnT0kYc
3zCiEdWRYj40zNEoRHoNkw1/KZQHrR4XcOTzaddRsMC6T0cWvkvd4PvGUxHfqutl
1016eyrt+f53irKFAHy3AEo3trj+601GwokKHwCuZyj2l+OVH0irbBxsgkcAPoqN
9QAJDNiQjO+XqOOEVL6wAJcshiZkMm7ZKokpXxVOEnC/eZmkWJ/AnA24YxJTwtkv
27oH2/LNWy+0EhnbGEmk3OISY0LDZw3CPCUkB+s0HSzOfnsbQb+UtO7WUuDed6JW
LPKXuDqUfhXCR4A+3oRJZvyr2qbvfpNBY3IsVzIX4ShN89PJ6AejIXX3Vs/XZOzV
ImWZkTUWeLzMz1g7RxV6Czp8qqo7qQKzkwdiIinOmz5AW2Zkjtuvb+i+E2py7VKU
tSx3x02tJuSoww/tP3TZDaLZFSBKBPJXOuGik1+xYeD7eIbSvVE1hx8Xea1hla6M
JyeIppLWL5ugX9LYHl2OCUxNAGuabGQGTCF/Ka4lu8UGYvGYebKUrgzYnsueKRlS
lXsjpr9xf3B2HqDWcEnPZw==
`protect END_PROTECTED
