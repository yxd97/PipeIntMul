`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tvS050Raz5Y2PBo5XNDkKWLJTe00ip/yLx3QZhnLiyWEP+PA/TQ2nMZWhd5ngR3O
g5M3/nGPIpoMReC344zZTafNM4GJxB2wlDPo1kAjxiC77ok3ZOj0xG5k0vJWiZMt
1mYvKlnYkjUIc6ss74RnpZ/lDzHt30byOefhD1hUR7P96/vr6Kze+R/t3373jmSg
Ds3gd2Y9q+EUzalCvhPQgzvQPSIK8tloseAlbfgXef7giPaR/VdtvBWWz11LmuJ0
xvTBEkdk/RRz20Ma3o8GnnnyUtp0GJKvVzCvKq6QxOT6/IRQKBVHu9GsfwiBqxxX
GR+NMAFE85mHXDykFDo0G7a+8YZTUhYYI/alEEPMeBLnAry1149xDPb/9ZxOh8xR
fVKTSn8ekGGBAlV4pjr8I0JvGcEBzekRN3yLXTdZp2kIKvufM/nh8QftT/vvW90a
a6xN33NwRqfHUCXTXwmQzgm3cgXY9RAeFng6Nt0RXnkMOv40E6TdoM3V0x4f6b2Y
FeXB+cPc+fnM1DgTr7xrz5TexgMpPP81MjLgsSPzHuHOICmzJaL132DM/7YQnWXQ
6J7XhmjmeJ/qNhJOPqUAiZT5hFmtGJi6SemEFSgWYaLdZCJAC6TRBWua11FksIUK
y2gTZT8DrHyC2KFqsc/ZSRhxriHOga1LTv8H6z8UkXdeYaHfJ1MqJiKUNkID5nRI
M84HQHiW/2tNFOuzJCjD4n4aXvlCvF4QcLMeugkQQWIKbyW0M2JTjDrleq0GZVHt
AVSscSxr/7f7WOJhKRovWHh5l8n6sVeMtKVIkNYBjqrylNNAfWPXRb3dtUQkJ5H6
2mE6JKvN6G//idWqJ1tjF9m5JOxi4afD8+vKmPAaDAyo2hISeV9nU4PcZs8uRB+6
C1mmdiClKTexTxTU4eVMkPzQSIurTdvEYSyJE7oMOFcjC9LkaI0nzpdoLLykWVec
a8q6SksSDBvGBtdQiZXmOs9bAePr/FEtCPKcn9Q4UxgiED0BOpuF2LJvSbN/coij
QmHjHK+KNQe+qUldhN66jws6Otlt8Ex3ZayMh6aRs/Tx2Zc2qWOANLPX/3ReJ+Qz
UXOkDEglUPmkgd1bO5ht9OoatKLqAbqg9z+n/0N/9UGePbwlQWGTAksp8I3a/D78
JzvKH3jkFvl+DKb1ST3PA9u34rJPxiTVIUaxgdI2D0MuPKlQ2+r8fCVMi+aPnEpv
n70YXZe7jtxKTw49i8UEru0zdby5805RyGOJmIhPDWRtByC1UTwAmFlq1LdfJJHu
48W6KegNcI6xCx9UlQcV1dv+ZeiFiY1HG9AK0SUFkzL+lNxllmAQ1tAluSmHSKfW
1WnzoIRaO1bflG2NUG5lNyxKsZrVPi1PcDysw2FKQ0PmoB0ffJ4eSlheLwIbOfhX
YLigF59aeFS0B9U2CQVvD0Ecg3IFKuwCh1SZwfvCnjsmLkx92VxPbuA/1+X1A2OT
2HT4F5YyWtxyvlU7joujFHBz3YZz+nbIGgd88s0LdoB+rH2gM2JLrBA+FRrUPLI5
7bOrInpvphWYgTeYUHI+UL0E9hNxFh4h2FkqXLEqzk2qaDfI6sjjgdkL2XAezO1F
kh0IO5bD/w9XXKmtNdDcf1h/fFLT/mXGcat/6zLff6j0vehEtbQyHE51AhkbyiJo
QhT3hj2QyGfVXbyyKPxKGquQl9+bCVJC+AdQRGaHpd1D1SnBtjpQ6FEeFDZzPoDj
uIVIGSBu9gs6Hc6+904fZ3Ay7uBYviGmdTXbSI+nIPX251kkTGyvwneGAbuIKzcP
PAEcB3iHGRwjY5vPtqdcvPblTFFFBKigqHF7IegE6WKbb9w2FUV/az0StuDBxFzQ
i7UoLIXEErgxtip8ztR0mQk18vaDdEXAT4qN4Vfr7y/UbM6eQ44+6rXAqb0IuVXc
Vjk8rEI2RsHcqQHvyXtqGVctOFYD+RVkxoAX/Dl9PaVHj455Ecp0lWmxsp+umAua
Pj5DSTCEa+qZtPlt4KQfUEbzcArQCUUQMxAnMJo0K0NDtVdvUXYX8WruybfDLOn2
aS4RczCnUS8M18nJjxy5azPsZCK6/oud2QFRJ5mwN100MHhcNNjviX4p43WeyIWZ
8kgvtLTXfwQ+/rOTpoewtqibgyAfol/SP+iVORzjdxc/9CpbH8n5OpQeVYHMoCVF
j1wCYvfIF2SXXyQk+U/7WLxtgX14dEiQKcfzNkn865cAvgJuGufVij8boJ87esjo
B0/Wbyld06vNmaHpL1h+Opy8I7SGNqLXM/rkaAUQxp9i1dPD+K4P+Kdx1aupSGKX
Uin6SbcZDvMxPhVZRnrV26dwxuvEgXOugkf4S2mTrAz3WTShLLBQ/EAn6Nhb2x6S
iNn7Eu3XaJc1SXmdQHguqnITfjns0BP/uSPGK1mdEuFeNKBdC0cPh4nV+RNKw8PV
bL7lgTvB+R1PZqXP2kXoDNpDPwGZNCpeKZbygroU5d04jb/ltWRkQijcOCClKdfZ
bJXKU3w75iuul0vsyH3BBEls5m3jgynhTPlF9AE/s+0KERR4OdXEwucMVxWQOubq
x/ZjZqUUUe11xIa25Jt42OZ9i2iwE2lZTIMWLvMoHs5v9hBTeyejP2FOxtpOfDtt
Dbx0Q7E6dR5MTGkAtWeZKix2DVEG9pYNnC+93QYVugeiN/FfJQjta6Z453uBzbHT
BRNUo1s8Y95116VVbWrYleMsKjgmDK940I7li4+O51wJ+DLn/t3RfN25ClgSj8Sa
82tZzMlGxr8LOz7ZSK2CwM+EjqIeJYWhoheXmfMqvcUigML3GB1jdQVu1+TVAbL/
FpPJ74Fn75QSiAc919dSiVzWcFu+4kuIMOaJFgHHA80NUng9UpKcwvvcoH4fkCN4
LUlw1n3R/URGVemcmCBTuFOPtmrXF9hJSkQ2dM4tlV6JjICaBJOiEoz5SOU7PY5T
vJYvFXOf/IWhWLSmHVrJ1UUGYK/aNYF22PapeKAlNU4Fj+mMuK+Wt6+XRhZTvfBr
kD40a0+nQAUmJj4nov4WdVt+17smpBFYw5h1c+5xegP0uI1KMsyiLn9zD3YYHz9s
AbXgmFISOBSsVacyx61bBEWGIC7t2NVMxgFqLvCyUAhzgrozHCjg5c/fbYFG+ott
r5wsGvki4YfXhTBVLNfaXIq55Jx2CrgC2Zl9p/Nu2v00eHnmnTof4EsPX7VSnxIG
YaEU2pVFeMn7sBn5wr6b71poH5Su/TbPf/veUVHbi/Z1aUgi/SEHcDDgWD62o+Qc
9FMlb+i0GC/TRBy0OJxUI1lpdYX0RJdUAXRb2PW8V/42BY/mkyvyg2mTnrnmTLfp
70HVcmfe0fIUgoTTFbFR1PNhpAaXF+kOkmCpB3/VOtjXSxFPFS+mZUmkRDLGOG37
TZZAG9ZtouKs1NbvuARE5lbC/nE6FY2bb0yBs+rMfgdHNkWrXMtnQEGrGk4bkvKC
5zia/6zKGMqezQtxZ9aZLkt4mzMRe9eeFG0CGPKbJHp7xesl3CFyVHolNu+julUn
UlItaWBHGcQ+mWBKWhMe9dEMTO96e8zjdaerRwkeJwznNpPdgMjz9BGR7DXNHat0
T/zlKNk7iQuAywyPef3aSDkdOP1th8Xa4JHOzk/pUr+3FDgMTV6po6HTyCMSK9jn
T+2EF2TTORz49DSudp9kNaKCwgUzLf2HVmJKWGde4Nm5Kclv7yjM6Gw52bvQEfjg
xrvZDE1aQSe1VXuNuqiqlRop0FfV0kqGWzb6OH4KKQ1Taww3qeiTc7qDsubFEzkm
EADk8HjNCDl1eoxomK4Yku+xeBeUIulE4XiZ1ETJUaQs0HW1QUssF8oV0PcDBY11
Yz5jpsrdmNpQPEUZSfUWC+MJTMgkCVKe2aVe3IdUcW8DZLzc1jzDEf11mGONSH/L
7GrMRMEIxPB9Wxe810YnTxwsMvEa+0JyeRi2Q2TwDMBzAqoLrBKX/rOSU1Cn6lez
pCDB2AL9Q0gUu/3ipdZnzId00PzBvVG9Guwu6Qvo0pJlcD0TJWnm8NJbIw+0j5PO
ycn6Cld03amdiOpBQQ7blPgbcE+f/Wj2Th255SMXBiJbcl6v9/QvOPAXhWnICEBD
Tu41f38V0GzxjH3Grzcp8J4lyW/VMH6QHwq3o0eAkpEF4g5YuWDxe/bhMGYa87kv
WEetKP9u2lc/055hG/KUxFqxj2fNTUEjwMoF73vXzdrzMMgC+OUByEw6WCiNfENm
8a22k6XbiWrSJ5/I8VgeOUJKmCMwxGzOkPzzZkJA7J3CV8ycGGMn9SNPIScQSSKc
GjZKC11BgXhB6KDDjFBmy1Q5tXpZTWpMf4G5LxwL6mY+5gOOXkkxO+/BaYq9CZvr
HQf/JXR+ir1DwTvsi1G9FqZjztZf6b+91k4PEURqArFFYisnjNNyKT58BIZN/Z3s
ElTcSu1niK8sbf3uQtW3we4ItM7UMXF6YaaXWB9vJ9GIyItXtmPLI9YriKqYuM6V
oGoVjwiBl40f5f0/TXR8XmBf888kE+AyhLTxSeVj67pInft7ocAgLg3iEZNTq7D9
MduhugbTNmq67phjZW2YXGrOBvLCTkNsXL4dY8oNcy5npHweGQZNAWhMk6K8AJdG
+xtjMxYmlIpxkCYSx0988iXlV2rcy8jFYnL1udiEwxam9GjAeNOXS6ZVW+s9VfBa
jTumGi+OL2ibY9Eg+t5P6i2p+7U/8W684Bm0S/O3ZGek2rj/luOCccdm7hOf4pgU
av392XlX17wDhzW1CrxM7gMKTowf1Zeiov9Q+X0KOfqU6VNUxhEIOfOzpEHjpeTv
Cp7MHTqDcv+bW4Yt/WD/y68v0TJ6kwAHLF1fZ8SuQp2XtiS49hO6/bd8lUvonp0s
RXiv4XBAiVaibM4WQZXtKm/if1Jpb9ycOhrQJoyjCs1rDrd5qrQreI+DaMapRpli
dcv/YD5PInl8JRdFiKhkuAR8x7yiFMZ72QmVqfZY2ssUm5eMVIYNdLXPWq2SVWXH
S17csmqjywdcZEPQQeVFer3gw67b70sKg2oiwqB40cdgU4UQE31zl5jVizlOFWM8
fpvbMFr2rXpSgYSwLQ8Tmrv8wdcoGiZmTelzqn3eo3P4w/0psKi6+EcQrsKPnVJJ
EkAc/sodE7JO81Mi5Fs0ffQdsySLdP43oiwmBiKEKaq7tc6yiGpzEHdOw/hQrv/R
shth3/g42ODcuEuWKve7tmW9Hk4s9rVy8CcizXIkEFwezIndCwdn5BB1lM7O4uG3
sECOu7LbzELWVoNAyWa7xIKobLZzfLthC1peXVnnF2xySJFXBJRoFL672sgQX3sP
CJmPP9y918+6CZbKKqqHhSZdbBwchbCWEOXy/RT/XnQezihjLnrwIcqgTgHlnAUp
/whLIg0Kk2/jJpD9xpYMySYCeiInlrrIqBd8UnDg7NgTNUlA0i/7cFCFJu05Fa3/
bwhEUazg8AHfIw645lv6PU0sFUFmHbIYDcr3zpuAOnw5CyePXgXdoA3oSowm/5uR
eIZJomHkoSwsH7m6XgewmocIYVuRW6QVLPCCxfWZ5cdutPH2i3IKvC3CEPbqwXxc
HF69+tiOI5vfRV2jAYhLN00PfVIxZbG3/w/bFIz61lliuiPuWWIpb0iDb7HyYe2p
DNkUKeSrBj5aw9Tdw9PZ4ob8pGDtHKN0xmsB/Gd9rPkBtsfKMDj/ooAkhu+Vcd2P
eZltW40NzZogrMRohyriGs4iRYxM+CjQIGV0DGVQVFE5NPFuhiGIa6z9GVKw82eK
SBFXgkopJ88uw3ckRQR0Z2ZBHYw3804O/1Wq6+7woNHMBOAXkUjCopHFO8InkaYs
hRldt/zUA9rmrfRurpNDCQblLYiiyHI6PuDefwgZ2YOovujjXU6O8yos94LA/EfQ
QhCQKAcIRHR/YoR7fTf3gD2HeS6dYfPjB2YUCIHxfllT25YcHAl001L+tJePCgQP
JaZUv9WIcme8VBKmNkCFYDv8dywfTlsMIReRpJ/DqURQwzMGyitNTIpU7uNoIxFN
hxEftXQdDBJX1RQjB5uhRQRDnJ9UmzDhFvm9NOb2rJcBzs//Q1HGYC0S5QGWD+Tq
9UFsYdQDzi4kF47TtkmncccRN5jVs0e5OWJrorw6PIBKwQqIsnJOHw7y/9KPmDgb
eLppvb6cfRP3W4/x4MahloZVVAncOE4mjGUw4quK+bT0QRiUeAbJsbp1tHoc5EjH
KKmUq2ZlsYmKCr52oJeYu46ps3m9aO9hEQiP5cKgXyj4WUsSnWHqhLQiyJ3+MENa
DflGWInWv8VBsfbZqjF/rJQwPsSU9g5PE/Mu5cvzVoq80vsJy+PP7ERuoIMZ5IIK
HkbSz+kHe9KNn3hW+GN7CksTo26bL6jVZ/fL/EEOanGXLk0A8cOXfj5QTJgMpu1T
PXDCjUAiJs1ISWEIaONxcDIDhJB2o4uRV8w02PGJCl4o1frg1FFlFbIX3FJopCvI
mgVvGdceJvWz20YhAkkMbKazMNJvESSvi4+P3u4TWT1D7TdXkIVd6A3gYqx5XCGa
QmtnPXJPjh0qRJiSAoUvvc64y/1P9U08SsqENy20FOxRSRFVcV8GYFE+AjGABYeq
O91/FhIzcUmcKp+NaUDY3Qr4F0ljXdM7uUw2SzcqALFoq+2Yiv+pgjSBLJZ8gXJT
dAvjNEClhNIyTVbW9lbumT6XHGbN80PAk3Tn0lEzqADg76krIUZKMII7eNZdIVJq
5ugncKAnyssexfuSY37DgBeZWLHQkKwsM2/L8IEh124k/vMqviU2SK8dG+N2EPsk
V4mjTaBQS9VKYn2eIa/M9mW5bFUPlUSDX9HiLNY3R64YqZOazGn6+Bnjz4YFKdgR
fnNh8xUCXXlzCiuTcY8MzXGmBC3r5a9OCvi++yBm7MdfAnhIfJGlIr8N8ZVwiR+0
Zo/2AxUkIAUZH2SW5YuU8EB+LSXBXMjupBIq6+IvlVBfcx2NEZWIIUdwNTUwxN2m
ajq/NZwmD4ne8ImLdMQInO1IsShbJMbQ825D0t4lLRAddisrjQmvkLdvL9LSCKzJ
CB5TcoZ/z0q9vWWKICtxJkRH3v2bSjMluIrup5wnSoBJYb3mS90dqBmWrDqCbMQi
VLDeQAw8E7oi4kIHVMsnNf+XiPt9Bdjw898JU11gl1q9urx8Bi2CcMeAFYpUbKaT
reJzowkSUFOIixJGwxBvE7pfD07ffFg2K/aK3LMWgo5/GsvcNRaXSHISmmZVj2xA
EaWW4NSBWzqSLcmtrcw+uoLfGZZrAMxfFAu/Ejfq1C7AxomU0f1jq+cUb0iNx5x3
IwdvYcLtaZAFVTLoC1rj1qogObjfdjxKmMSXpGNCwNrEMeWKY5g1/J0hEfgreolb
pLXeY42U0zIpOCTKhlWUvkHvVSTHLaNbO2iHai1wRck+WX/Mn3SkM5c+d3vsEXyq
MjvyGF+kuLYV4ooc+NMFBHthGM+6pmyZeY6V5FLV7zSrhs7LcnPT3cnflcqlyuqd
dYEGI+NtZ8ePUnXWQBM2w5pSHUOL1ijvcaNNgT/Kvc6oWXSzTy0XKfINDxV5CIZk
RxSEP32W97Lse0v4nAjEGSQByCqukEKElg8ZqUz0yw/CPI3B0yLf28QX+iXQc017
cWuIj+SeipzLS5HH+kUxVeyy96Ahjuv+hTPtxibhmMn6RPDEgwc40RjNm8FTjrIg
bQxCBO/ySzyLzxbmZpp5I3d8D4bMDEYozKHVu+PJ2cL3/c4Pyo4VJO+DdoKCOMmp
0Xcul/tdM4IdC7p9gINfTxMghK0WHDSjBODgNJGvpNTAdffMCdm7H1m/2y5aEq+i
4Zsm2mkcVkScZf+DbGRbj47+oD38xWqFapUf8ToZneR9Poxb7zwkfgQ3BSs6IVnp
RVuSC9CJGJDUtGP4im+w8vRSdHDttXavZURkbcrBPXSrOWOMZbbPVmVoKfbDrj2D
DWCcbxoWvXVVvzoRjl6dBB8+O8yadSxMqvsiM2ciW9cPymnTz180+LZaYjwv5ylF
rTAgltMH+w8SPXLah2j65gTbzpGWRni2hILRxFayEnw9h6u73koCowuYhG6hCU8D
4febngA/DbKZsMKgjgU9vbf3WIIVrDVoog7/R1aKNTUFfMX2GHciW7IEtMLtUHPV
UvK2MLMzD9joy9TNk2clAXhNsvRg30h/VYsSpRzR4cUM72vOumiQ9duRFCQ5QZ57
rB6W8WEeO0FXhpH5Q6UGM/N6uV0JoxQVFgop2hCep/amHnER3q5Q0hEkeDE1HG+o
IhYQ32ULTty4Zi/7cAniHZ88ag4HUjfGDIF6VJqrTPO8FyKq6gL4ZSO/pDOm2s9S
LpUJCIVLgoXl49A4LIgHDhY8IXSEz9trNz7QQ4XHYSAWIkN+Cf9KuVOIJ0dyMOck
GrnS90LxtFBzNjFWh7JOQZ58NoMKtCgjvMwNIvuoBmhQDB3q5Hz7u4UcucDGKXAt
KrwP0y6P0uFLQL61lC7YMdx6PUxCiTJaIO6fmrZ/UYS4Rg5XCn/+VKqdhuoA1OiH
7Q6a5rf11nub0PIzJu6kDyh0xPCakZa9OJHmpqdLuftf0Vfr0BZdCwtotfH6h3No
2pfh4iGre6D0CevQ45tGw3VmCpXYFXQawIAAIEbjFZAVwSgv6fgLdZE4WMG/ZpfY
7tqYwvmkrb5gnO6azKbo7t+pMBzP4eL1qM0evl2vzOkUabWQyRsKdtE7kG4LcV3d
a4Jd6R2QyKFrvEfEAPGY/DqhWnP4ME/uf9gSMSiSsnsgjb/TRHtKbKnbsFvHMD41
Wy2j6OFxfNFqJPBJNWMtYSWKbzxVkcAovNng7nTpPmDdZcERuXwHaZcEsVAZA+wl
gv73mA1Ek6CO/prEWm3EBna0aKV2s9TcBV/rr2+Qk/+imO1B9epg2rCN6ybVOlha
F5JzYfvAx5klDlHJIqjPuvGsfq7C/n0rPN4Gl8dXnJUwNluGQX77UWLet1gWcXOs
Qnw3RALxR9OjLMouc12piOFQaO4uj9vPIbG64XsTU2YnrEOG7rfUlWH2LZmYxB/E
OpZfsh+9EIcDhgDYe4S5CdivAMBV57+M5DaqlrYOeed1fwYX/7cqWw8DFvLp/eun
5fz90N8QpCpKGMvUNcAIE8QhL3crfL0CyAONDlurm6o+nXTsByFZig+Aqn+/zlTm
AjNQJn/XnUZA1JA9NgFEQR4CGGmIk6Cov3Uh2bRiAB8VddSk1yl3xPfGwwvV/+gn
U5dMw+reHoCFxF2bfV9ya9YlxksFK2R2A6BEkm1xwf912zRHcgIAI6/pIwatQZ+m
UfbT4/djh6VsY7l/AmX2nYyJy9gSrj6G6jLa9LsPL3vOULO1/AnncdNOkFyafKmw
ByBgDbw5+vEeaMGqaOxl+4HgBPpa8HSFh9bSTU8PltXq1s1Zz0pxePtR6RYdeUJY
x+u9OU05xqUhETFNTLdTqizjTjUxuC5xXhKYwHfdVVs6bZajOgIxR409tKbIKc6D
ucXE+9xyYkSHrXt36eYVRWVsVwyYRAE+4ZOJ90TEkXn6VhIeGdGVdcy2ExOd6++4
H3VBJAF53oAflMBXJK3Me3T41bLQ8fNptKTyVO7K/gdtkOhwLgjtqSuFS40TvXV1
LEnFzktFHKgnkSN6OYKqmEoLxFC4Oz/BjGawRWCT/LQB3/HnixjpchM/qAU+6kMv
oGOnq9xOo1tMFd/n0nfdojji2xnv3wFi1zk5dnGSGvvVTVvcUlRZ7/7zDFOXgfP9
G/JeE1JzLr3CaF6xuoGGCx7HPeS3usUVNmnG/Sqp1YOGPhZAYf/MO7hEb0WLhOhV
L/pF2xMrFK15dst7elEmSkX0+AP9XPBgtxJe1iJTSXYzjCpCei5l4U44OMs8JMjN
YAZ5R/1ZJFuvSHaN583ClPrrVBsXbyUqH3Uhzj36s27AYg+stDvuh0gdrkdIfcjp
9Z0lwBzUNXMH1+hQnJRAce3crwY8f+jMA0XrjjvBFc/P1Fgxqb5o63oASmwbaI0F
UVzRzzxATn7/7OGbrB1IJkRrWvzqnSIpgTKB8XKzraPPfgfsYb4Eh/FuhMxpIALa
9VwHyJfNCpxo/cHWul2HDjyJuu24lXpovI0OmSP5gPdwuRfBazuQ5h7mECCDPLgD
/VpMk2gfWWdDgqFowqTalfGE1beuFfnPnYXyt7vkR6psBUuT9MlealyeEwWj6V/F
B+TTuwjBLRYet4JtcUdoNVoHg9vPYk/3BJC5FsOGUzDYk9ukFIv19XsnN/bPrKUt
Xb3AJEPZ7mbp6eyprZGtXb6IHfPSdbiqI2mDu2HJ8eclSxezNCKu7AsniSIUHCNw
gqe0g0FJVZF2G4NAe8pht18vRULnrC1+iGolUSXU41LJWfgLynwqvNfq2/XhviPT
2Mrs2noMoE12qFCBy5T60EprzIP5E/RsyPlZvs3cYTHZUjlmqKh6to3QyahbVN99
3gtiMX+YiTkPudOHpzJ4m1+h7JIZrWANtApXXF3SoMvDBRPnj9uX5JC6XVcQG3Jl
fv5DXsgCoX2QQKjFcEtxbzrX5yy7mdQIi/GZkdWX8T24JICcXa93fDepBXx6b4vH
lTKL0fQpse6Bz9ysP3Y9Vlje+TkR9TtM7kGjQtxoLadrb8WKGTR+v5sE4tzdQN+B
s9VVHOPi/x1PuwslPciJcKOC5zcKoh8pZkRB7wDPEpu8oziuFcThOs2SNXOMB8u1
YAAGQ+KFlq8kYJwsBWqG1PkBSCNb1WfmTIZ4mm8+EWILz92aBIJPNTXtet/UI7BL
ep5E+2oNWpjXsKasLHUkyr1RFWPuIcwoSCdHy+2/EzA9nAYeOQviHw4pa8aFy1Ch
Qnj2Q0eMhrVbnTBKL+IZQWqZZqxvO7YDTFLBqOdxJIDOPgJoL7ghDxRMEoD/IcBJ
rnjuKM4XU55sijsS941yPbxr9qja00M67RWhDXFXLIHcx1K67XE/yyXVHoxhoEPI
Q+jE1rG/4CjVbcst5tLhoiPVbbm0wM/MlN94B0dSNW69VY+COb1DSOErx131Hjo0
u0PTNMG2FTgz0KYCeVcd6hoJmgo/KJwsv8HM+aLIIgnx8oGA7s0ZQhYz2V8gwyx/
1lFVUTZZNHOMKXFExe+zPQ+XJkJH6GCKTHMI9/5tgsUTGV41fQ6zrXqQAb9NRnuh
1zNZxAHbYD57ClhYE76thsQO5Yb613ibcnaxNhjfbUrll/2YctAe4JkYZ45SduH6
Ed4djlmhW52G9Ku5CSLV3awJRujeLp7BS6m2crNXXQUiP/mcH9p5aIHYWtGupH73
Y2fnVnKr1tSINmoV15FCmqnUip3QGiffXMLv+t5eZsMLsSHXEFJ54W0Iq04lrwBs
SDuEQi+zvrRgPN+E7f/ggzkAzZsWsBxKYYpxjQXKRUnlB6dEUJupkoFq67n2jl2q
mV/oewc6hwVXNlzdnevB1nxTamPImjBkdxjXrDRaeay9VsvgJ1sb3hSY41VvG1Aj
cXahexoJ2pOa4pdi00mrSJHXsk0GqoiO7/YYdvXh9eVgyswESCfAQRmSzOkN093Z
NE/cuYLbCtRM0cfQulvGeJ90V2/sE4I7AlSRgbg/URJubVjR0jitpJ9sIQ0magCM
8sfMgSt2TQxh/B0LDYCBR61VnyoF7zl9TjixudEmitjGrvMpOJJN4876RPK4yJna
iErRI5AY6WfVXozVnClxTWH4gsKTscAPswuTkQwEboa5DbACqGRnaPzugZE8Ov4P
mwM6C8fon3RPlb803k5ZNZSIj/3NpNDbwhPnV4dxKWbj7kBZUh6ueORsA7wTg5d2
Lqnt2IjVwYAGEmjHHBc79iZNsKhsQA9BxBYq66wvKWCM2wSXcVWOt4VFlqjD693W
scQJ2EX3apKE0FFJQcGjAEwhapp/V7XLExD0oSKF1Edy/LXdYWsUHAas1DYgAqmX
WC/XfWcTWapSWMecpaudCj97PkuiotRw8AJYQaVUQok93vsrSKozAyiOsnuNP/EN
KIVzftzMVyRw3g92e1i3ivhdSyTJ+RpJrSxZHLPEfgSCXxxszisv50rqunEvFKua
EYvOGBZ8nNqvKIY4XmcHeDRNSPzW/Sql5ZNhyzM4CrCg6ilnLvvB7/YfltuDmIIe
NaNgB1ADic3gIm2COO/ZCQCJJqSXiJf7TmEE/hPxa2o=
`protect END_PROTECTED
