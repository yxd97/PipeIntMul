`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGNlv5h/5PWfSA05F1K1xIYJX7qLS58N+6MnoiTVPaF8HaZp6K9tJecSfJjukMSm
78/SRA2OqzpwAwzhWteM8D7NBHI6IiRTdVgusDRhhus7w2dAZpMbtrWiqM+tjBw+
0ROMlAUaU41a7upQOTPQRSdxM4pf6WldF4ogopSkssz8zIu/9hirmmjbOWqbB2MZ
IJQAzl1BygzmLOycsM6Dga/fDFP/19Z0eHlZqybJCYr2wfL1bFXEQq4C4utpZK0h
olJ3pVxyaShM/ycutBX87Ek9jSbKRmUivHA0YMjM9WLeR9vnm14OPLWlZGI9IaoW
lt8s03J2Teb5QFk+K4IbSgKGj+GG66G31Qw8px7ZFUGSiblKnO89RwfqMA4dhwRg
Q+rII69Hj1t9/ApSuV/JiAcZyXbD9jkp8ODEw8Wp1DYoqSu9cC1nAap3WwMIl/Cd
Q4TQ/IJ9aweoZ2jS3P25sw1rSMuxGxpc/tai3CJAPTzBhgA6AZUAza8FLGg06wbf
`protect END_PROTECTED
