`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e5AaJMzHevtYqZw+IMzBhJYsGYrUNzZtMxZiOZuai7PXndN5+rvLMcTUooNIE5AH
kwMFl+Z/ut6cohGNUOs4HMkiY2n4F13fvxK6r5mRo08TTuDFRG3p6hHDTWdLP7vw
l0JE5X4Z7KuW2s96PShrYb8b0eCkwrysuMK4WaG0EZjixGSZ++z5koHAItwXAzGs
qOAZf0Xq52wLMjMG44WgTyLCLxskOtAxRavL7v7N7G2P9BHucro9DW1c/MAu811E
U1AFPtVWguD3UPHfEQg0cG3gJscavbQyRWMn0cvizl69lqrp9MiHFxv5Vx01yq26
leHnEsskizHN+SqvSAmRR+1WzdGx3Gfg3eHwhQrDCrSNGyaXarB/G/TiH8dKxsu1
Ggfeq9yZSNn0N9pY6fNuTbYqPzLmHjqxYI7UjsjfBBSQ8RMFqnk1qcuaRVWamd06
uZdpvrlZ9zMCn0DcMqgDqKNQvb/eOQxmogstGoTOIy9Ar5854CsjCo1lx/VI+aRf
rd4A5Hf4BZTr41wsKs1B8wgssOmhHcXrL4ArJbTf9GA=
`protect END_PROTECTED
