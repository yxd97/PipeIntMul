`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dyKE1uXjMXMyCT4Mo/4ingBMcroeiYppiVBBnU5cqT7o5CH1RQjopJt9z17OOD4/
kzY0nhcbjx533XLg7GcElw0FpYz8s/5138dOKveMsmM4erkJgBx9UiYzjdd78X9k
X/wHMBTCeFNDlXBPVKKrqc7QDQjWIf8F+r6wDPizfFFfy3clOeIiYxbjbHgeea4z
OfMPxgNyNv51DzqrTMpK+4H12Nv5R7lu3pmyxMVmoThpSY6EoKBYoAKE/Uwdjpqw
+CUQLEjN/icFLfBNQxBXny+AtOQUYcg/wMsCPehr6+c8XlfoWJL+aD+AnzRPqjo7
AThurLC12i5kYpjYvHLiSvRVxRgh7AzQcSp97vY8u9w7ZjFosY1xcHvg1/AtFzkq
o7Jw0Rpry4KIzgnJYf1Iq1y6IbDpzuuT4eMrLFjXNi2bUegb1RbGwtaZ7BWlskzJ
xQ9AYii86OM2qURvsKhc4qSuoI6vKcm4NS3EXNTPXjKyXbPLuQTlYdexluFm+IGZ
WxYJ5HL9PJ5iiGo+oTcEdqFEsD2xnhCJ03wne2il+RIc6bkETGtU4cgiSVbjinFA
SDkhEIKW5qNZSo1Vw/OyixIxqRAh1cq3vPVRWqw4pWsKqm10ZWoO3GYDem/P8pQA
QmOvDNffxmuExu+idRQUfONFJvoFnUVOOSRtuOW3Bf3w1tBwwE3c3rOVa7vnXjJ+
1le4Rrrmw7zvINrkhcc3pvdejZlnEETEzeDU5YH/NoaWSCiaHtiaXDDixzINE3tF
Cb+sRt5aFsFTKqzI0+ibwTuNR93zGqMfbVM8lfZNhyGJ7SXP03Ba0DJRV/W/IPoW
W+UF1dAZtm16dRZdjz6THFBqorRS4izCmeSJF5Pbd61iSJt7ebwDDavEjJSbn4jr
lJ8G7J1gv+WPUDaE/e/fluLheBKBGJC7KsKYaXVLuo09w4ghFWlXB23u3CIrXFkB
JmFZe3BSdqsnh3mPLtjDTCv1LlclXAZmwuELaZiNNiNkw456Cj/phS8az3McdKEe
cmwUTlFDSz5QbpeIEgakI+5kgmjRRB89IxaM3WQZrrn8qlwFFOlaDuCcrcNtZ1MK
VWRxeSszTZLkW7o6y8MsyrOwH7KN7TV3SrjvaIbn3sbvv7Z6N3X9Q9uvpseFNCl/
hi2t1wylTEU24m3mjZ2QOg7w7eqpmTsVp97jk6Y9NeUx9t3D7CIFGjqV1PwPomvq
+z1zXfSxKTNPNozhwPof/+Ev/AOzJciuWdsNujLSuC1GfLuG0I5KKVW+IFR9tcGz
woQh6QjTSJ21wES5LUO3TB/CBkV08PVC8vtWe2cMu3E=
`protect END_PROTECTED
