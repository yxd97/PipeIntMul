`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VOiEILJh6g2/Ak/acCsdaDYeEzxm18qYLBEM/vRuiQBZucFFxDTfx7/U5lctI2Zb
9/Kl3I35fCtP/UL17/UnUh75KGg6BglkmyYQnJYB2Lt99ACapeFDOMKLzLjrNSlJ
SvlLYx79GW107LrGMiuvxWYe/WefLp8x1Nj3fBQ61afe1f2pt00HcOLT7CdkBAl+
zTdQABkvEc30m+8C0zTa1WJlBD02mMrERpsbJUbYKw+VBDp6eD6SzLSPyDRUziD2
OxCpx9p7vPX4IwuxpNd17JCyetgMNie6FDjc4CTDv8YJtO8rJAPM93R27fylOFbt
KfD1e5PeRvyorX12a+Row+MruxGHEVkn/pOI0UVil90j97gHKLztx/KS7CIzN04v
F7+JW/XeDD7IfgsrNoZlbYp89y1HFtQvCqk3VZ+0Z7dvBn0y6h5iOj+ME+pPocHK
`protect END_PROTECTED
