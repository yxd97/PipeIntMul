`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Woa+VHD8CUg9EahBwlRJk56MLBl78OOP/xTxjHcRHG+kJohnVXIpCDsN3ztgCyeA
Efl5KaKKnINMiORpsRSV2j2GKt9/XaxDanpozRAhogdp9H0lOW4btfWeC5i4SYlI
d6lLmgN81wNCz5I8PSVqk9xs8fMYdA7LUlTqipqdKNXhtemJ1W7yCYw/1PKs6MQR
/5TV0mB77o76JvMyzXrqwp47cYJvMs8Az84Gl8bQpq9ZSQFh+MiSpimemL7Emft1
8Q6eefkNzqgJY77M8wAw5TRUSGDsY3cdZkUWr2MXxpIwdlFG7smJmXznEsmwBl1f
nd5MyqZvPEPy6hjKfAUpyoF7RtyDpnym/ehdjTQWHjsqY6d8zTgZLCa4eJN7DQFZ
+xxC26Nmu0iqk4RCzftDWpHBaHB95aZvtkl7SoGeaVXSYaxqCl1P+ChlO9Lq9otT
A0Q1UGBHNM+6GYwM8N84t19wwKbedXxDAX+kVlPSy9Ror2vXQcg+NcgZkyEB0tkM
MkSeDY4YnDRD3dBfx/S5mcqJyfoHXPWAc+qSLC+mQHNj8FqBrutt4U8imOuwH77L
0761amfcG9p8M2UhzzgXOJzq6adIzfG0xYpIMcmBvbI2PJsGzaGUC8AEXE5NNeOY
pYhE43IPkl3mseN8YbUHUGPBiEBLyYH8sGAumB6TKsvV/cuqI4tW5b4v8cRfxjWT
8CNvOuwJY1DdFBm9FNbg1taRwGnPOVcMmlIV3A9WpvFTW/cRREfeki53CITynaYi
U9+I4q9VZGyTCDF8BsAoSqhKzIV6XZq9YlGlqHrSG0t7jCGDWEX9EChvfzD80tTX
wLbBbhr93nCeqylsVI76Pt4OacttnRRJHCpNP5jwezhVAOhnW0X6HNfJ1HfdvaMp
wxmtlX8JSNV8x2YdNT057mVagcWPiR1BRBO68Ne3AM9hlo+md/Qd118yFjpumqcb
nVoXu0HofcYpSPT7dGSobwghEYHC1DSpfuLf9y2oBFZc7FLAAEEoI8aYZayM+MWO
eCtRBSliVpTz5kr7mBQwrSW3gX3Nls7Gp/fALndth7QLhE75VyQXJ7AigoBZ0Z97
664E2jPfiwJ5TSZV5BW+hxPcWNgHir4sDHt6Yzewq2mljJ3LuBGI+fqK4GqKsu0x
uPGrmMmWf2N21AVWriegYwr6U31qy6ACQDE4XL0Xkv0eO0GU/KLF9LbKk7K0mgiP
z/McESgAIBOec506yUeD95LXBrgGNC8ZHxBAUkgO7f6lhYkEK/5S8RB455leTG4B
asTCToD4GAiCSqdfrCfVs9Vy1XEZWqbuowf0m9Rl0DNgCvJiwlNOGD745rhM7Q+Q
vTwzIEXmrtwWb9sKrCrMQowgoqELaYngU6oRgvGkHzB/1Im86hPd+djomvoHSE4/
AtkZP8w+d2STFlLQ23R4YrivjQS80vBNydWCCvoykfmJte2rbu+VF/U2X472KhXP
uk19OOM5WMmBOLzLrENl/OKwVQ/P+QcNVwqfjhHi2/0=
`protect END_PROTECTED
