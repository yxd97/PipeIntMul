`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fS3nvLgoomQ9EQMcicI2bMIptnATRGBabXrKqiMJAKozXXt6KRjXI5VZurAShp/Z
JPDxuOR2wGDKhRVMf4uutJaf//jOmrdJRVZ+ENLVvWhgwwlb6V4Uq2ypNPLLkm2R
6ZYHj2kvUByHQC3KlTpRSS+87a1XhKNTCPGsU3FvioLj/lBlmJoxnugOgC/RzZK8
gmBSQvXJEm2difp2vQt+xvxZX12FfMWI0+aGeukBNw9OfZMJ4wlNUwz4xikrj2Li
dgtrAoQeBLXaCjmTk6AqEXcPEdNeczOF3gQzOBQNvG/u73ZTY6z4SaacbY3UZrEq
phc8ZObrxY1CPMlS/mI8j1J7R7A4Y1qVWt5f3caIWd3AxFPsR5FECbMzxhuVU2VB
sEYuJWRlgsD7Lwa28rGBmXdsStDVkD8sLpI+AT789/Ahxh9swYJH208GD7wr1B+7
tNiPe20Orcg7H7PD0QWrcEis7/M38yCkr9E4q+ZDKPRXTHvVolCrndlCQc6tQkZD
`protect END_PROTECTED
