`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eorYFxITAVO1irFdxKgoXlDfZRNxQBnIp7/Bo+6UU4uAemR+NenZHKWcRXjSWuZ
xIWqsjVWXgfsMy/QvjtzdpQQALdrM56gaXjlwiJqrE8D/Xmxd0Lg3uUkPDWAg/xt
tOjIQdHfQr/l6dEIzqePODuhroWuGCuJOVpT57vtRnjXmiN2YaztE8bYJsYldNoy
x7jIIDhtgTrMNRaQ9qwB4Fy6Kp60IOgREhb6c+AbRDuGxzg56kOznZUZ777bZSYA
OBIP0aujNTAP0xkRauNfKOiVzikvRdfEHcTVqGh0E06LlolpcO1t+d2g51CO7U+2
+dAve2UDf56DD1C4RRlBtRAWP0qBzoK+Ic5MLjq9gkIlBlqGSI/Oiyadw/vaenVX
QY+NX4EkkXddTN7QfU96WMBB/BmVzLn2Bjh/EWDSsd1XBF9enodUXBhQLhVy6Y4x
jj4wqwA0Lq63K7uH5ij1zii/nTEECp42C23vNLzI8DUa8iZ2+uNIIUm2ySDQxFeY
0btessvhQ56zsn9rf3tjg1csp1XsEFzUGOhzZrCNB/KWAw8PCJY4oehN5vnT0/Hf
6asvJZSMTS9kB5fy+RBsBa7HLfQG6IlP0eaS2sTCBGSt2rdqQN1smY0TU8bj1eBg
nGEExL6sZ98nZoaAdV3vmLRrfahdm8sO9FxFLUcRcXTyjFxrnxM/HbmqQx+XJrpu
asZSqC1qBzKUPiNtZxuqx+6esyPFqLKTqWI9gcg6KLrFT+56oEQWSi2O7HHWXEA9
6W1zXPhE5Rt+ptQqXYmwBjukm9uMqHC4zua6/sU0q5peeSoAsYVz1+hgdcvVHqN7
gYMVsEYCnJyi6mB2xgf4XErMOr/h+RNCQIYMs0Mp2i0RY+bk4klLCQ6G9kwMaRcW
Y68M861Vkl9keaa3AIRR7xIl9UwnywbSH6Ixx2Ubt2VcOcLAk/wNm7JOUGoATfrw
/EcvG0aBpU773IvpQ06+fmvBR12sxLBlxlEWgiXSpQ+HAF0cjN4p5JFN23rWxSEw
h4X4EDJpq82qIocE0Rsdiw9OxXZwC8Gn+LTtKHutKgs+MSL4OpHqUecZvAeFephp
zm30A/x7hUocI8liqVz5x6Db/KMVw23qaDiB0rgUPygXBnjl9EExu2qaR19UwcG4
8Hzvma7QCktkh6lOJbncQLPYjsvgt+7QgFfaH3ZPnfSa5AdwaCnFP3Sya7iKztFO
E8LAgVRH7wDWayMnCaFOcnA/RF45uoXYzu/fLIWSQ0pCTQULZwEMgutclTcSB2fr
8XZn9d4vYClXUK5mPfpI8AXpH5QcKszQcM1RqrjJ7Gvs3AYpzoN2vJ1YuTnoJXFN
UZ+C7fCG86FkGZYyHY6U/zWxEjRyxzBc897UerFuFK/oyNyFh7fBHo2jwYtmJ1Ii
zCW13ilnjRHefFgnnM+Kzh/u8mnuREf5xlKj1Q4JbJeDvDBK6hZzCSJvS9qN/l/f
p0QNFll40/dbxTBuE7kw+Kq0lnlKyrj0lY4lULhIPqqy004gXosYOIiQzOvI+vU6
cPU9pBmp/wOct8j0jTSfpZHxV7vaBHCdz/qpWTQxZdcZDifl7n/GhLVchJAvley6
ZOFS0As4CNCSkIlRB++KJgeIMqvo2JYTasMoTBCh4S36SFpQmHgMIbiWstg8JSmT
W5vz0z99DOcTULQm2+1o4A41w54dNuONHM5kB50SO+aCTq4syQ0jt///CRM2z8SK
KTsHm6leeIPVJ1BsGG37OxL7QYTBwpB1BwgEfIO1YCC9sHvr54K12uKRK8RfQBUs
80KyDamTFp1gPjibBF/ml0iE3c8zDDl1ylLpVQsk8CMhS6fake2ry8G8jYvhrF2P
ret9z81huEYzJLu8hW6JgaHbM+h2zOGeKmnVl1hl6Z0bhgaNxlt7+hW+7Y5xR5Gz
BGCQKXX2mxJJcjU2WlXi4XKKlzFsiJfQ2pinwCS5BjaxBKBK6Rut6ZDHFR6hXk+m
rBuAu8hPO742z5Pa9ss9bxrF08eQvTSlrZgiXlDyiWGmRrbah01ieuA7MWMDdhpw
q51bOwt00ewaJ+4MrGH9Dm455qm2hTdWn3/nqheldy6v4mdem/FvTh/xKzdPz/a9
xqQS+P2hTjaoPBRaOvih0L5TWKRGxsoIhBR81K5fbf/GOm0T8VNuhU4kayaHWOlH
d5hCl9icLHTC4Er2XfR8PdfNnpMAZ+sloJJ3nPpCqBxr+FmIac4pISyq2uGaXMNT
vGlZLJEgbVx+t2DXv4s6Ra4XKzWrXRxMlpw9PNo7zxrtyBckFCBlfAH+8e8Az/Sf
`protect END_PROTECTED
