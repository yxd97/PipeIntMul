`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKqIrAN4sFt279PNE+vrqGDtvT0dPcQnZ2H138TZiDiTI+Nrj+CaEZ+3FCDokDZP
5kcAqXT/N9mTA/arshfFfprCEGerJHsd9XH+S6QA9clVmnoDkB7gEOEPiGbOAgBq
cMuJqLwx34jjMaMo+skfD1u9p4ZfUTj3swft3jfrBfrNIeJbTvsR55TQ8rHZoJkD
YxB9mPrTDbaZeel50aoV6jQ1NohcWMQo0PrpRHFRRf5sjND/alawUSHQ+nwzDPxN
DO9Cberp73YlomXY7rI4ITkNBjgJYiFq3i8lVFz3VeDLsAhM0P4v06A1Q1kXfHPy
7P9VgYTuMbVkhQxIHcEOhJMQE2lQRji+oSDQlcD++6683KknS9HL8Z3BNVeKHSj4
fciKOIKKJ3DyCMQ2AsPN5VCiP3iX7ABwdsxfz9844/gUA2NU5usH2If73uSse5Cz
Tc8fP97sz0JR1gqUg37f+qQlDmcGdGQW3225CKrwOCc=
`protect END_PROTECTED
