`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UF3QuVZgM3mLD1PCOpPWzrlqFocPQUFsn4mbvIi/siB1g9LZGs44ZkAse2y/EtUS
0xDVn/H93Fn2K1WUFffxTtS3bXCxAKHZGEtm1g5M3EEWo5ZbZqcsTJqBjYhcgIQV
zdbNFaOCyGFE6LZVsZ1xGL4gs8zpDC0Caoe1GreCfssua4E3zJWH7b83vBw33HVK
I8yw5UJY4MJuWy8w0kwDSvN9U7VDVlggVSMt4Fmtlqb+Kk0s/Fkbl7a/NQ2NuyMZ
eA/9URFkyNO4EfERm8RjL2iEq0LJu90p2KdItGfjF9+VmOU1C75qw8FOEodziCr4
ndRIQamyE6kS/+OKh5+AWLonpORM0V4U4/WgAcu7YOzu6vUVj7QzmBuoNMFRm/sK
cWLla6s+2jPgYsUAU1Ji8UTjFvbEs3IQDRWOkFQBCdgp9UqdoGzfonyE4Pvj9koD
r7PO6AQ8Di+s/1rrwb26jH72SgcXAY4GhKPS73wXK4/EPFfgKG+YwJdM390gsE1a
5TV8gWahvh62VHBtakiY6IqDmnkhzU99AfMGM0JXqSbNZTlRYk4+pcEemO17Dtn+
8G0U2U5gYOwM1rVZZCajkdx4kRfhyOu+DhFcRPolNDbw5397Eg3QOn9iv1Vo0wqn
HATNdROs5VPzOd8EnFx20814TgSKDWqWhERldIQRrs6ghrGqD2TBOir8PPA3bkK7
7R8Be/NIOBaFBbOHyGkMc34kxX4bVKLJ8tP7k8OUHPoEUpDPlKOWz0wePzaSQUJu
YZL4G6kezee/zLZ1q/azPTr7JZi0BQig+PQhoey3NGEhlWA29UrDHXzIj1jl7AII
3Nt0xlPhhOQdo0U/d5Okj1iw2n7W7m6lAgrmjaBQT6R8EgqDf+Kq7KgGpFw60s9g
vcEl0RQRb0tVQVPah58TpZryGZtPb8boFINEXtL8zQLlzhAAmzmylyPkdKMjzmtq
IGmDpL8T8u/MbuBuR2lnesC8iCv1YD04e3KLQ2I93oo108fcOKbIqe2hFh/7gt8+
Kg3x3LlskMjch7sEvZiOupzgEGM3nCY8IqRKL8/jXHdJXd+pTCjuPjGd34funUAj
ao12aazek8RWqmdk0UVZwOUNTSX8Gxv4d6Oec/xLxoF8N/JxP16ERCYu9ZOmnksv
C7kVTH8KwdmniZ/GfjmmGT3SODk4p+fKBif8ZS51oWFxInKBJh/TqPrtivTbHUVz
mA8RuwtO7v+i5lGnsbpCxhVEf8VgDsM7ZhZQCZU6wpkK+jbudC3IkfdxoLBczEUl
`protect END_PROTECTED
