`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Anu+b8+SWDMbCI7an9rRt2ZMHkC/qt+5KRmV+KB0qLj0ZLa3wdr1q/o1oeU0wcx8
mNVY5qKhG32yMGv3qLMerflNkCqLoIM/Gv7oqBRsXO3Tt3nTIIUTmD8ALswvcOaW
0A9uuWss7LCOleHjvbJrRoag+YnD5zZuUqdouzBK5uQulP/I1FgKeTZuceTkTXaM
xZBnwbEj9gpy4Pw3Doc/gpZs0nszgbpfBX5btAr/BNobYbjjE2Ixnn8K782+R1YV
tQYhdxqiIZIGsn7OMRgeMOnDAjkyLbLQpikwdjBwAhS4Tu5bSu7J+2fKEPUmFTXk
6NuFMzJVTfTYivedudJ4wZisTVCgqWIgL+9LLywvlZheBNPyOPLghZIUVNiZHVCp
Ye6Gd7FtsnNKy18v4izkQKmXCwPhnk1DNW08TNUrd8ASlHrekSHP4Gdrd2HJB8xa
JUyMYtngSGOxgIstniI1nK1aVI1sk6gwgdVEl/rabP/6Jykt6MWHb0sXilPVGaB6
6+kUzcPrzawIeCzIKPiUREl5IbAAvfV20wOeTbJwICwif1bhrw+zA8P2lSK6BzaL
4vhMtUTQZ6xUBy/E5GCFlg==
`protect END_PROTECTED
