`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6Z4nyJwdl/BvlSX4olgAWbPtM3tnAsI/1zZc7pwFObJvv9We4cBGmKa4uLGEOVS
XnaoRDvWgczlrx3b8cYdi2WBidBVLmncqjy0hg0DdiTJKKc0aJPf+/LpMHmk/0vn
z5rL6IGyKxUbfnORDyTR0U5C0/WiIbGSIjx+SkaKITVO7bGCwukHNew6o3iO8I4C
8GF7e3dznlQk/Jr2EYs2ZgrMuh0Uwr0CB1Aess5Pr1UhnuAHkFLyJJNgUbUqlgQz
oXVNanSwSTsaL0KSYa/yRQ+PKyLlDdmE2GFC6E5GdbEqgmkX+OxAJew15COnNA00
Ix88mCL0ZqBgjw0dLJWqvFrKvQJBIt07nuTKmh/+PojZoYzzomvlm2f0+WWHM9lT
PHgKfLwcOkZsG/xUCV8LGwXIvzNAEhCGd9a52VHQZm63s57C1n83zcYaextXHOF5
kTSTXP/Z34jRo89upynqRsIWsSgTiE7lD6P5/8MEFrZ6imRJDkf4fOTDSWIKVoTc
`protect END_PROTECTED
