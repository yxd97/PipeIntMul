`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tPoRtIzGtJ2y/ZW39ZUY01kkB0GyeBSf40Vz4c8dn3i0T+2/OeWC37gNXGx/qyCS
Vq3mwO0O7FaKP84L0ASX60G62us49zJ1q8aSsO3D3c/Ub0EGhBknUmmXdbyUZQc6
wm9+yfV7wL3DXkoTPp1Dn/uKEnWnAYMArh9odIB1nT3wL72LglGqjg32uj+rLV9I
ffXd9uvV9/sowL+hBUKFEHNh7hL0XgfAcr0udXxIWjyA7a7vTQqVpuNCL2X3MPFb
KQ6JFT0XipqU5v+dNL4hsrx5bkJaR6v0vyWv9hggl6lrJ9/kohDIywwXk+GW/v4O
h2FFLd67Q3hqcnFBnGVDKcpKxUd5wm6CugvfFSkaPta+YSxfFTpwTn6XITPgow6V
itKoX76nPXnw2C8HRy5qZHsxw/sdG/nehZMVjmPo/n6n+HdnFUmj3AxvSTWToHwQ
7Eoaz32ySYc2cLnAtf3zTjsq/f+MPHZoo7N3htcYGrZwnarv7MDFj4LgYm05pXBd
NJRKBviZkDLVb0D0X6B5BPSsJWZZeGOixGBJbNV2PM9DlrLNkgFQLN+Ikd9PM24S
`protect END_PROTECTED
