`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+09MXyPeiY5zF7ut1lS9ivRtxmkeMpvVLj/Z8YF8NarGq6yMPqRsl1rRpqQgNwX
K/+/z6yi5UUzAdHootNMJjOY1bjczp802euqmuccx2jOBVsvn9FeCkRLRyM1svv6
Yjvj8EEVhBtVNCKNd8qXWZpkDmiqAsJ4qoi09fBI322x7JCOph3J3RdWXpSxnflQ
V0SEsFFeXnmAuw3aJ6ZMAdyY0WDuEK0Bf9WWSfDlTo3ZDN9ibrr2yLhFTtgnZwVl
T2Cn0zJZ/UiA9JTCzUIsvw==
`protect END_PROTECTED
