`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYUM3Whgrn8H/9RU8fEgJ9zUQLcPVQfDQFhTmgJGj0LnmGbmryfOSGtq9COIp1q8
MD+Po32P1TtZ/RkVe0vIIX5QrDcTbqaOLyX2JyC8JzMLT6x0L/QlXvgkkjpgmXV6
K26B2Qad4Agj9V6OX0DKV9pSVqDbRpzKOavPM99mlVrRLFxmHZoBE6qm5NNyxgK+
/eT1I/3l08O9SeYrP6ezoTxd8XiL+qpKdrXFTunrwBASrL1UxTecJO5kiFaq7AKO
WJycNaPDSRS5frI6xjG0w2tBzOOIb+gf2eBYq059PPLWWZt7Dg4JasFvV7qrL63N
EDieWkJCUatW5ZtXxaSL+vvj1HaPrLsxneOxJBlC2sJU3e6DWLmAEvAlKIENw9Mo
UbeIBix1IMSY4ud2CwnGcuee0/6WM/kAg3l5VKGe9yzxxgKWRwf/NAabKgwxwsPV
`protect END_PROTECTED
