`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+L3epLjUs27Uo6871A99GUVPgf3woGbZISz2LqQbX/Y97ErJy6t/YdEElLrqVsfy
iTDoCCm8AMvvjPIvyyCqfOlMhTY7ck6IHofZvvaPjdzO48QCHHTK/vqkxxYdVVPg
Aq8otQk1g6VW4hR5bGDz2dli796O8e1U4BdnYWdfnZAx/UFL9Tj/sgoKqttmFJod
lc3nQs6B+qK0puNbBRsr/frfSO/PjshC7aDI11zi47pxRpeDjWev4cRdcF6YqjNe
ncTGlurSaEkP/8q1Z0SotFV7SqHW24k7H67KfpLNaVLc+GVG4Ddl2XQPLBNXgp5F
na6vU3TCTAdlZ6XufYdJKQDjvdtc01UCRk9EKD6csoQdOLOna9egseHKDToRpI5f
3rRtezVLuU7YDDtlj858fU9kf2JuDfWMBk+QkmugROEQXS8UI5WWbeLGkyu2YZ9M
rODBpeOCKNvOtxh6RRfV3IOiIocscAY5i5RQOlop66oPisOuAEVZmGgXfTW+f+Wj
+6zFnpTbAhRqppIHB08QO07XmJysGo+L6plXUPoH8lEdfxUDapCSn9v1IvgfOt6O
jPAYa9VT5TZeOaRsGV8pWp0YiKgotVaOP02AgklYV5kipi24h7k8qA5g2Cu9Fi1x
PXe7IViRwk8ymGrvaleo4lS+anCBb60IWSmXcjZqRRz6q0M22FXgx9IO6YwN+Dcz
Gy9uGyVk9a+Rkoy6OIk5hKoOAbCbEx44h6Mla+Bby4hRZyBWq0zjTw6640Qzn7F9
PqqC5j/aAXut13ZvZnwybC2lnDg56AuG8abuiGJSAcQ=
`protect END_PROTECTED
