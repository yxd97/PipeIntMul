`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+mZSJw0xl3/CrYea37fiuHdzEA/QAgF/j2EkYyY2YBXwaMDF1UyrJrjDx6OkDtW
8h9WQO/5IceJ2irp/nxCV4Vwr9Ub4kNwic9+A+vJ94EYcqqr6RR4IeOvtRxsivYZ
m7JaEPsrjbBQHD10EhmwI62ZwT28mnMWcsOCcJ3lgUZoXgaFUyu31t6jrKBegEWC
UVLW9JI9xORP3kdRxXKcRnPMA8oCbfxiUIsg9pgqCaTvoesHg35vA+a+3+hfdKL9
dTmxYCAY+WWdY7aHv3eNA0+/7J7nhChEOEOxWUCfSNehgK4Hfa5YrI9B0SJfxyun
mMf3qZ++QHTo6rZP1F7HnCnS6K5EXLgPdxxg49VyrjasBEEXRvvyIU4mFz6pmS1V
p+01dR6YQjj8Atgv2ErGSe4ci0Qp/Up6YyCOPg1Um5pr000wEdbKW/gm5xgLX75s
3wNeiMnEMAGBLJJdoAp4hJivIEB2LrNVGwZzJAGuoTcx4q9Qwm/VpwZyQyCrldz3
Viandne2nhbdG9b8xrhTPeIh+e40b26f+EtP3GPPvxGzISQSYFgrJx9b1fUrHLqS
yZxhu0sbk7biLQxU53CUi+LjTko3ERZBnhiNrhh53J7ihxgq06Bif0c5FPyVlGVV
L7QgQpqrDVXsYI9VTtIxdtd49Fn+w37FUEEmBalSgmbIXbxyIl/HvxSLbeij7Zn0
U/dEiTqG2R/J6xUHWcx6VZb0Fth8uBOjVS0R2YUuXvgGJqzksCS8CXGOOsIrR33f
`protect END_PROTECTED
