`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxsnzR8Why1KnpgoUdSoBOIHjDik9VHGYeK5zvkmhgmawGvrqIB6rDmSqh3Ae+hp
V3eNXbI0XgDDgFf8guXHeOfusivBTsuMAYjzDHY67HNiJn0vgg3ij8JjaGIO0GOt
eu512Ei4ZxexfZoez2a8PtEuLd85h4JCq44xBqnl5IAmeDZD7aFj5FhQ0TocHKHp
ybYSGBRk8RghiQfzwsoOhzDEnrn2aO8sPHehQEDLDJ5STQkn23JfWs2jHCLEOCTP
1N3EIM7P0LjI63JbJXZM3otMGP1RSKe95ZGKR7W0quYXJUs9nB/7k4wA2/mGqCr2
vRdZuNIq8y0xyyjfhiS6Zdu7N8uiVteftzt22pcMIZdwdDKLNR9YoTAC2+jrphru
XuWELkuW47R9/JEGBAjviop65tHm/Ek8S69YyhnGH+wAI1cf8qKrhKnivI/ayvi8
ksNaGCl/k048ewUK+OCPcwaJWZVlfz0E+/iAw9eMUYl1eh3YWkqOkiPSY2wOn+0D
xBC3PXrzWz71wdFgPfrrLK9hqcMe/BiOrbmKLe8+U7T0qsdOStOWgVipwaIcea7M
65womgR0HVKGPvX5xpapf1TdJwZgAlhCYB1X9nD9VxG8lDY3bEgDTQO712ErDuwG
ZKhhhmPOL8SLo51QHpBWHA==
`protect END_PROTECTED
