`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p0nq5FURo+k/rLwWUEursILvMRtj2de/T+wPnKG3lpqdKIbur2pKTANevmvGm1iI
6CABYQqYrcaoXeIb5BLvDpZaa/86QWmVs11a1i0N5Df/YRHWqW+zd22ZYoCCC9t7
1K/joP/EL+Uq9KCAMKAZVq5i1MVn9iANJYGz1qJXiiu+oLb9jlSVykdz30hXeP5R
VkmVkLjy8GHMGyPUjabiL0MBULUSp73WqcVczavfEHrammu69qBvFblm9vwl1NHw
2YDDmzSRuGwLLl7yCMRKF+zmtq1qT/KavP3VoVjgLg8=
`protect END_PROTECTED
