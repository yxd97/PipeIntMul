`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2vdFVNvl7hIvuOpWRndm/o7DSWW/cHbtuogiDbmRifxzrSQbL70hULdKLfxtXSeC
mvlhLYaHnksjEFreX47WE9WaYHJTwHoHesSWJ9SpF8T4p1seOiDbFNBzoOC80bU0
iiN0X76nUflsvct9WTRvVdbJIAOLXyVoa7Vn71nVKk9wuL2+5rj39gBTuQpEXIPg
3V0xnfezZoTOeGCXliYdA8lR2HKE0i7CLbECri8jfeMtMQ+JMVid7RqrXCHLk2GP
HroRHePkoc9gfHGOAc3eUj6XfYUeLJguBdrVUH7ez8fqsM2Eurh5JZr0A7K5PyQ5
nK4PTge9sTYP5I4iXaE3EW2saQ+7ZVsrrGXQx7b6wRP7eNNei0SiQn6ZE9Xd1ruA
6oqyL1ZKYnSXhMie/XZ5yLGQZbGAZATUji31oBI8mHjNDwNUq0K/gSTEW41SUeoi
CKne6LqUiHvz901BTCgXI2ts7syXRVNhpTZ6NQycFojw/Vyi/7+8xOAdzchU9Kh7
WWNQ+WTCXjVzMF/zPaoyqsdbWnUP8hIFVKb4Ryq8xOgnrPSs7suAcZbjW9OCJnSV
ZUNY2z3dvGLiQzN5UJMhDw==
`protect END_PROTECTED
