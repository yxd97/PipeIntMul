`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IljVhLb0JzaSfMhSF8geF+h42OvxxgAy0pmjsk+oRha7j45eRKPLXJofKXaqwJY7
58pUKKin3pBetA2ViFtiqQX9ToPmSg+cTJto4/Vr7RwEe1kIHgIrssYwKr2+P8re
NQpyXSenxsiX1mHO0eJIW57Mv3h85WvkYonl5JN64Q4JWed8PYyvvRIkxK6orl5Z
auePYOQMR++vddvk55CWdMcAYRHhgnZh6bgUlNEpdrzw4tflqB68v+lb950vKE6r
rT0piF/KXH9+t3Gg/KCvHZsCBl8SXPH4kjpaCKPTUgYN6uubwhJns3PzE9XtEIz6
Y3tFZ2jGz1hD8RPHj4/60qWfF6txCpecwkPT8viV++HZjavlcKppu76bl1BEcViA
LuGpvaeO9sTalUA4j+CcYzCUiuGIfMFFIqe94Pfy9QCIl20OAVkwHFWBZX9l9Bqm
1hhtahYn5M6DXTcTxLiMeVSXe8laLBo8gUM+hWGBr2tqLQdrVnGSbWWFVin0Pv73
u5KtV/ND0dJkslDCGS6zMetVSJEMGky6EiJXwknGWPZXxqmog9sENDUOfaS8oHkz
NlAXRPxfAODoxHgbVsXoL4W8DQ2bhVcP00bwQHE/P2GlWPsvQL5W95iep6cuwNPU
AcZF8Yio+bJe2+u1zo2Xvkjf8XztmJSOUUAJINWuoxKBDemMekkBDS4Psa1svMft
822gA0dm1bbsxN3kiMBukjMLZ2xg7pSn9rJelEEUuoUfgyIeKii4DNp3PzRrEUHE
rlsIlaRtD63BgXpv5gobDioie2lKmLaHH2/lh4KQ2NaieSJ8FhjOj4tfYXhBgepK
Po24Acz+fiWi3RbgSFfQHylyjiAXyNdNC0a5OCTplzRMqSi4VNxsIIkjQcnprzV3
qinSU56jHsuWde5Q13AVLkFJi4Cib4wbIDCegZNEt/cB0DFb8hpDXSSfpL2+5IV2
EuwFPmV10HILRsL8PzKhzhT98cPU7FKiNExk1MrmlHW191K9myXSHPx7iPV8yUwV
qx0dvByfrYKGqfTPBgVKGpFzMTryGijO1KBjjbqG86eJ5yNWbUyji2zpm4A1tL3V
bsiolrml1Cy6dGbtMKNkyb3sdnUqHpPcliW1ipZ86sBwPaA9IyGORuNEeJSv7DxG
+A4a3jahvQ311iuLjuBJHlLr09Q2hUlxKe2D7kYCeXTYvrd/Y5G8HY+mdMXhzz8b
f3ebuMtt8fmPBkzT74ldtv4XEAgKnr8A52Rh7JhG+6M31JrOzkq+kwgu7rxQS4/v
BAAyodrVULjTzLc3SVCLFragoIjPmbn6iEADGiKiJbymzMYyF8um5BVEp+cGBfjD
B2u61V39u7h2aP6Ro/QdnVbprFD/Jp47ORo3kvK+Ja5tszuHNCGRYs8HGqYDnjF+
Iw/QpuidEQCcU6IMn+U7GnYO4uVS08esO68RXDxNTYkA7q7cHjmb0a1BARkz8JRQ
bMqSEiFbJUGPDzmfzcklK7ClDwsJsx2CzV9lTl3Zpfu//IgYbf6WzzL9tsW/shiv
jJNLQxXfZUE8XfFqXkwCo/507uHFeE0yizZUnc57ZgPwOvbja6AVkaCyFLbv4DJf
Uq9u99nMMlzNyL3O4QXFVgGv2rowZEX05pUdb20exV2oOlgtu4CGqStrmr7460k4
klJDiQUJqsCHTwTWhrjFs/Z2Wl94vdAgA78CHq+82eM2yxUTkZQeLcgZA36+etZ3
VSsxc0U1yCF0XPvwDUCiV5VVQya4uBVy1XNjDyW6GMoINwtHmgCAtWSb4QR1k9wK
cMfF8v3IdfeRhzP1pYF+YH4t8bm3w15ZxQGc9LXPc5xsEKzQU0poi4ivmQuV9LL+
hMSn8Qiyd8oH+ZlaXvWgfeXp2wWPIBZOEF/JL5N/UP88U44x9/MdZItRsJhQYQZz
4WUv7CtlDl99VgHf6MiuKVojUPRo/6a2rpfgXZrb0m0dhp6fX9+FgCuxRyuuGKHN
9GqxDvVMgJU2i0kZq9iUuonE/yiSRo2lNKQvcORZjxjywMdQR2KsaM58VapZxZt0
xz8QrrV4qdi84neGxjzl21k3+oy7V1hMXP5wnasLR0iEZocGzF2hdj5WB/V0i0qX
hrH2fpmTlXuztaC8LDCaCTms2zXakICgiUBQmnUV3S4eG6hYkYtbID1hlGhV8Czr
m7aW5QRXFCwQwB5ViXixEcWDaK7saTHAi7FV2YjmmV3VciyjFTrpMTBcZtd1ehSQ
Y8mas2q1bFI2pvidoCB1VbdDbCtFsmz44lD4hxVSaVdoYpYKrypxielipC9kOVF1
rRwumMRpmOtMst0Yg+I4FcyeagHWGmBOW9pb1txDIF/ORwV61M9X/94jhndqpUas
5vKdEUapHlu4nNLRKfp2NhNrsjAI98t5qUjbd3LMyYkXq/MEyJENAiWGByMOMyPI
CBnKkPYkVmSsAoAjzzOLqowGsb3nQsloawCr1blY9jbN4tv0McwE86fZ+n/CXgjW
E257vq3V74ao0HtmJs14brZl0ucRcBZOvo4Sweh5Thq6b99EDPc+cBBuKSWTciPd
aKrStjheD1B9fAvBJo00up08g0EcXxbYiDy0VYjX11zUXD0R2XKtRCtm1gU4R8uG
QnsBBjbj0/IkeMg4dciN1gaBVEDenmrGMp2nZrCF4o/MOEufEWSIW1iFmmhY7Ict
ZuFb4z6OfsiXrhHa8qF/YKQo5pOvs8WGXHRKvp83lae5Rre490xI1c/gYtGi10je
SOtTNK3n+4P7NwSwIguANB1Y3Wur/+NVAd7eZD+AUXv69CrJ4335Mu2IGHXyHUse
BVsqprmgTlRohcdoDIDBT59mzrvTWZo0soU8LeeVKianNQVoXVYc+GAbKMnYOhAF
1jFS8XASQyEwEPZBUC2DQH0NtUhuDiK8kTHtDvBMGC0NhaWl3dWAWCKzEPG0iNd/
uomzCc1HqoURmC3t7yKVyz5U6iy4Cg1qTiHvr8KcJXbkdtR4AibcGN0+mSz/FIPm
Yc5ixJNwE3CbBAsmMQ67/9cmOUZkYQ30VPNSHdngLO4rWUB1hXYRoZNjtBRWJESK
96MN5t3F+FcIv9wBPRh3aYY2EXQsS6MeslyGgzZnwXnLfx+TGVTv0vOrjGTTyRhq
Tf9DdCWQ74wrDPSpxm2XODG6pHL0P2oNZCVjjqFTF2aXdcn3RwMbVWH0EfPtzzNb
h+RCPGy4QIDObk+hUE4jAnDBfPfSYcLpiKl7phbmRl2HqS/dq8Tdk9Pz+KdPt3YN
LDtshDLx2KICJPIM9TMuPoFR2YJeyHlYFOSYo4RlCKu7s7E6b4lkoFvEGkjg+32s
5XFDgRPFlkCjk42hkocW8BW0gDq9AaXFcwXwl8hl45t1drlO5OsbxWT1ioLjkrD+
XNDhikaKQbFjSlkMoztYNmNDDi7eLKouyOfnfzdaT+jkXt7TyhhgBUzfCMXGs6tv
EEv8RhEZ/uVTqZJ8sC590uk6n0CCaTNzfzXVnSshTNsCpedjEOSKLFN9Y+xLKK2L
6TXXdXHlImsHx+To3SCfv7RpH4OoR4mNylcfd5xemfEX36rkvpK7vHT/FSJl4soq
xTgkxmPBSraikpqJh/66cet8zVbpxQzSRuZnT1oVBu0XP3Pv5JvcU1UCAlV/nkGJ
li4FCBpxT3IQk1NOYLrEklIaR89Z7oEzOwt1A/p2amR4Lz+iAE92EsIsx9bJTKgr
VRdVTYD4hWTXaBF5d/CN94vC70fKa5QapVacTrMvKO2NT7kdKiq5if3n+eLlaGdM
z/TZhcbaK9hbriSJiWMftN3/FstwNRwhW8NeY/XNW0XSJrFt8OXuripwFECOpI8I
cKQ/qgvrKYmrq9qg4KFSWOcaow9ZeqAslxfh96DaKjWDBmHR2boRoceENviNBoH3
Tr1lxk4jRAW5A9FJUr8wB+V9k8TjtjHN3n6JLSnSN6JEXE90Y+ts2/nqawRKxJ/G
EYdHAYbgMwUeIy44PpnWJ7uzLe83e2fyNjBJwxllXJswh6zEwsDzPGp0g+uitt2h
7GYdyoTNqGJO1sU+pxMVLinbm5tMmHZK0g3b9+CK6kN+9YBIRIisOipn2GfGI5FU
1wGh5AH73AbHxTkSqHrDzvrbxgH3lSOq3SdeI44XCsb8PKf0nqVLBtYxC3qE0XK6
QAeg3yd+J1UNsN/INka0U7QhHQ90ul2y2H0tIKvGp/BmB0aqDF8795T318XvIjc0
ft1O6ftcrifnPlbx7kYiUthTOgSNe1c5EKTbxlMyf8DueNS3RrRR6BcX/HBPtG7d
GU3tIA9PQ3z3lXhaA1LY8OUc8IG5GhulTdyYgK/cx5IKpgxaFjbwEoivjqfjBI5l
ctv+dsAqqgyG7rFyfSwDunxa53pRBGNFOUl9SiGrDWWlSQ4+cSCpKqbOCIkVyTDW
f+vCUhW/73wNM9pJECSPqDst05kmk72o3vVMNl90gWT+nnRH0VpMOGck9Yy3AiOm
mCLsQxp3qzIpgdXOseNjYG5bE0sQEswcxsIm57i7F+s=
`protect END_PROTECTED
