`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z5PAHXjbuKTcYLIcXa+Vk8u5UB60uT8rwKYYa3T5U4jgqmdJAnGdSy3dkHzG/1HD
Av6ZqtUe2VA7VW+si4XiSmj/ZN4ZcJ59Q3fx9hXEFSQ8bTbWl2ZNL0Ye8XiEnq7a
OrrFs/UKVPjbVAHKVSTtgngJ9mdGQGhgXB3NmXZa6Rk/5ZSOXKfz9TsfG/sCemWr
2tEJMLsuQslQWNx+VXzw17bsOsy7ZZZaTnHepijfi2JhiWfnvT0zAyZFgcB1eLRF
v5NNnZNaoLsbyIkfLm97wO3TIHjbN9FKrzhkiHrYq3AkeUgQLaCLFKXB0J/x/n9R
UJCgJurEMmjw4XmgebqcZ+KqdXBPsgBNjgyCFwKUvOQadSkHUO2LTSDk3rUN8ctH
m2XcyPo4sfy9TmrX8ly2R6byGCgcoRxkixxSB/ClLZ9e6Fyrsy9c3VBU+z901+KY
ybxHUDD2pEdp44l0pUIyje8rg498BX7cE00yelPoiOGscltvRMTGUo3ancFDcG4B
yR6EFmg7JUFZvOeWWyjCAo1DhzN0wWmMOMIdUd9XdVWfSAhuQ8J6NiSqkoLYtfox
7wBY1WSvqMiXc0zsMoWzEHpmfqgDzbwyR2WfI+YVN0edQbI3H1TcwovBsou5vnax
/gLRdRCR9XF5y/dEHXOgQ9Fic8pGJGEdLn6ytFxc+6WJqwJGOlh0kYmQvOQPawB6
RSQLbT3J90Fbtw+bP8z+JBFHxwCzlh46sbqpqgrggk8HdvBdJhgJMU/qEsJ1zphC
9HpUDuFUutyJt1pFNKx5stT0hLrfgwowKmuQJoZLRUzN2nPTDtiZkniawa5SBsxy
pMWaKivmEC0ZbWVO/TY28NiOvPkPZVLS6Y28kORD66bq5hks5pIASKRKo+nSfIN+
JvWxNhwh1Fch5X7vqG6Avpkpc4zyfGiMIyizMSnFabZ1TI5Slo7sK/WXrbj+b5wb
BPsN5YuLqAaKyExmika81YquyVWKBNOtwMU+t+g7LTkf0Qqf6+3mITvcsOKjdIby
cpx6cIw5Z/oYGhL/NOaUrpLt5H6euN8h1/VkdJZTMh0YQXXtfSJzok0yuSJditJh
ARfh7cIGZvhbINp4jEWqDG9+1Gg2kuaoR2wuIn1JhjhHG94bEshYybmQ2o8vmwOX
v6sK6U+K2qQY11Uvlp3SyyimLVehTVIREnWFUmDBw1AnVc2kzKITaYtqeI0j6aly
QTgESMeURTjRiZfq5v7PLTdG2MOsS+pwwMhP2XXF/sE+hcZvYCC3Y8TZnP2ut2Ep
yC52HkQqT2i3vC0CriYKDO7KXV8VONbEtVRAxeO9c2yUB7v4jHiAxw5yMDbr/0zH
TrI8Fx16ZUKYjcTrHuqDe+SSA/T0QF61BpVR2gZCAIv6kz1E5wsc0PnH/Z8wLeG4
HemvUnvcK+y/oRA42E0aD2lQi4/6YDGuftMP/rFbO4GOy+EJyGndV6eQxH+R0pif
Ngoo62YSUPgFRJAnfi3Dbn3LvyikTWYx44hPXbzK7bDWR0Hv6eSSR0rsIqghuuYO
KW5f6ZxZ0aiqqBBeDSNMiLd1Og5o07lgZzig0d2OXwMzaA+2Kgw9YDtQ684VlrwY
IAUa5USv2uMI4f4N2PlSfoeWz8Iy0/ku7XgweKyyGq2VTvH7qXAA1uzqUjVn6xu+
hoB8e1me8XbHKB7F2PGAAyMjA90nc6EFeQCU+PVJZ1aSYU4lBIL1n2rcyieP7pfO
sN8QzuNttnO5iEU2pL8i2dGXLOwC9zni84S0DVvoGnBJUZrpmWxmGhRflc5HFV0K
+/3MUBcdjoHDF4b23LQelvs4Gae7zh0nDBpzG16O0KK+zeXsF48hiHFLXoc+0DV1
QI6qlYBpu6vCR6XnyKrDDaBH86OLm1XS0npp9xbu+GvOnQDoOsNC/MF+PUNABMBP
mb/vuqsA3TSIFRrQJ5FzVIASzODqsk4lm5o7ZGBVfzyUvYyBm+TpY14xmFqhmfjG
+sRxDJinQ5cy1Hw444lv8sKbtEha2rnvlxuYU5Dz81zjXW+Ir1GSO33uWqdfNjgE
7Y2KLuzon2pvfng7On5Qb+aR/5haCRHBKEo274AFuoI2sVu2TMpqKXWzU/c8Skka
dVKOd3OeLCGFzy7KHeExvUFi9dn2X9twO6G59GkN1FsgKV/gvK+CaqYpA5GS9FMr
m32lqM5ABLThoybU5b9ap3m4wWZTdpPriKcKYoyXivitlfEA+EnmlLNeM9rubW4I
SpioS7CZ09dNjBjXb5IfCby2V70WnxmmqikGgQaRWFeIBb9fa1b3yaiUSZJ3lk3u
uDyFPYyq0hD87ubGuvNM53GuSM3zb42OLIOaH70OatmVJtbyD0HkpagL2AchKqFJ
9KN7lg0S9WfCBRiwqOeyN5Y76/qKS23XlRcKCdddieSaD+gIlTHpGs9unojR6w/J
qVqFZ7bW+JuVTU46ARoVNQ==
`protect END_PROTECTED
