`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Unf8GKIRLASHLVei+QFgPhdX+xgh4Pt1yPRiy/+9MTQQjYC3+O/ej/VInZ0W81jf
7EaAbRs80KaY3BzcOXEtFS2tLKURvUkuvj13UffP1ot7erKiE2Eaxt+jed1ndwVB
TWL6TgBlzADElZUAKtXPA8N0tpFol/y8/Z8B3SdU1gW6WdJc5vfTBg1xn62ngkZ7
VmOInWmK8hfspjkFnsuLcBhGq8swVzLxY98eaVKcGJlgbVFXlirwkTvWDHu1Qe/f
7Oly7sizR0qWH8lQVxU8HN6SJCQMSK4blZBBqTQVXcZrZBqY8PM1T6IqCNXwBD64
80ri2ACBblFcH+uNL/SpJVQrG1phDQ0H/prD2oJk8fend9TnYK+K1BQ7fbYTu+Jm
u5koTttyxHCRjt0tlTvZu/u0m0h1kWlIr7y1RN8HXt9RJNSQ4W1Ul003TF6V5asQ
EHTpMD3mUMQMbN9l5CU2EfdM3u8NIy2iWu1Jdc80YsN9SlI6aeaXdJx38kqH1/R1
m8869i+tIaZQav55nHSCfT5ERzoUOJwWpuNXFSPhlG9BnXcIGUI3FWa8p4r7vBGv
KftTyDj0jlfiBHE9WP6TOWemvqkhlAylaZdxT6nxJudbtOC9OzgD34oUIGdEjhVj
UkChUIqzTMMrz3yZluZNwA==
`protect END_PROTECTED
