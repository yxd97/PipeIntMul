`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0WYKCCGFmmPIbKXRPTv/G7gtB6V4x4eWUL8ZQs/WE9zgdWg+GjZS9ceIlx3FfYC6
4QF5s7MWCkejJxM9lIKVhtXa+/ehrEY7fWNd5R8B0J59I7Sj3874Ojz2Po2qdwF6
eu1nxw+Z+/S3gUiw5eLPMfUK7/fmSIjE60MCqEycrNYm1OaxRUfGq+Ol3ibRU1kP
l/b+ak+le1FHc4RWo2RznH2YOTP57+cttklhskSTlB/IGsu+yqF9Pg/RbyfObCTL
+63wEzeKqpvPBfsDjEr2FsHR5Sv9Idy5oQrjTX9FYrki4JLtKyf2SZqCq5N/hW7B
bWISF3Ti3bfzkTM590Xia0PVVNb2Ft9Hoej8JMD9EDO4oW2kMNnf5ARL9dZf+asJ
guQUF6CiRYO4UWWnPweOMKfUpmXZKRjJuTBGy5/da8K6V9m71BRMHf6z/oDcOota
YySkG+36RM6sQ1xo8DBX45UrBkBjLJaktkpwCIw8SeU4gBJCl4m0IQN+OfsWtUNZ
VVcXTQ+hcHtGQ0BbZEoiMa2vi4z8gioGv9vcXUhYJno9vXNlt+wV0Fnhrw5NLGR7
nUWmXoi49SO6pIBcc/dVEjarKVqXHcGAvxljXEftrGAw4sUizIdne3WuEtDdVieU
OX2x7Fw9icetNdd22vDTtufLv7lwS7TQ/O9jA9Rx1TEcfvET9LhIf9rxmYLRChuC
wfuF2+j9W/cVCX4NkiwJg7GmACsfnFQuz4byO9u17fY1z9NqB7GftOmDLBq2SjHU
QQHvpaKwBiLz4Ugnrh8nBZ0VoBw0aIqpQOvF+UvokYjrJ5N6GPV8jB2Ve7HMCDRL
CLdhJ+aZdjnXab9WR7Istn+7AtWW2h4F2M0CO7nGl57LLCxa8TqmZh5Qm0ph7aah
mDzTQF10WKPTi4BTyhxcHJqT1DrWm+oOdbfDp1pYBBIvOIO0nNXrdmbqLJ5ceNjm
4VYhcqLOcb/8iZ/7W9vjGTh10fYDzOovuKy2Jn3O/rv1qXSVAj/0bOv0Zc27BuGf
j6opS1qR+PxACQiD371pq8SqFHwsERRqi51snDW9dgnuSJxwbP9ICSZu1J5e+g+X
DJBBPrtkKA+lxSCvQ/pMQkLjaCGe0pGPHLvKIsf6/01vCUImEhxeZb0UseN4H3n5
335K14eAPgs7U2Aqgbk8VeLMc9z7kOvumYnRO43oZxf8d338zKY05U0MnrFD79d9
TCkccsh4qZzx2oLKOtPAlY2TS/iRqhJQTKT//VLNQmS5vAP8YYkqpiLuS+PpogzX
+oMk/CfA5q8TmsFTOggot2n8UPQfrRX63smDhiZbR+FXsz8v4G71a4/DZfa7l5bx
tAOS/q/rZqsDF1OfqUY1bBgadJaBogONv30ii6qDCX4dgmoG03rFN+NyixRDasKo
6mq5rxkGPMb8HGQ+QRA7bxF0bVi/22f0sRByVZJRF76aIELx/sSugGQwoQ655EMC
EHoPeTytQuLy0boV7h9YpK/kx01DnlQWH5D/8z4uFkdutyfCReLTqSACyLLkai9i
IZheWLlZaW0G7zUmZprR3bEjMRo4BkZ5XRmbuexBCj+q7Hd+/q9gC7U0boW/LXID
oNGsaFxARi4AfnlLAxwjaniBA9KOZZnB39YLwjVcVKHLBZM1u8xBMc5WLqkbo4Ew
UmHpoBkUXwcqtgTnm/7izjyNwK9wdAJEP1kkhR0bbmcZ35SWP9vn0+O69yOmrYIt
obiLav4cUChqemS4+oJmhJkyp/XOe/zad77TsMWaFkTNofdixpbCFRA3JGQMv39q
f+2iftZTSExds/9v3wk9l9a3l3yG/WMHoXKyxGcio0ByDSGsDUpQFwl2dnNiOKxs
Fmg3sRzEYodAoRkljKYofob2OCyu/AHN0jpkAHa44TA=
`protect END_PROTECTED
