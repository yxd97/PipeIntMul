`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ekiBBETzWAsDXcXnQTBF6zFsb50nazPw9JuDQI+c1BRId/TT8mn1HC/8jWuoQrpb
XDhLuZer5xJsn6xrOtMpXpUvCG6DysAjudoNetD0Ur1s8ilZ4cDgP+E8SMgcHqxL
tEpdXfhHPDtbfTrg+LSASNu8t0BOdmcfRt+vjZ1HNnyTCFtjYNZF6wyCa+X6dJ+W
30aOOBd/QUSpaoGp9liUNjkVQ/vtc+AxhYCA9A2ZIkfW9c6ltw6LYadmV1LCZmgW
hLDV/sBmjNuvUWchDknvJzS00OsiQEs0J1DnJbkCeb/xf/VFerYuOC0Z66SBr6Az
e9MTNlmPBLKKCAFUByncFrm4qrUNTOEyGFp2bEzeRh+XLFK3+DtBpGXvlDVh81LQ
EudICrKADCnY35C63gTD7zUeE4w3Xr1x+WTDN1AmDZz916+v7x83bBKklJ4izLfy
zcpOaQo8nezNFHM5/y3Wkwd5nxzuauvjTiqZwjj8IyxDI15BeppPH2/mKitvS13p
`protect END_PROTECTED
