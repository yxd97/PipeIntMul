`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ikl8idckGAjoaGBFAcgbiMZVB3lFnsk3TQqBhgggtYMLjai97MwfLuItOEmCKE4D
lsBUqG8s7jVTT0vT19OImUWb4Bx/eHVsBqBtx2dDgLM/pSjdyQU5GVR4Q1anGlSl
sjm4DFHJLUqnn+ZaDJXKbtq6+imj9E7BmJcxZ7FpgNxHM7P34XSxbnkjLkUkT1T7
HCvqkpGbyhRImmin1RDZqkxrrDrem0V2oz/tXMVJiPjZqvznl7hh3Lfi1yV8wtY2
Xvp8Knz9x+2yqvsRED5d26q8cnv6pier8RPC6a3PBK/HpsE+ocKykCYGWLzgp0KU
nRvaw1YsjvRpURZflwEBaUa7nyrZhbWexRYxeVHLVrxubQRqtCbwuIoB9gG13/c8
SSItjUtm1jTu7A2bikDxuKigKY5889XcW93hxdtiH9Uglx9VBaFmbrE+cKyyGasr
`protect END_PROTECTED
