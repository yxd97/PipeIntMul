`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5ExWoTrIoK+vyw5iaL3y1DdCcvW2HRukwFgbgra69B418CxADmEHNTT8ptiKCea
smQCZpL+ILo1Dw7Kt8FAxi5LqmDBkCZ9bhR/wcsCPx7QHlUTVjQdXUnnueQUnn1H
BQkY7cacrI713I7Dxl4cUjzGQ1veUVh9PDiDMrsoGiXcYreAQ7qSU9YNU1FOL573
14+aYznKaIzZsO6RzvmdCQmspq1gTn9ydQmo6jOqBQXXv3O2DYAPsd9jT8bQRz/V
bpYQmNMqbXmLK1yDEiYmv03+q6QkKiURZFYopgeid/Z5h3/B1RDOedfCZlKX538y
kLIn6QwGyGHUOiHEazWrmflvnCRkO2t5xZP6ZAKjO8Z0gD+Y4wx7nl+bN062BzLo
5pMej6aXZxWuGmk+98xVntiyUiCzdPobX9R/JI4GPPRudDfimtI61XUlJeP2IoB9
csgR3hhmJ9LB8Tf+4dlcjoW1zwPxDnv81leKRIeQi+2Q+aEonYdDkogY3OMlFygI
B/+qYuftcbCaQgI7qtCirOS07L43UGU1XI8vboVfyrVFN+T3M2iult0fKXswrg+M
qhWyvD78YTV2BhKRzke1P2Ea7v+8Sadyg8BgJoEI4cD6wwAiIftO6FPVX0ny4Fue
QRXSlHGfSdhoJBESOXnM9Fgdx/E/kjax6yHUubBx5dO9+6fbMkffK/Uz/JAeNRF1
EawrJ+cN7GKZ1ef5QdtbpiXcw3lX66IMfRZL7O6Nfpyzhvcm/h3sG8KJ0yN6GLHx
blFiE9o5u3wLdpyTDSgjL79NCbff5UPTyXHcP30Jd7IUhhSSsJG6vu2lIJbO5pvo
lVj/90DqiimLdsevJO8Ht4QY3S1BBcn0kMLD0qyZPdU1JcWl8EjmaDRzkyKQRNF/
jxUuTxJ+pmZ/JAaTljWfcDA7rLBlXb7IVCs2+HLV46rghWFGNqJa6A3WfTGNX+o0
ktI7LghASiI2My8hcKBLM1nomS+ggv99mlojpsFMtfz9OxQ/JHVTTJAX3hHOvhVh
31alGw7tYb9dY5O/bcbLXavdDQuk1o0N5ZH+PD76VdP5Bp4oWS03sr/uxsHQ56Zu
NPzv0g2+jQan+l6u+Q3m0uVzPTPoFzhHXdhWV4SfX8AbsFAHZFW+yas/hxj2NsLg
him23VYOHwC88gxKd6jGzXCd0OipidALoGEfsvMKeMiuJy9gLvwqBNohzzet4asH
rlvQmk6yJxzGItODL1G12CVsDz0dtmIyi1HFylvyD26hVSkk8HNN31gXLXHbMbi6
zjRasYiK9O5zxWix97ib5x4ZDE18rgEXmoGZ/We0EhV5h5qUe1fxVdkRYomOZaOJ
YD8KlWFi3vrveC4QVCRq7eOypuGvVuzOn+2B/qBGuaBLOUw3dsqyMR8p3cYey/Gd
5WwGExX2TE7jJS+Rh1Vm60AK5s54ZIQwybMY7DM+1amRby+L8f+bQ/c/SmysFcez
7Y0NuUwlWQnbktnnUvgwIEf/D+VJyYEWDkiH9KFdiQl2rp4eVfc2YWc936J872FA
TBwJ/PcTvF4VaBfreX3saAXyunVyP+aEgjPvfXrPqsKzcLQIgx6v54At/XQVgpcf
Lip3Xxwl1AVa9ZpDg4Nr7cmWnvj4eZicimV4UgvzYcSRri03WK1cKKaEAm3m16Il
698L9xRbDGN/3dJ2Qc7nXrbDBQHb1fcAeyOMCfOcJ4hcgsRrBRsvomnt25JHoIM7
X9xr2YjtasPS0zsvw7KogNteI9qnZvp1CBPP80hKk5mX4UTnSpgPCCk59+uBxzEq
H/qs9ho67eTkr7ZXVMQGUWspldBpDu/eWMRfbqPaT7Q1KB1nMsOHhPNKmi6Xx+oh
ysWvjVty2p16hiWjACnk3XE6nRvOtnr+N7BqT4aygOZzbXOpgKLtBUxn65ztpVYi
Z1uM5M8kRgNiddZGfu8d2tiy1AvP9yW7g9C2jYdGFQynyiBp4GADkNmepHuAEj4q
qd6ga5q2teBQ/Gli8XOcwZ6QRez7RDsj6mCuEoany7Y/kIYW5KkP+WM0+VoQOY/r
059hRL5V1FEm4ZqmCRilfZbuFAzs6vo4fQAwg8Qg0alVv7Fv9ypH3iJ1TO2u/1jt
ZMbpb7ANI51UDeApeVbion0HPOzUHPJZ+y5sidg75JZzaMWZzCj97A213s6+8Ud+
3EAEr/yPWo34cj6f85Sa5FO7ayeNk8lAeyeRPvfJv0VguD76KTG6lVjsptyNU6Hk
zAPrshptWMtSLWKyK/iye+JQNocW7p4iY8s4zZS21p2PrgckjE6Pm76AYBRge7uJ
QkcmZM475v9RtRG8d3ApE7MCJiUhyr1YDOWLyQAF4GcqLra34PPnRz8MTA3Q0e9h
onr963/3zkZJoVpNbyQyi7WbCpUynqggAMVsPEvjkT8MLZPTzOZKtdPBZkd7L7QW
wGLwYTc5eHAb7SBcMEn90JxXDaCzVuP6WpnKOzJioKSOSPwQQfbTqR43oWp9dtjz
Ek83chxJAPU1qQyelEluYwUzP8664JRaV4qxPAwW+x/6QjnTFRV7V4wDsVRTLZGr
4WzX4F2gZvQIGpSms7ru+UrudSBRpUQta9wDim9msc0tNTUIwiERjYmSR5+N/DRn
Qa6BADKS8rCyXPqvhEon2eSxHHpiUdnECc/TflHMvVBaIj49DWGbXOwsz2ZpNdnG
d9LmIovfcEyNwbb0WG+om3O1CqA7R9adDEUeyUmC2KDglsyXpEnStinFtUSbsOGb
lYL70PKeFSd95pBc56cZt6rgcqLg2VM7pON6bDMwTzUrTegtCQWbbHJgqKjto49B
Hohnnv3Ml6XhmoC+Li9XJDDlG53A7ZPS613qpChzI2Japb0B+fYSZmhrkoXkqf3W
JJbTVcw/VO0r5ysZzkUmMn9U2YgcLyy6SbAxu1ai2Q3uiT1RvIeIdfnbSkDh4qdJ
nvtiPz+tDgwFxHNqyIV+PYmWgPrHAhddrcEgzLhIySWFiSHtr+1xTsdLSQsn1s72
5mVkU7wQZdZnRAuuNq2s0g0qppWfIlp8CzaFL8WLuUz9MlqAtIwqzcU8gy43D9vy
dH+ZJtCHhSDRGN2pSVR8XiL8TPr/vUfNUZMyZhKa7hJ/qgq2Dh2Fn35XwqLxfvGv
VW/rYtQgBp0SYnkprs/K9pDvYMPH/YpccqO0wCu9DSWOvm9G463RZsfDvI+R8IfD
qR/gfHmtcHEc7tS9mlqtdY4BJ9U5AJtO4GvglTl+jzg=
`protect END_PROTECTED
