`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VnzQ7gBUfzYV4beSZlhXSfGrhAQ/LqtK5iN9hIRJt/yRfwLcWidzKJ15Cfkb+qba
JmF0LaWqj2SK+8IS4CjaObIQTBgdQC6STgK1ygnGyB/DzUbyc/xKNWcmfpjaCXGI
AK6hCWecB3ybiycqNBATqgS1n5hxCUfIh6q9oZHSs51LkeJyVVZQ+z/VfVDVQrDB
/FuQYTBY2sWiuvUCUSqQafrOMDrR1nUpIgg4X5dzH2Rv1CRvktT/qXExrKQETtSn
0CkL8axl7ekheQmRScHYuQAssuWKW7uNi88Q0VLGVx6SaVV5f29ITU50UQVl1F9R
bgpWs2lkmn5yOUpq5NIujdWqQKtvaAraMemoOuiWfqIr/vaX8CiXt5SyrLH8n9KB
ycw3VqEKPkh1tL9K/LayTdkQXf3Zxr+FBdnnKBK+AB2cdA9PRjAIAs6+r8JmxG1D
bk22PrPnMbGBxKbWyURXfOKnH5c+lDLSnxzT5hSUuyU=
`protect END_PROTECTED
