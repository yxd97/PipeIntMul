`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TlMY1dlaRLLeBWotWAzu5Ic0B/hoP1KgVBYph1wi2Jdow7kj0DyV0qRUlRnWvakC
PBNw8nQ7EGhZsDLQi/1fNbAd8f2wd2CmdKcMXJisNyctO17AyiujEJk/XUu7zi/n
yDDqVb7QJYMSymVLGXye1powdByF5K1t33xBV0Ynit8H0Q5DRDVPjZAIFHmhKQwS
EacYs3qpVqStNvn8Roaxp4xYM5rSJ/RuHmnXRr7upbS5dBJXgYR296g2h8qf3svN
ztX0SPWedMy0tByqxZJ53mMRwm6mRiC1KQ5Jwe0zphfB4rsEpaStFkbuysPBdniW
MlswbLr4t3wou7jl9mgGhuOUwtJAO8Kpmw0Vz3wmzz9mI4I3kfw4QWO669JXLbtP
tckKkW+7uE4nYuuAfgYx/WlV++R+NUJOORQ+ZNHo3r3cElsqaOXnxjuMWXZqBeyq
o7GJKVyg2rTjpEJL1tQdcw==
`protect END_PROTECTED
