`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7CpEATADA1jIobrQvbPtxQa6ZZX9MCBfCLckvq9H0gmPltSPC0OZR595DtKbwqqD
JdbQa38iOwDp99njDF9CXbBcWQEgOfzaiAFx0ZpjJ6Y62caK+PEngMb63/vx0IMA
iXjPEyQBahUvljxi5lQVRSxSF2MRaHsehYfrOWa62CMcyM0uQoDhTI+rM8w3FZnF
+miR6ZP8k29JzKegU0h7LgCBx+gpjWH8SWJHTer/IMyQWta8/bLbwJ25BNKVFM6B
jBCqrAyt0Q45NCqMc/kjfYrFicdBHfbQAdyWSzKdoC9hlpLNzEXjLZyD0feCvh8l
XYqJyi/kqPTLFtgNoMytJA==
`protect END_PROTECTED
