`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ys6BQynFOI2ZRpfdu7ljvwkiCW/pstEG5dLjz/jW0yo6EtVRgkC+22nI4C6Y8B5e
f7LN1otj50KNabc/p7VcAhK63KlG0nH8xjPxBBKmBhABqc5lmbG47xAuTZSNVZNc
NcGfBFsCfcLrfpOP/J3+oE5QklYp2PHWyWeRI71xK3ZWiFG0+cYU8Cks9eRH+jGA
aLOj16jlXwrfQMcNw70FzJhZQdlKT7RfWZL1iNxsmMAZ+lBty8uZdgsB7DvNIBMF
L5bJBDEW2pa/vtciK594AITcN2XSHB1DCHsgcgtBHCRyVaqka3i3uC6w9tX3qz//
y3B51+9J90x/2N6HF7bBL9vJm3ajtvPVChI2WcFCIGCeUjthicbRHscuGbIV6f8M
0ueEPeT3N+XWhJyhhV7+Y+pe0uSmyMw+Nze1zpdgn/XTnV40Vi0Pnkr9dGFnEJrN
uCRSIfdFc8oqOw/EhX812W5ZgUd2ldyd8rq4nWrSVtkoN15rZSPNI7ElJcLx9Iw1
u8iIFu0l3L79gX42gCeVwMaCQfvRznS8871K5ITX0I+oaKugvdNx2XVx7eNI6LJ9
2u02U0ecwaDjDMgCVSU3X5COD8WH+28UG0SVrM8qkm606nbabvMT4jNxGpufGbCa
WEqcSqL2S6HtS3y35hRUcA==
`protect END_PROTECTED
