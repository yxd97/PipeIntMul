`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
89rCFzuWZMiyBFMqdvQdD601zXp50gHpEWMOvXfdrVaXJu1S27yAlAPW9UvEIK/d
OcaUr1G8t3dvwid5wpKq40wjoEUMLKt01zX1VmbXyyfVoGi2Cy46q4Z8zbKoXQJL
Et9/emJ+rp4yZg4X2ap39dDSk6MbW7zx55CKtQozzazWk0gn7obSf4ZrmBbI+ap9
WJCqU7ChPkZhVOIxHMGC0T8ecl9RsTVgeeGJz1UA/M83t3YMoIMkPff/clZT1bS+
1CMFZpzZgyVSh+2P/UmQeY7v7dQgs8eoQq1FZwOWXUcOIe+3MGtZ/lUCCWIy22pK
afioqyjZa7gUG01AwJLAhf0/5EY+kaHbXCu4pcKMR+PaRd9ZENCTDLs9q5fYGZLh
fEAnSfDin3TR77Tt4DskQHrQIiesJl9uurtATtDQoMgXEFoSrKe048ccOsH07N6Y
Xo6ZZapD7XPS3SC2BP3FDy1Om4ifq1VmoG0VB2GhiUtj/nr2Cvp5Al85sUk8XOu4
9GSi5M464hFh5BOcljcF98Qi06bgjzjR9IBhGszvJSglwB1ZhG5uw3XXuHVpXYQ8
lYWdyvqo2msMqg2ettxj0/mA0cCMFHxqkDqHdflA0gJf2X7dByjF96mjI/OnzsV6
gKjVaoMoY1kqsQpk25t0ivTw6TBJqeMLdzlrOdGir7dqXHUxczXwkoQtp73MQZgR
yRgdXqTcJ5ncqXhijFrxwl7uDO/n83T58CBQTEyVQcY0npzIgBVy7B1CJ2jZX8LQ
5akqF4ccWPRBlH3REBDe8COg+onWY5jIZaoTL2/R2RuMTntWkIbhhLeURc3zBOyz
lTZYgEkMmZutm6tJYzo1/99KIgJfWPqedRvgt+mYblJNH6IDBrVho9PygdjuYsh6
zvrwwvHQPFbWPyQDgsrkXxVqaA3hX3WA016Z46RZ/BDUesy1Tj54mrartnX74tCp
JE9hrsWi9sa20819zSUkSjMydUZo6X5trkFrj10WiJPc+KLWpyDxI5TyaK42Pa11
`protect END_PROTECTED
