`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
etlerXNe7Rz0hP41W/PGFoqEJsvGYJsbHEVIhsxHYw0VT6eWAppkYNT8tmSFv4eT
fC16WiA2m9ZNEiHHX5cYKkdUhmT6z62Ou4vD3PYeMnEdVCFeIURZ6aX64HnY6s40
294SdoXIl+itKJp60V+iwNplAed31WHe1GaXt5CFISVnaEO/hzUNCMyNDJKWkWgu
xA2+9LtJ06pRjdUyPttJVkAYOwyM6CjIbzvkacD7u/80SNvqJt752farrxgU1CZd
wIZt2vQDmThQQaugBkG0sEgGPf7/ykSktdE+CUbQy2NbQO1kw6JhusbbJtM8hlee
g+sqH/1yIyj3QXHSzk4Vaz6rZJVVY16/NZoE2XMOlVJsaRz+mmIT6TMPyR9xSWoB
6Sm2BM1t44qoGSAUeRNZ5A==
`protect END_PROTECTED
