`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETS9KpIHeyd5nXAtXJ/4SCuezS43Fln1QWAeEo42LQh1P1NEjSRJuA/2pBMc4une
WKtRNVNLaNTM0FBdvszaUiXxWIttuVC7BsISdtrapAoq/S+Yvg8i1M5dHOI7EdNI
6VxvAx1BVaNF8VkTNUaqG1nnPxtUgEmwjkHXbjVOyjeDrvzVtyQQ92k0svCmPOxn
zv0zs62jb2RpskKp3JwNk0luNc7XXzFvMlRWykMhWrcH7A/+wzUk8g+yITd48XgT
HnQxFKUlxfk+P818OXN38T5uTihDaH2TQGlBMUDJMna57q5bDebqD5fIaPkxN3yC
uFUvVvsljPMBlkVFZRBWoMB5XFFuXSFcWJBrqH8CAPpU21XD0wHQlXkyqPsvW4PG
D/rLOxgOpTWat6B6qcqfDgNa8Z0GHKon0Wi5wNLvwOjB09bLiUKTpLINnuvceMyD
2STwayN3o6Dq3+MFkyn69at6N2Y5aUH1MBkCJgKZ3XH5pjTPEUp/AxWU9PFG/fQi
DDn5FHJjr886kBmSExCINfZN3ZOKuHgjNTeEwLuGvKKXLZgpN4Eb/RgyZBe6nckA
`protect END_PROTECTED
