`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BW9inAeJ5lXwZcIkrtRjzm6ksEtsCzbm8w/ub5ip6rnTbLEXJ+OMNLhkSXiz40Sk
LhN1i5IhYUPV0QJv3psoS8H+M/EpgtJrxYPHDtCVkvEfBWbfvXKw+BdiF7WU62rX
hX2SXyR9Vj9yZVF6dnQRRFPFniFdXwmk87W0CZUVkVlfVpR8w4L2LZWZ5NXCRFdG
iCEdioy07F1PCTauf9T2YhwD48/+tgnVQTOVjXNzN4vTKRyxNNwMAtEvMRPrlz4T
63GMMe2BzajR/RLE6+XDflIIINMXc5xM1ZOEWN8089xN/z+J8nqgaIaHRIRpsLZV
/mszaCT5g+/eQmXHJletPJctsAcIeJwsl5qo4U8OpTzFt3zNr2Bco8Bl0iKWZLmP
kw+SctaoAAE8GFcarVNy4U7ARBQRxdcRnvw5CTMDdih9/sDuOXW732EHP0XWJhdp
r3pFIMtHd2xNjcEIQSqVlhmrlWDtn+mzVcPiRDpzLItl0WMLjtDYqo60sHx3z/tX
igU9JEc+yyrLD6N5HFsU6OnvRJsrrZbgrE3eBr1RJdNIle3WWCCZwSkJi3tPLlLm
r6oNIhh40wTLPKVZGkPD1tT0QL5gKRuj1JnWg69WNO9CyxfdpxVdWOGt1953XFKn
yTwtvEo7xUWj7bF687Zpv2TEPMbQnoQHvYbNHRYfclzEl119Z7Wh9uVPO3/un+xT
`protect END_PROTECTED
