`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
14jmSxTCuRuwLz85bm3/Qv7F0XjWtiVVzzFbm1/+uRJggFh+zWYFSvlzqVsrPv+I
ux4orO/cmMLa9WQfzRmdyCr2CWSY8gUi9l+KO0w0/ZmiWcEr95GciKzWkYY7iT8v
DmkaqKasE/rViAhL4CBrlQu11lFS9PvvfjeGndpeGIvnHS1l5CyTnm1/tpuY4BJi
7Eiw7iJdbTuiH2C1OSdK/qkK2E3/w7d6CgsPEolvOoBesstPs3ciFdogdztEGkLr
BnywqDYSO+qc0b5KMlEv3N3TKWW9LIRws2fr5CcmGmXwgfQcUTqVfWyJGqLnCS7E
rTslwPndS3jPZ7E7Gjg606BBQ1o8KW1msAMwD28CqNlwqqrsC4qpWVGBmPepzVga
MQQOq5Z6AtBiWNHvkfLlNJYgVt7nuqYuM+eHUm+8eh9/A4fE+BgwpxuJhw+0YzXE
o6JAARLXcDqYCapW96CZAh+EnJxCyktNPxoHsJ6oOG3wHZ+Kw/MfKv1E6x2oM531
XRcGfKKKBhopvlouTibKb0le1sIbmxdwfVi+RNlAVSYQPwmkiRlGNkzL9wDwcJcX
4qbVpiQMw/JEFToH/IQ3koQ8NWcTDSbhCZEap2Utz72JD0Nss9Z7Mjs+ryy6o+kB
eWiBjyBa2/zEA4aB3mL+5b16S4yXeMJdqExDwpeyswiLamjKbV1+LhWmt95WvmcY
mAYRHkyq8/0hqSQ3ZEuhQ1E8rnTrSzSMXHvPDB7YyzqgwYFCUHuOVoGzInZesCVn
ai49G+rzKe2+r9ZemBtmkzZGxvNX8mlyd6504CHbEx2dU5K06MP7uSZW10JGsWh1
YPS/vrKgF6EIsg7dDDAUuyXQrYIkKiWL5shPr0FWLj6WFxPo6VBsqDvgVLjbiUcv
qXqBAo2Rb8igyGxaS2phvCGEfY+x/uZe/9mMZHu/8K1Go+w0qrZrNtZckiSSZzmk
0CEWcsU4eENY7qv5aK3KAAnCHAxpqF/rRrZZC/Qxwk0dlUPBY2w82AbVkZDq4VJs
vcrxtHziXxl7rDwzIjHzAaDSkOJzklW/JPqYAtXxFy36ArSiPHiH/o7Y8/N+Ra6/
pcx8CuIzk7qKDCbcQ2GRL/kRU7Md8qqgpJ5SjB9bzP5py+WZulB76UX1WmCyIELW
WAJVK8TrY7/3jGYcP5aA6nqv/cDlI4ZsVK4zAi69JAupiZan9DuZDWs6ZKT4hJ+x
F/LrO8aZdKOylq1RaqfXBp0ESedLT51WMPU3EjaebCafAWpDNPaYDO5/ve/owArH
b+3TwcGElHmpeAKx5Qo9BuNycfoMrZWdbovnw6/wiHlnJ9OeCfHJF75zTpVfQjis
10q4RFAEZcbvu5XgpmroIyB5Xf1gKO1ngMqYmlUPql30290nwwKmjkKQ8TdAq+Q+
R1LhGQjlPCPMDa+fwu4aagxm7Mq8Xu2282pQLrsbXLvmf01CFaBphQ/7b2EqnLJ6
Uik68a+A9lbzSf0mgIn/9SwPrNioWgiMGh/j3F5qbFs=
`protect END_PROTECTED
