`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Af+VaUknSh4D+39Ut59Grl7+b7vN2Ud3JxFDuCBCi2ZbcJEKi7WPj+U3Kj9xz2oI
Oj1l4596XiUWs4sl1vkeOtdhAFflXRN3V6mqFdqLe4u/VxWzztaHbJGbyeYW3Vtk
3dBqYjyEd+0RYQVZhHnHbQV8g8b1BSEs4/kXCFFLeoFmzz5E6biqjsGU/PfmKyiJ
zLGZSdpPoxX9inkgvwfDv7O2qcJ/FZJg3AAK7a829wiKab+SYAodKouwsOt1uVuB
4Q4V7CoEqJ3zPGYfjoZx9tSNSGLDJLt0mtyJZM0OMhnL1T/qIZ4sod8NQFfWn9u2
Wv59SHGmuLnaX/vCkqXM995TkVx0EqRJsKhi3K+Ic4ZygklCbuzAy4jKoSNWv5YB
jOEBPdP8wcKgb/vKJZUr18Wpcuugf1fC72INtH2dC/gVeSyOmb9CfDai0ZSvIleo
vS65yyJ3rKiCMG+axOQYXxM6sWZt/DpjhkzDwZwWtgQj2fTRxcXcbJi9oIuNMWf5
6Nd8JVd3dmEK7e0qOsi5FQlD0o0lp/BGAw8t1klEXxW9G3MKEvWQUR5znX32eA2o
`protect END_PROTECTED
