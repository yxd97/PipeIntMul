`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DKgrY0M1UBvrARLq8ZQUO7imxhSqUeYdTRUcMTvkuOc7v4y2c3GDEk1KhFq+UW2+
y0Uhwgdcq+YSAVNta2Fc7xXJdwO633BD9mmxLA6dzH38dxdc/H4PryTUmtE0TMNA
YNdq6zhs88Mo11Ke025A2hMhw0cn3l6Tf9JfWRMZYI9yTMtkAnFUh+Mml0ZoURr+
2egbC1ukhxJqKBUnSY3Rp2+f+C1VWHNG/8jG8qjVInqS8qW7K3kqo2bN/Jsxa77g
d4yOBw871euI/5eG+6Tc8doEDLPJK35yOfyXk2y3Zz8b3y2r+1BE2+26jVfx0RnM
w7ChkYMpQOmwK2W93wVU8xS7Q0YZQYAw3893mF0uqu6rn5CWXC70ET8KVxWdJJrz
sLBU5I40nSFf6HFz9IEDTcML8goCkPne29VYo0rnjzKtTgrz7RGiP5T7R9Itrz6T
MfcIrg1xm4ilNmw1Qof2/CqRNx/iebZJ1EFVrc35s9Z82ZxFF0xcyaKYwTlKuaDS
qIsxzULviZc7PnnWYtbH7s+Z6eYKFetsbmEmVTFokrYHDzYVEPtDQah9oBvnDZ+k
nYzO0Sj2T4+hPS8/4LxYCuXWEjWc1aKr3EfnfDPVahlNzNe1TB7XX3oIoAYQvIXN
eDdLePPzw4p39MSX1d1PKFDm+9yCyIWqH5ad02OU28Yy0P+q2/xbWTODN+kLrr+r
W+xlUypY6QtMM+cxSXIhTYHEpQMPYZfZADNt91ZH7lK+I16gEuIaQSezgvgR9zWc
9s4vBWAGDSx97YBtVQj9FsVWo+FJeA5aJymaUsSKxFsTlzTGkvy8LUgTGjfHPtJW
HO3SrxjDqfi1T1oUpeQ7Vhi4u3XshVRNPzsym+sIXw+7pR+aKS7h3Q+F2pdCmwcK
GzgmRdA0NNOnONl/voJwVWZiBO7HLUhIIPAQ/TFyUT+nFxGToxAWdocC3wLxwmwY
I8RDIzCXgOnUKmZ9sYlrDc2YJ9hYikqBmHJtaZ7voyn8e1rKPf0pqHtzHb74Zw+h
pg73Qax6VJjEaKj/zvMkp5hgp82Wa7hPeLFXsLgrbHBCrzHAV7qguTLyi8O0rOFB
6NKXIefqbgsVd80rOJjorUYtpsaJt4pozaIsY4D5GXJLqFKIKKBC7VgobxnWa+Ln
l2Fb4hZJ8dthnyJ1MHumuXm9rixUtQcnE2rcIoW/hUZH7dGSERP+EPntxR6Pjgci
BFG/OKNQmis/pL7Yfrya9vqn+PblHLxmwYi1wd4bzsnfQJ+9KNPG+GlLADbxtxOC
zGQh1hzmbO16+oIaG0M+4ecSXlMA+hQVqEItiexON2bmbI+p84YWSSws13SUXtvZ
sBvYLwgIV0UWYpT4dcSh5CkGgSPi2bLS9AHUohOqwIW5ZrFZr2Q2CyUEmgeYt5Rt
/517KYUq05vbkAtQHyEDlQKo0gdmDspgCHKfB6norSzd7qoUcTiuVn9z2soL2lAX
muS0U7BX80Dek8m0+qAtx6GSpr6t4vTQJtiuengcRx6UxOulFhB8+nu5+4fKEpyY
pKEoDVZUDmPDzguN2yc1WP8jyW8/gdQfSxfkUzlk5jPY9Qtn0PS8UoiSmhbtcVjT
pmfzzcloTxdxr7oU9jsCXZF9EXIZkmLf8PVbpO0tmaGVrcHk4rq0ciQMLzA0SGNz
ZRx72ryC+NRB32g9ttAvT6Ny39hkFRoqAjKjc1wtK0TdqOrjObo14VND0v9FO+fy
IgTADY3ULAgZkNq5r0MfjWTz1hMx/AZcwNm7t1mcGvD2zNjUun0wfeG0ZCaHy+Bs
OtxMFUkj97PYVOHME9qYmDoyROazSMapyh+JB278y6L4FbJ8HDOc6nmtJ2w4NMYn
FFUmuN5XWwossS2DWPlsogNea99BGX6ErptDD7MGvDf5QC5rs+t263KuBoHE4d4m
0yJkZ+dsdNIB5My2CrZWZwaTSE4sLWQ/sbpCa/dp6k+QCyM2dQuEjiTUF78OjS2O
7gZYot3mvkHfMtT+O4vxxDfloniH0+en6cdv4KocvjxQpfQ0B3m4Mq73W+5SDJfH
VUDPt38aX+E3qpck497tkvNTT0+V/WaFm3UeYaZwO+CRgiq3i+P+VJucsRNlwOsG
0f+AvXENREVZqea94Sxa+Kslob5y5Ga83H6DYt3SVVntg1B8zpLJOxEf+jlv/QUQ
VX97ByDRCRv4h4zzbOvcFUH35ap0e8UynVoPqHbUPRlh7NcVGtPE746i9VC68HNf
BDVsPcCKkXI2U8a1Kp2yIfRGgotfliBkPUsm+hmj9isSqIUvdqL2ectoRz/eTHbT
Bkb1ADBZLk5v9WqFrDzALRZlzGvDpWFzsw6SmHtHNTXVg7Hl/T7X1MCvfsJ5JsvC
D12qmMEQlv7xNK0VVFkRXTmMhuR+rdV6fflY+yiYcGKoyS8Ah3g71xfKE0iHuUMB
W91odckIQlvYr9CKzn++J/heh+W5YOZ4He26gSXgdktwVyUTd7Ig0EUtIFoYAvqW
yL0FcwUixrUZ0fZYt2zw+DPvcXPSpEPy1xnOuSHCIanmUe1Dgn9712XwXp3hFnki
IXh4wJVri8xqeNUepZGQ5oK+JSarHm57nMzX+7890efuEp9b4gPM1Ikq2g+AwkWf
HL6fYDarIgJM30Eric+a/lysDlb28qLZj/vp3lEeE1It+31N+vsKFzdGt/Ze7koF
SNC2GxUYmOnLqUGVR/ld1g5Ygx7BH5Fa9jjlYlq+EgrTPVfWQVpLYRVL+PbSg7bR
i/ZvJZ/IkivlTW+8QwVAC78W+ze6B+JK8AqIZRpaXpcrMsmizc1fjFdBmqAwEXOT
FBZeLnbBDxGfGynbVI5dqZ/1gIgqb+rkcXTw6g7KW9K/V84N4ILTLJ67pd8Hzc77
ERAx+WJEaPtGcgZnyQNINziYLHrde+bScf+uSl2/7Gm+9CMP37SZAvLfi5hu719d
bR6C86SUiEQr9DxcI1nqSUtYAwAvToWcszDjpLAHLN9EdvFcemHDfgWzqAnzIRJg
m3N/qng4UqQ9DroIpMFhCgz3a75Ct/KF//j8ZgQ0zmGJ83y7nTldZZrCmG6DZdAw
351oVRwnT2z8PnD8EcseqqUq210eF+oOiNYJa4v0Sxe4CVF08G9fzFFjprASNrE2
PHRYu2zo4XLr9oDf0xwMZQ2S/h2law+8ZtD5rLjyfbyQmvHlWrfT1eDfUfIOwYo9
n98jvdjACx/QviCSu9EGDdQaV2ccHou5l2x4LTLvJYAau1/GZN0V4DV/TIj1yCk0
yfSrXYaDlWXwU9CSpt5pehgiHST/jzB43TN2DpUMRjZlsLEOVwQJinmvqpoByRpB
P11H5pz7FbHHtaNWBLQRBu7Kfa7EI1vds61JBaIEoBmlwPcPa+xCJxLSH7F0T/J5
Z4Y5vRaigxUuBnN97XgzcUMi1eirFx6YhySbi6qn7f1IGMSu7D6d4+IGb5MT2+5g
2spj0g3A6M8MfOrBHBTWsQ1RDD2dYtzSMTcVEyVqMSIS4pMd2JhPOfhTy3wX0s9g
S/KxrSlrjZ9lietH3KnR07TTaFBEZvHKxleW5FHA/EVoABBUScN6DxDeKjZR7PMH
MiubVRx+uJLyEaA2RWCUoujZaT1Zd9sUi+dQ/KD4usJlU4uNDF4NVLuGfdNEfgJm
2oH5H/z9VTguGwTuNxyeUvtGOIsoKQNV4C2gfTpadDNczIGin/5JD7WUZmyOdy0t
8wozSv03b/T9PeTsAHX3iwp4VqI1RYZ09m8kXEd23BcWIlpx2HYPZOn1Nioz4ajF
aHxQzEb7Qc+brLvo9p8qN5er/UfxTowBWzuC6cFN+n00N8zM9nO10J/scRg6ke3N
cuF/a7uaaNsjLYVQojI0uB8ZjuMpR773qhrOVdfD6MHDNKJ3jpxynGchxVgSQFiA
ph2cQNaXkEvs6oe3BjP5bo1nxhzZDT95hT2Wv0qy6vy3/k9oQjg8qIrQfb/hMml0
qd3hy5dB4Nf6w0oqzJs6W1w6ApLmHZ7yFd2gteJ9lDOpykLKnP3buekFXLjwtQbz
/jVANowKcdxOO+q1fjLsS1A17VDeKpQrm6WU3LH0QfhZ9ZY+oMhRSxV9bw1NMAk6
NYnmKN4KkKOOpgc3pDoa4Jjz4EfsoJtxDwVwXz2nQfvE9E3uJOQJQT2L/vLbtsSS
97ZJPqQpiAkSOQzTtN9v2UWeKXzgOQxTN/F+8z7PrXdA7HKMhEAUjRh7reZs67fp
YPUNkP8+IrHYdtUi0gvARQU22AFOs+qUUYatMHnqehRRSRhWK95UxJlItAL3xuEI
fXHivxOiggeSL2JoiZfNKZCaS5aZBglSVK+NGCjbNEpRTF9bfeqpgJJHykYvE46j
AMgO38HyXrvCOVmhLDO4mjLHK/IQnrGjVeEyOUXMUVUDvynP6LpAOZsCbY3BWo8U
lWoDxKEmCRC0YR111U0i3EenPfpLoNOD89NtRwj0Nn8IbI8r/r2HRbETf/UANayh
KJjcpDzCDkvdcfinNCthE7CmhOHsO+Cfr4IvBJ+qa5atqQOtcyyNRx81RFXCbcg4
O4WIzYGYXBgx0ZfzALZvVU8euRN7BQYYzjRelFMydcTtiwH7Zk2MMK4wGK6ZU08e
kg4/ryrHAA+l106YdEL1TZRrIphPPRn4vynbcg2HsvShiFG/qopyNIDDE8MX1sYE
qx8KzhcOJ36C4pmZiqsIs5+1ZldlVNj3JJdivB7P0MuR4BCs4ak1Rb3Xch4oACkc
eoJQvOoBJ3M/NwbiywfmQMcl0dtbOsIsx2wGMojhEeKIYl8Of3JQ2vWy+S5hU9s+
Di5NKHSsvjAcJRkL2IDYAlPYMJKx68quX4LEPbIImt6/1R/PnTmPSNFdPd10mH4V
rsYTWkwcEB4+wSYzs9UGxumHvSb4Skvlowsa73hgCmPosQMB40V/JDcB0dhB5XyP
D9F8EE1HkFISjVhcuj/bmmLSngJI/z0ih2lJluorhbSISYqYqg4nVaRj4cr7RpqQ
+NjxUVzZwTgcAu3Go1Rtl3RA73RdK3qhahwhgHBbCWdpe5KW68b1ww4jDsBefO3H
szMoph0YgbyxEiJTKotkXgOxC8mnV1RVk8PcHhKKjm+LciyzvKYNnv71KPO6EdMn
Vu06BeflJ9KEKcvWVngamwuIE5aGO+6F7l1bRJxOixZSGCAnCsf+nNl/vsXlWXyh
YE677/OOMvYcHjFgzshaPdZZlURgw/DSsn8wkHlvAVawpL22POFGOyxyki9rlk+G
Fmv3EMruKeDkdAT303Bwb8HvL41X9f5j7Aofw7EJNyq+4JnHMJ4yVTUuEj/UAnXY
JFFgxp42LnjuJXEJoofShBRIGDwoBt/0duDFebAVBU7MxeaF+Kf7zkrIH8WuegaE
ZiUbbDOoLx8ezEWITUBcYPBtMtsKwIOc9skwtqMFy3ZyqyCx1WzVttYz923ftf93
tfk2gSYGUhglUAq49PypbnN0dUyIThOvcrxPVbw7oqDtfE9Yzjh/CUAGTT3HSgKy
Zf6BUFpvMnIVBaAilG27APD5G5vZHOKYNSguIyRAdAz7n+/u3+qDr+GX24SfZAzO
+bwPoVRNs82Ra3KeMAI0uybVw4fNYWx65K8ktYpMsZRGzWPFw0jaOG/g4CN1tD60
Gzzo3M67kFd5cdQxhhw37Q+x/eZekleNcKIxlPn9F6QbSYn89J7dY+ZVrKGL0iNI
sTy8lVVHYvjTUNZqkdQ2BX2jfk6ZakUjiZcvQ667DRJQo45HwjspZffNNC8ftcxl
FiZ3j0RnZ4OzkZgaMByz0g==
`protect END_PROTECTED
