`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLUr0e3yVmZfOQ1VazKb5qOSnRwxeIUmJORlvJZ6duyHD7JIxggNi91RQREc0588
5CdISz0Bk0S985eMKHGL9NbJuSmrST2QHgH512u0CvqsJv/RrjZ7+0Jgs/ceki8V
kI4nWGfYnu4i+V/bzTKnot+ntyAQ9sIdloQsquoGNVb12pCU+qEeTGVb4Kdf6DYa
704ONZrigMdZsDdG9tlb96D+8PO/Ll4ccCrvwsOCtop1trAAW4upB5ZzzAfvLLHJ
61F1mplX2CH2CsQ/GgerQ4KkD/ni6TJHvTtkf41MlyHCMB6bL1zdYONKr2TqYNnR
ZlalJ2RsLLBGO3TxU5kjx+g3L4pN0PEJLg4cNOKCoYyKwX40luBYohO1qfJQz+BP
zgp+TlfvFvmaoLEai6maXBnQfEXcIQ6oCCRBXPhLcId4f+n6anoLCd1KiV2LXERC
V/hlf6Oa04hg0n3zFZ4TGvEUZwQWbVzkk5br1IcFo0EygCFDUlFynh4ur+3EKWSP
5wg3LuJLLbHZ1c3T8TH2FXJySEG0zJh5sGMcekztMezlM2y0g9C3RcwnDTsyg9qS
aPTUO4Ihve4mfZpne3/p00wmmWTzJSFXrYdchkfH2a8Mh8/1QeNoPc7TnCYwfM74
bXifcCJn4WujfyrruW4IYfonP33ysOVeVDAKosvXlb7gabXxGqiaE9XUI5ix2lVb
3Cae+PW/qGDo8pIJZN+eewe0p+nj0ZczKGtckLZLtPnssIH9ff6/xE9nNXlsdCcP
THtgjGbYTkrm8jqdeO7o4Q==
`protect END_PROTECTED
