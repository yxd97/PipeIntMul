`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ankOEZlrEfqQ7fT3JX8tIKoydc059ctmax1zY0ItZndOnqSazu2BMXcQy1LVCjpE
tbINnSxw2Mu1esD2DVVYOWqOV7wBMDZav1HGM1klat/Pyp4BEXSOlVOT8+QnDqqs
9GJ40Zy0NWZXnrJaSBc4/aFkGpivY880ZJyEC/eAQda8P5HcgIU51UaezmRHjM3Q
rpDZFeIGhJTiOGuO9Tr+bxQVRVipwdNcPzwvOATg77BHSBytGPie+1j7e0mPiTnn
oR3HIvduZpZ7lWcZTatfSJj+L4JsO7X0hB0p+b6j1GiD/Bty4EbFVk4AHCrP4QHH
zspdloqrPeGqNX4pWrpJtj0di3oqI/s8/+1w1YY2XHKLjjWM7iAJcc0Od4YXfZxC
orocTFfBHm1cgGyAlC9LsDPizYCuxAl7t5cE9LJ01MAf+Komn3yHKbu4DlIzx9YL
xi9C2Adbm86Y8OzyQ6vKpKIIHMA82PaGxBkgtovo4w6CKvB5fj9HKVJ10TFDh0Xi
l+5/RQNq0e/ISis40KJpM0wBdLxQCm9WadsAGMS20Eb8JtGJtn3F2GlLK8jRZyG1
NV8E+hQMm0HC1r+uqG+F0d7YJGcnsFeuP2F8wQnPRVyLvVVSkDVYWd9V2r7S6p7y
kPWzWoXkgqtlNsXpsWgpjw==
`protect END_PROTECTED
