`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
psBE0kH0jzZ+If9EXRPUj+Y868Ab9GOH2QnvBc6SKvCXnMPcjgfegZikqBzeLpT5
WpQ/kZPcO2CQpOv+810spypyW160P3fuVwx4de0bDrhwtaPDW13K6tplSy1ijYiF
KzU1CuFYQfncYKqxl6CyRudDJtlHKVe817ymN/L8XlgP/rqrR6UDKGIzEaXf77Tf
R6NEctl1VQmE6yyo6/s5X9ua7EOLikd+SgamQgQLZKbLfi196iYjfMUwQKjRcroH
uaAdFEjaeIPcHN8e61CXowajePlHghLxiqwt1cKrwF+5+cf0Ecsr/sDJ50boaTX7
V2ibgL5bcJ31z98N33n5YNMm7RGEbgRrIqNCHN9Mv6NHhuvie1omMhkGS8EzTfK2
p6HZc8GT5MGTlmFOe2kwHCoJZZzaVu8uP8mDZ8q5LiouXCnrgPlraXkYfkdoTXO1
ijeNEhz+TDpGabdenzw1p2Ov9l2mVIoQZAdmht0yuSizhLTOJFTHMDHCP6xv9LUD
dddIQAv83yALSuoyxdHd6OyAexPHgCyaeiQXWj7T1y3JpsLjav7nrzeYedbFYaoJ
14CKqfEzO85i1sL0kg2p2s2fQnV+Hu/ka8bAlUKrrmP8wBcpQ87FaIeOPNl7ZImq
3gOT2d2A472ZiZTy7NquueJMsvVDrSHudGTFwFG3tTyVMdKFce3IYruH2jEmrezI
2vX2zrela76Hhsnu42v3AlPs3cektee6xErxoOl8iSasUvsoyQ+Lw/lb9vKOGF0k
CxJrkhDn7jRrxQYvp9U/CeEdkFPtqQfUpng35PQDA0CmkMU0rocq7yCHkRF9Cd6f
x0dk+fOEjIODP4k04nI+BGDwNRqbjJxfkvSjh97TSPQBve2qMGynFkXCLyXX/DFe
pI/zC6Q/Oeph/XrEnF3AE+2ZD998Ki4Pllhq90NsyWjRlakCGycP/XWYqO4b1gui
b4oogtiUtmqL1iczpf67twvQdMEZ6rv3og4gpgLd91XcxKEph8doV2myPw+EYCvN
uiuf4FO7a3qNK01B/KOXUmK2ODvcHb9r40S8/N7xYVMNepbE7D99MObowcbd8llu
E4gIfJDTY4CCXYVgPXfN+ymtc+CZK7yojKCNmseNqb0lEs/GMza28wBx3GfEuAQo
KOzZBjg6D3y+QAyKQZ0891rPu9pxMyjEsN6kKXVnbMH0lTAIX5de7BXQqjmKQSTU
DtRAqJrv75WC8ys42bFOCMUxOECnwqx22rfvL+UcE7TzDDpOUH3ALNKb2vk6qpDI
EEQJYafWfIcTdbnW7nC6ROEXrdL2dnELaToZO5aKfB05Ngva2+VVnFsdJV/VOawg
z4VBsMdfsh6unGN9FqRJU2cHlcU3p2YjRosiM7yv9Vx22G9yX/qABeXmjEbUeVLq
CPJ214Fw110Ly2UWNyuWNjhC1ikosmhoOYptU+BhgmGtnnFg86/6WPXu7rfELQDY
aq5gW/6l0xIkLR98F1LcRqgoJh3GPS1J+4/eJl3UyLBfPnLS7pjXnj7OFwRo+GFv
zmW7lJ5rDch+EwXtDrRUcbxUh2yChJici7hm2ud2nBAsciGyHQrPCAkvBwYN9XNB
wXT7zDsva8xNQMRJXJwNzEsEstaN8eSVWKIdFz14JVX+odJiKmsHdYWBdlbxSndH
eK4UfiO9xJabmEM2Jm0EFThVNw/fIewbvS4560mVQmE8M7QBDB7gyHe6CiZUKcfn
9FPi9XqX6B7TJjBXnP/J2gBz6qK48BmROKRu61n5U7UvQIrrmSmEgKKPKcnFzgQd
zJzzmr8JmloY2W9cCUZMyY2SCeb3mSkx2Vj2E1FEha5JyWoofhO8HCvQH9eAAugW
UZwbNGEDTq6IjBAa+ffN1u+jPPMNbPpjB/FSLywGNHi3CIgZ6Dhqnil6trNDFPSc
UcLIwlhqn1nQZ4Hqi0XlQ41sqsI8+XVDoE5T5gBETNMe2zpx/fXu/Ih1CFNB+qoW
/hnw0s4HmKmG3dkcYsF2hzZ/PBwIvvesUOPRDNTTSB5uyfORkMOCB74Lcrn4xPpr
rzl9juplmw+6bs9OYUmhZjZvWBikAhWlI03q7iWk9Bo3EAm+3QCcrly+0Qmn1HeU
pMpc4RyhQa997bYecrnbkFLnbCJMNewa01RjZVTvLsc6aP4V3fGvw4Oi4E1Hbx9s
bm/OFcF6Nmbr5XaRA39E0QD4NL6NG/cMDTzTo1qkRpCbNFThbjFmAoRzpNPEbyrf
h9GdQt5OEm2ma6WbcRRM52k2LHvkrKovNGSh/upA0NYVkVnU9wxmeBp5rBdENFhQ
s7jzcIU/Z3KZFmaZsYFOJQ2R/yBcypLAE4NoPGYC0te1uBb+GxzaGQq6ewPPCvU3
ehUDJI/4XB0LH1tjvHxbPUwx93WJK074kgz6xwyORz4+wa5mfqeC/fEbRmg01wc+
ikk55UErrMEpIXs4hbDmixfvkGxoml8Abzvf10Gy+XBlybp4CyRgueC9t0h0edsj
Ul1gPa5xwS/YtZKwnwPvFDDrK5PW+XgUviknF7CB17IqRxt1egVejqLngq2LqgzO
Yz67Kp25U/D0bJ4yvjs7O42FvG51mKeQgvTPl0gSzXzhge9bbahfo52Mzkau/VSE
ea/1MJIfFd7mDHZoz/8tmztIj8m+lrROMJLIYyk8KBV/4ud19VR8FKTdIqHp/RXv
JJXlzTaOsnkhbOyCml/CWyRlP93bs9zkL7+LiCXsv8bg7V7UNyiqEHUeH+CkY2ad
QzAGc01n69P8rM8vuzfJoeovRxk0imqahem4w8n/NnCUMK7a2/r1eWYWsrp2hbwv
zBDDtNn/5A3yEfYt+/ENP3P4q01GMAwK7Vkks/RW4bZwvw/42Y6A28Ntulq68C6s
CFOpSz2QtE85ElyxHFDCcEL6aw3feIZa5eagIoDpYcTTlC/gfrKaqBV8uswkveYT
EHCevOD4bwj8IguY5OJ/IKioc5r+VbXmVavLFOb4zg79OVYrrbtcrg5UwSLfcuJg
M8MtH24RbtaIGJjgteGCm7/GZZO4kIRpr3kNIlBcatvYNMixKYKe2ZThRUoTjKAJ
pa2vxdsnXo4aK8v9omy8oPZRfG0elHJXCYUvR1FQKosSr4T2IU5/93s95SVKKcZj
sgVUs9fTGHjYU9hAPItmk9Dt9l96WHgyLbt6ih62nW3tPdulhUPSJElXX/F37yk5
pnD4xGdxE7nrT3giOM9Q/enjDbxWnXZOAvnfQER9yJ8dit0owhGINq8cNGrisUnZ
nYE6inONd+PUVQNqVR/mVS3sFqmTA3h7PrfRO0fevOeAtefkwqZxlO52WHO3qb/f
aMd9ShB4JqiNGIK7y1XIpqD8lv9ft06ZGeckiqKyrmfrdfj/PxjXMsvJHztE7SUp
/oBK5BCkQ4uGqb58OFS2tJZVa+wxY2uZmY32UO6o9dI1GiPz77UKkIHk+AiDd0TS
O1KtwNLdbFkGvg/XIxud8PIDISt/MZuQX4TAJUa9E7jbYZXn/JEL+7a4nr3+25/U
SfW0t6WKTkF51xwoOCPFZptT+rjVR9uul2yiCdlhSicd/a4DTS/CO9tlOfHgwX/A
dKNEVHDkJyO5j7GxQNL35feFMhoXluxkNF2DYnTJp580/KMQqkU7SB6EKrdZ7BWD
2QkjPagVCNI/aAKeYwVhZc8NjZ+rm9ecogyyeZzmvpSP5Ty8WXbChjGMWzwblUSE
STbMWikBqlcO+MXaMo+mC+NdBqyBgMd8LvWTfctafkJtQxVw1mIvfLBy269YYiTM
MFVugCe36lg1I0/0gVmlokKuoHDqhnrmqpgI5Xu0vSHcuAEbVrvNz8Ii+HKGU3OR
PxM1sTYlYJDWocVouBrzxztWiUAx3+n2zTecRwprpKNzaWjxYtITp7+VuvJRr2Yl
iEtHdxCh0a1gl0nSZC17PiC49AtgL6I+4PS1NJ25xb9wffFphu4NIYrHy4lL0jUe
gS+3IZBVexMZyNC4PKlIQ3IF5Wtxc9++E6Jz6dqbEqlLRkAyu7HM0/AWJlQBiowR
m6ll2qJKbdRYBns8XAuALftN2LezVTowcQ8Tj6hxgQfqUxirDDdtWdQfo2sCozJU
svrFuhfK3T8P4HOf8Owlx9MjrdgGqrLZTj2v0o0l/CtGudgsAF2mlIY3coYXVHBe
PrVDV2bLrHiYCW+ruhvEKPEviHTtZrZZsD/UGqk3D2A1JTptRRg6jffV7dFedAHj
3jPHeJ8gmYFZ8pu5jLWhmR5jiVreq5NJacbtkzhRd0D+gC0dy+qtjo3ce4s/VQlm
y075QOwS5VK3ZsNhFBpucHag72iEksy9Qb0aqA88gLIZfT42CIHotfwe7xImutdo
fC9oXQ78hqESiPKRE6IhDSpbs8kiFz6M6jpztdBZnpYqPaEiK0+3ncN37tr+H+f+
dmLA+RcrSY6fbnS6QNQDjp5pyyuLGACQzWPfavtf1H4b7XjpQmfdZTiu/Ojz89iC
byX9eGl8RC6KcjroGx8Tg33Bbgx5IgMAcrQ6AbogFQfc6nsj3ykvf56/lAkD9S+X
QXZ/5CTH8iBfw2jxdwTMQ+zQDjV2OpZcFk/8INMyUqEdPHhula6vdXx+h8AKvuPD
kVZqbr9aW7zUt1mGtbJ4Y2jf6ZRyJj5qH+Spd0Pefep02jEXQHZQ4MMUFhz5s99P
Bqm277AGCoaaUqpNjRaIouofavG+0q0amQP38ypIQW9Y93D0EffO/MGr3ThuktMA
+47x7e2tpku8CmR4b7RmMgPR6NYHVgviY8dHoZnoB9tIr3ipzS86pLK0uKdqCjx4
ZbtOWshMAnVb3S/07mRkOLXa/syiTgkAvzBmwDwbnPKGyi6iwvul6cj7bBngbQ5y
GwErduc52S4hRR0AlG8HLc8PFTGlY7dg+2axDH2AMQz/n0vvTKO4kz+plhvYUjUH
zOdeax7tTFxYzXA2TdkpBxcPGFVfsBUTbEVAYKypQI+t0KJFqsun9JAZEo7OtWyc
IDKxMld/PE2zxima18Z+W51Uuk2Kjs/Am+mPWVjkyumiTQZkuqV0QFSR9gsf5bWy
pdZTbsG5WLPyATZc35z5+pjRSMz6ZS5UpN8f7YeceWWCJ3KMk4IkwoagnZuAFGsT
MRADkp7fKY9KwPS4/1GKcBq6cDkNAoX8A5/zYHsD6Wx8qWRJNtL53hIzfvlFpQgh
q2eVb6pUM5lnO2bYKKL5JQebknFGmxagFPduQ+M8xF6YcNjv4LQ0Pmg0SjmfnzJZ
pSbVAK0ojSRvF+y/1MHvXEvDNFtzhderjfbDG8LYRucLVHN1Bm46y53sptWbDRz2
8KBBPclKd59luTHp/aAJIrhpXwQaVFmN+lUJaLI28074wa68eE0KcRa0/7AwCGCg
P+pA/IRxd9MlFvMfG1KRhsGEu+i14/gordHaVeLfNh57TnDXcPELuoVUQFBXTSaJ
BpF2ncm9b9feZ8DEPs6ZwI8nHIIrHqMCPs3DKDN0Jr4kB1ZAbIbWZ0w/US/sLJ5Q
VsFVrvC5t7U8rq6bXa7vWRmzPF5TmQ0rHZs0l8cOS87qbyFpnBnKyS9u7iGHf4J9
+XWEf/wnjWO8gXmL+bpXTEd1rlyEse2ousLDyasFyTE3Cn5GjTKLl6ZOJbIh2CpE
UcO/mN5ZMMAv+70MlCu8paKAPN5QPWq6GsP1x/qxtwpTx+dl+W/pmC+3h6nx3znC
dHyNtgkwMJrvxJF8jPw7lmLevl8CZrFp5zr7aV6dot7f9D0Ks+oS4A+tSvPb6hZQ
gSaktfWGmJVw3t3y+81qtgw3FKBfZ3mqHxSCHPJqHOPeBQ+XCkKDKAWWsjeBTYDm
hmFqbEJV9ZgBbA9huETpTCYkb7W2e/b0qhSlEj/NuInrkPPspgkUG1CF5pVYhR22
w83fISth83xjeeguHG4wmBcW3d6rCTQdadRMxOOK1tEhlpaemZ5T5LyhQ63hoCRe
aykCVyaNcxJZlGkxVJizAX/ybZStAUnwfOI99CkgMXujdFkp4YNV+E4l+BC2cQkz
35GVJbBNu1SrZqH6+Mx/30q8EP9yZF+y9W7qGAgZDcKzOXYw33XiQCaOsIQ4jMRa
32e0jvU4VLEavhzWvrElXZ+QH8kCXZGqqZ558RBs7LkgMRgew7gw/9u39FmkQT5k
PVeW/t5plcTWRvW+4wDF0JEldyZQ1fi0sQgPrySESmsWOMG2h9RvMhMWmcjSWsQA
oOofXk3wDOsdo+nIXRcnL5ieOEhrHrFwgpk1WXke0wUzDWwYPPDGtZCE1NnQ4N1Q
ilT+mMv6XXPs4AwW3zdONLr8VlMzt37u12lLQgE6jcDr8lPXOKaJIT5+xmUKEO2/
Z2F1Yfj90UjTRbcmnysz+bhIkq+mwPvaTTYti1hloIJlulKY5MQ46fOhgZ3Gb6dM
OCecmNL8bbE0eFAX5KJ3W6iL2fG5GfRo7qyFqFUrPNDEWPNwDGQ45//WnWrQu4p8
wcESFQ+pA7RgSIM2SsR2Emzvztt1WTgRCgoRfmPtjXqoFs6oDays0TcPzz36mB5A
bfNKh0r0b4YC8snu6ZaU1rsCZ7fjCcUM7QPCAhYguz8otMzLzK3hTFVDj50xD44r
8btSdEi7FywYDYG4ONmBq82IgCdyHNuPFMl9GIHhyeZdK2SWh/B6MftMAfARBbqt
3F9NNnzpdGFKGwudgRUXiOThzmhfSWwO5VFW95VpBv41+xNjyUVYpfqB2r+oruic
wGZUeREVpGHTswi+EI6X5qrboMHsbCH/yjyMlrepYZcC0DGgOuw+OyXu9TgkaUza
3zOBbs9oBQSHyCkrpsL9Ggs0JsRX+UslASCGMch8eobg760GA849mhJQkAMA/wCZ
+EK6+20FN4GShfxJL0KaJHMykBu5zGW9dAutYLcoY4vv5PlN4TK6wN1yecqCJZr0
j/wEfOwKtcAmvicXH5p4oR1J+GVIUYyJLbwTwOdZBNxvE5MIoW11CK7tU9cogTMG
PFnu2SlWoQ9NmEWCrQL9omcq5VRXhVrwtgMsbEk0OwgxxkiDTuLn0sivaNh5WSsM
e8GhusPVRzgTorilV1tMVY8XLP+meY8kUyY3gmEf7rM8N447XrK41xKEybEFMfv4
k7/BKkRhMV+BW3FCIWzsIwUQ0C6R+a1CZ0h1Gk/qDiJ64ppwjP9aPOxUhl5C2X6U
EY56n6lITJD5xB3V2DhM/N/I4Tmzi3ReVxWf6sxZ7tbkWzmjMPqnlxzdP2XTLMlq
I280R4Iu/ZPhinztnmcoe0+llBgB0MWrdUOW0ue4nUYV920oCZspqyLE29pkPWR8
AwtREnmuFmVgUtJcwWDYfu4GK2lMezC7f81Pu/WjRji6cYtr4s0bdxemacZWWJFI
ysUZOgLROypSOP9j5qAtoI89bwqViXNsMJUDJz88bepuBVFrwYCM5MBsVVd/dlQy
3o76UIWIgniEo9G27JCr528OLn5GmFydAoStOCP6qo85Ve3i2CC6Tf5w8AXu7u58
IUscA0DMPsZoWKtO/50dBsN+ySJvkSZIc0ePdNTy4CfvFQfuXgJbF/tNTgzgcOg9
XYsOifNPgKDqHwYu2gBpKuXaHrOh0DHm6X4Z5/tA/FaGyt1d8Ltp2IUAxso0uEOy
N1ywIPb6VBpaLOWn5gCDxBVqJ49oFI6sS3W7EWUC/C1KgdHYgABDvfeAWyh2O0vH
u1qw48IF974J5yYu9ymA6TH97yuUrs3VOByO3KqASXz0utijkqh5SOIK/cWNVHqW
UaoAWfQA1LQmpOEmxgMRFz79rAfLdz+sqvDEDoyqFMtyNpCBl5bWC2qUrJCdBZWh
OsLzwgQ30OFYAno3ew9k/rNbxTWVy3Id0nfXIxCnkanqzgeCsTYSBMLUQMIcOX3H
+YZfY+MCTBW0g+YaGAkofTR+zpSv5qrFq5uUH7CRsJQljoAmIFbwzas+NciJ0Q3r
fzu4fOMIuvJp0n5uFZP3scyXySRRMcKZt4TX/IbSy05cCK2/Csk7cawqkpE2O+/p
NHvzNAZYdU37PCBjbEHq8YkhttGgSp5gbC1ca0Us4lM8BAQbK2BhxUGsc1qJeJiP
2r0qRtfR5tbz0uzuT3qcyXwT2FSGb8WVb58thK02aisfpsXO9a5VODApKp37gHwn
YR2KEAItX0bmaJRwEWjgcmAgTJntmcx0w32f6aM/GeuDpMl9ZJNUWFLA5mTgGTWi
XyZgnIk2852wFhEMA50GpDx9N9VAWk/QsnJCZ8PCpwnZUHJt4tTVVFKKM1JThgNX
FZmF9yEK8X9YulJS3shWTjGUf+uSlpYqC+2vR7PL9dad0VIUWq/DDWYdXh0vOyhd
Up3p6WbWLRpmRvOiX4Vt04IsP0mgP3ad9WRb5hSn2CbaMROdjnoDgAJxfqf/jGxR
cTMCbs6/lLNrwZWPoKBExW8o2jqzcEK6ZvKwtYKFhI5s10Qcc9k1D1YximAmx7qr
R8MBnGmdbAyb5RU+UKT5oKDg/qvz/+vmX9C7NNLQarlscmwfIdtN/Gd+RTpirTEe
EWadjy0e6HcqPagCrMqMMfQ/d1dtwsWISUAcD8hnqglx+GJ9auWJVBBA0xVy10GD
/TxSbFML4FjcYuXSw7aPmcv7eDdu53RXyia015JJ4ozRr7Dt0lxK88owr4lSj3a/
aJDu6kMSVFiVwzfatDHaQ9DXuftYV6pu0oQdx9Ms111/LWWGKzo0MNKXfv7qLTys
A7GRZHGWaDY38u2QKKl0N2nMEd6aurYUxlvOjWH/wrKAvFDe5+HZVidABq2mrmEG
3+iR7S/Eul+xL6XvyfenFhpiDNgBH830bjgqRnbYuZ2BTWxyqjl7kxOo+pxSB1Az
wUL7PzuGJFTIRfPGlkSIZ6JCKEOSxyZWcPlpY7Mu1K2RiRA8eBO/yLg1dSqRtVvM
S+i+sjGqWpgyYaguu4rDFf0Je1mmdSyYnHIjFHEEbMqN07cc96L6qTNfttiQgC2X
EI/9n+ftgrKTeuK3msZaAiIs9KVC5LVAWq1dlXAQLaJ1/1aysn6Bg9MGRjdyL44M
VqRsuvvhYS1Jnw+n95O1brNWoHNgY2+FA6vvTQ9+N6/Vq2mWyqMjPxy076PcXToW
jH7H8Rfz/4XjlvSdcyBqTtsKnbIR8UZcAjGZFQq/SILbkVPg+x8g3EuIt/AbFFPF
ph7SeIKNJZx4MyQmsszzP9Lj0nhUXrIIAr8ERIHnbq7YYAshV0I2JNNDUarAgUL4
zdhZqG2M75NCg2ZSOngpPVq1BepQff1BxZICcYt2DTFybGcsZjclN0FLaTBUs70Y
pQl1KStr0br6Wem65TCyJd283XAkXsATaz0gk2MSj4kvjDZQRQqnfX0vmwxnWRcO
MaYZk1KThEJi0UWAtkW5zNcWGjAiymmqHxQX388Wb8QcH/CDB+EpfPSEOcn8xQ+l
5dwcWVlx/pZ88bp/83GAm/vtzrr7Eh6TX+2xhFbnYbj3Plx3rppT3cnmvT3eb9Ob
k0dM+VdDG2oMXxELfu69weUOTeTPupW1Onq5fBG5KV1WATJ2E6NM8QHKN2g6MV5s
YWBjUpzawiSHZqUtjAe6xN/VVk9QWKoIgtWzh8HgfE/JmqVaHqS/jvDzk1j3YUJR
xP84fZsSa+sHJ66JhgNk3ptmfvxxPkbDj9z7cGn1f/NqhAF3t1nm3J3zmj9/1/Ed
HPqcaN9hvAmN8neOxpUv8+GLJRvjW4SCeJZGT9xe4sID2hZPLw44BbjX3YZRzyPp
T2Dj3+AZw1pS7xKVHFrJx6j0Z/GQxCxeD3NGpAxscE5O1EgDwYY9ghdHUKYwixmh
q8Ez5FHsNf+wKnyatE3Zj7RusnGPaDuP6Ln+nLtJpeeW7KGM2Cx+lbvYNwRnzcgy
eHCOL0N6DbEdKBeu1AELgSY1oK4qp3LWDlzN6Bbdp4AjZtIV8hk/1ZcLTIxmK2ob
BFy+Ij6mc4ey1lBLd87Cf29a5gY9J0HFaTId/ySb9HiNOJ0DgWSadFlTmtCrsF+A
hdoQpgXCXUOVr1keekPAmcRSIYNpT3OVqg835Z4C82x3CdQdC1mMpWrCSJD0XzLN
uGdHXa15n3pR2TOxxRmq0l0H0s0LVhcATGqFZH+Id+rC5TzNrFysyyFyU1I42EMk
hThyBWJ4+8ppC3+p1oDxi0ev5kZefxQqmeA66CiOJYphkkY1v7p0ADqQLUN4L9Q7
yFSbt7LaKResnZ34s8Hb44fsjAz7a2eDOcc//mUrCZ5RMtcqOAenBUlfrCaJICxh
yqiSnjEW4K3g0QrYXqQF/iRa2UEGrzy4WOWXGW9NHE6bEZTMgVDOARI5FLpZbq4E
UIbeDee+8pPuOYHL0eyOAHQG4B253xIW1Z4lGbHsr0oPzA9AtCY/8Wmue1tiPDxa
pUeaHsFYSGumvCk+ibtPzPMEpZZBgkfVysFKYJkielK4EEt1LEOYhlPJPhDXfQc7
0+zIislLMmrWqlFsfusu2ggQutcoXUyyV3SLDCft0DsSRU+vMFUU9BDy2TSAM3X0
QTBuQ+3q4B/6bdXkuq2USrNSh98d58CxTXf5+wNrJx3FFaITQtbPo/BQ3uIU+BGc
HH7HiVwhq6l7jc8mLan/GBC7qSb82fTkKFXeqw3GJxlF7tVTSUUA28+eN4JWu8GX
7Q1g8bNrjGC2yac+TGIL2Eos41xuOKk/wXPovQfJC/0W4R6rtFwRtF6GV+Fgdtx/
VO+HnaNiU7370mS204g7UBOVURj24eP+GLk2SBVwM1bfXxR9rfK4gZzlu8TobiJK
xk1eM5v37Uyz1spFn6TSUinsn+OE+OQdBPbw8UG6A/lVi9TCimgMcZaDtAZmKkAc
LET7en/h3Zv/1X+8xw8jy8hhGpFcHP8oI1nCb1G2nDTVmj+pKGeJHsdikaZYY6S4
464RIpWz9dlGb+hDmoRZMWBJqA3jJ4WRfNMNwhCphTXjHooNFP45LU0r4TVzROJa
aDNNfFYH8VNT6XscKGTI4R1R6ofok0IdubJ5vFrcsC4zxkd4pzacrh3GdL2ofI0l
tOdGrHXaoJayhs+bXa5JPjthkqBV+XFumqrNOZLyK7i/oS18877JQUBxl+TsJmeG
uyV58dSyKTxVVmCfvqNPROKTjBsSUJnNfRrYcHWP8Lfc/zxxkaJ8rfHv8xy9HAUS
xqbUw+3SKv5AGczHEW9f9SEJcZP2bYYSkh6ePlA+oQnM+APlVQPbphB6526NyQG+
ueXv5yHsdlYAY/AlrPpiwtey0ArALRWjQsWzChNcUi1gG2nnSiOlNI9DzYL78kfo
W2hzI0qRlc6IGGBbWJHtf172O+kBndfTB06Tzkj0huCxy8puoMV4/jp8X717kEmF
bh7GH8f0Q7VKqQkMPI8NmpMK7CZTEpeNUVUsnHyi0F2e19E2kVbAF8ZA9b4seuG6
lToR2Vj+dKyyOCogz/kGDPQLrFpW3xYFJt6A077BZxo+w7gBKjoy190lBS5gB1rb
4V9yx0l8Itdj5naZdEJuf52I5Gn7pp5HqavZ5C8q+hIKvdBWh38VsgtZ0GzJ4SMo
Cab5XaNwWLenfvXm921MDFNawWT1J7+e86rNviGqhlEUxsgqs+8J4YoEDNVgv+UK
cbqj98smkKAifWAgK2zwkfk+wQaQtPqj0dwbfEBDJLshEyUe+alUaufPFj0uS774
zTjN6eYUu23vUMjRUeGnD2li6vnxQV7A928btt9snX8X9IgzOMM65hHJ80fRBi8/
Y0C/pFMVRG3d5b4fhZkHUbMtjlfQgbHJVLegvLzMbElK4NehphcQ9rAYZv5fkWwS
XyOWDPH+4BRT70q+dvf4NcGlTWIdEte2fnP7IXI1TYC8bSAoP8vmCHfMyFCfj/zn
xTZpRUspcflBqOQCAoqsh4yzp+y9iWHSRMRUWJGhvC7WhWIRb0rxJzH6BiXVGtM7
79tsLo31t9kog6WfAI2EPEMADiw3HjYO3oWpLyv1LD+esEo1Rwne3q7hj03DArLj
VHzSsiDgSQNcYnQI1LudGWIwS6dW4EWKRmQ1fPVDAnJzVDG1yihkidZzcJUrYsQl
hJRnCznkQlf9ZXeBL2krMceCIo73HBaAACrS4Czu5XNy52iYvRY69jkW8oxMkcdQ
1SaaRBwxB6u6EIthfIJj14/aiN1xn2Q0kJEnt86xMR/8Wln5YB6PXZZF/uyPOECz
WEHG6q3jGc7uZgQvDT9dFdDKIMPO7y8QYDVLlOE9SNhB9ZLfcV2pgunoqKcgtwUO
I2CNbnl0hZ2rsXtGFL85WaNqStyG7XFQ69EPj6aqqkM2WtaLZAXmUYsv5ZI7jrqa
pB20iNptkCsI1BS1L2fNepTK6IaAv27B/AGzrOPHTlVJ0sQSIa18wSfll9fEqkRz
IkVn4ElhlY1Mw+adu9vw9rQzaRQA/KopvzYzdE7/b8xbwZ0S3wKfboK0H8Ezt7Lv
E80rcAshSOCJs3Z1Tbg6fD3lsrMh/1j6z47OWZZTZrnd9YvWYb9ijxRJA3FNGzee
uo/Cma80tzo09rm0kQzNYrtHhsBbrThz/drlk9hWWGmu4hv3TBz9MaUfj8m7/Zxh
sk7ZBM78R9qtSUuUshOSfe0xaOiXlSusoKhhdzsCVOywjSUZPRecOCvy/qNzK7cj
1PtNPvkePI2vHNOMVQ2Ud2kzL+zllraFKpm4uqMt8Go+LwF0u05oK/nUg71pwa1/
LdjakVK0DRpwoW6IgjzK+srSb5yK42qgtJ0jhy268QRI9RP5COTzkJKXHZ0lbGVA
tctre0aj57fOGO+/o2uASmBS4QsYew0F36hD2NzktJPmH+bgYPfSjkWqAWfrwHKu
AZOzcte2FrUWIpOsF4r10bzFIWk43QtbI6vIezU1hfFptPg0g/KcD88D1+cgLzFM
FeJ+HH5HNV76/KH7723SnJ20Dah6YpWbnc5b8/ESBXNkxGzSSwYE6+xLAc0A4MAC
a6rOu2YPzt6fAcfD7aOmQzufMEWtNjii3OTlqS3LVMaRlbE51Ag0BZ2SKdUBbgYC
wOm1zIjy+jiloDuuehVvpa64nY90bK+p/LHUQLWpayLk032uOgWDQT7FrBT2ymuR
ANiLAfNTfSY77gxw4goJOffNQVkFyHYxw9jYI/mYWeRTnn046IF62OR1rN+HsLSc
xs4gxjaBx4+ORqMPTzmU2O9Grk8SJ/YxS8OvoP9gu4H6VZNssaE0cZZ8cp1mVx7S
14vpgJi+xIrWZSaAW2bYUtJ678minPpXsjM1JkZQV6c4wyW9p/+9bDaVRgSkxEGO
i8iJreBWaGUK4adfGZMJfAzR/0MGXyF79am6ad/bL3eDg3AEzApGuAX1UiQPlSEh
nEwHdD9FRmhAWEGbH9as8cRqWVde04OtxOjEg8Xu8M6KePBOgR1cq37Mi6PHmHOb
g6nTKPWo9grx/bGX5kJq2ll4Y+hXejVQkiyEbu16BLn5KAnxikuPWlClPN+LgG64
4Cv0TM68NhJCE8O5uBYhJjbzrU60htnHT2uQHay2yqoWLmyjA1jkm7ZzAN2hM0XV
Lik/STu+mGqK0fS3MoYwCP9Kjkx0y10frkWrgGY2fVf5FQZHMCNRkbXkcIFUDa8G
9My9r9ufnCcob2+Wji6hUAzFmyjuM/ZEqIwbJ7YAXXefik4ISZ4CfSVcEnjR+G6I
hQbUjSgMvoEuHFvOjvretWbWfI+H30nXeC++nymgPaBDgKLNelPpo/lKGm5NY0qu
OMNo6BNzAxZKJpg4yD6AfnksukZGLDtdlZ4HfwpVa/jopyPLrZqF/4OCwS5jP6C+
khzchawTk1l5cBnbJcBZw0J/4HS/hURG54g+fMEdutzl4hRXLLYBNsV9JRV8HiNE
9TlA99bAe5KtQyYnQ0fQ25NUFm+0Ni30HgE83RWTfNFmXh7DIU4cysO6L02pc7cl
ZHMH7WBIaYdsRwgaoTminwqvTqhM5Smu+3gAoHjOt7s9k4ECfqQsVjuCwwM+H+65
`protect END_PROTECTED
