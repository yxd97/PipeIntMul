`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvSA3PB/r68UCEBWnpsYh74NKTcA4711XJgizzpVQsnjpUa3xReIib+2LOaSvlyM
GQr/NOeldSPNQIgYWebiXySuiQ2HsaE98Y/taAe05NtAhYcNLcxAgUlyF4/LJTyZ
Y5UIBidcBOfCwEa5UnyogRouo0G0TxSxnJM5MxsCgRt64Kt/2as5GyGBivisBzda
pXKza8PPfq3tmEN9ZGV/XMVtTWtGs1jlIRzRY4rE0SpkhJTEL9Ny5ejbrfeQU5Dh
8eh3mrR8dPuA8w9xJEID5Z+yohwgucmFcapLx6tPqmzv3bE7t7VPLKH6FNyiYHNF
diuFkLGFpe6Xe2htpTMqCqkBubeI/NfrgO+1LFc9flSmpuOZGG+Y+pFWz2x36MLz
hFqNfDm0GpFWacobcyBR3YKozCJJo7tIzQrKLuVEZXjbTGQVcorVlODNx+JXLr7P
oHpcfyu8kt9HcsMdxE/T5MXvF9OYKk/R4uKb49RRDLVAizvdgNfMiBPzKV6PAmLy
vTGyODxOFvNmWdnUAo75zb5QoVAElx0Uf4pZAnIy8J9vLfPtb9wSRCIkP0JiXHTc
mdxYzwCv4E/akHomiDgYv4U107l3ipzBEtU9OSEZny7tmHbo9Ypmql57ryLmphOy
K4OawCel6vvUgqxpYutRJrvrtOia5KkAluMQRgMBLUMnOWfeOsuPAnT0sFAa8UwZ
8sZmPjBh2zj2dHofhn00PWeAvYLoUcLe3CWDJnciSGVmErv8ebHYstdgaem+Eqld
W+vUQmMdymUuTODCEcVkMdV7WYNm0PBATwJ+gZEKbniIyXFUksTH8dWRyapm2FS9
YOLYmTbqS+v6sHVF8ZadZwu1gFE2C9Bw/YSwohjNbGO7X0419bDT0bTUKLOLQHdb
t5e+ObcbWxkT8u5NquO9/q5zQK8UcT+Mt7errhYK5cqZxRVY9xW/Hzy+lnsC1+Rj
q/nyu2/5clLDMv8ia/CXU5IuhTf0x5oif6BoHcR3UBshcLRdDyWsLS+uYpGvcvMB
oLUA7i3AmN2E68i+nn/7vIq0fRYc7rEq2G+E9nS4WKZ9MrZ2pgzrG6tCG2Y6eFUd
Mz601Ek8FYNH58KS1PDjhWq3lajzI3WKzwRya0o2MTvdUY13zU0+IBy/k6LxSfEg
gjl6uZ65PQOXIHlS4TFfzvzLdGDaygGjNV2nG7hKR9WtVMZNKMgIJgIrD/r9en4H
BPWM9faqtqtgz4xxyhSfhH+gBmzAUUO8UEfEopgvv6TSlzN0YiNWjZiAtnoIG6/w
+v/6umS5JyzPTgJNNZdlip9VoZObyQOicw5oRhuugq1gJF/fHlbpsNEb+HRhxPLK
FobxqDOdnm30YmtKR1EWOVeJpoU1CpGeELvFIFM1ixYVUTS3xr9ntIZXeWMOtWdN
umrbmEjsuZtwQA5N4hyLMh+bkC2wgniQ7m2OIQwnyR+YCe6NWrxSNThiKfUIassa
KooxhEIOLFcgn2csutR/Gfrvw8h8UuwlAiLIT8Pvs3FNRnKsF6t0eE1z2MQJWKUE
7ioUOys6FoPZmRW2ehqSPNpe4IWeZvD0Fg0sNJCDy1LJSTQFBlMzJ0T+n9oqI70y
Siu69f7+kNBBi6+Pc+QGNf6L2J2hkjmncnUZuai1b/srhlMPEHTAwErnL7Kz8YeM
Ps+AyRLzUFE1xSsQIm9HYUflysjM3/mFJB/LlMX/2Tybe5qH9e4CuVqIs8Eyfkve
Sq3HpAUbVx0lDAPbhw1jvrCtv9VhlW5sKZpDg3M8+TYvJ2DV6JrTiBcvLDVuTvME
4X687zeMxRTM52aIezwDKDiOB4mgBGXtT4MBwwBM3+Y2sqFEWPQQO+Tk+1vxLesU
S/7NqOrY6on2tFNWWM3lgJ1Ya7ct4N6e875JyLnYDZfX8SWj6BmxlcKNZ+QKOpk/
KrX1u64b381/+MEtle8Z43Li+zVM9cT/HHXy8CebJFBhHoQEfpYMFNlTLgzZ1LVj
sNJ8pkMO+rY5aR6E/Ok0LYw/IjBuUUlMM2D98DLTmF0H4pz5iE9c3M7U0d5c1UW7
Q2vlrkoEh5jvd/sY2VKhCD1pNmt86Mlw2ArI22OppRaAmGk0TtpX/61Jv9lUt77N
6G5JzH2F6ktDf8YykRjyiayZWqgrUNWtsa0LVTiEuZpZkxW60GhAQgnw+j3vJmPg
qdIqPYZPTj6w0zhLZWKvTS7YtUrgM2ZvJlzY7ZuAosi8pSRtXMnF8nHFYIpBj0L/
sBs7WiUrM/sJeOuKdQWLJxB/+r38FYP2Xbw3Vr/tJ1t1R1Eq+hCkD6B/c7+L38K5
uxCpVGYDwjz3HUpWz+Lh6ngAzosUX/JPFwkYrs4s0REHAI5akh7717glZWoXySSi
/bpQ3mkU590D/baoRhlHHWSWD3Oj6eWtcjcggk/thDLZYxHpXGZeFuKmCWhx/hgx
fEXEexqVUwzvgrExePVjAxY0QsC9ZdwabT3rctU6h+9yy2mGORyx5s31gw42QmX5
yG9TAFH3lBQ5TWbj5GMMIBSa6JhZlB3bU7Gzc2vkLg3YdsMnAi+k0QcRQGBBr0Rx
w9ENY14jT+Iu9edX+XDtToFnzG/CEwQCA4QPnAeECEqjnUYPWnzMdHdzwHH2/yYT
dUgR4CijkzAwa/beFSHqlPCgqNX37NtrfyP+ej3bIkXI4OzCd4U9dSpw/41Agb1U
wE5Ged77T8p+Db052AVSV9sKzrJn6LWZGAmt4MpUAAS+5e26XOOSEP2nuSf4hjjc
/+SDtqSvwnzoGrFtg/sHAPKfQBRXrOTooqLYz4O+5PRoKgjQgi8pVXPc7o1KvuNA
PQ4WHwOTUUiW6y38gT6QbzqlaVLT4Y7JAORg82Ovx2uUoo8wMs0RklTyr3Z9hPEp
m4xi7mhhq645r0qN1AoagvR+Zn6E3RijOOdIoAbHjg3AzVIPqn9o7lGiXWi7qnrn
hA12o7avgurnyqYEuuZhGgvp7a33sBJLJE5bikwoI3FnHDgi5pr0Iv8ajVuHn9Gk
2mWlQigQvAiBX2kQ+KQuoXaepKGC3GlQJfQTnoFi1yJjMLLXY6QQ1vvW3p1mYf77
g9X4kKKzmWUWFspZOzOUTtL0U0rI9Nt1idTckVIfgjFDG33qVfAh0FS2fKeKz7Tp
mM1L9v46o2CslO3VrzoDhDyT8/J4hwfIgNGK1dWO+9xzBrhEpmyWtKcoHSiZjx8y
wKqk+TEboCqdT2ycXF4Vkv+mt6MofHea0ig4fe1IhFhUtbzjMDtaMEGeCAYneZSZ
FOZCE6whjxkr4ZQCxUC6zRVUDkdIIATDL/jCaZ++gRfN8pZGAXy1kbPjC3cAuKfv
1a8HHt0liekQtoTRXD0vlG6HQNJaKfZxpKGhlIjBjoYBuE3rh3u6kMiDvE6GJ9o4
KRiv5Z/Zi8L3hCTKqg16x7Q0Y1UUwXN63KXxRknW+F6XJLVz3KQUD4A9y8xeQkN5
m9wSzGkRGVxSejUuOTdL/clyCn3GeQfdqI59qNZsLjaA5DHIym+H3knq0B48hjTQ
cokAgUeb11oA26vyh0CJpZaKyeMJPFoT2PSQxnoLGH9zCWmusnsEuha3XU5am6o2
155yHur2D8Jkq62NzfmeVGRUpkAUj+hqV3YcYo1ypmqjS6638uTGSIoz57YDmgb3
mSjkESwqk52wTORi5TtmErdbs6KF3Ytw9HUzTNj4AmwYvqeWgGIEs3gexKP5j7cm
QUvquo7hwdpmyfiete+T7KkMxGssYUE7pkVntl6KlWyULrGKrtYGzHCPGpm5j2Tf
cVcRFCmsuLDW4tdJ1zlcaNoT8jyNPqY5mIrKzcaKmnhOIzDjRScltZUmQT2Vo2BW
HvaSIwuKLzp6Y81TQS98eoZpSRTuV9W1cYMWIAb3WwQ7s6KarHrJlLLcpaMXrDX6
9aqqrak2Is6F5nO1vDcwBHcf0ZbeusZLVXN+zdJHr2UujYTvEVMINU0hPgVm1evb
RKMHbmA8AKG9CMxWjpq4pvg1sSLU/N3ayJt4HQ2C8A3DGPHFPv5vpR66RWw+U9FC
lBC4xuoSiK8jGRQ5Sb0x6dzcGiDbAW5s4ARUHiucxoLC2X75uQl3HlAfpt4XvhSD
XmsqYISf1J3efbuV/uUgqGb2nagczaB94pvxpL01RhqxjSp75yMN+XRvtSKb/vX0
Uve+klhQxcbkZWZo5q+GwNxP7Dy7xT/Eljlho6NSiWnDsHi1/p6BrNL9DA0WT44g
w2daldc74PgfZplwyYa/vYqimMNFWwwbRNxgyTtKU/yt5jvQm40E4bOnBIrbSWZU
iIbLhzuNAo+tNeDm5wmsMfvEhN3YNs6sqI1hAJ7vCgPAag5LyNFBztycxlB4fC+u
+uMeoc08ySn0+FvzOIn3xS716lyyabxcPaubeNSC+5x8bbtUbAPtwqCnEmPaaWfn
V6dSRvAj6CVeLvZuTExdSP0AqmVSgmnirhjXW6aaN2NrmM8agpoUwEgtEXkdjDZn
wyVuEbuZCFFLDnQzFipqUDMwzkRbf6mKVjTDDU+fl631p38RoJ1bZF6YCXecH7e1
SJsv8eYBaS+1MIKPxtVBNwI2urvZixRYFL1+d7lcV9//gkk/5DlX/o8nYdugeeoe
shCjkBB1d6RQQWUViHV649zVbAnixtTkgFeantJMp5+MR2c+bJu+gkKNT9+4Hvk7
KFAiUWW02cjS0LAK45J9QWTnVorS0dnzNJ5R45/KUDOiFaaUUNdgplj9oamwEFkE
HexoAjYRW9SLKds/9sKkJzQuCFENdYQQcE7kQzknMcjUf5XPDcR98RVMPCH8thBF
EMPWS4cXhu5DmOj8D6IakCo20Q2RHlmPSDyp/I8UwXtUWVohm2GWCa10K0rXwvkP
w+ZD/bris5Pmsg/GuhFvr1nQl348v2MFgjOb6qtJVLAOoY7t/U0R3Ozh/8NzHH41
mkmBfbxN9bIbV0y34dK94DtrNrECoWZN2WS+zS8ISSjOuhBmFKnuPrfnFEUWudT9
sn1Lns4EBT32zwiGnM6KSlqgux+3CurS+BMcu5lRUGtG1VGvFERh5cgHD1r+BbPy
Ufvu5xaRsQEYO55sPtm5lpFVk4xiBOiFIUxjMx+VpNC3RpnwRjH04+5UB+nehHPu
f07poIPLLLCQrs27qZg5UnvYUsf9SjdJsBo5rqGF1/1K6WDx4Rnmb7j3ctwE38Ie
iFFZ6whQau+wtgFt4HmdIMT7IsMOkSvwsK6hKfC6GlRPuc5Eaz+g3E6Zp2nTlWBx
bgLKwlrTUV3zSku1g4Ul9HcJy2KmaRuc4Pf9RayOfY/Psq44kcx+wp/S+YlDkK1P
H68ru8LX2/DTY6+FE6ZXO18dtLysjUZiwyKYp2AA+rFj+nQJSSiZD2PEjmhLZcvX
06QgsHxnXyHuApsT6xKWaRG9B6F3NIQXThrBYL0B11SiW07bJBfI3IqoBsMOc7Wf
TK7cZTQUYiitq5ifU4VHqqQM7M60HJm2iUf2Qht/E2WwbEO5S+/qh76kxGWODD9h
OUeEMQ+PSDV1YcEG1Rj+jJ1fn/ukelJ2dzXKgA9xs/4aZZbEwhfOJEhLOmWwiU9o
R6fXlf6ThsOnvdiN23V5z7CZbLltz4NyF1Oo5GtdhnywA+9C3zgmLc+2+jkDFxp3
d5s+aa7sGTvJSGwPd06QDwwZQG73klv+Up15wrNEDJ+aZdl7dIYWfxnYpGcK9eND
UI5JU8ZTUY3WGqSAJQ8S1i04KRzEPUx4PUCU9751wgNJ+G+oXXa7zMVrYusdl1IO
LSpYPdVJXo3vn/Fc/moy8cSDSoK+UmNgnot0fJgkbNBs7wCsVF/yIy7eupKdKpA9
5+iQcEan/hksxnEhl2jwa+Lo8oKcwdoRNfI2yOziysdY9nohBGBB4KlMrBmLCoKb
HirCzh8Tg99/KO+Dzr+DmKR/ceUB3NZ2K1l80pXhHC5VmgD5IQq5eClMuVQEiXlW
JnnqRxn155p3uaoTDoL67a0w1dBn5yNDb6vhmSMhWVv39YxRfjT7tnZiDm/46A9I
sCSzYw0+nBqA7pB5jOIb1L91LZDnHW/RCN4MJTJJ43Za/YYxh5O+wsi7KjG3CCTW
gOX8YT27d2kYBa+lTCH0kfBpUUgZk76U2WzLR4TSXyy3iA7umePtdS++0z8PtIeX
O6RaKMbrh44xOi+WI3yuJNMiBxfQCLh9Ww7QKAAlhKtKIQG9f5jZ2C01jMIY4+oF
h7h//EYjNjyv3S7BpOEtOERNMThVTxpA9+M5bgCNQKKkyZgPWtRu1FThDzS9jLNP
u5jfwPZUI1+oiz0+n+9hxDqSUMEErEFVhC4eaHS3mEfQvvtjlf0vMCWWU2OSvgHR
fZlUynxkHS3sIu8QVGJOKQ5N6eQjRjUWZmkjpBYeX3ucUyML9VOsKkj4hKclEJEN
k7IMh9NAijpA+u5cnsWRHQPuhUhIY5I7E0Sax51vsRKiBFOJ4IcGZmRFeM5pFd8J
LFokkt6e83bVjDMQWEq05X3OxAShjt5jExKg82g1ewLt6lyxHAQZGOtwgI5yVdG2
UaFtu01exMrKiKqzULsO6DK+crTZn1/OecYihP2PeH4wcvvqimZ5n6eeKVi70aPs
PrRbUysNd54zU2r77A+lKGtbkUGE6mykxHeeqnCyB8n63MWHHVWAQoJJLs+kfD2B
Oxd1nKIKOL3TgvduJXHtvHwh56AIVfzyoha92Bsqui97op2rzkHkn5MmXoBb+/y/
/gVPe0FOkUvznjhB98gmWS7EPGsyhgXgA0Vx8cVIKDqKsYEB1jBg0ZHu4nWhtKu9
MMVgaJd+6uRxp45JDLIRvcnWIL/3HuINDSlc9/QE2R9CXy2uExi7wccoTrmGdVZ/
kZ9rRQGfpCzBTxoLlWMotx37enwk1jv8H8vSZH/EhQbc7h4im0l0VkI72oaodQJA
Kl96J1RVrn8Je78zOKtNYICKThFahf7MBlQkzTTSjI64YPUw9LV4Hw+ONa0XgUOs
QrL4P+Y3yopIMHc/5M74RQxO/wrWzBYl+XJtRtlD41VNyKH8MWgZhPgXUvrxpkJN
/XMaeym5V6yHswMuvbf+lcujNert+zRgq/tNkcfdmTiMwKebTQVE+D9M8qFEyVGv
/8TwVsRbJGodbjcTHSVOVcOhpjnjQbdSCRKYePINvNRI6JkyFOucu99KK90vfGZu
xtgXmuqoyN/VwXtb4W8TOkugZP/cJYkLJt8Y106G5IgUZGswML/VLKCK4FQkIymq
AwkdFIf5MMkfPz8ExLyOc2EQm66KKYM9A8cUSMDuBTXOT1mq5vYDwIV5qslStoM9
4WpFEgfJxTQ3F5Ah8OKKTWciCp+YfNVC6BTMnp+i0qurzqj7sy+Sxz8apDLam737
ZfET8++RTaYXWKnS7mr3FlpQ/DT2Z2lVsMt5clMIE8SQaohaPilVtW5+NUnGkXlF
mYrN3FwjnenfrUsgrn2THTYFv+PTlFmJnTiyde8ngTjrYSlf5rx1Q2tNu++lgxyK
Zm/gEb6QvhbteKOTT3S4GmJqu0kehG6oFWesO+iFlmE8TQbVxju4uejP5KxhU1cq
Nt3eOwCfAnSZfesE1T5bojSURFeJMZuwj5WY9bXHWlBphTcEdBebtGLTYWucz94R
Xs7mDAMlC9wxoO5ScfyaKEaM9rL2T24tsjRetK4L3lawfRRFJYoH+BjLDxex5e99
nBBbBxwV72symARIWYAlS2pim973YrK2d0wgTi7I3IaHxpp7f969lxhkdoMsVroa
tQlmN2/zxXN/7ctkApwJfiLV8kjz1fK9s32ETV1lOjhRaX5fMi4Jn17t013PDg2u
CW0lM22kQz1qHxaNzJGSdLjL2y4izxERyCK5k4cXvZWdRZedc7BTpFRyXxhSovnH
jE4WfLttTthsz+4G/aJLKof8yMiZl9+aReAOON2i8Z6kKq/7qdli94JuWakkB+tL
RAOP88jllIxUN1O9Kb800yBCp4XDui3LUP6zMg/02MfsRCvsldxs5DRqZX7Jt44N
lpRbW84rCUnL7bIWDADm3m6H1KgZewN6lJbBjOKR9fF6prOgkikmjuqpNGyMsKVv
N4ovlnz+OxNWIoTSMkiZHmtrCh/nL/QYlC6khIV9koT+z3Mi7Y9J2nAg0PSXqcyW
0zMqEW1viIfsnzTb0dAz1IwRx/Se3FRyJcHN5L1fTnExwgztK3BsPDEf/aduyxwy
Z92c6Rjm4Zw3g7AXw5Nb5OzN+mPZ4/aZUuTcWhkiRxOF4BluFm/Y6+FmaLERq3jO
i98dLMMefJbDTgmUgOOgNdRzk7UnCXgFVtjRT1lvtdQ0I6ZwqWj/uraF+dqY0bs1
5kslFlSfwWkONJ8Go3ws+mLT+i1CT6i0AvbcS9Tywu6tZuEpEsP4/IUPvW+xPsiw
DpGWLL4ljAQBQoOiFnw8S5E1LgGE5+SMFhWPr4fKQwu1Q6ywz4JvaAPrmlu2sVuA
w/4k+CKxIbMENo8yxpQLGl8XOy1vlQLSudgrMQgtTEr5or+xyaVofYHU1Ij9E+RZ
HhrFym0mLH2ZnEe1sZMcVpBZ4/Fzt4pW1/YL6a3lcu6J87escz7VeUaXfdftTWm6
eIt2b7mEJkB7IftVgIvgNWOsDbqe05+k5bDxiZnJHP2f94XdrNJfyjVuh3kbhA5w
BRLXwE/t4YWcDIA8PPqo2gki32YT1YrmGAlNHKnhItj2KvIUhBDHvVQi8ywT1LF+
YW0hAtsbvLA4I0UyGS/nH0Tsux/ZYuhA7nYtsyggD/Uus9bSOdCumJw7x70Szio0
f7/vtG8XU6UKDkf+WcvCPE+7pbSz7Z3y4BJPb5IfgQg8XydtQ7uVq3Vox7Xtz0p4
JT1POsvbAOYoDJJ9Rm4uCXvPQyMKoPZDAk99s/ib6Q1tzQ84m5aAZYn9gRZTAjTX
j3pcbSzzY/HaYJUcEhTqIq4Jl/O0neWq4tLE6zoRPsAKjQHVPMw7Ka4yx/haudqt
ujmjtE1futmiMaAK7LAyoeFpplJXViiPBXSl3gSeGB9bHl004P+3wqTBBcUPUZvc
zeTuD672kPQsIzKtGoKPP2eeGRVCCeVv2MiqhuEj6TICFgQu8Cd6vbsu+uAvYnEm
MT7dzDUHjzEzR4d6EX7n3S6hiWUkGdG+CIm4yevjzY4bedakxcn1YAYE7ZKX37Vj
LBO5s6MiwF+iwsLOrwlDXD64d3JzJGtRYop0xfLlx0/d7zPwQbWJgKPLhTkHzSj8
AZV9PBTUZA/yrr9PxXXU48FhnOnMjXpOB6hCaGxL1YvYD3kJqZR06n1/lCzdXmHC
yr+ObkU8EUi+jiHkXiUP+qATzJgt2eKXIIX24SXGzfZ/iyD4FeimVZVRYayt62dQ
/fQ4DOBxvkOBHs0q3ZmdY2V40JcVfYvR8Fjr5uEJ+tnFLyCVP/mrqmc7O9IX4R7j
Y3WiJOskhW0VB9MCwUvmlwv1gMNHIoe0y76quR4h9ytAUNKY7uP7FEBdJtuE/xUW
gW6AgvC7K8t/bNkMLx/NPQGaBDDeXhKaesQiwsubFEdLb2E389T8xKWvfZyQHnOL
CCTvdXE8TksOWBerNIqMhMJjE/lqJ5coYHsiiM70ae++DS7ogky76MmHZyFwPQyq
dKTd/ddpnoaSEfLAZ/iJhlxCSoV2538VLCieRXQnXdvrwQhAyI4QMNY+0DaTj6rw
zb3jw0VtjmgqRjakWJgTIu/LO162wvBsVFA74xLyPHW4o1L45Cym2YiirSghf58p
xeDMBujNHqXxU0xDQWpQW6TayNRx29QebjAaSOPkTtRQlnU31DLtZzPEoa3WawOT
IBBYwluq40AOTWJot7+0obw1aq9HDC0rlXMgqOVBh3OehPdIemvPp7NJkSl8543B
4VeVjUXIbantw666nrjh9x43ddFnkwvLSx/mMGoG9uDbtXJRD4ilEF9ociPOi0Gn
8P5xSjCFMW/lNfAVeeHVGioakNhCY3O1xMVcFniQbpngPswZE/vo6VY9DywSY0bW
r52Lb65DhgP6HA3aah+vD4dwRVf+JBRSFkMnR4PW13kIXQd8OvG05jf3iUiXznFH
T2RxxAN6S+GK+6MDlvrd2dHSm0Cib5Hz3W97M5EPRFwUtQWfiwmQ/erSpr3r1bFP
nHWSVpzhmytLvbBfNovL0KotA+RZIYkFy7WDsi/z525elusAFnrEtVI8Fi9XvJqE
VLS04MXmXtkhK7wROFu4H90aE+I+x6r7fJ0/e6aXFtQltJ/prQRngk/lq5YOXPna
4+9g/EOiwPvxKJ9GJlKvKC5chT3g2zL7ND4OU+zKaDrqUidhcDlh3ecH/xMMTR8v
FuSUf9WeOSPodHCq3FRbakNC/aweDft9P5mh6RbofRRbT6Xso/mqOjIADnQTlp5+
vfrr6Yjvb1shiXzszIQl4V3Gc1gfVK4gTssMeOd9o6ekcbOtl3mOFZ6fAlWSya+X
Z35kiCjQSl/0eEy85g9Dzxfrnd4myH7MqMf4QULCHCjQ+EyNxcmwzqxZfF+SZAyK
SmRn5MgDUjyGiwOuaecnaaIsd0eJRe9iBT5I6r86RoWFCKvMILH3u8OZGFzcxCyX
dWLp6MrRfaSXewL2rEgwqpx2eD/kxGlho9f1pUisakCDjeurHP9xuDbJE3Dwwvko
dFXT1oqFSAliOhxMsaTfXAuPgYpj/8GTowz9qETbiJsm4bZWKbmg4lcTtcxf4ltF
9e6eSQds/djZ9JBFZKVD8YTSExsGujhMn2kSzxZS+GmLj1XKYxTsGWtkUFTTUILk
75FZP4ufJLVgFo0nW9Qzko/i5a4Jg0Qwv+X4Ex4+hX/Sdx+mxKY5vAqutmXJ7uQO
wn6zbeQwJ1KK9QJCJntjIxaOzWaGrtNGd+7qrZLKj6zYfgKDNDqKS7+Om+e0Sc+9
eppDEGhddJZMbrOeLOcuVUN6g6NeSixNLZJwmC+rSxNjEvvWL627mWRhH3JiPvSU
4NMEU/Q91sBW52Y4y7ckPZx+cg39tRy28zrJAeYy8Uz12/ZRAh469VTXK0MWTBbb
29g0R0IIoRXXM9nh2KqiDDC3WoAhi4BrpdA7PCnuGSz2L9QH2iNEUObuu2YoE2CK
E4il8EDY4IUkUwwmaBxsOO0TzXlrEFzta0kS93Uj2BtrLzP+haRTuPW6XAreILS9
iAQS37XDwEv+ilIt8JVh8Zj4c9izWU5FMptfBPC0TFAqAIeOlSLNLMNDY0UamFUW
iGCzf4wU1Wb29Awmpip+uVL2g/eukIvF9X71zj23jso4IhUPHWjKun7JcaOB9IPc
W4Mg61/1d+s1nZuA9B5pmt3R3lfyWuD2qrq1RZAYLIATWiIyLfiGKQQVaTBA+2Wd
xbveK3yaN3vPOYlZDRtFPqLBU1q/YqNgTlCxopBGUHLLI1RUmkUz8sMUUrEqTST6
6c7RPIXE7tGST8df2NalV+cg3VpVbbyd1nBAYlse3unVTDKXPiXnjKPan2TmSJ3x
1wyglw2Ma+BbJ1mAZ1dSu9S0UWods1t/F1F1HtwRe56T+dLC/M56gjWHWvJZU/H0
lR/hfS8EBw+Vt//4q+AGZEeAzWGwp3/RsTSgAVTczJetVtfNE5AEuXufbgqzVf5I
JbKxdwN95B9hMwM4ZeSuWMric0kGE7dc0bmMqWy/7a311cZA/zdd6HLs4paxpsJH
+Ct+Y0fE2dWJfKY6PA0QYRBxtGSq2oFppDgn5JfECdBjy1pOLhfKLMEt3cKu1iJE
NGrNLCCQWc1IGfXTAfMcHF3+AbXdQRBTY85VSY66cdSEDVstSBPpvhOSag8jDnJX
Vmj5mvdWYoyKxXeBvzMF4hP+6+qq+LVPtUrY4j8PuXbu6RTQj2apKpsONPY3DE+W
gsUlbQc5hMCnUR7YrO+crvWciKHbLOlTDE9bFS8vzV4St1E5o45sQk1tRwa/C+yR
3muhA23HnU1SObuZ1Ht6FwKs7vI47sMFco2fB9CJ8O/yctn4mZOsjOHy4sFoi030
dZ4oDa2e8SutAlXbm6twAdKdZDgwulk/gly6flKWlPqJlfZcWJnlVVmIHn/H99cR
pVcHevMtQw3DItH5b/yld72OrXAXrAcSZmnLdZYuMSgtUBbaYKQf250uklRwBUzU
dkwn/T9MCnEp9Dw1fEXE9ve3P1SwVWKkvnDnaUYGeR6bqo94PGRFJQszC8bgIyfH
0k9z3UCsaUgN8nRRYJhVIj0kg/74gA3/F9T8pnsKO7IwLqOk0uvEZmqEK6Z2NVcY
v/HASHNa6+xeUTKGPt2u3yowGyDDY2Lm0iqstS2o4DXHR1vPAk5k1LpyA2WSitYz
5YaqE6EOSDwrYF4c9tCM0FwLYmnCiUbl4krPlbWbWuBSgb7l+afT/8DuzD4y75nS
Vu2Fzej8FSsWEHQeHI6ANEo1nGA6B2fUQk814suunqW1dzkTBJZ6PjXKsy4tk2Ug
TOXkapKemhamMTqLMl5U0fZ9nWJTzCbYzfARGJ40J9lH3b3a7yybqkXBNngRRBAS
Z+1sForZ7K/SgRCU7C6jgdRBXwWEpLlX55CIXJmDQ6pZV/wMcfoLYZ+Abos3yKZG
7J8Pok19TQVrRjZruqdatE3izK0xhVdzWxxhE+QibEa+ESJmfNMma9LhBhMKjWbh
Eio2+p/5I0J6qIdjxc36ghALtu/uPC1UoLLw3UcVzDeBqKVU7pPB64ksf26s5nkY
9G2Fn2QuBpJopXIpP9F3YpcWDI0LBt+Vbz5982iKFEaqbhpvSRh0bXZsOinFiiZt
DZedD5FRAArqg/2gic4LMe0gAclOyGPNtQqmtF3Dc/gbz5+n4O4EQyEYodDazipD
pQuiBhpX9ycH1QPhqV4tc34PcHTeey0sDmQ5bQW5LeuotCQhjJbTgyPNHngU43C6
Eo92QxoRxUUNTh09Xe4inB/6MkHxWDW7dnXQArR7FC5Syb31Q777V8dJEeA0Tepx
20uq68xMgeGJEULLGuM//MGhaiNl+HqlKgfZuWW5Zj1XfZNlpErlQyjbcoK/D2JG
kg6CjDxetXHqFX8PX30NCJ4OFD4zwAKHHOM/MK8LclZCzOTE4j0weh4syWML1hX1
5Kf8H7+Wq+vxgwovIyxQoo0I+CSsvy8ho0xXcQdn6txvNF/MTCDnHPSIOFKeFeOt
dRP8fD1jCwBoVvUnCteaTrCEkOadF0Ty4xi8FaRICtfDBg6oUIUHRZyMIQZJXbv9
9mRpCfaM1px2TEA8u6Bn7UeZcFqRdBkH2FQKq/FEKaBHcZqYCJMS/EddjeaqrU9E
V/nCrTHNDpgndyApMGj1et/AcUthcuMD6XiCGWUiBcIqvDAZ5heXfgFDsNxDxiiq
gu4EwxmK/rYLw3XFcTZ1UrzeIb74Tzo52PZ5NX9WjWHCnjLuCjY8D2XV6DpnU1AH
oSvtxgR6R/uGGdoswriZ4+qYFOLYpWqow8kcUhStPUljBKutnoG9ymRqaypz8c0P
zhanHh4XAe120elluVhgx84UYmqRD8RvBDsYbD2/aI7W4lGk0jjXVaSGRE81lCAy
gCSZoI+xXzbVwn1Q/Mjl97JGGfpFxGmXoOK3eMi3qopY4/nTzn46BSILMH4BbEiU
YKf0Zl43CCjCbGvhZ754d3MP9LKr6nLUjPRM3oE4TueV1gpr1KXUjWndtZgYlXOj
4BsUGtk/e0EJrToqRstd58Ws/iWPc3QpVOP/4VTi4yKZDiZ7f4GfuiaENI7FdfhY
j7Hv0+fIUWOTGaa7vZoIIOdy9JA2Zdo2K2EcBXbCtWUbAs3BoTqgnVBmeOuBjhex
ty1o9M9pcB0T5YtYitfUNIjJAmmTKZEUaOIfEihcIoabRqFAuGebHcoDJDCd/RSx
w9FIObVHgQGiUw7i8YPlMPMboiz6hnkJQwluZJbz7PFTCXHp79XlM99R0ISpXaJx
VFkSkAbooNmkA5KC3ix5hEs259MGhPtku5LgKzfN0XKNw68tLJJv5oWfTlPseboF
sza42HCHCZHXalUuuk7QtUC6UGcotOJrPTb5TRlb0KEjc7qn1u3vAkQjmFjmzQOM
hSegu6lnMSTCKOnydeueYlp64vVUgElsjKeT0xg0ablymvPArr3CJzuycwRfXAtn
s1KJiaUB5eZ/j6ubiofoK/rNuFyZnYWaasrjYIfFLWoBIJ+szcIQWlaV8jL2U9aE
J6A/AcjlvfhTbKXlEcfXC/eS7dMNDm2u5FBjvNrTv9dyVM6Pr3T9iH9o3VuneMRi
SlAX8HHM5/2eK1LZk/stOqkmq4m8cB1fMWDNVUaj7P+KP9lcADnsePp1oHGwHYxp
L+Q3P36ntVqVaP6vmlC/RQpRghW6YUJEro5M87XPVV1UZNCwLkOI1E1ofy8BOnHO
wabYEbbb/AinCsxk03n3tmgZAMgqz0+RTiPUGY2IUjfgBuVQR+OpZEjh5D6hD15M
tc5crCXHiZiqBdK7Ef3J4Bif/neV8ITk7tANfWMH0bZZ2VvmaARxb7AybQUbMcVG
e4dkVgzJgRtBGG4biYaHy/xu0Mrn2xo0et24aQBFm4bQkylAPw6lT2mbIfS/bvvI
ZWUk/L0TJi/Nz9IQMQ7MQtVKQt36FrkNhNcKT7i/urxm+Kf1HXTW3Ps1ltsNFfHr
BwQUfnIDtlxjEUSkYnxfzjDNNFFFO9cB326XGkVVpOu7piVQ0WOqYV6cKlJgY7dk
z8xjKGkXShVYHV0+QIAtTsXvZHG3SYi9e2c88yqbHMGP7EucP2sGdV37Ew1AeQV0
wkHqlbeaD2lgoiJeXFuabKNpBQJ/KHIAM6EhyFa4dUno+AzbbD93rTKi9Qmq3nk1
rI/Z6ph2UAyVopLzYZC+BxVj2wzDYrD2DfmrHDyDqykesF+VdXW4oKNu8j0yZvzg
IcvWnUUQSFXRjyTYRsIcbHT5YUfGI2AKt9rdI6bO+uWlU3S1cMwPotqpEmUHC9Wy
m0Z+evYAZLilErdLpxVUMpO6zVaqgYVpon13FShrynD80Oc6hVumQii++cieJXhD
Rb4aJneR3fQz/LyNpQ/WJ0ZdBC8UZwbZ9f6uXakbsU3t+7FZ/CNGwZtY+7jU8DiK
G0pJrRou5EqunXlhLa9rrygoxQE7TQ0/jl+HaWHXdpB1eIXAbMrzNVCcFuBSWatH
zSX5PPnpm1XNZXKphmdUTdhEwofCBCVchxFAjXpTSVQ3WRqtdJulvbTA8Vv3wa4E
oXJTyz6n6MhBZtd5qSOlKlUb8C1zDL2A8fHYX4diF7QbzLdb0BlHIapXZPUWDzEt
9Pr2FM5HiM8n6XpiAA2LgNf9+jxLze67Qg7CWYsKKFMrieuNgWSUHVqOIrq4CbmQ
qN5LSI6iDeENJMGz/Tc4SzL6g6H5sLtU6nhCRFUz28IH6qZQQuOGhdwIAo9QtOwb
Zqnw0WHevXm1k5pfxBKJVs6jov2RogBDafkJat9vRXHflfKqRXSduNb21DNFAAD7
ekmAwxL7PmkUHC2/wng/IrGHkpxMwtr2o62SPh0WIWOBFrB0qGxBRWanTu8p2ma3
f16GYzpSEG4hmjfX/BnY22NHAlwFLIe2+a2RUvJC2dE2fqcTVq12oKjck0KFu5HF
K2TqqQyKq5RQ5OLAB7//pidAWBZ2sHYkLR6CjCXoXvi4v+GOPVw24l1I5tXx4H5g
2NzjT5dGnBxLzKP+EmFnZaa/A7UCRzG4k1FCMCxCDdSFv7J27rKN+Nmmo0W2KVJ1
9A4LKZ+HMiUf/IfJEiBB+iUmCVIWBjEFpxpYqGiuMcxWMNv070ruZNmF2SjvK7O/
M7HfkKGkvv2R7Z5oAs/pk2+b0umpmDL7PaogNLwhCf4Ky4wyPqqu9MuS7uLS87S9
aEjaYRtae7PGi8XCrnl8pKTwvLegDzkTo2xBSCzNToCLU7CTgLsaYMgIAwKYcFpm
ABbMQIjWKgd6FpbYGe4xNmsQIxftKqaFh6ReQ4+RYa4ePwte1rTIXvfn1fSbn+Nj
U6Gy6AK3Bjj09Uyz8GTY6GboShJmzuLnLwEmF4yrSH+uK+X8KEis/D7jE10LBSzX
cWLp7IleG1YzrvSP0Epzmm6Cd8zGZw3v735ckxCQg/4RshUfkdPlkZVufy0H00Zu
/Na2RMuksiZ8iMN3+xUhGE5v9BVvmttpMvvPQbQz7qi5jyEZXurD5fVhxcGS6sru
eQLCSu4JLHzVfkflA80SL7PSRdn/Y2RA1wA09DcvSi7fIOaIz2gXIGtx5Kco2Q5T
70qrw9OIxEYb7Vk4DjIiCIEYB++U6796tZF3db08b3hbnXJajtV/x9l8FTtI6ziU
B9R5YcjiMO8OUUKmbyzrShSrvMF/G5SLmJoxhZg1MUIp4pvoCZe1JGPC1RfAsm0o
hBjgT01zJYDZvODR2twXVWuNmfSiQYzPqVmeKD58Z84bjQibR+wwJ6+m9mHHTCOF
4qPy9rz3fokNA+5IrgYBRYIM5N4MN7c9rCSe6vvCOsPfcgrJxq71Cy7kAES84UcY
GTIA+61q4a0zM4tPZAlml4jtXYydyK7nf3oqP37rV88Qj6P02n+ipSXJBx9KVN8/
vPjt0GEwVY8euNcciiYZlOLfDZxGSPqR0OFfQTCYUEJFucc5pJflUMm6LrghCtPu
oStoK7g+bsaUOaBo1in/pojA54BXMB3ut4X0fwiQ2ELvBCI2ml6/sLnrUTn3r5OI
/JbH9YDTQUhVTlGI482BAI9PfwPHRgsHrEUZZWA02x1gHTZYAkBILHD9Qh+L/qkn
zQ+0hQIXdj9SdcXL8yZOLZTFjS+yYQI/5hyuv1DWP4m9hnbSI8lZNeD99IP+aPNC
cW41Vmkdiko4IFe3HTEHEiGCnWVqdPcIYVHtR7gqo9dai7XpGPmPhJZVsQVmWCTJ
+kHTWOQr0Za7fpVb0M6yF13zDIcU/Bx1DpdcLqL2LZaEeNJuddzBcOC2uJVQnvXN
npaCYIf5jo6dAKmgDQLCHK8+hbBCvYAzgUO0aIip0JfpjKPpdwI5ZHlbs7WFxAXp
jRVK/UkQlG445FA/yMWOZtZNcoh2qEnOQRXZf5bkypIc3wc8RGKU+HuhmiM8WiDe
I87mQHkGQdTzJhIF/Hycgz8eNJ2e+q4X7GrasXWZCYFxc3VheaTm5bhP3nc4RLrq
XOSfZyotDig/arV8tsQy4XyBxbtb1snBMZxcg9MMFRTmKEOKjKnhuJAnwbpkwqJf
9MLKe0bOLfX8lYEjSQ4PN8f1wrrU9DUZgig9hDlfxPKNaHYU5+C0nbWW3PkaPTW0
bhUEoUE3Tw2a0hCyl3nrVoI5XuExH+flftyTlts2SYOK3QNAlOaa6tp6hOouev78
+pgrLGvlvCTCd8au4edKIKDiTDEJYele6IdGpsRPwB3/Y9WGs/E6imrD+VGhQaIp
1SxTAZGit4ZHYvkHhJ7C45OhgUcjC5GsTUtzs6h/kLtnW6KQXd45TxWbdGND4OgP
k3sZA0eZrnCnmRtLuTE3xj8BA8LNkKJSOf34auWLwmr5CBL4GVq7Rgk8SS9VXNig
nsfctToezRyi13Yrhag0MnkneUU+KVHwGyCmHZGkczAisWotKSO8P2mEvUzHdIGM
W73BgkRUZPoaTt4EUgDtGCNniOHwVeJJeOAYP5j+C2yZiRadr40gFK5voA9z/5l7
5fTz3eppyVYj31/0E2fMgR5ugv86FrRKi4Q2w2BOHaeUvzeU2GG5GuPH/YJVGuH+
6CfMUY3TpNgdyvUbemATdZyw4Q7t376UO+Dh8gZi5ZkrDj9mixqmRt9H0SoxOCqv
i1n5WB2IrpqU2mwlOgYGr6vEPGl+CNXamErHYOqKhkAly9nwgCj9RAxhPLYRE94n
JLBCrxvAveGZM016k0kJgoyS8/F1AcLIE7zE9RhYSFdOrn6NkyjqDVoVWUWhtI+f
tDbf+eRK3PEAWubpLb0s6UaEG/TDgvK9zWCUVcmwqnlw0Dj8E084vm9VK88eBmaX
LhCA5WRHaNa7MvSw3HVknXa3OHjf8ETNu2kT8aCHDDE95NWVDoEdIzDJsu9kfe5S
Cx6eaMkDVocf6q/3u2LYnJ4TAw61cSsgKHdqJeT8dZwae1Q6q+iTyCUcV4mRJ8I7
UkpwVaaGrPX53EtoblZxb2t/EYy6aU6gh6hsxaE3wsHpXMFJpinx+4Sg9Qgni+8S
drQHJSJIbzmcqfmmM9YyfRgTSoCzqNToNNsTwmnPBb5gitBZu5UTmDpepupNfu2T
vj/F1tInGrBlZSyB4Yi7Wk04+9+NWt/FcZX5UQumUT5hsUxZM+l73M231C38pPG7
s0wb0nnN8eDpdgycDZM9kvDuWnRNYEMdDm4S3DCkxdcch4hWUFqpyZDnqgOAm8vW
7kQDmEb+/ztQBJtShN2dZQ95+qR360gMBgJM8wscnfJz/34WWZE+4I9dKMcuBJss
A5SXJyFjS8xRqUgMVGe2aO7d8OAccf8EBjvCPnYHHp7RkHB0QE/SRru/neWyWseR
AF1iN8OmRfvplqFjXZCUqsMnfjpgOpu51u42qNzhTE3bezz8APqDOf55KD6A+6Gi
/7fAq0KOaZ/27iW1Togg/Qa9GsS1EiJtHFIgGnXz8htkUvNWdxa2+Zptlj5jo1Je
cIjb8qBT52TGA+PbT0n1EbZW+d8hKQubBunMcnOW2IyFzUsRw9vmk0Wtt4l03ARs
DairYwjitZ9aXAFh4Y/TtPtukXbnEzjKjfzW22zIf8DEmYZmsMXr8nmXR1UhNRNV
vlcWoM4rgXDrUybB+evZdGFJrLcoWkjW1fy1MljIENDHlAk7gbL2iACyXcTwDROT
JFB8FPjv/1e9vFRk+7m8fZQNO1tvVlpclaL6ZZZBu7nQHXB3PC2swo/4nNxi72y2
JYbL04nib2p/xPsjHt2H+icZ0tyomf88oUmREitZ8mAc6n0dNquphw+lNHeEspFn
6OkD4FQnmggvsNdogEJmR+JiJM6aN1WS8BAqJ51ZB8iaPI90TVPkgvW86dBIK0iZ
ZpHLBauqpQUcsnzTtgywKy7ro8ZnSW4itv91L4/ZxlNBbKES1PKhQyzUDAJrZEQ7
7qJVSGPP8If93XIqkPJetZ4OY1XmS/XS+IsDhmritj9UztbUprVgos1uCvxxHOkW
bcLzDqXTwXXWyh+gLFa7JqSnCItXxbPBS9b1wf2Yz1GO5cCkXcbml7jKNxaZoxTB
6XvjgWtA4lnxFvZ/k2pzzQYlNG/HjCb/8A8THAK9WtZPPApMwx0vHCSOamydsdgo
bSLd4zPiSzgNUgFkDlBz2kSoJfFCIWwdC+zMcSd+NJ+IuGq13ilfjGUaC7rwuhAa
5EkR7wH7v29wtzSh5MKNlXBITyHrttOqr7nCFn1aUgb3NP++FVN3UwiNARdBIaN5
Xtma0h8dmOjN4DWV50MAVwPRE/HDOGBs6KjRFhLDu3RB5jurdjdEoODcqDw6VUcS
P4avOD1r0aM7cv5//qnwOtJgt8gfl1yt9XWmVf/XARJHZ2ly/WcyDcGsGOyNmuJv
DicLAkabktvEO5FIYWIDgnoO5vUbmUYY4sWpewPD1cQTGZxZdGi8VCq+J4MaVF6C
ohZVQbjFjQ3JZyq2oyyzs1zomFn3i3t5wLgMRnVB74yjlKdH4+YdVaQs8+2bbPQo
yhFbyrlwk97vnQKv6AHtDTDziWb5XbVxsUQQzVKFJkpt9Gq8OGhdyqlO6jhtx+xr
DWvQoiWyV0qZ+Ocurakznr+nqe3fca06hOaAF8gHNwvkk2gXqNPV5AJBeHVZSlCr
xYhejVKzPfCxRviBYUyWePXeaz/8nopuupale6jbZ9DmGGP6V/M+hrJZfgStq40n
ro7tQ0fhqenMKhnjOxywse+IatkT45HD0QrORvaPIAAnemZ+SEkFkczDEkpVn3o8
aVN6/mtv+3z84Ikoj0qeYIa1gqWlG0xBIlwhhP4JTHoWq2rQYiyxlam+cnITIKhr
hJiGV4fcJEOXonbjhRP1afUAwrXGuRYf0RZu6s9RKoExZ3v3dBRZrqy3Xl1v0JxW
WGc9lN+Fo38k5Xz9TlUUO5q9JDEJylIz1JNHAn0/ro5mEvKho8g+QStIA7g+qRwL
WFE1RGEtmzdWsx5y0uff2pM+tk7qAY+BiNhqyjd8mYajExD20zWzuDRGhusliyju
ViGC8i0VLvUSTbegTlEs7nyp7PvkCV6jw6pXnrrQ+8bHH/uQ6IukTmgKuIwSRVza
8rBL9q2/NldadEHpEhE/61GoAbK4psI3Zcb5FljXYOkxz7g9aoMm8/+yrqxlEt7h
DIkVnf57+uGGEbL/Sslv3Dz0zY82WeBrzDJ6WWKWnTwnhd1evmIjENjDWwMd4yDM
HMC1YoscCtDk/8imavaLWmSrALcDdPqMbtdNBTNQKlBuHfwPJ6sQHJc51yMT4tX1
FgAg4poyOY8dp5Iu2Se5BO3qVgm1kZSIg73i+cH5xZNF/3z5YMIANt7iVBkD/iyd
LZFgt29Hyr9XYPXUiu/hbetEJViCGqKCO0SD2TYbnOh96wcZWg7n49lPZyXRswLm
RFVL9rCg18IceSXexsAThCh38IUq6yHUYKZvdchK2CY9jMYF9V8yF2Sps34x/tqH
gaQw1WvIJ7ilL02ydvpdRcVM6zlcXSttMp6/jONxQDi1KhJ/g8bwUr0sp65XfdSW
+SYAtn6QNEjILnYXHh/2/uvQSAc0gZLi3R6+X+jAoQ7koInYAPRGxBQoqQnliErc
+9tdidAQ9UwBio3QC+ms/yh/une8ikpIfFAhL9m/riAotpz/V0bLIU6WA690qQ/O
NkthMcChv8puCgGlGqrdNrmJPAH/6Cm2SepWSn7oeWG/sjXDWivjHdRBtjH9Mz/w
L6IxBGn81cPGOZzHlzQ2yc3pzSObWECCCRDLwcQ6suP68QjtA8UNw4xEF010owdv
TtS5IigpxGG8TuDiW47kxMySbOOQtniPRqhRcbR70WOc+WZwH2ui6DO3Lm+KGrrT
Db7vfli4E+QULcxb+LCNDer1GEPGmJsrw6L5U6kOWpZ37TgF747i/rXDRpaO2mLZ
CVhPIhEUDJjJoJ97N1mcMrEdx+mhBuJ3lhOVOS/SwjY4GqiMdkQCCZ79efWINP7r
k+yR2eHsn4iH90dSaKHu08b6OUMjaQYcAwPOsIFm5D6CuyF2TdyZbkQXMQkju6Y2
bjwq+7JZ74Z9wVU8Eo1vWd1+XUVvMbzab5sRq4XuuD2wdh+DrSnJ+J+z0YC8jCy8
WhydZ/M5LvKxpxZa2+oVeN/i02+3UZJxO8UOlyMqQaJs0kT00MvStHoNYpWGO08a
ei2jpt43xBELHeNKk+LSThz2LIuiTGGyDnWHZytHijgp6C4hr42ox88kfpkN9SsT
P0sFG1I+JO5Cn+I8CfaEN6QA5CKLpeYiyUH4NskU2XkZU9IRBA7wckMtSWFAXbTD
D0W7asS6xmPaZZBNx4s2e8z6Ldgky4qJDqb0SefpT9ufJLiIzWKps9XJIXoqa2N1
Uljuz6fj/aLjHc5jnilXVMTGuoiouoIIJzqVtE5wrhI2qIV/xZ7rRoUVUnmeWMOB
QQA8+IljuwDk+lhMKFLV1E7ppwfS4xmfew8XuyPx/Z13MrsVpov9GqZKgoMEjdBF
gg3SYLUaUXshLGe4Z0D3kHh9VEi58lxlye3v4rjIcs3AGjH3b4d7yrRzMvZqMFgG
yz5BOoaNtcCPOPoy2rj50df6ACBSOsYKwzpY0LAt8xPb3OaQ9uKcsniQ2AFQdRNv
Sphmf8b4vlCSurMf50g/Jaj667eO3WUD6bFf2pYOnD870SkFi1ahhdeKMQ1/j4fi
ICaRAQXCZK27lynN8f1Fm834ofw8amC5YB59vk8WQ68vStBDiwTv0ghkoV+5sFW9
+HKsQr330D3S04fbFgLAm15ZI0HZlfIgTyN+3j2ce48q9LXLTU5gblIw4Wh47vAG
1my5CKmJA/S2LHsxTmOezdm3QQTqbCRYw5ge6AjtYCARYy0lerTrpi8F4pzrUD5i
HHhOVN8UXQhaVOga0VRQf7VvfTbzJECV/nqn37JFOnUNhSQBTlvsByXVehwr6g79
enwYoi16fW2hzARzT+lnMq4JEDGrQXTqNHlzBphUyY0/uAK50Vxa5woFf/e6vLks
/Q8W1hP0Xehp6z+ERHwh4KYqHR/8IchzHjntF4EPlo2XwGIEHnQLCZLuGUwu/kCc
ysoctX5wbRZhRos90MOGra8Ds/LldTJ5WC0Q1KAx+bz9Bx0wRfZ5ZKa63aHPxOXi
qav5TI5Bzn0lJgm2MhxEvPrivWrGxC+/BFS21jDBhb4T1uM76f56qSMJQ9JeWulv
Z1y+f4G3/8xecNM0bx30VfThUc/+fwXH+2TesRHZ9z7QaVdtUTaOTsfQb5atr3Cw
w7zhdx8PoN6ZAtPrxhNRU9QjYt/YLvDr9cbJtY5vkM9JZaCZyF/UjhoMHJcw87Mk
VtVTgzkUTFrM7z/a7FSt7kZKiB4IbgcWq+p46uY04MM3ggwAdeYozwmDi201b9ct
HcMN0nG3i3kHk4RcOj3Whvpnp6Vqfr4rLMWCd+aNc0pDGyWb2mwVaMk/Mc/4eiAc
YSte1rkIZ46Zs6RuiH6QZlBP91jbwV7MWc+X+et2tyfQsb3Z4lHZHF2mFeGBkWgJ
LfTO9oOr1gjWbAssp9TzT2MbWAEfGFPlWWFlGyC2xTnGy9Z1j+d2iJ6InkPdQDhR
cOj4VjwdUbWaS5iVIvV+LP8SL56Tb2s9dNfvjMuqA4Z10VMvZ/MMYutHfYM9seRA
XavKxNY6/nMST71boV/nCriu6Oyyt1n/c08n3szghFaLJJGptvgdoeFxnoP4VDVG
mGF523t4ZvEMrKRUOamB3bx0VY4io08d8er58HPE+4ld+a+K6RqYBOQfEWbcPWe9
RJ9u7buWdloCjN/wwJlG79ivRMKG9cEfSjj4sbIQ4fhffQ5+szJAJah+iqphzSI+
FHyZpmI/XZpaeq5t4zP4DyyZKy96ZPFa9uaaDW39Z4LlAPyIS0btS79ZHGmUALUH
lO4Ze/Ye7iGQu6z+RBt0VSoeJBQHxuNs/J/wlsJbpoU049z1axpgk3Ggtqy4VEz7
bR2dRrZtmxhmBn9Pv09qRoF2nJKeuq/ZYHmkNyeiu89atiTjWwF24cHktESvPhNX
qgCAAQVZaoHV6c6ClEYR2PG2XxA3SfZNfDRKGHzYS4r2/21UPcYl140NlFBymF7x
X64HxugoUigYs7N7hkjP9ltyOIkk6lnIK/35Rpybf8yp1E8YPiA3mLFGJyRI5Ow9
GqBdjm26iwbxHzXBLNcbm8RfIxEiAuYv8K04t4aWix9NUso6DiD7TQpGkrAsO12y
l8pcNPZ4CQVGcOILaYj+Y++iN8qUll17u4inaLJmsCU2qxd2LdxrUElkh6C5/gB0
96pWJc0ftoV/T+GU/ISKPVJn8hzuzROHvaqLqU/sHXmwX1X7c/HPkErEv7y0vrxd
guEFkwGbL+M5e+uynDQwFyv/hs2V5Y/D2zcjDfcj1YKI3dgCn3+BtvQbLaCPx3ib
3UzuEo8erFhWaW2fQJGTOD9qOGjvXR3sctcx3QwYQ4gHb7t8TdKzWpnE2GkW7UEy
RE/plWulXVo9ZuT+uFKGw8IONxRcPwLHorYHwvt5zj8yNjcYnxrmkoeTUdKJ1Z0d
A9Dhl6qDO26C8eEuw/1+DyFIkjUOyMXXKNamBqdBw/wOZURLKDUlxMQgfN5m8xj5
2J9NJulAYOnK+5iAd0gTgnyeDg8mYg/XjXfLYPA/0II6zKlYDBIc3LizMmTEjxjX
K+T+3IS1bkLiaIic1VhlofrCOoMi2uzQ2X51vIuw5M/jHNaPAGdBb30L7j8lj0G/
fV6QbSTrWI0bnQfzRXE226LcRks+eecCRleynZTt7Id1JgPpKuzHbr8kjdLOKGml
Ss3qRAJO76jwikJDV2rYYvEjqXvnUy70vEAuBcuW273VDhxFY/N0Sn3E7Q0CwhVS
DGOaTlLgPISKg0jtdYf4kEw0+GPLScmx9zXe1t9hf9hLAZSw9sIz1BAXAzOF3wpc
m3ZZEPPxWDi+K0B2/O5bsRQjjWm9DMez1g6Q1aw2d1QBZ5bk9s5nmfmHWyLU8mQg
GFCdXgM74n5EMpdS+juzoST9OD13lykpGfPIyk+fRXlr8RWYBgL9LYQK4JgvrDfA
tcEPzvgJp2RTF71QOC2j2tUXwafkI44nlOlYW2HFQwufOxLZvkT9Wl/i1TF7U7wU
fLDKzHaAQ9rSNeDcLrFC0iHJn35NkVpPiuS8zQ3eGR4PQrfIVcVaWQALW8KnAcSl
BDMBEaAGirqn0ze7KETulxL6AQhgpsig3cP0VQNWuicXyEvnkY0D+VhwkWBxpwSi
yu05fgQfx6BUjDQeyCsAy4FbfpPUj2QVR0yB0ToIj/c++384WwVoXLvbpfVmCGEn
cqCcFid9WR4Cvs43BwRPstu6t/41M9JlY+6njdSUIJsGwE4SWKMTxA9LbkVSpqJ5
Aup0kjsgLzhnKu15x/2m+3RaIlwOlMqq2gWxXzMk3PwWIyj+izwy52hwhBP5GUZU
uTx0u8RA8cXdmFExCibwo5Q1BUvI19QUraOBpXmIMnNjNnPQINOfyq0V4onYkuEQ
0XzOS8Sma4dCOAuwQ5giebDtBd6CrLVu345fG2CbDcx9bNSMEiVQtRAZXVoncPKr
5wQgmHGcUrXXvX03hrRM9TTYkteKpX5Ii02YbTwm66Gno2eLgI/15lzmT2On0Zub
aSm7q+vWLWFynkAx+c7SHmOuhIh3t+5Sqi3iEbqJ+SGvkbdWAlr+xjwCRZwtoFtj
QMgxySPPHSAGcJJRku/gR/G+4b0AdRgH+bZ9oNQ5vojwEU7gV/iO8KcI50d6aQDp
tu4ZSwMHtJtD9tUE0x7r5SPWR5wZGDQJnsu+CSzTASSvjcXXjZK3zqPRiL0mDyRW
ONDjCs7NlO80vsBoFv6I+RB8xPuzsSdS0oIS7xhT2M/ZX07zHWwNEgrFPOquoLHs
XZWafZmuDl8dJtiCMIZgMO72IjFhcFHbrEmsRpysw+ubDJfzfx2uVM/g1c8uTQyd
EmUlom/lNT3s2xnLlGoMNq5kNxBWQOC+vp38EnRQblgu/ifT/kFZf7PQwNt8H8qy
B54p9PnAjPIuzYP0YFlO3UGaDlShdFdho6+Y0LzVi8+ttXneZFmm2lISJqSl2WAu
9TtE8uMU/NQOgqFxnDaw56EPx6wR1pyGyL4Y5J9CGjy1znjELtXwqi9Ic2qYw5WM
0UJiYUdhpdcy6/bRnHTdvPrepD/CKm7TgJ2RCWfw7ZHqrEkn+PMxQ3Dw3wxb4CoQ
k+Ci9XwXfW8c95AmG9eOUHFJ6+sYdett/7midLAPqd1VrgwYjmJ3PzYTTBNvwbBG
juX1RqOCKZV/4+6FGy5hfMnXIT7XQUElqA3RF+AeUla/k8o0BQ+sOHZRbZIzvCCj
myltoy/RREzCuc7wPkALEiKGkxwYhB59QSUDJMpUGhInz1gHCf/GA3CHjW7MwchP
Zm1Ho0BzXi6j5JhkYD1f1O0XsA9LTdiWAhYnxPvRjArYjgu0FCicgJ8JMTolmWY2
SA/ZAYKumzFlgYF3aXNWoFmIVDcXEzN7pMEmD9tgEGMO+e612BM0GFqL4t3wNwvW
qVOgaiOWJSVebySQ/N8azsBMwBc19bxOgcJHKcvNmuISSoVrr/TkahFgz2YcoUwD
HHuEA789VrhX3C5wrIOkeESdBbSZg7lTGSF19ok3zAXi74rvJ1QlXVTS4JCCk8SN
Y35CjTmHhtvF/qRh8kPbuxEni6xSs6/X/ibqanxlb6wECEiFM6NCicJdE02H9H63
TesQYZOrtPSALIpdRIpHQ4VqEJKYslrC9hO33E1WUowr5Erv79qgoppH5YtvIhJV
7iuFiJHZ7pGNpNYXxk4i9dzev4LuW3830MZTbzQrZRgjbuwhpydV5OX5JzF8pssF
gIZ0cOl2wKmLM1h01HZesH49zaGGP6/HLek7ZIigpsjbabxI9i5nnhnHvUYOJAcU
4T8WjaNhrxRX0Hkg2BF69QsA1XakPkRo0LN07fPNQJam1vbntaFM8zn78G7CkeKM
/oBvpQEBY+PXdj3+iZai+hXq1vKVQcwmKYrTkOrcl4za+oV5nhkvcA3wxL9LCbY0
qp68gWNjLMqTSy2xD9Tifrz5NtU6i3MfSsnXfwUhkWg7/D77oCj0CjZYAzuYjkpR
u4BRhveiYMOgF+b+7ieyrUeMdAaPWPGRFsYh8zPGvg3InBbEs7atsqK0WNHbMqTR
67zuIwjWRKsObyNokyGxwO/Bw554PZO8DRbB1YFsW143XTF0QFyobEKQlCME6gfd
hC/OglMswRehIqaNpoI/s2drQ9HLAn7WQawwcRry6Zi5pBs3vel3Y0qvjsDFOfbR
1LCfzhk4DClEUqGpOzTEmpd8kB6lP0mM3M4GKhiKaeblPsXB3noiOyaj0P08Gslx
KsEuqcOpqhH5zgp9OLBt7TzNrbOx6siYy9Y02BjGo96Ysb3ClSMctsePyJfQPO1b
SWCcs0Pc4yBxkFf/2qS6+N5+JU4YOhR2pepD94rsvsBz0Q8UTeGeidSU0wUfoVuv
RjaQ3+CxoVEoOVL6SconLI8/ikuMvKreCqr7j7g6SLyKGH2uBP1bWgYlvl/UeMu7
AT5S6cy3rIYs/icX/xHIoeQN27ep1n/zPOJGXE++Jkq6+6RYNUgHI9eLzo4f0FYw
ZBNSZhCvjkOdU4qKgjoMQ70uFSArdbUwK5v3zDKt6t+KBRvuBE2zDskkTZucyW1j
+suIYkfnGo9gXk7ND4ry7gJrIgJy/Otp+NMt+9B77bnJsvwBWgAP0dCtz9QEBe3J
cK/22XLlrwEs7sp2/53w+vKxfhfjz9DHPLpRzQgS5uLvJBCDWYFcAf6kq3CiV5uT
qCr7eIl8Fv0rniTTXxkFo3muX5/lBfb7dJlUm4G7dNeWW+tWDMmQ8uO0BAU7gZsk
348jYeDX71Kef1TwlS+5LPZ/w3y//M8gixWJC/mp8FJif4SwTub1eW4aO1y3qVWr
DoBHvAoBV22W5JPe5Y/5OHObHv/GVERKNELqiaED6hHf62ndqB79qKWz09y55GlC
w/fe7bNCtmAbNGdK7gjfLj9VBucEbBfosKCvoTztYH4Hka+TmOq1H2+LCmcwS52U
A9sX8sZIeZJckttbw+TG4VlvRi9pc/b245FyOmw+CiXK6syPrROXUgHL3tkypyJX
1bwQOYVUiedq2OWXcIu7g0dIHJYKa+N6Px2qGZwQYKQLhJ1IPYPBbesfscuowTsT
17muY+SBOPYVEQz2PNixKYqJdbpYT4xUgHKuUwsnqTeUiSop0CGdiqbolgVBavwG
2waA1efP9m25zvHPzb51PQ75Tp9rQlYaNf153a/iyKMqwoQYw3YwudyovMsJRZwv
qxDbY7v+CFQF9doCmuER8cZT6stcgD+lApVZ9dYY639Rr0CSrPThgSg4rOTMafke
Q/Pw8YgnWQG1mS+qmBu2Ags3t+4Hgwz+66sKHL64WDxsGfbHnX8ixHQiSBn/qldr
qJNvxJSH2u8dz7lT1DHGOnSjp/tQzTJHRali+a/j7aCmkRC8dsqgw0JOZd4WdKJX
OR0WerNzpjBZhAX0tVo0cqOQjfSGwhcn5panvYcBPLce41z8kmVaq4UpJKfPeziU
DuwzdnHgYQBpWeLhFmDMFzEaDUkS6tDkakmCkBHzVejQJAkx6l8EueF8BXDQVOUe
klWvoe8pqaPoBZ0TIjILvNKpOGNXWBnRv2SObBa4IQv2dZgBXAvVQmLLR6P8FItN
WJnfaFMegm0w5hZ+zUqulp/9hVq265wUEIqn6OucODDx9kGJSRorCjkboxRFPtwD
wRZgORYp/yKTXv3HMqpuGhOSCisuBnPL5UULXESYaRPGpE/KQXwAcok1eYaSI9sU
StfSgdIrDiYtPYQe2gIHDwTidDqiTISLvTzwss1M48tVusnNGyMTXVi4mh5zuSYI
C/ZfIizzKQIJ4pGzjtWr/X38ox7LqMMoJPxryGpV2JYFSfRTXlBE9yP1kBKnQa5M
79fRlC3DXf/zjKKaTMwZ44M0qtz+H4n/jsP80VtlpEtRCfxmtIDqbekBfnOw1INs
0iOIPaGOFfNGn+gMdjqTrpY6/alx1esd4XDa+Hxpn/Ta1w0OWcKKn118MlPk8wzh
xs7Fi5nOYZPF15TZJb/eSVuKsctAO7Cs9iDJQka9A3av+GPUuTyboovJAhkjg3/t
8mi5dBJkKxnnUc3hMNETQvPh1lLn1MMZHt9sAkDvNBSkb7eTVi6Fln9Feib7PbQE
sNi5tCqY/frT8qzp7TvUGa/yQGhbN1AJhSVTwhXUHbm1bi+QlvMdr3GcpICiFlzo
d1/Es78CY2EwgVyonPUyxuk1BpzTJVK7G8tCT6QOhaiCjHD7X1j0uKbEQ8M6zliP
P3BPyyTj8+2FiN4/UwSARCXYOVBu+mCTHLnQb4D6n9uRCgSF82b2UEkx5bY1U+oq
5/gpW47ALAEwsSpwbtySD92L3g9VNJU42iNHrsAjEodQmme3+10+jhiiZMRxFEG/
od7KlsYEXil/QwxEVQ1/b11spqEu4zqpBV9LRHBC5hAP5FtihKPCdQ6KzJKma3WZ
hRQ7/wfXOMzKo3sNeqtHmpsS5cDkvNoagWpozQPxkypf2aaDtNa6+7uecH6c+KHa
0YFgBo55JDAD/NbtI/CZLnglW3jjE/sXwjrURUvcldk6n9QvRiihLXnCpTqU1mPr
yIoafaBD4z+rMBH4EKuji8Y01EMJxNuYfbgzt/yevx1XzDQU4qKEcIW+6lgcgFG/
d2RTldzG4BND0tJKwcVc2+Fbvz1dzOB1/sobLxD2wZtivIhSBL4gN2CmiuWszWp6
wj1Ktfk909D3YQgyKho1Jn+WAMNURaPA8lqIc49QscuiELrtlPULGFCe2X6TdYpy
G4c3bCr38Ry1bA279+u0EevX7RtG9fg7UTujG6lKB3sXNbrHBg9nH4xlUOLtwtpj
8kaq6G8lFDZOEIPg7LnqVuqPng/HmSRMU03MozWfFF4VmHf7xKt89dcs3AypMb1Y
h5jffqf6e+Zf9wkR1N8AVTtV8SQ51SQk/jVk4ylMPmoKUNDu4+hk402s7ikaDbKd
lGwBP53TqhXbg0yxb0v5mrjAwec2QnAQcGsnN6Z4n0R01otp5hDYpsaEqoB2YPBF
mkl5sxM5yK0TePoh8awQ5f6FnjzpxuIX1jIeG5EmDkZ4kA6Wj70E0X2D6CzAUmA1
G61qMkgAaWaMl6DVwUEwB4+81y5RpmhL3OS4dUqruV+mr+g3/oh0/5cuv4NzfD57
m69M+U2NTQ1nTi21WDUp6/BmK13vfTlCV/slN8VkamaVgp1T4uVRJkENbcpr27tC
5PaSN4EhGTxXL291biorptsxUaRaZ5M6JrQqJJ9vLa1n+06kz4Bzq+5RiPXaeETL
NRnY9cOSXrqXYOUCF4+d5YOOUTJ66szamnlfOnF7ZoUN7cOAjKec5fv5x4JbG4BB
ZaYglGhSMjvQWzuT4bnXiQv2OgTbXv9fm2dtrWKbIZ5k7CgBQ3Xr8PXwqWtNcJVY
Ey/ochybyjqrZJeVdzQxuw66giKlIXvT00P/M5faO2Gnbk37LQ7aLToEnH7X4pnM
COQrdaYMiEc1DDLLqg/ar9y7cLmz8Czl9omtNUymaZkx9v1jiqdltvnAIA5wcmgS
1D2Ni8gMoc+onFR8ldyKkn0bG8VODkDi6pVLTon/F3UDpAHw9k2ySh5Nwpj4qApv
39Smcpc/SCsdbdk+srKkOmp3c1e1VgEJlaZ6tv8WtMqpz+3gccWMLw38pwIwUUNS
H4w6UpBkCfyZ3AwBI/zcw2teLlvJVcKp3f6PuCm/8W+v580SGoor+5MibQUn+Tfp
qCOwAR/Gv5YqEBkiarkLSvNAYSIOv4AerP7b4kKvJqX8edQv23AS5cZDMKOqyw6r
/cYF2hYPtce2etQ03K+ktfJ8O46SWVNQoZOkdLkaFdiDomyp3mEZJfb0ZNWqxO7F
WcH1of7KzOzYmoXSqZ89HqBVu6yLWLNCjoIl3h3qnPe9gzYZYJ49THDFf5Y0jRHd
Mdoc1HNnCotX1IIFajygoyNxsFmijirGwVQy7ZaaWeiczwWrOmzCwrIfQ9LUxrLw
cI60oCgBJqC2hS9Xdni/2tzzCWQianqhywW2ytIvPAdH1acQz8HToCY8Q+oso5wi
HV8bfdziqxnGtsOn2danUwlqTynEVQ3oQhfP+PHHoTfR0Id+WCqBuNiFpzhAfJhD
FmI5vDnKNHAQE2zajyTj0LFVKfc6WkwvX0lv4q6+YsLUCr3lqS+UX7i1d0QC4mXF
bTYGncj5oDMwnqd3QskjPm+6PmHnG9kpYLa6vCi5Gn21P05yr8D8CTbSo67qFijn
M5PajliSIAMgWpAWODvO8St8rKrjTIknh0mcXRGolLEdYofMj2vSu8zoRU7XFc6c
y9F27Q05GcLLWMfo/Z0UGNbt64IMwaHJnownm32XUSY1SQ5W6f0t+ZD82eVxSYG4
spFbYUhMMqSiLMogIJfPSHSAG06hUaxJPQFXJumcK+GYGpF1YOwd9dHd+R1TcZMW
nhLF+ydOHQNN3DXmFDCJEivE5OSu6O3Zlatw3A25zscHWQA276fVcIfEwtDyIRii
ww7RujBjSJv0vU5Wn2SNEDtQlR27Dmp+jAuhMjlrczfrUwkLHH3DrSftaaS2FkNh
SbUrU/ZSEHtM0sBS4jvz8zhCYJGJFSBh31ulAsPey0PITTLFi3Mbgi26hUWgkG2r
Rtkyn7AGDbqauNTMXWDxoqmKhZJ8tWmAYR+fqhpwfvM5Pi38MKxPWeKOOayZ0WBD
6l8jvVPvAxD8fAUamMFM9YgQozxP1Y315MPi5MIZXaXgTpvwSlHapuvoiLzdWO5S
YiYDmpfBSLOR8EM7/5sivJn1z3ZBhcJ5GfQshoS4ge3vxTH8bC46ogYFDDa7tSU2
A8Itxp6oWFPziC4vTT7R+0secifImjb7TmY7SN0Jrm9MnrQvo79uNHDDe/HJSDfQ
epE6z4PVfi8Z15zIxdIVZi4zitMEEZSSGXWMNWdKJogQwZFpMSUddTHOvqO9OMcn
JhlPFwGVaJaAFBt2satz/xH3uDxoh6XsFUusgWzR5Q0zZ2XA5QqIEoTEtkY59s3e
Yf0pNDKjY4mRS9Eh/e6uaStMXt3+VwbiM+5gRMKUESm9PblBbR/qtARJcGaonhR0
EUuLQOz9Y7AlpjnMTDptI8pqQ6O3yttZK6K5AMsRyseyCoxgTL4EfWnnsMHXwyFS
GCmqtWhfMNSzGKoAlqfIihnwCXsnmSwpkM1a+z4Yr/2sY9eomM7rHVEp4jh9vCLh
FL+lFai3sISvoSh5zpcp+nwL1pfG7k0sbOMFHDqQDbaRaxFslHfKQF+yDNskvS6c
WdoevGshNNbRZrIAclJXGMXAD0Fq3BQLpPupS7SHcEuYLMNeLERrKU00QbPb0TLK
OuJdN4vn2CPYWIicYNFThvm6mmEZYjXUPbpupioGEHOmDj22+SUeHXSCK9fjiZU0
KAu2pb9CpWqoVVvKhTjHP7rGhsHNvdaXVnQ86j4UwYRSKT1p0tmUtifg2Rg1LdTD
+B0f15QOrj6UOuPcucLzZndMLtoz0Q8YXOTcetVg6Ml1VoJ1kIJ8eLzsrR9loUYI
NB1QlDWoB+NxhI0+J/zwXSbU0fwcKq7rTrFhqmR15RMc0m2wm1IMtw5GYGqNCpnl
Ujce/grhwcQQujT5gEPB1u05N9+6QzQ/jc9Zo0ev8IRqpdLEWuHUIeauGK6KYqP8
j5Cvza9Rq2KteiQQ46G3oEO4CWXv2S1tbMxjfExuoTaes0nFwmC5mpE/fWWh2cHx
pRCB/YB/08qwbBhBJW9zWLp0Rid3pI2Q7lmtKkfo5pDjRPiPi5FT83o9GCb8cM/m
FTnY2EVZi5shVhgZS3USkC9pJzzbycsjfmiDfpWp+dob5/vYDZzbCmGtm4VN5e27
E0S8/PFPiWhVmMcyAZ9t92BOyfeWvPOaa0rKjT1f+TfHg128kMRxvEf9mCq+k426
fPSX5/fnHZFy5+cxZW4r5Z86qAO30Q4cZvrJ9UpR63fB62lW1Bi4jgtH/k/dytE8
KdUnf6XzCqyJXsm0HHO5Abkpz4U68rMVcNFU9OylDtU6Yl1nLAcRlnM+xHZ3IQAd
jiigEU0uZ6RH0SYaOMDd8O9yeNWAfXOJGBdaE96lAFTmf/4zJCBj1SJOdqtjhv/h
Csi9pUSycidFeWT7ZaJW4BNn8oT+PMzPtGDJURo5gaJMFJjh7xAWF4MPXfqFyDcH
q8KcONBc6L+IOfX5VLv2BTadbmzAEVnFTmm1rYeYMcCqIhKQaymg8nkPGn5/iJzJ
kVJdEKTgt6QK1GelqAUpbikPbW5LBLMzpu2DYO5bSot3YWvwGpPBI4IymeSETQE6
6xEFbADOgTjz21U7Ec06yFYUCCUmj4fF0j71D6SHTQ9jAljpKpMAVieg8fbwpR/N
VERFV++sQXdEJPAOxAT/vfUvYJqfJujW/1DJsoBEYEVF/Z4imkEZZ6u6WT+cx6IO
e3kPlW8rz1zi1o/1ZGmi1c0gvwePQt11VsTgf8GnUt3YuQlitaXNFIhqdzEqGhSu
XFnFRfJMSsrUW9dzAd3CWv9BJ5REu7/YorZnRM3S+M7Bej/3vFw19NaKP/IKX4EV
cKo3Jjr5j4eEbKJxPWlhIBtvIAMrz37W8+GxFAK19sn5loAlQLNSkOk05cGlsVSf
wl8IWbcaBQS7NnlaAfdB1sEWGqFH0O9XC6QUOrArutwKRAU1IwAUVQsGj+MVQIAJ
b10eyJrgVctogwj1bbfAixKFxJ5xrqJ0PE6EcbrsUJ+5adIQlc77fenduiRaii/r
ZodJrrLBxlU5Aq0NLP5rWaJcD62cTLTffAFTv0RL4GLeAxGf78LBHnydesSHrsQB
Hpoq8J7PT4rMuuOA9GmMcVjP5cPIMlwCYtLdm1a8mfeC0q3m4iuGSgEyAvRvFDQn
JujM5N1c/zoIJ+VNJVnmsc/GUiiWnwOB/twRI3jQN07MOuZPp9+bGalOe1+T5/+a
mwEfPxhuCbOG/M5K7G1Gr9h0Wk+U6rheRCocwbuNYoeTvSiaB+VDx8I2Ij1xxZNt
QlE6OTs+kGJZxoeZEAv2Gvkb0IO9eeMsCXx3yeI74OZFY6TcbjU58dLJOF9pvwp+
pS/G6ZUp7xy+jcVRKOxa9kWXuEoqfbJNuriI6YGK5/JK3G2Fpkp7yqNiDVvzB+qs
VMVlNL8zwvhPHszgdVEk0G5NBmTf8R/xbxQqW5xmdR1FNyKBgcU2nUJ3cV4yZmhe
stbR/hgbSg2/BOKe5bqxyGmoWC8Ais2oIZK0i4zKTFwlP3S4hb64NBDtbVmke+J3
QINJIuP1YtdlbwlqZnwlA/3O5kSVaS8atUtYwLkqQakH9xYIdjeKkTUvMpOkMsk7
y6KnmdRBWbchSpxtCHBvLYcNqoSIJHBkIL/5ndV39/4kNCtbKAjwEr1VUI5wAoLC
GVyMQNeYJrt7i3/DLYDY0d5iaC42jqjBPD/jkd4UNz69+b+lQ/MPxsGDQkuPy6dG
Ej/eBjU866NiCmPzQNk6IzatZQRlw8RJUeM2IZ0V141BvGYcH7t0OZZW+1gjYyDv
1s5mg2KOD1sGzeLqSMmFz2HVAQI/ejvFTx1anAymMJgzzOjsJduJHhQ1VEHhQb34
DqkwClg0e+kTQHRMVDr0eG+cyHYyowclaV+xOGr6CPgV+z6VK4L+Px0YXwv45au3
xBBeThEoR6ZVBGL1hLYLSyYLlTXzHqW/s798ehZbL529EaEP2ABJZe07wQTgtz/N
Ugv1cbb1ZrFyz1uhiI2sQrZ5bckqFafQw7US2NYaRqgNtcGwjBXE1Fx2wk+xZnhO
PKEQV+KH+ZuD+UDgKAXB6paYmG+A/eXM2PYb0dScfvjBenZjmI8W8Ca0yPRHkfe3
OEzSPWnv0S6ZBwBxCgnNx1AdiEwikWwFhYN7ozgqTM6ksXpiu4AQR/fPijq+/fBI
n5b0XCEWRycW1LN/ZkGEA2paFhS2uXRMAUPz7D+NtVxm2m81tbdUHq/Joh1MPufD
1kG7eITRH+FnIS4oFbldhJ0uzz5QlVbr3YDnbiGx5K6Ddbi0+xvPYburxBon+Gzz
Lhdxhcy8NQX8KlSCR2oZn1XxO0w5KCrZ/ma1LliQw1Oz/RB8BMmPque3dtKT7y4O
DYLaIubpDVcGqdPaaHl7ZBzSBHKSVGdatLBxo7nXosS3CoI98fq8nX88UX8Gt1Qq
+sKAsYfF5XMrrXczzQ9WhbK68rh/VoJu671d/PiixX+NRZzvo61gf7b+g8sBAdP5
EuJrG0hyfy/6MZmQ4Fl4I2/Nz6fNzUn7gHhMx67OVOAxQhyp5wRojs2P8ligvXLf
O2qjVkh+SeUhNkx31EbaueGe490E9iOZcMGJZR/bGgwdNInif5bZKfp97BbNasWk
3enKOufSJcJh0VtIkJu4Ger3NycN2fKhALy4fH3TMy4YrwKxjDFM20ZH7QzHf8ao
a6+aiBj6gP8ZG8/o/1HA54QXVvY/128iufLeJHj2/hCMzQQMShp51Uq/1VBln2Uc
2MRrcoRaYs/dJPHpzQbnB8jp4jjM2vMJapx71RI1AsH8XviFIsyjj7i8RLjppJ00
/gi7wsKnYxT7pR0k6E6ZHQYDsejsCusFSGUyOo+5J1pQn1Q8gs5bBrWHpFZnk1HZ
1datGDUGiuLi0GtGJoeY7/POWFvGzEtLCPLDHZUoiC6GC4sxan+MhmHfwLYLO6ta
YDWL+IWTgTJ8JwpW1DsQ8PUaxfFp0duSMInpQhgGh4RHKJ4/aAET3v4RbOTvpE+l
GFTJXpri8SwNXU+QUGwI5eUCiTSk77W6vxVhWaO2c33sNo84JHXQuL+hwO4PnfsZ
4H+s/AG6VvuSeRMqM0cfNqybbe1ZngT0ZIn5TDHFOAiKFBJ4YGMfzy9kL9nWEmt7
HIaqCHXwsEZwBl+mhhEEDPJzeR7MgaxIlMAz7elKfyKloLdjJ0aQyW1MSZ6Myrpf
rqYoQRadR+03JWBLlTPN6TK6gmpWknmyxkUOsVKaphdkgZzgdAq2tYTgN3OsCL9x
BDTFYmbMme1rwP3x3kwStA47qrLiOcvEXl2uj0dNX4uwnyejhlmqgu+8QmW2c54d
mNyOPAx/P4JhcUMXTAiuv8iwPgDXZu46reD2lAAfSSqp9mlx24SCtDx6n0hCmi/0
D2iIH8gr/2+oC6QrcRF8EaRSn7aO/dbQyiudYugw3pW6YfJeAd3+dqCUY8WGJvhK
pX7mctT98kcSYKbAW28rW/DFWWc6UgQg53WKbKlREcaGQ/U2jntiuQtC7TYLpRHR
jWQPOUNbAaz6FGKQ3R88WxMirzHZDPCARS/SQPAiVGUp0ZfwKMexNZ1HKO8rw220
+UqG0guji2ARX8cSBK/uTb6vvoYiVf0xxd8Zsb3zoq6FZJb1czJJFugDvauEnAuf
1yn4pgI43fey9dRFQQ21Pr2RuoqamfujmSLyTVJOZpsK9OJPADVDMVE6pK3qsSsW
jC84qNALM0UHhCFZZYjWnrTdn8/AIh1YslFxKy/XxsWzML4qUT7K4b4ZxIzGTSnf
ZNJz44yBgBLjmudc0nWLsFxC/NoUZyC5i/CULZ+IkXc2q6ibWwPQk6LozL6E8/HT
koNPDjzMoElxWagbTFs25BlhEiNvIAdzVaA2SoK+gvIAT2/kjoy00/fHhvowvDqc
bGcTmHTYdi21ub4NnqmdOqg8Cmbr8E6YF1ZSEjvOFFdNAjp+i9/1IT682P8VOYtX
q4wjdMw0c0vakvqCtBPTmdmEpsObutmgIyOk31ghZtH1QtpFFE+N6xDwamdHjOJu
EZfpoqcTfus+6e+P8aZSm0aFX9vFaeERlwGK/jb5po2GoRy2JnjCieOmsJdsqTLn
YWLrXiZc7DlI4d8rKYXeDlPhCkml58FydEG+OSiWL+KRxyb6MzOBGj8X67iNg25T
ZFF3pwAb++oZQxM/9D8duCjZkoBrGRxoLRMfP0OP3rHtdpLxBIjtBwQOy9x7SO1u
TvogEjS2w1fsnGEvzeVv+N/jBPNMKX2vH/skYrqLysJEs37xhy82bqiQp7mR6E3z
QChd2OBuErOF1K9T7bNbuFsy2Fkzv+uWVTQaCJsXsO4D+4I9TZ6xcSdZDPj7iguu
Y7RyYGm9vUDIaw6UnZ2usjKAerGc+6w2Attk/Ky1XdnIJ92FVoqZ5tSER5EcP4S/
JoIiz55b8CtFQxfH1FmHci+QnVFXmao+/AkDaqZvIleFjsz2V2he+tGR9Ejv62fi
aSSHRGt8jjenzD1enLiNrt+4QcT/gM861sGPavZA1ayva3sLrB81+is7EpOy4dSV
kWzwMov411K6iQIzQ4zkHK+E9MeLH5xHTpb/b4U3i6U5T60m+mlHiOIUQOAgH9zg
EIssFcTIB1I7aEqw0A/VwkuruNnaw5E5HV0e7OHRNcGSbLTx9SReAhVn4UIS6ZXY
ewwWha0zeEE3EvP9ub7LRyquyzxxXxmo/3eQ2Lbh+9WkdLHTAq3Tj+MtK/OEw6yo
tGQKY8gLHDACEHEq5UhpXrGUJegeDqxW8vi77NhLt8LfG/uST6hykwmlLXSy+TPL
qYs0mXNR28EH6zmh11wEhoUOiFncnkNrfZyAxm9MV05smMaR8eLdjoRtTiMmpz2j
kkOPkj9AEYJ9R/kTPoEVBVmvt8rvWq6MgWBAP2Jii1FksJjSIcct73jIpAn2lTQe
7raQ3Z/UYngCSrqrqPMdeLLSXBjZdEUCHVruQ05savwsdWcuQwNfrK8HDGORKXTw
5KO2oPOxLfwqrjhPA8+uGwbIgKYgkmXfkwTzzgBCaZEnq38NBIEmZr2uUtV0V6qt
AhAr0JUYHJ8Gjk8KwlTrCMVI/yDAn8vy7sKJYMibcLvc37XuLUiHC9VDLm7YKkGU
Z9bWQ5sKYjqTRAsKhP+Yk+5uaKRJ+5ymCjFdEzWTJE5EjX8U5yfU5H7L/FBzw9km
1Jfgl3Owxz9g0DKzIcbh+m4pbJwipVP+dfXbRKPbLjIDw9w6D+NKPN6Zx3WxmnZK
YOhFKqjJBIs5/DE5pluserhue44cSl4wgbIo7rJaqQd96umlyQ7IMgsIHwFQsNTH
3wiIwIFnMKf2JywYgvUKLZL7u3D/uslUpcJEcLzT3rGzBu1p+9UABEcUEXq/86PW
uc51Kt30cu1ML/MFxBMp+wWr8lLxRsgKj9nsJ0LxfX9pctFuQIFGY8cm6zRY7IC3
bS9G2lbWI7mBjZagA95MAKGoyFJTE5HTTOr4aHAvzrvXhQEA03gkRg79Ue293erB
UH0PChYoaryV2W05wWnEfJuj1jnoYlF/eS60KOCvqOTJtPvF2iKvnKH6+/3kVISI
Q87w8TevUe0/REUpvIzJo5FKUNzDVkmDlJK9UoyvudRPU9UhhvP4J0vNlIWBtjW+
UVn7cHC40DcLat7+FcyqksjpjF/WVez/0h/aERZexd7ihVnSe8EaBODvT0yiTV9g
3SGg9zOHmsnbSBHkk7dnM1wg5CiRwi/AaT3MfgURrGj4msT06OW8XQUItBPgnwWe
Jrs0DwVzzMg6O62uwmglkpHYE3+tVHEXX0m40on7sM7AqdV6VVKhAAMwsjzkFr92
CYYpJSsK+/q67xca9WjYzvuI6Y8NEFgmGcpCyBq/f/ZLNHQJaLVZzpaCskGheMd5
3ai35m5uloGHYpROLduvhD4sz5AZ4lTvP/hMjBjTzC8dY6o38xxXGluS4Cj2SPL1
wpRXG+/VsElWU6z0WOy9MRILF7W0conz6u+INR1PRB6ueebfQe37EhmzPJn+VqF6
ldKS/Y6XLvCEtBBMa0S046ZxIi5xSewA+ktE3/apDqoH/xER2U4L6POzumNytBkf
FI2TDBVt8js5iGfpmxFLN7eDY7f++yFSCwgdscepIFpFdBg5mOQwcSn00p54Qh7P
zdzJmQji73mCF1YZkoxGK/jzEo/kicw8OhVM/GTfo3PKR7gpN5RIAlArnp3V6lEp
n9EUKnY1pj2QW8oM2J9hQLCaKZu15KZTpHTZKV3QE7dnwJcwiFgjvyCZzj/asNq7
a5zTK0IGuMvH6TDGRo0DcLNncO7I1bhHtMrlV+jm+/n9Ho+tAe8iJmtVZiYFOMZE
Mz/uvP1oQb6JKBQ2nBHOtUez/0a/R1FYU4JWBCny4UTXzjLu3rMlo5OTV5c70b2x
aO4N9nNc27U28pxUJ3lqo87LbphPVh0t2Ryb988tkdA2kF8oIHdSJ3AvilCKacSh
ERkxrZhQNT3snE07lY2KxyLJuiZb/UBmNUqXQJ5ZMkkpQ6lJIiGC8vfkJELmk5VL
nSNNPJObmzNTjFeU3jakQB6AEP0//MuOP4JwTbDoUtaNAr4BfU6j+r8Eg7iIa/Yy
7FWSG53tSO+hTcOUA5av6TnL5e6daXrCbxoBkhTZuryPmKew8YTM5wofR4XbFSXw
dDXaz/Os89x5FlIv/i0hU1RKZi1oAb/EGr1pmA+2xWSTc1Jr5K9DnONJpFUYiTB1
yxLD8j1d/zgC8P/spN+GDMqRk+BghzpI7U8k+8H1ftr+dOQ0rAT3+2PsrTb/DD78
a+uUqrU72bM2H0VHa7EzCeDmY/RZHFnXI/it5tFo11D25Aw8TN3BwPZLxYVf72uE
TPz8oHi99IB8NJAAz4ydq5xRg/YOlMhRP79V+nbPpgu6mXqbrdch72on4lz67FEj
ZfUd/89oSF5o9Llt6XCr334XEuRAXJsjtWZfA4wh+hPgLu9+Pq6lv6R6aLBB/Smk
pxBr6FwxPe4xaYZF8bNS3Qz8nPttdV3w8+JWHcUEfPIYoSruwa/+ESAlTUpSLIUo
2mJps/STD65Pji502Mu49KTUEhQQcrngAEvrXETGi+LCzDIQHMQF8wIAJuQVjOZ/
Zx6DT78jHyz31kP0wLkLb9jMoExBPXcHnZ0Tqf3P10JF5IE4Zc5xzk70o6N3BMq3
O0sAAOsisUNR/9lcsyiZS0vDX3ts83ykcO4ags3J+nLYB01dQDRM2uuT4iN/UxlV
IZt2TZy2ac8EHDgD53ZfMceE345mnZC01I5YEJXGjQbIyCA9OsDpuiFFSUvz8zYN
N37bkE5VnZkInR0Bq7czxC2vKNVqbqIr15NCJfMC4z5NE70vqZL9mdRX4OC4ni0t
f4jLcqsYs5f/vuvyAPL+l8dur6NiFvBKBfjiieoufHTNxkssWns8pGAyBiVxxESx
6ypiZBq8SoSdKVjlhTSyJ5PQkrFuMKt64jnJh61lPmP4KKH5CC3R4Mfe6pGMtgUr
87vg9Adit1v3YYAuTfRv26oSvR5HNZkoP41ilW8ZLcQREXYdJt8/5NYtyeXyFaoI
FojineiR8id098ky4FabXSt9PZlQqb56Hmv1O44UBIBWaDkj6kUaJQmUi5/BfEh6
dW34BwQskFF9vN/Ao9WY6xS2Thofl97vNIMllKumPTobZ9h/0PnKfebao8DHaAa6
X9ZamKltTfEsXZ73KJf3m++6l5xNHW04hbaAR2s5T0lTkB6WwHtQmyI7QSusV+kL
+VL88Ph2ocgC2CQdoYOh0y77cUvMdXQTlTIwpeFYnk0SlaImfDeKf2cor6xNyqN8
bnqDyk087gd3bahs0gsGFAcciacMypaGYkzm7zcSW2cy6pcgE5rakRtG7wdvUAQ0
ID2rZjYGKaFt62DOaP+gHF/hNMFFIEAP9/UpOZLuOM2MPhtOBmH64s1xx1SfYaN9
Opl+FabI/OqCuJ08W8WxNsVD7QddPlLNUEBwINT3FjMExf7BnBAlDxM7b3b/abQd
AUbokr9/dwOWDPngO5N/OoKJAJGdN2Lk9pON3YEgs3X3hbY/zaKgopqYixhxfDJd
REg8sf5O3/4l1heeTk0eVmdShF/EEUmwO/koltFnokMckNNKV+wjKuPFnC+tnR4l
mIVx7TVAyFLHyh9N/1dadY17GjPckKnu42ZVFz+806pIOaQjhdgYmMCrpTJk2IeZ
IHTk5oTttBzka8GH/3KkWezE5GEW9/w2NsVCfoiM9QmvGg2uxQU2QQ0OOasXzpeN
WLyunG1axbiv14tRCZK2cr4CM2Ty9kb6kFKip/k1V94WLIsvVRXXXvHusz5mZOjc
G93lnRPe7PnOjxmabnF3s4ObkJWqbIpEhfPyaMVN5e3aMqiZ3ANOe7vZgSkzEMEp
ljXBjvI2ZXaLPfYxtaSEM7fRuCepVE58R0kY43GrAyQnmhOzcsk8PJLnyOwmL06V
Symam6oI9wGi/Jp9nCrD2v7P0/sAR0SzDjzlXzredH0i1sPbAnP/+oDpWUEXiOHH
hf51sM2aXTOYD9eieXHaje+1iHsMG4r8qUHq4inWMM8ae2rt4E+AQ3TAKRDeR0+N
8n19jM8A9fmwH6w28q3b2lXsTYUBEtQ/LrMqsSZeL7XQxOH9UH9X8ooyZYXbeylN
Xe6EKURVfm7W0gIjVD9pbCCET7wpzBSj+qFbqo057IPhgek9ZOsTMYq4uSdYRxT4
dQC1RfaeQxeYKtSWlIm0ZHcE4119wXM/yqFMNpRjMgdDO3WcPMlckJiGMToNa1vx
CKTXUunyZxROlQcXoaNiWJREp7owx12iZTKqmBwmdQA21uhyvB8E93Q/dUrSHA4N
7qKOezF4sbu4Dp3Mz7cUSoU9zMtN9W7ndaGp9kMBzVXOeI9MPwmJo29syDcyNfXM
cZDBZeShoHeTGJAkiHzFOsKYtxV10Dt7ObOnuAl9W9ckLICk3Ei43Igt2F9MsX+k
IE0e4J1CGs90DygZnDx1c+0JJ3QAiF/uGeDU0F7Api2FY7IY8vdv9YDBNby6pqvz
XRwPaBlp9Eg0G8bp+cBokmftBQWI3o6yPu9gIQCEANff7I6Hq1QNlkASKKDuD6Rp
XhCchDNLE74kOEeFB8DdB90oKeIwAi5Vkh/uM5D3Fi6ThkoimuzpKxNDUftl7tEX
6b817lwgX0bFzTd/Tg+4DoznGtXISgsfgLTWOTzz9tek3jHnnZMzDMM6hgNszFG4
wPT7T6I17ZJ3vujdID21ZZJafH0TNYgvYaGDfotuFCrTcngpoZATw/6eOq8Hmvol
6p64cIHdDHNYJN/LrRD76azcYc0H/RxWf7N+mARn1A2NSMHil6WodsHDguTUTOZf
G/BNJZicc07W/GLZfBnekbdcn3wgHSeohKHuLsbVc1rCmjNyqtID3Bg/qkmMcJjP
FsnrTFcBOEochKUiwucTlJH6+ySNytn3N2OJA1/neLAP5/LKw2bOUEQR903sUyu5
c/UYTijdX7UFXBMENMw09NcEGsROv2gLILDb+YflNSjDP49tbKQjqh8uyiIq6Fnw
EMhzJntnWPZtTAZXulik7KkUe9hiNRQklwde7kBC/O51iHsW4jclcn28n4i7qGn3
m/kv758Z81KN0T6PKZUSTF1XfBpghPGffYnFocG/LYwTXgPaXbIAYR2ufpmplOji
FmZ7Q/yFaYwcjYrOIVMnU63/xzvSV5j7weWXooZvNiqBHdCux+UsQiX9UlsARDqY
KfgwQ7INj3t4hEkHB9E7RkP7i52iII2N8SNc6QcMyeg34egFTmJfSj+YM0RZSbMj
3vOu5numarHMJVLuO9RnFfMpyZC/vi34bDBP58CpKTK8XNB2Y22CzOPHGCXvLXWP
5aNnHDJb27GlCGmetCpxyRQwjP5we9zD7MYtQgesgSSmGS8Dth+dMgccef75YTzW
X471mZiS1u711iYsSg0oo7vyhZn4El8VgN8H+BVEVHoCtnQqHGIKmpIWAZlOuTFC
Ufj34eD8O1qepp/Z5uxs6gpBxsAqKnl58R3pOQXpod5Ev5ECDCFsHyKj6GFP++sP
dfkal0MvJ20iduRb2zRYTzRts2e2MBatuMXI5I2Ra/bpg+9G4VnBp81KOcnQsNM2
WKu1nytCHZQSCht+jiTW1jD09QhWFdIvPpXnjuHt+w8PLB84CzOdAkOnveeU6Fnc
CXncUCp0dYj+/9UFJiD2hy/ByA3o9+6qhARo1gf80To42PSJ43PHnNDocYp9yEWA
yUy2j+srQbJ0ARKZw7IymL+fYTw67NCVpgWi7n5eukAt2anAnfTrRg1K1/6nytFv
MBK/X04UVhNf8XdwImM0wQFchafwIXVxqEU4l5d7Ks9BDlThK7X93/k0pKTHhtmW
QdvUJvmLiqvNx0ZHEQZFEBefyWhEFfzhAcbYJaxNwCZJ3Vy5CUxuFN7HxWNjz2UN
2vhdd4IiWo9S2FqU9j+JyMkE/WHqakbthBaRSuNYw7J4D6+r4Nx+qhok8BoL4CK6
NQoYgtLTTPwsVEaPz6ijgdXT9tktx0WdGczfTLeLo4U0AgyCFihx4z5lIhTtVGAr
LHMW8QV6D18KrzwhsQLF1iRSvPbS3aISFp3hfzUFkjkjeRC6D7cS4Vn8u6+fQTND
V7HRvPUSHirJhPtZvtUzqLERzhJ1vBgqDZtErvrAS/WZ8CmRTrlfS7vUxn8X3HQh
vbI2Fzt6Op9fXz3DKCTitccxkJc1acJiigNR7hie3hnJtf4vY5ca5VoTuUPwuwZB
JoT4ZBLeHfoR4p+xiLDQk1XtIiw3IAIRgLTLzpGU9A2+1uFAqfDZASR4OMJ4zgmY
j7qIOVeR0oJR84klQAFoJlRSkiyvcQS0R50P/570e791SwUDof23aWZRqWImDGdV
tdEtMECuA+9qpRTQlxCYDeTDWiTSesUZYgsDziB6kSUZ/puP7is0pYAW0q1DEEEF
Gn3K5UIC6TnRtcJoGY9yjI6+ZN5hm0ct7gM5EHJkxqEIjlsQFoHr/34iiycgukLw
xVc4E6bAz8UHG/ztJqbmZNGNrv9EHRBJ4o9ea1cRo/u8KaHTqucF7FZzqUG/hqpe
T80AUu9uYS7seNURp38fJUEgAljB37cBoRaJ9R6p6LqIDgbbD/E60vcTCRe1Oy3J
MM/2b9yNinHv/gKOImlaMZpXjZl+MtVtlHT1ZH7i3RIYaJ30FpCh6P4gncGGDnap
5QaXQBHnnIXOPT+8ZboIbUZnGmDBz1Z6/MLP+Ap6EDFWat8JWrS+LUGDqPqe++Fj
uLXTtQqtPElkiEYOotkZpAcs41D9n+EvdykO0Yw+tDeZmizxBd4CtppkZU6KMJFM
+BdSsSGvnfkg4w3QBFupG6WEvJm/4PF6sChn8NrlH65yDutXFC8VQ/PDSg5VhwEz
y3h3ZTnagI9YvFurUbqIb9QbeM21I1Gt7uXXcUm3mv05X1t42yIJcwOCGUag8SNE
guQ7QyApg3QT9/FvKnTXgjYG0RI6fhsJ++IrwfX0gzuYpZyJFIjHDbyXYmvbUIWw
ctsO9rvql3bLfrb+p10BSbCdS3sK97/D8Akuzs0nihxxOiCdKSATwCeTwHT2Ewy7
MKks9BxEEupjAvbItzVNiZm6Qo+l5tITwj1W4KqYvUc2ztj2YL76o0ISq+afm2B5
y/ulATi+whBiclD4G1ybJOFLJGvesv/C/naViCc8EZskeyGvic84t81w5rXyQyV5
HCmOA8JuRZpBSMV7Rzcn55HNAzhi0zVK32eCni2CujqAINeVkQ0Lnrgcf1/km9Fl
u4ZExxTBOTUfANdFQacTxjEmk0mBWRi9HzCvbN8Vp7FBDwQ2gB3aoH2DvDNByj+M
/NWB854Osnt7xltnIuEm4slJpBGmbcLr4hMxQ6d1pEATq2JfYJFs9Q0DzoWrF4o1
vAjB6Zy6173030y2ylyK0iVjZvubEmwJQLiNIDKd9yVDmMPqnlZjEo4hs1qbiZib
Rp5AzFZX9MSbHnSXsRgV6sNzV0o+j9BXguc/M0sejyWlOtS7GOWvffqltsBIUNxC
OrE+jRMsBlNtTqK4KZFFkC+kU3HJ+Xeo/j+EBw+InnMlTcbRrfgzwD78uTsEZFFd
vvNkwXDKtygTg2iq9LlxPMkUUOl/8sdzcYHZpBozPXME5U56OsIC4ONwVBk+Kynn
eHcy49iusbBbhSrsKh06p2PfeVLY87rGnV9Sr832N4qDhQYLOVFmNTA1Bz954N3u
gxsTdF7f4DARCViKFN+2z1TaX2cPMpfn9R4D1VgE/mkuibDx/+oRxohHTLaBJOOs
OF+NrhpnTlB+7CjBkNF0LsWoY0MaRlYa53MXAkdSpm8BhOEtYuF7HYCxg9XhaLj2
F7ovsE7zXMPLSBmERrKQ6bE4LQGS7vB8kQfQzhqDHKg89yiN/dmp/Wczzx5uDNjs
i+do5C0MjEscUNxtDViw18YkNzOlK7ov32skTM9ubBpkhbay7CF0sqLM7prFUrlq
at33zNFhmYnovd+T8b0fHQ+VGg8OgmdEnFccAivSxvaa8+3VCZeMZtO7kJP/5VDe
2+3IJwRpYz3kuzYKG/XMAQGp2kMeK32iEsUpBY7QBed8gSacSsIOk0RF1HYE0OFI
MmPcMBL68V4+QTp1oPpcqg4owmHSPps+z9Aewe178vc5t524O8YAtb4QK3l/OnMm
g3djzyfICyGAJyywM+WhoEJdINdIemu1ZlbhUVzihqtg+i0ZZD6dseFeWvAMnCMC
1Fg/lXGm0KKUd0FWylukUAPXH2JKe885uXs0YM8eA9nT1vZC8Kcw7xzFn9UBclxK
lsWs/vlaOZrkkbq2RsToALKLq+sUkT1+YpJamnqh0Avs84CIXbe0NSw5fFPXHJUm
lKDe2k3gMVyD3Cv7HTOUs7ypVAATMIfhFVMwIIDnQ0dVfa7JdLjWShS9sI2853WS
DPgT/J0NSNIYnvyYQ1GcVOWq5ETn04qzFV7tRQI6WFLmynHpNDpv/NSF+twOo6H5
CumPVT/UWQsuSWH3aFZfsOwVXWao+rxZ7LkCatePt9Xt83ey4ltM8kPo9vGENsQX
5sJ97CsTW96GSTzAEtBP/uPcJ/BF4O6xpxvGHKbNwAiH0zHa4e6VhqjNJ4nkx4pL
pDOt7gv+TNagcey/gPMclfHkC1Aueh4TUL2t8of+VsXTcIkD7skoqIO08NWCFMsy
soCU+GXakxDW6O1sYe7LdbX++pe8L9lbV8fWV798p5rCvoIyX+Ict46UeUOe1twH
LeUMM0+socrQWjFb+pIFLinCsnNgljvGaM+DWJwZEpTg9xQmYE7atwvtQ6MDG90R
ZhhbOfmlAfmrjbtZzIzynAVuvi3GL0SLbWPKVHNKEWjBSGiLo98tn33WX+6Vhtet
sAfpClsmnRYSn+ywikTRzrMm8y/2cz0T4i3EiERbtewfmZYIoO7BirJ1219/fDw8
l/DMeBGaZZ0J4Z6eLfqkO+edIyrLVHRW9B3jjxlDygcUAFuqJld6iv4DUq0gRucO
WaloUALP0UablvoSh0v29yyYAzGbVj06epxIXRFqUR7Cq/+Dwgk+o7uc83KZZ8by
KrzfOTa7iqI3pVAErs5gSisedFr4ABFhsqsfZKOHx2xeNtRnjPVgaoYmfNpYK1L/
Va04oNK9lRGUlRG+/JUVqaxAjdro66pjPJFxCFIArQ4jkmErATAjbfsVJJNgHSe+
mUv44ouHoGJcUZJapSsq/1LMJ7usDsTogE9DJg0DDXJ6kLMwp9mk6JMGsJWRGjaW
QWsXJaIg4CKlwsAAnG+b1wdG5xaJ67JIPrNis5AfRSohs+XcH2sMX1A6ZE37TnQM
wfKuCqcIqESRcDdXaMuefNB+oTP0Jq1WUhr7zLdgcQH5DGdTv9iBasC5+GIzr50o
lcQPWweVSHBQFE4sYkc1RtPEvASOM9+8O7bdPh5RxVWpY2LPUvRLa9x694NugKbT
TBlIDW1aOYn0/zbKEYUEZjQHjyBWq4gPneThlD28TKUhRyjpKktpGjhfVustYOOH
HF6/rKZwGSyTHm8GKCAJZBcOLrhOrwc/SOVEoinIbsD78o+A3NETGOZ22DrVGDdg
rxjASTWlHJgZaATc5bnMQhATU69Qy8OC9i2N6j+Jkz/BnT+LR2j6uQxr0hA5KqDY
Zbe55wNx1Dl54gf3sN0QHbk2YamAwB0AMmHc9++kk/+/V9n1wJphj+qqtaTrqxtf
E/DLxfqyMhGy0AI9gbrBWS0KrBMf984PifclcY5NltEp8Ho5vki2ItHFI6LFDmTs
mHljEXRcOgjT6mn+mFbny+xKCL7ZJVjgKfFlX4IWiL6xxyESdwt8ushsNpUC6gM7
qSb0I+WEneoDU/y4q+pgo16pKMfmNsQQY2O/qriGgCDAA5Hkj9yfVw4wfuF8xJQP
ELhTGMlUuAgNs6cu+vT3xDIsrE6vrOGR2mJGmaj5WHmkP7dDtE8eTIOUv8dkYFeY
LE3pYxozzp+2nnorK4lq4DD06KG2TZnf/jB+VVY0ZYAdVF1LF6fgqycZptATKmac
eNQsodV6eepnzLntEYR+H2fDxMstA0HS+GX9N+3Iw0+juSQ/EDj9Wq93XEHPL2ci
Vvp2nSVF8dLgnJ3H4R9dbbWr89XmA2WRd33MOQ0ZVeQtgi5lZTXomkjoQ7MhbR1b
Ocnsqa6ue5ZhTd4A9dfW+LXksEJXNrpzv/9qm6nl6LlAFeVi5xGufbtNWiu4f5MS
XfX7cMzfQs2YwMccnD+dzbMTRF2+u++qIxoLr2dNCJXTEx3DA1JmZLPN4XquiwR2
gS8LEf8ESFh/hR3LvLHXhMzu4g4oRvX7IzdKjySCCCVfLSablDeEto8fgiKGHPUO
++rU+khdido31aHeHJ68GQ079wjoW4jYNM4kF9qhpsfZR7DOzoSAw9vbDbhOIhCa
u3DLkKkdUUBnQN6hxwPHTMTmlhVCQRkkFjP/b4ob0fud9VXG2Z1zA+BcSGhKBAzj
zrCFWyop2q3PXl+G6g9WogKWXVaW9ns522CGy+QyDKKLX+y0yHHzSBeQ3Z9Ky2qr
leHBgAJRCPjEh5gA5pqpmdoFgrKjGggVlAirgYAjyPPzxUZGsueUk/9l6MAEs1IS
K17n6fRHE4+noy6d7tDujQKNfDrsa9Nv+iOQShbjX++RX6WGecZ6WpclB8S9FL8L
Frhqvryj3TBGetKcAYH6gU7JPfziWTjLfS15FfQRENZnnO+gubmqb6IWV/afWP40
QtfRfBweF/4KCAJF+wPdmYBWgLVnXe1XV9c73NWz0rQEmcqeayiK7sw8M/16pzeC
vasecuHjeLbqEKjDexr3IUBlcQR95gsJh9X3o1LS2jbZna/OVpqPMy9/yBL7RXtC
qlSAYCRg+EVjRwAmk07Xa3b6EGGSJVlt/VThYRk2TbCzugmVHBZ+hjT2Bzs3N6mB
cbgSqVmtCt2dpvf2sO2y5tUyLTe7V5uvP8Y05eydKwqBOlac6cgFJ27K+pd7wIDV
cYZxWlxDfYM1BfGFhmh+9wmycfPKFTMm1mtNxCTFQAIexeIvFuYGmRcsRHV1FBCk
/kjs90qMDZIGfprFV9yNQF4Q50HqgAF8lJF8DRZAnfdjbBCnzhdpTbTxfMaIcKCF
Mz5cbf5Ldc+/7j/46cdmg5Nn4e9R5vm8FVwRIGGwp8KeNbdop+5+gajC2sZVq9Ot
0ltMNoDLFsTVtfQLxpxbZ/ifdnqAgxvXz29of11YXCl0k+sgFmHErH+SccejUQd2
F+zOandOXli2F2wtW7oyukEqOe3+l7n6urCoUkbXSoyHoHnDAQON9O5LpnhZLK9l
oAbzwNbQwMWmzhNVGg5An8+2RllbR2FCnQZfeqOM4opsJAl9PWjQL7Gzbs7VqiYt
uT3axy5FB/HaPC+fN0gaTuBG1U69ebm1tDSv9pJh72rJxWJ+r20P6yuiiFDZ9xA7
S7rk3bifT30C8r1JjgpKLQXT7ri/k4NnJLCm2fZ0iStstAua2KMUj8C7jSJK1poo
YesDSliAcHmO0a0YxsxeK3KkLPkCxvILzQzSiRGKvc5etKlm4WYD5HTF9RewclpH
xl8YecKm8ABsTGcISQRol5ONBA1XZ/mQF9OIfBQgKswJszeDcfvYGUTZXa8mjTAi
78je0tE33RuR/Zw3fZFRl1cKnkd5+h/hBi9MVLl9fn/bVWq/0Kvb8n0ymmL0SkS2
UEFriBRiOD4I/xg5AcH8TPAADvOS2PDmJGmVz+vVc5svLlCsy+HrJrULQMFu6BKY
rN5tubeikmhOOpIDOU7rscbvHHIdU9bOt0zM2bLEQ+yunEPByT4MYXJxEvi3P6Fu
857wsIP5jzpAB2LRQku0e42rbgcKbi2iibbVPv3Vfxf8fjkjgMa6ssFUG+WaFfwx
3+k9KfGoznT7D81P4+nRyUwSafhF8P+eYhJUEziP+kQobmavJr5uRnNyTEQC0yDU
/ZrKAcxHYKhFTs9MhmHXLRhwYSVNtGYFZQOJKuymLok0HldPqK+S81PFqNBvfrfx
HlyLqC9TECkP68PgICuiUjPlB4w/Ty+8Mw0gryHn40xrMHtrSBjeuGupxzIIZGyW
NFagPvzxs5+3eLBT4dVvUdzzY20jPi3v6ObZHxxf43Ff8O+ua9IrqM+MK4hySXYo
KVTI/2tmOcJyW7lgd0kOFFlTRgTQOeQBM4o183rP1tChXH4mFTdO1yhUt7rumhRa
cLPYqInNCklDKk/DuTPxSo4jB78PGoJSPC3iqQ32MZa0B4dRRW045yyUZUJF/iS5
MnJOQBT9LOSM6kamLOcipFN4wsFZ0F/P7/BY2lBhDwv9rLgQ7TjsSrpKRmuMs6Hi
etez/sHb2SKCa5vckE4WfoGpvoCArS/6kKwrAWnAboMMDsBdkBdUAal53vfhuWSe
xX1qRqpGliemNe/tDvgCtbrgG4F8+jv5NcCPatqj2+3nj5FGJmcWmrbyQbNfVTWu
uxVX03CpiIHCSc26bvkf2D/fZpF50FMHEu9m3voXAlq9bptNlacpD3PqYF4q3VdL
IGRuq/dyzJ7kh5pFDSqKc63BV9ZUqDjZHc1tp4MJ1Suy4ThukkbM6aq7ckTe/l9V
mmJCo15HQojYGxWCUK+/Qk3CGhlg8Xm3oVH9LnM7awWzomdl2QznTijaQ1YdGCec
l7t01+5i8nwdcz3Ycatjrdhx8/0s091B5vVxSAIU3wAEWARm7LGFHyrCE16Hkr41
Oz/ytokdFsb1Nci+XZlY7IPU47l7jinYbCbRLc84UdEcSUq3Qp5eB+7F+a9uryMw
PrdyxXkwxXednFMcbGBzKSp0/Kj4T1KwTtDALZFGb7ytMr/4BYyDfsUogF1Lqy/T
uAOAC7fLTnhQBaSWYDozlowtsxWKJJplL6ouofbzGK8KlkqYd4bBKT9exgW7K9gA
uBG9SEukjbKWQbgusGWcVG10TLVuiZmoquuFok1I1yIw7HdurvP53738CxrlO3yX
h8eIwkiGjh3GPUS6JqY7sqVYz23URiA6EZpGWfRxQNjaO3KlfPUsPCbB6cNVjSSY
gpGcyGNkGEfV3eNXZRZOMpJNCHSlMFQ6clPu5lhPgCQQ17TdjkqPjvxTcDtBNxTo
Kas1j2wwtCjhRQp71Z60+fmzBLPoTPdPmse7a3fd9XW/tQsKBWDRPrNmNXTBl41/
IOhLqsUYjNkD788MmqVFFkPdK+/B/WaBdIR4kr4Fu7lCvm11FS8wHtnQl0Pg/OIa
RGE7Au7G25HtudWYs99SHiFfPCmYqniVxOQemcKvEM68ZyUU8z7UiCgReUt1ahPh
b/uutQxczJLIysWGxo9n+gykRB6skEopGAFZwxpAhyBlj+ai2yMZaOgM2ZqYHKbT
cCJL/WPPdV5cTJFhuGryLdqYhPI3gaw/47gcAAsns4b2EOxMfO3GWTHOhzww42kn
qrQJd+0ybDhoU5bBg2UUoitwfNFxcVwoIHH1Ddw8sjgfKEwyvbzJvspWIO8JzOVJ
aMF+ZgV0I0iQJEk6Le7zviFbj3nDxJuMs43VWcOrw/AFY8z5Tjf302dfZPOcEQKs
7+2T6eqKo3M01mfIDWG2TkmfBg6zXMXYBmg4UiOrgHYpXrmL58H89TACxe45Z8Yc
kHNuxSm+Zo/pHJNFIQxqpJIh6/pTZ98Y8fyQYHNvH+if2kCYJQJEF8quDv+emVCi
hQCsrxnUokKvIuEaRnHX0CZnoOi00y6akr5BQEjkx2Nf758C0q+yppKw/ltzeMn4
/D6dCY1VExnrpfAedpJALeNdVnAIVJcIbuFfl4Inbe4KE4+B0iBhzl0xCL6gMYYn
0wT93f9ZKCk8czEC9MfD99Lz8I9BJY+FqW2dTuHYu8yCcju9PLcvkfBMaSRRthT9
5+noqsBXZHpcPVl98K0bW2CdseguW4RwNrCDgH8OFQsCR3Z/OSjAv3YaRpp699ZK
lJPtKxO4F5KJFkj2an+l3B5bCXJ94sZuIGVIXyb7QhoNfWyzhbTxvzW7WjqvKO9Y
AmJRT8DW5fqYuEXJxmhOPFNfvd5MzsWpPvZbUm8KSFgQy3CuzKlEWYjmoayuEQBm
yfi0+IwVW7RhJIgXbri/Xo45TiisenVSipPvd4LSmAiuYK/l+7QZODtyeQ68vAUT
4+QtEdBDvraokPbwOtPrVUlQgw50caB+PuTUd2hX8Mb4U4lGDraJewyroTGJ8Zyh
xjqsSpxFhxHejNtqfWXeza3SVCPDuR6f79KLEVrgMqw7x2Iv5dsoEQAnvoRehQWL
rJ+Yid4F1/czf9DOh7+MuswigiUc3KoHlcEbNuPX5X6uCutoPHdESmPJNHZ8ydgS
237zWbOc1zum+HA+Y9b6Kw1312owD6ulJv19abyWPwZz29uy+84bBxhEcaPfhpxa
JFePJg267CDvsYAXKUa9Wk2qt3UuAO+9NXYHFwTqO99DdLuTPcM7afiH7a8fB/Eh
9KuMZceySYeWqxlBEzGt+dyA3YdSL8oMZ2nqet+YuzHxLDCBput2PmM6+kAZY+1V
kXJKjyW5db5qrXUJXXDz4g+0GFc1X+3ntxt66fZzWjcEXjJbZmFoTfhltTibfpwk
gXN6AHgKpblg4MaaRPmrKPiaWIWDQ28s0SsPbJVLhrqd3Y5YE06ql+3dbbA6RO3q
HTqnKDr52rdmNNL6GjlEpCRPqXObH2J2Na+iUU/hsUKSrHSkGNalEj7OdUIKwRyo
DBXWTydc8dLXpTGvmJxsingvEO4hPP/+Kbfw48IFuCecmOFH9PXie9dANS75Klzc
8QUdEBIy7iYAWc/eUl1kvJTezj6vWigiHc6ZWRQcFPJNlt/w91rfZSwMs5+dJr3I
X5CTySfxVKUzw1rBWUxCI6k5Z/98m0v/pGjHiB6caoHmN0QuwEt47o/THTALEpeB
ORUPm3XoizEg+55QRAJAZD4C8MGpdq1yfYyOCau1D5KIB5jklsTYCORdlAfXXURF
y4c2XZ7/pDZqB5Gi9cqOhaKubuPolNAP+VNWerYZvkImM6iNyO6wrV2ng1BTDP6T
6h30eW7+v8BnzRl73ePyjWW1E/WvXmS/wSgBpx5h6PmurRYTBWZac5kI8gEZsEKr
GNEUtau5SUuUxp8f+eHlqTswXO2rSkQHMv3Rb7rpbyE2kW+E2ITh9DthSzs0gu3y
zssZy6QlqewGQKiQ2LOfEfTMmWG2Jmtq95vRAoYBKpZX/szdCG6+uOoejKnnRPEm
R+kLhI7/vzR26Vz1nxGM7ecknmcQ80IZ7jC8z2tNyEwa0A/zjOK0/hXB+cIvGQh1
cPriIEMzHJoL+ehO12m7y9ajAd2kLK0dBs4SxExETV8mLATtpJaVc74tuqejw0sH
ePXo7oYrNmpFWPTUSZ7spF9PX0+86aeBlX5cPOOZpAfdMwmza9hlJ+mZWCVeXvVM
djUPTO8JuyUv1Ia6QT6kAsiweElcLGNTaWx1juWo7cFh0jWDdsaF6m+8WEPf700n
hF0IaYXFJJf6G+EGLDOQUWAPRVwifuMhPaoxL29SuOQXgWbNTYYIYQZ7auiHTMiW
+M0tg02FZg9TQkAnqvIV0Pifr13zJuI8mNmHPI3tEHQAmSSAG+4mKKAZR9AF3Bl4
evcoK81q8ZEABP7QJNIGw7UDWV9Xpwd5JmEyxZrOFsOQznKwvhKQG3LqwCtF+ywS
tLxlQ+lYvbfjTlfOJcsTPu1omK4ZLD/5WSO4UF3ZqyqirWyJ5xD810k37WnLoLgS
RcJdfGjup4jZ1sCx5D6wgMgB+GfIv82hQ0+n5cLNQT5BsHwnFS30A47/4FjoSIQL
2FPcsIedz5HOh1vpW80vDDXCqojaAHx31GWYe942L5BkTw1YDyCFndysGS09SLwi
3rPmGicP35cLAQGB01m9a/B+SM9sj9+DxX5Z+NscYLksxwD/DVGIRvCgsGl9Y77g
AdwZKjd2uU0Je3dZty/2U4fj4Y3G9JPJEjYeydktjKXkMWNZN4QA/ARA6oVW1Tec
wv4XvD+kk3ggrIBfXqColJca6juwww8iS/5/KeJuKGt+AWv/iW1XcMAJ/Swn/Q7+
Qpyhf9/X8myvZf4kLcd3aGYUeVDS7GasMLslTiI4FPpqr6AJg3PZVPSMRN+83ESV
61+bZA0SRkqNW9//kgT6N5E4lK/5nwCvqJLGiUfrC0i8h6HHkgGp6OfussTmTuvL
Eey6jQA2S6PxEyY/DEpSRF3R7tOf4Ka2soEUyBR87KUfNKOeK+UytqgdphpV0pSq
U1W7/hrXvlSaaGMT3Ce8DAnBr9CjLFKE40iL9uMa16bGFKaMu/E2OAVUSq2vkpR4
eHk6SLMFENMEXXGI/d7o9ffR7uz71THgnAb+JKfQG2PGFTT0V84m/WivAlCV7gNH
jCxCmd+7k4S358OHn1AgqNg9xxJ1oVi02xSAub3q2jnrzbaTz4YF8TGAQAsGNMGu
1jjt9RRPD7DZpLLwI2npiNnAOVroCc6MdqdmfUFbxeTsCjRpjbyKtV3IWasCXC47
QUpeDPoGKpjSRAtuvRGzQBMuewHFxXPomQb2nqy4uG2XbleApN4hgJFZzep7vGTG
5KyfuG54qCnyCTYT8G+TKt08Hkrb1Zt2NFxhpmO2zZZAusJpimSVWr3xmeJ8lpeB
c8oelItc6iWbf7TZcSzvm9XboHtsVSDMw8Mv/8Ik61kjyFNT5/cZp0vdk70HP+9Z
SrpDawKbBTm/v9Ihl4tgSRzqvCkwr7RJJGlazRnKDNOf91QQrep5ruViUb/BTmmq
hWqFHmpUID2MCbb65HZABGYLx4fZdORQPAzm7CwlnuQr9tmF2Pe1YhhXVqANDV6z
TZBXP1IxkbJ/uWjv+E2Tw1lllI2U0QH49DZ3FBWWo/AH7kNY0g93H+veTJqYq0PY
e1NZZSlMCW0zECZFmQMKIEhmavBZ9Co/OzzbZDWdfJP3RTGIknEIMRQf/Yjx5mS5
1j9dBpOA+kB8qIVCbs6K5pTqsgx4sXuyPIjeQl8eZR4soqXR3hm/lheaGledCFSS
QJT36oWzWwpGje8nPSI9NAzG+SGagWCyYNo0WUG8je9YUdq/zq2f2zAnBOTK4nW6
QVGNzGq4KZ0D65vFp/8JepkOb/b1mL9xRLxsv937YhqQMoTiR+Gkk57/ivkLzAkC
nCS0CAXRUBsEXB67/PgsOza6zrnGgpB2V8oL1O8lX6HJQ5o9Epq0hPoFkT1qNOvr
adg5DiXf9v5INnybPIwsHrrT73BZLorCwKoLyDsArtr665m1N9SUvBLFcgHybs/E
xel2ITg0NYULdjfy2NMfMlC3lZIOFHNbqSHHduBesvp/wVKXYnxGx+kCv4IaTunG
CBaRbBlhHNf5YpTJJNh6MCV7UKmz+c5nvg4dKsMrFppc85M/nPJ7kfxXV489wmLe
djfA5h4Bk9BGKHu8s7/8fDTB1WmFyLOxDyfsYPS5rqPUwodfJuVzF6P+bxVqvmg9
xXz5R8w4Rjh3Dp1Tt1O+/83s4uJ5Czz3YNezmEaI5CAzulCg1t4ub9Rbcss1PpVQ
fCfvfCSqssdFA8GPJlNIF8Umy13SrjStK4aau6MiqlgvYkyx36dT4mcxOQoLtq9C
EpVLcLUM5MOLOPhe4TvxWNsGIFv04hGnKeeyhKdeg3Do1dvQF+GpPsOf/O0EQEsh
EVfkoNutyhCemXy/25IXVLoKBZziB6GOMERvzKEQOZkDDo6bxs3uZ5ahDiyOr5AH
J0BCutpRDIob/fDjFQiLjzlOapg4Gmt2uZrtRWvhihp30F3U/kWXcVpjtOVvqgyY
8lyrZfIX5xNd4xULbD4owa6hIykBJpCgRqypnsa3Yg0sDKCo2K56lR/QBNDwOOko
SoKKSISUHVKRmFoWlWZKMDgdwe1vQXV5qHwd1QeXoWGrdUFzCTSyBayaABaDaNu/
MKUeZ/LzcHsjfiREwDKXMb1Z7ndVqhgmHRnpvrXZSlw71NNKFEn5yIOXTxZWWKpg
vCE2FU8HPUhZZZ9WZQIrWJAG/G9tVsiD4BlCaaYBaThVNn9xCR03I99oPyLv4eyh
kvKsBcmO5yD0w6xg02+KHSCoW+oiFvW8NCwFQr4L7Y32pF2x53170SkbWTETZbVm
xyVNm26u4ydhYVORmGcvk1jG/OdS0ieetPSFfMCi4ZQs5kjwtyHGePcPl0da0bvy
8wa804iIITxfh+SaGqQcgNC337YKHPLyKU5eIHndYd0bqf5P0bhD9OWHaFsXsCUc
zX82fwbLm5/Y8ITHzgw1ZWmbepN6UljNVzXJsSPUWBaYsm4Sn3AVtexhqHwuyUH5
Sj/qkP3/a5TtIL/RKmt2CUaT/xPZf+i0OW1I268lpL8Uhd1T7sPldyp7Y9MKONm9
tuGRK3V/FffKGLQp3llRTuxUBPTtXAkbZSOd6SHINNT1g9nm/wxpzexClaBTxgd8
1RALWYQNetge6QwNrjG8TD7YucZgbEQlN/+sD55ZAssgcrgsHF9FBKzgieFQg9tJ
7vqcKpUwyLpCl3pYbMZ22vrjlVG0+F8zn5DX0mVAedWJbLkTxAzFH50/GAyEko1R
H685kntRrFZhogkqoNRSLvE5JThvk/n33ZezdLFS/U7Jmtzyl0BtXc/zoi4YW3+e
o9K2rSAKV0YeqXRdD/WFACmY9/CGFkzmdxIGgzXu4pPHqLGDUDE64G68Xk9rut97
43IN2DcKbk6MfQzxQ4PEBFnIKhPS/uO2CxNolyTnEPlf1yWl0kTOkz213EsuwlG5
XF/QWXtxf4kkpuXzc4kAIS+ZZhlnkfDnhiLTs3b4XfUEnQtT0FfXQ+VfmZxcZ+M0
LCUqsCY7idVo2sT6WSMIzVbKmoyfct1fqWruzOuAG9rmXhFXvgxtjiaNIDjiZiMB
Lw+VXFlOiFkEOeV/lrcRIJK7mOTsmeCGWSjFl9/ZcfsNiruM1KBQJTE930OZrtAy
tZiGjOY93Sb4JZqRZct58vVuGG3UkPU2VSREYiiMwXXNJ0ryD50cLlYEcjyIxk4+
kEULqEg5ibQQQSAWC7iIHcmfwy1D4tnddkJgmPCyoqPV75AjAhntOtyXMVvPf+lG
pMhVY4C3ZuY1K26qpc2tbO23U0ctjgSTg4B21kFT5BLYcMWuNrxpFGWdevXup8Zu
tUKxa38gahgnVvaNdMwBxIerU779SBWnjORWbZZ0AasWDP0Nmr/zmFLINaYS78Ox
yO+9B0dB/4bujpWxnxRgzfqyBtbzmRrwO7tklgSaocMqH2ZdaOeReLRukbiFUOcb
Ot4W+uWwHQpvTs2SW6p4bpklf1Er4bi5Bp+YY7VJZ0NJ3+3cKBJltx1s2jKjsq+E
lhBa9JpZoLEkNN3iv0/7NdPEHJ5G8+ka3v1ngBaIky1xUfbCkzsZCv4eFDUruu/d
wiIUZ2MsyF+nnjn+BamTi3vC+OXL8yEOCMLQksB8EAPVQ6DtZX68GeRP1uLm7QHG
anQO/GIep1Fu6h6zJTq1knPP+k2QLjRN7FYL0fwJj5fjjzpt9YYCaFVjfoJ2x1zY
3IQN6npN+YYJjhjdPOGoH9heKsl6TDtzn6WmCbkTuu5fXJxsfN+Y8WmAAR/GJ4SP
+txr4UNwvYLhrGdXcDyY0x1luDs+ZpTyUqlzMoHEsqnawtCBvITt7uNCBgPqPnur
TMWOBnz2cOOXJ2DGP3yJn644sUoU5Rlik9Td1VfdtTqiggO/hKS1ZURo5/MDtP8O
nM95EnzLappZBXeYUddrpbNtelm/MnurNsJ+s/p3UeI0q9KN+ISke/hQXIERf7gW
KFzOAhcPsTz9bZJxlBHW/+bILrXytWXiNGPLnt84+Im8m5aTWGdLiB5GMS/iIF8q
gkh4edfRNFTsIttKgHqTnsRLF1owmEV1pz3s7ayfmzV2HjD747dkumL9uqB4BakT
dRUlcJzlNR+jf6OhEtB0rCF+7TtVOvDyPaHi2asHd4VAMekxNseYf3KAwjq0R8nJ
X9fe9R08Wr/pd5VrkTzxdO2UZYo/ZqSi4cLhnnMf/3RMoCUgp5eGzqZEPd01Sn5U
89HI/A7viwwU9zHf5Q9ca4hDuE7kNYXGXoPtILZNaic5ZSVKCP60ijQ3i/4OOlMi
xNBLl6Zwc5U2SW2kFll+Wyc2rVnb8rIFFJZkeALC86cbbBTQk6v7sneknBPik+Rs
ZVmNbxobOlxErbZDc3yraCjAGPq2fyKTa4/7hVtRN3LILT12wAlOjWcm+Hm4PFl9
pjdqF5iHHZjz9dSYFZ9XUba8mK0XFVShCazMi2NrFLIA15PCcboGL+LLT0EOjDmz
ZLS1GW205ECmGT20EXRpG/pc2ZVtcojPP+pDFQ9myWtgwP8apNBFE2rK61who9hU
2x5RsPv4ZQBs91sjmnjWysZ5Qzv1PYVXSy8g+R5PXxcBH7udOWZLXDpY6QMmgWQJ
001Q7mmGkRxmYQqDBH3H8vt7Dcu3uwQoGRuDTMiP+IzGwjMVMWupgFmNO+AAcFuE
jfNEPxGxAB3ECZYx/MHZcrjwB2DV1Itqy3KJ8uD+AGj4cQjzr/5UjJndBkRA5UcX
8bI0hYUVC1PcSJzsuJbBAuJrZBPQ+7SSTCZRSFylFOkNkhnMGakXp66IoO+Y+TqY
/yDnqrxiTciYBd1m1VGPy2aj46wuFqtnYqWsM9ISYOCUTFakseHSJP09vW+nXMRJ
BkzBOnNn7Dtd9tK6pUg0k9T+q5mxqu51C/IONQltReuCaeD2wTxpqTLWnZYj19BM
8usWAE+iFaTzzqrxLuRHjBgUl27U/Mf1bcDPJ7N1hxgZ9qri4gOsIMSrI1+u74E7
l4v4yjLV+RSLBkaxy1YfFq4X3f6SS0zW9xOed7aagxyvfcFSxH/ysD3ZaJqc0QdJ
OGiUBUd6PIva4rX4zqQ1LCaRNOT+qQvQkTi+u5xQ9dULn5FUsHD31YXeeDcMXBAP
vLZnuPBf093yJ52Duqd4K5buH8De0T1ft7tqtDUx6PLBbYcGWmQgdrnVmEC4nsOR
7pjxOr1o8rWpMJOLFY1fEsf3Fgni4cDckLTU90/o+1ENqZZh6/Y4oKcxHj0gMB7Z
OxmzaI7G5Ok3xzV+hSuaPAvBWQSfMe8WHqFHJ3iyqrT+6xjzLkh88Hp8CdBfBOaY
LQ7kc/HtK6paV+H3GdG/UjWa4lSC+Ba/OCCLWb2IUyoNmnZ+GvHWMDjZJq5NhbRk
WPJb2hHjkvVcAyUvSjG/j1032CrmcRI6kQMgk1fgnh3y2Dx96uSLtfVSZ6NqlmDv
spfLEulXwhN14u5FJa2CntYeQD/2SmKrNBmes7aGNcMzA06DYH9saYneX6QflKvG
mvzfxqPVvPQu9al0Z6ZG6z16J2Lt4bo9EjOTHtnts6tn9o1WP0FkpVvVQCC4Lfgx
OgM642qCibF8TAs7d8k/tL1r5Agj+NYLJCwymzUF2ZPpGA4FF+MrV+4hD1AP78vF
vp9Dnx1l4B0cf0rq5p/Qisq3pSUGPxw6img/RNWGfs8MSYQpchOs1daT/Is9kUNw
zDJ1LygxBr81bXGVy3VNOq9cdbPi+sSsg4QM4i+jgR3HVjeTIHv2/kavYuUCxgZf
yv3xY8k9r9VEZ8hjj+zM0ql9P8UKLurI/x6PaC2C1Ht5k5i+6SDoGV+dAJZxGDNd
HgeHvD5c4k48ZZoeHNo5YDSCn349ZpLjs7ToJOQZqTwQ7bWBfwoqLwE4azkJObmp
chHn7g7BT6598s9+EiTJqzdosvdLddOAVy63nr9acJg/xnEk1CA7GMDZEI4pYNbG
olWgzalJ/poNP2YiM+NHl4YuG+2A9MEWA/Tv8YiuTKalArYE6jtHqu3l2WDoKmTr
IdHSBRSCeNg6WJ813g5PdOLPIL7ZPd49xXAs7JQTPKmnHeYQeFDhoQe/7z4ATdQs
7gokNYb/ztAarebjok4582s2V2bJBPvXS8yPsXhPcd0+z8DhmZcfUWKVX2s7iKEB
/yI/2KJxXzJbm8TmUjF0WFhJS+s1ocHgeMq2h9mRtYaSv5Tem5qp1Ny2QUtte6dH
xWwybM8X7HGYMhcMC9BYjJwO/wUSVaVtw/ivy5EJkblqCu21ezwmRB/iJbhr0+lC
kjQwNYkWKv1OtvmBO/aI3ltLMvoDYHPlM9+xQFndD2PlIm5C8j9HM8ayg5p9W1NT
f0yValAl9m3Dt99gZXa5iyh2R4fpd07QJn/qELz6Oq78obZs91nZ8aO4TSx5jr+D
Tld1OR35ce5dmB8fKe6uGi25+dGg6bWsKOpQYTwLPRG620eYLQJWPSSVf8AVn+Wz
JJQFhFpo+Fj1wP43oZmMQmyO2yaIqs/1IyjM5BuTCgq7iBWXFLxlAWbCOQwgKdAq
py1a1EVdFYDPAwC+58Du+6nr/eP7L89jdkht76+qYJqB0DBFH3Yck/Pnym3juGli
uojUbmwfA0xcUba9++k/kaB/eG8ba/Pwdz9ZQWW8mCBq0smaCG1wJAja9HcctubS
q1OGxjHikKKLtCPHx3CHHD+gLV1UOoRxdjThDBNohT6QaDCXHIrZjJiMgi0wOHPI
vIcgPTfDdqQ/g1b4K0mkkxy1JJZ6sKvUSA05I2C9gqOFSlfS1MnCtcr5/0dYcK0Q
5SATRsjiW5YfzbkA1iyooipGZpTxmvHaQkUUFbpL8TV5sq5+LqGNPczRjcQamyXq
Pnl/40qsRW5OBUxbXWKVvKdO4cVIWPjY+21ywFTsT9M=
`protect END_PROTECTED
