`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uH0vJKLfVycfyEiG4F108IjWxu6rbWw3lGg86jdHH4cJkmEZwY3xTat9pvvdrhsa
/7CZ29Qf2f/4e0x34dRMzt2QxpVsB9xT/n/UuG6dn1EucYNR34+6Gd4uwdMTJNwG
RQqahgtpgfIX76MG7NbTLiWc6LxQlJi5W/+u10gmPeOQi6Ohrcdol7T++HJlgviH
dEV1vFo5a+eTLLdFUZCFSTgJs95naC7quo7/RAZgkL3MIBSCIetqFzRhAf9Nuq0R
lS37ilWWT/r4Rlm/t3ixbcdiCPpQh4ak0+aadoJj3Zmizku1Gk1THJjiMiNUQHaP
okm0hk3aEdhE1Y5a1DRLyDqsHAuUHWJO8mYzvx10PWqPpfiCf0ES/xrwzVOUImD3
VxDPy6RcEvhQ1jJv8tPRC1iwXYZJ0t1/mlwrO+Keuq7Dg32GrJ87bb0e7zadhhLU
jR15iEVyC7j7tp+I2A1TEw==
`protect END_PROTECTED
