`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4HYO+eSkswEsnGF4/Cmbs3RDYt2pOntmEAyf5Y1MBvmp5B9VNuCRIzLc/9pSmsv
MteD/1mWjdNbYOezgOKcgl9UVl3Y0MD0m8GpZ+Ow5svE8H1FEpbOLobA462M7KOd
Qu655spWDoUkdsGYpNCuat4E3bweRzqTgTMIGL2T1irqEpRZGxatzqu4k/ObHgnY
jRYynpgXiTpP/w1b/achm7n8Lh1Wpc9qnIc6MHSkFxbNOSwwabO8XdlQKa4Gn10A
J8GYlTo08w8r/UMMxnMgkJFDs0gNvFoHNw8Sl1e53VSAspnFlq+nMrRYZh7qWjk1
Moes/t8ckD0R029QYzcktBf4AR3uah39MuX23DY4lGI7R1IjePEXMduYPnLJz5G4
Q0kvUIP5PGnB1R3WXZMn/TDBd1xN4rHA33uLGTWB+tSxhyBXo+5aU3qNpHSZY2g0
bslhYksLTUYD3DCXYEyl3/q8ZQO5FQUe29PyUGjNhyF4tPxHbpBNgpbIWdSY27PE
bOE1WiDo1VbA3csrHpdh2R6lRbkoa9iogy9dmr3wVbE2oHjUXR6PsYUD4C0XMM5G
65XkFZdOqBQEzz8dPX5+qEtr8iWCR2EQmaiA4evSh5xc2dB4H45g2GM722PfQn9t
XaAMMD2LLZaVKjSMRjbFCj04ZsWh+oFSmcGyyp4l+arReGpOyAInz5IyAVX3FXod
OLNdhMlgxwlv1bu3pSSWZ05PrQ2CRFQkc1l05+YDYINa/wCCfxbFozPySoKiy3VU
vf5WyZHD+lysOsKXmk0yMMIuddhb1FhjFyh/O4ZZ+tu6tfOnS4RanxzbzgGkY22k
Y1PvvUBR7UodhOAWoiIYyl7QUgrikkmiz2wES4cFHTOoFom+lM50NCfWIqihdjQc
BPxR0178L9/U8MTjSW/jXp1E//4PWfRgjyegPwk8U8mDCqzyoUFlXReueRTnQq4D
XLIcZpE6aHtpdk6j28ozYD8OvFTNMSznjcil3rKnE3Gvxjq/WX9n4+3+zB4IngJ+
abT5nU0VXycFtME9NSo4ApqUb7JRua/2VXYMMprOC/qvI5FqFdKnMLKjWOkRQe7u
1GuSpcnT39QG6peIpF7ikyzZG8LsQzGT6iMHBuyjtrMWDBHUC9nHuocF8+pgxKkO
cN18vwRNbB2dpiD2VX2w7/7VQ8J2DYSLTwhV9BzjTDtGyYlnFinZ6j+wdjSyBFDC
6CWcl5+skhSssrXoDDlw6Kn8ZzHDKLORz8pspGDNcExs02mITQFWMt5QHuOk/icP
8k5ft8ani1IerQz+lhRLXq11G7Nsp4gZ4QPQU+ql/o0gIoq+FgjO5jS59qMYnife
ThhRXxcntesE3yRkPS4Q+MQFCxhowVCPt3W+3rAjlU8kwerBLaCxM186xjv5Ru9z
ye8dO8BKDX7ZYhR/sxxjG29WYgP7EmMeRF6TgF9zGXBEDqlkPnxamP/VRFS6aayd
QaVS+Lmm5P9JPYbFVJT44WFweentgG9YsR4IFr/Vt56RMYXpvQRSi4dB0RUFegJD
uqInD14t7U4cgKOuwJYgyOMiqTRboJH0AI5/EoSdnTgu+mBMNz/CA2zO4OCd67EQ
MKUc52Q4VGKUomiZNfIGM7fKO84wYBm5jRyliiRhCLOlsKGXTHRwt6C5v9Fp2F1H
fsJULMG+1wjaSvPI46F7dThqZ0MYkcHWC4IZj1ndonMW7d0nPbUkNss5LrltMia4
MezrzX7HYCRw93g1aKyrMBvDFR4/TWkZqpQ4KrpiEwK2nd27nvzLR6WLXU/5T5FD
D3dJSR8OynFz0GLZbeArySrIQspaQU9LTms2WiuZmFjXyLVszObWgquf1gIuKbFo
W0RRGSGrvrKfIHHwPpNxUDpXpGIWBVrSdvFSV+gFiE+2ruu1osBUqtUo/e5ycwnM
19PkCSK5nKZdl0/N+XY4i9cyNdg9VTBhW+1hZtabOr80N2jAO07kf1Z0rKk+Xl4B
1F43ph91t3RrIqqQzWLToETzsX7E9QlQWLq4XZjdf9N0VHXDjuX9Zu4vfmAHvnp/
ob4J2UG9Vt8Yih7Wezq57X7rIdLTTz/za8kwQZoq9OdTwqEVdFW/h4akRpeAbjQH
RfsCEH/Xae8CxMtia7C0xIoDjGdFxV019w1f9NhUXjlUZMRe0odrQxnx6dPNwpDZ
`protect END_PROTECTED
