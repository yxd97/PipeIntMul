`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbhfXJ9Q/Fqtpz/E35yrpu0ugMLCJ9UcN/ACFKrHMQw+eEHEbUD9VZd3XqaSaVaS
g83jTJy0YVskxxIUQ6Ynf8ERyRAoqqe8Hde8PjBSPxQ1tMX1qQQvERFWZg3D8cR4
NREB7JoG7ISOum6tzknrXQCA/TG+f9CwKFGG3IC6xAaY/kT+n17urzPNjD+l6m6D
T+3vx6SSseitCooJLagN703P8vfGInwVJZ4wfDfBaKybpvPBQD67AV+dL7qYPfrd
QUNQKw7ueRrHfSIvUeEBCVx+PIcs2wJfM5RaAW7ubphooN1omwFHMU+HTr6o5Aen
PXKZt/wwhwRKoaITRWuber5F1KgliNNMogQ1e1AFb3kPU4Y5Hacpg6Vb4/Oi4L65
MtWnfF6r28PoInoOsgpe6M0AfenXypwXho26F475aH8HIK52kEHui+Li8r3bdVGI
6sO/4SZek+DNKg/Odvl8t3zp4R7q/v43hnz6rdRkOFxd9wVGlHk3FuxHtrxWFSW7
3rLM+9wxqarUrY/ibbZ9faHAuT8WTFe+x+HmWDOFmPCb7YE0507qHWisZhYs+ScJ
WyqmyaOv+rrKh5v8MqfG+Yrc0lbECHM9Iq08TXLMp/0ZtCAetUe3a9aU4MiwhAum
Sql3MD6hDkjQoVDOQRa3hUfXjGLO7S5ZohATrW39+AYM+GH8qkLFbLmYV+GEDLTc
wnzdozGbdzPPwtr6U3emXFS5plwAqQV8Pcf+zwUQNQef3XKplNJY9pwVKutBl4D9
0cysYh+0sFvOXJ/py5SFMQTfgCYgTBiLIETftHZaolK5uPxPTKLZwniNHRSmBh50
qj5fXo7b9bqkDZA1GaNA6zp8ILUhnuJfmdqBsv+VgZjucU4fe+xUDaXD31WqXlQD
AEiWVMULJIAP+GF+k4onxCNoZkr+AQw40NBhwqG4SjsxNzTDMGF8NRfHDFOpx57/
m+LCjvMjDVFF9J1bhu+KQ2uiyJCznmIqjlW6nn4P7YJFe5/DCio9yNlvyOlgg6db
3FraWh+OxePrF8Zf2LF+foRnNyPg9gQITYqnBNKzFfGR6tKAMqqcSwENz0t+aG5l
Jr4hz45G+QtFWHJh8VgnD4Q8L+/ZvZVC7Y5OwNGWyW84oXIsAXE/aEhxgjsiK14f
ozLK71yLOWwI9FM1id/rjxtHWh7GhE7zU/ZDvGrJtq26RR15PxXABZTtrnLTKlIa
SZuAAeTjYdoRSyKzZLK2MIh46RiLZ/6IkDBSh/SuR7T5cMJcDixsIDNcJ4bX+vgU
dQ2bTWinD/ka2bZz9U91RNStp8VUY5OkAJVkP9Uq5YNHqAAd2X+9RdqPjq1C3sgq
rdnr5ivoHEltEJ8c7LmieSPVvO9oso+GKz0AmzlWLeca0+Vmg9E8JXaOLWDDoNNJ
Yp05NZGx0fxYPOjVbIvRAbCsFDBdn3hUWaAO+JUmh1rr68RQRvPHuV4ak6QuhP0S
T4MB533oMKFmiSra2kcXhWiFNsdykr1G0DZAuQtiyTsSoRahZ3N72KGih+gSIv2A
YRrUW4kkxmjtsGG1h+sD/7eJpdVMoh2c1si9CV9UMSxUnAsDoZMbOo8QWcLBoKjd
aXmVN4NcQvfFd/hrZ3IUyBLVU+rCFvBY1sZkgt7/D/tATCoffSKLv1e3Gp7/sXCE
1AquMqkuXvIBog3jPp+nsVogUZqej2oP5HSFSYZK3jDy0WoPW5+OzBFCd65t0GqC
K65UQihtH0Q4GsdW6o5JtRvZ4dHOHLFwy7vT4TFgghZycwg5pOxyqibSMzvGxeQl
qgAozI1E5O2tT2xvZznsBdCwU/Tk2m70dyZ35MjlA72bAio2YZ3hd20Cf47cammT
6aoYNr2gfaAdJ8vnSObT9n8ezRao/1QF2bOhoIiqa+UOiK2UfFaimUvzAnghWC4a
VI0rsjg8ajahZxpR2vGL3wsOwgQsqF0OaCDX+ncYSrShHhq1nB+r3fsbj1qFpjVy
d/arL+17+RwGOVDK5qh5jnGlpUlnmAkYofnPFSuaYgyBZxawcaOyRAcX1GE+o6wM
9FN+V/nC79VlMsXd28I7YSPJw3hZ23eonP4qht/FOtJS2hi7uqn/KMqiOcbT32Gl
ybOoszZRZMl2QYzQurN/H6S1NENSb1tMHCm3TGmxeA/CjC28O4iPzPNvDLW0MuaN
N5atuIWcb+Owimx96Zo/HDT62siKzpl0U/na9Iwot/D9UJRwgGQ0xXRQh1lE3vBd
SWPa9sSco1m+aC8Ww/2Z2OCpH3rAZgfB2MmTfrXOB8OqQsxfmrODeVJ/IzPfLYi6
H4fm6I0PjJbQxRFq2FAQ0p1k0nqNlkWX6d316lmw+Kx3O/or73ITkEihYB29Tpjl
P0g152lM2EZ0jVY+e+35M8dub32M2zhU8N75drl62AsAGMwjlCHVBDAcYLE0cLE1
xq6TIN50zI53qvNLkEz/i3AKCJ4ZL+Na3SGYfiERj8YVHWoakwAzD8ZsL3WO6Ut4
ZZLCMVFvNabqg4vM14veAL9/EWoiIZV92+saGmYsGnh3YC7zMV9R8ZkWAmh1YZyc
Rhj88PjOCYMFAYzDyjN5WBPVFhi9SlsgoC032MzWb+MDjjasB/HuWTM/auPmM5ni
iMNFVkKdOVSgRnto5Rw/ec6h4fmAj2icdWXjwW7zgn6hTGuxOxvVDrPVGnTTwjfU
aLPDRYgUwpEZbKAnU4GQfo5kwcCaWLdrVK5v/aMYE6SdUrujAbtVBITM0PR+Uapz
svFWPW9XiiRvGYRZ4AXLKUoPsfWgPhpp/VCLLE3o/ruleIXvZdEvvnHyoeYmwiLb
tYYKmnLcNIaljAS5mK12BaHnRfvLFw6HYnctkGknfvqOKXXuC+GGpV2d1rVPk2gL
pgjzK90n2xTOn305oXraqIJAWI1J6MObVFfH/VY+E/6siweyR2nbfFOL+eGECt9g
mUbS2H6x1XjmcVRNmevoAlZCqyX5JfpjSdYELuUoHSPgXCGEm3TrT5G39vAADKke
gLXvlLavVBMAkXNixTeTqhiHhB7QjFbyiCYCvMz8P0Ho/IDwD7Zj343efbVjJNia
`protect END_PROTECTED
