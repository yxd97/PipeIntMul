`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PSzUX3MpSZIjSOWqoJJzcKWsl89+LFkKOxLd2DTLzpHWKyQDpxGpRey+ROFGd26k
G0sYdJBDC0rC1Fs3bIJB+8bDyHZZmbW8M2iFjYJfvbEhE0F+GA2THWXEBffqT28Z
V1e/HkxNrIuoBcNNWq2dJbNifIACqJ1rP+yZ0F6YgYRZyco249qVgWEyyY4UwJk8
mwQEyNshMx74teHy1my+NlMCl+gk7iGi8Q0UYWU67QhhhK+LtNl6Sw89IgdFqax/
WKCyvvdVGl4xQ5P3q/jEeGlD6x8sWjlgL8xayem4kw9z5jfKilNHVoME+u6hfF3Z
KsFNs/Bx4oDYrpzt8dO4e1JFwSjnjHspBe82kg+xsh587PjbRB0/9G4BgAkXDL3X
rK3TTeRMUb/3spG8IjkeSAWiMW9bibEcd44Fv18+1p2+cRXfeqr5fyUscOqKbxO5
t6TFiL5nnA4HjX6LH5s+iJVtz5g3yoCRSHQ3mhIlAb9haRtfJ1t1bEoSbRr9PTqB
hJNqytNA+pHaUcorRhEhLVIxMwI72lKenQqNGb7Mkvfs0I/s4rwtWKy3pqonEmDH
pPE/wQfSn6SeA4V0wyFiU1AS937LGrK7XOzbisN3vXdnsaHwPEeqK54jox9pfH2r
PLEEEUAj4gnzV0a/081kVoPt6wssKCgOU9r/WGrqDI3726A9jezeOzqd6r4UPMvG
zqIVFBYuRDSWzjOACC9u3J/89J+Htq4lJRbd4vdj1Y7PT/51b1LlhIYA04WKvgCo
K8CtAWOwIPUks6i1kIsNd3IMpGlHltaqRLiZFddoz1PeXnEkVVlEnCwC3OXibnC+
EIR7vKLXBBZ1yRRE9YBkAamv/ypgo4ncncYjFOOH9ilDMwUcIFIA8FLaIO1qQLQ8
MdWkvvfqo5ieVIWiMWWwztOMYlWLxR3zR/5Vru+sEryscY/kXZHLhSlT1STUDub6
IuwvTGVDsjL+xK2WKDqQOLR5nflFNlt6Of0eHaNGDX6ahdfFa7vA0YyVbRMTGVnR
bZXEdY7IX7Qsrg0+6UMCPztXVHmFJ4QxKKWF11YdahBbQPAkm5LCbjWZzSKQ4qlv
yORxLjPk/Xn0pWR4zU4ftofeb/nMZfK25oHqmQpSVsbTQ0bziqXszOSDAMzPr02p
Zvg/r6FUFWe9iArAJndjAe4u4sDnuGTRTqCo9FOS0JaAZEsJApnWFHuq3OpTdsFP
H0rHumiON7WgkOETEZWARNj8pc/1Fc+8CA9/No2akHMHyqq2RJHO+GtAIAu3Xht6
JCyz++ti0H/wvWAeLbBCsIXDkvF1cNoCT/AIXyiRDNjDR+JmPFX91hkA/eLqXvTh
4NLr8dFmriH0Gz/ReOnwOMEkYvFT/xgP6iIOtQ513YoeOVRJBnOmoK2asEFKnSCq
14FsVWh0gOZhphOCUdinZ4Jt/1UxE6nkbxx+VkukFjRyIjDU7U3PSsmY8kSG+dnL
3/WtMf5qFtvm4Y3giCGHe2OmuZTEufmZ3mGnKYIcyFwuHO4dVX1oGt5pX7ATB8EM
FJMFxevjBiKwL4kcYP4Bv03Nu3EdBOpAFBt7rgAMqRpBU/c137d0Ztvvc4TIkmAb
jUx6azPz6zsK/fNzZTSjh8124cqMlRbTv7G3XzaD2uJdFAwLvvPCD43H37Csk2DI
yRmJs5ck1fP6IAomNMkP7AYYxTUW2vrL59CAt9t7mCXk9HlQij4MroUUAYDh+VtK
agsLY+/18B9AA39b3KWGJuSreSsPuzgTah0fzse2I/fhkA2fQsO0YBMn38EdVuvg
WsMOGR6+wihv93lIpym3fsOFBOWFxM1WG3h2wSglenC66ktfHYKN0uiChUTNHVh8
WyCA+/liK639gbh567gjs+Xci+UYQD1eo2xRqF5rygwryKm6EJLVmW/hQk9mQO7j
f3uZSDaPppbTF7WUR3gi9qZJC0ZfuoBOkyaUDY67OX5LQSfP+qkeh8ECVzd58Ne7
NDr3mqsVvmsyYo+JImdlEmvLCyMEmXNWdRmbtE9YwYv6AK0oFvoVFbU5sHOZ2AyZ
qZ6GwsqSJWyVAc69MmzPo90jzuC1C8nwxTYaYIc6npQPU1xnJyVM3CnQehtCRrd4
ur7ZB8H3AuoJP3dDn0Hq7cxSR/lI048Mby0j/IRMyUqO34KbwvMN7p+Rpm5tb9gq
KA5YTHAB8RAdV2ZRjh8ELki2AZjfroOeiRwu/w1/S0hOW024ztO85adN+VoE4WvY
WxjKfvLzo+LMyw6oSvvJhZXFsAOr3usAzlVc+v22dpWsm10FESiYfQ/O55++pK17
pRV0FVrwjS+kApgq+UICYmHurzVCel/idE72xp7Kwn/3M/xagJKusMEYu+hBwOeg
yDT6q1lU9RwOYaikURmjQ0js/f+ZDsxTa2GVj47qwJMn1kcNN5aQIBmeE11vEiiv
8iQ8WrMy4C60WiiZbjANpF3ZPrWv1Of6wKfduT0adCZ3LwPp1uSXflsexijUML25
RfSJUx3tPPFCMtLnn6CNLFTXk81kA3qFlBefbCZBseM4z5n1566qi9WEhW3dc8qo
bOnM33iVRfcHtsrwojMgmOiERuKelkEKITWOZkErJ9ibKkyMpsnTjjNT7StATAnj
QieZE2YcPd6fX0jxgzkm5QxIQ2oPqXDiKaaLMAqtVvjuR0LbP6Z9qHgUYBpNcifY
Njoa1O6bwdPvjcV2COW+MOcIB23BHVNliwyqGvb/D9zRiS9+uKMhFaChFEXGC4w7
Kv0l9sNkZMhPMIXU1MU/AFwWjWHWmAyRqyrYynJ/Wqz641Tq2951d0U8eApCzPG4
YOSDoyz4zRVxHg6Fb01OsEQH5T3l70S6wpaOVfWV/UVO/eSDUbanXa9h8sc+nIdk
kZS2nFKaWawIzk2GERU81ozHSIwb1n0oLRAMLeUmAeSKmsWQ1NQZjgZi1oj6/gaJ
p+LFDcrvlIk+V8/2EJb8Tb4/9gtWaZRhKBI0CplBomv43hDKHW/6XydriBF5cKI8
2zVAQ/3/frFC0CghlkMpXUoZDqo8aCIsA04vFTyH7UjzdP5kzp8RadoEEEKigWgu
LkcI1DsP4cgHhR0rMmTZEeetOnCwh2u5AXfQP7a00/Zqsae8HPRh51U1mlbFWJAP
9Tq1fo2MMBmDpAnaY6AN7u4VaiIY1XBqp8L7aacaeW8ga96yDHpzuhzBpusW7gL/
9dkntOox+DhwtUksNUTfBh4Mh2uRvwto8sAXxEg2kt2pL2gI7PIcYM4qOWD6nNKS
GgNIfxCjDicVfDNPpyxFwpP7N2pU2tI+rhYZaZuIq0TQA1X7XJiNU6R8uKHL68fE
wtOnB3SkND82O9HM5zT3PHd8d0SgxQts/HkH4zCJ0j3mNKzxBJRmlHEnVeiJ8EmY
yHYM/NwPA5xn4RhSXKpCuoYL6cQgzATLotFd1w6GpUL8FlkOeExBvpxhJuaH83dI
kigjd1mv1rRhEIqIjoWKKzxA0lVUoyMzUDqmYqJr3F9bZgFII3CgubHnEC97f4Kt
5h5InGzC7YZrmEasOTX64EqsfT4WsZNZaqoHw748Bqxl1vx8Qv5I5JTfFCx5O9/3
vs64yNAo+APM8Cz7MuPtUKEXPSldGLGNpTSbMjW7Up4Mr5T6wV8Y8vbhUgob8Dbk
AILWWmf7AqSKCm8z40Qq7hSAx8e8D29Snnep07xJn9sX8lzgQ5SyZ/4pEDVPxd2t
jNtQtRudx6QFEDydQh5TIO6+uPTNNV2yWrllOvhr1oyzHUWiN/XX7YKcyrlfI4kL
iFkoFWroFvuveYRJInbVf4+NQYbJRIp2GMv+YXAv7vTDCAZPhimjJO7HEQEVSI8N
uB8YLAEFfoNGwh5kUapR8D5fEehc7YdgifJNCBjK3oPeFiuW+t8OniIiSbFS+FdJ
WWM/pVfEf9DiHq5Yrg1OWR4JxarOMoQqC6UMgUjb/Ei6l6Re+wIFHCuLQhRIqgMR
vSKJgwtyUbsGCxY2S5tP4PCaB5jeNEWbYDhnK0NLz1Fddh/L5prjzFwLEzifF1KN
VOGmynSG+jZMffUqSPs0xrcPRrTtpHq1N2K9FdAqCyIjwIRWqHu1t+XFrltYcd1e
v1nQpHRmUQStENyhzYz4C92+tpEukZcjvIRGWCxh1nxb9ifPjHmH/+nX8s5jhU2k
hmySz6V5R8bx5Bohw/zH/wykuXE5yw2YLsH68dlYPa4b4/3PRxOGRYLIf4euOs2y
K20Uas6TWh1sYPFTHz0fAEiZ0N3BabiQErDBUPj+xCp4xF+uR7LgOXmYw+hsV7bN
H011McRj6cJbVXzq+a2AoHzkx+7ZAtBT8bToCTLmYcTPnm9Zp1jyzaYoptXct+Q2
9SMzaKafO1uu0HFWg/PW9zncVgoaI4MAlTsG2bqVQRgL2l1Eo13aLLLc8NtpmVM+
QNhH1U5G+z6ZiKnbOtPQet5YcwVzRRvsmdOr+vbZS3cmKV8uuRN1LM0H+bShuJmh
r09gNluzvO96E5vxZ3M982T6CP7eVk7vsP7zddwtzTjARGmok/HcOIt0z5aQzI4i
mc99S739V+t8myHhdwYXBk9O1kDcdFbi4+iCwFJG/YxCTa56wLlOmuEyWy3pCAlu
iFwGaY242UZ0pMKRyFN6QJBkDt7dVdCW66Lky8ymYCKLGDFVrBam2sZWLBg10gHH
b+2iVP0mWpmQjrE9cGpiwmFXUMA1FJbudqaQN1kRNsmg7cHKsBeHq58yXkcbjBcL
ZamK/oOkvzCLGv8xa7uVX7AxZBwrPa40TKLNgf4pVY46sAqooXbxkjKUHB7fsA67
341kfraxKrp0xkVpEEpqTtf8aNkNPUdobtqRifdNy6QTaZYvzqSszLu4uOeg6FAq
NCMcEqfk1+P02zSeheSuB7EIt+Ttat7DB1B10QK6+VrZOAtVSQyE8gcw3n4YudKg
nUOfaLW4J4Ty4towTvF//NJYVcVFSglcnmaQ2gf5cWrWCy05M5ELIFlxIzkfndFZ
4tORHBSpb2O4sLhXRu+Jkr3qJ1cW36piyCrAhRMihBmBktAN3eiSkUyvhyEvja7x
XhRVtBJxTtRK+os+862ZAyhACidu6MzQGJnQZj9mV1J7Tg0m55dJ26LwfAWygoJv
0G+c5XRzYt+/w9ims6avYRK6lBYCh7oFqC/ynWQVPX/x7RCH3dO3Azd+EEn1Rz3+
ifsTGjnX+kykAmGNE1KmxKKCXJlANgpdNEfB/5224KLoIzQQ6J/yJyq9FUIWXqhq
pTJE16rv7J77gAWJyYUeFbmRFs1pwt7ZzhjSFCrjF8s9J/S/hjPXp5KSWf1Jb/Nl
NVo3VLfZXSRDH5D3vLGUQT7n8GMNkKyZR1b7XMp8iPo=
`protect END_PROTECTED
