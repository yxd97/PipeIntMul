`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
On24MWQ+6aGBvNhQJq0oq+Xm34oi6fkKEI9qIADZD5l9X7quo4b9cGHK4ES/tDnH
os17nJiY+4L2QR+W6QQnC9rFOKohZTJvEymCEFcQw9fnnUALQ7nZ/VKY5caybqB+
kbK7hL5iM9YAUZVM+EkihcklbpuBNmA9dwNLWbQVoVceKl1SnV6Rs8tz7ho/tbXj
wMPVJcSpAygU1wxmMm/SwFy4CxppYSDRgmpx8x8M0cO2xXMlsFtm9SVykyyRE0EN
VPYYlR4zg8gSuGRn+vMaSg==
`protect END_PROTECTED
