`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqFca6BFD6Rc2sKd58+yoi/fvkvmlrYwpXvDZVvHoE5z1iyvSUNGovA1KkFXqiLK
jrRLU7mzctE+9OQGDdh1debUocYJ3M/cjTjweldWwlgCwCWBQ1B3GrKPhHLS4xTN
TF6oyLwTs0N2FzO5N/YU209RogcgvgVCdB4zos+zP1HZma1X8CHxT3jiWqkl6/LT
2kRmwCNzlyfj5G43qWXwRbhbxIuWKHFe/CrA1GjDyvKRnAwjcgrTvYvOzOrH+NGF
VaMsa3NqolEreLAFmwBtp22nw0Jt2wR6s725nNEsCuTF2jPHHqEojwaLdczBP70n
rdBZdKJYOPy403jp0+jSB28o5zoegHKuCJWQ/0CLV8V70UPK4NTsJVClEKNpIv6N
i1LRcD1RiGiYOMsFT3rk+WZkm6h3v3HeEmV7mpQ+JFKOf4NvDMoprW0vKFVUZdpd
piV4xOFMCP3yWq8vXECvEZsolZmJqf6YM48wAV8pL5mSFMvQN0ppYcybkZkfiNLJ
vWPOTsY2972RGGhxaEDiC5BmoVVA7w7qbFLw6zljW+aCwvm7QcNHpA4lFwtIfbLk
W5ITVkI7QIIWrYii/C+pjg==
`protect END_PROTECTED
