`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LspPokGeIZK5dNqf8iiwiSW2ICAPsGplgpZ2cDXMdA93PqbxNZSI1laVxiS5Zuka
aS0KAP0oEjc1cyIE+ldMukBM63J7sHflUjUv3/qvIJNx3AYjMHfe8xtiVBNPo6TW
GHlxARfhFatM1tO0xQKI+OK+iUWt01v/Af96O+alLw+3q6hDTPp0UsP2pxJnOOKM
tk76nM5Kc4AJRu046hixXDdlKUkUv+dXmvTmNig8ANLXBxEFLUXhZxyfpx7WVYiu
zNdWqQakMs2ptAO3Zm1phbinqQlDuJkTpY5HYYU9dmCBmKQGAS7745dIMvEQ8R0H
JUxemjnlZh5tlcokI2XRl9+D5NcCI1FoOtKGOKJAi3yKBpkKH8NOeq2UDW4O0QmR
ro+KIJvXfJv8Uyr81hSEz7yrbOqXM9+DuE6kgDHkhM2tGROxDbitBWfrCOTSnFMq
evWMtvnpcYn141Xw1XLqAOvSi+vXL7wRejMn2blkgHVGolMnjaQuAxeibyr3bz2w
QyM2HFqgMV+I7z0cvyesmClokiZ0rcB1V3uwUVREHp5huq+bGLj56cRIrponYAyJ
ErdXUiGPijgLXUlTWsWq8ihls0avWxP8PRAgPf/zfZnq4I4vD3zM976JWSh+1eRA
1l91oSUs24nyY/BcHXZ0EyCoUaTy0PC0yChCQL0KnptstgnoEZ9mmTpuT0DhEZSb
rB0pBw1qhXO2Orooxdn0u0PS/YOF5aS/PfGT/f9xpm9l6gDkAs6rJbGKEPAXcEhT
nAiIjoK+WzlNL0AO5nx85QBEURRKgpiBt8SYDHue+d6dx+joL+DzL8HE3fmHKffI
nRcWb8cEYwRNd9Y6Q5h8jWIH8FsiyFFEVLO/6IiXMY1ceP0Ucd9w28QNgluZHltg
PKjT7/NuGjuRTKE4daEwSbWKMaQua580gfGV6SLFT573Poz+vEf0YYIY5PlFPGqj
1YBq6vB2PGUdyzT67nTNFCtLYpT1a57osTXo9x5MzTilPqZy9KshtOqqq252V9zz
Kd7dpwITpscu1HIY/g6yT9P5AF0m6zkcH2bdGqKBv2uBzVcakydso5ovmbzB37Ui
I8v9TEP6FiPwiPkBGjKc9mRvTV2NFkM5z/h76cJb2GWQf5B4iBGisqo71ekF4DwU
Wh186kh63AV1C6XB2HQbO2q0IXH6ORejB5maUw4QpFPB3Kb52O40v1f47QXvEwRJ
`protect END_PROTECTED
