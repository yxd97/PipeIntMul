`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nLRV1kU+7cAFeNYaKrrXpqU4rPN5JrdzoCDZ5DLxyhUtJllw7yMJRc5uRXx1pLB0
v6/Y/QjxZYptFHV8awFhnWKvMDmZLKg4yVx7EOFyEUVv3u2+IE8lJLyy9H/u/iXe
VwE326ycAeaQrFslVB5n6zLxh4wQ/R97FnqAru+WbmyZZakTz/QFGsgEYckVl3RF
T4zTWToEv1T4BBwy3+5AWE/3XcwJuBKw9aZPb51YZJcm0D8jPnLOEBqaUIHUlcJp
5s4ghvDshXsu3Tlb36TKxdjcrnvLSbCW8yfbSYJCeDGDbpli3MPIYXyazuNlsZ+/
4Ic9ekGtkcAk1Lhd/muKVdG0qq8oxOBfcH7nz/LEeQ1V69NUK43g+jvLiEFo3osm
yiYqZzlaSr2+m3gtgMm1sUZD537ayYYIeMN1wg+39T60kUAgqc4x1qEFnCvDDf+n
pazgJDH6v1qScugrgTnp0TO8rrjZxUH6uMXGQ/pR4VyFqqBTuF6cMx058NPh70q8
AYuKH09MdWUsX/dCd6DR0i6BEdMXYRoBZPBIw6gdEHQ5oxPzDdy1szy2FusD9m9e
T79DakA9yOxqySpaVMv2vY8S+v0kRY3OdwXPk21D1BaHPnkvKnZ5xlfOG/1XJoH8
teHmPFFVOb/IOC4poUqwMw==
`protect END_PROTECTED
