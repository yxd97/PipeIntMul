`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xz/SgvSQdqiFHzx60tTUmRH8rSRyY3VUGEyVkv9vkY8WX3wdWqrVaahK9atQqLe
YQ2GWDxbDPUUFk61gwgYh1ozgHOhVpsE8iPLUs4KkD8+S/TcxCD1aK6OkxTgRhMQ
lY7z/QH5HC7oepGSI5Re8NgQRipaeXqpJFaoy6QOg+ej87Qq4/kYXGDoPFJNECCr
8Piruydge5ZuVGdecuqBjKsrZn6wkNbwvbWdGMxPt3Ye2newBmnyM9ecw0nQQ1z8
C6HXX18oWkArJXcA19oxUrIhsr/UNrfG2XfYdd1kDW3fdyNgt+vM38FTBNaPQSAs
b5zWcTzfiVXgB7gNjweanpwVH0Sk+yw2O/AsznwoYfA2PatIcfYBshbuptTiKwLB
VP/iOc18EoVTob8ycogpNpnEbwWUFUkktvO5ryvuuuwwywFzLJUJ8cfl1U9Mkyg9
bfRuuvG5yE280OGEkhrd1z/mCXOnKKxZZRZy40puLMnW6zWQBI4r6x98+YXmL0Pl
TX1ZDcgu5Lh0CrkTFvcr5dfLEhpvh6N0RUkkKS32xyNmWEq2fjl50ejijqgfpvfR
g1C/hCZkqgmvZi7e/WE5CeKF5AxLyYRlmLlKA6lbUs0=
`protect END_PROTECTED
