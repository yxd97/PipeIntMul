`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ktCHPrcdcu8fwcrQb/KyRB4JnVqqXE2Es7TbEsTS6rxbsaWZmBsiHEp5MB+T2zdf
dlQbR81L0DxaKEjhhHJ01WkTjFvHDHtKP5RnskZvJKnZoDvT5a6mdwBT0qUn8zSQ
pGlWe2A2w/2EPgDE7clcqmVldaQQTpcRwP9AGNUZyq1BRQX4Zr7b3flPV36b8wix
Oj9ePaGjPtJHGgSA9CT/62VQQe5nqOTv0a3GZAG+hjd3ZZw//OUivDt2JsjovGvE
Q2UobY/u+o2vYe72LgUuow==
`protect END_PROTECTED
