`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TN7zHwyanm1zcMWeUvy/xPlXyX8zBTKOwAwPPDJO0de0E+7YlzBG7gavbyDCWcmu
qZ5stVmxUl2NlRnIs75kbRJ7FMhm0rlxvixuLapYSx+tUvthivLdQc2kMT7vZDos
2lZ55KjaYk57bg4byIFtqM2dS/GlaObDLgpFKgqswCmWIZXZOMRPq/wLwJ/dTcTA
BlNypKY+UKxChM34dvq8RH5KOy8mfVlzjn7K3XdGFRYaF9uph25mH8WaZYBhL4GU
mbch056iBuosGzL2Uwchkfv16ELMaRsUkzmNEg5ZmY5LmqpwpmXi2xEt6nu77H9d
klaYXVZGepmqPlIR05SKoI8ayxclwdAZUMBQlozl/LUerA+2mZFs9Z8d9B96CNke
fYNN/kUm7sGobkMVT8C5OUXf3GuTTDwpcBYPudoWJfRALwoOZKYKSWXfmVRRArRt
JPWqq/bL5U2I9SZkCjCz5gTICj9dGgEp2qEWnUd4zACtWnJsPtwMI0mxu32CO5r4
RQwIi4GV/izFWFAKcZBP/NkXjyOWJb7+yU3vvdjQk1xN8hmSKJEuNIqOgaE7bYsX
S6KSBr2GZ9rxgSNoAd6Zi4cC0aG8Ddz9DbIxH7bstS3MMOujsKQeexMp6hHYXTK8
2tB09vsxAkFgsEHAgC3RKUGcWS7byXhmGuOa6feqYl9EcnJqH1HzTM4EzMQD1EXp
kIQLD7p5Huua6cx/3FZghI9BrvbMJAXUPn2vdz7VBQjW1G0aHD2RNam/dyrqKRlR
IMprz/YYnAGsYpJqu3nogBsAVI/jUOeONZsDTki+sxy+mGaitk426VD6i3pN/lVj
icZhwSfGkLT5Paij+cPFbXQstgrmfrTIdwn4canqrwbBcSsWc//alpqkDpA9YAAa
7FuVM6LKq/6vaQMwrE0D6tcHvcFW01zk8kcTo45jRjg+pcD9J20zgzQ2uxWKaHGu
vgTG5/KHUUdvJImClT5Dl8w09ddoiXjBqiBoryOi/LlUZQxkffSn2a7mAnmBi/uV
M9/rx3UsJfaJrPnYBXdZQncoBlY+U3yM5iRm04yZhA7wnfsY59jecaPHMRhnXMN8
N+gbSou+x8W6kUGQVb2TezQx6I4BydAJVJg343CBfYjZ1fyOUSOwYTTy7UPJLDiu
5+8OLor6bRtAjyYvF8VJvQ==
`protect END_PROTECTED
