`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dL3tCuSc62cOWeR4f0Fls03Q+ktGyLRAVPEFMkDahSTe/ZCXcH7tfjiGKKRnGTPD
M0TIfhXV+8ESz8WLNGuuAeYTmOn6YogLfuWkH00GXyJdO0oXwRlXK/m1dYW48ICl
ZaNs/UBchIkb8qSM7+nw1cQFziQiQKI42BVNzQLVLpBh9i9594MWHAaj30qzTpk9
hV8DMbdUagL+/zzWdFkIs6XJILBAR0g6B1HMXFndvZztmNbizm4yCDVi2+DHxcLl
wW6WGoYkhmBrJ/osS3w0W3rTvml2Q7ReJojnZKMETcwe7kmgTyEaP01FpS8QDxxf
TWiKbAHWv92gq+IdeD3qrLZd0WWwsE+ftf6doIGCCk+IlTh1Z/y/eyOjCkJMdSQT
rEf1BvC/69FWuyfw28EFZaz068PyGETxmRd7d0Mmi5VZcqGlEU5ZCA9bdZkjftEs
tm0PsfddfgPJWrDE+Afwoygiftr6G13y6StMggKFt6+e3TJ3D8jDQqB24BW+9tRY
Rkc1+TI+RamaEfeH7n1oSR8+RvosC3f55dqsF762aATBMP+tgs3+MfS/iltY7Fcg
BXrc7LntQ0NBfJkSo/0R+bXKg/kKf5vCte6CWTl4mk8=
`protect END_PROTECTED
