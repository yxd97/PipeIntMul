`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cY76pagswvmGwjP+kovCa0pMFwLOZWHhZycUuJwHkK95RvpwS0Pl1UhfneqSMDhS
coI4xE5fmVxMKn4qTJZuka17XXRNFEEMdiW1exbNIO03kclt72x2WDzsFg2dMiXc
jww0C7XnUP6JKwaFGcaeBFSgxqsWFg8fc6g5QaxeFd5WPr19zTsCBKtZidnhwn6a
+wrwgtJiuRMYfBG55bNPX0+IZpZ1+bNXuZlfgM6FJlECYlKMMBOcPDIFo1fee1CF
iXkK63ZKl3lPwP0hD8K8wbDcTIaogexeoUYe53fi6codG20Y6Rf1IWGj6uxd6Ndr
7lpnV9owdt31GZEYq4Ej7g==
`protect END_PROTECTED
