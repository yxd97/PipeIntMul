`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0khvOdf83s6eluskDnJq+lQgfA4IMQjwuakaS4smxZDrB/EPGbLGNMgswD2u83Ty
TnkSrS5AKf5IsVUFUy9K1IqL2dpk3E8I9vFuIHK3JpY5gCUIih+qivd5v9Taiy+P
dq4gVgQkt6Wc9tyGQEZKUXq1/OnoGAaz5VmhZAxZifHwsmlUscvuqKyy4KGHJDPA
UGzKBYwteBNiJBvml0O7/9SUvfliM7Agp8NsdjXdsbmmZZ48RtxT3LadfGm7tJzE
E5u65VSj/no6CFAkB0hXKwkK8/8dhLkX4fzPE68+/oz2hmTXOJKOz+f6zjU0sWMA
t8qJh5bSm6lFZy3tBdHxrBlglcNQUeyofylq1i4NiGwxHjsgyneV4MNt8+tkMpGc
oO5VEVf0L3U5URF6WZZGEzGSeoETW7+Io0bSuMUQE7PxnuiPZEplLtRpZZcl4xhX
1rSni69lrgPPOTgqPysKQqfle2ul6WXZ1KX9Jo6o0wHQpKxKH+eNaZeeR9/G7Ij2
kPF1jJJzbPCSVJXZjkd3KjEfqt5ehBoeAErM/6E1dYyB1y+I3uThTvKd4dAig9rv
LzkM9g7xCHRFxYBbmnksn27nt7sFkzAa3MHe1kyvGYa+SVhHcPPzTgQ6KKDokk+j
uN+0dDXByMxuvONQLaifHo8R96zKLDjymtyqwxFez3dqx4WwmqABmMdgl4cxc71d
ZqRDUzk2TOq2JwUq0Uxm8sNTcjyGmGVGM92kbRTTj4X/zuSlgLIhwrzX5ifcHSM8
doujh5tMhG/ohRQtrhItg+KNRP24QrJ3/eGKa65hQXVw7VT9y3rfVzAt/xL5Mqxh
4Xv6SuPTecKTcoxpvRgfdpjzDCDvCxQ/YqLAc0mEBa49tibL4gFBDQyUfCiv9Zcy
8CMS/ZK/TT1ewrQ5FsBTP12pmu9ufK3CSKQku1ipAi2xZze2hMMk/jx1Jo6Mb5v8
EaURXCHb0YTr2Kp1fE7aEpyYqg+pYK8vK3aAV/vtPibzV4in9udU5l4a/OqnSW9q
TRRbXXczOoXYGk1GfujphDNQBFEeUAt9w94bIL/E4tDelFjZ0cPpfXUNhXWQtgw2
Uqf6SZ4jAoqxSFqMAl+JRDzVhm/W91RGo8rBp8su/ge0TRbTuXhVxCOTNIQ+k5vu
5JLchgnt2bs7kGBNi7Cxq2Yi0+W6oM8WehOou6+M74c8Pb8IJgGOIK2Z6jtV+3An
2SEdK7u7PMWbEq1mijHF9KHsdGvFOQEyvv0KulwXOiHlliAzsVrXE4txRBGrNl+j
`protect END_PROTECTED
