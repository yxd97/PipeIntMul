`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evt4e++//BHwVBvfRYBlmh7Nyu/4DqEMz+TccZpfi3Jktn4TQc/JidySpVorIPhA
4Bddq+3WOI5ZCU2QhVZiWDIr0Zkl0mrT9TGK5MOiC59LSWg94+Oxxfg28CoL5Cbp
kS8oLQL126c9lzY4WoLGF+zDsvGyQWfzdgwc0BHeAXHLhKWg5r8VzkBoAi2aOTP4
htlNCwPdPn5m5iPqFBkhQolXTFEnM49SOtSYQ8blyof+Lc6AkYArdAgQy2S225Qm
k0JVqhnbtsw5iVF5FrlEEiGV2kQOM4Dc6Bw9yufLvJOXSbZlzQIAauBWP7UALA0t
DbnvhfyJ7WZQ7GDYlJEHgzfq8QVm9Gjs2l4MXEo+VpN2YQywzNMtPk3i4enfvIgt
9G0CysY/WzPySeoZtyYYEtQAKRDpUSHKqQZ/Jzddocij3XO8i6Ob8cgcj5wNB4oz
vExoHcHN8YSm2CclLy9Io49bPkpY2Kp6xgIxUgzW/EU=
`protect END_PROTECTED
