`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qykdo+TNWHCS+uuqC9bajAnaY9cJfsxpIWKhtNdC81m0XT/Q/Dd0muVVqgslIdIH
JyW8hEeOlw4rjBYFQhobTwZDd+dhJXzCeu5aO192W+K/o/Ed+p5xw3Xvkin6vAaU
QWem8dRLy+jBL6XH1LIByideGfeTM024fzI5W5SHV9CbLBGp7hv1oWhgC0ajwzsQ
+VgU6YyBVl4Gq6H8xM5cPQqwABpU+CGb7ybDKdPRcn8NExT0LNtVKoBoYISSEStq
584W14x7vrAFZF6X97TmNAYeQ4RI5ziIntwk1vQoQMVDd2MFsZj3yriFEhrSAGbr
fkW7uautLLuH19f/PA9rSYGzug4w73/t0GBHitq5s06pdXvs62DhtREY9iOF25mp
8YYosiOrQuevtj0KOHo3Xw==
`protect END_PROTECTED
