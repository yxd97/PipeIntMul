`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6c6LbyojEpOfNgA358V2uAXimF0SrzJiosgz1nEIc8xgvW1FOio07jMrxUIBRSt9
MNX8q+05BMvIACgrTQU8xwoBx45mWehrm2nkKznESUi4YuQ8EapASJfqLYAAzznx
c1LtOOi8NYjU0vTYd3DTiVT/13AwPrUrsgBUEVJ0TdkQ7qj+3wXMgMvrK4NkzkF0
lxOSbv/IGVWWYhBi03+YF1O0Igsc8ZpqqhGNnY1m19FpqKa/VoYyigdg/JhebGpg
KdoXGNikb++dv9WKMa1CHgpU51d1J0ImfiNQbZ4aX64iNwwNoSm/rHzEgP1s02Zx
qgXPNKWqGp3NOttqmzFYZuSfRKdWD4b+lPcPzyQaRfP21hP6CcT8ovKjP9le+hgz
IzMpKkp+7OtK/iVZ9c19B8PGaF+tLM94ARiN8UfnZtwM9jUW5xnlB/Mcfh4vDfD+
cTCdBmKXy+kXD5Mg1RIZ0bv1R8nUhaQfItoGV/3sDtK1ck/fUll992y3XSP9vpvm
T/bpNNTFgVCtlo8gsW17vyCe2sk/j3Q2X2gM3iJ3Hl4IW2fHW0h8CevVsHXjo8VL
S4PReA+UYpBkhkWs4KHI9ztQlkLC5jrY84Qo+j34XPhyC2jamL4M1fNrpp0IEEiA
1IKh+hlsnSO1uoZUR48T+5BBIopeR4mfDaDFK0x5NZiu/7vkGoY+UwmHJtEuXMKY
gcYlchIyaKLQF4S9TtZO+nSiLl1fvnhxEqtT6A/pIfZQJsjzNjs2W5j8JsLmzVXX
OYvy9NF9pnQLKCExCFprQyjWvmUkPYkleaZtwQKWMAaAXyhXfcphOSKuzK3Adstz
gk8SxzpkhpGZeM+KiSW922smHZu22JCUOfnU308I9gc=
`protect END_PROTECTED
