`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G1SztpYX5yVIZcigvyPtdn540l9Th6uzbH1uFl5uYAwtgsaF0Ntve7PVqnyyxs0I
T6IE4c+ZM51wTVHt5ZtHevyyQ5BcODNO+fRhsl1RmR0lLGUt1Cnk8Mx0+ARJ5XiT
xzc8h6oWqtQNvcJNhWAddm8SUehIcRL8vbgvRqHm9zmFEULIoo8Fsg53JgkvuT0b
JjsDyw3sg8PNaKltLjAmhNJkoQDdSU4V6bqPFNoTUkDfs8vTQeyJR5q9dvqFMhxI
n49LAfXEqlxD9gC3pACOrWb05ZmdGDqsqlCbEfj6ixTbtx73q9yFvANLklJkTREe
gJTkp/PqcHvYymBr/ld0dNRgdhfOU76FikG2K8t8y86dP/6PaR9luslVxMHKxcCw
J2478lFvfDpx7o/KVGmEVCFr7Dyt9LceYIdZ4mvvThLjVywDs033e7LlcihOeFpu
VMc7byWCgv5c5/qdfHZVHV1GA7BFNvfLQ6dduGy64SB00qR6t/ARWaRB0VBSgIdC
XZhjEaIcyB0gFXIBIJk7hzio8eCHGTQIawVDmSOfhMtlgoXLls258Vf8vSwpGKus
OOa7j8w5DUozwHQf7J3gIj6TIpLS8PaRvG0PJPEasx+nmQAmFvCYZVfmZLlPxwkX
gdzHbB4OTWoLo3IWP2WNIQ7V15ys6aUClSCF8Bzxuok5NwG6pZC4/JEi40+L6ef4
EEwXR/kV21LvIu4nU7Aa2KGDzs4SH5leL7/0cDhqJi3eaZqXRjXRDVxf4LQLkipH
Ipzub8BG9ddk+/T0+rLvVZBT19Idi28TvezomhcZ0v5fFOHGB32VDSazaNL44wz4
9j+Pz8uhuQrQCTqcgl5cuw+uL5lzx5KswJlk0i47LUGhmbqSPn+W0CtswbYlcy7l
zAfF/Yk5p+UW0HOpZEjK5P8Y/sNjBkBKL2xsDa22cNkdo0rOA9uKOhRTiI1zdMwb
LRbLQWXmQb0+lOHUyQgUrdCUBR229zlfPoHeFyyQbt2e73A+fblTT4dS+7gnP3Aj
TLk2VJCPSmV38Lh70XgSJpZFiAST+Gj/4OSz2Y9SM75nh9KetaUxivvwjHVVqduF
kfnXjsEeXNSpwUv/Qlfb2h2GXYbezRzlPE90Xo7MbuGKPsW2ztpr2uWoWRTFfC6h
wLthbI94bxeQezqyz4nGnYexcH+MGQQ6hCkjBM8l3r+9wxQ/tiOOIj7uCRoF0y+D
6zY8H2W2RZWs8DAuderiqLQNfzqmBmayMFls/ZISR+fQPkNt4OPAw5mQii8l9aNT
sFRa4/LHHaEev4wZPPAYBbfoPtd4gINO7ywQ2gqJyOgEkX70sSm/VST4FQMiNi2B
kj7WqIHEVSWe6N3Kmx08JESl4v095qUFtf5c2wVXLZjLKYjPrMzCNVBSyQsTdqnK
WwWLJRU3dooCBDZFyb3wYZXKBuNQvr8lRjy6tQyc4VqvgVCBZ/jo9R3A21d9ERxx
A2m6DjKiNP1eqkTzrvpaRj1cAa4p4lHGnPyWdRRoZAbz4aHRWm/uLZsNmq0rnmyy
bCAd9bYcM5llqdnVrQlF+jaXcdWLSM7jHjmA/Is9TA9NwEbdmTMGwdU1+OAhR5kj
71qj/TfUsKNM09l0m6+XfKd5XYlaLwesElUKvcN0/qbkJs/l2k1Q7oYsxx14/clu
mxrt/zw+GGSgmRX6vofrfrYBAJFQQc1kImrNM/W7ePMAtRmoSjIo45MnClWy3+FT
4gpqaHPrk3iC9T5bFvhP4xQENut8ys1VXPVdboScV/Ds9EL+kvJpgy67u5rGwpPt
WWL3qMd1iLCd/mYt0Ub+j49m1MO443W/2MmNd7gxGDkrka6aQTU1ucOnXeL6fpTO
h6c/vnLY3zbcpYp69G5CWzpagxbV8COkCwpwpXXGxwVgNXKzlmoJyus2kjQYRPfA
BE4pxslHiQz1fvechOK61j/AotwrrgzOg7d95UoL1BnYc1E4MzRTibCwuQQcGbFB
Balje92dXIGpSsMxKkKyLNDbssPbU7hUEH+OtQcgdE0XggnUXmiStRuOFQDQWpT0
g3pgXx3Bxn1mUdVgA4CIPDYnACjkth/l7eSbzZPIASMOdqlkRFptPPqGXmz51Rmd
Z4TQE1tSoX6Dj53/UMUIZwB9zDKtI403lFpjdNGq6MVgxFieB3vPi1bBsfUyCxPP
`protect END_PROTECTED
