`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/LounLuxuh12kBRzW81fMwRoYVQAXQyO9gJdTGvy8ddjsvpCvoVSN5n3Pf1WlC0
/FTiH72BuIQyo+d1donZ/XcLCHM04eanIfCB7FVc4YJ/7n18gqtprnoal9v5Siy2
mf6Q70i1VnfYYay4i4HI5spCpqKtXDD6p/7lLDg6rDyTr+QmLIV1ocwTyF8QtjvY
kPsv+21mDFtGeMkpi04mqZq9CiUoD7E4B+zJqX4eW3BpY/CahcPr7i5NEgwH3UEm
A5jVbviZ+9VSPX83uutnh0iqzF6ehXNkYDJ8Z3sR+PSvgvd7bDl12ljCuJ6nSxL0
3ABOu9wyjpU1b4QyRsSKnTZM6KdIDRng2AyRyXyT3vJo75t4tMkvcOZ3IH7K6Tt8
rexF79KINHsog9eJ4v5kISlnPIlcn9ELDmMLtN7MdN8idwYAibW9IVaaGN1/rVTc
smjfVikfWzrphVXv3lVWMcTHmbhf8WUrSci1OUH8XhOqgGWIThvTiTGGsXVX8COc
`protect END_PROTECTED
