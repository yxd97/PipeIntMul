`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QS7ZNomJMl/R2iXDGpFOfc3Imk+4CcEbI9jZUE1r78s2Nakdo6XZd5dOCDlHud6X
Aiav8E28PXIlOLukm9TSLLWCWlxAlcyXTuUl8DM9eV9ofXV9a/2baLTN7a/DCS7U
p4CKwnqDECuDuyAmDPZdM4j+EEUccxdzqM3S5BGe62KC88/r0/kj49UcYMH+M2Lq
/lNSrv9JCxlLXfDwiGzA7dpKrktmoPDqLUeFmogElHjggJ51noOSW76cLSJytR0x
VI778J06JaATObt0KRuOQ1HohkX27zHEhCH0qh8GUc31qhpfjm4ceyf851V1cTWQ
ToKvmLq1oYu78t1mRp4ysfx3HSLPWwNNYHGZQBCJh99ntVCiYhRL9V3ls8rw/adO
LzrsJTHZkST/rNVlvbN7zMEJvwAlyGUVIYA78D8hKcRCTOIRMilaIwUHIPmIe5PP
giF5WABQJZxAdGO7DB8Ezh7MI4XICj+ZDtt+6xrrS/PZsl0dctRg9M7eN4MVGi5K
rin5jti07UCLYRz6mjtA1dOZ+qBueGlnaWl/jEeCrBQ=
`protect END_PROTECTED
