`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LREZMrtmB5NotDiBSEdlmE5Gz0iAygVfyFP56LA49G+QuBVvbnjKILoxzQUpsLXL
CgcqfF90DFWltoS1c5k31R/VaWJoxCPG0gTzhS+BSmX/AQ8m7TxWlECCqm9E9ON5
xqjE0OKRgI4C6y2QXm3oCk7lLvTQeijcGRD0QZk83RPonvQsse807KUs+1yGBk3T
Jf3ukjLJp56qM97YhoCK7jom9PNtfOTRPYdpAnbTYF6LC8G5sPKesX8qzcEV4FL4
NqrOZAjW0TpjjfnOxs423L8lj0mW7QWEZ4gEE3pc3QuNpI5tUHjdr69KQKGwHZXH
9EOh5+5LO5isqSjJ43GlFWj9pLHoR+WPwOLoiTJ4FJ1aLS/6afSbJrXBJGRKdHip
JuVSDBa6U6qZ8I8VMI1S357/Sib4XI48fq9Jp8lKF04=
`protect END_PROTECTED
