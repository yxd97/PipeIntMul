`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEj5K4cspqbTWbOunCZcZP9VluAuMpIYbx24I8/l2zih76K0vTDDiILgTJfSz5Mp
aRwosMa5hyE9Z5lLeyqDVRIPnKj4jkM+qqzHoqO14wL2In+MkFjKn2Lbw1a6aV00
2pxhd3XD6s0nCyWCirQG0+CXIiDXVz80AdUo1kTKOnUGxfr2Udy7o3bdVvmuA7jP
19L5gzKmsILvuHD0EN32Qnq7y3zQZ6zTX3M05QUgR+edn91i5LN45EeLiS1HLZmu
nITuIpTDTS3nRoUnX4UimgBbHn+fzZ4zf287DGQ4QW1K2zz0s3XfUjyRaG2Y2EtR
adPNhY1jWDNqCXjuh+L764K4qxorzO8xv3v7clef2eLZbZ0dn69mkH2OSojFhghW
HrkM19+qwoHsxU5/cJLO5Ve0Hyvbpx5+Dr3RSF681RvNx6w195k7vkwAE5dbOUvW
0lsW6yDcyoiQbTjxHuChEG57VDviLDP6nUIvGyav5+G7EI/RfqcVLzpj/N1PK9Mc
BIi4hEMvjiZAN5ebSqrJS3jLoAC5czzwG8p1z2hXhy8R+u5f3MIkNwAMfV1YfqRK
SrQ87+PPcrYpIyrIoGpV//0zktRUkUch05c9tn2XQugwt4wyVRl83k4Jvurna3Gk
LB3ESj9kchP6Aj28EvBvsVmS9yuHvMOBrigc6nkfMwXvmBo+ORR7AvvBJ9PmTCnm
oK7zg1tHByA4h2abqg/TtPiUDVNmcIZ51ySwxb4SWrafdA1ic9KqxPVIPirNA6KQ
Z+XdZjKf3Gh0n8Mfbar3NMLWkZ2I52VciXsksGgWJrZXH1E1dmltsdhRsm6KlhhS
fOcbnrEE9YTbvpoJS+A2nsdY5LUw/QEmZ1DJ6pjld3pWGuPIvOVA+x6ZtFRfBmhb
AfbLMdh8g9jl29XD0mvFeJNLsdoyDackB1EBqRkmsuXEevceOvOF/I5sIsb86ZgG
cf0oZGem+kEHAACfL+gAODXr1ehcu5cNU4FtmH8ey9r0uEbsO7dY8HtmniTrHcXX
4htOG4jscEu9NuoIl8qwmMGFOBsQYmcNsc1aoAcXIRoQYNy61k2gmNQhRdWIdhpp
lEbhDnLVxx+qw3c8obg23iMZYRDTQ2npHNEFiMP6ABS3q1eZgOdX9fggN7ZHvoS7
5+K3rjPyir+RxUUmJNMoX7LZX59uV5ZxuiB9s4UgjZxakpR9ZqJtz7rTWNSkdSKk
I/YGLydx9YO0DPdgQI3MHWI4PC125+wqm5VH5oDcTj324cixs0YABApyDuXBg7pP
VgJZkE6Stz7DicWF8zdBtdHkqzzJMesD3foL2IT+lPobvwbo0mkS3xnB9HrIkn4S
5Jf6bv/BtJjER0hjTxVnKGZy8tvlUFLDm3g1pyYv0zYjri44JFflry9eTBsJrUE0
ZwFsA1vjglMjziYu5A3vUCs4C6flp9Rm6KA8JfWYp0FaJedrnvzJ0BElV8e7Uqj1
zKL6dLTBni1dyIYezNngV6aDUEr1qFzRUq48oz4BfC6FdxPZst3mz9DRXCpBJbFM
VS46c2LFLhigfVceAGbVBeGmh/r/ZjBf4Lr98Tuxx6px3tu3HrfWAbmY4Nc7Z03/
2Q0/7EhnyqIbv6caOKB/Z1TsgdcC7t8ZJWD7CnjxnydAReZnY57kbZt9+svooEkf
wr10i8wZ36lAM09RvtTYl7Wr2zErdmucHhfk1h3LFbZzrhypF5H97YalbqoOFRn1
7XGutlA5vOGfujMBxTrPK0mGm0w1EAfO1z+j0p8DJ4Ur/PcY06ay5F1D3XuRmYUB
6kgcf2HSN8nxdV0o2zfH5UiUz2HRotNmkZzfrMlnRj9fcu5ZwjvkyM/ZAWH9883X
xUZ0eKeaQKesE1AiDzbaccY882r0dLTqtcAjPyBP+cpJ4uMzz4HGC3QlzL6t3+y8
`protect END_PROTECTED
