`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KI/a0Xe45PO9vykWSRzjLo2F/QRUNZtD3+amiz72/FtQV90h4XsG/6vwHQPu5ZTj
M/mjcFgMU4l8IEApi1hBGNTVmrbQKr4NOAET2RgMWzwqXbcc9YW/OfxZdRKmiAxJ
nu9jXCCBgJmeINjuDS79EP7QdCC8xbGDMkea6lCJEv/1qbH7FA4dxw5tzQ69PaEr
se5f3Pxu5J7HTgO5ugd2mk+HduWYdjwrrgiJTHeKYAM0Qel7LrXNDFgvP6Mtzv5s
Mt+xr2WiUt6Aiwsg6eJzON7WEKANiE3qr+qkNvCGmo6NVjesx2iJe/ufZ5neHZp2
uJ1KqaHcQ8PF4PKboTlwVgmdnzoYvhmephWK/qznbIiaEBxlPpznr2FinXMseqPC
9ocOn/Y5Ikak05GmrjDyTLbZqhPlkf82od7jCMPmq2dhCaYqClPmeJhtoGK6x1zL
o5w9M8Pdg5SQnQ1dF24AJamVwhcl0EbmULYzjR4+tnnKYZ0GVHhgkeHRrXdvUAhn
v03wVR1Zx22umjZBjTMPmDktvfh9LculxgT5yaVLfsTNid5dM0C+GYKLacyVk9dN
`protect END_PROTECTED
