`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VBo6Gv35x/BFih1tbOlbiUxuoksPXgYsmwV1i2ifA9U3kZVeL/wMtArRPFsgVuFj
cFqGH1JxYN1rteq3X7HiReB6TFkMsHAnXc64qL0UgN1+fbx0zOKIq9M5nuN6p/sd
23kzDDiyjv9bZ1Ohp41xxqcazNFllD7SCWc1SnVZxrPhpVwDG9HTY6omkY049hA7
IgByqOWYd6XmS0H5HPGiYzBTxDm1XPcVmDDs3xp2DPiXmrNF2jrewyrjbofx3HPy
QXjEvZh6zS0b5OeRVUUBtcxLFb27wmREN7yKFp4PXsr1uFYG8jqb1jTaZQvrf2iV
1ejSi8zcXxQy5fZdJSUHtCEjEO2bYrOwJeTTi2Ds0pLUF+yA0eyyslMcMTg6eK1B
pGzEEkgiKd3sCnEQKTxtu9XWpCzFnQyX9BNgL/n78W4=
`protect END_PROTECTED
