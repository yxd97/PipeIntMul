`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yMrcAiaJxJAqfv3cAUB/FHeKO2zxDcRDRh33+G4EIdLvYelsHRwDcI2vCSe5dzz1
VrYQkaIHfWlwO3gNskwn4Sg9l2L9ctYXgnuvSaAvE7Py5zecDBSp41SpBXbgyxcN
+FdLk3XGo81tMx/sgDzw70LrHK4TPqH0Rcv5eXNAlmJqOXvwz+oNjZPcpctfg47T
5DInNT9A0JoBaih3zn9raegOni71npLqs48g9uOrjykssyYs7LjFcYzIMTx1SMfU
eteN+8OtkPDIM0cbRoxqdpDAN+xc1HBH1k0Tf/PivrQEKNNdaBdUEE2KIu0F2LsP
sQw1UWBn7KHANquSBC8hqe1Mc1bm/4rSIIljt48MYCs5t4btYLylVjPYbbeQTKre
WPaSN3Zz76l4dmM8FK1XNKJb9d9eRv0lwvPzoBpOtFsxcjz1Xq2tPZe14ASO3UZs
OHRu3se17IT631YntrnpEhciWcm4GA7byXWPDug7Tz4FeJWrj2fxC8kAuqmVYrju
fXCVEJjWigJ0Zb2VX1IRYG+c7kevUO0oStjykqlKVSnEZSWTbafwER2m4mviCBVy
TyZ7s7MU875Le7MzZ+BGlRioKVKu8Q9uc2w+VlaNkt+bRt8YavFzjTqdiaTBPio4
Jmk5MVuuRNnMoDXe9q2Mwra+lx0un5V+9ubt18JOjxiRVW9dbVPr23+BARydjKcZ
fJZnVg9qy3RD9TY7QcgyEwwDMy6A2l/hNAPcj2wiBS+yowz8zZkbm8EyXTMH0jFr
kgBgrnwqmE7rCDLBaWHcIhm5pFYoAxJbxfV4A2w8N59kyW/X1VoHJtcLWweh/2QH
Cc1hvrnH/Ha2MKnIACR2shKxpRGY2VH5LWojUSmtbc/N/gHlSFsRGCviJw+mbKzX
2ueHdOBuoDoExQcczRNjNaXL3E7CTYTbo4hqDdEMVThHperHPZpm8rYU+p+w4if4
ejp8KtlPkQKxr2mIJ7zvTPuDTWqwKvRNSoPl0F457+wMMHtEbG+iMluIa6hI691A
4m3utmYq9dMXthED50KZ0VyWfoEoM4b7M+BEdqRosgml8IUEKdb0g8NCfgEc9pGa
V1ggFGzh/fE7DDRLpBwdDCtDUw9OTcGF2mMmVC8rr65WsmdJHX/6ugKaSZXij8i5
JyxnXX9Oj63kFQbSfbycB5fxny+CShOmVH7niF7osqXz2UHVpUeHa2jIHcu6Za/C
xqC6p9zur8kdSd/m/bMjnYPYNgE94yMRjJ6m8Tqjmn/xZZPPgoMiUUZf1x8Sz+v9
R84TKkjhfxcEDcI20OYiX/xGovkysSJt8ka/DH9jSvKa9G4A0kUcrQMEv1/6cGD1
mQFYDYiuVrVG2zYVjWVSkwBjUt+v3MTMsKVcSLydt4huts8QHbauIprchal99J8/
rmGsuqTfe7ODyhNao66XLOn9uB32H4/jWnmyeAvChQUAr8Rsvd5TEIJavD7G1RPk
2B7jnd67TUD9F0v7DPV2pusUsQLToM7OsjdMov93Rx53sehI6xkVLr0E8VifYh15
moBDgpa1rBc/kJonayJMVPWhopQnhlNNTFUoTgUuLQizX9+pNnemVft5wIF7dcIv
gM3QAt9eCjI/XCxRf9vuWL63BuvF+Cla1+X5+3nL5sjKFr9H3e5MsNCFcu1FIEMa
R/N/e/Sx0FxgSK+ECAcb4iMU8sfZITKKpq1VsrnCcwOMW7pSYLzouR7mLIfaY3xj
alNHgRfANQhIeLu7AWvUot+O1kpLr7nofAb/wY16VYCHsk+Zhp46WUFhxyjXAgyg
YumkY/bzeL79X3wfEuIKQ/NKYiuHpcCM4UBqD59oaFK4UL6RdcmVOgoeFBwzhVK+
rIhl4bFAfjV4W3LvBNBAIDUgpdZ90XpS/I44zHWAJGDHB1Wc6pO8QfokKbhsTOPl
eKiRoCLyTpH8Bn84G6sQYslDfJzMOmNniWTxsZueMOyABZhec9tTQo1UQPeXod5z
mE7ojJmw0p5SxDrVvSnXd7xOzMaAR/BJd/UJoJQPkEWBmgnqitRyW0UGWYbU6oB1
NFisKCSCXdk2dzTZtq4tE9EStcybXWz/dDaJg3tsuBfR9AIWhYoQbftIzEw/+aGX
H/6DrYC8pToddJAabr6FDJQF8px8JqNAE37ZWClZyBXe1nTOkyavRHLefRP4G67z
saQhuAZkE/ZXcN703aPxa0n7SNu/05XMDJFEb7g58iD5PlI89rLqR/hMD0vZVVoO
aIyAfUvsunf/T+SHLO1u2+6fy0o6VqEHu6DO06BvHjP3kLqIjl+0Ty8RdIpQ1xZf
bwZbjlg8G1AOwJzTqLy+wMpzC8NZI8UkCNdn0ImuwJLH1/pX+1GGpKrdCPU66r8i
xFdVBQASeU+pW0UVoC2oIUh1UczL8DyRdg+8I4xQRQxww+0VSsMHIE/UsH9OYdsP
zXrBsqkF7USKowVFlOvqpEwM3+G1kcMoFC6mPJZ4TlXMcwOdyDaYSnxqD/0N4+93
MG5CCMJPF4tWjeopyPXyjEdqfODNu+tttnRi+Bz7o7cdIxSo0mKZU5FqUodVIe0B
QrW9JfvCYtrck27fWzuN5/SpK2tVwza01fw5DhGtquTFe9G2eEfG0ijLvCXpktUl
3eJOepsv3Q8LuiE53W74BVpNk3mPUrPyfEi6m2SY0zVhhCiEZe/VXnwSz39MVAZv
vXEIWMMQu70N78oWX1pYe3zEUqZjhS0H9gDo+XIFwWOht3XrMqAXqsC2KBAOzxZK
9OTc65goFM45zIPgDYdHk1OsYolrAx0qsxU3Tdki/JuGAJzO48fq0ULB3mZP5Ng+
JUAAyJvQdIdadJxLFEvLnqcZ72LkCB8vvV5V3MiQU2L5upSnXO5LKWQGFnluHOHY
xuMZ1jk53AVwCSzc+luscskNh0ZpDR1F2LUoXAztLw/ls12iuxSxz/irhu3mG3VK
aLRWPn9WN0YstiKmJuNFdWT5zBYCpkxnSu16vb2FehOteuvz4tR+MoqZBNA8GaY7
ZciA8mvozChkaV8GQRX496UdXaWhCEbsn85pF2M9J/0oKv9qa99IplA/WStxelH8
WXc43iakYfk1BQtpkAY1l6i3CnmTY1lU8bfPLAXdX2CB4MEjtn+UwHHQfEmuuWbC
By+1QOt0y3jUqDHlObwt1cj5vfolMtmBcwTfciYk1hWpuk1TSEuPPy4EfhT7fEL+
YhI8Ttx21wy97rMHOZd3C5A6yXACxg72Ul7IVGCdRXqTgiIXmxrzErjoA+aeoTlY
ncVkEOiF2Z+nFNUFTdw9NRz/Xq2OOjqanaz6mtErJ/5nOmi42ytpxW24CsX5NTw6
nIsEWsPimoIxMS99np6ril4UqzbdM+dMHJJriTv+Q/noQnDuhcwlXfL5mcVtmK47
aSC7YxcYZzpylE17GiQ6yX3zvXszImI4VSzu3Ny4Fyegaf7Q3A/43H7y6Pin07og
/HTIdJ62QM3bbKPWdL604qcCjSj1prx8Jw4zNfbDlJtAgTaggo/XF5+W/AQKfL2x
QApYlQTP6qK28/zRKfxxkHGBetuaVpLGEcrrD2pqbKAsDFrcD+jWahjKrwqqwczx
ZI57QEc4bGnblIENwCwJFCeVKOWXNuec/x3idiNXI+WpLIcxevG8407PDLY/gSYf
AjdgxW7Io/SmNJfJpE2eiwMLGS3dNnGz9wP2EwZOzIM4pQkOparQIhzweAoLJYRP
IbWs1N6LsOOXESP1Gh+h2nCVl9Ij72ULTLsM00m0HrKpZc4efHGIUf3L2R6dYwbl
eN3fE/I5MQ62QWeuETC9AyQQQ8DKciYzLsGbf+DK3jkshChcKIqXUEznr9fJ9Gui
8oX22OJVtXPeQmYAmYjRFvRBlfVQoJNesE/6nMAxhR/gpwp4qjEN35MFOJgVm0TQ
NqVDtQeyTeKaz7d5y0Q0nRR5si2atZT12rMQOCBPJ37kelyDG3MU3RqBXPAFsXAW
GuV0GtPYSYko3va4n4ZJkaPfdsQW7/pC4s8XdyZFeBZjvRH3M6PIx12Y5wA15wJp
wQt6vDWKM7uaDJ3nj63OQ6ovmE8AWbaWMLpS5bopY/LnXPUJojyvAhdXP+W2sQ37
`protect END_PROTECTED
