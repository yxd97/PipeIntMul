`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jH133mIavBzM6Sugmgt4YiT5HdDP80ax7sKjDCwr7/Qn9AQ7daHvbpwPkHBG28L6
vbzoN3NudtRSri9xR2xRomn7SZD5fFTb5oWYecNzmJ9Goxr304gfHWL9iRLwAf2m
QDYrBRBc5qSta8YrxYQ/El1H8K1Y+rFbIFpUE/gdrSuD5as5pwO+Wb0O85ZaMlTc
Zg73+r4FpG8SUwqDBSZi3lQHGV7b80cZPEutPCi8Ct8isA1C/hW2ZHk5PLOJ4+g9
KdsI7dSAsfnFENFSLDkaB/drbHdoHiauXJdbR5fr3SC2Oq9Rkq8BC6/P/zoC/QIa
Dr/cAkNDJwEG2KgaLl21XSkR9nEZMxgi1ba35FQEHoDtDOSGK5iwDXpZ/4NlmpLG
V9YEgFM81qGZiWo0Mvl1VCUhFeaKi68bi3/Wsru8UrDMNfLwYrfFn7qzSqfRVBO9
EIfQt9Ncqfd/ta1y+CoSK88r8gfSwf/VR7M+CnKCsdJnztR4aqyNo7Zcm2FVFVMy
fGMCa0wcUFBlzQYOfFpsWYfuvfV3dn5biwo92JHKkq/ZCAOUdtPqqLDoGg5WqOXC
nGbrnmbxaKb2d8lzptwK/7FIo4OyXXnqgwwSw34DC+EutEzrXyzNUUyJMOdiErmi
0NDo48Cl6SPjOTPS3NnFVxqFa8kxF+I/aOlxc3+F89B1d4n1oMFBxsfFxA5N+f6s
l8W4qSvN/WJ7X9kwwMtenzrkHvwJvjqyWH6jdQ3zlJ8m8zoQsX4yTF+FHM2+0NG5
ZKLlMvPfGgaidQaRrO/PmE/bggd3Sr0IBhUAsNryxFN6WoDpWmUOFf6Z70bAD2NR
faA2OnPviA0vaWzajqBqceaymKvi3GB/ZIr+bFRfeqRjv/gpMR2GO0pDygLzqdls
T8T6jB9J4N+Ph8n14RXf1u1Jisk0EniRlHVxFb8CS86ZHRXmGLiM7r8dRxRkePYK
CLYql8xcNSCJ3QeTmdMKV05ST+Lh+nBui5K+5d72KkrZKgs2PVyBsk0J26NHxs49
BySocjNfjeEQsmDau/Tg2qcwauGoGi6k3h90RTOjVuFAIwilpkGh4J0PnbiC+w9U
u/W5qhZ4xfJb5t2kc/9QD+3gCietU323TmnMxPrNVbKJgPQF/0PZdr/owawAYlqw
Psaa5OtGAr9D5EDyV1CnarCiumfxxxPKJaMX2bsHgQ4NK4oCzXAAQ+1idyzDWuYq
VXF8fS4VOPxA9bmurXGgtw==
`protect END_PROTECTED
