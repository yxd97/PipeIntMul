`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XF3b+Wamke7Ew47avZEHzLmEx+88Yfy4LTDUpfursbiJk/I7Fscjm4emk0w23M7
t+A5Lw0Tu01nPDzLmoDwkiCvhpbQ1JQMPGQ0ls7AWW6otdv5ycj5C8cEH05NrsWF
sgAMlA2glUA/w4tT6GygZS1utkUU9xzhIw79SODSvYPMbJ25384xpro33WS50aqj
ZIipO8NTf237hZkPg3nAb8IWus7/yAimJ7KmQzPDzdZ+HueeX+86DDdKypXHQPyd
Uzk+BLOvRP8dfq++g6gnLA0NYgWq7Bz7NqHk8tLR+q6hPV/qCzv7ns8wfsW3VnId
vOP/VfZOLjoOTH8PVY/yQ3kD/NJIyXfcoIY0pGqwguWFCKHynlGTU3pbpNWMjAlc
pJMGHGL4NYa4ts/iLSfLc8+gKyeHN4cTj3ylz9sfAAEH/QIKe+6BwBZYM/ROx2cP
zvZRAMQSnekPdVker8jxZOvV9JztvEBzz4AtLkmwvDDK6tpihKlib+UOV4tcfCPz
`protect END_PROTECTED
