`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b3EfnWXregLDbIx8hmmlUBL8DgTVvedQhFid6Y/Q0+0pA2wOgiSrqCIUgcWo9fih
WOGN9bEUItmnzYka6dKJZOH05UXjE7YWU7mbBqFmYyeH+rUpRR+6It2sE9GN+mJH
UvDbOLFB7pH4NqDvkQsHwdnQtxEswsOge6ppFYXVqJENFC2FKdlTzUuh+Swg5fJS
0L4FE9jdZCai6hKtuAmA4fI0QFT9PSLhXFF0wyjvUxECrbkoqkt2E46PjnO94J7N
YJcaF+eS5ghKaMFW4TO6hg==
`protect END_PROTECTED
