`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KpCAdrAC8DetZDU0wKD8W/w9f05gFAyhUvsmN5tybfdH+4Rf4aY5oGXh9fGOqxYK
jWUHk1tkRsXvtvEmnCMIxUEwc6vl4VANYAaBskFs84nandvqDmSI9BFuk7Cbn/I9
XVN3F/HpowNmAsIINDm63h3NMbjxF4qfbxkaSUg254ZCu/Z+PglgJPAPeFG3Lj+7
MVhkY6azGBUCjAweF3Lov1Zvu8l1hgvYPFZ9fc7QHg9X1ycZ4/YUNi5KhiP4TYLY
PksEYsvdF0hGV0B7+MG9Swa/+6bxbICdppVBw63vwOsh4d+f0LFL6ncFw8uKXWHh
dGI+BSYpfPxp46kTrx2aW6UNP9HJExzgk5+x1x1Mw8OJgxxSRDxJgG6ealzuxhDQ
M1CQGV0piMaYfG3UZfb4VGtxgvddLeqMHNJrYKSlcfb8SZarDK+UMKo4darYN9XZ
veULZ5J4UbDnOzopy/h8AIJFNZMV0Ayd7bVNW6WSx26PoKa5dGfP6uZS2KSky2UK
rL7LwMIdxFApEkbjo48Yj9pp4NCeKMrL599rDBrmOUYnoM/IXOcwFO5AGmw5eWoW
qQgfabCVTSupmVTC15laQGC1b6vdkunrzgR68OjbzDjwE+DN6gjIV9W1nc3QR94n
+KN9Fst8GnfSU+hgjzLQcNjwc4V1ZJh8aN+rgHzUHC4fNNh7A1zE9NruTwwJHXVp
qdxgmxP5P3M9oeewuMTlkw==
`protect END_PROTECTED
