`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9qnOvDYVM21SPQ/UUvN2ByZTVftviNgXIDfkPp4UZLxx9Fwqyy1+n+vjthkaakjO
mcY52OlqTIrbW2Eg1392AgSa85NpPKiwP+CraWwLochvE9YJ6ol2ceE8OUniuqv4
SDjmehqIicrYUBH0AhVyngDvXLtSsJwM1jvlKnkR4XFWx0HtEBHH8fJoyaEqoYCl
s2DUyu/3fM+8SdG5JkzhfJSg1UjHL+1MQqQnJuFxP13P7lNdWl897GWt7HrQ18FN
5NScByBBTlA1/mu6D2T44ZPIHBKqWlx1AlfiBJaFeUPXXOsPzKh94gYzKDJLlw6B
J6gT7r9ykw/UCA7wn5+F7BTiI2ybcYBY8WRmb3/MOD3E4JXwjjWNsVhJPbEbvBXe
g4ACiQE7rLtv1eVwCwUaH/2L4F3T0hqnj3OigJeM/1aX4uV4GkUiqBg9Aba7jDq3
l/M3FKFjCLRT0RycKciDf8FpZDnertUFHXCsSZ3sZtww2+9TJPS0nV0GRS6Qfqq7
4axvcoeXwGMPoPCw+2itdatDzYSNvDNCLQqOL/pEuE6KRxt34ckgcoWtaEw62M3U
EfOaQkCSwrBT/t03grF77/MWLkWnkRrZN7RbBp6IDgQaaxDUFv/UUH0+kp6L9siK
PwNWvEZwsRiDWZz0kULvSrI7j3WQL+gj6hPaTI2nEUVkdYOt+g0SnrJ9FqCzrsMA
v0WgdnGf4q918sNe1eLXzWZ6esSLQvJNaFJv+Wgrel1V+cV+MEv4ffGrqiNrapve
eeobVTtNMZwZI5fHaUu9jeFzcnY/gq+c0qY5LYxXszjb+MaVmaGnSUsS7GpI4RPG
SowW7nmKgpZA9aD+zSAjmbicDqVUTHWQVioN9II7FDgz5sSAJjgmj0c5Y4uOAIl0
+B/rFxYnU64vPx/sSR/150VdoNYuaP/vYiT9808PCedGTXcVWXK/Dcp4mHxPPhKg
PFd0hidOCIJ0tvkcZLgH1wybtGCcbWhfcVMMlzyzTKFKYt1ukGJMI4xWAKm+NHH6
Rp5qb0/tH3LwxRftMslLA7vg1Hn7yoEMyml5hi5D0gwtIeY1MxiaZfnyPKl6vVbq
PUOBhCSdd3zSjMtqg2BniTLuwK/G/w7lUTBGCOMJQdmRnDDVuVJ4szXLx8yINzlI
Bo+dq+OVqe1u8z6XK0MTu96lqQwLI/9M96iawaCs2hmnP3a7xvhDP9EqhLRRM+o/
9FDBqaBV8lOOTo0jGFfOUUj3nTxTvSjOPVKOfv2OLGdCsJD9wBrKGoKIlGAQcKtu
sJl1PvvLfnHEGk6jzJdeQZlGsUNPUmrSLoEnDZ4bfSzcKFiTL0hJFypH+78xZUHr
R17wwtrD4QiTpUTaFKE8NVEt13UVyE+wCva4mczZLLfZtIydVv2sN9bS7PXNlPUu
RJe9xHBNfQ2E1NZ6Fv6bpk/Rlk56waTvMo5Syyx2OIyw+ntH7Ivfzmx1HDeoFKh/
n40Euq1oeysvDplWQ0qChvyERBPxbBcdg6fs9ZzXv4U621uMIotBbCr6wt5kGibh
dVgG/WmNl5pT+B6aysaMcH2emrjEMq6V4+u2RmwVU5EHoUNNnshC1UaoJZ1zGm8G
InMjmLTDBHx30UKmc6mFQ5yUwHLAWIO4PGL14OpCCG/7Dz+++/FS64AenS5BoJtR
7BPBO2esmfWzAS77XvUSYfCet0X82qoX1NrXFdJe0yGGgTjkiCe+REyN2hc2TVTh
vhx6k2YxAvt5nFC/3gdr4Vkbo519S0BN3PkMKkCOxjmbm2xR5/BXaWbcN4CiZ2KR
u4qMI8mO5WR9HEQ8XvGTKW8IDaxI13fhmgiBa6KJOWtOC+JSc+bXkzG6NHB9eLqa
SJ65bRTmFxL2H/2O2NvcqHy83L8VynL67gB2uDPlIYYmgC86ek+h+7dXdvx6MAeq
c/MvROk/AeFJyl+U6aZRP073TDbrA2jQTMDumZB8wPYD/5kVaHGSh9ozadGQKuJb
lmvLva0ejmA6c7CP3FRpkszooo1h4nolWN6D9yXd1KgLkLD/K5lwhpmA9CaZ1Trk
rLLfQ3GXJVyytvNRlA2B9blKzd2EeP/sGHjGD4yZuGl6A7iFDHEXCfz3XwC1rVcs
R+SZNcRN4Eu9i83W/UeZXn/BxYNsiiqAaojP04Ko8A1PoIbgf2zO6A7Yr4JBV5fK
J58k7+rmtIwkJ1mbGCTSiCU9gpMAMwNiuKbIFpQv90cjScLuYb1fwa6vDcwqtFgr
ksKWSNciiu990cYG2+l2eqaOkLxMvY5EUK7CH6Gsi90TFRQPfQLOj9Dv8lZ8WsO0
bYHwTnOm8m592srLU6x6jMNwTVqL1dZScoFv4HQNGDtclM6HznTFabemof6ZgiKf
8Rgrkj/ND7AiXDpBdL4g9Pb/W6uTzWi2f2gYcN3jZn/AlzMGA5Y7GFck2fTwrnXX
2//i3pTWl/khey98dn7NyYyW8OK9GdXh74OgW7/RV49W4hGgiF/bhhUeYFPdGc8B
DKsnxpan0Mm/8ePRfLbCLS5fCPRvNLRmJduH2MA7DPqEA70JMnncTopvz5fgceJc
4XC+BC/TcuQyu8oG7EYL/xzEj+yVGsG1snuuaUTbTFWe6nNDLdzTYZtps8UFocka
wGRhEx0Gf7oIyJUviiPwzeXrR52gvxC8R8RS/yapqD7L3y8D/kSEv5dZTVCYPRxc
DktJ11nBecxNfHpaKIdGQHQMWPOqxmYdHRz1EH9q1fPk4l2hnDaoYXZOMdx6H7yc
Zg88HoGTGD3uECoKRznS1BE9DpNyUROaWdg4ZFvoDxS0MTyMxItoXfM/0p/nRfkP
gUm1+XfkAA753Z336ylPC8azGePRAS0z2ZxLK7CwdnSUK9A0XmdpOflsJGRuUXQx
m0U9a2imIZZ1MBHVQYmbsp/IjesQbBqZtnNtpjViFAmqWqLlaWW84K35buMeiwOJ
g4vBYDEgTOQfTdMXv08MBfX6d7jYO0NCQSKrZOWmYqhYE+K7zvxDDpOFtnp11TFX
iCoZwQVz+c4FixZ2l0CKzR2+tQaUIkkkeR9CsUzNr+e7pBx1SgS8/9lQgE/wprdx
uN0vRcaSXJE5VgyJ5paDOc+oNJ3T6o+qHes6y05xSDofOiaQUBf8fWDYOsTV71rq
y70bGoQw3IKFq/fwVK1qaYKvOTnNvbWnq/w9sZlzbNEMkxEu4pMbJYOeYFBs88tt
UnnAFXRpB47efWBjRJId53dOrGHu1w6MIC/tv369jYU2jkcqClmx9AAyapHN02di
IhWonUGW7TbDHS3m4e1cPbQXO+1sDFQecVpWo7py2Qy9u7aDHZb+UzsMUKS9yCaa
xrIhEdB0d8ULbjQRemwKh2eXeOkBNxJt4Tw4zXhFlQzKF/a3sOWVYPiisJG0hjzv
zwSqvo/+A4uHfmHZkuhzOz9kfXwLRhjTwh3ibLuv8ts0ufdyPkjgKJf55pW38N1Y
tCAo7gIe3vHI32BGxgfOK/CgqYH5UOrZk8FDbQ35czKPSnTJuaSGBIybH+9+sWpZ
umk0CX8cS+VF5ygAKF1Ux6qRof+4tHBlZl3E8dK28No+Qhy8m2Ay0Cuo62ypD0co
V3F9CQR4wNfxkmPVjylN5ac/M4CCX5yqxuZRRoy70GR6noIw5NubM/yuQW9MODWC
7tuXecdy7dl/wcOWNeCtZciX9EDaBchlhA5c3t3mS0S1FXr78Kpx6STxUkJSw8mq
62nNwybEajEANXkSc2o50XpseOVDQTXOOR/KFZqPr0LoLEJTM+koFCfB+XkVbZ3O
7t2ZHRuQWMxwTxZcx9hkkIR2cjc2G/wuCNgM+UuQyeuXxS4G7AyCBDwsNMmg2w6w
5ap6dtBobmTZF9x5OqTlM2YofPByQW5l36AEy201OXstQXcBWSVve1BzeP0k8Hd/
l+q2vmfpy134x1eQkjWMs14aTH+0awr9nVz8ti3/9CP8w5/gIa26b39VwYXMsPXG
zpC8BT3dkL1WtSQ3Jviv7QxZ7yQninvB2JRJFI0Cb+Pps97fpMr3yKy9ffbH+IL4
3F9HKsV2zntFEQZshg02mFDITJ9Dl82rb+XudWxePmHMZGKy1tb6xoJCrNSR6kwQ
K2KAGZZf6axf1wTOCODG3ppOwQ3YUl4/rXKs2mDn71LOtEP+LcPxIdQ0Fr0lho8l
e5UFuMJAKFECikyVTT5o7tYUcex34dBWfWX488ahJIHEakOuOehdfkD0dhc3VRz8
E0g7iMLTJeqT4hvVJBZctjGoMAYgsbnU4dhSIkgfFu2JKHwl9HQgkEN4R/IKgWOO
BgctWHgrLLvooknkBgiv4j87q5CHxf/5A/oblUO4r8ckgHdemSHdXm2MqmnSfw4d
wjPJ2/UPDB75C5OK3GxI2c0vn3ZHVo5WVpW8OaE4seeenEg2DoiN7OCZvMLQwNNN
kQTm2RCfejRS7a0y6pHrg/ePzxT2t9Lifge/zLtNcnNA2YYJldXI3ZcLSUd02Rgi
wtNl5XAy7ro8POL5WLbxgqKyV/3tlWdrSm16R66/GaFglHt3b3//M0cFwAmhBOcN
jvxzgiUH7P+UX2qwlJpZsg==
`protect END_PROTECTED
