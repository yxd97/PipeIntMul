`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yaJCsv7fLeEu084+upLQ47Ta0f5qMr9yV0VN+j9Tc6qOdZqRmuHUqsQJvoEhhGHQ
HHuQdMboxfgP1n17uoQwv0XGUa5EM3UYUcJZnWS1FZIiyLcDFNZi1uss6Ee0uOtj
byXb1+20UF6f9nu+fWQePi/NFnDQSkABBceXo01FctCNsjlQIABI0dIwMrem1///
ezl1/uUNOK8SFjNswUrSwJlXeq0rnT6FUtOGbRKIOLx1iAYYMUZ9lKHFLaEXOlIv
YPUnhv0gwBg3XFSfVgxDXiJQtbvnbo0cC7U/T7PHNcVfvfSwHtod/56050ZZp44B
b6H7LJ4/4elh9YwQxGsmQ3GtmGzWALPtZVtoQ1tABrute3mtqaEc78Veayo62H2N
NqknRZhdlxBz6w58TylbQfR0CQruaczeK6OAHyiepbzk9g1b1FFRNIHSiKurz3mU
kuxypFPfrTVGDbHmQJ0PM0wMa5MZnPnJ1BAqHpa8mRT9yUP/oY2mjszje3D0fFjO
ISBpjYQAdZwZ5+66xnfG2GIIWkqcxm9xeufllE+Y8KUS1HJAzgk8h82FDiv8nXSU
b0ZGeBYYtXuJZ6ocbhRhImaZmqm24W7XlUg6FvdkEqV3wNF+bH+k+kdEqCgKmnJN
Sr3RVJ7jr0LaRjtygAl6k75+vuu51ENd0UJ7W2gkTq6lJBv9KXqMvwVfhMyPPdZp
JIo3DmTkwMbq9JooV3i9J2saAid6wLjaU4PRzDVe9uhJNn6Z+SgfVJBEfdM0QVrR
4oAt6XNpt04BU8BB/3ddrDByr+xeDSfPnxmuM5nBUwFRBCxkhxfGM8BHAl3EljZk
p+IfKyIHzaDdVf7piaCMPAEVPDRzN/H9vSbe5/I8pM9ZEaRUap0cPPUhB7QxkqD9
AU1LVwb05XySxUSRrXzcKsdF54gD4haLn+kUW9BJ5Teiw+A0NlZ+7kOKRuqArt+8
YzTInFsY9koGJTQk/jNvZrIOxkPJm1eMpbL/PBHEs6LjugwxQCez2azfLrf8/2nn
U5CGA/E8CDasafy0WOVFj0rP/ixgWUNp0EUDDw6I4Al7VGT235Qed9mxEwWVvjj/
8Kek3Ab52XDAIv3MyGFcqHiP21FMyDh8e7ZgGiFFGVYjdD+dYYYXQcpAXHsQQmTw
MZcpjiytDHBSdS+Cq6+9ugseGoBM2pUz4uSyxsa19cqYRTwcxGK6zvySl+WOIe7A
k3/FNZaSIskQZQstuPD/K2axyl7E+fZ0DDjtlVx8nH2UmxMZkS6zeh5zBMBDSG3G
P9MWaqOrLa8vZwVjNdIahAs6robSpiARtc42EEVGcUQOB91Sr3/CyIy4qwvDLSME
x20WyFjsedYr10iGUz9DZPgLu3+rBI6R93jVOVs5vjeXcv8h43wK3hqgkILQRCLd
mgqox1GEY3iJ/wEOjzBtPgNc8irDfnoMDl5ZQFj9guoNjTYl1ck0Js7T5an8t3AI
Dxb7uw9Prd9bsku6/bhFvWXyNmrWf3AUHWaJZshW5U4=
`protect END_PROTECTED
