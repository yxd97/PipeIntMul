`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hzxD62LBaw/OxNEqp/M70vxKGAh3BTrdif9tMhtvw3R6tokuecBgixNy49hXxgMe
gI/tpR+4QjJ/BnOVLUh4Iyk12xLLvhfMMrKLx5opt5NcmsmCG8fLYaV6mxKAj4tq
umrEKE6/sTVCfW45xh2m1rSHgs23AhggNTZ3vbVOV9gFiuXp4LiNRbcks6vqvL9/
XPxjJYyDl3NvLgif0VyP3ZC+BTzPJIe0FJ7FzDNDSguiKh4ta06c4kOoUOjUkqSJ
cFKm4IS6OW3LbzUuWiKoi1v3WDuMsvTWxe8p2d3CWTNSah7oCkE0bCyQXgz02JG4
9jvTGa0nHZ3v3vR4TKgOmoPEQOjG2ZG3FjLRepcpyQ0bwlQNRg1ir7ROugapy6dd
6PYYUWIUMD+k+FoWoUiEBxYZ1CZH8rdDuKPIAkTsTaC95729eSAEF/B2yOFxEcgt
A+2TnhXZMbwGMWjSPY7PPSXtsfaT+f6injOsYcpy7p9yPOehADz2F/mnhD7w1wZy
B5tWFh+PSudxoevwo/+QHc/PaKEGsYyA+Kd7N9qdCV8Iv2NBbML/ZMMKXQGOZyGf
zRf0ylqz2i0iBs95Hf37k/a7iHs+HTBHI53t3b/yWFiL3w9gOgBK8Z88pAQyxACi
KSN/GE9dUKz6Hyo3I8rg5cXuGYZetqIQ+kgi2/zzQjlfTD/CejT3zKYe1ZbMD4Q2
RkGecdMTyIy8P8U+0yStOExMfGs5Uf2AznofMYfFWbNCSiMiVAcekbzvRqgSL5kT
KuNixIRKFi9CUjQJNdThJpALtPHnTsq4F2JwLdKsu5OJwwR6h+npTqp1nGGz3xUX
gqw4QJWlsCy7sMoQsWbJakWUwKfgRupsQSOIs8WdSP0YHgH08ZnZN5yJG5izmMT+
gdR7hqem0LPvuhMSOLYD+A9RnrKzbNUo7A0uJcKlNqpPUeMO4XW/G2ehIr32LJEJ
`protect END_PROTECTED
