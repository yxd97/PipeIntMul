`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDfQTIbn6OF/Drls2tEO6FF+MZdR+B+l/pwVTt1q2LFLwSJuYOF4f0Rj5AXFpH5t
r9JHRjRGCJtQwWzvpjf0k/WJ8qKfZbTAaIsWntBA6s4IIm9GxUi5BSC76ElnQ1BJ
OhyX4Y2UsO9f/kYminjDbcqaNU4w4mSGgO9SFGAKuPt5IgffKMbgfduKaEwGb+K5
URgRBKfy2g+XyE0b6WNH3ss0OlNRqHzXHK1dJ+SA70DOLRYSoC0HqmNOlwr0ettx
hcx2DvNcqGAMo3Ows2Yu3kCd+b2yeEfXWBMH0210JaII2pfR9xZ4gmzwAOJYvWfU
7TpYLbFVAsPkYGlxZzjRNd01sU5BYul1Cx0FtxcuoFkfNk8F480Zgw2G5HMJzKHT
2hV8LtT7z39LUC61iU9Ru28+apGaoWt+4zo0U9IJjUoLbcX9jRGa0q29JAarmaFo
9EdsW4+Ar2Z4NiawdbfHd7rAOc30rdFWD9IodPG3UYskx1abWwgCexeyBLPvFcJY
o/HMOR+UXQuPJqNGCgzjHvivAQYRMbSvlj9uqUDnVH5DuJXlBo4wEI59ehR9BwlT
qMG8S6Rg2WOto2eWzFVlPnNQu2SpWHDBbkxOrACO5+eZ0bX52XIbSjIvoBUzzm0h
P8tfQxKj0hnkWpTM1h1FlnLX4pB306eG8QbxxwStJltNsa6dDvsFquyqQS4OvZd6
xMyZm9tr/zqHm53nq8Mrh9GhTJYJjnUBnMNpjRgfhil0cS0o8rbNTldK3ks53jZl
ed0qELzm4N3nopIxqULIueI50BpHnOjk1krrpszoBhxa9kR5dCtA8XPJu1XTbXI7
PEyeLPlCy3XTdhanY1eK/UKsNh1XwJmDOQvu82cz1CtmjRgx+UTltpj+e+A/X7dc
r5DtaWf4dY9XgVCO3WdQ+9IXOKDEoQqua0rbgfW4NTxvsAxmZwbBlYNnujjqZsef
/kr7dU13q5PL/p8TlU/mHpbjgjSYRN2uW3S3B0ggmCrcFLnIYry6fbmDZlAVWhTM
TCFcnXOzmzL3mZp9+SUi9E80ASZOoHdRWU5DKhkFU5SDFrgYHbvvkDp1AZ3XU5yv
8CnDXG9IrzTpeygsAbmsOvZ7y8czmf8VsydvEhLxxaP0jR17flBTG9ycrA6pttgU
WgHW5heojfZa9Gt6tNgr9jYkJRrbM5S1ataoCKdDephmk1+4rA0pL01EXk+AYlrH
f5q94PEvAsyU00e2xuI9cpmNVKqWCmZ7tHpuNPFWE34CjJYo3G80p7+bOqNSzc81
+kXDFNUqJTVSnfNNgvfw/j8CEwscA8eX1Ld/59rxlgbyqdtmrIcHT5a0fzfrSmvF
U1o+9iiAw+OqxBmVlv4CYDDISzkSBTh0kZS9U09mzS/Qs7aqTbHSgCjDf44RLqh3
U8xPbpbBLFDTDFVOpNuLj0UKjJoW7rRd2c5u9nYt+e8r7lCuaFZ8Zpo+l2/SC0EE
SvED5nijnqxAPqbL9SjaJ2Lc+wliH4GnqXmX9+B/KQXJSjabjEm/9d7hCNLVt/YC
Q+pOoq/P5goEpOjte2yfoSZlhob70M3JopdZr8B4qSstJ7g5wx4NICGABIb/bpC+
MhR37emCAnVV2eKR2UlOl4kWhAEqYbnk7unNc3tcWgkJrn90/DX1fdxZ6qSLctEE
pCTAnnWag+mATGKNnZ6hCQpuFqR6KU3mpCnoFKSTVSV+P0F8aO5iy1x522dfH3/9
j45xc6caK/lNF4WKH1C41xPXbawyu9LgzFNmRU2Kn93woDPCgEoAho2+gtDKm0zN
U9O50K73K+lb+l/1dSvHlS2BhrEzDck1nsCNijgBBAtYG+lpFl/2s0YKKPpwYZqf
YiwZlkz2CHE7ZbKZccBM2eJZuXInJPS0J47ngnpp4V6unKS7DErXtrYW2eJOPR5u
zXT7KT/zKsqEkojkXOTv2SW+Es1Z6mWr4lZ6ziYaPV8xgiye1ZsGBXo791sppUm6
CNaoZM2hRw/tdIXAkH5jNW7Ea5BGqMyTgCDPL5XmqfaDd5cKMUtQyukNpEF1b5wq
y0W7PMHbAGZKXHamLkiH2kxb9CoSlfH3wIyxNiJOQhpCsAJIJA1x2nlrujTVb+S1
zFsCW93bmUjgdZToLVLH84k8/d+I14j7TrJtEFDp3441E6oxPtowOu3BtWYlnGra
DevyGuGH79osbrSqG6/kxyQBuqk63f/n6mbwMiXKcSAKNNlFQTwPm3uuO+8SaWAq
N+1MtVxYS/nt3UJg0dazHnOL4wfCLuisiJsp1EWAwrhzohGd75DulGQNc+bcB3p9
47QPo2J4mh8Xv4d/dHrz0R0nM7lFGvYIh/0R2guQlXFKjY/dtKI4UQYMHPB5IrkE
DY25njCvXkifSxM5dn6+FT+wsOTFgzOfk2I+tucLmDLnNsHfwmrhcoGzgqWixI7k
xJOPvBTyd1ts5l/T7MZci1pBReaH4PmNroe0Yi9YCKeUIPR184jijANPzB763TJY
9atK3qOMfQk6KCh14BWGGSkG0H5U+ZUgQRoL6rE6Nvo4mbuMt53wZhfJISooZxdH
9FBXGgI8KDdK03gE0guzPnZE6VfBxCxqCkSerIY0zART0jqVF09GdI0r8ho6VTi4
Jo3iu95fRkl+/n0Ck++C/dZX+z7rpzkaruMR7Ysh8C9lh/yjn/WC1kTJseR12p6e
GDaNAzaca8MY0j+GTq8nYNYLiMMBkOUwv/Wqv7DrlJ3sWs2KOmLORqwmkMkiq5U1
z7hZGM7yApjJNxm53w6Vgf8xGkcWVDY+9wGpAGSMsW81aNT/NfnJHhb2dNsBJ1Rd
rq20BEK8N2kUHhOnz8hx+w+rLJaLuLA8ywOYTq0JoE5OX9LvCq10x0ulKcCbB75K
QEqhTtCHtOCP0pImyIu5B8P+SkF/yaYwK3BaHp4zBIbkVMXK+dwHNmQNqg4Tp7ph
B8unc3+f2HlB6dy99KzAVfd2FHLHXTYA/fNhNLNV8bOLnbew+138LhdANIv/tRvo
o+BDKR4QAUom6DjcrbOmWEUAz8LYo9iajxdlJTqSzgPTYjtUcN7kPfn1Y19Ov3K9
T78aJMNW92lg0an4Xs0kJE0rkvpDKSbF3IBX5zOOKl5AntarhJULTTPlaDN12Sv2
JEPadm/c9X2sWk0+olyRrAd6pe3DpVEzONiix5dLf24v6ehFs013YYxHS3CM9j8E
TI8la16q+Xkd78JFioqYwgLKasuvLdY1zjjWrQjgpeCit+rfSyYrf5c/8EGQbBEl
v8FlSGseG4exTfd50pK5clFKvcNRgOob6qMq388095mesFX8y9phIDMbAD+8nNfL
k3BFZSIwlPMRy5VsuK3ltrpR2fHw4+7fPnW1e82hyDFNJKbpNjQtiN+4FLp6UYof
zMi5cyBZtnPBLbCbb88dcZQJZJXXFUrlpI1QQIJAI7RBouRyOor6hmjJuj/rUzWP
VpUv+TyefRSaNe3jmln3mC8AKqVTb19/KfnDZjgq1QprDAHvx3o3FayhVtkbyeE/
noMYi9A4iozmLoSnAsOfac/xR++AB3xNAKGwZXyMmb4ByCsfoqooaBIjkanBAUxn
bw3WCeT5LyX/J3zuW1fRRjhvaTvUVlVCXPO4rkNkccQc/Xp3o+t9041p3ekWD+1N
XqHvkZh+wtf9eM2EMIz4g/vrybIX+R3IgAg5MZHCBcG3DhssMeUzwI9iCU1MZZQZ
yR6ozZQyZ2CAE/mU5Xj+9xTZ8ZfywIEgsWTK0bzmuxWLcx45x1ysUCF8Ux15eWHU
ZWERQ7ojd9QNUUN7onUoo5yXc51omkXMUHPkYwNG/Jeblm7m2foWjlvCsEsvgveI
1dfQ2q63DBMlwVfcaN0Pq9U89QxTGbZ3z76iFWcK+MBrfuI2wBKRud9XxZQ3r9y0
EmDNXj271OnHmrofSwD+A9SqqYnvP8xyOoiLBPgx99ZBSdGOW1AObegHbTPeraMJ
UzU6BE1Dfui7IJywNvsDpl0rH7cimD0ZLIx5S4K/AJB648QcMSwGv+3VHlWjnJNm
Mt7mNUXvD3jcmrKR43cU1ll114tblD2D/y2nOrLBwlZIXkMP4qxvpDfEz89ZFJrr
CEbCngT1U2UBhFoYP7H4nD3SH9YcINdLmw5NE9Q94M5GOhUO6ydbIj7IQql36Ces
iN4AYLRH5JBIXEhVlhchwejJ/lwFWG9CCn/UTj8H5t8vVxxfeDk/sYmhrzeNgeQn
vf3ox6vQ0AxazV6grE9mRMxmikvoNW4dsqIcY7ruI8hXuxRZzXfVYqn7qHiSyb2R
EKLL0xibWAsUIW52eJ4Ei34xIFVAyAw0GRdSoU5qQB7YhLMG/uKlrG2xtBvueRzW
ps4J+B/GmZ2+BIitqP72KMVglRFRsLGBHT+WUpVmggomudpgZ6pkaGGs1dsF3MbW
Uyja7eg3FpqVhTHb3tJxJ32GIYYtqeShkvktScyj9qd5T8umLTZv93BWTgy/RNmU
2pI3hnolZhDD8loSGD9ZG0ZzrTdlRhF38iVumjp5DHJFnuRU7a2zsM2xT1hobQbv
tZd6Sx4dxKKpBSLYGV+RsPWqNpsIQGeW+2ZmCYo/Ogo6iU4d+lMJmqhchWjKNJWA
8pRojVm6WnEeAZnapFk+/Qho8wrh7OMkY+N0B0ynO1SQMkU3tyABZBBEeKPA10PO
n/JPu3WPyb9Wadea8KpEhTloOFb65AB3wxEXUup/rfw8acfqTwR4hIeCo+0IERDi
THRwVZa5VIltzwrhf9C1xnqpSKfP0p0/SrP+SySYhFQ+aTegN+gH7ADpUGZey5US
UQZhSqepLFyGaHz/00ZBGRTWplWgJNEpUcK2YYaO0d2ufpTJ1J2gfJh++UcAvqfr
Rcm99OYSGomZJOe4gMr67WS0ljHPbvvTJN2VU1Yr5FtWE+htxrs/PEnReQL0oKuJ
iWBAeTWDIHbWk/Z4k0rnDQ13d8sDvXzwbcS6uQkUtjYPyUJGj4EnXbDa6zoYF0So
r96lr0SgTXvYueIKiutGEY3cwZpaonyu0apvvAkXxIqwTZqKJadIpE9Azm5GDvJc
6dkhViL9YBudcHF5VLMMRL8KY95JCtNqFBY9RCv28XZxpI53d2OVWlk8pcsxF1Nr
dxrKLSyPgA1t0qHS+ZLUm7IDGqecVLp+xs4GFUpuh1ysc4bma8geaY9rNlxu+rZy
3w0a2oc7fm+AW1RneSL9/c2iZUTMm3AB5HTKEqPTwD8+oS03vff2KckzE+M/GNCK
TZZ4JLp4/C56k/Tfx8DeJCrL754Kn+BmD+f26yUfZ+bSm+DpLQSsG22ZVUzto6k2
MxIQ9IGBANZiKu7oHl9z3ByBMXHGOG7WjI4JA8Wqx3ZMeggWpJPDffBMRyzF0xCG
6vEdDPfz8apjJYOroRq4El19pSEP/KtYL1U61SjFOGjsUehSlHlRNi2979Gg1oGg
vZLoKP6Uzp63zoOHoToberkB8oInheGEvStDub9UCQvOXa/91k7mU1GQ7yL2GHgE
7LH4sJ3hUZNGZKEJ6N5AvaP2gMop0NAM2gnDKT/0V9ibuCOYE2Wsfns7gO3KQwt/
sGK6NaKTCk5yNuHD3CxkJWNfDzlB893b/Db2r+e0Lw+pSq0XUBxCTCkXKa9bS4X3
K8wcU3WMwi+cxT1Zf72neAS9Nnxi3q6cgTSarJ5Nkw2asx9pRSIBFay67lV7rkzE
CcBQuY5t/cJ/BgyMeGc9ArtY9/XZAPj2inN+wnXgOK70ik5rDyTZ7pzw6HbxApbY
YoVpB0ThAV1WDfFylZqv3shEzXGZGieauloAIq5sslCH6E2ebHJb8RnRGweOIzYe
0StuNPBmVUI5EpY05j42f57aghChx0DbZGX8oc9pzIq6oyMHfT2ejbmbOqfJzcLj
6KvyKPELHjFpH0ES6k5JHygmeE7p4a6Gmq5IeY+YXqWl/DsBRglj7REAptYxc3Ky
NA7ZFQydDAk/aMSO7E6AbKWoj5DgbKl7tX54Qdhnt6y+6tKRYUqFl7UpWC9j7xVQ
wP9XRfkfn+CKG/u6DK66mYBJSlJ0i/XzrGYdvuMmUfoMpq3BomnYz6l4x53mIPDo
CoYOpHWGMfVbcBN420zm/+g2J39rnUGgJA1M1sevP4ps718cKgCAOEDflp2XEv2t
2TCN1FdcbLEYbTBh2f5E9XaXTcW52Ino1Juo0DOPIfe7ocI1t769++BeZc/oWocM
EUgBK78spQhF2gEvQT0YbmspaTl/4JC+JUchxNfgR5AhJA+MpanTpxOG+etD18cV
vLPRQeP930nHoKIanCL8D52sPOhtWdJJosL/6HQTKZL8ckZ6AMD5XYZx5roT/21a
dAqwTpiREGDyixuFEQa3C8mzALCZdRru2qdumNcMuOlUXlhb4L73z1XlfEPVi7YO
BDuQu9hYOPx26GKskMNvdARd7FYILp6nmmwlD300EaZhD7Dw5puZQwnYgmJVj/mH
ozvU/81p8gVJ+AOmUr+1lD/Zod0+eOrAjVwHCD7a59D+JA4OUaRE5SQ/QFRQ3Hw1
RrZgOTW5VmOOp6aOBTHmrt1Tj0ziUpyElIynrGceLJhqA3jKCPRFW2/btYq4UQoR
+JTCoarb5NHPdFglgJ3mlZoLXYDsRr9N6fAeSNaKX4NTxDiNkvRatiXjU6VO3NCL
o26+ayqAf1nb3MIcXz+urlS2PVPRlXju75tyfTMynMQgSMZCtpAj5KJCcpY2iv2o
F7XS+21VT1g4xzMoZR83vCIQzOZAtf60CguMh17FV4HwdrVyMtsvAvVETVZMbzq9
SAhIghQvkKWzHcgOj71WQcL3ZQc5ERY64xpR18eP636ihNpyEAv58zXrUp/LghU9
fHr4ezL0c1nquJSxyCXX0N/CaFMP9bxjR/QsFZg/zCIeK+632muAN+U2hiT4chLO
zhFVxT25S4L6r6bx7KjZqPN0Idfm1NQJh+8N0UO6yiS1cLv4UIvkQo9NjpMBtHeQ
crTpuxCRShsiL3vMfDHPuIjTLc31doKHCJ7lQnbN+fCEGpW7ZTbQxCkFeyAXK6uz
YpKhc0Pg/u+T/HIpRnasz+6D2x8Kz4IgkzIznc9p4Hm4tzhgSx/rJRwHt38acLXj
sNyLSll1sZrc2OE3XHcq6jjBLS8ReUHjiszOU47v3rKReb5lHwWFOz6WAyoBOg68
shFxLgMjatig0TJbzsZohp815yNy/c2a80jntcbbG3YzbUKK7otOQq/tO5wqZ0hw
ud7wHO9DjqLbcT1hxJ+ovNxxph6je9knBstUjL//N7yDe3pDcxoj/X7s03Lyh53E
PsRkrJ8RV7GK7fShI6jDVq+tweplcDLBNreDKreJb8NhAbWLQHb1N29/WsB3sE/y
NhhF+DLS/Lqu8pxBuKrEg2CRajwQCR20lMVkQKd4IndnXaZp3z7TnKcUcj4R+Ps0
5CNyxa1zl/TOdMN5Ws2R/3MMkdjHw2qGzGISIYyOP0qbELXA2viYnT3+vQLgTk32
cMqlQYf2smjEy63FOabXGvRjvSAQLBusu8dm/jEKBafAmiCgKuwO7gp4iA/9bmAT
7BcjoIKFPEyzb5jal0eb+yOzPjgtfSNq9qUYhVZym2897wKt0EshaidDQGsIiq5X
wgK8IFMyzByRW6fPCoPOePz/3W4o26AJwA4YAysqvwJ2INxyZkNExCWUOnYLqcSN
XgJQnRhy6JhMtY0M7OA3MJaRw8DGv9E/6GQEfBGXcAGUB5bZln8cPbD7e67QoPP8
clQow8rqGUxTuc9dHVq/MNvY6hd8e1JXzQUI84akNeGwKQCnn++3xG3XwXLvuJhR
fCHKjdELSLHgwWUlCAIedn9BvYaLJPNZpoUmLFoQ/vwoMkZP3wqsefO3XdGAv0Zf
Zowm3FvCBl1VIrcNu/PyhULiEgl22QNHYeh3UclkB5GCx3YosJSFxioVAPss9gua
eSfH/luxq+11myeeENunf05nHX4uI4aM8josswSfeQ6baCOncPN8/Da42NlDm+W4
/osVkli9xzZ+fTAVnQrtdp/soKT2aK4Luw4XGR0xvE9CZV6wsutBC1+xvLaTcrJH
dOR/Zz4r7Cn9nuh9IGOm02vr1JITSvLG/nR9uT7maULZiELekxiW7dDnCKEv5iGA
qPW0x3/mSCJPB9q+9hAi3kxsPhW5ZHmhtBGK2Y4AtnqgfEJkAeB2aKSD7ZsBYv5f
oYK8g4Wzb0s1fdiAjbuToJEjMEJ8b6vfFg8egVNwHwc2PMz2oPwJvsxmVFfTJZSc
qmFzgojbl70i/KfxG2cltRLJosKsXQu1JuzW0JRsrGitMVq0X3wS/U2b/cBLXYKM
bjz75BnPsMMju23YE+885XW7ntSttEGm80E5rQfMmcQkrktwVTVtiaEHslpicgV+
H7AjsDLTbmAdApNhyAXIp541mjqJfrITwUIRTSmYR3DWASN/OJrDsqLzhS/Pdw+U
RPFwctM0hOdqjyArArBmpkD7004WQdkrElaTNzzvJRK9pcahVGj0CSMduPj0CZ+W
K4K38LP2oEJcuU4ULi+wY0pLK8y7vXxxbgS5sl5SHII71m+Lu6F8iA5XTYHk+f7M
Epar9LOjbG3N7JrMll4jIkH5ELrWZtDj0JtvmWpfyCdi2mP3oyrkKWg4SBcjt6e0
NBCdqTZlUEcOgQhD7d4vglOyx+FCJVx2W+uKBkgzcDrmuJmLv9veADfiISRIVaam
+0rDIc/R9gB5lN4rM03guiIUVOBO8Cl4ll1VM2tNaq6ivJiIZI69JbU3dF+NkkQX
lwDwxGtNiK93im1WU+0qpRYcao678wBT2Z204wTfMwNBl1+7KPRlWlXuO/FXBCrD
uF9k2bTydEUxzHiEp6XU0ugf4IzTh/rywJaIpuLodyrX70NUOr6jZdspMmzvp1IU
2HD9CSAYrZe74RlO0LIuV7BEdVlsFdlJnah1VU7I6ufOIVYgQRIceQWk26nmMpzB
TunCQSYXXfQS3zM/RiI+kfQTLIjZbWcY6sbm+MMupAdqOfsPUjiTjFsIXybaW213
9nuwBFXR1IlYyNK4hIuRQmpNA71+hfKYksGET0WyPuWR9u5X3H6fHyrVTtoApa1E
0d2c9iWYcve9FefM2IkphPtWj99KxNJayCHSLnacOBqAtD6yR0yLSH/0ZW37NsEL
/CpY3JQPlOEMB81TMsSHP9wqDCRiPEK5C75Hs1SjndHHdxjtZUSz7wobRoaBRaTH
vgD7PmESVHjZ1h95lhcVbzfCR9BEHDaUZEIyM6m4abflMnBRavpz04mbO9d5OsRu
xXrLHp5ylYUSgVgzRtePdtejIIPM8kUO2VSj41GtZuvL/c9pNogro9aheE8/jowD
dE4bQaaMP9jqQsUtGNwxBJlE9TayfxbUrtdRiOnApiXjxNzIoMl5rvROJVDIqVdX
gg3rlARZU3wl1akttuZaZS04t/TeK4VEBGQ0deRf2fDalmqSJD0LtJ3AcrlIKRg5
gs0gypNb+RB86+FJDjkgXE+6lvpm6KzEwXLGgrC/mnxJZWrgn36eIgYw9mZ8a1hA
4HpMEu+xhCjTpsxcnacRh0w1KkVnDeItV+yT2Vone00RmA1D9aU51XDVKkoB8YWz
ByRmIxw9Zn7GDM85CEV+/aHiOo8KmEXsx7nvCZL9nV5vcEUCuXjmCNqJUbVkZqX6
Nk4pDC2+dLO1HBDtcH63SvUqg6dwMOxhN5ZWuquxc8h0wCcwVsAJcFkAX0eOxYlr
ibfLG8S5AOKPgK6vrwYBCCPGQhmKRAhjNhdFfUCEv7DonsiflA+ViC4JuBWkLOHr
wTwS5ZR0e4dwJiZCJZEKOk9l24mJR4Ra4rKwg4EohMA8BKQXonnHelq469IodAEX
+opsD6OXSm1tkNT6wkEyD2gxqBolMFXe2Je/7DBOlpsU0Ngz/9T/VZ3vXgSwstVf
jtfxH3s2vtn3XemvAs4J6DATNW5dLQtQu88/skcQC0qaPXemjcXiVOC1OIYYwjt5
5+URlw/2CVxGpJIDhgft2HHTZhd8SrXGknd9hE2Wfhdt+as+rDD9WK6FiQfTDY6q
G6ZWTrheoAGajCEYWEcm4+V4gk3xk67nYc6UbJVcDtgngosKjZja8FOH9r3F2u1m
ciK8r5YUbbSY9XQLo02kimJSheC5c0Jd0DKvnhljrS+4SkP6Y3hHApNhg9d9/Jp/
n6IUYa5fcdjReJymdnBvhXrZchJFpKOXB7kzT7q9D6anpOF4/d8nQjzMAf6i2L9y
hP0HF+XxRMmssrXPlktgKME7neXxeCAmBuvqGUmOoCWWkIL4BtGtl574j//o4bAd
+MEayqS7W+Y7WI5itItqxyJxJGq6W4aXUPw24HOc8tncQ66L/MXofbne6VQFzyI+
qrMm9yN1AFBWlaGe0SjYUI+mvryGpUqRxEQz0U63Ug02darf2mSeF2xrBwlXlzgu
CqyWud7giOY2N86lSc+qQRAJQAe+mc3JTJMfNEISgobtkL1cjTU8otcIFnvq+x7q
hZOTYx1PcE5lDAYc9oCHaupZc1a9ltxtZISBLgNQ5b0fEv0OGmwqFphcEw4CZVNE
vfklXuuaEBJjIAU3y572zG+KkgtT4/McCXiaZUZ2rbJhxernkRBBaDHyHhDPP78q
go3UYBbCtRpjIE2pGTrf/vrlfWT2usigqzdCrYG2o9rjirSl17R3HNjJtDNSt/T5
YjzR+vBoKneJgdC8FePwnCfzDYXcxKYCMUlqBoEhiZ2YIB4ivSeg9hZcdHPx9nV/
SRa81PPImUorKFJwSZHwPs1F1a15WBIRlVx20gms9m8KykF4uYiYynZoZ8ex5Gwm
M8r81lHON1w6g6pzGwQsbHeXKx86I22xzDsakAktj5e+j8HXefRr2mtQz1mUapgk
bCvWWIW6dNz4tTUUgiuQh7D0s3oUedoQkljPrSBxuws2+JM6QK8EcDoQRwBrxAXr
qW/V/GUS8lH765wWaDqNYNC34l4nj9mnZA02+TmCIzhej3ggAWigMhLjkb5mFmsM
XP7+E0DW2X5W6h1sUDN+Tm36DTnFey8suYY9p29SO2Wl6XT67alRw5RyMT2RGn1b
jqrU7BCChhCKj45Y9J8bsJWsdsFt3elmPq/mDpCHu5GHmVWQcNFwx8VnRm6YFijq
7tLAvUpo4n+Xj46C4M2mKId7eoMm3wcw18pFhI4x3I5fiJa9ZjaspqdpDFy+5kK9
wUKbe0t1qjWkuvKvW0iCcG6WOYljgEYvsk6dmr+N3pY2cRscQ9DSUSiVR01IW0A1
EdomQkr0dlfqMYCnU5P9l1mpdMiIZeEvPrS9aNo6UHdR+N/VmjD19aocdk2MiBS0
14vO65CUgvKULrPXD5HZ0VLVvApBAxac+2iTBP7E2lz0a8wPrE0DRimN5ptWmJYr
au9UrkQgKlqS5fhjWLxdGeO95NzbMtH1FRZQnwKGKnuuaBvPk4BHnugsd6SeG8dX
4hVmrvPJmjPdL3vLe59xikTXj1LivfInFHlTqIYpx8IWP1o6MMXlEu8+kTovqeyB
VIanhpnOVgOwc1WekpkQGvkRCTfGKankMguN+IOT4T94N8zwwhzVWwxNxJJPReV+
7KUoIt/mqOi00LAqR/668+8gEriLnBeJp3yGRkaw/c2HM1iQ0qCQRa6G7K/2QObK
qHn9Vd39fkUJqeuLE/DKPE6thc0J/jM7dcRjlDqUo4dHVnstGFRPBXudeMtsC5M9
YmwwHpuKfGKqGv0ZzORnSHXp8dETAZmclS1Ob9nWFkrqSlZjW74dxnwHSdNZaqAt
zyKXYlq2bEUUkem7GQo9/d4kpCOzD7I/xyd/2QUeM5oqjcgqKdrVh+ahe1itcg45
6MtVfnKPbXgCHhG9JpZ9vxLKKct0UyGOAFa6gsSDpRU2QFXHjXO/enig+7X3KRbN
XnEkXWnAdB/4by1srJFIQ3ZKHOjHFTXufjQ0ftD+NTdvyzayqmFCVlg/702KnFOD
X6v22bq7E7cqVcOuG8HgHQr3yZuiHlzJIx50GiPQJ6ST0kBhFPdX/vPBfZWsPHY2
3C9B7Db3GcN3XF2LDWVt3+pmoQsNuOZI8Kz0BGp3JpFuwqoNUaF8AmmmwnHBVf7r
3D/IEcGy9bCiFE/2HYGpvYbaOtmWUtfk2xgbNvmg+pzmAG7BiQNHmzRDX55W6D9J
CbXbSDmFwBox+bfrj1ALg2nS+/CqISKJgdENGC95xSyNUtoKX6ctMPAmSk6/Jiqo
CwpXkzYP1i+h9z8TgWnGhn+ed6WWJWF9HBrlNnWg6n3F2dneXy6weMu6qjZvdjg1
sHif93O5jMprRrB39Khknm+k7vJMACLUP/R7IpdCJ5M5JnJHMfoWKbYjyHU3txvW
6FABzKBXX9cj1TdS7HxpR9RXPNezqZcH2qiDxK+3uibKAnH/4O0A35ZS1nO90HUt
f59cNxYIjkuWTGeziZamKl+gTLFvANQ7lQsQLIKQsTuGJ3nRYCc3b9MjcBKdJjqB
pgHCGK9+dfWuhqWBEIr+1Ms5J1cvj1fFTB+X2qHkBOZLi16dZ94rYINamOFx40qZ
eYi1QtkpNGCjq9h2SUGcFbNB3Wn7TGEZgpAtVVZsPN/xW2H2LnWJ8vhiQ9nvtSH2
w2rIhk2pxB5aQLPbaw8KFPJVTSMMwRQd0Kzx4xxKra8I+no3nh51KKUUQ4XLvAx/
OUso9jmSpojLBtZIK8+N0bZfAMEtoq917vNVNJhFO+mM2JB/dhvrnQw/+N2FcV6e
uZKxCSG2WGx9ofzIas01qZtLkDR5xqWFh0woY9uohInzHzs0VCWS63jVvsQgC4ZV
0KUEukWXM3YLSSgh9MMaZdYS79DS0aa48aQlSi2WKvnNbyRQZ7G6foUqpFY9qTuv
7/cEkN0+tgjf6pwFWIh1KAWejscztcdDGDkJVhJbneWXazfxpa/fhZ/tsWX63lw2
1VlHPIOt6Z+JK7qPU00Ze0kIyrlucfp9Jpl+kkamqgZX+fWFBkXHimejLiGCtmhP
PsKrPcP4VXRZGCcZXdpKRgaFmwVO4091EX7NxbHLH4dwUtuYjOCQB9v1YHn811pA
hem+uurDo7PEM3uQbUuutBrsyrVvY6UfL7AChEbwHBJGMQ9WCw0MQKTgQQJKBKlZ
yyrjNGEfR8QGZddyM3VyUAFMtoRVYADLwGiW4uLP1LpIOm+D5C4efaGoWCmh0G/6
hiwjclMe4ioMGA1Ga4oXc7lAPF2JvDXzoAS/n8F0O4q9SWb+/o7hWl0JPcC8l2op
Vrsar3h5DUuBuIl0JzmuNieb0eHUdrS+jOOtCvUmdWVtsu3/0B6VWJb0InSo5AtD
gHDxn2Pcx8IK3E7YniqaAu+4rlCrBSvVSjAbTZteqasDCqQjMgGCCrKstkKQL/2/
Iu+AcD5xtkPIAvoCPH7dia9MmSNKPtN9hrUwQl9TrfgKZn6wMx/JN3+xOSinCV9v
aDbOFfHXxKaAbVclMwWjh8x8l0X00cF9XOznnfX8+Gg3Qu0Ns50dv6rlHdyPu8Yw
IHTSQEJVbfcQDrYZ1dMWrXU5IICRvCcnlnchP5oaZehBRjJaPldmhBVMx0Hp1fGG
xkfxmpoNSz9qCTt9+zqMl76IWpItLSWDemDs80OCXyzfzkoNuSB3JNafU9ymrdTS
c43pXceZqnIyNSCAZQuOEXHvkxPaACWzca30k2rX+Xcpv/b3tz5ndlFsh02cwQBE
R0t0U1BLgp6pOtciH2JduHM+8TOriuZntyVVf49mvmqIu7mJYlfvXMo0hUGyhAuh
iJlwIE7TIzhW+/E2mzMNvfkk0+YsXV15jwP2KL8RNfK2vLUhRBdrfHtxsVwr70r/
9aFhlQdYPKLKPUxVlwvUqfVQ5qNQAnztSPpl3N8O9hEqBfGQt5U1SialQvsgK8VN
Ju5VeIiNf2rQD2AyewnlywmzYnO/qwB6lg92kUIgDdYMq9OjMHbbM2rJvAsCVllD
6Xo5qXfbH86jl9IxCDN6+9IQeZAhKDQurVTQsIZj1HgNJM2SdSdtloCxtAlyPchA
vu5gFjXVtbpwHPblIQlkXt2dttoPslLegRagsmLLXte04U7+LPMcWmDRoKF4jrB4
uS1dqcwipMsbEqYtcNX1ziPbjtnvrdJDkw0JIIv+Cb0XJjFn/86bh+j+KmmdY2Gy
Up4F05cN35pWQKIPwpmvh5Wa7n9r/HEb65P9pIHbS8jROAcf8sM9pfGwcS2bwmqM
g6pNnaxUj8ssasab5oDYQacP0QoRKuZyVPdT1umtBwFl18jgPY22/qEeBX4ldVbP
IHedDGQf/Qi+GeOTCWa/88mzu3ZsFZOtqCQUGrGqtBbBIib4EOyFhBYAqqIj/lSy
70OsVwn1FHnLGpSZ4v89lbzsBwENTFs9KYx2I/RrwsrhWBbeQv6p3+9NjsKkSJ0c
80CeXkSlK8q0FW2OO97zrvQx545LZtvobrf9DZYaLQudZDDDVBI84pl3V1J3JFA6
roR7RI1YxiUFRB8TVsU6AmVmdTtlOXVShwriP2a0DaN6u+qpbPbRuSfomMi/K5AM
/MqqD1nx8CoBkhcl3AIju4tIduXLSDJGzJN7OAOBWW5+0NpgRO/B+LXg1Pc/FWG4
OkyoqoKKALPyRauEMa9Nkf6TxDUt4WLHbilvjpdGxnqz8t19yeu1orKrjGxRI4nn
KOeQH7U1KiDAA4JDyfYcepVrgB3N+47nZfe0G2cwY7ZLxmvoBccQzMsAdI6X2VFx
lAB7bDLVZQp6U9kYigP1d+tR184I7fEP0XLHbeQaMm7UkSjEjBHv/C5XzGyGagcu
VUVY3XZP5lZNn1qRVfvSdShWvyguIWWpmF0JCfA7LNnVKDDyrglGLEEfe0A1KG7o
uDGd4ByEHXHpZbs+ONuqSNos7QGVjYx9GX4GjdXJf3S8jcxh99nNmAFgKTknjuGE
qZjjlsUkB4KSa6+Hf8aSy+JniNQqnCr520307jD6vBWdXBNW/+A3x6ahED5MKhON
xno+7dP09YmA/elLZeWkMJxU+dEoN7CM2gA9gJJs/XmAB5AimW0iAkArtDyOpl5E
fnNSeUQ1OQgmnvvPfXmmMQMNlxrArma4j+LgFd3eU/UF1tCbJxk47YoBjvExcCAb
Cb/HmozkmFGMChWMfgLPG6vZmk2xpAtvyO4EQIKdkiei63EBMLnELtJ9gbKIU0c4
Bb8OatQpvKpKBy+seyFKrugb+Y2G6JF6d6BOITnKXgM7UO2L8wBRmgs/mCM/HPdv
kEySzbrbRGq0HCp+9+5YBFbwC7aV98OFzojBQQvW9LuTidiZJMc0T5pUbFk2LDRr
YJgf0IdOYChzAi7nOe9vNAN0G52yDe5CxaRymX8ry1Z1ZfZ/UFzmP+kjXeFJbZUI
P69L/t5hBeL9R5PvAuP7AVNkuGFTodfF5JarD4fUv2ifr0b6OVF/PSrEuwqfWRn7
pitKAtYWAMeRd4wf+QP4/xkFFYZt7mmQx3US/YBleANr1UbQHtC50EJdm9j5cvXE
STTC0ErOJuw6SiM9sEZ1zKxvDPs7wGCxdgjmfVrQhis5hjriTkflze5ENOEdYmTw
c0KAZ7cvw03rCYStXJ0ab1PiJGH7sAWyHM8IoAqBjoQEBn8a8SD4FanzHiZO4BbL
a9toupUYnRjQsiGxhnBI9JOF4tQ51Jhy5vVYyXWlNzNzNyWyk6bC89ejTBa4/gH3
TeNeBZLH2VzB2JbrKszZsJ6CPPtCkpTg+fHGk+zqNvyxpJm7J9nGZ85I12D8yKgT
g8gFMlIG/EdxdYbQ/pqwqZI+ClVs3H0fJ/jhtiM1IHGHZhLdjcj5pW8VMHmKRFzQ
lUhEL8W58lxW3WJodQw7b5QcHDm7jee7gMriWbgyOnpoXgIYdbtVXnhGjzwXVeFh
PFaR+6Hotz3BQyETI6hkf1M5eFgW4y7Jls01sTAkLMV7fAIqyyF5cta9Up+XhEMK
vPKNf3mw8wQSh/E6wCWxCH4eS/Zuc2j2COWwu1BKzFfR8dTo3dW23C0F+bCHQIHD
dsRHiPnfchz/5pKEF4ym0kuwpX5EMdOwRhzR5pxiKWLoMgga/ZbmGOLTHJgRzTez
rhJbvLwF4TE4zE6dM3a9yN4H6g+QH4iSx1XvzQZpA6b++8rE5B5sqMJ8M1in8/40
Ht3eWh7/PVc0/fR8b56zY/+FNbx4uPeQwJW5R1c/+wIJJkFII+L7b1bLoZ6F34vM
IDeaqTcOou9AHjxbzjBYxeDZQ1dMhDQVlxQWqcnkYj3wzBf0nUAmu0e3Kv9vdMZP
+gcH6kVb50qnMR1OMPNXY/2FgRIiyEnKAv3Dy80DmHHPAoLXGpQ4Vpqh1UbBfIU9
ronC3HIr+S+j1Wgw7c8OxOqMcDeQaGTri+hqJOv1Lq4q+8zI0u3DYveuri7GrnxW
b4lS9vHGZmOxpfUN4LASRDImWj+yjxKgnKiuRUAk7Zqwa6YJWth/QP9UaqX//NE8
JuDuttWDUq7wgVPM5qLsYUzpQyqyhA0T9pTr1cEUQjTMQWnurNcWJg/o+smRCrX1
hXs2TEk/6keusyCCnwXC7gOSp0lFBAE2ZQYIpk3WJb9YSd80k6zCmsyAJwYcp6uy
ESZXa1jmm2BK+zqRychubTHmxWZL6oichnS0iG91DBf9MhSA5ftzTRXxx+X79WC8
g8t16AC9b3WVv+BIctsX8jblIgz81OG9PAg0cLSGaJBogf/f7+dfX8gyKMxE5ikY
duzOVpvAcTcUdMnE3A+UKIJKg3r1jd6XCmcFhx24GW48Se2oPD/k8qMze5E4HOv3
HuJDHTCvbcPnDX8fHgwStJtLzJQIr+5Zq/7u8p0iQy3f4IcBHT861BWcgJOWlI7Q
/wWRoAN98g9KTGEN/JSpSftIKcVzm8hNQLPKGe6/0KOXp4egE1VbZL1L4xkM7RMC
kcF+viQ27Qva/oFFRbQz1HqNG0hE27CQ6mIwXo6uWccBHvSV3Z19U1QrU62vU45f
EMAAF16nMluRWNSkt1Tq3owQNXbYNlh1fQDZhZAl4jjwGuu0VxGrl7u25WdJCK0/
9t05g1UYfPhH3e15jSFZYWxyLsbp8Zngr2eT6RDCmraGryk6XVTW6hJY0n0GPSCn
r+5C8KjjkXqx5h5wxcTCMRxBV9g6v1RPUKp0pPmHSNaz2KR/gDI2eJQ9qY8s/99k
r0IlUXcmSP5cpzkX6dgcsQCK2rj9/30D5f9UYzXZrEKLAtzPCq1BbzJIXn+16u90
QlhOq+L9fjX/GXRMsAKjnwWz5R5FjVxNiJmDPGD79asIZ41CgTv0GDZbXJOvNzFr
G0IFg6ZiQDGqLjEzSBsaUkCRzWjy9irr3qUKYNyegCgiAAf0nHWS+FKp/19/gSlG
vwSK18DmVbJTXTrEF6zJ9AoA7hVZAn3aAEMEKxU/Eo/7F+MpZ8L1TPmgZbNtIvuP
wDe7XkqA3wA509up+psIFQ6M2IHreKJ/H5wlkxcorXunD9Qv/Geb2gvWa3myUpWQ
gE1w09fwOWAMxv3VpQf3NoDt1QUu62gEjHhcRXCNmgdgv1KurJmoMiHSDi4FKU7R
5uEcwqNgH4hV4fZTv7NROLF/CAikQrnFWFoUjK3isgjXu2kPfdbpkaa2JOIk9boP
3tv+REvG5L6zryjDuBDdELEsvJoNLLlLKWjaU/JCQQ14sHAxeTS2y7p7FNltHz9u
Pg4wO8huU9xZ1bYIaQyELjI52k/Afl8HjrkZQ/QKatHIeDWdwlIPz6ZU6h/826oA
DiSX0dT/k9fSdsgtmWeP9OVkcIzCBKKLf77tdhRwBn+6baWOdjErRya55uNxOxs1
P2pRIJ9Oa/Wn1rG7OZih6ot0SlL99t5WYKfimMD/+CDppmIzyOW7IOV41qzvYh1r
8slBxuMRL0H3MdoYYB1lR7YqfAMBHhO9JyD6gVTd8/RCy+WWcIDFMK3cojpWp2H6
FFIOJP1TKrt6IhApwwwIG0txbAHFT7yruxTK5aSR5qwrQ6DdyVyzoyCMQwXIoHzP
FbMsrasi3MUIxVrWzNvZcJY7+M4nStrfya6K7GTIzNDXzeaGGWezp9vOaJ9fo/Jn
JIVbXxinHQKWikL54AgaS4muvzKqcAi1s+Ge1x1nIeuphNPIQ9b8Q6d+SLSyv8b1
IfjOC2ENEBUL7TwXzgQPd/sDpN6U53XIJgYA5T7CATVq+eg/YTZiozQmRRrjZQkL
PuiJaZw6vfiHp2KMWi19+uIgusa0SiaGQIdXYjj1/tWH5elDOeyxOiiE1p+mtMsN
mLEbvUPefPLmDnXMw1ZXVP0WvG0pdRKEx+bg68zvarHKAbxAjS9gk9X5UcP5DOeo
BJ6vBIoYNpLy60maf2nlhbTWLT94HKTZcNsK/ffox9vaiGoCjIkVGvPbNFEbhU9c
KesY1HcUuAYenUZNEIUt8V/PkY1Rlf9zc+zmufCcUJO74xhOWiaSHIuwRTu8JXBQ
/egcXubD9rfzrVFYfUCPbCUXPmYs+s6gdHwgLKIzQ0W2k0zEByIn+ZMEmanjiBFs
a7sv0ghw6g/2BFune8kRqrCNXIZMhVZP98toHhJgnHNqdaJ3Tst2OuWIwEptY3ht
Ydh4ME/BiL2eWSAQImCazCc9sjyZ5pDWN2So0d7O5pI9lYNYdn7FbMSUMUaQ1mrO
opSkcvAQioUB8adT0hAlbC6TwjaveGuaVLsP2kJ2HToR8AotHmUVc42/qgOCrkDX
qoN5iwQkwEe2azPODIxXO7m8nhs1tUDHRtmTI/0cZRuW9RUOZb+BWoPnbWCyesrs
g8ZxP+bA5pCOAWuV+AHj5i1Hj0raVtQx9GroiCNqMSEW5V8bPX9PlVF0yC6Uy/PD
LpFrmTojUDJ5Bo1EE17I1JaqJTvaG8alhDc56IKd34pgFTHgslVVf6XzFL9CvL1n
JjZE5ItGMxCrTVCGjmLG/HwxV3mKyOneBf/taGU9U+z+I7C+2LV0YJUKHE8+8XhV
ZscgvTmgtc0AIk9nWtV6cdz87L3gvlPwSn8UduzvktL6j9qfETA3a5nhXVfd/uxK
p3Nj+JYPa0GFUSiDOUNQMUzIiMVKAMEUT04AcMcyqL10k8PIdfqRBgxat62tPqXv
n26TxQTls0ftgEqEwETrJwxWCx9XGH8YA0A53nvArvETJkrnZ8uH2cDXe7oUEnza
XSmpNGc82WTevFMrkyYZp65kB+tm0cTD4XPA9n5dltAVBF0isDfZcYP0NUwiZUta
POyX6jjmFlvtpM0FkOraW7ndv6rihuXvIzucNwEkHoCVjcwtP5qVAnetLGwb8dY+
xXg1dAegCxre+bHDJhHfDzLpb7ToeL/D+GNMPtK3XoylSBPE9Ql2qcWtcNvBj69c
LDoKEj33rsJucrZr3UfXlqlWV67J6y58/gO3qZcEMXPmIwOSxKESWukNL/Qb6Xs8
xGU4fMlXXz55Awb+HBwNOB28e3r8UTXFQCG7G8ukQ94/Imcv3NwE5y5TKjYQo21J
q8XVXCSYJoJo/NR8zbN9E6XT3jUGFh4IJO43rIQnUZ1RqiJNzLV8XmYW0ycPDsYr
OdWqnZKtw0FMiR5V6B/8VxQiDdr26hKIMHhm19wMdXgqGpE6DBlSNTyApfb48r5P
IZE+aEWrn+zFm0dqbxXFAWwX3gp7on0e0FEz7DHpxd70yqh+nxeIUq09ViU/UXw4
ul/SyDYsTYyg8pjhaj1ISUKYrnqbBTClc/rOi8g0WcEFmlb/szt1ayzsPfgdq32v
tbPt0LbUCZmsZ7V2LBGjbrVwV48x0lPEa8FMZdyTma3lEXIU+ndPV/ZOmOXGTFpQ
600Qecf/IHTDYFRUz2RMESMy8COuK3X21wQeQP5CQUpey5C2S8YJwBnfDSKYRHxP
QunWufqwWHuW3Pdt91aqznzk8IqacMRhRjAR2YQkb7DfnAps44WDWHE6P2kWhuwP
hRl58LUSqeT0+9s9SeLV7/Tr/k5Hqjp+WeTa7B8TRPN5vGh8XQmLhx3TK2Pdfw61
xD7l5RIGGIezMr7gZ40KfvVkFIZLj5/4m4pun5PkjQp0Or2TQPi4Gk3SOiBV7uN3
tJ/+vMBE6tk3OS4bqzjSoFLxP3op53JhzC7J7FmbXxH8UtieFzl5c2O/GjVpXrkS
mHcJkwMOOgJ4GUeOjtILOm8lAE7fiCPT9lFOaEaMjkOs3FY2ZWXUvm1Yk9mZZToZ
wyHLyUtfQeXVjKS++XznPp83q0WGpN+Ao2e7WqWl+RlrRw9qd3jzk1yasZHfjQf5
65m3KVmom4X+7k6NR0fFneNF2CYMi1IuK5h3xROdbCywdNC/mOdrR3C/lRwom40p
QhkLQ9ycAdDfEB5X2xPwVup2qxm0ELNJrTHjeQWiL/zhSh47GOaGDkFhQAWBfGlA
bocWQ900LMz1EGwvEY6g5AU2Q7quIAMd5F3OG1xLl8UVtgHaV0ZvvIERGE4/1Etg
wnL43uT2X8hx6Fo6LR74StCJF0Alairu0OEAf6Zppr7m4ocgFh3vccgYhiAUTcq3
khPywLeD/+CJE0OATaytB7OlSdw++ScZ4QJEg+G/PZm0F2myw8Oxd53VjMRtoiXx
K1I+gLP72SQIMkOPFFeO0HOeXQRMQWSQUxjeo1/ror6S1/5NeI3KgmNUJuCyETv9
RYPf7/BXg/1iXM1ppNoz4ncj1dbilTOQ70U3cTUzIiWvnq3+JmS7YSu/JWRAwjK4
JAF7IDa4bjVHU54A7mgwVctBr7abqAmJbjKq5p08Hp4uwEXBY4x366LOY6Zv3nrN
/7NlsTKbPYxgN58LX1KniPe3zA7p00+s9FtfAwrInXEWpGKcRgf5Ke1cdszVf5TX
3v5I4wZFVpPdaxLQLJvt1FRfRPijiwI2e1wxq1idyW5QQFP01pekgRPmKROH2JZT
YxATwi1tweT9XG4PKKnFUgKKDqOQoTSEvXs3eB4g+eMbnBhryfuVAZZv9KJGC8TN
6slpV2NxRdk1okllzHQAMF8LtCWhFz+z9G4cPasVFHD1TXts9WgWzIhAfmUlFcuM
wFUWG7QXgMMBfhn57O1djXjOVhV4XiLSBcFUKCM+4puh2QfpoktR2NkcVNGAH6Ah
Hsnn07RQKDFNR+cOTZ/8k70y+vmQFSdn0xgPoYwlWYXNYXmosIpGBvYQGOaFNUlA
Kkiy79ySUKjDyrxBIqU0AnRVNvtx6UzQW57TfjdiXofijh8o9YgfuBzoMmsSUtXp
Z6mI5NjCvXWNQRL4n+dPZRsGwvTFC2uR8YcoTWp0u6zWh6JvfqTSobqEU86eaE2c
zd4e+Up2BYrEqP4JUuLMyH/MTwIGRWDBJIIHLfU45dsEHpy0we4FE2QNJ6BlzYIA
l1CZYQNGK1f7gYBj/zyaAlQt0hvFQtULRx1pltxKLWulJKaJBZNOzm7bt8ZoKmsy
cePidu2iiuFbzGka1BwyFTiCa0Xoh7ph3sCt8g4cTwABeL7SGhrmYzJxYHHLuIlW
KeS4XljUyQbEZPs4I+p6yCthOP/rr5W+sewIbjZPI8NjCnvBX7LGxasCUIwoFliQ
pQg2PMkEdemORHFeybhFtWgfDt6spjk0SyC04nHdOWK4CVhxbfIecGjvwL/ouINq
X/GnMGAsUn9z5iQe+XUcmDAuBH2sD+3fImDUaD+BK1LkhRMTXBxHPP6YykmEx/uK
`protect END_PROTECTED
