`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1GXKhDXPwK+uxTdQqdmrAdA1qEPsx2byZRS8FyjwwxOqhTs18hzfcfaF98D4d83
/Vb6XW6Bc8cREZ2aZ5ACXHh98dY9U8fux20tld6fCObrHDq4uU5Ha00Gxp94WJN/
jhVzmTnepdsjxj27YV+4VsDpUt0T6AGSSWpGkMnJ4AYb5Y2h5eVA1WB3l/Uoi8AL
FvzZMCVfcmmJQwfFNUgkTfEnAicZMleo9mzf0/heVeLSDlGRw/ziSr9a5oT4g4Xo
1grUj2MJh1fUew96UUS5F/KFpX44ZFLfbsCCHso9sLVB+J+FE3uFdb8qEfdmLPbM
JnsrcT3v382LjM7RrMP1I8jV1cblFRINICclyFggsKxvey8JBrhtCVXmeMbYDcDg
T9UQCiSxQm2rZPuT81unCe4ybbtinOREL+auB0YqIIBw3IC8vHI36NmTOuBpp/P5
siwOXR1gVOlUlXLedIZSMvkGVO3c94IZFAaJ0jXbSaZgmXO7VFKZCHYIrH0bV+vR
fL7TCrrBsAzFXaCnmxJZCKe/mHbLguNloO+MQT2BQVzDqo9qEsinP+w/2hpRq2ed
60w8aZLhHPHFLscELSmwM1mjuSrJgMzKnytymMcSSK7Af2JM/sFx6JyDnWWbyZKu
ULYwjwDvHJfLZbQ/2RBobrg+BSqQd5JHrY+SqRxWtEiJJjNh2IdlgLEpHCKkk57/
t9RvO7HMq/BsmAQUHFlUQCpbseA0ThF5AcaAC9OAcfT5uOlczTFLnOgl6ZUIcyKe
KGBfW//IzunArmkIHNuJqELGFg7s9KxFToUtbQGQN8gLj65NuUMe1JSiqtHnciMR
`protect END_PROTECTED
