`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRDHToZaAZzoYEUIdpbMW6pJa+8vdXybwp44RAsmOZrd7hv6HXahHRoxUEJH8KDQ
OyKN9NqqvK28F/+ppsGYif00EYeYg59MGhek/7yJS03dba+bn/giM6T7b6tLLGbl
3qljU4iB/oM2MKtu+1wTwZa4pcV6xiuk8XiXKIhkUavWmnVMWx/RfA5+6Z/ehf/Q
CrFX55PxQaBchp3Cly9bIZoejH67fqTdbaETX5OdxghOtbu3ho05T0f1K/XjF1xw
YajvWR0qhNEA9sMPkUFmdFjwXuJwFSQvKUGEvLXSk35yYwGh8kauDSQPYhE4NuOH
RdF87q3u1Q+iG2SRK8fXiDmKPlxiQrzWMJOCYVC8Vsxg0xXlWA6z6oZ4dqMgABH8
qnsc+8OW6Ad9AHc4F9clkODHOb/EohSivEIbBGYYLppi9p4IWAWtOcnheKNKWyUb
jwc7d4Qi7XovF4mvyF2Xl7xHxwaDOLdBrgiByfwh2uv8LJo0QuFq0QESBtnm2yq5
MDFbaVa4iLq8ijaq3jNmUV22cbVGidQtW8zOZO5BaFCduaPA2gfY8hFBoVWAbpNW
V5puCMRMrwQgcipuEeiYPc2hfI/HTy1heBkcZBA8aWALQYilTTbyKVKNALWhuMic
V0ztdRnPwrq/K5RN95dFkEbqfxzcxhR3FskdEafbxURqBjUkrLVpLfKz/yGLucQt
YOAu53QdDPho4WMMZBegfTTTA1QTl/Z/PHUxg4i9p4hUHGo0DkeNguAIOcElBzeU
lAW2OGXtGNxFNjJFOYexCA==
`protect END_PROTECTED
