`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbxTvKqvqgpD0JWHWYlEPgxkkniSM34TGLu+dFNgUTAQBrAMUANXlL8b+XwvKdxi
B7A2a6dArlERfptGdghWjQtN+viOgCJOvRa8F/jjJgw6ni0+ck4A/SyY2WZ1Bgpq
htHP/uzIr837S2JW7lkTghyFwh3pXX7ywxd+qTILAGdf9BGVMqUCPptMyhhndp06
xbwr1H2NIIMjFBErmcVKIzqtUphP12lgiQU3DHlKnmzzoMYZ8+Ao8HX1Zi6GIhYP
4u+7jtvcEEtnM7V6vVz0VwJgTNMscy7C2gJx+Ow+/jZ6KA3TeVs3PnFBL2kSQcX2
KfJrJG8MnEt12sNMADgr0w==
`protect END_PROTECTED
