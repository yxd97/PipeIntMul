`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TkMYaLBjbfQV8+TNMguAF9LhsKYFcVjUn6xHbdM7Oj1mMKwBGaMeNxuX49viKj1X
ZaP2er06Fb1AXrqRLv4EH5Z0bmqjOXPEpvBT7/NNLT/49pFSmusZrylwdSLfSKYw
GRSbl7ySxfMDn4QHbfyonV2xwBBTeDjf2B3M32Giq+oQ4sUJyjEfyu13EkDi9nMO
HyIUELUO+WdaesZWtDJtDUWL/pb43zHwa/dn8QM4W2BLhjXKE1OhkVzbBZU/dAEz
3m/MHP5LzvBYLvBAapLUqCPD7jaig6VTJDLTb38vosOU4d1vwNYNotH4sXnmcDBg
PzyEtLa/Qd+c9BE4I1kDWbHR9ksBCeijNXiC/cgVG5A=
`protect END_PROTECTED
