`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ctRv6oH4ey2r/pvDQxURyi3Q/iYNK7uj1FSJ+EGiwdEHCsI91jqSdWrO8ZskwNH
ZWm2GjRPQlBA0YE3dk8uE+VGh8mHp47+k65lQOZt9IFrs3KlZtxQUutEMiIey6YH
5beOUBAbvhLSARrGhXYycxR0x+jPThXUTzsQqkCy2R+TVOTk7jamH6udCdBCKRbR
IpApP05eCzD/99ZbUL98D1ByJ/G0l8eYclibWHzEpQPVO7jQ27OrY/kB/zj9VbGn
DZRtWoajw9FTTP2wSwke7BeWo78a6FTL4xcUe/2pGPk2M/GqJORU2HQ23R392/8r
bUATdlc5XqnUJy68fKoapN6WEzLe2Va1ivb47voCKmfGDbVIGQgtng5fuH8OVbxl
HmQ+bNVjG/MBQ1nNqR5VrpjPo595boBP3dqvcwRpJi2i+agjKbGrm7MBnwvuDcpO
YN8GMB74t2r12tXoLGOB4OMKTSNODvzZR8BnIpGigsNNgRHQqlknd6XKbAJAL8Pn
1nJGJYi9RPCkx7P4VWIcVMRMZi9VD93xOh0HCCQyOvQnhHvDVKiJeouu3LxheZc0
6+Txtka/1pQ25jvYfXzmfWWnxnxqrCLpsWC7af9O+yLVVu0YEq842bkGyAeizdXK
eHOinEnewXXDNN8hvo1/nvN7SkCco1os9vzUkozDy76Ro2S021SAObobIKZts/kF
+oUkOPjBevSUIRrnlfPkRBfeaZxWBuWYI1Eu8woHByo7nQbrLX9IbmXPDEs9nq/U
q7pMb39yB1/a5L3hCZYFhw==
`protect END_PROTECTED
