`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aV6TKilMpkXCGoLqDJvbTkMvjbfzoy/ZKiSrSCaySvZaU6kOEGr2aivUJpCvwsEd
fpKgxqemm9DRmCuUg2pXouGUU3d0Aamv0Gd391Q5Ci0F7bR4xxYQIAG3/f5JySzq
r6ZpXODRXFVxXAMahAbDWzS18mW4AecelnDu32LN+QtJxQQxhzx4tFEfNUO/FY2Q
YSvaB3XoejXjangz8xokLjhCAGkrAGtbVTWUZBEIoVVY8AAt06tDi3taIx/VL7qI
AZeoHJBUItb/fXXRpP9EX4UemaMbv8T77GGurUUO2+I=
`protect END_PROTECTED
