`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ki5ck8DSl0T4zYNjM/DT9pwfiLkZhBUewLHnzRfA05n9FcuQCvsVH2FGcZL1XO3I
xtrrVZub720wBktVf3/Tc3Nf0D2TNgmoi8AQgDjgXMo9SfzMknjLgHGqgap/fuXQ
KDuTT5RzmT8oQ36+J6CH0eQAUYbGNFfnVpZDVtN8oRr3xTYhclE0xvoLDcb1aUzv
vsfH9pIjHrYNqfRtR+m9WAX6zb0HTjfHOS35p7oaCHgIfOS5/owuK9lrMAaAMxdV
KglVGu1y0vMR+vVP5vT7VQAtKJgh1QWoLc/L7+8jDbIja4WkdWOcS5tb9U7aFhoS
at3oNsPWWkVa53w4lkBpSNaZg2WTVT9rFAr2XEOPI+QHWmmtYenfh+Oc67LXidXD
OHWvP0KsC7EKfWG+GSHAKHP0N34//En4Q2El9uai5e6crFYB/NgLcLcGZ3bRk1Gw
wSUPM8B5QTUwvvNexX4cqIo6Sux+YVPfvSEUKurjx33t8h8/djzsCZSgS23tWoFJ
5y9HqgHxk6mmUn6VlCrneTurSpx9tujT8jzECeh0dQHqUVhuEdMRI3ZsDDULSOO+
xkzKTNsa/0iTH7rFiw2YNA==
`protect END_PROTECTED
