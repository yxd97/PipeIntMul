`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+pfNjprG14TMOjE0InZzZwpQbJqQcOHyelLBYXpO09rfnZSIGPKo1DOENgZ9+gb
AHC9An8egYhbHXxqQBKPY8Z7xEifmTCzAYQ4FuZAMW1hrXmxovxmMZmw+r7LFoFe
fOc7warGO+886CBVHFBh/EsurlVMEfCNokEDcOGSiUNmRznGTvOJiyG4h0Na+KJQ
v748i7Sqk2tc6tYGvF78Bdn/Q81Imd6ETTS4TfXhoF70itHIER4r1i/GF+8dGjIe
DUv//FcpbZvDLshNO/Z0nRl2uD/xxtnwAOW98TjjIHQo6Yb2lTYLmC/Z49CinE/x
/g5lCINNqWXu7+cKHWlCxWoM4nC5SxmFHzMNsHJqdIcan/EJGjSeCCOO2EkY3Auj
FYUJE1DZOsSCHhh34iyp91dqtXcwqvqjjtSez+vuadQfyl1OwNIuh1C4zsbyecvu
qyOqlazCCOGaFIBKRt6o0A==
`protect END_PROTECTED
