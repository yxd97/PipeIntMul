`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
37JWqS+w/e1yzef12izZ08vRBX1xg68Vzrvv8usUKpGYYYVy4ztIGBNuD/wqNCw+
q2V0UYJAVI4Iy8l+0+EYh6uCQrjjxuvCaZ7474a//WeE+zkZM7JeIU1n8OhFGas/
txztRkKsKg9ZCPTa8W+Qlscjyjhmz7c/JwP9dQaFYMn1pRvbaPsPau74ckQb3Kfq
IjJfld0Yi6tMajrwxP0EFC2LMP/cR6VMTNYo9XRLzCbVLKQz115Du7QzioEmmXVe
yVM7MbSbnCCjJ9QSgWKPFLTdgRGlyd/5kgJIgfjTuWNqyMbBZoyghOGK2ioBPea+
xanCEJW0hwMUh6blY20dYGuIGaGb573PvqsIF+U5THr9dcYBzQsPCIoiDS2B/Kax
vP5FDTU9MQw+mCQ8RAivquE//vaPi0G0PrpQzO5YofUpEWA3jkUlW1aOQYlmh4a3
1kbg2g/k8DK+EQT97EP+q13ltptwPTqp5SnnAFIPeG419owJoUaH8dUmQ5fbMTHz
1nhbsf1/OK2kFw9+tFPhLkeITwZ4ic6u5LU6VzDul8V9LZOqShmjQ3PS7rDMDLW7
O16/cYXd76sIzDHNTbT+26IbJ0UYL6jfDzRdC0fk3pYssQi6mnaQkigC7eCRTEDD
lWccGp3QgvOFQye82w7ezozWzsqHROAZcGJGejL7GkdxzsPoWIKGC7JX4F1dR1Zg
aNDOKE/d0ns90CTy1OYoE5B5qRgBenbrBZ51iibWYGJrpTALjzjgwC4kxlGE2/gE
BSPedu/CiPYo9J0P/a7ZD+UhoALtLoLKsajsOY/k5NvA/WNFSzxsFB2TwwOc9mjD
orUnSPRWEfalviqHp00Q7TNlyPTyUnlg6B7Fx+X3PBtzhEDP9tQ7l083N/8PG0nE
QuDOAAXg2GOYIPFIGuWK45dV+O3g98UkwtNW+Vsles20QQB63IWv50sIKaj8gsFq
aJMpkeekki4KxhFmorhSkBeOWg45KSv/7Ki9+XBZPEohn8icEp3p2idTzmRKNZtx
jpsG9GJtCUm/XZBHsQybmM06XJLRZRlTubgiA88zIw7yuNqGY6YsupNbTddSwEpt
Rc9pUL8YrHTa3NXDGvMUDbSiSqvBmNKkRxEUUYF9UPiwbYyasDwdXb6fUDVAznTC
v3Zlb097YO40YQn63bDFfYvdMNdkdQ6xRNChO+XxAVTjqbqOCxUtWypqvld3iMwR
zVGrKZIvlIy41Cqahou/hNi4cbnba9Oz7hXBeKZel+lxF8Uhe4w8UY0g7HqY4hff
e63RkUIfson+BJ6VwMxdFGV/F3eDiPLWBoE4P//ukJlfU6j1OneauGwyWEhcfh4Q
L6oFIsxBdqw8pdB5wBhNv6Lf4BfZ2MtAoBXvwWEC+ZujuorcH9+7lthurXzyFsqO
Gqr/csawGchPDPQNMEPh7VfefhF8Wnzlla8RcqeIosCpuAJdZc+GqbsQJeQK0veN
djDvT0J0GtZtClU4eAaHiKZ/L+3wLvo6X+zt39svmZZq6B/+HmOFSVs2aP0nezBk
w3RgRjNIjZsCk609b4uH+hG/NQlZJ44+M/eOZydWXs7fGYVsNrldxkFasI98gZ3X
ZUNhSxlzgw5x/B4b3lkI00T6p/OpBgHbNhEC66vh76dSfrVdsD6CQqIAA7Fr9K4z
kJ032Tl7lLMMFxYBhX90cGPZHopWaSN45ZwgWnlCSn6o9WQ4FlnIPK5nltnm2c5j
XkbtsMMzxetKpghES7y5JaWjHO/GaVOM0TJoLx1uM6avf7nlq53X+aZM1fqC/et7
AdT0TkS969ngIg3HxqCLrd1IWxSdXytQG9MxVNvzJSgCNN5Oq4/rQCQ5BMH7i8pE
NBAFbEel8uKUaxF1zh+hpd1NRHGARJocUyFD8YQj+i4sjVpQ/aVF3KS6+l6fyfmX
M1ll+malTrpCVZhpAxtv3S1ioxuRcYFvqnHE08pqTIAymMIWwa52a7jNcAZClyuI
70kR0zAgqUEj6nw202zNv7Yu7HrM4SrOHFBHF2GrW6CCU2L8fJr59XpnRHbJWnd8
FvkysxL3mR+NdnDD9d74yiAs1VT8kSTk7EFAChwFPld4qclR8Feb1FejP9aIDoe4
6K16bVRrWa64nQBaP75uPv/uwTuaAhwB7S31F2Y75DHUX5gOJSc81Uxfy3Pf9jTE
hj7N/uj5J09knhVOh4r1MCud0hM8aSLurhTGis4Z+HZs7bujlFf7GSJfnXxfgbJU
TBc4q4wGB16V/N8vSq33jyaH/iwXg9CcmfHTLIL2nDPqTPuS4BQsOOxEOGTt4T45
jaeSKQw0PHEZGAvvWTxUlYp6wuMvDhrE8hb1sk2jWK8IPGj66aAYpn+Xpwy8b+tF
FxAYcung1y5J5Hu+AzVaXgQe/UwZ/6OSA4ZA0nOvPd0pzW9SCj2mmTDrUWz/sVxc
R82JqO7a3LzPlvbOTcRKNnHXecVNjoMWS3adNflnAspaeBSIl78xIymhs3GmJ99z
Q3qjy8CwkVNUeM7I1WdGVBcb/7vOm3tBAV88l81l0dDhxPSFJ+TPI0wxhr7XmuBj
6kkHR/zWTCa/6Zfh1HpNDYZvY9uZsH7oWOdR14ZkVeGhaVDyKwBVICdirV/Zm8pp
8XYZqBqjrFafDJzfV/wOvdCDmAHlxggjOhV98tT2PiNJW1FOH0yqk7Kl0n5us72T
9jhFEQKMNJij2xj9YuRiKxzyjCIbIi7TwXvmgI5dP/dnoHiiH6W5EOV0knnPBJsR
Ck8t6WaLNeN4yx0hqL3iMOKdFvjClWqwr3GaKF+4dK+UNPkE/C45y4xQavlb8tA6
laWaPKMRBUGRH13rkSlwJ4INac1VSqe4GwwysS9D69dQTB4ftdoOt9w4zydx2Hav
kHyHVUea90GF+yDwtVglNqOFLOd2x13D3oR18R+Pxve19PK4mdsMmTgD8Xcme8fm
Lx0y9B0G4tSOXbejDPD9v2sLxrOGB4L4I1vKhmPYlMwwSwXU7Uw30vZvDoxYNEbV
9vBcn21Fq7JT7uwAZkYhmDNambvcIZ1TMQ6ZNwCImkrI9e9u296LxISXHqVRIB2u
hp8V1N4fjlP3b4+x7HC7hKTAhKbOiunP6pnG7LeLY8K8Y4REY6lIEH2NP8sXYEx0
LE8Cf4JO4sAz56P7v9TQ6VY3e7ak5WmTQmY6Fv/viMGibbWd5+jeP4A0SjO9s/Kn
wKpjahvJt+eCCN1NWhBHNDPBjBDsx+4lhcfWpJw5/2ZXmObjknp2lzyPFC33M1RB
fjVOEfbnXaP0w+oD4qlV0SHDZvEveRQKyWC1Uqd/+qP9QBWjh2qj4LOZ3VRy4f/t
Xv6WKrutyGjaTLntjUvUAoFnaRo3dVq1FomKTk7VORGgGwdsALR3WOm8qUT3ZoPg
WO2IE05Fel5pSAxVTeJxV7FHu1cX7ME8UBW6EyiCdG2VF2RSfEFIqDcCCkPNxFMR
ZwhObY4I04ncwAZxgNuMiWWLvvvPyNhNQMTFdqFr4fhoti6HYj7rGe0S2bT02fn8
M3lNKBFWSyv7R95xJLqIJTi61V/WgBedKr8jqDSZLD+XWY/bpoVhEBs6+U7CSQZd
DPhR/pdCZNJ7COsuxzjeWuxgau+gUl1oX6UYE3Afgf6tXHNnKBJ1ueVWVX8LpB55
+6Zxwopzv0VypJfhYSdMSalfkgw4dJogqyLkIoVWZirVrhB5uhrO1Teigvws9vjH
BqLMW9DiaRNL1IVFmRtxmtVVWYwabjKDH1nQSMTYHFJmFT84MjbqwyFsF1rT7O8r
Av5q+OuNJ7P3jxmbXkPf8muLnEpQKtLkYoHBXizCj7Xp098QQs+50yI1wIv2yZ+a
ox5p9moIhOPWwbYYfbnI9GgjXjpFir/yic4fCY4p6uurOVyb40lQf07daisEZBuU
jwijSUtQQGA8cyWeYtgIlSf5Qg43x3m77zhUFctTHWsFz6/1ahbYNg7gkdO7ckyQ
oIC0Hw2RKfKRpNXrLmkukuxvj8cQ+CfF19M0hDHYIS+hmUASs09uu/gc1Oy3YUmP
ohKjl1YSiRs+4JccmFUMwWpi7upFRP3nOPA9bBYtbRM3cbxd4LEm42KfXZL4rAU9
/ZeP1FKEJmERybMm530DLyHQCXmf8aOeyBrQKwySNnya5s6fATHBin0g1sIPwcRG
DbbWm/VNZTc/ZVGXgshHtid8HBLVBbPbV1pjYr50Rci+nd9ZwISGgS5DonbNsjtT
H11fvSqhrCXpvtH82FOztYeQqrMYpUrsZ4v2aFTWt8lxqDObJKefkWFcUXHX3oTW
9NWqu+OFi2PMkb3V4UOz7nwNYGoN6bb9td5V1c00RuzMZzrRw+yJ8L0PUk7Bwn2s
CRA/vkM1fFEJvsTBVwGqJsBzz+tD9fxvF391qZnVzWWx13c063TUQPQZ1dNl/p61
opYjZ8N5tafIrlu/czbVGcc85wVIdcSwAqyDIF4nYfNIiYuhj9pC3UqBeGjOWWyk
w2wayyFm6SCXImNhJiOIQOJDNawHgjMlY8yeNh2ilPr41gLmgh5a/lewkqnnZxF7
DJ/LPIF0UhQDuGIHoRw1VSXLVg2D9l78ZPv1eIHlDXctZvqO51567ONxa1P0VM50
cxx6F4GM/K0NB3l/kNOehHJYK2p/DCpvnIgpn7LBIcyUz6G4efgMn2g4qMwfZn+z
r6bqjduJ973Bvc9Oc9sWBrPqDhIJl7CrDtVmFhPZ1Wf1RQEBWjWEbpfghIbBNkXh
jtm9oxwN1fMe1+CeWnYgdNSyF0Lf5NpECyigrX/4CpUjtsdf10wuQ36CAoknt/d9
Wq8gdvOpdGDRDtrcS0pvMVCnHLnf6tVCEpRt/9VpNm6E89wVmFNcI7dxMg68d1h2
1fznKm/YskqjH3aX9wTMMHhyXbiWk+jM3a7xuJvtN3Y=
`protect END_PROTECTED
