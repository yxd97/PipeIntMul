`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OC5OKnYrXrVi56dFMM/OR5VdXtGdhLiGZ6xm6g4PzpqoziZqS5y1qXakv9XvXxWo
6IaQXHWddHBp+8IEqp7KhDzlSqyeN7hYBL98V6/+5XRxWzMBGjgwQBDtbNKzwo0B
hzKNV0AQlVEmjmNcaEp0zI8uRLRCAFXXIxcOJBIij+FuLhVH/tMWmjXMCywEuTq3
nzK8Gs6yW0Q8+MF9wZ+YmA11FdqJ7VXq2KuUWzvuzCFpnYUdm4GpmgUm+taL1LfH
NJ12OfyuODVxJPWdHVY4jwFLwp0SaK+NufmrdHC8QX7CuvrCvB13riUXcjW6WeWA
tLiWTqdM+qHuBk5T2MQb7IjZhDjM48W7RX8ClGzutgec+9SZMDaPiDxWkYMw0CMa
0EzrccVLO7cHkW5LJFId3w==
`protect END_PROTECTED
