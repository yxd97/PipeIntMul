`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjalddPe/HZQec4oefLo0ArgyDP9OhvRzBWA8hSeRg5/YbVHxjf6s1dfinEq1cYr
03s/0dX4df9ixgWqI8ysNK4EbHNC81MQpXm6Ba5W2M6zjs2I0KipVMKhZH+eJVl4
YG5PqhrPnaCn0jwsEL8ojVjqJTcKR+KON4SE/54SmAptWxZ8l0rmUeRNWctYwfWN
VkadAyy7Yv8l7U37c3VltnP1964hQY2yptvosy5plX5SpDvYDI5Xe2qyLmmF8kUd
YgX6zLow9+yVvoG+Q4CJPSnbq7RAH4X0MmiJcsN/pNclMEBwp50rshf3czcLSVPs
IxGwd7oTP1CRzuLo0slOvrxqcDrKERr+Xbodnh5Du5hOEOmM/PSkqKMWNzSvkwl3
SpZtmOZO3JUlpoBcbv6KCIAWqak1g0b27vDIhR2bzzxjmPc6qSZ4J09+Z/1O4aYY
HiwKqU8g28eEMHzjiUm5K63Xkx6T8jiptLmLpxMuE2h46VIKquR/LCr3cSF0nDHE
Pwmm0Mm8qwgYIqQV52Mo63js/arXYwzDBsazJmHZBf56hBTswLYoDVPhhiJBzIv5
kZgpqvf2Ou6+Q3HcAkqSFbOgjBiVZHIIfE58RGEMGK5dmcDNTYqfFH827Z8KySQJ
QpdlNy5SxZZj0uQkNSI6kY8B0MnEMYqgJNFmrz3nS8dxqfKZobyn8mngciu3nqPh
gd5FgMtUwUnvT1Nulp1lbqljR+KwM9DQ+cptyv+7rtrUNdYYnVENppAdTNNlzpXg
7wpYe4u/XDne9WBziFdaOR8pqK1k8jSZ4sYFOzfA0WnVCF2SVU3YNNnu60Ov3tFS
VawYS39B2v5/jrFTQwiSrMQybefYtRgARsHmq9/YKLYxqD6Qxpjr/21jYHvkrKCL
KMMu6r+8jo2JFXjGyQCrjcI1IqvoD+qSczfCVqOSVoLhLeqfQx/+IDav90U6FCGG
ybbivfGK9a6O6NggPG+PFhIc+637v+yTKhZW1MiwIt3TDKepX286gvapE25UULEx
XPCiKrz1U5fNSTl3103V45hNS1dizSuVBk70zN6OwOUU5qIhySLE99Sn0D4jW8Fq
nE/rhAt52n5pYXEfDi95kuX9GzkkeuDm8twNj0eTOED18LwzECUP16ahS9RmUrkK
GuwftR+u+PsStlzbuPV+E5HAR1csyauV02H0joyYapym2+A7wCyedxCxvl4PugE8
OBdGZWbS5B/sdUkYyCB1nUo5la0cdKMwyxI/IjE8Mc6pp4zrECLmohl6etSooHnb
`protect END_PROTECTED
