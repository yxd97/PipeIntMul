`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DI0nU1ljtPALUH2n0T1ai2bBVwgHxJ0w9RNKQYcoDHNK+IuKiC7qjRU9ZS227pD
heMh5Qoa5uZSBK+L8y/mDQl2t7/HqQD+RfPze6uQt0LYkMTk2vvg+da+5C9dD0Mc
zMRfyHKcH62a9nh34LwTYfktx2MNmMHnBi8pC2fLCToX9WMQ6G8lpwfFu+MMz2bZ
aGMJ5yT17lle0UCqEMTwc+D2P+yBUFauwL6x1gFuxHNUULK8Uvjh+W4pEA9/KOqZ
NPIMr6u2qQ3HEhIOc3jZqVxtbThmLeyh/q0VilRDAZWssbf1Gk/HgTdoJgoHNSGs
yKi1LnHjbdH1kUtSk8UhskNaxjIW65tUshaxLCaWmjWVpPH7H2iMcGungyjRhg28
L83JNChjSzMwIM/NP68IEpnFsg4pPFPGu4cqJocYAKl7j9OxkoijIhCFGAU3MJTx
yhVwYd0PITTp41Ups0pHbEiQEEmCIItcmizDYQKvbZhBjcKL6/no6gIhxu1nqIaR
cGEuG4/2Dg+IbqfVIepjHM9zJcEwJ3D9n2P46wtKU0IiG3b6Y13qpabvoXvOEsX3
k05hFeYiBb6TBRw+itC+TmXxfp32ANJfaHqHTgNotRmkg6r0oiXXvg2jRwsDj5IE
VpuBOM/8t63MLIUtYI4Dsyqubl/KXGBIyTKfGBg3t7tuHfWn9UL6taAABXqFkfwm
lLfJpIszlTvYmSroY5We1y16GBY7NGPlWJntolz8CI10bqcGhhMsk/yfqHnDJdhR
0T2pS6vQImxu1uSRRZvhe1Mt+ukqy4Z+5GFYk3Y3pCAqltarO+ZsHlkKcP9PZFc4
RgnQPP/HRWmRS0W82+o026suKtksIPFusvHPMU9UwyR3v4hoD7sdK7k5eE1h/9Fe
rgd54zs27sF8vmfLEHYwnoBBRh2HsL2bWgzg0Ff85Ih6clHvFF1kMil2tPs17vPo
Z9Zh2yjSp/EQzqMXtPzzRBkX3eIZ3xRG4vi2SpWwgEqGCHXYXj6IRgKWVDqJBAcj
ljWk9DAN8z0vkJ16vhxmDFJ6jqsZqgGPJXNMXLUcCAdI7oxZv3ns9XeXrsZ6O/ol
kzi+coXyMl30Irtn6nSBRW865P8K3Tg4PCxYa1pnIhg586I2BgAoZv1Q4GDVgTlF
hfA5NsdI2GiZ/klyamii/Y5oVpW1BkS2w1zc944EqfEU0r5NZlDc9mRU7waLxIb3
MYR0PgvvGqAuDqJwFQ5iTd8q7O1RFoxZ+4E/0QI246UuAg1B6xRTZe+3dusZ5xso
YZjKQGEIatcC8lWDtUkBDQ==
`protect END_PROTECTED
