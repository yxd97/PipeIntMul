`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+XQTsmkKlwB+yE6kp/UPChRZGbKM7poeGhXqo68yfjh7K1n08jvdXMKOjBrNYmyz
9iE0b+pFgNarVihnIGHy1WTAeS4Fv8Cv5bB/jILx9McLMRPVixl+Zt/GQ4rCiqCN
9C40ib9CWGVf4hwBAsGgEVLF5NOU3ahPCPJuq3BQFS5HSZd+0E4lNR4FCK9DaGL0
R8urw6n04LZRK+EJI6Xb1BXRrI2SMgerfaNmCvnTuF1WjFDQfeakIsNJAmxV17wE
mwV500dGmjDqW+c4EYRP5MOUdTSNu02SCz5EC3Hk3pJc2QBCuIMfVHnMyFb/xY0T
aBgL0tdKzjP12prgjXMMNMM4mc6x5A/Uzubk1VQboflWVXRYJKOXQVDuqMKPo09i
F5i+0Zqd9TgiFeW4dmNQ9vzXPZ0gUE2WGTAVndbI1r/Ko9DdNVEBQ72ssingR7vM
BeaOQ++DZS9ZVzSxuxsWcfk2oJx0dnuogq7eDFwvJWt+b+Zqt8yAQ5/ig/x9U546
TOiocgmslqcsPW6/oiHtSEcp6o++rbByZA1+12jaYmf61I3gAaRfSdXdgjUnrMo1
xV+4wqOu4BJ5qQlAIyb0rQ==
`protect END_PROTECTED
