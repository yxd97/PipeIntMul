`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Bfj045qHzcUCHSs5bgFrcLKLCHSbL+79q/HD/yHkwnn/SRChN/o7kqgbilRu+ft
lNy9auWSQJCRcPTZWK8HdwAQmSzHGSc+t8D9u8Yzz0XH7+Y7KiIPUQXOAYrF+eRu
hGMmrAouivCmj3lqSVQH6G4XVXZCpXgTqCwnqeJcIVX8uQA0Q92vxjTuqg5HgIRs
POLlmEyyHS4BHia9p/Co56mvJfdob/jqly2UBsxLPj2hBYmBRS0abR3nuM5wmYFx
JBvvwkDK2Sxs8qXqhgzXbTl5rlxh2YxB9BqrA0iHFb1s3ukBQ6RZtoBukzn/qZuC
YLTG/AuYaYVGmyovhB8iYqlUisfG6+UaCxGJw4CUdPS3ugi5z38U0dwJ075FaukJ
XC71OmTYSkgN7obLQHKjhAHtGBFrbQgFlXjy4EmOwCKYHOe+HbkVpPBdLimjuF4I
xcVOLHCbSgXJAf4530dWqJoJuiC+9P8uxYYc1IY+C7ZS+2x3OAX+CzANGn3uyLuc
SVu1tBSOf1yVzknIAH+ywYhp94NzUiaRdRReIshdb2mblqNMPvYjLth75Q8IqgrE
OJ2PQpTZtcnzBgVTwZY14jbr21Q4yU2hzGsC4xwG+F4iiZy50VtadF7vel4Cvsl2
o5LCV3F73yAhhp0jCJd6uxZpM/P9gcfSP7nhZURuPZLBNYBXTifag4oXpK8rRDSv
dcQRhE3GLVEW6UDdM3nyKbMYpPq5HyWcAXQ0U7W+3sdOdWSwBkaWAos9xBXhSUpw
JvgL5Yn2210E+Svxb1rlr2EEDFI2lyxxmzjUs3vv75a2AeruYOzEwUmTBYe2/QUq
Q/kKqDARVTzjZw17u4EREczv+uNI0OaM54qsBZlZGvz391FiLe+LLX4Q4oCDv8NB
WEeNxyCYAekkEtURKjC+F8gf1gtewtrjhEIFY5tH9cHvxBjPWuPklDiy9YGQW6qD
erSkJbJbv2fshI20ToyzfVuKF9SkF/9nK91zcFDJGo+2Hv4wEGDiUfj5iOpHU1q0
A5AkVncovYlHFKqqtBvr6P5GqnaRNVF4omrQYF42T8nD/hugZZvbrn+RLQcEQJXI
z5mq7v4nQhDoKjnDBUfX0cg0B9V+NRc+XQtLger06QhzP5AZzzd93uG1QU/rNlDr
6fOFl7+RDF61uT6oXFIIPqmUBrzpEp986Ub8HnWJSgd7X30Q0M+QUpiyWhD9aith
0gsP3Sq9lqnQRhlogCm1i1i0V2BMdhphX/10j5XlaitiyVioD1M9XT7I9yIwX9C4
GtCOlws18kieR/sgmEeSU+sr7sKDF7DPge2RY9QQm3QBOQcE5h35fYnA5nDeO9kG
VTMWusmhPyfsZ+4V3ERsPl/1sk78f0Dzvp+geWVJiSpzFtvtrnPFfkoTfr96AkJb
8X7IoMK7S4GEY4FhxmOdXmy0sr/9zNaYxKvfxtDyaOaVj5SDOiLm9YBn/Gh7q7dL
K+wyq/fTBtnnwVg9ktcW44UTHSAmzdpfs9aWoP7cqzHSlYOrQRnoKtV3DPq1O7mQ
kldyQeqiz6zhBI90wmOfBaE2ZPbJjZ+FVCYZWrlSYD4MZeuJlc6p9scJg/XKN/x9
31OKZqMsCzNdC1Ygw00MWUcZsbch3AzIjwwJb7alAdiP8yxizWFRssjWng/2QfcT
NVVy1rmTBnD2BV8RhXP+iFRNEsKYMmwNvBbrBcVikDphGU8zawdNeOBMzzPpQvjA
A0g5/n22d3TX9RW/+LzTFRsGUBjcquNynUiGHhZRG91IwpYN1cvhrHk4iGMW8V2g
4xDFB47LR/yx3pDL8Zlb1V8vG0wymnUcXdw/oWn4uMbZurHnydNZg7wcPyOUc5dA
cXtmE/JEgRx6Tp8Cf/GgZlEPyJWYzMo60SD1kz91qJi/6q5mNw7yn6S8gBQH7Hn/
leY/Ga/42xKZR1DNziDOqxB+Wx7HN6INZ99KUJO8EDnpM6LFVPpV1B868nx3+izp
volMUPB4nRlQq+FVLIvtNe3zAorrQIF6vxqctdhU2g5ZNupEW671+vCWjLJxx4Ai
0qK0oJLedNRt/lSmx7Bhd2OUJwLFkk5HSFDsi3uvaYM0nF39FFDIQDXI9NrE9Glv
nvjfvR1aPkOyZPh0zdRThPnB2P3/AXNyxgQxjE4wwobg60Mt5xdhsDYNtdIST9vH
kZGqFgsvE8rIEo0vl4aekDN4Q1cl5+SMeqMdpaDtcTFLwGHQtWZR4lLKHS3UggGX
VZNxX9MZFlc0shqxFi63ofC6hwu8nJtuSq483hY3221oR7TpZq1NipcYEGGGrthG
FHvbnXLPu9bfo+KQXRxLdn+kNuhJCaSF+5oi52SnLNoDlSdD//ZWYq5jKehtnIGR
bsZhlhmtNHWFKPdj8aK33Giko3JBgDsE0SuHh3RQbLE+/WMFfME47ONcdNVZVjqz
+P5GWLJYebn8W9X0W5xCPbPTSrZpULafh+LDaAK1Drx4UoFmvlk6iLCF4UuLlC7x
pRlRXGxBcwp3SLDXM0HmNj/ozrylL03nvwWzAsZyDWSKk3zEjdwB4inMgw/TIQBA
wduh1cxONTlk01qGxfvpdieGLv/zldQJxid4aBotNnIGNqkKkL4Zr41Qfrv2HkFl
ThjBEqihvAYMx+WOga/o2fnKwPfnn7cjOpCJIPpeMFyT2N9uQe0NAXZlfREO2kSd
eJdEueyG54R5aEHFe/7IU8CKvgK0ZIvbJjD3seTk2EqSehJMNv5+ANHl1ExyB3vo
fs9R0TNUb32TLrd806yj2jOVYEu1/SgZTBaHXymavmKvarZP97D+OD8gqvIid6sB
vnX9ya5KpEAPiagr4AGuyBmiS3/XGVM1KHMFo4ipA5E6FvPf/dkWweagRPpbheUV
x6gf0DKXosd9GP5l53fLfP7rwks535nN0WIp0RmsNckCOpq+90ve0HlzbykxER09
7MDqSFpEi8KjjQVQ7cQtsp0pHiSstgfyVvnTIjvQ8WS1YcSrcpIhOI04KJBx6N+n
RkJOCQ0AP/wO25GGdbPwCC+emK8qtKDiN0E1uWUop1IrZ8nQb3VX1WPFFhMcuEl1
BpQECvlmWzceWMW3i0nh3t3TvLCI80FfcbXJV+abEHNqLAjSoC44HM9LkTsG+H4l
EWwATuFdqM4rD+RGAmRu5pA4BSxD+arlLSYpoW7XkSePeON5EgqxrBMbximgnIFL
MI2EGKgZ8FlsMl/ChsR57HZtTtLzg3d7OpPIRKUoAaJJFR7DGjIN70F1Fa2IwFRd
Yl4oJ8Tua+xAntaYLfY5jX+FscfmStOW5NOJPrFLKg92wjmZkq0MA/ASfUvlSBs5
ZIEG0+h1iFQWT1rOX7nlO1xOnNnsHRbGDlp4NUbmwDvcvAVume7O/XX56NnIuEKA
KVkQk5qL6nlVYZLXrlPv08jErLg+YhSx3KqIzxJh3pnBDXz4gFihohfKW+qvtCHT
Az9DnYPb+G4i1tnznTHTUXdWNcKnio1i1V+o4kCTBeH0PgD81mBTE0CY9Zzpbt0a
nfosujSax2zwjmRVS9etolz5nBr8WDipmTTb7JGUY7kQl/F4vyzUeqYvUB7ETAw+
+r3LvmYwtqE91slFjM936Zal22IqLZxohGjlj4t7L9fHGo9pQOD/y2ipBj3mzkOl
lCwi5Qc/PrrvCQQbUHFQdMUUA7e2sG/k1iuI8cbW4j8=
`protect END_PROTECTED
