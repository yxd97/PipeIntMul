`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AdT/wRqN1J5tPQlidEBsA4qk0XuxCHgLe4ZN7aOvaRS7gLUnyuuN3my/+avuEogC
XQlUGSEop1vUzGClJYgI4cxouYvGCAv6qYQlCY0Er9P+kI7kuBm+XwtHXTTpEx4O
poeProDjzz7gJknfETrlpgszPvg/pvUN7h2bf++5wQnQKjvmesRKrkq7bn3OKM4a
P9Wg2tTRAeqE4BbapY+KD4QhI9KftRZGH7oeDQWIUKEEZxck09ZOv7a2fwhzqAkT
fgO0y8JchALnOOJL7wZ8aG07Cvcu6JN9u64qWUW5JONaDBzg28Hr94Rp4kQYo6ZD
ATEYLgGZAR0Cj8bDtgRPo1zAUX3Bk6SVbMokhR/YQzMIzTGiIEsb4eREmzPahiwD
4sYxbjrZ5fKI1paPijhI+ZQI6zNjLxgzxArxHz5zLgRpEkAKbrBScqo4JIArs9BV
9G8MlyZSoptXa5XniB0776m9w0mUVqUoXIm0nVTBu8TjEIcw2tNsx95opqO+z24Y
pW8L9T+g3slewtEzELRKTwClMdVF0+RcWYNkbQdDqZfjDGBQCd3534+P75M5hoXv
gp1iunfBcfKX2jNmSYKG1Zj4KLViY/Z/6g0T0xoHmB2gAfjE45r2S8N4+D9o4SWH
/01kaUQBq/NvBxjP6cxVStUc/b3Yj0ROX7JipSpsqzU=
`protect END_PROTECTED
