`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yGL+UK9eDdwvnnodOT6frvIKKyDvdICFMqJdJeevFJhV3PXhs4A6qBVlKdM8YRMR
5wpD0aPRvQwfeIZLPuzN6yBUg7W/KqjNRi44HN2zl5xzNlyeqwC/NZPFg++gJvaR
Wfxph4dhFxDDDX7lYAY94uUBZSjoa93wZ9aXgggE4SyTY+qLa3S0yUDF6sGrq1AZ
Jx9Zo5RvjaB1e5UnY7PQm95hNh6UMFtiT8Ewlutu33gb6JCsfSM+ae7e7U1MNrHG
lPdYfslBHxrzee/+NuNj8dWhGORr2b+SC6ky1mMGLe1ucXl+2/bFTrikwDmVIql4
ijTt100Xx6Z6+dgc1BlXtRiozqZjKD8SQrU9at0kmZXfZsXO278UI1e++P0Rblpb
HEYiNOZZTq77VaRFfxpyywhWwS6b92aeFgIuAeQjpvckTXyxcyew5Y4J8FPva90M
zX962136MPiPE4aGskgljd8AkYwPiWnq2gFh8lvsTa6CFRH0eDIAGSk64cXLMA8X
vU1AEyWhsSMwVpYsYlit0EzWAmM+bSnRaZuNVVTjD/Q5+krnlPyUZ0Qm/eUCwT0P
3lj2H/tKxE9UI92s/3wX306ZaHdIgSy+ttVUXQirNvBaOpdvRhF/Tl8EGth6UhuT
B+6cLVnlT67w9rYdFpkv3T0ZCPZjKOURJeQdTTfIve2utdC6o5jlbDnD1qsTF8xi
lQIX2s++pYyZgPnJbrsKJ0K7gH8rjJZXZZ7b+89cebIupXhkwkYw98EbGLv3BLnV
KoRsnLqeEJ6Num1ZTLVnpOq3N3ooeoQnRJt3f9NRA1uQnb/uwZlN4FdZXuRX2YLF
lHlpH2wN6vXkMkfwXQjuSWtUfMgKujYhd1Q3xW1t5i0xMoah8PAkSqIilKs42Y1x
pwpLWYq7nRAX+G41CstIScsi/ygP687PAK8TOJBJhtfeCcb8QAnXWsQytrwmkSP7
zzZbj9iXWdruTtz0WdKAa4FxRKKK6Dd14HwNedUWJJ7Pq/NJWiimW8S3uAydyUKi
cV3AAyZvWyDYWLE/xPCeFSM0rOQaLBgn9eOxlRxC90MAEK4tCq1lQ03jPLlDIuCw
+0KJUwBnu3l3M1iHPZRi4FYdpW/PnMcU8u45bNOj4/90bjuIo4S4BoqqTbXN8QNc
pw83UmaAKqcphLgqxWhy40daHE+rP+QaVT1vqG8Uu0Rs7WnTOFVsiQMktBnNkkXe
Zc8xwXJwj5WTJDSAQVn/sCPSUmoBtHealvBdYyRdNb1fwoN+bdwDg1KagtrcBxQa
9C5ev9ElVVw8LLP4T2XcUWj0XxvQlxYOIP0OHy8Y2l9cRT3ijLe4uGSC5/gJFJSY
WJU/hCN/KEJIThCkt2lRLwL8gMUfanksU9dFOm/owqOm5Z9fqvaPVXiPsmaitBvC
k9cRHD/FOfPI7lzM58fyIW9pEa/LgzinaDhS5c3ZV8CDP8NomQ9120WgeaKvCC+6
qI33I8oLS1xJB/IH8jRMmAFUH8cxOGZTPUaXnmCJvBjhFYQC6A3pEumOGkXaNzFB
3ztLlMrMyoC4nCbzQkxfs5yxFudMraf49FeU76qvQShCgsUUMssJcA6mllVOdCYm
4ji24PqeGqP5UG7gpnYro5NHPpMk0J2zP5mZZLd5z11/ycrUrTP+Erxw+J7NBcer
lPer/YP+OitKyDdnrIkZvhdDltADOtT6sI9s06xAVqy/E3vuMdUOxXP4ebHe7fS/
Ni04OT//bY+b4fbr2iaIxdaNptG4qxmPztNirn8QvdH3fvbQYx6OQfcDlf5L1enP
UKQ2SXGYSOE69SZBhNel7DdYWva+ts4vzppHA3kvdsbgGRS3YZIiqGiUyiWEtZ9G
Q6RbkctQT+noUdHcwa9jdDAKfugQJmvqHFslC6bH+Y/Oq0LqbbLU4IdkHdKG6Fly
R55NDUso45n7U8TLoCZe2Hvb6dDgjd3uRSFytK2SZwp4mkSsESAhbbeDbRlIUKt3
x7Jy3hDZp0mTjW3vmfyFeHDm6+W0mks34GlrN4GAPwVaLKgyvyqHv/FOw6WtHeCH
foD72Kf8zYqoWbE2PkqNXv90I46p7NsS0f6rGkmT5FtkdvFevO4kZOgUo5zd1s9b
Hd/t/0FQvhKkCDQo+wIVBp9o38OYKcebb4fgP7AIxlsqrkC4wzrDOFigHfioWW+b
ZGP0nF/dCCbm9qM2X0E/UZR4pogebD1ac8eR1cNLcFwjhvnR260c6o9PKWN+st4+
WidUzQsnylj2XNZJUkqAmkyQ1tXS5x7NNR+5mqDMivnK6JGTlYxENH0JqB7S4xb4
RcJskxGNnZpU/j7hsoJvs7xWWTYBsOpBI2BF5l3CFlNwJB2hYB+BFOYdXfEGPBqO
LtF192JOvf4x6hXz8JvvmaZ2ZXqZmrMkeG9d4e0h/Rx8fUMUeHGLqAc9VPcgEbmc
XO8VM5z1fxwIVEc2gsQTI0zvrlJrwzX9TSRLqGez1JnYc5Ybs6fIeKXDwduDmiJx
2IKgo+te201GoU5DFtG7JDxVAoUT68uHw40VMjwnNotaSp5c3pytPXKDu77cwHHt
PPV4mxDfb3H9l7f4V9eeWOL2/t8CGfvmYP2NU8X+E7/AKWZjPwpB2OqoVk0dCPeG
pshZomL4hi4riEsDoOWXntSD6tcbcrXDK6eDCgniENEN+0v3RBCxiCT4uBJdjWz7
J89FLvPMx5cv0vA5sCTl0GkoyuvtQKD2Kcx7NSXP3wgclQ5g9gJOqklTHr8o6Kcg
KvRsvzRC0O6BngUpM5rfqLDWh7xiWUORB7+kMpzETNyEJKhBAigNqVbgfuGSKIlo
hqWOBSsfK5zpwDTzPnkmjl25fdvLk57L663673CnbnUA7LTTkpq1Unp1JagMoCIq
jTbNOChDbuL0J4Bm191nF3qXyGdZb+GFYw+ZXcU8UIv+7l8CDJ9oFH/meYr56cFg
AwxO2LM0UEOnqb/uUVVnVvIZf+lPDsLhJNbPTLOk5CxH2Qsyptv2SikCkCQ904U8
kDT+ngH1cRTguqqWkefIDssm264XbgxBV+rGq8ZWsTC1AhF/E9T1GNFOOQj+Mo6F
V/bI3G1TZUNX2C9ew80MRjO0tZSKopWbatIMf6U+RyK5ZPKEigrdhAl22+n5d0Ug
8PaVKzD1GPS7xbc+TbzBdQ4I6yKKxS1ks8+HBtHIG0jd1MklwN5e68ooBPEDwlRz
K6N9m4Zuetu1EQJmhXMBc/vzjDW4NPQ2zDs14Q3bP3bB64B+YBfr4U46Z9zSkWEI
xysASMe76u496dVdnJ+gqk5DlSY26nOPobtJ4rnJZzmw3O4K4ivASFJB0AtQHBCf
9e3V6POiTsslrkTvLZA/O+ohLlWlLJek96Ys7mxLSiQLsMG6AGOGleXxAUwhKEEB
FBZNR0rXSQJXbN4l9I30B1D6e/Y1TUrcqPYTC7xb6B/wJu8owgpoIzDwnKSAACve
oOyowvpiQvCqjlUgRcgslSXYARDu8R1xWd2uHTuzVpuj6kVXeRiw4BfuK5KgH0g4
NMAzIjpYVErh896focy4gsF9pc2fOrZKnBQOUC2p0OmhWWIF+ibbXpB+a0BBhLGu
xU9beGIKqKXFzBjdX8J9T6IvFjrLPjek/3HEMR9FUBWliM4u4MXr1vRjCjetWgRW
aC6Q5c55WhECrLVS/a82CBCrQ7R2EKfsGLat7MDliOOa77jt4U+FVD1IDkWSOTFi
u3RF8oVekxiu2eCarHMB0WSqlrMde/FNoqgTbabNyC2HP4+CiREfZ8LyKhy70oRi
k3ZHKhKyO/ZMrSgIfn3kcZovm65jfk+UHjTNiL7MS4b3eiGZZvq+iVT5shMomdkK
8kQgL1ywywqOaGixnJd5qcAuasmOlmKAMy+5BT+j1pb5A8Bb/4y+wUtyBSphGsx6
pnmwaKCfA8me8iSyyiNRVV6X1CeM+HJmujzQ76yJtlVEp7YADEZuMj1mUdizr9GF
wdfSV3wqec/vJTFH402XGEPrUU++/fx5IE9ozTvbza3evDc3gvBXIrmVV/jYwqYf
StIJbrQIDhDJFleipDdiGAmIlqmwReuXyXaGcDApdoE5CgJZLnvFrK1/AwOJfd7a
f1Nr3suTs6n2mc963wP5SeGnRlG8GNrH7srQBRc0N+GtFG4h55JIQAbfiqwDVdaL
e1ySbbriF9/eK9P/0Oq5J0+e1Sl2uUKI80Z1NkHA0kvgO6V2jxIKkpvlOax6sPRw
OUZ7pK3SdhzxlOVjzFw+JwQQ4DzT8oic9NgHFQsclJvhRB8H6OrmGP4HzG29eRJ0
NDqX+IhoKd0nq1gfXQt8++stO5L97a5UkxW6ytYhST4oWo06HMTsu0u07RR6585L
rSLloY2AMStbOofgI8fOW8sXAGHk+prySgfL+4vYj1jKYS5i98s3w3AN5sRvZAvw
CV1E7CCVu3c/26Q/NPLXrYA4D6dK5HinMSGWENyCq/V6j6gP2FfaRct63iulrKD3
EYN1Nnaymi/ynfjiLVaecMUKApPAyqGYaWL43phg+d9+1zANJ1fJWcpkaRO8ctpk
SDrdD9qvLkluqe8ebXvCzwCXHU8rUypd3nBXwOxJPORsuqgOa8vH4zaTn3HS5iHq
55F7A9PpPqEfp1aiAjU9jTm/kYpHtdrBiiEZDTyYL6XPBsh9hTLzo9gkbxCq0tAx
h06WJM0GbJWuBYsmPWy2QfD3ygVO+r3wU9ex9NhSgWcV4z0ACxEOzdRltGo9i5an
xt8Zhs5d5FlD6mSXUqFxvOlzccKUkB9nQH6GbomvdujlHvV/TmEA8kpFk2BTZigx
r58Oj2zbdeF6ufF3t/p45mO16WtfKW5fa0J3EXvvKsW8S2qrpL+OTcnoQq8l5j4A
UEFP+VHrM5F7VRe4YQmhOMwhL0VYz67cdBZbwcek6Ix3uvRqS9c9GRncUGORbw9Z
qMX2dNASWBttiwwjEP0npaUST4wZ6Gww8an5/6Fb0BQflGI+D/6xDd5BPQUSdYWl
7kNABZyOcW5rmjmskWs6HjyVYCSfLGryCZCX4PwVp7FyYcIxvWW0Z4DpLamCIHSG
v2N5d11339OGOLX18nCeYvd5lFfdFr3YlYnmVJXNgsT/tcabt1sjboJP6iPIYxUZ
8edwSphdFhvLjv9/y8rX+kl9FLkmOgqdCmk1SjMZivy/nu1jrMaOQ3L72TEKO6lN
jgdMJLSHE8e8DjTUSLZtF1ruW9Zmea2Ip3hh+RPAEm3QHDL3qHZGgJMJ+bO7p25G
cXqaZCWAN3B9oakGn5C1y7horT3bL0mNPlzGIx+UGOEgU3TSuQ9/Ang9Q/YzcWye
gjzR/kqrLgzX7byk6yVKVXt+IOLaqLB0le3ztKBuJto3TitCgGXTtK2gjFuM2GP2
U1OEGBA8N3/bpTLTx7y8l8eMuwmDEGYUaYcgQ7Tlp540uly41dVOAGG92osKJ60J
lSmeNfV/W2BmKBeNR8r/2FG2Sxqw8CGL8iswfvr7tpJCoHgHQLwqRxR5CL6oqyyc
bFC0g6cj71cC8S4geVt/g/fGo9XFh650H5ZyKPHXimA=
`protect END_PROTECTED
