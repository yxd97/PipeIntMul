`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgFF9D2/uwkNEUgM2Bv2HuoxDeM0bwgD13eT+ycDUbkQ9SRKIP6igXD+bCxxA5ny
5ILTMZRQYZ9EmiR5FlKm5znxrvToBj2WbTwNwCdRXm2FWo6nEtfaBSAJrdjnMaWf
5RdlW8OvuGfqM/y2WZ2lULviPFUyMXANi+pM35paFHFPyywCMrlyESstEcRYy2tp
GeZbW2K269AYQ5Mzol8yWqVANtEvleSgcnfnTRfOHVtfJIajx7cvZmakm5f0vifk
4diu2+93hOFXP1TvLCvZaYsy6IvkY8L/XUXZ0V073q3iEGuoFrKMiQX+yY4sR0+5
iMnhJMUR5VYBjWDUx7wm1yqM9xvnDUHwYVPaa1g1bABJMNqqyLn+y7k4LuHD7cpB
PfFFl7ZF9wnsth6L+e+cEuBl3gKIgNg0L4P9AYLWulGsAvTL+OLz1a+kMG3WkzOR
5z3BlX0oeA+B/AU/87k/Fscs8ZDYQEi5cCgNl4JDq4ntf+mYuW+CCEBgOlBmnqfC
BFxkM7Y7osgnlTG0zL0stvzvpWf6Gt3Vn7MT+SO/OPA9fY//72yKCMlCPOY5ETiS
zW5Qm3G1tZgYt9GTncJYtOxbltuC6h/S8dGWcp8v+61FlH3hEFNf+3+zJKUHKacT
/ljKGgdf/U+mIIM13UMUxpq6qVlHlenD3i7KpC/qkTS6zR4K/PhYG2s8S0GeD8eN
QYl6e3e7R1/nLAIWbTNmDECrz/nFuIUzddk12MGarcAAFrHQ9e4JwZJ7qWgwy7gG
a5dbR7IydO/ULWKhLfJ+9PxIqrA1b+tHLLJsLXGI06zNVTboDffakvHvfHyax+Iv
daU9ztrUeNbS6Nz9l30aOC70xxDq610Tg/lsdMpoVQHZi/yl6ysvvsZ0ramA8e7V
nFiD995nvVyX04g4zlHZ+0l7yi0/qYGVoBWTLjMPaCdoSLUkXnHvkdE1jnI8+ZDt
`protect END_PROTECTED
