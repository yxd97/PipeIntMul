`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9VKj7QPNFjZxFp+5kSG97d1yMtsF/w6eWM/vdxGfSYKZFOX/P2DuV/m4//jRN+z
u9B2bpWVH25siHwVn1oVO4kq6DKih5JY1MsxwRPjdgGtLrFM3PqB4LVeF19turTt
4e2ujoyeqgleL0EpdarubWAr0wU4BE05P0Y9h+LJYua3QUJNbYuWNcIkWEdLp3hl
F/gEgQgI3ZceHoPbIqBAGwvyam04L4RQ6ksmWRtK3J9IA3dsKy+4EDI2mPttC2bp
F6R7W3IFMv0lR2dNf6kl6p0F39LhmyfF4jgOkrB1ByvZKnV4DZsCB/VgoaOsozG6
Wp2Kv/2oPTGmnIBGCxiP5nVC5aIOhFDWaPeKSiwh8slZlVhWFIHeK/rVOvjzGnpj
zUdcIRfnosG31bg6yNJmz6xi64xmdmv1tn0qrcTe+YY=
`protect END_PROTECTED
