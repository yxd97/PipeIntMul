`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yEJo/+/euRYYZLAO0cfFE+yBYxFalILUN2xuyEYB09XKvvROQP0mEv74C9vr6Boh
m1NlhdF+D5iyf2H75c5T7BzbubUuiiLN5Z2vDg78k/HhVFUAGnxV6sSaoFQHdtee
AqISR//ubTL7Ljivwa9dv6GQmdTi56u62zp8hcbUKPac+NYmBweEQMHlH2J+Z0NS
01m5PAaxA4a1iSi4G1ysZRZpYLEuJUt3ABUdxcWspTlDG36JTXjmy6uB2cHWuQLn
Igi7p3k1TM2DmvMEAZscqzIwt1vcL5AQzAQ1EtrvJpQFDTMKFJFYhxX+cxobJIbn
kWw0k8VRtdNtTYaj2JcgWuLiIMAMLfQ0/RyLVHc+KB4O+lfPR4mQBXJnm/ZfBCjs
cJ3mCLyvaMZvXzfBTML2zxUqjeCKa4mvb8qqaa+9jEpc/cxI1V/j4MWgUmFHr3vB
Za1aYyQEhHFaoty6LfdboB2k1eFDtczO+oZEHCb8/e0PbMc73iiYwKvDQzUII0Nh
dpC0PdTT9BsTbb7RyLKrfC980JBVtX+YgyBW/8W/QTXV4ieHGDAzG1EM7PrSGEiG
FVsShY2yoINM8QEPjMbHmmCqAAbFjKW4jeoJcuRfSkPcjBUHgrWDbJUt1yKUVIiU
iNXL5qyd0OoeJ1uy7KdwFuBrmdxnIJXEJdEEnJBEUplbRZ2TwJR1QMH96W8D3OBu
WI+Xvmq8RtztzanOd4V0bcO4onLkKG0HZ4TXIaq2s5OttpPHdkBRHkDtLN85J6ss
ybvA9DdI0RRB25p6Az6/LVaBamGUxBPXkT/7TbRLQ6IZnSIVpmeVKFe900c0Gluw
RzHxLBt4ReCEmH02GkYwAZwXd1Pyw+nTh7hntW+7B1uony6Y9bOlQfmuzXwsVLrr
Og2e52ksBr3dssUrvKZmvYzF9QztY1r7mmrZ4ILdw+VT7eeXGg+OzysLPLLqBIs4
zSAnBCD9Wf/JSejX18lZ4A==
`protect END_PROTECTED
