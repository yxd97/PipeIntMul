`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naNw3S7Eg/JDac/YF5x8Ig6TmznhkYe19oZiOGYbFvDysh972Xr82TV5XJ8Y7O+F
caPN1QJkJjn/daBatEsK35vqEijNY90Y6PZavCLfOR5y/O9lch3BGE6xCs0zskOW
2KHbbSmxyNHxYuyOWE9n+upegAOeyK3VZB1CX3kwwM/KOg/rCwpcTBPwOTE+WXGd
6ScefutQ0Y8Eggr5JHm9HBfZXCCjZjbpTAErGIz1AVHoll6hGquv46I4CdZ44GTR
9lM2/e+WFxKKzn70PknLnQ==
`protect END_PROTECTED
