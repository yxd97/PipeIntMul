`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/svTj+rFc1LOd7ENZB1qf6h9JYhhDvQRQS+/jhXcmOiOaJta2m7uchqxaqecJ84
bePjBOAjBRXUiyG4IF+I5+ot9zTQh+AXrkrmyaID5mrN5R3EkuiU+qPINH5E9yeK
RQGAryIOoYlyairxJJ/Gk2UaLGcCXcjScEk2D/laaJAnFnCOemS2mErtlAnePbZz
cskodmUT+6eARLGM+XQaQkCubMfpSf07CxoCjp5SB3hqn1WNjcijgdBhvqaVze8/
P7yGA5I1xf0HTphB3qqpVgGBgxE7d22ZN4R1z423F2v/cLeZPjW2MsoPFh1d0fo3
26pKL/5Da7pdV9J016b+xz11d6Jc8gKjWMDLxuj78r8KnWIVGU6yUFPzM4MEABgP
OlnPD29F9BuAVzRiXjv6895pk+6px2GkPx0eU063vAIkpRJWF0lH5akaLzd6/5Ps
aoXWWEhjHqscX4mPcsCykEi/QIIJSOOi4d1nIWp8NPn0GG/DSrpPWY27c/mWdiks
FaCu5b67+IV6ncelYTVDZ/Fw90d674RC+kHbbCooHfMl5GE4XvaX1Pz2x4l7RhIT
5K1YU/RuwyKTO/bI+qm6ltXF5AYb5aFNPRx8+20mfi3bR8+K3dEwbj/6111UbJP5
0n8yKjG0h+HXVm2vbfwwFikf1klk17LqzgmK+ErvJdQT3+7HSYe+3ZMzitvZiccZ
WxX8bCueTxR0PrTz5dcJWfzVpE9NGvmlbHCrelsBDsjSwZZEaHRINE/ywf8/JP1T
KRcvOAL0B+gcWuWGsUV2eG2GYCpunbKaAIX3+HJ7OL934C+kF9YF81w0Xf8BYBxa
pPI9Hv3HSBNo+8eIKAzBP+NYfXWXAcUUyRn9rWIl6Sjvu3EKSGqw/CtqVhZW2h8P
5nDszpTJI5LiBy92iGA0bQ==
`protect END_PROTECTED
