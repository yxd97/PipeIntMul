`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CyD0ozQoScCGB3vZ8Aa9de1j7UhYaqkIgGV22RWrncHhN8VpcfQs0/TMZcn9O4ee
MnhMaE6bI6ijCYFvgJJdvXO5m4BpePZ2OglmffoOXqaRLgLbdq8Ub8ugO0+d1IpH
CZhRnGSrc7UYVV0YJCTcy38On4zL4EuQwP3ory8fS5QjA9SaWylfOysB9VdouJeG
De8yIRldBgpIj4G1wyuJlPvaGZNAVlUJjy0HD7AQoYLy8yc7zeKteU9iqYwbhKE3
/WKmn0n44QwuMzL3Qpw4/kR3+pdKiMokbAAyeyLSCx1+MmFYpzHUcM8t2ARRu1Dh
cF7GF1tf7UaDmbYR00b5ozvzA6st1JcIQhJd7d5gXMfFtBNCxCZSWP2o0ibpGBsq
`protect END_PROTECTED
