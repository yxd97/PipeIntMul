`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w5lAfsY+xLIurWpCCwrllQvAoMEOnoGB8CfE6gysPLaXVduPksrEIdn4HHoJca2q
Xd4Ivgvb0Cf9GZbbRtUnROvdyJ/pfgqalYuzWdh0WVct9P8GLQXd2S/778kiUnFZ
DMuMcVJzJdD9Pgj9crDccb4/H0UYo9km4sHLwbmmcF2UKZgu6aXomC39B34kGXl/
jhGOTHuzqUWPH+pkIdxmcHJBiQCHuLc+SRcUVgJkXKR/38nscKENgNWl3aMbP0Gw
KHXlXbJ8BEyT97vjSCmIahUkVeRAwP/PbFr5ksEQP1y/UXJaQNAWCnzs7ushRgri
080mZ7WwTnyQb0SXhHR7DeI6biWrjSXnoH2EmYQa+ahhN1D1qgHOTXdlaasu4Dgl
9rdil0SwdVc6S2vSXZeTQMbwGGQqQ84hPtVltZe6ZwaaMpzogEzWtSShBWYkKe2a
AiQwWzPl39BGvVwaFUdtqOh/z6lDxbVosRR/jHV6rTQkgWLpEDBbLK6ZuffGPTNE
`protect END_PROTECTED
