`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3pjt38x2D5iCEk4UATKmxyPBfaL2GF/boWrZrA2o8Pa4GcvM6+AYmjByjgUsOuRn
9oWEUT+MTcva3OrG/Z6+elqMQbsMg75ndcxXYUl0ORqpEfWL9CijkwAJaks6S/up
JKKlsuwj3SDmmNkGyyuZJJJ0b7i0d5VtyHc0jBmZF2IQnWgtMf+RsSG79b3Y24F+
d/Hvt3pDTbVFW95uc1IaysATBIhCIzJvvaIiQdFRLbDCkDY2S3YNsM3cNPOqpUYw
Z9Bpt6rUvO0dmIe7MzExhJbq0R7eqEmIke11FIzgqQffJjGY1kcZUIRhxkEsjqPK
UAT6bRKe1x0PH6Jr8hm7FQqCX98aJrOg3w6Tzby4ENW8tGsTMnMBHGv2Noof7o8t
Zyks+CH9FETTbJf3f0vF5PGaUzi7WOxsBZRSzumrTmSkedp+k/Fd2bJ5HpBeYyO6
QlujbIn4nuOEsB/bmdK+9dxEDqaL6COTDRA1KKSN9Y4zTcl4hjX8OElTXUYFUsbS
TAqob/HOJGqvCFTVgXPbLi7119Hw3HTtLbxNF8oTuj6Ti3tLJWG20JjV3cDOp3vP
tlzm8wy8s4zbvB7Lx/2vBjHVysiBlDTdleV1EMqZNh0pg68AYj10iyz4RCcGrdrG
2ZgRZ6FcxjZdp14rpUad8pSlm/d6rEhiUSbsb9kPr736QuTBpa5XQxIM1CsCUyme
bpzvGaK5oM0JdPtK/cmUFCqVRmyZY98HNcDx2pLeQva4Bn4EdD3kPnwjwCY4FFj6
+TXOYJwCV2lS2hQtDLjd9LtkHG9KtCr5hcLvF9AyU/LrYn5tFIA8Heu+iwy90kyr
WhkBLPC9lPil3m2NpHT1niyVS26CuMGAuBwyEudaw8Z/9zuh3F3rpC7uEimtxsD/
AwNk+jxyB2CVC1aZgzq3ZEvbvBVsmSOOIyJhjbppZA4LGzUYouKkUIdYUTAbztm0
YDF4YH94DAuTOlNuFwwxIHCuXWQx4hABVIGRtF6R3Ix4/6LmrWilezbc+sScI11c
iqrHBuFpEVs+GSRrRonPsvH87nEMBmVZsNz28XTYRbrEzcauy4C/ycjbnbAhwncd
zuTg0UnvVxcooCtd1L6yGjZec7hsaUa9z4ewBGeX6QIf4NMB5gf8NbdpFsx/7FWy
1BaSDXBax/3rnnj3F8+daiFhimCmhUoqcOJ8iwZyRTNdgrkAfjgX9R1z+9IltcsO
vFm5Kda707kT2FjIO8ssaAycnbEUmXJfQyZ9lmjmF3HIR12BZGin1fJRhcVZQOvL
XoN9mNlrTsotsKxafxArJ7nOHZIW8F/6arYCLjl+9KAufmuhOLZ4bBd5nVp3QM7j
wDQNc6uYYx+mXDB8yrYLtxcv6Broh2wu74VNLdy7+KEKOesVmpyEAx9jnqNZPKFC
id2JM/74C0Xsoe8uWa8XrU4vo52zdP0VvRYnneqAxS0D7FPntk3Ezz0n8R4f0scg
HCOfXPe7eYF+H6YlhCNar1OVUkaOPYH+epUt+rxoh6BQx+vcrE+ybUMXSlcdiazr
e16bTfy/3bL2AkZFKX4RBQCCC/QKKr8oqefT9hqH6dwq1AvRNglKbXP8Gn2PGXLp
Uug2aVrJUG6XPU5AqiYnKdLyGZTPznOv1VQ0DeJfBetNu4Pg7913+QUecCuvh5l+
xYObHffm0emT/L5ARyLHrPTxxRv3lyKhf/9IBVjTVxW/1E5c2DCX+jsb575kyLQY
mn1X8L3AhIdDLJBMjO6Ax+tYl5ELFkTfJIT6eMh/z//qjfMcXC7105yOlc/k9xml
Ks+6a+KsXadxHRPMKPo9HGsnEcJdB78t4F8iwT+7x2A8v46XYHPhiXc9IdLpKQOk
ICFAzXU38XAfr53sw3ryY0QAIZVOyd0hztcBAg8HCWkGfDXVI27tdynUKBRkDm4Q
W8j4rT2xctdJaOt3ENeR6vSLxjxYCbRnq1T2wYHiBfDCyOeGrhnW7GAr5Ri1BWZY
qUAcMZfX09NbkskZgjpVcGlaEZviBvJUP16np0MZ2I5g0m10d6W2AUTgKhkCUVjj
BAvaVcaxDp5Y2jOvfYXHr000enoIp7WvxWzrxGFXaZQ5ksAUOz8wwKUBozSUd9Mk
ZgOULuOqDcTG5q1DbzMWWq8zxR9GABviJrz7qQVBZBqYsxYOEzRJpndyLmV9O0aP
M0RXltVNfvQP/PZuzD3BXAaqRKmWkhW61fzQawx9M8ZUVXd/7WaFckcgMHyr9oGK
YaXeJTNAZlMd51XqVw6oVvih/YSyZR+emKMCW58gVVLUgxki/9R63pOUkbXHsu74
1e6Hbejujw3ZKz+Wmfg1Xa8I0bC7/0z+oWCz5ioCsxHEL1KlEmA94S6LwI7oMUMs
1/+mgPboMSW38+GB2e2yxgDe0+Adh4os4EYb/x4PRoXNHL5UV1EtjTE/CpEhKPyU
WLup1i3ruaPLNPmd11E18qc3qluJ9PXN2uAgi23Kuv61YH9X/GTy9a2tLwtGYj/W
PLgyEJn446cAdkU9bm8ztzOUU322iJCcMsIMm3RkQCao1hh3Ra4jjlb4TjlsasP9
`protect END_PROTECTED
