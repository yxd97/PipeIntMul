`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LGCOym63nuXrx/Alp6cfui81SrRrPfrMLYDZ1kmH5ugwxasG99PcZFd3Pn4U+I6e
+yVwV0eIBZe5fnARwaeO9noYSbxxutybPlllMefGUFlUn2RMdVsN8/XQDWshr1Wc
IT5INRUUpQPUD0CG/DofcXpur4aW0U5ATa1jX9DUVMUEC6cgGTUot8kR4MGQHMIY
46Bd1CxTagwRg8iAX473Zg/sFj6Ynspne5bHdk8Z4AkQ1X43VooP8Kwvo8gm4ac4
oRsFAajNVqanu8esgn9DDz+UAU6zxLQxl/2knUkaeALrswQd0TwF18mX8DHe6JQT
`protect END_PROTECTED
