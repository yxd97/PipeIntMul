`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
krYaSMZX9crNB//ZIvyRrlCIi8nucP/qOCNrcGG0JJVWuYo/LXQbLS0Dd8qTnFXR
pB6fA4Y2gv8DxMz6Gx88Z4ClwhItOx+tJMWRggrspoh0+KYz7Cx962MzWADLM5AL
cvkKEJ50w+naDHbwEWsvW2azFnZli9ARc43Jgx5w+y1qQ8VXoz8bsmqBrhzW472A
SozWhTbBmlCSl6X/Qp+reQcF6GpAVw2Lyz+b+wXLKVbvL9CjAvH0+EEoPh+12VU0
YRIzXjK1srJwGge2uoe1REob3QdpTyW9zm/SQf/KeuoBtvZ7z85j2097y/Vve4lB
xG8NoGhwV++Npf2g0qopjJgB+P3Yb1y9s+EIMT4FFU8888rnZ3azBNM/2G2sOoeo
ayq3LEwpNdYe583r7wBhTzprmF8lasDxIH+zsSYr9VuJoHHyHKZqzjRZkJGqwsNl
AWoax9TjUEjre8Pc0tuyP5qVBDGQUP9Y1tjSuS/9IY3qCsiQo3bSIyQMPGH6p43r
aL66mlgyOFuHla9bviKvrpSOOVcJPVvCS5ny7u52TKkGLx+WBAfpxzp5P7IfPpeZ
qBQ/GDQmmDWraQBUsIpU7kyXwcmfsV9uBm/nNWBBruZANQKcqm16mbjXif5v0Klh
zu/+xI3CisUZqJtEVdT0n/62uSKWx5bJ4BRx7HJJzUyetKAUJ/mVaGqk8RrwtV1L
n5wQ7AbuhHfr6E8nPyiF8spFzKUSY1MnOyQUuEU3JznxPou2qV7W3LD5Laajnr63
dzyMlOp7RhPYvvpYTwz8oVjtC64hjfzDhvkhhutMbJzOpdLwtFnQVpEOTI0I6mh9
5Sd7ObNS/t48QQBBVIYaJjIbklyr82E5R90Dl+rlFP1OH26o2xCSMDgOYipElboc
l8vwq8Sw1JclP44Ghm30h6DY6M8PkSv6EFIbo5A/x4eyN4cmlB4DHDLWkRSXQI65
O6cvBfN8ihpCkyvhbGltXGsWVVPckFKNhlX/Jc0R7cyOnDao4wUaeo5OEHAittd6
r/hBfa+D3//jE5D9E3Wlte/DeKY+9DXt6oqR7rCSD8GPfot3/gQZsVEVd/IL4Ruc
v8OD677dh86Arm06GlpYgDeT2cpwMTnz0I7/ANvyEOfn4R9E6l4p0pkuUI5eRMHP
mE4CdLi9XF0HURAQhhm1IYRcJBx/Z1wxi30qcGSxzd5ga68JPKUIBFEEO0bDMkRR
VHaweLyR5Mblb8KX0XJDcWeT6Bd2k9YVElNM/gtEQfbDmgEQI8cXSWvFm9xGfdFI
PP3KcFzwQs8Gtqg0zz8SSSPU2/1/ktno6j96BfvhQaBiguHTCirBh4dL1tQJqWvm
NVcLNVN3+2l+LI1v0yWr7wisur2qoAf188jeiwCyEYCEpwUwpHq8Q7MADyYj1ZgU
ifQBlFFQl3l4+9zncioIjXHUjXfxC8TmKaeAnaiQ4RXrtRjzEJKO0IEctkGFKh2n
zOev9IxQkMRIY4qBrrOGBiGPE0o0hhAbRiNLS9diagoj7e6ZLndLjeT7U9lf3AaT
UYbsKeOrCLpZK1/lxwvB0HBsPcD6aMyp/JnKWqbO7wZWm4n/vU3l1ix2h7Guvocb
63OtH+nzePx+fQxhWMXViJ6zieBF+0l7VGxl1/4oSt5+QLJJEob7IZFb5hZwYaiV
w0gOK0GlD/blpcA8hMrirwLEivPVFN2E/ARIHj4bC0k=
`protect END_PROTECTED
