`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bvw5rifHTQalBme97dfQPI4jo0QmQ6L+lLaDplC1mm196irNu4BDCo4XFOakYUeA
BeEQiN4dZRu2vLfVtayjA9BnQcI+B6rkhBbLDJo4yniWnFF9Wg0KgmFoTXpJx8kI
v8TXbaNCnrlEVEHXdif+8BQ3hIGwV9S21ilQ6XPmsyMWMGUSFpHNkXh5qqpGZ6nc
fBVKs8g/+NTAoHljwtiQCg6+Hrvzblv1N+VSYrKoNLRhJfyGbq6WBCBwbUveeSvL
OS5tDzX9+OsvuiEH14klLeGN94kgrSwz5PFhQcACVeKSfxAIyXcDUU76qGGFhRye
oYLEgNTMe1VeYTcqw3I5P5CCG6YkUIWdsx5TiQ2GboHB648WSvTz00l6pZ+3s+Zf
bZwl86CBCGpk7Cco0j2BFRj9ndUlCoLSkCCuHPzUqA1cFVCxeuVU5wAUkjjyaWm1
4Zp76mjIfpZiwHBQ2t08w1DemygPrnL/bX+FOy6TDZk4WChCErVHTIcZpDqmpCg/
`protect END_PROTECTED
