`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dNZpTcF/sABk8CPter1kWYWTDuxWTZ4HwADv38wJaIS3jLe1lDbw23rGiaI4EOIZ
NvewJKyP6Lo4ZsLUtf86+hpEhTpO9m6bR5n8TlvYRT9wxhtOAnTfS2ZezCm01mxE
tE5UpvOZ7NNgeRbQgSj7k9nIpLPSpJG2Crvmjf0yW7dPagwM3I0uEIUbyYhedVE3
wutO+8+UE86hsF9S0gnuRE9ipTLyHsFSe52rugf2B7rvpzAdv5BdAFwiQMcXvhyd
uUFw2KWLRrqnpAMuej8DOqAXcPU/wvcoVPmCMfh5Jwb1MW+IjZE3VFqSVHbTodbD
HAc0oUDtho+sDFDyMnaMd2BoeTZXaaVCKiccMadp8YTdsFHfqCyz5EgRl5h3BT66
YPqqd+AgVQkBQh11qyL352/dSjjQ+Qt7rZlQotMgd3tAPMgGTesqKbNcL2D+IfAZ
d5eq+tIDFlfSubqJADlA81WNiXrhED+P31bdojszgTPeJehkaY+U3mXxFwmV16aB
VihcmSP6gNSSP071cL2KtUjMMyTwG0pAYJmXweyJa3n970w8eRyPA8NDVS1qqxL/
RU8uhd3bwoMBzXhP+upwLI7hIY1HjOjpLwtWOxiY/39qC+CKhbKtIt4d/YYGpOMT
+ziuhtYtNnxIY6UPhaFMUdx7zt9PJuK9UCC8clysJLXx5ksq/TIVV05jakIkj+G5
MWzP0Oxf7oZ2DYm3R4atqTvHzy++M+zb5D+JTXjo6n05QRhlzdgfPpBE9KiaqGE2
iibr7wNAULhJzsBDBj+K1pxqH/pvowsQqxwsjiJUtS0b5Uv04+ZrljIKb5SA0Mnl
SHpW0fjMt654pddlX7yrLEZD1k09mJUyVzWzXLFb1YWlhN5QcaF8YC0vLNfWMhwa
/u9oUTkaK/NY2LAp6fCoHdADD8mO99PS6j15UeE1BO9JDA4ntvzPDoTGwEBtiCpy
LN+C7NWkfzSKAy03YsnSvgoTaZEP9Ig7eYFdXOAskaYpjytU7fvx9dR8oaZW6kR7
k+acWMnlg0BAg4O9lVqpRo3sJyZLZ33dk2dFGMBZ+uojqznMXmHghwvEVG47K6Fs
iusRNWDDErrOS3E/7HZp9wS38ugcvTRO2Dte27YZc7NXxKNS19B/d+kh35vaNJnS
HmwbJKUzGLtYObZX529I+9fJG8fHvH9xVwhGhtzMG0Vjai0OfbuR64DmNmA4AFDf
XeO1EUEFtUv7hmwdJOPZMsS9XMxt7ING+VfGW6Cjp8CliTw4KQWZtnhQ1Yb5ORhD
OuJhi6e+vDqeYDNoBw8T0PFF2vcmoTVpuvlhqViF7d7vK0apYSyI78mhxB3Eyr/j
/Zr8t+/eGt0GtakPCIU1wWEmnK4NDTH2iEUHxXmVPt871/4iC7lSNJLKYT5O2mjk
KApq9DjKOjACQTY6rRVI3ent7MS2qKqSFRnSw2uR9z+58Lmrv9CBTrY3rGmJcb/c
dnO7veSaQ2ZHaf7ZrZaGxxlpRocRR0ASbY54QQjEBBU9HblWR+wfBQiizKJIO1bq
V7Sp2lYI72K/aPThhT4Qm4MWy98jvBzLs9hStBD6NQhhDzFqsi03fDm39Psi3ndt
iemPI1VkqAkLeGYI8vhhMEz7MzI9W4v1To+2y0MQ8v19vZtedd0knc72W4PORvf1
Y0rLIQBpoXyWHM2ip/hBj+Or8gQRLueYjekzUC1HzVfdSSrcq5czqyZozIzvUgHT
Zs5WG40Wj8PIijGdVwtUSzcTNKM+U0pTPet9F8UUjvYcMK5bmUKzlIlHnq4gzs8d
B1rO1fIz7n5KUrUblYur/PTH1vMM/ro0WvpYAlstak+mdB8ymPMVP+V6yBoq/zHT
UIw/0CV6KN0Osy1LYNNSR4glleQkgDLfBFxOStxShmk3FWtUE6tq6XgTLmlQTIkj
i6zjRzFqOQsHRA2/Ul94nW9P+RNeh+wn0LcySqaGYtNMoIlAmXu7bQjLygAtsHpP
aCpI/R1qnpBe3DAKLxyEXWFFtRVF2bVQh4F2yzJz52qnzCD6p4qKvlhZjM1ziDk5
Rela8MYkjF2/4Ixlk7e5Rfzg5c9uqR6FtppOlmga99nzIvBQuM/wqPdlQpgMnIuK
Stsm8UWBSCCwa18rLStNHOcp09bXFGv+kIu8kNKIaZ0/11z2WuJAxuIn9VkH+PX7
GpWPYA6QMfZR4E0XEMF0bHsFQRX98vJUHNnCnN/chiAa8TVzXao/obKHQDPWORZP
Fn07RJnum+OuLwqg3nlsnAUK3dCJhszR2O5lmoT8fP0UrMvT0YzopwrhLCr6h9im
UVZa0+HVZJk5iA3bvZ8m/2BkyEprlfFHReH23sSmDsEvETuBuC3SkCSm4CFL+zlY
FOk+LfUhsIojEv3PNUNTQY2BgckM33p5xu3KNgf1zlLQLYb5G9hafa5mrWKGuYZa
PiXhRrhbB7w/lvxzCHJwETj1oSu9890otEq3tq6kfWnLl8T3PoCR0WEoACSTYAt3
c/xweYymwWsVE6CxJBggrqQHq7pHsNxmV+WklP+tT306juNn4Dt2oqGfPFnGZaTN
xsK4cncflBPIvlNeJk/4dS57fANd5AxN4RpSuBUwEPZyZgoEYi+2LAu+FqtGvVaT
AChxEvAXdJNwelTgK9I+xJNyJZvWgzUeEIQwaUZDgDNskGhQX8hyxfdcwHBOVDTS
EvVJlPlHKRRbBlS6O7XNJcdkjBxbAiw78TYJS1qlFR15jjK4rDhgRjnyJfywWoeg
SlpM94fYEb+0fGEdiQIaxE3/VUNaPR6BaODfPIU5wJrP2A9ydEc/BfxpuJ+SvcIS
ZDV5E0hHtbm3wBKP2FJ9P0nXiZgSNeiovkaRqsHPhfUTPR7xbplTwImNMUVELkDv
Z7LhtQbAJjNryzxJpxMqPQ/ufqvJxO3d7ugdjYZwQ/q9JzbZzhQu7i/NMIIjPnZP
84w83E0+9828ZI4kdoXKZ8x6SxSFzXG4gMsnZO2n+/APi42Ojj+5sHTRpCiiK3yc
Wh/oq1akTfewsozx4g4ftjKkEEO7RdS6xq5amRyYd/576jvN25OvBB9Jp1hFD2sf
z14czIIWupaIzjdDASRYew7lnBGxBmPa4bHDPl7zXeFjr2dIRnjXIJjdXbJbji7c
LK1oiwfvRtsoLUczhRcHjU0F6gw4/E890nRFEiaglxI5C1X8CusF6VXeEUWfrJtF
/DHyf0OoxjS5Ypes0wfZ2orhqewr30zfFa+XJ+fnMGSK8GA/oP97CWe3nBVv+tez
SLl4czcHrN2xbvfpHPf0+6C1h93y89Kfe2Zs/r1PUI90QozBFbhYrXjO+JXT+H4V
DnfvL4mt3O1LgKmS9dOdhNQsV6ZimLHUJNovibiM8ebtCK1yvsLalJRSSs7hrPzo
W/xCsN+TBAfiBAWh34W4Yxcie2pOuUKl++360cuuDwsSkWQsy1gFdOK8VUvn9BC5
T4PsEjFwDO6FliLcfWMF2Q+lFMBzRVRz6Qr3Nc1Ovkst+KCUrEj9ItVzifNSu0gV
WV6LxkEiqPUxFCXMCW2swdssVc465gajty2JLaSf4Qy1sAc3084X+KSWPIQXsPxT
TnHJ4MxKQwbQY/p4dJE075GmGkz6Er/ZjzlNFIOsLvCNYUjGbyhPH8AAjGaixtGU
LxlBjjPu4Q+1kf5k2GxbvYJwLEBPUk0i8VhBSoxTlGA8zhPSoxLl/UeiM2PUQuBP
RhflgkknM6Sxc1NEyXVEexfIH+boeQA8oPdQLcsAREeJyzvcHRF8k4wsYGB20mUV
6CoL+mptBu9JX1BrtGZL5+6WwCeelGb/0RKBVpjdyWXLW490lpAC42WMOS5TCVOK
Ow1qig5j4sNDQu+JtBNNxcdg08umXgAW7X2zGBgZk7Il4Bd5ix1rmPDnlHg+ldF5
Zkc5niuYBhaQfVVYbO0ZK6bgssah32mxyjs1vfYUKeYzO4ViveSg9lxH4l9aNoyq
htXLePURnsagokC59P23FrxXK3cyKmtW/K3mdSVsYm80wJ2LNEL2YkIbJnSk/Tby
XsbKUbwmwuxRc9S46PUBqwETRPCEPkv22YKfaCQdNqIQV7bW247UMJtU1smgkaC3
gPRxEvbz+ra5KMelCen3kvQy3FvUtyscIDfIj5PGQ91p9BQjdZPap4x9yIyNjPuU
XtKZOV8PaxHX2VD0LXFe9iFv02b0RItN6s8EutQKZpw+DhTWLV3eRPiSdndFuneA
9aaW2pOGNED8QYCFKzMZCu05NPlNJ2LkgO6+8jsx+LcOMjzV4DFI9nazfugtvat6
imUxFn8Wr9BpbXze+pnfXCVYPTI302mesiu3MvmH30FmNWUiIhQKh7i49yd0jaIZ
FtliBWMna8uihlP/6EQNkEZpxjHXXUoFbtZ5jiHP3c4sFOLv62/LOWfbXpLfYjcV
rknOoiBa2+o632nBQui+rOLFeTGe9L0AEcW6VwN9ahbvCGG0pCfNZrzafBlK8RpG
Yx4a9eN19AQ/GH9wHL4GLiODsGiANqicrGBTxnpEjzE5HRAcQoWO2FtCU6Yx6ikG
A5W65Sir5fREqqKyYd/dC6jRBbym69Lw7TMrOETCW5UCK15q+vlLSm6366i/5mZO
ns4y2HbMUwLmXqvlytKhqNaZ3xeabqfpfPdj9s1NgsV29tdhdfhj2D92SWbxLeme
TyVNtgO3/wPnz3aQPpFe8ow7MszM9YeuGjUtDlSQYqJsVb8PjKpdbb/2k6B/L4OB
DDYUjSSUtmlQD0zstkxT1nVL+MZCBYZLLUhy1CqokxNY56PHIdg3cUHuDsn0+VNJ
RJruFYgaLCZyZYcaClm+1UthJY75KNCLT+/Zaprb4YmWs7/Z+d7KqZtFCuhcyyWo
Zfoqq+er2PM7ZF/Kmr4SeWJb7m51Zal3Kja5Uw2brT67Dgs0D3s98jMVvTUte+Os
JVgZVqlAF+UvacMpDd4If/zEisgdsYm5D4yXjqNNxsCIF+AWEcHVOZIevEtCHd5c
IWM3HkLHUBF0nzUQ9+KbWo5VpaqU2v8NbuG1cvYje+MK2yyb1lLG+9+quug6fy4H
fJs3Y99w8cSDpQ1B2AK2OAFB46P/l7UW4moT4JWc4FvEmljYGIABYbfy4v0RJjyE
XC7Vdrm0cm+WXwVN5l4Qwt/0Z3Sb5d6QYP8RhiFETkFpuTpwFjw/Bp3e26KBEDlM
m7OE2i0N6PHU2Xqj023LNZtEnllwdH0cc0nbzAhenFeEEfdJQdlNAd9/s6Qd//OM
32wKnmxzKDrch9Bz44VHcsIHRzsdRP6sbC62tCgBdnJG22RrdSVGAR128vMdVVBG
jQM4fd7fVdmxV9YnMwBB2zXKSWeucwYdmmw658xjWj89QbcZIx/hV57DJPiNZfFA
QqFGB1U4IxgploIHU3VeYezVLr6M+whpfx6zZtCnAP46PpZCmhOrY0x1HgVUPe90
ouxcssluoAP4SwNU+u+A/fn09yPYxSUyt0d6kZM42hjN7HfXO1Vr2PuG6XW0xAD3
PKM2knoHZi4eNl+eJdLntcsvgR7/djw/skoGcPgzJXVFSTzJ44cc8wfmDXm0a0kT
U3UmpR798upqOic8YJYz+793FQablAbnz3VNGxHZLSBDQM78/HG8UjO+rnyizJ7D
JyOdyuoScm97yXDn8B6MxQCHQCI9u6tdOUxkP8s40sOeEsPXlkgrefDMCf9rKDBI
QeWSZTrd/keuSAC0m7VFCg2dOdpXePIduw8fuIhcuDk4Xrj197NZK/Pyd12L8bUw
cMzuVzhhf4rJmRryKCIUvj7/56fLOMwgGsExjDH9riM+4GvLJiTDGc9SvxuYghd7
JM8ry/s2I7To81HPQVYToefeMQ2LbgIUM9PRb8C4NNP/M8Y1n0bLjO7BrAnz7uTI
aCkQ1IvKch7Ef+sIwXo0Qj6vRhEVMMpqJGL0fdGvEuOtqKFPdDa880bW/oSUxIBY
iU+wRh2NPe5dqW62vl9msj2GzMmp5nOdXTMsktbG8gh/XTRnDmYaVdzGQCj1K/Hx
74tladrAT7PTzFfMFJiacpKERO446cYqrW2ohfzrj1Y79NdBF5Rv+Q9KOs3iDFzw
nR6eJNj0bAVkBUWUOiKI7GWDZKP3VwwfTlgHM0FhkeYQ+/IPtotpv6iDmD7xoaRr
LMf7koIKNdRTxgVPA0Ing4QAb7p9S2B3zVPqh/w4w3f/bxGGpz9eiIm2ax1wT4fN
v0A1giKN4V1hrj4ahuC98gMrea6V2CvJm0WSgFpIDBF1zz6camAVZom9i6isIcon
hB9TTHJkiuJ5j0ZT39O4NiLmPyBdZ3XwFX/OlGt8vskGOOriUvCzLGVb6X2EwadC
1UvtCnV2kk3QnYEJ05DtUye40n05OojEz+cMkRpMMV5/cBi/D8080mXNNqkWc1OS
jiRx7t3+XMu63tebP5dmy0HqoTz+x2yWKq2Pwnap0EtQSqJ5rWDyY+bPagrzrdZf
E2G6QMbeg3hISeRG9qb+SOlDzEws1SL7d4Yv4Sz/PPIAEJaP/N4wb4UjOZYZO7y/
bvcbqkVfPkk9YZSPKjmnGH4M2nRuz6LjWKGrRCKbEe9T51ZDktOLscyRRO6tzeA5
zPkyCXahZDISQzkqrmCVt0R87iTGYg990JXPjopCrxnJlO9RRUILPBgTPT0/LCpx
sylmroQcmYOFqpmJIh27cpuYibflHxQshpVSrq1W7Pr/+7mgAQ2pKNhMs2lMKw6M
+15C2D9Ll1kXxhx5ZjY8qck0yyZjf/rMQvqsVR/GGRMNuPbU9/AYcEfHE73penpc
d4QUUe1RhEfhIPc0iQMV1TYUz3B3azwnDYEC6q+NYH0P683riiBnc9wX8rMvYsna
BcWkwjsT9yFiuXSi0gfFy+nb6twTgIXeYH4CYxlDg5XY9hd4BeVfVqudM79TlFX7
4tr3P6EquQIlBDa8/5NicoXQhxv5FZkr8Q4UxB0inc+hwZemM3sBGs/bQm5L5ITJ
WJ3NRSFM8f0bnPojLhkOTzN8+u0cd7UDvMXghGjGt7772jA8GbgaqnjPkLfrcnrK
F9yG93kR6InoHNepGRahTSlw3nnmCod1KrgxHYB4QhAHzBjjvgI6rvQ2bXJux2mJ
rj2E1DTSxwkNVL0PdC32Jl1whb5pyHqL/pqjPWEDAx7IM+IAuznBRTDeP5rw9dmG
U1k2iuCnQTHKX2OGHh586JLvcvTPIpWPPjo1aXSzuV7aOnkcWDuMeRljUvimpvCk
+2hsJ0x37KZFU3yePE5Udk+FkGLIticW7Z7tNupxrGcLJKs0T6a1kkqNUW3c+bqX
MWDHlTJIZMU7A2ipmY4L81jVJNyrdrQNw5wW5HfJAcRPKAu388EWMSB7ntcTLR2d
vTuT0PeTHSXpMEjrWpnHCkfA1IlqGvjnufzdIhSisNpBwTHZ0aikoHDZXZaNxjs4
yF2HG1XfMjIGNh4alasEmK5de4GLeM5fKylMWNkhfzN2r+JA2fz9LH+B0fFBlO7e
42LM9ML/6mRLy6o0f0DO9wWAcGPzIdQeEwnng1zxgqKLZl0N/73Yg+Ccw7/ur6gf
lQTTSfQZgSVMKIgRuamQmasl5njT/DPT6jf6iJoA1YDL1uE2RwEgupgHB3dP3OsH
boNs8Ci/5cOTqUq9GqNqQseOgs9R4Zs56GEAhgovovv0ZEtPa3VTwNs+lE6qd8MM
S0UY/SlFgec19X6F3353iuDDPj7r4x8hE8eJxcExneUjEAh9ixSVVJXIWBp7qGew
9cXfXW5Ll5bor5e4hSL+qkQnsJG0/hTYHDJrDzqvXlCPS0xnoOONsX2qV+qFum38
sYCzB15YWFKZDlRj6F/zgNLz988khD/B9FyrLLiviA6imJbDVJFRQlKvFc64+EDg
e1BMDQuUIzPgq/HK5GDhYOlIiNB0Rw4Zu9lT5GiMz3U5MJ7PaYUeu/51iXHTSHGh
7mV6UbKfsnFl2RDJ65WRQc0YpPkS2T5CL2mGG/RPEmxG64A2itYDcxySbdPjVByD
1Aev+Oxp+73kud0BVDIcFmb1vu8kRccMVEMfpFbb5RZSEr6rpjqED7TTWve85sjN
Uv9TXXXvzZ5EJLdibZruGR4frvarcB7rrbQCSQUTCTukdv0rsOmHtpLSz5Y2EYX7
uywFlJRPoKbz2BQnd/6qQJ44rxJ0mgXxdgGO0C4zVt+vY39AwXJibRAhrLJDv4T8
IiPgbrOPVMWBlqmGbgBlA691tGGLlTa+83KkotQEtiISGJrMZEATMbg8ABK/bpx9
pRx+tBbCbe/i1Rvk8e/aAYU607dVWDljqF1AfQ/7IR5U2+0WRA2qjhA9YrLS9PhF
q2HVxiyzyVfTF7EE5jzm7/fjzeQhVZdxZDLMzvfuhPP4g87tyykXfpWNxcak6+6w
GNwsTFPuNz5Jd11eadFkNJ9XJfQutCbeHjgFyD1Ahf6BIPJ4LG7KeIljLpOxN8me
brXeLFOzP/6AfyMS1iVxyq/MMzNpezYzZdA3skSmWTsmPCpxGgPn41HOLdAhbXtP
eSsA0Eq3yTP+GZ5e/dz1ObvjqutV7iBC3i6+EkEi2DoGXVXachEjMledXoZUf/5f
parC7uME4gd+9XZ6WvP4odN6vSgo6SnsAIdwiCfaBqygo2J+NzinN1fNF7kObuSP
YwMLCCCBlcBNal9alj6FTwM2xc2dM51fVP/OX4BPpLUQtZ/702LIZYsLlE+JdDRw
DaiqChXXKj7qUkuKjfth6wZjgEx/OmCo7AsnBUbMvlbZK4k6ZgFT3xY3HrqIlW0q
tHsW03ZAURqfD8s3T9I3h4oP+mLC4eXaaHlf/bAgXgWUL8ITfOp0kVxwFXfBM3VZ
TH0XAyxQQBXHrbikmjFtcV0LHy1OnsbnXBDNYbs/9+pnIGK451WvCJsZCSi2k0ZI
6/0apbBPzoOqz01t+7gbSouD9dtP1zuDQdCKAiZOa1Qpgfi6GCkJ2gizKRgpKzTs
Q30W47GJHVNmlRFJIc6h2MX0Ugl6+xwpCfHsoY/ewjXSwffOnT1JXSFN8PkcctcE
g7m1XHZ8Op73gu9yWjN+88qkBm3gFGetr3Cw/46fjeM+RNDY+YlN0Ll+XW/YacwQ
tCLyqEXWoWCrvYrApIK0oy6VBz8exM4ubHemYzvAVwP2RMTiyPGXLEloKTOXpjtc
iIgqCTM+vawxEScsA22QRHzHYBPzbsYWVeZnfIMUSMgqThX9H5oBk4or1xI+zksv
nT3T2loxF1NIIEdjUtTVCylmhngQch2VaZR2lt8neo6x5x6SDHDoRTu2N8U4ymKv
KmbmxBR7pPdomiGGId2Gjkv/YNx4Jw8fMiM5A/6SGXBqkkHmSnoBlcbzVS2eW0uP
zMqeiXDCVZJM+JSVNLUvOYJ+TvuGE3PGsvT0wka8/BZzTnKjcnAoqEnsxQa8doyt
qBj3wYUkdPygTeWhgTLUfhH7dtLD7m6EDxtFPBrRXhuBhS2UyZthfnG6QOMH4s8s
xsLbOmmKqtqQF0PniLW1xX6LvgqNr1ZmLlol6S55Yo0LGJVV8CQkG7GRuORekmg7
74Z7meBgKDmXy9pXiwdBryMwkMNg83CrBecBk9338pPetwoOl+8QIjgmJk9Xjuya
7Ltw7rPG4I+K2EsoUlOP7Fr+AAE+ZE0vneZIAcBmszQp/5WOkvYAvu4kxOoM+bUJ
rAu8tlvXWOYC+h7rXA6y4/XUa9jFLQj2JQSFFy3gHhDCqtMElSbwwPmxh1LrEz4P
3mgWJXmgimmfzwgpmhnJf1hY46L0qzvYNlytOJbpFmB/MslfV2mTucGZ/a/MzZKm
47LeJhcrDVMQ/k70sM9XcmmAEsJPjwQ7uva3uuhasym4MgAXGCM0tAhHsOY3L9sG
Cb33LO8ripxRvYxCXuaFCCtf+pThhGWfRPFpVwKmlR5RoY3GvwtsN8Gmn5urw4t1
nCP8aKW/glqwofTQHEP4BFkACgYLPBw7vfW6aO9GQJ7n7L3haem/yvj3CsIpKM3l
MkS3XLQlXLA5RsALR9B0HqBEnxr+Na/TXIxdvrPmri94gMmAtoS2H0DNhU94Uasj
iYxW6C1L4YAMzW2tGcSS8BQCOSvn2MKl5fxoRdntwzuNg2zjqq2gu8LMBk85XZRF
A4HKrHjaZ+BfjBqeP31ygb1gJO++6Ik1M5rqki6zXxLJ0rg3W9RaFoPEAH3vlYNE
IPx42IxN8TLPGrYHk09OUGzSAQcDfYIQ7vAQbjTFEmTr3sL0shtvlcI6IBMhkJO1
iHeWle4RUV0ToLGTVJhKhY82zw2Sg8seV9wvWYY6Wi6DQVBw/zFhpvfThgAvvUYd
hcTAg/N/TuYqsZGRP0+Lf0ondRW6UWhQeKJZRZaktLvdYCweYl9IGdAsexHLG5Dp
bA0Ma8J+NPOrqwuxOBLaSbRp+Yv6V7PGGBRcI4Qs8G4sI5FPEmt0tvkLiRi564os
YSYYNceugPLGy7CJheR922uGoVGev0U8sChT/dUzoYFmaF+sh1wsjzCUerlvoPHR
6/ahnsDo9yFM4KcvInHh4H2uOwK2R4qg2jUzfgBLrgqKzgquM+oXVPgOIwL26h0z
M3ItLA1/+RhJ8WMguqXMDwNWf9P70IKQE7NRCgOX3Yry8JycT++VBWTE5SzSBdaC
+ZYE7KD355ZcYN0zHKlvNW1loo5nv3qRHkBygdK/0K6/xKOCgSX5Da7KdmMSr5Bn
JifarCn7eD7DVS9QnElLP2kJ9z/i44JewPNVXkS0TvdFa7Nu8G2JiDrqjwojHH7k
6H1ha+7jobezcoXalR8hCf7LAILHxRsXPCmEq3sDd8ESVVmaN2JSWiiLO2rdX6T5
lxo/v4KhXHce4WBDyP/YE8932EYsIr/AmvPKKpwMcNlTlnPeb4dxsW3A2kjUQ+tg
4nZx/guoGwWmuCbKKh1EZnl2a/qOwYJxH8o2RBlZMJlNYJ+fnxrB6ivg/7EiCEHu
9ntJ6YOehyZd1tjJYOtIwjlCt4ZJi7511qDwdcZUSzHRFu7KNizIKFSEIFAl+n+F
NptATraLgfBf3mkhs+m3E01vbVmKyzAjIbqIGQtvEfLkqnKF96YCx7vnds+uQXCw
2RlHUipmggo3UjjpbzySczaoFB/2Q2umvYHlpqENEefLEDMJxTs1Zu88y37LblYD
BA6Y1sFyVoEYXepUvn+KxK50v/x0F6jJj8DMTysM2xpxITznZkIXxEf3At7xG124
UrqdidRbtuSxTVCoRcbv+Yq2Dgxc40n7pU6cndrD+qIymWz4Q3S8gFOQgT2KiCti
gpGAl0Agew2ZV+srwu+jnazDpsBULZMSFyarrh4kHrX/vKFy/aP/9XRZcp4wQBU6
2SYLAOTYuGJUnSKorRdoP01x6jvGbmA57Tx9P5ogoWDs0LwQ/2PD5kdyukSqGGYj
DQ3nZ0RkAkoC8j5rYQX7b89L0r5naI4XDgu2RvvtLzCp0fkCiBmo3W4TOOHP/WXw
MfCCKC1kV3Ma8g40Oj43sGZxmbvTL/dez/MHmMCgHf7+WBcSGDS/NIOp2KtdAsu4
mJ47/I7ImLH3ekrfrMooYNJS3N26scrH1n5G3QA3+2VBcC0vQbyOQ9JOg9a0SYBc
x65LTVx79bjz4glzhnzG7N17oq3iwgwkYugxwqjluOByFmZeBaJ83+WH9A78wQLN
BymPfYXpxwwUqLlayzDWXz+4tndeyBnwj7xHIL5ygzRYJcLXu940BxUjRhmZr8cM
ic1B8dbhq/eiI1w1AKoUcmWhMir0QwuSX//JM28uEu3ovlXRGEcH7+yqBeoiyC+u
a7d/Y5H3YZID9Tx6C4UDtd4e1XPbi9mFvbUtlj0hp4HR26l2/QIzD1YYTq1NSoRo
zHhYfCHf6R5z4BkJVfq/WVVEXaBOK8u16pcRJAATKdM0oiVUTrK2twIVyZED+LrD
jjRhbV8dBeyyEWroUkjrNuBlBpkjSc91AYckKHLQeWca5/y84pfNbFfJavbhB1zM
TaHQ3uFNdTmtKSBiyQ8xme1vL3w8JGP9W0rl4S203rZSIMI3RbQofOJmeWNHb8xm
dIDus1lPev/pM2IpAhO3vDZzfnD1GqpOf9Oab5zcxf9K95HLNi9jhYB2zUaVhBP5
RHxnQ2xQAiBL9rX9XbZaBhA3W6SJfxk4OHyeOjGIlOh1PVAwZ/WZ9AtgNOYPd02F
oV80KiW6Y/0AnHwMIFgLvGkTWAGycagepJo3px2Aw6MxYnUkQOyMduWIZim4fkvR
j8dWuZBy1eCxncUb2DBoAYrdGtXKRWa2B23x9gDU/lfrSir+ecVj5m2a5lq3c+9w
iqPFCT43h8O9bKQqFR9LQRWeU/tan0Z0ffbgWE+yxE0TQgnDrb9jx6+QnqEioNUP
WaXhwa36PrJvcoZDyBmvT39HId8/OeHXZxW7FUKx7TW0uJ5kk0OwGoVtw3SPX6hD
l7RX6ZkI5DBK+euQLzH9r6BdkHkMtMQM9d4X+HondRnY3MOJJibLx7T8PiaIOC8O
nUPAgiOSfhnHUrxNUjK7qClcOkKN2GVgDVW4spwE9/o3LU92MukD+fZr6vjAfh/1
I98vEhbG8KYbFOS4RfsbkXY9PILWms1Pw7fmujC+lQnWGB2ex4mnBtjRyvyGMNgq
h1a49w10avhR6hsy/w1Eu75WkygQ4rmGejZjT2Cmu7XALGvsm2KcbdBdxxgaTjDj
jEvn6mKtqFozAiD3IjN4M2ua4TKS7ujoUFOddTAh1dPBBsq5iQ1tyWp5Vsunuc4J
fHhcnkqIKC2OWJP/eywzuTfR8kZgxCb4YaWOktjD9Z1/I7e+yxPUsolmeT6p2LsT
0UGfE0ByRd6A+73xVeHVZUhx6zBwhtDOniYu5/qVIwULzhfkTnera7YcKm4XtpNX
nSjaNhu7qV+sWnHPdT1/OgHdb2yVWW3EIr9UzzZxU6BO+XcPdxoT4l6LTimOxAax
zSVI29axU47T+YE+ifZNsX56pPUuYBCF8J3Xv4sqa4XhuGlLYYFRCHW2Q2rTy1b0
ld7IY0WnrXEYSVy9BZWpPmjMHGmV8PtJwqYiEnMI+GZnbihsTZ3dh1dqGXtL3+Gs
urWXGLfo/r7GxzP/fxc15t/B2dKMtY4lWy9UaV8QDsrUFIc4Cznxm4gBAPkkXM8i
6wkgGwIZ6ixu10tVUgGjldY0G+jtLcF+35zWQ4Kmso867SDTrAGmsDWadOanZe8A
q6NyWRX7/Vvbm+W2vU+9Ic2OSLXlfbuxO9K8ywfiejI+jVpXf5ZKiiMNRPbE/fjk
HIhpKkCMm7v0y/SbcnaaWcGyIrKvpXdpchZGxIQiKlH6yxcth0z3ccHk1Zh6YUpm
knUa5nt0oG3tCu6hjexP5wEY8DHIHRPvnLU2RY4eDMCa9XvEWuOX19OGyftwCB6t
I1/ARCsXSWBqICdpD52t4xgarPEkvK9B+ZntECyreWVI1aHlZ3NiZzpKWKbgoUCT
tN3d4pnRSFm+HGDwAAIvSwBIjyNvGEPieA7Vt/SeoUmZbFzN71cjcGoabPrBEVt6
BUhMrmLKjnhecIXOSAnQ9HFFcbmJqHKeqamMMJSDm+ZM3GNG/sW6YyvhOwSc37xj
SwzKnJZedHX11sIuGOKuPOz+7cvDXG8HHmo/tVtLsaaw2teRYE75g0A7xctXdKWj
G0lM7xLAV5+vCa44x5sHJ6jgfUeYfhOjM/Tw0QApNAAe1QmoL+qDF0krQUvfaCfy
yQz33l+2InItrKxvVPltxDBWkbzoig2VC4V2qN6o/JzCneYkb9i8cN98lPxwEQS5
P+oqI4BpH5Es7JuK70sqDM4I75PTHjHystCNBB0Km5l7T3/8Ls3VlNl8AOfJQMt1
qgrk4ZGiSBx7cBa6DlmgyEur2+y3oon/ENMOjakiSoURrcYDWQBlHjXcwUWa5JqG
/la5NtlsQhIRi2pJN86BINPcY+XY7r47JjUXJoZ5yxJx57jtgxjoD5vd5znZkwQf
83s9Ibom3b0TKSjCHLgNEN5EHhNZ320XcmK6ri2xIS2BHhrRC8N4WVkENCAeRw6W
dJ5XECZ6VG8xEaEMVyCNBJ/KVJfs5v9tkwfmKL+Y5lZvI8UImxgs1kQyL1B1WLHT
Xj4QyA6bMHk0817z6PfIPc0tJdhRktQa5bE9oUvLxizZrE+ZGBMtVl+V59GbMlz8
tCNPK1Qml/IojDs4mq4E7uDZ59jTwFa3Wd6dDkAekbBFZ165vK3qO/KFnOxIAWae
jjbEvcGobZO0cfqFQwTFVGKebb5ghQc0b+w5HRIEcZPgQd49TRLBqCYh9ytHnNe8
U9a/Fw+CqUVfyvY7tVUczsoWmfBvbUy4Igc+qjB32g1hCozWGP5KwcIXVK4wchPx
ZNayFV3ABd5CMedPHP1S+eXp39ZqE9hCpEYQdnVLQmsJ32WjWr9UPmS/no5nFxHj
LHk6A8Lt2Pi6iHFF7+sGOfprSLxlLiH1A4yc0LtNsoWXnatr4jgK1+cSfFb/Pxoe
KRbdYYpmp5KbiNQox702sENs78MpRLsPv+6iTSbKFNF7RyNUjnt8mxLNinE9nc7n
PnypTgkgJ+drsWpRejMZ16LY5XjBOTLvTRhOPk/NGV3gcbz4yHaHvuel/1YZ/Aqb
stbNztc2BTaEi4LiKYXZWtgqbl7evmKspgkHh/9ESb0vHbHU3/n1JbUM90Toofyj
aLuAjGaGyLCPpMCf9YrsdiXNw4E5DFNZfHd/s7RjKNg4SWGtHldgwxw8aXM5Pp13
gHIomG6rESh8SpSNhlbmPXlThxUmXf2Zi/StvV5VVBPd+z45S951m0Gc8biNJJ2J
o3MTpi2md6LhfwjTaUrY0d9qzRZcOz/9fwcrQEaUAPBef5Fe7gDvdEJRo/0ebu+m
+fYbxgSkNTn1vgeMfEtD35ZEiIguEyeVfI/w2rjQWhhizniUoWqtyFMR1XzlrOGf
OtgeP4SVCx/m2ATQYmxgMo0QwBrtQxp3RBd2mxEpGPufXitiKp7XAZj4cpEjMZ43
UHUuPhHBjrwM7N3xbD1z1FRMo+Gao34DkAGyDm490iTPgyFJSyEA6HJrVShQw48J
a5NRy7xBqLBuHubxFjx4P0NkfrdcTnFfrWi4ClfeNx0mgWa7XSmaKwtQRFJR8ouq
GasRZR7VaoLc9uaMWxneenwonckayFE4tUZ4HT1bLJjfvQN4NrMg/2ORxdA1773k
TGoLSRDtJpMZMusIV1oBq0GDNQJGj29ywYQtO+k2gHUd7DOrmqiqVDt5XmJGegnQ
B8LG1atwB7YVDE+KdV5QijSUnyIzW8hW517S9k1uDeXJuWpj/KrVEPCMu6o4Uksa
cUMP76OMNAI3FjWlyFDMni5FHkpYgxwQXTGfHNVh3tmgpG1pmD3vPzJawxGCfS0w
Id3bf7uxf5Q2RKnE5xTlMJKwHxdyANUPZKZvOhjWiSzF21GIfqKTgSVQeOhNaK4E
9pIc7sDl6xlh0f1KG5U2wjDHkQSScayulOapDVUxwmKewqsDeRbLA4yZXDor4YuU
fxMIHZfj++kxbM3rH0NfcUYDbsQGsKJO7PMZ/ieEw2LeZPOSA0vT02FN+tR45xJc
hRMKoXvjJgz9HlGlrR4M/mOtVBAT85u7zNPfPDB1oW3ZafxUCuNmS9SSDqK7APZx
p8fAA24Xhu9hKvjQ0LFb4xLHON1jBUwap8nc1f6vb36ylkrA4jsBYHAl9dkASIHU
mtMTrvjR1moH23yVa+FYFEa0wevpmeZVwWGy5p4+cmqikxyZdZR3L/ASZ4dMRCZe
dXMOWEKu9oPYR2LBHd/Y6lfrZt+i4VyIaLSIpA4At+A+EoFqBnJgH/pSjMH6psmm
JWB5d70qngbG4g8E1eztPr4cBhdJtHrsOl7qT8KVkYHiBbgMgJ0fkOxO0GwsEjxQ
iI9LXWV6avqZiVFqegP+ZttvT1v0REKkyPvdBFUCljnwxYzWw1qGimxNlRi9tHv/
7cpG5X1GBSmEdAIOH2ovDGeCKacsFHT02+2k4411EJMFOWcf9zHNxfHfvyYYvt4Z
nUfkppocaZ4Roic+ObDAvlLmO4URpnVBUI7R0TFNuQlfdlVas2uyfLj6Tr5K/gFT
oJ5mCz9cSf5YVAdZQsiv0sxpxZ8nvmpbbKHN7//1zlRJpdMmMlnzHs5IYNKkYcQ/
holEcIrUTp4ZPD2Gb3n1JeUpLqiUPpoE/JUx+paB3PnAO7DNoo5O2Ww8d1/C7b7S
GY3tzFyPj1CYP+AVOCLw/XGFyM9Hstp6skJ/16K+MsQ2jTPr8knCRZe7sAnjatyc
zSHDcSjP1AaLF/Bv+mcJTVXNSdaldgtfWZKaxo+arQOf0IpUukkYnxFvf24hFyrm
9qo3fIWqwVBxXgJrFDPizA5QrzVCF32sxlWkvNo49tW+qb4rKEV/73TlQ5nTO1ut
xbsuCVjbuAhn6duJedVRV7VWKxPom+m2tWYQeUr7tWBztw5AoUYtFhirOF1llcOX
Q79TyuImY+XpXJSzXRmtOt2WuRwcDCfpWLhEIfbMBetKSlFyoe6MRJk4wgjjka3x
u/DEvYxq9rEdvm8A8rrgujNcGIUqXBKKh2TwlcB8S05wb84+TwMZ2VoqojWqcgds
GwZrTvmnS5Xif56bUHI06odeNo7uZUPNVtgZ1ziQTNVUbHTFaXdP2kgbOuoa18BC
wB7ThNfwKM+yWJ3Ncyrm2kgyBKRh0EMbRzd8Ttu0lKeZDIYcit9hG0FKNhU7lIZk
OcNPsmXl70BmpYzenJcao5wS5P4IAIMesn+v18//WJu6ehkR5xljOmcalJqNfUGg
1fX9tjk7QgnunMqeuGGC0B9nE42Nu/djT2x7IYEya0uhgez1tnPFuXSG1K10E56G
cYFm4x3Earw82TaRbc1BrxEDtEQdRhB5B2MFrxAYfeE50CLURZv6nr2H8vVmI4Ea
kFoNFbZ1t3LGvcS5Jmvc95hekS0N3u5ZqvEAfJusOE8OScQB2rnHNSU1wSl7K1ov
cEs/yCiyWQ3BSC0anl+LnXzJdfUyiwjN4kRmx3ZGLKSWT/KN1/ZLS2pUp/GS/lzx
1oM9yW6z132NeuEuVupkoY7dYeGGQuc7I9kH21I/HuSpWqZY6z45LOsKgwEZ7UcR
MGWlFrAou7BA3XMP/2AI3/27ZsCkkXVwJFMXIitfD7QaOaFmTIYPwpIsSXQ2pQ5x
7Xy+vaY+bORBXjhiwNCLQVENLeN+Nt4xqOOTufWJAFt4V5f8E33zO5eegjZjfzad
lZUNxgOjRadBF8oE9NIxgFMfGvsoWgWuMimgId76tI/VAnZXeTUmaMLEl+XjTEI2
tjsJNYwvR4wssO4xijhteLfPnGrQvJrXNPGN0TMaXuaryF/gN2lq8OIqhz9foJ5F
6aBc+n4A5IUOf63ztOE5HJlIUo/Mi0msYVUkEJQj6dB/7C9lAmrfFxsw16Hl6Noc
vUynh6DleNBN3RNtQaXSQW8TBdSJChW3vcNDi/WPGpEGkSpKg7liRiDNdfPHukSL
mQ1hu9Xgo1zwfi+jj7LwzxItI/EOQyj+q9l3rCXEY6OhqBdxfYsYj4PiL8Wo9xYm
4ICtoNfhO19DSGxoybpjWxU/idZanFqKuWllA5jYCIF7iUiiiS/W/4YxOCGRKjlB
EAshypBoi7zTwpOJqwWdYQMBFbHq2bqsvRp7mM+EtWhCLLkFKDWy+Ny4cK5IQveR
k2zHgBkk02Y8TAU1fe5iAz/dANi8C67s6vhnGxUWkGb+qWgPs9Ty3SOEf7fUdHdn
md04E8aFPLg5Co2cGPN/JVhpa+GlhFINvLBwnHt6j+GWu4TEyxG638akyxrIJXfU
NquVsOTcdk6JXNPLtrA6g9SoehoNvh7L1c2yxTcC4L+XzORBmiDqQUsk/ob6DOQ0
hHVNAH9TKJbdLuaHd2AyHwnSTdnl1/Kjw3d47T0us+HfqN1LumkXUg+gwq/wvuc1
RAJZVeEU3/ZKaLM0sJg96uwfhTArO10nCeGWxtISDgiMx+mWsP0iqKP+USjEgq1m
X2AcPjEPTh/ipaHhNXI1y6JXAEBIsOYUpVcL+w/tJZKDshe0SIJ4vTLkaKLYpmtv
G3NtzaPSxvphqBsroR1XvfuRdRbaKyw9tRj+RIKHRuTQQfhFEnylHq9AeZP3LCvE
2Wdej0nGVX1MU8TnQZFGeV6aIHlgU9JtfEjApjnh8gx8AiLxGGYoLQirmBI/uwK3
BlRrOWu2eMQyvDgxPK8FekRsf/m3c1c5G0Yc0UXldxQEEkhMoHr3dCJEILvbcEwS
hEjg0PTtOT58bAvyH/GOjdltOkkuWjQQXxjX1tkgeWx4j618BybHfvZVNE5HorJP
tRTqG/8Mv58pBA9aLoM0e0ZUd8g3k7olK6lPmatDrHWZFpm3fypqWeYf6NeIt8o/
X988nb/4CuvPCDYpGLztTdf5QYsYy5xjEAQ7LSrZUKk/Rc7LoPHcFb66iZuVyvpv
F4bNG8gUrhlUrF2aEsGHquey3OdevadkKgw2pyo0Fjvxy07NNmFCBYAlRlMb12bn
MCbhEwRj0hWP3n0WSMRUwUwZQ//LfK9gfIvSUW64VQLDvFsniV1Yr0v+0WAw/jhW
6C38muICyEsUDKJfWVnyB0QTW5P0PsmBJ5HZJvkPyidSuRT0ObUhtvxI3ye0yywd
nfa94xMwsO+BguVARlSX7MK8i9CefAcwPpe3HRATl9zCUC1fZPcIzOv3kgI3mqaV
kbtoOB48frSvSs3Jgu3hOL68dM7rgHHG2PWfo+Gju15zXhiL5dnfRmmCZTMUFCZn
9ofvPRl50k+PoKr3bWcs0uGfiIpyvmKO8oQcRCCIBLEQ6C3fVdIMkyu17YS0sAfJ
xbqxuEsxuq6l/alle4c+hDZxq0mBkeuBQrFnPnLWmHMrcB+Kz/9W+vQ8VUEN4bGI
+zUKfIGvfwkvOYy0pMViHP/qxor8UfjRT1+QeigAI8uY/JuZVIMKz++z9qXYQ0Gb
mQDuHiWXquO9QNbPVVaSf9GPiT7wKhKsGspDbrqHHih7xtqVpSEifF7k4M4pUihP
XqUJWEr1yc0cSLhj9GqIjvP35bKqrIcxlz+s15XfPY0xB3NcNIhseCERvjC0buzS
Dqm/sVe12x4WwNYrw26ctcBTGWfwVG3NPhnFMde/zUZ06LBqqPYPNr2M+5saYkJV
qERCv/aeRvTrpxYzfB8owOyFWxe/nT95rQZosEpZ6WR8aN66RYzADR9KajFEWgmS
rrQznnoJx+uGIXDBkzPaPL1O4er4Q+2a+cAjr3BmitzFFc29DQHIj6TMqPcGKwpj
+7pldmCSkIdOhD2bLM4icTd1Md+cUMccQDV5JQVO1HOvFMsetTRVAv/355kaOIWy
XW9kEHVeS8DGH+nSxjC9NcLuopMCe9+7/DiDJNbgZa8EoAyByZFsqghg63dSrieC
OCxdxQG9t/2u1ocJcSV3BjWFIIk+s5AvXLt05grJpS1HxXC9U6VBhTluR8nqrvtG
HHOLAWjiUuo5plkbWHVFay8XDqT0Cjqokxxl1aTCBEAMxudQwXvE6LtzwMdfnOV8
NxlXPxrP3NW2Gm9+Btu2F4YDbb82/lbDdJ5wYIq8acepIKeeMUBH4rGVkhTJTtq4
iVmAp18aV7GSC15JIGGbm0bYFplX0SS1BVHLPhW7kUw1gfnjsuIVThls6uk6eLq5
ZTzvbAkHfOk8mK2gyNmEhFiEom4wt6OujW9B25MBz5Wznrf+FSNDh9awC4aiwhV/
Y4w2vxCyyUPjZGFZ3KOQJFlJfYpshZ+DJ6hyz69zti6AApLwrovytQVlqqtu6n9P
hZGwh7T92gN33NM+qAF39VttsAMXOMng7LiTeYKS5994C/wWKCwssyWxn4cM9qjB
dcJUpzgcEdac5pch/i9mrcOm51somk6wbV46Qw15oqPjUlPMqptnAdii2O+cXHkT
BqR86sAOuY+FseE45Ft/Vhs4SSoQYHNJIYVOACoe01OBWj4kLU+IkqKcpDc1+h7y
s16l3XZ1E4XGZw/BVXlxNs8h7wYVRXYpaKCFQElZFlr/hVBmwLZIOhmAfXkbkSZG
3NttR5qEM1Kb6ge3v3f617iX7lDzlTmuG1FNoGpFCS5ngFGNK6tIwywOG7Q6lJmV
rzHScYVe+RXs6euD5LSV7NJ8pCc56jmVGWmhhgx2d7WuJYTNW9xJTnNlrUueYeOZ
WGNUMskwlYOdxvuVRBG1Q8fa0ZMBy1DIN2olIGtNbqM5eRnXUa7JVtSylJDwNKMt
9lhYN+Vs4/a2kh6syV+LHvD25UNyEMn/A9xkgODyXXRZLcxFAH9uXHmerY8jU5R1
CLWimAwuXLSwSgrkuOalu6lIW9hGM1VvAf+GnvMBH10YdmDzpUCXok5aRJIOylar
ZNNCIqZKfitHA7BHQBhomsgZmRo13uTmpAZ0t+QTctju1m1MIAktNK1+Cp0aQpJC
vd7rxs7oBEI+HpEDmJqgzxRa3XXZ7N2i9RaWc3ygo49lTYDJYCGu1GhKa7esvwtc
+9bQTkH7ylcLAYy4WJQqZTOqvi+TDfZZpAKBddsH+z3IHQwEPemgq11qILnaxmeZ
yq5Jp/6qsR4In2u6hEY7eUf6XbvcleZnlJDnp43TqrnDlDVZU8XEv3or8wH4IthF
xChJLtLIzBbecfnxkXY4QSeNEkmp+wXzMhfrwut49TcomNQD6AcRshEqGMn9Z8/y
hfZ4vodiqw6tgAO7SVpW4vi/n1AzN0qq3Ahub8e1IZg2hbnqshvv9O+TK046VHZk
2OhEPVMFSYK6n4Uzy2uErEAyFcXmdGIJqQ9HFMQgEMmn7c8egmFtzdRFuPDBfOty
RxJwcR3M88g9Tkb6eJBqoCFCiA1o5AEz3ZWKaneCaTUM+P7PtyyA36G37su5sdLV
D8Yxvynvd50KVcWcSd48Z7QqRHe7wLR0ivacxRGu7UfrPo48R+qJvMuyutBunt63
he6z+01DxL/LWG1Vf3OlNFz/Tw0/XlbBg/PPvC4TWs87GMpmDwP1K+gNTsJsw99s
bPxU+tNUUbfODHEMaExlBE+zn996NssGJFxhchYtfmVLck19FwRuTXnAF7MSNxu2
WSz0D+9AUNKi0nEIP3/LPnElmgNbNi6AtYiRhmE2OB4WVghvAdAE78Bm21Gy0WBD
NuLl0lJM61lJEhKoTuBnSgSxxG5IMY+XbEUdhrh9N5WW9yoijYV/X4Fwev3EZuRk
SmHNTkQLL3YIHBx/Z6e0A9N6e/m9kKLBlYSzBzKLNBFxcSldVzF6DkQQwogBMBhK
8i06E3oKVo7ZX7L6rVP2BaOl9iKvDl6pJmZ/JbPg8MOhMLY3vYemgGtbHb5hYsIE
sGdr9dtNyuUm7l/xnrZY0TcHE2P9w0qkP5u8qIiWimxvNwD5kvhnJOhDgamRmhYP
6xa44ChZOKXVRrOMOOvKUpxE4aqrv9fWUz5O30miaAVCS41X5CrzplyRr1mGP7FX
zuaqINZ2jIiItXUeoP72T9BaHgn44ZzFWyqVMg3IGEp3jUzIUW2Dn/w2o//bdpi7
wAjNbJOaGwnDxvOu+4D2YHBBk9UCA2ceV6byOapMUBszn4K87JXoieLJXks3K5i+
6jOm9U6xeG8Li/jVxuVfQ+DLI99BPygJ/cPT2umdmrDA5nvOWNKHhL50/KLtB0Qs
VsA4CEosDQTAwVdOLvU63UOkLOjacr/SyegBEfgnZpXS/MtN1f+Duqnk6/OjdzPL
3L+DDX9sYxxRXn5yNG7Z+PrPuE51DYokENozZbouhL59vV78hPgU0Aj6D1qsL+Kh
EdXyukHJXMcOPLISqUVAy5y5a4oiUZurhGnjiY6YMss//cyWzZr6/RYk34+yDI/i
jSy3Zd9QV1gH7Qvuc2todyA4pQ9Kipqj18k5YUaIuq75J7kghLovMgq6mpNXPbqA
DQDPr7w3w5+Ib25mehftHuuUaafzGLlnPvwXcOHBeqQD6Br8e+mJnyyYygbF9ize
1xyLT3jP9IHJ1yKpr2QASapjAfGO/9mumcO+MljUZQOQgOOgC4QLoCXlgEZjJoEk
97UGyEdIW9Y3pXrhdwK/N/vQLPO6gvW2o4IFoZzQtuQVNM+0UR+KKOfmnuzdoJMb
Q1t1oevGmSWPg0SKOeYCtmwXWBKezCPwZB3XyZhnOvcA8I0ZBd4bMbhC6LYF9Pgq
2GSDVoqcDbna9btlze/xBdG7Sn0RTFIrcio6RS4hIS/gkWH6r95vdAabejMYMLqy
9rhSMYgB+mDjXlvUVtAbx077+8s8etar/IZx1+KHVEtJ6tXzXVL+APv9iN2dJVds
gnicRb9JwsaUiUrA+6h+KkqlSVu34w+d0W4hqtB/VcqGTB+fETlp7xEFM5Cpj6MZ
bkIWrvrqsjbu9UOTzxPYCMWbPZJUVu0OorXiVfF1aUAP9ne5XWt/thjezVPNSK0Q
BEEeJ2ak3e208+MHkUnf2uaQF0VOqhpmQGeew1Lr+deTeVnIrEJW7kjySyQCITrh
YxxI40Z0gdWFIaaKfPtTS97f3wptJ2x5HeUxuyH8dcmFpl2VQvVTiNUk312LoR+U
B2y3LyHHZWSMu1mpFRiPyxi690RLSwbBSLTBVUaTpyk7bWqJhqpL6S5RQZmD8Ae2
fQ3Y0B9hEikOCyVdBjpFtgTRnrZYcSoOxrkg1N4603LEkUQsViQ/mZgInwpNTS3p
pdGTmhGY74S+NK18owzntBHIs5fHUZzHrYTzpCZdY5WiPMMLlSQuIWXjOQw0vvXc
enlerMCwg6iYIzgzLpYmg0xSdlqIBZKifDQKy+8KtbufOG4vXy4WTwOrubaKUzDw
Uv6Yp9QQbBLDNfYalKoExCePs9M16wDSt4xPpOJPcVRVL1Bk8CVe7OG0fVGSFGKH
WbKbhcOco7XVw4AElN/m8a6rSzCsVOzxhnE6Cb2ZLK0Ijn/8ZyIic3wvHGBdC3qT
4HGyUF4+j81eRJpIC01xZLsdZwQN62UQ/5WEkGfgSuYY0ifACqo1lyeMdEmgYTaz
g++K4l8gvjv0Od2Hi+0jm9CwhaK/FLlL8/hxo0cKpDSeOgAoQajrLBrmAa28wAjO
E9b6sLOASSp3QUA6CvywQV55njpRgrKCHr2k3eESlBOb178gH3FWhau6EvFg5dNi
3+Jfr+rsEV3jFNI2nfmin1N+lHyk3odBR8gGMKu1Bj0mRTTAIxNayxLX4coHYrkf
qVrwjqmqzEZi+rvP7ik3My/rHM3vdp90JeWeevSbCm0lkQEf8psKyxC/0SHcM5t8
AsMONB0yA895wXpO9R7GU3CH/ZvEZ8ddY5ulWqwOWuJvoduChXOGJQsxfJu18xXA
CwA5pEaKb4oKUBdcjfzcX73NuwzTx+f7/fD9ACYDIGemitB0vKyrjPnKgHXk/XyJ
Aux38g8wLq46GkGTzgreJkc5r7N23//+ZwyrscCNh6/iR4tEqeyzI5fA2Ql2c9pc
zAwpmJPxOaK/e3TKOj4EeF0lU4edLp5kW4k2LneG7rTCpXU+F5V1Qi8SyMTQ+G+m
bxLf3gH++4n31Mua6EuO2DedzEu1kl3FOU632gBCKmR8Kl/shMr7wXpSUajNvJKr
o6HEcaGEmYyVhqKnlrb4nVctzN6dXRDbtjnLHxHi7AeXuGbGz/zLkY5/RY75mMJd
jrNdpSP7My8A209CcdqBnYe2iftJYOTTd1E7EXrJzW4izZkDRJZC/CdTeNaYqBZP
PPQ21IWCm35ALmGXJTnkqS6Q8wb+yPwwmNIvPSZxSq5Bywaof2cH4R0rFWBa37Wl
HmXNEAGdfDJGhLWS8eanVmV6AHdPCiDjvxlU+4wubKorXmC2yV7Us83N1pNeRaQC
udphrMil/ytBVpQB+3EDEBIkBVn2t8KWTsX4Lu02HP3CofGyU7PwoSOmr2RYaQqT
2gKQlBnqCPu9f/Ise9KV0TzErj6LZW3M5Y/ntXlTsLQjnIasUtYTsL6tJMCuWjmX
zOtF6Reu/LmDdO4NJ/Np/h2NlOk5W+BKEHwA2EYx8jz3QEi1cLXGrdqDxv4EAwOu
h1E0+6Qi7ZrdcNDdSX1oHR8m6MJqYF5dd0uKSBDnUR+o+yhlR8YP6jxvzWcwvU4d
S42aky0EVpYn0zvQxr1fvO+1VJ8yerMhK3+ucrhtkq+AxvNpRCog4J02kxTq5+qH
5+ZmLCyyeiZdNQ6pwG5gvrcqvep/Mtjd9rgnYldc8wcDILcJk+2uve1Rvb8b2RZ/
lidbVWIDb8ejgXxje3h7vcqDNElTwCaD2wRHDzfJjiIohMIaqLQ9xi3b6T1lAlp1
fizPFsQj+PyF2WlaaKJo6m5vg5XNIjnA6tld/iYmJiFm+mJLMSswl38x2dmH/ydT
Le23ZdMyFzeXdliWAUql/slYjncNzga3rT1HP+8YEEAL1bO2kBzBZ79QSojC/my7
W330VS7vyx4uehER1h0ePg0pdmBbNX5ApP3/+/FzShclWuZ0orVnZ1iODMRcXLdl
L+cssTevBIeS1qW1LshYW8d3NJXBEK8a66pmiYxewWM/vxTo0ymBh2kjOTSCnYDx
M57EZUDw7SNpMu2HXKpA0XWG4q0I55qzmxjiGkQ9VOu71SOAV5ggnQhIuOWcVrPb
QuYfOmNSRDHKzw8DGbpHDfmpSu1wZyVMFoWfMdfgANCiTUWyR8eU5MbQjAnaKWLQ
NlplWLibHZwg9tubVs4+EYaxCxU6psNq58h8dZywtr0kvqjVfoJyfL2ZLevrrHxe
zhDzFBqKCDUORhoe+uJUmVC23u6CuKJnDvlJ07kETC+4ct+9AYzAwVHiWb8SSMjm
2IxmbAa2Qs7gDKZ2F6Mu+zv310PIZNBLhcdvo/LGyyCgLvC38ZBQnnx4s76Y+Mhw
wnD87vqA7ctHBWrQvUuoAJWimWHo0DVRdNWN6olMfSel10arKzlkACnPA6BsbBha
TTYsddTRhAg6+VdcsucyxvKFaKZxf6FZNZQIQA6tL/kt2RDQyaLcq7g5zFGI1iV9
lvvJbeIupHfIlO4CRjBBbbz4B7ZC6Ua+rhI/5iUBZocxR0tPIjQR8LjOCb/2N/tm
Lq/X3DRCeN+KAwsYeMq3m6D1UHvwfSpAHG0StFvJWyrzxhRUBFFM45gZ/Le4cSsK
y4sAjdLkG81mnnYSZR0gi5bzNWvO0TuJ0tbL7Xp4eAHMLMEzx/jvdbqcd+b/7aEV
N8G6vg5MB88DHxiXWdxfTi42c2nGYlue5E5o0zwbivYPk6nj8C+hrPBe9eX/Sk7g
4S67p8LVQwx4D5WZxJvBJIs9eZZ3qbg9ZWUzDQTUTxm6Qhltss8iNuz+Q2HXL7bS
qvTn6JtAzjGa8RrgVsuF7uW1+ZGFsHOJ0vhuYsBGXWwZl/Dy/fKbe22WrDYwD/BH
xj0MpdEVITIhZI5k6qPbrG1QZ9w/AZ0jaeUK3L8PfSAN1heaUjypI52mYcDNWE+m
zh0D9eowz9fpPmsPU/r83E7BZp1eTmCKZETe/5xrViSaEeBzTqoELEyJctnwe1/l
bKkYaHFt+ru590xwj4Kx+OdsyyCg6XgDO9tQ1aaLvLesUr33SaKvA2gNDgFdudGJ
N1BvsNJImvwlbyhT1EKX1jCSDOr9GR8GlNX/UYtd5bF2ijq1RtwsCgnaL27+lprQ
q9J5LqwcVIGkTFYV6SyF6YuJlN3xIkz6d2UIn7IiWxRlb0zT+qy1DoEHojA62HSZ
aMdnF/ip5/HSftuDNUGAVl6HXWROUbw3F8KP3ald4I2nZBV7iBTPrPqsR8+jxVId
rmV74YyhvCBkszI5QL1iVfldKMTPJgzUILeCbhxolGRp0JqDgOQKmEsQU1Td3pfw
myl5qICuNY6F9RZXSqFNI/9q0S7ttH0s7FWpVD6SVmKH9NQa0alDnQUrmOHRSAFA
DzzBmVg38y6nxKHhTutWzCgFLaTN8oK4GeLddFdFFCWlc1SF8Ol6qDowKfDek1IV
IGCa3awky65/nmnPS6U/aYhvL3HRgy4a0M9G41xLUsC4M1nYv8tJZHgCzygOiewR
wYcSLYDGsYnUCxsyI5FQsG5IEYE+OlOi4+1WYsURsJ81cyKs6OJ1GB7hlrW1f+4V
kOB5d4UKXxDraiiG2R08TAsjgk9r9SkFfjxb6Ja7a/AEg6lHlKi4nwKj6X6jIAhm
coMg0l/0IMRJUjWW0JiMHdksNm77qOci7Y9s5WqNGnw69ZkcuKszRa1HDnOMK26S
wSquxrh808dFI4Lv8KcY36iCQb9r7TC4vqMSyzygLhy4De2u8AV+qZhMlsPiSFJo
DQgd4peuhQXu6YoTXwqTt3rEPwANi0JsaKfxnuomZDBpTU8+3whXj516oAA2wYjO
Scg/kKYTmKhiljnXNn67Q0DvrbvwMIqFkAQrsq6dQ8pygfhID0ZaXn81trEyO6Nr
zM0S0aETJVPn6dU9LFxE2p8tEPWnX4UY5eCtCOf2iYadBnMdmzpV6a1nFKrHtRRL
3DiYQRzY11b1Z9joCzpJjuwHIPO/TvSgBBHEbzQCVMaMWN4BoebUMCMI1Q05yjvV
YqbVKAo1Vwycy21FBrEHo1EqQMwjw290zxMjKQ7m4QuvI7lnxqzlkU7uAJGq9zXv
E7HXG+gBbgRDrpi+HTuan2QvAH7hlATAjiqTIhnSmZpPCTfDD5luNayHIllPFvLE
1B4eGLL0Cm5RQdbNj/FqWnSpRsA0XBuN/TSf6xKkn1Wi/TlQzarEPlaUuh62c8q7
eNToQfa2NVO9JiGaxlM8KvNoj63u93NtxZvVT/WZVjL4ngSVy7QAYSHabtHgPmAu
KB1nVrEwk75kdv0vG6x1gWLprbK9nSVArnz740a95uEDUuNiXSaHmXOJX1AeWRqy
3uOoz8ateXi29WkOSVyKMldIIVij4eQaxLE3jA6qo4saXbc7aiRY3WuDTAp4o78w
/sjigliT8C4pqXcKZK5ShDiFTZLhQK6cUfhrSoR5LxOIeSYAsrYTkZi7YROWaCTs
cxf8aDBMZVCsiW0I9/RzBSWnafquvg50mTPLLb+U8nmg5tnMEJaFxmQVVtY140a5
ruB+ge+PY0mEJk/Pc7d3+xS88+zNDYd6ts7E9JcFvRnzXwwMNJsrXau20gPQ/fGf
f1JXkaABCud3JdQWIincFhu9hNDF5Z0Ny+a+rJjdsgGPikdf24puMbAsbH2WZB/m
sJp5zud4jHD46babkX85UeS9j/b7BwewOncbACkWWB5l08xEFuF4tDNc9sBsg0aM
ms4CCZbOp6CX6na9LFFT6DQ3P0nXTrdwn/RN6nOCEYaDVMTMd2/1bgn8+AxoLunH
kGDxdjw94zhL9aue2RP0QClMe8AhIaSOvvFM4ESzg9uTa3EgoNc3Bs7pfjdQ124A
LQU0VG4h7iw2NtqKSCRj4AAuK4xVf+6wwBKygVhSDV8nscX976AKFc3PDP+nVnqS
D0AsROp7H1I/qqQ+VRkCoEXgX7m5XjM29BC840yHAvzFqJBl/gdBGYzEaQ9Nk8Rs
9eox2Uev5zhvW8Oantde3WeTJZNpiSTdSMm1mhyYOkmQas7h/EpdnSPKuApR+hOB
eHmElo8+LQE/6je/CopZZlh1sLPGu44gISfGnwWjjXly65TlZsydDgkiS2WIQerN
xnZ1/NipdiPmFm30Y97VdWs6slIGJxa9M4xVUP9G8xVnASE0FQuSNU8pXj0OqPP1
vnyjt80ZkRUw/UCHEVATR2wrJIWvomVjcKvm9ngyP+xlbs3Loixs+4zm02TxVZ7G
vlojYqdWC6uVjsOd3OQPdJgsjVQ+Zrd24xGC2UIApvsoKJzvM80MEyWH2ryFdlxQ
SHQxisv0JuFQRKJecvIFM+ONkr47/UVSGUPvcI2EbO9nnf90ol7KSuZlHolKLJrS
n+r7aJ4fms/aGnnQYIz1PDhHVL+vy4QuH7NxvpPZ/1fW4FoqTz+8eUk2qB5EOpuj
Hcf8e/vD3BrgqW+PePtGXzBYfotql3G3sRobDGZOgyHLWRU+1tLndbHf+94d8f/T
baRnvd1iC4JHxK2RdKG5xhsxoJNaGiIlVwGC+gbPpMMBYjvAd7iTMxv2ybjqen80
Rbgdu/2LyYehJFMGGWsP80TCUbmjdVQFIWUyejSBMhJc3OaM8wiODVMl+hm7i0kl
bEiz2FH+TC1gEduFfxbNzIlxl3S9lJzKKT7ix4JNiXnuy4Kh3i2LfxtcqAyb7xRd
hGLaKHslmgQ5hfarVMEI1QKPvtbrDAtbjNpcJ28gFj18tKfUjXRnMhAr9+D2wrrc
xjjVnpV2jeM3mHQrD+i8gnr2/8tsvwEjwKJbtGUAd9/wkbXpMV3j1GO5CMkrBtul
AWV929UJ+SifafwKNkfXKtXgPtjlB/UXG0DIg3w4H7QeJNnGHSTmigLsPY4MOPwx
PJqgTU7MjHMhfMX03ut25oWcmj7ZKFp34jThj9Y4Qgn1YPiF9QhRUYn5KKx2XwHs
T0h0N4VkpsYQYrrWaANSp1P+kA50TiWJ2B7/KN4FeuBVYb7q2pzsaBki1K9Z+Cbs
/pboC9f31MGZreBSKa0lLr+a+4unzIIHxMwIHmvDIVIjPoxY/cl18SetT3tDx3Lj
pbI4g6/yBxUTQbzFxoNzTTzLFiKmLsnTH5Wwg9u+YhKsLylZhOHroiSGJgR2kbvL
xNhCtrTeqdqk1UamPCVPSLEtpyza3drmCa63N/5TkZMMhRV0IYxJxsVptpw9kT02
cFqpEpG3Q3yRdqjRmcn7R7JKM8VfAoA+a0iLkkKb5u5vExS6PefMIYTxMWU9yb6q
Gl1HYS8siqf4LQCwxMZDdaJ9OR3c6WvjFCru7w7ieF9JHurwtpd8W+uZrzVTS2pd
hKd9DK69LT4kmbv5+oiQmXffpUfn1OuiW7DI7rxM87Qdcj4GcraPrUH8x52H7S/B
oTb2SC0CWO4UDO8NACP4xNwBHf1tJJ5vZCgcieksV29a/jQm0mDwKvm6aXwYP7Ne
48sq6zIxNQsXuywOa57PasrHfdJILVMXTyAO09/+odFp2iqOmuqUzaJaoMCbPRsI
PpcnUlPBLAiynNXtC9YQVpEsgfn8PQqybxzGZvAA8uhwo1aW0H5uG/x2eDs8DezT
6bf+Q6zSp7P8tkxG2bMJzoEHVXKh8PtBBseYr2ds/JCEoXvXrqPxHsLIcpnTC9L5
t8Nz5B8shIyOey57CDHjgNQCHW0MVPRkm6xwvtnBbUXtjmNf0wUOdLz1dYUsYFeM
m/0nmfNwCBvsYmZCIqCUWwcu216W/Sh9dAduYtaBDIfYvOXA2iqjQGflEqM3vPyB
aqmuk8m7DgwG/NxV00ir0OQ9heOYotHfz2cNmKWKP407orU+6wiJMf6RIRv9EBSR
/h3f9jbrhyNjlcoyMXmUlETBG9PkPUqBYWiBdNpLt2coktVnUDBgGKkwKJ0nW/8R
b+CTK7bz4vHJO2Z1KzxA0iKsGtVjCA0fW4F72JbwN+bSS7OxJKPtc3BFM46xV2YF
xMP6F8M7SfCEMtMNGMGNe0M0l96+3vVp9TJPWg2lizjsafTK65ASl5tRHn4hjuRE
yr/adxUtCMBa1FvxHHMPGveiZ3MoBQL0LpDLhiYQc822CW737cUO3JDK8oGubkCD
/VrxeXUwuFXqPMRntxYG6uKi291sV50Q/b/guF4LNfiZNMlf7SoC2L2m6sxYXo59
tM5ho6Der4pF1z4l07D6c8j5YuS99JNVJgugcIRihJiRHk1Wv86+l4Aohz7/N6y9
4CuPiM+/pVTRYQt3EfxiylZPZKxfcG3bLKd/YmWwgl9UW8ahlagJDkP8WdJEyOtL
hSsa81GYVDpsuBvKLJIvc7zrLtj0QrdMSfFv54ycLz0ucxPR6qdtbVP4LnexR6Di
KLyfc6z0oHYDfJIHRxI+ZcgSnd9vY2aMH7SKBE2WWDElqQl/gckLYR3Lx9hs2mnw
VTHCt6lTcJgDgBSLByslwRKf6fQtcTGzS6BqGYdLEX1yU5SBe1E/Mec4+VHFbuYe
Ij6ZwdqMYZgEqTWxhtuuebDNEmC1y3NQkBTTM9jDh3l+S97L6MzdVvJPFJ31Zj6A
YLJdWrTOKUN0soR+D72eAgKZQNtO9yqTbQtcRKhYSj2FjeKyJM5Zb22VmmluoOON
/RLgllc+wYwr3BXFlNyGZGqid9gJkyBCdmNzKhoPvVnCRufCr8YeWDoaHJoKYio8
l5NSa1bmXtnHLy8UDEkeHQA6twrhkiBcpsR0Z3FExBoq5ub12zbRFCOQAAyX674Y
PSzpoI+SAF86HxgkC3aFVHR+j4WwZe7Y4K/MbXAXutla75kdIrijwj0XZkDvgzu6
j7vmTbuRL6v93rDfaC3paLnnVTLAZSMFi2hNCQlICb4uy5Ls4vyVGSEELRrrwPsH
M3a2Xq2qSaPf7j3jnp7tkBe3HlWWD5cWlYkv3c8HQ0wVG/psf7x1rZt+Y0F9WBC4
AZgAlLX7f2ICSa9tFy4T04TaqoIgTpDc3ELQX8e75Ai/u2jG7koOGOjtVjg4akez
At8OQSRmoGCvWImiycO/qHw30OodOLgxZwMhaTQm7IPjZF8qQxBUu42d+niyZw8o
hD4JlPl9SDAnOS94iApL43plW/7esuhCWwKOE0QR5h/ugPH+1Z/+b4XWGDzwPDRh
A+pdJI5xh8vaH9qMIa1eTfDr/AEx142GPiC1yn5cjwhC4atuckekdVfRewcottlV
TsAWLnIQ4zZZK1A5VWFsRoHYFdIIoFIQcB9lViumjPhBlgtlz50QSN+jV9zcCP2/
uohKbvmeLf3l4GHgLL8A/FC1XfH8wLsiRveoewSFj3L6EzZ0NoTlap3waIZerAvP
QW4xVYw8GC1Mf1PrUFFEx48opEDA0HUSSPknflxAQIX7VEK/T7rFOFs8XG2v9GUQ
LUwhHdJLIEWjEUpvm/Cukoj9yftnV4EVtzqIJoveS3gBZi23ENLsshwdWymfpSZH
llIMEh2ZKiTKwlSsUyVKJJSrjuVWgu6Hkp2m3+ArI65h6G2UrUqoIv+FIkq78TZt
wHfFEBUUw4S+NTj2PYqjtB8ib37i34/tatwsgllhOULyBrWQBLBXGkT5PKpYpEHg
FrzFNOhb4ZP0p+pl97Ypp4wt8ERuVSdHkGyEtz5CvhIlIJhwENW2AONw/vcPm76T
/AOIS8WLVjorcqwuGVn1nkw9ZCzhHXpjoLvQwBzZ3HhGaIkgcmNR4qBshdoFzYRD
9W5HO31ylIbWZm9Ud2iCURcUxklR405NtIQ6WmH5tkPsN/CqwT3sepdK1Adumhsm
kPFKpP/Ld6rCj2Q8ctM+zQ3NGDZtGfdmrk7iO6V9MXkp3hKDkTq2XXL9OjFOa07K
7pWEabkmKZWTXavtDFBjIsfsvcKzlarLMD/JGm9fs9VSZqFa/sFw+wZ/4/S2wL+z
+zwxTATaGKNdy091lZsOYVnEQR2jpdQf4fBvzQrwZUb0i/0LYYUYrE9qCcEWcfDD
GLPMzSHX8kPjUgZPyR/le0l0bvp6iKR3a/WWR/09RlOIvXdFqJWgvzaDWNvs+HZr
zebnN86c1z6aa1nbfJP38q2/viuxxV5zjLVTZ51P3VWm/24kvMzmxr67pUP/EjA0
n+QSEtmVfQCTShZ9tXsndQg6XS8eotIjwG3cHEZL+sA1R8TaEHUSTgabqCGQbSb2
/EYqRdmqr+ssqFT982XsfKqErHT6xvP+fp8N2Xb3Uh64nZEKQ90SROs7BHvlM4P7
NUtN6o3/k/EG4D9E43HDWiwJVt0AS76HC3/L3f1WzSq2gNXFv3pLWoWzfuEJ6n7k
2z6Ar3elBNMcBsCFHNL4Qcy++3HXBXr4Ug3NmCQrvs+WVlMNOGaTnGriLBECFjKu
r4/vUccPvdP2l9+LQEqMmpQvFF3xPfhnrMpREoOXfbEi8pEk6Fhp3ZfJnjIZn7Ag
DbOGfo9wJAcJ5ejhpThO+pZ/SB08LLqHxUhRuZ9lrjs5Wpx+zaFYBO15o/PixiSR
UvDz6juoQm08u+IJh/O6FXvSm/d34Fc/chgguG8JrJ1+7KVak3D7jx1frAufMGPn
DrCDtiImaT3VsvRkKhwfd7HLwcBDgU1rrSbYFFPj0l61/JJ//am1fpl0BGGdbjLt
2QjIsag87f2H30WQKYXcRsq9lAT8WqimEdXUyOuytfNfe+7JpeK9VelmmUFllv5f
VWVpEbvAs+3CCj4jUTYFbJnZ6WC3LVcAbalabFRQspOTWWBbPBCtoVD91SDRSSFB
cXUpOds/iXaGbW9Hn58QcrmznWNsoiBp1eU7TWxXeoKaVzCfKUCw7RdP9YBLxK/6
o6/1/Oa09T/UrYM3vkO3Msg1B/QPi/YTG7rjnIXvoXlSDBaYxUxZANIM5ujjvTcq
MyKEHHwedrWQvL7PbjD6C2IfjyKmskTCone4X3qPI8yw4sph5kvtoS50nfU1j11S
6A3wrjVXKsPx6Hi2xd+iTOWUX93g42mkt8TJY86awiv4CVaLhQMBnTimu86TkyeB
BqABT/gLU2wUUld4CCSybGy4zDR2qkJxUDlIMPpS8+82atqjFkD6enYch17VNi8L
wt9YoZRtkL4hVv4PCLIBFVcEdjYQpaIqI010oZfXdVluDJIwbYbqgILYYBIdoqi9
5DKDHDutIZ0UlbWTSZAtjbFx2zGy1HMASxqqn2/ovC2COgi+8mUocXQtTkwg5wqi
AxGoWKmn2XwZJnJuxQV2OkPCCB2IfFvL5fuzmA7FX3CWQXblbcDNdC+yCVhAdRTQ
6oDBtV6Ccijfx6109dj4+dmwZsD5QSpNeuPmuZgKFwWCKC/a6Pe6b9aHxVuKoEhg
Ix+9wMf588egoftB73EJ9k6xjppoYzCTNcPFQmttmBxJiBjajNPnuqhSjrhKdaWd
BoIGx6MSsQVtE6bGARzPqaS1IJrxRhwljyZt+XwfofmuU3h6MHTR8nHcodpADtAm
AocaFkqGmaBeW6rCcPjeGM51nl9Mgm3J7U+n2ja9tXaaXg4rYUQgwad4+nSmWv8P
7abtTDCqdm8uFnqc0UdGoiSR26mEy/KxYLXf3xoLrH/1BxNT7EnWElsyifJAgML0
NbeqAH+61D6lDEmnaMTO3R80WLV0wxqSs5GRtrIfNHZPqIyXJos/l5civO4cZTpn
OAPlR6cy9e9oXOfR3Vy4v1yThwBPWvsAKhqOyHgPk0h2cgNmn+emqsVX5b0L/aCf
lE85aNkneo45xZ1D/SWBAGMOXEt50c9xHtzKimrtLezTmZNnfW737XfyMQaLDent
mo4bMHVbZH1z+/sxDvDc6qlcTF00VP3CEITKiIA12u0i+wkRVg47ZpuzeXi4+NiC
a4doltWFX4dhWXuUBFi+nVl1clVnhrhI0PxOW5yIcVecsrkwvCNvrsESmS+R9OFf
if+25FLmIJYJwUQInPpS/N/dKAx0yyATdwnZVOkTk9aYS5hvqDPr7XIJ7mXiKx2W
JkSvmxJJefvl4EpLxTRu9rFtlyS2oPS8Onwc3Q5WFOdkUvMzHFUmjjjUY02Ll647
pyY22kp1FCOzwe8fcQo0Zqt4qa+LOfyrr4aKAhkiiFw08aXkaZE2Sb5tRK3mNH19
pES1wU9TbnUHuWUXHgAQ4n+RiRWX9IJ+Zedeo+sk/DkZ9jbGjC75UWgW5AdrN7Ch
q5nfIL8LhgZAQX1Nv9kcdx8o7D+HgiZgfJYpGMC1M0vRWqcqqUDnbwTOWhYTYY13
QQmLAWIzi8YVDa0iWo4ni1ZxBRoofBJObfbTkasiWFBBt3Ud/zioV7Hn6SA1MpMM
gRvUCAlgp6ApPx/EJ8pidTKOxuiNjSWFNfq9mBMeuX3SxFP3mjB1l84iymcrkXxI
HpS9JtN7AwId3+Mxar4E+bGrA4byWL7DCGj+HWyo8NJsi5Vi8O1XhSUQCavFjqVA
raboJlHqKj2xFshqhXMZlhfguzCVQ416xIq6+m9W7kd370fbdEZu375DAt9BJWZl
hvrZtndpkBZ8+ZRDC5nZbfjkwgbv3Bl0J44MvgZgi2wNrfmhZlUTqWeyyvDqNpX5
bFRtgWos7L+3hPsNpjHk1mJIzetPs7bWZStMiNiDvUCxk1+2E+mGeeDMI/dVK60b
ae6jDfuTwkZSDr5nJVwczOnicxN9MzbRzIgkKsIXqQW6NDtxiynncWpiJdzzsPaW
vcyza2aNFSvP8XCl56t1qlMZRyHo1BqaqY0teWFtY1wln3yIU/q5t/urvCHP/OpO
LbPBCRo7z+rWUzqCoFILefu3pBBh32NOqw4lJJ5vaVTt4jPPvNFYeDa9xpeSd6a/
C0UvxrH1ehlgyAkmv8k7SGUA2/LGHyRcTypFwTG9zc69Gw7p69nNiAWzOh/4naYZ
WFVXp++1STZeRh3pqxlCFpYsdP7BdyWHNOm0Zq6r7PwhMgK/AJCa/5/hvrDescE+
xZ8fTVJRl/aXOV+0c+tKy4NacFmrnzMFm+Zu9KpunI2X34vbg1j40LODZoKKkklQ
9jSTl0YviB5QxH1aKQUWZDpizG9cLV5/PIiK8/xGsvLvi6H211G1MTcuRU0IUauh
QdOZkuQlv9PuB62G750p6CXxYSlylaiseVZiHYiAogeyFBOONL4DDDeZTyjXtxe/
4znQJ0sp4xjV0Y+7+08Vkljhha+Xkp6Fs2vNuvdF9H1TMhjul4IQaU+rNnKYW+0B
IqZcAMcdDaTWcV5ea+QtjfcnRTNJPUsEyMcH3rfNrq5gUS0tzOauPvpY1bMb1dgz
QmquoZWiyvy9SS69cHARmceStMw9uaGoj3XxL5n8RWt/SOucAz0qRyKsw8XeZykw
k96R3g5+NpcPvePrE3DTLSNqFjSCcl7WDYYaJjCxIhqB5sHEUDyRUAv0oJ9Nj00S
2YYrZDPwm4JpyeDM6L0pKzQ0+eyA1aJ9ev6PaG5wB5XYj823an7cGfQRUyuQS5M7
f6cljAYj2ZmDH+qvhvJhWTjDYx4GwNQPXd9su0lyF4rUnmDVk8CdAUxNxPSdvb5i
N7KbLtBCXQmVj5Ms+qReVFVZZTSKm3KatD4TD5fYGpbuOdxcKgZ8Eo1NVL9/gzs9
YzF/w7JY9MlFtgH0+fxjWQYR4yxovulVJ+XY/eqAQaFYJ2NXwKV6zPdljiMaLrM1
gZQuvy0UNcM7hrBA7OX9sLOrjY0pI4/rEo5NH06BDiOdvJFOf1wHY4OUQzDSe6+M
bpj2c4ZZHH9Bl/KqWgzQDDILHT7si+B/vQIEDKHWLuhTTn7UHfdjd1TyUPORxTuT
DbPDHa8PbYbh6wLIiiX5IFWzlo15n74YlJ+yuLVZyV4T041FdcSI7kRw/tzaOByI
G4XEHOIq1S+tAQ7Dteb2oQNZ6Fa5gEYePvxoKAqd6773YWsG0mw7xDxMXhKfo/fJ
hJQllQi45/lTwtC3ZDA9hx3KuRhnUYCVJ2JL7lzRiyvby303JLNtHWfp6vSB7bho
tHGVBWNwkDZM6ibRg4rs8CujWSTkP3kzrqIBnzBjJS5/smsC+/yMwC+cWvjoq0U3
dVXV7Q+0PLId5WBt+f9Ydkp+MoOE+hwx6OkionTrWnGdm0X1WD1qIqYoWyQIY14O
5p1QLjWymhx7aU9DD0LwZiMQMN4vwzgHZSarjceq5SjP69qV4jo86IvsVEKX8AIt
JV2nXCkSUyUIHcs3DVsv0FlTehYEBcWikNItpTR6rfrcHwjU9/YgWfjQi72SrI0Q
QWXu5HmxwDwccpX5j60cXaxuEPjcDA3coxvr+TRLRnT7s6UDfCa+DOdvSuKLa9lA
KWHLkf1wOm3mMd0o5lRUiwgkP4GjneMTd2rGslH/P7RuiFmostMP7cHd66WyJdJc
xQjLZmQecxOKAFRdBKQ9SE2d+qUC3/Fo7hOla+YVwk3kyObDKkdubGpUqhCBY6k/
JB3rRkWieRL7CGMwbfr/ZQp7DJq4HCt5Sr/HfhI0lG49ZtNku+GLxTbgqkFNYmRh
Q9M36ThxH6bb5gq38dM1UrPA/n9yjJvx3PedwUXe7QNpgeFzkVBXkPXvpaHDV02N
qPRR3E1xOHzgKLtu1yuRYXMh1CwKf9eOY1pvXoaaaHDcTMtPDMx3BUMADL51qB3E
NC19YCFukWOWCYSBbGD/biIhofi19rQJwfpo5WzrDPFYh/C8NcWsMj7h/U+bS4VY
XtQe93FsRuHsJQLqOCrbRLI2bzB2jfZ++EpRW2F51I3Pjw5tt7HXdPc09fYSmM9i
7X53lyaZQeZ3vHpQgi8dU82PM8riFhmqrdI3XacLDNuKxEP2Q0neysSqLmy1kwOG
SyrKtheN1ar0pR2TP8KmdWnFt0wxRkzPNmgDk1IUlyoXQHpr7TnWNN262JmYL6g9
bE6HKUtzU598ylmQ8diqB8izZ8hm40jJt3eFqulpqymPY8r2gmEKSVOBiVtiPafU
fJpOrsTCzmmjo3rqBIhw0wjDfwfZcK2Y4QSZtEo4GWpP2m1aKsuEYo93czEAaWMF
GnRSqsPy7zJkQfxG7LlHaW08eh0OV2DVMGKZlFm9tAyGdpjRDdIH5jK/Uh0iC62z
9skAcxKrNIXHbN9mMYdw7yo+rnpXZixQ1zHMmj/5ByrZiCXB6dw7LaR7Uzf5u8nf
citfazwCkhe1sidTygDQnAwgPktKMdSxbs4SeMA5mnCRrEuYz+Nyu0jItK7c2RqD
nJ+tdFjSCVdZgfyEMeotDjC3O8EEFxLs3coLLCqsSsFsM+YpHGkaNFUpYVYVIRLf
SZsCsPo0mhxZZZrMvEYJYWPUnQ4iHD8sW0sEKG6xmQ8SNscmET6LTxSdpsow/mQ2
T7HbsCGophFbsryMyQZBBtfl5FPYPu+Iuty9b/3220rjp2YrunIPV/jBtEax9pEY
w4o0wevWkXafOJrGnp2/fxt8KJssa+zsxnQPuj7M6fPxPW4kvfU0KcjanHR1OqKL
Z72dirwcQxV8/rq6G+P7fG1rxLdA8uLeUZDATzWVjeiRhSvzVWkwRsm7WqECVn5v
lDulR3nYoZuCqTvFq/eYHzfeHj/nvGEOWp7eSXoblR1xZ1KCMQNffB+PRgnROOpw
w2PdkI9Z8AaCRl+AoModGjbWt+i0s8jxOhqt7PQdKxxmX2RwpKTmCCZq3frVgJU9
lNOLzfmwhMtmoYu0EHdINZprDEepjmnyAtCoX0i2PvDqrbQsxlsr1Po2/UQeybiL
6Ho3KTwhcjB9iyhMALqW47rxpfRwP0YxG2peddExIrLb5R0/iMkDPr11n9S+h7T3
WIMn79faLFs51D+qxA42SYXVCmc73gZIKUKbqVToeLJRmgD30ClVu4ExZlWR+pK8
Cj86/Kjfyxa49HNqoqHNWJF9SQ6/q6om0q+m3zZR9Z3hglYtGojiHcLEdYh8K1+u
6779SS0qObuCdq/i6Scn2kbEGGxFZlIEXzFWgP1mOuRYoGBpam2uxMS5vcuEZuW4
blv7h016qNoX07MzUURQ5/lYEvwxlnBj9uSRxpp8JlGI7INPzG9Nm9MyzlN0boZx
1YNem+10K5nDVhP9mqRDZtg6FlSyQgpDGTmJ1aH5SAENPHDtE6MHw9NQgXA7dfjC
DFHLF4Xv9kzOuTrNIVwTzCzked/384nyDX5f/IwKwtgPiQgSNPGKhveltQXj1GWU
tNLr4jgXPQkjKgt5jhfmZPgi3wIA9/Ep4ee493+2PIRQVL2NxMUMlhiVhLH9BsOz
32ZFWs1usiaYeftaTbqb1w6GJPjwgucOr0Wap1v2YoNEDSfJU7GNLFhO5cZNIhEM
9HG8X5B8mMJ9DmOud6E3NnU63xJdZrj+ZG2RmDbg/UR95zVb5D/jPfyLGq/msjDe
aBl7haLRgf1dEd0U/vFJm3JktEJlKzpbMb8MWkOn29TOdTR2Ld00hr9PWka4NeGc
BC3oTFNKpY1LJm7RQpmkN+1NX/O9a9nwrd8Cpbz0/ee7dYL9XkPyhaP48TXFTeNY
yGn+3V84KxslNdO9wbVlV/cITew+2epS26NDAn4/lczTePBEpwZ1xIJXGCS8TztM
zfOFtLqA33ZFywxQJuckGdizs5YIDRzXle3gcGB1JjaW2sJbBYJpmhZ79/0F9rdy
T1ioD/BEANzuI0Z2B3ebhIlDadOS02oGtEmoVuV8n6WptVwvMV+ZJejc7wvWdLCx
V5ztrTDV2IwGTFXNrAgy6HIVPy/pVzMTyLU2W5/+v7oaxQeUfdEONVKyst7f70jA
ffg1CWc+PkX8cVPtFw4x6H/0hRyJWqK3OjDVw1nqh5Up2P3ZO4+LWWv3LGxa+xhD
kJsHTWnkUpLtv+7cnGHPDEibfezJfUeLBv7qCJmFLuR0s3H1HZAO+Jb9lPO4jBrg
muTwwDC9kVnBUlfoWQm/r49wIj9tGqUcM/DDaVrQtY1L6sSqz3Vno+RHbn5N67Bd
cQHx9770jAfTkXa52ksZEgBgrSfpCCfk2aq1JxfrrDvpt3WA6w9saomtdlP6YdXn
82fIdpbqfelaViTF7uBJPFedaIYPOK7cziktv8aLygatOsZV6cR2/yDE3T85Dm3F
Jm90V6SmTBFcbRPTh92waNT1Ub//E+hnPxEMl7oEmvFCZM/toCzVkU4eWvcW35Zd
wqOYL9WqI3amn4lPwqXQz03ZmeSEQGyA2OM+AVnnBqXL0ZiakYCMEkzb91p3vLkQ
XuIF8MSX/2Ahg9GnBV9X9YbVoDSE7fDrlyMX+uug3xfKjr2BNrukVGQv3XuQCJhH
VlOIJ7cxRYx+9t3pgMymeitmweeH3rqEMI+5atX2r31PZFRwsNIZGDIP+D7PRd1U
qlSMBcrA2ZPs7lli3rlkP6pFWoW2u3SapM//i+c1fNykWDxtEGWer5L7Csm9E99A
I2NbfYw5eSsAiuX//EDO7L168bQ+a/KTzWvl778wZPY3Q1NTEjKh9qTcnMhFFVoD
d851fDlfRwjINrYL9bOhPfQxk9obfhTbvQQ4R+XrnUDKAymdFxAOczg3Q1hy6M+0
E6zxYxuHisAIYrmk8CEIBvXhs4NniEGlOO2iFf+CeEYW5qR4sc1xa4PXOqhjyW8I
sTZ3shh62K/IZd3D/8OiULuXyUWRLwCSACyE18tEC+Et3iV2HLjudL7WV3tk+8S4
kNYFQl5ek5LRSwRVPAmbsuzJJWJGv2w4j717MlwffEPoHSAmX5CMLizr51SwutPe
HG72dkjYKvVo6cRfqCNsyijp8CfULDQQ1XyFRXrLFBo3kvbCYLJ9msJ/Qz8ibMIz
PMlVlYC/tT44VOE6wCIHtSqbDS7KpwQLXlhx79o6jUeqWgA7aQBC57KepuDpMC2p
WqDLo5KRSB9wlusKaJ7N3v/tnn9gxHEclwVBmr5MYrmB9J9wbrXvEWUP3vaDrH99
m3kSZSZvc6DSToxIzaV6yuxbOoiwHPLQKvvWUEthejSbrzoxfH1k1Py0WDGLcvKa
reEkISuIVvndnX4zDoYMtMUrSiPqVf5vi0CVTnSUlmzUqrw/CCQuUq2eA8i0LTc2
AnBrTn4rUVlX7IfpC1EL2PZTH1basGDjTM4gIb4ajQ95WAeW458nAuyssU1Hlqca
4h/UoNWPEVVDhYuduNvdRxMWQC4hCtYv7AZINMJGiIVVmDvQjax10wRcFR4/Isle
T8l3iQzcadSJ67PsPT0Kyy0rEC014O0Ou47ZwPAW6JWhDCQLgEIdOkgK508advU8
5ZeZNUnzQ6JDE8JKKG4wlW3x96Qiptc1fdfQruqSPHNPUbiU3DLCQs7Br24Qa60u
eqXzL6HdWvcVY2f0sUym558NXMsY9jDeHQG9btHsKdrJXol9M60qqYClRsjc9NDM
DxiKPLGqkECMkka2+hbEg942Kc8r07Mcyygsou/bicmAN9+D5f+5djOSX1JOQbrs
ZJzFcMK84sIacVpG04CueSx++YsqZ6lReU11lL77F5Z+C0p2AVnLGeFvEDuH6ZSm
OeVYSuhlWZXgutwgbdl1Eksv0V2ALRDUEDqOuK+CbEBk1RWS+VRmnUJ0loCHQfI/
oTkfSs0/lhHbUoYvpmhhkWgOfxj6VL4FwBWILMcwIZpDOJTXcGKaLcPxsffitLYR
+yB97V6rMx6SQiWUw9UdsrTgBBi+rK0GI05g8KYP2nBaO7KHaK2SZuCDaRcf9stc
4PMlTX0BeMHug/GqU39VjZfClXrbEXolw86YHESi+gfmMM+CQzHgbgA3nFbCr05Y
wqBzT3YzZgMxwy8vSQxRmHL96Dr7fqyRuHUFJsLyE+hWe4GTiwgME5VBmJjJhKZ7
PVO1hx3V8ryfer3wYwl0Lf9xb8InFF5H6cYwiKjhAmFA0Ht1BQeLqzyB/2ScHqBb
34NFVMG9f6uwX7Q852nXwwZ5+sKQ1WbHvQPmQR+0aiOaM3LMpGQkGFkDzUOj5ni3
OejG6hLE2cqotUmFG6DM4f8StdPCKBU0psVa+/owpXCf6PRKO+0De3kS/TTVzAKk
bPzPZR9VeG2G50LRX9spEeZmxvQWjt71rG6Pl9uCfPYntKYmc20Gej4GEvEQM14k
nMEmnEAoyFaBwhdpBAeaInWpRfJAmJvtUMH2dEFydPeokgumAOTmi67lgmwl8JgA
ORCr6aU2UYlW62y3rdrET873WCuj3uFeMmGA7Mp63VHq8d1OhPN9ymD1YRn7VhEz
AIlClQkBlGLxAGqgYFo7eWed+IoDp9G79KqdOvW1xFVH1ks8dApFA44W+ki7EYmK
fOGWHRFpxYk4vHTYUWj7JvfUk/eJTEbmNpsBTDvPK5sjtwCeW+FCLBBLN2TbnWV+
n5uhq6QBUMVRdCKF6leLrIbN9AqcRPKg3qm4l4yhR56J3TH8R5qb7ZRGPdEQ+D61
S86b785Z3qI5AfCOQ3HAbq/HRvvWh7QOlMYpDEFnrUYJxDnIRUFcQzM79G+lvZi9
6tjTy0oBNmdoHP9NjAcK21KO3pMaN4ZayUauM18rRC93x+RRdoXmeJJ5/rPl/zNe
M7BczBMDzC3ismgniJqdG4vW5RDCJz869gEx0wQSa+WIcVlQIhxLd1H5Wh3lueSR
jBnaZAdyUdczJsAuJdXGL4+ChQILFvpCEVJF+VKgjsgElO4m8UK0F7MT0MmcDY/U
w/Prqoxu9gdI94nAtz5hrpLKx6r7wwRZa7ydPgGTJGTpfVSJ7W7zbeFjoNuZyVQT
wphg07X6t9C/hKuzfU2t+e5B8uCpMOpHV3x3unCMC8aTfab1gk6vqgaGt4+FWMHr
NITbnRDpjuiA5+HGhF+YSDFVOBQ14HKFBAhKOAarsCuZjUml7SI5XzLAeY65nrn8
qSHd926yr3ODMS/MqSIRE+J5w0XtyJNhGxXi3O4FcgPCY4jzWnJTWvqPfz+SG9BL
UvP8CDX5MiKyK78IULY4S2NCBSKHUfQVvZWkyXVNRopnWvnFZ1piNyq1SzeMuCSa
r+jtNlkbADpMexz8U+7rYEaVbToy4AltD6C2eHIcyB2Qzltu9jG7Y6sgJncWhUlu
CFcsO/OITra1S4JN8sSLSnJ32bz654XW5SI6irCq78qFGh5BWfQipWBm9IYzbLjQ
co+E7ZZZqV8utrleAVwBL92oY9MWUQzkl+LZWugrd5V2tprzcyeskemX46o4a04A
Fgv0E6wDaktC69bOPfny32yxhb+6V6AjpHD9zdtQHGStLe+CqHkNHOARb2wad6x0
wMz3bZePj5YDXa2qPZoWyQYdwRoDYgO3Vy0aAtahHOxylwqw/g8Z8mDpOwYHmFVI
Hg4ejTbUPZD40RmeoL6QuUFJANSamqIANFaXYpoaRaaqjhA6Bf7UeMWBOarzwgE8
LPnfykpqT3AnB2Trk+g+5xFOytvaPV7flDaR1PBeGrgaR75hFZjY3zgn+j8hGof7
D9fZmVvslvKjYtV7wLnur7/jrbuxqN1tGTxX1qYdofO94CqfjXd6uuAHsQsTMsCP
7ZPpAuS08WGD5shYJquSaImGg2mJYfU+rqZs4/4INyUNSZaQ3XpdE1/qLfN9Fc/d
xt/VjRsoeTfB9vOIBYLubIrD0abW+Wly4GELU3nLrMdy6Bgl2vLpuTgEQtzvcalN
1R6nOG814o4UIKsLhbsGoptAStcj5fRxPGfojMhZ/uK8RhhRCO4HGHmCkGyCR/na
/iL3kbBG+uahcdlOSeov1JJcD6yivdaSarL/dIFn1lKpGuJuJHMgZs3j9hQjOqF1
CRq/g3PY43sgs4VGMnEXVe9DfWi0c/J/gzIDYdrqDRk+DEvfCOGrGLguCVhTgLbC
S8caY1SilghIkGISiwuotDRws7jG/F8x7vkh4JkxVwIHsRytmB6LZ8VozQ/NbJto
2F9xBgvgEOzFmslxg/xBU2fjGB84d1S7cfzTdqS+SBWs16RcLe9si0hO81eBkaIy
+cXi1rkHFRjn0ueqoAcghUt2rQxKJmlYZv6jz0fdssj8QoFVmGprfipzg3TP5snB
3aobgKfpcToDdFyquoN60xqaF0tIafgnIS6BAhvJyDKgAgHkqW0fCqXkg5Luz5UE
V+pDNSCWTbYa6bP+sVQN7S4UM+JEkcThJufLkDD/ul36v/NvyJSIeeVAvoQsBadx
Zg8qF5fZux4yfKCgjpXwbitXxI3FZavCUeTf4NyYxBWuQbnRK7B6hHnCSLfAP1XJ
vvmrshSU2wvlRf9vqJVo8gKzAbuprrnYpp0WS1BzLQO0LPx+tVuKMNpPoYvVxJBj
WpHgppRyOMDmKr7Hc4IWfHkvddJPkyVoZ6PYWiJl+lPdeLNjfgul+PriA65g79qB
kTvdJYtnwG01bvVy3DSQJ5rpU2jQzhwnI8COWmi1uc1Tl0Bw+aPur9ca8l3cWZMI
VctCaEqqJNToFALibPXx5sM6CXY2ULagu3Lt+AsvdqjU3BmIQrF9gNmMN66S8Og5
4sKHYfgdyXFEoUvzlq1c4DvbBc6MhXhvGhSzE+GljXgcOk17KZiOoqxC4JjPguf3
RdyjMM8gOBSWE/CgjceBLjdjLVX/XS7tD6kVEGewJ9ZGJ44CwXw+XUAFiOJkJ1Pr
E+OZkZvOIJEVrYmYSO4Lxm2vNiawuK0YbapJ36RpJMf9IX/HT4rIPZ8VulduUXFv
Dic93+ab+z5RUoOSNI4NMj0qCZqD4eAeFVeW/FApCeDGyoF+WnJngsWk8nJUtecg
USRtyt3HpG99XKFtdOx7GFLuwI3cGfROd794KHcMgcNCtdbdqOhUq2AcmDODSk34
+YP/7lQH4/vJw5ooN0XKtbe+yRjGaR602jXRmeWhUzEYWx1EaPav7UYyfQc7xeDa
HkHd4LJcDM/g6mbSn5xOJ+x5x/vaaEd877NERNCej3uPyAylQFQkJ4wmRSjHjihA
+LC8sm3yjRIFWPqE/30VKtnzJh3Mucu5RbzMY/scRI9Nm2vRZujGuc7TvVQ3vl/I
P8erSv1yGmSAereMtmpBQGfJ1OlsI6jKxa0xXsrcuHn2bHFjeHGQ2tgV6xIky39N
YIW0U+Buu81o0GUhw4ZXdSk7jNVLSVq8pleZ2lmMdsbxAmo6RUoHQ5Q6GxhOVfk/
sfYc/h/TndQ6223e/EL850pWlddIysarDdNybsJcQZSCrSsmuMG9htntIRsT/Czj
9cgHnar00+AbTIkHpmjovX8uSooCuUci/fL3er7W5NLNCjdjfxdCpIvAOC1AaTlF
LZwPdQ0ApyEI9qHS3PnzgNPftUTcDCI2LtrHfItbqAtcNfzoz852ZBVXk/r1uZr3
YzsKHvYkxuJE8ZySKKcH7nOqzv2rGrnUaEyKUKyOxV89+2PkepBBYIu0dPAtQM+b
s4HSQmZFOER/Wkqz0XXI970F0zye889aHs3DgEaqd5oSmtegnMBnCjn1Gch4jkzE
B9SJq0hPBnJaIUWUgOl6ObPUB8x2F2hPdkXZPX7Nq46ZVYacqWC55PvqKlO0KPal
lKtJttiU8OnyzhCLQKbBTrTpYAHEd8JR4VXOrS61fwvb905lwhvrVLd4JINEX/Gq
VUZ6kVaNGjO5mqihEa2RPpaZnZgKwdNd0Jp5alZrUWlzL2BQSKvAlmOOMjl4tfEH
9PwG57HPZB9iYg+30pWzUnwuoHgbznqVMv/bKBOxooIRfhcITQmoS8s0TpoU/QAH
sbANcRwg2ybglGKDpZJUMkBrZKDaXlUbZxGXLeqewtAppd1tajvtTVKs46fY/ICV
EWQpgwcs44pleZDSBlDs0VasWOxlohg8Fcimn0YuV1pDM0W/iOQ9wWQj+qyN3oiC
hfHTqzvTMTuvSyd71fvBd4vi4+2G9Y4lKUOOdvh6tl5lb1qEApGaPbqTPPROgVe3
+zqN+6w/6X2Jbm6/KDsCZd+K+uoJU5taWa2WBvoTLhjDdHMItxeiq7HnYlSJKkrp
m05S5Kbyr+vQFJVpNTfmDGJvmF0/cxDEIp3qB0lXE/zLjrjUbXY8CvGoRIv0vd0S
F5QKRzc/i5KWpyc3LxE79I+O7Q4NPZtqc/s+Cgkc3LAygl3RKfWM07p4h0MheV/i
sLL8dBrHWT1ZxCnzAZgRri8ZYMHsuKNSLxIbKHWkQe0JRpsyQIWnKCyamY5hZrqV
iTJluial/yZuWrgFsSPRbQHtfngscwf60aSfrovQTvw+FxVCVdBAvvITimT3UFWg
8pIG52wgTMqKuFIuNWK2SCnGSLlp3EcOz5xDN6tKTVDBe8MR9CezbIWKMgNRCohg
t1skSHHe946A7PfCt1NtcDvJX2BA7dmJXD2Cx3TrYgYIo4Adgh+Rxx5sLrlpBEml
rhj3mul+vVQD0XzrcJjo3gp9KNpxF5wF6MKRmPFsTpJ0NEYruZV2zfPFRYyygMR6
VIFEJSq85mdILqJEtTI2fH1+YcpgJM1WgehnP14wd1qdD9u1Or6+2x3YhATgEmnr
+WYdLRmf+szv2nc8ciOGzShrvZXSoa4jShN05bEQRE9ibZQaa9FB6uQ8UuDKG3wF
FeM1g688tHV5ualw97oJoWGckpkAgVMlq8kG9D5Um6YhJ4D+LyfF4ITwg9PmqWWu
RMbCcQtI9ll5canEp8oXnakTi0/LQeJmwmFP9GzXbjpbZ+zsfeK2P1HfNen6C9gN
L28Qn49AXBVSHArz63S5LxtSh1TfUJZpeZiYcyTL3LgFG7MB8jdo4r9BQohUzR5J
YfEc6Z36GJBaJXZkE6bHBv35QnooVOQ3RCyMTPuN8G2l35D7ETVbcdkNVw6jz4eY
xL3EgGV+ZrzY2O9llIDTYCnmtbz7be18LC9IE3JgNjAaXis1dfmIyFwdbC8obBl/
Y1HkjHslFgDkW2Sdpj/Jx2NxLMqEkdkrlMSY/7f+YP3r+gHEYl2fhWU+bQTxtYI/
ExD9nepTniGtYJfyXODTWk1Y/btH8HwYRzEd0mnkc+L8JZ3VRL/jcZDKYmsq9Ghv
gFGm3WqB0boBvY9BD73HkF4ZZ4gPygQP/jJrCzMglgUdHvFWQAHfAg964KIwVmEK
REP+CFLkB3kIwYdZA4tCD7SxCnOOOCcL30PNGUFWjFOjuSImuWAik9qUelFeH6lP
knlxmSG26IFASl95utOsudPfDXPpZ1nXO0vQIykG/Yztbso4RpivK4+NvjwWMaT+
GMCdh4ItzIpEVi+SRVFYSAxRP+Vprhhz3J7lxbKeTM/S+/02Ufs7c9yHDxr+K2ue
w5TmCZIJEg4LWdCSgVe1Lx6/qHfNGLV4+kHcmUQ8qIMWzMrxvl/h82C7XZVpReQu
sEZB9T3S3O1oTY30pNlw9pJUWZo/1t+gyj/7Njhm62ptACKioA7aLp4D4Nqi6prR
oAOQZuPzyBxYTREsX/DyxAcNs0xjibURFj5SNbVQGnE/qiDK4pJI+LyBMqRClnIT
EHvv5+rMSlmNYhft9PH4Ks9YqcBIYR1Wl4Z+HVqE/UjCnuPIgnlbD616NzCDd8JR
5rsj/zR76vWDHRd9w46gxTbmbEB12XvFZ+qH9PzfVJKWKxvTvjYaN2Zoc98+msPn
uVA4Nms6zg4wRNrh1T7kMAsP9iTq0r9yMGPBtgU1g4hDOXPOqIxHHAmtlUh6f7gM
R871R0TkPbAgY4WHk+8Hfq2rKtVu+KNx2gEDZTZ+YkH/oyNJ9r/OdwjjGaR+g93q
es2mcGuEc5+c5faWSCLfQsDTV5Jgi3MDc9efnKq1QHzOjIaqCIJpOOF5XTuElArx
GaesdWeIJqKuFcnxgGfEPpN3xwhkSe5TrfmRaESQ5ywcUTYRj8hfpapsulNY77U7
+yVptnk2aRfh3VCLfZCywomIOoJBv7Dc+P1Pkvbqb2R96Gml1aHVljrEAr+/BYBV
IwyyOJimqLs0u7ZozVkCHCxFvv/iZruSW7zX7wigSeang47PbFHuHqG68oavYqzW
CnkI6G+N7eBMUFyI36G8t7UrHfs138XMZ/Yw9uR1apBQXPWUsQexE00PKtQBSaJs
bltlcXoCGI6KhiYc5ZqSyJjEAeMkZfAxNbBsDwOkM7AuTYWjDoQQb+PCA2e1PqfY
HvRuQSSPC00UCFsBN60AvH7r3ul8iPaUY6mZyt8HHJBmz8S0VQ9QEAlLb5jsul93
2eToFlLrIcxNA4S3kBzi6fsy7ptjsRkxlV+gQVgCkpJu//Aj0SjXGS3irw9ivBlp
6apoAb6ctqulAidbLXADcLw/3TZShY9wXI8SWobl380KyIMv1GyX7B/icvOcBZ09
RNDZ5Oj5ZaQEK6jrZU6V+0JVDXkBVJbGfy4tndPPR2oBDoAbA+0m1zi3yeaVOpZ4
4OWuujTWKAevX3kv5hitNjO7OjI3Ho7PVphEQNsfXVcD+14DG5TxZ/361X6gSIWt
so7Nyb61uRpjRqdggxcfxx9eUDy3w9v9QJ97sxPkGDt34OnpX+t28LOvBrxBAYmg
8URfqAFkK+0BpZFyHl1B8wPwmB74b/TqoY4en6TNNltILrswon0a3/bcGMFy0Rcn
FbiAesrrgIdhFR8yASkFpgDuOTCUetMITCXSCCTWFKy29bim2/e5bWK2lvZrk6UB
I+qWjj/5TkTuhdespBzDyp0Cjl06T4qDQGErl7eeWhGsaAR+YkBBfCO4U0zEBUMK
PUX86ReKJWrZnQDDv5nOoUa3ZPlFDrvJi7+6DdpBwoS0YRrjAlJdez7i3p1IC8nN
PjZRdeapO9/vM/V+SkRSrs0f8ONqP8XQFtiY1/mFHWtbWDZrmAK8Vd2CjYTwWbWq
nebNSrhaO8EAMHVTYZXZD/mbZrKNLJWkisLO83QKL3ddCkKnI1U1lUGEmY6FKg2X
2GzsU7pm6d0W9B+tjRLnflgQGXfwGImt7opMBQz7bl5ZVdq6WzqJB3flke1tL1ff
SKeiebaGTfws1fS45n23NmoqBRylVmksNuQgYe7+/knLR4Lk2L0Lp6vk03hkrYpc
rJeWHe9q6gKXOWc6kAb6HVFFiNDD8liDiAfsEzesv3UdsOeBQ5CZHI88/aA+xwgY
kDNihwggVzzmL9NSQNijmyQ65RXb58Wv0qtKCRd10auuFU/AwEQ9SffCwxBsR4aF
FQRtLuyf/aubL75Z87aduFBF29Qht2VJsec3dA9puspy7crzgHvNPM49G/gbf2AK
llTr8q6EaCgvZh3rdtrxlNEHCerUMWupPZSElFyDIQASHMRGkKceRVlHnl8aRDCB
C9/r5SizXm9YlTplfdNf71rHJPRHpV25+8L7XLqY0/8xl+VVzCv4e4g02B30SS7A
nBjg1cbPHoXF8MyVTnoA5eJGdun31hoc8Ts35WuKSQjX7bn8PlNsAZC3pZRYOswT
NHEtoFk0lwZ9dKnLgId4K4pYMaKWKh54g6UeCce0PmFVu8y49YV8SYJaq50Gcngo
ACjtNEYrxeBQ3f5dVzy5VKGLwBJLsCAZ3y/frRRgYEka5jq9VkBi2hibrzx4GTij
snCnJaQ6edXh/smRai4R3zV5N+sXIKIxNoT7tmDyl0Qxy78AYCSbkNoBiaFHjcko
9xMQFrvnE6vuaujI2IweoCbj/7CLtb9eHURKv/T3HdMMdIWe71n99/369zd6ORKT
UV2MBcawL5+L3RLiq7xcmaPegKSyQ/qBRfd1+3Xr/MhMFkqV0d4AnZXHQQ78A62c
JCVFOqYSj/mm8edobQfIunSSVZdW9+asJJX/pMPHjoTF1Sf70jsN3rHMUBfkWzWx
6nfC/sNh3tC0bbUyzs0W/9vdt3mfIT4CXD0lIkaHTn3UKInRMgfB0PBVeU3Yw4sy
P+DXRvI9fEtOc0FNt4ZgVR1205WF9M/uYb/fMZpy1qtwtLBcUMy7BoB33agQXR7b
PbQc1Di7c6s6Hh10mOB9Qn4SRGqAoSlHyi8lDA4Ni4521bbzrYfUKOfVUa44F3l8
THc4IDMw397StjE9qjkN0mdOWCoGE9UZJvXZc2fM5klpsd8nIwAqWZxPweFirlO2
DsI0LdNyRad8OPFu/9Kj5A9AMaHsx1OaDJ8I0qotE5E3OIK5o2SJ44Pm62VwdfOp
rkEPNNouHkbWl+BoCuq/CjlYTjqm6ll1sLyeEwGsTS26Ma/5vVaJS+4mNkQOoWuZ
Ed/uTylWj4oRvcHcxst6HjUJi4agA68do9/PzqQs07g4oqTaUBTcnKkxLdHCPXKL
Hh+b9CrSi+NQ6NAxuNmyfSx/9zLcj7T3DVNkrk2G/Kg9PPfLclV7/MEU7aD0QfxF
hPv5T5KDjszsRQYBQqYwl5O8VgSYc3OywWbVssgKICIoc906AX0ZfOSB6wMyK1ez
1+6/QKHncySTCONVKGvYkXg9J4iliojfqa5zGdqRn5dzLf2WVXvP6vmZaaR9CJIa
POM7PaMgFngTOB32LekGR9cktwsmE8+4Enh6O3rAEpuVUEOlJeFjXyZsm71Dd2Hx
zX8wGGZFHrYywUE9/axu+vm3fBfKR2GEYEJ/SkhXmoBsbULfB+0KyyM7cFz1kXK2
pIagdFa+5ZN6nYgf8TgJxexDDau/D0Ar9M5z1QGkf4JOM4P/v7muiQ7nM9QKBqhR
SpL0qTO4ebJm3NLVKnJQWkKEujm+LNBloDl6tjZn17Ifu+IgvgXDOdL/43Yeqpdn
3EpYIyheKKfN44gG6ur7j3yArOeV2D8I9lSu01alGrHShmT29J5NgzJyo94yMZbX
cQkVkiTwmYo4FIaspmgyVQJ9/9139CmejODBhz85Wqu8IgzhEyYPSdcTEqDi5CJF
6b9T+eRvZTD59uq7lNtgw6vHGJWDV+/PWAz5PtyxkQd6++plZwuBjztV/ESEsxjr
iB/46Uf3ciHZy9ELJ1+zAMq28NNzB8QZedJyO1LBMCJZ7PJdMqowxohW97kJhNjZ
LcsriXJNxg8qUvjpXJ1mhtRsxZkE+QNNfhmSDMl1WNPPpYIrH4yprpw9VT9g4xyF
fno9zLtO9HQ1RZQdpAkJM2hyzr/tGOqvlu/Uk6FpB6zXxvFTGjaUiFvdrX6/TzaJ
RHbv2tjg/vPz5L8TQfDWIxs4L5tdy2llyzqm1q5nhiwcXYLN7a7mXbFzwbsenulR
SNSHWDH8MJ/MvPnZpU3tPCNL/2Il5ki/IKEdhiiJQjyG2rjyDfo2e2N9FzovvfBJ
owzviG8CjV8iMIEva0Srnx8+ajoaXCWf+eFC4YoW9Mu9D44X4SN3L9Yg84Gf/KXm
qPQxDi5nnfGkNheObi6NvoVIa5qEUoXrWqjudMekpIIsCGDMpOD8iSdBthrtj2KG
/gOPLEMSV2OALLm/UQSWfjnbh2TTK4C2avunH+1mXD4ZtHNIeYdp5i8dfswxoTvc
v5ZJnQCxvjNYTezs7RGPdSH9DtiortYiJ1dibM+baZPm2j6GnV39BeNqhk27aQck
PSIN5HraCaI+O+FTG2cgs+l4tTlteHwmswkYruJq2XTHeAgXSj/osKY2DLYbFymF
8m4R0+Ufl3QZ76GHG5tHjJPJ5OEloSuqCVQ5+NVAJwy5eBpeZhptrZ25yOW3vciN
tJpzqqpe1GL1nFCqCrzfq0t+qpVOlAtIJ9sY6smFeHNOP3Ib8Xw08GrxkVnaoH/d
qSSORYqE41sszknKSfQZD8Rp1qfOnTg+2L1Rggf5gAPXBblmXLBzcC1p18w4+bt3
KScj6AdTQCn93dMsptBqW8WA4uRXWroyNC/NPYvYe28ylU2yKvB7RwnSQ9qoiesO
RTXsCOB5zxbT8PbzO+mCJ3bD8h7eDZXPOjCr+Aujur4/C4WB5znE4qhdrG+vI44m
x6jtGGpxuUsGIXYmBLTASS6mLxLuorqLR3uzuPjUYlyjYtT/KAj7x90fnZPIqw2g
E8TKBbphI2fPjOjF2QYRUW+NjbirSmBsnBL2iEV2K+5ayZsPP7g6DgsqpBVz0gdc
4JbJnc/rxhVkLkT9BF/oHiN6XPDCq+gStN2eNPMHU5lQIrfvJ3ffhoBBJ4jbq214
OhZtXy7F21rurMfFFxBOeR5d9c1rD0WLIEL73By1flqQV8nSO41mIliIWvR48+oe
ne2RbhDrJCow9MjniwW7TbKaCt1H1vFM2I5jKgy8wFFbVnrDJy8B6xhn07y40jhD
lMDGF4neNfW3+HMp+kRqAsoVhqRDkVTqLbsWP3JEJA99uRX6pwUadBKibXSrxKyG
k0C2aPxsUzKjKRifLOJ/Y3bGNV5l6C3Ru4WsDkGoVGd3E+VAHbZ2BejPSgDhFKoB
q3AOz8hsmyKbqmmBg8bnRtAkCNGV81HslCsPacrGPUKdrb9Da8BMTMmA67Rz02xC
O+IxWhg61f2sj9QaFxbtXHsgDTg0diF1Kitt19SqGxGr6Rrz7+BykNZnksWUaalA
sQ6acyOf1LF29K5j7CpxvLKeSQMeW7P/v/OQWGRv1PlSDIM64/7YID7B70wpD6Nn
MdVyO4RvyEdZ2QZ6mRv7aONmtadUiALrIKikUyaKfXz1kImPGVf5PaRFYnlTQVG5
oHlgu1rYXXMJ8iePdivUXsu1CfHoUqwCkMkTXnf1M0iaFXalQvQpJiI5GnAhlIay
XZ1vdEJhq4Je1mGUzpGtNl9W2i6Ah1+pfN/AbcNTnknaxN0MsDZJeROT3sPy2qea
W9h3+kkvIqr4fhDXReiTlpYw5QX5GlvsqYZvNgqAUi8lzHKYy1cnpDV8JqjXlqsG
BgtkZsnt1faH87Oo2zxKwOuaT9uoOUq/VVveh+cyqGVStjKWDZdulC4Ay/H0Pnbq
yde8iPdXTX64tTpM45BVOg2zyWxCgGx5bk9/vtvwsTpLoah1g0LOez9XPB7zb7fH
9wf4cZYMN02BUk9MftkPzwS7ruCfLdP8gvkQ9Oi7jlUwsDFiluhmFve5AyC6k/pc
HnQRRhphIPDiYaJs8Ow/0pAvg4cy4Kyuiwbwkof0arJjtFhkHU3P6OTPxoJN/yXQ
2d4oWRZykAuVMtjxjXpKxaZjT5hNGVznF7v43Ok2fqTho+m4kF67MdVKuP6Ha2Wu
f+6b4odZtC9XKWUIq+WcBTgLkVR2tK5Yy/bNkZ/2/Lv2UVlNXZEIXp5WKorf4NkR
J3GnK+eRYuiyAO7XB0xtNw2o3UzCdnCHkwgwlCjGiXFndYs9DjWUnhoJDwQXic3V
WJltod6zPHbeH5mWssgOUA1bTj/hJYYgDX3//flQnAXXCMmNppKxnBa1PlGLIl5i
YDWnAhH2CpaW5Puzkl54Uu6eIoKnBRIb13yK26INg4shtpVqctWhLw1Af0a8BYbm
TJ9EzVVOXrsdB3cjCrAqUNabA0xza0iU6CdfmtMmk8kgZiUHSPUjUw28AD2hklt9
cH5UmrhV2BgmhH3JLQ0UV+Q6z2cG6sfCFuCxLK7hCvIXQ3NA4TdM7T1ntdFDftch
yIqfijs4xFe0Glpo1SklIYgcv/CJMWDWh2U2PuzoK2TPCmcfpYgUNQd5AIt4dCWI
UOMuX2YwRvj5I+BDxhbFzGwsUVKxQo+qA9XHjWjmHtK1vH8fqE7bAglFzn6iN/iI
7MXt3eBraJjdrMtJNUCe1uDwJpEPQ/9VkFb6y183S1pXJDbL+Xjd08kje3HqQdyP
Q6aorqB4Vi3u1CDIulihYOg563nJJf+b6S/7w+CvJNKuyTZdaCEetBXd3PJCdCtw
zipIyHqj7kqVqODi+oxoRuRID/zMbtGhSCvUn7KFdjJSUcEXyqYh0NLTxtHGVRbx
Rwl5RpiWW5VbjjmEoHrqfma+IegfobreDyTi2iZa8EQAG0TlC709cEkspsFSdVb8
3Tsyc6iMQ8I7r4ObboG3j8IxloLXPfKVxIpFYSdr+JVpC/g1GTK7loJadc7WIWsf
FYeQCSI+qI07aKCZb6VLcNA3UwN4s84mPDbsF5PnlTvMsV6NqUDIeXbJyaZi7Hbf
SN/nH5CFlyQUK2b/1n+6wdCePuzK8FTNBh9moQMLDFO2QUkebgrRy3d0ilyeSDoF
k3wqKp9gGcdG46MwHZhsQVoc+Oopq6Efm1BRAUj5yxJGuZDCRIXW/XWTgN68FkRL
ugUUHY51lD6FcrREWfkrnnk9Mr9bYzxIFDd28hUadTtKTFH75PL7LLegBwdNgGzq
J5yYWq5CwxKziK86XNnJMlfHVQQCjm9lSBMbAnVG1yyluNkqMhxbrvNmbX8n8Ota
gFPAAjrA4Y0o5Ok3L8YpX8MWPcMuxogHeXz7EqvU1acxXJyikShhfvdGkyNSk5ea
pVXoA4WZTebnvQsQrrZMgGadw3Ioixdn6bxPop/ZBc9JtVIvMnkz5aVCRP0/2mV9
gAyuavhHDZnal1ikl4qh4eWd3/5WVrlEtxzfQyLNlKAyLhhY2Z5rzjfO8Zpug/ci
Fo9icpsZK1ralhjg/syufVTGL9qynu2uzR866IgNG8a7Fov4rcqk8Vrrwneng35S
wd1WrlTBAUbTXuwT00Zn+KA3jIUdXo3WosxEceDt70MPnF/EYS+RRH9iV5mGHLbX
4xeUfJwcxmCEKIjrMjJsZuv1EMhASB7qCxAFej3igPFNvNjh+vILW1Q9d0a2yHCW
0kPs+kl7NCu/nC26bbX/ri+Yrx14Eq5Cllaz429/7dlUYlFmGaBORk8qoBQkdau+
p9p2QswK4zO6JhwsZnTpp9G003Ne3LPifZQ7YkW/ydyaGuqzGjwb2fxPMW01AAsm
FVJd+3LBpaWj6Csve5s94Hq0kdt64WA5btxfgckoVgmbHpGdzBjbNuVqpcnh2ZHR
JVTILeEMHo6ofatgIvumUvlZMssLXKtfRWpUzHHMVw2wiiGPGOYndi8DovLc+wKp
dOy/8550djtBOSZOB7BKZn6MtkF1WvPEAta0TFhgMwqD4ei0ucw/DWLl80sahiHm
o30BN/yEAVe0oQDqMn+LTfh01lMI2p3rKiB5nznyFaxYRXlH6V4fFLpaFy1k5+oc
CLQVx6sq+SZ6T6+caAaRVYQ/FiTaY6gXgc0oqZvPq1ergSu4DR7dKYME60L/rZe0
/RxcMa5M5xc6ucSYjjEZtQUnGeW2DNjOJNTKPvANhK+GkIzQ/oEGrPiMvoS/399C
ckD0ChY612baw3IrLiALQo5UMp74ccTu/PZNXiRyD1dyFkT9aUX2i2xGAnUhfB3F
bVobify8azxOkPLc340rj/zeOyn7hr0rcFuZcQUu4fqwLQYyHroIEAGvuRB+SfE1
cAjUl1CjL/4PEGDIgx5jzDDJwK2RXHiWmgCo8ujleuqqYP3MU6S3zQx7RtEMx9PX
/P1rrqOY4karp8EvOhIzrWuoLmXxDKQ4Zv/tPLpi57KSlQyaLY7E/Ye9iH0NKwVp
B7cVoFGEdA3IJrl+dYIPTMw29s8l73VDf11a41FhlAZ4G6a8BosGFhwC1qHsqhD0
LMxMKxpaZM6t5LZPA3M1TyR/ePhywfMbb+lLHXGkMRM15fmUyQfMs7Jne+NvBkE2
4Au+f8BEbbbnLPVFU82OYuNbfBKbGd8Imm4uIO35JRt5Opy4hYUkZ4yzENqHEbg6
U+B7jsaKtDeNwfCQixhOcBTeOSq84r73cugnrOyAl6ljCGoMos/gCiI3eBpwjlow
oHkzNYjBMFpV36Pu3NGx6skxFvooOMGkIjf2c+sxhLEmUXy0agYY5NhI3yd07Q3Y
xSCg9d4kZbS0QmrwtfzBRxjv9zH3RdnnBlJO9z67cx2xHyk7hAJOynJ4oi+1mhrk
INPRVjIdyHSDxBFzLQY4GlvOZprv410qeUDWZvWGyTYcw3UhlzOHJyQ0hONo3/Dk
pgQp7DjiK4DZHTxvJCxebzMjEImwR89TZRqD9R6JN3wEYRMvpOxYuU7jwKjoKkxO
wBCWu8Bgf2tH4W77+5kZrpXwjIm08DNTZ3VtCpv8VSM4m/nH5ZsUaB8M4JmeEQo0
XddesZMDc5WZXHr7QmuMCbFvhHR5V9PcJuA2BJV+JcZh3o+Nj2JpaU/UiPU0stfX
tGTshL4YSvrEPHpISPCRfKtQhlq/pn6uSaiFmEzJSZyGqQPgDrL3UxX9Bl1uVv3z
iUL0hxgKP6mFZrzn61Ser3RTULZ3Hxq5ZfiOUCBXrsm7LwSXtndpakFDFh94fVwG
+RnGrDuf2Dd6aHemgUNhMk7Wda5qjrqSDgwm+2kzWcyQlmoFrjF/ur0R5sE8KrUc
isWsTVTVLZC1o3rREx+pTBHa0TzsEFhk4EI2y7xck/WlGW6cOHc8luaKDtHsvPF/
nJI+VOpC49mpIaJ4bhvIbS1tpCtfu3en2W1OritDIhmQEzb/1w1Q/CCiRrGvFBga
BC5dsuhbFfiL+Mv1axpGJfW66a1kLMZWrXi+9tEFbvUBGZpmvmQPYPYEmoPp/zDv
n70OTZv4pRu+oWkR6TY37zFvYERwvfX1Ooyq8u25HsUp/miXmYDFPwPLIG83ppRN
WqXcH3noCsktxtHmnmS/ua8iGgsD7MhmtVTXt0KkRc6G0Ebmhp7O6medaMQmD6l3
++nzGnwryBNxPMqKYRgcMhIgwXbAZjL/F9g4On3giSAjBVyRicugCUlVawUNKaQw
WXtbDF2Qp7vJmulcVqSMN7xhOLIJLMV79OEYGgw40GOW0UlVg8kLiArxOMnTM4mv
MB0FGofXww6NU3bfEUZna5Z0h4hzWoprPaY3FhrHeZKqcgK2ISnfYXVygrdVlYd/
9tnsVuA/ghOslWi4MfV7kapKuEbgTL/IKEpXFV1cBAJXprRHNkGhNUBfnUfQQzZs
YAOt8Nkr33yJBJ33IZbH9kNOX0CbjdASn8FbxCil41xXnQijIc0vSy+xGDkNPSsN
t4DxJgFVU7V6qyA3MxRtRaikasKOEBjNyn6cC/uxQ32BBglyYEcGjW2lfkQNMl3/
wmcIS4nDbQy187t1shdhZh/vxD+RxIRCQzu54fR515my/umqnvqmoTYOK+yS2MYV
uIBcPdN9DE4VOilNZWMyEOls1UFE4EHThajcNrKnjZHEsE4QrPzSXan5qns50dHv
Ln/mMk+7a1rWUr9D3GckJ0JUPfVPGt8qW4n7vqFDOBDnWaEWFA8i08oL+27du/aa
j6WLNrcv26Y6bHJGjxzntC+MaAXHRB/a0fB2lYJkYS3htmI1kJJSMJXfU7GkANKT
hKFdRhV7R1MbXXtiku9dnLxTOxlEZHfanFbKm/xuTkYwq1rkJSMGcERqyhMm+PFe
SktTpIgUslrRr3TuOVht6/JvynZMQ+Y/SFXW0w1k6AKy4wro6OhKmGNoY+jaHUY4
lUR65OqWE7b9nsXAHg+Ky9QOZsgSAHd3PxK6Xjt51VNNReeRaGJOlqxePj9zKOX7
iGxXSgR22yiFm7LbLDtkJKRwcEp7wXgw/IB62uS3UnkirsW0Qf9BBasL98klksnQ
TvSClzfnIUZ5hzou21jYHWfK1HWuwXJdw4YXpWo4cAYyzX8vdSXd87hpOFjJ3Qdx
pQ9k4gk+eQ2buIJ7L0ne4b2hEnLG1uEL8M++btz8b3a5BC5mZi3HyVff3lJ7yrUZ
MCnJcq8cP4Oub5sUUkoYZP8+ORr15vdpptDqo315JnYEXMwvtoKL1RXEuLdZWIAh
O/I4gkpMCf7z2/bV3DHiz5khlmKHuByNU6wpTDQHHKfi8pl6iaFt2z/466+X4k+N
Gt/bYJjgRBbocpQvQv/wKg31s415zj/5vCBOfD7/yN5BcOeL7pRJpR5gF1fNkPTE
BgKbLB+s9TkSubCVT/BEJvu3kPIHsdXMBUCbjMs4kXEV/KQMzN9JxSJKUZIQwfmh
uKYtp+Qt1ao2+nzzwlAl0th9GpPFO02roBg/ogBqaxowBJS2QnBTnvVg4TfWI6Jq
B2gIpuzDIBEPhII1D9ZT64OqXmtjqGZblS5dHesTpAhCj7NZhCaTXCuJXve/8mFQ
YkiHy2WwIItpfhPvuIBZBfZbK3cggwbkuL+ZmBpKZctsH9Y24df1g11f4Q0L5Xis
yij3JTT2U5ZnB56Ui+9p7OGCDD1QOQ8bdjenLwf7w9i8T3Z9t7E0d4ctxWJ1XtWx
39uyneDwg1cbCvkowf1ohoD8JOxPQqpCSesXzrGs6XuUNNMBaHEuoimVsZRTkh0u
WP8qR/0DH6XCrG28qGuJm1hER5nvv+graOI+CkfXDGyeMlRo9nfK9o9c1NgX1TH8
qgs0CaB9D/OkHK76J5Pwxdp9XFUh1sQYE6KQtyUheOkxLegCHaFrg+DxH10uoh/z
5/+p+rnsaQsCbsICIY6Z2WtnIHFTfdhTIQj3UTiYPd74bZL9jGk8RRfxLyE7s+Mn
RMnJM4XGtAYaxyRoonyNh9tQCEWDzgbKvenhtajE5skXHs2y5MZOufux4nOqSrQj
igsYyZe4E5LF9MPW2UTXgVUASGO8wJ1YpbTBsy5poUid+6H6VlEQkT+kFBZtWCQU
mv+zH1cXdqIGnuCGzkr5a8pwGDZjXDfSyLkhRAGEcoogotA4uEgnq7m6pgLNP1gR
NMyrO2L9lALNOuTsTusyj3G6cBynKfSuY0MpjSQ9qVd8O77PMpdJWZCnXszqIRlm
pdolNaDOMV6T4KtIDtm57z09DWBYoXJE8GAUqFwc8N0atZN/KDOgUdBT+ea6bPYn
0t2EcO0MTKqJ1YtuMwdGm58tBY3IdFx9FHBp/+cRsrS6UUd16j2H3rvT9rcfYiwv
l1Jq2kO3nJspcy3mH3HTWnmUsri6VvNQ8mYXZibPVV0jhAe1jOYeUEYjxVN7RvO8
FCl3/laML6pqyHcODs5/6J6l9Fa0dERzj2EuTaMMveq01dIK17ZMvN2a3ijeUa7s
hJ39f0k9Br4pp1v44CkyKoJFZPHDxfXKqST9XKiWghoycdZb+dYy5cu4y6gvKH/X
SefA56CCTZx1hrTuxGCMCo7YFkl24iBhl9FbadmBJ6wf+E4mm2aey/Xq+QlHvt6S
wakWLVCYQoKyqCrI8axzk79rzzXeGfECdrtHkfPRQ3AG4GFz/Yw6unrnJ/HxBrBc
yYAYGJsb+z0W6e/K8+w1FoApVjdALgiULx8wqQAvI1+qCeOAdsGbLYIJFtfgg0Ua
jN4BB9Zf9yGryydlTS4xFoGWhg6fMAYTLxmULcD4mk8zE0oj/nOA0OWFxpOBr6JN
t/z3dfFNaD/aUUxNUOAj4vJPk0UgDZGzMz3pEKpucqt33u4NUAseZnmtYW/nwgAe
EG/jlwQtf/MFPQTL0oMwriZ46KY0FEPyLOOAXhw3t0azsTh6QAsga3nu8vCMCwaP
E6Wi37o4ZLSoBiZrZYpUE44eNRRcaEAVBH5QBaSPhNRe7o86U/Zo1Ps424/DgbOk
rYjD4ilHU477c9BwFNq7XLjphRxTXmdXJPCb/noQjc9HK9prKEgZnhUq920lgaMc
WRCJHT/CDCksvyeuAspQMOR4aXRJzsB2RQL0yFl3A2yNfKOwDHjhc3ii9icVYpDM
DkcX4+TTJ0zR7T9yO/zsHlNJtN1Bmi/+lmKndAQJiPwqGuUsORJopwdIHFPWz7eD
id1GnmbBh/4Q3emvN97Vn37sp/Qy2Zuby1izHLN1di2GKjlIX8/8PKERJOIrc/p8
glnW1Xlw87AcLA5VUNhbaJ5e/3rMkgqiiuliVD/pbQmPmjB119afenceIjnGre38
x434skGbzKxIpqD7gVjCq8xtJgwuH/UibzJEd5fC+o0TSZw/KffFOdsP3yp01/th
BbckegHdr269VXYGunzNFLmXZU3P8AIcGJliHvJ3sG51L4WKQQvOR9WZOiYKUmpT
L6bF5KAgsyuxt+s+beuK4tIdMiyPPR6YyTZ3ZhBI2gVKHV0fQseP6JDRSo/vd0yF
dJiDAUwEpzx7Pkol++EdTTQBPk4N/7GqhaGsvxoe3r5/AmVOgqiEC3OwMU7T64nK
+jNggESOwf/s8hmHn6lK1x2Dwm7T02vM/3J75Kmk/LYRYjmH1ChoClsOiTwlhpOq
3i4Azh+YdVqjl44ZbNJcdg7w/7HB+40C+p1Sl9kq1KgGbzISm80fjGKKowBOnriP
sSy9p05UlcjWp2XgM8OQhsoil863f4OV8stsm64ynrgB2iziaHAwPnJHMj32W69J
de2D7WagLTE3U0wMk8i1sh7dDzLB8kkQkQJxjml858xOu1HBK+YL1K8Bd0D9PpaP
yLp5TsmBaw8WKkaxPZDgsyhe1QtNNbbllRX3gLoVxZTEtWh6+k6UUxHz3FAFOkVn
a0s/F/HIgiXQ7wkdAKo9NSG3AdwZmsBGgdcSf7+yzq2MvB0viiyodyRd+lHkkjPc
yQ7sCHugB7qPBke2rQVEhEhH8cZmC/AqXE5H5ngxDOCSykMTr/onlrOVpHiCZ8M5
DOANvt5MlWjmHIuvc+LEP5s8m048n0OBp6dQ+YU1kn4/TM2QzQc0RD2YHjo9p3la
QlMmYsXMAv/6shaSbDp7iYA9q0ZjOPdLqS/uzufQnvFNbhJqLHNIgxUVRMVYgrNm
DlAGIwYIHycj1Exv5X4PB94IDJpZFkusdwzfvbq5fzQg18JXNmIWAW2TFpM1Z3yU
qv/VwlPzsN5RaVhjk7ixJ+BB00Hu5X6EZuy4fTB+fXNyC3m42p+/gfKPzjnTGoF5
uSoOVRRwMs81o2FwjyLlhvq1swqxKuMRJsigDl9JxbAxtMwvw7LBoW8rAO4EP5oq
gHc+4zA6nsH3QX8qBCd3xW/qIzmPPLcLDSC/jgdL08Fe/l+icVYiW6aD7mrU24z0
Cx0ZxIJVlytGG9cgj7If8G4MICZJaYQrL2ojsun9Hnc/8hLHIZPJ1MKtLBTdzvgs
JNsHHagYAECnot6Pxy6w44Lmp1dT9HuLyYPZ3pdgA+fppXKMPHYYK95J/KLHYXy2
Nv5jioD5USZFaEVZ+bnRxuyklRTswhCQoTK4of+gr/DVRohVEnNTOTDvsgD6K7il
36KxufTvSmgjjMMnVfS9RUHIUwLsKHijJc6gEW0EFeQQfVAtTQCUzADsOTPdfMrO
oq+CnaMGpe0OfUEkv/P/46MBFItMU3L/Gg1puPeG/YE0nc1t3ahRhb53bYip2g0f
Mb3RSYfaQW3oaCmMbu7J7nxeV8g50v9CuAqWQnNY5GR0oVNZ5LP4H1NvcNV0srA5
aCZ7VFH3QjapKdFnkG06TluWlmmw6OveDEWZ19nfJ8+k5h13LfOtQxW+NyoeT0Op
o6DCQ/DaOC1/r0/bqQT+l/XGX+Pg9GUPpRxTYUVghdcnIC7+BAIjPjQ77d192EgV
Ae0zzEXMBoa8yIGjy/RrAcWBEIKJsrwCCuGaPFsvahPuXD0jFqXHqOcpG8zFa4P4
ODiB6fEYlMEdPQ1aIqCJzOVIL5zmcZw4x92Rq/a5DcWj87DxK9QKY2gN16q9RU4t
HQVjqwugKO7qLp9lOuuvsILXHs39r9i6kzpOqDCIyabLFqwNArWLzinFXgW52VgB
b6JQ734fM3OsTOmNZ4iFNDDXOOWw/FzjoTnCMQqCcOxSxTrCCVVjUrDmiz+UDTUb
jJfoTJkUGP2gWzObewFyyDxUmoSqNzIijNxrqrAd3r7UJAiLzTO9mKgfIMGI+s6U
iBdFtPxm0ncJ7PPDFPW8/SUTvipapoGL5R5T59aNTkhTNul2tl/k0lpMlq7a9iVF
KK44wSk7lah8w3sUw71euywR8MSYNhL1He7YlnFHH2xqJq6ycNlsAfq0doliQXq/
FePdTl44BBXJNJUI1J7U0+kn3WpZQC800s+wdgxc6tzaDtOT9mVeDWGwDAN8L4Bv
KurJ39+AtKs17H7pW2gMk9qz6AyBW7B76b8NZ8ocBrIho/w7+m7Z0Ia7lBlETf60
dMsdK9ODeDp0ZJ4KtrWOf2Tf331Y7vIyW68t/P+EdgW9Eow+8E/dtrYZC/f3oC2J
pt/lAxCjDZ0338uNar7P6+LqGxxwuEQtP8C9nTMhnrKOWz3vR5uYhXlXkwoHZUoi
wosKsGczRwXIlD9+jYl8Is5FTcZuORT+MYoYez6yIZ90EbqS4ra2gHEdBwDf8qPC
D/Nz7AtssDbmWkZ8vhtNc61vCmUvCouBdHLxw9Qsszfu26CiiR3wZz2D+jEpjLep
jsUCuM7t0h0t3p+uu3uWJtN9xg1MK/AixB+aFiJ53Fo5VPlRtFM7qFWO4xakg0Rd
QOTcB4z9qkYfY2b6iu6iUodpx6T41X/QzmjbLOdqQoRvd8A1u+6B6OIgEhiccvSv
C8HAorKcljKgTw41gvSokqb0qZjDiYysCO7nnyx3BBE1lDY2CMdpuDrBlLo/L/5Q
kyr3jx+CDKONmYAFmzZTAgLCCIxrz/cdfZO2RBio09t5yfltDfHU+D48lPXqK6mJ
2SZ9SJV0SP6wY55ELnXIbRKgTs1KGbl0WIDsMtfolXlbjBJh+QKN5HdYPWN7JKzu
JxYMiP3O39q10zyYwODk2d6Z+sEY7HXYCmyGGMo++c0v8/uhjAsg3G44WvL9EeR9
uGyLwvywgqTZS29kc3P6cPRxzG61vyJYu5bV5YlMYNu+C9vNcUzGqVIM1/CZcXBc
phIMI1s3q71xlo94O6gXbGGiF82l3UGytz6mwHipLFn7e8mTrrIF60KjwZDfdzu6
pgWYh4o0PVtZ8fi+6lYp10XH7sLXHAKucAtHLStTQXGXwTBbyhZzs0ebg0cNj02z
jCeM2HdUCOau1lkIfbqek/fEoc/wtJpPXkJe6AdQRPVtUD/nUtC8YfiubQx+GtFa
AEgFdJfmqBj/SR8Xks9eUkHwdlm7zr5eidcyr5SXBRagNJgJ40XhNqk3ptQCLBLi
Ccy6ej57qy+yMNoOD/E6gzh+r7cOvGnHcXwokWNZpvtj6jADTHMYEIybo0urzMyn
84w9oMzlzUikwzjzBpKGFw9qSqo915VUxx1/nLPMh5dLLU6xdnW9IgzfMb3JT1CW
r8NOL35ZnjdixZLTAH5vy2Enb/JDSo/4Pl8M5Xp7tZ9xmioa2wxIH+44rZkdNjH4
bDfpHEZHblOkkDcU5syHHtn11DBp8OE14O6jO/xQPg+KdH9NTkkKScAmrQP6eXQw
mLUosBHt0qkUiD/84xRpFT3F5nTdnlM12WQtjBdP9zJv55I3OfG0uwAbiPh6xSQW
8vRpTY9EVIZT0IdMzTgVC0dm3qU1MhkEfHfJelLgXZMIyhRtDb+Z3+a84yQvQNhf
HdMW5Bclr4ZSCUMOgRRbhtbdb4XcmG/Xi/5oc9SGdGeQ/afBt9KjtEZ+sFlYYWdO
Fw2COAijUivqeQrsvRd9HIoqXxViVegdaQu1KhdCpioLUz3S0zBBk8zVbTRVZpK4
0Qaf6W5ZCe0wBTXPKtgyEza7umVFfupwzrcfhwXNG9mLrbQGEmVA7ePXJyVYnDwZ
XT2ZR26b/Xx1W/jsrds3eyE0TsSB13vq+KFL/MW5BAVNqG7mlYmrNMdhDtV891zI
jEsFt1J613GupK6LErJY3TTTf6KwJl4dqircBDUB7iC7Q8T7lLdmKSnLzjeoEske
H9+i4XBv5r/CYtd3O3JseD60vb4W4bpMmLIMw2Hrvlgz8CZ2BZxzkMjVPS+WNL6N
ZT6r5QOuvNI+DrGebonMFvLUapM7xsVh0DNrm1W5HUH8QpR8jLS6Zt3Fz/jP321y
OSVKU9ZRDLWjFHSI9VttZZfDGv6KFKg8NmvAL6OGhbrK+Cr8b5RAOGRATGkexYnJ
rKQa1iEar1cjhGtlb5DXNNKGhzbCVTMRfbZKr2oXYpmhi2TbYJJ1q2hR8j4BSG1g
Z1vV27TCmHz8KeiYgc/3KQIhTNE1N4xJTbg1lO3WbK3hWVePrdPFlKMW6pOMFzwO
bKpypqzJte5dlNdZePMGBEMKwoz+Em+g+wIS+iJ/WkyUpWmvnWR48zwZv45+N1/N
SYgdkUB3U89UYyuEuoz4SkuPEF+x3L6c39hR65yyetP6FzJ5y33KgJ/0NOh9mMjl
UL5IMDTyLp0Z2I1BNHU2kFtv4F1OZfmuq7Am5j2q5ADtzdTCU1+mxOvtlIq4zNiK
Ec0CaN9ohCEYOZEeiaq5mFGlp5nmcqXGioL/NPJEQaCAFYhTVXaLGspM70k8h0+G
70BNnCesm7/7A+BPwJWIWXmkRct0fxMAgTOFmdQxb6JrGJ0NOsA1uLG+ARnQ6+qC
eS5ZCVq4J+RNqRKKRE1Jc6EBBUFd0zc9pi7SG+vpRip3FYHgNFtBChwNvO5udoBD
+eT+7z4iRPM+qplenPqI6qMwItd4pMgx+VeG8WWl2LvAg+rfVdMfwontnSEgJmX1
SxGBKqQNUlqggZYKHxoK/TiDtYg+lTQopaEIoBYx9d8RJzVe7V2k/dPz5ZDIXX3E
TMN4bY5irOeMDVYDH+oE4+SmBOdOMkXQzl5BSJbrdQD+okufPSlldhmgEsD62X6n
ckrk4JdhhToTlqa3rFSjfpewI7+BiqmeQ3M/hurlrSbeBc8zsyYAfttk4ki+JOoR
YJmh2e3JtAjc/PAqYOymKVWsaILQQDzm6EvkjBD2+txIvEf2BvJotWgDmzUokDwl
rdgSMESqi5YC2YhZnPwt0VL6QwAnpQR8fNe+jMDHSA9dhXVcCLdhIgjYl/lvsD7d
DMZktvGwOhNEc67ua9Pdtv2g1m0+sraVqYFBsFQshdHzqDCmgWM4V/rye5cv2gSM
J01Svd/h1EsTacdyCbk/EelQ3QhUsJCpti6/27iNAeTLqEjnEF2Ll6b6NTiNJxTG
DvfqFvdQEGmvUV5VWFNDSEXJFcLfyNFOKkQy42r1ogTdI+4kKWbXVkZihmovsMoD
86ogbebzZydL7AoF7bb8Ncm4J7JpWlePpjOVWsO9ARLy5jjijOHkiW7L/b2bX9lX
SBXQvO4ULnJDSX5XFhSHe21WHiPqfbnjuQvNFZ1qGPiqYJwKUb3QWjAxZL+sKxYE
W1/GM+zaaPMMs3pRYnE+Cxg+QhFUjBP0/Fq4R674Sk2IViBBMW+GnpmBOIFPSgza
BOCiTvORbDk4Ja8N0WvP+nSO8xmcl176dBndGf7IC5cxs7DYbQjxpZarTjlpHImL
mI4fUAY9Gat81ymZojnNeirJ4b7lUMsjOo66gGcAcMt0X15jWhwy9suGAfxMtjRb
JpZwZXOu28VMQ2idrjJSCtigbzqVBd1LzmssRb2enACYVAN10RNjjf0b+tp9JDNx
1Z+h5ec987XL+W7FqoldHibDw1TtL09V2g3bvCwIYTBxGWOUL2hZigkpGWhACBnO
FCUFLGy2jfyMori/Ouyi0lz0GPEH4U2RSa3LmwOcAqVDAQG2G3ZFkebZG+8UqoCs
CoaVtZW4fcI8cFxrGJHj7JTn3deG8zTkx8F0oPuPMeRMdsFOzVRafcS2Kokamfpm
QFLBr6Bpo6+R/xKvuKHGLuvcWSc68kW5Vis/bhx16pe1bpTPlM8TJz0dsZbuI3np
sc0oVpadjibKvb6q47mnLw==
`protect END_PROTECTED
