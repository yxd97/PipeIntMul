`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FnPXxH+Bv4W0ykLPklmry2yH5OVyTLc3+fdVXJ59YMZgBcuoyc4LHfe6K/mkVVW
rN5AFTfidQMea+CceUjYd+RNzpm4Hpj1RzbprMu3YDzg+uIKeiHT0jDTRC7iwL8h
Z/v3F1+gKIVJjAd4Pxdqeha+8jkypNAdZH2rMIA28cFv4k4lE2rgjDxEtg+Yd2Fn
aA5bCmh/5xgDya7ZbOSGEZ3kpoeLdOPUb4kCj/JmhOJuGF87OtNkuCk0cHnSOvjq
res0h4NAFt5lWYETcsx/Wd5N6ckAEZ7EMHQipY4cJ0S4kdG38nqfzsVCgFRkubZQ
K89LvNlIJAw9BPabFEw1s09NChRrrKZ7pNPZMEZlyt/NAsllMn0StkU9jy0F+lkq
rZDyC5xfu66hmHIlvFsyfZc6szojhu9pYwgVzWmPaKyitQRPK0q1B3f7iYmLuFqO
kPKaB6NoP7kXrMCoQT6P2/BWB0m+j1MuXoFmsmuOGXY7Oy/822/vz1mkiw7+hr6H
Sq+kXGvuAfTLppODPSq2PB7REDEiHtwffbcwaSZx6sdTfTVIBWqv8lb46wZbVh5w
UhViDiejKpkUt76clFQtd7mEPz3jRKV76CFIa1onWsZfCNf6NgyloTGbaiwilJzh
1+ixRpzh6vCm9jTvueB7+79fjvRiZFyH+3R9xSC4RX7wIbSCO/bHugfo5hd4lJn9
7UdE7dS077H/W4/3sqa+amT7WIPRCw++qOlSi9CDdkQ/5z95Jm7AW1kleNqFqfbs
e6PfcpRVXJM8/oZ8vkKNDkWGFO6r9qvM0SubClgdlgAvdleCTmQvVxUseNLGDI9J
vTAOFBzHTm/NWbw2bleViW4otPyMUKAEfHp0FxWIvNDGeufTTtgvt0lYdCuYeec8
tsaDYDwJYXoDoGZBQZCPRY4+Gxiavlsuox8eaAmC33f3z84aAvBok62j4tmIMpmp
`protect END_PROTECTED
