`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Llw4+p4TryMOh4aV9bq46YWKijHB/LFWB/uIRhRptX2TcOMOih4hbVdPeqQYbHhQ
ChrO69WgHsLoKpkktYi5fKZ/8Lt1a4EZfOuEdgGWLZAZJeMVeLqyK8eRLm2Ouplx
ZYpfNI3J95gBKLnHg6qjYALjg3RpEMTV6UQhhiB2Yf97RYeZYY2liJYSpTkmFp91
q8NfMwwlV1HDzqRJthlGKNhEryh+1I4mj2CajMOJW9IdWSDiIT+DgkOBTol7zDuD
GoG0NWNdtX6KI4IFXhFVvbtzadCGtJLw4HqOs0SgrpGUD/QswrJATfYMSaHStdXM
y17aM9w92qudFE1wkGz2LuGFht5MFeT/vV1opSBT9NjD8gkxybnfYAd4jEZEhoNP
OLcWiezkTUxdK9fd1Ank6bdRnlaslfRceLNwW9+HG2Hihc6vquctFklO3DGy1axa
3e8dnikq6tJL9dwosOr9FRnk2ezQMUkcDuzhpk+DJwqDEHPLEfhK8HfZqTem/qaK
9xAsqcu36ieGhRULH+bi9yxoc07Nkte+A+k1hVhAKxnozIP50mLU0dLVP9Exp+K3
6v+8cGpwFoIRBFscFsnp/hYZ6lKWyiE8/aW550ANkt0nFDiYnF2GUqWfTPefDyyB
73P2jXHSlVr7W6MpT5ji0Gf/0HHgRaT9Q5VnsMkN0YbpQmYmwr0CVpbLFLb4U6pj
hZaFL6wILwHODqNvH1SptPC6avqHVqqGAh4yxQ3Bfd5U2m920Sdgqa3iCQvx6QxH
KQsv56vKICJ3cI1NqRcmStFAKjCoiTo2FuJBEB3wXgVDxj1AlDy9PSOoGiazmBDQ
As9eHvvP8rmdBy/ZV7tBx1K8rs+p37sIM7RP0OiVDfP485elXVMdYFuUiAt70+FF
oaBWqjjx3bQOaTNx7iqzdniq3zAey6kDx8IwjwOQ/TMtpNPWRl4NcFEarwyTGrEH
GA6G8l81EKsU4qE96RKZqC3RhQ0uQFxYjITys4GPGPbSRGhxbDlTgStVQOB3KMQx
urktCEJhWwijRO0xn8JRQGshT7LRYSzNcKl/GpbuklmgiBW/DdOWM5a0OqqB901e
jU/rHeIZizilRjRcXqJetVi5d2hVKlpm0d6KAO39hjEsJvJfsmoNLW466Igc2WWE
BOR9CmRWU02mJVk2bagnq17L/VQ696oYtTMizrlX85YeMpKnSYG27U7jMdEryX94
vYQhA41fEcWivkyYYossAhe4/fd4i8UfxtgcBH8sUk8r+Y40Cimbt3463j0hiLz/
7ZYRdxJh2uBW4va3YHF14+tHUygv+A2g1DFUGFiB2766e8rYuIu+YNH1rf62MpbR
Chdyz9G6L2fx8kqWRJjs0QvXED6DV0v6Rx3q2yLrDxrJd3lxBvX3TWyr22U+H1+S
QGekhLgcN48fo6U6flmmQF8gkT739NCFR/sm4Og5o429GO3W/szZBjzfW89Flave
UFurtIfjahobvFL6g64ZcWFn71Kurgz23MweUZ54QyHuvXr6hK5M6A5aYv1l2bHr
BbIsVykHoENMrXRPyNIUDu3w4CvDa+QhLv5A8ZGHprAp0NCqzZuOgsld7JN9FyYE
oBMgPIFd08Qdcs5PEDEzt0UtG6ntXaA8ZU3kwskhgNqJXV+U4wkjFYoBgDGNZ5LF
FfOqAPC3xcuFZ3Udzfjg8PGxB54DWsApTn4JyMNn0APZTRCpQwyrUbkVIKMWk1PL
nHSrmslW2JxHfTBQjXxcRqOSZOyy338sMgh3EFGWFGtbA2jHXjNDT3vkwcOlF6Dz
+6DV3hFAv9opwp2UwVbZ7HO7iDlUS+4wKrhvVwoxYVFNGWAJ/77VNDeA/rcwAGQp
33nq4JEj/UPy458aZJx9o11uTx7A9hyj1gWg4ku03CxjtfU4WTj+cEKCSkzZMzqA
5BBdcuJLORaqFBi1xyTbpKa/7c4Up9ihFs4viY3iMUIHA5GBilVdgAkWlaXc1GwA
EeQjneOXto6KWOF1nNFEMgh9tlYVQQl+KBD2lhyT50gwhUeTwsjD9/EwNemSSdCw
d0R3x0rWr/Zjsj5xuzqzNN+cMboOZgLh2ZPHxrkX5IGm6GEqxODXFBXvGiE6l3Pm
okFvSn/UTwgB4iK8sUmAg3dlIV3kAlVzn6pMrrnxUbgyXoIq3AABQQZkkI9zR4KQ
N2GOYdW8Cy55hMSWyCoKqZ9193Mma3MY65FMiwGQXescTbudwkLsUtK6H8puACge
tJexAApnacnX7kU9Wl25oSn5uTg2XquWVLBQgMzbYGQBv9tg5BGpOwj1mpADwZGy
yIXFRCRkvxh9N0e16yvUQUzp19B0MrYZWMSIXabR+XlcSNUn+51zgNaOrSVYN/5k
MpuLuW566SdJim+InpQUgMi0t/Sci1p2Uc1ExbC13gYnDNZs02YJlN/gAt/lFOC0
pvETpxHe6UArMO+VpF6m2y792bBoEPahgAo1HAUNTmlQ8IKk5ECtIvwV5GTGATW0
yNBbvhSZArBbgUxgkUfLw1QXc2lhgSaDwl3UATi/9lmiFNOQ5d7vpT6/Pai6wkwm
hYyI3G1HSjIoutcnzYJT/r8i1zWx4Kzvm674bO22+cqPjat8o1uK02whmkbP55E0
5my8QahRnyUZLSWFmEACwQK/nCf2AdjXoEgqHlrCFzlYe/c4SB5XvaMzQ6seSSV6
XT9ed9WSlpqUmkArQAhtuL9TYZbKD2tWWhE04KHEraQm36DQs4DK346LQi5RfT8b
c2uBdjgwSlWYGz9H/r4s6uGrAYlN0URPxRa6y21RrTyu/XhpKLCobiNNvW4RbnlF
wpgnkqngff3FLYzyIFkZAiyUZKvAVl+hVWk5aF8WerNfdayc0853c3olnd54y3Fs
sQN6VlK7BzRvFs/S54Y7zJq9EaP1RKxs5g41HwBpjQcvbC7phawDnjhvP9O1Z7l+
P7LyrvWV/Kvy+MFBBGF/enRiatRDuzrlSvsLctNGw4NPauBYs8yS9W10bYWlkIdp
uPloQGMbLyubKP9J/zgLfDolVkly4oANfqjDBVylFgULGO+5znZG2viA5DKS2QHF
HHzPP1v18rY0MG0PwX8yn98MkCuLje3oLOLcWaX9tU/Fzs+slBJwmB7eF+N+kQCm
NqNR13HfSHVu8X+lZcO4RKM/IYSopbdfn26l/bnvv6p3p9PB26woCaH7F0IVp22U
7Hlqdc/yuNOFTldrTRySYzm2TwbG2BJog0uW0wPR7yivRkwQkwA1GOzJ/F0X/o4v
lLcX8qPpTZG8AvG3LHwXRy5/bKs6tA+rw010gIqtbITerWjTKgrn2OzB0sv0RtdE
zMOLuamWtZRVRrcdAzdtfkZjkegOK55YvqIipLZ8PQgcC7+5H1cD/xHcKUmRtRsF
/tUwN2VVh57TQXZ198ys4WAyTH0sfz3AaT0/OB4+d+aaLFagEFVIXlwLYxqRjHV0
hbJeA/t4nC5UPuBGdtUrNGdKr0OMx48Dpbq1pp4I5rkTmgsFVYXP2aLjEW1CBPIE
+/7HJ+OIK0KkFtCqsS46DfSrLuwLEAKthaM7kWi0JdYu9Yw5RrKi8a3ALcpzMv4U
2P84PK5GeKoLE4eSgHTK527wKaZPOW7gvHjhb+djnYCjE2n0Y4T5Xm1eEF7VEnhM
5/Q/hJpnrRqg9T70tANx7ihzAAdVulA7SFnMznNqCvyAWF7QW9M8b9MLNjoogVnT
/C+FnoUQ50xjMjxT6EdAZBoWZNDi55gOOtXkGM2cYBVlE9JJeWJFq5Vj6I20/q5L
JBvCHTmeKLHl+QUy4HL7rKwsJMfQRLW6ihPEXCDXnpk=
`protect END_PROTECTED
