`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBjnM89v6BkmVRCm4p4ro88vKf61FEm8JO9WCk44bgsz8DLV5IYb22AevDzk2Xlv
8SordeSdHfJiSA/+T+KdHV9AysGBwESdhq/Nu1PXaYZvvm+vXAbLb6A+O6JXNg7z
xE/7fgzjihq+wi9PFOWFZLOfr7FlkyJM83qyqBgHr/1Lml5l2HZOtOe1BN9hfZLt
1o9HRxkJCN79gQDXRA7Kldq2EvszODNJFlWe0NA+5+IjXSTxPC6o/RY2RhBGdOB9
Kt4LOtQKGFoJvF/ORVRFEDlwBhkG964m69r5jWTrhIEx3kBAJ1juzFgmu5KMwoO9
+OHjXPuBPIwOPfK2D4NZHzjOB2HoAl/UfqhBgYx68SsQJRL0hdiGiTPIA0rU4qGx
nrvz0na0UrKy+OpSPSes2AE8f3sLCs2WSakvSUUBXYV/aHJOurbtGXrQyq0S2uvd
aKbP4voKtD5Oc9rf4q9CJ9MTndtZ/PKmWkf5SU115g6ZsymOIhNieX1NEFn7iBGj
95fFEblMDNECs1zAfCdAON129KB7dS0fuNW1x56PdyZnU52jx2rKRmGHhm08uR+d
8i+q+4uTZ51F6Bz/Kori041wwczhOU4wIqFrmSMYPjkBXksP5r9ETv4pvRMc45DT
8BxgVoh/DhjtXvhJwmNZ4fmK++Sh/rT5F/9ybIUfprIvVezHrgF+osBuPX/gkzkE
cST9TWpIeG3UQqyTARxF3w==
`protect END_PROTECTED
