`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QektjYzKNHyEXEi/DQy7P6GuvY25D8/TlE11UfsGKLe/KiZMbBdpGrKZdGsfMIbF
G8YF7lV1thD8alrp57OLKSX/GprEYrsCQlXeJsPHloqgEuNneP8or7kfoaNaeavz
UrbWJZ1iyps5xsiSAvHFD0EGaAeD3NhPqCSS8HiQv8NVTvIA01cjv9k7vwylQ92/
1IkZxh54nfSdtamnEh7HFSeZaTWanQEa1iptwMgqJT+saF7oPvxh0KzwcBVo0eVN
kt0QLr4z0YrSVeRuiDhuRy++9d6rjgwxm7I47IHrUVq/M0n14xZh3ZJl6ysO01fg
hb1xWymS/6Zbw34A8RobqQBxz5GZSH1ZPQylUTicy+d6dbtueFQVzJK10eTsj1ID
GzvRZiPB6OsnRu0hnzcfkPlqFhi3uAL6WDOsXnWADcfgAcBiSN5ZQ/sP2Txq+/Uq
LSXDAGTzW6qm/HXirbMXEchxz5hTRwKSc+pOvqR7HEh99bhr6ZgCQgUsx+WRMmIe
brwMRC59Db/GeDH5/ILKqTePke0Tsn6D2jacWQy6r1M6fFqI/Ey6mo+PcRHGrOg7
G7L3rjR9nv1Njo9RoZ55F/q5N+7Enp3NUnECtxDFZiGS1NeZDvTaQy1tZP+GIuO0
Y1NSMofOJw8BrYixkZTl84OhbZm5Uu80w/nLvxwBxh6hxWL0HeAaBPEgoxEXO43J
tAsDAdzhbxb9SwXCDdetYjxunD5DZperLuKB8cjSbbR/WDySFL1jv81irmMs4dfB
xyVIIpghcDNBEr3hu/AxbhUp/Jzi7Kg0TGUfh/orWoHD/1ZOt7ll6wYUnaOY014M
htpE3tNVz345riZheMw6/+f4R5NecVtIdkhvAWwhlf01X69hZK0CFqlLWVsqdZgN
0nu1uraYJiqMS5mCSdA1qBqBpdwArCboX3kPFfKyNS9RLa/J3mDtXSj8pS9NXcc+
px25zrYzICwXrIF6VmretXiwaxoMMCJjUMS9IfpFa45g1JemWTftKw68Ga8HAEwJ
oHQjjlS4J2S8RPH/UE5LEn2+FL6MnFWTfqeXRTH9YwdrcowMDOibOTexKetHfomb
dx1C7xlrREM2UocISo8+Un5a7xDg5MnuuC1Bx53uQgcxNRRAEelITmr9Mx4tPv7C
YzmGeV2O0i3SlZ8bcOHEJ1qtM+7jCKMOGvVdxuX8rfHKUdsTsNtzRNfBnfF5ggW5
cSVNx+7+VX37NNAAw+HIvqnsYADZ5Yd9WN1C1lZp5k6QCBxJowMW2MU3RphxaV4s
XOy2s6oMRqHMX+s524TonKcjLquxn2VVCynZic42H17MUw+J12z2gjTKRVDGXG5o
q1u504Fm6/rfUGABq39vANMdjwiQQwG7Yl45qpCgfRYBkRnXDsPF4S/2bUqtn9VV
WnVEOOvSJ3wokwJMPdeqZfIeXFTG4gzUEcjOGYcjwzvYaTlG3CyCFhFa8SvfTffq
tgX9nmE3MJ63LvQP1aKyYh7yJOYu1Tr6UcaxH02ZpLE09qjyYfxY4lFbZnpu2l+q
8SsVaHA2spKWCVn12dzK9vTZy7PP78rnjSUujSfwUkn3nC6RVQWPB8uzWPqYngLf
NzvKS+Z4agBh+Fb4bflg1Qqx2qMwAAPDJk3JBOAB5LKM4J19atZJP3Kk7isOfqsB
iEyPkocJVGMd4ieE80843vdnc5WsOACrl7SvBeOIfBfdh2xde1rDcQP/PmUcEljr
kM7je0x+SHSj0dIUzQ3EF+yuQ7mR/+dr9dfYklxrwVkgHZ5wAPWH/EEkg+QDVk7t
mK9q9oCEot9mB3iCxcSvV29Kbg0iEKONX/GqndKYlD7Q1zZlM+kF77Q06nwquTiT
i9tK1D7hau/InTKxATq+DHOvLkwI6R2gm4+lSLp5qfsuICmfSplo5hB3ufUk+ypl
SWqEm9A9slcaGiDReJjodGM74BL98ZPse94xyE5h13NrM0IY1lx3/HEuux0D8KRL
9XuruR4XpmJCF5Auk81znQy5h1EY3eX7bNt55nICJJshYXF9DaUg4KEXetE9gR1D
1IpAUXVQ6pHGkKz8K0wYwObVka6T1HJHVIaqxTj0B+ijY+Rzm+WdG5U2mMhP2KN6
y0uKRJu9SCg6EqqS9QCE+ri9RBoW3uA8P25Jv+4uX9Ked6HxzXoI/sz+glJZVBt1
UueDF474nf4pyqsuIvt6+I/sagG0UBfDP16WFrG6R59c11OYLyWlnJWAi0zbiceu
TD6ESw211o6nCOCVYTcUawBRnLA2iRuvF5PkcBLBXf3cEoFQoVIoeiUwiOtgX4jd
tPEt2Hh62k/uklaZ5K6+OijfEhBwAB4wUJYdWyd/5xW0jqtkxFEzquyTERUlBIRH
fJnFVfK5WUSCW4R/SuvOkX6u+yFe264Bu7UgAz18TNsZyPHt+gKyCv7+UHKhu1oS
Do5xqq7aDpbc+biVrpy1oidk3QJSZqIP4NwLmit5oLVAJl3D+hATPDZj89DoCFE9
TPgW88gLhyERAVWZqeFxqDzwuoEAlQ5uZON7UGeSMyX+FFh2synBDzmVSKRSvNPp
z5vsFDEgSpczKloKl8cGKNmHglx5h0+CT6G7HtJPNc0iNfEQ6HUbRKRdNHlm1Il+
ZBFMvNbQ6+FkuAh2xmYuL9lQ/uai1YMy6hnxxT7XU0yCatRXrSCWTTluMp0O6lq5
8lY+INmqhgMro+8kEB/j1xBFTamQs5JppAa3oIluNYkBIKrSjL0wgIcayVvF4Gtd
6RUSxVHhEsu0y5gpFrZ+euwj4A9hpQ+9jvpj4pXjAnIRz6Cc1Zvn1pNUtYWI0o4g
py1iDnXA5GOYanGzlgWF4CtjuRT/rHQ8MDz5zqaGwL0QapuvdqSclvdjCrpRbC/R
LL/9h7Uv/PJj1wdu28RRu/UXXDHOSx1KjeIHkHQZHX9+4bx1mR5D0pfS4hvlYcj3
oylRfj2AYh/vV/JPUuGBc3yYMkDkI0FV6V4rRcJzTH7Bhl/sfeBBhIrFzdgy3QcE
wS99lhn5LIi3SQMuOEcqiC/x2uJWpZ7B+dL3sp75N01CDyljeU0Xa7IWX0x27NMj
D/1FunWiUUI4tYKbCym8z8YCZpAS52VhOhtkMtvUghWOSVEP4ROedULdh9rdJ67K
JWF/T8loScp2ysTrGYiIQZern3e0mxdiiY2IhIneG+O/zqqQyfP9gQhYp6+SF/cb
KZ/2lCwc10fElMsAeKMtzLneK6FdT/MmwHOyff39ggrRuV58H2SzZ+llrXbNf847
EHZayyu86/TjbeO0TtS7Z2WDkFAsA4kTmBevZFraDutcMfAPyS80J3nuKXNBzdwx
FfZ0KMigXBWP5vJRHpqvZCXG4+61CZAgEbptyprKYQfWc3Lqou00Hhes4lbwH/+f
ub1G0D9UzEmrvJmByXCPYpG765VL9QMtwWHaTqgWEq45pymIxb0+BPWNEQ3adXUR
4iggwjViRXWmKebHHB4EUcvJqnct0Fs2rmU5tNHg8ZTT523a95MZxF0ZkccPtIix
qPn59JEpViIn02uZRNCAkT96WqqugH4Xg/l6DsFswZAiQScMAXQHmD1k6mypR4Jd
BLhhMZrkB7NJ6tHB4RAerRD1wPbyC+VN/z34wYDj84c+hFtCXRiohbMfVYB16OBb
zXpLePal6DTV7Bc1bDG26FjT+uYDN3rPn+EhmGsa8BuviwWM0Lg/JhvCdpl6suaq
HmdlD4K9xe7THEqRRFPRs8344qUWarv+BOo2xTWNg0KoVfHLI5duogvSccCMIQhj
tvOmsBnC1gZ+n5Gwg8dacTJIxWROhfhgDzVTNGFhOV5WvDYCYdkLTOC1cHIcCoO8
QtlowNufAV2pSWQRBROf4XmRHCZJF4mRYka7T38wvsyy5OGCzUYaaCO0U7tb7tP7
TZ2ryiKfGkBDItdG6Az0G0nqLxwXeN5o1bjwTzFiwH5+6Y3XEe4kaQ7pzYwQWipO
WA68o9ZZwKx8H1Fcj7ijPKFuilW65CMdd6Z4V5Pr7lFlwfhZl5/ausNAY5Mor0oD
AcIWyviwKBO/zACQ4cY3YQy2opyAz0WMb46gZkqSmBb/NPWqz/yamgN47KzBmft7
qqqSGLUv9w2I1L3oRivUdDvJ1zZ2QoaohopcgaOb8lGgrHny5ZDbETCwSgPb7FRU
rLXga5PddRTlpMaJfrmR1PEA6T5aNBcXKe3TjWuHsr1g99hjY0PDOrE6qgUWPfbL
FUEDxorHxYCfUuO5xVcOLWNAtSYww3zwGUbTxq8jfPVWXQZIRwfkpOyJXHtLTmRM
bV2jPDzirpUx3drRs95D9/stAZVlo4Ce3YAVNRZxQxTcI3WFEuMTI2R11Lldqj6W
JNrwUL8x+ShXWQCqjJZ3W9uTSsza817Er7QPLH26lBC094Mone9CqiV9exPIdCHl
a/HQDspxQrT6wLMhdc8nEk09+UwX6KusuXKLk67ktc9p31NA6yFk0nD78F+QUY8K
wZhWTFHmPgOOMid+Sir+UzPMTFipAePg650vonoJJhNOKHjpmJnmslU7uTFdywda
uBxoq0BjwWjqlzOjtUqRJyW9TbnHyY1ziI8sxXvOjZHVIgJXKSghmgPyp8vlSNSo
pW4bkfkY4D44j72xR1V58rrcS6wmnvvYsTt9cE57vm6AzXKYMUfcfWbm3kTmIqXS
IupPqtF9mT6NUx7pWQfCD/tVNGED9/iU732+ll89yYocwylxQT2ME5BrikfnttVU
Pl4jylYwVbac1V1B+z4L0KqcIDqfgBtHLuZI6nBuTJ/1OGvPw4JxYvYyP3XipDaG
VBR8DET5WMZPRmJJIlPLj+vXXUcjiBe4Ry+pyIfhFwX3SGa+EXxNjTWavsqMzrFX
XGnRL3f88pU01h8bUP9+9GVFdFcECNhpQcqUMtsbvaEBB4HXR4x2IfZZsniE0LjL
ffv8hzZlOzFSgEbL3N/E63KfwTJAYL7AQT/rY3qsXmuxKMWJmOvLFpz0HIolRKUt
yl8dGYHvU2HBVLO8Ykub2jP+Z3jc33Vl/Up7TeE6AhcdOTGI5PKH2UjBBCbtorXq
FTqSHLenB3iyWAbvro9368AX8skJhbLYrFRmAF5cpnDRREiYiAm1Xga0f4SgmuFP
mbpagXwbW+g/kbKy2QgeZWeswwvjhwd7lVIuHaDU+Rbr1kTO+BOJ/orJ7a4YI8iN
UZOMoLucEFoSsgbXZT9LrlSCf7mDPYqhzrJpRFRjkG++n2+gr3zBsOdKKRghneKT
Lw4Y7HlCS/9sYJ4ABUSU4VgdqSydVw5sOTuVHLCpb86tFJBgcc/1ZYZWFpbQpleA
JjZJ94GqJ4MFK/Z53eVJKiyTh7iO2gQ/QpY3CAwhd0FQJ+kC+aSDUAp8jXOPGt4n
DO+LBbTV3ltGIyh3CTuHytfx9cCWIiWGkCBSomQ2vb23MCLDst4g3CgBx0Zm8yjB
KU6odS1+kwy0PkyGaFBGaUOs1C0I/zNbFK4Vx773HI+42j+e/XVQUqF9uzhoCBlQ
JQRyCDjR8MFh9VlnKvUuuea3p4S1JMUyqymQsinA4bvKYA9IDcZElZTRnt+C63OT
7J+6bePfclYtoLGNNzn53/ZFF2D+Z8Sp/LrHeqSmNGOQr2ier9pXjXh5OGibpjre
Y7L1jf1n6wGt/qolhYLEkluyLCbboF1JBz5mEgaF+vIfounmv+B1jEr1p/xn7a2V
MW7CD3eRyOF/A3YFIRCgKiZBfwBzM2G/RQTqcSqcRDjhDZ+SQ7hdn4vIAP7juMF3
`protect END_PROTECTED
