`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWl27MmXY1bLAyiNjy+6BLFBKUeWA9V7VGmS6Jm8SSOBEBycZP8Lkll6ZyinRUSE
q02BRhUZ5CSviMdNnpNiK+1q5OV6YXv1oSfcrfPMo583qnO/rW8pYoMeYTPrJkzC
522prlTDk65xUUNvVOsf8LAuk2lgMzFJGy/FqRmxyLcFUUoCOH879JaR5neMA0oz
8eySwH6OZcoTrzAGRhbomv0RJnbKppp40T6y/TbmFqKTEfoDqZmBgkwNltrXQEZo
D5WLteWfxEIPKNkHTAScktbwO8xN2VqFR43qRUMuS+CGGsWkTywDqVD9FQTa3YxS
0k6mzO1vnrlmR5zAf0QEC94xOKOuoBuLQwpd4PfjgzlJbJCQxFm+mujDXefpOtx8
INbwPsFtZ6druH7IHs7jnkhlyEbf8TMavrSf2nvJ2wQ=
`protect END_PROTECTED
