`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAy8hJdOLyNUBTHRDdtomnWoH1sQ1F7XU6C1mhQ/Jd7SytvSXPT3E10A4W8dVk0i
qGXtIv3pP5OrXaOLNm2yQWSDgnmcRGn4WI7dcWefYyIRVWlaK8KZ1hGzxLVDB+JP
qy4bNKWecY47z9hZXMCba0omcC92qBPbrYoPEr/pq15bsGFG4knKL+fc5IcJhBju
K75gv4IrRvbtxn3rRldcldC2BLivRc+HRGGzO8N1NqqmlsgqYbn5NP2NHmCONkdn
qgHpgCbG/9d8c7+Dt2N3v8f4KY1yucVT9bYysw/PcIjVzsPoNFq8le0B/wpQALRr
xLss7zaNB/OWVrXw7GiEBPIKZohWYBKq699tyX0GAIDqIXu16j7KEyoY9a3vKHxf
EMGwtFSwHSdi2zfPxPGmzQ5j9WASwLy5YTJxJCi/jOPV40IG4/S9j5X/e1N4HfhB
ceJ9N0wr/vZ3vktMDi+YTnFV8dn1TD1uqMCn+rIlQFA=
`protect END_PROTECTED
