`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLqLJjaZ9RdM+hRTnoCkiybUOlKXkNvr/0oR0eiyImCyvPV+83wDtsIi/eybE25+
LDq8y368sBqo+L7oK9hHn4OdAB4eoVJyXYF5p9panAY80DrzcNiPcHjp5Me8t5uV
RgG9Q4uwV2dB3nEA0A9EvD7mlwpnU9mhIUV8DDnwinfqTdEEeJaxsPZZZkPlexCW
GcMK4JFm6dtHsDDjfrzRuFLMiSdp5rlAgbMdvXymdbskq2bWrT8P6fksIuRicDH8
OM9AuPL72JXWLP58xxUJP0DfePLnSXQzMyvIHU+GbEWaGBjSAy9XBDAV8IBx3HrF
+s+pq1KGxTkCuKh/wnmqNUwtQyWO6w+eFqhWpVVArBQK8pbQwMwsyIL6lE0mozkJ
vGLEDEb/ThfH5dJE3YTsJ+dozVfetrJEhl0k4llCOiQVpLqhdfhMeV+hUaRsVE1k
8ACrpwHBWRtAi9rfMJWuwAspcgdnDj/bBUxZfJR6VQE=
`protect END_PROTECTED
