`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TftqqfCQeoF4XiB6O/7bSTZrNIogoKCRYFcLT17GuAXzJsoznNV7cNQsBuIseEzB
3ISjAtFV56Lylbu3bVZ037+6x8JWOeyNwl87EDeDPJ2GlMtw7rB/sLAWEsO1sIbE
HxRONTFdjF6WdWd+QVU/1soREak2bG759DRb8vU2gRngiwus9MjEirXkdtihmOyy
HhtRGMvjDTDX0GnrJiVq8D53xIBPGfPKgydanY+Vt/seNl5lbCQ3/PxKdBBoEgtg
GQbvO0LKm355U7anAo0T7g7o24JSQv1esupNq25zjGcbELJICIa99rfsjzcJ4er7
B1ySA7d3H2+fkcM5g94VxlHU0k/M0J/QZadxHr7SUhCVF+n7JWFV+tCkeWazC9Rm
rI/QcNktg5asaqVZjzzR2Sh+mekXrMREScUCqKaAimW5zGTcn6ARuH2dOraFMcao
hOccQ456CvRzORSNukKXHVY7v3CgS5G5rpxZlLjQZXqLjyk/YhANcRqgDzwo56GX
2ZArCDcqU8fy+Gc82ZG4ilPPl9UjRaA61SZZywU4GHyFraAJazSm5UJGHiNum5M1
VhVNe6lqP6YPA6tSn6IklSTquVrmA/7JjfkRe8VqtLLUrpKC1iae3ahYyS4WqqWC
cpuCnZEQMxFVLd379OGQQ+lS565LIS1sArx/jy3qpWNH6026aa3jevgJQWSlYyu/
oa0zpiSM/rKmz6Wh0b3H+8vZUq2PgnbpQldVy081fct5GhtnvGj0OqqsUOUUqzaG
8DLOj0Omyp31mec2SVH6u5FEKOfRq/HxFFqrxRIaf80EQ7Z7/rgWL55Ws0qT7Nx8
fK/4xOWB3bBrCE/bSCUo3Q==
`protect END_PROTECTED
