`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXqf3uB0SHeBbelcXTvfOO4ZPc1zUeJEDJQMJWg08SWGN4GB1sDLR12VM4mgqcYB
JHp5jliBKwvB6l3YBI6blznsjgSJwayYrx97RV2LQv/XlLH1TSqNTRCqHDvtI1Qp
E44V52o91SHEUWUb7RoHddvZacY0Y7hSLAsHXSZ1nHksKqJ+emdrvF/yzdUuaT1N
7dVRBBatoWvifZB93N5eTvK3zbkXcLSfnaRJ8yPjb3vz8LCQQEyIq7pCzb71NGZz
Cq4CsBOPP7GBSubszktoBUybuIZAybqO0FRkAWxBtikzR0LHLN0budx1oYu6W1dD
`protect END_PROTECTED
