`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9CEhplqI5FiYTOclJXjTq8LN4nxdElGCNqDd3JokacG4AbYMkrxXoFelHsX0BDGJ
CX0qBmpSSTv2abPnxg81Um54mffwcMI6M7AU9PKgS8fWwwrob+Vn+xJ7rUq5Mg7A
KqMrizht4eBdcUFaRDs5kV06J6eyVpo76MDymcTuE3HOow/qR9s8baQZOYA+qO6Q
/C5tuOWTuD9G4RL1hKhkPxR/J0DzCNViN/yd9LksmS736smQViw/k0c8pRf2GYZk
XHiDoz/v6UJqhYZiUecpJQdn9MyMg3pkjoZ15ey/5F3mnXEIJIuq5Ksl30SEg04u
5RrvsJy8K7jVHxFTlaEybLQ1gsRheLUCzHXHS0S9xGqDh/ELlI28tSEaE/vkUdIX
IouXNEbrVzVYtRu1mWdLHRyZxO0EBlLBCn7gDD/V7pRMekO+I49Lfsc8cSFTx2Be
LzL2c1CTL3N1O3OxBRv5u4RXe+YulH8phXbVQnUM43vbiqI/1vAcXEkNGNwNcyEK
eQ6ycfUJRnhBqAH8UZbBCymvMlpzZJguwCJfyNm8y8u7wRNS0SPvAmX3L6eIzBj1
wKwqxQ88Qpvse36q/Kwr51pl8nyVXJcYpAVGw+vJcBImP1+IQd5mn76U6yk9zcRN
dD7Xsy/Qq8tVTkyo7IcDSjA9w2qXWoOAn3E2X8sWkFnuo5EcxdSj3oBKlfpZovYJ
SacGiknQAVZaiUlZ84QbURxdbje5QB+5kuho631yWQRtiBnbp610Yev1ziRwA1eU
J/8Ko9g57lkM6V3sMv0LL9NhgKGA/c5vnZ8VHvuu2Y1y81uCFE3MJR2o58JNyco5
Cv9CLKl3EFFlAVkrd7Q7VaffKKgFGB+vGXTslKAkHfyqv/PWMFcA9YRoPnB5aigW
`protect END_PROTECTED
