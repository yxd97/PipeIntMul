`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8EfllcLwy1EnlYsD9bfU5uvmcmn5XpBun+xHAvWQ9YpqkTBoPvGks7tebO7/fXQx
fk9qeI8Hndu0mBrXFnpoAOdJRLiX4mRPrhE1ATmEdttR446Fmhw6yZvopBCTOakD
+uNSEKGk/MQlsl9GA7iPPHWL4mUjPWefteoIsxxjfL0kl3W+viDjPntQ2auHz0zF
NP5plYMwO4yhUO6KFzVUuPt0Lf5UFjmqT3R85a0LOiQqkP2SL6QhVPTsx49qIq+i
P/kelz0nW93VyfNpyutTHUrVat/oepGYrvRhp0RFyGkJzm9x/PJn9SrFhYLbDZkg
t91S7pxuxWXhPoAPVPxLYFEkSlYQRYzzwoKhwxuUBjV2WDQ0Fpgk6jCdmcnueWnX
UfRqSVHlMRHI1Q9VcNR+iyreu9ynDxm+yYb5XMQ0fY9ZWRxuqumAVI6hAnIgo3oC
+7xSWu6R3EebglHjb3BGUgEPHZ6B1swBj3VlOe787Oo1Oyxzwd9yOg8sAevTkkkX
wFtjaHG1khpp9vNzHaC2tLx7Y7wS1s4pQdYhZBbFm94MMRiAFJd+86bVOwBZaMB7
BgJQ9Eij7MxsZHbbbSWfdOGscXvpGOElw+lgY07/lldqG+FOfzOFUz2ArEDs6OS0
kwgDX54gqcSYzPeMIk2wBUfYXQpD9jy/vfv3NDdCHTEsKZuj78YTDDoCQE3fsCJ/
0UL99fRjIZaiM+mcHsNcKl/xQj52PRih6X4r3gwJ7DpQr4yMZz7vITcYL2bLZ4eH
nAvWVi34Mt4mdxq1/o0cqxuHajCywFBCyWeQ8Z2BKOfbFCeHrCdu9Xo1gx80z+OC
4TJlqihgngVIQY6DZ+HhobGpjWM1uhjPCm489K1ep38XFNH75IQPT/ED85PL6Cem
4XCqFH5YCFib11QtZzBvhKNHrJbG2WZ4vWknxj1QH03lND59EqJLMEDKS2aTDYq9
6Of91HiQhzKmMqLwKxvs6MuhTNAxgCYYzAOt7jMuu7cdyNdDFPiO6RmBfQ/8iVFi
aFtxX5KrELUWDu90750cdDSk/Cf4xC7b49KdLSswTCSLUZVCy189J7SCzk2++bi/
a/F/ezi+tQPLW1s0BOETClXkixQb/ZspL8uZ6St3YFkVC77ECCVNoWqi4vXdcnBy
mzP8e5JB3oBgdvMqjXiQhLZGEK3T1nQ1DtZxZZB6wBo7YDY7dCEKsckzisVFMFGH
N0gmE9NJTt+pPLI7Q+XjMmQeOo0TIDOtdR8t1YUZclBvWLvgw/hzQ4n63o/MhNb6
bMXApvrKtenvO6ZW7KKvZB+lUoIQvjlGkxCPj4WzuOtGWaMmNCQE9h/WSL3jkBlj
OM/dg1KNRJepzx+bKhipy/ta1dy/62rSIlB4puTDTLr9GOxA92v9sH452ntyAe6s
MMi+bfSWKemOmsn+QFH71LoJwYZ4SvZR1ZEhrYPC3I5dtJ70EvuXJj1fP56/MqDD
XEaf45331YvF3i8tqypVBC1KSFfMQvwRyz04lDg/7Fn39HGvurF3xjr1WVjxVyvP
K4X/8/7juVymWPXyfY9zHBXioUiNgGD2tURoXIOmam3udzqnx+k390JnFqfbzqIT
yIsjarKsiAIVzQBTK1W4szrVBtChsAhgg1TTu4+dh3kazVmyHYNbyAv8g+htEMrw
CKKk0qcIHLoUTPf6NHgyLCVbq+9jzkhsP6KQz4qQ9Qv5QFAUXek63FmWd6hX1J1F
tsftBWuOv5y1nze+P9JufOZXfropJ+8MnQwPXn+PIyuqaTTPhD7acVOMq4zPmEs2
110oxSLYSp3f7dDi7OMs/eU15PTeCzRYEtKZKI16aTbMYLFmFQ8w554qQhpemMPL
`protect END_PROTECTED
