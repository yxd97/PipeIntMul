`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ySKK7IdoA/58OVIbpr6YzYavHVZXVy1d4ZjgpIJOWCKv++fvnx1Y05NGZbTdLBqX
mX95o3SwERLA8jSGirftLJTQjD/j9xtfBrw/hw0QYNFekIKYHreM7AwgojOtCvr4
/0/jv9XJ+v81/zwUF6cKR/wzZvDept3pE788+OLwi7oAdDCv8ZYDpNjrreM9Q66O
QjGKjsFjWSibLukHwTlO2EhSpSrfQk90eWjdmnj3khgMfmpLlWlopkZzqx/ZckNN
DIPhNViVU4y4Ptf9/dudtGdTf7zLM6uRtxk/hORgQ48nDhxzr/aanJB5pnEf6Y6o
yaC4NqHP92mdc39S1mYYFtlo31QM7SaXSSjPH35HFMeUYyINAlGBUKWPeF5zmllI
Vrz316IVWWLL62Ynwg7PdL4vyfOh5bBCilpKVRZhx1qvnlGiXwZRTbt9EgtNAak7
QOyGeNvIqM7IvOQltnuV/J93GaKjOyExcpR1hx0feclX/Hr8lEugQVlzDuMC9oxx
osV9mYGSWpjXpe4xL06subXhMWwEJFiYeLIq4vnKP7fgOy+TdJKlemf3JzzjcyAc
2o5cgLtm12q+IUXrHUupt5W8r/NNLTIYlAobPciUasqr44XXlUtosxUBDZ0o73Jr
MrtrZOtwDFtu03F9TDOSZNA7tjq12IlMhu2Eb7Oy0oZ3oNCF9/hnI9jxWkSv0iag
KVVTpJz5LYLDsbu3Gtq0O7lXeLNl1RoK0YAuVtPAVCs6GqrCNbjuWS3oZb+A7jSD
nrvFi1EkmOiYRCQkNLywpwEvfL5qjwVMh5QN8OPlW63BrJ/gOb1b7kvYjQgdV8lT
rYH/0mArVgISRt8+SwRWhVAN7E2kgqx4zqyUyXENJubeBvovEGaZhbDBIs9FL8vg
hqz3WDLqBII3puK4fWPNbSS/vLfHH5pS2dDawSUFezmaA44xltXFGLYBNF09iXe6
GPxCpr3/fguLrX9YlrZP+YSCgJkJShviBToBUjEidEI1tAzLYri3RI27kt8DRxsz
lB8hrVmGyhKI3Ag5SEH8RYf3OQV/8vhroZR3nMyjxXUKJ2FHhnu823FGOACZnifB
uW+/j4nOjlNGJRX2BduYMIR+fzEAoc6bWZiqhRFNDlBXFWIJO7pGGAIGC/T+ld5d
JE1w0aYifyooxqCFxyj/1DyyiEywR9Aw0xEkbq4dtWEBHAzMAa6GIV0ksVQWaEiP
Aw3ilFEEgen3JXktZz045UBPgFdCQltRf3k+RXyP4/6o65TjEQvnkKLRLuQLqoGy
`protect END_PROTECTED
