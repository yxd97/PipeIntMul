`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lagML8YXVOqxDr/1cBYzsFhdz2+ehjjEul2YUwGOYmsD7YJwXSusrQdOnECMuewX
efuNVmZ6b3IBvgSPOqI0ETbF4umVjUR06Ez6mzHS3CfCW48gsR92BKBkAR77z4Pn
EBANwjs83akPigirkATDBrq5TFFZtV/WXyQRusnwsfLC7VAuN/LQwHTH4tF3TJAl
kZ+1blD/T4YbWEYgegc/54jiPYiDMCPtYYxezRO/7Hodh6mkzLFIWub1V/1kT8ep
pMbtgiNCMiFoWHxcIQFOvh/QrR2axfHLmtXijk5i199Oow/zVEEpPujWZfAAH4bU
4vqnhPDTAi2afnMIOVByYbtKBK1S15AHijk0UIcmWNfJrxKfN0CdsEESO1AY529p
CXjzG2tX2h6yWZtILU0x1Q4daVHWjOxyIHIb2MM7SKQoDeM72FMIDz9m0+W6VhVD
VcfeE1LymXgIu3x6eD6Y+ULyEZ2hp3UN+I0MtGZvTABga15AMFb6Sq5aT9GBt6Q7
qo0nReQ7AHzTnuCKWV3V5GRC3ztMG8uud7dO4KrIPGWLal7wEnIsboZuTc5mOuEI
C0uqNKlx2ccgGBmIFNUb9uSBKD5zYqaEze9dZ/K5sxeiRaM8QRQtWirfY/zQ5Cze
IwhvkPw/y+mda1IhcA50DaheeVnoViYBren9gVa5WAfrWypTka3LRcKE6/nfSu2q
/p6pC93dQ2WOPWUTpiGH2A==
`protect END_PROTECTED
