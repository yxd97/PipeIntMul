`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chS4o1NpF+QhxviR+43A0hPijaieaUj8uxpkTBY7E6JNBYbqMiaqKxLlbxNluVcK
tpA0ozUoOcHYHBLjIRBSXfQNo5iAD5/sVcfsgp+7fPJ6e5as2iyGAPEQJ1E4Gctq
o34Vf6MjgYwUAbzigwqBF04UCkSLcbm5CNXJxA7E+hfc+niBY+wFifmpiIEoyHFN
+cWTV74QPa29CKia9Eefv0PI1n1rsXdMDp4fk2uZAEoJbIejtc8XLs7znonr+tni
KdCJ+D+xEsutnZ+mhKlvrNLRMFkdsLZhwzAUMfCNSZimlqeGWzuyRlh0VmzE/H7e
vqa72E3xV59mk17ciEorWlakBcplFne+C4m6Lm4p4oCPwKZnGLNeout7phMepRDF
OgjK3ScFMN/K/MjV79WNbGA5y74JN8E0s2D30Jw372t6Hi1l5JahURhDeJo1jNj3
JxaxTk/ECWlcKwyoUk8bb9pupyBoKE27zfzW9U1VOeBKelkLA1gmzcNI7uSXeQ39
w7O1hqR/GjXwBPK54m3RAkZbgak6OmXieVWuW+B3KorYWsmQ1ZxpZg4cTl9WCCxx
wIX5IRkG21w8j40ADlMfUS3iAopMhVsUdoNFuZg7vi5+X3+/bPhLt+oX5p8Xa/C7
LUuNHZ1lS0N8lLdonOj2HZmJBwvHzFOu3YdtrSPMtB5dUCLcEWcWcEQEBBv0x4PI
zuLN36U/KlEtdsau6EQwbXiBbOC2N2i28BCFQjUyC5+AQ6jQ50zPti0b0oCi6lw5
LT7u0HU30LeMQuu2dZM8SA==
`protect END_PROTECTED
