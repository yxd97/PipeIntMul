`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4J4FQg8W4BeZwfQjRIOrBvIrlKYJ5hmwAUsrIh6O95FnyTXEgxF/wcJ6Cf15HzlS
SHkRzXKSQBFKcJeDeIaEr87+BjO637byf71z0g1TBHWyZWDLAdp80H97HcEli9DL
h83lKo8IzFCIb4lNaBNyySTT0c6JNU/gFfKtGiZoCG+/6cr9zJVzv4YqZkAO8wnS
Cy5jJ7DmqaeSmfYHrr+7TPJZQnDEDHp9yhQEZjhlRKJ4u2lOPEoUEbqvEZ33T3+T
YFQMC7d9ADXpIn7St0ci4Yq2BoPMX8tbIc7gXQaQneW2tjXZjtcIEtnCh+mm+kaV
iOoQ1QGo2TfyNUd1hI+zVC7zlu2jsD1edIveURVBUKqVCpaIk/4MwuGOKuWQiBbs
E/r5p6A+LQuwkoHYIN1jvVcOgO4PVjOP1gNCotm+Bz40/GqH/v40UK3rIzjvdey3
n7t1PA4SWKyXr/osN7IH0msOhvgUN6tYdpOjB0HMAfo=
`protect END_PROTECTED
