`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2J6K+WuPOTsmT17U6z7d8QB5lfQxmq1RETHdJ5JQmOnIJPamlCvvLyYp7UkMJCq
AjeFqf7UWQZAyIWZcgHVtNT6Hvq+q9o+QS1ocLCX4+mdG92iisqKZN4LDcBpeLI+
vMfZNJ1D3vs58TGq/TD3pV5MgG8JhmCaWRhZN2Z7fMcaDm2JNJK2PRA3JLRStU9R
SiItGYkL14ohzO0RZ+DZSVPx9Vp5Q5J0AipLZaKH++/aHCUiFXfuO2peLyh16NHR
9qONYsO0LPdntxF/18t91aBDLe0laPaydK6gEvITEW0ssMiFdZ+cwfCcRSD6ixNB
w0TMXQ6bvFad8jcYIfbPio2zqhsUV1Ia3uUbpxO6GdlYs0yHdHP+wLJS8WIKUvms
`protect END_PROTECTED
