`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NFCBztsubIMBqkmsT4ha7SmFnJjQZl4Z++JY+44Q2iD6obXEr1bpJCooy3InMCN9
YXPPDmxuxUDciUMZdbQ011COvLBAHhwYv6obrF487pk4oHoAzRbVCg8IIFcqbLig
ojR3Be2fdoFdq7/ZpnBlZXjRGudqXRE3yBkvAabgo98CsFd2P9f9pDa2IVxtbcpw
QNNGgsSx4yZSc4Me05Im0bu0EFNPj5FETHjcDMK7BCRTxRC/wDrFcExda9WOfaj7
5vH5irKtfcVOZMrXp2Co1f/I4HZdpXUUQ14hgHFTFM2xuynp3vxMKP00ASyzf6Lt
09I+p+JXLGEgHKn6vg3CCOzlDHYHrhls1Yd3dhTf95Fgo4FqDlsmfzVUZktdzdjf
MHiALP0fjK+okQ07llxdlkNiNfbwLJnP++K+PR8qEHpf1uG0TbIZq5b0Ck8+ZsXT
WYWFt3YpdMVMmKr70ZGNxPN4wP2/OJ3ETUiQnXOnzi7sPtSSzuOo4JJYtuFzx3e0
`protect END_PROTECTED
