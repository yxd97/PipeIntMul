`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
USWYF9HMb/KETJuAhzCIaxfpQM9UtESvyILpC4rkJQFhghEPvPFEZcIoGFLPJVkg
jipNXXhIDrU0TBRqsCperkaC55danJnZmwNpjbVLTaUpRkvM7eKTkTBkDiJYyyfZ
2x05leuoqeKuQtszdy4p+o6UM+wl/j5Ar5zdWFhoK0xiI7hzFJ3Yh4nLEJC2+TQT
OGjVMAA+1IwO0ArXfVHDyGpKjF0RvN+kyeR6o8GeGU9u2HuoJXFWlkzFrSwTD3kr
N3W6pvnNBkeGg1qJdi/ZJJ8J9SpKsCDYw0nEkDC1IXx3k6hpOhp4u3KVaAbzTo0h
rj+WkZUi1oGFJLaJhNRaLAsdnRpJizP+pG4A/uLzDclmwJJQ+L6+XrkYYqDhvTq/
foSjOAAzsdaqGrT/B2r7SjWCaaAPIVHaaRJe0zGsVrj4OF0T/mkNzIaLmXLBdmfo
Zc05Vgc3TukVHlIFkC1qu1QJ6me+MX2IOgjbIbQei2a0tD6RnBfdMf2CGX+gLEQC
TJ7p+WO5uOaQ1Vw5UOqS3QgW2HxQy3/h1zMW56N/nq4PY3hamnwkg6dPnbTg369L
UTEMsuMVzWFtTg+juXPv34H8G1VJUrlSrE16xsbjfHhGOj7DLeCyMruX5qKE6/zx
EtNC6M+hiHoI99mDC7dJvhGwDC8NU3kzE8+QNVazmI2eA7iMyYYwQnRGpmwD5edp
s7i4S3IaqdAg0+GHIB9+uuls79G56ztjMV27r7xxT/9/OhC0dZlS2bKo/6mXZd9j
4CjKlAPhJOoVTn3xGfcgrNJEGd+RklMK4a1bw/cFux9WNltuKP+GCNe4lw2duqgo
WCNckxTw7d3YCDpC62BYNQ==
`protect END_PROTECTED
