`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gZopndEoF47zW7+0C4Nq36oQYq4xLY2WpmNNIZErgMU2IQQyRfp6+56YpSV+V+TB
9O6PxyqRwon5uN44aa/Nla7Kw9r/wEHst/tZITS7k90diXU5B9Q0YtbikLwzyKUL
INvfXHTs8SIlK2uXQ/kAY3HMMrpP6uxbIBgXP0R6uqr/7YrNL4TDqX9b5+2g7FZ5
z6VeN6Xdizp0R8RHQsJd4WQpUzxuhhf1Uty+wJeUuQTl8Qc0azO3iJjFGw5W94KZ
5Teu1q13Mnsc2lJhXcNwXqFmeg4Uo2yrGs0j4o5qwqM7nxie/+1TvHN0CO9P+e0k
dqgEp/eTQybnXPphSU+vj0225OTpPzu7lMWVO71ttANc/3q1141wO+W9fj5K8PjV
2P5/VV/4/RgrDmXQ3Q8d8tlqpMgvV+nXwjKqKeGuCuQQzn+iEhY80g5SttlGH9vY
ZrP2xaHd45vsVFGIHnn+qyYdhL3rib8d4nvyQG5JypnRPOQX8MuWocnSSOQbPLwY
5hAH8k0/Ww4bt3gtmHS8Bwk1O0jsG6pJzeoBr1uVk+yzwzyL+M6eJjdBrdiuB2+n
`protect END_PROTECTED
