`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAzHk011kKhx8x6BflbOiDdTbsQa+kQvxnr/e9+hM/Se8kOhsjDka8hZw+qzC9ez
m0lp6e/42ojF2KDawVOQE5AwEAIfCKjmVCcJdl/XGqOA1u+9bPnkZTbWRG/LswLd
G7rZ7tg5pSf2AS09yoISd/zTXIboFuoYbIMPzhPRFAEFi4/SJYtULR5GJDqw0erY
ofGP1gbSVshEjV9RJ7tPVoGuDYFqrP2yz+XFwEa0EuAV1xTZ0yjo2Iw6jOQE06rW
2rX7lmk98nFy7cNou6edD0cU/OF0wgY7j8Pxa5FUuf3bexDJmv4RucT2EcRd1ZTn
ZQO30CukIOHsmMDd4+jK5qaNMuwnhCuFL8/kBuG44RByrBjdoLJ6IZNNjoVAE+uS
J5LmGrvh7tq7qLFWuu99/qILuOSnym6maBrNOnUwGfU=
`protect END_PROTECTED
