`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxsfBp7XRgMOlrRwaSHXbxCJ+8g3VGpCH9bqRRvTu9bcP7kmh741PJHs8vCPP91o
JsAFEaghURnmK4YX2IKVkMczo+/UljUfS8fO41b5CPhdyxt3lnaHHs2Uj6OLpiUo
2R+V1bTpGTDDSA3lOzhNnzaDCvzY6S5Wby2u/Mg8W4gi/4LwD5sOf7bqqymZDZ6P
HCuVHKXWDqgJ6iuvKsrfkigrmwgn2UAFPIz7P3qVcpBzm6w8vTA/7rdyCfNrzlnn
HuxqX6F/hVenTFVki0SvQcg8RAzNxBin+A57n1BSyWK9Dm8tNEHxgmo9+TqI/aQI
33OLccMJFRt1cSFnBkhMiVD8kCQVeO39+9itJp5sRJGiiMRNrzCeODBGMB9y4okj
eRcd4losLMzL4LRsH/yqwyDKUICO2Ag42AfgC8zTzPBdFIeaj+QbJqFeinSdNMuL
imM5pDMUgRHxytZzu9BxkXezIWXw9uE6Wc1VE2rFPuGnW9eazXC4AAzqqu2eO/XM
S64DosrU9bEGx5YSi1Wwx2FIHmdQVMZF7w77MvDItU1F1yLUNaPes0tLlNwkO6Cc
4rPvX/XP2EWL7It9TIfO4ddoDPiiG1RBpb9WTvM/HE0Mt+vTDh1kJC7OtDDtJ6r6
2Yq9TjDy4EP0jhjioej1CO1sFJcm7AXRDcgNfLfR9mZcJ4amnvGGV7KIYV/U1qJz
GgiNxvWlMTJHRdeHHy0hQvS18XiuhLAVsHVbqQF1sRZPouRV+wdtYHIFhKVJgU6f
kPQ1ntokztEwPDTR1n00hYs8A/guuOG942Xuzr4jtMsPgX4WCbi9yTvTdfoyxAJC
882OsSKCucOQtqQmweiH6O9RZsMWN0ikkz3Xt1Z/M+yRwIJXobV09wzO+Foa9Ipi
Jk+8uT9LeyWti1DINQ5aTfuNc16lht0oSk3q74lG+ef6zHwxXxxknz1lE64xV4ng
EIxpZqa5kolbjYBWLw9o1JElUSmIBVrIp7RczeIDwRkGdj1y2b9rorwyAMEt1Elf
fDO0MzCBg0VhxPSwbK9YezcyiNeBuGvUpVTsSvHbABVswHbQry2erMVu3CPJt7j9
q4d9ei0HpooAy+IMAjqYebcCycLhiCbjuX1GR/sOA/f8EJq9t6Bs+W1VLVg3dMFu
6VSXgppoJa27pZPGZFMYpOrCei8ElQcQ0W0TojxC7IS88CfSkn3GNCh0K+gI+dge
gDEioTnvouvhk1m/Ue8RcoZWN3pQP98JOg2KPGpRFfz+cRL0WqYxecbwVT9u6ryf
fwZmlzUzzu9UtonXNQP5r++gPDVzVaNX0UDi36Wbpwl6j1XkrtjDgI/B1+90ftf2
tjX8nCky/4KyCeZGqQA4ZuQWq63xH69tSxTxXIXla+Rt+vgUxYzK4NXDTZERCxg9
kt6Wwsb+tuFGN4sUGnmuwznSiEuNjSpIFUUVYxD1Ds+6Di9PA5E+g20nZHJQaRDp
14zpb4pBl5VtOpM63kLhL8GWWfavqD4y/aKOMWuJduO58DaWpe4oA1Z0F0KrIU1X
CpUZnNQqNfvK2y55wjJBADO+B2002pow+1iBkZqBrJYj+zuA6Vl2fE60t2ThQXf7
hQsacOBkDTXxYnGinme22OBqlVk2m9jm3Td+se1sl3Zvurq7phOQENl/rx5AsiwG
JKsi/uEVy/bg9Mf5Lbr2s3zaF02xShuzKCyWoR7Z7+WQWgAnJ+c8yrKJ/Z1i5gjD
o2SzY3Yw4Mfz1L5H9lIBCoU3UBxTYrVX5W2Lus6mw4FmSo3B8FVGYcMVMLuxL3Bn
giBZlwzhj2wmPlbtMLwP0H7nqXyjtxHsoZwy6tYhi/c3L4j2yuDOn82c0n2MEws6
OrHVpYv0opv2wtMYNTLXxPLlVc1CtIuYOpjFqCy+8ZPAwDEo17lrv4382blZmi9t
mRwZ7Vru0GxmeIkJiXgV9En73CMxmTc9WdjwABhiQCV8t7QinZjxmgS2cc/8oRqC
Ptofg5M/WCSHPT5byTDIyDItCzzqzyMBrz4mPPCslY6Q4owoTK1XpSP/te0Qp8iH
DNzxkun0U+7zXmYyuTRlZ6rxqI7QGhDMOiXmdfK/lIHcAMBM709bxXvCTvLWh51x
jrAR5lbQyGzIKTNmuyyeFiTCkuw8tz9TphKBeTvRvWGWU9V4XsPtFC/Mkk89EbsA
ET9ExzLu9cbidtdA6pqZwK3CoYO86NBPcvyXNVy2BkSGJaF6vBgmKPTlu7op4C/D
/E83qPyGxStxMSUu0EX6WPys91xxLU9gOx51QbxjJ0OlJsuqoT1hnzmZ23SQhYvy
+5SlEokGpP27Ufbx4CgaKntGW/Djy4MEXepx3cNtL/Vv4rEp1WtEPBw2PvuR26zv
7qC8tWpBVMLMYjE3fj6Ts20/UyiLl1Fm0xU8E/wEE5lx/WMy0kyJoqWoUDwimvpQ
0zQzX5t/hVuzJt0nd9p96XaqrrAmkW+F3atSWzRC2d/fotM5PndbtVVx6QKUc08k
YB03EZ2OTAhY7OkGPwvhl6d+v+DyNDWG8sOfnsopdASqdBKDHsssLMJaUrE7vDau
5m1V8m0i29KruMiXPtjH7WvMtYRI9RRQvOMmL5ACadg5Gse59/hav/PVqtR/L0Bt
kUgWjSarxGf9QxZQXP+9IfC27JPnVgBzLNunW/f4Q0of6deOFUbKpjpFOsiD8NKM
7W8lrUR/kha/FfPHcTJuxzH/y6EQhuqKk9lnpd+T2SvkLCb/DQ4pCQqKx48LUieY
h6HNQCOrmeWktwX402btpcpGVz8+OD0IAp0eh25fLDx/Y1WLSHT5rl+26W6XJFTN
J+UPzhYtmHlnOwVhUOutTc7wYD9d2HXxWmyljYbyKLQYWQWTuh5/LFb77eQIk4xO
mRbKQRNR+kQExq8rwLDLqvRTMeMBWYLDoydFt+GPoFiAAWEXoDh5dJP6RyEspvM1
ze3W1rLq5mxZrROdq1oKcxTbBxM96pp8rrCKmWHzajT5e6CJM4dZSrKbWPPaEZPL
WZE3TGExbtaM7UYPFVC/21nowWI508uupmLI/U7zg7D18XsKNoCCDQVu8Q3RwkcS
V6KiLUYyCUP9YHPMbr4ihv1aP6ZwNMAHLuZtsbBfSw4evJN3ohc5ukqGgOvDhRmm
7LxPkhXyAf+klVINyS7UrMBTgD3Fp9e8VKXTNmvpd6IHS5d7biQil1HPuNcw0ygL
ASO1iGFyKeM8E/OJxYINXNT4k6Sm077YuWfBcaiWi1D/gtyiA7u8T4UOyW6lv6a6
rEjCpBk+Qd5j154thhKzyiPlzCFyJHIbHibm5J5PsAFJ2yckE7C7BMmiY3loDSsP
hZcxhGqtZ50n2Rw0PldMidCGhWHFt4qvpAqbgmNDPS27a4eqNJx19f8bQ3/jzaxD
Wy3Y2eXjEg3A9SbSUKuNviCwz0o9zfBJyyuF84GMWnwsjKLh2C0SV/oarfq2grOK
mgy9PF8SlZeoJhtZqGaP/juUYDMptrtSOdAFOSLogSIwiHw03e4pPix+QNGqK2KL
d9aacxmGeh4HVmXyTKXH/NBlGkja3HW8AFApja73vlGxN7BywXzBtAPc76YOiYrP
8EnkoihlaxfrlS+xTaIlalxaqmSqIdSEUTV3hSHWu7TKpPqBxd843hsL+yxdSPpO
p82INF6hy7mre0ppNOlj7TZuMV+rRXzl0f7JcIOWwa8byW8xwusMk9zS4BwrHwYr
SchehDoXIX9xB6X6GQ9rJqc4GePdN0O5HYdtOupgwNR9sPzuNLF4Gsn0PCoVMVjI
2nc8CCXUEYqe2xB1twJbly9irRtn82ypUqX17oBpcrtNxMzZs/5RrnqXtnKzrkZa
aCdk/4tjhpGcUEzlLBrmfW/rQaXHbVSnUVxk9Np4+VAfrbOxKBCYF8ilwqoNH+A5
Wwj840HcrnfJlKW8ehtgn4lsqbWgPpMEnPmcPmGdYXuoTWtdU6Kk3dCTTcYRwkGp
ROi29RQAAi38iR1LX1XHh+3js7RKyQEJhhu5TYwy4rqBcFujuZCY8hsQ2PW0FTe/
DaPHTvSGnrj/QnJNGIBpeUVdFFQj7KQ9ldN/itZZGvfu+CaIgNSxS3xnK4I5gax4
G5aGjNa2iSHs3tjA18QyX1VXm57Uz73iZC9Uw3RLPJutEvzRsH3GQ6ruYkdA0jr7
gky4ma1L2gxpAB+bJ0lG/RWrcgbtoYT71VCvAW4GoCixvvQ6GhYN5LtidDYxqoIW
ZEFMhRf4HWgz7gvpaOQ0g2moGXQivoXIR1gUmvRqk58pEtfsesE2pKWuPmMAdLye
QYQjyZAECT2A/Cb12g1kOhbzk8i15Ui2IhJmYAy1B6dWedHrYl3nHCyWl1sb9UEo
H9GH3YiTKTI9nkXBPPkLniheN90uFfnMLzpeFZexwtVt4jNLtQ1xDJJFl7EfT9RE
WMTw5Yut72GCZL5q9Fj0N9Hl6R0H0WbLZ9Gw7gGTBPFeyQFBlUmL+DYT60Ydzqvn
P2may0ZfhY/GdSlAmGD4TmGNHzLHpqjxmJAaxMjVn0WNkpQ5wtcKioZWyBzt5UE5
wvb1RZtSashaHECFiXvlePgxK81HnFr/FbGle53iox3F0MxS/tWe2xlB2G5gUIta
mnndQyXMdRUZWl8lPrGRcm4vxV4qluqvuWUCEszcpwImOCxZVgPA7PaIbbKpfLU/
5ll8D2hNVfZ7O1SszB3+y4oTMAYcDke/raFCs/LR65eo1QRraR2J2Hw4waHoTyvN
nJgbBlFDlCWckcGkxp7ADiTrND5f03Y3662panPX4HEbF8f41kGgnh53BPY7FX7I
jpBtGZtGCZxfMZ90ezdWUcA1+ccNSrKRQdooDN2w3PcDJUkhrlckYLOvcPYKxHhe
uRdbp4VP7BS+w+v5ATtbkvsHvv4q5mnO5TZOveP8zmYrAhYM6vSEzaH2iCLnnHYy
WF1d+Exfh7QUN5BVDEl64doo545IX/OUQ5EZjX2t0e//OFbgEosybH9Znp9HLfnx
1jhNNBDIqG001qqw9HxzwC9pWI1jLzSSMuMnBL1b2iB3fwYDZ6lK1q9959ntqOtQ
uc9JfGU7nFTNbLBh61KCfKn0q28MtS28TQ4Lo3dM7dHX6k/H2AmS5JU3S+r2EFJr
y2E8N2L7F/GvZ1VieoIWRrsc5FO/b1cTJlYukQVuvUgdfG8VMsLNOqacP8CKkjdK
kkltsjm4RDyFNM1XnTQmNMRSW7FHEmchCKe8ww5xbn1U5EmuNYl7MtFA5XOfgSjT
paRVTlrOUp/o4MBzcl7CTXT6AFyGouGrWyxPUCpFn22ht5b5IkRiDO9qHFAJi9Bj
fWvJpjUEPsOIJNAHpea1YeiiwHg94c5EeRNRYet8THzt7Af7ojTGIsKyroj45gzu
uZcIYOk4DkLgEW4rXY56YDcog+JU353EdLIdpQg7FmPcD9AeJfLKtdgvwRoZtsWz
oJ245DvLG/JyV7SkeFrc7byJdox6Pzba/libYU6G4nmhVvEpELlcULs4/FCIWbmn
cy28OZoj9f2nosTaDO+fKeJSBMEkX37ZMfvOkZtzZRMXqanHmYqB4ZRFtyXih7RN
+viqm1bFgG/+l0gFoB/amg31tdnbZWViKps8KRTYnPFeT0wE2Watntmw22ALCFgr
Y4EQGz+wdMbbQm0b0hp0UBhGk7fCZHWm1/PELMZf5sa+a+jefpJCak9U7ZE70as8
DmFhLBf9wzLkBfL6ESDYA/jR5CUrahzBnzFlz8rXg2LS1v6FhzroAunAm1lQ1D23
eMLwbENZNkeMgtb+ogzYdIveCX6yIo+L8bREtwZJ8CsEGHa4NJOqQvmt05zMjQ4q
gU331mwfNUhkuLBRmnqNFxLl4vPIu7x85HiZ8CGzT//9OB3PLtSn+NeXQtQqmAXq
HbWRC3TS8Prl6Qc8w5m/fNN3+RPRnbvnnFm2Vvn0B+Jf6X0/J24piaP5vzZoUFpU
T6+rQITyAcC66o7Jo51uwS+qZZW/G4XgmGeTRDaZbXJVA7sKMZE/MLBU9yMdzJqG
ubifcdpUMIXEAfMuUXH0WA809I1JOUrkQCSEQl9KjYg6cImP+jDZJGwVUAEOnhF3
lvsPBJes9sa4KjVv0CPalgl5iNZtYYe5wfwsSuM7Eo5rFaomdwEBDw8VY5nfwo1x
jigjvq/i8tCfKWV4J5+DPVKUAFvAJ26tX3OyNa90RBVDe9qTOwyIXG0+pAZG8Wdj
0RboMOwOVSLv24dgCuQ3Nj4vJkj+JvvOSKMwbyOF5Y0BHyjFqsYwU2PLejM/1cni
ncNBBH3mHVAVQP9ObNCGnPKgA8et3EsB2JlhEGrux6tyYj9Osy8jvU2b4CfxSnhS
KhFf2SajqK5JIUHG0dIO2oBv7Ld485/WHb0jALa4Aiak+r2bdo35iKVJe0pPrmzQ
UVFFMt09FIhgxJJlsEc9YJ6/b0DF5YrUfAhXobQ1zw3QDH2BCN2W+TYw87yy/W1q
+UmBlQRNUtNaUefbU5KrbBiD9bv0C2oTzeRG3hg8tpGBYGX5YtXGeTPWO9B5TBoq
h0X6jUIx6RTAMwaYB6qts4hZ+0dP0AFZcWzbzDQxJVEhGlWVbQ0zjPgbKGp+l5Sw
QT8b4LnylWKfTHR7RiwtgFENoH3fFlLfXJDzFRwSl6eO46JDOYShbPzbVkuhS/tc
p+zJRSCWjvPb/+FBrpw79kcaWGOotf/s3U7ZPNjMAgZxMavTLdxN3WT1Qojpvq/Z
sQ/KBSU9wdz1VFmfe6VbgQk6w51aKtiQqxEuxidhPWtFmgWiEKYW6SkCL7f3HwCC
txmZmvPyc6XcnFGQe3rV29h5YtkBD7g3xajaWYW2GLjBe5AynxwSsGAtVqcPa0eL
W0An9+wvIdPyl/hw0c3K27MuSliMh571pkWy18rM+15+i8fZJkoVr6aVkB6v4i0z
t8vv9fosJymZYiy/kvyFAPzjsbTMDUX6qi61R/alNRe+U9FxTPsHYk2By6tERp6x
UBjg0ozBy/GHMFMoWmW5IEg7eYLrKgExjJyLyywS0ykfdo0U5qgiYJJf1sRhPRnm
V0Xa+qJmApFlrakEt/NjK6XBZEaLegBe9v3oPitieAjN/agTmg6CqSpPA9ykJAbs
k/49m1Bsr9w1zKquCYoM7bkV8zPWN4jVblJB9zL2r7O5NP2rXWxiAUrxtCQ4rd+d
YEFEKg/fD7GSlYd0KgInNA6qWHOOXXK4bFMx1qvFQRT0khxur1uXOzA1fa9u3Hkt
Nxd7OZ34gqNnIXnnV8dHryisDLOfa3ZbBqMPmta88I4C1jxiO9Ym/IoiMEgJ14li
S3UTft5n4AaJERWESjqqevhSQ2koYPifDinR5xuoVxYH6gIO6kMDnWRjda7z8aPT
XHEGvVV/jrwfj90qPHFbv3L6+S7C3HwFfdAxU61iuOfelROOKFJ3uAC/IHUwgPw4
x4fLxcb0PH6HsTIEAsUAYesaS8JcFNC0o0QBJlq2KQnCjlpQPKVk150AIdpH1Cnt
D3jWYlB4p8m0WpZmsXmn5ImAPtOF0y0uWcmBddHx1RFyxhNCk6ajHjfNBjPAKqbF
u/JSIXFbCdMokfhLvXDc5meL0jL1pPkWNsho7Xh8PIKcqFRjAP+nkKn7cAFuNr0+
Ez2E2OvpTfwV2cQM7FWLCfAS7RDfiAj9hKe8WRsaRJoyuuTqdGb6nkSHaim1Sk9T
idapDdHx5Tf1tTMM9pvJH9ABnCbm7mziOb3hjkMnyNogDVNVO/8pJzQAHyh3SfFE
yrb07RnUZycovXl9CN71YC4CecwafVhS9reV+Qph1TPfxgki+eJSR2RCWis217hE
XVGk4/DikrZGRNDg1Ybx01xsJIRdwX6KeTwicAYNcliBPZ2Z+6X37wsUrJVzV8rr
yUluNExmAAg4AMYhTsOjrUa9DIzvGkKDE9j1DryWccgjgKUdFRo1TFwo2hZQD1tm
ae/HF262hOTUMo+nUtgCb958fNBr8v0gDPw12Ne89Lxc2G/4NbvNstGEgkOiRX51
taicEM5F3EP/huClQRifo9UpjbBOuc9+Qe/st9caSKmJMY4mkg0wygBQvJyvKlsk
LAaSN+4YIXx+eI6yyAFW5t93xufK2+YAFgtwUoZ7twz2a5pESbgVFNX7WwYR3iTb
CG5ZyGd78AT+X7INgrwj5V2Vj3z20tr9FTyhmi5pK9IDN/2DBixPY5t25PzkIB7U
UBj8t2BVdayql2QhOMcrUg8UMf0jyh1eHfGedGpL6/j15o622YH72gUy55KX7SL5
2asebnsxPbPeJ1x+SucQuzyVhhMBSMOCCxQRdv7eQvbl+aX2nMr8CS3h9KYMuuqi
rClr0Tuo7o0J4ANmiQoxAh71zLKx2NQdgXfGYnAESDD+XHjr7lQngfSOnnxaqaa4
ivJ+R+kBWiP25sM1DFrqG+Jcx9AbICuZbA+XfoZbmjow5Zz52mlNmgzy318rd97I
3kTgsQCDyZkQ0KbouSQyVwwoKZ0sVQo/onV9R+GThwLjCT7P9pjPVoylcedP/jDj
cpgal3m7ncqSQA4xi56zxNwm5Eysk0c/4TYQ6FYObprguRaHwajnNx141NeMcl7X
24Ana+EwhuLxo9phyh3AJbCgeTPrzMFIDV9uTsyL7C8YFILIVp9ugdO8r5vJAe/W
Hjfl5tR5tGye/c9Czd9bts/EovWaO7IaXVPiccf9VEJ35RhP2ICGKMt2zuzFOmvh
Qf0SEG6ucKeqgW4FFaYnjYN9guXkqxw9aPNndOLH9UC8+JeZbwTfHqd2cUXhnliQ
81zQT597PUgE7azMooqAN9RHKiI1EAmcCpgkQnSF4CGfCKmjyOj6NF0z38/AEjx2
WiKngkRSGm7pcAquAqyxU2F+hAouHDkFBWYNpW4RqCVy+vx6VNhDziUO/ic20Rdq
NDbay6s3Vc9azjZbaqNtq8296JMBrPvWuYhERyhT3t7O+k0LM4996Ii5G3oWc5O2
cLXpYhV9uhDZJ150ROyZ7lnM5370yHqi2iiMQWBiP80cNqMfCHR1cajlvb5bLwHx
LZWVfdvaIyoO7LNa0pDXh+ClQKK57AqhkLX89GMAqhUPdK0jH1nzoCG+C1Jinroe
QmdGAdwCdDf7V9Bmevh2bNmfe7COgpLmoJb61x8lJbxMD/4yETatguXbxVBCD5b7
DGaRrSJKLYzpjlPdoyXNnSxeVshIbyMJU8f+O8doD9Ectz+AUAhiG8EShjivcfBy
Y99+T5kcl8L7zy+6sfzh5v6BX9HtBZlqHu3O5ERxct0kGUOm5RwB6ovmNoUVN1xV
325vWmknUzlZpp3yGdR8vU6d3+yBxBHTIgLVMkeI4bKD4/PLXNCI2T+9woLcVdu1
0fPkU8z3RmgXJdfljbK6+3F62e1UpZKmM9ruDk4a3HfcIzb/e7oHcl/Bnmep8dfQ
ZMT2CT1Sxz4obidXzitATvnY5T+LbPreuAZlINh0btOPACjaobrY3dfuujcxHeJQ
TuVquLqqvrssTEnOCAV6XITHXrsNvQbfjvWw1JXo6DdKi10SpqL5otmYrUD0ItMM
DIGxGoH1S71gwOdx83Gbpb6mV9DvcsttNdh3PimZbxC4hs4O9ZAXR57PPjEcFH4h
QTBTwMykzpmY/euavbcz56Exu+QdDwO6jfe1r+e3QZ22e644P98e5wiHW9ANxeCT
ohgvzN2B4m5PNMb7k+pOkMTLl9CCLwgflFgMkx8/KeJLI3oBCbCe5ayshxB4+tjw
OznBpIY52dmoXTYsy9hfatSTtWiwX8+xDVe1UOhBfPjkyi3/uglyx8w7Tvtjx7nf
uxPNPvsu5iSocHdYZTMtQ47ZKXbm6PoIMFVj4wQQ2sYspMBjHTFspo8TOAJ17O/5
6ncf2ZNetD7SxA2KKiumCfD/Ua9JQgH5iLuEbJE8IbTXQjGPqRICV1NLaArAukR+
1X4jGlKxYZiWHJyXbcHr+s0qtz+oCrD+getIgoBr+lSlcZEiR5vsalMabLDOTwzM
zFDf+8Omrf4ORTBqyGZ9iyblRfSpr+aRuFETqXhzJG6xFA5+BSUTX7evoC7WKIob
tsRPMIP4J4oceFCbvokE+oHXtPd8cE5bJ4PKHedD0wuGmmkN16+HIjjATBaXKUH7
HKIrYnC8+zlfYS+t+glfVJ4Gck66bYnh6Of8uY+Ap0VHEshPsnj7woK8PNsJtTQG
m6ToOfCvnoqsa+271ivdKNQaX6gI3aUQAKFpbpUZIt4A9ds35/9gP8haIq5+Oxsg
B/fi+KDGnHB1FcP970HJSIWACTKOJpPTFi7wspOaB1AAwLV55f95KacBCJcCt7A0
JmnKhz006bhny1PJ3dy2zOo8wyFl50sZ868k3jNAEzsb9scnLOG6fsGW1yLWVblo
sUSYhOS1oZKWDeW/mxAW95CFNN/vQ4p6A+fi/BIGiGVZ30NxcB8rxBRKovnDHSlC
7hOIbcDZgBZh/nY5M3EOYbetfr0xkAl+2HTXDSIUHeDzwU/3DFFtaBiND9uqAxpB
CLkOSskPjKGq5R1+2c8HXtxy4Ggu/K42bOQxqCDBrxVQv+u7KQbn58jLvdXuhKDQ
DBC9f4KkgbDYCpcF23jiJ3wNRJPaorWg7UzKKyejUsNUyzgiG7+JWSzQSdkMbZkn
lqxE60mA5H24ZcHk1FHXXcIUOOpvQBM9ebC7T955VPR9RYU5d8NKuRasQf2n1rD3
uLk9FKHcMLSLQxP/jsGA9DE++1VP2qLxlgMDulReFKj5k58jnbNp13Cc0aW5GlHG
PmnlvSafSP/MmYQxc4BIblTs+KIt6UUJFQYZsL/5B7tvXMo/DHCpnO8BtYmb8o/y
fKaAGk1olckJc+kWho/LzJpROdkyajRgsSvAesAehGMEVSmrsHI0hmzw4Gg/Jhib
tvcCqEmbWeNkusmqgtoFEzv0lB/PoQCzJTG7MWlsB6BUK3RTLXezY+VeWJc0pj4s
fhBn72qZBrxG3qTKHC2s7EQj1ZhtzopO4iRZ5IunLH0CfZEXEgPWIZhju484EAvk
mv2vCHMNJT5fW1SrRPoFs7cbMRy7CwwzPUVaxyT7fPBNQiiSyXFor/1zpqVzol0r
38MsL05FGcFT9e45hZnXj+M+3pzmOfiYMgGX7i2O762EGHH4NWGS9/Nzyo+zcCAI
8EpA6trA395fCLInYxU81vFv/K0YNufxVUVLFgwcRGRYg9FNuelSHqqtpLiXuYcQ
zQa8hQipHcMpasE0vCt8tm+Yt7+NEIOXWqTG7u1xOliDJPiP0dcq1ZNXw+yHboma
tqE2qLPljv+m7gDMWUxOfSSzb1Akvba35szSU39gmI17WTvicJoGOg7g0uOw3S9y
NR1vT0/+xs3UHEha5yF44aYFvkLV16n6hUl+jR4VcpwSGh/iCRbdFQmQZW7xV/UC
rxMUX8aa3X6fTfOp/67faYQFRAOvTPszgNCojAfbGTGrF2Xdb+b0BFTrWhlpeXMf
t9jnwZb8FO3sw/6dfiOmVj99yvpRE7DU2/rr/aiqQliMYhwiiOf/jwgc7a6s7YYi
bXlqn2kQMo1XJLjcYah1k3FjkZZZABu0W1C7xLw6RcvSsZogLCPP6ThuPrrLKA2V
S2++FeQ5lbNTsRaUyfA70AOKoaEO01BYQr32X2r15R8F+MqAyQgnHUfS/p1m2tDZ
3yy4qB6YhOpPtflkDTOkMqZXmzKXXU5GuLgGhPcRc2w9HXySoC0HmIbJx8NRaDkx
0hbOO3y0xwEUNm9S3K/7tgCkzcb6tq/FfyYE7gbWWV4P44ywklybYu+TEy6GjJZK
Rxh/gXHPqFxWxsSeR+FfmjqXqZFfzvH6dZ7RmhKeDDj31d8rC77gMvPrXC4aqdcH
gClBrcN4mITzOCwHrmWD67blFj4Sprx2YLgRK7KsWw6XqN5pnr/lQyPqsm2hHe5q
fbSIn+c5Wo3HTQmSXZmAKyDVoVyOLzStuIRAfwkzLecVB/SXJyebvdXiPqcEWlE/
FB3BtC8yGr7oLkohZVPTAw10WMssWBmRbIFVb0HfglA3vAoFAka92RZ5fGAl1O+M
QwxlbGOUucYKIcj8kvRYR0n1bT33l47eX+sI9eRqtR7VEbum3U2XPcozV5dIjd5O
UlhrcBqey7RSBL17IIoiokfg60cAFzFqLboVw8TimfQY0U30R1AWAzihnpvYeQQy
OzRalNZXaAubYo7Ajd2w69bi4U7R8Ox0ySPMTKVx8iZxmeTavW/DAnclY7MTkLrX
9E9t2cA6j0fGjeqUzUxI6pEvdC7Nqf9bnliObLsgqLTV61gmJ+VYlon91AcKc1Iq
ywC9JbuzTdRo8UdDOvLThzHqrWAHDuJM4v8U2M37kHUmMZb8Oe8FTj7NuG5wyfTd
tJpkZ9YGD/cOR44uhC0lFvPQ3pRlvws+d+qmDLWGspoQMH7BMZ8tDZMkwN8AY+og
1MBUo1vFuZAwkyXWq9szX8CXa+JsWVtU4CDhPuxYr5PxFSagstiWGQgfGfX1FTcA
ihpKfIseZK4Ry3OcQSSp1J30/vT+YBKtSsiJ5UiA+nMCsWQGfu8YoeDUZuSdWohj
1jLRs5zYUslWImxcC825o3RkL987nQ2awnGUM7TZk86DUJcmc4bXLONmEy7uI53E
E0SCVyc2TnuKActcRvFOJGb1xrDqOmlPgjE/DVxqwzrFZwP5PsunGWM75mJGvlkh
tlKbSZJLoSeOeXQSnLNMwcCUxXCV1W3sxYBx47QU6hvQSpYd52gcBKCcuDc6aTox
zfMqL2eNHRQnMcpJraKImJ6erCyXmb37P33N9QhTOmqgov2lSOjGpJNBFpuU8170
WLhRq+xPdm5icpDnjh0zS4fQSVrgfD5Kabo4vFVq9rYhEBqE1Y8so2K9z7EUc/sg
9363t2pf1ygHO/hOtkJqUq2gddJfBdAkmbWfjGspGtKtGV5/gmJemJlNU7b4UFXp
BHTSz1thKZoaDzr/fA9fUQEgxKLHD5hPCnjX+03hRHP6jVlbG5Rs0o7Os0aOeI57
u29IewxakCnTeHrkCFwpMQkUWOFV1Mpo+Ibb6JMrECQTKdyEOYFVVpTNLTfVRz3j
Gz/Xoq3nG3c1RRj2UhtBWsmSvzzZqRB6+G2PmcLsXtLLphyfuQxRYhxHJeEo3XzZ
k636qGGqPDwCS/IFzuDE7EphRlGJA+hnI3ZnnarvMpIaKQdOtr3cVWGRdRpqEOQg
jrc4lhrVIMGPZ3K9Yq22hgLLCEvWwI/lJy0CY5LnyI3loTVwYrWuFdm4a+VcJH3u
c+QYnH3HE/+Z3PDiH02BFhxXgmEFXIpsnb1TSFqV6ighXNsnJQYKSKQH7rpBSKwO
qIp05SNGOZ1neuV5w7QHmmGhZcTZWPDMgo07gfNSA/SqBhGMs/3Gzi000GKaY6ey
`protect END_PROTECTED
