`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xNV9P+9DqQp/h/eJVy9P+TiquxtuZBh0XKK0ItjZYi4XLxFkbusNBaAS/6iIqM7
dg5rE+Tv3wFxYunblfhdUCTVe3zWho0EVo6FgOTMxIsYrWXw0Q3jTwS7ORYgbW9m
Ozf7F/pTNqpjBoDkalyUqJVE42rRvqiOYid4gah0vTIrZekHTPf6jIxzAbhlf7hW
JqQqGpCJC8w/1D7HAYunfiFL3s+XlOao/gEWRDOzQGTl3z2dPzdFRB8JwSAlVjpN
H+Foeeq1CBFS+geTjAPpm+QLmE/CpbPgCkJwGyBhiPA=
`protect END_PROTECTED
