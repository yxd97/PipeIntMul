`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+M5zriOD+9dE+4pIycfw4Ekor6wMHzUQ+j4QA0k2mbJvafyhcOS+8VMawPwBsnz
r/amn5Fu8FmDAcchlIBH3gM4YpS5FNqH6sZJB1JkKH/EexUs8+7HRcrVECC0lW9s
gVAtLcO3aBITTqwk6jsCbc+0nnw596JbotuyxyVQOfKLm7jRTExg1mjFxMety6hc
kCqRsG/qzwO+u8iYs6ztnO5bAaAprjmv9KSPI9lyoL6Tpyhmp/LMJRgpTGdBfnqd
3sqCXIeLrm92l+1eYFlSU4i47nA5HMgTgwQ/6t2tJhEyxq6OgC17xL0Bk9E9JK/R
otl5gIX7FBGo841Xh9mV6w41eYu9303ah5/EImBJMBfQ+MChPONZnO4GczIePjrj
qb5OKylP6+IrLm/gvAtWmmUl5CrbTttmHg8k6WuFjqb6R+zTKEXdvF4W24yQfSxo
`protect END_PROTECTED
