`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7P5Wwu+2huhdqSkxcNrDhiCv9w4LwvyuU7I45eWinjis5dR1lfmin1OrrYWwbLZg
o6FngsiSNoc7d04sG3NPb7QN1pjrDdI6LyzVKznZBCZIJWKxPzM+ZwqlzpkadrOT
uBQgGzD9a03qpI2JOI4QTi4SMFTduEKAf56SGriH0Y2UqrHueIK0Q1T7Xo6TMtuL
lY+0zKKqBGmH4gcm6stLno7Gyrt/pPbWdDPJcUbgJTdWpj/OJSfoECC3Mq5iy4e2
WayuOu49uN/rUPAHowiAXlmXaOjZiXw2FO//2izikK87RPt/EzAjSloLNKTwRps2
9rS3zdNzRkLmL33SuVuzvFQsMep4WK+DcEzVd5c1Di+IiIp2Mh3ifnY4dXwFfoN4
gs22yorrI1EbRM0XTIeH+lPOLCeEleDltf6aHvK2gM18Iiqvx1XI+HjbqP50A92b
6ENhQWNNMwlZaeR5vbaGFD0RJ1EPjMo2pF7XyoxEKkLa+C/vXMqZ365zrGNmrwLf
/+6UszLKUh33XFiFSI+quZEGvtVPsq92U7YWzr3sI/T6u7NoqdIBa/x41szOhpTA
aaXeUlLCwVDnERG14+IXeLghBgKBQkVY3Bf+inQPrt5ctjUSSeuMtyitE0MEPmn+
ZbaG49dSoBIw6jzLlJUdu9KaLLb5Pgtobtb8kJU6psZNjdE7Q5tWp7wwxvGrIi5M
EdVUDLdOYo0ehV5iBzawWFTSh3Mvs90gR9bNpMWFroJHkl9A/bnq8kjpwrhjstl7
Moy8vp8P8EJqkBQB/hoZuWJU4qyW6nlY8aLK3UqWvQg4Eh8LItpzYd+usVXvVb3u
bQ4D/zGvyY9194eFP4r7LaPLu6FJiPPKG4j19dbhSDU=
`protect END_PROTECTED
