`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LEqRH0QoqeEVl0XHlHkahU5Y4JKWRs/DLMY5N9SLGuBDdHAMzgAYUmJiChFDjaZL
qfEchPREgwl1JsXihmMVUfUbmlbOVc0WpA1kKepifjYUVcxYdyL66kyhBQIKdkBZ
o93GbwXw7VGvDz6YTx6tsByh2lmBpP1TtNZSjr4+1CfKnxRDukqOpBDj0MLYWZlF
u6iQLo0EJPNBerYRzuJun+m7/B4HtEgBbIC1MGokOwGw0Fgn0/NPNzxZcyo3CxR+
Nh3YBc3mDTgT70PJwgoIuhshQauLyVCMQb9MVnjlHFESBETjrO/615BZVxlerWYY
u12YAbCaPiglvsZ2bsa+VAXTHBCi/wSdbLBlcVc0wAWEq133768miHQ3pQWVBzoh
3D/M2uo/0j4Q84DMLfaM+d8Kwhb/HQGxvhwG+g2LNZjL48jakjsJC1f4gcyFo87d
+mZ+Uza+H+fTMm263tOy1x/dZF9Z07XgglvUmkhSTXMGnoe+Mij3DUzTlgigrdLv
L+rC29fBTmNk7X633wnJzMsZCeakW/XRCR88S4bPv3Y6dY27V6THG6Mjd6ZbY8II
xd/cHCL8UEmbLptyq/mtoAtXpmu8TAbJaOk8Mv1g3LPpA2sqXaW5/CD19Dv+DujI
HUruDv/ZtmwgUUvTqFPEqvgfn0ilLJG/2JKaUxYxw1UKyYGEtxeiZQppcEozI9cZ
ACueJTyx7/HZkWAKd+tFvjkOdsjpKDaZsfxOrHUmtMykVRie20TkmvzZZmYzFgYj
HmE6Wm8sQ/vCkDAWsUkDkUV8keAAJHsT3TAMPqnAuyYF3wO0fAfzXUo/jSdtXfrg
aNrkrDyTjJ8Amw9ZVnA1Xq+bMr9a3Jcdvgw/EZLQSI4IATs4f15hRHX5W7Eiv4E8
UbfaF07OXhtc/+MDGj8Ac9Z7OXbes5K8c4u2SrsojwgRyTeApwQRC7sQ2yikKSE8
Am9+3ODhkj6TaNSELfy3qE2Tt6URi6C48qcy3AzdD+f+7EF+DV89FQXw/GhatgXp
LLdOiJVtpVUEiU6MflxibuUDcBKc+QS1RhiEw22Mu+I9sA/ud32X3pzfmhzzLwxI
wJEtkHWW1jK5czII9jyZjg==
`protect END_PROTECTED
