`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMg+izirZ6lM+ZRfgBQIHvl/31tQXIv2AVxa2UZxkNt04n5GljvJkLoTNINb7Ki6
rCvWlauSwfbVFLeo+11F/csq2dflY8qGQRhuSoBdFHH7bfMaPikGdenzW3+lX9iN
E0aodAlxZCvCkPAPkc4QNKnTZqdE35R3EZhQn4XYenLM8OboeEZ7stdkUGSIG7vq
LWymxCqb/9rhm556gSDujX4vfHecZFc7ShwEuE+zCYzYFXxAYzd7yX6RurLx8234
P398s23at6CviqHrcYpPquUx+b2ECSitnrWUMFDvnX+wov4pAagMUvgxLiTRCz6z
F9fnils3GJdhC9Qsiy3jS7Mx6UWfxdgP+V7w94gEfGq1xI1CtxP0h+IFqKhQpVrR
Bc/tTYvVVfetUFjrAlAib+y96xnjRpkhpo/D9SmE5Hy2xCMb6KRIA+3fDFOCbO3H
EP7HnD4UZYAZsC57O+sd0miVZSxQk3IdwD670PMa0qmZxmu2vXg2XNGRzFnDZl4X
B4OCjJHBgf9bUpxcJxjEUqNMKLMYPn9PhPfy3HA0KefCTej0RLXKejzKYgNfcz/k
bcFgidX7LAMAcBhbf+fpoi0he4R0H3G32oHPesSmKsp8zPY1Z6HejcfC3YuCgyjN
VmgdSqlh0VT6WNkDNU+2FHqU3ol+RCER7Og6BZ5nVtWhBu6FXRvUo3XxsfEY/Mus
1xVrO9GBVo5moGYvA4AlXElgiBr87ngR52PzI1q0/jjOZm86CEh20HIGKoWiAFtE
VIaSQzuK61taVI/Htb/0a4pnRyA+t0uPL4eWhC9IVbqHjQuNkqjMwjwnbmMXzr/Q
hv/gclnvemkjIkRlrQavTkVTrJtt6VF8RWahcADvcJJZLOsRRn5N6C2GQymk3Gp/
j0ylD1h5K7pMKvusPzVLFg==
`protect END_PROTECTED
