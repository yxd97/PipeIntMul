`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvCXAZgzzAFYDEVniI7leFixAcmYFLaWHUlUe75Ykt/mlzr4IJR0VXZmeNdg+1u/
6bjW0sbxJAF0III+f+JVOfe/XheqwcWEYLuc/wTV+e8oRA1FKUoKemWKJjqliAek
c0ivRZX3r80iJJyOgh5jmEly2yx7MeRN13UEt3zCEoYivkaZEVsEi2DvnaivHMck
7Skh09c9mOz6w3rpf8//UK6hMSru8orM/lHHX0hEEm4+U/giPZLBwQHjMVAAo5ZC
N4pdKFg8YPpfeo8BjUWhf1U6YPM5GKrMziWQxttntnLm0qkJnn1MKvxvZhTesQBC
tRTZNvX/M0x6AvRHle9GhKEF3csA/il9U2KkGyxqZSnE/KIoZh0LaLcMqynKYQFw
KV8VT7VNFRrR35Y7vosK0UrrqqhkIUt5uC0xtRSPhGVUuHTLLwRPh0Ci2XGB2XOg
jQIv7V8UZBtx/ihJFd9krmzYMXexbze+sjFdthoP00JQlhjorqEuFFGl69vSK08s
kP3uGCbfe9ptMHKpE2t6y+YEz90L4qGvii1Hqa6BQd4EKFB1ivelrWOT80RfoCRT
niVt9WBV+ckyDN+7hS/mZB+YmtoQ3QTSoS8hZAquay6ttQD6YJUxOrAXRrepy6Eu
va21wr5pOtO43ecAvFsKuWhfVXmTxswYT9HJkWBqmdyTtDthhK5yn4O1FiGSlP0g
Hu0p4elnWTLheYJ0SiqjEhq4DSPlKGr6MDjP45QzqwYytMrLGzaVP/T64tgaZFMD
mtDoXOXoghjm936ZQmUnvXWpMQx4iINSWAZ576k8YvqNfpZz8zoEYw+xSTpdjz/r
VtsytxgDp4vkoEN18c8eWXRqi6N/8HsTuTZPqpBeyBPvDVOQjX/Gef27MWdzZDnn
ow/gpVXQSryPlWiYgSBaQ/HrjuiZ5RikcPwjkFzfoOQmUiUYb2JXNz/AFs+RXMMA
ijiZnaPSJwJ0dxso1ZdDbf4TFMHUg/k/HdDhcOrpLfCxP2Lu8VPB/7VBhtxcpIir
yiqCj/7KP8/pTLha/4r8GoPro3lpdit+Xps84RuELOYj5XqgzgXdoG3/oiqbXb3z
ejWhTYMVExTY1hfqHRU6X27+yVPIu/vU52KiIgZVcrU=
`protect END_PROTECTED
