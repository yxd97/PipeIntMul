`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fxFuehznPJdc6EP4Mar1u5mZ8x8iD9LYSxL8JecqYSkFbvxmu2+V2XNsnLix5zV8
gg2A1ude6qQYH+3zcefzREzGcry5xkmcWxXR+KuH1GpYT3OoGkM78Lj9o+Xql9E4
L9zvbm7kBY+7xMM7ae2J0soDEw8fJjzdwrKe8653nXnyLw7S7dHjVdP936nxMImy
C/ftmQC3JzmkKuiTjzmFpEUm1GLA5aHkXEmYs0FUNcqRNMGRpstV1/XdjZJTPsxN
BMNUrrSxm90r55OqMEQunzT4a5cAWhBMWqGDzrW37OYBxXMk5W7CV1PQjMP0yBeI
G1nbTDZTTkxWmLwaRcyAYKH6l7XTM9F2qA5+oaeLIlhMMlferPp3fiui4XdaCoU3
p4eli8KZDLJ9Nc9AS792QGVoANMGXADhVdQZQGB5GVuY6l3Sf4wGO+dSx8l9f8ff
`protect END_PROTECTED
