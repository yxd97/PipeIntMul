`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EFZed+RzpZ7HEzA2wlPjOY/VziyzOTAZo1I2CCCeIwaNAp4w8r5nrda2A1N5iElo
Z3JG8tqwPVsaqWxtBSBj5dwRT/LOQUDm6GXsMPneZY3Ba5iDWxrKmMKQbwXp/cNS
tzIIcExVd3ayutkcXHZMs8VUG+Z72R8auOhx/S8uULvJ9PjDtZIV7/pV8eAH/OSs
MzF6AkfnfcDUTpdYrXp6uSRAv/6JofGRTAWeDrwdeYNM6xPS4MA1gDbxCU/xNWIM
JGBNa4GX+AjcFHNYLKnCuw96pvKm18ZYRwWTnY9Dz5w3rob3BQhaSGkyGTX5gBvL
mkxReFY2kYYrf2a1ihgczOLe974j8Yof5vtViuwH6RmRuO0X0KnsUFiJiN7Gfd+e
g5E+N1zXieRE/cmtbAv+OkDxZJS3o3EioU4+kYQUMpWILyO1n88E0YrtZnVb0W7v
Xv/6Xu2AIIHe7OKT1wo2VlCr4VwKg7bu0GoVB6S+aR5EReX1x6mz6lwzoi+naJ+n
yg0CPF8R/uOPJ2LJjRUs1NYiqwyFRn6ebqF1U+aIP2Ptr2Y2+cSo6KS+id/hIGX0
V/5IREO30QMUU6eRUINrHbT/j+oAa0zqCzBI+X561EyaFfPHT5HfmxPKpdwzim1V
PcmQqTXN5QQ+QoXr28MXKQjx3HaglfLax1ff5wfV3SAQD9WGMdl2qmMlyQFpQRJ0
f3MJn6GicLkIbA44y8ZfOfNAChhu+8w9SRXwJAqpTI3VYSKHyW6ZFZM6TCcMkUT5
PgsiapSJcCpDVtlWnuN0B5Kj1HCVWz31xgmih/M7+GxzlT6PZgnhZY5+pPjpD5zr
OjFDCH97F/FxAV5e2beBFl3dECqAs8RZZaD4ZbhSSXb8bOO7Hkg1JPk6pjoB4tFo
T7emr8mP05QMitnUOZg+7hg9IHel3U7AGtOZ/4f8/eWdxsdS5djwY5hcqqOX+TRu
wO6HHRgm9h8CjANAEGzgKQkeBMhibK5BsAdZ/3Z1A89CllHgDrFQbjgaW7VdxsWw
TCSNRIrLMOdC/k/iegy5YrnNGT6sfpx9PiSH4KhP5pM2a+230veqgmUFAU2Kifvk
+2q7uzHQcOKpBzM61RhElF9Ox5DWKZ0PhqSwp3VfXx/0egQC7q0vytb67W4+Mdyv
WTHqlSpMMEJKj3imRDWUUmoxb2DCzFTL9+d3G6cU7YeYbB4/FPN3Pl1MRg6GhbUh
OfWh2nrmTvnzVQLs7FCXUDrwyXSV3+vzWLfnXChDQ2bjZ9waF89N84rm37ILUhEM
bagsFT0GmeGMzCLCXqwvqNDlnk8BK3h6B17PBpQ4QZHR1HWDMC789PmBP6WE52tT
hHkwIOEJMbbsFE21rmcPtJUf3epWs9vKDM2iYjwIfESQ9JyF9Kp7N0IcjBtwnJk8
+ew6ORa8Q5cD7V7IYkNOD46nd+XJtx5qHFPZFtO4N/NzWLoJpWC4omYBzQCZ6Cs3
Bd5+fHZQiiPoUGGTjewrn5EKdFgZAcPFYYLPRK2fz1oG7f/9b3wxBbW/p7UXxWuk
nRmhnsXoiXcb6rwsXQo03rEl8COb2lXx34pMMbdaZE+OITrX/0CCInj7KPUwEqqr
qMgos4Axu71G1NmWAUqQVcqFB1Nud1k1Ty1JzWykn+8LyVIAGPzSCWYP2tk3uzbr
KGgt3W7m9o1zf1DGw9/U4+qRZnF1ZhvcoGf2Auw5lhmvmnbSNc7AeVuE2ZbKBQkY
P4fHiOuPIk1bpq4eUrIkZ350O2TJC7bkt5fQZV/SF9yfHAxm6msnNBE3MCkrhL7H
hKKLU4M15A/YW7kZCq6899NNoJ5PoZy7UuKMVTdFhNpjMNEfHVW7QSDY+gD9liww
zhshtjXg4sCvsXQ+d7pYioEv6j5ypBfolrqlON6Hz8yuJcOrhBtP/CexIvEyn6u4
oo4NrSBo6NE7vSBEnfkWeyXIkMlGLWWIcO1kWUB1T03r6kr+3Q9Ft+5dIl76F/1J
rS39RmhBkYQ/lbluw6AEQXQ2SFBmU5S1wfCB+Ya3Y3sFhaxNjT1v2TiUdozpfZVa
L2WGe9wEfDuQ0yPvwns97NAvt2frQEGSNMCAhKbauyGmj/6BDlyBUx/2o58nr1nr
HdslAoVMZlGvjc4SY4Q3i6bHDXv5UHqCVAG+L2Kfd0s=
`protect END_PROTECTED
