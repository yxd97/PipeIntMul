`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjyQI6G53rjtc1Ps+K5IO2+sZAVB7EjmrL3kG+7IMecDoiGdfFEvUIO7qOqQ/U+A
4tfLYtTlV69aGjd6+Ulngn+aEOLMYfiHcuMPJ8/VB4SOGkRMNsUFWOiz4dSmFEnl
arRi60OGyFRHwXFSrhnT88bwjubcW+Wcke3REqhgIY8U7MUqqYV4G9HPgJ+7OxJV
okbNAoJLzsv/DidFLkL793x8hBqgbMzApxZGQJPieBSSQnjBHgDipcWkYlA3uTA2
BDGlmmZFlKmpgQ5YTBG1tQBdwsjrUX903LjfOkcDcIzk6uJqTaRqjZW/Lsk/c/AV
CRdGxViLzbiOO5OOOxWmUrNRcgKMUrqYa/ZoY/OVBNdxy9jaSKYlrUcAGN81+Qa+
oe+6sEd4LF8HZ3KlrTWI69L/jCG9zTgGyFuYgYcRo3HT5atEZOzdO9ealh7GR7Ph
fKquujkJywhjqDQftqN2Pk0vaLq00QBTqp8eEm6bq/ds54NC6MxJ6wP531ZkVTNZ
niRubCnrSBYwocs+JxgVtPETirOe3Ip61+Uq2L0XdVUVBpHXS5e2uQdAKEMWsV2f
7XnEa5g80szqQaPagxJLGkT6YXmQJfzo4eOuBEQ9ibQICHGL83FnWwNDa84QGrAp
dfWBY5ivSJlttAgtCLA0r2HgJJEoD/5gxR5jJi2xEQEDjnweU8OBYyNtfCgV9Bm+
7VmwRPoSXP//U6n1gQFIkiLZvGAEQexen25efXHTgqLrENVx6yfnyWHioHvXjGr4
Ei7Cw/eZSyFJWzkRurKI+TJuSASz1INS6i5Nh7aGenyU3LlkyWRO5+mgWNPeTeAO
5uYTpxGeWYsvYvo6RcPUXd7Chew0kvodMt9oKCBtKTjaIe9OGjCZpZ2f1HO3sIt6
kGxsKKOBmrr3Abc5Z2NaHYDHgVjz4EROLrX43ddHfz1ZhQjdAnTwZ/AthqjzQoGI
tMO542ATywbfonzhJQCZQz8ApaFBcv1/zcW79UOH45u1OkBAeaVU/jJe6evPooJd
XddeVg4pBDcKqr/1wOuwXtp/M1dUJQeXnRtO5Dn/6yBVdTkMoqefcjOUsViOMMk/
62IngW8q2G+NbuM5yGLrwLvloEK0UaMnnHyNiNxJD0ilS+19d8N7eAA4Q0haNIKO
b16EFDnwzBCvXm37QZEmebkFbzoN40THsHkXQxF8sW2JAUh9b6h8AebjKQcHRepm
IgvXJaFFjKFZN0hhhgu5+wyYvlFX93b3sBYo0WhI672CEKtRUW2uERYR9MRNlqUT
JVWUeKbAJ4D73ZgcbnJo0vUeTu6EDetTDfiNY6JRGWNu9EuMAu0la+4WBpB5sDKW
QsOrkOWbN8RWc13LcFFsVEgw9htrcanJNG8R7vf6g7m6bfgiTQTtWsz5/m9+MDbq
DVKY2qae//Q5zcOIzusRP44Y0Oh4yAlplvLLGCWK/u0rRS2uGjPbv8fehBRvZcn4
80ObWXsPOWqQiXyUYeIbGrGEylYy9o7laV8b104HhGA6GKPbEVR3ayxYxKP8G8Ok
4QnoGv4wAl4WgJgW56/+hHLBxZspgNxRO65v0S/h8BIHdrQMkkV5wLxuN/RblhRX
ICdJKYJdhjX6itYRFn5nSYyrcJq23WQdRpzwSp2X3Je6CcQIl4CHJ/AfvY2vM1Ce
FI8jK/b8bbW4CdPUQmB+Wk5lO4cjgeBmDuUNNHFdztUZF+cXHITGKQQ251DoWTX4
+RS7PlJopx0jaf4GSs8OPjR01yXDq78txxMaB7tv9NgXhH8/DAFlC9d9NPTteLCi
PPQL6xg9QYGl/UAU64zSKtv41v0rj1EgLts3AINuTrFRB/XttcUU/Ide9lMrH589
7SzKSPyObB3RcKxogJ+g6I2MLLNedKlhwdVogQOTOm3p9qcz4+dkwrDU66aovNiY
SOSQ7f8pJu4p2ziI0b1Vzto86UHQoCL1UAuiBSabQmcPybcO3TVWk2tZvGXes1+B
xzqnEtS3ljnADoZpHR5ahr7ZGZJBSyvjFAxJjtHBba4NCj7WhKQyH13CFRQy/toE
WbYBBQm6chfjBW0WxfvfVHPUFPH8pomoklNjJLCrMuo=
`protect END_PROTECTED
