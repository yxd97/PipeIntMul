`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTTLYviyeE3wuY9D02DYmiWgXm/anTOr42SSYzM4Af2YdUkZlNvtkmXL3jQhQUvQ
a1gZRwZiiQeF8FX7Rh2el7k4nmx9/sK6+G1x3FedLtVe1jv7qry2Pwk1vY26RtY4
jqNfxL47gCEoKmaTAx5/fzBm73EvNmcjOxRnA7by1fxPGul2/3KN76ipuIljstvA
FSjjbdy6R6KRqif6KHUmnQkw5+F5KULcRRuGyCbNaGSktxjs1BXSiHpX/AD48J33
8Vx4kXwEY0XKtC+J+H0YLG5JASMayh+AY6uqXK6wpVDaHnAAqZKiDazRK2j6BgEC
hvhosBnAjLQU0cTnoYJY0fxOu6MEYEZcX+Yk1YkfjFd13FTh0h4+F/Q6d1L6LkjM
Q7xgTbbmjRHhn1JWFrFukjhsXn9iJyILChRAJGSKPeSUcp5J2QVY3Y7ts+HnhuoR
XDftvB9ePVWRmMjxO7S3HlXHQ0Ew5oJAA7moiLo87v/5wAT+moBheCeaSiPVnex6
9hiJYhrdQdSGOE0dhNKsNesVQtn4v91jKRAiW9oBNlSXJ4pVUe/FK0qeJD979N66
0P4Xamt1wQcIMrS85Ftl7LzAirgMjh4bLgsbV6msJhlPBiw8wNnPvN5CSRnaOKeH
RgiCxLVSPw4zEW+JXi70EKMgFo0EHFVO1S17uF6a1uqdCGZYu0K20lnvBHY/43eO
uJfBGdTu+vyocPwFx0n+uRaLFfVBiUn0+OqXxn/3FLJ7F9SA2bXQMsKRdoNnbE8O
aHAQkWTG5ztlvCNLDCMfdwm04ZrtyaDt81S9bwTGfG1vF5SY+xgYlZdUP670DV4z
lIpV3Fua7LdS8hhnIioEgSJTHlAmKQfWO31JrdQeLCxl/2LimH0oJ3ERKoxxw/OO
txZO0CiL1BJqlxffXEXC0HnPuJsPr4mhxZkCC2cHzPN8SCeLe4CGgpOqDC01qwo5
Qj8gTD56GxAaDwWBVe6NXhoccXQCynCb8G/PO8UZhqWXqd1NAQgSRi+EH8I8DzGK
f3lK7uiq7/6xEHb/tLbVNLqyKISY3dUlWv/NYcQYzHe8d+VG3G8T0mk0VxgDh86T
9l8YHUjWPE+AUI7AOyBOtgb3hiQZ9JG41EJWpu/tRgChkv8KJZlLgccxupPYqINI
`protect END_PROTECTED
