`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6X+rYHQopgNjw2eT/ihz9euy4kWLi6JAqZyOXiv1aLvy5gtys91K3sWgaCHLrENy
FYqQL1B8tBf4nAv+yiYaOSlRciMpW24lAdyigi1/FfVVqOjMIwwQDXiTugEA1UZu
5viO3uuXdvQ+lpO4BgQ1x5cUn4TQQz1maw7qcDWIjE1Dtb2evC2wuX57CkWkUR1K
PG1+kjU0jyKTBoZc3U+QoY9JNBh2gpNAdiJ/6TF6JLyADKkvezSOsyXPHQNpCzl3
qyUBbCLgYkoNJrP+ZbgVHhaS+Ty2ViUZWIdMj8EoGGy4zFGxDMg2ePff50fUdMPz
kQncXj9LTGCqGRvxu4xkFwrIHS3qpnbSlpgVVayAGDA/vY08RlnbQJx54tm9DFGL
`protect END_PROTECTED
