`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8CcNYC3E8qTHonPiYVJl0irpLlSNmE4pjcuTY6VjmYWYACGhUHWSl8DTR9rrN72Z
GPnK3pA2KkTvQUDZjKg3BpC/UsAYVxob+OpWNe4HPvD9a5rIhqhr4NhbPDM65k8z
YKmbbDzJhZZVgcLaQLRvt6gl4S+hp+2R1QgL/1pB7Rd+crUS3BBpXurZUwjUyyhN
tSCk6kLtVUyPoXdSLPybQ99mAVXHXeP3/1yyg+5M90JU5uluDHyFF2hqQ7ts2W+J
EZorhD4KhE2qRs5OC+FutRWJ6+fs+UdJv7M8FBh66MwxO0/mVHUd4p6bfu87T34h
FdX2ZLB1665CkZFPiaYuo0ppdEor/vQzAL3ByShgngizSFzvFjKaXR8G41b38AJ3
FyV/NplsFZklfxaVgZCivvWaYYqT5iw7PdG9F6a2zSSr1Z4ChJrNdmRyzWAsSWMh
Ut88avwRPjy/Tg/ktnc+RWktbJEygS1c7tZMVUMhK5sYHurQYusmtI3LQqgelmEj
w1zWAbkicXlEgwocgOUO//joQZJuRel+7nNYxDdcjLWIxtFL81535+Ff6BnEQdyp
5g5rFxMNg27hhZ1oBAC6bjBpkDBcWloyKVFhj0KHkrDgm5/62DNA5RF6wo5ZVTdm
B0nF4rE3sne/cFHe8qDnEw==
`protect END_PROTECTED
