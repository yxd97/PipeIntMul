`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DC60cNPAKmiXKHpp4aenJ2YOBFEZyCV5lESzK8nhWwSU7V1L7+hEMacD4y8VeShx
pLe2RfH+mvLIvdlSduxooANLDJ7++qlDbbFgRNyf47JsDn+LdCMYyB4glxc7e1gQ
mTeKKzdBn4YSypvVWqFh3ML1P6fCmi7DCU4wa2NfzUBWl3eT0tE8qiT9nJHQBBOT
vo6wyioLUWVea6k743FPxo6u5B8aqfn878xb+TuLWhI1k5AFLfj3DLhZHsv5NAcY
nHIhe8I1aX2z6L2NATFapC9bmuqdviLjce6UnJoEyA8r+T2bRf+BsdwTqwtWdM5P
rjrkvGflWMDsBmqzRblv3d8f0HBfqHg3IRUZiHySfBSzz0CGIgwrK6ILSpybt93h
4vRp/71cqk8jsGMOLR4KntY+RMtbTKuhn2w/YjQmnZb2hTdvGqujUmW2JJuKDW6y
nbBgAAW/lLImjRvJTJ0s/r7Zgp+KKtc0vasZ91Uiu/ybRqf+d/lRa61MVID8Kivw
q7d25W0Fr4HVj03mtnknn5m1PLAtR02guIZRPNQj3DjMkj1lPZiQFe+va+Er/+tK
p9TPAdjfchKlkMntmWUic77t+GAOBQOsyUV2lPjIBL1vBbedH/F+2b2FcA85Iiht
`protect END_PROTECTED
