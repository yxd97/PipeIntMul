`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N5k1T028ul0leMAYMRYHaVZC3PVoJxI2z4GKzbNTmJEggQNRIp5CnQ5qiKNjieI8
JviV/yjoPFECXwaH3gy5hv5SGjAZtkSz0X0U2P76tx8ihWJWkFYNr6rT0lfnMRkv
/H8jqTpn17bUw16Z9atadGahMscqqQFLAy48w12e9YomvRIv1wZ3UmoSg2fcvOAH
Y7+myk7k6NcT52nQyRB2pknsCRDen98MEmmnzEaws/Y7CMPFUnTt4XGf4FwYpyJz
thXY6Eb/EnyNUC29czR+SQ6I4/E/AnkpqyJh8e+YxX5JO5VCR55hSnXRanpTmknl
Adym1t3IcIWqWMwHOHzhYbHHNW9Kd2g4KkpBJC9mVHA=
`protect END_PROTECTED
