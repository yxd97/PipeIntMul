`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npdLTfDl6mvEwfbbfApWCdhGnS1fD++FhG/AUgNUTuLiJgN6FS7dH4ecNmtcZqfy
J2ck6niR6G6PfUaHgUY/8D0/YFEKn66+t6DVN/YfSbniyCZPZZuwozG5EAp1idvt
aHL/7ge1PHs4kmYleTc43LFW9Ntwj4jABHFTkizNL1bJr+BpU5hdASSUARdJrAA4
L1H5t7chd2LZZB+xuG0OK8/vExNX3F3C5RaJkCT+LUXNlhyjtUfMxMNTwBQg6n2+
y54HlIQTkCjBRRO22u9f2EBB6SdRdUBdiIKnPPxx6ZyNtjyuakkpIf5uOrZB5EKq
meqdcPIu5yaqeGIA6AS9X5OVDon7WVeZg1+QPo//lLmPZdAqI0X3rurGcNTdY/Rl
L8OksE+YRo4A7tPPmQUw7y6PkD6+cOmOLCyj8EsAlXP2JiU11BQWWwKuFUjNkXUN
zf0qANum9LdbDW9EJO6jLlR7lzrj8pI5fFaE6kzCt5jpoefEWTHMHMIyp+2ArLVR
8ZXBjCkQ8TRRhW3lFloibG0mttkiB0j44aD9fqZtTU0qCY2p9IvVAPkPHislCwq7
gpFfxgA7G1FnTCdVup1iyMH7Zwikpc0yPlEIOhA01lyQnb1R6iD2Oo63/b1Mluow
Ne0xHaFXqrWn4oWMIsTjYAxO7OEkV4XKFs65oh/Pyvhojrv+GPhsTsR+YYyVCdNz
A89yL+b6eJoeT+IJUUUsBihMvYHyZaFgM/Al2uaRHAdQi4FCbuTtiQWt5L8xC82X
Q4eBk3jr17lpR87Op9/jeQk/L6E7G9bx4nyifft5smcIuRdvPMJAtF07F9dpzb1d
QZ1fYbQurYq42R4AcVMdd8cpQ61HybUAQD+Ep8EHlURFq4CWRwY27AIb727H43KI
jgL2wwh5K6317JPe8WE+YRUyQsFegnB5oFZDswPOU40=
`protect END_PROTECTED
