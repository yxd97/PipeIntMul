`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZaQ6s7aTzxYZI8kzP6hAqvRi+ktc2EJ8ChYTWafe/h5F2HcqTal2YiR7LAMgBaB
roKmUmIWs5qdyMcNGOvfmGNsegPz+0hKDMRGuoQFK5rj8OQjAkI62WauTcdd67uK
DX20h2QIrbzh+/4/O4Pfjtap08btDzy6AtWVXswt3KjTnCEN3DVEsfQnV52QmHb4
WcMHYqGF4bO0LzivOZwrpJCZAW2UL8VmJuwXYD6lmSLtmu8VZReCkUxSVpJvjT0p
mt1vRYNFpNbUV3/FTYrWxxygC3Dd3A6aX7YAeivBGKyAPlx5Ljk+rZrSuOWw3EZ6
x9kqw4qrA0mBRsO4NhUWGRxqrkNTcyvUpEsud0ptjNvLtu8m2lRZrgnOtx08TBrH
FoJQkzu0LVXF/RRlgnst5lMLE9+4sUkELY2dvMNMhh2zdWbFtMDWq91LCBYDtvLg
07bu3NG0051nbjgIzhnwhLM5KRoSVBHEOMU9MN51R61HV93UpYM4LPxrMWRkKTh1
76LjSK8kkyy09iuPbV6KWD39tOhvML+f/4RmgJfmyxGtgcTQXaieWWYTz2nYnvm+
7w2NdGbJVeeG8lGgbyf+jBGD8Fk/vYXXQHht+F0WP2YoNPC/xj5LN+dblnV/v3Z2
cfGB9QdHsS7Im/jN1ifhjRFKgXVGECG1lm1yyYfVvI/Ti4VkHlRpuHkiQTm5bdX5
ER1P69G1Mo6vitZx/Vt75T/szJSC7O1+ijuKthmRf4E=
`protect END_PROTECTED
