`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gj6WHj+B8pd3TzxHc8UHEDPj4XLNtpUiIknR2kcnhPAqeF5IpUo5fAL/9tPGNGXK
EAzKPIH6TDSUKJgGx2YqDGVDQwGlKR5lVt96hPn8UEXcMxnRR4o0SzckOxF31oTy
DO8G2mnpBsvHDwiA8ftCeFq0//2AKBc5oVrS/sITtvqAK1sIMnV4FGAhsDV7/r0K
ZzyDWAPGBoydRItiAFcrS1QztPf13NZk4cwmmRzuF8YvL5mSSk43ckKo30JbpAu/
CjYPEiJVw7hSIwAyRCwBZ2U+Jef7QiY+F9W7TMrbk0o4uTe4qy0Ots0P+BoLFBig
+xPwEAQArPtLj5hVUTMcFtFoKQ2a2N4cUj6VtjrLA+axzig/FjK3kC4Y8gHRx8s9
TB8UdND9eSHAONnxj6vAYJuxGDvuid1vLJx6ho/goNPESV6uA9uWtHy3KZmFt2N9
C2nTnH014Ev1hKAB5MIP/2BczBE3iuw3AsTw/HAKptHojnaFduZN2V945lTs7UPX
bhg9wOKcUE/UwsF+vuroy/vPg+CgMh6ayXurUAGvlbQ=
`protect END_PROTECTED
