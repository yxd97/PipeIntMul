`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KSTjxoJ9M30OQKnyOpy78wo9ejkD58GjuzYzm4M+I+IROhBDClakRcBvbP9+R80Y
w7oZ0QHd+jFq2PmNIj5M/sQ6IkWpv4bIFcR5nJg0vgoiQkklAmHXZNCZMxoz3vXS
q2+9kqGd1b1yU0VhCDJX97U7OeqbBAtSHOuCPqRclAGeobdCp5uWxARqE0rfhFxq
Qpky487K9nDZUOShBIMw2N4lz1KHTvgSJ4TzWjN2heNG0TB2f7BfPjD7i4va6Gxd
S+mf+rsJKu0woYR/4LtmfEptzDBU0StzvTiJ8mWyqyCmsRgkuyErnEl6TPuQWWHn
afE2nz+PJ3zT4shwU8wu46SIPkWOQ+N6TaKPDsGWDS8HnrCTABII92NCg9GYmLdP
yaybI4+h477lhB6z/4O5thFtk7X6mdgYI0LZb/eYV7+5UgP7u4QF51iQC5vUu8bg
fwEmMFiDWz/XCv1QtwXms2eAO7Y7MNqkTTCQY1Hu80A=
`protect END_PROTECTED
