`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9W/prxHMXXURbqzS5exARoUDzNnPi+u+NU7hbd/yxiCBkGfgafPAcgb/Ley8179C
FySW+2u9bx+iqfb8wqi6dnVJh06sh/JHD+ONvkuAeIxEW/sdmIXiepxap8ZooFmX
JDE6AET0GwgD39nfXGn8HChQiTAVd7XYA6RgVxg+HPxhLBeVyIWzCEUSHwN13IVJ
Q3sQSVXNNuxQBzy0ix6HhHD1dYCFiLhp+AAhDnQsTxF4F+nV/WMFZ52Pdj153SKP
r/018WZOCPdsy228h4a9r2jQtlbLKH5NlogunnmCalPxm2UB2Vibvr5++iCib9BH
/wUFwUfTvP2sA/M27KQ+L4DTOroHqb5oCi1fut2xPymPzkZKeDvpndUocGQUYrRC
Jfb0NClukW9+G/nqgJZT3Te2LNZ/YFb8TedpVRW/sFS2alCtJI3xZK7uXJ/BLIRM
aBdaV6xtfhbtekxn6nA/7davLY43tyMmN8hDcCnj5EAvnVD1ii4fwXxq4h5o09h5
By60LqfmOQKg5Leg8jmjiuYOhHFTJoWvgi8f9WTHJ5BEutxNxKdU7lpwkF7rmBBz
OesXAG99l+2FTRS4d2sGHF+S4zDKDf7qOriVetHgOZUQ6pk+PCRRO5mOnZ36rbzc
gT3m9aXpxPsH8jdlfeBWbBqEbRdj4skCqZrTVCFwKUczyrMWFfgLp/oXmvHnLjwO
ccCPu+RsR7tybph57kk3TuVhdgJmD+2oyJigRT5Ce/KJH1WMWAjS/oMYTg8UY+wJ
d99kKLJjWSnK1+CkWcwA3g==
`protect END_PROTECTED
