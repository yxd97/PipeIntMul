`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qbS8ug7ezmm9FY4yjiCcmXwnKp5zIz18aX2xmchR6lbPE4rKpQ8ynP2Om0ULUa3m
gBrFdarosn+hxXKKm0zs95KTtO2GWoWM+3Ema7oypoAXC2cmzY4s0DohDhCgBt6O
qP+CqhuNMxyCENmryBxQE2XklRU7ejNUoIlOXDOBU8/r8ce/2jpnUvgSH12X5c0k
FrZZ35J15tjvRlndBYqw8rPd/JDeQUf49WFnNoNL/YGEexrq3LDg4/1qZGjO1vo2
84Gu+wLHu7BRrwI55tZ+CHZ59PH83/e+KIxi5+BL5TVuz5ltewVcdoVPlvqLJIQt
z40Da12nhmqsoD2AbrhKjhqyy2r2+KcHWA3DQ+qYLA2qm5WjNjb4MXy2dHLGbz8V
rsJi+MkOg1NN/3O2D7AFMl4lPfEOt6lKhZlkzOuY3O1dxGRlxf5gNiT4iD0nZPen
z4o7ID2TZFmEo8fCTKxcWp65aViwUsOUJ2VZYo2nB/AjlSrrTRzP40vzWQbEmgT+
P48C68rVeTCLw7YNYw0b5qc59XSw/7ZaJidEeXFrc2ZzcKrEhFM6U8RZoeLN8ZJT
LPraSscsJKdESk4iPP41yde/nqfspct58TqyNH8hYX8Z6roaZPHWl4Dsx92Wf7oe
kqkjY3QG6JIOEmtKMauaqA==
`protect END_PROTECTED
