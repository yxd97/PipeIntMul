`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CfQAsr9CFByvKUHwYZ9+MTYLvN9oTRnCl44ng/1varDGn/y+3opOteOIikNcxq5e
JL5rwIVtNGX5HSI+PmWqL6KOHrhPVaCNbl4m7cOD/oJsIuT53aNErU8/+y+Hsa0R
T4HdyCjOOVp4yq/gQW3IAKSyvQtkGeClr9JE6BIcj3uDrq3KTinKYFOEbuKLxsZN
yS1PUVfIBIj88e74mzfS+hv/cTaXc4gvdXt/ppeWCAqHpXuF+0KKAhi14Sfk1GGa
i6jz47aMj+tKKlQW1E71RO+dSPje/6Ui95lhfjYrcOPzu9pWCaeon8CqUhJX+987
9KMFR4ZwKSBMLB4qwh9ERxBd6JV7iKCX7HGSFUlzLRK9TzXpUIWsv/dkknKPQjWV
6io4gpYJnpqIMbNe8SCO5o+YtuUgKCIU6ZDPhkj2YA8gUqubZPBeIuJNP0JNeyV8
bjvDRiMphlGfb2jzq0BzvM+dN5OVHJxdtnPAzjs1DXRPU5cxGNuP14ngsQKJHPIP
5sQPkcus4q6tuOkx1P71inLT3ymHdtpp/2x0JAf+SIqcErEQsU+B5cbw+c0OGBac
9IGqunVa7CzG7aq09QjeSkdiISjpfEpwAAsGMqo9/aCNtBBGZSZA+NMkmLWXY1yu
34m7KOCL29FEGghj9J6M9nkiC5I8ua1piiyZdigDiL/bxKJQHJSmuo3quC9Ptk8j
tdK3fzJ4rP2q+mXdNBPousHZNije8mqewUqzd4DgzTeAn4UbGqaF/LfcaSOG0wOQ
BtqP54fDULmv1wE2whk+s24NQzV3a6HgSlESeH1+iH5jzLSRKR7ifNa5M6gcg/Vw
16x8OEHk5qZmwZtkba9sWg5PRx4HHORJxfnMiPTmJv/B/pzbP/hX2WKu+8hAWZHm
GTitBACN4JNN/IXUP2k80Kfhn9Ncy44Q5wWQGIkocnIM0/5RWZfk7HVfgetMnJNb
zi2t9b9PolYfZ3+Z+P8QMvkz9sOTk7kDgJcniC1UMMRMKHgPz15VO1STeYg+4lEh
MfAiyYE7Df0sqSy6rtl4Mf5IDTBld9oiukzCY+hR8jtIbXCw8O0LJhijGa1NqO5J
m2zrvRiMCLqhTRKCBGRElYWEv+EffaNjcZ8KZddgGi1eXfigk749djX4oRo8fGxV
X6VGZe8v1VvymgZKhOAMl3R4uZ3g1eksIOigZ7mSmli0YIksNpO24ZTReFiWlTJT
9WU4PL47MJmKHZo/lnthI30YAvw6nE4t6k1O/wZ2GtWLND+8AL/1l8iq79GsBIVk
JpGBMLb/BrrpW0TS+chSQW7R9uJCw4+BJvfddsABnhmT+G23iLzfjJMJsu82ttOm
onwtmnTjwJ7g9CvXwHKwMg2MsmBI436aSyW28GqPxiCrHJvhe1Id4147A34eQBr4
FzhMz1x6Ggy9Cig0iIRv8iDeek6jpMufz71fijdeaWfjMuI4YsxGzNjXbU6URaLc
ZLu/BsnIJLquzVvoFarFuizYCiYPFY/76qKaIGCpvpn1SamFw9rKRsg/oItyXCJs
esiuAuI76/WEEcKPm62QlDCHHrdbjOGWoWW7EOSDzb+LhxC2sm6AyFmDLLq+3bwG
70xcQLk82KwjgeKxgKtIPmyuSx0teLQLUOUH+mq5PxZifxtZD6F6MkAmcyfY2HM3
tUxA1KijokZFncr1PiGHZzkntOXgpLDRAVAsSEV3PvOjzRmCiWhsrS3GbSQVBHQz
yU35BBMeqHeG+n7pzw/VgWpexii9JWgRmTZcFVTojjPqpl9QFyDErTFPuerJkgi3
eenMka37gIjDKnldnCRmR+oxtPTt6jIf/xvvF+mEdY7UG88XavHDaslqnO5d3I9N
ODXbxbUmfqHKZx5L+/2MbGhX6kIQqBlZRWL9MSz8orbrGEYmBokinHqzOYBBt4Ko
M4woh+cMrQybPMSdgPKlqxQBuBeXx2ywSarxbS/59kWL9/Hr8WTI5ZhpFKTnm5Nw
PBRuLnBqc2OFqVOH8erk4wOU/4YszJInwUhXdH/nTBBdLBqpD6MVt+bTyU8vaDHH
p+dVt5R+qLkmpDGbUXKozfJRX2+oFuLDAbQTabrkP5mb106YcV82WqCGk0ovZ4U7
g+y78pEVRONFK7/KJebh/6jJ8WOVX0JdA9t+lXfznjOCZsE7zgpVu83rlk9mH88c
ugmr40LWIhSQ79lzuzQ0lS3n8pZ9ve4QkjRsTOglpFVH+QjZPUV8rX5BYas0RVZa
zynb7ZnupcWKHSaxn8q08cnYJz9KKF4Mq43QXDcSBLTjXRAxqmpY2+Ek0kQAiYTF
rZit6tF6qzvHhy0/unJGIbpJRECNYF4ZCkVzJc3sm6Quiym5WX6cOi+xtU+gzRpq
SK7BKGpxv5d8m9prfgt9ElPFxi0YzQ/ka1StDVt81bTSQk+S07m39wicvEdVucZ3
ENRKDLvqSSFrYXSWMUhFPDFpL4b+ni34HiMZ+JZR1DupEdn5SB2RBgVB+mmYYRQu
L4ysyfKARUiZzECcSi9XSww/DJl0VNoRSN9N3K4ftT5QuOXQsZkGHCZHK3+21uUp
+f5ce/cgtYCDs5GHaRiMuk5yGZpMtKkMip6QoLaVZC0KMgwxLKJJJPDN9IQrwDRw
8fZE6wlCyZDtNNn/jRwm8Hn+5tc9tDPIqchp5kkOKRD7y8eNDoMiboMDz2zSYO7Z
EbNpaTH7sUBOrv/zh28wUtc0Fi89YxMZSPiNsBiyhGRVLmkVou0SdwysuiVBlzkY
mwL4Qpc72LceEjJAKdR24msMC6PqJjMC99Gu3xXzkYKmYbiqny+HmyyKa3gXEQhF
vOLQJPt8YX/RWV86Dzl/X4/oiSx93vgvNLtwCwYH1mc=
`protect END_PROTECTED
