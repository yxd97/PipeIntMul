`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rryZ0GS0m51PByUdIvG7KFdoBn5xAC30jAVpeQWhNdxX9TuADVbJ4uru+1/nScAY
XKTaigcrBF7B6D3S6/GlIMXaLDrNvKj1dkNXt5can0F4rvrWFbUcVfghTjbZ2p4r
UGgihvI79U5PUW7UVlWqgCjblsYkMBXBpF40sv3AU08HUohO9DUgqFa1yxPmGSyy
c0KF/SKzce/lEpbhEieCfVKCHLYzoDsKB78lNLOn+jvheY31tLyx4PrnOrgN5IH3
UjOVmWIzwVxdVT55STyUb39DziFdyFpyWHAoiv8+d09yUmCR/GXi4A6M09lLKMZx
Ymaem1LV9kEV1RQAp/HyypAa77ruZ/fI6dYHs6TOiMD2+2jqVU/dZ82ykkHviioW
ZnJSHf1G2Umw7asU1En+DYO/27dBU/I0h46J4ynIJpELfqRTXhwzOYkYw2P5VwDC
llAcxEjhUKCN/XByAJyBxrJtKnIPMeSSqnCwQLRVAe59FbORp/edUv179xsG6DC3
WrTSvjnMt2MVMOquuFXEJ4MDd/oeGep4hIfMeVLQZeJUOvj5Wq/opAZKW0AYHKKL
LN16/+8EuSH5e/vTSf4CTI1guuQkcwbHDLSkpd0IvDNT2NP+ofuAXI4yupG0hjmf
7QdEFLpiGA4ifR60TLP1tLQHzVs2+/Zm2/gGXI2i/xuKBW+gKrC0ORxi8HDF2AFX
U0mxVndhBlpw3e6tkp8alFp/9KyKmU4sf2MFPiwv8ueLuXD5+YsXlKgtEGmVoM4h
s0U7r/VZuilbb9cT79AFQw==
`protect END_PROTECTED
