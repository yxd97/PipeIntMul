`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+OVV+KbK4knvL3PNMB2GOOmRD4NcUkqLYrVXMdaJUid7p/E1U0ntAS8Vpx1QRX1A
xf4hT6KQWTU8BjBpvNTRHaZ6ulX1zxV79cULCel+9Sw3G/yDBqAr0d0QNWzP1Gz6
/Fey4PWt3Gw1wQ6jvcROHY6Z5zmo+T46rIQ4D3ZfGCH/b1dCf/54Hv36A6LfxW/g
wm1wNJVgGrYRIqgDwm04M8XUwHxHwHR/LRV5pNb6o/4Ybf3XV+vJi+2pVhBhgoCt
wDnVrLFwd3/7BbJCqo0vloJddUFbN6P5BbetibCLdzAffxB1END3yicUFaXufxw7
7Fl7HZFS8IYzwQzwKalq2jWrh52dEeZJstMtBJ5/K4lp4S0VIw7CcalX4yTenjqr
PslOtwW3DrxcR8Jhhze42OWzt91IPeSe3QoQvg3dICXZTIVdoetGuIBWz+dQnlTo
KH//TurYahQ7wB2k7eKkVNLesta7ku/BnLN1Qa8ieIk=
`protect END_PROTECTED
