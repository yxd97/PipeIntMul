`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bFnZ/u8XZQJX314WJKHVmP1PtRAV7a54eQkoHdVPwXaTL+hPjoMdc4swevDZkGf8
99b9Gi5/4d6Cn7Tf34vlgX+5Zcx6BJrByN16xfEm6pMeK7s0GcMRE9At6KnoZc/7
iAjCRKv2lSnownKZyez9R0kcYGtrMx4crj+E5qaYftQubwejrXOBD/sVI3G8lOCn
SDLwP00oeL6UYcnw0PWjPuc7Gq8M/G+QqwbXj5NdQhk4d0s3OnHRsbGyqYzDF7sS
7Unt/wcRi3DdFpIXPPjD36I9QvxaFGw3EFJ6A7D15dNIyOLmXPNoMoBy02VerhcU
SiYtInx1RT17n7f7sGNam3vhU1JtfC6mM7uOF7jgGZVeEZXJuWXlPjSWF0en2ylm
cv+eO+zKZZaNHhKiRXZM6Z9XOX4nrrIkH19U/Bf5gFIV9uPMcrg3sbTXivq2taCa
w0gm/VgZvUUjP92M18ODuHejlfbn2Br7XENBjp0a1Es=
`protect END_PROTECTED
