`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCL5ljCmIHWmnXSswB6jn1j4IcpVpVzMHhvm4bGweUJbIGjMT1oBU4hYQxTotyVd
9tkCigOLKXeEnfw4/WK7M8EwYF0VYqilALebXtdR5FMJgBSJerRoBTIy+pB689eI
wcV02+B7tcA0ItgWEBcLtDS9N+8WPqrqvbEAt8eAQN0IoOIr6bgibzPgXxwmXWA0
QSDcsH2VYUP1P23SWVKGoyWXHJDsUwCKOA5VuNnv41tYmcNH7Mizx7pEFI3nW8W8
W3EaiIkgyU43xx3zxmlmuDHIBUrfOEmJVBm4aMavyCZ5xNpJEcX2BHtF8/n5w7Nq
b2AqmaWaSnk7TqN6bA0AXbM2GSd/M683QCMxbINo+ojjZdx+Ha2frcONMeJhxu6M
BO/NF7qQU7t7GZO0wpHYMmtm0hRPd1e7CpPtym5qaWUkeGGCz0fkZ87RidbOLKeQ
3vUNfkqL+Th1M+vezeti8UNCIBAQpmYv5z5WKJm9i9eS7IUxhZguLiz0nifby/yO
8lfDA6g8h0Ncovnc0nlrlhoBi6jRBJeGg4YJleQV337u3B9jAM9fDN5HU3fxgQKt
6YQr39iwwLpgHvhLzVX+lIXIgOO5XKZHr18LzMPfyiczzNKq1mvIDJIwpVrL+0ER
Fr+6sF8R75GztNH1pSNTR+0Z10JfR7Z+J4kTOyDtwPnUAMmxYLCmb46n06yNQp95
NA15BdtnNnM+0nsdmRSHnsXArIwRx2D1DTpb7cXmiWI=
`protect END_PROTECTED
