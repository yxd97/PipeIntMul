`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frb4gOHzECoG50GTu3/4LBSKwpT+duCAfwSf4JyE5/8inCtdD+UV2foH+GM4hwHB
ob6+gjHQDrdyoSPxFoG1M5hdEMgy+rFenPldPzSp8md7j2gqL5KICVrj8+go1v/m
YHMWtcOQYZYNCzc7NL40g3Kot0Df+t5ZPMKtP0FQsXzgsTH+Kz+hf6Uwu8+NWUg+
Kh9b9yBFAJIj4G2dpbjFXMvD2M6mpnNziBp4VhEsNpfFO31xE4YjXbifwAxNMfXN
9w2D69zUIX0RTegVkSzev8ZG308lZvptek+u+JF0xKUrg/yqMx29E++VN0yNEfO8
rlRguT6etRgPuSE0e1rnBPDRXLuy0cZYcypmLO4OxXmstpMXLNSVPgqZ3kdX6tS6
`protect END_PROTECTED
