`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cd6hOTgU9LXlHeM84WgEeTfKHGP4v3RRiTcm6MlrvRv2YvzevgvK8xZGSKCQNmLC
0RqSKU4g+PrR7hgveirCmMt/rRXATkTdHasrprCFYhj0M/IAV54puZ+3u3AxP8QP
oCi2kVpFhKuZYFAdHEDHgzTZtMqWc4pQluGzoM1GqBa7dxgZCDa3MfFGiUR5BFaO
Q7bBxJ4fs13fLknfup3/xVuXqTA9or2bYdr1NCiGnsxPPw6fxe9HOQTN7UZJyz3Z
PIqy87T5wVC+7G1D6+cw3TmJCSt7avuDb5nYcL5BCRtJjAvKBOhzkbUqLngIBAPb
4dQ+8WpM2lx+Aihy0htD8ugG8DRK8r149LoQl1e2Kilm6v20e+2wCUn/p07yDZL3
APuLnZg4SZUNS/4nwUMGP5+Tt9maez8fya+daF7/++bfvyQx2GDetyLf2DvSqHTu
2wLjkqio22y1GF8r5V9xT2NwTm8m8y1B+8r7X/FMW0a+4NRxj/zC2zXW0hG7N7Wl
m5SGn0mu7GbQxfrNjgvZY4yWwpVpbTJarfgFt0nn8uO6I1tc2PdVa+trVz5oG91o
`protect END_PROTECTED
