`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0g/PkjbrIJuQDoFZ4HweSGpwyez8f10FDbTOLP/YbM2UH4FS1QZRZPSxXvLqGp/
LOEpVIKUIEj070YXwlZKVTRRKKnXHzSaAYZ+5tLSZvPAteVY2KAuUVbhzHvmgFZx
RnWoW21PWvK7pAhvDdQVK827wAuU5IH0HwIDC6NfpaJvSUfBawYoLFqBMntH9F7Z
BdE7kaeFr1p2JwxQmLM+RnEHvpcbkX1nwlHQKldf28tyN6WBZ2UwlgHuyBmkI39N
m1prYBqH6vyItAM6oRAVSveAss47Phx+X2n6eoROupYtnQOuuHXuALkxkTxHu0pt
eMsRYi7llpUOfDyMSaWS764izDj10MEQOlqbj5Up7lCes9Z9X/5BBo1XE1q4Zg92
NUhXeXTXa8KhZL9LcJ9O1sRpjasnxqrYxl+wp3tZ4dI=
`protect END_PROTECTED
