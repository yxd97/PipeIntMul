`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMpht+0zRUFvxj4MsXiOl8KUb+Y2txJQwyMaZh2yNhflO2+821KWuPefeBhG3fjf
rwDfIYc97inirJZDAY2lmL83DE34paO0oV2wLqFWV/FcdyBEj1OuyfKTLeCzq5Y5
EQFpreXLJXThZgbHb2jJuFe6noiqa2J0OtijKpmwrEaJjF2hkos3qZQFK2rYm6DG
MyBq+Yt+KJW/QrM+wAVcv32fXtT4RGuGVliKXRRvZu6pni5Vhk0txt89FwXDkw6p
AdOadSpfSr5gOt5Bkm6OOC29W8naR1L7aNyoPNik23trm1ZlZxjoNMaCMB/Lq0Ho
jHoJ+JLgb/uW2TWaT0KYw36NGR2mmGYXl+LQs9IWLI2iD2X63nJP0vC+UBXY5TLS
eyeTYnjjTlKvuR9YX4aWQeZuoDIPdCwiqwpGSWJrwJ3RC3C2hGvBEZL1Yc7Ygb8R
vwrfI2TJsjVt5xurR3Bk+2aTjRQFtU0N2+XWlx+XVDp4Eq0Lhp0crbPPaKvyTabh
YRoPvh1mgJs8/GbgnVk29yOPdPEb5MPgnywKbYv+X1KDHlzqHmN7BaNz25R2XsYe
/W8Off4U7gSswvRS0x6W+qg6UcPWnxO6gQH/jqRmqTe5iLqYxCD/GVWSPDp1T3LW
khmIrJzv5FbLkbIWA8nS0Ij+zdJO/kqfT3WJHatVHh2JVR1DeyL2wEhUk0bsYhkx
52GUeEPe8OxxZB5B656brw34SHPWemCQTU910s9zxyajQWIuhtavebGgG53u9H5H
b6Q/cWtN7NG3qCL+HE5Wbdr3eFkyuLZOHZxNwBxf+8b4kHg/VhfZe2jjKqeW6vWV
oWL1QxV4RoZgg+xIq/SbnRghfxyS5lc7LOhQhgYJeW3N0xcFV3PgajG3H5eD/aNU
FwS2KiMxFKgEn15cDczEGTH/y55m48SrVcC+uTAFGxz60wtuN3ZfoV5QTpgTA7KQ
4hg3aylr9FOAxEDmWlcsk8c38kKToTfkFoeDdlKaA/TaYtcBgNVhf2fp9qmRUdmM
VXyjrTF+agshUoF0uSoacVv7t7r8ugbgiL+P1Jr3hJ0EEAgVogoq88gTFup9x0FD
zfw7H2omNq1j3j4E/sPIsDo10HWjIW2krC2+klJ0AE7mNNO4u1fMfxsK5wnWueGu
whew8jzNyn7T2d5q99E9HNgT0+YQjUQLsRFVwGcF7l5ZRo6XTY15BwqUXEExynha
02vwwf/YoVl7yW+s+AtTwEtId0EHb0Y3JiOqGMOLyVIcXK8Cew+PP9NsAIfcu4XJ
5NHKADTFK6JnEThP7vb7gNsvOjmMRjlm67bS9dVZmSYufk8GCZXXDh3NisBbXn6W
rKNzHVaf9bZaVW/FPYoR5WtSx5kqphneIWEq/OtYiUuNYES/p0Hyum+N0bcrdKrT
+vD9nPHPEb7e8HdcnEWsrMT1v9LxMO2A9KkL1dRCeDNS079pIyYyX+7Jt7e1I6Yq
3UUO681wKQ45Vz+7/UiOtSgz4VUkPRK5ulfMoAE3cywttl2lWu47sVn8yHpwtjsI
tL0Gv5PAbM14Gq7EQNeoTOnAJQ16SwViT3MaWzG8chd44Jd4Ee7wiYknownvm0aB
qk0fC9axr7+LeJAkAfRvn4ceX2MpslGwT2Q8QPNC6+2Bs4Jww0GKJZQWjmqjC6Cw
SBLUGFfjGplkGI9j/lno/tIvUCpVgou0Y/R8T1wrbl1ECu5WQXGxobyT2bb63HXc
DZqRcNySdYfMGnwmgjT2BUCtkWThhnKohmRpMAXKzFycJZ6IoHEq9zuRRReYbwoS
CVrLk+yZ2aGc4eJLKSXiCjdHiB1M5mJLSrHRfoFLQOT3lfL9Vg43P1fEodUuH9gR
SHCDn6183agLlyo24DFW56xs42EBPDvDTLoQUBsmMf0jwAQUg/ULnPofvkXkaHnP
d8NFyBGydFdJInYyF0yh0blyRh+L5U0+0hlE1bDim8eEg10WOzMUwNkFA9KQp+3S
oCJVqf/LrO/G61UynrcC7gQDE3xdFmGsSHuQ9nBja4pyHuB5HVfZhN65m9buhGyJ
Vyr6PlrhNrAlFWwI6XEWy7PlCa33gy5OJ9YEmvO1/azEI8cQfXmjFzpueKl1jED5
YrYK3NsQO2h8/amG7e4VXDvFJs5kmKYEdFobg107NfBRZOWbdf/ffu+3l4PrCj5q
7n4lC4AHFpO7uGOZ8bwOIee7rYSm4nEwyD0P6HtFb4p+J2/MNp109G/LnjwxyIe6
za1FEBk/CAyatKQnurbQnbnKu1wjNDgaSCqaVBZOj48Tac/PoDAxLrlQR+tQMLj0
3Ww/b8WTRpF5Iw7uEmoasQ1ocAjDQp43XhlS9nQDlLZrXtPTIfGEOnEPCQzEW57A
fqB4nTi/b2JaXFdhEXDJDRmroGEFJmjPX+9T2CoaE5Rw9h/cPr1zX7DCSe85rmsQ
5X+BK/TOD8QsjnCUMbu7j4j1WJAbcVas48xNjHWLJVFrgJhuAgEC05OoUecO7tqP
BS/xyXFo6BnpFJBfMAHEOb2sQgjc1dow7m5Fk8srmQRPwwxLGx1Pj5g+QpSbLuGe
158a7jW3Y5TLX2MuHHO1T6DmGF0eSvsqRN09wRyqyVykAcuQjo0jjkC5+V9Q9LXe
9yYg5k1MxwQHu6AmIlBD2bWAfmeVV4LrDvlvVwAJWcjjsrV+5uIqunet+M2ZuTjD
3z0awTVMW8aZn79BquIBDlhrMSDEmxEg9Ml6v+J9bnXkma3gLyT7NtaJnmpQOnT+
dPEUKKbLI6WnCIYjXWZ9FqiExQXKfz4BzJ/cilH+gG60l3RecZFMutkW5esSShTu
prJZz2y2UAVyDTPFVkgEvvw8epjpXTNkDCAUcfwkS8KyQosRLLs0dwgA/Xm9LXIS
CgLFVT/sg9TJnvlW2xq0gyIJalt7oTokyAESHBH977ZesBzA34NqOZEanVzrUPyb
fcV8FWCtQ/xr9GF3FiirjV5J76t9FlDvH0HyBCA0pI24bdz0xakfShLMp8m3yRVN
0GQxteYYGhaZBt3DIgPoqow1xyYO6Q1Qngergp2VFeAZHh6OW67wDqYm/delzjVa
6DZ/DvLl3WYbMiNE79J3aspn+Aw41+yIk1E3C9YxkTaOxWZSAloCHgQUHjga51R/
cD6W+854Ew6Ktp2T7J5no9xO0nRojoivX1CI1822d8mTf3rTnE7YR9bd7BdmN0Vq
CicVYnScN3UHUWeaCWoAqvJXnflCqRVYwTffjGlqO6tzaZD/ggdYq5Un+6JL7KnT
EEbHLBxALBt5Oxz33+8x0eQoG0Gy/qSqA9cw4hUURqHC/r24l9Awqo9u44j1i+AR
t35qA+KgBZ5loyx5UfbfKOZMOCXeGNXMsKe+evEzfvZo6zoxrioCQmAy33RCVdzT
RiXwCX+jc5rUGH6unLo8ZCQMgIhe5X3r+s2G9mG4iKC2WZtLdFnux+mVNPZLIrFR
QyL0Hp0oU9H9s32gUfNHW64VdKI6SDsQrIqYsRm9KJ2AqPQfDF3Lsp6U0xXDFCTG
k+4HUEslz3CEcc8fFmTZc9SwTZJcQ4MEqHTcDuRNf+Zpb+PHghzesafhjfx2cie3
uXvSgGp3A1Na3xR8YUiE4gMsAI5y2cf9KKBIPO0neXwRvxpKKI34cNPWTDIwaU0Y
fxYBFM4d9jsEKpUHCp/D6HhT2RueZUSycZ7VnbHTZUCv74tVZYupzZN8mHyJuqUW
cOnReMYl2N7v/IdW51xPbXhxFoyH/ulHiMWxJtc9mPplk4c5J5ECzD0X8jL8MM4v
w04ZOygSUI/PqI/z6fXfikc0TOmYyK3iYTaRTG3/sqzJwzcqm632HKugPOL8zyJE
SvHSP08mIMlKOBVTf21x011Wtow0K4EUmzqyfjk8q9DYsrtCEojU+95cGMZ/g7Gl
ysJ7mGlsjU/xjQWcrbnc6wR2l/dXCmTOPBCSsSmYfyQVFsgcAn6k4yZUoB6BPULk
OXP6J7+MaUi22QLRV4gf7FBm97q8VE6zL1bF2SvVzblHe8rTf0Arn/AIHAz4r+Qd
hghABGs0KQBTrJAiVa9z5p0jdLlOO9oNZpBtV8D/lPMJHipyh2YuUnk7c/ve9LBG
hK9si/BmtwD/dJz02aDI9/S4IXsnE1qVPj5dG+X4Brb3lF4AeW6bdejmRk0BIFls
9ouBFgrGkq2tZeMx5y2N7AHCED2PBIEG/3FrTMyJaw5CMa16lTgUBoCRYJJyYmKs
1bxU3CdTqI122qbL9OL5G6QS5Mr/YCgGmefBejuNYyPaQv1B5WqmytTw8oRbTof+
0u6uuhusyTgJEkjUiERekUlZHwdJVBd8Urc40sVwpPcoSCb9bcgpA8Gm3Px9dWAj
wTh31gjuM6lLCSzcN6hAQjSG7KFdp+njYsFRwM9ujnMo/FfldseOLWTpWqNL35rW
tS/GkLLXbeT84L8pq9OYtWdDCSgdB0qMiaHrAMpeesyHqLSEXuBUnFRmCn/WucdB
NK99Hb4udZMCYPv2qIWtitSS+EKVHgWaC+oYGjL4kQIwTGjTh0pfCvNot7DAOkZd
yv3JvpB1Vag5V/gznO3Exnmz79LL7vjsvR9ltQp4OrPxwjZ8H++yU9pSjjBgNP9E
WZUzEFSCW34saVwU+XHlfqDNILO6c4N9ENb/fkBCCQ88+kGBvRSmIatOl8CKs6+O
YkrPYmSW7FAKgS8yeuGaefB04LV9AH5cqqFcZeRChEwLWKNgdHPP6vSsyZck6VoL
RQ/+ERJfWoOdV2WMyyyjPAp0vJQ1cOcVxXjDx8E2OiCRobRwIxscRN/j4ol6FVox
UaHKLkrbZOa/2hJjNv1YXgPowYoWtYS5PIjFCVTi15dCVUVFFo1C50VJgIbWw35p
fafox+ET3yjiP0ItpHtbdVXqPcdo9A7HkL7JRy4l4EDO9rNXtDTttOZgBrvmHM9e
Kj3oWYN3zMm89uX9J2Zk581A9TwHaGDpRF4q149t9kREXrZoc+C64cY6eb7Ozbop
7VOjgQDAvAVrsigTTEIWV/v1i6DuqDJ6AuGxRSEEzGiaxOV51LL7xSJNOwyYV0Hs
dBVi82tG8bOVSpJtvvos+p3fW8tveIkQAk1DnM8MQzWfvpGjmr8kPLa3TtxWMM4l
mLXnQgWLFMZ0lRutx1kBIuAmUJeRp2b/5sD+Vj8dCy+c+f76MQlklq+a8gqIbzoH
tLAcf15V0mb42ShUnbUCVVNLxlkzahKxChGcsuOUfAw0lX2syvwvzUjqf6TThsdE
L8naYkKf5dexqtjTNi0OtUGwkS0WqILMyfuISBc5ybJ9wjxiPb0kq9nsOvFmK92K
i69e7YlspgBDtKqk9Tt+TPN9sCpk8kAX/8eRKlZ3Lc5sR3UTIekkokMq05FdBs/E
JbywR/a+DHzDJX+At6qYLSzYLaaCOfAcUXAgq83+d3BFkTVJG09/0IBEOCYbCj/D
92RXidL6wLnssmDGHCX3eVRp4ojlk05AkidJNpzAo4zv7FvAfyr3SRTvI2Kz2FnB
eixckMlnFhGc+qrEAB+TVUyhFnfzWqgTNjl+dnhgcE+qVA881yAtHV1oBeGK7867
TTajJXrD9V+QoH8YNBPb164sVesAVDYx7zsy30FLmLEsWBMtp6VlTAdZckTpgqwV
NRyjWcwi7azloh4U2+Cz34Q+OLn2TEOoy6Ji02HkTq9JUPS7d5HnptKNJBtmhv46
+4oE4l0p+EfhdSPIqDDiMWtQUvwtfikCUCB/0y6yLW/KTiTHwRWIZjeKLA7UdRug
K0MODo6/wmo7fe17DzjjQCmXnIQrMHJe66OEVFT10/3wvvHeMOBvdh5Rh1xBkj5Z
kFaKUMnx+jImxOCkF8VNJqWqeHYd8L9GcCacKYTT21WTJQVGMx7zG/Ib/cM9HPUA
G/symvZHEiCIJFmLJ3RUEYqJlxxTtKUIJL6vHhfDUWSnagtciBHi2ChhAufegG5R
1+jVNaVhAATX/qQSGXF97umEOudkcApdL2VPxtA8wk9e1jTlk4KKGO/k7Eky10h2
S9RTOgeI5EaBF8htKBRihFJSo4KMSs9lVKYGvawOjw37HaTnHJi8y11GhG0h3b4c
B75nZWbeIeHkRegsgNaU5brrE63rHhO0L9g+6KYtOT8ZX8mKwmUWn3UgfNQeLedI
5/StdBccp6EsUKZA3HqKRxmhO4L9xdiTvNmxHHC2UzU+0tPUMalCCZjUOoyEKT1U
QrtXDnXJZmy7JARkicid1MNS8deDKZsxlp+ZQz9LMw4NBtvSFO+0qaaEU7Ec7oI9
Ch0lceVftKTe2IfvTPYBFsW5tzzoRHPeXNTruMRQmHmlBoaywvcnDkYU7dyk5ARj
bK7PMqOCBNqLy8HLljSpWYq50NIwe5R/7COGcbF8v2og+i57nWzlzofR2hbGErCo
YSBj4yMINooS3rf6xctx6pF2b5m98YNvKJcOFsa1yDFLKj21ZylHlIskHAuwvaQs
SCnytwimf/nwH3AhiDOUSxVXLoi9zDtIeyO1ejK85E7sWZJ6Z3huFx0s/i4Xkn2V
W7kjsdoXt9GTPcWUTQn9l2S6wb8fpF5+yA+e1/ic6l1QqqMWfcquOeGdbpjH6u0n
tVfUH6DJyYSLVNFrz6O2YAbICTeYniMS4U6FyuZ+UM5r5WsUZ+RU8K2z+lS2VNYp
Pfr+qK16hwUPadpOHpMvv58gEPWM81RhZhFueTCd8+1s4iGtdTLAQ1so0fhjBbaQ
7sA/ARNJIq14E7dqhaSiKngzxdg1p38I4hx/LzbykkkZo02FoRPpcy6Z6G+sbdP7
sysSgEs+4g0oKo6WvNlvKaXSJYc35Kg1E/TsjHfYyH6aYWLzE4nlorHCjZj/jAFW
6sA7Wnn6aRrfNV6ruozM3R9gaWgFigKvqMdONb1GLSVCwQsM+k2c2WkoGCrP4+no
ahagMHx5shzt64Uni2QrkPZMmiLXByhrVHsUktlDDAr3N5rk/navx9HT1lIAVx5J
bwpBkLx3KHwV2AByWVsOmpQHpNxNMz8ToxD6Ffnh0NBHYMQoSCNiY+fAaRzZ6mUs
x6ZopmK9t5j6fYqwS+nNdlhHjGzpkg2athWhlmu6NgZmylL0ZKSLMeT3XXtfA4qE
8WJ00/MVXob22JYo5G+rqGHgGXkBgS9agLrpwAXDGUhyxV6q+NTqtu0Sr4rZYZe7
ckpqCCfm9o7qZ4sw2m81IuhBBF3a0sdbql7oW/iZNXp1ZUWIZ4v3jYJpME9qjtBv
zus+zKES5qFB5KS8kEJ1HfCWmH714ShkrMeg8qxKQHn87T9NldjlI7gE1upihy5Z
4ceKgTZ0FGs7Zu/h+IKRcOhXOsXc8Hx3uiyH+6bFL6Tyht6rUzoO3NBUzV9FFKgj
lzkA96Y/FVv1xL8x3S1oFmrxvdY6bcRmMUSS3tknGQvoRfU79oI8EmK8971sfDQT
FeoSBd+LtJXY1t/6kBcSMYysA7p8VEW8j+0oxngPOPtdfJfWaFuMUDoFwpEYPj1c
jpBwDenipgJUg/doHmqCE3KhETzdSmJVvNOWK3TvArKILyFJJGZc33huplVhYVi8
8tcW/BVykLLHtNLbdyGvPHvDcJ6FiDzK5QvDSsq8zAmykceX9OTLoGfq8hhPRNfw
JMiYXz24TGO1SjWLH3U626FYn4yLMy+qJ1fHgyKGBWGEyXJqlxFYl/9Y4zTMopdh
IewOOcblXRSBImgcEIyP/B/ubjLHjRnIa1jRBiqU00DI76sL9K676Dfjlhk2icoj
5kMOB79O7v4Asni26bf+DmiEtUDK/EOboSvabY2jQPdZduD6ecm1vTrxASZvcQ3O
LiJZHnSJswDTnAIsAXVOrwk7zebcvsGt1U44XF26C+Mfh0sd6ULvsWmju/4PEjSq
Ovz0nRrI/P5VjStyqy/cCtrAby0LGT16g9v8YStrsNOd6Ii+m2WatzQ3SaMrotV+
3e9+/RGYvTRei0M0J8xOitmIpxZvOoLH16shU5SACwvQuXWuFDWm/jW+TjLguC8l
q2fCwmBz+9PPqpkyNiY9zQWEneFslxUe39wlSgP2HMg5aPXRPxl/pTMc0Ojv10i4
DjLHRIEyDijpMvY6w7Icg1wAEDDI3EQ27g8JFzXj19X0A8hFBydB/FT78PxOdCtw
6VJXgmSr9NcPHMqRl708JUiqYtCwYpJl4/bQobC5PL1/06EFvKnOxZI8oxCBQEoG
oTVj8PAWHhoNUkfKfMkLYQf0jowpIQ+bXaMgYejNda09m8i7d8p1iRlvaUOpPwtL
XWEGyxJsIU3jWSoLxzWL/jdMKC2L5Z5qZVpHLtS4kHvCyhf76dl3cAdy82XEF4Zj
PlpUuCupPXVPutS2UZ1DkeTjytAa7iebcMaZhLlKn45vpzkx7EqsawQwEe2nxQm3
cVqghDq3v34V1ujHQtZywRdKYWjYdnkUGnKBjXgaX/3UNWThI7D1pIGZ2wQbXNWw
WPUT+grMOv1CbDt9lmdqzzmqVx8QI6O0WirdDrJ9PF102A/y8+l+Uyb6m7lkLUxC
E2cFDMluhQttn9tO+n5UdHnY+4gsliicVMYnbv+6v2GwZnCVZwat7jTdyFnOID8t
KZH4ddIf+cjfUMzieFsWZGbAgrXvYhosdOcWM9kQ2NyphCDs5eGl+t6jstbH35bY
v8+orpi0ZspiS5MZg3vUMVhDdH3acv7UwVxP/L+OprzcdONer8VLP7VSvD/IGACy
yzvHSRz5p3p15MrId992TZHuRKDkbjj0FNnYaqhnlQAwIEJG5PyQc3iZIqCgmYNK
x0okKkPLm8oRR5Su2IdjmzOAQZLvQFXDFQLOcQdDaT9GA49j4yApEuiYqVycPAr0
TstoVado4tYBqcHFrMhKsECueedhSKik+pAbhvH3F01Kw8/L0SH/1vrYMdepXstW
J3mTJcacN8Hndfsk6xYkjmX0uiHLMp+dRe376jpdZUPYfJCZpW8jJk1nCCFxVGg7
4o/Vh81Y3PrQMYk7uEum3iP1f3DkKLRvRhG/xzAT9U42Kb3EKcgqYzSpfK5nAVMM
SyNSn1YCrYZ1TX22OMOZSWjLeAhLdD6e//QfEkRu2Bqnqx/DuIY+I57eF092ykIi
dYH95nsv25bTc2KSpsyFBRzXU2z3pnpMbekHCVAjvyw3JQcYtFVJ/qClpKXz8UvF
kLSnX/e4f2FiSVZO1JMv1O31RvBZ2QEeq8gWgQwyWLaMBHG8uD0q3n47X3XJvc+k
v9zVwm3Mkp4I29VmyOYO0MyzF+84sgCVq4SYpbav31f+FIIlbXWe/UYJuCWJOAl4
xdzfevstYq4eK2jzMGTdrdFxyhw8bj0idiVX2dYgcLYIHupiaQrzG3Vt61pHr/kl
s37aDlVsiPqur6JG2v2k1CM9rmraYZa7aHo38sa6/FDvsSKSZzPN2iJsytzcIBYW
Ristbs72aGB39uYUS8GrtwGUfbiKFx1xyC63RGeOzWobvHditk1dHFYCLRfi39Ev
OafDULnS0u6t5kr+XzqJNT7UqLF49WAGzBVoWFAdr7Yk9lqHQf/CZ9p0BagKoBgq
j2ND2vtH9vZwd1CaXG+9pzRYAx5BQOXzQCgi8ePXYdqEv6ramOYqlanz/g/7Q0xh
mE5WgUPk2xH5YU1y/rNop1dFYU0svEE9gbnYIaCrT3W2kScAHEyb2yYGi3Mf9Dak
ggYqgYme96wRoaRJw5P9WODQ8rh5V03HwHhyI+KGXn3tM64KK/P9m5uVe+cyuCNz
bkZlcGRn/Y3RQ44NftDlM2mGfeuV2ctcwXzE4L5isoifvLzyUPG69bfHvrWfT/a0
bz8iBqN0zLUDCUjN0vYa9Xem9wrtD8E66+WbUYDZupLTNNZQg4S6gCw7RyYWwSeA
XTQRYHhdVbHnFey9pzSKd9/LI5DdQjT2/4mT6bu5kAevcqt/IqteyKTcO//KHZip
3Pg8tnWgu6aSUiD8CMqLqBPvHY5OY6JI0m7xcKFQ8TumBFKcLLsn/aea2MoOWW7l
SqUoUigJNYZUX5DTMzQMm3YVo4YlMYUb30MIMJK1OGk8CS/wW5WV7L0n07+eJuHR
DmAIeOF7vLeVgLmWXvbr7aHP1bAETgVMJYdO5tOv4M86V7sfDqiW8dnptzbA1Ik4
oFRGiCGThTOHPOBq7lqidRaXiAdl49P12XhG67CM6g6RtG8u8Xrj4hYB8sa8JIJ6
KtRlQc0oV0EfpWF2m+F2YoFs9SvSh7Lt+j+/bDaeGt/Kf0Iu3jIeNEw2Cdg6+kt+
enb2M67BNDOsjnxqpFspTosUOCkVcdjOFQmUMScTH2m394K2nZLKrRr5ARtFudQo
V72K8AC9t8FQOsy0f31ajyYmWj0WZnNYlWwwNLKlWl3dEELh2XAXvNbOSiCUMfs8
GZxbX8bXSqPEWK+loA46LHRk1dfAgmKILGniRLRpuGtXu9mpT/T0PrbdKydtG9OC
d9XGv1cRBecBLvyzXlpqJhorSCQmoj61mMqqm5pNSoSOkMR4DcVMzStyFbf8bqrv
NxUExMpUKGwGS1MdUsl3lo0EDumModTtLuUkZyfpc7yc9dB9LAmh5D5IFEJ6V/iZ
EhUM6aKh/cRKkRxUuO3IRngQ98/TLZYZi5vDyUf6+BWJcWiwHbGN4q4mZeF8TQvn
rxqHsIJ3BHW7YigKzFLd4ptCScce9DaKbZ2S2yUaxFGfeKUL8x9Y1e8tgXCBB5hT
sThS2UaE6Tj+JKTW3L6OSZiViAm8+JJXH8qoNqXFYSxae8QNNmKesfwCPiF34KZV
VxJ6U/yZaUHWpyOoL3UxC6dUpFfjvyUlsMcCKkXd1mkXRlenrbAW+ZTc+Dm3kAR5
Bu4icj4hYviYFCo/+7OBamscLOLO0CTd6UVfxlv7SS35cZmvNwUC1TkiIvf1zcp3
ihQcjQtwZBbjY4G8U5ajZz0Fs2hffoCFpwYV/I7Eb7hPPfTDdfoHipFex0L1DQxb
pAE7llfHV9yMLJOwmf6/s0EFYzUlHnn7llccVFR4pDJd9MCatEi1CHqcE9pyHpyZ
hi9/WgBKEXf4FkqOc1/XZfJNS7doCSdAsQRc8wLkyvYPVjV32hCVbhFuV13Fwpgs
suqSkg1Mto9g6DWvzEFKOiTNgGFGc+d/L5TiRNuViPyDbczvoF4L+4ijma8E7TA1
lQVO+LC95evETvGQIHMrERq99LYKWjhz8gnuSK/PbgiPmvEQqHzZ/PBvkiJ3gZmU
wkDAjKUlitn2SKowYa6biz8D42pboOOyXRVWdDox9NfAJ4f1NBaz3b1XT/DggjGi
yVPSI53eI9IdT2Ter7yVp69Z+AtR9bJBC+E4/8/CRh4g0yoNRGSqMkXjGQYl5o/I
y4AIeAltJhR46CWvnV5LX2c+tA1O8uRuEc/4x7AfUFsU6LuAIfZP1+qhj03Fe7d2
mF3WZFiAZkLbvN1C2qSTCUjqUiLJ1bQ2x5ys0AnXDoIaKbg31at4OxGbWwcyb+S3
6BzcAXFTI9QZ45v+nz1904Ub2sbYf37Clvxj6A2f+0jHQm9WnfWHbBQaq+IQ+Gdt
PcOUPj2xIIxUG5oSGAkNxP4pjEI3a8mvLbwzTMXQNXJJgf05bWFaipntrFxFXThI
AbsiaO/n9ohZuHsEyDnLM0YltrEIt8TiZCsqHIqz0SiaTn53cZ6NBz0UCdqlLPqH
1CKNSGvW4huJCa+m3z7erD2pFMz1s9WKYS3oPxOkJa88JhfcMS2fXeheGMqzMDaA
x0BXAO5QhGX3mlZPstnvrQ1FM0/HfRLRbzYdY7U93CHv6+K2vbDzcRi2AWwx9kOC
z2lP8s47jkqxgYc8B4S9tdMwywOOCNVcklw9hxMTd+uJlqtcDumh+02PbzaThHch
58eOGsnE+n/3ImidTAsu33VJAhj8kZ6gLdQfs7mH5y61JUwq9fF8i47VCeQl5P5I
lR91+itGue1A9TUCAqUU48jujdTpjdVYVukhGWtA3AjeEBQjas6keTFmYyTQ7fma
PGO/NnLOBr47Qkl8q3Sa/VsIVqDB5tDw7D9Htxy0IfSGlQQ6/nnvgmbncl27GJcB
cYrfZ2sHm1z8Z/ONg/xCA0d3Zfq0rlGqAhEeP1ujkO95o5S6OiYHR5Ea1usvvFV1
oK9g6J+9ML+inuI76osHjOc3k3B9zU/89DgCy8eEOEfAgkk0la5+BnKF0lI+nLR0
ucqjiI7oryvQ3DgMgk3aRGTkaErl4ksRja4KvnAXnftxvAhbTlvBUbNPowQIKfBT
h/8/vgJ6zgo59SCc1Ay1gdkZgpQnB5tt8RVpialM7jOwhzlIU7xTxAshYGbztVRP
BONjztAK8413VmoCVNoADnASckYDMzoiKQjy6mEcllN/881FsP6fFak+VEe/t5sr
Frh2+jJodo3ELGzMfKfulNoN7vF6H2L2rj0+eaZo/1Gxoix4s6f+TnczyTQ+xu53
u48l/YhWxc/J8eKPonvPTYRaezVONZFKJNKCDRm/99Eb4kmqU+4qGm/lyP1f7Eiy
kpWPAP5bybkzEj7mka5iubUMV8FN8nMo6Q/6PEFgDMqqxllzCeN3zrN8+3L54Dt7
2MvP/Bxo3jZ6owwVTAQmVSNpgQmwIvoVjAqk9g3MCN/e1CiK9H8wr9GD2OdqqVfx
Yxi+/ENuzM4ZmxUOuOLR/PqMsmv+5TN1towATzLuM/rNIGrNCABIRrNpidm85cGz
nmt1IXTpyt71j4LIBMnzdnRYx7IZZI04LK9kjxsdSybz80+b9EaxsWemFnvtC5Gb
Et12htQxFuJixc7h2mbTl9HlJCEqNKzVfBEafuE596Ad868CHbagD5pUZJc0X3ss
1m2Bjrs0Qt+1A3yJ1X88cdpKxelANi+4UTdpMrT8ywdIsmYVYvXo/3IyZ9eE1ohr
wk6Bo3sd/jo80p14CoSVU9/KYrOxN1me/kVHDGt4gziyIDEwNyBrq4rWxcrY38OO
rwhlY4O1aSa7csJ90IKWC4pq2hQ6TINEUjwRT2/oN8/D0MBWgbv3rXHZL5jcNJAE
S5MrvNP0wIPWmRK+V/CJUmPKr2TdiEtdatlBJGLoYQr6HgFY8zVFccDV+XTSuz+c
u5FEVwQUSXHfjsOJV8hSkw1XKc81v/8wdLxVwOpPXpYPPz7d14FmfDLRP8js1xql
nTHyQzpwqjbH7iFmY+kEyIc2ynP7YdPYHsypBAXQ98UXjWMchaSzMoE3tO8nlGbE
4fxHlrPc0jTZ3/FVQ2Ns7RndO5tOSjgaCu76h8eixmAjyKbFL2rcLTG3d1ocThQf
1NcC86gAtUjqTlE8U+RCiwm/F00jUl+kH6Ne2fszpkI/OkNkqwMxLeGmeYwGzheD
S7ctal7lBauHiLzJriDluWLroBP/YehdYIjU6kjhyZFEXJgZFdDbwyXQko5gvOKt
frhXatCScrnRICS73uPpZnHZ2+2q1l7n8dqoN/65iT19gUpiA2KWAD9qs2jPCii3
CxETcK83QfhbNBLsZhXMO2I2Q/qA0VRE4JPCArgOHE02zU6oxYXsY2rT63gyfJSo
2bARcR4KvtGIlpdlNaHUcWFA9E8IGmdLAC3lVSR+A75ebFtqIDZpCQXhJRd8syVs
lu3QQ150koqQx6pN5gMRkS9B6xh5nsGserOVn18i6vktEYGWZozoQMRymqNjIiLt
fBM98YD1BIwGO8Xr3ISDQDVBW517Ma5wzmONRdByko/WmgVFXilCnp6mB/Ur3gkR
ZG36bwx0Ekoqc5ziFvAJxHhb/hPH54KjV9q0L/m19TWy17ZCdj4G+V3ClII6ehyb
h4wqVjisGG5So75ytZA04hp/DYMkPzbyvw1Eonhy5/T3ehxdqW/CCHO4/npEKQX5
DIcu2j2EQCOI2y5irJ6+n9M94OCmBTSQzNxACYBDE9hbGm1FNUeu4VZbpDj1ZnTh
TCYVwYBdyQHp7sF88/UVs9wMPR4DxUJ37sB1nPUywLyAHiYRFC4PcbRoIITimAjR
yrZn/9W9OKYBaSxXjFHT2Lz8XxSGtVueS8BQHtm5dTHfe0uwwyouUAgLAdPYnqTE
MretqlNjSFgOfKoohBk7wz/MiYoeVR0KTRjphZCmgQ8K/A2kybuC0Vb4LHg/8QQ0
yX3wBYkSlOucpKytikVigdP2r/2PDYPBS/kbjHo4E1YukdcgnA6vpmrLQAQPn351
nWVHUKO2T/GjCcROux5UGRnLkfYhuOYWNEmzSyL80zg1dImjX+N0Nhh37uNPjoH7
javFP1s85F59iliPHwRLjemr02UiDAZEF3rfA8Lrb1200/KrMuitUOS3P484zrrj
MNE/fvEALlw0mSInzgMDT1bWy/x9zi1Ux96N95o3fv5oL1g6NUxJrK1HvxEox4Mj
x4oR7EYoelMXYmxLL52G0izuvBl1jSb3mzwaZE03T/pJxu2MmRbKOb7l8l2mlkJI
KMHWK8pfng409sb1btlgCsiCemHMHn1WS7B1cLs/U9CPE46Mo0fbAWJfqPQ/WwLf
iaf5VgxrZlmO07Zy2/fEhjyVTJ79fTzG4suzzrn5bbkcTMZ250499kLbKdl7VTyJ
9MxniHE/JXPD3z5IqOkL67z7anWH/VRfgtCCqN0LjnzvOxZGBkvqL2GSgoxNPIWD
sqnnRIiU7LohnGj4OFbpYyD/AeiqxQsH6Uec8kSoL4CWqhk663IzlLukXxgLH0GR
++D2v/pr6InSDabDUqYyK7ash/vhGMTzWYpkVbVjv2An6Tv0H+sFWeTRPPLv/JeL
wgUD8QDqtYwNuC1sZRB2d81Rj4QZfHENG8WdIGdwrqgaPtEMEDZFhS8tMHf4d1+n
6sRu5G6j0uS69UFhLfylsAmYjx21WJ/Jf9tb0yoGBtCj4a5HR7RVgJVU3M1BHvEq
qCSXJw//1uWwiUUxyyj7NsWCpMZC84b/jiTEpY57djV5P8axrgqkpqGRhAQT12Y8
fyaN6hGAKzDJYYI0mf92Qy5r7dVKFY7b9Re6F5dhB56KBfyiZ6kAmOVusy9Ivftp
0kEhGYqvmG+e5eXKgx1B3sMPU+PjLR1OJ+AZjysKmLum2g5tlu843Wiya8XEWJU+
RCccmugc73c9OmT7DGx0FQHD/GVCHhIIr1/4oNAj/fBM4hoLbnalaQxduk2RGjib
LxU8gylMhTOg1/AxPT+to/GgrLmR0//z5FWb5MMvlcx5hRg4iEufFfQ65odZKsFn
TuLkQzm387SXdyNeN36YK9c/jcNdkB6fGHuviz3HscKhesppvFFvtUt2yTfSrjLT
NQ/5PjP7E2OwcVEXT+7lABLyENHXLG444mt4w9aP9FuEa+5h7FfuxNUPBQL+XC5B
gbKUm/x01S4gApBSjnoKZvv1XwcPqefRg1a6UQpGpMVBFuwwKzxH2S0E4VSofXkH
t50JUBFcJFAj+WZ2jn23z/KOXuvuiACQ3lNZqAvcSrEU/tBdZzcdn1a58omlylMd
JQ9BQPSViow6RdcOVdYza76+gAA4bC4WUjiiOTBPbW6Cx3jzn0OCIs/FQsrwAYPi
7cPD1IkFH9hiDoZvTIG6vyeokd0AfHY7MZGR35yOUsS5ZqJmlHrghUgBCWITeoUU
bJVvZmNnzhozE9HO0pZsOnibLppB6lOtiM4I3okwZce9IqN1INY7XD0bGLl4N62O
SP5wAujvkN8szKvb9WD2gEMh92KaSp959tyYfKRUJ412qBQRRlXfiqvjhjQWzyDr
j3TkuGMlNEzarYCv6UfMzoeY9f/192+V76tRyLqRHQTUgbURDqCFwZ1+0kF4Xg+H
VHKvCjjZCHi+S2uSCG0dugckaFC/5VcUbQ6Mi76pATryWswb2FUKg5pkBwZwt2zp
I+oZfOUZNct6DnTo9CchXyKWW6JgHPpizfYsFVmXdEtGkxofuAhV9Qx0Leqhc9xU
fCKTH68997gY1tyDUggLYut9pzDAxMrq4RfQBZANglxwmuQNLdP99pEHUr6tJYG+
GMQnxfIwbQDvFfV4a3BWWTcfHzs8PCqlf1bDcON089xNH4eRS1pqKTzH22HrCPQH
a0gR8ox77FQ6yglQ9GYmcLgs2nfaCORriOjND6kpzWD0R0+G088YlNGKffAMMZVx
E8Z+kgrh05aYxmhwqdwe26F1YzP2tg3cG8l0wRZa739Ez2x0sQD/tp9tAdVKtH4p
ua1GYe2/CU5Yu0gMU3qdDtM1hAJnIwuWYSvs38ueCsozckOtXzLwCqtJKNMOM5T9
WHrd/mOjhAlo34h7nx7vhtzdd8EXZsicL5QPcRNVC9+pfSk4ZCPVoNMCnHTmN16J
La4rsFf1latLRqbyHSmcktQ4tpyoFIkkJ0dMK7RUyBxCelqbVgBQHOMaX5TSR2F6
Nd3uvP7gALLbqkC+Nvg0o/bYn69uSWEh14qK8NJkllMFqhnezWRExCZFl6/PGDm8
uRL5s697Ft/FKr5jYSb0Xz582QGm6gcES9P0wWiRBS60qhIXd4+XQGeSp1oU8U4H
HyaqKEqoytZOH0Kc3gf7OnO48+th2GjOMSBAKtIODe4WKVnOCXuEd/C12k4wVsHv
4sjOV0u84Viey7rtQ90ne2ISTOs+4mIJIHMspEuMUbj1vQAulCqmydRcX6GhlROH
3FMmQdVETKkB5tghM2crKmXGfvbHI7Rit8kneVSiOpKAGXYHe4HXGc0QPCETw/HV
Wxp51kjOmq8vK4rdKZ1ZpK6tNTISp0PY8aJRr0M+4kJKoh2s7ZLOkDXUan6rPC/W
NgJRnFesoaK6FnL7jAGEW0f4YJ63kij4y+YExKQS8vW/6UtWSQi/c/0gus7VuHwN
YPOYRiRK1yUFQ0fsdL+Ol3qk03WCMG0KnSNBmK9JqlXyTc0bAATxqsJ1chNzW/JW
5A5bJzo3dn3SagHBARElZnJfqp/7QJmOKUbWugfoy+Yjo1NsfBEuEZuslxfKW6wb
aD8HcVKGQcP3sSj5RulJjxjf2t9rlRZkkyA6kg5AX/5h5Zm8uovfhbeuCPBwMWig
lPfbc0DOicgoes0683XAVSCeC0IrKu1JC+ki+rhsL+EpQdIDh1LXQ/EKw1B8CkDo
VcO4px2miCzNeQgUz37aJdOX1Qh4XVHbaQBvfnKNbp0sZsTkRanJT+ObLeCMe+ze
S6Je+up2mAOpxrywpCkOgyeti+brY5LdHQILU+fFu3WKjqsVb8te9JOIVuKnlZu+
9Ya6DQPHTAz+7gUR3od35OUuIdwNw3XpKuSFKe2xM50VZ7nd1ws64hmoNeEyJO5k
HyJQ9lsSj7B5QK4Qj0FyV+a/Bqp62ItWZ7HEAAGSmQ5gjyLyDLxApi2NZo6srXTF
fGGwdK0Z/dV5TfjNCbbAQkJzqxlRf6N2FkcfLiFFtCuqr/V0e1/Fp+hGHs8GNhDc
LXGXqFCjjlGfL6r5hTdeOrZ7XztQy5h/LyeIuzi7cFt8ED2waoQy/vtTXX+aIk1V
aCiHxyEzijEjRzHXV2iggRfhgw8yoOvsYUUgv6gQ47NgkL8OebEPabMYin5IXHQt
HkZKx2ddKJS3UQ3O3UZVPqxxl1IpcBo5cPKcazxyrqHtylE76uC/o8p+CHuQd2QH
LyjGYrdMd4iJRCXhREe+eOXLzGeYejWHh3TVjGPqrrerVTuXPkf9fp6183h44Di9
shm+Y8ffAR3hxp7ea5L9dJHgNaO+1sY0jAjuYMq2XO1AE79Bx3TbNuN3FCtPSPz7
54rlQmRlQVbYoulgiMEQ8zDwX/CV3FZJ3/xkQIyOfbiqWrE9ruVTv4xHGWQK8HFY
EmLm2xmOAJTGhjnxgnb3UN7RlQMnVjTDx+Xesvkoz2DYRQZz8zcK/dyJD9NBRyta
OPVy5h45jzvBwsv66JDb7r8XZ9Zp2jXB1ZCrf9nWK4tfQiKQtBWq9ODD8JneFcDj
yBtM2DjQjlsm/IzgCBelkJylxjrwLDcjxu0LF4+OAiXT1g636mEmvvx2BKJcXTVr
cjXcR25c9jIiuDkW7gRL+XxfhxU45GJqg8g3gRObk06WmKbdR0xEc6HBgI1VPrl3
NDCZQ1cMCZRxRUBdgY18fyHxx1VBbdhGdU79BFgKebpA0nUcypbL4CGpFRD9tWrx
ZUEFZDA2UXEDnKn36oqFmDCC88hzlSjjT5ctfkxdmdPQ+IwC6NYODGMipDOfbkV2
6tSXXJphmCJ/Nuww4usKGPLZUlHN1Mx2A+nX9nUeJKzuHaNITrq95mn1P++CzaId
sCnf+L6aZ77mYHCR9v1hqXfid3hOdyQkaNbgENIqK8nujyQaSYM8i3W5A8259rS/
yX1CpbnsEYvaR/yvJfdQzt/vxG2J1z6pqEluKA/iEH47sUZuTkBLBWxrnqdrVHEu
GqGc87wDL3WlBQcc/THVWH7eSDONAWRfv1WvqVpr/2EcDZmF6ak6MCDeY6E8x2n6
zCUOoy+M0PGocz7VD9RRaqJT+9z4s6IM7ZihjH91OpW7ApaHVo6hWQ/iL4Ns9LVY
/Ke/y2GS7fq0lJQniFFwk4hrKEBRGbRjpvahNTixLUXrX8G+cAFk323r2Nx9ldIy
pvyETSw29HPIhqT5FmjfvKHbaQdG8M05hu6gfUluiHZtHzkLdynu7Um2XMzOSzdV
gat/XcAaYjCvxsbMIp4yu2M3pyir1qEXMPAQ2wvdNRSfnVKdEf6/EmJEKQuBMOzb
FWcgJ1h5dnW9PjGv9wOkA5AvOb41NlnffOKSwsjtL+KFA9Kqys2R0KdkMOWjs0+M
B1k53YB9zZM0Gj26ZbFU6RKKKbOhgFcPLtpjz9DNpyAa0YUsBZFEzKpwGF7jMWw/
z2StGEoMzKPEBbsesbwl+GAS9vNoeg1UhKRcukQbxJUkP5UfbIOG+B+BEES4rL9j
kWckdp5ee/czbnqRgED3ACrPtK8bWWTygGitCRyd6wVHKJLBP1SciIW4Dx9n+48m
XCXkRJ/P/Ds4Q8b9U4fki+Is39D/9awX7VmDrKlamRt4pksxcbTtOYvv8jVhuiqN
RyUM05+rCMf8ZSiG+y8iT1qanvtiVoCL6BjfIWIr26XN/5Ct4573vMdtr6zm24JW
`protect END_PROTECTED
