`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfLkagFX5AdBCA27jkC+Mxbr8NKwyhiba8ckua05wgR3L/v6wqwOKBwsf9FQJGVF
AD2T3d2OhZ+ZTFJakKpc4mok8I+OoOGPcfvviiCSdphdxTw43OBs5G1EvnvLT//R
BrEKARBePhvLFyde2weBrqtOwoIwJt4jqi2l5V1K1hmJE0q8hAwxsD2y3+oqAxOd
CRbAjnbjpyupX9c7/+w58tjZUGqYAfMx0GiiETXG3WQ4XjWC7CsuZHrQKF17PX79
W9eX0nAK2LNPPpDGyPJWMvO8UsWD+ODPhoGOKapi3WbMkDKnfCH4mg9AdRbNdMZl
SWdJoQigl55grof5L//2q6t7UZpbQVpHI/jc0jQXtAwb/lN3/Oi5LP2dSiFB9Rua
`protect END_PROTECTED
