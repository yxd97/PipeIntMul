`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
37mmrH+D5koF8FDX3h4kNZDQPAlS9LOpO+T9gARHJGfF0ezweJ/slPMD60G1A3fu
j59lVQHZTUsQNS9GeuWp6UyhYbO8sRm0h/jiK+EXR98NvMP9XEhCKZf0ARXc0eNJ
0sjf9hXKtAADmonExe1oW6vNzd0/1YJi3AwUlIjlxwBWnXRFG0KR8bCZEWNjJrAL
z+UANA5bfW5X58saqZVn3gQ9OmBCmZBYvs8dMcfwZq65nQmCYhTB43BRH2Xn7em1
iL0GD0IlS0YHp+EfiZiIu/Ld+Z6HMvgA2ehurOw4VjTN+ggF6AVOywILm2mnCyd6
Wyie4aI4+J3FyJ5WACLJlqelc6wfXs1kkTwZfJtv2Z56EQGJVJCQ7bPuj90bZWhu
gfgFV7YqVzu075ULkD1BtjbrNk0JEb+50baUu2MZ4ru3CHWq9CyWYZevZwjf/877
M92Kdw8SmuR7NqwDQL0W5PgOeWMLG5r9EC35C/CDih59fkV5T+qb7ElD0F3/U8kb
WaVBzxJTD7EMDu7zkclPMMIVSxk9OdwZqKxHOLLbWL4HwTdH6B1ZfKIrSGeNkchZ
QUya3UrkNq9fnBMdLJIvQgsnjvQd9AChGBh2hZZhpzZA7agjZAWccPxQqxypCmjw
53OiKiPB3RjW45nKrZaYvYr137ukqcY52s0CSI560PchL6S3KRqnWsTK2XlrpprN
POZxvlHeJKt5uUbv4fUeIA==
`protect END_PROTECTED
