`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IO0Fb4M77sMIHrS7jPGJSQLd+6UjSMUHd8PLUJbmH5HdjzHtI7ByIVlxSIN3RrPg
7Dr7tlA1o1g/NfPG50JznZPwNDvRvGhPGnZHrTHBAOorvYqsjn8LSJa/UdC9uxxv
/BEtns7QrXSW9C6lUXBk1Zun/brarQUjbRd+JEm5xP3KjgtMeyXL0lxm++VUuJY2
QKe+bijJHnfhFJug/HOFmqESdFCeu+fmVR8blRtzi54A9ncfoqcHTqLaVYtWH8sf
1R6kKgPkoBPsVm5CF+5jcMHtLrU1mbthhZxQgxomoT5tNHtyIYKhm9cXdYhPj59C
GXextaI8e5db9uC5neMqgyvQXTK+D9fF/ZtCV8CYH5Ui/pSWJCCCD7cDHF/UDLZM
96I+9z8ILvwC9wmkem/o/g==
`protect END_PROTECTED
