`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oeA6YPIiqODmam5cyi0bqSnP3DOTsYCOgqCuXi+RSdU/aVPwVqXodKnWmNgspiBC
O2Ly+W/iB7Tt0wfePu2RAYbV2/KXV8D8piCLiK6+ZrgWeozK/QL4FcsXouu6Aml2
748Vh2/0DxkU2mCmkTxcGXOK7P+A+di7z1+24G9dXmC8SIHPjAsWwU35g8dHcS+p
EjliygPvgVk12WdBFCvZdxkjq5Qz89uiUeJIwFG4898cD3iE2iuotuyvNv2cm+g6
2HN5+qKtVGHjO17bcJ+WKM6+tRaC8HkhiC3ss2k/ADyq9648AlyWC1fA7ncAEwqj
WGgaD1qS5CNsdLaLPvuxP4h1fxE2sIp4+8M6LTrhLHy4ZRgOfDv40FtybqP60uMB
49jusQVCpoc5TkiuLtdvnhTcYeJzaemmfaUTrD0/v+H/P3WV1RD8q/sa3LbrSJo0
`protect END_PROTECTED
