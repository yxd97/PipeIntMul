`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7ueCMo2UPYuVzWu82C/OpHbRGHVBX2hxsnl3+VI+w3muriN89vKC/gmoK+j4BjP
Nz3OWkh1qo6dR0UV6TLjxZLy47FQk+CJ1uPz6d8hTOOyEtcUkA7P4UXlAiW6TIn8
yTUepDAErT5H+MOXLxHPf5WFgu92l3Xy6N+LxAnGyo9KUat6hXJU2YUtRevY7ZS8
2XoPqdbqRAkomL0A3RvQrXOXoEqoA382LjtnZKGetfVussy0/VjN/QXqc5Fmbfsz
2341K+i+qouLhdw+MZj5fojJDNMmvAiOyGGwhrvk2HiVsEPYjsw88nWlKK/vDbgh
hAg+xqM1uF92v4MhtewjHzwaeIp88DZ+JFgciiJ4k+oVrRTyNfcEQxGDE4tyjt4m
X+87OLpxku4fEwTQ2FMycqX2vrs2AW8z1uZqrbNCLuCH+2/viDq757TV/reVbAEJ
`protect END_PROTECTED
