`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmCK8vqoZGHsaTgomWIfmLoihcf4Ttz98NHHeceKEH92tQp4I/BW4BYKuxGX4ZN3
KN2l2CbPpSdwA1P1j5FIBT7QfSZMKxi/drjbNLb5v33xKmbL9K93jEoHwE7xMy5H
gx9A9pBICBed1Ot7renm5jzakvhu1YcdXczwFw6yJeVXNtIla0Fx4Hp7H8umptyw
rCQulmIOI9v+mzpoWzokptPXcKhDRe5GblwhniisMGvx/SzFIqn8DONg9acC+rAH
9G1cOhVLfCCOETD8tM7mqCay0mEUScJUx/8V83Dy7VFrfq5hZ0zg7dkbQcv8ZIvx
VGaDdjU54x4GQu/7SZnWXP3aBBmdKZ8i4wfoSBldToeIZQb1YF0GoQpt30sfzis6
i835MLpragtu3z49KWGnCv/dgG5Hlv+cmu8id1k/+Ec=
`protect END_PROTECTED
