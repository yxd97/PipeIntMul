`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JB1cAy4Xa1jkKkQnorVNb4+bNX0rQ7kGhY3GQPkP5BnVs9VxOPSrl7JNL15d0KxF
MnI86p6aleBWx6J4CHETKF6fck4zS3zV6/+T2bP2SqgGP1zI3IXcTjIQUrMIYvV8
g1MrAA+K2JxV+2oKHT3UP3zDtUcxxdRnTjHFSQDi3aMwMNvcPX/FgjcjBH8ez6EO
C3F4zN9As2ReD7JNNYVAfeCuF5lf9Tm7eKIIyXcHNlgNPUnc++9n9+i5oembmCuA
4FhJFEVMxqJ84+ILIlXvWrLpFvoIF80hkqNG/HWsq63/zQGkRaUTdZT2ZKZeS194
KWjo1UB78kVYMyBEz09ytSCCzbvqiSPlzjdaYgzszOy/N/pKaA9O9BSnL0LDutH3
AQfIEehCci0UPseoBjdLm4pbqcNBe9ZZTe/MNie7MsmxaHjOpfWPTYk2/lJDp4Xs
`protect END_PROTECTED
