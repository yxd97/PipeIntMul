`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WtnpcCNxyx/AWQIsqxZD8y3G5LhxtXQyB4wNW4zTjQ+mawobTs5i1n8MI72cx1wl
vGRxLfelfc+IOyOo+jS0Q7u7il/wry6N/bnR4kdKiELPWKuo4A3RJZ+GNpGxfSLU
yO/f2GklxKzl2YYWarKFrx70zwQoJFiLM8ioCzzepjOvjrOo5ZaaNfcM+qTug/Mz
aQjXwfrG5p64U+z/iLyi426HQTN8kr2ZxvBqvngnOjovD7KOe0pAc6LzxcZKeyX+
`protect END_PROTECTED
