`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9LU2DO0+7BVjDivHcW4kR5a61bUz27YCQsygQQ2aW82uKidIarZNLiMi5ltkyJZh
fqISysFuGxq2jZhzRf1mARvaLb1E5EXTpGxOys50QdjMC9Pq4M4S4id+hWDxkPs3
EDq4wQbpW/NnIhVaV1xl6nSdEDo4YIHDJJRGLWt6FNXmhjGDMnNh6OuFGAwN6TcN
3fSXW58cQx9rrxzpnyFUKLZzMDFnZDMBPOUMwfRb8F2UK9N57KrLJYUXSmBo+uRD
koJ4vmgqFawtATwqdii5c80/i6lkiZFiAO/87zECLiaxPfZ5S1ymLF51U8XjZPgf
ItU7xfc680OyXqRTAFqnFvHqd2QA4KKR0sn9veJezO3vknU5zrt6nim43vMZuATU
rNEC84nHdBOP4kAk+mnfpcoqaxasrYyt78JaOjT/doAMrnk+4XQvBjU02KCnlA9g
DDDMO/EHzrX5AZXM6g0pY0eqsTOK8zM7vjS/9hCqYbq7roVA1BkGBe1NPoqR1MCk
eImoCKYvdqUcAV7zFYHtitnEp9r8WKJTE1/f4yn5mMrTSWrBrCETkz1X/iK80eww
npBq804+uYyye3p6rqQN9kXEzMYBiWS03Z9+aVDiHgnbsnEGqs8l04jnaGf+H0kp
jnTcpCcRcI/OocmVMuK0q5TGqP+09iwB7NPURbCwJUElR7JYerFk6rCTf/Be6xjt
P1SW1EUr8+IegGS4u+TY8teZ28ZPNiX/PIkL4PNVEC+zR03Kn+RQrDhOeeJPb6bA
jAgGRgMs00j1qO0cWOKS/2ZeOMC1YMHUF66MTyQBIix5XYh1o9CTnNvlC2+zCkND
47ZCm0z9GRDjhY1osBOmFgPPL18atMApRjTHiJncwDnWBAi5jPcRXo2kbOpI5VrE
0W6FxXxYhYY4A01exLhvlLx1Zywn1HBHsgOR0drTEnJxrYrYfY+eBc6bcn2LcOhK
IEfWMf5ySYjLFtqNlXl3Ttw1QdJNkM7ymLH5Ca/5dXjNzYUuCMZsvVtb0Iqig/Gz
`protect END_PROTECTED
