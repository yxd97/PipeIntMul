`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bn7+YqlVpuVDVSqoQF92bwqVQDtcLgN3Tp4Aac9uqIhWyH3igc14gBJPW23/xisq
VsyfVPnBUBJSfyRCzsm0woAjdaC904aId86DJ4cwy3/IMIKGet0/36M2JPqBIcXS
MSrQKjtbuxuAJdaw4PJsk1uNv4OmeNkqRRMTEYhoIjRtRrsxwMGmQVzr0zJU85iU
IfE/wgX6Rb0tkSGOPCy1TYwA7HA1x4NhDIEkAYrGC5hTA7BLsxDmAKU0Ngmc0k3R
ugTnrShf61GNjnqSwY17kGXMuvYf4JWug8LWZZxMZ/CTYGKFxfWBhAjt8elhz9/g
0CeebpBiJUhNytyWX6RUDSFbIWXVLa//WPaOmKB1J0oAIrdxSJ82IXYNPR7mLn/H
/77cg/zMRJN/FlTeVrmkIK625gpEKtZTg6maVRqXHPJ8/R3sdVSSBoJhWcwTBxnY
Ozs/rOhwauesgmH+hP34UGqQspDbbz/n7KC8wWvQjbo=
`protect END_PROTECTED
