`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Ct3ZmWxmX88lY/OuL3PkCOZUEpSQcRJrGmE+jwFm9eI+e+h9KsPrv1ET6cCehGR
GQto551C3VgjnbVKogtCNtUt+ULnKO7kYLCETvsEEqDwEmYAzin3H+DbiI/VUnMV
A8zIKe/83rp2eoRTgm+M39BQTQ+JfF5Gvig/9S3Wgexe+utnyqqwjahB9yEhZ1rI
q1Z/kLWw41lxhKSbigPDEdSYhbRK5G8M9roBZXBmaOBDiniRbEXPs9OZJzywNOCu
1gyaOQrYqZiVeRs47ZJazR71WOG3lWd02IXmzhc9Bo1dbAU7TI4vRPYHPq7NGuvQ
xHtoKMjCezEDxnrdpYkpa5qBpgMSCN0pJnuGUIsVO+HGxSriQgBkj7BKpumXLzaZ
AB3k5Nis/7ficLLJZtVWnZjbfAN5ALmrESmHEQt7Wa0/bTN+gU21SY2gpKweNRu3
QJrJ3CPNyVY5LdRxhBo13l5me8S4s1N6UsoR/8RkaBkeFptaOYEGyJrGsBMKT3XV
c7P1jkdahXoX9RkNxq/EtEW/6peFhURaCjKXf5qch1dFgJUKx68uhltSHRyb2TKu
eWDyj88ARynOegg5sYHbxsu6b7S0kzyI/esgJzgmcOKLwvLIhMbBAV+3diGijVhi
YGzKYbXAJ33F0aFKgqZYWnPOYlYYVNmcHEm3K66gRi0+zy5VviOtLvuGAZVvExnK
2Jdvs8xYCCe+5NRVwDl6s5PKZL/DC5V3pNlaS/CW2i4Lm/p0HIcG9vajv13BLreQ
0wKPy+/67Z8u1x483C3sl1wYJQd5glS8XLRzpIJsHOT7TAoios2qFHzAF2FIqn6q
BFwpB3ZlT0fs4RW8jKlbwH8Cs8o+HMjBD7DEH/NxiskyKfZU8f+NtaacByXkdnLO
DWHk7YAXepUBybbOgBggG9XVz1h3Ub5fA9Wszw3bew+3psob5SFCA8RyGtXekQOB
cGocgMa8Xd/cHU/dv1HNX7KTrYE4l1nN8NR1ediKWDk/hI3XoVw/FJGwEK3MJMZd
qldXM/k/mLHi62q38bSNUqwQnLKIlbKa4QWJf09+GaKcjxGwTxZZlNCJmfBA1TZ/
bFDUrO8U41N9edb8Mok9PslX+yB5/jDgKxfiN2hk8PBAMGc8DBkxPyQzbetxGRpX
7itZhqlVRjCMWk6UjIp+qqptMBVXmX09uAGitlWZp8bgp4HkERDciogAzr8TpvCi
sv8ZDw1E0cEHrCwCeQyg2qDKOGaaDDrElZ5UUYC4nDp+zkV670euCyFU7qldzI9p
wUcNhBqU+IsdTrrSWK0lVTigvoIjm3rm21o0h7XtR8Axo1n73Nknqjhg7wK1ggD0
tqr+flbX+KkEUogVB2qqMVGCdipmm7/z9cfRuOcaTpS28ndwZ0Ke8qd0kaGyxiH8
DEXJsHlf+EKBDfrp6sfgPsbg+g2NeE5IyQujYj5lCY7s31AU66R6gOb6st5ITu67
g/pP+dw0ejzHdgnymV2ShXe1Pt/Dlmy2N7OTLkX0H9vcJzXqrVhcVl4rnxlvmMqw
bmicoTE/tEtewZBZuetuG7kf2z9zHHs9nOvXXwO9UTugdWQOga4NuRkW0EE8yyTl
FMPiGkoSjbWSpJKe5uxaYu+q29kq08KlxWs6+xe4523FveLuZFty5eroXPSoa+7i
Z6Fvpvs/4gdSAuLZlF3eftSbrJxrMvU1iiYu5xBx5JIm+Q20ijyCl6OsCeRLeoCC
+1kF7JSGIbRTONzUEH0/Y3qBS+z/htUFmugm6Z6k8Xja73mJWBfNJXaMsNawabnO
YqO2dBLrp6bghvOyrIS/b0YHdEucdy/tJTdShnGP0f0gl6kgHdyus0EktzFrRUOv
nMSfSSQE0x+hyfaRdTrOMjqSRUelnJ9jf1H2zxz5U/hGLK7CxVu50pIg3yqYypmu
iBoxjoaMItiLcHovR/JMi1xnbryM6TCXMCt8QFTxe9zc3LluDQ+cDtvrupilkjMY
OqoxAJeqjMLnUecOQISmNwlpJZA8hfwISzO0yO2eUtgPfWfXt4i6AoWlVH/xRGcb
XNuIJV5dal1Cg7/vT3b5k5IWmPdKNIQz4kL+k3nghZuMDkql2xagLyArDV+7SbjZ
FQzNNjPku59bkLNcLGQiazEJ+Opj+IJNuFxDq9j6ne6mGuTdeUly2cZBJ7O3fFvV
QvQ03+uDrMo9ZQUzSCx6IiSd9kJz4zSFQcQhX7DP2G6Yop8u3GBIVIJernfXDT1n
y2A15duotSUVXPNd6yMS1maEN73yn7EJ/qT1DQp1kJrk+fdBTkVRBoI9tFHqDB9t
xJcsm1NC8EBqcOnBqVlv+0y3v6XcTlvMmWNj75UqcTRZ7LnJE4Lg0zfcBfCa8xz+
MSpTa5FZRa2cWen0ldfcbNEVim8AiK1IsWatqe82Of6GJnsYYvbeN47UpV1LhNQC
U0ZNtrj5QkW+4voYsnQ0Hdcc3Yv1HH5rKs/bi25zxIV42B+mqTXODprl4TkWZCQt
yHdqkFgXXwbTE6CHIPSamm9KRgUQo+W2VhonZsXcYpjbfD9zKjCJvvAVFBp1XSiQ
1wcRppgNQ7gsGFfhUnGmUxF86vcx73CxemPKRtj5qxUcsOnMk8Q1DA64qyZf3o60
ItP5EhhSpdp0etpQt8x9Yjk06fOxv46JvhTB8WXFPHPVmiwolBQgXpp+WsMZhPsI
w8cIWQEQ1+n/8BL7P72NDDnVqWoT0yL0TshZKWk6BK5gpz5KpsIlYmQcpO6qcaek
Z5Z3h4MB48NX1wZIomZE2U4R/SYFRYI/unXGKA+lajcDq07JuDMGFrdLZPxVfMs/
pKSu9eDF5gXEX/fqqtV+YtD9uGv63OJ+X20BS28ZmLdAXNsPNGuDw8W9ZxpRVj3q
Co/LpjjxX3+we9hf3cs62c7TU7rEGUo+DoE/jw1nPyLtXqYhmN4zcDyR1n5pIwZ/
mTrv+Go8Es+nxXqMNePsjFlQzuDgoqeGbLFM3Cv6piK61GfPCZh+Sb1veri9UXhD
C5nvkWmeUaY655BbMycWVYG3I/s6x4aR+Lr96E6BvV4k++IyBkjbYR6wcMnxrbK8
SqNvaSVmZhupXCQmz4WBUUmeGAgmAyGlbsiOCTlZ7LS+j70q437TFd5vWTD3bM3i
2PnIX29Jpy3fMUxsKxpa4N5gqquj3F02PvhV9fRQUGY3UapTR4EwicXpw7O1Hsy1
AmBmxMJiqKeAGIrVzhuSM1G1NX4RP/u7vRr2tYN2fCv5/xXCOezsfdxfw5DOPCvO
62Z04TKR6rdHZsKjM8eRWzd3D/gGS4MEu+PVX7bRSiOmAfB4FfSd24iRsB8RTarb
xXXg3lIVyKYY5vFADlg9goUOu9q7vOAgBXIHW8qD00QqNgqbqOmBk555m7W/NSVD
uW2qyj9w9yEGwNtLD2UrVx4thNQ33AvHCiqvqPyzJQGVDir9XdwFfo+M7JpN0Rab
j/bb52dThvVfvqtv/zw9xpZLVupx8jtclJ05bVgjkR/YiGQ/rqWfI8txCZ9/rvtB
v54RlMZxKp6uo9Jg2u3EdURBa2phXtwIM27Vy2npEhuNMnqyV/aHEBsKn1NBX6uI
/TJGP/JJiJ073+Sr4HIpmXYCEDQ/Ym0ViINATgNgUMYrZkVFJ1uyuD1FLhHNaJ9H
QV+XXeAaDdYfPVTs0EDhu+DX01s5sOBEMWZ5FuZxWS8lSha8XYMVLbXIqTjXnT4x
JSA+APNOuJbULwml/lqEbxGcLUvWC6+3yNoQbVKpYoazQ4OkeKgGil2R8GVjPA7K
8NbXGtr7BJTr0RG6W5QNnqBJ0jMFL7fjf88C2+IYG2vVCAQXyfPNLs00uogJzWE9
IGciwUve7p+pa4MtkoBb0JAqJrpZkrPHCsN63TBrk2jGPL8G+Gkj1e4m6yGN60TZ
yGsmZ7+BMdLHss9rQlco9g/C/eVWWLIQV7CF68ImbaJtPJyn8GrV8qKu5f9LUl8L
3vm6s/QdDqto17qYL9nEZl0OCPujCz7qLsJnv8x09ZaZ7v+waMGlo/2tILHGDkD2
VJBtwOPo8ognnxR1UQuLXYncinqY/J7CT4dGtjjFo4SnBCaDxFaLy7VC2WX+jbka
9eVjlI4KhzFSC6x/i3sGPSg9aAbcKupQXwcKWJUrf2DG8w/epf/McqEGaFykqXyK
G8z3q7lhX7HiaHqphOrlXseWF46a4S2i1Od3iKkkIiS6ZnsaJ6ea0QedIj8ms498
NUv/3Ur43cSRGvBEouF8+NTnINCqXVpVmQM8nJ9KdEr87bkUDmhpoq/AdhUkG3PS
Y6pufcXzJnkFeta1RjaE/CTGlYGJ0YdbRZPkKA8Vd1Plcgcic+nwWoCYOtDR35XV
Vc1b/NnhBV06Ib4PSDwQnWN0H/dnWkzuqqGBiGOERrRTG/+X4vHMll/6B+mFzsJe
FtkICgo7Z0yV+AP7BH1xaAp8080VrHpvtEDRybpEdNjoWOGC2AcCaBDK9qXLp84C
Yq9i1oBqyQuEMAxUiHs1es7FGw0NnXpXb5hb2wJ9B7y1/W7nRQPzjSkaLH3DQxr5
adDF9XCYEW4BXVmYTAZJj/sEfF73ZB+kD0+sb7SB4WA6EiDlpSppLOSkmGpB73Q+
SPIHxS2sWgDtwskMnU0EkzqbZ/AbqSvvE7iLd+7E6mlWNU6QS/+U9d3v4ClX8PpX
7DdztO+1HyJLBV0D+tsanDzLuPdNcZ9RkbowKRSwyfg+Hvmcfa4wcA/SZpfuijDt
UOvGmz+JT+xiyv3C6b7Vk04OuXc5nxVfH6xZgc8Hibtb4xD9pd8ao6DO+YasmXAP
qhmXzZwK2JD2czQdqjc2d5/7j17GmgS3gPoCMENWsGc4oQ2kg20oqpXQrGSWJHaj
xccbZiuHRFp95L/NfvxmJKh+hm8iADCYotmr/5Z/NrYeSfxsDfh250mPB86w2pH8
x4rJQFP89y6xYk2n9mD7VWyyh+2wrJi3Uv7iEXfKVykxKVMxI0qxKf7tH+VQuwYV
bk6n8bQc/qosnstXEHSF9xDV2hinIcs+ioBY6qF2lOmWSY3SPNvrXjnc+qKZL0Bb
+DwE1S+wgAPAMTVUpd+xmfBfQFj9O6cskYtAUqW9ZdwiIt7UF9Rd7uvF4xTfeGzp
IsDIHD7gj4RXDv1zYbvQgqUseZukwvaUSqhTZL00gN1BRpUupJNCSwVpRgEcCqOa
fUZqwWll5aqPPATgVqnMDRVAQ3dakunSEcPrn+uVq0hk9RSjkHqX+p1jyFygTbX5
DgZ1TuO+UylSCXPE3D7VO9oMH1po9EZUHjviU46QJt2NO4upp8lGTjD1xc9Qyt7w
qoBzWoxsSyR4+QuK5tzXlzCYbXArnpAfNS598z2suTVWME9uBvgMBAkZqEnq5QEY
PouiillUGEpnMkuSYx6kbz1E7i0ZpVjSZQO/BrK3/KS13mw69MRMoJqdzZK3Dg9S
KH0LysJNBo5AJHKm+ok0oLmeh7wt3Q10nVAg5euB6Pmtzrudk7Bup5b29ed1RGf0
I9CjIkc8YsiL71DirlCMJ79E/MKYG7nZporbHapoRmvqe8OzfW8aVG9Zt8jPEj+b
lx+BTIU7ipshVVsgSQCGfBGu5dDtxcA84b+goMVyxuxLjBI93B+jGJ2Z3i+MpAuv
bs8MCNSpcTLjAd1M/OF+LVLmqx3IoytwwBOLyA+LEWsvbzXUAOxSY0nOM06fkMHm
7y2rfYkn87R6GqrMqfFTfZwfLvdSL724aEDcfrPoNaT8hwECeKX/ocfAaD3945+8
nc7Dj5TzNifzwOjyl5kYVuwoRPRjCU4XGa1RxE5OGoOtx/RUMGhW/r2xqe0rVYab
00FhyqcaIS1Ztjfx0FYCmm9bm/oFH3Fx7H4pD78xM2u2rt6KNH/YMLw3SbV8/cfH
bhOAl3ti5f+5qQmhl2K68Ij7A5XTCV5X+qGNPihDzA8UcF5LcdH2m1lHVfrA/UYl
2M+3JRbc98KSgaiIdf9no9UO3Z21BcAEnVcRqI05Vj8qv24BN1jzw3/8x5mX1CYJ
Oc4tnNYmjBniDPXyx2jLHdSF2Wdzj52DFOibkRljnlpfkAeQRjn292Dyxaz4z1WB
t8GXU5CRrZheNzom6rCS/Eolb72N/L4VgkFmNV7CHZyAq/Mr/Gl/ORL2rWVfVCch
/kl+21YaqHQMw9mnWOnWs0X7+Vm6VQQUPXqFkNIIIscFhhKs96Dk5BYqCEdVF1TL
M9pJe2WkRxNib1kfijvZbE6pBwo3YT+OV33atvkyjmomURYzB3voCAHFJnTOAvla
+Os+9WUNDcojn0MdxdMYgQqycC63zoi4jODNV/ELU0W6NWcDvM+Mq6a5pJFAIL9a
p6zuDy1JXpo3cdOuRrn+V4MqWSspIP4vQ9h0rT5orlGalci1c6ZQFNWs1SWuAlSz
PPweVWmAbznlpcQVELON+PKgMkPafqgU2z1eBNsWZZ54/zGE4nIeLMhgRQnmyIYO
dcUNPd7cNjbqn1LOOmAj0UhGVvJJAewCSccwNTZ+6DlE3g1tjuCdt3gXGtjPW3mW
ZHGhVnBzD+29IbAw0LA6W2xXosqoQALb8k2kOdYe63dGEJi/pQuD0LYpcvqnXv30
oOgL+nZYw6bJ7Ubj+NxkZLFGdZw0viowrFAVAGCQ1G7RXxJy8Au4hCAUzlQ5IHBF
dEjK7HOsxu5kTbUMtJYXURz9MAzF7Kw/iyP/VvVmJzlgas+J9EKxsK4vbA+G53WQ
bfBIt/H1gGQO6JUJLpKWz+ToNPHy7ImZyb6ios9Fsqr6IPWmv5V5OZh5XeSNcRFb
a1fczpfIl31FZdnzAce1EZlxCojJD09rhCK5bQWY88GmaYfquMMBLgh4jU2tljXn
2/m5TJVJm3NOaWszafgDQfmr0a1p6sZrprIi/3ZfQbRVRKIZsve5XcZXP02qQcaz
t895wIjao8hJigi9OQQToe/3Gzu8R4uFOK8H4q1TYbr5EZeT/PFYuazknxejBOJT
emalO+M7pDUI0UiCiVNI9G60sVi4U8xnSR0+HyyGO4C4Vk/5WkXxclHykxpq+bzX
yo59iGGLptFdWkyQ9ygZR731gDgokNnyrBVD5Ebxeu1iavqTIDJv8hx9TQkd6Q9F
kurFCISn+HF3/Q9f/fSA4uxhWdGSFazIFJgxLMZ1dhJVhbJKdPAhyjEWluC60auN
4NogWsBrcXnUQwnrQAqKGqA5Zhhd/KmSknKWFSyoNjFZQmpC6ke3wPNzrXODW78W
Pi9D4s2oYPugfbFCdTdyIgFCWPCkuLndklGF4wvhhL7ghfYNnFNnI92kLpYI9vCw
8vaXAVlhaCB/VBNfh+DwrabtA5i42pFAqkfqtrsZg18FaneTgHkW+3LpVAyNgE8t
MePTKCeeDjp5OTxojWVjxAxWQhYOT6+FmTbl2ZU2XdEb+rGXog7JCILbqPpeydiT
RGeGIMOzMIzt2pZccpQXtTJ5VrsizJMaJq0Xgk2waiphbNGQdV5yrw76WidlmgWL
X0CoObTRnHlefcNkVjfsBSvzN74sGc0r9dklHifQtBBg9qiJlIzZ8xGCrIsSY6hy
Zr9fq/mJd1nXf+53NEULWyURVUNTQuA1SwlKp9B6Is2bZhsKLDms/XkbPfjbtJMi
1MVfRqwXFjgjyX3VFt71QfWJvFcjLhvxfc3a/T6699Ot4qQMLJgTBkQvMImhZa0U
4hYCzOwjr/8XmG1y37NvVT3J0X08ZJniGCWLXb6iW+tDVcKRKUCDVcKltVtn5itP
4x1/R49cBHVRGe+Lehz8Gq76EdBRChfg7OluxMlGl9+Q8iidiedIn+GYGsYE76r8
MFa2TyeC+7+voFj0u/DEzYN4y1gPPqpdjQY0LWR67HGIwn7iV6w+Co46xJQUZlu7
2XslvfvcHUuBK9sFBXf10xRui3p9RwV41DqUOt0T3YQV5ki98Q/fgLVphI0ptUmP
E54aD1VFRUoyj6ukFX8go2cO7Q0iNf7hi/yeAK14OzQx3zwAZ+7dRXLq6Ijlwto8
RkuAa493ltChs4riBOvwEgxTFBzh0KZASYHXCh5CWCSancPpKGP1ZSkLiSglGllx
BF15c4QZkxpzn+oUDJ7ETVpHr7j6wGTgp0tJc1dEzi8Oi4CfprtiZd/yRHnSLFwM
OJ5iEP444zZOAoyJ3bRLVGWQH4+1IvzOuy1pYjuJrwN64jhHLqbnMaYAEShlfzjd
4HLzivQbedEwxR9ag6UEWYivRPGnpjRTZBvRjKEH56sxxFLIPs2SrRtLoiuPn8BN
XGZIGO7XBygJCeZtfx7aLZv8K4HPs5eUBwBhHlIpZdpXHUKAM/7lcn5PeiHYQEF4
vGNyLNO6mMHpTW7p2a13UIUC+WHVg1cUNEvsD8fLLBgKqcuuVXQhaKv7YEde9MGN
wXNHt9RGGEJ3f9tUOeGEsws6yf7KZYQKkvuuctIGjVhyIbvnbX22nwI6SXGgB0/9
1HyVcPBKa8OuPmvgsMaqvnxR57k5vYAbj8dAwv3tpEXBO0/a52wJ84tCM1eLGtOh
dK5wfxr+1z474EsHk18NRfMDRA0IMsIOB2w823dXl/aI4RBR30bitPkVnZDLvfrm
+oNU3P/7mjy59EWWoCL4ezT4OK5Qmk9KBLDzlyCJKumYyUmUXF04vih2R9FT/7Xg
26jJhz7YA8H+QhBvNYusc44EKSjBJlog3ZJ22FxKXdTMiMjZ7s8cqWd8GStNGN5L
CUwZK0cviBGzjbodHeB2SYppXytTA7Tbp1/NqD96f+r4Ti8D5TqkNWdd1OGrG7EP
lCbQ7H18RAMKMHHbSfpVTDp/qnpVmsX8GLg+qGziaJs7KggbrpsCOs2xY1qzLqZg
JVI7dyWIXB8KIOB8p0jNKR+R8tgHWm9cNNqIxEC9B6X3jl0Zf8wwePy90PxhSmWw
OpXPzC4FFH6nWO5/VOWwcYBLwqYshCXleRQLp8uHr+N5B/jNEV6BbvfEUUCRNNuR
PNGxzP331PUNCSx8S1flNklIAOPzdmn3RCykpIZl8R/jPWhN+16j0iUBBr1/B1gA
SXcADCUQTp3hVYcAIzVvHWbquGZh0eo0HeeNRbvT4xPxU9TPiGrBVFwmyUBs5uMG
OjpVZcE/w68nx8fLNYEZfrtHupCRYBkYnVbwhdfKyPI=
`protect END_PROTECTED
