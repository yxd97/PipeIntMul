`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBemZrwC151W2KXbAnuO+p5OMCnre+zdWDDnK4YAOb6lOYFRwjnW5SZ60BZIGdJN
Fazrx1GA+JJzgomMTclYxYDTR9MaYDUKAm0QD028bRICO1PjElDz7HCtwZ7/FIR7
sXxYGh8wqpji9YgHnUbN3CW0/zkk9h27bPRsZCYWe/CIttwoowo5NyNqXW27l3C6
/kscwlVryRE2e20LT9ZgaShwixg385SvPt57OCIl1wbZQyY8vlzQgulltbf9Vx90
MJ0f0kkzFAGGzv8wTwGTL6/P0nhsj3+ojQMfpXJqHlX+9CLYUlsKma8Rc3601lA5
TQfFecKACoy8E/cTzeXj/LTjsCwoHOa9sP8nQE9lXAA=
`protect END_PROTECTED
