`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rYv4PuY6vin7nuc3eWCGzjN1uk3iRfBUBtHcILzvDKnNaJuD4MNK2QJbcnp8bmm
Rom9vaWvOOiWMnIZOZtk8abrwZgbx+pR4h1sGgELHhnDs75BPDBRhygaPv9SAQYC
nM7OYtnvIYiV/OhJ9vvCDyEw6eyhcEgxZJ6wPUJIAyKh9KMRtybvWYWc9aZZ9vRV
YOcPB3gDPUKHJrE87ADF/sFoiHOx96zF5vHC94WIiaA896cJGPJGePgE7orcw530
cH7m9N0hOY9zG0d7tduJUKxH9X3/2lCZKsoimkEFeig5oD04RMcmy/7o5eTamz3M
UeY9joJ5gWyhTenlk8jeT4yfoTfHQ2lDegxlvFk+JcUrzKszRmgT+Kwv6fCntoQ5
cikzeEZUIRFZqmTKqSVJ7SJNKLntE8oUKvW5AJzootiLZKE53g50iwWsUCu0YIRy
YzIZlVXoFo8n1rxCx5qI9ycdvyrfTsR2b3W3Nw0HuIFLTFBYK9BUrC0ufT8qIwR4
gmJrWB1yxA6aBFQMZyoCJI+xXEmwJrL6qxkLslQIYxwajgHG2rhB/Uj/m9PUwkG9
x+Fx0T9ZuEjjZzv/XR2CRbPdhGJg30M0ckauJ0lAKbxK8Zq+qZpCFy9fXhXY4fWM
CfEyUp+vFLvP8SuaQlPCMZbPgjizBn4C7/BmshUOv73BOPvhKJsVXfTWaphTT5Fu
AMW1EpFBY0Shb11TERbOFusJFnmOByQKk/2Dekl7K6wCD9UA05hMDYHAXArT0/KT
8Fa9xfJrvyq9t/pDvctaJiWUIXKlSTKzcB31pYOZbdUpWRyTxP5kdHK9EhaqV0Pt
5PRInXAOvFZs5vJr5S4uG+0Wd6KapoeRh5k//2+1EgRW8Hizz2nTuTQgOh/aGSHP
VB3Jp8QCCSbYP8DvhTyFylTxFqzWsktiBaOxWtGE+4F2FTSD5f2orA7GnIplWSoC
jpz74l7YLNCCOnsgsrIlwqPAG0KRE31+Nwvh+rC697wG0pAyDGTKFBN/xcA9QI7r
csVZgDIgYYthl3pECLteFtj6KAqJFFekD4LKD/YjuQ+Ts1F/hsuEucrfs1wluIng
dxZ0zNQ3PvqfbLAlKcxhQdLYof5Xu+OacuUad6fJ35hDOCn49WFXNR+Zn7iJjNMt
uxpT0Iv3Z3BFKLxqYLTO2REaFI7HcluPwr+wJY6ZeBPDFhCY4Zz9A0iM0GJShFi6
77kbsl4EzvNhzXCYAwfgmFuo4xC4JSM7pxVXBGgex3HJQ4HZZGZH9BNbke7c/lnq
ofNjghhM96tT2VSI2XQmoPlQ88AsxdCvWYwuYlzayk1+EGUf2JjPY5Qpskay793K
wTot4kx73os15RQMZibhVG84v/7OizGAoH68OKtB8892N/ns1EsNO57tUDwq72ap
rrdQ0UyN6JyFaRe/2eBPnGJq0QJ+C0d3YWMIBvSbEG41RnUUeOOQEo4JvCl4Dbgm
IfQh94bKHl36dau/Iumt5lvOWNBVdIz0esMxTHUdFeeONLJyu3l9cY4Q7QVmsjU/
l4Ebhy68OO+o06DVc533HsSbC1BViDuSuJ/XMFxwyR7hWEYO8AjFB66tkg51bvhI
S/y+G0OKHinDjA443aPTOKAkhWiuw9JGa/MucPqKAoi/sL/lCz63DKav5+RBciLU
NBPZ8z/M4lPZNINBnWMhiu+5tEb73QyGFMb2p5WVdQ2qXlqGphhaoVaePVwc28oa
F/c0V8143qEWgxrLqIPWQj51FrcmrPjgmpvWKV5rqIqBhocoOeSUdBGzop0mqaY4
wOa+GcnNEZXITbWJrPjhgw5cQWBYm2vuoBUH78mfcG+DduGpdkQu9FNjwY3OJAzK
H2oWd57GgN68CXuuFJPWFqBWvu0L6t8SC0G3BZ+FE0i1dFSNKrG6TIyPEHJKepL5
0fggB1eVlkDHT1xbB5YD+Q2kG5M4K8yudkCAb93LkxU6M7lkH/5De10oE0CAvCCA
gSuAGCTJn9K6CpmoA9cXbFEm2gDwbb3jTlbD7jbLBgdfRc/zGV4FBQSqBPOYaA0h
iZkLvryDQuA2q07yLOCxM8Z6bRSq3N/7JtGXHx1vPOTUvWiUpgvYpwRxh7xrHwg0
bzhXDcW0j21DOL8XSVSDa1o1gbr9C94Sx1kMTDF0XqR0Qzzi2TY8esbVtfvfzUFf
uJmjJj2EIQSNxDGJw8bnsLbzv3ZEaH+JYVObGeQEaOwLmJEtRa97OPVWBkGlWvkm
+fjhCUnlhYVyhFl1MWr2yeGMwMF9VzCIAmWe4n4yE6deUMAzfwCeI0E4K29M8rnR
as2P5eZ/lr4riEe0HcivpX7x2YxQkegTSu7zwo9PmHekp+8PucQCsTTcMNnLIj3m
5GRMoYTlFylo1dBVph1B76Z8bGAFNpoYx8r4xlV3pP39+MDC0hNWgSbXzDiMsKCr
DOcjSa5C1P26+a7iz7uPJEC14Ef0bTGfCv2A7uDGAGKkK2zURwY8wLlg7gY1NF/X
nRikOL88akpIsLDQdKP7Cw3k5AfXxyuBlxtz4yElVNsbBtZH/OwPQU/3zNedP4uJ
M0dJv3myOhzbh0OOq1+/P00FuUUJprEw+kIUMnfPc2MJeH/uWPKXHsELhDQzmalZ
6TyqyPZ11kIOWvHPicslLgHWzV8gjo5VO4BCJGwyPDhPNMWgOXauMhkMT8MKf0q3
jTM8iOz1h16X9Xo5eha6199hx9L0f46+7wr2MPj3vorkeMdSh5FUGzg+k0PNCCDU
En8YN4IAVb9DlFyLzwFtUA9hdxbCIypNIyOCqUTrv1VuyMZDi/YAwhN66W457j/r
NRpCwq+SVhFTvAAxrZiy57VfmYMj8SMqFKSQ5J0lbIdCVzP7/AHCFGeE1ZbK9uBC
TklUCMreEIgyOdQlzr/H5nWvaQqtntBCiewqvjudjhIIRdT0BkaXhh12n1mMvwPw
wHKcSqf+bHiufH2nv/YYEkwFQqEK+GGEUJ+Y/NdXh9hDemcun+6laG0Tkc7HUMtv
RVTy95oGTvVqmBtm3asLlwnaJRgV9HaENRgpZr48LASnCp9Zsc88cOZWTlwwcQbl
3R6rFOM/7akrHU0osZAYbyjJf33sKCRwHlSNgFLoRxca1afyuhHM3TAHFVsa9uEj
CcYS5LacyhDp6N6Nr7blb8e7YRD0hflkQoO7OaAYg+zewY9WZQdw0HEsOcOB6W9M
l8d9o8KsGmXjwqBt4R102evOhRtppfdKEjz6Sb3fXkFJD6hUdzfnOzXX/2wAbP3A
Vklg4v6QkGUdNac6/Lms+SZ0D/BwcvAYjX/2SNR7AlJ3QIzHBqDwmN+Gm4NeP/kE
LPT07ZMf34FEbFxRiiKIodzMFTP12DKJmbpbpPAG6ehnPhFpGKKNEcyzs81eVrhB
xScTeAuk4InMwvYvBY6UsRCsTPfFLvZdXUFZUIeleBtSpNIG5eO3vxfY+ABaK/i5
zg5oN/bwLafLmyiXsYu/TnXp8zobFPewzB5yrsp06eHsS3bEfpl4NLaZWr66FSk8
9UOAiCUdXU91r9zD6UiRMqHgJkqOTHnkebgvojWc56RAOYQIN75rSEGVUKcYynwF
JeDPnzmzVdTPi2j4WhgN2K0lv8DTppl2SAt9qWpS29SVqH+FStWTe/vMSqY0WYNg
egnn7Hj4V+RMx/1VZ5ccvP4PPJyAXU3n7JNSUpPspVzYIvCGjjg5NV5ZKPUXR7xf
CoJj0pD0mLjBIw0xPXp/lh09k/ntjoaMd5M3tILrFkBU8n/gRK7fA5FD1xgFP3bP
cLDAtYTYaBIbU/7tLZmN16mvegpXIX6qpx0OtP6gl+tZ84FIAAaGhyKD7hFr5rDM
eV79+XTikmPYUuxqZf2VE6DMrY8EFjK5gIthz1WE2jjEhbDD5RJgPgWAnwoKdexz
zVxfDDqEDSrMyUdJ74ih2pvtgP2qwaERu8qfnjyOEWnKJER7i3lWLpbZ3gDfNWWA
HPDgFwsl9jnQ873+qOQ3FoLr7kuEeicQ12seR3cUk6qo0zXnlOXvg9TenXOB80VL
vjHrd0gMVl2BPXJiqhOqD+WyIXbSas6cKHLH+1RtxqIMQXG0PRW9wXSfYkpnIw84
8Kf+ezGJM765t5LcW8VNy340lcykaCNMhLDVTFvfNP7VnaqanOviyp1X21V5zQ95
fPaVjtK+sw+FUwsKXo4UaXfuzkODXYv8T8K/H4DF4S7lpJ/hsBmUV8tzZC6tyD8B
AV3N/Wo9y5PAIpdExlJZ6+TU4McEJ73H4jOQnI222h3sjT1QupcAi3xk433sPr/f
TPjy+kTq1HA1ZkGGh57j+oTppgSTBuLJ5dcWTqJp/KJglFuk2LthF2jdjkgVkcfc
4vC98fxTmbNHOh5rDQWDHpsJd4HzspIPfmRt8F3QPAcM/uc7MWeWMudqJFvwxYbE
bCmvj0vTaGtLEKh90cJmJMQLLhDMNtJH/RiLMWcgecTeK/YAiYeRjCbjbnjkjEqY
1GgbiwjI1CVax0YibTkdVXiU83nCwvTmOuBOonxHKo0CY8CTxowxMdv9bxYzG97p
pdcJ5k+to2UX7FkwO2f7Nz3Gr8WDom4RoF0TCEACgmQkrTV/FkQEqqCwNy38NIV5
U3cKTnagSrhNmq5xvf5Rn4MjnBS9MgrHQZM/KkV+oyqF+571zCzEhm0LOb1ws7xl
1rJnfXgS5//04Odxo5CSnnWcv3HdsfH6IJtThgSTahRh0bJefnkdcT4wdlZlKJsy
3ZgZW66EiLHaL7qmrU3u1y3z3uct7+EzivRK3YS8eto9WW4kjvfkuUD9DRnmpxLI
i2SAdNnVSK9wbX9luBNv2bOuEn6t5WLzDBfsciFNHAtg5JKCEiUuYOiAgCZ5Mc1l
ab5zVfY7Bsj7gJP0ZUTZw/q+fcjoGnqrWGLjlg7g+6HZCEgeTu2Zlu9ZVK1OaDTo
uz61QbzlRQgT/wUtp9cxaYOlzOENfG9s8g3pMJodUouvPa7gJo4xHMprCZtRcLs3
/NAyNCWGw5oILPO6E5eXsaaAlPYq0tj31rmkWh0BrjJ3zRje9a12Dqj/rNudm07d
MBYiw28HedNhZPN+CEN1XClCaKlfKZUOLFf/zkZXxC1mMIRkc6D1Nys8MaJZjmfp
iun/oxa9LQB6KqNGWRHPWPpy+qkCwGmkPGR2udvdL2zd00/cNr4ECYqBdJbx09TO
SHT7Bnum37CJ2gmc3iLJRDgek8qYeSfsOfqt/ydsrOTgXV/TaK1s4ptD7vuWqEea
9UeGS6Z2PEarRqFQcb2RVbfejBASSWlv0rummYThGZ2Nh2pI4D/TjR/AnfDtFBmG
n7nLkuapNGyt6gPJiue2OlH9Is8qZcJFGNUvDNS/DV4mKBKSMSR7d4zWqXhx89Cy
qzQ2gcu/7tHI3XiKOOx+V8oOHWPlFZgNzLqIb9jo7pLvdqKTWDg6rErMCtN+uDjs
IaJLDatr+tV3L+HRbPdNgbrDq/lmg3hbETK418/DIrkXaZHrIBB140IZtgs7sfr1
OLGYg80rZh6DU8qHIXV8/EvQOkUlLIhJZIkXwXG+NFdUp1kixCymuUevxV538g1u
6ZMjA/7v2ra8YAfKjizk86pjWD3p1cAWFLxAyxI9nSXbx8NOBUwffEuhy4XL/lMs
mowUg8BEi3AiUhKY0+RXOC97DMqw3C35JKLaRVw3StXZFd9MOPV9wklrPvFtOANL
5S+Oup96rP8Uv55FxFS1BxyIWTdYlomjqsA0oMz7WkMn8KeIGwz3UGbxAAqqt+LY
c6q6OWDyYtIb2CJwfm4AuDdblHID4HiCUMw7+uO6/BB2a9DuKURKFBvndWW4I7bF
zqZelmCCEvCe4nKUZ+lzu5iYRNyF8DTGniySLUDMmQbqKPkucWCIpOdXLEOtO+XS
1bIDJQYp8DVA6isHCWevf7+yJjKmD5VqC4l/YGCF967wiAbjUDOSl0BdAdEJSA7f
kmlq7v0hnqnvfgTAGqpiBLNLUXTR0CXf0m1UbcxxaPDJK5bGA34nf3BCqAjYBg6N
p8Lihu/OqHnpq44ZcrrlreFLKFzauTXFffuy+M/sFN/x3Wd2DqYiNmlnGhZQBIKh
MxaTcyz1tRhf5E8GHS/KEXtI5gjk2AeOveiWKp/TThDShBxE+41BXIY2GevNgpGP
JAV/xKyoXyfOs7MhaWG7y/M1lQSlFO4phfbEN7ieeZuCRURur+fl81Ilbe2KMzl2
lnH2ZxyoHsZo5hyXA92LOpWKdQ3Ia2RupQf4Zw/z3AFSQ4/1KkukFIXik/2HX+9Z
rSTimAEiDG0LCoiz+LSCYZLJ1ZA9ziRXkjBd51sWs9m1Vh7B/7dYv7x7ky44Oloy
SzZeSaS5WeEtisi624Oxz9sUEvpbP1dt93Fw2nzfrcGOkXPhcGojLpHSlAEh1E2p
8U6I9N7M0DSQvMP6dODWWNmwrzT5bN4YqLqfA/zELuM1gLdH1lfZuRELatQVPGR0
/Ah4hKRRpoLwPh0iZNZJHF8EaebBSYPPYW2vlFDqQectCmICrtRkrIdgVaBCW5ab
NuuBo3A7W4aBk8vS/vRp95NeFllqV1cY6wAg77uBIVmda7w88bPVrwAkPxjDpTh7
TrTOjE1ZBnV+0K9uDtdNkHOpIy54xQif6zPwGy1MRHkF1FpCVbITQFshST1/PqOj
bZhgF7Mdqok2+4wGwdlD3xtmRqhnNmv3JSIKSqTbSO3s4sB3zY8gfPIIHozP9Lc5
IFYCztEzgah03zurhkryemXE7cMCVd9tio9aE6GhyJs=
`protect END_PROTECTED
