`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P9NJZYtGWfxDPDn5eITnTI4YlWJRXoPqsCNpxfWu7i1orsyN/dYTMJjXBDPN+f4P
iewfHq7+6aig+ivKNDUuXh6CM9oS3dX8yzGNFr2vTCDpODwycTPnAjb+PI2cnj3e
wQ7peOV9mEPdFg1vgkP92JNUpVgNqJ3Z30FjNSACh+QLxzdcCmp5uBX8ymfJjZEf
FS2996w37mu5XSNGJghxJPoPf9FLXFbd18gHGDndAqHvYSI3Bdx1wE+mkYzSZEgQ
uCU79WgWOIUJRZeWjtSNyF1rAH6Q4LXyzzXnIXvSoyWIsw3i3XaFGZoAe9SZMQ/9
d4oX4UMShmeiuVPKw/yEwgvv0zyWbuLvSHnCOlVxYKU4xH0SJYXWrfoyhn5eAFxi
7owJUWUF5Wp2JcPAhIXySYCfbRm1MKbEFB/LiH1VyjkhiJ7fa4wzz84aZnmmAS/U
CD+xYLavSpjC7IHDsOwMvqE4TTQ8BanVb6YwVzdKFW024urWRxI+j45c2TmWDkMc
Is/EE7gAJQedddXuFAVBfGlwcgzkFfUhSpQ6dF7Ryg8bBttoeHbp7mevo8/oZNMo
2WpRjWPPQnAVf8W6EpoLyC3nibI+P+Z8MRiQJs1lkTLtznyE2cXo7EDrk6vjhBYP
+5vfShbbC0Lzk51QmZ/DOrDnocB7WvDWy0bxZbaBlPs47djd9RFNbKrrlsQQfa21
Nd2CBqj2LvaMtwN23T37su6aYGp7l/1EzrYqD9WbfQshZKXdudLIjqRhMu2ttlSa
eEv0RKOTotvjiceOEzmCx0xudhtKAQ/5oqVzwmFjKBJJgPsjNaAccYBSdMjgQzNX
evjG6zygE5yvOd+YQPvMUDNKAY1Je8lDYmWYDcmkRtoFTgF2NtHgyth7UlYbX5/u
hqbMXlr0PS/W2SuPCwZuZQcgS0dmA1R1pQzkeIc6R89TEZARzJ789KbmZjfv8QXL
bU/WKBpbTQ0fflj8P/RnJBmhVSwq0lN7cDmbRs/3O4kcVsX0eJHhNsIImN4tCdZ8
pVrorSs5WfXE9YqZZMqAiE9u17ujCruk+evdP4xUekN2BCB/STuQJ0LyfSnTuv47
EJOfbcCIxRFDYuzwYtdUx7OJq+/OCgSpmKnl3tXdzql3HjS53w2jt9mBLcEN3jGJ
6KJ0ljeGjuhxCek3QpV7OqWVB+k9qsCJg5EeWdelEeuiS/u7M0XPCjMdwjL83rDy
HmDPAdFYzVxwLkOTOsyTQDgYHOpanhWu5QGvrTlTMpZaZ2AbtNS7evzBnyZvXMb+
u+klD7/iVeAmNokuvxBBkfak2HUTe3xJJCsBHpJTHq51arKDxlQv9sDu15BVktoJ
n+1ExPu5AgSF6WCbDsnwh26ByBo1boBELhkTAs1LbY5VS7WOmU1ex6sATO7Lila/
x+8uv+3Z4JxuGawwdKqwJRpGOswEo8L4XU0AF0iEijuVnJ2IqEkX7Dl7V5xFb0PD
i04XpDleZvWFgyWpk1uv9EPgcjRjHEj2gDda98UN/lRHQqVwYzo7ZA+4+auiNjYK
oQlu98q4UyaODX66QTdA0O4QETS5b0kyYvIH4LhWXNQazVL7dPKP3xUWD5F6QJIK
MxyUkIQSM7jfq36ZcW6JtzN+Ht92Qe10+jx/0X/oNet0Tbv8rdsS+8imuu4fg6Qx
wdWm+yeSQXLmDh4d5uASZJZyAn1OhKWcoc5Wv09RXr4fDroupDADX7S3aufvdBwR
9St7f/QqGFdQv33nHPU4oYrkgMjLvvLjxTqwN7zUbmA=
`protect END_PROTECTED
