`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5grurnMBsOhIXLjrE3jJNwrElqTEw8Wh6UqdGxWKKJmRhVixjRY3WI8FOZpO4vRo
P9ifs8KHC0V7EC/PZrhXBN04LHS715KcTIJnkIP9gaiAVU1DuhIsrHYoweH8KTuP
CXbr6KKrOqzIPJxupoo5/TpbWv/mGa0oD+mfRsGlDB7joylNQltUWM9sG3dHxONU
sP3UeFVEa/ahHbNgo6y+g5xguJjy0KHNEWcrCOISv+wSpsqGTMjo4ibiCHyz2pCz
ZuMm7mUt/wZ5J71iYqKNhi7niWQKcOnrCk2e64TP1czbZCu5ZQK+zL9hvxQiT0Cj
BAMC8rcIsgjBNckq7ByVY7rJlKsiFfcXX06Q0cpgCKD71olDWu5Y2wo1NrjdsrLc
jfikfu0Y9IYQsq2iAFniame3wdQ1UcMjkshsQDb7jyYUqCGEWcxUALtg1PqiSwFJ
JH5P+nOncq4ofBoSlR3U3/CQ9vdOEJsh/IJronKpMzHiKHSNXYW2unaHHvh9JHTb
`protect END_PROTECTED
