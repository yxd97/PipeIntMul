`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kx1HM1xVCarfpvK5LlF6ytBv2qJlEQIargL3+J9JkY+FKhEzqFBBJOiXISw9hV/r
OCPlmtZB0J/gfXhyo4PGPxuP9P8RpcRP0oFcrZvC+lSU/fsa+8kS+yCGAy2hKVmW
1ssT1RZk64vr/PCfcPoPGU+++7cgl+MeXe+TG/NDiIZ4PAsWEIZNHb7vKO6W76iT
V0WF5BQDMm0645L0aG0ik29Ri6ZjT0piZVrvw3xxOjSVGlKY/qhZ7E2j/gSF/FOK
JSPg9zhYudsDdegzny6FnhaxOTvZVFhvFmeZvwfku/mTuUIBnGmJ5h7lGg2wBwTw
zTrfoWjSPELILXVKi4J89rOr6xCGyTPdhJuOBgFRV8ZZbyG/IV5N56J1TFBdaaHb
XK/5mE1P7qlWJ4i84q3v849rcsT1ORMIqh3WKMMkvt4a66U/n5wHyXZqV4NlYKhw
`protect END_PROTECTED
