`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWTjyDyyHaNCOQkDNm3ga5+HGPx2ZlAbPOMh98S1hzS89ECAzkJluiFRF5uMhl/B
G53mujLhunZJmqe8R+WpNln23K/M0GUohWz6ThLQoSX579phoOcvWtbWeAWirCUZ
bgqxESVZ5efGTnrISip4TUOl8UT87Xq2XbJTshmYU3qPS5Vf3kGCx2ia6oxDIQto
wh0mFbx94Wd7mTJX/KSw4WRmhUVWOnw7QmV88wm8jIaiuA9yUUquDbE8Br/5CcDa
B7pL1tfvAQNuACrDxI2AqacI2KciJGdgMSLTrbNkJ5eZBvXao1dmo4gnickrR7rk
IGH20Vmkkmo/dPaAvVJMuJ0xTXHGaI61mdlQsbPN9vp/ifRLFnwpgq/H+X3vwwHN
M+CuM0p4+brTCiN5h2UaQyK6ifucx8TCH/JFsOG9iR5m053QEhR/CCIodBhdXOo/
fAyw9piVRZPPsKk/N633ksEefXQLHDv8hCbL4dv9GKABhllnTlz+KvQWw4sWX7RF
`protect END_PROTECTED
