`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1WciU+fiMnpYQcF5e7QwZO0XRGScDmAYzqZeb0YyfzwMfqSWroUnlar9ZOYVm3ao
S1lBkpsXkW0skVRxrYIDo/05kckxkRGjUCb+L4KI9h18YvLAw9Y1wXOSWx6UE358
zJ665QP+BSJmx6Z27mXWJDlh8plRfTpD15siYbZ9sDyNG6icrLzibB108J9td0Q5
+E3nKfC50MROvk2lX+NrRgPz1wFwUFeV40o4KBWhLRYe0C9SJxC8sfGc+skXRYMt
h/R6yg9tYcOblzGD8TKJE0Peqp3Ldg1cw2CYiHZbhzqGh6FOsgL5FLD+yDcufp2K
I5fQQpHcPrAS9dBY4MG8oPA3NFer2QDZI7BckSjMjf/AiSWr1FAh6bV08RdefIR/
jehUYmomUQVWRS5CbODuJtwi3FzQ7emxKHxmTTWadWI=
`protect END_PROTECTED
