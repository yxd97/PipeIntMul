`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rBCX1N4u88LE2kO73ohuSNawaO6zeA/i9nK9cjWB8u2uX3nCuLIxk1l3cdnxSicI
s143cT5fjtGll3DBbykPnReBFvybXj9/8LnOrWCMevClwUjnTSuYBvc3/r1jUF3e
AruwsJeCxeev8h4Jc6XuyY9bhPJiuvSgr4BthBGXg5xS4H/Sh5pgRQdeIOwbtotS
sJWox6k/2YotpHxL7G1cS9e+cX420f99JRHYb+lTy3oJuF7UkV0eKL//AcbIHsFW
4UCmrssby6gyDSGh9AW0+nzCNj0AtNssm53GqzZEjihbNR3U67EXrpqnRrZFRzoJ
4eCk4weKHJ4FrHirjMH6O/VxF3WIFWZ6DzUiwWQYbGdbGuaHEgeKPQl1MNwSwpLC
t4D3UYpwNxO2872BAy5cPMQCs+l3Xm9OSQf7HB5iibY4zP+HCGCyasDVspDDKhBK
Qaa17ITTBxfBTUdNvdiQieIaGPKbJHBlOstsb/TmHEc=
`protect END_PROTECTED
