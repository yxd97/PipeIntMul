`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPihG5b0BHnpOu7YwioWJksQ2z7qNLQq6i3XUD8jPAA1Z/aFd4dmdOu68w1k3cnx
/TxiWNSRwNu2ojTvDDaLaGOseGi+LJ2EBqPm4+e0S+7c69PCpuBJJfyTMHgrqn3H
7ag7mRMovd8iat7rpu/i7CyZjVf2HRSwXNl20ixwjvNI7D+AVJUHQatDhACD2Ypv
SwM9fnxKoElV3T1rfVx1mUXk/NiSN0c8cvWAdi1zhwzcyW5ou9y6xxtWbKCNO6dI
rlLw/Ykb3wM62EOfavLJYjYLabFm+v7eWKPaQghviW56l9ezGK+xmfCQtggW5PaN
eJSim00KOQRoeS7TLqo53Bld31hn0fuz01L/OEhGnNHHT82QqDaouZ3/J/gq23Ci
TxgrXSk66LnVO1GgHWndjaAGHV4LL5oFxKg0Ng+udLF7sE3LuAq0iT6mBluq8Gyo
84WJTZtJapZf4+m6AsKnUkdeWqLbpxRhxlG8lzZACIW6k4S6EF2AuuZCE9ATf91q
0OFbEfuPUml3EVgISmzUQXAuiSUM4BOPZiHbE5X0DlIv2l3q2d6oQfV4YdL9tE/b
dLmH0HybBNfyLIQ613ZeUr6QIidCuqioo5V6Fe9YIIWQN6pdL4pPJlRafEXC7hzD
MZex6TfAX7EeUNqvJbbKxbpijBllM7tEqODgiEb7ZIfJefpWtX53/2ADExPRO8n6
oV4k1r34PmcE7WC0Qhf5V0k67C1H7uhGMIYKDW3SYqGgWHNOePUg2TC/lcg/TB8I
zWgpbZTIxzIcyf4rdimLHJPglpLLZqlQ4iyxzl4OqrmDF080V4z9j00wgJlz1BCd
rCJ5KRLppbRQVX8Lf9YvjreuZ0Je1ikQ2Z4JFu1aJYqGZC6E4sy+Ux/6BE1mVqcN
85hVK7llsOrL3EFnigMIKRem1Pj+AeOa/IjjvjI/recVNmvwT2p7Zxc0iIGhZzx7
56keHtKc48Ubr7gzY5Mu0QnSylmdP5zzEhbxBofzvHJCYdK+iim9ezFBais5svf8
I6368p6yHW0P/v+yASixHh+kXAu12UVmH2au8/BuAD6EQQVtDMAiKg3594bp0QQ6
3LqKZ70G74GKxi3sWCIooGsP938Q4BqzFWOGViWbvJ+XYRzPoKNckzhU8d99yxpO
cApWoXdbPohFt5NQPqIAoEL5OZtCHlmqIZX4ZFyuSyZYUt7iP8ZiXCQdZc5Tg2Ef
TLCFFJg47wdF15BgUJtl22b7FyUAYlpZ5i9frGiI76c5GU3tIz60J09BWh+Mofjs
+HUwQI1G/5Iid2+LVBP1IwR63WjRS9ay75+q9TqtGq4VIm2DPU3hNBZDDih44bPZ
9t1s3xW3/ocXH4NYAejec0yWKCULpB3skE38NCOc2TeBITE3BD9nb8hhdLUI2o+J
Xs2zrN1S+8tix28+I6ydR3OHaWmjOjT3cF3O0aqL59pRANsy8wsDntZYTKH0VRGG
qon2tBCiEOVIu3V0RlC3qFhkr05JTKbaPHCqsFlQr+E/7PDPVI5R5rbAWNnoYxyy
EvNS4L2IAYRLcKL9PuSoIwAkC2VY1J5VbK5/ivgs5BWgAes2RrOglhi8sG4Cri8V
GnGoPgiLBRrSTkO37JDu2cpwjhCqx5gBTnzyahYVxyaLVB8iMXTBFYjbjz+UYmVB
XpaEhPoJUIOomzSi1ZgHk+ybBlBYzeDjZsMlEt7AV1/6NSIFOX6EHDjD3kPhaFZD
weRYtcX2tVvhxKWelEbqsQIuclQMhAZnozSKdURELBbC7ED3TkZtFNzHw/fw4DJk
zAiAAUU13A1PvNGOBRkiqCqDjQu1vSo2DLjb80F3wm7rxdqAeozFeA8Da4y/hbN9
ydft5vcwzDUNYPQGM/s8EEjIUpofX7i1XK5kd+99bMgmxPgW+Q3gffCKUTM7x6ew
BrvFSW+qEPr/ZAqLGau+ZX1NU5cpCLWgO1Oc9HzquiCjHB//YkjMZI/kMSPm7LBg
GUf7JRlS9IlmAP5GxSXMNZnwZS7NlMUE8av18hX0WBf1t6WF8Igh1Qbh1jwGSnCu
1B9ihq4TMilU3menquVEUADYH+GilkST2/uFFIZG2a40MvDJ1HhjbdaZmtFkuKi0
k9hpruHqzgEum0eri5X9TnvsxbPq+HiqOWZ+BAjGeYV/skfD/K/S119vFxQ0JvGO
1bwQtVI5D7AmhemlzUlG9qR1F/jlSz9OYvXv26G0LtBjdyjdjQzq6OFXpGkHkaCL
8A+vkvrFcHcMPQ4CECiGdW328BrtuouWfQ9EZ8gb1SJdHNcvJoZ23RmSmGKbfeRv
v/CPPyPQklVB/lvViWG0pMV8Ym6eTB9XVEM4yWAlfqMXywEx5YWB5lXduREhY+7O
xDID38P2xDEPsamjd3K2Oz7yzGJTuiCJks6j1hCmF7V3qWaK7SNJ46PNV9iDAJY0
yRt0I+IPw1yr1HsdEIZDwNzX0OQRw26bYF4NgQiZrb4OfHfrPS8QV82UiQFExGPJ
nHOg5MZZaJMT7Fsk0maDmeQZlway1YkgzuF3HcRheYkTQfKMJUGpA1OzvoZmjdmo
Wu2W3oNzSrPRJC+/w1hWcaQZeTaJIKYUhB+vVb4/XYN6cVojEDgGrEfZEMZR+wZw
juVZst/W0pf82u5DK5J7snwI1lCxY+gZ2X7MOHiVZcrS3rhuoQeb4nJau+8qIwqH
bG4s4I449V0MuFuHTx3GcJuLDvwOJz9zObymxyGYqJ0axNBpMaHDP0ZUjrupjN5O
74a7dG88GivLWYgq6TF20loyCbj9E5qeAiSlWuTROhgEG8VCjUtNCzS9WnVhNhEQ
G5MkE1H+U7I7VV9j0ofTRhAkJcbo1+e1DzLJAyW8JsrJpouRem3HxaJlqK7EnOhl
nj/DIV/LGpkKKA7x5V8yF1ZWEhh+wUa4tQU1VFSxYc6o1gij3nmdC8WsG2woGKzB
s7waKTzNkmj+8vjLjRZpieoMlh227XzMJa1/N0xw13nbBGxJnynWD23gR9oU7rhO
oeG7kQQsxFx65JuyE6DGA/JLmr369BOxCJe+6cU8CjVV4HYo8WYWpNXzJMDJ7ORt
9AI8gH2kwjx2u7hA9eKXLrj0qgXcW270uYPfx5uEGD1unLSNHuWK4p2HproBx02R
dKSciGQEXmd0yoYF3qWDnxnuQer1p1UlFWs740gI4SwtBbxJQUca02VdIQnGL4vU
+yHNop5wn49dQs2/owBuYp/e8wH9FVqWpsy033Wj4qmwx5umDQ2q0JcCvIaHaGrY
5/FE5SL02FxaYQPiYOnUDSLra8XBF4Z9El6ZymJkmhvyL8iBC86gEClFfJJEvqi4
04lRoh+Ty7YMXfEZsOOGMJpSVLJo81gTrs1a2viIbXpw0o7/GiZQ/4FH8TIqUoIQ
lmi7UvcgMhmRcsoWJn0xn7uBhvy8SbIn5bWria19xmKqQVe3ab4tf3/mQA2yDCqU
/bLzhc/m404/4/yhi5aSFTCCrkLHNa/IqQdQw7mri3Cs3EGK0XURCVPRCDdJc8vs
Ch5TSId2ipLSxQU6eKSv+rUx5TTjIdBdFKfQ8Za6Lk4xB0Xrj1WE6yXAyhq+cT/Z
jl1yXXC+6IQRDfbQGFekvsDlkW637mvt1FZxJeIq0ZNT0ovlHjbTOGQcBenj/EOk
4C7wiAxs4LyFvG3GvhU21XLYYpgpnaihfAvUofy9a0lOqeXPzt8+aoXuY+6yo4Ei
sL1x19sWn1mLeV0WatQj7uPJ58ECMBcqcqHedv2LLqC3jRm+Y8d0AI5Ojh5tIdny
J9bB51dXWkk1d82uWdc7rqpjDfvSG318Z9iQGcCPwVBm7BXiVqbY5aRlaMonzO46
SWxtI7arMR4A5gafylgqyDF7eVY9f7c/D4bZ+/Kj2cr1//MKuvz8M2bNMaFFxPqG
/6sGRTmT+K5+oyNhCVPnJnpAdrs/+0bXeFrARGScEK0+JWGf+AWR/3UEgBfhPX26
hy2UkianvdVfCgjpfIZ8XCVveZEw9Fdg3+7+eYvsFYiPpizaLOOPShWi6sbi0EU0
FQmbSxHwF7vzQLQSa2SIqooegqbK5M1bTJ5aeKCZ2tpz0ji5jbcXnL1HTyZlZqFX
qkvuBe0tJfhH9xe3+3NGT9qD/JiRU3Supqi1tRAKk6GfaqyMBKi7U05e0dwnG30c
89QGOTc99E9xExpAw6OGtPjTE0JgNvfvkLNFc/n+nDvpl0L27vuBXroQZUk4h/5U
W/oyhHelu810bccrjNYePJK/0ZtwCbZEI6l+WvF+/UTBiaXfhBhUWTiy2i+8AkDx
nCcxV5kraysm4KXsG9/sTJ0i2DZEdUgGJKFwIxvWiyDoVsvLIJnI5nzFBdOUbExj
U/E4V2pc2kPu+cmdOLP6hd6wmRa56KNWqOZOazVFj8j+HDvOVGTyvlanb8Ml4vtC
KIdIOUZRyQedMh8BqQ2n7XF5oJmksZLXnUK2XCbXLmJgr5aTqDyDbr5GFFFCmgDr
SP9IkWFDxBkEXkRSZtBjSshvg6WSkiRB2gG8gwPHkcUeJpq2AJb1+wp1P8lcdli8
jx678wu3/UFwFdpaOlqRSIZoAVjvd3ZM5ERpXEIrb+tsu7ohoqFazkC3AK/gsZh8
8ml5Xjy09qdZtBjF8Fh0KnRP/ppxX7mZNnK2hJoQfxZXJPbxBA0/WQPCThF1YtPi
vySErS/W9P0wxcVs6RrEEzbXqo7J4jaeU7akcBT3It1awdjXFxkIKnCJK6bsvmSZ
UCWW51iy+USHnGa86p/16vDvYxop59wUYBe7Daymi5Dfo8gpnKokN+N6hfmQMG5M
hqLKcvSTWgLT1ePSaMbGT/hbY8RLMqxrKOH/G3Yzci5vHgyPOmR+kIY4dHH7dRqz
4wd/ZPu2QCOhisAFuDpDeS6gw7Xs233+ACdKf0ECaUCYPMOQiF1SymQuPcDaVya/
dOBNHLOoRqQnWcGHMlPi0Zb8BHoa7/JpumjKv+HKof28MprMR8VuD2i9NQ3bPFl+
qRrC8BjSaSFtT6PjnD8uqlrhwfJt6gWYneg5LILcFi+J2APMWB7YvQP+eVI873nx
51h4nk9l3kOvnPuKfvPS4GzcLah3MkpJs3csdgzlmANpWFYmRcou7jw04RsatK07
2+WTXyEYTA4l0jHpXGLa7hRRuCO6E6htP33vRh/fmfT8cpTM0WVOg/1ru7Wt3wbB
L1XnLJGQObG0TnP2AfKEl6imYzGZe5cyh9nCaVBLkpN5kYAZTl+MAmyJ9bZ89I7n
5B3lz1+a/Oe8sl4AhkZ/TfSZ4+RfW+pKtWSQcT7Bie85aWtUXxj91hWA4LziYTfu
YLW4kQRf5oYAp9juqCuRz2he6KhTU7SwA7RD8ok6Y4wL8TzB0lME7MCCh44+8nNO
SOQMPVgDzzMH/V+SHkxzz3R5qEhDkq6uvNnhlM0lyIi+yY4ygCXnmmvSe5EoaaEQ
7atVx1MvAJlBIxFqN0oI09MlGN7rosdCI2ZdTfl7J9Q06bVjrnZ/M8+zkrCBkNs2
GjGQJDw+yWnRmRo0eptvOh9IHo/C9YBuRc8sGyaR1PT091ypzIeWATn3SGi1rpSd
kxX6JS+IRCWfupgGbwedkNLTO0u30sFTapIEgU3P4oAPjY5t6/pWW25CWrXR6eVT
SD+ysR4SM7F+MorJueIhn9bOY39+Xg4Z+9DY1pV9XykbL5S0HUoIEv/ShBwdfLgC
jgDXxYPcLgk+sqDEWPivZ12wlimG9aUJrtZ7Am859umFVj5WNN24uFzTXwUNwBYy
d18/3zoy1I2rSmpjc76JFYETURnYohsW0Ca5mjGReZ5wp0yxdcxKmrYltWrggo/d
SkpYW56TOPUAbtE4lZhphtY0QWiBc1b2zpM2T908wodi6RDCin9fUmcSbna1lO09
2sCHkeVBZY6GQrJKBrI7b5MFP4gWHRnynbU5j3y9F+hu0y1mco0ywS3TVJH7IXHu
aOeLxMG8QsFomwpb7/Z28htl63uBFetgrvT+B3rOXob2i+aM4EIZpsA2+S+VUzIL
IOJtKSEZ+eMA8ta17wXhJlSbFGTnWUS/3MAaqr2xOUNrQ33sDeiG5OU/6aRSgTOF
SaHUrg6gdq8fPwBuTJzLPJ8OtatxU/cmngYXaul9068BLYJYnfoPi1YgYV7PBph3
cWGOnw511ciKt3pqxym51k2j9onhNN882gkENb5kqjCI9bcD0FdNt0jxAxLuSZHZ
grcgKXFWgG9E1s9SaxAjOPYNUBqZvHX4XwoUrusVRObplvZAxPdSJnIueK8RBZnN
tpP9qXa5owhy2pxdJ9avlaaD/Q5OM/pkM+G/xsXBtg8ZD+YB0+CNAzFXDVhP127t
bUY4fGgg52Bqs2uQanMp0qF95azhsdkyRdoWIIjAtz/DsItruDZjuGJH43Idycl5
rzr47+jVafiMIq7j6BngFvWzfyUYQ2JzxzsRka1fZihvyaLJJWdzsU42d5S1ZLGp
H0pisATG6XGyVocOVqShEPl6R5CRhPrvPYeAFiOrR7zMeNQ9vckQWTFsW+SxPiYd
/4VT3Tr1kBIThlxnqmVrUMKjXgP9V6CtUYFcra9oa+bir2sPJBPdjQxcJmWMfTYW
IWWeUvPttyh+Ds7J3VYXIbiTwgrR7lp/IhrNJGqeN4bkSoZQ2EcC46ZwpOj/wjBI
oGfoEQT3SZh/yihhgajmUkqEmci9s7XkyECGzWGVu8JYycE1ZN9c3JdklHob20z9
kA8U0z+fsfwXraIBmDdhwmScSMm4XUS3DvwT3iSRvBfyV5CEB4/H2uFBbFM73Jtc
y/F+Sq68Tqs0GwBDjMmDBySsA9WuneEt0xu6e+V+GqwoHF8jTrQ4ddegt00KlZB0
2lThHJ4iLBMBymqHFnVXddN9f+mi6+bb7xuaDOdHtpoLIvFP62XAi+xUpit+4PQs
Q5QlNL1ScW4kNvtua8qpTobhcB/lBCpjLGYbE/siOO/Z151DGku56GqhwtVuIqWN
9KCQeAWDLeZ0m/EjGG4vJxuxtJjgPwlmi00KC9QSncxjoNNjJk82tJaiuOI/eUX9
qId/V/MXO6jnEnIadecITkFBw3xtn+Vq5Ld68D7esrMzemcpEeMlG2Oo6NHcST5j
R3ueL8gMhs4U4qjqwu2GIwoG81X51B0834bu0RSeDzgz99H16dLAGVor2G/cDg3h
5X12C8gj1kQFhfD6NE4lAIoL584KONlw7fl0o6caioY1IjcrV2Cvpl3hS4boiM1T
NJwPAx/pmbDt/Jwzj01Tunudeq+kNhtpZPNll2uH7PaUlGgQXpnd2mmxgF/8o8mn
6a+oxivs52+EP7Kd17zKB7/hkbyUYUklJQQQlo7bv0nFWFtqaOAeB+2z3UrXuDnk
+V16p8Xe/OjmXrG9eG6oKiTNQ7pOga/p5P8VqfAa8tSlnPaGQSynDjXVj6P+wtSO
rbpdnfQ/lW0w7XaU2MWP5ylfh4WfxJx2Fo5OLBOgccbuPTBLkknoPBWTQiEFuFNC
bDfnNl2XKfUeC5hPwkdJImgntxhT0KJ37a3ZMtMTz4SPUyDUjQD1nXARFEuKWf8o
yzUpGDVt2U1bxVU7yCSnIG7uMFj3lfgy3pISzHmeIpp6eGoARcKvEYxPH/Hv++xa
w2qUkXkykCzjnfcvTWoHcPUshBovBuARoW5n92IMuS/wAGsCxbJ/J2SMIMjtgCrM
xqKm4il4EDpdf2yNz86oMsThJNNd0kHS/F4SEzpCIAaLdrdbaONN7z9mw6koWJri
LRXMg9Sb9qfJEXQXGmpcJPDKncTwNTy/thFSu04GEa8LVJjLnIEJyOQVGudb/sZC
t98K8GeuCWVwSb9XtYAXAp0o1appBKUAGV8gQuRNLtihtMBPAZ0hSspiyZ1c2iAg
L9XcjUqkxaJaij0MyJj11a1vIxSqOKfnKKLnzK7NDqz52FHaRzIWSK2jgEaj1lIi
hLiRbY55swPnau760cmr2AZur7uemZ2CZwc+YxVrxjD4D+KH+OcaSYRaYKtaXwF+
Y18Rne0Zs0JmQCpokzRWxHCDbFDyoJ0wSLUKQLZB2O3p7Wn37LQfolDZGU1PNkYU
4kUQhyCoqwGyksvl3GlPySXIZtr2+C6JLcWcYd87K5CP4yNnTvMJEfnUaik693zT
R6w9qIkJzR5hlXGP+ETpk/K9YlN/xGRt9E5w5vhgs0mOi7FQahbKhXaZmrLwhocU
zFjrCR1FpWvL+DZYTgzYVVW44bjaQ2zE39MRbCjsVcGFU3YymAlWlYIi9iGCr1vV
xuu8duQLsGfxr/D/EeeCe7Rip4FDhi06Xn+WICcwMNKQy9OddxWGOm1peOLAuEXy
nb1QAg5vwZhoenz69q0HJJvFZL03ThJ80ZaQdeDNDQCmBTfgzUX8IK+xk2I8cdpV
9oPb5fUnIALrBGatUDh/mpwE/vZo+ao90lyCPLjfRhM69ZsGBTEc9hXxVk8wGwCA
T4H0Sm+J2pE+MXbqr+7GA783I6CL0wNZGwRDTpVhX2ZAKVnexvTxLECUujFkq61n
tztqsSPap/Fvy6DxuBm5bUOI8KKcIKG9Xz/9/s0PyDMpjAkt9Tym/e/bK1Wp1M9Z
GHOzDoCGjNG8a7ylEMW2Fmv4QZp8/XnfwDpUEq7+ZeB14kiKvlLitRBnAsJtNFEt
XJ8p2NFuffqw7dgsrwLMTHpFLWb5c4eqSR4SJUmhckyIJ6a9RwpcmhM1V5L6aXtv
TD8PUv1xasTlw8XE7wenXksV8sOSshNSBrqLdy/0UPOmjadp/IUHtrqPdZ+YW9Mw
xu/GyBtmjL787g/yYFojZzEX9iWzGvqTxpKfSSvFzYspcHzpWN+GiEn7rYbBoS9I
yiTBl1HptliKxVviYa2hVOBIYmzDzqyFrxx7zhFMRIiLox9CRIsYC23V0f81CgKg
P24/r9QQ1tSpJHqA0KKiakv5TPnBn+/7C6cWbJ0qKQlEW81hqdTShIE/4Y/+jpI9
BZK1AIExF+RGTmq10qOYhcBx/+5WryOUpbu5yi+BkIOY913TNgYe+0gKbqp+VawC
YgbYNhKIgIHp0lkQ7lctYc8YYhxntsKaQzdnv5lFJ3GFUouYA/W00Gxi2TUxNwnQ
xwACMxhrYqEQUZ1YZLEgKrGTI3Agf926DKAPmOvSd8oIdWw0JKlicxv/l+GjDM1g
WXM0TFr9fyQhj1Dqx5m7S57yOchhJ9ZEg64kPJ/Ad4ni4aDa/inAUNTtFrzWUoVk
484b4lRs7Sp/CQgrBsxJ7jYkz1SU8ZvLTOk1wVU7cdS7Cf7NaFQwvSY6wrV4e0RK
hkuwz7HM9caJ/TyqS32U0NefLL8T1nLJcLphEY4/Zq/yZOiafuwVPErhrXwSKfar
3sjPZoStTvcAMT75vVhiUOtD3K0N6hqZP0eMxRPd1/YRq5P7MMQhGeQVS9yJrj+R
404mDxg68O95Cc8wukyUEKr1B0fpokLhqq6ctaIYDBt1ohLosZg/F30ZLC6iTo8S
SjQdwZwm6J8ScGVV/y1Jd12YPvgI+EIpfih9rSmMT4CSI8GoOzK/51O6TdECeLe8
s/Ucxjdrz11tXT677vq663IwvDSSyu/49Qg1SX3y2qS24Vk3Ek9cCU0gVIyUKYLC
q/jP0SOJ6A4sF6CtD1tVrsHfamEMdNtTcvlvOlEo4fG0w78zVoYNMXmklyA/C+xX
X4Ygu+AcnhI+MvjZ6uddwD/pypbH1g8lnNutbQY+Azi1+RzFzACGHDonr+efwVgz
JIbvTpL3YdiqAmvtpUvYxtAaTlyxK9EJpBfcxY7/byhdcMp6A7CQubijpqE/3lTl
HfsyH9a33dfcCI7H5MtR4WMYV1jMm3HN5wr6YoxgFCK4YnCrirFWIdTomWtHMKha
QtcEuE/SuLvqbFtp5+WRkII/iw4z43v92gDBIiD3jF+ldTGs9WYUm/PvqHZyKxle
KCRBYfbR4dc+0n8CF/KWUOo0IR+gW3/4X/B3coTHTPHdrL4BdDw+aq0JnnsaxIUC
STL42sf4nC5h2L+kkMPgtPgmFUMSmdzqeK//28Nxh5LfVnIx2/e7vCJNrIrLL2x4
S7YmLDQ92HGYGM+711XoYcxomQgixg8jRsLaKjRqphe8txiQsFF5pdnjTxD/ddHy
ybJTGXyxvZZfSCLdmcAkJyB47wdlkwj3aeKH5asXZqdCPqssQjdenyPW62pAx/CK
YY1+GnBgvrg0xEgmjL1rm+muaU9hDhQ5W2eaoFtnBZ2KyX8j6clt9U5oeldpk6+I
2v2/Rx2ewxADFBXZUfugl5kETM35F/O2gyqz7vq6V/mIxo3ZwnvZkAwdhvlGRWyQ
8yjt7ERpwHF4gD738YUc/P9f/N3noEVpOeMopIyBbNT8S0XsEBoCQ4O0j5xa7cDV
v8W8kvz3rqHfQ4gj4a30j5+s1ZCcnJYU1KCJso5Da1gudBWQfFxuPCzKDcTvY3lH
NE/dnT3TmepUsznz40eG0KhFBP3dCgqWcU9ThpD6GODPqnIJI9VylZ3L18PVBh6B
ctv9qtq6RxUbf6AEHA2RgkyTqr+XJdkWqpE4vejOl8d9O5LUIhyBaJXqvSjPUXNB
hlhiloumN1ccF9EenVhp53RXmpOKqmANlKoKTEybCbrixFscVJqKI2GSPvTzGQ2U
v3PAYhpWeLsJVG1phe/BSTCnRIdbiAQUPQzCSss4uHDJsaZQQpgF8ZwYDMRM9Cis
4mwuIvTUUIyq9KfDNoxiG0MWJFrKMcMkS1SEyD/s1YtGpg6XkYkXG6sUmBsHOg/H
U5qJvdzbc74DmtooVroDwom8lMOTIxHUCFwVBE/qJj1PKZQgUWIaSFNMDH4JNcY5
MUrj7yzBO5mh8J73NCjAECNCC5+jpVgkPOJUFp7mijiSl40v183yA46ZruOExcIR
NfN92/CQ1A1r3zLHmTBmfadF+yeNTqNPKy5Y7Z1NZkI3/EBTD9L4UZXdtzqt+ZyJ
dI2+99teIf7ZiNZgYCiAGNqFnYC4BAFG+ELIQOARx2V3/h+0/HmV9u48EBYGHdPT
jHMkNY3QoyMIp3l7VuexQOmXsu3hiu4h4NriPcoIzqLVKyI01b175QjiHa+PxGxi
z4RNmm+YwjWpbKzkYXhDh+EktwrXjSQeFinU8AmwpIK1w80ac/hvnfOieOOXLy+P
tnPennzf6Fra+sGw8QuDG4uy3FxgEIhQo+ga/ZPchI7Egvs4yZpHacJZFUEjSaJK
SMNl5M87pXWrv3EQ9S16uemPm52BWNAT39C0AWnZb7x76QXNspZLb09u+jXux46F
nVrnNhUuaAwSWphAF9/UvLEzyOb63IQ0WdJ6mH4mEzDFIkkI25FC7i3YujWJbqiW
08aSmO9uJ49eXy2YZ+a9co342kdIHf595v54HTCPeL1j22nOlThw68uO1NBNRNwY
mIePJNpElUN49tvXe14KyhJl9QS7I14zKr0nQfE2bolNKpUk3JWH1NOHprCZEfa9
WOfTWfnSLZxw59rc5V9PgLQO4IXdir4EkU7naoNSf3aM4kFncx04st/6Dj3j2kFB
BZLJ+XxkP7iScoBBZGSY1k2IrHiGxx3QUeHoV/Of6hNekW4UvONU4IRcEmWcacFb
cki3bxxlbc5VCfjmxGm3QOqOkPogbgMvw2WhjegMZ+Q/6s+6fNUu75af3w3qAojH
JciO8DdDrXylqAAcuKFQALzIowzolIxHsw6fWiVQYC82j2jtDgJW334qac5DcsYo
bchBrx8HfDPjJeIpdz5CmsuVHsHiNsP9wMm+TZgdUOXKw2x1RGg8VVbPPSNUxKqD
3BpN709Dyo3lGI4Cz43lnV7Oy+q/ZOzSciTssMV7Kpyk9jQZRwxNvDz3H6WvySBT
XUZ9Q67gJ6aQwLCfuSFFFT3Dw4NRUqBcSS6sAqOMQgYl+yd045otNCM520NemWPH
3LXhxbDqhNz6grW+uzaiWC/31mRZgv8Rl1zchv2sSxRcGI5pdlxuCJHrqUEMLAie
W47as8toK3yYH0Z88PVsvkm3JPOF8lKL+b8eBuAkvOy0Q2e5Vv91+c1miUS2RAt9
ZMEO1dogxpnFukmG9tQ56S2IPBwSUj4M8meo8mVkUHBpfwACw2aV9RibLjEoJUYj
ZncbBzPqbj11NFIqu/xB99pDi7f81VqITKsBT4vksiSIdBI9rW+fEyODN+zArzT3
GQbRpYpILSrTwIGZ/JLT1bfmb9cZcdgkVEe61A8D3mO9QWDOD0M3afxscXjodPwv
lGp/SruEgj1hQeTGfmEcHJZIR3VnyUNk4xFif/BHNShbvG1fidN2U2EA0hinx9BX
eN1yjgRY7RLUHJw/Lq58vVjoKHOCcLIZPQFoWN3mc1rvJwdmfkqB2t0iwiIccK4h
B9/BI+CDV/dteO034iOikN/iEw0iSLVCdX5wzl+fBu5J1iHLHaFVizxWeRdcIOaf
L1W0kBVIQ1KhkNvE6RE+/omdmjSEN70M76NQRrWUMkQW1duj/SfFI568LoP3GPTO
bGUwejJh/UP2PJL8hhFmpzhhzEpH0KDai9G5u8kPxH9EGl1me7yS0LzrepbgjV4d
e8fc8oasOuz4eCXhTypGhVynRzwxCUJLjYkvHx2WRtetWKSSlpaIs+Z/EBTjbecM
k34HGAlb+UhuY4AXYI0eQ2tdcWfv9bQcU1q+Ht4blhCasEAb0YKLfSvueA5Ajzt6
XzQo6ofqOzKcQtrbCdSXYG42LFShqRfAO7BaH3cHh/YID4S5M9JNRFpd597LWQci
M5nub0QyCERsxl5S+KeElR10lRGaAQ+IIfjct29YgWOAZ5UySInzPxz0T8v6E7My
voW6JCLqtV/bmOsmFDSiohNqxHDUr0GOUL1zN9rW+kqtVSMLXqd4hNJfH20wS7K+
Mk9KnCMHN3I09BXKmaNBk6ThTxfBC/e3HUBSQXullEdo1QEo7KgtsodbF1HnkFK3
6FbXbfZgN5Tr1fkIq1/Clb2CogaWJL5gs1f96mkdMo+c60N/UkM4+DwyhcHK28tY
83TxAt/j9Kp3TiDFXN+8L6Du3lu3gxGWT2cY6FZeDasHTo8Cn3OI5bKs8tBIbsQN
NIUP/qxqIP/2hayb1dXDEnuJIhqCfWNOGh3/l1r1sITX5+Z564ntH/FxKjo3jxOh
IMkj6SAmC+1+Es/pnHCeBDferGhTVlUFQXzXiFojXwcc+yHsttR+AKLHGfOVweV3
+H34zFtrr6I0QisYANEDAT3NRoHUodAhdAkQLFvkb/z4tdJRRvtelVQnY+GGd8PY
xIjHSdhlqtS2AAvOgmcZA0L4R2DX1ImMA+0Ir8z2rGhqrVjz8euj6FrWOvtROJ8t
y4+IlIVqxoMPz62EzWD9zwM1V2g2ZPZ6d60nW8jL01xE/TmVpIkrHRAIgWMOOBcE
T8c1V52C6VtTvaXnGBD9YXLAABm7bPCBrKvFEm9XzDl2+fLhSUTLCsGOGVInawMH
461BxpJHRShyc1jUKODKfB7YBuxREhnMQ2BqswPAjBYNTn67WlNh7Zvj/l4kV14S
p7T16KwGbTxOnOLFt00+IM0ql2aoeMYErhu+6Ynq4PebXIy6Pr8kyp8TkgGAbi6v
lgV0QfeBUp/sEVN3Udy5+0wNVhDUs2k9FhDRwehpINsIRSBTBdGuX66ctttzOAhT
9aArpqgJ0HKsXEqFIRvE7zacPKxbu1ecNstT27Scx2NBbL6zgrrdscSCqTzC/Tnk
gSIp3EYJqB+hgTpryLTidbfQtZAyDSNweRpUI+EgbtfdPpf75yRrRAPRoCcgFaad
HrkDOtitViYdEitqmyZX6XXsqKzhKdFjrjF+QMVnenQ3XkHXTzjeHzM0+Ahj+Fkx
+ALpiTd4ELjioqWXuyi6tc4nSx9lMLxGfKBhAbzJtHQDM3iMlEZXB1JLY3+ddEza
6WIeUHBkT7ZlENH+ct9eKkrp+WxTNtDlakiJ0XFbl4+QO/HDRHTRjd520Irui0ln
8Q68tPu7JKpGdF1ZY5CMewXdTWGURfk2y/R6w+sCmAMJlip2BTQ1WbOSovnN6ONX
eP9PTc32y17m3Ovu6OYe0GCpjydQcBfElbod6S0n/Os/P3gqLJPfM6xLxEW/BZ00
+B8MvklA6rB3LaC99mXDfTmSTrpGyX+imSnoi/v0+kmSVIvxfEG1JkgBvWSlUr7x
441lq8M4l67ncMhcDZK7/3t1BN2P0cnlX06oLEqc5EHFDfmLQv+rfv7j6xDNibkx
tIqqzoxqNeg2TnAI8wFFkFxve2FNSKylAiBcNzDrC4OeCg3iSjiCF3gqTIFLUbYQ
Mb0prkOS78yi+CAmiafmRMEKIPaoJmCm+J1x3p3x5YdZXJIsObnkE6q0sT4Z/CVm
INRWLBEsfmbD2dMUfYwiH3QaS8LvAyDZirsflCf54uXxh80QuTLoAat93GuBPhtb
D2gm6COag3W5WrjPy3+LgUaFNQXaL2qqz9EkhJT6mzBVqQVLb3GQXDvRYzyc7u2M
Tv3CfT+kG3QL4zFpzFLd7IfYGKysj1bxxVRu9BqY8j5BDSrexB1fRWTppzF3T1hz
hf6l8F2AiNKcDDNoJg4VA50s2DVLS/eaKobEMFpJ7yyM798L62KZZmLfh4t66e6S
XwQNR3h2P6hzF47+6VSilUtrjl1HXOYOhhVx9pPw7diDllpv5ake3DPwML+BwmjK
JIm9VOizOalp7C9G4RToK8X/eHLu5jiZ6zwlTVb/aP0KB/fVzuEYlElwDi1qOBjY
kn/QCbniJTmruUgMkouO+gcrhEs4dRqIBSvZFQKDFTftn0LYu8AbM8N6NssPjFTq
OwUkQbz8BI+tYmqMjNxVJ6+dMWDBEMYLct1SL07TDs5iztN9GPtZ+dvshHBdWUia
RDQqyDLCTfncjvtoYkcdLdd6wVFIqyS9SyxVVGzCkLbBL2UukryKvwefZVaoWtrd
GjbxQVlhJyy5aq/KlwMeytVrG8OISdpAE8NbdRpyHUJ9WK19+QgO3NnMkrzg6ddT
YWpKAuvwtL6nar/K/E4FBVPUjYlVU9JS60RtzeXL4Jx3Fdmjs4wWYYAznQ0K+1+D
JZDBIZT86z0FqTX3teNnq92zuZIpf1uzzguC3NLEOc2J4Sr8xFxs68wA+9SFlg9l
zOI49kKSiBy7hu7A1agMQrrEL+3a8cqKWB4JbFOV6jkEXLb5w02RIlZ2AbEKprEE
PslqW5/b+dMq0hOHiXMqO2rZRC4eELh6m6sv2Xr9MPidjYOCPq+FcdKV94MD10hO
doH7Z93FyHCpu/fiURRAdQPfxjmSbtwCri5uMIj2m/z8PXO1RN2KXt3vYnn4tRu8
cUxM8/C+OQn9pG48P+wvnsXLZkW5wxuVo0w+4YwWVHeo3CR6rzlSNgltZOasrczp
Y1Ekvck8+8mZ2WK9IhIVK191gLN/E1WWc244ahvPWqeAJYq3wOJOvSvsPN/58oHw
I0pzvFJWp0dZpxO11Ddhy5goPlJ3emnvcRet0PVtjMIRwBuMGsTUlIFt/0loLQOH
BhFYodOhY0X40tWjeGO0RwTbtJLq3eM1oBLnTLxFkpppgTeB6I4ZSMjTWyH3Nf/B
VWSTCmWA4eEOKz6nppUGO+D8QD9nRa062YTF9mwhiYwfALM1cESkwLNzvHINPLBu
6t1KuI+0fYr/IbvZmbHwQ931ndPWimmt/xo2cIALSRdaK9b2xHhDgybGGysU78up
nmD1Scl0NiNsVomWKu0b1bmWdlnNwVroH7kkbrZXWZOKYXm487FcY9ElJTNp1qpy
fD12khgpExWblYadUWFgTZwG8q0VZ/yZO6giNKQqvSx8jVuyMuuRhGQsxubR2lAN
w05RRXJw9gCGBcbi3saTsgm0pyBl2W1FoLXBgMA8d2fS9s5lwUO4M2IQMyoQoMjb
vD50sQ9IQYZGWijjL7hyh2qPDeBLEboNu4j1FEPou+lFhPF29KJ20F7ubisc26Kj
9uUdEfvkl8SzvA1ms1rBjs6WaaOiDmE+vRNbJg0RXKQOAubs1B1oklnOx1eDD6xu
yIaPbNvw/ZZW0foNoimB5KZM8O/AloCidcPHQKGhVzey8T10ahPFQcFdbguZJ/Ph
Jk87eW77uYfbojBHWv9oTOJhq3pf2z8xrjNw4J8cMffpNGYfdP1cNx4suDb3Fi7k
opLG5sPPF5Z5gsDNfNnTvx3RfUtv3SI0dekgHEiK9SbtJx+iUJ2ZZUeVnlVfBwWz
eMfXaL7fbOeXSa9pgpU8Rh6H/ZMbzuyCCuCY0ZF9ESHQiUVfOODUcLF4Q9mDUQdj
SCxUFeXj0yDBqnC0c1w548dDN41NofkwAiMCKs7iALocjGMvd07tjpdoGjiJLv4X
+dDAfYlVJc0tBmmFz2Y5Im59uDMFy01t0AJGgNPMrdeNZgqmboRX1CkCIkcmuaYs
tteS2o8K5IcVtVYtbkwYNpJDAf95j0H443khFC8Q97wfLvGydLNbO6L/+zrAduUp
UJ1lspGYIwC2kWNKYfSagu720Ps9pt3iRo/2w/s9G4Ej6WU1763DQHRSmwq8/TmO
QbJUsYQYlOUQCFWJ39mR6XszEILj4ca5ygWtiZM6iwNWuDB3R/BxlptOgcjCcmkt
Rn01Dxb4XqPGvpgXVnEIppRv9pjHaLTgzJGSWQDfdszHnxVhX1BRpRGAXM9VMQqV
CzPdS6ZoAKGKKmGALHX1GSewSe6WWN82aVk7ftNRdL6q1CZw26QPMVECj6hPNEHa
76sOZvCq2LYeCpURSriz7h/eTZFx/w9L/wAwKfPmSR1J/7T3gYhfcm1xvE+hrYQ2
nq8/M82m9tgBYZLs6cdc0pHQwPbyn4yaUIx+7iqU0TyVEtrPCuD5h7vKQXSEsmDS
AglRQ/GA3uuibYMibBq4NSt4WvUq55JuZXvgnQdrdoR5KrGE0jyDm8arTI6AlTxJ
NZEqS1vhFIkElmQG2ZmV9fD27BTA4COqrTHQ+nEuroYnEqsJuvEJuIScw/61BU1y
1rLuUBxjFJbvOiB3i42EK4CDO6ghQ99hU1PQLBQJDJdl2Av6K17Rltpwf0nFqGcP
6srvHTco/IrYGFNnxDlnAEfRv2SDPxqixsEzh8yw8yEDq6GScZ56taQh1gEWPooh
c6KlMJU8KgcDOURo8z/hn/s4Oob+G3YUYyWWQQp9krOyMSWrVyBgqq1L5kTOmsVj
I60FBfrEj4c7RqqFGuCqxRVZg+sFOIHBylLwBjhm50RkijSe9Zz3SiWIx3xoyLTu
JFzCRkuCnmyZUrTBHI5bsM82kOtvwbR/ATNpJCJulfoOd8Hwp7is4+9Rv1oVK3dY
E1bAtG8C5F7hPjulN83gRqp/is7M8ydtFeUL8lv+V+J726qZQ6lj495SpD8xJndZ
32td3JORibjaXY4kYppqozlNfKelQnSz8XjD9eIVZqyUwcnHJ4+DlksCDBXbFByu
Y+U7R7F7II9QbqB6HJaPr5AtCEWMyFJ5s0kENR0Se2ajNMP2PqCdBnopRv+J90gP
LoTDZVs545j3lDxHyC5By5X5HJEMZ974i8uu6TqqaO3KW26vJxlKOH10iH/L+RaQ
HLYMEZqGY2IckYGP02v48MIhDS712uG+AzXJ4SCVUyVX1Sx8lsA+EcsS7f6yT5eg
m87lJxmoxURpso2yRBoGHWkQuuE3hBD+QKmzfB3b0dWLxHPm4Lz2PKh3D3JqR2tY
BM8FpLhMtpjky7K359DCJBTKx6Qc5R976meQfMHrfZQl7Y+fevSipBhcNtSn7k2/
+pap/DF6Xx596vIlcDmlGb0o6AWVtYrt8rUKzr7h/agyK/LDMqgQXKWCZgKqCpuU
PILJij/hxU49grB4p25mXxGtMiGLRVByNg7ujE83XIa9joT3SngEs8Gx/pfuuMXQ
24D6hv4FSTd9fSEcMRnrJ0Jo1Cik8bcmhcarBiG6Py49BNCl8e6oVB7/Rh+Xo+F3
/oHAyHNFi4DgTYcqBwtjXuR/F2/oV+60gzJFDw8C7qEMYhD3reC/9ufQnVf4ttIy
am7xC3eC6ZH4ce1rEPZhc6e9OoZNnVVYieI3UB77DUTFYb5FasZ2NA2YfV28jqWA
MGe2d/IFUeMeT4CQHNFOkuY4Onn9MGgEVUoBJ63KNG6hm+glKV9k9TRh0CYJTzP8
UyJmGWkS3hAiZoOk/X3VKxNnurd1ts3JNYUo1qM8G3onVUzYw1HNXFmx7JipklgE
+m+SKzNfk4voDLAioRwAoZRL+1LHVOPR/wdsuwPCVollANRXdEDjPfOlomkWEa/T
+RvCQD8r83e+vj+6Y/+jQM7IN1JauLL/eGFYl8hguhHDc4ngsVV1geLaRyX8NPco
KIH1SbiGz6JSIfNt0zLf2yYJxIfQqc8vFojtgue0AzgRtRObwRQl8nTS8svLXKQM
hyhcpVjedQrJwGSs1LW+koUqFE3MtxD6q6TFBqY2KNo2kTUxUJTBSake/kPrY4wg
tnDK7WnbT/ePmdlPrQD1IilCPxYE5mMtTBaCby96V/xbb/YMv1o+eygydsGvSovd
09PrmzlGEBBdSeH8Gn/ZPsHb3RT9JopaPgTdlUKRCo++DHSyzzP5ScjsH/sSBr9J
JnBT+lPSDIkcN35g+HLmNzILO+O3jiXMpOcHHMgRCWmDb0E9TdXPlTycckk3MuPF
1g3Uz+vkWewavxIf6CiZPE4BX+JeJkG+Jj9Hi05Hu7qmQcoM4fQAZo0ksgbMF9PX
dpdYl8UWYCXp1E0rkN0Ah7/5c0BLconqv/OmxzYyETWKJJ7aSROCtTdkamTRDlnz
gNpEpY+ip0rJhEUgZ4I70YIpXeTEC7dpz+RUvJRUQJvIVj6wGs/AmJJDPtOueJcx
bL8+mVIUOmSZulX24bN11AW+GcNzrU7pWxO9/+YQdNH1DOQwjrQJ4R9i5+pYtE1l
RAzQ2tHhv+yYBL7gZoy7c094Bcym3VORczcvUTytAJewOi6PMeJpWMtcNGcTX74j
BTx6zE8WfxT3RusN4SizWUVBDkU8BO7jOrmUAv/T6jhnFkm8H7/dhdfogPjiKwcz
4s6ZkevWO6gtwpHKXtdboOCJsVWpLQ/RQON2WHaCFC0b0u9lXDKRXyK4DEhAaYnd
ZuKsSXX2uA+B3nMm4sLtUNzQckXyiQ1m2lEELfJjXpCxNV1c4aGw08im0q+BwEf4
Yu2ROHY8GSXayY+3s+3Hvr+GqXq2qXrTKUQVCFAjM6avkUUPKqWS/WcG9MvsnV/s
tevC0xDFJAggjBFxmgV9ag==
`protect END_PROTECTED
