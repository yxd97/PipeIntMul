`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xSzhWc8WwzPjG04/KrmnU2LokcLrgs2nFAYJSvEPej9scW3MhYk9tsADwmKop6jG
IvCa5qWE8b3yvAoulq3Qz3+c2SBUPafwmLr/QPOh5VU3ItNy8wFeOGbjp9T04Nkn
EvvBwZx9B9AxA2wgSIMHGNu0pLd62PY14a+98fdIKgb/FdJc4d2gUfYs2zouPlyx
UjLaSzDyBQCNIjsz9NIgnkGTQ8JPcUjIM15XYpfJh3PqbMFKEmxXsBTNURJYV54c
s1z3Zo0e3mNdx/A5QNpoTg==
`protect END_PROTECTED
