`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+/ri435J2Wf1zl2h7zZ8iZ95qJL6N7kvxFRlo7baLzDCQXMgtA8ZVG98bhDDMUlT
7Pl3qVXg2vVPkMUAkciULMqBpEWM0hF+BKp0t8dMxY7qL9dXqx/pTK8exDWnG+L4
1s71dfaMHJgPNFRbGUaKrbIZrmJbX6z6gfJdxYDt/GSrOfPEJ4SXU6QGV6H+IGST
huLE9KL5STbO6iNWpSNFs3Vjhs/aaPoXHreSjJokoPY3DrLETxsjpfjTNHIfIF+u
ved+lWSZcQk704JUByfVgHV8R93KnbLvdh/n6cKuqQdxGR+siiFhIli9YPmZ8foB
tfnj4XjptbgLTe+o0sPaewj8N9V5kgVg9H/a9Wd6/jjDd/Gbi7tXml3LEDg8KHK3
RIR8NZ+pRxBk+pBX8q3JrjRzBBMm/PvATLbn1t4Ps55tCL0/wMAIArggxGyruFg5
cly5uCZKTyom3/3hxCtNdRExX+4cD9r3jreqRZxzNg0NAOwz41zsYVVojnrK0NsE
4srCN1rzIp46JHofTC10Gg==
`protect END_PROTECTED
