`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JY/k2dVqVZyOYgmJqucoUtg2cKVExLhKN6ki5AkLFYi+c+bWgUSPM7XcpePC5FNv
RVou1WkgiYEPtp/N4h0qPQDVO8evfRaUvyCwVCR72CycUwHZlV6juXqM2wGR/Bie
1+VU02u97yQVpgKm655C3+ZCg2AXET4gQ2WfC2dmQbDo5lI+oTfBQc6IJPt/GC5L
ujXvkdHtTUqCUngwSYeN0/LJDZoUYBSjVlywcvkNIzcX4yVTgsSZOrK9qORvq7z9
w+Y63D7hhPdK2bXISgPbPJW8hXNi5TNE/MnPY6xWy9IQdzI9KXttBE+Xen0hNCdh
NfoZkdQR3DMJH77UfGf+FZPSSxRGB8MPSNFgRzcUeUvAtobt5JxZaMDd/3VRbNvX
qOrmAGwQutyrNyK51M2AhkBId5DEBdAchmLG3msmIRMkGfCKg0USes1O+t606la+
fQ4JeoD2XmW7w9jOAJloajiB5rCmyuAfIQ8p9C8e7OMi1OnxnQwMvdJ051wgy1y3
7LeyuLor/u7GxaVwC1M2yjU3S1AXwEea6d0vv6pz5HOva5B1WcypOROd5gVgHDn8
ZM22hFJAKIV6deuVv4LUbn/JkJ1DaltKN8aus7wy6nIRojDp7/4bwTpSxSPDUjuJ
8xRwpephufb9xmIF8XAtWaupfwr6/Wtg8hPMyspuIKOWSJQEaGxBO25g5wx8BEl0
EW3s7eLAgbKxu6sVBirm5xAio8CLOy2cgpMGcHFOPO4MxCy0U0r3TaOz5g1jVMwW
eIuuuhIyyGG+oxeOjnHANHhs7wyapjDNSDhtEReMEhO6LOT2TunSd0tXp87gggsf
goS4dwgT45pnYmRf8ppUAELiAIA3pyyKY5MRT3jMVNCnz461u7BQ7arQwbBe1yHk
`protect END_PROTECTED
