`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tXZ01SqcaQ8TIw3n5jlySa/1k8rjd6zOpardpOZBA5sMCYMgNB0NK+0MY1RZ4CT
jrbAilRoMMK0dmpX4FUlDn4WrT/D4OJM7dB4zjgXQNSgt36kN9WlWQGR8//JshPN
K7MfAF6h78HxGXkMY7PwidXyDhUKsoaLAAnKFhBaI5lAHnTOZltW+ZaOvWHVsESJ
2E8815Ea93r3xHQ3cAAvSRgw9vtP37gEclv53xs7eAXsDKqFE/pAiS/Z3uq2aCCb
53/UgkDTrTCUUJWmnoy34awr5fxpdIXKYud9mXoWLfAwcLbewNOnRZq1+3mEEFED
77Kmo1aOAhtgCGjkNn3RDm+N++5PW1002Swx4gwAAjTmS5vKwwsm/J7KHsPf+zh3
ink2CVrXt9mbYWO2W45XwpjXe87RiFlQiJxqzqy3G+++gU+mJfp+6BmHPY4VUGwb
vQgHbrfLelsgCyQ/sRjBLVk6SvUcO4cdmOT7Y+ysv0b/vw7CFktzyOW5I5TWuEPx
DX+5okasDHDW5Dv8gvDkY/mGu+LbH9dqffSJDQNCO1sUDfNTv77GqQnK2SlDd8Md
8M7ap/g8Clw5onZlEe43jtSc3ZuwnKhMRB7RHgcBy4ns5rZ5GHlkgHiVwX1EugiQ
c48BjmhuavAzNg9B6es5qkIhkeHy1xaQxlfljkdqsiVSRTuFLY//dRZAZAAA0MoX
uBza9n3W9d9AM852X71WU2Fg/GZg6Un3OtPQF+22B7UhvSBY1a8BsO01NqqRnBd4
/ZBwp/MV+DWIVNX1bfU22mX8h/pSVEHw5/fXwGmfh6LPhgW5pPzhWZlSmezxH8tx
vBSJFJw7r+/Ehzpu+qhJhM7XjZuAXEBKUXtV5I742M5LFTpo7toE9RD53dwKXmra
seS50ZzFW5kttrUmmaYi+sfWP9vMn2QR1POXtH1B4pATtgIeDFfYIOjNSTOFIjrr
eIibqJTnkZJxSPaya0BWP1/8oogbmjxrS58sch+GgOqZ7OJFJr0R5XSm5cKZ+XG1
HSnL+GU/iAE347VsNFUs0U76pRmSiO/MPjNySFwhTq3yi2TNnDDJ9ufaA5hcz0wl
hs6U5Ffq1AolBITu4DlBf1LxMVrvYE0IiUBAynbqODhDQ8HOCj06oScbL+6KNhZz
MTLqiR4Mr7IMZuPfz8gqww==
`protect END_PROTECTED
