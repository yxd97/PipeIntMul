`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GwxXnPIx8nnownIFuU5TxiyH/jWQAte3vgxgMa4wZ62QBm0VKyY8CWH0+HJMgc7o
Im7G1FNnrE0E7jucFV3DiFtp+UNjP0uc8C3NLMl3dLf6N0T866jirKDKsp4Zw8GH
N5mJ8tqJNNYLS3BUSIC6C2iESLszo2leErovWUGD4ixGHlmGen2nzoG29FJ1p3FG
WTpxZmoJsokRkTrsjTIYwAq585qbmPdIV3c4y7j2qEVRnhGotCdSFX+NZSMQUKCB
n9Fod7ohWVcXZ6dXIFLRLBRhQ/JBkaANXc2TveyPfigy7Io64PQglTpVxBXukVJP
Y8Ecallb4jndXig36unZr/cdBiEQDXayYnptyuW0jWt32haeZr+vwfC9+HdBZ6vI
rmiK0YO/6D9yHjWcBiOc+kDslMbJnfaOnnK6zDSSVTUE1qGlPXO6tYi8YZpgCpVi
zIHs9TlTA6l3lawL9KU5Nps7rQf/nMg58twMB4fIX9Vu4/kCpPZv35+caUk8FzIG
3TNh7Mg+mKNcCiMRqpEQJDI+2tOOPSI9WsbS0yCwYqzXWFQiDPAY2ymCOIU7vqw7
Yh4oU/Ug8bTEEQ7Fisf4vIlD1gKWEX/mzulZXOprHGw7juJUqB85FBRwglTkUFoJ
PdwDQ6anOkv5ay1SQx+9fGt/QsmBymhK/q34+IbCcC+o0xKE2z/7DF2A+9qgqzeq
ibn4bNASaHnW3fRG5fUv3HfRnPvALwKj56qfNQz1mwoTvDBwjBNFSzMfdSA+2flt
PzFyu4u7wGqWSMZCfJGvj1UAyKFOm7CQ1ZNJ8Jj2tlYCF3V4fC5r6ktGfgYHg9aN
j/Wm1fxyk7bB+ZXyw3Hiu/fsfb9eJ/o8Bqu4v0+QGgS/uXFIPWFZWxi3w4pBVsB4
JRTma1mDGR4qzQkmsyk5TGchkii5UKiF2gsYYbhEncUzRd6URI1KjTGzlcACq25L
J6La4yHfE3n8SHpbSb15QvzQWIwKjgrzVoxrBta7h+wSvjcqAWT1EKQss2Qgq3C4
VvoNo/SbK5G/ZU8WYbokTBtbiWkwdI1UKYafVxDaXh0teGgPeQrEbY8ApF+FbvFO
QmG2ZMhY38bgPgsx7WyKbBx4F1NzMsaWapqE8rE48Eg=
`protect END_PROTECTED
