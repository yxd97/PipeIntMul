`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBewq2lw+tKTlclKMkbZGvOcWz4Dum8KJ3nB2Ho0I/icwIcNZ4as1PB8lGSR5v8D
irHOWwXblvwCD4Qbw60Z3vm3AZq3RpSOk8Dbx1bNYrd21kARwuiLJeoSH2pECN3h
W5T9yXIGBZmNSWWhsnanm+NZL7RGobJjGn1mqhhmsWQNAEfH2QVTuzsnPyaUPsF/
aqlhn9L7vUlYt54VZqRyQqFuy/kSj5pWkIE8lzVesSAEtdtq1yB222uFpCCC3i3g
pS20mj6/BpMBLG4WI74extNlzi6BweX8G/ZSWVBpKqght2ZXlWlRRvQCmC6FU1Gl
6IwNmVqNSSDjJexW4Yyr2QTgbp53y4WkAYQOUErjZXFk3Pc3gWL/7k/J0b/nbH+8
+bmkSgHhb5Wsr2uRIx8rXAA7xyOgW2Xb2Y6XPkHmODvdKyCkdrqzJ64U+Hjjlwch
2ObFcoiMevHnMzNg9g8dGGsBX3rPF6QSjVb0vANwwEK8L/zafyb8SVTnf3uAneQ4
/0SxiBfabr5kmHaJ4+n6ew==
`protect END_PROTECTED
