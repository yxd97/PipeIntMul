`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7JBzldIPNnrP0XlP4Aq0B2r9UF0Q+GHNYH+wPX2EZQWfUCGvdbkGnHxrtY9RVvJu
2TJt+wJwgyrwyx9G+5pUox/U+EFqzunAogEvRJa3uQ1VriI+rDoQnf+hbudJYcce
STLegq4WZBq/7wvEKVBkt5a1nE4jIWP4vq4LD9hwjtxuYvO3PPuH9KShVS2iJyjF
FUxiKUrWWeko9tCqnTgmdq+d5JG2/niVNYquK+/yHqXvRvJdIXNrDWQeka9SQn90
2726HrIpCArgPgWVXw7PTjVbFCzwLl6D8Z23iJNrR6rrm4nXFgV1zvY5toBCBKW0
f7D8wNC2FZZX7IaHhqRr6OWxuAipRXRS19j+puvwlVeI1FI6v/aG6S/NR48IrgX5
OpG+NeJyrsnPrqn3xGwIUQtvPVhof6lbwNOakH5RqKoobUjMsJhodGPQo8pWcv3U
BU3hfS7AlLVcVL9KmrFxJ9ZMbRUYNvVcvGoHoFrtHfS/mRGo4ZBXHYwNnX8aEaXj
6PqqEsqjEYDsU+VZEm+IlWIR607f6ED7/8jJbv2KHizhrPSQY6Lo0iwlKyYWLnxj
EA6TOCdtZ3uFB29+azvXCWXbKg0k98QlQyK1OovX/SQ=
`protect END_PROTECTED
