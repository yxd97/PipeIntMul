`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3B01jShm3KqKD5P2mOYSpt1+PMGEYKzaV3wKFv3q2TdM0l9OwmL4eLOxaw38JUU
KioFRrUcvc44uNm8Ezghidnvsmk6q4blz8jlxUSwS1t0DAzGdoNjP+Z/JpJvR5h2
mVuBjaoGicEQaMUf8xQHgVHPW/OtoT2Xx+d3ULsaqh5p/2BTkhxrRTargCkD73ei
XeXrcqMjptNouq17B1gnJ5waQvEbhbzN7jWSlC1XVWzUoJ6CmAXTMzdwMoOwY7jL
jcsjvD7/7v2QuIPOeV8S7LbmrjFE5huC65zDAniSa7FEvNyXlUZvPGCUubM5YL5n
5Zao9DL7SEUROz6wbHKNUGD57bYBuXMqykAhoKgdbl3U7E0qIj1YARiI3Kasb0zL
KYeirUHShdSIyOhD0ZFk4lkQyk2ZO/Gheh2SCnUYKx5AJsRk2DiNHbAyoTk+OKZi
tP+uMshMcdz+a9iuruDMfvuYwS+5YAR1ze32eS87+LW3CGZKnT/ZVRvEFc3ArTT2
T60XZ9TyGTZj92mld8QRibhADdcl/XFEgXCXqhKCYAJGsHOgvVatS4g2P+KYqauV
JtikEghfGK6MeBbCzs8KCyOe0rVVMPTlkfCtsT6joocCYF2LViVCc/Licdfv+fJ0
cgYddgUeWwOi1jE+KimMPfMY1bhhX+DArnVHIre1Kc8qcxL2T8JG/Df99wNyqNYi
paSk78idoXvSfu/3xl0+zF6rhIfR7vOR8rJ+mVZKJ1khNzUyNR5Jj0SaN8nvkGaH
HONuOX03+Gobywew+bNKhJ0AVFuRmsX8nGXF+abbXhtSB/nSfNQPxiekFfNdjzTD
rdyYLNP1FLDGJq0KOM16YT9QLH9XbHajzqY0T8hcbm6cm7xZEvGJqvubLztSa4wS
LAC34oHzN5li3v3WsrRGDAHPk5UUCOrUfYnhiSxB5G1eHpfsQoI12aDQ53FpVM41
Z73D7SUeUP16qgw+NpW/MpfD30C+7E3uE9L1hG8htNcH/5M4zc/9/L7QjYTOZ6pQ
NqfnDEfWM0WnrPMN2RlA8DqKNqxVy7AVr9eTnc6VOca1EFGJAUuTEH0ZPVRWX0hw
Lrmf4lvHM+tX1pBdnTn0O6pmca+PnkmiD/nJWaDwFBCz+fdBWbYQ3u13L3jDjmGE
9r7W/xjFTtOOy+ABXJzKO4cKCr7h3d5SMvhRp9QwMSSJCr2BrltKfKPV6rzS27k5
Rkd6MY8ttBWT4wB7O5QdqmI+eoEE55tCDosQegR3GiA5WhyiwLUbdLC+z0H2fphk
df7xDblzB2ReahL9cKk3UBlD6R5CA8V7xykYCe4XhBxFMMon1vUVwVDbfVygZKQw
LXk3Qbsd8DGNOCUcsB96MGCddkEW3qkx7wp5anSyAFcne7iQ9YLr538oTe7xxodR
AX+ENskLEnOqIM6LkwkPgFAc+T37rlxaEBKuxCVFVP7Jolc5ZPGkViVdyOcNoKwo
p4OrG4USzohCLWPDbGyBlEnBQigpIjrxEAiXQ97kRAho+cwMOZIdi+8lMY3ihDkB
Qhxjr/EMSWlHqjvwLuqP36Q7hLwRDrY1bj4bhNkzFOG3es6c2itNUwR7HjOIGVx8
AZHL464kYoFUIErVz54G2zWhQ6L8erJyZm2LZ0MJxb/m98rksmw1/6shRRh/aGZR
sjhqV49SIIwd069M4z+kXl4LfOLTTIhLWCYEExMr3sRR+He/VBXj8re+rD1sBQFH
2LwXkj1/bkh3MdfBd26FqmlqKGy4stZk/zirGBGnkgg=
`protect END_PROTECTED
