`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iL7PzwxlNJISJkk69awO8F/S+ktXvmMstzXga5mvfxK6DqgWJJ20hcN94HEgzuxc
16xTw1lZED3Hte2YLKG5Y7ZyCrpR948r/iECj3zZUskLS+dZR3JBWwlYYxo+VrqG
pNJS7ibd8k/XlcyOuYcZITiivtXdk/9x4pdTL/WZaYOVat82Umb95qhheWjxjedq
DnOg/jUmHM0LMlMBLve1DiVznoE1tt6yS5nHNlReSQ6EZmNLGkcCFengYQW+QA5C
+mv4D/KJS5C4K5OqBSUx0wFtWSXA/vvvYYaGGQB99bXA1AZ4W4zMBst+9vsWgEr0
GN5V8KVfPFPWfK1FKUTNDZFxOa18f9m6LopULkR0dEE9ZzHFwrIkLugW1IB49RjN
MsFih8m7D27UnlBbYA5lk+36UDbqorjuIJdfeiA9I+uGJfA6T2AkCmzzhcg546hE
XwpywZ2vaOfTbzApyjFjWAwmfdCZ3ovWYQjHkGRZsi5hTV2W3ZYdBlnGVqL0c5Fw
5XZeYsnu5k1wy2fYXXRq/xkFPhEXESM/njaBjmIYgsV3Dqx3zNLxmKPO7hXFvIXV
R2Cl7HME65Zwnss/9I+1qbBbFrtBx0wr4P8F19kk7N32OJUVA5mzCL1hMXUXW5XP
xDFlyyy349GzOqnG8D+Smrq2vSibO49TwY5lpZbFQr61hTFh7lx1O+2k5DMwo2Pf
Sd1S2JjP0SSPcPyEDhDeyu6ek0hIRV2vpHXgsha3Kl8NitVV4dMZCLKdehoPrar1
M7xHfDrhTGOL3+pWIuTCstB2M4gKUOyoz+Ye9c2oOMtqU+29t3R1Xhkx4h5CWaU/
yMvbD8Lvwbutvo38mPRw21DHuA9vHqY5JpaVdlEMNlS7/lWcdfhcXyF5u1zRZM04
jYXWMa7nxLaY2nih1ooJLYQDfskfe1PGtv+PTKNLh1A7wgkAYtQ/0rHJBT16aXc5
qJec1Kp1fJDqgwfWWxODwLq7BgLZldsmqCDW/kBZruGYiCcUgeOPZcNQwcl5PSlS
CDpQ0SFVLz0e1YGZCwHPxthh7qK6ycCnEFy4EvD9Py21N9J6dNMKduOcAdU1r44R
0SnEtR179wGlMlsBnp+8R+2MLGqeD8gqZZe4U0VzyLmJ/Z2oRZuB0TJp51PMWaXO
bZEEuSEZByBvHmD100F8FMZDtn+92GmpNcII4QLWGyjjZiINruPCf4xmlAA/ZYQv
Hypor7BqIN1iI6V1tSFJpNJUH7CWsBUhtCn80NPVIFIN6SXcKRjjGengLj37vHQC
Aph/68u4COmM6NAVMp5KDkYfvnOymXuLoX8WJmbZHjuibIdIRsy8HR77nrr6RaFR
VSnXbuQv5vpv0s9SHGSNDDrV7n/Sa5vWkPCCg+5QwVfuYNk8m/Rr5TQwNRXdc8Js
`protect END_PROTECTED
