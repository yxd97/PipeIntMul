`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEkJuJCf2zNZK02sJ1hqNRq7rbB1QehXgY6GgrqufX50TCExm06NpeojbMoBDC01
olZIcPiR9YUSxtHRTcn6/+fE/5N6ipZHGkFaQ9XQkSDrg/3/LqbvJ3jb4kBBAYHR
4MrKv/wFu7Z+/ZxBB+R3iop0G0ROnWn8VTiCuUB76qG5YdnjOsyf8qBbSGvbFK7D
0w6b590yTUWbK1zCQqHVeB7ZPqQBKGLvN2hJ5FLO3hY2lBW5uCpHA5I1K3XJT2rV
O3PhByIz/IRJ+TTpA39woReULzdiIFW91g1YTHaCEHBYee7NbxUiLcs+gzwAF2Dk
OkG3iNWEy/9W5oqKXS8s39OiOT61H2GgWzPYdS3FH1DL6HNyfUmiklhDlQ7N4XK4
oP7Jb9FUggb0E/TAWLCKLQPLD/dmTYgi++Pa5zaki3qeC+PfsbwjbNXSf7NahlfP
cdGFW46/Bfc2MzQlOyjH/EiXyl29BbaC8y6De+VRlHplXVtv7X2KnHP5gWyBRcgM
QMglYcT+JcHlZ2HkH5Owt/caMEBJRKa13BS1rpK4CMHHXwTOIzXya4+2F+i8Ux3O
b5xz6KHSzUzP0ULYC42qreQqkoqkfospGAO3vO2DcQ1M71NIQr6RGFTVwKhC08Ay
fxHgNZt86X1BNaBjsmNQjE5Dssr0cft4qpmboGdCYFhhJICrXseiripkD5lMmjUz
DrkW3M4/61gR2NeDvLyR55MrB8Xk/drXJEDLV3hve++FSO+VGHIU7FRbG+0wxT2S
lapXVD+cjWM0RldPJCF38KnaivALVYCpyu/+K6lLICpUmn+AIgsxOAaCbV1i8jj1
lUAcPKpkZ1rwZHCq8yYvRb4yeLmOBDrFIDu/IotBTqqys1JLb5gp+zyjoNRJKXsl
q/vpsU/579tAVReEFrdbOGkl6eXpiM2mf+nr2M7O3SF7D91s5EpHEgPgWhhXh7/x
MmAcovIDhJOmWhzOgsciyrTQd0eq1Gat0qgkd9vpDa/sCaz6w/KZJr8CrqO8VGJI
juhSPp3I2Hcj5EEGfONy5y/ZTkkBGiNcR/M60xoQYoyQ0YqBDjxBGUqznmVaJxbx
xyDhp1dXSKm0tj1trz2HZKvKYQk8gkkWCUsKpeQfohgPzMQBCZhGyGdpcX2bOLpv
`protect END_PROTECTED
