`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vd7LcAe1n7BhimsguafSrJd25FNB5b2fZuzz3HuU5EO7snwBaJtdJv3a+yYv1drm
N+jGqMIwMvZA8A8z1cskNX+5TP2iLLmt2jr6DewQeqDsybD6TN4u0PRQMq6eSFCz
e2mOOhPZQxxIzELUkMcXNLppbVkPEnWL6ZTg3ILS78q6goPXnOd3EGocbbXE+TfL
I2VxDDS6B1w6Q+xcj+oXxE1uBFdllTca1tTn2k+8LXaEiqxs7Jj1MxiqrehisSis
1CrPFHosmtjH2k+Y72Kf85LsDRvR+K7WfwcKEWX8FiAPHcg9j7ku7A9FlL/n5sr3
k/J3W6xfAB6btFSydVAlWULj46My3jWXNnGjYXOMu/1QWRrR9TJkrABH0GrxVPVS
BhycM52Ue156YwKH1iorriK5gxMMJA7DJZaT4NItLhF4s2M630KBAcPU+lm2KnHs
kzJwzDjtleOSrWpxPGrNIsmBDpIy+8kLrIb+M+sY0kCWoON7PrzMfuzJ1C49cqsg
JUNtjDLjz8C938zjWP9EEQqwhDipqVO5b6q0hDikziFsw06a4rJW/6XH3f1+pH04
y/z6depQ4Jl/ldFWz9dDxfRsKNqyXPqcZbhD7Izf8moG7luVCyywVnmaSzx/xfT9
aRg4VgkmxQJxg7rT+w4fMiMBJENxe8nK9bYElmG+sJFxRgq8S0punvSNKx6D3kO7
91ryIBKXBY492l7oN0XSWlBvLUhLDGWpVEPblqc0SPQ=
`protect END_PROTECTED
