`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YHGWbPpMje7g8XZhY1LRE/SmbAZ6YbU8umt5xqyJ7Gk4pTFv5Su405PcOq8pq9pU
n+rL3FNcAdKTkXE0Pe6OtKm/NbcF58f5rUFKi8chBfZnhv4jREhOrexPpS3wSsHy
hY+KjwAHI/HAuq79SzVsEmegXI0+hap+aMHSy5wt71ecElajmHRdxQdRb2FWs9rn
2A7k8HwI3ePRJKEwPWTty1BVam0Y7otj1vOx4/KGgk7QKNPtSXTJh3OjXmTN9s7J
1kW2HvkJfaMZREZJ1rN4CfTSenisSGWREQ5oga6XX1kHtQNzrFtKNENWV2aB26zC
+StviLUksXtnBgx1o+0Ou4jBsEzLIY7xthfJWpja76bKc7a4c4xbpfyjPoe132yi
G+W5ZyOTffUXiL/P0v7lz4fJEYUtsfAVA4gtnfSfrUVIsf1PFh6uCvAxv/KowwbK
RNZWelqV6MJ25SNXnrh0kmdquljsVnQXLxs7lxc9qwRAtpRPJ2jRz3OUYcKTjFRh
hsackKKcKQhSXAw9ZKxJ2ojqF7GypPCEFxiVxMj54k7okL6N+U3VU0Y/mXPexxZO
r2LOI91E7q5gw/KvEkFdVm8G6/yS0aVySG4/+Cnl/hUQ2qf1DfUteqTo8kAAkynu
DksAs76oUzIV3ldmTge/oVqVdWrZ0ExXthHJVDrz3zYH0KpxIbgkZ/3kGir4DKDj
l4MO5OTev9eAvzFVJLId6g7LhUtdSxrcXBzTeo8tcK6GS77Fp+5QpK1GbQZOcsXB
q2lbxJdzFnxUi7BDSUzNcg==
`protect END_PROTECTED
