`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WHFKlMCzOVOpXFpnlP67qYflesG/suEhJZIK3Lv3PIw13++s2B5S4njykmkSapfm
/626vhe3EglHnC4mVDrVhFWLLFCn6en/7BjgFrHQ8ebClkc9xulFgPVX1KAS9Eh4
LazdektG4o2mrRhCP2mP7xPQ8JDQRGIpiWk+UoONTqUHhdG4DhEsNooRuW238Ziu
x+ca1Dvrz8pbLQ05g20j7zq0yGPD+9qZSpjvCajidsZxLQ0YRYINSTbltJHWJuz1
UtV5xIiM9JRhmDwM4LfVH1F8NsRqG3TD/mUXXQxKt8vMvuUJKU3eRJKBvxynFkl6
WKyfrTFhwLBh8ma19ja6PA==
`protect END_PROTECTED
