`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nnc3cyp7Qp2eythhSuGdLCQEIsKLugdHEGxYbj997eByhe4EGc+oeCh2wg24zELm
M9ggxApTKLCk5gm3Cl1dgh4JrTVNbDYvNqcNs8PRChzsEJCKBUoJvCZF6AoTOCUj
+eNLByDZwR5d7hBUfeuhjCtOUXrJ9DBrmC4pVTwosdeF448ehQTrhJbTjZRSoxMy
3oODpKWVO3f/a3BpJvD6n0hv3V9UruyHbexiF6IcK29HwiVZ3/SJbdnwi8meT6WB
4UnHi58+IXus9Y7zuWJKf2WjwtPo9BSw/7Vf5iIZ784ougDnI0cVpQeIQkwEBBGS
92gC1W4t75u+PwpSbs38jHd5R1Lg+B+atSMqDjJQBwXfmT6HLpe4z5DKfHz9Y5fO
PJGsQbBtCDW7jfGn1hIukp9KYb3Q+OXd6QiWOaG1fxbrU4oH4jBIvGd9YOjY4EBt
qNRzKqlTs1geCDkk7QGJq/IFu7wJC8TUx7xYBMdu9U7MAkFIXr49osEGsepYk9Q5
9uWalDSTxIhGYU8wMpUFpHnOoY5WOkpJeNX7T+3E4YOd1S50QsBLZDNM3LmoIWjn
`protect END_PROTECTED
