`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5ZaOM3x++ViijoCHxgt/4wfMhx/2XbWjttS1FJ9SBSKbEMMhCHEUL/d8Ou+48uk
qYk3Kw5udqfs7992T/g6EoUO3zDHbSpjpWiPAIGKo+l/rl68cOuI6g5/C8k1s+pp
2BHgPcRIRI+feXcTHNGfUtAXP/lxS4/+bA2qM5KhE4Uli6UFbJVvmLKCa81TW4N1
sa2IPd36Ke2SeLWvxXoP0g7+UJaFkwjTmBvvT2A6vtfcQdGigRn74zcekCCbimFr
C8CXXrCDpxpnQsZ7pkrep9y1/F4GJ8cTDgZCq6DC6MiNRDDVe98ny77nCiv4sTi3
VRhYHiqw2Xj/OA6H0RxqyT3jrt7znaEbNrvGRlZWKADcxvAP48csVvTWQc3pys6Z
1ytaOda9MB5ywID4BvaV8nXQgU51Eiulqrda5kE1xdxb414Goxc8Emil32RVPVfU
tTXbvETDeilXzzL2YwBfo2NNnWKZ4LgMvqejP9oOTQ73msOvyW9slNfEc16Yffgk
+0dz0AppkRjKluLtWNghLqhYDNwCPtcfuRyZ2R+6G/tL704Anhzooy2OhPNT8gE5
9YN2t4wrI4bTsmGLGcCMsmgn6pbpQqJL3ONvkf/f5SSGLqZA/Aw4tzvctlqB5CBT
5xNGbKq1zYTn9N/fZ/SvkQ84qiOqq2JIMXuUbVdGMRE=
`protect END_PROTECTED
