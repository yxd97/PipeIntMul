`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9kRyul/7w4aeVXkDQMGVQBpZcOcZTyGuRJJ2ztbHqvKOJP7VCcRJXy1UAGPXEcZ0
a1eth7XidonplNoKGbN26nFjvNrmnipUBvj1l4VOJx996gDcqj6RvR+rsylBME7/
Oc3L9P6d+/EwE6rCcb/uOQ3cWxPLNDeiEYBYWKARyrhSXEmPEokC6oLLU07nqlKZ
N3p4RFN8Oa7u5sFiOvRbBPf+g7xntoxFTIrNAW6gQB0ItZ5vwaBkOyPeBY/sMLLW
Q/2PJCyBxVUd9uae2/rOIrDwOnLEARYTY+7o5TIefkiUleX4bycphrTHKd/HAADx
fO4Uw9BM8sfJOShm2Ls+/rD728Vpom/dwR3NkCGBc5EgOFwGtjiMWZFw0dA5Ftgk
GrwRHGRCid+Y45c3dFBRMQ==
`protect END_PROTECTED
