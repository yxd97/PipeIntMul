`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NV67QZyy8WhSzRvlD0W8lJs2E2B2uIddp2j9VrH6EQEErY8YUG6fD1jJUMxqHcXa
Oc/8uqlWZTrJqfpv/FRup+2xTqMXhVGHxTVbSSqkuVNIJ6djs4qFAZoiUTDSZQLq
4JJy9Sj8aupAR2v8VhbqfSAl9bdEaFYyhQtwKYvtN30kxiya8ANebzDWbSq5leez
5ODMDXX7IDN9+c6HIgdsTRTMlw+GDrGJWCMce9eDyM79d2YFY7CqXk/9EeuNkosZ
EWlAD+rB3cX3wrhTYyRnkyZ6BqDY6ZDpKpFBVoSEqv8wZUtCoYWfAFqw3mU+fLN0
RubXgrziGHr1EIFlKu5L8V+HFyDdQCeeDdI3mGdYNjyV76m0AYCj89mHhCmorzur
xJctUvPFfcLhs9EQSwXUklWa9qby3CX56UP+X3HYw0OviJcd2R/TE7rI2PGPltaC
iupJrPKVCdqn9Fyzz68nMLDh4uG5lodAC9PWcVtgelk7dHMgRPaMFQ1xGBLYaptW
TEmyQs5j8RM2KNhgUdKjcF06ImzuzHvw9US/H0JSpWPHpd1z2PNsKVVQm8IssKPj
KN/lqRa6OzXvvvwAY6TR8SWjcnsWwrwamBeFqPraqMyWqbOSTOmgYxH6l7br0/8p
2w+MkvVAO/nP6PrXWgQ2j9WIl3xHSxgshySmMoIoQ2wak9zl68K1mxBDewmc9Omf
rzVqRj0IKhbH6YYo34CPvKJhIInE4gWNoU1DPwkm5jgMJ54WwzYIKNime28zNAIJ
N9/UxGuyfOGq6MzEu/C0l/C/t8ZR2LUUi3C395TNVNOSOcfE0ENgbzeb9gwOJ9WZ
hyLiB3wIp9A7wBWgCFfotaAp3j8PWyPTli6L04rW+dZXt8E8ky8DkBVD8URc6RbY
iJRL0fUQmZJuhzxoVCSYj4YzJeLza/VkX6oiiWlOIawmSliM+sucJ+eQ4EuQLwPd
qcWAQcoiRblATc7nSgW/U0jdAJ8ud/B/ng17dLYIoecZ5XsxfG1QbMpK3A5r4N49
jbjXs1zH8/hT6atR3ZdRz560Esvm1080hoJKi/RugkIae/rQXIOJdYWbsAGv/xKS
rjvkrZpsd6wfxsIaYNMt2V1pizkdh7ZtWRd1gsH93v6o790skn6YyuvbtxI/2790
aFrrW1P8AzhdtuV4xF3wF/eBGOd4cyKZbCqOeX+kuJaHMiesg8VvuPgclm7R0K2x
2cIm94jUHPrE6LMngiN/jlDngMLQFTXCF3s404hA9mTll7HcjvZGw5V/6wTnEQVP
cZhAahdGxJJGRzznV2Jfb74/NkbS1UuD5rAiXH36FUR0iry6Gd6Nrbp/TURv7MG1
AhaIAbXmchXcgiSRscHOtlryTx3uqLslt9/9Oc1b4zvt/igxw32S9NyjQIwBa6Ic
+MrvFt6okYPlVsqwjtUSJT9S8fOlsgf3bIE2U97a5z1dNm06wtrVmD1D+cgtTlNW
5Eaxgu88sC0pbyjge7Ja27tLfXkguMJ8Img92aPERP8SATsMoS1wXHPXHyy/4vwm
ih3BH4jwRRuCCKJhKkkEwgMhxHH8WBGDhwtxbxfQHpsKllxOQr/xPDQqiyY84Nvi
I8ef5Oq6aA5vdAa9JAYnQBlrV8xEZiMgZTFzCPvr4oxYGodIWm/b9sKhnqsgC2Oj
4YgyPQgenG5KjiKirY7Lhrvyna1RrH8keIiaxbjuAtrzyCeQeAyhG0B3zg90lvS2
gP9A75PIHklXt8aV43/zgWK8L8VczavL7BrTCxoNvtgo1kkr/30faZZZyY06L5j2
tWLAOYDHbz1iYPz9TuxIMYdSuwFyI/6THuGU01XQyRyS07aAqx0ZTtkidrg8TPA2
J1G8nslM6hx+iGF9/+OXRVGAvr0y6VKQVG2WDC2CNkk=
`protect END_PROTECTED
