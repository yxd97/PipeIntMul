`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Da/y4yV3y05yvdE6PGxAPaFcMxkbpgxsBDSuzsBe4Ffki+cJwDbmMKNcMpaYfqxf
B/E3f9gkXoYgKXPyeCEFEbzeJpEHbs7yhTNNiTxuhPQ3lqKK3ENuT/MbLYnRGv5C
QJ66JKFhwBEJddWdOeCxiGCgFL6f8beDYI+FUGc5iBXQU4CWdvVO6LX8U20H0T34
aRipAYcd1QFOtlSozr3YOhRQ7nDnd14M9/Iwb6TYt9d0z+gDJxTrJE4IlRmcWqhU
78AhU2WuuHHlcVXb7Zfg49c2Oxr1tLi0BRwJ7S9W9BVVG9x1obR8IngIv+u38Dyc
dk/nr7JzB/4EUTgCTkbOCZtD2wJ3SVjbZrdO5ManIls0Hw12Vs4ZlAuY1hxyxPzL
+z52cT7cmKAhbMS+4IlgoQR4DzTKwwwSLXq20EKV28vTMNyG3O9tXwSfuoV/eeCE
`protect END_PROTECTED
