`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXHqU3tpWH8P6spKNPmT972YEqWG/XrRmJuRwaXqA40cj3U73f0Hl7/a5r3mlxLw
hPJejt0ycdfj3m0gtiPfV29P0O+wz8GkkN2Y+ELQGRsGmaqQitPRYnOsrH0xU535
Mk1UeVZaOm3JUR2XcZmZjF7l0ibKmWqSZtI68SMQtUqO4idrhn+eJePyq2AQfQ5e
mEkLWZTY91OPAfwS6bD4IjpF3iSo4tfKkacXe12B+HknO1F+jOFvURqgVOQnD/KH
tw+KbkwH3MzEWUQYnQwAeXX46DWcgidJzcrJGgwlwyGGhBIuPm4DSk2kL3xobc+L
WEtCkOYbs/zvUIW2k6Fayn7b2NAYnOOOoWE0OgJLosjdSmSHeEXeStIGw60QBgWD
LKt5gtar+SeIVnXMqHzkj31ihtqPd8ObeWordkCPZfY3t+jNnivD81f0lmJEIgSx
1oGzzvdheRYDlaEkhz2MHH1V3CTVnyoD5HKE5O8WLmppbE0f8wG8HrRUcVWGzu7m
EkABLAQnHutg5msbAOH84eePytWK0qfuEb1DgR01VnopVRL1eT3WXFsRiWSypx5h
jc74w4u4J5DnIK6cL5eNKmXtBklGKYvFjNwV351JoGVc0fBp4rzh5JYRGNXuGq3N
bEHrmCG0HUPVydtN/aH3qJM3aVGnCUtjZUPob4SoxlfDIWzq5OPJkfEpjFSnSvbL
lbQPZI0zhiUfOeYpTsd3GNMGysTH7Uu/KYgMmKyDijZ1Z9rA8SMTYt2P60sMbX1t
gkHR3kGpGc0woHy4iHBVR2HbKDgAx9T44s+TBcceArXmjBXAolppkN1IKwRCSucN
AkKYA4RNUuzQGlyXk2kdciJPBZn3NV8oMMzrH9cEQB7jhgRPkxBvzLVLaq2ANxpb
o98Imx5/DeCtcFwrQMu6FRAzPJrhpJvlwjnW9RIdHFS4WXswfTSNVOq7c0Widi2W
j9gveb4MFmkjqPE3dpJQbvPtf3YycR0Xh7AXgAGJIe5oVe/ayhtyCiayFAvepdgu
ODGJGoFmpc7EDdSU+n2Yu6TzNpzC0b6VZ4OJMus5K8KJLrvGj146W5TSozXSzUrL
LBdukAATMN69rqgOw3kJ2WNO+QKoFDZc+czVIKoVc2A1JXma3G6JAupnO+ZY3SA7
NgD+L6iknM+CCpyfc6eTqMJTpwypCiR19oVtggfQqFXWmVhy6hvc9o0xZU3iLqub
gaDKXhqSqmE1dccUmzC0NQfCvxnKloeUUPj88owzp8rZ51p7VXl4cHVcbxLkVYok
zbg4vA1MZnFnzRxJ5uDUBcJlQLfguTLPHmdnt7F/Wfe6e61g7h4veO1tpzoYUcq+
nBOFtMc+o3KCGKSpqBrjSg9ILcf/aRMgPBsI8LIY0vEh3hYlLcVI6bvo0l4B477w
CK+jSAYA+BG8ed6Nd1r14pwnmaKsr5RZeohqOhZl9smFVc+D9dPGOU4mc8P6nqyp
Txjjrgis21eYcfZqJGZKtaDX26z79+7QG5BWe5DTyW0lHfiT3DVcPewAFSV+gFpG
6aEs7SNe43C/sYoSTdX1ZDQpz72IbnmALI+zVDi8iU/Pj5pUyMu8AW75uB/dMko+
//5PLCqqDK6JefKuPjGZzzsKTZRmyFKMBTkrgFgp+G25kujT2S1LpNlxXRqUown5
avEGhndyqRkdFM6n5kSQaJhGE1p/YptkrP12nPtNGD0Re3uu0rtdauB/T/6sH9ij
+iWruLUSKXldx+D1UhYqByQCvomDXYjyWXrtPzs5y3yFbSV+S1OOBJgcuwhcWSI8
1ddUbkcv5owZyd3KtWEcD2IHFok0sfrfUO3SPF+yDb1L0ML4aa/H8ugk9paV6BBS
`protect END_PROTECTED
