`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T0TvPS7ObmKmDsUXwyRK2d+UEqpv1BIokwLlkuXjtQdHbi9lUIxO9RvYvNGrzXbm
1sFFY+9Uh215VRCo9HAU4zfSOateNhx3DtadNupueHRXbE7R0Yr/oJ0wCMgw1WbO
uhyATddLYgVaRFAd9YeQevkoEPepTJ/MmlY4qxhnKPC+PrgE6K1SvxI6SNnWBJFs
rHMq6cJzrhwszZR6urpi2mdI7mBRau13o0Axcw4tC816UTrWGyVHxHYwCgXO869v
Cqe6/vMXMIi+frY/gnLVg96q1D4oeJ+mLwHMNUp/DnF8hOCwdd0OHVUWuWCEGCSW
DK5JFFn/jmb6BqHaLRAYGHrvj5etivhqpx5DxMHs7fbjdkBBi8Ju3ADefV+n4h2i
chfECmdNKozyEbY1HfhmRQ+Bs+6tLrgaIhPBXFOYd+XyTebfeiBCAEY+vcwLEb8z
TP9KbRrAfTPDL7exTTbAOmpPstwSivUuAylcH2ls4CVlodOguHS8TI+HUU+UE0KC
JgDJX+1wh+pcXUaUnEp1jEEd3Kv5Dgx6TCWbCD2PcizjBzotsCKqwkLRws26qpXN
i+pCjLAk9rgK/dgvdzuU5pNaF5Z7dXFv28wvKj1zS7vHWk5RJe8AtbZIabu6f7Yx
eY6TbuormgnC+hlgr4CMt8y0DuEbg+zuUZWe3RxMvBhhMTylvj1FSzrmxY0swchZ
wWF+r+quERHLpBqkgA1+NMY3B3YKAU58XyLceHmnL97/l0o9WD6XgpwDah9wxKwo
t60gWiPau25BCTRC7+wQmGFv6cJNA4k8zC+9S9x6LX16RbImAfoIZdGHhucB2C1g
E/iOBR+4T+CapjDzxbWo+E0cXX/RzPtq1ltpqKgu8IM=
`protect END_PROTECTED
