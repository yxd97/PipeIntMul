`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JTckNkL4K1Gp7UP/73i+0V2PPTRIcTlyFAPnZMO3brpE4UjVsTdHEo0OLohYWKqs
wHAKW6mkodkDSM/PL3kCjjFzapvhWYzZVFN7eOw0TScKSCKE//vgTN/3+xioN4Fb
2D1OfgilhlwmdjQsSM71/sIvgON2TPdaY5p9oUzzs0tH+IibbeDW4C/jFipsYCMp
dhvetoykyp/Jxym4GqTPWtwcVlgHO8Y3SBTgN2T0SP2utoSkIEBnKSrsyOfxftbk
tKwyLa7ew0UhZXow+h07ggQjddlv5Ff13aSnEw2nN7vvOKkIcYvBnQZtR8ZcvEyl
xrFFbLXYfVpUwb0CbTsnCBb6IvuWFgUw+VvDBhSpfWxH9s80/66Z44nUrRYaEKD9
Jd6OCccFwGZOgVQCATwTd8qjEd8AMP2N/MZGf9KZCF45v5wpLSIchvQs+1+RUncK
XPd6FjG1pQMI1uhWnI7FVeLMGZCnYbQ0+LhWXTqcA7+aYyJWK55w8LbiZXxTbOel
ZfZaua7LAvMZnnv1feELx+gN+UThTFNyLnHZQk9kX5f/7bycGcx7wlCC27YjUzYo
Cbcfn6hm19dwg3w9ijC9BQU4RRWTKfGwlBCVhJdP3K5SV164hMC/LCW6UtLDA8C8
G/msJEEjL9EbFaPIZYaJJQ1SsZMVtmFi4m0zVA+tQnYFV7AA7iD2uC/wPP2TTEiy
EVoHcEKo5MOKHk+8WVqeJ+U1Zqdp/PH1HfN3fZ5dzzT6QvLxFy3mXGP/TFV6KfMB
Ad3o5i5oDZTdErSeQnDDhH2UgRPy1GgAPpGTQ2lgJG/h5O2eNVswkcXKSHwduc/v
1By9joX2rXoEzDfpA5suhBug+W7bK7GyUECQ1Gc4XVfa9/mZmMMTvkO4O9S3qmv0
+GndDQISE66PLk7OLQ+n3wJ1C5bcKl0woVt6NJ/bplkXmB2RcVFlAF7Gm7s//zGH
0gAF2BmZ0j+2RhJBTbXaGjTyDPGxXYXWQkiGq7lxhTmT3D/yGnN+EIUZ13gXjM0F
j1ET9bi2b3vxtCnL+EoM0k1Do8qr9X5Mx9rfpvDt4M5cwGgAx9ghh6EN/mzfUCRF
yecbkdRMmTAMOF4PVBW5Qhmqy/0MMkgbPTfC+QJxq57JN1+hkAiry8qzXa0VecMR
cgka4h/XY7btBJWIYRVdrio74+1tElBMELvRyhf1POWzqUfi0dL4I1aV1A6rSf34
MtofHOEmalQypenGgpuRlU3VR0IPO1IBlzsehC9hvqQ73DQD6raHkHB1jZcO+J1G
7x9EitQqTA0I72Fdj5Tt8OqixBlrkcXTzRynx6knNVYPoHAo0xhsWVhbhflK/qeo
DpDvg7UUUCtlh8VVgzCR5n8UDl7ITg8D2lJT6gvWmIzh98aJ/FZE5SclQAmnuAdc
NJVyzIPYifb9j7KvarBZrWIuO8/EsRfiZgkwePGUFFcyzusZX/dzQubRTeMl8uW8
FWz5uGzWB6xXqJLW8kKkoJvyQcAQ/i2xFbbXYl3UjEriv2+VU49k91FEuKlpQIit
AWxxvYGukXqY2m9i5kBP7lxQEmCyZDdg45VTXPvCkVM/cc7Q/UfhE4FF4RQw9va+
HrMIOTDx+7LlXwNltim4+7/QsoixIGJ4eAXcTDNFuKG5lZGReoOZikbcdEJOFIcE
7kOcXJG1TFcgv56M9L9OmiJo+qUJG+/VcGK1x/SXBy4Z2DNPn+5nXLj8aJWTB7vL
6HAhjAt9Z9LfZH+E+ePS1xLyKb5INVmtzKlAkgTQzMTy9ZkzxLkRN0D+kJeTOYRC
Uacot+yIlO/Ac6GPUIlH9jDqyIqL5592lWK9cVu5qyWLlZYEkPVAmloRq3QJvxnH
WP72scfreSeaZsBc98aoGS7NrhTgby0qnIVZzNmyjmG1rMuzbrMTEJ+rJlcAYB7f
+QDroztKERjw1tXBOhIiNF/itWBmbEA2PWJO/0h/LBTUdWSu5bIGHaWhovwadooa
SBpwyKP8f/DT4DTxrTlXdnzygp4DemUslHmsny5ZNpeNQM2y6yF6mx86sxksb3cE
cHaJgI6FWRzFtCMitSuivUSRSddf9qijb8TtJv5jTcnCo0yUEbxIkUsZviURrjoX
asI6t5/85jzC3eMCwIBuf+dBQFcMsdEJ8+2R1pjUow0=
`protect END_PROTECTED
