`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUGyF4115EVTy42pLalFHOD4xpR2GQkv+9VRqcCCwklwhV0d+o/pspRECjRFwvB7
Fr4J7twTIsRTVg4rlMq0A5vbnKW6uzt8MEKnPwT1BONBmDKfpsOjL3YkRykbXjZC
1s9GwRHNjfDISvHJH/Cl2mQcrQSJzHPyzbG8iPn9FkUBE+eMwDttFPlm0jfJOXZd
wP/+lgXf9lvZEZ/fgPLuGFfvcN3aP8u+z319RfP80CwciMxZF8mTYTNm2RGWL7op
IUKeJLn4ZDnf+dR1oNifDKIU7NbjRhf4rIllIuXC8h8Fr6WF9RUByfUffDGXDyIr
Db2iGmYarsasawdSmN+OU1mgwvzP5JxXMN24GqgcjIeNDk8j1ZBiVXgEWcJlsCYO
AGdhrkVepDh577Ik3aJw/rF1y2fG3CDJXcpwYb2nyGnLatabJKAQVv6g7KT6Dhsj
HwURTVJNhSEaXM8bQmNUfJASBT4kn3xGPzGh5emO/cl6TNYXOyt3OOMCBf4YnZh7
8ecLmimLN97XAKUvW1H6VkCAw+f2vSBCdrHf8zojlnktCD61mx7RcKLOy0RwzmIe
XBjvIge+N+LuRnRiDpXllAtlzFBsxBrMRup/KuzUP20hOv1N4gmhAiwkL9/NWJij
vGXpOUcxtk5rE676vLVs/gppmoeJNsfMUFjsZrcWlg1pzuu3nD9JkkOFMQVYFzhX
R+7B12DC0WNIaw8aSpDmnw==
`protect END_PROTECTED
