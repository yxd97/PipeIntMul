`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZaOwCuZ3YNkkliLwewk3/gi/pAHme81SFLzV5zfpqY/9AMuHrD5XNatRdOBvGGT
mwVRPoIOH5j9wcZszqmhzSffkvkLAFWkPQXjjmiE38y4Qbs9tJPrWGyPFAyadVbT
I0pssPaJjS1yDevWWPsF8DoHMBhFkLTfOz7AZCvleJiqjJjJeKtnKLtDLgimxaJk
kkGqEyK75fgjq3oyEOq3P7FQjPUifJa/eMq1ssJyVTCZsTaRLV7rIF+YcTeUrAlt
UenRVYZjhEwwkMERv8YDaFWK2/yya4SmJm7jqSxWIWJcraUVXQDZ5EenecE+7lus
PuVZuoP3+1OZtN6N+M2WTXbA2gL88ZMR5vMMQXG6kTUHdadF0Zm/i0YYMweFCkqb
KBCkwarJMildgljsQ1g6kUXQf3Sl1W5SJEcCGfYlRAEZin4yiwq0Am8YWE11hS7s
hDQv2zLPajU0fdrb7magHf/yQHcQWZ8/pMX8P8g+PziQVHwy2gmrCNuTXOa5pp0r
ZN/iHfEHdLh+LO9HTUe/wkCMSBia4z4JGQdzdB48NhOZfWeHFKeMPo7pHbDVj7qG
jMYh5Pgw6xNRE+Ej2dVR6F446as27glIiQMXtZeNaHH6Pfx/aAEkKIjybaXNJdBC
vYCIZ/Zsg3kyk5zPHFr8DJaP/8u7EEtcGC0mJDmq3PE=
`protect END_PROTECTED
