`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ojedLe5tqNJnqWGRGW/qmnVNFR95SAvI7N7WbZD6IG3CYIvJkdS6Vl4/+icsVq1r
K6mRxEGWGwsVbhnWzd16HNusZ+HLqWs6gjZetUct8ZE0Kr2I6G46Lug71C/hCDAK
jyoVK9WJ1mkz77NNtk6lKrayOEbT1rYcfUoroXsgZ5dv3UVHfOkOb6T1OapmiSmb
9iTmBCHX/IekeyTbQE50iOX5EFTM/+ScgWhKEsC4NSaSzgzMAN+5hbVMAkFSzo82
7PcUiMmSFP3R5JvDVQv1T1QOoQFmwJCNVm9E6R9i6xW1n3Xhv8MJULBWzgc7OB15
8caHO5aBodQtYGf76NneTxnsJ2/iGCZQgdhorhbuxQQxEVQXTs2Z7kzzRjD8aquM
/UwT3jhq5rG/RDm0ePUFvuQa1aBviD4cpGYLek8hIYV+wNsizmzWUXXpFIZ0TeDe
Vy/aBytK9H1MpFCEePd9qMzzTb4P3iKmSaDcqlRyip5pvJUlcxmvYe+Qx4y/X/Ij
SYKNorNYsGjhmNI/cn9xCe05OaqcndJ1u6S5PRuTFcsZPH/VDKrtVu+lVbGFf5RU
fSYyVWs27QONb0l72wxFaR0sp/McAl6WSX3c/fHxmkibr8trq2MbKFEMquqTzRQ+
Uz18LQzQNKU6JFrrgBFVlQecf1yH1ywkRNFHfZmjTtGUeF4mqtRoH8Qab+06ZOgt
hCgkTmE6wLkxvSvjH9YLKFRFdmcO1aPRR0HOeytLMyUk/IvKEKuwE5xvsG+UMYw6
PV5jxMv6jTJi8qd4auSy5g==
`protect END_PROTECTED
