`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IzdO11wKu5Dpw+rF/FVUJdoEMV2XpI8e0YoTS9LxHTj4YqmQSjyac1QB0abKaHhD
3tFOzmoIpyY0Riip/tF6B6JxUK1pm7Y5oPxW2fhzOZbVQTz833uPKQ9lgH9z6Ori
2n8iwYX25rXYDeV5+SSDD7CY/bcXqJKS+OG7uvctSpuFFgY+FBjWMsKlP4fUuMsB
ru5PlzOr21tU7QzFji0HlmOSEv+BryOQVPwvBU2sNPa9A9aCEo61Su1q5bf/crDU
70ja3qVmdrxHpRrRhhxigPym962kA4SQdnWphTxG2VWQzOk1qNXRHGRaLAFc34SM
ohKZrdReMjUURiFJOcEOU6Xsie/Les3AjissRHf55TzA4XGo83T6j5zaRQIapOsm
F7+iiROglOiQGyDVCTkb0+0bvvYPfYDNiHg5hSwEarlzDHm//uIbqWWSyeMsndR6
BMKN6lwT2gKqWzCGyBFSABiOigxcCjadtqI6ugwAzxWm5QFL+azNQuT8Ict2JUGZ
`protect END_PROTECTED
