`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qpd53NraQ20VaPzoeC9Xtc4kp4AhPivKItS5zPF5VmJ4F0Zw+DHWAjQ0p31lGrR1
xV+SySA9cV+muonbihH11T1RBx4BUhj5w83vSNE8SFZ5yd5lJmcSj69u32cXkDSn
4+TM9Tuxm0esVz9zAHgvPsynGSvCalgQqLMmTaOI1jjLQPFSpW70wN8jb81IrYIf
5IiZNxOSqA3rjlHseN/cJS0XIMFECuJNsH52CAp9hAdfR1UbpFg26+9G6BdwREGj
l5AFfW/MmEQKQTJDf27EPZ22W1cMN/P3eS8EwI9W9VIKEKyPTVyfCTnvkUMf7qEN
IGEluQ5IG7NYamLV1+t/NXHpLruuZogiE3AmzUNA8h3hEx9RbvqIqTMl9wlKpz0/
NBqOknbef45yMB1w7/ZpM7288Qf5rLn5RrwFR7RhW6BTPFsx6eLrwTW/lgn+nn7m
tLrEAblsjnvH45wO6+vZmGlydnrxtZ16k6Uft8GkV2SEmIDenJFLK9at/S11ETIj
`protect END_PROTECTED
