`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N/1tiHkjDeUJjXtIBq87RjOs9QUGYV1E3uCC78wjNadHcP/KjuX9VeCihZa3KVWr
sN0wadaBwwT8wpAxDnzEhumGZtSyA9S0mQ4vebB5XhlxiymCmxREgPA18XDYl2m3
F3p4H6HM/AzBP7yQVqpheLHmQi2YWA7LLfZ7//5IRoVNb4Oqis+XFpjkxv5vcu0l
fkTiHc9SRIDacbhXV0JaVeGFjuyWeiCiWZ7h3wOMMx2NQvRwXzbxkM3kW6tL8xBe
26yZnoke8V+VxlSqX0/Y4ju7EfuxKsmDDbD8TYFFS+ji7q78lDltN0eT48kxbXMx
rWkv5q2U3C2js/0AL5c0MB23Nq0ku43DtKO8mKDy/0cRdQZLIeoNfeev9OCAaGaT
WtdIdTrMGl4SnQB47josGmHD15oUAMwsbiWKzg7DzKel6EJMpcSbN4EkPIo09AFi
zarY+gg5nxrbEbeJGmazUG0FjeLVvyE4TIFVBSB3y2yo2XHj0Km+peW+Pttzp6r6
vI/fSawbGdbfT1hEdFuqSWMY6TM5qcPy1wCylRiEWpFuuomL9U9RnYLONW6qQLZo
myNbo4DJH/2eQs5iDCffLsfH3WKYzKI18kaC75j/2tHHqf1rnzjyUZyIBcvqevtX
xoQrYAI48MuuJZ6XlmfpzZ5k3RtyThe0xwsdZMi2IqTMTu9mvNp9QlIzunYZgifJ
xU9L7CJU9RbE4Qnutzdqza+wxxLoZNaXcTQMt4JJH9moYFjLYM89G5UvImE7tkHY
M/KICTtma8C5YlZqpYp8EtB/4b0auYjYQJklVgU8upuwXl97D1qvMBrdDK9PJFM2
+5vLPIOtf2lUoIZP2IYDv4yfNf0TOocYPLcVcOiI1JD90Mo/L51UlzE3XlBDT+FE
NSLR4Cbfu6pLtD712biG1bjNpHT5RxbHmb2pZwk8crxL+sfTLn0+nmiNYcuD5xcT
+nVEOQvDU7RAQJIN2FG00C8/4euV6ODDLLtxeYzTTzmycHRIl57PPIKTILnXlgBP
QWI+BG5YK3O0AOHujE5D4tUB6/7+MTmXkrvACY0Hfpz306WPnYkpywnhPb6+jonm
LTP4jAXEV8TxmN8h9X8/YB+upQg2YSxNNReSBIjsj4h2XdIuPBoRTHTXsAaeWNkY
rQIWkTBqUxtm+0AMHgJuuO8IiMfZUpjdZTBJEfICaueOtkzAL8PQIM+/tvjwzZMT
dohZOpJSl3AvhNjEFk47PrlUbxsRcfFE07e10Mt0ulpgRlgaPaRL5AsRd1S1W379
NqHu6yxJ29NVMzsoQDLkyKkn91KgK/woYGrjMJCux/EqN9LKKJvjdns5x9Uxe1+v
JT5ymVyZ00SOnUBx0Fvzm+Os/pbJAty8NNSYoW0tjZIYzTCSYTleZDiE5yOhQXAj
janFKv+TFgVje5rDZgv7XsNwXp7PYws/1a+AYuxERClhIDDRdGRchDXYdu+xLfuJ
u9VgYU3YdLzQHOyEw9FpAw/tJn/jPSnPTKrl3HrKNZdM5ze6O/c7F3DVcetQdKMp
FNOCfzGXk1Z5lcb2FtBO2DeaCHcxpnfhY1RtcxftVFQV02j6e+Mo0wB6EWV5Q14C
xu09O4Gy2qkr1mFGyzSjYm/AscMOGuqsUdEgb19ER56dcu/Uko2Fai5UOcarnCLF
j0nuMTbPX93wKWwYRqrtE0ehpH2oI4W1IWDyrKWhhuQxEwOWaS4Aklz32G3Mtpsu
kbKfs1Li/ZVc9A4lGTdltJFEwNMoYrE7KKmVfgOu8v2Rk4TBCdvWiw0zVReVJRMl
5/p++s3XnEfqre7bKHwLe+HBHYk5h1m2uV95H+QOZwhBVJTAKNNu9tmrnm4llIUD
OtGYuvP1Ohi69IV82CZTj0Vfal3C+u7rRC0WQ/MFgb/MxWrad4uiCK5ELX+56UDF
huCxK3MKKR9PCawkBDSihsMPfW/NzW+yWOfix0lebweUB9EjACfyBUuf3khG4hvh
CUEpKdYJSy4Cg2s5IwVoC0nQ4NRZxHuyQ7Fvd0Y17oDN8CJ6nvBTEVQ3dnUwx0Hl
ycHxUmJleiVXlWL85AeIQHW/EV1uOk96GtxCnmXGZIfor7dc8P8catMiBGCzVYOt
VfTY0HQ4sb/+y8Z40BakpHIiZzJbVkUJcRI9HgTEwv4vqNFSZS4RIxv06iOz5LBm
8i9QuaScImsm1gCdPkGJJhWVPX/ltigZLixAmAo54ykA89lkYlrkbFAI9sIsl/Ya
UW4kAKAFXR1XVQixaMZWDkr0ds6oO3av3iHHL9CEwDoLD6m3Qh9HaDexUIrh5s4v
HGo57rN+PmwDc2IrImIbLKs+dAalCCH4O0UXlkgwOdBqz6F5Bt9BAL/aiI72zrhS
fMJ6hnfU58s6Xkx9Z9hABrPqXv9d3CPdyc1yA9EJa0SfiaUm9uOfnst9hTvbNi/v
xzDMBn89VEWw4fNkGhR1UzPc+YorFBmYt+UmfWamSNGTLo1CqoSh7zS5bAR8eAbL
EOyk19C8UERL722hVsg/4ZJQL/d9fWWqwJPMWmneK97J+0cgAfe8n7rU0bx1YVpN
ST6etSnlot/iHeStlkwNdikUDNcK19QZpozcvQG7C9TlDm8ReNRbv6+kuxaWMjdk
bGGQ7EAwvgm+iPHwbHn1xGJ3dAKE2H3YwDnMJW/YLieCKSlTMgVbHc3b1iXyOmAm
uhYgnQauUfO9hIRDPHme8/eLo2z1jPEPpYlgiyqB69MUS2RJwngLUiE83xIKr9Iv
B5MKNa46KG2pAwSD28jpZiaaYrjibUEZ/9imfOrombhgLu75mHowD7j+ShbBnTqa
icM9LZFFMdFRgRicpXU79sOE+ego6y/2NY+VTdbRdbGvVAspUdDoaecHb7GXRez4
3ekWP66ydM3jGxTCqwZtfToldNc1XJfPt43Qe4cGLwCXtpcwvSgvP5baOuf4eMqf
JDfx40tTuTwoPC9pKvlPlpYbVPtgkgbOhedF9+gCtxVPq9gQ0UYekL6FthVE1eyW
rCKmg4SbpLbDCciFNR+IhyvisBiLyzELK770rbghWq9Dp8oDe9BbxsBL732Fwhn3
S0ravzkqmRdlzOC3KVnDrA/R54iooKlNHT2qW8JpMsTUD47RpTyakSbLmLbAvZCJ
fL8xLroGS5ifdAESkoYgb4le7OLXdhJSxGJrkmHW6gQsVojnYXWlvvnuz9u0odRK
9qY7EnH+aUqJuGrL9nHHkV2roky402j9mO+os/TSeNP7HJKX9K/2dmM2cP4mfo/k
2/jyt+7+ir1gg/i0TZC4bac6oGkdmh9tu1Bhz/W3MwroJge/zn6y5AxNR36tHo0u
ARIC2UGzFlsGDxFzYTEF7ZSFAQoaTZ1JfyJRUsziDoxu9YHelfNX9efbNQkA5VT5
5RKu/PZEECRirxKVwTgc8wLb8jm7rdzH9msDP4cH6r4wR2EJScXrLMtRkt9p0zS/
FwoK6BaLclPhwH9XwXIOE36IvbKnkk7RvuN4ehQnuoR2uIW8N0F41DG1/GyQzgfP
BCzYU6S6PzSjWl6ZR983Lclqt4uqCLA7eE9lBYAAj25HpaBNphZMx3xsogJnNL77
x1WqloIasU/eH4nRmCStoCSqHmrF/05dnkD1OJ1uX67tvxKEsZL+JP/Gk3jj/rGn
ESq3gunObRSnsuyxShP5RdokcK07Xh6QDIcZD4O6n10QN0svhEHeLhfXOFxAWQw/
bSTVWBQYtopye9HlTd9YuqWcIZZS2h6FpIZUNHfg+r+q11+a4/fakUHKFKgGi6a5
EBaBGAGHK7nGU/1RmKCanml9kGhvwwt4LZjNfZbpTUCfdrKyAm9xThbg1WTHczWk
3f83p4b3Jfd4XKBz/odIO7xHLgfvwseBTCMfm5rq5vlEKQz4Bjz4xuDQFl6HIBRi
/9bTtkrkuKIq8CmH7wwyOo4OHDuZfwu28bwWxiyw8r8X3Q/dZFAx2iWb0Zs/gPZv
q0EJyzggEUqjfk1wOip2g29QYwVAfEqSi3yV1aPSk9pykbPZ4MNR1XTsPC3MXLhJ
HEYDt2k8ApGszW8sTT1NuLzLMsRILQXTUrSZWGdgFzFxZ12/ESCIjaFypm4oVDPm
4JcBzSV0St3qs/OZ3Qp4XuK6RllsXW/8P7XKIErJIaz4PzT4unOFbiF1XUSG/o/O
x3Hzm5HpbtM6DYjRVseYw5rW+u2VDj2DacpcDUsDSoxoy3HX90/s7aHPyRHEKifU
rJMdp4ElnFjCmdSb20FC/oeP8BUEOWxNRyZ7f76dNRtujXpNZkdS/XFudq88llF5
xSnTjYKQ57p9SxoOpXYyKiuQrbme2M9K+GRZxZ+O0C4ARqwakUCFN+7xHBQu6ZW6
MKzeaIwwJG3jelY71G/mTFB+S2oa7+05/CnZ29L4MMtAROM2N63P5nIpTEDdUEtF
rSAvUjElovMIjayZWo5xGGztyCNMPqiVehRJnv4GjLvM5+wNA2QFelIz+F8M5o5M
g/9EljVljepgWtDJzDBUTgKyq+3vveCDVa4MQipsdun08hAP0Es2Nu4KqhWu3Oc4
FQeUerk7w8oqUJtUoGTL5mpSc2q32+hvnXoZQ3shlh07GHyfMnzH/54m861fPo4P
z42yYp1Eke+BAwOYkdK6Rstnh7mKg83Q+QlFxCxtRLptYI3PMggXPyr+2uBb7tpM
vrZS+0U3H3LHwYwGs8dazuDABUXJPx9DuXdRTapll9vuiJNzRdqpucGQB3Tkdz5v
zmfEzctNKbfrWPXyfRbQzMi7F/i1N/lWDrkjJr9oH7I7P3OhkLHOKP65GAduI+Xk
ntiv6+/5aNEgaGDD4rHruDtNUP9I0x/qQ6w7+kM3PA0e9IBVlIrSzU5jfRjKz43e
WHHFiec8L+NIrLPg7BXxZROF4rm/U4m6sCjKBAsYOPURh0Hc4+QpmbA382tgWEn+
iYzJwisgmH8PNNnJX50LCVNsUAtJg1vlFSIVGMYHzo26XkdT2gYpecHlhow53VfM
K5KByp1mAprX7QAo6OFZAgR3TIBHrIc+nvW71ri/x1jtBL9QTg23Uk5YA479ZELn
H2bHffYyRiNOu9pZW6jMw5h6rJAY8dkTxCeBRASabPEHK6dWVBPbUxOvaz4M90Ax
qi39fgoZQ5+eXDzV9VIHy2sxV6O0ZyZdfnqor9s72HgPfekVxf7QyYFDBnAI+K5n
0pCPoTBWiX2oShXJRkhMX5oFf9EIDUVpksTdDppyWE7Oe5EdDpIX24g6WXFObtvm
p2snK8N+yWKVLuyCmQZwO5Ml13ekegBVSutilQmF14c=
`protect END_PROTECTED
