`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NnGSZwBmg8ajW5bfAWs6fxt4nFHFqMJIQvOJ8py0jcCbCIFVTBp2v3wpwgQPqpKm
AJlFlEWS/F1trd2rn3dj3yOJAsQWshGqRYyAxy5azaEDYaqxPqye16D2u8pvRUIn
l//CFOvEeBJIQdkx64Qa8xU3XzlgR7MkNqNeVu8RFpO0Qu7wWLx4n/4RuHWXtIxt
vmZg0m55gEZoaZEdGc8/S/83zROhKEIn47tyxxheaB7+Jimel3aBUUI/gsAcXXUQ
il+Iub8i1esWnuBMU05Dx4Zhxwqu2AcyzASvbTUkK1Q3SYczbo+ENyLWlellCEa7
+vh3yS2BxCg+6PsWCyrrCZ5MAXOhLRZRWxEONZ4tgKqZS8t84QQ4d3mln+ZioaXl
0zT3nzKdhruINHAdXM+UM6ySMKRthZttqMp9TyKhZILXmOfVbKPTNNPmYWKLNIhI
nuhdQw04vYEfLmebMI+HDg==
`protect END_PROTECTED
