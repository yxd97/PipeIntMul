`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zapafLvRcjgf7pbhb/LDlAl1DiErcpnSeXJVmBGl4rOOE1tWZahNMOjvwmDI70m3
v4L6jgsDZ+jCrIDBrlXwaLSrLqzBaYjMVxU9EzsPDN2O4A6DvrK2X95tfQVkhbmN
lWbjM9byyFOnep4HcX2NVfYQ/2NPXK3pYkSBF6n8FO2BDH6BZOYTcoqsxZLFrMVT
OegpNtttDAoUNcyLkD/Rx9w16WdPaVioF/yHT4aI0KIm9ItFM/k6V9oYLZAUJ0LI
Mi6GgVIiLywY6olFPbN/UJj7n8mttZIhZRg9P9k3JreBaMxUpres2U+nFlT2gRJT
nUjEFL3vjN2LTnhW2f9/3sQUrFhBf5Y40wG2bftKDoqVekXO5PvZ8PFw5ne0BBOS
IaJKUv02U1e8FaKLJ1QO8L1Xdl32AANJgbPN74uI9NM=
`protect END_PROTECTED
