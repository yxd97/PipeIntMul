`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7aAq0oEIWgeJ3sF74AXfK/GVl1nbumUz77TztDFrfM+36VPrb7uuTrfZ/hBu2mKw
FVY+ByIjNvR9uNlCoJpBHzJCsFLfMbW5v33x5cW0JejH2N2ns6FSrNZq2eLGO/dK
Y5OpK810iUDnLrzh98KJ6hhTL6OLQA3f+noDfkf93A48x44rYVLJnTIdyAOgP2NU
a5Y3P/9RdOKoXGVeCKrjXoY48BEeFPeztRHhiV3VpBJ800se7GiRXplXKKA4I9hH
lJcZr8Pq946HBHZ4W5LpCewxkzzvoBeMUAEVNcouF+7rCgGd1OoGUzrU1pmOebKG
McKW3A9nNA3boZ7l5Iy5nCeO52LrQczejPHNN2CkLHs6P+OTxWYMG2e1OKjNXHgp
/5BSOHTg5RMh/Uzk1qsd/3UVv20aJzgTboKdM/gKcBoQLStMeBOhNYVZL3J7iTP3
DJQ5yPzNPnEr+rNMedAdHfF4aJCBMptS+VtRg7MBnLA8z78rr7zuMv2HIXXImrNi
EdXHpFZrytl1EwSVmkiquWUNshvsPkvUh4Sor4L4KOqbaL5tafLx97mt8aiwWL4I
05EPtbz2KvH7VJCJtjUgwzu2Du8mRxiY7SzO0xlai3VWcjp9q4S9B5YAmfHa87bp
YpZESF1VF6Mf8s6Z5NZRbiv9RmrB2cl0CZDcuW4pjPTpnDjD5CwsH/HXWHOmXIKc
gGjlmcP05VtqfbkvbYgzsguv76A7bZtOcrhyPjCo7JZacHtsetTeqK8e75CJepD9
kK9EMXWv4RRAJSVyfjTwm+xhNlQXnEea8u7VuLn0oOTM8pJGKFxfTCspVNrxcA6r
FIE157jlVOM4aMIXiHb7HwexLLs+zqsJXJP9gsPwAsmWVllt02Tl+dc0sg7w1tLU
yAAJUX/uh9kYgP1+sT5w2nckBRBOhXOofvYvhJPOh83eZFMFPdVLJihWJi9nOL5W
dPJk9ztS6XGqK8fCke5CnCGqE7zadJyl2/Xin0Uj1M6OcpLtGmXQlDEfuC8KTFJL
mWvdbTOK/IGt3tuWatLDK+1/ORN+M1auaotqDeszskp+nyUasHo3cqd5XMrDTKry
/nJjXgU4HPvNKG2XlZ0aDqCO6Go3ishkaVPNbGgv4c+qX+0f9A7+vvI4l6lXueuH
AkUX5Qo/KNij+c1ReW6VeKqstIAISMJomV0dJTeSIk25EcnszT6in23mHZecwNCX
84IWedP8MC+0Hw21RXHIL//lzHrZHE+LQlMdj8mMZw7dpFhkTeKzWOXJLk3vFIYV
c40qCZ+qP+coMc8x7TNyhnwHumyvVGFD+N/dg4kuhAaFApK4UQglSK4PxgyeHgth
Ws3YIB91Q8kJvZbAtDnsZqYIV7N+JrvzcFgaVVZWC74iJ/l44rLJI/S4wU2b6cOM
qYt+ottFPsJEjpI7+n+8ojXBTVDrp3gIGtkGWKuOr76gSAza86xI5E46sJuvkimK
UE0rlKDprL+jlJuoTZMxC4ly3tMzHKod2Gn8otwpWz30XLH65zyQhOCIpsF4C+Dg
PwWIW7y99E1TLhTD4LpNSRt4+WEmtE0jpV/FHodrJqbe8FR1XLKlXn7q4ovKAygq
Afiu+dCNnbY9YthZeH/9t9FgOXe3jDgnHWBF4LcBts+EiRlMCuQT1bfFEMZTO8jj
UlHY3tXzD+m/GC+tqRtGFNdZbndNNLTo3i1qLmvN2UkyWKEAc9afB25T4PtgoGbM
rzBiYeZZpKQv9lzffmM7T0FO9daIiEirAlxfc8uk6aQ66qMSUIj9e1GaBo39T+3h
5Trc3ODaVMqz5ACzoAcw9nFIBQChcmy3pzptZIod2ORbffmWi3Msweis8V4HkXE0
TTMDtFVhFVZLpK9T0bOUu/5j4p5CdIpg6qhPKVHXCSEeDmMMjMHGRtJP2BdjDAdX
z+PlNf/6wj+RZ7eYIk98o58VNbC50r8WdY161T0U8oXqKypYB+eKojHYOzeZ8BM9
bG6VoAtiycXZL47WkI3MVHaqBqhXY6WIseB7lHB5fCg8rWNA9iNIS0bZvHzsQ4jK
Hfuiw1wnSWtZemQncyIaXUNrGTz6EOzstJXfBRhHCRoP/PUVP+FdnYS5+OeI26gu
OVyPVpNK9b7d8PNwb68Pz+kVWIgue0N0DXj7nnwU+/jNZQexdai0tLeEcXto1P1R
+LX0o82esQoEqYbRKUTxStCbyqf+7gbaET1X4WcPuCGpOakd4MhwLw0QQifLz/OK
/qXC/dB9PdpUz0zP4+OUJ51IMXfCltx1GtJEty0qKd7FefzF8olfL1jPFqqFk86g
Q6kJIoh/JESjpM3rsOJ689PB8usen9IAVt8ZneWWFfuPpyPTnJBu4of/4LDfIXI3
NhnDsHPo8TFVmwLv/Tk6ZFmKznAlOB+I88/AcP43FhzB1LZrM028ADu1+8SGyhQK
kbudNxCFLZIXburmW2h6oXrUtbuEeEvpuzKzPwEYwQ9pp+sl44FaSxaFMOhmDDs1
e3jnNjl5q8p2CmZ/Pc/S32IO7+FSz0gNySZ3b/XBleNY2T49YLS3KXgi9KHxkoVA
tROdx1VTJkfhKgsr2ZKL4W3+W6Q6lP876QGEbuN32Qnf8BLey9WgcA7IyLvB57c2
`protect END_PROTECTED
