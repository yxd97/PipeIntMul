`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnGP6pQo6HiIAYeX253GrqvUrXuMJ9jc8SOjp0AiDV/Wk5hcrWl5DMdZk4miK/BM
UCLn1TMe4ICSYNDtjF7TK+nCmSY4+iw2L++eZXymJLqOUxrtqNFaJgXmbue5XL/L
JW5FfpLPmy9ExF2RWYlKe+SP+9GA4jQfvwya+FrlYfvoNkkvDudB8o1AwWbFwgZL
3DwOXe6mBDcjTJ4Dx13XiCPPIhf5D/6BOi8WnsjDcqQDihu/e5mDmYD5uIztuSJO
R1/6iR0LnwyH8qfVkHzPQZaadGZweqM2Y1CQ1C/8Ld6c36nCEVF/CzpfkbGS6JS3
T6MJM/lfFXJei25hNhbqV+6iTp9aBpKn1eQbrWdToLzIiLCqYvJ4MKAu0hFHAalu
4edXIgNSgJDdH917uvpPoZj96K4jkfzEs23Un0PGmJ2MmXuz2/cQLTrVZlpuUv05
sOBXf4kqK4kkoN9xVN8yahVHIPBUD+uFERsC8witugSDy0taRdImCLmmPCWYLGKZ
65ajqLDXxZ7KATm7UQJAC96fV8WHuUqBYU3DG3X1W9Dq/medcViBZl5Ljk11lvWK
g8bGWdUIQH4mpc7677PbooeRMJrTj1k5xkFtvxfsO4qez1igffo2/u6zAQU21UNR
SmBJvRCBbrU72Nq0nCJ3gLYI9Q6q9CD6zu8HbAQXrAbuiTSsxzhdvbrzSqwhf6id
s1hdun7ftHA4L+wjiJRojxUe0aGI51lbhmjyXl8pHtzS1iLHdh0SBDAQewT5IQa9
n0qd5xmlmQ3KpWqcpzt4AVgckNCozLRly9WC8bvBefI/zNHhBrZy2RacqvoQFFqd
WljFxr5DFtfGz2c9hxGTupk8raZMTiGJaLs87T0DuteTHQrQIC8FeQcmjPHeU16e
IjcJ98E6ehh+0eANnXbdZ3SpLTSR4ir4sYEYnNz1CysmuHvdiDL08hSeUgz3+l2/
z8RdSnI9izIHc3CU4+gOoicAg1HwdsQo1Ehx8L0PlfmqZWSCx6DYNzZBDedXXL8j
A9QcMHwJRTKdTb6EW8MoAzmdfu4TFgab/bduC9gJPis797BsFRKkSpsbYb/8PUEH
LUclZu6m1GYMRdPMZy8hUulJGqQrh13SQZJCv8AdFbKr+ipDquY6Hf2rIwMAC5nL
K4bIiZBiGCfUDd/AQ4WZgPzz6pQ5+KZmw80UXQs5l7GB+8deR8AykekR/vvEruKG
Bh0xRSrvDwxjHydUtLWE0K8gq5yO2VhwSlrJKEK8A6bRAJJ0bdmI0f8HB6yeW5OE
gn0DYUDBKWu4YaX8vhkwEhfVfh3iw2G2uVXzAf4x9As=
`protect END_PROTECTED
