`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dE6Fj9G1r6w5lsX3MIpIwYcjDAYu1dX0cQMWD3dddr3uIan8xJBuP9Hx6qKCHEVx
coKDfxpR7ofHB+bQL5MYUpQG3uQ4pVmxR9DyqrOWgveJmYzWf23VxVi7BIPoa6lY
0shL+6GgF0Lk/kC95nPak6yVhifyUxOOgXsPt4o+Ydmb9/u/TCKf2wHnWQI8gJ6q
U4TbFoKgJEQJPXLR5d71+hlMNuPnjkBPilq9434dL3qXNPCY3xhSyz+nwZLDy5gG
K+daIyTI1bWmGB6Gsl7k1pLzSPwnSFi35FaxUO6Ef7EwQyalpBZPNTZtICXHg6Js
HNguVz8tZkTKWv1XAWcEBcnCySXe07QZiTjcB5sCKEL5h0X96SaAy7mdEeaHvw/n
qf6nNnsz2j2mAUrUTfxWIKIooOb07jT2cVfsf3z95vVgTDD+gZBvL1UL3TCMD+iY
sh2ya9r8O01VdJjHFI7h+tSF3mRdPyn6qHu3c66ELbVrAyZ9OpUF7Fu1fJGbJLx4
bjNN5LUYk5ZIfyPY7LAEaHtvHKEMsMlqNLgxijzNpEWh2C+GdwCqgg+NaEzeUgJn
Y5TTWqk6lx0gBSQtoso0aa5fJyIsOQQsf/kbDTVz1i4=
`protect END_PROTECTED
