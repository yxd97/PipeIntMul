`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8WUsXhhJpmcNyl2opclHv+Oyr+Md/zEsdhS2+/rq1yHE7YK5XS3VHKyl0pVDcydp
+YsVT6n+FYBw2aDV1wVpKylzre57QMKm5EfleTKxmfDqcbDrMh51dRkrwlxm7VGR
gH16xTnq925wF12/8aGatqSRZa0kDWkWov04mgSeqoKzWqxUw5LtoO+jwKmKgPgA
3K+mpSTCkegBNd6Tniudmsp5l6GYEhmYRE5Q+dpvoCZjO4aft8YZ9wCpAhkcbLjF
vMZRevTw3sRiFYL+HF16aAg6cw35Y06hQl2PDzo9D5Lxh1xwTw+A2g6S6PZcWmun
pagDtmWEnRBdxTurlcuJNXa8K3DAt6fcyHi5JEoYZ2hQkHrOciafMgucU9SAiE0V
Fc7UEEy/n5nPGrZWqoKzQT32OU9AK8oYdwdlIUQ5RUF0KOzconQY5l92hjaorPP6
2psOIiBinx0IJ6b3RHFiKe+LLkPQrh4BGv7rmu1DIA8jUamyglyEsYh5zaE4ST/b
/CeJa9LqUZzi0eAeiDExy1/kaVnCaz0EVpj4VuKhmVPtUrAhfMJcRjn6gS3cPZTa
Yr/LPCs7gZte/BFXG3gFKxa2e4DoUreVgsOkyZRhcRYF74XQlmz0VnrlqHOcljqR
fhV3p0m7O9Va0efSWySlODhOlTk/ZA/8h5Oq2ovLhhAXvNryBYAg+GUtbO590gvY
CMEQAf/pTHP4u0yWYCIKxxSkHHJWevjrS9cXj6LHtp8E7VRC8pgTLFaiFQHgQSji
0X8g4GFbDiGfwq8dzEZfM6EGhR7ptqky7fPdy+76PBp5YR+37Vpd6RDsuiszFWkq
WB0j6MzMdPVqu8TjKEorAXTLGqqGt3vI4LkSEAoml/Rthtwc1CmpoBSniERyBNnb
djOhJpf91yt32lODy42zkxUmTYa9eEjMwhvQ5IcYBZCTDLOIa7RLlFqelrQZKzSt
V0p9glKA2jcq8icvAyTMNJB1Fc3T75NLTyoKDl6kyJow5eL34NjR2KpqoW9xNB8Z
gIaEKXmWwX9WZUfhTXk2/NZS9cQGGgpf+NnX0o3MDS9QWpWV9hO34jZVjQJx1hrc
HukBcNJgkQEiAuSNyQpciUN+6lXhH2nmVsyrm0mTI7J6yXmKAaMcO/XioZKTpVAd
YtMnPMu1/CevBOxURGzA5JQpmiJUv824OlRgr3x9BySx2+yofgOYWySaVVAlhgCG
KZ6aHkNOYx8mL8hATfI7vbeai51EwIr762El6vf9xldPnhjig1rp8oIT0UZZ/mxF
rXwr3xI+L2RG7dRGiF7BQ6xmQzM8tsUCq+DPDzoPkmje2UQoqJ6i1ymfN3u+Jt91
XN1p7NERQwA8tIuj7O9SSiy57DAgXKa+SNk4mUtrN1cFqa1SSEHK+rzKtvjchBO8
hyE1kK4KjolLVL65opTwsw43kZ0pP8Gt5YeRrqS8x5vytPCAdbMYkkUEIqJxyncd
5rZZJaVep6rH6L1WfgYgCZ+xUsDCYKRecLISnDQS2WydsdYRMhK5X25J2iM2qfhq
ErHCuTZ8ecN2xt6KzKg5PU0zMGEdeJNZtzRWtyVCr8dO9NEcSAFvwCmJEU4V5txG
bEN/Om0V8fMEoeC8tbV4Gc9wjR8moEkwK7hTkiBZFA4ip/nWLqoGpG2+4x5ZX/xE
AqomRgcuVq6EZmoLEj0lHeYdWVn3jl+z9D+bTletl5WstrPUyd9xn6rvKiEdZVe/
B15fA9EGxAXnUwi7DCmmvO3Jy0/G3TVmq9+mI5hUUoN2wU0jfpSwohSFU5rIkBCf
CHrek7QPazw7Zt3Aa6fapJ4NkPCy5EnKGsWALvuRHV6ke4dUNyPTp+im2/u6CkpL
9bzmsvbgcvPdIJxtTd50dVkMqFMiHXW/OLCucdJGYPHenGNaHza/rU23Gn/ZmQL7
mhLFlf6u/B1I3izbU79bhJFS19xzL7mQmJsl12INi2FbOrBhNkOiqUp+octAhsRv
mY/lBb/ftdoiHUK2homRjE97uao00y6HkDMVQ6iKH3TqN3hJduDtZoQyOEENyrYg
tgJ3WHIpv7Vr0uAeiJ5lkmtZBrnHP5WqJU4NkwRTn5T86SDBB8Wa6DxjyKIqntv/
zM0PKxGfZuBvi5RKFmhqNknZi5anrSZWLiY1I+uWYxsP2Huv/bSQvknP23cGgDwB
9ddJbwf4k+HX+F5dIDk6voIUobowGOIkN/bZLYD8TSKsFgM4dXRO9lZPuYiWaEIU
gBP72qzwvF2E0+K8IvJzXq5ZpbjpVwraiVTRQKhHxcTQ+R6JbfckOvZ+bXRMcALk
EretcIgQVJhC4xLE8RAnffkIOCSlRy9sEOVWdS3x7WrQvrhzdFyg/3vwPBnqpIyp
U9nGDAD1CrgqXrI+V57lGE5DYfPgt01nH5OBlFDS2hXtP6FI3JIo3AIIFLLt5U1D
0UyZu9ARqFYEVMeKcQgf6YmuKMqf2M+IqQBnkwrvF1msHpw4Vo/yOXF32S+mEgwf
mRJ9J/sdSdH3Kvt00tCBXwgGpKqhHEVHX6zbolyIbQXNeNqchcgJcbNWZejJIHkT
v3NpTb3LD4UnwmDI9e5RTEXt6m5+kyfJri3Cx5KTc5qIiCNoVZNIJoHgidyQCkM5
h5rP+bkSMNiMqXAyzcuLUZJslWJtjVZ+EtYPUi6c3N8K84UaFdnb5eeko1R8bk0b
xbDnPnc8ntP0aT3zXe5AJOGZU9iydiA8cEX2lT2mJhwnw9aghASdaFWGFj3d1Wev
0bLciScMj9TwgYlYDjgH5v3i5X5eNVWTJXTrhm+GXxdBs15UwR/+8/loDSr7jHhR
gIE5xJ4T0cWfl1YpvHwIL6Teo31t/2En+Ka0H9WCG/EbNLiaoFz2ItvZZH61zJPb
eAovgAuwElzuRHZIqQfByFPII/F0xsPPfTMf2ul1KZUl+jGAnuxR/Uin3/93CDGS
hy4Rdv+7sG70VuYp4F0llTnrxQ2hErhyOVEHLQIAt8XxPiFLeoxAg2kh7Vtdr9Zp
n0uGeHxe7ilIfDHWngciEErhtCSQgMeGTFnpCBlAnnsgdGTAIqajkCiUkmzvTGLr
ZQy9EiYCxpfA92lZwtqz/srOY8fHEgpQ7tJaEiY4JIXPQ2H5Yq7KZ7hY4QrkR1vU
Blyyv8APe5v0nWdQjg2hn+AawwlawAEAkXexuIshyh6JnWCGHI6/ZzfXAmz6rVwZ
EYJPXrdzM/0VfWwYqlqznmNK6H7rlqCZlk+/PKeRMLkoWcv0AbT06O2hTPXW81MR
mp0ZmRmRj8Rg5Pl0dtIKyRWapouGrXGldQatc5Jc5E/3e7/Zip+/mTsT18ZYd6Yz
5IGgMFOgYFIObW2o1ySS4p39OEUJQARI+vw7yDdcLShacB2FzP1GGaFKte1SZfTp
v+D6YK7GuNgS4XX6JY71KkN2ydrc1tuBX0rfs6HllbKCDkoLovUhJo5Zvk8Dpx5k
VLWMiG1HR+j5RbYBqDv46VT2JBJBOWJO9po0JWVDR8UZX95QialqX65/2bEBidgE
MDJqxdwhIvOgSnFcfM04cI8h7k7tDDJB1bmCHe47dEX2H2XN5IPsvVN9O8s80MaW
`protect END_PROTECTED
