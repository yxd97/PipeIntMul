`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHSoEKhqa+nUcV+WpRvB4Z8xKXbGYHG1oWpgZvxQ720fZDSbNlJGSX2axFcHbRTD
/dJmfb31S08N/ktOnNEaE2IPngUYJw4eKKLPT2AVy7SZKHyQTfiPbWQDZoxfWREP
i4J2r7jVEEp1cnhn7P16Y2efCZE3lwXvXTzhh5DYdjPVkfhEJ5B/LAIpBhC1eqCd
LsL0YvlXXa3o4kEaEzwMn3k+LoMR19S5+nIfUcp9jOX+GwsiqTqZS+CqaXEIeY+E
W6IeXIGxyjKjXhYjoO0MudtaQiOl1/9BPJBWYhgPROZjHVeZbzB/7dZtqa7jNb39
nMrx4RvU7Jmj9g3npwUSy/cEDBmKSMas+5jdIvD18kqUVCnx+ySLXu3CXeDXjD5W
r/ExD29K8olP+HtuprEcBnHqneIb6P6ZSXw/IPAPV+8Swbr6sDN+iBrE1APO4IPV
GYyeYbTEd7TQy6XEiZMP1I/DRECw83uDkpboqYDuPKrm+G4X75botyfA3MEEJY4+
x6nVpVYBiAtqfTuRrpkdMjqQMMLNX1Q4RN1cvhXor0QK+dn2JMlm90xR+nk0hmlP
HviijnugKe+FFEvfMOViKLQL6dxbiG/c4wszeGuUXw4=
`protect END_PROTECTED
