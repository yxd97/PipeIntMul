`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3VVX2WQcqZeVWQm3L2wF7lkFVBIeQc2McGz3G7IfsHFTN3KVf4KXAI3Z8iy9Lv95
qPlY53F5GpXInU5hMq9TH8C8Hs8pC1R/wP/uD8FFr2uUpHPOdQ/7UO+Z/2J6t9Rr
nZuxWBA58y3O5znEVQ6Oa1ugBJEjPtnml/A3UTyCu4EQi6cyukXKodVoVw7065Gy
eZyBvo2x/U/HIpagvc79fDq4oYyWpjYDnpyKMj0iA09ZO9GaiAH5AjeQpXt/pSy9
K27lu5+QkBwVbvUfwQSj7ytPG/w5Czq8jXDwmqDALI6sVwRfzKf28RHbxqRzzRBB
XFmJx750L4rlm65hubdLoHgCztxDzXDYqfneEdTkxQkz29/8Mmbn6AaMecZDX4JF
5wgssY8qFb6bEhdjAR9N3eWHJihCbCYJrp7vjgV6XS7NoXrT5Y4kZddEeTnFyJJN
ipl3hNKaBeKWnUHlFcXSG2+1ATMk0uTtmzj62lOJMlGRurwdDDiyIMG/vtrzglS5
tYXLm4OXDeoAkQxnzw7k9kBT3y2AKjV9Me2WtbuVD08HaCeD6SHNdU+S3OYMZGJi
iWrS5cj1fLLLBJfLecBwWpcNEM5fbemg2fBPx3w1ajdf7YS9geB86xg9AaWFeMP5
csEZV7jgkmXijvU6s3+VQoGTg4TfY3G1zZbzkJJTRIbpRq/OWuDHrrV9QMOBkCjj
vdS9H6kVN6IM7kAfp4bp26myqtwFdK3h++Qakk9nHoF3FpRAviRqbyKlngsGvv82
OLX2Koxa6O+2gWOEVN7s54najJVF7u4g0qrpPLNlcKjjYs4H08CL0omxHuuovfT0
`protect END_PROTECTED
