`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhDoneKfyDPpInZ0zO9t8i7df2KovNX+LYIO9q5E0cMMKz0pRPDH5d0YSMYp2ZlJ
rRHcpl7pokVNwPSUkQC1J+NPt5Ouqq7iMYRkMIiTf+25UepqeXCNrdimAy88Zuq8
a8a6zUi4qoFD6U1wIG6fVcaf2/KniriapZvDydcwxmkWH6x0JexJthQHJy0p5hH6
Ibz2bP718/jx3eKfX9kOY+FMadDCblwZJPXRertCWvL8NEVduhquoXHcvy8Tz8pR
GZrD+HZgq6XWkWwZeuotNx16p5C78wfR7mmUvMKwFrOQH2rAcIlLL6ujCAAnuANt
leyIjEuC/QHgIiaSgPH/2KCj760PKvGZcZixJx/9LFsjtH6A1Lb9QjVI/z+mQ6Gw
r9QozCcnHVFhd0BaGBMQQxGe8hHmWloozb1s7oZ4SoDfywiyzf8sX/6DPEBOEpJS
7fag1C9WGEuRX02LomDT/ujO5SYMwmb3s2/tZZKaVCkG6tkS///GXiCpTRKlalTk
PP7biebr6htmMNVYsdAfz8haqPCcehMXBjyFvCgEY90=
`protect END_PROTECTED
