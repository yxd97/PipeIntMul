`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXubQBasMkoLP4sTTO7Bg8ROXkBkhUa+EQVRXJCiaGYLVYb/gmhjt6Y7TuiEsfik
LiMym9R6YUH2hRd9ch36hHpftWdpToVzEV0x1rdCSzr7WgKbXQDDzGrXd52q93zY
6BqWGFwegKJUUH77DRnO7PpLkSdl5mPAgjCWjXUpy0duSMQ7h1Q1B5c/dHGpmBWz
WlBkEaJoY+scRsZ952UE+9bE23kg3JYc2u8mdKzIbDKLriQnSHs/gSoVbXL37Bk2
QkqoJhirVpINs5NcbrXFmJTxwqzC+yVy05X5DiSrOQBhrnLK8dVfykIveiDD1B23
Lnw+CR9FPATfG7eq1PQkBgkoN1J2jC8sdcXKwjwvWnsoK3Ws0d+6C7o0xi8Z6893
7OqprGxVYamBvXAZi5QTM5m308eCm4sGdwwQg7OfB+ahDgldr8t2k69/SpDZIELM
y8iwLMrXJIUEXZv/TY4bdZ6HSS565B6majAzQvWH9jKagTG9hXTCSAgozMB9ljtC
0AU661lZdF7S5sqRPyhL8bmhzb9HDG3jSDLY8eZdOKt9djuABnAE6NE2397HlBmp
M1RJw5ioFKoS5fVKu3drZs0sm44eyKXWGcwNvAdVbqCkR4yJ8Wt4gtpRqDdcG75a
frKbGoLM+WNWEEkl+zrjsLSsOApgPn4roD2J0gwGgLfQfabeoUzkohXL5gDkphOp
CQU9u6nYNiW2EbBMiBJwuSw3pOfPxgGbzIDvDT+tJj4=
`protect END_PROTECTED
