`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ESBy9zaXm4cFV8spdnTgxLdbUKviz+yGutm3DPIGHFsSd/YYb3bRzo316eg/QQrJ
BJZaA4Qrte1NqI1OGUVDZeL42769/ItmpOWxT+FdWkuCbqiKuLOCiz6cpb2+1Cj5
f0hk+4waFJTVVxRLlzHtjaYfDH6bWNlFLQfpd1YFO4JPj15CGg/7FuRPcAbVblsB
KCkDKRpFafaDhmTwHfLPFE3WL86khKFYC+vKZdcOUo8g+8xM+rJi28SnSGID8ogp
yjwM8IJ39fc7lalGZLCPbM85XJ5Q1rHgIUJVx5hB4/UQyeT6JoqATyl1ffiSsXWl
Grz9HDCvKcD+FZ6N9sIwA7RUfxooRPxVv2E1rem41JI5raqDJ0W99OZKh12ZKwsN
tBQf/1IVcvzFJPrdWlgUEZcA7OIh5hEa64xyL06GphGYOp8IOgjrgFHcRneupqxo
t7GBMQ2U3FSmOpgclTVc4xebY/OjjqiLmTnLuhrw3lP0dT9YU1CrEasr1GiQVPgQ
G4ETX6laac2TPeCQYmHnR23qipS3mZL+4legHpQAsHl6cMxJxI6L2imFgq01JNU4
luc5GaIvv9iCllBgixg4vbI3ves0Qmn6rbJHWyuKH+1yBhW62CAbHXY6Sd5EgEeI
bxUBJU2IL44okxAp/hRvBn0KKstsaxTUZbxvkKv/t9jXIRIl4dY2E3vu9tS0yR+D
5q6FZEgZsxZoPOpNWssue3FyxWK856esh2aGqDGNMOfPKf9z4Oy7uY/44wNK7V5h
DyBZLkY0PVgoHMmmAJz375ebDS4MmxeoH7YuLUzpSHfqnHLPYPWxeCW3StkkER53
QlI+1H6EzzPqu8XMNwLQk2JdQ+XK6jwOIMK+7OhN4AjOyh1cauMzfDBkX78gdKgu
3e/GUXcYOEuoPr/OnafgH1p2pnyvG00TR192Pr2BcrF/scOkmZlzx4Va1IqZK/VS
TvqGWGxPLF+Z4cz92mK5Q0G6tsk/6rkfOdXYmTudH6Z+2iMU3fGopTQMqqzvKPRQ
CfVT8SfCNm+VpthQkZSfSLFuAWV2hK+0TsoZTizxIvmRIh5lNq0/m9ZEniizJKX5
N4iiLJAqZNipD50xAxzUQTJdX7GfD5zVYRBBEOpWQd0KMqijEH7ZwsgZnkQAvaX8
1iFHLve3fR0u5/t8clXaRDNg7K2/iv84pMT1nK3cejS/0+qvm1ldl2Tbr4LgJJS2
rqH5q2iadMgWgLzADjhe/iSFNDHhVFCXEZyWjkfv110zAFY5MLQ6tCfOJ/qOt7fr
xrhvD9+EE3IHXf2cRrT4cwjBFIlYCw5ZjE9iZzCCvGoZg4J1u1KkyAN2ht7BBURX
KWwOdNEHChmoK43HBMIsEVlBofaNIDESGP91q9I3fi2H8+gr7fDwv58wYjgZdzpN
CgNm+xKgrafRVilz9fqc3uK9UNhsPO2evzGUzPZZNJ4L7/xAJQJYiZfpkISE+9dy
lPlKIVwdRMmlsbuDGTxW9acJE6tJxln238mI1GjzdihJZ8b1i9Px8V6loejO61Q6
6n7U83UYRm7mA+VvMF+1r9bweYGjY4EWyEtNbGkNTlIeP3mpVCIh6CzIsbidIKMS
MBU7l3cJT1jmpcp6rbd4vHfCB1uv746GRDlMt1McZabnbCWZkfLSn6w3gtMV3+Ya
p62Da8qVcNGYUybSusfE0TH42ppswt0ku+BkNGwLRy3jyWNhn7BNyrFCPGF/X7SM
mduxBwoCJiQnX5SBPVUXh0tS+O0OFAKyVyBmAMu1qn4qirPUjRdBTmzkRBgcy4Nf
5vTdIjG/841hJ33kUd13uMx3Gbf45/FCQV8xSLb1TBJvW7Tkc6gINq9lTpidMZVK
mm+b7VpaBSegJv5hgW0+MozbPXH6b61oncT+nqKseKr2UaEobCRpH8Q0XqtfHj/H
SsCiBxWcT3k2rVvhRSgwf1dK6Xl2CS3mjzDyfE4lRrXZ3V5TPd2eqHdJAD7E7iQ1
3+ULZ1SwEKWIjl90lGaS/rA5t1Ox869SKvB/zMBNoe7u2s/hmACOyCU3BQYnFbh2
nHsrHsZXvRIw1LkVqFNXTW25BA9a1XhGI28EJXVGLYk9gLGos+m9DT+cuN/a1rqx
7Cg6cVTPcfYwEMiR+uI327jeslMXQXXo8DhShvGDKk57AKjBfsT7BGVGS26n/ot7
8LkbqdpW6wFfnLfUiG52zHKqrRlxOD25VWHmB3k5FutT81OYrqQ+d0ZMIr8ax1aF
XN/TBtUvQoOhYUlOWzLtIog/I6xAwSWsD5106GqUeIf8cDKGAW1QelHBIvN44FlH
bx7G+Gm1BtWJoF7b55O1wNOzBdJR9ltasDY6fy68I9n8t6vTf3sWv1Il1Qzu8gz3
PYuCx2jEvM0+ApmmlbLtd8O3MmmpJNkx+vzHZSTPQEpslhDKA/YL+46QYEbYL9IV
jXkJ0bmPIa4tqxtext6qFG7ZPBjZfVcGqfH1isDYwij+yQ7VkRTwxSH9Gsa+R/fn
UCscfvapiHhnaXadyW/whD3c9rM8RIZ4VYCoMrvOu10If492M6iazpDnmLM0Sq/Z
+HL5F2UXxDz1Nw47Oj2IVWs9k74MsRhYmyujmS3Qe7HQ6H8LJWNVag8kIc6X0ZJP
WsOob6Wdn+tt336vkrzH7QpDCtqPz8KGrPT+mV/qvdu03nBAcHDsFbmvbP3BMhHQ
T+pPiBZWsPub8n0RQ0mhLOFCmNTldUDwA+fka7aA52fkb1orI0DNHFYdch1rqAoO
tKVZqyQMpNkAIbyECK+tzB4rngpWmpjDUjsLOhBYZVP3ZBa6LmCc+9wwDBeDtPzE
E/HXYDsGDThuUT6Y3UkWVGKyHzZiAjC4otgkk5csjD65RuKMxZWwtn33jcVMC5Ca
GkIimyF3jjX8e0hZDMBgUwIXqhmWJ6YJkgFcuV5Qy2NsucuMJYafBtqDPRqCJL0A
AzQ+dDPcqj/+LZyTtqFsZPavBr/Xxp8mOxyXdJF3WCy1YyJM3jdkSg+yv8b62ZxJ
LZ7qc8xrMSjwP+UenFr4AGs3LQTIGGUcJrNDQGj2n2jjndQUXHPSf+yc73Rhlh7T
/wi3bFQd6RuWgNLFtC3VzyuMJd73aji00XBNHeS94l/kwCJRg2Q9eC9H8fQ2Lxhm
yfTmiypfbAhsSRiO/F0RJW1cdmVC4Tl8RoMRYbJ+pLVPiivgBk3lvx2lUjT8f+lN
4d40HUfrZLxq9nfVkfNDmkQkHS384bbWXVJ9fTn90xNrW6HMCufVw1t8GRubFYf8
l75fHV0K1vSj0V2wmNlXEw5I/n44TG5qs0eIwaSiydf+NMzZUIhRyFe7UY4u24mk
voQ2iUs3FOwzU209gHiwefD5kJe62u6C2FuXWUOjYheP+uRSbFIBcovu8W8oUdgm
X7N8oT3QfKC9h94J+0heFg476ng3LpXttQSSPhxSU5c7Nj2wm6n+Av+2r1rq2NS+
QbqEYFmDPaJR8P1cNvgyx3BkgWdQ6QYhuppCDY8OYILJ92VRlgYJiPIWYTfldu8P
eXIyh23D6Jb1TCNRx++OTIbtMoI3WayQBwbpFxV6zflTV6d53411Z7ocQREu7BFb
aRTASlo1bKnDnLbMbiT5mFIj6rDANq5AbpTgnEWMlPHlPnHD5uxFAifgFDk0zmw6
rINq5anltem+/9W7qKjkzZiZuYGEalQLr/pUP4PTYajbpO7BU4jSQcncY5iIu1+u
l9ipv9vutFjcJQeFCqU2lxONbdH7gnye76Gu3QnorYwSUdNmzgCNoSLCZDRopJWb
DRu7gbzTe/rxhf5zF/byHdP429ScyAdjeHyVJSfxQwoBCbJQgu9LeIwy5RH6TL+r
JAMcPErj77m9TnrRQ4j0B63NGzR6sQhkBHjIteVi7IqB+tftbNAjW9hhIsM1AbGB
+pQfGmhA3KJgHn6S1G0BfzS/PAHQhxYRfaScUFnWZQfALQjWhRfb6qOKyDduzls3
X/YCnqWoUj00M5CDegs5RE4U7YEeHrHrQDv4t1ff2Eb/drd1sV3OtAN9WM2ZRnRL
mpvUwrlDfuDtpQ1vPJd7gOQ++iC/ZwqsOGaKqanPRn6OjhaZ3wxcS/p4itRMoyng
r9KlBsfQfE7mj8/LNpHxCR49ALStpsEdPzyvGzOTFOMeipIcjsWK/3/A6ZrScu9K
qdg/R66xjnf7xKafHTYvDX9Scbe+7pqFIxvx1ArB4NFqxnH9typo6NYAz/O89BcZ
+IUjmC8lUGWc+J9zp3Zdy91b6SeDgErk429jHnBZxq1GXU78/Y6oGR352XT6/6Vf
D+sJ3P0/m5WdkdCRt/XiA1m358Is8nuyFsVSkxBM2CgffELlCIfIp3WGRWu3Yc48
Zb8IQ4004QS8w9temoRfeeM1OJgUjb6c/HkrfC1U8H6TY+XCqcotsk+5USYX8Unj
/9MUfttyHYwHvZPaKfTMb8M05WG/hSOhVliirzMDsI5IdtGSdRioZlM7h71geGgw
aEqEAUIR8at8Un6zrqbBy62RCj8e5XmotZDbe+gsGYOptimhf54COEW1bYKmEf86
2G1msxBgN7JQM4mYCXQuv+GC7D01TfMSYcDmwGdT2ilkNw/Tq4F3iC1XR7BJVfQh
PF59UXK7OtvyfkSIdKz1N9rErPMVudBg6DQFSmi6q2fnhXLo7AWRNNubyyzX7jfy
DKBUNyDlrg2J2b8hs8oTAE10na3FCP8olZdLUbOoOwvCDby4tsHz69B1pGqW9Q/W
r0ucPhfIb3IPrJPO0+6CFrMmMD4fjVdynldD0u5ViPgioNWoEr597YU+DP+nG7EI
r7Oogo6VTTJh5JTkoISrGOFRZTDUsLWICR8J/YlA9/oTbuAPKSOZhuKkfizLocLa
iZI0/lt4wSZutmKb2Gx91fYJw9MH6kfeLpyhYxgFYwcPPPRaCwkEvaYPkBwLQJsR
JIUKQmy0IQMnCuUsAO1KbpFEv0QQDMuhU/1zHRuXAnMZkBnqMjtfg1WIHZ9RZ5Ya
6mqoaqlbqjl3JCEbTKGFHOKRp7/559NtSEaQK6jfKrBE7Vv/Qd1umYLFym0e0hkd
+pSsST6AAXKI3DZYasLlWmw0AoraxqztButBHacvMwNAfoEQn0g0M/WwlZHTMT2N
QfqnsxBLs8sgp71SLlCVeLe2fWI5ciag/YdOaq8hGoIAbh40n/37VoO1Ltg+X1hN
vrdFHv+YC1SA2KBY/4uOnvbuHGLoJczlJ8pmRxIeMK1y5/D3VTxC6Tw2L6pRtNL3
iSZlj7lLe0C7cNcN6klp7SZeYzX40d8tukTArolbSDGTh3+ITu3V7ZxW5Nc6y71k
dqqSFuq0szyaM/Ms6eBiUbMWM+LSkMvuLUn3IS7ijN04RrPzXg+rwHV3DmnS5lgv
94k2+iVZ8rKQfZstvbVFy89+c8Lm95bgWxBpePLH+IhCCBb/xdbaK7P2SmsyxwUd
qhdlbjk8bUAF/JOYK+ws37RNor9FCCovFniWgGgQbM+y9RSijwux9Mzl+UDkcMOI
Ceid9201v3Z1ZrzSOCUekkTZdIeJi6Lj1T4QOjl5W3+AsCZ9eqt5qJvzkHseZaRr
WpexMXf9bOjqnnTLGQcyHiJqdwPU9SnX6swshpsqaBy0WwmTcgQhDj+8UMhhA3wU
z8CfBVcF7VpJVEK9a1QTTGXPVaUdYLfGItKawpRaLFiH+nqD+xuoyqm2baimXR2P
GP8Vjl6UmqW8+ZTFkJEe0mcr6Hs/+DU/qzM/60mNdCIfVj9jH4NUchf0cVmFW5/B
3GuNXpFHeMxyGNvp/U75P0xFgBMmEEOZ455lu1kZ6M0p4MF3P9FsloADBt5XVfvD
NYGTp4dTBfu0upUIQpcuqK+ihyc+v5u4mxTEXHabnTbAUCyT4tWnl3jQL3APsQwa
t8lXGiC1Kik4eI+WK2uuU24NkVRBz3BBmJOa241qLkKhmoJ2RX5p7+zm9n0IPc7l
QtL804xO7SASmi14hexyHE4vxRdgqnx/u12KvTPSrlLzUEkACm1JkhomA52d7iED
rzDKIipW2bo0ESJhXYB4bd1lsnD61oL4tc/Zh8Ig6dPc2iyry66Lf6XaDxAm20Y8
r3f7GaGbE3CnesbkIizUytVavSV6zJKoxDPhcNWvgenA4AE+/SrZACA7/UYvt4EY
TrQITZu6YhvbtzMd7k+tKpDoTgG1pjKmkBfH7u2fEzYGAB6BVTMQY5HmYKq98hdO
K8ZSgAYhjjt+T0XmWTfFwIP7ufwBW4R1BlsMgbKMs6T64gMKDjQHL82bv7WOEUVT
Q64ijHib1nbLrF4BM2pFVYNpXYSAeQDsYSI2Id7UPpkOAzuzn6PKsT+eBkpFJtYu
svVTqDkx+I4CbhTIzZy09DJXeKWuiAzYZ7JJfthcV1T2YaB2Sy5PK5eL8fF4n0gc
xqPuXGY7MRaUGwmNYYz6kX03vk+6TlbBHO/qgRw0ZJx2RU2SaQJcnnUcMePtbbrE
6/pcqHu+TPa83Uu3qxBmpKU0ae2vfPa14T+BHBgpzf1P+tGQalVOMljO37K/71UA
PlyH6oiUUYJLuF6lo91GXLvx9rIadQY3b5LgrF+UTZP/T/xerRdm+Eg8+Lwevr3c
19Z5b0HlvJUxnevrlP8JQmhkpikG8kmRjAiadTPm/mEO6pvp+0RGJb4X1XCONNAa
YxZuyL6WracNu3P+JcnsK3iIAjZTJV7NXkYhmx7/b2KedWKgxJKjCurzhlJl2e3E
tyR0Il7fvIERMIqEmUKzyrsDLbY9LnRJfivj5fT96Hq7yQnmFp5ZTQZGnicA785P
Lb116DFVGLTwzTkzueKTArvz1UNJHcJbURtTxRnCt9A0W+qoHqLiNLJvZ4sBB5YM
dBsJ2Yl+sqPJkoTXox5cOZ/MhYxAac2iXRTZ7/cC5BddA3qAXR+iDJJ4RiusCXgw
x5garMj9iHaV+cobPxXs0jd7573JMmFn6w3a7iTUGSSiMTQXaHB9ZNsE0P4atuWo
S04b0Fl5cKIgJkqlWetrI0i+M/WGmmKBWKB37Wit37RKLz/yVmxHN4fB/KjCRfTk
T7haUPPq6c7cChTrNZ0QKA1kDYZ8xReZ5ZkfYU8wi8buB8TeLz3Gsgh4mQV/OjpM
GvtWC0F0Pe4JnBg1dwL1jDpkKBTbXItGbtL/vipN1vGO8ikle++n5hHYHvt3/9Ui
T2r93C5FMTdYJyITthUdJnrVoIaCotB+497aIEuzRPdw6OkINivNziCfwDE5dEC5
HYSt4HyZ4u5Df3AAYJ5CDFyiRMhd6Lh22jX6Nj9vDgDzF+1YiM6dMZT6o4tP4Vjo
q+xPclm+SxEZQ/jw/Jv8PS6pz1O5EDq1pg+U/ocUEDzBWkqnbCAwqE/KrPYetyaj
orBikhHlF/YQWjTJ5/S7B4RK3DT/EBAlLUEsVsdwfOhV7WyEAbwMRm3rTYHorv5P
YdYR0Mmal4y9ILf/Ap3Zi1/IFLWQDvovD3nwienVsZkfPkbn2V6XAPxqt9BvXeTE
xkeeMNWWt+Lb/B7KhknzXWfAgEI+9b+XIKokmn2R5U7Qrzb6GqgcQ1ZxEauZcrJx
C6zxK3nUEh09abKJtxDUUy2787FN18MUw7W8hSxgrTdi35HTvxOO+1M7aZbf84Zp
CDRtkIZOzsoW8ybABk5bChr+O7t8tCXa/Dg/e/mStzhuOnyJOpHOWFB+JUTzwCq8
hw+OXKAiAJtpcidH9Cgk6RrcYYdjaEsTNj18leYY6dPuuNF6+q84Pw4vOLxXcoSH
2zhq4cljulpJf8Qwd+XEr6FF8ODsS99hUPW0kVGU7rey/4VJSULnkr9P/oSK2cpI
4dGrptM5C4fUm0WdFbjCN3xeFHmJN7wv0k1lev6C6rvCkJVrKocglyYHYBWitG8p
uu30pDIp7LVG81ZqJ03xKW3y8G5+rru8TQq78MYbaWXFBG+fautwSx5beNBL5spL
PTF94s0NKVa52d3ymZTuhmh5pgwx52ASBtwq3DYAuZ0Zfr0oQs/boGO+NUabAlfY
sTVk5N6eiVRRVIkyl+Euibv1AID8dPPEPgwnC8ClJN1T/jfKkUQiRUNL5Edmfkvt
jlOYbLztfpap8wBalbxGpKcX/DXtV/+fOW3GlkN9Eja0zuu5TuI5NnW+WxuqlpUh
jkZFFZw5fFlajDlI9KcYGuhU462BmLoQoYXH4gKmihC4cYqIlCrlr53x28i9ijkW
cf7NrP6ToaKo93W43mh50dBJf/8GsFfzjjxo3d3DdlCB0zYmZbl0WKkDsAvi0sSu
wmfKeaVWJeJv/6TIcFcXXNcOumVBXvpMsqz/qyWyQ84PRPGGa0uNz5x7bI9t2v74
Eo3TL0J14fbF2fYPIHYRrozvxp7A83BdiL8IyXAr4SCc16nTuRq64KzrdM8frb3D
RCrGh3zeMaeHc6VCBY+QKFPj5RHU5HwuVFzdeYPdYdixsEj2Qhhle6tUZ+jU2a62
AgVwGsQYPzZkGZSaB3naIbtmX7tP6ug2s5GrhxXOMPZi7c1RtUs78S0W7eeUYkOO
7Dm4Vh7HXDBku7S62Q7kICOOh5LAOeJrbYBiqGpH+tZxtmz/nCcDUCbYS8Jk1GJ+
TQ8AS3fYdXjeKRW7JixcdXIg0JH5P9T8IfyAaANi2xvVUAhVvH79n3+aWZUwppT9
7HZo1WG5mZ53ODtt/ZezbZizFDKhIB85kbBEM7WbWF90EGMlmxCahW2i/I1Atjvj
Dhb9AnR1d1gzYEy1o4ZZidUVp33MFNyIPblDnQLNTTWP+oqLqi0dV0rBezAkSPNm
0a75rEV/dFqOiLqaxoL1Ia0DWDHBg/a8U4XkQvroviDWwoLB/3p4K3oMtpy3rbqR
YzFaqmpCkIhocMtXhSjgZ98LHLb20sd+BX/0BLexk0PwW1Mwv6weup3I4ShVKqRg
UxzJEpBAza0mWvwhln93VI0uS/MVHV1VLClvWRUl2S56/NFy2gSxLPb24SNQm8vF
P3kU/FD9CCNZl6FS5fGPKuVkmorMCw8b5vn8WuCtZptA/N1QYZnrBO6/xLMzV2H/
C3y6vKcYaaYRTlLL6e9qLQ1kLDJlh9oBgLZ8xp0pOXdmO4nVL+BhWcw2Ju0HGb7p
+J8EBh5QjHN+PjuOU+Rv6YnBCVLgD9Yu2eS6SxOfPw5JAwY9bmuMw79QBzSP9hE5
JZcnZ5Nd0yy82P6jI7KYXcK4MrWddWh7bcdjVMsJOlrUpVhVW4/Hcn9w0yfAvP5J
BA6G2nHRUYMN/8fDtzW605xznAordJSv6ai0DitRifngzTHls3OCnK+SZhJvLdAg
1134qg/xHsSpEZHQwTkcQBV42txY33cP/thstCioMf/vYtgCugN+w66ek7jk9vaC
I33irNw6FSGjZw6FyNUMwxFu2iOYXHW6bYsu8G5R6pyVaB4x7kuo04iQMkixIFO6
pm6P7NgZgFZ3FjPdLcfSBMv1XZDy82jYWnjekd2XPbLarhRksiLxVz/Y4os5o+N5
MdHiNdZNoKHloRT27J87YI9X2aCn5c2PbxzuIi91yw3FJHoZ9Tvv7HyWhfz7kmob
PIv1GyZIuwVb7xaOp21bVFjoqAnTrpSfk149UUWQkciE1D4FCP7Jtq/hopg1e6t2
soMC5JOBC5RqJ6AMh16/betzaQBJA0PsZMzsKyQVmLr74X8JlCJNJzkjxMBj6BnB
TPh/UFkYiRgxeEEWiyAzUjs8ryFMnuFunsziIWzTEhDdI9cwv+fWul4GWeK+q/FT
D2pWLZzeAuy5PmqraZow09LAiSxpELx04Yl8mvZCWCDktrP9eMa+D/775pCkoLuG
9Dx+L11ix7jdo3v8uvi0ZFOabn53zX1bIcjPfzhfSGCv1PSVyJuBWplCLprETO3C
eT5N7PxBAElgb0ARnaR9Ifm8VWDH0uMR3FmcesXJBptSSrjj9V8/DMDx9gcY4B9I
PmyUrw9SEQwF+MJk5gieZ/GxyP53K/EK58yDcoXiNjff1a/30N7dwsRh/lyhqUB0
fXDCqgmWxwhu8pTF51KM30WHhCrPMs08Wlpl90dTQ1qLl74TYbqV1eDm0i6z538n
JPSX5KQ+TADKHwl3E9RtRQ0p4dYCLBZVwb6FfOQ6020JIp7KrlSaU6wENNK6bnu9
Rq89hSqiop20kCKONAa+wAawbmDl1ko0Y2uZSk0u9hCRRYAYX8FBbovLdL5jNmBZ
IBQpoJex3lSFN+AAiFIxx3cIgEhCSSKsuYIci0wOxEimossifQQEY/ajwGKYl2Lo
ErZNYxaK6ThGY7++WKlJA5ERPJoLPVBLqXI6SsraU4ZGWxJZ/V3rSo1hQ0x5McMU
BjJDRWC7FaPLdoPyPbIazJ33nKjNq28wlTKVLj05OVt/chQkVhhEj2rR4ujTbDd5
njKZYBQGLv82nTxF+qzn4QUgoH7Dq/nEx1VDMPH5GmHgcS4GeH2iQuuYGiwVe+3u
T2DonBFAWVxwqm6k0tib1S+2TpR2tIO+LLGrIfGITFhZ6SUKBTVIV4cT+/MCu35b
pMrnbToUS0TFnQ2odRM7vxwc55yDNbpxJYIJRTnoCeAvqTGZSwmJ6WNI0JBp+mXD
A/y9f8qloxva8AzYIwR1Htcqdlll/16uD04hMztf/s+/1V7IjmO2h+dFvXpgm4Gc
JDrBWWAZuIlRVoKljNDF6GCiwAoiHWD+y6oSXEzwxO9ph2APJiBp+CxFynVmb+xf
8ZG9IJ5Kneiax+VrfDZ9m50aKe8KoD2Vz6xoMoooUdGl5RDbjQjsJaN6dJAdoY0a
cAwh4LBUofSCJLtS5/Leet2P7cTv0ZBnvgpjDaySCri8ddZ/mdiArC78G2vBLLq+
84BCy+r62GNlkOr8zgKbFlR74ZwhUavw2nbVOj7kZ4lq55x1pNHOKUIJgS0Ksbd9
nYM/FZAr5IGnvDh8JnFa3+FVGTtJY7RfEZFvQgHeQolduJUaeIkHyHN0P/mKr9j7
+cN7RhYsDPaM0hwTxdgYIBSgr2B7XqIaWajBHEtuTCj6UbdaayB4nZrXLSrKNunW
WHp0qpFuM5hn4bSoaO7wHi8cqnSvFW5mMe24HUcrVvaGf2WEgu8fb9biF3qp6yCQ
8vW3Fo0EuHgzI1hUwbyiTu6Y8Xw0mDdHzgcIl+5wOwtUZ2ErixDGarPWC1Lx2nId
Ut14gmO1Zxmokj2rT334MmLsRhWRdRpd8ivXqVdQyKIjVse5ja6oBDdAPPcmotET
CsEYWbN7sgrDw0LGn9claZyeTiMVLzv7yy5/jvK9o1U5kZrkMHVWGQGZ+AlN8FLh
ZIU1yNhWRp6gHF77OGXStA4BmZv4RuWmNOo5Ec7D1KiojhwPx2cnIVDAyM+tPNDI
jZPxH/+pLjmzobnMEKTdbbFangAeUDZDvK81QF1N9FGG8uJKo4pnbV0W81oQZ0+T
YWUSM31gLyVrSDJBBpul6oKkG6ySoJXZUx9+hi6htwBYV0A+M/0r72ZGlmIzyr13
Vku7AvWp+Tg/lmjYAw+hQudSXIEvQ1InN983NFcq9ofAZOUBAWa6wrrQYb4QKFx2
Esatm/d5mVcYztZNftlTlz+ph5wMXTdzEF1Nv3beJeUBEd7q8fkP1NMAj8hxErJg
Y6lqobVc/rVNOsCgPtr4AVMz788hkMpL6WOo4cgMk/+twUhyMGSeLvekMKHg5QKm
Q1eocNH6fWO8m2rng+aLLM9Hjnj/eOYyUJ55q0waV44mPlV2Lg3nv62njatQ1KHN
Hy3KM+pK6t3pb1I/hxhQLOxB9XZSmP2bihNBr9oneK1jGrM1AwfP0xcoO5PzsNBH
wV1BQbR3gUzaeq27DjdRY/L5kGTkyVTSt0N2Povashh0piN2+qPji0qnxqn+Np4n
BRIaxlbaPzYDvFmvWm1WMpGk2SxgVLNdFqS5JQhDiGwD9Q62h5y2UzWXj4RO9myK
lpX5R4E4dXx7R3Tzf21ywCzgczFcGiWqq7L16kKuE8T76YivgJ5eC4ns+pUYQAz1
e//8mNoAIj0l1URY/GykwReF7jtkc1LrSyCKEoUhCsHpVfLEBYn9hwuDx7yVoIrh
rIaINUDiWSGmq+TQS6p85Qywrpq30Vk6TJ2XF7pZ4fUNZ74yk205csMAu6ZIdoT3
SKul3lNQZQ7+mzMCY2Oyheq+2iI1rbcO/cGBpXaIFYp+J5qmHPnzQc2FY3mroJSY
2A37RtXdtFswoHFGMRZISrlZjUOEr1vf51yoF+DlR101LB0XFVG/WjClRd5miZmS
+hVKomh1ToubNd+U7MHTWZ6kystgIZaD7JOxdKO1LR272HtkeZCyIf8NxM+toyXl
TJ5TF33OP9N+IjSyh+Qxb2dup+QgGMINOb76L8TMiMcZbFzOsqfFxlOawSP3372T
q6rhYQiPzLtRX5+Yz/eBRD82Qh1mJH4ceuioybXfjTkvrXww8IYNqzFkd7FI+HgZ
iETa+u9VC0eOZJPLGfAjWKxKCVRfHATPZUVkw0ZtPZ1knjyU+KgSV0zpzlk6bS26
GJmsHTKlb7Ztu2m5q6gnmWEt9Vxr/s373AGlC+Rx3tcDESIKEpKi+d17DdCplBzH
SS7Ps1fHbqAOPp96k8UubdaEV/lC08U/RjgMLyhqx2AO7f0QSrT0KYUYivVwTIVL
Ge2b5PdRNV/3V17EKscaQ1UPuNZevEskLFlpHKKlPbtJjTaIkT6BnHfbfsHMCR83
nwUI4kgRXjftDvHLUvLKCq5SzxSUSSSjwzRpz1Aq2+WRe6yKIbpVtuqvf9kF9WdW
lvMaJknMwkbLCYF8P7hCCNvy0i19URB9k8pyPSG3ZNEerT21zmwM8WTCGuQh3ttK
72pULYuqyklW73nAmBMFirDEcOXLLdow69nC52NC6Jk1DTnhtCYPM32DAFfeGHni
Tu1AKC0BIaIsSjPs7jwnFks8CodZcbLoPpdVZAs7EP1+ecxbF06EWSTXOE/o9pIp
K0nxvE/P3YvGwuEtFzNRcNo5CLG9vbEVfZb53rk9vNBMoNdFfSGgj9fgvuJihxyI
82hx2c0dlBG8f/w4A90rluEmqPjxSOvTkaB13mHhtrpMsOYsTBgZ1l56ap3yJ37x
awdRNxvTVFwmVPQJErtQ98zphOdK52/zNDRtX7BtcazFaIPPvlFHNXDOAhMY/vAK
fSMI2qN/dUmG2igwpOsRiDCIW26fAffpRDeJuF48Gv8Awe5+RvhkslZG5kwzqy5d
SQqSuau1khLnwvon0qtrfefcoAuMdDo3p+1dlLw3ZhsmtzG5uagjX7t/9pRtGlbB
7dHWmKBqzTtg3AIwGqIcyICPeYMPTIbc6kWAdnMb3SQApgRN0jKzB468GqCo+iwm
k4Jh+7MklDWKjXl2FuXF2Xqh6HGVck6Q8G5pqyUpjmbBjKao0OE990KR5qyobMl9
x15rEulSayroeC5XpgkHiaZnxdz+7uuM1cEaNmlWJJU1N0w5WZOruZHuOj44JVcN
io48BimV+tVmEiAiLVfvUS5CLE/8wIaCSUuNwSHF0ndSMZohAPPefNeF4wi+KP1V
ueumzaoBg1XXaIRr+WJqXskUfNs2+P2Y264imRwQOLWVt5tIwRXuhJ1INI2mBZBg
5CiBfwY+KXbiz3wyaJ9EZb5V5wcxWlTZsjvBlPXEMWeNh6+Ne+yWy5jsJXp7uRF7
htZZS0Vus1V02gTH8b2GaCWjeAlmuPD4pUjF7RQ/FWzPV/BGZ0MwFOUvec1GY9vC
/63vJjuG0lIHkFpupm5Z2nsF7AFB6HFTD0iGDy4r59V7r4RxuTld7P8JsqpjhVLd
JfTwH3XZJbDUsIdu+1wmaSEI3StwgQJrHuiYP0UyRs6PuP3CEOHsj4waFogOecfd
tG9J2EfI7+N7eqpvCKccNmTKugbKUaFIz73AS0BOjmDwTz12YLecZf20iP1yHbNn
0GF1By7qH2KLsAkMZa5wKZG0fzKG3iTxe9afArFxbBXrUolvKZ4/zl4msIYvgrrY
YYsLuwnxj0zRYziryuOHFcUCgBq+EIfiumZzO/HuHqLVm+t6glbfE+AX0uJ4qf9/
J8jIvul/s/6MYmM43WltEIXJ1jHBFz8ErEPfic68mlUgT/LszrZP9RU/WltROn9h
iy6cwbifT2g7RJJg80pWP92EVxLpZf28R3VKZV9Ja+M9BFe98TDRcCM5mIjpc58O
9KLH6/aM1dvz0zhZ9RHk627+WV0V99+BzCx7QueG0u/SpEma1WwSimRJddcO2jie
i/JsR7sDAp6TVGpKLXypEIsF1Y1uvKElgTg0SwYylyUaC9OU2NpS8QDWuQg7PE3J
TrvD1b8VG5MWbyN8bjW+Il4UDtupyeAqxkhVsgTEVyFjEzSdF9M4k5fs3uYaQk8e
zh2OONn1XvH6rYP1orIwuFkk0IyYJEKfyy4u3pnTPdBKUmDCG9DT82xpWb/BB9cB
04d8T/Lbs6sDHQ5r5QdrdQrZB4HncfAPahNuGxnXyvpiPb8fQDcGpa4KxbB+jQng
yCVQU1Q5pTmEPlJn4K80vgeWpKhv5UCxKqwkMgWAIGle0RNSR36kLj72QibY+Sk8
33joZRcEFVMouaeEmPVLZgGh11ibC+DFlNyrLv4KNLuKcA6Lo0MJ7FD8+yYKt3SU
ZVM7nT2vEo/NSRGsAOSxC7pMD5fLoKLiEVJePoV1Vw3w3bHuYDYANbE5IT5Z7rBF
LhRp4Kel6thAg9BMdw7cj0vVTZTaIyjO7ni15xKaJgHn09JoDG/vcanEGP7DFCw7
74dtWNlxnIC8oj51vDWZnz0/5YoTmWFv9dRazfca+jeCTkNZntNmMnEamRXYTZ7y
52LLLU/2r73x3WaxL0fCwaUq4j6mXG06eqxsGwo5cZuCVpsOuBaphgXyY7rcMMW5
Qebfe52V4ibiGSy+0NaCyZxZnWzFAAzeGG54iuZWFIZXZGbf9GZDbJdVqXqmc5lz
dxJxpROIBGMGTryc1CKhQoSDRH4kPxeY9Z9dYB/XLCnSS75gFg6PZvw8SvVGxxcl
lBCf5YaMUZAjC5Xw2UzVEut7nzyVNa8ZuHH0HIVLDVbxYt0XeAPRUv/v8iPtFtEs
JEn7bIm8ooJDO97DYNFuai+Ngeq5+QOGMBT/UoYkmxJqL9haE6n2y1Bwys/07jPG
K04OpHStie1KNPDHijE2IvrBICp6AncQNk4YIJ/AM2KUtdrkkk0cj55/dZooKW9o
VjmWybtbi43IFXxTggxpZfqnxXKukN4svtqBeImOo1Cn7FdnI9vzcD2WLA/uDo8e
4rEp6krlTufsvKyYLf3c9/7NNGTRs2poRwoUTICFrbVQqkuVJ1s62qYdv6wdK4tw
X7bEmDneZ2MDPgYI0cwLMODOUmZ3u3rrRytOj3PK/vpznGVStgO/78gW/Wx/m79K
CiOZC0mNr6fYtsaXURemegUnjXLzmj9vPwqpkr7RMJ4cJvICXZ7Q3zuafx4OKozt
2MOJ2wCC31HGo94TYmQxFOr5tHNqu5mlNvkiJkV/SOediJ41wQZPpwNVjSqSwfRR
nxLaasYI8cKtprP7oLaeu5RvSeitlxokhbeWY0/9dhymbUFB/WZw2mp9izJxOb7b
dTSPiwDhrHPzR80GVOZmK1A9XbfITnVorwo0qwL6XieI7IXCLkbFkDIOg+wUFWbS
Mop2iuSvihco3ipyFFrQCok+UZUnX6ChAMx7uyzHRgu/EzzAL7Rc4JLhvsoy3tGa
tThjzUFOn6eqCAeYJG297iYdvmK8i+xuEZ/eYMXxY+7499QOeSImYg9rSfZntDrg
EsmJYY5lWSXMw4qD9RnDZP9I+6I6jef7RQtvaroQMKix87UFG4khOhIB4bJi0EiP
+64ev1KZ2k420QYZGKd8TcjfQgW1DgpyHkZRdjm8fqYkHt47MgHAPfIJcuP1R4Fy
Pn6AU2hrYXVAiaK6CFV4R1ApO5j1GSmUqP7GpwOkp3aUh54ZwXVjvJlZt9P6hcav
vM1wrAyWewbK1/Vq4sdDtrVleTYVJxbc+4ZLWdqxE1AgDhs6PjDDsSf+yQ965e/n
u0ahaJN3yos3k544PWZVmlFtbgY9vE4J8pjcClozl5682FAtuXOoArTdHpxp5+d9
Wxn5wHVjtouLzSNzIZysKkUB02OdmgLriquAnjRsRWEmw0qeaAzvxXUREJkvlKuo
9ZF4OXWR1fn0FwLPcEdL2xY+hj05rAUmzVfYj2fa5I6Faw4JfzclUrQuKUiCqvmr
DYqe/s7Kg8MXREtu/Wohx3e9Y4QlywzutroPQhDTvhDSh1ss+NhvPgZiYVk69q80
6/hFhJq4gN5kH36fYqMA6Gq2gaRKUTEMhsIvTXzvdAZK1SdaVgQrofh80Yds7lQg
MXVVaTd6xPM//3EzyusA9ZdycQZhxxiIZU8Wk1UUtuAlHYVjUH5idPSAf0PrzJBR
OtRURtTiz0ZAagqNJKdLsJ6D7lvC3n6jJDXY9wDVBw8y8WPQrep91Q6sE+HiEUb4
eVA1Q8t7t9mk60mgtGZA8wUT/6ue8o5j5FndCZc00nRu0uosKdr9Pnko1NurtJrm
Y2571YWyQfX6KqmTRcPLOntIRVOeaov6jMj1J7mLG3aeT3gqYbtIlmwAotKIYphm
LaPdihtv7wXqDBHPe3soYEj6CMP+uyHDC1j1xedws5jpKs1jKXZXl9+xv3/HedCG
S+fBw7iC0ud5qQEv4h11mDMWufHX5bqWZ+h+5ppDidVvYL/dPgm3pkzGa4Vy+mz6
HTizCDZD2PWDwxD8mPy8958H8vkLbHRI7QMAH5RtlXSN07UyCY0jPJgPDftKoPQR
nb3TQ91ysbcKOjAWD9lcIL7YxWFcTYOdJFmlDaYV7UoChKvQmF874TAJAPxjZvEw
j3YPWSQPBRD1BqV34xAfF0AZVaZ6MNio7IGFiRhEbFB+hUYTORcRkf7z7yPGN5/O
ealC2zyQoKjfseH26MdzFnLa5CDrKug4V1tlgSJdE7o92qVD+4Y6LqRi/12vXDOR
n9AFLL68mYblqimjF2VyNe+AQnPfFo2fQHlXSsDy73Lv+7CwBOUer2u9bllULWMu
xzL5lAJTZmkf3uuurTAWKHiRyYFAXOe2m6IQK5xFajwoaelGRv6TR0fvW3hWQ+WD
LSjd7Nsvftqsuz7hwvO1QftgswKhmwbdi3o21liQuuoVBRpANt/IWOSbkOsLPviE
iNqDz7IOutbPPAwLJn7z7w8gUVwRlds2c+ZoAKmRnaDKkyVV759wQ6XFlCxFciaE
2vqvld7v/2Ie3Ov26xU7R94Psj4UI7kWsLx4OPtFW8f6QWCT3IBUxot7GJXj5N/o
KFQ08tMqthvJhUIBeZtDn93eulCvfb5jrXvmldQlbYSMwgD6PsVC0372EsdJo6Eg
4xWIg+VAOnDyCnEAT+zRPccnHUK3J34Z9ew1r9eUuLX1T5XK2XY0v8e2yjCcWGav
TBY1lKJupJDpdSg0RzgUx1Z3zVjsl/2UbNtXSLLy8+HYBB+AhUDEX0Ym7Y7Hsglh
2sKe6cbkKbZ+oGdEZnrYcG2DWelpw2x9Q0eDh7zSqm1x4BP1BkUYxCyelqq1Xbtm
QVlCxbog8uztmK4MrCLzVySHFCTOdogWDOLO7Q5kYix6FIvixPVfqOpDUURGyKf2
kuEY2vvkyT55Gy1UFHB7wGVHVeF93dRs2g1T320Zn0Lztw6rcHSonplqaUG8GEbM
7Zw6uqPC4TlkV1LdnqnodlR0/sftWB7hOw5kgfnI0FTfrK9niX2P4VjVVCk1nThY
TSyP9pmulOJKQoHio767hvCitbipB01AEyre4D8ZF9vVHy/ZCSw7WuOZ0OOO69HA
nHK8jabpvlUUJ94w7oaGF4epWNSxhE9T6pRqKcwy5tCFpyFi46Q5wK1g/db3DOso
lL6N15KK6yxCPDZs7lldNbYsDbefMGmgj2YNIE15VzWcvqI56TJSiBNIxBaY4qVY
kDPKpKxivSbC/prEtFXQeHrEGQKz8DtnDKxPjisgAkcTVLMy08z7ekWxPcwpwgff
rYZ3MaN3lj2fICCg56dIrrQJEMDuIxsILsWCqjVxWzYJSxdtRsvOXpKlLmeEvRh0
HEHhzZyC1GYlJusNkvg6zBOkJmdSGV5p/KXNQaT49UFtMd4kY0dy7GUFwkUkKn23
UHQ5O9J3R/aeHHG7b3AFmmSkbrv7NAAK7poZxUfKramSKMvmCc9/9sNFwDnMNPvb
y44M9YK7X2aME+2wpJg8xQDdg3kyTCRRYFfY7bJKPLIXl3zNYoR9mipzivKQKxmo
xyobDWJm8wjFCJroL8fUgpEM2FV2BuLFDtO8I8h8OrZFGKi597MJ4Jxw1SQ4Tgj4
X4QIhV+VDAxkqAHfzL5iuA9OsCJ3KWD14/qRR1JmzhFHsXEsy3/dLeC3nocpFXQv
/fcx65OqlirraFVeab2nZ/BGLodzb/EuLA1clBFMUbYmP8Fu3gRCHZehliZUisTm
Af9A4K3Xdpoc5i/soaiP2J/fDSSwBmb67ZTcq1ycaZxJMdqrq8M9sWfmLMaQmS/E
wxfIRJyQgMThRr1JFf4LAmLfEcW5auzwWxiMIxffmMnSH2kO0A84hRv12e+72bUA
iXx6eZckLGl2R4cVTY7P10mjZmclMrZGNwZy5oLGJXNMz0cI9wLqQ5didMit1/LL
LdiHH19F13ttnuHyAUy6rcYCbGWVj5UuAzqQqHZSN9W9T+wPIa8Pvtyt1UiLjspJ
vT5uulf2zfKQCkTOvYiUQckS2kOzLE561DQM3YjbyxfUA8sbk0sZymhVWvR6lQEL
7Mvf+W8WdOD79X5lJATPwOMEmZXEBjGm3j50H3gwI42LwWTKAuWRSkO5s4J8SCl2
OETg4jaUimB6mJ3xa0CqG+W5GV1+lYxxSPBwrGzGYfWoQxdy61+1hWxApgJPVf5+
tcPoonZeeOup3ZoD1mm6nvcaUm8ryQeC4zsTb9lm5a+RRiFmLwI14hoKlNErDO7Q
q1f/MpUrjIaECOie2wXs3mEAvkLB/DRcf1I1b2SObbDyb/665tkZU3VvwtzQAn5m
BWaTlOFae9fqHf/3ogacWUmxrOD9GLaQS3w3CkxsHDG888Tz4jzQJI0+ELBySJlx
aaHn46HPAbf8Z4XWcsGgNBRHM3L92tL65Iqc/+LuZejb+cGc5cjvAgKkCGbRG2QR
8+kS4yooDg45Va+4PJ44ZncE4RhD/gwipJSB/2DFkgM4/bZmMaEpbKTQrO56Ri4g
x+kvWHP3Sl115uytJ3bxxB9Os1OIdu5xRYo+8M51JLopzBzys2WO9nw/3UrUDlJx
4BohYWZMCK+avds67FhBLaG+Vi2p2C8AvdpJDBPWCJ79v6XAJpz916cd+u9X1BiA
YI1xu9m6ELzy71gfidj6Aj+eERqmJtoJpYbMdb7mheM/dW5T9SRFMNVwgFNNieqp
XlZxdQv04L2f7SaYYIMn0LnXdzpAi0W/8ZBYgocgpIQRujd74urdqfaBG/pT787y
T66Khpcq+bwgbTwnCr+tUZDLgh5X9HGP1rvVn1YeNIC+nWhxb2xVFfMKdoSMmUjE
RIatyAPQhj0PYzMbSEF/pyHf3C9zBMIZb/diuxeVspcWoIi3zoLIFkAXQVglzl+o
6KP6QAxzM7iuv99tliubO6rTHfL3v1WOdNUgKmyEv/zbRMcOro5PD1ODCh3emj01
FXPVOO+0XnUbNx9YLLHgLmBqxULsQ6HHrCrBNqy9ipI/n4RaKML4CxxiAeBbpSfa
X31c11rW1CXHuf1BUISj+DEwtwnEWrhezuJ8IKUur50RM6jYq7P7dRgEeFHbV14F
9MJNJ0T9YsfKnqhrtsHoEgMeE6P7vBcoMnqKZJgZ6w/Jc40hjtwELb6j+KS60t2z
BchlzSGD/xBu0nHP6s3AR4OsMr76I0MLJMaVU2odNqGHKlMZsbo50gmDXxg1ufzG
i/QpKyfiI4WZjasiIbc3EYwROcn0k68OBcusuLGdMUc6UpV7bGjURC4WfcQD7MF7
uwJBz13hW/KXlZICoHP0RjVdr/SO8h4U4u5D1oACaddQ1MprWlKXKMpEXLo+RDBr
k2z9tF/NmBS4BvKJgUPvO7j1uqzwsciFkjSCMB31YOV+qG94f6fe+o75WK4IvKYk
LYAmOvaip3xonZIBxqCXyeP9AdgSNU9MqaPm84AtuELbS4fMpbTtpEd1XpXkNa6Z
2HaxBAML1HP63CuRkiW6EDS0YybNvh5cPZ8HQK/Gk4CTEJxKZgR74XfCWZNeSk0w
cjTjaqGLYI43XSU7aHN8ntRh4tHY1Gr2fe4a0LEy3Ez+51LA+Zm0/M++S9hvtunV
KB3tAtJUAMZLNcF+5vwle5ShXX7zxR5F4Qr4ow39kXoTzr1m98rQ4AylGU8yGKj7
t8Tidyauqrcq0P/WqrT+YrKV0yRajwsTNKFG07ealxHI7ib31rcNs9m17GmcCUkb
3HbzxR5iGInCFT9cTcVKfV4CROfX+T7LLlZZnFCDYQPZE92OKHPL1z4RTjX0okkA
IJV0tqzpQKjl2mvctc7GMft30J9pqcdKV541Xt756p/Sh5Ro+hO6toC4agP9Lonv
767lx1pkOPMPFCzq9FhmO0+uO1TKUqMNmakRpYCzvNfc1NMo7imWpzJdqJvgG4to
Iws/f2EVRiuC9MhlnDVaBvOaZZwFCYQWEtyUzpLYMPmHHfHFasHfmF8CSnGVHmCp
5LQEkErQk6UM/ji7sm667iZ+cWEmMWcqYy8e7WzadKr2EO1pabmecf40O/YFqk0y
3GF90uBbxxCV+ltbZ96nZnClIgn55lIo/xdm0kqsUIJbl/WfnGBxC9eb5v5n5E3d
Gt5Rxicaqgr2GKk/cnLpMN8h4wG+gticJX6z+08bY5Ct2398nxmHaJm6XrZZjEsR
dJqL0056jIb6Jia2Lk1wGtsr8hM+77RF71MPB2p6uQw1ciAoUakk9buAi+sgQiL7
9mzI2fKbD31QheZilPmv9AS4i8rFBBfNczKRUtiKTda3/2/bY99jw8RHTJfzI/V8
MSg3K/hvrx0c0nN0NA3DEwtnV37gyCVD05yw88j9SrOwSHo/si9alUP+Rl8HUOrB
QpJizvMsciDT7O2MZvuED0UahbEhcIXpIslEvYw/a0YjvC3dCsb+9FrT08H6isfY
+uCzSgbR885HLjU9h80+2mXywFGLadRXdjPSsEmf0uPneBHMu+qkvuRO2XoYsDT/
2+Q3xWHwacOg9/kgMqTVDRmqE+QKXQ0mpeVAh3tRGT02q2upZy90J72t3jzu2O1I
4pVNzzQ2z7Y+NXlCq5Y1Oc93Pyocd4qCfp/TEA7ZFwkDnd4uHEQbWgEBqmXhwP97
kmQVhD614DqCeBKOkGCczTyeOvmrsKHERZqt78PXyeoOat8zgeMOUkTo9MM7tMcY
WTWhF3QV7dDjSltFXKUmpUT9pyCqNQfdpuP1QzXAitXiFMQq/TeR8kFx92O2DtCN
J8hezrYIRd14trRBB+BNuWVSgwc5zEQAk7rx9eTxN6b03cu8Nr0XpiLfGV3V3GvM
Gnm6kVAgeXVgiP7baO8c/E4ZYoNckR628nzCty4xeiBdI0XpyEZHq+WHbTOrI04k
BJ7Hbl19rWVNZL+UTAZvxl66ZaesOeAUGvJRsx0QAAjfC0TOIT2H6NwN7/o1nT3o
1PzdJuaZ4YWNK6knOOnLR1EcOXPG9rdxeKewq7GE5BicecCbNPr6RiltD9dzwZ4h
SZuJJVASBJLbjg0SW7hE9AcQ3I1QgP1GLRa3Lt2jv+zalxHwi6zd2PHNwlUkZd/A
fkNKzo5QLSg0qXwTIZM8nlnPP2AM91s7elDWHD02Kr4B7n23LRW5Vn3cPb0dQWwT
sqX9xfw99IqnaKX5iCE6+bLjfY6biNlhQQv4gFt54ByB/EoMhup/G+4pFfTpzpxJ
+VMOWa/rDQ/EKQiA3hBwY4yktNQ7HBM8wqxaPa81zPE9/MJt8mBrQGHJ6+7xUDEz
4Zf/05r8r6d/hz4nJhu9oVqhcakFuyfMG6R1mmudlETr5pF6mVgXXCmPjXnJrH+W
dTOzZSVfs1cTzbqFn9m3a4XAMadV4GSOKD/EfZhg8+PgN7wMLyzq47Vq94Llv7QZ
jjg99B2DAjdksLel6C18g+p5TjQuDu71On2AxpiZ+ehyZkAgSazZ9kxe6GenghY/
iwmkwk1HCcxtVmBaWJ5XD0LIDwR9tZA1DXGxqxWPDD6o3VttmlDYrOXQPiALo3iY
4Nv2PIsFqU0Lk7mDB6VgcmGDK/o9Y2cihx+w3PE09JA3RJZYn3KEO7FiEGyJUAYC
EiQ/glKbL/Cmj6NVJUCTADwZmp78a/IHwCm1Z3UP8aWr+5PhVu0zfGlyR0xDdA0c
BZ5H2VmW11EZqdpFQOp+sDUCQ0Q1SmypzUhaSMae/wQKDDvr1dgjFl2UmGP68dKn
+JRKGVBOjwhvGZkRhpeFBzg4AIsg+xPTaC6Y2n+YVJ388yQhVElzmnxCf222Y1JU
68I4uL4RFuIsQNJH+s+OKmXfwUeYOjCltjpPnpSBTEJal4XW8YWLWfuLfZAc/nm3
8juXC3kgwjzITY4DPCKvWE8zWO0ESgugOI1ONLbRV9EDZyTjtIqWQwCcgAYa3Ica
4VtXuoatf1zYxN+V2TUvE5OdOcrWeIG+eBuIkYZ9bLWX5B5j0KYTKI6yCoZgpv0M
5lbDjGSS3L50jbaM/ZVHAJCao0bBvK0ldwcHRtAizg/Xv23W+BbJtJ+cXaBOEmzx
dAp++yOzXhEOxZkYZUJlk2szLOzrxeC3azYBDJL8R7b646V1146mykwnUcEdRMKG
1+WOPSCRYT73xNAyyLCIZBcKo0SNWHeoMrxIyA94X+mKEgpTdaUXsFoMUNN2ZpVH
TqhScgPILIq8cXh8mZFGF/8bk9K/EOwgFxwDnlvUQXor1ZLJnWfX/VIadLwQ4ViP
u2ifxalGDSp6fs4rNH2Zr2lhjxpjDCiMp4R4w1BUyUk1QkQTAQbStiufQ4Df3WqN
tjaGOe/SVaYzYUrNQM6KpNI9j1AKt8gnOBVcvP3HSaWjYB7srVdgrIvOrlR4j9eq
zE4Q/ajBKdP6FZzG5rGwFHj8FIqjmbdZmQB5SimKIukHeB+r77QGERbrRcymGGPd
DKUknsG1NA47bWd8CG1euS8TOQ3Nn9oV/NS4sLRBTpzpXHJu/q+RL8aB/3mT6OGP
hvNEUljBF6KzVI6zy2tJMSsW2Ag+K8UBbypeDa/JrG/omYha7M14qLfUfBJ6k7QH
pAWkXxQDYWjBxktfuL3TeIkUZoICaaeZddb3rlk0nDj7OnCOeQ66vrRKEoChMPXm
PDNz7xvdI9l2OG/wfgmB+SvaifVcZhxCU68Xe+JxUQ0P1ZTU79ixAAnU4lS1O703
zp/Bbp2YJcs2kujyDvebUw8OrI+2dAz7lx9aU9XK9K8GOe4IjWv3fus9t27yiG3g
1n1sjaLRvTyZ9I1M7kiEi/LQ08D+JKylDeMpXWZrLqUUPfb6bL2iRRFJa2cqzTXo
YAoRsUyVqjPzEXxvmYfEEJbTMocT6dWDurs1B4wVQ+l7SYpK9B8yXxsINi+s91Z6
vWxtP0Fs6OTzkEuaI7+mL7UMpfBFuialt5QFxTccl/jozWcUVnkEEhcJEEZU+6vK
AIGFC4pWIB74A8UnBU9N/Hp95UtMJAniy2oHC9oYLmfUMcLlP6/8VeRNOrgAB+8m
wvmSBj6s8lusXJr1wi5p1wztkOEbq3/jO1kgWJHkTgvEdpkG8Y7TlDnpUhKzo9F9
GFqufcnPigogcIBLcOV6FAXPFeZih/VxT9Ut5m061xNAc29Pe4vHRuYSzsR9xwXu
wDTUTkIdkHvHbNV1yqyaLyx5XAXqAz9LcnLry4unLsmc9vcqWwyviaWh4NsvxMm0
3r5nVsxQ/0V0FtRi+r5qyvElLZFOnYemvIW3R+/hr6/4YF2yxOo6wFJHrezYvZVV
b8+ptJdGu4inLsGx4WSUhbYxqed+unh7fWoyWQqu56M/T8ymtWAc06OKzSGs1ne2
aWfGqm2VgV9B5vA46V1/G3M60oaTpqXQpaqJRmWvgPCAEJvFXxQvOtP7j88eG3p+
xVglV8lDSdpNlXX0kKz2Gw/P82nOUxSX8TUvQ+tMIHBW0Ukixdmmz+XWI89pknM1
PbmP3NxBJZoBRUDNGweN31iZ3s6rPe3tr4b1hqJ/yh84GSfU+R+16Y3BVgTi18lP
JViwYrue8k/TKskNcW6r4HUxmr2+4LP4RMweKYmXBnVzb9dbFLxksNTO64hOoIGu
XlI57layb0SUYgxdOm2Yj6F+OtYrEq7/uQlu8Wj4U+o7aCx4YgjEEKRE6Dv7bI0N
MdaUSFsxQ4RnEPvNljQPLb44qRs0+a+4sQsY7zgZpl/J7mmJjOSGJyT29dT43JGR
92zbFMtHXiX6L3QxwLDomg86luHgfDCqnY5CPJYHWIYQesf/16w/CZzz6owKqH6m
5Op6dlBCbzFbR4unt0EI8XXnUi9ql8825pRqvIUUiRLnoVaZ40VpE4fWf8pCQw6A
L7Fw8+ZmnXnTeqI/zpqaCnZ/rUiSDApXkR/rhLPAIFBgYeBMWotD/sGc3OcG467r
M4oQqntXuIejDbai9hzwkDHNMouWnXUdUVlDgWZows2VtAl+XA7Kkh+lU2esQE3h
Vq1XYYP2QKGwTbK6FV1ApJyUYm3g+v4RJDsBhH7nh8oRHGJ7k/ZJy17XZmKa4t9v
bH2pctvt5gTRyx5SHDmJHCttrJXyK0dxcMKVAjYRuDQchV04MbLUpzqzdQB2/HFD
CW8rCSTQppzhBzjc6epD/SA0cE4T+6tyQcQI5Sb0kpXuqRZjxGvAH7kAGQCiH77c
VPjmaO2a2B7VvRnpEsilZeG14NhJlOD6EdoBNkpueE9VlQM4UICju4L1wuFOOGrO
09/AlMmQfPoBFOD9YDRQ4USoX0AwxGJshuBlSjDZpyrvsfS3J734egPdyQ+rqbU8
W13Su5DbJsD5tntB0nv11x5pgn7CiBJOb/UYGph4xJK7FlAColjw+IPRCnk3d9jj
I+5Yzf6cRyr+z0pSkL8Amgx10hdyI6ghbku97HvkQdd6SyYPFIFCylRdA5c2O2A/
0HZ0S5tvodp/2n2k/DS1YocylPqdioVjyo2h52g+PkPQzwxAYz+G1EtcJLyl88uK
JhPzQMsh2FBFxOOmKUUXutadbtvas5vbsWZrk8MlKXvkBYSn/bos0jDg+LlAzhpZ
GHzf/wYnWf18RgEap4QNn6X+SylgLJlbJk7x3JDzuPkwqqV8GkT6meAoC3tRWtEE
JE6Nuq8//1wF0HBXo6bNcfPMnx6AgM0kV6CMgZdqgiVjOTJDUGpt4Ffywx53g1sP
MtUT0h2BxG/dOaUFFX0t0yCR0F99LfwypI2qyonFG0nADxiF1j9oGFgZ/5ewpw2V
HhFTaU28iTB2cCxQL1oKxevhADDVl7gz3L/ZkoHz4YLS26dDTC8pEmLHXD7cVjnf
Bq76ErFR6eMGZ87faPYiq3FsDSJeuV9s5b8sRnHGPuG6xWmHr/aDQdcAIkNlBCcf
iQMuDKvuKNYspM9ORcCM33kOPvmKJN0Uyazrnu/zc3/nSYK38hzAxixtomHyBApj
h4G87NKyTjIltTSgawkqJDzCdeJj5xXfEO5KRF7xlOWRZTItuNaczhU/FPm8YYci
UWxTSYlVQIAQItGIcQTm4Wzdls0wIl6VnZAOnxkbTRr3n8jmHCPUzOuiQqeKOa7C
+dtDTxwrV0tg4uiyV2w9LquGSaLT5A/Jn5+vVesb13sqOowJd+xzcyeVtOj0FsdI
yoQZ35Y7hMRBQ7RWbRqgLBlJo1chuoSeTSsXvI+MIwecUnMre96hADoFG7QGRP8o
/s2Ur5OBLBHejxDk8Udwf2zLIjLDBRXkqJpvEx7gg1gnvfNtWQ9pLn7AiipHiRea
Z3LxRwr4nSK9v/EOVBF2E8/2yAblm58Fx91xRdUi05LMNy7ipcQEUq3IC2mRD97C
KMMg2V+UQm3pdc5s3o8NwPU3XsrvRbvFuOYdCVXnve87lzpODi91NZ9uSv6TTGcZ
dgpzvaOmF+1cP2GHhipdYBP6DWR+EqmwM0KNXiViCs7nR9exZ3FRdDMO+u1C3S+8
e6W8Blpq5/fL/MZ52nEu/2Z4VrEw9Eny9XM1hBO06FIK6yLmDAlE1xI5FvEb80vx
UPDH4HTwILAcXXxOP2oVJp+tvNAj3L0znwSDjJuXh4j1htgfDTvB+j20tA4P6eAF
Y4LBenuJigaHYoKENxTHBI0zQiBcK13rFdgAlsXXWnEaJMGQ2aBJ+1bm8ZVfgD99
IckLPlZ1fVBdyxEIhESjoDuU/f+IF+G3ufRpiWqeBOyAS23zFzkjbNMZkVicyxvV
aHXw2jtayBpEmi1ctP1m7Ymy3n58XADS4PV1J4LReuiUQ1z4afFG8RZrVgEx2+ga
MTLbwfkRvtbq9YAZYW8QanQv4j+h80b9f/lmlKHO0Fb6aOIjAGhCBuQVBtm7cVtm
onO9HPw2m+kXRx4bTT66eDNSB3AdkBr9+Shdu8+mH86wEyxL1hvmKGGktU3uUC/q
/3Xx5VUJ8Ou25cvJp1an2pEztUBjVvkqn6vwFXp8cxWL1VDoRODa4ahfuwJCbKwW
o9ZRZWLLuanzTJuDnR1PSClzZqUpczkCDBB40YEOAxcObQWK7Gxa3/NbLigoP/hZ
TDLBOR2GfU469v+8VPfiI1KrFzJTeO3rLUyheUj1I/hEPZZ5YsytcD52OSvaAZEg
oZaT6W9MMNd2kHmtC5HnklD4S3Y/OJbaIsf9VHuFuxjc0lPWUY+x4OWgxqeTGKsf
sIMB9G5KsN0LQhf393V8NywZxr9/dUvrZIKqYhN6/dQrWrPs9xQJaM/KEavqDfua
JT+iHjOz0hqnSxnVPmfUkPd6DYdPxuBDJ34T2yQd0YHx8VVFQoK6ozpnIllzAZCW
f0vwP75JkRwLbyJ4aKUnm7ZtTW+G6CAzx4LKgPGPo/AFlMtz4QbCyZslKFjRXbZI
GJX3cRc+7+vxRREwZMorXdJaZ9u3xl5HMp8pqV7XYmosUO0lHjK3Jm7z0+SEShXS
pJg83DdxUx2JvbqUNqwMrZdUW0vcaErLb1wgPRCd2ONdIbBx8xTl/vIM/HRlMEiB
AotNPQEX/mlfKlgMaA4k23R3HQAckpDTzZOn4EYph14MJoOtDdmuiL2sNrs7+QHb
UdpMNhc01WIYHEaGlu6yVn7XJNPcvLeHgoKqpsGs3cNsn6Bh/USziP+30c/7RhRR
3e9R4mo2vw4TVOTOga4HNceCMJb8uzMImTovmUYjMlxSq0RehsjYho+ble8NhugF
vABxrgS/efUv9VxjCNlN7b/Y/uH+2w809sV3tVqToyr7yd3j3GK/4NaxgY0/wGdq
FDN5tNQPSEjhulg1QeHVSkGvaCjHWnrsmRG1CYco4tEdL1JmNHLBiDyChHVhAM+R
LhYZdrQx2dv0lHpEADZ76vMyVuJ7U4zl6Au+gJham2Wv2NFmPCtRNCQvuGujRwBi
EciH6ZsZ8npNtFYRgiUWcX2sigHLjyLLaHpGC5+f/mUS4m9LvyLX2hRnt/IPMx6D
/5g1Y8ZfLcL4WbWn855RhRe22TioTOLznIMtR5ipstpn+Imeb5oIpUGko+kybAc9
/qZj07lsdCVOzxQAH0GlSoVaPCXgPt14O1voPkeUIW6r0CsNiIJhopvlJVYU2UYQ
CAjvS0ObXzNKz75QlhXRhY5zel1Ln7xm+2uX+thT+KmxRyULhdaMY5ZC7ff16UBL
W/P8g+NQcvRNZPdTqp+C4dJe1dP2aDN7QdOEGsIDOtrZCpcxuvyNImeh0aLVi1l8
p3YHXj69SKokzetfyBouZxkT6Y/9IL3nEJriK4UdskMJMZ8EmQPEKlROQ/FbNEbq
fQ8PY9kDephh7B0iLUrhl/2MpdA+WwOoYzFJiW9sWRLM2v17uEP0LWkYFB2P+QA8
ViOO6FiiU9a+EFT0DKQv152qsQhqUk9lcRBc89YMOYLS+wwssUd00/92qRwR9Txn
OEStNFudGizxatbtoV5VfDsvz2JEtBLnKiPJkW5lk0iG4uNQ/xF+0U9MDptRFBtd
9uTLA7+Sx7KpodqQEXKmUIhAQ75Tmyd2nQiPpJJ/F1h06aPUEfBRObyTFXpqk+zW
Vyq2bdCsJVd31Mr/WqGEERjCIA6yIL3d395FZRpr7i5haYYjw3QlsfEcEqC+8qGI
iKcmac7MfyqxFoLfCpcg62chOzmrSMLVVONuPHSVDaBsLWcJNU7ve3WH1qGPBPNx
hjpi6OUlNLyChOsxrsIq1NzdmZPchMRmvXD0yWOOhEvfV2BXol/Tr6vivYbZMfwm
2u360DNZOHvpKQeKBdNBX9TfsKf2QrXJ8k5kUEOGv2Lu01+nN9bOAl1j/mLmC50V
DtQ175Nyy2miESj7VBfwNmDjClTRD++QTXs/nqy6md4sdFO+2ey1/rXsa3/8q085
M81MNKLKx8ndg9TUy/szG0fBL5gS704X08dz0Q2G16NVwvFlc7FYFAnq+vqIVND1
c6bnFMDZkYkhZ80IwZp6O9dQCIqYRpdOXHhzWJvggZtb4WwKfEd6V8L7J+BfbLHH
DDreDLoHMcEx52Yd5XpBYHxjQa2vxbdtUwsCn3BWAZx2XleUeGHSJNX+ERv0wdA5
48KUiooaGGTvhFHAs9+lfFfok3yT5DMk+sscgoNujwByrkXD1oNRkV6olZgZs58H
kh/wSy29V8i97kXY1KyJJ+B9/7G6MLP9B0SbSMJBCjdzbCs5Ys+pDB+fHxuxeJSN
TNVqVt3GSr0t8vVSBkf/owJg56WPjOk3kg9QxJIl5gjjgn+cB4wDOZIVN7+5sU47
EriHtTbb3FDMlvQBveP6l53GSvruItWkdLJVE1ExIQ8ku8pDqpqB+yv47hO0oQk3
zCVWn/K8FE4NJXq0FFu8P09F4nIjVs1949dtprsSarxjShjECdyVFC6Fq5qiO+Le
4TuX7bHuOBw9nOnYX6MXKH3BwUcXGwVIAvobRj/jtRjpod6aE4Uxv1MYbgTjyrET
ww3qeT3Tv1ItqxRL/hYojLg5ZQJ5YJYg7H4OfyA6SI2cfRCsixFVltNeKCO1mw/1
j8tgVDMHjzVUe1QWenbDdyxYoqaycdgYrpcb6f1/d8UkwiRr7r8w7riNieF1EfC2
QHE47tpe0l13gN0X2rxG5yzTKU+oIrW7fiZ7kk94ItSJuNjcozluR2hdFcNr5EFh
JYQv5v1Wd9WQFWxEjmzk5s+xvJEjhwtksdg7yO4kLQWDU8NoGrkDlZWCPgE6N1FR
lck9eJPzYMz8aGvDaMRLiGsnvrcI8EMRc9Czzkelf2JI5DUFKyL2hRWo/uRFzUH9
TXwDeLckhm4xp+L7rcGI3JPFd651ir7VfTfWSRr0S+3pNQxAZv2QPkw1bmkwBhws
bK1Cn7vJ0UW3nt2h80HK3jBw11Eave4qRzSL0fdG3tQLhbN8u9BdZG3SyLJrcQvO
DgMgorzR0qX6v8bNCB/ZHrlm3crRJgga/QGefkR2+zjwicR/LD7xCedjvH+DfMbS
ILqJaYKX+MXlLVJ2/5dCs361Qh+XnHgI2IgAhF3r7xQLfunIYqOOBeO+y8X8ZxLF
yHlw18V4a8SdGNknFFbEuK/YAAMKVF54dhetKG6Iv272eaWQvnY1bnpxabmJu6Ci
ks2pWHe2rqVfizq3N5hS5/Xs2jdbjcvPKhbmbXaJn4GdchMi87urnF2ws1cto3Ju
fyZK4wCX+Vf4sZrApV/+JnUwTKT7aBkTeXQ4oyvhDHYM1wUi9cRSU+nF39vTd7OX
saIJJLfeh/yr3PYK5dbTlU+tSHBXR7mLzU3pOhH7mHOafpDXG0GYVqpmkJrRxrxW
HsaV9GAC2x7vE4p2qVXPjWdZoN48Cn/b1IkKNevbk5qBIU2b8MHH3PuvhOXsIwak
RXOOZ6vtgXV05tISwPYnFdglH6yGbXcoGBGKEjJy/0FhnzOes6FPFrZ9XC+s++L9
owBF9lvggKuYxnSTxIQrs/ThA3J1Tlcuo6Jg3g9MaQRwjnvhxOqAHU+p5QLMy5K+
pZ3rewr/nS4ROOHpDWywO+NgG45JOW6rZr96If1q2Tu5/VKlcNUhoE8TMnPzJN9W
LChnxrPbgxPT914Me5VZEXaznGc47lekvV9ZFM1LBYlhoJ97fW/0fNOw7aLiAUWC
vj2BV77ubIc0IFkz8cHQoQ8El5+GfeRHS3P1yBCzeTVE/VnGEn2QLwObU7g7C8Lb
r6qxRrodpNJoI8Hvzv8/suRYDa76CF1w2g8ft3TvQc68N1fk0y0JUTuWVfsvcH33
Ucsp/z66Hej1IlRyL9COKmFN9PAbQ1NzrePpmm7gOCfEj5oFAuLEv3i6vbFIwnJ/
vq7taZJd7qObBPJEG6+naPQnlAutIp30kTctvcFqKw2pQkZbtmTKwBrUQDDxZIJa
V1P0LmfgWZMF66YxyjlD0SLgH9+K2zrtqfpe+TPkNqyp3POr1HRdyMmA+EnnAFeH
x4UtMH6/clbZRpgqFWQrdfm0GtEVg2KyixZNE+sx4x8Shh9NaY7g9vMDQm0I7PKi
xMMshItJVAAPk3ZnAg571iO/MU14qfEtwM6Ln77kxt7kZsT+GROawwYZSgp/9nML
nNwhmxWpdkKBaYsG9mf7HaTwO56pUtZx78LD1GVMVqryIPNhiLpUpu6oIkG6zDHL
6AUCU1CaXloLPiNnPX4Tsf4uni+F7gITUkZGlrjDI9+mullNwqJ7GO34z4adf/2Q
xPOrZ/vqCRUizRuCHojVuh+DRHytMTngh8w4+zKc2E9BibhIOcwDU+1YjZoIVIhK
hBUxLVFGRMPWBm9HhU+l5eXogMchz4iRFJsuxycYbIvn9CBq8+BeDbuBdOnDB8/s
SPwXUrx+sRueNQ/7w6S9rSSIZunDFfibr1n7WvTEnh1Pd45gLHqpW/Maey1XDvIZ
12zuQUEqWNpGhvJaA2683F3+T97SPCwjos6ePtynKvT578DFO/V1i+ASpdwdNouq
OMUZv51s5nXaTQNnDIvJWVOk6l2Buxk2MtfjfP2sd50LwC6kMAtnMbSgVvUd0ipg
OR0gbGhwMh1N+0NkwyqjvLZZauSaEI0Y3uypIvyanuabDWz1Mcf19XJj0Wurdzr7
LXjhwLIaLnLdRU3blnEgd+IP2xaIVqB9FSyTsdVgc1dAEsRWsQXKi+nDkQ1St0ij
9fVZ2OwtR0h1P93eBGXjpIbV38S4U6O2+vNkkSXHTOHG56iU38ctscOu0gvYbR+5
bqARYLyd8aWpi0IVyqsq/2vJhfy0mz4hoGDI2+JtzcqA5wwZZAQyPb6NzlQ9X1ZG
xpNhF7M/FlJqEpK0NOlOJuXaOrCN1NlSkgTYBBtbPvJEZQY72yUPDAmBfK0FYtxz
wZHofkBcjQrjCP8AzRUovjeIuJRvXlXhwT8XXvg5TEaQ8Hin7oISO1W+BA6M5mnP
I3TC37SkJOHgRWSzqmFI9YI7xbvYmNHRn4LdS5NsQ2vb06dK+q/0eQdAK0+P955b
gLN5pkx0AADGoGEslRmjfFf0N92LYDk1ABTqAXJDCpr1xm5yek6ee17827Dmlotn
yagmw8A/X+P/Y7ih3twhuvBktqa4JgdRdg4r8sEONGq5uM4PBC1HrGDgLpSWx8o8
ZQF/dTmguFSMNzP501q1Bnjt5W67B7TVdv8NubLCBfnIaFkigAPAkaq6GuO5rYqD
L+SVA0b+Yjm1hpKAQOGk8Z432aGQxXNFRrWCFHeQD2oGEOPUDlOVfHl+6MISZBXU
iyTm+Jx5IIT0o0EQjdETXi3kQbqVhFhtGhhe6smaLVp0GKkTjIOt9lgTyfM41xSN
chqHXq52eSQLyaMi0Noji1OhSVSLTUkuhT0wGeLDt+vfK0INtLNcuIaet69lAsmL
QWirFO7ECo8LebypfGgEXJE20ROqA0Oy9eYHZsa4no8YxWbeFsdwyNr1Fr7c32gE
+Zs31TrsZWRVmO0URWLpedoAuMg0hRAhDvngI3cHV2YU42jvp6oLIsOIbfQzmZVr
KW3dP99zJwNvtqh6BmgwVubPowM4rsVW+LTls7wKHeb6CcUeWkkqQk+/KsFLV8Mc
KUdRJiB7KPmRe46B7ewI2kfljyyDSjr/bcYuiy/emJxY264eGuMOoudcwjyEQF3l
vn7OTY9WTcAEdBmAZNTBtsdkZ1s+eHxJ6Lmrv4ulGYRSB3PRCRjDutue5asJwpDb
i2rsOpamwnNJ+aEIvzXxZsQkje7JfSWRV+hrmYqSm+JPpHJra0ZoR2s1TlFtkUra
t7hhWeK5KF5Tj4n+clzdmevw+8GUVNGCb4bVdYuy3wQMfshdOtSHipDMROYKcCtA
5aNq5cYgUWXcBpS2FyLDcJsCsHzOX7YTVzEqJR1UZwfk1Nnp+BvLBfzkPPFRcIu+
+rm8QCALwXo2Lq2eu+CrjTcTDhRamZ0d9Po6kVsdX+rJnoY4qK/3QfXs6mUSoJcC
WyvhaR39f7yvzKi9j4hrZSNOryh5Rk64WiUTWpM0FhJXXYqQvBRvVEnwAB5eXYSX
Dr5NjFYkeeUPKALJ+Pv3wtfCSy3vhspvxdcikFbCQv1P8bRA1l/JmS6qziMZ0O6X
861+iF2sUdQsSCCKfxM7VDMW1jQaiqL1C7zWRXERLMPuRyRqMFcEIasDB6ZkXQI1
bIth/gyXHAeyjfKXan7ilfTDWbdSTfNnvg21H0MiGasuZWYBU2rCjPGmRM1XKhBQ
bszYp4ohXnS4MXXQPlUsNwiCSUv8pOrtAzfq7wlp+q8ie8gHGwscVtdxjo+waiTm
uD2SZgBoSSljBcYo/bSLw1oaiPq2Cw/grdCAHk+DE1GwJlm9gwGsbmTc7uqlRv4c
8g8xlpnQeuzDrRciXFDuCO9IXlGDkZ58nxZv8bcgXXuezM3dbee6a7gdmiwvhw1I
i3uBipFWld4Kz0Hcb/uLP7+T61NrI7KGTRXXkrVdN0EyvwbsYXMr66LW2vsalKDY
YR9PDWAxzmjSyPm8ksPzYSr4xWV8gdS7zMbNK0RvWyaVossso4f3tlHobwkLTWLu
zDHUPvW7uCxjN1FzYWo85Xt76RSCWhfyIc96nJV6LblE/Gt/d0Z50tf+yH2miWQs
LxtabaVsZ/FtD+P183ihuYU8JwG1fWWqHSAh3vU9R+R6dUNg1EI5gJw919FOK/EW
+kzmIpB9I3sqp6vtbxl214eICHo7IPRUUo42WiZHA+j9Z3PYr3wZelT3A++sGsn9
xCe8+wMMDrCX8cuni1A9f9wEUZEKENdfqWxn1TyUDpLtW8Yp3EJ9HPn9FiwtEURU
v2KiLopELqeMehRHHhIpR0+8r9yhwwVno5CC6xQM8C4InXAh3XroVPnMyg9WeKpH
voghyexkjfdc2flno6zCwxguQcfPRFY05bsWBA0sCpZiafGFOUCYsFklq7J1oNuU
mQms/KsDHMz/r96vP3v01mvB3bkCtfnOEW+8MSiPZcB+fAZY1HeqHMUKUxriUMlm
iLJThSrsUr6hGu/lkNPh1eW0CLvvj++CmmswRpm3C29RHRsVsSu1wD+mnvZYYmYz
as2SO83PCWATo8Fg3sVcXoRpmBwhikbi9bTnLszqDKmqGYVq9dbKU65ZCwdKLgff
XBdgxzLgGvqBpEuiWxJhaoB/lZHpF9JSTnfcD/LZZcV2w4NVjgs0iN2NSUKJZSe9
lquS7VP2Tj3ioJGK54py273Gz5MvZEMWFJvpISXcb7jWBwlDMH2aV/pPctCvqx1T
XKI7Gndq1w69QfXaS+ySTT4Rw3R3CibMmYPs8ImFDv2WXYwz385WezBIKss9KYBU
bqP+MQaj1NxWkZ4zqdkX1hbR3dILPCAN7aCWI/qq+cYz+gi2VDnOQpEi3ZTDcwFs
cLEsKSg3tZQ0ZDpla//g+xZ1kujjuFv+6wFcz9RnoPgAQWuEBViypHdCZKio/BWU
3mWfA53Enu9nZV975XqiAu2SdPJeKOQO0kfNSyQb9cPUCN4WAoOv0QW5e0S7NZ41
34r3u9mo4dxsS9dVXrKgEMQL/cAi1EM189ctZwucp+mXm6D15lMpqfWatcifstMm
3O0NaxBjx4UKEDdhblJa56YTBJxEpsIf5KDZQ4R+hnE2Bq+7VN8QpmshmlIwLXNC
Py/ZRNY9U645dw/GhWkdPZWpn0t2gnNTZEOTETk77oSE9QW4sVmyoot0vusIHZAp
or94XPcCdArktmvA+6Vw5qWC7OCDSOipjnvTyY9M6ONKwgJ7DXJ45s3jUPK++m33
PDi14UqaNbr/jcAKrgvJ4Trovqs93PyHscDa9eyN9goCpEMlB/aL6sitL/fuYoGf
Fg+QiI5foxBGfSSGPvFV68ru3KaSlwtMOBheKzgRBs2RojHNn/8eu5JLaKVNsnpv
9hGyZTUsRvsmPtqGnPlMsIXujOC8exzwu6obgP3gGW6AhL5ioZEVIJMGRNcCfpJh
aBfUDU1Ckau5ESS5fQRBRBuEZU1ijvM+CSJyWYzrVVoF0b5AkBFEkMGmgvnqs6Op
YZHUka0hSs+pCeGVvsqehhn6ZZTgklUxKuYj6XFHUHcDczxQ4Ks0hAt0BSGVEs/K
pRYmIKvyJ7dtnmXIUBCNWdMyLvO3mJ03hPwP5JZbrDe/Sh9eR6l0nkUwfpeuKcyS
U++MTm0vHRo0FR8qqT41heOjhri+O4Uw34I5kWfjwnfsdlLs41U3UMtgEvRg1WJa
L5kwfriowyFM6A4qbcCbVf3LpJT2SOU+lufMIRYdYRtTWJiln0DBSjGOuIQrggJG
o19kDPCLRMRALvvoUthBVooPjwhFpKlZG27Wx2aZZi8o61fTTl5fQqQ9rsjBa4ji
iRApVqnHrNUDlBykjfAusW9uJ+7w8ATIFYX4OGx3EBq76Rh/1DaDXWFLV4sdxhLC
x8sEO3mL2ozTmz8AYo0lF11mRv0fpIAhbk3Hqqs/mubr+yNOXzGjaT1Vc5Jnn0YE
7Mg6gKl9El96ddb5tPVn7r0SM5UJo7Zuf4ivSaVuQ96ujhZ5iwsJoO3e6Q/yWbAA
haqaCoK254pEDcpP4qEFkXnqxEXMkKmmczWsyYKARD4gWuwuxPg7XlBbN8oBa8Bv
4hNkot3n8msb7IwEvNq+irIDqrxgUb0D2bpxog3SDomv05BiyOxcKMr77J6on0ee
eJiW7IGTe9714/gWxYxVNCDL+Dcuvjx5BNUYVO/d7xGJ10Jtx9ZlqAMbZn7ZpnDr
CwohdJYyGmUy15zaBqN8uLAm6w37rmE6lwS2NTIdvkzHD2b/Bme1Pys5LYxWv9kI
WhZpPI0anuoMb8ndm7AoOU0LCscoLk2/iCeK6KaIGEAz1A3UDx/yE4AobzOEtRzn
3sRROM7PR5LNzQfIFzIPZDSoWOff8d1eT40JFLL9Y2F2mEl2/rrdhQmnM0tiXGak
wfW9uPgh5NOrhfbR0hTsX+tfrMduFlK+WNoFZsPmNyfZl5hIHELHgInjZQl+go1M
8wMBFSaJM06777BcjgowNyMiIMig4OTZelL+cDbJ9AHF+S7+MuJddtMt+hgibvyj
STGsUc7cOg2Ct3sgPvgni/o+2lpllEa14JMtrQTPY/VDqUPQlwyy58HwlQpeD6b0
IaiS12QAfxisEU09B59PrmszNsG+1SuPfBgHzLOm8MlWFfBFGClUHSUmqXdIogjZ
G3CAItqWrC7gNZJKm0azF/bd6h03zHniaiiGRipxrRKQXtNEL1PE7WmDaGqQzv9U
JqFlfqbyc3PjxLV1CGmsRw6FZOF3jsqqYaWzGls/E5JdVj+IKdR7X8IxNbjrt2IX
wb0TgkzlLqoj9t3+FfTsfwl2FM6xjFfLUZKq5qeHRrWAxSmLa+32j5kfwg1J8Ssr
1q6eU/lLzQAlftSdkqczNPgpDaotojPsQsm8wzdHuqIgVQ3mW45z11+vtRQF3mp0
+s0ZgpzpBc9fQSfqgkH0GRc84LzbewprzEyn0BGV/D+Y1gUS6W7svkg8ejHvLUlh
3GPMPKImy0hwbcR/0IjS1RYAIcUqSsLaFS704jmRYkG60/DX3MupxISwFZJJ4TNw
HirNqZS2TiYHICt5hu3GJ4UqNwJJlAW1D4CMBQyc50Cs7uHxviIez9AQdaO/KyNZ
c5l6jaNkU2uVO8/SM34FhjR/8ba/qs5GW2K/56kbUah6cNYuBbP43sTTOYX+3gg6
S0l0SbzooFCETB3J0wfkem3+OlHFh3xk0kNASrTgW7si1pTTc3nmpOdWi0fjfkvG
FXXEzcps/VnDHF0b7cs2KlXB3/XuDxT5SWXJ3UgRmJTxbP5Qgq85NeQn2MBdR/7v
U37SlSSCR0YNS8Czd1yYwNqZOWya93bLOlZBcVVwA6zx/qTdPGbo1qBJ+TBllecU
er5/7S+XBNm1n0q/k4pTkiGkjcbG+xqMzIwiL1V1g2W+B3J3AgUsG4N2qNi1z15l
WROpuZ6tlK1plcXl26uIEDZcWLNDOFqTnBwTZh350cp5Vr658Gg0O2ey5z23gVfY
dqCOBc48PepwGJoCoISkgLxYBEmRLNrElw9UaSHJTBsXxSd0jVo70QmWeCv0zYrT
vYCLAlN8WpWhnc9Q+LSCEHtDVkv6zWka5z3Bmo3RJRGcoFk55kKaE3nYBQWAZiqx
l+ILQnB9OGsapOpmBWgo3lizV31V6N4DC+9NzJO7iMe+U6B+xtcC5UxInpGFBamH
yQA3egGXdrfwHjvg6XEjA8pP9D26vQqCN+a9B8ApTho/O337zgYzTtCX/5b4C2jh
C/SyFc6fyRT2uSDoM6hXx37zuSBSl9MOvcxE8u+SfdXnJ/cgRrIiUj0wCNFEBkuW
whXGvNpMHW+ky4Ohcch7FIWnvoJ5zwTOajY1oLt62zTI8SWmxm9r4ZveeUTRLHkw
zZJDn/BqBzq0vWP24tDXVbYliJN/IiMm/VQIMf5EJ7oN7pOSYWX6PPrfGhX44bBd
LmviOlFexWrX4bCkq6jESNrZ1iT/XRzeI7BXT3iorYjJjQM7BoiWvkm/CEbdPHYs
6AAE9cF3gFj/N+MvUZY6idKzbxoQTzXvwA03ALAJM5ljfMBDTCje4hijkjXyDalb
az9tz6OVXBblfQ3hsYC5CpCMnlJYO/mQuIzM4Xd+M276KH4n1HPnzSihFvCn6xhc
Xe07NCrG1xDJQj/PjdINLB4GFtigZQAWiitbsx5jH9zbIbAfbjHgmRyVE2UVnDBr
ZILrNCBPoH8j+b8KKA6YHHJ95c62MjP+JfkwCy1tzmCVsDv+tCaTkNAw6YY7sF0p
YGHtSQcon2afaM85304CX5dYyr94lQW+lsCZW9cVdWevHCen6OaroXeCWLMGY5gD
6kkkGTaQTOdM8FvG5VDI0z/KXi4387miolLUi99hlvY9BqwoL5oRiGfvUs2VIhv6
cd6+MjIiN6c52TESEiPU2MpfywXp3PaidNTiYp17v7zmGhnACt1uPeKkZVxPmfwG
4yIGUhzGkPy+5xbjwrBWKFW+1SqXmhIzpOXxuZKZOg96UWVMPdH6Xl+CeV9vV0U6
55NYlsXpZJ3GlKlMw7M+AZfiOr1t/wDoNFXQxBt2if17KrGruO9H5I526bRURWvK
UGUVjaheoF/sTT1fTDox7vBLp3PXNZ7/MuC/pgtM4w7To5DvAHtZ9wMIDibTyZMY
O5W2kJtHliQxYY6u7+vQ9yT0zUuy9062Db38+onS5vAtzz6q8yRxLCS6CmXYeqBu
xiSamj0QqUuV2a/AogJEIEc7ryJx6egPcuJxry6l2yzM4s3pn5FnsE4H8SyYGOLv
r2o6KC44fJVKUd2a6UNuMmLMtzv+lL2QwSJcoyLC9YC0SSQOHPU0pupBZLopjDNO
Z+x+babEgjzaBv7S5XAcYNpxqksOJ+eZRAGtmxCCbZbAF6hpTwd46ChUcGez5Vs6
vfuN7zAISNq2XaydZ2zTBhF1Li2L4Jp/xu43fQs5kCpUU2ojJhPOMVv3VrMfHXdA
jVeQgoGmNxFjFWbgU4GXJguxvsloiXFx750gfBNqfYEVL19M0saYMUTd3PizHDzF
ntfhkSLMhCT1azZ8tK2DtM7u59NiFXbVIHNRhuN90jL4QswJK0GkapNddWNW4xWu
xfAezFrZpMfFu2jLPALpESR/uWuZLBW+mnyD8GQ3thR8ORZCq721ucbe107Gzr8W
m91MKNr/Wqw5Oh3ZXb3bFdplNCspA4WqN9Z6D7VU1sclnWlqxXizmiMkHcqi9Gpw
Bhol6TlxQDPwCykRahvJykNEp3wg+xKatxjjBJIrGXn5dtCAFpQewGTPdFS+juDh
DL6q13i/8qxKPplXT3BRg1I2/E/wpQtFuDASco/HlsDVMac8wDZAl3I0axlPt9L4
QkgOtCQxFr/hkyNkk1YqejACnUJizbBPfGk/zioANNO7Lgf4cp8mcUbHcvDpeSX9
1nhcDWc92HnLv09Nt8GuuRERbP8gnTR3CQh9Axwnb5fsSw+jL1aOsck+ADc9yZ2g
IHwIpHCnZ3viTn5Gd4hHT1kz7g3cEb9iel62ScGEgOgCTaeCXRjOpx3pk493g4Gk
FNbjf/nJqbDCZ7bgw31MBEG4xQl641IWqwJf/ysm147334n0aIjZn8xhIWt1yu1R
2KTHnGlsLMt8LFIwoInMezJLAFlvLfbeYA1wb7OyVLRMbMGjBacmo53U3aGRudcm
cuwBIjtpXaCpfgfrnhTOLBvrW00n0F3RkKalgOI9VUAkeF7n/Kb5nwNISTwTxtgs
rFjdekUkUWOglrfs+y14r5YFl76iLsziqG0lrxNzSiZgGn134iLY0xXsEkUUQ3U6
GDb/ZkeRiPm1v/H59C2+eImGws8YoThIynWhcvdOOJlhPSLgYwlWHTTgCELwhF9U
I+xU/LoZKhMHruNDGqX9KYKMIueu2jfn8fEyn5mULCywCQPjjGGhvnu0VzRh3V8U
wivO64pT6n5wEEt9LNUhMbFFXkfBlve253IlqzbrTJMn/ALY2feeCChuev5j+wBG
MecDeQ6TLsCM4+froDmLqKr+1c0wfiIJ+zpWfUfPUJ9a9hd6mAPmjfijOByT9rzh
bAL23vNjUkZfGwg7/RDjhMgQKd3q6WeaqctKtfbRFzb3B6T6xF3lgf1VCr00T964
qaWbUbtI3mc93e+GQ3d5b15OfdGmuPAhNSrt3132C2j1Euh9NNpWECKNpad7Yl/U
CVoKujqQT/5Tc85Lau6jfmwjKbhInIw+ItkrXDC+UgmdAWkI2YQEsJH0wFueh25Q
zByNVfKrAJCG5I6nG8x+IFKc+W7mSq/4jwY8gVcQ+QECVTPbALjBnsh4a3ZS4JNT
NyANPsQR2iHiijy44wl4on5wEMAT/9pgVmbhg7dPU/cOxETTfQUbRSG7rSADnrug
0DsFJ2IYBnqUYcnoiMtjYej2JCdP3W+ePq85xZ81AWM8/OsElTT+YCdKlBk90TNa
aLLI4hLx0fXe+nadLZVYHgdrH/StPWWo4P7cUuRucwFWYfNNoL0XImprWWfd5vGu
Mf1QAqLHIB5IFOKetnzebX/0jVfC4TtO+pYWc0d+Abe7fv5Ss1D2PkRLE98fTTWJ
+fJZeZ/4T/GYQeQQnLsDmUZWlfPcjgO2b8f5+qjmYzEcbQGM9GWv4RKGTsSopXHW
UBI2ThFwwEnZ1LggwFVTshwViVMVFNtqKC8ST+cCd8ILFex1P3z2YirJj3AqVnl6
AjpFdo/xYwFoUryBWfFom+QZPrshHdP2n7wZylZVNhuk+vpU9+1SeYmBBtTe/CTB
xoqq9IkoaQ4IbZRqwVnKNgXVnTIU5E+R9vb2eJwbFB6SN6WH/iU58HsKCqQi1IOw
b9+055XwNyqh1PeQANZ+23A0fL8zVIhxfHVhqmCUray5dr5+rZnFzOsHfEjfsUa2
lKuSxlKPg/DDAs6Tio/X0xdJFEU8mu/O66A8barXQUHoeF1ymz2raL2I9davzVwG
zGVD4VOO7Akrn9KfpFxCR3m78mTCllmItK0H1YNJZD15Qy++slrkWuW17/7dqGCP
lMG6NmhAkSaEfCpWPV0dzyJpezTZb+lSYYjB/PN+RO78ALhaUCPn8+0/fY2MoFM9
gg5vamFBPuDJwV9QrEZm5oati0UqLC6tTrN3Ov5OewcDLyUmcPpfwyKzOy2pI6MA
pOYemMgKftCXVVQKaaeOBMSVwiJCBoFhPJz2NZ4/ZilVpeTuTT87uVYH07YW622v
Gk4A2sFzP0altbQfKxJ4OVOEfv3GvBDjA1ODrnM/MHC3dpJMbhuSQzw8/Z/SvaIb
CBkWMftpEth7FKcAsVD4liJBtZ5xxa0+9xnLiFiZyPSZHHZrDtLesjhTt5d2TY+X
ES+dtoE+UsHvJGCfO9KWNbCrAq7AcBTINfA8yCvVoHPvQpkX7LZx7hM9x0QybBzL
WIO4H6AMOXxgmuqD2ca1o9ybS2OTmEYvyKc0vmG95A3A/pPLR03oCXLarmMxZPI+
BKg3duuQyt1AS4VwNy4aB7RwjjWQn0qRQyPiCQe9cgwLR5/EVQT9PBkr7km6SRwx
PCLZImOluUIWoXTCjrSJvGKQV08qR99QEcCElujnJEt9xFjI0Bcgct35oj9AWmWd
oN17Ji5JTFfcNujPytpiqSD376nsDkcObTk7banYintx1IdND5x0YkACX2rthRTX
g8m9FjiiUE8TVn2/Ut5W0v2O/9b1G4+tSjEu+I4T3wZLCk0UJ5rwbLJahyBHSNhn
Qt+xi5ZyK/XCG2JxD5KxLhTVuok8Z4T1KnNenBzDWT4yOIEZcI1+LNeCfsrNiP92
aJRl0da4tj91s2BhCs0/fHTSVEUL0ZZ1nrr8H/3j5CQ7DKIo/is62gysPH8wMHQF
K9EBPlY5FnZRMmmiEfillS5m7YashCO67XP/pRtGKOwYkKGVwxhc2iSh+6sedWjT
MW5rozeJDtvF5RAo3qCXlvEeTswmbYMGJmg3yCRZRY6SQU/f73T28ZJEjGnXQ6Sn
5G+UZWALzZMLBoUgDapaCDuVPT0esWqsDjUa7Je3Px8KkXDOQU011mWt6ufeiR8f
J5zfUTKTxb9lteaqtZ55tHt7hEsUPXaf7YWl4FABwbk/eLh20Yi7g6zl11VwAwCp
KP9XyZJpswd9bVUFUijeFjI+3pzSjKxSzmuRvDZxg8YDUuc73eNkjNHrY+W3yvoG
a1+VF4gQvMaL8B9IFNayacLvsA3sAIuBnxxyL7ZyMezgpsiKqJqt4Zu3Nfd4p98e
Y/QVI+NedUkttLCQnPtSGl89MZitMyTpxo0q121HMxFz9Re4lTV3htKPeknlny9u
Vo4eiV5B0mMn4z1p7o+4gWJa2sHydbbvBhZC2H0dfEVLjVaGq17o6a7BknkcKWiQ
NNMV14BqU793ysxOYjTzzAbKkU4vCY4K73z/5p9cCzSSyJmMK3mIyrL6VEN/E337
F8sIEH519jL8ecRxkDtotuRFWiuzh7qVtrRv8cBuKQ7EGVbwRFIpFWvy0W8jkVXo
PeygrZYv3m1eL0+880XPvndLQFynfBKtNXXY/7fdZZL1umGGmpUfjol6LjbaTm78
HlG66GAHe5QIHGVjy5kpNOtXV0wTXwO7jLWb2VZRvIQ=
`protect END_PROTECTED
