`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZxBSTjZolYg2v3+eolizCd4rP60b+D96xV31N5ZPwqhmFwb0NydGkcDOZeMJKQQ7
QXQdwH7R6XsBGzpDwIn61/MxvJow7Ih36uwArmEr8g1qNc7csnHvpbjk3KUP9WdX
fVsSiL05VOnhJEBTAUMiAkIe09Y5XErKdJizrct9OVlLnRNURqMUwa0k0FtbMNf3
NXEeDQCHEESN4m32hq//Kq1vO61lbuTRjahY3RrawvUmn/PBm1p9jKT4zijcXYvg
8qaVuERvzVfr/9tNbsYjFa6D7s2qkkSl1KmymyM3RLg3UQ/y8AJk95G2SgQSeiCu
aIJniXVqOA/KoRFnooGk9CmS6MvcBjhxunEEyunakM6Rjw6MU6QRWdUQCKd44yE6
QZ/44Fv56h9QbzQSus+p4aNmZa/ctGhJdFEq0bfeIsYsolYHzO1RHUx8w1eC4s1V
Dm9TPU8q52M9ff5c7UFL3yC2NYdcUiL8nzGB6h9H3/1q6s9yDvU6OV6Bze26ScEu
qr5FOGg/w5cxMfyrP68Iq1KtL/qIQ7kWWw4tKsqvidHzgjwhhTJ9CoJ2H6WF1EzC
tTic4fIGUdTs0syYD2DB75LYMd1CeHvs8udOsKXagQLTrC6DuPNq8UQhN/TeI7b0
fU6PBKG/1nuwSP3dDecTTsSp9PXZig+hjzT8PxdUksMZwhcpQd/xD2oz5otOqpFV
7sPtdiUeSzmeFO1Ozho+GdMKX411GVr+aPQ/k/ipWf0rv1mYdQs5ZCyVSJLsJPjM
5NCixUwjU8lpFeRWqMvTaA==
`protect END_PROTECTED
