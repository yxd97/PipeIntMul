`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vMkNhnRU7SkUon3c9ZNOnlJZBTDbHYwX6UnaXHm+eiyqHVrDGPwTsLgwpk4QOk1x
ORFgmwee7NWm1i+h8+I02nP893BWkzBqEeZX3zdmK1w+T7uhmAO+sliSU9NS9NV0
9+aYkNUUrzmG/wgS+1Z+izmTJS2LXuT9fJ5yTTeLWWb0rqX1LhEcqyzWBZ93eOPV
kjZiR8gjESrh4DIi3gnF0VbD+VeCogc8L4+nhgRAH2VvHON47Q/zuNpn93PhSVyg
x2qeAhjijrQwOfyAh1UXkgZyuotipOf8TdKrWHQBqC1WkYWxXsEEO7/RptSQn0r2
UuDVjKZC66ZmYrcWJrWa2m9XylffyCWixFEckZGqzE4dVxkmJa+4EzbaMXU9jcCA
acbJl76eJjrcvbO8b78Oz6wlUVMzksoVWWfXf27GKsUfPv01VClGH7pjWHc0y4L2
T+ijAjjqRV8B7ZdCno1bES9cEy1W4KhbYg8CLtTEQ0LDOERTDrBwJJKR29pNbAI9
am2atbcXM/8bZvvXdOcye05PzUrJuCRdmbDG4BOTX30xnORYYBd7SSho7MMP1M9p
pUeI/qNZLQeCEkdFFc9Pry9Dc6+nDlFcA3Y19bvAkB2MdCeivSHHhsA7MgARPwpX
JUVQeyoHNXzBb7ELfRgiOrocSWRTssaINJ4dlEiOXf+rzW9hfaz/9R6BuGfno+8P
jwbA/SfdINjYOuEuv6faLLeSSrs/CFUeI9RFn30PSCFuJJyAaImWsZXjCeNjAfJ7
GF7j1AKbO7TFHaFcePQzo1isugUQDXMM9XfS4pL1O8s49EfyVXdTxhkda33XdALy
FP4KfX19WZHpzha95aPAB+NxhAFFNB/LfqWUSahMdeK7UcziZ1eDZxfLwWqZJIX4
BpfLOHfLvfJUS3rP3ozpoDBxVyItej2Wjw9F/oZ7tuQR8YWyu0hjN9bVYEAF9hU3
lUfU/eYi7F1KYKUq4luzM0teSI0ww4GsatZpXQdx7POi0iAw56EGB0DFfUxZijD7
mdZdnc7KJjkpjdWDWH5M049Tt3WY0pT6Gdh0sKpcQNO3oNSaWI4JTMKVl58SC8xs
XBaJqNzuXA24Sik71uTy9aMI2hs3TeUj4M/iVKhM468XAgbM7Bm2NW2E1ACrN22Z
JCZPzxMesDQT57vQwfyVa5DbVsV63lwquYmv5Y9VjWNJRwDMNqGqTPwWXsM0Op17
oLBn7utv3y/o09bO4yvW+6yOUQKXZ6S3wGp4pZsSmD1uJty3ZPFz29GORtY7lnH4
sdVS1mzActGvts4Yyzk/2kdcmjF5qDipjF0dLLQkraWkmceZLpR7ynqctlOFKw7Q
YfPVfpRwyn0IaU6dV7mWQQo/OhvXjkAg7jTxBpVur1xidyiHkwjM1c4NhRUOTLho
HLnEEICwbpr2KjwDBoHxEU2896rCjygFtIxLsrSUF+O9xS0aLm/Srqm5AOeDXWqP
BGWHr+1h3qPlIZBJpSYywr+zB0khaowwlF8U2/C4IME=
`protect END_PROTECTED
