`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWQN4SY6wvOdKhMO1ZSxsQZ2KY10rqdjSA9v96bisfP1Cf430iiHPXlHiEfTDtN6
E7YCjbJowkZIarx9R9DnwkMLnyacmS2idlrAI6igqK68a4WvmdkkO+iXdJWFrvl0
uNdbFCo6F8aAnXeCyCxOU4VzSyGzILuYyTBLiyUiybZBX1HYBx4v+TJiAwscaL7u
nFSOqmKJoN4CkyukPPs+zRksmZYO28lzhinDoEGHYIFti4IjWtWdv2E5Y4o76TmA
LlyEXC6TF43HLsCUqRTcv8x44hffK6vB8s7Tmarbg33fQDs99/AAcw/otuFwf15t
7ZkO1JiRjXlwLGKW+72mDNlKyWym4IXRITy2YLDeZ9tfpPlsekAn9Y46jtBuN59r
`protect END_PROTECTED
