`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOSpBVoDbmao+dowpK1tsXTHTQOuitbNyr9x5hscdLZAxNIHVpTKiJZA2TkXNJrn
RTZwgcEkwo0ClTm6BWI8dxp1e7kghsjKXM10ZiuSlzzWrQPgdHB7WQKUVxxSIXxZ
L3wvd1UVoLvXTNxXn1hX4VX+aEu2fy9lvpWudyBevpzwuS9H79o58ivOiiY9w0yY
tgDrJI7rXhQjj4JlVclHJhJaX2q+ZqEYL0jDmUXLOtqg0NjUdXgn1yaEbFghQ9fN
OfMIE6pjzN3VEBZ6vjNPeie2OxgMiHyzjJ0wz6xP08zSmYzKlqxOBEl6V/XK32nf
zURnmGDE6s/7AjVDPhRAUides1GxEVTjlA+cO8NhAwuVVIUtkRoBSK7Fdy6XYcRo
ABE1r0jtt/n0uQ89R3NWtDdG3/kH0Vt1PvTfqtDrrNhO6Fhpuq45uZdZi/AZMGbI
ZAS05nAD8rfDK9sWTdE9hW4maR4wyGyOq7Ns5tXy4uteznmohdbK3gcLyx5YB45K
98UmI4ISJDnKQ+rnrB3xvqwv2Ylui0LryEpSwDAIubktRLbyP0JIjJQSQWsR4y2H
Kip2NTzbBOgcJF4Qjchipp1579goWGzhBbu5blTPJaHXpVDAtWq/n9faU3QtDnxC
QMpsTziCmnBa4vMuN6td3Tbmun+6no0h5NF9DW9ODawt1vBwMi+6osMZQxLyvTxV
pOmKIAJdT3t+6Rf0SDRh75tbtlfLnGizPxcKJZLfKwE=
`protect END_PROTECTED
