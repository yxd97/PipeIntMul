`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dRkx67DImrujz2HCEEonLkqjWVjvp4hGucgsIFI3crMd7CNdWW3aCNVHa/ntdnqO
kKkyOqAXFagdr0Lq8AVNUYVqf+y49gb+6DQE8U10RswSYJkw8DNFStI8U/MDHDcf
AC5J1bYGVs43Q8mafL/Ca3GGfgTBAWNmS6ZuZ2vYNIsBH5J48gwPSoTYhAkaJz5o
+PISw9G2tYdp76wnc49dxS+GOAVQ+ZCpSbb+2WuKSNyEz2PJwfpySgJffaMbWMXd
a9oV2IryD6af0dMWPvsOttPB5XAWtRhUI11nphZTFJew4IT6fbmMfPGQyef3v5g4
pzwvTtSCjXcrGfra/s38cGDaXLKOrlb3oQAPrhlZZVZXr83nRIcJ24eA69QyaAhT
Nb/Vpo88h7uenpIM3/Riqkv0ul/XPA0Oc6aUFO7bU0Y=
`protect END_PROTECTED
