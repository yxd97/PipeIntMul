`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uaNxg+aW0RoWuhpDBg3jWK7EC2yJjOIXUdnknyNw5ASR2zzeyEAt611yWZ1AATSU
HwXsJIzHsD9yWTjOqveVpSbCZLxqE7PMgxDIWkm5T38JVV4tBFt9BPI8w81jczlq
vIQiw5w+zx3ey95wFkz8dzSHFQ+wRbb9JG7r8kfbISPQPHfAwBaVpDNsPYHB9S05
AkH5sF0QlTofpV4iBd0RvID7dqM82EFhbDAUfC+IwbhX/5lQZpt0u83UgK3q54BE
ccT65d5wZTP1p2GcBrI+PCDNX5i4jT63dEHdOLVZ1uvl+//1Sg1w05z/OjLJ4e/V
NVEMhouqAEXZBkzjZaelQUStYT2tfLw0AMr2ltjBstt+9sJ8SC0x9NkNSu5h4u1e
`protect END_PROTECTED
