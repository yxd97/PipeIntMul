`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xnWLKmsVW3nt85WAliDK2pykZEwZOjJiVI5M9t3eokULvnGzzAXCa9iqyEpFK1bf
lDQdDyTklp+NA8AGmdxmvDAYkQMEVAQAG9zJlq/z9Z9r4svKxoF4nxU0PzoJfs+o
qcHnuo5UJIOkTFnLa4aJPmBDn1ahPaeNK9PyFgMNJCkUNc7k9iZqc1iG654iJHGi
672oOelhqizbYmv24Q52ascNlj2EG1m4DslYLW5yxrzEgYBGjrh9FGrPEviNI8ny
7miNvTquTsm363pdgX48NrcGWh9wvfn8LysQC4X+QuhpPWBdmC6tA0en6h8fmqtp
aCMnhv3LAZaeggBJJeMEIS+6nc6OCcQB1/IN73TvK5DCyARwCiNscnmzDceSgjCC
SSeQJLBUawNfoMo2ACBHoZnsO1rLu+fdq/navEgfhyx4R4qvSXu6HlmAm7bfR1M7
DLjxMTFQx8PRFnZIVHRQPbIyRQlzBPlZymd3fggwg8KAesV2fKMDlQBJNGKbqNQQ
aFrEa52PDrrdgZDBgZTI8D/6OE80IX8DG2LgrG9Kj9tuZ7o2GEOfyTuEfwilj/+Q
gheLht83SwewC7sPfydkJBuDrESavzoKxbwM6oFA3ozWTniOPQXT6bls/WRB9s56
UCH8h/DAL/vh/Kahyzhu/nQAdPYJIEmbPxW0ZgdqVUPsext72RaJ6yxk256PaJQB
89G8kvBQe9+/WLUMp9u6XYBVWoFkBkkuGsIiskRCyFcOuAn6lJrb6+d8/l6lW0Fx
9BTtNViVBUI8robFuKz8Seqs1fCvoVU10xa6ZRAMdt3CBjF8Pps//CkPU/Uf6NMe
nhG3zXq70HX0u3j4/215Wa3f7pQ1Qdavy8mt+2X6+wG1Il5MUd/MK1FrMJwKy8Kf
JQZbb36Rv2uNjXymkOcwbmQ/lj2a+CJwDl3IwnCNxSiGtmWvztQW4xJWVYqQidJw
hBsDcl66awNir7Elh7JutGin48bB0Z6k2CZsZ7I7dFzStCEBO72wPME6EDW/Z43s
xIlT5TcvsFrOGWsM8nn7ZJ/4GCT3zWwdH1R64P+kh0ifweZyluZVCz1qxjSvO5UZ
QwQtL4jo9xcgrJU6GpBoJpwBrS1FaWiQfA33GYO2EcxnzsTwECvMKFAW2PtJm9Ou
tV+D8as6ji27ijsI1Hf73GOkkgsr3jxMWwViYA5bn5in6RYqXsX904fcBD1rfp3M
eukjzlGEFb9PpjEPlg+HMaPpZuEXk0ClQkAF6bUwd5bI/mA30b+Bjfmyhm6iZato
e0mHbXegHrlszQ/arDt8PnjL1LEcX8uxkM2AXCpWipCct8Y/A4ovjIgLizDjAUTr
NjRtbKJImIU5teG710vJhYZVsts8nP9jXxx0yADeFlFq2y74Kj0aSybB6tR+t0uk
qMOpaMh2dDQEqActWSi/qUGusDOnWMWu45GZKsyybCy+E9cd3rT+S+KnwIcU6IsC
Z+vJFtAr9KsVnZwJcNqp6aUDkiFdabDG+/0CPu6UzN/AsEWAzENVdVc2bi32JaeE
v/hGOOCQPXZKudJYrg7hyn8SwV6PLwXOL6hTytqSL//JrpHnwzH2Vab7dD9yl7g1
hCpTcTBFJMFEsTQcizEBUnzk0kAw59NUHHzWhqlcHl6DQPox7NFjJtR5dg29eftA
AM7UHu5mL6T6kW81T8bThegvZb1TXpySihYRhBmf19BZwhS0wpe2AeF3y44ggBEo
XSiOte9u18djRCY+t6lwUQkx5A8ne6Ryt3DcSUhpzgxC0c+aVP6nXlN4rcxDKHI2
MIWKpYKYnEk+kO/1hMjoK1nI2/9dlKn3lnM2gTu8iNsWR04IEgpkzXrpd9/rHhPW
ILcC5HQKTNUPMfZQJre3gmzQJrsa5ot94kkGwH2XgOoS8CtW4d7NUybLIAY4syPq
oAIS82YXzhNHvRB7YAebvi84yYqSF0qT97edIO/bIGTQUWQosbnqMHV1tqnJJ7HI
Sbjb+ScWdAxJ9JOyyujDTcAotqOmtDFzoxj6eu9y73XWEvNXyFDBhA4VdmVqj+Y2
kXsIP1EcfL9Xmg+wZfKVlV9XSFtHMJvpOkxU1zhlYmqhIwbJbIpB7t2KImecVkVn
sgbkw3Sw5WxQ23nD4wrCz72R24Xp++B+G9dZEU8JSP84yGot2UTR08FNo4hNjbrj
x/XXr2CxV8qPAQcsVlDM/Lr1v/MUE4z45QM6VPMXbVn4b/MQxHDPsLDuSO6h/ebv
6kkagDAumqvfCZ3HOVbV0xBemYI1JERPRrIPVEnuFOCcFA9eB6cdOEOdiwLZjY4V
GG+m8cXAUWRSjPYuAVPazzliSxNX8g0r7QixNdLfr2OhQSN952fC2i3qb+sz5n1r
nZH7Rc2Y2UasCjp1751vMU4F1SXAL8C7137Ey9kjEpSaN7iA6u7QN0XZ3Y404kZF
/rixGepnC+rOYDF6fTjPa5nqxMbZZUsiJp+aEvvqcj+fy9arhIEzhfkTFl4GFcOk
wd5js15eMtU30LriRyuYOd70jFNOjy+v5GcNQk16iJhVVNRdFOj/tPbzC2v0pEGx
qrxLl/SE5YaYZgnIn3TUUT0f1OeylDBx1tLFk39tJg/yipr7rb400aGTyTkpGk8A
m9pBTehQcdL8ZsRe7imRAE0Ds7w66yO18KEkgJT7EY4uDaCzlhsusr68AkoML53U
mBoWXOLgGY1aPcAuXmL15kM34ZWeKblaUdfGK9yY/2jzwiuDJuaz4jI0qtTmMSAi
LDzocRJfqQjsLi4Nufar1P1LJit+tHfIluKh9UDf7rQwg5tdxuPAY3qWJ1MEEjIP
RjheL0cwToDpJJ0N1tE8HWv1GJiJVNRnQPpY+AGUWJmH8KMcargkHQbdoWnYlLyO
J0w/sXLxSBDUKalercWBiUNgERpfchgnrs0kPny0orFNsRBaxY8lCGGPnmXVHzTi
trzjYU+uK/+sk60W/8O0hUhHquPHMfL86OW37a9ysoF2O9bc0KonNHEvkGLPfhvC
/xBZCkkvlKDn+28iqGVrpggOQeI4FggsQzK9lqMTbEJ6MrGeVXcTxUy2JJ/d6+Gs
jb3xLepNWDqJJYN5fvQunOwoDlPGH+ylHcX0YPieb5G+oN1/gQkeACiC+55Ui0gp
4SgU6ny3HYToOztDHmT6urTYwjH+JgMhSVlIM16eh5FyMxoYcFcBnkvn8vIZ6Ouw
WR3GlvyO9O/8AnjlhCjR0B7Xf41z34wvpGVwFV2Huamb3I0+1qMZDIfswoSNnAbI
16Ce/F9vuIpvac7CVBIY+bsLMdsbyFEEcTeUak06YD0k/MVBwWIcjnNAM5iijHST
H9r171CI0p5mlI+RMUJyaKru89MpFzkfxbNE32kBanwFRBpaYsb4uiL9KhqaSfqH
eJFZFYaYsBEYu9yaEsNatVLLV2HTzZmqP4HGyu++V4GLMQ0Uq3OQFJJ1IwWii9Gs
onH3BjiV/xzetJkkg1L1iCw714NbJQ78ovTB/rdFSgsUmcLXSxHMea9TpvGgDgLU
nwxeoD5vOFAbwDkJvnfxF0vq8UJ80oHVomhNh+a+ET8gzhpZvcvIifE1zZOE9oqN
FW2DhZV8qBPWHxV+sPXZhrEmbjPH7ITNameZGpAcv4EcpqSJkEb3Zz6wqdLG3+dd
OcjWwPX/Crc56qWg7qHI/vFBKz4EuaOS2Pa3dSjRCGM3t/ACOEJq3SlXflHVCdao
IZjXkfEcQcha9eJbuKRz21BUkNwZenrP0zrnjOcsxH2RUPxBjMwdnST7Xs836hMl
JokDR8reMLzuM8BAlFBk3MBtxwuoxl0Gog9UDsvnjfMUoswrdF1Ui/4rUFIDETe9
49f9XEgimM7/fH0OxSX108XUJZNzFol+zDmSghd2ypgVq/X3vyHRUXBM8Kr1E99/
xdfTAYetS6lTv0QhvAepDCeBY5JA3uWmhY+nXtSDKUA4Ne8opXKOMuX9fDGLOnbl
gsfc5GYNxmJoYu5myB4NyX/f84RK2V5rdD5Xll2FH337gaOlPxM5Us1pd+t8+tCr
9Q7gi6cyIn5eQyQP1tw6RD3YQOn0GRBWSFsxglnguewW9E06oZLrd0GtCEfplnaS
NFOx5mS568o2nvGAc7IVn+GXd0HK5bR4duK4mixTkfU2qFwm+46QfowDIKrHScVE
8HggI6VPDg89RwJwu8iynqs1k+0Eyjm/80ZnDefAVZ957BJyasWANFHG1IP2n7Sj
z65kiAXeuWzks83WMjXo43NHLNqYlLYl0sgSGqwCIBjaZBvVFgMQyUgYBxcOwZYy
Xfm9DlDiuG+2M5KJdDG2emQP1xxSeGnzJxXG/LaQ814ZWbOREO3DEfiz0mio1HAD
4j2AsxCpNNkysr11OHTGWNzMVmwfxlaR5x7VYU5pdqlIJByUtuDBK9bVfkWCcmwN
kENdhBpxXP4vXKh0Zz4tUW0SJDZUt9aokMvR/utweX8q+4uXFKeZKoAZINdepqBv
ML+hEoPK5Ril9WaR4cQ620bBePl9RcvWUBrEWjdHvcrOqC/JPjRr4PPZ4xxUFgAm
hUgKKOg0syGRsIlWPUQN0DhDqzN2YsOX1I7yo+Od7HNS/OnVyM0Frs4pif2HwLUS
39fYuOwwbwIfCe48DK5g7ZjzpsoxS7EKn9NrBMfevMDewQ7g/0tn/7rSRtkgt8b9
HEtOyEU8jT8hx7R9oIUHXG3AmA3urSheNpdpfOefNEmL9s499fUlN+roTPe+By0h
Z/ncZgDgkoMv29WcA7GmER+dO/GnPn/bPgtXsgKtvuzRRjyXDMZL/OsKJdlyJ4ni
eKS62c8NHYv9zryT8h7t7+4bmbc4OgR7RQKSqL22Cs0IyP7bvToxpeo+iIr+55rY
D7uaCoYAl7rbM6KaIut7BR9aqxWRpm43lmkY/2uLPiTHFqa0zMjnElHlaFzlqjY9
N/I7o1qI9YEunhdA2hhkRJtURwNFLyZvVpRTtVTj9j8xvOOqbi/hLNVx/vK1/T7n
EGiRW77C+bfC3VSfHbYC/aBrwsb0BIAKnJEvDEZ565KDQJ6ldLQLSB0lr3Uh+xWB
hJNn+oUUs+6dNXxPmXCFZAmGX2ANVhu2m2abKtkQvzOyguVbnNiwNQDq3zLK2C0s
Ohw8032Z7HPfjqi/fGh5IoNDiio4JAKULEjHVGaoww/t1zQybxVbLr3rvvviFaZw
BL2BkS/B48kZzO6VKr5ilAisZ2ufoSFooRDPLHfpAF1K245PecAcnDWGRq84PSRN
LGn5WRBCoF14aPxd732LZ0jJz4ZjiB5M3fmHQuuMTP1beJOv7gqAgVO8x69LaDwi
GQbDH+hPbuurKBzqB7/otY5zQW2B6Z7XgP2Tf8XN8kBWLX7YXL0csMUBtr4iXWJl
9Fnza9rSODIrovyGCZqzlvT4ldxx7uHN/Sn0IDYHyIlKSX/IaQlPK+YbABg5Oabo
aku/ZDef7j0VJ9/hxZalzWMeATXRDzBgfdtyyvgVaReZ0CZyqyMexV/9tVoIEI5k
oQWWEGNMdkGCfK2mLTk4f5QZWdna9suXtNNb0IHSSXkEqWtJIqqc2thW3UksA0Pp
5/wHP3GNZM0dIRaTdDM1250EGeQXQQU739eCfXneCxjjTN1xS7CZ0S82C0Ryi9j9
a+MnbrhgacqN/3aDWfoXLRtpwuhu7EernlFCyjCpHENgMGGRglN1zi8xbW+6pnbs
WI0Vy0xn9cJXoIfVDglP+sj5CaE6XAP40ckaq10L/RenNUFmn8o3f+6KghBjz+PP
V31JgVqIOQDCZzhztU7QIE+UI5PBnUBVVOwOm5SibP3aE9I+FhAFHq+MBL1t0OOP
egpjgTZ9+mXRXgvL2npFAlbFlFhXmgLvkK2jaqAexFvLbrerZqwph5tx7b4GVzj8
+EaxN9F8gveE3E5rme+swSzKuXhI2v075M/bQCkLAT22rlYcFTSiHhaEmNNv/zCy
Nwj/em+UuWykuOz6V9fkQJpws1M51EWa3JCFBtn+OMdwucZJw5giOZC9koqeZN7v
l1DE/2/JGYyEgGSvbnLMXOjupdUGq4ROugtFnA+TPdm0/OziMdTbRuNu0+J7rx+Q
SdzczdZBE+Ejr8W0xE1HYc7TvrrxruHPxlxKdkJCKtgTKhmPTjqAYUKgC+W7P2jN
i/ZPJuNK1WvjOnnbhvwzgc2ikGiF3Ob9IvW8GB+6xbTVFn5TdTbj4gW0EJoPWnZf
z3F2V4bkXgMIlM260KVCy8pI0+qaKHlK9O1uAP+atR7bixbSxCR0AlUVBCNco4oi
ePa3D4LLatl4AX4Up3uaWJLS3Ad0//cmAGP+XgkkMx2p6Yav7GNfK8qP1+yOaQ2e
tcZERCSpQ5jN+YE6m3cyQKW5JyOVv3RJNrOPEJzQz8+p5ebJzR0PdtOpnHrObo2Z
hiF5Z+oXfqkpQinNWBZL6ZzDtE5w7wtYIZzorax3Iiin90FnRMEBDCphO7eUbRo6
lyZkOOiCpxoqTuAe7JUOqtsKaaRNufb2uDEr/vfIXOGJ/Vlrm9sk0m3KxHf3BW/e
MbbiPVypAglDnOmwt2ybInlA7wspgNSdJfiqnfBbhH0ZJDUzIRDs61ahsprIelex
xCXpejQGba0LxlbbsDS2VgydwuybFKTeV4IdNh4M/rIQWT86mLY+fh9PZY6hGcKC
fEcYJl7SJtPO2zvmNr3nY9Z4Paa2D4mQspY+Uc6zFLVIbU53Cuml6KmwPndOKZtf
OT3KifV87ib4N5CMGHDGlMvbwAtpDXgTzUtYRPNBTei8VB8ivbGfWhNM5ZF4fvoF
kZRAxlj91LqYBeCoKE4CXfDQx5sqY20WRs5Qu9OX3b/V26WE044YUCx0udduQ8Nj
y94x7ClhnhAnFP7C5b/7JZASGKc19qgWAoLdoS5GQpIZ5KELp5JuIuBx0/oSGE+N
wjL8Xb3lF2vhv05vmPrrPmEFZwIuaeTEYhLiKLEwXpD81y8350xpQBvgQ1CAba74
ZaRFZ4ZDxRRckZ49ORRr6awyROA8kGgQ2AMOb3M4L5Nvs1hISWm3rtjPKFIQde8c
Aqtq8CI02m9qtoIxB7wrrXf2xyAASupDd8Bc6LO++wjKOAgaNCHWCuEz4DiatIID
bWAmLSVsLilquEtdN8bak9eKf6rjkMoJwbSBobVh4k39NzVrr5Z9s5H6tsErSuYd
33Diq7X2GEu92lnQ8QWz/us/4nj5fcVmV1ZQzyq0w5a7FOIQDilvCWump9q8Y39o
J+HX5N86ut+Y5/LX2dlrPPs2gqoCHjOCVOsuVr5FGWcWfPN9o45OirJhjKxpSN2N
9VeFLuif09tyUZDCi8VlMDMHNX3StFLvNu8tKvjVin2JwpRfdCg+iiVXuh8g9Qd6
AHgRNHOSCUDqa3BX3JI+0CdMwarFIs58TBxgWEf8nXfapb6kIoUCeECzB6rz3ffh
RB8ytcshgqk6DY3yMPqDxivHkcsSoD0t+5+kI4A5EVIRLOEF8I7jllNinLkI9hWI
sH/Bcw+9LpjBPYevwswd/1N9J7I0sVJd3IeuSNkSqZmft0bQ904xbwTUD8De8jEb
OlRZs0Y0zMmoptMoBgErtLip6H6MWqdqN8stdKYCzOsJhs4/hdqrjTkK23C/qlCB
xJeFx/3sxtS65bal1GG/Q0EEtsatq6YJvaaO260Ouw+UO4mkil6UHWC8M0kxvPFa
Y/nkBDfnJx5zEf+ay67cBN3CIa94HJH+/ZX0i64qbCDLr/RVA/l7kiag6cNO/C3k
jPCmyf1dnIVySc420bQDUdENYtVxre148qg2+kYaqnGp9W4pVEiGycHBkxGvaCg1
F+ussI+t8cBKBdSjhvsvhsii1jtKFm5eqvxFMC3Pmq0UTOTlAWq5mVAR9JGjh6qu
Ch7sYzeW2AY/BdxIlhVOJEjVNCLeZJdhl4K9Pyc2EP/5O+0+/ndbKLA9FpjjCINa
r3pkGBjoYW2rxLPaq835YDwKl/o2tPqleg1962gKtu5h1Enx1sIfg6I86UAWmn2L
QuZazhouHe6SiZ8TJBMdFLbMfFnE1W+OYYx+KIbE7OED7mEu7i874zztpO1ffZmz
lEss4mACxXk2DNJvsKKMf9LYoNsewcYkSTTMfE/54mNuXwx4G8KhncGEea6Pirm6
GYGshWMESmtPIChkI4mX3lsBYbGyRaBueWuMi/5DwA/LVbhrES6CNKBzaeqT1xPf
MZG60nfms3a/jqCxWyfqQpJQAocmfbK4/7pZwYuFwV0+EweChBydoDDJKanLyMg4
4+8NMxkk/Tta7skUBAVQJW8F7MdchR1YpbOb9ruWrRjkenu9q20iro9XlCccQ9lL
ikXu4sOzhY1N120XmpXWlFA9q3gbWX0AASKV/+hHIYGo6o2cX2tEOtqbBnjkICIy
iipSsgKRlk2vuuuVrQJWBewlcd/KvohCInvKBN79J6aoj1WVHuAbzp714SEYSbeK
2TXHE1x3+DUfTyPBlecOCw12qhqV7pCvs9iFDz1oirnp43inTxtGGsAWzqFlwgk8
07Ar2kDv49ZaxDw+pi1HOdYo5h+OMiurksqTp4F3yISKku1QXmHlrp6Jw5zf/Gh/
uU7xjMBCaAm0rpcJecmf1MqUS5FlObqA89HDBv9iOFqs4nvQNBo90Ka3CU6QyCWy
MOgGJJ0dEl0lleqDAuN+eYoCpiarKEPPJKIDGuVuN5vr/DW54CqZ6NjXHNW00HEy
AhhUeszQn3hy6q66YvetyQkn1q9Jn0Y/A0y8trLr5FqwJJTOWi5nN1etXL1Jsmcj
VFvM0zWnY53yz2gCfKNr4xdH7imtMD/tjmQ78qQjkJUi/OuLX/omGHmd+g0jET0O
RtuQ4LutUARH5vevZQy3PPBW4Cy+TpQZegQYrwKWVNIuRui67vc4HXxfB1pTFI87
oCx5ZpiPDgzV9mFyGZcXS409NQJqVsL2sg23Xma1I22yVMNd716u7krHR5G9SDYS
zhvpXQFfaeDyoY4ctRAwyA3puSCrRo4fysHQuo2q2vLnvTAFlWmB8STAcaMOnSwt
9NzT96T6vEopHpnSAVVznuapdOIRHZJzL84BDidNLZXz6yV6+j3tbMeZH4Qg0/rc
1rWEGtmwqHZBQIh60/XAaXm8Oh6k0tw3HW+LIwov3my31Lu5dZsd3/GxCdSxzyJk
04FBhnI7ujD2Ioqd8t+CVQIGZAxBbVW9gT+HV2kcJs4/8bH4x1PWovAMv1tQq4j0
HgxT0OqxvcMrkTgv8QuJP4V5yfenwtUA/lvrjyQ55QY1E8qn9Z7kCTkWdtFapurw
vC0/AEo3w4OHnSUsYNsvGa1ifoiuoCpKVK6Kr4URzmzrR80UZ2jZNxaZ4o6aHaDR
1/BYxwmFCuVcP8OBzYH8FMZEBZB51VY2OTW5E4wdzt1YoYgsYrD1xZyDiI8DiIw+
yY6l+eWIt8T9tUgo0/c3n9oZ17lTgaTuPyA9HrvMudNWPlYlrvPRMu/6Vg46bSPU
0Zq3jOEvlkqIH1hsAOu/hAyjsSnFm5xDFBsM03hnDrtFpHct9CSvo2KfvDjnKKyh
Xyg2EyTeJ1cv3eVTFgs/KJNLygfV1OoVOtr21MRpF9SP1uEZ89JUV+AL2N1ttTp3
pOzteovTTDMR/cmtQsWKsp4BKeTdaxOvX49Sj0kv4jCpiLYZT7hf5L49s+Dq3I9i
XQJMu/ET+BAC7H9HQObDNmNPdDTkJ7OIlijpTG32PbxpWF/HQLnh3FCEi9eDN7RB
2twoyS0nPYZO50Bln46PzMIcHigKTpdOwZUApcCWybcoJMizkz3+Khziu9CTtIPg
uCGXDayrAY8KC3r12/r4VZtwOoYI3QnGfe2k0Pg1MNs5BU4iJ+uSvjcuyaiK17h0
iP63UB7H79tJ/6GpcK2DBKs5kef4O/eEudndhClpgEFwn32PpfYy9G+uNfIf6rC5
9KmeF7gpbw4QwnghVbDMrHYTBv2sAWRZamjF6Rj7ji1uiehl6LxrRZ2shGobbiB1
Utkc/MrD4G1m2+iCClIRRoO/16XJqKkd/WiPhvP51cWCwKy8ETOAKWZ5k49kcK8Q
c4G+F3iXl3yPQ3iNL1zTxfg+2du7KMxc7HYRnT0GByZBA9x5D9d2nw6RTS4WjK25
gdLwWqr0EO8bAdMVlQyDEoPXIt91SeQ5BR2sEIecCUI1HhkjBWe6h6qfvR+dpuJl
DYZB4Hij6NKaDvKYCLO3S+OZii0C2cGjB0RaGSTs6duDoJgdVW+aIg0NryKYQBvL
RAJOUDW1ZS3yP+OZP8jp1UVsTKoBekIT9ieVFBrrEmCAN5jXQOHvk8hnPZC+sZmM
2xGR6iZ2NG1UOAJ2ocHxmx311SqnQLwHGwyZVHpg4rIia3Hb3jedhx22vfX77xYi
Uybfqrax0wcsIPWIM4yx6MvtgVVeR2TOEsORrmOuUY9soPCAMhzqZjsMwg+N0ULa
odkpWRa9J+u772jFHT5WSVuWhH3q/eMRDqduT2GMjRVkZRszGkDYXkJ5mnMwtfr6
YK9cekYhFZ5C4aj3M9wO3fWw8Qwbkg168P84ahg7i0v/s9maHhqWLiv27I1YwgOj
0lmmlgDaQIFD4qb9QluTjoKtbGj4x5yAN8z3W2LbZ7fuQpQtSI7Kn/KRRroDjgW2
k4D4wMx2K2mD+bKjjYM5Q1GqKNiHSyX4QM8QG1WliD14sAbQyohaq/VE2Jmq2VFk
efAxgz4MYzKPKWomCq2I8WK5C2Rfvve6lT3Abt6Kt74P1ws5I4OjY0ZObNpfN8q2
VBePB3U5QImAeYdvCYHAkMNj4fPBmJaBs+hs0fKAoqkMcWcS0cau6cLF4qMpEXRn
ILO0Di8AxcMkRa5Q70D+yZOeO8mMZNoVSLIJxkC34NO8Obq0K/AUzwglbBmM2Qtm
gwxOLipIPNEoV2CPKldbSTdpIZp7+7mQjMf4PT5bpHalPbqENJgVNjObTRZSEnkM
v1kZ0OUNmnL+JIGVQfUMFQLWKfJskCBLRY/ISiTLy5vdZQvPopc/L2ng22ytuLP8
UN1tqzy2fWvSRsvs1zUushrRcEqmIxQBQM067M+fqLz6vol4gpy1A4NTqMMna2vb
AZGi7aTUHkAYozmsb+y7rwpkybx7t74dLouJ9CVzQqW/4z7HVLbRyEA+yPFCz07l
xfho+S2u2lQgQbb6KxTphPplmLOUK4Rza+L2IOOncXSZ8kzM+IjlfuGh2/IzibC+
q45N1UmygEb3vo0Qt13MgMA7R46WDQdxci6AXLZP3Na51cfXIjxwevdDuOsB/coy
0phgTs3tn8aD+KOhoNtRpJzGynJW/WY576cSgvWVzOv+26qDIv9sERsjoXHabYUF
W3L7k4zE4UBhn9x10r7w0Sv8RFILJkfyT6lpw4Q/+DIM5cpRFviE6Q6afgl7rVYt
Hi6baXXZFaEaXC6bSkJNhKHmXRA1JKJuVX/YiogxgVxvQbPOi4Qx9ZCWvTghuZEj
9z+5gZntRRouHOC1hXQIH+bzlasR6Y1VVGLmoxtsaym207LmSSCOWCWasaIcp7p2
UwFtcIhn3vBdmhLxWJd4KUF+5CxHDua2GL5LH/XhMDwXZBDaCXTVKvCmJ9hs5Jg9
es/mucD1N4EiDaJnjUiFxjkxaUcPNamWZ6sJMFx9wshW96AvkTeWX0NRdE/eQ357
245px7NNxLPMf8rUeMKGTmMtU0WPiVzkjWm+0iS8HBVa8usKu0unCNNga9pDxFsA
0mVmfbsMDjBdVn2hHKYnJEFKvYyFqI+mEBhq10+/bMgQWsX0B5g+Q0lE0akn7+aR
RN0qBDUVuNomzt9cZydR2aTldES6yCaRo6PX6KVbz0FWN51IG2uDG0Mg67ddh91g
q27lYHx2XYpZTsQBfyYHgrNByJ6gRndgPgrpUhvCE2Zu+OOSNcKnsTqQ50lV6tRm
1gvmAYD82Bu6NdEl0g++z0J5iryMIhzXIqM514OCgxDx86+AXuQZU9j0WuY98YbO
rRc7K0ttgxz/sp+a/rkqFMP4xNBQw/fQMUi2Ntkr7eYFPioqiuv3UaLSOl3aTvtW
D574aSRV7dMFgIQn+BFU5TwteYF6P2J4iDF8JFjZe39+hH1BWmJ0I/renDyk1flV
fYhen2V+qTb2ku5sxKgJxDhTZu8+UQtHltm/kqc5riPpSnD7+MbPE106C7n/Xl6q
aJ5Zp1maWXkagkbF+CzEYXBF6w3pgWXhEEOCcKCLrJ7MN0odm32fjEZY1PDyskgA
R+CxDDAiGYXcv3voIgzOL/qjjfyFSy9EhieJAFkHPK7oYzHCrKJMzXAK5bc0gJ5h
fYXwPpNgEuwODKQg6iaR2VLwXP2sGV9vHpP8N5cWqdJ9cB8gPmePc0czXGGXAhve
wXTmgd4D3AVyGzmh4HOjmLu9grkDOg4CQ59HgQiq0ftUs05HZkiyf0FhqCGCACiE
zeh+X2BmCBTYcNVqYIAmJPQk30CrnFrSx4KtzZWO14uwEF32gFGrDmxufbyyRnii
b5hfitCdlEdvzczu55Qyij2nStWcGwhLi277Sk54/oNGvkOEmcF0HVL8XzgGGHj2
kmH//eGOvEwfU1e8U4KNHPhaH84QG38syl+G6gMe/oUa1ZTdWGlB+dgb7jhFV7y4
DoqBtZiffjiyDN/9laGwhDIyr5xiVkmTzH9djSMl4QYZkyLLajOZeQ8m1P2M9Et5
irg8UPcaz9HMdppe5bY0Xz9jYKpd9X2e/GaQJPtpPHqgLNKDKnxxR+40TkZGD91f
wuTKO9SiVBqDiyRzWpzMdmT5jP3nMN8tiDeGSmND+x1sUKoA4i6Exbz+XQEOTb0d
EyZUw9s+9pHapkLCfvNsUkW+YqTWnjnEUZ6mJqcW/HHIDpknU4PaNIIUKqGconJd
OGF5BnCa5PFkDEGtgec6nDYCsVa2R8tv1J2IzfKdrQ+ZyYJlztP0rP3Ta349ET6C
0KkDZfn2+3Kyqn5Bhv4FF7iVzVSD4pMQ/xdkgWQBmTODIduczdgaMzoxjJPSeuef
7pU/FsDId6tGLAttftfT0J/x8SA6ssR0XkyDtYh8qmWQIKyjqWIveTs0+oKmyJMX
ZlkP8fUg4JoXLCcrusXCrBNz8OZshomuE84QOJKGjtC6P/y60iw2fCUvWEqhmUMA
xcCQUmu87abVkr3NdpSGCHLZNibZCGS3mdmTBO/koGdlIs/sh/4ECbxSPtfcztra
gZ4oBMcF+lsvQb6bX9cFvF/nczffvRak/IyRPOmEeMRKRnvsh3ZStLsB+j6xldJn
bU7kEYXlkTbQ0a5z+C42YpFV+bpd7jsa+sEsdADikPFdjCjtGqTwWVlVNrCTiF8J
letY0OBXLImEIieh02Olnkl3x79y6UkPJNrelKpOmc4mb5nAG2Eye9j6fmwBIgZ/
rMv1YcYqy3AlKZJESRcH2laemmAljImc44qn6c1PWr7er1skzK/Kjs5HJ8IK6RWJ
RWoZVnBQBK0K8SNLPpnvywR45ytufZZKMLedAQALE7DinArl0ayYy7qRTbGArn/b
md7Zu4bdYAaUE3srDlWICv5D7jEA1nZEepsx7BOOdKxF9CdLUv1i/PPHz70c8you
3bh6sW40+QEjzeG2Lz+5Tuv12wWOkcJfkmkEMXciUgauKGH5dQaefUjt0H6gE4eG
llKCpEvjj/nK47kAPcpXpNjodowfxgCk5d70gYOCbrXV442QFjl6udB4XqqTww0c
H+xVwXO4kDEPQM5d/uk5EjBb6xoamcVboN2DEvIFzxVExWtKEm1AOc2y918xKegx
gYxEiuQRuIjUzfDxPrk4OrBcxXA11hXBjhBs4Hb+p1YVaXwmm+3CHRlS5tAYcWJt
8TFmAm57O3glGUcPcjvuSoSuVhPoLdnw7d8cf/MNapnqzFHeEmMUNMjzgpWL0F+K
rjfldNwtz7B/FxzJmXShqD9Em4K7JnI6lu1c3/7gYc2oQnVyO4Upc6r9zpqVYLIv
dNSKwpLOWxxaJNhHz7YLOUis6MYeJTrvKDpGAs6hOKC3kKUN6sWnGjpoIQclZM6I
UwxoGFYJZ+zqVK8nWfmxrxqDfPvJn+CouGIK8+fl3ulxMciyHu5gXtF6Dvk78Wb0
6wdOrh9ZNRCyy26qY9u/FvZh6PxxZC1kyXZog3CXA2RJUColHT7QMaCR8Ql+X6Ef
0pyzhDJekD4Uo3mPaADYviLOmo3Sub+O7Q0VKLWIgwcy9PkT8yePc0Z3PIrElFnq
RKOUBKAM4nZc5myZJCdRN6qsb2ThI2C/GLutKP9KCrihNxNpNVfv+bfNR9F7ajTr
kOpv7e6tM59qWC77RW0eQuVI2mQJMuusbObIk1aMRTZW15NBdCpftgwQ01ivBoK1
nZaF/YEpvCBRg9ilpSUcm8lG+wgx/VSwYo1NXbBOuZYn7blFsSFM/NMIvbMTkqFn
AuWOkmJ64OiRV993cdpylU6uZk4ZflOEdKhZgLU4e4CDIRj9kD1sC5UzIb6lZwXk
Z/GPmf+2yhkIJXkqh81DjUTG4uy2iQwvVBxytz1tD8cNmGybg49fV8PHWJwLM461
uSa1PTZS/Y2QzEi40MY6oz/xdmRIDlkAMM4urJVceBKXvlvIR2lEDqN1dadv0Hx1
rAlontytKnz4RKmBJVn3aAY5XfaM0p1IUoCRZ3boUIMShbT5V+0BTtHHoidSOOqH
kXe+YUW1PgmatFUxDirdQuNSWdC8D7Aw0UDhwo6f5RLXk7ht24OGbp4Zj4PQ2d+A
ZVBPfW7RK03Ht+yJQMxxGjvSoJQsZOmOhi66xhzhLt0XvAhkwbIaPHEGSOszKJ1d
2V9b6z4XfKkpu4J6QN2USDO3cUhRJrKAxqk1HWakk4VF3HTbEOrO7LpdL8W8oGqK
7fFkGAN/bniVi9P7LDvmBk/Q2hteYlPPhgFRtV6GZ9pDQPB2HY1iGQgoUbnetOVj
UqyJZt/o2JFIAp0xuSSD13l2gCKOEs0xYrg60V2+3qSnphsK9oJDdUM5PY01GSnK
4VsD0DBpepblAaVpDqmw2AMlaWhA2oKveiQk86wikLPBOYFNjV1OGnkZfLnFPBjf
QMz8ZAuGNJtTX2mMGGRd1G5fZYRaL4y1kvSLp4PkhPD0Kol06HZmTek4bOg1pfBC
XAB0ThlqFhTW9HrRdEq74OirzriuA8FnRMqdloDmvggeNjDzVRK2cDHxskQfsm1J
DXcB4aL5HNEEnUcGQICHa7VNUEIpx93SKYMsBg1kDlKmu4/qV+RGWLcIF5QLAtPt
XpQzPcJJMBLBEuiVUPwTX6uS6GMuLUH5rM9gkiKS8wEcTfvN1rt/N5N9GxIqx9IO
2tB8ZrUCejYBHGrwoJv/Z+wYha0chHhpuvbuYc19OzWG41QuHcOU7qPUokvsP85G
6CgR7M1CoyxHIUT6DfP0HPKutxpwj+k5HmaTMTfUcoBGLhu+xNqMEh2zwcwfohRv
XFuPYROxO/Vfbj6vIpxoZtYvrngXPjy937ZeaXtaCZYD82+XuARVrPL6ULaGP56c
W5jYBDsWhkUElUHcupR7OG6OerFVylx4y5zJUa5Jy+eGru3yVEzrpoM8t1wdIvkA
YdSKzQ+xqkBEX/Zwl/CRLxJsiJ8m6BNl7GDt/e/Z5x/XHLsO+HpjiueGUA4KNRmS
zqk2ocpW+iWg78Tr+RCktamP2V4kB5FBPYnD7ab8l3oeIr81/j30LWLv9MYJI2Q4
b7QXKwM76yVL3vCG3sPa+J+Qp5LN6RHCfprz7QR+W/a6RkUqEbG8s759m6grjZo2
5V5gFB60HutFjUYoosP6i3CXtXaJgsBDfOHScrP0Fdv9Ndgjud9SB1EPGDgB2xDC
a2elCW3dP+GFDNahWInFeSUN78FDIclZiu2VkNYciD0RSN4dNB6g59auT7+WoOZn
OwAs1KaXH5PnsLMtyu3uOcXBBEfs0FbLRvGFlcKwSz/xyRw4fYduRlQMIZIpvASx
/4bd57S6U/W3RFJfgC0YacaEyPei2/6AeY8Aj4EaaFLJJ9qrdUkJMlPXINFoGWZn
+XVq2n+FL4+nDl3GQNRCC88V764SemafjI4RcKrtKCXnBJsZNLpRJchRf5NSmmvA
d4SlfUYQEWU7u22+QtYK2PMYItUI1FkzeNZfeaCtprJ19K2akmpsVzkn1x8oJJpA
jfNzcydco5wDJeiv2jnMkVCRzXALfxRrvEkbVNhqBuxBt4/aga6AthYncPpWg9JJ
Db5laUGTnYBR4caVtTBITat7ru0P7E7srP5cNWlijRQ4fBwLXdN2lqnTyh13F0ci
DPBr1pSTT2akixeWx2dX9WTnAnTiQGJO5bdsldMeQ0vbdy0NS+ymwGo+F0feEOk6
sS8wQSMy7MDYCLaEvzckwHDO7CvY3JeiuCZRSqnlureNGSJrF7CATcM4NwN37FlX
Ar3O+y+EH9DjCydjMZnM0Ics4yQFC9xLua7B5xLFK9RI1CCInc+0YAHaV9Q93fyS
caa348P14bNJB9g479IbXwKyY8Pv6Y6xzarBB7c0A//6+x0VBEuq/qjFnPk1OZdN
UAAau8QM2czLGdwP57AsJdV4MRP2aZioonWH6qp6to46cOBKGdxN1wLkKN5JAdpU
5KAB2sPr8dlSXpBQSHayeSVhQPf+Rkza4t971nDxo8IbvHb5LdKiKM+nfRGoYsj7
ud5JyhjhwpKbj3tH2bNjSYqcc20muR5o63wZ4IzYAMit4yBJzVNHhDwiwHUdbZqe
pmEBzJsX0CuouXzM9pEeBsX1fxxPCl0UzxNXZW6XQCr2Xm6Zkvq4Tz8LtYRe0CX3
rLpeBuLX2n/OdkEehDx5IOaXZKBgbFjBouK25gCsoQi0/8Uq5qR3JM9eXgmeo/w/
XBlNTfkPaAERHY8lTMYMP1g3FbX7AdrGc1vs4vSIus0i1O8BvV9LeMR0xp4qRc0F
bHGxWPM1hNz3NX1BmCCZYz6Lknt/3C6sVVVLCX72dZNw4jtWMfTE0bkLtjJpA1Kf
VE/AwdAFOvVBEB8ants5nDUfWogVgtEXkhC436Fs9VTCX4SGM92TYDJ0XqDzFMmD
eJO7jg8ttfNC8KH/xWXLhjGEUTL97P7L1IHShKK4Ny7LqZDNxHa4ivAScdQ9gA9s
ojOZkKXtcGTCvTPxDFcsVgwXL0w8dbrlVKNkjUtg9JLYy+2qwy97LJ4PNahBTf+O
m+6z9GIxFUFMajMBZubzwYf7XLF1fnKqteVHpOMXEVt2igdqlgg4SKmgtRmDxFvi
+3wLwr813b74IXBJK+z8wAmT4fRcD1EjnI8peOfXeQJQDwGuo1FfF8PUBuH3bQbN
+vDNihJmN0RGw0lh05V0ILZkWSGmKukgz4XnUWcbYVLXuYPm3O8vn1aqRiS5iHau
wnRLMVD19hDfRTzZ76lGqQfK2xxh+2UP9u5veNF+8OvqJgx1PeZkEK+PXa1wnN1T
z7+FeJe6dIXtK7ppEkwICjp8G0j5iOXqxupTlg87JkLNf00u9KCZdq3n9KD7w6bX
gHWxPC7HvY6ErBaZuz5h3kPl5P0VTOsnvsBIovfZBPgsnXnBB/jYQrSk3du590dS
Yib8nxO+0IflQxQb3ywlqWymwBrPcGoYL/K3V/LqJB9YJt+53sHGIVQcEe4Vvj0J
eLdsgxF5Gr1Aaq7pzUu8WL/UHbmh7pFZlZBDUyuQYZ6VEtGkqr26YHeVPnSnH6sn
e7NNZcnlMdjjrnQHfJuYGbYyTV6mjsNBd7DiUbL5aXS/eutRQmt2lwtXbFv4We8V
Yuf35xBzZOhW9HpajKYcPE0PdB2C1jC9DYN9slMTtn+L8B6LOXUXah+aA8sGPEuL
ySUo9Bl0fsgQTO5AdWFr8NzHA6HGu1ZR0DwX1fDzJa0BNle5RCBhuQPkz1z6640P
dRtIS0MHf4ZF1cr5Hy8UHUu6BfkE9G881fHKtERmkCwB+g6jzPl7b5Ufr+ym03eK
zKsPa5oxCxCyo3lfWOLP7dCn1XKCOq0YeogrJaDMZt5NJU5ybYZa2/03nC1jWsMq
EzyH0eJbZDuThDhfBh6/BIE6WwfnphG4mSBlNqGEZeAx172RgIFzqXiOBxL8D2c8
9dfD8P/Z4KodSJQyN68155lEeNrkKsVmKLP58WASAt5mzovQ5FJE3QRb6C43n6l5
fVmJD7gfO7eERqWIyP4F5JjyWLJ4v0ktwCKJc2X5c7uWKi8NO8ygT2crlYHYTkHm
6Li0vxlLwCk9y4hhw9g2vgacn6GKpy9LKYl2tARtbDSAX9G35O1c11OiVnDdsBoW
Vx/z7Swj6c0OshLZcdEAUoQ4LevB9aU/WvZJ44dnpg0QA/debVgmKYGlIXZZv+IL
cZKBoSYp4naQi1avPF6Ev4zhwLIRBC+TEeGCw3qM5DPWL//8xpPTXTUKGQpaRVjw
Thsok020XodQhm4hvHPyhdSaWoezVd9NebJTC1giBM56XMmCdlNOsr/uHPEt8YFE
iw7R1v0LAH3UeKP6Ndjn1swZGe7PL2oYlHxcelmiiF+vDG/EFcMXQxQWRPOGtUGG
BGLTuy3NXaBQM45895l1lbA1VZxCAm2NxWF6huyx/b1GY2egdZMcEYrxusmTaFmI
7gZorx08YDAlMDEQ/XWKB/q1C0JEEyiTi/3lqsEIxe2bF9NG6nKgtd69bQ7BRLrH
o69N7/dxia53FqJz8jPi43CDLziSp39Ugg9kAC0QXdq8EKTxUMJlBeAEucCtcR4A
1d0uL1yd8wJjuFAtDgd33P5/EP/iumCB/3W4PYvSefAQIQupn+AM2pFqcfx3i6+r
TMfUF3cGsTZVYf7nRZbqpPmOg+Svhl58+QeSRTzuoFfhPJawSKoAKRzLlf9dULCC
ZjztP1q9BomnWREDd2JJ2RnOXxeDmQsaCyePuubzpfo7cxzlxE5D2FJG3K0sY0wE
dgONgf20GMJOaJnL9UcMuwAWbMZNlnqdeQmRRf6+r66Bqvd4tBOvxmvPffUdBXhj
KV5sHVUNnCcH6aQC8rRyiG89WabHwZU1kE5ylqxa51GkPdtKRrT34t9hCmFMhPQe
mc/EYrMBJxSX6R5/mXCBdKXdGLo8A9l34fMYKJyo4LFlY6XyzIPmuSEkLSSQXQnC
JQ4Z0sS/c2PggPFANgwW2vTTHv6mjdF484EJUISI+hsqWrLiEappqbi5GC7dsH1+
SoXNYPs2P4YOlYGZ7QfPp64Eh/6IriNZXO3TPGnzH1wMyEIvQMRxu+/a6a4fNb47
qjSUDuMFMyBUrIb2RPdbTgWBGI336n/Vi84qdJ2jPRouzmGnkRJwBt0NjRjiqhiL
HHVHKrqxfyJyvqHXyVRmPCseOj6SDrdTJ4WxStIUd32wq2QBqC/H3eIl7tvajlak
D7HobooM76m8D0/anmTzz09V1d/dsFNGdbDgTsdoes8Yesylau2g4ON2RPf2/n0A
0OK7gUBv3BOvZ3+Wg5cAYzVJylFdz0GsIaIkiVds+8h5wfGpRXHKeytAO2k5/QPU
mOEqV2rgIhmwrbzmfAS0IaynT/0shyrGRZAWKi1Zxlasj1ZBiHDBF7XHLgT+fUpE
+aJoBBRt0yREztmtZgYftz+d2BRASgAeIkd22QAJH+8VjRNGT9j79cTndTWGMOHa
NCiVZ6JmSuODdOf7NqSphrrSAnJ4KugCBkEV8wzwKNj8bROPreFn7UHcJgbn8NH5
bAkTmL3O+N0hQJBYWLYD5flf6uvSWbp9frvvqcy3F/CmSBCwV1Rx8IbOPSSCmtXf
ZT903SUBuOM0CoWxlqgNCHWuv39BErDp8NSFGM72TSGXmiCjkX1F0Gq0hskOQ87N
0HawA6oOiuPCxOE41z6ulS7Pirxy04Q8iTXEIrFtcuKdfFAwmEBA/5L1D2CZrIAK
nKg9FneGX21iZufVcNp01jP138crrWg3W0drUwk9Zr+39v3EOPCP/3GhPfPSmbOo
SK6L3prU3PXEw0D7UCm4I73HUpC0hAsnqcRSQnCDHQtShdQKhPgcDJkYvoqUNdLh
ABGXSlkH5NRt2brq6frzKH5zm7cmfQ8bNjST3tW31nmUjFFVRBoRksxfR2p8zy2r
NgGfLwqMOoNiODoZ3Y2vln/XUsAXKHdURpnrf4kgx1cbl9ZF1SU7jPTg/Ixi7X0O
YMh8IuDGtMfeVtgmbXGl8Jo/C0VgAdSJabAVERKBniXCWCRl41Cu6XU+WJ1pYztJ
hcsjyLWPqlVWsjb5qaVUcxxcVmnmApjs2tyeFli/gl1qY+kGruNoy7PVEoWyeZNe
n6ZjcivTC8bXX7DvhUfVPWk62ynoJ2VItBiLcChb8qdzwUEtEtIsERPG8e+RPofX
B3kwmS9XrkrUCbpsGC8eU2pb/nl6ARXyTvyuVJb/cK1uGrDa69SS+IqzU9T2WaPO
nxrm6ghRRi+Up0V3vUzk/PvAilGbtU9JAcoEFffo/znwUNH3X1y4DrlM0amrcA4+
Csf3rC35ltLbwl693zSIfrosUKt49pXAD/yNBeJaOo3eXLwdG/lLJ4JKDZL0ISU0
jr+eOZNPlsQCm2aNGHUvsnqNosHAvRSSt9+jgIZ7kx9SrnM1KiMKvIFsCbwTv+r4
tHeBC0KiN7/tgv/y/Yj8r2jTWcXREklh9kLZmwIQS3pnLnbaH16OY0iYWmxTSTZl
k2LMbcW/mF404c7z6sSgQ5wU5l5Ib7Cuq6fdMpJMY78h7RGWYwYumnXadaWZQNxd
sfBWpV9kjIJU7E8nnhy/g3+vkmybQ5HKJDPJDXaWY2/qsiefNg9aRGMQgru5bPN/
IfMoHPk9dQMbluRJXiTEzNvCe8MGBN4r0MlyO0GN5KEnNGfAOY2Art6B29LSbjrl
FJipfbi2Nfkpth5zJnyy4eSnex7hIs/RolVck1UEG7XA4kkFWbWw77A/h7oXcfV4
3qVstRotss6Fqa3y+vchUwWlmMzO9/54gyocqP8dcyggYEXhl6O7tnLurCzYcyFu
jyD2zQpYdAXIXBXA4xGaq56YCxGKDIcAt8Gvco4CHD+jQ/rcxP6SJvNBijDTihbG
HmXFlWh3sAlb1tAJhY33UqrGtFYim76PrCdZuq43k+j6D5dkqGgmYl4teM9hpFM0
6ZfbjRToJKxluprkxwn+8LMgsshnSFjrMYSeAP3U1Qd33qTECyFaz1sZMkO/w6vL
S90RBjuYvyJAaQd5wd9hblS7fYYVKhnz1nOiZ5AydYOOdfQ+kE2D/IEj6t8TwxNG
ALizDuSHPW2wp24KqG18oq9HufTfKVRCGcsDG6u91HLKE3ZnkTUWqofrpLSdqWVa
rMBnh8ltu0/pUJl1nSgaA+1R3YC+hzqGOzNxIGlrPr6eAcXMurPCw8NliRmSrfRu
cU9/ZVlkuchsDWuD4GLQMRtGl4BbTq9QbZCZy4hCYe8jLBVzJ3Qfn+61pMq4gotA
GL35NdOXoWy2+qPwOzmmnCmSMcTXrjW0yfjZZMzP1Hph6aP91QHetmdtoujrDivy
bGyQTAx0eTgDV1OY47j4oObjkD2WsDdZggK8lnl3DPGhEPv9xIGv7p7+YJXMEUPL
QDI0MZj5NH5JrCOkFMMpPtjOlCItsZEQ+5XBAW6qDv7VGUxXRFu7dWnpGj01Q23r
KaI/ZFdsMZHDtKoeTe6sPVUpyRP/7xF7eJY2g240X6ZVGd5gMj/F4vqwCFy/CkSE
7Q3C7LtK38zBehNKz0syr6oXpYMIh/VzXVt0Pn03HUxOHGKpF1JgSGZS2mc9ZiFp
DqAhTsrj7z6xnxnEgMuxJOVLqt7COND/WwjVACpu9V6Wy66claIj1a+NntbwCr8O
2q0ptEnuzDxtm8zZwlnntgT5aviwOsw9zTheIabNPYpukA0IPl5oJyI0pNNbhan8
3UZ3aRgYt299he8LgIwNH7w5PLeHOOSH+wkV6ePkDG6elwpito6vwFXnhOzv+QAd
5fjk1wz4TIoBlmKGwaB7EVx4nH1p1GLYpNyTAxotU8NLPImyzXOvSxBXgnbNgZkn
EIIO9e1BFoPShqDb6hhCMWeXjXb7DD8Cj/19hCGvtSsq/Dxh5ncpkW7HYppnaWb7
n53iWbyuzRgV3XjjBJt357W5nq7MeNy8h++vAht4HNurJf0Rrm81I8YJlnPG5mq+
efRSlaPnoBF6pbFNQnIvKHeWoO5fKv2GtstJat0iafuzYoSTessMsPFCoW2ocaFi
hnyhDLxFI59gT/r8xR7+IBHVnsFNrh7WBFLOEJffXZOxnzuP9/Oh7KO8KboyIcLl
cddzeCKRDE5iYpMvEqq+Z9xhgd9cGPgA/JOr9Wl4/gK7sevmLkmzJJTAdYEUuCNQ
pmuurD5CYSe+MAV9o70zSiFRgLXBqT20Xxe7jdvBFbbtQo+fRgcbSHKHTYjRxref
P6aXJNDSpUKqGxrDcI1o4jugIon45ePqXiofAfPxXKU4EeNVeflDwDk2/gCCZTob
oMbmduQNRMKfABeueJrEumbmpz6D+puqHtp8Y7gzsZrrEpaw06nKSrG2ZqlC/vNw
T2E2Kuz2nJh9z5cnFooxZex8GwNzll26m8SfrSdFtrAQww++sN5ads2I7Y+mjSfc
XO04r4SddQdXLgCDRjJgvKvyAneNLbJC7JSvBztbwR3goBlC7+sMC2DNEBgUUEBy
oJG7MuN96lOYF4yzvHYEC+mbIa1urJJpyfk/YjCm31RemCESWZL7LtlMOfWPm2oZ
66hqXWguiVSau25tKfX6yQXWvWKvrNRV74p+s7f3Ru+yMeKRZDqZfK1j8DY8lxz1
Dlb8NqSLNOdMzx5K2vP39t6wBMLVjnEzLWeTwOyQIZuFZCatkj0k3n+eLxIft4SV
Qjw9Jz6WCVy/ETWZkJ3H6FyDWVLmxGCYkh8Vu7PA19lIwG4MZMrA4i4xE6bhInkt
ayp/WpjqAItVErIJ1j8qorvfnh24Gwzq7S/C3o6mtshuY2YKNBWxc5SQTThLxDvY
Q0Z/ioeBw2MlPcxbpqNdgWwZB4EqTMR9PLsYuoGu7UQWO/uxWpqeqKPeB6th++En
9fLpD/VRSnoTpgir0FP09uVjnnvIylPyH6vky4u+k4A8JwywJYmc0qwv0dm0zDrw
Ge/s7+/AMKaQhRTBABlR5Df9Qn4qsoCK3ueGon/e2AaaqP5TxEY+6o2WhfcMp8es
hhPgOIkPDPmMeevhEF3by3/LAIAPYkU9yiW1qfNmKdeeCOQkaP0s2VLPpgnLxCjK
CPirffUiTsMchYXOP6YMhBI6Ds0uXdoohkME6aVO83907xK3IzsSIZmAktoO+EUK
aw8ChI13xwGxdmpxsLkhfERrCN1UEPoqr9N3T1w1gSt2rocqAqwxdAFxfHodYZOg
KbHMAB5Bfb9Ylal2u7SOXFn9hoy1FIknKyAjIglEb1nHYRfUmpbHPKxb1IQTEk8I
YM2yL0+QaYzz0PYbOJOql6d8HcN+HC5rw3K9ckuDG3+jS4S2ljIFnQ5D+F+5TmkA
gV1gN92olfPZlmXBC4LuNESFttbBtYnHenQbFbRC5casbEFX1Wz2SL7Nxv71R5KS
KPzF/crfDBXbbUGi0vULdQMHkazamiE8zcEEH7KAKzkClvKRVTgaKUWs9/I46IUJ
6pTa+2JgU4Ai/bRWPbbu0Cw6o2241Lp1sah3wvoP55skef3kND0noOUPCLrePfa6
NqFsB94fArPC6i+DHUTScHvBZflPheNZWn8h7qJxrMcrpZywVclbIggYHS3yfuuC
GL1OyGb+jy8EVYrkQ4CnMdiqTZe24Np3wqbY0vmjcwTZYVw3W4RTqgIUI81TrG0c
otk6mzbv2eft+osaOS34bxQqxKjKXkXY1+DN0qpXM6NzCg2ZnLRMOltrNWDxmkMU
cxOvhv4Ek8lhbMWhb8QFXOKmps1/nILh9zWgxgTLskzCjoQF22AipNMTinR9pmwa
8/Z4E1018dFwMMQ6oAqrx8iYbPeaxNDM1K9O/iSPY9unH58qzm3oLfLak9n45qFo
VohCUEu701HrlDkYJ20HSVGP/ECpl4vJKP4fbR6sb/SK4RTW2F66wSnvyISDevkG
O/izb3xEXXHnGS8Vf6If38D6mPHBj0q4DMUw0QavhUGTUDyowIVhMW/DzagEysDx
IrQJg/KvE/5iZ5Cv57CfBLabVvbSpYCfhrtFWI80FtYO1IwhQl5I4U9Cw3SD6qrH
k9YYq2sdfRNMRbOdpfOH7QHReU+jEOz9lFloigoUzyRQgl9KYKd7wnG/a36w9cB+
hL24StuBUfRwXNpN/Zd5b1kMhgUqArtC19+Q2QWDVU4ZA5q9a4ZgYlIMUwfTNz6r
kJDwyyDMh8z39ztPWNW8Ngz1k3I3IT/KsKJSdh75CfuVb0GwrBSWC2UUZOMxaB2X
wMsslZ4xUOUHbuh+A5oBW8qWA6MzksNSQy/Q/lUDiMXpynJ2JsO+2jUoC2Y+8eRn
EMv6UQqol97od/z1q6oRnr/MvbTLLZMkPo/b0VSS1VBuf0/t3Y3GT0IgBJ5vAg7/
5twF7Nds1h1VyQ6mz/AMzNncm/lp8PZFblPQdp7YPspMghKuRnm/QWBMqP751Xco
oPAtDtUxc2QWh4FJMxzLQ/+zwpf7kLXGfNsXG5xbqZ9FzMHvW8t4dwZ3y/ZrpcAD
jgrOiO1oRzvL1/bc4WFWz4H9wvzXscfhDpsKA4L6pyOzkMafb6tqJVlRX55HcOR2
6DJT66E0VDdg7hGVDKf5uMikhKVcRE9YJhyIZ9sM4Kt+HpUpkhWZKkq3DocF8Rhq
zGYQymVG4HLzftrKE+KqGkK5sndFzT4tmZCagQKgb8Wv7eAD1KYHZ/kYx4iGm2yt
eKPIVFaTueTatXHefJalY8RmjicNSc1yhS0MiU+VEEPEiQE1FemchspLDM8CF6YP
ha0lI8w5hiYIcIrRG5PFc8BQ30hWHd5bUHzzMZ+vSeYOv1XL5oqetmBcKkbDuUeR
8Itg+WdR3Em4bBIuELjjoZ4fXs11L/pnFJBaILFLsIZbFsU396Hsr87VUG2zpHDw
g5DGwejWkrOPDd20pTwY+oiotx5/NixeXkaYM8a8WhtmCiMplUSads0/Xwy9XwsR
FDJD4ZQVd8LwHvtTGhHjfjNIMsIXxERCwRk22BRgtwWA2z8A/c9N9Sh/yU5h460q
PXegfuVEaNKRXxdoT5GKuAynGXo9nr352Aek9IkqISLLzODE3mdmskUMUNVGBJaa
m/F4JjB8JVgp7cDdhzDT5QidChXYAh0gOxMiK0NVNqvGeRUDwLe9zVS/AkeQAmr5
U2/nzT/o154/UpVei5NDlmYD+2K7Qsst7oRGE6hIOrch6nF7iSi82BSi/JZEpX/J
W2A7AkOKtW7UXujVbasJBcmra1b8msf7m1EG3a8F5v+vMkhLnLgh4QcLuQes4C2H
ow4eEd+vEmSw7bno/cYi3JARAlCj+2JmCQ3i10+rnROtxq6naztFLdZCV7s2Tyrq
a/8BcX5QbhuGpv8kUJvAnG6RkG+HlAjovABGqj7SuDpZIZgLXq972OzRckgpymcv
gnqjHMgWGjCpMYDxACDwlr4jQRMPopqMI5HZqxUGLdDiOdNi3UnpBrulIjgAE7jf
yG0ZJXcVjoiLbx4PmT9BJJRpTxIIA0eJzvo2B+eAf46z6WV8bK2wDeYizeIpIDHZ
22tqWnscsyqAlCy2QNNYDGohNtf7DVT/GR0OG/Om+oG4fjinKvT2YKfIW05Us0yZ
bOD0BEhqar6eBFx+hLz6dkrf5gKho+5wuMPyXbc+q91e/bqwlk6dGOcb+NU93kfi
YBcefEkTjbKzY7Ry23P/EYs4OHOaAZ5TaZD98MAZeLjdewmjtmdYH8VrsnAajLYV
iciGTdeag7nheC3/i7he9DTy0lMVK8F35RMKjB0kZbij8tblmxfoGOQMI7s7BgLk
ZTai61iu3feuxlWUkx6u3Ja39ox6B9tM6PGpAAb0RyjzMQ0n5MItl2nSyk6qBTFH
f+R5PAESfDMOvIv00a5AKDdzJpOQzn+ioQeINHh+DM8KtVBqsXw6T36UvQQLO1F0
+M1x9QLRZD+2b1zWYVz4jhhWTES7m9BpPbf9/rm0ADkI3Q/ZUSM8RtKCoi/W9n11
Bv/P5YOkjrsKDXgRLHFOvAp/76LBKbb+0MpHLy1nNMm7oH07envu/gv96qESPQze
KYuzrF0J8uZtDv5YEFJvtKdTL4TZDwhtEC7opENAatyaqfsiRokr9gkDR++484k4
Jrh+h9iHmoqrBQCqcjhI/15JzqeXUVg83fq8vhhpYaTxvVNXKOhaajTuI91HKVS6
2IZdFGJga3JKsZ0TN4fwmr9ifR8in1cE1UuSMgevWVimAOt7HMlgMRzbEjihBrJV
BCBeNFuXkokZTr/pLrS8QIy8oRMccXSRdBPS2wPWM8Jo3QlK2YnxSdTKTY7fVB5Q
TteQmYugnhlNcn2U4D+afvlW33HzYkAXFd+l816VeWt4pN+wogL9PLC/A02TW8UM
iudE/ZTYFxjGkAuzXZIV2/ux7Rjh3U3iqcLQIcE1LwOREpJPlV1QpNHDjpDzufY/
iI8c7BCokLCkiOG1lzP/z7Di40aMjdNz+jdQ0k2aAuw7lCo/xZ2S+bP7sXMeRw57
awIF2qoXSOWLt0sKHRDBMyx9bF3oTQC+sFKJySzZ7Y7p7klNMGHbb/AWcH5JLX9R
IkczFabjUYNco9/6989j2Sz81x3Qchl+ISQO8c7fo+psLE2kkSAfVNWjl5HW1f5J
UqKXVPPpgQFVW7OhCfpMm/15b3Wpe4TgkGiCkYrltSX44k/JVYFTCpl8I7ReXecc
V+ehFzMGZtALuzXMBjpcJPdGIEfkLq60YIfctGX5lIvLf63j+tdmB6G+pwT/HfBV
YYB52dr7nP6Ay0BOctnXxWGo2QzB2QaG6FrhxuqlOFIPCOfFOYxQFrXA5cDRLXfC
ryNx6dv5PR8otBR9gUv9RCti9elZCCMCRIDxGWfH3EdUAENJec6fUUI+ZklX4uf0
ft0C3dyuI35sgv+4z3aYcN65UizZwZZzxfq1Hrj8qHzNdZixp+DqiELu03gMgxdI
8F7ZwSX9qsXSsxLRUj1PA5LPk6hshQWyK42hjCMCXgM8T8vF9B6hyNpOorFP9Ksr
gXPyCApWEUFXz61TMF1or+dEM/JUSzJFMt9h4Un/4lST5vpIkyw8hJnyP1nwqbiF
ZVlhceyvEhJs1f51Mkk6lr+GWxj5H62eYdN/g3anqQvcogqx15hDLPVz6ITd7TAo
k51c6FCWdCTBYsmEZDelvQ5p7bF8qEAd0ByJWkg9mOntYBkKlzR/XGMkwbQsKqcD
CRuDt0fRxwFbnMlp0PWwjNovhn080qws0KrkJFMItYTC295q2PJh+70wn/8gmUp/
Z5I9z0z82oDYTl7UN+OPNdp7uZtKeyYLz6dINN5/ip54vavpvR4dNubFtIsrsQPg
7z+RG+1QHTzjZvPAHI2vxH4KEOu1Eq5JPLv0X/EH9f5rDYAxn7G1qG3jeuxIPBPS
vRwl7aVHn7dwn6HRbzI2JAnakpOAz6utKpoivupeQngGyxoBBtQF/tBmUUbBSFev
S/PuMLCI0hJiI2nHSVIZ9WLxVZqhRPXXKqsFk0/X53x0HKRsqVv32qg8dBWEANAc
cFy2tzFHLKFWLMNSwKnDZABwu0rz793nkHjVd4xig6M+bxzSYIWOyPVRIFIAbkr8
a52Cx7+xYXezuADfzTsA0GKHMrJZ7y73IXRGvzCS5Pvuz24WjFUxl/NWDdhGW+5X
B1sm3Vs8iEQ0W1n6CuscgDnw9bg2zkDwkWqqzo65pA9HxrNFHzJ9tsijx/1zMrB/
4AFjafJLQ6oKprD0BCMHfTeC5cBRVL/E5e9Vfzk3Go39MjdB49lWbW3bIUgdP8rC
BReERtv4qEUGHAhxUbYFYA1AnGT2rKtcb8sIX3aU3IpLehVpfj391V4JbdwbfSY/
cIb/mtIY4BdX7uEwICAgmVR3C4mPWLbNW26fEfpu3V8hWhGaD3I4mOl02ku9uO2I
nuqIfgMSsMNd6io3UrdFw/evXwANG9vnXc6xVZBUp116N7ZT5sN6ia2+MhUD+Pys
QwHwHw+flPSUClQuUlFiWxdeFc/4c0EN3PJ4+6fhV1CjsGPRzOTcfRwdXOg4os4H
LGgK+zzFKy2wMXi4cJhzRv86cubGgTNaTouTJ0DSQ49wL5B5rISjOBNxavgAeunp
ai9NrDokP0oOzWZ6Xvc6lOA5pbs5GTqBMyAUjnZbez7SLENmT0jUTIVnapNZ6lw4
lbKruZzVkCjK641zcTuWpoPUr4JZiYmo/teqB91IhEIBB7Ig4pP8V/YCeidNY8wp
bOVDkcRdM3AMBYF0Gs+gmDVqFt/fe4eON4GW8IeO8G1mT2fUDxb83zV2FS76ja6Y
iu5JVTdlEBZQ+GTNdmeeRx1KZ3Zgg3Zyi6Gno/tK7d3nep7pXnLWkvXJaFOnTc/Z
I5Rt2s1crIvYZEn1qoWHkNT0IZIFhBl9MSb687HLSzE4DamWWxYnQ+7QbO80+7Hp
uCu2zdx46spkUmfu3OVn6F7FgDVZoMBE6rSeG+DuzbYwt8qpGrIDUjsrHNE3hMfD
64p82zfO7EAuY7Z/hRPRxttcoJjYkxWKsn4eNvccJv5F0L89/fAJcNfjfvYcbDdg
dlRhzYuSwUSPr5kBiUjvjPFbSaree2Q9fvBU0DP1YuwcrwuZmoDO/K4BrvvGtD7S
WHasaRHKclcuMvQKyI6ueLl/A1UcSujlq6qPmQ4MoJ8WuHFP4H2bHw4i56ZEi9Ch
LlzOaYca/yTIFBgH5ujBrLNNpvnV6D+4kxM7jwlXBccB7t0UczpGDeVTPw/b16WD
WGQX/+80i7B6jzNiHkbRDKXsNKfmKOVmkzqSOJT/QF8m9z7n8XnoGp7A8BSPP5KV
P2OIp8H0fvDSGOZTkBteDSbnWgII/HaOeo9A3eR+YilP7CthIg2y9DHGqCXPjbr+
/PpuhKM+4U900A5M0Y/vxVpX6PLtPN8V2Rq8AkjRKlFITtYN3tLgtJMlhCZDCy0h
I98LjkkllIRWAYA/4I5nUH8logekt+LoUMXxZV8IHnMZi+lGauu5xpWEF6izT1EW
G/2WejCzfupi9tjd1cN1W87+0eUII/54Vp3lXZv6f19ryKnPB4PScxhoQPkFJCz3
mKrXEYWzNZH/97X6y7wym+wZmsnFgx3QAKBZ6t3EtunubN+lMQ10iP9dkPATAn5b
BVCJJiacEXkv286hDPoW83IsM3hDQe1HtkcujBYbKveE/i9ChPBKIJE/gh/ci6kF
MWQpxXR8dXeOr6sanKI8kbBHARPvEVDTJYFrjWfXalvQw/tL3XlmDsS2STvJkKMz
rPLosCIkA68fg9jlxySkta1stM9wpGe+U8hrXIshOUnIBIPazuUwyRx82r5RV17j
JgzTUkWPXHCA4WsEM9aTa3OSqDYcCwyrbwntSWYDQ33hzlqA9Ll3IXSkz1kwzwZl
OH9mpQ0O+6DK6Zv85Dd+O6jE+mK3kQoJs5CwkIpATO91v6JgAIbkQ0XhU6E/PRPi
9YAGTMvQok8kuVgh+O5VnXvM4zA6shtS1IT3yTCSTbAzZRS3BGblrT2JKLV+j2/I
L9o81GbL9XZE0yDz+lXMaqogJmlqixoZh00bEyWon7az3qhqUpEJqFU8I++433WJ
zY7niZ0R7DcVzCUTek5EmDhu2wDKaDOqsBFzVf+ZCopFQEcvh+Hod8O5WFt6VzQj
7sQ4QEjICuGKLjTV2TsmH1UNKcRK6reNGoFUbLFBuYushmToGit2V4xaWvUhNJTn
QrCmkOFCjlxlJVJXHuR/kRQBgCJZKcvGZR7ckGdQiwikL8+k0NHGYJh3ZZcMwyd8
2Ld59PDf6OOZUkLES6ASj95YcRgENIML9chORnIsP1yr1O/aVCuaPWhjjnlguQMh
ueRVywJUFIBk90AynrMvr4p1sXaBbh2WN553Dx1v4JJpGVRPyd3kuzvBEW8X5lFX
aDmR6PlygvPSpz8p2xj2m4ZOBf7Q3WTIA52wYjbpMNoOsgOSc7kPM1scJl0pCWa/
SidKF87Bren3kdf4NghgJwIOgzGS2OcUSVONE8q3iNjLhXYgxtMJfiISsepXfXOk
RQnhXyxaqjFvQFzuuh3Dpz/kpndBEfx4wtIXWud3F3IISz/a+a4xv1VgJXM9/zZT
LYe/VB99X1TX0Rxy7nlfOs5TSzq+Zd5IWaczIHhdPbf2DONVA2o6Yms/EzFsrn3g
gRtpHopcJJtlvOM16Dxlv53ysmvf53MCh4DOCfW/bYFvJI6I5v246c+diqHxpwDG
KkeNqC0SzNOpMe3V5xTDgytFkF/xYbOO0NEtg1sMPPsl+lh17yKmX+3CpsGNfr3D
0n3sIxPgk4fnRLPU4lH+QBrzy+Kz8UvM8nsWuA80KW5sq6i5Ynr7ZW0dJfc5wN+C
dKai0oWuk3gwWIViz67AWnzVqBPcEUnOkEwW1yeZ5aeY65FCES4bFX6EEJOuOFcu
yO9KMKy1gxwhv+hIO664MSKPlAf77+D4LxjAlm9viWMpdPwlDwUr51xj1+J/UqxL
OmXVACUpkalDY+Ncx0ztVSdugv/NQ4YajZ7Xn8KzW11uxF2UE2LC7QG1g5waVE+j
2Ggv3Idz6pIBRgzlkhBBsiPx+bDl7Ahr6eEt6c6Nkhk78vDbICkIGYeJTB1b/9kT
VvFcnYn/TsM74blz4LV+93o8sWmXvwBpjwWSGRCL24NbWXE6n7rXRvd690sVzqeO
vNdWj7T1CqxJDqzxIWxUO51B981b7r2oz/OlK2GjrtQnmJa7FnHMnD1yKZzMRT4w
hr0ZF9fRbxHa+7nMu6RSt/rbX0k+3poRlmw1iD+oULnFSOv7fI+3sbjh/kYv++0u
vwUAkNoiiwbTuuE2glFoyAoX04IdT25QBt5fzOfEPDqzvZ8U8P49M8dCxCS93q4Z
iUc+L9Qg9LUF+1aJv91nTdww0ozOmUjG6BMuqanNhpABAaz1EXpDKxNjfE4lix2D
XMtjOmB9foNt+7B9E0DPvsqFMKNIA1xD1yUFUvKBzlJSOboALnjE6sL0WUe5qoNY
yA+Z4hkSVB/2qhXsyB0U8coPOe73Ga1TYCJAwj+cOvG+UiouwAlK5Qi6qz7D41cm
tCU65YJvE1I8TS291yNJL8PoKPUXPc7mgdYw/0jya2H50TCBOrlmqbToxH40bP2b
D9+Q3mzjg4pfJSIHXWfSvzHHyfHoHTSvDcStSGci7GRZQbulx4rml6N2aIt7JjmP
1+0vnTiFI/zLk+Gw86ZMZq9AU37G8WU4RmeudOoUH/qcm/fe2OUzaZN/rlJzZVy4
gYdXXS2fbnXuhPH0/Nr8S0jKlWGM3aUNAHL/eNzwQSCedswDZ+CxqO8ooWs9nTZR
wi1QIR1QE79yBRatlyWSCts+LwGDlHJJve1CN/cGVO/BA86PsbgQqFNx8Yt+oIiv
mPQy+djR6WJe6zsJSvZq21qgkGuvclvOSCVj+WkZMs/WvYuQamt6Tkn3unc32B2w
Oaq9SHTYO5YtuMCGGM3CHRD1dCbJzJWiV3w6STa8xxiwtSn3qdQNT8/rCYWRfshT
k0Ud0nm82OY6MZHI5BHXWyfwAQstjk8edMI2xtDu2scCeAK9k1gp5Bh1eTIB9Boa
uGnQATL1xZnSBT4r0lddM8W5jmHFSMMBBwUtnhKTVsjg3/GAnL/yQuS5vymXTgRH
nnxyLU5eACM5ekO7Oo9egpKhCapdGvMM+qWZ1Izj6RMqlEanl+1Uxp8pW5OKJ+Tk
KWKZ0VBUK1AD/Of0mzSRAgnWSQbJQutgd9KDh0ha8FYchoXhfyLvBgPM9SC59kNR
xBiqTVrO1efF8GU142Z1SWwWM5MKi4FW/uQ9oKRqeMpWGHbMfDfNO/hSdnzkFlE5
NpY09d/+mXMmO8HHsrwptybVoPu9NBx4TAnVU34YUyHAiTGcuTioI+7hJXCW0fv2
jJURBvJSINZPWMDep5HCGjN24tgJcx1nwsD6G+bSReD/nTv0mkuJ5UzlJxpjAutB
hD2KRU7c3Y0UorJFcsN2rth3H1Ukr1XBdPHgCEBxrzHK05hQin2vMb+lUDRgfFCt
nTjzRu8tgYOxwwaQ7bkxZ2OTIdx3Ik7WdOj3d9qRouUeJ6THnz/oajbT8F/gcRPM
jbi5T2fC4/k5L8Xgw3KuJMymlVLrwzlMsoj4k6Hilm9OgNhk810O4eIJRvpzf8e1
WXtcyEmb2LoO1q1dB3BvcnBt1pUvVlsFmHQXYyl5ym+R3O5K1sHjEqpjZ832JJmS
JeCJnDWgPzpDJyW287dK8OUUWpvnFohtvPNV8i9qZ5G0eHaAmuf8qj7+gCrA4a7P
MfhOh3nbnd26SFHknIoKwbHWHDVM9chPnmJl+BZ0/vU42QiIJd+SUhUx2PWn4DBN
XRmwGAdWT1NSoN0iO/OcGb0bu82L4g2x/E2iJrq4uLvQ7w4xdhShkON/2lBiDRb2
IBWBcwDWkULC5gUcagV2Ahsth/QT1Uhj0OI4tugZi3hBCG8D692yaYww0ddaaaAu
mTbiG9b8/P8LyvNM0R5JQYCW5a2TuX5+bQ1e/Pqv+PAiC6k4uB3SrbFfu/1aPZcP
ksG8SD18lSDafdNvYlyQ2hOFCsrE2JM7QBicDIRyaPEnupDxmGihdWHZ16afgEhg
U0/jF8EdbHva/gju6Ymv/6hRX1EswACxQoZr1InFWAredkeq8noqPH7kxhLFXIwA
SMEmZEEVRSk1BOV7o/Vcn2iV756iQC0uyIEdWFzylrs25/dgvhVU/q6uy0F2Jyg2
+E80w3JkP9e5oczYhsh6C+5OJ5kgoFiHxrNpQfINy/SUzHQ32iOoM4Txfbl9hlnt
xwG9JQc2pLkZ++bHdmYGsyZ3L0S5AoZJSpDdWjUXW1fTWcjHfjxYGrespxRPxk7e
JKqXExpnLzzjESekS+YPlRuwKyauT36ITjkEV6ea18NhMazuBGkSKnWEe9yBYn83
0exrpmJp+vNN3EZgw2axt//Xs1eZL80AI7M8NI9jyzVFm3vT9CtGltsEa2QVphfM
fjLwnXY1E7vHIdYL3UE8CGlvmk4qk2zC8pktceZ8bco3t+2NByrPNI8/Cgty684K
5IuSGqTGRRsHolJgEk10U7FXSCaGXJyvaci0xZLqCg2RUi0WGrUlg0WwCR4iem5X
Lc4s24NunPXLCr2VVSG2YINjO4wTcyLFnv/VVzTjzQ4AAxgPXFALajIPydlQHUdd
fnEqYWsYnl28rupSR+RrQKHLmvQXuGqFzRwBEJlWtZNmTDdqWXtoBFjomc/LkhN2
ezSHvHgkAWyXkniAljjEAzOV+26LdvqvxP9luCoLl68htk6vYfg/6A+o13zImapa
H+Zio70ey6O+n2mMLgVgHYviM5zquoHare2UqyAwLQHSO0a1IUE4MitBVMnwf82i
W6oF2JePrG+OVAz/Kp9WVZJbGKxs2qgSKwZWmevjDjEiL1/QzHQpRFCHGiJ7TweY
gNZ2tLL856YHKTutsQTMRqRdmWV5SEw1lLD+Xzny8qutWzfvGViwh5tj8bhKrHGa
4nQ733tNgEbi8upyp6Mp/nZE+WQBynDPltuB/Wqy9P2JFmwuuImxqi2w25QaspZ/
VJpFuB+EuKghoGR0BlAGaQ/2AmcA13aj42CtGo6MveJ0sioG7/fqLlUTtV8ay7y2
8WrKcq+iODnDsbMMGzxjOl8gXzLRzo9755jxFmjV3dQ3oWdNLKF7rWOs8ySAG4up
JSUfb2iv/A+cKe4vG87yzzXU+yDk6FcmOhN8RSQaSznuh8C2ATqKBIrKLueUQvvG
nGAEkR/nOuHhjy9z+ZvBlKv1XxvNY78ga52McjXm9SQIm9I7lo3f/+JWL2BIqdTj
GTTAU6TVUHZWyR7Immh+s2X/31OyU8EiLSQ5cWXgW6cNqg37n0gPl5mYO60IJXZj
gBRKmcr8FjKgLWid1CxrafA9byDucA6CKsoGfERS5vUeIlENbHQOqLL70w6yhmsH
s53VQyxc1LRzuNZ4NcpWMPSG3gZMYhE3kfPlhFrapbUKyJj21sBcvWvvChtrmDg5
4Cc4NP/Eg2tGVc59JOq6cMvi9AKK7XihxA8raq8JJhrwZ11PnaeqRc80J7oe8ZUk
1XhEyXejG5G/zIyqQ9YgRlCTDZJ+7XJ7g8i9IK3F77+GyKc1IKxdc0N/zmQaY/rE
YCoA9uHvOn/YDhz5UCK4VSUZcI8WZ5e86RCk97KOs+pd0DmJ+sDTv5GRxoewVSp+
4NY39lXB+f0/+KIX9WfKayj5JPd/4y5pqzhvfCwwX6Deo9CA+v9kzOBJ5P/w0r48
jIuT8Fry9Odnx4kyNEIJGhwCOg5sJFnUqKDaiVbvhp+g/WfMWXuBHB1ayA1Mazv7
PO00tT2Mx8m42CQyaHGZDErWLxquTdeWPZ29W5uxhw0EcP9k7QcbhRU97zIHLmTV
axT1FuqJ9JD1YHcRUU6vMnGQpgxhIUDYB4Bx0JZ3nEngAGmLOF3604MalhahkPzS
ev6A3qrDC0Pgd8XS+XkVMaduK4jdfX3WzOx5fjdC2m+yM8gyOsQrO2tTIJTg/SSY
kM0sLc7/JK7+BKF34oi1t95qgUgsHP5HVLjgETgHE5TDaC7bms6hmMXnjpgyP8+2
zc9vMUmt4bIOM6+IPGhZlMQZEBrr64MvqgYE2IEBkqs8UcAemdo7VqY3bMp3e+Kk
SuuT+HzYi3c2I1Rs4/2mX916peoEVa74z3ooNMOHJoqQl8yVT6tMVOgbw3DeDTIR
SX0T5Nh+LCe17jRR/rZa7VXdHB5LNF8YWPd5s74OiKgAYJodYO6LBjmCa0Y/z1qV
Hzy6i44gERbgupgrgPJWPv34Kxgv+peXaeOtRMpVMU0XwPxPDYrH32J7Eegohx4s
OJW3LJc9xQmLig9lB73mtSiN2tezdqdpQHEra3H67saEkXvEFaXpmPx17OQpCTvm
7sh+VqdJTXYjMqqdlX8eOwnzAM2a/ATmFf9b0crl1jOmPoM3+QDZBU+yHYXbVwQC
xRWX32eUQjxI+d2ed5ljKQB3/dhNlydEzGVsVPKEZu/a1xSt78gn5yUVO9mf+Gqx
2XEidoB/cXD9OcaDLbnSfHFB2hYRuzdbuANhDU3Q4ZivOfiUGwdko4FU5YjK/YyO
1w1PFL66Pr6y6hSOIlqg0BdBgwbLGlxw3pGcHOJrvGgim9pn79qftVKElgUs5Hf2
JbkRD+CkdxyXCzFpdfPrOS+2m15GzdyG4zT6les7OFJTyKRQLeRMLe6/mDjz313W
s8spBhqDNsMpaGQK0Q0Kn0SbrJzTZVjZxof8YxGyYwfjEeOUlAO9thiYZR69Lg1v
qIktqw8Fg8Lno3Lb5k5eNbLOcJ0IYVJaU6zkz+KUN26df6b0ZHvWaJTz6kyA8WsK
sExbMyIUq8tTIxeXkZsMdwpxmGRiBUigfHoTTulZ+E60VFyhodaMmfmlIqMdGaLv
2cR2NgTkDHB7AMiUZTgG53cd1hBhJaJFYov2cyYbn9J8n4C42GTuPopIajgPeJSX
UY/5u98/6f2wQttsUpHh2Xos21wPiQOpsABLi+RRJ0L8SO7f7R7lzR4GRxGhb8r3
PpcrvbhrnAxJe/qRpR22tJuqGu8dJ3FDsxb3G0BPAMH7RxpN5FELWfw0ugnwdN/L
V3b0z7EbWDOM3WRCBSgU/M/Q4Em6XrJLslMD0hfb4iISKSnKBOl6mHp6+zgYfEFD
eAf6+lT31H9xR8EeHhoKtAfMdzuldoE44lUj8NDWq9meUy+/WG/3juMwllkNSb/q
lRUFWm124maKBoVMud1GmQDBAB7MZY1+nU0TCGX/sQBlq3ZVyp6ir3ixKIgloJ65
IvtOBAzSTUg0kKCFPXWLNMKr0Uq4mXjHyssLrxpQqr0z+tBIaes7Asr1v4fkmX0u
GyR1QYIUYcnilKtyjQcgYIeerR5On9Ai+0rbaR920hhwyQwq4Ei496qgBZEyAAfY
AWTV0KfUMTu+as1Wk70LlEYu/AtfEvb08pm9BmlQlnDdQKZ3o/BO0IBvNZRiZ+iG
8z4a6/mkvM+xtuSZe4UUpP/v0qTqMFdzSii7zLGpsO4nAH46+e458eJZ04AkXw3Q
NpZuAlnvHt1W1TeIXLQSHpXP7tdjfxgMdsNi9wE64r0R1q7f+elTym6yiCFd99TL
k1pDVi0Qj5AxZVD+2Zd0miNRA30/zK+WYc5VL4VwpsHwnIIFQGCdKUOYgkCwkD38
gfXzLvtDlal8HbRWM2tWRuceI/Ftv+dX8rBI6s9738uo4FQQLN4Isyq5viWnDXAa
lzkRRuph/PDDRsgjiMJfFsEXENfGiglHJi7wBGqTdNMNk9IpOW6FznognehaZQcG
q5jOhrYdHz80Px9I8N7BYu2AYaoeseI9MlX85WX95giBFLICZuYrxJSKCIjO1Wt9
RmfJMriKcPR9Wzxjonb4YpIrH84uHSB304BdFMIM/zsqemtQHREJLfH2ARr5lekJ
EXnm9MbXOWrPlBKcFKxuUfZ7/ro65wrh2kMxZr5k2nZnQWeG27WIVsL8kA/Nkab2
dR+lr0V8/fZ6Il3zjd3xn5Xc9xKgti4A+olyE4Ds7IWU+gNmlPwcEfmdXmF/ceWS
p8DARPTm9xXqIJErG+FHkQAvy8vAdvXaSgYGy8ue7ySrpeaGGSsJrEhxvFlc6IRi
w3Yo4xQkS/UxdJwtGjw8MTyP5wvBOT9huyf6kjUUdQ3Nyh+8oNSBcI7bduqTMvqJ
Hh68K2Ru7WQ9qqpLmT6MiDzlRz8kVBeQ2juNYcHeXypMmXVhO/B2TQJdZYwOaylj
Yjxcj/D0krZrHIB2QIXU7zV8huJ82WOjP3L3QfFb2KwUJMSJDts18Gjv31MgPxl2
/ve5vJl2mcqBYhwJW4al56YrErhX+PmEJlgOvY9Cj5PJeFnYbgFbOilAFAOYPfEP
H5VaCljK7Qb65MRCUzw0Kbe1a1wdkLqAdYq/F8QVkARwiCUuA6DOoLJFRNKuJapM
pnq0JGghAeDC8hXWXPV/aZtYXlaWh5VfYBi9DRE2cUOpZnZG+tlkc8dsdGLvMa90
xQoaEicVEMGYyF8nb6Y0uqOKGSarjGmgBf2xHYAOYNs9/QNG83zSc27xZNA+CUgY
05S9KeC9FfpBG1ffSBdHGZKprgPdu/KRBoWfyVsQ6vVkizYNsvkNVlJ0UUKBrSxK
JaLyy2D2hIuPXhRQZxoobIPxO9zlIb/fqOqA1DO3wP2dK6GcCkR039GtPVMT3NYm
w7S0suTK9kcZ924aOUpZgUYnjiHezxB1BA9ki/ZwQb0tACwSTdeQGmURSSnrcMCY
UcIvGEaN+90pziC1is42bf6I8FfhDuC9mbQxntAt6qGuXgGgSyBBdDJ4UA5BHWuz
BnZCRLpE1IhqCySPe15ojaXWF/i28pdSKeRO583pqfZPiECfLzCxpImbDX7afVQf
CPLy8pOUJ1COYEuGLf7HqIJguckd97YYgyVdi6IIwxhLFA7oOm01t8sRSxBeYO9/
riR/EviZE6v1r04QTH+0pc341A9Buoz6hXY+J6nTUC4PGOaNBZxYpbmCikeoqJvm
56MatR3vgp/yTIomnDyi2maOiVAFq4Rs8poc+zwGUG5SjbZjxZnDxleWLeLUivcT
WktRrIXMNlM55GUPrubMvNr0n09k10zFHCZvQyI+MRsuNdWZ+8afyfwpnc5OOs2t
4nOSwJxgRkKLwF0Df2qGPSNvmwDAdCFBTT/EijQVLdh0add0XI41uy6BmwNJiD51
Ul4ewqSQMVmlW0IZt0Hc3BWuWlDDDzTx2K0xL85TBUmBY+qteI114+V3tnWKBXSq
TaVdI0p5GpR4xB4m4T2UwOzhPbgSzIywmDalhbvNwE7SAeTDkz56pNrzkxswp6xk
MFyWc61DVJR95a17eQWB1+qqE9uOY0XSElhMmI459RAbmOQlSdhLfJE6/AGuIWUK
rIf0QKZzEBiptTDA/1alrCyZUIj2ipoiuN/CxTfwvBadbjMIomif+loRIPfeapKZ
779crMxKcP0ub3ifKF4FlYZnDJG32Rxd+0LCLfNtWrQqtNICZPxeUA7Ao0ZptEha
JvxCEt48sqZwme6vXOfN+gAwVeckLhMR4f/AfdcMqXej7kM1H5FTq2xeMQRGDvK6
yAUDg1bXc67fAYX4vBYiygslqk1/go++I7VFsV+HbSwXQW7L9TFdLc6BM5U/ieuD
r4tbjiksH7WAPA7ADghvtG9bUuda202JXZ4BFW9RYkvYbf4gEy0nV1ZepxjI1O8c
hvr2CooKKAulIgUkpbtajlOVmykN8hwAWfkw0nEJc43WzsmDqhD/FmpvD8sLoRsm
nQFWWgjZuqsY22hhEw6GjdE5i+XijUIKmiB7wJgCSEKLvHA9iIvBlBgHNAdruZpJ
/ikTBsKEbY7CQFQ9wdCIKOogTmmBsLPLzdsmiKF8j/hAUtwBECQ/c93eHh6HFFU9
rX76e8nJAE6yyOtt7qxnO6q08GMOv7x6wsDedXQ3WwYbHCsXgALdCTOot/1NQ67i
4oB9hE2MBC8lHQ19XNX0kJE+djSUNfim92UcDCtIQvGZE1Hdc0iKwHXvzXsXURsw
EhhIeeyH70gJUfud3U1rSsHnHQbfioIq20q7vYsDD1JeZuANlH0plToiQuP3KWZF
JkOuyM64A7sJxJBaqQ5rUzsQ3BgnAUgdBkLdtUQoZq9X+Bzo5ZS9n1Z5VLqAKcyY
KwLJnY6rhkgIarvt0/5fXN3YmGl18Rns6NmmvEB9c4u3z/xgwEK8mqn7gSZYlfQ2
ZNvoCCXZ2g5ro60Id/EkDgIEe9BGTrKF9mOv0dhub/eFaBJyB3zNczvOjhJixUyx
STRgUwuD5mSfndltlkafgiLIMxMtvo7uZh+SyzbVom1ZoR9ji3KvRdB1vKsGVGX8
9x/tdjSAQAiPbB42RX7SCcsWea4+7hqiVlgFiNFzkRFa3JJNqfjSSRNpagbVgxHI
mpkTt1q0N91UpyNsdsKaix92sgN3UcC25aD+d6Y9I2gozvYYzErg5yZvYVdRzgEu
+Xqov7Q907OlqsVJ0K7nY7SfyXgPSKp/heq360RbkIfsL8tUEhSdAHPA16hLgc59
Bmd/a228BMoQr0ABKGMrXZ7HnY67XgSI1DejdR8JocCdzBdly3fI4DmX9VeHq0uJ
2tnE1EIke+uKD1rUZDE8XW40vt45N1I2oKK/Q9PHGqywKtyVsdphaqyX0bLgNf/x
+fdpv6ZtCYUKzDOPWM5rl9o3UE6iDkB6bejDQ7orN6JbUZmGv6a+x1ytUvlgcE7/
3USWeK/fD3r1iydnjW7LW/G9xNIdtLrTQDQD+VuMb7PymsJycV7Wr+XNFDOXNtLL
oOwXCuZ1R0Iid9XhlxqPS1T+wVQnu2Ydd94Fuvo8bfBIvOxlqPU8y3lXE0tISWsj
jb3lwsfKahq0za7CoNWXzVMfhSIcBMn7QjYGUeSajfHSJC587iEWX1bOG5E/+cYU
yelZIs1w40vXkevFoHCZIvQn6gWnvygha+juTD8xwwDk7K7+XbSSUSPN6wFTirlT
Wd6Szr/BSrV5PJn/xzGCp1XU2tVLDizQb+prjXQJt4cWga03wnHxBvPxWZ+KwxUS
l2JGPJH3brCktW3IlbxF4QfWYxH/AK0HsjE/rI1p10TtAU2ZZixdZMZoGCNn4mNV
B2Lmxn43jv149PRZjo0ZGkOcO3L+0GLQh4jQxWTLVPLYUCyTm36KyGBCnu6tA/bN
M7b7gJlqFaHeB2sfvK1nqKP7DTpAkhn5wIzWZU8k5/dquM4+fbS3sh8cmMw33skZ
Qpmygvb0xSgtQk9ue93vjs1Dxa7x97G7D74zwGH1iIJSJSo+YFKCWj9NvUnga1no
bVAsiBMu3PcaMLz0+aymmcQX4g21O8Or8pPT1hUCR9sISoAIk8oCz5AMfjJE98dJ
+qmTqOnmx8myLupN48u6kpkaQ4z8ZilWxbj7nwvbjyD4qHIoHI96GhkqzBHoHewm
CSxJO9+0eJ9hhvrpvVrqJAWItuj+R353Cc3ttuMAVbxA2saOMMN0Dg1EGHO0K5ho
bgfL3Pq7Wp2RA8mDVkBMIRV9s6hobjQMi6wkoDwHy+vsmNqB5PS8GvbbYHJeFsRF
c8nuldXW03SFOCuW9IHydRmC0uxj/+PpOLYz1EG8SOC8tJdwW2F9acCq7Gzn/v8J
DHgEkMlvIo81/CAei45aIfHkBWwjgL2P5RLIRiVhkOomQuSIZ6pLjqe+jElP3Ptt
qx5S4D2L8Dma+I3FikLvCRRVIT8oktdJhrNfiFAd9K166hqta5AXDWurVDE9O/3G
MRh9St3wZoQxsSBSI3VfgGUHweCBEnwuk1IDTUcPWId2CV/6/C3uZqNhKV4Yt+mc
jA1jR78bYb8x7xdLjW5nUYqK2LVEYi55qhVomxpUrBBncUcmISd52x60RgF/0kis
Km6CyDFO7k0wqM3tcjcQw9herPbcJankAIxxwvnPsnmZeGZ3SVaMudheAoQbhxoV
gZFQxMJzbO/1dX+8ZHSkI78FE2tT57loa5P5LWk0blmqZFgnK1gkwO5iUPSKliDC
gxKvZ6bk1iIuhBbk6asT2ZFnBwJ7RRG6ciog60nCfJBoTnPIVQnf8q+7oJ9ByWih
EN2QxD9Q0uozaeyseRXXK4dPOn/dLyyRTeP1ZYBNF/aauLPQ5WrmBYdIDv9FXkgN
+qWo6HmR15/87ukfQHd9uVSZGeqxUcXud2kcOeWg0MhKn2hQxVI20Y2QRULP+J5M
JF9bAiQpkVWSqpG/3YlDp0VmUmMzZbgKfR2BwLePip2gvoyO+RLJDFhNh4kPfK3Q
l8D3NyfIX8Ek0N8dwCJgFVm7KtjG3ZVyIJ0e4WVRhL5ntN0rDwPSxsYuAGCcShaM
SZ0hHHjytkmuqXWhHsV64fyTzod6GbgstD23GDqTZUVNSKhLr32wZn1cJLrxEuhe
hTEtnWXodf7TdNZIyAIExanllsUYgK6WPR9Hp+BKZw/Uz+xgK/eAdp/hUhxo+07R
zwFLpmmJWlYsOSalJR1feKRkSFfPHxLP9pfm6otwyNyLa+H++eyDrQ5Dz+zj+oWE
BB/ouYbEuyrzc0fKbetDDz37oxF4pveL9LX/n6Q6MqnzwR8He6tFZs5RZWZX52n/
kEJyhkJ4ZX/hvvxMoZX8atT1sJlBzqx41rq6hRsTVZo8i4KrSWXNWjgPEqnk39Gn
RAAz/wki/T9AYFkyFKiYcVKN+OE0iEF93BvJHrPzOCbjpjg5aJxgXZVv0zWHFCMP
vEBaJd/oJrvCYCVla0OoT+1oJu3wbMfaG2FK/AuF7CjzIfcnLHZWUYHuNH24RS2O
EUOuf7lGVbE8PF8wN9CzTSjehWKrb0D20e6OSH4RTOBeZFnAq3JvPI4wYzZLIhKE
QL8Z3/bXfInD2G7j6mpZDCUd0giU8+Vq39S6lKZOxrsP9YuYzwLamsq7/w3KFTvN
kc20UtsTsi+dBV9GMckZLVfLW9a0l6d/Qs0RTn/IUmQ5vZLNrn7DzbovpSwgFv/5
Bm5gptYAolLDa2cWXYAMgSFZZU03oiHmf5rO79IB4Luj/7EQSAvPIF8KQetrqMeX
d83knADsc2uy4l7/c7O3EXn6p7fTkm5KT0qzfLDOQ9ojLNJ/6/EPrlayaEbiV5/v
HoAe2sOohR75gaT2K4+haFNc5/tu2itg425mC2yTW5dMVFwu6UWdY2ZEUrUd9t4H
EqAUFqlRLLx+UEzJiTPtAJNJSUGv10dFtMWkY/c6jDfV+2hQRonn0Goo57rbLxqu
cmFXK25mKuW6s0gU42/QNR+Ty0C6JQlCxp9Mm+3ffLipkHmRNdGpb8gnYzxuOp8G
OXcLUw/9BVHZG19K/JK5CyS++hd3QN9ooO+9YSsuFgFj3is6VOSpIARrtL1x2fmC
ExKFTXeidI/QC1+UUKul5q7brAgl2Tuqynw7lyLAjYVwof0Adas8wVZewyX0Lnve
EvqeYK4fh1JTURmAYNX8Rw6zFHWrQqGHHeDusjK1ZGEdWp2NSEqpSimTxAdX+6ED
Q8NTaZLuSgdLye+BwJr4BJoQcbbWz/Z01EPEcvIsWO7gZCgA6PhYeVFgAiBH2RZQ
T/s/LiCj/mZp/AcG7EPgZob5I78cpaDHeRyfv9joS16V+hsKmYoo/fmER4km+aEa
M7yLEjXFjiJ6G743xKeSY/26PE6HAFfkHmLptNdyozxu++NQvZOJxt8WLT+DHyoA
ZDlZTSUQlWy97U58dwJ7kSpVMeEJR0tqyVAhL00VmGYusWg+6CQ7g3Y8CPW6NXcj
JMiHscsJ+UsCGB7kUYH2iF5hxsI7v5G2J/97g74y1YbBd8fBVBGtahP3iRiq03tu
xkmxj/DHigPcfzyWvDPXdqAgjpjA55wRqdWkb4RAXy91JejWd43FVSMv3uWiptEs
Nh73dvdcE0FOONpnLN3dRtHdGDiirjupkcPrdMAKaZ1TN82NfaGxxjUM70T1kF+U
5QYovKjGcnps6KMSj9L4O2Oj3g5bCldX8vNKxvb4tHIdL20Qs21Ycm6WB60ehgIr
IS35loDeXFZ6JAk+heK8ITdfCM09ScUNGGRTGB1jXW3cnd+2U11xp4DyDYWlD6O/
UK2828/d+9RCDpwje9WXT3EnFN+2PVdOLZq6Eg43eZQXF4+iRt5mqieqxChTAkO7
a3Ejk3Tp9nuKXw7EX/JHDqIr9oOOcBU1Ov7ql/W4ydyAlkEQpZ/ahXR68Ir9eV9z
QarNukpF1vD1xJQ0MuPMKWIEHYmEbod3ewFEMnOJdVDi5ctrt3UaxshZCug72QYc
k2XOyMd3krg/9R48IKmQ0zEEI70tl1UStvR/L56bI/RO/p7BFDESo5/Ox7YRHGp0
QiaIwxM0xHlcIpf2tAdskNKXahOkYI5XrBKG0x5Jb2eI6GraMyGjDtSmZrRMGee+
PyM2V93QFf51iSCcTUsouaLV70w+rSVdBUS+SmQdmGLYcJpOK6x6sUfmzkBVpTUg
l1jWnw97eoSYW5a4sW26df+Eo1hdEIR3r0JvhkX+RLwpjzN0EqvHFvW+ybtJLzux
pJr2FqZvUo6ryTZZQjFt5Oq87x6pr8skdqApIPCBrVkaryJrkh0ccBHA8mgt+G0L
O8CKuuJfdXtOtFeNFX/lfOm8UmoiYmveAURHrRrqb54Ch/MBcNq6Uz4XNnHNoMfI
yG+L6ixHGAC3Ea5o/YmGWOcruUH8EWpwQwk38oZsSfBOS1SjHK5On5w0jmMXFJF2
Xkf8a0wxBkebXtDPTwfnGwBqNNyMpq+4LZ0M0wITtlIblpyfvQKzsNVGDH5qVbGk
X2XydHzEb5EESjniHg9yJ8t5xJBJCCnUWODw0mfVxiDtvdQRQrtocIcA2YSwS9PG
tVHYIkB4dK7YlPxcB5GlC3Pbn4fupKLpkx6rOryUq03Jk09E7tzceryP/yYoMjiU
H9DozzZlUSdtL2O28iMXFb/ziCdt1RLuPniwxR3lYitEUTikVtj8Z7qFsqv9Z8Fd
Ob6QdPnbjz7t3/1ig/MxcZpHLFqV8ZVjHZNbRn0jeU30TGm2vHvOW02/Xx0QuiMJ
77RD94py+KGnziHxB+3g1BBxeFDq5AilWPUQRPAtGlpOhfepW5Jq+0AeuL+47RKn
uI3P88WP35wbdkJX/+/bOWccKCrpoYkr3HO382WXMB1nOIJHDgrpB+GrQTvRuq+p
Nb5HcMwh57oGPZydP4PPCRvM44hjF5V/UcJGDrsnzdS7AhRNwqbw2wfdAUHQjrpP
pKIaYhK5MSRAslJR07tOthq97mSceKEe/HCbcMdHen9c9d8KdAcvafljTBls9e2f
vdpU8+p3sq4beY9wzjsaUV+CliirNkiift1V/WgAInVqMLLjO9QiYf/p1403IofT
jwCGT5sxygAky/7N2ms98aKHCugRwCh4AdIsgTZ+Ycs67zZgBnYFu50n0WRlQLTY
jhGKHXyhApSvlMB1LW19f6Y3E0TlXljFZqqxcDCKdbpKmFcKeSJbyk6WtrmNcaFu
TOarDub4qDPmRWI1pX6Co9Xkv+dYEUKNPLsmhiZ58+Qy795AzWNy2O0V4lk1nedp
5+c9R6ZgfpV2+csvhFCHqsIUfpaPkEi0Ok//+Fn56cQ4wUp8nG2xNfmcePJFNf2P
mGg0j7XznAuufKOq9Zgg3kJ1c4M0fCoOVydNrjbLIWWNOtWez8aMR2pShMW8Fg9q
3O5wlFWbo7TRng2Af7//X1MsiwUgaxFRI9B3vVsrRivJxciU34g5OGDBHRfICziL
Jkghhs6FGnTJHaHMpSbRV9hcE+U4fqaOBQ6q1NgqPce0q5Ch5XpAFjFLdS3zJA81
5u/cow3hjaHWOP02+gCAcxdCqWDrWOT6flCf+AclxFKR/yuVwiGqymGwUCZfgTCL
GrT9U9dXcJ2SzFHw0b25M5R7VCi75vuuCOXudTUB47jYj+Gm655oqal+nEStkbe3
0rJ5sQ7fx5U2iqJbBI/XjVUWCbhSZc+EFlZvpv5jxArD2XG+hDuJYxqeOWajBOqT
auEO8THildXfWBJMuuA65knfKkIXx2h3+iKlyYbh04prddfxJxxnsDcKfXz8pXmV
1wLagqG1D5EG+bfdIn2xJfB4XOHwwmvLBrgofJKTndWQPF7POecE/CjAUYHryoEI
lAmsF8kMSlpSVoIuldWy9wBoa6TbF8iQY+K8H8zlxj57oZzYoxbRlvt+rKW5DuGF
fNvaAc6JEukvY65W/BALm5WeG6vi2URknqvvRAFN0yfHDW2kHQjlAdBFw2fuh9Oi
1/2ShAURmHl35RfZPy0c9nVKWSUyUoOEwWN3I4/QOtSrgVdyqq4sIXcC+EyMBgDg
8k4T4TThMtLN7rqUNkHtqWP1e3AggOD7hLOMtW60otr5IzpCcP6Rw8aaHs3jyDTD
RTxqOPBA0YkXnMbAOILnsib7CmWhiCb9buRFeOvB9UTmgYFgSLXP/u7KNOx+WCFJ
eEhDvQoq19r2EVuKNl+iwEfcQdqpB8Vk4QUjSAHGjLcz/Hvtugul6W30C0RsDeXt
i8k5Ht5n4Cx8qyglDYwN1+bvBOcw95Wu6RXkFU0Wa2oI5P3PalISCcReX5BtxQXs
yo0iE4J30Z7jJTtfe5r5mayG4bVUWxqIcfpG4Eotc/fhCi1dxffWrctcZiAzDDSp
Hr1A5K5V8mKJtge1sAUCTlOoMFaQO5h26qiDtYTBaPGQmWSND0xyfq/kHbHiq2r5
ECtKsKGyRk0sHrYWAdPeKk/zv/NkvVoP94DgZT63mZSx5PJn3bcboda6n5EPrPwb
rGgrvDbjQdyS+SeM92G7dPXxb3G3mPZYRI21ncHSnmjpVDh4d5J+xGcMQp3Sq4Wu
uRNhZaHwGoaiyGbpwtzscWlVDdhSOiP8hDn4X4WKyZ5futugFcFixGV99rLCAZB/
GTx7fbudHpv6TLtOM/3oGqHoNgPEscFL2atWAQm0HRPuv6UMrTOmgASq9ZB/OaZG
Ta8TNRv4oTPPAeBW7ET1SvYDcz1nlYJmEVhijVPU3WkjhkMSANxSYQd7dmKI9EY5
paVHWD3FO2DhFvqIbGYfCvlfvfJm4L6kYqju1bj2u/DvEHgKRjImS1xnBG1106Ju
QagpAFREouNyZ1vVmuFqVCFddVAy5wy6UpzhGU7doqVy13edRMPe/nWYaAQsMTf2
1fV1rvsVZvpBz3TJHoMq0CfwtjQZfm1JJ/CqTIDH5/C3Khxjpol+JjZhgTOdrCZN
Hhn7TER7xJsfubnBazBtmX8ZEVjmCRHS0/PdejD3bF5gezIB06ei7hOzuOJ09KRX
r4gmnag7ailbdsPma50uzzsgkGnSsYM5sibHl+8dX3pdvNlMIxPPSRSuxr3vTmA9
hkzkjjtgtKcnVy1Rg1Q5ykh2KfV0dKPb/cZKO5kZqGx5y74vl2sR5MF7S+8F8+aS
nfvYEsj94e5oz7dUFKtLJcayWpMNo3cmYTNJ76P6xZyER25HYI7IStj+rTTPeC7s
B6CD1oecjTYHYmWq0FeDI1ehASEvjQrJGb4o1j5QgeMizuBZrNM2UHOLAomO6At5
RQ2uVY5wrUNCI5VDfLGvUcJ8d1Y1UcGE/fuDrg6o2zmXwBuckA85cxTNrUl0AikA
TJFtnhvloIpOzQQ9wXPWGgl85OE7UZspIIkUSHhY384AIDZ/rgxj4jP9Nm/kEqbA
7bClWQ1AHpmO8EqEYMGM9iY9AcklndwxnOpq0+M73XLxr8kV6cCcenLRc0rTsrRS
vOqZ433GRBbyClD4UuW34AFuTL4sdoXHPF/hFk6mw16vp6/Z+hRIFZr/7TP+ucUb
02RwbAuk7McpjGguFOFifL9YRJW7r8DGdKyk+GpYhjXJ5A4scjeZiQEfov/SNaYG
0uSNtWVwIdInkeofvrlH3ktAiGm+hTNXYIscU7lyPsA4zWUW9rxDtfpK4ESVeNm9
xd5P5Xv925wWW0LeAan1XwRsEopFx8HtrBij1adFkYT2gouX6dsP+V0nvGlvYqf1
wXXKUNVQ68DxnhdTsLPg7ZfvtkGCMjeqA2t2s7KsbDBiuldH7XSBtBNL+XNzWG5c
GA+V2fufsEFcoGPkVklFt4xlZG93ZpNaEuePj9ruJMruHGh1pYWQHS+1jD1Ypkwr
RbrHXNek/WQkrhfR3kPf+J9rqhIQr6xfz9ZEzD4rJxqL6AwrzALr5IowLJow4vB2
tHqRCtm8U9cOviEr6zSuDkifmaUYC8aNoJwXVpcdt3pzxe31pwDe7omOzofvVhrk
DVcGDBoFj8YQejPcHQTOmxZVxMqv6RQ2eAL8xr7wX8ODONhMf9HUe4SzGMGyPCsV
6PgzfNlKzvPyme1xYrL8ViJOE7qQYyI6oRLrEDbSFRBradEVAJUdSgb+rj/oYpI1
da7+KhBXoDVJMKGMm/GHtRpUR5UVKfJT4WqEL8Ioapogzi8HpX5V7l3K+9Su/0QX
CDkRgGo4xlY/qXi5eWiNAgA615vXFgpi6032R6eZIBJctaJ+BY14zm547rpy+kFd
38iAbw9px5be/FXX/Y0G3Qs763zUkg/p3kFd4lOZXb9Ck9ZT3V8VuMJBo7cVKAet
/+Iuml2NQmSq4ndK7gcWXmVABcqCJkFt/YYaglINphIDEOz2pzlQxArBGZoY/IRC
rMen60cd8xhqvvFG74lpQUcVPbepfRYyFQE8aAXjHc2hr1+L1mH65cVaqRNmCgnE
FMzp9tD3isXfxqT++pteO4Xx7Gr8ja7kWEpykkeQN5dts+OPQTHZW0N0WvJT2V2Q
O0tV2Rui4zKhBxwVFuBvzMpa6nozeVX2t8GpCUClewfOZLyHVy00dwf+rVzz1umA
ChDdlRGqpiynKnZhc2WNyq4ZSAMo3bTKq77Vy5tefYaQthtHHn/MtbAqvUHQ0tiM
oxO6b2OXNV+D2L0r9j+t8mhQQooFAWbWqlQVZDFCJn8Ip4hQ1+YzhSLgCEijff9R
AGDpePPFlUvdQ6zIL4Sk7QZFVKhQIXDzO9XKMmYmWKQK2xgvYqYMzcpThMdcGlbe
yo1gR76atvGk7mY4XveeRzg4c6fVJSd4JNu2wZx5MO4dBbo3NRcWsAxxp1yKeNZD
PKeDfX7iYzztncnH9j89Q94dWl3v8NUs5Hn9yBlrEW6zknK+rvlOfbvrS9UBWxNR
jLpvSQ7R7ZoTmDSLMiWpgXQpYApdNnokNlR1w675pSDD0iCzrB0wll46ZEtwVl8E
ndB2Md+RRFqyCNBWRtcKK6s2cvwsRadciLDcNBIg7gVtJOWqieyXK79iwyJQJu8T
AJeSXhpjfDUM0FQwE1QLC4Rujpi9bJ5cfP/J8Jlx+8eWJSl0Bx9ZcutUrAuJjcXy
Uh6vzNU7DluuUVNIYqvWtvi4bWjuABBBw9+4io1ul9qgdyg4aAorFfagRg+pkh/o
eY8/VPZ1VShh+CqJzhX5wWFJeBymSdd6c4kq8GSvIA26Rrz8GQh+xCu7A1Yars7R
ES9qVL+MctfyuizxN/9m4xPk4S5zeic2Esf+1o31jhzRluJ/MyngeAEB8qhkYoBK
Y0LmyqbM93p4D3yoe9XxGkwoeqnl5AnL9JYf2x3wbnAq60qvhXj9F9VLlsmWHO1f
rPRUasrLQHE/WHtN52NVZTEHvuF7MzVIlj0Q3UuC7Xy5LBu8jUppih4ud+Irn4+G
2madNxbK7cNsfPJXj0567LHMipLEPQ14Qh/ggMeYtfL91m3HlUDvw6rRrYYS8O36
0I3P3b1u+Bytyp0nb4hxQaG/Vi7yCutGAI/JnZ3o4WhQNVf5Cu0T79ugqKyRND29
Ob7UsO7CNVGzNEUUb5j0cn9GaHlUplhe96cLYJzS1aCRbvJLd3xQ7r5gnnPpNt+n
zu4mCZ9dFAowmJUjErZwCNhpTw72BE50lqyQbvJhJtCvbVAU0M/g3q3LlmcEKVMR
sLMXzMA917fgYpXEZnw0XB44yUSDElT5nqXrtAlSxoqhL4vBVGHhf8RDPOIcly2k
8P/pUIXMNbtmEcIRmLPfCSx52knbTjPEce7tQrmL9rchjRUeC2VT0ASmhyzGyvpS
qeQ7hecNvw2Pmm0gi0aHFWqb59GWq1osM7dG5Fjb6GtROi2ckwm968ei6AuxJVrR
lfEoTKAG/d+29slzgwmBIA0rovI032ot4atwl/GiTsNCH0OgC2f6P/LYql5EVNn0
WnM86PvsVSqZjGJl7wuu7ReqjDcBUro354bAmq2I4uzJ/GWvRyhhR6vA66u7VrqS
/bnykN9ig51ERAMOWO0kgdpAHFhuz4ZJCA/0jaN2sgeSdabA37KJo0+Jq17QBhhN
NctRgBPOnRNLQZuNWSwiVE4A1LHEzJdvSPYvisc40nrSxd1TVseL3HSQiJ8YxKmr
jMKZ4tQD1Zl4GSInH3EV0AAMs9rqLxQrZDaa5eYMGh0Zhf0sbDk/Ucz7++Gf4+5X
ivVfsASuoViUAlS5xkyr4czwBqZ24c3Uv4YS/4UCBBdGC0yYEUO1SfGKle17AdIB
eqVJTL4MkgW1PxUmDvwk7V2chxBajIuO7jv/w31GsBnkSSQCBIp64DvWJet/hY2M
s4kOh3IVSPuOh5ilLXYdX11KPiNp5/S1DnkBIpy1b5AmALbGsYxckQcruH0nwsZH
c8dtSIb87TbjQq54bzNJeapZ3lyXQOuqUxwKEln4WMdBm7o21tI1egjslNxH44DC
Q6m6kF8UdhS7l2BX/4ZK+r5ngeEvWN/+VXN+/WTyD/xwq244r/DeFNc+SJOaPMQQ
L8qPHL17shvVs9s0+OcbwGwJRuxprdWI5OAsqSrTttW8SCJmTzyCnQHnGOwXFHNd
NdfrBsF0odh2q6u9GJ66DLUICGl+IgGW48uC2KEpEQmG47aObqSkGF+r/k+OyXMu
hC42/JAIB5x/L0tdcxClJKSou3YA144cIqjaY9n06mzySn3eq5/RVB/MIrIHKFLP
JYLt+MD6t+8p1frgJaJsd64Kv6Wi+6reFe67OCpF9c3Ie7++Cn684ZIFpp7Yx1kQ
RFdm3ueLDZhChodzh5/4p4kO46klL5aLV8XGERLVTfAuhH98pPqtii9eVqqP8qZM
mBl4SW9ebU5zHV8QMaPOWysCNDpmLpVgXmP7On6/uuquYzhr4G9qzDkpRERJpWaC
1eq2YG7CGt2JwnYEfgDIr2WJLadDcwSEzNuCS4VrNUzfS2XVN/Hl1hc59UjBSSP2
VPe0Tye/g0dK8Cwl0myYvF/SbTkJSE16ZShiNe1vF4e2HV7QGOTeNJje3AsHmmXm
CGFaByKjUnrGOaLJIUm+sG/pWrw3pmnpYQQaHAhnJYzNkBTX/67krQutTBfmNk0p
kKBWmPlvNSCR/wQ0lFFZb5gHX6JJ8fVXCMcgiuqW9PFu8qYrgZ+Jxpl5z09fV/V2
o9C+cR6XpRKeQsB6osSIRvcB9BlLcZWnicbmQ/N2uNIGbaJa627E8Ob9XA4HOY+u
kJbtuknuFb/tgHB2fipsRcEuHGfOLnUqvvmQP2SJRjgXENKbqFOkao0UyweEPcdM
EGn8OZcZdV57zPtOQQRf10tJv4O8K9dy+LZt05nVbw2BNYS4nk8b149mPiJm5oUD
Q26E93ntylDLREKkXlFYIQ8J7LtDJ3cS68OSsBPpIxEQq//jJI79LzZvIUV8pqgu
nQ8ipN32Pk1FSGddXUvJ6cEqDjRbj3cbZs9+/s5482dpCgMQXWwuxT+ILbS8LLAw
4MhZOzdxJarrXhPeEJY8US+AFfs1ZrwcAYX5fxw1ig6gBebxqTXdz0ig9NUh1hF/
SNZZ1K6mLbOURVfhlBDitTB8iw0HZ35HaR95wcAbPz/wZ+UAHLweW2MC2idkrstj
boTzQDQVRbir06aR/C1VrA4w9VxcrVYTdnYyY/Iu3VrsnVLE+3BU7/B/+SldcnGL
HXfTHbfEIAog7Oj1rtR0EBszxN9x+pUvKjIphkLXM/Y71x9RvzJeb5yDkk4XqgKX
B9FlQGEWQ8Nmc6CIXtPnMo271U0mYY0sJsRM36KPGsp0J1/mUwWj6DLrCunPtNSA
c6d9KCiTLkqrESqtkJN65P1WRDt8jtd3+NvVneg+A2wjPXb65p1NOjuHUCkPNIXO
bQ9aw6ZniwreoC4KOog8faXv9q9ZN9ByChnwqPmYZwXKQeJAjm3fxfXkwidOb3Fo
1WyDkmgKvD32i0Muh3QHqAelbv6owBG2DHVdA9v6Y5wT1KBK4HGjZA/0jTI+DPnt
Z255hgL2LZ5Iez9jJt5UjD3phXJMR8T0imr2QR30zN10avcLJ4hxvzxsEafv1Nz+
v9KKsEwhXOr1o+a/qDVSyqGw90VYx9VWtDPGTtb4hWLYBw7ht7VFwCrNJI581itM
Ll2/Qf+7DXKLI4/5EdfOIc5foQCE0FLiT2TBadCCfsyILvKL+ZYfs75f9f+ZofBY
UbhqsOPot8L6MvmJ3vFjQCcMs9lm7b7ZmSf3FePsG8/5cYkBhTyRWSWHplJ95JHY
Zj+FhaIyvRdO/BiT7LV32WyhcKBs+0LYea0LSgqur4XPuLTLkaCuaw/tM1DhVjOa
XpRlbTKLET3vT1kOtE6pS8KsMw2Mt1I6m/rWu9zqd6qyQeVS+sd6U//mgqa47gXG
YiMR8c18hLEqJ73HJ2TnoWErEtGjVZ+H5VFYGabVImFCCHkKRRMfC6h+nRQkAwBO
H8Q6Xy9zE1vmkq0UXS0nPxHbwRvUyXJkXH/u6vWLMR317G7GTcqpXu1DXj7UJEHu
+jfA1v3QtFuAQWk9WGHEpY/5/bd4gHcMFP+L23bu6w5L9hx3AxNO93x5Q4gi5dEC
ci7LWz2VU2n7JKlR8eVRv0qFv3OiRaGDT35lp6m5v5tqKqNEdErjYKbI6rNbazSO
8v3YsmvwU2PDdg+mdNKe7Q+8ExG9+7bbPiAmlLu2VbDiKQaQqqrPwsbqwkUU1V37
Mt02KIE36v+VUkpoka1jUpsSvbOC2pkD3mK6+n6kjSTzG5ivs1gB7YSWc5NRhWnp
qgoc0JXlFHYS794ri0l4Fgu2Ud4+XkZFCmpsg1mKtCZlKdP9Ldz9lAEhXDdQHiqO
WuDj6lGDsRKHxD70LfeKiFMzeR0WmeXjet9r8l+82ypdFrQ1XOulwDeOTCfvYZVR
afyllYzRjHqaCXGnjwL86+puKQX6rem4fkvhkEnsZAWiVMK2huMg7B6EdjF9xaqe
HafiOHG/D/IDvTZcHtDwPFszNV6RA8r9LVpimpvffygqmnATGs/pbEnu+r2ak1xN
+mZB18M+Pdo4THw62+Tzje/+qpUlv/ixcUMfjNc9xpQbhoKvmnDBrmx8XjO2wSf5
LmY+E4Vba+r5ARl6X85xQvGdXoE7z0/+DgP4z+cgY4zdrdwSD3QrFZR6e80jrX4M
VVOrkHZQIwoEHRuSWQBcF15Es9Y6KesSl4bfqsEOGWKc+zlWoWyAUceZRnfR/GGT
a6tMBfPig5zoRWeyIDxz0Fsu9q8QerxEkx/22++gJLC5wxB6EDneZ4CT/GcqOqeo
AItpTmSwM90KMWNfFQJ/ebdkm7s7mhLCDHgIHiOaV3UmCbMhUfgdjBVgbiYgf30O
/JZxTWHB10TgG3VMr/qITaGS2CKwc6fyhwxSVTPHVdv9X7tpWlV7rLNMljmhx60Z
yAndWSmaYCS6vgSD25dhwhhBX7hv++XWUupDG6AJG0SlxRPJ50sKcIgc6YXOHpv2
GFBDLaLrJcFKDt6CQo4XSp760daxQuWfm+c8RUmxDqhmFdkhdT4gcBx8pSbO5GXc
0Zkvadb2LBAo2RkAvDG1ny7i1RGI5yetNvaNlSuQZw4Mn1xfdJFGOtCBXAgFhfDl
1MJPJQVjnmwNR+uDBJgBTeQUaO4am70liyJJCzD1QKk/vvtj7N4VIYlXaElv9Y3+
haiTIrWtVej3hoyOa1aYgqX0HdZqvkXdd5XYyQTmFovUk4BmMMxGmN96k5y7VtOr
ZqP6XMRNZPWKyThTllJD3fJ2h7a1dq/Yh0qe4hh5SYVB5g7u5YcrDKDdJG3RHFvv
CcswcGoBuJmumPI98ikJ0HbgdWptSNeRvP/C/y47dDGSoKI00ori05e4CKkcHZWC
tleD+o7YCgSsXy0bU76VAWzvs3tjXcSxD4Ybnj8H6DyeWgLB69G7TnLWEpsdSiNe
UwDLgaS/3ErjPiEaPF70dqRFYWJE8l6oViRRW65xibMrqm2gBo1rx1sfVTG3APqs
/Zq5TcXnW/Obh4QekJagaoz6JBrRc+9oWXYPW/ltfXJYxhBa5IY3Z7C4xkCZ8Kcl
XGdSnfFC9Th6qG6jf0KzzkdHpWfM2oKm37bXnXiuQS0KdVVqZOdka6VFp9fVxQu9
H8LLJcCfmmXO5ZySIbFzAHx8bfp6eP1n9EavzQGt6e9a3ljHmvbnArwshrXT4ros
SzzR4lLz8S/QNZXFD47AtX6WHbiI5onXMwZg5GyzxajjUBiyrI3dda49T01JZ0xj
Dtzrauul5CFfwm6DFBvNY6MFUAJ/uP5mMkaHTDVp51QpgZUf5GBhoIsOxA/2PXlP
XPRqYRwoxeni1Kvw0sBK3Eynn/K0qcQbeYCkAskSrKZr0n1oDHPsrz/DLfPuPWzE
mnNadf0Y4JdjSbrq8ucAQFGsoYvcqZEGLfqgjFjFgc3sdT9jzgxOp7KWLzWY5o1l
1lVwF2It4n/zkpMrnYnexwVwnAzrl+tkX0a2L8w4bkuDSDq8qbUijzX9KO+LcMtu
0mhnbGebul1OCiu/GZSpfdSqkOxE2H30W/RM2rCmIuxIcrDd2JONJJU2oWmDyjgL
ZM55dBsHzDC+gIyxratCL1VjNV5MVkNDisT+PphvWRqL9r8mKi+zgrNNHmdTfSHW
lKs+Nm8kzYrIXz9wPs+F73476LtWsF3WdAz0dSkVMVYSNVrpnw3lnbptHySWtUTs
9j7DZW6fFxD/xvAO8lRfAnVd3aW9gW5Drl3OZPmKV6DLcK/7ZfcijmyP+f7FiTlH
Nt5cXeuQ/mkPW22pZYLcXztTR6oGmXBopRHOImRU1SK7DqH0/cNmJUpyuoshK7yM
f2PAtavqvb0885+3OsruK+Ni/ICXN5kCbt9va0r14N7gNTnoWtdD1s7kpqOe9wsb
i1ax8ToqKoB+UNsTYlGJkH8S7m/3hGIajuV3IRGXfjTG5gL046EUq98P3iQI0FFg
X1co0MJd5byqpLp8ldvHwmLNxYfNEeoObjYWfo17PZv27YIJ3fa4pTfBi3V1Qaru
RlpcFuFjmkkwXn7q5+52W6DODhNjUsnTbfTIvDAEhy1M+3KBM+4ltuLtAzXgAW6j
f+pW7uc56xT7IbuFhZK/6JxzArKDrnAkk/xLSAhNIZ1E1TqLXwsWyrJpSGNPFb8i
MF98XZyoD2iMRPt3wPHW0mEcSpc9N00zQnUDOwyBU96DNut4YmUQrnnmCn32Exmu
noSLfhwIhep5IAwDfifmcZFApuIlEYoMN+c+Y0IuHuXDS2j7X9HTY33aWjFEoCAW
5nhXNjXO8wjz5O89HeHVDDuuA2sJYBFLXuOqT96i83G+fnr35QdbbEs5FnQt90ad
+2bR4k/A4Mkv7TOw2lmKlvLh3Nqp7Kftwslwt4ZdzuWZHJf9Nzr8Z/iZRO/tLvRw
FDHNJcporoS8bQvQrrUI/YY+0ODpV/NXfL8D8TNF/n/F2Ri6DR2C56vR98ZF2YIv
nanMKOMjqQilqcSwmDsmFAfMa/UHijnPY+V6W+RmzFQNZJk0gEt+VYDN5/5BfHM8
lFKLG32fU1QODu+BwSmlEOUW9ykl72WFPZ3enrwdc+OMycPISqy65MBrNVwJFo5B
Ax3nDKaVa8oMHxsOF77K2AfKdHSmhb6Xsw4Z1XqTv3QwzG6i1d6b9egG7N2c6cKk
CozTv5NiOnKyT+dcy2DONQkHPii3tt5+U+pIucq38rtL5FfJPkHO4P4mb5YrEc9Y
jTEI2SEBZQzZ138NV+J64rHmgJySHFjSOh8Zb5DeUzzXrUDetC3BSJUdrLPElEFJ
0kKVhdRVIWzyi2P5yFlj2HTV4Wn6YdnQ/MbW8TtvUfphorzAT0vJsUNlgcifaoNL
YfINpLYE9aD4LDFEJI+n+fGE//l7AP6XUlPCkTSo2opgQ5i8UHjxBmXAG5LYsoqI
7JgWmwfUFuNV3wSG/nNIqYYpwWV5p3BezVwcDADQ6znvJ9pHLZ+HXBkLjmN7RSwp
IBt1OQ8hneAPczYoO5tzryf6JKek8K59jiL9jIem3Y4DsR2VT6pBl8NcqMnTXv2U
HvnV8VbV7bajjOZoQcYL7z/ODkwvRuBRGhvqRDrASV2bLPrvpTJmhi1/KYADk9Br
c67TzZ3dFuEbhfbDRj2PWW0JMfVnh9IlWgC8h8cU4+6tyFl2yZGmXd9d6qizNxyL
PFtkBjcnjn6RXU1Rv/c13AmoqCDHX86wKOk/F9Ov05HQTbNBnuaCqgsb4HnL8PTO
eRYXlybSjRZ2BX2QQ43R1WnzlRiDHC7HMoG8xEYIRubLkXrlwHumjd0G32PAV9s5
04zmVdemjSxwh+DKTnovEqOuoW8SxfMpBrHbn6UeQgBHdC8Tr+NZzCwMi4WMcNNy
wEukCgm/KU9N8ZjZYOt96hlQjr6xW60JowNp4nqvInd7leJJITMt/3vKyDYYzJm4
UaLlPUXVWsjIebWC6SQ0FhnRyoDDVhlLmvOBgQ6BgxoFZVUjmN+LKznubwHLuZ+6
oeXfRT/26P2B0TCvR8Zvsudprr2v62+L95ocphnFQDl94eDBRR0s4iujQeLDT6Uo
0d4f0floo/EfibSHF1tniwXGasB6asL1oAlxvQhpVGxnfEC3VHSadQePFKqNSeFI
Gi44E/kRxK+ZqvXVlzx04uoeAKI1tTYWhzrVNkEnQpWCltimVfqmaK8qDgOufojY
Wm7L8QsiXadhH38G8/Ml8xI3+m9gXfHqazKsjhdQ/bikorvSb7U55oo5s2hJd0RF
5ueacP4LGhOvYHiRaC/tT2ppMLv+R6fRW1/gSgWEiDT/vwr7sO0cdRbX6bJ+Q9bb
2JDMrmc8OxXijrBWHYPYe2hF2gfUTlgN2TT+wsy4BJmAJoasFrbUIK0yoOn60gQ+
G2MNJGdS1nrtlYXn7UpjlvxxgjbpEt+vZ2HlgM4NYcnE3D1A5ClHxmflJf+gOzIX
z0fXOr58E01cNLhVi4ASZYSNOu1JVTZcWsATb8JiZNsK6yZUPiUtOuqGKsfcNji0
eiGrZ0wfzuIIqBClQq6sfS++5C1sw7w3RU7V4TNvRE9Kpjpo+x6dmhbALLGvEas0
yFazDHOqlkpF+XdDdFY3z/FdElKUd2R3GcX3RtpJUgmnbk6wiKcj8Ky22bDW4dW5
y1ThzVIUmZfen0rZzbDg/oZzCezEWecFfV4bEeW4qzDmhmBS7Hi/xjDk3kHazi+S
M+REG3v8ip6Niav1LbSj/c4wlspmNlGejUT8lVNISdd4sr6V3ZanCwpYYnm460cZ
8T0COJTuWc0EeYoLCDgDdQyzR7GsnPM3mDGckMaKvnyzdxi3ZyiViZTVq+c1HvBo
LrxVQdOmCLfxROtp4FNmzY+co0/AXpjgj0eo0hqa/xnKWYTyY2CTy5SjXuU/GqUW
QbbaQ0clL6Grjds6DL7RjLBSrL6KfgbI0WNkaCm8m58BKx/bhbR/pPYTAV8M5jah
wBRsqMkKYpa/nO3OtkJhU0P0nQuhOD883xrwIBizaSNwV7SnytThZe5LZUPdDVhp
+yBJKGEHtctTJqRxgykM9aBFY+KT791GENMRh+r8wK0VoR5l1hyNmHsPwvnMyOvd
E+2pPXGgr1x1lj4OWBJWPQjix9rVR5MJ2rFrsbVPzxyRUBfs+kpRU5bLe709YU+y
mqoOjrwus9UnQCCKF4naFofVP9ie0NXHWOiiiL+VH/TWwfN2eL8Py1pz+wPCFj0Z
IiNAe2uHWXSiH+nOf596AfG+VoGpkzSOPIM43xb3qyEKlWVD83QC4fEMRclm10Bb
mpJ9yzmHB+s81ilTO/RLBgvz/bRJh0BcnRHlnm1wfzHV2x1EI9pwZByY5hBdsc9H
1ZsM4IDl6YpB54+m7P2LjA113oruIzZbhv4oJWM1x0ldboX444FuYvhB1+56sJvx
eLSxiX2lQoFAF5OaWQBEz/PHvZkceTO4EZs/I8Q3IPZGn74NU3o2ziiSntHN5M74
TN+9HSSCXsjPxJlkNCVASUS0JLRTjBaQfkNQmuGZG9AByD5GiieT0D5GslTo/9a0
IpsqWcay87oIjHDh6kRdypKJ1J8lJ8g+3A/evpPmVYyXZPW1pEiIENQjCkrHXTHi
AvxMJfrSsGfpj47Zfm8KpR2RtjzJwxHzbrlbR0KeHTAzVoAjqwvVqfRMjKd6MQxW
IS3FMSuUwZbhGJWnkNi9b8CPQ0MBNn83m/e1d7JgU6FxUKE4f52QDg4Q8x9qfY0B
KN0seLFVBjEipBs5XfEg/KZe92B0TarDfF3Ki2YPYzHk0vD8ph3btrA98pKPfUUB
RD2nRrDZFAI0WQEP9hHV2kna8PW6ddnmWN+WbIgKaIXHDpocztFR3nj8fxwzTZ6I
jaoye4IaWDMkp368Dhar6iOMk/nMkcB/G5CcDLt3r0GnkCj2gtTL5IpEdQuT1Ma1
/osw7jcYocBIUgc4Gqm768M1gkKliRtRlicxz9dOhGSMxm6iu1jsKf5A3EzjUzKY
Z2oOKDo7hHn3L3etp3aAWoBKIifbTlRnCpNOwoYgOKTJXbtxTV4Q+phleQcAjR1s
tZ/3nYKAjDdvX9BhbStmgLdXJPXeMDGVsy5rpzqb5OPRAgHO8Jbeqj/nEJUZB+39
s+PZCgtlkt18pYbuCLVwKpAKk2VVJXbcLnlleiXABrlsWkaLG4cdNb4HZZI34dzP
pEgnma+b+ezigfU3SNAYi88PB7xSMi/C2curGkTeBJNNEADlzWOVfSlZWcSzMXc1
4ikp2lDhgJ/46UEVcvMV6sx34xpV3UET8WoUC8mZnjX69QZnpF0mdIFWtl9IhlQ2
YT45eXNElRbqPvcTJOMdUOxAQtMuuZbNektJwBTeu3l1Hy2igJU5J2UiT/VvOlNF
XAD1Q46Bqumw742sAJCmG/vqbJaCzrCp0IQaz+lGe3uNk+IqU1fxIwEFOe1wu5wR
CMITftPxe7TmyNf3RhqnqZ/KCk59AjIYRqobnyV8+f7HgzET3nUj2sDJfqjtGf/v
hXlAve1YVrIVrhUnN2ATkkFedeKeZKFNkhVzAgKSInprsOqPex0tYM+shQd+m6fu
b5pR3U5WaXu2Akb/JY2f9fyTm40YefvQP7KypbB5G6dzx5wYe6O+DL/SYYHo0l/h
2AOBmSPnSmzewAedIbdY3S10UQHtp9oVuXyfl04Lk8OuU6hg+5PvhcPcAog3bJSv
kZl7Ef9o/zohwMeLcpwK2LTQl6WgXAv3O3oqBrsGTaS9XvJHuWuzSJ+mTveR3RjE
SVQ3fwBNuWEDJFyyjwJQufwaCDuxZ3/jdCEmViN9040F801mlUdlakjSwx/O8qTN
5tn/LtQfRgeRKdsM1jeiI2U+pYP1B2YkcPrx4J9VzWUw/6QoHEERs9oYsDQUAuRx
hZ6dg5YYScM7D7L91McrnV+WJBxq/O1Fw+oHmS6kR3T0qalyDzXPQbA8Zb9WQj7y
tpFBq7n5VbEpDD465uI1IwHhGdiHUYncHysmPSSbMtTytVk7kEvdATZM2VeazhNE
yzU2M7dKpnzMdupDP9BAq5ZkJf1YeKHhdmDyK08KSQiZgaNIkn7Jbo++9utGxByd
Wwrcps5TNMU6yIf2llk/1g==
`protect END_PROTECTED
