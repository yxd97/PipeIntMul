`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kn9EwoiicYGPMGXyTpHMOrc3H57VICXldRchDKG2VYgh4Np68YP4Az9Jl19tWolU
1QdG343x3fZYu/jCUv5A8bAQ8KV2b2IjwJbr8561/8D2WkPevduKDOzwA5dTg0SC
62c0o/eqY+IyLobrU7ROGWsN5YAuxxfoCFtlMpC/zaYAsPFYquojpedzd3/Rjtxw
QaXuV5xQAs/hBdSVP8VdnhZwTKyH2dTAUOgRIJZTblHhbgmGYhnn0JHBZLlkVeg1
hoURXDjqGpZYatokV9Sz3oNlKONVfj08NK9xj4XxCLmZqcUdOTsFkcFy6Y1VRX0X
ujIhEVFrTlVrXcIEZ7A+1p6Y7odV4tY/BI1+4MadymxFraXqo90CJJl4j92KT+2N
fZx4lmSut21fjxAa1Pmc3jRtqLxIs6aADMkR5qt5V9hMC5ZtzLKcONV29aUHJxwT
DiatCCEEm7JM9S8+kPZ6eA==
`protect END_PROTECTED
