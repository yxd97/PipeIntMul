`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2zkKzmq8BQgTGNSrDgzd5ph8YUt/qoVSSVA/I2grULP2NqKuZF2w/b8Wg0TKyt5
A0QD25HCzmOpz2luPkeEMVAOJJanuRbltKRRtBXqPYnq91CccLdKKBoe1QhsnQK/
+MxB4duvfEx9My9ls/JIQGbF/baIMWAHqZaAyF8DUWc85KeIqFo7G7HGfOu5mEoX
9q6SdD6RK7JGRp499qT2TvHq1g7h8SpmczOXkytmGZKR/NAiocQNt1Ql6pGYaJOo
I5tkRQbylSpH+WmdVhWfpg==
`protect END_PROTECTED
