`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVtF4/Elc+3he98aJdB9eBrY7FoB6nUYcayHghZXGO2+fMzkVXVHIKzkQgfVvly5
AtafA/WepmHCiSWiNyad3I1D/hXTkO7wMIyzUDsVnSfNp4YHWPUcb5TrHcSmxbL4
Jf1mWGOgqZ8RKENmBoP7HGGGumzRvRc6lOXg5y3ecrY+Jp32e5Lv9x/6udirn3iP
mFSs56Xh1jL5Xx84f1vogltU6Omxlsio0DHCXGhsMcrcUCxrlhWvDqyDUgX8J06e
XDOsTaJnT+4s+76m7ok3gfP/fiGv01+E02wmNGslvJTVU0y+EQ/mH7ZLaQW+ajrN
OQIJ613DX0HoaM9p32pIk4C1l975XlxRw6ZFpksSGQq3Flk+xDFqHipt60ek+lH/
sSZerPO/aswCUgC5MBTy3B/tZgjwc7uvTBszpIB4JBda4EagZJPs923NsC465Ep6
Nu+WOBaFvSnjiaZGTX7u/WId+MH85Y/wepgcwhfp+3suBzJkYxlkBpZ/UWnwLWUZ
`protect END_PROTECTED
