`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nsMBCu09azN8FAPpQ3MZKcv3U7PlOdE/XXf5wOhrPuZOMEd4J2YfmyUo4f7Exdxz
FvQZtoFV1iFyW8h01Z+BszNK/F4vEU0mB7XbNJobm/DsSwWUeVYpRTp35u3YxkML
AG0ueQvlDgRLyHT+P6IPAv74+Xt5/jFOvKeoibdYDS3LH6KQmMsd44/T4omrII0o
A/7L2VZsHhSwAMP08U5F8ToZ/CzijGKUeqmc82xCY/Hdd0gL5rjZptrUtS3lGqhv
0uvgxTnxe4MlFNeZNjBonGRcDuF1Rkekxtzo0hh+gHb6Ph5nL+2WqlE46G19RXiM
SZI17CC7xtYETr7TxJQb8p+4tOpoNmSeMIXdF9MXwY+V2JIaS4EehMhF4eBUT/lR
qmAfg9t5yknh1vJHNhyikyY5UIMFZGCJZw+Nf832UbjfmRlyicjf4oJXZ1gLzrGQ
VvIY+RFqcUUZPq2cUdII/eSJxN9W+DlbT4nT+mXtTh4AOh8DnUyEG6zWt9bqXcxc
CG8+WGbdwPq1svfHEFabXpR6lm0MqEgWdKn4fIgGbuJfD4lVCfpt7DnuWw5kOw2p
Es17XTNkIuBRRmku3ZyRcavR7/nh8ZM4CDi8Zg4N997WmKKLrGHK+ed5BirgrytP
MwcQqVQhASTT2nIBcu5G2wlEC3sl/0DmWtTOHl+AdWJ2zqecqxIpzRbUCUpHigUg
nWp+qBNwLlyMZBjNTaH9J3k3amCkZY7VYw2sTL8117KzWB0XjXll9dtIEITfiius
cyupiCY0+ksurtB29jDQnd2I9KWwIARDHrW95AyEkwy4OdzqhdXYfZouFhHYm/cQ
dDiSf+bA+BhyjTo8toAZeA==
`protect END_PROTECTED
