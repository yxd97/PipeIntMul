`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6VLH8/oIEXxY4QiIKTPgldKefRj/+6Rip2BzWXRhOL5axlIb9jgLJ+Mhf6xoZxJ0
XRmpHTxVYgaCPT2cqRdT8efUx/ONtPrHeSVjgo5X6JL9hCrH65xC9ZnSLP9Qdetw
ck/JuNaZQOubVGWJNp7c8JaMP11nwRD9xD/1PUFhFKAVNUDnicmVuM1bwY1ZCXpl
QuzkqkBRNIu/GDk7xU8p1UAEoyHZAqqppzPktdtEGJLmB5vzOlayIhfJ/G7tUJ2z
bOGehkWtpJjDzTqwU17x9O5jChHYBtkkjHaEg/BF8JnjiCGk0j5GlCz8QlxHHzgn
inEiwvY2fZj71s6UTCVQWZc9OL0nB25un5jJ9fUK5/oCjIlJnU7IMwHOSOn9SGYa
eGDTdDumjCmJdvBbUiSJC/mnarUA9GBcNZScKusvoOGaukEIugaoflilHauGmXtX
DygMO74LwR6Y8O9Qptv9lcgBtYWG0tqXUZ6D2yGHCHdY0S9C1jDiOWbqN3pLa0gv
3wJ/+W9X6ruFABouukP9QJSLi3fm9wKvqVP2C5auZFTAKQ2RNQ5u36Lf9wz1FW4W
xb5Q+TO2gB8/V4SOUnO4VtbJcTo4En5fKjJn4bQDEO4hfxVN1hfiGk3B9XY75SMI
1p7QKLTR9ihO/y0wT4QCUQ==
`protect END_PROTECTED
