`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
raOk2TcaoydRImTk2vjXoF2rAFHpFVeQ/LNGx8du90W/WMWy1+eGwsPA/Z+DILSv
SsUbnzj+jjTYLZqT3UGE9LpsVG/sr6F8GomNnEAImaqQR2lnECEQDPGMJgGsvNXv
3odX1BJdu/6XMDhFAQGy8ESLRqxxvaRbd+HnEjpGwH5ovTX4rrKXaKV9ZrYeFJNH
qHWPY/EXhN+nBAHhpStWhr5QKeQFupxAOBRwRXUyq8SJQNRY0LH6LP9UumcieawG
ETGDJ6u09xmYY5d4FNCnbG71h2HfSianX3wNCBRx74rIoCtEfOY+HOVYw8P7/SXB
JwwzzFdDaMNZzEVJG74HOHALWdAcZMlSSCSZtfoDHuSpjPGEIZMJH9uZxrA604tX
fdPlKmaywsFY2ncpWgRQMuonE6biwrNossFvYbKI0d+9QkOGUihT4WhSlFzVOXT7
BiRifxuBBJbR0kkjkqYcICZWhzj6pHsOl6gtx2kMGYSZUlvOhzx77La/xdcxr99b
a25nenaIRl45wVfmoYxYhXmgYG7P69QbKYTBnyvRe/l/xNTKyjN2hv30AUH+wH28
zXGFVu1/z9Fgor4AqSmQlCGLTzYjSdzE5ebVqO0Zhtg2YM3C9aiMY/LVPal18I9R
dhpjURBSYkxdUAfVelO0iw==
`protect END_PROTECTED
