`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/zloLsX4YV7yUNqsGPGKjhhc0pYtOK5X2JMjH6QW0hdXFD71ghIGY0oLnaGgsm2
uRm7GtgiKR0mtL4/GH+104gYLHLpwk8Zj4/c3Sm+EAY57bk1eiJzPwklCNTejbJQ
YsWD9Et4YV5SttbWgNulDCaXxH/pqnBDv3Pb5UaX4huZnK1a8hi/WR59EqCgO2S7
iEvaR8xjwD1R5aJsnWfAIaL91177a8cR09KxUaGpiiH3QvjkkdLLgWQBcXKWacMJ
f77V0GAfC7VJA8Zw8AogvNBxby8nnX2jkZgDsDP/rEMauhIe1LHb1KF4gS/yr01i
4EWSa9fffXXf9UFLCaQXQJExWwiR5o2/w8tdEZX5nC9BvZ0RTeiC1TZs5not1Cl+
LStFdrdXX5cAU6HlTu1Rypfc+Qtj2gwLMfrjzl/s2Pxr+Ie5LaiXiOzpMSQ52tbK
waJMzJWfFefWjfK3Vdcd7XOn+MPygay269C4MjYFj/Yy4zpLwZ/ET9Z+o3vfo1kW
fzqq5uNbUq8/MnLzJsKhEajGjMgXU52Y6uJk0bjLkFLbv4auwljVPR5OcbIK8oSC
NkySpCxkBa0qI7PpQKR1TpGSltf6gMaIJJYcR2CEB27Q6MNCSsjf0lPX4ufxKB2H
drTNQXvn/yujNdV6pY0QAYg2trB4SznAeqiUTvP6OT8bbhRu1B+pX+SgMtqfIqAP
tbMsOHiPR0+jYpjhEojuAAUOTXhv8R9pTILhKNPV95Z0s23c4MOaMsrsVPY2hT5Q
yoeBbmV83/iyp1eVrwjyJdJISbs9wwBh3B3cr72F0W8Xkvql2pMXwxR5K93t0t3m
9lqtKalcfPTepe/6rrdlMxkLKEa2YX1cSXV5PLkw2bTARF9g1TzDyZ8DmqqBGHYc
LyAxi5rlr1zUusA5plhSU3QHTBP8123Lv876JmXdqFE1O17tydtp6MOkI/l1Tke5
lNlcdOwt+oT1DUlNUQbl/YlHGEejtqIhIxVSODFeadZW3zNUkfB4bYSHR7fCCxg2
I297Cxjx8D0J824BzKwiBoP7OvHcpcmZ2j6B3qfK3dOXEmJ7strF2iXBwLh/0yaR
iqV+w3tQdIWRqQAo+OQKhQ==
`protect END_PROTECTED
