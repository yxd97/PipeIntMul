`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nC4RDby4fouedT58OkLI1l1GbL51ZUpPY/UC4Pp/a2BOIKIsTOgyksaYUj397eqh
BwRgp2dflR2b66ynyNZFScZ51Ze9c+SRjzycmDAjelO4nLd4cYAE2+WOsMtlKrUj
8d47fUA4F4i+Jmh9oMEAjg7W3fQiBTnn8DC7K5B+a4bGjFKp8sSJ9khq+OXkkmng
4ZyK3+VI2uFA8hArVG8IE749sU0EImjgKS1q/8y7dbvCDbXvQemqD0pcs7GHvj3k
8nL3A7znf4liA2U2oPgHLkGTcgqtJeEP56gJs41P3sLLUjr5HMeKwCH89Dlixtor
n2Lft+FJQakYe1kU7YSgQN8HjdT5po3Opk4lM5ESYI/YwBbqELEG3WU54TStp6OT
N1oIwDP3KyCWPuQswnTTgW5EoaS3oFPYoN9GOMFXk9EzvFP/bJtMadR7alqrTJEq
cMRMNuVemCub/ubq0W/F0ltli0AjJ72IOkUT0agLG7HTLrBEYcQnAgMHayOp6nrS
lcTB8acnVjEksa8qy0R5JxAKF+Bfqtj802qZS+hpm2Rv+m+OoKm1ts4B49/OsFrG
NX48zcKtQrf/31iMB6r0UMNQQYdOApd1MOqK9//52ftGMNjtzr33XGbRWJ4fENQj
0ATXq0OESTiJ565010E4KsbD55DdwbmeycttkHPuaYqGB16FOHOVwux9XRnsOjvL
j/y8+q+imwXSiGm4HGyCNsPFWUn2sznBkktJ+ARBUIqHK4mLUPWUmbz+psCW7VAd
c98n9aL57Sc7MTwvzkFgb4JlR4x1sZWtgThTWF0/Tcr+oAhy9BNOUKZxF2BP/BwA
Oka14iG/Ed+XiPYa+LB5yUh11e+TAUlpwnfuByGeC7tuyng+kRR91gpp1oEZE8gr
Pu5ipVueYMeI7ZIAm2iIkIWTok5AX0bD+JFMsYU0Fhp651SbDq8DSBwQxJTyO+sQ
JDpZ8W8Wb/XcxdNhuEQu+eKrpayQPoqsVGTyBrwgd3ZtT3DwdvBic7gdaFcb98yG
ovnZW+Kd+DzohgiG7vCiLBV8XGmIzWFFRk1LqcsbYkMysut5bbbaP4BBW0/3DWU1
pcEAw29S1q2MN0CsezbYN5h3iQZ9cl8XCvMXFfMnNWLHgyGJ6HRmE43G1/jkgRwg
6i/SGAdWht/axjCdZu6ltPOOQtrpXWed/ilqdlwNINkX8sAeTzqqOu0u4fF5owQt
/Z20u03mI80RL0N4n1mw6rsMzXU0KICcPllsdgEgjdXIwT3Q4E5JeSNdu2EnuvY3
o8BLGsF5C2TQJj3lO5W3bmHY5ZgPRv5f2WLo6ltgN3MGY8Z4MyrJI05zG8+nTfJ/
GK08VL9xG+nhtAfD7RtZ9/PDCHETV8OfSsB/wf75zyfKHs1b/ZUmln30zqA8qAqt
y7VVMzwycVoDoiy2Dx3bPQgc+LKLOs6k/do9/SwNGOo/r8MlNOkwz7jGnvz0k4ej
6lHVglSFIX+mpZZeZeaHdhcnuQ4OdpflzOUwawMdgQuxfEkPY3q6Y/ATUyM6Jihw
auRbQH6enirQA2y4cCCg1KWMssKaJz4ZFR/B3L2DLmWJX1jVvtgA5uWZxGwmPsWC
o1MF9MJaoRSvGT2Fe3DD29MncHVqvfauO2BJODXC6Ex631uyW/U193hA19ETEOoU
5w1i/o4xlJREX9S8niUQj/5bA1BiIt3o6AQNnnLaJDRBTMmxVjfEQKA5bjlf4iXq
e8aALQ6NxoFsxb9qeK3NZuHtsK4/jTwoVjGalWpNI6AArPBg+hFIqON+HJ+ldEzb
QM21oz/7dLCIlysQAjOPsf+s7P+wrlGYIiB25saAuV4xdQjMkE2oCDWHiaYOy/yj
AvnHaN06U+hKHH/C2KezQIcjBD5Cd3oDgfqgDhDmGdpwEqzpTslr/jCersZPvQ8k
xEzHgmp6UKTSiNcw4qkYKp01W7sZYrRUfHsZkvxtmh9sqOgUBn7RZKbIuXfNQxMK
PNAPH2qQaEqX+OdGgDn4MojHIX7nzN5TxiZPyVTfRl5wjHNB+OJRBB2/xTGadn85
RheUN7UWi2iCHLrP84/Ttz9b4i9A/D9NSbzgBWTrLUf4/z6NT9zno1hWeSJE79GI
Zo8Kpkn7RYv6D7Js5v4GJGHrK3lNLCTE6X+fTh83NSt8CR9sumH7QV5j+jfIk1V7
KdI4aBNV4wyu6Vj2B6/rFKRIJZr7/OmCaKisxNKmrPXeiLiIfHpA3OzOkMvVf1r5
MrtVzSoRKiqtls66K4pHxqfeXtGoO1MskYd/4r/vGisvN9qq6QFPVN7Sy82MVht9
SbTTu12xDDDR8WBIcYkcW7BEVkEijM0b7Gczo1z9a/sjorkgIoAsVl4LE24Ce7ja
y23EvAlW91/nygYuluciZaj4qKPA9/3+KMjOi3baJX7amozcFzkskSFhZHY7yWLr
1ZSn79LfQteI3i+XL7PmHjnfqZyWQhKZ07tVFCeBSy6w9kfduwQy7xrcFvx6heOu
gsDUJK5eCVmbAvkVhI0kuvipVpPjuf0L4me228dnderojJ4FtJORrKi0LicGZv5G
aLFX5OCh42gKgqwfZP3EPWLSSFoMI2hG+A7OjwyQbO4b4PDjWbThQMD6PnqJ1nnM
rzak3wR6CTDvfbX/KGToI8TSJSo0xhOeWhifAQOgaLF03aqY2i9CF0hoxaYd7WCh
A2CjJnUsp0Zzi2MYY2pRs8S9y4+4w3Ykahcz4FulpuySquQmNy5/n/oefK9mMdvk
d404ABjxTaM76WSdJag64sWXbapzChCUF3YYPGbG5xi1OqBoeq3jXYXTsH7CzlJN
dpJT57OuOg5kCQvcCGEshLJIeYfjrLg8r9zM7ZL+ItTQ4UrAycgcI2xhVC4PwvSd
JKiaYKvSTnzZv/xLi5s1CjKQg+LAyNP/y9/arZae7n+ulcaMVvXyPUROrudU799b
L/LPhn3/g5GPEwgkLI9L6K2CEZ7oCDYqigGhf5bLurI1HO2/RGJlCyfMcxXAcQAB
0g4/0/7Oo10unYJZF3G8ZNrv1IVAJz/9knsmnsoMIDytdBx0aooSXU8UFaZlDOp0
RNiI9kiVPXqNya8fYLY+wG9CAVCNtp+tfF8jcb3DSvzQjfpeEKTlhUGBv1cLCyys
sdKQv/Ax0UdwGRSxlMbCpEDjMcha/w1IJ44Ijrg3Luitng5cfjflasqqnET4AbmO
P1rO6/VIg4jAVVVngfk1peAyBlWv/U/82+Zqit26ihbeSXORem2BZNkXFH3nAmx8
r7XQMZkTtzINVNBmiBtSuUQCa7VXlW6DBA23KTiWdybJbe9FO0Ag+DaekoZDUnkj
xkxK6U/DZheXiaiL4mk5w9/Cz8sR6AQiX6Vy/sHVwR2tEt9RAhPefAKy5VH5Vt+X
M/Lje03BDw5PO6EOyE+fn0Lbm5N7PFAe1sCUnLtnMMbPdAj3OOFf+yX3etDVzvYq
ogQonGH9yhdMnNsngXaX9WfQIs5Yw88f1aBdGsBRWVVKaCdlPnsFjcEqGkhhX80b
3yvR9Ioj0bH5TgyLz3+giPkOD7XMNep+suYnkgtc7hzOhMypC3CfAfkxr+G04VXz
tSE4Q7CRMzMe2OAdpK5GK+6bKmAWN8vf1Jj9CERMMx0AA+kY6f/DVa93sfeNjj9l
d3C3sBMWtZIdxgSpFgG2F8PeDNS1prblXl0QcW7rNq5X3lBJzn5ePdBO84WQ8cGO
GIqrtGziU0VvsUFYd9/lbxPN4q0On4sqGnUvcTVAbwsmQDmU8CfCTkFn6u8O4+0z
YiaoF6ubFIGeE1SXDfi2Ch2GbaY1PP1tCnbwilQosq0edyHwuwIXv4Z/kkD+0wCH
MvDD2pyy+E3xQfIG/5xVRnG+p1GeMLzomGHkWOHOytLBk2VBDs6jguyRsBppb/hK
7mILTCHk3N9NzEBmvo9aevTJokvpZEOAS41XDQA8MQcvc7MEIrMdmxCKPV+kSpPM
xjzKwokXP2gdpkbEXserf/rqAE5AIACQHmHp1En/04IwAwuc+ivXXEOnKvaGQ4/z
4HH8gZWL5Zs1c2GRrjWnBb2Su8Pn6ue1yKdzX4WO0AOs8SOGWNxDRb1BX/+ERdN6
Bkv8oBtNOdPsi/NJSPNUY1x+eycAFgLovIZS9+PFIScaVvndLQgtfCXkylwXgyO4
KNy5UDag7Kjun2YiILxTKS7TA38m6b5JHt0GIRxbc4dPHb3fhueRXWXd94t27ODp
7JNolzns9Vkx8klw5hfuafSU+iZTE8A025ovQEh2wzkEweiFTP1B3roodcZqMsfd
OvpB8JvFG6bdDu1fDqjDghgb+F+xtll0+UaM41ECwY0qsgiYjYytAx7T8mVqFhhu
OFcKVwo9aF2bfyaAuC8UYzsCh9XVWiLxPPytbtbe+QiPDr4tudMo2URy11Zynnpy
f1YNxEWgSxUxeo0Xjgt9OTpuSE/p4U7xUFaRhCeh/UJK5jqt6xVClzqatvEAzLVG
EnQqJenPmAAO0IAVOJKMFP+pl4FCvmt05cMKSBRmTunY862PJo8mOR8zui7vBwyw
E1MPO16t2uyq7F+Ak7jPIJos95BupggISXAkMkKQBqREeW0CyrKdxFNfkSnk0Dvk
4MvshM8Xc8ZsyWOxtSrzy+dSDnzL8dhJV5mC9xEufxrhUxZjFulUyrX0sRoWHy/U
mjUKHmC7Sr0vIG8+vqh8kNoamw2TaEz0utAotFY7h03SVtmjh2HCnZ0gUcAgtz0B
CvQ+m+na/qTLLObybTKzb4qeURqMl2i88IoWs4QcFasHNOTQnfEpwN4G6sOGIYn6
IarlvsXGOeilUsIOj9L/1ZyZQ0YK9C24eCsZGESArxc9AMeqDK30a5VizwRAC4UC
6GGRx2M8jY6fcuxPBfL1icYLjh8X6IpB0slom897za7jPQU31bB1AhvoNUrjyrkS
FcRhPNd16xs5Or0/XvSnjdQz8amtI0kxFYoqJUhyKdZTKiPX1od1n13btIYpQoeZ
ma3J+lyW872nCgp8F91wO4dqNRsziK9BRi/hvUvWXWALxEkmsWK07K5V0abKIgeX
5+KRGvx0qry7qEz1XEJ9YzoiKORdAZvFoaUMkRwUUII00JiG+L4jkMbSvvBviLjK
y8vOhLEKaxkBi9bxr4Y/WR089VdShDCBdQZe6iEq8JnAeiflB/ryCcOpn22GWdu2
1UGuSddn0qLLjbJt4isPs1Gsxlfnupxx245i+Px1DL+ZDCHdWM8JzEivulZzCD9h
pmAquFZhFffqeeHppBmpmHy2IPitPJ4PvQNQx57DNcOxKVE2iv5F1Xe4g94OXcUZ
I3JW9g2BH/r34bf8iO0gCoRbWRsLlYDlDRp8QvZ7gsGpnMq8+9W1GHz2QBpDFaML
O6AGv+k7xf2HI9v3w/e8HgFOFUlLRB7fuVdPu5Hb5fg72j/3zOiZQD6GY4l9+Nr0
ctr9uDu6aiFktmWLgb+PFfmUpYICpLa2NfgYMBdfyknakb67KZ0TGPu6qCufpf09
sX9bjSbYz9aPe7N9Rt7qlEPmWMVh5UtxKrbCWOteBtQtqYrrkO1vjxXq2gYxJcP/
Gj+S2AatQttIJ5nbdh4MSUSGpY1IOsZaMTcpGllt5eKN5bvEN9dVoUt8pEnlyGKN
7miBHefLKlBJDOjkddj2k47rg03lU0if50xQNHpgBJXG+l7Z9bv0RvzLSgBkFEeU
q82jb4X2a1Gsvx5ZCCrU2uycOSk96glUPvRgp+O77uoInJVoGMHZUvGaR4kmYPsx
n1wFDYtToTI9ZFp8gkgZUSXU0MICTUkRm/IIZam5bzzlhfMRnvSOTDGfpBa7KNWF
kAbxG9zZALuFLJYqW6BnCQ+Aobf85e2jfmcTS9sF1rSPHQQJxtUg1kCgrxkdkwOn
8O+FtpyOj2yN++vWrOsZt8u5qgskqImNX9TZSv624OXzQgRFMKeLd9f5/YZ2VXMZ
Rr4Fqp4S7ihCWKwHqAGAbes9ggOBrhUh6m8ApgNop5pJEytns0oo9Nylul7x1AGh
tjkTlTR/oGcWzomF+ZDyKMkPTs/4UJR9aCaZY5LMlYBGA6iRAQ1VaSkFQBePUMf0
VD4ooogCAt+NM7BVJGbAKCUE3rRkYA79tAlUmiXbkH6c2Fc2zTCWYz3QDw3b+ZPU
KB3Q2/egpfXa6ZdeiMS5Dt2wcqKww4RpfPeYeEIHq+WP5L+vTVCFCvIam8TiXD3/
aluuB4MDPvvnLg1u5UOtN+zBmYujWNgBB5RbQHgUd17w7SAH/wORjEwN4EhwJefs
TC0rekVX/jov7EaSrXTcRhQLFGBgg49pyaM65Ihj+/elVBnmI2lmr6JfOFOb6M3j
JAT9sPkNFrprC0yATFazmQaiZywAuOp/bdUVjL+mwduou6R0ywAOi/ZeZPl6opIy
ZxAFDHnqbfsmleTwYeQhSyIANYofFBT7hXnhZDqo+znE6eyNu1yTUNwRpAHDfav5
Qjcp2UwMx+TYcWPesSjaEHSqZUQBpiyoYafoOvhJku+68UZ4EpIxDQnWDoNasT5E
QezCJcFCot9ycbjqqQtodVwH0vaXp0O3XK5lXpB9dbbP+9yQsFPiZOe0g43I0afV
wZKEronu2zWAEhDdOfN4pKZ6AMWUH8SnzAjf+KSpkH/aEHv2b/dg6heyntUdYVse
ShWVaYXozsL5qGu+gH3Zjml1PVpbOZJpz2zh4WMDptZWCxlVo/SES7OUDGriSHmR
dkEHv3ke4p/5RLnPNc6amjO5oKsns404UOx3nCWE4QvnG/4Vlzh42KjpiRg3dDWC
IX5X88QGEiAbBBUWm0uLA2+GtBxi48tWS/R2GcxwKcQIikPbyHvNcPO0LbYvLGvu
vPr/jG6nXvPeRZTBkjUMlJvoYX2wWk/Dmdox8cSi9xv8cy7ljpz4DTKB/in6q+8p
LUz9nl6EeAl+rBdxonfysYG5sRkpz1/w/gDYwyGh+7n/qQh4Xz+PFReHlD1buCi7
6DoYani2yxNCYesUlhX7f9x3wNLleDv2do5VX/KaNs5OY4Zwfz45kHPnOU/zOxU9
I0T5dvZ7CUCVGibjqm0OzheGf1Hj4FPEpN+5FLc6F2gYXDMzYuMHz8ZI7UWrMdcC
GmHhB9fqlf+mgkfgtxuDYsZ+ptRLOKaGwmg5eEUUP0HmE/NjCxQgs8PdE+DEUWS5
L/bwyqNOxOco4vD2cbsS1UU3CcalwrJ2DZ/ovIu1G7wWXggOMU4lhZdE+OUvntTb
YI25UDbTSCF3/mauvf4Vyp7V/+zdoriXMfpU/mU+TwbXJYyDWgKkoQNCYSUQB4JC
7Bmw4fG4Xvy5q6mCvwuFShMWdaUNE0+DH3ZR1YsEP6MNJDgbj04iDNfvSXgyNhk7
LVIM3Qs6QvjMykVePAU/DjY9226t1VZ8DFmifIRRML0c5fPWjUKayA4fBETxu1JH
XZ/fvHP+U+59Cs6uFdPiQSh5ENZTHumsibmjKXR+LD9Sk5H0AgbpQWjFs19I7alO
KowjU099hIcgeU5fk94wvx1kuP2VjaWQM3dSBSfmrAxRubktdxMPSr4WUdtlT/d8
RtN8Oj1eTrcnM+B+50yxygxyUwpuoOUZ2MuLJQg3T5q1Jhqyy2tzvRsp0JpiVlNJ
iUCrxXdeZDzxe+5tmv38s9kZ5wfUtXlel8YIjfx0iQnkcDj20lsYxEPiNs4pFqqn
wrz8NknsT8EOgK7QFgcr9Mpg2Bwg+lKPhy3Xfog/OILKDPHnqugie7+wJRfJ41Mw
tqehGBOP+0O7MtcmqV/gbaveVcd8a6L8YlrZZUkfTE8ETEs8GEvyOIQ8T0EwnncD
yaN5ybl1NOAWQ+1ljjgoCPgqN+zqpW5oVDdBEDdXMUDo75WUEx3WRauv49LUZRb2
FupQCnnsg+ti7BnZ/t5at/lUKgNpWn6JGaUeKjoUP9W1wQAu7gyGc/dwMaheVI3H
TaiSsBxv5saqSsWzkFojEUm1mMizu5u+ueBt9FeXymBxcVbIUZ8BATrK4BiNhG7x
FXkPm94xS0A0Hwy19JPU0KiAqA5vEqbh5L/DEBiN9Rmu19VL+2OXdLqOWmXHbNwH
pVl4r1I6o8QGwTGz315Ce2Jb0vtd/PD5Ap9XJClhsTNlMir+pVsB1gO0MyB7dPJ9
N7BHIYZz5i/oCJiabYnGXSfoCRUegHEvOfVufOxz+qbGSQ8aExBnM6aPwq4W9luq
sRi8meeRe205bl+vFatB1GI4CASRpgxl//XMAhYNiGqWQnn1vN0TmdK2IOdhvBLQ
XgPPRZw5UYqoPpDCCD4IioXQTpxWPYr2xdYhQxlSeYuJqbZYFCDh0BC1sSTy5r7y
hqFqjw1iLY5lIjXkOoCTKQENiZNsJyAvsAgIaTCXHuDtevTqYkCA7oOnURNc/WcW
sfSEexc2e8eTVqEvVBqF3XN7H6e9B7n4IIvVE31HDpaDhAtSvqEbuUKUcZ9EMJAK
3I0GiZtGIw+TPjE++tAV4xfy3V8fdMC4sjEg6xwSF1RSSLAZL4JdQF3AqOAOHeBP
OBbwVWhjwcM19KEoPwOY5Sbs8P5xuYmP2+6jTpbXx4EhWVrgzdj/PkAWgg7w0nWG
G+sruz4is+dHcOCYjtv5eO6rQCSpW2jQj5xexBoHewrODGrigb68ofE2KO8OuCus
85RRnivziqBPNH0umLJsqLDk5FgQcOWlWgUR9vvOlJCpuq+V1PWk0hAL3D59k/rK
1SxZ4NalG7MHSE3ksbtx26re+TAKA9zEzr2z25cW5Isybten1WkELie+Odg9mm5l
WdU9/zZK9tEQBdf3bGhwAsm9oCnCyIXNEMLbBkSihVcpe9GIA/dV1+C0G1cSCGyy
DBVlRpq/NQlqJj24IhhtGyclQ2Hpy5t+FbGzJGOW8gpMO6t5E+UiwwrGE3Fzn0a9
ZkomW7XBoUV7jEE3prYRqHCgOicl2KCBOLplTK46IjZ2Kg2sPR+SAPY8AJn7oue3
XOBQViQSghqbsB18QoP+oilnkphniIP8RAhm3RdVRnha9GixF5oxX+hUBqbopdcV
ncy1XDZyi49aW7mqxANAt3B9Ht8hfsUXwhiWxobfQXRScV3g8GpP2QEx6GWlflol
gQMuFKlj5+LQvQqsUl+j49WI0cOh0D/5YiYFHnYV4dKH5BVPepGsoO79woi/ydud
u2UpGCHl9McnNw/Jl+cKT+YcPWpJWFGxK3NFcLB6Jl6VTgtPM372SJEeV11qoQij
S4XwyXa3b4obxC3w6DMtNVF0AdLYYROYShJ6vBQYED8jcjWlnsvGDCr19Iha/O/j
iNm8QJsFFaX9FRr+/Bni/5DdXeQMOiPEP5XiwOX3ZHOpA2ZRgIQCPjpGy7g+VTZa
1rwoJV4d3dozT1g/w1AzGPPqrE8mz1zZE7cJyubm0UtDG3cuk3qqearyBJxmvOb2
1BcdU8dPVo/Zrv5RnGzYw1WU/j81Byf8Bd62ciRN7cRgBbyJdCIJ97mCIK/8i3Ac
uZmHNXuV2/8kvWSNo3C6zgFLaf8Tm830fBk8BCARiHR66vWV0eLJxVRq0W+CPxaZ
LIFxu9nEA59mU1jMuu26dKhtDeIJqqMKwwDa+EqVXNmtPgD/QZFtcIAGKTkRSfaf
luekOYAKmj+XacqM70ieaZEQso9ADrJwIWJFkhhhLMq043PwJG7Uy59/RtDja5MN
AECVuXPUrNak2ImqIiys2ogR8NMMxX2hIaIT5l13YWIhkmzGorVtkM97DZ0csh03
ZPkN/BYRXlTW7d7bz+NeKWlqY+I2T6I7WCGnIQQIoHOyBw10yZHxFL+UBLZuLh49
2lPIzLuKmkWiL/vWJNAkRDkhEwywkHX/T4SkaF+PE5oqakkR1DhQmGc9tG5JAa1G
y2CDN6BQzRu2HN09h6qS4zEEYkU1VqyHg/OPkYmDy92QF9AxyW3FQBH6HemWIEmJ
EJzELWKVWr/MtD8F/bLj0Sx0DIiDpjT0+5qULyQ+Lm98/SvqRU2VmGCRzvM6vwyB
n4k00oMzM1eSPYmtggh8jAjRtTUX3OcMt5ucos1gPw+Zj27cIsV9c7ognCm+1Zu6
h/dBizAMHvtKyOjeGd0/64/ZTL6AJFdSZmesCiLFg29zs+lyeE9iYKSOmDssktye
E+WNsSeDqDgm+YzJV2Yk75DRsbVoD7CX5a3NpQkNPO+zLulOxZh9urObxhzx9huV
sw1J0Qi3uucFgOPrydnJCGQt8iezXmo4vy3NVncJd1iX+jZDK0ScwS8rmYL8jaWj
KaygfpVlDI6Vd+4Ya53vKWuKjruulnyZu2Jh3Nk5nwr/xaCrUnhkK5IWziRZN3Uz
LY3C//K2QzWMlnQ8gK4jZVpSHjQDLAXom/Gvw/OCcRg8Bm07gFatCt+qQObZgFPg
f5tLCho7B5x47UOF5tR4yvVPQd7Dlcsa+WgqzTspkRLvLI5Xm35QBrZIlW2vgGBH
z3tF92kGIu1QFz1n7R9CpDHY4ZXzNADlY4TdoMi+Gt5SSbCv7VmpQ6oazpo/DZtt
eAFwcRUlNtRAJe9jWsueSm48cFCuC+07uJaI5jk5aeGCqn7SG5r2rj3CBiXdYPLS
1ldf8D0Ip6LF2PgMD5oSkBOiVWHpiz0KiFaeJisuXwjvqAI53v/uijzfpgNMEy7q
7H9p5yHajbeqWYzaTIORt4quoLYdssV3Jqq8OL4yqKT7pszZpk5mnEqyrklhSYB1
h6C2WgKYjM6eIkNPoGKeLVuln712crY9qRAJU3c/LOiK+LQZUSg26b7OkKA2Xi2A
Uf/ym5b1UQBwaB5aBq17zNox/ugR7mzqU+vzW3PnJttaqOu/wPBJF4GoezCNbs5J
xj/b6HuqaenomqawA0FQmEZ8doXEuzkSMwogBTuPtskFoo+Cms+yOSDqpdV0Si59
OOy7pw4NsycDXaU6dH4/R2WyJ408s+MVrS563ymdB58y1lZQ8HCytmlIStIKbAsx
y6j+fikMiSbTY/gd1XJ6Yw==
`protect END_PROTECTED
