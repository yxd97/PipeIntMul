`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltLUebPYrSn3uRHXhuSjQM0KTFpdakddgHRMkPP5DikGv4J0vyKpQpIwAt1vS5QJ
n60FqgLqlOfdK0YRZ4D2U1Mb8dJtPkT0eboUjK302/zz6IYHDRemccFwSBen8nSs
IZbFyPRGf5aHDslKwkViEP4ErSIUwsBUGK1Ar9rU3qQW75e0ftBvMQbOMS+71lqu
a+g+u/C6Iq4kLkIpLC51G3ob1TnyTDD4HSvXOYoxZD9ToqFhJAqJm+xSf0D1rq1h
YUyLo218dtrqws/APhxqvSZJPnol2S3iC+LZHpOFLdEFmjdXWQuokq8g5pGtLCBR
koD19dZEwHJvaoC38UXKlPihWqzCom7vpVJcDos1qfOEhcQjNfWg6t02GF/mUR/v
EAE2sFnUcZjgK10cI+WMVkLhX1uqDYF04/oJKPpc892rx/kiJmw6ihNfTG7ncMk9
`protect END_PROTECTED
