`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yk/wPSra6hQOcha8748OLLl6CDXiB4aogyjZimxSWD/dMqmVR8wWNXOLkzPDnhbE
/UlIZVZAkE4NHuHQYJCkAsiT+znWpF8cZfL3dd4Xun9zblfNJQnHqPFer6HJMnaz
VCi4xLDlLEh14nIlpRwmvH/XYjCDWy5gwRlFV8bwNx0+yWxqhM/E0DvhvggTO14e
C9is4EacHywtzlMIVcFxQVRVW4F3MkFTX/FOHQHQwMQOr/5YWUS4D/BKf07mA9YW
2QZPonB1C5XkkFfe/akQ1I/yUysAZRZCY2h0qeXtkbnxpCFR4i4YyzGoRZ20OG88
QJ/7wn2lvnIoF2B0KunzZPGHS0GvVgZdkXyCY7sDH3cRstWlO2P9KRQNMJP1hHyY
M2GGockrXKnXvuExTszkECX7mSJ4IRQut9c/EQsS0tyKQWF2vejaEEZsOtC/Bike
+Tdio90NYwp6rX3IVFmLPePPIMAkAbyjfYZtdy4R3Xg=
`protect END_PROTECTED
