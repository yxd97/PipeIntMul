`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LtQkfRfp6tim/+j0mE4iEzTe7dtXD6NkuJRPGHSI5SbfyNbSjAFskS9UdBOoMAJ4
TmZoEE1BopM1c6d33Z7Wh1MoqMNfy+4xr+O5ioJCsjwSmjd/nVc1rC941c3HvfoY
Ogr6AX/34Si5QRvEFRxuRKFCmbqyRVpwKWDaPBfNgJhRVLX2NxRW3zMNEM3P/Wb/
lxjzOiFCLygryAE0Ca1ExPxAwZLNEu/+RRfMBmvCYHZIafB4U6i2tw/07N1ZU8TW
p53p/Wglh1bgK/g7PeQ4m7dUbFrbZR6zPVYaUFyO1TREtl8XbG8Fo7+hN0Wb7D7T
X4giGcJ/s44/2ag8s6rUKl+u0uUHU4i5Je20y8yFA7Q+2OHW7H0a65MM+dqeazm9
hSiMOi847Dl27RmWQWuSwpz+YXraMWpTM//w9G0Ho2IKdpVjGn7kAxAY2lTKTNXV
6DMWcGw5hhgXtBSwGXrveIoE85QYGObeV1Una6H7cGgWK87oqBs+vPvIlX0KxvKP
KHzCTC0VVmPOO2dhWd7pcUcqogMNKKaIpQv337qoiWMZY6U22eaO16tGRuvdLhza
0hrLVvgGl/BI1RjhA1xypqCXbZiBDMRmRIRoPM9DnsviGoi4cysDNeJpSaWdgAR3
zUcK0qP/eVJtyCxSYd6qdJrAd4LM+oltIsLgmVn3+M2quIQqAvqFSz0jGulFUMzx
BPSiqPqofIXvcOCU/dD8t1NXoeWZTjhX9AJPJSnZEF7pweYxUWMcFS2FL6mwwMcb
l7FjsXXH6oE5cqRBo63Mdym7OYLK355qshnRwxx7bOZ3glc+dgkAeMwW85ml+92/
bkURXgPbC8B0D2uc97s7QPr/X28FgN1pNWHi/NedOkHDqjxDlExHVcLajarxicuU
o7qWlFfitsi5GPLhcoW4qNdrvjqWTAOZDnCKP5SYF1gkdchNuycPyyndbaMpkwQy
ow/+hs704/jTYMvxPzY3JX2azN8nG5ysDxd1JLfoq2CxgvKZBaTFID6+HaeDg/zg
bYnpGrj4Q2LmX+QOZWzvhK8jT4riXaKAxkbX26xb+HSNWu7wHtobOrOBAcJpq5bi
iPkBupvvCfopffdCEkCfz083ts0iskmp0hdqk+jLCAXD7WsVU+TJZ/2DQ8GcqFCO
zTnpxf9i6e35oKC9QEStAgsb4u2HDfXr/8hXkY9aAj+VZvD9IOSQzTdyTrUA8Jxa
jJJEhGapR5Te0EspgrZQlG+0r58f6nXMmgN3ZkPbltwy0QZTvkH74wRjK2FBLeSl
yM8nnQeQysCafBH9ns6w4NaIzf0RdaSYUiKbGRwq0Gq1/07fZjgQBSMsKRqquCXf
GW6wVleVfmyUO3r6SvkX1qyVKhFl4530QuaVP2eS30sxNlacqGnuEQQYooys3L55
soR+9PRNvGFUtxZIrTBJ+CGrmX5UqYXe3FpYdamgErNUDa/B2tspobTyhRNpNAkl
lgbUFeDHu4FlIleYKw4cmBp5giafUdK2XIA3B3DF+keOInZK5rUg6+n9/k3qMAjb
T2gN5VM13rOkWV6X+l8ywU9eSSbp1klZxwdT2/Epc4SqkVvJ+lQfx4cfg57qTHN2
BmreI8TDxUN4zXIVFqSLuLf+IZh+HfQ3ejKaA34SSWIstYuqDcNJBsZAOWn0DPiY
ujcbUFZ8hB68VeAdDcAe79FN1mrZqTOKWgpaK90ls+/781CHWbqF3w7lljw+ZhM8
OBj/Am43rcHAg13Oxk+f2cpwA8VLhZ+TS4wGDe4L9RkD3rnjD5p9q8vEUo61VNZh
fVU6n0YuoyA8A7NlKJF8L4RKhDYvTfaCJ7BBQThx62bOMrsMl1fAnbtZfXtDZ/2B
nyNyhTjwjujQFoePi9VHgBe0y5rONtA4EML+VX/WwCj2Fow5TGxQHcVARm6SmoHy
KdjZ56PUYY+743LfNQv7qgWlWHuUnH5Ju2ZF5DiTstWLMDti4kNFUzrDTstVuH2v
NZ/qIxPwLUbktcetfWgRZtGmObvLTBhIYk2Bm+K81zq+WAvNKKAj/UFSewSeWzna
4TLPkC/jMH3yQbu37eCVY97fxmy2WsdSOBX/pIpaGLdgPspfIc+TSYVKJifUHYCu
hB7DOpvrd2GK2kBETBONlpFqHl7eXb6Tq/CiPfR6lPMMdAAruzy+zpvCY5eBUc2I
cL6k/tl0H3j3eq2t4IC4tVC4GstXRnummWrqoBK2iDdLt2zXZIE/dok3j3thQPiS
AMreNfliOqhXlVxOd6UFRYKAiND77uCWSa5Zul7gHgjd+KTAzL/lmnlnISEnaUk7
OVmap+HYl4ZNAkjs0PtIJ25pCQSxuPp7uf/jISfWliupGDXGFwGP8GMpLtfkBJJ6
t2xsl5Unh5z34YoZxKyfkYHO+9eunrQgnPi8coWU3Q762VIq1RW++7fh3Od+Ue17
Wv+66f9AQIPTmEPS6C8w0KPNgkZ5IEe2neWjuf40D4qoZwhjSm9ZsY9WUVJVJ08p
V1sk1IhSVR2D9NIgfak5riAbCgipQolUqb1V6StDJ/jx3M3cuuNaXqM/SYFdhcK6
RkjLfIzxth0oY2F5ulJDLXN45FA6+SFR5OJRczk1WS24cAXIYrrn8DvK+7DqWjdA
5lS2R03j/4fHtA0vfpk4Kmyr3AxoEicVYQTXVV+HUPg=
`protect END_PROTECTED
