`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PFAx3205qfU1kd52qLW2usGxIWkih+n1JjakJ6OvOwJVDe0lGcbwwfDd6Iec8R0u
gdkTd82rO55nQbtZvDHq/0nAy5q/3xoDfl6hiVbpiyssngzESQHbbHzpzzh85jOU
gio9EbMq5902+qfjkUTwJUerxU90lY8LfbIMtwt/e6rUVvKXuawFi0ZKB3CRRYRN
zVcKVAgoroqyWedPDEp1wSFsd+x6GCBswKFPnORg3yc+hW4ki8GzXQcrgW5x8v1K
ZQ3dw+c9vaFzaDkwJQOqGcfj2SdMTuR8D02K4ikD9/oBJNII2xk7gFmzf5uuMIHz
vZN+86/fa+ysZLw4kkZn+3JnCVSMYnkgxi9X9zMytH636YKxi3Rk0v4rfj1FKtNf
R2H4Xok3ZMWF9DDDsltaSY76DCZiKLQVaFv7gqwm1QyMXmsu3hUWEZCJoPP4mgs3
oMe/m7jfvrWP9JXIzTNCplCvbq1+NmixFBj8Bxj5p9l+QdqUMetZspN6yWpmi/Fh
0okS32HvSK4n/hY+Ii9vRdGDtnOt1JfHSfX9jJEbm5YtUKpcJ5E2FsG9ddsLkKKB
kM/tgfaf/q+IroYjrfcKTRLJu/H4WOc2OdVAkyTFFalZHH1ApLo3IRPDaNUgd0xa
hxqPmsn9Xysw8F9rBkzGtMXleZhVH+Nv1Si0rTuSAQTioQ6TTE44z/YmzPsABxYO
+gbzdyzhWkDzBF7IZHGHBsYrCcF8lW+P8f+iEIEhS6jt4LNi5q5B2cspobYr6lPu
lipbQp5pAfVBXKdEF0gtcvE6ylO9CenxjWtmG7lyB0QEkwORK1a63Zl7DWYUG4cs
Trcz3amrDdtlHqXLhDEB+sXmWa7SdN9cN5UaWb/K90l13BOwxWRwl1ZFQZe4zJFO
qv00egYEL2VRt+CyT3dAZEr7fePQZtMXAGKtHFUcR2nPQZ5gOz0qM1QQJ3t2ijm+
LE4US+q57tIIQc77UWwLVgK7sEDE4Ko3OwitOLBnuDdRYqr7aL6d4jioYWyFVHJf
9R3N4HLDs7ZHXpwMpHI+1uhsTHSdF0JbDqsoC/xkBXGcrhwTvphvKQsEi9AjCoja
ndrJIVTzyw0hXDEUQcwKgg==
`protect END_PROTECTED
