`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3k+1hfFrCLbeWjR9ytHT+V6iFsbLlISXQ945vMvokoDdJWF30FsF8hIfZxTfpgwK
kWNdnaJtoMV8OwXeAp7TbhO/v/Zbb/xPRhPeBExwieDSUcM8maW5jiRftcN5PV/x
LUQ1kzjBRcrIKbXJZ4NpRFnB2Wh79BSCbIMIFGS7U50Wz/7NKAoBkPXYsIUE5KHK
MMlby6dkaQY8XILcXrq2aq+9j03ucuB7qxKKK6cKa8IiiRpVDJvvBVaxjfRS/d2B
IYJ4Xb46yu/Z/9IZ5J9J3R2j0krtRtAFpo5u6K6HHU3s7/AMRgsot6bgqMPZU2Hd
rnhlFsDsq53LYugf93eyUyJUapN9oOnFfDKPMvSgMrHmJT2Sra4oXv+ESW1JzJp1
2MGDxAnLFuas7eYg7TSyP/T9NHs6z6068qT8AIJo9KEneBHl/9ll0niXLAdCBSZG
`protect END_PROTECTED
