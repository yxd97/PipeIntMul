`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9uHU7qRA5TYnfb2tGzqCeWTpfTj3MOc3WRs35I9OhgfmYnXYa+eeNynl6hIFVzjm
DDnbopZo2D3yBAA4MDPUiwSG+YqwjPDIBrnHfQctdnHUTX3HcUBIX7Cy7jU6HrUs
1c9cSzfZ+wLR+vRlrSc7y8+vUzVNJhQKKXBWFphs5tbJxAX4YZElRo0dj2pcuEXi
/02vHzbYp7Sjdz5MPdAzWrelZAncPRoMwgSEhb+g3jgsO5oB8ATlSKBidr4ptStZ
1f3EsaN28H5oferQLvjWmyCm5Ih1CmzI68EeJdTxTuv/Tn1iitbWTd6aKjEwPNQ1
aaWG/06eVF110tVpvuckj1X3UoMcnseukzjmuOH8sMAWfMpTmTW/IksnTIEvWLll
v5zIoVwouldPrSVOJ7V9rvuqs/ejiZhLivWBXbhqi2dEx4kGeSCChgc8hhdQG/14
UUgrMbXg+/ou1IaP9+sSIwvJPeTR2V21a11OIKCdkBAtHb1j5EjEL1km1LK+XGTt
UtVs8e/f+QT7dA8pqBNT89odumeBByCZC8pQHBBRU5FPbAdV47wE7fyxaZLmA7fz
LXU5ldYDFn/D0+T811Q5wGc02Uhj2aP7y573kckh6SKWQsjTHOdGvcCRLWgPKsvA
8lyqRNvfpo+RRXr9aC44tYkJc7e6U2i5InGyW80SL5sAKnEV4+LJpQb/i/sY1evD
zH1zF3xtslndEt0HSIOPAmiNLCtOyDDFddASFSdCLJAmVhgT2aa1j4zuFaunYlvx
E53ubeUR5aS/e4/zK8wIBLYcx1iVblEB9qyIUSry9mH3Jlqk2XIvS0b+hnOKNCQ5
D/7ocfjeKGhf2RNinv51w0743z1w4Oo9FbSPm1wf+rvtaXp/EnaqjORu0moXNQNK
oy82oJT9oBWH9xzD1mvxMlhkRXrdz2Q3B4AYtl1VpHIEH2Vzeic0EbabmVu/6Ign
JQ1xKDj7PkKvVYPNwsqhw6cmsZunU3Rn8UJ1f1LWb7M=
`protect END_PROTECTED
