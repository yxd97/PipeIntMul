`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbC2Rg62W2QhkzSkAQfjxkc0GpJgs3/1CVqsRJF+o3V1sLTZ8qwbDmNvv27uKh/Q
kRVq6oUqBruIf/Yd6VRbytwp2IlglMp9jcfQisWtjMRB1zwcZ5BA/bRbJYec2Jhl
rgR929zuQcZd7LisjkXKWXkdw6ec1iom+BBWk2eeuhXPp933wPg3PpObIiaDFQRs
QIgBBkacGugyNiLE/MVmaylkqJ+jtZ7BJAtYvEW4lGJk7iwQX7R354BpZG6SCiFu
h0hsUgTni1IlxmuzldXX5rCGuKYZokCdTfVfOKE5ej09nTSTSt3Fex9s71Fqby0B
8t9O5kgQjCw2TxG5Wf6QRPcmUMmzqFxQcuO/jRdVa+62sPgp6/Im5fROT0GFFuwa
VCFzB3+U62ow85GH7RuROEtWGTLTWSGTvpMViCT0gQqlc+viMC1Kv7JvaLlwBNKu
dkf3dJGresLV9T6Tec1kMxn72IXlIKL3ZCmSOiu5H+0=
`protect END_PROTECTED
