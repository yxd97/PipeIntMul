`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r68z9GM6LKw4MPwtCt8seZRIpWi0jGvkSd/mRxr/tIGmElmrDVpLreNvt9QSLCwg
h7FWd1zZOQzQ1cUgPRiRyU4YkTYuUZ/z0Npf8C7W4HuaQLWv0PlAljSLtGUoGdbl
pp5+5ONyOhBnFBHwsCT4eQh06gJOoorIm7yPlSo3kmR/kaF7RYnkdY4Ct0UJ81/9
GtEZ3VcLJDLSYhxS5DBXmx3Mvt7xU5o8+P5UPKCXhHClp0M7tKOAcajD1MLZ70MM
SEuuAOfah6i22tCSdmVMJlNfO0RPT6UUz4fH8spD2dARfDnAC4ejoQGwTcG8ndAf
zh90wiAQEeA9Ngb2MYrrcuV9e0LTnbzXDO9WetNHDXD0zgWnEuVRRg9Fy+3y0UKe
z/u8H1lhCYeggbV1fCil0fgx5Awx67AnR28YO6a1LPNuCfyVnDBLv3BGY24K2sKz
H1PGtfq5IGU8azYDr6xPu5s3SbVNueWo6XDEIOUwXtGr838n2FgyGwErLJniyC/w
GPA3YPcakBRrTQ9cpSe4GVKWxgOENKEvZLkMx+xnivvRjT0whgnlavURg7dK808z
8VL9fsCSY5o1I7mUr58FVVMuYSEDWtfhg+O6YCWvKsTN3AnppbfGbR6Gz0nvIem1
KfMsu+bjWtng9A6XJYDjPQ==
`protect END_PROTECTED
