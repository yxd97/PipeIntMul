`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ENC4nbC/7/VTYC/lB6e/mk5Pi0q2N7riqW3o+1yaG7FX43tvN2OQb5EHpzKs9ewM
XILAeJDo7iqiDYvUvAD9umMmwU0wbsiaQQSWS1zzP5So82MselPu/1Z/dvxAkF8B
1b9Xeg6EeWJSBAxZx0BoLG+MTVAE3mqCbv8MpLbmbzg/MP+/tjSwpAHXyyS2EyaL
Y/QEXj3j+0H0wQTT2zOqYbB3ODUTMMacwH1SILP42YjeftprQGHqtHqgiMYoYu7Q
Gl/QACD/LWDSVpb6/wWz5TYGMhyw9zeTO/6yZSTSmIJlboxVBO8tGQAvX2cx+ubN
xdixbc5jpexws8AU4B8Pw82WZpNwZp9Li+qYya2ZEkWVX8kcT+dwQJQnZfZeanyx
PQz+Z1Y6wd4fGSiLsT5EgrIJlyg8/oCd7NN1p9KVsrDIvgPhSheB9KOmteyRY50c
8ns9G1v6ombmrixBrMf0n//KFmQ07IQRfUKX4AwjMRJpG0cHZ9xeZmZEHLgksBa3
EP73Shrd9JS0heXWam3KwYzxCRg8v3atMevd4274WKoXfa1hiJ9npS2bilrSE0CE
Brvn6+XnfPmJk0+9rRHNNVFU4Kn8mRWY7qFc5sbqLJHhCjzVf4pZP1dfp8/z5iCM
RbErh6zsLT8V0PVmSDN28ot6K3zfviER/jKCpvoHKYLdri+8qfswKP+YSboHeuW7
ziaQUVLMECDWH0xl1zpGUWLptYtBfJJqClrElQrfal3dKBVJ8jpIiuNNEG6llgjj
aKkXvOSqi5XRI8w8wyooo9fg4fbqOdfWRP/yFlGocCql8oV92U5hTEKBsJ7N7MYa
p2t5hLI4umjJwM6sh+V+1tlHm3XivZrmg2XS3aFzEZroY+GnNI43YeCIYnIEDe5M
0tx9+/fAQDX1kjkViG8mF23QcKdAHety/KRFE0NcaJeU1aQ/3mDQTOf07p2xkJC8
Wlnbx5Eu9Zz3+9F2mbJkeWEn2r+y3/5UoJHcp+aK4JNUg2/W0wRPvzvHB4xoRiGD
CLV425F1SQqswA97aW4JKtosAB0tILkBvYMPdUlaQtkdubqj+23v0FPaerZIu3Yw
o9MCOxR0jgjceJbD1sPuYr4bYqrrrezq75QW4choSeim9Wr8+KcDAqT5Rd4CzLru
cTSPeH5O/2il8kuPO6E97MdSJGsruJCLrx3M13j2dIoWFm4t74x2XUIhYWdsaTyj
geWjbDOrrYIZL+m5SXCYPUDGiQM8cCqigNkseHauRMZ0ODdxYqJgS/xRkQ6XIeYb
iAI9cJ2cnfpDWpgpnPtFGufhOZMbukb85Horvzhb7DXUIVUycmhjUUrtxDTWDULa
P2w6rgBXSAEj26kSQTYQbJR6JVHBkMRk+R+HUpMBxj5ZR/JWF4T8SamUSVrTt0Wx
mZbffpViJJ/4S7SMzR8yeWFbg4BrgqH1YT7itOODUZAkZdUrstERmhMvLzz0QsTV
R3Pgo5L0wrzppSty2MBTlgBsm+VMATcr8/H9PxwxYdrOrEsNO05pEcwW5kyhjpZ1
30vMU3h5fZhvxCQYwAhaE2ugwJs5Fr+nic0PbcFvTdinh/pK7HmacGClROHqbX6a
symHWV5o0oh1R4NclY9UdhLDHswQODArl6yd1JVgvrt1pSM2O6mhgN73uOS0NifT
g9BrgO6Eh2jTm26/2XiH7YtwS9f88lKaqdOxirvknfaXVr1+Yb8DEAJ8OKEmkf92
xkKnPH4RKQF8Y/PjD55RY8kOw6KSM4VYYeAMHO/LY1R0cnrdx7KX80Y9siMwA8hx
ovuJrnV9G+gOYzpllwyfVimOLcumWXk4BRMXUskw8xqno3apOU+BwwCo4tZ0732A
+yeNB4qMsbEVjB4j0+73GZ2yQoGmFB9OD+5DxWN5x/XOdn4bjUNQ5cVoXBCtXOEa
2TQXBBLe5waVSz7n46FIr3f+EfO13yE7xA1wM5XG2BR4pSjmORlv9SGLVng9CJus
+ZN/5/kBP56LPNguxl3xuxBy7eDl5k2BK77Ruc+zd6pqrw6a0UvIjuZBtl+HmCVS
m2d/36zOHheu4RttBXzludZZHzMo820/w8uW2U/t6FBkqneW5EG6c1ARlObw8aDa
Wx+jBBD7JrV+pDrpbT9uBSErkjq81UQLIH8MDUCii/Cc2pis1bFeV/CUrUxH4J31
sotCT6iux1SRRxlNJC2iKY8aQ3kaszv8bEhtbmdkqOeaekmXXqLIOSu/p/rRSNZ8
iFkrlAYPTulC0R5B/btfYzKjFh1dLDWgigU13LvxmeGGyckwUMcXzcwipseqNtWf
oaGgkzWvKYPHpVh13mqaFwVNTwHDPWL/00dLRrYtds82spfi/+dbb7f2cyBHUvTh
vNzCQuRg9pAeAm3qv3RXOtbueqT2fzd9ZXT9JU7OgBuEhqLD9flKHL/4xSGvMQsK
yAQpSeirICHuZHIK1iKncjpC6aRFVUI2uyUBVtb2WDQVxpt2EJr6E0PrqePitGS9
1qCjA+yDFQrRIn9iijiYLUhtAA6dUeiorIko49O4qa4pxYGfSziEpQuUMx0t6FVQ
0j7mQbMC9RQbusxAh8f7EIKDptJGrhfiI+S3z9HNiQ/4TnPnUtzr0j4adALtjFAi
s05tNCE3hKgvqKF7ns1HPHtFvBTmJ7QZmJ2uQCWkAaGoaf9RB5MmB8LDXRiJiTe4
HLJc5MbxX3PZWcQBTag9peQg0BfMj30Rvfl9UyqPjecbDiuqsFrf3Zt0CUrE6VYN
52YZ5o66eg6R3pVcEi3Ncd737+GQJ2lMsq4wuyW2uHDzYqGRcSY0L40mTsr/VYpQ
NILoWl+c5DyH+//qgooNuNWdVu54sMJ+eY0YdwhjXw3xw/wx6y9DyGrmwCqQi/7B
w1Wb539hOznnHofg7iHGvJz1zocifeHdGuX5eLrmQbP2hGJNw52f0QEGs8ai+Gz1
f2R9O97D1XE43wtxTsB4rySbViluhNL7KFvJqoRXFcsTeiiAQ2aqEyGM5OLGmWPf
eE66r8BLwto7aUd9TEr3xsqxACQlhBOJdSiTuCScXCq4Iag5VzBLYg3Kdn13DsDL
kY3VGjfYdI4NvCs6M8aaG/SdHfeCb+phbKVbju+n5U1zuVLmq+B6xoi4SKch4HPj
Znd3HhXzU/8ZoKkUBPchUhnTSLnAmNeINPW/ACSyDNIderEifHP7wG4ELupr9Yis
YC/mSgO7AF9+Opx8uuyRl0IIKtXzNtkiEdNHHSXBaAb7fzqSQmIY8QN79sN65E2u
9A2ZSW4CgiVFJugL4FcP1GmML73wP8kKzq5LzRG921tdkO4cC6aFOaCUOS/rs3bY
lboQT8auCRNbDt9DjqKnIVd9cmsXkYmTM+eYDKTBr1An/u5xWvyQlxFam0sxzDxX
Lr+1weDJQuvCGoE+4V99KgtM/QQ7tn5P6+2RlWpsoX55X+jxXWy9/xgTiY7gMQnD
Ou30PeeKpomeiw2UhQvnQNdFVKRj8i266XBHTCTG9c/halPGC2lrO1FwC7QChh8o
7EbebCgZ823DCxpdnTNLFC8rGoITu2s9n+l2DYUtxjqTuON2EChJU7oEk8t0m6rQ
8ld3oJvokfPYHNQv3hHJeU6r3nBIz31Jiq2cMXFX03VwIfPP3tQ3PdbmEcHnuNvc
2PhICuDNnZeLqa/67zijSwEeSr0mLyKadG3fJvHTKgclMpXFexpt74Mc/ozyNoRF
6eyGPOODzhEvV9rwEWAR7s9Qimr6eOkDtbojQImf5+ofPAuXpfVVfUqSPB1LNiNh
MoTcR2KmwzRz0dFvQFUs2FCocSE2bb6uxUi0eSGvCg/GRLJV0/LHovnZ/N/tIh2e
T5/ZLgcKbUG1lM+PyPwXF8j+BShJbGQe8hKIKbacHaEua5s3k96cY2cMUFhqomca
I0ws1KXGDFusXXCSSY9ZwbVS93MH/YIulnEq86xA+ej4GuYcvQRoBut2SKPEaXBs
f76vU+bcy8jfGMdpAiFhKKhWuSAXcAQZOhKm83+fsKHiiKXpFfga59qHgYBO0Vd8
QyzPsKbBK/lsiVH/COgh9d3eag1x2Vgq/1NrmlqC7H8xN1cxP3A+tcXJvMRTON0T
bgaU+DLF9FOaDXKd4874PS5mnlfN+VEgMV4t2DfOXEoZ9BxFmnw5UiDehVwTEH4V
B6FXOSyriePqAPlGh3qrfXsMi8NSSPn7Tu4+I0JN3aVZ5wansZleUU/cIRYtinNw
rfpMVfcS8yHTiB5ry7B4YYfLuykdFqho8VI00JWcmT/mdMmRuHbvcmdLeIluO+Uy
c4VxY4qWFMl1WrGNs2DI1RBLYt32WkNC2ajQnRXYDGanwd+HvZAUrAjsgGncvfkr
Ak4jsyYb13uYRzbaITdxHCbCTMRtOtejlVp6A7S0pX9udH2t0F1PCP1U9ztfm0BA
elqtJatSjgb3jyL59TZCdDXhoE76U3m/h+cN6bvr/DRXscrFSFbpez/1X0QXeRG3
yjnUiAp6CO0COrsTCRyzDD95IMw/x1fXbZi4Itlvk0Q0If8hZDb9kzsBv59p8Z8k
L2Qi+Fg7ISo3oY9H+EXCWOAJdGT48HDXXrTeeaVI6TrKHeiJzWqe1O770Z+MN/CB
dJG3A+KEHtG+BgF4FvUF0A9Lx8B4erz4CdelwdhUNT8tooDgzLFZZnyzUzKT48dy
0pQ8lrT0d54tFDoQyjQPnbCrgDDuGov9SnQQQbeM9MscfuObb2GCdrH/xPNr0ycr
MBzNFtSajGUX0pPFox0NELEJ1l+6oaFiZbb4iHIDMDgJrepJ1QxjapM1It6BCYcR
AFs80srwH/DIw1vNbhejKwtcWU9Pm+E6Q1VBKpjBoNU4EyZo1jSe8u8Ld6UNmNJM
G/mQUPHruVW9nL5r5yvHfkwLXbnpcB9q8cA/3FmD5kaWcUh7qC9oMnxXEOwc1Gxf
mcTUH/7gm7W4zhMtxp3bMCrLP/PZgYJssjRRgvJfP5MzN1fy84NCyuASIJF9xCk/
8OSAP7B1bXiAqS0+YLcPCXmKhCgiVtL/019xDczLtInt+VpgPNgoTLdX9memC9xF
CgLMEi84ZBKTK2C7IsMLwlJclvBRwECv7xSdago0l6ZxmOucK5XJv2IaSRvjQ0Jn
rHSmq7JeXrOPcDYIXnC1vnyHco57W/gUTMXrgOvR45SQfQCgqAZwtaDYNxif/Jmd
tYWHPYt8i8nUd8usf0J5I/BqvF6Er4BXSwUFw8czfJhPwEBVn/157M5v3B8Xe8AL
Z2pD/MIKVJZXhHox4qowxtoogaVZ/8S54xKm3ftKwVKvHfkHGp71pN5THFvGNN5g
GpJmA1RN9efKopsUZxcZ+qBFLO2fe0lvU+mghNtriPRiuGfoZx2l/f8mRyNE5ARX
8nOoyknQMLf6Goqq+jJ2UUtpk075XpPRuWXei0N+EF2LM/J7ASVa6X4o6kvt4egk
0j3wDo93Vj3ElXyM9O6yyvlThJtjrmWQ65sky/BVZLfcyVe3czY80BEDg87pFhfk
EERa8Ao84C203gM4FG+DuXb2TbRJcDXxGxUxWTFhKG5Vc9PKwwfV0kp8A8SpUSEH
Zn7BhE79Q2lZUP5YzD/vXaaaTCJ9FzRsD5uIEYeIRGQs29g+LpvgWsD5SQO4AAoE
YyMz1n9OALmbdJYlraNSWBlHQugfPVP0XRvjzuXLIbJydZrEaL2ahpdCqVFdcKDk
tHkKwYYjA0DOYKzembv637JK8Y0hqPr5l68s3oU8jWgGfFv30x3oh4vwSE/UQjCl
XxM4OGtLcGtuoZ1ezUb3+v5YcBAPAP4p0+yEM5lqkP4PsJoas4qWyFkJV3gTfmdU
5oADigdj2OKvD1GVz03sTbPkseX+VXD1dNYOAU0Lzwd6W4DZqWpgPsDYWZpq0PY+
i3m0bg2o5uqcfpVJhpN43Qn2frqR6XTCnAFfjJbbn3L8UmGamFn/MO8UjnuNZM7x
HTFnJOFBC8Pv2AmrQNPi/mMxoEfScTdcF7vDlmNNrcV4GFMOBidwmu6YhgN2IfDS
pVVIEgWQvdJlUbBcMi9FrLkCg9XDwQZGkCwWjS4HAyjRYvYoYxcg3sWBbvvUb4ot
EldPNWIVVthZw0+2D+V99yf1U/DhhffDX3xtKLjTvYQExEStJeJF8SLc0rGN+dQr
m5mFlG2VZK8KYKl34jMRWQL7dJlKnFDWxEHyHkoN/G9/B0QUbd0VuKP4wxO8Qg66
xMy2Tbjegl11i28lWV9fUYy4CB2Ht4riSAa7gV/vfVT+9p1KVMakHdqiv0uC10ha
x+pK3fIOgAi/vHlH0t87lZrWUnJ6ULbwJrhFli97oyviiuT099rQxfsW0mpxAVFo
N8q4sQ4trE3Lc7ewr4FWdbO9Ra398Xcq/dxDxC2SPWAiLE2mf97fKKDI2DYtu+is
U/8gLohl/xnd9zhhoMTCEn2Z1l0QNeU4glejhj8Dp9XItdlv7qjmXDMftGQn1Swv
fasJWPRjzHInvxgreeMoR0OPv/ynAXfZN4g75yZ3Zw9JinBOQlasOYmvCUdX62+L
gBWN1frLKa53CqxzBG5uJaoG+ZK6IZIqLhvH9MpnRXeH97lV6hCbr8ym9ZspVRsH
GoyeoFz7KYn4LP44AqD90dCCNmeS4DLPpvT1iGEYsZghb4s/lmBvfc8pBU/U0RD+
Hx9pEGgFarMXgBhLypU/2QL6L1eLz65EVhRb3aAn91k7mgM2zcDUHkJs1OzoI5oP
numa5A80l8pPm54bUys5banQtTEHpNOeR2TeOiqw5MowzytdWgSYI5mq0VYUokc4
5Vbah+ZpCOjviRz6VpQeinwDr9XphgEm5Vx69PvPQRYDCILOmgMIgAUq/hBIC+xQ
JV070B4fpomoZOHZ9tyMeZsyWw8mFgK8tVXIBTCDthPkyT39Whos3dVCgPp24Ps6
ZnWwBFwrEmcZU33JXe/Li3ZnIxp63kwFAk66Cmc2q2YYwvPRHe/cNhJYoAImVQa4
0BuEnFlfNiQDB1MtoBaO1EfOqyZqcIw7WaPqvZIUFrgTOGA3qsEYgdp/3msaGoEF
ShrYMuhfWl8DeAU3pUMPYMoBeljetmLDKp67IAIr5kZJmk1HhTfW73VxPQbBvLpf
Dy6VapKUeVZYyEcwLc0hzJPwsg5EUm6AGk2kL+VnAR1NHAn6Vdl3Wf/V/H7mCna2
EzoadHl7EARc69iuZgSJuVJmfOG4Mp0vqGJrVEt49B/l7PeKJFkhzU0+Xd2vhKCw
4b3MPfKkwkxvstf1Zep1/fl3TqVs8jxbjq5tiMbrnvjmWywzE5tXKEWWKqgOFILM
wi/uFjurIWYrzE5gSx/qZgccAeX89wQuQhz9kBRmN0YfmMEUiJZ7EXun7hpnZiOI
Osd4eW0MUCV5iuBa/+q0ljgfOuunXfQQYkPTR4CkVtsPrttQNJ86bfIHA286sWhM
5RvQi+rLtvnkFCyjdkL/g3BuKvLwOPUI2o/6n6Wkw2ODSIiBBhRXVe69hLh9Sbip
TwXTDF6OZrWNP0zX63Toeqrp9ZqgQLgZ5ZST2dv8aj0WNp/8cpOOPL9Tgn4QxcCC
ArUQJjJD/wC8bSK732ZdzYaEOpQr+20+gh57W2dNzbhwMnTCWo87rsUxEox1zhdz
RFNywWhs97tBA5i4rJGgGgmC9hecdt+0YY76a5PaXYy6H3hsiVdt9w5YoOr9Y43W
FWLq78Sg2e2NVJw4HuwlrfBOIHSHo60ooCkOqkfT74t49+qKl9QxUXuGmpgOziVv
ggbGk5WUQkXB2ScEoNkDkuROwuLTKnh9UBWw6OBXjAjq68uTzRzVFeEcuPAzlRxH
Mzh3iTg6r0WsTm4RBkBRs/LgQ/KtgPJCHmlzaaRlmKng8v7NIZtFzghdj0aGlRp+
XI7Vi+/9FZ5WtUM/zD1oDgSI/Y4vqoYWB+3aPGrAIhTsYkjx3xoa49dYg0RrvNT7
WUn7OJKkg63X5wdTz3dtew5oaHMkZ6MdJg2j79fiIsn8WT/ejuMx6aSu25TmzLYb
3h//rn/fW5ZySHq/cHc/IHkhPJAK5+viK41PR1hSOked89rmLtBZGtpTdsufYJbh
OipwSKCrBM2VYslpyDS/Q8XeMkDjZRNUeAyqDFbEn4JCoClZJzJRPnWiQt8q+/uT
dEsS9b/0xA5G7rLKL+9Y6RCQq7e0HLE2r6xkAQoAGXJXf5w3qUERQtGNNJ0eK80p
BpuX6+8BWfZS1ZyH34FIJK7WsI+wd04S88tiGVwLwaar/KYV7+rqYF51i992KSFp
D/WHdvObxH2OutC8oyKX4L9HaNtfG2KN3K8aGyRQX4rBcHJxsPCzwqLrMz9ksXyC
gqjJjPA9GpTnbGz+HztmcddfibrMCiIgipY0KeAuVrttGdg/CHsx9YiCCwa7+exH
2UdPZ1u6Te7/Kp5h2JsmCAr72/dGK0A66wy22aLfr3J/NRpXlEZOOC44BvlqiBiB
O75blvrAo19a1Z6lCUdV4EZ2QvgG3/jT9JZVsDFx366YMbCg+ncm60PgWJkilyGx
yKwEeiF/VPt6D0rpyq6xQp3VpNJonpP4yyiH0y9KwoVZaX6A6ZG6FuZeKIh13lsJ
KFGXR7OCv3d3UR7/g+AVsyxx86v+dtOmlo1DuzM7l90WmnZzV2tSxDkW/1bBFdNI
Ja8+rDv9sTExNIihXDLQ9W5yHe6KLBCspq29q1SY419B2YYomt2PxSQstVP8f914
9X4y8ewkvpJp6Lz1MFqYs7Cz9cTbUpgSKbpW9ATyIsVGJWtRljFNwZSoPVsCIDeC
/JE2DmLBxWrIlJzYFYih7Z8XFGC6Fy0ww0yT+XtqIFC85+i4ogw7jy+kk/m32R1E
X1vb2leuRXSHHaTCWEDvsmqi5LiwNX79F+3ebYqfON7vbeID3BxfGwQ4fHa2iRA2
KLYFYLX0l6tmwZbYmIoWt0aBynRncyukLUhfkoa5nKzioEzLHKYpA2LfufKD26Gr
DvCq0carbSzefaDwv+E/jjq9haBE9ixW+NUPTe4d1nL4uH/CCQWkP3v3IiO0VNFp
uZ2sh1AFWWaZhdN9r/usZJc2kZMjMZKT+oXaasPksM/xSPJDnphLteMHLeonsQD3
24AFUBQ9vmiYwsHjGvEXtGYPynCboe3a6JST1OtXLQ3/yWdVpxe8+2Cfg0mc+hVp
zCVJ2SfpyaejTABhaaNB9tpdw719boherjXb1HKJBX10i2uT4iD04ZvtQNYDbGep
YdHCCe+eBCnSy669WjoKcXO1v9mV1RoehYpvvyUFhTl1C/q39OEa73kikUhZS0rD
VUZ4IXTK1OThsm/FQ3YzY3o4Fqe6BsN5tl1xFv3bS4fVfNPk4eFpiXYxOrCIM+p8
RgpKx7RlKgp/kHJweQez0eYWTQISfwJs/F7vmID1Zu6fwNwkTTCguQUaplsM6L2F
XM2+9bkcJn4UGzeiGIw24WbVIskbAKYlHtnWcQfD9jWxleiL4IL0AW6hKfOQ6aiD
d9wzwsU2r4gfKPPBdiy7bP8UTK5dcJD8AYpafYKl6zgFXaNFrrJeoiu1Cf3DDUMo
/7Gd6BiENcmOX2EhheqkGxZvMunee8XdZt4Wnl0ovIuirDOin/0FXLUqG6Ktjf2X
U1waPhhDgp5CwsLIVTdmajLCj9PUa0sOjUw+I/se1Xxznyt5HBETGxvF4+8CaqOo
tyHTZ012duCjaoPiLP7CXiQCNWSucBfEic2YbPAZfZ3XeGNu44OQaic935VEFMh7
YlC/MQQjOPQOOWlg+cEW8eLbFxKhy2IsTnStY3fbpqSgR0GRr1xJ38tf0ibtc8d6
2agmjbpxTcIWGMI9Gm7aMHpCEjW3KVqK6Golf5BQ5t26Kb1+prJ1Mis0Vy8ZOMul
ggzRBWieWMl28OeGelId3XG+EDikmZgRf0x3FVo95SMOG4rs6CJz/JYpNVVR9VAF
6XFzKp0Nm5WNrFKokG7p4d1FvpopsZbGjejVPoh50OsqRf4PT9dT9yIsHv4TNn+C
JjsbK5zPWyjJyTTw6GmGFtSwXao9b3pGmYNFd/IHSJhMYQbRr0WXvgO6nNZx1iFv
uZwUcxJotSMfwwcSy38+KTVClbZwLUS3F0QBSRzfvMGmVUJe11dERLDQd1mtV3KK
FjKMhN5vwuDjUZlL/Odw/kyKHkpLhA9iFJQ+V71xrxddsi+lLpHQ7bsM9SZB7JSH
Ur8Gcsz6pdgPWbpttuccbURrLscF+dXB2rq+a7cWmSxHTgQTsoEHJ2auI99eMeu6
P+RrcSY1UXCtvIByB437Q4H563PFj33i8jotDtfAqARZQS2TTjosZirPNHOB6BIp
UgyXsNF3Y72Y1B7azGm9LrKvmV+trxQF5IE7E7nPYmaorSpvYOvBdFG5Lj7nOvNb
sgCDp9SjOHMw9HzWUuZNAd92eqaSmCuEJFiDg0O+CYg=
`protect END_PROTECTED
