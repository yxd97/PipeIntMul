`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6TGUwpPKo92uwjJhkrPu06NGOH0yrMhDEYek0AIPrKF6oJLG8D58oouJm7IQzSzm
mMNYwquCWhnhvgWU6lZuBSAW7CUs+l5obvan6CF43cdGG7EvTIBkCyqZMxQ3XU0P
8DS2xelJR7mNBTN4KI/Wss/7MTUm7W0Qb9XAir+j82xIwhBJ2as78Cydx57/4kVE
n5EfUKPe/GyinxBbtFAMboMb6HX09caDOl01De+9IvW5zJnUgCkmYMG3uk6XVIJc
3Xe0mLYDXO7Mvi0idyDDOvV8C5I0U/RYqKMgKYn331wTLxnlYCJBnCo9Dvj3gSkA
Unz6duGgzGTfuMN1r7yexFp2I1gsThsg4uOndfstZ4c/6dnRUVqUvBBsmMbuurUf
ucK84uvnJrBebb09Mzh6H7NYdUFAikKCU5aRR7sV5VmhnY2VJgNgAXFM2ngNMRco
GLFOBzT0jd4XHVoZ2QaSU67EUYORTClfhxRThLu2ETiHo+nfEcE6fP5Tyi/42DeV
GjZcDzb7RijAF8iR1fgrhNvG58qqJKy5rRRDK2S4EpYQqUdWGxTh88xCfj7V6hdd
3qzOHgsfp316wRMB5eWIGvdeQVEOEgl/TXaTmqrd5GJBb03yAkhbQJpnjdbdV2sV
msl5G4HWY6zNZuLyNtm2Agf1Oib1lQFRUJKZ0NsEjMdLMfejOlNjqpiUdhftVBq4
+0vfZSVFWu02LHTaAdp8RWpTvF8Mg12v3cXd+14ocgLa16PTcCfWxe6lQX05wSwP
w0R2rJlnRq0k6JCGI31k0IDWC+WmlNXijzHwp926g01s9p/0WUl4Febo+6KR6au4
pi4q3j0+v9JU27geUDVbCqnKqSc1HPNajKvSM2YdU70eND+dRTnqd4s32AVzIrpO
ctXJ8d6irQyrvkoNXjs0rf14boRGEHWsmNsrwzOhHLZ4fKhQ0hEJspSP7f4J90w/
AK8hAUuWflaFW8VfcnFIfHZkKnR0wvsxgSTpwQFbeD4MdqFPohjk0hPD0Aqq063m
ZI1kqsbO/10HqwMIUT4wu1laBaLz1sD665pRjv+Wo0GlJIJIFw38QWimjiL7JDkP
y4MBg89QHorRcFNix7vaR2FTKzIXNr49tGaIuv3I7ArWf7fvu05Z3RjLW9/t7TF1
70c1onwHejoGsrn79gCHgbgB54uczoagHN6M9jdSKT6bYNbEDQY67BHi9VF5zw2P
VsuDsNxncRntBlB9KtNhXzYqFLOdUwIXJyM5v7grCyU+hTXlCZoQ5VQfbqvKSXqg
rTPIOGXCkJ3u5D2NrQohwICF+AtCkczfAHgjQ/IGsflJhfkVFsOpvPx7YKpcKCEB
iGNumiWMPZDmI/zUEV9AN/hSz3EzkHNtTgOZQopP2FfES6zpdc/Kti6OGJ9FRuHd
E9zCKowtb+XJzn8Eyvpom8Fsvb+USXTMzyuqYeXryA9QV/FfJRMJ8SHya0+ARxSc
YAEy6s0kInMslLy1YK9ATDsm4MXPFBTCXKmEe9UzEZz33JOLaVSlJjdtYSLB9y3I
oES+jvsRo42xRi1XlTWYxf21HLKDO3W7eaZ5cDE2hlu8u3iL2OGnhPdqExzZNqcm
Z/cHUVRm9BEvnbDx50dHouxDqcElytfUSbQSBepG9wA8cC4BGQJeWNZjsMtJEAoV
woXX/PIC5yKpJY4pfsh/ahRQahQPD4rxzgaZxuNgoNVv4lMz8XjTjISzfVwarYhu
sLlldRGyJbtCV5Rj8BQ1GYHhm9Vz6d/V4lXzr1ZdTzvaVOTyl3IbaQ7oStXFRcup
993SpqtTO99fKSetphkmTSD37opsO6WNLij8jJ/S3++z+xDLTkOL+PwGpnw7H1bZ
TdJT8TnqP8wfoMXksC8587gde3hytlujsbNFzoBdLxTzIxMVL9WXVdEsDI23UHvf
Mo52U+mtxBmClE14ZdxENOCk+PGfpqPF01Mlou4BbbCJNP5cesxZrCcEbMQqzxVJ
G/xCCN8F6T2lCmwUYekCopHHhPoYPnHQMaixUpqTxwD0+lHOPT76TD5kfKS2/WNg
MMbxQZ6Z4GQcQV25eApmrgIemG21AvTcDuRZWjKHbiaw1YARV3mgu3qqqlw3DyVB
pgP6cqLv9wQlV6iVrxkIo8hi8A1Xtoo6b2/jIWQnJNXTE1l/vTeC/FVDHLyfqEJD
OaEYwkRXJarmocHG4Td3rkoYafuGzmlF2pjNszDeVgPXlx3QVuw3sRbfJgzMpsnn
th0ZbA1wGKfCpo5VlHxG7nTl1dtu6wQZnK0giVDr3QmYoHGuOfZe4bNZfMWBqCci
Ut4SHnBcUu394QnNYuMDj311f9yUGRs8OsM72DeSATQFY4L4eEVepSqpXpI/x6Ep
0+niHizxNWkxu3jZzATi+l4GMnGJhlb/NC1fRRy+ufVWaQV6wbMfVtZLIk/PVu4T
pu4VvnQHYdX7qoqVVu6Rsjn7gZASEtZ71zofiyZXK76x8IR5LDWvZxVeeQWXxLLJ
k4DhDOvRT0ow416g4RV3+YcLWJWqNNQ17fBYsTEeAsdECSITs8tu+cozy7VABG7p
lAvuO57Fg5D4qNmA+nzAl07XcA4itrUSjVVvoi1HrWe8VjVEHOaeuqbpQMc0VC67
XzJTVK/E97K2qzNm5k7QLGoGK8LaPX/MtRNLt/Mi04QUzd7EdRvAss/LNTx1Q9Q+
JTnahPzEBby0a3boVdwWgwnSSCLkaM22/Aq/u1quyZq6wVB0QKrGdbgYriXThlyo
XHBruCKv2cq2fFFBNSIW4Y2VK6Pano1W0McRmZa/zTxwd9z4+UdDaIOu5C+yklF3
prPtHIIVVs5YyXKK5IqFAzj2oVP2qcpbkuRvnuMBOXPHzAxVV3HVRkB5w8hylBJQ
mPhVeCHW769VIfhUK9JlU1inEokhO7fM/oMAs25pzZi4xIgtBQlKoP941vUHg7d/
0ieD6Xzx0YhjOK3uPjlrJnaLjGEedXnH9fId7wM54y9jHi/tRfl7ROM7lCSnOF0z
zX7dB7eubmjM8dGdWsZZZ8ggD+s70A4u1jOUBhq86HBnm+rVPxWbdqgqReS0uvca
JpiOyCPsu25l5NNNUgJfkQOViWNllJai2HKoAav93dS7n3ZoqJ8R5xlYjlYRCm2B
z5JZBVjPRZbh9vBV1WclqwDFzdMz2hWESwNPiZ61+KlCcYpBykOwHpsxZYC1Mq2e
Xt8orH2Y9s6K2vHBulTY0c4LaE1wW2GwKOp/TkxdJQpxz09GvuShOJjEImPLfzpc
99eY6RnZE6r/mwpPvVnyhibIEptPeJ3+wkyzIFCOMLSs2TawxiF1u3reIrZ3q705
D5b0Q5wtRJo8897+s+yFdUmHpp0b1aqym8A/a3cdZA3Imsn5qrs0Uf3JVgmODQFQ
mI3B9vqAlaDSE6khPsLGoQo04Yrii3Ve2VnXQnV9oLCSxP6mJ2TDZiprkAbARhpT
VxMdaQAUqRAdXrXqPCgm7OmmUo/A39rWze4sf0ex62Kog0okngaqpkMl50hYYA0z
3IbrFMWU4e4RU3Rm70lXtpiVQdnNmVWe56dfEWlNqjsGLdupoC95UOwoAlGqPsZY
yhHyP5YYy7hbT/0U00KPulo/CHY0TtAdD1EfMk348vskFlIiRk4f3HnerPhMF4P8
768E2tSu1eaONPKyYrsgeI6Adix/wSJcMGXHsmSUtFThwbyBpPvUUjn46fHDXERt
P5RzXVCX2WMi71AmUd0NCgfUzGsdbrEvdR/bv5b/qOwbde0d9WTyGw7/EUyYpu6/
xEjP6592se1zL4yggRrYZWCpf9DQ76X72hjd5c/B/+sgk2Yi9hQ8Qe/M58SqKIfY
nmoMVCU/wy4MD2VguSBo8+h0z9V2vQOHa399cUE73nQNZM0qXaJaeAQJF8jNiyvx
Tn1jxS+Fge9T1G90lYE1vKj+YPuWEvIynuW+gEfTTViNwKtfaQLi7C53u9nEGfVU
SDck8TYMnzmjNlABpp2vik1kB2/dgg8zATBSGdcUHh3AVTaXEsnwmP5/Pg9T+31b
XpgLjcEFoxRtFb74qxoXvZGOL79B2ysgkRfA0xoD1T2yIgcVO5sCle5zgNV9D/cv
hTRaWekvnWK+xIt8f5bbqbboFRctfSWzk8Es5joUgupDEHVU+2upMX5uuJlCSxg4
wuT3mvG9j6wq5nM4sawlyZTPouceHHpCr2sbznEhvCgMcuHb4ZHKhcuAX7eeqO/U
QYEsdUJLzd93rJzx6vxqP5fcAx7fDzgt/KZM5waVhT7eJW/gKqC9ZjElyPKUUFqd
ChM4WE8fHWovQfE9KDdD30162oB5M/Hi8Qswkpmem7IrDq2yCUMmdd1rezcVLB62
Pm2O5EtTdmP4Nc/iCal1btitYF6QzJpxtSEYX/2oALe4zHGyMqp7dUU/+7vhttER
vagt7ur3yUlWRX+Jj7ere5J+w76WU3FWZ/vWI2gHwR+kcdneC14u50iFoD/rw5D2
ykxrnFb2OPalsvLQeRlx8SJdkgWbaBkDZ75jHXQuhntvmBGMAQW5g15gSZKdJ9OL
HPkfVxkCtEz0tUoRvRqpVFR7JL1f3fvwnevQIbyzkzE=
`protect END_PROTECTED
