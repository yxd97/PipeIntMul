`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1dQENKk5h/XDwhhKGaS6hnyxLsHiwTC96ZUql1H89Wxicymi/B4+QlAmbW6z924n
Y/02hlAsv9pBJ2/ecwldDXTb892PTNeTt/bZDIzTHuSshjtOooXF7ZwgUlspY6TM
rTcd0OqXRE+k6uaLsv326llO+Xj/hf4MkN78K8vPcmx6nBZWrEAPx5M7MThdTNyT
xUK5NawzAgERouNXjeWmVv3em2m3M8yT2n9qqVDYWjaCbtfuKe9fzHQ27yNHJSe0
7xTbUr8OZCgnkyVsBtGMh11eht4wEFigsMrpQ49Ku1BDE5G4Nimutu/r0BXgq/Jc
o48yNNiz6TRov7e5llGL4PGlRRLxJVBKvO0ORPCuiyv3zQ+xIwFJGZTXg4fTPBjb
x/UTiaYKAuU3wDFVi/XyaQ==
`protect END_PROTECTED
