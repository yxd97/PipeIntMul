`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4HocKGADfY44Ibsb1pCiZLtWy7ZLXlP3NFx40QRLOmCYpo2d9w/+NL4LxUa7DA+2
SAcW9V/IWNCz1SZUUX1L0cp4a3IIeTkWeeCbOS/6bvDbhy4LC2BAQNmTmB7uNYwt
B5KnGG/DJA7lwcGlSJfsMtFCW3YJnIKxWA6om5GN1tfCQYQJfId/JJAyb0l3Ceno
mMZhKTho/7KTdsY9SfV+zxn2DniQJqJ/5JsH/Yg1JbEq0zM73nluknLweWwAabpj
pqGMhVjRZMXgG+AulVdhoFku75YACFPG0ggGy0g2JlW6nyx9CVTIJ9MhSCgEj9Ld
ePkGAa32b8DKi68seLK5ZW6lmW4u0wg7/E17+Ef5fgOCxmFcCaUGQFIHk5aGxGl+
lO6WeBxBQyFBhnWBVEjgntyhHTzlRnlqyGZ0+MveCTJgPLOxDUMqLF3eeU9mAn5B
u+4Rjj7tNT+qkv3XooF2xhW/MUJHsdeEGQmnoYOU05TzIJ0Fq63cLaf0hX3nHZOV
LeXcG8Z00G3Rs4KHtjaNzQIuR6cDd81t+Z+DX/ZCaU6V+ILau8Rq8oLanb2edcmt
KZ/z1hnIW5RkmI7310JPDac+GCrVnajukFeBDtX5z54LpwtuIZqAMiYe9PhHw34+
8GK5LiGVt9Qyql1yuqCvH51l2YUYgwD6dWNbTaD0stu4KPrvoxXbd61gStmjJfjH
h3jKY2Qh+PX8geqYg6Z73DhxAn1hH9ZOBYrKU+6kgUhXzQMeVgpoM/hZBoE51ja1
TdMs5D6xOeCZUHX8ay9Me3eRYLjGEhwZVV35WDS02lkL0KPj72xlN4Fh1cTfqZQI
NxvCa35Mgdndn96Q84/ITlVUK8gM6U+ol0PrNh1qesc/v/9W9XnmyREX1GoVgQni
4Dk0JyvEs/xhF2+KvPDcWkXupwYMvoepXXPBq9hHmgS9WI9sjIRs8MMspkHdixyX
20R2jc8v6AtLy3WBgKNUwEFffyx9KUfPDocPxblBnyceY+dypuiicvrhL/aq4wHF
1yECsVxspVipibkEOe2DHw==
`protect END_PROTECTED
