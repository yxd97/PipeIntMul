`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbFf8aoaGlNzleZC7irxMRwTHeINCoSrNbL05Rek3RvnLcpRN6tTfUfbDKUPciQ6
YC1Dy2o9HI3YWSuvBAEu8IRTHIxWp0XZmAkGQU0LIXnaa48BJt1HhtQb4kwBQuQz
aGKxJ4r9t26Xp4A9VDYsvx06qG91A92karG1jC+igSg6s8Qkf42B99FsS3nDMYz0
H3yr4A2PwTxcjEF4hFPaS15/NzyhbDdUunkmSERU6vsmpXqDzt8vAsYCtq74KmeP
I9+5cnh24370YPbBFfFOFC4urBIhH0yDAGhu93R5S7s+uhL2ubo1IWYOw8RixOzQ
ZJI/Uo93twfE8bcem6khpQgOtmLU0oED2hHKDt1SA+omSAGiDulriD05t5elXDBC
JVdfA3tZgCay4eyiKnbeBFXGDYLewmthmfQsTowo+OZQ/83fTZjx5uUL4Mz7k2+O
HS1lI/Z8gMm8kLZHyWP+PqPvxyUjR8mhq9sy98RhDyCoxN6xJOlOW4T4DPABwETX
G9cw2txgB/ltmnL2D6u1TRPqDmIq30e/K9fQ5zUHEcbKhtbOCMBdyP+CA8RDdcnN
2/o0BdG2ztwtpTF5hfA/Q95QNji7GdunhecjOk9OIR0pbT5oEOhXaMV92Zho7/SM
9W6/cTEvtIzh8KBhRmq6ofxwavJWOgBXp4uUDE9WfjcRmggNcAogX2WMmWKTwCe8
4l+76XILXBwXV6mhv64n5wjw+anlW1d4ZJF0C9cSg7uv97bbghPHlGv8u81Ru/Q7
G06KIZmK736JWI98ClRHYqxsCna2vU1jhYOyDKliOZHH7Scujo8h5TNqAEtbzBPi
`protect END_PROTECTED
