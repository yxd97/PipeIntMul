`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tcc6wl3r9o3zlWgsspKdtQ94n7ieh/XpP6P0E+62v9ySV04R1N0g5BQdSvq0pB3C
kHMbxvQeqPdXzdQ1M8OjcjdabkocQPy/dm30kmWFGCfV/U4pNQpixZa4XZ58HPFl
Fxy0IrUd3ve8arOPZplGB6HndGpe68puxAfJbx2lzKMVXkuL0AOdt8OhDrPpkrlG
mybduXtROkMRtg3elrZDSiE+1hhLRcuKAJkiWedUfsXV0S1xbMmXNr5uxn77UAHK
O93i49jvlGD+cr7cZvB+aZpWRBHRO0ESJOSo5RRSqsVLPmTMMVLSgwISbtXGylN5
40VCWUaQgpJ0+iUydk2RTJAhZaxgQ3tUoPIKD8cPTcKwEIh/EesevBk4WkAuOvt5
mIfwTd9Xcntst4KrvGxaWJJSuozUFBFQCA3ic0X2kTtuGiEt0kpJCmlmLaAqQP8m
G0ebK4rSAuWOlMh1pxmIis1j+1x0vXngmGuJzh89VOQFlDvpey5HF1TZuxaCzp69
2+O3Qj6RU8DLt8y9mwmDF8LMoy86QZUDgQT8sG4lSKElBuv89FratBAFtrhTtNM/
4zs04TImFk1MFSGJ8W0x4DB1XoQJtuMItny8HnUYFvumzx93zTAA5hhlsNfvQi4B
oM4RNc0SLF/3vT+6hjkhzXCF8i4LSLatSjTy+6vbMh0RbF32UN0NIitLO9dnY/fG
SClgHvgYAQLc9Y/Heg7E7+kjHlGk7+Pu61uHvVtkQ1J6hS0sshJ2GGuY0uWD6tF4
xh1NlpV7bOsen/cUThiSbrehLkxGD1Hb4tNW5mGJEAlNKljJV04gm+wZcn6RoPP3
nTRoZ4lN4H1dfcdq+32K26vJXGdc8UQ7itnh71r+mkAIOVqH3yVE920cGClfKJld
wNMpVdYIgerxDwRLtpgA3bd9uzJlYnlQn6v/uypUztFbgcu5nHNYiZEyJqB5gg3I
YABj2QhtHaeo4+ZwQ5ROhLoS+V6RpwnKXwADVePNpIGXi+hiD/GvLRXFIxApurtm
/EjkZf271zRRysLNTH3/M00lSRviI07n7VL2KmuKI1ZxqZEZNlYtxVCdCMZHTB1e
/SJTfe7KcHrpg38VMUMchEeRi5OdKlEi+VyHRmVlw9NrjeirV83bpNS2AkgizDPx
/0btIg5Ufi3RhtN0tnBagaRiZqkjXwEvEiw1v6Ep6CPVAZZ/+vRFTqrkfdzErDAg
/qap3LXtACtiPK58cL3WlXgjPKY8fRqiFBOks2FVlFN6UpKONdr+z54ao6xvPY2R
v19ac6GKwZv2WaFs+UQVZSB0vN6pi2dVgYxDdcT/Dy05s1yT5V0E7A/iw2fFQcTH
/1imWT1n1jPcLvTCuu7j/b8MOpZJHaWpkXRyWgADBrqTi/kUo5GRV+E4mjBLryxt
QETg5/XHDbAQeBW0CtLJrOQFZ2rOSPZNMg4GZWWFUN+7KV9FFfwKq5GrzMGOZHBE
poq4SI8QumtnnJPK0ClwbWPiodC0qRjBbDGhROWiacsGJ5ffYKOLhuXg7fzMsJJV
7IqtA0Qcaczcy9jkpY+qjDnlqIBmvp38RE5igzPJ8dTm7P0G98rCHDo3nZMnsgGk
K3QNMGtURFwoJpRCUAZsB5I9pxh48KCd22wdgGHBpvjf3veVx5MEwTmb+3U0sZHl
Ih7rLKU1YnTLQKL54ElNFADBqu13eJNZMvIHaHEqh3EXfAtuAptnEY8oAvjoAyZB
3qrxz2aIPIB6HvstXRZ3GPpM5NNrzM51KMJe8yg0r6o+iNJ6uyH1sqzAiqcJVyI3
11xlaMi4959BuMBGqL+0uKflABcLRNThUrBIa9IYBH2Kp+XGSU5/MaNdvIVCzN9r
MP9ghILoaviOED01RnvMniDVpmuStrsqkjnzU/zTJm5p0BhWFbbbZsN7uW+vtsuD
opOHZ8pHYWFcJTGqDxW2VZNBJs6uKNCceaml3PMBL2sAAJdFsdijVWlvH0MY3SQh
NJVG/jGO69WTbHXgrImhy7+gy8Ib5FLKSWMixsmzAIGVF7nRjbthPkho4/E/vJG6
Bi8Y2wPQWyvPk8ulisncuwq9cueDW4BQqQ6A8LbqdXGxSKZ61weP3RbuFt1ZC83I
VFCCNwwZJCNo+3gCPOtkYgb0VeL7pjxJsSQNMyxjfHKwoFPSJ1IJZqiNvw9r5/Rb
0wEi5CZmWLJjqPoQiXck2EO89KaxpnHn4gYYSiraCzbEPY+Fjfd0jdLjWzKZto8o
YMemHDFTXUw/c5NYItNv52/mpdIB5GhSRiL5kiBBaSyQhIVqhmDvgedByFLXK3h/
iv+IVNSsBHOqnat39oVMnoEIyJ/ylkiNU76cYS4OaIWuNep4Z535ZS65jfbQPF+H
8YWefLYcmy8q5KkYeUL1DGEMuBFaVEsdJ5hQfNjlZFw6s+fpDhAxKdjgAUbqnSTT
jKQetUJB+VCfiaCdNsitiGdYKng33L6E/hj7FWdqDw9N2pUCCLPAS20ruFf0zqUu
xo+1wixgG7ZWyBoRQewzL4Zyw6lgYVAudMUYWvzOwaLD3QnvPCo70PSBx0pUHoto
e0ncMEOtvX5x4CjbBRWcsyCWiHcx31mo/B8veDj4Ik3YPrY5mwcg1qaoHIoB90rs
xUzs3BTE5+R9YAQ7x1mGtWKh5q5uZAkct/rTxp1V3r61MeJFeH6Hhzj4Y8LcKj9C
dmOXB9fW+ckVR5/7qAyLvRiZtu6wO1bWT0IzLqcp6TcgZf7zp40jQftBDukWPTJI
fHxdvpAiMkvekmMKpvWWubekKtwN1Edfy3I6Kfx1NMRVusDDr8ylvZGZYsnqXuOr
jBVHXajnQ1tYp9y+tI9tceI+PyVCMuhHQ3SlJq29w2KgjBEBJw8p9ZkfPH3Mx6bf
/1qcMR5kDZkiKYXAPYgmAiNTEd/Bu5z4NcjNUyeF7QRBVzlhw12eOwmjAEmPIfu3
s72eYPWCAP0VkTUQYOmnXZTKTs0JBvKC9FSucdqyunEIOgwjCOmm9lHOYVwdn0MW
gGNiZhWOh9lHpSlNvABthOtQset612V4s1ts3thlq7nVeMAOGdUyrScKda/Y1wJK
15xkrnZSKxzgLJ6LgHRbIAYgxuzaJw+YbOMQ3MYXKe9fIi4u5lKX8mAup8+AI18I
INP6FTPJhi/Ix49otcegEp9IccHk1v0TCU7oiTgMXuqwmrPLd/L8vC8GjC/KPn8l
T9deJZLidR/SsswajoTHfoN6e/6SqGJruR8w9bp/6K4d2rbsokAHkGSVI0wz418f
+eR5yQIardljwqldgZPLk8wgptC9jiR1RoRc5zCDlQZaafV1S7yaJdZz8rBLjvKy
LdDTIaguNBS878OAPdPBlGlOjiacmCrtoonx6yhEJtYk8dmFPYpfN9LrUIIWyO1d
S54Oi3NFCG85s2sQ6P8c5MpPoysX2O9RAC5/7ENonRAt6Tp/r23aamfW0oKxIuAo
ULO7WxoQzXsmvbCwk75u/7dZDbFxKb1qCwkjN28BbbTMqn8eSCwhFORbGPHft+y9
rSJ93iIH4cmM3gV5pykhvYJz0HYzEnZcf773dQxXfdDc1ijmcbrZxXQMmXebpiSv
zRSQIB1GwUzfBzdiVooGjUw1aEw4+CR0nU6KNCRboB439HCgAQh7TUaJE2pdTGK+
3XLIn72uzYVy5WsqacF995hhn79jWYdWFytj0HNUWbxXI2Gg8wv75O8WJr6kxJWh
BAUVNabYRMd+exaGLRWl/c/3e9XrP0Hndnk65Ju92hXR5at6pi978CxtDvUttsOe
yReCKGtFGctHUJgrHRvpzGLp9/t3svQuvX9tY8jZ/zBqxvmPHhaO92rU+5q61gRY
Df+71Se/2kGQEPFHNUGqcYQdObjadvgj9xNmykJ5lQ/hOOF02JFSp+vPZ95ovyk4
z0P7wyIU8fAzZjr6TVNwInUpihoz66ITeJTCnnnvJRwWdNyMs4tKF1BTJuiYwHKJ
jzQ+CYpEAAS5vrPptBHrXzt5GQA7I5YMS7JRi3AyxRv+8g27r8BRJCEUWjOVr3MH
C2J/cVNJDL+vYCD/YiiqjhCxycXbz8htzKaCobHh3qjRZLQHE8Tx2WGn9oVT20eR
jJzO4JKmROUK2KMZyypmkfr2PpheddIFu/5dRxkGVguvBbM0ejda2odmQCnB6ktv
kYEel0FiCFcWpYwJiAcHxKuZX7vNjUz9HRQQL5xH9Y4/fgBc3JmeHwEneR9cdCCJ
lTmqIgIYEYvDYjO7XuazwoVZFe3XeawPm1zw63XYmCiaMY2xgp5Y2rnSe/Ok49ax
q2qO3nREMKk3SiMDiOXnd9aUqqz9eKaCIo4n7Jq24D1eIgIuOst8h2dcanG8aAqy
Wasjpg5GTnQNVYOzUvLaZsNORsDF9A7Cy71zRaaXi64OPw7qA++JNPk+v3NozWVC
yS2IPjvTXo4RoZAF1TEhrrAWPbe1t473uejqxnXNrWPvc8RQ8/pYts+Ik4goz1V8
7/CJvHu/BDlWtV1tqdEoa7Q3QXmBn3+eRbE3wM9Gw+cSda017HAVMog+NVAr5tzI
079iW4T1Gbfa5G9iM1alxCyAKdd0mg2CaNRRReGfcHc4kaojGF1J683oGFdBk3Yx
SBmnsd3mIa4e8ghyjyAqFfOXyWVYxs0yeloAiO6igwKQV7/Gl//fOS6LDC1ADKQc
mQXPWEx+SfSEAk/1V5gSBw==
`protect END_PROTECTED
