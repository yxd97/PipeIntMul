`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EuvpXLWosGqvecD3ccwb+ncZvAS44aNTrZo++ljKVEetpCsmEsFVIchopSPW+5mW
BUDlvGrcV+9Q+W2IGgE9zBIjevVVP+bcVQ0iH3Lcfged7d1J7xIyou7tWSSd9idd
y3mLBWBfJ7+1dnicVlvX930d3/oPhFjPF/rbu+4spvIBT3h+zwAj3XWXwQGJ2uDT
wfMz4Ym0WHP8MzJnk4SeVcXc+HqfdZWIMPRTp9KhE7rkNlaX/xirjOY5eV0zOiTU
0SDLqE0XZbzDJHpF7x6AvbIB/g7LondU0E3WvryBeLyJu+lo3/W4S8Ca99rBRTcR
qAimZ+5mAwacQ1iLwxhcetJItlnCxJZNbIdkSMOaejdjMY/ClVBJWS7P7W9z7bO+
KEHyACOkUW/I9JmpNTrMKQ==
`protect END_PROTECTED
