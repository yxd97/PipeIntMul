`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kUNDBy71XqgNKfB5iMtrOv0Xy2iJQcYhdNcl1v35OQ9FFKWGPLRw5y7NW72i5N1o
FNPe4tqrv5H1jTkUgHh74haiHGtEGfDbWhbK1TsqaTSL1snMwsS1eHMycgAPJbMW
DLSQAEzcPNLde/tCV4LEgBipYObbJAU73He/67QdQNj8ohWfyq8fkAr4N8/KdaKB
+2JkJbVPLejCe/YRqxvUavpRS7fLDppPcV573ZCAF+LJPZaxDL1rMJeGR9roBPjy
GvVzfmlwswsCFzuDo8pRbPjAtNsiemdwkBqkj6+EJQqNBQTvc+bV4d5E4I8kGV60
Kxa5tMWbbTPpEAmsFmZ55dqSZZU1sUOzDheKx0HoR11l010RzvTDLnMUfMcr6yW/
9GeBrKSV2KvnR9qPMfDCudrJdfzV7WO+JYjtSXY1wF03E3v8HFd4v23ldmq8KeYI
zmDnp+VOovxqeLmlIwmuGaTpl55uEuqFcWrnKQLV2Og=
`protect END_PROTECTED
