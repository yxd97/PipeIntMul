`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xA7ekBKvb3wl9uA4LhYXQOCBTzID2yN/H3jlJtoK1Bx+XcFwlehAWYjsWJj4OCaK
Moodelx+nis5IuivCOCCD1ytp1yS8ITpH7uc+bUi+0IgToUACPKSFwiYQwAPaPeG
XNumeFOF0bwHrnr2tyDZyKRb/+BpkDUxZHxrVvlBhrSlOIX9xqPZJ1DASzITs8db
+VaD6wn36qr4zkMiW3qZBSEThXrUq6VWJ+O4RftKUYGmxGcSACXAlw1FdPw4y0VC
biynRQn3Lpib0EsQrYemr6yCDa0zKg48lFA1ukJkJhChMYlQZixYDkzfWFHxwY8e
Fgr1G3VhVgjgYUibblV7XPCrtXF5OOlsKL9rcJGECPX+UBMBq8KhUMNUXp+doUXm
kkibKoBkLz6wNQrFWsQgaw==
`protect END_PROTECTED
