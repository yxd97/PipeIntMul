`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mubiU+/hcKNkZz90roVnov4GPczsHaSdUMq3gF32QPFRAsAXMqvaDe9R3rbnJYss
fzOcQ/fzl7PFncjzJ1MieCeehTVwWV7DJbAOmBrHjEDcIzul7kRlJt+oqEWqv71K
WMlMfwnNjgmL95KY2z4Q0KmvWhSxSE2EXXfGYcenaE4zWDAeHMG+ZQFn1HqdzvTY
OSMFE1HTQ60Tu8csaDaFTL5AVaNxB7WR8PFOgynZ8yvyGjes3av16777UAkM1Z6X
Wno9oIyWtWcwOyF5CKT6ZCwt7jpi7kEbsHv6m39BaA4=
`protect END_PROTECTED
