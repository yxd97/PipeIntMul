`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T8Qw2sMd1m52UD2Pu7i/jrmQWniuOcj8ojqW4mbetvLB+McZ78ZJBlAZyQqvFGpX
IZbxhaw+TYn96O37AUzNdcxlDP1/8bxzjAeqNOs5Rbp3i8IslrIz8LHz+NBuSrAv
9HPPN+bLgUYdW8yG/K4oVbOIq/PTySE7+9EZLBcKCUXNApAxvU+EuHC5WehaxLEG
ULz04u+Xl8ajfHzHtNG/OVIr+dPkh75ejOJ+JoYUsAp5wZHgr0ri/QVxlcPrsiAI
h2Nov+Tqne+F8JxSEpt/EgJ3Y60vi1kxP0gVGVDw+LbHGA8ppUdLfQYUJp0FDJTK
JHG40Fz0+Luj3V1Q+3SY2ME9cXD1MLlHBziou9JX21bsIXk6jp4M9dcytyir/AED
LL9l5PB0AxOkdO2O+WNRSaYnMScCt/qHm9yQR6Z25SGFo3uSb4yFAWKvytuy+mtt
`protect END_PROTECTED
