`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yk3QrY7MgZTFhOVV+EfcE4gEDc7tJBUNJZjew8BAci2m990tArqJP+h/TsBcIA55
1E/WW3bnVRMPTs81BSbuKv8ajWhPvQprt70Wzifi7z1JsylGSJ+eRb9Ct+enJuhc
lNb3iqxdvu1QlgcfGoS2Tesktsk2JZsQB9l31E81vuFn7TE7SL1y5lKYNmK+cfz3
oDJJkg09Z/l7hzN43zOF6Zd8NSYQoSIQPXbvnMxbbA+7k/LOzEMvj0ibIl7WLZOq
zJt73P363mq1Lm+qoX/auHF/Txm+9iXXirC5k4mpFm3z8MwdRHSpsQFs1qi9HSvu
4ueRahetKDuCTsUskQj/+XMlh93J7QR+MhNEFWm7OXI4V1REtL6UkmVOZZdC2WuS
4xtVkLJEW/XMoMvo7PzoOm7UH/RUQ3fwocdQr4XTSKSyV3aZhvkEwmz9GQjyytRL
22En8GmoAba2KR3LzysqcH0YHyahhFcDXxDLnmNMZdPzUi28x2CQ3ixMM6Ygr+t7
0XKPTNA3f8Gflqms4E2QIffwoj4v2OgD6Qr4cUTMNprf+PT1AjnPoapIYDsozrpV
8R8TuOyqKuH1BeP9Ge4YPl2EvoFuJMTZIaTDjWYVugOPvQJuZjf3rbRL2YXIPV3k
8bQSeSZEB1oPwrNfEMhCIWvMuEJ/cIBagctrKzIn3sF2uNpzFTjglT2n6Ix0+oj5
`protect END_PROTECTED
