`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F8F7CqvnWpBK4OzY2OBQVaBTMGAYyv/94wEJUbIS63GhjHFp3WvyABmsmKzFZ/PF
5bNkjVdn5aD5VdzG3Mx8NCRt0T/yWIfe1VQlcKakXxgdBsko6JCPWGSjdqCaSAtt
yYlq/NP7emErJcaUEErtgvy/TJjLXgUGR8M/einuIwELqVPVNGTikkuo8fX/9fwO
/43kuq7Vt6Tcas2R7S1bXo07Lc8WFrEx8gLjuRbcp33i8gl3jKoo/Eextud5daiN
RQW5OBgYlbO4zp/84bi4s/f3TNIuKchImbMrZRu8zsVaBCEaAZ8DdRHrdrodSDJH
aQ5vfxBMuUYEGwyN2sMaoQbQ2Bl3LtHF4LAX87vJMVYqANag+M60PambrCkFRo1y
JJyv7gkpLkJwhKCTqq9WDO5KNoo4QAWxP123elxRpkswfILdf0bVAtFM8ps7rYg7
39wzpVeaqFU/yFX01WPiVUrREr3eD4Qon18jMmICMYQQ01gWyAvEgVI1Ba8MiU4b
PWH9zKWmpI4ohE42Y8B4TLMqIZcW8yZPHdoGA9y7H65Y4wDBTinxfiAVT9lyFsmG
YvSE3+Y9JLk0m2sJhXmCSbz2QmsD7OrFGRAQMs7wpvBfjyoBpw535qPRAfgA48nw
u9rMap0um5wM2to30O2xBWbqmP7a9f4evPbRLdkt9IFx+kxGAi8BoHTZCwqKbZo2
eIoIp91ZrGSiAHEv4vsflaOitHh0cGfoB+Z5TbWDgVU8xMpx/1lIcy1mgTBwzWpy
RbhrETtzPbgd72cORNdHgv/DT/jM0Oin0pK98HOC56jyVWVNtNTukY0aJUKWHsZm
9h9KmrzR677yRYLr2IIRyCHezEguFTLtPb38JtEPfegYR8ttcxRgLWilzX6NhMHi
W4gOgdLCMoGUQvmaQQ4Z6jJOY9hDycUUGHF78zQLTB6FWIYoCiyfBZPUaucIpnz+
pn6rylGdQIi1tZ+eWnlrnIUPvDsTgaV78TENxTqDl1U2cIdf9KSFOChohDxl+u7C
v+LuJoaqJGEuL039AbvpaQrXk7Sq+XJr2ULNj2xeDEdUl1GlH5SajVHWQaWUX+Qg
dWNNZHVjEscjh8trWRnFGOYyOoCEFt13ZeI9h8JMlkoPZP42ouABZtVHlxDxhQrJ
QxMLbQ2ucBsSSdxI74409HuL6trsDpjkn4XZ6nVX5JKqFnTgCGz6pfmNv7C5zvJl
o9PnX5utP8KEh1KljeHGYfoQY6dC2vzY9keQIxc5wQRxUfDo7pq2gSwqJwbSp4q+
iJ5lzy04r1Ji1S7JD095Zlnw/D/2K2O1aVM2z1o8hDqI+KwGJHYFlasxMMcARpBA
pTt/PsNsAOq90h0axcY0LDYstOofIXuou04M2qrJPuZ7KfwhgDc/0mtyFabsdWoK
Q6jS2obHHgTMIsdi/YMFs3T2olpAWra8xBf1BSO3Y+EeXHZzLPnyEiT+/RYMLKtI
mL67kPzIJdhO41TeS/gsGQ==
`protect END_PROTECTED
