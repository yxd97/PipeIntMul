`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/NZ92RX/b/pnz4tvVlShFRPhsp6+jTG3uHt24dkgNQzZYbHp6Io1oeOcB+gwoAU
jo0WQ4yk5ndznN/vOLo5sxtZJ6ZFSTbIBLTWxId/42nsZD8c0zR9yUlRjnJWyh88
QWIkPJxLR0aC2030cssRo8Bb23KvQEA5NP0Cn8G4UKfFv2eIb6m5ITwROFMFRrLl
Ss+DggLGdRQYPHN+i4js9UdW4yAt8w2+HDEfzKESV35VDXbKeytD8ppGBsCeSorQ
N0YDnTTsMo0Z8avQyRBIRhBPl1hhfoOjLmDGUux3qUkLCPppMxmlA+vKOKzrx+Od
WmgGcuPItfE0Gqj4wL8nXGZnCUONoq2NdBmLFAGa1Ze1CuHiSYS78A8c3gsHBbwo
poO2JnuG4Acl9ZsIiEPZyQl97IYctrX2tBQecTlHIcgjXC53k+DeI2JuP9i9VNFn
1e1cGBMbAf6Sm7vNKxmmDQ==
`protect END_PROTECTED
