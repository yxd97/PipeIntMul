`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OT4YzyS+xugFtveQwjSPCyGSN0cR5tIj+m7w8MBCrcd9vlB5t3FXVawu0WJ1vahw
sZKg38gkQUl3jy31WJk3Du1HGhz87Ei4QvaFVupC28wK7pTG1wMbMNs2lWisrgCK
dU/KBrpQVjSqF80I0iItJmlGOmhup6Or0FZd0hpJn0NbIj5oInW+0Y7Jt9WOV291
YsvLIsDcLFHhddijkI42sk0RexdvuI0jXQLetbrHK6mts/82Jtht/b0l5dcChZX7
GHk0cWfX099cB3uAZ5EWXGH966HH+Prv+JRD+DNnGySnWaeBx3LWlG0JD3Kbz11x
k4SrVDIfXmJptqCu4YTmJQRz2GzthYxRwjKMJh/9Q1YIdtFzsGZiGvsdVxQmOFgH
votfS2CfXKOSPocQKBP097eAeAtTdTob74J7frk/OLvI41xX5HQ6dK+rEVvDI8vg
fefPmrvwpMq82m81UfxJvtFxLAOXonhL/LvmNktPukqygYRJ6ErrTMu2Ow6vWN0x
8FtglsQYGx/Z524tQh5yz9+mAtgz3FSpmOFOS50AodqGWgYhtQ4bqIb5gl58Bs7c
cs/IpGKJ+O4bA9fxK89MjXVquiTNI+TRyOshX8TkzuGVNloF27Ynwm8iy1Vd0ERk
EBpCT+QZBqXIND5XQ3tvUlvHm2abmgxoreZDFjGmqRWV8r5IbgKBoTrtOO6avG5r
`protect END_PROTECTED
