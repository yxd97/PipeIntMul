`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Onah2DD67DpDCLqW1BDFLKD8e1NW/5RqTImWxDA2h3MBSaXILaREScwSdeDBPJmg
cAr+3jZrZnzeAyScuSnubQ6yjXf4H/vwpCB6tGszBucyJ12ACUNju8IML/wv3erm
P6pkBOeZLvK9pNl7/GIZKx76A9a58INaFyjV8O2wcmgfd6TXbajytLNZEqbj+ao3
IuQxbZPrhFyeRNdaICwLALmfC4vCphDlwlb26i0WsVKq0k3SzhrjrTi5lIPj3AYy
Jsc7U4larEWQaiG3SJS++g==
`protect END_PROTECTED
