`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QHTlRsGC1VGYWMgTxTaU/AGfHzaGGZ7m77guMoHWn4au1t9xjEB5Kcm6OynH8S4b
6G9Q3SU93EVndwW5bTkE6talKwvjUD3IyuEAZqWryEwTCRV7FtoEa4HqvN6X8YRf
EcoctKXIeKu109C9nBKMU9ruur3Rwrd1GThm1Qmyorb6ONAeE3v059TseFgNyapU
9VldKl3jcglIF3miQ5bzelsP1GiKLeVjT701Q64bZnp6l0z3k4X7WSIZatMO2hWE
f8s1b5palfL2m7IBQacGl/MBYwAkiVbYh0AVXZB/wkr1lBcz3BVambupNgR8y2Xf
vv0/8Fc/njUUmgmdy7/enXZ9GeDET9BDhEKlLjRI06SYGSC22074V+OhUvMMv3tD
LqMyxQw1TEVyGS7v5WmhPLEkQxT09h5kdC3a+VMP6zyxdOjTv2tA1wqVa8zbayPS
vplf528zVmhQ/xU9LA0mf8Jq24rdta2sEkeUNCf14ao=
`protect END_PROTECTED
