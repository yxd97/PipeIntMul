`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ls4HYfRNgraZozOJmrGs7MkhYPBl1b4uYQY2wh2rq5tkrqV3lMGAQ+HbGBOrSVYc
dkLxdltw2PDGKeojmVOsBY1RCzOl3XhsZvIUXAi5NwFFsLmTbC995XwU++qi1d6h
9UXpE55UqGqysGk+lMgILVz0mrk49R/Ul1CIFZnMMDBEhCPdv/iMAxyEyh3+6vtG
spi3A+jnBJGSWgTsMbtnYNhzwQ5sVRIO3q2qUGF8KEhNivQ5ITQZZ8rbZ7dHaq7r
cWptsdZ6KbUpv2sFzXKm2bHVfC+3pmVkf6EEweO1U+inUfpoJqqIxMjwDc7qLaYS
qQtE4PVOFLDQrFRllL4jRHH+GH2oPN5pPdJWSjbIbAyG+TlapLAhKSBDJe1/MZbW
HB/k10ALHcj7Y95HI7gEtA==
`protect END_PROTECTED
