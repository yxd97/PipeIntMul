`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0M40eUSQUqPMgdaOuVPgw6jYgtE/mLGmCPKvMCltMevIo2KesPU5FipWlFcpdWLE
k93xpeREyA4Z8NDO3K3TWegOO5g+7mdL5aFlcCamZdfAi8l99Y1x3ZW/lyUeMHJ6
OeqZru2EdHoqmaTHLZ38M/b9kpJGGNWBkfr9C7bP3f4Ov4BDGvoWUGBChODhM3+F
3LDSLTV1sQCfqmG1dN7gEcSm2+F9LypX7KVraHV3/WVQYw9dNHwaVBTfupqocJ3R
TIaIgY61dlSuIiE29jnraWUDwX1JyWacJ6N2rsBeAfW1z9HrAMvSxGPBJgIhBp5x
V8vee/T/51jgCAgNIN7R7w==
`protect END_PROTECTED
