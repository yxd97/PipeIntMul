`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhSKarZB8bDF2AZVg41V/qo9sizxZDyKe+1CM24Gw9zMtwum0hT2zB6ZZo5EhYgi
uG3p+AN7/n54lN6jEUO9AYlm9zJ+z7P0HHmeXdM+Cq0V3OvnlIxvxIifYhsUE055
f4zgt6ic5TfRvz14lKJAIAK1gAqgmnMwXLRrwm0RcJ6IPI44Ie6JDL6/k/+WSGbX
QIkhQJgo4KSBrSWxt9ggdZ5DHgamsod34Xe8VjpglQfjzG3LtPEA4c+pG4hWObDg
RszQIpiGaYK3c3jyrGfrJO75/c0J2TMONQuyX8DqztmLIY99BvxJ8gUw1tQ0PWhB
UrrKJWiobSZE6HkNLdwCEN4Snn6eIT80X7OcD8QrKD0KNQ0ToOxT21CgOnC+EmgW
tyP49QqTpDqbpxZZCM1QsUqR2WUs3k7zHHENpFkR2WhhTlngr4vcBMSP0DTmJoqa
XA53skaFaC+xKWsD1VPgJ5NP6OiOhoDIZxRWQtC4eMjbLNxjCckE+JHeuMVV8Nfp
vsAqh/kbeGpfM9dONgZmN/qjP49iFuxI1v5LLaobEPrYLiJ1sue7qHl+WmY8sPxJ
Mg0aU6V6kEaRxA5CatNfvJR5B8sNaAI5Yu3KCEZJepT9AGuYcITFGjlNSQYA8aoI
NkFL0HtcOOkWKmzJ5GAzhJS4UAinov+5yVDacKjcbLugf7wVceHEa3lTonsj5rRd
VI/pccM7M8Tf4inRJwAt86kDXms42uDH0OmrYOaYe2oJVm+i92Wbz9Ef3C/65U4y
DGe0JZeEvkxxw4k9d3AT1Gp6qdw4jReZRR+6EhM/76J8E1Q3uf5f/lmntN0PPs3b
jkzlDOJbB/B4o27/W60LSMwsj38uCfzblIuWf6x2hhEbmljtU5H0GQvIPuuS5Kk/
SDrCnToc99iTjO1RIbEQTfjL+td9xihWmPzIx3vgEJamhHt4bfBwSFR2coWamUtJ
PWsnK5MjBOqYgWQXe3KjdfyB0asIMbrVSFLU7qaaEaGVrfPPNl5Msc6TVujggzcN
qxlOqRMgEt3GK/01VXe81eGq2gF6ftcB4eEMBKq2TufIv2mSF4jFcZ4F3v52RW8v
PdvWRVyGf2ih89Q04+rEUJmdAXyYLzrtxHZ2ELNUeYrWdrgKzLYL8MeoY4XekTNr
GV8yg2isZowL28SDcqvz4d5y9rWq13k69/pMslg92dIuXIfiXqdPAh79FcJjHRBu
VzacDCNUM1xp5Mc6D46ifLjkL8UWR9LoSu0Q9ACqUaaPS4vwzr14ukmFFcIxH/by
YYxuo5OMK2JwRJa4Uq70Ks4nc09YVRNgiiMzhPsqxG9rkQMhNyBp2lL2P0i//IDN
EfsllzOTgX1A6xPlsCv84edg1Xy69P83Je/xaoD7RpkZhC8uD6m9NdUZ/Gwi5yOe
seSJ4Dc5ow3F40p/5J1/mqVKo4JeOlH0wJ+KNuqE0+d+8f+XVNvLpmIUGbGig2WZ
xel4GDC8qepVq5QgZXvuuzoVHDoeb3HxqldzyjFyXDDvnvryKj3nVp0ZkHa+AWaN
BRnodl0dcobEjQMtTJNdqy6MgihwCOSZ8dAVUapRpmPepG/BynNTixrammFhuPSy
QxRPuLkQOeMPdm6OuM7tc7Ne+YYicEmndqzYEZuYrt4LqSJbzeZY31whG8odw2Lp
uvcXGKiAjdcsEPxM4Jtm5PFjP3zoJhNIp4EpcGWgC3t9OaWf3QslSaLpim9mFHHk
lkfb45ooGkLO0EBtO1I1bzftfOqb2/cbzCqJKc4t5I7oi9E0h7Ew4GAwzpI9hKoP
K3tpac0Uxa1AL4X/itNN5hhLyc4HfglTdDRuiJxIr8fOjlQ5vaLFL3uagN5JYVhg
ZfkXsuY8rNKERMDj4gCZvvEg94fXKSYvlT3M7Y2GQTzLIVYGB2xFCCFa8NRXw/Dk
CLPPJlb/QUH0Blz2LfQXOIAEVOHy+dVThMzFtuCJILaHZmGZbguzitPFDntFdVj8
TUnPLoXqSV8l13INMWYmqk6fcxRV24lBXKWlXZcMTMyKbXfNwmvsawDp59OxLiS+
ym35NG46IWoOR0tCbJsI6HKT9669qN5TfIBbdm/SYbvVYwXOyKwNSLZz5hzZ7HnS
Bbxj63MiuuJmUqDBnuS8vyi+PsyntoMnFKStwSX0lhbjveSw/+VDO9oRr8UAeKZ2
mF2VPOu/KXArjKwCIc2zSh/qhaNHNDldC4wwBzk5BzvP+ijL/rzBWuuTTfJlTtBl
YHSk5I78uMWX6fQmFzT/Dc+RiCITMH+1oJkmFsEdniZXXPYIlTZ1U10x55LUnGej
LEP/BZ5LBSBmRGkio5GD8oHx+J+lrAOEVAUVWNTis3lMFKcW21yjdsYFipNT3r0k
0cqv0hGHLkTcu46wsTCZzYwDb/9twzg9nphYrGbRMzDflUuv7pNX8cUvaE1L1voc
jKihzr8msznyAJP+Tj28y+4g3jAtO6ukvgcQh+OHKzEB3l6Z4KYnIqdH7YlGnNjn
1CtWT0GH3QMCnaG3GWnkUf1X/0u6DkQrgVYjToXoiTbkyNTSoQPBcjwW+37XOtaK
l6suk/admTGSBjGbpU9teBDIWrO/lTXsDQh/U8WUKvkJ1ZChPWjSGXL/o9VXSB6U
CC6TmuJ4WJLsxtDh1CEdtEJlzHKhcTfGGb9owd0v76rUmLxp7daJXGItEkvf47NY
ky5Ck8DVrgaiiUEiXP/wsT2KZXpjsVlCQwaznwkJw/TssGfdJeF5FG2LOFQeEd06
pwKqWredTfGpX6KQiRuJ/+dmQSiXCkQwwWUWOkj5hgCZnIqjqR46TPlzzHcDuiDp
TtMmOnUTDS+n6FwNnn9Qk1xsNROefft4b996knYQ8EZhLwPsCRb+AK6dsjvW28F5
2gPd7WocQ8cbQPdDUD0fuuyIWQl41AgVqTJm1LTYiOlLWYnmMH/y447+PyCYvKTO
`protect END_PROTECTED
