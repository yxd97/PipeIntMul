`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ms5p7PymVcizhMMZmz3hJrcyfA6Nz7N8snqcsd+QFGjjorpZFda7P47YzlIyyh56
ljOV+gziuJniaQeR9HWyFjcKraXb53faNv2sD1nmtOF8KMjCm1rgXvAvPG4guPKL
jGqGcjChVspjgbU/rJVjqAXEyHYxdbswj3L/ULeqzQeSSfgTn00hAQwI9VNptFBS
3WEP6s9XRSASyCTgdP6TYHsKm0pk8LXr2EQAY2X2kUTvzHCs9Lbm5N7DsnqT2iSQ
IYYpwE87e7hCXtly7KggG0WueXKwDKNBMqZVUUuk1f/im++50DL5Nx1Bbw6jpXh/
oLy3xJB8AqZSaLZurVbxMtklcRjZuhRTrQvyq/yFHTO5DXTLTGSsz/FgFhP6mI9d
+OT3vhCqnkBWQ9liqKakYvgnk89awPbQKJJyQrM7XAZOq0wucXGIrj/P1vrvdDvb
vnNVIud8Qrsun+OHnrHhTXKL9ziKZpSPUDjdKNrNYOZ8gB+1RISQROrob7m08ODq
ZQ96pVZeNR5cjUvsJ8LTHXGYoriwUDHKyeMZYkW580tI2sD1jPtQC7JFgIymOmMe
yA0LFHQpHto82Cjj3Jc8+7K1h9nAze40bmTUCv9jogswXks4pf4vFD2MUThw++VJ
aq6/TyYrGhvVaKIxnBRhLJn39d2POMfjT8Wl7Tt2IkE=
`protect END_PROTECTED
