`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUEmDkc3CqEb8qBz6ojcq3pqEvDbrqSjskZnHV1UtlHJ5tSwOgf66pEsRfaWaCXV
UAuArvz1VqiZKuzbI1g3TfpWnZciwFiihd84Csdzl9arQNfghmmEUkwMMU46N3fx
bpakOcNY1svOLUO6ian1mXnz/DSJVrEJS8kMH5vWY2gDo+ArGKmpQIwMLpnBp+6J
RAGRbxUi1JCai0l6PM3pS8havgDxq75EOKaSVKQTQnqW2yGE+nKar3q8LU5iKdPf
rAGxx1/upe9GQ9WGWXWYU0IeSQbr2fSXKBaK56L7eLunaUlRpxpdGwML/NclRk4G
v4XHdWbor6jduw2Th8KRRpCvLbc5Y1vb4A8AeHZAEFk0g7CG6h4ihJSfVddcmPp/
E9e96IK3986PLXBBS9/ahObTBFakwSKjf+rCMAybC15JFWqwpR1BOx8jZ7IzNHf9
uY/od6HzoBKqUh2YnXIqu2xW0Y+4mnSB/EsyVbDlKDs6I4wv9ZDiGROMsBv9RLDw
23pweTtGt2alZtwU8NePA5GiBatO1FMmuPAQlRQCCAFY5FeUb7HNqUSvM6qad4zH
eaPsYJKHrw8uZPx+qoTPNEDQWywz7kHjwaFPsuUCokze2lS9PQNlGcJXIzDH3HdD
4PSfsl9F+D1b8DHwd9/wDJSOKzNB5dDc19eI3J8CU7vJ77gYZVdBHSvizIKE8xQ9
mhdUp/ZNDAwoXX+tLg4TXzBi372ajieLjSvS650GYD0yymntKWCDRHHtSHKZxwZo
Vpy49jX8nrG73CIReENGc0HC2uiIyvATg7Xa6bXwte9BuqFYBnVA2oaqpi79vJaw
JVl2JZBLVCEiLzCoVzhs1h1qkwL0e4xtnJxcKwMftJb3NQYUSWXAzy0FJPIpLtqt
/k2GxRDuA7x13G1CW4WSpICxxfU/PnJKvN8g6/mau6X3+j5DujjiSjhr7jknz8H/
AJCe1qxw98fJjq8uWZeqK/RUuKfgoXjIfT6fC6FrXBN09+ZkRx7GoR/9iswJN9T6
Pxd9PpDU8MjOnxMmRP6MFgehmu/WXIsVePs+LFeltoJnt2KWTJR5Y9TDvLGhePkw
pDUQny2V9Mkly2KyTDWQzlSTQJ52r93XgAtLtrSrJHwOi7sPXzVoUdmbqsLJAeDz
0qDPzhCUC3Tg+VQrUSuglDFUmx+HIts0zUoyP6ltnSZbSzSExaPquB+OTxvLFSjQ
gDsL0khSN+sLNw5accFiL29HPYuc25VsCrAI0Fy17pU/n1ivdNTRfi/rNCo8rlJc
`protect END_PROTECTED
