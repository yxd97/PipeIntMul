`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NL9wXV57o3CCF4KwnrY+3FEiGGHoq6SCnhvJTyzOkxvUmfzGgJ3YwGNHkrG+pFKA
dXFhYkNBHX/hEdJW1qnmXy6HDSboq1wrOTcx8XpYn6snNneE2XXhTXnv+1/IeN7n
KOOqJkNghDQFWqOIq65GQ7HBkR7qsZ3FR0hlHmLlT6vvLK2Q4EqQC7wv94A+Fi0z
i2sNYHHL+92wwrZZzr8LrtH/Txb7WCRbCHi8b7daAiy+PsF119OUcl1ZKQlJ3aTc
wb88EXYJVatdfywQdytUX7ijgxwCEPDrRA51/En56JoP4G3GaRB6EDozAcsAxtmO
7Yd6QeIAeAWN4sGJEBJtbGSZtsuZ1/RvH6O4WNIXvSybOmUEXdOkVxlPYZnAqzHW
IUQL3pr0pLizo9gCNsz1SiermOlSTaE6rWg8lLx6ujt4/gxYxw/MfMCiYX1zCOGI
1I+P+0owpebKM2lRnk6AdlbEpL32ztQSHz54KyAjH7cLcbAxhYYkbl+Md2yWlFGF
+VS0JXDt6V3l0xzUf8KXaEqyRLvgntIV6urxx3UttupF53O8EFM+U9safwZH+U8e
SF+ehBA7cXn1UAYujgX+bcFlhV9CMTkwx/uvr9hWTzuOLj3jKxHjskwaMwSwub/j
c3KSBjmYz/SeiI8T2+OYH45pw9SCVb1NdfH49hXZvbtmt36IvUkLSggGAViDR5Vw
40/HtyBuNdB+RHrOal2RLPapu4gG/nZeFhrmyUOuJ6hv+lrHOv4PKb09kOYrmAzj
5rVCeaBBlZDyYxVbxMEGUBKtLHeTXYxvkbD6lTFOuly2y50JoLyJRRi75SAoy1Gq
B4iSE5GKDT2Jwa0TPASwF+BtDDyv+FTpw064PBLfIAEtVaYYvaf5Mskju3iolwei
qiETU9cKlQQXmfSDTtdyvNuA2HiMQbEY5riT5yJJVoVqGXPPJmpN+2Xtdf+OEknE
fsQyjO4hXFhzM0eT/vYKGP+XBsNc2n/pk/yMCQuMNUWa5GG2BubbOiN00JgCb/ev
/t5UXS95KI5KJWgXnfKQF4GKokHdfvb5AU1fPbpdXvykDEg1/pLhOTGq5u7o0q5l
TVCyuB9Ha+jxtIEWlASJpJRAGYa8T/aKReYrgBC1FFgZuVYvEu7b+Uscbb1x0Cki
i66wD/Z7yRCTaAl/p2bChq/DGDngWrzLXCKqTUFdkasmfXra6vWLdCZj49cGAr3R
F426TlFxEeCfvxkU8VwRUIRzxEJYgNwNbSbcSMWR20d7kqVaMSmpTG/DYUeob+2a
0N1gE2ccIZeSDdSiuLD9MDz4nJS3iOE9T12YMdcwGS7Ex82c2KBb7tmnDpHxqMDC
AI/CJjhgMdgZET5VX1YdB6rH3CJKVXsCF1EESHzuOaycQm9oEFT2RwU1DMEOcPDc
ddXJh/xMF2e37sNdDEwB+vfa6lrN2hn4IHGym5+gE9Xak8Zx6Sl7b4J+bBDOGpjW
xDh4qZz++A2guAn6zdZ/Nm3qXk7ux/XeWtEtXk6Jj3Kf0cdBb2TzXxfCYV3p6aDR
i1bXJdbr8mr16WsArSCGiNpcYPmpynhY6mX3lbqUStfZ7/VygmgjnaUfstKB6keH
//3mo+pz0uWR5QMlTTdfpdM3GF+ZnQtpH0Is5EILNS32p9uh/jPPjYIZELsXSFUE
uBwGGAqdtaqCD7PsE/8JTrvAIjfpecnP2wPGbYhd4FyoBbC7VGcfN+E0x2rv7KoT
sj9OG0zNCZnRpiLT6qTG3aoFdW9f4k6SMEMH5f7jl4UTNnTWwdOHloa3FZtqQyWd
cm18eBo7Rj7e+73Pl5UTCv9066tU3a9lnUJOlwtH6DRHSvhVNOJoz0UGvNNkyJY/
lYnMgAERTmOf2qubXz5EmxD8n5lmcvaf+wKORsrKPfaMZ4Dmc4QJ2Q1QHSBFbHmI
tq5WyGYDZNEbA7g3CdqovJSa92lUdr9HRqt9jDNnUvuFg3GCzKN1SehT5SUZnyyN
GvrSuE8ouW+X1/enQpRRpAy0rxiVkaWxHQVqAetJsldhyGxYuHEee4u7Ejs4sRGV
ePh81/LVe9JQWsstIaQcUsd+ZiOPPTvxNgrwTaxEp1OJ7qetfwmcTATN+OjFQscr
5Bt4nqKnANt+d71K5Sj4+vmVbreqktcGgwgywB28SJmg20GlRUZIKaXYVOTq0b1m
GQSzS/tI6NwSBykN2p5whuhOqWN5kQuVzCjpIfuj+Rm34PIHibtBnlcSlJgME9Rw
jiWyjXkKaf1d5UzPqFFCV422k9fcgiz3GOKjwT3QiE5EE3NZQkPO16+illpE4rZn
KWnw3B3JDbpvsouyZJfkUGFK7y5wevyHxMAjukiTZBQITu1cW6hKbXYnXibFGJtS
BSW6XAOxW3ViBHG8sYc4GB83EfjJbXvXZ7WQNrzEcg959FQtJ5hb1EbfZqtFtcLE
y/aQ45qoPeILud0kHWUSg5HGxsmiXkMAHFHKEVHT4AEJPdoCBfkR/5StcW18fUji
z+if6RZpd03OeEetwFZh7R0VmgrVC2nLPfDBAD7eBxlu2gwG2W9rbh2x/zNI5lkp
evSVtM2pUz77hgahmT4+YzaF/4gOAw1g/0zvOgXI23IKDlK2OfE+ArIvkqGQdcXw
LtwYNV1ISn8givDLX+kDgCGDn0CZdF4lw23I8hVyUdsu2qAOv405f/MLNyeVAf9n
dQH4j6iQ+PhPaBrZjsTgzkFqcV6Nx72AlM+4C6i9MwoHY+ZjRrGOvBdOTll0iyei
qTLCpI44H1Zx7fM3mMgrKUL0CfPBJf+0q0yOn6grhuksxrgUY/3o1UTqZ2GWGnpO
YCvniLFT2W0GOHKjtlQGq0dlIfYr3FlXdG89ZuFwPC0w49J19MkhrP0TlOQXnf7/
kSvrgtjHxXK15kzDWqysIafetcI1q4hMiGQGWmMmJjTL5PSU9I+dzMAwyPgqt7Yr
eZ5X7w0gxdIFSqLoYnTm6olvNQU3sh4fN0yB9/TBKqPk86/KoEDd00+rjJKG3C84
HNj9Qz6yNfM+KyAMjGgTVHJNiqvxtPqJn762T2QrOP7GUxXKG1jROXSizQlHh0iF
yUki9U81ybSZWEQUVPLr3Zewk+mFyMcps/JHe4RAhXkpvp8Kw360g2SKQw9Qv3Oi
D2sb2eWK0WODIuvvHkgNsyic6LEAVscSLwbXkkAp2b9VgQeVQ7Ix73IXNOsAcTMs
Qi3c3WNeHbhMgoTlDhkjVS944mbt1ngBWIm6oIFt9KI1wtpv3V6WBEVIX8EHkv9U
MbwyUX8/ZzdmSeA+2fa0/EGQXzPZQeYoyqE4KgFWJq5TFWlOt19oCH6JjihvuAs5
VfckldxBbRyQVNdxHh+p29M+utP07TAp7vScSj4BoeIWbhxSuAYSC3KP4ahmPAjK
X6QBEgUdfr9RaCQAz5JBtq4nxXOI5lRgKyz6K1qrH/M8qVGOisFXOon0Ge0u2Ycx
q+L10INQGZ/qXniRMLIRNy9wOgZ3KhJiPFRo7gu11dj+7WET1VYq73eixfFnu5Y/
17K0s26kaJVifrumXrhPS6KslHRZiaycWLOf8x/JvEoTrgNCxwalyKCDnFvjbUyL
iMRqRs631gSc5bF3oGEsvCHSgCS5PrZiQ/ctfFOLNDFqFdJSUtecT980IRjOM0yJ
6d/1HWgbTa/kZVVUstPchwyBrkhkrJup8GXWgrhFRvH59BxmIY3sInBb/+yw2Nv3
OaAGcg/ywbsMFItDC2yOd6h5J2HFq+y8PuhZBHbUQK1qbh4Y1jmX9DlFWFM98OZR
Zfavp0RKzqQmx1R7x3XKAeIWyhX8vewznJrc9zd9jbKjNcAZoial0hpdhkQqA0TB
Oxh4ZDH8AGSgoXwUAvRSGYcNBN2uZfdra1hZptgkTcSUKsZZmbouOjmNJNOC7Jww
IyIdZV9ARBNTthCHxbPfw3GR9f3NRTWg7EACm53bqNG99hmSLSqEUOdC+/BdAYVH
M6EH36/608xC5IbZFnyx7UhdzS4yUJI/QafCi9whn+ahCirnOjtJI5PgUEytypCO
XozgRah6LcDEZaIjq1BOUxxwKOwPPmg6Fn41bH778/dyeJH1rCy1wXYJ4/Uz/gA9
EubAnOP4CZHW0SohlSmTjxPsjxDYBto0QswNAa+ldIZrFywrs2K3K1ew0/HyPZ93
hvU/fFCpNyyVHdf9uwyAc09dEF3j38Ew0JhkpjpqhfFO5IWJemU1SnfbSBazp8Ql
VAdkllb0bPPolz72EUat+xk4orNJzmVrPT2hhrpK10LKcOwdVHSrmAQzriBDxyGN
z2ugXOg14kffQPPcoMkwdcepLafhOxhS733PjuoREM/pwMQ4CU2lYaEP1haQoeq8
pQ2O6zdGggeLZfXLR4nckqCjG57fb6Is0UmVpsphAPelosAG96+EfNsYi1S8vBuQ
V6ipIRl9IX+UFlJPUBsmoXbtPIzwRZPZH5kE+DSsAt4XFBaqVFk38nJHLuSLMPOj
6hwWdL9t/7yLfcQJjx+FmKpZZ+/pot6oTxptajzNsY0wiGlMENsDG0SelXlB8Y79
k1W7JQDzvbYBvpi8tDx21Pkf9zy/8gQubrwuL4HqW+Ej8yZUyFpIN39jG5m8Rzpt
x42QoNd5XBNJOlDLJJ7PMqGht8ZfpwRhuvSJc9OuGkBfmlKpB8j5RHL2T7acdDya
S3xZtj7vBiE4C9ivrIPmfhY/nN7vkxnCR8kV+D7Fwb/JqZr0NTE+OZD7xODaz/dM
16qRk5CDX+mU/DedC44nZckbZiHy/0kgfmHRUi/c+KgIAoZX3+kJXWTdHBb4+xcE
jasIj2D0g/3gWavbsjAaT/EqkzvqEWAmNzT8XAuG00zB+v+Vc7/Q4tByTnR/aep/
d98Bah9j+vlzd521oU+GdbCkixCdA12nne7Fi7it3w3Np4ZYWq98wf6z9TnZc10n
YsMEfv/cj8dW1IbsF4hgmyxOQhdyQRVl7oq5PeT5vzh9XIOSHapjDa1ajNOMGty8
rFOOuIHX89EdZDdA+cH8cMVubHIZGa+0K9Q6tdmuxhPrh+hZqZ9ibh1eFYfJ6qA2
o5x5hf824wNmCiR+ONuA5AnTyY8CytaKCPgZTkdClFNTd5a0tYed9IYW008OBTLQ
K8ocJIEGbuNdktvc7JDCOapgstYAeejZTvloQ0Ckj2zC/2zLSeFRpOYomMKb66kY
nNBf+4hv6WPKFPdfj4oMD2yOETfEL3ciIJxfRvZYb0KFWVedB8Oochd4/WRxkrX6
cl59TlU2evy7xEVYWJwbE6dNzOJ/r5kU0LABwg68pAM1Flr9gaeUd1iLi0zC5l7I
nnnLourrfugcvHp69q5GRdcE7cDd6TBJjh5liN59F/XlLk/GfQCVCwRS1KmaWhDP
vI6HBD5+qDR80P61cTHvKk8sJBcqpyt/g6XDw56vjo4jZeJsR8z3y6xPT5sJoHnN
kyN5v6Qn1m2AXbgE8/4lXpWpGYAE9ls1djl4/pPMdz3VGGScBUYAwHKJVSbLd/05
fjZpEXMIXW9/LYQYYRuIS4j7WYpAB/PbO7w/RKbAGTUPiPKLDnpbuI8T1CHbNYDp
1Q3Nwjkxf+0XAqCmCl3VTVb9LW1Cm6CDH66oLAFN+n8z0oQzLltb+DWefpClZ59Q
ck5QSlvyfsGL+BW2Al8XyYmsgK1a+KysYpc60pFPtmmUFmQ9ICByxfsWYQawNDoW
DQCeZnLZjUkOw7q4VlqDTB5kShKBEFca+QRW27DB+qGxIVzrGqf9YJRlkn4YSDDe
pU9o215ocbVAj2weFDK5jqCyh6+OJFCIi6ODusGISsKQheTDhNnQwi19rjMjhEEj
AfoftlcEKjTnGhU08xyw+P9ewVb2789AuzFSijZWUORYDT2L8BqQywDVHKEmc8QI
X4oUcwJKf/zSAclpSautDR2LefGT1SUxhjS41yrHpkeGKxrDGif4LIrVQ414Ffo1
lr8/1i1qPA64ewYQqSUxQ/DjRs28Z0jZLt2aWZw1f0blnuAhggutUNqxfeoS5BgG
lrn+xD4ZqavO3UIqBpIPYmHkxbjGkpdzcasCSR8JEl7/uvYEjBkjq9HBJzYuGJow
XD0MyokXTO+ibiZc5KYMoXuO2+dK8aiEMOLDqY05AqjtauQUKIDALatSSh1S68MW
Eo70CJ5uKEcY6ZE5otL1zHcpEu283UMvEW1iewmf1x0Ise0wQD9jioma7V+FkSQa
MQKwB2gw4yrDZy6DDYXYigsROZ76+pODxOc+d59RQGL2m5ACTiQGJ18u4vU60Aua
Se79J2Jf525CQYKPvMx3iiyyPnByFe9DTXvT7WVU831GPl6KjkSxdbOe6FT69e7t
oMX9HFFj1qNRAOK3iYvPAH3K3ibBonfBWhuX94Mc7h1+R/5R5hKgY9wGFI0kHaS5
nD2SZZPmu/dYkLBo980gZqUmZuR4Us/HWC+ub9tkqo2AY3G+YOg9hRYcudynRvHS
/Cn2oPShIAezg0G+GfVSpshe1Mop+8tBgeM6VP3ePu5HIw4fKrruIJxxAtQvk/3L
rDNxJevSMtRah5qBdN601Sq2G2TLJwG9+Nkk+61yYZs81e6GS7tFz2uJNYAz3own
pXsucoAd/1ubOzJMP18mODqRdxGqa2TPRdgquHm8sswxM1Hyy2Ej/UeMHAfI0XTM
u+zYj11ZZxOU3NWkYNeBYQ0n/A9BKjyPGX/E6Rsg5rmxs22pq7d/bwkjunRsBtMJ
yuajg9lc/GrvBMiJ+KHDutOvinHLMkp+JM9lWzeYP2+JXIfo8aNUA/L7y0J9ZEOv
4ubhwkuVycl06jXqZC+6ewQZT/+H0kGbNKLXjiQHVolQH8YDfTX+B9tDClRV64cG
6A74s4+O17TENsQhby+1QzuGx/AYhvQ27n3h/9ndQcViT72k7LDycjwzvqn79Hhb
MOYXU8Th9liMJ+BDt6VPgqFZppE0/PpJ7hnE1O3hhpaSvtnTf56l70zAwzRM4muN
ywuIELMR88iJJEw9xZpl/YIHr+ZQQf4BsM6lJcvJrS388BF5BxbFnemjAH0/gk2p
fwyIRYbe/wBzi5kq85XexcFLkXTtGeDTgN9DB3u4FszyoFuiSMoimJzA/1vhQcZf
4DWOXYcKtsjimN/MXh8pw6DwvYXSDodKX4TO+ck8ZZIZC8yTI3UxkLV/8IqVWZ36
OmGfRFdfrDxMyq1FWIYKXt/3CAGyz95IJYFDNqehzliJ0w2yc8k7qrUWPSu9xqoX
yTfGIcjMRGguqhxYtTSfVGgO7Dvt7bh8qyDEzQwG5Q9ilx/yMmUYRZon7cyAPwXg
JfJMum7EtMFJtQgO4NSYEQZ5cIKY27VMureNOlJ+cslUx3cUbsMWyL2L3hXECL2F
p2Q882WTudYgLVIoEWtghuPs8PZr859ARXYLyxEMTI4WRlpERL+w2DSWMka+GKAv
Ofq4pE1hyy/FRRvkky9tla9NFzXnR70qwmq0ERYVlm7hs6Lb8pAI6geGADsD626V
WQ8b9y6ev+WydRUubUVGDUS8FxJXgWd+S8CSpjc4Y4wZYiBVkDHUxkOiIYOzYNe1
QB74ToN0mhVEKham1QeKoDOcftc04+sovCHU4dD70ApwWCcrzXVS7pcvAivtdWFf
/vD7JOF0k58iwa/HlwFSw9/F40BlJTWjiMmfP0ksaNtkW3czTnQ2kvNrsIUmVz6B
zqo9lW3gs23v+GOhqLAegwuXZPXHXLuR/XiaZUHFayg2p7uF8abjPV/5dCdvWQpR
OttRonGEvmZzgLQ8PNJouTeUuyG0Vosdl/5JdJAtdYidwRNg//GepfLE4D5B9Mfg
xmtbUwgBKXdFNiWUyZE/xHXYQ1H5iwrFiu8EBs/shJkYeYrYVRZKu5GTW3ad6NTF
T13ECQoE7j73lAPyXaUCV0nOOQel00uOsb4zuCwq6UzH0sc7a9hPc1DzyL3r8HI0
lb15IoDFF4KsIwB9WfUINWL//USB5TGjM6t8z3VAE2amuLeI+bnr5KDNEtZdWhMa
DFtJc/NrSBMBs+tj0zDvQoylEvl6iUcgYdrO3MfGBhlDEBMcpAJcJGY7+LGAujOH
fDVxFjBdN5JuClu0sF4JoDVYdwdkS+nG+wlrUchInwBPBYfuV5FhJ0ZkKefawTYk
5BDCi+RV2lgbB5BOFkIstrCyN6/2F7srtGIK5pqQ1xy6CddsXcCPDxAgZa+7qjOx
X0cZul6gNjXztj4LK59W7dXPXc7wUaMoOChGjwgbfe7lYmQFLeCdLl5f/7BK/5iD
MAKcZKcL7U+kNMZpXGmy0GGI6lBhLfYLNiMIzNf8igFU61CNZPBF2G2OkkOOWSD6
yO2FbT3ElTHNBarqQ0sf8hrlbmXrz857RWgbE0FTTyCDZI448taRQfb6xdjIfhR3
lTg3P/L/IhI9TDK60hM/grRWYZhGh6PVYdXrYnTOmcSXYdzSD1Z5XwGuoj1THrAo
zVFcCvye1Wq4dZoKswqaLCfOL9WnhOkSH0vmtFmec4fSg5lKRO5uydzs9CJP0LPO
Q4arwQHSEngHC2WoBx21AQtYb/Q+KJBnx9Kawi/Ji7cHkIMR7uRbVbUQHIwPj+do
Mfl4Q/fHAbE1Vnaa9fkTO6RU99/lr1ZrYWHco6A2QTlJvFauWGyi+9Pf89fCD8d7
jU8qvQXSr5i/J37h9bvwXgXEBChpMfUsLfEWKZLcbmKdycdmz4ArezB2cAP7ZO4X
gZV9sEAyicTXl9jy7Smu6xe016ZQz4cPQ6zzkx1+rLbH7cqBMQkhYs//46cDeHsf
06BxwbWy49V7/l5btSliqObkxJvW9ne1KZ18qbJfSyqy01gYP7BLH3Ie1+V9Q8Eg
QiDCExOudnZdngxzy1F9f4w08/uy8beoXdZyPcgbnPyaAwgocJe5SbUoSLodC6vq
wP6EqpNstwjhGh/deOj4xiEFItTfy/guVICZcl0hg3hHuYAkpIA+Gx7bN3/IulKd
ReI2KSjhHCz+zVixiyXm+4U4SfWr+mz64NWDtp8hd/dlXj/oGR28kr+y1eM3g2Y2
WraIkjEQuj+iBFdYDcUVVxCHvXAjjtRN2Q26V7EzPCXomlA8POKQRCMSM6w5ZvMw
zayrAXtgGvfaQjXk+NzUrM+ipobloTIBcn+swGGo7BnO2HviNFskHdtLSPkIksbP
PYuxe/+zhFU0ttEWx+GovYGgXIkxrPazrBWoApdNPeNcBQSNMO8zgffZX06XO5Hi
rjccapUzc/Ek9sxAZ/uEAp5ZKNZEgZwwIopFZ0CGC8i06ExLfYXs2rj2EgSFB9bJ
tjrzSRrJ3o5Hu0ujWPljZkCZqIUEIVokrG7BruX0Dq/xVBN842A5reT9y+RtMbXr
ueXGyUN+HYFZvoyrPyxypKtqyKzJFCyY9HLQR29npSO67BRHq9o4S2bSBD30xbNi
oZW/nou3bHmxCQnrkv2nZxQ76aIB5NpwAUKnwMHOXChy076v1eG7LwngEpbkpuO6
6tbEmstjRoaD1Iuz+TBI/AyohXbI8lq3fNuXOQl+q8KINBXWXVkWHBFcPDN3UC1y
Ldh0zQ6Akts/P1SOG4wYYHIIaHkpnT3A2Q+PiJlLnMSQtLkw/d7hEo2UwN0ymCs8
3Mla5VenAVljeEKvxBuScCZZJHyuU0u89bGYjy0h5CwXOsJwDTvWiVSJTg+ACQ02
as8P9zvNHB6dvNnqGpb9+eExeGrAmeHzabE9JMqFI4MV6MH+g4txZt4v/CR1kpou
bCHGTNAGI43Aq7M+dueaUUgmf9+B5W5yIScXCABBXNrtcZtXGloU93zeAupekCsn
QFC+/+3j2LKClfUFTSOxHOU0eYBdcqp/92jygk0LpKwH1Wh/Xo3cZmOLFlgNeKBG
ku7UclrhKQM3k0NzRIOHcCh9/CUJ1H+T7H4jw0gLk/plxcX5XSh08V4usuWcDxYK
5BUytF7lM/hfrpW4c0H7uWWCytpy8R+qINrhZz/c17y1D7JySZi4W+Usj8f/In7E
1CUzU/TxgDmu+SwZb4SACcnDWHgqkNq79uneHrEJuEZJpkrfwuxBfBAKRX7o/YOK
/Cl0jn+eg3QtOub19XlRitxKAMd0s3W4bfcfdClAO/UGBq2PkEc0MNP6yaM9A2aR
qWsU2foY7FHbXsktqcJojkjX9AXjpU7bVtNP/LXYWUsq/tB3SSZ6s3taHTD3XO3+
b5kxd1/KounFXkdjb+A2FpEZIXC+U12zSZOLyy7Ge27nOFqN9yvwke5+V6LXyj/Y
HRlDvnz5hoicrv5FzULRAPFteXTno6WUA3TZK3eaWZwWSANiptjN6IhIdPKksUPM
ar8bwqfXrprN3lRm44S0CaUZ5Gq4GJ4mnd79XFs1jGxo1jUrVI8nlAlVtsU89WMo
GimxzFpVxKyFQoa18WnUdSwIrJLsb3F6cR5XDSOw1C03A/4do7guQd23vPFAZpAG
v08G0yxNAInG9IQbSpGMYisXP0lgapmmkziSLH6RNNvR26rTbfxzUsctem/N82Eo
237qz75qpjJRSwyPizncABMnbKkoyqPZ0NIVHhbagkAL8p8ZDDiVmbIlDkQjvYek
rkqzQolFM3gLIGkUN+q7RSPtTERzxkcJ2MZerU237WWE7dbvtXaM0Z8+QXqPHO+7
ta0kzM7UlhTKxkVUeNOizQH4KZnDXyD2LXSQrkYdQILD8BwvZ4Oh0jwVyffd08mz
z98N+v2UXLBaYkFsF5GMh501/MIy1Re81h1fKMZ7F2fsvUwIPMARlnVleFQ/PxfM
PFBL+GDrxhcrvA4brqA5lQ2qIU3U4/U27k9sE/IhLodF00qItUGqu0zDZaRf2s66
6RTf3OrOnlH6vYZJZnOy0asT522ifnMAzv4T5Q/lTg2ZCCdWb2pgTSQ3oZIGhZgT
LnfM+M7inC2qGw4e9Mg4unNMXqYsALpV5K5o7hGRS+fycWl/u3i30O6RFhArkISV
Lso0cNPqDa9VEtg4PicHk361oyXqNyAk0Mr1J3bqMR4t19l0uj0mG8E5ihtucrNy
wf81aEQZAva3MHjY+jqru332iAfFc6nwDg1Kvep9yFV1oABvQekLQtllxvthWqf6
4YWWWmgppb5d07RFlkr/hkscnrJONlaGtbV1IjS2uDGURZMXFKUxCRLjhKLGAHIV
w3+sytglIAKEQYCjQB0N02xp2jvdEDg4qYATiQNe2uAlLDfWKW1VzrUZYz/fO3lx
/Bg+4QtMih7kB6m+0rl8ntpggOMY+bN7DrqYrCPDCRYLEIpp0G3RWjIb+OonKnJB
FDKgH4a/bU0eqMkCAMjzcLtMCOfAI1iN20h7AsyrvNo6NalNwbpUX5XAntnaI5SV
+cDJ/XDVusVCzXKn+DrPJ++SbFoYzhkUsK3KtyMtVFhrijWJfcOhrxKNWCNb0XNo
8BVhmx4rlskKYqqyQVm1uLiyHYIL9kQ10fDZ7NGuJK12/MV4YMTGXmAf7aVS3b8N
mDg2iouzscsW3chr3uZpw2ewwjFiyz4K7IDR5kRska0gmS1TSqOJfoOl2DingcHA
sRG47faPfJYe2LIXkHKAtwZuVDFDQu47YM8H7MJhMrlyXppfj75Fb7w0l1xmqUX3
iZqiveVi5RPWjwQ098ZJKKBQLnhIVMHvg1hvFIUlg/GfMb9sbZZnmmyIt5X2rU15
3osEYDXr5KIFVpL1pE0+zwI5uGCzndhU4IC54NqMO4Q4QLC37PebyWZQF2wwyqQo
FTU0wOPCGbQoA/444/AWayAOnNE3pr8FxG+qBHl98iyR74l4rmv2RFzZ6mvT7gL9
SjQs9VD5hrvVBQ9cH8f/E94ZMGjx6+gPOdDz3vQqt0YzjJdPIDLoomKeZhvRVz+W
yvfUNRYXA13EG8IC8fUYlmi+lWc8cPDljPOhnKUd7F2R5rE2mwcvHo3760rMjBLy
5x+44O9sDWQm6SjLkikMzVe0lki72v2eiTOKvrXR+Kq3PHQdCnzsQMub8siWttaR
wWq0izLs/2j+OO+hoIofOwP1rY0DrVdnYV8d9T51Q2AkIc8+r8c4O65/8ih9/RK4
N6EDdjda39UIqFv4BYxMc2mbsNMiGlTAeEvA6RCFO0u+SM/Fq/dsnoHeatefoRRC
YTMBDdaGQZJHceWKShNhqqc04ZzOnr96J0EPGbRnC0h3a+e1moDtHezdKg27Eqsi
qvf8+gkpfhyIkO72rYNAvrYEtN5HtPdfe7APGj4pRx7KWLwrHtSuKd4Tm04++zZf
wYwuoOjthVzojJAPjsKT9Av5e3LQaY1pJdKCXR7e8ue+9dx910C1CeLoP8p4NJEM
gc4cDnxQuNJR16SzV+Iq8E1R52qvG3wbV/bzmITbb0myslqEsNkCo7RLrxh6sQYE
uqy8k0g13kcR+xsfDwbJyztqQhLz1GifDQlQCMSoCXjJzAuFlKTFkq1iugcvk8Hu
S53/mzHz0lk6FvKi86C6Zw7kNqvImjqmpQBMdDz2hetO+zVbCfzdyTN8EGIGWxFF
eTVyNlogVcKDEhJ07Gnk6KVGCPdm7ItWrzpa/kCCr3tcrHQUlzFlF1n3bbDF6CKi
77C31w/uFQwhsyC+W5+P+pddKjkHTFvj4iDq+In+4wZqWSP1vFEoiUpmbs5wTMvz
4ttuMUcuphOZO1BT6so+8cTRQPWQhBsP2TfnUeSPKhh0hoI6rpBu93V/1dOfD6kB
U0EcAGHNYgy6a4zXa8Sy8xSrEl1YyBMM1/ujtwvLd46jAJDJ+EJAYo9luwpRI9Oq
5LuR0rCD2TeOhktOQyc4oVJ8u8/qjSyjKpnMxTEPoNFOqS3YUu9jj11TPnb7s9tj
Mb6yLgM+EAoc5GdAjsQcnui2qD7i/MiGk29BO8ItDE8I0uCf8TyGcs907zGRi+EW
7sJec5eYoKo74MA/KA4orIt3lXipjqd1F5r/lPs1nD9w7n6JbzfdhH6pwyqrvRhL
qxg4oZSlct6Gw3YOrYfftJLnceO9MV/pTUl5d1qTdRlA0nihCb+i783UvVqgPgT2
wCGAgvhc8zzm1c9FlH24tA+ctH5Kwq0ghXvX5k9XPPm2KorRrbFNlZ6HT7JyqFAf
i4+FM0Na28YTNyKFR77w+kskIs99ijDAhECZnNWVPA4u5QCTS/VINHggL5SLoqji
FFX+pTwN+xHqJ6SvaggDDFzrfNK/rIaimiCW/kxKtanV7nlAwIqdZsT2n+Z3tbbn
lBpcQobCHsC+nfiIhQujIxBTXOAxIShRhCL/Lcl92wRiz1MgosKLLQ9QgKk2LOEr
r/qjpx5ULNk+M3YQvVzPG1zsm6oG1Vi3/JyXUM2VJyE0zJPxB0s89a4D7BdEnoMP
hMYgB0WGNSOSlbU6Q6ZCt04Ssabj0mrKuoIqQ/K9do7EzObADX6G+psLtu68kFrg
k5CA2KbanJSb5LKO+r7EHhcSj+qEhcTGIy4exWGtog5EJC7v0drZ5ai/LRGVIKdN
xvheF151quF2h/rXT8RDwwtbcsS+sAixqqqm6WdYiwSFvIwc6WIubYWhSvbFIdNH
RPOZhIFqEsCt6lnKvnYSxgVRkD9GarS97RtW+Qv+CfQZJiYvTFkCdC+SZiv92Uff
Ck9Cbj8lxmN1ojwNQ94eG/6uYf4zPvBTlSLcDXmoL80x+fKLIjDgUq2b4sX48jX2
n/E8A1+zTxJzZcDx7YiIkqf22KtSWLUXshtOL+FEUQ86AShunEs7uP2YWhCi0DOk
o9a5nYJIkN/WWCtASoT86AqA5+gnXN2/CCaCPB2ls8FQPkfh6xlKkwXh5pU1/Idd
Is53zUAgqcyzKhdXY7HyiE4/3ralWHuemWv0NB+9M9xlXs15bUV6vSzd4YztdRdb
2EWvFbEvXQkFfIH9nz+FIRBWmHWr4uXeg6dek1YXoVJr4B/yv8IUnMxwtrU08BRx
6q1t4L2CsNcjmEpFJ440VmyKiD76hQFEZjW8FBBzWSV9vKNQD6nsKMwZYYUbQU2k
rNpOwOCVkt9YyLDzGklyaTZOT8/zpOneS01hHSeYbNCuoJTpi+J3Z6rFG3wjQ7lW
7jPPDjI/6I4TwCHnuLzUfxeZx5Ib4O6PKBYz1RuGhI/B4wHGwirIf++vQXFHykhO
sRWZcEw0eHsdCPkXZcX5Lm//ZLtFDmNjMUn3dBF99s7/l4ooKv0lBoA3ofPOiqZU
tmpWdTvCmjP3IJhALpebmSt5CyIMISnEqRRsJJtVq5mT5dwlhF9PI+l/uoI1ue0Y
hdqyfdu0quWwFrbw22yHTd6Rm8GTx2WnP8xsGDuxngrMmnnz5mAG1ECwQjZqho96
GwbqOAApDpT+Lo2ROHZ6smYs1RK3pqj4wNveNpSRy1WubaU/nN6js2IyYcBhHLB7
pHzgORR7OYZHuJyNwvRJBDxYa72usqbt5a/SVDKJUbPy3LlIhqZ3Qo5EZpaCDfoS
aqE3rC3EoBBW11C+apK574/yc/CsqnA+HNvl6rRlh0FMJ0wGVZNzqGMoiK1NWtjF
mvVPiZoVhEWEwPDLagkSACnBHQTPFBpL29bsaW3r5oy3k4KZXAfbFmrjL2Xq43MR
uwL1KR7ioB0x8wr8UXKobioNDXEHnghBImI9j1Ia8WrgwnGbJL521x39tNwI4CBE
IFHNnHYMKkrbxv4/bdyUmQAVwxFH2MvmNtpqzXyYSgxqFD7agT3l2LftIkOtsKaY
JWhITVz98lQSY9uUxuQijHd0POjXH28J+7LmGDqzetXmtTv/Z2SgFcbJtTAWQc6D
i3uvM3hE04vrpEb7BDTZsgMMeLDxegFHziLE4E18rjdZIWzIOeX3bvxRaP3npOk1
Xb+VRvgOLnuuJuSWGaC3La1lCz7YLeDql4WLxijGca08EpfWt4JJppE406Jg6YeV
19mwwsLqQhit7yJZKY4mzt7+AJvZbpZEh0JrYp8v1C2vKHYv/IWwes7k1kH8jFWF
iwtaeiaSKVq/GyVPqoBUaEO8BxQ1j6iqwME0jAStEG2Z59qhPKSCJR8rHx7jwXV6
ZERKiX96f4h03byS155vFPYx4WOVnbFJpAU7ou2D3BbDUuGDsZGVeKvkdLETvd7a
LTo6391HWAbFAUfTTDVcWNhWFLlKQWV03XXFnHSbMrsMDimMzL6COD3vQI6mdsha
gH5VL0ZHvs5DSar5lbO8CMZt9no/5QoMil2u9D3GmeP1Ih91DtOrv3RSNo4kkDAG
uAloD7f4/PolvVSXA0h/b/Dc8WTGoNH4544WYwcdzFLlzmSe2t7tLKsOUNFntG2j
JN5IMgXYRfrt8x9KEosxFYucBOkKbuz7/fDllvKrgjaVdubn0W2QNxteQEnys8pt
8Eq8H5+vCJymt9oW3WNMB/JUYC7XdIL4Ky7IEHaZ/xem3BzqY15/CuLF9cX9Zg3v
y8O8ATXog6rRY60acLBjCtzvXagn/lQzznY85lMoAjuB7WuPI89Awao+SWPi69Q9
gqbs34T0CJPIxQ6fFBBclLKdgFM7s1i7J9Wm1QDCX15Bc6Z5bBlPH1x3Gim6rABB
UYhELvTSOAlGmEe0UFloPlYi2IlwexmIBPhr7W6t1nN8lbiJ6dWeJQL0otdg3Dk1
2TdNwOokRP9OFhaOH+zP71Y2EzgH9t+oLzd/HlGhKvt6y78V7xCsCG2od6oIeSOk
I3mcya3jmFQUTqUhoUcqeC0OLDPoOVWMe0+bvr19Au9SqQhTp3TRWt6Wy75vBSAF
bsRiNGD5y8BkbJD3TpTloHcPG97A8zDeB47RLD/hcXDLRMsLo2Hwlv4nH3mKOJg7
Oca/42pscNynPzdadActPpDf/K56CdMzm5VK8HbtwjHvSpe+0yiW1PaA/XeWOV36
fx1rjEpZP75MKN/ldOc9l8myUAg7OTzYdpFqEUiLCfq4kph2/LwqNwX2Vkwz7HmA
l1GKevgqmjzSBQCONwVBfK2KuP220djz2sPFihNbTU7YV+M0u0/z4S27fLAo434L
ZDZvGt2Pmq/upQGU6MJOWnfUYoMP1MP9y8gC3LbAl8TV0HdP82JrQtnJH2LXkq4e
loY16VkNwabkXAfMw+cIahJOJVm/FNUiC5LvK0b9TqZnLsxLw/ndMFAQWduisDvo
OMFYss7+7bK2r/rcHR2/xBtbZQkGSg7eGb3osORlc2d/tGVbHloiysHLGZGCxFLn
qsL1twlLQkEa0AdUFesJBeIdwJzFFu0DLSk/7ZtD1fZTRlCvVDAuej8rEWgW8FNu
18PqhMOzleCn7u2JdGPFUYgHeVaXN3g5cMZZSO/RrbZzaS8trdBQM2WgEs+rUzk/
Qe3jnHBkRThCe4qBaxIU/5MAfUdkwSUyi/czXexJNnPwjuXYDysGMICMR+KcbZJR
LoeukBzzY+UEX7f9JD16HxvNho97vwDA+GxKdXrkcSYUvmrUoxSwt9pzujhvylNs
2+YLDMKqNZQr3r6ywK56vBTK2fNOAnpheNOzAy9qkSUrm2IE47epP9woMfRJQwpy
gmfeJ3WKqiYGURjl5U9Ac2nAmlxemsHmbLPTF9kP9UxoEon3wYu5H1B520LuhIvS
a4VXUPpmTI7K0kBAhPXcDDbPupM/9BMuBAtb9ZhFKs0uN3pzj4Lg+CJIL7RLw/L8
6BXaHTLAPn9UbDKmCMw9NdYnGvhKYYrgNeExKs8x80Ph3K1rcXcf+No8AzAB2DFn
OLWNdxZ+nNcWckkoA90DelmtuubJiB3iiO3lftP0mB1aqIxVIAib1WY130A02arC
Fs6sE04LgYuGz56OBPQrXUJq66vlmB7sSK7rD+JvXofl1xj2n4wFVNQHS+5W10B6
WtKFYq/IV49na4ctgW6eD5JJjZrf7LhgEVxcoolsr07Xal97TcMdrLFBTRKY/4n7
yeDBOfmZ15+RCI4wDGbvfINpPvEcVOD1apt2dZo2n6J3WuPgBNlihVJZHi5tyAu/
+YXoaiq07rB7gfnxj5n93DjUt5WFAK5sK+1/98Ur9w/VYU8yq8xYPgv/U3wwcSw4
rlpun7K2vIjPoxlzEiVCB8AHrHO1QQkRqgPwLyjB4CXB13PWdhP1NxNK2NbTGG3q
NhfHzilZ044Hyq9ZuseDC0b+tI4m1qcR+efKhEiM05VkmIF7/oIyEBQDVBs5calM
91cSzC49tY7uX774hijtKk7TA/wYcDbX93eMIEHejSfTsf0UAwbQpFi+KEl4OGXG
//zhAPNp2GzJ7t+oHilPxAmOFCymAXuL0l/K+/T+MUhD3HkJ5kba9YFftwJ9E+wb
w/8nQlYMfTD9vHyCahIj7jVVxLmNKinZSaew/d9Zp3Ci4/tIP2OGWC5/kw01bIl9
Yl1mv39KzNGp/mKqmNbojXLRUGy6UAQDu5Z9ZHOMZ9jKeIHzTa9UPHSuzSLPpR7Z
FW/pfUXDh48M56yLydsrC/ryDzGKq4K2Y5bObwpARKVT0U7xodZ3FiP2hQWQI51w
LyP4iZr0Lamy4U0RaN+pCnj+yMYPKEIz8qSBAaWsY5ce+OufkEXINhPDMLT01v3J
T6UKubpQp+lkxiWhZVqJTpS6IX1AdU5vCr9hZfDMVWdAlMcYNGDId7nhhz/HjVb4
Dav627+TmiC8q1ESVwBwGKRb2V9WO+1PPTQYY6vWOz1ozNstSq3wBfUUPhHaB5Jc
jE3KRrnE0kSRrobwutsbGM6KBV8RyPJXS+WqLryysO+Q4RPEEfd64v0ZRABKwsTi
vNTqZ+u8VrwMXAnIkZ9zPQPSQ6yUWzm9yG665q616+jtFdLgeWBpTWPWDJVL1fPj
VaDvQ/QBODlcc9MHOEiUiK/kEeBqOHL/O/of4rzS2Pd08M6hGn+DszvQueD5Iibr
0G3hFAJ1RX/5SGXe5Im5We1MUHBGMqW+j1Cp7t4GvpFkXzBICii3K+2fG8yWV07J
w1HHGHWMvniYfXbH1L6nLXm35XYusjTBL3sKwvjcKeLO9eleIZ610BMGyHzwxy5U
8SnM8t3asNlHBINHVOaTxwTvKaDVRGPGkecWFH0lysdfXofunxx6EevHJzE8cUKV
mWycq5yfuPH5wBX9+IrDTv28gOoLYICpsJkyNizk/CwFKRCLsAWLVgJaxgmCBq1t
U7IgtRb1CoqvXYfVD5dTMx7XlYB5AJ34ssm/GS/wxdLSTCnoRn4C8sH+i2PoAJTB
vZvt5W7O0B9MjOtj5AvXOYExlrLvATwBpTRaw4Jdiaxz+P1mNwgPiIxKk4HMzl9E
xGIgikX9AxYoectGui2WH1tm0u+rgHeNVRQ2/HDJE5WoovK70+dRsS9KP9mvamd6
SqgfnLwIrDNkNbJLJPyeSVKHSjbOBLffcchXtzp69G1sbaIekQnHssZ3/DikLwpB
o4mND/bFMSiDVK06aUxlzJ0CzoFL4omBMqIaCj5neYjKRWPFAsbWUMnSWfN2v/sM
5RtAWvtlpcwlIN1MiiinEu9ZKFMjTB6VibK8QNrwwIVEFz6Rrdmxw0lPpwe0Q1xF
L19dvQPx03XGBFSE2rOtyVSFGG9wWq7pUHxtI6pK9ERPgQh3diuddyp2HU8eGAbB
p/yZXm0ELb6jLaaAI5e2kL2tvU6FVj7lNGfXbIf9/Vl6pXVorqIltMm74nt9Wq2p
aUeMoFegaq/TKTsnezjoIQ/Chor/WZbA44O8ixPacc973RVZsU2DYWxhoVlEIO4S
rD1c/gtC5/MvW25eLlb9WW8qwTvAsvNvZFs0kmBQkcdi9VwXm+Aylt8S+ejhTuX2
5W/tewPrn0DV63KAOA/6ACQq7eQsOtTRfzPV7Hv+ryVPwBWyy1AfO8cQlocBq2Hg
1PY6T6D0I6dB7fdV5SHg3krq5TAFwPdgkDtoW2Xk3kqBKR5ZyAvDKdj6kEotu8M4
LT6ACcP6h07DSmRJ4PAAzw+MYd870sCe43zwGfnVJYmdPnvAHU/b1c+5hZiR4c2t
teoGjwWi0lUNOGm097qgCaVQ23Ls9N2dAWxgOhlaBhJwVKFT/IUpu5PAl0dtOaKV
raUMw2A6ZuzjlUEFxvt9ZBiWrwaVRh6JgfHSqasstCxY25D/rWcJa0lttqWCjugp
1vBN4PKDGMWR5eW8hggJ1VjJkqaQnMAsKev5cLLs3YO+MAKD2GXJwLIHeJ3ugrUR
Dv9kh2OBTyE/2YSUvYYMwi57IVBVNFeDNO8ilzrC8SqBw9FgltbsdClMuImMvnxB
dSld/rs42gvEZmDtAsoThfolWnj0BnQWuKWz511FqN6LFtGpTDpzkkiiQQ8MOb0u
t9heC9qsZhhTAZKkIO4irJGtQjiDHyHq4xtMmVy0X8Iun++5ivnaggXrdukEFXri
eElYT6hI7ASj+W3194XCrlgSITY85L8BI00lUjls9vTqVemQLbFr0wEXVpxWF/f+
ciQctQMPlM2dsw3i8VlM/uDjgkPNUFPyCEKr6OTdTiaSY2wcOmk4Mn8u2suR4l+w
HTIHpaD+ZU3S970xqb/TtmdtieZiuz4YC5gt+rQTro4XEw8jJ2uxZRZ+2NmZ4XNj
4WqDSj7hrkUF6MXPJNBzS9UTf5JR7XPrPJegyoXTVBpcbMs0MEKjTENyhjwNONGo
s0cvK9RhEYg424uMVTyLou4pmk2snE+9cj10UxFbtPn3rewaIKOZKk/F2vSoh6eh
xGXl+Ww6fmJVKQ6ljK8oo0gxPfTX2A0a/qh/KryjCpNBE3fR2q8w8CWTvXJ0aLzx
o+kJvbnIXGVRZ3KuybmdNyvX7zcGaTm4o4vTkm7mAjUa/4VzmV/DhPvOXMXGczWQ
oeDH2u6jdnx9OLOIYMFYJvbMTM7N53yukiBYwIrUK/o0913Xl1r30gqaBYszpMhN
Xx4kbq31xrq6dODAnOOP8f6r+YXiwLq+0/+5pUXvsHVbfsj89vUxdDalpbaTwwdP
owZXAHD53vFUs2BgdKOSL3Yy2pIoLEm7BqbMdgNJP9MWSQEpNP+ZrVF0WX20bNF5
DJ1UQaxVtTN1/OpAyB9bJQyzv/1X6Jo1oCLqykU2PUq3qqHPJKD03XyE41JhdNjK
XlT/238mfjE4G02sqUb3uZuRSvtahBj1tkMZokTlJtoj2XYNpaxsfcLhXCCAg/6L
Onc7IYtwEAPKSGH59uslQcE5zzsSobn/QsZHeCufDz1kJYIufAeg8VjKOqN0RGya
KuPK2U4sok+ITdzInL9sVibg+1eF/LLXwrfgaz7yn7w2RL3HNowCzrsUQuO78DhE
HjYgtEt/weZI4URdLVEG0S3YDlHy5LV31LwnCYz44w9kksxSks2ivkVZJbpvqte0
lBVfd2TwtegqA0miaxtNY9oLy+R4HFGMjRLUKRQKx/0UtNKN+bM1D4afGmarnwlY
Uh2e7VVStqErJuRp5im/G3Z7r/KeRrxtLa9rp+oaOp/rvcwZIskFy6oTKNEyk02y
JM6Xbb0Q11UbrfwmFTzdW0eLHRqOJGb/wqgo0oUtTQE1qSAtkD0PKe4GkPTnw4eN
qVnLajgly/eN1RTVUNkU50253XWWH2RaG2gJkBbrz+PrX+WXdt5eeXwLT3YIVY8z
3bFq2RDlGAwDd+vfr/OagubKyRM8TE+82WaL5vwtArF0Al49fGC4YmGZzW40tbbr
NUxctaqTR/lkWBlc7kKa28YNf9p7PajrJ/1466y2pjoQhyqWMWzufKxUUaee3Fxl
0FopDFbbfV6n+PA179L5Dg9i3v5En0a5mDImg615QaWlJQWWXcezdovtp5ebSf3I
JittHf4cuZhy4xcIrDWE/TRBeSGZ74p+WXUYw3tkJwei94gvEjlAvi1iQ8hyrPx8
P5C7xIhDtQKdVY11zUdiGDchNC+GkcykB+kDoTpBnN3VeJwjH8mD/F0XxqNN0fEd
c8GnwUlVHgr5GFSr+U3EnOobLc6clY83y4zkR4eNhkHuKrI7vZmgHs4n6VD+eB9J
wTWdfe7/gdMBf4sfn6wu8nPK4fd9P0qOeNzhqg2OCkSnoqURi6UhBbX3hx9ka2Ts
GlnIN0lUrc0hhA0nf8kMI8EeG2ODgC4dnWcVkNEd6snyJsx1OWL2ggLxCKNbDWnq
/9QaLiKk6nYqSMQRvowdU4qrf+3xRfiPispn7oEatgaXI/fFgKSeGtgpkpEG2Xme
UHRy7rtMaGGTLyk6BCG6srylNFr/3l9Zgpc47KIFCdTX4wxNrKB9GHN4uaBEvBmV
iVoGth72oVQJdWFMQU0ij5P+DBELOt6oLRLFs+LWv2PAQl1+Lgn4TPqSoLKLT2v9
mSaRNu9yR2YxMPC1guyeZwIM4pw6iyhPR/cGMHnUEHur7fXg1URIaPXFs7WPU8W4
z5ksyPP3xtzRyG+8Fv/m6hxG8WYRPDto3DJ3y503vg1TI0ck76VESnh1TW5Qji5R
+rjs+pSn/Ml3hF6E+JydpoyNcjc77U+CxcNXtePNcUuCo+8cOMECCqQgBg4gpKc0
0a52WVjCMOY3ezDWvdQicbAQnEw7iIn3RFuy1trNJPGNto1P1tnLdQf8Zg1bk71v
Hm2UcTTYBnHQG/Ylxho6IcNUVG9sQZeHY5BipsllHSEsse+i53lD7nILsU3oVViK
qIuYbxTQmrr4G0S8eou0NOexeT9Qw8aO/EM3c2ifyPcEAb5Iv9N5YjtueoAeRtm5
tlasbKcv3ZtFkaq1wULKcAz7ER6DwDZMR9DUvkGCzV1kD/QFywAaA4a0kp0FIkDw
kXf88PfanFm8QKqSzu2GChNijDFudnsifQY14uJ2B8XMDKI2OWnYLdgyvn2W80jG
uuYDpl6aPyDbik4Vbq9L6ztmnrC8fVuWdZtKujBcZly4WDoxjED5Yu2l42BFDXm2
mC3rz2pVC2O0Az2u7u3W0bAFHr4BfGxZlcs+smB3xXzJoUzw2M3O5F73ZCucHZzE
p1R9/nC7z6dFDHtOAxwZBZNJAQKYnN8dnPLvsycDOkJOs4yptIYQOS4hEUH4WC6g
qply8EKmhHmLVz6N27Q5g7G4q5Nw6wqxnJxrrVU6yp0A+BiKPHWG4AFGqPE7Lp0C
9qdptYgfstPDOzEh/D2zrwif4rLGEB7BgK/gZWTdDLIWSfemTV3AtrrFGXovVe7Y
Vx+SEfAck0IWKl797okeXdHg9NgLCDPGV+UiXWiIg7gJBkmMfVQhA/MT73bYZGv9
q8MwDs4XPwKp3l6+wh5h2ByiuSaRfXbDoPem2oZTEOaEISZtmTubdxtzysZouq/B
isy3sIUKMvRjkfWAzy85CZY7AibcR5rG5sajt0+gnE1acFq7Hum/2zF1MeNstYV0
gZbJ+Yu+vLSWUSmqfJ9tZPbxyo58qvvB42039BVLkP9F/FakCWpcBtfdrVkz1x+X
zES/nWsCn1dfnrUQoDs4tUsrH0kTn2DnVMv3wYJmpIL/gK74R7NnQK13MsVukxuL
idrDsuW5B0+E7Wmgcnt+op8WPfJapcvt8kxEHbujPFd0URgLIZQHblq2t9VSRu8M
Xo9c+M/oc7h9qFNajFr3bgvOucXEbvM2vLOou/Xvz69GAqoMXQQdGj/t5+Z34Ezf
jCuXR0IJwcIBl271NVIfDeIATea27+aQ8Q51nNQtNh/BTLE4vSnMHuCtqN8w/J0B
jH7OasgO6dFkNWPO+0p63Rta+bIzWt9cunPWmu83TWMQz0ywZZQCbzdGLy5aXVJa
4QmCadxPRz6gkW578/+UFSIOInMGuAA28PZzvP64cDxkIOj58xeBEkvtwVtXb4cN
zlCmxUvcuzQnbtwWuIMfOn8mtBOl1oJzeHq7mUATp2Q5U9Klv/utIlLNbuCCWGv9
kzXrTHs5YkOL/TxA0L4MQ/ie1eb6dNCRf2AgKbmqJfMPpPfV1bzTupS+02zDc94v
VbLFyfwC/TS+/oELQ0mJCRFBRQ9upmN9ODF+LXDc+Kc32H6yYu/1R6h02J6Dihqv
PyZTsJhHFay9tFktE+DlfVTWnyHtNxehdT2FGLnpxAaYZ4xoQy+xsN14ZgH7r9R+
7iFXVEGeRtrtdHmdgmOtaVblsVXaxZNXK1yhMoMSFd4nr1vq1MTxqxJzvzesfcKb
UqA3KgO3t9wU8ShrSxon7tFNzO1rn4rs+MfhutCbPtqlyRSG589k/7F8cl2MAfM7
tpaE6UJLYej7rT3JufcLQGODahIqjCyBnomN1FvVAbjSfmgbLMrtA7HXxRqSTI/Z
tLBtaU9kyG6bwqb/F82M4g15m5p0i56tKUR7QJzdB25+tpbBtLkgXR/LALihITbD
S/TZiZTNbrVDS3XSPNvJvjNkXEIwjUQ4NomPRo4Y4rhPHDlmKuX3tom6DKrlxkT7
52p6YA4nH5R8jZzk6UMWQYFBKRBYMFeWhG1ufu1djAFrwQtVExUirDKgt6r3GqrK
L/B5aJUneiDpG58sqTBTMOxPeTF4DDQ+BONMzKIWnUX+4dhpWHtdQg7GYOzvjVar
SR1Xrpy+6Zklbepz/hBWDOZSDMCt53f2RNu8SpJavBS7fHf0qnY8/QoGSYUXCzOB
5qqx0eqfWSoimTc4gfIXAonyfMTNR6WKEOGk3nvbjzakIT/Prdv0+O6neqYj71Mf
oMGQrKRHvZRw4YV5HDjwZBs9znLYCUD36QczFvyRhPFXVlYal/+COaCMoN5/wsAO
69ki1gOM+/r2tSywgBH6QqCB3qNjlZmnRLwlkrY4nLazIO0ImTolKQjQ6SaH4tRm
b3omv1ocGiLGWrRIEVzdfGfh4jG/xxMP4EgJnd8iHVeMKuG4rqTeXxLNcnkz2tkT
54qaHFUGquOaOoRD6J8KIS96rMlTGbaw6EEPysSYvolI3Wj8M/UK8sFZ9+O6hq7a
6A0/jcBPiE7F8IyN5l8mBNQTP8uiR1yKZOXiN7ifQJGBjEaFVKnne0MscU5pjHpQ
wXnILc+lP1JZay4VZldpcSkSAsO4zVGo6eLIKjvADqIPypVUoXaNLTdwdRwtv1xM
R11601Dsc+sclcZsd6Uw256oRYzevr5Do5GkrXLjpgmTH8qlECqfLxWIRXtliTn4
4Zx9sxvXzzWZgIQ1czOFw0MYnETjscnGKLO/Vmkp5Vcw2kG6wRYSPLyzuvZVYhmg
5HE93Uo5T8AdowtQI6Nel/GgwkTwelpc33XSu5WS5BZ/pq6Elf6/pjG0FVh48cJx
sJyT31r1Fe8vdP3MXTo8CVdVu9pfm7ED5+gjn8Nd1uBm9gLo5+6Z70j7EwBrnoJd
0DAtBOYXD3XeNHPnXPWZJZ4vMxAIHk7xOlVPaZHYKph7XKOQs+rlSJp1qbrYHUhN
/19O4jnAdFkDoXHT7wkS4dbnztFYz9aWeMq5Cj2iq8o4MV0EpblHMpfFIIgqwufF
QBWSnzTOxNgunGOscuDxexDVp6FTCwP4a9mjiX+PAqfW9cKeOokoHhH72MX2ip4W
fOJLkqtDTanOg5ExniTjgMb9qamDQ28V3EkFYfObf+SUP1bIz5GmnH5Ae2kmVWCw
tDOW23Wk+NjgzNdR4zgXZpE4dPJWqJxUiOHniQFU1dp/GINDfndZytc9B1RluAqZ
pB/hAllukrxyAqnJC4QYYBBUKQTSf31N2fmvq01ckduyqwDYxkz9lw1aMoKR4r0l
ie2z/6/lAphs6quowncJdoJRInGSAGYCic69jz9oCuT2lBtDRTUUjFIJd7PpHx7R
h/fC80C3ux3sA1lWSbo72Y0+OoMqiTTx+ng/2Air6b+X9myFa7YbfYsnb/LPLFGd
XmralcQbBKgH54WNnQVM9MRl/JtDRBHXayUDM3YDcyJhLgY/EZGQ4OV7brV93OIy
t0zEkITxDmmUhKo4rdK+zXCSzo1UjUVw960PMjLONUwKQ/kBVXglVLG7S2bJ37Pn
KMMMrURPM9Mj2WrJDA20S4yxrM64hx006yjSasiEmK6dSblv1x43n9zP6xKvpvu5
hXCmxnpNf9jYO0qlX3foMOsG8OgDA2Do6TbkGsJe1OWAxkXIzIVQuaddQEPBPLGS
CxriX9QhtQ7NMSuQSGCOF+wGhUehAuwIyFqeJboJ5MyTTJU+yTl1x3nYMUHMsTa3
Bq98cpDRfLcTq4hYqnPluSPcnac5MJSwj5ICZ4A2/GfntebKi6CfcjATmP+hXt38
gjUC1cEj+e4Vge3ObXlTCuugbMp6DZK22+fx4Yv7BUStROK68BJ+hrMuo1W2Kjcg
1wFEgUE5VZK3u37VAoAV3IEQR1b5eMM3T6nc8jV0O4AxhF7gBqxRCHamEh6Lz094
KsWt+vUdt7ahxDUJBipyiz53+cjDdUeCqBBc2d++vzQ+sDDe5Ljv6XKJ0limnAqS
cXbLhwwCyxFK5gjABJbsU0W3pw7ExhzY2u6ZuV6mCWpKp71LL/8ZHaAZfGsA7uIV
uh02P+ihxFl10cV1KU8wqAmQL9g4FjPjRvTk3E3Xw1NWyly0fU9fXLzYb7zqzF7U
DlJI+ZCQ8gouBvLmubncziwzH/pNJ0DFfooiNFr7+QhIBN7kd3UqxWwcWvVCQ8Iz
Ut3U6NnL50vhvWDQ0lYf7h0IqQ/Zgrmf4k3YIjkj4GZIjCCKS8KN/2TZuAmu1T2w
dHZFw1bmSIJl4EwEvTS3dWq0AEYQURAWcFyARFlEJ7i5sm2C7XcVecHUowsvTx1r
aa+bghC6YVRwTyKurnOapnyEIc7oZi/9K4FIarQIOxjFwvsvRgKD8zzynA9wvObz
OLYTgcKIOA+IkFhM6zCPauZP2UIxlSA+y7HM3iOGc/M3FKnlg4gN6g+AFiuwG1tE
T/YN/HZ/GPglqfB91u2sb/uuyw2wG3pPJJtqaaf6+xfi6C32OmxIecUOBzyp0pAT
5siwBFBzwFnCDo/544WXQamwMoAgSluByEazdNTZdBJ0mMub9guAO4zuBojBk/U2
wJ/PiIyQRxvnK6+B6B2yfMZRiU25bMY0G5bDJ5Evtp+i/QtahokSvhJQ1c537cYz
IllSCQ+/5VzUXwTuYWoTIfUeIRqVk1o+qKHvnRmD+kSrgXT3MHUtK9T9E1Ay/Y5G
lrrIXvhc4cW9y0UTyZwqWFLI+9R02npwPM8W1dKQqoohEfhqtHEAewdmHHugAXv0
NtcdCS3YshBPzjUpUEOmOAOOqIhjpjvzbOSVuT4vbrSytlhoPbC2HFvzQ5mC9MdM
Dxl4Py031qNW2gAfQARvp37iBZLjldRfe05t+0Rl8D7ac4bfH+MO5FFPWUjfJf92
DgwZTbpvulTVFzVsp5vajn5BOJr6gHaluqxacJZYPV1ccpuER80wWDRpQWBuH7q1
J4TosqLz+Ikwm4s6vhQd0t00iTObVgSgBq024LDnF9SnyyBJRYK2pvDU4TiiFc++
350schlkMj2fhlg2M265LGAd+tQPUsdCQXwCJZE4pCpMCaMGsR4e6WPb4d4tJzJL
it6yGclgY0kVJkAygoQGEDOI/iw8tOER+Nln+L8QByIV6TTXNy44RQpXv7fbmjs+
Mc1h1TnoXb4aCQqLFPQ5okSuFtRHEs+2H+L1bfiROsnr/czOiP7J7efJabaZ6Sjg
N3xxfOAOZaDRHWy1Za2CFuEj9auEI6mlhtiNFoXoVzdV5jqV+7ptx/rqRO4uU13N
tAkzeuieIdcE92awMZ4QCD6A7ztqO6wn3reFySI9gN34eWtuC2pMMpB2dF4HBkw9
ZCwEuBt4G2CgIQLvljFc4OKFi6nRnd7szGYxB+hEq3E91rbcc7RgayUYVFgWjq41
KRm3WnL3vlgpAu//P8/olEwNnqvhcUj3mrdM7dPuIIwDUmkPx6yFNRozqU7VbW1d
G/LWMzLyXxF+EAm3TNt98rafrHiRQd2o/+nhATvGYZoEiUod5vtkFOVy7j8cIUsm
ud047EcKrNS571nGD0imbTYgCpSy9+zukHps5G/nXgNUpEhV4wP+URx8eUwOS0FG
fDz48X2cPA1K7xoYqVApABtdT3lxhY40LZoKws79GTMmiUNg0oT9bC8NM0+ItDFg
jgkqY9jFhScuyfcXRqMxGk3lEiX2nrkTk59OkHEVtkeRPbc3wJaMou55OhJ7KcDM
SVEAZzNBp6+aizKBksThT0mNVbCMXkFhmAuu27pulzo+RO0RTMT15D83DjMDRnt3
dkc+gxHR1noygQ/ydBdEiiEk+FxZbEqcPiXaztR5ky1uO4HPi2/0LL/21u9123vm
gb64S/XIXRrAqHnd+b4PB8L62gcjI/6Yp4hgnd2AFh5RVVKwziSfVtQae7FlaKUM
TXSwvbdd99MojwoFfgdZjv1IZllTJ751+ywQcB9tOzK3Qr3P4jJ7+PJI65IUOvw+
OHh/E47hrOq3nmT7XHfL26gjIJYN7gQwcFRfpXUGvpO5EpLJd42lEg3A1dFGJSSL
6FC0wlZ3o0Sp8hedxVVI2X4h77uKTwqr3MAlMD4b+UXBrbrIWXoV6AXvLa9+Mceo
LBR7Jg2HNA+Ys4hjnUV7fFAfqcJiBkJH1B3ugJjAP7r1xp9QjuWsKHtTHLdVXeTL
7uXYfwT8YVwH6yEVfYFhAVCks313qxICZyuC4CkT4PhAr0sNmElVj43kz+CfnRPD
nVoNsBAnGsE+EIvMw941zcO6OLMNd5I19zmXCW6NbL4WM2SHRP7gMNTxen17qXab
Ah+ctn37m9odSNi1TzGHOqb0QufFHH+3DpqxSdmpknwn0ia0tnGWsL83A4Rpcwyl
uKRouTiHVDp76XlhvUF49XAagmneRpnE4mG7XG3jdLImB8M0HcMw0q/FU95K1Xof
pJAQlYgvUpOFQj6nbY3e7khN/1v3GnjDNhEiynxanKpmKpX7lu+ZfFASqUOe9j70
vJz3bljbZ1RwmsNrV2d+ZDBAFLl9LNsr0qmgORLraEWl836X9YyEQpbkgT+CV6+b
jY7U8AWYyBt58j0QepdUo9A1n5iRMzX34lhtG1fK5nwHbJ7BtwFaB5bZiL6/ipfP
y8ix/dCCbSfxNnxOY0y7sLQW0AN4E2lnKedzMYz0Fgl/Xv52TPXcw2FXFn1YQFnl
2frca9A29kypGfQjayhZZ470+aB0IaSwvhzDpBKZi8fK2Y8ypCa5nYNyKwZlhuls
36jjRevh6r1lnRT5SqxwX71UM6vRon1RuLVZ9ahvOWAto/68Aq+F4zL+Pahnp0pF
PTQNTbvGzFX1aoCyki8Gn4OI3Y/LnHz+/YUz6s0Ywc8c7fH4qxRnZDfJtWOwuH+W
3nDhL0ph1LeW6vr1mZGsHNRPqHYAqfPTClQcP/9EtFni1dKo1uhhhgsMKvtfld7w
HjrEa7jUB5b9C4Mu6jAAxs9NnD6rRCP3cLzVoqtdBhuLzNVAgVnjd7ZUELxO6IO1
T8dFZi5D0Xad6cesoDuF01ObpJ9qU1hztg8T7SGXUi6++UG9iKIInZ7HrANgnfmS
28Qks0W70bcGQqDnz3agvOAOj3BKFUgA/omnrQm8T9uaZZ/u8If6UxHcfcnqTpPA
FKeI3wScyI/RuS8gzSqM2HSRiAGT9t7Vd0quSOW1m0yOhNAxiMjLZLdXG+FN088h
fl/4Symjk6hSsxn8muqKf1h/RaRF9nx7m0SopoSrApYyeOKM911BiNpcevyhsBQp
phZfui5TD3yfoAaWrzTxvyeVdnc1LVDaY1J5vozYS1Fxu0Q/N7Iv+XPh2bhvUptt
s6ES/u1cbblwvkWZkdXyOCKOYTZYEEjfClAupeyRsV0zd9vmiAFdUxmlfSgcANEN
kQy7m+oack5jquyRBIxCC/mLxIiL3IdkaMJ/GVRjGTXj9QZ1m9EI1AFUP00RId8v
hEnfxVK+1CIgp7H+nVq3M65lyJJi9OEYoYGgSoDtOTGVIsKopF7j7Hnuul2neJVn
7Hv8spIjwK4hsDoTMPex7ld3Ap0wk+QoF4udnzoi9yc1pjfm0F7zt8gMkKOvfz7H
W6vKhXskjZkBfW84P2K+e5FlMVF5GHO57yG3eRwUPWSDWLfcRD5wIB5+xTgUoV1+
atph1zdapUH0wqSPo2laCfuPL9jjnZdIcwQ6Uxv0Nf3e+vWTv0Nt/jeLmF/r9xHY
rf2b1W6jZv70oTiXKAWPAa7ayDgnqsLs12DMTlBtlBdV+ozKCo23DXoVhD2OHKA5
N+PPt2l3/KyX34hVvCFQTJZfcgrZ0FBxRLG22v/3In1p8TfHjmwkVWJy4I2Fg8na
wMwkEtyA11V4hCbvzDg8YCIIJ7RLNLzyAJPoqN2GX6aew9m44ks+Zanm+7oJ5g02
VhHz8PX0cVQDGCnLwdezugMcndKkQ6Xs3MnCqvGtmgXDyuvQS0epiri7rLze8U01
WWeHa7m17kI/chIjFi7lxeYB9IdYGR0vOxZGQNy040jD3npmgW+2P8N6kHGfk3/B
xNkI6zsw+r9F6547Dc/LHHeINZSt9iDC26K3H8+cq1+DsWrO78D7+pugTqDXdCcM
UfL6eB0Ua9FBu0DNLgG5zFq43Z3gj8B+gQ8v0hgum91yHVyZfXqD9QKmeG3hpxkU
sjGTUfStnW7ov1hJ23KzrCzyfHX+y1oFWiSulOaOnx8SOjFbE6s/Hiq7kvzQU8zX
yJx5bHM3EiQUq+ejhJ/jVKZ85QdAu54L7+Jw7/TlCkmm3g/sCHmz8FSIyWa32ZPo
tPjkGSOPKtjn0GcTQeptnBLW0TEFqh5n0oG/29f0bDsakpczAEnemK93vr9WyOSr
HSiI9arxgN2Xazn27gOxrld0nce0GQidU3j9/dgZvyfBRk9SysLI2Y+FqAxHW/XS
b+woc9vvK91rrgPxAVMaHXk6IGbfWXSg/xuAEMFfftq+sRaydQ8qxckK3oB7rEYw
pT5rAWGuwEENK3ULHJsC7tzBmiuAD+AdHNXlC9h5MICWpGmQo0899vjZzxSMje+r
IgDqXL9Vlf/jVCpcUIErkNM9hrVwYzIGXkaWNn6DZDSh6DRcXc9CaMYGAKa4flTd
ajpat7eB/E2lJRfaObI/T7hzaQ3y83TtOEUQve7TVk9WUSmNU5BmGazKRBDin+NN
hSaM4qb9s9GBRglGqtvTdsvyPdT+/7mIV4NU4vjyQrgsj35VJ4thgzDrSO5FavDC
O81zBDNzEkhSA4/uktcQixQjGZGsmatbolnUNB/t7H0+e/wcJDESRn17FA2Px6gu
LLsp0BXLAh1u3eBV0UBqHcWdwVL3k3QnZnx4YlgXq40e4L6EZ5bi+FqMzQvpTTwk
Blv9TcI12C0YX5gtr8pdyDBGBQ7wGv9rY1v3sbcn1z9875VRdnAf90s4QMQaDOQV
kFF/i/mZxHNQ/R8x6AX2kU0BQUYFWrJjfP9fJjd4wrG3cghIt9fTMM+awlUS76XK
erqnywPUHC42UfhvMmkXPtFX1+JeYvlz/x/+kZFZ8MDrHaCDVPMFuy3CZ9FA63Dm
A2vhF4kQHjPbm82FtRW6AI7h9FHGfdM+t/lCs6ualQylDJ0zFndhFq573/DZI4Nr
og5LbZla3L1jM89IYFA8MwEu5kGWwp05aJKWBuFZzu8CDOLpF6oGxl+upz1UcnRA
+qydGt9/TVraR6IMbh6lp3gdkXa3vDaJEFLGbfe/hqzuqZmN7qT+04OJRpGM6pkQ
rZrsiYONZLZA+zXm9onckP3qpLECtFzi7IE1iJEQuJ2UXX5Go40YJuWMTQpolp7j
lokMsJey152QHUk03hQiYtdqaaxNFRKPZLg9YCEgQ9HLtqxeTQM5EY3KwPKwD7jQ
ZHYp+8gn9Coem1hmOMy2M0ePZd5y20lCeGfF0lUp7j+/wdWxSlNYmIhGLTYXQJrN
+3l0/OnxLJYuM77GQJw9Q7INusIB1pde0i37jKdeFB85f0Aad5esEPyjKRMUnk/G
O74Undv48fXRetrByltzfZx6TlYGCU9FZvJKYfbXFzbvsxePQUZZF0PMYghYjMz4
GPrXwN17j4F8woQ6fuyKN+tF/AyslQBB7pzscsuZV0sVr2tXTjysPDiXXmM1/BjX
Pr39Hm/pKadwcd9XNAv935d3yhm1FwFUPLZaJPSmkhEdqMfaI4MMEUpolANbAj7G
cz2Pa0eijuxU0LRfs6+NW/Z5rqoHm78NvHhiMdc1nf7V6kem3LFdz8xa2zdnJ/hY
cv3EBeN/Neie+4B4w0r2KyeMFdVVHN3u7VXqTyWznZ/y6dFi34UuwTosxN2Dl180
8AAcL4FPoQmyPo67+/bY/yIc3RqO5PbD1w1MkFKB9qag1DbDWCkHMNY0q1I63PKO
qPEnu1YbIrjChhf/WcR0wwxd9g98Dfj29AW7vM1lVrp9nSWy4Ne3oRwPylBwNwtb
OxltGw+wecv4xWCj1pbAHrxDuWJd4hE1kHcKJsaJjYaFmpSNVRUe6fbaiHfp8Co3
uB10mJp+nVF2goXovvmyVC4n6fGSgiRkmwmyzKdQ3pypGGyfTYXVE2Jz5pY16RUO
dQ0r8cqz9CMaOQFjyVii/wd5/41JFPatISuRU1UZ/Z4K0D6sddMfzqbFKFm1qy9X
jl7+9s3v/jveWK8mhxH7v94wcUOwFN6mC0istovQeqhOsZK8VfyHHJKtTc1BsPTZ
bQz98NVpZBvjC7U1TKV5ISI0k599FSUvj2lohwNrLY0PakfNUdYv/nwuFrdFy2HV
HGKD645WddzF5as9W1nBn7+Mf51hR5pum/sryci51MjnACg7H1Z11g9TqtdYkXy9
lDlQ1zq3gde2ycnJtuLfAfumnL1fbX5040s/ELvU4eHt0snUB743ZDN+AMqbb16c
sBNcyH2Xk6B9Qcrs0MbXrZ3LxM1oFo1SEb/zHOpkdVsyXeO6YoomolcefouVsw7o
/feCFnupUKO+jbSQiX5Sg5qYnckoxYrNvOjd1XTlDgyV3b1gXiZqFZfseaRCJBqF
+tHv/sopFp1IxUymZ6gY7NSPbTlaSwxKQVUMe8cAQlL7Crge36PxT8VESlnnZ36+
dc6vFSdrDj20Zg3Hh8WUnWe7Y8w9BT/vFYi7xkKyTSyVCk5QEDViS88UkSNg+ACL
3EqIlwaU+egQvh/Uzusbep311S4258zNQ7BOE01HTBXf2GOjv1GrL9ux0/gnK0m2
lfntxtsKJoANHy+1F5g/TKXkW8bH1WcR59dQ9bvP03XMxpN+MDr1P6vq/1mZMILm
pSvR6HRuE2osq6vYPie274hJiLDvLoU4I95IVEVdneP9rMFuIPeKSWW5jnGFG6Wf
CAgGe7k9AR6WaaNebDOMiwcFrI7Xjo8B+/T/7ABmnFffEGUDbq+wDikwDdUO9KL/
Kf8x9fTUn/DZ/gbDSJ4IMZWBdpkI+hlaWBsMRb99Vfd8PNOePSr64TulrTNNEg8M
GHkYmE4RVsBcnZm9Uirf3m5hEuAvqJQFlmIXFamXZFKTgxTf+Pm1IcPZSi77ATGx
jnqgal07Nkera8iZoOJoAjqDoUERmrD+eSrul9+3rxBNfxTXmYEhnhUlzAgCsQIL
QRxDY6G336EKEgNvEy5e5UgzS6Wj0T5Jo9CXgzE37jXHy++9zswwBG2dcMEF6Ow6
XB9t1wGBa1gaD0P91kRbxcneli64Gjz3UQdFHeyqPQ7MmvrsQWykopd02hnxdNsA
JPiDL8naCW3oMcNJwAnJ9RditsQuIUiCxlqej+Vfzb321SiusLN6zkUHMKQX3yUZ
wc9P0rwqYTRNHcUAYLrtOBK3U0GRHwwMbMqjMEceLx7JG44GGhFJ9QG23Fy1VNs7
yxBUw4oclnSDFThqr4+54+IKGL2fUrKrQleVscqEX3La0P4Z5YzEUqGxbCnLYv2O
wuRht8BnGolFUV2R5TWBbujgbhUKrTOoL+V5+5TZRrjtzFJ5pe1aHY5bj+6dNN4M
9w1nVYHqRglK41Hsxif2odYPPgzsJ/EvfqDsHw0ozTOdWMPMO2wEp/L6Cp4UvC2k
fe28qhW/v/d7BttSVyTjMNGpPoN9JKqTiZG2e7I5ycWbqSDL3ZGzxCH/xkImeDyo
8FUQCdM/FnZNHDcDXTZXdJvASHZizxWADLajkPhxt1Rv6pODgDIMWI0LapsvOT5/
qd8AycvvPz93gqy2CTwDRPn8qL7frkYVJssQvztitmkKfu88aCaRGx8AClTSiKjw
cab/JonZ2kaWJBAEEMHeZqW51RIIh6kv5ISGskNcyvjyr55d8m2kD46y9utfwvJR
DWwBOB2xhZhVtHEtzq5lcx/d+Ji1pps0WQ/24j/btF04FIuyFT8GvTnfmTr6IkI1
7M97RDYwJEbMNojYXtCpNqaPBx3/0dffA8jdCItVRkRppEP5hjwi6g+aSxo9TJz0
XcAfEeMVRW0KMw1pqoJSYR+k1iMHje0GZkgMhnkWVHnrfIFTNYrLDqGtDQTzmhzo
q9X6CcCo+vDZhNiszgztR+8MV16DmUhlP5xjwLD0NcLPW7CzkiWNZsiMpTdHhIM9
bOe9mlyjWFHQKw0VuD8hnfEn9AS+XHrqWpMJCvUn/4w8rGpo4zEAgJ6CO/at5vIh
0h1fWyoJLthgo/IRXo48IE/MLqh31rLI64ZebpHnOT8QKs9CJc7alVW5n2NCyqeK
fUc6IFCEIxvitKsNfYqtG/fR7Qi6GTepLTwitNS3C4VF3z+h+rc/+4yWOaJu2S9h
2UdjSj4F7jmKKvN+3+L9CQb3ow6ZTE97Nj2kHy1kLVs77+sGVVDpQYI8hg7Ucu1Z
i3WICkuL3eEqKb6H6q1Fey7fKLn82o24o76lRMKj4+jJgD2UIO4l3AhdBitErqGz
IwAcgtu2UqFiVNemsjNX0Wqm2rQewQQ9Ma8kScAnOLi9/rDCPwhBy8faBN51GSac
N0EuLpOyZ2i7IShmiVzhKfENLvE3+2v6R+sxZ6g1XYiTpbzjfSwXX7tR38WqGT+Q
mwJneZ1C7kQ3OPfv7UxpPqis89JkRq9fvWNWB2FxNKxDe1yFwdijivqkfpKP8M0+
BKU5+gD/nZK6WELUuMRczj1xkMfS0Wbe8nnGRG9rUVCo+culHmNVcK+2QEGTb+Hk
KslKcloR4zv+cCJtg/+2PdxwzCc8hg5WxG2NusdWphFxMVWwAwaqxIXyJnabhE1c
/Hw5CG1FKDZSvbhOyISX7mzlmjX0g3+R1YXUQUaRrsvXRkL2DcqvU/2xpZLDbKEk
7VDgIB2ZeAbczutBdBq/2Ng2iA9tKDId4pbu4qunsZkuchAuGoohusHSTZN74KRM
pJxWsQpDaU1dDV+2/8q85IgYeMi8Mmun2CBsocS90HWlF6gofW9A649Q94EabWCb
p26XxPR5sS3/JKK3s5PmmMGjl25TSCd+JZsIS+FD9QZqJ93fDxVpNtP4XkHcryvZ
7Y9BKOq2GnoD6kqNYrJUJ2UcYpsaLQlu6Ar/Bu2TcQCRtigszs/Cd/thZ/AdgtE/
vIV2n3B80XqjuO1epAduj9A9wlwaEvfAc5eR0fH99O99PrV50oa4P/B7qoY1tUFS
aAfz4T3q+uhP+49xm5fUFGNPRHAm5vEhZrdOWOlHJLsw9hlJ5n6zLJI6zc4KKk5K
mJIlXOP3KQn9XQElctR3aDGhcs0IcozIfZhzUj4HyUjxlRDF7qnlE/Pp/H+p1NxE
qsqO2Fk41w98iZac0KwJae5t7bCAEuJ1jwmUjjXVNJEx9fhjXh0y48U9h9l58yy4
TBvsIhlPRmmFyA7pPMFvUb4/dPjSnC14HJox9qQFMTMXCOgR5yJsVuJ6gY577YNl
qyBDptv0f7Dta1AyRw5zt9BQVKOVcL2KmVt628SUlgzDz+HChyF9YZS2RjB4M1Rq
UJ4l2WzibhhQ7lqqIOz5tcZSgG8nuaihJvVw50vD2kwfK364cyLKfgBnq3DzbAUG
ufv4IVYfCKyHHZs2X8PaYhlsQpBt2zYRvnsYJCKILYxfL96ZPRBO3ft085v+N8Hf
s//NgqGoioHMrB6PRdmeDJBxbR5N0LCAOJz5ku7E8PqAqXgZyawvR2PhXi/0W/Bi
mRBUHQMGA1Y1WxRG02Kfa+QRp2jw1iISSxXRzSz6IirBuZmvnUTekYVEcQpMySA9
QpT5EfBRcYb741hjPSU2o1YwDJh2mWtsxbpvwJB8PcByeq26w2aSt5w/JHpe2A/W
69x6MY6kUEVbLpRyf8APhjVLdXBNriJjr7vfVPiZneYrnu5+PTlY6TsVykZvFbhE
KfO2ZiAQfRwYyuHNKI9+hZMK2oqIdCa2y6QjMh7+r0JMwNq+1ihqBBj3SaPK4vLE
eTPMqD/a1A0wEG/tlDu2jBfwCvTFwmivF0PCj4ml9plFpLSFbcyLYXnX7BKclq12
fjqZC8n+p+hAtC0ncLfW9OkftiY4NJ6X5iHogaDH6FXpWm6ZCE1Jq+/hwCeMZ41a
RW2yPUInWYRTseHTxOpDdbRI9RuQRId3VITfr1W6UBDWxHFNOQc0q11uARgQ3LGQ
5xljMTLyFEMu4nqVzNHF2dvBldvBy2HNGZOvcKeqPHNerOb1nzGFw1VZL1QHBrbR
rpvpmW7tHn2G7al3nZ+XX935/Jcc5aHs4c8w+NrQ//NNj5A1LgEjKAv7rg+6lMRr
GNFMnqZ9EZvTHNmoPan6ZMUqd2beVyP7r+st/OqnNc0tNBIO+NDEz5g2UjNG9tHv
tOuTU1rxVnKv0JIEvhUUDrt9xUKquIMPfQOZld1hh0HPJGk7y7CKtJ4Z1w+f5QJj
KUZqg4kV4rQNNPivmR0hzGGnOKIFjBzEXFuLwvX87LajCLZeaUmWxBopb9x9di9I
LjSrdVNt68Hd6xfb+4dkHJzE4ce6+n85sjNuAL5eNcwK/btkEstts7Kj9cPvWrTR
u7Cavvm8FlESL4woW0CjIXp3Y7IiDiXho+rokhYrklC+lwCh4ncpBB2AEDPLAbZT
zs79X5i/S6EHkS0WTZ01BJFW4cDwUEGtjdbrbv8fQwgGNPMP3b+fvpURh7txOr9s
ywzIHn62msIACpWOqkP92v/doydb5AiH/pKxeRf+Z5PQkeQBj/YLRjppgYH+fcEz
/O7amRIXpRl3uhI5iJpm6xTiLlXo0gdTwbjye11ahBz16Acq1BBq6RpSRLebnmiu
rl86LN5w7AsuCPDj28lvwIly1Ob1k3QdueLwhsqN4VbFn3LW68rqOXrKRkAQpobC
Gua+57MhwJLzxpXZ3Now7otaryuirpLqrfKsXTyRaemP/I+sWO/GTSnzsnM4sYtX
YNDYQyF5bpMQDG429Z+OoDocXMx77mJb3r+ArgCS9QAZsCwpG0aBxuhlmUjVrJU7
5EwCbnkiOWf7cgw3C0Xm/KliPd0fk0Go0QYzG0Huce+rdwLLf4X+O/hzPY+URNcT
FVdqADUxU+dwhy5ufTFfj4KFHzDClefOGG7wozfEEy2JEf4cgc9/iZfSRSvxUhVp
GOutobSsmFd4pB6EILGWNiLVP/ntiLHhNwdGc1HpPTDJHZeexIsRU4DP9WT2tWcf
cfPAo1YS4IYlOP+hfpQndEjdOKpJxONOxGXWBPNkI1yIS4XB6aCSWPpcnxtfeOl1
rKKxCt8hmOKWRLlGhNExDd7OJ0enXQDUNjUjqtXzETxoDGNHMZclAmSO3UxeLgcI
Apl5G0wLhlhFzCHUcsjOTUXNftKS2WhZOFmNRPH6WC+fYjHul4rI0EO/u1j84b08
3QOKxdh9OKK/H+jkGa6+oOFxqENVwihBGWqWZ8aHy+CWfPA/TkN3W2IuMvS1aGbx
OW9c3wk3D1ytLXPpOUQ02NzVlmqXIYDdfb9N1ArYzqKpgxKYJLVXWN01++XemBLG
Bc0nP6eeE/LNdAVJI+PnBmWIlUaSOrU49WoTA7HsKw4q45aar1DhCg93Jb4ZA/bl
TGW376ZXxkeHAlefqeHV5/T/rFOJmXuscaAsA2R+jUW9OXKtpH36vUSGhz4mf4Xj
QhPFKhtQ2hoewApN1JeitNgkN1sLpdeEZNP8u2idjcts6dbChecNEkCF0QPYZScA
XDYai+1dhSpwinzvIpI28Z/lCPU/mNi0ym3F/Z7q0+djyK+OUapuj+gqmrnZUpHc
/xwv+QysAkujlXJFCQv+LQQnL8mwKkSnuYBzoaVIIbV+Z50tPHdBKY9u+lNaAaBN
g9Ri9Y2OvLGB6WIOmjgHL/Re4ERFumRKaqSXbEqiXmzR7ORVWnWC0SO4zE4ANpgk
f830fXlvyFnKXt073oIzISOBFvZAEBGqjoENU1TtQrrJDo9BXWerDsitzyO7G9PG
rtoseCdOaHEE83uylkFZ91CWx7NUFgsPMkoNb6R+UvwuEjzglAXztKdd9C1tL3QH
Cai/pxlwL/7eHhGR9ccNTki6DkmPcOtL8O5y/g14CPdcQH8Rrq6dC0phcnap449/
evQ1DG5blFoQedaySoTUvSwWCHwkusCVbQhttI2NDuvA9ER1oRw/DPrTgnmp+7cE
WwepOQaXRcsDPCn31H/gZvNeEiLHxMywIDt7pXqH+KdEotSQoxQZ587xnWmjycBj
JFvbdbbeHwkSjpYUpDEVx2K5WTtdyOFD+cV688o/aOTtylB1Orjritym/eQiT427
CdLJBrNnwRAj6sBJCIpfe7QCGd123mt97SPmndC7jmfnswo8ksGM7xzFXXUGhcMo
C6ABZRc59QJUK/gpFDHFRmkPfe9JFEH9MMfUonmMvu6yz97POvL4DxGZpQBVnVX5
HXpzz5fy40OFO7f5pCwbLUgPg37p0yzfVUfWV+xotfAdKwjJZ9nZsNXn9C4x8YDH
Knrobd50kNxP1AbXVXOp0VSMOUskjoL/u21gtH8T8VDVrey9P7uQv4RahiU21+n0
Mp2VUVVq03YThvUhKUXgUk7TBTpGI5r/Y9nqup4iFgZvila4BfqgQ/IkBsb3j2+a
K/gMfBusC5FeC7d7/L/146yu6on9H+d/Ugou//F0hnRR3BdNUDD/r3ZDIuMBKqoX
z4dY6oWtwTJx1N8ComXZG/SzFwT5h74nfRdoS2nucDJhWFL7kWOkQn6FRgAOfGeG
o1KiyzAPqz28PoU4aGbLIAtdh0ZDVx4h/JLmGBh0JUPmK3cK1qU87JVmxTQ78rJ/
H8PrfPT6zwUtfM3FVOFUUBIBQ8zF25musohGd962XHXTIcfoJZ3m+h8ORUf1vxOZ
Pn1uvAIsrAxjAqWe4OvIJ8swrYG5Q4IuL55J+arj0bq4cOPDJQdU3YOoDj4BwF1c
n9nNpc2yNZFaasNGJd0r+yah/6fGqKrNKBlUaVTCotuegDpcXmkkR9UDnu6SUTtK
Pb53umYh2oUZxPboPPuO8gxwdbadx1S7Yww9YklIyOauvX67Z543IBM5N6NDWT6i
23LgEFe0xDFxVNW/zvqUsQgFipodxxuGuCIag1EPgFpFH88zUD2HgrZ/yQkBPTxg
3huQlIjK2NpAyrfqv9b8YTOqoFX+I9sqZugvOyEBtbEoqut5wzVHCWYERAlO8kgZ
ov5PVToiCFG0DqnDdV638AJPVvrpRxUij+XJPXzoPm6UAkNdOEHc7lNLIc6EtLkE
B+F7MD/L5xTTptMtnpj9hKTAkw083VE7tLrb2GhmiNgcpoJ5zFx85nSnV0nCsB3t
XrtLNdwNd0UVe/4fVdbIpaSgOdvMZ3/yVtcj9fEOvu1qg43BU/xOgKuD0b7gL8KY
cqt4tHa/+oXpyCXb1JPXjMBxnCpL6lx+YiUp5h393+2cvOenakTbL+rzLoOh9iKo
mbOgqh4axxvj/e56ip+DccTlyuaF3G6P4TL4xP5wdC1ILlq2aQ0S1bWH0J5AdyWO
G/Rb+ajW6fCvvbHzTfFgBqLNwNHE3X+P0ZcdZ5qMdQXnCsJcGYoTRqLDyUHABoT+
sbZgheb6DTHwW7GGf3oW/1GGW1ObbiNrXMDWwACea9s7JNKSEA19EPkotVNQlc1C
q3x7rKLl6ng7Kb2AfpLGNvEwi+4ORPQ+qH1LBgofC0JKTFAVVyrxwK7+CMHb/oIm
UkSd+VRE5+RCM0eb2+glfoOOnCU4OEYdO6lQtTmuJPyR7sIslTy2KOs01VrjZycA
G3rS8KMo4Hx4J8bsNUBIZyKD94EZKmSUb6n+rwQx4uomVwjvkZFPlC6RQeUzgEZA
41rHPHNObo9aXMYONZCHjAxKCnwpeln8WwA/Zs35nN289rrvkJNnH+OX+k0GR+zu
ptmp1tgkuCA/4QBGNv4rRSNQYA+LtKsRV8eK7WhEGfvCh/d+GmyZ9tESMvy63lxI
x9zW7vvR07Zao9MftMsXYTObVtewPsTP7zq+Aji3rCFY/snvtGWJy/18GlVkjE5Z
xQKYq0BvEB3yQCh3OnaBpHKNQ1xTPVeXW1lC2gCaRcBMSfDeN78uaAiApa/aOcOL
VLm7kegGUUQitVHsir3E87b7BQP6r4y/fyVgjQLWAyKA5jql1pKyqweoETgXw+ao
D8zXus1ISECLj4wG2PWIjKCz0rVPJ+D+iC8lF1w3KJZr+NhgVW3otmEysVl3L6yc
InOsMuzslnMpM6SMnWKX9csqHWunuKKXgpahXrK4t9GLBO1fCPGbPsKsFW/lbjTK
8/e8ZF7gcqrGqVoDau/xxbX73J9MTdH4Ltxmy6O/diExx5wgTpgIIqpBTF7kfMYb
rEgAx+sX+rZzPJaiB1R2UiZcsRrFAhQswoO0DKi4wE+KooZ/wuyWqO6pSIPeEA4A
ijRU1cMK16H3m2nOW4n6Bqv+rMJ7BkH63j70EMmKveC8SnIY2Qy3cFgxVu2ymQsj
CnUn7g+8iY+TE82eAETodcXNZskXkB//oJR+wksACcLd/vfKEGMCmdBG++Dn1W++
FamHMOJeLUHo3KNpjOX7jagDnbqtEVu24ssNSUccSkPoMjy1wXOyRL2B5oFScbEi
2iJOxtTFU2mXOxDjZEkQynQthIC2odJuGaWZZmtFLlOKf4p5x8xYCw0gqaMp369C
vPVplKTX0qGaXWMY44tguSRFSOR4FnPMUupRbAeJ3MDAMxG6aNGcAno2mDe7vCWM
jeroZRicp16QBHUZF82VmRfaRtQSEqOOe0DNhAWgnj7uiu3o5/ZzCFfASDsDaUbS
GQCyCCOEkpBZOKwsnTboNz1bJoGFx2x2nfkbHslzpu60583pwIZ+4c5l3+WBL8hv
DKDDzXboANNk552S2Lwl6wtuqaaLo4hgORs73X5/MisQs8xqnD3H/0iJ57Mklw+4
zMhSh12nbPd6ky6tVmzTMYxXZN7cIcZxF+UA4eoJ+eIrfVcrhwPepcwQIiShB97q
G6AWyj3jz8cPigoBGpdTho75AAowU2ZYQQHwCLoBmv4WFnO7XwD/xomV/Js7e/U2
I5GXQp5ANScGAlKO1S3mDW50MRGW8QyuLuBq7WX8HOWLxTl0tt8rgMv2q8aSZpf2
f0EvE/AJZjh54CuDYElsSKku6Ky+gaTJlLDShEbGEBZj8XLeqiLeJ6+s2KK9mA0/
sRLGJ8XQgergbY4lnvCXB7HVm5vy+qpRO3SBODIq6AuQc0qwZ7rBsjMIWjfMXUyA
N8QsNnO4B0bgFoUQjpx4CvWXp2S8JhH4288UZbziVnAVYbkJmJZKkxNt7XHyEgI6
sv/b/hVq3uyAPJxf9F4H82mLZK9XTmS+3Kx234cAwxSa5nYcCg+KcXDIPJh0Uanw
YoREGk+2B9bjbBGbjDQMNueiqLqtvL5FTh32U8TafoiSJZWYPu7EXDuQHoj8F0bn
i9/3RuwD9K6+ssoD+pcgFGbmU42bF4VE/N+hB5x873aDQH5meR7fZnK8y/flz0gt
bDTSFb72vdv34MLWcO2L3/6wYWmaEUEHidlual2Gl2X6BSnX/z4H4M0mD9Wlp7/G
1nrwaYXN+VHxL1LQ1woe/SmVmJXu5WkbzvDw9og0hXv5MutivnmvEkS4Ee61gyrS
5rYPyH5PXh2DNEqLUXvIo4VYGn6LmnRt8eWCca+fRvRK/w2xPBUIueUDQepuzHUp
yNsH+Hw4D69MBDauH8uT/ncrpeotG3YmmCUXYWqOtuI7CQIK0h0EKO6BL4hgu6RI
gWyFyhRiUy0k07sOHDSDuV0GJNEQnRfvVEa3bCFN12L7bU1WknwfiJ1FCosb4dWm
ukGluYLu2TgJqARwQvjOS/Sj1UWy9k4oufIOYDnDwHOtOs47DwMzH6jFVBwV4vlw
l9xunPeWXub4+ZGd4TJRQ8ddtHE7jOaKxTf3JLNbHrZDQYzJl8nvqS2q1+84sEyh
lEE55+BWKHk4xRQldHrZaXZLEGMw1M/VePUbksaNzFEOoibcGA034JJTtG2UA/Xf
uY9el0sXXJr6VzCA6HxnK3+uNkhEg9cFZhnfb25T73q8oa4C5RbN5c/wJlS2tyHh
X7fPEYpL+XlbKclJRrkYpjuzstD5Wh38d5owElAN1lCUIIaahJoJbxt8o1YO4gzc
BkgeW6BrvHIXt0oNFwiRRov3b8dDPot8NxGeaXiUZY9qJ1W+HZDJjPjl85UCkLtk
p7yHFYGhbbNJ3yz6oCpiRv89sCuHSPBKm197YRYGZostxDOY1yOC5MCvgM7ep2Bp
UWutixGpBu23xk2T9NGERy59hi7FBJcUfnfbh3NiaAg6o5XMFc/K5WGn6MKhnieX
s1BGyUNtI6Muo8mxzJc2vM/FZIWmBazG04nHBwAb9chc6/6htAfFVp8w6XfTTqWV
8KD3iECG2/NLB0PC9fvDQeQWTwAe8pxuPHm6xC/eUomu4LnRaeOOZKIndkXXWt+3
wUpR9pmIxN7pgu+YmzvMpF7zigG5e3/O5413Vk2Qn+DRHjZ9mqA24liZLu4w5u/s
7myjmt9Sry1xBQupNGwjGZE0PBXmoOyo5r3XV7T8xq653mix4LXaG+UrXjDgeRbx
ECXve9vMrIfJXCcnT3dtgcEwMeMR1+K3O2F3YvmvHgZN1RLUWR4sZRuPaT5uFbZ4
amVM2I9+HuuYTSVp8DoqnG8lyqnLu5ciQot5Vl1zv1CKXm5+S5gfqUdcHxiXMG4n
CC5LrvMr0fQkn9GvK0HLrUDl2QQxecxcMCzsctwHL+IBXoA4UkVzDXt8uxmghluA
HDmKe4FT7ISwco2pOpFfhSo5h1dxqYZtgavBJ/IspICrOZK4LnSi3ePCfAPYcejL
wGHkEY936X38WPrITOU1i2Sn0syuns9GpPiF5FUoD46XAPpPGfYcPdbRyntUxiyx
UjZ8KK9lrRXgEy0ujKTFtiDwLKARq3P9+UtyoBi7lFyOnjZRQYtbaCeZg5oXq4ct
UHlsDNVZqbnBeSQgeh/UtY4sSw2ALSR5u99HWqrdAHGA7ka3WWtQXEpfFJTbdVCD
sXZFdWydjaiPLme/imZB6venJWw6wHX+GjOk7IxOA0Rsvym7N/5KMZ3r1HE9NB47
4sjhZScOggRz0VPdIbjmRKZxhafNH94+Wo1zdr0iVi0Js444j+iSWwAdbcAKCugY
G8sK5hS1ef2iU/YeYDFha574UrxOnHgPn/H3ZmkTKKZRHpx34oijrEi7imT72j8l
P2x75xpc71aMPFPbAwf/mX81n+LdccZqHLr4NW6OFF7XF6nKQK61BTSsyOFPep42
6Oy6uVzF1VSxqBXSuOqPqtEV+055Ks6LYzkW3rcO1jHRXhplVl/nNzBTIsdvsyzT
Cb8ZR7eY0Zs3OaPlzublrIHVJyw9aFkj1rnKGVpMVUs9dqMYgEN624u3dIkKkt5M
HOOXYT8QTKAO52X0pWfKPufxqxZDzIDNPZzvJiobybUFEQvX+ZuT809SSZp2Ff9T
HWj7WoYmU0UgHGNhzXbnII9fE2y2BMGXUGHCoKZPPx/reeiwlFt4k8BV6D6K639u
WugjsLqslhTXJmBZRUC7IztlTZcWWm91hnQGjFj2q3bnYzTolJb14TUJs6Lus7qi
CzzuU2azJXXP+eXxP8e+6ZY1mwdffr4WBpiizTE1rmk+C+RqTaEcBnAFI3m3qXmo
7X6uEV9wADjGyvG//63Pl6pR7WfPo+cjPtt1xmPmpQVjykmOJYHk9yBRy6n83pX1
t4fN7I2afewP/IvgmB1hsw7huO5QlB1Q1tZpd5C5+mexwIaJHMafMxZ+MAmfcj07
h+OdsHu4K0IhUdmfsf+ZmGV/DQJn+Tt0sgNnY5iAH6soJ+S2hAfdcRQw7nZgWk2z
hzFEjkOiTOD01zuOnkIWw8/0nSlmLo9Vl12Rw2gQdlLEwpTitqjWdtYr+VW9Kt80
GiuVVmj8cGby1DZ8eSy2Ad5n1Is33S1RREXfvDwqnbr7TiAfvfyAzZbPX9SKgMjj
vVqGGyVfAW1GI+qVSq2383lWWpagB/JDHNG9A/MkK73BtbeCZFCsJHdgBTOswSmS
ATnHthfgqwrV+fDmH7f7rg7eS7XRTpGoVePH+p5CZal7iSDSsyOUUSdcsFVyijCm
zaT5CHHuw7M+Xb/zh6N3GPm4z/BaXbarltH9uElMqLTN419rGlYMN8ZHAs8jWAsE
9xBp5p6YpJkQnNUM5LGXNeoHUX/iM5xSgP8A2efSJlCZxOntxO6uJ2zQNVwo/xIz
QFl9DwZ/gnnuIGVlQemdP6pkC/kE5X2MoEGQJuxuMsuSo5nPowJZine2A4aBn43F
wkJ/VvaRVF3DCA6X6tTDLsYcvAvhrcrYsR98hNL+f9x9iGJEw44KFqe3gqb+W2dH
+r/eJY1rOuXZQu3QXaqUUKiPomowTsShdwecwwTf6dyh4fRl5MvcvxzYEuyGiGKt
ndyYvcpDIuPbve3EzJGvXEhRm7sV/CVVbcK9RlqlbWtlrVGA1IhB8gkGdrE1NsaU
IMEi7hz8OaEh6f8qKBnF83c7v3V4L4vRHvFBPG6mX+uRNbABwhQPvW3YDHBz9JNY
8xd33R6kDSdWS4A1F0xSYaNjxlk1rGRirAjiYWkWFsBbEj3en+k951DaDyQTa65w
hfHK6yNHqO14Yp7VZLBtPdNl9hrJ0uDVf0Q6HOaO8KPdL1JAHKO/Vpu6Z3C3xdjU
g4znCm6sZIZIaIdbmnpHRCXMCZSgRC1DbAXiNhdxWQ+bsSacS7AdkPM5t0tXWoVc
4LHbIf/9JQUPBmrpNV8vAp/6dIW6p0ZLYcqcFDHSBnr8la5v4OpiZeuKVi5SZI1c
Kcj11fs2HTDU5UB40AOKVViZtqTbUaFGbFHEF3Xy8gTJWNB7RtLAk/KVX6LJwuSF
rfjosXmO+SE9LTA62VTMEk41q1IuFSOG5a4Oryb9m9r+af47aTuvhR0Den2QJY/C
T94FljPnmd5CkuDwiVPO7Oc+HfYKx4HNIdolnZDrFGGSrIw7/fR4sfHz++jCEB9q
B/AGPBSFj8igrQJGR4L+ircMjxA8rD61v3oQbbZqqiSwB+jeX/E+U6g59ed7FUMW
iqV4MLOul8wYuCJXM09+2xUGlgM4vbn+QYj1XU9P5OcVczJn/ZmHc0PhnYg7KpfQ
9iRMSpgiNx1m6FFvoa/sX7tI9H8HwSTTG/3Wh+2JIfeMf2IXnZ8m9W9NrFfI14hB
jFi5/XHIhREnM1WScN4UiQ6DQ4WinWd+IUmdlhIRyMuV1raHWCcDbDF9VQngngqF
dzpIl4ynMfirGCOr5KPe1weMRfTBDaQhxEy7UuNGE2veJbKEnmSUO2NeCofs1i97
S0YiGht8mvQPLPT5aTpvLz2ubF9g81OgDk0CuqdRBnYxe5xTlQS8TsLLrcUkCNa+
abGWlwy1ab3aii9ZHwKTwXmET3OxbRNAcXOm1+Pu8kq3QuZBtsqXkqztNQzanfC3
7kyROJnjeqrfanEZdLPsEFasBdCYducqthF4vdQ6B5F+fuODuPqDPhY18dkERsXL
ovdYJJ4BPD7KFRGsYjtayik9kfK5H7XeYCwOvm9dHuAkcN5OtLLY5M3qUz9lpNt0
utL0MQhI7apD4Oc6GMeNDvgKUKf+H2wNhQOHDqYeH1KJP2pTuT9WMc9tEs6OVmZ+
fcGjdIy6/c3vUFWhY0C3F2t49N/ibSCanGOlSsaHBFWe17YifBFl2+s90FWxEdcP
FcSqaSGtIo0kbvlBR8gdDksknlbqwKzWPR+LRV0HXPH53aS0AN7Vqw7PJ3v9LMTw
YJG4Mj5SsWNONULxjL4IgQwIG3+KrQ51+5Ot13zQYJwh+vWU9NMz+JQH6mEMm+DB
rUIL0y020dtYAT10+i5z6XU+lG1Zrmqw2CWzKCHr6Cqsthx7JWBEKpknk4ib0d1/
IF+8UAzn48AUJiA91E3I9CKATYKUlLKwYdlomGbhebjR+CRR/2tK08FCAUeIxMh+
wfIRGdPxhdQsm24UNtHGw6SMaSbHBZYatNfArG6BH+VdG+QaChcgEtwD4uBmkeJV
FpMq1uICR+1gyhIJKJJD9gJVZVvIS/a217KNcpsqZs10/yWE59R+HilKYA9AELZs
u9zqO8TUGppE6w56b87jQRMTI5zVyUZRPhBMjRcgYf/nBPc0IrXQyRb5tR905FKA
pZEubpML0Q/nMfcojxn+THx5aKxV4hbAfp0bqN+0F1ACKksFLLRdWy5CGSpmPeAl
E/xIiSk3ZZtG3mebGeVeN6Xtv60MpvsiGJk3H1+j9rVAvLlMEQbFCTXOMlxZJGck
lIkmKXaCB6kUjta+EqUQK/6kl8T1kAoOLUltVSdaXKQfb9Xh4pi7UjmbRtH8GXXx
9BS1duWUgDO92AKGZN+pTZW/S+K0+YN0af3H38c2wivvqy5kduwBq05hF3MB2Ftc
HoF9ToIaKLr1onqTwI0nqzjertZ+S5qlR5sp5HeYjSJYmiRi0KmgcJomO0rAeDoM
Ne5JLUs9O0ZQB+So73sRZ638+A+PFOTDzQM7aoEX3lYUVBoSzwfoRvSr8aEAwQZ9
Sl1VrwjcrRvzKeX1kPvXWfhFVXGmQhekf7mTsnMcVUItUcepHYYOaKSGZzXDKYHg
wYsDtbnM413mVNeJrZpl+30z8l82+fcm9fj6ktuKGjJVKw0KOfpqHTcAwePzDMcU
IlH9YxaPvOGRxXBM+EVpeX5S9TV+wz2abDLOq+oQz4saOgCGlbGDEqWrBETVvi5f
sFiwVCkHEkHBfIQIiCQJapeN0yfjBkz6LWFQ96EoSsy+sN4gDKNeV9AW/FApDUcw
06msK65KjP4CV2LQpBy8FG/tsXoPXaIOAdCC8yXNxkn7rsXr83V6L0CIp1OpQGJ2
BDqhTtXPPprSfk1ej9+Afl2YRKfqhl0EyCheSI7PBh4sUi51RnRam+9I1w3/5uSg
KzibOHTVXej1cKpdguJGFBXMxmuBFcbJpR764hInlzt51olImTNtjTn9ZG3xMYzH
tSfOic660c674z2OWseu5BI0Du6FUCdo/YXcExQNb17UpBm8T0FQMx7gKDLxCUVi
VpMFYedERADGmspUsWlRnnLPNuGWx5uRfCaAg53VtjxZuVJkI41SodTu2EdgJiNJ
MaMrcLSmC0KlXkoXlYCH1ra7aLTRbHtQMFmeB2NtfGtGWBHGHYaaHxzz1Ljm7VnG
l2qTo1zocJFXz37ffBFVc/Al9tZSauFCwQgB7tcZoD29kp8aRM6Z7wbvJkT7b3Fv
3Qkh5tLCR0cVrsO5E7j5p0/+SLKfzEFxnD+dcckh6TbXuXhhtcCWQRgyIniz1+iL
Pc67hH2AnpgGop/JfsLq7bT0/Hvct8MZr2bMo/Xqb2RQtB8Qf/lszZRDbkCBCY/T
CLBS64wRuRUH324uhO5h/JC/tl64vrAkh8mtHrCqI75unzSxJWVZ0Lmuynl36+q/
qbRb0OY1e7Opyq3udjHAPW/Hkr3NQCbhw/Ebvbyv6WO8ULY3szI/tCcMagFDAzSP
UKMw8jrttSvahGxVZrFSSW49QD2tgRLZb82pLr3z5dZLAcvav05XHag5GvlmbHeL
i6vz0yzwFGW+4WIWzf6Cz+1mF/ortevBhFPhOmVpI0tu8ogqPGqJmfnvSgbVrciR
DOvQsD7yH+YlIqta+FdQPP4dNhobYNxd85YF4z6Gnh6YNqxegJ4cSCNC3Dwtwtgb
EqfTzHrBPSXskVlAmmz/+XEamKYzLGhQ+nBP+gmLHhfDMiE2s+IbNC2ABYanVW44
grZQhIg5/6hnw5Ln0C/iRNTmOpHFrBE2XhBfqOUMwZYXahA7u74kVV6iczGhp3Pt
431VVNy3G7TS0bPykT2x2+plG8LCF3V/g7YNmJ0H73kiKuyex47Mh7OND4xvqpyM
XoeSVkhOD1kBsyT/tWz67CyzulNpvh8alKiKTmnAUQYpN5uOsVqnHIpkDr3pF6zZ
o2QOypzRZtfnEVJozjT1N0MzkvFmjR4rL08xDHWX3Dh+t/hO7EGJzqk5s+msfAyL
YEblNK8x+/M2Xc0N87SvD3cBNV0FlSFIA19ukzyI1zAXdCiu1JvZGWKH1o8UdU6t
/G4pVnFpEWcM1VyPug9VS1zX1Xgyfm9RWcsAkFeLWPHvUZHFb1ElfQIolT7yEzGr
WYP9rRY/lAiB//TglDOagmkKJ4wLRZ3pCbnbriwTGwRWufts2HqwJSqG11ydFaFd
Z3rpQaYf0JJry/NP6rgtYCtGGnRnbhoYwK+i82C+YMCfczRB0I3QOBw9OQ/8Gq0R
T0HBzItKvBFLDDLEyl+JwzNoXNXpbNaZgjPctamlltSFktulZwONO6zlNr0Dxzaq
EjOG0//e3izCduraZnWUgPHp9WTba3FkalFO5lQi8MxEJmoCxQaoGrwCnf6a/im+
zxPIFIYdgC7EjLdqGJedCt0u3soWsAaaHb7DSiOaY85DMVW5UzfY+BgnIjj0Ksbw
A3Cf2uptQ5VjrDqxZARL/QPdsUFLgRExnkwPzxugJGrpsKw5GeV22FDztfbc02Lv
1TVa6mEUInH77E8VVBnpTYAXpfSOCWX46JyAYminn6RL9ojcDK5zPqvJabcI0lv8
DOUJl17KYDX+5Fa/YMZXXyJiZcVhDAfsu6v8IZgGFcySgSo55zmN3CND21HfNSa1
DsOyRPyUc+qW92YqGALPahlA7dbIG4KKpHh5ns/pmKKuQXkMvo2Clqu4UfyxfzhN
ze8YCF6TTTw4G3wMjH31QUjn8kDSxDjTH20c0NFf8FsihrGP5fTtee7ZSQ/fqu7v
8ctwfFtLTNbgHz2ux/uTQ5+KBJATWWu4t7bhsRHWH3hTcyyULgSd6tnZC0Sviokr
wAtSqRuciA18j9bND3J/oyNFktGPA31RdpuDpXcpI7pHJQFdlsgL6peNYoAoJgKO
wKCDJRDc4fzxLh1XxuJ60H50yrwcAkRbzA2jyDIxsayJneuiDLUc7jPBdpWu2TNE
t8DFeIZFkMWPXLVJKk+A27YOQadvnxt3dnjEtiE/DoJb67HY68qWu6L/OVjFjw/s
ZOGU/HwQoadbn2F7ZlNESySQ4DIS88Tyru3kH/SlIQGq2n+FVzWZJ4hxUrQQTp4M
vXTC+gkF8w6BCje0yCYtciY4qcBRpFT7oCsEIAW+0NexLFUVOGI3BSuRBu73htX4
d45U6CN9PL9l04werh9nmxq8MllhevJdujeJMjlA7n0LGAuRzkZ4EZlTeR4y5h81
y28H2QGFO7SmN/Vj8GikIxWcL0Z6fHoyCOjYz98Q6j08c7NUZY5NdVvax7IbQvpp
hx/CEcviTAX/MTlsKBn9tBbvFY6tK+NFNPku20fOUQOP+1NlUkJmvXI/Pf7gtadj
L8kbTYd7J5KvEwQ/8+DUHpgcKXM/SxjT/kVQ4C1tm10zHW3hQx3HoOw1YlUFZ9N3
IIdalql2yBjOTfrHUdY8iOYl35Odrna/vGz5qWhW1Q4s7mX6vNJqzdOoj9edS17c
UcJvLlloTQbz1GczkF2oNmsofUkjQU69KyYPekxG2vReOOiz1m3PlMsZ8aUMMDdC
yxcfPWBpYUImTQA1+47MAPD155XguJqBU+kKdNvGuAGhNVdTC+pCBAq7EUUXhmXt
GJLsEFw9yCdSF8P8dCA45Ve/cHxALStFrfX2wdQUHCi5BVRIZiYljn+l60IZQGHx
mbacxJq4lCm4geVd6+Xk4WC4m0C2SUACIIyZpa3QCyt3564HD5xKq0C7mUPv5Aeo
ErQZhEtgZw8w2Yxna0lXFOhQesRAMvgIPTVDyQBYjDBLu9yZ7JzjtF4taT/+NDfP
GP031jLfxYHnBPDqXBfNQNEcLr//7gatIS6uZoxcaXbMvAY7gJMnLzQF/5qFwnE3
iVuAlp12jRU2ICZo6patvQoW8CZivDxxrlL4DxIrRTkv/RTPCihqBM6GjNR58KPr
nFm1VTeqXqRphV1isEn3gX1Ln9I1Fy6IJeaCOkhj+DInhqZFOLJdLMuCWZ8XuOZn
2Cv2vqZhyhG1NKknSNcqwBkLGgdxrVuqECOdNcRJzbowKtAvqH8o2ztPyGQETj5N
nNH4LPPkRSpROFMUBroyRwhvmCdI2voTIhbjh7+y9u9RZMPyPI9z0AbB1ykeIqJW
zLglyYX0qXWOUFzu81AtdKLm4QLkdsvmik6C/l2dqdpnvnmuERom3601/ftko6Qj
jWtx1hJRFIBC8ffDT28YMCyx7puzJkjOvJHfSVf/d7YRjLBzfhPVR7kSenivLCmL
Zdy3968T4A/x/UJClF60ubDEwfa+4Kg7msap8++KG+HoyfzSnDeOqm5wHbL7wOqB
KXPcSzwRHbX/l82ZbaNMmX1g8rgKQI2QgUUsfzWuGk9Elq4WRWuBDnREZ7AleZOl
vwLcFZPiXhbdUpsnGXXC3wwnPkTuHBPBNZCEjIKMap1mWr4RrJFtScYuwppIBdCm
C40trBIVGYhcuAgZly+yU0dwYHLKUv+hXtFlOukNCbKi4w1OezF139k2EtHxe33A
WhnkAeIBmQXDuiIvh2TU3UU5nqntor9CFd2n2Ouo4tUnT46P6EbmYsPrL3o1tDDY
KvKvc9queB6xxeEZpx1+n4aMT+oPwhqOqK+AeYWvgmxwW5PvbI0+y5I1zSd4CPSv
HyybMHPoNqTQhRm59GS9WKc52wENxb9KabuGmVkdCgMh6wOrje+6GaB2dITz4xBs
68LHqXio/XGFqe1RpS2QvvKyVpiakAgmONR0vJyoUeUNBY1l+cF6/q6K+DsV4eyW
2Z/1XAB27nYto2PyQwN6yM3/iQnnwf9mwbBCwmXeTKTI6CPG9MXgdwWrYyoWCC01
ahhciE2B1m+DsmtdKIAwyDXys+K9iNnUCoCaIwcpyEsRyqi2eOYc2+Kvwa/V9EqK
g3fuhedvBRFRbLBlHA17nyLUcJvGlN2ZbWV63g3moCKCpXDtORf5tUrA9XmLnhLZ
ydefXPCzw3rofUYH95PgUISQbvXt/PZCcmuYA+D8dRBwEmdaHNR33Y1fGo4sjZ7R
VLyqkrbOB7FQyIpzjXiTN3zchWIM31RhkMfVhg67gdY47SmyeE4nwMv9Y0/4qmhb
JtHXxOnlQWcj5LXpzH7Bv5ijSVnNKZZgS2PQFPkm5401IMvwHxwsp9cPSpBcIrLE
iruqHe5e88mx6wUy/hvX/lR4uCRYGyEqQuv7sEjNgYL1+l3jeHn16BQAnaAp9ax4
g5W+zF+vr/KHyAtVtk7ujMO9/zcnqbRKixeORHsQO4pO3fhUNYe/C19swSi9DMCG
gBAdYyGTM6Y6bPV2RYbGW9SLzuqsM5xb2YgE5D6nuqga8R/xWhPJx4GI9kP+N7AH
5hy0fUGCl86dLdFuQyHXaX7tLXOu8nkoumNZ5fQ7HKpdTnIHiZWxkcrMzC3aNp5/
aCAw8ZCw2IdpKuLs+VF8kQVyjjJWsTcs8KWfHKuwpIn4IUYeE/+EeaNHliAGAaTg
SSy9Fdk2xrS+WO6XunqSeUyICbixypA5Sl5c4uJFzl2nz0Im0UdGRj5jBrxe+oZE
5/JFhTQaHrRRQv+dGpnmG8ueAMO91dPSkM5ckSVrkmM2M5aZgTJqjEVT71u5MKeS
UXNw3+KetxqVXMEFgrTbF2523XFA2vY1TrLgTSVIfOOVsHxaD1SySZUYweeOJhbK
SUraSHEDDkR9yaqubVg5KjSg1mV5ADUFzbI4uVfadUyX/dghwaXl6O5GrZhQGHe8
meVCxyL4Y9bjxo1S4pKAAJ6DUF0nUMBIyLqD+W+SVhw/7+CzN1THShIhj2mpN6qn
F+ge0UMckggGTF1aM+BPIE91/4LUicSC8AEqrATvlTnvBptCfJWwqQR2hzs/qVzc
HcNMlBb30LzmNhPRl/EktGbXF3XDTH4I5L021hkF2C9IhKZWdWB2pUXjtJeVAvBZ
4d/Utki2Ex0FlWi7kMnIYirBeB6Z0ye1wGRtsIoHSjnsdPGyAMNbrcl91junUG3u
XPG/lp3xCB30q4lDKaoHDt/Q/dS4ULQrySE3GL7upYtZQgEEqzombaXNus1m5sRY
jtK4Hfqxcd14ChX0Obg+7SDqp5M8HzqHYmjVD+VG/fevV3VEYVpn3inaH6a8o9ES
+NAXFAXl4W2Es/w/Xd44aH+Y04y9Lb59ggwCwAh1Q+zHZnOHqbUjy33HkPZWIGy/
WentxU1sP8Pcd3/C9noVJIqngXPH6oAP4BLHMKXCMXub5UzQrZk+XXmXGxKHRM26
Mm9mJhg2YoW4/T36CYXQfjhcUhXGB+M1EoKFpI9dun14REC+XYGbwsoRd+6hdEud
r+qjvBx7uRXSx3QBHPZf+RaP5dniIl+AzFiHN7QCLr929MA7/YQOU3tkwZDguiXu
bZHv8gn4P2G4pbbtVHXpTCTw9Rrqp1OJy2B1qpQJzVOmlE/HY/K6VXsyaFWoUWtn
cCHsNxOu6mLb2mCyPCbqqSz5N5pd0Q6+Z8mqYCgq8Jn3p4kcGC2zyUxSzmkWyCS5
jM2bg/zfY/zQ81VVWcSfufUSrNyFwEmkvT55f8PtpNEHTRt3GDxdtYrp/x3vJFCK
ktMQAPjqei6Lu2Hox1Z7dkHzH1cRUFJiLy3gbv93nItA+YuHOcvtuvelqj0tGjSw
cbAViDeUOCRHQy/Ca6lYe1xVnmPjLtJzDrGvvBW/Wvh3eGRC2tkII8ZzxOlZ424I
jveUB5VytOwM7J8+xdFYfbUuH0OJop/0+GFYXq3ljNjRQpzTRKGTjZr7uXZj222M
oTZOGN97hwKodB1znXwWO0IE9MKj9uibg9GpGgt4niTXCjYJQDpf/BAn1AB9JCYz
QWuDpHX436YNeryhflP5GkER5sZSe5wMKYFVPknbNeUsKpzqVdUGjtjRLHtgt7Gx
cwGrN6xtTrhp9OgvWp/9VoU9Stj2TdV3XQCBT2G7gSPaGj1ICcUzFosJK8YjzdI8
qCYwAohRdEIyq0Y7VP6J/2pbOCbWylrGLGfBORmdC18t3NZKXXAxUrBHU6hJui9z
+AVThv82so0fxEm1SfPaVFCFA5Ub6vjP6nguJMjsATdqHleiyJSm1Cocr7zlEju6
A+LsJEjWIhcYS+nKSxGCOxezRFtZRTZtt7xiA0+gfwrdeYyo10EsClEi9Ke20/Zw
HyCpxS60784wSjm+FksFtDnPE1xYy/MKAt9PBeCfZwDVlYbgKmdHsQgoC3ZowMhd
a4M0He5sHMALZkzzE4/Ir11eFvezr8AYAE0w7xpxHM+B1K4F/lKfOo/lC9JKpJ7+
i0kpXI6zCji2iWHVFzqHiXVxFJRArzZwBmLV0JLjHOZntzcHCmDiVaNQrZYvTGUU
i/gdssYH8Yl1wZFA193U5KEz2FJHUiFerYUd9yZcnap8+tGtVXbWuyBVArpUufbv
OCryEbso6MZgwZv8grrt4xul5NNI0O8dGfZqfGPRjYuY0LjVF+xQ2ot63KEiD7TS
ZmBCE8R/RFThYWXBSqnaVPMA6uuQG1JL3o/j7bjAvvTWSLmyHADptroQQ1EGRmRm
UaOPKZoqqX1wgoxcvibcwVUrtZqfW+HuwHxyOi7bNSNwElNG1r1hsQ/0ipNQDY6X
BcaPtGwjoRoVv3kBRWw+FYWIsmuLRcpR9rmQtYe2ml5eHyxdHQpUoDgU/nctP2Dy
BCeK/zxhQ371pgn27tShismm4ogWzbA775ka4BC6AWT+5FHH35UOJWASCCZw9eph
+OLiZN2MkPBx116aSMhz5FAK/6278JOwUFo4aya4MHwUQb5Jq/aQjts9YG9RAsav
Lz7sEevHgsc/pRiY6rVCFQLrIDxVSRv0P+3xY2CL5TrR0JmECnWr3t8cHxWMjg06
Sftaic52SIp74uZXj57sQqm+lJ3QTaSqVwxJuTX7ynOMUVF0wpdjilruhV7gKifw
auJdyF8qC5eyOy+j+RiqMtv2RYvQB/LnM0516sYFrtFg0mro2zkhvc9zTZQ1iJRn
4MT7oKxotSk1l09m+tUGgicqrr+cfJjfhHDcHO34AmZVQ8BQz6IxjpXVNiRGWav6
MPo7hPJw+UnwSfPio3oeOtaNlKb8YuZy6WVe42WkdWeqD0HboAkYqqcc1gFz/H++
q0NM+20CoLVZGr/Kn3RomQyZ2rwWoI/meuo+xsh4AvKDqJuaLdeM3rG/n/9N6Kvd
rYSAd3/yeQ1LWF22fqR0JS1ULE9O+wyIDTaTmiY/k1aY2vjmtTaWDQPjXEFmY4fW
T3tgczp5uUb/ONFfWEbDqO8Zw9Xi0jOn10cVqulUND4pNsya2iUmfNLG6hNa25ib
bQND4Gds4MAuAazj9aQdcg63UfLInjsg0mIBg4uILrEbi68i6cvHQmbRVjsvynrl
7zyeO7kkNc/BQLOyQWkEzmPqD343/yupEhpzyrPbGfmiQAbOkmK7QG55jc4cQKUe
EWsrc5nN/vHE/Yqr5+uSo/vxk46GuKoKK1NJeNx/iNmWbUglQdRZYOw16z1zpPoU
aeQJvl+EamDat7ZuqiAocze3UPVCOaWQfyuegSO0v94GDmWxOcV0/Ho3Bojp9LoD
RS3FCcSaGCQMyZqxC2IHxMbdA6lBOIgv7JpEk4V0srJNb7Q+DA60FTDPXo/CS09i
b2nKu6V1psoVbbhxahuCHVyJVpNyVW79yctX4ncA4BWwdw0DV5BkSevfujiJIh+U
NwngVUuW4TqxNDhx2Vtb9aaQDjiA7bodBSexhX7uy3qSPiIy94/eRPO7X0SbCBtx
vw5QGqAHYTpYWvCTdBOx3eUFhLaKyW/5wwwnMLpVrsM4ZGhN2c/1NwBqqII2ZNrL
KUr0X7rfph2pEy998WPLg1BsBsI1e1uRLWyYixqFZyJR+0ud31oUsaU5D6GMO66o
AdMUWIHVUM2ji4VR8a7iBfrG2sGOZxpQqO4ewaKcseWHnlaZxfm7yw8eE3WM8kB5
tZVkUgSIxazRII7CgAsxbKKQqGNthogiGtAEtMsETCGLXCFQqvV5KgzG2XtgZDeS
cPAosHsHN1QQRCLVuy+USfRY1ZZfAIovTcaJm6n220IARyyEt9QoKIvlE62O9nr5
Ueo+mjGZCkv7Ovw5ltMNUQGJUnFgGBbz6MvF5xSoofUgz7QBD57l6N37kFbvlpcr
Dg2ptcpqGsHoaikp3FTydT+szNsyZqgCz0LKFhzgxOv2GL3Ld+A57Bx2zv+yqr9s
j2flat1gcg9cTT8M8ndXmiaRUl7OvzWVt/Y7PVkB9NL73ZmEeJJQ7PmS2W6gLGLw
bvygdCGCPmXPXCpYgJo7ht9nAqyIacLLTKaQ8bGllyeLbmAswTXsEWidOXZ3IjPN
MeJvaaneGFvQpVwYlC86LFkRNfP/QiRgdZD9Eyhs0YdOLSTEw0DmkjK+wQGyBq4v
s0AXlv3XO8xJEc9I+hX22HFVdipcGdFBio+r9yMOPEIKskAKL0uDb+4KKvO5ZGds
4Ep3/EfGRWSLFX1GoXWL2z35h76pP4gVXKPc72YBUmxje7CI4k3Pkrqa4koAnB2C
YO2eTUV8RTB6UuKxWMEZDNGL6fqY/FcXz14lbd58k0lEn3BUNFki2YDVx2u10fKL
/fj2OWaalHgKRmTySg2P/FjkzcyRfbVSd7p0qAAmCp0uYtuL20toAApoB81NY2jZ
wRT8Hwq9xwX1fHbushyp6jurT1UQcaYBqs6vZeqUWoAAXwGz8mM6i1okEwuth0la
YZXmOPBDUsYE2/brjwJYjDMVNMuGvRDGB0uBSiqPboSi8JcypgYnuSl3o9oNlFkm
9sQfygq1G//E0kGNyTmM95vFrRdvSSkvkPZCENb2dD27FjIfvfwugAtm9rp0mJAI
ITl3HnA6xjNncbxsT64hCAw6KztaeAIQ75W9lKcJH8cKxyPmQOgrb12SyOrJb0F9
8zvph3zJpiWDwBOBOeTq53jWGoFKy74Z7pF2grt9ifvUId9Gt5tiFKZsHMhf+2jd
eB5GFGTdbkkFC+BbuPKeddtpFpinelLf515HI3373wkei/JY5NGdPRdMAlYOLFur
nEI/T9TSVpPsV63glawq6ZZnynplckfbbDvo4B7S4H3alQ7sLk9ib0oKlakJy5dI
/gTu3BdDHaFg1ADkOeJLeHQjdaBQRfv4umAytY7MuJmqvI/8/E/nPpHpg4hw3aID
yeTj143rxUVesEkmUyL2dxLNIvQdhSWxBlnRWocr4RtZfn34YFhzbbcsJGXABa7v
yjm4KX95mVkNGWc7vM5bybfpUnYbP9SJKsU+y4D4INFoiqbKGSFr2MM4+/QCNuUa
Wt6E9da9x6lwqYVzLI73GM4pcqUuM8NAHQDS5o074GaS8j9YaX01j6vMAeVxrnDm
xL9gAdtOuk+gwqatgWUYVw59wsPi2X35gm6PF0A3oGjavOhtQjOOJEvhGB5n46eR
E69f1sMGEjfaVvGlBbaljfum+q/uc0qB6LLXBjPlhC+Ka+9rMdsfSlemybpM1NCS
bLvMP7yf4nodnED2zcnLLbVpd1nnsB8Sdj7P6b71Ciiive6yaIs19f2yJVlcd6Qn
swK0KbBbU8hXhZJBQoJ4vmql+2N/GQt60mqUwpzvstdiBlc9OGU+KLw+mlNSw8JM
Rw34mDCfpAyy7fyfseyCEO3IXugtzJbTpOu+0wYEd2+sslx1Tl3yQSvzwMzOuPJ0
QVR7GF4p/qT5UYtI1ZSvfYwyy0Hxk9S0VWM1z0qT6f2raDXjntGphxIJKK9DuqGz
rO3AqvS5+96vRlQlkwJ1beosp5CSbxcD9k0siafATWbiqqkYvYci7OtY/cGyXZFq
aV/LtGy2tRnvgIyXAFdvEfAJgHk/NiHz6fJtU6JMrsvcVgJPpEDofgJ3hkTF3qV8
W04WCkAUGIwhxbX+euBlYNTxdGs59WWNYiQtitBT4zlg+MFAge2rwRKlhUNSVJ7T
Q7nRM8uChycgYeveP3suYcarP72qpEhFOLQJmzo8xw0Vdtd8vmrl6hyeGPcrbJPR
t0mFL5byGiwRUTr+3BCDqKPlKOLi8wRwyKk6ktLjwk5TYIhD8TKcufpjmcT+YtfA
xXHOyag4vHUXaLsyug6oMH1B56mfBS0hFis3ZH8c3wDyffYU2z+KSRUBpKbVglUz
S7yLfjUhSfm6uN8q6mYCdwCuISDw1pNxa6+4zAM3jYXr3PnJ4JhR1VODiTTSWqcq
jYVS1Z928WtNICkyWUeXUF68toqo2q1SDPmGxZxk4QVT78gjpRxWyDQgp9asDbtt
7YtrG3IKU6W9wTT9wqhPn/Ix+hwoXV0y21/Pme07TqZcoM4Of5FfylOgMaau/ZKv
jvSgbaMNKCtfFiRP1QfKXKbS44bAUt1mLfziYeU+opdVAdNWnPrMvDYGfuqDv+st
UnV8j6jZh5IV/ByCtjioCrT7uae801rnUipOeVBusATqRZVPVteM09aUAan0GOdd
0ZXDzWX4iQaqSq+w2bGti+CB5K22EOHA71Sq6ntI+1I2ySxosnVcVGpzWlOKld3j
MA/ndcFm+DXbVxYrEtEqS9M7//OJtb+M3Nt+ohKbKoWzQrf/W6NT9HVXT4tSW84N
/S9GDmimS8fv0v8otzVNSLlRTS6NUPXnfIQZaa1ceRRRyGtWVGqGKmVylf9T2BF8
PY9eBEIv1UUUefjykC2hMBk7MCAluNf/GZjAyDP31Kk71GVa7YwCj+FsHNyezZd5
Nkg8NEajF6p2TqzYynMjwV3FhfTz2pxvTdsSARDcACQACTXTj2KEHNMlwbNZebcu
sh2g/y6lnpIN7JmFFtuUdgvtGsdzDGR7JOED2syWcePY94JtSj+TlKISQwZ0VoGZ
L/60EAc2xniquqE/tPHOmyxDGBYiIrqMqDt0vOdBeUQZMvKpL90/PSTs6ZyPIgk1
NxogcMDgxvIYqqI+HgzGapZUwtO/yrhOXYzfYhhhrYeMbAPYfP1p93v6jzniik2z
9ev3DLbaH6dtBjT1xNHzi6IeEOubGQBKRtXFm0YWyx3aLpkwWpgZ6p5LI98rmOxx
ZXVUhxmLdC8a7CVpa8NgR9NOIvQLTHlsUhBQjs0a0fvWcrCyvUooNa7lhU6p/rux
8WmGXfurZiY3IT/Sr9A0CdQfixpLpAsAAdnCPi1PNEsCJno6u0Y4X7kZ6LujIbvc
b+iIi8fPOk7fqAmDLzJZVLLwNc9dIPIDdC+bi2GKwG/wMkttwSyRZj6ev9uSeAyF
xQPYK3146VxH0K2jGVwmuuHKSnkZEDPoCGt/kLf8fJuhA9viigx04786tzjeCPBo
en6C5ZOPCWxMdNSGm9ncguaagHpj0fmWO/gyoK7nHHUlmnSHzviV7RIlcdtJi1LX
1ReQE45/G2bP3f2OJsKfZT1Sa+Aetc5rY60Y6lQB+CJT1G08UIJKMOqXbr35t+s3
IBtlYSryW33R6KqdAnYBKnAvonVuDvRPIZRA7xmmg3Rk+z3QVp1qjaRiR0vRwGHl
eaqKknjx1McBqOH0qkcIVuFwVMueEbP14CtYX14KozrKZTxvvpWcDhx/D9mFQ3Wh
f4L8A7w8U4jS0M0NUovkAOhRVc/GxUggvwUhnqwHZ8CUNOcdqqT6Wdz9FLP1Hv3U
F7ItlH9qegpbrIKv2EFyfCAlWubyaNnklUe5TdOJpzrwzN3o+ISuyJ+wXjwFXs6f
mvgjnbWBQGUah/S3PZtRSDz4sL0ZQvvkDMryWNa6DmixDJaXnXi6ArpEepGIZq/o
iKPKE5/iAiTO/SgqyXFoDALavraSMGIGh7KdzCxUFLQd1TY9uryLyhWI4AweJVE4
1iNLcPMQ8T6U5GdjbspR/PZ9tTJlvGuzLZ5WgLxVYcC6hzLMBEs19H/zDMS3kyyz
PUx/WiwgxfZA8/LwSgvcwxdyTfWuz6erZMTwrfH6yZkOxIEPf7n9ZgpOvEP5Yarv
8bj+hEAQamW2jCJl4299ZJoMwYVVNYQ2IqNu7P5sQJb/Jp9iJOd3qZ/4rMPGs3Mv
JrsaoY8BS+QPtRa7FpTEgucdg3SelLAKXQBWw9oPSg8XtOFHSV/L7VzD8AaMq9zH
5foYiAv8btdo4BGi6ffp57ZTgQ9PgotsuUQQShX9NoNextJwwBnRHiue//d+BwyX
RCihvZa8v0BRyzDZhT4fNgm63s+2LDZz/+BcarGOUId6NSrU7QrVK8cjbIEYepFK
4O2/FLlglcAcmsQQd8WmrvHR5r8cUKfO6YLO2O1Z89nzU71Vux16F3OOsfVju8DU
GaX5wFzUDB5BZOwFPjoEeVkWqGGTovU1qUZ3c9k2lMJUvydL2fube9YJor3Gqz7i
vXt8y2792823gMUpcxv5R/P5FqqrZ/+X1+FJVB5ujT2Jk9yjf1jCKCyUP1nXtUKT
Bqs780csH9mUkv1QzAxDvXGekUD5PLwjBLLLE1eMa7euAopy000x4nNPxmITgZ5n
R71i4c/5HjGjrkLIdm8X2tErv5AecUMb+rjUOCPgFYuioPjpMocr2lAP30BxelEp
igY0GjqgmIaVlEir5BIycpU0Serfv/cFe4pe4jQ1xgOEezMqEz76gC3Tp2ZCtjzS
PK0fNuHoX1zVTkGvTEueL8R/FGiz6FDnoOdo4zTXwcoFpz/KyH72IezKf5l2ODhK
5QcIhTFGdhm1qSIdCdZz6EQIgeZKoGPV/tMyZzBKgPG0xNXRRg3TYCUWoOAvGjjH
82T8L/VQwz8uGiN63SVgWGId79WJLjPBS+J2nK7UCNuUDgUM1FjTTJ7y8iRtDW1/
bijZkH0Id6dMbkTDW92WzBRiwBMRXIMT/2fB1HDeSmnop4dw47G2b5yOEabXnjkl
jSLvb8S1nC178xJN8N0Fm4UKzFMDOLQw8rBRb7NASaNUilChpD9XgR5XuIokqqOk
0bchhl+Pn3Cq8p7aT9g0NVpZdzecSU3ts5k2sb2XxNtYvKPllYxwLjHiVM8bJVL8
IF23CVwnyCRz7LCRg+eXhBi7N8kOM6IymfsHTbvgpLcHsJ4hsqboGw07Oed7k2H/
6yEnkO/hR3UI0Z5CmnWY133PQHUVy2YBUGLc/kVBeC5LOKrMUq1A94gqoWq6+h1K
A7hFM+yr22i9b+7LdlkgATcMKeHfusifG0kvVkJOYjz5Lu6Or+zIOqTj9Epd9VUi
6BboMgiQVAKEPG89tzhx8nLAZDxITa+kYuVV1/cTlk8ErHj9PmleQy0BsZju2NUT
XaWF6AxgvHAG825hGSJEUMksmYWMusTyIT8yrRVPnjSflaBqE9ggm3YNCLKuaIzJ
iIGEuAtjQEfLXgYVZ0XbBNqWTUHd1QTWQiDsqzLqMMq9QFlUqmPRm0DOS1O0IcX1
CvLqfAMeWt6bymH7ALize3dVptQa9uA2FUSQEJ9aITwSTrDxs0GTzEVehgXGlKn/
LzUSLm6q22IHuShLBcsvfjHiI7d81oL3m+XGbnUDu/JBpJs9clySMC4kWfzmvg1S
6UcfNyxjjiuLAUt3wzXIBSwcp7flvTzEi+gGQwy8ZkOlhvfuF9PITVz252Ok/khW
cU9M525lmvhRjRHk1Xm1eY1UG/6ELxJAlRmXs+GPXerMFGP1zKnR4W72KQ6uJXwo
4mGQRkbCZ+4lDsEnHUONu4Lp4ekiJAsgAQnBZKkJXi9/Wixueu1gOyH3+HyszBj8
HjQ2G4mP+pLI6MoLAX6uVaOiEgiwehJ8oLQA2tNA1m9l5pqpnEIlfNjxnGlIxOTq
C87RhIHsAmwaIqDLgY3Js6SrjWm5Ab3AOWOp3Qqc2BlaAU8Rr9DlM4laV3fSwmgE
UBXxA3hixrCiMoNIRci5dDPcYlW04GIbJbMvIoOQebV4VPQQ8PHVLUwaHA5Mmton
6On16ybG92HOi3GdBb4KLC7hBT1ySZcilg+vb71OEg4i7i310DTosufAb1HYsELc
a2yYj3X8xFXpMKqJ99DwKI/Wv3p8da6XUMpsJLpd9wYFlte5FUylXjHMlyV3xdrE
zdFljl+8LriJdh7gE3979sMPiJdlhG4ifcjjYA1PkylykJ4+006QrZIrBvmXTdm8
Ngmh2sOAts3Jb/k24coHsbiy0zI8GO55rWJtf9gunB4zxLRz1ARJlR/TL5qFICDt
mLCFCWn6/2DArakWC5YLDrmNORWwbtPecqNRnMKuBIsgzsNq87f/h88Irep2r9Qk
BH3Qv165JvPMsNtb/1RuZQ8YGZevLN+3VSbtOLYZMqjyilr2nphKAzLt2/K/fbb7
spY/JOqMPOVTTbzKvAuubrRHoqWviEozpnYPngWQYde5nsZS+OX46RIsICgYWNCK
3El++l2Pzij+hUuu320XUxC1RvuZaMELxUdBJ5bVE9HsE6otBeuUgI1+51nDN/g0
HEX7e/d+RokabKOQyVD93dQcuvp6kCkg3YiYvrJI06mF7+TcjD3QWu+eVNKV+BCl
u+V7VTIDR01hWW1t1XlpUokj6zsJuh2XVGEFb8I0QFe7sWV5f/UTnB2+MWD2BOVR
YvA0daGzW1kQJOTxz8n1RS4EV0T8lWryqlpHuBJKGN+m5jlk6ChCbuxiE2mWDxeV
hmOfZOD2YJhWXqWvEaApK3jK7ysLg7hqskC4w9pDqDFhFsmBXXEqMrtqaoR7xRPb
NAc8gzSZLC6Y6gItG4j4udGSpgqcrVXyGmeG3yIBXQRymBkk9aDeDo3DCQpyOdmC
f4OPFy7H4PonnjpKstm+yifxzDjKSubJ271y9+Syz18Fy4Vq2CRp6ZAQx89M3sFc
qer6t+oBenmGRUCCXyfLrIQImFeltnyU8DQe3clkyogaAHmn3IImilYsoyG1zMCq
pkPa4Fk0fzh4FljoMkB/5m4x7Ht43Cirlq8fBBGrceG4wHbqiI30mvzljhYTs5m5
vBT+VwIhfyovLoTXy4YxUOFfaixuE8z/aBC+yz/a4RSk65m89kS3cPXBqkU1Lr47
3rczjNlDb7WDtfMq2ZNCaN/1YajlQwK/LFG0Ws3YPY7rvf8ArLauerCDxS4csFb6
SXLAXeFBwdQM3JDAffQDRMblSfkM8UPHbjFCaTb3oOTBhwKDruBMNOk+PBuqN/oD
ApsxqUfSh0JaO/dBE0xbkdqnHj956npOIVW4NCzFGJs4SJy5RqONfSga+Hrmu/Zc
7/Y7evIw+VlhBiJVsVwff5uMdkmLYO/Mc13/yW5DgLZ74JWNO3vZUuIa1S+nMpjn
auZD2PXzRofG1+hpVsX29I19PovAuHy/x4Fg6AjJO3O5nUAp9kYcngKa4O4uS1y+
oJpztgMEK9QAn70truv9O/Z6Lb1QPAhO//LYb1pn8vxU3OQgHergzM+DIsaT7JAV
8JOF/fFtlgPW1nA5Km69ndqhaj5EQDTMkQm8LVfUw6/BKNLWrt0BYDAbprcFLVt4
lK4ZFlU4nIjPESCK9AZ4KbE5bE0x9WhXeaO85K+U+wvds0Y1UA56+2mjM0xn1ntt
u60Mo+xmZzOBSul/2S/wWXPasMcVV3WkhKp8Zp1U6UXfx5H96z+ZzRwZpHxkK+iI
yLObibm8ZZ8EqWffogcd1VPlh0RYk50hdapcfHeRuyH5snQFL17xXMZ+IkzuwqSC
0E1U8oUJIEHJwTmxTUvaCf1K7O/YjN3CtEscHrdMWfkz8jQ/EGxc8lLqa8YHpKO1
OnrlSVvcD9bdwBF74TuKTbmOu7ze6FWLfMm3B0sykrtFpwSRKWMrZwaKR6yVPuDB
NIrtdlapyPFhfbiGR81SXroO29VzTZYXSWtX3JHTagZvSNhkohbSXscJgXkVGgXD
6/CHguqiJiA3gH0zr7HiJdM4B9ZeBrM8AgLfMwbTVPp8Nj9QDUQcvwOtvCGgrEnw
vSm/+r3hMNAVrslkhxkLdDMjTa7TM/XUDk14otMNl3P/PnaC1p7+NKkJ/+PoCVjr
IkLwC7byjT88i4debMjKtZiWwDhg66BeuFuONaBHfVIyVFGkKbNpi3V+ZvwnrNIK
8CqjW/nPw/Gd0Yl2XFn3QP9V8SwDOMUvx3+m6eh/U191N7eKG+q8e44lyfQKhDuv
aoeHR7dUsHpY+QlCzXbbJ59FO9GwBwDyn3chwxRBLZw0tCb3n8wXt0lub3aQ84FD
FPBSCh/0L7lhlzLyQWrCfT+YKVr3IF5y8VRXq77jdsOzizPKXS15olM1TbqK7G/P
niiYT7X3d14AyGL6ZbuKzFQDqZNW3AjdMKBF8Kk+vUfi9JqhlNzix0qzSiYRH34Q
OhdJejZe/JVk5quMNySOAqnJYB8fLFdK0qsZICNptUCfTZuac2iE7rLxH4o6DArz
c8bBOCKz3WlA6l/Ya5HRX2pCmd08LnQp7Vduk1/gvFASlH3mVM1cgSPfDKylNmUZ
9iFPzvTCZ0I3vwSF5dPYZy83UZeRRkpBvcPM3MHKhpquDkSmEZSdcqnbwDYqqweV
M6ZgK0kqajUBI1+xmROqMkP7ZKliE20o+JWV8bph0pO1QIyGirA6vkgc7rfRlYUy
CmWbih1OBmGRABQ8qLiOuc3PbBEXEujodfxW7nbXRwxKKyRiMGlNFoDAFOmMlOZo
+TOXOPQh0hx7//KUS5hqW152JYloBzSSVxahLQuKIwNpVoE5dJCOJHcxuwfqKBGj
/NH+fd2WYk/0uGGkKZbNoXgl0a6e3lHbtU0CcSWbXGVk6pIdu+O1AITU8/TksT3m
RJpkAY1PCqkBmM7jCVAXGPWEg6DN85zwFqNL+UjtcrmRJU54R+lqRD3SBfJcLidF
+HZgQSDgtbvj/iNQj0fC08bEM8hQJ8kxmTmLf7e4llZD7n2MiwgOWvgcUaVkH1Ve
3d7H81vTbt/Td43mONSBpw3RqXLklpFTHBGemjD6ymaS6+Keu7ITJ0Df8Ahr7RgD
vr5+foR8y757giM9BRm3nlDxFrAjRAJ88WSjfrhQYfAdDROsv51AxZ79Ku4hNTqF
udaYpqic0vGBD//Oixscg9d21z0+A5XOkQGsQ839CLVJePh6ORnFoFCmf3M7uf4O
L6xTjLsGsdN7vwDp6Xrd3ri7xNt2ubWJYxbDlKQRWjK0xotwzGIeeznuybhrOKSx
vVi27bdIM/yTiq87b6Y3BWpNkQb/0bD8qGYIdUxXxJIKVIYCayMMc1XVV8zo9sce
WnlwErjqhAiycdbtcFe+PaEdgfOeCFWCmTeNr2lyQriPKl8TnPQtzgMk2OrTD3K6
TjcyKvMrnKV46m9WcoUmujS+tvAtri9ijvEaeaxV4gYkUHpv07ThIR5mNTOCSQWY
fSiWuZmY5cHhBeDa2ydkNkUtjKxlyG5XiMEUOwnpODhkdl7myqJLql9nAZBtmu6v
breL4SuTbG1vB4KEVTplP6iVDMDJllECNVqPPsZfyR7LknQEDVYCRKSj2AQuqA6Z
WNc3rjjNRTehYFWWlfnXZ3y0aq8ceLvZdogPwMtQG184sA4EsyeySgDiNNVirxLk
A2a3RSddYzM/IL6ulq+DxSBUTxyV1dtROIomaw6PLoMhx9d1m9L40QpqKa9//oB9
jA1JHEFiRmbaE19Plx4INfVoFQKIMizQRE/Hzrb375ZSd89S3+CO92ye43pQrpfS
/CELlwvQDIx1xrNEIQgo9oTbp0mAhReBvunngwmZvbymA3u28xmkxafb1ZG6lM/v
RMHJLsQ8usCerBMtt+Ot9udoKP4faXn1EGWkGWed44VT7mTzLuqXb9Tsa3eRRNlb
/cNesAPsKBmLnEwrOa+8K/DDxZemgR+mpo1/tSdDxz48M1Hridlb/7rZZlDx2yH+
jXshmEPBPfw+t2tiJ9kshU/4ed9J7uM7agvq1jSl0WrDQ06fqxi9+DRsYKYEs6qu
+6p+TyNkakQDyYJZVONH45UbMrmXQa0Zw94uIu4CxkxQRc3g8ld/W94pgiijtMtp
FElIHyqDk1MnsOUKvXoQ0WRXcgDemsXjrBm/6cFqEQmLXCDU8B3lImhFbWlSsLzi
wq3N9mIdpXkPl26nKjczQ2ZoyjWzUrOBKK6TdBW1LHh/j3GtCCB/r0r525ED4uaF
UnncsFwRdzvxGhDUnOG8M2/QqeUKjtLm7EPGJJoHV9CS5cEDTxtDIQZBBgA3FOS8
V8eLMERiEZ0K+dVs/zMHITihDl41rOeoBWGDNDrYolp7dfakwMgkkkRTs/qLH7pY
FNC52WK99VoTLuxou24qnlHZkQGfqScoiVmzMa5JmGoFI+hPKFQxbs5uK4fHj/AW
p6GiCZnrXvqxr033xTw1U3brP6kk0Tops8WjoPdGpN4gMJioQDL5xN03P9AvroDm
C46zUCHW+lfbmClKVvlZ5Wdq0K+L5CuiwOnxOn5XwDldVCfz9EV/yLMnRDZBzl4w
GU9If9YJHvjDU2Ro6rEdtqOGBZBMbkwn+l25DCwaYUjZR9/swArEHzKlPIePvld5
NkMgySUsphrtrdBSOTy/7lNibo3xhOh5gm63WqfYv/tYadokIj1q8tsQXclF5aVH
oFyjupB3ubvMEIJPPAN7n3wf84dpl8BWbuZP+WBF+3IK7aOCi+2YuQ2hKC7vfNuZ
CMjJfQCqm31X78+KZnZkV8Nd5WnADTE2QPbphMYJp4Sa4AdVXV61EDCAWlqYIP43
SzFn97KcdIsd0v0ajTkVjtGSMH2PhoI1WAXbARowSO0SCvb9sJ/Qt35DZ3EZawFb
/ST1b3Vp8nPSpqIkE/Oe0jkdhQnro2CbztgNeCeUsZuuWbDYqhIi/dy3nrIpwRQM
77RmC1yzpn5yOZI3o3l8ca8SeAuu4rHwyts50V0h6N8UTnEoP2jNXLpDNIpYEPU6
yohEe2pyP4pK9AZ3okUf1n6jnLHj+CkKfJP1vhsmOU1Q3hOGX4QwAcizMMQPK669
V5TtSyMsoaQaQZkMQ9mb/uNZ1thDiuPKE5LvNBxnkwZAN3uFtkmWziw8v7rOUBy7
rKqRGSKePbUtgIzJk6DodVNfQu/AA48Tc0unGsd6nAf4axcnBrMdYPrlcA39IU7R
xY6tWT43Hq24fq9cBebx/nA3MdRdRtXiGy5sjc15q/1eTBxiOX1ErRzPTQZYpqnA
sfIgSoHewoEeng9oJSK0dmjH+mNmdeS2Z+FcVCLWMYB7NkA2/njWGFd3aTddluic
+cdO7nMcEIUJXpfGmXeSdVdxB4wjbeePvQzfDpi0LJXyo/Cx9Ccf7AP4bhgZg/kG
fgwsNm6a04ubCr/yYVnnHZHfu4mGqdEGAZCS0nzp4trNFHTRv4ZgUbJj3M+P3OvU
+b915hQgql8EKcRl1C79aDEd9Tl58I7atGDsNzGpwEX/GEIQbluZNWuHMaDNsQT0
bPwN5nM7ZgOeoxRu6mwi8JqxwKqCWwjuApDJDlRdzqmaR+o8zHy2HjU888mCanwg
sRBjvBBZKshXIBAhPdJVLoKBRjLUeXZYf8Y9SzuKcNI6V1Elcc0Dv7NE3nIlC/Ne
S5MwQTPvccSOBJSrGw0MlbSAv3ZBcLDrUHmjrPjCmNEWGFYdg6gYIC8oPBNZCZIC
uvPq7qyvMj0B0pmJ0QhCUKOtSsad4T+N+bj38hfdqQjYQNYIHtiibB9fm9/jRPF0
meDUpRrwer6e7NgRIp49dv/xeTpIK4KTDUL0kJ2LFLf61KM5NprzVVwN9lF7wHNM
TlQzk/vPAi7BNRnlzgJcstKnG+63EusoYyXbSRthOuZrteYjNVlOZxno8YumnCRA
R7cmrzFuRibVIc426g7j+XZNB8p/DsaTZanMqmJAOtvcWGtE4P5VIWwNxXHSYjX8
KsjZkhQ2K0Zh9NyRIx/0r8XLJxUO5Lbsd4lYqeVUT9xaNXoYVgMmraYU1O1kcrC/
+vxLm+Yd2r3CyjXIijYt7VmObDqDQrwSe3Y9T2CQgKZq3TOyW2ANNqpTlswfd40Y
hlFqquMlacY4guViFo5yveiRhpRLjxmIKz07SaAnhqtP7RZ9pl3nWvjiFxlb73nY
so/PRZ6riSDsM1VSmk1S+OhxJb45DDCQm1GYeqbUT/zP/EW2DKTzNawKex473dA8
tGB4fn0riMvwqoefhIr+XpMLvHft/G+9xj+CsB1+7sKW2UGSy4N+Cr6UUR/8qORv
bCNOs3sqw634hul9wJwy3GJFt4HS3+7Kqd1jEbAtqGATumHhgqFXSgFSlZAv+zwL
bRjXTOb8XjsrpZiENtTNgiJOdUxBz/8KFxDF+7LFnRo/PJs0XL4Jd6nGBedeLoKN
ceXu3y0+Qcz3ScKpU7K7HusVcU/JWS3OGF4ODovqNzGyNquAc0+adRYyGU5cXkBP
CZwe+pJLUWWeJ0u7s92ePBYL44jbdImdFVa+UtMSPi3FDOJm5esdkoILPR3AM9LD
+ILng95QYMD5/btE2bjaX6KLczEIYU5x5+F17dFBOh7OJ+Z428nxLqkL3XoAKtgX
ahSlWAsAioA8j/aHbS6Li+A2HW2e2NRpxsKxDSUPBXG9di7YAWoxXmELy6a1GU1l
UffQbgymokqC39ptE217L+AA5NpseQc3qOL+GuSwBey6AAFpNe7zIP2eTHuQSfVe
AvAeBuewiRDX88rb4a6iPCmM7tTwocxW55wcWe/ad9+l7BpWou/8HYT6j+jNms+8
DkJoc9qzOVq1VNgypQDMmdz6C5Kvjlchkdb4YdetiB1gPL1u/M3naMWG5Rjp3xLQ
lokzdplUzK7oeosx7FsUz6cCn8FBsMo5WTDobUKm2waVZy76LoKJ3qP092DR10LB
hdBsEu9CZblHxAjQw3pjhd8+atfxbJs1xPzCY2MzU8/3GWHQXXT9ZlNUBPwfpnap
9inxkK3bqSA4K8wSrtAD6aLYFvmZSPMyTJYIoNPqg9Vb6uODrtUD9DMtiyhYXcOM
IqmCFm8dyFHA4KoY86ohb5RycVf8TAKXHmAjUpa74BEBOnZpB14M7oXk0Ebb79OI
AICfhknLcsHTK+OOuInG1/S7pol4COujUOzjcPaDWLw5weLA+3tpwDv+qHlvlRsF
uKikiGmaA6ilSJS4owkYxxbsyz5/7W2JNEJW3IZflDMdh/oXkxOmsbsILTQSdpsI
7FCnVYyG3lgjVAANruynjUDaS0PNPCAVpJTBVtCqT3xG46Cps5fvpQQkOAsoamrP
ryRFmuaMgWl9KSoO1XN6GsEYObVtpOwqwtGTq58UuTCo+Zhyj/pO8TEoJ9GW2BF4
mwAowsLXVukVvy9oZ2zMCfTUSiu60EoL1rEmLWHfP0Fltyu+WCYIAP0jMZ8koJ3e
sjLuxtVkpK0qMTlUXkGYzdq5dWFYYfhY36Mr8Q5Uj9iMhaP1u3NxFXPzLGgcb5g4
DrnqWWiwO0wr3AjJYs5Z3pUqYOv8jSe8Jjyy7YFIFoaL50yrF8MvkscNXLUOeggI
PEB3nOOgmV0HxRnkI+XCZJPi3Hs08eQJDTI2USCbyp9aKBNRe6c76kDF3FJFwHsY
xE0y/zX65009MI7K221iybV4dRZnolTgc2VysPVUAWf8Oo3Tc7e4oXF/rFcKMEhM
MdDUTd2XQ2flQPpUylqla4m9BSbpA/ogIDuPzqAeRq8VW0pP+YnbyTYHwZXzaqK8
v4MtlfOpiGS5JjwG+0SfKMDJPLOqdsgJGhM2/cIFv86lH4QDbBPq8q0rWuuZsD0n
1pbA5q8RtXiMfUahJjS1h6jBfUd/+uoqzYL5XKFEVKjvuP1bbMcUrhqyeA7RlH6e
U8C+4ooewK7pDJIe8Byrb57lFLV4kgEOBPSe/LPgqudBwia3GFzjx1FnfTUNUdRa
goKbUcs2TWW54t5rIn0B8cjk0ITOPclVrKWoPC4JyRbelckZBo0Xz94iUhUkqZph
YN6Exsb+QYcJDdqr1ZPYyD6BJqGcDgMfsnN+y3dvRe745zbWszTGTamee80ffX7E
7xd/l6hufuvYRgqIwR0ntKhrL5LUdjC/UBETBI3d7G6rIXu7qzoj5mOVGNKtWPmK
ghflB6h/66tuy7fbaadz6oN68ZHBShKk6MiSCc7X274Us5u979Eg1kLRHrAWotUK
z2DBusb3GRGPbeHdsr6D6Tlwj8+HwIqFn9SG3rTmNGQF6mS03WHCxBFccV+YPKOI
HbwjcqikbxsCYI2V0OnOBPVBM3lCz3frAYLXSC+aYsV9bcYR7K5UkLpkhUj3y0Wg
D/gO6bNuXjSOdwh7ctGGRY9HdIbg2TebgiFjgfvLNeIKanXJYzPDf/mUF6JSSijC
ogeZScDhn7WokB/nNxbO7qxlxPZGvqglaZxW1Bgd0oCJG+NNXcTBVsThrej9V1Ze
mlTqySDeegZtplSWSzD11iCqQe/uQpgpUReE7tDwBGJMP048XezQXsUsHlxz5kN2
/HpBRPd9yluqDbuNVOFUwhw/sytuUAPTnkVV/iOI6EW6zG3DKKtxOT8T5UmUPi6D
71D8t1UAWuofSmGyk83A9EgA5zZf6K2vj9elp7YupeN8nZUX4CSTJbOuejPUD1Ly
GDBLzKp1wfO6XnRF7biCQlLCELVm7p8DMuWSAPMAfRaQ40yWZECbL51PMgiRlalQ
5ZnLHryR1hn6vbYPIxIW8cypLaAuF7NaLD3aR5gFL68e3dqsz3AjEih4gf/GkWS+
yVuzayGXkoRZa3LtCXsaCH0950nwoOvrBIJSbsc3ozIEalctKScoyICZyel5LUpw
XBIkForCGyVjOVeYwFAMDMXjDGu0HkAc5cwzmY/mqml5DeObS/WcEjhwes5XLNUw
lKN1ztxZNEvkfvDnoqlv/wM7aOOmNWwGKVjjmF6u9/yMLbANe63kLHWZsr1Odtuj
rmwzTCxwsdaGbSoZzwMzhri5TE+dBasvs75YOHPci48MrzkqdP8K1dnvq2sK36Dj
DfvQraa5qGmGeAaddjh8rm31gGUus9M0hL0YcZBxFc5aAziSLWvvKOX3K87BGB3t
PNRNw5O5GIWE1zpc4HFwYQZbvn0JVHY4B7MhKJHAKL4abtdDpb/WMoMcZXIggmIE
sHaeMq0fHvYbP3kvHE2vJVVQOMepwKdXhdBgxrQ/fd5aIxAuEUCrNLTWo+6+1S7L
Lubx272YQt0Oxg8m0Ed0mrlpSoikgZmGT0gqHSWjcSiqTuAkiJgd35bhtw0Bb+1D
wXo+pZGDef1IczaEWM5WSQ47rFU+w+M1bH4RZkkRTjF8KPdIdPeIPchxxWqKYfkm
GVkjvvCnXsAx9TY/kzGcqrrTTrIQZNDVYyBYJzVpGSHsVD4lW3tiEsfjWHyZSZTz
sXhIBf+uERZCHwV9fS5UnSJHOmXIhTUIt2mPLRsxdOx4t9WcG3xuQn8lqEaYRyqs
H0pEeuWmgUgOlPdFi8QuiDkQtciGx1cCAYgCFkxF5qqU2xx3pPsGJoqzh7zRlwQ0
tRah4wnK2lEmHKtx2pvsFP7PcEg39CvuuDPmpcsOtKTdCfEvJBkdky/YxTL+Rl+c
MFXtFG7BDq18416U2vNdZ97XLg9AzabD9Y/cRxbZMzx+95a3wRrNQnCICyePt83e
mKnF6hE6qF4Q+k3lkI7wHFr+CN0aI/B1pdA2lMsavE2Hgp89EVjkNn3P2ON4eocc
KWajD9toLfImTz0r1qqnuECrgofCsWNHWWZ5qtx0sZdk6RKX8WPXcIRyO+qLwXZ3
steBSGwzhycr28gxuQJ00X8zGTI8XN4RSwP3gG1OfcgUfNSEnyX1gTEeU3EGzUjo
Auqx7chEiNgvDLCy6ugxcpDICvcqshQw0hmDSJdYx5bevXUg2kgshHZJD30ONu11
H9soqG8z4av92JP0LIraeLg2s8DRoqzNV6TKbdmd/NLBWBuDQmCGdfso3FyPY3Ae
6+k5hMy661ir7BB4sce152zb67PkxLil3/THy64AZt5MGCNcsnPYF/6ziNwcFh+Q
MzMpQh8kmI2rBeV+IofZ/vXUw3PUpla6fT/2kjZqUqot4E9zK/iSWTOg/R+Bw/eg
xPuk1O2QHR0Uc4pHFIy8101si26YZLlvyWH9caKZRWDKOsVtLlRlvE54udqrNmRS
q0JVGhiYqD0c2gKKCAcd2yGHygkozYzDb3TWkXII2TO/jeM1KBEEyPOz2gb6I6Bn
T27cbUqLq0kCVu6JQCsv5u8taEx6h7xxPFxnP1ocqCtZZggaZfSqD86iHOw2W9Ae
6tWlgWROk0kHeEnbG89p9nxnAFehqmtB3hqxEK9HoO9FMws0aHGtz3DIbfXPj5ZB
T4mDDt8sy4wAWKlc6XRMuqmeDjPZJPAd06h01OODexjFg1gsilHyItLdNfoCbh75
VdguR4B8sWrfmuRDTibnJk7T53U/PI4m6Rm6jT17bAU+oZAR5S5TPgnH0K+bcl7x
3s/fZAIqt74cUjLasi35moTWc4dJpZEPeK31sm91M9jK6pJmxpPQ13dTEKklpvjf
fPGvsYrgp063xtDRD0ZLdvnYNDNIGcCLXaziZanoCI1lSWxGNf2vf0Ierk3CxPRi
k4NwO1pbubeibkuBM+N7zmLezHWNwrJdgUuTqrazNm6putvmFXz0aE+QljUUtKCA
rUs8gpp1u5GahdIGecbI5gPpYroK7afKxg70igdDvw9K6HZj0UFa/4S/5ieVe7gk
DRrEu+BIfkMRifB0eMCLvfBTfUv9slUqgQe8q3Jxxxrg3pFoTv2azIsSy9L75v4S
Xah0ob/Nk+abMpH+cKOeSO9j6zhIIfZEbsBJABxGRuFFUOlH+bmgues2RAEio2gf
Oiy+93mNb52bPjkdyD9VQhWKH0V6GN0+5TU3SCfFwgeR6f1fFcs4101K/M63tzVb
0bTKmDDfwQdxaXjgWmhLvQQr/+WNsgjcu09dPnKsJePrrgtp2SbaMS+LdFNjFoz/
uHV1pC/2rvA8d5x+PeTh5JsoaNK5+Imx4eH4kIp8DAVnW8f7zPsDchoKXeZbOrBv
5RXWP5VDEHLh1CVHXxB2aOT9zdMZpgWg3MsxyGDvQs2LPnoyW+GUBoEXqUndrgDj
IYImNAM2eFda04xtpXMzKwbBsywVwx+1BE8UBwysCfOIuU6DYIUa0AzObBrf+zJE
OAYuc1U+oTqj5c/5XLJloZNpBrws4O2lqoedCuKaPQ5nnzEn0LfgOoXmn3q749ia
v7RJRXojZqZBz2SAc902a8PvAQ9olr8DM+0sq3SpIdouj+vYyn8NwsvR/ySNx67t
wAMa+qt9vth8fVtOZJ/EmhQzINRkBt+kbjcvXYdLHkulQvhgU+ptQzuVfuiQ911I
1+jhh5vT5Mdm36XkY9B/jHU+FnImEobz9hZUw4aOHsm3p/ev0U+N7U0oZDCVtY7a
xJUDKVGWoxsMRfpl0ATAUvK9nTNpuMfCzq2a3i3C+st1Yoon45pMBMvuIYjzFb3i
/jGkI8s6OX1JMkZqdw2Tbm1V/TF3g/lerlNZEwNIBYST5ak4AD2AIydKH6xGUBaV
UORmU/mbYr/397upWW0SzuwM1VQCVGWaUHz2OWNKr+En+kacalzKarVFKWgZbmXK
L5qC0ZxSgegDQLz5Gt7QCnw6fjunEL7gaJ724tAIpFtOnAPlJmVDiAt3tpm56Oo2
TXPr3jq95p9qk9OHBTb3jQb83LU90tSBu1d/6DThOH96BxJrVAOljaaHpx++FXzU
By1ZDr9b5R267o0X9kdeGuQIZznlZuCGurFmEG/tZVnU2qQ49m3Xmf9rdpnvGlXm
9D9O/+W7faL+on0wykOYX7bhT1qDkKSgdE8P5YUyx4zoGPypZP0APBW7yVZ5ZpZM
79SZ7GW6TWCJOWFU52GucUaBOr1cerN3FXxFyRrKJ2wgAW2MIQQXcKNcDrA4FTxf
jrClrgSXMmeY6ETBdU3yGiihFp309NMNtFSevld/1xt8OF9PwQdrMbrv0mKMxQ0U
gCKVMkkH0cTB0t1JnKPZ7FSXGHw2y0u5gLkxgc7oIqQdJXJFzDpKGYU1lkFpUAC/
Wfuzy+N9qOW9MaHeBBcrK47hLKf69ZwVwYjmcy6CNt4nCaEnNZo8YIDKGiHBmy40
SJ1hCnSGJ954iSDCv5AK6/AQWin4D2mSZw422qosIGfB2U8DYcIT5JHA1nNEbp+P
HNTlFGTa4RHnBrLJatVvwCi8vikZIgA8TOBStUFF2+Qksv7ClDn3sJJbLohALkS+
Uij2RF1N1m8d7Y8qmoLPaiv0vmrMUMPPmn/K3L/s5Eqq9XZiJfj6Igp3bSLoyeXm
PIQryl6DzECu3dFxc+7+8vrwAx5/lcjVvNaiJTe0HQ9jHRvQz1f2W0/vXdTJLet0
ycNhctfBqM5j6DQ9BFxzJGIz9RXteep44m85lyPUi6pqUmLLvVNJhIFOhZRUiUYQ
VzNt9koIBhkXPzddkHX/h1wRSV0NpfQXK8GH3+7c5BT2/XHYmhAlfE9ylvs7y173
UjgNI3G5EIC9vrGOmxcTHU8ytcrYKJQZ84Wh98qgAu4np9zEWOtrnen36D/q7/AJ
ZD9UyYATvg5KRPaLnFqMEx0ftFZcjcBmrUzI4isLQzqWeWJjRhRP+uXV+vQx2/Cz
WPx41RvkFFTRPd0K791LSZdgCG8teBqdtbhWu9PwMbRAue+Q4WNUV3/MlyRzIL+U
x4aDAfeQL5TSJekHTCvYoJ0yPQlOFV4ZSlcMeca5EOmdFrXlw0RSiSD3DXW2nqsk
4ooSWWDi7deugQ1x4kEUDA9u3mkaPPjFwn5IeWU9WJFsVZFMJLXZUJ5410iCOEA5
Vf2dLNv4kXSbIkyFESseOAOxmlYiR+LBE2wrcRoC5uO2M3M0ta1oD+zCOqs3LP2I
O0XVrlq8FkqQeBIRypNc/+XmzrqQAy9fPUmDig3FHPBoOyU6OfXxqCYX2X9P7EtH
6CTxIBzozheavmO3S93b8sBXEzMu8HqplAdRDZmUDlgABr91RYw+b18bSHsq1/8N
G1JOMfk7ce2+emZG/XwqlDtd3laqGONNIwfKRsCjoyqCPNCjgsqqxeK+Q3kzcMVr
v4UcJScnl4KbF6LzT54MAdsI3L9C8lUpIlpGWbMYAKbb2tQoQg9ScEy5nsZ5d6/n
Ki0NPEjq0+vabWNAnA+II3yg8Xl1zkA/qSK66xzFtKz0AaBQ4z7L5Hbt60n0YyEu
rllpvdNG/Ry62f/H0qLzl2MD9jfCi9o8U9Umjz8djK9sHCjRkzmcRwszQfkiOT51
iLOJBzbhYZ8ZSTVGL///dhsR9hjIlSdB0fFDqsVJ4C7b2YdhRYblxz10jGpIJP3Q
oGF/eQ2WwnLVpPV2N9vkBLqBq25e/PJS4PFZyD6gv5FUeX/2xWxOVRobPNmNmyDU
mLGBP7OFNBhlN8gs5bYgVnT7IRkGkdDU+SfsbOLMbLUwP96i/pBdKBOgqru3Pwg6
4hXv7qGSHKes5wbLtfV2aJs5rwIez21U3G7ZZcAmaDZyn1VjlwTIdY3GLqUcyMaO
sajpu/KjpovQe1mC8cIv7ogs9ggHe6mZ2iLQitk0WhlSMpOaAIgkRVt+NHLCvl4y
vD7Pw2uBEiSxCxrccqB4JfbfIyAbUyh7ZMJIwycvmQosj14sfWQbyo3Cfi4mzu6N
yFSXb0tEmSeCmNThD5N8NxKyO+oUfcU2xXuMypVy1CZ6EJg9g6Y9yvEXZ9TSRed2
gOaewQzTz2KZIBs/dHnZzX5YIArwDfYOm/UoS2Ti6VJktPr0uL/8uRdMJGAd7/9u
5cACI3JiJgnJF/EKPqRTZ73c5D72mPi/yedBfGlqrat/lkmxVAtfydupgqPGRzij
IzWk6BFBXQEYWHDQE9GL9NlB+2bOLwAectRM3hDmPS/94f0tHEnNEopLNwM2XTZm
n4AWyXdgrBET1ICGPnyMIK6Q/BmLeX24rpmLuxyy1nHTiDpiDDlE867O9uHshC2K
l5tasOdEjOHIeUvU3bWf/KY1vveoMSlhjGzgvMi4bH1aphtz8n5GvKu+OfA0dZCu
t0sz9iCTV4i2fE25K835rxUJfTlKoQiTAtjB10D9hqxTUkHJEuynWqyLYaNoSC4S
TVJqmLA0uX93UhOphFlRgLyk8M2oz1Vz5GHPjZEXMHL51YXxpQz6Z1zrnr96YE3V
qqnpObvsl1M21DhCQrQ5XC4qUAFH0Df9pUq3z5EUyLJXvA2YdtObWTIXoT3km/+j
TUfBHSYJesfHk3slOLGbiqTo1Y1qFV3+idG3Va+j88114l0a6shNmJ7/Nfi6MjQx
zbjafM/ZIaft0BtiT++MMrVpssvX81u6VKq1CcPx57/i/4CiNVKrxSoP8YrhgHqk
UdJycVcfkHAA2LFqQYeonbfWdXmWna3MjG5SnfDibZFsT9WOpEe26+3YG4LJNMsN
x3LlH7u+LvJf7nzHFY2vUVdDF1nJR7gB2c7P/XS+21SutbYv3ZQFa64VUJaU/yCE
neeI8/QBAoQhNiigKgUIsxLJhbGeVHReGKMX/1cMPhzzLKdX+bIwlfLstImbXQR5
EusiSKqCMf0eb2o2btNbBuDsbHVEzfIPQP+JkXZRyoeCZh+RNk97YndLm5U0uCzC
+RTM6qec/FSLi0I00ToNZEZIbu5a8BSCCW051TkfK67SdompnFkoWM7eBYaQjX2G
2Q2X5uJS8XF0vNizLBMneDB5hXnoHi5J2XdfXuzPxVFjukSFbivOzQsKfqhpAf3L
uzl53ofkIX/8CBPxMbyP8+T17FcZ5bSGihxCeNmKzzziFWIcJJKL3ohCuxBNr7wY
3OwoaD4JmAP957/bmpdUEifsEIajWhShaxOgAFo+fysdzWLC9JYY0zqWiiJMucrq
pclLI3EUUpuu+m07pPa5r+8m8iX8YhkBRJW8On9TfIclLOOvD6DiN/OWE2DhfD7x
FtlLVg0mFM+74yS8CE8M7BYaV09G7nw4x39hzBXhB5QUfr2+KIuHRL4dfVcrgph2
K7HUCpfspOpzcPFA5A6mQdz3l5gPeJQNFNgH9Z4uLlMdNZR9HeepYil8p19+iDhl
uo7pVsYFK51SDqyLvtcql1THxhkpmtUgLDSusUygA9Hnx022wDAGUN/55i3PA4my
CSumojtkiZmxGUfzYZ7k/LPh9O1RGL7/PdV7qIRhmc2L447p6dblgjDCDbycM8z6
XPdnouZUsyMD4OshOmSizQ60I8DxG7sRWJrT9tciQkfcwlW1HVU3aiRz8NBf9iwL
9bmNya9FNg0LscYbE7dSvL6ek6m/fOE904kH/VjOYPog/UsR3ZafFzaweYgnCfz6
Sexg4NhPb63zjPav4NeVt++fyZi02qzf+ml/oDUjZttLV1FA9lxSEes4ilIO+Z9n
u/mfL+AdOjOcJESu2megeLJWXzr49dA/Sxen6i5SmqpYTpy2XRNpWQcd+HvXqu3a
9nJEpDC/iV4mPfUe8de0VNXHMflWLeMAyLd7rRh6+SVCWGci1ai35ThhaPunYqpy
+yZgHXiUGZS2Nf7PYfuAud6oW+Zr4UvqiS7GLG8ofv7RLrZqyVhEqpEX2GqH9WS8
NyvhMEacDgPd5WS9SsPsgT8Y5djRm9jQd+RRLpWS2a8U5sP29GNLFtHUHtaJxMOZ
SjSpUREcC75o7YK38+sWtnPkMINZTK0pgadA+XH9JAHqvpuvga9bAI/j0hSCvT+j
A+Jl80R6RQII/qSwu6kN/btIOkOlybyte8Ru8BJqIha4DshuCe//EiiOD533oLe5
WCi6zfCi1eWopgFDfZ2ulsYxGRNdx3XYwtoiWQH9z/gZLsX18+4XSCvnBEe9DJur
0n84nwOXqlcQIqDlTG8oKURZFhEfug7LCW4JBJ8xVGAdsH32u4htCc2JLJn/DXEe
7//IQ6mfnRAb6b/BNvV57O7dpsNe64CaDhnKT9dfdN2TTAnO2Z4aOaBnnalRZfRw
t/Dp95bCzqNkacPiKwzcHWGwVvpGx4LQWvxdBRC/ocbuOUrImE3EeBUQhTRsM7e+
bNGleKYy9CJSRMTaiHGhrIsUcl11GgbE3LArMiO30NMBVCOHkHqw9gJ9b0BxTaUr
S51BfU4lvBJhdEmfWeoL2/vKt2F+lR2CHGxoBXKaGSvuDYbXZtKO31VrU57/pOp7
tNpBYaSJsBqMkJBWQ9VSwI64u8nmBQW4pmxSEYmyDHy+iuHOknrgYXd94phmSeIX
2yhlk7W8ATYaOI+O5e0GfKRtRs4WzoOHnKbnG/mnmVPihIu1j/j86zQm7dn/pZaB
n+J5uacTZBSaqP2vfjKDgK49HCAj/8nBqQnU/RciUI98jaC5NLIAESRAn02cv/zQ
O6C7BIKNFbhqfkQ91hMAJ0E1CcrrbvfCJA+JevYUZtbIVOUr4yoJTeoEo+UDrk2g
dQuzHB7isCPEOp58AK1Az4uKeMXx76K3DZDuDvu61062CEGUZi0CRxqbO3/15PrV
edTBi3g6I2zxmpkSOVZJT7ahPEMkiOQuUJnQb1wiKauO8npkm4EN6jG2uTdrEtsM
FIVtFTgtcx8khsqkvwb/kkqGsQQvHwutzVxqBygxrNJuAmXVufg5HiE/3IFweCD7
Fl7P+jRM4Rp6//K3T4xD7eLhTlRmYYO4hsUKW6APx9Neboxo60H3uOiKKpgzS5h8
Q3hb3WXDtwHXezPXV2gVcC+oJ7zYDhFWb1q93tPM34A/YyrKy4Lor2Ns6WSGDulk
72XwPy5G4pEEkFwxh9rmJwqv3kq8KpynEMS1GKxlWqs3gihxW9LELl32qoXH7FRL
Jn5oBUKou6LT7Ttzk7ejvgACBLT7LMiirKYiWELx8wBdxCZqFV0MIMrv/oTzd/eQ
HHZkxorj/xx8wPsyunk+IDRM05OwE10/9cKG669gmbrSWOGGAa/T4L5oZj/Nr+pZ
6stDWSkDfzMCTyYNvXKKnGrQx+KcN/FGpC0GLxSyNPJ4nIm2Uhk6KZxfW5b1U/++
QFadSM/GfepggZborFsWWfcRJC2q8qJuLIPuX05Z6NlaliugFHPK0wyvCWUvrSMn
itVtocrJE45ZDCq26CIMY9TMnLaWAnhViyoHS3T4pRWT+PDqvIH7cC81iwLl5sdE
M+6WefkaMW1AF9DMWoIsFbAnPDxJzqHjxUVovVD+dreoAfoDQ+kZ66oGqLmRp9g7
sg/NZ8k4rtDVD5v6p3dnd2PVr3ZaM0GQnbOq0jh51QKLaBEcHpw6c6Z2OOj+sV2A
2u+IrbAyQByKMlEFdXZtO6p/4Y41DByUXLGdaMvjtvAderNfSwjHiyv/6Lhbj3FT
kIOLKKNeEGG3THzCRBIA5PAlAgSXmgIsmDWmjHrCUTO5e1h+YUpcQv84JseqDuNs
Gg6hQI7OrxrL0jWXNKD01oi2OZSB5/etnErpz+fh6zEkRgyZz5KiaFMfoqH5gA7I
078/LzRpSiHuvXke/g5hqvghlN/XFGYUZxxEn2yVv6pQC8Ro2Pso+vWYVNT7E6lN
1i0jpzXQiSPe1SDgJGMSX2Mp4lZj7ytPH6cHB4ogUinaQgDydWUg1SIqUAphRGcK
AxDVujdKLKDcRp+oxL71v36AuAjqgUoZ9046UVRh/7YfCeJRj93cQLikkKE94JuP
UiS+RNR7/a2CUicLHG4xFHwKjID0pcCJN/NZ0Mpj106+5k0N0UM58j5en5W0oqG1
qwiQ/c3oZU6PJXZ4pPhPOjt6PhSYUkI0ETPu2za8Aqt7xzdtEy9aCqW9jMLV1Yw2
t5IR1D/BZX4lF1qt8AmoshyNEE4Mh7rHjGPBi3BFyHqTfAYp8GchzKT38yDQOEZ8
HG9hWGUgYZLSTruFLP+HR0GwXn/d73d3Y2qpcuTD8EprViy7wk4OFNLptOrd4f6X
SBUBJoXI3kUHmn11MutkFrDAeRj1PhyX5JA9znuTPId1vNgSTEBqwg8z06XpacPt
Yn69V2cNlzyRjRVPCRipMHA5p1ytC3sYmYQ/tXjGgkqpxghId2akBjVpiEWAv9FK
EVfgW/bDRc2eAUAYjeFwVTd2mAFb/uw4aTXckXqoj6LkUdfopa8bWiQ8b5ig1TdS
Yauy9ci/MM90T3hZTWB0Zn4FRj1qhiQ0dgUPUJ/MirwcaFt83jmJYR3wS1ThgB81
orZiO9drmEaQhSkBqJfw03pgGEfoTvLXBSJpGXEGAurXc7MtCUMXvuk43OrO+86j
bkSr4no/C3bSLRHqGW48fz4HnrmUvwfR4QFMp12DutT03NzNwrugXiu9AatDWkh3
VV9CgWU2LVaURk/ilFWynKrt0N5BpexPOh+7Kue4NK7PAnqmx3lvK8b68xDWNGB5
O8WfXDlW8hoZu+xAufLI6468mh4STXvaGaqIQ7RKy6TzyGFYeN+K2RYKkYF7GZHu
Jq6at2pccT8g2A5Ln+kKPiVc4DBdBGD0+WLBw5FHyVOF+Xs//rRsm/17gdZTRjIm
kKN08I7Yc2TgglySWbo/WkKqx53ldhe5zk4Laz5JuZD0cUP0vVSALaTZIZOCDQvm
T03kydqrJ6B6lz+4HRGwyhxqrrXlXpom7xD4mh5dX3vpFzpLXLv4O5DJTN6gPdTU
H0zlCOmEajJAPfUcClvslgZG1oKXqZU12L6HFDhLHTEhhv/yd2Nf7ak7hUnTIT/W
KNFucefsMGlDVIYBkcP87cCO2yzykUZVFV8vXfQfELxujvb6QHXJrszzaWgZnhR7
mrZ+Dz1/TC0LyXFktHNJQo20JzRNS0KmStJXalQ/FViVMo/otZ/e5ND08TAY3aEy
6jFu4VrYGg5aZB+DABQ3ojijq0oQ09Hcswbl0X4mlwRl9qgOOiV9dLu5XyqZf/La
i2flz9fVicQdWk0MUdBgoghaxuK45rDcOzX1FK/2JokU2CW6xxnFPmfFPofbMZ+D
o3jP8dFLKsr0st4dRoDl7psUog8Y2tolKRlwptaRZJfHChZse3qNwWXXxi2PYqCO
q193L9IbeJrjib1WcOeTTVYk0O0tlZyPtxdcwx8TFGNH+WH0hWTDMY+47AZyre+Y
D3w62VGA9oLpgDx/R2dKO3INnXJdtc3WmHnSM0/aDhm9tnP1GaXr4pJcbzqGKCcK
Aj7ja5YJ8IpBKTyuPZh3e9ymG3sA1beDKvAfQkAnMkXrqB3uyFSlRVveqCXm/eeb
CTtTs1Y7Bu/+YL5/QLbXNMktjbk8jHfMv1FkUw04fjP4IXFSDbgk3jJJMuYs6VkF
m78jXSF/XpX0zVk5wBXth79lTcesrB6WM6312y0CPj6s0OiCv6+/5OP01euHNLzW
Wi8b4N4U5nG7sXNwBr/WlS7J3F/tgBO18D/yKDPjaH8rmno62LY3HvA3dmevYp0W
RVjRT5T6b4ReFZgRVMX5k/xQ0R7249VrTKmIJCu1u7L1GUujOxdQQrCYs7efc36Z
EyCkdhSybJNf08/+VncJS6smwTMJgAQ3AnobdtyEeYgIZdl0+Bi06BnDxkd3ke08
fgcZdZdfFGX+8yiOcPY5gmL03YdN0jEtULC+37x41mjT1lgkwLkjPxphkjDLQawx
uzzb/jflmuIAR3olbLsdL/6PcWTBUhlIia68j4aL4m5qy+TynSA+cFkNTKQbIHM6
AjSN/O385jOv+Y+M4sEwLcPDtKgrDXrSv+JmD8kRCdnhqdfk1XvWqnp8Qd4EXqrD
gXuqrFb2W5dGg+N8mfpUD4eqUjRtAVv23DXAVE9k+TtKhJBQZi61oTvYT1uvPwLL
m3VA4NWzanUsALajmJNbNUqkpcfpw+sGadAe6c3elZpukiLVrY5PvDlDYK/+p/Zl
xJxjmHNh6zpMTHYsfx7PZHMTn8Nj1xOzr4vTo9RwGyY/pj75zEazhBsN8pi1GbYq
g95zUdJouCk7QKf+2iFsgWLZ+uVRDYH2uCvX4Y+A8OGBsEhELXMUVC1Ff4ZjGO1x
tnPC1LAdE1Od1ldPLBQH+vnIjM0ltRLKaH798+ZKi1zSQvJNppIJ6GDN2nJeWIPd
hPOlI7Z1AST1vrnESqRbsXTgCH4CQh5DnVwpxug6k5C0oiGgWMYbxLLZY2uOyFS6
BzQ1HCwdO1lAkg0HDDjQ34rtWqQrtrJ8jbXi+3sbY7HV76SpjF+s9eUJ8ciqyMyK
nbVwmmJYXCgJf9mMVkeyamlwkanLX54nfKs2ujuM/WRSeF9ZLL/+kd6dF6KPMeII
nAPe0o/1u0cW0d/qJJ5s4qV66knmvCh0aXl6rZI9v5kmTy959SWsdJDK32BBa5P9
g1jm/mdA+TI8B8n/LAoiWyAIC3GyvaXvN55sEGFCr6+X8Im200oe2+oIx9CUS39e
chM5lHFPhvB32LQffOk/jAm806K9CfJjybWIdwCjivc0wlkhDowxdTG2UNcf+Uwy
fJbzgFxEFyKLYSdhVh34wQmDQSrkJ+nGeJi91+j+ZsDrwfYNRr8kOd5mfOD1wBV4
etT5yVVx+a0072OikjbIKhS8gd4EOe/Tkg69T/yQ/jmbx1FjWhNS5FKVKUzIvTA/
iOgPpw0+IwE9a7f7MZtFCRZMBEYotizfGvPLXKHDbWe5ci9yZTUlMLjeIhmhAXbf
K7sIwpeHCH87b5lzn5ZEdFvpNYBPDy/MkPRtgRhQ+ruYASGHETVQq2EAgFB9FONH
Kq1vE1nL6wCWO9LpL11qXhRENJn/ZY00JRiBG1/hzhyPLQXRpVqvaMnTnvVjk0m6
y7mROryihkcg06/W57nXWyBRt3y8UAFCmZEJzksnmWisrFvZFtvMLsKu9tMEWVEp
4BYAmwj7PmYYvMw+xT8KPF+PcI9f/j2iDVi/zEFU93ky+YcR/Ce03y5ZfHRfk4YE
oh7k2JfHc63WKOpm3MY3jadfqwOZaXO2zPAjtV/6EeEDqZkoiCoKRU44LU3XcXbI
Gl60I0VHJppLkoOygTh3Wjg7P3hkjNn3iATOCLMynV/OxFx+1OxenDcL/xDGOGnX
lLFAWz99w/8kVbxsk1svuv8sDKxWRCrUNXkMd/uvKyrryWEOpXkVcNAS4ulMfAgQ
wQ6CX1rEAcoNxw+78yCAuMClR6VX0Xl3BPFNQQY4ysD1aVIc0fSPeMkTJFZCXx9b
hAhsFuPmQv9wKjboRTr9DqnKOT5R73mjRGAvHfFzmDA6/cPDjhPknJDOPIjXYARX
hlSr4zYizdaacJN+7VT9bVXLceOKJ5n7wSAdjk4PXtMgYHhDld495SjvIT3DXGzE
b9b9YPW5lXLfEqjiHy7Aifp8vnZz9M1wevCYQU9Jmr8DC6EiatvyA3uhwYEqAuwB
sbSOrvgY365JiM3Bc3LRKIRevIpUTixw+7bpoPRFFp/qQWozZGVDXWkvuyMkQkLv
JRrdgz1By15bwiImWxd76KM1fxIwyydf0/52LZdBxYnz1Z/xLz+nSf9sGJGuW78u
V9J3zXSTLlFZeQ2t/AZ55+mDCOgj0N13+jVkpFA6sNKNRbphBazqz7lX/cnvoaNi
DSJpDjSrHM+ty1gOjHCBaqjlQEpWzTW0tbkDxRao2fivfxbiLE+5pdKeO00r5PFs
kQvRXVb4rpklB6BKRomQHk3rgU0Von5VLDTBI+WO/13de+K2z5VIE+V66NDSuibw
+OReQt787THMrt6xAjOluMKNPKnxmD8jbMo9AkXHSdYt/y3w8A1ovRVm/AUCEarj
bZMUVCcGtR+BmEGOinjtT4o8UtYDRIZc0ZSci1s0Ht+axwcDddDrItz1DUPCzfDv
EZaM76AeZnFbqqH42ZCHoNFTkNcur6m69RDft8GeCOhg2NE47w1vc1q10RTMZJel
pZzCMANey/1x8B7jCKSVRjyGd2Dhxzxun1B6rFxyHZs5wSqLAKe5XQbjflvtJSWq
pYnU8vrm5Vk7wb/3sCTLWAs64oKGfXvRThAfYR7ScNQ/cYB46Zeg9GWLjpz5hnm/
qTVrVWYGjiI8FpkFgTs2siw/OU1Wzxtiisn1G9Sqr6XcT1fCw+GAjqL9IpeCoev5
RGlDKbyednn1KErPjT2pzvni6udZw2ZXzI+BmnGQGSV6jLwz5zgwWcP3UzINLCO0
seYj9iwSrtvtmUNAGbNE07PdsMWsszDneSmkt5ax4o1/oHim280PYMqALp508CBB
SNI/oaNaK0O6oLkbgOBbtIFAC3Mb6iDecLxJkvEuRbiJvV6zmPKRMuakJPhA5bdu
Qg3u//2PZvI7byPRTRzxvGo6Jw/uOONrr5bNDfQa3fyNBhYUoLLEks8IxBqGbTZQ
ua4zwgnDv8jZxb+6jP/vLfpb0wlg12OOZl3m6xk0AVZT03NTtZ7txm3xfrelSK32
UOYWxwYGG53pHy2JXIrazQbt+EB4/RUodfxMUsdmtA0ttiDRh5STdw6Rv0dc3Ide
PBubMAorpUVb/WMsuYsI8WVFRKyXvKvt9O1JZovmSXWfi7AcqJ9wP1/MblfagvmC
tLEw6jMYQtXEGq4Bj6dtikKLZQxDtg+sbjJ1hrv5GiHdNSMyg+y5EW+LFQFpQMLJ
obmGcnIDC90DS2iBQ3WihDkHm2GCMNkW/wcxc5Y7TChBCxjLhNMDoY8Y0aEwUSpA
xFp+eDTDetZs95Z+ZX1TVqFVXkk7wdsG3K7OdiCatYcphRp4//tpNVGXJEZj2U6B
RN1kkojRM8VBPcAOauqhX/bzzbJemRxi8EZ63U2U+XzAF4p9h6+r5lOxWuxQ3gh0
gZvLeaSItE7//BVwzWiSanbBUZRx8FwTJnOnk3uqlIJcYoPclsBPdB/p22alnDEV
LLUaWyKApRruEJdhkRYgwLi2iCQ5uXWdCtMA+TgWiYS08dzodnXizqkLthww11/8
lM1EikB8w2YmYHnEj54zW6cjBXPt1vCqf1rwPLZUDPK3/hjBt2LHu2zq5wiWA+bL
x0dqpVHsXPzSJX9/KDUQOw6BJhUU/RprGQ47ZUxY0RvQbumNuvaJiHnF6xot3IGO
fej/vhKUbcpKkbyAYVtGpIjijhJTfyg/ozyMv+vbqOX9JlYz72YPE5VJCExyMkci
x5oz6VL8MqSrPk/Izv4hJazFSP/2ViZYgmiOYQtWbzdKOrcbdqWSB67qtmPvBmUk
8HXEx4SiKNnIVfMxG0C3kFvIsdcdIOa5GQV2oo1FgI+unDuMMMuE5e0VXdCUZ3Uy
v9mTo1AC4HZkitf4s7aFOv2MNsGOTn0wV3r9m4gfS6dGRNbyxUR58xmD1/z7OvAy
r6FU2wPcdH/YJyJxvRe94aBJHtgh6tFRU2drndudCM+K/ba3Spod0pXjTI3QnLrB
uvanLLsvSD3oEJpijMAHoh+EmKGw0zqA6lucBVb1V3zqnJS3aIB/dV+zKNPPQD9C
eCe5Uaz1tQRyGQKQ+h9wxU8zJ6h08v7hVNNuuG9eXIEJPihK30iYfPiGbFdonXIj
wlgcEIBKHJuRRCfbzd/AnEN30emY9Nfy2Xm/50jdQVI+edPxmRNJJLJ2sjxvmHet
EeDvcKvw0A33gtCkss/2H8RLS0TFnuNp9ZmPzokO64iyVqfJPqn3JKFN1JsxYSYx
NWyqjApbvphsAHap+bUlsI1SnIWbWS+wmGKEkYDyIXVbFgC4o0aPFjtN8n7zi1nf
vMEcILrqblAkgD+Cj0lZjyWmNXmFf/eHvvnCcnEIKL5T6cMMJ4NvhC+NwgLzn4iV
T27pSjSEQJAF0Ja0sAgbMtbJ2YK6nTTZ+wyZGS5FwEyPVdmlIQZ3vm53+E0X9oVf
/vaPG1sjH8La1QTXYOghU8ECaWgwBfdfUqWROLR258YRsn34WER/dGkzCCmUxHMZ
3zmfvH5FR5m59DpZRTVIUdgEI4UbqTIOZBHU0Ty1Tk3hPqhYwuQr1fZU8LBeH/xP
c1wzuH8oJNkUEjyqhLK1qOen+ANU+6hgRrHdREi0m7Jp30fyvDlHBlDhbwXP7wui
If7w0ynGi9ttflcFO3KOwumBnUlXQRqdeJRRuvUrv5gEuZxlkwE3cpLWfmo20Za4
CSnSRf0SDfskJwoXbcgyZWWM2UkYWr98aI3T4zblpRdldAWoL5soem16ImHNKUpt
yAF28jN42r3WSc8EtiWL7FQcpumg3CD7BMCfK4/P6mhQr64I4LebkxSd53WKhJh+
QPQeOAhXAXOEpwV1u1rcFukymfZfGtnMtEaf3DIgHJKREFVMgDwb3Ue2ZP+ZEOK/
S7jjnaG3lozeDeBrZtarxxmzzwyg00Z1fGeHeWvuc1aFNQPpgLl+Ck7e+vDRKpq9
IGywx6MAo7OyC2LAaeKW1ELfo5+RJRO6gUcMu5pCUyzqZSh/eUmePV5Rd0Y7qiwF
aa2vhapJ4uLqz6RToGXFMOlslEMcJIhfTjSQ7xJl2pP7GnuARSe1JLvJoRPoJRC1
81kfW7s48w2SOriEMGh0fO4ooIRRZFPZaRrwqBfXzJLF6doHexL9qaOV7LzRK3Yj
RHlidZZPrk1r/8odBhuRe07XtExNAxgAzsaxveVoThOaolKb7DIB47RAoW7nkWQy
xfBaFG3xqfpoiDgTA6DwhH19kH/XNYHAnM6u2dWZuycRg2zfcac0OuztlL+ScLhn
pftfxLAw/DgrtYLcT8fCTQB5JB2qQIaSwNeaS5KBRRNUW5KaRFLlq2ETqehpOfav
3qo2ed+DpBWzgs5M4plWCqjcH1Es4W7o0M7/5w/H+mLelE1DUTUOPZu4iW6HmemJ
yIQy/TK83Wtpp9YfepG84dH/cxHnnhc9IhTeMnf3xy10souh+rgsg//5t4Ku0mOC
rWLdAdkdDUeCwKC0OFwJDkmo51J+QTeMaGTBqC69ZO7BQOiWKQkjMwN1ZKdf9mA/
jszWhrCUHBWOgx6YZD61udIFOvjxB6Jx0SDrOVETERrEK1RMkmvaZySbOlBlbgms
MYsY7/yyb1ywFknSXUQ1mkarMEmfYIyAeI/uV5nvvR+ALOT+20lo3CPNpoEVTpcb
xoy99lYcxUE9mXXGuq1I05rcBuFLMEe8GtVR285OSkB/487I6col0hF3geiiLbcE
39wLdBveuxE9fkAgq7npenBqm5bpibY3+/CdDdLycL658YyVbDiaYgRfVsp2/+Et
i499xWlGcnJrxvbOHHWxFoVg7SrCfZJxLhP/Z6WvklS5Y+1wnwQk1G5RWRnE426C
F7g1q+5yZB5zsH0+bFuz76uy2z9/Hse0xYUfaVIQYigvLKHakoV8HjPby3oErVeB
SJ4szxAYU7S8+tnPXNNRNgg4+NOT1U5GP5O/ephfWsDLvmcIvw/CN7bxv1P9Cj6F
45ppoOdQfFw8BgCkSdaDVwCZfYNL0pDxGJ1xj9iYUMM1dqpqVgo1FVWpfWSAETLQ
Tzo7gUWmOf0Cl6+6cVBLwSLXoUdQCO2zqIn3toc+MNkY7sFFEnVqkqJ4HHC60IBp
kLmUYnEeF0mnKdknidOlU0JcxrMxY93GHovZxHyqkAQH2dNpFANeho8x9dgZehVt
9Zg1J7C6wxlX0uOniCoaGrZ4iZdoYLkYbbjKJdoxZV/wi1dp3R/qCAaukCh9aBTU
/I+t5pENI16h481NxMQotwIEHStLUEu9IVT+7Ba+6gcC178ieMT2a280g2/MMjOs
ku1KKE5vk7McAX8VUNL9hXhMTzGHHISpwcCTvEUxnCcBZqkXLGhl/+FOT8bUvTGg
UKcklp/aK6OBQfhQ2IpddM9eseJclbFCvhB0HEcsK0mAd6wM2UXrKjakkSzqMhEk
oVyO9gRAYWM1MQau0bpmHMdbI5dAdS9khQAcJKvrb3z/+9jK4qDA0Uu92huEsy+r
D98fOceaOMDpoTgqzg+zxsQFthV6RQv9tLw+mLVUh6Pcz4f4hhPZd2ZYAji0ZtmY
XtAagX3Zo6V0embUzu8VTnZ34uRguobXW/Whf9b1W+tutawLeTta3MOvSIVgjsXr
PDBamLrLNFxl5yqwC+uEgH2DUBJDIozzs4zoePWyP/oilMeu7iKNkn2Xd/HU5sQt
CzDTSUyfgaKJP/EFnFp9yeZk/o4BuQE6gM9jeQvWe5TGAWL3HUXTLPeMgVjtxJmI
CmJFM0CXDYFtgmTBPZtxYGTtfzY89z0+FjCPNXaJW8pSjyK9mi/8XXLAiWcKZaa+
/ykGwK3uV6h28fkSefSHFH3VyhxtK3N20N6lsHuieDHvYWW3pDwZ9WL9/YnaHsJ6
/CXs87r2FDtIOJWC4QbFqulT/INJK0iYts76F9EEf8OIGMoX6Vdk5xJIXxLnT4jI
YGVX0R5MHd7YB/xsQR/C6ASAZ7RhI5dUT92rYbJvNNKmxD9qG2+/F0iX10LaVOtM
1tXsV7CeTN86Yh4tkH2KnfyAUicSJqwZt+FA/641ixCnlrGfR0u4Z40AFkjufRj+
2n9HWvWeF/314TSIvlXLYCV95ppM6SwDpfGcmWS6PSzUElvS5EpcrG4PeXsfCY4M
5kK6rYmZI0aHHvtm7uwPTczEAsovMXj4aT49DlhNWtBqQshCWMkUmuUcYyIdrvus
tZzXgZoU25FAdajvOw+rT3psEl3VcQmxNLE18y6qY8p/YYfnb+i3/vNB4YdseM3r
ulDrcxfypDPDiwXtv9IUj1ysGR2BU3qTbCF0CjW0WO1T+c/pd2m9YIbXpgdAn10j
QScRb8w9/N+Bwdg9oW7zdu7E3iHKuHkUDLPGkrNzSVLaHe3HfFjccUQNmXT8lp4h
+vVOeUSCQe+/GyY8VnLS6pFxKoGR2+4o6rkOK98j+TfYbAeAwYQDRQg/Uvb/XPYq
WJT8oeGcJZztjNGKSeB82VqcJ0xZHdisGGRIcQ1sC/RpLNneTi/A7hIicZPw7prD
50kn0t7X8OA17okd6u5ujr2iXD84tYB5k4UX9seCf8d6TIBWNYjaFA3HCY3YUo4v
x21BdHYQOz0arqL+10KfslGmeH1IKVC2wp8nRa1aARv6TIG6kGRmnYYOojbH55TK
ShBwWxPWX5nIKpQakrprGnb1gWTLscGocf+fPd0Yi4rf97lGzQbC0mRQMgHQdFtO
pLyawK83nTBxWdEjyu1mcc3khzMXPC/1ZrWrOqVImx4WR3K8WsKKs4JEkRQOpboD
HP1znmYE8aRn7Mj2b4PK64UqXATfinAZ2M2gLTq24kYQByd/r8Hqtoq8hinMlryf
+Oh7ozHR2XvRr8JeTsMakfKU8PjCbD/hF/WHUr0wnzHsK8uepLQjWfmtqff0hpDq
QiE8M3qHLvVQJvOCrgb0CFFriFIsgkWN0FHaLvQv1TvCw2TRuVPPKGo9AVNR+MJe
JV2z10h8vrKmnZd9FM8sRf18AQjmnvXaNvtsz5ptLrz0B1HejxetFrnF82oi03FJ
sFd/XqKFQ3RRzW2XcHJDiyCnai6t4A6SXmKCdq3odQfzyDuiqlZNuqWCo/+i/JRb
dNESsaGIhPnVmk1UxJFGYvRV6YsQSMbc07tnRdbju/lrj6wbeI89IEI6n9jn283T
4YphUhg3VV7EbcHrjg0qESkhduH2J2lz8122N5HPJLWdeKCs3tcHulcffgZls3L3
ePQNJtn6U9xpM6v2xYsHvzitFIFkMQnjA8nGg2vedtpIkVps/9l7wMV9GbrP6Zyz
GPW1lpGz0bJwq6hiFwlY2yf2bzuQVMVGVZSVKkPDQW0KnzNEUUhkiWXbtgmZcpYU
41El70y8pKdUlJz2GeolFze/0BqbBoX1EJPX7T4uSxqLnDad72TYDbJfsNI5OPkN
b06kOU7WNT1d8fVLQ9ZiFbtdLUm3P5iY/5qht4P+r5zI3mIducwBgg1YmBWl4Nsx
KpOnq63HPRsiugA+8Gfg+C8DgymDAPfhAHnXg8MMPCoR3GKunTqVzaw71FlPHv15
yYTijlZJPKL3NY3zCrDse7F4hh4UP8diQizsFLGP52Bc1rnMGthkFlXdX6Rqfpni
RCH3vHiP/cG6AeMRDodnqplyhgZLbYoijJWSnS6AAWm8QDKdw4lZsJi2SOqbTAow
AQMYHedX/iDkVeYauEVmLZ9PSDKjl/4OP1fYBHjIJOdYCJOasgjGXyzVusq7E+QD
usSEnlp18bohrZg3pVSlPHSSI08Cg6koARxyhYnf+0jN0o/1ZwEEcTtaZBdf1Hiu
sqVPjoideWq7xFp/rmBzoa/leGvNYVjJobJG98piu8uNbZK4EPqQgijQS8AumRf3
LRJq30Zcmlne5mCc2ayh+Cny4mr5gilpLGvWqpTVdiqbZTgGBYoX2wRGvsU/pXpt
Bb0RzAnLAX6AjGnl3gAysSNGbkAzRt1Jkr2MlGA9mnihCcMczyOcqiRTBy4iCJsL
xnqTqYXyfTzc6u+mlhEiEoI2JGoksfNU+/RA9FLRnqfd3TEg3+S/k6srRU00Sln2
yzrHEX/fuHK5h6n8OPGgZDSvdtT2+2t2LOZmV5tw4pEtzqdjQJrpQjwL2ctemYeS
VWwBguFCJ7ygpk9bsNvDdHB9xnPyx3AocMulip9mkrj6dcdwoivZ4+65yeQs/ZJs
RY3kuiUwhhgfAQlG+skmPug6YNG6peoFf1b+n/a3Dwi/rEVfml9/PgKxK3uZIlPD
1Zeu+GYpARjCazCKDwwOYKgmxl09wFjgHUV0Ai6pQm9d3+vAoJtjcS0GxWypQSr3
r2olfJUhIRHqKCNplrcwPQf6goS8yOz+sNtioj25etXWy1gBF8yp3ps7AFVUMDb2
L6Oh0dGYXkUmsOSiCxE7Y6Tyv7/4357QYy1+5AXNWl479pz2FmrLCY12uXorWeeU
kNSVp7zXLV80z+J8Co8iy75UvYpPDQqbI69RguT+vVaP3gtyFJ7yslTbm4HdJcuS
50dA6RoqOcCDex7pJEWj+hHouHu+Db2G91ILbnnb+ubFxHj3A9hiLng7wKB/PUE9
MGseOJpjIWT/THb4ELT8UYjAlJbbnMjK9gbcC5LgVTi8yjI8W6xK2aDanZDwyRe6
cy6DWKWaEQGKNtcbJacLmGizg/A3iATY+gHgYbNJ2hOzBm4ykxpWsQUZPgyjg5Uq
qCbrBCX1+pmKKYb6ON3gGCl7SL3P3FouTFIiwWoxlBKprJwGyd/ddXE5rSMlGuVs
k6+n5zCh82I0C+EKkMf+rWVU/0LmS52u+xyQvlJ5K3YNrFVS9rfKzfZmNzR3W7Fq
XuWx8tCIEyIWayxmoq8vrOS+g7B+48cAUR5ssRVd1cBWQhj381tMxJIoIz7riF8V
OHbB//GkIAEjghG8e49uQqcjrRigt/p2hYGzTU/onuwfUxxTuFFRXwhrPx+HBbwP
eYSDwdfaC37Bl6xVkMYiJbXZt/ehR2T/IsC0fFxxM0+JqFtMYVLvRk9ADAlAybdo
Vp9S+1Nrla60G68kzHGYiCnHCNsH4UeN1UNeIHkPW312VSy4fmZ6YJgIy8LgFeTt
3Vc7bICNL5X6IsC0+q5C8G+vqLo4mAy+WgPsKCXj20rCz9Vix5hQV7d1Qbg3WBBN
if9OPtMxWxp53fYvZMmFSwPttoCQGecONBdtfs3aPsv0azmQ/TE8K2RH4WxgKQEP
N1RijkuQqiCqVvofvt7bJuCqu1mGdJgvCy+SUPJ7WZGkFHAXK+I+tyQ3cVr3KZaw
drTXBDg3+5Q8ETF378WmBJhbu8mxz0iWZy0FDEqmL5wGW+2jRvo16LJbXbaeWVw9
t6Gd7XMt0K06g/oOp+DczjNnebNq8Ru0x7c9AXManhlUswSRwnbAy8H9iPDd9ikA
mjWjKF+qkboxeOQW788fcHe3FRbnCA2DwVxXSdppGxY5RVQrDFYbbpTpUnCmwQWq
XjTtvFQt7e+gERdgvNw+1G1uR11Lba6u1V+2ugLnazrSwz5u5IIxms9dc90Sax6b
0dHMyqrgu4FbrLrJQFFkVrjgWWAidQHilZzrWDFBYiwv1gMJcExohR/UWFF2rPwS
ix3SaAqKD3raWdsaTCU95DWlGtydK00YTFbwGiFvK//+ajvQYeJ6bAKFHE1VYlVV
lx5wR+yxOB2pYHo2PNZIAOZSLGjbRoTA1Q94dEYcnMU0VTqIrpZSp2pX2gs5ds5T
aXSlrCu412QzItvDM6gjBFeww7Wj/N5VqhCogXUZ62T30QlUl+zATfb8NN0KCib2
10KTD913miyHW1ez9Dnhd2x+3jCgiCiYSSv2m2b2L0LQUY2VEgbXhKSGYWcW1hT8
0lS5id9/WiFUNif/Egrj0DGJ/jYV4jnB7tw+WlXYYlm+a18sM6ddBIILIPZ/txyC
GlGxV9h4CAMndszKqVPCX5lhpgmpHggpA8JOR/QpDiLzEuGUvfBBpaPS5YEy8ZWM
zgVmzjQTC54PAiTTsB2f6Rn5KZ82/oHcSwxjjIv/uRIkizea8A6lmLzbuOnW7v4S
KC3rGBBBurUiijPILNHn1f8R0oz/Ip+y7eLfir70R989yHsDy8RlnWXilm2ry0M5
LXpEKj7oE6JLzBXO9RIu4XU9PkNWDk2uw1HI4FV2m8IcuNTRVlz99rdEDXOMTyX+
AHQ8k8YZkRS8lfSCwL7/SL4mkw7YfRD34hNvAphFdZt81OB8cP9k/f6Al/8Zyeev
6IZoIJBiivpW+5L5MwmPv3Brh/0suk+5TA2Yeo1dPYYs3w2SD5m5dsXqiS6OLcmH
ZXSFIzqXW3ZFQCsqX7bTGNm17RfbQF32BZYF1CnAvbeQsWDTCKpv2yxy9pbjaxGn
j6ctfoBOppjrHAkV47L/Sfw//X9+SpJWNIdjY1kkXcIkORABUwlR4FW6gSM8kqrd
gclTZeKmMnaQxm+3MvAJ5hU7ZQXdF+05ykSdzJhC+zMLTXcFsgz8G4akElII2vaa
9oL2mGOJTKXimbAIat7+R8c5cAmjvi/3ntOrN1/fObi4FErKUc2l3v4ClXmkyqDp
Dvo16hS66dUfzfk6Z9iAsAXPg9mxRTrxmAUdy38V8xHrjLQyXC+1CAlGZwzDulX8
xBMudq8LxuWHfwM0RtqHEl5y13LedhB2yAG75Uyl+zOICEDnwCtFfMpi2S1K6BVN
usNfdIG8ejJYpC29Gwz3jVsAqIPCU0CbA2weAfnHOMXKP2q3unCM+SkN8F9ud2dV
sZxbsTYLBcm8a63uYW6iWuSA8Ypp2owDfUueqUp+5m+mu35EMviNuZTskuZ8Eg5X
o0YIGD3i8B8jjvInpP9YnflWv1CJQNJ8YFhvo+rhlcb80Z3NDQvdIKk/QLNbeNRa
AOyhf85suLDb/cx3V7zXYX28NBJz+K9ZJ3oWWxB74wKBVfkZrRNk/60avLMDHUKC
1qPnOtUQgkKjgVZIOZCUwsOmoemZNOLa0Yy/MTV9umeBHzzA10jVw1KGT5Vu1q9y
3eFczWZCnUvZeJZ3onhIURJqe+xeU0pQ/ItTFA48vSnLuTNQ9t6bEr8ltjmiu9CJ
jrSQOh/9yN04RJL4oZSdJ9PGGYxfV1252B44YjFnsuKW04DqXQogIAuw2tWfAIrJ
JCewe0vgGHAwCIKBtPZ+PTHDNAm+8ML4S5T+GdPMCiHzIvPqdoORNoxLLHm9d4C4
f1wfxEQnVNY/DYJy3jlCcVdTh0S2YzCy2j1hSA0P44psIbVVphuhbrYF088FXuHA
QYfTO7v93jS3NGMxBl1AFzatI+/inB3e8+EwfooJQbswAW1akCrbXNljrDXryRXP
mRjk79L0DVVyfCrctYSllVhRwazKTkZF9wdauvqwWKpefj+Z2bHrC0eRLP3nHQWo
XcTSy6qmxPQR43Fxa1bpzItZEjmDebc2loZOsUtPgyDMKRkA+0DMXSdw8ArlPTQq
YCRULhDGC2b2QUU4dxa3UFNXnAlnwBtsH78LRkaoQ5+pmTdPigzV5++QgCOFTRpx
eRNbAoLnbfClU0kpBwcw6LTCZm9kIWNI8EQ/hPugqxWdTqAgyz/aGdAr3sGYKY+H
9L5EFr4s/IzgzrAp0P4Y1gSKrNlCvkNpulkAhUYMi4+f9kj+dpDs+ixQrc4S2Lt8
KR0ztMEzBmtE3NO3do4Thf/cBktyjTZtpUO04dJXi3IGjyOEy4s5wmB2Xpy73rPF
aVmTRy3XlohY3o7qCpIZ5w0ixiXs+RfXpphlsNB1CNNGDCRzMnPshQepoPOC42WS
1IVono7RhLFzwLninzU5xEV5wRiulAIaJe/MEy7m0qjtWQx/8IuDmFT2evIRd5nv
QjI5c0+7wkatTaKPVGR2POyvZPEBRIhGEul7Obv+GWLmBZDwL419ffA9iS9HXlsE
fcKdRwBd97cy4RyKVtaY1sqd716B9BdmHqior/0u4fYMzGPGXmhej1IGhDdYKBCx
vHA3QOUzz+qskD2kAH1FRn/KkU7kKR8le8Ej7X24q/GGiF24vB701SzsI4CQRE/V
KsnQcuYoiVxrVAxstu9qm+CC2ouvP7FrFdYn0Vlwsqq9NQyBRX8Z+MzFmN8ZAV/J
FfiQ19uW5tuMvB5H5zmy5CF2qlMtn4tw6fuZ0D5419ZgeMbVJqO9/S7MhhF8RFA9
4e3c14WyL3VDFeDt9MxlX0P2EacHK273ZO9UP72R6fsvXKuQ8zxTT/S9Kro/Qiwm
9lVXtZlQn1x0n6TotLP1uvn1CBr/QoP2YQW1jJ+dJVr6MjmaBpc8+7WpRX97ezy9
Ak+LJAhbsjUPPXaE4vqd/FyBAfi1Lld21N5ETOsyDV16qeXa02mu/h/kNngyfI1G
yke3oT3d8s98vDv2jBp/MhUE4l0ASYu8iH3+AE19uMXXvNeOpe11sMoRHWVUtExL
MvH/Upoo+fjNlrbVU95SQzudenb1x3WrxfEsZo6URcKM0baC7U2HF4Zqv9ZtNKPD
gsVsT5GqO122oKQz3RaS8UOYDfuLNz8URJNvyzfbzG/6t/FJ0z2IkhcevNehdZEP
yPpbv3NpkFx3H6pi0J+epAjhlSlc0p1wK1gRarMd1sJChFfp7chnkvRg+Cm63ybW
vz/K69h23MkeAANrDVmaa2wkblw0omRHumomPjMe4IflWJrRxww+Y0m6+Dzcjied
rdjOvq/2r16W2PWiLs9J0QoMYgK/rg1hy+V3k514zw9ewz8bWMc3NwSaVN8ae5wi
kMQBs5J+hiDOr29uEEDGfKremx7t6+4p3xZUoWG9GT6Gc9VRZqCdYfhCQ8HVP6EO
da9lq+kyb/wVnhiAuK1b91mCvam8fUogvImPtaI6hHQWBd/yFKIaz4Ua+TcWk8iD
4PzxbgeY82+Y70PR8hlamwnllMBRmarv3uMhXmJ5eVPzf65QK/ANeuF0IqrBC4o5
rIOyJsJWbXHoZLdUA0Nj9fPtcsT2G77tJjkUgLJPfsAtpxgP4CsX/WOutQX13Wno
6JUekLREbPFZwLXZlE3oqKuJJU80/fyvKjOUoBWG1aYmyISefryVulzFX4AR18M9
gmQS8pXbQkRTNRodLvylx5hINC7pbSEx1OIchGD1zj/eNMU1dpHzER73C4vvpBIx
EgB394IlMpszycE75FnTpvkvoLzYAu8EfXaKInoPsbFNhU5C9J/jRfTnjw3Wnrnp
4os+3lxeKCTygq1GHcTlBQ26OPVudUSY172+LYDceuqv8fMLOYYBNnF8wVgdJXnw
sFWlI9KpVe4IfRZzYHng6jqSr+2RmqVrWsOnyCDro6jA70FEJPnzOT4b2Fl2sw9M
P0k+Iy3n3Pb/f/nABTGwF0tbupDqEZzu29XI3wRkiul16u+Ldz44OONu6IE9Bk2B
3e/hTMbSfsEnSoGFYIBn5c8lNeqwKs3TwZZBXUXJnMC/4CtmllE//hiL6xddL0tR
UNDFS4/IyB+Ir+uGjngQB/prdaRfo+p2jT0whLl/CiqQjVFFl2u69NEp6u6avmO7
HqOESPK2/kowJsUxvHjj6b5wo6zujry2iOMm38RAl1N/FouMfzzncZxKhpG+RUQv
I36wjPn21JwbB651yD+WzJeSarrQPK+PLPsFYX0oDSOQR0f9t+A9VPUbSZhiDT+U
bklWandLKnRtEVTmhxhJWjndsvaxcHKHFTmeAd2xfBLIF700rIG3ZkODakFMZtL9
CxsGG76ZWBBxYsBBp03ym66zEXvSBQLcbhTC2pdqhDENY2KYptmPQV0QOsI5GpK5
mwa+M3LWJxHYp+gnARfqfeSFOltu+VhYQ5Rv93DwQ7nRT/ZrZbxtuyJm/DtL06gG
6v44O+qMvln6WD5jCfJM7lknAPYu975ktsBFhy8GHm93hNmQjveXZFeza9ypNdcB
94DjvXxi60FzkutTkzDsLnRzbxwMTuMYMJvvHtKr2UYydPcErb2TR175erttnxyc
wFsqenOWLkUx6bNGnvTMc14GlLXUqo7DUicwHQwfc39NfKocNOw5scdHJcMNQ7dE
IDyqNZMKsz6wChOAYJSx0givtQNG7QVmXnvN3AT+xPAFNLMTM1GsxpGNsnADzLon
2cEauNO8klDW9ZYJ+nhZmQvS4g9e0EyEyFYmt9TYy0i8CAhyE0pm5CBFlfZxokER
DjquDwib8x91TKdxtSEt57vFPzUDbcNpBa8ExdJhx7/HJ9CAzPzb70DzK6IeYwrD
yaWBg5cl1dizVHX/hTN6tNGkRElQuHGqu8YI5DguFjjFcrQIqm4oCuayRJHExDqy
tUeobivj6Mgi5imj9tEv/W19LD81mkI2BdKhzs0/WVB/JyWK2oBtxgXr3hE3Wbq7
0FKz7GoXPbxjQi51ZnwIUQ9uqDLAyntefjQx1cEQcRxg66m+cypsqRKx8YaUdY/u
SI3Nv9Sj0wJheVdnIpLtk4DDCRi0s3w4lxSOXfl2lyUFhENmj0OMwMfg/IJuM/6C
9ennustAvkqjDLdz0EswfBj5FIdPPJQTUjlIO4qU7q0bjlEW/YfbkFr7Dlg4rKOv
b37iIQgTE+iIkUN84Vq+Rrh+6GI/VQstmAGnAJJeJOQXeVw7dsVKCzC6vlfEdRKe
ovNDMAYI+VDvndQrZ3cWKUi/Bo63njVwj3oq0p+Wnuiw0pBtPvxT5g3HFdBmofI+
nrBY7SErNBsOV5QTbfISmFPqF/ESnqNZHS840m0L1OZvx/GCIjfLvFVeWC3mkMYF
d6pr+M6veInACdjBWVvBU8kb+LsjLA9PclVzUfjb5pmCLm3uxbUt+Sn62Hl0E868
D4zNM2/hLC00YkBxVJdq6+k7ojrY8d27luQBD+BcSBSja3d6nkSiNX1KcFUp4m0W
Qa87OUTGYq/1Sml9CHj1rU9o9JC58DzRE9jiBgfBRkrV487W+Vbo9N5vBlCNe3s2
pIGdY7iF9ecDGY/Hg8RCy1ntK2FQzzZt6QpFnctd1FzxiuGZUb5rDTDGIZfLs4rN
YE+ycXohScAuoVp15TJiuJBDm9K/n+7sK1EXRQMN/t8Ph29IM5xiHNTT1jAhSn+f
UvjiFRKpwdNDGQPZWO9KFylTy/Q5LB5ZDDDYothW0c/jJWft/lUYuckbn8Gb3Z1a
PmSL7Wm59u1vaYGxNyzaUwQllLA9loRwIDqU5byL44+GYRfPj5kzZUj4AwuGVu/N
mEzIv0lyMxlA/aEc7rlAbCVhVF8/BvptZghYs/eLlDkIyJFZRtLVKr9YTqIR6np2
7qMjglH0idW1asir/t3SnIduOV4qFT+xRQQ8PWA5ehDFfViZryN4RnJZzjFs+qA4
QfJu6sLjHClyUa4S6SRnIxIYsoVutlaBNSsVB13Brd2eIlXvdeVUsC/6BJZZXOVw
l/YEy6VwFxPIEIguKstpnBnPyfZ3B1CktM5OFfMg3wSFTtLMP8PPdsWjl89rLTxl
+4Tiw0CeBtkT0NB3o8JjDJhGVCZX6rvE31lvo6lmZFoHDy1zoloW0RPaSMPYaYHt
Qz6M4SduN0Tg3Eu3ug8p/RT4osZpfxu5MPGLd2CAohFKC789IZn/N1INFbSXMgBa
NnJOB/cm4ZGdJZskHOkjBPzabALr/TXZPgnDvC1f6HfgG6uCIIpnb8HaSEuKKpwW
8GVbT99dDQrhYVz9zwxQwFJX6b4mFXGdT+ZT5ndWdpF9szZ4v3PESEoqPWDEY73D
Ni+qjENhsjFUwEJjDVG3qEih4rdz5EO38nsI+YuP74FlBfp06mNJrmzGW32eiE+Y
lsTg9FtgqAAgYOzVHlRYrB9cgKMOs0dpaPlrni3X6vevigmiwSOVAK83B4N9LRuG
8ruf1kI0bNbl2K6ORhqEoyH8HGnN2AyWdZxMtSasQA7y3NF0bWJtOKZZTg8RWWzA
tbUOYfyXmuVKpfVzjjkuoTjfHpy40bprwttwFiua3EZy1tpQOm0++M0DPwaNIMmt
MzWoSgOHNbZwTn12q7/abxDPCgUAVtGmudPpFhulsrLZeXLblYOlHn5C6GZ6J26a
1x/FXReIi+KVBwUSsLGb8EIRE9l+RNzNuTBrR1vFf02zakKna2RXkGGJ2ScQYwFw
3I5txjLFqvAS5xyB2+BSefmDTtzPaYHEOhETYL0IaBuD9lDBa805ku2RphxdoZSu
jjtma9x1Il9OfPK22bPYmqdadQbHrQ1SUuH/QuSPt+9+lSQLz9puaY1A8w8Mf7X6
EIJskmj3kxWnw69Z1ftAhyiq8RgiEs2ZXEttK9k/OAje1iXbyBAUdc3bklls0VcN
K0Q1hRSp75Hu8uzj4i8o7K1M9LmgGM/vTa6BgJ0er1Ytd2Gia3qVJQeRCUGJa+pJ
TKgZ8gL9WkMLu9mzt2CrotySDxR/YCoLBCpe8bihZ7s6dNFEOGCRL26nEHmAINEJ
O61MMFvxP3KiouC8NYBWi2vD7otK5U+ssT5bPPwIvozLntY9QPrqjV/SY1UFIYYZ
OKK/zPxyn47XPWmaI02SCdm+gFke7vpd+sGk6+L2enIBqvMzCVtQKQq1IIZbyB1t
naLPpbMl5HD+nNTrlSVRBFy7qnhhDe+yvV3wRkuNhf1X+prjZ+7T2Wuup/qsa3zp
II1KNc0yY9kiUrL75AnIXgVlIAdUx1q0bN1oybrYmMl4Oh3CAuF9hiT+cS1WNLoD
ETcGF71IIXWim41+EXbSD32ECHr7X6ArDRSm7eusBK7k/vzDkTzn9FhQk2rux6Ib
OGcZMtJ2KJRII5N14P0JqsOM4Z8+QDIgMLBtHuKp/R2jcorUuAZkJkTYijhEiTYr
+UkjE/Y4DIwYe+rmixMVwfiIP+GMlZosG84kRnOXIwEahefBtsec8nmYb03oAQKx
AwNLLh9uI+HB0YvcMtEdyLYQingYgw/oXj44HSB0VdqgOxMnrbmhqpjpt9+AQiBl
O6Dr3k57AnDDFJ5AH624XeFtKLJ3QpUZqMhzJvNi5SrJBHahg+FN649+c81dT98i
d3SWTJN2eskTg/ZwA3qpAM/NwJA805aA7vK4OeVviHdK6M+3p51yt8EWuZR+1RJu
WTB75PN9vHDVIudYjKaukYoWRJnM4hDw32080emEBNzcBvrJO2o8AlKYND4db7rv
L7yjkEiNTA7/rBJeaPNTVKY/9D4NqmhIciL4M3AkyrdJKFwDM1At3m2k/7Bsf/P1
3XpaN1ueMlVZYLuesMuTWzpWuNg+rjd9Zry/0cf5pjnxD+OZ+V+sGqZYbaTe8M3k
Rr6d60LKHdhAV6uMjqGXDHH8H+HjcaOsRv5ZjsNeGzVBlZp7oMWiKN6NCAveBFCC
ZrmVLiWMq/82UOFg57IFcECFnIFDISWm49uhHi60/9MJJbc+ILXzdmdMnmPxbJn2
BfElbaqcVnK2E5REIZtml8fLXFh6mwMSpTp0tKpt+19qF7BXE/zgVTxuPc2DTPpF
iI31b+q2NGbcFeZYzC8N/EWNyGUI2wSyNYuFu85KZk+SZUqu0tKUWs/+41pGfEZe
WzmLaqrXZd9mr97Fk0LhozS71DVo61qlqiYLMx+rbkGzfEq2+aRKHfQryKo1G/+o
t/d/2LKIrjjy1DUQ1dmYdpnZjwm5uTlxW5ycG3JRk/6kEiKwS4PFUDuUqnxMeJtb
t2bB86ttMf4DBnhubW0jheDqFuz68sCOaoW7Zdw+1zkpr1TGG2a8zT/AE6XW/RrY
halnBrV2ryf0lPdRm1rnglrxOaeB7GRofJxMERaBvlJIaQzpnLIkj8BU7u8ZlVJ3
871IUOiz137fYbB0je6bpPHj2jsTas6VivseHFpRWckWbWf+VqmUKXJD6ZgeFpFi
pbpTtHy5IJfAPZ4BmCYGc+2NsY2dzFTnjwILRA1AWsqinSElx/Yv0No6FSmo+JQK
yweXPygiAIcNcKRDrT59DKT9BpBeMCrEwy3m9/12M1+H9sMNt3qgmClQYCywLKfH
+hkb6ninbcL3XTkey+w9eFJZp3h0iDZ1t/TGfdJRJE9uQ8TROfA9DnAgEF07a446
mRlSON0ql54vsXw/MC/ThQj10vddrxNDDqo0HMUfKtadWBOvkK4M4d9mZ9EJL4pC
iI8w3BX/AMcwMDvoMxZVt4jrGXLHSJiZhExI2omDyFcf7TcF1fiLOvVcOgfkhapq
VTv9agaWS9vHsDhtQZ3sXOZ0+AsK6ljRTwt1VU6hqz8gp4bzbzcKBV/93QmWcAov
drntgz9mvzVNG2ZINeU1Ntvt4wKd7gqupv2BKiobLtWqwaY07bsLYdDiUVTWSH9z
rXvImNj8UJQcH9w+/d3Skdr6MgeCc1e/VzDoy7zGRvVufGg3WZfF+I4idY9WBZKe
k4zJ1BrLMEidVfQnjO+WZhlcxjBV4dcbWYma8HuNKBbEJYKSUPDyXw7lXfNh+aD2
D9g9gA3X2OpIW6uo72AGbZkJkrVOstzGwTWr3xXpyuZmhC8m1GZbS2hbjUQLu/t6
sFA2BVIj2Vup3uW6ugE7XrHWaYywRnRGCnHCuzfE60bRAgLku/SeA08UnPodBu8e
jF0AqdhjhFlXFQaBhD2zHHm1AXqLm3f2ZeBx/0DSNc/wx62YImaWxXdc0+ZTmKsN
hEvD/Q61kdY5Qne1vC7Q2qjBkjJ9lu1x30rBXIVyoF0=
`protect END_PROTECTED
