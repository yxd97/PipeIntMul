`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+FAZ0X3AA5jhjkNxsFDVAAF2vAU/ldpWZIVWiA3ak2h6pKZe2r3Eoq67rkGa+qpS
olaW8H5QOdUQbUiEyJT8kxcd70pK8TT0IVnvzp5oJoVDN8QgpCFApU3cwmlMZ186
B7lU4dJm2s9U3NHy6d9VjFw+3rWSelvYZSC/oPSjCv/UMDqr7Kar3CznsBHJFG37
OeXXBqQoGUYEL7Wv/tcLnLORyg50IQn6UVWEiWqEepgIW0ZwaJFab+iWPixFaneH
`protect END_PROTECTED
