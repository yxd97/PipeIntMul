`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cr8jaRKhOYBtmFFju9wfwAcz84LZCAnaPqitsdpBgmfNxh5pS7JFTI7cId4UzCKn
xUGj6uTF/UrZ87hH20tYrKoOimPrGEl3vVkSZcOR04sdm92kUqfQmMUogkzhr7aH
TICrVOauuylrCqjA2Pt3veHlBQCceDF/TsI7lzOXsQGT0ayryyxAhBrm/umZYAKh
s/6GA5Z6moNl0+u5UGfyOk/cbtI6ayVtsQGg5OnpEEvieUgDzG71PRe9QZeRfcyt
njLLKEXdsRskflyBJFO/s50q9WaWLpiOtJSl+7Qe5GjI4dnr5wMDH98HSUUmbvGa
UZcPcCI3oFPDRbTX4JA1ayRKT6hEEFYvZAUz9QwCnNyskhrkjx8Ha0p703qwf2m7
eA59HLX6lkUUfmCtknPooA==
`protect END_PROTECTED
