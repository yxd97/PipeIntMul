`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+W77IOFeK95RKGxQr3xXpp8qiv05ztJ2iSZKY8ZbP0tDfJAiLBJG11jSliSIe3xm
Dn7GT9aO7xwxJEF6QZJfrm5xucGB0JuvshSwTTlk3xAOCLOiiUTjZzN5Ouce1z6s
DDlvMZLRSBAUqm6f1NjLF939LiPckRIjp2CTmwwQV1ExOmWPgpRKJFZimASxdhpD
w1qcmgwfALlgY42+KTTM/3dlTySsWURxGDps9pPv4HcisBNsHkGpYF2ZrsKQd828
a2BifMgMlKCY4p91/zMhZW0q8ov21Hl4fW3T32BYsWxzH7QYYWMR+oma/pPiv+Ep
l5OTw9z2nmX7PIoQ5hGk3vvG/iTw3/NPsT6M6I8+Jm5eWlx9LgviycbYJF1LrEzP
xodQxinxUyeZ8yDVnfdAC88aQlVjElLtlcBmfJ4D7PMdfjTEQUoyDCZng+hWAA6X
23dFDXLkBF6Ba3cBL8RaGbME8b4gxNvWNrrLHF09E9B93O13rqPri5zPYLTRTQoT
xsfYsIulJ2eXCgLEYKhDRduVQhqSfyxZgGjSNENWAg4/8eOBnUyAQboiaJ+eOJUD
k4Vz5l9rwOWROR/HUL/K8d+7psph1Ua0kYNLqsg614bHePWKgYcFbAQY03zoM6J2
1gNezSJN34rkQw7DRUnYMpy4bljXltv6isna3PALKzpR2verbgZQxUEtzpT1Q0uU
ZOgsGrAB2b9tlrB9YRFRi0TDuTF9ne3dkpmZ4VFk5qXHELnLu1ZbVfmH9GXMDMBk
p8WdkuFl1Zo47zkXaMPEeEAJpCZ3jpoTtOVIX2RrVnqf7cA/bNnaSjJSdFfZnfEk
uIO/wtNZwFlc+dgTe7CfkRf5gxGz7/wdEtK6DGxuN9wvljG9h4/YElvrUyVZCikm
jGHdlzos6PRaI6lgwKYeLojXDf2wDQEEYBs9PheKWsXMc/WS+FtAO1GkI92bCanH
JEsCB9aEJM36i3TeVTH3C/CfURgC+LFmWrjjVRUBEJfjlWwPYB1SJH0Ts5j7k9Ik
BXOauKcFjjc7V+FphVxPDYom9lJZU2XOFwtFXLkovZlr1WDKxFaFHiQK4TfV5I21
V1oP2G0oSkGJWRGhzdZnlDYS8dAUFBfy/OCzTJx09lK7muooJlfvqbdbLjwKQQIN
33Lpx5cA/+iOkXjVxr9IiTqpwGWHDWM/Geh6uLkyXHcYNoU1JpYl+hVryduLdZWY
QDuKb8tQaC7VO9Qq3Q+obhs2tNnIHjcVcMpcAg1SwpbnChQz73vMlipnDmt2G1aH
hujtMWW5L1q3AcxAeLa7c5xO54mtFnPlzjDup+YaslD/dRZ3NQ/wb+LT4RaT7Xyk
Rma0QXVMnIU8J1II/gsLsQ==
`protect END_PROTECTED
