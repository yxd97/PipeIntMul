`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cIZ3O7MV5rwYuX216SNUmleUA5uljVTzUY2iYkVrJ62jHN0zd1NuG8ZAA0kYkNX9
kt6KgFc4cw2GyRE8VzETDLRpf4xlaRr16TctwCW7dvEs3NvSa2dk6Unb/e/k3biH
jRCjSvx6HolSqWOOiuxVjvPGwFpeNVMX9hLOuve4rVrlvYfjJTUiMENRaqsgAVNg
Zv6B+jbgZhglAXdB9s1NNUI7kxxOwwQBeO4Lc/d1SvgxhhSKk8mrlE8CLg1gS3ZO
8Gs1CDSKVIegVKinTxIBbw==
`protect END_PROTECTED
