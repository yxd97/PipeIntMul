`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MInUnJTlf9LxZsybsdFRbVCj2d9nl3BABZRbmFqRZXebxdS9hsUnP7xBiMmn/lZu
sD1WoJJ3QzdCD9jTwzkjOPKnThOwKAGcw0+N/qLSI+cVUh/pmlb49mWSMKjKml+J
aS/qQbvH62PnvGdANwAhxy1BQNJbfBDD+AsQkGj0TiM/AxtLJazAQxo+tK+YTx9Y
zSFblQ4x0sw285v2BERckvShOstjstCBgt9BaqKtb+utbKVJc7ebPlima8o97NI9
xzh+fiQAyodq5ctsQemYLAddQWNOUeOKJXjmBYZ0l2uCpT86AlpcYDGrUknmlKfY
CQ97tKyIEhUmkI/ztdKeIRj0sbPy8EKnuuGEGirtkwj7G5/qjWjsto641aTqhWrv
oVGjVJ0ziAGQVPtaTmW5p6dB2Opvx4fQQJicBpKKydNW3Xn2Im6w+11+11Ib4u/l
yMjvh9cTsNTDOP+K96Um3r1iwlvD59re4ZQr6H40zY0pd2hwuGg0s53lY5MCaZx9
`protect END_PROTECTED
