`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YDBfY4xWxH5jEHRDRkR1cCHamP1K6M48I0eujHz9bjVCzN48E5TH8erkTqnO0Acr
iM2BSXTGxoHDOJoOtjiKItK5il8Ci6CcEEts7c7OvKshIGMXS9jMlRrSgVTWHxPE
wCyQFUJ87Mx4aS5u/6McD3+98NXNJbdRbcr+9bGj5RlKRegojEzf9GFusePbtgel
oWZ6E4xhJ3BREGFxkc9qwWgn/vfZh/jPDMO2nLQlCNTFD5Z3SwJ7YN+K12wMp99w
ocp7LigsrgeIOkOBlsTmvQQStXwNQS5H8gfPP5mh2Y9OqyIxp9/Tunb/vaJU+iql
kMCwCL4QHDGPgo8o19/RAup3Lrt8XZDlrVoF7NWaBT9hly6uRnk+Non/ICAPXrSW
`protect END_PROTECTED
