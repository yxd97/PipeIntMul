`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wGP3ePmm6iQjoOTbYYLYocCnlcEriM4ZP9wao2j54/NO7M/hXNZttrpgHFJ4/Wqi
JWiGtkhYp44Diix95/2g92ch+yhb64DxfEwx/gBr0qe9injceSMpu8vXwQvLM36S
WFiM+kt97WbU2mT7UsKJdYwE2G+h41Cvom2R7sNAPr2QzXrhhVP5F0OWr1vogMil
XXe+zb7Ys8kpzLSNugitTnqYHiT+AfUa+H3OGH6Af36D/6ORiawwNvtncL8iXjBV
tagNtg1404lFw1M4sc2QSAh7Cgo2Om7QftAbfHFW33N33VgL9D9VVPIgkXRPrZCu
Zw01QbAvKuLRNClgCWbmKUhvYkKrIhOfQVz7Da+krsQ=
`protect END_PROTECTED
