`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jje2z7VkLE9umSp6wQhtyMlLcVJozBGojAy5F3UnYuTmuqSiYtmmufc3bI7aViUB
cr7oPVAnYFIIhgkKjZpz6RWrSH71OsD30ckvQWCvfjyt+j7S+yJNALPKdjYgvcA1
xMifrRRIDF5K/64eACtyfcrxgFnrkxYx0UjXzgotKFwktWdpWh79YKm4imROsYyD
dr6+1xhqERHv/5x06Q++UPFUWD2/otbeFsOMidrGEP1wCX/kSa44JNWMZpt/Xl4M
KXZgOUpqhxV39i30o/+mPicrZRAjw9O2jirPjdVI5eWjF7ybljDoFUnuZZLz8h5J
zBmj0qNNKhtoTEt+OjZeBCJyrDaXl9sBKUcBaqs4CBIfHymsFpg8Rl6etmgwfRIQ
DNVBr7J3ZKSx3RWcFQO0JnaNWn6BQOEMvqScU2XJ35eov7zbM/2pJ6XVI2t2wHo2
Gqp/Vr1Jj/2HC36ukE4/GYoJdnpIM3IXFR3M5a8vzBUu71khNaMmWsec9Clq+izb
Qhki2rCeoCURRvVgM9reU7bTkAqn9JdqBhBthJuBoEQUj2fnLnBAb3XRFSk/8ds5
OKebGjYwgnGJYNDJyeu7q2r8zDvddjCAisajSRAhM1vwWeCVQd6dQG++/DmogrKT
N37r5HtpltZ7nM9CefVYkjiRCgTScCDY8RkcXS0V959rJQDFAMDPN+i8NmU0vl2f
wX0kDTQzXw2Wc+WpnLgTVtQzOosJux2oVkCx7m5gA5vZcqYxCu8baxJREfpGveCY
mFrgHAXiNLEWQa8owqh+mhprJ/N3l/Rji5q7MA9qA4droi6x9C56i4YKgqw++qZp
EgjOONg/F0ZzKDywLlVFLq9Fn8GbmfdInhyltrlhHfLBZBgz99snJNahqpetCF/j
6gxg+/mrI/YkOm4LS0Y8EOcyeJD8TN4LgGKkTnJWDQi7SheQ24m2j6VQjUyb8JMl
HaeXVPyR6BxOm75VDGBFvrXAbpNjFl6pmSw4yjrXXd12+SpJ9FFFnxmGfZYIsq5J
JDq8q26plI48eb+VB0A6+bFg4k0Dzfo01Wp3qCY5HeqE3vxw/FegSPmUmD6Y3/PU
AeS5SUJEVQ6anB/GHVUlyT2DBHPY+hve0vL0gHn4RpqnbMFVOESOnCfxtb8bUEMi
VNRL6d928n1HoyuV0wS92s5QQna/X8hiZyNYUsXtIx99vyf1YfjqQtLwHIqTuae1
ILvy5+DbTI1RqRwGmmc7f0h2fBIF8S/vTSgLvCv2QyuNcY2VwiCtP2d9hovZLFcu
AaogP0xW2qVriJVLwSCqagEYc+Zfwe9+xrFt/LscYzNbhJrq+9oe1qQC9f0oy7YX
mToeZFO5g4PVMs0XVAttuUdoaxuIosU2I1wF/ntmOVPfPutFC1GzoCPNutH8f39y
IjAo2RQoA4ysnqjinS7qxgPQHOZEJWGoMNbaoFS5yp3N5ogfScQoJtpaZSnsduKn
5FQQk+LJ8DMJLSX9gzbTFFHXuyIns21Zea3r/tJrzyxYvgjwLTRUZiVJjID+yeyo
sWUAIUYwR29ndEFsoetiatQrUBFMHkZsRDznZKEaC0wYTobAInpWocfdHddh61ia
z9SMfR/uFwr/ZlsGcJA6tEwKDWEP97iKSnWFwWnnI0qkpyymyS6uKenGZVuHG0/X
w1wWRWdTY2NIq7CtUKWDxxlE7u/J/WhjVFBnFV13jr9gU+tn7EE8PrYDpUTi+7f5
w7mE1Xz1YbUo7j393viqbfb+DsaECnnYMrj1W24eK7v8knskmenZfR733WXfxLJ9
JnI3xhMrGHnuMmTvX3ziUK4ib9jyBgwahJgj//hD2YlAKmRNAsd9WYeeqN120hXv
Qxhde0UURle4coQuX3DpR1/ufSGpJzlkXKYM3Vtj6tzKmbgRVjz4Br4iJtdJgZJP
0VPhehzyPZSh5ZCYB/t5sweVhlny8KjImQQan+bwiPHqxehNyrNNObOq4/89VYEm
vfg3hJcgw9WfEpepZcOG4A7Afql02RbA/ML5RDEU+IYscAQQZ4N9vkm5el8Atukz
+5FipVUvFa/O9fOrONpf441Oscy6XK90WJ5xGroELtHQcuEsCCRVdlP3XS8sBtc6
APK0HqYlTvjZcIXaIfJQLHpIJ6ZA+0VKlro4YRZXnAjzc0BvbB88ZF02TetEIR0o
Eb3xmgcVSg1KyKumw/kKG9cGH37q/uvKldRHo5mmLgiN5JzmGsRGOo0CNmHhG8HO
VYNlI1gWTqcKYC/TUycIrLxolNM2KkR6J5ORuABxxMWAmeCzSCY7yfSPhJ2w7pZe
b2765RDIbkJQ8nb6tCYoQQ==
`protect END_PROTECTED
