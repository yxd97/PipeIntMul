`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9K66ekwUEnT18pa8MoFfu0LXWruUTQGv4hV1hchl+T6GMzu5qAaQo5KtKakZF/nD
y+0Zey80FsXYJ+GabEWNYAe2v61GSuQKipPib0jj0gLzWf6SkbL3XPz9IHLi7m6q
3LitCHf8LMcn/Pqd4gtTJY52aVCcApa7tdLOaKdNa2UC7eycRC1VCyNgpT4olg5X
s57ddktq0eaPCYTlYUdpJcGJfuPlnZOcRzZc/vCcK2AAy/Hlnah7kCNAnFF7LU3H
E+Fpr/oXnZTnIyVO30a7BQ==
`protect END_PROTECTED
