`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KSn5cyj2qcjitBe+UowadeD7UBfn4v3+ax00363GvtXbUQwwcFb7EfWIgJD4wrdc
9NJtnoEVQsN1i2+STDP3qvf3FtXDyYC2U/155dz8MQ0p8n9soFPMtZSqdOWFfpKy
O+vy5Anh+fuYE/PIZBLN/wSeUC9GJQD1KogoptxkqGWh/aDfqVZcueV7o3FMFxNE
1x8MvEqaLIs5jDgGDUS7urMQNgDdQu6iS3xw+RPU1oBbHoXpkyhFNd/i5IZm1oph
kH5vk6prUPVOzYp7HkxGlEoUdPwjUhdgDoxdRcYkvyt048coLNmaHsjPDLZAVhPe
gxO3enPa4jLV9p5bJHxKS4Am2EMpAUZvTmawckLuRld0vvCJHHSvsqCCY9Z+t8vS
EBPcsxARJpWE4FutkUDs1gADtxpvwIjrOT+Is0MBUpLJm2qzciUEHqBbbLMJOdbK
FQ6oBg69Eu6aF2GiSZXqPwAtxzKUvdGkNQjcCQW1iTQAbyVqvgz3ZpMnFlfcu5cR
`protect END_PROTECTED
