`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRsl27ljTEUY1EaiPn6mNmgyc8zXcpCyQij18oAbTfhtzTBdfldPI3IGXzuw2hR/
KhZq/wA/orYLiUd5jEuCV71YJ/g1thGg1CzcLr5s4CwMuEcaJdyS1cbxuilyIDjg
HYAoKAEfj5PvJ637Lqw6ZmQqXNxNuvs9S1qFoNRhUBEHKel6H7Y72ofRviGaVmaN
c0h0dVXwDhe1GJQvIK/4CGGXI9yGwpCoOV0Ah9AuS4yPT0/CGxnl8EKuAw5kkPBg
VRQ1VweO+L6+mjmWOPCO+g==
`protect END_PROTECTED
