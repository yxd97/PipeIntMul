`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h72DXscGbAAVZranYXECj3hTHlrvRQ7FCCEZELmyYZihiOLgmRBDpQ2oAysbnPDH
yNqZa4oXb2RHC7fjh3JcM2pBa556T0Im3X5qAqLh7jKd7mnLirAsg9+Mx8bChkDj
swdkyeL+UFB3WWRT/+ZGzymLTYNNfPtDhI07ay19U7lJRbDuBAf4V18CVzaxJw8O
yG7M4lnyMsqUFznxViaulHvjK3Re3/+Teg52/BNrbHbwRuXiwSut7tobrE5dPmkV
NGlQqKTHsO4w1UKHjIYB8oBd4yg9OJQOT+k5cFUpkoE=
`protect END_PROTECTED
