`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LytOAKVawTS+cEYRe2aOECmRQLUVKv4bTctGC1LGntrUTNG0+D/lgWTJa32G70AV
YqFd4T11iSl3D2r4LxcMRPYFceREnZ8WCwojGBUZpe7hXFrpLl2AAo759cQCGh1L
lh+TBZF1NiZrO7grEgga3Czef3qgT/KLuPODF4tZ7jzie6i9YXOaMFW3pzjEDAwi
OaZxPMjLq0ui4DUizr3VwTjHH3D8s+LbhXSTWfKAVstHsrhWkFDmYHhV+nahmeZP
PtJ2dsO9vRrpPJdABKbyDO6aLS2jSJpKS3F6q+85+0JLmiYYwKCNBmF2Sy+PBrO3
ROQ4w60y8MCUV4nQq4I0L5O5kZvpnqGwxx2LALCJaeSHzzzz7tQyWnehoPlimjDd
FYNyQ6yunpUkk2WokJiHd85q+0Ecf1C27OWvFt/5wWs=
`protect END_PROTECTED
