`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzFepRJpg6OrZgm6jx+BLnk8DVoxJfWSlzs5tU0C16QqIzHohkQq5LZtykVKyqXN
+GQyaaELn0d8ER9/iY/4VoXO2On5spdq+ke14lAoT065S3oBtE+VlRLTFDqqumtO
kxxfcE/m9lH4PBUx6S+zfrsAC+K+2DVGQSd3ajCPdyCS2mAUxxV4f1jmT54RmkNk
Mg/DeaCst8ZkJaDRzP8qRzI1G/TmMPu2E21RM1zjU35M6CxQ2ofoHfgQLWJ5q/+D
iCuyBSgungrCAJ7Olq/KzV5IN57qoNlEeBiBQR5CZdUrZgn5JFwts/rSwd/QQlhm
XPJ6fTzg5PHrTvF5OVFor2OcIheNIUwu6lDet1REvnu9cd7LviwTQH/y/naRUqQ2
avFXDYDsi6DnBwNkpHlem9AitRcDTdGSxkN/iPJkyTHXVhOQkJoZ1+xNgKR9TKv+
zBe7B8m7ZmfOMKdyRrYg/o6OPNhQGE8K09UZcB6K3HmT4f5i03a5mFYN1zoJUTeo
`protect END_PROTECTED
