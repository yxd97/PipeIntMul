`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uhmgCvhTUi2cL8iPl6H8mJQOuvkiB0Hp0TQho6KmJ5BMbv4/ITOQxllc6WG2iH28
X9ozBnGMWMHs9uSmDQGoOgEo0YGFGbfSHXNXXTuxtD9QCl63pP5S0RHDlmltr6to
J7XCAbvly7TIg40x46BawhZf7PKBRlw2tQVg5dFPOMalUTKRRRcRNGmOglzrDrgl
xt877cb06A2E52sOJHTU3A4sDQHSqdt04J0P3A0Caa777reo8LI6KiY/CKfL1qdt
vuxlODF+EoBKKGL01Ynas5UTRYl/MzWwnCGi4u14gU5P8Ep5sw4gMOedDLqdo+xf
IeovhJuZCtORGUCigx0RRZDCF3rSIl4pKuQeUAmmRfzdqpFQ+drejhYmW+GJqCoy
9jNAD0FzOrwb1CiwntpAAANvY2T6HKlmp9RhL+BtnzLUbUfwggiwgoyq4f01kIcv
fM8trSf0FA3U4BTaUDHPSaBgyVaJoAJvmw+Zc0CAubFqZEr9M094nDOJhCF8AmKx
Ld4EyPJWwZ5NrPPM6muA+GO3Y+AQL1XvIvOUiHnuZ9Upy8B+KOy8xmVc5TeYO8mM
46yuEOGriQ9DWoSouv7gL7/jO4Q20DFH/c8/IqAg4zf1j0rG761WbZ555lS3T/0/
epPMOFmLWz8tbmQP7A4GlztPLedGN8uLqbyjXCHNcebWqPgrqdy0vaYmdw9IkM9X
IzHE+3ClITYyBdzSwWP31MWszv/Mem/aeGROcvJ/OZrbfIrOZncmJg7dHUMObP2M
7Uci31xjM2VDXeQFv0SjRsv7ZPRVh/kromiU3i8nsDieuxelZHQoUK3cljhsWGOj
+M0ebKShpZNYBuvgqoqTaCJV4325yPUVTyX/yph4KpHPd6zzQ6WhyvTEIY8f95jd
98s9qBcQj0TwSK5tvymAj/YbRlqXavZ250Q9Rd28MykjA5hwcRO2Xu8xGeE8rARO
TFVWbFZHpywrg79r/SkvIFTTsLWIZ/WY4cK/TgdkOOmYlY5WSJsCdvi66p+sxNv6
W+W1/w6hgf+L+SSZfDiTUPuDA2MXn4RplSZ60w8IxQVN/pRzodyzHe48pZ8t8Ynt
2OFNBgz8FSiHzF120RxZYaEPBOqFj4RturPGuYcgH1ATD00/XHfN2M/hVZjP9MCx
1saTnBcu/kI+a8zVUsqIuf0HMIDlMFPyTMGzkJAYZ0bb+PviiuT+6oG8+ILWC2lt
8WG7vb8cLOXcqkCgKSjeEoCviMFq4TS1jZzkU0Ib52N7kjWf0H0gi4yuojK7Qfqd
EGlFVju+GTETOTyyoC5s+7rqlhcmG50JKv2WVUkxRPZWt7pVoR6/0qWGLzDtnKxl
ga/0bHgZucJWzkQYNFmt9gq5cPIYnixHUlJOlH7iIe1vpJo4GE9OJfvvzJWC6SUi
xh6jP92BdS81kaYNSNKCr4XfYWAGq0GTFHG+XODDXh759eh5IpSLy+AfNofl+TAi
RH6+WnPrlmuOiHlKOiSncBbt1i4eWU/OzIV9lWQMVp17bziOBVm+lW5RX2T/TrHS
BBF5tpuq2H34448ARZrd4lILrpFuHGgnElCjXXqG8FqW1myDKTNOelLwrndy8+Ph
8ncI5dpIik5RYDW4NKfDWjiK3Es8X51d+VGuj862C5AWy4z/xs6i4rU/mJrAtCqV
202UGLTvf2cmiK+5K8YR1jroi/aMXBSGdkbwseIlDOZpX3Xik5E3/38ADGEsKaNg
G51R7hqF5vMODS157vzUQiaznShisfyy16ys62ya40KbeC5qC0ES1+OH1xxCEb5o
NaymwkucERxEUv+OOGBUkmT8saFRKERK2hFgFlywQKJYK4ccPLEjXw+vDj7JiS1R
ziWdrqoKRbWYGfZ70noJz8cxB8Y+v7DvvsUVBUju93qtfmmKNUc5bkPTru2jXut0
aTcZeEBfNa4r6GI5IqgaigZDctz+Z3vtPWq4cMgDab9L50HCcIL9yk0rdloVNXol
K857EN7tMNohi5iyKQavgJrEN744HwspKg+OWyraujOGckk4FMUICMYaN58l+YPO
diZM1RnCwVn0XQDTl04rXB7tfA4WoRFFmsnfE6nqs1upwORGefp9uQpETGfGaLQe
4RbVgZBN+G49rgJC5D6cE3b49DHiHZXYgzmngmTaBw5Yp8jhKVGc+kNyMG4l8lii
rBcfm9CWuWn3J/JWpnZPtfE0mq1VIyQ8tYtr99cjkpzPhNo5P3kZ/Hw3wwyELY6X
xvS9UTjSIGghMRYaDJaClJOcKIuAknWxixHQUbcF5peQyHP+MJYN0DWhBsQTtGjp
bK4J9mJeMCh6reojMhYR0iSOPzOcgrO0Ap+yqZdpVbk6YSbc05q7kNTXHRSDJDG8
a3aKtwuEAfOGUuFYLV0Pju6GTYHsq/OJWvm5S/7ikhgHjr0RV75TyHqIEMkmwSoN
gJle9Jz+bMFOHKwwMtFmpAXjnt45LM3sWogNq2EGc+z42G4dSw4fp3IeHcc0IcGp
uXBBanWYd7Kybjbb9wyccKfpGCroAYMZiQDZADnNGiJfSTpzN/WpaWjegDiCnNl7
wMzOTiv7Es2GjHoBGMM2bV07P6aq1yW3Jkf8phagW9d23T8uv99YNrbuy5FY7P67
g2eOhZQ6G/HbtHtHUyYHvyVGroibyb5akdBSjNEuIVLyzEOYuwhcA7xWCvs8eGsk
mAUNMu/awZBWtKrWjC1msKbNWWNmjdQOqYNLb0kyUaRNaKSlLVwp9sTbvBGwxQHL
tdThqdt/PGKOiC81FILHS5lyxDx1e8yIsQxPdFT9jgk1UHf+1vTC40MhqTIHPMHU
FgwITYH1aLnn+am7nfg5oo7bXiO/7n58G4VHgmVVsvAKR7CujgrG34s6WVY38WL4
wsgZpqVB7dIzvOYeE6tXAPjlAMjkITudfunFLR6odjATXyqE2Vo7C81OEji+pYTQ
oTU1CEKgNoTYY8adG15rVao6KomPBZtPbEtG86p6Fu3UUVZjYMd3j0WAKFURD9X3
+KVc4OwMXBQYFowkj7UkvcaupIXXXXj7RQdJ+fNstZ4M1GDXN5PoJJDA/4+Xb5G+
yTnSfAJ8eUMYibYj6ENHOsp2Gia7YTaao8sDYctQGqmEaJWHdSCvvsDFGQ8tvXq2
AVRttrZkuUlrle7cyrm1nH4jkewXOHMwbd+fA1g6Itagc0IqyBm90ak/5Q4Fcxas
leTNM4ZGNnuwVbnlDt9JULu1FHxN/3elBjNx0accBhTw9pcdzSjK5VR3RRwbw3Y1
J80n5QtT9pREugK6iMNhYPh6955o6ROjbzBKtej+AL0qBa7wfB9l6+sqTnJoQac8
y1o2t52P7oyWwYELKSBb5OndN+ZxtW2GBi7RdQgl3GzEUL+VsfTKTg2fnel8LfJG
SYGG5MT2N2RRMmUPGsfamc7XvfyA2Sd8CHXuR3j6ak4/+VxBH9UNsmbGttts0Vxj
h3DZ8JkKtYl5w4cNlW9K9r+Oge+l0gG9bV4UMCyIeGdhQpt8BxqlEiIY43BQy/2o
4vdmawCOeznNLCFfecRts2u9CS0jmymEgvQsLc2FvATES2cbY6WDw/9lMQf/PUvm
TA/BXk7zvy22f3UWPBHuQC9NU/q993/AgX2ffBVA9s0l8xtYq+f3Ln/mkm7D5qoV
tMtK6rRcAeSwDlA79LQF4F1iEMl3+SQwAO5y7iCVDftxhd454dgk7O9H2RsOx8oV
zMdw9tPhN8OrcXxw43wwvxVXE1pP3Tyz4B8D00NtEwsaotmy6Fgryvfe6PowY+38
KdYKCCyQXWMQwhngayHTDVHFd/BMYR8EIftjqVmKz4EJmo9Aat3X1nMGjdnRXnq5
Rixf/UFd/xtN5u2NpAHUd3SnuVMmkx3gPOsf6R56rUiyrMMTjHj908T6xzay1lOK
Hjdl+IQNcWHnyxvLBR/7lKcfH8VacAryPgX49ObyvoqIw6o/h0L56gGvGKVdRn9p
LgQdrUlpAx12i0+WUZRVCwgR5ZL6ghOlYnS2FR35WcZxZj/VfZQf50D2w53d2rH4
rCEzpTU+nkt0YvbDKC3tQvxc5mnqjrnsbio2qo9BDm7Ytaz/VSMauln4KZGHcyuU
nm1JniuJwUxX0bcj/UDqHURzvCVcVFGSZGnrV2bzBNjeSEBla2bBCbAdHqzroMTd
Au6MjlzZL8vVLISjv9V2tpMn4E1aoYfDYBTey8fiA8uJowsyvMG3q7QqkItJQ1f6
c9VPzdW658hAQMEiE+wtLOsudbhAfruuFWO8cQHTegmCRJzYJoJcPdT4Mu/LFY6K
fkMnDikE4GEjuPF+kjIoddhkfCDLYjL9aPNzs1px45p0yyTlQ3W5MXz8EGjKr1EH
sP1FodtF6R9W64BDKIfmVg6dlgX2Pua/XbyRdJ1j4LVsE+DqDgqYQZpZM0btaSoa
n6gGAKlpty7r2X0MjTAFJdEsEjrlcF+CM3S/EyK6KqnieHlmFfP3AUHnvb0BEAUk
BCyhs1UxSs8bdOp8v1qXcjRAiX2a/IqUs9ptxEo+JkOE8x/xfZ1Ee5ap6ZFvw3LM
MbVuHOhiCJbFRc22SRMqU85mjATMU7HAEdQ59eTHIvYZrfpimQOjFBYsZnGIdXlz
UMlEBarRKZh9KImEvD5Uh2Dd8Pqsp31G/HGwoqDNPCpuo38RHq51v4wAGHLIvTQW
OfEEcv/egSaaZZ+4nJ6m1wanB4tGgltcjFkx0BO7VRaZfX8EzqJsibh4QfgzdSiv
RP0xzhNHkxP3F5mHJdfFInSBh3AfAwv9DbXPtwXzkdYzhAotsGuwmWUVjW/FuUMh
6FfkTtmzvD0eYVmylnFMIkVTA/NL9CL55Mvo/v3KeZuT7lsuu5nvYaTTu8lEAjAG
tJ4BVDWVyV6Xwk5kT2hx+wq0b9qHX7WRGxB/8IZvk7pUilTpSFun+pkrKPr5Xxjg
iegoHdDhiBQQ2/eLN859WgAQVFmWbHfP5rs2WWq+IaDKv5TT8ooVi7K2jYh61Fuo
BNEThmsRAqVH0hi8MoZCoPbH8bHtGmyHALqvqEdcFrtBPBKYst1bwEGhvGcXyXKr
UUf/actyCLnnKR/v6/syAEagh5ehodyM2NaAzHUDuPfTKTxhxxyfQiP2ZPu2vb7e
vh+4VmS86zKqHodrZ9IiAT9/5Fjm/LLHtI0uk/S2mE80Q9nV2JR6LWX+O9hCC+Kc
whRO1zebKMPrgSeKgB5shWXWOVAN7kIvVHGLT7s23mp4m5agRM31a6QhAHqAJiBJ
gL0LYP/hHcgoYfTAqay6MHGW3T5d6zNvz4TTuI61ZkBdzDKywzwD0GVbh2syJIuD
VCTM07ihKFC0ld8PefIBeOqv122O6dL5kFtp7wNHburMujhh9EfuxQg9+4F6APT4
fm88cOb3ACDlNo9/L0nknAaovEDq/zy5Cz29hN57tnHrJz+ObOevJYYLJj177Sov
pYmfvTft22mVlZBdu6uOkLmaS6CGXAPHQTpggcDNldiFKLBw74WtB4MTSdOVCRuQ
3upHtIeDPMi8W22TamaqXXVhMbF7XsW55C9jU/dTFOGoVmIFCzUuUiaxbcjJK1t5
EC/D4qQJdeXp4LaaNlqU2k5FYk1cReMKoe8otHh9wHA6HU6nBB9le4/BV/2+FiW/
LrWBNgWrLaiZjW9xDrpaiVscFnlOd1oMUokxJ/MZefp7zFnTY9UzAHbbFClYPIWc
Lshws57vLAuwsMzrXvOH4oOlvDuhmkIDCH9uwn1xFerK4AU1Pit4uvqt3XB4OFmI
sGRf2AWveEUw3ZM7P6SXpdzwbPkLwx8eVjlmYzJVsvZuUYwbSD+tYj28mHztyh+i
HAGkHufpRm/poDPO2JmIkUeGFwReUIiwEsOsH5LR+UH+p6QCAgsa0/TisXPgHZI0
ayxWcdNvLMOvZt1PuIrwZsJhDw7W3FbIR3jlTBrZ0hYRExt9qG9D5Qu1yn172oX/
PJK5+wxGAsMUlzAtrxGUyoSjgAhDDa2QDOJIHR8iZT/9xA4XHvt0sKK8LaQsgJ4/
dZPVXE7KVhGVzgmVmOtMzZSH0zYvxCNHG+XvUqJfREqOzjypWACb7jYH5+tAal02
XU6r19ipfKvaEb/pLcaJNIrtffjAI1SxocUmVancd0j3x78uTr3ep79ZCrBpK/W8
O37QetIEKYO2RpbV3Q4j6oEdjxtsr1GlM6py6cTfQZcH3RIinUR1SoHyvGWCcR8w
HdXY2D8J8v7WATwevNwYS13raLen37WpnYfWVh7VOVyK3lHJHYgMLpUcbq5F53wP
9exOXh/QQbDFV1btD0BTz2otkRcIQqoKYw/QxhY/h3UXcDgQZMeRclI/dfpkjw9k
GA+O9UpTZWMlwLXoXof85aPVBKVfrFSsqTQhJVvJOE7rnyOz2VgW5SH0zte4GZG4
UaYYesrk9XPpLgJH6hXUHvJWa5+uNEX63kKTYiLkT87jk6+bbJU5zLSG5P7EGTgo
ibCx5Ap+Bycpjhk8hYDjsrOStlHugQMY+a91pFQXG593m76GfQW7xSS29eFs3akh
4rfsy9ifDrEihAwSll4s6QPIZpx0hmTLqrwaYDm1EQX94/3UA7MVza0cOlSFA/d2
iINEBA4Njxne88TJvIsKKiVfPM99L1reRQiHEwvokQNBOGfpL8dQ8m8QF6StkUAV
apkyZEpSSuaa5HgU1mAyPukbm0hXR86dc8Za/P+XHFZ7f1Z2+IH/X+W50THSaINO
CaTbaRvncSCY9idh71hSsOdZv3zPnff4//hdJYosewgJBUuTgPxEQeMIyHfKt/UC
TVOb6kaAJuu2cEM8u0PRfOySJyLCzgxSUqbOPqI2ldjxjUvgrIpD6lDCHpZUprGT
ImtZ1VI0KJFPPAcOgXrGIA8Kig5VVS/eOx447ATABH6tMpBjYAGlMtRyJ2U3kmPp
iimSlLatLFr9twGctSxIe6CxitlY6EP1cIcN72Gl8OkoyE9hBMi0gCUwv0S/cQrG
FxeHsJXSFeMHNkxj5XJPbSYTcqbNjxEoycnfUvoWJfmAXQ0rr+LVG069S7JlfQ86
QWQqMJaOk+ivxGRziLyJCBnlNZ9FFwUnTCWY4edJ+3wRvfcY2gfpf2xhiYpidE/5
jJ5ibUWKpG4XiLgpjjWIaZJG+L6jtM5UZi0MidAwuLF+/VMKan/c8j5EFoCfB8vx
YPCNhNtl/aKQ7y1oh9Og2aj8qyHZZnaYc1gSmFR/zNILCgFOwVuUScbW7yVc+4q4
UBTP3FOr7Rt+Bkqauy27e0N04J6Z1NF3HwYNjSYbDxzEqeZg4u+p8dh4BQtpBzSr
xK/oZHdSk44aj+x6w+uHzIA0DCUuTreC2zksK2aQH5vlO1tEeCTE3GBAqbhdVjK3
m6vmqKY1qHA0LJmuLj5NKIGeBmURhVc9jnCH59zFsB/UHWHunzv6P9uAuLufAZKX
AYAixrcNdL1zCYj8SHwi3pjUZdRl+I/VtQgEcAOnxw3jksfuQ0T9jVsYtR+wGRIU
LUlVTsGKobnFsf4sNxk21zZ+5MV/K3ZQE4gPvdeDnz3mCGWnf5B0KfaA6I94qWQw
U4zL4/B6J2tqcbJuELpZs1mnaB7POwwQw4YuP9e+/f2bdkb4DkH2zvLddAg3/8LK
ZC24l0HW2yMOLu0Kd0N0UElxYbzLiKO9t3If3dgfK1MeJF1/M9IlyZar7yksWBP6
vqF838cvC+5M/XSnwWDgG3hYRWs+6FVOCbmBEn/zGdgKccJ+If7Os0Sk9HTr9VPx
i66CrZ91E8FD+AH+k4u9uEI2lD4UDySGwbKfKOEGTRR43Kd6I7NdXYA3af5rTSTC
YBz2pBHX2UbWD6gmlH8zKhNqwxle33jAaIPLDiR6Nllo+0nGQ6FIkN8oiwO7f0Vs
F7oH8kgSGRnhF28MNjPTvS7VOq3I1NYO5F8H3o7Guy2W3JOwG/YonoR+j9H4/DTB
/uqAhlsdTQbhOJHlIeHdwQxCHkdNAFrZCm+svton2Bs+iJYlICgeo+w49qNTHcED
8R6fY2m4Yw2FUrUaIGkL5FQemZlXKikcsPQIHjRMmZdsvuuzX2UwkHQv1JBhjhJz
6BnlvuxPC0+tD6CT9LEM5zCTc0PFrXY5H6WDKxxRM/k3JaZhR+1SIVLbv4xldCeE
YCvfwwrCXypu/AtgH19eS/qNH9eTp4OpnanVBm02sGoCWzX4NeLwWljSMwoA5yAg
clxGXaifzO5TzOf1b84se/rUqy/+63cyERKZ677HRVYIGuhT4knRfBZTmEu79zF1
suCj9oHpeDJGn01TimjDPxkvoSbKgWjvmjfajDLoZiAoiHJc7EYZgoVYkhWc3wRA
gFyFNLRX/pMa4qGkosdEFi4kLyWtq6plXCCn6Ys5SOT7O+pAumYUr5hq6MKzJlDg
HS02TVIZqr+XFp8uICLTncSTsw4XpxjVxzq7oEiITJ3pEB8zR/aXP87Z6CtunKNU
O8Z4NK1sbFJplGGO0x9RSzWn0Qprpe63rp6nuuqVFe3lqPizWb507DTwB3fN+yv4
RZLZ2HY8bIUnqpUoV4XCy/Q/AXOq1zyU6vVFtGnJhh3zovNbOGwiygMq60ksA40B
mazyg3bqUkYd+aANC5PWsuqAREQoD8eeXc/vWps5aHft2sEqtt2l7zETe/6NK1XI
j8NpODb1g4P4kkIR7AHmWIDmIG+NVPU8mVik/U8VXp8qua5O44w+Rb9sTsTHqbfR
lCX0Zy+OCxfIKQYYqyPbz9Qhcd3ZNGpQgvLcu+xUjlfT2IPhxUWqKYXyJcXgti5f
WdM/JjY0faKHTV7PM3RstHihWp4oPgnVz6Z1QQxqwyufaS2Crtf4VqFCdCTGC46r
q03oKrISOejXutmQvavFY9G01TUNmiKzXF3lMRZdLqMS307ItQxAfv1N34BGV2G7
aVvVWcos9q9Yse2OD95L3F4jpnPx/mULMG/XkpZahavq78kJRigeTHkNshiWZhbA
SKpFbIJuKLbxMnXEEWUnYb21cwkEtp7cro6ZHsI6Wq+MJ4bOMZRbjY8XUH4RV5Xi
hPvXPYzwTOmqxK6n77ebuIcJk6tPQu0yBgrNRNmerl7avKcKRUZ0xj3VK5W7qRBQ
gW04uUlE/9f8rgb4SMFcJ4GdNcEtIlz95uJpC/VNltX29Dhb8+gcMJ3jIAACZsov
XEzpRnlF6HPsndTfPeDUzQ3vGGSakZ3z+OLDrIM7HCSpVMuI/L8TPimF6dBH+Wfv
SnEAbtCoRXcgEUSHCUE6MEwE8YgVaCXspcUYmCPFpNFYYFJZ+fwMa+F8rx5Ge8Y/
WvnUZlKCHYJS7nHG2X4agIiPIFnQAbSSVur6B5bowcf6XVqHyTma1khUnqHEMBBX
cdV+89KZwKbyRQP1qxN/UKR5i6jw6dWRaxBPhY5znu5rcnfCtR2ADmuAGNsThxvl
xV9O3jIG6sOisPla7H0HwMGN3GgbLVSyfdCCVB/WMwgoDZzipLDctGFbhPydcoOR
h+CVUoCJmoc5OHsjgZ/3ooSOLZjRSF9Rhg+4lyiQYF4EJKAhaQv26HLT0Onty8s7
GgSwzRqhD+ukHQlo8cOhy1yL7dYy3B+dzyU0BedyAUoRbiEYK8Ceq1SopphAPlO5
YpNdoApIAMufyhz9NVq/40MeH3AIQ30+FNJUlho4UcjgXb7VIrUFGMuYFWrCnogj
6r+pSnM9K0yTHNivcC5l5LlqhwcQ+VkLpeUfeawW/MH78hDWx84uMzVyjaZn/3oS
LpZ89frlPZ1IOp9LF3fp4+n01sCef2dmALlnAiZCw4fmd+xX3yveA5y3hhAT6d4b
w9q4zIvKc8MlG1dgZjICDYiOa1Pn209FivhYpMdIC83zeWZZL6jCof6LzHusmKCW
u5V0utO/ytr37PvQYkjPsOR/vXbXjz1st556ztWuvuEgRInT0J6g5sXc3wSdpQQD
ilxhC2wVCcA79H5URHe7h+c2XGhLgkTNYmp0WL7iKqQp3PWxkEGdLJIj+u0E3BFJ
PO09BdsbNNzWDnUV7gyhzI/e1LLF60n112jz6Kg5kubRFb5sz9upvBLOiiwUA//j
sO4iGUJrkqE36+oWUHeovmx+yZRtrSU7462sEEUb3UYFDcIvHRWLSSQZd/XsKYpD
y58Ayidkin7u2X+BwwI68KnSAscTr32YEtmIXAoKYS1x6XK3e0L9+oaZodzePFMz
o/nQX9RaY+fjrRKJP8SU1emogSnirg0ME5ZEDOLhdkkFUsrnv220vroJp+KfBjcW
N3YetyQ5xNzF+xlM4RIKMYv2CNCRdVxVis5LTPfcRR9BcUCk8M28aIfPyk0kKm2T
U9PU2K23OzdOR35J2Y9/0QGl9scw52SpqTyEzqhcXhuISr3K5fFonERjkla/+Ohg
7fe9lTeOGrEcaHeSuBH8gtmcyfhreMjOJzoiru71haIXfbRixgzGg/pfPtk9QSDE
hb9eu5nX84YI978nA+Sriw48KSGQcB5wgdIP5Cmipl5S/n/hEk93F+KKDmtfNcoA
7SsNJhpYF+k0CsYNJMwJS/ZlbwzLfGT7SplHqxjvZSsl1F6n1bYOERO8wAfmXQue
/b3AdUaabOtnK1SucaTZaM2RPyHf+ZJQke+mZL2RVa8iR7R51zET2aK2zrWhwhqe
x4aSPkb6j47Ywyru+MFRDHUxx2+fzk/buFpa+cBN65ciCTvMvVYh2z5nOoLBDT7c
5seCIGs02PL3abavzJdHerwa5mW8OPgp1PBtc0GLLMb67jte5VO+jZd/HJIL0Y/i
EkFxacqllxD1kTy289uZrHynsfnmcveskgBcM6dpqpbwsy5JjxkKQlkmJPAVqaEN
Zvt1Nj/Fsf5+2dUzJXt4qb/GJlPHC0wpIQ9krEkay+a4iZ+9whjf4ABFppcNEHrf
xaG0Gn5fSl+z+jekJfBw3bbZpZ1nSPSVEH3X+tKKxTUWq+Ezhnb3vkxZ1q6xXEWA
NOkFaxabjt/EXFFWG7Arm3J2YoQiYonss+FxXIzmpPFfESfANTd3qrjoTwySF2CP
oV9tni+qBZhzhtIyvcxnCD+dTdWOlXiXGM5gsWNr957auwIXN60pk9945hgNXug2
dcF+z6x2Aj+ki2Okymcgd/SKvcKQzEX+KGwo7H+D2NXd2dM2YnZe+ZABJ8vTRebz
B2QCtcmhaRuiTO4iffRPpoLIA6p55FrFfurX4rwhwHHeA5ZMO4l14uwvvqeYecqu
UT5qqol6G+2dfG6jXbKrGbTDUuZBRmBhCaS8XTCXXhB+MFzE3d6+IsjvzVEdHYSr
TI6lfZNKMtvJm8aCv7rRZhIEfalTjdLIQXDytSnms91zTNNReSiZtO0gcTUK3jLA
t0BcgMo1Mz7HrmbYvZHnmq9FAZdShtviFvTM6ijPXFsRopk2Kt7nx2tF30ozKk4H
BD2+afasv0j+2avq0WuiO0O6uH21N3zwiiHNrFcKQjYA9kHYNjBxtUpTC5DE6fwW
QegR1EG2fGAO2i0J+T7h2BVXda6TUwsU8mxvIoDLL7ci7mz+cfxS0Ah8lfN2AvOz
2sXaX0JuXtu1Cw0LMoY9Him1K3A3WkJUQ4tQUwjbxMjRfRvw3EDPjOtv1oXNF/0H
Zu8+WQQMWHPbR1U9+JGhRmK/MpnopaMBQNFz7tnynpy2mHih9zLEdHmM8pfY4Moz
NECQ80N8d7GwsXRsOARpjyUUgUztIi30/cZAq+nfJHhNtMl4acjOdDsh/1yvrssW
EIJMXHRPwyngw+0hmNhRoaDaTqG8ZOJ9WKL/ZlH8ir1CWpHSLoAA2ULmfC7gxMs7
MzCH5Io0lvBir6v72MsskP3C95GhR6FFTXB6iUq+JspgL0pPtau09ctETmxdhSEf
xCIgxiI6vFzyMMh5tGcQbSxpXv4iC3Yzt15sskQk3bm0OSdB4CY3UoCS9wKnLb5F
OXAFuJ0xamZYBQZWGKARQKDIOqd3qwxpWzWq00ngWF4LX/z3C/siXEqftvVVbgED
cnQ33N3kJXrfNel9GkSz9uI86isydXo6vts73J1lNL50P/l1ej0tXUDCiCzEtyOZ
y0tYF3GcWE/ND7fgKGyrbOWaRjRr7Mg9JS0OMQwmHWssCJtRUr9PYhlzjh2XXzw0
vrBTna/ZDruHmgpRtjjFaZdMfVn6Xmlw9uJrmb9cPkxKgqWW3GxVjS79YZdOwrtB
5XueziyRPZ45w7/xu1CymjDIzR5DjVdGoSsHrGLo/QaAVJtcIry+TyitHN/vbpVa
uXqM5K/5T9uRIZe4UkoeaG6N3v9SWE0Ps4FInPUQEOVN7z+AZczzXQ8sIT5HpGjJ
2wuioVwFDNQPRi/WGLeqQEgNErhWdyUbA+rg/FQr6isn6dns6lAOCiQNyg0v4gmV
ebnZjunTf0AvuGpIVn5Tkps8Mbb3mKUiC11PzqHZ0iiS1X2a+7zDHmun0ar0MSAq
6M2beE/W7LnFKdDr9wmAvey1rcJQdbIfuuEBc8ZOikifONlXHoyay7PzoO/57sD/
n9wuowIxQn+wf8kMT7GsTRulHtKzxbAU4vpy1reWwMgRYbtklW4AjuGGcXPLy9Sj
Jh4Pvb7IW6LNJo3J0Zhu13M5sTIMJEK14wnutJK7Na6764RdOMAAV7+fWY/orYGi
8pvFeFoJhUgofy4ozbGEnGRzigLujVa3mU3wNsnvUzZq6AJsZyj4+IGKFWu5LOyQ
aJlJEQARjuJcex8jADgvfGScgnCM4GTqcA6RZUQe/GTYD+X0rPmI+nh+W2J1f50j
Qs6MpzzFuYhwnFVwMM7QBm5dTOwacB6RvX23GBxF+Q1FP+S1IqBIOo6F8diLuGEu
1i2vmx39n63JYjGVOtjS2qR63CmLYUEX/QYEhoK4A9usiCcH/Znm/bSO3R85zJKj
3oA0DRWxKoanEtcGXm7SEKG36ArugvBzjKsYeYAgZJHu1pXPzYWYVRO9fRtMVSc8
kYBuzrp98PZ2qNcsF24RCLbt5fctVwagPlVvCn9LcSsLZ1z0LDCx053KCZ47Swv4
rXf9ZbEAPbKsVsygJlbdZCw1l0dLKLCXe7gOKhjp8+Xnj+TexjeGFUycrJPWpmCs
g9WiOVBrK0JGAg46/KLwKVFrfR7KrxuTksmeeav6bnrybMkHyjU3d0IxkrVdrBO6
HS8HXvhFDpz5NKyepBElipRAa5a4znohZNfzM8BPl/lkGEl224U5pVsWPlWKK9Ky
EnqcPjrCuesPVeUSrZ0ak1c0y99oPk8gUjbB2IgPxTW1G0UtiIuM5bHNTAZdhjW5
yVW9JuWI7pIZCDwwyELfX7duFBMBiOSmxOCSpBDMqw6QFE6/uPHqcff4uR+g4GIj
GqSt19fvOJETxvC69u+hzCGdcYd0CkmdXfwu+c4xGgfEdIXMuvXN1kvhyKcrILxH
5A1WqcjZ7AR3kAefV9bIQwU9SU1hyminDQIWAw+koObxVitaPISHn0gPrLNSYPem
l60RIiKumwFvCfatwFVaP2gjkxcyTpyXuuxp/seyLLrq3XrAHjtZopA87/VFJp3l
k9A9Kkx81th3pCtqF5P1uOoR7tb5cz28mi1hpZmj3fdXO3xgztsRr6jrgBckn3T/
LZrdBx9VoRmLohhv+NnopH9PfQvG685853xv7d0Lb9ROjR+rg/QULblzL5Zaym60
eDKZ+/h/w+KuCJIS5AUgiqyy3h80g8U1hqUFx6vpt6daxyNlFMUeeeX+YAiXhoDo
PPGwp+yXc1qWdkmFLSP2/PdDdh/ApklTAJOCOcHx4mIdIxOBH/z9mmziFRT1mE7i
pyKsj4k+C3LJ/xxEuv9lbPdMgf8iyhLGSJZp5Jrdh7PB2p7ej5w1nXMt5O5VjetD
CPvOtyLOsu2qEQYC2Utv2BHXiD58UnDBJmH3Aa7CXco9vYVbh0d7obK/S/AK/M7/
ieFPNxSrqfPzBUyBYuNWzj5mMvh+cwXYHuPgZsPaOsVhawBn+508TYV44o8eLrRA
vISzH/VaeNdIHMgmKzSHIPJzDrD37gF1uXdBzBXTGBDyAI+sYBLouqrWVcPWRHnd
sFH0ysusyXDcdUl7FOWy3be3EkmgNVrZR3GSeTU3vUSX33pFE1ui9Pq7qhxfZFoZ
qRPKz2XPvXGe8GH+bj8aCm84mNhtCCowHBDbx6FZ1pXnkW+GGdSHggK0Qq/EWvls
zU4CpRuWxd2HOnppB3Lvb65rKhn0/LUZSmY/qitl8x+N1gY1YqeEdKSiCGi494cs
IBxwuwnvc3JKIBWYyXZorpaaOiwnQGidLDe2MZf3UYCB1hHUBjV35bCC3NOg+tPq
oePmb7yWryGA5u4N032audyPMZOe1s+f52oxJTEVvuy/q0ul74JsC1yQWOFlWvfF
Dki5pUPGnMcvbjchr96z8On2QMEiVDNAZkmpdFBcjmMR+HcK1AXNwlnl57G5cY9g
J3LU0Bc+UIt6YESsOYwZECWLtd3cjWZSeFD+ULTSpfAyWS0Pqfnuh6leboZDyufN
/evbyHHQUN575DO9e556K58Er2Asr18UzL+arjMlarPzV6NT7mt/NVk8VcyD7EGi
JKguDN9+4QQUM1vzuPM6JWth9hDQ+/sHCw1EZf8Pv1mxdXfjIMogpjvqQvAKMbjM
BRsChuzxupZYxzaUavsEv8ZASAcOrodpHdXPLcWv0vQbq+v2ykT9e2diqX8Qxew+
eUDN8nF+Dodr2YjFemj8d5CJABCPQ35wWdmoIaPeTX746GUlAuF75ODYtu/RrSP3
mKXxXJy0CGvPsOcNJCcRPg3HL84cri47eOlBHkz1lKL/OVwtH/goFLFxlulHHf2p
5hWjGj1ytnb4rYDIJx7axn5yh+0/zZuz5nobASVuYn0RgqJKnYEF4TDx6r2A5pAt
jv9pEhNvOm/YswQWT5MqItsz0czHUVfI410nhqvhSCULLpMNPHQQ3CeEym9eloms
YgDXHvoCvPy1/1VCfi1vUTzCIkP9y98buWTWRlMSAgiAcCuXhKiJgFp4Ss8E/fQT
XXpI9sVcUB18+FvIlgbyEhAlWgj7meE+uk9gcykUnwXuFDzAbj8Sg+Y9bkIuJ5tW
cj1YBjitfDG08JJBXHH5PL/5Yyg4FK1CixQ5fD1VUrMLGW7wt7/5uLH4KGLGOSq+
PW/WvBH6iltuecFiIEFwUkC6bL4tu5uyri86RvX+d7bW7ZDNwkZjCZZAOIMeIsr+
38CAh1Ey5prrcCtBTDasYS5/CiA7B9O7lH6UJfAvdose3MgikV4jm46tVBTf3Kuu
LEpAvbAbXDOYufBVv1nFUpq1ay1pXToWDgG2QMTm4LHBoqQ3P+qLWIUmebeV1hwV
18SuwloGdpYEHfkfk6ZBbCWs2Fj0qLc+YxbraQsHiWXDgIOrPn9lXKTk7ZWGWNbu
+hfUfRxLOyBvst0mBwIWFEZ1EPNk5C7jWvBJXzRuxlZtDe6tQjFP472myBlxJMWL
2CDO1AowwajL/rVzuGIg3UMmhTtlahqsxO6zDSsr7Lti31acdrQ1DwmNXVoq7e5D
rRgIEl5Cu2XsnFCFpcb1E7nLtvwYZj4lmDZKcqdKmKAbRCVFfsXxBDQV6Gs20cHz
EiRAogo+8WpaoFW4SLZNL2CxDjyAaUsLdMbbXgHF6TA9VhBfAQ2X0gXwRCAXQklh
v6hOQqkKtAruvGS1cbG3oZjsYVMTgiaY2sHUnaAnNEytaB4sjkGtbt6YVS/Lm3bW
ZefC/FUb7uCB5SrYxsaQ1P4VPfV+PIn8m5FGMf64pYWjQcPoQKBDRGB7Gv19yJq9
uyWWmNDtcZfEqc5jNtb+onpHDG54YQzF+T9CjpRQlvzoCAocwCDXePSMaW6Q0fMy
93vTuNHtie4/e20Irs9wAahGZJph3ZL8exSk4VtT5qEZ2dftQulo5rU+KSnZY6Me
3b8jsbDiibWQebaFjNSPRYTEfSUTdq+USpPUKGXpXQ2gFKCHl74rU8SjoSvNxnsV
5MDw4fLFLfH02AWE4mdS22PdnLtIQ0sn8v+NDfvSyf/pcwngMP0O3mJHNhdi7Uz5
pSIppDb9qJtC837R3dvzSpAlrHTsm2arKjEMi7F1oYl3AzUxZ5ReLNyE0YVYohPE
T9w8etbKWbREsTga8ee1+XpRhYGnGLWsJTB7ftzgp6y7afFwEk5HnRWoZNH+zsuJ
uT7wPYTgQwhTfE6cA8LbJz946Ox1HJIEl4zMJ7ms1yUe6OM4mbkAFO9Xo++z6qVe
tD2XTsKKWaSvkHHj6R9qElwE6yiLkS2BgApEhAzeXKTl4IdMuSIL9+57JAt5sR9a
VIfhWudfq56wbPDyrRIJBowJh/dQ6PDiRPQ9sAWhc2Ei5lO3rWzOZnHF/iw3b0B8
jfwkOSpu1puDccWaZ4wrFe7G6ezvfAhHJ+qAqSo+s8kvxJ7O0xvaVenyI4jeT38L
GiMHxSC48Sbl18VIZ+Fp+d6onZgWYhwTARkr4uHPcdHP8oKYLFHMZzq0kiElukza
b3yMalDisICJWhgVwAIE8k8Q1qRjB2Mt3Ql4whGcCfts4xpx2zUYHODO7waaoAGp
7IyrZcr6XXSUs6WRIPf9NrXioNjKpg1FJSZycLUQYEQZUTLMRggjSlm4CTuorESP
SrOTsmsbuAGDeBCDhm0h1YCmSxcjvwdAumXi34JRyd0+7qrXw1NVzUnympFKaDda
hok9Jbc+jmwS0c4OnVv03QDoZc5dcbEhRIIhagTGGU+vQJqTl3wU3bv34iOJ00O6
5DNDlGQ66TxXditwKpZrlG8dLSKwyJIQqZZ/ak9UfrbWzDWhLo30Mydb+M1ubTTA
EXx9+YECORANo6l/O4/t//OTIzhsaT93PlYW/9ZeWFGBmLsT9qp6OVdmV14OhoL1
tdFy2QMvnzvyknmpH3It9pa51524ykjKFXScwUuBFZZjxi5qOkvrOqTi5zAXx3Oe
Jq3NMljIguheP2PBYemyeGUfP0RLOvhhO+2e1pL/gmXQFMDc5RHSNJk85I4bEA0t
MRlP7KoUVl/Aj1MNIoLB1pprSsS9Em08MKCQ0KRvxVzIlH//M1TQTAlxOYVdZUn5
eQA+nn8Qa3KQC7c3HMv76fCIpPpmmbSMMI46MB5P+SM4vapP2LSMj4YvlGEufkXp
AmWKHgjZgbsZ2m9AV7Lsu7FSv8esQl8d48BWSNzGRkFjvmmSDDEeYOWpH+D1RwRB
lJlT6o6Zq/WVk9xyHeVH8qgZr4JZX2VLztEcWh9kC7YxIONFbeIZ5W4aqw5ZlzT0
/fe9pVCX7zxfjIkeenDQjjCWQXWaCvi8msPTha2AJXsbzQgbGzMxR/UAwlB5Alzh
492FCjFoQS5DZSoKwEMWG09SgpkeE3m72mSISwdr+HrFOmIpuc0FIJBWsT2jgypJ
fTmJB87YVBNAW92sR2SS+p9HExpWKuOcUiXQXnguJYuaq3LDq3JMisa2UK65JyCx
3pGyGOX2gGjp9hP9sy08S/X06iRBHw3S5pfXMJgrS05TqzAW8zeMoppxqFvpl6w1
W3gDPs0c3OCq8LaFBEdLY7dPjLlyA/WcjEEMIdDr5292dfFLLKVfBxd0a//RyMPa
mTUJGeVj+yXlg6tKdPTTIfnRNY5+R3J+AfngPwVG8hZdXTv/lqa+xQvKRQdwIhsA
xF/z9idfepXW5xdEQMAFSJ1y3VI/7KGCxID1wugcFCNWtkYk/cAQDGq6m17g4lZz
bh98i4NkDNEPXyFIc09HbeVGsptU/cu3jY6N3aliunxdx4YtpylhVRp81q2aAO6k
RHJcH3utKyQUtqrXerp3wzt3jfrnsUVEdyqnNvTpcd9SjSOjL4g04WZjSinaOSSs
RtocP85s9UudNXY7c4zcHvY0beO9RBi15jVHYn/cHa2TRiDQtpmJBhcTs8RpHjcL
lyybKsBZ0yOKEsmPfWjeLEzKhHJTVpxFJuvvj5f6ngj/RjK+U+5Z9cM0FxJH/ZMh
Rkx1U2HB515x8+Q80BudyUDC5hT1CH6u2Fq7pOoDRl34Rx7Iqtld2Ms9V9UctgyF
dseaSBlSK7TWgjg+ti9EiDRreNfcSL76n8ccasB+mfhBgljzVs+jJBOrTnzrxJ4L
M7wwFe9FIGhcy/YrtA45xL9OERCAlt2pWvAmN+u6kaxOHJhBph6xO3FKn/i6qv0H
MdUh688rAuHvpi8LufoO4OmI+8TUuH16ewSTguP+1MtwYjUZsxLXihy3Te5BR2P/
iA8wRx1Xu51tViffJh+jwxqn1ebdv+QgOHySA+MhVdbOpBT6MhB3q4DskbeOT5eB
wxc33JDOV7LSnccCiwHgBI5rRipdnVvDBxwmz79AOc3cx3K3HwOSmuwERgf2mSX+
axmK55ZDo4o5pAx+N78h+RYhLEXTQHRZGge83JI/64mwpZaBf9B4wkmONlIZnEsQ
NlTN39zus6jkWKAIapUSE6t4wxXprzFvQucDUxzgCoi62mw+7s+1h9ry9VEutzXl
dJsahwWv/U2LnyHMcWxESttR+CTW7hZu1UdkXDzuaj+1NJcY7zqrFC4daeOJKR6H
D5jsJdWg3MCeQBd7hDkGoMvtfln3ATgicL54yOlUW7cjSe/e7VQCUEw6wSucX1gb
NIWzxM+9lviZuRyUY9CnO5e4CRZwEJock4kp24+gTmnNIpsyz9Pd15gLfseelNQU
8EXAWK1gWoEM6iJPFbhrcbY2L4Nbg0oj9ytycGe5aelBuaXMad99SzSpFkLxYRUQ
aNG5KwmzSnedLiHKNNJZLsnk18y5dYf2Ly5+8G5S7aLXgCE58/D2xOKyBW9HjV9h
7+DzTaOIFap5pOUrJR0sn0AkmSTLJycIZ3vhehtk4NwEWTBEMPmLpihYBXgQeqzJ
l8blyb3q9w3KINePdNHbv86P3eEQXt0nWFp70aRlKMsJX+vPt8wQk6xyJwRi4W/P
BJ6di4kxRUBnt9e2AgYR7TR69hwBq5SVHcZlvjzFGExel0iDK17kYO9UqAnfDQnv
zNGqZTBzviwdnwtD3iWyey87DVhVHgJr19CB+34kXLulOPYbo+QSdh45g/SRqLSd
6Xsv4VxUgdrVtIv/EPMlUZYAPuFNHr3MGziApH6cgbvZYOGPdoEbcev17r2PaSDW
BuQepqvr4c9j4Nnr0yZoMcR3iaKmJtaik+FTu7Z9HH6LA1If/px2beAt+VvPU998
KpfnJ5XSsrkPqU7NzNBC7rmGIfU0uB2nblr09goauFXBgnZ2q8OdrSdLsvC9LiaK
323QczuPBR7I8R4FlKjd/qAxvUyNzMl0sLegzQ9o96CjXIUP2+f6YdPjnbvRlxzN
ZIZhYtV4o0r3Gfu4w6ojjhoaNHqC8iWHCLOC+5IQysrdTJt2eL1tTBUrdA1r4eqg
aYbiSVJOSHIiqPZE+oS4ERL6k0SzBWyEfUL1OXawcZscT3aovUOxY8xZ+Ryxx2Le
1fAeLtL0SOhwOExM4iyyNbywIq4UApb9QU7DqNTaREHLWhNX49/bW+0WDlwZ1P85
RgP5Huk4OaP8d/zORCTHAhbt5PG6g3BnK2UvBpBi0FJ56bHKfpRVrmZlu91CFHT7
B2hIXL1peHoOqddzk+/OS2ll0N9Hs2iS/FfxjoSKbpIciWwiR9wkSLVGDGGVjJnL
TcLhw6Rkoro/mLJmLgMsujo4ZwEO6W9t7u9JzIufk7CfmhuCNDQoPU/oBcRA4YIG
xAE+X7AaCVj/izO7AMXUjlC6iwwQtpyZPq93TArmaU38Dm+Y8PELUUw6AN6imAwp
fBB6N/GL55FowbCi7NlWwcdnG7w/6lMhj7Yp4Qfw9Y0XZGBVBq0Bm+mHbb8m9ddG
4FXolCCsaML1bjlyoXYJeJxzKVp9nxfBoBsKRjR1+TqqFR+XsV0a8/jSW8b7MjtE
G1zeNzH7IcVfmJeCYSctPcdbgHdPxjcgWByGxVlAWsuViZiVTX9pd8mctAHkWXg6
vRdwtl9NJHY4yOt1Hd0JMkKEebnr+sqTuxthQIErGPAnB62KsrhGIwPHzpToZa9g
ehnDiC8BZ4a3op45ODCdOD/1cEgZObFxbVHXHmU9OwwFp7NRtNZzLLpjjfkf4vEp
Ni+AnrX4iLNhKaKzu+KnG35WjRPRDUWezib6P4gV7tVgn713Z3hWU1p5klWN7Po2
Mabp0arXo9Xg+vAlvrxV3COjJV/VZcF5Vsd98RVeAL18wmrwPggitgAjPlD0sUty
lSsF7LacSDw7O9rySJ+7ZSA3Bo/gIozDZ9hJNmcXAhHVowwDSpntke/wxsFXdCAA
q5kfrjD0gA6hN212E0vIje8AACphqvle0wwGxtuc83GoxWcuQ0E/I7p9pSZcLRax
nGz568nUK6kin6+qo4vmgIkY1LwSm9+vw58P8a9Q9/P1yGKKGZ2VZCXaB8kabJR8
1GhBvYFYDeL7p9rkDb5HWKUG+y8nYIWe8Rc+u6E7yr4lCJXkWdeLkCtsc6HUMi5C
JCnC1kZiNvBH7qZGsDIHm6nH1YSI+OyUyTjk1zgBwty0uZ2tpWX7zLyZaJQowzxV
b9Ke7HH1VWuY5EIX2HtW3X9QTfZTuVG79G7fKgGtWVpZU4Fhhmy4EZCyL6z+Bii5
5NZPKIfzwoSRfclaNimEf/swKkhtwIdb1xzK2t386oW/YWOY0PtUZMH6SOdu1wpv
KdwKaXcn/wOhBr9YfFH+NFldyx+mgpW8QhraUXdz7wJTaS+//0x5Xfvh5+QkF+Ms
ZRSZdDHylr6MQ+1rI3a446DTZBVvhqO+nW1OndebWDyQVHF88A66fGw4cGcZ3GuD
G8RUeehJS6HrXrevqYq33cuXIVcVa+QIU6mpzveKcH08YAgIyRuAcrRdHdi0zUzO
GgqaZ/E39jKUM+refLOxEPFjO6Um1AwdQduaNxfNQbFK8SSjCJPgzfyg+sgUyy4H
IWm4ERTGsQlG0dB2ykp4y/iViPFOsXfVHvvkqeySGAqu5z63toXBOff5eQGpFnH9
0aT0tbCC3phSxtLxeWkwj+dYBP3eQHaIybB1VC4LHJlhCrxxsgALiNECPv8sx4eB
+mALnzzdojlJ3RvJm/e3IvGkrxVOwPqFJdriT/SJ8GMJCFCtJ+DLCZSFJLgHS5v8
u7/gtyFED3e+RCsxAPey3lpXa4vr8RgApgmB36XfCeHiB1RrQs0zjlmpQRKaOwrc
SRlz5bGPqldBPY/T9Q4qlOlLSzWJAjbSVc0HWH634qTCXiaudy54tzd/L3bqcgx4
GLOa71WJrT/lyMWhfstNgcizJD2ohZ71rFUwocBG6Zu9M5NhUwT3+Z82Q5VbHhin
1jSwsAdih9dH6oNELi0MejptKm56k/CYd2FUYKfNINz3MJcnYF9sIGgTu3F8tWRS
yW0QjyHeVMtmjZsIeitSU5fWco6ApDmJDFqmLslY1kU3QAjWcPwKF+Ffv+64rVqe
bubwor+o5jDxnANcDjJi7T2CKf6MAdmqOqMT7X6I0Uvis0avoZOF4uUU1DZ11j6F
IRibHFWO8obFl06JRnLQl/VVeo1mnKguHXXKtp/aVeAx8QkdngndS1BZlE8zzmqy
3b8WIvM589E1kuvj1er7HMcUhR/QgMf51uL/lpsxTbfv/xLZCZfugb+SBPtih8Af
sg33NfCeY1N4u0A1TwNPvkfnziN/rZK7Y47JGc378ZtyE4koR2B9Fzvv8x3yunvs
zx/rxXNz6V0hWZDEn1EJ9LjT11RxJ0ByMGILNjsq6nqmM6Ud2xTwR3KjMVBhcITE
CNnqNc++JVT4FqGQ4bOCOGu/k5+sduHrscqCIJPhjZq9j3EfRqeM+C1RpzKcM8b9
9HeGRi4mcSTxjjdd6ktWPPOeE57qWEm3zlKCxTWRXUYY0WWWjWg+IH5oCkYpwimU
xCPsbp4yQMDPFLUBIup0qplehKDdRwE85XlqqaDDZqlsVUl25tt0aJzXfUYg0dKr
Ah7A7CBzsyNlECry2UagPSqkEgnZTmYI8mrR2FLtzHQK/x8BMzc4YDj5aGaDeblW
FPMCw0Sr8cYDHJuYU3JfmitdQ2HKmoXhuCBMOiGxAu4wkEEpU4oX2x40fieZCKg/
ha1TxpzrQ8AFSPWUP5Itew2W0uiC44SLy83iVthSfByNwdu+lJYFTPa8+km5G/tS
d8qlUgf1jWbw62XIP2MErIAwckQZ9NzKXiWuAEUvN3UTNaoFv5UQAjycUmbFCnLF
C+iqjKHAKgNgGuX4EWYjX0fUBiwnwqdCdDx7buWz+3OEiAeV2d8DEBQKmGQw0dKd
scshe4lfJ5/SlJ8CgPG6D/24aPMuUr3IJ1C7v/sdLXGn146izFS+B7+5uR1Exujq
2VI+YCAo+rti+pa4oxW/DRmTCp2DN8MgozJpGwpPp8gKFazUQrwlDXexbJpkt0aL
kCmfPGWk28sFu7qHrhsxnQi0ojtNDyehtxHGOos5nCcmNmE+KGdZJ5ABwjHMXFUF
y0nPsbUh7ZihHnpshp3B92g2TfHr548FYmWnb6ahqH5ve9g6dgZLeA8SLq2otj58
uUsit4+9m5IMVCN1SpZE0ZmZxuxzRSd7zo0k7tzjIo7mSGERGomSVQIDER6lQvTM
dG9NWFWeHUMvnIaXr5+iMqFtNkRddZiJI6fVMa9PsHMCKgFXOuF5rWqpEDx8llDs
9xurdhV3dgz8H4yAeELOTLS25ccmRTpnMxQXj4zQJv7fJVaV1zRqZPNXd2FOcvYg
OP2raN+WSEMBRLOT4a1MKK3+u1NuI8LkFub3BJpiXHv7XeUDU6CpPE6Fk23s7gVw
+vy5/1taa2b5YTNHjPPhTQr4JX/DY6JZ5drS+Pg4ixIb+oIgIK6bIU26LWp8BnBg
MtV9Id0LKG+8qrP6GE+i2//c7BBlAehIVQK362SQCfvrCcOViwqMbhdnWvvRfJ+i
DFr0vq4LD32z82w8260/aMn1uryqNzX+buBELMiDm9hs68gtFZ/mAXtjKyhf6qQl
n22CldTqmsbi7KRjJ7bO4Mkkdj7/4sjmHuXNEi85ioZdUpvv+Ev7Ke9maQO2HCCV
2zDkLpWLitisD+QtPAtFDqWSDLKuEQQ4Ef7Psyl9DHmT4lXZN3sCu4dwMw06Vge2
fzO6Dr3RaFkB42j3QJG0SQrQvuv/Zdt0XNPTWplijMKkYOzMKePtSEPPAjMPlEzI
n440AtqNxXi+k3tlluNPDG49ojSbZ9G5SLDd0usMP8DIgP8dYPv7lGg2HlI2kz6k
0bCc4rgMO4+OE7oGDtPn2kvvJV4kgB9uNTnfvKXh7qPtQvr4Et/7a2iLeWGF1SKV
9JdLsliqohIem4M4rm+M0mRrrjb/0xp+2N/AaVH2YnPkblTaNB4WMFLp3opm+PC4
WBAIkuo7NNRq7l+gDsEzMHRh1s/yfJvHNWyUwGA9tQ0zRQd+NVgrwoLDEflTFNZv
sUDIn8nAOTU9IlMN9DN7PlNUev77VLdVHKowlDHft3LktUIM5ueTxBkJ4kT/iZD+
81E+kVwGWnWkNkvb0tD2JrDN+754EIydWiLusorojBV8/Grk6NMFr3j3FDP83H0l
yYGBSDqkIM2gXMeFVMFgnWXkSJy85wJj2HgdqWr++NRa/eUbk1oiy2c+lAUqsi4V
GQ9ApyJcI0IIoh4qu0CPILdrS/msByo0ubP+SG3N5gW3q96nZofh+obxP3P7zI9T
ugI+hSZWqMEiFiDGof7GpyCIsL64B953JHnHkl63PgvUcWQ0F09CuMfLf8qjukRw
kuuYTAKWsPkVDpI6IMW6m68V45kJNPiAb73srwgBLKtT1BkmiF/n/Yw+nRicf/zI
hOT99Ov/2no+XqoyCPAU/3x9ixY8FZhFrKkWaziVdRhB71Y85D8Lki0ZgkckgwXD
W/uLNthg6zYQcnWH2YVAiBkqO7ZfJKrJNf+uEk+owMvOJvn1BdYnBkLeqZE6j1fp
L9YjUnLZsheU9i+9Ib+lGjTbES8X4c93Dj26no8reIV72xhEQrdI/ai5zBLU/Tjj
gYC8QAcYqrFJ6k8e4dmOsnVXwk5jR5+TcSLLBy+5aymnPbten77n4QRoPh2Kj9zl
FaF34fl+A9LDVBDDrHqHv3/Y+ydUm+Yvpug4psBx1lEqWPN67wt6kalYbZk5QsNM
d8acsIHB/kfRvn01eTKjkGuLEV6swz7DHVWD/o8IVc3Gf1g96q9KYLpnvqLX4o0M
BOHGG+nAK58bKX1A8UN43C97FPf6ipMWkQpctLVIUiRXpaU62UdZyccTVnzkuhIM
fNLd1aoPKRYYmTvDgFoupc8gGOtdnuNuZ1+Fabc/FUOz6hBnheontBczg/qQyI9C
ZyIM30Xcq0jcAHGm8ZZ6uNTTjjqQzNj9ZELxojivYGvVtNJYE70opu1eGN9XU+TL
/tBDk70YLierCxnAWF5q6gXvLGMh94GaZTxiIOCspJjMDxbejFWJDDPU9cbbv3l4
XE21wDzekLLweS67tJGrc2GO7LvuenmOhdxU9SolwZpUy+iYpeIilOGHCooIxCx2
j6+xo4IRAZkOzhTclXO50Ka8/RGbwV7oetVDKAOqq+XuZQkJXnOhbWhp2b8PFHZN
s5rQrVKt3JP2mIpyXvaHEcH9ZKytn9lgYnuxkwz6Jybmae2AMf86lYTiFiSKRV2y
/vAo8/noubm7aYpFL8EG97n1iCkvkmUU5EaeeMPRGG9rtpepa2rwdN2m88CO64NN
wtKcFnqTRLKDwMsZIlohDin8bz73sV/qBoPFRjk6jH17u4ri/rTAYC9TKLV6+rnW
DrZmpMohuxe4AULaw0WilQYHtM84c/4gmys8sxLjgce/X3s+tSGM4ZVvEvgRHnAN
PWegtmwqp/PHxinqHkCmnj4At/bG0PHBVRqNAvpMK37HJy902dJaMCyk8TaFtjmO
/bkUlarx+98WhE4kXMkOTBBCuW8gVHtDKVdlZhdZylQaZLVUvfmNJd6nDTjgQk3P
Sus9q0MktSZu/N/uS5ZepCpF35yyUdU7LIEmK5CI6psrxlbF2EGU4uzHykWnFjXd
q0EFTDGnJVGqC34IP0Eg3gPNspOwL/sySyDBBO73RkMndzrva0XaCdNGbvKh66sk
7KX+tpoN/Nf4lR3zeff2U1THe+uGwiDKXhjGroXCh79aeczI5BkFmWaKpqlaEWFd
c3yxx9vhD94XrCj0NE/QUP6pinEJJb454B+T3aMC/PQxAUaj44b4cdLAvitnxC59
TVrcg7uXLCR/nNKYZGWBd/wU8PdA4IU+2ygSHMDzqTpHGydNXrUoCQ/ZYgF/SP5/
1IItjx0VK44d6XfhR7b78Gmx8Q78XoK4pbatDakSRH1IfqdaK/nML8+UH6Yy0eRr
du49qyldaVQUwRUhhHud+1OjTMLNlUvmIY9ot0ZvVlwqlQnfhboRZXpd9OksjAGO
/RkDreBaHAQpphiOqaPFE4Ldl0B+WV6h75dPoFe7UjydUeEYUNtqhuxB38qveHwJ
Csug7d8oooarXzVoWVHGNqQl1/sszCidoKilJIUIrG2sZyOQTKOsZp+1rK+xUfzM
4d+jlrLDwaTbQGZ5RcpSYnZdLpvG1P+jqaHrFfpypzMoWgvGyLBZDB1qx0Inq8CQ
kHQgM6FLp0DF0vj1MUK2MeMVUdDgmx9LgIv7yyOJhgiYbYDmfSuUZPxH8Zhc2U03
4VPwyzXaPCIHDyD4lwPoPiEs1Zut6K7+YxLFp1tmzBVFUQYWdlEGprslvsiDTqi9
nBUJ+ivpyAJYqPzqUlXuNPaQTIfNFVTf3e8ROpID6OpC5gwiBG8a/LlFwXYcunrY
Q2w8jrRnH0bxbebBF50rWWw+Z5XmBajLzOvu81RI5IhThz2mr4oSp0z6IlELjihf
HQnl3pnOZDdJQQ7Aqc6p46XBqh5tTBm/FDmQZvibbpMth2tDMv0sP49SBoaWQ6/y
FmrECytHHoodr1Wt8DdEuaNuGsWf19oW0a2kzcOQ4OzEr/b42q5E8KoqRTmkdjab
wA7txk4gY6Srfb16i9e6AFmSBe7WikOBwSYVFCZunmevtUIn/m28uthlwooMoe60
LERpSvHTyO2ApKxDHhEhg8I+jStpjeR/EGMA4hRNkN73XovnmTxWqFGc+VYuBrFV
Vn2WzLeMiRY40WuK5WqxNoyOz/io/Jq04vWgGsTRjIH5bwuup5UthqWZy6zFUKYo
kltHamksglyFeoHXPmErxijBhHNHl+MU+e4zskiguPW0c4iduqs+EhVk32LCcORh
nAg98GBcGc9s94kD69UTdqqIccjdAAd+RnjzJnxfP3iLPamPcTq5bsqeB1w6H2bw
mHM37eCLkNwvaplvWuE4Lkq0caDmKTPRXjFE1/wZ1aSGVSTgA/o9UPCfY1XCrAy3
MyfCOrq0Pd1Uvwa5XbXgh6lnYXGXCMSxlsconAnH+DEc8Y3wVGtB7bsC7L/go1bI
DB5DIKpaeSw1kZMsUxonNytogH4LxW+7AshB3NDxBchxcCKD1zSbqjStihAAHiW3
o/ywT0y5lt+/SGG/Mx+I4/kCA2KIKtOb56KlKdCnsX+aqoisZGEPJdP2LuDm7btv
RZWV7PPCEA9bH6lMZZexNVyM2eNXBHME0Ews5IPOOzsK8JjdC4DSLFMz0DduUFsx
Y1irUGJllLg54kIb42qJG+VuqVqjPZd23236N11aQZR6rJG6q4mSYykUHcPQ0FBa
VGGdzqzPfFxBUDPAhTUJe22ONM1zRiwIIpLh4UtU4v3v6SCsxIYN6YRuki7sM0TX
GHSDqTa9QaV4a2l4o/Z6zOlFUIS/WI+yZC/zUnpki7pPzykli03/iTfoPSSeplMH
KH40XRanETezgsxArnOcG9ucQTd8VCUFbigsHvM2e9tY9U5ZLOuFLzL1gMXnZ6Do
/h4H9+bowvyqF5H0nWsKjIElGXGPE2dcBQlbcMUh9YPy6hAA4lWJ2mWyB9KtxSmL
ukM8JSbEn028xldHEFYyyaXx9wP4mFkJHRLNl0j0qLX+ETqZE8JGBFinbTn988he
ByQlHDIpmB4mcYc2ZBeaBrNoF35OMtW6TJ5+D0UsqYQCmt7WuX1NFObja6ZNJPbo
btTeSq1p4Ss4UIn/ikPZO/F5DaqZAAT8RSRLi7yKeRSFtUVriPq3+SjBgswzr/3L
W7MbjWXq78ILutBSRMoqmxzDciauQVj9PFT5xAmrf6ptbGgBe3JTI15r89Db3k48
CanhZzg4gNIuFgRSDIoWtinKlvz2mEUuK6USv9EG0F5DFhIaE/TxTY9RaAC2PdWb
sHcGA+28I9+VPwUxFW/SbddmIttyBDUQZjWor+2NB/1Odb3hRl+Nn54i181sXcA9
TPIPELiqIF6uJwaw45CWNkv8uvy0WvriaP3G/gVenKW/953WSo7OrFM0Hzrj6wKC
jGlENqrU0Zr2YTWlGO/+nP1Rn5DIbXNxZwh8X2NbNTw9nAbF6PH91taDBcrRkHdt
dylkVuGuneLyGqkSJ5SDDXi0Z8W79zdCDbVz2uYJnAAQj8pXgFZEZhUu8qId/ony
T/BXJ8XXuhEhxBL0m/mIxn5hSx+6wGxtxs+xkKMEIt6BXJSrTyNRQTIEEOKqPve/
28Q6aRFZcNR/LLkGCDKKAdlyIAQbihPNIES73UUjTYR1+fIsgDayw2URdGCXMDFS
iLrfXYcMYHm32voKjEccg9/Nc2TiSlPQvNChTsiYNrOxTvQrlUUKXG2PFUo2b7NN
oU0n4c+tf1Q7LTZMT0fTWFZa8+dD0vMV+FeX2gJfoMutSxabK176kAmDST3eMBo8
VeiA+O5BD1IEAYLX4bom+QrvzHW6SuQYZifaDQgCd7OxHaKtaVZ72l/cGClCMdzg
8Gk+qiTh0wx+sf0QK3Rti0BvcLDCet6U8WKyKObV3vhsgZauZ3x3pSJJeBcn4JbY
us4hYet/qppGE4j/8lR0sewEduT+8gfa1kRR5PFpl6QY6eK1ZhGTml0TkJJoYSZT
Ilc5lLuS/QGFJEXgIp2E03NCvTRowzI7lzibE+ekPobfC9mHDTXCK6jrZFKTUdvb
KYYZBLAsYK3sstuX4geOQaw09is2rD1gCBh5iRfhHkc8hNoxFRLWWhPAdauiOoiE
JkfgypGb8gcMdReSCIOtEx1KT9sWCHaaQmKNg4cTnwvIQ5bWAUglasLH+r9tPvFB
p+trOaF6o0CmJbmr/mQIwbfDNbksfoBmgMdB2w60SzGIyng7tUTCCsnn8a1GjYYX
GUQIPx4E41JVGnw/ZAcFs9Ob1ygPv40QUlaL6xG38CSiM/zqAezsaY4hcPRymx7j
ox6TW0L182tjY0yNglKbume1d/UzQSILnaD0MkSj/otn6MvkE4pWh4GSQfzHpKcF
GeA6houwp/dYqRMMqCsc6SdGEP9I3To1F5sxfMKsCyCQLi1ff53Nl+4QmiLdDaXI
KxpoGpSbZs9NuI6UuWVhwTDjKHibci89sVY9ph/H7TMPqXB+ovAVHEdufZqtU6/f
2b9YRgV9heJjgUMSYSWRpCxayYvL21yXMHVvHbNEKZnUTHdIrlMOpndY5htIO5jW
L37JgItApvNo2EI5fzMffAuITXKUEe4NDs9m2bNC6vP6GSSWiwktiDhFhtfkaIaP
QmXVAfip0QupGElRXop0+jHPC1snVhR4wjSyoDlDhVRaMSwIsUCbZEtUujFdKjJn
RyRwuiWqnQVtT+9jaa41uIJawwfCfSFUBeneQj1YtC0vpeFcp//zsPx9wNLZa83Z
EpTgNiq4D5h2baeKeHo2fbglhb85iM08qIo2UfME6X4BDFYrx+IASkgA8FTaQvpZ
nxB/PCKukM2Z0i5bubrFUiJ0wPSjWOpdCTgRyWN0P5Z6KvyZA6GQ0g99FRlylRI6
MXFosouzlmaKcwhbhDK6bkEEiEYEL6mg0PAYFDBTsDJh2VllElRiwb4L1boSVVsP
zhjhqnvZ2cVsXb4HKDa/mJmusAM2QzZoj76tp0TeNon+OVhLv/QNFM2MxRD69RrA
1PbrhH3gJI0s6RF5cMBHYlOH8eDcbscRan5VtzGpDcWUeBLmSqbw5MZ9MI5KyQ73
+MHZIkiJEFlZ5xoPMD7X0xzdTMyY7y/WzKaS6hcg8VWwLhL/Kj4h6liorlOoq1Mg
rO1MI76wQWmOFcbKFTyQoFO6h3iEkyRBA5Y3MJff8E0Ly9rhaihQU0pKRsZDHr8m
Fv6Y/BVzll+RTTlegD8fQvznRXdC/EnruxlhkxLfWxR0iKdcdN13315jNHUqYpiH
`protect END_PROTECTED
