`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gw7Op/S5wP1kXjpembXEp2jjvjxelIjqHyFrM9kkNhoY6+zdUHKKp2RU22HNrMkE
UOvJkfbA/HdnQ9JN5xSUt7sXWdyYkKAAYpOc6j16o1fwaQxtKJ7K4MRf3Y1dkgzy
aMO1MxgIcIdnrB0GuRLXn1iLxGqVpBweX157k+VzdBDyDMMjUIvsfQb1eSAaX0ke
K5hR93lAKGSAOlYAZ42zC1Cn4ce3aeM7X0NjLgs8CyysbF3zpgqzdnseHS9+M8mC
bQz66CQyNVVJ3f1d8slz8MR5SMcTVjPnpxmCO1MzESM4J1cWpV/RECAqLyaVO1UK
5+gQxQFKAuWl23bxg0DjEQ==
`protect END_PROTECTED
