`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zjIe9VCuiDDWA+MTsEgGagWGXYtdVazRrlTko0Ww2tq0DADE4hR93RenaCgLwNzi
skGPqmr/g0CWOSubp21btFmAeNB/ldtOVzEyPwvhawq9Kxl8GirsK9ZzgFoLbdoY
fExo3O3bGACV7CIOYzacRLkWcySs5z6VunOAikPGZaO8Q3eH5gtahkQRd29Gnwxa
vSf7eQ9LevEb80sdPTkRxQfA4CAqldQ6IByuvaMGmpryOWvy4Q8pN1dTxOOm/6y7
Ow9oNRrjXebcrMskS4TGhB2gvNEaIppngLyd6NalP04=
`protect END_PROTECTED
