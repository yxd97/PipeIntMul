`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7mjkwZXcfLRv632/60CPNEe/Qzznu93bU13+eihdMCQcMMGIHDNmQFf7jVPAIVS
mtYOBZnUeQd1BQsDVHR889qh+sk6NlFUwMM5jJa/NohCg3tDtka9IY9KNUkn1B4p
/imgiKH0ljKbe+Iaw69SAZDRaPFTQzvEBaXjVbt2WBsjmLUx/GLemjwt5ONQu6a7
gTtRQU6L01P79dOQvyQGLGqJbf8Tnvaih0hDQWefWv5RBFj6y5DxaakB0dMjnOq/
4dpUNQYLaqLdFp7wnKzdKlMBKvOloxn397h2d85KReqYoPppwapJnaf7ZW3cLW/z
59WIp041ArsZE8bsuRX+C+8RAaBjP1D1TV8McERPoIXca2TjnyrTyOaDpbT0r4i3
/yMNgEz/YoxRY6XV/Rs3YV12zHrsaW9a2O9bNEoAP5OMvYxcAft4oTE3HfyW8TtW
NnUVf9V4E4u816e5TzJpfOPCECqfI7sMp0LJU9S9C0AzYzqhgkYrlNaa8cgBg5NU
O0s5frPpJ1GNFqnry/uF4Odpn86hEctx6902/Esdxu5+m45fVU9nlsriqFoY2bix
Z8WhbNPIbo/G4n6z4MrGwg==
`protect END_PROTECTED
