`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0+RlqIoJmJoezwm6ZIcLMGzJcL6X0BBnqe+4sNqfG1POI143BWoi9GNVIIQJqT13
6hhkb29+mDoYOkLKGafuh2IRILztjc7s0dYzuEnhIHmc7SJqTUoKU6t7IxG8+Te1
lZh3KKoe7qVwFku0+r+ek9L8w5YrLmk+PNSQx/j24E4e9UQRdJdTIrndrvNpy4nf
+Hcmv7lL61z2J4oMswjsg+aC60GLd52XGKeZIPXmmMGdnCdBwOmSd9RauBJRTkL3
MuOrohoK/q5ADN+xNoFHpKTM0lzO9IBNd8zxRwKqb5MHqvMA07BsoiawQM8fQ58Y
BXztIO99Cy8xy1YOvAM/oA+2FsLXhMmZx+JwCMAjSt9q03otQB5X3rSIIPMsJPKv
lJnL7cNS10TEt7RgkfeLxsIG7HPJDnz3dU3H3imJgHMGseRagem77PzAPiKUr1cB
AigIxdFzGfkrwr0tM+PvjE9fns78ss6+RG05R31RX8LOM7rKgoWevDamlarVj2YZ
FwhswPsUd4TYfdqUuSWlh2TYWIMONEiiS8UfGU5aOCvNwcK8udgEKVnyihb75BaJ
FcVD9QlonYKkbO/KLnt2ZgG5mkMryJreZ8kdHTdxV28=
`protect END_PROTECTED
