`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHllTIR44BWW6iN8FB694fEsaoaAqJlUzo4ULiTCfp1k7vtGkW+26JHWaR38Ec6m
tGKgpyrG287qxOXIe/v3W4SEZ8DBECthbClv4v5bVeSK2ROjKh6gy5GoKOgBId9d
vj6Filcss26tSZ48Z9Z5PYjTadMRyMgu8aAH6Or0CvSk7iOvhrn6R9YWya1ElU0j
s5GI823D9lzKwndbOi/VJAMwA7ljC+RSO+kLkx5ogRD4R6iYprOQYfLbHWIUzSeB
fBGBXzcCv0qBNuwW/1DUHnZ6mRlAZN2Yo/9S36rXpPhvqXjz6fFqZAUOM2Y6Ufd4
ScffA7z7PBaSC25mV/+w8MUv9wqmWsPB4k38z7qg0Qrr/TsXvOgzbBQtpDP+a9fl
+GGF6z+XeETCarPGtc5lIGZM7W0hKYH9e6V5OoyoMfl4EKZI46asJuN7RggZoN9C
sSVJjhqY6COzl1eJXr7k050uCMV+/0G7I/7ToG/pbjYnp6763dkCp2hlE2rObNzF
uTPwQ28b3Gu+Sr2tkW2dL7uzSy2RWeAD/EQp10m8b/4/HTkf6uKCnoZ5p/z8XATX
rsTL/p2yJwVbnJp2npN8tlZ1COaVzMlQmMnz6dNOjfjfS+rhR8U/ko73AHC0Gnd2
6ykyQ1MTwl4L0DTUJm9lDYExaSotuA1Aj4/EUA+/MA5GRErTUSq8kPbHkSZ3ZEY5
z87yN8uyrInhdoIfjR+0TiC/76/bDu4v5lavmsa8rznzw35qv1fgrtA96tf8DOA1
a+wAb1kpU0hcht+AHSZNp+3Towlosptp9drQMvztclJkcpMALEGM35RlKdRRIX/l
na3jnAKvEHNvKDSvzbx0Q+J+XLHI8DTQilzheDHZdGXF5gVKNVqGM2HT5SLQLMqU
Rx8apUfEOFhyxe29vup/kxPBX6lDpSj3etylmdwEbIM6RpmLEvmDPGSg4O4od+W+
OeqIIDxQgi3n7p9W0K0esDi14iTB/AQk2Kw0QzePhKO/EdblkwnXCeAUHRPiERKa
PaI5PLsb/x+Q684JcVdt1yGz4mz7TKi+wFFg23VfhMEkKkO4dQkc4jzCvtXeLWtz
0LFG6NYX5eUWk6yZW9c6ztlX4diIc/mte3Hk8K5JlAfXHOkKpORr/lRWZpPOcH8y
3frgM874vAMBImUbASophw==
`protect END_PROTECTED
