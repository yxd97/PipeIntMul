`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+LYxrL+L+kVY0NHJJz7WtSI04vZcfC0KT9np647yRCXBVAu6UnNhSkDHtRlhBMo
AH47SUvvxsAPHd2Sx8PUQkU5fGLHPk/RVlx8mcrytOyZ7udnCHqd4Ib3EP0Qo2a5
iU5eJmBNYGOzXO4jdtOI4Dq1OhUguK/ZtHE8tDXNvIum0WTSSwqJKcCqlWkcaK6K
/2ssVx8vNXsUwNi+DPrjD7NEkqetkcUF9bwTGpWY+y/ieBgYhFPHaXAP6BfGUboR
ZrruG7UyNcy4p40nWLAHexzLjGH5oUwh9cQxbiyxSP9gQKUCVqYenci/Jxagu2qh
U5W8YwXRHzWs7+jvC8w0zzJMUJ16N8r+XzXJ8TwbLFYYIt2gmZ264gR9hnZJ4aWo
`protect END_PROTECTED
