`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HQtKYm+qJLedboHE28uWTQ8467Jq2f8PY+4NDj6V8LtSddUbM0Sk2rb3tnX9MK34
8EnaT+DdIetZmRXVpEmGHGx31p8omFs86Mtct2A83ykJT6cZ4AFwHbT3HASnc4ug
nnZ14bkZ+uahiNNw42xQmSBxh2smU3Mad1ThyeO8AURO+PEVifLB+2tViSX2G7I7
teEJBtmiGPG/X/NsmjxH5lDPQn2WThX5M/3N3nMDJqv0eOPR4FIUd4vvAFBoZORs
YtCpk1Vco1OFRob2B3zYCvRKF37wq/mVtyu2lqYBoqRH85XTF7ilfHRa94IN/YL2
F6JtzYlp3srNO55/2cy4c73nct41a+qd/bcWM1w9MtKN0FTkGhBVNKqL39jn0UU/
8VpS9Ws0Om6Atv/2uGURrufTjiKFgo3DxVR9zrg/o4EUFxYoHy3gLfX9DEDvwQ6G
`protect END_PROTECTED
