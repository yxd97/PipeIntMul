`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
je2i2jLbDNIv5koXEorg5GTrMx8t16AVLBNLf9TdXxGh6e8WZcAxy2nI8elcybJ6
Q5iMLRp/zmzc245HUpkNOY9f9VsH2ICusIlmy0Y7GHV67JG0S3hUn+Z7SePFi2uB
NVt5szY0wsZDWTHVul7zIvKvOgn2Zd4KdZ9BlzDygYkoYn0phWJPpgXEpSQRhI7V
ZRqmxfJWha0YzF6WiikLGsyHLbpJeJsfJjwCw3WHY4mJJqvfDileUVNKFNGigs/1
U+Y0Xkrefiu2Zi21hwO8kRcVDsvQl5zR3Co6aoyCUJPKk2vPJRjajLvoTX9LhedX
I0WKFqaZZ3XredcsEKKAuRXAQ+fZMA4+32tB2D+xkH+cdkRGaz6BWyyEXBrBOALv
RIIJnwMfG/Seoa2qB1YpEDR7ECmEbx5oQTcOVQckG6dnezj3B0Ioyi2Ri/XCRd0h
Ev4LezpNCjSQLMxODeFA7Nu5pXMghbUeBRJo6e55OmTWf5h7Hx1RDEi6lfa1uOhD
M3b3lBv6SshgDhx0HtmvRApHP0Kjv4R+MrN12hficr222j3cWQmzxHdEydTiZyPS
8lL2W6JsvwLJf2nn6OwhbIzZc1KxK8WTy56nZ7whrDSCSpeR/HC6BYMjO003N1jg
DqFlZ3j2RjKyfBxQchZfwbK4+3uy2oiO5EnhrxLXLHMAaFnU3UjppstIVytM6SpW
yBtIsb9XbVno/ZK1AhenbtK2FKIdi74p7zXnPfEeYx6M9pGTSFORVcdg+R64Ldv0
uTc3AdUsgyKssYfkHrM8AXmlbAFlG3zDRMzeAsEE+ew7VJmcykLqflTtAUzPWVvV
3cFqCtxrKs/WJnAVBpnOIvh7roK2eGh31oSC/+HllJGA8Cp5A37M4v1lsxXlUn1L
76qLrf82tp/l+JTD/HwKvUqRhtTrMgl2YS440Crc0maYDFOKIc82NhYp/f8d5Ul+
Wtvbe++s37/k7k3Tu75hkbCdUOyobdEyRvuRruHDx3r6TnkHm5+uLcJv8oz2snPQ
qRGa/pEDPmmSi4AUP38NHB8UDi1QfhrIwtpy/I+IVeEdWlbTOWo9r1FPwAzK4sAE
lM8BJdNy8iQhs/tRE9wRtLgq8QjxhqjaMuNQLVFpvtKD0XTPoqdjdWMjT1b4u5Nx
x0YPRl6Te9fxsqoiIVcYpxsu6rSLXTIRUg+OCwc0BsDHxel/UySVlFxcXz1XH52u
yCmfIBfRUqukBD+wmnsTLf6M0aSTWcS/kGx19pUZmqhQCq1uUVyAcV1aF9s63wxx
skueRu3SojhaQmnsqWVmlW3wIrLFfR8CnU8unhypDwmme26qzhk98UW6OKraFWB2
tsDlQqhILygacieU1VuPJHYhbTnWkaQbtVIYJ0qHHXaT5w2nFbfuWzlIZ00eFmef
QZilz07wAp7Y67DZ2qEuQFjgnTZ02MG0+okGo7B6kV/ccDWO6Nq1uaVjKNMWja+s
llAKEGOdNSJt6cP+FjHz+cnTQq5PBPqexCbBumsTyzLpni5xNBXOqmP0TK6emhtq
Np6vvGBCvbwQqgPzIcwORzWkK+cyVqMh4ZiiFWShbEkP3mqjXkgFhJNXgWv9Hixi
QETl06GqL9uMHYbEUga7mCtg+3h1KdHfrNaj3gKfjvKREKd+j2X8McvkLu+BYFUD
ugJrDNY6kp+Elv0ZgZSkchqZJpbM/QAfxTeMvL4kw5+EoHL1HKGu1GFbyhP2cqUu
Cuk3xqhdamVpT3zRdIaO+Xej5jMNU+3PE3R0yYX5voZu4+P6EfCwRs4WJa1ZFT7F
MEYcJleYqZNTVeev4tAaf6FagbsGg/yOQZKWxGPoPapxZEmfbqZUjZqjJL6JahDC
t7UvSW2hPPUoZHFTCxufnUBG6CEFLi36ADkiuAPJhzh4g6PQRdnr6+BSWr+HpwEd
N7Rv4lLcqRlCnLia8A/YQ0MbItHQmcID30KzOMI6A8FIgiLbxkIB/ogw/MrlqgVI
R+fZtwj+e6x/e9s2fsj8BxjFPgxT72HoDgYdxCjhRVatPsR0HCAEBuQBXWPJNRIK
Q6s640gkQWPyCfHM2j8stqEti4VMgybrbKcP/jzYgaOtQCEdBBYuG1z68ISu9IMQ
m9EXoLH6QYlRSYatsCzcg3ilLD7Gx/TJ/+lsSY3NToY1RAcDB3YCO224D4FZdZzQ
C8j0rh1yDXV1waPNIy9MQHdmH/TGfFWYn2LbofLadypfUDGSRBw+mi3UntF+sfv3
Vtc5m/EUJi8u3EqhxLlzfFuLRHseQHooK6JFELg/z3ddXU14q2LF+J8hzGemBlsF
ytC6L2/N2i4NrY0x76zIIRbT67XJ50J3L5kIQ+1muunqFf7ocFKUqMwCncJRtgSL
adVbZZGnw3qgb3KCvDPDJJlCO0IBMlk91FZS6DP4RqVEle8uRYQWMd5nic/LfEsh
9AKM+CugiGPDSp5QsTu1y2CahGDSk02tAfMrGvP28f5Y7TaBYoK0uSJdoY+ho06I
YNGOya5nXKJHyvlCSN44OLjNo1CZB9/SmcCHMrINd2BniXTgHd4s6NfFnW+G4fLt
SgBOWmGvC+SeUH+iWkJX9ACu6e3F46A00OM85jx2aoxmz+Q4eNAAttpfQfq4NxxX
JprQLQbo1MjsdSKCFFKeZZD27lyQP9YlTNCkdjM0RF97XtwvobzJD3aGvM9wJ68H
1laEpu2lDvm8eaHsiDV9Er8Kyb5EjAfX6/aYiswegErUzPfgSLpy5biv4qVNmNLD
3kWZsnoh8KRCSWb2I8uno8+V8EW461y0poK2admg9tZXeruy6T7azKGCPtC8JXqz
AzjSStigi4ot6kZH6gq1d7xybSdbQ+E6aUtZj7s6vFD1GoWvhxvGgTJBWeVPQNLh
B0euhEMuqJUbwUO/OMVV8LKMuPbdNZJCXWBN+qdVL6CGRCVS1RDCJVCucnFdCsX1
Q8tcTxZtxh/tY93DT6Z6JH/u36U71s9t0b6v/TUtMZbTM3O/LPYgVqHX8yevdxOp
lKBwBN09GroaUawQxHWFa/BJhhOxGVllIGWZ4mfrILbtiTkA3yPx5wug5dF4hjzD
NHL9u1V/lRtcGbbveqcO9G+8D4AVQrRTZ4WlXg+rfLBrKkcqjhkaBI/dLZa8qXuz
Uh+lspQvUmfiT42cp/11OBn9OqVwtKpZozoOVRCK773xE5MFPT1IncMCvynCm+sg
K9msOCQfXa31OWDLBI3Oxs0TeChkhC5v9ZYTk/yUuMxrBs62l8cY7CLxakkOJsfF
Kn4p8uE1mJd/AnWVqqv3vDxz8csqbq4g9hfJ55umwBlTY7jTadLBX7a7pJfwmypJ
QOnvVV3DH87zRi6bm75Vaw==
`protect END_PROTECTED
