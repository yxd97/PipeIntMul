`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
112tBpydLKrb/pQNeQkfzIh/Rx0RsoO3+AyUNtIU27HbKjBYlK4ty2zX6tOBXCeU
IuNpc5Qa4X073+katNwVuXyj339cTcUnjVCxO/XuU5b3LlpwHS2zizPlQvsvbxXa
F1mqVBSNU+gcyfzNrA/T7BW4nD0ZlP5MkOf90mxWl1+uW/fhYTc5pIYpBjpmHZ/c
fKFTvlI+kMUOGFqbM3a3iyFFz9kwpb2zV4LmO/4japk2P8aptd//fgeyIts4Yj/3
zJQ1mJ+u8GRjJfbe7pUyTSqhkxp7Aok+36IzP7/rXRteiNQV6leh0yQ144UXOMCO
fqg0IvUFKUg/Tg0aDr3A8WoyKdjy2a2IobuM+u3oFCnPMUK6fn7gyfeiPt9uHfV1
m9X5X5RtQlAIc6Rpbf/4yP5aOYJHohVaYtbkD9cnUB6PCqvKut2U1zcMF0PDBNZ1
B2caILFh2t0NXtdsrrRqwOeyreMEJya7GvT/Li8rKaJtUbuR0eJ+g78k5x9cGGw2
3EKxdxdPsPhFjP2YGlP7Yik66dMfoQ/6hFZFtm8SXrePCsgkFqgx+XMMPwnbPv37
5YZqBaVuFmmIlQHbEfy8Oo7BaKm8wWgepHz/jN1KmYf5O4cckjDFIGcpmvbvnHOU
QZmGKV8CkrGKTfbh3d5r1g6HwJRNAIhuNfY6Di0HFzMF8O1AWQuIOlX5yH3j0QfQ
ONUYh72ZvXz6H4VyA+RgXYTnAWyzqqPHtvbK2wv3oIDjBa8+ww9g2I7bsUBMI5Y3
wJWowLZHEjD73k/pYeAN4nlQ1NqM3lgfXfN6bZ11n1fPnoF7yZ9ggaBVFGaCsUWE
+i/MNh+5dvAWpaCg7M4xEvIixoHNZFpNTRBZFSRkT7/z5hGePg8kwIgs19FOKJr5
IdmOPmq4QGenmy+UkPQkVnNbKvEyVeZANj6vRmVd48I=
`protect END_PROTECTED
