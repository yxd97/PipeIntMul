`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FARGMzN/hRkzyjGSezAMYNotaF0BfVlG8b+ZxeRlyE/uFXGC3hM/Gm7g9EuBD27i
nFp9t3DvjhFu1+rfZO5PiOG068ZAQ4o5wDY/+WZ5kA2awzB0pZNNtwpKCL9VIfjQ
2wwCoJtiydgA8hMi42A7QNJ/EZPYq0LUfrjmlp22yHvJ9KOIsi2QkHMuOuvyt4i4
B6LDzsXi/Ga8UHT2cb7avSAvKJm7BchZy/ypmRGdBxsvqO0wXEfLwmwZkH5dt5VH
hnQY5NqNM5W1oy2P7/3V3P0A1XraFj6qHPgxTh7qBAdPS76OXQIaaijAxH1Tl1nb
nbviBI3Pl8G9jfEZHAK66H/ObJZ10Sk+7vq71THJqsaTUWG1FiDcYFWtzmbPWeVm
b8e9i/Qt62SsDIGtCDMul4aOkV6LKHZM/iTtj1QNl6FBE+ywGRrc/taepXmdRXc6
nX4QPnSRhNzAHIxne3lxy/30ZcMbnyqfJdL6yiy/mDVqM9TH3tBkeFqohwYZwIc1
9fYoa7PhAmMG7eSXBk7vXezQgmIgQ18PwwlfYXvXEP5R1SuN30MheOFfSFyn27T1
0XuXDRZI5Rt1i4QP7GvQl/eNkpnqwA8pR1yM2xTji1kOP1ZBvTu32bN/SaRUmAZj
cieq1t04H1rsf2BVamUWdXWOdiOXRbNNM3DlOFtsKHf8Oot4uFWWKNpJKmpDjoh3
XCEzOnFDG/V3VN+LYsqceZl5g6PpPIEsdnPplnsfW+rAI0apGTlzHtv4bDqJN8kw
Du3sY7BliwIDtvfVTNpK8iDPpXXj/y/QoDj8v0E5B4MePCqSkuxlvsYVNhztEJ4d
l62iXcC+Kazgw0QbVGhEgdrT/lNENBM/hdzX45sMVmpIkKoP2ld2T6qFY7zV5NDz
fIiehK9Hhi2JWWS6FqxuIZP2cior91J0xzcxwkO6jBbpW5lSV7rHTi3++4J0hB9A
dPl4Pw3sfGivzwREU+6MwAWnZBtanEhCSmCy1IkWf4XarJ5Pk+eN18HWBDZCs9Ss
FDgUlmYkAnx37vnXuPUWAZE62v2JQHsp+TdiRZp0RMPlcs8OYK5GfOqBei2pjccn
8Al4a1YY1RVk79NnKLJOGRoEbHs/wK9D7oEGjd1JYUlauB4hEzvn+XfYdDZOx+tl
TgWYyy6cjfoR6FVm9a4fxMe+wWg60LwxNtByMdt5vb8=
`protect END_PROTECTED
