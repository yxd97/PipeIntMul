`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DhSxG+Kmz3UYJQojYM4+aS76tx2IkjihKlJOl92j/3yQ4fnDMfzim9zICeAv0nGW
CZa9ZGtrGhwANCzgIeioSfE1JFYfU7u+mZo9Ue2u2u40nvQUipslt9/1xpBfSPSh
bo23ONiYiNBIMW4Fi41AzlhddklhNY3nNZfZMRIXPtTDq1OxjFl9EHj79+Yvd3+a
K7KGZF0p++FP7rHlB25po/fIuJYYiC8MibzIrxDIp0a/yT+qZr0DzynOPwYwr/+P
KLOBREDRRGoHjy4uzc4nmpQLNnYtdSBo7l/xwrXFkRm8pGim3onfsUtpYju07VDd
3V9JSc+jbYJiOptWO9UQyKHU43eDjIlq4XGTFQlRvHmeW2sAwXvBU2ek5VXBNJTa
+5BvC0f/PJE5j8EXm8tmHA==
`protect END_PROTECTED
