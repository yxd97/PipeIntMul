`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7p5dE7rrg78jEAQKFZ+p/1ok6PjFviYBSw82Q9Kt6bEnBvg1ufy/lBiTqVMPhOgC
sRFTWR64c8RhaY4h2yMAzHQ1flmd7n/l05gPgVTyUK8X3huQNAS4Get3s52Bexv+
kRz/1HhTgqh+rSInJn9Fswul5SV6oZhvwa9DbwhT36TV14G2xAs83tkKYTk8Bc6O
4Ni9T3yYYRdNi6JONuYtyp1YLqGTl/hBoord5PhjZZsNvU6naiWRS4+BTQiddddv
ctr9/+cPFalvVePKz405ukmEVuLM2CnzNbnjEXMQupkYj+3+T/59skH2Qq2Rsl7Z
EQvVh/wvCa2R95oBt/caWDBCiKQm8KuA9yvOgQ3waIFAc04UL3RcMmmPHiQ7p4eG
ma5BMv4yjGrWIwV/RJcPvg==
`protect END_PROTECTED
