`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cPfp5l+gN5cqlxtoMBSzErhY4whz0JX1rnSnQjiQRHjr/skW4i6TFka9nlfWQjdI
hlUGqkTwFBP8ktfTul/PSnVjgd9qfT07kg+iLqDB064f6RWJhPhGM/HFZufukXmg
V8oOJKzfq+L6KdIozg9sDMjc84BV15r6LbHybuf4quRPPvsrwUx/rd4QopUHAi3D
+OWOq8JNH1HtNLinG/WzYEvHGGUyou0/2am4272LZJDzOYn2GUNY5wNLF5SyzrJZ
XZHc8UioSLfr5TW+LghCVQ==
`protect END_PROTECTED
