`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cPEvlvyjNMuIda3L1hqdpRTkuM0Db2zLi5FxfuIxqeU7w08tqM0oi4RTaUS9DDH4
SElsZMeJtxUFRD/FeCE+0e3fWWCUIAW2KW8Z2s8nZNJ8f04+oZIldKeWpW2mTMcq
QMQ+/PSopf3/1LwVVAP2D53rDLjergapd6ENdzzM4cXA76emnWF7yZW5B32rudIC
97lqnqrxft8UOOSBcqzRoRIh5ZBWpQ3stO0/NswhYBf8fxy7pvp3gFn1ywN6UkWQ
GT1tpm72zk5TztxKPAQzBbgNZH90mtOqadXvp2EchgjneYEi1D+6SomzWTqY4Yd5
AfRYlCKPytn+hj+4JZubzjG/auHvh1Ui6qSx8VDY4V5VJuDB7FHzKssj1hQx50ey
hBOBapjMtcjIzR94GQmoa1QFxyrm4WHbAi5hClRe6ag9eksEbFycrX+A6vxaV8R7
fjzhpg0NnAtShA6ILqieT4q8l7uymQFKcwA9Ts1ybXajZOGgpAYSIinfj/+4oxoY
0xtFopvMdgEd+LsuyqANL+WpWZ85HqoZ1Y/Xqjn0voEZB7UFeZfps9kQKFb9m/KO
J4NOaSts1tDMZIsbwCtfYKct6wse8fD2g3x1GFI0Tf0ufM6RF1NbbvSlGSsY588I
MOjbc4Uahv40ZzoDSr87GFXdhitzAT9Xcaxf1+7NTasbdgg/Az86cv6l5CM8RXUR
yzRZant4rP2Ho3cHwCEMvUIyoU0MxWc98hxH4snp5t+ueu++jFS18aUOtUuTOP/B
W9cJBusk7+r5xyW0RqF/+AyTB9eIODixKzGclBJOk46gGRLu0K1GLT5pBCQFg4rk
F4KF7DLa98436VlGcci4HxLetYGMHQatU/2R0UKWuzqt9KuZ9wK/OLxUjyeHtXUT
7EFB6RhHFUSAcwOF71DmfOyggsTNmnh5pXx2OOv9M+UPC16vM+CNfGOp9/Qe8WFI
MpxvYQBo9B8GcWpCc/huZDBXe0SKGCTqCQumhw23V0r0oUf381zAAFvndRsD1X1g
umFtB3L6TLMEAOvm/gDwZMA15RhFLraKe4MV6ppWdF3DE+tmUfyGKVDtF/qEev9m
0L/OOD8VfW2DoUg1KYiNXdo3L3xNRR7cRETYPGUR2VgqQ2dS6sciOeYvyiXdk9lB
NPcmkwmCJnSgFzji5EM+NtTsQAnmp2XmUz8jzqhVz7Nq8ivPiKaibypyYHrUooGa
hWRGN1e6yS7/l9lgV9jZcxOTJRCgsoyw2bsbjlyjyQ05tBHbSrMkc7DMyCwXSMsh
2F9V/RnAgfe4r52fj3v4/4CJTLKX8elcstjnnLlLR/JOn0QsUX7i7RZN4Le6vsGI
M6ZXT5GsRO1kVn3Kz+6ATI8RItvjnYXix15VONRRUjrcneVWP81IB7EfpZxN49y/
bn0ZXZNaCR+b5M3aNbOd/f1qyMWXT4plBM3IgH3HatcxegNcca6ktyxyOZDi+PUV
iiwu0FxnQaGYzl2cAsugoQ1o2ALX+sSmX2/i9mfCXnkwE+atn3gPmhYEvoAE3n6n
69jM+/MO9jC4J+W+LQdi9R2GpejeNUJVEnaULGjBR/hbG5lk6fIsu1YjfO8/xTJ9
qlWdBpXMRrH3VtH+9fZ8osLEcEQPhUWpr0EOX0lQV5Np+XJaITtZ8XZipi5LVnQj
PVfOhzf90sqb+AX7TPRQRW1/kjhBQR9ZNp7ByhX7U5xMnhC9sG6vD8pTn5eF+BxY
ODkhaEfkzorwGWWx3yp5iQj6EPbSpN6IPJ85lySK59yAI/2utHsBhTHmpSNu9xWH
edoZsQSlAyd07IvB7nxGAwdN2Jvq8jAAcuFoCd5JJlIX1eD+3Ho29GkPXV/N5VLy
/5q4JR0ETH2A3X5QOnIHqgXrSqTYippFUH1Iz2qVHuTPvsVPgkvn4J/HfeuTwqCk
iAwnYt38Gsueb8qIfkCN1Z5cYGbbwuN3yAotZtEysy1UT2rQE+RzpHUq5ifMZMaF
Vkpo0y5n2DTDBlwCKbEz7VuIUvIv/9iio0fnb5aa1RwsWE+t4qEDPuOa+59CmTRP
HFVc5j1M24SMlueLUkKSAqyd52+6fFCvTnG14N8Z/GzemQB6rwEnn0JFD2+iMizh
evC+W48mPIr7AQpOTpnGEg/XJNjUCqdIGqpxMbmd3NqRTnQlc4Wrp6uOnEUz20Qq
0W7LlevT99r6x5ppa2DO5XaB9hLElXDzyf3rzUcyYl9wG/tOy0G5QRxdkKzL17Gi
sKYBl6Thpb/6/0uADQQ1dAqFPEle9JfjveTC/yZzd1plI98A7MZy08hJCLHUajqn
/FsWVjYRqjaqppGI7zHyl5tJmI2Zxj+ERIyswlGDmD6M7aroSMHVBHZh/tbyStky
bEC5uY279qZOCBj2+Khr6SKL+77LTjagn3qT4ocZzK5y6iJXQIvVwF2r0Dgo6kCw
2yO24YT97U7/sWSupKJk/FVLR5QJQFelYRKKVB8AFIz4cdyYJlOWeYmq8Dc9rJ0O
geRc6mhkelVynj1czwz2w8bDfsuT+ECtsyusMTZZMEkGHOB5Cu8JiLbSKke/u9k/
fK2Trg0nGj16oGRXTOpsxlZXO7hlG7RXkPNoEbD6AIVkFRl3qNPUe//ZVty50cIL
DKV+jC96NJmD454J88R8qf+N5zVFK9EIxsFCJlkPSFwm/iyasdmpx454wxUd7kqP
REFNCvdjJ4i5Zg2kBFS3Hn/rbH12derLDFlRSCd57reSd+T//pcb3c8L8bGHWhbu
pvOs3+1uLMpo51V21/ZSdt09ivNDmZJTilQF3HHtVlcnN6jRgGFOsM8COwyWRI68
q4RBIVnpd9s4CeroG3CoMc6EWAzY8Lcn01OFjkmA8ieMJ8UBsnoBCUVuLQnVPD98
jFjyq5t7fwgrXdk/r9wCdNxngv64dvvLE6AuaAWrACig8IelN9brKqzMOitunF5E
tFhxw810jkizW8hlaMMj+9c0nGjgkPrcfAWt+SOG7BZAIFQiYom/xqATXb+8hInw
tg/MfIG3/cAvHTCV1lBA1n762tSMD/TqxXO9subvvvV5R3+q0AJ8c2iRvBJEz7vy
RNBdoKuDMInZiqnggAmrYYEthBSp0UQX6viiqkl6T9JwPGqO/OTgcRe6e/LUBrhF
oc0antJRiakYGmXyh5paccvTfhIs7MeXSi30Eq957bN62Jtd1aVoKwDH66995cL8
1kNYBzn8LM7m87xy1kI6VBjvYExqApQ93HeSpwdJnqE4zljcXW3Jf+79Pawzco+/
bB/KRdec63PndzAsBxvB3UT71+AgLC30QPE+tfQNH6n7En/v8u82zGE3PU5irww+
ou/PELb9qdX5TL85Us7kPfC4nJH8Nk0xe1xf4QZ5OYheSsWZxJdUGwFjN7/aSGNa
NKU+F7nWxV6O0I1IWabojniyRraiAclTY5JGr7m4LxkMZzzRMCofKL05RYeBX93u
xScumSFCdPey5bT+BTA4dn9w/SVNE2Q4cwQMgYzFeSTmJQJNx2tLb/M0+2jdvK7P
zM/VAjGRx1IlD/tNiHfLetQAUtXhbuHXcmwbm3PB0vWPjZZ/GKTR3wuU29/Iwh5J
FzK4Mudc4e7QkqHD1R9CJTAydo9iMwZUlfPr/W/sW/xgi+jNnVAKC0a7PKsjqYn5
e6phzq7kW1O6vQd2nreQpZ9nVWqnosNnzHhaQqh6L1r1ph4vjHceHUvUQzhqW/QV
IlYRnmQyYBfIKZW89XWD6SNjIqubbsaILo5cpayf6pFjTAwfJ0ghAAXKpIHyQuB4
UW6nU/Sa8AC02Wu3ThZmN9EnKejzvLI7R+qH0ZT/cdOoomTzNIDDZDISp6ZxDoMa
BWK8j5GrRCoBZtLqFuvnW30Vh3Q7Im2QXrfE+bscV2FBMPbDCnxWxV7pJ/bkSh//
Ta1/QkbYAnZlT9w8W9EP9PyOHzF9VIZxn8uQ32DofVBN7ZI7k7ZWzG3oEfRmct0C
`protect END_PROTECTED
