`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3gWv66nlBSW6IIL7oFq1CWjCWe0o1uodekYoq2mlNMlxEY5doEVwFb1bnVCZ9SJl
O4eefL4+WmuftGx6eDrTHE7+c6zCiX187Lg6f4le7XPlb/rqjUa9jWTcxaI/aPGo
LeDkJqeOedbnyuNV1YtcTbdQHik/nAhd6vbTT04lOPRaA4dZub9+rf/zGekCp/Ok
adyTGP+ytGSy4h/A9NXtsTCFY8+St7TP0oa2F4OjXwBZhOQkLAj8JbpKFYNDPQOK
VHdqzvQ3MLzFZAJjT4EAqlZTtPRUbWbrUvpP2MGwNE2re9S6TUuS79GqBTxVq9sG
hePwBDjwLAHNt8k/snZVspJelSAPDxb+Psbq1hOSyL3WXXXqT4ZDcOWTsK1UTVo8
Kx8in7sBbL9zQUowGKtDaMZn3fSCl9hXy1IFq8/3/jrw4fLyqEs3yBOYzXyR6gdE
72pYSOWuVsm2qZrdMyuU6TEYUwXIeuNEGm8YI1U4opTg0erBvWe37wwNWUOQwbrg
DI3u5+FRWbVDDUjYDUzNvEbWxE8hmgnD9taKs4MvMTW0tjD6LAI33iaEoArBKK2Y
gN+CqfdN4vJYvJjz/My70/VsCyNhMPlf/SZ62zKqOV7uVUUQn0QAgJHxlq59k/Hl
+p0GBHrqarvapSU4GNJdG/ILyCZ/beojWEAsyRuFYKf/moIMO/fG7b2+MQL3KZEJ
Q6l8CPMpYHla9ua2sV7LJHzA2Oafe2J3C8xIugq6DwwnLArdIzJJTXX6KQFmgRo8
9PyzyH6RRp+Kv4i9dUS231/KBwJVzP+X8kd87HMCMr653OFqsZUihUZVEx1olyhQ
9TM8KYbFYHBDtW1iK9gSUS+g1jUnUQZdXSBU2LXKYois9qptFfdE0suj77GLPH2O
jaDy3uffww3ft8y7YfbqPhUx1khMEc+OU/h7X7WQvKMx8xFepfXGFbt/lkEeJhCm
/R54BUT2r2G0YO8ASxJOFKHKrWG9zjfyRUhTM4cTbNin980CqPGrsEssOK71DfbC
ZFOE0sCcCRloMp/Xx3EWqA==
`protect END_PROTECTED
