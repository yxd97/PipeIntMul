`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DF6A9EyhHm7gk2grZ7Bi7av59MFMGdKM+oQuuECf/8Up7USFOK70Mzx+fqgXdWzX
h2/zQPVwqcJG2VgjUl5miKsLHlDuTnwriAY3aS5DhiAuRy1d7SulJn7f+J7XMNEh
QaA+RQMCmZ71WorL8pujo0bQzFZ1zyrqVE992xaxIoyKEU217qGSlSZAy5v3YJMk
x3/y1USyQ6sbPnpxFXGxKETDx2UJrSfJr+7v4B2tiR3ctvlA2yzkJq6pwf3qp+Vi
emaqdIPeIMhkld9d+5oubFPRhSnwaVRNXyjVVycM1arCUcDtOB3DNCVk6QJVX7YD
oH1uwGo1uS10x5YtOlqcKMpsgl0jvnFU4D5LsKr4D7e14KA63LlyKPjeskKOkJSE
mIJDPkNA97+5dbnZLbcb3XadupofOkYmmttKr3tRD0f9/BqV+r1VddjX+kompt87
LGP38sKpOlAN0dg1a5Hosw==
`protect END_PROTECTED
