`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
at6zwK44y4w4LXaYhVjm28PRGvKeoXGch2vJEj0UwUeRSMHFtOA2CuFsN2/WzgYU
sHLgxbTkSyNamN/kqxUYeYJWPb+5s8pr91U/vY+f8ajCLJ7/t1ukctGXCEzhNlQb
AaK3xXbD18TyArIjSm+Wvb7kMMFOTZl5av7yt5Ynz4WOmSl+o4N/t8yZ5ibRMOhg
4f2DWAG5y/6JQseFHOceu5QRztFkbkMj4qr6k6Zu4kPyc9Yj6eES/V9RwWUA0uj/
zveM914SevEKieEFCTtnud9ZZFGaBe98jQ9UgBCdULqfhLehYsCegsFBN8xYIQjj
AatyEM4h9shJyx+J1clbDliD4rtC9xaWU52pr/i6G+Hdb+P///swMX/Z1k+JFzsJ
G4MvK0fKtigY9lZeElpDRCryrsZkFp/FtveDEVIvUMfTzNWEOrCZH18QGU2vkY95
pbFBw0q/6Ig6Mi6sQNKEvbh2aem+xTEJ/S6yL69diuyRAdAXLwlMH2V9Mt4sIsRg
7Od0V6vRWQf1KpBi9369lV70aXGBOiYODE6CRp59xQjng+5PcUO9IBApGxA9k0mp
9VLgZFlkTMojze8dprCMwJVlrUDZzDmmuw6wjDt1QnCQs+DcxTM7fF/a4OizBO2n
mluDBexv55soeLZjNZilw4Q2wJznr84PR+f7S+H3tVvMlh0Qc5SUusplveI39DGL
rUTFecXp2IzRfzvJOvG4RY7d7bJctJKrd/zZ9GLEMbWSZ7PcKNyF2zYfSCps7lcE
tagpyWCCvn/oBOnlqtaZm+q6rgqbqhJxs55iHAaOgyQMX7mLcWKXjTX5n3ukl6nz
ZoX2icGZl1OeJi96RPrjhtVQEefZChbbxwMqy/LnTjsRj1zix9RMYGmZE74HLrWn
TxH+xbyXyBREp4xizOF8OVRiRaQ5edVv2S+5vFnL5eiTOk6ZYkPfDmS34WJ6XtLq
PcErFC53thyA1IztMGKRgQ==
`protect END_PROTECTED
