`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9pbhZkQoknd72f1+1/Cq8p4Jcp004+S41dghVz/Ufz+WCfKHix6uDKCP1QtwlRV
HptXAjLfBHL4RiOpqQy8PinN7B95wctckGw6HHcx/UkV7Qj55IfWeyQtMY2xOwqC
GDsFjZjTjfs5WFBKKsiO9LLX06zET+97wjUHlt8BVcEfpEkQoOZnPDfT8uKbBebq
J/TzpZ8P9ze68cWUYxQJX5m+HR+P97hM2CggcZdey5pbxwrn1HUp3YPsJIcwzR0p
0W3ZdxCd3Cfy4qWVeRdpb0UEGUC8KDsZRsxyjPDhEhVC4TA9BiNC1+dtfr5aeS7P
nfMNdrjxKWswiY7WVElb1bwNCBQyXd0ClEO+94WiL+YKZXrqUT7BGHMjxd3r6fLu
R4JbdObgr6xTxooJeON73t/Bif7eQCvqQj1DpX0+GLRWl7ROPXvNjwIlCgpQl22f
II0IjQfzNHitWMgD/4t6esg/BILzf3MnQiNpm2nC+7leD2fvG8sV69eICdkYL+Ew
hIM1fkEhhqA0I0Z7ZcHT3nEQ7+hM2xyu4eS0XosXYLWwXr8Nqmp3f+pbNCt6j5+h
Qrkf2UoMVNhPefB3dIwJJyBLyZN2UuRxCNpg4AIB80K8i7PF/yHBSFw63CqaaDhO
MMFSaSieqLsIYynalDWxir1T0Re2uFcjeIv5YUtnYDBPouh85v08oS0XLITHDyNG
8GKk/+lNBYnh4dBhtJND4nGsOEOHl5zqVVmynBkNdjZerDz9FXNLLp1UkIAXTEQ6
Q/D6ilVhwuV67Of40O7W0Wzw/zOhMSbU3Z4BG5yNUvf2Zv6oakJQ4OOkJAGeyQjE
yPbpiTUDiTkzkANVdy/BJg==
`protect END_PROTECTED
