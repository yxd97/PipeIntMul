`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qysrqWj5m3+cJfqiZsDULJPcb5vT9sA0RID/sHZQuz0xmmbr7hVGC4MQ1SqV+4c9
Wn9K69wrI9ZfcAehuhNmTlCE4xkFna2zKKc4pjcj2xyQCtkeodO9TVVo+xrLgk7d
INnki9Yk4ZcGwy01Yo1lcUL1mKFg1IdkiBGAafOtf2EVi5HBRvcNEzJlGO1nn0fn
PsjWueDr0t0XAXwcLhUePa+mFw84sVOf9qCPBvyF+x5mcuZuIydHTaZjuBAuOICD
Kt8rY2rNn/0xL2w5+OFfoIBqNJPfh3QyTkJuVBvTdk6yZgc8rFKMnJ/SQXLF+F1x
IPx/i4ixocHpr9WO1ttaBijzB4tVbiIDXTV39QhY0kP6RPAuFT9RGbMKxmoWOYxr
+HQwyUjU5pRvFCCE3mwr0QCADPBxhKEL/RGb0Ghyi7a0AgLWL4fWDC4BqusXaBj8
oKE12BPTXNlFzAjoQD35WfyOPWSNsqty4wMyigPfm2Xa1ynLX7EpnkwXCNBSeAYf
0LOScadHjo4P0E0/YOpoDyBfNwD782I5C0gOXlnrl8lzteWQrIbvfV72c/FGgcx0
iY+FqwDAn0R1ttHemye50dIzV5F1baX4JoaMasKLWj+jUI2xVBBKoYDeWfdtS7dF
YzBwSHPmJax1Ihqzy+hILQ==
`protect END_PROTECTED
