`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k2y9etRYpwM5Ad3GD0R44T2ZOrjwW8pn9IIQNBSJWVZq+GXNSZK9OyVqRkUT+Bvc
xW2CvXk91RWg6dDngyQlvdMh9W4a8otkIbFEeIMqw35ypwC4hRoT+GurJYge+vSl
5Jvmm+DprA6BViD6nGq8PIrnG+THrfgAkT6d8lxqI24HgAkGEJPqit7NWOGKdyE+
mjM+2t9EPTv0Km2AD+0hNwdKm/0+ZSNfufUGCmCfDD6uTc1/+XUs8k9RWLkVVENH
xOHtVgXgLG4qCP9+eKVAr387W0Pvkh5OKU4ODFSUkUDdQOMCfL4flx45uEOTM14f
JIR1Rebkr3cHDVLHjBVPf5GKh/lh9nC3S+HK3gmUO+M=
`protect END_PROTECTED
