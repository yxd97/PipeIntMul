`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXUR2ojf0aJXFYL1l5Ew/SD6jHTAK9fcnRQdttZ1VpVJySo+3+XrPLDhHGYQIVw7
WTZofLlJ3+xnJ6zrL3iUg3bn166kcdSCXWsuFt3uVyC60R7ToPsBZs2vhIPzZf8F
EMyXz2kcOiaD+vmMrYyfywXuo4rvLf7VFpoLX8fLb/ZtF9wgNjLYOSVl6K+jLHF3
ovPm/XIs+fG3n8PJLhiEYs1L/xadWWRUSn6ZxxKtPUTXfU8JC4eQflYvQPIyD9dC
s/aAArBrZpAQFF60iW2/BI/HZK3ni1GqRC1I/y/Zec3w2xokoddoLCRIYlF3HFB3
Xb9wTdifbY4oERAmokL/n6rnkwJtba3NAvSUZstgWDR51X+cVvhDU9n37WplR+4p
FRFEUmEFRXWtKPhXKJn5EMcD9hj4eQRUKh7ixwUopXU=
`protect END_PROTECTED
