`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QPhjdYbDqQaWg48GP7DLSsto83/XtQpO5bfLOT+/GS3guhdUV/lBzaNSB6m1EnJx
gTZf8jMLOF0wWwPxe60aN62cxEMiz5+dABJTOU0IKh6swUUbdLGJQNa4zetVHbFd
78gdR6mQK66NdE0g8Ll4E9bmnFxqB5dsB/nBazBfB55fpS8F7sbpjyagP1BuqM81
6Yu2+RMHFK2HmLB/6+4QiqbYwIqP9OxqjDiBOm3I3RjmPMrp5+pntsbVAf0V+vhG
bYWRWNWOChAZxIDQaYBwC5fKPe4/vIhpX3zFNRRNpFwmJ0YwNzpxAO0AopELqvgN
U+ki1bTQOXLLPCcUVxvW6H17c0sXJ8/2m02FDoxzbogOEyVAEmgTs0Rv7G8UEnZi
T8RXURla84w+WzoUQP12XYAM6fpXqS0nxB+3sDXyaVahHnmYlJf/0ynJ+EakNMsM
TGp37B6b8YmbAaB9TNEi5BohdRuXNm+Ys+RyXTowYiTCE1PmlRmYSaOhguPvYvct
bX7Re0hthRssXl8IzyHJJphpxDj47oqJFfTn9/OVUO/a9GcsccjK3e5kh5BXZHHf
gA61cYvmI3Sm3TMaU/BESym8btxECrPl1C7rBHnw4x7d3p+m/5IEP608lvMLsX+q
Bgq9545UeLNOD2vs8zzyV5seWzO8AB0SVmUJ8qGLrCAlEKbUEWlfvrghMa+SEzyc
b5CykHuFxzOwKP0Zc6ConHHaVfWG8cPQJQY9r5Z/jOzP/OMornSCpfLIdyx8/WLu
6iX8d3om//Rn3x43LQutuKEvIoIoBBKOGlZytFDMA4XQZd6ErGj7WJ5EvXIvfFXE
7sh3Py2MulFfQRc1mfF/KP7d95M+63VXbu+K6gPYFub2mWA4q1q9PKztmQrTTGi6
V/F19HTXfQ7iyG0inUjGEl6WIEuAcyppZByiGw1/JQVWHf8UznkVQaqeSGHT4nkj
REH6MozOIljt25c3RrJQMe/hNgMqEUWWH3Pnlg/vRVypbkQaXN1uPweYFYqmm9oI
XSDCI3Ab5MfrP87DU+UEDu9PVpmYzI7zbrF1PG3Su8d0E0un0/zyMHl4qw/ONunO
h81ieTMsA1nIstWm+svO2HNqqO0DdqkRXxbY8SLNdhx/0CKA2qRz6mLAmCM2LFG4
V6Okt671TklV9FyW+NjV3FQbETM3rHL/9sENEgUqD+6EEV1JNYhTZ161XyiEGb0/
7+Edro5hfrz86HpvDLLGAdc0pkBNcV904qBPi+41xsPFfF3Jrssg9D56mt/mT9Eb
6Ug7aqFRsNdA6NayqLsfOB41zsmkgjHVPFAAvq5g/GLetSNVPodWMXmKETRXUOhB
nvydVScRiS6T+7r1KZsEUnteLDdhEelnOV5gsLfYhmwrW83Wj1xK+weI9qpTljc/
6XO6PSu7VfNN8wTJ1xZWlTaRZaSc8Zl4kYaJqBYVTEPVIjMU4a/2X+QX7KGibJcH
VEyCdWqb9UbJ+C/wwey5Ty//yPtUhbsApoBlnyu6c83FDR/ocQ64Wghr74eplWFq
iVrZJQJu46gi1kBbtbqGCjcPUx0oHtgSKmXCvPT0rjvTp0JpK6LYPkK5sGc6vfo5
0AQ63uplWxz4M8NsSZzXEIyV1+6xMlYtnoz/rJp84sVmJWqvJwIT3ZvigAIeLr6x
S5a7eJt0ZfLosnY5OcqpUapqFi35rnfZN3UhifwPsZ2iltajfYZmGksxfRuLRMIH
Am90Ic2pzGTHFX2GrQrXZwDyO6/MvX62abpkPRwKg2V5JwnoL3b7DY3DcDuuWT1A
Xb9wjYIStz6nEPWvfAfEIVy3+p/8sHbxcy9GrZ82lsulrGmrHNy2TZGLXkIE4PG8
Z0pb8SurxiN+KV+Dn7lzu+5XuJJfzndSIZ+7FLSJRp0AW28xA73zinxxJF2nQHao
YSdYRzcsqr5Y+hsmWgINUvLG78PzXNnb4+Fpgk5A8G1hOF4v9auIJ/jBoEUr7ulr
W26E+JCFzHvY7NUHdY4kLtSK9N4XSUNkAtm7SoPf+XOWWGfLYEgysKBj2Pn73bfv
SA7YizFVey2tGspH0RDJSBpsy9CrRVtQM00pPYBlFXdTERs/terR4QRwRh0SQR5x
QgKunIO9gwbhWDi7MSqgmx4wJ6y92ANqRPkoYwRicdw=
`protect END_PROTECTED
