`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M3Bgp4CfSieAcj1melTBokM3Pt/bg1Ja3kCG5O4TiuKJkY2gnxMGbsZZOoVrEdl
URo9ccZaz9TAZYduQOoDd/yXtUMTfPhRJvppZX1DoWZlQcjXgi74XicFRGDe8J/d
HUzSsUX5YkdNzuf+IwDyawXBkEa6AFFoYEEI4ugTSB0aluRyNQK/YsHPp5Kgfcpd
9XlWVWjlrARaaWSOUxySmXvSrQoITDSlS+Zdnz8l+5KRLdWSm6Ua+EaT82nWXr/J
BEOBBVq0eU8VY+xtgks/WMh9Ex/Rylyu8I/HdJ7jHrsBC81v5XCnR+CVZHAAP0vW
cN4+qgQlnPqrgQl2dlFqT/scZqRwzkw31oElrg4AclE7prUMSxUO+HrbzsGfO7OL
nyBa8JD6xn25OMOCxAHIeatLPNX1LSvX2U0ocssL0O2whjmrq1XePCF0Zru8kfbV
LaU0ypijjmsVidUUpEiHJnUi++TDbu5OEqoV5xdHll4=
`protect END_PROTECTED
