`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qqTjoNiUYEDCWzyuFPtF8bAoENe+ZHRnjeHoGrkB5WG0F3v+9D3JkZXGw9pODI6k
EEtFzmN9hOGPC52dKHK15i7IA6YoKCaeErcQVPs7K3RfT1TksaTT5jv5hnb7QxfK
OW8lYd+LlLcId3Q50xCwMekMHEGCVjLpJVyAYkRXdZU5K4kpkycNWyJ+lQgEG0YQ
GJ0XMm0sGNAdkYNAoxDaAHeHgMI0YvJgV7CNLD17CcgYKtmCm6FS9SICVc9Bz8UM
fHyWkbjGAmDLH4UBagxKWByHWF31Dj79Y8an8SxKB1Hh0JwM4lMfPyl8JnzsirWZ
XtQ+KexSaajSHbYCw20iiR0dK3IyFsNwwOQubEfNUykQJxYtevr3CrEbggdua2KR
1GD1YjchSiouTPYbTiJX3nqfCJViLS8phg7reaVc5SLUwYb2MjgBlbDiM9YvihmC
nrQr/RqmUWyCnfPDWj2p1FYDWptAOvsLTkBvMxMRItXjeL/OMoRcHaTbg+abrKF9
g478BtDoMbgi3jizd7FzTLwSUXJQnL1+84VxJSMMBxomoUmCypP/GlNND26iJ4Ak
fPoc1c8qqc7t9cEToep7Vx662n4CTFaKJdKcRUclSElNkpSXEk5OowI0v5WXGif2
Qtsnx+XsXsdXLEFYDsUc7w==
`protect END_PROTECTED
