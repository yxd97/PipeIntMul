`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CeouzJzwftaGc6+02+2mbjjzqnqpqLFB/2bpuj63XYGBDmitjnFCHxXIU/Nxrn7o
i8gvbOPUNhFH0k64v5YG8XCMzxW2keVP8LS3MZvnYKKYNR9Iop6RpOrKY3YYvsM1
UgpnXj7Fcthqr0flyzmx2pG/OlUlVIgwp6BuZRsM1JfX7g5wwNJF+MokkiCEsyfd
gbHCIzefBa/2poge0jwnSkSyBPzzXBchV2y6kCVet7fcHNMEC/dI8Z4rkiBYNgpd
rMt9xWv3J9/VLesiGM6wNQvGT984A9ZewpfrG7NRMdqGrhPMOWWwoV2aR7dWoLbW
jChKdtYrMC2PsYLfh0lBdCEgzu+GoqVlK9sAJd5YYUmRiHe3RXbCHPiO/hjR7PGk
GGB6V8lgM8ZSPVfiz+rlDj0I9yqw9oD4kTroLce3aVve0a1Agy1Pqb93DDEl6QfK
edexMrgIMadFRfyfaSj/zEKfhDu+TsY5YbrXlC1ieoJaOBmU/7qM9FR3k7NpzZfh
R7HTwS/LIA8mhjo+g73Cha/PvRr964eeiIaUPGBAnZB3p+hgCpN0soz/qNM4LApJ
RzL2QFN2PkSvcJ+TIy3YJmwffNkiIA780NkT5R6d1/6ilKL6gXerOgshFQkDODqL
cQFFMO8c5JNd1W1jJnQPpzWQnzbb3m8WjaJccxHWPQjnxC76jfJPAbnu3oMeMJeK
yxwIkegac06zlclLTDH4Ie4GqeNqfVlgobswVVLKcBlSa2xRvyfkxO9KXHLaasRW
CuuRBY6qddJhE5TTRhxTH0JnBodoa5G/b9+JnYgSsVqCUeJ/VeoBZr9fqcutULhz
jplOsEpj8GvJBdKLESK9Iu74/QyrvIfmTCPj4VExq1FZ59YL1GlxWHDq1dDPwRoG
HG53tGzPJ4Fjogv0NzzVuicwOR1/UzO37S4GZIVduvgSY2Yr+SpLi3mwj5lWkUEX
PQuKYa0T2yHOrmyvRENR0t2fn1P2rG2VkILjDeD5vPAoZGiXieCa0G4QCHK0p+rm
NUAQLdhYQ2fgsuuduzgBoVpY/nuSRu4pf1hMNb4s9DrgqW40V8iq+pcHA488sZIB
l2M69rZ5YJhVJyxMZ3QXZ4wp18Px14rzEViso0MCvbM5leTWnKie8Ygh2Gih18ov
BgZAHbXi8CK+gW3VVNzmH+bJzRU/CrEV02h0KRUDC5bI3Xdvs63r92WkMh8J3JG8
91kCJy2wzmfvZV4dIeBL725JTvP672693VaC9zt+yXM=
`protect END_PROTECTED
