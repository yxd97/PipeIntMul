`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rFCaU1Wory3IUHUZVVfYsD1+Ta5KyhtQcWp3pBP6doz4fHVUsS+x6mOqarPpl6kT
CPRiMmuepcvssjURWG5l3q2oAph0RdJV2DJ0zgQyVApTZMGv80JGx443LBegVMki
h/EWFXLbXCtk3TVcMZQWkUuswTeAZOzmL/PDfiLay0ACk/MlTAknJcBC/yMb05ee
1DAtBOAPTF/kvxnT11XAzm01+C7Nsg5QPNiqI3Wsv+uY6KOrymaJJrs/QXHSCIfz
VUrCOgF33G6f+oKLIciHp8YbUN2H2meowW8SfIWZ2PwcDBeYknVhM8wnJt01NEak
RQzM2UKdhk/q9WPcw6ieKi22p1jCG859hqNycQsOrS2Itb+5ZAGsAjti1750VsHL
a0hxa/Mx2GGSAe6Sd1f66/nRDFC5Y1MxU7aiqCNHAUkvX+BuuRr5cTr6YvY7fWyy
DbgKzek8S6xlrftZT0PTdg==
`protect END_PROTECTED
