`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GYTuaZRhzLiYz7iwTaXabC/1MRzZ9sp+TLx0gecKw/x3alj+b2+iPVyow044Y6Nj
vCOqk9UEF+v2KbaTo64neKA+JcLSV2m24vRCsrwKk3Op9PY1AI/o2RFRDu0ZYhVZ
USZfglovmfpEHYwE23kE0El5AG0aMqWn9OG7S93vog0xTSMMyheJ79EXq6E7FdAA
2he7uUa/gUz5ah3QRprtS9Zr4riuBI7Gu06I8kw4ipqFZ/N6EIPjMopyU4QaHgjO
mAknAm400WnWFK3aEnQ45A5UHP8dDYGDhamp3n1d2AuD3BXgU+3NslciMxnBqRVs
nEntrVQ+sWZPFcUtYscwZOCm9/aTFeqQ0rPbp6ot5NwfrT1DsNyS7DZM8H7+/7fD
+ygolba/rfgYpjmMOXZy5GEKfkPwI4grWD9pjlcVN2B2M/+E+OYEZnp8xDxN+m0B
vdJ/dexaanHeZTf0dMrKMqv/RI5M5PaqYOqAMOoW1Up2gIa5wLEWqzD6H1tqyB+K
XMnoJUAPnLkE/LmztboWtozoz5sC/CFOQskY42d1pqj2eVPu1/gF1IdkSHqreoQZ
izfjV7UtDkVGJdeDhZLkblDGOk6WBUXODF+FvdZkcrp9xZ/U+tjWrbfaKEwVL46W
YRCWYZ6JxnTd/kWigC/4CU0SLgW/vogPFrbCMcgU8RVkzwWQKAUKUgmL0KmwWNeC
KVQbXiSWjrTcMsYEsCwE/5q36mzOnn+o3HURB4cszTJrva0RC9vLOCcO0HnVdgnH
A4+CNK47rMNCRKvUDAwbIaiPwE78fkyYEkXWW9RlwEYF4oagnlxKm2bO6VYD1mui
0R96gTuYczn8LfzRI8MTCBCtQt5+cQC0V3A5TdGr4rDdVZMJwUOG14HSPsZC957F
b2Qb4fjImBmJCA3S2qZr5n7lUtoCSTYvXNKtl3IEnUHHq95IMh5wFvBOclNQnYyZ
z5V10ycd+dnCKMVMygGtzty3jg+uirRwcM4Y6SpQPu/ySZXExSSEI6hAGS0Kg19X
yUre+v0F43NbhYYvRBDRyhLIUboloZfUjzfsCM4aEtcYGlf81vA/0faMHhIdoDlI
xHNf658DEjGRme8OfOW5kvTfgzGuee1GaelUmOJyatU=
`protect END_PROTECTED
