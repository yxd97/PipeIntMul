`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78B2uoyfEfM+CypAOjjuZ1S+438O1lKWDQL+uOkbe1AjxLMxnDzK/B+x1HQz4NbR
ly7r4ogXQGcW83qQnoSHyyHBbalU+miX3baKcz9+Olr27AGBL4d3L09L24TtRw4q
6BV/m/SNFaY4PqwEpCo4HSWUdPCSsPCLJVvh/RVyWRsefJsY9/h20rXTi2+2Xhpd
zUifGpT2g4FFZiP3LMMX1WaFrn7qQrm/Q2ivvXdxE65H9sa/Hp8AFbRmJxeVftvy
rpOibERHwEGsTAFppX8Lr4nyrE5OPeuGdQB6q4jvy2jw8ye2LnJgn13gGo/HptI6
Nw/GEHSgIIjuOG3NR+YDbuYyBxPJSd4PphkCT+RO9DUP9176MjKPcA0YzaJjSH1a
s1LrNfbfuC01r/tpVYJp3SwlWkaJxT0PqaC2iZd3jYWDi2P8njIvpqffc8Ov1eYL
Z8gXL5acndkqoNdh2//pppXUZFYezCq5f823kR6pUVPUnc3rfGZcGEDS9lSMKtnS
5525+cKn6EU5cBrr5fx1AM+n+t7sYrbsUDDe4ojWoA6UldnuHDqMrIq8ZhPER4Bz
Yuz6Bicz3+s7sXSUaY/ZhP9UoNztfPDuiaE2a50yKE/5zzC9aBPzfTSU00nGc5bY
5wCR+YVvc4qXcP46xWWGCMRLxnYrqZTj+d0SXy1c4RjH+sacLvYvOB7nwpmGEtTl
XoTuK/bivNL/vBIOUD9D00kA5OdAXb/0BNY4cq7vNKYWlaVeltM3OfkEE6J28I3S
pScoU3U5BPf50fG59434mcKgkF3Wvgp3vHioMXNf9FAQykha9oTLvDBfuzlWgOen
7HSBG9r8/hmYim6OkLiAAyhMCu75p3uYLxGouYCtbA8LwmmN44giidh7kb2f87MY
iJEOjneD+EcRrmBienzTvR44vK51BmNBtRRyWH4zU1QfV6eR/YyW0Thdyn9xKmp6
Dqx9tjr896U02IsPIKgYWGZYrI+EXDmQn4kwflqgOFiO9pZN0s7pebUjD5bu6HlA
9ad0Vcmy1ZPRfORCYwBv99lWaLQ0kZ6wjq8wmna5b9S1KT0bgfOCFdL9uQ/UJpcF
GjGtkAzXObITLz1jnWW9QR4h6y9X/3tfkjKF6hjv1sqDY8eMcfeUh1XVc9sqxaoE
UhOGSc+toD0vsDcNinvpnIa5e2zBNEbynE4T60veBEehVQ6lrUmSgm4obinx2tcW
lc4rHiNy/FbyVvUgVgjbP+7AyoMBGOnSotjGtAyV76DWqgYG9F0T1Qn0/7dR0dPx
NKUCU6cdsVs8+i+/7fD7WxqzqhU0oAVD/dbBQp92SnU4yiSQmmFV4tDfkaYrfkqX
RSd7g+zfsHaJIjv8NF9HYWxSpagOZFDQOoDRg4ZK/t5Zj8gGwcrbfCShdxShrN4W
OS5Yo4cP8Eqr35QCfgSPmw5w/vNC5T5KVrBMrbVPyM0w3JeaoImWYDeN5T2ksxVB
JSzROrHWwEXZdQCrpoHGJDfmriXtL/EF7nYcv6qRnl8a3Nw/rylpg+VwkFOcUSd7
O5ZCXgK7U2vqm6ZtckEVnh0Jr9veHPLyjX3CIIshqdxpYt0cwGreZmg8Gs6kfots
v99PSDv0m/C0BcZnRWzEjOUchd7Z+mX5lFJ5QPNZHMf8UxCLKz/K+mkRafy5PoPy
J4dhFYlhlErYOiQmmbj+hzEB3qML6c4HIHkp/utoSf0UZz5TYhTVxxslZ8RktzSk
t8ZJAgniYcoy9G5sVoeNcrLrW4dLwBC4AjDI/KvO2jtT4Ea1D+FKXHw7ENrLOc4i
nBNi+F/FTvvFGVptIfHf9GW0JMzUzeSA9xpr0xHCt4plnW/SeBUFV54fdnSSqFxw
rmAvD0vSSzWUua0YsvQbDqr3FJFilEcTVorT0RSftEjQVzqajwMuRbM6epct2x+1
WJY1ItoudD3u3t5R3nnaAe+cXhzsmIxEqAFkxBLt37tXa3tED6Ipm1dIa0LrYI8j
Hfoc6zp5Et8V4rnThER+v4fjZAbDl+Jcxls1370EdYP7khvoj8yx8Pofk8aGqILD
8qw17ABGiNpdJFkaY2YjzK0YFjxrRU1PRl1YMAIOUkJdo+5gyXhYPKX7Vhi4k0s1
fkgCZPNRXR1xY/BCktkB6LYBkVFeMo4WpqeONk3u/8o42zYJ80NhWztBJcYzDFcW
ozspjYCUDZHWolTEYBf3gXgUVsXxDdr3b/dvXfGPsYQKC8Vmt8hLDoxXImtU+4Vu
SnC/uIwOqSzPlKLXPKt90RaD/KzYjZ/8U5+kwqNd/uM7zcmbkb2npYv7ew0wGX2v
siPmawdoayNY2ClaY0imVKLpCuD52m+wnyoRBiCi1gCd1ZR9je4ZKDXxXjIlVJWB
mbTwCOwqloS/7vv/IUWbAj6XnWAHHqTPoqxh/Jk5aUCoOoxSgbnzzkMeiT1BATRx
2DIeL7Z5HSlqkBqKGCkUOG0+75mGDZ8lE82MmynG/L+phLffDCGfbMhBCJG+lKO3
OxEVsyStWoXfoIQ5e8PRT4fHcDY+i4+gKgJT5EBjdkJtjIvTsSytNkLDqPi8Ync6
OwSnnkAHlBGTPLBO6BxAXIpTdsGUv4kk3bzev5z2+Hen9kJWMTWTOF/AGVrZGdg9
98yIDkKCXRP4aP6yDSkke1Ik0Qty/N4cwKVbeaC+9NuIaggOBU7vCTAAW/N4UYnJ
wdyt3FGPGg5MRVGEKgt1oemPsC9RSkjIU512o290XUb4EaoWCoIvnOXBlxWtY9WT
hCQkXYNIuVtzfNRG72ZFUReyTVr8tPU508BhgSKOszvLIlT1ipLVNfewf8Aw2zAu
yRjB/kU4n49Iacel+3OwB5rrP53iYKH61Baec5PxRr58YPJh1SEX4YA2kWl6YGdd
V0m7KLSz5lHcxEGOoyJ4K3lYMkXDbuK6CiHsWtHFWPB9tdZEf9Fe2cHivM+JXVU9
uNHK5fSU67YTstWKLWefSuNmrc17tcS5K2dNY76xeR7SrC/ea/2fGzNsihLv3Q9c
XjPiAuL25QYEWxfjhwO27Nyo/3GOXy43UX1Afk6/6vfXWMKen+gQMXRRFZPIMV80
CkTTc6Bl+do2jzTMoLEU3qaDH3JGMYxu9gSMLFA5mzbjRoRLaEor8HrjNn6J4yKq
vkJ/bHtbw43icXMS1AvpBF+0dTQPV+PiFmeUqGutkhsOJK3Mp8xtQV5qC9W9pyjJ
dZhfKAGYRNM3uHJI+JYcvA==
`protect END_PROTECTED
