`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GDLHdq+hc/3khoR30q417OLQSWgLHT23+/v4LR9HqhkMHpSS/idZoSHbXudu08pV
tg0MdfYqNQthi9zRrXyyZl/JKhbwUXs3Pz6YHl/BDTPw2MdrjmM8B+a1SzOErTAy
0w/XYXQ+J70eVMfv8WLFD8t72ojLif2mStGrd21J4KQuy9u+EsPpDjLZ9LiTdZzS
TYSgjHhavzJqs3YQ5AS3x2sqPanFq9wyntwMVNsSnwLEUYhoWrRszKK7FYVAi8Vr
rlpKfyd7hderXi3DF/XOQU6Beh6WNlSLvRrDH3/81rE=
`protect END_PROTECTED
