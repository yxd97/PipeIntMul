`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fg+LSyssJNKapBKcZ6jzbtNqHJdcOIUGxFp6COLHr/YhuBMzFEVuNCxO1uimIDFW
nIdV6wDss7vqaUpCnjaNgtnl8zvBqEKMykznjv3/IRMV36RbKLoH8MeeOisgePq+
mLy4PELDwkgJ+sus6y6QNq96HtUi92StUmY4M5LaWDGwgH0bqBPmFiz+17JXFxiK
jrUGdBhAig6BAEll6jZb8a5yx5du83XNduatEXwbzWZGruOtXzEwjQlUqqi8z7An
3k+dhFbK0FD7ai8x2kDm4wvEL5TziLwAc9wpQqFyUCsjmrEttyhuZW2l13KBv3Vc
zGDaS93czJ3Eb8wbS/5jTSobUMnJtCcERI47CCL73iUxNZOs9WAui64StFs4qKY5
xWLKp5caGUVYFKK/uM8wjEkxxVCijw8wD4IOMmUhYmk=
`protect END_PROTECTED
