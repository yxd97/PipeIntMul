`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+K8xp2u27p1I7KgTxNHo/kEp+9lzoeCdRGM5PnNfNThpxmpD2eXl27DDVOEqWo7Z
imX/9JgTSrZ/AlbIgRPYYe2OqLxxuRrGCeb+AjO82eDzEb2WmqPXjqcoQAP2tfcz
6mYZcQD9XHCuXs3TfVkWig2SmRbuXc2R/bkkLkgwhg1eO+sjOUUQNePyzpKySHWk
kH8DNogpuTqn4nbLP4JS8d4ckMR2/QM2gcAvGv7GbKQEbOHkpIxU1G3Ix+1tnj2d
rLRClwSNVIlExukj/+ExIhP/KHWURXtrDDUnpfAk+OoOI3ix6Il94cjtYeJ2B47w
8r0+fnRbhZcaZWSodPj/hc6ZOGlaLHwcjYZ0rH41U+U=
`protect END_PROTECTED
