`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQyrP0U+1kkBxj1NSCgBolNd0yKFMSO58whSsjtBdFxp5z7bb31ZjLSI3LUEQsAm
tUeERYM/4kc1/Z1gqx7q/sLdRzaQ8RQ6H8LZSkE9yzxGv0yVfdCbYJSLMy2MO71J
TgEqp+VrX4bAZ7cTtcAz7PSl+ovf+9Yi1cByaA1gdD0SRWhErq1dwWAs8kBj9Uem
C8JAD70yBmaotznZtc7ut/l6w+s7leQmH53jnUxVvY9WJJXxT1d+xUlXb/htoRU2
Dyb4hR8mmJMgZTfSeBjkjRl3LnR1Nb4ULXTlnQdBO/G4E8MKb6TV00hL7osHS79Y
`protect END_PROTECTED
