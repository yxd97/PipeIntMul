`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1ibM74xbKNsxc3CtxuaPa7e9U2Px+ZvFjwdwdAd00b2oVr4tfo4yxIohfJdpZkP
I4v1nzCWjj0N/OroT85TqhLRQSH7uu1QrrfA5fSdsHXFPfuPmqYGxNpKnihEohym
tsI0mkj8yru447dVGruGIYgmltWMeHzPz0JK48wAbYWRgXdRSu76HAJaROg8a9+K
jw3fFGFx+SyE5rF5GtMAV7vuZaE58xIep06a7phK1nkUJ1nfo/rNsAM0j7KHmpNs
fOCRAoSmMtAGoCER4FrJr8OVDOlOzNktjzgHDvNE5K3EAV58XAXCWUaR12h5f9Pa
CVAKOXh4IeZZmsueLVIbHOdabA++syCJLvqxcZutm+ds23uYxQi7abKiYAEdwJqn
P7Ycd1bNOTgReIW2bcqYEvQF5CBnV/3/VP4U1LKt17S34VK/upLQbDMtyeCDAlZU
MQKR/yZ4ZGoK0sd7IGsM3Q==
`protect END_PROTECTED
