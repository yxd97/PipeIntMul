`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZDIHFCCGQpiRWDu8Ied+0Ei8X/8Ck1Wm53RL4Gs9fZPdA87hFMky98HeTtHXr4w
p1DIorGQYXZB/YdBt1z9+gw9x4TQgNOL80jTap21dzSGmw4bcQytN6f3to9oA4uF
LsOaZik7fD+OXijCU58Jfk8cNp3ctTii8CtftxDCZaq+woih15SFNhlcjc5cTbo6
WJwe1CbZ/drZX9vSi9uGvzd3Wx7BhoJSKaxl+eaGULPBlq1pUUDn47QPkzou+J5w
0LBqKkGFZ4yuWWtgPsZzR60tYdV8bgHLj/guaj9xpzFMMi+Q5pnT4aLMUPiGlrov
iiPmxZq6b+hsPfhguAzhubtzgCgGfh6B/B9GoflWF1uIpdX8ds385M/S7kolSKV8
k/XGYYg8e1mtjostnaZSPzZEQuMfUdijmwNzTUq9EFT+6uPF5qZMbleAQs7FVK6n
u/beiCcTodn/TwH7vT4m1gsbljpUWexZUEKqhtPNI+6HbuSHzgG30abArkjGY+s+
nCLpbVCqA2BHRQZdy6GgFfTX4AKPE7+pCvhO5w+aCo8j+y5+ZUN6ggMYYQd+R2ST
a9gSBE5obHb3tEVV8z/fbLq12YBZRVue4U0UYTG8NH2dQaKZdPi7A6k0QjuF24JF
UtdBMhvrVoCCp70iFywMMw==
`protect END_PROTECTED
