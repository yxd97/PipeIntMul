`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aQLDW/ypY0OX8+cZceivyfnNyt64pb5QP0XOZLmHzstUuh3bKcDeSY9YZ8l26IvV
n/NzbI0OjKbKWnF60B3Fh0YWzVBX/Ol/ZZJEYyfY3s2KmYhhljWJclsUuQDt1puQ
1niGn2Rd3NMg3W6b43AUzT+d39T7KE9Uc9KsRVyUI1/vnRNc0+I/g5/30ncMkmSU
T7W82LxDM9IwRmz5HivdOLTDWd0PfJcIduzML1uKZ8yM5q1wIQd1ZOxDwao4ecu/
mLBK3i/nQiudd8Y9ldY91vQMZMbordHwESwnMAjnTb7vXPiwdVGMet99hHlkphcQ
`protect END_PROTECTED
