`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THOtdeZ68bX6f6c1Ixf4nxBmDy+fwNfE0brCoynJ8Nt8zHY4ibiKk/rzO+YCGSg3
aZZ50yoFU/relzstFvXh5g/DdXqHKEmnY5TNsI7vtyXMoqxMV43/s8AugMTHuG0G
MOwZoWEBeCnatDi9QAW/3fKW4zyAW7ALYRT812qnBHeALC8VK0pc+mQGY8A2hLwX
YRSbmJ2T3GRl3fSdHNqQxyfiPmcuJGj8lImViU2mKoBMd64+yCt8BqCWjvtBn3OP
xpArQYh2LHXJSlpOVcEbwuvst9iKx1uDuA2a1PfmS4hABlNO29qF6/LDXzbiPv5z
1TIsf9++R2UoDRkxRxZRfwSbzdMIzeVMHYf5RBlhe7Zl+vw+LaGhLeLEsIrqq40X
n8KOiQlTsIwLDrxQ8oXWoK0wE/OfkIyoJtTDs5Uj2yjDO2T/aTYtVCt1fK3Dyeso
AHGU6BjeHmr8/NpyZBsmetLaOA2u9B/pQDfcgf8QiZ7UD94YlbIkZ5WQPOv5BjCY
GLo413NLpAlqro+mfSG6/I103iWYGyMUVfszTM9BidtOEqVs57omzU8UoNByPTm6
bx+1LNZ44fiDQDqdpD/sp9L2J9lXXlvQZSmLpayyHwzGriX3Q7TaCWuYSDgVFub2
+ke1zG3tthPfyID1HH/XZj/R7SASWjsKFFqaJ1m6jeRfVpXP9Oh1hJAcPukOZXRW
ZBcEyLQSqGdOoXGxcYrn9u9H5RggNqMS4oKWvqmu8rkvvi7jC9yKkWql50L4j+YT
V7Q81BNZ52kOnEuwF1L0JmxtkP0uz3V7R0LjJo1NS+UyTvQZsFNIRLr7qydMNLHg
S3P0++NHtvoIU57MSlewG9L9ALBebEzo1v+XPTq8QQwjuYE+UpYOxH0O3GVrV+YF
VOszuidhW1p4DlUxYDc4IFWVYlVxKHrF0qufq2IU7PKqMmnLGegzLoy0/2nM2rL/
28knqrEki+8b0PGtLlYkqhIPhl/+MmM/NRMpnKTBWe/336ib+P16x3uFOeUwQ/xB
A73yIJ76nvV3b0lS+wBe0GpbIRAAxY19n4xqS/DnzhB1w9JL9mJAZiQ/FPiyhlpf
5NtdxRZ2p/P7204MZmRSyJ2mqiHiFMUF4t3ESGiTqSU3nw5r/wmbl6uWfZ/9xqtR
KHYU4//18AMIdz8XDFzTr7Qm/CeRZOLcGpqaDN2Jotx1Ao92h5fcv7CZaOVWmv4/
z3SKSV+owFdHTx07SuiBCSCfiTWaNAnidSWCq5YEnpOUh/PkHLuwANBl3yT3zDeT
6Hwlg33JtU8XJEggalG7Yhe5XbL2yvWi+Wj+PdetYStuwb3jeR1NyWa3WvHEtGaD
qraUArsePBWLhSQiT+Gcvz4Nnme4eIjpiMWRTE6GAJz5Pt/cpqv4qDAGORltL3Fr
/5wXQPbiteJsa7lOA8xTu/s8E7Cuzv4Y32GL5hLuv8FR+vwfRbTDNjO4T7O5x/pn
P87b80OX5sRFMcBlesJ2Ui6KELWp+Bsofx9Sj1DVTgoKADCnsi9k+xeLYcZ714li
+/7AYd+D8yMRI5hdWEf30OHCnp1KvR3Acab46NJKE9bzpyTB/R+VyCCAkPlxCvGn
QV/7/3DtgnDK9ZkvcwsWhl4PTm5GDdIe7Q5Pp0x4xgKVLUYkhaXqf3aiPsnQgdF+
Fstw1ZsaLH6rmXqShKv+COLV8ub7vhhh+7B0vQoRbK2RBvczfGR9ewKYexVTeRhX
WPA3b459yQZEOswMCRu/HkvLiXnnCL4UDWDITV4bLMNBDfp8/4nze4XrFp14vDZg
QkU2qUCsWMVTlh1A2nppcycTdb8c4i1lKgLCR8oT6k0qdce+cAtZMjRqEeGuguLF
hIQyNYifRpLVcxekB1W7a2loUiwDRLnF7fnuu8Qpcc5zCRmMzubBNfj4N7OWHKST
afL/3TBTdo1TS1qEqb7tfyI/u8eLw8N1x2FCt+Xfflz+EZ/5OYd2FwFdhJXvEdSD
HiKxjmpJCIOHgauwoITfmCRnyHkX9HOBGQVlrR6MqnLKXHSZDY3yp6yl5Fh1JtIO
Inmvf7tae9fgbUa2QNE8CT+k/MAZPg2QOfstcnNL0cjqMmLdn8AHEgz8vKOzud55
ah9S0xxfe3fC+1Ip5TgXG+umajI7LKHdnMXreFzWBDrKE6R63N4w5TOJgQ0cQetM
5jTHxJ3RMZU2VmHsItzDwC1eUgAwag/xVwPkT8nuIAD/EU1yIE4xDAQrqZDKOHUl
h06hiVB6AK1zDtvE065q1Ij+K3D6KKizmkyy4WUVVFezBy+zW+BiowCWneihCOvJ
TX41IbcS8+CcS2/5/9chlbv7aAywBC7lrbcz6sGf0s4g1i0sQ76z/fTOq5AXsFD/
xk5eOae6Ief68GXeV9AtLxGwSLEFW3xIo/Svh0jOBpVbnZ4AAEuGRBphdKRU4sNa
3mIhszdrbBK1jpcNixstKWHnr9DyZBWlUjVylOJUppfskC+aZcXyB00em4TKLH2g
xtJtydv467JpVp/wQHV82w==
`protect END_PROTECTED
