`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bKO3xzheK9WI29WO1TB44FSGpMo723Tjo+3RqQfIwB4ksGbi5BThUehf31hM/VXF
h2wai4pb0ddjGN7yE+Fj7rAL9DtCJS/NC3Mu+icVp61PiqPTB9QUTksfNFRCr5hr
1YxN5l/bttNkDeOOQHBs9H7Texn26Xx75anskvKGprrv1QVp0hzHzD6VO49mWYVA
gvefeqtzwmMoWG14li/DQILN/jnSg+VOEUqqJB8LOtJTJpCgnN1pNIppD9LKCAw7
gxODG61NBeyS/jyyY3PsUQ==
`protect END_PROTECTED
