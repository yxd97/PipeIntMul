`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2H7K5VUkuH47kUafVh2sKBjxMAGIRTGK3mTUzcfvCzHnqpOohRFGkBxp4+YivvQ
TICyn3abuXs80e8Efz9kSdjcDZCu3HaZCcbGO0dbfz+IElaYyddzrIqCQ/wC1/6E
xLGs1FpTr9amvFpJ38jzS85HQmO3ksT6xHKkG1Zr5Im2jn0OnqKyFQwejG62tk7v
GnUcKPktOv1xr+TGZq6TXYWyjpbYYKmq7ArK4/VY63GMd/ENQTxg/GiC2Eq5s7Fr
dlDlmSRi8vMMm71o7T+mRCfE+etZOdCK/mA7GywBPnXVPUnSnNZRzsmtidkgBv6m
1rl25J6xUxi+3+n+SkEmVyapb/1VMpehC/iTiJcer8M8REUmZTkyVs5mpXMRmsIv
RMdl/DY+vJYroxVv+WmUnA==
`protect END_PROTECTED
