`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUwlb773W52o09yqYCbac9AweA+begpFtMQvXvUu8G/YMPCQhbXIaFhG1vBM57cG
T+OTL+HJqmBgQp9iCOI1g+hdx9XnSmu6AzQwirsXIS36yy3ddE6RvyCvT2+t/QPb
Joi5uAelWxKXKCmv31dk2uRD0MErXLcoLtsJzan+oNtzdmESlm3MefBGE+v0k3VB
KQnqZ+DaFI9q9sxoV9PRWBHKdhtmlCVBkKgIeqdk+Ocd3N0u720iSrQ+bQbWwM4b
`protect END_PROTECTED
