`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3miHrxtv+KASltY7AZJtR7RbK1XGBVy1NACoQ5skzTID3wdsfqOBTlTQJhn2SlR
aBtdp6fMUC4Zj2Boe3jyJAZSaBCcQ5JDWIl2CX9B2NFTxfS4BoQkeAkSxAq0UCMH
a9uMsamO7T/aHmAa8vzdKEnJo7t220bdR710LKQSzVHQhLSb760L8usLULRlFHKL
bcjE+Shu0d2kzdcnVfQdxC2yDV7NVY0WeLS4QZ2b8hxIJMqJ6whdeRb3XmY78qES
A7Cu2vDiVSqcqPDfsEWfeakq7zi5W4KXVOW6GP27MBRqbtkWM0M1FQy/Ua8Ba/pH
1nK8C9eMHdnrvYds+OzQ6v8YnjqM3INKqVDGI+swbVQ=
`protect END_PROTECTED
