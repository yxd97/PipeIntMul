`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5Qkw06gjjddeWtG+bnVDOTYCa5ctkz86x7tS5wCt91OVaITi8KJwON/NfN6wr+Z
8CK39z1UECtbezNmy9JZjpIeQ2OQqSPvfy/YkCah8ut9TNzGGQFE+h5K1UcGRw0r
ovTLlkGrZzBhNzYaXw/3x4EMPXGEL/cVESGeorGlh6ZZTS3BDXX2C/z6FtidjUer
3J7AD2vJ30TYEAUD2gmpqG46Yi1kgQvdcmIsv1jmKA5pXH0S+CSbYQzPrQWZOWsX
+fsi5qBHEynG6mG7IrUTG/JZN8iWlUZ3Occ0WexwBdHM+rYylOxcWxYJRMLyauoo
8K5qvFQCbMvTAQBY0p/f+YD2QV9I7N2NWLXr2w6ilUeh8dTcpY5smq3gF9TG1hSM
7HS1jWuqp584w4HAHTvxuchTHKJWKcG2+KEaGSIVHICJbUkIYdBa2FxPlAJSixda
cLfHc8MbDKPwkat9qp8VVPQqyLGGRm3/wNqI+6lXt2gSnjakN7ahYXJaMUgRAysL
tswqblmoS8BacYFhMKkh0aTUk6ymEIZalIb+yJ135+iKFqDBQ2l1za1lnaqnn+P1
Uvqd3InCXZxA/J4rArbUJBxR47eRVGIz9jGFI9dTOaw=
`protect END_PROTECTED
