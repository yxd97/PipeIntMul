`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24LevC1nT+Osm3pGzde7KJHQ0K1q2/M+J+4pYm/B15x3d3z+BLnzrz9tRNKM6x98
gnJfLI7m1DLEeIZnoeFjMlW58svo8HJYX32s2p9GksVqfu4ekF75iI2ZfwZtntOp
3Ag+GLfv/hK+qdG8ZDyRKmhR64Re7UHHCHKF1WeRbhgVh0pBWGgZVk9NRqK3qYJu
sN/U10Mfb90tfyk2ee0YDgJ2MZVU7advvdCmrF+VE9uIGaoLUD38Dq4r5uRkhbcR
11sLJSajVrs1DoFa5aoPWg+TLBhhlgYSdI8TVH2gaiYHL0GDqKy4/mG3Vq49VlzC
zv2/ShABTFBKCl0LUBKn/zisn+1ZjyCRJMBs1H7OKKcKSeFA0ffRu917BoQwB4CI
NpWi6Oy37bpz9PIvuiTKZ73gpjhbuvpTpwx8D+w1lUbMm3Ci5jiohvKLEk8pQThC
GOPBJB7OSlO1IhuVR7EZOfHaGdqJtIlQjU57wLNJ35d76tGllE/mDThcGrJ4/UQL
1jVpd+LCVmKyGB7KxZvxp0HP0WQf/egU1ufht8Zjm3TSPES3VuI8c43ZoMQTThIf
`protect END_PROTECTED
