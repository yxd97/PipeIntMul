`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YLsamAuXetNwXHcZmJqnKz/jhPJh5wZh6jEoKSAKQRstWpj75cIauOsmEJo83Khw
J5JsWc0MfKCs3JEHjgReVVMNtSLGfazMIZl9Uw7QOASQBRunVKP9lcDnMdxK0xdH
2x1VhOs+BDU0Qrqa07nKk8KS/+UUAN244wyk+cN4A/W193GP3tJNEfSMw9X2PeAZ
tbXM1ZuFGvSm8C+m7Vr/vYAh82kvmZdPRSWzeImnxXt6PPHJL7u84VR4LXWfBkik
OLumcqiTw6Fn0JwjqThTiw==
`protect END_PROTECTED
