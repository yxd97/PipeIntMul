`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Lwf0OzIuvrkdKUnmXBOOAjTrvksTJ+bLr7Rxx0z5n33JFeCEkPQXMEtg/UJzzf1
afhiGGy4WrUQS4zjCq3geRh+wXmOp4Qh5HPsBc32j0KToQJOO23pnZYsoGCTaTLs
SxiT0AbSwyr4RY0ImVjXP1EYtv7Kkb7NzDKo0jaQ+RSlOup2Lsig/06z1kYPmNPz
+RhjvyhQV/GKIHf681cmjkpWx97J3DAAzP6b/apKZFyM9j65e4F8OVrTu4pYFu3G
CJddE8JsAzLau1xcz4TSKH+ab/pXx8hZj2gx51BfJJxFkvk1+q+huinMG9W1pc5d
m75fQsprJgeTMgFifo8aBPaQe7KjEVVVG63bBEz3UXeagJNjZbUejTjkqKFRN8Wz
Vp1WbTJKu3wBZ+PnAKM2Xiw5noNhHOfnEHIVub0UHMsW0WiPQTU97lrxs0aK8DbH
qA2kMxMko4XJUBCuv4hCeBtepzh2plqcL+KnMIQWDGb7pQncJq5ilqtwpMikYkai
VsxiS31cVib2/rg1kHrzwY7R5dda+w3N8gqzZABTTGeihoL40Qsjqk3dhCTLbaag
RPEpQsPjKeVbNhPap5AdNgIb70dXpth/m8mFWe33/vyra/hkilpAK/+CXakcwuD/
X8SIlxr83Jme+11oHq9PVDFAM1J/sT0hgcTQfIty5cN0q3j+t4e3lUyuIxUOiaDI
D0+wY4PJnGeXRm+WHrV8qX2c+P30gQkJc45NEbPGB+pZ/QSS3eQOe/pLZJ3FPYJ2
`protect END_PROTECTED
