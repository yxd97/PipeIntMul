`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6f7K9VOmKoPv4J/p03xbiN8hXMw3146RNmzuc3XvEDHv6nm59dIt5uxCEs5L5w5Z
0AuhhILGsw4dy2PSO5ypT5B1erZj5MfvTi3xqljKXzHbfVY4OBc0P12Y9TasbDNq
/2+bRDFcrkwvfUd2RiQPRcxOSm/kVbfue1r0ceuOuJTLSIsGh72M2yQ+1VVutqXe
qRrVYfgyXXgqaidYraVR70zkQXs6ybzMkZzUHRkN2BNVJC1KXoPlqvBtWvt6FpK4
Mb6hjCgIzJ6iiGJJtHw5ygvZABrgtDv5DMA9aqEuJhQbE0//aX7eY80omamcLlXy
TQV5zed0vMJLK42a4Y37oxA+EtN/2VzY+j0KfQX/rFbqGNdPnIUTUgbPE4dSCU5K
hFeAWeyFrqYB97QgSqjXIfhYnzVpp4T/KPwdSG9N9O0=
`protect END_PROTECTED
