`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUs2bJFp1naI+tyFlkvKdKktYNG06EFrtVpQNDFgK8fuKYlWTN99tOcvqyktq3pi
Rh5VAm9obIzo2xqIprB5KFZ0elLFiJp3VAlKmRYT25jOFZmQ2RvZcBNRgE+0pNQc
Az1gWLwM64i1MrKhQNZ68ZXivPaoC1UqBQTryNjxBzanJg5MOZQv57lfDTLAPQLe
MOHY1n8/whYG7/FhAAsSwq5MRgWZZlRRpirDf92Ij3tfFlZlPX9jyJpefgHPHVfk
ds+komMzWiblyBTQ35RmZgcYcG8aovR1m1+HfzAJLGDA8yvgVVkWkbMsaM6ku4n2
JIuqf5YQ3zAmpoCgTkCnqM/rtglzi294VPF2SLFv/9O4Adx+cQhH7FYva+orbZFW
jItf80XpICxGcMh/Lfo2sCz6+KeneNadcQ2HTrVAyow=
`protect END_PROTECTED
