`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYvIUz2SjsgfM5x+Fj6kHQBkBRWkpmLdEGz35XJH+CcnlimqIRDpqdcUt3D3bT7f
17ZicVi6BJ/JC/PJLqTc0aAtB1/gTyKB9/gUCJ1eegjr+t42dqjYptubpPLR/TJ4
d5LGlS6ya5VC7J8h3QZPQdVoWwyg4akz6sAOMR23ZwAuNc8RdmNRvh2ttkRzlP1N
jPpBQRQYVvs3LgdirtrEBjo0p7Od449JrjSOdO8Xh+kqJWhEvL5v/OTrveKYjoov
uQZNTs9zwGV+vEg8p48d4uwvQiO+8zetTtGKvBg9Sf+U4oeGIshLthptoBebd42J
iCEF6MxyXBX9w6LNpXxa4+gztCrd0qUBSzT9Ag54BUJ45NYMcroaFwR/aOtQf5eY
GA7gbxOaWMC48p1K9m4wKZyE/9SadSkQUs8eB+JLRYc=
`protect END_PROTECTED
