`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gq+zL6Xmr3ymfK88Ab2JY6mJk/gpR4/RDjM2vd5R67MdC3q+O5qkkjJ1kmK0ZAqT
UkltFI0NuRbfCCfHj+ihp+hTIXasABy5wmjPBt5c5QK27WkOlpPBNB8Oxncn+YlF
HiVVoVUuF3/i1sBz84DZaVhxZFSCDcnXFyMq+B60Z7eAWauWtS3muqgIq/w/vAP+
nNEJk7G/LY0h+XduFzXEjwdOH+1nDlH6+zkjjbTQ25yKSn8nH92IdEegQiIXNwsm
ckEveRyUGM1ti45L6ScXUbYxnYlZLnPiGWJq4G5hdaG7ux9n31mzIdpLP7dZRrU+
pkvSYeu4bdS/kMoQOS1I+pM6hZNbg2/blZz2/D/k6euWQzlMH6Aa4W/S5g4iuG8e
qjux0tMLX511McNjG5drg4kQbuncIJod9smOsiCtqzRv1okmDLwG+Od+cr8OPN7z
o9+33uoLPLZ386YIPcfYdbL6RyMr6PEELlMfvseTxlDfK8X4/6hfruH3uPVtc69n
22nMN8TwCD+yVqkIrBsjYQKX11QBpe2SHb4bqu4qh4zbxOFpdmLnT1ZZgfRa/l4j
oZ3jDSzdC4wiTTP+wtaKqrmOd+E2PZsb5CjwnOu2oOsqZjkPsDJaUKolWw6ceK5W
5mWYlX/r6HCVbiin549E8ttQHxUfQxn8oTmPlwk904Nv1kp9dhUGtENPDuqBHU3Y
hAqYNAPHJENl5RTP1UDx1VWuLEGEp6Qm5ker744a8FWYRlI4PStGQFcX/JnNfO62
8mgSIjfcxLegagZnMiuJvbVmjSVo2bjn4M4qB1MwStYCAeP6vtp78OJgAKdsJ3Sh
E52mjd15X5W14q7xiOQJ7ckekR+FlmNeFBDDjewQpRdj2CO7ZC7BZuNSn9jHF5lx
ea4DtKAArR6JDxFeO+RLixkOFqq8ukzpIhJYbfG5uPgZ3Pt0YlJjRtVbUtXcRTU0
0xEPL5McyCskMugZRa0qUnN5IRZwzJ3c/m7A3K900N4haT2qZPWl15i6z4i9g75n
BSyblmZKuwgWsSqfn9vBVvr1DLvhZa+eDhajQuaAYUSj1xxn6+YA5C+IIDORvgX3
VRjWkxioiHFeQJhMA8dSvjF0sOiFZHZ8f5JrYIbGQoqfgIAKvjhUae3PfLfaATTa
qpLTAVJ890RdJtlQYCbcIA6K9AuXRnuS6KM4JNb0FT0nbV3zhqfdhDGFNaFMUI8W
8DjyjByyYIDL1mHp+Lk8ogcsOWh2sVAGZyRzHfdSiLt60agO1jTU163OQA6rkHyQ
9wkGAex5cm6epNbqnSlHz6VzuwzZrZiRdRP8BqIRvIxgo9U0YJycS8EHRRDrl5Po
uwwnqjpLe/1gQh7NXSf/NxWAICAO81q93CoFn6y2yUmMdidq/LtdXDE+LJyIiGGA
oxLx71KFIzqk/som/G1JclP/YEAGSzPqt4JkTQF9IqHdriERJANUUWDv5gImGAxy
AEwXPeFxiw/j0lF1UEjwOa6VjvrvS4ZN5gT51LfkOewlGawUH3nPp2qoo3Y805E5
iDGMpYS5AV540NCi0W6roDqzcF4W8mk2vKuhw9MYVZxbpUgOFEdPrjRzLqPwIlWb
9hK9kiNuBClalm/afFX6kJycIr+2Eb+HN/FdBt/mte9cXxSeTQsMEzP/Dk7gvVGP
d09i0UcQe5dFzAymvL/aO9D1oQhAB4SBkrmKoGI8hKHj8HSuI9UzLNz/6pAUSqtu
/auG+bxtYqFX6KxV29CK2HzS/N+uaQvu+13kiX3geco2aqASNPV2LDfmzf3Dm9Wk
rBvWoUcuWO4ea6lgdl2IJ31AMdmSUquF2NW5zewtTZT8jCc2G6dB2UQNEktaqymS
mXZ+BtWi7m1lQm5YL91KTzZnRm96e21tXZT8rIJHHZS4hSmCo+hwWvTZyJnjSOHp
RwOFSeFSQy1BHLFNILlPPgX3IdRQEDl+KU45jD0pMj7dRInXl7rqkNlM/NEHMO1C
d1G/Gx3CUFcldHCHtfgiybp0cLMS6CtchowETSte4WMUBBNjZXsw+TmcBynux3xP
guiLwjESRTn7AauQBBI4A6UmQ3AafhpMOEas80J6rwCC11QMMfbHT0lsfL9uj8Jl
8MJFGFIYGewv7Pw4HlVm1gJXM6/KNzo0CeSxHyWXxs+/Qj+yC6X5nO4ULRdUjY0U
EMVVZ+/BoYur4jFnIjzIWP+pVTrscv4lRaRhdj2WCShWXlIYiaWqfin6U5uhttue
tUPorccn60Jwecj0/4To9pmYuAD6hONyM7yXrIVPOqVON/HM5SF7TjvJtxPkKBTx
gqI31iGLpSJ+IDH53Qnrt8RxXWb/4jYl824LsG016JYsvAaqwBJJnyHhdtRbMxv7
Ctk4GMWB8IZAsGOs3IYbAMi60gFpAMcdF7dp/ff4s2SKNyiGHYwzpU75cJLw/M/M
RKDHe3WzTUtCh2ZnSbD55jHoPbAtIK8cecW1sdgi9GUMUFPVKAxz/K2y7o0w2dXB
VWpZuh9lxhPIZYT71gtVLQKcIQCxlqxi0wYEFvm3AxX0HFusFwlCuQ7z7z1qKzLx
i/oXJGjuqVtj61gH1bcmI8V9kRhyxcfSyy9REG1TxzU6+tsiOJfEpnXwrDNGyGA8
xazo0GSWPZpQ8qrNPlTSE3EXzyupxCpEnVIslvu4tSkiUro4qiL73c91kcz7xTsF
kQ7uLithoFpn8md8bN9yYgylQnT3uwz1+exJ8u12bTkkn655KiDhL0gQQFcV4Oq7
6IxOzKli76klONzONXZiUuDcot+maOTE/mFHpv6Tww6Gs/w688VivT6VO6MjON2w
fwh1oqcnq2r55Lv/KaHDAW4Exy+YllKy9VOcI/ZwX2Ee+ENH7cx7bhaYBHw5X6VM
VqlzfhQ40B+ecC3yTc+GxO4xjR8CyUj3wLJKXWVytn7fKdwVtRTe7rUj3rRnzM44
6uXXRYxaptT7hGyQsLnfpmp3h6jd1mTFfNlSmfH0OaDz7PY4xoHE2zx7kWsOCwgO
68KsVNZQa7WH5PjumpMFZSjOy8OubzrW38crd2juLVSqJdAV81hjGOIzpj9QCL4n
gg/G4sjUXy8E7HNFO8n9FWrqHe+7FPKwPSdmC1f5Md6BDi+Zd7DtO5i6QRsUE0uT
ZnhMe8Nayj7LlqA1OcEEoKatz18W9W9vqi1269bNuzCYyBz6+UfhG8hzA2DEws8E
XYX+JwIVte7sd8rXysu5W21p8e6v8usB1gEuNoKUr1cqbUIpRX9T6rMQfZqTZxrK
eQakns3Tl96dbBJJ8spxZnkPmWFBYxoTlBFQjgX1Y8lcvfwnp+KDxxGQ0XabWtsT
tjIrdDwDVwMELllhLfrRSld03Fy31/QSssiDj6JPYePrVBC5P9ULBOPVbRPQ1H1F
Nphx0lm2EjUKum3wAOYGm4LnbTg/EktAOXHzIpkAQZwyO9nzm0PYpNa4oWAaSlrO
6SWicWIRgoKcuXaPt4GgRuld+cY56w7eVOFgVAys6C1xyd7zdl1GPSki9KGnY2Gv
+r34vTohFM/vOeuNZkameVIoPefVwwdDLCPN6xAshNGcqaySjFMWVacqjCQRVzSK
OhK2bDQBAGAL1rOY/VrXUDkDERfwdq307EdBZCV4oM03tfdv/wKU/XPBqZ55ua+q
i2twVSyCyXqNT2UjOdNIPkakWWE5bBbEE2+EP5RWtG0YfeIkstrJujCE4o/2gth7
3ZU7nSprIyBml5H+K7i8eH1pxROebPeyLdVX0YLFJtGko4WTGTIihAPlQOQksPcs
tVvKecZ2phhv2MK4ocgloePFQstGLIl1J09pdT0hBPBxjBCmyhDAIrg/mN1nHhI9
4f4yOMb1TGDjjphbQU/+8eMlSh1JcS/RoubYa7zyifKtn+x7xiVrU3qTlqaP71q0
+JCIGQIvgdZJlzN69UyAtg2T/NTyJAEDjvWLwHhViAw93JhyGqCmcIa0vHObJ3oM
`protect END_PROTECTED
