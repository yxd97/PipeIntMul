`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/El6i/0vj1qg52T5j7Kc6wS33QdcmZwSTy5AsQlXPv1y766O3+bHb9tuelqMrf8
mTgrQddvt7Hz+Pvd8ZU+DDpOb8ab9BienJD/56RCVj1IgKCWxZzuag4pDw2Vh7bO
QVxdynvtcRTVmpbe/YVFm7CJjHA1awW8jm5AdOwNthdw/PRLne6lbYIn6DT/f5sY
W3OCrJ8LN3VVArGFOiJ1tYtaMVr7wQ5s8cupUjvMYCuhotyFI47nKnvvte3A2Ii5
bK75tkefpjU6u/uR5sq6NyjYOFvt4JqFMpZkQISU3aKJkSmRYreHwu1RoJqgPSep
7snFY1w624oFfwTiiBYDMRf6NcSVZpbzBIRUz70mice7ONS1b9V7tRr7YR+L0EOb
lvAO5Uu87vjnNlI1MMiPoHphyBNtJkjwB5s+3S9fyPhiz+bLwryTlbKbvFilw1qI
`protect END_PROTECTED
