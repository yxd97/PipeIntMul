`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StI0bRzd+S8n5qhtbod8tO0MVpM8eXMtU/umZ48f9Neh2dzSig53uDmQ0Nw0rHY/
4TcJe90jEYxkxP2rCYyvee+7w4Kwqnair+LZWoV5t2L1T9+99jLcrf3LdKo/Fmcl
oID0D5BmKnpCJypgyhcxz8IuQw7vEbflJ63dvbWFVj0Gqhz+QWSbdWbXSBavzfDv
PM69kf5INc8OrlI6o/LhqZfITuzvM3RnXK6L213/oD7dnPHeaBEnjPMFpybGOGJ1
tzTCChb3kdnQZjeNb1lFk0X+O5EDd8Ou6baUYL3C5yz3pivHy1Xl6WMB5PF1YTL8
IMFXj4z2/BenRFe+O+45mTPagDswO201LgNd65/aSzqqE/oTLEiZEhPnUImazunU
YedhW0zxgfxN4XKG9gSIhxxhxcR4eDFZ1Ioye2nOr6yYm+Lh9GbK8FGiQzr5PYjs
L31ybxkKuMgiS7NI14ZK0SfTJx2xVwWzzvagaZD0l/LRiOu1I/lZPEo1fAHE5r9v
emZFlS5SqSFgTLhUYTWwUApEYBfGdEzHCEZwuy/IMkxpgXuIrOiH4dKZAo4Ptxun
S78T9/l6IacOlsp80YEZBcw6MnX5ifrujeDB/Ix9e2ke0Dp9aOgmWWxM0RNz3u3p
Ae1Rnw3FUWhIdw7wYm3MEL/aVl16QRweg7pbp4BtVvVPjiyEeHlg63loNmx7bqED
e2liDvL2ouZO+nxxmSp696lsngsr799fRvutfhxdYhRRfVagH7jXdYQJYpWnWme/
Qw+prSZpYrQ5XrHVNEZ5+JrRt3lIsze03uRVxCdOcFCgSg28/HSIsC4AHa6Ju5Hs
hkBNzAPjQskMwU2fmxRG/YivzQS5MSrIvWImt9/L4u+0jXpPIS0Udyb5WG8jRdFc
aq2UPEIpwKGISnYUh+Fd/xAeZm1qghwIvpBGuYoQ/fg=
`protect END_PROTECTED
