`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5HalbDTZeTEG+/Olht+K0KZJd9brOEShwdNlovGXPEviFZ6nK/JNQyF5XPpQF3mb
KQirsaInSB89wSCakB59qm2o1Zg5Z725AJW8KwmiwEH5HPbZ6qlqMXvh+rkMUu7g
yDDM22Ea0wXFJAW94C7jiOGQTjGV2+oFDcCeNv43R35OFdpTWL5Kui24Xx53YCnR
suchtTnfuBtcRnUJbzgvHOwaVZGaoK8SD4vC3+gXLiRG93W2+G5sjawQlr7X2azD
DUh2SFi+hq/hFZHGEW2/YaX6PxZeWhYmDqgtgi3BaS4IfJ5tQUMdZgugipapW2jC
0Zjtu/nj56FitQe3fA3/G2sEjWvHqmArrymfH2qV6QcQR/hurtIo2Zn3Vno+gasO
/k3u6bfmnA4eqXL14WKdW3IpK2ShAXuGbQDnfFUtgdMfJ+bv9IC+xbacEDWiM9z7
zSrppHabngOjz3uDD4xrlvPxhs758wjSRd7BU1+Qv/1cQVwOCYvdEZA8Yg/xLGSD
Bcf2dnRVMK9OGa28B2qEW0ZQ+Z6rqBFQtn/oJIJBp38R7NGtkIo/mwJdMjoAUnYR
7QKdpDhBBa3ttd7pcBhIFkENa5tuzGld9bF1evSlxhyaa4rzdmHzR3aPRM5ojYOW
wZWZivZLIHzeJKEtCmSjaw==
`protect END_PROTECTED
