`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSm7mXZVwYrvHC51/2SXF2hWo6/Egw+5GhT4s4GF2pTh2B+jiK2aPEgNt0ls7q7x
QmbgHFmCfp3b4OJzUU6RcFH0GQOuz0cLXDdrO473JizmC7ShPNQ7cgOL6jOOvQs9
g+SmS6D77RTsmHorjkwXT6RfznkIkAZSnjX3gh0rtkCe0SRmegbC4strWcKsOzTb
xWrukg9MNWWmaDP/XE1ikIJPoc8jwOltA+3yW2RUNqx6P1Oh7J09g8qPg3FS0Ycf
sroCkI34z3tmBu7LQLFwoM3HDmjYvqhHowVxxrbctqFA2B5javZPVOKZLa3uM50R
D/EaTvqNVaIienkegQXKPQ==
`protect END_PROTECTED
