`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5kbXhfgnX+oizK/njV6L0rfdB0uxkFk/z5BjiIvOrMkkVpXG9Waoc55e1a6i4qn
JUr7Ljiag0odrcLIq7H2gmz9i3djWRwJuFFCitsokOLmpJa466HWG35JvWUJOJCf
qSgG1FutldjDa3DeLVulxGAoV6/vdYqCoL8uyyymUNmRl8sBcMmzQFMSfSxkIe7z
mxQfnTZ7ZurU5qEKh16jNlTN88fynB/msVRojbnnBVQWQMVcJT9kp5NBI3CMWHS1
E5yW+A6PojtSUiQXasS7nJrc6p2ivOe+SdsSbSzGdnRVz9ComnJYSFd30ZwSCJdF
JF5nBiwHDIWLA0uTOrwCIbYknYrZtPoQgNmnI+EhpgLdrBhwlEOEZqryXyydv2z7
zu+AGCy9Bfmd0c3N+eZyIcmDatLV47wwzj+z2v7O4r2CirvgZabia96gExf3Tf5/
vgznHg5igFW2cOlLWn/TM1qNTshvB49V6QZyiPlsuqvyD0ICNEwEVQVLOjvfczXd
KSSyWkudof+JFzrAyLSCE/YXI2zHLR7HVYxWzP17PoUBDCytob7A/rdhvGV3Y/t/
Kg7A9zy1oB/ll3ym7bUTUtyLou1tm1pO2QRIPfHOMaH1w7KaRkJD3yR8e396AJTh
X9/wFydm0H56+xkpVSx0Kg==
`protect END_PROTECTED
