`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V78tqv4KpU2mkiJ8ktjAYhOmcI3YBkkZ385RUXe3CMeohDUE/u4fRQaXq9WSlRQn
Eh5QBfW9S5JeumF0fWMz0xyIYr+ZbRpFTYY8wr77QkumMSijoRGAsdccsDi33L0b
xH5puiy8N6ax3wdTStvFYOfGov3azuHzE25gi9lvVJZwxhsSpmEwh3eqMUQkJfqj
I8QYFD2fLsShHwKddxnwVczMUPzeIlQsHOSEIvozAdjXx8xbCOBVqnXfPL5leA2g
riRBwlTvihxsUw4BjZKoNkQ8y5xE89zT8SGXiog0dUVywAU5QbWtIpVaZ7WgUnyC
3zNCR0cVG0uXSEZdqzePk1ZEGYmRUy+UeeTUpnHth/mpt9/1gC7mqccNtmJ1uwZU
QGouTYBrsK2J/6QSPIRQHnCOAiR49BfJMYA0ZJ+FSnMfYj8hs2GZbGJMcfUdg+nw
y1MpRfo61WOtKLvhKuCLl9AN4CqE0z91focZluEY5jymw3p+sQiwXxBv2155+IEe
ZnzEt06i6KCqo+yVWgoICUSTyq6CysXgvVhssy7mk8+Q2v9b5tX/uJ+JDblfApIG
v3FUdVh9Mr9G6g51ZTbHKI8E5A5aFrq50iU20ErvoZk2dlK5mVsm2Z1bMcTDd2bq
mxaPuLWao/8fiyoWhfVu/2cF241lui1i029gN4xSNI0NcbG7asDdYt3IfbXCZ7u4
yUhoE/Of3gRL1rq3resXUhZy/ODDg+wocawmvCOHeOwkuhW4bJZeovdW+ivbZDcs
EClpT/Cv0oapOrPLpoziE0LRLIMFLV44VR71yiobl+5eGVhYLzMJHJ//dpZQ9gTC
9ldkVTA6ldICanJv50jdWoZfgAdzTetvz8hPQuR45wHFI6ITgpmakeEl+901qKpQ
6RpjVVSD4PxYNRbJApwQOCzot8ZeRxvS8LhgmghGNeVzLeUOzb3pSotKu9IB+j42
UTHII6uz1lZZVhg7/XBOlAb9RUgIGjcjuFC4RYzzGH4aQ0wyNFHkcDftGqX2M9o1
Y7zindwjqNKDALFYzuXXUQ==
`protect END_PROTECTED
