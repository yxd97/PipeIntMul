`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKR6l6g5SvKFCEwHPUeTgq2ygavL7Ykv/nNBI4m3P+iJjO8IcdAr7uelxXr///E2
4ukKgxpeWNNzXw1SmrCLAcb+Wi/2lt1hFSPnUFvDSLB60y1YS8PCuAUQMuy74oAT
YGKjxXAwdv165JuE/kIWiu8K1bnd4WjXABU9WwElCm+Pqb2ku9tbuqDLuHMBb+8G
dDsShaFw+76bKcml0S3B5puxGuNfpTeOHKghfqjMV4MNw7mpLLTMv0Df1gyjQFC7
o5oYP9Vjpcs0Hs4/kQIzcBvPuAp4/8bqNgeGcNawLKlZ/GG76yOyVi8qGAH3e163
Lp8iXBmFta80DL6mYQVO4KS1oWCam7bH+EVfk5eKdDflMos+LbaKtitSqcTXICVf
HLyBhTa7Kw4ThkHzLz/XiN8HspWxZxo+Iwu99hpM6UqeHAcPrVq4c9+8utDvEtXx
TGSP323TzhzBtjaz6+HLNpWAATUMmOe1dmh/NVumRdMDCQDQkc38zayGYqc4eZ9E
itgGuV/cpL7DMZuGI3UlGuAgR7kvpe1Zn9/qN6aozuombPzj3PB1S3+/MamRtNoR
jjcsvyn9R5iCt1CfNTVJG8Jek6jLFVga9mIo3w1IBDyC50+WUCnFNmxmtsWThVF4
DnlPnjpZzpT4P1Ve76yokP9allhwR01/L6m4B4O3P5cO1by1MBvNDsWl9WKZ+KU+
fQcLu6ugCSNg33D7KB5M4XdpTotosbFncGe19GsxqhKIMbJLUmAtyMhJOhRfDGC0
jHtv2F1L3SwpVw0bhXzqdX2BRdOatGtHXVR90a3UDSPgns8rja6euc/AWdceFirB
vg69gUYnrUoT0n8sDeRllo3cgzo/vgavy8nQURZvz1JKyuoxiAKc0UFt/p3sEK6j
+eIciJI9iQWxWZNMDCVdWE2iauWuWPrjGMC7cqJBpfeIKphHNGTbh944kNN1T1nv
oHNPGb/Wp5ubgPwlEdVRKf9wQJIi6/h0LT1Z3+BK/Jdd+iCw14YyFJR5Y+DY3jqN
WwyKoevkGvMFvJhLtWfNRhbKjG0ML8AaVh9XP6aQ9mU5xyGFFQqgNuQvCFrvd+vm
m871OCu+up0y1C/VX7ohagvgsuetG1gT6OaeAOop3RFrM6M5SD+yDgoOfPtwHXPZ
m6zlg2YMMIfMOIgIIz7uj5MwFkgiBnCWMWZlANF7C4Uz1M8rWZ28S6qQjc2ng4zy
cwBy16MAEadwoD0wn/q0WF29aBIbqmNKgbWeu1tIIybqbM6znDIuOxer2gkrXhgy
ovs8zQQr7cxzAjMWz9UcLkNhszFayIV6hAaaCCdJgZ+7TFlXNwWMz5Y+YV+JeD6Q
QPYdmzkUU73Wqv9MViLq0UwqEZ/nHD8Q8xUQwde83WBmeElxsLoWJPoyuLh3pbv5
6WRHHV4SWjSfjcAgEDz3OvO+2RdIm4blh4Hw/x0JOvVpMsRbU1wZ87hcV86Oqae4
Ih1/ZZdIRJgdi1xTzdeR5M0OUPssvhtjSWHqkX4UYC1yWaAOgaX+Tb+QszWEAeiI
wjMl8WbXzt61n9Bs8eOLcHAwZVz0vaNZ8kAjFJ5dhOzsvB3Gys12/3Kdkdm7k0BK
T6WeGhTA/VnD/c3VnxVBu+ZuG3dWDNttH/a5q8wU8UCLK/c7k0xXyQnc3NAH6ILf
PUmD7QZUEqlDN6W0GSPSzVrX2iQzlYNG8viSDgYcJ34pB2925mHKzKBrWCfSGgFG
BtM4/AtFKwq9G0G+pzfbu1leKoTPyU6TfjIOPSUCKapQwwaKLA2neyCpF/bltI+I
ap/GoJiXhF8CcIwhy85QL3mccJXx1Whf8pqjoLppKZ6a8ZY7NBYDgdJ9cW95XVqT
v6/BOGk8mZtcL3zEGlB9K94jSytSAUk3AdcqZwdGmomYzgXy/ILuBjhMMSR3u19E
5eUb/uR/rVyFxJ98bNQDkS5FDRilRXyPNOfL6wzKDt5+FAmxu4oNhkfPN5jmL8vL
/cw4wc037B7kropGe8EwhSRu9lUybrQ3RYTSrPronLNU5EjYW01CZmTFf2Hy/xlE
qF/z5IHt/RVmL9EVsA5oQLJ/my7D+YoBW4iq18FDukClgzCNF91Z/01CyLcQXxgV
25hh/oHvE+vDRCrprDLIQMpq0iwGPQoFB26cigf4IlLvZVbjO4fR13RZ3UP1Cwly
K+f8uKc0L37ODelnJhYxbamtTg5wfNkhAVqEDwdkctDLGO2/fst044ULTSyAdNFI
9s5lhhDHVkxFr3iQb3gHhJlQmKx7cmbGacolRH1t1mFCS3I+pJZYl+NXnv7R4R5k
az7YtcYQn6nKpbgCg61TpIet0OBWjK3EMB0XtBgkhr+/VQiZpHgthZvc/Q5oSit8
0FtOfVIGMxfGioB5VE7EjBXPoRXpktEBi8UTOARJd02NuBZmW+d3dvo1uZVl0B1P
jhGp8z52qjugcemzxSyxnJx2/xSLuQEGiGDaG8q1J/8Iqpc+75UK/l03boE5vgs9
ZPPeZTViN/drtcS1SnYmoUxfK7BaXYCa963nKZT8Y69EYMCftGKNzswh1xni9cmD
fl8BXnUwtXmPG/WJ5qk4T43MfUsbMS9KI4GPZ+0HWestJA4mTaRT5olTfrN6UZFS
97LrPt/aes6Uvden4HuC1rtxQNroLL2eiUx5RS/eiYUE065QJkM7pZOB+4YozIZ8
RpIayCZJ95/5nS2yT4SCG4tpNVWfhZfmL1z43Ge6rcKO4hZ3295ghh4dkmeI9BUD
mmKdiEolnybgNz7UzFY8s3egtXQASVYjZ12gDp8ipQxemk89prXBiAC9ZL7xCsQO
qo6mYaCszDgkJ+/lq1SZ9Tq3phixJQ6oaUD74RwZlnDyocgChlnO/v5s24CXYhIV
dys+dY4ymDCg2atdElQrM1c/u2UPolafn6KMy7m5vMLfs2VccYUA/yZIQ4m8vzKz
mFjKnVFX9eDhRioZPFM+KC3THTxqBYUVQSRlaYljwdW/uyY5aoTnZk3FQDCxXVwe
gLtwCN6WUk/3lsYyytJvc7AJSYeXuQFHc3dadwvxK8ADQ+2HmD5TFdVT4ODUV7lI
uXQl86C6dw996VasJM17W7TauePOLKMrHDwnUvyZohsTuSaS6BHzMd0T0dvF2zep
yTh3rZGvcqAcGhmvq4/VTmZJUNIwBbr/pH3iCEzcy5cgFgKajx5+Nkmws6MO7jEX
kbDwkRDsmL2utAKyOIzU92IPsikfk2KRKxr5hfvOHSB0NsA4yiA7BF6Ef4/+zpY1
ct+vg2iG7fdJUTQQdzJBfaVkWU5uqk8hyXE418Fdk7TYW9dbb8M2nMpucKzwky+l
hSYngtDr5sngiJyoxJEBDue/6T6AEQzv9rMk1IWveeYXgbRnYvs29+yQiqexL9mh
ePj+P6QA0pLWsUHDcKNyK4kjS6SvK0q7h9zRGYJzZLCPgfBITxGsOSpCdGhlK+L7
Zj2Dox+1ZhpsVXxZAcqu8JohSORVcGFGuYGGzfPHFJgR6WpxKEO7NHIQrEKso1b7
hSVp/01pZGSfXPY917CqYQlVhRI3Z1W84OE+IvdBbFAOQiXU41rfEwdURCfEU3Wp
TXT2gISkrf73LIqVMzJBH1BSSu/IP5EuAbRgJe72D/Ik45M7bcZ7AYZpO/r4wKIi
G/c2pfBoN/N4DGmFusAWamTj5HC6w5t3/5yXbUmYa6oc/eTLnjGFn0riC7Dv16pD
QScOSAerymI3+sK4jTZtayLru30bOlexTA53jdkL1fuIkQrB9zU0NP9NI83n2HPE
jozFe2e/4SfzgLna0/8AUlTGk50Lvm2BsllKqCorp6YpTG6xNsBp1nvVn2wwt6/m
LJ55n5XUcqF7xSEOaG9DZtzCsYIxJH/4mxbTSK8mBlhkJuob8tiGBU1reCM5P+VP
Z+SmSG/zcuTGSg0JvzSF60p4c4hLB5tQAcY/iZFNXIqidwzwLNom5N0EcD7Fm69U
z7cJX1NyjTSwJstN6EJXyBHULc/HbyOTE0GF2IWFKp8lUuhp/QZSTVhNkn4O1yqK
GAecfj9C2GKxM1muGJwyYXembZog9bUwDY5Ee4V0l79NSvWcxaiGt4oMEJ1/wdFm
oC5lRHfPuo6ioOK5MyDd/ZwmPpy1NTKkaKCrI9TpksRj2dq+2+4syNUxw66ju0jC
2+8gx+GJZ0bGnHDMKOwC/VAaN8EriVgqKQAc5AsOKWaBD6NJwA2m8VggQYG7ljVV
G4PoLIISUyUXTcogI9FKR+NHgedVihbk4yAnvWRcq1Key9cqFYMTWk/tI2VwhMbb
zP15u2FPKMfeiZyYeKAhiaxZF9792mEP3eeIpZFKsQcvNf8FX4+19EUe/DyQ/q9p
PjrN6uVZMClKx+vQpsOAFrjN/Hdd6lY6Dkkykf98CygdM9z4W0sEECquPQI/H2zZ
rXLuN/tNBmmnAwyyCrfsRXKcBwqolbumzOmRMAh/jxH5uT62PV1AvmYCLrcGXbSw
WMjKLEt0X66h5golHwPkTa00P9ZapfAeKaFhLsmVHNDTYpPB6tB7qqsv3rKwSH2+
S0DjN0zqzhdXc1wjnRzRBzRuRpDAsa3HXyPF4NJrgeqt9/aRyNGlD098jvZwbjgv
izpojRC1TZxzAB4oRURGpA2OuHgM9MrAqYP+AH1F82P322z2gbL4OPCmT0tH/IGG
pSkIz6QKNfE0NCawGtWEloVTO4f8CLKcjCac5MzvPLk0xzJD33jmZAyvAewXYPiB
ty9oNe3tlB0G+mVPrVDbXeeFDZYtG17tve8e2QN6AmQ2xjEvQXy+dckCUMB5CO+/
DfeS4Hz5JUQAvsTK6Ybzpj2N03nvPobxxJFGkrgmiUo=
`protect END_PROTECTED
