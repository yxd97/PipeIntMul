`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNsWkEAEkfJMf64HA8OFXsv4FJnHmU72HsGNB7KsJeFQwrMR59FJDq/z0/VMchs7
+ya8XAwOoE6UA0yp4ZaHiESZynEkquRojJtSsTtS7+WH7wD9/FCJfdVPkQ81YGB3
q57rEW1dfijUY0Zc0stlQnj3QBJ0PSZvkFyDT+QAnwQWkeYSL31G4JF8SzRCRqWc
DT2ALvycyZmGq7WV8ZyFNc9rPUvIYzf+hUWkVqa50zAxmBeX0QymsKFZRbgsdvdG
24GaNV/tVhLVxtBt2K3eSeXs98aRXHk02ONehoxUUhs2Z68EvXANoUT2TTxAI/Fk
HDYsNgbY4a49/a16F6N/wIotTPcE4n39Hh12Kn8XEd2SOTMYz18dNVheV1mXNE1w
W15qjTitY8sKeBArymSkU5nvJmyXjWz7aA2LrSummRBXEDTMS70F5VyhlbyxNYR6
wN1wd4rF8cXqes08LiKPBcEnsOl5oTFCz6iXsj/PLob4SQ6tfGfPhDgk6uXwEGkh
`protect END_PROTECTED
