`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
57Ucv03clpQxoqvvRTMCf8ztSDC2/9pQDdcsNJiqJMB6ZTpCV7sSGVZq71lNW/+S
yGTzARqEl+BmTw7cDYCBTREWXqgLsjo7t0OYXv2QThF6y8VVQ4KN3k+Ye3Uibx/Y
R44mHIsr1d8jDmh2+Jva9zen+hsVmkkT0f16qoyHiZL59DeYVdv/3U0kjWPJHZsJ
QrWy3B53najXJBEBWlcPkrGyu8KYPhI9JTyfk/Pvp0jmvwUjthEkW6LhJCXqdSAs
epEeUOcmiYulFCNN5CqwRx9Jd2P3e56TTEC6kNPvCgwfKTBIJaoPcVheE4vK5ukr
2NyuC+8OkQvTRVW0gXDwmDpromAwUBxmo2blwCx7QYF6SvoZcl3oqqCuADgD+Ws6
InI9tgFWqUpH8cs+2nPWuInknbFmbrZ14oBUzAQGSKFvv8fvasCt0DayOeAyIDH6
TKIpNn/PSEE9tAZ+QwAqWPbld4fnaRLyjXukx/QivzMFwKy4txaX/P52uA2xefUe
tcRdy6MMWkmhg5u15wzx28tfc7VRJY/e0lKi7nQqFRO1CQ6rmX6OQyQAQqiyDwaN
GvydUwCLlG0edHIs4U+g5CDj82+Fo/6zClucSCH/qdXZlaJumG0oqoUSalZpGnUz
WCLttcbj2vvOalh6doD46IRnSq4ZKdES5JCqB5ShHj6ZyCNqXUfAztBP/G9i9Wdg
1CPiM1GQioxKrSWR2Ju624m0jolY0HUN7XFCJqTQMzBHxi5BjutZ13x5dPjmeBin
z2fhBaU3G87z9WiW8llpAAUakc/M7yCJsPRaC5QSb5CwhFvG7dvmQI3+BuH+4QJ1
P4uN5AzVxOIT09kzvDF1plOykoSYcoRWP9zA3FChZoHzhSIY4muVTQJWJL2YuMpo
Q/iK8FsnMzhm3k7mI1TLNy7b3hvCRTfNACtEpFJQbDX+BhPpkR8h6z5Gv2QNVV9u
Cec3hJ7tQ0rBxkol1a2LSJTrQLnRRoxwdulWDvZdNKp1JYlLIcWKdjIwcvJIZkdZ
`protect END_PROTECTED
