`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bhvv0Lxa9lR0eVGPbjlJk0+8BdMuOzeFXeU1s2t6bEk/yQMlOLYIuQf3lbN3kS4L
DiADgwIGEofwMJTbuz37+CSB55PEeoPOGYYlHVlLAd3rY4Owq1E5yJOOEGpSmE8F
f3w5yyu+I/lVwYMR5MRKVbXiZ0qVbbVoIWqAmiFaGMP6v5Zgek04oxRYGMD2Tf8a
WEFnS02ABcUZpH6cE2RliCFyhLS9uzcofHrrhLE9gFvU5cg+vbQzhh7cXr8sjHbW
eVTWkNcLXHNrP37Q0GtBzsYmyF9NfwE6KriXHQGGC8g02/38fWhsTI757H5qLDTk
vpokKcdOUTSlnl3ltF1h2bC1mN8nln31pJMSIuVfMDZH3GTVNS0iSIbmL7JtpY+P
2F2zmW86KfvJmEF6QHUHyv1MnYzpdV01bPaw73gynOaiuwRM0fyek2W6IY2eGnZ9
`protect END_PROTECTED
