`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
554pRt+V12Way7quExBDUunPrUiiNa7zdIyazUXUNfNhQ9Z57AS0TTaByVMF9QUL
kH+4MSsYcG9OiLL2mS0pObH71gMDaoYj0ch0k8pJyTHiRnAmlYfnXxv++q1xIbGs
3h018UWAEanDJj+QqxKsbYuVxlW0s0Uc7/FGlpXVAwnmuNd95lyIQpZpr+NVJOyh
ut0jJFKNvSRuuSda6pMEJiZIoUgIbjd/+SjnaTVVSP11B+fRzpHp3a52hjoGWf+q
aO4blKi13cUoqG3Sh5Wrlw==
`protect END_PROTECTED
