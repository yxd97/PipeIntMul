`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z5/YP6Ryo+M3xH8TZTI3w5FZVv9diRZjdwo7J4tOKAjMaM7DUZJqRFRZnH++b261
opVu8CznpL3Y6DbUFtnkyXlpdSA0Lz+X7JTBwDiIO51RaodEHrr1DA8Io73latHS
gVQolvspiT6v7Lebblt9l8LXhc6S2BxKY6RluJp3RLPvLJCiUhPK/dp8xZkP6VzU
fnnCALIquFlOGDivI9ddIQzxvuDV9WZPnWqTBxSLrjNCGTjtaTVg/4j7S9eJjUNL
EMpDoSYvSLlLGfRt6gS9y+Md3ix4U6rlywYLaNKPiUzbc1HRG+GU/7E45YOlSrko
sOlUSVI34y48q1bUyqe2gbWL8xJA14isIDljtbwU9aLAjcqrVMuGl2KekSqgibEI
GOzu66t/cHNt7tF4yQu1Un7fboGs8PjjpL3JHX2tIo+rcsfVs4a0tAHG1LEuTtZj
+n0BcEwz8ZCj0qzWc497gPBmiBHCpqzSqZiwz7H8EgFfxxqZ8L7ar7TcclW8JmYB
SyxDDDKmxy9mRXRaL1Z08Ej6f4qSELR5uTWRd6VpSUlSdknYikC1hj4lUxWUJGcF
+5c80UsoAGNnFP/KvGB6V9OTXK2YnI+pQ36xjTxemS3RxOKDfdvs1WLWmGK1psan
ZtfECab9jbeXye4Uh8vWaqVC1Ts7NyoueFqKH+vj49WP9tV68EZcXWJoXj6Px2ZG
2TuY7wkiSDBtBY01OZzinDbh7Lf+u8ubUzgLKMemgz3EmS8Wp+lk+NEzQl9iDnLI
z4PBWn+t1gn1hOA2QtBo1QdnM8ui8eAowDyOnMJZzJ+P/YLObYDGVklr1PxF7rdg
pnjGH5IBKoFNNvK7u14IASij3MStBaHw3iLfTXYdSSgLnFhqf9DnL8RLfnV2LKkc
zuLRnQmtsyRbf5QTZp03Rh9IQDrFgdOcwhImPjFzz8ioiU+lkCwWjJ/S5//ox6Hz
pxH54hxo3eloyL+7BJ7XwpURB2vqrEQvV5AnwS7yYR6VoKa0A4fjxiMam25o2Hna
cwq5e1FCYbR7cNy2i/v6j1+WgVxxb8MAtKCJpnRvRe312QmoQ114tceFPmvsrJDr
SaBWTqyUlDh7CNfTnWE3zQ==
`protect END_PROTECTED
