`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x3VJKo2cc6k12EO2RCcxFDUifWvUMcXGwZid7SuO2JLwhMUEHpfortjw0CcOgQei
cw5YAU7Vdd210D57KCQqx5Qy/3yJCpp0rTiFkmR8vUOTp+GJCEV/hhvsBTMr1xit
eNjBvSsXvrdlgLNepel2Se49/QQToDp0tGqjmdAZ2RudYWqobT+r87PYpu46uPr9
HRO8JGf5SrL6J5BI41o6Dg8JpbftQmAe4+HWGbHu7KHP3VhNCs3Y8JaEB5g1PpbU
D8qYKuit+S03vOv2txYhLe0aJTRFzqZS1kVxj+KliSiUx1HAJwtgTwJNZOAiMLxV
RL5krQ5Yroeb0tCl27E6E2yy4mfCeJCEdzPR5bPmkg7cENzsgZaTi83P8SMUASjE
57rgMwyFxz0lpZo8zhoCx843FOuQYsX6D0HFRRVWiql6ukDAzx8JZAPTvsGIE5mk
zM5BAZyGoVLd/lLbZULEZL21FPhLJc0c2lr4sorq+t4=
`protect END_PROTECTED
