`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qr/DuBzdHArkLQIKTRJaPLfBrWrhmUYj3c3r05xOLcDNeaLj3SdaYxlP4I3tZ3Yl
RFcXqzsfNqSMBEuvtO3ywYWcUimp7JwlFKWmm+RgVVKRmD0XjLeF4RXEeR3VU+GK
ZkcTVo2KGjXZkU1NVhz9Pl84BILYXbzMp43EaNb91LiLY0DYvCE376LeCJ7pJPIv
b3n3MVtwM0WYAiqVBi5bvb7pTCpduwY2EUT6JulaexGNGMIpaUbcGKf+oJkEl5S/
9chEmGElZ41N3VREikOJClz0Udh/8kxSrnV+Nv9VJ/dG9Xzzd0FNOCDbiCju0eed
+J4WqG8rMIpgpvyHtFkDm1/VCvT+qtCnpyWYpNlNNvKtf/b4pLp4Is8YnqNfhb0k
dlk3SUxv0H/DzeAlUQLxIEKxeNGlUQcZX4vLm0SVnBMU/Ulee1p6hwdHK+IIeR/D
mdNtmsosigE7h9yF/PED0lxZJ4uUYmDzVDM4lxL7M3gAfGGQk/3gwPcXZygS+apF
vYeYmlXrASGchfgPyXJEPC1nLjEAnWzSPb5kHxShVTs3O/vFResEvwezpqOHOE7/
8xWrxjr8ma2lN/JSkZ7pyw==
`protect END_PROTECTED
