`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LoaxzM95MvWSqmw7DqmskjvFwdBcZmjd+kAQ0NrPgeoYy7heWVcd2HlL4TdRlIdp
MRsgH/tnGqTxwSQ11xrP4yTNS7+kAS3THkcZG6u0TTaPbCkr6Ln8wa+fhjcDQCpG
symqGBnZvPypR3KZ7IcC1EwGYRJV837g/DVdHNLUO92xto1qt3HRhDiiBnMXuZ/c
VBQ3dhF7ZNZF9iyFbb3HkHNHvtqfzMpF5G++Y9f1FA5xagUq9o60co+P+UGZFTSQ
tWS/PXVF7PuuochhQ9WjSrO8uLHIOLh99kWxfqVQcxzkBs/EjyMTaA2bBcqgv2b1
0OYBsDNCvsheEa2xSm+ObPp6V3NEu2aC42Q0n/I0VIYeG/XyMjjdUODpUAzXjxLL
acMnSJWDe1BD34o/Ajo27g==
`protect END_PROTECTED
