`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n23kvTZCQw4ojRuonVKUX0dWLDa3ia2T1FRj++GG4BPjb9kPP/S6idvhMv79WH53
WUr6Oz8i476JGywiPyTwE/BJQRtwu46oDQ3tcqOodACDvvKy6SzYnwpDyU5QmWOW
jXgK7CPePqvhAGfO+t6HcPO0tXAQhYGR8Y4i6mgrQ7Ct5TM1Ppv+bSupLvWI6NnR
p7hQ0/yBGOSfNUJqIrL9QiELyO9RBD0P01+605FVfz8QaeTOMOOfPFJK6OHNokbq
8RFqLHMV3hubxaYft2Bgzt764f4Zs6C14g/JY5nhHLKV7BoaBmTyC1jfV7GzzH45
/ibXoGwcKZ40wz5wtjibPm6097k/7SZRswuR83kpzeXnjT0w+kSRQdh7PemV9qWr
SZcKA9ah36CL++ORqRMojxo7utAQxPgSsXgY4Xt7Vx58wueZj/2MNB2YYzza6ner
UO1U5OL7/CKMSw1eT55glQ==
`protect END_PROTECTED
