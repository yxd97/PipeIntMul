`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aur1q7Fj/MMp47x/A/EA7ukf9uRgDrx3QlPjffQ2jPnHCFtz+IWc/itF9jpcD1aY
82VHXQe/eeM1DiMasdxvYm2ZGwkJcRfv5HYdyzsJ/vETTiWKFpfhhSHNMgV5Bp98
jpzgbRq55O9lKNuKomu2BPsfuK0cNFJgyoPN6ZnNIc52zWI29vwua+Dx0FMBhewR
hbRO2hh04RCDhIWt/K+5ChzbQtTeROCu6GD9uiCDKb0NeYsKEK+hDuMz6W/0qskE
AaBbv4Jw3MDR23ubi+s6QON3JM7oBKg9dRGcdAH2dPBj0dqvKltfL13nCuk8sP/c
2M73RJktybVrmxrZ93jwAQ==
`protect END_PROTECTED
