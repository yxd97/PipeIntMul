`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGvRpmJQYeJ0uYz7B1GDoj1QbO+iqsGA365qZgbRmNYky9TtXyYU8fbkYEj3PDzd
s/dPbgkE8xaMwnxkGGqDxaMf8iEQcDflx7PN8yRaPEq6N+9I7fzSTM9BvwmqQWEv
bA5g2U38zXKYjRrEzihWOZjjF6LavySJNU+LIU60aE0vRzr/N918v3n2Md4ptPJ0
ZnUAYEEpaotWfltrYeBmIlQv0IzNGn5CR/KtsUAdkIxt1SD8AdaFo6SywBbhP3Kt
ijsh54tltpHYgzENfG2x2m/2w66/1uVwHxEmYWLgsf5+QkPQiQKLLlRn9CQ7do28
PScL3bxr5u00BJ3C46xOZg==
`protect END_PROTECTED
