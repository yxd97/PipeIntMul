`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iPs1lNlfUTuNM/bgUFYsR20TiuH2IoHhzylnT4sBkPiG9kPs9KOFWWjhT7O3lK8n
TshD0NJhp87LQXPfKytlQ0vk48q7GGJsKLr28dyXdrlpPAJ+PLMY0qj+x88br6a1
I6G+0SKZEqG+FRONTXb4pi30T/7KnJREPZ9NuxWeXemI+1tCqLX1krW4lLFLrU2R
lfNebJ2J37C4ZDJTizH7i1IeLjMKbpP/ViRuHw1bTlSzYutJtcpkIM1ncivkDyq9
SJyF0S3YBFCAkPBXVRy6rdelyC1SP2+CuMFWQAb55mlPx6sa5UlTZ8qb40gAZlFY
0C2Rivt+m5iAJ0K7luWptg6Q9t14bQUdST+Rm8CA2nyQ/jpl+bnZ4fU0WwNDkie1
4TJQfDqyuTNh+sZIw404AVkJoIqNdGnjU2xKHmMXj4IA8KC5heMYpBHEs/yyYA8F
YTuWPnM8inPSmNcy3MaHID+LCx/adbkVnYZnyohBqohGHp3ebbnsgNeuW1YiKa13
PZ11DZFS8Pdzwx/UjXUoMB5W3eSoKvMabQBMsUBft5legiXrDNGNQBWj91rgEFih
YOWD6wPeyqxtPY2OO7RhiLPtQWl5hmx51XjwqrQb5Jif3sqfbJhfpR2o4tPZi1F/
r0n/AUSgRb6LoyP3dSDT3tgzk/LQs6w7UGByCR0qOWYvZtsxZBwTsMZX5pkktE+U
yG2/lcCn+rY/VrTw5oQ50GZI3fRpexL7vFl7qfvUlX9mctvZq8pHIgGg3MpuIldb
z3D0OySyaGvoyVouY8hY2G9ypHD5s1rkN3s12qXGYEXsCcMjOXVnDKPL3vYKFimR
GtO5d+NRJ2d8u1nl50qkgVccsQPHP9qTbdLTCbsdCP8jEu4EjbUboYtfK9LsGJ+l
cKy4N9+WzGUW/wgsDdtiHTPYaSMxZDRiaNnwlxZQoLbNkLzVvRbEpuwFoD1isBPC
/os68rtLY2kwjlsjoZrJSyCSjATBQE+vmKIR5DWPME8wEMT3NXJCKUAeJDoCjWCH
qbJizPTg0Pj8fEwtUaf0BGn/o7OpcKdeZ4YPjitHW40ATHPP1+MmCTmZl8O48ds6
pF7OG5P60pal8CJkrEm76g20FgQQMWwLU1GLrWrscXuMRumBgd87yY6hzk6dlLNr
1GWjT3vgH1DSP3+J5X+dDA4yQ3OmQU/+/Bow9ZIIOCDAIXHjQgt1+F9Jwjl36kpd
j0CHmJtReyaXfWHvYYDdPHe/0or5v7X03VWYjBL0ztaWPwcSri2wYw8TLHUevfDW
7hv6BJcx14I7BcWuIBWHcMCS+yYMEr1AULo+EK40Qy17fhgdxseII3ZMuWRg+DHR
g1GvAg7O3GEriKNJ5alMzRGxsLGaUs+hsn9C6tJM5uIWkRrLCSZZoCqv/MUtoezb
lWtpBAqvA0QcCZC6woPDUNHpkjLEd0riG6jwUqZc41fGsgOEGYfTfBmQwh5ZGfdU
GJdSiTnBktXHHN90/8Hb5bJVOdFjcJlRLYwcoP86qVQ0I2buxvg9z50bIpQumH/o
hCUUq1869/aE1gDwNaeQ2jns8Pj4crPc3JiXS+g820i3SEbhKh+raHdnAqzQc4CR
RhijBqezJ0LGu5O67OJd/Y52Ex1SlxvDaNMBxRoYWasn5ea789ov/6TT0t5J+wiY
IA75t0iM94tBIiEFeT3Tw22ZhrGqMf2j4XDz9jhx1A8tOV4KpQv9+eSAB1qQ/BP1
BAtdziMspELWWJyiFXDYOguARYHLcdj4Kn1x+h+MI9xZmwwRMQ0DAO+E38NllPBR
nlt/rvru3fCtfN1ESb06DG1PEX3H7MEyVphvHf5tquMXynRrSQCtAuwbQgyMK+qp
0vFGDX9eqZB82humoCZ2F2Pkpy5c9GG4sxMGbvKNgxb1BpWAbhncyC+tGfVaS0UT
87GiRce5njnASRK5pOONOWvQ0r2dBKdLj+qNwkoCeSTQsetvbk162KeR25cxm53/
maM5mvYlYRMYIKO0kmA+kAOcwtqMWsslWlxu2L703ZPoif1yGEnf15i2oBmyEBzq
Fg3t133pN514c31TcIGkJAnYySXOCN9B+te/Z8fXJJ0RWi1TptikmCTMnWuZMALc
I6Uz6vUrXWmrN+xcFnWyjzS7MLp1JlDkgGIbNb6KCtoy7NIZxnoYB16l2xqPUvkw
ZNDtM5cxv9YbF6fo5vSEIrLuGHPkURiifHyORV7vU4dlPTtFTartowu2xoi4oJXg
O4IClUA5rgUa8lHpRja0860VYwLKxLWVm0OVtVBncJ8/lYwVS2AigC3GDD/4K+e3
oqOBOBxTV+7GUFpMl4b/YYOxhijtVsL6zY+7h9XiW9VecLvJWbIwYRlCKvMnLui6
UyoXZ1QGDj2rvNSX4Do8DULbjhLetXrrl+kSjuDA3jgmnC97cp6+sGMNpzpE5I+q
SMvUpwBLxld7CvfBmQ+sOaRuHETbzAgaE7XEqkcO4rsT0S8yoodRyjPjQkiTd1YN
88w5p50Hbwgq1M6i5uqozi+WLHYJsjGVgueHPn1GTp9zEztS7HbRwwKHZQdpQJY3
jaByWGA7BV7dnVkJWLv3uzeoEnQ7bIyz2SzmTh4Xu0v7LuV9SxjfMaEvEs85CD2f
IUjJQlKE2+K4RZsH53CDydr4/aFcuKNEIcDCMUBdUi1oWdOmf7yy8TQg66fgtUFj
qzkeX78zBsatZE5HMsYXAGwSnK0kUJgsL8rPeGtnl/3gIL8PH7IOoqm+T6DnVNSw
T5EkxlT/u0Q/413F42cqrvhjMCof6CwLise29znteGo3DiDLuwidliQtrjQh0yhj
Fww7Txw4I5xklBRVM1ipKBp3qYXmE0ja/t1qV+K0HvatRetTs9cnN8CswiktM2wa
S20Y/DxnaWjdA5uM1MQat7DoX4cWVIE9b9W4GkGhZ8Eql37Lup/SKjZkk0Wb9yaZ
800jrIQE7kVTjgoknoQ1WbWXQjxGl3s6FKNn1Moa1hM3/Cv7k4j3PSjAN/v2zpyc
CdIUZtlJ6Yzdsodl+gc65ep4eQlASMLCPdTszr718OTLJbBb/igqS/0N3AAnAmql
w/k5+UUiHR9ldoMX/lD0kRpq/NV+H7MGHLLCoqme2tLvjy9RsT8ms3G+pRyIVow1
ttmjQPQpUF7L6kV3jTmoAv+LCsXfSM+7aQq8OlG8u5lfMmqu/PAzAZMzDTVqsE2J
447E6Om4wt5C4qMtvG+Vu8bHVwCegavn7uZQtsTomS1pvMMQhmi7BTh1cXc1rE8t
lrfvsfNtDT4hKRqpLwXiep/fP/hsDVa3J1GVu9x/CVbcZUDo83IvVq8ZWc4vJkP3
t+ET7RDsOtmtJdNRdsXkzRpHRHXMnkLdnr4/EZ1mLRPxUDt6Gbz6hVEFC2LBA5nl
p2agTJp3eyWE+oevrXhajm/6gr0TwSuJn0BkWbCd59LWbXrjRj5Q8/eO6t+LfbmI
ie3kMv4/Wo6XJhXQkaLMRcWnd5JJmapBAOZz/WrOFV6+pdM5TcGvZkMij8pS1wGW
6Auod8/NzpydjDghb7x8wliZpLxIR6Zr8qpztEm64cWqVFRtM29Xn5CfXXJcYQxm
4CNSbj0YAr7ruifj28gW+Xe/0PCDktiNhkMpYvlVaXZmRULbJOxEu4r9jrgIZyCA
wJ/VV8Qbc+KCH720AOf8L1A72d9VwQBHW5p01Lt77kDmX+BepMnOwKalNUg/1jJa
318bEyoTojWAxEzL6xTbUkIO+VqshaTHxj+7ceKlQuiicMNOdWWuwWe/dnJ0UFlJ
CtRRYoAfN+nUFF6mgP9sGyXMeSQqpie6r3w+uTjineWq7CVM++rLsf/sy8p1imyO
C7IH+2zHFFe9GfH2haxTkw==
`protect END_PROTECTED
