`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r0Bo3i2nqgrr8Nor+3ZqjIWINGvHgc10mjE/kixsIGIsBCqVC04kHpZy1dgsPGNj
rlQ/jdzthNyqWpr/M+SiA/50ReyvGtWv8a8KqHi6a9HGzdOX2+32KI+ECok9NAa6
n7W7++8TyRkP/u11GB6c5aeAXRXi4x5a3SJ1kupgGLCzabgP4RpdRvyUxA80QRbr
Ow14m58Id3XGHsLO7T/J/PFfcA/q4rDM5vlxIiXAZ5HmSVoeM9BE8R0ETgrX6iUr
cc4QSdvf/+GFctyLdzVH9cC2mlG3hD95uJRGoDFKzf0=
`protect END_PROTECTED
