`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKxfcTzGFCmD9xIhyR9wChdIzB3MJFM2uKAkm52knbSpq9el5yV05kMj+8X0w3dU
Zisf1qZ2rp6l82PWHD2k9WSrl+skFwJzhqbKaTR+znza19YhNM6uBcF2VPu13I2r
aFMAefSC/+KF9+6bszZDj6PX7w9AnKgNT86EBOaxd447HAm7x+RwANuH7u0Fp63o
+KyHtxGtX5MRXkzRgs1At0I0CMEHKxOe4p20unvBO+nB8HOhLwQ/3TbVs8ZXwQRF
rNLrP5F7vtAwvfHeWb/6zRc4tXcal+QtmXNsX8O76Z6p8mCGv/HVzM/TCfQDKMeK
7QsyjIsM9ZRBd74DOe5PhWa0zNnisF3d6qAW483XbJbDyE4O3cpQO6iEEV4fTkhy
asTlk82Gfg0VSV1dN80crjiR84Bj4B8dWT3LeaXZ42NmgjFdOQW7Pq4Zd9EC0sy6
DEDi97JrVHm52ZADePN6XwghdvTdgsr/2EfsxDvUaDNEfxdtMbgfGLnNaKLBGr2q
G1EmegzTtbYqbnDwU48WpzD/IYAyGMzgq5a1yB7MB1IYwsMuZs3C6LjTnYvwBzM5
mzVUMv+/S3ano91DPn81L9oao7IcLNZAMLnB8k+SQ4PDd64stasgcvz1g48Qmfqk
ZdgYaFajz2x8daVdIjhtAsbmwNmJKW7e9fLaToYDzeB4w0i8dOzo1ogLNzE4MBf3
3jzTcXFYX+0bi+KaPmdc6sgUac4+8zHFdGWxDmMxQzG91X/PCs2HQJ0mweAeYrN3
vqnCN7SbJPyP91GT9kSZJJ5PzREP8xQyQZTbhPKCNRUdD4hqL46kI8QaLRFhz5dp
iVOxfGHRIZOm6CjFcZcJc46vI/NCqQdpnJgTctz8CTVTYUJyk6RaCrUoJqb2p3cq
ysn97yJS6dc39heeFWlpMpGdHQULxYJL215qBxnIapav780KyXToiET8GSlv4qIh
9oMA7gVRmb95aHzqhpgYPl7S5EMTQ8Ra8U32KhOVv+JUPQAJO/GS/VUNZ2ERS1+I
zWuRdTxKBMeKm7/CbFFv685XU8vJuuBV0/aWv16UHJY=
`protect END_PROTECTED
