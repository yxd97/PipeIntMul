`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZE2Pc7cQWTAXXNXHGp8V4syqg3Rm5siYH6B8Y+ktJht/FnDhiXFV1LKfIORS7zG
exAUSsOPsFamYBPhGgi+71GL4iHE2NG+ulCnT408Y3WzLiYMQbxZ7fwMENE2x2Gm
9Tie/Kykj0VBxhSR70AiKxZGZ6rR8epcW1PYdUvIEMRfAtmGXdfPFuqHNWKsN1RP
NCbxaqiOjkmP/hlRtFVRvTql/vbEdeY2eiARfdFe98Zswr8xVo1GgnkqR3fiKD8j
Gmwc2sYdr+8JWYDZxJrQ6Pu7uCsw/gjJpGytBmDGukubRcg1AFQSBv24MLJLVuu3
i123ToIw2/cu1h3mi/akzvWzsBEWpTPhCFOrsLF3VP2hjFRmExvZ8ufUkpSlZJu3
eTVNJTdgmBDXR3zS+GGz3ZAE0EMqd1irxIqeGXsfUXJevPfsF908h8BJ1po1wEIO
R3x3IFRD3zf6pJx4bBGCMpzM0khgPg0kJeN6HgZnyCkwFI80I0j/kBvqamxHZ89a
aCmsxzEamjIADqer/NTWDpbqnXl7H4hppkZD/6wwCjpkxr7jFQKvg0rCZ82/ynjE
uETL9LoS5ClwvulMQO7fezoniq0kEJXCA8PKAgT00UyNx5z7cA8zKdl5aFU287OF
WtzzrtX5jGGw/DjAl011yP54wzeY1wrS+djbzu6Rozn1dNUTy70NTm7ygI236iyQ
9jDRnBS67AiUg6tdM3uehOelTkIue+OKkSqFcrOwDtX3TA/dUpQmu75T6YOJIKWw
gzCtFJbAYMYcyyQJHx7vVy6toqkn+ncameaxucE8coTN0f/qcpRw6PAjB0NGbsE4
aulDeforOPz+DeE28j8BbQggUCDtO04rTeMxifThiQrB2gkNxbiCu63TLUoKYCxa
AINUferdzUNeF+obZEk+MVYZJ8wC0v9kLRr/q18uOonvanl7su+jMBzY6LukThwa
jrqA0hGoWxmSqQEtOHZSfHE6MEHbsj6++LgiIEi9YoawinhQUrgEdRzxYtb8qrLs
aqbUEH4mdeYCQRDvfSsfwrxAriZC45srhRmICE1T7H4EOMh7EpW+zZTlVb4WDnFK
x6FRm4M8P+aMyt8YvRORtcayqBff9MALSAv+xGU5yVga9/V+hDhkIfruOOJe0nYH
farRQGfEmTTOrbE4lRXEfV3880y2LuadLzsOr1fqHPdfZICxst4VP/guuvJWSLtH
nrTN73UExfx7a70k0Db4o+Q07d+TCAR58Al5w920R35HcoUHYqH1eQx/U4Kzizmr
g8A3m4sq/dW+AIs14IyiaAgR4AykTY99eW1V27nRlZwIBxZJ3+QS9FJoGOJeqeMx
+kevRsGaYtACn5k4IV38DUw/b5q5BKg+RekhiKDCttPA5jxID8Wd0dxIVmvtPf5S
jOrJajvKxvsdHVuMNB8XAS56t23I+hAZI56dGk26T2BWXRVQFlC6EIaYhMR+At5Y
AZ5Id0xOUFC5FA/M8P7CBym1pjfVSsZElfIOgE5/a2IZcy0Ah9wEy/kMQaW5kXSN
w4IRz7erjD5t7BKsylHYO29tYYN78WYQmuz/57BrjCJdqfvEA4sOY9x/JEV97OAF
ezX4yZ1GKqDyJ4FJ86pc2gWVJLf6DjB963W5HeCQde54dAz6LS3D3JWtucFaPGRm
ZVwVgrmregzQOrbO7O9L4HF3sRwkLel9a83WjFza2fRND4W2YkSLyeKu3ZAmorMj
wT5fdiGBfIz8w10SzvTr+o8OL74ieruKY0wpyknLldJJMKOAI7Oq+EW+PRyfnfVx
rbawaTxiOM53UsPxSj8GGx+TMBwQmwurE99O1NgQxcN5gwuhnwNLsezEelRRuz2o
SPSWdSGWmVjJUHIcuY0Tqs2/yETBnbJ+Gg6979Gu80/U7bpoLx7xR+7T9zZIjrGd
7XfaqnTZN6/JC7iHDIIdryTHmAlr2B5Ydgh1dNWanNyOjryewjH1tpSA+PPPn4l5
1/C1DySOmY1hblkrGYlPgC7QiGauWntApnsSgR2gMLMt3tHcWhymZgdFmquiHNqK
+afdZq4e7iiuYTFRuXV6ukehEbeMisHXvy4SLA6JHRuvva7IdUoLbmymHLmNeoVe
PaGauQQ8IoIZh6Lm+Ll0usVYXExbhW4qadDVRxjswEaMEt+sG2XG54a54uIiF7DH
nsPrbtpnE3mFN08oiSmP+HD6f5XbAgCuH76NIaIIN8CgLj8rmVSQ2Ps6avsexYFY
gRXSjj9Ish05BWlVbtFHDsV9dPvP4KkoMUizPKMDwgqYMftiE28tqtLoQuN65QVt
rSOx2//oYuRrDmb2rlpmVt8oifb3UiYiX1IMLfOCE6Ky9f6gyvtBRPpZL2Rniaax
sCXev2eS01ESTtq8d8k/7pSwZ+NCFK3mH9rdnz0C5xCC1bN3ydkU1RUBkvxbflf7
z/+2x66qBvxLkp0InQNjysP/DR1ZDtDrcQAbscPOu0UuzaQJgqzY+LjHHACS04DA
ttB4LxG1RzpIpsOqGgIomzUJci/eDxFvds4bMEDwE9UX6+WHybPkMTrgXr6BQ+ux
brIi+1XkqZf6+k5cuYbrKp4dfqOuDheWqgkWvIdMkppDOYFem8HFRLaTjGKSGstv
qyW+0dzoq/iDNQYCDtvzKkdYn3O93d/ty6IZm962ZDeOrX8+ZdSjtKMRP7K4E66+
r0M2fyHeeucAvOgGgB/d7nqM4iM03YwfJMqQ2RT3uRQxsJCV9K//SKAUBm3jO6Ac
Gr/atmhGIVBuh2TAh8QxuBohq+4aWrhCcUC4+07HWwSZZgTi3593tHkxifOv07eh
GEJFZaAg2EySYS2AbUK0MJBbJiTQBm/bcBA+g0tB8QGNDrHZo/6h06++UhArJD2F
RXMY5yw1c3paLktP/mH9Ddz6U05MhXippZ/hZRI5B25OIIfN8kBvtQLgTvL/kDxr
jPltdJCtFnN83N3ISqw0GCor9Cro7plN3NdyegFWIiQTj9yMX7eJc8Gk1qYrq6VH
NocSWjxEJKxuHkwYJ3eDNS2k7bzXznhr12aZBc+vRSeXnNoHLIynRUscdaNIx6bG
sVa51RkqOHyTCF5mLpP1XxWl19lycfujlFzDk3sNaN3ibeS90rQTWbhR+2LB6PAP
YW+JPTFBrcIb1B6Gx9xDW188Lx4PYJg50bBik0hFH9IKOEQ0JoX7BZ9Q1GIjuQc3
jPfR1WS2cJWJrwAoY1v1GbZHnLeC2rXtIWCKCR5goF11PX+fxbtXoKPY1R5qKCLf
Ti+FlazT7ira84tkBQL+AZl1WC695GG530eZUyrmgHM=
`protect END_PROTECTED
