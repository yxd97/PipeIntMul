`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdcj1WlYM/oBORa8DUz7jheok8FZZvkjNekGDT39cyeWDxwaRV6zzZftpILesAuj
1jABYk8690u/EbuxktaRfT6GhqulHnAVk3f01URt1juJXjjO5X6hbLO4uJRQPNu9
1XH2puKEexM51VQWfSg3y15VB75m8ctmDW1GIiZ6Iqfr/p6NjT1hgrFQS32sbaaL
dZRQnovDnGrFcQHYISl7O+RUPgNagZVkGcXpMmJcpweZbgt+vXmJWAWfpdZqOKOU
XOyaCGPz7HkAFxXjKTSyS+LrLqD/6r/UvP/cQqNnqE+rzbpl3o+s9rmA4M7LcO8v
oURm7HZ+0wbfQRzja9lLJEibbopPBHPIInhBzsFT98Ru8YYncq8EUm+OxllMZ1xe
46mplnqkX1kaHbgO3FFPgd4HdxFXUZmitF4gI+zUjC6JYgQH1cJpWivvZV1uHi6L
4WnjwnDa5G04/m6t8wTlgTwC5OK3m+Wh8FxBMKqEtz1ip3O2jTL8ez0jc7KuA3fg
SK3V61msTg8HMQ7haFjDH+5c1IHQzNJVWFyHXZdqVwvTQgiheBUaxcMbqDKgBd2h
fIKBi56jBWDgcMYZM39odG5IeKg8qQ7XBhh4Xibw8tfQbg/Y09oquK8qEHVIj+tx
hDyY5boA5dHOouTqi5vshtBFVrskomcU/x7lqkp561Yn6nK7iL73eppfWjbicC26
n0zDDFiISwlaqEATnbqhIbpaw1g949MnkuzQem4bOwD9Gg6oRg2tGmSKwoheP40i
VCIZrjDBnGlRB/vK9JAj/v2eyfOIMgMxG9fZywmoZCkzdo3ET+kZwGrzXJKcRJAo
DtKuPzfeaTqzUh8OdHS7Gvviy2Fo6nKsCF0Dggxad7XkSSMKS8r8wMnOFA6jy5xY
iBpaRy4Q3/7uvw4IVX+210Dh9oSqoQV5QNE1Eyr6oG9ZUj1tZa7esNVLnObMco7X
c3wre/Bt7eOAoEt06T+UTCBSk1O9EmsrKT5WG5l6jrld15WUSHWu1e0U/L/ekb/p
8WAuZlMF9onHyUKdQRfzFAmXzu19qI+BN6Qv3nkyOFhpOEmz2fgyS3TURGxoqMd6
qpKelXBQ5DyIccH6nNduvYDViTijitd1Si0BLqO8GF7TKWQYRAud2Tmlrf7dSgeG
92AKZ5VOUMQG0WrZC+KAH6+sbSYFVfBFB4jvf0x55SlMv4CQv//Hpa5S8YABk3Ko
+vZBf/upAr5Dycu4SwtXFzJTkqzNEa401AarYvsYDNDxVYomigZNewLHWlORIrTK
bRkJjKZH84CkLeFYG53mDYvf2wfI5nL871zJfr8bYFbEtRJFTs6eo4MmUHH57OZL
H0BAUe8yJFRB/uDsCOtfDfRaX/EgmCN8UfsRoQCceLZ6X19MTFHvzBvWtP4kLP8V
BBpkyAyQ+4KVjBS+YxjXwhL7UwsccveJ6zsjDbtnYeIVSLHezOryVa1p6OV7z59s
FD9EFAiLqrHcjeZSMCihWabPjwuFW8Yu88jq4N7+EJbbHgbXpjXjljqCKlgcELa5
J51exZEYng2WBI2hO0l8qD89giHU2ZjVnWWIQt+dZivJ8x2A6mtNwlQlT4s+184g
UhvS01WrHAwXCTXy3iwx80SvL7A+7qbAkmxQAXZQ3wQciKLOKV8PzXkHSqtdAeS/
v7tCKJCsH9/4b4DpQ164bQ==
`protect END_PROTECTED
