`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
weyfBdOxMk4tN2+DIuPa9+fQxf5I5TT+1Vl6n435SmmbTF7nBmFSKZcRhyNsnE94
2vCHFwkm10ZQ/OIXcb3GlkYOe16+0K++H8UEvy+7Jvw9S8Ul3Y0o9M54ise96rtJ
2aI97xIVyksBLQwmN4bvgZlttP5WqcvF6RfJcKqASBfBo/kw/pDqi34ogNJdtHWk
Ojn3G29VQfd1ESLhAaS7UmRTvWeJEM+4F/VfRmlmdafpJPgLZjj4IGxSapQheA9g
JHIsz3aiLV37C4z39rVNzfRZaOh9T1MiBTAPnCG6JWbKwLYOzxJSXjBWbR6JY6/s
kCilgBMcssBcu3qrFUWr3hM0E2RjHDPrY+URAch6/UpMU+gudRQplQX+hvlufenw
vYTggkP7/aK5Pfuup5NuuAWBr1KRQT30vH3E+YfHZv6t/5G7L/gsarc/xCG1UJpy
M++hmoohgjfoxJGCBkIQYLwrSq7qWloWUzm/7uU1QLV1nvEgBq+tImbT4bBeSHMT
VtzyWc21X6QV7JXIB6gxLamu3eaz/jxEfv0DED9NmpmXgCvmYgLUm1sQwmsrrouS
9VCj9UTDBAK37wFNX93SsQ==
`protect END_PROTECTED
