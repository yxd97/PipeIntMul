`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7VXQkl3bB2clqlU8OSsvdEfeDrG97OOM+4oNB4jj0Op+i7iZOSBI3YK/Kpw4wwHZ
LtaAGObZlbjOZ/BQIm85uB4izpQ8FAppla9Y/9OKgSwFovujhZ/FeujKmR72H0iT
0BM9JQ7+xHa33AzSbsPOR8Bf5hXG68uoFr7I7AEUTRzu9sAIK0qCLDGVeabtAYTO
Jn7to4JYdFIkwvwVHAEflLrsuyc9S/mg4e7V9svWWIQJVAhLWeCRVZUjyt8bU03h
MQIMNgnaZXS0UDEPUcP4wPO39P5X+xRn8vDelDK4/9bURulJK7cKieMKOEIqpsM1
A5s68hcVQCKWjImRhIarVgK5UDH66oGfyE6W5V/RWlmp7H0Js8MrMOgpeSuYllXg
L9d36LjzJSh1wpJnbdAqUtaOPl8mSAOXRKzRqo5zCA0d2DU2+l69ZYJgtbOE0FEC
f8oyTeDavYNZcsKIpWBrtMdpgoLnzSUlVHmlSqN3f9ft+UcF8QvX5g+v6gwmYltB
kkxt6Qm2T6G27l57TukR6wQJ81Gn8o48GtpzV401pOyGSekUaHduDWF8Lz8hyttQ
ZKk3F5wm+W5TAK+BgkyCygk6/3MsK8YRqgoJOQhYLBtcF7A0MHGvv/lltacgWN4B
i5Q70camo2okReq0IvZlpPWIiTWj0rFAZTZIuvrhQdrVbDX1O8w2iCDmHWrfXXOi
`protect END_PROTECTED
