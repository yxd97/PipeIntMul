`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luHKJE3sTOnkYaH2+nEWgCo+9QfvcOM7hqJl84tLsOlLzic1FRCTRHuQfc53crB5
74u3VWrzp0zYiFR1GIz4eLqk/E7ZFskgdjGdJE29FtRUPsOJPpZOr8ad8Ta+2m+z
/IZSRPmwG0rmb3ktXNdYUY7gPaRLWljvqL5y1FWNZhNzHEme2K+SazGH+8nayAD4
/b/OUEpOhAZPSbMEqn/6g0vLl6D3Gqh2eZllnWb6G8KriKvNW3HuVnrbR4BseAVL
lVk9JQ9KcZi7IGRthy5t4gYSbD73DjRMAe5qfzwdxEC8Am3SZ7abYDvDCCWfDK0Z
9A3eGl+Ld67Vo9AsP70gc35z6rNAu/lbZX5IopLV7NDKOUL6tyCynr+ZDuptEsjC
NgsEYE0Mftr1Q4PvIxgi0kEV+O9nJQyzNMjN0iDNykyWBXcHxM2XBPO4lLZQwAd5
KQ4ov77s1ctMtdvSAUd8NZyxX+2CzIVvD7JwZXwDW1mcQMIrL9nK2Zj3Fl91YvzI
r/dcmIAQcjUYTVlWGrNuy3McPT1LWXoZ8KwE5i4NqzTlnxlJN5tzMx3n5/dWVvut
A2nsgxs4t7RZOmCiplCM+Fzcmpr4zM3S938zr8SOGpmnvLUr/iGTiIC/PSwha5ey
rL1X44yLr3dFai5wqjxu2MLPwYjQkJR8R6fAWZ+kRoml4e8ZA19gSvz7iGbgJhbI
dbNd38cZLdC4R4J2jttdvv/RGzZHU50H79MKRuMMyFxduvdhb9U3VbazjzuItclA
AktuzQwWHxV+GLTDCExvrkaPoEh2iXYKkHMc+sHrjaXgOpX4IrE6ofE0D9k7jn64
7U0MrveM2p474wqp8KaECNttkc1063bx5stQGMOWep/9FFTRlvinh+WyltBdbTHm
Wg1hjICcRzVHyU4gMARGoUs+qerejCvmfVJQtNulVyETrtHqAR06ieh89xDJPTxQ
0iDpbVvmCV/p3oOe/vzW3L1mc5RZ38pgK/9ZrULflIi5E72iOg+TfrKS9w2TZAOG
Iur2djb/6XDgvPsP2lYbS3lmk18zk4S5F1Szio8eKUwLrCea94UnA1e9h5l00Tin
T/rUykVqTEUYoTftyOk/BiODkKl1ws2rlbqcsoegRZ/FXJ8ziVubzcjedS8Gpnub
mbxFJESNqHljn5KRuE73a0+Cgg/d9OukAcMeADG1/EEL12fvS+3LS4mxHlxFRFIz
1KP8yJx3xys87cr+ZBecK2BZ0LsG8iI9xQTQCACk4biPRx/CDq9IlS+18dHyCLsu
svPxYfr+nvnr8oQ9ydcmwkJ2LSClVrMO5WB3QahdXQhcXomIZta1pjzdY4yKqvEf
nKum+Opv5xv16btfOUmKIVMY9GhDdWN8kwhAhW/GLRTLOiptUnUfbvS7GlN9Gnuu
U/LgiP6kB0ky7aymXagxEmKa2VCPSL1R9/r6Ff0Ic7PsVZImVPfMFid/wa3MW1Sc
b+Gb/zQ4X1Oe8hMMOfPl6g7LpGhn2hdo1GeMvntVHtrYD9MBovkqf/ywN8kKQpDU
e55dDvWgwzT25wTL5+2Tvm0eXH//qEoSMq9z+6kt7Q6Cn0PcAaJgbphItczttfbj
MVvW9Rzf2dVD8/CUl3h9A8BIcFOzbqRleSnLY7ok1JoOm7V9sQr/cXY8FaUBtIBI
fsZLx/FzdTACJ0dXHGLrR5TmeFADkDz55JjArZ4Q4lCrFOjr1vcLta73lLdHIqtq
0RDChKhis4NLxBDgpi3rcy77/cmMeE5SBCWz7H+i4qjX66S78wf6kJx083/jV1yI
/kTdsEGmlS7+yD8xLtDxk3bB01ePiakTRwPCfeWvBKqNVmcEi3Dc3H86cjqlJKk2
hRPtsF0efeBU7Y+6yl0ZIG6l0CwW8whEkLcCrB2sxJBsFwiM9IWNYWEfKLbWAGbl
61PuSP/G/IsZnahXtQoZLdaNnBcUmr5w3BnH15tzcqMCprL0hTfGb3hMDheTUlM2
9TE+jTTmzwFQK4XGaHNpB7RhNT7/jfAhwgTqjjxE7Ydvwb8Yp9IPVQXm1J2jzit7
HsZpfXFuBUOE+GpAdWaZzPeCKBhhBtFAM3giRMSvKQd/Y7m1iBn9NX8rG12ReZ8+
s/zMwMpcqCvfuwLfWqta+ar+1EQIyscoL6bxIZSUpRWVQzzUrFVZsjZQinsOeNxc
YCL3Kc8We1dzYP2fxVItUJXKMYxBWhk0Sh1Ci4vqpTE7V8C7iPxHPpGzU+dd2Onx
vwOrDaNaUI6zCwVHRu7X8piQvCL/CmA0nGa0qgPWsap3B4zOhTy48WdBOX7qKmxS
xEUC/xmCFbo4NoM/AT72Q8WyZ2sG6AX0hrVivgXiTbIPuqeseEwySvWosAOVKqBe
qnSqUxNY6YtHQN54+9cpIFe+HhJZC9G7RS4i5SFRLmIgEbzBTi1DR4qNblBm2ZfP
xdTmmjnsfANJM6o9fgwVlXO1TTF9nrIJOayRu/s+9586WJFaaN8+2gPbEhHM+Evq
BQZzllZhk5D62AZBEjpg+jP/+sxz5bGlvyZ+sDmlkRWe537rwSd5j0RnQs0r3pCU
NtwvAJIBcjVtXQ+ppK4RngMZ7m7tky9HJXhl7cwDH03M1bvY6rmL2peY9b9xPafA
TcyEFhcmDYfARUvwoGG4DBz7/MFMIGic8tqE768H93O2W9yObdG5CydyaFuHYhR8
yrWckaM/+lWx1htRMOwLX+ZtsH5szHEH4kn53SKYRfTeXHVbncp8yIqpQv7wVF9u
tYgpbsERdeDtZrV/Ra6z+rYZD5zkIQMOEK9FYzVUyfr5rWPI9tJqLFOBRVfE9XDI
iohM3rk+lVbpVA4QDtStdSArNVuZfwtWq51rFHZlMgdopo0QZ/fophgurfkEZW7y
Jhb2GICU7LblsxrNS9mysu+hun1YjSYIuq5TQ06hF+HU/h/67JCJXtx/WySLatK+
IrBt0mI+Sk2xXM6tzj296NL8FkkLvRIM2DKmyhXj6v8LboGG0hKgWqOjnfGUslcf
7ZLubtGz5jzltGWnPR9537bE95qeCq9qzcgsOuvZGb2paeC4beQOEm5NKjSR4DZB
miXgbqxxS1k0i/N6rN891hqTiuoe7A9Abgr2TZudYa+ETwkJZ3NKgNcAjItCJ9iW
v0tOy5BRj6G1C0VKCRO0TXafnOMJ2SZIXX8+/g8R3VF8dCenXTy4W81/Uy6ChzCy
5iVyOiVqiXUMOZZ6VCV7uNRVwPYOrLmPU1io93IwI/sSLStYI2r/19cmq6S5LVgM
18etNRXXHQETdMKJPKIJtTiwBViDTKoY2bok8R/wYSTNCN41ZoZqhpY6Ot75yh0N
HVMi2MbiTFjy3mo7LpdUA0lQFxekdUcrLCjednPmYv2wGNnlc0LGZ8SHNpuWMvFG
MgKAc3mZUYcIttdciESwn6AFxRVE46GJlgUXx9Rm11GI5s+gEPq2TrnL4FtR+Mba
mDbMpIUSZa37Gzh35lsWVOaoXFx7Sj31uN8MPKWiB9bbjpfQwdzFtSLpJR/hNyGb
0PvphrsFwq4EiF11DYP5R8u24U+NvF39sKTQhaGGV0Q/kU2un1XAtaAffwlCnFma
s/10yAIV9eIznwrP4BKWJqVvSt0SBTZO50sWgvjcUITAYcTpbF5/HNQUP00+pQWf
MGWMKH6AnSODfIhCpN5U7BRfb0s8gMCsOEN/55N/G/n0pMVkbQ7WDhmIU5OTdMQ2
lJasrUo+X2iI3oOPRqq+I9je7mBQi8W4zMGWuX4m1vNKqjw2jqFTHrPUU7uyJUrq
9jj47wGwfI0yxFmTuWHd0NZnYDSjRoQMNAK7QC6MRIOS1D+OnzzV0s29Yic62BfF
Rvdoh74dOJD9XTomnk8BFIW1gbkH+zqjBDDQtFrW4AjXovwu6A1D6XtGcVTwaYhq
IzIKOK74OGZD3Conw+tCL8ippRZAjuWMzTzsYPh/t3LDlT8W0vm+mlSdhLj1DkBG
1X+nOWEpuH4upAY+LoRefJVGnQfvEbsGgrHtiaGhT8QbWW49SmPNSm0vpp6e+t6m
r389sclZL54K8rHKsq8lfeLsElqDnf7HwNrv+ivoFCj/nes3hCOnTec6tsdH/4SS
a2WXhQVouWZoFqUUpXTM+Mzh8j7Bn8rQ5KOR9LQLAesZDTvSK4eEJj5Djw00C1Xw
yCJmh36HBn8hcItYliH5olSIN9b9N+f4Gf/ykq8lFyJJTjZUM5JmFJj+f2JZWHpA
AOCeYgBg7An9m2DrzWm1ONc8Nlg/n3DEpO9LZgc1dlksZtvKU4EG9yoGIP0Jn0ex
iTWsVSCQxh/P1KqKuYZn5sTzJuL7jKoyrlVoqnOFs8/hseV7P8MuFnQ4weQAvKtq
unCxmV/7K+SYS2qFosqIfMdgRgR5BXxzGNrh99Q9ysc0BEYSl0Zar3XnnAbbG/7l
WCV6a9fb7sB+Zavbyqy1v4jsPjzgLM+UmQS9F0OYCMk8uqW+nprQZoWD+apn/dO2
xmyeBTvkqZZyf+2nFCT4JJjRI9XocT3nKknqXXdGGV/ZVExy4NGn5w0c8zyEFT7y
hBmpcbQvmkSKmhRjkH244EizboIgiive/+tFT/iEjfAhZ7pYdfwL+v39g5yNfUTR
ObxMMh4KoW/hspL+FGjF4l9MtOPlWNalo2Z8sKAcbB4P9ZTH8g2VyIcbdrP1/xkh
rEw7MmdnOEb5RdP24lnHA9wbll1sCkyIKGjXwRJsGaBjCth1y6rGBRZvaslaHNnP
6I1ZGuGWHNk8IMXokiHSdp4dtUMcDY3+7m/YaS7G+VpXKkj49kyiYX9+pDABSjD8
Kb7Q7ZRv+pX1OkY/LO1Jn6fScbl0tKKX5CSwBM7PkLn4pDFICYCBi5ybxYQ+10ua
hewm8IDR9nvA6K4NS103LFOPbkW15fRqq65h+sMMVtpq2CKa7bZq77VTyY5VD7z3
nVhRKLW0XvfvqfQqIOfHtKuFIQrK92BNzlh9aEvHxWiTX5xN6ciI4uZ0FGkRQo0o
qVBa5w6g4iZMaeqSazQoDnPLYFE5H4Vt9zF6ilTs7ktrzvevzs3pMYbAPKiSbOc4
1rM8jX02GWrzbWe4/V706cUtkN1u3yAzTgk7FiZs5W4cPkGVn3f72sEhNAFjJ3rj
95s/stXvdpZcYSbqYMZ4ScKNGkoKRKlttQnFpjryId+y0kuC+t+lLzgqgFyuMS21
KDFrzt/jndnzz6xrj1v0cplzDdjp/wvayEtYnv4tu4dTNBN/+rELdJyxrp2IuEU0
Fjf6AvBcU96p+2XPueqjw29Oi3rhsUzGjThXvINsrjRSlGYli6ULmApTWy8WI9CI
Eg6CYh72gYgHgdKeBXEFhV3j4SxL3JhPnOpdpTukHxkZQakld5+gDqsxb9v2vuMP
Lg1pR3P4P9vFFl+e+6CLjOH6dpjKrTESm0elpmlNsX5zLUinvWb/Bf7QdIOnbMpt
OfCY55zHIMQe6/dA+9VkAEcIdqKrmY20tbjMyYwI8C2N5jAdINMaWOeTUGqJbSQr
1nQyOabD7lpW4f3AA/g/zx01e4rGFKTIlbk3phzeO/nZ3qnxySEvjYzgps+y6PQD
M7vwcA1ebJdbhikc7heA1MhrTTVG8QvRJzHDRQmzQaDemD8LNdHZDEvqJozKQhW0
al/KHhQxpUGniVzgP2C8x3vlABRu9nGg+VS+k3VN4RHI9msVSleKSD5+ebbKeFBw
O5Pw8QdZBCeop6dBAPRis8Uu8XjQE3BJZbBkC24WoAp9nRJ2VtRyUmTnQcpnZixQ
mjEbQH1QtBFo7HiHJocEYn2aJk/43kWQurr5fwf5pxacIlAF2y9gsYEffh0s7fFo
C3FpMM4lX859kE+bJb8IJxGRWpGAJOb23/a0b85VjjLeBiydFwZ3OMu3XRk0mdQ4
kmmIUVP/0xETDACIaK2ISDiGB3C8XTo74ZInPtiHZ9ZSD3X/QbOApILtlx450e+7
JkhMFISgkPWwNA08PJTiHgZe1+abQAqMTXu7XLC5yug/CyteH3l41ntOE4/BbW8C
x7rJOAt81meh0NsENP0YK7pe3NpRom7gbxFD+CSDCJFMTeNwPRDyXTTg78M6YCTU
+FtrPI4Up2BVk+Up3TyMPKpAAU/9fIsHw7OMhNbMUG1VNdMT/vSEAGZqKhWsIdoS
5Mp/iTP0+Sb0RIFRAqZ28GoPFu9GUHcUQOFkUnefuLSPD8aH73EkYTaDGAiecjWm
H2NBGMAHeXn7LqBUGhHQoah87lI6KGN+VH/AdzriJXJECLZ+UTqgomArTRFlDONu
4pYUmTjq51mFTFbOADk24aolfPjyuHXt+7Sakm+TQtpY+fmNFlenju87ScXDI6W8
nqo2SxmNuYE4dFTt07IdoKDmNY1i73PuBAMGx38NuueYIhI7ISv5rUmVtYZBh2Jn
jlLjoNDOuROdpgXE9PtVohTtFMovOJ2MTf8eq781VrGf+680gjy/wP09Dsv46f26
w4y7a9F/4D/HarQJODiNZpeZcGK1C6/3NZX6WlfbcNpy/pJH+06n9eCxm95B4LNj
ZAiD2C2yaYUemw2ttmo/rzJBt5dcmQLRarHcbfw6+s/zYY07SgW0azuAgFOaizwC
u3FBZGYqlyNXnLRZn74pZB9aTSTdy+uo56qv69sdVsd4LwHwaDMxZqVlQP8cWOKC
dVoest4zEZAbbX1sC8XBAXLTDst8DoGiXnt7UDo1DNyxf7J/eD5fB5YWlVTBimzT
Rp+Rgn5BGie4W+dW18pwNvFVxO1KqF3AevYSTkFM7325EH43r9i5ZAktY2vT14RQ
MWDtJ186GOUjDBNTpowozpOftf1naom981NOygav6Fmk82imj2CT4vBaSEcrnzlh
4C7BOpIDE6Ga0+5LrIidLJKfIp/CRL31EvdK5wpfFf2pB6qv84pqfOj+E9TDHwHd
S2P6IHn52w+qcxpMEj6HFAtl69OHz+VE7loJtvCnuvYCsT4tonF8pTQlKgl+OmUp
kMZ/UZedHYD4zi6NnBZnLKFerUsR6Ev+vZiDKSoMyxgwH8TQoKXOXGRqcnaBD+41
eFQBuu1wd7RHEnhoaooWFTHMvLgQzoBOvO776gE3W/KPmDHIQJvk9oKz8U7xsd56
iI0S2JbiKLqKIEWMs+G+NxA4CS30tQH6gl4dpjTxDH9YQSdpibBpIDhRiHifIkoJ
iDCUIW6iY43gvNdrvQ3JXeJI6iEFiWEqa1X0KWUnQCG0x1efA4DEU4Cp7eKMODqc
KaHLv04/nW/8UkGPILSoU9kFBjh6axl+rskYxhq3zTXwFoCtqJmA1Fr3OZNFsiPe
bkPNdIhGaE8OqiOooBdSq8mCIDora6yh6VFaMU7AUmp0vx7Co8YJ2jkmIkSwKEEW
w8khnMdhZq2lkfJI2mattROsmpOtu/XZr5fKltdeVBDFhs28HI4sFCzPYzFD6pwU
9KPQzlHD3n7YioqUoL88AUkzq5BQEhCH+U4mG4OPqsTiqthHAOwg7QKb61VN7G9A
MPQlF/uXo0qdIY2O2w+tHV9yOtKt9wkyYjLzapY3CIsEemhaSukHA4B0h8UOt9Sz
7MGLI0wwnnVpdz5ShSYiuuv3H8y0bgzSDDa3ESzKdl86MWL89XDYNzMufq1hw7SV
r35VYmvi8pbEk0dyDh76cuJ6bjSPsZe/kWph9IGrIKvm3nE+j+kyAJn4hastkOUs
Tp9mJuRRiwoOSip4mQBP6AvIcr72khvfZ3EWtmDtWLQ+/ZEptpv7++q7T8aBmcFn
SI85/m/8R9wJtjdqq1XBjKWtT2IML8g2roFmPtLKGeYjocv8d1FWJusaT7iNzQlk
Irc0zb/QNrCxCG0s4gfQIx5gPM6EFLwWjtX2LzpqjXSC4XUA5ULvdPJUDlGcc3jd
ce8CMYpM35CrxjBaWb1icxO3V8jMoqGqHuXvsycyQMDLba7PtJYDJgUL0IdMFizz
k2TWKiR23N9LcuTAVV6jYQ/M8PMrkqyC9YYhbs2ZOglGAwfx2KidsvXPhAPGUzDy
beA+5ujtVtuLPPXavaX0Fq1Rt2HqGyyAO338q7o3Q0IrQz5luwYolUbR3K83c+oI
x/PRKTErmENmhqtNkrzfWJh5UKqNB6pKlXLSByRQzWC7j7nCMey/ZBXTsfns+sTg
RDsJFZ/2P76Ok4L7AqDXXf/UVivpcUCBuiwLPFo3Jdw4MIvawJvMF5CFoierOQ4/
rALBilwzMgrRuBmmgEU5ytl6jO3Qu01HEHL6jTL9x69pMeZ4SPpOX2wY0dv0013w
1b4gjnYwW8qy7W29Kwsr2rGUZYl8ajS4eu4Ga9jd40PK8B4Dd1+Wgcgvdd5nsq7A
pHlqAq93bbO4K6G0eAaoXn15PT4OsiKXzTHOc1oNJU+fnxmauUV4CbNyHjo9wiO5
vW9AtJmzq7KITtxukNSQ915y+WU+2WKUaddHY7TjtZz1TYnwtNUFHr7i5T3kquZr
eDVotoMjA/k6bPE+8qvsTlNTRpx7iIIerLIXB5OW8rkFScZ81LI+I1DILpqV5vga
Q/gHMdBoee90BFuiZK8xyor7ZgGbOPuuYbFBv3JQYHL6FPOs/7KRWmKnklU1Vz7K
mD4Cr3q1FFgtjaxZGwEP/BxghnrddsiUo9jlI9NBk/eOtEMMWtbEqLiNmPl3R97R
ZWgrsqN1TgTmOsBv3BDnpK1dUbfVhWzi8XFMjxnDSk4ZtxQP/DR9Q+r71c+BmYbu
2FSU3+fE6FjgKtFFHmbPqJ/axgG/NOGmh/0I9t+kcG6iW9DuqhxwvRZ9CP/vgdwV
byao761ygfD+Z+hORNi/2Nttq9XLAPH0O4H65sthYmzc9mDecEHXyvs6uBbux8Bo
1muNM8/Zc3BT+jezxU1fczt3LKDWb5z328iX1BKlLj6yYZEnacGBzcnDVcoMyTcl
VETRCauYWBIzDe1JWUCDRSwBSm/iHWfYTn3G/ea5TxNIDbGcHJLHKiD71RDNAfPU
y71rKUuB8mhMoDDX1B3YOoPE9OS1CyBaqGPx6lJ1LEVwcyzoG1iTsabzp8pJ0BVN
w6zp8aa4jpdVJtR8Y9huejn0sIMRG+WG2eCk9D0ofqt/XWKKtFGYL0TVTRsyUZBG
8LaWfUiwggEb+UBa3PUK4dae0dXi2pNSixG440o08+/Irq3OCH+dOMRBtK+Lj1yh
ve+2UgSk9Gz0eR37amq3klKC4BwwBNPM69ZHWwVe7ZIBYtQNTE1kipVkFud+HZse
wPwuqF/pB85sfoFnkHBnnqTJX9davKAwZv/weABrDbI9Bp/1pwHX+b1W5EtF6eOX
3FECIaas5fsdCcpJxK2WuFsStEn4OaBgOQqYfefgjWJgwCTHmpJzRvLQt3+btfRx
Jrf4OlYT5EhmvNsyIo9gNccU1GH/yu6vO35TGVazMX//uS5hMMyKKkWjLjkekWLH
0Az9SywT1D9LPI272cSlr5s+7DnUpn5O3ARLkq9zSJi51Mwb+HE8kljpUxgQKIyE
AecXAwIuVteTJSPO8wM8UjeK6XlNJfQdiZQ7OmUr5Uwyw8IMnoH1/BpcIcJmp2ow
3m1YI3BNBVHvU/m+8KRyIgAWNWWKxjoH1Femnf8unqlf6f3SbYSMYsEZGhauMIpd
LlbIA5PHUOfFZmWOIKajT6pWB4TJW7H3STo8KAV0vzB3ccE9VZh7+jZoEfYI8qa5
6E2TrftS7SwF16cCSF/9BUfmBjMGKEZPdz+0YW7Jjq2UrCdkFEirqncPY9C0qzvV
Cn2pIZfbKmf328Lt17DlfI2ADSTnseyFnP3GE5e6REh3UNh61zpFyU9oZcYJTtAS
4oRTzyFccFOtaxpOmR0Ou8K2prYkqJ81LmLydghEmr63y8+8tayd9iRgDjVXISnp
lWoRzNY1TP6JUmDKLCuSzLWcqLn5Yzth47SP+ehUNsG4TscqMb1hBNaUPaB2Tgz9
0k7er0EVHquuxJR3Q2tKvOnItY6cgXiAVLC1wnnl/61xMazUNI8uoZqiKuJyKqJ/
5TKvm+GCDyQzwVh7U4rcb3t9EoOLoR1bUodByDYoXrBBLcIXs98zKPEjt4snNOwz
trkiQhz5GF1cvWtrdHNcNhbl2u1f4DWd9uUb+K+U5E2NE0wJookoPz7UAXw64KZu
CSVoh9Je3BBuVLUcjn19r2AyAOaoB8Xokhhn/h8JCfbWrUcdpjpjIp5uMUxKovzZ
qlOQuL6BMdkFQ1WlxK2QQOulixz/7ahtuaYOC33oo+GrFseD6Si9zPcaZsbGBZHj
pyS8yZcUQhCMcP+2CzDjAioL/eC0y9cTlbc03Hxs4LMMBPAB2lEHljxZZHnVFzzh
mVYh74rEmpD6EPHatdbzzlzsoLfDrK9tsgr3xIbaD5LFvMiyqbzz3aY4T0tSe13x
rKVJBsrcuRIOUk28peVYSffXVaMfH76MlmushrnJBOfKtWk+KX294rkatRe9ns+c
iFa+gCGe+12si2CSw3Hdq+sJXQXsg2cDWxPaajJFCrsMFgMR8RJ5NKhLr6hBQEWQ
oku225nL9cKcZc0Bwu5Ql2WbBJD/ezlAvoJgeH4htOjJtAbbEpzqL2dWZXVrqwHj
sG4PmoFvsYvuzIs/KNJvOPHFOlZ+dFRKdzDRD+CQCDjje2+1Hxjn7x81x9+VlQlw
iAl7rzJOehsajxhtraCmYQYRfLGmBKWcauuybBmRB4cbevglbmRFeHCY0FHRJu2z
z6KTFZegGKxHF+qBoDmANKIbrcHJLJ+GETdShjssCEhxwmyN06zZ04Yk7MqiP7kg
FXgTwA1zqhz87QjvM0W3tA6v6DoH0ezKeNBGx4DfXbLlm3iQR//2sIBKEIslt9KS
bPDJIeel1WfjF9b60nzFSwg/DZhcYTDOni1g/XVzpOAvEM005dD2eCAFAOevoJKq
PhnvJS8kWxS42lVI54SX/rUW6fOJlqlxgEGstrv5ASFeCCa+obnddz++vcdSKvj+
dfOofXQQ7fk0MI9lb5zJ2C8HI8OeqUQB8byH5MdeOZI1rnBDAJE8NH3JpbCkSjM4
J6Ywq67oFSrZsMG/7512VDN16hk+21yIAfq/qpj66AZEXOR7giVHmk2gdQTDGdsp
EELHPp7WmAFFqG4raKh5OQQ2YF9WFxZpQEatspmXJUWq1LeXvQE8EtH4YqiV+OsQ
xSUDGm+PtzMh8d4W/5KjFBIFDLH8gs/MeG5+6ge71xiC9slSNjITV9rtAs82ICFX
ZA45SEoK92zdTcNTFmd/WtXT0NJg/Y8ovolARCAX7t43e/B/IELtFI3UXEytfywt
3nlGn19diMNRDcfGEsX/tPSf4O0RNc5BHY8M7fgKq3yqfxFORWtZtLA2xwPphjbp
1EPgQ8g3Gy61Xj41JDkqZZ5e9lQ637nLUNOu5TkS4rrqMqFGt/FIjihyDmbwWg+o
SnwYzkKkPg3bqJnEke7bd1MGNlg1nNkZ1ExQ8l1R+q5cZAK9kO7zU1yD2WRZGUKS
DUa/j+GBk52rUINAM7ZdLLZzXk23sTshsnjMBmsfWtf0xZ0WEorv/941YlODVstN
1+x+eJf9Pj+oVVIpJhlS62eJJZO3vLLVUFmU7cigzHeHmS6LXA+CRJYyQ7AjSX1R
EM2kAYa5er5o4wqmf/sAfR68ufTJkoDSwwi0nipqa1y0NN1CX6upuTtZ7njmIGYp
WoBqkB1TKCe6thZ8pA7+FNtuFCUb/9J2a7NiBfJicJP8GjdwehqmQN7hq6xHgZTZ
TYioW7NmfmstVepIrV+yR6e28iQiIpcjKCqQlVKkLxUpTvgJafFASK+5A8hwBEn1
9GQPn/PgJFbRrELGGG2xFQzlGlfkthLATANv4wN523wORNik9J3eYvSu56P45b99
ihT0yNKdw10/CHX4W1F0x37h4K3YVcFNgxwqVLfHnd4lVUJmZ2ZJB7AWQNSAT2l5
r4naLKeZIrkQGA1pIPl5z0hNdkkUXtdVAPGi1tJPaAOfhgS/thvCYIUsHLNIND5s
b6gU4ca3yXIh/wL/4lGygwSN6SXTjOhkrrOl9PQxqQB0zsavwAA1L0GbiQfIuT6U
RG7BPw6qEa6fQkP36Ny2Obbp8gTp6GLtoxwkV2oUY2iRAize4qV7QmkHIP+45nyM
eFzN+fcWeMlXeCiUF9hCTsJHxE/AwMNRZYA2oHo0NSfKHBA+wExZC2MYgyrZEI8/
dTc0mxZFmaBQv6R8HiPFT9WBqpi+2tvuNrMQA/KV6xzbUsJlVcB54kQ15JTUHGFu
BXeCopwtsIhjzRLgd2VhKHzYbPne00UR/R5GC2/+2CgF453zW6JslBFOaHocGz6T
MuCeeqh3re9i/oppFtBkGm3lCMF9MAZ8gIBZG3febcbKoR7UVGFod/nb/nZtcGiY
3MF6ozWXFBJ9vOdbeGgPOhSotYxt8aCH0OX5p4RM5Qu2gITmaBMiRuHZek/bBsJX
tOr9+NH2WFyC8V/cj9pgIYBF/U4MGMpUZbQwsZa4pA+e4DrbXYJo61KxUEHAnnXG
ubw47sr996ujjvQOWHpM4iueDWnxVhBoQ88fhcbrShXydZhgg2QPdAlDH7QvWmx9
UkesLUY2D0ihH4Ij0uXrWfEvucGapSInVZMRoRD9cK/TKFdrJGhQzR/Hjxw0uOvv
3g0aTxN/a3JwYNdIuaXzkakUUX5kpBWdAJCJGmz42NkO196Phz8qdlPl139Nrmzv
t4CSbgBFC/Ar1HGsIVBzVnbn3KLr/hXp8strCrqxBRqbFUd4+6XZvv9q/WXlf2Bp
lg8ujfRYefLQe3w6LCH4r35gDpwzTT3WKKCS92nxIHN34Sy1hDivooj3zJJw893m
5nq1Ghad0iTa28x2tWRg42uPn/lSdHdFjORe4wWURcmH2cRoXyEso8+XYpuycyTu
K75/SwRTbT5BExecccbrFS8ySUbYJVh9tU+diALhQ4shJykS7LiWLCQNlSOgyqUu
9aoMrFNU3wWG2F9WwG8m++zNVNjddhN1JzlyOk4WsWBPQ09aPsOMXZdx22dN9baD
zi+pdxHfX68q/mUbJwR5IpqRTnvABKW9B91ld89cm7drzTEBiYckPQws+MmlyWTb
C6/oKNzuc24DpOmyC35dhGrkSPxRfLctp+3ne7KmNEyGDVqpz2VWY964m+sGUl42
KWz4FToH+Cnf3ryWbnvNzTFXYovox3ECQJanl1LXQySey7gS8Q5zqggwHLWnoyGC
OoDYyrSo3W3fLI323H3tauN9pyYOf8+QTEbfTuWXRnbMdveGfphrJ41bp7rf4xbS
532GxSr5w3KxJv7ODZkCZj/BBvHWse3fUAHD/8bgbnOAm9I7IeYgCcBX1egq4xkH
gEBh68I5JhMzmk9vkhU2QBEtHsuu5v9TFryZmtjE9ISpWp4By1ky1Zlx1JE/Mn+M
gOJUJ9ioSrMHwTXkjbeLS+5UDBdaNW3uDV9c8gPJKZKbi+q7GqILwGMNCLpnxPH3
TwvS33bGUxX0v7xv7ivIWmKGLO0k4syWgNwqH3/LO1DqU6aVxkzRG+pHXynfSZlC
AxjPcyMxmMvlyDfKnFyEqf8bw1/lXLZnpU5cWUjyUGgyWWLknRGSJfAJN2uHdHHo
Y+5ML/NtrGEigmSPiy9GzNBQG1Ak7ULQv9dV5eozXsVsgZpZoI55VuXbqE1ChvT+
pimkwAaQM6CKdNarh1HiD3sQeC3ZxPmc2078YveWD4Y0z+QB3fuvWC9qHeDyR0Z7
M3L6Ut80hZD0rgHQtN1IOlqswMF+pWhp6vE6Yaz8RW4QF6xRytlZIEPY7rhcvQsn
g5eUE0OwbfA4K40jB0x17x0VI4byrSVdzT4I9YQK9gr0paWvWO1kEXidFKie3n6O
0oGSreptpFF/uDq/MqzKyVYWq/EoR1YsBNf9QI9Api4tX9qIIMELYGaj1w0Q149M
AZUeMoD/eKTJx8HN0s/LFodHINFBjoLvrWOJUBv4AgXYuQYiv5SsuOFcsGnA/P6Y
+g9S7fwQgwCS39uB+fg6k2GogpS2nAEU22Oq3PzK4zswZo2xqR9c99YvqAvpykAp
Qlyv7zOdt/q3a6Dmu3XSjJzvHkbEGgax0sb4ZJ468uLpvJGrJghseMyDy9umA2WL
NYWGIvMWfV+yKuGC9MmfgPNZHK8JqDYIcBwCk6iX5oMP1YK5dQXDvmdebbqJBLGP
hLYG+nQcOqzMI0J5TffO4jT/yr25qL/2eNtkKP1kaKXyVtj7O423VMpSj8VMBMZk
aujtE7WDqG00CDW5XPEuiVxLFtuSP38q232Fyo8b3XmK5X5NIsXKvlkecta7xesT
8ifoMImvfKjCOIhWRQLq1NICORiOQ0Jgppcb0f99ZPi0YnT/QdJlqxvd3MFoQfNM
ERsr8uA9QGIg50iFqk9/sCwcyYn4315v9WtqyXaZBBLy+7y8bYu9roXKB+te2u3j
VUhgGXUMFysQJHSiTZjmeo970DBTVIYTvIJYUBJXWcW9ai0r6lssOnVidBXv7UbH
n/L/edDBzRfWcEuaJquOPdlgmU+Uz+2jCqYqlQfSDoday1dH1j+mo6apPtc2czI6
4v2CPZsW475wYbD39iVgbtad9qcKqNNeU9Kk6rW2DvPhEfraGngNY9AfczlNdAC0
fqVQuFVZt/Ff6omyfMYeRIcsai5RwMAE9xgajMkVGuAabpB5hKvr6MJLkE+2S6d4
3JLs0NroVHOZiWePAHab0FwvkSM6byM2pYiZ550AHSt+OX0qjcbrvH1EzGSQVFRi
N2FbSuJjxnyjZdLEi0qFd8PfDZIByPr6d0Nvi11Ik/3eoGXv/LJmfRRuk2grbOxD
R9iq5ee9c54A4gWzuT1YZS3rZMKZzTV+EDdrx9emRQJfUW0tFI8ZYKAreyMIg91I
r4U1zDe/kvoHwlnIbskTQ65kzzYuk/Ch3T09nBx/iivFOS/utO+i40lPCVLI+ALS
bwUJsdAdWDKgC1SMN5TGNTYAZi2gQecu1QzBAy5lKA0ZiKkX68exC+3bI1QehdGr
hiEnyfr+7MccMHtq7hb2wEjOk+M8Go3hGVQOMn2sfOtRY+G/KYYojo9iyjybnoLC
CR1FzZDHNiE9pbvnVsEPJK1T5VdoDEoQT7oQakFqiBlgEdMX9+6XDl83+p405Yxm
TxEUVl2yTDCbQ69FJO1uYPgRwPdtOQJyojb64fHU5M9Ap6Ftp6ONXoQcXjXOrBI7
8pe0i69s2ZINJ0Qj9f2X+oqRnyxRuDXgKilZ8/XaKtGsSR753ABiTnPVVevxz8Vb
DBdhwZw8saHKrmPqFzcilFe4ANTCTW+hlOydIFLccG9gg75e4VVub6dJPwnwkZhu
g/nqAmJSMI7udxQ3NfL7Rw4JRUSU76FjKsfiXMcwI2n6sQsajGfb4aFZXLFMQiwL
VUvLCs9eQP7B8p4BHzfk9OZwc0DAtABPt/8AfUM5pjmso5Ry0KVUbmfrgNzy7sPU
6I3TyArPAuzvc3VUKkG0cMU6AqSEZMcAiLV3qMhBGP6fQ75Uvhl6P8auiQbLrjx2
BHdy72yRhNmfQSfRzkhH2xohGY8wV+7+/jqzlaxSdGUnFn9Z+7iZjVbx5eu3dvRJ
M9GqXBgvcYvL5mVVKTcbQM+PJaJo2fT+j/OaW5/0xqmu5rvvwKjoGDCNsPcQ1xm5
QBKPMCtpN72xH/2lEmM/6M8SLlU3COvgEWojFR4PvjhJ1CGQoYpd7W4Pr6HxpiQK
DWt7pq5HgWmJqc6uNNIPWj9xxa0lnJd+cuIGg0v3BXall8NB7KLw8eoXXAwqUj8n
fr5ltpDQEwvKW1/eZelHavLWwZxjWPvcgYK3gu35iAieJn1ZI4tfSWKgMFgg+jNd
5uHFDLsCsQoVOzWY6dGkf9NeKmHOoX6QGf8kqH6VohFNAB+mxPJYcsyinUwRS0+F
4HFA247MDi4qkcTk/T2nCcQ4QB32BSqq25ck40pop83Al5sOW3AaAN+xi79okOKz
a0maFMSHetTWxdkrZ7SmtWI7Uv8rkjdO3MV1ujNROhlZr4k+Tuqam1SKv4ruzgRo
XJGyyAZEgarZXP863xtp8wlsaEB3NZ/KIFuj0QqOPIGzgU/tl/ZQhqJ7FMTL/ZhM
om0lBzcD6JPq8C1r5nnVa9kE5kXLFz0CxZiQ/sw9MwDTsp0dCL2wE7ix6AoY7Kyp
N9Ldl8g6FpWuR9hxSywScbNCzuNOnfq01B4U21ldHcNSpZ8Z0qkziiivJ8A7ZScB
um9GXoJdfjM7uLvTu5Nz7Ah0hAGhMcPVbUHe/A/TE0uCjjVRwcjMreOGzICCpD3T
Ynbmzm48XEq7ah3fokuZWyFM47u5xqoQ9p+W6F+r4P/xQQTx3rNO7fCY9dkGhWLu
pUJ4KZ9F5JKB4awMk68tAFBgyr6PZG/TdqO7bSfxAx492MMCjOR43lsa4BsHHprx
FvdyDEMh0GaBYjH9xe/WhAzwH6GkEcJ2TbkRkz/NZzs8T8e3fhvEiHt5+B0Ukmxr
HUzv2fus26yxmAuByHJCRx2CUvkkIk0IAWXlGrsmtgJfdFKbfevJVXUc4Nmu0cdk
lLAWuXomjcMif1hwvZ06j4jaDikrXv1iMS6kXTlAbMzNc/nWwmBpf1ZNVBRpYdcD
pxpDlvftiWNYADySpqO/KIirOSJSw9SY8j3GGmTnW0O/p/oFPDsP7fjyRaChPFgm
vD4By9PfsEf4YwuX70aZkd9LcNHL5V6FxG7ra/2WllterAdNg6aLeCRn5F1+yABQ
X0/UymYeHelxfLQZTX4veWvmaopWqaXF76QSsMExYmypIV45+o+V1rsstulQw+kB
w7po4AimHjAL2oyXck75XYO+/EiyAxRW5PNyOWYXIktnymyj95Q++Cd/QY4GOfUt
Dn7y7jyozxBKRCz9P8SkR0YMaf+8L51BMJTLNzi4H5E+IDfCm3ROjZdk6lSH6gSy
eMpx6tbZ4qo4ZtElXnFyRXyNRZOzyn0swtK91oU4RSlMz5GX9acmyCbX7Y4eV3iZ
rl3/M3sqpJZKE5eU4Lv1ed3hIfkYEfjVtkd2dyONeNruJMHMn7VNZORaPoF8wqka
LePr31qgfZHVcD7nuAzh+Pl7yPO7mEGDap0ZAu990N2oW7WxgORCHpuxojXSoMpy
DTk3CrzHFb5SemOLrrZZkzz9GlbzdorqyIC28F6QUZlidWx1FnjiJBAQlFZiUtGs
5Tp8uxeelzTSXnlB5ueBZLxeCR8eXmimdjavceXIYo1GV2W4qSei16cHvUJqgLzg
a80XkFvx5Ui/d0XIV8RZS+cicA7RkapebSyq/u7PWWZihQEJrJhms9/wybSbseLX
jrwcxKR8BOrMZrDKXPcxGI3AkT+6MJ2GYBDi+gWuotkRRg/oC6o5/N4J7NckAEHL
LkYpL8QX4ZgdBNchuI/6hMwVET5xDKb77XR9IT3vaD7Kpw94VoB4zIomAPKQERTh
m9YKSxvPVW/8pOw4CxPGi+FP5ypn0RMv/THH0GzBiNFJcJEK3aZO/RHecoRK7tyg
PiK1w8I+jdIxTa33+tEDah9ls//28SsS4hnb4VbOyDSeHpP9wn8xnS1NZRAKpSxS
kbWpKRSG5hwcTV9tqe9JqXkCRIvVm6WhNueQZagyDFnye6R/f9HlhiDksCkW1Ou5
bl4xvhiMl+dTRO3n5b6/DdU51/yDOT4ejJXc/E8OMeiqImhCE/E/i311GgITs7mr
2UoZHkqJeTBEcaXY33j8NQd7DKfroEMcG5N09IkyK9v1oJFPigm+ZowwZHXNFaFu
mopMnTWRzSH2uim8NM0EMR1k1lILwx002jeDsTCjyju/SZrCKbXeNYxAFak5pI6Y
n3I+VB1LIW8naXnKexn2pfrg4L69w/UNBBRZDTChOxazdvpzLjGvZYPFSchMemzV
yFOxDzndd1cicsr4VZif1+PAEAYFoFZBLTQCs3HPGlxY+AIRPr/jPrsXA9c8OMYO
APcz7omcUVuFJX74mEpOt8J6dBb8zkzrM1GHNKwsLK/j40qsqvkx+SdkQOxuJ3B3
A6CLRINt1QqTTOhl1nghtB4Zmx7PIciThbdah/RBGO48u9sKUr2Ao7U+d1Mx4t3c
e0mv9ouhfis8WCHFMnn4m/kWfgzPDf81WwLdFEfniZk8C/YPQqIM9kV7/9oXldSz
VTmSZX8X9tC7wFOK7XYe4znnK/BnXc2cZfPsuH9fCzHfwiN45k2i0UUfGhfRZshp
KFmqbOSm7gTo9m+89v6nIKzQXF/rCPMVx5CqmbRh8EPWhm2fIWeOMvOCTYfRLFqz
CO5c230aM6qO4AWYC7ZkdkYaBAgYydCJnlk5ngUG+NQo6WdJRYwMU5xxS2K7dnfS
EAsGovTbFpkCQLHpZQNZM9KLYjIUVhyUwD5NxBce6pyeap5X1lHNx92nq0HKmbSM
67rBhKGZyE2uCW6mdRCkCElYJKNwZrEq4GnjBTIDRNbZCQCSSr4s7KNfoLExEqVb
QlNEcB1OFj3JzVNOKiDOl7VzG1AVxcrT23tsnT8S38RH/siSeTqIsF3KwkXF4UX9
Fx0H56EllaO+5Gyrk/4Wzm8yV9whvgZf9GG+94F/2EVwK1aquabyoHWjjRgaIlTt
60jRSQRZ5Y/sP8AKJWfXSMxpGKIv1PBmIQ1HK8ENp51ykN7AqBDC1T6hw7+okrR2
V8OD2fg+6ho1U7S5OnvAqQZQWdx5hiZAKumiO/+06P5tOcpOEgyh05+wkmEbJFd7
O5cF6B+FHG8le2kUpLZ1qr/SFreMs3QCrR8yRgQCmFlwiKLHufkQM4W88n9QYVaJ
W/3TjjrPKTRamjHDmO0PearQTy+1pSJ9WIyZstX2QjIIqw/u/OjdRO6GZoQPl25a
NNDDNn9uZPZr6EWEhrHYRQ6HM6OrgFvuH1PRhEakqcxLKMbBEhVjGcT3mLgMj9ve
QeECg5mpKG99O4P8gcaOSmlbOGtSr4ipw6tvoxNxSJTM+9MSn2h77ZuobBfHryug
/LiJ8PRrSohc9jqHdWSfdBOPWndV/3h3k1y8pWY27G1gJDEvF9Y9RfPU96GVKz8E
XnP7bIl6yHxbeLldK/3knRMFQB8PuaOk3RUnzpDLg9KU/1NM7AmJLftj0u/2ROOp
beHea3aAnRJR1Q76vimKLTOosrPBuy//kTvkS1fx7zJoCKkYF9hdLC26ZflDhXWx
vCD6yvBxbOUKn+yfg6ndQ4q4ThcaOFZCYulxLf5oLHYTSDmUPdHdzhQirfzL2AnG
DbXyNNYC1Y7ohTkyR92Z8xyo4Pb6Qs5b9nmJt4gP00euHNaJvzN3WGw8kFB+srNS
ejur6RUtGcd2reGU6gxJsG7lsiKpy7pQxym6shZaotgyQ81eFaXsBS3iDyVApFAI
HvozPucDiEVLt9Mc0J8UuWdAgBPx1/Vard7HOJ8L+WU8dWsy61AodbrlFPPheiwD
mlxvrAB7g1ex24XFxEJyuxVN5KanqgreSeg6Eh5ETgX72rniiVCb9tEFQJqzxYJW
YGucOtZhFeC/3YXCZsljH7+lfpeAiAK+QY+nI7NWd0UuUHwWirI/yGMWycEI0qAz
B40rVjLu7yZTe2boxEUcMAZt/EDSDSYzxkZEd/FK+L09hAI4JDj5jmwL8Ejw/WC4
om968PFQ8B+y4Jf0VJ6FI+F9+tSDXK31DP2hkwuiyKpWvtFG34X6WVK5rPq/iAPI
1c0yGWvb7kSwWyjyCKJPKjGcDpdZdxCl9Rp9wRlLl3nmjP1ZFeeqCuNKkiP9r5tr
30INTET8woVxKQ+aXafEEDF2AcB2Gq2iNUALU6VfuvLYfB75UE80wDM9GoJHW9pA
1lGJnfra6H3pzUOepqUaoV/jWLzEdsC6/Viesfd9HivhZsK2qMGArTQAwg8xmyfX
S00YsdIATIcbFCj6S3rZKUhA1Fgtd90sadCbBdwt3y8i/zRVOFO/hsxSK3iIbaZP
brGUrj7eGuZXglUamUZoOmHVwkr4KpQAgkoAJHmMWPycUiQDWzfApGEtrtZyh2zq
PtmuGmsqyhyK+uPywyRKvC+joL9lEADr9qn64Kgult5E4m7RrnmV+qF1/Ex91P/R
ieF395nSJ8uibeVOB7ttrQivbaorSeS3EdPZnn8f9Ho=
`protect END_PROTECTED
