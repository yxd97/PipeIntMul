`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWQ53+VnfwODAc89talyGBIn4JFydKl959a7M9w1ysIwXGFna8r9PI9X4w/roJjD
5odOHVJIM6D2NaSttNS2WuWlcW5cedn4YvPmScV6Wro2XhvpeBdKz+vjIdDQWxI/
2oZfxOUIX3gTYFSo7oSKijQMxrhoJxutrzED4zwksoz/NgpXccR6BK/blgp3HNOG
SVqk2Dsjp1+79MN9r+G4cBo00ihcbvWEl8n6jWqVZhyLiOLatiuNEV+8GihRTDBl
egf5/TH+ZZzp/AtI3rQM3noApvycJh2tVrtNpwnpPZ0Nx/wrdEsVHu0q3nylnn0T
onjwxtu3f9+TmeeWDhsw1MNovVysRHT7WYY8Ok182omda/W20pJD9O1nwUKm2Xwf
g0Kq+YI2SrwgQjw0yOAaFnaD7xuAPQd1/CSa96aYo4ttZMmjwCHFddzjVrlzGYrQ
HJuRbBR+YYP8aRcMw3loxxFz//yC91mTwFJi+1f1D2gQFTZI9Re9VRQsy31QE/PA
O0uJJzqwxYrWd41IekAD7FqE1SxA3b3y9P6J1HIh+1JTayjiRQe/rImDefLF7L35
PLslTmFnkpTldoclNd8tAvmh+9XK98mck9PwoZhldwymNyDe2hhLsj7GAraqkl74
Qrc9kdp17C8lxEnf8aFhboOdew7VA9gnesbMe+pTtn3SXs7jbQLurhK+ACKGDbsM
WiCWXXcfVIpyjjDD/qaRnITaPLnNseS1aqxak8BDFADUutZN6QjMfVf6qY54MPDX
kOuI4hKbUqQvDDvu7tyMEfttMFgI+vHijo9CLqzVq5ArSJ4vYU6gmN5dLMaEBrD+
FjGUGw8U/IjaaXQX33JagOvn+Nj2a/8ltq8WJhSeMWrwooU0V0sm87cdWBcZkz6W
OlDuicGiNXEi7Zjo5GQJOUgVuzDzwdNhxoPY3B3YZtOzvhHfoySDQHBTCcWvjnS2
lrS3KR56E7eXlYleItXIP7CQVDYyYwn4SRhhlDxqWQ7bEECew587YITIpDlWXZQk
ZXtnO3eQcid0zApEvvt7OEkb8tllVkom/gK7PLtoQfesm3OxdmkNJnDHwyn/9MjE
vxqANyAxTVNDr7lS/jPMgdSug2rkPsqznF1cMa94mCcvz9CLxOWpAFrL1l2vyR/g
P8MyWKISi0ADVeB3/Xw0ohYZR+coIdM52CGqQmNjRw2E1aZb1IMIIEM5Gtzmte2s
KTK8JCAfRQlLXBx668jOWQCfetJFhFSMk1HLWW6T4IpQndQkmoPk8P13NNVPFmF2
UGXDfHLblOLq2JPEvsgBBm4mUvq8uEBG6qyrG9BAADATkhPe9v38Hy2/HPvPSdUy
9UCYhqboiJPDsdNqWRmEG14TadiH3l0Gq+MId/dI9Vxbf40z676W+TGxMPxxLPOf
bwuFg8mM7uLrOBXzGA7RTAULUa1KfngSV2ftrnWOkOc1G/raLXQ9XivcatV5jMCE
8gquUH4o0j2cckoC7xSE9zYFH4WC7HNWnoS5KwwV8v0QQeGNvXsC2wycx2k5BGFw
w6ID5xxT3vATpQKOsQFjlfY/Deyxn/Pq4s4MbwsvxUyRf+LwsNOoO8Bl8lgaz+GS
y8m2wKhqH4zmGhWEw6kER8l2wQ+yZGk+Z/vm9+xzcAjR2OKBWI76J/eWwK3C3xGo
u5DesdC5Hr9CwxfeXupI6fkYVs07TgGPd1wZn+1WzdI9AHTNj/lKmsfzNWk0zNDk
d01Ooo7JVMAyw+N8sh8tROElKmWUBbVOVTVCpONSTNYrq3xEIXhkz8erFtkU0p8l
C3KxTTAjutfUZN4iqYC5O/b/PCJyXxStQNUxz4aqW9WIxm5gywABLkh+Y0bDocbM
zDhuSuWg8ifkOzt/9dAm2bW8MFqdUeQ48kqj71D78f/CTDeR84OcBkZ1xqQwRXVS
cJyLSNcS/6l9OHTLrnHcigkkfOSx0ncUIzJDg8JPYwvmNb2X08FKFAweLk0lhKRJ
91jM7UHFXVr67mrQP5StjeajemRVl+xsAVsa5zvLQas7sG9f6nlxBnuJdm0LZhcA
mMzsvV7ky47OCQM9eZWRlKlIfqSM/WYEGXODS4WtqCetnh6MWcEVkk6r89FMivDE
SMVbqBUMRVW8Hmr0D3+Znr+3tkJN49bStBj7pOIvsHUgMEClHgH1ctEnEooXgBho
YGq41oOn8wElCe0pg+QjaaQ5noR/lkaKjiSzxjLr5vNBX9m4KSepCiJpgzEiyNPN
hmIeSQ6/Zz85lTKsRJMNkPpGltgcd4UzemcZw6sYqdHlU1JHVjug0oH3Bp3eVFis
+RJfa2wbfZ/r8XKw8GgKOV5ahHtg+HVFYIw7aIC+XQEzi4nzSnB4SVpE899qfxG8
fprVohosfG8AJbSXn+znr0iQCBOTfE4mO/mcFT+1QOc+9x/8gVIzfECo3BrZdqo9
bDFExoRT8wR2/vvXr6t97XjZCMwxGmCuVHND4n6JrxaWNPlN4GrOgL3+RTO8EIIq
2OMY0lC+9G3m1AE5o8eyAQ==
`protect END_PROTECTED
