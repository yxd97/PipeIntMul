`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r/gScuuGrruRKf3Z45q/PGo2NTo28yc5slf8s1/rA5xFgUn7hQL64H1iWRyptlow
+6BiRiCP0gTpscmzlmo5Ek0yXEhotHy3eV8XZeTYDSTufC0rx2qgYYXWstcZcSox
8OFGIBuL1i6N6HnB/zLhr4zQBBJVntuYl2tPwhCFQTsaGH7bgzsbb5pGoeYTixPj
NOovnAT9A6WIFr1h1hGQsmzw8Hmob9Vx/vX73uzpHMSF62EROB1Avz8bIM3oS35f
3XCkUglP8Db3k1miIVnBnXMSgwt4QSPD7/OcAmUOmYP43xSd6EOIlLRJUlqIL2jv
JGKKv81SryzQAXipg55YwPUnaTzD8Sh/v3bOHtrRAUeHcLTnVgmRKnmF3+iwfD4C
OgijjMwAZP1p1aW8NS9BhyU+1L78JFnrkoVZO5fS2KjYZeshYHbKLycE/MI7uySV
JBXJG/Ws/kkmyKX4UvLnu38E1Zl4cqtscluLQlNYTOne7Vkq++9JuzcPvvm+VIxq
jq4eHACgZaDCQD9+6bTPdAH9yfgOyEgM3OHJwOd3/N4=
`protect END_PROTECTED
