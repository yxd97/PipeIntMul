`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pD3rtjRooa8nkBHikfd+NP/ZUMbqGlCyVUhLqnkxI4M3fKfiEv76txPrgLW1VIA
lHwUeCN/08SSWLv/awbrPPO624MAAkiaBoMxEujdLhxvgbqipR9HuFS0tr7ko4ts
9+MsnvikqjRiV8JlxUNeMGHgnGdy0TVzaPB5SRrM2lvt2wje0E4zUQLWPUSR/GS9
r4lG7Up1raHvbR/vQkL3HVVGtuieWD9lX4T3STWMO0F+d0GqoZCsRIN3d2/uVHzf
EBgf1i+m8BfalVzl/phrRh3hLE0yW+iFFZgBXGNEKK9kzatG6tIRAL/uJsMRqh6a
cMw9AjfoV5ydz/ulwF7XUhokLknTKZv3PXIUZ9eFZGXWhAraPZ0zm4Sdghror+Kc
um16ZsDxD9E+VryudfmQSLJJIqWA9gQla1Cer3DBnWej9PhcUjGduVaNH4ntDT1A
TbAn3AblyGYfcYy7tYrJEGfTbX5+Qra5DGsXuMP2H5Mv0C3ihuhDUQX/G6RhDIOA
UzwmAHzcJGkWKVof3j9nT85eeKoxYz1Qv3nU1SVh/9xX6XmmL6F7VdXRp3X/TuO/
DokKIvphE4peOiRxCnY4qRNzV95yZoJJkxkUSV6F5rMv8kLWx5ACWkQO486VRi7E
VwSMerq/oIjisJjJNaPkqToT+PrJJcyecTwQFDAXTO17dZdrUH9vZT6il/vXJdaD
w0+AhGcUucghqn3D3uD+T4M/WxMpCJY6dBuu0ux4gIc87NqB6LFRfo5/23Ogs20E
+SmjI6KqWSSfjp1iBtOGSTKGBR+H10MgRrawG7+UuxB3ZN2Yym5zcEE4gxWgZchO
Di9dGiQzeYhbK4SainUF+PS7gdkQQxxpbn/ZesRu1533gAOxR9Cl7d4fuSBRCs+V
JCyb8K8CVtVFwXSB6Y6QfT0W6BRvRECqiwTYWubp+Fhf7MTQYB4vl1ZE1ERRpcKg
lRYpLOGfDLz7YowVhnpje/gVmnkDkEQ/Af2BGiqndz+jBzdh/OhprkLrlT/GRkTa
iIEgLjTNfjcMaijxeicTd9qiDXuuYONzCYCP/VmLJLTuGSK0Duc0gPlkzxDSdB20
V5dW0U8+BnyOOxFR8qoJFn7sZHlAenT1XuR4qIZxX9LMucsAJGqoXK7H5IRpEfZn
erSQvGy/e1KxzSzWGz8ESE0AVgIHEXRtcbHGMpZ+HkdJHWvEHj20QmvLo1wwA34B
gW/Zia/Y9FGeKyThYfcVO69Cy7K95sEgZ1DoBKY9HzHttjLKZQpQPfLasl8iUDXr
CE9skHxIp/90EhBGrrLD19+nXCR4XosuVeA3MWPI70gtgxoBDFwNzjm+CaxWvulN
dDAGslexkCYNvcpfjpeyZcn4IE2+Lk+b/ram+qJlpKaHa5VonPXgdx/24X8gh3Sj
q/5gaoE6t2YO23Iv/0F2rA==
`protect END_PROTECTED
