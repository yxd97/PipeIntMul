`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdp86iSNLi8levbY5Zg81eRJZ9rBcU9TkE1eioN3gvTEcMTnwl+hq72ov6Ui4i3G
lMwrXko/psrjWO/+p9oNbClgJgfituzZBlvjXTuXmqsD0Tw4Lo8Ar+6mi6xt3oPH
8fEAkJ1Ko9Wmkqv/7FnnhDHUHsmXMpwslRfXHbye6qAxeldo4dfe5ZYV6uV6vonq
tot+t1JVdQEtA1PxbldeBo6nbBq9P6rI5sPhsGSEjqTteG3lhjhCKt1KgedYbVNO
ARANAZqGp/KoCT2uA5jKHgVdc/HWj0R0S9ORGp2z0o1SPGBs8XaAhp5qkvMpNPdN
nctsow65TxIeYcqm3jSHL1B6UDKoXRGAa42CS1hpl2UzjrgWRxJzWgd7bG03CVzK
y1TQkTKQsbxDOo/RQS48JaiJ5DzDw0K9lf7QqEQeegGw/CSamlBe/uRrw4XDFdLQ
XmV+nboGHXsse8BuqOYZ8P+CGqWK/FnkQD+h2cAuVKOGXWLLbnr7D6S4EJZA+YqP
IQPlvdFHlXV3aH8IHq+4fYYwEOzjIHEszmfuVAbkObvub9FfwKZVtUCY561y1HJv
9kjq2rijoqx8em9VjZuZrg==
`protect END_PROTECTED
