`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LQxZilNWxGkrNcEWIqzQiHZnHZt3yjZuDFkVUUQ6XQXoqblX0AWIDDU80MO6iXku
68SVj/EkghiOnjypUSth5LrA6q5liyT5XkoKFaf7ulONx8LRZyfpvtblGXWVl2J9
rnnKML/6KgNP1QqdiOnEO0KW41vVIiqbY/OSwRqdeBIsbTHpcBTUEz5Z3FG+zmpI
+IZI/ht75mLM5te/4QteQhu/SJ7pYq57OU/dXPs+DGFmepQRiw4ywnylbQSZYVFg
IrPsTu8WoG3XY4/XGS+uVkZ6fdDr8DdVPHANnsZ/Ent9Kxhxkr+RjkrfY/uyGogx
vt6zgV9M0QlIdkLs5+VvaSYrTuiRHKE2lw42PZThpy1VodKae8pON1n8djpkNNIX
rKcGhcqGesaOWYoHauvoAkM5AemgprcGFEVsMYVTluYAbxol0CXe+AnXB7Hmxx/s
eVAjWdUO8NT0x8spkyoNQqmfzdhllJj5y4P6KtB5lOCkgMGHKWW2X2Wsz7w2k1wy
jfI0Gu7Xs12BQ9nV2QBiDMAGWyi0fI2mx+E58X4VqmH9aAJ51tuyKA6g+7000IFI
VGukVCdCZQFp0JHkVqI1WSNX4Y2hiceBWV29PqjcBlMzXqcOl8pAhXNBbsmM1YkX
2Puu8byXzeq64ceSGgRq3/xqr0rSAWN5HJ0cRvS6kTVP/rsVQK0YouFvCwBwHOHZ
`protect END_PROTECTED
