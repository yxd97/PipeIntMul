`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Ns2831btpPHbNTvHfY+ujgcODBXsmm+QVvjW+G/cAdqhkEWRb+kVbqDVKBCJDLg
QL/HoT8rTQrU5hL6a6Uq1MvbeAkuhHI0rp8kaPUVE76JE9Hot1rpWYTOefehGkcO
FVBEuuAhZzfCHjQi5KKc9a1h6enGesxUFHYz0DPm2XuqOjmr+kvWhy6tAFxw4vCj
eCG9JczwW+JTxOlwpywhT4lk+ij+QErlB6LIyQBjjb46252LtySJa/U+/Is/zgTS
3yUXRtrEDMUvjUNJVN6G1ut2mjeWCKn+e5CrrNZjbK70ZzVBYjhQDsUcbwv5K2NN
8sXG5uJS0zHmHOspaRVR0TX9q1umGH8ggkCbwMw3SVdavvIXFd0amR3CEaP3hAbb
`protect END_PROTECTED
