`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/gPcsocDw+3idzg2mOo0eVVRY4ZzeXRUmpbBdrFUQecaRy1uB0m374cNIOUf14Q4
cF+sp0b+WtZ7/Rza+YBvwe0tYq/keJ+g6Wi8rUFDMc6v22LnZDBs4tUvYMicwUzd
AFkRZJQthQ6TmWTKLnibxGtZXG89tQPft0GlxFw3pRrtcQjndQib6SPbc9X7+wDV
7u5I0hVx8jA4J4BPr2OIwef0OOG4UsKIm/B3VG1KNrSLunwtnyrvZvwdYIYTr1p6
vcB1tifE2udJ8OR7vW3pwmqn2ONiDbO6r24BsgD4IDF7i4K5DKqyynB5arCNKPdV
Ksv9rEsgqnunPP12CjoPtw==
`protect END_PROTECTED
