`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHrpiWxzHxykum25hudoiiFVq+kRx9NtJTpb7U4/IlX/HXoFI5bHh1T96juXtQnn
KBie0//hyB4JBTILAcJ8Hsp7N+/LoWdm3KTvJm9iQmLxZJVsz28hc4yrgWginIhp
50pZe/CSLyMaNoxZnJyXiTcaFrQx3sq/eRHn/ejEziohFNQbqjiIvtHgWv88dGiX
mnL/wGI71X3zU4kvsgXW0YqPyB8voKIMWaTmnP37TU1gXWRWfbXzWmZMlhctkieO
ZpFENKVaCXmmEU6Hv2q+z4ZQJjf5JlDgSA3hguo5KcdwPsa1VKQXFQgzWj4aX1o7
X55cEw8xrNFwjGpFv1WOiyLCPWcWefjOEPzyA3HYnzA8pSdiULhs8PpjKtV4o5i8
7u29/6srToeZZ0heoNL5DzY6ApGUnOdtX1zggyDnhwU=
`protect END_PROTECTED
