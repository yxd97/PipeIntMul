`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WLm7hGfJmqPwdpRH6yDPbOiYRmhu5b2XslbI11k/oRdMyIT1Bso4QUVjV/CjsCsx
nFIp9406bLBGjvWTdhWQ1x3FwZ2rDMtQOoTe5BDcuKHNDfNpDiBPCoMApstgfY2k
CfwRM69vAOYLS/hrQtNvjSRVYz3xaHG6IV52TaO2QUL7Kd0foAHkjQg64Oi7LFRc
iSIA/eMiQtcHg+eQTi+WwLYExTrJPetwQKxzdqo3aFsoA97qXmykEuL6L61EvHoQ
3nn1v5D2fij3ZC02Bbe+ggHmos+GCfPpYV3C1hi6uzSBKen8OVbp1/rBTzlhT1kU
+yb9gvux2/npBzn9PfInhjxhW47NaIVIR4jFNGXjZxRZ7t+51Af4BvHJBEVGC4DY
N5D0B8mDDRtyObRxlaIN9T88m80Lhhg3Gg/LvzIOZNXKMeZD6+OS8YerOsiloaT1
b2CKssuANTSxV+bI/mRzDMJY14g5GuQqcJztbugc+yA=
`protect END_PROTECTED
