`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oqEF6yKDQD49ZjPSeEVtphBsH/pbWTotWvgFzlcvphdtztZXFKtyWEawSqMMlp3W
bJk0Wfn0tkl83pB+jlvrZgU9EdszwHu4MO1XJBw4QXygjfbnbf6FZUO5SYIBplhN
1Ns6i8y03NTXe/4g4cac4ZYOEKczo0Q2Yoxon/lztiH+T1fTEm3vnccAuVNDpV3n
EtwChpg6nImng/QdIXregggYl7qQFcLQ/uIfDhjoxnlNB3w5YQZGAqIOI5kQcpwe
`protect END_PROTECTED
