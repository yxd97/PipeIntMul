`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jTo92mr0Ic9t0X0nTS/JgG25YBzuAjBF800kEFFAQhs1AufCR/OsOGJ3fbPIRDdd
Tx7+BJPwM+HTtmu+yy4lR3uPlCLaaL4fk+gCunKLyuyUD/tkxJG/gDWUcwpL4HQ8
a+1J4qX5phCB03AUMcWHcIRr2kv/fnbPaVlYG4vtKbWWprzmmZaU7wksclBRyrzN
PnIGIatjb5F4nK0qiQ1bqDQXMC2x/Np1w8vdXZvh5ErAtrxZbxgwwFPWnlapwAzn
sjwJn5CIHe0g8ldPhchqBQ==
`protect END_PROTECTED
