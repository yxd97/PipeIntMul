`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EE8Z9bTFQK5Enp/wERhuvAQobkM0g589PtN3DzwNDiYnGfn4LfOwLIfz06RLzX0L
TRTX2yQnYmJnuTCX9ueRktamhtHDT02cSVhqz6wHkc6A3JishF8NpuJTwOInnwI8
0EoFKL1nEZDmvc3wpNqaVG5D9zycOK7XFYcwGJ0x0F1yNw05iCopM4uuZBR66A9W
Exq+87+n3GLcS/KRuW63JNhUwcCuq4mx3KN+zwRNEPWeBnE4NbpZQmP+agYGahoz
bytSfWlwKoCyEC27H3eibS2Y4rbY5tPllbh+38iWl+Bs48KGBgIOKoxblI7Xy+xU
+Mk3v+lCAlP3REbF2coxd4SfFRQe0dUb6mVgaJVLybLniYwYDN3BZ7UtCPTW7aBk
+3IWBBAGCyNC/CffZlIvGqPeXLaX449/uipTbbLx21VKShAyc90HFtR3806t37ee
dhfdJLeIDDsDqJaYRI36pEX9Ut9RTnFidXObjfUN+kU=
`protect END_PROTECTED
