`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3XiYtGRxRJ2WJOlej2+/7uXlEBQAavIP0i+CAg57+g8BF9q7wan46V9ObWofioKx
8tvfZM2g4fjqTag8soBtgQH/9s4st5zS3RIh5Wm1BmhKzzJ3yjzBr/n8K8dQdDFT
p+b5OWoHLm5iPJBTMNZV4OygV4RQPUZ+VmJGMV9vArnfNaMPp8g0EpAjIRJN5Q4R
C7yGMW/o92i1Z34+H72KBy+4tD47j5mHxB1M85YQaOwxIsC4322GKKvlnO78zYwS
9rYD7Z1aFZWPA94sjeP+uohV2e50RchDoTPN94sJUTRaqjN+NfWHisSrSMRN016q
b64OxeCOIP7UvZdOQUWcr2U9o2x9oTkWja5D9C+Uc2koom/AKfd9L0QvgMLBhCnq
D3uYL7R6FnzGUjEfi0o9+Jvi/bS+P5bk7WpzkZRO2kbBTbCkXmPybGDOU2w26RTV
zD1W1FmnIslihJgoTT764pLTa1qcB1APSjNhTvGKYIqsYQilPs+/x5762HmE90CC
r02E9hQGa5XQBVqC6tuyV1sg7v/DO9Pf62bj6deCSvLReYddoFNaDaCtajACDUTr
iWY1cGfap2Pe7E4DfPNjSO/EFAjx4C2FRHMVI+WQDnbeKcR7WfftM8EMwEJxyjo9
8m9r/zIRxfPl+RHZtaHrBA==
`protect END_PROTECTED
