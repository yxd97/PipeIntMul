`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8wHgJfrRy08hRJCW9157oFxQKD05IZ7NdtJ/L4jjCK7ZlVFIT/NjYohVFvdjdnV
euyv9ULk75yW1yVo+OcorpIoanmy2GhNJPNjZ7ZLkuhOkp8hlTMf9PoeAm/0uCQD
jjdLfDdmxC4l/OlVW8/3OYR5bym+I9MdQxsgAAQ6yb591a66LUrMFutkgQ9hSrS7
ncFwEz0chHOPEw6/iaycSqaJEAabQiIEP9szrDLVjA8ESDsKYcQbbIQtky8sE9lQ
lonOjQVENmymRqzyglauaiQn+mdF2ryKx0x4l7QO0AJSVfHsBMGTqFMlzZPwqQgR
Lgse49zV+VlUSGS5reeKzE8cPmf75qZ/Fw0EKR1QDQ4tC/d5EEx4isOpbmsOKS9N
HB9TDYsqlsJc6rZd23RYNvCrATrQkm0gUqoUWkeLa+a87QsF8erhKr4B8Y2rNnrJ
3l7j//PLvOdseCW+ains/5FuDa3LfHvJahWMruWHoodTVMujXkHkF5rxOXsyt6gg
Qe4EofsvFh60tuRgx+Hcbg==
`protect END_PROTECTED
