`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwueEqfQgi1pBPNJemO2/IgWd06DSFB/gS41os65JXJJbyD1KHTQHs/3eeJX7JbG
AoGlFUvArbQuxEcpgQcqfC5Av1JA3sogK9GIABQDQrvhuqdRz9VO1H3R253mZIbn
jXj2wDiCLqFusnhByEWzf9/wtgCULWotD3JMW8EakRhEFJ2E2L916iYHQe1CXfKU
AgJX4T8smN+R6vhrU0AhnrY1s0Y4UCZ+rsLEv0fm0R7lg78BDMKTMHoyRAf03wA7
zCTT3h2BHFoIY2Zx/n8mC6TYHpbwhaSr57foTrrmvrffxoYtxlpx9PHPuTjIxqAE
Eki5/lp3LwHlyjFuw/jhf+nmNuFWE7sI59DoEREWpvKzJId4xRzldgf/LsYjC75q
reOR7CaYYZsiuvYKgwGMbHLo+PKtjz9OXEHlZYmpxYORBC/txWt5Y8SOHQgDldRH
CZgAf6gqP8+PV7xIM/VZyT+uIfEzmW+hYYpGHpko2MnmjEVaR9v7ui5Lw4d7h9NO
hb2/2l3M9CkyGGW8epff3myDE6rwh1Sv+7ylnteaYVC48kmOi1iVVzD5YIoK/f00
064ispCp9iYgYwHTTCvLWepZtxv1s4uTzubkEnzjUMAScq3caDRZq1KCIbgsfoPD
WwBrEx/mYUYseRYXQqMXUYFw2njLpvNZ673PbnCJPspTCnN5v+rT7ecBYAeOEJ1F
e8i2WtdeGYXPVQAQZQ1ye7gCbqGdu3x7igsTZKpkDPzyx5FkdJr/vbKWoRCbf0x6
nZ/Tltr1YV1EF3+YdnO2GqhoeJB/QYFcpgtmdnM4W5OXAKyJLRQCtOQWordSchxR
PCZcJIxtVs1SpQz3KjuxuFCBEds3WsG482oO85WEqE3zkdw3OAuM1q2QAcmAapff
gGdfT6n3VfJL21m+kutdJRIAi/pPCi9HzvMXEeV+qj+EPcgcJoh8F4xfM5ZfvI/X
aSVU09/WKT5mF3gXUUOd2/PV/EWSnla6yJTAfeoKjczVAE7Vj9eeXOHFho0WiV+I
3DzzaKnC2Bcw+/eR2CrRiDPbxm4EDIDlV7NGfgAZEMku07NnFrybp8EhuTR6B33W
vcdCYcez1O5/mdJRCQ0i63H9fFwX8rnCXp5be1dPvJLZyeesSfxt/n2fgcfm4IAa
42m/8cSNTLddE+aSsKUoX5YlAmMIBInQ20LwYtWF+jVQPZ4LejNsihjX+OiUKwSI
QP+gqxfmUQxc+5YqEy1sEl9V+Ut+m6unQmMYkO0dKMaGMHlRgBWzZDoOyXIn2qEd
IZYZ8ccOFzgaqWaFGZOkhJ5RmgEXdZSDjLm5TnfCkJuefkMGT/y4OKjFrtZxFVJ7
BuYecc3c5eb4vca5c0RyBdnFhVXpAvXbvGh4R29QaDMMo1S5IYtH+WU5U132R7VL
bKjB3Sv7HGKuZzwyqFMoso4kRBY9fW9YehXb7YXXZgqc9TvsiUIiEw3PXEH/eNfi
jtfnOL8d0xMMf3lRtMA7jOe2+N7TGY0YFyfAmd1IbhcEDR1VoZPL1BIjwFZKpzMZ
CCQ6w7JmDF/Bmuy8NP7MGLpWZb1wRw/Z/S/OrQphukSbOMcKQH/MR4rgv8eu7Pze
ZnlShYysVU2vwFN/0CmWNzA10xrRoKgs2oFL5mFkCyf4i/3m2YRknF9suufQyRLw
`protect END_PROTECTED
