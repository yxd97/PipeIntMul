`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PILpiSjw78cvLmGn6OuyaovDW71debe27bYQr2ob66FUWl6hIdnaqyutvq7xLHA5
n866fv7H+9mHgxx5b4cklyeMNbIfdrydyOp+v9FbonCUg+Rcj8ikqAVdO+fCINPt
q0sgonf29DaIi05b1Iho/KgSEN7ZRLONQnPUsuGq4WfJZfqQVcn8Cmynkatp6uIl
3/jv/sMS62YoKt1DavC6QfmeBwLqPzhhFZ3TwAgx5il8caNUmd/CbuH1wA6rhScY
4fWb/bwiaaXYHdfsNKT3ZuXEOs81OGNCHDzqg1kCdAYjSeuzgpu2k+vcqHrG3g4N
w04GU/wImuhF0UxrnpmO1ItxDuB0OoKygg76ADTSQPXtk4W1bwSHvPNcN48gdX/N
4gL3Ud+GeRTUYEYGudtA+JDRsZA8saPeppgcHgzno0Q=
`protect END_PROTECTED
