`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ds6u5eePBLKAdEmDyrZTcoRLvLCy1K61aCSbJbp4bFnOMV4QpXwpdj+0sU1UQOh/
Ug/GpiWSf27URXqd0z+BTsk7BJ34+imQUJacxt1icjjcv6cYEsuXKn1BciDnEpjN
Ym9o+5Fhas8Mgjfao8Kk/t4jmNxFTPAQfCQKR+JCBdhxDxZsa5wLpCgRrxkVA2Es
//+1lQEUOANtuil7HU8kk88OoUkhZ028BF6VGzv4boDMNmGlBH25B05NmKunDF8F
iupPnULyAoX0fgGxUlLVLyYk6iFMKFbFovN+2SATRR0pAiBzLOXMdvyz2ynIoJ/h
eRi/AAvUCt2k6FKQPGvc+u+/yWmvQnEKKeqLaucm+2wcmwS2K+4aYdi0nRV66lY0
2rykWUvAlzUO16zE5Ob7FposCxNVHdS0HAAac4PndBWNriW3aoqBNLZEsYSh8hKB
`protect END_PROTECTED
