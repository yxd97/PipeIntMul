`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84I5QBIQ6DCMg06gmSsrGeICmF8PNrYhnYInL5wDm/4Z2MaPOezUOQsnU0RJgCyi
Ooz77EVQ5h4XSWXzTjSm9w7HoOLVk0S5vTmFIAVNT4fZE/0z14kJooUwaZNNs6Yq
YVJRWPzFZcQRqB0azgCmeayZc3OSHBNgH4Ale+cqCbf31YKWGb3NuFhtD4IiLpi/
Yrv8+nh50mPPxHqiBBD4loSSYR6xPphME1ymP0tuYmDWHZG4lF9l8E/XddMlY8ub
iX2ny+8ig7IBYAaZ9zkOuranrWmGvWTf/0z6eWKqoeYj4v1Xrisz+XUFzTC22Isu
wHyKPqIDVzTOxhrBrOmqpnRKAKW16yuD7z+uSDJL9aXnuutRrFFFc9EsHxv31kBQ
75ABbSzAvTNucAjPbH2MgotZNlWzf7GXdp1E4GPHAePWYz8A7+/ruaBQCoxxPiOk
`protect END_PROTECTED
