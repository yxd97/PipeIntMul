`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gn/mLQO2JCpS6dEuGCD1d0tNpmuv1hJzBP8OpFAJFU34fFZ0Tv4uoYpgAV0AUH1t
hNgttu1FK72M/SlqDeCgZPrDG9i2UQhctJ1+ANUfKF5cRpt5cpG15pyGLODiX7b5
McBzWKQlujHGM3pi263j0oWiInK+QMMdbTG3A35+nYPzXRU2AxxqAs/3XN+klQVB
cjO5YJJUtB8rFXM9omxYfI7ElAvDxv7hDvxAKjSiEmi8LZQMU9vBwK5If1zFEdGQ
gfIkW+HbYDacrl5hjRJJho8z4FxayC0AqbtGND37xyLuwB9A/ZpGhFFP/LBA/q2s
ZI4CExXVRMyhHvreiAr2dljdNgBxYmzDp6qg3HQsgWmSaMCOSDMf//DritECyPLk
keqqwabI+PELI5QwKse4FQDs3dfzPgh7pX64ePQoId6kFfJKVmsJWqEnngEMSc2S
z5lV3akxNYJRZhgMTFxHVqh9d8J2l3is4Cw5yOj1z2W8vFo8kNpPk/RRm3s8tgvl
uHPc15r2BDMqxwLpFIwggky6qY2LCTbHCBQG+jwLNZ6PvzMnCY3fwVwAPqZ8rN0x
1dZLGwA0LgUEbWnbDJ7uGkfMW0VhpRzofOc0Zk3p62ie8wdN0yDJfLNH7W+m9iuj
CzaGBpKP0mRfvieuhjJpAtafVVG/0FDodbSG3v8pMHRyjN205ybNk63X2r1tFY2x
i3hZpWVHkIO6C6nPiTBcGNmgnmJ+wjWPCEArZV5shi8=
`protect END_PROTECTED
