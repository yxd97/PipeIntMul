`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z46fVaraS4mApul5Fr+reSFc8hcRNmibn/iU6Q6EL1ytRGb3qRtDBsIgNR4rf9/F
gCSiGKp9fCgYPC8uXzMQKsp1iqJZqLLSr5wFpAYcWEbjXK0Bzqrj1DfoEIFPgM5R
++B6XZsdP7YiCejtEkyYuxxzbvje7YodX+86UPnVdCo4l+mK+uJcPK+x4W+1Hf/+
crv8mlBWWmYfDO0UmOfTAlmJUKvoTMgSub0PzyEXzVp6E0pKhJjaR+n5rlq1F8Y4
dqTAMvSWBljeLVs6SGRCTkAKKAvpijiIg+Cz5KLqqvg9wH5K4mmGsCUpQ8IlxbFp
M0V6bZ9W1tqD8Vi95m8XBu/GbPZLMfeGZqEvzaby/MNYpmDWLc/Fsoka2csxjpp/
fSVoDsfE8cX6IES7k7cw8uLOuB3Q5s/Z9W3yXN0R0FIFXPdQx9HzATZf+AvDaJeJ
eqaE+GVk6n96FA2+Ao7cYz5ZkeTXEqXAI7NzaJNahKO/T2WRRGlRjDEe+JipfUqI
kiVL1GuMRPrP9tNvLA3s3In1sM0ntYAhOID7vciYLeAW5Wn5rkmMTkI6VVHctYnR
f/b4wx5+2d2x7eipRoJJ8fa29/aGAQrBUHCrwiYre3zdVlH58AwR2H82MVn8c0fr
w8B/4LIBJ4tTSTTU4mxkIA1HTu5ZWZpyrExPoDNT2urgqT+kG9qLvNDQy3naRfqN
DMl8Ryslvo47DxtExMmmTxQikW3qF+8KNw97WcdY93pHpAH1epUNj7UECGADCXil
sQq09LvyWgsnZJpRs1qZWfgCX3LUpNf9Qpu1FCmU/snL9s+ebSGWkGE1eo1ng9Rg
DSVAloazIC6qMKkItPffE4rVm37AhCtvTW6fG45tkQ9NzJJTre0gr6htddylilRV
Rn1TJ2pm0AvxPc+mvyD/WGh+VUW8zQK1nEhQhjc9GngmloRmehJb7m3yQSh5SIgB
mPnhbJPgoxzAVJcUtFUYpWg5yGrS05JCEgVrIgJivwxoLYBkvCLR0f+T9gn4ADXe
e3Ltz/mLiiaSLp1ZAJPdyDn4SVh94oLiEIrw+4n00173RxDdhdVon12xd1H4nmK+
DEaO8cmxxl6M5ZbW96S5dUBIJzqrv654IAMk4dMSyuO6P9aFXxR1A0k0IDq2z67S
C6f1HyvfaNuVJrYIlP1vPC+ikj3+orYqVVZpNDAjtKiJqaayzV+ubDeXAvSR5Pza
tY5TJvEGTKYgkLCduOIkRRzHq8DDWM0XMs3CAIW7k+zZgwMLm3WujwtdjMtixf9Q
Nw61CFAb27HRU4JRQuA/UeFUqX55oYWjRWnSvuiTjFGjzzz42c2cN/t5s0kjQ0w8
1plg3cuE3jWvx6Dt1wFN2ZeA5gFQLJiWDrkIGVWesYRjBpBM5tLrnp3CqvZJTn/n
Oe9o8+FYJDmOcrIlm+gtz1bMaZCXHHNbP5YU1swIukfkyJI+fP7akkWlmltFtswz
Yf59NyNxFw43sLuFSSePxQt8u9DJAD+7zYB1okGOP6rwb5C4G2E/EKf1Ji8DtFvF
4WpzFH15x4wF5oajWLcbCed12/jw+rBHyeg5rvfXRjFiSZWjrXRkP4Ww/sYMwE96
Iz7Nk3M4Tv+56Vuur67bRqcpa3rFzzlC3AQ/Nb2rTFc7Bn8EcE6Z4waUEwrkqDG0
QuHJOy9F2OLzDuwZZioaiEfe4emwcn4T2cUdpXyRxIzYQUYxPg8Wz59DkM7bVKY/
WIwIOxrX5l+Pet+Li9cUxAh7DJBrXNmliq+He8RQcjWlvkS7xnEH94a83WgmJUL4
ykL1uejkRU4k/pNGjG7SD1UMrKH59VMYuqJ2duCvXavpMIqfyJQyWkUw0Ba9uCKc
Shp9PTtSaV+ZqyLKoxwIjlJ4kFFregd6OLBY9VOHwVVPVzM8QyPPhNxO+WJb0nSA
aKFb1Z1Ee+VkOQ1UCvZZOD6yTDe2qohV+52vZU1GuqrY2dKkNUFYg7OR/LXFqezk
S2IaSnantKWv2oJat22zNqZahdjXhLp84xfSP83G7PAZOdH5vSfMBuTG27Bv/J0l
D58N2sYCgutAioK2fHcipUkTQc/2klNCyT30/zAQah8=
`protect END_PROTECTED
