`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JOLPk6geQyyU+VYLnDb83rRmEl+/sHfVurO8QITJygzOQ7VwdW6WH9okctVWgLVV
xkAa4bc/J1RvF2AjgJZUBwBX5KI+vVwqosRcBycEuosxxjQhezOBendqnkz+6R2P
NzDMlHUbtBKEvo3SrV8yV0l74F6Lb5paMO0flmDo/jaHPBHbpusKUMVJ6qnNNRTx
tkJgPNSg5ytISW4ejGaWmLVIIogsW9KY6XvomIB6es+iLav5YDkTszedNw/3k3z/
sddojouInZc/Lq/PraeckOZLd2YmxjGB7OO/zcO1O4JOGcJOpM3dNZdryMigyW6J
A+UMRapYbR4hwWbMLa4DzHwJcRhd9tuycctYn2davLF/rjBAXSb2S+boixalNzfe
IDvM5LV25h1oZXGsUemLwuNZw5cyGMF0uxeqsa9H1ZVKtpZzTPe4kNn7fv6s7Q8K
DArA9k5JUt03E09a/v2dKD/kYLMBCj6nJnsqAeRzu1uND7fsuUneYYABVuvc8ZOq
rbw7qq0vXJuLqi80ClV7CAF7NdcFfLZXYJJtEG5WcsTeybdGrXCRgCGLF1G8BRA1
cQaMh922Ux4BD8rPK2q1MAHYn4z7/QAe1YGaADfPKv8KdUveEbSCTIl4vC1EvYRD
cCYf2qnDpSK011nqYkVv3oQWbEPGt7ADAa1Srle9t2a8fEB7r7NbwzvwJQH8trDF
RFobQSk28FDakl/RbBmtgWo+iczWp40wlDZ/P0iAqDXdFwffwEf0+5sYf89fPiCV
CKT+21l8O3h5KFyrygxmHmIJTIwQ/sS24AzNTDVei1vw4rGf0nRgZ2k7krqe7hx/
LEt2P4BAkeD4Kq+14Jrd4BkKs5YvJePAWuQxdErRkbVSqRzNb6gZxOMfmw8FU1sQ
NXFwuIOnHMuFNuWSV0+KZhscedpeYUk1a/7A4PhkGTOMLR1gbfDa7zrAljn/uzjH
`protect END_PROTECTED
