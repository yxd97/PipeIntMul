`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DpcsUq5awk/AsA9xCnxSylkyllZOZbZvYIrs/OjZtgK0EWD6ta3sde0D7uKGJ/UL
I4+hw2PMo5xOAcVQpHYoC2F+JZVrjbCKVQAt8ZAZc/NqdJgHMCl3MOifRejmIGFF
DkS3R1ka9fmRNKPsCbYQ6mjp66SI2DN0NOp8rYRrkzzRb0oB862yd0CkYV6iG3hl
PYvaPF+mMIjalJfLclBgt+fbxh17KThLhAhqkKAsTty8rtipxwqqP6o2VBalbfXE
EB0boRgb/kIBfODiBycqf7MYyIn6xTFGiH0ipsgTRT0=
`protect END_PROTECTED
