`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3avMuIh3JP4gbOX7+xAHK0eicUnuTHN3pjuq35kgasrDWxfhrQyTCxElzUdLiCyd
biPx7jt+e1MdjA0oXOEdAf+yuTGrUOQtyz8RLJaxSik4USx+M8Zmmwt6fF2kIWrq
ox75hL4WJ997/guCnFn5Rnne4yb8Dm5dxatjuLeKzFGNrNRy9wm5PsbvQeHozxVe
N7RVNK8PDKe/4cvoszMh2MD99kaj3FMI3TdegSvjzR2W8l71HIfz0fuV3W+48Okj
2whitBaHwJTnpSu+l95rSKk+gCGO37QwCVkZRg8oC4lfGOsNgBHivk+anfLJg9H9
mUXtLAJ5fGbYfM34UQqpSMyphG8K5q6Xve5sAegmcHTFd5i88bDJninKUZK49gtS
dIXB6taArvLPJu57fxNuboNj6mWcfNfnJef0PRsSrRZ4keEe/OUz2x1Di50h9mnv
`protect END_PROTECTED
