`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRZ0M2ZGVRSrtObafn20HTcaa1s5Z6G/z51MtCTRdlhxwvODyKxBLY+sNYzqz9XZ
yGkhk0M8go9Ob+0I572uZSbLdtLNick840VjcLJXb6dRN+ws5uTS8dc8jH5XfcfH
wtchoP3CiTS8FsUb2fZ1KrJu1Mf6rV63BvzclRJAWWtaIHm657Bf9gIUZRSD2Zwk
gcNXAMFaMuBk/j/ylRKiFLQJP+4dRiSa6EWUa1ZJJzLSC1ESpLwrw8Sz7WvI20ki
Y00uDExWEtPvATHBdvjgOONU+jg0cjbuVUBpMwDkaq29iiDczOrddIYMQAsT9vDc
mXmdE63nf9XPj44yQCK/6gg79YqPB8ELlxU6uJab8fk25QnQB5fSpsCDmXl9sO42
Oi7QJLPeWUvATo4vsKSxQsTY05HEoc9Sse+m/gzGrDEMfsqh06jZwF1nh1SS/Rue
dS2ppZ2xH8U8X3AVbXiPSJGKwbE19LU7yL/hV0/ekFazfleIvc1Ec1xFYlonC3xy
u+W94DjL4g+YsSwiVLuLd90tOhwD48ElZYV4SOOZ/IXqa9R6WjCgxDPKVtdK7tr3
XdVolaPxGasLWlImlMmVgp9CVMgyrJOmMmPr5/LEu1p7ru3cfBJtOGJxIb2Fil7M
J2QllqdvISeerlFs7REi9rFi11j1yL825JDx6TkFapRqI9vpTdqe+yDOitf9OqUX
`protect END_PROTECTED
