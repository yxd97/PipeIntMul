`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFqngzTRqBctrzz2pnS6qaYX81omghWfH6t6iO3SXxb7YI+Y6w9dlwjODvT1lBz/
8dlzXBawwBzmj9l6uMKpk5ODK5wblnkoqEEQPH60scGJmqLxJUhBCTI0WOUu+nHE
zw2JL/Go4n8sSCqv4AT1BfMD2wuzg9M4xUlraMfpwqkqPFMy4jS0V9+JMqHommSo
vGNHVRp1L0o75Sz0Fn1uJA0/80m72M9SJ8nBZeMq78Igt/HIAXrG0UcBfxF1ZNp7
tH2HUsGj/lwJAKJ4nNXhy2A5jiGf22iK4zyAxI7S8FLDS7joO6gsEpwNapJHnunP
w+n/xffePLhnC64TirxX35H7LtM9eze7Rff0DQCnqKX2trXWavGDKL6pCChhOxaF
yS1viGGYwv2wEeQRwcRLGhH0BeBFVjF7k5Qz+KX2N5By8KA3Q68QHf/1Hp+bX/XY
5DxHgVEy4sG3wXGRZ5VSUJknODLKejmVWYzkzmdsyzq6fvYS6IqT7yR+HqhBVaSw
ZdDJtxSNlVtK74KqMTkEeXasZIabl5ap5ZxuCuwKsA5RVvgMESS+8qzR883GsB+O
dZ1v/W3xFtO5+2NhrsApid7pnK7fls7rkveWpYZfg7gwYc+FxSakBsX+E7+6uHta
M1yl86ZHbZuqu2EGdOGgZYJE4NqqENno6xmEb6GspeGl+c8S7Y5aF/TpESU0Omu/
wuk74dv341DXsdI1APkR8hlJXiSXzwvLQZgfEbctIIPjH1n3TTVSCsOBLTWxVeL0
k8Zk4QT3W/0cGY3ByD3Q5/shKqNcNS2/dcKi23SwcagDpYK7a14c401DY0lcH7To
OBA5i/I8QJwQgQWzfPfshzDpqNDRmJmntiXsWDOl5G/hsTnZTWknwFhWwV3zIli7
zn/xJnL0OEI3nXsF69ms1FPMs7gRlz+Df8dnzpr7oniYJioctNF5jDTnZDlljlAP
kf4whuTZIYpdQzJH8YNEwpMlnsdEgm3Yhr25HNwmOSItlRcN6eDnuUGfltJ+y6Q7
IqBehvVYe9l7xZ3jmFmJQWqkVGUXVZlvaIFTxxGjD2VqFllzOX2o5xg9+tVKXivY
cLxppnjXmDbEOHRWB9tEmCFiw8GLdMtMPoIHY300V2o1Z9oD4rejgDrViG4/Q+qG
s+JT8ACZnn0gDVPCyiwy5TVoUfS8Qeahd264DFC7poRpHOXy9QFNhAfWxr+Qc8Vy
bbuPPyJnCkZ7vRuWVDrRuKp9Vf/0GAHlsKkxXY4slUCHTJv0RJwtzp2GJkSMKd9U
Cgm7GzLAE/+/khBg6sbeB+ECqBeRYw6k+z80oP/XOZdLcFqrw29wAfqDhUajqW10
7SbFJYV+ydnkpHpuWzEGZ094Ad5+a+/wLLVGnNKvSDZoeg2R7hugO+l1E+v9QLFp
gKAnckXvZzKJjBchfX8RvpYS5c4pUynagu9mrb1awVsbve8AT88EmpGp4unW6uVA
5VZ8PZwRSdgOiA5OEHC9grWWv+6AvMAvTZMUwk/buEf/lR7jv/5r/WWuueq82c4/
AhN4a61WMjRfsyhnVOBryF78Ct2WIR683SjxC+ygscG3DV1KGuewBj77u8UUE0tD
+x0jrMkaWWuldUmZ0v4yHwg7+/tIbBIYrqBZtUrO/XdFFGRY73THZxHb7jtbwzdo
/JZ/erseKdjfXnfBEm1FKRMzLRyEtO9UOG2WVz81gqulwMkjue2jGdv6ZUFGFFYi
TIFNPv3xlLkIqUWfdB/HI7WBcINpkCbSRhQWqU2h881v/IF2NKetCS8lYG2XrhUx
WGkLbQbz1nXDlQFCAknHMlBRKrC89B7OBBoE8lvHiwk1lIJBWX7nGyJffOzI5C3l
DtrW2jKuuldRS73VEfz7M+Fn+EO+dQLvvug0s1Z+3G+VKQnx8OmNRl5cmHktdFSc
k+jYMOUBxREjhEMgRi4bpzXaYkkABKnf7D035CgNps2TjSv8ql5CbDYCh+/0/57n
qqsdqqH08vLZqvF5U2/N9RW/l2ZlMPvD6TybJVY8oZtR4jJCLSWWqZmBIL1x6m3o
vXaFErw1qUG0BP6uIocsf4rEiiGcBEjAwA3t4dNx0Tk2GqRObnjfCU3yQHM6BIaI
1g2PZ8kueUl7mK9e535ZXgmnLGaOAHPwHLIMmhQOIv6ozZPcmx+QPhj2c1Lu94CL
oqDkjhWbuYDNTj9eTN9K5pCavzgSgFNgOw0wGzfrCu+l7CzBPedq/uZ2Alm1x3RD
gGtqinEW1LBCt3gK6GwmsB8WG9whfXiG/ftUcrJ0w/o2Xa8AXF3FYelkzqBbc/Vk
Eqh4hB7JaVaa0Hm2LbINWdl/oXrhz9HTM2PuaJfIrbl4pLl5Y8NRwJWEocWvJ/Wj
rFRsrUP57mxVaxnJHVWg21uMUZ5QDIOtjmwsIwgtxBIdjoMK3GYHkrDqXB0eOJdq
fUXv8uw42RlMLwljgJyJ5HeqVI+psD9NRan2gX4Uk9xtcckpBCkCNSLnvk+z+XvW
/erugRx8dG4tWY3DLvh3cHQg0QYn5su/0arRN+0gTh7c9zLyEGdi8u5sTBYofxkU
jlAhPgnRoktZbvhuSxaaDg0cRp3GAQ/Q4l3LaWnVM5cZ2H5uC8w0tg9TIHVp6xGx
2f1TZaM44ZAyWhEF7eQAgWY+bOCCwa0C9lbnXfkzmOxQezNwPIZvSXs1OuA/5MRN
cCHxNQ5j4NLDhqjsy3LQ3EiqGrbjyMzD65rUZE6uI8q+x8uQv+dWk3o6I31AJ70a
tgbbe44EpkfMMbEmuTB+HAspfMggJxmEfvCWEjaJJAVbWXYV8TeacOVzLwIFJew/
1lN+TOF8i/oMHODRAeh29q4za6RQGS1zyveVatUK5VdD8EX8SdQbuzIVK3H0ZNFZ
5JHzSKn0mABLjQEUBQTEEXcgk87R5eTmSt/z6Pb0mU57Q+4wBcy59ErxJfPwYspD
NnHGHPxbkWB9guYDz8bz41j305zHO7c04WUxI5uWMLH2yh2tlLOenPle4DDs+K9g
ACeXFdeFqiaJYYu+N6QeebE5PfOKccrQPsCLjSNmpeUi0lxIiSI01hMHlrJzzoAN
hSWK4JaFcXcFW4ra5l8eAzC0GX9I6BWlkwyoaGgvGVeumbR8qhorCeoWI2O/Jv1Q
6hJpvOrN4EVoWpvmH215VNwQ6Ax9ZfrK0S29+YGG38TmSZk6NdQaoPaOwCycNfOK
DI3LNIPXt8lBhTmHTbBZV6RvCbrNLUQ+GrwwIkiWESu9qyPp5+RKJl1JJd7Fj/EB
e+Yl7i/LKS05MVI3NAPOyqzwpRvSE2l9UOi6vbJ02FkDaNaZwYAUu1h9ICucEmos
hLm4xtDwzvNNBurKJibz56/fE3lUcEp2LmSVizqHVOE8IPnYlDeLj13vyYmpjSiS
HH/bqqc+Tyu5DAdDVsOm5Tuh3sMJX23Rq3UIfxRDcGKKjlKedJWD896NvWCJ5eIN
ZntJcuvq2Rl4VSfFSIlFfryZWFPisk7Gb6QHw5gQQ1BfAtNoutJTGBOR3d9m3cNH
Ni5bROb3z3qqF5sfnFWg+g/GAuQdhdHjsWKDgQoX9r/MgU35b7uBoju9NFK+ojD1
tL+gKyEw4cSV/f92YpkjWBA8ERo2IhrxlPMGj5B56cxIaARdH0Lw9G8t8WuoMvhc
GlWquhCGCDySDhpWKRhLoOAs31n3768G0L4e2Y+pSGHmx0u2Tz7TrlOg8MB8/7QP
tvU/44J8b/KCcLTJ2N1XTizdpu72azvsgmgwxmH6TCjhBtsylFyFAYrU92SqD9ji
y/Lw8qa3t64ruImzV9YKKoPPzAwentpn5a3bACLfVrThmB+fXr3NlWYgBhGyDp1B
0fD2+aRbYI2dC807plPd3A3BftMduqL2k83N1lvoLiXw50iitbOrfEwGZnjRT4Ht
XSaG6NVug+BRWXrpfaM5CA3mLAyHAfaROYCy8bSFxt9qVzeZKooXWBF+cc2BUzg9
xOOzlRH9ijqXKaunXuS7hY/BEm8YNaYyLNFOevXMHnG/+nfz/uP0ZYT2Pa1Sf2nK
uj9D7ZqUVen2+JE11rPN5T9QGkEDfOXhc0VtneRi/mCaLzuNOm9OLCpJBGwUB9aV
t6U4wIaKQngUswq8K/5mMUDr8v1Y7c+LQ8fPakVwDU7NjmG5lYqdDi4qFtvBUX0Y
Jh1VSoTM4uYVA/RrUKnozx69qlzDKpVlYuCvoZIizD2/CX1UZTV2UqJaTQRDQZQI
bwBRx2TCP6R7hN9RsQ9uc4M4469bBHVDHak54Xfm4AqHphzonxfFgTeDWamUu3A8
C30AWSod0jnESnIy1u+NmPFIREMg+5aymTS19GleTGuRuwcvc6C8MW2YGRMbCW3F
HMis4tF/UfcEjtwZAymfUYFAiCtzSI/pZgFgw9P4CDjFvdjpBm2LaAAqtgSfvSWa
MTZgwAZojFhx9fM2PcZCXKVpv98acFhWEUJAUlBLJ0hc63Chdzl0xxG3Ffji38Zl
CkSaw9L09DI52hz2usVhcgCdTNCNNh0Z+2DO1bMD3P27mxNC8r5VSWPo35T82PBW
giv46C4JIgqS/H9AFp47t+e+bN+P6G2l7xrJZiIkD+bBiKd9VG3eCdR21Gu7Bpzf
ZQBTPAsf9RASJJtIotxrcCHLIJk1OnXT0qoECsvVW1vu4yMe+44qcuT5sIMXqzIf
RGNWdm/rLKM5vZoGBl3Q1ysQx0DOpiQBHvHorFSNAjN0J5EuPB6D1tXSzMhKKH6o
ABhuXX+UKq8D1R/R3ZUf7UfjnNAQ7t/GjXAeRWFempytoHAiCXBO10CBk1+V3UB2
zovxiV+riunvC0rGyod+cuSp37XPMQtb/Wq9aPW8Ovz2YpdFSFqhKPxsnd3Xq7El
e9bw+e89/RE+7+gfHiYs10QFp/Oz/5f/rbTxKJ7RE0TRTXImvuXFrQrWurmVJu/W
VhHBlp/WD4iFCFquLoX5F5MtNX/BIVRYbqojkoPBX6Vtp8/uD6t3GeDuF8mNh9YI
uHfS5mRG0l/M8w0LR1dS+1duyb6A/qtKm5+bizN+1f0mrA53gcc5I63PMhtjUrLd
aH6/c68/zgiQCZsWf689tYHJ+6L/na66tbKaYNTG7tN0HSp806LymH8RQzR8r4eb
1u9hCLd56kiiZasG0Rvo6VBrjJFkJk3otgqqthMx75V1G11cO/FkzsN2bFBUkSxB
jwhQKnXxu+8skGxz5C56Q5I8lqNQgfZIK34IkxOFRE+jsA8oRqCrlcvJOxno+vTa
DFwqbdVYKXFSo695kJLhxA==
`protect END_PROTECTED
