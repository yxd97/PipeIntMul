`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gIfrS76rdUtsymupYWQiik9eTstBJc4hFrHQ5pcuLreeDtsV9DLMWanxY1Cuc6Lr
OHqPfYL/5/1gkYo53zjzuc1gZbKfi24Mo1LRYcxxCuRdNF60N5UWz0ogF0rBhNSo
iPLRn6dr+57KKNBA09bbeo5p94YD+VbUtt+ExsQqhzDS56ugAOe2Qa6yDFDGqomw
ZpnsAtDN0rhwO0c+69G1nanhyPCBhv/+M0CObL9+GO8SwbFXSH3nhCXMXPPoy4t1
UFB/M9RvX1Xh9e/H/XVVlYwgoBS0u0sMtlBVjHd7VIlw4FsfSGigDqX2YRbtYqQa
HwqcUKEA+I+Ky4f1KgK0R6YlBHKA3aVpI1tdlg1Nvbw=
`protect END_PROTECTED
