`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPNLz+DuEH85rr28aEvAzKcl3+Q1R1zJbNTs6fSR+sIHzHBbyBdhxk6Sq/zkz8pr
PtTFCKqJBzbkqQ4zc0Fyn1laEA6J59+64L8SM8vRCwEcdqXnRgyySprtMU08n9ov
+rjviKwuBcPMXvpUWn5D+4SjxRT8vGtUqsH3CZltw2C0ekN9ZaEHyT/bY8iXupgc
t9U3n2y3wacx4IoXYPeQ07t+vbW8LzzzVAt9DgrC8Mckv1Onqow282ZzoraHJaRu
Dtcbsw1bTF7cE8WRgMZ4IpxZErMYgfCkSPS0ZT8vQ4uWV0rSp4ErvnY8b+Vn9m/o
NbH7YBe/ULSXF2X8YccsEiuXoIWn4k0Ib0zjD1bNQdPNMLAd4NaPXy0Aeee2MMoK
e4S72S3cDBEa8Y93ukeTsnkLegnx/3Lz7EEjgGpmMYhfPpFUVII8bANztXGodh5N
UY+J1PZh3cwmQ34KSzOggKvP9VVvK+1Dw7etgkynzi/2F+l3iQ+sIlQxrRntED+o
dULIc7ZA2r6K6ibs7pDO5+8oqrr0Cb3W9oE9o/lV8lcf0cV2jyvC+85ODOBSRoKZ
4alYclEP7ns1bFZ37Rh7kjpqgBwbCXWt+tUWD/yzH0S28mo9/toDJW928ufYt3XD
xDTy4ItstEgeRc6zWhi0Vz+jLkOQKWem1NkSq8zLwsc3hpBWyz66IakRPuKdNTrK
VBQVoFpU5T/XfR5h7d4s1j6rTYlkEplqsfkLvh8Yg0ixF4j/KwN5gvptQBLwIxXv
ZhK6NTMM1u93/xCYt92BkufF3g1yt5aivhKTrOcfQAmSNSU5OXOPoECZ6TkAGNyU
F86ukg/Io1b/OzRZ5CxjTK6up+3Y2F7fJQQgOF9VgHTTvF8/w3RaDOSmB2GOGTLE
sDLkM/hbvQgDMB7wfcZfEPJV1b50YdWUDQhRyBwPfbtIqK72SJ8ERTdkAWvrs5Jq
6JjSit+N/STmDWkS0aSOQU6b0tn+5+SUFDacdMzxXBqadeMUqmHuOvEPKcAaqUJC
JNpqL1Lh5YENmI0/dv/QMlSunyDIrpZ+N9NpJIDgTKEcVVeLiDSyeRYoa+GWszLZ
37cDxR2F1aOuDjaCCpn8qvE9eodtUjpwn77AKo1Hm2+s/4CG003W2PYAUwoNM48z
EJrURe96O0CgC/B6Yjbgz+TxlXx2dZcMcu5kXJX4UmJegWvAkxoA9UH+sadWOoFz
b4lj88BQHm91UJspz+gKB6w1fx47H8e7ciyQoyfG+k0w4I6O5fxd/3xAS2WpnT5u
he1/V1dfVkg4LLLyvGHa/SyxTpRALDrbjVmYWmHjNOe7x8AekEAAmFOfnbfYsJ49
xnbmYsV/pDY5/URgmbd0PKcDpXMVFdcOUdNEosxOQJf6MDV8w6y2CpgoZtRqgevS
7hp2Y1WIkagy0t57sUqWKg==
`protect END_PROTECTED
