`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bv50zRdsxXd8UqNC5A45axXYOMzaK5nmblbvdjUi9lCX3nPKs/Dmjm47cd5Nm3sw
PoRvKUKX9ViKPyeM5zd7qIPt8BXkrV3EUse/eh4jrzRCBcEYrjkVI4HHIFLOSJdh
wVLHI/klO38FQTTNRSUSju688MXlbtaDvG/vT+VSBR3vriJ4qbKv3be5QeMhX4My
XZvJhW85Qx7tPBI8pTo7ycKIAf8bbJfnNY17kI8k45Ni8SEvRozEsAYfxVkMdLy+
D+nmzyFsRa1jBzWE+rFwV/WAi7YlC2p6S7SsUjW+2QuGzGZo7JwgOMCgFa7KVdkA
hL+fRzEdf/tXgYytnu2CUbhtXWa3M8vPyxQj37HcOwqq/Sk7zPUEncA0EKQ/NfC7
4y0dQ/4P78v8j4PuJrkhL3O5cbnjEZsUKfFumJoWTdeSCYGWA0djySVhvkevKILJ
v8ubJQ90VT4i1UbxsmExAA==
`protect END_PROTECTED
