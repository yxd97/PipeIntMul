`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EjaCkQks+d2I2jdouwOzXty/iD+Y6pU6rucNxyT160YsUhw2Z6eokDAnmiBRVCZy
CtfqOvFOUog7dmA1vMeQwniq+o/4BMlOfoCI8lPDKQqXFFvxDLBsiBLXE7qt4lM0
N7Pw6NhOVGelLXfaw6+1seZT7kPfYkt8WHZRnzU3XUhgu7AIfmuMsCuyH2xrkH3p
GZpy8/1by8tLWnFstm0gcI/AWaQqiWAM+4+ASUUT4eVDk500m580J+cV6RoYy6+j
zr+n2MhM3Ly6vZb3Jff+oAMZNmMsCuXc0LNGQwsK5SNAeKD4FokawDVHs5HaZ68s
Wms/470aTp1XAex+91FdJcYdaNXRKHpF37iiTv0+sSgNz7xfu00gG7trA17z4Zng
2V9eOsPlzypFFV45uLBVxUzsFYiDCUGKhwh3Vz0V0VVggUWNqhSx9p7gr3HBGzyH
`protect END_PROTECTED
