`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8Yg3sHi7NQNhwb3Mr67Hcts0EPwOB3kLRbQvEdCZilZt/D1yqsvMt/v4CGtyIaz
fWG+7D37JKrfJmrq3ylJQpQD9Ra/wZD4AfUv4Z4lJJfhUyviUZZbg2YwGuJpdbUO
IpvihZtA5BDbuZGtLD7vRUpKwzbRY+s1M5X62z6fuDgo4KmUuVeDbJrYGBE3AW+S
ml9oqsnXod32PtZlp+9VfUS/IepFzW+cTlxHQGm+Nq0ElusHMEcUmVmMSpzZ9EOM
yacv7HaXyAy+8aqK3v1fJW/Z5Gm1kN8k+gVSPzupjWLH50ejgs+MVFda3hxW1XPX
Wq61wANi+4K09PCEDznprZhtpsv51rivYk0zlC3PyG9u0XOHkVCDxBsCrLC1zSsj
B3GOP2P4zUEo1XrNXN6bHUOm2ydmBWQZBwk1pNB55Rvd5uog2CLF7HoVHj2Pvkpk
1UD/yWx1D00eOVEAa9c5XrJHGNMrlsAhyKC4EGCXwsRViGcHLrOdQBHuRWoI1lH1
WoyIsgxCaXDnv37traZwFWQBxQYoMIO0VUaT54hZe/WMkLdfzQvf6HHzRVwBP5IU
s6gQPcBTMMMZPC6WUOo50aoj4b7uIS2faFfgeQl1a6t6EPedLUIpsnTELMbf/VZJ
mwbVKnbd8ZPKQW0hFib5EFQuuyPBaAqO5284X2/3T8SU3t6qmbbZAmlDE1kXI0OB
tjjln6C1MblwiiNwjG+T8yliguFhOqqbHCvpRg1zbMKjOynFQtFzjvCikt4qDy9w
0+jyT6DI39kVtP4C1Cepxg==
`protect END_PROTECTED
