`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6H8jOSRxFVxoL5H0FS0ODNvgUzbFd/1t+I5+BlbiOZYsfIrlVxMVd6KTHdV4UhDg
bHp2FJTtJCxGu0jimN1GjfcP38Lo0UA2FdsDI06gowHqe8RVBp9ypy+6wsR8mMNi
qMRR5zuc1WRXZ45WF57+v1gVLk/I9b4MpGdjwgc0ovJ3KFy7E77bzn1rnGb2nKRu
oKNHKrJP1ypw76A5n+nDKCqaXcUqx2enWs1/IVtJ614Oszj8qLTwg5nwZY06RJHW
F9huKl9bZuWDF4aiGuVyXIPOb2GBmBhKqOJ0Cdmbj4uhaZvaiGBeL43W8/Lov1cJ
OFxoYjy3sS21YrDJcnTs16gQONL173gkeqXCjfUqjDdvjMerJngp+iv5bXmXk67a
VS0POltkFPV0nkY0vNnzFp/wzhtyjn6yMmB8JFEjIekrOhxtgArOjBCuzv6Pir0h
OMCJo36EIMTM7oVcPUnRZkLjYh2jhwurhq8E0wVcdcObWVBRekVm2Xk7aZVVEjC2
sQa4+m6OQrZU1YPrT7LV6elsA3pKNJKcGPq6V+7q4mIg4ZzeIpFdc9Y3fmoQ6n89
jjXdDfMp3nS0PonMDUrLOSaKzuPbqG2MC446I4PTs7Ne0hReVBO+WbI7RyAlSc4b
FvThMRAF3g/J95qC+h85HKxgOQaVV5KGKqpXksd/nR7EmZSKAHa00+zzrvQdJAYZ
Bf/zBDVPE3zFcGybp+jDFmz/Gwe/hedID1RMXSyIuquJ56aSsqAuexr+n2X8OWVN
hvFHuO9fkhfQECaaqNaQ3YVNX5qVUUgVMR+lnYTEhjs=
`protect END_PROTECTED
