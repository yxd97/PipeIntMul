`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AKF1T6zcKSTGrc1Fl9IPVZ/g8GbY0DYauNu6zKbUzlQ9cqPwKsAtQHGLuSboyYbH
bANEVSSgGlamGjudi77HYyXoONXVm3nqC6CeyA+cOv8m9elrHDpyv9mc9Q42oDCW
Ne8xI8IOgxsqPeq1Ulp2Qll5T88xNGKKwQ+PFtj0taiqH8Ysxo1vNSNu6Av97PR4
zuA1jzQyVJFxb1yoEU1gN+Vgxt3kMUFVtfbE75VLKZyy2/OttjjOYAi6Iv8ceeJ7
Q93DwclWZwo9kAAVOdzjTp3ny+KvFFTYH4KBg4fC8d5Wk6LHsN+AUQ6c3MYe+C0E
euMzUoevGO6VN3yCGelaD+3dhObC7rtZNHZWxAcDo8u0KkB11TTGvmoshRRmDSZ6
5o/HEkqqeidm0cDjm/fFd/vEDsu2Ziwa/FbAoHDzbpG1HuqM1wnYEihMD8MmUYCH
MQ8cxJUVAf96PqFkmdtmTbRGmi3zt68ctPT9zw1FsbSyEMtaeWlcCXgttD70N2WK
/crcs6RvHHxVgyxs7pTrqA1H6NavT2e80ijdWuWw6HcjdjuPOnyJEyLPJsXFU+m8
2zT9oW2G7k8NrFUiOBZO0qbLBCiRCDcqtgE709X/DYiz/Ntc1oPymxThTcsZBhla
YcR+dcXTFFPX6HpPNbok8IJingKe5cG87GNondiL0kxlc+sLYyISDSUV4ev9Fg48
yFGOZHpZcvBJbM1ITLHF+Ohn/sI7Wb4RPHKEqmXgo/Te0KBZKRXOUUnNapHgxFo6
LCZE2aLJebHWALlmkc2rGIQ5tafZ1IH0p4xeUf64lSv0pCMxpPE6KNYGcSPXQJ0A
AabxaCi5H3HEmLhl8VhsaUVcMCfAtI4KIM//KFWvAkw/GGUll21azA8vKH26sjdW
RjY1JZ9NFSAimwGtcGeGOvNXqy+2MDNOVHIDPbquDIj3/ngJJVKTjbQADrI2c5gc
ZL+LJhXz40/35nvOKwRt7Wf3aQ3KHeS3hoEC5Mpsb75KIqiHaEItHaDlNDYY4ZkC
qxkByfMFUn5M9/B37FNqVDOzu2qRZqM+pJqO95/L2SZcd7uJwcNt+W8kxie+/fTi
ECxGZXs69yUM0VbWfbLgmOcYBZL0/nsCl191qF9UrvEfdF088iJUlX8HvlYQojdw
n9eO47uF+HgIGv6qhBu4UIoY+kl65EcD0zzKtuXDdg+octyhnY5GuRbgdctB/25s
++NNCZlQoRxe3LbQyzYdYr3mo1692Q9PYCFtHVmGB65LArBRVThcnw+Xa8eMiZtZ
nRRhz5sN0dX+eMoz7IxdsKGdc3RMwogm6p/Iy3VJ4BRYkZ9oLQwGg5Mry51gfZb7
e0aqPbu2i23AcFPCtijA1msD8J5Oco3sWLQPphX9fq/D+kR3baTUWTQ+UMJWbzpi
soyvfSBEX1MZmY3QWzrulL5ftlYcrnUFkiS3iNmZTt+/yIwlLWktgmFr+GYr1iIW
jA8X060IduIewz2Vt+twHeCKlywT9GewEgNvkfDP61fxQJDqToz3UHF0gOmqZWkU
`protect END_PROTECTED
