`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HpNi9A8GkIYRbpAqI3osuWmNBGLQ316yhE0VGSEcjwtl68OxJbPZTfMcABQo5X6
TBOOjLQx23YPL0phHJ5otWfR4ZqwxWr6IXR7wQyT10/YiSNrByUEpMVfi/6177EW
QT65rZnQBsjn9d/lwfbylLAQMeNo1hWNyPvpyeWVx4pB8xKopz45pIx3vQDZ24IT
EFhPklbPUCnKSW2rWSHFtP9F1NBdoxGJdrD4MavafdIyELCFhNZiIJlR4/ab1tDl
zFm36AN4Xl63mgmp0WvwkoP+oyAUJJ/JN/OEHy9RllWLB4pW6mxOeq3UsuQShevB
QWJpNbrc3nBjcnXhns5no4QAvor9GdJ7T+9QsWf7DcZN74eV+yudyeubalszTXJa
gLMfPP3gxtqzcDU01c0kAQwmG2ylXF8HCKc1jXYxYLWVTaRHNu73HmU5nv3BICVX
8rXU2Y5rInkKuXGlrQilnw==
`protect END_PROTECTED
