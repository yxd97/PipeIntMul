`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zI8aniCIC8JHhoWo0X+O3+h46F6LbxPD0cJQs+4u/jXKUAKmAEnZDtS3Y+iq8YnX
nbXV/Rgff9yDRpnLz7T6BmJzo0ipWc2X9GlwQYPcOcLW84MxhWzSC0BQszE2CeKq
/jQ0r7Du0yZQcxiaWrbL2Ree59QluHELDcI+zwd788cz0b1kuNBS2v4GEUWo5M9H
M1ZPR2Asg4NjzZD3/16LKJeF83z8G0didzOP91YN3e0epOExkBukBPP67xDJ9s2Y
DlgJZ6rycDrRDSn/Ka/y/ScHbrwU/JrdiNkaK+MrZlNwIElkc6A0R5HLpsxti4ZD
l3XXas/KIUdJGPHkKGOtixcgDyMGFQnDKCRRvgU+ru1Af6kYLew6AwmqrIKrEyJI
CoEox+dO+EwPCrUwYKGelT8E1wSG+UmJUeivuLNijTSbtxuFhJtJLRRmUlwJFt7G
7FYaUsr6KnVquScH0u2CamI0CMSsrzwz6/cE0SumYDsCEbUsEuhut+ohAzwG75WA
RO4VcMTdhWn7424Dh08/zMyLA6CdfhDzkVJckfZk9NNxYeiiQwxR0ccNzh55qPcC
VFss9t40q1/XMbyEzaEmfEf5GhZ8NalLO/fsQUQ3jNnbJYXk3snmTcA2cxKfMvXn
O4+E6CA4mjQDCHzuMMdKir4+36Fjx1zcAi1OsE5zH8oJu/kshajFYvmdjqskY8Y2
amOwzo5vHiD8GgGxTFd5u9r4e6nKV/skfkJiC4v3hYh8TbuFgbQfYdyToskKFbko
ARt7e5MXkbTSAgO0D0Pemg==
`protect END_PROTECTED
