`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npYTydGHNO1rFQt0wm78VNZ+vdSvEUN0CD59ZRLT8s6yM157hzhNlsojsz1hZ0XY
OcsY6X5uohSiAOxQBtu+1avyo9G6RJTLPSD/H91aGSpjL91o2QJEAmBURYxSQr9r
9UqBrcM4fdupIarGVGaj9cG9+KAjYN90utE412xD5XRa2CUc+m1/byXgXiCY7K/h
CiUIMYVtQTMRxUVIOTP0OuHpDDjLrSPRNZtomoNbhSXSClixwE1XTH9Mu6nvTq+r
cACiElH2TxkxJNNc6EYeE8TcJF3U93tcyYnwdQnznG5EgUx9yRCLSqghNtnXD4bI
ZPdywMx19F6BnJcRkF5jODWzYUE6Nf0ngFKy/nKi3lyIsRsEf0ZpAo5ZKKw2MZ2m
dCKkAy0o6jwtKZIkE8CQf8FFctT2BlL/9boGBpFB8jzB84OcQa7gwk2eT7bTP1U/
WLI2rhPlP/DAOECOAdWMqmC7toaXCtF9jA7Xn2lTjxbwbx6PAr132CnFv6bb9jL5
Shazg8S5UuQGT/oGxh5V3zcPBrhDYnuU/UekhuX4DX5jIxUgKRns0s44B/hHvpWD
kTCKWuSkSkB+ZT7U3m1QxqOQhm2mtld953OchT/aSNZZtAZDn8GEp3pOU7SSjp9M
yiCBMoPcKsouupJZbk8dU7gJh06LoblonbXiYeWIetI=
`protect END_PROTECTED
