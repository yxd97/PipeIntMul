`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypRumRu4bhS9DOf+Z1X/IhlLDEFLyyiI6QzqujKhizUwxiGdENceGIlIFgje4RGl
INdaaNe+fbZJ5DduBNX/g6Qa7xp+229DiY9KhxGHoe+C90X8UMK4FOubDkoWS1Jh
RTqf0ZeGkF6841TzAajzYDe0bj6TZQJ9fFa/9du0B6TFO1LO0wPpzlyj06xryEyD
r+EmC8dKaPMgUOzU8qiCygd1A4mOUbnIomT8gkjJ4jN6bPdX/gxx9uNDeR9AP1Pp
KqmDUtv7hTdDeSO24cDS1GpsCVs31gBejncpVTpd08LbhQc1hkv+Nl68QUxek2Ws
V/2G+OgBCryBX1Z4rD25VFdPnS3j8rk3QoUGbbdPULiDhRhWMBicUPcapTDO6EEC
kP7goKNZjSwAv92nvheU3Nw8Cdtib9TRpDWC+1BIYcB7bC73VuCHwP0WmPysTjV5
jGnUbV7OpDegLf75NmD8WA==
`protect END_PROTECTED
