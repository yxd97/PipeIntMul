`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9mgMqVVuESEaJK5jfI8tZEluCn+vItxzVXLYQM+nzl0h84ezpvvrt15zVqhpO/I
qKAWsj3Ex7i0V6NgweQW/IwmuYFo7+aXLW8BOTGyxI0BNUJlZq4jG4zTgoQGzD6u
4LwF5k+qj/9zYz1cFSvfryjwJAZ6ZFrLpBDvZQCB3Cn0GZfm/Fnvl3QMOkLEAD/V
CHCGK2RWePMTMhn3TJW+H7FQgi4KHBCuFvXXjFuu0yEYKvkxIpKijmN9VcXsuapR
hK+W5AmBeZsENBhtD7vBo2fKMMpv+IbKxGn1JD6/yUYYKaK6pWtYONPrMzKrVVTq
us0Mw3u5OxkbTDEFVygvuED0yq/y8YKyVHj/h8MaonZXX0B8jjAlsNW1pJ0uGp7x
GkcPzyJYEuWSq9BlQHeh9kWIR6Hoizz4GQvDeTgrMg4=
`protect END_PROTECTED
