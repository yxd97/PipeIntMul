`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qq8BkJxcshGWZBm8jYYBw0FS4dRiVkCLHVGbzk29PPncAzYxhTotaVIZF640g3Fq
N8bhNgI+bWEF4OQq59anEMJ/Qe6M1eCbuYoSBg3VOTjppGqo84e9nA5NRkp9g8vN
QLeJHIVQqfFOdkE00F71a9R/jlt7HQz00oByDmnt39ZlgFyS7hY/+cJNTsWGRVHI
B/d8jmVkQU+oJpDSIiG4svFhsTiVZYeBvzuIp3pZp5fMaT6cmcjWk7qjoeGBykpS
JHd/NPeEb3SmeTk0P64+MHy3iBZ3BqWg0X8KjCxVCUI9oJ2UuI/xkt1Ypo/Gxggy
`protect END_PROTECTED
