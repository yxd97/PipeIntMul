`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nZcLGV9Ru3LfexVxi1eckK3/ju0ZcPYdG3ApHGaHKhzoxAvDz6Mvr/RLZzCURMzy
p6NV4v6gsgDGfz9Mm3Eu4dHCqLjX6v+DtOnxyjqxjMMM6MIRAzoB1cBKMilYMJHF
sVC0x7Aedhps2xlmR7uLHn4Zqor+66suf8kmUMF0B/EcE3KT65kmpaLTxLuiRrhZ
5u22jXMV7SMEXa2ShaEFR/PcbHP4v/LCMwDDBTp+OAb+ISL8/DPlXky/DQiyS4j2
Iq5Zz8CnXAjP7jlVsZ3EvmoMuT6/ZwAIlwNZl0jW/uzBQao3J2MTc4zPk50R8Rqd
pF5Uzrc6syOhdY77i9Cvdy+U6Znq+AvQunJQYKbob11rdHZJ9b3YJexDsGyuAdaq
Ydcxf8JzzeinHzBAhDmt/2cZZL+9SFd8gROfPbAMzpxm4vChofY/i7BWjKwL1TrR
nAbx2Q76prcDYlPJgxUVKJoS5ChNz+2GPZEj9JQyq11tfUjKPlrOD/taIptyHvlD
PRubuS/1OVHw+szB6wwq0wi3kf9Jviafa2kM8fWVFyDn6w4pRZfOPDw52UgA2a5/
I9TCkb34TXExZd1jHiBzKfXrdi/rdm2Sf7kOF542xw0ACaJQi25bDvYsG/4hWWe7
QpETQbwr5Yqrr3AFrZNRgHS8KmABDpdvkS3Dyk8lRIaPx822mKXADHl7WQAqpec/
ZFpb+RLTAhiLIo9V0F+Nji8zJN4zKKN6AWgEhOFS//XlD4rCVL6Bm6J98GeKrvme
q0X3fgg4Xsz8MnJ38U0Pnzy6R8ub18iNoNRDXdN9lci3LWtQ/Mgmno+Acaek0+/Q
CY4DvOmMXsVsnWzzoUnGEhIG1CBNso8kY09we+ZghqNYITU8CZcSmDphI+iLNMA8
PL+j68JbpYm0sOP6CuMlSjaSDFYsPtv1lHslkF8IrTE=
`protect END_PROTECTED
