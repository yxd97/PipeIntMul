`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EvfmO7L6dkfjzJ0sTGLI8TBICTUnE7hbtMgT4wPakt0KQ437ZPG6rAbHSPkScIin
5mmUO1KFmE/20G1lh3GIXWg5VcFY96Zq73IU0GlzJA1+aHU13eG7Awvs9wyw5VrY
w/U0/2S0s67UyyxpGy3RTBsfhVI2KSPat1rLbd9yyx80JyM+Qqv4Yq9jyGjyyQU0
239bgw0ifZ7kwmJ7POP+UNNjo2w+CGQ342Z7LjISrk+7B6YnwSe7DFtcvVtuZvJF
jFXZe2MS5wCVOiMrEBr+oXzxfzg71nblWRrW6EnXL0oXzNdN8SJCGdYLxg8mlHn4
E6/QMZB5UJy2yGFyu+JhWmSgiY4tmEkfmGqMdsOA65zgIvabYqvkmO7UIB0eMi6x
ntC9HLcWu9C1jzH0Tz5Qu3QgJeFa9bkAEFvyzyHHhJbrrEcfutJpQl3dWqCCWbF9
/Y+Ygkw+lfXo3aENUo+AvOoZR2lIg0Q++iGHm9m4m/lJjbFu/HuqueqZDY+yK0Ui
ru9VMz7NcXWouqNo0Shgkgh/TOltNr9pDBuCMwIr/YaiVnOqX6RqIajapCozzVzZ
gU6fYy1o/GynpyZU93k+nA==
`protect END_PROTECTED
