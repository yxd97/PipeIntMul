`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZKYzafQan2t8I0kpjcPRK7hP81HxckB6nlEC8v8+kmmmPEzs5ttHzj8sf6EKXBl
f0iqZcY77m9fcv0dnzTrFEJQ7EFF3S3cGOwvbdgaCabRnbmHQvQyosN73xCkIKR3
zJS8W1arJp7sWfxfApsyTfLTjWUkGB553dWM6jUgMQ1ZlQx/x8sSHEmUro49MMDQ
5ENFeNMfOHJftxryArSM2vLje1ddoZxmUL7gqIlkWudDDmIR52RdkjzjhQuOA0gP
RsUAT90TMkQN7LJW/IZSQO41pArjHRcRoQgbXcOdEj8d2Znl8YhXcPdPXCr7EGCP
7GdWK/IPTUYhg4CRFaubYYoZgMN8XF8W8zzfar+cMgCqc+8zsuebTpQ1MygaK59Q
toiUsQDcmvOgYPpEGl7C3m5ZgSnnYhl9kzeUfD+rh1A=
`protect END_PROTECTED
