`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kBpp2KknheQw6/ZgWG2lNEwEA9is/Q82m6XwCviXOeA9YDAwmUoVNpMD6F6MlRsv
0qVF1NxstEjb5hsP6MOFsGRUbA1MGqQnCu1CNIFcKFssPnpf/giYx+vhQ/dHrPbF
g3e4udZWd313HPNI0EoO53hcFy+cbFTZ8tYNgKEATrwS+GdX3tyeWdMJDqYp7Rog
jEFqafcjEYdJwrzcCvG22aj1MY0XLYhsHcOjF3/4WG//8Qk5tUjq7421mFxRkO2O
uUA3ltgoWYy2i8KF8qvU1q7M6nQPFpIKqi3oqqLSKR2DTgq+zRtAPuSKqe5Y7suQ
B/BGFF9FT6vN85uIQ32/v9ce9BgssjvNtPmpyZjGfT5hn7fyA2T7B8pXCLBAyuXI
u9tYJYzBKNqCmz429Y6FU7taTJvvTzidqaODc3Q9aV/wfC1qJfGuCObQSvfh/wU6
K2ndwT6f0UoQnA2KBGXRvU94w7oPgHXEWZYJi4qdLb6QqaqzqdJbywMwYycdPezA
LoZkt8Nr6Zd+cfLqKbHsr2+afooDNE9x6YbKq+xrNJ/9t0zKvu7yDrMBJO7UbsVw
zpG900DvQ50i1QFOzmmtPBXcznhfR8I+Lot2+RjQ3Difw06w/oOt5QKJeDE5odhO
RLGGCKltL+HE5Ksyvs9nRA==
`protect END_PROTECTED
