`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSP6nmFoVUM5qDAqEN9ZpKAzjf+odWL3s12TjrsQKsBKE9BJZHkV43yBjmh7WrR8
zM7tTf/RcOSaj9B9AziXsZb8fbt1955y3ww413GlC1KhgPMsngyX9S8mdaXLYhNR
CZnZD95BANgoSO/SLAvQwnAn63R1Cbx3FgdGjTwm6MbFfgYT4//Q9CXmNXugExzH
HocwFAseugy6aw6AA5rd+dDMp30PWjd4OUdcfsognrk=
`protect END_PROTECTED
