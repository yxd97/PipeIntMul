`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exiprfzhAGtxgqBwNriqDY0bqG8TX+pEiHyouDJxBRVA3//wAG53gFiukTmIic3H
loZbYhoT4jDxmgD/iJITJSEYvxc+veEXGVlE8yiOtQ34FWTbVvfl8/fCSRLhEdM8
nNPHLOU2n1QTxDWcMOO3dkwgd7j7E7cWWOm8JsJjfzJudGItzweFC4O8vaoIlPUe
ONCl7Vk5jkuEwMWcUOf5gioq6RWiW8LJdvaB0O4260TpRN4U3bsp+FxMgmbFrYK8
kJEbk9JpbCH8tbug5u9nmw4lwqirG9dIhJZtL2qgUFuDzN1eBoABVX9Nck+sYmrt
53oneY3NV/aWIsmqHHUKRRfU5LsTy7Du4mWV9epl0Z5S453ximuZHqyrTxkn/2pM
IiCI/chUB3e31B/uvqCVXoW6rhS32rQ6VwR70dpjqN/pQcuZ9B9ngKmvOkiaOWgf
Qci9dPSs+F8JdVxmMH1XLFjG2UJbRLOWV13K5v196RqDMTAMv4a1wQ7ONPmybDBw
RBnbNg/gSCSbFMh//KeE2LxnIE4U4xfOPWtyIDqtf90TG5bLBd9sMGLNwiGnqPmw
`protect END_PROTECTED
