`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncfs5IGJ1QXY8mnCbTlfO7kDGhzfgWMjULyglsq+TvzE+5rQrONIdFjuAETtq+rV
E9cydPnx4Ep/CIUpU6W4VnjBh9AFzz/zEfEi5vzJ2+hedeNiXJ2hz2Rq5Jg8/TjI
aQzpE2XtiNsTnZ4iR5Quea0+LrAko2BRqSDtYS9iYPQyKUOSC4goiXHnE0ruysac
glBmm3XvwI7nD3TCvohVwClMRC8dW5gfOMaTMAw8v98B/2NqZLvcmfC8UvD9tVSt
AP7ojMqrV69zl6j4gQ5xtSV6ubZWLMKQzaGK+eU5nrEmI9yIYCpc2KEtdENPBtr0
ireNuF8ms28JaGWKmE29jCuP02WxiXvPX8ya7xhnhj3BUe6f8wvevzhw6J2qBk1j
+FlqNpxYfGDzPwsBGktO0xH2Q1vUr26bMztCUbY+CoK3J90xLmTWJwimvEYhlUrU
IKd39qSCKiUXL4XRd/v7Jt7c/12YjWfWnGmJ8H/uhi3z4q/vjHB3ZIpqYpgnzSlJ
4vIFD9Q5R1iO3rAQqjbzOyNCrnE/01Sl5i8gP4yR2zzDg70RtKsi4uN8uXAHECjD
DzsO2WQpgtGIuw44bQkhZjYjBy5eO1/Md2o7dUtYYoLNuexxvjgdls5QraMZknQo
JikU5OKXiH3Xbennyn5FfQ==
`protect END_PROTECTED
