`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1kDDH0CLIitcnD32oo8gAyQFB9pe4HNVmaG0S1AxnbMBrpPmiK6IHzgIsSnuBTF
NTYnZ1PKoSevRJDDCYJ+HmVI533Ljj0C85cAMsuh0a0yICLw3dl1cQIxneJ12xtl
B7MPdKDyn0HmrobFtwwQ1xOy7UYK9jiHoPy0S5bAIHIVPIUOf5zPYQf4UJ2OpJBF
R8v0T6xYBC/usRAjLZFhXMUMPjs64T1ByqEUHOscfLEgF8+m2rYpBJbbQX6vFAc1
7YL384kqfCDow6n57VSF1vNg5zwrW0F4sLyl6VfsFDa+REu3qHCRhxUgIAXwaIdq
8kl9LxiRf2Aansv5vRAUQhM1b7xXRmQzzy5w1zjuQS4enRzAO+Key0fB88SObjss
WfoxtU/bBbxMr3jSxbdL0K/T4yZPTAW9L5nOrBCHUtatc6uLmJWEN/aWiprP6HtS
sZ11QjSyl2Jl9jYLQXfTj0qu1yueyXPOn4jWCizJVw5MmvjoqQJgZhjuz+H2/tV/
znMFG4sPPlgdzDYDYfKiA4FbSeNbttcDydobJxVJMXnTFz65QkhjfWQcQtJVag++
ZSjqc/17koJ4/FfSWE1jUVWn9HDne6i2nWp0M2bd8OmCkWNlHLLwHRmtlJxkm85G
`protect END_PROTECTED
