`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9e9hczaKCZ4DiBneHah3Y1P+XJGAm5d1dMeBssy3Y5nUwhVwOx06nX8hnxl/MzZ
0PfyHNWCe06i1eJYjdYRI/Th6wsiyTvwv7VkT6zFK8qsVZ1LB/Oj3GLM7WJlyQpZ
n6AtzTvKG/7ma/JWsiIHNCzC9YyLrENmTvW5Vda8ghH3fPxhujIl5BipjXZiF4dA
2F7eTGkyafxiH3vcd21li+6JIhh4GEwww7uigerUp6nMO00BMLIHdcQWfxtfnWG0
uxoSfgMt4BIPOoNv4HUB4GiexLwSdwh4OcaqaI12N6gqZBZxo1WZfDcYA2p90nKI
RU2GD1o1awKtCaWMbhNrCA==
`protect END_PROTECTED
