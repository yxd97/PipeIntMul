`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AVlQKPDTk4MdkcvSq0o88YNT/8LwVz7nB/+MBVO1KEoK8tL0x9fgbtvVbZ0Ub/nd
9WUpAPZcdLgVkFBci9e9BlnoW9w9RjVCUWaqSkiEQvsdhlFe+RABfnF2HKONcwog
eS1EmHnQUKTj/I7vk677g13VpeotT44t3O4Nm+dQP5Kj0JfbDyQYcsNMo0aHaeGc
/o+ujiTHTN9Hy7hYTHUpI+c+iA+TWu7ZdGfgPIrpNvWBBi36G/RZd7JVzYJ+qRg9
B3gGE6/+3f/1ZiAcZkKdJ7OZuU2o9uodR8SpQl+0I7OCWggsr+tfqGcOGSLScSBP
JfyFefC430sv4aqagvXrxUK3qQLnI7xzkqnKsCBWzVIk4A54jOCZASpG12gkAAbk
/ETy+e3qelJD85Ueb3Dh4Nza/glIi1sB5ALjq0lsXxutip6+/YSbXiUgYAn3f2/p
76ZM177KnzO9fwUT+J5tNQZTRrWqEJw8+uwdbKXJjB6MTnorQ1oqX5GpwzckqzsF
j/mQnUG9dfiRtPLneq02xEY5Lp4s5Yn8wShriZKRDaZBJtXFYpfazncH4y75tra4
73VWt0ISvop3kUb7kU3ZKf+2BHDcCZbYyR0F3wbFQzneJZebs7pcxD8AmfzAY/Ls
Rh0HWOQLu8FZXNXoaXojIbb8uGA+x3xbKqJXIHQGxgmh0CPiyZa4rzUhEdJKq2LX
X3DTv2Do2ulu+OZEDfoPnMR0qOJq8IWv7zWWiuriuzD7JAF3elGZ7fA0xV4u7i7Y
t5tG7QWAvCKXJvpZv2Zn2GcQ2ANCzJpH4ZjxV4S+E582DciTZZJlTQJwttZ+UqkD
jahqO/tId9EPgxkMUGFnKFXCklO8TZQ8bSjPHmdGq5NmwDVQ5tCVVpccARFPMzDs
h9UD3VJVCwfOTF6zZK3FGAosGW+4DKLx13S7ESSt8xQNkyu1qQ9cbfq74i96iC7I
0jI7GQz26uxZKrdA72zLmf1uQ82cZnZSnxBOyvLL8+MSWHvSvYo7dHpycmk2XuIn
r/JrEKxb8KVJ3VqOHMRR8xDFsVF1WjxxilPD/j6NOnAT0pjMmlDG+WpjOMSNPo3I
Q8K47drv3r+jF3jrIJN7P3ZgSJeXna0zTi8Asgim+HcgRrRdrEdiPOE7aFhjs1vR
rceLdvs4Tq8WqrHtCN+Y+hEcOKJjEx43naqYj+xUHu71H/xs/VdOa4afgdQsTb42
SH/i91oYIl9J9rZKLv3L4SghrPq8WEgf8nECsUJipX+li9asotCp3pD4QzNHGTFW
PPQ6b7wG/oVTdwPtlQaJ4kxA8mgDDI91A5cV+uM0wf3Trbajkt9pEzbmu/0KCRIX
ccrabecdbPSngg/cGLXz9+jiB6vQp1bqvW3j7KlA/0ScbjvmZjifUEXbbMcklkCw
K/sMRbTvtjXl7x2VCHmFMNTHoJ0axCR6gKwfLH4QHjjuGC5tLUrVsTbTdOPrrZHU
ZLE/oIFrLb2jKB4zBEBXoxH5Tu5lfUzoLe9zyv6O0GjLdNE5IFBfvwStRm0djSOY
JrC54MNZf8yqb8I784gzHKP6MdAfxgZAZ6iB4qp0ZSpNMZX03SYfaPIeFvtfdi2z
A9O30dufPaC2sljXQ4nIGevDKXNuK6SUQrMy6GBSKH9XHvMWfGXOhJiia/TDeRep
t/jNRH7NmmpS9osiZFrWXGiDj0F43zmDJ68lQzkgcggSQg6xxCCPzYUtstCwUTrT
AyZ5DUVoht4nZwiXJ502oHm4EcfzT8mfJs9E5fob8mD/5XzCze7PDsPtV1FHLSyB
dkoL96JkrKdWh1fzo1mJXDKuG31ARPGD1cJFaTQaEl94P4nnbhpd8yCb6aPHKYSU
phtI0WPkiPr2C4kUMsDPs8hl6joN8FrjYsZ/IbDk6nSP8e9GeHVX7ojVhgR4QlNO
iziebVPyUmL9KgcSeSspFl9E7clETGCxog/o+xBu5zIf6BCXPxDZqapwHBWBzvMq
rSIT0mpeu/mWvlr7EYSR7syNE4JoTbErpbRxWx//Jl8JlbFlp1JAxxZlzVYqplQa
reYmn1JBRDnv8srrl74m4mn7kWx0qnVo8x8qVKVRs3ZLwHWeHjxyPd2kdKOzWfyP
7Yu6+HciPwye+ztFvbE/qu54Birfz1wA9qxZKWl6JGWgHtIWSn/OZudX7pEJ8+fF
jGdL58XDF0/eD9R/JcAnJtJDaDsE7GgH8YeBDi3GOcyVMVwuNlYVSGXULTl0/r1b
k3yQ3IFuxQArnl7UuPtB2CcvZ/O8ntAtSBvMrpOO1vZEKYjnBwFhfaRAQOIQiXI4
0fE/ZKSWVuY4CloR6TqcqAVUDv5LchoHVhBZzgpHvniTxQDNKNxDYaIwbEVce5nM
UIMsARISciQZHg3yVXCJBQgUIidCA3KvTDWYwm48TYsA7ULcGMwkyTYeyDJDIj3r
cApISSBNHCghFLXcRq6sezJ69aezUCVwoCpJL56YT9m7omeaa65h5nZKeinv7slP
`protect END_PROTECTED
