`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yJlnuilgjDkW7enEVAbWN9o6JA4f/sL2gmZ6LelxaeF/BvztZ4uEHRFtE+KnK+Ve
LAsIbWw5vORaQK2HfE3XIdlh48WD74gitSxD2Vv0JjxsNAbSWE21X64F5u04g52S
gqHQ9fD+xQB4SVworzhRCjh6PhyB6c0jJCbpgOD9UrQnDjb5szcqgbKeqWSXS3nN
dOw/TIO3dHwVcrK1TpqdD4NsB5ougIG7SlWhvGZHzttnXqOJuPIERkF6ECV4gBEq
6hyi/7Iz+XZowXGw1SjSg5yVfaHGqOf6C6Q/0MT3ymBEx5jtbpBId59o7P1xnYW9
wS7nDPdaxxGBgPE9D2a+IzUPhiBxHsww8XCzIc76t4HeyFxtadYmKhg31rrQWWuL
bDaiPU42QTw6HlYo5axbztVk8AaHXCuxmq7wKxua20X/abq6K0yACqcPbevHVZyf
rcESnNsq+/FIjIPXIy6U8/+TeAAtu4uQ3TV1BUoCZSvs2FjxXlJgDjiFRHVzSC7Q
SOvkR/aGwvv4zzHGUtM5T1sqxPl5IxVHVZ9/jvv95ZxqCMeewFZnYjY3sAkdLDrQ
XUDeWJ24PgM7Fy/QTvV5GZjDuu270Vd0pC9WUmHhzCH7TAaNs8Fiz+ChvWsS1n/X
TF1CIE1INrZHtIBwu5wgOA==
`protect END_PROTECTED
