`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgXu+rryNh9fjGcJH3cocxiwPSzBDCPgv6ovvlW/nV40NfVw306bMbRJbSbo1e4d
LYo6322OE5dlzJmXNfAEsCNgfYSi1XDOP5Sj+oexeu28edyo+EoZvu75SNJFQ5uN
lqPC66TlVU+6YaO8+Rbe4A42tBs3Vc1t/ll722/SUiBzZtSLWxDS0rAtOySscak7
Z3/jS18JVoElKnNyNS52wrkvM1AHMCWYKiSZ0QCTg+0cGhqZ4yqepqbDikA9VBGE
G5JBVK15aI6WjxBJeKKjdRmO8IhnDTOdxT5OAxfnJGNEscJ5Hi+wU/kW/10q3O+Y
iIi6admmcjKAWqLpfgTgS1FBoZL0DZpAbrHBRZRiejHqzA88exhVu/eEL2i1h44x
bGsz1cUki0aSJqtok5TpVwBmh0VCN0i7Gumw/aIxP2vGjJ+3nYuJQNIz41tzJ5KF
V14Ij9cBswE0l7GsDATLTLhF7BpRvjhgbvUAqZFVC5eFaBcCib8tsQ4/MhAaG/y9
VziTgj+eS0Qp4kmS21o3zX6zYW7Rm5eDEstDBgfz9TN6jHKzSIbBuvnXjv487/6q
dR9dIsYOTfwZlyrIP57EwVs/obd1WIw1VAHLQ+sa+AsKf0ftJGEr57L08sfXG1vb
Q3X68kiDH4lFB01E5ncktVaGil/A6fCE3YEEyeEJcXlq9e73txQfuFkTCpkGs5h6
5xSVJIke2VOzB1xLpS9JUA+UqJOsZG4cpcHz/SrthMXRc1Wb7Ta9QN262P6jpu2P
Qx+Yi9IucpO6xrUb0w6QQxpLkta+yrpF0i+u1c1CS7la2AYkUPHKH+l292jfE0LG
IKMJtgQ39febBg6DxWJYdSoBJ/O2b+xzJKchAb/EzNPZ78s6WEdXaJRzPpEQSAOh
bbxMrODjITlPFPBEnc+sQgZBDhbZwQkKoINc3sgJIXMw8+/QDZNNdzWDIC4jBcdi
EtkFqK3VDhijGgfwPViLKozUlPvt8L/bzCSbZOyMZrNOFxyq4XHzlYnb0TTdJ+ka
`protect END_PROTECTED
