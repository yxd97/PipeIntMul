`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2JYQJG6p3qeMYByV/vasQtIQEz4zwgPMU3LdHnmRY/0TepUvqK8mWJLAWIMuRaE
5AndPFq7UPu1Lmv2gUCRJdNbBEOfHleK/YKEglXBvLgDvaZYIGSg1W8fZ8c0zI3M
RvdC0niWl08LQklQ+EJfdXhN2MlulQf3hfzsgOE/W04ftIDija6PEAomKjQmg4y2
LzwBOi/F0qvi3U+i2CAHpNVSOxhbVsdxufeddwCqD/AyvYCi9f0HlKfdFrtoQNdZ
dfWaPs9/ymRUG7VacMehs8fLbwrpqIf6LAmoGJDZPtpJLQSWYTPwxDDxLPmQWTJI
rSKkHlp2qG7S+GnR5APQWUDXPyjHgrPZgaybHG5xvX4DMS/ktlAF116a/EuTUSEP
keJX39qZSa4XWCRHk92vRG5ByTC+GZdFHLJs98jZmWESDZpJaroSRm0yUaA0Ju6P
qSjTc6OOls9Tp6MGIntCPEgUfWIjugVImIYlxUjW1GIh6v/ehdGccPT3q3s0zmTK
w+BA7WrCiJ8ZVeIbSu53Hp4WvrwxaYhBuyB2JmJPFlN5dsgya2MRfcGhOXoXXVM8
uoCUpweDd9JWLkw4DFs+s1cHb64CRJAPXGdEURIdSomqiEJzImZD4h5UF+Oeyhn0
qVDMbKN64jNaI/yeZAtiBQ/DHes2MBnR1Oq6+5hib+dgTHOjvfsafu+aFy9XP49k
D/nXlqY+V6dDvQEWk6D/H0A3E2dG7CAHiLduBDSLYD3284GAXwlLmGkrPmpdWUY7
euOWd8YkVz+OngQpBLu03jI/WWimrnxavVaYN4ylQyZAJF01cwfK2GtsqkOKkluN
79SjJ61/jL4FHJLX96ETbxC/YudhueqSH06M866HmIDKtHhyzSyBdGpzrYdUatlo
d3EgcPEZk91WS/Cn9j7Di60mzFkJ+PhIZ621SHdjrJzN9ipMgv1SwYpDU1U9r739
forNn4jDSFp7x1o4fMcL75dVYd1jnHGC7lMQ3QvdBQEigmv8GYs9pGQjBwyn1737
Mqjpc8cyz2F1rVIPvkfjImFd+AbLz+jSS+g0d7do/WP9g74+CQSILcoA8Ws92AiF
fhh99nF+KM+c9uDSi83BrpzvCVJ9HqBaswm8z3pQ/sGpcqWjySuvqBMc+Gf7Esml
sASKPDwo9De17hhfe88wahTys6rzAUi3uQ2lr9L4X1nW+DD8BVksgFMOHUpTIg1Y
suqTONUxfReeVwr693Af2TP2jBg4KrTmqzdoQlTw2a36LTBJHeGwM5EvseTAiq3V
OSTyHQoXYX+qcip2ki/HY5FBcs/0SfHTdWn8cliC6UzXVtA4bTzLpbUBDz0pkvSU
u9zzSDjmSnUO2PdbMJTHy1LRYlmLETQ2vInkjTIFwPJ2cdEfWuJb99KSXhez1kll
SehaUtwOhjIYUfGE0Sa7hCB4j0RFpFA9O37if8IsC+sh7+YD/qdZAS1oTAt6h+Fi
T8soWGsxfDnaBVCSINRf56VvFA1iwLapXjQ1gGCqoA4EaMYvRJgxbZm4dp7q4gYj
Nfj2JIitGPXIsawXWMBKPLDrQrkDdYFuX2865pTcJFd22aezm11a2lw6EcgLVI1T
0TRzjtQ5fP2/VxC0Tf29eqZ9OfPzaa4tt5+tDI+H2ZifSEPQgV9UPDXGEmTMSSMN
A7MpetVmK4CsdpEuSWPzkqu9V2mc1uS6ryvS4bQKKy1ebbChOD6OufTvGDIdRkS2
xaDkmu/WAXiRacuq4w7Zye28W+4xuTAB3S05WIQ1QSDIP+Umk8XqK0pfA0wQXKu9
usJIJYFPlrGCy/GLoudnaxv1Hp8aLZmTEl0C+3f1yEM2Mb6LLn2uUFci89nGqQAq
r34Z5b/NsdNJ1zZ+YgcpnjMtvfoDCfnxyJJDX7DoNHO+dsdrkdMJt3vOwpZw8CxL
4g+c9iDJPp2IIsK5Bj3LDlM5K/bH2Frx+P27wXXgPb3Yt+NPBJ7RcuYbjbgwZwzr
l83WOOfJbiolF46nYC7vfKOckT93yWLD4t8R0/MoMEIbBuEX5I/GGvS5IVHRR4hj
55qnj8q7i6DCD7ArG2KMqlRzn5A2IECMjZxEfn1MXwrpUc71m120cbgukVd4s6TF
s5NRpteVOsX6HkUSELHpo0m+9p/kTfiMH0Fty8R9ZrZEPnJPjV3rJn59LpH4Tj81
YkGrc7L+4ywWUz+Xy7cbUYMrjOtmApDreOFynmfiNd0=
`protect END_PROTECTED
