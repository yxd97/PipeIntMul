`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zM5mATtAMkcsvRwH4KsqXCuoyLg+noacuyt1lQxSduiNuaOoZum2ks2b1gn+BLSE
8yybGcO6dqQoNSnHDOxjqrNOnR+8YMckMUUkYZIux/DjGhjw9KoTznIJYeiqMAoA
tkU4ug/QgWvHqq6ZLGNfhRRHMmeIZtWXNr6WnofNamByDTcYLEb+88V5YKdY+ob/
noASxVlTFdI6l053RaU6wjkI5rAF6KzQF4GQAYqejy7HaML0im8VkxHGlyhbtSkk
6NQ4JPBCbVo/kvQt/yPn3rrB80FmDSMMJG9aEQGpoXE8XrCsi4RjEX7AUMhq/rVH
fW0+rcMtSa163WzDjq0IUaRSv7q+UMSXjK5DwfaPw8m23KRwafYmiRFwPPyKuVio
frA9d8sxG9SCS4rV4g8hx9havfOf2DhxJ4tFkOL6lKIK7aB8NsvoJFGc5i66Vn4+
jw0eVLPuKSgNhuWQs3jKtbC0c6uYXn1+vAs91Ahuz6+StANZ8eaSdXEHJjoLGwbD
JCZNrOAJ4B3ic+xyrhcUMiSaXt5RCKEf+ecTPgdWbpt2OIOrznaHvyJ36xf0B3h6
Zy6R6dw4xSBZHPPQUC8tmE79xNWIITDd4nXDhCLMXBYMjkDGKjuKgyImoz9erWa5
/k+h7cZpwxsqrj9JORCQUCfv4yH5UdhUZogprfqwmW1eQ/KIm00CLhVqoGBg5Cw7
Y3P+Uvl7q/JrKUKo6uAM8Y7Yytnre6ASZmV1HmCDV9kshZqvAUcJ2fOJmAw341UO
LSaCWwEEQ9wBw+21jOKalu3f/YQBhlm9e62J9x2xefXmq6WKqaMUNWuLSNK0yqB9
+BeorqSQAOZJ+a65afwRA2YM+mRXRLhFA+S/LUPwELLvDV1Ciq51P/XNOQ0JzeoU
seZW2TUaq0oOefLipU9M09g4YCzo/VpkqmA7e8QR8CsCxkepdz1arfKxV/yn3ONi
LVcIqY752t4SIJKW1Os00Kn5NqEOP9TUNPVmSLHz5+HPqIiIsul+hgoqvKiDVosp
IfV2HjULPv+g00z/fruteKKbyJGfY8GHswM0OxX4MSCdTr+hW/MKiiwOWuq977So
6fj1KcOvaF4Yd2yTPfy1Qapsp2F5swnX6YdyjIjz2s+2UBqoCBCs1hiFi+kSbR5c
SN92zG1h9Lpk6vEKKMadiVf9w1OBifbfWP/bgwu18v5qTi2C7idAuvkmaU+zXYgV
UhVmnF9WlG9gsFZbG03S02mrgCBV0G9dJ/UMBllMURiV2SYNCLAWR9fmVDgE6gWS
XtMat/TVjCo+bFxwFmTsrGU5pstOEN94M5S++1WFICfvME5FULekEOwf7JNSzTl3
RqEONN8BdW2As6U3Oi7w+WApkdndWwSr4R5N1OnVUFS7UpcTxE2pytd8iinRcvDp
BYEtxzP8KFvvg6Pu1z4mRiXHIElHK7o5+KJIzUU0Gm+Hd4TIPIRRcHurNVjx5Jbn
f2oHfWROlyg+h/BaBf4kvasN4HfEoztBPnQ1soVQI8uO9jzxsnIDcR3zOJ6bmT1K
R/apyJ5TFQxHqnQxMS0wMQY6HnnnBIETHRG5PHUeyl4If8TrzJAF/c2Cm8VZ02ss
SR5+YJXEzXcPgPv4yrArpK/OdCD32MGUQ0PjbB+eShRl4irlDETQ41CoC31AfkJt
oFy0szXEvFRk+8HdXFQn0bzfpPLvkGFEAt7EEcBiLQVrXToGastQU1nSTeZLpNNW
p5Qj5UM0IQJnmAjhuNQJ22ymdRkTNDMDnDEokFQfgtTraiLS2S2GAF5UuAnygzBA
V+0PIGibYItRvyQz5kr4JQfGfhoh7xD33ncPN+PN+TgxC7zwVhlvhyEcaX92Qk/i
OGPwqMMufhrAz8jBAUM656WaouR6AfNRNoheOGffsQry4UcxRC7ji5GymsqUf7Mo
iCPVJhkrExpWt1y/OdOLN0d0Q5Jq6+/RkmJYOVXNm0iKMf+q6CQXKMNtiDgtTEiq
rXd5rF+r2bfxV0FFl9tZuCxLoxU10Afty3/XZ+zzOYK5qNFfKl7hVWPiuRaRzGEE
fLpaWlX/wOKAsAmUM+DOxR2cQTUTW1nQjnf4qbaTvbVavH/vnINIbaMZ0tEGLf1P
UmBjBUQB4Nm3tAo0Ih9uunXQ1Ww+C9urjLVVK7IH0qcFRkku7duhrjedQJMov//h
D4iVEmqI8pW7ap4Yy5EAw60tTCzwLlfX9vNL/OZ9w5+Xl+fo/y93Biw9/ao6ytor
ExFmlOrSkCsEk7Q0D3i3YiduhuDxAdzTFr4jl6owWm9cKythtX6sXA6mNEa4a5bJ
ApcKnYUu4OTA8diBgl/ld/LfnOL3K/wY/HMEdqw3HcZRJsrmCHDQBKLg7dvvaOT+
cAe8gi5xO+M6yNFq/CaSzPSzHbBdRToOuX/VbbcNJCH/OyAD5Z5KkNlZuaoqKqL2
Kq/KEBD6EkvznG8aY64qwVybF81RFdmlQpIj5pviDgCF2zJL7G9yXjcVCcwM4b9X
6HgA+E99IOOaFtBC3YFsXLdmhMLoFZsrx571dpsVfiZmITxIXyKYXiiJI53w1Om+
s9rQyMPhmOovdQExws9m6cd7Ol2z9QQqFEhrDEMTY+zMc34gu8Gfzr8sYXAD67Ju
ubYBva26pwJE4U9y8QWAMk7W+7xG2Rzi0MmQOCQGuzIpJkx+0PiC5MEp3J+qv4xD
JJFTnfoCBVKE4ei8epLCjr+lXtCrqpos0m3kSP8BA3wN7n+xOyWa1UDySxxDvbTg
nqTCNDwVdBuIh3pRglSaw/tH5S/iq4IBemRHdK58gnO9kiIEUwBmYr32IS29fTnE
sxS2I096EWEDlZJZkMuv1xbAPWeI3YDJHRv1245j0vjxY3Q/RaYHqJcyyiwmr20c
nCwpr1uMVqYXCjCBnXpWmpfL7baPL422VBa4OpyxGxSuZAIIBmuPxBmkGZ1HbPSN
O3JA5k2dXooepQlqA3Tkq6TvJowgfaUFse1/PojOVkuFf8r9CNWSlHmpFV2ZmmPH
ndw4C97SVRqMfh+xXuxV+d1VGq9w9tDugH/JVmPlXkdnHtzxmdlDVqE9mxzO93X5
bVNfCMg1qcxfZwmYd2NEDgBKKx0EZtGW1nftA0sL06SsrmIYvikB8XeGsWHLJ0FW
2Y8F3JEHQAXN3Qrz/Wp1IitRSRY6FlPw4BKXMY/xqq3eaI5gQz50oBChLiwepVb8
X8Fb9YHv7B/3tJW0Q1PbR4yXCK2StWcHfiHZ7Fblt8GU8BsJVCdH/D/inBREUpi1
eqvzHZeEEdr5cK4BBfyBnVINzW9lHe7ajraL4xScc0Ykmjnxx8wqkU2VC4Yq0FEn
asckJkzsHir/uKNhMZhku6xN0ejsbLf0Ds4DDIIC3LNdstFeb1RXzP101RTDD/ep
dSD72HnMf6LU6m7/ROnFysl/c4QDTzi1DjK8j3d9Jizyb3cZwikKUMsRePBbVkOE
gHq1XoBpW4zaKxK2vYbknCkjnSiYx+Ofq8ewWHxRVz38TK11XqR/tI66e6BTs+qu
2BEGle6H0S0mgRAOSYub5rAjOj2KSlgi832clkai9+jOj2mLilzOJ2gKziP7pDox
H5EiRqimw3ELBczn0H1l49+ar6SRC03r8Hc+tKbJhtFwnBody2gOe8DIGDEM8uvy
wmpkB+VbvLMKd0I+15ma0vq88uYiieWqa5aAxnnoqqxKIQ3Kgcwo/bD6XhqhH3lY
Ca4bqUkkgZa30vDrM3p0IV2Mg/fRe9MbvJ4YI5+M7inDdo32DOjTouHWEyrgnklp
FmwZ/3nF3TrKZEpk54rWbxUwhSQo7t0XF34UCrIy8OFsoWyo7y2wcAQRgjhMMwrD
ewem8FxrV1LLabli7kGDlb+yWBUNrvTwnYkJjvTWkCW5lxYhyquUKrWHm6m4uhbl
Mf8S6iT3/ipwDcG/1imd4rZx9aJlpnjgpzlnBtGz8wW0sMuHzGKYAB2pobf+trHR
6mJ0zaI5R6XEt8IY/+x/LO/rch3rwwwx9h3Y3hZXRiHxef+G3Gm7NH9xqRB5S+u8
MTNTulZzd6SkQDTNFNaFMmgDJwItfAL3lgFQCrSh1mhfqSiKZj8L8V/cjfFLdaFp
gGLdUut4quwFwrXWq9nsgytg8GYCIfqwixQvKpjp++BdtA+PaJHRrX3UjsDGsVez
dJkCYzOgz0NBdcr2olz7I4DsE+cRTDQqwiZWlvlcij0rDTmtfw0XlixBDvBBDsfC
//jF0+A6PCDTi5FAroRp9JJ5sIyoxVQrnxrNL9Kmro1OJhLJI3p9dTQ35Eoo2p81
WsxYq5m+Ady4QcmUvqGbbTn3726TjwHOOAdtEa5Hiz2Uy2IkDdF2IuBvDPswqpyy
XYvCReU0earCH5EX5268Edf8F8mLx08nLkixXzBn2OQmZ6nWgqQqtC0m4ITQtDw2
Q3Dd7pOCxnWYHwfH0oodGV/To/NmrUkY6G3oTDAiUvbVB+kML5RtQTse/J3TVNdA
MHa5RPyI57JoZX7LclQkIo5Yza3bH3N1gx9qeSV8NdRC96SEwmG1GoiprA2fjE2R
j4gmR4XK3SGGGtWOD/pCz7XkiUtqlVSxkUjtmIz0f914FMzzsL2v3zvigu1I9sMH
Z3jrzHt1EzpNBPGMZdzvc0SfFvsxQM+57DrUu5Z/y8GWceu9p4pe6xWjyzka4zmi
yWH027YtZJP4KaYQPt0c09ODahijz4HE2xZ9UAzk5m2KhVqpoMKCi3QvgYnHsHb2
QfJtkHPN0w8ciwNqXQXAvXvkYX/3Yu6Jtopcj5oNHuQS27E8zaUKb3lhaJFLc5nU
8S+z19sT/FtN0lXAIU4mi0gNQvvgxVaIzGfOIpimGENixbC2GudnyTCCHv9SsxZx
Wx8UawZcj6qY/fU7qWvJMlnDe8fb7gFjgqe8CjWTXSOpKprnnNUg/t5LlAeNa5+d
vuiIiaahkijoQ3jSHdd+CSddIQy78NezmuJITev+nPzKZJQsu+bNJO4KQlDkat8p
gofEm7BDj0sM1uUJaSaUufB/8lBijdTn2mf3iBX0yEg+JyX3dOb4l/4RV8OOEZw4
mmQb2Yk1JYOX3M3VWUhAtcxq8QVTh+3U1oB7/CH3K4vVMOkh5Iiu0UiijdqfU45S
V8+T/Xcoo+a8NX9H99yRgfRtNJuOM97CkQhv4E0B/L8OsjzSB8VEaLR0wTd3T5j/
+iKs41bY+PdLjM3bpo4U7YTxrWnfh0Op0PkQIC3AhlXoGanC0aiTlomEzt2T3iag
kr1HunLwklT5ANz0zJwxgyjb/9qI9tdJ0+IDgEbKYKQwB2drP8XPqYdBEzhiViuK
HgX1v6nLsYMrgSORn/8aqisO9e54PXuw/rwDvuzEaoInSS8OrbKYSGunk4ezzTnq
a47ReY/QxLPrvl19PccsueImEpwViEOZlM+MZwQqeRekiKinT+hX4UFKFa8gsx4T
RdZkO2INDh9lwRI9pEhk0xQDqAR/N+OxAeuROSg5MDlXaRu/x5tPJjZLdqmBwuy6
2G8gHJTqQWXb8op6ephUafQnRRdlhpWZ5CY5cFTuk2pWq3UgRxSgvfOP1/aXg9+3
F1ntG0P1RmDVtSrLpC1e0eSyha2FnFY10rxyxocEqsnPXLQH9+4Kol2A2DqAs28y
FV5GpwF37tz/qI5TM0gg/WB6W558wjb/IyyTDTXKhxxHxrx87kQpzmfr9/8shmcz
/WNbrN/aFE+hyE9JKONil9pMds8eXSU5ZcGxhyJcojW/MJX1RUTpbJU2eKUiIB4D
maT6DeW4XQrMVhpzbvf0Ru4WzP8SsAi9tFZO7XikOUn35u5ZUE5yZOBsTJDCVBIE
F+3YtCYNXAN1I1P6JCy3XN61bNQrV33lQcb/54J84bK/bJOXj3XOr4YFDO3ED/2Q
MHtKVwV9YZd1MLKilk5A5dv7uuO4IDub0f4mPVyP3z4uvlNqS9aGiNm+kDqUaFBw
0ZlAz7mY57F33L2ViUO++EQr6L940wNdGH53qu/lcmwsXoe0av4ZeR6evJg6JpWf
o9c4YTsh6r4F1TLrcqgMUDOQZpLyRYwG8SF1/uPmvy7TInkA37yRx67FPqwFYtxx
sy4FmtHPbgmfuHBSBCTwvZfG7uTrJ5RZJZVFFMh0XZS+dbgih3z1d1iDpgiVjVSO
6+jxWblxOKywk+i36OAQBE1wxIggnL/wr0Gbh444K6NBoMbWB9eJJamPHzHDxNW8
jyMNhMIFJBIRACVbNTnd9wIynGduf4P9a9ZwnTjUcRDo3RtwqqNS74dVFU/sh2+5
5baZ7jKI3ox5PIYnirsx2SJ78MaD5LdjfJ2tHWCimFu6LGx+DeqeQS49uuKtClPe
pHpXi1VlBqjlBZmug4howXhA4TMda+QlvsFFSqeXwGb1CxhCqburjXqmncaQsq+p
6kulClgESWdf8eaHyqVnkmev6AghXddjUVJ0jCndzfZkNfgL9bQIVAFpPvsYjk6H
XZ6Mie9FuacUCKy+ekFv/5krql0NkVx+X/KJe27fVO4Pad/RDOX3ILNuqSUguC7V
y8yvR8VCwQ9zjQ5pB7c8BoofsP+azn5qpuNTBdWXNi4Nkw8jgdaTDhGjlLkALCL3
J45fJyD8+pDuhzP0V1/s/Ve2aZDKJ4fRTqiJvagLxtYEQWXEInMuYEDCscyjUqot
MXPi6Lsej+9apg4ISbLrwzGQvGPSi9K6rJ7T3Jt1A+6BtOxtWvV6ow6naRsDJjxa
XDQ/BHzd07Jo98YZF9latzgFbcoV9yLPfY6jFJjycStlQ318ESPc9RiislBsCsW/
TYtc+IhOxh5LchyHpCqbP7xlO7stIPXRPZBQqI4lDXoAbPpGqmKAtJMsFZcFCklv
n8/WDykHb+Nhgl9TfFth+h7qx/j8NDPVa6/fmaK28J+nyxsYC2nnQ/Kmc33gcRq2
Y0vLbNbyht2S1IZLXruLBBYL0cIofWUdgq1fnbTF2IWx2ouIs6iqBmurbZLIYmvZ
jgV20sZVqXcmLfsJw15AjtlVC1tLN/wuHLjwEhykVcetKjgqtnPYy5ixtPLiCS9m
zuu9Q8NpSvsuxyL27uIELf/E9K8xmyTTkuIAOoNGOXb4eouwjtks4fZY3CCKqL71
rkSFwAukpv2QaTSsh8G3xqiXHMVXzwOhJ9rF+WUyskuGYEcMH1F3S00DuRFb9hD9
fX4MSyIyMSB7U2swo7Y5w6Nn1/LBTfmZSnGe5c6/6VT+fHJz5x36riO+UIpEHiQd
AgyJNczhVmOxQMwC3xHiwHg6VhF86DlHBjuM2ANriumjynOcWbwXRkdL9h0KRlFj
XNLhbTehWvWZVbHkX6aqSjmj0UkilAaSEDMx8F/ITXeJCVWmVpqLJlHAjvVa2Tx3
J69KOiJyRQ0zW+o8lcikM653CtSgJYFxrIHTRoln2VYEjr68vKZrA1kndA2dZvNr
p1fA+Hd+hRaNA3z/wkXEEXth2ZCVtiu9VE782MgNdGcBsGTdmI+Yr7Jshy2JVUXF
au0burtN6/NSpVYKqySbAId+PPBgCHb/rUrxAKLp4ho9x6M99hERicezte/c39bp
ayeGqI/pABKkC90PadlKsEqaRX/gjC02byBuK+0u/MsUNZ5BK/DRgeteSggvb0hp
6+DOgxCBgxB3Rt76zzRB3NnzvOUMAbg8nGaMn+uCrctNRSkIl1ezUVFnLJEzmNqX
O5lfpgDv+mJMjag6KF89IMy3clWlnhGh/PTDOsvGha2gZ9Ul+GoCLv6TNne4B9xW
rfMUW9qSWwo0Y/eo0h/7R2lfqrvlp+HgahTd5m2z8ZgBk2n0AFw/ivcwgrzdE4f+
7Gn5K24rVO7xCLrA0fv+tAnpRxUT1hv9oNee4dLmbQudvIZTS2WFILTq9bMFTunz
m+aWQECs23itxHut65EK4rqpWy7zvgskpaWf8viDNid+H/PifNh6IAOS3MffIMbb
tR1KDGEmJAEmth5jU34hkgGqqCFErYTd4aaBkwAMxRQaEnr7TFe6BdMqWPGQs9I8
kyoph58rGoTuxSV8oJjxKSRi91i9XEWNG30aOLBdzL62Qjy0XB4zZUhntBEBMVWE
eAPATvKq19cmlgD+/99uiS98JgL8CEXsB3uEIGzlU2WmSdwQRfxB1hAr3lVigwDj
V1LMItLiQBv4j8w5PahkiywO/4rE9xgiifhyMcwTKVoDHq1exydOSJJwvHd0aab0
RnMnbQKItkTqTd4gZn/A5A1umUSWG1R3m4SX6IGLNzczJhgy8GMra4c9Ncib6U3I
7gz0knBi/tIEOTz0bzjDGXpWcA3R56P+md2G2CEyvOGrZyZT+BaB8YIjhToTO2Bk
NqVwk+HQN3WKtfga/oR6JojUi8YxPIAPf6R/hIZEPyNl/WpCbyv06UfpwHASpGdQ
yW63bcuzYEddeSwyhV7ylZcLO5LcWleQQ6VFWiBoSoACDQR7IEbEJaPMC79TD+6N
xfSGHlzMv1PvGFKM4y086p3U+QE0Ktrn18u020aq3RPm69j5NfKexyXRNUnOg66C
AfKh1DSHHUfxv7bugU7AG6HmpHvFA/mmhrEndRG7q1h5bcaFdjDkyB7K/sDlfi1R
5TCfSJfiJ8PuDJ85H+OKRukY/aU34M0UNapuLC9eRL0oB2PvV64Qt98zOJrVmq46
ZDhN4v+4zXniWU9BhjEGfEg8WuE/cW3NG9bo24dT/ovxoRagNBhUvM+/KwGb54Tt
76MP5J7oeBPCDIxr3Oy9/I+EXHAenzlRZcg4SKtTwaXcWmj/boHcVwST0sJxrbWP
xmEOkD5kMma1JAG2dvzwxogz4IjNab2pOB31YfENrWjYuVwrv3AXb1v04cvjTOd0
FBKcbiE38tYShpyaPtsxMB7waCVBE404XaR+thgocFK8CmZ4xmig4b39WFp9D1Zg
AJZmG/Wd5IDyBW5/NYCTjG3QpJKiEkf/DepfiOUZU9ttXE1DyKnmIho/sDSF668t
J8eHz5DbnwqauLXaQDH4WrM4q0KWFw860i9eGEuI0CnI35lzZqUPlIV7CAVzvHNO
cRlHA6VVEQOYxdFVI2o7nc6YbbuOa/8OrYQdhFznNv0vVRfXcnjlJiOzfkEYFfjr
czKvmeYkKxlDKCDrov9dCHXUuhR5XW3QB8jU+47IMvfSPpdoZmrn5N8v3JZ5jSrR
0JQtWuq4z92drNlShsCX9KMQFcSHwDni7rJSqCedNsYLaFGLHu5JOvQTOZpf+CUl
AOHjoJvNViADRKq2x/BpFB07vmXHkeyowEMpZJqoiUzXNDAt7chXRYuKBtDunm+1
qXseiqpP9XybH4gLt+lXnlzTs+WKcXt1kKletfZiCvXUWG+jrLpw4+BwHBrILpYs
QgJA6JxRTNl2Ds0d0Tix5xUjeeIR4AU/1X+QeSFwnz1w+YYzyFfXn08KTpI1STa9
ukyND//DMiKTiVPJt3H9mWNmDf2bxtj5I9Czykq22yIQGf4CjIjrA3oYSP7VpxMU
aVgaut9JpTkNhGi2iwj9/ZTSQ+aUyqCF9iAIDNU+SP0BxLUfhjT/1vGhyq7KNjBI
BbnZwfnzoHjXvqQqK8B7Nv1dvKFy2plQWpzDNc8QbrMpTo81LSe7VEtXa1jrfjoL
ofpPuvxVVmOUeWARaKVuXNQzl/u2pjWoSYV4nfEllJJgjFWWCjErsQQoHluBdCpm
SlSnT/qZbC18CR0UBByYkibxK9mHAkTX9KAbAuR7MKm9ldqH2rweBbUgeG2W/SeA
YgKQ8Lg5M2BlxT6t9xBKnH2yaUjYZsiIJizsFm6+BK17ynv9sXckJNJTdwVslyC3
epo22wzqptJ5XO+irl0BC40e0XsmTXAiai+6F+M/FvgZy3eckilGZDEnDOXgCxYq
NsvH4E9iweKfzNvXnZDP25Jtmjjz2SXsyStuhtt7KbBNHnYhljsL5rPKXOo+li7k
PF10g2D5AVyH7caXSEoCEOwvpjlrwfnuLP7z91nWAWVs4dtb1Ct45/OCVU4FpyJN
zRKC5JqdrcGTaW6SOC0NMEDtS2ujQryXdkCIl4071a3Fu8OnOP45W0yxiTlH6gZU
0DfjvwoJo7NPhMOmSv6c3/ircPmt7qsnFK/1rlU8wsKbKW/wITfEmwA6L3R6nUmb
WQWDFk87J2fmO+arSEXGV7Z20obWO/S4msQMyI/yjBCCjiTq9aA3jGCxzsMwz0nu
gilWMogOId0cHt/jOoYcHouZz2XcE/EKTIQLVdZIHXJ4J45c9bIIoKYxP5oDP51f
WB5A47Wl01At5UFEteo9qUqETrkQClIKNuGialBlSJeDez8Xont7RkYJW8/fdDRE
Te02bzBtqpn1UboU177etxPNp/5q6E17q56GliqjJaluOcNVP7VigZXFCYjNyfXx
skOXABC4MfiuAzuZmqkXFsD2nwVTeYITc0lIW9aVpV2cVq1gq7ZEn5nr7tl+ih5S
/6okfDy5V2rwtquAgw98PwG00RECR5hD1Ez43a4zDtkIj1BInB3XEj3UvxKWJPr0
FEoPUKkXL1+ARzDIl5PK1tA/iMZ26d/etmqp9xj9mz2sZ6YshgdJ7JbwzDWDimv9
LNa+Lory8y9do42dw2gUaELAvuh9roBNyPlDjajsi6YWZ/GfyQpbvZaKuVJ4D8R4
1wNotpT53l+/NphLdideUS+0OmXYfmv2UP9XzL4JVnyDcfV0a43f/SD3YIttAZ3Z
zMnG1WUaAle+DvnXZT9wb4ilYHStBGrIG0/bDPTts7UW3FnGnQ6ibiPAg2zYv6aW
gUAHSljLEuFgYTfBqZrcHynmWj6PbbG7ZT3zrWsIoOQFF4gD9MDwaDORmZ9BBfbD
jkeHXEVFzBH8m2xhSxApP2HdHOEBlQzByZmvJf15HVpVjbFFKyB5YXny+UnsBSxY
Hh6L250gULHkCKSzZ3xAxvgsk0jvAMJikyyyze9tUGA/97vVDz3Y8yBMMrEwJWIP
fG5LR82+ky/4t27+VfK91PhMu5m+hlmSlQIYwYQj2qxyTSqdk3ZQ+38Ivjam9ypy
UUKSTNPfZs9p8pVy9mbXLyhWXCf8UiBuLPeuKi4QeveYbNdTHeqAXP2w5EymCXbp
OrfrlkWtFhP6yHIljlFY/HusUwXfXHBBhzAArnFkEPyBLh+r9iDB0ZJx2rDLwcjj
Np1IF19MdnlTzOGcdddTXzTyBVkQa0VjdmWgLq7ts2sIXNoXhdkyHaw64blD5G6C
nCI7sIk74pgT6EonYSh5ih/prdW6KtQUIn7UX8XwPsbLPNe9qaQoAg36VhTlyu9u
PZ1ZIJXEqW4wmitaIGGNfVRfcJEdFzI+5GkAXTVlBokpYQGdDwwNudag42zfEZOs
j4DSV3kWoclbs9vT8XeYUNg1OAglWIAAwz0vDrP5FzjdDPAxMDPXduVLTn+aBwLl
hvyAHaf8iH2U/9K4wmv/Me0jmVM4znLvhgWZBMnxxA5ya8Gd4Xaz52jkxLyE9vRt
mbdzdjaAYAium+g2rySWBtjXBPTFvUyqkEGDLJLiS4AvnjLduEZeZOhlehme0XL/
N44EOu7qq8ExBoSBrQ3wn7XzY4sSogmnK5HYT7uCELXnboqYyuobVz2jZJJiyNlk
U3Ai0c6QDeGSUdSdCn4Z55Gn3dDA507wmVCSGC7G34uRQCFtah8DaH7lTUtkUJDT
H+9e1b5pHgJlKa/yN2eqYnCQ4uFafP/4Yv2IefAAmJHg1kOfyM0zpONT5+Tznplf
S+KsZnNlmMowCzkO4W/sZMKKQNLjzScQhHuljecl/ZrUneiUUoms2q9NENecLsXo
FSXYoDJa/4Wml0N+Bq+ur5Kmx8hukcgRtZnZM6rQyuFGom3QfS8iqQmMVeuyrNnJ
perKHAbuPDINfk6hf2a7CFA2yAJDUTVQlnnjFuxmcMCHvWYmw3yfkgQMk90t60ma
X6jJQFSmITKHll4z3F9ALUkGnl2ic+D8p7xnK8y9NmHE8IejfU559BtgA5uEniGW
gWI02iinMEkmiz7rQ/Skb0uk1j71ikzWNK5x2Ss1tW4p/46RqOKBsNmjn53UHE2w
CP2m1/0KZUKmv5PcLvAtkwLZhDkiKDh1JjXBjl/+8GIyqDJhUmW+Xuyzc+mfRQej
a4QjR5QI30CJ3iAVJBZnh9pNHHhT+EA5JdSsIbJRqQafXS8eyW08RV+lluPbTNTp
XPGrB0axaGdtEeMDS2SmdJ5UFuf05NK59b7NFAmO2FUll+F/ZboJ1zUr4qO1oeeq
Q8+uVjLZCyJtaM9XkUEi8yMrZJRGqpq0kt7Vr09jlPEWwPUloMzUXI6yGKPUvACX
8MWWnLDPUqrz6rylppITcIwMGUVko/OLZoeSQTD8QF0OtAEzATxthY/NVr4uq8Zw
/UfuU6FzGz/DZCQMVpQbirR8woicpV6aLKv1xQnd+uWBR0dJmqUKpvucc8RXtXQN
gDKmYRILQ/U393wJ2jlBBaB+iRgfl6WZZmbR+PGhfeumne0gr7kob6y/Pzmx7vwF
hPG3fpgQKWDErkgvgfqMulEo372t9klTeIFKTj3qnlnbZA3EDxBev/JMvDD6S6cH
DndxCE32FbJQDV1DxewULFO6nj5jxdJdo00UO4uC4xOnrF8vY8hse+/0d31MVX8W
5yvoglMqi8GJ0A0vyx4lVDIHaULmurd003xhSVFXUefwAE9aPqThNS7qvFx8xhQZ
`protect END_PROTECTED
