`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLq9KqfJU6O8gqkksekRzxXGnaHbIeVCzlo4fGDvuYdOF1GkaRwMarIkFl2/tod6
LyZfkJ9Z72lwPU/WoFwzprTJXRyK11AHgkWQs37ZIFkjs964zHJaTPo/HSsHPDox
DiBbn5IJ41tZLUY9BVMNhzmdQC2lbjTI6sxyh7pt7EuAfxmcRbZlKNDjrTM/4vDX
736YavPMN7ZgB0I6zGLD1umEfuzGVqjPiINp6WwLMGHmO5Dq2npTtEoQBUZn/clb
TCoFWkx/eO4Uh32tp8PcMy4p/so+R2D32V1RI65whF+BS6IX+4G9VxgTFAbjIq/M
P1fK7I0Wgxpo2+SVqoLNVBppjS2pzGdnHLZftYuIrZx2Dqts1VHWaBGhJYVGh8dS
eN13cDuf6BuoSG+DY5mGafNJksdnIhne/4m7M42b1XJNfj1NMcC1wxqf3zYDS+G3
uoSS+ZXPcaLun1nSedAz1I9kRj7+lA906ChWyZqhs4lXLCbibhGlWmSXn1fE8JMP
VCL9ekojAqszOalM5wTyzYNF4VC1asaSb9lSu98eNuK915aeaNWl9IsEBOzjox9w
4Okg28pZ3nZWWPFd+CGJc4XERNXqpL1jgvZm7qM4KhA=
`protect END_PROTECTED
