`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zyhX/qGJ7A/2HckXawWLDMjqpDr0U5e6jRJrD9+65GTix8eD0rXEAN/uEp2KdlzT
lTyUJjp6S5TaXvfdKx8FOp+hmzwK902qsvSBF3gj1Wez4YB6516pHBHPEMlf7Wzl
zasRxPWtjFT7ZWzRKTrkNxaz1jNnUohDqhfvYy87eOw8utcN4GeOK1hTEhVvh0rv
163mwcXd+d3Hn+TuR/2CTBmb7WYEvkFipZZEWeA0faoX0BWWtEzq3c2DETDcipaF
IFJKJ5SqHmbkymYSUujfzn1ajrLloarYgHwEm1MXyjyb6oHOIIleaLjgcljGGyrV
tzNrAJyaVAJF91y0VKEMQoqp+d22D+zz87i6mlEJ22NiGGMImTK3R0vOGn1RCNhF
`protect END_PROTECTED
