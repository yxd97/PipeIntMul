library verilog;
use verilog.vl_types.all;
entity C_ADDSUB_V5_0 is
    generic(
        C_ADD_MODE      : integer := 0;
        C_AINIT_VAL     : string  := "0";
        C_A_TYPE        : integer := 1;
        C_A_WIDTH       : integer := 16;
        C_BYPASS_ENABLE : integer := 0;
        C_BYPASS_LOW    : integer := 0;
        C_B_CONSTANT    : integer := 0;
        C_B_TYPE        : integer := 1;
        C_B_VALUE       : string  := "0000000000000000";
        C_B_WIDTH       : integer := 16;
        C_ENABLE_RLOCS  : integer := 1;
        C_HAS_ACLR      : integer := 0;
        C_HAS_ADD       : integer := 0;
        C_HAS_AINIT     : integer := 0;
        C_HAS_ASET      : integer := 0;
        C_HAS_A_SIGNED  : integer := 0;
        C_HAS_BYPASS    : integer := 0;
        C_HAS_BYPASS_WITH_CIN: integer := 0;
        C_HAS_B_IN      : integer := 1;
        C_HAS_B_OUT     : integer := 0;
        C_HAS_B_SIGNED  : integer := 0;
        C_HAS_CE        : integer := 0;
        C_HAS_C_IN      : integer := 1;
        C_HAS_C_OUT     : integer := 0;
        C_HAS_OVFL      : integer := 0;
        C_HAS_Q         : integer := 1;
        C_HAS_Q_B_OUT   : integer := 0;
        C_HAS_Q_C_OUT   : integer := 0;
        C_HAS_Q_OVFL    : integer := 0;
        C_HAS_S         : integer := 0;
        C_HAS_SCLR      : integer := 0;
        C_HAS_SINIT     : integer := 0;
        C_HAS_SSET      : integer := 0;
        C_HIGH_BIT      : integer := 15;
        C_LATENCY       : integer := 1;
        C_LOW_BIT       : integer := 0;
        C_OUT_WIDTH     : integer := 16;
        C_PIPE_STAGES   : integer := 1;
        C_SINIT_VAL     : string  := "0";
        C_SYNC_ENABLE   : integer := 0;
        C_SYNC_PRIORITY : integer := 1;
        tmpWidth        : vl_notype;
        output_reg_width: vl_notype
    );
    port(
        A               : in     vl_logic_vector;
        B               : in     vl_logic_vector;
        CLK             : in     vl_logic;
        ADD             : in     vl_logic;
        C_IN            : in     vl_logic;
        B_IN            : in     vl_logic;
        CE              : in     vl_logic;
        BYPASS          : in     vl_logic;
        ACLR            : in     vl_logic;
        ASET            : in     vl_logic;
        AINIT           : in     vl_logic;
        SCLR            : in     vl_logic;
        SSET            : in     vl_logic;
        SINIT           : in     vl_logic;
        A_SIGNED        : in     vl_logic;
        B_SIGNED        : in     vl_logic;
        OVFL            : out    vl_logic;
        C_OUT           : out    vl_logic;
        B_OUT           : out    vl_logic;
        Q_OVFL          : out    vl_logic;
        Q_C_OUT         : out    vl_logic;
        Q_B_OUT         : out    vl_logic;
        S               : out    vl_logic_vector;
        Q               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_ADD_MODE : constant is 1;
    attribute mti_svvh_generic_type of C_AINIT_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_A_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_A_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_BYPASS_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of C_BYPASS_LOW : constant is 1;
    attribute mti_svvh_generic_type of C_B_CONSTANT : constant is 1;
    attribute mti_svvh_generic_type of C_B_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_B_VALUE : constant is 1;
    attribute mti_svvh_generic_type of C_B_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_ENABLE_RLOCS : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ACLR : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ADD : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_AINIT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ASET : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_A_SIGNED : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_BYPASS_WITH_CIN : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_B_IN : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_B_OUT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_B_SIGNED : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_CE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_C_IN : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_C_OUT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_OVFL : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_Q : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_Q_B_OUT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_Q_C_OUT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_Q_OVFL : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_S : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SCLR : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SINIT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SSET : constant is 1;
    attribute mti_svvh_generic_type of C_HIGH_BIT : constant is 1;
    attribute mti_svvh_generic_type of C_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of C_LOW_BIT : constant is 1;
    attribute mti_svvh_generic_type of C_OUT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_PIPE_STAGES : constant is 1;
    attribute mti_svvh_generic_type of C_SINIT_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_SYNC_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of C_SYNC_PRIORITY : constant is 1;
    attribute mti_svvh_generic_type of tmpWidth : constant is 3;
    attribute mti_svvh_generic_type of output_reg_width : constant is 3;
end C_ADDSUB_V5_0;
