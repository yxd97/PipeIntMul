`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fiTjMWQGehiV7QEwr4N3XMhmxFvZIhxv1e5XPeuixosKWx0siJ2wEjNR2rb2Bbxn
qXhK9/tSQF/mTxU6/2yumxfoyEmkm0elQ+w5MCI3pnmY4nr8811Sl2vD4K8+Q2C0
nZrjDpFNpUiEI6l4NLUoX3Y+oI5uweqzUUsXETqbmFGJx+4AZBDfHJO/tMADey1T
3hSr+eMckEUwUzTtYaG5Cd9eAkYABbojsiC3VrXrvG84OtYzUOT2q22QB9eclqy3
8VQQ6s/n1ti7UMjyItfmQI7OfKzuOnUoyyqg3LTwHwBw1TT9fIiELT5DcSwUz68E
Pvf3CFKBgenQx9piAVsQGkuMFKseu7lip6CHqzDORVocNcp5/cyRVvK9ofTp4c43
`protect END_PROTECTED
