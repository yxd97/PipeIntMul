`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FbEXqIzsoP0N6+asbpsPaaZr54nPr2WfbfmUhyhe+K8Ze3iR+ZziEJpqFO9525KF
BQ/X4V5HVyPQPhynpaqY1ZANSkmLezpPQ2Ih3d/l67QzpMNwhwJKMHGBb7W07wy3
CaS6j006GMfx/+vZeAciaBHT40x1CWwiGfTvmf1snRrq2Qdtvp0SrVina/UtfOmF
al9PM/d2bdG6WGHuMvLbRhNaL2NsNDmn7ek2Nwktp4eQrVKL/7bFBTk0oSrkWtGc
Oppkv47E4kNVC0p1F0Pokfq8vbP5ZeZLs2GZCyM4VE83MQpyW/zEAbqkTlPgETRn
pnTrC/YYyB1PLbhK1lAGSoPW9rFnnHr6tcOHIpabhn21snTg2WjWSDnEJtW0HLd8
2O1fDRlDqQOZm+RcH57lwvJccLsizmjHuPIDoB3gsscK3khBPlybhpCO+tRszuNB
toid7tVLfag4uZit4dMCm5hRXdFj2ltowtnhb9/hnL/liwf+gRAL7oHBj+p+UNKV
JtSijcQUxNhSwGzdJnlyyap4s1NGxYS1TBoNohxBw5IDZg5Iakuj5SfW9Riu4582
9qUCd7Wr0BIcD+Y570Kmpv2i6NJSqCKjVGJNZ5V3/OTs1rL3MmML2WrCaAwcv0xJ
1pHbYK9RN7WdvziUHZF2KvPjkMBsFtD/1BTdQdQyDXQGf1tVZscILaJt7lDji7VB
ekVgUF6O7MCerFjnWywNDI9Ma6ObVUyibuByA9+TCna/pQHYxvwY1+dM5kiM9+X5
genNkEZb8ACD8FVQrSOuxZrE5yAteR2ARbWru33s0K+331WT5D0LClWXPNOO88oT
7BjcHWCzxXDq18XSHpbP4AP5wbJ18sTXoSARCnpFS5UxhGMX5GA7U+4EWcSVSwHr
6bcDJBC/BmVtHPHUV026IKXVo1s+qckvf/mc6V9rSPjzm62D52Q/c/vPOxPiFa7I
439SAMoitGkYFSNEI2wuqPtGx5817oedOuuRnu6roImAdOGRuU9vTHyuNCuMckpA
aUWUZhzv4Cdnty3ush69gORmCrGEqJ5CxSNChH5Ll7Ij16HqsIK3wwiXB+2BroGx
cxqhrZJzv/Oh/KlBDoqdrcZDNhWruJWAt21CGoL622uU2DOYRyL9tGkbnZY/xhki
qRA+pD/3G6sy8nlooeiMBjDzvFK2wwTZo3m2ZArdn6+3Dhp8Vb2rN3QbUBC4Lw7A
UU0w0JE/jdRrXTcGSFsmBMn6wM24/spVxmUSTUePbXYSdwzmdI84uSTt+n/ZwCKW
bsl567J9/Xb993Pwthe4O6Y5Zk5u3HWC1sG6jbMClvmHBgToTtcd/87QSaIoM8Zp
x/Kj/+uk+9UszZUxgSkP1w4neJzveVoGuiqj/EgVdcHhw0j/EulvITSquP+eaFZQ
ksyfYuIOlO7hhLs42WjHVQ==
`protect END_PROTECTED
