`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mCzDllZQsXNB60vrIzfGcfNlO5TmuucX0kWQptI8ZgNFrrYC5kBb/a/v5854sKlu
88TAVZl80zu42FCy40a4EXUpAUHmlOJAXs+RCqxDTkny4MICwcgZgGfZRKy7sPnJ
TPGseJyWuVl1y9Pu9bQtv2XzhiARiG3iFhWSgYDtQLJy/W5sivdp5AFr/OVPhAtY
9RVZHwDRCkvdR+jmyW+DHYLAsDvAXZl6jqHH76N4usbHOTBwBeivqIPG+LxD65OU
EZ0aOIoH3JOwfdDhO3ngtrvfjqYp05CHQkOfb7OewAYvJh4lVNuUXMZzpwxBCxO4
WnYF9cW6bHdg8kPklwHE9tclQR16fu22ncXDo5bySCezCeHGdirKZm0uzP4bz+VW
lijFdk7tPCXACouz/Hstn63W6cwTyNb/tKmSuiexP7ZOXIeTIJB3325bIaKpo4vM
`protect END_PROTECTED
