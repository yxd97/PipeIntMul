`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S90P/nJm3Q8qi2aX+nDbuALq5txc1iMKmzIzdzmgT+cuTmqGSDQWIVXdpzqiKnfm
sEIs17pYJrK5BF2AMlZlBZuYFCP/UIppWpFIH+FAGKUzbu4jly5405wOp1MkN/1t
3A4hajgj8dZgCz9mtnMF+db7RhSYS+lWbd7yMyF1CqbhU39zrwgyCQeTBmpI5Jlx
vYFnECingTzYemRrecquo64FDyjjBwwYQEz/mHB9m0bLCLyfxLjs5sTQTWxLQqJb
lEoPI6ZrfFz6vpjBZLNDm07rIhSsxU5Z4X29HlN+AycrfmCwLaGJeOrmgQNF8UKd
Ig8xXfvdTcDxSxOQFobK4PklxnQGZp4yhmFj7QAWIKd0JgR2m1pnxpyoRFVlU6dX
9t3ujUH9M4aofwJer2x9i5IwM6Ga6tEmqFd5p8IUpC0S/UJ/mw3n6h96MmnLuqGk
41AHEhe5m7r/WiLXYvHeZ6H8e4oejnDwUPuVyHM0nkupnqfCbRkeBL7lFau4shXs
HPKHUZh2uDhl17ohsmmyFwY8SQQ+1LothH86gBMLum0=
`protect END_PROTECTED
