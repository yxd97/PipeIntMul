`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGhP+ahqKx0YSAEwlRFn6MIkpijaCDAgLvJkfWdeRxK3QoUjQ/42TQQOE7s3y7z1
LifSmBWRWNmkhUftejVoBmPb/9yzMxFznfNZzdv1uSSPAvHItbicUJD4IUsmJX+Z
YMfvpEUat7tOW0/tikXr3Yq/oeM0/FqzieqyXpPLI0FxCZu/h9boVqoqVkvoWz9p
U2C2wUnCi0KwkMmfW5wR3oQeUjCKvy2FMiH9N79rrMfTB08tXSDh65BwbEIyEuHA
CaXWj1caf/lLqkmfAuRNZgKofks62A5HKAQbYX/bBNglEeIxsrbPsOJOp29ktKM1
cO3+TyZo3bzCfrP9yxyJeInW6QfgEBNrMgn0ndn4jYY=
`protect END_PROTECTED
