`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9DGaeg6kBwV1y9mYD63kMvymM1I3JSxA4woyQbp93pRIe9q5m159HfWKHUfj1/8
i7aNd/ssRzTiuKibHFa+XFD3MQ6v9xd6fE/9cgyAo9mEMfVHGP5FngG6y5ypBHwV
1jHk5Ty/VRwbZhxWs3QSnhzdZ85QWh/XBmJ68LY35WEZmjnYamMiKSNyXUYihVw+
npCApznMK+G9zD18nLfRz2Iy8Q/m/mAI8MLjKfgTc7kle2akADsZVZy58rUA6qzG
80B36OCBWtaCU0Sdg+3Y3XBHDNypk9Fmt5yxqUa9F1z2TaRz4UHVSNqpixcvUw7s
rJS9yIIPT4FlkE3P7Z+mKHMDr3kWUB4nDt0hmLEga5R56NQE5E+9Rxe6/t/EwfVy
g0M4HRVo3i3Rz4qY/shBKugFR6QUqBJG9tqj5KYSw+FLMTS7B6kQvU0Hb5LwTybN
0+XqYKwUStrvKHSJFVWYqNLlrupkNei2AbWvXcUgNqIGBrx4aMS/1JpINOc6m8Wo
vkP0NzUiZifaBhN8QOzqt4EQUOUqzyJ84UM6nK+UIIc=
`protect END_PROTECTED
