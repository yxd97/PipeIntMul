`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bOScZ087yvhiacParLazeBnmEO2osQ63aoQK5F3bJCfnZ72x7r2na6rD/aEIZdE
raWY4Mho9hCnJWc1QDevrtu4cJiKNabFNWcLJS6R9fu5gYjxEBsffsEPHvSky9Wk
q4fdSVTx4ds7oRxzCgBVFaYeJABvQjkv4zgLUJUt9f/zLNsE13jDoy0yFojpH4yz
CsCmAKsxHizyewm0KajMDGDCtN4zg2u3ZW5+vF1bTS6Wj8FLjidKEmW3ly1JFOBR
VxqZSeaQfUXYbaUYEz8tfHnMWqnj5cDF4dUPqvvRLiERO+fpdzNUs5m7l99gngDs
74jc2y+o76q914lvEgRvNdsOpx/tLHv1nQIQu2q/bOP0gXwkQaMfkP/SAwfaQ9h9
+KRJQdENW+Zut6nSguaLgl3ZQtk6MGABr4zb88GQYT9Gm5lpz6E8fyPX2Gy5DKBV
HE4Kz+y3KgEERt73eRX2SSNh/bgm9QwRkxDa5cu7cBmakBaRh/Xt89OcKl4l57o7
oPqRk4IO4t8AAgYbLLfrjFQg1I2QCGvXWLCtoUN288fTBxu9gGmbWdQyRM00WnR4
8LoOJuJWp3cCZJWnT8gvoB6vl/swT6q3z2uiGfTrF5zdx93EfloxUJ73usMp3r+J
C6l45wKmGv7Z9Q2PkZOncN+QKyWaRlsRdxDE+/QlVzxPm39SphtJQmdxShDSSMPX
DHNktW1SKMsELnulIP6yRPhleyjDMzjdfxoeCJgjy6UazQLY9FeryXpV2H6WAncW
hzVTDTiFscuMOwIQqKD2HzM7si7T/KFAJryLwQkwvQi3Kxu2pyumgUJurbT7MvLJ
AZGpiBVF8e09ya/BJ5a6hwClE+G2tySXLjSUEMFUpSpWOalhKa6B1RXQRF7WB58C
Yb8d0bQ35ItqavRXpV1nI36NGziWJ1JQhkgy8zCFCQru5ksHCIAjGf7YulWKbZQE
ifE1OboggKjP8SAVacmVoIsFOCacWUOPLdUWXBcCALMS53Kp1v3GOf8p/PdkPlF8
Vn+tV8NuQPgXzwb74qO8OpepYJTGkfQ6t7Z+FrVUDzp4QfTvxBzj+1Z4E6WjYQAn
Hy77jR8TPlE77fvhE4zG36UB88vs6MrN+ZQ9K9xhZFWE32WV4QGFi2uGQIWwUi1+
8GMgKYBT+B/b5IoKaEAcpF9FsxzWdtUbNZuE2SI3ih5kTVcuxVqpSQD/UWFL4Hvb
nOVBmT55DQhM4yESCCMJuosJ2eHohVU1Y1ZCxj45bh56+BHroIyYWIDoVjuXdHj6
K6gctb0kgbM22X8HFvfGu6P08Vdq3y7zkU7nMZ8Auo67UASHDrxNcoosYqWL8/Qs
Zorv8PeNWLjWJVNIN08sGW4z0XBZA6OMzilf4c42F2DfSwc8r9vSg79YVoIIA0Yc
xtTaJpD8F7f6L0kHa8bl+A74GVBSZ7vN+0UiLri/k9rsQ/AhcMHgX7qyS1yyp0Fz
C5teTgsebXs+QbrVpugHAxvwvSKtDOiBrijRfmuCeoTeTqZjtMDZkf6xK2dH4IQD
KcQ2GvP0EHMTWWk2HP99uWx8DnlInreT4KYcgRAlE+NMWpGekaNSnZxmPEfPoHoW
I/zDDJID3NyxMY69mIi3ghHpmGk/nMYBnTP0yU+8XDrr0yTZG0TUQqsBFv/M4LBJ
7xYttuv0dCpBNXfz3e0nsV8WfLuYW5ijRuvXH9/+WCMZE2JIuNDM6UGChhVXZu4Y
XOikaEOPggaoctknYgmqUyNV6E6fzVx6P7ogf2sogv5wUbKg5ov7vxlQYo4TBz4C
WXpk4ELWrYqc46s24l18+00MsOuqygEExsuNFis/+xZigsdn30NX7emvvd/TGUIH
gZoZ7lVLTKhDr76ek9/QNzbAsXrm6BvBFilW0XiPsx5QiOaMhwo9oKIoT6WpDllu
PFCLMBxPjL7oyk5LN9W6HCFbEj101Ozfhjk1qSkRz56XqLL6O5uNiYdV1WMPYhzX
ZiBEYZ0mUheThwahELPKTY3lXNCwcEx3NqJC4lxCWTVlL/GzJVlJPWgs9i+pfoJ5
B72nEwfwsZ7VrL3fXoFBKdyudTlvbowvd7X0/t9m6ZWSAGYb389W+Jz8XYBzZIQR
PZg8zQrRdVYTBg7i/7kl7Rls0bQoUW5UXiI/lVLbkxyenJbVfZygLtnOAlptD+iL
T0mFjYTfyjNuddfk8mkuHc07W9KXzJZwA0T/NYkk4GcyTfXn8gFjZA9nix9KedDB
w8bzFO0sqsx+PETiUoi0/M+4uejU133TGXSbEDVUU6f9gy6w9PgmY3YqdyTS5vdz
DLY7ptntHpFcw0GS4+wng2mX1wfGQ37O+J/Pg4dvqjdjwP93ws3FVlbre/ECRQhs
nSYTjsYw8kp8DNXAPq7hJc2yUAAv5X/DeUVOgdskQerjzCmDbVutBXXVmf9jiMXo
EnIle01bPQvzwxGPR2i2PU8BMtAjmHnShb5momdTSg/Vn9GFdY7KNjZz6GSWTroN
q+IvHBA+N5odiE+4p+f2knHgdirsBRUfVfHxPifNwHIUu6182o2NZF/m6cuIX29a
hpm34EW/w2zi65jGjVz0Xy4CIcHnrEPlocwo+OAO7Mx0JBVuHwgFQX1wCCs4PUw3
ljcYlLq9YRfqSW6eQBQuuYqPHHeL+7ar58GB9mWYZQzKUPgAfWzMjAFBVR07vldL
vntiOrHBoKozmuHHoAkvPLmBatPSGGDc17eOL1YmI2Xr+8Q7/ERnO3GCRFRUKKOV
3pg1vhMa4fzusi8lwBWzPIcWUdJ0qoBHRfFEi8Biq4ssXmVGUziKHWMDLtNuAUhR
QNl8YubDtsJjcD/eESVjwc1V4EDRwTDX2GCAlzh5SYHylXQzuvCBoG+74fNa4OUv
ImOGzXt6kuI1CBUvFSvAu3J+TnS3bEz1vamq4RGq0ZcLRNK2OTOS3QKWwRBWoght
VV4wn8AdfvLAhzHaZF86fzdbIkQbw8mk+pUOl1/oQYcxKJFAYyas7P/BbiB8IiD4
XPE2a87eQvVrv+fTgRoyVaKPkP4XNfHKGgwPfh1Ut5EH8knApxMHQOhk5cIpP1Ke
PPVyd57VPSwxLt1HjK1pgzeGSCi/xuEXieoAJrAuCRA2RgXy6myPmciCkdtbAwOC
I2jRKEL8V0lK81Im9SyjrJUciLKu9UC+a3ON6M4y/UzsD4H1zlkoT/P60rR9d35q
I7DhBznwZzXcF8NMusML2eO6+6qQL/NXxZFXuodMJ+8M0AXAA5l/8t5yKHSI4utu
37qQb9rFkqZ0FlaWrRkJ9zMrvnC3zxBMKt7mHaAJP3D5B0VpqkhVQ2zH7/ErWbYJ
mvxNNiwvboHSiT1SCFoZ523hGV5WMIz9vftHBMrkTISlCMdi+MMMFw/hk/tB8fqS
cgzItmiOfr2JzGDTmF84QHBNUqx9Yu8EH7WARDuuLAo7z0GIFdjN98DpJ7C/wmNr
XxnkpEwk4ChSexpofDrzCITcUWVIhndU38eQGvvgk8oQZgulws+qrqJ+XU5dCYRe
+XC9jLcqEIdxMrfNYQQKnYQuW4iu51stewrDp/BaGs3QJ7Cq0f1hT1j2jX9Lzp4h
GTgG3/eH51GlL4uBaEpotjSMTJNfN5S5HgpPmULyNbso/Xt2u+K/jf4hkOKuAovo
IAcgMijLII6A/2qDQKmoQgfAjKZ1cL756xGBaCqAbApPIE7gy49pQlaI6Syi1Hr9
gCcrUugKqfjAhsY6e8Bk+vSIZrjeT4LqI3IrPLTkOAzx4tLNaP8XqtoGlayc5lvj
PVEOrxjhqwDnE4Be+/bYhns93xvXjDoE1u5XQfDKYXXJLYolVscUd2z71aC14AhT
ZYjDzT0vKRP9HvMUXPVAvabKcCuTfvL05YRTrFRL1yE=
`protect END_PROTECTED
