`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Scr1qrleQPWvq4aTFLDDfEwAZU55xL39fjoWvWSQDnlt9FIE8KEl4yLOHgyHA911
GF9IBviPMMguKks2iw25Peh2fWFvoga1NIDpF+QnKrGezTFXMuugc1BAZ8Pam8eI
+9LRmPiFnMirLf7PTUgVehvhmUC0En/cX0Uf9eEDuTJi31GskbsOSuAW9fRKPUei
WmwAmqIM3jdSHyzX8TpZ5oQ7JPGFQwAAJidaO7d3Y2VojA3FWrwTJB4EgdwqePnf
W3U7sDLwMZmcKFcoxALBz4YPYHpjLfEHvrFiMRPjL+WQir1+EJ20ERuheI+owW90
nDR3myXcAxSee3664I60Gmga7olqYvtL3vBUDNel+m/opaZ4x5LxIrhfWQL8QZ+M
/PPjKfc7YWQpTxe42JotC799f13bagzPSG4bZpNoM4i83Jez7Fkk6YjTBgsBuF+b
iFlGsLRNyzLUqmovVtTjvj+dLuGO/ak27kY0c3ZZFJlsNE36soPljDGMpww+0JrL
18otfa0Iu6EfQPxBumvFdIqJDlP6Dw7gNmuE5U6zyUTpJa59Ax0I4eG2xLzVrZx9
BCwopWRq2KAuVXTGefeysQV896ve5W+/dVSl/kyHcw1+YtzncnGBuiQQa+8krMxg
F3e6XNarJ1nhNCWkcVmhAW1GSyV9Y957SKe0l0tubyg=
`protect END_PROTECTED
