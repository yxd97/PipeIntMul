`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TMyGylz3DcRzjZmsGumPT3L0oWlvK5fQp8RMWw14DwRN1f4s8Z6K9LU+vMRV/ZD9
mPRGGm2x4LfGf3+rwh2uVcEsinFsNOkdmbR7+igTAb3wnzuO9eIt5AJl46Xik3pA
mgxCz2am/GzcRSZPrVYwUriaIX7yOSG8mJYQM2KkI8RyhcJ/hpg/EGm1QD8dndr2
BX7zgqN5r2uiMpQhoucHFKfk3FpIZrO/2RL3B4rVn2GV6izic3rIBA7XytqCeDei
F02rkG2XdA5Dfx2rTeCYPIw2SNJzN8r/VoPXZO6BNXMZy+w/SVS04/9xFmlw+QLs
yZTY2gh+aGRz8/cKJyeDdx1R0G1vN9npRwBfJE9M610RD+mSFY01/U7hOwvh21uW
YY4RcgEsd7b8zAPUFsPfdrDOj97xU3MvsoQ9zNuCB/WBrCgVUZAOT4yeHLQBcNFC
`protect END_PROTECTED
