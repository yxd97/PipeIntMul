`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYIMWVD5iJL1FOKeeJR8T0ZPR+6gY3jxjCqlcUFnVxsVSLAH/vPrLaeCCSIkpXw+
ZBfiKwn2PX7bghc+c60R6xvr1Wh8hsNOppE5GIhEIm/xoW/uWs55+X1OiFdbkx2l
/4fzszWWo1pGLgdW7KN0OGkRRDQKVMgKJTNQ9abE3sUiyP1nzLouWHN6S8jwkgZe
qNYjhkKUPluQgKuuPsm5cp3yO5VF9VWsZX7AvTAD/uljrxtiuKdmCin/gvpeNSwU
W5dEkT80W+fY5dCRryOnMfUi7epE0zQ4eGo/80sJjDurXb6Fna8UHEnmNZBqZdHt
01lTiTFMo2nqpzOATU2a1KrMCfeXXEFJST7ikvye/7+UzMkz9jzu3jRkATC4gFQC
XZRiw9ApatJW5SVSQhVc+XkOk4bReK9/QfbN9g2HaaV9ixK1ilCgq76w4u6B5Qpy
9/eXqK9U034J2Kt7NKaFHfebUhAWWtZ2SR7IeOvloGUrVNOSY1H1a2faUOpXIUuq
luV73xGKkMpBXw2IJr7JRC3e7pkJUNnR7a6BEDP/FT5Cab1bKdyGQuIg7OK62GsM
zrnadAsoVqzHb9VJLM7tkimSWsSEkSohXVSFcoGQlBqLYrW+dbgw7a9c6aIPzx5/
z1UNDbBkIzPsP8xQil2y3pXNGHjsVsYW7/qbSMJCKVJbMK1M2SEYm3AXJrIMe22U
SprcCZmUuf4kctFwbZbdUTBdgOq5IOa6gHMt9tmL0Y+4S1swX2qRwC38U4jWJfO0
PtW9ABfD09HaAmZGVP97I+65Q4DqUqa71529zymarRg2Chv7c0q7JkxnntgGSprZ
k7reRNjdrOnxrs4tnpbWMoVGLiDuNJoE4uMnp41xNCZ1jq3RdW/rsjVCQDvbpZN7
CDnfCpcCccCNkh1mnGVJET2O8VIx9rowqNWyqoLmWng0zODcLzqc99rqKJ6XbcLO
FgsjLgBZceVMnz3MvmFx79YpB5/vssBBhVUFSuuvQunjusqpIhjWB0p3CtSzIyJu
JfCnkPPh532kHmjYZt30cFr6HwV7SLYYESN+PGRKsarYYNX2mwbgO2hZhhmDhf8b
bgPdEmMpJy4metxsck1Ozd1Aq1DiuifWstVJDOFeAKW1tpxvOsrzz7Le452bjOTW
FxrK9KhBUIw8obrSBic4bb2KgUvzlNAm+0KnnG+siHaAMHjG6Vv6Gei6VZ806K6C
3d8+wwIuKQlCJ8ipQEpIvqXLTDPduNa8b+s9XfrmAK6hWrOBNbVb8qG53pzECSLV
WAM2XbzLaBkEvAi361JAXZbb+iU4ufGi2Ot3t3XmyctDQcJpuOIjXCL81TsgazyF
wgu3COHV/6e/QDk0sHNk02WKu16QSGxX4W6WrNuZ+0Gb56bvqVsLCFQPEQeB2UNY
I4Kal4kuuqXvUbQgjSpzb4hkAWxddGdrrvzikWDo4OnvEOEtnJzld2FkatSZyaii
nNZRX5cX70l0XO+ucF/A68tvtLJsXzYJTb8vyA6g4VYv3vrrOtKBmERjGhsfW+SR
ieT9TYEmsSVncpo3Dbn/gOywB2MNJS+S/c6J8b9RWaU1U3HeDFWLZmsW7mAT+rxF
RL6mFRCZG5tK7zzz4nJFE1q7uQiWNBZk/MVORY1mloYur3UaXElkn2o9aXav7/um
EJS7zabRBckQkt4+xNc5RSS/rQqsuns9PNExVmAtU4Yuumqlx9ewaS6ii4SQ/6p4
rWmHsaB0OLJmK77b5c5V388Q9PBQyI4eaA4fn/9j7dPqFvNXFy9BPubwBSDtzVtX
adPfZPKtgZS0uA+/to3ueSzTFx+0ZFyD2E1GDUmBTHdk0HYACYpO7uYsS6WmcFIU
ucdmaHtNQ7lVdVvD9tv+CNWCrKrjQy0em4nocb5j4LxYI6bHDwk03xaAPr/nl+pC
QJzEXoZbEq3Va5lopQ73DuXOjxMhib/HEhEBLXaPovn9y51jG+LTCqKKCfCuxtnK
sUGYRskvlCm0igiIRPzV1N2rYbgOJP9JRiUEc2NVTZ2GJFsykgXO/zgD3/aLzw1L
za8I74Z/ulyiL4WFmdRo5vhUOy1X+HJPWU74J0CnUF0oJNdwfRBDym102WR4it8P
JNBFfH5+tvLYgzxRsfnQMFw6QQdCK9giaYXxKdoCNx7J85k+0yxezTMLLPZSAzrM
Gbp8dEkSfe2ZPw0ytHRMhdO8apuy6CHYRLmmy/YhYzBYAk07VSgCMlPzSvYznEhV
IZc3n7gtx6GJ87pwg/GMMWyF4dd2ArRmsL2wTNXpuW4QF9m5TSDkPPokO8XZwfmh
A93tG6yQJDSpEFGcTqOf4GE3Hn4bECU37x5o/KCn0D056Y7NtgxNt4RjlISGkX4R
CGXTr7eiL6pX6vw9uxQ7VSOJg87ELicGoDUI9VvlTd2P7Lqx6jkKrbIDM+iok8lG
uRAaRCFnB7TiqYyqBTv+N+b7VckVtVFyOwuQvaEuNZ2BA5eCh/e5zp6L71E7Aih0
BmnUXO/2Geu/w0BNIE4nZ7qtNPtienXXhiiTLMmPMfFWH8xYOPa+aLrcwRtzIz4Z
urj9i+bsfE/TpEf3uKAOYPW9HoFPf8EojlrxdN/rqUpqc6nVnjNgFuvNwkL1nUSC
B+pSXYVoDMPALrvGVTb4KrZXdUdN8GZH7d66Pi85gnV3AKu+Y9BkjZK2Hh19gyrL
0IpQSANx01gt6RXx4HgRA0cUdMJyC26bKHXIlffP+hsydzTSXbfbYqoB81xiyeoK
H1F0dCAHIJ9wRVxywlawfSGlB0FydSuJ08egzfhC1MH0UhwcqdoLaoOINe/9snLc
Dq72VC4fKJC2ZbkdTmBVGTHqwG3q57F6n2ePXroh1sJBIbTwDGVWpN+WjLzwBATw
zT5z1f3hy5wlhuJk7xAMTyyLmgtcFP6BVvNgwZtWiCEZr4Mc+l0WNti2Gg+Pdh4C
3585PiWssUhzqEEJ4Qo8UIwMN3KPkfPOBeWKOh9/w3VqMhaAD54U9AcO5b8heIFf
ezuJYDET+hXkm7AjYD3TUKnVOiHOW/0A6tuBZUpzraZcsljuswCrmVdnQLmY8fPx
5YlEGv7JNcHzpc4wAeRJDvoThRVMMmkgrNlGnFAHn7OkPCFKFdbFQXFqrToVIv5o
EplUWt12sDTTAE5v++gph4FOjOQ+ZfkbkrqE9qdzPXIRo5WP6Ne1On9etB1sKwqc
B9ohXBWeUvPo7Ur27woMtJs6vR3tt0icqYicDglO+/OOXm0+wxGHsy6v6eM6LKhi
6qZD+WD5m0dVSOQV/wrmnQKYjyYsIQS8gaWImFak3zdypBXXqLlnqQMzlAMRhiDi
NTjaMIcJsFj0N0CwW1pjKdaMkzDP1nF9ETsHhQP6/uClj6UoT+ZeMKHUbcCbZM5Y
lvTFY7qbfGGYuF0R+zAvXKTlrqj4eF95rk+Ts7OL5KpYPmJCbLgAHlZVCX1tx7jH
S9DpOcf+e+hhxB+Rb9kHI5BvJ0n5AAsrcw8ATHX6mKDa47a/MozjNUo/sXSPDGon
XK0E1I1kUZWESPZfQW9fisNEnIGBxwgzdxCWiDNKIrSsS1c6zj4lZEoDwxfuJkZA
k6Xk9ZqaOWh6LXkvwb0nTBvky9zopUwwD9d84SljwpXogDfOKJ5Q+7UUc6QUqiI3
2LlzjUUck7tUH2BE7Pi20K7fz1hmxSfnwFVGLLb5jI305d+FBfJQrSBSsqcf6FD2
t4j/R3N/WIGCmj4vcwZIw+ITeqlnnd1bM98Sc2P4yc3ZnKqRUsfDVttziBCVNguU
We8AlsL5Iigp1pBzdSAGDJ0aZ0kCJ71vtq764cHWOt3X/USnWZ/gPWepcv/C6D0X
28H+CoGhXlfgovpgceNgtmo0OBl00iXmRb6XQn+dZj10SOYI0xsiQNbFC9WokZ7h
pgKAXrBlv5K4rg9g6JmnNoYtIIUY6Cl6CsxGLly1DthBHQ3oIYvc0tQHwspbkf/s
g9u0zTS2GLp1n1LqZcNkCEcfFVdcSODReGySKpSmxnSbQ2clkUAIgpED5aT/3cDs
4fXvPfTXV2SvqZQjSJikytNsv/fvhDSl87kYEtBEKTrKL5qZ5ZXatH6Gx3sDJWgU
3B4mvW76BWtWL3uF+dvQxCyJao6YAfL50JVAGRDKg8rdQkbknMuAC06R7V9sHUsa
/HtGwQfZolCaXPdN9P1SvC+QrkIjY6HDf06Usr6w+LNVgLOXH4OAYbCLKUYN7XLu
5odUO4A4LFr0QE875Mb9JcALyGaoROWsqcVS9vYivE22CNaGP7mfTVK/hMw1MnoR
G7QCUwbkEVYs57/hKrmtchAh7jooggZ77AJ6xkJ+6WcX99iPR2KoRNlZfsIBv0+A
HRbn0p72hfF8Ut9EfOA+F/An3dPfjHW1ZccWyxch/iIa1UwyJRz948aS7DuyKU4h
4Q7+E+qyUOJMRSNkSBA8i4+Fd8GWkOwYkIjhu4F7XE6qcIykDbeHMbUYUbhO44G6
Pey981wdsYtlQcfATQlv3StwqR7NFEAzs7Z6Jz+MGymrHm970uXTwxghiWuloj3+
KbeBlklwOurv/rlBOzlerkUfEtPBLQFvNUFlGyfOzH5bWh2t4PNSUCHgJAJFNbRi
RBMAvwCvg8OUP86GZfKi5zFyp7ysGfGzbAwcOARSmeIZdtS/+UBPXmkzO/LToMye
sIoI0cU++tIfeKllztPb8ehCTsYskqEll6d13k8e8FwKkieE5ELLg022hP2bjoKc
GTX3hJFVl9n5m5dt00+fu6FrCBr3vUs2uwQxhTiTGxDCqBWVdZjtSrvHTUuzkusW
87587+ZwKSIOEbCSMwH6QY1iwAacCblgc/kR100MzI64CPgFi59lcYXK/ANlq0HL
5unComDX84z+2BSyeyeREaCuLTwDAE140/YIkuFR/naCmDr4S2yVeQnoYnfukqa7
/CmUbjfY5oY6M4aXlRXf0qze2L/c2f1ye+b/w2jBNPwe1Mv9bvubUw1GPcEL0fP1
ujIoHZAMR0nCTWU6D7Vf/Emx4DCi5NSD/JObDoV1ibMxZRbEqDU/QMLX8vH7YimX
s8hJHqobLKfog+VakWnvQ8BHb2UF9BQ0TbdVmwv+ok/1FSE+yz4H2d0lzmjlRmXU
DNazO4CJsaxlzWGTISz+girxoYjtj7Tl9e6uPMkdhCkl4H/kmFLn1ugysVQym0qA
wIceN0m70xJ9FgyTSnyAhN99hTLfD21gKGpWjKwvGcc1JeCTssZDHw58XUkrWSMK
G3aHMwF+FpqgisLApU1VwzScfnbp1RX5ezDf+QhO+R9yZDQGrqn33PorL+UFIQIZ
zXYLVC2m8iDw4VnJszyt+GoaOU5wC+wMJI+yy1s8Rv4/FlxyBzg8JaP54AePt/f0
ux8ISdX5009ltb8ihtR05czODvl7n7Us8O7Zv0Mdg4VAdUznZ1lC0jfaQrjcEvAm
hx7Pb9mLBAlBm1weqtL79zONoEfcBwk5QO/7eK9fcHLGKo+s1Zrp+sr4zSeaH+vZ
612B4K2QMxPCmLjR3Zlwls+8c9/JwNathG8cPQBgstBTU+jft0ns2WTe4Y4TM7k5
kBZ/5H7zOOY0PXbYZqyQSTvgSrvty+RtfukS33SifD7bi23ga0lhfYHlnbOswmJx
avyUZe32QMfteRSDb6pjhiyegpMhfqBj+0095map2LavJopu6JazyMMtikQmY/wl
cCKW8of7+g5KMl88MlyICkHaXcDBqc1Y2ZWTJFg0iD0NhRS0q52zdANpNTJ+b4/v
3pjz8oj4Jv75KZO1xlViexvF+Zg1ndk2CZ7no8ZeyXycrhKMk7mnWWVOoER63Wxz
9v3uQrF/XOuVDmnxaLbHdgOzv9rPvC3r54TAJ2POM8EzWib6qcodM1OPZM5/DJZQ
3yplcwfFzOTJzkAbFkf54kUEVdIJDt5e+ElFNJ79wXYULrWpiUL2hR85rjN9XO5B
pwVL+u1i4YdNTpioB1D8nU8MeAfv/N1vb9PeXOiqKWJK9nTWjeYUaM9fwIMM35cA
WO34y6FfZ3CQ5ipRVJssCYy3SyIFMtn3fM38WumpsO3xyJcDjp9jRa0iZEZMGie2
qMPqtmkrNlF5hjaw30c5+7/trqYrW8lV3SHyGkIIOJECCopoWQxzT+5F43sDQ1lF
NEJxsemLj1QEIbVFpBWzzEHXB//Zxxl82ETKEqmufs3dIOnx71c1qH4w/xnhKsL/
B9dXK8EYRg9OoR9th/cHBgeeZQ2ENHnn49N/xBM5Xdz6P0GQA6h7w1vX2harnHuJ
lhKIGAe8aARaIu+3fO33WsGnk1BoTneePqw65TJAcU7529wTVwmJ1Z5J/XmAftAL
jVFyIMxpNCils/sMshf/4X8NOaqK831NNd8a8fh6onxXmb9bQBrqRKELWOjv6BAO
9n6Va2t5A795U4B7bHLmJ6ESnMqap/Igp+ILPisPtp03RMqGM5gWx+wyB6etAz0L
hpNf9p96lVSo09+AQZC9+ZsyUo1BRQW7RkOMkwctPwjPGcojwIVtEYwkCWUBVzYv
Hmrk7B1r/3jNwCIBQy1XL//1EEv0tDKZjWojEvj3h9DcZsgaLa4L8gCe/YWI1EyS
9K9MHskpbDu1Br0EkDwoSI7dOeEAwxvV67lW0bBGs6Oo7xuKF9ohOlM7p0F1T0BI
g5Ca6sbOJNUW1sXfB3dgYm10L+oS3VjAoGlgNDeBZXmUhhG2zSkpTTIPOghM58Wh
OAEaKMUqsURcnEHL0SmhLXTcxgk1Uls9qyFAC/oT29MILD5p2Ls44FXX2XoZ+8Cv
0GHfXyyqRgof8MNuP2eypjBufYX1LMPHAlIAQ6ZSGpbQkjMsKDWqaa0og613bVfy
w9a7OAzplLTtlBHgKbbyPeTeaCgfMarYmUyIrS/VflSalJgN90iOidsGBSYHsB6p
QIqQn/a5zoun9g+aAD2spjzJCxZeKZmR1DTtuv7DUyp7wa5mYCGQNmKXZIFdr6gw
Wz38JAgAQuv9WnD1TjgRjE/Q1TXh9UUiWVSmThl8dDb8es9Z8wJK53lJTQJNR1/x
b3YbAtE7JIRzENM2YGFxJYp5/s4k3RW+14gmKBz9uYfZaJ5ASgVhcivwgJhzxRh8
jhSytsQSHmHnsKmxmi7aAbWJrANltCC+hS3GlzgCywbLIKAk9njEXvgzQcBEiGXO
ZW+KX8rl0P1t7/DXQrET+io20H6iK2mlF8ANQ90pgGy0DsCrd3U4xftifZ1l9tcu
aMZVmlCdjQ1lhU/1ra2GG+TbrvLFCctv0ygA7GzJ5xByGN9tsTXPdV08D2FTaDjg
NwHHDSQOnULlHhTj9GSpTEOOQEDsamaCd5lehpFwJjEXKFXjkUjmfa93N5yJjnJh
dYTQZmiJNpOE/eCxOzmK8WyAsoWJBdr5DJk4rmt0mHSh5rVENg78OFLWZ/pB8ceo
81pn2EszU1PnWCnBGPiG/9OcsingvkG74q0hMwL5Nu6zOQBONBdwHuwSbJpgnICQ
gMRnqGaxwADTEmvCbSXloEF0ANUz9tmy2IVbV5ZuqnK9uW/rJpduAmi8q40Xh54Q
nuV2nBO3OzUGT/7FVgAYMyz7qsS3ZC7CwJLKCSgjzibFW6MfX2esityu/tFAcfUI
x/YvKYG+qR757ERLaj77yIgiZJrtpBQsNdoNd4GXms3UdsYY+Cj7NB7BJB3igHS4
djQdiNi4j1qItwwlnNsjRzOOQvqYPuVqiLBTS713sNtbAREcGMNJmHjHgejfPE/m
PNl3vZRz9AeOZqC1iWZFLR2H2cCsKR93ZNkx6wlL4a5AsGzjziOuO4eOnQlrCj/i
1fT6lmwkduHDasarQuqOmsr9fOobNN9wkIBJbxwuJXS1zPKi55cZZ0bXv7fOfdtR
zOJaCkC3pwZRzOojHqPZN2pWfVsqPM+d0ZJbzQgriR2kax8S6YtsouRarITskw5+
cl42D1xKp082pOoMLOoAvh+F7zr6Y9g/Axt16+5FcUAhQU34uzINg8uBc4aEovki
RFu56H8pHwjMONlLGbO2iSbgKj5vJeSj48+C8Rl9eCwTfx/pm77fzY82W6NCBhvl
7a++wFFXi6Pifc4pK+RIUSJbmY/xGReB5k8ZU6C0LaXBYUKHygt15eIQQFNV6pri
f5Qtc6YYP27ictzwZ4cKR3GRZ3UzxBkpwQaYKgLWblZ1hMuOXIAy6Xaylcro+wqZ
pKcOiJmSMYz2pUuHNTfG7OkFkOchHIGEuMMdkq8ILDydq9GDgEgBhVlz3KGN9VW/
wxRgfPE8XsiM0JxEuCFTzo/R4Bw8nlVqKuY2gXcXpXP0h1ogj2dh3baJuNGZOsrw
ovIxUf5aot3yDd8/IRlsdC8btCOTI7FztDBttjXTQKDNOw2BZ3spZ3vjrDWRtQA4
b7TbxWMkbjpm6KSGcXr2Ait1juc4YZfCf4ntHjLSgEMhebpJcCQq1vKjgUH94kJS
pNaQU1P2Sej9iydj48gCjc9My8wEZ36Fy7vs/+rudW6c/27h6UbvcD12VMQDV3Yj
nNg5wahNhbR9ifcaEln2YXFzP9wtMMmMu1OFUM1tkNyCMpZ3szMmwcq/Id1TzS+T
c1aZ68OvscG3nRHMsNlTI19Q+KLckrd+AxYTtXvg7ChrABplMp2ixgGPyxD1zvlP
tDLnVPDqy6DAHwQc98hZN/4zvR2jxZoLGDt8OFCYjmjAhLLPBcYuRtsGPA1iTo8M
fqazA+raDDsyzFnZ8aEFkeNuVcP9CSnGhb1fN0SHphFdd/j7rL6s3yddpFl8ceoO
YA/hXQiWnal+5iDk+YZkL2hur9qaTyI0IIsH4SDvm2e0/Ib3xefLj96t7TAVvnrY
vkhmbgkQNb4Lug36+9DPgeWxJOp1bzt3I7e+Mz9GivmOvtKQYbUwr3DthtRtY7mc
SZ2rbIzb6p2kpV8Z4IO8QV4g4vIcJSNd/6UDHVAywfG0fiMiHZxmK2WMIWJGGJCW
z31K3eP7287iYfrVDqGL7Da3sZ8qrDx2Uf9hMQA0LPUV7r7xZYkdm/10o2fXvs+f
G//R+J6Pw48trnmV7qn9mLbfSez0SMEHoZw/KXprNaw9T2vKSZEZjpUJumomQH9q
OOkEyZt1In595vnrG+JqNIMU2Gp7F7xk3UD3kHCST1TVWX5FgPLkS8++JPErwiwl
xcZki3zC4UfspuxIbtCq8253jjLmOBMWfhyRafznf4QzpqlW1X4yZIsRQz2CzDPO
N1XPcZn6rLGUuIk5VIZAnPAnc0ITn9L9XcWKXNQtjA5RF3kVbE+NRlvBRFzk1IBK
IGpOgqjmjYo5vCtlVNiu7vu3MC/bA/vnlaK6K/86onQQgfw37suWbZsCbkWV6hyM
ZTBB0NFDTCdcYIfxNspDFFPocedn0FVfV8edDKHpVvK7Wcn4vWvcl2ycS0UbSEP9
g3/rS85XjQzsrUjZByFsWcr3iuvy16A0oeOJuznbtEzWPaQkVeZt/hEL8+akveal
ON2tGXDynwmD9XUfTVIe3HMwBWmUOCS4m76f38J7qB7rNPAkwRGmwxemlyN8yHvK
ncVEywnst51MZVaW+KAlCe+Jqei/JzxgRAjzSm5V1tWCd/xYZQ5dvDWpfKcGWF/v
vhG853DPucoQ4PVNvVvx2JvgeFL2sqYnRK2c3JHyH6Ku36zFsLXOMDGlyaZcQzjr
dqDa0q8wXsgLrWLqBMCbiuk7m8KGtlvqA3ZsxIxFctNb6XYf2OKs0f8O9Hn+agIx
htSnSZr5eHPpZOiypEsiIdL3aTKJYCCSXJSrbJEdqMAPGLP63XPJDGokYuP98vkT
qMcZnj3vmWf2XE8cm27la0FYGKBff1FhXEVeZ1ZFImS4Dd1bas5bpuRTd/2mMFDf
9+rVzAijrRZjQcARDMI1i4xG5RLjyDaoYrGv+FQNnJukjefTq2HP8cNhTN3tf3z3
2onAuvNIw/2X2KFPZ3QaoSLBR9V+jp2f0bJP6gHRIKGOA9AoK2zR5yJjS6ujsBxM
PPIU80DaZKZJW3VReG3jtc6vLXW82vedrAVTcJUq9sLv83/Al3Wx6mg2dICWw/8F
9rUt8kuiWa4ESHBTK8bHvfwExxoke7YalK0m7GinW9zYnPHPuuxN6X1Lcjfly7A3
EAoYH7hHUZn5VH0/ehf9MlniO8DZV0QDJFl/TA1R5Fy/4T9uHk8Ephj2XNZ1hjtU
t+u0wpSnDsJ27jHgqnUI6wVzfCHnvRu8n+KN8ZabX6li2z8T4gBVrYX9DjewoaHt
6z8fK6GjYJILzdMZq8iLN72k87k8DnqA4UB+QR+S+8kFd7BPzfxERt2CnuYhW381
n1Yrfo+y+Nibd8BTUVK1ShBwC/Rh3C8Z9luE9RmL5NWw4EQkHddoJmC8wHGoHffF
s6JRkCrl/IRPIyydT3E3yQ==
`protect END_PROTECTED
