`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFiBlRpoxp1HClgRTsepn1U/jRUwjGTqJ2EYrkMINevSJsB93wGV5tWT2NXOgFj1
xHmrvXOmmF4pOPtCEMV26OtXHPQJKAck4wLPZJQhJ0g9LED9pgbJcBdT4rvXOzfK
UjnW4JVHOI4/PuDjdLV4CyoM5YGR26nVNq1LKP6h0O1kr3BQw0XWV+kkBC2F3KRq
L01Are82JBnq6RhiXn6d5VXiRJIHZAMsniC0KaBJBrbZierfgrBxahqj9FrMmR26
fY4e5cIDAO1PCRUoGHaNk4dljRV/EJRW2trO+RPgUpGQF+uaQqsQJsvrONW7/mJe
2B5UUrMSCZXJ78q0fyeKq4OllAirp9uoqtgfU9lVNcLKjtQVKSRhzOJETPTdri7e
2UAbZ3UJ/G4HXGW/Nb+45pedAg1RokeLCFwnW8LEyenFpoR3a54GpI7QvjbEaop1
qk4CdA9ZHdzRUO/hrGcuxpSCHY0AfupzlPXUFTcTJ9ROJuOtLKBmr+VSUrG13myE
`protect END_PROTECTED
