`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxD18gtqVphUG8AnRBfKDLkeK+HWRp0pzEHfdtEysdolJT1YMtZQME3N7Ez7CCuj
0fNzjEFXjr5aU+ShHq0apN2k+9vAF4YmFoebQMOnEW0t5/C9vXvqAoUbsgvIBwkT
P5h6Lsg5z3MWFnfodqkvLeMAsknZxektBgsAt5ac3dtf61k8YH2TWI66gu1q1P9U
f/1iaOb+kl4gkd7TSdVYhnV+HYA7sFTxjX9sSqEAZhfjm3YN6s4LYreN5FmY3lDN
Jbz3IgitmIyR5Z6Ox09HCJddcYXV7Xmyr+hv+RhaoatN7SURs8Re/qTZ4/SjuMiX
UaC40xNkyi3Su6WDHaZKUTjQQ0f9/xbrO3l4BualD0aU6qOsEV8r18/kv14Rx6Dk
reS0sUCsIfzgT1hrOZq4rH5ID7nFhYJmPzbz8gLqbhz4a1TIQ3bwhTptJQtyKHC8
hPMIKtCvSwfnEPsvjmaUSyNWucqv3sLA7JgQ5BrBEmZoFGY0pV0OlABV+GkoraFi
`protect END_PROTECTED
