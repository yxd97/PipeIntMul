`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+27CW+9JUSLAvqgnWyfL6y9roi7E8chAKKCaGiqcokBje9DpNgB7zIyYFMwMAvaL
fhW2cLz0X2Oe9tIJtPqM6mY3lV7WzfGz4v6Hz610a2EibpxegHT4QaNLzROffBHF
s54UPHNeUgp25xh87nspPvreRnbRngaxSSPEznJB9SfU3eo1NxcwG6nWJOFCB3/T
8xDFc2xGWVjZ0EqWeGHYNQ8dWIaCD7hKAi5JH+t8it2nMPWqCBem/niNnr3vuWuF
QKssBm774+M6oqkJyj6JaGI9U0Ik+ZpGLuWVyW+ZgfzJxDP73oii3h42+nFoyqYa
9I5F2VZT0WM74AG1vpLrcNVXMRWmPK9oRvOdvxunqeC5Xf1uPT0TeDfTYL/bwW2p
w1p3hLzo2/aFjnB/VuC7Om5E9jFvF8ZdGHdoQDQRX6ZMbkOmIFTKSMW+U2jPxzzN
abnMITQ8sL3K6yjQxGAaU6L4ermOJ28CG4h+q9EeRq8bwwoh2bbTniK1tuKVd7Ux
lBuJafdr0aVwGP8H22Jvnho0CgZoLHDl1KJUxs1g6ekdpyvExLH6K9GkObsx6IQx
uDJjVvwmPi9pvJDL6bE+0hwOR6n2S3G6wr/FCS/gKIxsE67WfIXXCpKF32euBuQl
Tg9vOceBKr9onsLm/zPCCtwojGylyWHkuiI6WWMWBK+JFKSMam+oSXi9FEVMcTQv
s1GIfoupN7neqGbQaxYDPAYk+LVBfxV4UXhx1rpSX7JXCmklVMq+Or9Xd83mwzwB
TEQ2GLRuFFABiwTxSVIxV/ccQ+qN9coh8XkkfzihJGsmfEARFkTvwBITsy3vLLMk
Oim8zHLyr8JZBKLVrvkvY0QMmNjERDyWk64L/x2yHQ/LheZS+09knNXM3Ir06OW3
TSmQQVS4IFLAqr1AAarQLB3z8p1/de5mKwBAtr+VO7YPsiHUYQ4hr5uFWfQJdTA8
7a1oX0xXvYeXsTy+KEvxqTumjJwmFVWnjQbC3iTcqahEhvelyTD2vswJ0AKll8r5
aFS3SQkqMpvnlDbGVGnVhKKpqRTscSKIlUcte7Fp18AA/2AEoPWy2zinM12/7yQg
ihMcWDd93rto3Y2nrB0ena2cYuzyXv9HIHmZPxNBuD8feDnfgW+sKRFJLOAO+XR4
3chZClJjQ+pRpAHRFN7l/2HoMxXdKQlcWU2eBU3ig/JTRRetny2oGETXlVAvdgDk
MSqrB3Nh+fX2cXFHKzPQCJgIzRoSxRT8VYk6evYasSsKBW5z/PJZoo5UrszsoOiq
8gbqZr2qqVMfdV86A7IV9IcGPouJwpZBxXtn04friPaP8yWJFnwxp7MMrNpRrjfn
oJe9iSpjcEME1Vp/tO/v9z1YMwH7T2BXRqzBZj3uFdymcbaz/ufGk3JgfEeznSYF
alJNoO3TmxioDi/L0VoiH+mYYgz/2/XvXtRTb9ACTQudAylnKIOSrhfJrCL8TO7t
r7sidJ2CkTg6uL3tS2mhxajlqBTtYQZRi/wtGsvhsIf68LGiRL+WF6emOUMbtTOk
ddSNDsxAIRIuWSFmHroigQV/tIkzs8ppQGwSk48wg6ZlaJC4dtupRYcym+paUGiX
kSAWommUignfZbTucSei3rMgvFaGuPt8k9g/cF/KLq8MiQfojmzI3JUjBF52nFH/
9+NXdcoYnt6WsmhME9CXLLsjsvpakZYIKMG0QaCkAK7xQYzsPKdczsICUPibZJuP
CwwhNliim4K5Urd1E1tLgkMiZFZxCidt2K/2toSRaoVDQYjNJHANuvh9b85sUi8s
QsK9F3PIf1g469wxoPPp03UNqPGlfxNW1ak/Kb1eARBZEjBFNsvk/cQBqzyEtFDV
YkU3AOOcxTS435yfTFvoYDntkAzEuKhkWVdu+LCfC6TESaXnVP5pxNQb5RnkCDHq
GR8AxRWsTdv13HD2jfSd7Oyj9Hp7FvBLd5Gs8Y0qKXvLxuqvKzfpLCkej07BgBud
ISd+7q/qPeTr0sbGpIVJDqG43aQjyqJB++U5dBJaMX4G6u1ZtGClpGjv+9IVVYM+
pjkltmCJlLoqMqVAkc3En14tRIHZPuP7vptAetmgwKhGkRXVfBmxwo354Phx+/fx
4c1JbflkiyE80LDYPNguNDlDenmIlgy6xbUrp8Bp1qJJ3ey/Oo0aIOe+r/qW3FoB
khEk3I0LgCl8A4NLWYyLutXzw33pikRLR8LUaq8oWGyosBwQZ457xLIH+o1IEiP5
N+QF9gth45iy+zJkyc6vbiaaSDGycDPduZsi3rNJF6Ygw1QJkEPVds55GRO2RijQ
/4pSFZVElOW0iC7OxUtw2UXAzpnMmHJ4m3rhtscRb7sQ4b0cnf3CUJ5W42S0tZrC
NnEUcx+5sTRZYYMESJoqedZvjOjHFhAxlnTwGQmiCTO09FZKqkdGb7w/HKd73BS2
yWUnqOEguAMgcdJmd5AMXqRWk0YaaUxKYCJICYFPNVzCpCK9iATPP4HTx6Wh0Jjt
Pqq1H2N1JfTR7h8pb5Le9E9YNyTjdSqzS3opsRwRqxSHr7fvpjRQCZHqSajosr6K
kKAp32Lmxk7MwVWbYc0KLWhlLoaijiF/aRdVK/ciAvTr1G1UAehHX0FqGd2ardmA
djlvfta91w+VN0orss7tWGVBJ2yKNWVADFagSHYTDk602vUECJ5/frxHKCOoEWZS
thraX8TWOd4tjConhuWDIAcqy8znIrSNDnBN6SgM7Gy9kCneU8bBz/UKVmrUtE8H
qwP+TFW8sgOW7kXunKsQsXHHD6kHbUu1toKJLrvzayy0MPiEDZZApxqAEuJ3vvT9
FrfjLCJCdZcY5g/c5paay2pGJ5PJUuKRAQE0/9YESwHVxWjtisiEwpznP/PvPP/k
6FUcYCry1KmkmRQJKaOnaig0IzMhAneNJTib/Onh47g1qneYWB3MabM+P5x+XLD7
vPXkapp70hrJs5p0SxzuLIGg1AV9OESINN95i0dLKZtsEcdXRz/9K1FXtl75FAza
XkYW4C+RcBtydv6xS+EBBX7NzBfEW9JUzFsFahDLc7Dx9bPe7z1cwSjqHv4hqd+q
JDumJTJKZ3bB32kSxDZr6B2lnu2VZIo04wu5ixPNgGIxvOOiuChSupTf5ocR8qLd
oMNyymuphmMt9eqAmp9wYaOcqG3bo1cr2/zMTdojXzWppCpGxuVvVx+BQy1DyhpS
g+B88EsODHlSwPtGwgUqLLv/6cZfZmx4lnb0QhM10/lZtAL4enJRGq/UfGxzJild
Tut8dLpm1vaFI6c3zKxyvb8+ggjcrikWkdZS3AfvIDgMLzSveAOtQZ8Tj/mTF287
dNezTkfPs+GxjDcvrxHELtk3jj9cvNkyJxHrrOpglNuEP88Qg+mivafKMPS7HEQp
tF9uKh97hFOrGdIc6cGua31usgIUiu+a+THZ5yHwjWKXG8UmZA8DCR0xhuuqectX
7tuoLUqW480dtoOg7w7TxzG0FKO2CwaTWb4efJvl8FcUwFZHe09ol6ll1K/+Zd5J
83Q+sxzZUF2EFiapr3BBbkda7MnSwLVX7usXvxnIlnw+BeE9IiWJ2+Qr/RxkVE0B
szi4WXPqk5dGDrUKaBXiI6uClVYNHlxRQu429JO60BnMwVVB+bAh7Nls6cfqRuDJ
RGwjvvgsFUtIgEzX1mzdt0BwMJh1w7pfvdgGAvwxKR1xJX424HmHSJSagadW0/hL
w7yYDv+FA3KAHm56iL+Ofp0lql8374ZROB7qRMu41q8VM/01KssASkogD0pwP+cz
7brXr8kIswq86IbrC+Q4qkhCUBker/LIxxY3WnI23gxF7NW7SbQ57SJF8FbwiGxd
eK9PSqJqxFaThTBaiQ6o3w==
`protect END_PROTECTED
