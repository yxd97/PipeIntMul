`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xpt4ubl7Whv6Bk1sOlVzYWhSW9xKH37aQjOQxi+99+68F6znc/z1Xi12J3EzKqMJ
ldmrrcDQNiIHeifzXsyuYdir3rfnIy3znOXEdXVvHyYIMZ81x3XUMEYkWI2QNhAK
NWZAq0r0bHuM0t1aia4Ceo7TF+LR+ypaoCWIO3dx27JqooMDaRDrILDmha2ymFaS
JT0JLk+SzTYsws9qUL+Y07GXVqwI9HJKfnqoAy1j8TYVOrV2uOCBVcKXW88awWu8
uhUfemofv+SbcTT4J+uqAcVcYzVONEBS+2Ewokk2Hr+LlqZeXnjSDgxw0CZPhPjX
XR0snePYRVmBCu8qIqQ66r5HmTPcYu3Gcfh5JNeqotyVZvoKKRF9J4se3zHYJqZq
pF53LVJErAKjq+seWZC8GNjmxrja0rVMkHDYw2Xq427xMeCj1lMDsdh0AEALymHg
yoKomVUc9lm1SgLL+hnYGjHxz/C1yfS2BKxvDr6o7o1i1dQ3UPczCHX7qMVP95oU
xoPSD82VrLklV+AMCvmEU3IkJ0z2x0vEQOqPuXdCVDQjcwNBEnIepMpmgCKo6A/P
HJW7zP1kYNT8GQESTsPmFhx6eiMQ564WM9jBaZgfDzAA+jFBneFJFpKhxnwljBOU
HZVpzdbDhQY0a88XP/X4/HZ2mkOuAYzw+UTcQEEfuxuGG8H6xrH/t84cnvvtBQds
mf6nfS6W/eX6usKyfoQLE48WO7s4CD2A+dDYgq028xMDuFWEs733UM861Dd3vRha
QATxSHUN4Org42nd78qQlblNclzB5BIls8/vcvttQIU+lfnGLnMBWJlWOS1BObRt
QWtgrrDOnJMkrbbsnXJcWo2te0aF8OsP+AQ6UgXE1bHZTIQ5Vm8178Gv1YX1nBfn
K9KgMwWey/ysSR/qX/1fW/+Nq1OhlkeyiKPH9JiVI6MQ4zP1puMU9bMYroBf10wX
/fEg9xyYMlvcaLMT5ornkT5K1pnCJAjViaCqWF5jeb6STUiz7HiR1dLzzhomd7Tt
YsSEXAL6UCEwl+62bHcTGT/o9+/9kdBgIMdK69lyYSYQQUHIc4qjLLek/2WWsVWx
WNluzZ6thWK/KX3BOCUcllUIrpGd63j/do0z66OtGTsz0oUdDjLAJOEq6k0beq3X
bhJ9SlCx3uEbbQWmDzh6bf7MHBO0bqO4NKzp73hlXdetvcJUni30ix+LnUmzpRKt
gcZamdwvsmqlkN9XFNhykD3ESYy9DfL+w+kb8mgwJulKmaFU1RSJoH+NI0ZL7PNX
IxxNEv+WKM+XxaiqAZrZyBOs2Uf4X1MNZR5zOAQ8NT5iiJIzairkNC64JnBapUHz
SlHKswyYr/43WKqtJ0cXZCTKwl4Oo2O7WvaZcYH8K0B38NMTgLUPRTWs033D9v6d
fKvAhJgfKKc3SLIX1o2uyNrTijNk/x0RxCPFzBQ7FIaFsQs0EJ/MaEJnd4I2G55h
8MFfd82KB+afII49WDGjo27+R1KLQgArgMALYRZTn6hEnkp0zOA5jcyW1CEIOREi
o7zQeDvxW24sacGZ4qvu4cTH0AiO1yHOb0cH6DdfIQbN20ZmuvapmXXM0tbUNjMB
FXcAidmr5UolpFJb5kltnjF6pE/0VHWtXJzTug8okP6kQhgaYLhQtxu0QxvPZ4sr
UmFs9p1ylzgryv3AgI3IyTB2nwsUjHEf1o7z1NLP59BXWPJCDU+J0OyWtmnWp9UG
U01osU5FOe+fpyOOqNBHCdmHb3zuI0Ppw58mjHRsm8aNISSEJiHFyKv0BrN9nn0u
SdaAOOUPsbs5yLyQsq+y9D6m/wn2yQ6DLLaSXeE75yZcYRIkLojxdAFR59YU4bCW
Jt8jPyGVQiA/jgmpvAYfEVvQMDL55Gwp1vyy94Apr/sUCCPqOwEvEttpCFBVjp4L
8PEkCwYj9KvjJgyZXIj/UIAXcO+OMf2W4SOHcI6LGm9IVLTnYHbCSzHnjRcr2q0s
P71J4I0FafUkg7LMsYRX3E62yns15KQ/1jd7ySkvE9m8tNwMkjyvzron152c74p0
7HGXppN7Qn7JfeG5OgVVw/du3boSnrp+cOQi9rj92VwFFjM1Kl10Yz0MVe1iZvd6
cO8A2kmVSDSnTlXqmBcgpO9h/dkSnfkVR+ugKvshN9WS+UL9/qN+gvu7c34KxU6d
UYnAy+NaG/kr9/gfTO4igTOImCZSbDrTzLXMhvKz7qlWIaBWyPjf414+AG7B1tQo
7ow+mYWBdFHVAU4UKXVqlKs0RCMH+iLGcIZQ26JHW2a59lZ60EEL8c5zQIRh4l6Z
0UYPcJiw2Kpmd51nBimIilF9XfPi8OgHVnnugluhhcpw/hRp9gbK85NduRIbJlSb
CO8Nhy+oc2+BnJ0HaOOqqdIUufLkgcG/hRC59rZTK3ukSAscAwdiDIt61tWPWvDF
dEmy/dA8/l9kyEs0nlpg8VyGYb0Q2e8HCc620G6zPGygI92H5hYAQTMkmIjgWgSZ
j6T18oVDtTwXpeATSNjTu95ckCyQIUrEHIj7Eo6y10NnQ/NMud7uw5wPhbacQR3v
NdssQyqLERQJ5Vum9+Yo+ywnlIQLZGyJf4bhr5c1J+8Mu8gmNiDL2o8p5ki8i2dx
qTAgXav9MopixzhsQmwDnj9hyK9AxHWM66T55pZ584WEgfKMFsijbionQWMyL05H
LgBmYwM7HPiH4/H4ZC91oz7krBtZrV0b6Bk7/sJQICgEVv9fX3E9TIJMyr0EhVgQ
/5rNG/UUc5HHkmt5x5dSL0zOn3kUVdrcTYmOfyaOAW2C9SSl8YKIqSoDK0oEpPhx
pD3TZUvPRsUylQvrGdkmsLxh0M7OKhCMCL99R1+WAXzHGNBBoMDrM4rmo02Fphj/
ir2OBQIOivydzX8R87tfXcVyVS70zDwy83W5x1cXwWNuzWiT1E/RBiAoaFOOssia
16aAxJ3tqZZvl4etUwvyDmzrIlhjdwPDPBwHlRZdKUeL0J1qg4EPdQOQ2/8eQzP4
zQ7u37a+RNPUxzGImxQHNnN5SxaGqcHKKVvZKIwY2P0teEDxu2vAv+ZURC0rnd1y
lJBGowO/zRmP4yEbD1z0gpPWijNxJ/AluvWTfScnk1jbLzStS/UDZJWfiW6W61Do
JFMRddKXnXqB8+MIYM7TgpiJHveBUbcbtgfPvidC8exL0aEir30xvz9FuIa6ZWlW
ufk8h4cMuEKmEvHewp92EO/D3uaunVTNCsFGScVni6+0HmWax9zM3KxLoczCk+1+
ehftZ7jXC/z0QgyAuDn0bIgFnVOdUWTjs3ZBYoOjsHYHIbuHluaQ6CLraNKF2U5O
I0UIiEmr32WTV0bLZUldqtA46G8QIWw1ABxsiAtKH8GAsMs1fw+hgYIU7XjBpgo6
JaGvAw7KYBF11/6tSgPH887W1wOjELOiV94g4myOeRP/UOo71Mz8BAoyUFgIL2Fz
rz2gda5C4A0kTx1cS3F4qqnpXOI/17Zaiu3Bv16aVBsBHOZBdP8rLszvs087OB4O
8/InDXbdYrHgKLWTrl/pL6O3qoxEAWxeSIN3f0JnAKb9WqAF390+hj0MSEVfw1g8
6hjwIoCuDCMpDwyUYc4u3ymytsE7plOj9wwvgVN3zeqvUaOCkGX/AnzBitHQO8BQ
xRlrAwdvu2byHVzaTM+Pa18Z9gRDrHIaN4ChxoXLUJ/jCi+GPHhitVeXnDVfCiFi
hAoXLTYtvcBbM432HgDrZMRH4kEikOzb7bLdk02sC9AcimyxDLPDD29ICDb1f71O
Vt2U61x3mVjUGKl4WXjq1YuQ6r6DNiKK3u9Gy+mxq1Uxy0v2iwNr2Rh6jAq3doIQ
eWLF2pf6ldl+RhvCYMSVDnjRZDxBAj9+TYI34ijrVvAzYYQAuMKjzJ2oP5hzt2To
WMC624xQATqTkuaRPW9fCQ==
`protect END_PROTECTED
