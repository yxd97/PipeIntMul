`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5yEc15cyX6fyl//WEc4Dazumj6be50upNbY1CJLOWit7nnfYjLXv+Q+MzEYC+Aoh
bl3XRlnTppXtTQhwBPoPmWBN+dq15sDVhui+CQzMtYtLSyENohalTNtYP/mKPrE/
6O+jdaY2o/ohPtpX06WDJoI/QL7chyLkq2S512Qc/sjn+oEWGsDxq7+KH6DiBnqH
joaFC+gHUZKpT2aX8TBrfzmszptd4y4fzkzuFU10d7HcZda7/lQJ265+d0tzJ+YC
ItsM+TBNPHOEsHCYjwdEkS6gd+bEuKAf4LOKwTnDUDYWECqcSZoVOJ3BmpeoB/+b
1259+6CMoepAAUuQ4QCNf0V9kA8SRvh0qGDyg0b2B+at1ImdcWQC5CA3rDJKPoNj
P2P7S/sN6FzAs+Wa0y4HQSoT3KRweJxWme/nMuZQIMSVWm27zCK+OU5ThCIh3Hd7
SJpHR95xHKwU2VKJLihSgFd0+8pzJEwjyDqsUeCZt/yK7mCfNRtzOh8WynlTuzv/
RKvblKnb6SBtHn4x+Bfsej4srpwjjsaja65WOHcFTkuq/RRKEW81TcDq7SBIu2tO
WeM11+6OqvjsX+aB68Gzwn/Wehi8dcYOyNWMypsPJ0l3lrxtpGP7nwIV0nm+A6VA
HvIIn4qR3grOeQmnFwR7PGW4Tm5DgtVtwn+FjGaV294tV6YMAhoFy8pr2l7Hve4C
U4Y5YRqs10r5PjOUx1HIvBsZG4m7KS2tDi4ySFvtC7Y0kRo9c6kyn40f04r+K2rY
xAU1bnngutszTyzLDMIt2A==
`protect END_PROTECTED
