`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ioV5XQPbsaQxMUwlgPwVleyPsH60pmPHBYpo2735+xY1eq7MpoKXZ9jFdeWGXha
ta80q47TDs3YAa/45fn39AIhjbqpCUGaqY8ps5SRbeO4SS70m0Pz+QrSE/N6vzyF
VR0EwZhkFpncVw048sYyQF5WOtZ2+3V7thqfzKiCaDLhWdgRm9+H+AGX1UHzTm39
uKfw7xIa0hM+p9Hm9+KW46mP0P1A13ul2eRFRzyLjWCPR9fRa0rvq55+TA1idbIF
JTAhWf+lj63R1/GyTZVLTyluN6MtN9XRBnp0B+3XOzmvDHLQ/MSjcy1KximzhMb4
iOP8hudPxuI4T45XOHBrlpLJBcGBNytki2vVnmdGb3QhnX0UNfQA7dK9hkBip5BX
mtfHYaRXjgWT1iaGzfkCdY8sNfdRB3yuAjxKmfETK3Hi2JGM+Al9iA9B7J45PWiv
gtMt6JIIiboznio6AnDqPpZK2GaR3Zd8YpirB0sSGSN6JF6ebU7NpUJnjz9t2oAP
delsgE1hsfk7oY9pfTX7GVv0yM6XqXnglVYl7g8GFMwnpZgoG2gkqpfkTIIe4vHp
46rWcDAxIPVmvT7t7Dbf4PMk8f+2slCuNShBRxUYhQazl4h6FHZSQhiJzHj8OwYh
Pmfdb/4RF16RXDtJAeUoFtj9OyxLtNvcKE9yRdC12LJi/8fNjaMKLA+aDzg1rPM7
Wg4KVmPUp2CSqsYZtp8E1y1iX3umsWfX91TSufkWNRvbe2NrGE8muZjnyY9oxubT
Mw9MwGMssp06jSqFDlwtGqtvYBz7hCP+csDsOGFk5EiDaJl/loqDposnvTO9k2YF
pcOKkPzGggTdpo/Co5gJyQ0UktIILA7VOWOA2DZsC7DvcDuaSl8GiQySdmabi8fr
jePR8sc860e7i6YpNKMjcE4rINkqjXYNz3fI1Vd1A78LdR4KUp4SDrbFTCAnGcKL
KEfM+JhM35tTRzG1hSf5Q9VSWCTa/Ylf8ArI7N0N7fyQ2hjLhlFF5VIngNR+SL79
JcJEnV2UfE37Ln6me6EchxPmV0kNi7i1GjHnEjzea3bCNrbpCP0Tf9CYCL1zrZU5
BT7fkpkqCsfdfpJbbaml/w8yMQd5vuRv+afI0WSCvw/9f0z4AhjJsn2AtmlrBxne
69k/QnxfjRfwZ4uWHYSalGqzqqBAinAz93SlGtdZZeNTs0fLh+vgcegsgl/5+s6n
wz8HeUHvZbKk1oODIbsSl7fu3wZlpGCIoB5ChYb7LRDWwsfgNH9Wr3ExysNRHdgm
ILGMTRhl7RTjOh5DFoY6BxDqbxkfZnQBk9ZpCqe+JH1OcN9tgD9nT9jrJZpB61nj
rfkQuYd8Xtq6gaRNcL2zbZ0NIefko2BIgxOkh3KJZEhKHBhJqIgTQZ68gNv6wH4G
WrpVQmhKsP/pu9ST6KKR3ZfPlFth9GI6zxIKLCPhZ+Xf1PavGYsp7rxRaW8kLps2
gfJm7wz1f6BaPy19r1c7nyozPX/C122ZKSHTqalnBwo4jiHWpVxkClVpfcwtaXVd
nMm4qr53oQ8Urlv+JrOhIXka/4Cjk/mVFCUnL+8e0NlrXTp7Pd+axzuTyugm9p2K
okEmanYHm1oFqwKX8XxMJcFGgxsD5IhbjqNyTOYK39TwQQNDnsILmaUvueH89k05
0xIOONRpoPsPH4cT5m9G7td2g63+cSKpWfCpT4r8EQO9/k8YHuQLRhBdjrs5SGSK
tl4bYIwyGjvXLMuIuLr/Kq3byvK15YF9PQKGsrAhJm2ICkd+RRHHuws4CybN6Zy/
SodXNmMKK8WlZUcBpT+HKtYGS2jA8WRuWKfpuFPY/HdSHxelbOlarSKfUjyMxam7
CIfBr3NXcg5L34zEhCT8VzQqH3QaVOHP7JGLVfXuAM0r2UGUS/8ttgP1G6danDtt
5OIeEjBr367Wb/iePGPfBbYmYuS5rb6ma8BjTfLEfrFIcinXeJybWGWtYWt8QUpl
pQMFDY3Z95DYY3oDJn3fM3uW4uqQfoAxd+8/CVrXPxdIwmQSEcLmaNla9f4DaY80
5R/qxgJRPwAWkV17cNkVkwPtXxE3uvLYRdN+RN1jkYvvDqWWoi+SyFvlkA9GCSqL
XUvGBe6gYvGIqtzizqd9RKyPThkDa+4PvygWQL8rAG4VCyQf1LDRZwXUA7Vlxb0m
ZYZ6/hJYbmWfCFwgdGnnRZMHraplhzKqDiP6JHMtua56qRhJhhtYEAUdJxeTVgjT
NvRruZt79DuPbDfYc6B1N6TwW9YLxS0MHNgrMj/40+aW3iwTNkAeLYgoZ7FWBUa7
FjoQKx39R+hDGhozeiB5QBRA8Fjk1VM+SQCHsQ7gwfcTRu7e97w8tbKxE+QPA2vL
6/pQYTcGnZhyRzAmV8HmdOFhifUu/9xvqR3K+SErS5KIzs6UJ35iAzPwOl8ei1uK
0f5Wo+wcCadg8ofVZ99EdeidpyTEJNqobq3AUEebjpCpfAUhe0D6Pa2LEQoMUrbB
mRZ0ilXQTfwG2tLINE/TTQBK0PQr5tP7gT6B1hslzHwLnSbHZGzqW06WNr36PMHf
eLf6lKFWozIMmRJ0bMlP8mAZ2azDwiVVcPdXMSZ1DxanEmnL67vzkKvQcR6rgN1k
BIURdfSH+MRvl1LQGFZ2eKCpx5Q93b4N4pmPJ2vhHmqFdNHa7UBydQi0iMzRKPwf
udnhP6EFzB0YKwfC0s5TQTO8xp78o4nSkJWYOcs7MK6FWHPkK6UzWNOBsg/NNPEE
Txue4NIA5SXkbG0uuPT8RMboVjDNXazncNvtsdsqUCuDGY5lA8x3rubmuBQgdje0
G3dniLlb60pb4wLZmp7o+/jCahok9mkPgyH9y0m6RCraEo7eZEmLjzVixOOShYrZ
teq3JZ7LVYQFrVW6Lhhs4RKc1SdMB/Gk27lXEhpzalndGfBSDI7X4WZcvTunuRuj
Sa8+EQIpvdMF+T+0xppq6XmJqrZ67zkNn9+w4k7F60Fzj88JO5DIttTzmWfbXvjt
NWEngRPIcxmTvoUUKIm3JHxHJ/mZSh8DE4FinIfWL4ZeiRbLFNAduUQZQwm0TBHX
oGapvPLTBh0esqRnyUdleFdonr2YV4WwI50nbmpaE88pl6+bL7ihe5BxX/Lq9iEE
BvfYWwTVGSpPlvlwwgBfX90B9ZeTkZa5jdabG6lR3ui40LbpjzzpUJBPy0D2l1KC
HjHCHT75lVH5YEI+ePKS7DWzsSd4aEfCVIt4dxGGi32BfLQ16oMsXjRWNLOzTbua
cDCPsxfAm3Vvpx0UlWjBhEUTJmU+gmAU3RJBZTKWlCNVg/d5h1ykl04FLda0YC9e
wB9YVC5H1SVxMnixTxuzTnU7zHcHVHegltFV0CrZB/zdiSPFcesBlVWpNO4AC/dk
XqU/osb0r0ocGLJmgf3yEg2YyK7s4MkxLaE6o1xVD0MMagwLF8avqqN+FTAe1bG+
to7GjpsyQI/6FXgdT4FW/qEhGNi9jAxlo7SrTZPswOFsyAV51KNpVFuV+GT0EyAK
YxG7BNQVzYcxdxCJSDivU+QQpuhLE/FO986esW4Q9lKYjzY+eha6xXE+OagnL0bn
eWFsghvC9lJSHQibp/Qoskj5YM1dCsewqTD/ZVuexKSw3wXHRIwQn/ihLcyJjOQc
CHCeTNwxhmVJnuyvoyeMKHYyy4ZOWPWqyQ/A7xkmUSFL92dGt5YQUDU5A8MLWGIp
JQbtAwYZPGSe9wV9zCWBP6xEROZUplaPgxTBSEAzVg0GSnB4GbSw4ChvCGfUfB53
vavgUYAwLp2aAyjzZbC6kkJkwtaivHW+akTpMHKxRElo4wx6j7PgNYXhG7uph/1q
t9mEZvwsJzS7QSCjKvqiSCDym3c420ldfpTG8kdzoQnqIToiD1o9d6zmQp3MFfux
7sbYqw2EmDb/nFsRab8RBwiiNdFG3JBGSuUNnMZXgGd/88xqGgCDgZYf4fCKy9LB
D65wBYGoHoWdzKIN1TWm0aLA2zUP+fSLYJvbUg5dI+A/TTrzXMey3xsQs90EbROc
idxXDyC/8FQrdo6Zg3ZkuQcT4eL7p67pRiKjqebfwTmBsrDQeiTtg80B4Tj8A0w5
EXxWxDciU0R1iRcQTuwYb5dBdAvXpqccUj1gLudBhyeCHb2sGjHGJcbl0Jwz1O+A
8sQgANSMJuyHiU+fKHc6MAoahtGjRIrj5RI8zTOq/89X9CVkR+MFE/jsVs4q73k5
MTLkpBkrrsfc6KjsWFV3lTEGJ6RcifEUFzhcDTIM8n3XNR0YxEkTCS7o2sROXspD
X3x4IRlQavUzu5EHHkkf8Raizxvsli2pQt+VIVSCXxv6iRsuNwFf6qCNTXz3wQzz
FX4f+oEU9gZ+Z7AolqpVoZE3W2U0GejwSPEjOt04I5PAVKb5Tug/vMhpXszFO4uF
C+80+tJlFOcERS2S39k6YYvtdlhADUYIxabyOfcg88RO5vviGDm7l//l/kXpvKus
EVI4kl4/VAtqcUHG4wbq4Rr+dNWAlnukjZi1WCusBZOMLVp27+71EtW2nVmZQVmU
7XD3O6tc1HpaYathdvn0wrBQCscnvRKrK8rFrbqtmjmbgN1xEKZwFESGKoB6lteI
0wa97kfBobV3zMxM3a1VjWvkdXZ0R6XXQgd+KvkEDFE9jyY53g+SDRl+BXFMrIHN
Ofl4KOyyK0K+dcJFtP3yz/jjNuZoa+Auly3FXjqEo99IS/IZtJRcbWCzIobLZMiu
F0qymIyQOJ0YcBYlqTUz1Ar5pvyfVn+QHK9LhsFM4PuvwSXWE7GDjHvsLOriZfHE
dt1X+qCN6yH2pTs7XroKpUQJvEasupcO2KpPwjaJbIdFie2EICcnaO2ls13Udl2v
f+ebQv8rJOPWjT0Qe1sagV4cL7Seh7G1XANcuIKxdCGtKLcNRu6P94DJlZh8gzoD
GPTFoQp7yf2jGqZ/fimvxInFnWnLg8lzhCFv7N1pX70aP8N1I6Y8ROkJ0f9Tm7Pr
88reg9foAlQk3BaisiIqiOLm4J3DJKPC3TXkzcWmEzgjwK3EaaZd3pEdwwWQflln
q6YIkZetHtDPAZfathnlS0hUe56nA1W3aeiyXiUI6IKCIAKRo0xuGUq6VG7R/mQA
bVejMM3uQ2XIezkSjra/xlCjDgnAqBVvbm/qJCf7rYjd3+t/kGxvyL9e/J7FKTtT
l9mhM8bfFwe6DtAXGOqR9wZo50K0GFO3qGcXp14j//oFkxJFeT+gefPjbIUaQR+u
TeEqQKkm9rRh/Ha0TN7zK6atRHCwwU7pK2z39jzfC7pD/qVz4/QLYi9YZQHFg1B9
1C5uivRo6PGIPZzmdoeYRW4QBguiwrbtT98/jfkyzuwhzKUTenBWE3QAL5u/rmMu
BRDMUDu4B+5trVunam6ZCYNflrctpG5aYkOiNnff8RIlccYo+VvLCuaOh1Jstsvf
0WVNUL8z8rKK78eQGqkjzmyEELOzt03+VzpmC3TISK5jmfq9VKzH86YabK/Qwt4U
T8FqJmC2UhvdY24VxsgO9TpB2GuveoPSa6LOmGqwAv934gVfImnWi8327pQbZJeF
62xKOxIOZxiQkcbxs+NQE1eITMjoOM4HSAqgLkIg3wBEHV4W4TTLtnoAI0v+iQx7
MkgtwojRsY/bJzlnFgdVmKoKdkSveW4Z6WKsMzknZ8joz1RwNPN3whcGiLPXR1WY
j9zBUtjGOLYY3jn0xHNR2YP4patWa4TVk17OjBqX7YIx3fc5bsIai4p8LIqy+oMB
xCTFe5fVQtktjX65luttDS93+PLHQJMqr4ftaSwe+iNfFgxG2QM5xGxd2pYrQswm
Wb37wFxrAuVDZak3sQjX3yR5axG2O4XjHIPj/Ossg6hafOkBi3TxVFNYzl1ixx3u
flDiwGhPEQjvuJrNDEUnTKVjDVBKuqst8VF7iFYtw+e0OK6uCxGlaEUAfJKkqrwM
lLct/Yh79yJ1oFrr3paj5gfgNXd4qBkDqqhVjQcr1MDxtv/0N2ZcQmgMqX/ddZDS
WDmgBBUk/fDPLqHy07TccNa/7BDcG3aC7yAudDRhd4h2iMQscM6O29EafnYVl3bm
btbMRua6lQFtwV/uLZXZZzBGNp0wJPcd5ZXV2RvW+gyVDwz94okzV2J7j/vjNxA8
Pn2PuEZ3WKLnwZPwfoePduNvNPFJ22YA24HtOO4rUr+GIfVa7hdpKXv20DU8w8bQ
H12YOmwMjKUkfk2G0BNpVq35j4gbZcJovFrrrCi3dD+bUHAqe9hIgF7PXK7N+kYt
gOR/laXFNROeiumRfw1R6Pf4XuSE0CsPgCOc7mVomIEsDr190yQDKrsqMdh1p3rU
jTawKPdbIqgTn6oJaCsaXKcxfrCFOJIWVrRKBT3gxPF1ScmcEYMngoAZq/gUVZEt
ipdx5KGi7yTRt3npbO36cWmGa6bT7Jytl6lYyvhzrXmTyuBm3THjgbVSU+sxHoR0
afFvYQoLj9bZzZ23QFl6b2mMvmpzo0qvr7c7aBF0qINXwtr52eXUIoM35XWDRdqb
HWZvtoeKhLibCfwo5AjwTmILpIXuwcEB0H8aUf1e3TI3kw3QboXxZe729/d7I1Jm
ynN+2qLMLovybHkqYffovhfeZgMFp73gbjOs7BeI8Pxd0ZZlNKkXBDv7IhHiqjzE
tyRmg/DjtqWcekgcr2M95PiuFXYZQcTHMM9eUC+hq93HKAa8gxWBJJovlAOKXPnX
r4hwuMQtoeteeLEab9zOrme0NzQ1YA4bkW3c66Qk8Eta6upL+AFAx6gstpjwzJOC
AH2JpM+EVC6GJF5+ZgHA6qnOeAKaw2WDCwVcTARy0gxhV8vAdfXlbjVPxchfBsNS
dWpo8DTr3Vg6kuyeYtorY57/xAGM+1+RqSs6WlDlaHWgMaDa+PBXMmQkn0zti4E/
yUtu9kfMEBj8dEr+naxEhyWbyGehZ+i28wABaQTgkp9xdT5VSyJUU0gITJzL+glQ
t0eAXKftCNRix0A/URR94p+20x86S+aRKypu50x0cykNedJA2eEZhfeFEi+QcW+K
PTTs2Ap1g95xfTRQQijHHy+QvzmG5YZtLMnSk5oXiFyT2JR5PwestNDdaWaAMjqp
uW/rdqsZPlOJZS0k5rHQ7pEPSMf6puw0LWZJwXmSqFMRUoRH2F4XSNN/p1VY83+J
fZ8VXDF9YwDewUw8kOezTqjK1KxZWBgpENS3SzZbayMCUFfl0veN9zjAt+/4s+Yy
eC56MFdqc8IwRdnczZnczFBHh3lk3oCzPvdH8NOBHQzL/mVGYu/LhsoPYcqZ47Md
mWTE8Uwqj0Nd8reBVveP7j0cmGGKorYbAz3cmMIqovV1XlRNHAV8KOnBv9mZM02P
pkU3jzutVmFMOjl/G5a/kZsUXXXevsnRWPlP10c6eal/gLYy4VDoN9OHPX9sPLlz
EH8BkBE7BShtb4+x5O2t/PvmTwQ86JvGcN3OwcFjpjFWxzXfz2iRHgrx9ehxWXxJ
5Xwo+Hv/nFKcIFrwiIolYK3jbIb3p14Q81qdnfudRD5MSJBvTQaQNnPqwJv9pYfa
ic6kXAK1luPXYwNgGgKRADZX6ABPqeXdlW1/w3ZUEyVmHhD+dzhRNElwiQv5HJmm
v8L0pIZUlGWcJXHBgsLVUW6xz5HrRTkx3O3OjEQ2D8zQC/jlN7xFj2JIOx+MVpCC
xIwq6BRG+2cl1vair9UH+x8OriVozTTLcxwLPGGFxgwxSwdHl+XHNSkk0p8lpxjG
Yo3RFGl3ocj9SAjZwon89ncaXyFeNjJTH0ANXpX42/VA1ImT0j4WEXZNBdRz/pQv
c5tU8DO303ooYA66UXbHqmyse+CsSLg9xEO8Q/xqU5jD+4hPLSfgLFelp6Hse6zS
NRhzvoPr4/PDpe85qrR9ZmDzy4FwtNr6aIaJWo8IovMM4qSjQ7abvXaHpTzuaeGa
Yvl/I2yvG0sL3aIWt3cWZECegha9PFqoK+mmuDHyVNmUuRniSLubjN5LRMjtlyUN
qlFE5im3ycwQz528/99VTclcxV8nQnrr1MtVOM6bTTIzGjFLLwRSG2bKmyTKajf2
1xFj/5ln2MOulJXT5/9r3jX1wy4We2wkVJHMKqqEPOM9Zs1NCxk7/Npks8bLptLy
zCs4v0/npTWfdSD5bpNPMRvr2AAc9fyhuwv4RPjoh6qC0b20Ec32ydOvv1tDPK9y
+xzlK+Fmwmv+InBNAsTpxOOgWTL3WnFfItya6MtY420dyWiT2w+ODMK5b4oaCExK
2lx5JNzdkBbTJV5ITIVgel6yKwv38Ce+huh2yz10+omPSw5DZsloyx3mffqUzNxM
kvusU5zZRsJVFZapQhs/4oy1u67wngzSAizLzjCvv8VHhiUC1Adot1jqB2DNj0ML
qJ6Fa81LFi2h3yVUQOaVhaO15Fs1AzMEylThw3OfAJjiuwSDZ457XOEC4S78m1CD
RzbhksLBzpSAfskcFjyZ80zzkjOWufniJlGiAYreq2QgP+irp4r20SyNsWyiev6j
Sjto+M0HTriUatlKtqMrLuTCp/j3EqYiF4oORpX/0M5sq6PaJ8yIGvN+I/Qf5VC7
Hysc55fWQyJF9r7TsxfqysRdIoePj+M7iOxEOASLsncN1x2l61ycs3gSYMR9S9NF
KNT5FFvI/nMDXQ2tUr3fNJ/Rn6i2wyUjwDtUA90M7FKQOdqsOPtKvz8Svp/5hcfO
zsopOBb6idPZl2fzp9jroy/PUB1+vCq2HgmJs7yjQO018B6OTeTE0jUxMnWe4OZP
kmSVugm77jBycGgTiHhMaS363tNwwbyKL4PtWbpjU/YrtQtasq2Ohxp96NXw9Gh2
XkX/oGUkE1PhuhNulXcly0m9i75CxG4jj9y3tYqAvF6h1C+k2Lg6Yg1kdnuAq2if
EWw4SQ1Ogjeqx7LcqHMyhFxNFmn5Rgz4j6OiJigguvpvrhyZJ7b1RK4oY1iGyepz
2q82MlVe1v7BaYnnrN9a+78PxVjs6KTfhu6iTOIJINLtiJvjY4kdXduJYxlgVyoE
kTYMoGw8r3oETi3EsKWrg32jHzgNdCKTk+szRfeDPEKKRCajZehUeaVntj6Xl9zn
+YZljPeUTLTYi/5bs15/IeQDX10Ckxii3+6qePS2I2r/OT/LALBbJg5aPTyxTqZZ
KILvqq1ZBgSD6A2T7nDx3vTqXIBalKhJrmihGp+QlHUcPgbYwcRoIHzoW6DaJoyQ
ITpco3O8kEyqZhLJszJTZaKNvwgkk5NnqieuJi+VC50CmWQGCrIQOjOKQZmaT7yo
zFqjNAYOpk9CeVj/LcIcFZhh+yG+49eXlt2gDcqg4Fh7uqipxaICTXJVoC9/qKBb
mf9gEEpCNNwuVaImM0IFyHEDg/6oJZ+zHt4cADn9RaldFtj/vgWAxHOQG25zV31u
rm4kdM6m/cf8hqW8C0wsp6CtZawrHD9vuOWDUlO6uBydr1L5srGqzae6YYBDrlh3
7T8/9NpK5kVyiZdqgwP1o1jd8YVWWjwHfgC0bKNCKbXQmBpVNUUUcJpydPsp25iL
2J0kmdIS4YTyCiJ7BHw2X0dJIhmNNIYnr+NuWIhaimfzfTLgN5Ts3HZL2kCueAhO
lh7b/c+9YSJ3sTNxm76p5CJxVWnD2S6LHJrQOgu51R23qfsLknmvwQ6uHQgdL6ZS
55WmTeFbPOuml9mxPXgLh+J3r/Sl1kt9Rxjvr9xE8Sl7OZE1zIXY6Y6Ka8aMwxuy
w5ucsE0etTXNfdE40TuZcsUxIS9tUE0c4M3xyy5NkR3c8BGbl2sht+e3A/DLtQWS
r6qJICHHTKAd+8W+78gMCz2C1XywrBU+23WgHvX8s8u04XEfOW6ERRZqLcCJ4fPP
zWT0wwVqPp/UkJNJ1trkKmEvOVWyYNgFuhexLRtF9uuxWQdlFCHy4zcI7t/ltGeI
ZC6eN9SPSiujCJRZ8ZF/CYs9VjwVkwzMiihtw5vULDmciPUms2TOKLi4hwKkqmVb
/8jTMg86QtnHU+wxj54Jv0HgY1HtKgN2akoHdXArlC0b7ZqaOJmKzzCTj6LuccoI
3/k+hHXoSDqrHJGztOnNLpIy6/LrllcggWRs8myweXpOJJ3e132pxbzHHBwpy/RW
Yh5bXaRLcmWsQCpPiTd90EV6BptcNyx+IyXz/EZTuAZwhWEPGUp5JjFNuDKUAr9O
LpnWmLy5VexU+1I4aSxzcUKOf+V7jBn0DUkej22tYOdzAKvTgkLzJe3M8KsXAwxx
wBP1gR7H++jriwMa3p6Ppf5sX7MGGVPpefuQ/MFUaI4tqKiMNY/Lvzz6y/Fgrxgg
V38XNTxCXLY9A1DuRXTVT8L5vTKymMWjuyc0pUTb+QDLMWVWJbPdTRe/EgFEHJlk
ZLpid+idje99gZGI2NEoJ01E3aUHI181cftlLaAHKwUhA03Q1ytobOnh38uOvWx8
uRcCcoCJ4DTX7lCbP25UuSjUL/ttP+wes2hgQo4ueD77/w1CcuxUpm5A8XpxKz+u
IEaSVaB4pN0J796u3pW9ou4zlEVIsVNRAZte19tpOWyEIXjVBbo78V0uFloGa3Yw
AkcMzR2JvZ/UFuUgyw5EoFzIinbgQMlJ3+TXaFHzMZNq5Jt45vGnrzb7aBuuWwEv
A3Bd3KEIIhV23uYe8rK47IwnRQTlcApFx+aTgZtrkpsnzWSGJiSZvm+ux56yG4Eh
e1KW8X/FkIWgSfvDpMOU0bdKX3e2gahQMXv6PddoO+TrdPSxUvfbUxhhpeOzyis8
r1GI/ibz7Nnx815dDbHZIy+Ku/FJgt6M/GYuCSoongpBRuxdA6fMfy7Oy1PE8H1t
8t0hfdOe6SlyPN3btxseKBXwlhMDHo3++oF5K9O0GsZAC94TCW5Hifk94E49xI7u
/1AQ6e2jeUT2889hfufDWn2hvT0HcbwBhWU1hJJKIv8mMH2/PDT2rsMNlsdlHHBU
JfSUJorlrL1n0t3UEBI8vurFLkcIYe3f88K17q3YqvLN5JCAF/n2ITUEWRM9a63M
DhrX5sMOi9WszxmL1VFHTyMkKIYHDhcJzVokXPo/gZKvVYJCSh9sxsLPOPRJAf0W
ZDWRGribpmFfoF94kiAENLxJWNI5Kz8miF3HVFbLNnqYhCHuUiPW+jzWz5EBBVbY
J+vataXxgGclpAY6lLsWJLZzCVLEQUwQdZlPFp15Dj1Ay7FJ+F3lXFSq2AsR86p0
r/Ry0jFs/beutcgLOFP1fnZOoxdwnL2nkFypaf7ETo0CnbQLK/eclY+kOgxHrchN
UIcSH2E0MmBwntlXaY0ty+s8yAYzUa4Le7Fg4E3zXUbtPrcxMz2x2KS9k6h00SYU
ttyoxbozPdO9N6V2NHa/EFn7NWXixXz0pXwTUXiChYBM9V0DN8RkojA4J1HSQ3cJ
DYyzlBTKb2WDlr8Pb8TS6idIONuMNy6j591LOdEqDiW8DBMuNZbXk2ddyQgbq6kl
ZDhF8D95825MC+XHy5qc8KUzhsiqBMXoAGgFx5DXGAr64BwM6eJwK2xWt+BaSckV
HsVloWfZrk8K4KUst4+jPGmH7N+ZZc6iBLpu55FmWw/BQ6ssceg/MI4SZL72acAW
3iHHqnXZ9zIebpPxbFmZSmPMv3Xo18I6wnAT8+fw7/pqsSQF557mioFxKDC9z0Kk
YHY0LGhugACaMOKRRDUf+oMCD+S4n4ZsZyrQBog2KN0Myn8fTVyfAJjGupbNQWCi
lFGVBqoYA9aFTUszELcOLpxih984OlvS6GDvRH3gL3NStQnnaOOBiuaBh7x5HMti
JKfrFPauPyE+3SP1oNWn+6aYPWwXf4ozVJv5W3jaDbaMjMmCY4VhR79HxuwUYFEt
r3sUSw0HDPmhlbyU2kd1t/c/TdQ13BZmdYWH8G1Xz3c8JNVGrZbe7Ic5MEcMfgS2
7/ORjXr2pe30KQffCUOwpYBcBTB0abyjLdiLipzu12+THLPqkAp6W3OPg3r6jQjC
f63oHxJKErWjjY4FzW57x483NPflLjSCxq/99yhGgmkB9pI9PQxIS3vIYLRlDd0p
AZlJA2ngFmP1x+qeXjwj//ZORJA5pS2ROvsgeE2rUJHGWYwy3dteMD7fIr7HqAhh
7M6q2TuDvS2hHRC/qB1gJYS1UPDpmS5QJXZ5KDkKB1FgBDlr8qhOZJYeSFHe8jMK
blKNGhdT/YsSpMXzEPHiknxzzmy0arK/D3DMEDSjh76OkMgtIUOAkksrNgVCZ4f/
pzyJGWuzv3phEMuy17nfLzoLYrMUVv2KARgH1PNBYNNcDkYV4W91dhnz+jzAHUgA
ShZnXqcFhJNXxR1hU2bwXUZci8c60l/w1MNzpkIFvWB3j9f3pbKQGAe6eTQ+tYYq
a9VoLRpejAIYOhCr2fRdtr4zHHJTBOnU4oMXW9Z8LPQoolL/8//rh/vnsKxNmBqW
Znz63RpBbQtkLpiQpW3glmTd4CagMPo1MH4hP7xT2Q/WFXckCZsygtz9b3fAWoAP
MSAzlYPGc+kp7m5ekO8FDDit4orlmT8MzQqxGgT8kd8Ha6UZ4FaW9+cUu4eHR3VB
it0YLPFnzu7pQk7UFkqrrqIrl+LDNkhNfjOSSFFHV2W9MnMDWkhpN69EZdcepzwi
r9aN7acHMPefahjSf4SSoBvmYd+TBNUf4fDPobEX1Pea+lCFG63cSuS2ZP0rdlqK
+vPkCsGbqqvgONTiEvBaFOidN5vhVfzt5InJWFTddsnxEORcCqZ//I5HuGfr1ZCb
9aUwsX6PkQfihwIllN8ApcAXC+m+HgxZTFOmBsbIhmiiz4Blk4K4E2WASj/hxgrw
/rcleeN45MpLR3x5oRrDu3EWVCfGOjb4g6HM838JbOEo1OP2gl3XTZNhh0sFKUmX
QKABt+ue8AoVAe3miFYOoCUghMUEVeysQSasgBMB4a/8rRD1JPHHCDZGgtCLzeuv
r13Ph94c0Cq8TtIwQQZcY6Hm2o7C+DIZwKOvhbfPBe3ZvTNhGFqKyPZA9yZnKDf3
cqrVvxFOUTGYFo6MXl4IzoStGt4DT2WxI7ylyOUv2gU2wSt2cDDRtu7d5xDNJ/Er
oFfqZoj75e7ytph1MCQ7xYhwfAapFVgyEjfVU6E671xiUR7Ui1szMOkJ2hK0+pfR
YhE1RYQxNEd5uL1qsqXvMLdzbc7tKcdc2AjQJTDGok2qcckk57PRsTw4iy5wEdRv
mp+bKv7g320kApocgylscvz1V/O8usxK8PXoTOymyMLp5usziingEdYYt5b8201C
7ZQ0xQltOJVlKmlkO21ezopPhATOdaKUz5E+XJ/+BjSfH8+hKV12szvXHeyN/br+
kjFYoc1OnYtHw8KcaEX8y0uO9VFrOC8fjF/5AWnaHITbgperbFaxSsYb42PI0yzp
1leb7IKz8pyoVZpCAvPUioVGeaaZNu8AvvDKjKSPAbJH6S2Z8Jzq8iYI+3XakO68
NPx9II/MTUoTqrg+u/feCvCx3SIML3ZgTGnazwcJoTuIaWw4fjjEqKyr3y1lui13
67p6Z+Z2zJKAOkaqZxjdZJMci4PyqdeBDLt+Sc+o1s5VTMj3xCXvKscTNljtzoL4
+Bmv4LXg0OZ6IZfwNwIy4K2oNyHetDldB4lXVa4vQ/dG66e1Ota5z6eMia/NwUQJ
PyM1lAjogaVoiuEfURLPDs4miWsFnwH3AXLp1DN9VT0KaJ1p1ip8rsM5ZUboYOKX
wBEF67M98rc+WEZgp4xcHJkyrgNTxviVo9NA3Blh79eR0ePzmt9bORTNCcoF+w0g
ytOKq6B39RkXD9xqUsCtYg2oDf9ckPIhuF5D5WP2QPxxNuhV6VpOSkKkHK/jh6v1
z6J1H8GYgmWWXROOtq25IyOCh0l1Uln4ti51BI9j+/XIxiJWQoi5bPj63VCxRKA8
+MUTQQHhl4Kg/Yd7Lbbb1KqDFOJGx9k50neMJVSx8ZzHmzJPovZNK6s1Q4OeSVad
ctluk5bgo7awhQ5jsVyM227aZbvaIcpq5mw1YGHD8cOECaCGU7JDIRxqMXkUkZsK
TDJlgwg7J6pa6J7yI6RHt7Fw+47aE0DTKJl4SWsrvhJhp9te4zgtgFcHPCRguHFB
3Z3JqkJ0mde6lb219wCiGQupvNbnv+P3NyjhvRkKIJHa+AGWyNBRmigauSs5UWSR
ZcZsz/1l0xRqSqztQlNxXlc0Lee+9cKmjKGTRn7i8Xi+oYb0YVbLsJ8HH51dGPcN
LaPh7vp3KJiPTBzUl9kwMRy+g5BOSEpN0TE1caabWrwlABU5yTSyGQqUrbNmPWsS
ZabEWslTTNgd7u6TbZL0NbFBYtrLmLkhXLhd3f2VMKmxTWSd6i70StaMP5J6HCpI
89OSHz/9DlD5XEvFKofRfsLB4WF9E4GIgL60vvp4xU9tyltfoudTwgBGjvHI1zpK
CLxZLPyZaKT4AvV23F3qIXACMr9gGL80bcBthj/Nu8kIThL5awZeB9olYg+8N5+f
nDR2klPeVwLWt42YAQsD1ZI6W9S9lAEV/bTOFC9HPOIsdUso/NF6FAIC5xkfCXug
4dZWP2oN3mkUElTKiFp6NE1YJDAE/6lsZb9mF+t+NH4QbD0Uz7rXbKRCjCwIFfhR
uQwpvRQgl3YdkvYR/Naofhsj2yb5HeUslDAlBvxnLRw/E/UKMZovLGmeJJe4LRRy
epfXFffGbwOI7Qyd4HrZar3kpyGZvUm40IxTfrxeQ/xiEDDSUr2EF07gLTFYXPcv
s4mFcBuBjGB/bgnAZiXvn4CAP7ENrPWyPhNsz/E2R28iLL1ooXdrZ6kw8qkTCQjf
nhSWv8YAn244hlEoqYDUJAPCKvJZbaJNCfgoDpI2o82aYKs29jZUMGZv9qtk0v4f
5M5xVrmvRjtJ/7V8IYBIdZSVV1fXF6Ck/gH3st2uT9g620N3+ZazqpqC5MC/G0nY
3zFQheyCWkWk3JIMWs0dIpC0Pn0zQ0gPBE/Gi7ffKEjCYSgCleDEg/glsDVZUS1G
+TTjsV2b5XFvIT3Qp9QiJ3ROVBpffKebEcVjZ0GimD2nYvpSfgMphG6wQODMGfZg
w4Z5l9Phm55NNmjzQtT5kQWxp+uvAmvJIfBKkiVhX9YQPFMxa9oLN/PAcrWDZIQn
d6N5Brff3RpEn6Dex2Dc3veovwff/+amgQzvqHv7NhmkPCcRDQ1uHikbecQ6Lo3p
RjUFijLLYS90YBtxWRFzkLu18R7JhwEpH6ZthH5wO61btCjK7zYl68mMyI3S0adT
L7Efrm6mrhp1o7qXfNw8PmTRKPTaWm88+bjudOsqEHRJB0WrZgzdAF+S7sGJX2bb
o2FXX2LAu3SlCh7fY91TXj3nzxZZiQkWhCFW3B5sjPT2n02wvj/mLUw5uEC23ZEh
SHUMIt1jsMUk18pRwW43H9BRZx3TtDxqZCJNYi+NEhQMVerZw9Xr+eqPmaG4/KXN
B1ko5MbpzQd/gvE5+vmpMMAmzAvU4vzpNEPXtJU7EEhMV9LGbs7mc1Gd2Q+K4V8q
hppWGcjCQen9kNBjV53CjdqJbdldhY/BjU84c7adYSsR1Pl7Ds9gkccZjxpEOBWV
YbGMh2TwFs5OG3WG0uxtYJmlJIsVzb34TZ+//pwghQU2HZ+et7YHuGCARf2E23z1
2N6lsmf7MG9/vZvlLuVxkTsX0m4eE4DRVv/rFvjZ73Ny5tTXipvOFKRdo/cTDiTt
3t7acxsYJMLzLtDYZ0ossAdgQHiR0u45OMjf2Cv9L4RTVc63W7TFb9HlqhpcRjz9
o4hK4RhdczIGQf37WrVd8KN4mNsbNUJ9WMuvgO7uu8J1/+lZbnKCM4Z5zDsrureh
LELnfWGSMAcWqXvPk6Ued4Dzai57U16ESngBmC+VyYCtwVgYl2yKkrC0VEIFiOUX
XH1WmAG/uRwfiOtYJQTi1fVpQTibPOaSAp0vrHHYcR1b1Qj/L/Ta2ZVG5qLMKbDX
22/64s+wl9kXoyWfrsC4/w/wKLpwy96Dh6nYAWuyuCEtc3zzt7Nc5sf4uyiOmkrJ
x5IqiOMliT+PB963Z2orr+sDBK2CRwKXfL1g4gkbCeyDbxjecoRuw3dHI2jGFMp3
6LyyGyww3H9zMj7SQnNFiatGqUwTkBHqeufFKe1wP2I1jXg1UDGkT6tq5MoovIpE
tqXX41zplZVDa810olB+9Vdlzmz4BlSxVE/dxHd0wJrNfBaLo1JJTyYUFsd4qkkO
3hOx64TzyV1f2yUDho43VKVexbNgeUI4xO246FkCroKhqq4PYsS6FIJA/q5UXSmc
Y3nbFG/UhpxQvIYDDZ5/+HsAPU/Au+8TgLAWRdwHVwHE+zEb74D4LUsJB9kSsEb/
Cw28iiKtqkB7VMY+S/IcvJ6D9mVBHF41jGcNz3YqyPtT+WK2+hz1NXdZSYAzVMfi
piHO+Fkdr3Zbi9B7eH9aThsAAFF2KZAzVJJJ21T9y5bWBtPaogzjFtUxV4MYvTYJ
85KNca/7VH729CwZbyLaqjVzB+acqRofyuwXaZEo3xh2/+f2KhBBKKdhn6WJBWM8
qboeEe22rM3cUohDNybpRUyq6LjstB7ZdQKe2g/yNXjazT/qzouKdo2rckj4cJxQ
LzJbMzfuyQs+b8nC1ri6alEWseI2ldVW3p9zRe8VeAm5FUETMznW7bV9b84wsj+1
hun3y7QkE89l0GHXjEPR9c+B7m5sxlWUnqWvmZDVbTUJt89xmr683EFdszy+WMEZ
XUc63ng94HmMJQkBSnm24T3W5o3xAaAt1qMBea5tMB5eso1F1+boB1QT4FY3rEft
QC3mltwKdy0GmQSc3gVydQZ3UdVaqJO4qHhkfMIvKZeKMORK0DDdjKqWEJ5dbUjJ
MzLhQe48wg2wwo4ThWEsq2Uaxfaam2yje36aMWsBTUArU6FOP47ZnU3k7bq9xVRe
TxQJ1urV5QVG1Z8ZEUkztizHpIVYFx6xWhWXI8uhYrwYeaK1f9AnK9aByCt7ulrU
i5WGNrw5bXc+AxTlDEXQWujLVsOAWsHqgyaCq8l2UofDzGdomY7YV3OdkOkelbhZ
NQeIpVZ2rJ/mz6LiuaYV54azDGWCWQX+ZSRDz9OWd+GnL7NXPXsv+zBxdO16K7lr
xUGPTd9G+X/YKQGdBKXwtDE7vWRw08hEJe60TwDo97lrWu7AB1fI7R7tn9pdoURK
NtSyTjiFv6H+f95KfKm13YdlfpH6DXIjerdZokwRB9Fc9AAm97WubhZJkWEDvumi
qJej7ZAaS3lVzJ8fGy68p8pEjiKiWXIB7jIyf0PJKuu/oxT/kS+Ug14FC9zeqtdW
fu3SUfuRROLh7lFkGKRMitOw+HyggakKrtZwp/CEi9NgpoyY2GVt9J9rgo8iZSLo
v2ojR5Jf9fV3y1yWJOvPKMuRw0S2L9Ul2VOjPZF/WvexkqFFSVSmqfQOrfPCFYJW
GZs7SG4sxtptS1OV9kq8+XE95Yibb4JEcdlyJ0SGPjvis085h8mG4GmSR1aiVcWT
D1IsnRnczM+L1bqXI5cBINLgM2uSGpAD/PM5oV1exdueD0e2/Iv89iSMQ5G10Kr6
mp3i0cWuJcAJsbM8ZkFKsOzuQ1bQXrTm6KpnFnGg4KgmZirthbeSrSUo0PUuy54w
XF9WfNnwTYn9LIZD7bgkmOrR1fHF7eY055/bxOPetx8nRDnRSlpF6UwxWEg5UsAY
VqUasXyjOFbZl9ncQErs1xtVw6yq1QurJS37MKDmzFEer3O73GYYuvlzri7kjYM8
KZhC1Z+HWbPw0G+TQ09CjzGE/MeaUBKXkwGBbzU/DrinkgHLPFWl8LKwXbLni8Ac
o6QbLpHTWpehlbcwZGbqsoPA72vQwB1XR7FQhsCCqG+hczdSru5k232SgmRcaINj
ZupCarXbcVR5tF+xGEFpaaU9Q15Bb/GlXDr9pb32uJA7kvQ/v3fR2cn1S1vptAil
xo0azxwXPyEyxooxa6SYO8JM3jH6SAK4+wy/XVyGeqZbQSf2bXuvOF7cHL6VDStQ
vngA4tvTUdVD5HUOYudZifmrsrouEtNlJeZTPJVPs+IwCj1eoxJU0iaMYRXrcd9h
801lrE8nVV8bKAMhZtDj27ZWH4C5ZhdW4wYu0kBSzy+1/lL0Xm+VFBRH2pc4ybYb
u2h1Mme+oSW4DalviK612ipp4+bgsQpc+pS58ZsFIpXwh3PQQx0VxLX/K0o30lUv
7AeXdXk/jZTX0FDVkLOgGt9kN7F8oJz75VY+IiDtTPOEwHSs9SbVoc6h0Fg+s+mz
V8USopcHwARHqBw2R+K7/PzdvryqHBR9harnTMmzlGF9ZrOfmXK+YxkWIHJZc9NE
8l7QUgMvjFM19JIw1IJ0sq5DxDGeScXfCMvEL8sQXbzV5xyQXmeRsmQ4TJLDvAQc
YLLELRUPT/kcU2uROd4x411WHwqOGnpDKIUSyvqA2hGFitOOukiNJ2AEt5tPG2CQ
UyN/ctAsnt0sJlmAo5EKgUNohsyqEdqnSWdwefmLeN18u/leetWJLMOgiirnl0Un
wW4J4qSTFkJ3nnfGl72Ts1v/VQ1gvE8SWk9Je1ZLf7AYdU8B7WUuyvgUuZwhKZbY
yFRaFOncsYXTdAI4ka1rvwlgwAGOsFR44Lsg3Bmhnt13PUchFJsGI4Wpi08eECA5
+0F0LYMihGe0hCkwkiIo1FgXoEjUmR6wf5LROfs+5VEWuORCXXSJQMRdTN7nebBA
poYphKOWkPNCy22Z7ZJzNKMO7yPyzuEYgxD/CFmdVOKPJQ3WR66tslduNK/I4T0f
A4HqkR+159pv9HOtExoHGKnrTVXOhrKuZwyh/iV7a0hnE46nXdd0QiCqNGMEP4mp
L/mHccV7GH1TS8MUMbAqBtnd1qh7YY/voISCXBYTRfNV9ba1aONbveOpvhg2Kc3e
GTZlUM9PA1AVLegKSuyGAW0b5ZG/Rr1693T0Q8QNv0HsABoBUwOjZQT8cZkLP8OH
SoFtzcyzB7cgDmYEhvknouzAHa2Qo3k7/peLjoIdNXmTwQEA6XvBzBF+cqF5ilqc
ZWAb7hemR8bq+68zddwHz/t3izFGyCGI2ZKDIhv3e+wIfqjBO+KajzFz/lwBsnGR
uhMBafbGxZf2Yj4IinwaBXcNEnexZxXtSxt0yKbInS0b5z60kg9m7pI1XWm0t8CJ
ke49v/O8WBG9JAH3/gKkAo3SXAbUdAsOaHU+jZcp8F9OtOTl/7Vdzc4AMpSMIqcL
sEW6LKFZ3DKMp2zDkxvtMfkVwv4jcdyX1gRt6tJcUPMy78SuaqWCC+mtmOHSq2p9
DEZSL0oeD76KBDVJtswtseiDwzhxCZ7ItzgfRHJdeJCv+RK4r2Jookrmz9qdbHDl
6NHeMWv85Uy1ShJ5uI7qEUaTg4NLxD5sqJjs0SoUPfHaZZM5PRW702fg9tGCHT1F
43I+0v/U97/1oc4e915qnE8DNJ0jvLnsCkZF2tWzoxOQxtaMHNtjrjFthM+BuwoF
OCtqfp2u7nF4B6U/ECFkL3t4s7H44xzGT1bt3ZP6xHu/RDaog8NqsBb326bcoE+/
72Ek00HI1gQnEm3QDPVX5ZukehcA46XRPABcviGsRINrD6YMlYrVLsrNq7quZKq5
/kLkzZ6a0y4gs96KZZhE+bEfRogCSKhAXxbaK7GFw6mS8bFIKSD95NsvtEemjKOP
RX6gsq3PvtYSWmZXKM7f0eXsHoQVfZ/IZGEbhpQg4z8rY8A62bRULrMSag8gZkQl
7wS4GK/WlB90YrssmAuWOuuYQvkXcRUm49DAMKjxYR76pAow9DhLIkDhTs6uL/u+
AVaf2PZLHCkc4xXa/g6m1+LloRDutnBdCfZ2i+YWg1JY7u/H6cxbRhzn9OwhpWXw
TBCtYWC0YPzzntpU6Bj1REmGOvLCrDkiKV1xuVyXofkLa+cWYGhkcDkBC73Gv1r0
w/6m9RhNRYf50UihS2L43GrO6l9xltXhoLHYRbsQfmnQdXrSNv2PlXFqu31lLgQK
d3tdNg4/yyiizPcAW/E6ZYaMhbYaW8CZLc1myiU3AFM4AQNT8NHcJ7+8PwBHGwFF
oh0Gxm8GwNBMGcyTiHux4W0FzlArLMfLyL8nE6F9uktDTY/Dcjau4qzlUTfQgDQ1
YTDqXKPINN8S2A3PXd+joQ58Wz6pm3nXIjE/HEq9LWrTTb2zJhfCPKOextIsr6vx
1ngZlczbshzBREB1Ps5nRMBpdk1taKY5ed//h8ll4b0pN+2A2U64WHbF2w/d/8d7
xjyzaP0S4Lv317Ka7Exj4eJ4bpWO6T4BKSH/9jvYoMoUp78seU/CuxBDbogHUT83
obbHA2kGvHoJoxdD+MwkeuxIlv6OsSeppNWYJRrwfsaQDTC/NvUvsZtA9t1b4D6B
TArUNZc9PnXSg6QXWPi0C4HrLHNicswfY4qMFKT9vU4xp5SbedbhVu6QQbO/EFIS
OlRL58aoJDrAA0RNW/EospFVRTlsfaArtuZoHEifbyrlne9RLJd1JkPKgNQ5Lkir
GN3DwBfGvQgOw2dn7l9eee9DrUNSb+d7+R8LtnRGjn2b1+Pc/SyR4wFOT99KXjry
JmZ4JMML54ZDS1VGnJBBtV3QPQoCXj+avKXUkKVT3f/csA0872ah0TX0DKG+O9Mr
ytcuwB1wIS3laXB6cd94ZoVz9wzJZJXh/LD3yNCC8hhguE8Z/n617Va+mc2tSsCt
lJ7ztuYLGYkqSpI94aw5zY1z++cFJNe4xMAwKyEHwlvHR3lA6IEg/mnQ4TPPw38M
0ZVS5wFTHcRBlSWwHnnqZ++8q5ENWZ5BsqtFBuHdjgoM5XRRnj7rpuglW9QQDEmj
EO20PzIK70PwiA8i4b9j3j0jC7fw4pWNSlG5Wbt5sMA1KB3qWa0sOpnOLw/epRjP
Mh7bx92Gilxe5e1a7VtIQWCXY/EBAf0LISgLGz8RuTI2nRjnRsqrkNVjjEIGQa7p
JOLquRhDLzD3+zWbSTuQj6cwFPQZNDAPO3CythmwBAp4QH1hPMqkDnqsmdcPOoGE
q855wANWRv7ayl0ybFJUX4gcFZ2g+UO9OudlrF0oSOip95RRI54qltxhWBmm0wOY
v7fC9EYggyMrXthj2DKTVgpRQGix2rgYU+yZbMKQm+6yvevpfv1hKx7xh6JhI+xA
zF+bvzbyHAgPfcb5l1Kin6sVGVwBaPom/wF5RShUutF2IjacormADpkOm53hTIOo
zizPnrkJGaskGgDNwkdjDk780zu34Z06tVHcCTV/WFCBSU04T1hXCW/EtpIo3xCu
z13Q+ZaUvn4yjuNNw+Ka/2n7Xr4DS6i1+/aqsLySOLQYJqMIo+ZkCZXZrUX7Z4/y
2VB3lVFSiUzJ5deso1PnCj3Sve2QRxH51HHcptK4cZSwDjQTte/IiflQXfSd6iUQ
Rdq9s6OzZb7kiIRlBbejWvDPHA9/mvBsFcvHBmIXNuGG3Mvdg3i0rl2BhQTVJlXu
O3PziLf/rrltQA1tAENv4TQg0mQiPM8Jc7FUtLt0aj4wpVbq+Xa7DHHc/cmiT3+I
dYMXMEpKOwgvCTkzSyBYxB4ZcFPBNWXmtVIOFwTpPKE2lc5zm6JRjbG3JvQM6mbN
m0oAMIfIAdjNXSWHEsF7I0LClE+S8smtaGO8hXfoM9PG9yfhECMzjf5abdpXg7gT
MVmJGi7z97ABXsaaE1bfRGyi3d6/TWT6uEJlvuoMDMAxZwSExYBkEAwoT3rfnGim
b8h06Y//o8Xgq5qumoI47h3xP5I6DHsIEM29W4IZk4bbciJzZHOJ3hRhRQGwFAEk
3340AdSakRyn2QB1Gd3LGNEjo/3cDPgjkchzDjXBy3B/j5Xs8CEV45y2u9cZnwuT
eRMje7VJLzxbY28vmNs9WweGi9ZoeFG/kR4mY7ibHbVprFeuu7DVGhpKWI6aW94C
BGuJ6T6mVdsuxtsDHf5mJTrLe0QnWU9KWZdzfHvY48IkJGZZ+ACMXqO2QeGsN5cq
zpid9owcxOKQwU/QaWs5Ix2V0Yz0yb2J5w6d5MQ9Qjwt7j5dJ8V9jrM/Y+6c068G
zFvRMsf0i8n8Yq/kKVh9gMs1ea1kqMNaSQ8mcA+FBr29qu/DSKcBus0AGtWWDVyM
flr1LwmS5nCRbkUeAaHZYGpcC5sVKjXTs3hODg8UgOlE8WVNSyI93fJRvzCJyowY
VA7SprUocKMasqFg9O/d7tM0jyddzYOI0oLivMuLDnHQVOs14bBn0LoGs/M6T6FN
QV+5eeuod4WmthGnrdtqmxhJvrmIb5janvbAeKDeNCVJz7lUT12AUIWLEji0TZuz
tQNKWqhJMAEkYNvvtdUWvfr2QKnT10yX7j/32ZGMOWgA3V2+1vIVSQ2CPnhrd92k
nl3pncNeLsB//rY3gfu8s9XT1yP2qSauwEihNRXQblOHBUlkEkKrFSF+tNWDx0R+
bJpeA00csev/oKbOGjQ4CSUVcQ8vBeZZsuLgb+r3O0iMQGZohTyhaRhcjfsbe8DS
nVX8DwfFc+Ddtb+u2lYqX0d5hNP1MPk3/Edq2yx8lR+PRZhdSiszeqdbrXGc2UwK
R416WGlrD/T9WYcCjhA1UkWLACJdzLfDVwVs3jNJCkjIzVVG3dKEVQo6gosMavvn
vQpjuYPaDqmGIVLbaqJXihmgNwxB9BzYL5HCZfqZ5SzmBPH2dBTpZfd9yqCxBEER
r++gRGXxSoziUn4hes1JjVdwNXO/j0SrviqLLYolgkMDEyToJmkofMWfcZt/aE4q
MrKUGLSKcqubSmaKmG5+VIOHJTbo0h17ttQcTQRnciuZcHRMpGR1Crc9Nrn3vZwZ
Mev78be5BItvKKznnbyvDaxTs28iiCxsnVghFYj6jyj8t164afg+X5sL7LWn5c4j
yKZkY8l3N/Gprla/w/Q9P99sALcxgXu1iyzE3vWILIgKBbPrwv/QAAzKKq6bCIJV
o+44R0U5pjf2jcN8zQdqZJEg65lhX6vu65pFdhjgH6BHIsZd70ovWtYvZB5+q2i4
naHAwVwf2KQYV0lfD6re8z+GivFPHb2mhgP8axbs6guzynHbEyT9xNZpp7D1j2it
klcXNSsxPknx9n+5mvJHsqxS3N0OsJo2zm2Dg2Z+mUX1OFr6M7MEkRkLibes6DMv
h1x3pvOGVoudGsV0NJy40vXyUOcvduxX6aARE4aMZo/tNB4KjQZDpD1MIzaIPhnG
ZmaGJ41OhkfpzBm+tbWoUDd4qiCJGzedvdPZvuFidNKBwLwvePiL1TbCDA1nEsgJ
GTRRUGrPt+YfRlkNGhbuXA3yb2bOJfrunMV+FEq1R38BjR5NrKysAhf+CR8L4azo
iYgXHNnEf8Od87dr9FhvJpYS13/rGGgxCiicdy4ijuP7bzsdcbqWA+qrN/GZbgYp
6REkIr0TVNoeJZNujhMAmKPiTEBZ3wCMv/W9cscKp/12FOnVW8NnCQvQ6s2O9/Gb
qQNmnAVPQs3Ime7sgXTW6w3GzifxEHISLSgJUk+lgqX+OlVzMXRhJ8EcPZAcM1B9
F3XCf33+Ogda4MWlic0OX3uMrZM4ekPU+HUZFcrNhHmmpk4vVkhQazAUJluaVbyV
d1sD9wqC4xGKyYkbtxKuzhTrGTIC9bQxLYc6WYQK6ZqZ6byiuQrNZaZ08jXWRQml
6XxASlUC0yA454QFAlAtdfQNY0sXtD+/FBiTzv9oInjv4nwXN7DEgmVDv2sNj9Zc
F+dgH4IaBLpqhDGV4/28xVX1MRwRnPq7b9s5rlI4A6VUPoclerDIkFw4XSxSEWyC
2Gi3+UjUvPEPVMEn6en+Cj8sJIpEVTZQy5F3AV+OeB88NJgpyyTttNgtIP+B744a
XTed3EaQZaU8ueY5dU9IlUi6b4cSxJRdJCJUewmIPGqEwb+mOehogEZnlk7qWhhQ
33As6R+HsiKLtE9mMoS1BGP5agdcv86bV2KYPgXD0DUBloIC7RvBs1dRyuaw0ZHr
Vaeeu3l9VStZFNdrX8TzDa61UN/PX25FxQgQxzSfZUXF/BREezZcdlOnX3sGGUuo
07aV/WFT3y9cnCOQei4lYPhf9c02QG6UBigLvn5h/bDNPVL2JhUNqhMjYSr8ws4Y
0vR4CCYqW29bQEX46G6+9rZgJeHjlncg7AlykfN1dy5qFW6FbFsMj+EvpQppbvIu
kL6DEA9z/yfCllPx0jgXds/MTVo080v4yqGEJMXU/a/u03C9xA09CH4xAhw/ypNZ
CBj/vfyfkNjua6OBq3T6up+R/Lfot5jvOl5pXbx9POVcwKkYEZj2NvF5fcVClDp5
1I79jrhtg8NsciKZi56GoQ+ZG3F9KzbAIChQy2zPSokrU6PLArG1apieq2QwzGlI
czKjGEV4n8Ot59oO5ZsYhrMJHbjFYjG2+D2mVgQdfD0IncdU/oVru4sZEzhz9wtP
nPfT91rBV+t05SmJe8FfVZvLLm8op5Lxg6ObGVzdqyKHqEROpV8IUe00bXgQH4GL
i94jAiLyzO9h+dsM9FYWjXDhqUJI7zv0Moh6mwWl+D+HdFy1sVgT3kR9mrdrLKy1
POGtDmCT4Sr4wowLEPAh6BW+p4UF/6M2boEvv/0finZ66j6AaaolxGuxZuHwQ9Jy
j8Ypi7BpgyERPdMYSy/kIu82hWZeDR4rEFaL87bUp9RbXLJ91b6SMOO4Pq2haV7l
BtwVAzerkoYM5iCcyDz/sYZ6sYQHC9JoZ3A13fPwz71ixVctRcF61xHU27/V1huU
ok4AJ7MTeN0sLAowQItVYXAEq7ZcvB+9/SS7LY85or2fUXeeh7gjcu5wZeVtdSaU
q5Qw54Lug4smaT/13LULICFFPpumzyauY8koZgFw4mkeSx+VIBRyEwsd3ubzNEC5
asmMiF7KVqTCR6/4z+PAlL/LIp/Is2KZo148Uuria1x8w5cpORbPpnEL602NV7N3
LRoR4UlVmjoehDz6knRbtN3zTpchpRi9CeIzShhQGf73bLICiEzNRNS9TkS8J8dg
GicqByn+hxbjtPr2LItFiI7edKrRzygWrqNY4Rzvi+89YCaGDrTplg7kCD98BoZC
cH34zoyGb9hqlir5q18uWByV1rfkQ3gsY/X9xO6C52QoNDZ9w/hywwof8j9VKTRt
7jtzuKauS1zZ7Gi2MoLSv/xxy0xRqck9dRCA/G17h7Keh8cYRPCTRdGoCeBr991M
IYemz1qffugioF91wOuTslUYjAnw+oMDH+FGIKHzNz60O26KtfyuNR04Vb4pAzgR
rS7DdQRtuxegiE/6Uexn+ZYRKueN325IMXC3NN2dwLA4TF29PqCSZ/cwTiyX49+f
wFjr2FI9aQL/thoxquenQmfDAKTI1ll2Z+gMhq85CXdB86sj4MoSmjjEgGKODp4k
NZKOmBgxdBmZmzDfU0cO/oKGPRpeIwBX7YT08L2F3diAVH2k8adMVFLyAwWWjZeA
FlYOc9xnr08ZGelHELVM2BNTd6nSyY01/g2+Yp0K7do5jqzRUELTQ93UpIZYDbP+
DUZtk3XEOyS/vBU/MsK5jlcyJ4zXun/BQCTPdr1qpeFYj1gk+QLocwwT/uBRAatn
EMbjNCEAxw0kMTXmUnkCoRS3UPB0tbLAFU18KLkmJYZWMpu44/t1/Ug+dXPhP5jF
1zHLfUSG9RUBTht9bByYU9wzr9fQjmdvk+FfF+Hs/W9IPnFobA3DYbqBKwVz7e3/
LQd2KFA6DIADkdmDI83+cUZJ1lFG44SxN11QCPoZmmHMhOL2zjJUezCBuloJndmd
qVQhH/FhPbqy+McSIJGIV6Ij39TW8jN+6/kiAAk2Fbyr7LZDlWBicT/nL8rajt0z
YIYYAhQRXe9Lvgv0WLphaeHXAh/vs019vEH8a55X2Vuk/bpHZM69WlT9rIcDxuWK
DtKu/BIkID+3Q2tEI9+Z0zjEEssMrBSSkuwk2ok7610qW9PEJB9O+OkxAkMcYl4V
FQhtZ8wYruY7A7MOM0J8TI8HBhckrU90XDxzcSFUeul+gXoMYx11sJjWzyDk5kfC
FtEg/wJBIEGdeULHYVC8r6jsNve+k+hoBSsN60UGYFtFbhnxRHKPNhnobj719MbN
GFw1O5O/xEVmjXH6tiiMTdkpQRPBnuyX4gebotFEU8RXUH1WqfT9Ef3EcsGlHSPH
oYOR8g/NhAC2o0qOus2FFhbkC4uZQZZZJOgj8lyEUmcss1psWyIARga9ozo5s4Dq
Eju0XYK8uRorOl22kTRrHjXmYazJW1KNbUNfRVAFyl91AjenwVuoV5E9a6J4BlOQ
rpty6MNBAO72Y2Gli3eoX/21VCPCT+fL6+Rnae4dQ2PKTgHkioKO7In57HDao998
uQhi/02IKdGr3IWO5DP9jGTWwUIra10jkqXrGdRVkrS7C5gGrx8BoMZ783kycUDP
eHyDkomLAlRKe9Rcc0AC95cBArU2q9A3GufKUEaTtNYiA2EkLnunACZOLGPBc96C
+LlfMSe6po0mun/a5bR70orKF+a553YOIFvKfUt3SopWgOLrwOLLI7nSklaSbsY7
GE6qli6QUdl3nle6xBNS/Lb+UpO6/l46z2PxyvFnnhuaUJo2nj6LkZrdPnQDj+ZV
Y/jHXfwUw8rDxQ5ZvKwQAPYW0W2aBQPuU9JOQ1MYulII/Jxi2SZyzfeEYG7A5CKg
gJJccOPazZU9Uqha1oEaaIx/u+etcpo8pzKgi8qv3p6Gpdfbkdkj4yxPMVjGRHFn
TOEteHk7fhI473HrFJsKUmyic6fbK0JpN1WC3ZxBObaip/cGPkQ2r5GNWNoo5mD8
S3KnNlErdRUIzgFEzlcm1CpgLBMx4xWoYnaF7gJxtgQkhF/3loMLbDxvnlq/ocHe
kV2quCw8j3OPEB/fCuIwM0Q4VPS0r5kOOldwQnpl+NoUfFKlXzz125q/5TwW/3ov
CkuEV45JR3us/QnRrA2mpnanSLnEXCUqc4RRjYRE9pZw4icpVQCUFhiTHwBxHj1K
4gt/c6RZS7a1WtkAPWOR81Bo/XK3Dp2ONmKNj9AOpsiwBQSv32b8U3Rah9Y9w0Mc
RLUu3ervoCpwXgypp78s917NC7YPhGr966DDSGF4VFaI95gL/TUjSMxD4HuTU94R
iv3B8Ttvuyi57Bbaq+6u9DTsXFGJS/qzE2ADxEXTCCZdAvupZxEkj8gcbLpXO56j
SLj/9rL9zLiEiZb3ko+y6i+A8G0gT8oF9k4ydGHXjDKtP+BSyqhLvVq8GJELyYsj
Cx/2yXAN9tWeuUNDcciTdNFbxtdBH5xkcuk9vUQAsiA0Uj0FZ43TNNr0xLTmoswL
TN+5TXRhlPe8bkt5+OusK4qmUVVphbcTlE3M76rycNLLibca7vFv0faxjxxk8tXd
i1Q23+FNmyYKW1rdQ6gsuA7W1ft64Vjge6W0NGe4fJsuPepcvRDd+mnbjD8y1qlH
QXDXdKf+G7+bId1JqbbasPCvo14qmWNQtqTWIg7G0s75J+6S2o+Ow8Mb5JAQ/zBe
OOz6P8xx9psSdMYxcxcYlUWpqh+KaYh+XDW9bpZVRFlPXFZvs/KczSCSz33jF6w6
RkHi0hm9/OoNfQrkQNKSHOjIChoyF8SxqP1zQsvDthmNN3EypyG2PAWkBIfHQz6r
UPvKNnkCdc3r0s9TIb6R3eAHBSL7vqokJIAY2SLODS2Cdcg7DBh23wCtDHeqXpDf
59ziLCys7ApZfAjmbnT9Wdkf+49blEiPrw4LByUZO6O6+QoNadw1YWlTetweH0r6
6HkBWI435K35TrForj1UPHj50am85Gs8qzlnogkWDP3ZlL3IsDBJi7dpj4I+V2EO
Z8Ze6Odz5ZzgSBX1epSLJbbru0gwe2bduz4zvuId8a19FrzaTlMuUjZVl7pEUvPq
JBM0Q5CGOneB+6LO1RunIm3ihhvuEUsIZ5jm/iMYN/EW0DowgS0hVae5kV+q+wq0
5i0lyCFHlXdPlBZQ5JwMjLm2R0wLGfZHaKai43wQm3OtkIDCECiZAUUIAxnSn3rJ
L14f1QVYz0bMeIj7bmsUzhvnDWTPwd9KsApMvT6OvYrXv2AUY6cWpxtwwqfrAGEp
buI5VGh9Zo3Pz8PUcnkZ9n/EYEMka0kPvA2KB8NShfJTcjZ2cXb/hc2ur9GVdGrP
fa2o5peg7mGlJK+LtNVFrrhUQhoi7fK31vWkwNa1swN9tjiPdMJiSrE/eEsBrFJ9
8zRieBfJ01b+eRPZgnt4Q99zktPKexKp4jriFEoiGa3A2CSLHY18WUpGTHpuRcik
N1c7NgK6YD6UiGZ6CaDZQ9dl9403V937dsm2397E1SkTC8+dVdQqI+RAZGniT4wm
ALiF+TYXVOMf4nL/2rxQX6KQdw6q/D5Y4t6FqGDz3GPreGZYpt4Q/Fo7mFqx42uz
l9WIzTyIQsX3Mi5J4QexBFTtRauD70tzbnV2pO9BlaWnTDTlUfg5OSNfIdtwRQoe
Q4CspHDw02CWZ/ATZNM2QVrec4z2ZtnmZvUNOFAUkxknIrdOHswAbkltS5siqd8a
wxZLduWjgFcEqC3jifXr/+9abj5bTfSLRZlzpvff9eaLnwnfYz+PJIXlpNG8Jxcn
7t1LO1CKuc8WN1ab70T4G++aoZ3Ib1lfTJgO8o/FcnuNxPa5Vrj4H7XY0bjeF5qb
I7rkRLE9SpRh3JHA0Ksixp8iPsy9jr7l5msFisR/uO1ZIUdqce7/WqD29b1ToDVc
lNMdewVikflu9P+/tsObR3PitUvvFr2eqfFZemu8W5hvxwEGbmzmPbXhfZ4g0XSX
82SoAUneZ6RhWScxL12FbQBsbIi4ZsDEzFPimZbwzKBrFTOD3RpLC+Q7exzhVMr5
xqcJWHMUG+DE9Z+MNPKufcgUaUPPGekMnXi7LFHyk+r5F8kJPnPS4YqRTsk8l/Te
ecDecU1IUCopI2wev6at1VF7UyivvrNb7QElYv2jb/rcM5csUeWm00wEdNefWCf0
B3kmlT/vkoJzN0bnIsjxE+0riyTtmozScGk9O/88rNOYj3hUtH7itKvE86M+vdbV
AqeKXRLkh67avttOHt5M2EknFWkh02+yGjZ3vOohdSNH1SBA0LkN82EQBXcG0usb
O7z/BGvqIKmJZ+evK1jjbHP0lku3Yy8yKd/bxC3UhnQPkiVaXLlcnU1rQDXX2ra4
qiR2wK80xoGGao4InLEeHq8L3AuilVI0wrWXNBEsj/Xc0twrTE23WYexq5k5S/NK
QiKX6JsbZpW2hK9tnvKJTVoorTOvdIw36Q77zsks70FyEzKX+KFlpKW9u9VqvSxT
hNfCW0HBgGWt33VdUYutWjln45+c3W2DCiWBdad/sjQiuKu4ETs64ogyxPOMmZjf
RIkDoOPhnqAcjXRP39tcRLLbDZ6DnU5TepvxXShrCqvO6LR6UCclK5nLyySobyg8
P32OGR09GWU+TfhHOSqPbxL41Tx/ePUoaByNeoz3TpWkB2IxKA442aW19dOA2GdY
U92ZXd5ZpZqvBCCPedcF2fZWiwTaXZAaV8HhLu4f54d+L76FP29rT36+xPQONwOk
QVhzWYtjkHietYu7DmH8S911W7BwOoeJP25VCWMKLmUMUNFVjfDTSa1C4+Zpm0ZU
/gL6p2m/yWD193N5QabY0WTmhO9UE1dnwekpzcgRQ5SAR7M0elBtNSDDEqSeJBrf
4ICsF5KqRb7rltx9mIJ39oCzzd9p+AiUXtq/2X5oEeo5Vr2/wsQVVe9ws803H++u
tfzm0pqvtbM+0oMEfIn9Hwn9OGgafeg7Ha8gXANP0/Kk32wsEF6s7PscJoxe4Yx3
+F1UfUTGwDFIh6a1qwzFRl8HnYv8ljf/jFpQ0KERQfe3C2vSlaQnBqQkHozU18Fj
fEX26+gm0ezFxDRTrO3V/WtC+hE8EbqX/zHcI+FBjNVFoENDZpoouNuu2c5MrnkI
kNlM35D/wKeSe9dT79Z6N4vA57cbR5EvNzgJTEyOvfyMKVufckmCOb0zsqkX2tLx
g/H9tjYkrpCD7VvdfxLla3v6EfZWOUoUuGWLO3ZJveELnPq4b2WDrMkhtOT+CwXe
zonDpDGF3Kai9PNpTg/w62F+LJ/btYZSWt9kOqvrnbQjJScZtwA5UrHbcbwkQSvW
FvKtc0yroxIhh1ZDKGGl+3SeVEJ0N3OMvPDftIk4ZKZ9eBF9Sb2Hvek/zMy3bLmi
bOU2KGPF98RvBROQdxU6X1QxtpYFSiKB70qCpTNGErGkImFgCQi1/Ruv/Yt348Wx
TrtzIra6B0HXjTEoAoTskaCtofjn2p/zDnDag6ni8SyuLuBU24tB9DRweee9/wzV
+4eIGI3GzooX1GcOibkCcGhC42hHOibCCtHpFD0ZfJ4SZ4K3vZrFPrKB7TMS29I+
reotDIhtdPgmrgK12GK4FR46u45dElLHTOJX2WIsmREsxLnbl1S4pw4g9MM8LOak
Mk4oKpXI0CIrGEmXus26+Yi6oFMfbEluxpIdB4qeamvubQFZpUw/B0Zmfk0MmH0d
C33FGH7kYeU4kPPJuNwf8QWSywZJpd/0HxP6EQwzq32ldiqLhquWEjnizzXW848/
VXt0sxb+LH4h8kC+t3Z+w+bG+Qgz+OYbmJhlLXj3jBN3JyTcLdaUfE2fpKFbeImd
dsb+X5o0gALPDeO0lmljKZnyPusl7946erfmSHqTJ4UhtMH9bjoheEInQa5UOCiC
9C+uBi3ZQad8iLJc168oT1kgRSlgWrMCnLjzAEA4HbraVvkYdPRsEJ/lLGEygN49
lKuEioMgkw6pS5Rb0Q7XVIqNWHZqkf1VjVYo07bJG6v9zinFabeYLYFWMS94Hs7T
P48Hf1QmJUXGwP+ygYZEXmDYfQUUwwtRLGu68X3tfipLsVSA8v7AofmJSyLghzEs
EsEPElxXvqsb6uWZurghr+024SwimJ/Huz3VizkvAztiAU3xcxySzOzqntrDSQf1
TxlQ5iG2KVXdnAwKQTnkj3z5azbWd0j6A8EFveWLZ0FhFSYLfKI6LU/wAKI6UDih
CYpgpVwmcuzKjucQlbNMmXjN6Hxc0VhdNcGU65tzx/SCEwX8v1TOSdZDFHGLsuUq
5UTMsUl6BrDSQtPARBkN96heEC70EfVxKEfHlRsRMt33y+k5QI/633rNuL8jztyO
ZiYAV1J1ZZpcqyEAfRLW21u0d5j8srUvHWUzdtu3s7HtRMR+Y+Q3Swduc46S7D5X
/8EeaxyyunLbmuTI0P03gmu417PjT4dwv98p5t7nEtAa4Al34sHOa07fTYsoilHh
OzaxbaPePxg2vRVd1WfvIN4R2JqFXY7PoRtFqSc7wny13K9wuKSD2sELadniSQYJ
FCwUd3fPPOCh73pCWB6gvz9KRU7xGl/LzWHWbnfNh+nvoSLLQMBVYEKhtyvfiLrw
/RbyHUf9WnWG4ibWC85ws5x+Ar6GLHJJXoT8PriQzU5trSRBkP/q63j99xgwp7qb
iiMyIaQFtKyij+YvasOnnmR43Nl4yXycKrQT1Xk2TD6tCH0bYboFyN14eQUnosHv
PKa7vCEBDipNrqlqwyIu4YK7L632pbszm3COAa15/LcKrl5yQ7XRQteljAyCH4Pn
2XT8kxCFHXsR3hPZi5efkSP6e3mzu2slYW0IgpcTFC3ATjC8xCvZQYpkN90hicPM
9Mxt8D83dNjK2vDNfUx7LqLwbIyZiHDgHjn937FYpVi8ylIKN1rzXWohxWCwhXUa
Yh2cGj3iOm0+nQJhv9/KeuvIoqelmiPwXzxM/asnze5HOel24hE5Ba4t7c6rwKe0
SjY2ONJOnWmqQ7lEPTm/0NbRgEoaz3ABToLqcCbcG3IosFKVwaV5IBKXmtps0oSA
C0dbAaxhLiW3NV7F2T5LhpsgrlbL4gjTcOXvS8TYaLfrDc2kCWM7AI0RfNwSdH9F
R1uudn8aWvDOvrEGKVibYaQeh3zn561ASSlVj7VrgQ0pB7HhPk+coBpW1TMqGOvz
N3SiHONAVnjz+Fhz71pbY3lESl/bHPE/FY9fTg66f3HtnA+eg1lQxFB01jfH2tmv
MlCnjEuWi1L0kC10kaz96S65TcmrEOuiaUP1SLVDI6F1jKz68pVJsI5hOlW9Mkpi
3otzF2MWM9Od+4N3X2td/Ti8BtUJs87/yi5JXqKBMyNznAxZiYFtNzcSzHKh5EvK
022NeYU1ptj3z6CrcWg5nDTVSK7imh0nDs3NdawdxUZYY7Mg79+IKHHufIp8a6gN
mm6Vd0rC4eKa4kUeQD93xkV89RYGNDqk2QvSD1ZYwhqaYwUV2xH4VLVuZptkv1GF
daCXXWFPFnX+kPhKnwGVWDupjBEAA45Myf/HUxsZ92v1Api1Qq3cx4SkqM3tLURc
T1ID3KZW3ZxbJXmVW1qctXo6Kd1NH9Y8DzCb/FPEOaSkVsYlbeUYaentRqj/A7GE
WFE4VkkpKoLoAB6cO1MmidSt6al5C8lCWOqXyucVcopZIVK/UA1emRyHIQK/TUQ9
S2fPUmQPhzK21JlvRh4kfI7VDWz4Yg2EUszGy3iAazNtrjgflWq58ouaDcqsVhDz
NY+kcFXfyubeQXYad0rW9mB3pj0jp32gDoiLiDRFIXmqyYpitlwSM4f954ZH1kh+
hpnlL+wVPT+qqDzfy/En3wDun1R9GFaj6aeE0IGMxA4sz6HSjg8UPua/1hdd92pP
1pc9XDQLqcq6DW1LLC1KeT2P0ycv48uQvqr5eWhD/lLd0/Y9PFXJOhfqHl0vK2Px
+psXIdjUzkLt25RwGCZj+sUEj9tePe86+HF3T+R7PY5+kwsPgRc0MH1vmFDM7UQX
UcItuv8tGEjFuXjbE1QOb1AIJUN4IrBvm4M0jZHZoJo1RMl8noxzLNUW0VVupStL
78Min5GLrwx6cU7oO24XdbdI/C14KHkQHgEQ+N+n6Wj4NdFHVUJg8WccHFK3oJBh
l748DGjSdG4PyRQQXELayZncv7AlPYoFqCM6hH6q1zyz5OJ0APXeOQUS+hXWDFus
i8MyY+6VeM95g+irspY3raNZsdHU9yWl0eaPRzRK2/3ieoZQ3DEjRSLxAa+eBpWv
2qRE8W3oDrlrncPIKjm0jfMp+/XRjk9pmpKM0kmA7UexUpcmsgIN8D8hwUlIU4vh
4yihGIB1xSJrTmi82CraXnnbrNGsUArxF1/38m0meVuigzVoMglMCAie8xLWFktr
6alvM3Toryjg5HXaAaWZ5gI11hoLeoH+GahO6imDdPK2KI3L+SvJ8tsMKVoD8k9f
TJPrcnOcWITjxZ5kDwWjFw5OSCjEiumbeXcc5N2g2N4Yy4SGtc5YmTY5W4OwZMde
tAyEact1HSgs3qV6dr1f0MY6OkewtaKCs1R2C1P8/MGOe+mIX6cMPDSPACRACAwX
j6sf/iDk5K7hBo/pyKNbOkeaiLGgETkNpDzYviLZkB6/euzsW9eIn8Wzx4GyPlag
46wDA3BEnVu+loLZpfiqDRDduedEqkdm/3gqHeowdr1zB9jLzL15ogZmkI4GOa6l
Gtnw+GjWSE689FUDigzSCFDd0QvMMMFp7nrV1jD/RW+k2goPxgdicOO6MLMCHVF0
2BeRAj9TXgPkfMp3FQMrOpaZLzionYxvSFboZJncKC+F0GSJjAilOGgsBDORlJb3
DrKAuuapXDwTjHK2tljWyuhOckFmcsDlallxUtiynqezdWtrim3nuQak/t2s65Ut
Q+ilnWLfj34wbKhm5PE8kQnlPfO4Yn0A+RnyBzIewdjxo29sl3egJsg1hEKxb/6D
h4jezTjijrc8Of7wo4ji5E8yX346J/g6tCWD6IGyy9wn2qF6NHB8uzIXsuVTAE8C
TjqbnO7cVD4QBDg2V2YcZfBXgN/YanqgOI1BBmFYNYxHsZthp8Gqo8GybmzmvyLH
8VDfGkEJAUs+ornlVLBlitK9t2eHoIYp5Sxl2Uu2LbwAKiPQCjsewPoVPci7y4bD
Xzlc6/FFQ3+Z4JscwiiymRHW1r2HwGhJsrIYPPhhSRjQ1snkFY8x1VWuFhcILHKh
VhEugGF3YEUSOcmmA+HRGDjrYH7GVTcVXIr2GLh5uh6aN1+quVsnCfBE9NVm3PSe
DoRCBcwTkTkP1x1t8wdvqyAvYtpxVXCqGlIElKrmv0PQLB7vIdCpEugz9ppzIZfH
9I1JF/fg5A/lp38LOxR9NtR9hhjmfun1/QTNyqCO1ksUBX5fwTCuB+DkZ7qo7tc8
uFEX3SYL7AjBKGH3k0yBawWL4WSRj+Nb9FhFY82wO7VX/s05rSxBLZOoI9lropEo
Lpe6x9j/8yUvqoEPty8n0HljJB8DepJLzNECXAfWJq8FUADjVRTcmqzHi4Ina2PO
4oGojHri6dZvNVBUxk31aBOtGRJHnFaUoi6ETfNAZ1QWE5Z8K9zvjkDnu5vkpzG/
VbS4SqNoAFu1G3EWvBMZiyuegbEWrrGi78lH83BGA0W/jyuc0/oQnXHULAkN1Qje
OXw59LooNEJFL68zdh9Dm8ZGSMQ7Zi+MsKVulV7f3i/zO1Wjon98PDQzdYbcRH5A
9gy9YkHq3gXUkwBm7jNCzqLyMiS2x9pat5HYOHRnz+Izi1+VONXsmA0PdkBstcFs
M8TC0VXfGW7xdC1kjjOj2DFbneaQ+Tfv47dnyYugNzGPRFweo1I+Ju/+SKZBlYD1
T5+6/eeS5y4BsH59M9HVhRwcIu/16ejoJh6KKRSYWFp044AjxlonbrAI5xmEt8e7
oyrj3PNVH3M0ZliI3DS4qbBMke5AQsewmTQt8KHyh602AThTUyI+oaY8jyb/F43t
yLoAtH0gdo6wNKS+4swPjVwJfTMLTOgdp2ehz0D65MATA+0pTqfKvYcK9Wch1C6k
0V6RVhZQ59qQ3KhQ9a8YnIwzI5DNGnJ+TR+XMhNPxpHioA2BbdyG135H61xIHPZz
eKp+5CONaS4oFC/8fh2E/l4xHJgOJR0Neug9Mj+pESRGk9VgyRBmKQPJp1KdCrST
7GPV4wzreMI+SeUT4Lgf/F781FvoLpIKnr9eqVAz+B8Bzz+j2b5bHzu4g26lLg5G
1hr0ZMa7jQNNDTixa/NGCjBv+8NLAkPL6m9eWnIJSFIoElE1Gvfv4enIcw6TzERa
b2GPDY1MjSnjm6BPo7w4V8PGyPoKnErYpTaA/BZ0J+8A5CzDOHIFhgVfUKMWlRJ3
IbxRV0Do5L9HKNBwnJ7OjxHF03GWchjLeHL/Sj4PBya5MEHsJQPmQiBRMJ78FMIj
O7pSgFGfI5lPnsFZlWpc+DO36Sdhlyup69UL/sEDuDXwlR1NAJPWGRWoYAdsZ8eU
7Wwj2JgBGTGaBUQAS5Uue03EetqhRY+wVUq0JYuH0OSyB5MWHhIAAaUtvisKoldg
DeszoU1TQPTCxgpeEdB4hfY77evqDkNiwRnH9TC1Z16ZklQ8hwd7sp24BXy5Bk+2
aptZC7ZignoEpKh0OVaZjDEyWvAh/RhBqEPNFyngCx8hkVQT/3HEwTa/9jS1bshX
5mBVlZ/5+ZQvZNu59tnVLmQTdes9z71R03+Pb3UvvaPLsRZlFGW279lHDI/+0DNL
dsmGH9ccNrgwL6s0y00Eb73znss2bFygrPK7Wj1YMBuH4O3nLt2cZdrM3T4oyAJ+
nz6w+pzn4XIYSP54lWN86h3sktv/W/vIgEr2QpXTpyyJmXzOn5btGWG2wK/JUfqP
xW/zF3TSLipKUYZ8QkHBr62ehF6GVUXLdp548S/IyuSa4ozkbvHDOuvLHdq6R2Yu
2KgDMv5JbQNo2xcDKFkJULcZieGbFANiWo1u43OuAZbjhewxodzG+QytStk1o/nQ
EIdMisai494MzyC3cU7eifDjkC4qMuW5DhtFzjbT6v41UkcOWq2EaDbBz14r7F7M
3UdZ05WvI2DjF90l0lBJL9FLh9BOxZ0iiTwePShidLCZv+Zurtjg0rrt1nKR2Lyd
lq9xHF1kJBjnVX2I0d14lGZ3CEqYG/PYjCEehVRVRyzdEgg1QUfW9hvWcyO06lzH
O90wb2YBx1tzLqzfQ/lEWbuCKH9Ll5r4Qy7ZVsVx0NNV2f9N+EmAbL07r1KuIoJV
CvZV9kGAyaRYKlMp4zZZB6keEvI1jkR1J1Z8jhbCnUm/eimwMX+MOrDw/jWchip/
zvc38dUOJa2KJhZTQ0OIo/oEsDbFeJXrozmTTpkF2sdJbTnFbqV/+RckmiwrYcOM
/LzvMCZiYxUlHmNSnHi7vmNR4sGrBICmvi8o+FIEjZH5DJIS2CKu15EQsCZu7Jnm
nVJKZwjQfx4BWT58qXjgk7KfTO28hMH3RHa+KI9F7pJtl6XLGxddTnyU2rxiSPmm
Bk+Ippbm3LG4MiDNeQEFr1E+B9ajyDuTMAle3k4fNvA7ixCin6lXsBBnuO71CzuX
REWwX9tX7SZqr8z/MrBzcfvPN6xlU2pFYX9O2tv8c7ST69TncxiJJF+1fbczKwki
Q6NzQf19f4mS0zTtakgc7FjlaA2jV3y7etQemBvWz8+QyZtdiT5H1vYkR5Q5o70D
u2iEZy4aGp+m393NLCVrRp2EX5zW6wN8DxIERIIoASjfmzTCmIXZTcQLTO0tfXOE
6o06W8RiXzu2Q7QCPDPZ2i8A+PkPZs9v9RwggGEcAzhajK+DEqMm5SmYWE/hyBzb
hnMQXXRpzcC5Sg+imVtderCmgubJPXfMeRNIZMeXFcGPvNkJvBF4qpY13EL1Izfk
fJ6gQ13gROZY0fjXdp7D1N4Ibs6OHRme28u+OAI2t/apsLpdSsqoeo2O9NhnClrl
79SJ7b7P1k1eUqoBV69E2hODxqeJQ7oISm8++rWtjj3brRN8lDI0wLWyYzbSeIIJ
+7pssQZKV0srxy7EGRT8eexaHnfYN+tbc4RH3cSW2O2TObzZ0zRhDbKA4LsKWycN
8GBnld1TVNHoA2Ud5q76xD92cRt5cGvQ0LTZekK+ZIeCPxzuWzpckjm5gY1wH1FV
IcrRKQRmcjhI4nFJMGlD7Rw2vATEvvo9xcAb9En6uO+sR4SoFc/buIkWx1CDl/b7
JloqdCYfRZAoBOPgLlAOH8D34wbTMZ15qcq56gzRcSIacOyi3wt0NErZywfRAZzw
iYzs+gwKPz3shXD/DLqSiICemsuACHDwcww7ImuFVwZDn/jHM9FZhyKJsbYbzsOD
Q2dJGsLntLPkyfWPvQ1LQrnMbFbMUp7bbCrr2uGxEGdFJ0y6G2XaVLUpjzjOhT3A
fJxSR/6iNZZCAsN/M5cgykDjOjD/U3F2d0mD6YJcUfW5oDM1Sa1kycSxK4lwHGaQ
8t0EZ3sS5p4zxIuQcftsSYNo2xAmmAaJCax5p99/Ryibme7lmMj0l6p2j2T2GbDn
znQOUNo5RT7WEKPpMAmhzzq66MFjmhRt4TWrF3SwPVqPKlsGLHSTXnOQHYGq9Hrh
M2tFGTW+4Uoyp+2JbyKBrvWGJFjGDBhy6erqlbNIGfBg6FYCrUyq85vv4sMopisM
2bNyK30wjAKKBPMF2YaeUjirccOBFA9nC2gCro+zbeC3vci59xR0VNUh9qdCyvjT
Ct86uT1V17LNSKyyFN40x9w01eTfNkRyBncIluaZ2ZbFfqtq8l0JDda1DtNLbAm/
zkvzOrvgL1w7o2viTZv0Sg4K+M0FxYaA2NcHlhah+waPmB7sOEW0x8700+rDU2sE
E2YyAPpYmVkPFRDd6xvBHqeZ5qw1naJvLK1F9cjcbQO//jE8nE1ITs1ShIQpEbgD
QkWROO4X2OLxIHQ345UgGrv2Rt57gwPVTLkEP65EtRu3Y750UdWs+RKeZ3lNXWl/
ZXY1EZRorRaBvu9dIrPPY+PMEa6jIWCv37q1s7ddG9C2nlAZXBtgu9tan50xIpGi
dIXBP9iAPwiDgNUbNLA+mnsm7pAuwtK+7pYUnUjDrDZJhu3gvdzRBOLRONqvl+2q
gmwxpvbFYM6Z8QEheIfFmK4bPpoB1MK0acjXljaqriqjL8O1tK5+Ckj8uBUtxCGz
sLDKvuKYx/6eXONA8WP6m34ayStZdP5+V3/1iCsFFh2S+aFXz6dUyc6G94BUWokz
W4D5oUfxDFoQAkEIIA4tCYR2KmOw2uuru0C4emLhM09sGOFOSja7VhL7XWc58mia
ezJOi5FbRIkDUFwLS5AtJlUMI4u9VOstiB+vR/C/gN6XXmCoVdZJJbF2x/IOPbM2
trq26S1qWH/U/j8hP422zDk+JoYXEnWDC9hXAjU3nsovFB1FlTGombC4p3JJspcx
mMo/PwEZ/3m8CSu0G2WGd+PK0gbxtjdRxTZumvTez7bRh9MZt0EpPJXSKkzNPmkg
HWrlXieryag23zWniRh+Jrg/zXU+s3qTPa0Qc2lsKRGq15nm3+6bWLLHrqjxIZMf
8N/JAxrefDVlmyPafFvdnLYhA/h+CDQMhuD0yvSbIRjZfuW4omskUJwLapus4VbL
7XfZHF8Eb4REE7t3P9ljZFT38zcWBTgy+6ZUs87Q7BVQ+45dH1D7RfMmhtk+kTns
4PTytwnSaz3CuBx4dE/nd7EAwECMRupV/N/vh5siKkFlssfP4NzXqVQ+S9IFQ4Yr
My80+NpSRsmfTJi8hKFf1zPC//CbPRaZjUJ81Fl2CE/arvQ3OLVxpuMB4TPVp+0k
52xRqXV5UYYGEe7K9DxV3JPdloaUOQJ7Ou+VRdr7Fz7hcJSLAsJvVnqqGNpquN0G
fQ5ek8qrkVh6ZrH0RXPyFZfsFALiH2+wScFLfvAnu60bLVnl10rdOVaYuoXTdXeR
VITaR40srYNwTxnLk0Y49Cc1qp/SJSIMe/OOjlwVeXHGzdEYyhJWAl/+Rl4R3rWT
FL0+lkrZIpXEnIlOApVXac/M82oOGM7C8FkAvbED/HO63/CSHrv8+2zgPLUKJ0YL
jZBOv/zOIy2Rf8rHXnUR8/jns/tEY0GkTYdCERrcv915hupCq4C1aLQsEH6qYB0f
shJGKIsBNlCvpQf/6PL3bkznPJEMqt7ys0gTnt/vbrBN+MRxOeC2MYlKijoFgUkl
BOo8Pw+TufbKSoJQ3emRyuXka5nZ7Y5FYAxjSz2dfBYF3K0Ga36w8My9MBITnIIp
oo7qny2F/1r4ZGSlCiw8i2dNsNbjRPLYShEhDtF2sH8u1KHWsbToPNi4S8PTJED4
Yh6Ls/iKCR9ZffuDlzrovMICUmeejQ4WVMLUvS94A9gui5qKcyGIcrpNJ/rmhNZQ
lWu45nNUyXZew7ZNjNUpBVjimycEbUXeDEKFmVScPw5mQsWow988TJV12HMDDjtH
Ixe4GSwWgiZ2PBJrdvf7hcLBK5Mp3Yqcmm/Hegk//010CMrzLZDdEuu4i110mG8O
PkfCK8+pNWM8j8iR9pPKb7HURUfSyGcy1ShvmaC+o8TSEHsR3sHFcEv/DgcDUqtM
NXHiBSiEz7BoX2m0roiKfHb0akLZf4HdMxKuuGECtAO1b46LDAO6JVuJyrqJvrze
+hDomRLxkfLz+OEOEKsc/5lKpU3Mbk7XQ6o36KRE0pDH50spFuxgDXpeiTzYlep/
swrvbEDnVZ23vGafX2VqfjRvdZaItcnQMlT5uoUN7COG8H8W65weAw6HYKGQJSfd
RdNvLiM/rHaZAVQX23vd0EhM6+xGhojvhakWw8453oe86JmYvIjMgeSXkQdwbglV
yYHe4tE3fNF665rNujVPPC8LGCAhEO4XfULgAK6xIiL0LNf2nT03R/CZlIPWzgBN
vJLFdsOz9qLj8kGFk/U7T4aEruzea2QVthzNBl6+zItnkaTGxl61xbYC9yeOPVYl
lBztaS2SrmEwY5FH8OoCgkYdCD+mHduZaB/2HksCN3ZKqkbLA343/Ntu2XdCsO5e
6foi6acikvSIhrX0kX4s/zg5q1fTyuI0esKL1pufdmLVH0d5Da0PjbuqxczwAvka
3/GkkRc1V1mNHrEKrcMdREhcv+lNOWfdmkpUu/yL81V584hBSyzK2gmajd2c1Y4g
SN3Pd+iz4M3BfzcblV9jTguro1eyfOcmWtdvJnnO10PKtdx7bBM02ElH0HgejfJh
F1Go7VizqPotsvuzAs/93k0IeHcVStHQ8/TQY0RuFBJDkCO7SpQhr3wnizyfFzg9
6xt2FtBP9WHXE+xKE88Xq3x41DiV6lF9BeQOXZfOi8gx06wFcOSewY4xwHDpXABw
LtD3+++KlyWjeNpCuzmjrer+fgG6qhilN4fWiRXS0EnaYUSXDXfAUNwDTSmX+iql
UtnpAsHm1inVsKVfwvxUfEqLXWUmXmec4kw+EH5Ni1flYDaN3lz4FS0SYGFiW3SF
rDEKXzyugpFT5oWICLYXiy38VO3JEE1AF+wsMcBwB7U8fIRvf7xpkIrpycBNQl23
ZIyrRX78QQMyUwRJmA8lNSDao4CU33Efa6ohAmMLktulodCTfYnoR/DgXR2Rpu94
xaR3ELBrTvLwNv4O8cO0aekzV4UkT0zu4heBAuuUlUbfsXhhu4M/pZ3XGhvzrJCj
YAbujbDPQHUzNiL0/qsxWkd7xvL4UbCztJaKFcg6A3QA+i897h6+bNZbhV++jeA7
lR5asLA+yaADtC7WuTwP/EEsL33JHxESVkKMCIMkDkhDLFSfKOtFbzoUwOmXQWaY
Vr1tohW9X5OgYTlJscjr/T4CqsYVW1gk7283uSUJA7/c8Lveh4fMsFeZ8tNLeCDf
6r3RSbd/30du+Q5GQjkDuE3bkGDgxDmxJuEaW/c2ZH9hjNZdP0KmA0pVU0cCnAdW
Iznj9dYTkNXYzII6rnWdjweCeNFgGbgFv0CY08LK5E3G2JlypBz1eo4fGTdU1Mgh
Qbn9tC4AM67Gv+jKBPZYpBX2XOHdae26zUA383DFPYK60jHKYxfAQ57/zBcbVm6f
X0jdi6PEoT3uaGMUtCITCMYq72SeIbnIyNHCA4MoO9IiiRn/sMdn+s6SBXlOBqru
PUoGAfDXQLSRkM7Q7UJn3KXu/qFHYNM41vmZT70gekX3MUXVMoX2k8GpImD+k4c3
genaed2YygIokExQRaNofW266eX8HLqUUFpL/rCciKtiqa/RbDgP1xBheyr1OV/e
S96K+X+B+Is2eMX9anRWuZoM1+KMEJEhkbiSqFH/S+rWtL0rUlUkj7QLsS/BwdKO
OLqaGPICAGOaangcdDnMI1vCkZU4MyMOwEr3tkXSpur/X1nOPpAwLFs23p0YiZRk
gnPY6iTATTjQnSEbumtnwzUmxo1UdOFLvqwdogg0rnb7ES7Zxrrfv8klAtQrW3DI
m3WqzwVDxn1l23S23rVPuz4bE9SGkFg/R/r3EbNAkmwFlsqkCeAXt6J3ZDZ/zE7s
PB8/zFEQS6Fu/b8i9jlmL+0uOxT0dZFPftULqsyDwH5vklF8j0BDGT1CMb3tHSxS
8UteqhHLoqPqTp6W7khoPPIRXKPNfMZBaosOrRbQ+z8OytI5KihQwhdAVyIcef88
rS8Ltecp1cPslBCL643l1k4QX6sbzmogfHBQdqXyJQbsmF2V2pDXXu5poWwQuMe9
wEK/zWnISK6Iu3zT2WM/1C2TQ1AIt1cLIYepSXLUMJXy6PU/bb5sMwzdrhbE6i/x
GeFHE/jMyOThc6uePdpmFaY9+sEm5poKWq/5pdr4qDFV+TKDbutSEaY0+f74iKZ8
KzgagB19i0Wq4/MioOyxT74pC869eb2AUyvhuRvqnzQlqmmpxMhcpOpO34K2FwJ2
8Oj2pezSJV07E8pbTDPiylJAoCKUXqFd75AmSS81pELPSS3lZKEZAR8BhL4FEgPH
cmHHScnHdDozV4boWyX6M3EpVnIg25uOSXpv4SwmTwp30e1TuYCNM4Wspw2RNLlk
Z4F2fF/tT7Hf+6+BqSibFs3DnzIPjGNj8KjxctDzMwNzZ5Eqx7aK/s2j9AlR6GFS
Bv/VkijpO+9ysZuw+obO3A4djdZN+cPVACJ1SUzYVYQ8pwQwE6tDtY9mDV55YhjN
vcHhVgKSq+QB45LyfspOf17J9b4fsIpORd8QvwIXfBqAbpfzKR5u/giuKHq+Vyqx
n1L0xyqaySxUXXtFr9uIrkD2sGSfMstvOrR2QMh7vQIdE24yfE+a2Lo9ApolrTHV
kCmtBNFf25aWFRn3w587+3q42vN0Dy49QQgvvr4Z8jzdsIegewrfYFFoz+UcQ2Jj
ep0UvodmhBbtJSjwOS32Eyx5hdzGrrnabQbF1+cH6yXLIlTW8xLrT7CmwR1En5RI
i1KR0whxvCKAHuBFa8IEVAEUBkznmuE8g+KaGvwpHTwM17cRgu3FaGtl3ZNnEY5d
EbeVowc1MUmx+k4L90ha4SuSFdlaniBKkMciBllY8A6hIJChp7B12BB28dT1qPLr
WYxCQHvCU1AxqTmHpHJCh/YWyTcW0jqtgw/xAHzFL/dBmFNdtnDcKU/8+IkeCLX1
kdmNR8qns9HsIdXS1GPXIr8gXnV6tTSBmhdiKN5Lp7zO6b1IrOTx8UzbjYRcf7wF
vVWWWJiCq4eB/3pHpaOsYF8YaY61MoLw6fHBdK5846JYX0WJ+g6hLGa1e4X9TjT5
2wlkM/Vf8fmnbu1LozQsn7YJGpshC7TbYp4rWPROH59/b46fIs7daHcaJVYfwHhA
pBGSmjUvqJR8kH0KxWCvhy6sOIs/iAv8totHICtJP24V+AmcwpErGPTRVTpMCYr5
+HD66ZyfFoyOempTT7GMeggIfEq5ZdIkkwJn9X6GLNvTu3jouUMj6RgLG472jo6D
lhxdbwbLHxUTsrmKb69gySngQv7ggMeTN4pvBE8B6dqqXs10AJ4ic7wyFpdkGKPv
Ch8kb4UnceMPn3IiKYUAD+P90HwBzE1XyujXmoD4vMwReSDEXtxqLFIl4u2qx887
Dh9z8AWgqNnnZHXymEb9ZbWAfkCKNkzZV2UbsJrmPfddHxkATzQnRVX+UWt8oojz
2jtTXl+oDhFq4kxr2J6KLfrTuPkzM9cOUUiPTzU1gsPLmRXd9/nptWGv/ROg8ipe
PhOxh2t87T55D/Uqh/qi1sYUdUYwGAfJ1ZkI/BamhZUQweU262k4fcsewAb7v1Yd
50rNpJWJ5pRn5aW7hgHog2Xq1eI7a0JLMuthuzwv0X3/7zmXcjDopBz18Q+3n/1v
0EJxJyEZJxsh55uaHaXWMR+xbUH3xBK32/QytC6lG1hpNb0eGeLlqVckvJv0blKn
awpFo2YJqJRXSbRbc0plVEZKeP2rCXuWofWjmYy0DX/t3RgbLuYnPrSvZ9rXmbeX
rb8FljHc6Krr28Ok5dEla4ioVVmM50q4sGXguRwj7JWWE9rt1ydPlIGpAwg7ZfnS
dJvVoLm6sYyWzJ7SWgQWJMVgB0RvRPN/kfbYYEXMU0ftCdh/pfmn9L26Hmz3CGwM
BYt2JnOBJ+gkvXEZTrr9Lj4Eq+yOY2j86TlBcZ09pKyhQ1Tf9sTuoi8VUu04xVlB
r+hzop7723ChV7AZ1UjEm/kKe+L4g/CN6qvsuD/ZLgd2fXwRKkavSImj+eY9vw9/
iOPHI1CXC0rSKy+9K6vcSC+DQpgbvsVaSUJrwY+H9TMrWwAFLE503dKREuhDFFp7
DES4Njm3ZtTDxucmTpRYQsMGmT/gKopUJ/GKSgLvoEGdRNZ1B9zfzG9pW94fhXra
OhdjIHfz5g9ZkNjLDXCAms/yRRPAODfHpSDcqzYKYJNkZP0exTV2nLgrMKucMafH
lV6pZlObhqTDXNHkuCOoNLXQsZEh2OpxPhXZP6m51v5a/16+Ib1dIKNYT7pxCnAe
MtDObbVVRzDpL+OwnyBFZyG5eTjLjrA+k4BBiXn3K7Rznb3uIwE/6X3pjA0KZeAE
OCayfY79LiILjoaQbz1IQ2572J+oRLAcYV4Snh3Z6YmmJpbV/4td3E4/zNPqCNDp
EQ87ZOpFV9Nox8tsmY7jFzZayT+EwF+39yXNBAyHGhckZoUQd9+aYbbpliqEMNTM
c40/bsrCLS1Ax++jxJoHwvYW0IZRpIjv7t1KtloGxKFAjU5qnbP/U0H42yiwaPnN
V5ibmVvtXzUEynnsnW+v2kjHmoAqIMEF+/6rl0ufK+tm4quKnwrBWAMuWBoZ7TiP
kIsLbPWo5ARmDFxvwTWOch8YPrO/eU9W/xQfg+iwEOCU/90xaXlqcNSub5g/iC4+
RGctyP4fhn9gaAOkeuuryNWMktGzGVK4y8edbKjjlTsDzQsAAdW6tWaiUQgnr9KR
qaDrL6iONw4cedPx6mfHCDdp3wWrJio5/lOtpXouFQBZ6EVmGREiQB6vjN5k0gnA
2Ft3jp4OflELbrz5Q0JQi4One+sGaqEbH5dibEWkI1BfbvMv7iOIkzW82G3Xtwc4
TQfYlmfb12L6Sm7ipvwYc4oof5kSuHHJuc/YVEf597oEK4OSiWBtjQAw/A0gE9BS
NvILczsqfVqadbcLqOAH0+XTI7KaeggH40aJJNv5FgK3f88rqeMmWiLr+9cT9LUL
BikBj+kV2ZmRKMTIylDSemve9adaLKCTEpyg3nYESBSGOudh9IKEMTVDZBkXHC4O
VH2k1uzVrjGVyZpUKMsonkwBLi14RJdLGdViQATYFmom78ZITLO5vIngWrrgHWyO
nSta2iAmmcdYIXlCSlMzh+1IHQP3odrlrtAcSBf4QGfnS4VVR5ApcHmxZClizafN
A9g9J7U1GD56UQ3g7R9hpTIrpY9i6k+J8xyNQVHkJ2Qa1hcJvs8G0IbvZs/EIytW
O0rXOX1lNYtINhBG6YEFylSwbCfA6hAPlaeVb+lNKxqIZupgvRyS4wLEYuN6t9wO
CB4hh4lrbKyMvTmtk63zOTpEF/Lh8cQn8EOFHwk/T9qwJSzqBpi6jJq5VE3dV5JQ
5Paj5xjVV16M+6ec7eYh8/b5dk8cKJeavRbU71nhwKeEJn8izjKAT1fblOAvakEW
z+FC+1o6jx7XUQ5/eM/Kd41yVKbMjJHso4mI9PW4M+0TjRWp7frIbdGtX3nh57wW
o1ggDTZCSS6SlwkqLiVbv5PF8QBkw517gLulRBXuE04H+qWB+f3o5xBmbukhkCzO
KBtPBX75UmIE2/ZBViQj6UB8fJQLmCd5aFQY95mDWTH1nVsjChWSKCslH22ZxvVB
rOBxg26OPCw9aDF+XT8a4PPCYnJfVdkWyWexVBq+k4MFxdWtUOk2m//0v2DBv2mj
07nDRpMWWQyWppf/tk8B/fx9yjszw33zlJTKy4YI8P2sPr+SfK0dJovFOS2HnM0K
+A10i0p/zCn388wJS93/eYz4rr+65JAyvplYZ9nJVD/2NvWYv1fnfsPe2voeE2Zm
l4YUEEyHHVV3Sh/JsLo0g73owUWoikZGSSR8Er8PhELS8ceTabg7JI/13pRJ3lOd
W1p+3aPWVgmXZ05n4542hUAEhznP+r4QoS+zae12QKZarwniBmI+pOF58SICnuKA
1/ZOudrH21sQbiJUoyh3x1zVbMihGIl2GdHgHxhNtfjrVWAE1EO98KchDqKwgqgJ
YXPpvPlfHfEWMXMZZw1qGlHL3SeQ8Ge6dmsbDybvlvf16tQxYkVKqDJ8kTpJwgnl
hWh2IX8yZ/Fgt0oBXsaJCmjJOmiluuY6aXLn3pJYBrjbifGy4E9iGKlHKChq/4Uc
L9mamJzNma4xnlV+fjbD40PrNOr9H+uLcBcQqju4GIEQVpP6awpxvZ7DoEGwdSb4
bm5onKuXKlTtZ/5OmDTeqWl4v1wD0EdKg1EeVW6spo92OeVPiMO9FGmATzr5gs2U
h3LGhk6ZuN/2Set07JYKAKJwoaYoJEL3S3Js14n+7dHy/9lfIle3DJaDZsQvB9DM
RWresVWrtkFVorn2Rl35j72HKzyrbsMNCw0JYfln2KC0o4T6iPINb3Y6LB99Nmfy
nVKgl8df9GD0ieie2g0ZBMgjlELd96vDdaNjyO29eIYH1n8mXvosmXt9lUqVry8M
f/0Sbt/3u9XvVttwch7pggpBF1Ds9/5rCotxtiRU4o+vjjohIp1jz7RioVYWZd6c
AtbGwE14tl/dJwAK0g7HDG7ljAK3Pcne1BgQi/TvYIMfAN/IFzrQkE4acSjTX4KG
WQbq08wrGjRIRSAUziWM8h55IjlraiLrucTjVPq2PwdvaiLdV+XiC6oPYnj2xWzA
c0gQ/fQrRMsVM59TerjOy7XHYIC8s9cNJMIqg2plZ1ssL9B22+a2BeI2MEV5mMi7
bP5FoexhHuuHYG9pLXPpCcLGvaznwj2uYGC5lZjR/YgGuNI8y/3WRTueLPSEX6T8
h0uChgfTUyaP0MAe3FBntFJDJNxjpiB5MEjQlpiazcN6FKU3+51YJrIJeWsF7lrI
f84YpbafmnkQ7X1ceinT1AH4/ed7mECqAC/VgW73FRdhC55gviMA6VMNhluEcP6l
kt35N+BkErXL4ik+8W49fYTbvE1f4rqca699iNe6CsH6TF3zOISWdrKRl2gLvxRu
7v2SMGAS7sxv7W2vh4u4ZyyZsvEhmdSJs4jkCg5QkHiOhy7oQGUi8AsGlZRHZ8Nx
baaoSJc6ak6J5gyxfX3VXLHg6AkjsYLNEMNBAHXvcSCRVVn+Mjo1aOTi6oqvpNpo
ottzkK6xaJUFrn1gMP7EzctXxPZU76pWy6/PMVaCZgr1SxPRqCTrc0Hj2beNXmzd
shwahQIqs4uapHeOdgcmDA8/yTM1x9quTVrqN1QfNKJ6k98DYZ9L0Dq9a3sJXZfv
HkrQjtQEOgmyd08r96Hz10/IQXDkmIVqqLVFtAHCsaoW98X6tVUmFtf+PqPsjd7E
2Nj5Gr38b7f6Au9Ysxd7m90FvMoVO97aHxWOzlWeyvdFFnPDqq5ZZuf5nkDV3QH0
xPCloWMufLaRhJy0ttLX9uzfC7WnG+8fSkIEeeXCrbWTJJdaimWaGynC34WLV7p3
d4y0Yf4Gy+9t+K4+i48ZsSBLT/dvlTaMOGTe5qC/pqRnzzlcTAdue/fYS2WbsZtS
vu3BJ4NqK3cWLhrANVPRgcGHPQHa7bnFQE1ColBKMPyi4Ldxa71Fat2B9pR6BJO0
wd31FKfwqR66OZAVNIMhhbAJ09S37WGFoA66jEx9VLQZT0BaM5lTEFLsWCtp4mp/
5RdDfOEaBB5u0k3hDcqaSRY8/3EZfcXNp299FvWgl04cOKgfNLHEYDxqem5/z8fJ
thEJIk2dhEVP4Y5tX5ApEy5KBDga46lR02U0wbENe9pIUKNUGSlRj3RbcrjoI7ES
85YLh8EBKsn0cdvpdOoZV0g5oWzrPmBCx8IzU3+9b11gVrVInqmsY/Hfe4H7RrRV
gydM9mqieC3tn0e+N94pXJgD1h6uj75pSIfZGp7Hzk0VXK2vGrAT2atrQRiq4PI0
RYzlxoRjFiQ9+V+y7+svE1jCWMgtPyAT+6LnkxQVeg2mOyfo8PvmTDE36dJP7+Cu
kkq2aH5lpCacuuwAQEjTfrugaKrTVk+CPaSDOF+DtOVtgoKSz6jCtHWjoNPM7rMj
wwLnLQ2BKF7qBdcjWIZv2+cggsXIhLDlBQYnqBGHw1HdnqhO3e8Tdj/DvXUekzyO
RgT5oAVTf4+d8CGdaiL4LInN60AP3hdhkr/ARaoHuUM4rjdosaq7d3axMXg7vtXH
An7UkixGY6hQt6B4LQ4D1mW/G7JEFXAHtrJSDq0HQ/WlJ6Z7cWz5C+fxwFf6n5x6
oea0vow4cC59KLxkjfgW+GKGFF16RKc/652xc/HRI0PKXF0atCDIa80ujAlUOwOY
pGQptDt8mWgRLGJxkfrNxO6lp0mP1HFMpNyE4Fra01ENa1fGDmbXltXuLwWduSzN
BH9tu8sWp+Ah+PJtHMqiRKffWIJ9TwaKhYPcGjkjAhkNtFs+HwbH3ysD3q0ENtPl
X2++QSO4m61AOIBdQg3AByK7uHblZlZKsQNo74YYqtHjtSYrxLsO5UDzscSAMejC
jvDNhW9w7AnUIpSlhsZLcVFjYSgKqKEzsvB/2jW3f+vQaHmvv/F3ZFce6JzJX8U1
FphqsEsDOSUZPiXPdY/JQqSPyw74i22E41Dey0iIZYMEU+FWI4qn5FuvXWFfZV7z
gUp9+JAbHp17dy2y0Nam0GsPDalgpO0trk/VrfGxNdFZWgk+q5QF+nbxuBSz+ZAU
oSG/UASazYEI9amdKLra05ES95E8eS/BqlmJUb+KXtDSQvkDp4azLtr2h4mkG09f
liEqwqr5Wxt7X3dVIK6ozQhn6+NvXPCDcflBrAd5ohIGG2HV/IXRVjvUqKOZwezn
tRak5aIYkAyXBhsQ8HQecxfCOEHgCJPcIhp/9i8zcLPP10gdIU/1XAybVxDmurHS
8HlEJilceVtWe8I8eQOk4Tg4np0H9lun1uA3SId33FZpMPOBsYuzKmTn6MLv72dF
tEBeifBv7A2A/4NvFr8KlxCZ6JoCxUDy45U1LRJf0P/RJ+SFuCD6YiVFepH7qMpX
yJm5neClnbb0ofVvPI3YXYdKgSyxMEFC1e8Jrrjz0eMCdlMPd+gW+XrSoecqUqXR
q1yj9fQhaYaT4KX/Af+xtBJPL6jYGLaEfWQ+WjzRKwQWvQbwY/F9cvbZJKo69xDX
Zaeo/jZdBJ6C6ubam6B/lgkQkhuc7HSlZKVjODu+KQ9Wzft+GiUjdV2+s0+VpGvc
bGY6NUFk8FUnlBjwGRAb+jn/SI7oTYjhic7K1PcX/EQiqkB29GUDia/uvv636DAV
GKMccvrbqOEqpTUbJuwOWTa2kkDqXZyG3qMdO8+3mCCpFItJBGJYyYhHpFAcDpF2
Xb5DeRz+TPsZEuugJbkKzO+76vFh1EihIsVWjeMJ7nzU2LZ9BSTuQAQNAo3G+UOi
2wS4RdKi1buJZuH+KvbnJd3A41uG3bwzvfA4XHNB9xFO/xjCkRirB/TgGyp47tCP
S/y/RZDF2Gp2TC54f4f8t8hg/ex/yU/Ho2Az1gq3nHjb3mEkBSJGRO7VHFw8Grve
PK44YbEvTQOGKEYjKpGpuov5wTT/pK+A9xHLZ4GhiSXAOoiq71OsZgQazT/6nuCF
ZJhBiK9wC/ADXaNTo0Y1QByXrGAQSfEUAz3VC4ebXrq6/m9x/LqdRUi3JtpGP/uV
uYYdNpj++EwqnuE8nGzxu6lfHJDAFwQ/vYnUGYpgM3YqfKg3nR7pyLPvSMKB+2HP
dt5JDdEZYqOyY8AL1DqvcSgyqmmSFSqXLXJPtq3rh6lzC339xWdRtynQu4mhb9qC
JIXgcrGmbqDXXTojecEom4X5SwRPc/RiinbbFrbg/ynNbZLT2gV4AHZSHdmhh/n+
7jMMI3JkJa5cu/BbCg81bKjXIiGPIxzsh0ztlA0xRsZHSLgomPYHy9FQFMRaOLN6
y3bzqddrIqvNjTZITZEUjZ4kU7R9Wy6h56g7aAj1htzEW42Idu//JtwQUGBmey7G
wDF1gB8n25lZ8nnu+ayNMnsCFvTpd2nYC3U9UjjdZpm4G+t5t0POE3PFjj6Q6eVl
D8Hw/OebAwJfeh5xh2zy8lZNwQNq6HHHJ5Fe3zv4H0FoDcP4sBSyuJpSYedp+5eU
SreF99hC7P1h/CdKA+iRNDliBbIcvizT/Xu4/UwKmaOG+UP6ruwBt/efO0yq0lEg
3OUfzc+6LFQktmMwDNhjPFCrbcTdCu59lJ8fMfzkLfdH7O+lfaY4O5KY8rsQ5cuW
utOy3QWeGfOA/CqygKO+1+VcNFEMOVHEBlJWiP0SFBiLL03eazkuSwNIZ0p85beW
xv6hcGGyykS5Cpb/69RM6fA+9rZOruaD02shTWxoaXKCirKVgCy4o7L46E6T39Y1
pixfFSNH6tK3eZYhQyvyErlubP3UJ8cH9HR7qbD4XfW72S/L3vlkhnFLDdbnwF2U
9FsV/Xat4Ril2iQrMOUUz0FjnYybWJJOENHbAF8Z806JYfz3ocrQanOzxLpTKiQG
n4uPyf+Rf2TQDKw67Be6UrsYN2A+idj+7Y0Klq2ZsQ4UpNpQ1uszAoX9d4eKgt7/
hbuXnjkVN04zpFvYUnTOkHj+huS56R/z9m0rN6uSGhqghQMmD6/1KO5ikl4e2f2E
HVcHUDewyEMrOCq3ciEzqGGXxlej9BxrB6/8eKDKCwfYVsqGfx6QEpZ0uYE9Hgc5
5VWQ2h2O3Vt25HrCF7u3pJpa3qUjUMM8hSSLTf+n7V0DAc5kBAen0tEKU/NqrJkb
/o8adGf5QpdT9AMAXc3MskG/GhQ4IzGtXPZD/nQP7I0GW/x9MgKcpB9g5OSPIFAg
LlBLHcurgYQnlWPxvOT5zStgvSICGgxijqnuKNowGaQ7bR0OUEiofyYJOXBN8dqo
S4ocp/6mNngHjiy7mvuDEoE2u1dKXiGzDe8KbyCLE+T+stIOMA5Vo7FjD7eQ47uq
qYke2RGj+9fVR4F0/VFcCzh/mh8mnS7OjxIA0kLn8yZR02G4hbIHA6kXdgpYGOu3
q9v1h1nZJjq9nVzfiKkEi4B0Ugpd+PAD+PGOgau0ePdgKWEzlnM5kZqQDj/cc8F+
TSU3wPr6DuU4vZZ34/NTjbXbY2t/Yn/GJNWp19Lb/nKPJXqiqCls90d9HxzLVlLm
UD1LTe1uqXLttaQIwg3mgHuaC+wIpCNNCq14MfdzYOyY/39wVDOWGY4SkvlapV99
/oWK5qLkgOYQkeTZWFa5RWhV+h7chA08I4L+F1SmEGQ+Ro6KbGoCe/tFUiBrVGMt
8mt90cVq5tJ3tSAS9OMTUjYQAMJ/sTCmq/trmHHt/b1c8g0yCs5DaUrBmWoZZCcX
abgm12lKYd9zJYqG8qLr3G08yzIbY3EMp1knK854NH4kpqXAYGpnFiemI/3DO30c
lu7TIJA+JdI9ghkkWRTr3L/EgjgRokG9pxH7cn4vqtCUIGLK4TBb4m+KbmmTqd2K
8oUvGfyHnzmhBq/l5ajfOtGGfbssSJK+AhxgIxmvfWwOES1F0CNq2O3rDbS0++nz
x4IO7hOQh0Vu+/ejuGNrCW+d3q5lmuM/NILlIV29khdq2bSkabObwKCSmiDHAt4l
oyeXVT4yNsqSCNqigffbuOQq5UVewE7ELyfhfLXdKB7g5JahZqzEKbM0EFZK2L+g
QiPboMbe2pPz9vl9Eq+TcEogUDg5g2F6EQZOJGrTMvzSfeQTXQr318PYRWUjuJQI
74/CZxfqKq9O6EaP3HMZpBQP58yGsi7QPRER5MPH/4k03lwdVhKuS/iNzqs0M2lw
dBGT1FzuPR6HPeSUnmMpkbt3CUh/NK7zAWmiNVS3J3aqZvo/d7nCacNtUe+tzkvW
KQbW04GkXmOE+nwEFSCQO2BEX7vJ9ZOylTZ9HSdddDmjUEtbuZXhFiMx9Op5d+we
LV8qoz7pEpphjXeDe9qfrIf8Z/fzMAiGhVL2OIQyqWXvkynN9KrE85CVoeDQaG49
Wa6vluLxGyc0GNzV3EaVUEwDBSowy6VDZGNhD2Ghn1tsSaBh3hY6BGG9veyeTm0/
S+qigPYnnxShmMMxJZwVf/5O3y4rzDLFwhUdZyWCOMzz5lDMP+MtQTbwDwNVCynU
MJFVKAHHEywpIeep9hXH/gSoU8W7jnGD55d1UQWjy4xUI/65qpHMRhcrc2K82zy0
4EuF7DqiCE8mwe1WjmfpOCo2x/graDR7GoWOun2qmZT94Yxaf5KjsNoHv6x+RJ6j
drdzNPOnO0LccMogGxUFf8VGGhSvG7MpaAs+JNx7ZOtYFwpYnxNj1goaHeZ6Eqcn
vRBa5otkjDU6DOCiwM3mKTPCVawQ7fZX7jITXkOhsnM9ltJKdIu+U/gubNW1AVow
ZJyvjfLSqj03C5vnBJfc/96hNDunjbzdxV5uzm2fxUu2A6FG0L/tS4PWbCQysjVL
iJOJOxAaiGTrzbhAC94OWaT46VpFKyhWLvPLtZ+R/clyKkUhjdye0y8d6+LcQm8J
yvnpxuGkvpSkvHU3BnwLpu7JIem2fbIf+pO8XAqadFgEGBFj2jVGyab9bF4v21V+
SbFADVzoXgulBRZWs8S7MJCkBUHCbrHthK8WLnZoR3f2YhFQm6ZPJs3LDyJ67Zzs
iwDUWEHfnqogi3h8gonB7PTk9GwrWxhpWEHLRXquh7CuyfaRAg4NC75dZAKG3oBk
HLxbeD1SF5vBFfqjsBMolWz+vPR1bU/Sv8GSBlAadHzgcssusYOIjLX2tt5hikG/
p5use5sUwXMDohXbB47DDMu0J4akJwaEwD67eyy2AlExYU5JCGvGU0wJz8p9rKH4
7ZWD+A+rSCg0x2EHS1a2zniDhjDr5YbUmqBz1TSBFADkhgnu+2HpCTYbn1z2EeI1
oTry6vTjvlQ3oC0HKPLRz/8HvwfkIsGsyX0BIrdOYpLXlLHceUS+LT09KojrJ1tg
v8UY2cpNFDtm6Za3Cwt/q6GI4maTmbIOmqvwIeb7fJGqtCiwULBYtZHzltXPpTNc
CraLEIzAYU13uiQvXvnv7k2J+wsrQpAxUgUQpYhNCJdUZgttjf+Cx8LAWdH87Y25
6EsG5w5EnrFmuefbUJuzC91SxG9ejNFs4TrKh41bstzWxJ/Kg2SLjoZPgaOjgC5Y
DFTPqeYf3Tj2oq2RceZaWgqSy7AlOMPBnQmdzyUEr4M1U9+fTWh2qIUVH4N4jZga
YN+/gDZHUGRp2YLB4b1UCdVHghGE5822fr/xf4T+R4WgPP8ttirTFaTzsYaEssmc
xi8OZdN2F8WXd0Kjf87xFmob3PHyhTjjq21uykNb/6jpnQFkI715qBZhpqN2i7Xo
eVT3k+PQqsVISO7OPy3w/5SjM6t21JgJcosOWr8tx12vT15dflqS1PlvjF+YE/WG
bapQfd452yklBagnQwiojDU3w388nDjzXPcttzvjt8K7pzqbhnxfcVxBXCaSytBZ
WOoR+MxDcjjZrVu/X6uyUxOivxtgVhkz/F3xV8h9FfvqmdBUJYY4m2Nh6L5WBy9D
bUvqeFAEiFiQSrYyDo0IVzfJF8e4aOsFvWCp7XG0IlHI2H/RzN6jiIjpAOOJUX5D
LlPGKm3L42ZkcOq8apSZzjJUFLVPnh0rCKRvhPFQIdP018okNhJyerG5U1TM+I5i
+YEN+C1PdsoONmOCJNvoko4ZaUCX9OzJ4l/UJr8IDviGU4yyZQxisHesozXDHL7b
o6Einkf2xJy1dM8Z5SXZdZCOn7X6+aSeHBCLa/K5gBkVsOG/ee9cd0ETxJoYKbZn
bNsOlo3COrEDKB3ynkYag2ThVu17kIdZXsfwsEkCvCeCTvRNSG39vCRbFzVma86Z
MoEWoxG3Dbqsm69AkyhuK9ICwWfN/0s9VMx8Vz2QtFVAMN3qTHRZiYzwNdEk2Obr
R/18xqDVGa93s4nBTm+3iPasQkArynUg3+3wpe48rJfss62xH881xEtrtb3hgq3x
WDw7rGaJ3dMqqH8K6VMr9k/ZRTqaKuNjWjU6Kjc9QAtSKOXSS+2NQOePKcxyr+Zf
vhObYhsOA7VKgSOsHX4YVaW9SNs+Z28GfWALmpLGkvFpcgYynCvWAF+xvi0sma2d
X1UM7Vs0Li3g1gzLkip/q8u/YjnmzKE0cshNQX9XeiPceT0cKp6wDh4TKOJVuMme
3JnCOz9e3NtKVJTz3yV+SWpk/to8j1LNWVGgk2jFE9dT2UPDIqXmb08BRAflVQu0
7v9EkiNOJPdlmlbIx4nlG7p9e+wXymUEZkFm1JsEBbGHgyKEeCuvOz6K2I0gzx2J
Pp+Xojy2bY5soVx9H9xGWyM4knQlkS4YLQaaS/0VOJygUuiG8yg5LrME3YQKJLE8
fzukHRh+3mJ2hWqpYmCPFh2DjXR85u7BrN8MtkpRT0GuiHaiqMf7NUb1t0FY2IZ1
BfJArXDNA3Xmpdtd/wqQSLafsS5KC7PwFNcxxgRG4v6p1fW2ywcWTFVvMrrYNvO1
KJcfYbJv66JDVgkqHUaiRB1lI9boj57KzBn5l7bFgUPoHWygltyqpDgJ7darO5fc
g5uvT4ZwFmEtMz9uv69QKEuleydDlu7UrNuymB+9mAju1lkSqTB61pV0pDK8k1HS
P4wSkanCSdOI79tmIHA56xhd6UcP/k8uFa6d35nPEqc+8oGalBRhzgSpfaB+MBzB
c3aghq28XpzKW26IsGwSAubOdZmkic0mK5MC6JqJOCtbklW8sU3FIJR8XjJB3irc
e0iFARwzazb5He5aLz8Y5I3ddobQRNs/OkTWuE2yEz4azeqWG8ZkMIxp+Fy9M6T6
QhTWE4/V0Pw52bVGT67vc1oXCU5igMxAIUR7yzUfD8ul5eDgqchr8GDm4bsC2B9E
iR6csQ50Wbe19f4oDWSJr/c8Yn/sqp8i+MBVq8vs85cP6XLzOdjMF+RaUWbAlxdz
LvMcoVZYYXMYFdkHTUAeLGmxn2SV+HHaeEH9v67AkkKI5T6Q7khhHUZrGDrwX3gm
u7wGRPC42eaCsjs97fkWRaGc4fVf+ngIqNTCcrI66nRGz7+lXVTCsrWDtUAcH1Fr
kttUo/nRYQTxRqzmIO0Xu1o4+LpXZk4hO2gXR11ZIl/QdLGr1aKe5pBq2deJc4i4
60wrJXv8izFggx0SEszUVRO4fTH18e7GW1PBn0NnLnKnCQ+6fsF27IUH8AU7VyTc
Cb9h8jtQQGB15uh9vaG6jq6z24eT0Q0/bwKkOmWAIOqdHgiGGvvEl0ipYcJ9JtN7
CzGTIhdQFtPAgwuQRwegJyuWHAkl8b0g7VdhJu7wnj8T1krMxzDSwnTIhD28Zn3u
7nXld4OLaey4vTdNCkVNbRrqYGo6+AhWTiDU6OnknBSrBN1EoVcDPSn3psiFeA+g
nOW4gI2Je5fQdrqITFQrmzc5SsGy8W3XvReVLNGt6IEUefT7LjUol3Oq+7DsByT7
SnUUArXUt+Qxb/dVkfYoOmmexOgpulysleQyKinmXR0otHmlIOHZH21vt7TeYLmh
eDtpnLHOmELk+H8TYnW3wZDapAWXbi4P+i67Dcw9ktkhsRRAPa7C/Ll2LF41NVUj
Pii7RiI9eEgQZFrhJ2+Ji8KDGd9pjWwY5OOT3MVwz6NDgF+J/MK4TESD5vWT0gJq
tF+X3v0IeIlnuboU7iQ8qQVnRaIasM0tkb26lHfCzbNU1uSTzOI8CRXfLMQ4Jsuy
ZtWTL0hauhhmdWhDUAIjzpwDMIDbqM5TkAwcl49Fpk13dqPhFVOg8dJ7PJHlLAAx
4vrGZJChs7bXXF0ZuMBJqYrIICUSYVNgZaXiVOLRMhR9lfBbCoJOCZ2HVI7mi1cC
aga0K4Zi2wdXfs52rtWlw5v3YPlpgOQGs8Nie+5wfbvf8FAgv5m38Z6o0yyQgyhv
CbKVZ2+Cu2ZEqOsALhl2jv/+9E1+DVTxDe0y78JZBCOwOh20I+kM7BMk6EdaOy22
k7ZNCvVzLXYT1cALyCJcNRFwz8mMaKksFVvCBt9xTGbL1KHgr0thOGtHpdq6y+u2
NaX4hyPHRfvxG8wcIaJfP6pSGddbeen4/jKuQ3ClQPXRYs3OC4yecDvzNugOQmrf
PYe+nNUNCSWdJCwLG6HONKyTILYOOID//hcVMe0ZrLvmnIIpAWD1jlnROxHD3g+F
PLeSLNaOFjUnhQ659IOENWb0T/CoVqqurQ/NgeuVLFSi6X1vZeNq3yiC1BeyF5VC
13qySumxqUAble91o532CP/3Lzve1Nci460uXsreF4vo1NHRz1Cu2jCEb6WbX4R0
+GWHw7SlvHztmcqYHG1P9avNWlapFVrM504tfTJRoe1rvcBfHjvPrMsxaxA26K0H
PjjnpghBVzJ8VpkEZ5H9RDcJiXYTWTa8z4BzcxU0xfBFHTwDvEjl7QuM3vsiN8m+
0tseEABufyut8ZAkIzHf2NEOOPihpCy1LuDeIEkixpnFZRu6I1OsxrfNphsKBT4Y
6Shln4UclMLdaLbs3AmlrvTuEC4VSBjMzC8T89FP7JwCygGQ2C+WURI6y6Ql4/rA
6+n8Nj1up+B+xd2xOohb01Uf2sCe7C/DnF+JRZHu8gOSckVEaO+O22r0049fUB7g
KrkQFR+vxoslCd52+oepwAbS6SIgoaAbBwILAHnWHGc+9EGLZwQvtA0u7GBKypm1
PpzB8FTMG/cNRgWGhtAEPsa/kPy3JDLL6x/EGbDA7Ar9S0w2CfxEeAeflG2urE0D
DH6FaVsGoGIvcDlj4Y6YMKGhY4btUNPBRnNWPSYd4mx3ghFiPWgMw3ReQDOkr3m8
tpnVilEW5dFI8ySKUYTOQyNbxsE6v6f+UpBjB/c0oCtsBoQ3+bo1vjrZlFNaM67A
QdOapxPUXqXzURRqMi8QJTkoT4FFM92XuuzW2WsnUb/2ksc/dFhPpsK4geLzzTL0
Hqa3RGlivisNgkYIiTWdsMVqm7ca3aP1lDqwz9GGP9u41EvSlLgO8Hx3l0Brz85s
aWTq55lcD2l+Us7IcntdkDXujAESefMXe6zl2B0ErugfaMd3VS9iHixIsWPONb1w
jM+QjklGuQiGC+ajnXD+9Le2KXLZxzEXo8oQ8kNmXN2F3QXEPCW3ei+yWJ1PvBXK
PcNNV6GXtlorPiafXOzXLxihLOaWVbbeSL7v5uy2UljO53FB66IZY/XMFDsYOMw7
owAhEYgOdNbel5IubdShFFxHseArNXaKbsW0yKY/y+YozRuMqrHhWgpTJh4k24FZ
XrM1cQ+s81kQG4uBOdR/o3wHx6fZ4l95hIxb9Lcqt0zTM9DkYNlVhgbUdXSM8QtE
GgObsIC4JF7U8iD39qPPTs82v2t1E/a5snzO2MFlI1inGw6ITMmO1EFx/driMZRB
FWN7XdWf0Y84F1PgfeJeSpJsct6R1CBIqzcsinoc6LPgnpc7BUPFhKe5I8QwMcXa
8gwNqljA8M3LVrlRGZx4Bvc4QrVGEIk3SWhz+Yly8OL/kP32AvN0VK1W5G4kNKH7
SD3UxGB1YUUX1ZgrvXDouWj69rOKf6qTAVyaLga3FIwGAMw2k6QvM5A8OmTHjuow
y13NIaI6mYCg9RLqlLSvkzdP/gyshjDRDBvNW24OGAk33BsbgJTPzvo7JBAAl+fU
GTT5tfIKDcGVQ28DClj1kF/PgOdQRhAaX0sHvAuzgMSY+C2QgltzZ+gLHjDEUs4c
kBH3Uuz2VkebIdSjjJaAHAA/jh1fBP6bXSHI9eRqXk7GJ/CMYqJKr3LZbvN5s943
B8MfYGwH8bwXGEp3Ic1hnmNpI3GuUl0wadEHuoi0Ip5gPYdcF1e8X9i6dANpVYex
cfGVNGSwyq7k8Rdtqltsoh/r1uH/0coeXYrT+YWZn4QRS5LbfeWvuqK6G7RITizZ
Ms4gwLN5QhMfE28U2J8wfl/PCoEbk0Mc6XrjlDzvFmISRsnls0BLThqat6J95AWL
lGPG8RCeGUiG9hV/fKuTL2A4MjuzD9SAm0aPQXjSCv8wDrpyhaKOjJkTVAJHX8OL
s1UC+cVvPYFedScqW4LDfTMvRomD32tFV/wAmJWSi3ab7phUnyxanVt8jyrvDFmZ
ZDIfmLF3su2QSmk4SLmDebVkj3rlZ6Bz1/62C1VZuVTVyH1aMO2QXBidBDq4isHQ
M1kmlh36hamYWEH3xgAqHdn/2LVklLqUEz7no3njnM0KErXgKN2cSM1i6/0ZxVZy
/qrE99vWaVTF63B47t7sFX6sddnvCWeHvb6y/fupWiuo0rT+m47PvQ9jgHzWtW6F
aawoSaOtO7yBywEfwVLD0KZhTyQkXAABzGvNmnH3TdACpnCwyuzvmVWntprv+1Aa
17OeCaLzSxy/q03zzGf/psYijXZwqxbmBDlaQtTmIvHqtmzqX/vlOq3XfCJBxtSk
fYW17/PB+teXIAYW2XG/21t8L3RqqOTb8yif5abzOJp1cAXK+TEbeoIx4fQL6UW+
s8d6lz1ExFyWGQsCm56EFwlnPs7orWcuY6veVyvVqO0OP3+htBUVfCJ8aiV23obQ
1C98a8oKYqvz4zcnx0AfSEMUBoBvQyoQV2SJy8ki4ZdG+jSR8CfG+ucnA3dNNqf6
TEF47cZ5Y3X8UJOHN1DeC7x69RQO20d+woYtGjtopdoI/F2g0zwLv4hU4DIc3FDK
lCq1MUYQ0vJv0XtCaGgncytjanyAL+Jt84WJxTmwHzRetx6AnLoeRSEEqytrp/ir
AsaTPoKUJ46BCQFwaG2aMC3KzW/Gns75QhQKOlGRB0LgfCxqMGPBjK3RVZw7pwwE
FJ0pM2de4QS2+YUFHWMS4f8UKtJoyUoDv2ydI2X2JW3AvAfhn9rJny3dWxND0+lM
iXMgRKeJ7oNJindN6jpY4vXN/i/7kMorce6l+pvsndLD5QmErvudV9h20TDG8zCY
4OsPVlunuaM0/bQ5K6aLcnTXm+sG7cZeygJGy8cepHZe+/fAIB6QIVMYFv7rI3Dd
kt3aEJRsxenaiuhTuq7USISdD/wkV8flprgSHwkBBT0Io/9XzJB6Zox98EQQy+29
wL9pVIC8v+8HExXrtw+fmDTH+BkOMT1cMDe16IVav6HhMC7TWZMgtRIYSl8Z3nJu
/Qe2KBhVczVbCKYQZqMyn/iqIS93dSXi5y+8RpZTleN6Pw1mcKXOkDzVtqtm7V7c
Sk3GX1zEh0LPaG6nc1KLZUYLrf9kRMXAZ5jQ3lZ/AV4gMthYA/QqwDWfW0aALITm
CJBptZFLzv5h+c8szZOXwxmjgyiTU/TTezLDaXgbsf5WV+wR6XU65aHp0mhQePhc
0APUSYKmK9i2L6z8I9LNxPnZZvm3YhKLZ8aXoVulM6kZwyfqyp56bU/AvLVzLhs5
1UcGfzpFK6KPYG7Gh/DVQg3jdihJSklghYce6fZb6vhCEstbIgqFnsdD2bcVNBUJ
jmkNQ045rVv445BXB45Y+4bWcSqBdOGvgz/wapuNpwG4QxOp/FeP0zKIkwRKMKe1
zSyVJlDjhoqCpLlpYAdYB66cljsiAk+2yKjDFpcjmpDIYP2UnNs2e5y7k7CDdazF
39gEtIukQy2t3RvJYShcnHPdyX2yHgH6/+ciQwiwNOcYKgzt27QEsrecWbjz0dzt
NTDeFcxfY7kBW39gFd/j48F0BjA4vYQljU0jIYLGqJIpSAzp7t89Qt3wlCyBFPZv
RVGgwLUzu6qG1C2AMTJPISFWqLM78FiMMASTxPEm5ispUUhDwSb4Wy6qVGzbTOmT
Z3TlfCDrWwrIh6imYTMvpAlniTJFwZQI3D8ZIG/utvURq0Qjs5r87g5GuQJBdPsj
FaLD7fV/tkBuJBgC2oGCgbt5uYApRyQd0YdudGrRjkZ0IGMqAMqs+P2Q62ARz9Qm
td551dAHmqZhqq4ZZlBPMl+WFg4pnE6hJFMocIYo2T8dyK5FE0eJu85v4Gpz9KGR
BsvSzm0u0v33DLtYlOhV050wpPJs2oXwZDcvgFyljhRQheJXVlXvyD6+bR6gg/yK
5CSZauh6nyPpDVAPfnoILL/HYa2xt3WRbyy1qB5Qf/bNwHlXiP63no0sBBJSzCo9
iP5A/4XEMGOvC0wbf41Wa8d3nunhkwbW/VRaZPhQKBhZd38aUILTiYFLehKG4/U5
rBPiqjqtzDPqbRIvvrIclqnyIzc8TGOQ5Ve/f1XvPCmwyEiqXGaMf8QkrVi7h2kl
A0VHPY2X0HQ/ERP2P31g9n7sVPniWDoZHedegfPXV9bPEYfcq220zJrWo9nT7II7
XMWA5nBXFy+chHGgMRK9qGjBqGNnK4K5fefCQywzEQ1FcnZbIMbNWzyeNayRXFBk
D1nULjEYOIUCOmqHvgwDBfDCSOf6g9b1Q+54eeq2ffTZPAfwyG+qdrWjDdW+G8+N
RmRZV1HX4JuMIRISZYGNaJzudhvu+T6NO8yDBRm+8gwv265W+qV6+p708va5gaHv
qsF5TeOhbyZ/uLL6yEwEH8tO1KS7wquDQzAwzu17846VPKFQRFuSvSexdyBZM21U
aNp91EmlLGEmgwFxom84WiZJio/+rZZ+J2R0zpMGZ+Vfc0kp4TwZbrRzPnqyyNQd
oZrhYJktuEcl+NpISSJUwsYnVBbMp/aqJUo/LK/C13WxGx+F784kgJbpIEntdC+n
ss0SXc0Q/ahk1u+BlrgGS0vJwmNhps6dNe9Vj0f5HasYiHJTPlfo5hLMXCzXczlj
FiXzuQXQpLJMmBXM+M3C4qUqnl0V7m7sHiRzx466yhYi0umaB3NU6UtGPPx1qCZp
y9jPbScEzh1gBIoTXPJZ9/EGTFcg//PLHu02EPj81O+fy85YO5LKOnHPxgAo1Xbd
dCYMyl+jl1hwhZAIO8DiNBz5G1aVn1ykVDT0XQlIA8irTmnXXy+7HCF7gs/IiUiB
2vzAfWkgeheDpI4kLR5RfPDpgG6nHYWZkjKQYjDhruk0IUFLVOwaWricmJAWQnD0
SakGFfvmMSNt9b1zdfQPWB/dlhyWU/8sdoFnymx1GnR8KXtkpBp0QIbpeLSHJ/tb
u3hI7lXMyan6Q0WqzcI0O5HJe+/Fco5JIbNqdMdl83oK4fWi3b1YM/ei4VokUTGu
iYDrgzYlWmmf/c0j/0rIEr19m8xCBW2fUP2jEGmBwkXow94O6EUCcnGm0umTrLdk
i2Jxyu+oy6EXBqpHw9zNgw+2rbniN255DmifoGm4gBYeiEGG1sl1ToK3ueOsA+IJ
YeoqGuSW9jFhzpSEvEgd1kITL1y1+SDuFgmPZ/eOPWMGuCAub/53VAIgpHrhUuCl
cIjgZUTpwzLWIuV5Frd02EwPK3WtUMTBGeeEVO6XIyzrAA6XWkQsJnZAQWq5ildl
YctZMvh31nanFuJJjOWeousomcUmERW8oyAADh27sNooxGh71BGuyASO3IvuwY+Z
Mt99Majb2eyCqi6flVvQD4/upgO5T0hb1DISmd50pJK/Xw2BWZMxNkrIni1QnjMW
YqAUjZevH4cqyJFEjl6LbsXCd+KvSaL/rjyY68VlcWGkekWFlmdJpiqQfxiz9L/3
ioEKnghWcjoEaEWLcwPReDaCrYegWqOneP/VGwLM4W3ZCA2O8obCTgBuifkfuBz5
/c6WRaxhM5jMfJDrqW4jfe/rLYRux6cQ+KzyFidDhPswfX1Fm3xz6PKrZQmnckbM
C7twvWvuogfPyFxza1lXlh2jpKt7Hd2Gvzpv+FBLVZ+1i114KQyzUbZ8/nbJIMu/
i8jDLQx6PRdCYgjkzEYqDxPiOlOuC5PjW2ZPTVyVpgl2S5vMRrZQgreWfKvAW7Ku
AiTW3U8UGmL7fq4nA8Uo/Onw8lParxr9xNwQxAh2KuHDenaqsNEO4HYzJurnR3Kz
4Z5plrm8AhB80LQZCIvKHp1U2Mb4ekxyS2glUrCiozyYesQQhI/ayR5bmCXpMYeo
bV0bEe521+JKksgFTBfoTymNOxMGOkAKCPkVyDR3LEB80JlkNFXZ0/6zLhpFuz8y
FoM4pv/GMoGXKNdQoQVwu1CY1uQHeBMqjrMjBnF4I9uaYF04T3j0YH8y/se2dj6L
J2wxAPZd7HOdWtdydw6bmjgCvycR2d+KaTOzay6FUI+RBIg14ScnN38ej6fmsu2A
57BzxOaxkGhjcvDcwLZmWBgPBd9dXQMFoNeEElYVf4PKJ+calat7fVAvoC3aqYwm
xm9mkLrayLLffnvIZG2TINWCxldIALeqCW6RiX3s98WFlbBd/sCFIAQ+KIG2tSHq
RUyTTwhs4FL/jPNvq/EvqZi7HRODyexD92T0QtLDZVEyc4Ged90ZzI3O1/KUUZIi
DN65SzDFCAb3251FcWFny++8fT2NMXFfoL92qESCmE5IUDfo90L3kDOcQiGbCKs+
jy2MTj5+WkSkmatov66DhrinziqUoiS/pSgRIgH8NoQdfaN7JddECRYXyMwlK3Bl
ZMWMABl77dN/IIO1YSZESHZwKaWWsM0EO4hto2Qb+GdOcWowMmS0sDv+A7qUtcFU
YeHS3xzrMvtDBvZ88nKwxc8u4Ng6Df0v8dlOacTL6pYm6duMf+tqT3LDuEHJx5d1
d5+4I9dFYcNwlCUiCOI1sRUQyeMXA98Ej1dcuF6UynKE87kwl46eRq28SItFJ0CP
Ix5yUntvMpXciMzMTud8NQLNhVBNyITWQRIWNKPjgaIMIqEi1gKeottFS1ace+IK
AJ4QlQVzdkKNB1Pv3VG+5/4rh8xWSe1i/jKdrnak0PNPO21aWdOOzBnmw1L9vx5a
n6XHaz/js+/agNqaFyvmrJviwnMRU9882mSpmVtIDaLZaYL5TfZQHM21IzukLSeA
HLn2j3GRzTZPv/eiLFCbydj9MPhiafiFezLpPXMEWAv09IwevOuIP7VxgLIGu3pr
t6+OXZroLSnQNyAc/sSm1uU0lA+f1CG1UuJtO/l9r+t0idHPRKT7/4WFeEnwA0lA
H+Ko/vfvaPbRM7Nd50eNHHkbG74zY3qy4UbFuuvsmW+jfWzEfGXl3yISptBA9MvM
etVPMdGpwXE2U3EapYAfyfDNnqXfLj2y7JQGTgn2KBNvfq0ttNvJLItVxtSskuea
m9p4BVIGxrJNDMJm9Zn3UY/jsokRJ+5lzrS0skWUqULTpBQ/12XK6ZJgEh64tMrv
3AWaVv6pklLEQqkLihg9qNydsXufv5cmDivPb0ALDH029RQkitUktLTAki7DXDPe
luUzU5JF6K11DPd+JQ5oje7zxPBIwnE+/5GzVdfcx2DQ8gRmzfncMOvXD76XhFXL
8OCtEF+cYEXIR+/xZSb7cU50ptvrIpNnEiFNZm4kTbLTYxJZz+wPCKmMOJct9Rao
meyW/m15uHJDoECS7/sB1y1ajXQkOEC8lJjKJNdwcR5CkV42sZGnLOXl2upN8eru
ZkyiQCFgqMK3hnWOdE+5gOxujnUk8xr2803pWOSy+NO/33VS7RklHSS+L7eoctJY
OwBInvsFts7oPTbk8KbbdXGPpx/51U/k6EK6BvX60/IfuRdleTajBaVP033f4PGr
T4W5dsbUrIeuCR7TWzUmBSeXiHJdIZvSWDfR6p62fJkXfLmSUuoDp2Wuwe6wAkmd
uSZIyE2nEmRjfsgzSKN2s6DlAl+BIzxL4Pm9tAYQheVHO8kHhcbsHNevlW29dQq6
aPSIzUifDaiulnOvk4nY3ElS6zAfpiy30QTlSVafEU3nNjNjAPvn2JYjSBqF6kGY
/xZUua53Bi560o8wIzpAPpIoSk2nReI3y9bCZlYFEvd+ddwtKiQfdMQIa5b50XCm
SDTa03hNiLmN6sTDbf5mswJpCEpKlY6EbvXYaVoUAje+nTDBesVEQBwLEN7eSMIb
M9ZJBD1GTWLGuSM8fM+GueZKK+bl0THR4GyaiGCdTh6rwNcZM1tEke9v+Z2Ud0n9
ikCxMZ+f+7Guf+AUveywmIvPije8Ps9NBVBZL1WCdtfiI+jXsZVSLXTKg9jaaNSJ
AndDCsX/XPqOZio846Rsn2a4GYWhnnjjnMdWB19Qa+HDIbGlMxhyilCw/uG9HFPR
tvKUUTY43VrFBLRJD9oJS/JWdppwgDhdqfWvhzYRbloeyOWsMDu2NTkTzMzpYkgh
pWZ2QO3YXDIac76oAuw7HflAcsSl6rSPEJeD0Ma1KGB5DYi+D66jLS7P20YzGeFV
qn72ljVGowyUjYgE2Jp1xgGdWSMcQPfkVVgAkNLB3JcTgWajOC64ls3hNaOxX05u
uqGwt9uDLk9BSLwbn8dcJAJIaAXtOQwKQzM/yxXBQEZd6pJQJ1c9Q68iPtwU9H1l
j8miy062mbV1AHA5oJk0WO/BKRSJSmfcETpdaij4iTm4rTwrhfp4hvHX0pXjkVUK
93jNGWkVIKb3WT+oG7JgQRFFLsEYdc6jUYtqQ1AEohuy/RTq2ICSCbIel+EIaSJJ
8dWf2JXClvxTo9mQWh5Zuz+UYNYNZ1ft9dFZf9D7W1HaSxayRyYehJFbOXSVm/OZ
lD7LRObKrm99qCYJej9YHG2XV+aGG1RjtZVFITzIPVy6n6BSeLtoLSM5ONoxscmE
bJ8Si2IlIQ6iXofP2f7DUJBL7IldHfgR+v+L94blYjJn0K4LfKMecl2b8vjfcxkA
EN6DFuWmyRi+8SjI5wu4EOWvN6DpV1fZmp1xzRWlvHWgTvKm98ZHkus6RTPsgdQD
aeTOjDs5HvKghGnC9wABGbHsUJEr8DD50aS+nJOvHGg6RtzoJIF/+34cI7Op3CJx
rJVJ45qPPYztv00TbUj8ZFZyjOsCw1bBdNds2P92KsHgj6/eVuymNfRIhavTdVsR
MlzeEKYr9ewFbvaEO4Op+QFdGuJGpKKGdDFd7+XaRAAXxavV/7019h9hJIrLlALz
1Kb5S0RGWHak2a/r/k8Tgzp7HJP3q+CNJKwuFvXohDAZOxOkev2ehxuEPCLUm37Q
99mPONdpUnfUDnZ4Nl07okir7LYyXs9649J7TyDJvrnh3Gor/wmw+QZTbKLyNnam
64LVtQztQI8nrO7jvCDE2Kbe12nJAMnDvVy88lymwylChF4aD23CLRdpOdiLXPTP
msGGO9FTfHoQ8db5k2a38BZzC6mgUINF1XCE/k3Yj3keZX5RcW9K2LhHgrwXhDp2
d3hoy/uqIZJpDaYDzu0FihR+XPaRB/9SmJeXJDbDOFWt8l/p3Ajr0zb6S+wM68u/
fa3goVvjKR28a8UZoi19FUAqdO19aHuwqZkHIXr8pb0x+hoH5Oj1YzBkPUVuWwAI
KQjiyyF6Q7ifTRulQ7o+Khd1aT67LIZX+Zx19NuF4fGYjj9NOUvfSYEJl8nq05fA
jjec8xdYNJvPWM8GHA6NYSdcY7fjgUXH4USdnEi05/67ziQBURgpPUPsXvtC3vga
D3O0+bfhD7nADAuJOem2E46g9k3p1IoqKy4kzCeo4XmlRRbQ16dTC3vJQ2xBZLM7
i3k3jd1g5e6iG71mhI+lrHESpE7YBb2oCXW/WiCN++if5f+ZggoV3uw00re1vjxC
hV8EHzOmSNYHp9TWJLpYbs0B4vLaSFKEdC//jBzpO9pxVmkGA/vVZ2huq0hWFCha
7N24ISZZLzcPwUSbRxbjs9lVoQJ14hNsKrhSVHRXCIJ2XN4/4d4XMQw14ylUe6os
40do1rf9L2nV9eOjejsBhRISxvqdiJArfpplB8Qt+bevNjXRdLD5hs3nEB1wP2XY
je3/2cHG2gjk5OMOyepoi4kaIVvrNzehQiIUV7pXeDL0U9fK95hCm0Pc9iDIMmDv
siH3+fDVh20XiCdAm6rfM71C4mUnKTmZpMAIYGnZM9i0PsPqmt3eeiT+Ca/h+NmF
62ba7EAANztOKkSyCaafSVEluLlf8VfTa87dZxhXAt8X1da4ZNtvtOshqu/D6C9P
f/HncX1+Z24blUcMdy/sUe12qBf3nqQlYAEa9A1aAbby7iqiObHfoAZPXsGFd58T
kwr3vV9TCeJCkfaHQBQHp+BkXzoG464a01Jq9faK72yluUaqsP9t6dpGyQyoD7oz
cyxKgW/r6BATOCA17jei/DwWK1QgWKyoxlIWRkcpRpD/E692B22vYRNDDZAWETEn
mm8JkPTlFq/kYsrGJKqIWNhirjbVEmmpe0YzyhVSoYGXfTPQWwbJ56RDFUfV7j43
QtrniJR+qgCs4auT0bewe21MmXmzwa9gL/aquPbBbVqpqfh+0ouL5g16Dcyl/HQ+
s+0uzkv/lia0mL60pGv/LaMtB3+KVwEq7KJAVwoDaBpeq4wGms38MN1/+rqqTu9h
2yItmb+cNWeHhKv5Zq6tie+TSU1nyyZE2+TP9BUOsBSqgGo0kb4fIn/bLdwTAsAE
JAtmRhDGHMzkqfNKTDr1de66mkoyq5KyufZ1uQNChUS8xvwqiiOwibaqVqmDyPWs
AQlg5qJNWFUx2dt2UMMRqXc+RmLpBz6O1QGhULBCXBrDKBQOXC5Zt7pDQHz+xZXP
GZGT2IuYI5P6exFYFlIj1Mr2ygHudlbV6ukq/J4WXGjEI2ZzUOfH1L96JigQZyX1
o/PXH9yNwhehxoInxnAHi10IVBAakZcQd7NhexTasq5q3Be53LtmjG5hXOuwUnb4
eaZdSrbJ7S/1u8tNywVKGMRw415DCM3puW+8Jzx2X1TduCAlqNy3WWowBgYpgD0H
AaKmo8LsK8d4dtgg/Z3GKBiZD3w5urywfnponCAsc8+t5226Jlg+0oHgw25E5Fsb
r/nSckSu9+qxu3aBW/wVdkhjoPdaw2Ab4UM29yIK4v8r6UUF25huoxfCl3FbDjpr
W4Hu1E8rBb/qiKKHc7lcVXribNl9JeYdMAqFSHV6nxEA5OaEHSN078ZyiZoi6U65
/yDxKC7D22L82POwJ2YGJqa43sfko3xCWj1mNNNaSdN9bljI6aYzUPCcLLwkp13y
ddQ1OT9NQCHGoLEFaoRxZ0jmi+xN5+8CZEtS8628NzOvzcKH/DocIJju7gma+wwB
WAkzqlTiVBMY9wsIvYyqlGx3R0jMOhjSgqEWbFIoWrtbelkRm12ISj3BPbbVJkHF
423DAr6KHa2l+624DfXPd+N7K1DfpQu9MVOzsGM+7yAbS08u8s5N/+WyvZdt+9d5
Nm50NMuq3u1nQOywXfi2PTYiuy1FoZXR0zafk3Y9GY+Yp2YW0HDmubZopVn1G5Ns
wJtBqIFiVPhVZGJWZ9puOcL7QiZc7Qx1+ofv5FTXRJbsgKRxpTfnDL0uLbK+OsaU
irys6fz+JXhT2g2q3vlFTesswP2IsTHMc7DFpBdO46o+yHoiqVj+/48IQhNCyYaG
ZTVfnCsysy8lM3ZorkS7eoIWagA1UW6a21ul5u0fiQYL9vw2P9THtkRSumM+3sC0
TP87SbY3N1sF6yVMx3FpdaSHvc153BPl5ggs/BLJeWbhC1olJyvA/feizdHnyL1M
VXj+1Ns/RMha3NOTFWWrc5gAXEDH1G6/aXRA5s0dAUqD0V8G162pf3doLpr9k6Lv
0aE8tHAzlZNJOwVnX3mUQ59CXrm52uOTpw1Et6a+n7VquWa12kA74pkVH8XXExKB
HUDsDVUsJhv3pHCUYi7AGIeiflowxdhxlZEImbUl25RldF+r/SmhYKVyNEy/vAee
JL9iWy7BUhVf/8VXlU/NiYtit9mTzfNJ+T4QaLPYxUYzf1l9EqzEH+tsHh5DyZu8
8U5ZyRiUup3IwoOx/U6AD0pbKnvWakuYZ8nptwPFM9AveToM0MZGWv8f7JnT5Z8F
yw2UaA6giF2sYFMZmPF3PnZt+ZLXc9Psq179KEC/quZlrbOMlVsM4JEsYJmHrWBX
QqhdFwjaaPYjcYyN3Aml5Bj6wTdrRTwR+uBq4zFbSVyx+8jrYMEuqfvB6iEsXXVy
IBxxOi0EfrbeAfjI/HPR8aHWemkwAtC7QArMgrVuz/HP3o/J4GWKh4FwyjLJgL5b
oBfRlE1qI0bAvGXuf7S3WYm50QCWrDzTVRiAotEMlkrFFYns4kgnZiAi6i6CUXSB
Zu+8y2W9dIb8T1Dq/VbWEhkokxzHHrhGth6FPS4AyHWZkCXqHZkciKTDk2bAnPAd
EmujsDcpGEVviacOOqhJ9k4QlxphC3tMnWcdcbxlEk8JbZp97QpjIPiEi1Ck51qS
gNY865k0WQfenbWSkVpY4M8CO0RQqIsPe9+O/MCGpLPQAWPyAUYNGTKuu+K6IXxi
55HWnITBCAzj148LEnK5liY+JdhSCCkAyqvfqd5TlH2uGLGOWo7/fybuUutlTwfs
XT/ncm+W13+DMItXD1RbMspriXdagzfqadKymJ/btaqQkNNIx98WCHRjdYfSVrIT
vTUBofEF1o0WJtNMXI5GAum3cghYHJ+GQw/51zKna134AhfjzMOV0CSM2dDaUGt4
PFjUgzPW/JFTtvbF0mzI+VNvdCjetDi4eaEJ75ux0QFLUak/3yImXrLUixtpGi/d
juJjmxrLl0wn/TQzmHTusfdaLaHelSQeiREVIpcnqMnFEBOH1c8eTkPbJMlpEXVw
FADG+CcM0tU0mzS9P4FlXEi0x2rBm3QDwcjFImPzs8LAwmvF8ae0RK3WyP2M3OvW
xR0guYp/JXZvmACGAmRbhFdo1qwtLNSiKIwJzujqmRVqLcrb1BxZY+k+KTSFOUJ8
lvy5mokdRaRpHd/evE9EtI3GEtvuqyJipN340WuhNDjW9a1whOkyDlUzV0PxQS8J
8Q1DM4y7BvbDcJe0xqeVZRGwezypNuiMz9h3aNTXbug549AeZ0dEy6ZexjETx327
AWqhEMBfs1JM6CoL+uxEDIKQhgFOKBDgQUm42gQ9+2E+Yzi07TU+AJpbWay56Jpb
6HI7txPY1wXuNlGLPNwg4Lwc6wUH5nrkCTJR3WSITj5kCMsor2DHEy3KyCAiTDeO
c3AC1B5LS1+U+2l1V8VYInoV/RY/mPjeXEenfF39YK7r06+gRVajHHuTvdgstzN6
lez21AbLBr6BhMRzQQ/H/7Fk3UcZPML2fr5h1MVPUjmi5rGHR4vgd2rxoR2pqRud
BLlnbOdBLxM1GPU0Ssyc1YAoTniubMeofMrgO0ZTUvxxim/psauEULb6/b///bba
ZPBgmv394j8bGwuvFEnAfdatPnNn3fCr4yJngs5pf6IUPlMGNS3vxTIF9rAM5rLN
MpQ7WzT+BUzmxCBQdAFhxW5WmJWGaoZoVIXPr9Itd73XwtEJfJfjv+jKxsfKziLX
D6neydL3bEUNxFoc9nY1H7GKOjOgsTNbaIfOSdcwl3yfUgZ7yOh+wQw6dLtzdL4c
tiIFxaQbM+bOV2uN4iULM6tejJ9Cwqd6YJiQrOsdzVp9LwfnbTNsBbUfDoAvOR7T
jwRRD2RfdfXEJqknglfK5gRIzvgng3c5cfruPMDDfvfEXdglIwkbAcwbqg1YGvGP
dvdSbaFzQZYpir/XA8aCkWlRG+x+/1KuXnSDi58CRH6YAPgmSUe3//ohbZY7y18Q
BcWwBdfCdaMEdmstM7gzKrLrWG9+v4ZP22JtyhKcfghMwr2WnWNB03L6Kdf6r3WI
MSSZ/e5cD2p2qaO0uQCh3vyQXYwBli2J994jPvHExEnniDIgR2Z/OJPXTBGkIIng
yUwqnFsQAgqSVlBYv1jIstvagh5KlsmXBAhtSOk5F4CWZQixxVenwIfA/0WlYbaj
MBo6qsZM4GXQQDhcD1RuRX3Vb+8k5ygveB0UiLkRBpPC9QyKyNR/P58cj2p3pOsq
Rwju5ouTtEHxeFtuixesO5Hi5up0B8lUB5beO0imPXseYdwFv0HzJuU4E4cdJOwR
dS+IdGHtjGdBFWaiazhO8wpEpPuYw7h/D8xZVIKPUZT36p+Ce2plGsHZWN8eLF9Z
QoX5XZeSMod7n/qO3sVBhiqiWiaCibNRJpC1lptdLwIa+mS5mT+JPeuuQ8tVpW+2
3RzifBG6emyyqVxLpafrvWh3vSqiMoSkxefHYjdC3z5YiYztRGUfBaOtcIYGEjeQ
pRFQsRbPYkS8okqsQFSokHNRPM03Cqe0H+ytddt6vV5OLeJPbCI7/U8SFQN8wyva
WF+87xsImIBi35DyayANfU90JL6Q0Wbo2BlgVfXjG6OAZKxLrzddbXelJDUcgTCL
MjxHvP0be1kmDl2s2GHsmJ2b/zR09feolOiAnTEW2nhexFVcQ/5AdK8Wuctnd4fA
djfnxdATVMkvxb5DyO1y+RPzyevToDgQv9g4ewQfzETCT8iHpO3tt24OdADmtB9a
hIEoDi0Z6dMs6+NdtvpKndeIfPADPuO4t3wi6IOqHBSac85gTzc7lAX4KRdBSPet
PRjndX4uncmTHi6Lh+5OYoVUUkFGM2Hy1mEriEU2sWX0ESQZHmziTrN6oS3gZwO0
52hvt08yfNhteyQ4Gwx6B4TMGRF2G3fc10H2HcyWxTUKWBOFVh8nPrm/C4CFkYY3
ncO1tF+vNOLFpruHZOAX4pFHJ1rYTCxUwlOyPg/9tNNSHrQQnd/egPq3Kt1ohs5/
iIXQLK6P59WHm882Hl6NUc6faEQlxwy2Z1TUAezHpPq9kLhHs0wm5bcHB/se7C8V
oEFfm1DgVbjntU/antIeCRQc8YAeAXyhGKbJjaFBSskA/1iYv2S2jGyUeW02dvle
1wS59IWpeaqPqMrIpfzGFWBjaz90i3BmYI4eMspMN0cGds9VBKfHAfjv8+poT7AB
WHLHcBf9LFb07mIFtlWfiwUDWN4BiE1eXibMJvE4jJD65dKdRZrXXiDaffGf4vZf
0jRB7HkoUfpQnJP3LfcCU3Ws1n9s7pjJJj/dQV2sJ0QkyBNmhKOLdgKYJHmJcWrW
lCEpwSXrKgi2R5HQK+nDJCwtHHRnfl5egB3+1teX3lGOlx6D04r5lCjJIUERqcMJ
ep3JX/iqfQ3Z/vyyIYGrTUkFBtO1qT++H8lXU5ZDDZDTHhnWKZpd0uc9REZ8MZXs
B/7qxcdRtJIfPep9dIlmoc5lqLY0uSzVeKAFKK22OVztaMCAn0xBRu8wJaZsVrKn
pNVuIpvuFGdkVSGA8VTAMqYAl+/2Bz0sIiG/6WoP388YxtwZPsXeZpN7iGlIqOv6
PJbwEldtEez4I3vBYmKljD5rq/z4MpI2bS5TfXy2y5j6Eh/QBQpsMcpq8pyh7FDB
/yubMJV5rXzEDyqTYdsr6Z6/ByOam4vCHvWlgT/BlPwH2SUsf80zL2WO4xKZoscT
wHX7ChcowL6I/2+nMT1j9rggtnvKIGXBZRQeySNp8YdlWZEvuwcmokoCij+FsUix
AHXknBVOr5ITVE6PSsfwjBrEQvUEabqwiH3FU0Cr7Rz2XqvF3TXEVQ44lBOs/alo
RW0WxS6ysVQVhOGCszDpImARoKOV9ggRIB57yb86vNn1/9kVe4sb8feJaR4FRqG5
yA/JVu9LTLjWrlKERJHk+YWmMZHHwbgdCetX0U8DFrcAn9Ahajrxv5pt+mEk25wX
ZrwS0FltI6UH09XqgSZ30PnEn6jX2P4gVGacI/zCrTEq0MaSvy3fdkbcB0WFVi/m
EpeCw6fkle6PfLQ6UgQ9twtlcE6ZcyrKhTjtLG4v2gtsvAv69xARP9cF1w04X6SD
w/oCd8ZOYh6XOjVQxyK0Oadvdnfh86Q+6pYevXCor51u/WCyYJ0w5GH2BbCactUB
jbMkcSwHrhI3dighaLph7fsWWhNJQmvltjewZlWgLW/yDukZCNm1fCakkHJlN9w/
1+3uDgVwh15izx4sLom42ECjPUXtMiHyHBP6Som8yTuAjqL/pbB11xIu0/HBMZpZ
td7fcC9HtHgyfB1YMZIw0W4Q96gnVWUjH++d4T949iBOhUCsa/hXbosHGYxvaNKC
kfbCVb+6j6EkXTAUqf1pzEpZWu8v2IytxQZJl9SVBmIItkXbXHdyS1rRYyRs7p4x
e41QVnns4sng4e11yaTJjU8Z7hHYjW3vX+rqliPIqeTGKUv5erCLw4dgnPkliRxV
2WKzRm2NRmcSHdvbaX4FICIWhI8i9Om0Te+OnHGSmdjaZ0ueUMkxTRo/tQGe6WXw
T6LBt2ZBQH3sXxiESpeMwwozvzi0QkLP1xKaKkv/8CzQLmnW/Mq/GOGFryA7dCkF
ms5u24rK76neu5Dz5LT0zHU91SENK0o50p+2sHc/OoNQEjnvoEH/bWTiQ2+wtfqZ
vTTLV4XC03z0vxBoIWztDoyD755vxcwWQqBx/HWygcJDTfhu1uNaPDSGI46tNnO6
4PrkjmffbFAOjxuhB2U3zfUPAOcdbqVi0abPB1Vx3iT2mC7PWS5noqbvRIJTJCAk
T93ClbqZjOYHVbSb6Sri35ALl5Y+EQnzarU2byjgp8QG1Cy013Bqzk1wHRX6yVJI
4OUto6xG44+Z/MLtwcVMgRxhnETLXfeZYTctB+kepLDq/16mQl6VY24dewz4zL8y
7Im3WE4WxT0AJX9LN1rm1bXyIE/hNeDwV5t9FpYQFX3KPViJ/E9jpp9qZYgoxzL4
9WNH5XPdx0OLLSdsOLJsSf+FvX1h0btE+tTei2oapuhCzgGtTSi3NsdZS2kezken
F+hJLnSRTUopdZ3ZET5tsfPL0e+O2qTe6EJ6F0k5YEV17nN0gyaf+x82lpSLjuDA
PhZ7byUcr5IvpOX2wEE+ujNK+z3jjRlYbsKpf92kKQPVwamEKybkY8nkmw0HXW9Q
B5xdZEeeM6A5PH0+rH1IouTy/EieulzE6WAA66ql6UHiFuzs1V23GaWoyJ5m4eWW
KUJip0MAEdVStl1w5UaZySXUj5Mf48EFNFj6+OLPH0JOS1+cFDEpeE44F/bPsODB
Sy11dulaSpcmrBZysFwETTnMnwiw4nN4emnxQ7nWG19SsNHdwtd3rKhtawjnycAo
zpNVgkjzpsR4CS5ObcFXnQSeCsqKR0coP//WfGQGjM0Uav91yr7WjGvCBOnLvzTn
qwer/Cvz7NRA6n2o/FocnIVDBceow0Loh/H3s0D9C2A3X5wVQSvhVftHX06Reehb
CGDN/Rgo7ycu4JsXhWK7mOXEIELaUQ0F306jaBM+I32pQ/uHcU5p87pO8a810NOj
/JSKREJ8kEhjY6WS1PEjPZImDj8od0217hO7mmyM6CINj3rCx0DXYI8n61YpgDqY
W6WJPBDX+l6xlVDq3ObKlFKwz1m6rsKO9YbAkm/Mr30sc+hJe9eF89N9SfqcezBe
IVeGy4pIIgiwotkzaRWOYx/lGwlHWzuk5X+VRIvgmcSR86PXxGdW6A/6ww4v0IUz
LcA1XJ0h1UA7kvBMv/BmCKNKHULVjI+yjTIK0+FV+46MfA1ckjy16ZZU9kOZcpDs
AFwRPFNqNmcmQc5u6fYsGCcWCCnMSZsUGV/6V4R9Ei51O5v8odAqHiNTHF6nAeuj
/gbnN1M1Jl5PHXmZhvvnM7CAaKoGb7zRviXGeays42qp/W8kRDS/37CTGZKj5+JY
EsfzvaZlanHyo6+I2k2+7gH9xi31blmTBSfmwnrtZrdk8BMgL1sZPJQ+k5XnIeJm
vTsQWRS44fQVJ+9Lzx7HWs0n0/PonNR2NJ8TLtPBfcwpzGKdjk3MUh9p1bH9vlVx
WQHcpDsgqikaFVOaUX7TXbMMkieRujnz98neZxDWHfQnKOOdTEbwowunDcG7j0uG
sL1vEGK6/hsO1A7Y+a5p0iWU5B9FT6QmCVcJYFsifxPhtZ+nMkxDjYO2ockwF+Co
8onYEEEOKgE6DN74hPrMF0KPQcR4UwFBq89WSuGcSa6OHjgUJjm+Djb/B2zH/a9k
t0YfQ2QPcT47K9q2v4RC70O+NYMlji0qTnENB0Lt3qxWZunoIG4s64IZL7ASWqcF
5IRtVUE4fM/MiAm6JOhf1vI+6c0G9aOB9FPELQp0hIDS1+UK50r+aCv2u8V6baZp
UBLbD8D33cF9iFFHdlT0sTIFgw5hk9AQ2IXvdA/krXmX0sBvjqBYeZP1nZwve5jf
F2W6VGopFcs7b78Mxisab92F8l6fAweSHuxDhObZ4zfnjsKyRS/obs5vgmubCY3J
wsmAgVnjv/M6R2HG4CrW0mLfKRl/V1DoL28TXLtKBkRkeVA/pS6Gy0+8fy8sVv4z
nUkvnyJAlVyG/7qGIlvexn+abNejHLxwQ1wzCR9xe4bA+4ECckQa++zvv3cGmVld
E4UZGsckI6pvRAG9ehv1TOx1+CY3upyDkp7XSX3LyVGqIUktg5BKqfIR0Yy/XeoO
L5rG6nG1B2LYEW3NZyvdzV6Elsgn4g1rKH8tbyiRAJYtnQm4upJ5843L4aMwm3h8
ER33qeTHkGLto9UNkpWz07L2jKMeP58YV2ykRXlrfIQPCW3RFAvd/iqvmu9rRoyp
Q6qZCmSaM07Q8fMN2riuizF+b2Ep1YM5r2axkzNBn0X+YHwo7GqXA5I0NgGESbq7
6rfV5UTpKtB+Jt83hNDcXILNJgn4Wu1PI9JhBTliIkpAqepZdwMhsQkKhCj8mrEv
W1d4AXq7zLriyq4BHMdWG5rZdYaNC2oU7f6EiJetdN2ksSNkbWyCy36XjupKdLW7
w00T07JSnbNVUogbVirDpHxDPrZOFsUauj6/UZfqEgmLhdWid0IBDHTNm0raNpca
Z4XwzlPfHO4KgLDJ/BCT8A9vyrHx9AjWaVB7TX7lKLjbnxNNDmpeM9CsFnnnVhkA
LERz06IxMWWxCCHkDCf6Gul794H2ahpacSDSn2vufcRuBvVSSY+jHFwhqoxL0gZU
Oehx+8zNUP4tHSOy/A4+20AL/Bzy9h4qbgzDYEkD09Ka/5ueziXpFtsqsPy3s1Co
HRPCc+rrO+RgRxF1nBzB8XQfiu3gK7VkdpmIifEsAiudqDKBm4H2HT3QBxjJoMj3
xwDMmnmjxADBON5q30d6lpeqXeNp1LdHyktVEExBdwubmXhQ+11Zf4j0Kh/NwL2m
VGeV1gDqqdNtkyQCLdzpRxtPNUJ+9VAw9tHt4aleiNnhGCiORm/URL8kOOa2AttC
5b5Jrp1dJLhAfxZpPtUBYOi8xcx0XoVxrXmwQReumpHY+0nmIXyGSTdlIhr7iXl3
f9CntUpNAdnEyclcwBruDvApfnM1HJ7kSsyUm9WcDjw/p4HjMROXfTIfjnbWJQ3g
zZ3BTA0O72rDvueqI4Vlqll/wMkWbBfXo/QzvOloOnHok6VHZY+2++7HRNA2/Adh
zIYdhyX9qFLH6TNxzvWpKMQD5nBrQmnW2FpnG+lUP5j3jwanS0DTQWN8h6AzOOFt
7inKMx8LtyJVlbHf/sjZiLBwsjCH0PHEm0pljdGYUl3A/1TItxx5GPp9lZqAy2Ac
9/r3KJXpOljTOnEUad9tKPZLJ+zpJZ2TCbLrLzujO7g2E93s5ojUgH+Qmy9t4RN/
vLV0QuOugqSnyOoA6sEbpHdUhZtpffTHqsDiqwCCybayVFWLrnSEpvgXowdKebyq
wq/LfDxMM3y+PnuoiFBSSqJwwAkQkGOxFCdRKuQTMV5pREvZFT+sLk/jk2Un+5gu
KOtNTDoCCiUzs6Aq87Eolljx9NpNa4yeLI07Cxbll4J0RGCDih/HoT+Lg088AVIv
EY9TJP7wBVxQWDck8/TIvRmMbNQsHBhihUDF2h/+bqpzKTtsRkDMNXtDP4EwfE+g
E1sQAjCz92tdm2l6WMKctit0aEPKU5bWWO2gfiFUbKXqVmQKWZoYzl/ESm73GTE5
N/JdIlT77aWHRxIPCFazBR23wnBdOhmqFYstI67riZGpIyQqITxSnJ2lEHBxYGZe
hZdQHmuh6hUNbul56KbW9PqLsUy+Jb7mk1sABBwb3NBNsuFt7g1wJEZIYsN429ak
69sbj9WuyJVMarSRtQ8dSfYcBuIbn+iC8QwsE5FfhXbCEUeY3z70p+wWSvHzeaJz
9MVzNOx22aFitNo7xK5e7KJ2twwgnwQn6Dv9Ak4M3FwCMWmvrOndX/+R2aBpM2Ag
HXWGgxkhR++gtBpjb72y23cze4oW9Zh19z2wCLsdcCqrVsV+x2HSANcHNGjMb3EY
b7ztwQ7AFu3+SW1WCiWn7otP0O/ZZhUz8NK4SZFCskJrhiPNsjefvgRSoO7W/LuF
T5ZQ5avk78ucx8WKdIcbcJXF+m9/ceOf7GCDZnOmWO5O+2PhufKsa6LYuMO+7Xf4
kxXFukOQMXbCpXaqPA+oSYGVEygODwdjY62iOyPzY84qt/17f7ZkISYKSKujR5SY
Nr0T6YEa6+61BcDWxQ0FhW+uX6vqOfCryqr9z1hvKYUJT/PLW7paf0TXItoGpTM0
hKQ2+kvkKOdxaDWLFTGcHovwmSySEmaHpi2gscANdlrjSjUqv/vYQ9LjETg5vFc5
6pF0rg4CsHBSZtC83RyzEQ+g6+tLd2HwGtPpCBnFrAtpgnMbeVhNlzJat9a+hA3A
287IC9OSNus6TrGerwU5/cKHkMkBLLoRLyh8kh7UHUjbqQ3O8NSGau+n3JSCgBe4
RYkcX9X2CC3ZmwAyQKURNR/PGfs+8T9O6RzETIWaGZLlduaeegO+Awiyh/ZAh+ON
qKJ5RQhnvhU70YbPxhmgOAl0VO1UeRHl0pi0kgfBnuabV/L+zKdebwBEkFSAGRdm
2IZwOnSVuY25s9StqbWkAWiB/0mzFCuTcyM655Gr1sbqkyhpql0XrPP4vDrqbFHr
E717f0KLigMkxYce51Hp9YKYvnPGC0CpZnt7lMD+MNK/dyrgkmcZZmi8N0lCRwz1
TDJ1P5gZWhwNtUoX9Ql0v+7YwplAVb6EiEllCEPoKgMj53jws8gktFNcFRKKnDCX
xbC1sR9sHN8fv5URtqvtW7+S0e6SsHuw/CLIX2+imD7vTfaqqSu2BgKmPvmxGiIE
cPsyLOUyUpEW0HaOY10z3tJaqWLlbFhHQBc9XIVkUuOnKk42QOT8F9f95gtmOdLN
GtsPITz9u4cZnfJN3bjRKpYKEvHqN2NHHrDddoTtFnfTg0A/U6/a84m44xbAJXjh
QUB0eoxFp8EwXCInydIk6VtbUovPi8xfAx5CBVo4LxsGNLQ5KJunW/VlCZl0cw77
o+X0lsjy69cwwNvZFwoukvHvdohASfGeiS8dp0nPa3EPjkqHzfZkt43PMNnjzOmN
L30XFZdCdazMAMRzWqPPsciqumyyujLEhGCKE62UN1vCoW59kNT8/xUSQMgJLJH4
HjCoAwNM5HJJ7aEyH5EYZG5sHOz3w+UDfFJf85jMhe+YGKWRrdTETF1OCwco2RaT
aI9wb6yysSsF1nMmTVZOtiJoERUC0ra5x7xz/RX5zDYuOUmHMow8tHfdhaPYZMZa
mbu+8aqYBMv9zk+ZLJbeaRQO4F6eYkxrJhNB0NuS9f6mxU+bIuaMdzxKn7REcu1n
DaECLdrN7pbxYVtEibg1FMezibfjvvX32T7l8X+NxOpg0jtDTUfKCbFvGt83RJco
JhosCPfTC7rMeyEjydVJ3GzLR9urB2UUMje4prXKSuO233YqrOhhansOQ3ITGj/U
QF6ScQnX+JkwI12E+WF9ri+N9jA0p0HlGooAprAgGxBZivsD9uhp7/jqE0+UGkGk
z96nXzsO9FyCmCMKvLztl8srMIx+0C6yYwJHzRSs2G8OBL3Ians+steBb6xCBn+R
chmT8YUbkfJrrlxrwX7IImi4Q3JECa33SyI17hbXFQ0Jj5QGOY9olumO9EoRFdHF
1pq950qEx0GHp1lxC0ooRvrlyjDzh7RvxalMIZmnrLmVYNs4PQBWZ3XSmY26iNCo
FdcJ0PtUv1WHWUKm1TENt3UkC+M8/YGOesa4bG4Vlb+niIRJVf2zdrsd2VBlNg+h
g7D4+L8WKSGKHzPS14y6GHGjUqeV+9hwFq5pB3QNLGOeyEcCW/u88/LRiBwLkp1O
uwO4WVKFhI07GGE/ns1nz2qh6cXPiexZobcQcip55pHidoKd3i4X9HE3Ru02OiSF
v0GYO1qchAYQBQfRyQGuJNQR+/oT7YbTIaTILg5pSFL6U6lH9iLJj6LPgDyaupIg
scj7X4LL3/gIv8L0pQsjtnvgQmzgZFLNvUFE8B8UXtXgux/UECh6cO6fblT5H4uf
mhqkH0rSbcNpbcjkFMJrjHi4QhiUW0Xd4BOhT4McTcRlJ0nNtQhXdO7JWdfUDaXo
CqeX/LWptDv7kChgyipXdV6zYBzbPJjoi65pDMYL59FXO9B4qLV86hyO0pPdrCoQ
jEUWgXbSEoeX6kXbKD4VKX97zcadOkn8QkEbdwwFvV702rDCHCP1j5j+iJi7m3t7
XvpNegod7DxB6k5Wu7+CTMviElLdRp0O+eDcUJpmAsRtU66kjoML1qiqnq9BKJiA
2myU7FrYLr4S9OoADnbDkJG09zt3uups84NfMCbHSW0TMcPE1v4kZV6jnt+yZXpY
E1FnsAKIognVRqQ7nQe6KrEK7b5Rz+oe2Xi4ox9icBuPXeUSJU2YQ5g6v5pfhtzr
zGkkvFJ5imbsXbAvIf96VPJfe78s+2w17F6NYUBfCdeLtAJzmweMGbd1i8NLvCzr
vw4/4nxcnSdACT0OsUcteytNMcMO5WlO9/kVi2gVXc50l4eb3tNyd8BTl4C6uL/b
vOwPfGq8/MnZ+2kWi63MdX4Ei+evuvRfJ76Zliw7iytknMF60L+ZrpByLZnTvKAL
owCWDwttLfZHO6sSfxofwfdzRU/TFacwGLXXYVmP+sGhPboc0H8jEdMhTZtYWabT
ZLfh9eqOkIwkBgiIz1kW5inTY8R4jn3ltwMOwsXYemgXegVpimxpgjNSgicwiCJR
rFsmijhxOfjJDNOzQ0RjZusxdYH7+8weIqI+wq5HjHyx4eoR+v4CzakmieYgbR0j
CFcif6Yc3kcG/KaMKvsneqbzlO3JtsTHgEdpsG8l7SeRRKQrmXCz5IcOPTsDe/mL
/Nz53em/b3JKfuy+KKm9tKj/Lzpx0CPRWn98mUsKi3SvjGhsjVOiJQkd/ZHF6Yak
iE+n3MKrwcQCuXfS7D+jpnJnkt9UpZkuBahMpO++n83lh/ZT5ne0TEah44us71EE
BgZ+aKRGaBEwLMBHOfTHMZwvyD/N6+7gvtxBE6r0tNahqhjIizCf/kjytAny5yzV
XpVWfG46p0ByHFqYp9eX3AhHWuZxHbYFkKFBgon92LUY+eRxL4L3N9pKVpX5mAmL
sBV0mxLo//VdachLtOrhq07lYaIXmE6UD8wCHW2J2b9ZWJHc1pAmrC7CZx4/bCRR
ZdHvxhzwNUIGxXH1HSmFeBwYQ8k6/JY1ptuz4rjMWeg1BZeVqQ4d/K47h/nuR5gr
bRMRavjHx4/GLdAyZPIBuHwLsmwrRVYzq0dyFqOhIaIP/opMv89bgGJgIgV0NE99
RrwDlkkbWn6SDU4wEI5BKARdN5duglzYxoiIR5wOXMhIXD6fokF8vLMcj0bO0Ppj
399z6m2hKYl0RGpQNK2ASBx8d2j3PYKD7A2OVTAV3pmQxPoDVgmB6APbcDakvT6f
UnFwmlG5/iql+MwgAzXZsFBjquh/Dgk/kOBrjIcInWtJ/EH8URKGCz8rUJ7M10u3
P2U4VAZkvMy1+byUvHtIx9L1O2v2onv++kTC1Uqo9KMB9w9g+Mnn/eTgNNMS0bjS
JjbkkSlRhPotKfZw0mVp0sQO3t7dfZWnM6x6R0qhvucOA4F81jMdZoIym/PmxyEU
NQKI2GcqdUOK3FsDteFNOLXpW2n0BM4qmltrPKdmozSL5ZMaPOQSqlMfi4vukWOI
nQNHBczmbm7p0u2BP4gBC1pVSqlKilcJ5GL3WdM23WKWZycj9vaVfOqTmLnuHnZ4
VROIzAz0M6enCcT/vEq7d6RURc/MYjt638ynX1hub3kU+nqcOQoZomGaMRPAAw7t
tnzD/npMMIBN08lT8QL+QLzTK20ha0ZTkz8AEBFW8m0PTIBAPzib4xibBwPTUFd8
3l3WpASk2Dgt8EfPZftNSg7g2vfHhgBFgdofdVlXOV++v+eiLPst81LyEFmo1DrM
oMpN+REOUbXkelcd5H5BSFFAshGmjL9edqOS7BqHVL4BEhhUMH4AydI9yJ3oQbNI
M73UKUpR7kmCH8wE+H9RkHohy0cCvlK5BxZopN3xOY3BVy3PzFXlqK+4nzNl8oQB
K9udpRmw7MO6Ex3/C9+8cHxuCKXcVS7TwmUcOFvKV2emfH1u8X5VeQiCS68tgLcB
fJ0EqH2GyH/Bern921GT5EtrD2n9jjr61w1OdbnaCm9e3Rwj8rQs0tYrK4XenYyK
qrUxtfhmjLVh/4q55OX9QsBzeOd7qTwZyTI964eJcmXdR6x/wrkExr4YPTfGBhrE
bP+b5GmPWJhqTxfjyxaEyVDZN+nphljduM9gwzw3Ns1K2BbGS1b/Bwe7dYT87m6o
u6UGSg+MmK2Fg9zIXBMAPS5WpIhHBy35AMeibFznsZVFjRu30HUZSuRWibiU84Ve
v5c0gtwI3Vuo/E7IuSLShbDxdwM+tH3T8hgdu3mj0/RCnJe/fGIN41J8OBaLRwhk
D7Yoi8Ui9NV73v8gYg9+kZfIDQGG9NGwSxHiv4TtM8X64YXjY8YGcdszxfxwGqnR
kAy6eyPACsjde3ihJOXOu+/C8bcNzZPYHz98KxZXNzDlzhANujhw3MgSX7PoaoEl
AljprBgv/E3Jliv6Q3BtVZ0t86NEDaM901n3GxZJcgTmg1Lo7cEdDsq95AhF0OoU
OtAEOwL1JAxA78GUtajCr94uXxE9LBQ6V9R2QbcNxxNriZgRNB0nh/7E6mEmWjII
akPKadFSObez56ryMnvr+nrFRyWKbLVICGkUqriilm2C+z4YWNEHfpB4tO3Qtvdh
tyYRp2k16gqWIOf2Abp5hchGcZjb7yPorXob0OMAXj4qG5h0KPsO/ACkXaPDImsm
SyHPuQSyNC81oR1XH16GW9tnjAgHJZussN2q4tbEUXNel/iYrrCl2uvabqDlyZjE
msAvdNRd6BLCi+MjWt6HYU6ONJ2TAMcgqccqnYvBkdp04fVgzK7ziPdXzk8dpKRe
yPGdIAhLsvKQ5ahH0R0Re2xnTx03oqaZ3rQVoTI/hoOHCoThOQHXnW4XYOq+tk53
u+B3oxKDi4kQ/yu3/AzFyDNcqzhXrdD8w9sJL3tRoSQdZ/P7yEmc9AJjzusl96ag
ClJ2sm0+0xYTJbyr7HqmY81xxiM1ps9nMEF0vN8HpQCesy585MazN7GgefqEDXKr
2f5Gjr+LQ3Gna5G0pIBwBsMhkH43QGF3A+6ogradFBLMdh29QVxF+pH0JJNrCdPb
lm5uuifK9ZnxE+enl3nSANZB8NoVHEwQPmG+MHtCuROGQMM0a9eX+Szy2hxjhqLE
2vU75lG/P4n+6Aei7MHp767xJdjLhAfm6eKVeaEDZIbFxmuCxseZxf9iIqbmOitG
3hZbbr0xpqnXYb7vnsNMVPaswSTE8b+eBSjVR9lutPLnBhWvXCE5/lUgcMCCNhMh
3+aBgDeu6ljnIuHquCOvYMRhfZ1jsjIKn6ifhQcXbqTcNn4ISsjcfKmJY9ULpolN
pE/FfbpUVojrechRw9Czco5T4lw5ymi+rHmuGAvVKqsl7reIrLiumaVtD7kbU6NG
fyajcrBX8eFcpjJ5H8clfFmjC41G6yJLYWvzcUMbehIpUzs25LQv1UvAHS3T6BQ9
zk1Si+sbN9ZA4RFAOOSNHmmkGdxB61LPt8TRzPlvBr0Zei/Sa4hmomv6+eiQbCVW
c3tkUH2fwJ+KGXYlAHHMUKIBy1VfPSK31jKb4Zu6d/ZcuBs55zpJO6zC1Dil/PDg
KermdGRATjyL1B85O/QcHf6g84lQpAfJmxkMR9DErRAOlGhOGBsFL+414uJMFr1C
LgGkC1n3Yo8VOpo09x1vGw0jwzrbCr5mhK50t5FP0FamfWwYf4UKibGYBBdR3bX/
aCpib6JFw3Zd3kW23Lzab0QR1EacOluSmLC+8OElgnLuntIZk8NI3ugMfXlxrfUd
xnPnjceF1GLYCJ6I2n3XFEHVrWAODp9unlUNXwNIIXA0jgDQ+BXXRkw84ZXlzkmU
vdgymDRNoVZoiUptZmahvSWxxAIs/ouPJpE0be4wCMd1PI2gV6hYlNQBlPg14DRJ
WjeWEKZgyuDUfH434YabHkDkv2qhEj7XBKh3ZD1m512eTMdQogiOc9mAxfJex0qP
kpvEYflfP5DlkKy1Jxm2Z+RBu300bLTHtRHHj7uzMxGzpxcqMSjmSAl848qgqI3o
cSnjdADAsdQK9+T7sMHFgafysSQf969+EwMsR46GBQwknQnE1XKoz9PUi8K8AI+r
MJwgRQkRmZxzINkkD1Ih0po/0boamLRVJLDb7KxUhDr+BAu6FFQjHWUhWkaUoigL
RtcppR62cceNvBTRVcioRqXNzDbCvuRB+hHoa8XxHdhCOl8PyOQX7MUY3Owmz9oX
VMCPkc4yjN7kPxaGqaGuux8tJBuUXdQ5G4p1dNIptnS23wzyNeAA+baQmgQyTz/A
EFF68cos04sLeaSfD0YpBkKgb5GH5db0TQRzNeGJfqqTAOoUiWSxBl68sD/Om2xd
g5r8VvoHrUOrrByonrBQ2QsadaO8r5d449xLW9/QvOz+CUF3CCfZQJY3L+gF3yRw
ojKSmCIM/nsLj8Dx2aTkbEUlWD/ZjhlTOdHgMUJrfzBQB7IYVgf+zUX1yehT/lZP
b9vGOS4OXTQV9RkEyIF1W6Ag+XAY4LtcikkrfPZSalzB5uUMTugPBxhzMe8YAb9v
+CMIdl2DQF64wtuPvIiC4ktV2Zk0XMS5XWiNweyozIS2vttdVy+lypjABgnGBXBu
gSm0lU3ruNYfTqtjwUhpREI8c/i83KqSNlbNjhl/Oxt0bfMhUbDcGmExKv/bzPnt
zEkx+YQrONZAPStL0v5r+HDE1s62Fz5uY/pDhKWNeOqJGdsi/g7MZ7jmA4aDroOH
d0ZYv+y8ZBz76TDR0hkd5+kn4qPTjkrklyRZPJuenjqk7exklb5xyDTKjdPiDCxl
C32BgWXAeK+YD6V7chk3TuiEhBb+k/0s1YqzbXJzGMt6Qta+HpPvkB54i6P2+Q+Z
//rbOqe/Z1bCup2VgUBxu+QSgk1g/Tdolyeh4c3lJm6IPu9Yl1jWjvMspxFNE3Dk
CkljwzAxrO1nooJDz+jeNpmejC8ndeRegpnWUmmZS0aklsaJp1ifEATKksFcqczV
ulNfTEoQlrWvrRik7r7UFDdI3Ek3LxTz3RSlBeZ66X098gnhybn+1oZWqXhHWREc
HhgduOrfz1WkPoUbFTt8aWsHjAf8BV4OLV1KoOjPxyuo0WOy15s0lPmkP2ZlQu0z
W0NcS4Rtd1HjE4aNLe4ti4MT6iMe7MVxIOCUUPCYadKRj7J3rVIfdGOO7X05Y1b6
Cimi18bViej+i5D5wIGm1AXP7CcLhOpC7XjPPbSbJdXO5drUca4pdS4+jbRoVmGN
cpKf0wr5NWVk0HhMU+bPmyWC/OZqALsjFA2aCbX2GAttjt1LNZTeXQS0mCrCZtf4
icqk36japfR5f2QQV84JISMViZWi6TPtHMTCS5eU21VZt39FiAxaRsiF9Ln9uEW4
y4ASMvYL1tXIQs3qp2izT/nNnd+4jEixkJ+ofJZAIh0WisbCHKX16vKCTDqCtCc1
SdAanZdVtfNg7T4JAueC1Tn99kxWEkvTmN+o6cQu+kBK2lWhDRv5pd91I8a4ar/F
04OB4kQTK/996Y+7GdoFYbhx0SXt0jUbeA7ZdQ9siq35X4wJtOdFULYwmAorcl+b
5tiIH5OtJPArm/txS6vmwfKrO5FuRDLoo/T/9IV6AE3PS8FtzuWyqDBWfnRZCDb7
qPIfaNDuE4gNBdiqUoDYvyLDFBwhfLpoikn5G0IIhBw9D9wshM16NUmkyX4gEmJb
iICDxwsmRi30i+1RMzL1e/d0bdDgLKAqn3gFtq+kRwE7nZR5qndSNeRYyDH78KaL
eeX4Mas7fWWmtKCIQlcfVoXa8wv6VWJgWdg7OI6DTb7Owg3IOpcVC5v3gLjUa/6F
Q7Hw4m+jcLdqTlxc4T9aG08gRysV/HPn+a6n+4uzjNJ/Z881iDFuVgBfrhVO6gZY
O/72zkcwi0e4UDqdRBiqGkzXpbV72oZnas2JIXONnDzCH9ld2gQuaTOXIEoBtFh2
4Jya04xXpTkJ9fjeNcu49je/8rqgFEEEr4SZ5lJifdeq9plV5E1WoxLOTTqk/jPF
9byS9q+ujS6AHvg1hhGXwCSHFsRpGec7iV6Yj2E25zodxxFcJcTj5gnWWIEibHPV
ZqHc8ZyWxorersa+gXJzS4NYj+81EkuP30lb5F4B1oFyWwnvs2NvA6mYmJ77Z/XN
o1X5MqeSnF6XTZC34hxq75n5OocemcBZh6/lzF7XZepnabU9AWmQ0CRZhArdvn4m
2kxS6/BW/uPzm5J4sgcxeOEkCI5PHh+EbqE4dmiaXhoStm2+46R6pBiZo+M/lLjy
t2tNPNHIMZCWQyjyS2MEpCXLxZxAbH3tWf21vDqMzyuavfQNPxd8Y2QoOiYqGwdG
i0R7x3oA2UK9pjhdhKaFW/9FTkCFwQUhzWIJP7CyULq+pgXLgd6OsfNKapJtE3qb
7Nymr3V2UFcGLHAGtwrGUBj7UcCCAWvCoZ6wJ/c7vuUB3RDF+FlBD0yyyTfT8IBL
OVE7UQJ1aIqohL9JGNtsOzx4QGGmk1MKJYSBtJbGUGUlXxFgX/NWkj2Nz//tAvCd
0LHd4OK+eWKXza/3jP/mByFmZVPVm3cg/My/+/GD7hE3OzOC1xnvhoIhs+FQJI2U
TAIwF+JVXlkIWt1XhTC1/MK0v66CUwyVqT93/5QXio7JIIbnV/26j3RKoiLY/8Yr
lqXbXfCz0JohuttZr/0vw65SQfy4ogaLTawiMfuequ6DtzGTe7OCyC6fUXzyXAs0
EQvQVEkYFQDb41foKijTjQxxe/c7vPegiufLOXz+og/CLoaEp4AnxDqiXB0wgWwB
Mr7rXzy1/OSAGiNaib6ZT7vOOFZRICSZJmsPp0G4DxrQugl8p7g31gZHB1Ck69tZ
wEwDNKKSlyRmQ5YbuP3js5PFZv+OVAsG9pto7FIXqk6SaXWDY0JWQ3W+O9SmePjJ
xWHOFKhONW2GEolK4mfP6bnH53VDCOLdShx7UCMYa1XMvZZknMK59e9M9LyJFduA
MK4xtRYFDJ7Bb22RY0S8OgONig8qyohhogJtCMSSpl1cV2LafZOx9PRV4c5MdsXI
4nSwqb7Oyre6D7D0myFzqs+O8O0WdgtXZX3212OEioYD2UH5juwOGHzx4NuY5tqq
liXAjMQRoEpXIqz+3pqZdB7W/sixjn6wZgbjV74/k1dlLOHt4LtguX4iOelijr8m
9c/Q6wklNS4mtfFlJzA2BkQuGqIirr2n6soqvZ4dJPVsPwyKd9z5NumBOKFQah+X
e6JRHEoRC5Dwe2hbBZb7JhWvQSZpfzLc1DHeR3c4PfABIgPPF1RGABNK6QEFo26N
VgCLMUSRnj+toJN2SZvEPa5UjfZgmSx4JLP8t1YytgsDbXlQUqwbEsKz8g5y9fES
L9ZM4SWVbcKpb/BL8VkY0Vry0fZOEcwYEiSkQOyOhVRQV4w//ej/CyyrT2RPtNsF
x/iyWwCK7M+4+P51uXJ3mdDlIyqXuzjLjRR7ie98AOIQ9UWbhLPdFq4fYibdycWG
8HAhlPvXbule9HKxfjwtqhgoW9jjZ8AqQ8GLFhgkL2biJY1vxW1NoQn9e8B3Zu+B
jwR1P70wPTUqjSB+uPASPQkOY4qXjw+rf07+l3qm+h2PkH1Lyb68iSCvYtvRBxIw
qLmrojpMyIRtpZHx+aaSnC5REtoQwluljw92bGomQzbv0EmBbcJxP6MMtdeHRusX
7q8DRGILsav78Z3zBM+8rMr4Rl0mmMtJwee7MOeyKalYySs28jsD5IdpE4ulWr0i
3FeYzZn/87Xlm9g7xiMtYs2NOV8eURg0319gAlVrDFcMJqXIhEewcXmEmWq1mB40
P90TJOmj8efoxOYkxRimpx+F+nvr+ji8T4trXuiabs5gzlZs1mLBaDJWK0XCl3sf
gCvU+UkSdf6y1Ob3hAjCPaPYer/LE/+0tMrpGdhR3F4B+l6U50dkLVfvdn9S77h2
iAutl2sTh1leZaHhYbhjs6ucNIcoSTFCR4eZ5khcYGnWJOmkOtIxM82jZep3Cjep
tnq46bc7r46tibV7lDEsl3Kas5WttYeKpFH9rPCTVrjy2XgqRN9qst3qdg3sbHqX
x6OtvGsLc6zGhBJhAmuy9BFAHsnnifAnbQfTGSqEA6wR5LwZ/rRNr3a0zlg3hPK2
HU3LP2aQ3PYcF/fK72Pb7epgQzHGQIitIW4lBKZiB813SnqAgUqTVzJhJs95064w
ZeZE5uP38X2ZSBjsL84mMIllX0mZ4Rs1/MgfAzS78ul6QPcmkrxv5NsMTj0bbRRa
7SsJmDZzbNq3e8VQ9Cj24Eqzq2Ei1lXeSLj3nUSBKt7SPCWzMj8sbdQg4xx8Xkgq
GdmGuYYD+Q5j6Jtq16kmsfFBH2uJuya5lfat8iZpdjMXplw342irGeAUwHJYb8C1
`protect END_PROTECTED
