`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pI+OogkBP/Wg8lrGI5/haKKafhXY7SDQUKCgsCaaf4HRqBo4rQ40UX07YFlnRhcy
BfXy03+n4c3yOCEao3DGMhaufXqLgkfUbTgPxZiCmwlU+4ArbWXPgBnumrfe99hb
Wnv2CamsV8b9C2VbZfYZWZ4SVpcQUzovS1Pj07D4oSm6DaTh8tAf65ymxIqs6Wk2
9fEC5wza0nryUdRMBYaLomi3p5PsiUPtey4bsW7pNDSFxKa/j3K5W7rZVGyWlxL9
6DkFuadTL5+cDvT1AF2ydNSbXOHez7p9hX0y/fKErXCQZ7m93hGvWR5Dy22Gu7R8
8twMUvzGscSNxQ8rjc60dKGHt/waMtWQt6bwXypw2icURHdP64Yvf9gtOAsG7ej4
FJnPtYw2u6RAICvoiqix4FISDpAZKb18GWme5I9kZA1jyvetKZcTYnO0hEOenKh7
1wNZ0LP88AgqDS59MKXmF0Ts9jp+wvnN5hnyIWl+L4nCo5C4dIzfxcFj0D6zAgFQ
MY8msN/Y0iGh1IGR/nh7SYIpHNqrS6xxzZ3afQL0ArBUzNtouP/E8dngxDl0bv+J
FWRzzUjYQri0aTIeo+txWRvvQQRuqdYp4nShzAm7+HSRsbK4rOTNCesL0UfZr7Di
EQoAQ9/VylTR5v7EOH1amBnnCtHdQ8+0XSot8D9yUPdlo6DHdNFEAE1aeogq64CQ
XpQgVeLm/wbXWhUhnGCxzcCUblSIxCL/bwbAArNpRs6QT95s0qbmPqkqTU/dIfeq
x+KoXv9wkNHtSLwRtFmgFfBVdUsKuEuuQiYHQbZvW9FHCgG1tFfNionbGgoUuhuS
tB398fe1ZW7Qpzc75/pNKb4migF/oA/awlXbjiD5ymaP911n5YCXFuNs/3SIFATg
ZWPu/Oq/aEeuXbiacj20RNZ0aJNH80TzyBXkA32Ykfq56DSflnSZ4HahoVqhWVOH
FfDZu3u29XM/NWXB4EDB/kGNka2q+VdKkwtsIse+KbgKGDJNd3I1KPy/nuTwO1jp
WBs8fKxWsM7v74Cv0oPyUpJWLKBgSzZK6j39K/w/g1uUTsqY4qWOcajoPQUicZ86
K+FvQAZccZX6x+WZ6hfM6SEW4SkaByZM5Xyh8Xo3mZ8payas0huEm/GKbbEQ9aNU
qoJjhAPjTH8qkjnSaPgsvSpH/aPSRosX6vVi6dlqHsTu3Oe1ZZ1Woi8tR25pphy2
9axjP0a7JsOpd9DeJZaqQ6vO6jRbTzbaZeBy6gkCPWCbkQWIWIWFG0glDPdL+FVE
YJ2E79U+QCYXIn9AQz2COSdEwppSMvt0F7Ki3uG8/68dtfcyNd+ruvxJg5EdTzzr
gbmfyQh4fmTHllGxXO5ixCXnCyxqfymsgoDXPrUZM/p/bF0Ojt1RX1Ku3mjQF3xs
4ljNLsj74EmdIvflV/cGqRRKHKskrUwsO2nhsAWxPlWq6AAgDkq5YFbYBXcaCNjj
uYMIhonSmE3QOdVfRlnq+DkeRaB5tVJNZM2xrsqoIFFAAs2wTensgZ0E6GBZwTWk
3tQP8NAvw6NlKfk2PNgWQ5rfflffeFzd0nJGihpXRgPL7kG4775fgyOXbWf7/gSk
HdUvUg7QaWy9NzfSnLCwkw1InK1O1o33txvbRmRD284YGFTNrdNnNISGViTgTvaJ
hviW1jJpTsxsXUjoTFuxk9hCebK31opbVKBckDcIRB28SVLUhMo3buRnyTVFcTj8
yoMq/n+Yki4o8F3xXz1kBlmpOz6Ja+iMvl5SC4gro3BEiQ3MoPLgZTyDsRCX+MmV
RwZxq0CC9jg6F0RCfAlcraOo49OzVhKFESfXyIvThxDn0huXU9sgYFZzqhuLAwX+
47vMCWa6cPo6tLjAzKlQmSaqjGaalq5O3aPyGANHarHAzuEZXmQQawT/3jN/y/hW
JMs1uKOfuN/CBj9GlxT74UW60EGAu+9RPPLLTZQAovyKhxRWWq8zpXHXL4yDnasK
oBu1oduqX+bBzwwP8lwlG4l3egCY4ACiAa+1prvvsidnpFuGBVtGHD6XPN+slBxK
X0Ff+b18OnF7baDDQdPsb2JfXDv3boruQqghprgIRqf2Y+i8bn6oajzCs0kX7qv7
99atuixsXeSUqLr67hABWs9+YblhXBzMzfG3BppG8LSOqIcjBZA3y7KT/W2QV3cq
`protect END_PROTECTED
