`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XglJ3qdQQnUn8PX+oYiNMRzP9mxe/QBCXfuTd9y4X/efjk3GBXD9H42WZwuTVDd
ozsQNQckGQ7EL3nhkSTe76VUbLT2r0ouwQG56uk5Bef6HqEL1RbWAYRxP9ROT75s
nqIZDnz2G9A3fz26C45I5FwUxWwli0hgQeF77ypjapjirb/g0yPJVnpI+wYZcFCk
VFAw5LTG3hvjMkY7FAG+2Yhoy0CLxLPYJsRMoG7aVYTYOpBJ0kkMCex/WlsGlCMV
KMlRLjJ3Qbr+47yoDe4CK0h/CA1o/whmf7rGlsdQBdc79DBzPhpu5/VDGunM2uqw
6tMJRFeA1Z+RUVvE4aopObWmpxCSlU1JoFN41QYC85WXfoHtPIM9+BhIe2O6PvId
`protect END_PROTECTED
