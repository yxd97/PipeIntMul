`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
awUDDdFnNxkp9UJscD2Trr/O37QvB2ASdMep4iutEIra82hJLr3tFfjK/mI80581
CM47OwDJl3nY0nNnLomdaKPEhdCnu6HSH+LQ9nOf9olLpCqd8LoslkSfHHFK7keI
Z7ApgOjV+sX5IEewXYfFfP6CjSV/rO927BlSmobZBQGimYVMtMfvLxnmnb+HokQP
py/iVdOeNzzpNAMRl7mBBjO9X0B4sP05y8uAKw0Z1ifi2EsdnBZDt1VA7bKXm2rB
2QHWXnurylrgE9L+d+Nn62xQt1tNfuUZx9Jr+KeEHEUhQql6dTKJ2jHnid59Hp1b
ffKrnsB7FX98zjC12B7Esw==
`protect END_PROTECTED
