`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64PVKqJSllzG4/Kpm4pgdwhB7I7gM3RC+QZ3u9qHRDYtKgst8EjUzRI6i7f+lMti
dWJ0GQ15VzCLVHQgqqY7wOf5sdsnXqJ470XeXm+ofzHiSajtrv7l+4C7BoVp8ydw
Awt6AT6PS9yaTgnV4wd1l3uldoi9nBAix/Z9OtpDjQmIxq+7v2HOm1Ed/kLgB3uP
9bf6uXaSu0H+V8gitkI6eMlrCFoUDbq0sR2SxQOL1uAhfEvwp/ZK2PT7vSbDgyoj
sXA5aS/vPpcWYqzEr/3jnf7fokTsgt8AIW8aPp9onHEQQ0RkaEmFOK75BL57oMnL
OELMFS4/lOx3wouCxAE/QwQldPEbEVIntCdxxp9XcEFLgvZhSQr6xT26aOfCHGij
69T5dIM+MqqH88d7UiUJmQ==
`protect END_PROTECTED
