`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vsPYQ8MDDlDx+mtxWzZDoGzLse9UXbPnR+oBbqbRq0f3gTUzac7gvpy5Br2UBxsc
xeGnDd6Osqq0DwnmR+snOgRJ+KgEova7xvoF1zyIsBF5hSmCD5ongpfLcxXnAQOT
Fnf9Hy/dXvzbDIctmy7QVW+mxNEgmEzYs9RkGyZNFiMCy1bKJB42tee/DC7De2Ku
yfjV+frvv6MSj5G+eScV9nXi2dsdgEqqUdWJpyucjfQ81SKmJGLYaGQoqukffR/d
nDgwqMpxrD1mIxl0OJFql9nl06NTdPx94p06DaWSO304XqRyHHbuYsXRb0oz2I9z
Xtw6wuuYQDj2vzaldwdNrQ==
`protect END_PROTECTED
