`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQ0N7SmbRSHFe7gcwQjN9u39SQOb6UMUynrMbxKxblWd9iGkdG5bXdqONlVUh+1K
qWpdBg6SxyV7suQlxbs3j2ECW0puCvw6imA58Vax8juidAdO7mxl1Ok9wHvUMxjD
I88uHhJ2OLPXnQ6xm9MxbgU802L0YWUM9H1t5EheE5mDMfyjgJ3SwzTeikbFCDA9
4E07LOC290ldmVO4ix/EdgThDrRfscUqn03KUOoElxGJTe8TvY7KIMa3PgQZmGPp
VuCozSyXNnR7+r7PtZxthQ4GmFh5JSPluCO6q9lbBdYoVyUAYZ6JLElE4eqA33Mp
tIBgUDy6++u7Yn21/2Fp0EoyFY0WbpWvj7g/kv5Pqv/k3sF/TwApxgjVs9k7442V
j84sC5N/s6+sBJRanBQ2Ou27tZ4QfrBancLdPy9C8sav7kd3CqD0Ci30LH7R4lwQ
xhtAHD7UnQ/uPiRN/5j+XWLRJbtIy3cmK/YNf0xdPppzUO5S8P2ftfJSRICM8bQH
mlDQgbC9ZvqjjUI7f7ereebsPxujwU3E6/tox0K3T25Ux1OnjDyoNLJl/oeWCRBZ
Ub06OI4PqsXVLEpgLAX052sBZ5JxvKr/APYscHPT6enLjFEzIozOF/gILol7p+B+
cmNd1maNrUX8+iB7uAE4jVLLgXBbHNfBd5kfYI4NaryYwj/9D0m+Q2/+KS0dXKC4
6B7YfnyvWC8fn4dkMtEUCLtc4RYON2uGAG9Ejw4/OyhLIqJ0v68GgL1SvfMr6+eQ
icTyQZFwLaQiSBf+NaIagaHv07Urg7sWYzaS1Z5VWInkO55eTU6K+deNfPB6eGln
zRzxWL1Ht0makqn3RLMaBGe7Y6zmZ1M89L3Fxe3IaUp1OdZfCDaUL5IWKx5Snk5G
ghNHjXTQzD2ALbcRlYTY8NGnPf/gzIrM0rnUswsG3Wwgwt2buROSSiaDm5efi7J7
X4IbsqaWaKyf7+GvysRfalxMOfKmf3DlENmLo+z2Gn1og77qBvANdOHTKoYN78IB
vVIBkwBg0MK2yDyYlqQ8UALsPZFX5pWfEcjqQkAyN+lYHnmo6Ezd7SwsBBc1EU7j
4Qo8TXLqzCGLkYmjnQN7Lsbe9ArAE1cgQhXciv0i8h0AO7T0740DBySbCyY/hH3E
lvGN41PSlE0tGCOWJuM84HNrDO7AhuhlVnFa//JCxC8EYkfh7b4GcqAYI8RNkDzb
KhDvmcsOSJNz6kykixel36KlnSnvqCE5ZeO5GyKsvsaI4Xk6yTU9YvV5dugajL39
toLCJ/XmzwMkqzwvJUy5i0KIYd3YgQOXMjtJJ4em+Lp3wXC0EUEJxG5AtUjENOxn
na8plHRJn6W0qdsjQavmgFJh6GH0UpF9WMvQmj8jMMNP9EdFlal3Jc0qTGrgThG2
W+1v2v7483a1q681XroXiSOYoqHrG4O0Z/76xg9flO2ab4Vr17mzrKx7yjjQoXsF
T9zMHhB98pLAawOUSLDINmRqWj4Dw5cHap9k7pIkwpRv4XbLJ3JMw59twYGLGr4Z
MDQWjS/xnsGsLHrHTggCKdBgtTs8DX74nM2DHk9a6KMqlaHgbdSoeXzHfX1ZvogA
WU0uUhxhYJpg8PWpDODpgLhzibLhI1Sum4x5Ck+a94N/rxZ12767GCBsczvuHDnR
DaSuMQk135YcJJSqW4EjjC43DWcJs4HUDPIHHTOhdB3P94bmftuCwuZroHSkwT0c
285/eDEqejK6T+JpYB9IrR65Xha22kbFs7J7r3FWiCwMgTgC05Wo8RjETQUQOVNG
u3RvRyG17qBh2bKz8czEmQKvL+NsYZ3eO0SgWt5O90/6qtmMg3IJI0vQ1xULq1X8
nAORBRdE62jRe4qM4yt1wrjT4Zs+HCAWSJi09xF4uFgrxGdAFV+fIL3TbaBQy91R
A1su3NcYpfCP1aiJDrRAEkNBIw3kmqf0l4LmhO1M5MRgQWrt05IfU1mxrvVQfPYT
aKVrXwjnnp9x61EaRYbVDlA0FisOCvhuQ1onQODM10HwTBgquq2o5Xgs3LdGZ/F9
OvkJOAQpkCWv2DuMf7c4iaoQvuaGlP6YmaBzLQ/cy12camwUb+PGdizDQsnsHwXI
bl+Qwa4EcRfM7c1/L4NrNyT5nQw0xJm+f4/odhyNot3btdURU3ZR0zlesjEigrLi
pbs53cZspILmC/DMyV0aSJb8rJjST393GRYmv9u6+DpGFzTySfZ6k8jvg/17zqoQ
Pnuv4gkOQa1T7chSZFnmy+DyfzLRJaN/nON3VVKZWRRPTsv7RSl7Tfo/W2ZNsoip
1Fb56Kw77udj1u/eQN1fisMYUHggLov7T7QGgnp6o68eLnnf9RpUbppd4CzTsh9D
Yqy0Tckal/eqH8yoVEqoN0dzgqW2yf/PndGglhc7IgSWLtD2BTnJNXr+9yUVCwKf
47K1s33sxeuubJJUQUaoUD90lWO5XTwcf+J4XhcguwniC/ohipiyXyqZtQYd6TXH
/4kQO5r936W2a2fKGzX+089qAO6aXdvWoa+eRws1v5Ks8o5INiopDqAtJ5XaYyTt
qO6N8/L2Bw2GhcRbBr0B2FxnKiSSWo/mrYQwrn4M2jq72sM1LstBaA68e2iBbQ8u
vVGXmmRZ/eMugBEEnfXc3E3iaf2ckxWGmr5sP39hyUmywSXZrDJCK7z7Lvs4EiI6
Zn1pu4jYj8lQsfZCDrXIkgxCD897VSd+9iV2rJ42gmUnS3w3TTIyT6tVptIIxiTy
Nwh0mfO2vGtkhpKk/UJMrGLElfddBMlUi85HeJG3/AlzZdCP9RDKyVBJ2tBTcpnI
lVIpCDzTzMf1aA76FCPTlPIWOwcAUt5m9CUHnJIsRnyG7caQO8R7VguCCTAZvOwU
eUF/P63pnKPdu3ZhgH5JfV+mOwBn9EGF9QiL9LjqAuY4fgsDvZjQKlaMKUq6KhPP
0br3LTIx3PKXX3nFJrhQxyoRItlwsacNGCPVeWoIQDLMhRHQswpY4fAq6Gt9UswR
VkMi+xcc0TCkY9mkKtQOQhwfjFI50RKj+8/0y8usiXnSiQOadj9NeOugkp8nR0s6
CGke/hc7BkkmVGNzpa4XphPF0SZ+LWImX9m3Idv1sXdl5RD5h0RDoH2E4+rqAA8c
zIKkSuIBtkEYt43eUFgvcH7laElEQFmqSKdtXmxNKoYVA0EzYJJoDESJouhueIPL
EmWICVublLYCtSNkj+6qyrMCtiDIO/FpxmPTbqgPDoZ9Dt5Z+1TISRSYlFn2a9Sx
bbeD/0RivzKw5XXS5w2WbguYUmxC8iacEgo1JV4v0BMlNC7yCUju18wH8v4A5aAr
DdCih/xaJ+Q5O/3CHnIHxGMkY7ngPaNE1A1ZRQjyjUT3U3I7PQrGZDtiMmZSY91N
wuIjChc++QgqCWegsuTW+ah0z+PEOGoEANk9CHw1KOPBsdkNNEwBH45rl6x2OxPw
gfr2JlOa8ptIWbzXXnbT4durXaba+QpB8sJ+/tgWIo3+4h4mPy+nyUXGOI4VvjnH
x7dvY88hxFYsA2kjxwODbznfar4M58slUlkB+rbNttjtpGkzPqO+Y07kiteQ6yVa
aUJCQDb46yypAw+8ey5MUAmfKz37+60j3esUBCUyKjcYKLF+H6Up0ZKbNkgyr3l9
QesNp07vYCWdepuSlp5Ninyo3O2Uq6C0OxRhG9TM62pvSkZnupnEe+4rwvKRafT3
zJMtcG7pVRd3M5NESe0L42FtnN/rN+r53B5znQxj47khUngYqcg7WFNOeabpZZbH
Amez3f/yEqiF4PZHhbYZM6yBNFXVjB+P03ckpu4f3m9FzsBGxSALYoxxrlaD/g3o
kQTUh5tFxVOkBHuXk90LQYyUWdDMMi/PAHeMgYgorhN8vohZ7Be0hxOKAn5v0D0b
zV61rR4x7QOt/mH/Y1nGxuU7seWrPsjz2HEH+H5smYKDJDeEJAEt1ktVGaxTLjWZ
dB0Qec2o2wGJgEGj+Tia+ic/WmfwBX+RFvtKIu0Iv+cI3RUNfCk0JO2rzMziUPck
ksizfc5NM0Vs6nJ4bI2aEb5Y5iN3GdUavviDNFRMXeWie9C5yjWMiLp2/yn7C3SK
f4dlBk6yI2oMju7EbsSv6dZXF+fjVo1RGqlpMThA5rhipsWAhsDvwUHXfovsFVfT
cTMyX5xL/oa7xCvJX16h18ZUob7kAOkPVrfuUV/bcwIMt3xFl3ZV/bxIB3hmx1Bj
CNJ7vgVmxMSXhNilSMtFot+lxZdJ0LLYV3qgxYV8ZF8+ZOLNVzpl9lNpxCV5e+8J
uzbQHnWJ9xp6mPLFoDSTiCHW6qBo+I/w8pntCJrfTqS8xbzYwhkqY4lyEldx3R+R
w0bLY9WhvQjqv3M1Y8bkhv7L3Ys50JMCfwm2SQX/of3vgYBrtqCg/H7Sg7Q1++Uj
iI/SZEheIzKf05eAR8dMFTEy9xvWDSjWEZgS4okrggjtnd7vIB4p0OLK+lTIoKKb
tceozJ8wgkr18pHGSFH19ywUJWjC26QJ5U2LLK9Qou7eRvfyB7w4cCgdmkyYpbl5
UAw98Km8ghUrbUkDe+QGE3n4i0dTh9gSaMqBbZgTs54xEYHcEF+fQJI3w6r2/2qK
nnfjt+Dl5/ntgRlvYaRwu2EBV8CCAiw6PDNRu+ch8XQYSKG94swyY0RBs7y8iEDW
E3OaJen9J8tqg6c1M41SIMyqWhLDMcxgvJrc5M68P0FFgq+i7xsgZA9cpR3wyjrC
2Q/70Nbia+j16kE36Wxc/l0NB++mFkuYEIKx9fN3DlITOG92iDsAmZGs6am3cb7R
kJtF36CbWWJiBdXEJqr8xFsJ2ymQavSfoCRP/96Zff8o73Y02V2/yNQSBIJ19twA
wPLlxsJpAUFrOeWQh+MeBdh1HO90+1WPa/8mCLFx9nCGS9tNYjL+4Vt45UZOj6LO
xLMSQ0lsMaMRWuXSWSfMt34nqOuw3F4hzC5xGTj0DMosUNjve7DrKoAVwXxI8Van
PrNi0lMAxKgrml2dFyF8pcm0qK2zWEJDPSw0jStdENoo+CX8b+J/TmZu0swWgfB5
MigKdaXGiWdEVrHJWiGlde3Dn/iVYsYmAPAIerWHcV9J4AZf4KfCakXkTPH86niP
xBGDIpZ42Gw20kvAZ46ILuF9Eo0oc9XVvT55EjX3/N2lhYsJsP9nwt+l8R4RsFl0
AHmJE3C2M8kyTqqBESw9dcHBdTv0wxq2lHMxJXK2LC7KVUQy3pziMyJjNYuNVEs6
ZhwOnRAZ23wSLkDWjjNvUws0J95mec4Eiy/xPYQLefb7sCuwGhY+21223Nl6JjEn
LEGOy0Y1VrYgiLv6ScPpSokTtYRG4WiWpJJjliiv39LdQycNlxW3Z/A+t+aAvKJa
pccHdBlMfvQSTCKGmUj3g7qJ5kdk/H4AzoaSAEMeJdtMXOAnGb46acdAwZOTq/ep
dPbfM276AOkoAsAX4cbfOgU1o4TJFLtpe2rrWof1GtCbv/1ZhY7KkdPt4o/sGQ0W
Rdwxa1D3As7Y1a5AcugCyobpQsr0SrpwlPTj0ZJtyQzESk897Iyuy5X1DqboaR64
+Gn1Z7ulPphkLDsn81JoNRT9+HGrvsnY0OtHPoQY9wersZuv+DrPndanuaj/Bllj
P32DNUuDqMwbvx20BAafuHTbrT4UdlQhZVlDFT3B5CbVKG8Wpux1Y1saLsLiDAon
n7B59ggvLYWeFdZoy07UCsFn5dLeQaABa9YS9FJkEZufrFt0g7KMF3HvIyKCe57o
Mv2csW1NS5/sXwFAtUGOAZZQdd2lO1ZuSDZrIbJ+4/CWRtNO+cYIlQ6YxU0yCZ23
ad85eRcOvH/sSm8/CJJzCdNVv7b/TmXitac784fp8ta3sdU4h6of6upRe9qudu/v
z59sJqbBpu8KJ2tH/r2tqeLr30hYmcwwfn0IoJ0zvT5kR0z0zG/jJWt3jZ6c5AiN
U/Xll6mfCrEKhh+pNC/bu3t3jOhj6l3rSZpBPXFsior5nF7F1fNLV7Ffw3GtRaAS
NFoitjbALZ+rnAZL0X2YzyMkiqHyyaFinPhLn0dAOjrAnYRS7HUCyGg7P+Rb+uis
E5E3Tefr0N8J/MhTBPzAgOHn/qR8VoAjKyptKWMgZpR8p+Z4vTuF6ugMQwMgPgE5
TtYi5cg2FQ1S43u2ugsX+lW8RoG9X8x8xQiH33dK62SsJvmWL2I9FZrDhT76buI5
hqjIO9IQUFFG6UdWUjcEjBHGLaDoSEDHq5f3zjrep2T+MGCiHwOzSD8u8Ucx9K39
eMN9JyVI3ARPuHK4SnDyh6YIMtMZhfm4nHaE7pynEJSKhcMI27rLldVOI4AaZRXJ
VW7L71ObyUHVDjUf6N0p2X7+r1/qlP4eVIjY21HB1IopnnAyZ18y5fe2Ct5vp9DZ
BdnxmLsiFQRFl/lb8B712IXqaFPc8Gq5MTDA/cuWmabg8Yjt7helVL/uDcGNyliA
z6TjfXgioqXSacYFuLFDDBPcDI2mV3Ofq5/ayWq4lUxCRvDF5U3DWMk70DgiUsDw
czfN7NXa+BvCd8hV0Qyf4Hj0dSjPC5bc/1QEUQ+uYW3trYolpoDyZeMLWOEIXJdB
fIpThu6Dv+S3fRGgb6nuo5eTtIrkg0m+spqKX6k2R6a8gMxKndBLzhlIWgfT/yGB
57/TJyKguaiMo5ZnNPTK05Da8H6/Hok/ObeFtWQQO94Xxki34Y+AE1LMT8wj+jao
wcnJOlbXAnjM31bgzX1z0/hx5QKkiQrpADpEJ68Beg3NPmUItoPoWwMgZLKHADUE
0L3TxhcHfppqX+gRZvaaEzQHYIpr/KG8882oONyCiU5jR0smeKWoVt/ICz+XdEZx
agf1y6M7zitWyFWPg/aGctEdvUcrQ6kYCQcQNc6pp9L2gdgexOuFWd2XhKoPNMeW
EsyMcpB4clWqhFNOTsi+MfV4dJlpaq4pP0WHuYnwb6GRi2eJwOwBglUjFhxQNDoc
JVK+MSF0DJ9XtdcFYUE+3VcJvi2IYp+/19T3EZaqzpwzM/eAiNz3d4gw0tPDxg/p
ls2GtfFasNY+O2PkwJxXUwEu07RnAiCvhH8JjB7GZciLsoGPOEvY6ySEeLU6N0gB
UFMjk4g4lg8P9jDqDPjp4Fb7X4/gCYFsKrjzflOXKbaitNJyFmdjCiIQj03q9Yb7
sb9Gm647VPkQJe0R/S34402y4SCUX6fMzoH6dStN/8+vu3TtIEWZpjkbIDkux7z7
KUsoXLrThLzDpR/k4LaZlcC3Q0ueYNLpKTHdvzuvaRlFk3YHz0Abf8WSXccWIJsT
iDZBDXcA8vFkH70N3Xr3pebk8kZcD6BADccUbklp12Bh63UvQHFyxvY6cATnz0Kc
QPas7qP526dTcJaY2gypFIKhw/07SGFzYOefNtOkuk332kuH1B1ED9iZOz/sfCFQ
lL56mTXuLnr4+Xg90lCDX8D1f21PaiW5rhHTruA/smTmvka1KSWm5FYMtQtiTMmr
TLMdgo0lzYR862+bPZiowdxGiU560amrjyxJuGGMl4YrVLYdxxUeTRYmgabWgebv
avRtrSyJqAwxifF+v9Owe6Pkbmk0CVF+5gbS00pPtqsLOLyOlB0Uw0JkyblYEcRY
bCSQYE7MSQaQrqPh6N7HfT41XAwoLsxWwsWjAc1XmLc2dbrfFEw6exmeEB29MnXt
1ROnkmPjBprlKqEOf+nP4k4+PuprzXI93hSX7TcV491zTW1S3CbIn+kZONXX+Kfx
eET1uuEfx8X3/h9AJkTNsMKU8pzIvoj1fVLWM6Ne2V1VXwiYBFI7sSM/spbXOCW7
2bAQasUYnKi3f2G0Ch64OuN7gQphzrirAxO3hHTo41imevGr+Nk7+5oXF0Mq4BYk
UZVRnlH4s7UMiNJ/RefFriuvR47CpC/8o13Ci0PmLJLGkGex35XevY3YrQbY1L6G
4rCwE6KFjn9Eh84Acxx4/M5yRdGKPByw3xi/nWm+/OjDbAspXdYkKja84p4cAjaz
+XoSSHbaWVqlJ98p4YUEGNDQ9pJrcv4oZk/fTeLo1Xl7bek4dYCQyXtlasEOdLte
JcpUZS4f/inKNwSRsxrINq4wEIt6BVIx2bghXG1XK3+nALGeU4M5YUotjvpDSEzK
Ri3yur8uY60auiTo4QSsaVgLGsxWouzoR1RXYUHyKEKdqYXO5zW0ULS9GWNdQXOI
AqvemgB7Dj0KTGGM+QRS3uoXKSxN4eJXoM3KCA3Rq48hs9uFuX/9A8F2VfeS41M0
3YMg+a94vHQRTZw00Q2tALpiHJgIeHpbPI1UAbITLI5B4fSIDbdNW0XoevSUikxh
ZycoL7I03GlI/tu8nh7EXV5htrOjdBzDeTLX4rd4XZVGyVIIEFtYyJO8vRmLB6bl
zwyZuzEKCfg7p+XLqGet7iTexThHPpqp/WeWD4aOgRaIKU3AsAxKUkC1B6j2A/oX
18xBK8TYzf3PMj2ykEGMREo0J3s5nbUtir432P3+yBqUi18oTl0Q+RedKKxc0zpW
wOW2fkYujDVV2FJ4bF8qiONW/7FSHBZeZZGiqBPbnZOSkmXpJhnGAaw4MXYIeY/l
KVb1GfvJA4biGoeiXc+IlzGBJxHK1KeF8eB8KtVAOYmiKDz3AlAoIFdcMCCe0hGE
dHESCWGO/OVPCl6QENr37YWhJlQkA5/rb5KwTby49YCqhb2icvRRE1InL7WGfY1n
2ADddJz20jFJKVRyKrbvMxun5HrrG2ep+F0kwX/WK3n/y5QpYnKb7hfw89Sg6G+0
WMLq8FcF/U6Xp/XOzBt6UXGnAnKMHQSAgaq6exsmYYC90OV5aavAPmYrN4eCVezy
f2KKOg8/v/oXWEZYPYJcSqpepfzwLRlpsJK/h8wwA8323LJbqs8CjyfYNIy663c0
4qW9/EnCkQR23YA+jPriyoC8s+0FHRFWUaNZm0fNQdfp0RRsoEb8A4lx4X6UFRDl
6q6RHLAUNyqBzO7d7IeXvbMjy/zPijAy7tQzNrNKugBOs6GiA/HOpqHvy2Kbl4Iy
Q4EfOEmxc8289rsuQx7iTx228oeZYrzw2BXwAY5reDb8x7RacY0fqSMsGRcfWoyd
h6sK5x9U3KQ1idUl3zs4lNfy8L9MDIvCod2HpS+vXUbiGIcU2iir7hdvPH2iLXGL
Vhz6Je6UeoRNoIhYbT35sRqVgfKDWKmQcWQv//CK2uLP/9eqAuyRni6fi8HAnQVy
FonTGPuYHlJuVDLxO7B5D/PvcJ+zQjRUw5TsMR8+9nZJUZOpWWy2wwjR2BS0SAGo
wEW45KAY3uJ0nEPxUb5niAZcitryYjRhS1PCFeXu/FfJmzz7fMqIYQ1K8ooD5OZ1
DgHutFbct+s1RSd8KZMIX2ipsQKaVvue3RpCnLHMKAJY/6r+v1WpZrLKl0+eFGYB
HMW9NxuM3NTw9wpe3V3SdR00ndP87ml9Ovw3qVSGFpfNxrZ19fDDdSUycUwTKTLt
vx66jc3IVBKSMdNFK3CF3jQSxJg5Hr2dnaOMnXY5Ut4MQEaWQb9su1rrGXOa03JJ
gVjEPfdG6HQEb19pXAmEpDAf/SEFWU4T5rWhWK6h0Rgys0aDcgiYjwDUtQ4YlaOe
G8pQ23amGaeybJtTOkOluW+JCps3ERRy7fhHKyKTooExislHwBG9NPalWfQNBGyY
VGpo1FoTVaCt/6GG53eOwTXaGdws7jhvgW0uSBsBErqxiiG83aMAVCrxu59aLWcY
yRCG6oN4kBoLT9bgRso+2fqPZxzSm3RSTNxGqXvd6KLhmbsQPv8KHFhZHnNiTzCv
eo9jr8EI6l4Js2ajX80FIIVai+vuOnuYZxtPlwcR2HTnd7tZnnqpL2xVrfp2+XdT
ZLVi+Oz5NbTUxZkF7bI2NF5vqB2791GfQOicPSpQ1Nokiu6xHcbWdBiZ+/RRk20+
QfWzKKUeP5LjtTsoPvfL1AF7nsFWuNEHWyHK5nXnhCOXOycOSfKBUmo998LUN88r
po47vJEdoOJXDsfe6GrVAHv9NRBVmaJCq3bvaShFTRwuKoqAdC1xCjXhYV9TRm6q
RNVGFhxHUQk9t7mlLujzFLTxYcxRwFlDNFRS4ZZiYgoKiO9XkxZ2MjW23YSOqeEP
aJf2ELKslCmfiij5t05GeI3C7OE8oydXImDVxed4LVNjwMp0PikRFn3KddryaNHg
0P0nbFwWsw7yE+N/wthWfeUIGkhXI8QXMJ6fphoKbKpq/ZTeKvWiJjWYjgdGmDvG
3ti2NluFu1G2DTY3YikarJ5LfI5AS14T5d80yyvCPO0=
`protect END_PROTECTED
