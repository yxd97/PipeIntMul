`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNCN9JiskugqY3TRH4YlYNjz/fp6EX5gxmjHKg8uyDS53XYaoRiAOO7BkeBrnP5+
jmC9DIqP18vh8RKb67raew6JI1LjD5RMQuuZWyzqLnoIQmi3BjytKcep50dmwKbM
rT6fgrVIbd7bm+11aEtu9GcTWq76lWZdvHxCGyBrUXTO2cMNKcJk5GdUfWrb6GtR
/ehqMMWH4sz7/aO/UgkMP37d8J/R+cC3S22y4PFqSoYwsfoDIdaw0C/r/OWAakib
3zZNPTiRIW41KGhB1eU749nd+QWjIY8zkNdwBRZKhP6JKA8Vy6rzacrCjownGyoU
CZmwJVQEAu3Q023EAVbmG/F7FSOjHUKO+j9rr+WH8F6QF90uLwfNYC0LP0G07t7c
+2J4qm6mpqy5FecXfG2p7XQoy9Mrxx7vnTBj9kB0vWCb05bmXq6nB3SmRpNPFE1k
WW8JSSi9MEapTPZcyNDfs0UaTIobsK11SkOz3eZSPE8=
`protect END_PROTECTED
