`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ocGIO2nw30CrJwzgJrUOdU3KLzzR0tXYZVKLcXm6vHGqMAWeKagCHoaQtHAcbJx
ynRduk6XYqkEZR4+BfCrQT2JABTSHfIQkcThGvOKdUdQzbboSmlX3DsDabYieRmj
f0cOXiddLiVi5RFAK7X9YpT3pkTf/LLA/vjjbIKcg69UNCNBowRp++q5Vjl9l2il
+CIP2RyIhUGYTBlpbYvjYm2YmYglaOMcx/UEbqF1C48yIDLyopopiXnSQyLunKIk
DzIQgZqW1gWjY47GdUWTeuu/f8fE/iQmastyWvR2INsOvzoh+YMvi3ldg7es4Zaw
GSCHmi7ABslPP4Pt/w9T4o3YAYQZ1pPzsHhe4ek+IgJzybkMxZQ4x4SiKqsfW9r8
nPqIJ78x0MG6C801inmmMCS0bYDm0HhjFPAZXxCuVuzSE53TvvwZW+bdOiuTnIqb
zQ+kvGy8mCD5Y88ATq7R1Q9autOLbQZpxa92uhy+P/9rhBIxQq7MRWM6EM3SKYJo
tPIXVHBgzNDgu2ud6xIj2EVgaLBGDicGUBku6mz/q/VuiqebSIaoBerrh2X/5yL6
fj+gQzoZc6oTHtVWuh7Z15pO6+Y53+NSIHudfv+XWfQ=
`protect END_PROTECTED
