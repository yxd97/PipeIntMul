`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuUXYXSTOyb5MkMoLqjbds9EShzMnPfs2lz6RmAVonqmW57d0fpMZvKnU2ZWhnFp
D0LBSWIQzK3cSCT1uXHlzKG/bHkf1YCil3QZPhq1TlTdIhPCol8WPNAhTQJnhAUx
icnxKGpVAOh00dGgAvUFnI2EE8JrNWn2Pf2co+gqkeEBVfIsakJgu5LjWP0HiJaf
xa7p69nfK+6GkH4Sy+BTU2FYXrvNOyebkJSuZWpwF3FHnNOB+LteaVYvKE5WupRS
S8zZnJzcnpl7nP69EzbkMA==
`protect END_PROTECTED
