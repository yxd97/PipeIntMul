`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTSxoDzcMrI6D3LVLTitTUEsf/qvrzGNZD097T4OMs+cVVlasg5knkmWXMxhU03O
ruwXo4UB6saQvpcFPkDUjFLNhDx7jCidJp7buTwxf8y7L2/+nDUPs2sRTZFpMM+y
GbLiovGi52HbidXdQdAnli8rIqycLgVu/cVcvqqjEjScPIcCXiWDTgUtjYipeztW
kU1VyFb73NdlqYYvikoZ9yIqkOLHHZ2Xj9FIFQPtfGX/roHUOu3gpfx91RIeUUMK
q2dX/GH+81RodFXJJ4Mko9YshonBsHHLVfz8Va9iQI0Tdrh1PD/ai0Y7T2T9DmH+
cKlGfJckmHv49igCA4av2Yvk9qQyqtNhlGz4BjvZx9cEbTxD4pxjKFKnkpZQPDKN
zWhkcZ2T7KuzSWBJvsH8G0K9xEMQ4NgMrg2XqaXpWX8xQfL2nwj7Z5ZSblotASnb
jY4c4JLcrKlBjp4RCTatjXvdBPwDnyb1AIQrhLa7NM4fgK6LDtLMvjpS9tKKOWii
J9nRf6kNDQkCN/lXGJSk1JyfSlO8XPEJPHGgHanvqAXLvMiO3gOCSlYeObiSoxMQ
yCzkBSXUCfrtKX4kpHgHrEn/K5wIuDJd6SLCxvy4bqjZgcikE2JHPcC8lDzIpSu9
ClgMl5a5TXOIPDimyjja8qAX/uTxRbFvxzo0IcPxfMqgO+BUkG3kThYRC5hxfBz5
cidM9aD1XFl2idRcNIiyFQ==
`protect END_PROTECTED
