`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqgYJ5gl4eD1wjVcCmsHYrSh6skRdOV7cQSjPM67cAHF+PE/cgtwiIoZpyV7Jw0G
BHxnf6f5kiZL3CZga0SioHKadoU70HZGu0vTPo4KLZj8HM7Gpewu1RVCj/0/q704
XoQgfFTxz6YY+3mZyq+FlwDJ/u/7vMCeRClaImBrnGiUR6f/WJtsOi9Le3l7gvNb
AYd0O5/5Mz++qUxKwMCDxOihLKJ7O0/zKM61GfuFNPq2FOdXNzFgF7cJPY/SBdJS
DcvtEOdqfcrFZapSfv1aOdWLACG64lrz7dKzj7/zvriZ6NpK99j8AlUNaY7bJFnN
c1wGfIz4IThO/3X7tZK1fDumBtTSKc78Cnbcv0hzARVd945X06IMGK6Bwcu8egxf
nMIBa7BqLrQQGkzPq2+M5ykuuFi13AOzCnD6QNb8548=
`protect END_PROTECTED
