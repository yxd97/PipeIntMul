`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNAlIxxXRV+jdIZ8SV7/348biXh7n1IQSdIq55fdEcrufZMfVoDBB2YateLB6Uig
mCITvpB30O/mmw/WcPKQhimphmU5qoa96xF1OE6zGOY6cYdHnSz6NMkbnQV+PIKl
vB02qFouCO3RzHM7MsoMWd74+QK1XljuvbOlmbU0DfTBbXO8Zg21JLHGw7V7l+HD
S14Oj2i1ZUiMTo0U6UUHzWvZm6A1BdOc9cPO+0cVKFmtxrnTZI4aLpnCVGRj3bOR
+3OXT4Ge0oqS8CoO9UCq8e3Ryx6lTvNpLUkQw5KnOtU9WJGm+fOlrlwmXk1+DlWD
j6pBC2/YR3QnxN0BkTKuRxcXHZXi9agPMAD8EwU1NafItgVRbV9FZitnfyPxcnG2
fwB98jwQrrl25T4T9xYt/cOsPo/vA6sh6CA7tSxV5nByZ6dtIKdztOyXvF7/H5Fy
TiiLU7OQKlGNi0d+m/h+4KCGdA6ZythGKOwqMo7TzyIAzVgJSCjD4/RuFAx5KMlL
uvJYOXq7wXcGIlQH9MolAUz5fJJCwhUdOHV9qCdvKC03xAKFoBMGZE7Vd4QfXZ2s
`protect END_PROTECTED
