`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2FN1Xq5sFQ6tJ7vU7Wn2MlctSWnCZ6B5vIJMqfqfasC2zkq0h3mH/xKsOC3QfPz
25SyLiUyQPCQ1eclMTw1FxopfqquBuJP03mdWPc+yFiQGI9/zRwiPB3VFnNwzjET
5THEaokeaNwJaPKicuAnTE8HUStPT3ICYgRNfhS1WSezSfJUlZscqzBgabh5O/HE
DIn29ns7JNkF6QmB+yPlH5tXBfvZHk+NfoQUPOiwYqWkSiZV6vi6A4Pz4AgBOQHy
VsD7IJlta5L6X5cCpkqyzKyBNylYf0EQRheiV0ygfYb25knHJRcrCt3vH1KIELj/
bIF+dN+C/ZkjivhndNyOE1Nmpi6pYlAtI47SWTa+KsDTi0XkMJI8yMT2O5ReKuQb
mJj0rke69PTqSMu6ib5WWKPtfv5UFyq3wvOx8bkhtLK7y6w3wdX6ays2tyEhYRBY
e1r1KVDE3025JGegM24xAEe6irUIPqXQ2RigKQ2H+JPG+Dx3fvVdfd7gHx0VAKkl
ek6E349feLTUlU52VFOUFzEmTFvHRPeEEDiL65mU/tuQwd75yUsu4+rw9rW6jHJu
GNGkxswXT5gshq64M5l5USDTIKGFlmrmEOqxy/5WYEfp5Z/F5mXww/aMz0VrK/z6
hYlaHgnIBDVVErlvFTFy/wEBSIA0fYbnBmKgwGVl+kWdO9aO3CxAo13cm+6rsa7t
QaBWcBYGaDyro8nPHBSTif6XyA9W6o23sahmhkmCyaeHSZLxfoqygHBpjHcjr2Y6
VluZrpXFda5RUSTUyKNuVccilqgobIgrNa5ABx78NPldISMfydBdsmnpfp7fYjwx
ucBw6Xu46nhdy/vRplxEXzRHPsItIxnTWvDPk/k9kmGPvvh61DcZkSct9kapBsYw
UlKeuJNzcfjlSBgIjXEFvGrLwnLJihZLWRKNpWCRv8YARiecsF8U4Lz+huYTL9ST
Ey84FKy8n762b2+JhMHedJqIAZIrvRNuTuDwIUDRv2u7Bg8IzzsCtA5L7TeGSEcw
Fu9aYhEIShcthdAmPg8yyaXe65b3y06FoFlasxlSc4KRD1a6ph76QwoEXlkWmJKI
d41FkiC7zSza4UOHNtIcK8VZWiL/Hm+C/hvYlLgpkXqT3zzpmYZNfIMKdh/L5eVA
fonqgrQkHb3kuOCyrFYU0RiD80wp7KpQi+cm0md/uDVnpdOLqEC2IOTY1kBqh7e7
CA5iwqlVFBNK2SrrOF3cYD8RkvxtWe1GlwHAFAI/+KJQamFtQh1aRbjXemLpOI5Q
LLZ46cWO4lVLlBUzB15h77E8n2pDfEmKQgsHXGd7zUjfpb6egFdhM/EPG+r6kE3r
0zlBmrwOgyqRwCsXqvBa+80v7elwZrz4wXDb+znpNJt/Wb5Dk1KJ5WVnPOrjg440
`protect END_PROTECTED
