`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IoKnKpw96ycoCPupcl0rrbxkjhpt6ksynnEHZPgnB8L1F15WnKJcj4VAqsUJBx+m
zdcQERUaQUJl0XuZQlzfpPFsvzg51GUJw2E6V/XKe6T/FCtQlDS2zLj0YOmZOYLe
F3WP1LP1PJuBhBPR7iwurRmKSwNeonj9KxmaUAedZp7ODnxGZCPEeqX2p+dY9YZI
1qqpGmBnWzCum+JL9U1b7JBlImT27G6dNs6IbyXbyPIhlK+pGucAl4MBPRleJ3rX
6qWgOVU7jgd0hrubgWGxGaSuW3MucJMUGTUClNE+Sv3kDS2iGCF4UR3mE1LrF3Ov
wO5Hn2HFp5w1V61vdWXTcgJFWnOcBp6J76bvqOEEhuwAZ2qvbPub5MRVhDU6pvVD
3AkVE+JT4YlU+X5xlrarDg==
`protect END_PROTECTED
