`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IPfKLt3uVOLuotaywbfHKJ/hI2EM8zTDVMBuFRuXfVCqQFK5AuASlAR5HHjwC4/Z
AOeZ8KXe4rryGaCGcwxJ1ETNKJ32ruADWqg/Ri/YQnvwqiSYy1ZK5Gj0cPqDN27/
nzRfdY7kQl4JVQf98a9gWTmCU7wNqva3yW9ck+LrvUUPPGWH16Cf1Dlv1uDgXU75
1X/dhBPATZnf1ycI1wA7MiMpsOpI/LTZMlM8RFc8c85YC7YanaCD2nGJD9iKpv90
nH2D16hskTH6NNVWcuef/yldj/16yIg6qMB2hSuhS8M=
`protect END_PROTECTED
