`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JC5IQ7VTed0/z8zb2D62O4EUKr8HkD1KfF9BuuodArAd7Bz8B4Fy4h02DJYNP640
sN4IR7PT2hK7JHoU38q40FrQ0yOpy5YT+g5AN+UNapIDHGO/Ht79XU0Czx/hQcNP
g8vfUDLr9pCIKV2keMkXICJfZZ9hv9ga9rEhp/+/HNZNsv2eZ77nuyjWBUX3+rjh
vfZYdW3436Q7etgSa8VJ7slwVvbRjLDTF9xvmx7joYrOC+pQrRu7NzWta3cyMBxs
Q6/Ve7gi7hh4wOYqs5vvG6/HxKP9MNPk/w30UaXmRzNcRSpZmgp+gPzPILnjwQZK
bCPdXu8Hkn/roB56jqbwTQ==
`protect END_PROTECTED
