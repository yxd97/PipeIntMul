`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cF52pNkFIGHEN4MH/0dC+HC5ND9uP3hrraknBlHJS56FfpfROrindI8zWHxRlChi
3bYl4w305BciiRKTSDNXwlXMXvTDsHdl6DUwlwNsxH09rqilqurfiSkdmdNUe9/z
5zaPF8y0GRwlej+lUle4sC2unh1FWcE/USSU2uxPipOv4J3Ewt7IKz/VM8XgbD89
OatfhNQ3HyPj2/6WUjg9fnptFu0ZudzDogJrc1fAeKPQIIfDEzQ7o/J35JtQxgqF
XsSkPNvaP5ecTo75KoJPM3hKAIK59picvx9HMHjfk8O3zyIFalEf9mrye7p6u/ZM
nGWYjeBOklbkl7pNOLcxnn8PwuiaSQnjAGJs7Q20HR2BRao8S5xMCE5MWFKY3pTi
uquz8rLJTpZxnEg3TAeZI5S2JcTlaZr9yH7ZrJ9f0H03fOs7g7nGVKakdMIaUFyR
yNUKeZyg2ouNyw1JIX0VQc5o9w0TmZYvly8ZNXAU+DL8kTrNdHp3M+qCAbLu1fQ9
LGEBP9LyMlXExSDgAjE5SioY1jCO1gQTxYTGo3aj5hK6fiZeMkwTO/UCAf2raiKh
8u4+WRkOSL5D1DUAKVZpPAyeqgNta6QJHEGi1liEJOqTx44VtWGALZnA4WDQ4RA7
W3TfEPLE92wULkbWm/VurVwFlsv4OdWO2X3IKLYyu2GngULEj98GK2Np+f61VjKp
x5Oy9/iAbTCy+4VuE5UzzPASxluooUGBygsPQQDrcXPETHzlspp/2u9CwIeurEwf
xCQCwJIJAz2nDqOFiPpU40ME3pffoP9IO9Q3qafd2KdG78RaPmHMzwvHOKO7b6S3
F4S1pa6+GxqqlpZ1eMr9huyhXAM2rY2QXnk0lyFSnxCYGC+PnwNC7QOIcISWFyOj
Kxfp+0Ddf6ijix/mLamNCJ7vmusf1Dx2+PCuF26nGLr5C86c2PuJzuWxjVjdZ9C6
lyMvIK5upJfbuhN53+VVKoTyiQQSu2F/QdD6I33xRfg5nGQzWw4gmpn2L+OimFXG
Nmg3qDgGP5ou1dWLkCgowTj8lnfXDhSrvGBiNCcR3NcFJmeZtXp2+5NxrjlSfnaS
QwrjhKEOZA3CL8Wq8Yxw4KO4B4RbhRgkgS4BX3GkGV62XZgPYFstXLsrUcA8tt67
il4xmiHBt+0S+myG8+2zEI2lwPOuNHvyOeeQyyDrLoxiWsz+rHfVCxJXlLCCVmkw
jeuuEPtevZIK7e9v3nUyKOuQ4SooXTZq681nINjGNDr//Wbc+tls+zbs2wKWEGZA
HMxzz5m0K4jOZp8Ai5yuskA3VeGmJvbXi3vllyvQ+C7h1E/rBinZq9MMbwQaCzsV
JyLfeXly2scJ6KyGxQejL27N2SuUu4nlmvG1VGiR9ipM4XhIW0lUJdP6W/Z+g6/Y
5SQ3lgrNkLUHmz3Gg667gqRglaKFdTJM6cyuHKUl271haMB7PG2PWcIC/ql1AG5h
MoDC2DuJ/UNX6t9e6mpAuIc/DKhgPYoMBfyN7kVyaktjrEvUvUhF6APycHSob1L0
NuwauD3UGX2bp58fAb2Tzr65lPdL3koFlvyOx0hoPhFVOhI9QsNztB7HsRYBBevL
Y65647G09xo5bsyOROap1VVHky/pvT+uhSqto/FRKqUFY2vNih+wzwir7tbuPEiH
hxbdhhWapalawzp/gq50yX5+RvHgYjvNKCS4x7xC66zdJ/9myipwLDy1YaBqQtbC
O/xFb1IzRPzW+apIihM++2JVezOw8VA2WXBEHqzYoKr3ahIzSFumIFGcrNp+5Z0i
GmCa5cOA6ElVo4SDmnaagg4/SoH/3jkrOv1FtMPYUa3d19TgzWgx+7PqnSohFPDG
vAnqdefWoBIIrWiaKji+Qnp/CkkO8n5zB8oBp2ix9GRDM6Cbwxe6/qCtkVGGZPxg
OQ0hAhNWVKXRbrYpaVK517cNaDNc1IJdqbIpngQl/aED57mZQkJZwZMpPjHEyqLF
5HQEHt6tMQMDTOPbyk+ArGbaWiPGStgUQhu9cn4/F5UOdlmf/BUVbb1ZZWMHcVAO
1G8Xd/x+/EyaS6hFYioR6/4TrxCHpMRjAIoPImXJGVLjl40sm4s7uBiEbrvj6bK3
cJrbi/yt5fAAEEv+ElGoxxXsktny1g8gQIHWwAtx0xA2j/Jtx8FO0Ld3Q6HtZhwb
noWeyDMDDHNWKSjMwwT7TicmzE3xB/yTVAECdTYscxOtjrDlcJu6F/1jW3M6lGvW
z5DnaXEqyRe752Kd9ntGu1HOggm3hJUeatHpPZV+bKJBxYfuctxFtTGKEi1x4kfL
9+bFelv9LwMTq4aMcamBjpsX29X//d1krxP4/XnEo5M+CR+5IkB+mdzYTEsVZIfQ
ipqCY3+CPlhS1ox5J7BCE0QjK05OLR8GXMy9JZphcagj4OifqkKVO30MLd2KenPF
QOWbz9RUtpCLrkzXMJ5ckFfDH1g7MQjphbVnBM0RF0qlAvG3+o9B6yjXKam7zZov
ewnuIur4n3SRKAxMJGYhn+iAD2VSRtU0hd18Sr3zVhh4chu3o6mYpTJlUoJ82vxj
J+BND8cDDx5/4GLpgya1OWOIsCUlEf/Sd2/pex6M3gGUt6xHERVFjXZnbjDdiina
YMwe7HZKTfjRXIFyqjJueqUKgu1ucSjxtbDizBdRJg0dvtGzbY2D5ZJXt4UIesX8
AhP4D6p3urf+TZyu5xqKz5NvgTlvQUgV0/Rgzg6fTRqpvJuETkr6aVjK9TwiDgDf
awT66GOyXzlR94pMuk9kEgRZjhgZJW+WO8xw9sBkiMqlX1c6G71WoFstw0MJC5Wa
cxZmiddJM0/d4MgCQrxwoqevnFUkfv7duwG1EEZ1Ut1iJY3TyvJoqsivn1Qp5/pf
oaDB++uqO24m3XXvCjnZndQ2yFPWiBMaWLRoVlasYFk8YLXvlruo54QjDYLE7rpR
L33TGwIsHbktiJw4YzEuLov+NGQyUv4/tcoLmkoW31AwMo7qOFWFHpizluvlQlCN
ElPFqlqtvs4bLgfQZQLviGU+Egv7/peVDZ7JsHz0ZK5xw/lIuLFoJKdnLtq8Di6Y
/OOguNcnQBxrtU/xo8Y+mLJrpc/+lkGNVWj9w/gjejFUdx4BwoWVeT7+na7/yGoz
mJXFXtJMcLQAjreiEztmItNSiGI6l/U8qtTANl5/a2+Co1RvgfPe4QkyKTFpV/kd
GSv1lhgcdj6RNvy9TzEV4Mf3+ixfHxeb7A62UgYQs6K2vvigQT0UVmEQMdyVmMtz
42ZmJiKhMLmg02sa8AxGWfjnn2xlqx8NhbrskGVB7/ymRQuFPL8euwKfEJ4iZTJj
CO21g0QrcLZItsCpMKI8mBHs7mk85s38juppJFMhWroA+QgR4ElVCo1GstJp3nJU
5B/Jk/F5iHKC/lqaMbCWSW8srfVI7yK9ELkjYVjp7zY4kTsedPqsa1xuohLiCfJn
Nkcssyo5lkm9gl3LIGEAx0auMTeUgQkXa3/p2EIMBbU17HlTBeET6WD++o39Szcq
sQ30L1SbWGgqMId6NfLxj1FawdujPld9EOpLQKuE+PEyxJpm4raaybpIg/mOoEWm
ljrcE3z+mrB0H66+6AeOjSYTTA15dJ1LMma2MCS/J09XEjc8Bu0XJgkIeoLJ68Ab
GxS5f7kC8g313I716jmaCuZsbcYyI8ISaspovz+E4xJ33K0xQ2Ig6OL4jkSk8ARn
G2bd+nJSwGER5vD+1cWfIgmGilFWXLq/iyJmRtqgHcspzSvBEW79VzagB5sTcMvp
UPLmUKMh4mT9Bdk7dYklAGNrOSQZ08oA689JNaKqnjXmyNlD5hXsU7SGy3Uzpj8K
+/8KUiKfoEpE0+Nh872dSxteV7tLfZp4NdzechR+TT4wVRZU3WR/+pT+YqkgM/LG
8qScZWkq0jGN3DPtX0jk0SkTMtAV3GwZ2RkzQAyyoz+QU4nCzbf77Nh4sHoy38dO
axAQyodODYQF3DW27yP3Gv0ntqGwpJgErtX/hVu+BOn3ZPH97G60jsahX4xx6X7F
Ct2zUQCosm9s2k4Nl+VGTaZgu1UO9tDiSHew8tj+UL3ts/L6IXp3s3n3uhWYL2Np
WPjdLULbiZcy5lo5LhfkZh9wW2XTh0ATEorGKjxF9jQ5Pif/bCSeL0BZ1+8YAgmC
/lR7UVDuTVtiIVR2cGuj4j62VyI4BxKVfMgnzetrh6uy5g1OR3z6oUzhPHO9dfhY
ny5m87s0hp/jsM5CvddCFifpiGNHQ8p9MMucg2yYJENfZRfFDHuOlGYJEDghKvEV
JXQbGhscSXdHoTy9klNvnwTMZ+eaPdpxdl+3Od4db1hpe322JfSTx6mzy6FWb/tU
pehY0hLP4moHem4CMaeJet3guxR+1v2Ve6Z1mzpIW+2hSVQwgd0xiHZs+pC0VzL0
c4KExHp2zuQBosvCeAyv3cA6hDNhbJB4tWlnZRpC0j6+DqkODZVcDlLGzL6corFv
jPzZTH1CQK7gyWTzNwhwYTaEZ3W367z0E5BWuHdZWmilp9Tij/Y6YAU7eGyzleT3
+jWYmq1VeCXE63Ogdoqz3uU7AGvZNXylNgKIQ3KPSMSezxF7cCjuTsLBviuW4Fdy
/3tBF8A4FKhSjq3/eT1HiaS917iwjC0OriYqpfm5/mLJqeP1qefnKld70/9a/sdG
lVbIXNGNAhpUNtBQh/cH5r2SrmusE8/3IN3jKAemase1DUlLGvHMPCbeD9QHSgT+
p14QHxp2CsYhiv6VaRpGXg==
`protect END_PROTECTED
