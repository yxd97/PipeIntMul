`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g0x1Sly4raHidhH5rCKGhDLVVEwc8KwY3/NAM46+VB31CtPFc7Jr7QlLezrSmarD
EvHUaUiZC647WVayNBaeFLuMIN/HugZr422Pd5JPQwjsNBjNGZjhFsS9maN+h+PH
TdG5jGXx3vXgucZm7XGdR9Uacll5r+l3bnTYWx4UYsDVp9Xwa8v1gDfNc2vjE56U
Z26sNNvKAXKfMNMLH7ASGI9gwFBsVXZMxxU9bfzMAfa0edNvE50BWD7gg7oZ7DGD
bof/Abf7aAEI5NpokSCNPE8BYBUgF7xWsmF2B+XcJZi1XWywPJoWSgcHfPaOirTG
PA7iC97eLg+/db77MXa/kO12CUaTIsdyYlYgC/dJMpz/gp+FLVr7anCGOO3grFpU
Yb0szgbWxOXuAziF261tPD9kr+2hDQyLoASgIuNzobXDUnsD/L9avoqcQrslfPCX
kZmeVz7jrlFf8LBIOrs2WR0nK/ny0+zbl3vFZVpS8sBJRLWpANIRZPZMKGQPAc/G
o8Lz1X79FbFYS1HE23C00p+MZyu6C+CZ1phOoBjOBa+AbBvJlwPHuJb16lkHEBhu
`protect END_PROTECTED
