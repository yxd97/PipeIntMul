`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axL/WpQKlsEqmpF+mIHz+zYp7QkQoHR9kHVFJIjlLnT3vAg1kJys+7uviIC6jLBz
6vhYCQjNz30kQo0SwOCcWPxI9sg3R1C8Sqe1CdJdTTxtfHMpGuV/vVKtsK2Pp00A
28flR1JIZnxMWCNdsewvVMHeF4GiZGgVrluOeb2G89y1/2PELwYwmNvqKIUzxnf3
ryjoWRGaWzSC444awDNKHiTNCz2MmlpGv2ngzhNrqJ1RHSTaoGyeuRXJidSOo+qd
dGPXTGD/tGxTq/Sdak+pXX8iX/HI6gs4TwjahdMi2r+k1aA5AUsoibS/WdZ02HR/
ZmEDFMwAr8GszqcBlkTNrQGdrpurQKhFcQSaWA7KEA3MQ8nDlTzb0qANBk/uEyyY
2GDWfUKavcVm+6TFVlcq2Wi0zs40A+RGFh6jegXOK2iRKK+UrfGT39T34UTxzHWW
PGO5fuP+FymlcJnUBFJjQXC9ItMpOiPsfXiwaPok/+mkpIvZcTeycs4tr2ulw9gC
ClklOjr86uk7engmfBnSp1S35MmtB6xLx+MiZVei3FQxnzJHg3ZRLZAX5z0RanKV
umC4+VQfqc6GikmqHhMLhg+QEk4Is250rUTG4uCMvZ68aYpUHvLRTTiZZ1sSF0rC
9cBjM8W5qUgnEIaTQOBDIKCkkcJtTf2nTRt7BPULfWlSUtl6ACs3/XX7kMttt86A
cOxopaAbw/RAsuv3f5DhjavFmSPpeQCboKNFSB4Amfd3c4jYPixeWRr3lcWXZBVQ
+NNjGtQkD0TZKI5LdDR85Wv+HrhQrcBz1j8M7r9r9AB7ras/Xng1Xae/ojtvjQBD
LGImd1EjwXWnETic7a/eB3WrvfC7pgvN438BUF/IsdDH4ZtDro+gZIxGriXjF8hr
0tVsmYPUNEsQ1adA6pMTLw==
`protect END_PROTECTED
