`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyYcVK5wt2+DY7a9qQWSO83oVX74iEV9N9GYO4OkN091W/uMqju/rdaqtz8Yj3qP
bOGK4/qiC/Dd2oeGnfdAz4M9m/wCwMfFpbpyvlf+cNew51uSIEwj1huCljz4F/WI
74guSag96/n6B2OOsKhnIEsbA9ihBdhMX5wJuVj+9EMwOLaqOWiNCEw6wPUSsHDZ
lzGsyfWuUUQ6SGHfL+F59DW6UKvXFKfMZBHQfW4VxgJ5J9C8BhmpD6X4XfLrg8JC
g6cDQOaZoxguHn8lV6MKPaK3bM4vjtADyVrORNZ8p1x0wDECNHO0QImKPm98BVUy
VjWvQFuMXQoRkeRbwXu73bgQB/22VfWWPQMHo9ZOzTBRQrE7K9RcvXYhbDfCCk+6
LRMsY/9YADMvz6bvml0NOWvzCCG6/lAcYQilA4r9qf4=
`protect END_PROTECTED
