`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZEHQzbM5u6X+ZrU8W4TuGIM3oVaX9skKnldZEBYvfS88jG52pGZkIU896qrzYLj
fzuDdiqfNWnchJjXtm3ByjLqJxZ/SKLCNz45GjUq/IlXpert3vMCltPzYcD72nFW
R0M1CKcSFbGTgDzYgLK/1NJywyJGXwFriSI8roDCB0wEBzAcY4F3N1InqFsUjQHW
tYUzFx6Pn439Gqhe+5iAqYDvCJBtRNGMIAnInGfB/ebX4Se7PssTNKpPAgNAPlL+
8ZYhKW9spd1zIsLGlBdBZZgZrl7rAwZTlT3KtxGeeCudvI1j01wEaUUvFSlW4c8M
YaKZwnvjLsxTLVpVj4QW3g==
`protect END_PROTECTED
