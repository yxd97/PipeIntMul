`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ATrbvMy9HacCpEqOyOpf8DDF9EK2jt+uZY65EMwdVs8XNohGm6whFLg54xcrEWKI
7rWM3sBowbj92I0sv8kk3ug1l+bAQIzj3yzuHoZHi6zgtQHeO19SRuR+XyRCPrY+
v1ekA20YjfDja8KTZ4kWkJjxVzLSZLAknD0k4iIGzV44CRJtx5ma7cTl9ZxooElH
CzXMI3TzZsjG05tUO0RpO4Mcu8pcfzLprlN1Ol61yE5izdgeWb0rd6CXAxeoYQrM
b9sMoM5hXQij1n3CLpYEd4f6JF7rz8hv1cN2HMxTUgHCn2BJ+hvMmIWuUIO9k0S3
xIkcZhNx7qVBLBPfCtyKs1EAwmEUxHnG6Du/VlxH1zwEBXOQBDfe7OukaWjT3L+L
AP5qwDQaCkwFNazrJdYe4ysL1/tpwecWSrJho306ORJYjx92A6kqRC6YZVzy9QVb
yDfhpFU4zyQPKkWa9XnxDvHFMdL4c4v29tHxN91Er4ZAXKe528leiX+y9cHkhY0Z
L1keJ9cTd2G6zNj2YpNrhE0O3YWnuJCjM2abyc8hHfl4KfxHs8Rfsj1UxjhkN+s0
W2F/gxYB8lvKiG9o+td8qQxVNLPKnzeXCPHWyh5119ai4LOuWH27Td8HAIfnR0nm
uNj8KLqYKjkxHmcf05QCLFp5atY3ZFPXoy+KmbmVrONwJtYBlG+DMrJ3kwCBUhrC
`protect END_PROTECTED
