`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oFAfRfJONDWjrLaibDwyHCGGe24FINSBt+VfqVO7TkoD+1o9IxtBUY6SmBl2OtxK
W5G/815T4D/WmFiJjnqGxdZyS/rsozcHLm72HaVLuZop6Zl3tXSv1vxyLh9Ik55z
Bpbvb27TxzelgHJ0GZ/8ZsGLpn7IqNfGoPUL1el87K01c7jbKcGG8PMw76rBeQ+S
EsK7tFKeAE1xMV2F412a6aYRx6zrsjkg/FpxxjYz1xp7GTZvG0RVh41zOkXzpQ9b
H0yMqcKwNjkltRlufH5cmALGuOTKZUfOXGv4nMJ6LY1YN2MI7XycwzAnIEMlIFxw
arJvIZhGU+JEBv/w6S9rbx0TD4SKPZgH5J/E5Z21/dgRyEnbWVBNFo0MP+OxEyVr
uEDFgevZJYACXH+nCML6zh+Am8GelgzO3RXpp26BnQfPoI1LTbc9OXYq7bSNg2aH
z3uQcIz2x5wZ9ct/11ToJ6GQdzqBbYZa2BLbsAT7DCJlbl3HJzlVb05oqRiJA5dE
`protect END_PROTECTED
