`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z82B73wfuEvnYeXUqk+wF5NqkOk9eE0vELYZNeLpCVn5sCe+Zfk7ZLHdpPsCn0J3
dmKohfctVdoI7aL8u7AmJ44KGgDWtGaRQv39+8we9DW6/Ygq94Zr620uKc1KAOQq
6wbQq0MHh7uJRl6Zywvz/n0DZyp5xjzV42PGm3SBO5uZBQ29ffQCNWtE5HF3NKhg
gwM+sUlCUWuEuY9joTcrqeFMeW8SXIs5OCnGnQ0BgjcJDL5oES54KOQNapE3sO3o
WIK/S13j0LVW+bcU/ZZcIhGJhOJy730cNRoOr2ou81BKtnfVKavVZ9YTgrfTdJi0
lpvLvDDNejKuOihqdrMSdZr2bExGg3PCSScQ2cEtP55N+EW0hRZzSRV523OQQKvV
PpD9+LfbPNiXV0vfnsqJOkjdN9so+tUjfe83vh3BsRbYGeNqPk+PoQR1S6mIGu5w
kV3Toj6K4chJ3XEwB+xzTw/aXwrDLBrYNIjBJXJU6sb06F76vxSuQAtqlGvbHF+L
Uzix+0TaoAXfyb2fAEKwIqT8UNu0qJMUbJw3/pT+KfXHs1lK7ybVYHwlGo3ZKrMF
bh5vOTgFZYRo4i3ImAFhvvZH9ojy+xGUk6mcGSu+wHkrGlVB3SrsYyAiyFg49tmO
O7bJ0U7DtqlA7rx4qzXbQA==
`protect END_PROTECTED
