`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TDB2xjuYUED/fQaQynrApFA03NiDRa5CY+7QlV/UXMCtYtWrR/8ctSxBLc49x6Xq
gBT73GRpJdDpZ/BxQDNLL3Cv25OaTEi0UtcwgHUmt14CwsinGa/ReBsHAGKPGBft
KLU8Acun7V1US5LcrVUcRDJOdKUiPF8Rz9deZoC4PCTFMqsAnMJjnOgh5hS229hD
lIbZSAEAHVSvDnqn9oNU0YQMVVY96BBuaazMroLfwtkaLRx2JQ0VpihPGewVQMtM
ZdvqjnKLTXmDoTp3fnX/aHzU5e2Ud7ovtwAAHwAUy/Mv5drLyeobX/8pfx8+vzw1
Gs7J87LRVRUcqK+rR8X7jvvHi7Ny+ucdKkkeWC8liKpNJU2LVHcQqB7oDQZtDOsv
bL5NiWG5HNDlGpNy5/qrjFjibFJJoB1Y1ksDLon55OvPRFtIH6ucz62qentOkdLN
y1vjLIBBgEzB+zAEanPoNAkLpWQT3y3L7LkEkoUYJz2K4bWcCN6B+uNT9uxTlMNG
i7GvmrEuHQetJg/gBlbCbigCcqoE+fOquLvJpR8vV9907mnCGvo3H5KzXaH7rxwu
DhSVnNrHSmCZO9HbOPMOysmzY0lu7ufavd9FSyMdHBp5Zt1uyzXrUoAgXxUh9lcI
bu2a766p3vmi98mSUvwtMWh1lVvyS83aPZYCoNqSACW6DJmwDY7UqnQfYT6SAFyY
KSxAWOK2aoeGcn6G6nDMve1JXXve63JrG3tQF8UCOaxTtyLjqhPri2CPrXMC7nlY
1w4DOqP5TjXlQTNHND/iLq6siL1BAQ4zeDtqRntXEnglaD9jPWt3NRpXoF2/kyIL
gZk8JAtOHvxUrwa6DsLPLON16ykuJSTQyf6oxMFpSdnNSEOB8EyPqb/z/mZ2uJh8
uk0mj8DPbol4bxqVgFWwdS/XcDhzDPE1dUxGF4coSdg=
`protect END_PROTECTED
