`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DF96tQavzt4BcJQvrY1AGEdZA1kfUIgrDSORJW/zz8yvr9KSinglBLNN6ZftCUpo
G6kGebtOVuLPhmR2z0lb1PBRcYXBVZm4G6j7l3IUH2/O5bg7kT6z2gpq5AU92gkP
qehpF86tulq2KWAqfP5GfTfEtfUK6IKWRIxx9nPUvJWcpt9tO5vXP3wmEcQR+FCL
HC6NWmT2rqyoTA9I6iv1WY+yVPzBYZ7SspwGqWYTgW5jSrI48SRpCFtLgcMJqSGB
X4ZNzUBh7wVCvfGZjO0uG2j6S6+0/0psx/LZ/qbLajPZCP3eW5bDkDiv+1sqtuy5
+0HqLDrT46XtY7g2gvicuCvmbLYE19qB99ROEnUGtlvJYSNtd9uTJrg8DTAbIEFS
mE9YrFgFGEGLzA+rLo40Z2Js11hbt5oZF3ZwnmJ1vx/Nok3eUBKhOzFf4hQWA9te
4ohAiYo8F1iKljXmIF92Kg==
`protect END_PROTECTED
