`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqJJ40cF/fw3VUjGALL0NWz806LaalHjwK/FD4UsDEw89ZKZqxfmEkhAhlQUkZcf
HmlYAMveba/mSjIKw2JpxSRT1zI3UdmzxNOju9JRTJZ+aQct8HKg0qvkZD//6feR
UdogYogBsgksjTFe5ZwuKRsfPoeqSBOp81PFTdP6pzajy+avtWiwP/+CL1YHUHjK
MP/ebCS5ioOUqhe5FTeqnERuXF2PLAJsqK2DpAS/j9UAMb5+urRQhpxZad1OzPJJ
`protect END_PROTECTED
