`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ee8JtD0SIKBxpAW0yNZUhEDEItG9nOYp6SXBWa8J5bbZmE0bku7Pmsb7fIBPxnbw
cujxS0dlwBVAvcxw+1glc9zIfokwjK1tyny4Zks60fMAabeSMrNl4z7gSBHrcSuS
j9m3WE0Do4bB5XgzXdTp+OM8v3FoCk/Ru+ehSEIiwFzqQGvwlk53wxUbW0MGYmVs
0Eu0vuV+5aXqXyIc+32R2KjZ47TfuS7FKSL0TXIYcIv/xtTQBEV6pgVt0mRx27bI
eHT/QTgOqQg0i6TFMureFq//8Wdw0X9kmOVhjeoj5Rq+AJD9fbxKhcqXwQqP4mhA
+5mgD6loG82Pl/uNh2t2hm5b6/gCvYUej4hrbtVlI0a1bARzo6hHhi3sDkUpH/3k
ylYXJ0p6AL0GdzgjfB4tMcWB2G98IrG3Wj+hSFSWDI65SEao4F0bWvpIbgKZngBM
AijqIW1iUG4JcapTwxW/KazbnfdM15GPDxHNWTOIKCMKCGm5UvAhdaXJFk9Ykocy
LT3Mt7A1ln3aSP50aStPAJEdhqvOR2kujKR5R9IDVp9SAjGB7VaIRCB1dnC1jcpA
GrovsDd5z6mg70d52gMHaijmevYrEMrLkXABlWCd3rEWv3UcuS8L7ldNx/tAXeDP
leFj2wJnhi6wa+HPyexDtZfSE5x0bCwaqQ1r5etfcJ39AqkW907sceeMwG5ehN+c
0wmX5BR4t5HBcI+DwtMdDFukJ30zmhiTviu6sQ7qW2IhOiQQxZMNbBTFf0xrjlYL
81+RS8OkT2p+Woo6hEF41m1PpsKqZa4pWeIc2qANBneohoabwehUY2U/AAeCBEBl
hHtCyu+J7lN2JB1aFYKXL2mqi19xgKuJDVXFtunKoDHqqchz9V7qGgDyzOXglJmR
bCGh2PmDqNvK4fHrGN0RaofOZ99SXGfzYi5iKwPSWZkJOGi+YEmW3bgdazCYJLh0
0AIe/5YywzAWt/DLK0zhMR5ij0SWJciFo8ji+djD9yXLCYD+Kt2c0SfF0++rkiPX
QFT/PBONkJJZvo4i8afPYUDeCdbzA7af8Yz03r+uTnW0YPq1Tb0fgpQUPd9VkO/J
6DN7E40rhd2OY2zvnfT/wPZPrHgsljjT7wa+tyfUM3M+uxkaLzKrOEghb5Wlynxu
0CrAK1DzCWq+7Ks4urCLqqWDCsRQR9ns4swT0eRNdGjNQACRw3m74sRGceXUs/rG
kylV1qGTcMZqEVh+UiTlrmCNi/3scXP8fRzXuJDxME0bcOktvxXe0Zn2m+okrwcO
ggpmkhqSG3PCpbjso961nuIA0n+9b/JKN3VDqzzWGNv4CQDUh8C6WQAaifv+XdGG
O1CCT8pHF+DMSz6zvffWggGM1KCVbcy57B5qHekTH5ZD3/UfrpufTH9Iy96InDw8
9H3N878topg2lqsni/rAgz4qW+ZAyXDx2HW2RsZMNVlyhouB5L5p28j0b0ZWsb84
BpiNaQzZ5kakmM3uZt7l+8NNWIIOcN5dY+NGuDO8b2HD3JrUIw8D8CAyhPz111Aj
s6tSHzsPULM1FRX+1tYyH9Os/AlEf9jEUQFQOKOdaeKB82do55npbIMiWO5bM+j1
MMUAPE4zD13EHlsUv9asz3u4mggoc0cfZq9qaEdBNIDroGMKvfgayWPTISNxzPqC
Be/mwQHSMNRVMWZNT0ngwxIqPi0dpcoPMH0AH9o7He0FHH6q25yM8tIvJZJHxG/f
rxbgHsKZ5rRoge5ZrrS1wHPZuskeuveRLGev0+ab4e6ZZGGtywnckAo77qef6Bge
7Tp7xjLvwQDFXn4oyvM+mIpQqsncLgXOoqUQXn7BL9Vcmcwztiw88RlordZPqRw8
1jKixL80DKyOhQNq0v5cVGey3jH4nf+XZSad7hL9waGlZJdjHNNl9mztxRr1ng6j
dV4uHjRr2t9V9bXi0KFRssO/g+vriFb+rVuz90ggjfjWEQYLmaBAkUdF6GXYNC64
+KgBJnWjhkWeZPZPXcjYTw3jOdhAvvOfxr+AKhtVK2VHepzvNaWsyS9ryW86csxr
He30GvLaYFDEt0GYt9opAjiRtrHwaeT7Ft9FJTnYQc6sGOWrSeWoxbSXtus24yWE
/zaXUZNJcFwPNJo1OtYbwvoSP40ikT8GaYZT0RHqbVl9+TSgJ1HIQKmz4HqS8A31
cn2IgsWyn3J1aokqdLF7FGR1IfsKnrCZgMWnShsXfFN41gR3lhh2kN4NYP3Q/hWr
rSNXpFwYXKPvjwBtZE/2K1at4VVTohyQ1hvExXAM5z37Dg8TKPWz6Xnda9xqRpem
o2o6n9tI8LqBQX/UznRo3r68PR0fhofj6WLGFgUbc2Y=
`protect END_PROTECTED
