`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZDY+ESw0i8Yb7y5J+fLTZrjsRu9OmQ+gAcR7O6F0JNpnVmi0Z5Z2KoikwzdMlP6
qS1eB3Uyi8xJq6n+RaZNJMoRW93dcOj1sAEgnUbJmp0jDkdwcwRZ9Nahzrla38YB
fdlkztVoym7OzFzzf95NrshF4rEiy+9eslMomVPDkzwAEi5XOw9h7eIfeDC61KrU
4RC/yBeEJeaRS0BYK6cH84CljWA8134Z8f7aAOKMwmuADtEw+a/P2j0sO8sTbfhE
nWmqPSOIDOsbr/akSt689esADLa26R1Pq8K/PPmn6zUJVfiwFx+B6ZnWk8mcYXs4
scbStoRuFHAK5F8Vm3yottvGSh67/dTt8+gcBQ2CS7cKqbPtbn7cZT5+O4tysYkm
nucfgcoUV201W/McUmhaHg==
`protect END_PROTECTED
