`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xGOCo5FXlS1bD/ObaTjPPLjDMJXLPooCpLRT9/RhG0FoaNnw04iElK/XT4tvgVM5
lQ9FuLEBBRIuUQh9fgSGo0vwlTEpBkyazTK2MVkLwq5/QTsRlKigk9gy5jLcYD/h
dlIvJaRf+NTlnIiBupE8XtOJ0gsYJj1u/PkTHwbRiLFnMtYGYh7bUfWiOKEdNpca
UNzJ8YuTrJOaQ7TKBHQriJyymWSDwIyPWFw1GYBXIaDCh6hPUySNbokrVut08W0B
gS46WG07nGSKXIPCgAtUm7ZlwTZJ5Lm6LnM1HWDLxQznW0rlXnOAdb7zHHOz+HK4
P2TfDcr44apH4MHddBryxQ==
`protect END_PROTECTED
