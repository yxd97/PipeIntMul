`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5TQaQKj23HM9SRuubk4zUqIIoExlgC70ejphwshbTydAOltG2ee8XE8I7nYfUkN
/Hl93GFTF2rGnYRlaL5Tp23tkTjk+JZmtA9dTIRuj2jIlk6INIAUaB++awvCvSiQ
BGsWp0Mv3eGNTKmdzLP2H3DFFs4u+R16sq3WT7nQFtDE/eRNWVVbsAmdGVvKwPA3
A22iTMLzek0holQ9UXKPdDyyh52AGxXUMP+Q4ymDAQ6Zm3JfxKjysNiGHHcC++58
OgRR0jESKFDfPPrGIZKBLiva+AUb78FLtu8S6BnRIQezdiG7f9xWOwOjbNqUn2bf
6vCau+Elzvfw8ZeDAfMWIwi+CrFEYppKZD+G9/vBa1W+BAMQ/M0DAzyTof0w74Gc
cmSKiC8+B1wnPFyEgGn3I+e1F2eNSp+BTNBq/8bFVXQFfGFA4U+kdFsqq/sX45JJ
LTBLrzhpQMrjIG2gmD3KCLe+bDwh2cSsOFmnNHbUuZqQuc31mZ/4PRfeSTAwZhuP
z3ubHfddmQ9Znp4+cSeo0mQ2toSMvYYs6pezf3n5TDSgGhu1/9m7Yl8/mE7Tmsy/
qyQ1U2Gqv6LfOTMI1LoMl9wl6gQsTAEjsPpyqbgPlRSbfOyYBVwUQ/Q1u9oN961K
bndSr3ba/491WBKQ6AmMvSChuejvBrynqRpqLwmjPydgKJxASDAgtkrX4Ley39Xd
9/Gh983N0UTiw2j2fgsmHdzgYv7p1hRyXBh9D1c9SKM3fBL5VMbDddVpy8H+gVd1
4gCnT/dJwSGEuh4sR5Ev9yHrNeQjgtUNNoMOF5EUmOqRYnNZFgRx4DVskBUbhUa0
Q/cifR6wYitc3HXxtPUHOKsHNHFTqHgelsXZYmBYe/dGm2wsXjeya4DQYzY710Y1
2CIHeXburNuEhnW4V5qVvH+HV0Nc9+5IjH5TYNAH3bmaIF8TQ1/kgcr7m4FNSnJO
hjCdYNDM81djlFmCznrsN+eWGK4/+wMsRz+ZivXtWxozmPdAf1/4k9sBvzd+PQMx
bh0vhQZh665qPDDxk68m2SvpQsYRy2/nLhLW+VYEZ4PLVGwDHHnfoX4itEuA/dmu
+aAqfsjDhzhvutCJYLaOM/lz3ADdzVEuj9bKHkiLsclt5LRHoL+SlYTY+/lHpcU4
XvwyEF6O8CPxr0gp2oxMQWSj2gnSHrXWioaM0/9ouAkQla4xQWMStAJCbRyVFL0i
2LV2wTOFiux5y/8zKXDI7L9L9h96vWfVKXszFmSiG1WLETAY+8HQ1g37fUKG1kz7
ZCkQpUuveiRcRwDo4nnfLng14+8FpN1oM+b8H/rpx/oqfCJ5E2TiVq8IPuzrhrl0
o6UNxF+zFXi+w5KjjxIWRNHourpK698Ye71mFmjpZYi8zbId/Bvp0OIyzcQsHPQ1
Ot07R7d6n5Rt6B+rt3wFMsizyv5kISu2TAJFWfe56caP0j0N2HKX2hzHg0xSbXk8
pPUOOG7IprXMebptHAjMA44mL7+4Fdroj6RST+qLw+cYsqoKfoic1GZ6Dr7yiQ9P
XSjwKi1mhiwIKBKNrfMxWWqA7wRubq0KbJZlXtyvAr7lk+Wsa76rRxkGmv/fRF4U
aM0XzUT0nk5sj2gE8yQutt88CFdimTvGnsvRV/aEw1srdS7F2rG/H0NQvBCBmqCq
OjAwBYT1/bg0dWSX0Gqo9yTbZZAN/+hIvI2BLXct0bdAYkHJ70Z7mRP29S2tAdIh
kFfXpyLY3++5tHu4qSgzqZP9DAo6vDdn6hN3MeSX8Nycas5WdrxkQ5QqPGwUhu7V
2J0DtkeY/olM0ENMauTkizwsSYN1XXI1/f8EyIQRLI3ZNhOWQoDBxC2uGnBcaK+R
TPgK6Akmm60Yo8A2Wsf/NxtTpaf2dnaA7aBKCziFDBiJhVUthTtqvC183jQEpdC+
r0v6CXsvhkNRgHywqs3I1tcStLeoWoSznUG7WfOQ27gDURMa10js1QRTpkTr5hMp
ZzGGLWZgDG+Naycu4F8bGqWdLZfy8zf47MFWavqofVZF41FBnQ4d5PbtPWrBDDx4
+EE8Lkt7hDyrGp9de21rBaJQf0xPP7NqFNuNAgxfhHnWfj+1ldjvdSqE8+HYYsR4
T7SpiQxejou1HcRFeKkRMB5zcjDX6O2CFaev3GT/aaqFjD9L/sN50RlYqwj/9tEp
C/IGgsxQmdaBj22wCrdFEIuvm4ekBVA9B/O6g6wRJ1e7kQwNoPyPBvWn0c0XJP5V
Tz2wMJlD9DnUKZkuy2Wxbk1EXfUeIAlrZfzohxVA4rG6StpV3YTZ/MDyfbbLBcZN
gat1lo3YZxZwrBMxi1KEEnIZgSEO5OCWB+lMX3lvRJ279xd3pNFQs5DerKinSCRS
RUhF/YL/Get1esTCwA1XBhWWDloCZDuFPEzn7odfaLR1X9hjfa6aBo60as/yZs0q
fKFiGDQo5Id3SGqDwscC1Jz54JtctgjB50mmw/y8Rqk2SXMrerR47wXptn5bhGuW
SnwreyxE8PW9JuAjUEtJPiPVvIuV8EWrRPSCD3ca56eUXAj/uK77HPm/cYZmryAm
UA4spmAZVEqKNorzM2hGun/9lye4EDbGPsMBGCOUbo4gANLmZ4CdjVWGkwwkZJ6+
fdnUMOCrgPGh4KeoAXmCmadtBitN0icQi6zM+hwmL8SwnsSsIEtnhsNT0HJ0NuVa
sGhgqrId5JEml1ommZdbjp68QYBNq29yVAzjAETlPEazn49Go6IFCld1NhyPg98p
md/zgz5mVW1d7FS5RpoxdPK7GWBXLYqfzWwrQ2hYGjqrit0NFyc+tGkcinASc72E
UE5dLiO2fpCqTFElbE6mYxFihZv+lqwenZdfxq/C82eNZnZuQELrXWA7hi6rCluj
JNTNQYHHnVwu73+YBbiQr+vM80oSelqY4BGKLqfju6PX4vN/Kox4unpHRXACibWm
/kwuZ60Iyn3/e4Xdag+VS9/PXc+c6ejJIBY3abTGXCbuTCVMPLRz/Mv4qGlvG9Jp
mnHrbMVivKThPJBOdXSks+POJMsbxpqf6zEwirbWVgRZpN7ZOdDbYrZieqFcDzbQ
OHUPggGT0kxMVZi+lptcrCYv6MGVlQyJJqyBNKKqtCMd/3yqbl/1Sm0bc2AzlSBw
Wv0rgl3ebK8R+TSw85nJshTIS5VWf3web64KKXx22eLvo8PPegMljknq3ozalKzw
6JfiddcEokO4j0d0mepnjaHtfu4AFSENSz/qj3cuoho2WZxGaUHlM1saI2RWtfqA
5lXiQjwRX28Ls7QFg7aNK2OuBc/xERIR4XnPn2oX34yR4OVQ3zdCuZK4eAQm5h3+
k+0LjlP2CZHtIY7B14JjC/K996TBCHvrLhVifVApMVv6chG8SjBdU3vxVYbTGLrS
BlE9awqnod99yx2F2+yUTEYCaWwvXgz391bnPA7EY0MMkUCE6kTS8YdhMaL+shKR
3vuDwziBQ3EaOe7aJlcflRvAbRnCAGOL4xpAQETkmRLt+55QUT/KEHpn/FjM2pJe
OqWJXcQ7fnlq35f8hBJZ/8cec/LaJ1NgiAtDgIa7OtL7BD7BQBihAzEQe+8aG0ro
BYp1GUn6sEd0FWIRMm3e/j+M5hh8qvPF2M33WP1ulwfRfDXD2q5/kOKiUwRYKIRG
w8pywjsro9FhJMi61zV/sjk5azfg2kgS+1OyCNSL5WzixldLbMg9c5v7BRZsD7pv
0ETJFBWaQyOA/O/VUEumzmG9y5YjMjb+wmtQosWkRpecjYNaVv0ealbYUGP97EgB
wvwsijRmr+DRTYP6scncv8G1MZkb6lWB1RmkvIlaNT8MNGvfvUItdzW6azBEluki
WL5xmAaQFQ7xpF1oEXNSfDFl0PhoVe1ixMBOGAiMN158raogr+cpb6fZOao4ywD7
hoE0Umx5aefRiRiE7ePl4l2g/zDthfT+NSb5XWLnsBtSN2F5T3h/eWtrGBNTfo9J
Ppnh0HiHJUrPJa/f3KZbTS406PJv9lOAHMu/ENKiATPSb8oEsyQy0FHRtUAtHFS3
b79B/WGMMMYmjGWgz0NxGI7OP9N25KrSh0STqqsQSFux+AIxrvJaOlLXUTTf95R+
RoY5Wi8q57ivHKpcpjQ9LmR0QuPc8PT7T/0yYElKAt77WMfLMtGPuhL6K2Pzj9WB
vviu6tuIvqw7VCWePTG+n8ezk1O6sIVslcYzFNPSZg089KJMz9WsLlSB980Cnxsz
ZR2cwduGeJD4x87mkmRS58aI9QjNMqE671LCtci6ZygBy6gkUU7e6pVicwAJdFzS
QadA94+9XrlGrMB2jH0yAa+0ZLy2m/ygXqWjfYnCBuGWeVTye7uVq6+o65GS85+X
vLUjdAyR3wZPAIXS9yzYv6OBqydoJcfoVkNLKYf2mITZVQ5Ip0HXhAkMLjUzKEak
jObfExVMQPp1+UI59jh9unApXyE2gWbGu7A7mqJRe+rdC51s7kVDM5x2GVS40MKJ
Xy2r7Yex/2svB1bdyYl3e9smZPTPvV6wgOuJj6nizmexhDItdYvFbSfnQipiMwQT
PIDoAWLrF0suMd1SbYrDgYfnB2/G5/ttIQwUgLo6Q0cun3tODjDSfpIHWiwUVQrF
RWE/7yR4jlbMAGgMmaPnG66Zf2qn24KQWTpXChWUjccLWUkJ5nOs68SCuBhk789E
`protect END_PROTECTED
