`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGkPTdg+EbRKqCkI5LLW/U8Rn+ZrxALwZ87J0H/ojniGfqfu6IL7ExPIDjy+liF8
h5SlVhjZ7TsD7tjaYQxKH8gwKYZAjBG+MXWsEOOhxyFK6eV0V7ozo0IuOZvMg7l/
EASUpl9L67d8vOaNU4oY6j95lv0KrpKgaF4qG5D5Xk9CmS6OV5ZSqsFnGet9vTsZ
bQv8tJ3OpryQTWjvD84FLlXQHbMLrPIcXZwenVkgekwwkEfi70CyjRYJvUiNOdzy
n2315YqDtXcrTjxFCly8SQ==
`protect END_PROTECTED
