`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rkx1mTe50WR2sh3QOMmrDujESf5HXlzIS1frNm9fQm87fjUNop9QHe8ir5y6snr
XjTNe5JcasZuHSYUY7rNPK4SijEWOEdobkbFTQgLPqSJXrl0CyTU80nghkDH223G
np1+8f7SMM1ZvzsTLCyOwPT6gF+F20Mcjmz6gIChWPkvk9o3e+ncO1G1T6SrSIRw
lPgyp9NrCukluDaW+1XrtxBgFI8EnHlnubmkcqb/je/toLmn276VBDTu9RhPxWzD
SmMiYw9PEP4qpF2HwtDOTlBZvNsCvto1evMQPuWjl7e8rkbLN5zX8jEN2u3v9Iu4
IV4YAlxB8Y2OSLuhSJtpIx8jD8Zcnw176fTI464afkFFIM21iRbG1QI5Rhi0Z+pS
L1fnyYwI8SHwASgvTziU8or2OqbWuhDKBwwzs1lUfnWrTJyw0vWrsx3xY9/a9g8x
noJ3d/c8IBI+xjFNLqPFRbh+fEBC97MkKlxbOtbRAIu8O+/2/rJTjghlWoJNVjI4
VnYXbopo1jWmCsgnmjnjftv6NuubvKFOXIt7VXbxE1VcxBWana+xO53x1PD0m15i
KVRS0GITK3leYEHxQvNQT3fFYVT0x/kDnGHxDgATbmc84g3+Ig64tTFNKX1v0uCc
xVoLusyRKt9aiqhEO8j+WUfdzl3Y8gFxXcd3OA4GhvE=
`protect END_PROTECTED
