`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nV0TF3MDBBx5fiUzDb4OHZhcXeqCGHjlQbW/y3TVcf7TZoox0V+dBK63KSZCBMr
HLexl1FQh0V1iJkyfxQOFR8kvmzBqI5QGOwO1YmeWcATpfKbl3haJTbYQTMEFcRi
CssjDI22jy4kV0MLE/H0jwHWwzsZEs0v35ay5dIbd7RgOdWBoXcsbQzP5e2Yp1tH
fPMbi3hL073VEAkUTiqLvADYCQWtIwLDoOTwI0FGhfE6NvHce/jO6A2YKDhLipHJ
Fw1JMq6/c93Nq3ll5c/PPg==
`protect END_PROTECTED
