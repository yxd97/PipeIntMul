`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NTBdvBko72NOHnbXtvGiW77CNtr59InYOGLYmTsHDl7LcfhbNokbrRrH30bhuzrc
7py630+t01d3haItF4r2a1AaNRa2VPo0kJpn8Z+XOD9Yxd6h6Ym8AZkAXf7DPn/M
reQNU9LKAFVLcKB//DF1r71TPKWi2d2Djmo2x8NiVj5C3le6/eALeZpMPmOxgbRh
q4WkBiKz/TFlegXz07fSoItw/VJFvxxgvxI7MSpAUmtvto259uMYVd2GHGX1+uCp
c7470c9BPELAIXh4bwVbnYoFb/eskE7Dw6h9FswLs0vLorXImbdXLWT/mc3QAaZS
NjM+jdpnBniJpCLQ2gjcfXf2jEAH7UUl6x1jxwyq4SU+BGZo2wle5wRO/L7Je5Et
UoAWLsS4U4W3Fgf2+0MtvOQgv80ytUyOyx37xsf6qKloea6UMraLg5KwwZ6fbgSp
BxfuF7iAaOs7jDE5npdtLOe4YCDwmg5UtE15i5U4qmTTeh8E3schxh+SN0neBd2p
vV9ZC9SnxoO2mxPL5brnyqHIRAsftfnyoZJ8bjqcDW3xzTvmdJSdnmjm4CQy0qIW
kp782Zm93A6kLEjyus6i4CsSDAEiI+0q1kdP6WACqFwamrGlz742N3WPU47lckzl
CjI6T4DJ2Yyk/UKqnIjsMJzKlYsK6AWSJC8q3jSx0r/F6bQfTgKMQeng1uMktm2S
Ycd5OpBulHDH+PUEKlxYk4x9ERbPV8vcILE84IR83V3OCthRcVZUVTwjiIKb5pvK
eq3aAe3QkpfTSis5zGdbtBlZLSgohIbNSQq/Q0qc8fs1KoIQtE2u5qhj6d3niq1h
HtwNhz518k58mtF2Y+gCmjFx6l/bnh8Sp/Boyox20pybbvKeNuhgi7A5+QoOtdbV
Lx7xYiRUZT6ISEqwz5+x8IC3Odb0jPoECVbRBKOBUaonttXY+iUGOIP3mcrxvCFy
Q/+9lSlzxnnWrz4a0ngTyCVVnBVPJzzpkaa7C0Csi5CGJ1pY9ZrIxwNzoHLWScPx
xDowD85gp6uXsvb3ccfia6uLwYeKxOUbP4o5nSMYPYeCq0TBwvSawzON308HB/PI
8Lr/uYmtXddhzNJZ3W4xKIrKNREmS/6ERJDn+WNiQJi99eiltjHSLxOI28OzUu9k
JAbSN7eOKO96UtuO+dGkPAGg09NT5OyXNDCq7v5vVP8AR2LYNo+S+hzan5vyVbdT
vAvC3ainxzvFIcBlzhmMoVx63roarW1IdBFrR3JAdx7BOW6JwMFRtYkDVVIQcCy4
1hSvvEsJet7slbX1LXZ+9mt0m7lW0eMhqQkiUIbktp7UyVQrRRtMW6lG3/GUN1fQ
IcUqCeSmUtZeQQda6xRyGJyBTthewznqu1ouNfpN1EOnTwK7ZIuY1PjLAEesXSat
SVskjf2kGKJOLUEpXPMx3lW3MJa6d/IILnmbdlLuWaOBrixDX2TZJ2sB5vmb+0Oz
dP52OiV6OqoSbOADzuz7nBfgTsZX7xJu0nffKQFzzpV7pOpffV4aqf3nJoKbjbHk
oMIA5LXlLuxBhKv3YwNOx4ycuwIzFJpZFzcpQdGmIOn30AbXE1SdtrS9AM3RPcNl
/6wHQqPELCKXp3hv8XUClh4gpfsZQaQGSq80dfyZvUBDhibHabKisVkKSdaGAdwr
Q3vWig386pNABSgGZASB1SrmkSPBCaVqkKi3/hRjTl9/jT8CASzJD7QHNvv/UEFj
3Ntmghnsc6oN+ydazAXVTifoXX7bERpiNAcvNQOGeq2LsMT28tyWUfhI2ugwV82F
P4+54J4o0B0OwBqPMkPhT9qaI8kCLXdZLhBQXPddrGQFT2VO8UHLIBCPKuUbegtM
NQByRCecUTnih3woVsGmVHS1MN+LURM9X9+rpOSA39Baq2qbDjYmauEzd1lY3V24
PPMIg4NyEASoNl83KJ9BXnLCIBMr1lxO1WUP3qjY+rGrnHSP9qHU56EofTWz1Gh6
AWx3OMVDLAwLmtItXO9fk7JoSaIeP/y8pDIIO73n6f85/fmNIQxYaCgVKPPwV34H
yhYttw5fRpan8CyEQzmrHcIuzSKU77NZncKjWcZGUYP3aCbRzbcICYBqLCDJbhXV
v/Qu1qy7v/dywOPpIcYqyikxVYFqvTMVaeq86ZdJClG7hSnjVX7fmy2LyENmBab7
dFlgdFWjpnand65qQgPaarLpDMachHKdGCN1rne0cf81VBpMTzK2EfaFlL3lgUDt
88QgP2YiCc6QeKsMJ4KFB2Muz+puDqaU9T2hpFX+3+r9WG7Ve9IPzGkmo9pjexsK
8PG3YwfQPz4C2MISm45enJ1siyR2P/2g5RAbg/U4iXWuAuf0n32b6NzlBXmeHtrB
FKjEkGVYhi1xHUygtMbT74tw58gdp7/aA5X7u5k2g/bH7jb49UH3sxQ1IJMlDBNk
wfeBuAWpm/8k19nQw/Vh7OlzLjgcrtMhFnZNXrN66UxPL5DA9SE3iIyDtW9ayAW4
BN5gebKqp41XPlD+T3TkMEPFjHoHjySXGQs92hS0zEYKt2LBd4dQh7Bx7saLlJTn
RrW2KKiY/U2oA/z4T20HpQ+9cFlGG7WDgaXfM7Seq2UAYS2tR280bjKHvDj0IQG6
dKB6qpJA2f4xoMez1wVsClfgZHH84L91+D0NVEHaRXb+2gr3uLY1YTZDzVHs22FS
jJN2SFtSluHY/UREVeVa6+MWUg30/VbT386yZOMLwoOA5Fg2eWKboQS5zBXxpBXf
nR2HNKIrVnp7WJmlYG84B3iwIGMjLjy4OEpTT7y3U2NxNYktjMpWL9G9ek9nyeyL
`protect END_PROTECTED
