`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KzbeGGWbD30zPKPfooMoc0a6CLpaRZhXuKuDmByk4CAzHw/BDS165SCFsrFpyw/N
R/0GAcKacrsoH0GE1+ABVkUv6e7tWolWb7Gox4iCuE9sJHqa8mnbwqnZ4bk8XsBw
n6MjwCHcYPN6JVjLETS/vlUYo6i2uxtf9q+yCSZdQVvzuIXlVs6Q3moWPwCVY2a6
tLAD7lh3xIIM0ywiYahpA/fgrsDmMvq8Rh+ZCq9KrPbdXKSkrnTVdJ6td3h/TbMH
njZINJK+25ia5HsMmojk6/Mq5G2qI5q1BfQGsPV96kpeGNdw4DhFRtadsywuhg6g
ozIxe7puOYSpmBW5WHop095kX8lrrl9TxIvZ6rLQoavxlI30UC00cbqhBB2Yd9Nn
VL/N3t5+eJ8VwtxQLeQUMfJ4tmqbEFo6Wl7AWoh039J6wQ17yyjZn34l6gSCJ2SD
/5J2ZpLh+8FOhlOc3vdfZS7CA9jCwHu+19D+Ce+156VZiLveij0Sbqpnr81CiwYD
`protect END_PROTECTED
