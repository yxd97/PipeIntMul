`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SH2Nby1nVMgLTtLjtVt7YJ511M0VMFHhr2+FOD1nsdR/o/HHkki9cruob2RGksSE
lGODLt5ML0XX+LLAFiSw8s8nPnpMwHUStrZ4uczaiB48jatBxyPGzz6XVMHP3tJh
7LnJXUzIN6h2TgqKTt1lL3mU6cyWeiQ4q3ok2ilAHvuwPOjFrCG52EZ4NgQxEHD1
ChgOEMKCmxOxAiJnr+CYBx1owkSSZFcTFTHfjG4yQDsCTBRFwQvpxmBZrpIpz6QZ
qowhJC6ZeJB8x/5eQSwR0ligaZcjGw0flnpwE3y2MvI=
`protect END_PROTECTED
