`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JYzPGmMeotLBxGjskL+Ecf2+qPDw0DrYFbHGjedWgRmqbrx2Lj/rBvrhqJ+Gq7ae
UO0qBsbLqujVOKuIfpbWGWHhYVWu8dn4MM+8LLYaE8lLnwd72+u6F/D6tQu8E0Ww
/Y8ketytSazzKDDkTfSJY4kKHidseRaVvkVCBnByq74c8PTbQYZJjzxvy8+7C3Fz
WrNr1KNLvNnbYWIzmFORJkq/hzppY3GQP5XXCZ/YmQmg5ntCzAoZgeJB6PXx3iRN
LJJR6LNKP4wWLfvm7bIYx41Krx7Xac1xCIwY4orgIRkPuAflJNzEG2OLdaNZfPET
u4InhZC3majn77xeF5NQ/5YtZ/HX3g3ZJdtzMDRs0JNxEnO9tdctci636CTC5eCT
mC1B0LV/BJPMN7MBC4ON8o17kG+8aIxpyg+8lqYvIrbuEJ5jm/pIys2uf96NXkEv
eaW2AUso48I7zlsyBAoaU5P42uDJS8SORE2737fFBxJb9iSHr+Upif61qOa1uEkM
J+8Bw6577lXvAVgwOZ+34IaqpM+f2SJ3gjMVfPC0Y471EEOlTw7+ZFilsmfg4SZp
T/IL+rdab9FwGf6m89Qkv3XVo7X+oUytnz2HEmGC6QBDAiIviwZaxbbSpYmglnW5
qOdVhHsFfXOhn28QfgzfiFdU0A44HA7MHXDp1ahaBQVUBtL25owKt6/hfLutwcFQ
5nE0lItyAOBOBxnQ5q7GxzF/X/k5fYkva1JDftWcQQ7GlbKmD3R0pPU0AiiBZ1Xv
EkPEG/kv9UziDVaXZ2CoIw==
`protect END_PROTECTED
