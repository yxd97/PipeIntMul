`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JpMiuaFBofj6a04s84HAUYkSlhm0FKm6tAzP+j/Zvq5ltYd9mF7VDiP3FtxKaKgp
A8dItUwCSdKqM8uqsTsCDvV9mGPhHUsEY32Sk6YY0/J5sdbbVnVeyWUpCEyPweSR
2tRAZNLdrH/8HMjNY23YDtsa+QAm0g8WzEsOoivYNCvDrweonWw9MVotK34mbQ0d
wxmYQBzqjsPb9tDprBpWQdF0Q/E3VB3wcwTZZu7di4ewSD24NN5yMAK9JKvVS1HO
/5lRGNtb5FKXsqhX5ZKnRNfuNSDF5sDbrXXkc7n1i4yMS7np1eGC5hnibg8yVjKX
tEbmxACIyle9fzAjskl5ivsjKJGC4ft0g7nHopndrj5M3noVZJAfrW21T41G3D7t
v+551qy+TWlZ2yvOFrSIDDYxQBoI2sOzKgNfRNkjtMHGa82I9Zq2f44PSC8r04XX
oBNpUE7TbXppg2ErjxbWqq6ERXnoTOHxpAkpn8jvu8RGQ4u69H0sFDElUEognI/y
`protect END_PROTECTED
