`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UFwJvjp/CIqDnIe+Y7zyweK7MSGiFwTu59PyresJhbeJ4Lj7Z02BGjodEogXmvTe
hutz4Jo5+yiE53YDCvSmBcjUhhcVqjH5gOHqFRsWfzB9xoDlNICtvqRH1otZGyu3
51nrStX5mvApwZVKiSWmlntULhe+osck78pkzIfMxkGwoOOflZSOiYohPXroYMlX
CxkC3XEl2bibmG0KcDlR+JfP0DRs8rAJs5QYZXGNVCuhhO4TrFjSaa8kZ/thISzg
/znpr7PTGcDtAkedReWvFpOXIjrx/gJbPlStSMb48kDB/cS+qxeaTuaEKwWTSQFO
R0vTo3rmIARkk6jL+N+qY/x2hD4KwtkTlWIkabdOPtSVsOoNBebV2SwKU3RTyUE3
aQQwLUG6sR0zUhbRhJxr5Q==
`protect END_PROTECTED
