`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6zNaj1f2U9C97cd+OHY1mRILIiGZoe3rTgAI0ea/2EyJvRIH4XS6IpK799Kg5yiM
hL1p/GUbqezyruCI/W6xr2qouEc/tnQ96wnn1MopktYSrmGmU1hWBX3vrIlCa3jy
AuTBEfDiAAl5TTZfpmWEyx/wZsdovbUyscpTnLo6ihpX6zTGoTeXlMSrnyt0flHp
oVsjeNr0ePyZhnEnBiO1vwggadKCfBdmI6RsHAzwbk5yJfyRu6GEyWiz4l9Xh5xA
cb+2EO7Hy9/6iB9jZOTQ2V6WkyFvlLZU0OGUGpvdyp8WL/xuJT0+NgKa0nbuJ/xY
XNjb2YaVzjlTyf+4g3cG9m/sWpobY8gXgpro/jIlBvIZ1Kp6r7LEzxt+trVL4so3
xWCbq4TZuw+w94RZzSMNnuKZqkkc5tN7xwgWdHRWAxitrmuanHeuCEEx4BY90IeL
gGR6N0WaAxinHN1C/91YR7wB6Zb+C1GdMdXgWaQhJCfgicVdgi0Zh4RX5E9jsWEs
ReP7ZsLO3FAfdyGz/A5LVgIVw0UXYHZaOVt7YasHeSuRcSjhmLABwLsEwJ+2ezex
aewTCRpVCGQydfP+4PN5bbgk76DFOBEF3DkQ1U4V+X+XjaZ+gBl/PlFp8ptVx/4A
JXBY7VBb7nTknbE6sV6gQN18cbZB9+dCir/WKrZfre7SQHmndfa/NF4vBU0TU/hU
QFgZP9nyOxEhgyuT1NTbj7lZDsH8UbQia3dOKRosrAeoa+xEJL2tzWs+w3WhLv5d
+XB+B08Iae1piXFZkFLLQWaqKk1+jP45vGHqAMFDlbAUDn6TrUiMmK1t+A5P4phk
kV8O6KVcrfw4mGAXOcx17lnVMXmX2jXuzU7xzuWPovIeZ+23q8Q4dJfBE7LdFJXj
2k6YCYTBkQ5lrEDQy3Qi0Q==
`protect END_PROTECTED
