`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4CNEEDTOlx8vnCBORTzT7FB+oNsg0UKUylELWb5l/dISzNV1vwauset3qe0pW5d5
GbC6ldXRdXZ9og3TbKNLqOcrddDHCfpj+o50w8FeZ9cviT4dWtLzs2PsCAeZFeQo
qKOVjAW62fT2XboNoPwxVGwvwdptCwg8wZAkY3Y0+gAaStcb0+jeQVN4fLi3o2zg
sJG7+QkdSYu7nKg/ufU1nAmX/Jq7Ps8eaOC30NoWnzoXcnauo0d4TKtlSF50xccb
mebnQL0FOBm4WAYxaMbp+HHXvd3ulMOGb54MZI7N2spJj2Sy8X2g02lkWOyGNZqU
7bsUpcPgltK6EHQKSXkeVgj+RyAOoGc4o8yvKgSvvJFoEjMbv4WVLrG9el4IBj/A
aPWkcBMqFvJpxmr5821l0EvHxz6iXxFGPbwODiBzhU9K9IPO0+f29lfsuOnwnLVE
FF5FA1wgthf91BM0ZsEk30NLYiVvZREyoRv2RuTr1otuGM5H9jkJElBEtrcEwus8
zQ2tYq6ChD8EXbJuKo32aNbdr2bSmXs5F1K4q5OyGio7C0rsyucUhqbSp+1tDbbm
nJ+/Eu7ErL8R1BYhtUIERcfFQ1fodi6a0RG1A7KHNnV0ya5zHsxK9dp7iuS4q36l
RleXtNn9e4bmfcdAIQWM6VJSQi779Bx+WoXQkpE/WcI9NSottwGUFX12l9xvs4F3
HkM7lj5Zsfwmf+JgZYxvMUp8u/dKKLxUs3WyomyYIsiroaPQMRkmGxTKui9l4IgD
RTGziiTjcaVK7SqgXWKhLF1Yg1F9ROp6hkOKcuHtaec=
`protect END_PROTECTED
