`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mWfWayDCO6XOHuOmKlirUBMA7pmH1GrxiXW+vbSmqaMxbgl+RmkKscXkenLYbkas
b7mmRxWIiS29rXR3gPPg2G6JId+3OJj88ZDRDucrkoHgWCjtwTg+3/lF9R0h4L8t
kBtmyzJV3SLdsVIB+vclQZq/OdkxU1CvCycK1J7lrDR/Kj7SjurHU/iAowvfYtFm
PduZTVdFl0IyXqoWLw5x//OhsGzykQUoRbSnV1REuOdcRzlwPR8/zSiW1hfbJ9KJ
x6VPtC68l4P7EIQhwD6ykOPaFjvW21kBrch8mG2tpVxv1YXUsKUKGZt/5hvvvPV9
4p+2A/apwmQXBtDdKFpcZgAoKpdsVJtgnyt/ifV9cJ0XjM7jjGHaP7+z0ozcgpkQ
bs0rZmQD3P2uTGnFh9JdaGWC5p8+MHXT4e6v2Ym7hDrDKLYS0UWGIn6IlzdtKH6C
ME54FBqJU3xzDoVk/tI8LkOJ1kB44hok2+XwDjBd0ehe3e38T1EnphRxqdQruOQX
5jcG/l6r0LZeAZzXzNfP3tumt2pORq+85tQsH+YKke4g2YLES26krs9Ep8fdHSpF
pNJS0Mrhunuh3EKDP4cK/38CaLlzsrZSM+k0mTVkZ3d653cQLC31z8bu+1TOvJFk
l2l1Z6dQCZFgTFyA9/XuxXcaUmsYuwd/yAOQwwfEXDFIg4hEMJBHAdit8YdbhaDR
yDmHcvN2Xc310tUDmjMPNVTIYiRbR425IM5p4GDD4zthcNpo9jZTRF4f12cqE+nT
aGs3dY+b2TdC4k29g3oeC9tjwT/zqegov3M9ujl8bIrQm8MuUc2U41aZJNUkbZcI
0TiLIZXOnm98NIij+Z354oXZDX3c8+9Np81DD8QeRle4fhghqZLHnGwascL541o1
7NmVnTK8VehrvmpKKAmDZV61br1DIV8hTe+wShFPZDGTW5xCScbziTjxw6qI0BID
R6ZHvmdIxtILwsZyE3hMsgwLm/K2HNkcPNH/xbnf+LPnALEkBRRQULuULhgQPDuh
hs05ACQ9rX8rBRJanFj7c7HXscDQ88EvuoERYKw4GMi7+coMuq/KswK4OkJBOiZH
AuCfcLwrlg0Jec9OvOh56Ej++XcQVrP+cSo/pNXlv3R2dJHkUG4LbE+VIBk4N1+J
uHrGP73cb8ginSlsbRuWVBvgfoQgGUzZWyiC1Ao9E1c4oA2193ERpFke1a4o3OQy
ecg3izmRPxjNU/GYfBbjT4yngE4Z6uraixE5Upajygk+hZ3a/fmhpp1K8AuV+kMz
Hou6plOsE3TCouJhMa7qniOjFHmfiK34rQaKuG8RJCzjk8BFHC1ncZCFlRfMrRR2
Xmxm6fdUyKoIdlmOx09npXfJsEplTMoQAPhcFCbw6rIWzp2QdVKs85iPPxRlAMSm
Sq4yconYma7XNhYw6+Pr1guOSVz9xFVzgU7oVzv8GEKNthoDaCWfm9C6eEI4vN41
/M0yysEOxeJPGgYduJ2tPknSPY+wquEi7R2SnkuzU1zpVjAnI+ERscSYeE55F5jK
K2KjolIt0t42U/e202qGoCDfZexsYV8+GvL1PVTeISGwrdoi0WLZKT1sLBoLXB0Z
gtOe+Oj7zhlf9LjnWjmdBi3uYBY/tGk3pfhm6ljzAQ3BVwZwa1b0TrhRgVKbU8CE
1OXFM6UxEpU3v3/U/M/k0A==
`protect END_PROTECTED
