`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GtHMb61JTBAwut6TH/aKcBDw3HoscaQA/WQ0xcjtnj13pc1oLyT6dWm5A3J1PM0c
LOKZECqWaCD0D52l8+YV0X6OYm2CqIGoDA0UEjUtR6khloHX1jEs9aDC4KYiWb6j
hv+IZYu4rQaX2cu/P0YOdHtnN7rMGuJyUsUdDkXNljWYCgmw8Z7Bdjw55Kd58/rw
fYkHMQ55FVprfhjRPa/7NkHKey7JCq7YMk6yHYqdtGiNzBAAZYD4GC7YOlXNHg3d
hVR9qLFAu78KK7W5HWavCO3VRFsZ1n9UM2rIcgVFPOr8XezIP+uYN3k0dFG2e/H3
rV98y8uGxHkA7o/k/GjUvk142WfQ4YXGanARzUaokYXp6dN/qmgZmi/96n+19cSH
o8nD/eK4Y7EyxSKXg1r7TuWyCJgi+trJNYjvVEXGCpQ9dRb2nFG6SKOOIv8ysdzW
mF4j5UHMJV6IGyD/0bzSpY9tMxmi7Qy+WFC2nJWdjK5JdpfM5A5Q5gsBWMHx9X9b
OFRw4wuyWYshBr2S4Oo34EW4FT4t0GpGmvHpCAOIGXFD9d6jJAxHlzTVm8lwRchr
Iu5ORXBI3ULEKf+Ou1zbvYyN0oQrTsliJ2u1FM8l+BEURzIqrN71I6dhrwlluIiT
spM9Y3i0JbGi6Xi3k4aspqyZTF0S16tfZG49Iz4L7x2xCaRAAZStU4xJDEhyPZqd
264ZDNTE3GYNeCpVaudUg/JV3OVY3bdVZ0X2TMxUZVYTLVL2v3dRn3jX4lZdPCl/
NcumLq3FdZDtccNFw5LqyhGCp0ckUJybVxD04jqBaGXe3ozalQXBY0WaojS9OLWd
Xid1InZ3DQUeVfEEDPw1Q8Q/kOT9dehKmjmnr8xfWHhfQCy/zVZKYW9hzvVaQL4R
+UFXoPyibY1PesgW0LvpT5RFD6eejjA/jiLNP+xAFaMz0YB15jIJm7SrXIe+Qh26
fT5M/ivRuSVCQZJW9byBVXnJuiqNjcB3M73yw10rSQD/pCT+wWFPvI76q9PR2FiA
VyhW/Akr9UwoMy7e1GkYXTkTZJ0aXApFrYjbe8zowZegb6Xjco08oPSmAOxZwXwO
jLQZ6PtE9UvEDBy/7+swfQ==
`protect END_PROTECTED
