`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrePvmgyge9zPnY06GtMWeOAqvH3dChnjl9REMqy1/nRqELA6Q1CYrf0OG6RYEmG
bY4ZDaEGFyHG0x1ziFeJQSGXmBlPCmN7Z5IOMIxtw078gke2RwiPBIuNIgl1Z3On
9D1tHsVdSaDHVIL2p6BcOnyyXD1+zVy+V1aAxMbVlm7MTr5a2BYmKYK06Vld5w+b
Gc1JPXkHxU/7Gx/L95D5HC9HDf3/KoFziWxLH4/Z8w+ntcXz1mxlfZQPHnOfWUn8
ZKCxBbO8JJJMBACugPN3cyi2pVdX7iEygaJFWvi+dbbd7yN/PpPKn9IQWhxKhzBT
NGkT5YpCthv0NdTjRlUTivQ8n57M0nZNN8t0yI2SG7ER+Wemstg4RwGSg70ZL3po
0IjM6f2J4FN967jmaA5VJMIKQgmif8cVTUu8otBzJI0CjmUa3foJr3eohPbvXjkO
wNHXmpX6jbO7SPE8QMCaXWn0Zd77epulEmUaSG1Uc2znFpNhIps+KUHGCSqlyj5d
KZFPQ1lKJprXBK3+uPzkPdqXQumtm11ASgTaC95nyg62GizsfsgD8BZCkBva30RT
Iqm7mxdPIOQf1sT4V8jzisoFCqN1yJLo8AH72z1OkkOjUIgIXzMCVlUMam/Hxkjd
xqe3Km3ehrn3BBrMGmjn0JrMHdOmT+9z1msp3+AHrrrxqG0CYy5PPbIiSvt4/vE3
iWyVriZrroq5gWz7h0J1QQU+3HZOxtqfPyeiaGSqJz79qRMtYCSns+xWen3IPjJD
98g0wtqyQGPBJfmlDOZamFFjb7sojLCb2VTXcA4vm2QWSjWsjjtz/dvrigObdhwg
f2k/v/lHjbGZ9g0u7to+qGkibR6IQEkcPZ/w9wad8dupCHOwBP3ZVRlFEn52CWlz
8J9PHDfyfgNVnDXAIjBkh4Ma4B/bDWhfJS4cAHBdR5YQ4+75FUNiTXau0TGh5VTO
uY/NyJKUaGFRXZF/R1cUkmwqEGDPhoUau0UTOyemtd+z73jOcUhyvlEOi0goUbAS
apMwDrcuLZICQqChgg8xkMv5aHFhrA/zMpKYPo0t+ARxf9k4iy3z2wJzedZClQ/P
Kc032JYn4Q6XUi5FymOT6UTaCe50Kmpsrj9NyvKL11zjTxVmeKbCwMx2TuP/9zEU
mWOlmFW1q6rpwnVQONW2Z2oYtvT/0aH4EHKDnX9KtngZ8iPHiQPpEsoHnRnPOTV0
/3wIZZ3x4DlfR3Uw0mdQGZYsflLNeTgpKK8S9qoB1nl2CqMLBWQoGQ/vU4EwObou
4I5vmkI+fpCFh7oVvS+3gJkZ/AjTZsIuJDgfyGHg3IywvnpdHHEeOaSey+ILf68q
tAkXMrUEYVYQM1eYfX4ayr2rXGYdo9Siaopl63OnZ1XCAijDtV8Lp0Gx1IW1/Pyq
JldiW/PSAYyFGT80LFf9X+NwBnBtmCJkox/f/58LqKCWprXYx+n/3xZEreqaiHXJ
54gjGwnjh6dcVfur6xSNUrUoaKAedpsTKLsyV3/Vkka2UQr3dxg/vDxWjpfjokMJ
7dBfOeBvKFow75VdBtVGCv7dJ9ReUoq1Fr81Nx/+SVkLrrEEOjV5n1wU9J0ztTEf
P7Han7xW4DUqz7rqH3o/ojG4iXLDnj497tD6DVSOO2yvV0uAhf8aEvib0pmRuA+5
lyCzvGDIDP1TAfeb9HblpE0gPqNf++cPf66H+/wzJ88Dv7qYTZsToD4LUg6Zjf2p
uezCa7dpBPiIVKumdZZBiBtdZteTTC867VHAqFXmjA41r4sjCUHVqas05HmtvO4H
+28fpeY4SJ9x1iuQKq6qXfIwAWYXDPPwGHC/k9OJ5LBfPzzC9TgolFdYjjs2ex5T
D06os+wVgMyuPk7iyeL9WnKt6uKaD2Ihs1Px44D1len8yAq0ag2uGkw8sHPxgdpX
5zbh1zSpPhSbFz0KbSQhKZLzgi64ATtibypAfZtQAcYgzFIHbFvVqVC0wzqqjQQt
nPftPFlk9cBTym+/gvEE66paFa9aZpFdawfX4k2DenhFuMBJgn97CmnX2kGEBpga
rXa9jDUzvX5n9Z51GrUN1IxrrxR/3ydw9fIe+HPYTi9HdfPB0gMiqepiBXGrqPRm
aXEK1/UrDi0qn0P2icDFF1jZvdvHha5emmTopxC6zQi85rmRx+lrKSnwEtvZ+LSa
JMSSXPBihJH9U/18GfNSOFx3AdN5ipRyqJLLmbl1VHUJW/yGzDHWROkW0/a0QNBO
pnfrD6J0JBVtKF+W/ZREZ3xIQcKhQt9Wm8vrdwBlvPeVsGBOhzdJDiM/N4CybDR1
8iIZp1p8AQgFr1Kn/EC0dxtvHJSntp6Ew/EaYsGr2fnKm6lvg5HvqJ7KCvJzSwDM
kVIudxZdGdirax/rVfucQMoVBoJ9F/quC6uLdihD8kkzaDZ0A/yL/rOVsz9v/qI4
Z/QhoobpbdDZnZyGfvBPyliapnMzYRZ2SAFc07u5LkVb3uw0BAjKxWnqlQVpGnir
wWde9Zsaid5O6xiGXV/6SwegX9WrMiwkjtLGqpgx6vihhX9s5o8dkwMpVh/oJvyo
U8UoCqtNrAKfqKYSSYtTvdx6AB5vq4cNYzNZY2xIJBc8dHUNtZL//4FgkMuLjtPP
gLv6mqHxX079rYcanJdLdVQSwaMNLttxppOSwhhjNfZMYuswYfEmVczP+Ll5BJyV
cwyvAbOzqhqSIxXAE/SiZpDG8o/8aq5U9LwwXKWdfd98GCnNst7ckOvqTHqYmK8M
`protect END_PROTECTED
