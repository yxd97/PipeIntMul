`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+KcE3gDK6bB11P6mAKeG9Jvom5DXNEuxptUPxaTw7OtH9Wj6q5IFsbysuujj5R+
AzTaaKNkzfWMvRCuCiiqI3sc3piGHZov/nAw1i6Lfutp4923F7+doQSuVxtymH4A
JUlEq6r8y//dMnL7QuCukuWpnkEeI8vrZ+hglaZgKdKnIC+2ZmEmb9Q5dyQe+stE
tFsvnSvj5IrFvqMdxshd0iS27jJb/X4exFWB9GGgGdXqk8YR7ZvfsBWhBOga8l//
FjgHbuxXgHa5t4iTiY8OgrmQ6VXi9/p0vJNLCyLy+W0BKlarXKckiFi/BtYezBVa
TyWaruHJNqQIlxm+rsPlGx/c/PtBX0HKnQ1Qvv+jTJdXuwmN64s1S5iAB/YKVmZT
G76b1HArB3kbtrlFaI/aPetSrg6wN8XJGJyfF/zMFr22wz574BGIoj6WVAVx6S3e
cjmoBqrawn/DktHt98SEDmeuoh51j6ZsS2HY7qH6XeAfNOGIWgIm3e+NpV5Hi8+N
EcxCGgh0Ug/A5JEC5A3gD82m9G8m4m6CXIBFf81mRbkcZPUbGzeB6TEnra98yeg5
`protect END_PROTECTED
