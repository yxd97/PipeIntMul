`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdJVeu92hCBwUoLA9Dj7mZgqdJL0/3IY1RFIwUTLq1krOP/Ua4fPEbA4fRVKc7PU
gFxtxBCqc2CYdqAv/wTivMDZNpLn8VrGG/BDsYdllSBuMBF+pJHTyOMGxuvZYO1E
Kn7koArn6q3XE7qb+e+q1m/t5LDK2PuGlsDNjJzybJegvtKzhY2XTSx2R6uLYu2R
hm6Jp9v8ajT4f8zYxtXamTBv01i4zwZOh/lelo6LLF52Axtn7pLDptod3rKRHl1M
gUaHAbeS6GybehuAUvjqjI0a39U/ypy5JDUsPhMTAcD0ZTE9J6Ca+vJX7YsXUmqd
fk63vfilbxIwHcg33EIL9Q==
`protect END_PROTECTED
