`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmuRXMY28qQ0HqlOa57XB8yLPDURlINUJm9P+6qqd4mpxv+55cxqv6jJ7v9M8eAm
dX2s3EsiuSAv9X92JwpGnN8avgswfXvgIVtVXA16O+THszSrvhvBBrwg47bgzbUy
Kr3CajCNoR1wau5gBmYPgAl/mx1KNX/mpwbXTZ3Or6DB6TDc4feKlpVE1oII7rbH
dcoKC2nUKDACjgN4PCVGZ9W7baOrtBDrSTemqBOUEUQinGHnxQruKdHj7k6aEXll
sU/dwboSRxlmnUzWK5Y4rLWi+IxYVLlYufObk4zLmJanF7dQxXk9gBqMS912qZXB
IIJY0DdzmiDbN1b7oA5XCqicfFEclzfLLNme+P2qIuCfM2P/7DU9fohEzrBWQCP6
yYWjYnblGz27+XobkLAptkEBFczNXz8mAeASbNagYNxVCKvflnpUYcUQ8a9vAO7y
vxKQ4tsKuverG42hrpgCbEKlNK1tEl3Jmpn8rwnUZKIbIQiWH4oDNLdlngKg0FdZ
KzdhifjhICIG55WPPqeGdDAQzbneMYDV9BWNIqs8trFmcxLRHuqXFLtP1V37R17c
4BRx78FfIbRJgaoBp84KyAM3C0zcXa877epOgZU8mbU=
`protect END_PROTECTED
