`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tv6ZgpxQhP0Lc4CRuQmx9gkQft6VQh+bcY0L0L2FVXfBta2dDV1KYpB9cLf2cn4J
hxczaIqEVYUjDp36+MGt8Mf0zkeLbSv/OyZZpOkIDlhmB6fuUb3IM97aoaz3GtW6
GPh/xd7DVSVC5DRVQ2T/MFbrwwWVrQq6nSZ6ZIrbmCv8bnE3Mw/nzROkkKtwVq8n
vW0TV1liy1Y2bQ+YpwxUA5ds62lq/bFC4QIR1AT3roPPtoHzAoLHCoe+QG8dm4B7
E2ejabu8CtPmBdq53X61FnpwMld0YmQtW0u7KJp8b6TLo7bGVKQpRTqLgGnyJJDZ
tqgPRLXSuuTeMIvnAjvaKQ==
`protect END_PROTECTED
