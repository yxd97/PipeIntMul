`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbuTjRBGuSNEinIZ+XxKOu54lGSWvcZIlKGi7yQeoFXtWiwVG04WC4EPlwfc+g9R
7/CKC4NstsdPvfepGVk3p9YFkcXqi54gm+iaLEuNaN/wAZztxmPoIeKLAmV4mFx3
tRzLVYRNwOW2Q83TA7OdYeboQao0WBeg4Z3ZNlr3SQic/JOVpraLIlkH7zDoSHlM
Moj8ChZG2kgYjpBqwxJa2CKeggCjiDHVcUeffBj5notdwPZzt3ENysSod1owBZpM
hh89WCWMZ9ZzqE7/GYwzAGBG32a5fdN8cLC1hO4dQ4O+kpMd0mnWxvDUvt6OS2Ar
9kN/4lpo71PtZyiIi4x3bSmmn31r8IfCSTJ950792rjMtqhSzlpjkw4BZJwQxK7M
PlpRIgP3JjL6/92279BJH5NR53/NCEHLXp7xHpr3x4ar7o0sT6YMeifNx6RlxmV3
ph+pmTvhcswiZO5Nq6vlI4UNpd8UCw7u7VthiTG9L6UBxlj9ACuAfgWPoHFPDOoa
+nBTVSxUW6rsW1csbu18iewXV5SmDT3Qrwb17P8O1aiRlNu+4bvZZy70ZHkMQPs+
lQCR0YAYNz082xfmpIFGZvYESQ+gpUG/SCmCweRctktMcCuslervs3/9C5kp2z2N
lPQ+r3Q3en5ZayiWi+k7OEzKpv4o/pZnsrnF9hadRsdQRBS08YReH8XjEqxi87pC
S+m4aVRVBTSDJBX3ckqbSJhEqJ1Kp52FHUqXnlznuG0ZudM513hqqBEFcc9mN3ri
EQ8mineqXp+hPK5qLmaaOQURUc2eZJULbag0/xAKTPk+ejpucWVjgrD/727gmrm1
rqWMX8BJ8qhjGteW4dhYU1QbW2suiOUxxZJq7Z/jHNB11bU1Ml3+wK6HUeZ71LlN
Whl5SKMlLQPDULKOgJCRC9SJV+Z4RuH3dZjip74YerM+D+FqxvEiiJD0FrM+s67k
HP/MbFiP15YKpg8gBB1GqyuY0adjR7wZurWDfwrVwYZVOASIZPTACral2yi1mdvb
orJUQBJOJhXfMyS3bufiPOmop9UkJy8eRyYJ75b9p2p5LKEhZ6Vh7EenZjF/aaA+
JYz2/gJ0ERznrUsX/k+A+/IHOIbTY8QNz4Dd/iem/ZyuY/9EspN9uV+V4iy9Mz71
Wz+ZbremkE2YtKw3x+xZYrYr7sv2Ru+K2f8nD0bo6XcGQpjaIxf/3bnLNk4vsf8L
ZylsfgX3EzgoBNHHbSl4cRqJiKcmCQAVLBEHJked8pDhBvPoRBTvdd9FEidh/hbG
2hPsxaQrjum/4kCJLs5hezPAloPguCrteQg2QUu/XXa83QfTt/azfPG0wSvrf/8G
GrzBhpa/BS0V9g28LZ0TUoWQkfiYow9JzyQ9mKXpHV86LlbkQhm6I23GKGH5AAae
3rXfzyKn8UE5PvJUOc9LOojBgctX+iWeuyeGfYCLgPveuDQblXBgZqNLUgM1AddM
`protect END_PROTECTED
