`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MWdDRwE/v5SOcAwftHoW/e8LXZSwUbt3i7GYkTcOUzPdCaSEFtajd12eHefI9qgU
5zqUjRwY3gHftVaA44SzREUg2i/RrVBcY+C/Qv61XbRiEP+3WNskPj+9mCVAfzqv
CiNEdCY2pM8Vp2jTj3W/cbwcw/Wz7fzoNQ61XWtoR3WjMZECTwYVRZxdYdaFIVYl
gLkEBc8cIG+gFF6K7QllocH/Aft9wGTAX9/iYvZtuGzZhpsXko6jiOVgltvaKmau
KrPYbGTy6hRR8OkwaJ3Vt87Zbk+b+8PnZeZya+foN6aFlYuHXqG5CxT8GdeN1bRP
9XyBICMqnxIfb3DDn3Ri4ob67zjxHMZ0BHsNqj2zNfbKL/mwhr9U6NWNKqAPME4x
enVFiJ6U9Ziw6K37dAFM5/w5a4pIhV50impSPOBaGAMoFNF6jtpP13SYmiZO1Rkm
wpUa6n20UI2W1qV3vP+aM5FTEZro1QplC0RLNoXrupLzsUxASEjAi7ucfH5Vyit0
wTi7X+be4KRXFNu79U8IfsHIhvbWMAUz1OaUNbkyFd3j6MBc9Gbnz+9SjO9PCdIz
B3JmMXj3NE61I/FDr2SXD+IHVsiYib96uynNvQKwjOG+4MPQ2bhyJYSI1kVfhM8w
tQGihE9ym5U3SMBu75psgtRXnVv0WJa1RwyftvYW9c87aMqMCNI/P8klALyelTYk
sXZ6pVB74QRK1froIK9lLlY/CXdsv+LPbTAHCOHFXFe1Rl+/yavvVF0IkpEmC/3N
Q5b4dqzHuDwHpeq8a2dK0TZqqT0WFNr/9CeBSMsdZCx7+xCd/NXPr7WS3SwfF+FL
WwqQG8huxrbBoz5yf2aCl0e8dQnJL60HRzLcfMqK0rKfrxJJp2BzGKA+ZXWlyD8z
ssRo7h7puIOiPi4fq5JzCg==
`protect END_PROTECTED
