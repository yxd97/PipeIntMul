`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XBRyFW8OlvsgHk5R3ncjZMG9/5+bvz48DKHl1X6akSa4uk0ShV5oBkkTya+bSWee
Y7wKZ4W24qrokN+Mx8Xqd7k4BBXHZDlmwe0QOW8GSgXTUxZJav4BTwcGzdiAL8Pu
o63OXRvdoPGQg7bLCi6cHDN1+c/2vYmGMWsaTZltPaE2pfGCFghAwamwS5VK+QmC
FHcTyzHIXjCvN1DI6faDrmR3Eb9mmyhwdG71rKibCG6nbCKz055zbNkOiSkBSu+H
03TuQuHOn9/pHwLTUhl2q0Z7k+wsJ4phnvu/MB0vkVyMsDKdR0ktE79+64J3C0GA
MrChMPWASJQ7swAWEUDVnnsxPzV0+lLM+ne2v9LUVJTdc/UMMZdxAWTORV494HOt
8W7D3kIouftuXaBiAOJgpi0bt1xId+a67bj6QcqtlSig9D4sfNd/x383MrbnC894
g59M9IA2WPyalJkYRVNTVE+yYpgfPpuFgznPdPpmf8fhWVEBkey1ZViAhugXa9pG
NgG3lrH1R2mEjv05UJpv6eCH7SZv5YmW/XWizw0SSwgqEfEI6oiJP7XX/1cIWO54
wWvElbSBXEguK1TRJobrjyFfird+dDDaVRtbJ9QXHV/2lv+t9wo+zheja2P7npwE
iE9zeHoShKe+BTW6sJLvcMOFNPYerdJPcjcuomWceksXacy29tHj73qSrMKsLvvN
`protect END_PROTECTED
