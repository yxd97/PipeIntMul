`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sSywnGFAJPmotluGD1y9uyYUZ5kyXdfAjCp4ssIGvRP5DwPXlCLppAHlQS6Q+f4T
PZx9cnqSTe6NewT37Zr4uKZRDD3XQDD2bFW4Hi38KdwQvSjk1BCyrQOTJQBuKam+
XTICE9TFeBS/bxh9JkTb7eL9ToJzPyc1eHTbI1wrZnZ1G9qXnZjWYOtOYZ6tsqQu
JQUipxLnTjNjKnuJC9MWWnGe6s5bv0Q5gV7+dsusj35D63I7rS6P/LkgTg6XJSLf
RwHMFY7rYdbeE4D4cjgI5SRBTT0QjSQz+7wwnGWV8koVe1CQJBvUPN98+qYyDx50
TXTZYGxYh2zuSnrcqYW46L0QpL4o+Wdp9mA+rqudCLNmk9JZJQqpU10aQgmoGy2C
h7pDZb3Z6meziaULWvZdlHO+VoFSPGiPMMkHbQo9o51uGs+4+gBVzxn3DXYk71n+
0d7D9OPxZlRsbq18QfdMN2alotH5KVjH4yMH0u6iFGYBfmpmihCoLzaHw8a2/U54
7OOQaNrYx2GLHAa92I+8JEPiSUB8EJdYqr5BUURTTuba1v8sbedrH76Fw8B0mf4f
85UdIu0TMIZmrfAd8ohyOQ==
`protect END_PROTECTED
