`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
reAWiVyp/0TcpM8uoiWt/y2veTdCZkBApKXn+gjyL9/b74W4tNI563yOWrCF4uNb
8a4U9HiOEUqKPjwvSg1JDX1HGBxl3cDwYEuD0Oumjw1a6WAJg1L6KOAj9mm/XGOr
2rU79veyAdVaINsJKJHhKPGuOkOEcMTlMVp2qS83kJP/xwf03bWQv+WYPDUSz94T
ZXpIzWZ8CbXa1+SymMk9AmGbzEOZVPyOd5WQhYdDrL4WF3w2gtNrW0lfmt4xd+D8
ZrcYanE7NrAyDcDIqkrJ7XjLBRxVah5Cgpumye6MYj9/UD+l0alhy8+T281Qc2MC
9oR7P334Pn0OqcChYxXlMBJXoH7MnP/TStVCFLrYm/ftmRczoef0zl6jUk4tjARN
3L1jtt9AynL83zVs+v0TldMB1nTnaP2rAuNIDXePTTKaLyV1e5061OB0ViFQJHNp
baMKha47sZ08AYSQb1OmFRK3fwhgBMgzSWJmQYOYQPdpAommMid6C7s1pSM6OVsf
`protect END_PROTECTED
