`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hF9uptiAhMvfcIVZ++Z5Zgr9Nb60mAWMa85ZJA1FVuGovAws2P4bsUA23PBKCDNU
csu8m0dVyhPUcDxo6xUnEGfRsmJ7u0lfbOBwfBTjpvBkH7L7WTuQhFx+PUmWhB4E
PyBdDdYf856h22w0yAYuL7s/tYSkxSi7gZtkSWT9Ok2SbxA15kMqO1N6Hu58YR/v
E6zaFZvkTqsA7OJxnd99qOgBZcKQDh9O8Nv7Gh0OTN3kUai7Dv1ZkSFQ/LuuiUoC
PgPiGszWxuxyJlxodxbhKlG8RyKBBfFGYgSIm7XC5v8Nzxst84qu+1Kt/PfKAbax
HSX3paftHnJGzkukWnbjTc4xOIGDTR9PsbUu7YR2RDf1HjpnKxj4DmmprAHGhpxA
MhFsP+0zyrdpx4A4Pkn4vnG8bDpisMJuQuQUefG0KyVMQaA0Nsydfh1zVB0WLR7S
4CXbq4DQxo8VqFG/p0Vh+ghpTnDdMIBzcCMTzqEYe/Y9v3+cakREKHvU93QCiX6p
VoLwd7VZ6wXrV0Rsb8TK08Km+2jyFW+Obu9YRnTRAr/+FIpe99c56JBAuIlAeqaI
0xFg8pf2Ed5Sh/YkQwxJQB5DRqAIvl3mKwT7gh7hEciyWUqvkNirLPxx5jIm1vcf
mDN0P3d9qdXVCRMzOKBusOi5oqsWG5BoNT86TNCnvLXOZtxBdKZZU1hjqBg2E0zf
51n3nzyZ2Qo0EfModXiArmdiSjYGiQNkaBaW2dCnXMBxGWgbnyi0sUtx9E7AsRgs
OviAyLuiGb4/tNP69vdjbt1uteMNLhQ8i7/38jkpeHn+OSt2daLMyyDvYUYznSMK
Svzi+ZgkQ4duuK7P5rTdU/zzn47rwoaEvrcmzAzBekAtOqQobAXWA9d1sZzhLdaT
`protect END_PROTECTED
