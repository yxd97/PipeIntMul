`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yVB9hp/xbs7BtK0HOn0aAJbLo8a1g7M+r8C1FWygDbaF49x6I6JPNJQo+tmbB/5a
8PvfqsO6ZCt8GmIQYexUjdr8TXNzdV5e579lIG+KiwOrWWLImcKGx5h20XhZOiAA
wYr9imJGNrTXjuN0r5eMJh50PnRcikbgkY1LqmC1fHq20ayRboTozmR6FDIn5YbF
Ze0qjhijniG1bXfryUmeYQXc5Jo0Nx6JIAl9QRgi7yPiBRpuB9A/nk75wxfyPIDw
zRB7OZP7oHtU0qGw8LfNiG5vZTrWf1SLjUayZvlq1O3PfGr+Bo8k77NvwjFZ2rvG
YeOiGsw8NEIrlyrXi+Jc6+f32KuZKLl/vVeLsqwsLF0CoIuteH/Q2hMRvEZcCCyq
J1NPLfaW+dAd2UXb9wlCu86FR8P5jjz1YxoK+GkQn1hRGihO1/ZwiThHKTRUlNq7
+2ghgdSBvBOvej2paD0AYJ4Jm5uYdUaIrCooXcNv1NxSAlImxDDxIRpuUexdZpBh
pHEzQK6Bg/GbsD0KKBGwwNDC+pSO4dBaK6GpvpW/hTzlTSTp3y3ubxmFYdnvLg26
jCw3cDgi0QI6D1pi7U+vwgZ8BlKZMU+Iwz9Ovra6mt0mCWKKTuOmkTCxf94XTZcJ
ZCQ+KbZxKbbGKu56iGWno/u2TzJPDlqy9I+lDp/xSUBOW/JLk1JeBchP6INVG1sT
j08aSPtFIx0M/joEuIAeHIb4m4RuMYkniPZC8IUFOSju3ji7vuc2Z32jykFwqlLV
8U6jfH0rM4f/HC5b16+Iog==
`protect END_PROTECTED
