`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxWWHtMDyWCcbVChkiCW5abv3GmA9tezE86plPBXGgi6e6S9+Vn2ZIRA+ah3s1UN
9rWX9A2JfZMzYr1HIkBrrJSNKDQMokVmW1WLOEJKHNpFYsRZbbFVofwzFuvgILFf
yuieWFuGOfhQq2sGNQ2zMQUKQmsZVuA2FNkPfYSKtyDymi+ITzJKGwd2nTNRc2Cs
gJbmifRi3mTd01CCVDshMMKj/nynZKNyZgzT1asH3XpN9oz3kCxzFPgumIH5KViz
uGGrTjeoP/b2eU7tE2GUQUn4XscpGMOTiddT/AsRUGjoPIN2L+dQ3NAnBtrgfRTr
E4I0ffEXxbLwho1i+fwr+28RzOslZJktTtjmVBq8/DT/FoFiKPQyMfuFqjDpXUGu
P+lbcwwgP5NCq3JIXDNJU2UcA5XRd8iXBvnh+a43s2RdkfvxCEg/OmBnTqGFOzpE
UjlO5M1smzj9ccL39FLGY31ydtIAu9qxQTt9lQOGS7QGZVX3I4XVVcoGacXeXgXh
ZWt1327Yr1SDNxOFX/OHsPE7giEfRCPgeG/Sjt0PqHOQisstgAo59On3HO+1RTLP
LE9MXWRNrnhxlvsrnYBhZ2D8eKISVIhBt126/HHEvxTGk+2p1TzsjqXUY6H5+gmc
56Pt0slNS5tcexsTLGqMHRLx5kmBPe6Cu3O7vR3eGYLTz1NL1ObVtwNjglE301/X
71prmKg6cwWvhor/Jr3KUA/LddtsjD2vHjUIaHRUUaQNQM+42aX183nXfQ0sN+GZ
IPOgZ9XOEx4qBo68nQHnyFnPPyxIxbPlTn/zkF4TA1GIue6BM3cOu21ZtRYWGWRF
PZDsQO6tXLhcDCyGK3E6Hk2jAbbCqxk4/6QDYYg73Wo1UVWYhCdinOwN2LWrmr3E
THsrxz2ONcUfuiwpTE03KL76p9Kfm7isCg/V49y0myG2LyzlHDFRgBTHKVz5Adyj
Ozqz5nnrb9Y8EzVw2D2k7DLm7AhZWuEADJuLwu3nogUchhZtdyjKC/+jtjH8Dkoi
`protect END_PROTECTED
