`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpnORGal/2ZEwHfL32Ns1zH9xzwbj3gfjJBzDpisdP6aIodU6oBUGzmhPrzEr7K6
dWXO4SDuT551W0uUZ3zNNPt/1gw6wZqj8m7DgOi30tVli7p9DgS0xI3l6ITFYl27
BkuxSpX+Q2yrWekSlzEpt95Q9UyhkcqBltUFyJrC8RjZyI8J04TqHbruN44afPUl
ucBaax+rFQUTKKph88LJDnzRoM8DK9E1x/+Qy43zcRO3E835Lqg4VrOBmeFyodzB
LtUzF0M6Zob/BnOj4td5BodTUXyvKP3OFqt8WPFqYOylPVUtCyfq6gkUGmgFkwjy
m7OtJN77Its4J+GSy9vwYA3E378FcqyaYEZW5iGo246QlX4CTt5gaKOwf8K1No/7
T9y1MpTylEQnbmZQb633tK2dW0fn+FbibdYL7eLOcaPjF0K8aGaNniUvrRNuxBHn
LTOVbi/FmfzdsOQFQmNlBu9pK45q88iMFL3gpG75ackS6byM8Ig2OSVdE896Yjbr
jgQk6DLTb4rn4wvuK+lElKNtXokeHxV9qpluSidsl5TMgxSpqKGtS5JvFM51QUsG
`protect END_PROTECTED
