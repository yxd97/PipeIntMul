`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oF42HMEr98tckZE/fPC+k2W/iFdu7qpy8J/yGt41FgHnWOhIVD4cLOkTPNsi76E7
SbLvGGsU3gHFRjdGOSJN118py+ggOJJ9TXbaX9c/yh7fNTQ8suxuxwaiSZO/0RNZ
CR4m6bVfqgxDKLtbhbgTnxV+T6LTmrNmI9YKJZWZ3xrpJy0kJTZ8Dos6JpPQasUE
aIDM9egROVBnKt6weU5B8EuPyocOFDxO4jzBx4/mk+4DoVC3Vh7BgAHz6ivpr1vW
znFkF0FrTiUKyghuOCWCHnoKA7EU4T+uXrn/AR/jJaUQ+MHkmvmPAG5pimLcNeAB
rSnQOPpgP73wfiKUkMNDSA==
`protect END_PROTECTED
