`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WLdt0XhEsg4RCVY6R1W3elxNjnBousIy0HvQ60cnhTq+MEdl0G1XGWWR/2z764QX
35D7tAkvlQWlhmXhSbj61lepzjTUXxW6RlBKP4spBSqCaRCo8hPAW8TsHGicKS+4
WPkihw8Qpk9M2gpQ2p3ebvlDFIoEzQPGY6GwwkOlG2iilKh+xjsTeZtIY2T461Xm
nqLcfd6mIjq+YRkJRkwv4OOoKNfIcv+xVlTKb6aulyrhysAnGRQJIPQ0GTBW9bzU
W9tVBN+/Dzl9M8KX0fG5kPRvSAhVKvlBhaubQcbWdkGuPwbSSFgud3DxesJU5Nbu
dWcBXgLsCildDMLoJqTbtA==
`protect END_PROTECTED
