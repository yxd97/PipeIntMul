`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jKHU948P80orP2YIC1JhhQDZWkghR86iRHFhWOqKISpbU8kJr3YvbcA0opQvpu4
BWuZb+gGYaduYqnTsuSG0z8K+uPsxmJ4cMTsD9A9uls+P6oZTMdv9OGDUvVZDPq3
iwM+BQBHiEMcE2STSG1gjJK9wChNghCjMw1dYXZTFUF4qsr6RwP4dczC1joTzCkE
xZAHkGAooU7/yQFS9lc3HE4Q1k+r+92Qak5XUgqOkhiWh2AkhPdzj/vMH+vz3WFd
UkSzSGnTn1o7m0FzSMD2Sdw3UUbDXzkXfxRWcMaEdkeGemQZiJWFlKgCFGVfVmUX
+xv5izkYQyePz8VkeQflzA==
`protect END_PROTECTED
