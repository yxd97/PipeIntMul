`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PeAv1JbFnxv/9bzwCaop4L28YWOp3Lk1BsbjDJlR3YE8ahcORdNaawe3WvVT6Vqv
Fw6Kd7MtemjWYQcPMKd2gRfB1qj8DxXExI2SZF0SSDXIZvKj2HP227JutEqVcNLk
I27DcrAeT6Xs8NKKMf63+2dp7QyD7xjESR48T7I8xWh4MTwxQGH+ZwqH4/yKQ99R
8sGKJF+m/IkAaKU1z0XZLNkfNd/Sa6tOg6WhJ8sra3YGhhO7LLHypoRFRIE2wKBu
XUNirgkvZC6yUWlh8qE90Gw6N+3alTsUzOAq5keVN2aAo5iRL57dyhNPmiSc8Pyw
EkT+x+PMeFaujULzd0IlnZnVeohL9mNUb+K3QDy+VW+9uJCe02X47MSzWeeJVRNo
Vsh0Lkswc+nxO7kZUPFr40SEGpChggZl5CkvhU2GKZI1UQbK2a0MgPO/lloyahuN
AwrzmWAcDkm/LFlRUXiEE4feeg9NjWw+QB4THVA1xxmkLIkDqZfiugwiLIaszeaS
kbITw9lYh/JeXn4TiAjettwgtvTUbX2uc+GtwweZRqJVDNwykFtJroOyLfyj+yjL
DLh9mLpNTuVjtRRpc2Q7E0i5gQfdrwUlEWp8ZdpgnLPYfJ1SWJXlqLKbJGWv0uYv
J3B/QDYzasdzRjdrKSHS0Vj6QkU+hxG0hQE8EA9NTVsYM0DSaFNJ61DhM+Xu4NNZ
FToewa4H0/o929ttsInUq4Qi4YnataLb55q+tb7a7FfJaYPtk2Jws5KsUGDDcALf
NdvY5DgENtX1eMvlPF2XwvAA61EHnsPQrOPkXFbHFURKXvG8UNQ4mYEjGO645TF2
DzpUiAcONbdc3i0dXx/TM/XYwpFUtwGJsVD/EcTMDBxf0toIbqAsOdV1ZElLF2E2
zFn/u5h0+O5Wz1upzQaTaEfbDo/nqSpVGeZBWtZ+FYVNwbgMd6w+UvgcrsPHCxC0
1i3IA1rbUf+wKUOIj3E4/UA/d1mOUQUw2jtzFh8YJcg=
`protect END_PROTECTED
