`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0HivH4JjDmMqP5x4gqG/r7g9/WB6SGdqpBd1WYYtL0QCVnQEIsiEef1bzCQlHnjT
loMFyw8mJPy8WqEchojNLDhY5XarbooPgr51mtNRDfSdjhhi/8XfA7czrTp1noNN
qNqfRdkV5IREaWV+fU3KSL6ytOTSqDCsj4w7DVR73ZEvsn0Y7urJ8fU+HfXcvBvJ
47Do76vVL6I5FUB2V5DTZno3gLfFoBkwSMA8epdPI/ph/pw3NLsxXh9UvrVNPPN+
PlUyOYLQqB190mqn5/MWrPHWfbYsBXMOwIwKbJYUlgjFTAnocoEAFmumM7MMrdtK
pwmWrhfqNT6JKxfCsk6Oa61tRs4schPUWUYtspHyXgWwKpM4vFsJlDgsFUljZwkI
v6Pb/O1jkZdIO7Ed/l/ZcSRIvLgvDmrpCZgEErxitl875SXcM2LErpvuw01EfW/a
+ZDWqW6fn3QBeD+BNGLPspFb7t0GwLv5Qy55DvoNyX7BS+XN4SbEj3DPq8vw3zc4
QDcqJL1ME1sS/OQVGK0FizCNFLq5tlL4x7L+mVx7XO27rj6+O0LvXDoPcHA2cu5V
vzVPjegEK8o2oz1Sx+xjSV7RJmXOFdyKlok/nIlDiOZtu0IoIzaRQpjyUqPcuf2/
te1paqRxOfOmRAqcdmBhf4gnDmNqNj8fdMjikXyhvirAu4CjUzq8JNyeDrtQI+Re
H3Ozozsj/Di3TNPvlcVMJXLXFWgOPaE+UAoMYTsjQsSRZV+KLGDqTAdRnGqi/gC5
kUXc4wmGpajLAOaMbcGh/+xXEA8o2y7j+yeVD1vu1bO/l4SynwTf6rYZe16XWZxX
mDveyg9YbLgNku56l6v0TaCTbW6NkaT8Ruts2sv3rw185D44Ceu6Dm3GBkucrG64
9wv+h3erkpuqn3Nxg9/z1bS2DHhnGI2Fq/yiaxd1vGGI++JEnm4F8BiJQ7IO8Epw
`protect END_PROTECTED
