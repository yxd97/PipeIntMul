`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTo+U1ZTd61XDMNKq7eXAyXpIdwZgbtB9aAauJT3mchwLib/M14On84I8S+cdtQt
gWOUPgs2Bg+QzSM6jUIlNxp2lhByJDHwPzQQvW2+s7UHc7aV0O8G2KSbcJM+/UGe
lSF7JHNBA3LdGOuh3sDmd4a+Tuka6T6WNwBIl0nqXFOSoqlrzrNUaZf6nK9EPRUi
OZXPg30UZuhhbbVseL26vKQzn5vJAAnqIFlMLDLtJCc+3oFpG5JrtCff1ALUuqs1
aWlaHw1A36i25d1l1KmfRm2F0fV5tW+QFqGZu1lek+ZNfGZLF2M/qIFhhkwODxPT
GoX+j6WFURt1q9yu5gWSRYxI4uK8BCiM+UGRotIwrBDY2ga4gy/t4vqWg4UidYlj
o7EEx2TcOglhnckC+gVS61SradSGe67t1fGtPCw4IA1h1R3i3mxwnRHz6y7v7XZj
lVpPqcysVW/yrVOhiJIcJsUymeJGmta9ehAjNeCgQlQimgYPWGKSWMXwaTiNVpBQ
wquRdL+tp0LOHH/0RvdOLKZedynLAP/MdVdTJ7gq4ucgTTuuXzYYdpyuT6VC10bQ
fnphLXTMROmuRHV92mfh0aU7ZoHNNt57su8azSTDSEMJZ3mBM8zqxOUNgsz+l/gM
p0mRVr7kxzefXG0DxnbygkQsSGns9RnEDehG5hE7API6v8Z6HBggCltzKztHCpud
a+GHy8wGlKKnAiH3bgDKP0IySKhZs53PevQHdLvEoy1Pvq8t3wT2DTfcxVYxbbuz
QhRUmrHYMIspf93ObINF0Yp46b419QX0HOICGsR5ar2ljlZmp/AnmO/RKR0zDegr
bf25HLWPZjN9v3dsf+HHhd2L21cBZvDG31akVTecrt7p5ZPOWX8gFOUb+Y7vfxtO
bUhDd//PtAWBjKqrmoBS7Aw0WvO8Dx4x3DYWHub60FD3LgxmQvjm7O+ab7PMprmG
eMGv2pggnTRWr8EQMH5SKKc0sKViePH+aV1K0gAygsVBHhXoll7vPYKdi4pu5yR8
OuCH1GU8y7xbqXU1/5Idyp1/joVb0XBCim5a/a/qL6M=
`protect END_PROTECTED
