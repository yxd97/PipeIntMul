`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zvx4VeMVEaZTgLY8xCQaEjYDsWb/zejbUcWKBAnahtk4D5kIW3Oi7M6FSvZpuH5z
hvSrnkhubI0HwU0dtuzVP4YUOshpyLSA1VL+l0/HEiMf7pXWVGKfl7/gDl/Wthfr
LMO1q8SHzS7Zu7y8wSPvZ+QjbbyXhwzO9tX7rbqSx5T14pW8iTgcdDk+QgdUm62/
BXQdmRWG27rCeo8MEmE0SFigLW/+ucJze6Z8Ib649Ng2MpYzXDITGzn+3wdxWFZu
`protect END_PROTECTED
