`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s1jvA1fMzSLKQ9mQZEVoCMv0rvSxvuS/hDvHYXdKmm3GDJ/IBf1CJyZAP58Uvu9z
KG20L+q4uuuv9tCskccP9C6hSkauBi2eCzvH0kCfyyY/kYuM5wWcmXwcco6XZhcP
Byl8q6N/WtryeP/iHi+zrnXfYwNuQrRoy/w2YuBvo5Z2P+iH//Ii7l/kT4MoygGp
IYviShq9BCvtjXdQjPU7QFiNLsEJp4dNMyFGelX6QD7aKtKYOioxuX4xVcstuROv
O7v8idfLmolLFRwBSNMhg/sw1kIzx7rQQ7oOTgXuRrIVYNbusnT5YrpcyCYPb20L
fdW+lKOAmqB4YQKmTOs1KQJtIM87gh0YZuD4KBhcVXKJvudjEWwjN7sxDOwm+nt1
p55KJzSc3SqBNVyfjgXs3G8eiXQdDPjcO2VWyFdD4SvVyhOXK+y7UxmP6q9MoU1D
`protect END_PROTECTED
