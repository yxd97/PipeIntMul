`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2a0MZMjYEELrPBMn9hjUtOeXe/7WL6EYABSpN88cwjvcO3R/gKSk3vem5IIZOgQG
qp1rq14T3ndjqnJc9/iIEKQCtDCl4drAkcBnMU2YrTAgjOxsMzHlIQ78JfyNbPZ3
8cR0t5tX26KP9KDTk180VCgt26YyVjnjMA+ATA0eOlqoQIo1hDvc6XRB4z7E2lGh
yXmFos5VnhfqEJ6SfQ/s1Szi9fLlqPGWF5ahbMnOfaWz6sTp0fteWZU4uM4C1TO+
7TlmmJWIDLrOuky0E6X7KzisjQ5oHCVzT1pqaZ741r8=
`protect END_PROTECTED
