`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHjDhbGe6pTcMBVvkoNR36qg5vhL732i7XIw0EYtQB84S0dQycczIt/SoeBOWXia
NpVh7+/RNoyIBHdWkX/fE0gMC+8Z35CIDI4Ex0H4Vq+Gh+btO9pTPXqIMblkgNx1
JkDKLtJkX9y77tLFSQgb4Qw2S0rYtwVwVtbJ5h8cH6YizBfZTfDR5RRBwUyuPvwb
ORHW3G5ncAlSIed2wRjoRkzfN+3tLy9q+vuZyVnwI6tjlQVKzg76ihzfDW+vGY02
RNxyRfHvhQYgMfzm35JJYO5cQbSVeqDyZ11sJMMvMG2J3JsDyR8cwiVn3zZHyk5g
DfeEjS7t0IwS2PrtvMHGDrCAtSD7j6J1L9TB8YXZY498lRS1ltf72M4NgCHlpRG9
tExAXG3FLk45QgxBO23JO33r2VS9JSBybB10+xuSW5I8rue2XPQiGVSfqTELFzkE
KGtB+e5iPKgZsWYkQRsCSN32ifzJ+Yrzpk6D4noEFKpco5YEnEji6JptdeKKXtGz
uKUvqQz92GZFjoW9jJtNYi32DBrHbRLG9pKNXdDTJk6HanpRDSXwV4JCyXVrS3rj
5itIZA0r6zTgiHhjyslauaSf8kf9oJWAVKsaRdwIV+3hIg4ZBofK7g7I1tzs5xfg
+RFVhqu/CGb5JIgH9b7D/Ku8zxWucVnKTGD1XrSHn+JXV7HzgC55CWzTv0pzVBd4
ZVU4/hk0iiAVJxkkgvoyPsRwouRMgFYTfMaKmsHupr/K+BGv4gwLVObUazrl3+Kf
xatkMaowl/N6plxnqq1IzVvL+c6EhDmbUE5E02sajquVCwQOPALDApeX/k3LtpMr
sGHr0N8Tgid5Sim2nZnMlpzqm9bY+qCuilFAGwJA1pmTJzkt8Kr+xT7QwnekEdA9
lSBR+556v8+AEPHxKzjPgBeAdKMV2BQfoc34JRGQqmyJmJKI9uQs+0Fyr88LFS7K
6DukVMWQ6Y4JmZonIwCxaRU4iOevohSuxijR+lBOQaFxiLgLYpFi+fvqNbU2D681
idTDSaIbcN47KYPmVg7H4cSZ7GI2RQUuWXWEzdonrSI/aw2owodgTEV+FGtFCVV0
EylPe/RjXAKhLQEQKapn533mpJkpNuxGxAiEJ9vGyqJctwWN1VhNeFXb1Ggf1GNm
O5h7Q63VmgGLJyM8MJiQs/cSkv0HpemicptNQxWFa6VBJV660p3H5x7y2K/tvnLO
0NaKkTa/CVI2eUDnnNSdzncGKt3gIoLO4C64XKnF/z0ZXb4g+kpZVJblvfu9U4TE
715/h1sns7WaT9UTfe0EDSzLksIJe6msrc2cuzeAMwFB284ZrlTaEMyjnpOJrrtJ
oOccUItElZi1dwRwjxLmsJbaTRRdljPjpJ/6ousJ79kNPRhTTPJ1ghgXvO8Go2RO
DmDfh/gS/pxdjlh7B39gz4VAvF3sJPHBObMF2l4K+x9WfLZ7VkYtgffLPcwY43+Z
+GSmiolhrtpJ6KAWsx/aAavQ7eS9/a7W/5/XOW96uzKeaHUEjyaXE3ACAaJO8ExL
Fl+bWphYpMvitCBYA8WjGQ/k/Sj89UM3tvwYytEfnpYonlq4R4L48PAtQpbS4PNS
IEtB+lOYxfNTa+oPmSlK2Hwp1iErRl9UliPU2ecoPn8ufi5Wai9mktMdtwnx/+J0
RA6fhkpiZ/cIoE3Ye0HiKqwU9pa0nY5SC9tGAPLzY0cFGrxeqOQQNGrwuuccBcUT
U8wli8gOxY+pl2h6S/4ijhO2AMbfPKtGRZTX9hHkXY2BXjVmxPS4vqVY6MsACBBH
4i2W0uBtekthM5fO0o90uuvWRCP6IPcLxZDOLFwdchsui7L1B6uZOe0TosCpJ/u4
SqAuu+8sUG2StHARoArs0g==
`protect END_PROTECTED
