`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJy9cknAFNEikUxJZRlDiZVs3BMkiBVseDnc9ONb2JspzjTHCfL/TFwKxlUUtNk6
enRU8nrBhIdUVXbCgGIUZt0MyeFPuTuhK1VP1O+UrQE7VwU2qdk9siPZrVHdT5el
fXmeiHN8qZL569q2EUApTzgbA4sHPW3Kl0gL19SS3/tyl7WlQ+YCGDl04VvMzv98
swbsnLm+z7omAvnX+4KMW4X5EyX10MNSIgrub4BVlt5A5favek2T5KmY6vOHgxw+
MN0ZfgCm9Fuvzg5zUNJrXPRMK+cbxOSqJXV5io2UlmR7LCPgFfu78D4gBRPq0OPr
mAp6ssIBdzQ1Tt348zRpkm38RMwsS31dAWMaWkL2PcKshttLuJ8X4kBQAB9pkcms
yvd5ghw6jd0/Lo8QP/Zr3+hhL9f6pDRXUfTnreX4jodpKIkO/pi2DgCZefMgTQhD
vpCdc7AOffyxp5JUaBvtx135yrHKf9i7G629kmcDwwW7SdAYKLeSde9NOD9NqOSj
3T3nvkjvIYdKrp8kSa9SvOzw6Y7+UpPuKQlVIAYxWkS9X6f8xEIYzIw6NE+aHZLO
7FG9KDo9a0jxx6AtaJMyTyymCmIjWCAHBSfS16ijNa1Hfdf+4NhqhtEy9JKz5djq
LcDcLt/n05WIRGLvH2O7pEhRVNb1D4pInfWj+zscHyKw+xv5MRMnvQaEPVoZIrrJ
HZRKSkg9Zw9wOKRYhmC2lZXH9N+7rJTLtnLzeiksd+t6Ry6SSdE5QHDqmbOhwsay
vphvhtE0tDYroKdy/lBRaKonKznSKWVSGLCPa+t++FoaP8G0A8x0pm2FDtARh9Yu
3VQw3B8fBy0KzSJQre9pWrEy74+41fqLWgxhB2mgS0VXNNNbXLh37vovvOTsZb9w
ReQ4y30BFxKhXEGOoBdjaOuut/Qq3g8+eNRlEiHFWpPLCCYacW3WM31GGlFvwRk/
`protect END_PROTECTED
