`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1cIJvCPrWhyrM4VHJpluzKTn+cmbMdHsSvmZqlki2KFeZvp/2lg1D8cWmc3HZSK
DKL0abzzA0EPll1LpcQx8nAVBaBFn7MRWyNvoZH/Be3bwEJGch3u1yST0SW6hJuz
NN8WrckYNZV/CK6FA/UV0+RPpKWmCTA3783MFGBUEyZe0Enh3OPr95ycXZuoSxLC
DykkQrnhnYwWbfUCXqymuJqjKg1/yMS7NHRwPlNU+/9NhhBQg2kjP37uuJ4zuRRf
YiM1ENCN8fxNDVOtRgKjTH5yoTyTgKdCgIZN1KuPiTnC9DiOZdIZJEVs/O/wm8p/
wy3DXoww35KVn5NwZsO+ulTLVzNGFlFq3igJEWiSQqb9HaO24udeQ79Q8E+zIAB1
Gd0en0J2/28GOptDtM0Vf515ITLuFVLkcKzL7SMrFhVjVAULftqP4bSnZJo5pLYF
`protect END_PROTECTED
