`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHf3uHBHF2Z6CG//05+cULMqqbFVqUmSa5Gir+LpXdSGy6qp0C54vh2mtjTgnfoA
dybZxjVXdCKoRcYOKsl6/0bcqlrErcCC/lrJ6bsjVYKqPiCypOSzbhsYAD54FlVe
z2NaVJy44XDcwPYmmXzO3xR8eqBumP3Gb1gB94I8i02+wI9laGCBq9speXKn2TA5
YjUiveuvDqT0WsSz17b8wEMbQYstYSOKaSdIxycasPOdsvyG69jFbQrYFA39ib39
QsDOwFeP8z5jPLQ/P6SAUneIrdgu3a48qa+p84alUnKoEoT87IUW3OfrF+j4nCHP
qZD8Vlg08ZCTcSRCBRV8tlxCI6p6kU0Th3/kUZ6tKfcJsC5S0a/EYm+VL0j+hA5R
1TW1jwHiIzrhEMnYY2d7cUBa19n89f46KeBLkKdXM+E=
`protect END_PROTECTED
