`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQvH8uoxqzKKmfiUSRkXn1HBNkkwzd5AoXNmJRB6xz624ucDMsY3vrA/pfTJdR7I
yzJjufeYvLVgUDxYQ0MZitFY3TGHKWePhnVmeEuzUYx8BojXYFH95Ac5WcpKXSLq
8+HYA2yPsrNefgRMxUlI/hk/NqJkl8cA7lSLaTyxDQgpohwzA58o0Jdb9abQ+OWI
NcE7+CXy8IHNuHv/E9IYcjz7/JXpdCzPduCs/BSmehfpGmsT6bA9y2+9EOg+RkIy
PQx1ysrwsTdbmyT7/HG3SjScNzm2fl5983a482V0NzkHNic58k98oPw8Uwzq3koD
vQSjeGF4lESiXKqQTfTwDBwVU8CXZmXZAfDvxrQ20hYJi7Q87P4sZhhudjpaKEn6
2z0dzMSmPkF6hZ9nm0E9H7YYiH9DestdrKHWNX3rb1no5FoP8+00ETKOzqRNQsDE
`protect END_PROTECTED
