`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vfCv8WSpzQnqUK1VrX2qs8vBeUSXT7tAR+wRgkvUVKoawMaISejd3Uej+sIYDUzy
NbKdi7cUG6Cq5oeR8JG0LfWUfeiBa2mVkBNl/M437uPrxi9u9xD376rlPU6ck0wT
ysOk+TNMifX8QaCMHV8zYnuySH6K2F1JibKAi+ni2m/Kajvnm8hqdAdS+THfZ/QM
/jpJIJfSQ5CCxL0M59ytaK8YktqNNZp31SG0iZvH00I03YrA17lohbt7O7hokPIL
aDmkK/IDPrbmUKK5N/Mo+lsb8PUFFDsil3zUlmBn2YpxoZ1D/1jx55CXVR5rUAiX
mZ+2E5FbakPM63dNyEqFLfhX3i80eNKfpqPEtQhJLgjr+ZNhzJz+Q3tevklaJdU6
3fMr+kkUDUMcAfYA9wx9Xsww1BEFOtiI2p20Mo8Y4aU=
`protect END_PROTECTED
