`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9B/RDtt2UpjxlpBelDZPyHArXDXzy7NkeOg/jVupkO/F+L5VBqOoK6MVAWciRaNC
Ua3+YhA6Z4RPFZSbEEB2JS+XQjaK4Vu+uFfvUJ+8XkIBlr/ceU4bP4zobmZ7BlpK
eGfVM8GytmgK2fXlsUcC4dpKvfmKZW4YImi92N6h2XAuJhHLeDECkFsp4yBvzDUC
AvvIRPuoOdMlvLsuXPDm5mp69l4NtLULDJA6MZBNc80XVEbXqkjxg1+FeAzbWl9x
RWpzCvZPfPXcQyorY0AiCC+OkfokkAZlivN2Mu3D0YT1FRprzo6YuxRvP4+LRx/e
xypCSz5uJeVue2Dm0iM5vaLPhyjcUgYg/ektkPWEC5CSWUZYltMYcBnQrPFRMFQN
KHHCj7s29PO5StLjfVeWC6hGThFd6R6zbIVaWvqjY/JHzAcLxMkf+5ucbwXDdGDE
`protect END_PROTECTED
