`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IA/qjS8BkhTAG2UCUzseMQqY5ESI0c/OCugyKQBkE3Z+g6pEhfqGImadNJ8yeIHS
4x+XLSGQYCElRdLLeGlWxu4Edd/YZmyCnzlsdsaVKxAp9yLW36uC1RpUaz+mCODx
lWatCg/t140na21pYrtOTdjlmEa9oqUZT7frG9uiRM7kFzzzuEBVEiqMqljxsM43
xy3P/1gnoFRHmvk08QsMd0B6UYsp14xCpZ6DBJh6j2uIC1AMV2pt+sn7GWVEjWWe
4syGni25G7wOvSks+vfJTInMFXwNHmEaNDY+Fd6kWkpyaCSJzfi/lAPt0UXukPwl
n9eKzH3WeaJHDgfDyMb5g0hHpFIMJ8S/8uAqb7IkU0Dix/5aAeLvZfcEZNeXKJps
d8C7abX9a9dCx8BKhe3RJZbfu4IRvwIfl52pvNQ5Et06t+BNthwSyuAWRHGlwb6O
VyBXN2zq+dizgwsSbgQwBcjnU76GHHPuexmoW08mwZY4cqYYLMSCBYCGf6F7EXV8
9KLhodfN0mCEAe0U5ivZYkWhpb5LrzHvyCazWNM2IsJ0f5MTXM8y0ikQxuzAsfVa
glGBW/ACf8QGfcHJz1vVBjlliwdujN1UJCCxH0XoDgSCjbbsMtz+6NmZ4y4AzIdY
zTTAwpNt2bLlPbx5PDr8KJ2gN6Vz9J587C+JOwnsO9WYWOKRGCr0PE2gnyx3Zn1F
TnaDU2x3UdCoZz+smJAL7Ow2kilsZ+yUNGoI2VivYtuQh/Rr8PoLOXeu7mxpRXTd
O5ZFItLwJ5PCERDAH5+EWEpO7BkCul8GYqKjGZChFafGHLKdA9lxt4NW4o+Pwliy
dIGW+JxiZTULOV/LnNI3nPYBK4S9+kr5sTKPHXSz5gM5eoDEY5IfmT+iaOZeFqwW
2JHsMLGCu+38SCVnQDLqYmK2SPRY5flpUCBh7z0JWfvvBQdXiVy1+KfIkVrwhixi
2YpY9iw9jvIM2t/PnLPh0WA3kobSJqQ922q0FYPU925Sfdy/rRBRxOISFa8y7kOs
BlSUdo0Gnsqrb7LCP436Tqwc9TCJmqBwCPzkeA7wW87pdJK9ECTvxHQPduYWOI4s
v+8fqceJf4bxmH1I7pIrkeHhm8C3WRC5tmsS2DBIbiSClSjq1gVUl98ulXdhsz61
tn9bHquJB2USlwFr4DbIo1wZkdtRj6joYMfDyHji8WAWVpcjfsELcKUQh94UkPsN
Ct6aibD+BvzeJbGkPKGcuyxWwcleo+MuhUUW8bw7VQeOmIvWamSXEo1xHB4LELQ4
iN21/T1PdNNnXAy8NJeAejHzeTRv+pEBxUD1rYDY+9yqLymwFc4ztYhRWws/6K3Y
qEEj/fZnNJym3XEIihS/odctWWnPTP4LxlMSDyxFBDiScAyb0CCxM1M7Mf/nrnYX
cYo6T3Rp2gHfWoxHJPCJFpMCFzb6/kj9CB4ZpLl3ekz5/tmSOyZn9ZXYIJGqyY7W
hvI6Tbtl4dFzd8jG6M9/Ya6WvQdbfS2zosJLpppakIPDc4t8KCRFi1yNBTdGbXC+
G4bovWiafM6dLA39sODDznEWwJ/LqAziGBGzwBqN7Qsbrd2o7OP/OuzUV2mRrxVn
3gb4jC+UMS9FyRj9pXmdBUya3DioNqHLhE/CiVXq6wOIsgt9dGhqO8YhlC8gbbDd
Lcd/TMllpqdVOot6dAsDOfm+a7mk6X5OIALoNj0eo/IsHTUZkqdOR/N58r7Moume
+X+dLfS5A1KyJ9Y5lfAJ0hsWg/EBcwC2Z/YdsPtVb9HIK1CaUbFPMlQ66T++gSGQ
imE8DpmaCeCRL4m4IXj0LzU43fn2egtFEk40AWH/9x3NKp7ya39C5smxCyKStIBS
aQORvbryI1IrpLpxliAsmayV5sy1Tk0xrtxMgV+hXnfk7F4eYf/XvL032+7tHbFk
XusRvRt2rmvdRClwHtfvRRRwN7XCrv6ClRjDoYUhUZUSdEpok3vxvUo3t50wWEJh
qQA4U4VpHcRIq2e7O3Nck/1GQJpOjt39d1sOUTDDz/dM0H63g6FBQI2+cdJH8Js7
GZKbh2Kr5zLSqz7L4BKJhQ==
`protect END_PROTECTED
