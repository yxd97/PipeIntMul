`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTzLlhNW50vp4RFgZiNz91ss2i4XlgBaXrBuMvbq3eQjaisjAqln9QerviPD05qe
gppBPim3lkH39o6qX1yK+RORvfUMZwMjJolHOBIBll7Ask0OT5Jt7zIGSYj7VhYm
dQ6Zc9kvBBHpOHxCSUQL67q66Wne5wt58LCCfEdZCvnU3ERi2QuieXW8k6016WZa
z32Md/AalYRQGNuf06iXL1vppO7H7qq+K0kdYefulx5r20VYmFnWlcfCnLEoEuFD
UGLXoBB29dGUdGRaoDMR0dDlF6LxDYi31+0JtvuZqxgjseJ8TH8SMGukfw1erLkn
UcIt6C69yXMphq5S1s6IbO/+N0LTFrDxMtrZm8Qy3ojjvy4qmb49zZwHs+4pU0sK
5UoHrY7WsdcAF0nnIeWf+JDWGwnF5fRSSMc3rOKSDT9HtKPYUaJB5GnVVuXg5OPA
0YLkl/c4t83fak+KyVuZELXODimCV7jxbdWYrYt02pPN2lYm7On1DEKKIeWDyRUO
N9212FGuOasgNoSwLhtCr4xpjJhm85xtb2vtSZO5V6IwQKfTNNDrdpToXOUnnvvA
ZUE0Ap+JHmBukiZR4uPPyQ==
`protect END_PROTECTED
