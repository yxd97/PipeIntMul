`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g1ZhB+laP/p0WiH7+HsVWdmx+p0SQ4o1A20ibGREwOw4Mvb9xG7IF/9uR3aTBpX7
NdhuRm6e17lmQNzcQ4qNsdIo1UWeUaFV+UBDoE0AXVHVoKRpP1Lww0qNnw2+7A1S
rjajBlxTLUFGliMdX0VC8CGThM8NfxFWtknJ5HLLbytU0QP+7FmVIxLMTij3HA/4
g9ynFxmtIVgM+P1zMNRdeOl2LhbCpDj2iSSyb09Wz2k/wZtzDSoqo0yoEROctWvn
aVaDLEKx6+EjB3W+R0UXqseoIDNjjGWUz9mJbBVd78Z4nP79FzE0XhPGFbDWUTfz
DYJC03rbsiDJKnCjGANXoY7FEPV36Q+7fGrSnJjmqih3sHW+kw0sfxf8zgHfwzBk
2IpKb5Fk5pEhbM2FJNUNTm55wNAyh7l9Ur6aTLhamJiE6PdCHTEnTEiZ1XOcnuZu
qCFfmpIc8fzICq/DLXykjXNF1/8GtRPcnStfGodJoTicLgVMkpurTs4qa6+j7cu6
`protect END_PROTECTED
