`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bv6bV9z9kny2xv7F2HDb+aW7yl6ikjasM+BF3KhAYDvEHm6Y+bSJ4oLiE43sL10c
4NeilerQCzr4qfU/JerK/w1y9k8iBe+j94CAYbd7iAwcfw4lVv1Eh97jaNvsHeas
taGiGoODeSwM+kXWxJaBTYU85HtOr2QjcbFKQjXKDdnNO+OvwwpzwA/CwgvS0U+K
Yu8WE82xKq+Dx76H/zHidxZI+z7qDwQGk7hQlezHJEZUKsBR5N5IEkT7njL1qy9d
S21t2YgEePo9tNQLMesa29546srk6s01/5mGjrpPWOsbKKhrArXqqstGYAqrRiIy
ZRoKv4cdBpRLoLTjXtQFRfRWq0IkV+HNvUh24Kpxu+PuVgmwlv07/zjQ2I7zUyI0
M3dHvgbypHtyACDOEh4MGEotkrsKUtHdfX2vEozJSgjGlBueEjrz0YUW3xAiWepb
AXG7PaabZVoIkrk1PgraCjQ8k9mDFpOo8deAdizGiqVoubpnt/eBDMWE8GXxOW39
wmY6LzqizRMU4EulJD6htQ==
`protect END_PROTECTED
