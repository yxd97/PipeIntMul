`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65pcQJ0I9nhqm3rRsz8YwZRiQH/MiaD+8O+89xs1Y+m5K2REpmLS7Z/REwMwYGE6
w2se3EIyiRZWwO1av74oSbgQKL9m3kwEz17GtFZw1UJVbTdXlosrEB4EpAXA9DJD
r0MGKvCSazJvBnEnNYXzy1lmufw6JfkxWVS9Uc0Tdxj22yyPiJ1CRBBLPKifat6Q
9oS1FDPtA2hJ9sPOpWMDMq4iPmwY70x61Xqd6FVH8yszzsGCNhU+Qb/Dt93CfxlK
5ibqRa0yieC8WKZ94bYZ64uFr0JAK9nOmdAG1xTH75kenh5Ra6rSbeCgSOYNSckg
sFSc3eT63QqObsc0Cu2KQs2XsiDujZGAEfqeYEYdKcJb1AtPGG0YWR5JFdS2PA0U
EAZQ1yic27yK9CsFdO7p0x7EU2moQkSV54k3Qpzh6odE9KJ0j5ZSPI3XuSOfkGYg
Ufs1X8GckXH42ZQ7ZRNAhQULub8/uBsjDllEIc5BF1mr50dDi/ThWcvlJSsoQ3Dx
cItrNtIf4SJrATuDUsYwSMKC7nVCR/iIs0HW++NmJC9RkgQul7BjI5HyvR/BjvVD
zunH2gQknCvLAJLaEy16IqTWm+x4Tzd6TJTfYn9MdS1x9DT/3rVKr4iqs5QCQRH8
l7n55QmP4Y01DxEhCxSQkIxLhxj7bd+IOen/xJXh2wnYNaeN9iiSG5kowrDFyNeU
+88QgLTndL696w2XzKZbp560NmcIydx0MYZV6Tx5/LItQFOfxxdDa+/v/okPTJbM
srWPJJmFNt52OL6qjgUL2uKY8TSP1/oDS5vbMe4kjmTg8CxjUOOXglwYqM2n6RAM
kdaw34QnqxN0jT/Cp30FYQ==
`protect END_PROTECTED
