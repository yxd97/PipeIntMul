`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eYFcSSbIG/DqyjwdTpMNDSoCzGLVIebuScXKftvDROPXKPTDpUcw/LkP2Yamipv5
QF4Gwbr2KhLXxuP+3/lDd7GPLPwKOhBv4zpkwuekxJseyWLCyXsBIIRN26feLieD
c4kekrQq3d9BIbe9h+p6yYg8ATCABuySh5PMFP4oSq/WzXqiLCjVCXiWxACcsRie
Y+QBQXw00VlAfVNBpccF3Rb9qEGjb1XOZxXCsNwcF4/MPdyr+XXfVTK/DGuvdQbA
ljk6vY07LPC92RRdVGx4Jw==
`protect END_PROTECTED
