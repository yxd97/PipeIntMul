`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9e3XxEMJ4s1dnAwVMkJRu5rYU/d4nICvc7PiHmqs51h50IcLeTkwEFQfE8NCCwK+
JXSJQbc8aG52esHMKyVvhNZkT7lP9lcLaIIagwnznZIu2Ydrs9oYCMtv3SJYjkDj
B4sxJ0kbuABin9W8PdvkcTXHSgYMsDCyo03bAp3jED+Qv39J3rrXnNZXJra1qqpL
jCXvfhmS4zHsLQEu4Dqeci1yTIXZuavB+w0Cjy3wizkbV/jKLQyFsCwF6biPwk1r
SWXlWiKu0TQTEYRfOF31opKPgoWUBZu6C0FtjRgMSlE=
`protect END_PROTECTED
