`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KbVf3yezl/oO3wGzv6DfSIHN7nJkRQ7hexT077aiwtVA4zf888XwdLngIBbPtkG7
m+Vj9M11pQaaKroZwXQSZlnexVcedNvSwilI2T/ewZ9OkSS6Zv2ov2eWmyiYsArm
NW1oHi/OUrsRpGmvX1Xg4NhKCMCD+DFmCBZ05oBRSqKnFFXUamWIJW/2wFC2Fxpc
14S4oHaYM82pHhkLhU49N5GRotfnYit1Q63urmkxXqZizlti+3aqZJ+ZnWyYo4jH
KrI6Aj36IIE7IvvBlnYJ4z3tLdSj6nwjhR0J1UVqKUYlR4IdMn3hGne/QSyQtHrl
L9pzMAhl3LvffFwb3oiEFVlO/xUi+zNHzPIyFZWrhWFmxlMv4Dmj6NHzYLnWRpaZ
ppu0h3YZm7SU2jtnKsXMkp09WV+SYR7PA8f8YVZkNUptzC/l+x90sCQsqehJLvql
xNcGJl7dU+85qGEljvcNSQeNgkYCsBS0J2py+BFyf8s=
`protect END_PROTECTED
