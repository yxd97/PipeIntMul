`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X74RHmBl920v4dIGM4dixanod8FFOSRlthxAk5T4zZKesVq7CYNGu6oRa8gm0p9o
LYVVhogvaMzW+Xr4wT4A3LhfywVzU0WkxunIwfAqxjCnov9LK0JOeb4/NdLaA/UC
K/66AStQXpsocNJqdeXyv1Zx+m5fdhbB6MgQPMmP0wmjAfS5ZN9QkLN8jdEU0ykg
cNuhrXq9DmShouEn9ks5gRLfmwL+PS4C9r1tyPPQEGsA8MGQH2WbxHaWxgmQwBcv
qIVKoGS1Yykdfc9Os2D3FIdko6B6SLgMxst7bkQa1dAYUQx+JK+PoK0a/l+qH/TE
kSMTPOxFqhiuew8xofpbX9/ukNLyEYsZa+qs89s7ev+bbyyWSuiIQpnZireNFdn/
6tWPKkUUChIQ4651nFelFPfxcIlMIuZRRGlLmHlE5p7LEk0pi62XDOovxOFKPhDh
p4qxpW4I9k3dHBez4Rqteg==
`protect END_PROTECTED
