`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fKCPCch7mUFyFTbhoI/Ah2T0oNOIIdvlJC1K2rpEjlGoAzOHGs8omc3sPXvtj1D
2PyQYsP5e8aSdk+ZkKo8D7lW52DUqP/dEWzcWJ52ER1GDJ0XIz1AzmCcX613yzec
pWlSZG1B7m2DT+6j7+xiyCRq7pZqbnbq/EmzcbMm2FvV0Rp74a5KK4EyfGZkiKmT
2WBE++FNHvYbdRIXAXIcWbQ4QzSC1+c8NLKZkzTY8vOFDzLum51TQgYJp9tzXOJ/
ihaiiN93IHLrdeGeCfYP3xsn0Z+mDSUcAufh936wrIw4jpFGyJa3ynTdWFHT1UXm
/OaONTbUOkYtHpshYYANaABw0VODPEE3fQ1WIinocKaUMcg5djcIenBvWhGZVdEV
d8cG5jrhWg22dOeitGFu+WDxVN2LDvQRG1bS9QpKyQLP9dXvn1mR4yxxZFqE4HR4
gfrALuCLVGkV6LWLi+Geb5EAvjVTXtOKqbaqJdkGix/2MwN0oX0pb9KIfA1qTNpk
fsRFTYxaVuAWX1qtlI/irIecxOiexaT/dVmZbXKe9G4A3BzHJ6uvMK2pwmjwxVUq
4ZvHVKQtLt6IpiNmX+03qSkZjkCYhGxfXomqA64ELQqtQwMJjgAZUXJCR0P69Jvx
x8u3oFOG847I6tfzWRY4oSB1TUIjTTsThjpsU1Q13socZPHka+f946kXHhCcObl/
LMbK0diJyZ0dl/qxE0owiMoNlJZjDaBlBViOd7YvU9REUOV8QYJ2w/aJQrkob1o0
IRYOpMnHVWKbuJ/bJvvsuQNwZ943VJDTgmj8xo/78RnHXJ2Sqea5JJaZhPPez6qJ
2A8fzhpChTJnuuhqAV3Y9ZbI8WU9h1lIU7LK/QXX9dil8WkuWE34Hdpxt8K8QFKi
1ZmQp6j7gDsUX3qeY4JbZtlKRPmOQv8Rwu1NgfBUSLQCTJs/rBhs4Pe4IQnvsQRh
pHao9VWeh23M0SDa5pZvu19jxRE7sUcojjBZxWs7lbSXg7ip4BspgzLEYdbvjeLr
PQxCWNFwqorIJ27C3eg1d+riV2FzisU1uYi2BsrGMTEp3lDr33tS03+oAP4lYJdZ
JqQFRaDiRCZAPv0YkrBWncq+IRGT4gh+qm+WgT2RUmryJyzc/3hN1/ApUMMIQDmP
1e8pN2Gzk/x7w//EKyDJmgI0Cc52CrToPeJvWz6/0RtANBMS8qxFMBaTKOJKHt5R
ThvUkzOOqesh0itYvr9niLaN3/pvq91UwtP7z6ZYXP0FN0fCQLKHmgqWKIr3d4JC
jqKjDtgbMLbxDalTNGwwFT09VBimvxNkrCWhCANmYVSncjGbszHluS5R/+/qE/h4
DCN34NvqY534bqphMl1VitA2ld8X0zWkSTHD+zN/HMgLcOrfyLOkrjhsuskWCj2n
D5CiiDkg9nJCk2l3iGORQeiGW2ilq5/Ew4YeRpVu5LDfAfZI8gERLm6grb/zSZS5
OjLSzankKWFN6npyBQtvO9Z/D+ujB10OCKAlxn8omQEYMnv1mgJA5i78J3oPd6mq
DWspfVbVrDcj1lN8Qdu31bYEZuKNhdHrL25oYfIE6ylxEnZ+e+8ApCqjsR4OEpRJ
9mQ3wwKFBAL1Z3Zb9It1l0sTIS9dYOL65SaT7aheun8/mtowrY9xcWXNJDXdk5Nx
77dBbvGPLQ7x/A2dXJQXGMNUt+KZWSIRQ74O5hRPtflUbYQ0WIilV4sw2ir4VIvA
vGDIJOt1zpzUTHdxa9SfPbAkzs6DRw5KWRPVbdCYEf99v72R/OE7276w3v9slqa9
sOmyc0QiyELUJfPkbwqvRAQX8x9d95OA+5JzEdxuHbQ=
`protect END_PROTECTED
