`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6ohyr+WIsAMP6R87nEoGu6/RWzN7iA8ODeqHWJWA4jX1mBdrh3YE72WswCh+t2E
O4kFybSTUP7/ztnB8FJT7BoERog3A6dM+d1/03UgaVDNnZhT1bjodrBT4HDENvX+
R/T10I4g74AKZWh0wrjJP0/xcnTAlzNBLupKFbzAszPBOZMcI+X1nrJD0u9gjmZW
v88wDaZi6JfoNQtAjwOzoO/nCKXaqDrGJWdq3gV0XLlg0agvTzjjFa33iNXzFpY2
qediybSImpPX+lqhctEMVem1DgKJ4rPddBUbkferA9gNQ9VNultHD7W2Wt4AzDs8
cGXZkKPmMc8hrPNmMcMDCo1MduvezeAkxAVi2Tocilx0QlBVMS/HHSg3ALjCCqH6
VUzIiPhFx4m649rFS41ZGaJmPJK96PvB9bZV+HMFMRfV00HKzvkWnWXV9+kVnU5p
58UIMOVcjMeifu1Pbqjp5IyjuKSp1veGgOP3uWijmLdLlGKsuEqg0oAffxtM/SHm
Q8oILeoVCH8heppRbQ/pFUag+8OzEPjaXjTLzgHf8U6TWorQJ+FrmGJzNGnGRS1I
od0IKfwJmX3LeMHUR+OuBQVluw9lYjKzLF6f0I0iewaCW2fX5tqGnnaXKTE5VQqu
hJWUkgKfyXGUisKsKSlWNk3Gnbj2Kqlb/R6h/RjF3wB/QAdOw7PLMflm12FXKJzs
mONDVVKqCgj1h8mlrCTbsmkGyGzKjhW8e2tmBLKej7oNBtVb1DtQHhPh2l5TQZKD
Vt5H32yXgSmPxtmHeEqU5icUBVsFh7VuHJHvUgYLM4IDEVg1qiBa0UQwC+YgGCwY
jJER10Hy1xDTNZBqHnJrXSVnpuarChQCLMbK03KE0EH3ODww9xtKeprBby26xkT8
eJ/jr3lTk1KUYRpcit5hQKTdGGPn9tyv1kwdq4B9qkBGQSuwjy2VuPGYcp8E0LUX
`protect END_PROTECTED
