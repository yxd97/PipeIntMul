`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gjkPpeIirI98kbTQqXkDRP1OI5kETMKCDzA6/wJmp/2XK40xbPGjNzZ6wDsTP4E
nrdi0ywm1nNEcxRR/Gka526xNvys5p+DKXnzB/4iZH7eHaYgp5gl8kyKH6K3TDrz
lOZrrDOkH3dhB/65NI5pCADq+LBz6X1HHzb2V4td+l7wi+LAxryi+TgGLqV455m2
gwjEuTAM9B4eg1AzFDsAhM+ugqatyrvrvaKyZA3B9aac6CfBd7atv4FhsUgQCtPu
Lu/DXyy6EyTyxKyNlqbZZ/1biYHUT8OHuvUHcgCbjORedKd38vE7PUEAr1hHqLRU
hwe6H8H0xmJeAw9BI3Mx0yzpn7XokaaUtY0WJN0F5zIkIo567vyvq2mbeRCWhLIe
mzFV0D+aHegaY6nNiWG4i7PgCq6aG1NqQokmhxviBbw8MFytFHdehb7Y91YpOYkb
98txBNrsMqMp2GE0NN8yJPiRtXMlEmZ5Rv9ohJRgdKFbiMWMb4UIumLKTiwbtXMe
TX6YvO9g2WVsgRxOCZoew1i6m/oDLqrVLfQS4RZLUWehV5W4o9fXXVdXuXU9X878
fa3wLqfLKxs0/i2atS6uNBYZATnKKImH3CtYbl4urGQ+E1yHqXZ0jKKPijW9Aof3
K2oonNgRlmExgNuWI7t+vw==
`protect END_PROTECTED
