`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZspmOii5bu4zTAK+FGUgpyHkZfck9m2RVpu1egekIMKmshKzDTM0A/mkSM4Gef9S
ywRC2vQaQzaaAXQ1+OXpbtf4NZuB5aOMnP3cHRb6uR8wBoZXf2H3FZxuoVtabN40
hrFBnOCoTNGg5Ql+7KeShAy68kE6ry+JF3XDD08QiV55b+BTj/QuP2fy46cqtGIj
wvrDWpIR1VP9VSRZyTn8t9yLBXd0ROFfxyPZqDUNuBAfT8yhT51MZyRvQyyB0/kn
tfCF5qO/RkwqG5fte4nRGafpbzIRtxYgMgVXBeweyxnBqlvDnBRJrtIIormOk0jr
Jb3Uo2bExAN31vagUbHrVQ==
`protect END_PROTECTED
