`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9+zjzx/bsKTxaEpdH4iMwllHWQ9sYJHrDckDjdq39qgwLJddvK05pN0b68xNf0z
Y/eoevw8eenaX3Rb/eKXIaaE8RGHp35Zm5cRi+lUq9c6acFqcfP43e9gUZRoQEez
8OK+dDhuUp6BW6tZX2M/I5z1IXGjQC+j5maih1LCd6Wj0Gl3zVuScSUJutQ7CDhK
zDkMakPxQVhenEb9ILpd/62bREFmms80+t+P2s551AIyNoLIxtuTAoquvSTGY4fs
37Y/JWVBTs9mXNOKno9d2bINRt+rU+awHfQ3b/qxeE57aXVTrkhlEdjMOXSpYvLQ
ISUZO1kxievnwTIDSje8rcsTYE4C8ruDPoZ1lS0JeZWVMIjHFIbJiyTxQLKiJ8MP
u3L4Ek1ZKGeOWZwvdrns3OY81Ozekh8ffVvadmAXxRGcQyRc7bfvMeEkxCICivrK
kUIW9TGvtNkYYBzxF63vDkPN/dWFJcWDo/iYvyNzSEAXAtACjhVJ7aElKjGhOLkH
hC2uu/VkeuIyCtgrRUSDWNVG0UieQIdN+R//0INfCyMlU1JmKP5uXFOPK9WGVblD
20ilGhxrCdLHO9aC4ehdCt0fdsDp8nKHP1bbtb4zjTHJt/bpwRQQJGYNmbIPEz7y
vRN8MmlwvlrFlvXlT71adVMf9oMi/isxY6e1xDi/V1zN36IsJfD2x8AhpMjUHcDJ
yzT5QG4mCmbQza+BTKpQ2hk58+w/W1ceKJkII2URANuQIvIqCEfAKZhi1XzVycC6
C0GhGgHeNRYchwO9vGqFL6uHrpkZYB73ZhRirE/bmIx16O9/nXHExycWAsPoQcfg
ceNssnPTzhdy0eQV0JJMcOs6MFCE0BQ7G45dMoy5VLg27OuEP2OqIzCIiItnND3/
P3Fhlc1Pxy0RF5MvygcHByTRJVHSsIRn1p2YkqnrtqX+6j4kkrwKIsvzjPh++aIw
ieaY53uxHao9dkRodw+7Dij61mM/VwEI4sPRyeXB5HO1gkwwoYXYwB2Qh+FzGPwg
RK4Ldj18Jl5gXilQ9yPKna8kNLS60dU2pR8jbw/sxDk0HxXLgPKOE7sttcpyL25I
+hW958R35HC5d3pLhCpseCDKgiya5wFz0NEuGNuVZWmI9kYB578uZVC0xqndGN0L
`protect END_PROTECTED
