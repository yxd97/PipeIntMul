`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0DZSWySZ/I2ulQb/gB+qeYgE4WvmCLQgAVbZIaueAdVk4MiCBWzdDNHGuPQmEZw
Jy/Qgo2+6cjCYNmhHqVPKCyWQ5nptTOc31C+YZFjbmGFuq93vRNhTwOSQ7B4TFp2
Yk1GFWQHmRuSMfgJToRFNRPQTkjOhzIh8HvTcobzX7Ul2k2xAh/WNsT6+Yc/IkLX
Zz1VRRTYDYUI0NqlvKeg7WkSdwK85hMwyDcjXhWtaQYXVjgeGbrQ4yI5w2/X6sC1
dqDvqNe11osZbT21nrs3yfs0sZcxppPD4P1BcR2IiBlcBbU1IOnB12RpJTCr41Mc
Q4PrQHNRwEdH2RNkBYAfZg==
`protect END_PROTECTED
