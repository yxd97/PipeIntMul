`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76cHi3+TWb0h7dzOwxIsc4+5Ylgbowp2CG9wqUnpgxpHEFpB/OvcSwDyTyWRc2nm
Ia9JRUKIggvwxP6u0mcofRmNdV0OuvJKJaiROlsRruZWxcRPoX/pIGYFgZAlWw9z
jsOsGbIY15d4qb1foXSqckUCWjFxCaZfILClaG30KnM9vhds6Dyyvxw6lEsEqW9v
K1T+WcLpEBjQiUgPJiPeRL2cdn68UcY2CW8Mel2k0VOmVhNnzdUayDwFQxDef4x9
FjmMsAPGeIz7CmL+NCPIoXF65Y/3BOwEfPu6LQE6Vl55FTyxQWE/N7I4xcpN7u1H
oedpb/47TSEDrYGgY0UirszTFH3cajA2MxQv9BFqxXh2ypS4aoS2xfYOminLxVXp
NQL82l8E6sMipOAFjRw0pnBHFgP1d97RG+NIwIyR1m6IntioJGXYIdzuS/9Hoq+k
/CF5/9ULgbldOSiQBk8n4R9PhGg0RdOp7YessuFMLpBMfWpiFI+7QejHR7Za95eP
BFczS8KiQltWDYQ9dGNwKPrIptDSjTmrrzsmuFU7mGPLzOMbpSHerZkbuk7IV5nn
0+vDUWW1g00EtK1Q1gocLBho6VgI0p8N1JSRPH3/XBzSi2UH6Au7IzZSezrxtyYI
tv+EXb7IAJ/UEDPYwJWz6+lw2ceJXxr3/erVMVb3j7lEgLCi2Fju26J574rPhyMd
EQ1qQtnZJQZapHunA+NXftN3Jntx83aCvDIhbEI/W9zxq4K839DN0pAfFvilcyjo
Zd0AJdmmBZJSv113IOyjNqiMumalXEUh+1gKIowv8DRK63JKvN5c+nAns+aeqWOk
bXBjO2Xg+ChfrAujmT8gSpCwf1gop05FsBdxDqWhtG/286kGSBJBXBCOuNa4zV26
zQZv1FRC5xYWDKifUdNkan3d/8sdHEyEeCflSrHZ51v+ifffAClDG7jXVWZmIE+r
5/8MVduo1vxyXUeXXVGfAjg0tuHylrhrGs+5vnoxYZ2wuLSGRuoc3kr8XzCBNRcO
i4kzefNC2uZu6hLUGLsonwHM/7Xznd1w3KSx3tyv9Sg=
`protect END_PROTECTED
