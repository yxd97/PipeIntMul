`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8HdtSPZTIxX3Mxhb6g14lKPUXwa3WhR/sytbh2eF1HVPXzzUCz4rHOVjam2DDWr
DHyz/xXd0FG5LiX0pV18utQKUlW4b1SRljO29TKIRtBof4F85fFigJXMUzSXdmC4
Y2VJ2VjNhEG0pzk1J0ByZQxWsrqZvJi19TGYgwguRyuFqB31dzs15LxIti/LO3HI
htl+0M/BynGsFLZgqrdLuzFROhNp5TOonZxYpIqag+xuPVsXGCCEQVhWv4kk6Anf
IdvNJO0DDZ9kU9/oN+/VLol6QI2Hb7Th9Zd9IEefSrJpuQnHJzSgpkzKn9Tq7aZN
YCsDYD5rHwMM+dNZdGA0M+acmIlrMRM0CCUHQexXwM1Ry1FIiXrhBnzvNVcURk6v
7GT2ts8oqoweaG+S8Zv5Ga5hCrDsic2aA7NXV1wRDvfuHlbyrtkzQANwCucYNYxv
ecOUlEX7GdZWvi9XIGb3S63RSqN5VLBFw0yGsC3JaAltCD1mGXQKrlJR811nYZAv
HkUpKdQ0lqUdbMbRLmnriG/i5S11VKtjJIr2FzSiHvGAZbvi01ELoQr4nYoYPcgT
QByUlG6Z8/S91j1OjjgSfw==
`protect END_PROTECTED
