`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Ct4VxQjEgcwTFbxF2I7jNkGmfNusGzwr1Dj5aX7d2vrLltTbVSueEfIUJ34XAbm
vyWjzTOuK+QM2MYui5Q4dI3/WNe/pi8fKVXxWE2mfUYQi8jl8ojL1Jc4lkXChAJE
sFJI3IcRu84RCH1g7D6lDHSiF0ZqBEWGNfLjXA/HQjKSIoMiCQNNiAhTHfVDr+K6
puG8S207VHNPhja7O5qGNzjftsWlT3oUn/lHly9bg/K8y4Dn6o+V8m3Nhv240yG1
kLGSfPHEZ2YmSAHjzWgQkc9hDSTpLSEF4YcrdGyFIAePRZcxIWpR6VotAQCb3+tZ
SnD8FgcR+A8CaLaJyRBuVAJcv+nW5Bt66ttZbhfYZIT0eMcZr+R0f5gI8jE/HHxT
YUSCQaa+6lQujXhnk46gGg==
`protect END_PROTECTED
