`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70D/zKbgYH1lPrn2UfVf/xUI3kxPDSUhzO8GR6/PuO+le2XsVGMSrqENb7hL6jKB
Aw0IRxGh65ft440cPNYvcbIRDzglKLqzfxTAMGthoFCE1ND7NrhLOoZacSMMpKsq
N2pWXF8KdZ/zxb2LjUgQPIm4Cq0hichP5p+Md58QHadWCFBBcdKcPfH5iu2z11pr
3hNOzK4xCza5ARGGKxBTQQRdHocJ2i2HLMRY5u6Porf2Q9zN+opEOzTxxxxXxwkI
UygGeIVLHwTZBX8Ysmz0Zek1g9BnFHokT62RSStu4IaXoY9yvgamYWWw7Z7Bv2eh
QI5CnQcnZXpBh0Gn+FlqXLFbcB0mMVZM4Cg9toZ4LIVL5Ubp1davyeLMX17ruwPX
wbh5BQ+J5QVqmyAdwyCeNqK247KspHt6aUg2qFER9EtBVl0waoRIGLdmF0Ky2mwX
EbLyGOk4eS7HYbLHuplErfJIsbEiR6rfBOWscuOqSl3PoeNViptokv+NmImYF94Z
Va75rgQ9UAaAnP95MI6604D4E2hQYYgK0ogVan3ht6BrounvRwJ8GY/JE/KIt8vA
zt+lVF/ZDfGm88ZFpPTIfCTmwkoKqtadks3KrwH1pUNKH04UKLftYE8r/dCXvS2y
Da806001FIsaJerbdY6WOttmWuI+m1k3e0GKqp1IOveiwnT4lyvOmiZAMHPWBDbi
lVqc58Ee3YrWIkjRsPzHZVGpw3BN4+t9ax6hFH6i1gXAT/7JTXYN7WKWJdI8PjAL
a0jYDsfyaJHANFdxuR1PgbQx8sKTaTP7gytL50aXJ98L/NybTlq22BtiHGotW7E0
9cxpdF6p6RpMxSwY9WZRxR6fjn3U2F4/oKoM+gX4z9wg5f6pb/GTyLV+v579AErP
pSf9UcA0xN+e0CPxy0bjFEtPGCMLKlkaYplZ6k6iFE/1uTXgkPu9qw9XQRznPexD
gXLRq5o8xCLY+ON4/IiQvDk3pO39vD68FLt6EwLqFDOyBSJY/sn1sPpOstDjVYiE
MTxmltRLCrn+SFRtnXTK9WGk3FdCg/nYWzphsnp1/Z+T+2dJXgI3mZfC01wQPFwC
Wpc6S/HVYVzQCqcgjfUqhArqUoAftKaGHs8SUJ3ECa8SxeDdKY6Y0tq2HBivCMsq
l/BCleYzrlJa7pOR/HmCumsoBgpy/ORV4fG8oLHkk9YgH2LWmhSc8tfncqxLImk9
A6XMP8MDMAqf7f0daqF8oSWAN7DP5JX3nycEbJbkYAhcFhS54HmMhedRjoiKMLX2
Jjg4NFRwZiqtxBtjhOBGVQpt7BjoMV1ks6dNvZy6CAP8GwTvZFQrQN/6D6xVMfK1
9T1F4ZhAIhoRVsL2F1W0zquprbiVklIdVC5p701jbal6iVNLXR8pKoBPZ1/bJeBk
tBIAKiNQaF5ML2uy7mgoGwLFHuJ7GQfWPo1Ton5SKFoICqztrdc151G9QaRSF6Tk
nKjjQX+aMl5X+hTVD/KtFd8/SsS3DLuSJwnA9sEbPNfb/AGMTFPsL5l1JQC82lM0
qFm6p6STAQ3DT9dyFSWMw1R5ATylCKNhKBovo5mt4O3HdQB29US+ubZxfoecQUFw
IPFay5N15+YFur3CaQIKPo1ccSFW6UK225tp9xFvN7COyOqdCmM9YmnnB37vYy7M
GwegN+Vcc2aScFR1uDR9ckQk8ZDH/sI6uoqCSWHROCwzaum43p+DX8Rn8FuBsUyz
KVzCZoHq6kM46rBBnpwyRbco+eIK6FwQtafnTeBj8VPQi8Ds6rc44ZKPRZlrhKGh
seigo336cb3g+gPEv0RmOxfxCEwmVSLUowJWHGyllKV6EsCr9cE0wfqLRZRM2h1b
FSi5INZgIHi0DtgUeNWd7tUXQftrQ5hkuhDZ2rZjcnCvWbhLXW+9Vw/THKQxFxFR
KBPCnOZDUWfzO8BTKR20pgMcMkI0Q/Y469jG9FWGv8G307EaGQaKMwNMOnXJsO3Y
HpBdYiXuKBaAeE7atS/gfNqhxIiS0xDHO40Ph/48ShI9+KYmQSP9+YIRgaXUkM1s
2372e8xfTN8owInjjToUaeUeA1YISu2koSDU+61WD2xoeW4TVQQfwDoHnjS7vXPf
ktdJfKqJMMkPPOvL9wPUT9YGyDwGyMNRr4u9+qVZz+8+Y8bFeoVW20ObL75HCoNS
`protect END_PROTECTED
