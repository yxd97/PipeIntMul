`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MsCXQBAaxV6EuuxNqFE7ELTmX8qrU41ENkkxFeeu+LnmSh62yJ7YQYaQ39SC4PUW
EmI5aB0el5T6SEbee2dqS6NjGGpYH3QducNUxMdP+oTHS+mGCQT+s2NgaPwsgs7b
dIP2uxVgv4QAUK9JCybpH0nJQ8OBJZW5SoHj5yF9Yuk3QmdUMn5aNp6FbR4m1L5d
gclAjGk0WfpM+2xbanrIorXuy5DE0+KVxHJF/BhYGV1Q22mp+aI0Sh4L07g3veWz
ImxDnVlbQW7hA6WvReqctDuR6zrm/h3IrOiVZUtRIvIxXCIhUWkTaHUS2hrhKNMX
XxJL99tGRMIfUPFj3bGi1drIDEAD7Gk3rgtWBzAxyjnARF3cu5SKRz1QqG5qd1yc
35l4kyDE8vohOqAeJWFxlVYkpXAPMtEroQvT2+dmggRGhiAjT4by4IFR5p4SYDV3
lD+xn955sszSehF+5sQV2Ky0BGnSCi8FGJZSXv3Ruyx/PlbYJs04kM5ROZUFLm+a
ZpaMGwTX4RDTAouGDHwIOQ==
`protect END_PROTECTED
