`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/cLvNTBue/Y4OC2Fg9c/XTzkcflqiH1khRNQ3qsae8FbebNE55/ZJ4zuoZjv1OJU
/0mHLnwH/t48vLgpzWKe8GvKYxbMNDHC5HbSzJz86b+jUGIXB/70TDPiCHnRxJXe
5CBy5uHWG/XSe27gWk3EvjcGdSI8G9NzhoqX8+pi74rWvJJ21SOYxzaM4IgWdeEp
SeIm1NKa/XHIQ7KEnCbvpU0lkRzZ0r3X87HTRbRi2MGlq6kYbFKqRISW9P3mRXeR
m4CmKQG8L96ovQ0Xu94bcTO72G7jowYFYZBcpFWoC7OIio+s4Hsd96XVOl/K1xb/
1tE5yW0+q0EeBAoQrbc5QfrhAz3BIM+ayoLx7H9LrrSQybe34BPon65wi3HAD1l8
b1lTcvW1GLXr9cleC6d5w3ZgsX6sWvWjrgCEam+I6awzqyXnxs3Viy01uSCTYD2x
+XQP2jHF6lnGOSI31HgCIb0UURLu8Xquo2F2WWpsKaUN4wii+780JmNDoQ/Bbmk5
0OPzhULjNm9O45R49ChKTjGFSV0eUXN3VkOuHNSiKSy6bBUPHN5v6H33TzCkK+kg
/WBj5iZQQ3rXxL1oiKM7iPkD3XizDxG9cl53yhx4XB2UelZmmt3VR79+gIy0LFH2
T+EANMDTTFnZZ1/ikyUeSL37iRHEadLjUqyukEro2Vhg/15Ah9LvjXcYtHgm2I4X
kffF7qgtfGy1/MQwujLqVUW5UFxNe/tXlbalzm3cZ0iwt4onSjRrivqzIQ1EExSZ
qa4cCdFl5jAZQ1siaE2H4PfUKucOWjftSXcPMGtrVcu1FJJI8kh2M70NCgivu4nv
0Rghydl2NhVe3KwN5S3sccYk4rmKvtG1yDg7jm/8JsjhmcGCTzwpGPf5+dkW2E5P
gQRSeSdch0CXG/IGqA5CQ/L+WNMGl9EhxdbL9OPp+3CqKG50R+z11n/tux0lR7lf
m/G/epOonvIpR/DN3mwKDRtNriipGXcwOmaqkKWK77Sso6CDjjHN6ZSaWU76lYyZ
kiTI2V3VBETkm1eC/j+MpJZYv7VyfC9gipDUR4mm35UCpJvF6kOwz0h2WvFdT6D1
YT1wsGcnddcQZuQPCkBGYyz8w91Ab+56sIz1VdRbLwTiffgxU37r/APckHtknel7
/oSCgDt00lkxxKIlVmBmJAIU9DJPYOzxjXlkI2CGkPzYDsvh32XiJ3Ci/fdYt2if
gJl31xX2PoVgl/xM/4iRtC/3PvDjqkD4rzkmTtJjNYmBdl2XB5eJVQeozaceoS72
JufKyVeuu1CN5KvdECrWEGqHjN3rHKSygADU7ocAlj28Cb/HXiFIsr8NEUsOBGlK
dfY17TlDcuT3cCaBLl1Cs7YhTcSoBq4QjfSoE8Q5Q+Y47VxOtBd+QV23h4F0amp+
Zwpwef0vyjkr6fqMi0YhYWbUcdq8Aj/i+DzM4FyLaebZt0aNAhIxb+tvmqnrKvdn
1WvfwaPtAAiaV1cPMLxuJlK3zoK18dDGwU9IAEMZdDSyjyzt2oEUDoYXzB+QJqdE
VriCj8sazBow58jE9xoxc96zAdd1rXnW+PBU+yvEbKrXKKKnYTzXWf0xboaBrruu
ZH2bozP1t9/VrcvpTGsSPw==
`protect END_PROTECTED
