`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMYxM5q9zSVjHHtTuCkGYtVclbbxHcYOmsTov5qtpuT6ghg76EYlC7sp19h/Rvsb
royj60Tbi3O6mXOjs0QuEnaBhX4szdzVYnfToohkoooh/YYTO3n9PBaFvEqg6hG0
ND1i+jkpYZNBwB6rmz0/QqU1NKLCAuYkJxAvmPJhY6pjZfjPQ4gnHlRK5s6wep4s
+7S9fgwif9+gTtP4oVo0WcLrz4BO1Poso1yBXfJQWvsRqG/xZGL/rYmeO2Tj88jw
Q8yU8+vuChlO6ch7xgg4GpKvbboiOKFBYqgdsZ/1FJSfPBgXo0ONplVJ8qbFXFyr
VYrZ/JIV3Ruqx4BQRN+14IYZz3uMShodHOVc0uklJwH7Yqap+R8y2sPrwAaUHfSi
160xUA/TbANLFOQYfZVsu/0j/XdJGKl1ZBbC9eV7Z05UHuI3QtdRiPcRq0/ilZMb
c/grYj3rtNtpw+axYwmMlTsFur8RyCXQaZZvzBv6SCgiioWWn/NFVruzbNQzc2ky
0EC248cQ7rcX+5oyaovp6vbGpmzR82u6gCFLi4sAV/hVKM+6c9zKnRi/e6HqCRkf
Xjyqcz8mzNTFu1A7QuGKfl0m5FicvQ2i7ZBaH32ReFeR1e0dJ9IFt/Ms4J7egpde
cgdc30NxGjxLgQySQWd7ZKGTrjSGmBaPn2IkENW+MaynjsPABDsdh45W0mfYV2ei
YZwPbXrYAjoF1m4RBsssYTUJZQIH4aKMkPhxUaUUGPrUpiw9zpMlVz6WPyGA+JQe
tNPh/LFLTeJ8OfX8E326+YSZqjxba424Mi3za3dmiVCHMFZnp+LMnMC9QWdyfqdp
aT2yvVWAGb7ORgYeu0LLZOQQi6LkxlS7sUvQPGCkVPTbgUg6mE+7Duqp6SBwdbXb
POc6GRTZE221I4k+bKXscA==
`protect END_PROTECTED
