`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2Br9GxQe8lKf05JqiGXRaAqhQ6aP9fD6aieZmETyGf9YkCsGLWIpoe+mP9yl6B9
yzxh98b1/hyYYKoHu7+RB3EigeN3Q2zy5OCXre4PTzmUBwq+UHMe1U90VF31s7fv
Ws1KYLMMCzdXCGn24kWaOGlEr2lAGxnEBN9v1fXdEtK8FvsE5eCuoMYTB0IPxYot
YDaxm8cINkta09KteztUcYXbJICWEOXzUnGFPJLH8yS7lEARyFfn4p90MnvS7C+s
Ks+VfiYhoi09WY6XJAwMud3Gk53w07JhlajDExPv+a6z7bqXqRx2oUbbD+6/kyGh
Cwm69p4MLTaMwdMl8Lj1D0hh30Llbdig/ByfThJkVXvp12wj8jbSnrYqvgcLSqgB
1S7grQdRhq3bDoKM0f+hSZEoCRFXMIUn1Vqr6lLgSxc=
`protect END_PROTECTED
