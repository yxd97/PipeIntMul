`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6m+15ev3RRyouMJd/fDiht/fPwq1Qe8SXhuaU+Wi3jjS1lOxjtVgsGwQWaGjhKhh
VoKDf0SAMfFOYL7mqKkVtzqwyhz6ZP4S3sYidtondtmfcUOjmjgDgc1YhfAK8Xwv
L4jqLiPo/lhbpkd23h/5cLmvOtL0xyyuYFfJMGke2Nwd50UEP8Wwqi5vDufafvpr
jhIscbRQf0EPaEyHuMK/JaNlU7Sba/qF8XDuJmQnRdLFK3xP5zB3VhkSpODRqQQK
njDnx1vwsCRv1rmvcuiVXo82vieSKVDsAILjfO1/q1K4E910nouZolAJj1jC1EkY
c0KW651r6eGL/kXi1fqeVZPZEW9++ZZoqqS7fL/JmpIU8J1N2R34/8OFSmkoC2Jg
+LrtqMSZ3Vhnt38hmzGizHV5QbXlpDt0+kEYYge7No3eH4zDuNepapU0n5a2PRRs
sr2xHXGanEtz1onrgykKE9u3L29l5HT+GZ/ix4wZLcHgP7JLAw9ldZCCiMYgvMMn
A0Kxc2qzINN6sXNEpM9DnlCNuBNbbuCUWqviy3rokGw1rfM6Q35vvypLDQYtYTBj
W4qC+lc4SWibO52LAkqQjw==
`protect END_PROTECTED
