`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNFip7QzQhI1IRPvAw3eica7qE0cVAanZD66XFWbP3woV+Fkwfp79OoqfDUAEgAp
7XhLE4u4zI91UFVHhImbn06YGzC7xWCzdB1N2HmB2vthjWOlXRvAQBfAT67Ipa6Q
4Vl5M/HdGQbF+/WcVRUaId+pA1yojSa7ZXYV12biUC1+C6nwfjDJ7OpRNgfK4OE6
8sX4xaXlOu4M5dSq/aA886vrIBxjAJbiOdIZQO8ll/vE65ku7jlEB2spM8YHdHJ7
gGpoUZPmcvxQgEYTWzUrwA==
`protect END_PROTECTED
