`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P5gR3glPPVdVimOL6Fo7souRzNToAdl+v7YPwOFROCCEVrwwQiGOOZNTbj470+K2
qpEbYbEzwGPBeLgLuUZiWfaKPOxG+krN72LbGZtTMvTvRNQHLgXVM0t2vtuaYKgC
lzyYRHIUDEaA3/fcBZoxBxv8utMld9eGr6VqToB6te5ArkrKDWhkm3q/BcrpD5Mc
55Xwfw8h7sLXobd8a2dyxe9siajnrPCqlDB84IosdM8jFDrUUjCoWOlINocCReX6
BRRrD3U4n4kni6kgtyR31iIrWMXD5Ng2sJmsq+Lja1D8MOuadtZxahxmLZ/5hZ5U
qV+okD31AVqrzeV6WzPVs7PsiWFjEBun2ip9/oORXNGZjy0vIordWVGtMegbdvcS
UUyiGzCKt5I4hgQzIYY+k5+wGzS+ysZdUa24mIE+TnJexOfms/iBmQYrNAQ2w3bm
t66+QcDNjWNrJZQyxZ+Dz5knvuuALbTeqvqx7g+NPCaEjkfLlZorJREZ1Js6uLId
APdtV6A7G3EDaYr9BI3Tew==
`protect END_PROTECTED
