`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ean2VDqE1UCrL3bR0b8FGp3g4R26tg0xSCXp4ORXjOyT7FwUBDgfbQuwbr4tWyIx
TUOsLF48Z2gxpszu3YhO2m1KJdKW4IR4HXAwg0fThmLJjuUGlRM35m4MPDyUXaxy
GOChQgzXid4QibMMG9tT+Pt2M6a6Dgk5hcdFAQSYSfrudKXWsLmtJGi8td0Z9bW2
abzCFd0Lt6JVX06B6lx7nsi4hs3QXZWIxS91ZjBzdYECl5B1mlQUIeRnodu2y/cF
MJruGeJ/IWfajZo/mfL0OstNjv/7wSkkhuMz0Bv83MSIXfAk/EFdXtmyW7ITsS75
0PPhF5nXvoyAz0JC2ZehDXbWVE+yTd3ruIfa5frNm9SL6EFtf200P862WPH6lRpG
kXV+6SLb1Y5+HMl7Jyh7v4zW1VDRLxT1SMDMFsrSfEo=
`protect END_PROTECTED
