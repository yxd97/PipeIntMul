`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YMEEREae7QNVCfpq1WMplKgMFoMdM9MAOw5jc/fpAZPn1IVEuFmwFYHSXiqiPa4c
tCPXFjsogiM00nOX7GqDANOaSIOHNDY0UKYXg5iJAsF3CHMhAHaSU9/50lxOjniI
h6/5XDJppEoN5rCZtQsnorMPoqxWtjmzl57utfCLyne1wKt/dupkckYBJNFBGQC/
Y3kiq2r3YdtlEv7RTrI386LoN438gg5FHQxLS/mbaptEmQwCzc0m1ckyc2P3DZ4t
L7thed6uaS5qUbYNYfioCg9at1XQdb4Ztz423z9RkZCS11mRo8kl4q/FwxEe3GVy
9jNJeflVIMQz3dd/UAv3hY4uwtF3S8e4QgiPlWKipwMsizTW++K2Ef7Kqct1BTKw
ACRT+/SAi9T3HZxt1CV77xk9OvSOLNJb/swCUySWu7A=
`protect END_PROTECTED
