library verilog;
use verilog.vl_types.all;
entity CONFIG is
end CONFIG;
