`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpyQBek8YLBDgl+JgUBSrpGCrxzThLOL8sUzrFVgAfr4voNl8EyJx/i2JD+5cL6y
SZ04y+ppI0nqaLHES/RYMJsLfJCUxRDgvndsyr1alxeaS6kD91cuJbkiRo+ZJyr9
wO8w+0bYsDTtoozECZ2kgnT662Swp3xkkncGWdArJ2IW1KL6k9JwG2eXN34sZfu9
1PvQ6y5uKflXlo6pBqYz3NWlkX7och7Y+RzVgGihEi2PFUmU3G6MGnZbfvBsFv+6
YFcShY0hGvlncZLoXW9tqVjyFvwBMskhAiwBjC8axXyWZPLhMwMDA+tDrLyvc3E5
Su6kTRTKlbdA2Bg/bByX9QmT72m35NWYLhshoJipXypQ2aKrUaGMcDI5bnWRcyqm
OkbjJrD0if/13xzGY7UUvb53ncskLGHZu3GXNQcf+xsOlDjNNyuDsBSKmSK/rxjl
/+aAafvfTP8LfGctX9eOpkgN8hACTqvmMwKCMnx+qeKCymF9dSWvCb7PoJyQVqf7
CRA42njKs/HYWORCw5I3XRLv9h/Yv+QLQmnaBwFWziWBuWpD8oNMQxJbgtO/s8C2
/H5uUFPci7WmWhFxLITtg9RDHarN5T5hIM1vV+TTZ9tg/pqqJqJzUZIHk9iDgLRr
ejox7/M5ljjPPhW2v/6VYV5b9KTDxdnrjskkDtiZC2HetRBK6Xgik4ItV5Y6dC0q
9X90mvWnN9S8Y98by46t+sy+ABsOBCsMjbuSQ0PeINGw+qJqRHOWPJLQE2fkFrYP
LgvcB12S1hUWN72HNl2cLGwrQ45yfXcUu6Hp9sbb+n7AdftRP36aWF5s6/bmzNPq
+fUbXR31vhI1xxemE/0vF/hiGbTyqvcAFbtxQBjhc2nVVk/XGCxkkud4aE2HtILf
+a4yGNwPtDLB7MZUYdEySwl2CHoo/2K8OAeutXQBZKRvVpnAvwTfiko/U9GrC2Ix
+DoHBWwI6K+mhILXhBv+el/ZW3vz8xx3zuyyHP1iDoFPTEc5Ru+gzUWRfesM+Oj1
zwzPHbHJOsG80n4RgilBDeF0dItmZ1X1ts3Dv4up76e/1o/GrLrSKe8zQhmZuLiG
56WmruAD8pYgRLrfcXMjTVMQKEP+LxKcO0QSgQfJKU9KK1+2t+//LTCv93tXa0wE
4JPr4EIs+G9I8Hiz9RUYIal5dLTELKOMS4jgsGlyh3DjLEvp1iD+xiCceVOnTL8A
uLvmRxGMRADPvd5RT/+HCcsyvhZJoLi9+pKy0G6s8Vfc40VfWz3TPbCaL5GdVNLD
1zTAnHmT94shcB+E053N2VklzVEFNCqq7RRaNm5Y6y1Lcsh9bP2RQU3P1ErfixEk
fagOC0lPftYHhIZzUnVEmyUXsf4W91uza/hIUUrvaJ+47pU1eq2g1Viicq1faxre
fOpVG+mLKS1WyxvncELbm3CuzlvXlHnLcVyNifwz6DbtU0tXPeK8t/sVDAEasU93
DwJxK2e4tFSWF6FzNfQLz3aTIdjt1PFeha/xf0GGjQeQUnAqlWaynhOb7DHoHDeZ
hELIcnIpHzv3HNtKaSG8n++xg+0pPi90Rq4HbDU+pdoK2WEP+lNMz68sbgh7JNMY
`protect END_PROTECTED
