`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZaeTYEHNa+IUt0DglrsZ/6h+3szE0Fsk1WOwQPt7uvGvjkrTWqhMBFvgNlcrkqxh
MoI97fAOwR1S8V7jAX2tneH1NRe1vu/1luqw9pK0UJ7GL9HSfZ1dxhOPT0Lj1vQI
wncR/IAYQQb4U0gRe5ODgpqbD5RcIq+NhIitN32bZrasvobgL6oESKc5qPn8Z9rl
n11bbF1LWoptSXS2P6mcBiR9CKGpQzG2DX8QsthE9wEISeSbIEB+LICTfzAaQ2Qn
P+QV5QsvPN/31XKyiN6d1yKDJseaTzU6q+xXFi5Xkl9VtM9k3GKtirrgcRhu0W3n
ciEg627LPBlNWSMdcZ7Yv41xWX2VjDnGkoGT6GZzCBauXtpPM2rJWzRdX5zPaCfT
nj4CylAEjjKvbK3WLANemuzYqRICBqfCEdbfbdqBSx4I03G+cLf16f7gr+EU4RjC
uBwP0odxL4SE5Mz7AwsvVforzLryuOlY2Xn0X7X9QuBRafxYhPdws9OQ23TJBwJM
bzuQSM1YzBF6FggVVhiJMVgN1DXqfRjWM7G4ZmIFEwzKJhXtMS+iZLIjifWA0eth
jrEueFzg44DNf/bmsCAdL2Wtj6s9woJM+vd2ci1eEGpiarpNvJ/AX1LY9ptmNkoD
qfWrjXHbBie11lZDFReSxWmocxLRIjKKtDh84Kth+ds=
`protect END_PROTECTED
