`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lzkcd1sT4iCkE/m5+4S8XNXPj4jEOLZ9IqSfYfASmyat4UIoRCA3b3iE2JpBJUi/
FpU3O/f4nnrPCVusDUjaesGnDNnrwVz2PfTvNs1CpyW/evbXU7/jfWmWW/2iL+lV
JoqnVVDkV1VOwfImLyIBTA7ZM7aJGckOlKPfYC9yTfwwbdGFFXiivm8H9pvzKscj
A4vh2e8SvpravakFgCTxwQF1mBOqgzmqf8QU05EgxDH9Eg6Fw08shtLrTfLEeZdE
glUTETEWVHE4d8F+34IYXyfBl7Yr+IU6SAOpn2zpCYo3mSmcPwqS88rNrrzyaTKR
s3eHTgxYoNlseBGJEDt+oX/H0vBn3lzOYFEAfzsPCPPa8sLSc8cuHOBTyqQ9F50g
KxZe3RsG3CfAigQaEgKUADvL8gmR3w5Aa85uRE8Zow80HjQb+eWZhMvz4LQNIhsL
`protect END_PROTECTED
