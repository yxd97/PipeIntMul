`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3lClhCSfvGEPEJsTZoOuAKMEjCJ6Tr+YvaKv5MzFk/1QjKbJtgSVj2it2Rdb2lZ
8DYy9kZqXA60fQ8+GH0MLm6UBcmT4j6zrr3tVW7zuawzrum8vaWg21hUUv9jNruM
K4SnePwcLX1PE7LM4m/zPbDN312WQ2BomCtlHq2KnJ3tsBTtHadOuiiUkmHOf7Q7
0icDpfbufCg2ikYOqqpAQINr3+GuwAHWuSUffUxdxxJDBiLSHnkjiwdfxjkeVPoK
crxMhvRehstxmsYGhz9tNzgAKugUbbnld9dyDWa55HLoOZctMq/pVhHUIRRLiRgq
zTpNBNz1u2uyjwNLIw+49Ayd0xZdHP/8Rfxk3kfKcBWgkSQ92SUrLbRvGg05WlPF
gjPWP3eIq371Csw/gq4Tb4TqMUaOhxK5p48vz385mes=
`protect END_PROTECTED
