`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CU2HDAalncyhqaVNEOMYpNGUMtvauO9N6+wKdhvOqEzcdS9ueDA9NkY4Ekic3nQf
i0qn5oGOlo6kQBs+Wl+ofwaVD8ZYWQ1Cx43uTPTS7XaABZDDrmUX4+zIOgjpmquc
zsDtoeWjl33eAqCnN/F7LcQjw82jBXAJUw+WKt5JEbXNlITHx5XIIEVQTNKz3CS9
v9yw8vI0uMbuKcOBdqiTJUOUz2IoE+Mm7d0eo84mlAm4VabQKuB8dmFCzztU+Lgt
l8XCWz50SjE1m4A6HD3PHtLPZTeVVVYfNQfd7L8oP3iPgfwoIihVJZu0WInbKKq6
EWixWO2NWdO0iCgxYPjOgg==
`protect END_PROTECTED
