`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MgMnPABg7TLhn2v8k30FurQCb69CZIaGon3Jx12ABhdNX6cb7+orOpYd2GsS+ubk
46pSY/Mj9QpsEyF4KQJQrpNQ0aiyYzm/HZ3nW5AIryW33zzE3tdp648co7gp0Dv3
RQTk3Y1pYBsuSPsg8v8MO0oVQ5C6fyshpgdzQYQDVu5pym8Ce4nNVqLKnwWuLxB6
9GGRViQox0W69N1mPvGHaI5M32JcJnarVFEL3RDr6LhmBdYadK3HEPzF7MxaBn8X
RR9stBA9+FhgUYNnseanN+BsppjduW1X9xQ/Ijp5ecYxGR4EilDec2JzyCbDhk/E
VCKbJSRWjum8JH2QjOZYLeiu2dGZoqnxH8edA/gnfcKDIyXAFm/VE9cIa7lpmMmi
X7me18Quz6+zKQr4Ce0xjp3wVm6bswgNGw+t67RgDG1iT+jz1f7HzHltnQwQvIuL
lrmFTB3usdEV8X0CNQbMTlamgRse6DlU1y5oK/p5Gq8Onlc7hHz4N1kxsdTu7tin
DfIBWlN9svYQYG/gLIEuPCJ9RWleJXb4uD+0Zq+8VXY9p6rkHSFR6/Wq01h7IWqD
BWe3jG2AuzNOwPyUs9hdytTbQ2GyShhAyBb7FZwzbSVL3kg+HQwi9xdEhzydkVcQ
KwS8hLUt3hjN9ulPXcZQJ6ONNy2rZid4JVYPNWdapGDtm+ftJXBBghsY9kceDRtj
WO+c5jLk4aS/ZJQxh8kNjDBUzGvPKksvb7S///3can+SX2h7r/QuCmPZxIhvCBDZ
GHOWZBCAsbwFUxG6LvNkb8zVSXjhF4bO+G0cUsO2pJBAQmMyW5jcqXLgEH15g8+7
TxV9U4nVzT5O292s44YylOT6vCjOax8svt0HqgGekKl2VgRc/+426S9VxrNURcE6
fRAw5ZO0iJPcWy47QpBW08ZivLEWMvv6BRKVdmOdEwz9D7/EVuyk/+VFFVPRW0y4
6r/nsXUUM6w0pzJCBg9OtL9k5EaHXDWul7hu6bycylg=
`protect END_PROTECTED
