`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XmLUjInnkTDgkFlCeQr57zf3T7V+zZRqYZ2zzNvuoFP7jtiOM6RxnIHHFzj+f3/W
4WWfjh5ZlBDlg0r+weyojpmYoH8+2Yn8CaTxW+1DBQjV6LlkkvSiztJMCbI+CDMt
uX6thwbXWMOSygRRGt0Mc7jLe4IVxI6KdYOr9uYAU7/VagW4pG1OdsstmlZCA06U
xMz20ltK+HGJKk6SXV4dhBabj4X6Kuq0t3scx61jEU7i27u/CKlTaG20MKy4lDfQ
nJnb1ighEOUUMkndsG/aIasUOLEZZwu+xizSmtGqU+tLhUI8I/+8zOECAUYYHHob
4G+O6iIFYetv/1MIY4Fg0JTmzKDVG914qCf668ATz+38GBJQVSzJNkeRDN6AGd1U
KCHXqfsw0YHU1z9E1LnyswMdx4UQZAJZ7t2uALEtNP2gf3HjNLhcrp+cPP3gdPhJ
`protect END_PROTECTED
