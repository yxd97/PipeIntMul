`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QE83pKfcZE1VubArINVMdvQhvJzHeh80gLNWGu180LjfYlKp3TiV8Y8XYoxSXiDw
1dnuxLB8FWXOZz9CU+EFGL/bxeVc11PoYe/TTTR5Q12gAvqNSalbyfj+B+tiQfE/
UdCpzVagJaThAVnIPGVJv/XycVffOI6tjbplGAHqQCwOA39jkzGXON5Tr0X6/nWk
yvogvluHz9AY9yDABRMQopFK76HjO9sFI5DLT7zzg2whyHlBOGXUiAnIdYUWyFtt
pc9kcGWPGHgstRYVfDlWKjY2b41D168NJ4yFwLvpUlNV6z4buYBzG/cFuhNrOZol
3BiOcvty+pwzzhEDb4bgiA==
`protect END_PROTECTED
