`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z8hXLbGO83GEX6mwqYv19GIfAr1cnUtgbnR9ykBwWe45haT7EUhvI+am4hWRfxkH
fKXkMoEf+XGbmeV5E3TNgTP2jc4gJKPR4Rtkes7mKeGmfiYBM+yA5UiwxVLUoFcb
9eiIz0cUHcrpr2JX4y3U+5uUkko3ehghKcuQkDxFceAi+NiDYY2SDI4P5PGRbszo
iqx1XGGJ2VNd/HIlq8EdzU6WDu+TCuHCgm+mcZEBZGgcm2wp7ZjveTAwJhBeOzX9
l387GYqxIqPJ7bgbNgoAXo8iwkiTJJklZLjrV5u3Ua9Z3+HZYOTmjxUGEZPiP5L7
yGfPdsHaGY1vWFohEDdNLuPmItaj/lulwgR0mJCBHqatkdWn+ptQt5+ng5AZ22yn
gfcqFwNsa7Et0bPq1oLuApsySD2Vvm9NpFcmnWc7kvhR56UXtU/nwWkEVwQU6Zlq
hIrjZtzX7Gi1pHTs1AfWD5kYZrWQiOoOfF9iIAjdtNdO5uqyjL/XSwusaxPG5Kgv
S8BSZZwt+N8KWn90Jum8i/RBKEC5AkWTOZH9c/c/zbsxr3JK2Jt4kP8JQlihCeBW
Gn+PbAKIRq6k6POP5dcFMBjeFrq1krwjZn//x2TzgIWJhxp/vF9xRMVo9SQOBvgi
H+vGvG6siwWswISAqvFfUcDiH7RdDf3PIru6dRPlsmjr9jyQEN0M+7QHHvnkGRo+
E9tHQMuOE4gF3ZxSDSkPc+bTVMoPmSqN36emJi9DtoRr3qMHZTCXVnGwviHWHhiP
OfZfqb1kxsVEtsU+XSZJ/FRMseEYS2ValL3XHXlR+ies9raZEw7tK5+/T2DM2EI+
8CDxdXbYi6LdhGwhNK0jFp8p15Bq2we0r2hlYr0mMbjeD+kc6kemRaKK4Kz3OvAn
DVwuiVkgPg/oefR1kswT/dWAY8NrKbe5dOHjzoN5V3MFPdxr/cTo7ynz79OXX5Ny
9YnyaylGq1QZQgFKzqlbf/cYBikqco02JD/Mme2uKQafNvMdzQNNjQbZoyELLcEb
rdfv2oPpgfedCqSuSLZ3U6VwqDV3//rqPSCK9W3dpTF2blss7qLUAUWm4HHU6CR3
xr8KrcsxSCDA9XvfZ86OyqLVG6OkRk9ApGf0bokca9w9rxgeTM9A6mK46POQg/Ng
9zGXVAhHw+2e0zzf0x4HOv980AMUPLpmc+Jy5RK8wHtbQu2TvejDpiCjK6nkM8Ft
BSBB5EEoM5DxrdKb6S0uJCfegyaAVGSKANl7mhURRK1vuDaMr5EWjR9W5CusgNBu
IGp8bHMy8EUGQ+RanxH8xVez5iKdsxIbUtsH3zLWc6aUHxo3lJoHYUb8Cw6NsVcw
OVZBCu82lpq5d0bv8D9Sen7nCPtJfjL3zZImpbsNksrFtQn9D7vCVK57pZTb5S08
FAy6t9Rt18eFoNUJ3+haKv9L00v1yRrHal+J6GXL/YCerD9Nbfblh0qxjoZsTQUi
U+hZPt0SJDOypuwbx1e5/IUpEjcXrrziM+lozu8S0+kzpGE2ZcQN2OcYqN6tgmXc
SYUETAgtJGke7GmTL1Q2/ITJPVSLoZXVbqYH70YCO3ms+U5Rf5BuSM6/TdHKgVoF
O2ZobP9NEB6q9iVcA/yg2n8ACvIxcMAlV2pkbsvBQtbqxI2eqXKzY30UEEIY6pYf
kK7xIf5oTV9P8t8rHu6TFs7LytIb5mhoVUajLyGPcsd0p4PsbU4f6TsLrMRhG2Ac
o11E8dkia2AehyFvxb9eiBb5SDwUPCBJGkePrzguOraQ4twLh7P0qq77HcAhZlju
niZqL2nLnIXOvYxu6fdpIWPt2ibz0xtYcdxrbEBdr3mmvEn6tZZP60nAW4wNJwW0
l/QiYvI9UsHOq1HuFlnEgJHLIsuARov0ht34J9DbzGx2cvsM2b4SPde22l3RC4im
Up7FKFIMV2bzmqqQydY/F0j6BaV1GnR8K6rRWQAl5vhk9Ib0/EN66gYpgvhFNxxa
g4rybwd7Vo4f9fbJunRz8uEha9/wIRNRGw+Oub5r+PdW9NTw7FaTp6penO692jZR
M687z5P4zBXMc0xBZ45EaxyODUGVxzmRCeZvRG/eSFgwoagLlL680U40lMfmFjZz
tRKts7fqdcGOrvHCpI0UuUd0kh6HG9h5cjv6nzZz8C2dwTaYQ+ZaWgsH22UorKpP
VJSHrGnQnOzZizQWpUyW/GmQGfsb5vVVJ+47kU5iDVOyTnsvFSgFfw2edKR8kMhm
MLCM2gx8yEbMAG7m6c1QE7kLEcWckzK1hYaS3Ilse/U1a0rqVTiS7i/IXsSI/wrz
5y0vz6LfxtbjPIQcJsMayh9AUGJEGdKo4jivDAXgACFwYi2nPcUnDHt5mXRh1GPh
wR88NQG9+uEGvfjS2VzWYYGD3/EBxhggqRyqMoDDj2GXmMOmTh14aDhCvWm9wXXZ
wDHWUS0uuj/id6ABDg+L+0CJ7IE70FrWkebGDHSLkyc+5561X1hw65DFWlrPuTYv
HlMorF34aIYDDdQYIy51gB9OL0Mg3Kgj+4Q8X+nKu4ey90Z7tKvr70hGYOzLQPXS
ikYYHjwSzNgcpfdCqKg0dz4lRMpZ15NQCEf0uDEbGyTd8JQuTot+pHB6cBPd8750
KiBcII2R53hMH9lxXnpfRYGqWHsxlDcFwXAFr1GZuOm5ZXd7Cym5QLG78EHty005
sghBETsM4ZSPVl3e9EBnshiulCfKNsm9v3iHI1a6hNHnYarVgqOBnW6gWkbnRlDW
a+1fezltpF1w/aPhYYs6Sia6K5EnDsVA+UgBWna1tSlz9G8OcI/cIhhcRWc9YaQh
KgWka9nS5gICNghqNjmblGBBKj0FbDuvAhBgr9kQr9AB4CwPnF85bOhM/F0LTcdg
m07jJgguXo9Ip/qnZ8ezSYUbhfTXZpoT5SzCdg422kBeBvqqRKB3w+tW8wqiAt4q
xCyJtSWc/CKBP9368wrLeEPn7K7X0GxV6qh3yA+PO36eCag7O/IIdPB39yhLNGGS
pgxPh/WKD+VWH8ceQRFb81MZB2Z0knbYNvmW2owWMSAMFv6bBc/YHrF42op0ZmcT
ldCuKMHTJ4lYXLYUEbrKLtAgXw4nkb5f0yjk3fjYgiuMEBOo3qTxkZyVzPm0XeFK
ubdzCuZE9+uNiR9tzrR8jL81iXuNrHgoX75mH1g6O8qJijIifxORFxffVgum9Kzs
Cmjh9zDERPQmDCFK3Cv+LtwkfZ/o/xMw3EvS6z2OMCIZqwa8E7DPoAIaxiLTmMot
fVB2Tr62wVrMKi5Q+6xhZKK4pVq73zr+YA02jC5YUhhpzLNDWQlgmNQMQVowYQS2
h+rx1CsLnwxap0qaTrfoyuZEJ86gDYSlBKce7QAohoQmUX8kNTx2BH782GNT09jN
sX6y5FRYCHlcI9M6VpBZR4qAYEZhJzFl21sMhz88Y4OEX+485/vGpy9y0SyDVEVi
+0FWgbWWajGB5dKYocK7MzrIHNEMANLcyDOLr6E5xKKobCnn7b8bzmWG7pDOhLEL
qOxNJ8fSFOoXNKzGH9W731iPjK9JcbM1D8tVLlXvZQA8SlblPQ7p0YUEIjEPwFkr
Dccdu+LKLfO7m4xS437RrD6FIP7vRAQSELkdfwt6EaydwdY6xrGAirqHQq9i7YN3
5tniAOHOXvbSVh0P1/skfCFdNK3RlmnkXL5J5vNQOZeU1b6sVPRglSYCnGk9B0cc
2b1AxJdxDKRYu3ClcbbDwoBGXgxuHxGcnWPwjYt83bERby++0kmPdbJVzIRT4547
p40MC9H45HzpN7Xpc36THRLoUe37/AlD8ojkLHo+WExOVayGJM3W0EgdBw8FXziw
7eAm42p4VqejGaBSpKAgXMv/+2MLtpoZr8l97XG9T+JTRtiLLYaxFyhOmCsm+sBX
vPR32xTn3iqjZH2n5LUfgtKSChLwR85APncTGAjtZ5coJBmrmk3lbuz8ZZYxeAj3
+Foxn5xWIP89aq09sqmoj/+8WJ/2XgIHGukQ75An+0UvhQwhF5+SNPcYSZaS84GY
g8UPdmrYfpKI2NkE6LjIvK6UmVVSWjBsgnAHxr7W/c1OZGXc9mL6xSNIUNOSj1qu
OYHauRefPCPED6W3GUAF6ncShrstHKa6yrHQGh+soKpA/YoQVI7QxBm/doIZmJ2r
hYf5dBu8buIIsUOmIvZK8/LR+5bvSzMOYj8qsAi8E3vys1YqFrUUVOBTHLz6UOk4
u2V1Mkspo0K+LH3eY3n2O9DgBWxlUI1lTnfmA2T87ocf71z0lrj3FKTfkFS8moUA
1NLx/PYRIisutAPO4F9Yt+GqaRmPqv3zgiheLCBfB8GWsnAeOBcVhqoZi68rYwR8
j43vk1mhIEbqDKaaxJUC073ZK72no59eZeb9RgkNHE87YLBjJGunktiHHq4r9KYP
qTJQC57OjrbOpz5Vze+AhOLh/cI9WsgkrlbyfVqGFyMQnxdVotDAYxg0EuCYwDqe
BGJjqa9M4CTkLQ5bkBp21zsftfYQXEXGmZm5W9VEmuu/XxaidbTz6xP+PHn9blLA
DUeax+TlSwZ03kg9nCw2S/utXiH9sBZgtfbThJqjYJfFA2SajFiBg9Lv5kDedgnL
fueXNLJCbMADWzvgex7Lc3i12/YGIWQwJzdiEhwKrWyW+VP45bZVKGcgHeF9L8yW
4+XGsXDwNHx52V7fPp6QLuLOeVx9B8S1zl22c3ri6QM9gHHAeYFvRDzQvv958t1t
QCP9CdmQl/1bukQS0J3h+cAR9YaG47ofsH89E6JlU1Q9GMkGy8APipZDpKSxSVMt
/1DIFSVovHhnvSXXVkovRiEbxhIa0ToRPi+kkGY+c72ts4lG6U4Av2SJr3S3Oku3
cAtWhcqd+C9osQKQpewOdA9q3SQ6dKGPoqM4r645CH6CSiGydf/LjljhmjSzkCTc
aU3Ell5j2QtcSCIHdhuK7NKT6npaBOUjzHjF1v7FH0YlGlJ7IdoZiR9dEF7kl96+
CPxlcmyQZ8AdHER1B5RoMDibNiVrwlSqKaQ944NvPc04GrKBu2iG7r0Vs3ZO7Hsv
okvt5QY/HTb7rvPSxPoQUYilVIgX7EDEzJwL8nB9mr7NAODH9tv0sBtGYVPMzp9A
H+rwdY7ksSbj3SmUo1ebvO9wjEjSJ4L/DUYfJSe3TRtbpbTZyR2ttyn+7ntEipDm
vL5NcNXSbnTV17WqXYai+RrDGLSKC7zB2S6O6zsmbVJS4C71N2WFHHxAazQbMG5E
j0NEtLY74DxgBVSdY9/3aG4WgvYDkqSqHPvf1FWUUJS5NJUmenBDgMYedXZMseqq
PN5ccanDkQWrs5oeoi6tLe4DVQGqHFqmMCLkeFOkXwv4JZDM+KG3Hlh2lYyxDpdB
1bsXnKRu2/2KofmwWHdqEI9X9VngKjuPcTXTxxtxUUEWdZfiI1tvXEpWBKudGoaQ
kHZLJvSLJCqrqVew8jMNSZVa4QRPeeP5KnWxs6X+p0E/qmjnhOQNbA/DzQnWp7bO
b4IV72idvUhD+PO+989g4/2BAUu5IG3zeE7py9jNnsh35K1H+NaSZMMMtLgqe2Ap
YrlCHw3WTAVWEuv04p63+KFhLV7VjyK86z7/ddJaok9OLfGW4qUvvu6paiiLCDhS
A1kRfnHBdKWANQcvvc1mx3TUQqPnK5hIQuTBQ1+3Bx4KicdkzlG2p8ug/9QyAPPK
4PXMMMOSzvdoetQr66kroOI5aDT9EpTVbSABFwOQIYgoYNiMrQlcTLFw3TB+0toB
TDbrFB6uOGGmIDPMIziu4Y3ohwJxwULuLBRhR95hcLnTYn8bNihKDEc+g3voyAyl
Rl1zoww7dUAnMx+yNGu5G4OZPrqkaos54nlPo/minCr8tcmDjO7ZtnGqENCmEAou
vJWjJPtvnUhBYYRXDvTpG65hqtgE6H09NOxSn0+qgRmTCAMvmgCYgumpDQilb5xe
kYqayLEvbDu7yDoexRLHdgQqU0mnyVtMARnwHjlNnOkMF5pOZO8knxtWQ7Z1NmNq
Zf6SlnI0rKciZ6IwGaX+yZ1Mi7CaqiXnsaOsFXIezwsa4D3un5VFa6wm4dolkTJY
ReNDzI1E/nc99t9v6cNINzjqGeZISu2IE+NXk+AKzZ3LfMLO6k9Q0bXqB+ArAyqk
KUWD9DzDtDgbjVdWzbrEziQBBiUSskHbdvaWj2GLnL9zGG7ImAvt+BsIXEJ/S6L3
bqFApJItTa5NItbSMUHAWWJhOSQYIctegYSQo/66irKiczVe/jcb7sGhGm162DFH
8pzQulI7injofLtf9TSdStagkfhOJZ6cNsBmztQjbu2lgMjWU5+rITqDeZynCJ3z
p5E99cdkD2LZ80dLp6aZQee37XW58Xf7K8v89pCa7wmSOiiSpZBiZfhX3wESVJ45
+a4JsF4jHCygLh8VLA5FQPEU/bcSHZmlrM+bK2eTIv9zYl1LEzyXK8LJLRhyLrJ8
uEPoNMyBe2EWQAxU8jpf5ddDTrr/vThQolVOOV4mJuh7RaLAaHzY5tUQcsnXxrqY
mMDvylAxYppD0zh+F8kRNoYsirIZcOPN18Osp32ao+mlYYqO5bY66LsEqjbUX1/4
0aBpTBwYHwHP/EyBGKzCthYXRjO8fGxbrntCEpdBNIz4se//N2qehxtI5XRBGaDd
GZexyupI8J5NFKaJvTE3kBkW/og5co1octunyCAFjUVzWJ4Up3OM4cXBPRqsFxCw
L53MBSMdABxMOHrjnGfomJpsb/T0u5WYBx+55UVtnTCbrRceNIeJLYOr7WlJEhvB
0weKPIVcc11ihkoZDwYYDjvc87p6mO2NMsBMK659CqSWcTK7ZCe1/Ok4hsSjJok0
VEWyCGD/19hvyTJAomJZU9cWL5pLBOY9uKrB8XJj7d2ZU3pmk6FJQ2K2tW4FhC5o
OO2F0P3i/DJC8z1rFudD82r/Hxl0jXkC+Uxh9e8v1e9xW4px63KPudl6qto9rbUU
q6n+E+9idNVWkJXaB5p5LeO1bnXQIyOWyN5LmDjBnyuuLCLMQEnx8aerUt/FQzIh
asaq+DXreFhy3qC68U8CwBALHmq8b/upT2iTq8nRsaGJBFTf9rhPdilfb3sBf2E0
do4zlzTaUhzg+uO3TQBHD87KorOz//hgv8FJISPuhkwzUIrM6CuiJOVJecWB2zVg
Z8Ylv7t81rSlemBi4cG5A9tKSiThNW2tTkTDcgXaFXvpWk4Eurl+cjt22TK+sDjY
RUyfsrcyo6tevKMIwMuc8fyzbXJ7d056wvXmhnvvyuOqYf7St+C+yPKvpYox/yQw
gwWtq1IkEZ3q/4M+yQw43ihL5XOCfjvCSFmm/UepyySPJJSIBW0cUjokjYbt6XiC
UeyZATIgHQ890H0rnxtzQeBBM5PW08znrX697cIE2FtWwoTP+lk/Z3kTkthM0Ah0
zwd8tI5byQkw2yOgy4wziIDEuTUlTSPj1aexpOz33RHUqhYXLV+/OHytxQbIIucd
oWPNiytASQICb5MR71Ef+IQCR1LCP5cGgUyvkENjr3RyauRV5+swuBIDWrCAzcqV
91eKj4cOZP9+YLmGSUAHS/Qf9cV754T5jnr61C7NK1pvkovEHK6KJE1QW2kg6HVz
VbAVAjC6x9GRRRKiyo9n7a+D5rcRDi5pYHIZOMRPHDbhtpooOoSb7kbK8oENSkK4
+JLCl1VbUtRoul81upHhr/iG+3VEA27OOtwTv7QWnaaBfiJjMxNd0I/ndvKSnrUA
rLUwT6iaQOBeoEX+3hQCh41DPZcXbaz4zQYRff4ZqCR5DN6sLh3wfeBjf11mAlRl
CB8imLvjz3Gyvu7rUESvWAjAPATgvVwMovEa1k6DNbefiH7RPrVJbDoyNLQCujCE
xaLp5O5H0167F8RIj1lfhyrr/wlYfmCxWsLe/2n3IBMlhbwgbveYK+tLVCetU1WD
ZcvLB9z1zHSyY/Q/n67mFLytfxPDV3pZfKOC9CL0FZlkNxmoDbxvcbbj4S8kah6m
9ySjjlamkSQ/NuJGniD0b45OxfE2iSoLON7fQL//hw7IwkKGD6TMLi5oEJ8m4JbZ
vZxcC9QObeF4JsWaLHN6Me2LDJIVSYCwTQGeGRhc5IU8tcGVibZyew58D+s9NUIk
IXKtc0yK4/e3qLoZrxZZ2HxdABnYZRMx3rUsjT4iKvLNK8sGvf4cpS9KRdwmY2et
pO9+WRBUgLrZle4MZ6GRRDj7jx8buGDZx/oXooRyjeq3HOAkVXrR8zEkJZUTdpLZ
i14Nq9sWqPd9Zc1K3hhJVEIYFGfko2xuzUmKt7SsFLoFlmoDMkfMly2lZCLjN7Mn
jRM69NR63LJ/GX7b/k9KlJkFM4+TBKS6PdDGSlBK6xx/1fBqohgGZWV2mtG9NWd5
NoH7kLMx7G+O5MQrhvdEvSnTKpSAWOZhsnT4bwiVCqt1IgTUGL53ruubgfD38StU
NGJ750xGaXpMA7cvLLUYdfn5cau1NQqc0mnvsjGYejm+piMeV1ibSRwF4OUJsfC7
4Y++mLeux2ijyPiBuNpKDHs2VSmhYbH4n4kERKUT+LRG2NydnNkGlZSpotEa6hmX
Fwmm6zRBpPqbrHY+uiH5RhIouY5nZ9cWKvoaRGxIIwegFqaksznvaY0DCm5mtMmE
2lFA+ZlngXKNb3sgh/3yPIYbxSwGnhWeGkpxcCH4+gDWGMuVHEOOIcEBR4oTipsC
dZ7P/f93uTB2VahPPRHww3SlzePqHn6i2HPz7t30vZS/Doy7sDKQ4u7LfRaP/7iw
ZhLHsDK5lN3gI8/kyN9wX1/3pXYdg8v4ucT7Z8x5gq4ZEBQhKFYFmDvhgTs7JfBc
JudzDdL9aSkyjPnHVrh0qaql7daq2ItxtYXjM/tD/KodIWxjB8mCCplkcqHwiVmC
AeIqrbsRCLDollcyz2UdyUp+UAf/W21n59NPsGMUPCqDiuZ0CYTPKSeEw44lI2ot
+9qEyEyPNlroH7ndYYT2uvSNQQPY5MaF4n2+9/9NJS23XuFFWkcR+RxZQ72Hja7L
bQv6HXpUoMjDEC3p6TyzVW2ZLJ1FS05F+fdeT/lA2nn9EtoP2QI0/scjrjKT4AXf
Ia5K3dLXfGVHiooOOaRoo+i9Dsu/aM2RBDunV+VxTId0Q0h6Ps+dI27b3UTZH28P
s4gKyTr1/nhryhN5vPAkFUoAdR49NZjS/lz3Tjphx95UbE8NJkq2YLvNqcAgo4+C
BmBoeAZhveYPdvpiz3fw4B24kzFRWRsJuK6RLxA558kSc8vsBvL4dYpn0jXTeFkg
9VA4DFuzZAZ+nI4K6y7hXA6SGUazwNald+zx/TvH6z/7RTp4H9O4pmpQrUyxz3pe
Z7A/5b4LrJUmNhejo4L7baMysVU+frf20jLKnSIDtQ1Yi30JG20kiYL4xkUuMHEz
/THR7wgEqmpXSS0sMmcBPcEWxpK2GYfQLbBkM8tB2fkRdgIUrEQTxnGsrZ+t86sz
AI8FDA6m0jJQYQBwNRCQcoXS63Mlt9fpuTSBWUiabWPBiyS0esfrVVEaViXlBbPy
CjtfJSCJL6IwsRN5XxlH8gwQLR6El0EwsU2WdSgQisAyhfqAga0yftJTVqe/HPto
pBIzoPaUbKNpn3u7/ZaI6+aI7kRW7tXRsDtJ5oFaFJ8xAvz4v1YC1XvqE/7rFBl9
8PthrK/+cuSjVWR1PhZpKW8qCdGWqtTvKR151jD5j+p/m6pFAIRul8yzNBS8xpjU
RFRB61Kmkb/b1iydveqYNGbEz+sXPpO8Y4Yi7KTKtrem5x3Ycc6VM+I62tgpsVyt
7z2/10VUlMOEKOYk+keUXZAsYEZeKuYL3OU1+8Sv/mH61KSlrJl5OU/6nVDoMw33
ZS0Mab9qcFMAkdRAFcKTNZzG9ZthKO0IzI55A7LKTjKzofKF4Dx/4urifSUZrhB/
OdFfSR0kmh1EpV3KwZwh0EjLz2h54VWaOg3MJoH+7EScajNFzXMAYHg8GnYlmXwj
mLi/POAZlwLIET57RJgCrI3SwjMB5irx0+fo+pRKXaztuwQN554khGprLOLCwizi
6aLPdJxR9KG/u795SjTx1beHRW7tBvRiLzhrzCYxef8jF8OWOrQM3mZT1Ai9DbWT
VARlubvkGTR/YdUOzMG767fiuDINIFPlOBwN1pa7DjXmFfBTWOUsYk4zY+Dh+z3p
99XJuasxvx3jIhKrgnBubiLtF/ogPQwF4kPo2MqZ0lpn17Og2CfJhbF6gVAx5z8C
9FHPyHDkUnMm/rV9UN8VSdM98Mv9Gmzvr185J+qxr1imhwMjv1uLOXC1QAKjT2r0
ePC+Ec/hWTMzFVbUbbd+IaXBSb+idIbRP8anwySw2r3z+49FB+a7gjkhPK1QF7oF
sQa+bBYyZcDViCS0T4cFooyeWZyg5FvP+bKUwBTq5W1Zy0PxCGRbgvyRLBJIXBvD
pH2NaaU5uM8AZIiHuL5w7eP7dtbmon7KuukY/HZh1L3W9XOOti84L7GM+fQdelVP
YVK1tUHJ8ZmtG4+j2tLaeu0a71NtInvLba5YQkbJnSCSvyteW2LV0cPkh6BvBLmN
lCeFLvtrqPQpS8LIqM2suzFo/Tz8M7O+LkST73UOR7ceO9KK6Uc4RGeSHj6pzD3E
X5m4x1H2L7Tdw2qd+uKiWIFP7NAYTVwC/my9b8xESFyIKyQs69bOed1bTXrY8wIB
A6WhiVc7/BP3aP3yHBoDc1I2aqH3CaUzGS1IGZQBkTf/fIhsbZVhDFnzMOoixxPv
Fubc8h/boEr7ManGgl4IW1p92lAL9MN9w0DXLwDgLcHCzew2VyJFmE/iAMk3GpBK
bS/uR2bUrCIpc/peS4tS7vnQgUv7X1NL7a49ENhqvq5JVxf/cMgAZMV9RwxME1Pe
1rIxKNXObRmTegUG8yOu+Jr2HTE5hLG8PALXUNCboHH4vaDKDMElqduy0AIyFAQk
gY/Lj+how4PlIVrbe9o4bAP/HQSunx1poz+c4a4yYk7w3psxh3qZYeQZgj6Dc6SV
3Xi8MSGGkaEMWweZOj80OXCdqnm1Mu40rWECCDJ5zYcUl8YwPJBoFWRxt6WG+lJ2
TrHx7Q9AwROm8HulojSBhRmXaZ6SRfswiw0UgoZ8KPZSMDPYYTCaAEgP9M9yVfbX
eOhXII9oF5stY1YWUsb5oK5IbrX06sf+t4hSE74DgkJYkSYNrlJIwsgp+fW/h+f1
ytyWJFo/tXjcyeEpXtTfC+BCMjaSko1AfE6VrKfrSQ/w8WV4VlSw3HhSccJ1feDu
bwvqb2dowJFa2zhlKgGev/0E/2zj/zCYKik9K/zxAiJU1zJ7ydfWzfof15COeX2S
8kD3TFIG+7SAOpruscDoGRWLB5Ah9+b0fiqZRWgQJ1Mt98o3xeyWvI4NefngdcAp
vxdDE8pHeXELQljc6kWGNcA2LpSwLKsrjoJglnGz6j7pFfARiewlX1uVJzImNpSQ
xYi4rfG0HUaF0jsfwaKMk37Ggej655mB50n6yT/Q8JbpdkuPn6DaOLP813qA/was
tOp5uTpZ79icP/vsBBd99cMVTG0Ct3pEM52A8Y0kAPnscph4AH70jxVbd4SrHKyu
m0HVrF9tMiXIjEIggtRW4dip8yhiD91voacvZ0cGnJvLKAqFuRTrNhtzQolngMuQ
XqxPm/8JSddWVMBsaupWjRYIyxk8KASm/PB/FmM+WqIkvj/9s3FCuyPk7amI4RgQ
xdRDlRrN1TqMeHP/CBI7Lig3kcAfDJL7AO+4RUgCcKh5BYrvVSO7jG4HfSPaEsk/
OGmEzM0FIIMldIcvW9tluB/jGUr8sA7jiji4Pmn8EiAKOxgA4hVRfIkBA93X34SP
KzM/WYZBViwcpW9mZ5cU6MeA/suItJrM3F5YfFNCnM3RZfncdX55peAHFKoVwbpg
RSHhL3O5wd95Rb9i5Av/OiAZdNcXzmp2S61ytryLHY+KidTvyEVlyIypQcQQ+Yhm
sP1xkVP65AXnvxRabDh+h6BIY/rpwf+tfB0ekY1aQofIfsEa7Bn+xgOsn3WzHhO2
CRo3gQtrcM2chBoVDDTBdKijtTIO0JrTC5uwFdjJThEUhJQtcF4GQQK6SlQ9bCkZ
3LN5ApZxfGRkQlZGLTluE/VsXSLPTVJHXZb+yaD5J+gUI34A+f6Y5yrJzdoF1Rjr
x2sSEEFTZwhKSxf5nhVLUjomdkryE2v11wDKnP0mw/5PICVwgMwqbavZKo/3H/4r
NgE+N7J1wQyMwNNQk+uchoneXQNC2BWLp0Y+h3ACn4pG/eUFIrKMmF54IezZkxNd
QBOoovBV7xEusPnAMoU9p7W3DJSX/jo/Xnefnibw2dfH2FFfjpRomf+ZZ0dJpXpN
85ReGeA8QtT5uWsO+9ZwN7u2j51hW240WCA0tQxZqUd1jWMT0UcdVlddYdoQiZrw
Clm1rsSm0K34RLmrd99HURlLIV8HjdlJcbIO+KVEgvqQItze5dtsloh00PrlxK7B
/lJgbkNCpd43rLD/pwtAd0ET7bl6Xhtzrqd9VFYAHMicLQyzpRQE41aEH60SZG87
lKv80Rka5knkMCD4BFC2esKwbOF5nnIf6dNNDMf1SKjg1YNYAIbbEuhdrrjVpINb
NW5ZGCP1N5z01Is1G5dZFl5/lx7W84Tj4hhgXo8/zaVKpmR2ek/XVjEfRL24ww9i
i71CowDvwFY/we9FjMTD1DVyg+jMjkM2kipyMNs/0TrE9qD7nMW3MI6Hc1N7XhZ+
eQSGjMY9k3PwbGHzX6VciNBKIm/vrjDdrkSOcFq6AwXnHiFiCzuZ+T5XO5EN6vgh
brmlLS/RlxF4Hox4/8/NizzMOP9i/RrwoGL1BTKyY0AKXjYFs7N0bX0+/c4X2ARc
FasYdQzDEfIb3UAufWCfpuCapky5yzz2TBK9K1mvPNBVnTFSmB+wJ1aibG0fBCCN
1eSnw/hW4zdqkaHYaNdPMOz3YxS0MIiPBs1Ot/F94y9ZnvekvMjfedqVA1CEOnFH
IVsKkuyrCSP3rkVKHG/sToXHva6UnKBEy81nANxUPV74+75E7MxmKjNUC1pgCfE0
zlkCLP+0qBKQTQxi+780ZrDHoRIeu+xEe5I2X/PUJJ1Mg/wOTqJQ67wOqJKB25fh
0q/JvRSua8AVycw7nJwC9lbPQT/txhG0ajYcjXFaUBvpngfhwWmXYvNEjIIFwWqx
9natKrczU1V176OL2rZE3xTsJicfmbxpLZX0Q/Bmo+StHUioOgQ3yPpPqN4+VG6a
GHXXhNt/ze228lqT+vEJr/bGhxee2EMorjECLypOQqKKpTVLveWOt1IgY3lfIPOE
e/T5Dx1rjAHNAJORGIve83wgbJnBSvTj2yV494ijVi8m4r/Bs35eA/DmfJT26Vyx
StWR+cj1p8DZwkHaOV+ENuU+O2asUmu+ELIIgr2rOzaoEj/GWu9lUzPZhj3WEvU2
OpzXz9pe7vGMUPN7ggXXhk9ljapE+D397/0DmcgkrxMV6jEa2UJ2jzUKFGDvkN4k
Oj606mXGxOX6sI2XvCmWfuePVlmbnAK/NZ7rJl0hr33T3NYvij+nWIy0H3gBsq2d
t/hVyAsNjcWgSh7FsVAkuX/CpSVOauaPDzrsmzb6JkUinBj7yE0TXDU92upQTMel
TuLNve8yqY/ukL5/mm8Tc+QREfxbpQlX79g8A9a1W+/MH/72GkiNTWU6i6AEM2cW
X2l24/eHxvi5z8QfbThuLNJDMsx1d4ymPNW6ZhZ6gBt51HsgGakdrRq+6fgdpnWu
OT/b3fuvgTmXmGZLNdwufme2MrJeRGnz/0RgHz3GGi56ddcT7D05jAlHdrpsYSUo
5sGe70D5rrgsEkjGEpIxCZ0TeIX0AQ13EKY4HpHi0GYO2/8cD3nW3WVWb/j9FRvH
MJREHAyM+pRVyM/dNlTlDsPkOWdtbpcfPzHEFpK4Fuc7MAc3OcKqZ9ha8K3NRVOi
/30vz+qL/dk0wHQbFqYZf08mPNr9yJTWvaHjug5iLHVhuHG8/t+MgveuqIWwJfL6
O0eTIEcdzf8QN3iKnslTkJ6PNknmKVVLWJ3as6Jj7Yt3NbwIbpYpTRxx9dKyqf2W
9hvEX0DSsaCqWvtg1GpJ3uZcnXAUjIe5WHOYbZ1mRBozmW4WufX0RlRkDMnZJM0l
Sh8LKvJVs8jSri3osk3VdgvS9qdDFi3o//WxIRvtYvxEVD6CR7CAEloWLI8MMN6O
b4MEzYTcqHFjyFaS6EniVTDkMKncZjGyjEe9g66JdLja/pQyE1mbK0BX3f+d8jim
MebVm7sFKg/ZGOrpy0C63aWtPiSmutoHT29WYNMGgBhw3l7KOsF642gEkkHS8+Km
D0VBjhuMtD6pJZAONmQ/qklYRuGAkxcP6VoE4+rj3Is9WdJ5OSsP/lyL+u2eXy5w
FSVnytE5eFSkImJEtsriUvlE/qnhEfEdavTrrfcrzMO/wIEgmnSbAdjf8kJGLJ1F
Pg3KVnitL51XCB3f5p7BFjOkrtPwde/i4yB1VFhQ6WsS3WST6rRrWfPN5HA9j6M+
Ue/xoYHW57Yf4aTsvp5TZjHVAB8qBWriI37GYOUZ8UUFTq0cWQjMckuTDlYfgOCL
0fDaCYYHI4eWxM+25mXcsuhF8+Fj9A0c5D1A1tcLiYWbmxcNJe/MVeURrqIt/7tO
igSk9yax3eJjkjrWoOricaCU9agu0oVzl19hOS0lmijri0yGd7sur6cUuBwzScIa
eEOpU/hHAiYbR7FLsUAlIzHl2VmX4oMknkTXzFqTbSxrTBpohGcc4VpVkrCrPZJp
oc7wMmFeSH8VNAxptcAhKx8jwgp5zwnyNYIXwwCG+naxdxVJS5TfnhSDddHE/obS
zMBsGj677SrN0R8OkQOz8u4wAMbO/UNZzqqb8rVA7AFEyRhAa/SRwISyaIPGpfsG
zYYmUTuboLK8ZWu5xK9DkAs7w963mzVRQVWoW0fjAa8IqcY3nBU9bABAbyV+pt5F
gqp1Vw+/NWwLhiBRyYG38ZRNokJ7JVpuUUKq9FBjR6k3hTXOSG+YGUoelQjVDuX2
gPGkt99kmVr4rfPg6zeeSen0KTvUy/ocQ13xs/xS+lzSbE0w8RrCv7MQIC6hZRea
odn3BY10bbJhLRHuHcR7wNTLW0p+5HEnDhVBEXbV6IqhrsHSe9yFXwd5A2uySUdk
u15d+jDj4lOWTgrIC7rZ6bQelo28pPk1HWETBa8qKdgw92+7KuCKMRB0INqCm+uY
tjzne7fHRh8x8hG1gofcbpetJDThUxCzEBMM+G6wogKDAKR2lm8pbGa+EyFdQaz2
A3E3F/+CQa70+drQD1qLuuK5CRUsvQL8nwFmH2/vmD/0HKJl1S6Eb5529wf8T6e5
WhN3bUL4M+c8h6HMTfxs3SbVLmIx7DhkOOa6z6EGRV/YQaBRgeYWZmrMzlQpiKzg
HefaPdGNZtt3z7KZhmP/FzzKtxUJvTzZJWSBuNwOrBZmRUjiSGGYSUR6L/h1cgui
wMKsVdJwSV40Br/THj5mG/N7mr+t6TJKGXmm9VUSUgki7BNVl1yvLW08SktTW3fI
YGQ8YWOVHd53+Xz1CdlaJ+rZabn0wxWqaZJiAMbIdVeElr8SNTsLjHEtWuLUPepi
3pKcZ0Jk9xT9OrqR1AjqG3F1vQwwrVszVETKbLEXACLFMjiiMoP2ynSYpm1ayc1z
MwB1cDq3iAGlu6nGD++x5WUjiKfQT9E+P25ZExhRnUBfq0EAWCKAKdGeCp1uu+T9
YVMhmDAY7GWz8yAw8ukB0PczoqPYlchIEvtaJGH28sQeA0LiPBhF859ON6dH6FvC
5pfk4QlHGWnAjFvZwTsEEFa3mDPHegcWNSHldYADv5qGOK6PPsbKymdlyUL8tJxz
NwwEZHzBdGWk82SXGxmds28M4CkbJYYbhV2lZh+u5OgcrbC4SZFy++WYvzqL5WL9
bGmFUdFtfNJJG/DQwK8hfdgPCM7GCYX7Ah9l4eTxbNUnaRM4qySswwu2LWWUZhnq
retoEiil8Nto08RZUETSFS1ynmqiXfJUZnttp1mSF7SSEtemTGYizZF6piyy7749
6FsX7g+ux9Y3h2zkgAA83jLAi61QFXvy9Mf5V4qE4cur3hTjcjN93dHpRZvWrfbO
fmwUmjfCA6QQbpgBAvTXCnsJRI8QMs2olO+YGd6r2Tut80KKqa8jObbnWMfkQ305
GLRFzv+x4wolaY6MyCCUk+IrAHvg0alr9E05Ce0o4y5W7lcold8+jgFRhsOAahdZ
JNif0BvCJ3k0/S+xkoRYjRU4W6ZhTxa0l8TmbMxUbRWYME2M0aPbDgbhW1Le9Mrh
nDdj4dBoAcDXmon4CP6uJcf0Qd7ubg8sO57Zvypv07tEM72AYr7zowYF4+X+QtDw
ipAWDdylUmTBYvpGzEI87YqpzMxu16yCvbJvxDs9sMEiJdYrVjXojzkHN9EeEGr8
Y5JAzywffqriROzrx9tfWw8xSKt15BORqcsT+tPOgdAQkdSZJWBni8ZAmJke9JWU
SgcWPEK+TsXVaFi/v0QRp+R30LjjuRx6RubrS1SfdOrgul2hJmhQ3Ij9qJ+VeP5k
j8gZrfOneGYhEEZcs0syM1UPKA2hJ9HgrXbuhVGF7501Z8+4Zs8bqlVWbfJe2hZ6
HGCv4NxbBwyU12eys384m33Ogv7IFB6sC4uMHlf+edM9fMpvFrM4+J8mASLvRt2U
8OW+RZErWpXpGKMH8TvfsPOoECJBCmaVdG4TZYmRerDRT80BONYsPIzPidoQEAFX
a2I5JozxOfN81ByF3wzoYePIFs7Hs1U5qeohK9wORJb9tkrUxZL0NFbzPhmCZFr5
1XfguHkigYQFWjimJStmbddaRnYg2scZ/J3kZHbsq4DXTOig/GRLk3AKQgGRsGrs
8ybsk90LWNmGBf8I5HrBGoZgJSgzZDWrvpjET0PleTkzdEiHe3k+1lLlbE38kUy7
HGTnl3M7TgjcrCIPJT61PkL45cddGF7fzAwX+N4zBWTo1kQx8QCJFy/kzL4erFtE
YDYGmRM9T9IES+dI6EaeYZizPCNg93H627mHPa4CjQ5V7xJoCVGsVX/SWYSIJHc6
SNmH9epQfrrjKAahdePd/kTWLaNLzljIueY+bKTdOX74XuExNO0B1JHchFIfEsUg
9Fn4xhUp5X1MCIJ+J7gH3DBdqG39bhhiXugP3MPNxKzwFUkjKqvl+bj0sVxWbhVh
UjO2rvjvSV9+97nwst9AzP64ibaHnoujzAHFsN0yueLe6VKi4lCVrXCGVJqTwqav
W6fXAA1EGPd9P+Y0cf8sUfolFNb2uZGEZz2f+xsE2eEywJOlK/AReIhs7Reti2Lc
FMrwdi3qyk3kTOwYF43lPVqGgzY/8golEHQyQMMXAED5RWA7gyoEbP/frZO+bjSq
KLCD8mOYbqcd7RlzYir+bZE8PzBLM6y9Egqp+aUYkXviVNp+81fpkZYoGMP0zBUD
hC8PfvM806BrQoGGSzzJzXH4/NKXarpMy3ljMSQMbQTZe14ewKcIeg2UwxaaNe0v
jRgyPZAUPEp9/h25Mve7ZKvvY4qO9f/wfCfGiZx8tyXk50zmFuZMHlhdKB0uhAlR
JEeDiGDo0pw4SOeZdosIZdUKote1Nho+p8+35AjBVuWGcojuqgL6P/IeRekr72Yy
kJyNn6gRs54+KmenGaJSAOXDmPNWju5PJXkKZsYUQh/tKbLUwvjh+DySJJ25svvN
53Gg70BKiTZ/NAFUI1XH6DsSPtkMiT1QmYuFzysrdMETAaulCpcnyL+j7UnLi6XK
kCClA+FR+eBBLhcpYl4kiEelXpc5aZpY+E7dxFX2TOm2mvE5FVdG+XQd947D+6Zs
kOXqig6B/ETLixSmAYNgTEFe3DE51qp7jVda4VY9qWSkgztfMy7JEtj8j0ARZwwm
PlkuLxqKF0odoo97xodM2cSu9zzOa3FIIubKNsvtC3htbpX399VqvE9w7MeuLjAV
gtivSO10gu30/XAkFdG3qKcfsyLjYzcpLFeoht+jldl9pvyn3eqHHU+HjL7butey
8zIMcnpqno8RfLD3YHe5lOtt1asE4tdMSwSCqBK0QZsTHY/MqHiYUgCRcCsfmAmA
wwoLrgwRvcG1NSTzVI88tQyJz3rwoozZglBRJagrE74wVNAkejXM64KcFia228pL
vT9Aw88FLaNBQFoP0couXsbI+Q9r/oSy1Ts4RT4562aiK1RUJ6kJjcviPavN+Vwb
WoUjA390hSRl7EcOdkwqiCoCUSSIILTmD5odg+U6iSdPhkt8GX0L3jCqeRtcUGZ6
u8Iew36pjumV9OBz6KDsONdqHqvD+jBatKhSsIXn/83tnmiANM+i17z+4wFBdB8W
g5OHknUZO/KXe7p2I0jtAyZg0aejOZYHeXVu4w+2E4g8aNIiQry08o0T4CcevrTw
Rq1ngZRnzz6Eq9Xn80oLC9fYrbleuM+T5uIn5njnX4M7uKZ9ytmNWLBPtADQ0QzN
a3cIplqx3tuW3zsrnu160HWAuzKmOWXWytf7VP7U9KfKqPHKeFJ5tHtoAV1iNSgC
CGR4Hn5c3+yduMommHp4ZSF3BCINIhyh9u2KyF7YFcHSPOggd07V27r37rabcaev
DR5MPxI7mBXdpYnjU0Bb/x0TOjLs3t/kFt/qlUUgnWTSr+b5TcbzfJmA5rTwK7/F
wU+Jf+OaeBqn5fbLhWoEH5JMWQLxeXodUjjPZWPFj6HXFbV2OSlSbZmKu/KZFv4s
wsNNaQq2u7e9I0tvAFTsR3icotRSBZGsDjb++o5At9UuySGlcMFdrD+Ew3u73v4a
M4mdZr4H9jJbmjiBHH+Gsr+N9KyAvvC76jTEdYfNOGLdHoGMDy5WlSH7IvX9IBit
iyp6zHki6w00La1mnAqN2dl5iGAet6ejwpJdPMjGf8aBETGqZ93Q4mta0+A0uDC0
EkyWIcdcV/R2povLHsHPLLtXjGR9rm57C7zYFiZ9UFxM9sZRBEJ2MFUW9jkSloKS
F014rMzSdv0xuyWbByLZBiBb0CFSxgOZrRitN64jimaM7BFN0bykxpYskcF2zp26
5Ov4R+v0HYvWzR/LrM/pdLv3dld0eCbiaVMmO5i/Rd5mP7CBVANAl6XzFybQc5Qz
wF4VlwgpuEsIVuJwPzSAzpYmWLbBNyYKRDgRtHbB/E7TI6DjdKMYKdKWklvCeMQT
J7/B6XkqIXLuAAXSGTvIZdQRYH5pUKu7OCSo3JdCXTF8cgBAWst/0FRxTGbS/gch
CkTObJZn8sdv2V/RI19ATWYeoNeB8WP6/TpY/g5LvIDpMysFbqQuVspSsdBHXA+h
IUcabxfeyf+sVb20csq6C9eewDV/pnhChlGDmDng1yv4TVAZH3ZTedhj39HIw0kl
Bvuhqpr1Zjq7AwG1Uwxvq8sGB8ovnTKNeo0cGY90o+fLhpC+7t4AjoTKJB1CnQxc
j3NQgP5B8Y3azpsVev8kP5jk/l2yhxwsQcDEg35HAzZuC+ws+127yihWBS157EFO
+zR9FR3fgATv/CokmlRUTRtwHPnpGoVkHTlhFlVZ3ZEv+svdAwiXYw2KakAs/Fq+
B980rMjix/I/SKEqUyqYVPaJuS3bgf6cRUOnvwTgnfGH9xfwtAg7b7E0RBZNIwTK
NWrl/8+sCaXR6IwFO20+p34GWjghV8DgGS4gZMZGMS8syDIEnTdWNvT1qVwjvq2Q
NJtsNCK3XNPNFFKzzxwPI+390qr+4dgyq5QwQJV7pzrucJHLxtBclIUrbcp3wU0S
7cDkjxAHyQ5iq5Fvc1rbcXtTCWu2MiOdIlyrPwHKhmUK+t5h5mJnsCpGiL4R450A
j0lpfv2H2u+wOi5WTJfcA+WPavFzk7CELTGCe5GXakGwvvn7g6NBL8uwGZly7EF0
S+oiLzLotuVBpKw7qg8A3vk1a94LE+KPw69UmgohRDZ8RO3Gn7mDbAEicnoJncJK
wPPHOS2mxWf8qjE/J7uDRP8v4b7b3n5Jwa8Wim3Ht7BaEdaghNPHeAg8vF8fD6xP
yy5Uc0FQi2pqA1nawc0pmy70Q5nC5pcSSpifTrIvq2yw/75jfphALxKpcQPaRlOq
fRSxt6fcSJnRnBbBFIHv0F5u/z4pXOv+uG6xj51tc+hbd8wgjTQaSVWFp/9cqIzn
qfkohp6rPxuZ+mWoCs06XIVp+i2X1A9uTobR90AQbuhubsQHTcys4BSPZ59r5deU
SO32QOeSD6r9sX7CKPFRM3nZKxmaudSbBkWHMXoCsAIizuJ7U11+ISzosMCsyjUN
fNDyg1gAJol+SOtxvmwehqDzyzYguH/kJ1bIVQOAb8V5HeryoMFI25vbPACwazEr
u61L05/fsOp6MQ4R+wUOs69zP7D+BJ74VBtoQ3X0JLrp22mCfWeqg2beLqLiIfRp
e99UjraFbZ5MaItKR0sZqpwUPZ1bhOmixcQ6b2lR0185Kh7GiTx1OhdbkUQFQVat
reYZFmARfL1Myk1WbnieW1rr0N8ys++L6REKsVegFzgGNXHpxtvupxVdtlwF+yHM
Yp53P0FlzKGZaMLD93XtEQBjdmq00TkSnBLvCeZHdmN6K0FBRpxlJcQc7CeEBC3+
W/y8vW5+uTkj+7RjCV6rRlv2UoxEILYb6E2yurHM2EMdYOxSpu5t1VuNcj/ftJKy
Ttlo3ix8LRUL4wkMfwcvcYoEBKxwwfFMWuBuA8MAb0XscTxg34gsHdCSbXIFh7sL
nSJn3eFd49BTVzll2tf6RfbtMmzs9MgMnpibdkDnokheGv6b00djNXl+jKbvZiDJ
FITR0tGvJ4hl3WR0GSRNogCzEljtFJZ6TlSLKPe20FZy1TJoEUvAAw7F8dMYa4ls
rHoQCMgXyJVBmpdmgIA6nlm80LaEYHmq/z7XtFSWYEE7wq6H6oMs+6ydET9UKvsO
1Qis3iTsRYsUir+65eLszzDYJuNRDPuobgRzODklUTUuqdr+lpVM1J5S/baFiLKw
Jw3/i7/CuGcW1aEJaFV6EGkCY07rcZjYTT0j7Av7JuwZxonfKkHk6OWXSPRsdYuU
9nxeNiLHjbn9gp7NSpKKl2t8vIaLUiJBrsyksg0FQVQ1wG/poK+XUhlCOtLEMbc/
oJkA2DJTAOQ1etPD8KbuATbI13CLzryl5peEG9F34a7JNyRLqV74G/BvcxGHC2RH
YPnZ1zaRINQ9VYpB3E36SQ3J9vGPwdeGA/Sjdtgx1mw2452JZEt8G7F4fHr9wihm
i4ncKLDZtyPD6Vt51UiK9pRqEo6plG5V7YC8vqDe0OFPZ+6NqLnHpxKYJIh7telv
JQKJlJqTc22tvdR5/tB99HVSGkNR7rc1jDfizWwF306H+UvnKz23QXL/zgp6JTqj
e7VWn6RcIA2Rz/WDcJltC3LttwQ+KFcsFhPsWCjvv+M/cvCADG/HPVpQXLCYtZoO
xvwMftl31H9D1DXX0PvTyrv+pxahhd+pxPOL4nQinTlcO/JhHybzoaSvsl1eGh3p
Zmk72/eVsOV5hlmnZukUrtazczHejIDxdYgEezI5mJNiHyXs8OoVOs2SmuBzt/jX
g7BZTbjPTiZXL7jdC7mAV9l1YVEJsoi/P7wMbSDxuVTohs+ajfHJrEk7jvqE4Utx
KZnsQHaK1KyLFKQvto+HPI9/dvdE1i28lknpDqnNnYrWJmsetjx2t8fVK8efyZAS
MOTvvnDPSM8X78hrihXGhnWMBJwh1yReI+tmlxtpwqjdzk31Ur13iEksBH5bATeA
4DcxKX5AbwMPiDg9CXCXx2mYJYGQyKU9EP0kcgH1NLkL9hkRMGGF5zmDuep6idWr
FwzJXGoQ2gOGdOasWBpvhrI1GVxKoR6WmYgpNQdDEK0uwgVINGqUe3YcB5x6XcDs
cvRLmsZhYKxWmX6CeVgzK6vzuRDLo6G7nnmN/4IztrsqKl+emIZUcHopCgrnAat9
dcDYQon8dw6lkfJQhCLviNNYRx2fF+Hf+t5SI25PERb3dvQ06vEgfddGu8qf122Y
ObvxK89mIYMTBE8a0JZelvqni3PIxB+1wVDd1I07ebFjN/Z6Z51Bi4hx1QL2mPYi
ASweEEfdZ8w9w7Mrk8d7h15scZm6J6ulKt2rUoPrabOdWVXhV06OGsgrqkcZ6yit
W0H2FbFfiSvGjL3SF+Ew5y4Mq21t8HmOrtCqJBj/LMUQ2CEzeZh61swPx4FdGjuA
R/4NJE3pIc6CZMYWf1o/rLYctC+Hhv8jAZnbj5Aa9lnvAdnHbBIdz+0wHIyX8m+v
vF6mgobMFPiioQbL0KWfAlpLBjbJtXThKoJVbTKDCqH3wNS6BWsncT5s4zVG3axi
uW630a4J2+1JQDCEEo99pMimO2MrKG5RS9lI0K1vdlFVYXVvFf73Q3rTIpcomvp9
DrQfW6NbrhLj7zbZTFxHIgZ7QbEwpA3FBnLh03QqyXb1DnatmNNJ6CXfzKs8M7Bp
NAndtrMzCrKQi0Rm1AEDfh7YE24p9hup5wdz4DiTBH5GRvPWpAm/yaQAtNwWbtn/
rCuiCnSlM+G/CGAA2mAUZp99yIDLKnF1nuFPQKvMTjLv21oQS1Fx8H6wNrzgJ6gm
dRoMOzxfxT/D1q/lzhpHqAd4SPjHNajH1eoiafapyrhQvtNIqxy9YXWTJmR8YXDB
uftDQ6Iy3vKU+esbSE5+Oy169irzbNCXS7pFFiUUZvN+6Mgu8QsgmZ1O4GGyVfPx
p9j7PU1H1c/4CN3IlazBdypdx9KNW5rPu0a5ASLo8GcUhs6mVTVsxIQSnsf3Wm7W
YL7a2Fnyf6PGJNszM/6lh4v6XOnAivMUOOAlENOV0axTCzgPuJRdbzKctm0jnibe
9RcA4iOJBdc1XtnClMxwvE8AZgKxJJrUmFMyKiYTfS9IbsseH/m2zQ9mhKTr0yAH
N/zV5VZ+jKnXflcLqEcea3X1QEidDLLrgWlLAmjMQJvKpp+8GDvOfYocLSqjTBjB
Wz7AGvetD+c9OMK3yYhoYspquiQR6NFhOUIapERAOSes0dErouqlkYZ4dpYTUxQn
98RLCcnkJG1utqWr1yTxzNKQFc2XBoqbJF/erdnl+yl/mS7xg8VLnIxJ4TZklE4N
BdGpgW6WlV4Lr2tzxSs3Y4dH0vkqeLqGd9RRtbdTJiUKMGRvinJ4lid2gkB5djUm
p9erB63nO2FD32NfROh6lmPucdeCZo35D6zFA41yFO4hKvd5LM8i3VfDSDRm2ukT
/ErGmTD+WbHqfz3W7ENIFdvyY4VTS4ys2XlYk/HtR8UZpdsIx85JEY0XMRXoFJZj
bG1DXcVH/yFkjXgIQkot5fRwby829BeWmcu/6PvKjq0Qc6TLw2yEkcKq4AAHtxSN
CGS9rd7KBiLOTL5h+emJNPRBeSwSwk/nQ6URmmKrN0ld611RH2Qj1BxSkkN28+s8
RXobMuVrRF+W/DIB62FSoeF9Oa9/pWH4wkrqF7LdPjYVtK2oTsRkE3+izUvXrtHP
VVf39FkYckuPdGh+OkdCdZq2gkucq6aROguE2iedT5CSoVcFwICm5tYxdN/VYmCV
Pg7J13wn4cOsuBf34YF5k990y9FjAg+06SL7YG8RLadIiEZIrFlNP1R/V56pvMZP
6HPILggjUonwSA+ei1xAs44/cse2v6mbQfq4mBhlHOOic4efuNDsxFCCdYx78lb1
6uMXatq4FA1Qj8kNJK19hubs5zOtT6VK2dkEJc5nBPs0yagXsP7SILNqMJUgzqPF
PDdQrS9r1pGi6G54aFMOQQV9qxZbVzsi3CVfuurJgMrrjkpYOwbSpkWx4xZYStZg
FxZvSdp5DEW4FMhn7wnKbeDNHFznbMoCE31tcyZNv/0C6nkDqoOmYc32//iqVi7K
kcTLK4Vvta7ifbG9cOhr8I9SpsHsef6CNASibhdBbYAofpksbgcllnEtnRGv9FfM
6sEJOd5WVBY1wphLERCGaELrkRRs2NciA9YrArdMjqi/MkItMAuJ4Pz7LIzFYppO
6Tj7ijkmjjY3ofB0Kzl/hk5tnckHUXxIWVttZ+xxgZWJ9GvwmiGqOE+byDKgC3pZ
tbM/FfzIffLtXsjGDF+ILUNHV6mNY6HTErXcXPbcodYplWlpCBNCna88H4HBSdWy
HZuc7uVXvAnKWkYTvHYwjpPg3rHpTTm1M61b/QaLbQDeDq9sp7r13jEM1tO0cp/1
czF+BS2v1YTHmE7haybzXIxWFWsbAx2Dfspe3eL7iOT0nTB8pUOXyxGB9ZYfSMgA
XIJiz5tx0YIvzQ9G/ka+/AFTDPv1PDXnGz/SKcfNJeZF6w+E1OLU0P3HrQbWGy+B
HrC2uRmYwIqfD+B6bZczWYJp1FcgEL2ymX+BxJ/zTAG00k3yB2QoYynT591gYjLM
DDN8eqIubTnwZro/DsN0hhHEZGYvYPqKBVyxZWtFAiX/CLucYBkw941aie76eXdk
CX8Xh+6314tgsKn2HnH0S1/SHbcv1snEYMo+hf2gI4LAZOJO3DWEUMTxrc9vAna8
+45ZRf4e6+KMf6MzIzoV/1sfSvuwYj/ZidQGIlrnSw9YLvdCTlMvN6yh3t0iG0xz
Mbd2yoPEclvk2dZtfegB7jKsImvAdKUB8ouLobic+lAv0AwAJ5q4t6+bbBPitCWx
LIAXOoX67zBIGbGrlLchBlQvdHEkWeDGMuQo0NuAwVY89HaAREEyY76pRIbdQURz
fkzm6YcOGlp6CBX1UZAr1HMt8ngQUfmLhlBvxCYTwRLnMgVBYLzw+KoQAxGd1+6b
CD1/AkAmHOM+p/5N2Bhztj2K3jrjn+aCvawnpcvXkeH9C5XPM/6eKQbm2qnVYRUZ
23/oGVryNFytrUH2cr5NE43KdAheWaHHo3NlxpktjUIANr38QBiQ+5FOL7rDUK8P
aU/j3JjNCYbhMH0AESoUSHKo9Z1XdpikK0d0ngQuWlFlbJD2vjZaeO/0NFQOTqHX
FqAX8LhqL6Pvu9yd5Om3/Olv4LBHawBaPaLHAd4GozVKuE/F0SYbVJ+o/RNwXjch
iAUGye2K5CkV21AVCZltpt1iiEsoV1BD1XKjPE5OXYiiy8Jk5zJQFwDcGZD23ibm
Dfi9sFWTwBrndzqGfROZzyFca1FvJbggyUk6pxPRIRRKjAR7+tdG5fa71ZGlrQlV
7g2LFK5KZRRCmyS3K86gnIla/G3XDNC0izU8fsTHSI8oxOSE4JEbwX/JhVa3dSbG
xPYQmttSuSEHtDLlM+tV9z4u0ecB+7PlooHY6lyt6hrVSf+2pozBIQrg1dLHu09X
Aut5Z6nJ/AJmlpX9H98jPFTO2n4ZIPn2Eu4PbwuzG5aBGbyU8EJZGEFsnHHy3LlV
Wn+GIencqOyiFLjUaGZGjZ3REMna5lB9EbFDN46cTrvzS1Nk74YlM3+FYBGg2dba
4RTLpdeOMN36udqlUaQLMfayegg3maHtHb4/yKl7M2u9z1dlTaVV7f1u2qnVuWgd
kYMX5Zj9Ps47J/rYCPOh/8MOaHxHYpTzclgcdPfJVsCKJNwKPQZZV1j7M3IqoyDD
azWQb5DCGFu5ojEMI9AjPs4NDctplYlziVvOm9JatMYvU8yuB0AMz6q8z47Zj2mn
r0I7EXscnEM+kt7qlH+id8VAROcs+pcvgVxyefAWOjtKUFZBti3o4gT4qU9KJ5Ec
eUtNUA5sriLUhGS3WjpRPJLm31fJDprPyeFpJyaGmp+tpSRB8tEtQx97AwXUIF60
aHSLRa71tZoduTr4xIPPGh4HD/WaH54MxocRZxkxHdj/l5DinokuD/OPro6fNNWT
h6EmM3Q7N2gMHWZY7mcjGg/UgA7Q4QEMjuPFoz0kNEmDtxZT972Y0Hh/3uvGDRhX
sqVGVJUwtMAwTw1X3+eaQ6Q/wYFQ4etRyOsAqL7YtcUAg16YOz30NNFDwSzXsoxq
pTnrfI/4LVq1ETI8T0xCS9ZNwiWJsSJ9vquVfj/s4AAR3qtut6KzmfaWc4ekvQra
oY921gN3lRgxGwZIOYJdbfAiYykL6SKTFhtyy2BD0FcYzoTTl9pYslPiIbdTnuoY
zL8Lnf+KSZzEuDr49gZ8tLBOmAKpL7c+rzAmXSsG5cHUfuCcmnX3/m1GTM7li7I3
RrslpOfVF0k54LRlRPH9vZh6xpeA0oK6Xh8Lc/VYKnnWmyqlmh3gmVsHuUGqWpbg
MiRN1Wn7cnoJfsWLgwNusUQHQy2SSmUvbUuSu6k6rPRS4mvunYOzAmL32RFf19/3
KSHpYqxLl8KOTaaD3yymUhS13LdfaL7uHfCzq4FsF/jNzztvUvwTPAFUZIkdg8Rd
G31LfU0vmmsjlQnL0wOzGnJgLWFDa/BoRWpFFYhAg6rNGMYkzax2PDV4L+4EfMTa
Vrbvvmr6UfGvg6JsGaBQRz4wvQTJ7SeBOwNygKTBFGn6NLuSht6o3Wgv0JXpEk9A
D8a2k6uDdcK+8ljwtWIOgSytrZ4MoMdJIIZuKDEF45v/bfYVK5Fot9FXxC6g51XY
EzCex5FHaYrgg42YWMkNJrpIb+E7ekdK6wnYNNVGI8PxOHF2GB5jjTWwJ0OF0fO0
VOWGasdE2ri655IL5tLfbO7jElqL0afVw7cbesoDH4TUtdDec6z/CQEHnPdQCc9n
XmdwPfvlpq145uMIA+eDfP3qwOF3EP+PbVuAohI9dW/OjbvR0K8PRqZAsbxu2udM
u0wXNRiqpDQR36f/GVJXD4iN11vvvy4X2aViabzhlVQkNaP/tLzwxm1KtDB8k3De
CjKm+I4ZkxIs/lZt6nqZ1+A8zUz/dASAlQdY4MoW1njLsI7sg6uwGB8EunZBZ36X
HegBwZwjb7CALrxU/CyLhOkLsFE0FEVvJdJrnLUffRqba+Lk4AFkQydcsacfCTl9
jWmzO8XMvWHOg0tR/X0ppWSxBgbe5xROREdo3mtKUheE5UrpobGLS/6na2pPYyVU
4efWyIOI/nCVI3c/HF2/CIY2E1usSyYR4B9v3vbF0445oYojAuSKfAx1gG1CCLqP
EypPmAszVVJVJJEEDyKm5PKF3Ba0iS839IOsgNadon8u5Ef6s/JmMBgua/mvFpyV
E/WpGHOediqV99TUTvFVOyRgoWgf4Q7q+MWihVl3HPnfKYrgWQFOSlpcbj24sZ5A
CmI4J9iQtbAQg5agk8AcsHN6J3SEzYUL4nZ72kaFCCqYwMsWNn2KXUSEkx7VyTmK
8ajhp5rKcoe7K7JflJ0JyUzhJ+fZyJgLeWOmSi2LtRnUYnTFzV/cCX9QZol6xQa9
6peb1zpyb18CBoiykwcjkWPhJr5TjDFte+oJEcgThNatNPR4GUC3gF9WcnMg4lxz
NpUmJzvve66CMnm5uNIRtcJjCju/F+TpHxuQzIdoFIklzMZMNO/N4QHhxgceaJD1
6hl91YkTmXHNpaDCInE11DdRWhEyNYVxoY3l+ymvsCj3hRU3qA4yQfgvdSf6aUci
IDARGWJX6akSI3OpK7zI07YfFbcRem1vzUObYUcm5JIN6tFduesTLZtLeKSTxIOV
vdgiHbQyy0FBiUHol7TJoicnxrqSIAqomnOssxgo/tfw0t2O6uMjXizCr9Pw1zVX
m74o6r3YprNn95D8DwsBV/59uAdv8n5fODOe54R6ZozsLPGA4zLisDwu5owcsc6f
KfCc6yQMu/Hm9aCe8ToX0Kn0+3LNCMvZVrc00qOdPLpoV5ubPiS7iP3zU1U/xk6L
JTseWlLJTkEovzqIT6+dNWPlD6RcIkT6kFxG1pLg6QSiikwVEh9w3pHDYDzC/Un4
Cm1BcPXUrFZecp4R2hoy0+bMgx7RkfA72pCgj2+p6QZYiR2XFDTKNbdXXgsUs30L
xroCVwv96aeTJr9HAJ6lhmPidffejS6fVzhsTj17+5g/duPh07kxSmtIC22/73yb
PVwDffhry2WW1UEugyeP3NvlqEgQXgAgcQ28JpKt+YV+cpOBQhaYjWOSPOUI6wYX
hLta3TZ8eD091ZsszeUyEojBbOzx5CBbakJ2xPC9QRsPbBNon4WZ1VqlOlgNbKFW
kM4Gj+zIloWrBaI9W64U8d6M51SPJLAL89hw6whUVOsrxUi/We2NoB5xFjw/oLkr
riovStPk0aaD0fVvsvY/DyQCJL7i7JS42APTrGxOcv4sYCYK3bUaaipZXyEfJYC8
71SuH3VaU+jNjXJexzW8rxeUDVeN7Xq6hAHXV3lPLgfC/6FLxqGz8DstN+GHiG05
Bt4ZYmuC5bYJ82W9odgOcH48ZeA5iO5uwWijZPAXAvloTQQqg/nahrFHvqHf9LAF
vkfypSmA0TXXj2i4CRiVH3L8botNfTDxhxeZW/UKj7KrWznzg28AdOwu0pn1SUTd
MtYaiwfCt0kgDTmH3cULmX9C8btBCNEHKNb0zOqs+iPu7nCAJ6StghTO0Z5MzXDT
BYmGVMgDvKkOyMLflQ9XgdR3+LbF0vnOKgeyTAWT4wcO6MNBkKthdrxEofIcZTj2
iZLzZ6uiDc3BvJ+uDbkXJmLSmVgRihxIIBWPQ2eqbAZ4w2A/IeLrNzt0/B2fZhzv
EXeGnVYO2E+OF5oyXQo+Nz3mY/hqibxSxFe0Eu/FbVbdrNYhwwB7aK9DphC154E3
5J2KgwZsPpjxGdN6DsVQZTYRS+lLkDzRl4hiCvWXLkCV93Fe1lIdx0vWIoCupr6q
SSWO0v/KaUrY81L95Wg5Pwlaqimq0+ciN6cnrz9O/Kskik/YifW6UHvurvBMmSVG
/zfq1WVH4EsC81uYbgHpe9wPrWGqGvHKgky0P9bE4BrXuyFS6NZCl87aeggMaZNq
cGGkHBs3InHS0jWHNhj2XWf+yrX0gGdqLUgKABHJ3O1DwggydE63zraewuEQzDej
LHshyQ57XlecTKysE+MKMpK3JNTDoSoMat7csdF+hdoDc+W0Tt9LgCZEVvs5zJhz
QtxK7TPaNKjvkeSdIoVwX28lIXXUMvv7K7Tav7oNGdSakqPUudBgd4wWm5mYGhYP
PSrzTtDXOREfFHuoNceO4mnS3e/dCqDyjSfIFL67rdW2qMpU33s2XnXytLya6iGT
j7L7ATml8jC7T2DDv3O4hyWoJF8uN6pi19/DRCQGCiqlFqORiLVmlrtpiGGSjNgC
vFlna2/e5j8NbAawW05eZ7aoSsD/AbxTQXHoYGEq8vCAXPJYf7N7aWIu1/WpKLq4
hhJts2EnC/8cyk3o+V4bjdlKUKzS6MHE+qxaFlY/6qAGV5yHwYzzTzs7642FXGFr
uQoshduMgsUv+VDQCDdRWiOlAOiaetGIpzc+X6Pzal9A7T9C2INmSJFGVnfR+gJI
S/1Xc+SqIqP0rWo4kx2HbpGejL969IRUiogSMW9SVkmXroz5nNSnVVnUHggCgSCx
1IGj+EngKhTbPOpkIcYHeVNWTsC/hPQfWhMRepCzlskNz/ZzVTANDaLmVgprlMoN
/UQrq/kqgSETvurqlxYAXFwQWhcPItU/578lvBqQKMAHCwBIpvkBwWI2JXMcONM7
aYDYWd6Q+aBeYFqZVrjCxfqnWi6nqF7hssCus8tcAUH7i8MI5cki7CAc7Mo8P+RK
S8P7MUp2K76vhA+PjiYIRULnLMyFYE/ifVepek4eKVAG4PcypqI9LoqPXRO/oV3d
3BnvxLR/BsApLDSsZliAa9QhOqpvSRBSWIRbPrheX3YjjmmTPeq+1X4yWAnNKhyY
m/lUSPnaxO0OEQYv8GXoapJrWNKgA31oeSmRUzmjsO9F+Q+zqhMODcfuBRY5FIRY
32q1ZNxx1/PxK1Whs598CGVvWbNvNGRFCQCWx+sZy/H8E7YvwIlH3ANC2kqe92ch
SgGxlVQJA7otaP1P5PyQsB21x8/amPDWVOlAyoSLU3E0ZIg+eJNaz0BpHTD6RGE7
Q3396x4Gc441W4e5NWPSVvx7a3sYFk0LIiUwXHO3Zu7aWOs8iZyrpoAkwuxHTB9C
o+IQdMsGINUx396b2TKv2st2LYg2v0CBwap6PzEAA46S5nVP33cO6vqX/f4TEXnV
a6j3TT/AVaMq253cULlldg0WSAvTCtXBpKfm1/tVt8AJFmukrNrerFO2vY9r0wet
GyRdmPklwsFG1HYvPMkKYqGn71DlM3K3cneVXTUlpAD4bp2sgP6B2WNwo0qWydOi
2XUl0T+gfSXRO4eeihfe8gn3fCfPfe2ErzQ5RxwZ81a94JeRjNjxmtTA26XVegFd
UTzEFNVEUhFP7+DzPwgy4JnWCteB/1Psg+xh5yMspRsUZzbqWrwlqESwO8D3yNhr
mxuR8ehkUjwM8fexQlU5ZGfsBJjaieBBqZ2vnYq7oO0W/OcHRpiOmr4Ep5LLkLzX
EmVe57iQW1M11O3E8HDh8a/GNBhZJMSrsIBCk6Q7Pk7w3YddJzSqMWRWh7SOPHwf
zvSzZU/igz565fvmOKFy2z3YY6Cqqu7XKA044akXG1FEwnUPWMS4zAneAHKE94Ay
Eaz9LH802wn4oFjrPoYPxFqK/NBsokhdso8he44Y0gbMBpRqMs6/XtVY30zywIOS
bPiGZgcCdp4kJJw3YdQ/qDdyVbm/Zgq+F7i1v4w/BWr/k43bmf9okT2WOC6FdAnp
0qcs9TXo/AGL7I2V9UVFh5xX7VWd63/vMLwlovC5JZNCft2/DQ9mep1SYcYrFOMq
fS0mATNT37ucfy+dluUjvE0K4Kw760e3qK1kRij0Zx2iz5d0x8gOgwIgIhaHfQZG
qtt+bP6nhTBAZIdyVOKtnHU7wjfGWyrIw/ih4o2dEmuBqwuqkEhHHTAxxYcePQ+4
gongRD4htYtyG0qBcwf7q1gsdgTCAzxylmwTsoLFe4b0k3wBm+CqU9Xa9sYTCmK+
/VR+w2valvmc/8EdH3gUIy0lAHZ3pKbjRm0IDLuwOMK1h2/VSfvixIEUmgbnWd7r
fFDQc9Y60DNaVUnndyEMl2iLO8cl3C1AFIKBe5kJoLxF1fR/x9rxAj2+xaLqOW6n
/VGS6bNMDhG9UR9hESpZL7l7nAFPRBkR+EhvHZvC816ka/jK9F1zKxH49OnwbE36
4nvYT/64WtJEm/WS1VkRutVHcBquMXZOc5Y9vECvdBhMnNnaBREvyqG8VfiUz2da
DtX/KuQwK3EUGv2UBDllCwSjnLGucQBYQuW6nkrcdRQKzxsRM9BMCyCZ0gqHvRNq
rw7vn0EXrEj6FMHmcFfAWWOect59pJB8Gpaxq5hVlerzs5083JSwDVvcXYw3H6m3
C5u/Qju4bc8vTEbPWmJAldyYbK5LwWeL3K6iuy0OyXt3AgbcIgitydKrui/RePzU
dA7LGVUHDrrOoUY3enNvAXShuwAdx6l1X3s2tKp/30JCF7JGfwLjE01LLVnMexMN
UV6/F0Kp2DiHlrOMhUlXqr6gJzuAErtcPUl8KGXyeIK0zr3OV/mRxb7v1Jji1ip3
/bTZmWWPORWQOQqjeuFCzDhdW33Z2X1huqSdzTmxs4dqYIZSvPwwJFcKxn7c0CHQ
cuu3ORIgGXq9xBIYcObSx7R2DRGHh9S5g0VIcqvpr0ViojoE4J+9NE1yg1JKq4vl
yX0zUS0tNdreMsI/9X/0HFxQ2jOrtFovYqkHYi3RmwyoOG9ypoRUTD98oQTTFK0y
HN1QcgItwzWSMcB0OI+QxgXqnyUXJTNrqcQCAwt/75vJ3N/sEm4WUpDBPhA3vf2c
mXVbDBfVH9hDvuasQv3IdVHM3U4sylxmPANL4clmI2uVxoQ2QgFs7hmaserNtnGk
wYIx7G7sOwB6MAEbRS6mU28Mq/M1iwH/b15RcCmmMxO2WYzL8bIpr/AkQAe6Yq2Q
7zwMqoEB2SRsFFZMUOs4RtQBSwPOGb73t+pmLPlQ1K1AA/DIQw+uusy5nfLvjVND
vWaDxE65/M2NCecJdWetEjFAXdvL08Pizqsm2kiheNWwNHXTECA2BZbZ7PdXrxJ2
l7uLdYus6vgJXe1OFIJzQ1Fqzteb65NuH4fpC+HQYsAsSPzZ5EvyV0rrpjc+TRHw
YQrXlQJ+MyaGBi8U/Mf7Sy9MZ7kyVPne/tzXERAe/w/CpDM2VgjQAAsnDBbXsvyu
4ghBXmZX22tA9Iku2cLHZ9ukcMWiBFJWZjCxaJAwSoKraSUk2DOwM7mZimad3e4t
bCxVZZBLbHoxVch3e1UIi5Okt7CHB6v8hMtTs7l1AAbdkze1Ysr+wGrmeN5TGjDF
WXtetzBQKfm1xl9sv0NX5WHLiOMXba9Fj3HBor7E2EghAoyVJBEnftRI4XpYRPY8
7VCnEkYd1NNgDMwzYhwIpFrmcimnW8D3mOhucDQA4durnJzlb5QfNznvCgHNubrK
zrttj22549N2m+kCjtkB4n6zG8JnpI1mn5EjHfonxXY1KeLtMsHrIXFKgqfB5HEM
0s7GozGpxZk1tIcRa4UgYegxm59F/8rGzpQHLkMzvVreqCQoRd08VfqftL79298i
KveQbUmn7ksPdoPP1V8l12h3AZGn/s1xpyZnk4RoW5rUs3LflQEPM2VLJ8Zqw+yS
zEVul6WxVQ4r3fFbA4L9ycnWD2ajCZ/s1kfZjHiYuW9IFg+EPhLotpxMYlg1HRr0
feCdJhkrtK53cs7s9pp4xhD/ApiYapMmM4bcwAGGCO2+Ef3IxxVlzhGpCIzmKgqO
nnr5FD5Sv1EZxT6xwF/JjY/FXyMDb/8+zaxBnfM/rmcK8RAXFOZ2FNuITm/lPWr9
x8Dm8aIivQYdQykG1sE7FZN/fJG5SlA4hZo4JOqyWkFuXV9ve0czYOwuDYkoJ8Hn
/lMvNOEyZ9kHA0Gq04RQvqXARCYVRfPRore+sGJEtaSxoQwbNGOBYbqHinFNK75m
MFD3zA6rjQ9GjycAIIW/KX4nG159k2QUZ0OlulSIViTgpKsnTk4r5J/Nzd5hBPLb
ahhB608SUk2OYt+9hS6e7xiqv3R6LpUGKVdhoeRWFqifsW70Vd8w51k8ddSfO9/H
tpNNf8mj1lim5/1JlhfBCWdlLc3LuQ2NVeVllQ5WSN6i8J5a/3CPzRXHtuQbRozF
HOgoQWlYKnHV+tJWMFDSvukyoKAGs9LJbIthfb/2l7X6vXwy0RyfzYneYZBY0Bzv
tqtT1BI1rUDxLffS9b/ksEg09DHMMGUP/HCNpvDw6GbfRARr14/LmE9yBcEu9USW
sk13nld/YlYvUHnM9VirQTXd9jMHYyCbWZ0aQCgxz3iwXwyPemQEdqmjBdzPV8io
1ZbzfIrqS/wPl8wkZxnBHx0sOzu/SRdkOrWDajnQv1e7PwHXm+aOqzo1+NDYzioo
X2XFLbEOpaU/sAe+vF+QG+PIRjO3OTUBIcBOXJjX3SYQ1q4U8N3PDscSgi3TK7fb
02LZna4HtHMw1UVc5qFM/6awrNxtjuTVCMnrrzzJpIMFEcUQsTD+hRCqoNN9hRw6
SHZ2sPH82YLopcnF0Hf0Jnp32mXJRhXn9898YcEeAxPhShr7GNGcjCkg4VFI2ckG
2qj84omxFaMQtRqbnXjriv7szY4FPjnKk9XBtkxk/2RNk+hrm1TNle8NvnCS4uHd
Sc9LCpcxYs/fgV4zgNgYZHs2Mj+AD/OeXWp1ssa9dA/7v0WXrB0IWDMpxcQiaK9x
n6AQkRfxqL+NMkJAL/R3MrDQ/RiFA9ofpel5FTFL6G+7LkmxVqlprZGyLbfowy29
uMjXLV74pcREB0/y7Rxr1IMWD5eTL/K/o2WDUTNJC+beXnSug5mdpVGEf6EbScFe
QHYC53IWiklfkBpGEZceFlNd06zB78QgdV3kxj9Axt4uFsRw1WNiZyomuMKxODh7
ZJol36AvTRYID+52l8GVvDd3FVKuNImF+pM66DyYK6XxxIzpFClHOb9Xm6EUIYQd
28Sv1rvZLsG4uNftkAsrONCKdGonMJ4fYhaLYR7ZKDa1IftRhzggwljCvXTXpaxY
tYbFiovNaGJhBTdhizYFCoqACeMxSiyfvhlFSP250cuasTETHuCyPP/NsfUSJnze
bAMLHLr3T+FxF9aOrXocMa5OhKzr2X5jv76DkqICQCYj9x5qrD29E1dAhHoFWJGN
HEWWmvismy29is55QeWof/GYnqFXjx38D+4XqSin92Pk/ekMgZC+fe75CjHRdE+r
0uV6viK9hAP2G2eQCxebl6eP06QcNOGo9REpJ6y8Ojjm2kilSKMEauMV6Gx6aZJC
libopWvrV2FuUSYYhW+AP93TVGmpfiuE2rs4FMB0G45bUqX0CAhnyJfFoDpb5khn
CcSJyeruTlI9PIWIcbgF0yB9GNTRi5hyjrXSPAOuOBHS4CQj0ZkqvRPjZL4fsfHd
Q/pf40oBFmCg4SNvWRYBin6swpBoMhs5fM7m7GmO19bnnAdFqIN9zC1z7tve+3Eg
91+QMuw7ELPaHRRKOBwOaxPnB1Jb4ZgjvJankP8c9SpB2plOlMpLkN6ziV5UlpKC
CxX1wjuzCMGE6osUOFpTu8gngaKVvzaxz5vQ2zBV6USZRRdqY77j0FxmmaPoJ360
9qAExL8Oo95jfMtPZiwAPMpLW1Oweam0sTfZ7/5+6oYKblYgoKNwwf42IjVlaVl6
7tgGf6LGTZKtD2Xam/8oZkuDZ3ONh47O4GJQkUPIxB7h2pfw/0DHBHaKma6p3Hzt
f/Z6jbTrr5DJmpBgd3D+zHDYNuzoszKugLAYNMpzsNUjlXCu8pnR+1uwotl+/XCA
Ff1ZQQQWEjyJGbyTEwlY6ffCBKqCPQJh26eslrzb3/9lC39Kyh/9QOqF+2MchtP+
SwXJ98kou9IVxTdh5n+AnnSwFKd6t8XvY4VPR0OHR3zz36Bfv05DhBi+gPedq2mq
4IA0UhYg2tpV2yFcEIB7mGvwp1Nbu/qNwTnI1zfluHTZN1sezWqXqMabtnQ4YW4K
SxhoqIIlIXr1T8bBiafHxonuxFxncIR8djM0K4lUB/QlbDWytPmnHyqFPXbPgbXn
yAApsKO5RwVTKcX480jyQryZtmWQd5lhrHzA8lfP46AI3J2ErTD1abISnY03niNR
FoHd89rd7j/VGTy1Att7wSZZJXZrvPcVOJLpr6jJnbDhC4fp4xoy0HWQJ37Dqz/S
VTTHN7JDTLjHP/TahiX2iJhJx5U05uNJzHt6E9XyDoTKlyv7Pku3tgrka2k0DVUb
lfAP/TE395XXQ3SUHwaU5YHTv9CjceoiOielzNb6ohfuCwZ2mmjk5FqQOAIR+IhN
nG3c6glfwlxcHn0dEMs+8wHrxu4asOr6J9wriN5+kVu9Xn5JSlEHKYyE0RF7/Xcp
bkxbQVp51jPNoxpgoQsVRRqwqlh69qR6tqiqASPjQDDfdUZnW4nwwo4sEGV58Wb7
KhrFzYb1QVsMj5LYDFzgMTgQL5eNGDz62jCoEoc75Vwz8EWT4PlJB6+j0dz5SUH4
g13nMNCzBxBJJRQfrgWQiaDcon9lSVWRpvdYHyxBoAyw3WwOicY//uzTOM+d6Rzc
ZM210mP/Jso64ppQLbK3NfEM+CQatGjmWUFKnIjVGAKt2JwvzP/lbBSPP4LRYNb3
VtpKkigwfQ4Mngd5Z572230uLPRZVvTxdMIET7/Y/ZXTl+FSVXCUII7xwrvjCEu+
NA9d9U5zyJihMiFQl/DXumHrApHn+m6nZm5dAWBmGmCMDQhBj5laa1ofuPvS9V5v
f0JtfRYHod2ukaL3sllTvGMeDShxnZKBl0AQEI6UcMJKBAwft4c0mFt6URPlaSW0
T/YYFsEQMqaeA5pWnkMOUoOu2a2rKRzv+oFO/P0xwDhrT6iD7STH9BiOAs52nbR6
CMTaNNuC9gtCdqcXz5pKZzCm87L3aUpXgkXnsVIZnozZ8zKDBG4iedKnvOa5YEt+
JaskoCfWE60FRtq/XwxMERTl1qh8SwDIPrGsM2dUuchJRifAcV2ljjpEjK0FcLAE
4iwPu/bUV+f0nl4O53tCdXzvQJCFT0BHxM5YPTIcyjYhfx8lsMTEejbssvRVnOHE
lmo1lIwYxiHaDmAsKa1y6Vu44xt0GwxfQUSnkNhiZH0QYxsGbWSDfZmm69W7LxGK
tJQMnuccCQvT6NNW8tuIW2mz7DztZpfyWUqRKioG13ujReOt9RnAS+P7GzXPDPgG
P61cHT8qpiYp3iHO45msDToVedGAmvxKxmaXuiE0LA/+WSBDZ439TInWxM5yGVLI
2yFOQYzVy5CCjDCGtqnHRpGJVHvSWEWFQIdq9Cb0pppkIwnCSUZ/gushaYBSIfmL
rhWE/NFe/yhE+rJFolKtTxTML3SitFqUikyqHND3eMbOlO6bmIT8G03sq2VHt0HL
li9LfXADyGzI1TLyFnBNREte4OfNl2sL3WQQLdKOHsARNmC/3Rvgkm3G9+x93sB0
DV75drgXe85usBDarnCA3wryuTQxwHhnkobINHEhkcs6ZpSOwpeUsn5KHayWFRb9
+FnHVJPoyHjicBps9i/MHbaje7W5/Hjzvd7mUYLjjJmXWMHb9hdrfRTbXJ95/7hK
0m1qltpz1Vn8jgWh5u5ciPlqScEABlE65nys4TxhxtL5/zNIoIUoGRkWMwVc7Khi
jqo9fcxUh0Q9XopFKr75eka72dLHe5mlZvHKrKzOaVml0yJ+QQ+rqhSYW3EZzbBe
rr5VBcqsg8RJUA+dmbBkp2W7W0tGbJmfv+gpWuOUYRAwURrMsjhunDMaJVg/2ELu
LBb/lCPU8l76FXXr++ZOJPpLRqCiJhr772iwBPD/XtwuGKSk/hSm1G505XgmpD6z
6Xkf4BeVEpa2zKypqh50TGaVOYHtrH9tv+j5a9tXra9P4ArHwD8C7wE/U8oLMwXe
wwSfAlABcQhLQlH9qvGrOZUyOzTQMbsRs719PsjXl38/OraK3jvoKU1Ac1asa9RS
r9xNiiFLnde0lMlFQy+aNlAd9r7BfH1d5UaUv4wgIC2ISnNp8YOM/kFo3pb5i6J1
DEnCk/hqeOa6bFm9aVkim+/EXzniWHhspdmnKueuEUtit/yOC64AeudIsIeXokzU
IyPhaaIA6IVnK38wrE7WJiMWmo16NzR1PQOsx8ogyekqwN+mJVHwIcx94lkt0uGI
cgzNWCcbuGWquf+OAGPafd2a+3NmUTGxnWkJZYSdOQHMmvPufrvQ0OkutX9mBlIh
59uICPETmXhIB0t/7pyEYn6CaKu/6YrL3zCzbAOa6pkrCOGbPZzvpPvMJibpH2vl
O9cuhIynbaeh5H+XQuoL9Dx2ER9qHRQ7YcBM+L9koC44kwBtY2lN0nYSdX/4tsq7
h8kbpwEeL6aYqbss4DlOjTsuDvJ5jI+e4BsdfW9TO4PXhHHpGycz8kjUz9ZHxSSB
edr8BO7xamON0f594IFBKPuaBnSbLfch5fZ5LcTUhjRbHSD4bhBCpPycLRcmEpnY
PQT6j6l4WiFeaexYNr9XhdZ2DSM7lz/P8WuOjjRdbMebgPiD30D6EJuu7HDaXWjC
j8u5QDIRswkf1QuOXsxWH/BnnfEoxLHQcWoxYVH1vG+ySPDBwc1XVe0YcXc2nBVc
sbme+knTfoOhyN7NGEmcUCxP25xtSBoW6drPAWUvA+UWq3ARxkHuJYoTeHaamted
dMHwx4OpbqpbTfMMJXc4AUbPi+q3CXvbtNPnYs1M+XE+uNKiarXnRgYYspFv0LYz
CHr2Q/qBy+7oz85XXxIoAcQ27SJI5M+XKHZUdsgAp0cCdsYhX58DLmV2TF+J6cwi
BhP4elxQGxggHbutsszubhgH4i7AV96FN1bNQ5h4hMAgu0y5KXiBOE1Yj49lSHAP
1301cVvhlSakLww6FpMPPLiz6iBaHjB/2yKLXkYZ87ZZi5VrqJwwzz8pNPY7+aoV
VBE7oJoS488GiHvIEAqchLKNTXDhd6dqpxveB+rfKAAgUXty3meF3tf1KtlZng7f
FBnWVCYMECFaV6avoIyEjzFgqi5PCBemeHMGKqBWXfHZvNLCzCjTOB1mRvdyDXEk
QrFwrMVbhyeVJixKHGtPcqaskgHv4PbfCuCGIu2pFMt7v8D9r+MFnUcF/1+PM+Nm
bKGzvneAuMkjcvdwBwkVAgasYGwHh72K2W3RICOsWJXnYO38ripA2Nnz3V9kcVFA
0jvaKPPgWGfHgztReroNfxbqJIKzpW/0XYdr9bI9NuJ/e0TitKViGJkFQrysnrkF
hwaYukiu2gyKLCm/Rykzy4wyGHQPZ4jmWNjAGX3p5ns9Dzm+LaQyvRLf4wnggesd
8oxNM4vZqRZQiReGUICzF0hFILo3eGHYV+Q9l4wpfrEdF8fja9PBWQ7x8Po4vUVq
NFUiCBG2wIFI4h2zVid/MZILMqs/jH4EXW2LHrMF3RNst4vfk8RQjDzGgEudOa5q
9TrRRmED6YRXYD+Nld9W1zT5v212JpB9gWuHAInivRJCGtIoZZaykiIfxTFF3eTg
kTlyG37FihxSHYtua9R6NZLHkmr7wf+vnwIx3KfUlswEZzy5miD6ZOhHB3ZUNnZy
TnM14KMi5pIr9t9fc3tI81HulQSEQM0lEexZN76Xh0tvf8yI1V3Ijmw1wvc4L0nt
jJz9PvMrAvlxVygDLqklBlBcIzmhY+fFf+zJFQtxAUGJpB2nu/QgKny+ztEycUJH
bm4OPpcE4o1miK+mJ9uNc/N9pAY02s0RjGZNGvOeVlQC/63VybnGvlYduT5DI2Uw
VSVh5flcKH+YI7CwGZBS2xr5PSEifimsHMWnsrgX+jTQOMUXssA0rxqcbaf+nBwp
iyenWesaQ+ig5tkEUzMktKdCXcyK7a9Hw8JioXx1Sk/qI1dxoTFwxJ0L+ppOztk2
V+7KURK8kdqFzVeedc5IloKiqfhNAzjPNzx+WfVJdsTZ4d/X4H77d/MykV8Rny1V
tavEU2nAd8ghlsHt3GOa9NWAdtj3tJSYdJIf+UXsq60nhl5DAqjOK3e/o2p16vRn
A67aCWBumCnUdKIhvEBCv8VTo00mDsniH+JOCTP5X77FbWqKow9Tlc5hj5u8M8Dg
ymBn2GAT93ryZHO35XnW/nP7iH28sHoXRXjMYIiHnb/04ZlLTyyLOMil6hg7pWZT
62H2vLA3E1CmHAjykxAi1DzzrNuly5Wz943LmwGapdOis2iGha4kI0dHhP5A6zZz
HMU6xTkDoAHBREB23WJtUSqL+jZuD/leJEtyjm8v5qvjWxV/IVWYLHxSp5m1dr0+
WuRCaY5XaV5hRoSwRltr6T2rFkzaE1ayItpqqusmiVBMf4ha2hyYVn+9n1dj+e6F
HHhQNht+JZ6lC++bjBAEtD2rCg6RIN6XZNlDeVwP3s750TNys3xpifBK36PsZh40
qN+zbv6JmKolGw9ZrpYBWYc/y8uTZhkaLN8j19ZPqaCuO31H/BDlpR/ZRi6r2EhS
SEOwfyMALDRV4ZmQMOWirn6C8qMw00T/NuKaE0S78zpql0HEgcKuCcCiNdwgkR8+
8ZR8NaOsHhFnzlJmxIJ8VO1d+w8QRHZtFZvZNDVXYKZH9tlL/99ACbN4HT6tCVTj
oeKAsBvf9yEv5sZo4OYPxjKm2nsunGUWM/bsMMdeewkbf8aEqQ/Jjd+ZMa+fitM0
p2o4LgeRa9EdiKp6yWNTd8QyJnintr5eRUhZf4nF4PgrYGuT+lU2FsWky/+I3NnP
De1sS9vEMarre9lPruKwRnrqZj94ZAMnsf539SkvJO4v1TqrqXN+Y8F32YN5366i
gkt7fOJdpmGY05SCRYqll67158KQPeSrojCq3y5KsEpvnj/VCmuz0QZjtUyv68Ck
L9vJTyn1AAfvV/VK+MmuaQ8mt/0wYOFG3upkf37VrFI1+jnJ24nWa1fXJjcvFEkT
+zD2rsuEm1tODuK219n+rZ6d/JX6/vpD+NDODdr7fzklLc6ty9gz64NbDTeEyJVZ
czdroMJjXExfy4bzHSHEhdLBK8IMyZTap2nfq3bjnXX6uCS3ccjENUFKIlkpaV8+
vnNIU2CS3j4B8hejyXb7n6VGHCrct1nISP6+NCYRk1EyXHg8CUhIs56h/zLQhKF9
wYPEguRIoB2642iCZ9zaQNsyLiSbdwByklFhhWvGf/CR3COkVM+dgZwcSFsrqacR
rwjaZtzLxufLSaM+foOWuKndO85J3a+fxtQH4RNw/e4D1q0dAgEhgnPwcsRn89Tz
BPGQ4UvCg/LLEeXPmXr8WvhdKjOq8XsWxZdEmGyYO4riYhUWRP1BzDaX639ucTYf
xLfLYlb9W2TrE6OYuOG0OiTEhXSt8MRNAS4TkVAd1h62x+lCCSmSawopmixadh8x
7wOctF4LXzO4VBtecSGASonYQ+O7GANIJjegmyBcgq8RtDZSnWdJIdU/d/KHxIfy
mcUm7W0PX/uw1Zoqps+t/vHko7BRGqalFzu7oDS+h5h+3HRI3R/kSNH1SIOzUFjC
EnwqquLOOj4eX9cNcqzT717atQe2M37TrPjPTD6DJSMXDsKnpifMJI4HDd4WoJd4
jlSEVof4WCcuoEevO2FaHYCVF6tubIqjAp4xkKlQRLPJPDRSjM6jaq1cJXdGA5iC
dJ31Nf3t/jUw0Z4Qu+02lbn4q7lFC/GrnMs3GbcghFazzqm7RJZAIF0QJsddaSNj
QT9IMXSkgAbeDQKkZQdlRg0Ea+t3cN6dC9bJhZ9qAy9hvvXwuu01xUTkvbZvWO8n
8I9/aTksrdPwB5MNgzyX4P2WpW7R5GmtLZ/VYBMSoT1cnkKQnJkg5MusJcUImJqu
0KIC40+McDtvW82ClypUoL77s7I73LCSXBadteus/zcqowviPgeF+CBD7B1TH2Ho
XthU3v1e0M6wDtotrVDcAa0KOVrzqRFaKiOlcq6UAbnFUWu4MWgAdiLtDlSiB2d5
zG8HKkn2euHBBXWP+1NMmD5uswGpoyLDHJELKPtUVR3pK4Asr8/cBGaMRo8tBzFd
V1doe0sYBmBLE5Nj3mbt4kOmwVIjUISYp/051Tt59smhQaX+ljNt86fNhcmrNi5s
+fCENULNCgF8mC9EQjVvyGwia6KMIA6AiMAfg2uDP7JuMzNBc+EelI0JBl2veKTr
G1Q4JAJD+fNrKVMCF+Zc2yaXv6WV9pxFZu2nBVlzQdeqEepFctns3VPqDall3Yqd
6TKvHz46M7E+h4V+RVAgflnpQJmzDZH7/LVDOQQ8PnQS4l8jLBTjsBpUs4+UteDk
5ATQEAL3tkZUI3PA7lEH+taGeYx9iNCl9nqD9iHLaNJnaghqlOaAufwK72Pw5c80
+hJNOznEgpny+VEulpVPuHbAQrRojX9b50IyT6/zY0Wziy0CgKygZ8Z/hyGDhuck
djXbrTmiJiE5Ut12AZOz0FsH8gLr00H7SUvQhkSG4zQDxFD3ER3P52avZppUUOPf
+eqg/tFEeGFfO8CtUGaiq0nCkhWciFrUaLjMsX/rbtspFdYaBmIItc+NXOgr76XD
0WHef6FqXSWCaGgduwUMtF79InRSs0vSbQLqjndRqxYztsjXtSQNUtHX2zTBak/P
fEAkFq4tz6EWIpoakUY35pA/3XxuaiYuFapsB3EE81+ay5gOSfOu/2H7y2Gg3lCU
239FAlqxPakK5xLCjzLuO+RTl1pKbVP6YYbDE/urndGMd26ccl2qga3CvJy5108N
PvbG3lZrcHGdvTrWOa1fPDxcwaU7jUdNDTBRuIBxUbAQw7mFwDJFVv2dMbuMcUWg
cJjM1f3mX16ug/NgzTbvvdq84cL6poB8eQqEl+OGScED9trfBU021BYKLJTVm6Qh
z4txfiH87dPa3ZPpgmiRy+1tA+rPInbuKarN65Fqf4SB9duBlWoBKgZjuH7wEWuK
4E1P7g1A4TaIgCJcH4NUYAvyG38b55nsEREJDJuaAlfpuAgDjmnD+YVnBcs5WbsY
0G8dhEqFbMCh2J4IfVpJZd5JfEhXGj+TEH3qshNi4pIaonT7e8DGRTX+uYwlvdBa
1MNnBwZcgxlyDBWcffF5K3Qi+vUQ7gqhypw0nUteJ0yNjYZpE8dHzi4h3a4UMarF
sdmKyn55odNWWH3qRnjp6GlZsrrPHzStkg73mZPYfg29kOkzJwDID6/XlC9y4mKb
OhfDShvv0CH5EEKkZfbvjTpDFp48zoSkvlfJnoOkm/wv5Rq66NBKLhF1lhDSdoMp
Hk5CwciXBWfHp23W5nYPMBWeRa0VsTiGRqfnOBz06OdP3tyLfQjIJCVSiRXP+ztd
P9NSCdf3fN1IKdHCISBMeugKX046HqeMsRi8YJTZiHJqclPKEW7bjhjLyGNu50GD
gRCblJrnAySmLRxtC5Qyas6Hk8+alDzsqfSULVL+SjD/OAjf4BsiFsfyMGAJQoHq
FMGw9WI8eo8oA+xeDBN/ocw6pm68adVOA40Q80u8e9akvhN1PBko/oCE1UEZL3mI
59683rucavHDxQmb7H6pG1pnpF49xHs4hWuApnNRAEx7BoS6f+axJQk2NizoaBzU
vKQKY1oCM/MatEwAXW4jBW1o2so80+GjTq+FAcqIm7rytPI+na1qzjxS/Xvza2Ud
Qwq9Dyd2FoGFLmkHCQcnlnOJHdh3JQNGF5VKukoN6VnvRIrWrTeJM2qdfseOKA6f
QsnFYnjCLc2bOnvl0MmOMvwNOXZPnEqWth3VPWUC1z/gf5mJAkTgRUK8IrmCfyxg
ueDH7y6Xsh3gmKvrltEXYBNufAymIT6kTCz7V4IWufYfmpwSPDKCaiNOvuxGl4Mj
kVogxq6zcFBTKXqieHhpPB+MlSFYNfA2txDVufGVehPmjKb4Com3M+mzSHH9dM40
W5sfE3W4orfUqpshHTZWd1ZSAVrtL1O3U9Ailazm12Xc7DL8EbuWGj6flXQZStWf
9mFPKfS55lCc3I32sHX2YPcqkiHcTdGkCpkoVqaNI1XlGOx6AwY0jzDp7xMrzMQz
g1vY+a8SAILYJGpkNoBH4Xlu1C97tU/2k5BlXUFQ1CQSM/QoKvNiY/wyi5WGKMJn
PRuPbmGtLS6NZ8BJdvGjKJS9H6jIzDmFLaCSxt+JGqfvmM2MBVp87QcJmYa5vN0m
hIL1I8R9j/yvOwXXwU+erIQqfkEPVeCnS+ZWrj+9UxMdCavLK5YXfkiFdHeTRzuZ
uLxzlsF49NeUApfBC8qvzEV0U8JFOklw9A8HLVEzhhV9Mk0kw3nEmmJPMoxQgP7y
ti27oLkn5lXF5EqW4JfXhoDN9A190M+GF10MLm444jChy6mDbdjyuMPSFXP4rsws
80p00Vd4PVBf2Ys4aA6XGr+Ge9YJqDNGc79rAhx03b9TN7cxUpkrkqaHM8OA4/+8
1uvddq9Hn0vAVV6wAfH/HamJCOpcUeNwdDO6OXQNCZ7qNl2AM1aXvcMZSlu1HrQU
9gt7dArp1yv0ezPIH/KtBqRFnWY5AuRuMzQ4gQ3ZV8aB6rNJQaq1NMa0so9H6wgk
bZ+5Fhm2hrUgrdReLUpIgpgYLmufBxyg9Gdwks+R4DVACcLnjxznP1DHtV0Bn1Gw
8ZfbJHQZuNGKH2v1DiLxMLYzp8wydX/7DBYTeIwFYH4BdUi+C6WUPZSQgk6sjBID
dnIIKYB9s9ePdtn+0FFJCOfSC/KmKjzpMLluZwOsixgHaTq99hxUabFGsHwY8q4U
Lk2Z+J282kogod+UNgANYVHS4uJs5ZcnwDB0ir0bcHVZqBjz0G87UBYy4NwaSFDb
/91BWIaPUaGGSTFM0qglVZjpaHlcLjzkM2EnbRJS+ZrvSLJIdB5vrDJnpmscaftQ
uBqFJ1eNODF/5W8Fas4LFhSpxTU4z6muYCYS/yuV8Rs/0K8VC++84RPCUqRQDkDl
jiw+fn2BlCLyh4l/C2NT8ERRMxbQRgmrHn4AKYNswUDVQg8t6fVOZgju5Uh+1tMr
sJ8a4pUCjYbFo3BUF0Nr69jBPX0+HbjyOtIjEKIsZoIX1wjw7f5rpQziGvncqRzi
G/YpklbY08tO2yA6+LnK1zDkRTgCoDR6BB1lahggbvRYenAZnlPvl1nmxQTqwEAJ
SXQo5OihM9ZVM14jCwaHf+oMOlhKPuMOQCwjXCZtuGhkvL/qLnzTaNd8G40qGA2e
vwPm3EPAGscXiefzVarMbAQgRlwzNrqTWMxVTXv/Nt3hCEitP38VxT6eU+5JT3bx
xRlVDbKemCd9pcaZ+ziN36lhCZOnfjT1i4xY3OD9mSLisaPxaOinGfeby4n5ZboI
1k+A/NQRDpShTlGQ9I1cfX1eK9oDtRx4gObxGdg0C4XEs87U7GPZ0F/SIm6t88Ji
SO+veOsojVF3Q20EZ+ZBC+yVyPrnpqfCPNvtlbJ5xopzOBIUWdcPJULtyqJVTf+w
bRTKDogNeWjOFcpBEc7FhJKbUPJH2cFLyknzbkqVBk83xWr1uw77aswVhMy+v2Rn
+gsBsLuM0UI/g87x/b+X3q6IDRiFAfelicgzDrTuLq+s36p0ScOoSbVrzIurEnOK
WFO1MXJLJ6XUozEUTytACFxcHCSsxL+MhbV1DzF9qRE5pxt+zDeh1qhOawcD0wI2
3TMbNxOozr5P3cXLZW1pE6A1GfiIdBmLso3d2rxNkSOR/aLSXiHlNcyXR3XkyMs9
Iu43xTiITj7oPrJuiUMCTtIHUMJFAsBnlVa42OIAqWHL43tj+0ACE+T+uBM7BETr
gLtXZTpA2q3hejxFueVaIqqnp19kxqEzDcMNfTAuS3H6Bs2QDlHA2j027ao4YlLY
ifXddOzgvxoHeXPm9G98h4gxof1PlJ9veUQsdyEONSiPqZposZzZ/We6yC9DN1ka
QELY6IV+Cr9/NRdcuwVWW88iNDfaJtE9bPbi+k66Df6FTcivTK0ZSnKmns3e5adp
FpxEYQR59cDlQJwqQji2tWM5SXf7X+LHFG90zwWYfPRisr5HeaYvPnIchkUUCi5o
CUcnnvJUnBqobX02TBwEMyiOj4BGwBw6yhszZRbCItsx5xTukUi3U/xN/EuUFLS0
DDlXLfAEmirRNXVUQw9mKA67EN5qn2zMsr5FGHEJT0eM7FiDyd+yhuIDvfZgKXAX
QiITxycba8BUpnMZmKioe0wrTygvdSGypq0R/xapVIre88R1Y35vWoMKfdpTHCBC
4WvBzx3wo2TTM7XrYVug4hPNUAHJ/YRvHN/jUM1hZKOysaC7L42w8Hbfd2T8zZYz
lrBt8DXCuM67ZFIwMRAmaqgK5JVzs4C+97hRW/nPylZhw+b0RvU9VpsjBxH0Wfg5
9dtgAUxQTpAthik84wRmb2RWehaQDJ0T64zaYpKjGKRZLzC1iMyCJ6scfSQMfwvv
EFpg+zxhaviqsqbRudwc3080fADW2o6ZdlmPFO2tZreaVHM4LqIFm67cLmAyx3ry
v+yXAKOGNYp9n4N3TZ/cMiVhhoGQWSvrUAkRwVyovkw1562jehCXVfMP1KUL6LYF
nEBZcE9TrkZ/ZqpMAs/OHKvAQAwYfsevzU0KWSCIcLAIVQnPMcG/VLjByLr+sAMy
34JV7HQHql++ZGzKb1TApnzdXJE/FZ6AuX4NFDmWlYEwGBGLd6HUGMWuZKxggh/V
6XDWwbNYpf63XLgj11iwo3vlIwTsRuV01JtnXVQLZR1TuQCa9kcLkCFFjJq9m4vB
ENH7KjjkrrNwh4rcswObe2oY+L36vaj0AYizglZcdmgD1IgFzF/SgS38ghhtP+P3
APhh6PIC33NRCCgl+Z6Szgk6kf5Lk8SUYp4cIZLzgx3QHWtHtPqEb56w+eTG5eJY
W2u1G6IQXyYAyCvlXCTy1l7uZy9HTpfmNWV86O/fs22gw2160LjcS3AyZoQkOqdg
t7SdD1DdO4IWDgnVJC2FkJ4nFm/u+oE8izfHWxZ8YMrLZE+EVj/BSIab5thkUu7Q
W9XPqqbc/K7kvZQvH9FYj4do+lEpwMoJUEJGAHqBQZN4t+5L+80QMc1w9jkZO/Mp
edYqOo4UDNdXQ0Dl9/y3ThY/PqqYbE5vYAAKVjnP3fUXe/PUtCmt9nQt/g2h0lQt
vzYR+ozl0wYoUXlQLFtEe40d1ynfG2h6eWJTsEv0a8BDn05DqZti5ycTv60EimEs
P9B+tTyet9iC7m00mNvwXcKwPbXmQhUTv9TUg2K4Tpiv1Fy8d+YyoeQLaHuKO+Hy
CBSnCUn5bPuUd4fSVEnorZ0agwRD7zQYoU4qeyttIQB4flgvrYwkPNUUPeKXILWF
Nrc8WKtGnDy7E6tb4dM8/HJFhzFp69vB3YvB/1HETmpXUCjKT/lbVeSzXFxwhW2C
hRtqth15AjUNuPZltl54ggzDxys1I9NbwhGMkCIey7/HBM3v2KHImq16OD/nXFw1
FBRXF+mmxT5wKwPMuA6sguNTsq9XqphiYyzuB/iPmPyIiv38UL5oG18PvjJcxjQZ
wj7ivcwjyyxQKJne6rTQCvWS8nziGVgyESVsxE+/y7BN2VCRM+a/h/7NY+J33b2J
Gko7eHoC3oeYlu9bXqcOdOmEcPgRqlyYpTcYwRucf+aYn2nNt/rJwSvu2OhvbydT
lJ595gZT6R2wHSJiRSEURyX6ywLhvcGQU676z8IjqXi8x0wL7p6U22NUhAuN9YQp
KcmXmVap1XXSf6cGDLCIKZWAEPiLxtJbXkmH09ZUfhVXxVfEDJG2tJ63y2+1BPx9
+8SIpt9zWgri1uTJpsG75mHSaE5US4QjqRILz6kWMu8Yp6xeON6tkameD6dPjKhe
8u0/CSa8rmL72CDPmkEOorxhDlyl+2Z4bUwslztLJwoar+sHXriwXDqCFgANXZHL
J/YmbQU0aXcCnFkkSGxWb7uE/mkAF2HUqSi/KiRr4oQkqJ5E7BW/WXiw4RH5WfoH
JVJO1v7wlwvZ8tRKoL3TmpKQ5nycSFp8VhUa6a8kTo0TZtY0krXxzsAawTmLLVZN
xIjtg3Y/UE14WEwNmyUZUOXs98YolB3ks1+zYjtUIarOG2vwSs2w0upaKLMDNwqc
dt3WUXeRzoY5JiLzqEnb9RPVczKsPn6mqAE6lAWTIjUYAnTWExFn6JiD7X/6yURr
Y4X3WZSQ47Mhq2UveMscziE0pHAoy9O6NcxvFWII4HCBmk2pEFPVnqMkevjzH+SY
eIcef8Zh/VAViO0lhoYGW1gpJPAuYCXkSmsd85yXtYc4euLwz45coboKe4AzFxV+
ORE6BJkXcsETI2yCR7osX/R1x4QXc2eyXRMm2dhHty/P/zjS9g6T+Xm8o7Acwnit
lQOxLvnQBW/VpWRPRKJGhnthhy4GFwJI2wcu3c1ZTBmRNsSvNhWZzKr5NWE3dvB5
Ylzz813dDZ9NScIN42q2JoYN5qbbJP7ua+fIuZEsmue5eSyFSu6yCIodxg+uW3hY
+VM9G3ROocP/znyAMd+D9LDZ3QsG7+G7bWH+gT5saA9Kvw1EA82/i8ODkBKoCzaJ
xP9N6RcGyvXYbMWuYptXWFt7PSM9PI/ByaENyb5YzTlGb/iOaFSkaRBPGRQilDT+
g20JhNVzSRmE1MAxg3qoHMMPda3dSemEoAIksmVQDRhJ4DhlBpuFRORTH7FdKO/c
HCpTrpISAq/W+2v8qYVRKviiVzR76lbWBl/0duq7Jpc4ltqtpDc/MYZQfgTn8sxA
/bN5dK2nA/oJ4j9yYqpr/mZglrnCmbXdP5UyxoCi86P09NEmCZLKLCBMETfr6Q20
QBWUspwWkmfLu06uV0uBSGEsqVipY2wU7EkDCK6dkkm3AXHVTvOj3/hpmym6aldJ
yK2EOvCCaxDgt+hRyUFHhRLxM59uWprsASDQ9IzpsNPxSik/6efrxQudddGvwY6f
K0kiuL/b8iSr60Br8mbzKEHb/wOUubGQy7tm83lIyf3zBJJ4TcMuhEEKKvITAD/u
in56fGcJBdY3FBW6T6eJN4URnIQnNYzSCZzcS3AYKbGhbGOEjm0qmF6Rfx2fz3zj
HFWCagq1+DOQccjX3reB5BrNl9U9ZsFoj1hMDCaB+7piCxdcjqzNl/PW0gY2c/lG
YgbbdlfdPL2MZcN3VQg6FdciXbDH0FlTe4B+fgLiRDKGrzicOyNqxABZAmhBfgo2
2D1A6NQtKY3fJxE+gwXEO6ClGInnBwLp1XVDDCZIaZ2KjfIFAghkx2obiy4YGPRP
+osflblVSWizymBOfanSIBfQ4luRstWcg1+UvRS+KGS/VGXMeIuJ4BPBdSZgCtnN
fLvgtmgzt4S0m2a8q5ltiR/C1vXreu3EuiRjSSj1z+1BTumRXsdqHCyEenJKox5c
tT3j4LuoB5UlCura354VboHYr3pUTaFC8DMd9E0aBn2nLCutVaMHCrSGoEZ+AuXc
n4npvnrk5hOM/FMcO3dBbfUh5s/sCQKteI/7ehxU00Hht7u7j2+fk2RkST/7Fy+j
qpby2Fsf0SW6FrFyqiC5DE+qAjeD5RPLkq1DYz19O5CmV3hwHK3ZfE5jCHf5X3gN
Db5ccLt8DrkdLvYGP7mDeucKH5zeekygXYp9KHBPg17dpgWA1Cno/BLo0BAS7eey
haZlMUFVx3m794FIw4VHYjk1Crp4iZGUHqkBh+4XQoLnOPjfszLaNUSset1pLAEk
pawXMrCGTn2JUidgV2m6vtVt9zdxc/jK3FmYXhSxPFQuYMXU/nUfLQs16XXbV46e
NQveEOe4CQXGxYyh5SVQ+Nm1TueTpLe/CUQGb6Cj5FUkV0aq5jnL5k2Itlr4/NSO
tWGW2MrU2mA69HctEgKc2KUH8znnEnhV0KxWia23mWo7gZcj518IPnWH7fEcc83i
dL0YznPnlr5QAp3YFDEg/KwZOHUOs+j273aZKVi6lCvipPVASGbM64YIRtbPYZyS
M5FTy6S6oK+oOPUytqiuhMU9YdGvMGG26ueGrqjxJrQs4OqR/c4+MqTb5QtEBK7c
mTUbAkRv1aRnbG9XxUWtoqTGM6aIRQYvqYI5WoWTg6fyf6yKCv3jopLsDWQkKrHr
xIfleIIvpKPOtSnyFUsmhO3Q3zEO5Gpae0S3yYsBBGEF//X2aqZCB5AL571tJmpF
DyOeuQHFn5Wue9xaZRikwwTqx9xdLl+Y1prol5wJwgBEdRW7uStb61GAWKxZSlKX
g5QckJnvjPCgysDKAMnzwiL1oVHZkjqPZ1LHgDwL6cGRThvyEaf27JgvNE54Iokv
yhMEHI+oRZT0Gf1A1Uri4VewZ9OYvI18q1f4eun1RLCTD81/VjlIVYiok+B4OnZP
CuVHOrvRCGqnmfG/1urCIW+rgGxTGOu/+LC65YBqk3PUWNmnhBEjBVeWoGu5Y3Y6
Qa8esit4O8wr58NjbVYTBvT+TE9g04bn+1J52hzlbbsG33EwG85PI/ZFN24cvVlg
e+WwUviXSnpsFJS+XeacrLvGIr5tbqNCYpB/sHMhyGXlByteZpT9C8WvLfuFLCez
8x2HE7pPphrkuIWnCZAda8/b11mWkJsoO8fVjvmd9Y1P5zLrsuSwiMAsNOBfrwbQ
4KUCMqlaJnM9Y8IjHCHBKcYWxXTg7ky66j5vK/Zrpn4AB1w54hGA+iey20jOP36V
GMm1558cuk3Ujj/LxdNC/bB1QukvXVydhCNOgZPvCE55AhWASujWLEbZ6c6QgAyy
z1W6xTZ67982OqgDCD/8E560WqKjZmfcOMrXZx50Exqmg7xGUyBYSPdvmG3hFuXS
j/K8Ft5Neymgih2Mv/HbM/+rFp9Q910YEP1DCot/fKfv66ViEu9hDlTJ+uRQSDwK
winktmA+kygDbJeCMdzp43qwrWxKGpAR8wr4PnzxEMoQ0PUpwaA1se9U6a3Yumhh
o3Io0iILWpF/YTk1ADK7s3hSK1aS7A88x7MXeNoTgUcyk8/NVkMXqt/m/4WVw+q5
gBke+3ktITMxmcct8yiJCHi6LpcMNPloV+kaywd8nND0UXsGUgJ5cuNbCzoB7kDt
Olffa6tCsBhbVooHAxbK7dFpIhvUGcDEQQAIs5QvCxVwUJfGO186eYITwlxs59Xg
7o0I50NuTE4mcLnlEj2PXrwZxvnRwfMmQVRdWn+ChRxC2O90gPJopDic0WfsPeNk
hfp+5Ijcx5TRi/ryltIrmccWu7XqxKplwzYxFInDARm+M/95D5MT0lDZdMuuGeH1
LdKpidKAB6XB7Huxq77pI9okWCvoBF2CtWfAHrCTKyVoVt8OYY0l3aglTWG/DTXh
PaAGZ0nmhIzgJUkhmJ8ReaHNIcOUWVUTwANDYx9gxuREJx7uvMHxFHrTsmtFvkWz
oKcX0SdMy0kxdk37isbMk/tgR67ifBLgNlGSd6SAp2agbITuK73F9jtA2Ayr4/yl
ewtS8FWT+nmbCdSezfkb/ALPWo4naFfQeou8OlCFv5eLK37mBBpuMmwb8FGt6khS
NUp/ZVVfsYghewGiXikIF3u5wqcl28q7cmg6rTp/3JEs/o7/JNUq5YDHQQbWjBKd
Rcp6v5c5wFwlUFzM3P7wKpvfEGD/U/izCI4JEJLZ5wgEZRw//kjqZSV06WNzVTgV
mY8ysih6FP0bEcN+pAnCh3PrbnTQ84Bnw8E7ztU0gGBW+XuaJQFoDv7qgb8DR9Nm
ZNqf7HKMPCnxj7UruDSspchIoyprbWYEFfyQQhefs9D371CqcwLnkr00uY0YqlZn
5EJjqXNymUQlCwl1UOR3UaZaP/rN80pPdsyXj4VZCzKwXtK18YmGEbq96ezljd/D
h0FxAV+G8JT34fFgJsPJbdJB0Yqn3wZExsahf7OOPA1nMF80JZqP0fLL1q41EZiv
hC0OOysQ3txqilyjTFh/l5vnVuo9BnAGlquqhFifO4HFanzJPDBxiUBAmnB6X7F7
HLUMo6nOilkpY5sFMD+N7FA4qtoiM1+rbEdK3JZ1oGuEs/PW5E6S9NBOAB1TlDZ9
k/BBU3X6GXqcx2D3m7yBvq5M0zC3KhTFeDFVuJ2vsTMwrjcH3Clpf0ujtvrmAKFp
RP9JKQXnHqSbRQh28ASkCJSXmCenZoBFMxqlvmgmbNyHntvS16cEqj8Jr6mk4aGw
0YOeeH0gR2m7m+Unt7x+RmBtPstcmS62BqbvEQKlqSmNrNS9irRiCwKXZAPrFFjh
j7TZXG6srPTejVCGk0kn9hVQ/eUzQhr8VUfPhoHw6QIyvyG9PkbC/p5gErmSSMWi
T/g40bmNZ+sX7IXLdtp45glVwFyHBh6GkuvyCxQxoVBswGm89GlF4A1rfSoz3/UD
nF4zkdUM2mOWI0H7gOz7Di7zIrj4iakU+aX3iGOtx9SV4lmg15VIc11nUANRFmmd
EAvyDNBJGWzhDfF4sHZvM1Ylu1MnPIa8d9mbZnp6D1xRntyUdYTTv8K9Ui3gUjo7
DUhGFKt8EeY30a/6K8tjPce4eD2swWq4GIwm0eU5UHyeT1GyeRyoTA8kSfEPcJ8f
jLlgK9nMx8q2B+vOUrnAez3S84JdrXNU/HzRVzBO5vPp08gK+vRVSV5P4fqCSK7n
TCKYprwoz3FVqZ2qIc4Fz2nx4bviclNgYXC9LZ9s0WEre7hER5W8T9St2OzLS5Tc
RRfxjE8CsBfHDIR2a6jOoc/0gLcz3H50RHxTJVGEKQJYxq+/HsW9v5nwDBGQ77em
FZ4a/ViiCAn23Ikh1YFcC1dLTXSgRk0MuaGG7mvgTKaDR+s379EkTFv1cS4QJVvu
NJuNIzbDN8DjIP+Vr7Vp9Cv/db5iDzXYG7ayZjq3ySuCKWKaCUxZ0NoNJFuYSZUJ
O2x6nRMH3mtBPOszWAGSrR0bSnzZP7jCpeaK8nBgw0lohvHefFBjeQedGxfzsQry
DxK0zwPIvh72VVkZZrXddYNDWz2Bzg0M6qtFPJ6jLJV+swSfjt6Kx4i74i8oomS5
RVJRs0hn2n41WEqCdnrgRvXYtYg+FNKDRpv+vSz9eePaBGl7ALM20uRe2EcUvAHD
OO5/+HLdQBcSdzP5jtol64OWxwz569H2T+o6noVFxbe+0e1k6mG1AetyWZ5Jfc/z
R7Omv5ordHZehEci5T/Se86RkQno22pu/cZ+FDo5M35QpD+vkxxN6k2Hg7GvpVza
EfiK/BWJjy9LFvKlZxa8NzM2P9jiqGKqzJQ2WEn6D5qVjndH84eie7vH3F79CU87
uxmOmlay5iwZIotm0PZQA0nYkAYmCslYiGB8RXZZXJVtPwa/FBQKGb2e+gqpfdOS
Z7u9rhjdfIkIoc0Ni+3dJRHZOs3uONiJMKZ7DyU2VJ4k8ayAfmj23axL3lzfQh7p
cNGMHc5snQbDEGPyxTXLwkCiu/qkHXd+lNO9naZH3pf9Q/CKwhLEaFIam53Araaz
tK+2gCTqtpKB0Z2aj/VOnvP5noMZMtt1ByTY3vzQgZtWq6dRS9FkOFmiZNECc4/h
NebKx/eYD78I7qWFyhNzplACjdVvlu0+kNZPfKSQr4bw7HP3KPfjwMRZTwyz/FRX
oITf5oRWUJPnagSFSIQeCgoj243TWvoS5wkPXON6jOgCLL/pJRvWbhPnfTfk+u0y
qSwvJ5WFM8nEWm7m9qaRvEy+l43sGzlpE3qcBIdme6zTF6NIHOgYczfoNg9hxaCo
UepQsNq2eQNRMD3rYirZV0Xh8BHG/XzPKsIxIGKFJtkB0dDunpNhZ3EZpTbdGDb1
eYuvrlZmgh4CaCfgvzWqwgISQjrFULGexhhpd6z7G8PkFk8OBRJ6SFybwr1B8MHg
oXcToYzJDQjt3TLeJX9OHm+qQlUQM3fPnx1nowlYAbmp34qc7IjZYN13s6ow0Wdz
pfxBcqUyr+AG79ZCTiSVl5ccxaDmfyyDs/gUcWCypE29N7tLozfNgwKn9hD/Dyfx
wl/ZcRLV+7QbYcOLuEcY48ZXNE+m4ONthi3680u0rf3qst4Wsk2CSj++r6P3BpcG
gBy6sVQwTcjgtsDJmQH4l9Pt2+HSGgFfjtMkVztuVQUfNUksOkA33A7q15XnB33E
XH9zIvKIrVDOLKH21S9gaEUrlt7jbiGeG2vHjhs64mcGXHIiBFiwg8a7UBZkVqqJ
AZ9cZiPoL/kwKOtMKiFpKqAKa1y5Ucwr7DkEdozTjqqtS/Do82pzm36OqXQKWGJ3
NUPxd9Tym6/VsT6+uUIigsghX2jX+lsxbm7CLrSeeDbTD9sPvTiNg3IxjTEircCP
kBkRUWNDYhK10q3TUxVcMdgU6z+2afzY5RyYf8GVDxsFCC94Xw3eY9wny71Z0KJG
1Xt3l4w0YLMqp+Z9WZewjHbZ/XkNSGy3dBMq//8o/2CMVnijCRYj0kbgAViRXOPb
LrmKcOZr/DZo+6qsH9gPM+rIRfU0bhKxPt9C72SKLsuXthe70OjbiIKI2KhuzV8b
A9rx559niZQYAKx2dMtiOIbYM6FzEBkLdCeTNf5hpz3WPL0WhVQm8QZReYmZFmog
fa6vP/TbucwM1TQvGjQssDkmNhPDplLZpOocZ++A5xU8w9q4S8pK7C2eJqeBOfqL
8dAOkDKpUyU+AoSVtiU0UhyQ79e26jKZteBO1vf4LMrrWnbDooIHJjkFrt+zHsB2
kt9FWtIWRYfbLN4peV+rbMWAFPHw9gjhXKF7aQQYF+n4VlDkl0VCNtZjT4EQMgHb
lb5d0lBAFT9npMsMcH90ftLu3YXKHg1OSYflSwhOwur0crgBLcD39Dw0NQtTGVHL
w9p6uVU+fK22B0rGlBFdvSuuzdbNrbxbucqd7+rWWgNwVPZL95QVMCk6uuPhCCRo
H613rJFIUm4KTer/7NYA+V3FeuJzZIN1HZBm3yXXIcwkhIwlo6OVn45TG5qBytct
AUtAJ9ALUoqvmzOVCJZ3xbTCk9YAFw/Bzmlv54DUDziZVf6SteMEST+Textn//oB
kAGbRb7qkdy77gy1QAIgQk1frLwq9wrftREDty1ZqPt2s/N0yV44ytgUoa540Lad
wJDY4RK2aUklYY1/ZDum2H4wHefM5b0DtybgjWl3yQ5Wq3XhhOdTH8QTy7L65itL
bFF98hb6QBuOPvcpFtz1/E6/Yj7ApfhZjNpHnw6Hu+gHJiH7BXkoaYzM3B76Pv8+
bcEq8iE7fOEy2iB23td2x/WWbu6zC8QVv73Ba/ojpdIBw+XDcboZHABVeV3W5ZM7
w7/Y8E/P1xGOXMglzOaXRldc6gynrUlV66m8/sQqUKxVVikW+WTfE4hUt9S2mbQ+
WTlbXJW9wFdHz6xVmeiqr+Em0J+iQ+moKnx3UQAwPifOPoFH142u/fVS0kWrVOJJ
lGXLpLBdXv67LvS0huZj+dVMFwLOpKk7+12oSBUteH/zaked8j7EkfcLMWbEIgeD
28NcRpmVBBRrFaDwdZhMutnXCUfhm6cVWR2rDrZRR2T17cLayFtGW4OAW2fxzTzT
uDBDdMmruFX6WgxBs0Ye81yNj8UFQE2jSNhTOIjhNXmvJB5OVrSb0HRZaDkOItjp
IMsIeSNhM4EfzgSznAURbS3D7Wq7HkwEUJla1U8dC/FIjAgeLH7UC40E1V+NRkY3
Wcrr+iw0+azMRgwrx7VS3PeCfC2OBC142gEqXnOQe0Hk0EO3t+k1IJOK2CVdDkJ0
3vP2/B1+xsMokaBHo8E5Y8LcGfyPRCKbvnxi+1fP8r2YGzHzropp0i7oN3YkJjeJ
zQM4vcUU8S3qXqYIPgtYbucqTZB3xGjXp44EpZD50LmGmUVK8dSiKi/dbPgx5AZv
TySC0X8TaNN62E7tbD6ykYQP5cKwumJQj5NAJywXTSGJ3VSWL2qM4jDEwg4GvFDT
uoDng0Q/SBCyRa6Yjv62O4K4DvCULzskn7dADaH+U/gPCzVGsGTK/sDBep0+eM2e
OeOgAHmelTq0agwv2vjlas0zzJvAXyo8RndEzKq1qelkpiwFE2BQ9u0Gogaui1+G
WhNs3XhpjOC1yiR1zUPH91HWMDAfMS0PjpTEapvzSzFSLJMV2xKC5QqfaJGzEXsK
t30kt8GtEQ48ruc/hyaykVA+hDeiXbVKX5O8W4YtlS3/6MAKkdOY8NewiKIHi6uU
KIp/SRrpfDTMW1jtjyY5FaiB9JDBqnG/YvRXvxZK7/r91iP5kobCZ8/kWvUCtGqK
Pf+K1Nz1SXNaDi9yHVkIad8hsZSFRB+0L523klC2ZYe+5mympMq6/0EA5NKiPnE7
aqFxUqpaDneZTnaaJLGW9YnfKXtF9eVUGQQHUnCLzkC1wDsZr+dXoHmxoTy/Ap2T
jc4w7UnkXnqSfW+qunSAjyQGediHf9i+s1f4xy5sVBtnuDxETj1tzh3FCS+uwt3Y
o+wMtSmmVObwJC1Aasq25t0jbUhQcj03IqMPHCvRBlGSzSGLbL/sX6Z1RoN9L+jt
1ciUQ7fbS6HLY8qxZzJr+qC1mNd/dUH06aU23M72bU3qgj6jOPnIZXiOehqeD9Iq
0fHcZ3/4jinsOwDEGmWc3IOosnobADHeRSdOGY/lrKNpXQ2Aa9S1TanjM1kEbjNa
BJnNu2rMx+08FXDtHKSyxpzwtnnS0g4xssbT8IvI22N8Sbe7UZ5pUybvvhdB4tqu
o0vQiz/IbsL5LgfLCg0gEwYAMVrZbF806rJPgKRgmpEsRxHGrZTIPwPj2pScm7VM
Qb2sgl02D58oVVAZ6JNxa4Fo3VOjJgS3oNavY+pxdDZVvzJiHZrOh/W3eZ7TnySB
wTQ5u9wzMKVYkwJCIcKFOI8Q4l0YrRw33ZalQsrY2bFY0Yv+rGLhe6I/Zb4Rjuaf
8R3eRdx/NipbhQoE9QuiI1G0aNbfBi5KhTZKc4s1LHtXp+yBhRsr5hT4APFnmQfH
7sGN/r+A5Tkf+AfHao6E5+zX0HICHDbSv8XKTw3ZH7o+Bih+cH9U00sBbvQClzMB
7tPGzoHVbGvAQxOhNtgCtvs8fnNxsIztLOdi0CrDvdEN203zpVIJ9x8a36TV/0O4
dxtfVBLwitGOY2xGYw+Si13MYUMFLeSNPcW5KHuzUKkEOA1sqAIV06PKeTl6NHtG
iOoYl7BOOruoQyL5DMwfo0YGnOH49dqNQVqb5WAyBI2TxCb6aOXwaiz4zl44mfpk
/OllB+6VI3bLHuOK+cMDGvL5I1hKf2UylUZ5mMQqhhnvr/P+93+QdvPtN5EOH6YN
hE8o+YPCvpM4DM7DiyLSYy+IMkrLRXKDPc/FmXvY6vAUzGh6OWWFn4ne7DqOAuD7
uGXvafg/qc895GpunDmUeYfg7lPKLf+6SEMGu3CAOkKErnXcS2g7iGGUK0LSKh7q
/z1OFsMCDK2K6oP1zBtrhxnpXVt6kXHQlxHHO1r8UzeW91gEt05etyGCR+E4SVXH
bsFbAB6OdgGjozMEf7NAKjYWt7GTz6JN9md++6auYfQ4HYq9sXgqTbDiYSmYX4la
pVvrZvTkg0lttgr4emthyf1TSrxcRPODGsXLyr8Qayv4OzmT6HYtL6mEIm1zmVow
YoGFO31gbo4Tx2hoBD013hjIfwhcCQCFyl0iL0w49sdHcOLSO3zO977EEOITvaAP
Jx+URoTMG7y0d0yCP0mM81xr0g6fzNyOlvFdi7JptJefijbm9zleRvt9J8IIYPvJ
ksyrJq52MUddam60E6MRPkHo/gx5t0u40o0rsS0RR/6zAphHXoU1pBs18uN8y0C6
EZdS49Ul3Q2BGHGGGJWHUxcTDsbhlOd8H7/lB2xKYOz0ihSLXn/TAiw0dZmlnXOs
YnPotIryDxefJVTVXvi8k1RUbLSXPq0XphApvrcVw1oDbrZwtDJpUWssMcNkSzau
PYb7euglhvJC7aGNfx5U39i8gYw1nGB9D2W5P6iy2zw+EY2rbTyhT8OFof1WTuUw
lnBGhaXxSH7IVkdw/4nI3qCiZJxge9vomeeKSBFHtnWVUfMqq0kv44w1weICglk+
xn/MwY3YNVJiLum6m6zfYYWXkeDnJBkKi/6HsTX8hU5VwgR+gWbc+dtIOKGOZKtK
eQSywvhLOVaZ2wCACpXUDTZ3Nwc7DqA2QI63H3+YOCgAWUCDTUAqE290RgC52E72
o76Ahzov1sOzP36meXR6FAs5ZXFcN0XchcDde+pOtNRJZT0n0fvOSMzbdRFz6vky
+KuQKD/t2vgnKP/bc53pl7/ja/gy0m1ieLK7nmOoWsY1HV4x+Hx1pzp7nZRryDWf
QBZO/riUSZycnctODv3XXjwhrddNedU7ODkV7wlEm8IoyJZBPdbulRdMOA0G/xuy
S27GxDyS90RJrRf6rhJaiQGjsSzX/RUeYTggP+ZBCLQa/LFyHQv6sd/sllb2XfF7
iJG5PRRVjy6WxPBHa94fBZSXstDMzU/guA7uxDmSgxMXTRvT+O7EAshcBG+bjrwU
vpINIcaGlsm1T7EvcO4/d8wyVqDeJ9bk+jthbTQu1kU5IACbnClQteMtmTvDkTIA
AIIMTFSfH2slACmO2cxkepePE6AIPE4M6curmz287GtuWMkGJo8hsth1Selr/gJY
Ino13FuFw+lM6P2+cL7VTyaCFqo+TT9A1ajObra92JjOhAFb2QhKc8BOdlmtSjC6
ABfnbNgLsAgN8JRRonRfmO3ixoZbIP5EsiLzcDpxevIOI3qvWf61zPwHeF11U5xw
sYnrw0Alax9lSFaV8GdLbvVPS2DcHy8H7epnx/ZaRb9LrXTFdgSIqWPNTy7DAHqg
93+24hrK/1KreUBRR+FCYzqi8RXjAe7v0OaOaVZ63ghDpqUm4Np8wgEdRvKyNjsk
h8R8ZBPgXtjQ/tzfgkJ7MaGf9lRBXjs5Mhd1YdO9mK/iMnJgjjhysq18NfHNdfSX
Kw5/0YRWwEoM7ev4NGFBWf61NX0Z878SgAmcfOWCFnHrHCtw7bNLgb/IE0c4zrMm
1GdsPG1nRG1cLFlVXBDUde0uLfX/CdyOcSCrIgmilYTHjf+3NxKZ/dqr8pg8EkRl
vZiQx0hGGV2S2lbSJHpDRBS1UunvBgsK0dMcYjMybd7C6AYObxD8WeeRGLHLhIKp
lN8AM3FdjjOusQK/zDyLMwvh6/PXBSCYEy1+cP2CZ/XNiMLsLOkpTODPYD5pMj2n
LZ6YZNCXtogKGssIOpIJ9c11Ffp5FyIMgc8oqhqukeDjJu19lhSSY/OjdvElGWBk
KSye+NdBCjzzAwvxlmwo7nn0qqkN2uXodYiFA40enEJqW5UIMFgUZM+bv1+WnVxX
OXFJV78qwD5Jd7JPSO8Kn8rrrboDWn58gY58vwFd+fyzaPoRBmI6x22osD1V3dfz
yyjeN4VEwXMnJql5hKkVO7yVAuNtLrjyJsOaH/D04PF0HPRfcJQumrExGlkBUhwn
/G8KjjfRvGiAQp9gaZsDcE3QT3X0jte6VVrpqKqDmFvMk5TvACT7BT9ylO/IMHOg
3PpUOQhW3cC6RD+hiQi+tK3NoUoqti07gpeek4pXv4pYj4pjp4pft6Bh77SanXdB
9p+DjWJAMqIFcIekwmNiBG+CT9hlGphW7YuK6nmSAMtzRompEkn9wn/ftnJ3G74c
MF7w0t5JVADCB3YQ2L5bKq4i7FsWkPQDNgLOxaCAUdF1oakTgXdkEmkJJ7VNRGzW
zw9zUMGU1hqzPjh9TOJHTFNxLj0SXUQ6mSi2wpoNJ505hgtBGVpELpHqQ4okcsgy
vZAmItn0sH3xnyf6P5OS9vW62V4rVin45mx+eqYKPAX55LPbDxiyGl1l1VfHhqTy
H1wS5k9rryEN2uLf6cRw53nR9RlhSo7hMa/qoBtnGyZ2iWrCyW4PRK43B2Ew9rv9
jfnS7CXmDzxhnEIomguIW6cLDBpz11aK83NDTS1WG2kfN/6u3U1gpl/Nqvhe4nfd
nwIyvczL+e9w/RJxK2PsqXs7vRjj3pcevikSWPeo+PGpF3ChKfgd+LstNXKaor1J
End7nFEhiJ5wjt13WKK+I7lw0hWGNIWbq2dlcdoaL6XvG6a4An1x7Faazg0WA/UN
iHPN+I0qp9R4NkjxgB33BO/16KTiLO3LRH6MO0dC6YdNxGw/M7LzRKAAhlZMK3rj
6WUllHllcxdvl6GaXvVwR384zR7AfHxmxscP+QkB08tNTCBjnMVHOHzng6Iyz5K+
FlksTqd5dcOv8oK8iL4Z03y+JLarysYlDvcOclMEWyh+zvRmA3JAKrWuH1TS2ncq
akjCpbvvrc3C/OIdYx4kZvqDJ3+H30BJEVkatcC5I9SXiar6ziM9EY7pZI9r2E/j
ymzHp2NT14Zl1UwW6WBPUWQLGZlA5s3wA7NJ2GEEgSiTBX9EwieuW/xdcOmjA6K6
Uk8dIwxzCF9gau5cG+CU0IkWVZ1OvW/p2pbjKElXEalygHxgjcA/4dClHT4TZ3/z
q/JbLyw6Zz3yApqdej/Zf5StZC+w4pP3cbh2873/49dJJrMPleGnYlKxo529b9FA
kbVMnvB0i504WeVt77DwSJ+h2zbkfkVW6N94DvnYNjBr01R543TKtKXk+WGRpG44
rmbDT/gutWGOKilqkTAEXsfXJGNpEp9VtGwN/6aMm8DfBNCWH+gphbDCQa9s1QDh
dE+5K9xRb80uj1GbtPPkPDAAei7NJ/dD6CrK+22shyLq67+tfdau2wh+8HGDfVY6
NzvPjCBWVnxhbQqP4QcnIdzxEkJjRKW3OaSdvNAmsVjvM62DQWDdZU3u4WW5LV00
G7/B6fm9oMvjZXhpkP3OO3iWOfOq+sWkJlpqKXLggOxuCZcLa4HXfDzRVnSKg31f
AA+kp1LQ24X9WR1v8TP+F7EFdFEpqwq20DjTES65knFlU9LyRnJJGwVFDCAAKcKJ
y4nQW7RvDa9NwwC4VS6J7k8KWukOSOUT38P/Oq+yltiF6gjXsalKeKtXwcar1LQ6
xGHuiLalWDLmKv7mnmxJ+G8zZ9UwJtkr8HmeX0rEwB9Ap1VO7VwOR07CLLigPs2S
gfjBf2q9pTuK1/UODnBeRNjnaJed2dbdUBqefEVvm5ycCvHz0qV8+KC/7GiJMDFR
+zaz0XBBpP6/iSr4I4Of/9Yju/BBrz6m4iII9f1q7ZWv2zwLsv/rLoLO3ehEDlXn
smZp1U1aeCZqj4KsHBtMfQjbb3gYCyxhPMU5G+Hv90vI42kOe7PF3LMuVAUDoLmg
gIkpd6vU6NVHX1zf/+FLsz6IYU907EIAyYqTs6iQW8p/4uT4srQLWO288cgqB2RC
lTFh4jA/bS5YMtidRQbqlqstiLEtCmY4R2jZx+rtS6pOAshLCiQhGq6/BS69FqPL
By5b1Y6Oe+KM1Vj74BgdD9TOFByqe8jOsJ4pS8/AyL7pRjkdVUJJxobX7GCkVOAS
674begUsCzcibg5abgTXxgOfKpfoj7F/3Fu2kVUAMPd7wM5aRpJlfttFEilQ7/Vs
BXULJGOY/0KOYyPFkE7KblFlnGp3z+xoYNiHQDkrvFncmCulkCFYfFvU0YNCltli
mvMkk4iJZZclRFfWQ7XWBNslDdRtUtsvZeZfNoVLHXyE+feZ2J81NN0FTuTDI+Fj
wE1mwm50KEKIsfQPPnYiCGNn5xCf43XvP+6Qdlw+8OBzrWDCtOQgxEugowitd5ht
ZVuJoJJKo/ANh5JRya5byWNN3cFRqfw8u/0zcbaf9s8C/JgBbkTkI6xis5cek3aB
A3oAdBFwouRCtDTUxt5geCNmsA2PNn/Q+4xYS3FuMFEI1o5D3rfC6O8BvGouYx4F
TsL8jwvx9MRF0kKIj1GfgH+tcReOaN1X2y4bsj+kEet7Y0RYv1ASRL17mFHPTnsO
8tFPRMT4o7+xBcaG0/il2h/X6VhoyCv2UykTmtibvmj/jm33b0xIir1he02p9PxH
4A/x81cgMjK3LjTgaTpMO8cQdBdWbbe4KjbYj4JxdsP7G265HvMeO0Mdtb/h0zMs
4PMP3U+I+VaTIcknK8TorJTikMyLsgkGHGpsDCCXgJqJn2U6p3AmFk8eKZ8B4dBM
HORZU7DV60zmVDaziLAKsLzgOSEfwhkv5P8akhC29gDuXFPtCsSc/hvEE0qZzOWE
hgFdANoVkor9eaiFfucm4u9LkU1loFSGulIelPz/gmCcrHClaUSDdvcWEHLxuSFP
qG1XmeZLX7g7gax0X1bz9rwvzJigs7mEg7ynZjZjHV3FIwlIjX/T1bYDvQ2/zBUZ
FhJw07KeiPDM0SBlnoxemZi23GdGqdTeWyWeXW0kAeW3hjTNNWT0yYCWBTxHjPQy
el8YeTP363olqDMe6akENyFegoPG/XgGFwyBryOnUGdACIoKLm5BYgWIoTRv7NK/
tVC1OKu0HAu59CbsdES3HU42L2OsPQM/KMLN0pI5uo1/WF6uzVV57lB0IIAhxtLH
9bXfTkmHlVe25QBWUobRs1UvoCvZ/sXdl4zgrkBU9miRfz8XmFLwccSCtr3UPtAb
fBd5BJnUVS3MvA5a6ekVUw274ObA6vSxIRr3BDQmJ71PNBSH0eYn+W3QgMtquU7Q
kOkeb5kQuxUFNb3oGz9W2FK+A/hlyQlEbmfUBv/gmWQPO0YevOgBzhf+zHawNcha
AOumIwcb8reWATHWXeBEDS7ZHpin9TRRrLmFV03IAnY6pHMVAW3rST6cgAJs07XT
spMEch2WKz9hgIKJnZkheWtqho4Pux77hYa2e8W+OZbCmzU3hlDx6KQfjIQvpez4
GUkwB+eMt3Gbt0wUn3HpsvVmBmiUG0BTGRIMq4gZRsEF972FkgeZpPolX/1jwZRH
1O97jQuE18S9yHPbsch8WPdN02O5DmUmcaQRZQZ6ZqjfdyoLILiVnzStDKyu09d3
0WjvzQzqxJjR9KF+YlWe0smUMDuVjk7NjwWfyOqSsIiIISxRd4I8NlOVD9HqP7RZ
J6XDOnpZaLcJ+z/eVPoUPgISsUj8YR5YtTR5f8Rwm6aS8y9SoOB8NFpoNcg53eQg
hMuEe1v8EptmKGkyk4BeS+WepYV2L44lXwKylBjlqOi3+xU9zQ0d4IT/jBlAHgGX
ySKTP8Cuh2voghEEELLH4L7pMXfO8fUJ/ZhKUFF3YZKG12KXWPQIUhPbJvqUXf11
z8meVThqhtfXOC5TmHMZ4TN2eG0AmFSPIElyS8Bt3AFX4BQ1zS9MqA3cJIWuL2Am
/DfTqJE3YncAx8fZGoDm8rf2i/XJ94ggnpZ3ioA7ma8lybk4klo9kPXzcltxW7FX
bfPbXpmCPluIwCrw7Rt/RnI9zZTPMrsH4Fq/2Iu0118oaWXR0SeuzbeIZF9Vgh9E
BWeggfqD0ehs4eePHHkol22gSEoWD5NABgf2WRyPFTH6yb+sU7TDXG4wlZzu3DdV
s3Ba2f3ZHtYf7zS5KnNjQaXwEIQygxE+F2ms5aGQMXIgNsVG9TQKLJsqFGuR6DJU
CO/6bW8gdMq+0nCM8n+QvX9q+t59WVFu+TkOpFl1361keb5d6ErLyMU4oIdyF9bO
uYyZWjcbLCJS6oMVIEHlllB5DvybiAxL+3DWM0/I+aY/4s9sm+/zG74zpL+f/4Jg
odGP2MCY56ocxQJucYHZbEb/nrg3WtXVY0QaHdL9QwJozaZB8cHFyiZJrKTQ+0jq
0hrPlOJ6gFleY5Or2kBzeUUNy0TGnhjlHcb6eNK9x8UChel5FuOKB9ePtBvrHf4k
1dMluiyCKWS+WejkYvcg2aLAKzhMXpuDvOR6UY7ttosW6h7TbsOXVJseJ27IX5Pf
h0MgUJ9HgqEGH7uJksf8GIwlxxkrC9OhUDLw+veWL4kne5IHqYPmWOVhH4jeEevM
VSzSv0IQcGgOHsN8HPre4L1yLwQ8r0Da3z7yjGj2fPJGghZONEmI57M7G8+qxXpa
HXvOAkeTb8pQABLSUuG92BYKfYjFqqnfITtdU7pf07vtBxvTDthIIftcY/ineJQS
hc5BHZHjC/q1lDkedHGYAlTwCP4mEAjj2IJ/PZfobapkOjqgXWOMRsBy+8OJxOhn
/VrDgr28JL+Mbp04QsK8FFwHm70j2Bj3gI8A85xx12OlLETz9liFl31IMUajehKB
siOQk9eXD/4UJZdHAEapcduWItXqg0YRAKU6D0JOzjSeZ1tGGUAszcUgLZjqxghE
jck/nakOc5jJMPU2J41mwbJcNmxLmSE9GzhRmcDbL5gOb8WFNS/GbBV7AKk299h5
hmvvZw5ySEkr+ZHLzZt4noQ0TVBxqfffKAOa6rLp9uLKSLnfanzletPIE6l4KReV
hS5noysIYNoQcjRT1TGkZIDK0NtbV6JO5rG0lVzp+JuxVm+7bCz4/4YmQmtytb7M
6HYmJ7H9hVviPawm4QpRXwNFisFAJ0zIqgG8pkPcT33tp/LS9UascWFL1KV36KG3
8bOun621jrrziRsWxD3bsG7wTMdyz0eSaDedi9FsTfpNh9xIDY/SKtCZVhgSl7BQ
MSq9TnjFVirD57mfX6H4R5WiluS+WO9X3mcyy39EqrLni/k2O6g/Vi7N9kFPquMA
hKQ/lOdMhdYUsgHAf7rl0C7Fd1Qu9YuAspLEAf1/eFVKZhwzZyKCRhx6LO5R8Vpq
dmiQj9E2vWn3D4Gx3RIT4XDuqt4J+Sa+adQp0THL8atV7Ri1yW41JSXgnrizR11T
OpXXHDleIWv1vtPNh+rypsTqV/Pm/30wzzgFcUnXfeaai44KyB/E+bBIYfmLJz34
5gzYsOo8lhZPw+spaeAcyno7ifAMJTdM78SM7lFmhSwgQDFBGu8Enx2Eq3NYBoZX
qTjgODGpvQZemdYDV+jVOrLoQS9l3xwTZqM5YEaXXgjgECwfHtUquTbugGCnwD4K
ssOIj/VkXDBHbEjLEXF5974IxYilSHGD92DdQ+1zTHT4G/IWnr5CbtfsUYVVfhYl
k0MmQDbr9+qZh0Gse6Eb+MP9j84DUqewqdZ1pqpabdOouggnOEiliKRamvBUKqrS
d8AoiFcoc4qF5g2ykFSzGbq3DthiiNHheEOEocIcXJ4fp0nYO+YXewcpveYyOM8+
/mDw1VgUdNCiIAgshMlz11fDlYWz409p+tI3/tfCEHLp8+kZgQ0KDlBA3loRfz8x
T5YzgaGF9Pw6hyajVu1xnZk9F5XdWjkQRRgC6n/FB7Nd7DMw4FJzAJ1hYThA487s
XbQadZorgZpPrn2liQ1IYuC+RXl+/7mN4aGpZ9rh7sDisNRcSByp+UddQ9wRjrcj
jCf/R22EZsN9HnEhXTuYNOglZHpfrL0H+EYqnnONVW+jqDUCL1CDw1835VH5S3MQ
w7nP9yciHFpF9b95etBhL68a5DqTMDnpCs3Qb7Q5X5LbtRje2J/l273wkFBphq1h
C2JSZfMg8VOt8daN2qdSydBKVFbdnxFb7/pCU5yEuazM9nVHazmb+nib8SN3UvBd
nDVkN99AY3dl1Xo41DkwtucsClQaKlwlPxNS460aPn7f2cD50SNrn5xsxxJMO0Iy
We5I6zX7bEyIfx1lHThfFgVSEYkt9+m6jj3LvXwDxSlPI+iJ3g7GgOuEgo4FE43W
yJB4Q2ybRJOZtpO9dkEFfgvxWxnuWShhDQd+uduaYPXaMOlUzI5KbXCf0+LSdziU
J0grU5ez3V9exJ3E4pmXgx/jOgb+OIiat/fn08W5RKWGwOgEbD32Sz28qHJvyJ29
3nI7CphxOswEPg2RyLSwM2Vh9T9v1fB/Opic+Lvcr2WjAXyVb3CGuviWMRrT6gXm
j5xesmv+knNF1ohx6kLSGWsWr3AwygpehhlXS9GT3VCNVOOudxlZtOxsT0vt5vDY
eWHwOdL1yfKy6yMRZ6skfTlzTDjLcUymcIhVT2e/n2ZVNzPCdWYRHra/s7EsNJ+2
Pe2+pUEwiqFXIwMWXecPv6q5HA1UxyR2OAFoDRCDJCrwzU+PRicaFkcDAwB546lv
MsGMAFXsOikC+v+MME1mlnjJq/8Zh0MSAAyur5SEmmLUY4YLEvTIp7I5P22ZZRLd
u0iO5GBax8Zf77Crh82eBntvtsFPHReJgmEWuVfvLc/ZDZxWKnXupiXzDL7iV4ij
l7aZ7FlmD8h/u/8amGjwlgJb2YRvol6xvAj+IFjVGTMcbJb3dOHKBf9hI7IaukQ5
GUFQXk/5oSTX88m5X6C9RI8X4MT8LQRvguXQEUXDcBUD+0jYO02c+BBVm8/KbM2V
hRrr/eq3f9l6kEjk+st0XE9Df3lzqy1DH0mwvquN8KUC1ZnfrndO9CxNHzRNObha
HHG9YUcLaX+HjHTbp0+pb0QUktWRs+r0jqnf0WRyOdsK/r0J2OHNbooTX4m7YuaT
lAR6280TkYZPXrIT1R+QJ43M4zfkft0uX+8Byvser6UHXnSGB//TgKUP5JDi/yEo
crAltsLS2dCmdV7Y23xzT8BVDSTU06nEQhMqFZmmrWvpEf6yT/Zlv5eiSclt09gL
Zxz3gUL9wNGjut8cvSJbGWzue9T/SYHTwVbCmG2fynH6WvXBcm6Uk+Xrh3uaCaEK
/qyNyz4d/2yxewX9aP/bMfBVB8SbvzR35y+JKkvBrA+Pjbdt/4vzTUORBubXWQWN
n56p+QiSHRGvHRbOGItd0ggbw4bZQakpHQIATFD2ey1k1Jj8RM5odoCz9obnpLif
XUhKW1s03yj8KqPpFFp1yWpYWufy/o9o73IBFdp7/rOKxPAAZ6zkz0ptZCcXqJGR
Maqrb/eqK+f9aaQG3p3Dh51MozKCKFfzyPAiUhwbE4bjMHIDYfxy38NGqkdcEjpK
DALibjPuYljL1NCuOsEsAUb9MF1fdrdnjvpg5W+9RCgBvZXGC9cL9KG1ByEV0xGQ
fOgFQL4ZPcB3HQp0XqB/+m8QzSARrO2raXnraHruyj7UbcJP7ZTyC+IZPMYZ37QT
BymwErgon6kryJFN+sdyrCMU9aGfo0amMG/D56H+9mmmslYMIBkzEFpjW7Qjnjza
CDorJwlTreaccukSW459cSnZ1FMuaHQeDA4Ohtk9OppksfR2opxWXnWaoxewd4yE
Qyp9cHvMw9qp1t5/7tc75GmaC5FKx6j0iY9BAY4lQcQqnRjxjEm7pg6/lCvOozmS
mv/MqsalEqMvAgSfsA9H0eskudkxjFCJr9ZOnCmxTNPpRmQXy8/MmLF6eSmGUWCm
mLu4/mdrTZd6gL2wIjx7i0kKIuUBTo2s7UIMQhn+dYMvHFtslRs5aET00PNKW+lj
ceMfKY9fD4QnGlURXnu6zI1tBRIojOLgeabQqoTCeXSoYUmKvkYtKlNdjIZO0Az0
SWNHpM0NwQmUJq2rg8pWDod0A3uyQ/J5JY+x2RQD9NSuTCp9jVl6eqBYIErKgzxf
RKEenLs9Urc+BqSmIuDzLn7C2OSE/6hzbrAiduHaYVSvZqtUWyudNPlKgvB1Mm6D
DFKUOxufAr8v+HtiHdhlbVSKhdeCIMyjsr5xjdM4eXqqm/JMGR7KJDkogV5yevjM
PXwXt8I46VMnIOuNVno6ABftEQHVdrwjIblqA4hAX9CXWT35Ez+LN5CxdPEkXR9Q
8OiqcbESM7+KClQgIGI/Zq0c8kRwqcxh4pPRcwRcrbfSSw/ucrTEc8amP35k3DH7
kMMGsw6c3rO6wfoefqCn4GqIzo2c+dMZ8Q3ZLM8I2jTmHVmyYmgmjMdDy4y6hEes
6qoXKoezFAjRfRo8tNXIGsULykPSoRWn6gNKpg+XSinZ2L+PxwGd0z3hwlV+kmTa
ovjDtOoJvnhZHqBL6aZxKtU8Y13JkQWBepTlmCQQeLAW4eeldsEMymqwxQr7O55C
2BFf7gDJAD4YAWaj8avxa/dJkeqN7H7ej11aeJAMaS7DMslWCEF81AX0TD/1f+u7
8tTQI7n9JE8gh8dqYZholJ+8tObJ+NfoxnQppEyoRQWDfHPeWBmH0wBoNWkgU5BI
NnZf7G/6P77dR6cA0vLOBou9KBugovJf+ZMpvCnbFPHrJ/mLC0uwTfGnHW5W1zR/
92So+YruaoS3XHM9DfCGnA/ABP5eYVjstQ5yrht5vxsAM963Xs73/hPwh+cSa3G3
Bh3cP188oMYcS8MhuHorRh3ShwkoI7J6FOmQG4+gzZnZhTu68qXInUcFl4lFM8u5
WldOJY0okqfyhVXVVL5k7Pbl0fS4AsyA3M+2mywP97numiwyao42c++Rmszqzu/C
4LMxCcTBnLWDjEYxNNUn05hB+Y8QGYNIDwOvovB1FXVfdxL9Xl0snvnWhTyKHk5g
D/sRsQb5vkhvq/QMPov6IpsSrpoNIwSjas7pFpkge6ovisF2K/bF3zsbUGrnekh3
NfHRIbz9XqFUzfgggE1wevpwpBS9zUEVwGzDEloahRzyv0Eko3Ld2+Pd1ml8KYlI
mjZEIh6knGmXOT4ofoFBk4cfWRTYyGkz2dDxaB+0UWRXzjp0P7BbQ1r1206zRntV
dbQYNQPQiIQHftSAcnKEOazLBNehe+KvA6L80K86fq5V4NzUfp7Rfzuxd8kLzhiU
IhWx0FOensy4a3YPIjs8NPhIflUpTWnnD5lijaR1HAcJH+Pu8iEbC94G/BNUcdLB
/EO2foj3ngxSz8RD9wkMX2cZL0iySGwnDgaFCEneRIxASQaKDaeQ0R+9hggAb/km
5u/NXkqvwZSww2i6bz8jKlxw9pIBtX8k4Auh1pBygTPfsE+fBt3vVhYE1OVGz8EC
FcPSucnC7aiu28ScaFTcWieDOB84bC0QlKFiU8/cgO9t4Pqgpko/aYTlNm3xhUWr
hkMgM0VmLKbqlp9FVaKB/3Imiz++nxMA5dQzfFXbGQ8Ru0lCtPFGYVbJ4zMIv4sh
9lYD/RqO/jcob3EVsyTn7yDwykqRqFxxz8GavfmN5/TpeuR7eLkY5yjCxRwia71D
9RGM1rgYHRjctQpHIMqyGnOU6Z4moNZBN2I2ZKQVzO7dmWYWOEINdj0z2Ni3g7iH
WW/M6S1kt/G9PR+NqSG/m2oxrX/AxBNC1Q/EUVYgxf66DOfZXqSKGZivbl6EFGuG
88ZVxIFKeqzUTuCbM5buWIXcd7tPPi1R37xPqUbVDraDDqpEERuMxH8Nkz4Bmije
TK6l+RfWXs1NeTo1Lf0HDBirHHCIQdO5qBuWJaRZMtio5asGpMpKtYebXlAwXayV
73dbkARgi3OWVibhsbMZFfFYNvyEllybBeJOgwNPXks83RHUmINNHQ71B1/Fde87
euxGsiADjece5Gk+XDc7r3ZzChawU3zbsslNtj996uGfIPfbSw7UJDPjiG6BM28q
wuOx5rn6VfPjn+aOoSeRX1rWrLcdazdgc8dviDxNr1aDjFXF6hBES4mlZARVW83J
gg2J2SrvaYE0z/BhQPBQRAbhqFUrhWpFO5la0w6vuOYdLEdxBcnXZz0LP1RDf12/
B73VhFSsjd8SBP0n6r2lO/aAfi3vNkVCcJycr/v9eH1QWQ+x/yWyMChw2vHaCBK8
6VQ7qdsGQGxq+DIgUjiN0RScCtyYUqHMDnUsXyemPYjc7fAoFdyIT+BLS8nFA1z8
H+UxUOl6XqYbAN6HAnmlLZtLApflX+mkbjF5WuNGHOp54QYpvXucoyKBXuWSVYvD
lmbzJsepW07uLiSLOAx5GV9L4HWoqGMvAakzBS+9taWOySZlm5c2dhT8FupzBlGq
tlBqYgG3StOAqEFNp7wzNZss4saAnnRg3IGmP+E8Y6B3Y1dHnMEeYDinNYH5L3Qn
aAcVlfHp+AhGQYa4XsayIPqd7dXdypTrne8MOsH7optAVP6Sa4LowHxQJRr/EjxM
uk+XwdiX00jGM+2zC7/tiTWQE+UXUs4fuiT8J5/7XxFtTbRlKFAfBy6WhrUypF7c
MbAhw53iSJHMpLDER6xo7l6PiB4K24LSJkUiTaFr1+0iRsoDMIJC+TefYeHerHdC
XGeMq3cGzEQNWtecg4lE1s2e9cJsnFEMBjSKnJU0Tf7gatMJKJC7OOEPEeALCSVB
QejJ06UsCkIWypivZJQq3Rhrex/0jmgz+6De15gbRxd23TW0Gi8Ej0PkNHCIfydY
IfMg+KZT+P695o8jvNXtqgZ84sPJ5C8geFNw7DxMlkn/lkMnn1O5swFdiFYVs03F
u1N2cyfJApwSlc5nId7t/TEwY2keJeXsHsi5qRevyU+gDbhZPA9MKr3FbT/XFH7i
E4IE4cbYUL2zgX35TS6WqJhug5Vc7ggc+axAsYABe+mJRxI9e2oRCi5ftLhTQQvP
HmjK0Ust+biZMw61y81X29NvgMwT8ZedokMiJxfQUdDaUs4xlkzfyaancjGr7u2v
nVuF+1L9zmyHiowy7q/PXeSQoPmcoD7TQhTy90Cimdmy6gVcghltGzYmDTASSVzF
IAAW4V5xbteD4LIR5CVYBsy4swnjTP11S48p3PJ3FrmyEOrOk8hLWD7O/9wLboqg
i9MBNrNx9NNlc76yBzUbZpR0aFmW60H4JR2C5eP79WBufGWmd9Cc5ic4dRycFldh
hbY8yFrxi4xi+bFLF/LAyn38t0K5JTx0HrGlQsP609fwQ/Ma3WE6cZxND0X9iHtU
wnZvrF88JevohW95h4E1ccVboYu8lKaMiOm7rplWA1JzXDAbmrT1X33eT1Xk/zLW
bp+Yp7MoZ0usALLt2oQhnCYrxJ3h1TVmehZbY1qiTsVCYCVwkP2gXpI1/mNbRM0B
Qqjj3985sj7jljOkOz3QE1kaGwgc0bWCr6bklOCvHPtoCGLJeDLlGSjtxXNr/lZi
1Og7hL9g1tLzLwKQmZ7TSTfwQVBSJplIaljCnITT4dbAFnfNH6qmVt+M1uWsRy5O
LzLsc8MiDHIF5wpYFcjnVOi/zZzJLtqFIVPDcbjiQ9S9udmCpJw24c9zeA84aBaR
gRZxy3t73Dq2nR0axbsEYoALG1Vb11r0LGBPqOfm139BWfPwzVkowJAeKuL9TBLz
kh7+ob/6fR64qOFYuERe5BkOgr35uGF/oL94j++qMdBCqi1MzDXddpxGlG4ZUmz3
dszGFdRlt5Un4b7HBcgQf3QWoz4iQID4E05zQ1IujexqQYybA5k73PvVS2hBTuix
ZPqFZwzH1B7AsbAc0VgtBVBwKY/2I1W8IxHcyC2R3oGFhZu4KpnwI1m8Ps9FOm1c
+QXjtRQwPHxZpX/7c1oiVB+z4NqsHKdFCIbWyCYfNfW+0cBq0V3SPlbhl0zVtUZr
K1vDCFqa8Px2Ivuuax8zYYTx1nDCwJJJHMDI/OOkPD2BaWZMhJgbMkcJREQTF65D
12XTGbSPVHJb6/eHcw2RzMu1cApOdjYozlserLmTmZU49EHL0yBl/TKw8h7zBZrm
usnVEpid824tdBTqJ6yH/p3fGZWEOLgB8zjOV6SQi7v6jUTvZ2sdrfVuZlOZsIuF
2ZG33uVZdfVjXV6b+RFb/FuR4xUWhhUDB3icpOFjDkf7SorRDzf3cYi8Va7PB/YD
BDfpItb5V9C7aJ6dkm/hcAvw4PFDKuer5ghBp8FQ3q+XvHqFOX/fJzxmINbax2/4
MLUSzwdrprjLoGVg7HUKHSqz+sL6r9jAASNn3e9rlaSqbzpX976CVvS51zZxhhlY
kSIMHb7bgLQhG6tA8GJTQhgk6lFSvtrFB3Bvzi0vAQzouo+e+qsbnSc02IScZWNw
gCkJjV6bEXz7a8OzDmd83+K5TGL1lW5PCeK3XcBGnqOAT5+bcsVhQKKKR7L8HCIm
UkK46uBToQimGHz8H43vWpwSgzR7Ihbwcgj2yHiPl52kAYoJ1IzAvaQk3b3MpPaX
m200arjmCgtqItPMqNn6lEHLln4ddqYfr0YvEH6U3xgz/GlohbKaCA1CEF3OpBST
9cUsPMFrFeedrWV1WkNQ2b/0ZqyQMxdThYskNY4IJrsBxmYbtJusM6bPQnwNC/Bl
vhh9Z7lgGj+VFYe5KVPRbnJWMSPWzAiDfbbTDtz1ecTVzJdDvrQxpf+VO/n5BZpz
PV/sQvk86iHJfLbVsVj6yeCtEv/vErhXFMMQPonXmSCIbihA9/ChxmtKAzUs/I8N
qUCVwJcRltxN49omQAB43RQgoEMnik17zbog39/bMoYeAFxskKXQxAYM9p30S1Mp
RwG2z8P4+dZG/KVqHtFsBySz3yz68NytP6DroyXnBb5Sx95qsF+cBwyBlDk5G0GC
MX985aaDVH96+hiYFAcM2VmY4oVndUvPfQfUbS8ZGPYdoS/lIuFh/Sv/EVvJ+GR4
xF2eQ2i7xagvV9fvJYWsssZub4IdOaKs3yJPpg7KyO/RzReJxLAmawL3DUOTQGxi
+el0ZIPKy4FD2xnoPWu4WWo6xuJaYY6rPrAftSl9SoFmvIPRdQIxY0w24eKRX+Ie
lInOcYcGKhsNNcxiYT4l+BBTd4jaUnDXWYaStANffEr4pjFPACJYVl/3vICRJj1+
VkujBSHcj6v26/rIhkaVzDwb2pdIgOwMBYdbnS125OIzjJQsdKeRalSUOWMpj3zf
/OZBYfWN/nt3onF4RLjU6ZmWJyLDVpQ3sCigviWGrodC+m7NnBF/qTAglG8ugdoI
mfclQje+lnzr5MWoUFZWQXfJTG0YXHZHseH1/t93wGuZvSbPuIQg3pGnYuPfruQD
V1u+n9E913jS+NcpnxqEu3I3zmH29Ld9MJchH/kxmQFOhVFWaFsid3sF++ZNKMA0
lL/2T2F/XZmb5WWUDMVsFfvj3lvhJTIOMpX8uMOg5deTwQHgwV7tJ6fJn9pNB15p
qirsaZR5L7vjBxbI8U6MwU/NP0VI+zRaUX/phJl39aVToolQutKorLtAhKwUuwD0
+zYd3nLI2/OUkmGvo7ffECka+MqxyvodU3TzuEbg7BMJacnnhPoKL65Cb/MEpfJE
eWgCMdo90xkPbNTUl8zbl0xRICujCAdTSp/TKbnEpE2e2QeqA3aCV/L1r54aVx/b
lX6mNIm8Sfx2WQBH3lFjjmjORmH5528XZTje2yNxj2w1n9PTJ8mh1a9OFumDcjfd
zJbZt256CyLdB+/AwvZzknpLKu1zXmETc1YE4zoClWSRzK9xltXCDMpKKuwRF4HA
f9D+Zv58mQguGEtGHlYG5CHFzSkxLu+kgSfIA2y7itxDxvgoAshr5lFVWvInQUG4
k2kW0Hx5dJ2HYC1SeW31agARmU5iGUxrYasAyHYsnScu3AdQMG/UV8Bid5Ec2TQ9
EwO8aIgUgZKAOZvMlT7KzzRTyWcYnvIp0Ke3ItszAl1FKIQ4sFSV88XpIOfmBuvl
d2Ijge83Mb1zWJJZ8ifgajtivTJnn/2bpiJag0EW+fTnYQNvoUaoRRRt/XExNT0C
fspLbt+tsxuSq8vh19nRIYFnTedHEixhhC0vD33/I9dRXdB2b8K48VYYwKhHbPk9
HX3RXG9nnJNPuDfkAeAu+2SlW4J5VPYJFAxSuDbg1WWpAW/4f8YRAd8tkkj55EI2
6+urLSJAejQYRBGooD1nh2ArdaYW7C7vebxMVi8oFg+LkELJnsYaqbD0RYsvXigY
ZaGGg9t5GhMPOk8bWloGL7QAKNJ9lp3YaXfi4XkscB6fuGwxM3RB6Fcp2/cmnaLG
Jz58iaIHkS7f/UeSBE44yZwlCdsOLIBvS/vBkT47VuQewhkz9sSn3EWyPqQtx2t0
v4AI57yPMmecrYMLtVb67NAjBdH4nUCdAqdro6seSmmtB3NQZnU4J7Rc1NuMKJ/C
Z5NkWEnNMQuVXacFitX2mnDZHhyFEgD8ym5I9ckBQnYrC6W36UNyY2f9/caz7eTb
CkcP5TppmIJ2w92fJSylhO1HtNm25MfzgA8GaXf9o0O1VAVpJumWvKnE8U5KhGk2
9JxX5LS3uuR3Kh7xZ9SYfW+oSHWx6e7i8M5OFFVNqj+A1zZEcy3fRrNoFUZpZfDf
YdCcalX9ku/YktkHHLHy5gFalFag+pdN0AJhL5w03lhCyavi5HePyUlCy5qSzjfm
sziWrPZSyMxIRpa+yjXz2sDeSSk/IQvScHTMAld1ZpPb0EdW6Skmw31iUOj+J7pu
5gYgtje+mDO8ULTMQrJt/nemyTzS0u+rxDEROTuU0NrQc1L2CXZSP2d65ig88zd2
dmdAyzZnofG1wqjzHnMZe02DBaEk1W4xR6s91FFOcAAIm+yx/gvOUGyyLa9Gp2f3
aHtukS8RsJn8vPChrYwe7x7JybIHl3ZxE615su9AEgJWwRjw0kpgMzA15GvTdUvz
U052+wnb60wDClnU0rz8CPM1hO63/zrW7DhyzfHKEwXH+B4tCdS7sbnwckFYgCJo
5vGFeE+TRFIuIvIZgj26ivTcLaI0JnJnRB9q0Q71KDMrDqoA3IOr8yowymwROJzo
+4CCT0ygLyOXB4XgDth3VS8EeAlv35xNP/Kt1CmvML5UvSExCitUhTm/Yfh5ne15
5wUQI7FsgZ29eXjshdnm1pgf64IBfeUXbAino+MBKadoACVm231KPnjiaNRsE27O
JRja8Ltu69cDOcXqdWHLCelyLIYGKTVlrLD/Ij9a9nzMbyt+iOZ7QBLTNIBfp96u
shZzKVhHZ7GtIE3AHhUK9zg1naLl52GRPv536QRBmDmL4S0pqNIsq1Pfkv0vHd4y
+7/fpoC1Whmy77JW13Z9g+sg4bWRIpT/03vUI4ix1Pz8I42qHj9MdzlxC3BzEMAO
iwx6n9e8+KmEktStqeHe3Z39c0ANN2n5XCwcTeAaQEb/29oVRkHZGO2EmhRG81or
hHLahOeEBVqn9aXjf/d+byvu2+eZ4GqyZFwJjR0Z4HdlwcDfoe3UCQY3c9uQ0i0K
W6d00ziziYQbKR9n2J9Qbw9zmNTVQ7iuiRxv1iVC4HhhOFgN12+7cXsTJ9jArz28
kEIL5cvv5klO+8i5OOAyc8Ik7GZos4Wafc4zuv4e8J3r8LfG97tx8+lJzSEmwfm8
mnhgpEKR8Zlbwc91UAmy3qk/KQlDMLK7NwLnA5M4HqEVgDen25Tau9SLxP1/Y1BX
UYqKuG0yEjEJlRj0IJB/mimgGGvn7OHbkewIMrOoFu/hjBmQBus7DywtaXxs546H
bg0EaERh3q2g1sPI0iacRAB5yMM0C7siLKbnnOOsKXyBzHRTeO7gKxWG3Cg1pMOa
AOh47atG7WhJ1UEZ61sqo9wsgamKvL3Ux6p3vjHnh+NhvwgPhBHqTe+Mk413nykl
fmIPhVZgswFeyR8TeqhW3VvK2KEX+0Yv6t2DVA21nCskX7bWblar4okd12+erWS4
8z5lTofKcBgdm4EDnNr8djlVARo0Z6gFz/jNW2yUeXLB2/LZqLdbPgF23Ldj4AuS
AtTfYTNIo7yu0Hg9tb6L4uXYSJG3qgaO+kHgbgSjNprN7+aNdKoc7VMVX4RTT+xY
s9PxskrWWq3p7qCC513OfKdaJCS5WCc2twkKmNbkcdwI5PtKGa4YFhtXGZIO8xXt
K41KmflSjnsQT1abx8R2rcxBYgIn4GpioHTFKfiRlPugaHhBjt1XYp+sd9Fpfu+s
vHN2nCXuJ96WUFNcmoqtSpvV5uLk4o7jQwQU6bTnk9Ky7fm+3nkvqC2a5TVoqtiS
3vh8TdWcIgzS3PtwOdLc9LuTX2o21u4l4kQOLdQCQU3je14vzAUD9G9DzQ7go7zc
p0EXa49NOVaJ2DQLnqXqkyJR4Pu6kPADIxcpSWq1lcrdUsmhzC21oHHGMbhxsFFs
yRyitQ5lsdc/2z42GNvWCGRa/ERZgO3NkZvmmVTE4UhiRJUOFJtpNhGpPB0+7CQd
v/a26gIqwxmbtKN7dLKRe/V3aBv+pWt0GXgiARIvL5c/4BPupXzg4zObd5nGYTEz
CN5I549ZOfrMgBb5t9P+aH+iDa1jjpnc06jUgc2A+vSwH3AV6Y0qQbeW+HZjXC9k
Z/A8WJ72ojqSvgeL8gJ+u6XoPau/ROXJOZAXpma/4MzOBZlMrU/9/x9CFpA6eYuY
yxqPmf+dptWZYW9Q8MGSyHSxG0Xhcm53+XoTg0M/TcFGqzYexv1YzGrb9wEk5cK2
M14QhIktqt11gm6o6Ru98iPReUynvi/FZ88UIBTRzUiswfA/UAEsRvyuW+0lSXO4
lvITRLBZzkWy5eAFONAnxbFLyQSHVGqb5OidrDkXWcv5nlg+pYmlGO+SpN9r6DJh
Yd6CyGzxOwLYkGlTlNPXy6du/KV1x4rJUk0CMnWnz7rb2WgdbQnLpo5jVkPet1pn
8bGdpdu9dwoWzJ9zW0nEmaWCIYlOwiUIlmVuKaoX9OzWLCHl0eBg9DuydhvtbNnk
07Naoo+yrdiV3Hr7gMJtv8oSiGDR2woBqwwFNdSovYloujEkdniqHB696YdeV/MT
THojaLXLxYTnOqvj+OZ14dSqK5HwczxB08tyOw8ORfpR50oT9ggo1IciHBlezRNv
gi4uIgjJIiWKueh3YKMf9BxOliHUhkZ5iGoSITB8ew558UCIDSbfa5tgW4q1H2A0
60qBzEd93ckVEDfheWBYLhVtJQuA5XeZqHSyG5LHPopIy3vjYT7NIpyP705MkjN2
0Ur90tOvHXjz6pwVVoQIb8DhLh09pkwsIgem5CP4hyWt1Ay0gY93cQcUeNnNl4Py
tjorSzXNyFrQBR1t04nruwZV2NYayLFQUBXzrqPof/+N1sFBwQjBIbCvDMPe/hwh
Spnz7jYP6Z5IsmLKuVfzJmSXLmJw1t60llD24RTnchTplaia56bNuvvL+TsILO1R
HLRoP/obGadTv+MaLABEEVFWkAPFogSZB8zJ/8KKIH5tnvIrYiUOcp2hYfMT+6sJ
iMry4JHHlabzLhpTxCUjfdgfJS2FIgeFZKjl5DjtZweSMtl3pLkhJBfArK9YIykV
/H7al9btF4/RGleIWus79Vvs3xZiP3NJ2uyJbh2AURT4pop2nCDm5Mkv8PIm/OqI
DtGPThQsRAxYGzyjrJgr3oXEWALnGZio0a8heVvN3AM2nwmuoTjD/9nDCDepDEWp
3daMZlHa8OYOEvtPGq1Pa6VH8h2hseA/V8TmxQJkohgHFsffFaLqNsHxAnrXQipa
4ryHqfDNMdb/neYfS6mFbFdhLO99OQWqDKPXmbMqYJC4eUdJqCPJgxgWPtp+JV0K
ScdiFRnsh0I/hNBzC/+2dwEQR8Mqui7k2XeraP5fHUVXzCxI+OpyWTWGKrPG6rAb
jq18BObRaZeo5RcrVPieJMeXOuiBSX8f9fmzg1Pv1S/I5cZYgQ/cKssGm+jPbpKx
1nQIUhA/Z9UcSFL40QqeGTsUZC/FAdCrOp0DNu5dugFJ5x/XcnwLUIXELgvzkxYp
gOYW4iaPC2L1f6w0vqGnTLAcx0k2vUFTW7gBHU4W4Sfl8M4gnJd5n7fbO9i2PsYn
DfDDfDxt13RIZcCu/YZIVbtBbr0HV47NMSxmOKKA2Yhkm/LrDkbnBSuyMkavykAX
PTZCV/oXjqYOOnE63ykfhsQCrMOBPqN+xW4k1cKuje6NYUWXHybI6onJqbjp8Efj
f7OKpWeKabT5TNfMYOotG2RZgmFT5m0IC1XIsJszMPppgGmZArdBuKSM8LplWJqy
btJiI6jvtt8+txPhp9jFNYL2Tl/rUhbK/ITOjgW3J53V8I+jElMHOebqEm36N/67
kvw1fuRep4VRBzIHUJ6pWXwKQ2tUaQ76pkhzGzkSFP0dn7Yns87tQa6s7QmfQGdD
BNOAIQyOE0YbN+b89W/akTLnOUNFJyHZuDh+HmEbwHCVvU57irzrt8J7tlDYDYts
oC/dQLx4VeLRyTykZZdg1CQrr6ypWfbhXeq4qUKh7MEq7YiBDpAZdqjI8DmEle0c
1JfoPqqgT78VNEBOCxJiT169FklhXk0AfSHf8XkywiBK2hx2IkOJBbZW9lUf2Qql
wRRnP99BCI5Yym3UPUXb8cef/W0T+Mj3rZ8YEdV5dtN9fNy4whHcLa/Spkb94A50
15k6SWIjKLXhHoeVlqlhQVvNm3sddQB6fkrBTklfl6/tr4P/SSQ0kJTLTi4aGxlM
ChumAgKbKNBrIObb/beYpPteF9h/DNvgoWsMOrphR8FKp5INlRepuKRBrWnQJr/j
Y7v7AEZyVAWQqu2pGBRId0BetN2T0sMZvodpPU6gNCcj19wzknHOO9YmEzExNfL+
QLJRBYVjGmkrvbV5KS+NAVeDAE0VZZsrN5jrAQR7dVlC1BnaLQMtdJmDHMXDdC1C
2hqNrL7gx7vu3u8Np8+kLq/jQFRWilILCDPai38s/w2DiIhuINmFvUPciF9suvW6
mrlODyfhIMtiraAFB26W6kd4BaqG4J/5b8JK39OQFxmCj7v9mHOP74Ri47y9utOP
Lh+WxHiD5ChNGMyxXHrEYTc54/09NH+MzUlH8kfy0GIw+8BmC5qpduepM0Zx//UI
vVtG4XJvOlKEEcYFV3GyAmusyJl9T1RadWKcaCXHX+H+acbyDLqHiDxfbm9P7jrT
82uaj7mD+DY9phBtnIDa9BWy2CFEt950KrToh8/3mWFHO41wWR4y2RhIICHjhS5b
ORZBUD12tvGh3xjzHSZ/yQkLAfvilmJtwIJm8HmxGD8SnYZI8+L8FEPURIH2Ks4K
bjxmA5VJefV9zIXeA94TBFb18bfLIclzB8QuzIaofTf17JghBlVQnNAdtPh/VtIY
eBWiEx0fKzDrPuuDQoUY075DeXpNfLWy95ZNU4ToYeGQtljLV3L4uq4IMCgStcNH
0hX6ApqZaH/eYjeEkBfRNzCN69nDx4O+szzwu3gg1nwQhK0PjDOQ2kYict/Gfe4p
TLTuLgiBJLDARFtx9RKh9smnXxhkIoRvsNbNqBFrAp/9Ay6bBSHXIj8RWzr6kP0x
x/g2M2cXBMpGmGK8n2jo1fxGgW6BW3LsNCLZ4LOv4H99rTsXyeq76nX/APMfb3mP
K3fLUtvmWksYsX1zDArERg/lwv7fnNZ2IsjcI10JZJeTLFKThtNc6jN+lIJiwPRp
GBa/bOhzlQsSkkpc4yB02uIWokVG7rji1Ri0thOqQR5LuAakxV6+zGPpVjPgmjHF
WlSBD6hePSb4gXhqiQC6rnfwwfaJz/EqpEkTktcP71++nC1QRbiqrJJcZRRizUhf
W5m1xLWcumTZcAkGrr2QkHudtHnEztb2F901VnRe7Wamfxc/c+5x96Ih7F647Abb
qlqjQCSTo0510Zk3Dwuve0w1d2iLUyme6z5ni1PC+sY88ma6ryofRacAJHY5Lc6S
n7J5rkEtj+nw8B82vND4Uz/GZCtAVZnx+XYZvsSyOB/Fi5lc4Sb9fDFRSgg6Ii+7
B4rB51OymbN3sGOZ90P2OLe4UBiLYx6uEyzC3GgrUGWkGg5ekTy6DrxtgaxovsbJ
ScamzdFvN7MzabJSK3/MQI+AzzatMHDCIU93YcOWB0E8x9WbuY28hrwiVcx298aX
juDzWgWS3t7Twjc4a537lLkxOQou5JtXXOkSXv9yx/mFxr9qXHh1o3TU9OqOtils
cxkGVGr8vptTBO/yVhaOmf20Kjb/76U3JcmCNsrqg713Cu6ODwGmLrY46iVV30n3
2Hv8LBAuIjHpHMs8uE3tNQLCuTAHUzD08FEVe1uDWhNuXC4mJtoaEOQ1YNM+t2YV
BDiGP0hJWgDPQMjNcStRbGO+dd+UyVc4840wnl8VO2FqyWDIChWkE9APIDPh5DFM
nmbVC4gza/0o4I06pN1LouMrVKeMYzPbWVbJjNdNi83JjZu4930tvXgmVjgI7KI7
UdOcKfxVbPLv1O8rHv4pVOHOGJBORB4Z9kvywhF1Flh19NtKexkdqfpmzXxcbhPQ
Bw6TCHRzlk1zK8NCXOZHBVFO1rZw26Tlx3oQ8U7rOP0G2Wn9CZuCEwWdGc48D1tT
fCDeIEyw6OR+WplKYon7hD4AxM1xjiRPOYKu9NS2a2WaXfpT/guN+krU6+je1ui7
DIfxLMGMvzB0JBUEE9c3FvC/ZpDcKcMEWi/1swAQRAxVp5yN8bT9+YRAQoDHNfdA
44Dq3XazQRu8y39yb0dVe9B7uvIIVn4igxVtmII0nJutElydbVDZ8mFfwOCQETSu
XfS5NiNHn89rfXV97eAhoeHz5QMjKv2KdpKudhZ+vX7E2IyaT6AxwIF1v5cfiDJK
jjylKtTo7Np2hOEynWKoSOZoXp3e+5F1TvTjLkeC15y6tzcJoeMhy4t/ueRtgkE8
b91oO/a+MSg0Gcv2fCPW2PBOOGONCBBryXrPOsyf0sYm3oi/cw9squ6rae4OHO7J
xJ8nrSBfBh+9zt0VAz1nQCdsa5e6nKDcopbz0DhiY1/BC15EdDnywSCs09gi+QfL
sVCfeXeFBGP5/VHrRwBjC1AZk812CEBvIQQv2ZLrHXy4jz7GkABCCTsNtAKd2Nki
/qc6rNgN7o7m+A/YOkLQklZMXZrVisCRSveUNVRFqZZjscbLapx+wN62Eb4qJO9o
7W5mON+wAgMuAKZccaMPY1o1oFNJI4RK5cP3mKBYoGpM5cEBfD1CIU+n/AOGzQV9
QW4rk+JKv9LkyzNmiKzsJialngmRK3RL9ezL7lPWBi0dW1KJOlfK+rqedK+B8WIU
hfZ9CFnhcfqJmrPP/JLA4v1WMzG8+BEIazSciRo2kIltQ0LFpqhmSD7g3auRZl3G
W6ZjhZJq2+u/rHM+Wms/XRD5DeheZ1/HuuOqo86nXPHNDYeu+/Im1HbDQNvEgzJr
9pJBWr7drbUzVCBKx7fZTFQb92tgDtQhMB5aKWA+S4VuU/lDgvi7vjw+UgSQHLsQ
hyrtNwnO09My4JPvoeK8LsBUsNhvCUllDrR8YEDXGJn9z/sBr855IF+UTw3g5q2J
AovTFqr8catu6ypNLXNM16u2B7XXfd4V8RzqOmH2Q14Y+WNPdyOjMrc2UmN4e++R
bCK9FOhfiTsUsTWb4dPnNBW0uJ9FQAQOt1+6KBmkEfIfbnTeymoJKgg0rsAFMTCK
nSaU1WKmjDxmEsMeXfRjWlkInsLGvyy3njh5bargC2Sioc6b0ZkyTlOLtxXC7mgb
t0j+fOvYzuuDYJQ0ErQIcK9O5NcxQmUGqmIqk7S5zVf0tDJIRs2ipy3efTaWnhXM
ejhHCoJIONueeJOlQIbFzCOwUZr7F6h30WEv6IZVUBQ3RmUFealMdBd8+fFKW4UJ
o/HiAznDOv2K0fjissHJ07NegOUysJ/E13tvy42YPdAlfsolfUdv01j0HM8jIvYq
w4tuukmsVnNPwy/23sl+affkbfrG23gzu36MmtoB31jbI3N0I5QFfHs59NmFvIvi
QhVXlKNZaBLPXCqiyeSoJKDeo0zv7fxD3gFJ4N25/vV3aIciyExUwnZopsQZv5Vq
wEIHYCKkjuW5adgEkt8BEj0aTyWh3SM8CyqxV9t1K3w5XpmhhvP5JCWdiceBizZ1
5qm7TGruZs7WOu05jCHvnRjYr12bgfORp0ISRB7nK69JVuqFb+IJN6MTipG04yBJ
btlfgmcmoxURe+j7WKVitjguB0nItg4uGISw9Iv4QcYInac8TBDlFZe7ETnRH+ss
naDeAWI/dD7tJWfqPOggOYopxU/wBgST2LrG+/S5ir14197M031GN5wWjBP7T6yA
2YgnsEcClKEVnqro0wfGMWyurz9ciUte2sfaFmqFPU3JyV3HpzBdPtzVeyajPzgJ
asAzjTWEBivDpn/onm9nChRRt6i70OVkwIpTGOKffBCvMA/zqQz8BT5UU3KB5xZE
1UwhHuPAQMllErLoCytrg5ml6PM2qXG8ojcSrtWnHJQgvXrsxoVIFmrC0MsAFues
Ox8SIGux7g7L6fRrs+Y0jXd1t76yqA+AnCfdJSINEds0XGddmwTfD3pj6a7gIHyX
tABFjdigRuZBsIwBvbok42z0lokDw++YhIimZHnf+aFpdqKdJFUPpRJ6bjvawCha
QL5LUsdaZWUP+YAV8DGt3ODxcCoX8FSFXlZMyF2nSSHA2ezYwtQySm0O/ohIYgIN
P6ixAw2wv5FCOYMZSE5yDGef8i19mdhQbOiTlYPkFEqn1kDe6CdVOYQQ5RZgoiM8
Jb0NxqR+lyJKjaauTG7TiitT7E24MQZF5l1zqNeRpBoeyNkHUyakJRwUWihvry/6
r+UeWPuUOsxTU88JjAlChriaFgKkkuWK/kaz6IvPrnZEAExQIaAru12//P1a5Fxc
J/LCWRHrQLGBUHS3aGcSqLC8mc5LvvIfMqHWItACdm4p1jkyAsN0LXfpydzmSKOv
iK9POkHmsaLN8aJ0Ssw4VybewM7/s8jw3PAnjLU1LBiEFTvzEUlubb8sWHdlJIlq
CcaCveEnbp5PrRbnatmkY0Z7GfBLCwotTu3Z1xT4Z73F4wwiFGLM0gVb/lR6yTkd
mC7sZ1GqhvAhOCrJ7FAVzivuGNszzvrlKzqF1vrhbB4mf2x7qd/eYLWmzO82dLv/
i+rdzO9bk4nn2HKMAvjFsEe0Gn2hkg8wdYVet5J/EMVKYZVxRwzZdzz1WbHcdKdW
q0wbmMqvp1IbeiSKDWQeRvHwcHk/s83iEtjxCYZtO5TGlZE5xRqZAa9c/4K9/gLo
+fjnuUJixToq4kFHVOkljA9fbfPbfwNC35XwgzAS/TO3dAchExV5xEfeW0X+ksX1
fCk0h9dzhD57Bl/AmlE8PyfwKTrhAIDCuILzgd1uwovQquZC7DbfrcxFBHtPYBSP
hov8jcHDhDzPkizj/1rYbhz/ahb+BD/zHQ4BvHla+lOse1OsFWqZfV99zjwSz6gi
j/Xsg/tcH5zE3v9lYw9eMD3nQAHUScZsN+ptIEURCskFK/ui2Fw7twnxxVywDMDc
C+0MKRoiYoTMN379FzOgHVQVmdDJrXTZbvcpeuX4McuuKoOIEicrRIcboT9kukj2
9Nt2ZRJCVte26Iu6O5rdXovaUgYdOOWWVg5WnCoKTO3IbU9FbZB/+YNSyrNuPnHN
WCJqwR/fVk6VidbKuYa+AQ9I9R2Q6eP4awStZ3ohmkcw9PCBIa2vz5PGzJri5O+A
K+oDOmpLU2aWiFc1wBLSymZQ7iffJ2T4qW4aGBn30XtzJhO0ngmgKqf7ugwqtp1s
8IHckuQoXbOlYheP3shq/6L/2ms72SDzRYDxMK/gCu6V4vd26N5XEs/CYKjF/+h5
lpXRYKzDWkx2Brjx3sizFX6Jg3XnurwiHBrXFuMXVhu8yZVP0s2WO/w399niSol7
2qFAEkYptH5xMDUMXIDnDAy7TV7sBDysSczfePaOwaJVGX9+zbgfQFyqJKUa9P2w
rSscnJmijggXuN1kxJb/PtaD1UKtoDhuGbyWCKOK7ZeLxrSHRIZJXr1mftF7ZOpa
O9LgriUM6vnbLbwnP9O/uQZLC3q4QKY/NqQhrGH3ZaPNGSFglJkXqtU9/6fWOr6+
/57661ARVZcnMEOEhOdfMmSjsW5/Z/+xk6u/1ATtuU3jQNJ2WMWNatt7n/ayslSR
fZZohrxnzGU/aUJNZQl4pJ/Xa1eiXKYJ1LwmndW9Ct0oZ0rT+JACK5aZoIzzagCy
ksJw9ec91wyDJ809GQHbAXTn0BmlU7Rn5VsS+WC/VujjnCmdaGW39fO7HHTYgD1n
4KeghcLjwlQyDlIeICkKDaKoEw/zS4yVvwQ7zX+Ux0645DHvtHytFpPU4PEE5bC/
IG+9EC/xnUvRUs/U0yjovLg2pFul3j9OKiWPEn154yNPAMq41vfTeQnHAvk8Wwis
rtu3gmJPdN6X2js3Sk2AeH4/q4VKBWXqX997czJTAGS29EN4jioGcXVzvy5QDcgk
Okck3A6kD8InOMZMPX0ujL5TjGpXcfmWF6Tclbw45WcGIR8hR9TcFSdPUUUgZvDn
faJuKt/VZVW+C7S7lQNSfjPhi4atrqmFk66DQdTxTA0T6di8WrM6N7Da70G4pHv5
KG6Kvdk7I27glevxl3y5eqS5I67tawtKBOlknqZ3Ei+douJB4j4NekzU1Zsg3kh8
FsnkukghRSNYXtuuL4hGWZf8qGH+f0MlrFz3nW9BLbFrMUixxK0lIfpooIYwRpO6
Mo9V8YNGW0MfbLTjBbmdfl5EXhlWz2Hvzo3lUA/rkEUj0G2FdjgL8rvRcojhxqMB
ZCoMNvXR198L8Zo2JbdlWyAmhkpZVjV6CE38N0zrSFxIHg0M4TOzQrzWYNCnMinJ
jrpb/hxzgMsS2afRbBrducZAvZYZuVdMubCU6IWlC52NvkEyP1/i0kUxb8L/EZb/
Lt+DN5s9cdlRMxH/+5DTm30h/LhU4Ui5Klgsl2GcMPsNsI/W8FLV0aKwgOMcP8DL
cfBXrKfYPwaGym4oH2hfxR4l/iB5j8ACjBBDIa54u37m5fLmkKV50hebmpfP058W
kugeaAM+eqSjW9bMHVI9fcJ8chhLOZ3xPYLZdM5QJowSW5kOUpd+LqVyW+lviWxv
j/4Lkk+NZgjbeAv5xOnQeSi8JKL8boHT64fY3M4y5yWgZs80CbIxF6HcI1t7gAcU
7lqDiC4igYae5Cj9UOAWD69BH2IBXnvU11PmiRuHfIVICN7pm/qKQva2k5s/mUng
t04NGJO4O4DC7EpmmTV7bqPtW2aQaH4xmmJ6NVi4aqU8+qdiDSXfSXZP9Ou1yh2P
4X6sSzELXviIiEbhO18kKP7KzSFGuOg58Hwov6okoRMZDIeh6+R/iqfX48MvX07K
JxmHebtYmVuWIHqZzurCMjRpyAys5p2QpVpLkSUX2Vg55C1qf6N0F+NtROZSN2+G
5j6+WCZbERU53IlZZCv/BIED+c4b0svNV39MoZxjHhva8wFgoudyhas+MCoXlO4N
DQC9cNMC34Baq5G44HgjVIXv1Dn5YkM7ymGfDctiaIuJ56YBGchpxusxdEgA9qdD
TnmxJfu+XJJXy44dHUnYXfGiPhPan12H6ux8pZqm5J7TRVXzQjI2TMMeiU1PxNoG
ZxzEC8aCg9NJnpxDhfAGQ2GU04gBwdomLP7uCiXd+2ZQ8O3qrH9L3mMDfJ2lHbSq
2JeNscqinlG532CnDxnqlusjWoFo3OWnOt6KxJlSyxmGQ0Mix9816igO1Lg9o6+b
pKc7ePioDaVFGpLiRNJetxwEhUq7HiR09LilW6jMLyizASXEQ1L08Vig7w68Pfic
IiH54fbhLmFshMZAzoP2kxL8yhIBnSmy7CgfbiriwT4ds/l8zyofmO+dTZD5Btfw
U4SmbHMUxSFn8ylMkwD0Xc+MBR6HUqLV5H4CGTjb5UWGCSTjYSPqSQSYx0kiUZHg
Duh5qi/h8A76gbDiQoXNLNYa+0cBftAHXQwCXAbr2rIBlirBpiH+3Vd7L6PftiPQ
4HRL5BM+1N6PsJqPN9lkGhk83YXw5S5Ih/DnWku/5nFRM8CqnXB8+DKAaQVB+S1M
jbQkR2EQhPvbj7+dHZAhxs+6uV69OCcWrVF9O/FWcu43UUukHYm4OpP2OAEwrMVz
GbvwMLoU+xquod+ltj/cijqwEUHJsSGVy63LJCYEOWjKPe51mg8dbyiolt76FtOp
dklufgkYE/hxLm2OdoTxqGaqQqaDVv4PBKKN853i60KNgkBxXhDkqCB/JlqQE347
UixS2G8J/tGAs8wZwjWnTTmZgYN2YRuCzMiduyvWu3ghb4waNZF3LEujSXv60QSz
qBG8R4u6IuI2FVkeZq+bhohbgzoQw2YoLFZ6ZQFaN3+Z9wr77CbUL2TMUbvsbAgp
nUc9IM+c1yXMHICC3P2beLvQhX7bHT43jxSACq3lg3Oezx4WoxOOsxhit4kjwDWy
xTwcN3yNstl8pGE1YGlTtyBH0ioltBN5XgvErb6vq0XK1hTC0C+6espYOISKZG/5
sUeUZyP5x4RzABKOvh1HovM8HBqDff04QmYPi3IMjXJqBNuVWn1KsWPVXt7NU3xc
Ee1S/WOedssJoJ/Gu9pNS1iBeo9PRarDhK1pBw+K/9cwE50eiE3t+VthBgmJaP0c
mXNNRqrOJe//PdwrBsOb1sDfzf/wTDZvghOW4nPVabN2ADFK0GaZqBD/a5nEONpK
KMi9gvTKCu9G+vi1yof7Q5xQvBlY4p2MMyvNO7mOA064/mk3A/sTszp70Gg7UT1W
BKAFDYGR3jY2vrCz62Sq0wqO9ZWFLiI/zigMw7UwuqaodK5DmT03KoIFA8vSQoth
N2b5X8jV3ZKDtx0LMuJVTloZSWVC+vRV0B9hXfniDdcuJ7zzRCrKGJ8H/PrymR6Q
wUlLZ6nSpc1xO3OQq/wYKyjI4kdMLyK5G4KZ0l41a4rvoDo7hV3QUnQA4S+ymCV6
g4Fc84Kv1eKxhfCJQx9L5dZUC/49C/7PkOzmot+upZ5+4q+8HeJrfqRBGIu56qGj
cxi5pjuArmzZQJ1o0EIIOAGbBSxm1TYBV40khzYO+lSve11B9yhv/2ACga1flh/g
18D0ZgVhY38QXhwt0k8/I32vpkOPJl+i1rejz2voECmFl6QauMcq21DZHb6r/uA/
4t0HEzxF3HBOYZwranFgrPlW1yMviiKLEHJIhM0sFe4cPdFBBcN12StP0bDsTCor
pjtoeetlARtgbLiBzodgqwKGCBBXOhwcQ0QO8YL4bWrdWkvgnYTmpQ2zjpu0rImb
UUmFpKtUQn0XPMMwyH2I38B16EoK3KkxyFr9NyQe7s8n7hsRsCOKgmgGciaXnrld
9RURXZ5tfbWieVwhwRAS5+8JSh+xzhZdPn3vhGJxeDdoi7xledWwKT0P8upzEBWK
l08+7kdlzbDmVY9TU5aixG+B8K72MHoylCdLazHzhxtxXK8dLUwywGNIVmlha6XU
iaJMU+HI/NRpl+1f6qIROipNnviJi26jrYEeULGa2TMapDFPJAGIn9DCAStG/0vF
LkW+8aUYJ3qPJEI+3fb44i7sKZUpVu+pgPsOlXLvUxxYRiKwP+edb0KbcHXzynIy
B/MiiW+AlE0s6KNbotT2nt2TXrjTeZVLHQhlwXF/LKf6Davlul8CeB6kG3uJQLx9
B4Rk8HEo3zl64RKY0DZ+bVimP+Y9Pnj3ec5Z3xp02+sYgPxKHtd2FYfy5nQqVgAU
axQyCGjFBFdgSxo0osY0TT83vt0t40WVqjhSwEFYybiQ2BFv7uFGVzX6G7Rh9SNo
VhB0kXgDSnIPESlCHsj0C4sYeyKSpKeqyOjoaqfR3yzwmhC+L/jqQgL3kB1ovA31
TZyaaHj7c2HMRrvhkBFlHdsuJDLHDLDsF5OVkS7wX1Yhi/kMQuKmC1QMbry0mdR3
NBrGXlFMwxLoNEbMw/XK2EK17cR849dmJGZR8XMBFhwZoeaPrJ8K2xghNtEFuqvW
uaaSAhFsvljbkdFFYV7iBMGgHIztDlsCxSFzCtEiqWSsI5ndGEj/YxUdZIfGvHHk
fKwnF+qor+RwHQfeVZiZjc7hEgrZeGXf+cfIw9YCcqp2H7t1/w4T2Mxaxze7ucea
/tTfn6eeRFSW6zPPwXQYANmQW6rb9c9OKxrxJAt1ouNxzlcmGXl27ItsYRjGFwG/
9Wzq90eQ13Z+i+NAr83LvRr06lkUgAkCvhig1C7EARUMzFL1lAd6YmSpAlfMOXor
Zxse/w/bTNeYfBJWfTm0PccTYmpHuQmeF8PAulbIt83GROXTocToz+lokxQOd5+5
2kobkPJxYEs3fbqwrtd0fPOR4ZcdKCgsPgLhL/o4fFhKNJezRzKs6tbswxP9FvWd
MlZKzxD2oIjo+FGsu2BoluNSvRTOHmTiakm4BqEK83Wa4JoiEgclHnLMH2FPvSqG
y1RxTnPam4NCCXGV0GgNBwv+UyynychOsZBqiqTu3eMWAQh1Hd63k9Q2L/PP/4Q2
YMvMukggLcuJkhPB6snrD2dRVzwmjhnI2YOq0wyq48Y2FMMqPZedE6Io/IdHLQw+
LE/nGpzJjGn/ZJDgobYpZxq6XjxcAhLLLHxewZIWJ6tIPk5zj7D5+ncnHW/8FaEv
jGHGMiLRswSQTEvG88fsZYoaW3pSFBQpv2av3w4tbHm2M9w2FfVkXwKSZyRJKg2y
6TMTNMp+wUFqIAHoeViCHgFGBlnqEQwSk/xlRfCipXRRvycNggAm8yGZrCw1VEbM
4p4JfN04F5/GNytZtuC7wNDXkY9mPI1IlJxLi7P2b6ZeRqfNdRTjcZQNeTYQQQPK
33pSKLv/3mOwQSg2g2qnSzZfy4hyBtMSiTvC6DsCjPSQw2Ohe9Goal2EAl5e3sun
tN7ImGYTVJTYm1ud/mZM2t+0OuKU2LcsgsRWZPE95PxHtyF8eZt5/BMXYuEsCGnM
7LVeXakACOWAy5dBBA9kK1L9Y7EDPrCZtWcSXQYYtuXasn7hZfuPNt0rfTTJLJpm
nyT5pgrOMjf8jZ5eYJEXfd5682LAnOVWw+y3R13+/kXNPdxWbPJYcO/Ys+e0YI/8
0ZeSs2b5kG5MGq3Q2uN29rCWuOHvqUd9Xwz7hhEkSX9JXgo1tii/OuX6kRwL4h4E
WOPWKF3lQgbnyO3ItQbdUD8uzZomt8iXcQk5cqADSPOW16oLnaqOyABeo7EGA0XH
h2Q7QDyZ0KtifFG+ms0aABTw32XHzW9wAl5ak+sq/FDrNtA+uYhs42dyS0rKbXKx
B6VdxB7V04o2j/kcBNnHroICho2fzdoCZiAh1mGZpRNfaPpEFrK4+W7zlX5H5g/O
iQBwhfST4xd5X6DOgWJ3X9fH+yYsFoaAQfhDO77to104r/p/Hb1pcJbrB9N6nwvS
DL3/A/g0kjzsIih2i7Lw0sK84oXGy9oPKGvUR1W4rkSv5GDwhpekeHsBpv1ald+m
5O76AGngsQuaPKjqSdaqQR2ILRSOgfnZd08dBQkfk90dDdn20aqQmy+VXt0nzH90
ZQ7wqHAANTknueYgKEDfNkp2Tu4bQb29mZNv9TIUHJchhMK7SFvKxKp5vsUUhLkx
ajfAIr2lGdutOIq68ud+zUpvneYQFpNQeaUijbQjlc60+lqmkI3A5B/6yt4NRyR0
KEyZmqzDpPZqLnc/hJZZcby3WIlHfYpgi06puBsyinULRWPvhNIWYado+pFNRvQZ
lgVI3qcRKNTnpbJo6UH0qS+aAZ2PcFtHCx2gSVoPF61+/ltO34fAUhxDIJub91b7
ncz6RHJcni8/XRodEbn+ArTXzbr+itwaXYGmjgWA4inYyxaqYnewmcCO5GMkyEj4
UITbPRcxeHV+kx3NQty70pQQEcAtN7py1wGGwXP/Em/DGhdDN2M1pdnNP6GEPoM/
PPXiZ3FT1fRB0p5NI0ORTndEeXm0EdClWfmLjI1qF5aWJOpYxM5aPabcOrf1uNYq
UqSMkEs7XACWlXgu9aaDMEtNrWEDYMkvUa5cLa69vVC3Zy9l55KOz4ejZtDZRlqF
3exhm1lwicTIz8WwfXUrfu5i367MRRxS2Qrnk8C22hS64Xt3DCzPI5KZnPJ833/e
jbIqDzSkGD5n8BJXNm0eCXEYFeAkWc8zghwVWkk7RkTfEYunUQMVhX8Cq1I/ErDC
wXXYsHUywhyMBZH7iiHvDDC1HkzjBYc9VmxcnbQUqcFenE3kwh54Q01BffOAK0Fj
8PIGuVcrxrgy+HNK6c0l05G1OppqeZT2tx4MtgRyM+lkYFE4exy5jNF1SK26/rP/
5haI5v/RKW/38Zqsp9gl+WkzlQI6hbWGSurKWI7nMlyLIX+NPk1uLIuI8gedoBHq
xtRhIDY5FJZZGqimTfCN8HlXg3h0g1lMJIhl4BVP+Hcy3VPic3GK+yFtXfp7TgLd
K6VTb01RlRXbe9fCcTXNCEUfLGnNR+QWC7SFvnRdFJKtwO0qNut6cS7+12xHsoXO
SnmT1jqhNvWupccmc2tZ4DJPTZTto+G4xDoGf11nOfPfoSKhFtxmEINoK9IxFpUv
ALfJkikifPpUpdawSfnm/zQdS4rv/4+rY3Cz4ZZouwJKamoOY1mqagZFlT7Qp3Ws
X+gery/Wi2bM6jpp5H6CkzgnFDwQEOfB+NL8B2IonS5JGqmxi5HCGv6osuSHOSRx
ykAlnren/W/G6LnWAsmKHWUAOVPX7HvuBn2QTTr7Q6/sQhxvLG7YYa2zwUrP8hre
UESzc8wjIDhlMhHGGnhryIGsjLya2TA9NnJUHR0BupU3Ty1rvNz9WcnjR5bCVKU5
YhDetrtbIqrgs/h8J1tTtWmVTKgAkrQAjjFjBWqi2r7F1BWIu8nCLF6bR/P/axAD
1MH2Al6c3Qnz5Zorq2GlEsQqqZrGqnZPHKmzhRi5vjvNxg0clM9QLu5cMi/gsh6j
xGZi5peZYU6yMXxzQepf1GOl0VVYbx6TJXhPqzGZjL2RTEdLjcxp9CMYzArgl0ga
Qcri0nuFxyy8p5w/EY3fY1M1Mkw//SlaT8V/a8d4Vro04gBypYuLaam/tQ03m0Ww
GyUyGZYXXUTTWkchjwKNBbdbeTuBB1LmKdwdjKYnN5p6tQK+LHopLQB/O+mDZWQU
d7v1UfdNKxFwr6RjZOt8tO8a2VJP/m7fqI7Srwrqb0jobGbHWAA6RD2nXySc3P6g
mbQYU35tUq4XB0OVqKKhKRe4J7PT5ckx8Ovply972giBaqL2mhP/UH/HXW9WU0fc
VevdIWnE4lywaQ4U0W4DczMd+7WCbqoRJAFbkkTWUWxtvQMcGk8mM7FXdeTOReJ5
zxzf9fv6bKwJrAVq9wTJKjP7kGIZ0bjrkQffVpmFSL5gwbMoqAneWlN+ccrR/H1L
q2WKSAnaTkeBY20QBuYbxHY4/AHeQDZQrH5FQuk35yMKFDlS0U9FbmzIchIzJA8F
U+/aCFWOCbP0ULPzMg2e+7niMKDHAI6JP4ChS/kl4HAwItUN+lDEIOM9mac2JYLJ
M6rGk0JZH/tEBqRuMUh/0SOSOTr8L7ZQ/ceGExMUV0fn3DcNi9nls6mLj/ceDurH
rlJcJOAMSL8n1R2fG3KVJRI2flGv+pA6beopYkb0z28HFbGoKCm1+z+Oxlr3ki3Y
mg+C0sPdzhiahZmSHFOh6Gf+R/+1/TTy35f6NnzJ5yeqiQcJIkkLsrvKSB0O3cw1
53Rp5wy11V3jPVxD+yvknOQKKsH2tbedjGY/MlJtYie7UlzUW5Tye2oPKNc3T1up
JPiIR42i3shMQBYbMhTCIxo7+jYENOMhSaxRz/LsMhgIWyNKD0azMc4RAfgSdvLe
OBjkY9N3FcLTxD+Hhl28O8wA+QGYvS8mrFkfN3hgSk9PtlqlPL2DEiQ9aSgW/9AQ
1A6Arilejdd7uYeIO95dhkW7+J5HC21aa2rsk70nkD4/ew87HrYZAC9I/8GOIUs/
RsV01Uyc+i647Hzd7kJqzlcUb1Lwnqa1eAkJDFK3CHVz9ZCFqxhg8I8hBlKdMHIW
xXIeSmkFyM4Rc5B+nMj9HnCOG84q8Xv1jGhrJgGJLKV2nKODbqiQn24ggpUu6HL2
aROhyE4R0ZHrB9PDJCdSbqwOW6wM8EXVUUCUXWwqg506LkpCpfWieSqBfFkAamjv
bjyD0bIjsN4GRfZTP9yZjmkrYtja+xo9oJSxSidGdM78MJTFpAnB8u4W1beTe5eQ
Vbwfgt7Ql5cmrRKovN9yCI2P8jpj4ITqxajEQX5DhPs6mT5rNBDZiS2WVx7YUS6y
ZjU68G878+bwmGxlWCBVi0EdlOVzRT8OVhpyCRp8G3vmjhKOFUp3vRmdg3EJ3Qfl
NHF9wa4YEPv9NrF0fd9GmWfA9SyasiCjawHMbU5VimQ+MRPoy1A8YsHzGEIX+7mh
YfcUm7vdOanQVOt3Kwgv+aWee3lA485yn5qggH1VX0QDfApRpqy6j1I3ZsjLZZEz
L6E+N2uxdFKbLfbRcq2i6aqbS5awIlZJ8IUN4JnYmKpPU1V7wqhl3MX5VJ+0th6r
g0g5e+g2MTvNV9gn69J5KrIexPKb+zlN5QpfqINZF35pLKVGDNJdqfE6Rsxu6bMx
1bd89oqo3VcG/MC6n27LEJWG91aRTW5uyw8I5JL3zDhOHLwKMIvxB9/Np6wZFxL2
o5idq/en5ps32uUINqi8mL5OvtPI0Z9iIY7mCdvxwBLi4yMPF2G6lexvOKR7D+hg
pC2NwznblUtnuAtzRDz1AVHXwaiTvXqbkcpOvj7f3sxG/ZaSOjTWzdeMwfONhboN
nn7PrLUga94r68pf2UlWV5DPh1neVxqaHHH3oGkGaohLsm1UfgNKwEhV/X7BjPzE
QEesOd225XwsVBj++uoRf/PD+A3629PSJ6f5+6aSN5CJ0w0bQqYoOaRVe8+bvslG
nfgQ0DsRUaguLpBk5mW8SQ4303WCzJ1oRCCeieEEm3D0blisN6H1qZAjGX9WoRpH
CW5KCKPTqvP/OZcQKedXHPDGtmOgeYynqNd5ESRrqnqvgmn2nASleio58DBvLkE7
49roBTy7Wa/rAkgdjBbd3nTJp4MR1b4h87aursGgzQjEbV2QZ3PG9HQ0EDdy6j6g
BujNWGzzGBY4ubKyu0rRrTAx1DcUA3raRTBH9NOCuCCXFymhnRXNvni2zLe7/8kj
U/yDFiy7dPF5J1KYdOqm4FcyfeWCTRsJw7nBTSpoIh3BYHPLfxSEC39X34Gqjjnt
8RDCxOoEwXvMyLJMSiT8hjuzBjKt5et8Kf9LrDSGXT+W9O3494URZ6rC/EdHS++f
2v7sq52Lyakzkdwj5SZ78X7SkTqKeT2qLaGAVK5URg9p5qDIOywhoBT/E5RwcCDZ
A5pKRGszFrvVOc2OnDYGDu6PLBZFmb4aDoEkzYALVJyo/CQAsD03NsTnh6pHVcrk
PV3dM/gQ8gZsSWAEEJkBxqfsinHUHAKiU0xW8XP8EA9hRs14Wob/cyXMn2kdyUP1
YWClo0BPR73Wb0SmvDRGAute0ysz3rdJBHXwKzn/eN3+neZ8Ly4NTbpbu/AjA/LU
YhSBskd/prxpoTWA5vAU3fxeAkfrxG+KaZ28u6J3jyeV1bEA5A0EW1YwTmWKpYf+
fTKcl3Vzwlshka95rEDwjsdsCq1BoLJ1QMoxTEW4pXl50jwph4WWdwsQpyIV5VgB
rKK/dUGyRdnabHDOCcQpGxFkNhGAYM/VONFeTBb8jxSlyJbNY4LtTRvugNKT6HX+
A3/ixwpnCl+Kxt41EXYzGu0HWkniJh5A5EdXk8adpxIYaQ8qpXWhWJw8p9PWrARA
BRkFCP/XzyvukJX3Hev2XOtI2DZD98L+QT5je8C+qkEAaMGCSRQHcdddCCnHs42r
iZJnGYFIMNo2HnJ51eMTLZzluklCkmpD+mVkuLqJaWaKAT5qVGywMvbr2whVybvn
3MwuEjvqbG6nK9ceI+3X1CiVUoI8bhjfHx3ho8xRekKDq0zXVBNXsQTV6U3kIeVs
qAvexSEUDCFxewQL3irKBVwBy9QsNCaqDqj4YHv0LqG+lJVlEcrXOqwC1Q+Qm0oV
5fFegzVE1shCfkEohDQpnCRG3df2AcxwO2TIT6KVI3V4JJL14075nj/iHZyI9/Cs
2fMb9pbyVZpSqNgRuQAZY90xxjXoBAEuXSawGWxlGlcYEaHUN42U8wVwfDtbiUSo
fjPXj3P/W81Rpoeo7UhOc9berypdMzFTmLce2W45ikkE5C3bxpl/xqvXBlWjRXMv
uIROqKx2/cE61uFAx82ejNENWXdQqMBAePcJhjSAOC52QIydENF9LsmE8dIyCQMb
8oi0a4aWoLvzS5fa34EtKk4Z5Sct0ACRTbGJw90OvDO2NcbBhrYGcfX9uExNNHAw
e7JdMP2IEfmp+Apr5+Hz1AzisfC1lmoi3u09d7JfDbOhVo8XWaUcSaCdaNGZjNTl
BbRfqM0QbUoDxjh35i9fl5k4lhQNLSu6p1VwcdOEMc5/CoMy9Xsz3Jm/MXI5q5k/
uv2dtyNWCRBIpApJOmSFvhdgVBg3zkE3DKSIgawjSaCdyfaG7Cm7xubsLFT7wC8G
erQKuEw3llae8bRcAXXZoEBFD8RtEVHyQSqZyX/CSDwRpMDSNvOq7hz2HZPYxwwl
IWU2MFDVO8T4WfLhSYrTGrf4GqYdorQKArPB6VtUJ6LNPQYznfxuZN7TWOw97LTh
mPf4tRLBWHB9miebztVsns2fpT0AFAQXP3qCBWm8YjrCQh3bsOHcvRaZGoVzW84A
Bv0vGuzHclbT6g0p1Y/Wmf8z32w+Vm/gDZGfyl3hZ159uoOOTn2bmC5qJX/f1LSW
fMoHB3KdDRFYbIiy/fqftcho2N1+7phqLagtPpmapvh+ohs1i29kIfl2OrIBoBFY
rUr9s0jaUlL+JgtaZxm7zvEdE1EO6U38oxGmlmtNbySf8ZE5agYYPIfdxx7NMPDW
9Qt/lSz7dA+K1afJzYPk2vUlrOGlcj24NKlhUTYLLHZUKN7Nci4IvSV1XL8Emq5a
X8B2hY1UoEbO+tyyKnNUNmf0R9FIui5pxw1GnnoMdqBJarEjM2ymTNUdR0AGEaTi
o4ZlNZSLKu/FZGHxQsirFF+GX+HA3YoyxoVaT5CKJc80vI/9DdHHZ4n+oF6MgmKp
QhEjR9652bBSp309s8Ej8OinSb9HTYHJ6e4AHQPIc3xd/UVR8fd/7km8srfgWGcr
SF1Xo3UdaUMlINv36i7OIugZ5MFq5voM3sj7pKKWYbmzV+LMPiil2ZCT1EnGM6NK
3lM23hPykeWsTyirRQ3LFL6ia6W4zjLpRGXdHRqkA/mnOP3tlZXaWbYSIR6luGhi
pg0o+HbJgtV/9aBuTWUXMJ9bevEjY7Xt+JxdJO5fKO7kHlxuJxf4DAoJlcZvz/SY
hX1Ur9uzYzwEhs+s8BbUTge6KPJh/NDqsr6SzSCA+u+MWB/wc8tW4D56fgjRLCCg
X6eHL0qgxAn6+xZnVmdGTBn0si1N+MFuT1yz+Z+jg61jF0E0QMCvgjssjnq6FMz5
JdVexNEfqJpTIRPZw83pNuMjQUQxqWJww4+dmFw2XOSVp0AmJ5R1sP/zZqTEJzWL
1N4aAqhF3AfGbbEDvp2bIhrO4wKq7VZyLOJ4gN/ri35KwS82uZ0QpdPvFMXOKPgA
WOJ+VS6VCIdcApl1Q6mT5IbhiGMhgUiLXqr7X1kj/AI20twgIDeS8pFV3Wm9cidk
+Ybs3Raub4KqLU2QCS/HNTjoK5+3eGUocrdEMoXuPYY3TpsJoRk+fsEHI6+FSyYN
4Cq/e8xC4eDaQmmNLvFd/Tx2x3ltrRxKcI86zJBx7q0e1nenV06EaZDqPvGlO4TM
WjJn+9JwwBQ5qYEunFbhb+CPLLP0MsIWAgB3DsUrPUgAKCoaFUHgkFpHHKNjExdl
NDmksDyUrGwt7gwhY36qHu28CiSa7mYWebad0TivxJUcEeg/Gmkf5f93/QxHnRn0
jLE/M88TFmDV/NfSE7R6O3DTl0K07sfxvpnHmGgquaUvzF/qYySKDXuRKb0yAH7y
JTwQqDzA3V0kOurOrHZzfgW7oerJAeqy+aK2RKprTc2xrFZCtSY7waw7Ho9qSz1G
cbXSSMuLB4BuYX5p+OzmPIONFnhQvTq8VkUW4nV5xNN9OTi2lH3cNBhskmGLPAEw
S6poYbLpCSKf25+C8Jh5r/YFBrcQ4LPIKAEgqaqbAS220KvRW4CCUL6uqntsu7H6
xCLcLgRSElTWkaXIFJhtwQqviydh0iDUtz5g9C3vdQd/FX2PycfH9LLTB14Fa8hm
4Lkq+L5rLV3FoO1TvtZYrnyevKlB5Zdz/rZTaYKmgdDcV5P86PoF5Xfm80T1jRzN
QuyPDH3A3KF8E8UoY+Xb3XcZL7zvsjkSW6OklmBLRSxVP2aLzCaff46f6xqD/P74
KOQHUkEngtEgU8h/oZTG4dLpUnwpxbr64aZPhEIi9vBmCk70Df3gvq1LUaqfMe+c
uMZbieXN07zOKpN6rfdCwmnpgC8S/niHYIziFkWY3Hb7WX+G8IDn6+INeXynSEnU
vWF/RIWcskYN4kNXjBN46+AakK3Hq2OSAa4uM8Yhj2LQirpgAw0qA+RJHWDwj6nR
myi7YYyhMN98qFezE2BoDv8Ydah6pdfZ4RJ8BP+kLISEEUluXSg46NbM49YeJcoJ
esSwSAk1w/20ZBFFcozxzA6O/WmwnGx/2ZgGChsNMhyYrlU7ZGT77oi97B1DMAqx
G/Qfo0WpZkztSPQ684alYjdRgUO9T/ZVzSDcTl0ydr3emrjynkGx819rvcBfv26d
yy77OSDtq4wdszP+hB4boTpGpkCTJnjquTrkIcO4NIFwElSe/FVoZ9NLfn9QSSCm
eAVA6fH2qTeJ76tP+v+Nww4G7vQeVwmPJ23bTeX88tJGLg02/873bqEjr/4530dI
bBQdapVWhWPS24pMjvbnknWRPuIC7e4pOFGGk/LsDb7aEWOk9sJyRMrtUP2aCH+g
dR9CAkxTX8Po318VODBCrHTZ2lHmhy9Spa4mch2Y4XxCBSpmYRzDKORzAPnCFkG7
xO2jSnrPoMNcXfiiPhyNE40DbIwj8hmcSYhji2M0fqxvboegFQwuzB2yjjW6EBTP
MEa6H1X2gTX4phkIS9BAsHKGmuUfE/XHnQHMxENG0PCnR5ZNfmI81ay3z7X9jRhA
z06rqIu/H2Eg9EeiqXp4U61OEyjvFDQcswFpCCHNq2LxQwjH7H8wob/tnpcjQ2Gy
cP08sHzC4sNR7WKSkxDfOHJX/HMqJHA2W1O0UmxaNDWVOGUhyURKRPalFulDYXwn
ReRd7WUDgqobnvznpRHXh38u574R7+6vKUmBu9bodM5/edOYlctrVD2vxbyPhd+o
YAejM3/HAjJ17GiTPmutNUJZY9nm9dlRaD58ftntOM1EP8N5mDSQ1PbNw97eM7mU
2aM4JJKA4sDlH8yJTrazv8cwVAXBfST6V/scRVej1o6849EVvYr8Ec3JxWg9n036
PZNVyPZydKsB47pS7RnCw6mPylLjT82uD1mjyZtsTGHfXWEt9w4fWmv6bmxU/1tT
rfV5JhUKsPxvYPsf25IqiL5+OC5bNn+sN0MbuqtHtAdsbthY3FJ+nJ2hbLceakd/
5u0v9bvFyPivSkaDQmqabX8bJQKuLcYl+QBi39AAYwY/tJp7J+wVcJXpTY4IeH+s
KQpwmELq+7Dzlx1yhNl5Bgi6zewL7cZcchR7VES0gcs3j9kEPlyRM/FJTOEgQytB
pnVFX3/F7NIyFN/i7VUXxWNUlW17IbHY69a98Sj8ik+Njoofe7MBtEjKNytYw9+5
JioRIghOdY8Ud+wdhT1SNb04hhttpM/g92CLd7vqTQl+wuMKxEdw/+8FsTpPVpty
gHIT2682IQ1JC8ULnS8KP7H1nJJ4uNEtC0/vznHaRj/gkNJIqb2pc4SwMPXkIH4h
Uq38wa9tQao9y0WovANeOowAsofkGfpinlt9v1Q1DjLe5tlb0nnrEJWEflNuuv+6
2P4D/dAIk2nurazwSbdX9CuJkew0xQ/aWQ2Hi6RZpazgc8nV/rf9OwWfIIh62zds
TDchbVTs/vaa7N4BavJ1RQwT4sHiKuu5t2b4dcJxCM8EcC6hs9LHxfroBho1Zu5a
jdQy6ml8tJ60RHvwgfSHq9rYHOLc0lED7fR/furXZsU9ZXD7n3l9a8LZLYW6hT6T
NUDKm7UR3DmjD8ADzBHGotfT6rwUiFWydMiRm5eaN/Fe0e9ZHrKz6ZBG+CY54/zn
ZfcfvQdI72+CLxZR6cgwWOt7Lx8G3Xpndt5j7vo7hr0aJdequORdL2YJAsnQ/1TI
S3evhle3j2wIQt1WyWIwQ3td4PM3AXaL7l1+X1yKTC/upQxj9d1RF2Dma4Jvuyoj
0sBVcR9l/xFJ/il6y+5gxfDm0rznh36pDbg/gg3mZprcUrRNeQbNikaM76uLgX/n
LdrDfQIRBLwK3d9Kt+ZmM5TFcnyQTiHvAnoW9xkgElc6sa8IvD1Fh9rjJ+MSxmvW
bQBMLYcX+KvaJNU3mU88cg386xqH4Kkdj1V882WcgRq7Seww2Ri7V2xQv3XucEaF
MLj+ANXcLkbfTcItnHGsDBQBxDxU1S7xBC1Zab45QycKM97m2NN7LNc6Zu7rSAHG
9bh1m7cmPGW4hfYeti6Was99OUg2LQ4Is2T+1Pm9Bj0NRMBzzwBYZPkPRYLUqPKu
1FcKBULnaHkuIV1AlcmHXC9bcGvyZzpDHoal+cr2F/+qAki1kpa4iMGL3Oq7Z5Gl
nsX7v7BF/terTyJtYAOiSeGC9y26CmcOGeYkGQLLe4D+dGYtxKfgWPz0N2XBwv7w
K5/PBlpnKbTzCtMkXqGgZbRcvy4yM1fyuP5Gsn2JTOviA9eYzF+jhIl1oLriZ2zw
kgfHEHZNer+NlurMoo09Ooj8OuRXO3kWpJylJ+IWOvgRGBUHHP9jabW1h86AsAAm
BHZdSnq+WFeAzE3zwHxsVWLAydQbXOYXe49lWUo9PtnJAr6bvaw1U5Ipx1YT61M3
VymAdc7hVx6XhZf9XS5w9CpF8i6YDvCzTWl2H0N7lucYESbAtAKXdIhMh3pxUJlB
ateUl5Wkf4Hs1DwKbpLRLNYausZJG5YxLoM/Hgt92HdQKldEVy+2DwaoW0cEfzP2
lf1ZZ2CHOyqhXp2zxxALgTRY+HoOVWjJPUperL7AxHv8OXLMLLXlck7ljxDxbeYB
68jBIkjmDxQ9J+zLtHpn4aPSs3wGlf/I0tsxlD1b7gIi5op7R5bmm1G8tQpdOrZH
TZjZ51XBpDSBQgZQBcyq1DQd8WDkXiiOrnHUM5tJ9YEooCZ7c+4+n7zq0sJVRuEF
TjoY2LU2NhG5n1yW24/tPbGLfGD+OTPVPa7XcPBUq8CH3TmXrd06jGfxOMHBWUS2
BqH9q1KCBJ9QUh2uQcF9LLqjQr1n/6nTSLnBza3C+5rhsDxyIgYCU8Tyl2BJ8KP0
rTBq/SQHggvQLy8gMmfUboNlRLrvGfCXr+aTr+WBPmej4whGyLN/rAydan/aVcVh
a90UxjIGO+hKlYWMcQvC8PwTddDNJWCQm02Xng6mIPlGgOz3+TGWjmeLjs7KjAaU
4mVkqZ4B2ZPgWEvA43QIGeW1aB2x6JVzFyRUcbL2JUV9Iw2t6aFJcPR3+NElVUAb
FZAtRSrKA+px5sQS17Zx5tSVgVoLOVANt2feAcN84jJzDSoO0biWRcmWbhP8U2TT
VVZSjsmggfNIHXzb5eb3ttlO9DLSYilANIZZVgrFdAweSOyPs7OunsDXnkdhRo7F
GWencOgiIpUWisO47reFkI/O3GUW2y30sEdNIGDP56yzQuDctPHZxCz2mB/EzUJy
PvCNeSf+GgVf7pWy7uikSxoQrJSYJmNwhn+bUobri7+D1ABhm7hGJSzeiwon3qK6
aLQwyj7K5WNAFRRGOLoWJydkCztTKWqp/5aDe/bEQVvTad89w0UCcp+V63CpHl5O
2sCK6Tcr/1MLBWbZ5vfKny4feAYMsuLvT1/EG/gzhpHRvleCQ7QaW1V2v709aacs
dvkc8wSz+gTlodH6aA2yvcjrENK108MmcBFIRp8huzgtbPZicbN2ieLNihTq0cev
cWTOp5hneKVbJ6dzbQHvauN/MDUWTsFZpeNfJ018n2KM2rmhM9R0H1rRDiOms+KG
cOMyDy5IyM3/44vwuK+DPZQrrnHnuOxW+qntco0E3J4137/Wd+RMwJWv6JtYFqj8
V6XDBZqRPkvqFIen0dq3GpH7EFaIPl7y4KfDlIMLk5950mzSAxvmSGwYIY5Vt2Yo
wZdonJvK7niCvKdZde170alCBMxEZQ1GjERaFrJVkdbBvFBPouf4jFkFVwEn6VMX
PU5xBPvO6Dk1btUxnGkd11jpu1aY7V/CM2iRFOnaP8rmTIW73Dmfc7x1GA0pdyMo
G9rY4MUbqciV6EC7yrlFGmlwALI2j11sgSaE32wnzMmw823lsRIoQ3Od/+5P+1Ae
q8JFM8Qs+qmLHVI6qzSJ41yURP2vTUAiSl6hEsmi/YoN4uQroP5Clbw2TMZiW2HU
sriXtRGk4exUxeiuHXZPq7294dA2xsVwFYM7MuOA1ieFL5bAEewFzP55R0V8aUzw
y3hu2L04CHdMKIkZd9IoNY/Ulq09xkpy8zbiHVKUiqLHRUKSdZSquXAkCe9gsDjX
GjLKBly1GbeAyJOVvf6yWTFjVxqQRMjTMDOx1UuKLL8FRousRf3lal/cOxDjT4jC
CTbvhajcawJ/95yuHPUSiaMQ/KiyoEz46ppE/u7BroxFUX0aVbGoBoG5Mk8RcZR5
F+qx1UfTR9irllC7zh0yhxq2rCCf0CAxwuQoCZ/wdnTRtKRV4rWf1ZQgFOzIhLM9
v7UJfSqT92l+LCgKaG/Irk8xCH97riQE2QNZxu/BOV/mNEr+Jz40eXb0N7M7bQ2y
2Ycci/Hflxaadd2Z1lbo5MlUHFe5XCdRhcwSDmC0Is8eSaWvorBSctPuwpmkYFNA
vv199JUC/fJk+IP5D/QYlicPNXValvFobxOUvbhs+q92s7PPTLWih/ncGsQkYn79
6/Sebg+Oe+Ywv7tqOUvq1JM14seSaFqOw4kdng+s/PS+BQsbzI1Bq8ZAhc7CI3WR
kQDiWA9D+DtJzj/rItbRksDULS/0TWm4R1VOdpwQDPYwpJjgjP8UZVocxwt90yQh
JRIJIltELclAezo0tmbg44rdsKXp/noeR/GJpcVh12Eb8yhUYYT6IswoeQiU8F+N
YZrKiwZl+NeElaEivhMMxQ8/urFtipR3FzwTLQaFXkYR/d8vacT4vrBXxH5nzIC+
sXzMpDSaPv3QWTUWEIMCV34yqFwYhwiAEgYqDhlliofcSb1LmFmsQXejVm0CPVME
OhFqGyk6mcLs8jMkCNUhnEEBTnpu5mWpGnzDKxvUOuinaMMlPwdpCJvBl9FUZb8e
gWtXiHsLA5gnbYVURug1DI1RybA9Uk+o4D6FFi96GFLGcUahJ99XfHF5SAcA/3wR
Pg8JyPo2EjzdLHG+q40hLPajWyLemKZze2nv2TPy+o9fEj8tkl1vJZoQu9y5DxQ6
4UCY0zUc5DqY9Giwtiere0DgoTJce22UQWBuiJUjoOPBTpF980Mygprod2ZiLzer
yREMq/x5a1+P1Mk2HTD3FV5Pm7uJb+MKuycGJYqm7kBD2g+dft1K+GK2KVQCVFTL
fOObT63794EfE+T1tfZO6a8L4l8uvh5e4XlOqyyeXbBVTe3YPOPmJvY6F6IxYf5k
mqFm9gZrJ+4Zi09JbSA99oZVGz1iLez+uTr6QVqgr3dqObx9n6kp+iqOIYH/RcCD
0o4muNYTl8Wndz2goA3UnxOU9haKYpb8JuxU8louf862/BB92cAxtR+5sZ/I54kH
WZV10Tona0vHq3r3hlNE+RIyELYNaQdpcoOz79TJu6SZMvTkzMDp9eIe/xQzTQog
YDwFGtGhkxuqcN5tImHTkBVSqxXEA2Eo0PcQhZRJH4uTLm83SI7dNiYhsAuonGEk
Gls8IK+M1QzLcqexHAjWU/6DJIg2GRp25EFHvapsB78w1kfdN4IyJAczVA3l2b+K
JWmr1bHZ+5zP1Zhc/pDofPfpUZEAjFohi4q0bZyJJDA+wcJg+kMyybUZm1A4/REA
b//jhAmeNDqSYq56CS2Xmz8EUEHjvJf9RZFOJV8sVmE+zf3nDgzDegc8U6Cuu6rm
7GqDY5QfjhVx/lMUAZeX0Ubt/OyUagIeSsYrmrYpH7TpMMZzKsFYHvAu5SJ8DrCu
pqTuEvuxDw5f3IjVA2prnfMIQpeHK/JmZw7FYCkSKweM0jwv3pXYYKTJTSMDaTQB
nVEWyUoJCxRPjMkyKF6VJVzBEdfPExrbJAVzSx68FX3IKdVpsVL/AWD1H/voEPJ8
zjtXpSelrhC1o4Z/ikUIwvWIRoUqkfVdXe1ojicFcRmKnDRJ66pNpkTx7m7E/VWx
6rFOTEwwV5n1+oyRzlbnJTJBJv8ODCAkjVDIhLpy55/LZTlne4kVNQNDzrQtRuQn
QHzAUdj0REbum8ikDWy33m7pxJMxDN12CJoPbK+EUYqJkm52Jrr8Y8UgIO+kOJbA
oHhCtN1btFh/fjqaGj90I7Obq6CibjJOHiyzgGrxwwGIbH/z8Vtx2C3oFb/ZQ+Jg
he2Z610h23LFhqg6X0eGhIJCjNSzDnrcnaXPgRr74bh5f3SuiBtMj1cikSsWyI5z
WBtJdES4RrxvBWFUYwyEUslQuB0bXDB95vEJI25TUvwdgsQKb6W+kvPuqZaJLD/q
frTgHL+NZ8RiEk3kSvgd2/+RGgUxNg8XGlRKY2uscLb4jrszg/iksvkw4IQziaU4
lWdX1Rn8TxxzRieaWyYN/YFHSv2auVHw/K+ZgwCZDYWkHq06+rUYHUxRkd+tYdFH
SkjnZnE+WcO9hMLC9rayNH35GT+1s/UInwUbBZWxn6CqvFMtQtfEk3fLqBcjoed1
epj5izXoFJCDJpMpkEdpW5LtGFW/VuNiH8b8rcJGEzNetj8aBo+z7D26UlgQFOez
eNhxTXxT1WNL5nBwefN5jKnw64iBEkaX1uOHM5wft9DysNfmwWrAZtwu0OJJlLip
6iRQXwLYCEJXq6LHj8kkElRKGtJc6Wa7OfKjQu9E4dSKgWrqBocaZxtGVM8wGrDP
lzpY//xArEa7JbzIwaR+oYxkjHkpeSWIbbR288WI14Ab0gg14ncqp5q552YXQ3Bp
A7p+sfGNkFAq2Dx//1V+UkKn2n2smDbhXIa88a6MsIrxuMzMPuURDtY+vdhn96al
PZr8/Wa512H62+9FOyA8/wusFFmvR3VVZjtOwdr8qoJn9Tday3M8qxD/jcQqWQDU
QKT7YaloRwgcT4lJVYLRoPMnJ4QrLcTCJzUn7pTGm34mbUsRpNKbA6rYNRctyqUk
FmMpITQCv2izY9FPNcLsJPsskoQ1UF2RI+kmc9JDE2jf9aP/ZIODY56YZV+fPwOl
RH+pxMX8zTv3jRlKGBUdpWoqZIl3+cTQhEZc5DeenQTeogAP97m1Tc/p8MZZvk0n
0aVSCC7diPWMqx3G1uhMzPOvSKQPxWLlazRvzA2xQ8ETrbAc5kGQXCgT+nVyMOch
XSKd1cRTTWntsukRQsCCq0offezMDkMyttJTr/M++j2yEtIUWUSDAhUNUMRU0fWu
174pvZKv1CSk04QCVvwdBmfWIiEXsEXBoEwlKGmzVuKRaIvKNLcbG6CDplVaMQ/0
eM3JDopbARlBGprd91z7JGAsrQ7MPijA+iWmyLCiYyU5KWVujIjoSSIfMJJFZo8K
gtCLZf+QU+d5YkYyKcdWSshxee6QJKRtNVFmIu4JzY4qChlu0jy2Z4582BVg1vwD
wJOaZ4mZTnXmDYlmStBkzfszPXzWXuyvSMXfzJDkPz33Ei03Prxr8OLqGvnewfIV
D8COU+fPG3zrpSc/uF2wp0jqzm/+0+FBHSxU4yXeTQ71SRMB9MLB0nlm9/wPQbou
TNHrT0NSLiHQ4tw4l4RRpDXbwYMft85bl+lDkM3VVZ5dDb43Xi1aFcQ1Mmiv+Kdp
VrbvG8IVTBNBEswJib0ZEsrUp1tg50dzOG40tV2usgJDOISfrapiuMfnrFOxasmT
F1N58ZAGCVS5jxj45LVYHHQsBDLLz4UZFXhsc4kG9mSlcehRqeYuZEgmN/O+c66z
FC6JRBhqZECEFOfNbXbhKmbBPUPUSdpOK+ffZqJnzWsxY0GuP+uJN/zLQDX4HHmF
XagcE92de3I1mWPbj6WzDbHmjN5Cisft7qgR4erAJoHWqfkU72cMORmtlaa0xRcw
YupDcO7CGs4Phw9isxnTlgM6LB7WIm165bcMo5s19aSvLEMo2vleapSI8sgKcEfl
Kz/hucrEwL4SxmlQIQyPu7R6xGSYeNCmn3tYhcWsocDbq4cgOAXjvCN0Yu64VFpN
e3lfp1NSl4hI4celUZyIq+wCZcPSli90vfBjb6Ove0u0LyluYMdFgO7syTUVJhpd
vtAaAWyARrc0tIczC17jX/L++mlB8zZkE4s2pp5nnFE5ruL4p9Snwu6Hwqhox18S
UhanUMfbpkNHCO6nYMaTyetejSiGnqylFaY3ZXlhjlngVjX9wkZPMqkvRDU6EIXv
UcfujkPZbKa2MhvkK2cMzqEjw0egsKgFLp+jVO0Q7rN4xfT2JitS3WW7MDQYm7vW
LU8Vy4DbDs8WlpY92rP18MBrm/n2k+DATW9uM3jy3NssWdrI9sGJMKeFmsvTg0Oq
FSi3UzZj5FWsbCsuRt6MPQX9uKKAw2+Rm8MtZ7BJ94939m5F3yTWKZ84J8PecT6j
1nlrdonES2CDNq3vQ6uycZyJAnrLRca7iJnMT5pomUBkzJTyNUPjky6FRm9z0767
lBJWHUy23ys7AflU6HA9XWvzAo88y/jYxeqZG3HbtiiCcwjb2y65sQeo83Pq1gsx
/KGeYpLispALyZ7y9ShWCf2rZVqG8Rp4HSQmLLq+h/9ladUdJvt8B8hL3EKR1sVM
P5rNuYIAS31ch2LBXzd/lBoCQvXBQhESp8Mfpn0kejj7BZU0X589Pu4b9JtiTCVv
qfzl0ayar7bnS1bCkIqDlqeZzUeuZukO/lA2yzovLzYvtJDvexwKd55ZOdCxN0Gj
4YYDvb4SBEOxjlefx14/jANk0q1RhY4/lU92R5MCbbOPmlcvpx04BdWCfAnsz1aY
r4aiBGZxEklcRtSrVJ9skiPdvZ/hPwAfeWjPkBfIzok4tihmObIQBVo4fLZPLPmL
XgtCCntQ3XDP/ajqbEgLxI35Ra3Zgs5n2QQ7yG4Kd6AeBO8j7YGPjLTKxgone8sp
MC+ZlYB4ZdnExjkzNEkSmZpBKc+fMo/5M0nVLtkwYzBKBKqwLBYNgwWTq+jCJjUZ
wB2voYAo/NO6FZ9PV0w3VsFe1rh5dB4fdVD8oSSLz1cs4/r5DlC5fRmBUgJpdT4X
Gz8t1Z8DNRgQLJYEpZeZb/+6oWX2QBA6KDpNZrrNXc7G7Q1r7G7QrDQ/Ecc7DEw+
6iQSOjWkSD9+zyi+q0fr4XIdMst//plcqqnB/jWuqRafF13zyjti6Dsmco8TMxj1
H02yS6mpH91CDjDdm8ZnmXCix9qWAJFjEanbP5BwnYmQo+n1+5Bfm05plaqcFwYC
yt8eGfnPNtva0gTXVA8NlWqFyAucX0Y5DOYRE8PzTlwjJD8qSSSlxOEyLDprTfLM
WvYaGf8XJ9FiwM0qg9575q+brx8sMRiZSHjaOaBIyRYQmhecixYpVNdwtv42vbba
juvUA6uXv8PiOvv2KFyK3/SAllnQeXnkGk1YiuvL102mrOOiLjf+fLJEKbl/nq0/
K5j3zMmy4hRN5+GXCBC5zvQH53FK+Vh1UZnp99aBdboVrEWnfh+qZ7DwOpOljCjB
TEVSNRDwUrFtmybNKlZDPyzuOLQiIVnvtr1HvX02n0MhRsdiWqKvvhzZkEx36b7t
0tdrdaWE6yxqrfHHlpD5PGX3s0bIOFMehWIAawr2CJEDKUJI8cY8Unuk2YMarAB3
udvw9mEMHCCvzjaK9mrnuOk57LfVvWQpieIiVzpJD5FSUFHzyB3Cq3sK0lt6Aa3u
QP1RR0Rahn2btXkyMmM4GbdvL3oiSc+HC6a1rUZdZFPPhTcVSklhOksfBbC4RY0W
ZQ0rc9VahbF6rm2O8Mu9od6slAM8nHsTuVFkM8A07mCdijibZGfzFoIioergHSsw
Y/Q48bF3hXM6z3FQvJ2tL/EXvK0kFH9OWY95adqmfX8APf0WpoCh0rh25mgcCIAr
vt2lyvi9VyYZgkTYxCCi9c3XipaQO7S/wB3VVmyL7BihCRtssedsVKY7Z4coc+sM
Xw7HgUd1SxpoWzqLNdADSlIsYBKimnpZWQUYGqkknb1oJBiAG12aKNG6TlQuMU61
HwqBmCTmlleRAdTB0r2Y3PXMNFfl+aurFc2TSEhClcvIW1+xeJIENuBEt4cc/1og
WzOcnyqLcRyoSTMG2WJK2F42Sv6ccaDifljM1bN0aZ4KvJTZ11TpdvUOBR3JjiNC
GnclOc9JJeIhb06qOoOm7tiIZVsLQOIMk5f0hZZfF6mgBHHTjt16ANG6x/mqkmg7
9jN/DqTJHIig8GiL5QqVVwtXp/Q6WwOISOzu+UJae7rPiJ76TE1A6/Sq8vOPNM5W
1L/oiCai3fv7Jx51KzAOT0RWMhSQ0v4bJ/VGhYx9YxgKmcN6GCVOyEyrJOCVMcgZ
XyhXr2q9Fw0nXmUjmZqmreYs7tFXc4XYW++URRqNEGaryjOwJsjqlh3T3B+o27VK
y23uF+MRzTZCrcOUJep8wBFrS1cPWOEbz5wRX0tEej6z3Ldby1G93YCyrqi20LWn
jktuYXE1xrLlaBbYbLcDOTKiDIaighmL+t91GOsqU+6fBYK+ttNtTDthpbP9tpem
P1ig4tevPKtfl2OIbQa2IIEivtkgVJEwqdinfGF4j+bqqiG7+Dj+D6wwAjE0/GS9
8J6Uwy86PmzaaDOfT9dERBBogUZ/aPxVJk620wd2HipOrdhe7cAFFNgKgBWuDLN4
XaOO3rixd+ZHlzc5BIjqarTjQoXcO8q3/eKYhZ658XSjuejHkwcGLYAVHZ396KU2
0iJL8klicewBEF1gAYOOMJ53Nup/xm98nNW7KB7o/qWs6GY9kbIS7EN6kzNLThuL
B8bZsC20GC7drAH5+tozfev+v5EI5QxOtxJkBL8z3TQzdfiTeGTNHhDF9mEFN4fX
8OWPTxAkjetnLozQaniOWVK1mIfMvNcWUQcwey5eiobfF5IRW1RGRXl1rLb6DaB0
webd83bEt6Vz3S4FTZRfqvgplSUFypNxZebFvKfq9XlomF7XL/CYWJGzXTuPax2k
bMP2OjT1iatxrhpc7ua5ugCQvzhxHouX7pdGzXJji+YtSuXxTaEW5jHygqezuIEn
uwwX7DeF1h06mOyDswImJ3adPdZkiiQpzz37mEDifI7b1q/PhIRR6M3EEyfpnx5h
FjZ9eBTKyZJDZalYuajGwrA6enBmtjV8+uHhro8frx487ar5a3rDUChDdZquVA4T
+2yq1heVdGgiv+kTTyde/8UG9a2wVijRXk5lifwNs3MORcXWPY0KKbKRLloenAk8
Glo/cmGzuCUCY1cQ7NIsn2K+L2b6yg8rXr+De5KindnDGot7KC6dcl3e43We218W
qfJdhG/Wyv4/ShjxQe+GYHk7DkPaq9Qtuh3vUUsjZXsmYeksVxTzqR6irj9Kbq8L
oU0EQ/164Es3D8mvir5zvVKhX3DnRa4KlsfZGvr2s29LMYwgZf5Oz1T/eTVUjYBN
NDSVhW4l+I39nI994PMP0RZ0alKMcvOJmPY9N8s3eOKeqnIL3dpjf5BicytYlHxf
fYLX8a+XPhMC/pyd4jCUk9wm1G1F7gQDtCmzKY8gbtTgM7mwS8DT3IXLNKBKS5BL
ozKMu3SdC////EfTY/QZaWp2XJEKjbxDFu17+xp04UN2pmZnbQLu7WgYkMaTfzHV
2lDfp8HSle3h6JmjMA3peZ8eP2hImns3cuLsHwrHJPpZRx1Q2qYzxcCRcdMOPNRX
yfIA3UeChSjBmyMISvsqhR65Dn+sNmJJlt7bZj0ay264d2PKj2BBDLFiZq9Bk9vL
k/L+Opj7MafLIj+Q6cLuxiLIvsDlkSSIY4XJCvgmC9qHiPUDFsrmPnRF5PSCZqpz
ZxFZs3OcYZNVg7Gw+7HHpvXaG1YwvmaS+1GzSI108b54+G7fRZz4LMnCCTdQ7A7p
6OFQ1tbSlf3MOO9Yg9EFhffvJrSy0bwgVNjsGafrWXABRC7rNVh3orSFLzJoUfIw
mN+DLm5ILgFOZd+AwodoeeX78dxu1nIkbBD78yefki/L06KnNe/kIAHqguKNDcxH
alPClNyYC6IHkYZgXG+0q3BGrwXB0mMjW2i0139BRKhrSywnOT+EuAeTEbmNfO1h
YWh/IoAz2zJArTTgD94tAJF4oXqDjdOFwgtfOu+F9lCibihplLfvoHvG2gCFh4jL
kf/XL2JpwdOjHyE2RsSlwohciqf19/z+X+USeY8+XPBY5cspMcFShvhSVxR8ufiy
rAnQJJlAkvG25iWDTot4tqy92/4T3DAL3D0FQBhWBnqTSLnJXa4/RCc/64EdBZME
KcJheqx5oFGT+vUzwyBCER4JqlMXxAhiIg5fVS2RFh7Y/z6jmKsqbrFsiD68eH64
N25xh0PVvUNbAdlok282VWS9N9YZmL5xBgRQGnDooyJN2fzzp+su6PXRRkd6FIXl
xm2ViGaKS6JPKzDVSve+X8SR0s1o6fsP+lTMj1gmLcIWLnZ2UOoTer9AbYbBUaYl
3Ew2cArYjBSC/14qAXuEzDcWtlOFYwvXqFsz/GmNMqVqgNUG4nRpckEheXDME+zN
U2AoUJnRg1rdi3HmVH0gSfRL4Qj6KMh4AwAnmv8WrPtx9GxXH1rzR6JwVR/3+S6Q
3XpPd3odP3Wg5jslCp2Lo2gfeMXjuFb5M/baSWiydkou7SbiN/2uZOS71ZCdk6rp
AXo6r1mrqutALu+scqUHJLk/vO2MJmFPZ05taxKaqf2l2O3cmCtRjC1o1aFyWWWc
ZpoIiR56NmWcARaQ8c82PSKtCJI5I8E4RNNWZPHTNwCRzLY3JXW0CjuSXw+dDzDI
2m3m3llLgUdl648Fv4GgErjfkmZHSbljzTTI5dsoQGTyovbMryIx+NsrRpzcBIC5
t+oUtdk1qRWpSu3EaFk99/i39ABj8ESMVSvl55/PHnanet5a4L/6ocfIb5CCI4QO
6E1tVPLnwymkIhpihRHpGD8vhG9NpUT1oXUgyDtZVATh4Yqqusxt1ncamdCjIm0q
brNBD2HzlP+P/Cf1McAcqDyxZE1IluXOPeAO+OFnh/bhLIHSc1F0y/S2+PhQIDq0
R+7Tol8eLTg+WbSrQnZacOsOcGhrm+QMdOuATCX3vXUsOmyDz3I8kWtq1UIGk73S
FZvtLD38qu37itrDEM8FL/YQQBe8Ks/NtK1KEwIx5bjRBG+0tMQi5MU3pUeU5BHY
TAvDWm1BFm/qRkkkJmSBBWjA9JRzl+vYwoPmGVflWAKCX6WQJyYkmgSlFT3hIbdA
GcaRw2t8ehLpC30ElIs6eb21lB4YOjXfV3DicuwPLxzRtULmOwIx//EnogWb7HqJ
g9mqD9XD7BXAbsNNlAqpmLa36daFd0KiYClD0g9/f5PdGtx6hIIW5v7hxq8/EGyS
n7TS2mCxKpsY9iRhQo17aoAkESX46elJxRdI0lH15Pirgq75T/KG49NWXzTKjy3s
El+oNVonVVLrDo2HT5t6X9qvAjDBAVNZfqw5SlPERTw5S6MYkk9gziOEYuyofkX2
WszcoFN3uNi5EBpS8s8/xwujVAwC16dn4ckfMO+zrdzqucq2YIp5wz7vhIS54qgL
C0ybuy8E6mLX4KQHnt9zZlTKySlfhu/Ec6FzunIYO64kg+rDU7anpe3pRvCooqjh
4BaMUQr72f66lIqsNPh+r+8tqNdW2XOA889R5yElr/0h5GmjS04RfYMNb7CoWZKQ
UeAtBOY+YHHlQ7SOBCBt19zuWbGepbEAQzO1NS6ilGLagv+236sKQJ1Efs4J/FVa
A5oT4gvh6m+ZqBE2hJqiIRrxH1qq2wWPD7UgHExb4ej+PblC9TIZtmCHr3eYBG5b
fTxbdLAlEju63KdpgMJcXeySljayn8mLo6jBreUtUQ1ZBU3Q+wY26prGXNfJB5Z4
WfYHu3RDRGXHSBlyTQT6EU40aZoAWsslvNRfsN7xKq+pDvPN1Dbjk52hRopZ6RRn
52e5LKWwkrBUrN8bgCLT8fnbCgP80WohsgSdBstxeVOzWqCqdvFLWijLjAsZ/UjY
Yg040oHndVd4hQ79p4oCdbDyxoshbqndF2ksdQyirlwx9QJCX5Ay14u2I7qBOEEo
Li08zhYb35zKU8h+QhC+BhoknTlsf409EW1tTq88t2DN6modUijCBnpkL1V2rCIl
wGY/njeLro84diRbT4VVS5tifJDWhSSCawHygUaZoGjpoOdRYg+PORV8bqMBQO18
rthfCJ55gPxrfOPIGk3cDHF0W5j28cUxHcjfCQYBePPK4NcZrEDXjwfdWDWciHgD
aEKc4MwNcpurQ8+M+iUswEOy5qvEtNg6zO49faaJ++7Hy/SnHqCXnQFjoUse/8bg
yTuYH1CYlE7XfwjQGBSzI4Ngmox/4WslBtVWpdKjDd1jHN52Hdpx0kSc6BxKozAW
efMHJrVbYrcZysdYporZhtOgi5oVLjdrabHvy0HXGBFRTAQyYx9cKBH3qqVFGrtu
m8XRxacIELiOUJa30DkytQS7UUi0CQKAy0gFhaA4Z4wH7V1FBqSJ+ZLT8N/8lxSL
wsYhgyoIqdXEZfPmIQhoI6zLmwKUDGYcle990X2KCHhdVj+K2iuLVtxvPjHr/wn0
eF5FB3h3xd17msIpNsdq7bSEo9RuyLr+sj2fjXAvm4P6UvWWfJQwrXZ2N2EUrsZG
gyeE7Oh7666hMtuyNiGTp6pvAMZEpUkoLC13ehdG1P9YSPbKUyf3r8K3ocuiuPAv
isF259RAjbUuX+x9Y7rNsvYBHF3FT5umKUcqN5lrg4+FM7kIUFA2sZBVdwlFgrSC
0y/rTHCwh9+piblHgBJ6eN19NObq3ZbjwOnqHdS1RLZ9ggexY/X1ZK5HxysWAVqK
wZEdAQT3CD85x4rWlfa8I+hvmLiuW1C50NDv9PI1Um9qTmJjJrYQALUyVL2wgkQY
dDk4mWrCcYXVoWFUniEvsAKyUuQwAesb1fL/cjXRsFXLM3FxcGnLw2q0qtUiC5yG
GuYWefotlZAEywxdGUVZZShcBL+BeW8XFLYU0bIor7QAaokINq7ea/bstpfEqavG
5hIYRD4rXQwyjPgUFmtLpg21axbD2CJf0LIElykan5nr1EuIi0Jbmkhe+7F37CTK
MetyJats5S63dqXFZ3plxopJOd+k5iAl8/Fc2oAS0N4leqaI6jnb20Xh77SAh/Vz
Tihzr0sPX1wXFjc3qSRWFrJb2115uDXAdrqDj+N8BoL078NFzx1ItD7C5DAvFvPB
KxMt6VHLa8k/nZ1mT4aE2VUKdcNpoqYQbJBiY1qZjdYRClAjIwpgGKmK6Q2KMuKw
JrMP1B2whdzrU7lZyPJTRDSn180O01m3ypjfuT0k2gxSoya9RT1BANCB5QDY8dra
VdmmVxzczHuTV77ZQm2nT48lQ4mxic9FraR2+rTVASzEhj/PjxcgRoKlk8o1H2K+
emgi1BlP8i1DoR7SpamkLcGEmdgdMylOY6aVyFrHJpisg0mYdHv0Jq3djtrcuAMD
6/2B6hapPGrV+DHxFLHmI9EPSvFiJUREeuK+XLNeKfckXgEejL97JrhIic7m5QR6
/F6cazOY8E2VtObqnQsZph6pZnbEKFObjkBqD2p92dWEXZwYMDpWCvEZLRy678DH
FVAxAb5Eg4KYuSyp7+QaBaA2sHGvaP6NC+4D/GTEvaPsq4/Z5x1Q09jXTcpTXdF7
AAxL2P7l2WmWu/2bU2qoHfVn5H0ANYWO3nU+nKr3QkQzGaJVSNkdHEpuWaf7Dl78
vDjoXebHV3OfS6+cufv14derpSonCimThS9invs32goi0mMAmsahJ9twZYVicsvQ
REPkKnXzZWLmuGROwB6CxI4tjQDlR1jgh3vt9d518lPVpCLbxVX2svhIvTWFU2fO
+DafxRYlAeS/oqu6W+nT8fjnQncvoUzW1ygKdoxiGYJUeusiI+ZfJTXLggCZlj1a
0ezvG7SCr3DXZMS+sTpfl+tiJvdizevobqbN/Q2zCIDYWFXCHYp/dKAkzG/6aWuR
CcZySLw6BWJcSuxfMWstVySazgBWJwpvqhQWuJQjG314QTk7SMI/K/pRaonf4sQI
nhtntHvoYkDBUvQcX0UAARMVtoM3RYCqirQAKR0qlMrTZaNWYzbzG0z3yVcQgqQ+
4svbGpBgpM4loYcUadi34YkgKq+lrkdpCJdHIb+qM/w0Jbf25NrPOm40oQQ93p4T
C3bz7X6caNLM35lxHiFUj9jbSoZ1+FWnT3q171ccXw/dRSqfvZi6i2uYPA5YJb2C
xuk0/eQwNqhB6PmWsbj93RBMoaN95n5ZQ92cdAwfG/UAss3f4GB6QwpWZMH2Irnw
5VkTRzquw8ZHGmp2I0mx6dM6EFTRcD5O65TYNmg5kQUVWece5nP/XF7dZFSLLWRK
3ICi9WLtPp3EFgEP+cokw1drEta6YQ1ImkPsx/z2jVIOX7/SbsPeOhKVIBRJSfbg
yygb0HsGzQ4Q1c9I0eQtYBJqwb+8/XKGQVqNUfPLdTvX7PWC8dEvTg2cv4JWjXPl
DLyuwNQ7pGBWDKj1FRFIXCfXbJ3AS9+WDP9ur0e1+1aeYBpXkz6efAKwJRa5Gaht
z18iD/tVrLFo96r9iqZpg/5EpUlD3lraq6Ygn3c96ULQUsar4Ilnduiu8MAidxyV
ng2NJdHxcEan8qRCDjLPOg1tz+wINalS6NqgJigRTybnRRwFCrY6mjWA81G3zZKA
uda06hdK+JFhpzsqAIvTK4JtPM/YTK7Je+O+/DK/UI2cCoqCucF/s5LSzvlugM9R
LQHhh9g5ok7BnPsC885aZEQXpfiOh/ifHMtApBfswljCSoMWCGG1REHOu7ctbnav
cSOR8WtTbd2T5O68xEY5xJuerFYd+WVcffpcUDnsMD9dBoXzBswfx43rlQC2JWqm
ERlNFuoQYXk560hPydg7YEWoAlYWg1eBxgsPn/LamwaThp3umxsm8/DLOJ0W/u0n
tjwXUlBWZRJsYtj/ZGgVvPcQxLr61FXEv35AK49GN6lRwnv84lmiJSpbgw2atHKs
33BL9IWuG5X+JHl+51wZJOvCXKDnuqld/OC6fgjdTKFZTCb2TRn5DKglBKJ1Lnix
B7jQSe1EkFpNLNkexAVQTDgzjZflkhPlb0nXN/GIYjL52FlgGeturvAdzKTKj1KJ
UlDWnt2TRbU1j460ivWp9XSLue1YkLEkBRWTh4lQ6Qh7CciBwNDovmaMzsClTQ22
+HgHLkjC0FvkfnW0xbSCJJnZoj9W3meGH8JxwJOQUSFe/WSzN5shajVCHVWQDFRZ
icbrDTUa9TViMeuxGzX+en1mA1BnZVcR70D1XVoUPQOhKDCfP1UTRKh1auJ5uzqs
GN38S2a9QOaoTcXQcErC67fOustZkAVVUKckcVkO/cLlc0C5ZTiKCqFwGYg0AHJh
OZa/0HNHYXguF5V3gMhxn4n3TQnnDSNI3WLeCsks45BMPbo1blmZy/v7UtQkTg8f
kB3NtEoebTwIry4wo9df0FH6OBfN9QLA1UbdJ8e212CrkfSlX3Zwwa5D7/jiq5II
IzyXUDOA5Bxlrz1MaQlFGjN6li/ewTzXjk0c2qL/h/CoxIMdqVNB8eZ7flfyi74C
XAITMJk0VmF9kWU8JsFSWNkmHjxNWhxa5UhlBUwZZFSxyobLEsvXLrYDw/2A+SCF
Ud8T7TUFqOYTPTHlu8+13y6X9xRGyQ7atjEREzI4j14lj7cHScjxxZ8DzrPpxG4m
+ptYNkVMLUWzut3gatbgE42SWVrQ4pgxr6oUvOZ2p8Wzp6PCWFhr9b9wCM+KiWp1
SaNYN1RQWnaMZ8/F/gLFuCQc642CS5P89JEBzB8YlvG67ttYiLVd5r+irWQsZEjM
BZoUyT6A9dvhNudNnxAl+tl+dvY+crnipLOy+ryfbbUj2LN3XfVVdNJPcgUGeB/R
QF/xDiBBdAbhbfSOQ28WAZWCOYgQo/RlDzAnFzE+o8fzsu+j5K2sSkjg7+oHVshc
k+R343xrdBRN8sXPY/OVhaD6G8O8CMlfjYtg5HwaeOdvbTauH6toZRrNH98+H/kP
Wgvssybb5Pshb6gzHa3eXd+HgawG37hFXIwJUvwRVDaViiCQFaMhzZkBWJNhUCnL
em4UExiQuZY+tuuZ13nh7mcktRL+PHmAGS1WDYaiShe6pB+k8C0Ml32IJT+RG2uu
tWHTzdnvaUgUA3VnWBEArG7Uh6d3/lcMC9JvFb0AewnLBbIPVgaX/246fvBA9uu3
U265iUEauqMNavNtpGbVQ1NNLXIAhaF4E7M5pcvaV24U1xWUBexdovZGOx4cyiN9
aTS8dM1YmuUtHG9KAH3HrziQ8dKuOc3Qg07e+sa5im48O/kJu++USsorr0jsZJwR
VBo2j3f6ByOVpbwdgzGVsIBNoVrk1LWMoq4jrEbIAAucALAVjBf1Bnk+6dXeLbfy
t3BzyOJz8hKupzObG0Dw1RVE/48cpqY6GHrqb56LrHiNW5MhAdjLECeka3hZMyV8
OWyNkkGKMCA08YMqAHx8QXAqPzSHUf2o1yMhewozdw8HFSQudfev3dpGfWR9QaPf
D/w9YxgaTPfEV3t0YOP3OML3Jez5OHrXVy0GkXI0Hmsmi/1sFhVEVsf+byCmFUTN
EfcwxznaIR8Ky0pkxrUUEWwAfaMXkWzoMFQyVLeQlkGHtCbXbM4YXCgjT78HYilW
9mQmwm10f+UD5MdJw7GtRR4MrP34j7ypeiSW1jT6zFuyaCzoITdC2pr8EDS9NCkc
HWH0Db5jScnWFqLwz6fvf+M61VZMvkOP7c9C+3V1nqGMn0FQtwXedUtT5WJAyI4O
/Q4cvHrvbO9vt2Eb+CU/Qr6KILXm6EiwEqA+hPmg02vL+iEVLbAfYE2eM1X8IfMC
z8g/tAcbm+BQnuXkCeOoKQU4FMXEPyg1/iZTUYCQYaTJXjXVc4XIZmI2JxR7495O
pJB37m/zrnsFoblUEUTUi83qoHPK0rV3jkDyyITkNRKv5ituycLQJqS0sEKG6VIu
zG+omeuKa4YRPhXMbtnw2BUDbZo8zL9az7Yvmy4mmjddFTZjb17ZjlSK3eCPLJyI
GBZhEYGiTsDSk3hnd3aBN9h7fWgATIi6LFwsKWiWx4jI6zjcHrX9RvJ+1MTjlUnD
0O0/4d9ar/Hj46TwO16SeSLcuxwZctiGkJ3kzWqhJyET6rgft5VDOMbF6BufUEov
FIm1Q8vVOQ7Fb1p61nspLNjsIHKFUA7LNAub3gtzYUHJbXqG+pzdYOGk9qpg948J
iQTE4BHDBeNUE6109k2p3gM0UX1jj0UJo00FKkHC4/rD3FMdaU2S4ZRtklHpQRcW
rP0HP6hiX8r0s4eie0LfAvHRQkwcKP2c1P9oa1v/Glj56kg+im2ppuQl10KEkou9
dgYHo0G+jH1rj/qgpAfaNb3AcK282uirlPAFqv+jtOzhNGUoHCzyRl2XcH6KF618
Ugwp1Lot+DOkdoUnVLYnZ+r27MxbnoEJf47OGb+JaB4dCpHi0d+8qy1ZBAsqyBSW
joM7XFe49ZsYEXiWKB0uRuHj+Oj74MIMsEEaHgfKmC60d+yFsFNLPQmdODlwd+3J
ljAWSgeeEXjbfz0hPeNW+PR5kugazsAwjmCmsLLHVe1YXS4sIMLxJEHBwXNmAOH6
yKBXu0EtcbtNdHqBzwKoDXAt72K7DsH8yjZv32HXsj0JqNBZ89NDvEpqPq2Mwvn8
gnM1HGmNPrq7Uhe82ZxNyl2h5AhtCCtL9izr2E4s3tLohv3tXpYCffCstFXR6Lgy
9WI9j8LXb5BvgNl0GxGwFdxZ9degv/cVW9B9goYIbv6gFk8MaXx+4xYs0rg4CvX4
IBgn6sutDsfERQGCYNwZWlefZH0jpqLLpkJyeGgr2pyKEiAHA/1mWYVpwmIcqpgQ
js323BYha++LCazN10DaYDj2gP6olrpdKSBZHYCfuGOOHabvUzdkhGoZyzn9Ast/
e2Gw86xrAAKFN9mZCbIjsp6XyaiL2dOqfjZRyxHKO2hGhtH5trkEqWbWABTqGTbe
crie2G0g/fArDVVitB51OAXbxFK9bYqxppIuHXaAdd2HFox8bPAgyU8Tw/e18gVD
yLJF1ceOL7Rd7HzcuWFLZxJ3gDsZnmiijaRH14VEu4noKZKxzyn3dQqC61qPsMQD
+R/v44tdXWE3jZ2tmlV9DCwbgox5cupjueMKOAWAV5/juoQc378XpWS1Cup0AkWC
+ov7cajbeRc7HUSL8ykHma+XlIWWtp9bpVUXhPZcuTuPTzqZLa2vG5RHnZ51HH4r
yXs1B/rgx5YWpKmlBJCaLtH6bFpM6Zitpoim6j+fhx5wyFmhFVwjOtlSe+538rFg
qCBB4Ib0KqMAAceznc2bLIvd5lA4lWnVw7mUM+cct4134fVd8uGtHFioqONssB7f
M+6j5yIVfCL3y6Djj0ffMWz73CxnfHsipMRj84g4Q1L529cHo64oYfLAU9d5MLG5
Bsc+VZ/bCvFAxZEKNSrhccRYjEZ+0o/GvRO7KCHgC1pfpWd+Qf2EIwPr+SgPTyBu
40NebGHE7mqnZL+Lp4dRClGJNe/TjOBzcSdEqhh6zULERFNd/Rk7zaxa2sJy2he4
IQCy7XUXWAk31/lCcUiFUU2MULBCwZTEMuRbmF4lIAkzSmT5zLnsYPqleU9hldUP
zP9kIg44hBYoVRlK9e3R+d9VmsjDX4ryphpEf7TeXlMEl8QwAxwSoMUO06qW0RQ2
KTCgiTp0PU9Qp1+qNQg5spIXKpbkCEqJlzSUz/vWw0d2vOdu0umx+EjwjcxQlIKp
4wIcvYuG0hyzh3MKVRglJ8N9C+kmYe8AcRDZ258H1+fpO8+ypxZAfUZdWKMtUX+z
8h4miz5UY6ZwmWl/EuNF5ywX3yyLDt9Ha61DQ5dUZ1CsnGXuLbab/5PXq7+jTfSn
zOxSOz5wRHuPm1QQe2gMkYd6pSvb/3XxTeRQP+FPeT9+6FX/+u+YRJkeOM3xxIWD
LZ+teSM5B+iB3eYxAZQow5MVc2rP++tZHxtsWqXnGMOjpeMqQOzH8aJrW2u48ViY
kgCzRCvx5oF9gNBqxipIbv/AcRuw/4GX+AGWif7+DNGprUdsKe2t/9wLEH+PG2gW
esbQC6vCn9kODrU3Y/+HHWTQVKMMicVdDn5/lRBUmBmeu4CgwlYLXH/KC5upNRkI
M8uanTucXrFvyVrdrPxZH95e8Z7h9JceFQ2l3zY1zYkugbFM5wOPAgHPyQJyjvKX
5we3O9X4/o1k0uOkd13eSJHR5QaAcyY+G3ITMaiN4Y041xtldEvkSlHpfVhxLmGy
ouhH5jjMlJsg7Oa2N2JRbEkwnD93DGAP0K+OnQeKUpkoRiDWGbsaxFlugWha6COC
gFrNFLtWUUZa+SMOQFHkzhvMzx+hqmEZ/gO1/iF6XiXNkIlkc/xVWsom2GuGMQ8g
J3p/73nwuTwE3B0T+2yzmURd7rBTiAP7TMdF08KUnoaU25/kWF0DlooVTVSYd6zi
ZP99YQ1Sxd1LmeKf62bJeLofSQnMYveE5ZApiR5wrA/TfIaRu6yl21dhwWXAMelw
zKEpQFziSDj1jzMeTNIIQYjRE9udlzLZ9mF88Q2khdus9KjZZOPEwNrxq+YqN+dA
7HaRmp0+FEHGRKbsxX5lbE5uDeH1V1KAMhdFCwmVlBzYVzsdxzSl3Ehd7Q+sgYo9
q19Zc9cRza3SUvtPXR/9v0XM1OW0pTgHNN+/glJUV5oOZBgcRWPbCh/cZ6Ts4jjS
doH89Ka3uHCGfoYLqJzUO1NHzC27TSSVXd4p3IwOuii4+KF0c/SjHAU3llhx7zJh
1zrut37aqWPPsC0pnzmQ3pFH2KDHXLqcr0tX35RK2IdAY2QwTjlNqlBJ2pbET9sf
ab/PNVX1aUTOWMz3c+vSVYr5W5BdUXd4z/3aXLuJwHWEXVHPLRksLwT/FTei+aJe
eCDNiCLy9FP/VjScLgtGkxaEl4w2g0VKUkHAqmknfkOjq/O9suUAwPRHUm7+s3MQ
AVpucg291UGMPV/PXZOZa8LzOkyTZYtdiIeQ4e/uP61lFgNCCRcFtItU4HmocenE
NFBAXo8octhkJtGyevlJj8OXhKMMjmxbYG0ChJF4iMDfcr6+Imi2OgrvOfVFWYJs
RIEIpqpOFLjq6NuGrdLiSsSmVgqHXC5Vzil/y1qLnpWcvbL2iuThqisP5Bq92kq9
94FYNICB56QOJzKWul2/IJC8aXpWuf9Wfx0oNdOxS7JuRHFJLQvQbH77B3fb/njW
u2tQ6/12qJw6zr3k6WDxYWM5qImXjnUgul501vyb8x6RnqEWeP26Tx6buXk11766
Wse3VtomBzHd75p2baSnKFBI4SQ3ItomxOcZweRsRlUD92bPI9nz5wOa2KSumwEt
EEtmNJEgmFYjHeOaSss0poovy2Xd/sfcJCukkBUXUoAKN3PJjplyBU2UYQphN2OW
p9LRB89+qpETRiPiZ/ngSmTSKyYnf/mOLPE1+MNxCeBUgod8SuvyJUTnK1dc9Hw8
RL265vKoY8GpzKUSaHnuc1Y5mfSsvfiokF7D0eIcmj8NfzIIrot79K8ptpkKXQuX
CBi4/OVGRieTxL0xP0AZhpbOeebn82HkesCbxcCvBmLYkYkWstkhGCs5Xn/Lc1T4
0B6jvkqRy+URjOOvnL6vcj3rhSc929oxZ+r+EzlmXPE1Dx43TyMib1IFMKp4TkW+
kx3EyVdxsj3aqMNvt0GvKlnbAyBY+g3XJWrDUNmlu7V+MKO9LCs2qM3DpUAwlyWQ
Mt7rgXgZ1nXv0wE+xfbMMXaibcOci4QuyTHKamvem6eUk/SfKWlL2CbJsZ6YSOPF
IxOe946xLkISGfhV3ZRrN22XKIJxhMCK2MpxByCvP3ZOusvFnMoCBeucEh7r2xSk
D4CMI4dTsKiOWm+UYO16VnhxlniaObyPqcRxKrTqTBFZoVpqMLQYvx7prvrFgh+B
DOrBaDE0U50lgKFlul3l2cxATC7TMHX8eYmm2T/L7UxqMID3OUFPvF1f/t3eE6aB
7XhkigcXU1Rk32DynNu91ffbxxIByIS9vmfgt0zXK1lE2YZ7/yHbDhMwK63C+l6h
ImtWe+fG4BYiuzn9IIphrp6h1IeupKbTnMns7Q5e0zXN9kZS4oTRYSJRmTPAMjoK
+TJKU2UNcAA8sLTIw5H3r5gAWE/sfoKUNA/JgR9wjNCyGiDaSDnkrrobbBaM+W/X
hujjBO+LtbnE9pkkCdU04JGFfSrQyyJXa2/WNC/JBWPP1cZstcO5E8JL1nM6Fskj
SEqJuaJK5yLSUuwt/0YX1zWXWcd6UDP/PRhwisCury7GeKfhoJFYfJcE1iAxYO8B
ELInCTsRBtwaH0fdFGPWFN2US04yBDsxPIAuT0SIgLaZ0wb0/aIeIcZznR+r1jLT
6pnc3+83+yKfMTnVGRTdBYxF6NrvJ5Re/awC0FT7tmW7Wx0qNyv0qLFu8S5VyCjj
ZD1BAsIgwG6RsI6RgOUVkIiJ275xdyxytA7xhB4ZphYCoZzuZA6Aianstc1wpte+
bQplKtYdXLeEJPpbn05YY3dCk6jPbxKmF2HY5BKRg1Te48izIFzEu6h8GAGkliPe
wjMGnO1na5m+bP0HC8uvonMtysAJbLyHVYKMTsIxQEkUPhRKtSxZDrqOvLlfARce
j/Sg0sY0/vj+WzBSX+VKut8B6W7IdVH9w3/MfB37SubLdRW4G3eAQp8pVI0BaTIr
JJ132EhnoYzMX+MCosonP4M5b+GZJPZI6sheDzi0rc6semUkDAAN7pAOUsmsGsA/
PclQQ9HmNFDpXj1/x9Offv62Lk3hPREiipFNSJAh1978RQ5u6ajtIN5XI8Jvp0cA
tNPJSXQzIHLIAQvH6qT34YH+wMMDuJjXMQD7D8q31iwBTJ8BmtcsNDiIS/Sb/KW5
1z8PBcN24OjzC9l17N9cBBqQtW+Jq87MiRREQdmSZcmyC7zGAVnglD6ZtZI+Exd9
xOmdSxgWgLfqHtPvdLuFYsgIJpOzlOOLzhzHTc75YwMR2kIbIivD+57avHegTL3+
txXWsxr88VDX/Wu2w8/y/5h3IgDq1op4c6uZ3v7dDHnLh+JJ3RXhBz8K44iPg/8Z
zHy9m1PqwIkfndOSxAf1PL1NcFZ/CCPUxPdO5e/TDE1UlE0OkZzj08wfAM8sFZTj
7ExKK6MD0t3kQYwX+4q6/8U7IysuExadTu/pG5jT+wO8A8Av1kNLZJnAtDH/5X/Z
eLImypIkVA1wHxmfvnROl0oXIjn3Z6cdXfKHx9j09KOGva2/PjPPWm83HpLiWmEO
okueQFUI7S5vqcmZnPD4sERQ1P+TIfgk+OF74wTQhmlAOAif7Csz9FDKW9jwd+Ss
HC8ZmGYSzH4Oj4xKtDTjZV5B3j6qFc6qCub9Mg1DpwNP9bdc/UiSTyIt3CHg4ICx
7TsXy5L+JmYECMP4dPsq9hP96xwvy4fpV69v9uIztssBDdEg2dcTOIbyp8iHrs1+
o79Jjw4tExJEDQmV+BsJUpmxLARJn3aB32SHR+5AB3yC542uJjC8ILAqxlrDoRv/
OnJr8aY6uXTKNk3JzKUfi1jwoTZsczjjKBpa97Ug2UDgi72IOaKbnP5XEgkFL19V
xoNFvGz9Sf45BmwhvmPJ12nt3HJOPfOYb1bfvonzcZxXAsmzGSwGufgDO58veha2
Y/cwdU6AefxI/67Lls1XyR9v15V1fdc/wehbDLLGDVL+QZZSX7UXw02OPgimMW3l
YV20iLkC0f2hzu1rMHLbgD3Rm7abRE2rWVzBbrL+UDW6+OAr1QSzNGcCFraZja1P
H4D4FJ73YYNRq//bS4iyHziT5iPYIJmyUyhYgR1e3TLWHi3USWYNLt0hTlaSO1Yy
LGztZAfenz4ugMr/RTAEjrXZSjUFrCKvrA2441BIRmWDHR5eFIcO8MsezLKsdh7t
MKGnIOThTlbZnhCAiD/TMlXiEfEkpAc3GEUhbXrFpYrbLcPbBC3a2HwT6Pm1Qzqa
P/MWP08iQ/2SJ1VXG8FkYdRtINcBHkk4aC8WB4zPTPRzpsu2DT/sfrvnqIlVrH0m
YzHINb5ruPG1IIos1tbqh83OGOS/H8KZswRiAY1FSEUah18NdCUtdhHT++b10CYH
ixUrhrx3efa60kugh/4xnlHNXPcS7w+yhUSOjhz91gkv5axzpHuUDo/wU6Osmgxl
X508CKpOCuTFUm3KGsU/NNt8g0/WRGJ/TYCX511mIxBYiiXOkvsQa6RJ6oYM+lg9
y45P0XIti2l3/60cWr6wR+8dI/gLofYNyrhaPsOx90FGUoKpy61g+5vvO6EctRk5
rx+yCZc35enyFrQiT5sllMBUZibhCatFJcagNp2KmIHtvECVekPv5LA6dw7biwKv
gGwHodgekSSGyQIbV25x2u0E8xQcOwmSFXS/mzMm6bqoCchHJ7hZeg7zKGTr5hQx
oydGzXVA47ThTAAe55k6+UFh1UEevNhMPUAO23nAxwRL20LiVEJcOfRbg+qokim7
x17jO9xjINoOiPMMCK/O7NSfvYQCg0np2/L7f5EHPA3Olo230NdkGPhXoMdfrjdd
5W7rhSxMsCTRaNFxnFpumSl/px/tIaYAeqnJz14GC3aW9Bs90J2KoirnDMhsrE7X
S4JsQGUYg3+H5m98dl+gMIF7bxPEUCq11OJ6G7wZQCWE8hTD7JyA+/qQj14o6shO
yFarck1sEI34BjXOSvkAQAGIOYFjDEZ8wcaOlGcg8iGypAT6raqbl4Jk+eZB+UCh
vUTuH5CTTFENagrpNoOH6SUdKT50OLtqmJChuZLwoJBmN2ACNhDRCGBKNfsfjnLz
aG6p1V+BpwFJC3kv4ho31j9ezrIsvXGUIWIH1b8Z4z8Jt6zftcl9E+DiFWZj8y7v
U65rswhSIYwXymvGYgE14dMcstt7aoqyWfyNNbroD3dMDi5Vm/+acg05tlBk7hVj
oJ2M1wRs1c/smMgFPVPB6hEffzM8QiAaXiyfCEQgc5L97fjM6ZZdMpqeLRc3Go/Q
KWJm5ARgQDbtLhI2FB+STJtlqhb2ec8WdvJphhCVhkiT61dnVbN5C5ZEB9AGXk7S
31Yn3VynGZBQmJpU0GaQGizq/PPaDiMCDc3v1b7CzL6dxnExnmhTeeKCuhNuA++H
qoOc8wE7KhVtrhogA3MLlKbbGqIQfFEtvXq7d3LZwr9aq5KfZ6sN/vcFcJtJfeBw
5Nx6xyumtUZCCTKnYWZ3NSjHP0uY/3XmQ2w4QVosCk59jabkS+1MFj3LsKAriLE9
oTMbdSg5VqoKoKA+sPcxVCGEvYCLjVkEsNqZ861n2n2PTfC8GzeoRVU4FQD6mi8h
hd06W/YUWKeCmw1iwvkIbAf1vmQxOi4RE5WM95SQjJWkhKA96H1DdM8+E4YV7Hf2
09vIRedPnDOiqk4HZouNUDfqPy1IcLiZmJK7eggqTIxNVb/ApNe1BIjVq/tLQpWG
OJVp0Om+ScPB+aJrmOIApMPxLChiLESuS6E4D7pr3mWpM8VhsDxUSc5cjrJoVtMs
33iVjzQDtBbGZs6N4FVBC8RUPzQDUThaZrzWOHvNCe++HRI1fUDaisKSzRO/aLad
P6rF1UlpwnpxRFZaWm5j4UMSINT7MKGwA+v5U8VmAiLg7sRxDMW2l0p5TLxrjiB9
2T6z1OdSgaGtml8ybp8SCGCvNlM6H1KAnWZiXsCVPdubcdv4uhx/BKXF0QvGJnyw
BuFhD4Li3G3To6kz8a87I5PKeJdmwlZE2zT8kfVm89DMyePQpCxQxk0sk7Uf0/lD
58xM3hbWcCXT+pJKR9ZYb3+H6Ks/gvWURcEYnO4zLkoky9dFEQHsmBneZKJMvR9L
ZJl0UYGR5EeIfg96q268TEZzhs53eZYomwCvgsR10p0fOANbN2ub3uOgPf3iQBKP
THi8HtYR2Y8WNIvXPt1pgWPvXMrQ+sTgGE3OooJ5dWDFmmCWvXbM+mPc1DhfREav
WOcqwnLpaUQ6lqgB0u43dqO9OkqIYKdEBpkQpb9Yk361Acw3IuntjG0DsQxOWby2
E5m5uJ+aL8y7gZV0elJQzNrdeUv7pDDCcD3K4FocZJJ6uKp7IkkqNvYrJigdeSQ4
lv9QwY7kNuBQht4FbWJDIUcaAa8ChrkYVY8t9fdvhiUumy3YYver82evD9uQrnKe
fNP9WWtCdO2SRpE/XMknnpTB4fHerPubc3FyqabGe254b0cQe1DemVr04FzYMhdQ
6BQz+54xznPoGvwi1EWfR2qjpWUjq4v2RxMen5hiyDZEymhVk9y/9E/OQ/xclnif
+Ew5OI8YB0ufhcHV34cp69Gjc646Ogq7ca6BNHjGyGIpBjI64Bk6J2zY0euOtzjK
97H3UeeLBrwzNLX2J42p+PpP/rJ8x5kKfh37Qf0mr38084dmWYiEt6eQDweJ0RiA
13pCYx0TzUClpuPsaQO5YlhKie54ejLv9dUorzm0oxKSc+I/SJefH1uW98h4T1is
f5sIqjG+kLJ8KFB9go5oebDC1t47epuTryiBPGTwjCrihbkRuAoLm92RH1GlMBe/
tHLCaPxyM0R3q1ARzGpdSkE9cW0ax8toNeTybHX1SKNFZFQWLFb6vlsJG+rRur/N
me3pK1MAyQc2za442RAuK3jbcnJM9Y1sMSrv2GpEkhyKu4/3PukPkq8GSj41Xu/W
SKAclhdmaM/RzEztoZHd5nbT/g62yLrWmQtZf8lXIW0A+iHUKRRdongrT/ppq2Su
xpN2J2kgy0KX9Hg+RuKG775344y4er9/LeZz4Emw+FFj5IaWUTMooMCirjQtxBlO
se0AD5m27aFlcLuGLabiFyRGcuesFvTx7Pwdg4nqgrmMjUdLHtTwPLG6xpOszVNu
BTUUrn/3+8XZVGhCsi1rH7E8TysPdKSF00RxHejMELh2I7rwqa9us7TYSOPuZFcB
lvg+lmYIXDFEcTLbxLVey0vTgCbOKvwQUAOuCdkU9jQOg5q30Nf6xgmQrpQhtN/f
Y5PRqwsa5yS+Dq08m1Gr7R9UmPuSwO6EpCG6QzdA/Pw0vguNqmU1eV/mqAxojtfP
2i7pkZXJrqfuKU2dGghGApjcMwF1oUZbbMur5TCg2EbqFCAwO1aOnFkwqwIVpU51
S0jF6+4sx6VIT/8Y71z1WRT6hVy7yOA95GzyUQdwblY+21UQAoLowKyE69Cn50Kr
bXLFVcTBXgMLjgiPVdgJkcg2I1v08boaQvPGlr8rWzD+mUg3m07e1kXrnslyEl3S
Y/3jpsTSpRO91V1M+PEkpmn3iWNG/TxJX89C6Egv9/zNI4xksm92pFC/+S80/lWU
L7xID7s6MuqTa2yNwKku7c48RHZQPlgAkqxIG7PytVqsGFJMl40H8fs8KoRHxFUV
E/39G2KNOwR0Yvcq3GDX+U3ukSnpj3Xef8obiwpI/0BjYO153pFWkyIksS9KNSWM
6DxNSzeTI0CUdcZCpz7739HkywFMrAYGkHMtuIX223ESQczqxMU5Z/MACDUeHAbX
YxsnHRYqcecqVGhnu5fF1K9zCDoGd13/RNXZDiImdM5de90bfNh1ghXaMUeU0RQz
gJPOJu4rvMf6yjYJovUytnIneqqwE8LGTI2WH/dOQFcLMyasiOjdtIRrkJNL6bt2
/LF2bCj2PhOxrM8ZXWYU5ersWLUvPjWj0q2yjVeig1Olvy69rO0LGqp75O05nL4C
ppPEsycCGGUa5M7lG96AGJ6vSIyS8anmrGgWgUN21d4Wc548f5Ei+AGqDDeJ5irC
Ym1Fc02iY8zW3TW7qzchtUVKdljNnFJvjFBsSShRrjK02AfnWDjelFQCUi9Hw0ht
p5/kPmSdaC5r31z4X1va1a9bKZ8QJnT8jcdF1BE4mek9zts1L2OAv9JrCCd92c3M
RGkWhyHFSTLtFICvYS6fizuikgxeL/uKpmbpn7YMO57VxjkuIgqUB4PZTdrgfoE7
EP0bYZ87BqI0eayOM3a86IiH/QqKb8ksKPDZAEx6I+XGFKfEyPDQwoBaXRBOHycZ
jqELTLjJ4yZVd99DZVXaNB0FS7RYYu4kS7Qp/7VhACVZi5Jw3G2OC8/29HS9ep3B
mSbT14N59jUl8tMd75YDhhVwQe/XT8aurnFuGNbXq1Pt6yL9RXVMj0aUI4WEggtN
WS6jkEczfhP/HD7jNmYmKFKsYwFxQvfE4Wy+vx4RpoW7qsPeovgRY1orA+MvK6tm
tyJ6bCgo6tHAsU6dqI3UW9JAhXiQi/4SSv7t1hmTDUMvNt9Qh/ju7phqRfpYlE6U
yP5GhyJHqXKAwoDDcEjP/bADp6O4dJeRkpSVThoZ56GO6sXT5h1YCf53RhOUjDRY
BuR0wjaQrMccSlnwQslUK9vbwLNmuJG0FKugJ1bpSBL9P73X3T7ftHxDATmRm1Gs
wA/hHFWlVl9HP+ru01gGkDbU/UCOsG6zVKtdNzJUwAjRFakf5C1Y1UtmRb9OeFe3
cUE7wkxDE86OYWU9OkB+4wCJs4Tcp0CBsBBLO3o7oGN5DmLZTt8b5FV3JaQWpkXm
GH4HoBkMvllZHItWHknolbFb8LsMJ0YygIjoBWguh5se8kfHIwXSAfhhGNwjL8H1
6Z3amjuZRFbIKfsC3DQ4VJjM4txEsEnvctGnUQLTzcaL+ML58qLRRdE+igRE8NCj
xU8x+hDasmfD/amsaybsQH+pczDKs9og7RjaiVGZkVRZOkKN4pCOggoo42aUUNzW
nEYW3X48jlxvf2itZ6g6xpnyEsrDZ/ieStZNyHQFWieDbbX772E9+mWsdhyvY6HI
PizE9LG3D5u4FZv5xQtZ9lNI0K5y/jjv4L8xTyFQ4S+yO9E3Y3gQmRRyTmE1LVUg
GlcVJj/KYgjgykFp8OwTx+jtCUkrct7oP+XtQbtp1h2VYKokP904sxN9t5Fr8ijl
J/Oxy7Dh7abFot1Y6ECUuzjpCPPQyf/vSHOoecTHEm7UEGeqmLM5tbDt6RJ09Aak
hrCgdaxMBM4XWdwFOp7USlSjNfKR1bI7kcoZRE8Q38xlU8Bs1ndP7eIYnYHeIydX
ti55yAfv5NgSzf/6aCNVv8mNk7Z0QX9o9A7njyv2VS/2KMq3iDvAheBf/gXpbiUS
+DLtgepVN+NSAK1EKuqI1Uu4jHhKSBusNxbe+yNK1+SMtf6RLA3jhmT2e5JnV7Ek
ant4fwtrnQCqXky5Vs7YkcGKcEYxB8C/J5tVzno5uqJ8jHzBcGIkIcTzW/agZ/sd
HMq2dyrIFH/AjIVglh/nlOoFO3KsdDJLnYh4lJW6r/smmhhxCwlaLKH1+H4fHhsK
20+b4Hekv5b6Nn8RW3B1bECVfPv0Upo4OUNURwCmnRojG2KE5uM4m00FfxqsZZYU
GBsjzYlXt6KXxk3NvDu3h9irGENPP3kyrP7CPFnJyNFkwpcIlr5B3u/OKC1rxmE8
IE7EWEHo9eZnmTxwYpzIkZW3KsXXC3ULIaZxkLzXAePRQpToz4wQebYfSAS0jbu5
ABhBWb+2lB7dg8Xc7ykkm/WD7BxtdqBZQjPEcxFWecTU84+fyEJwuF6W75bYTbAI
bFvqMdBjbRK8IEVem7DAkrDr8SMSn5m/x9Z3IRCA3dQq6iKtdRC6Q3dNfEaCU5wL
esykwRTqvESZeXKHTSJM5aHkgJKTyBV4cSqSOAyvAZ7vEZwqGK4+ItQdPg5pn1H6
6qD5LXOr+6LEYHKtru6GIg5Yj0d3q2lNlusrzcHv/ryq8xwbEY8qCKvQxqcIiFAK
9OBSBYbSCOPIPzCY1ttSE7GHN8EUzhtz4ysG40jOQ/y8dc/6cmlmClTEVzG/6qER
tZqrLBHZNg6Aumn+D1v8a9KoZ3J79APA66xZ09AWhIBX/jNQEdb7YZ9GXz2JiT+W
+Q6/CVykm1/j7sO/nvbHtHLfC01Gy6pQZ4sT3gzgErQFg+NeLQkJFjIDhWKLNNHb
BhlA0s3hM0XmjLQgbTZnGi7xGshXVTOqI6JcI3S6m8cqX8qOLPZ/Oi0uE4aoPGuT
DxYI7h6tBB6FQBYgJjSuuwKt6NohS7xiS0Pjs4JFRkv8ZfHS9f3TX/QRVtS4NsHr
fNUgqBDh2g8n+Plf6WpynQUwPMZ0uBpbDtP/46nGSpX5UJADX7zOsdpIGLQttMAI
tUngrbsZd+mll8zkv/A/+r5Yomkr9B5ohBm7q2/NDg18yPwS4PAoBtF4eGhS0PWi
b12GO8WXn2VKOYmmfK4VKyrs9cnxksIqZSTEcis+AKFCLo4ce4pC8yMDW7cJrmJ0
qmsxUgw2fcmEz7CQLJlvt5xFUHxIMPemqnl4Cv84WdAeqnxdcXjoqJOPZZVjTMPD
xQT7YVBnR+rjE3CCqNf2GFUABn0EwjxH08Zfdg3C/ydrIKn5b6MrtUeu+2iu9GMn
VzvCHYqMk4qMXD7r3bIyC3aIQVtBNPBwHiJBPVx2Ioa60p+pYNzf9WERfRUjjQ3A
Da9o2xDN8o0fLaOR0350NZIqU4Ld8N6V4tU2aZOnKegNZSowmvvzzKG5dxuWLODa
ecOFhBOz8f3TMZ8OrCQqiD6aZRO4+Ok3PtQfaAV35cxWEb/2H9rbSrLYgGcPPeb4
x3a8R+W6FWKqGOyYNmL5b+WrDRdUKDNsxcAX0G+eEigezGFGtxCXJRNkLl9viTZX
Y6NGArxOLY+rDtSjtS52YN/6hAe6KWP7IwEOHh32Zza/y3KtA80FXqsOhGW9nTYN
T8sAAvcQ+KCpFjM38BQ2cIGWCszQGCfjSOH8uPj25tTWqEjxqkm/FRh4BLFOo1ml
3jqx0X16ao2I6Ggc8KdhVJiuNApw+jKAC7RBCpn0bdzvsQIAtJNbedSSGv3X7hBL
9TysKmjFZLuAToc5XJG6qFTmujFVBjlzlqaj1Aclqr1Li0tMl5zLEn5Ap9+0B940
TqsUtlZkxoVwOgUYLQwc3XExR/Xv3TNR+9iurgNEFMnOc7xoURst/J8WpO8kmf3r
PXdzwTcZIIRyH81m3qJj9FMr0abiLB3/lCvdEgurV6FysevalVG8dbCzs3ByP573
VPSxCC0zxBGh7N4bm2IB93IwNnx3xb6i+PmgAS2qm9FNXA//QGXI1McAX4+R59VW
+TFJk+xlehvrADg0soV2wQ6nD2IB7C0vVmbB7LhfkUOLeoovkSGX9xTeK9I1mnPA
iGUOq5TF46cYm7TP2REdhReEOmckKK1fiPPkYvStLYwvn4nSjT9cLg+pSGqCKjhj
JHLkBYyV4VWGv1RCHqJwbAfefzQAY7/058gOLWWB3cCaTMRlNKx7ls747xbqvivZ
UgDYmqQ3ZdeTcJu3pFVln5BElde0bZ0evvz/ldzheR7+KLJuIJivLpDjyufIK0Lj
KrUZkAWT3nXaR+FSdaUW6Q1t9Xj0qDs2LwAf0zsIHjmQbee22OLPLIqdAT4Bb4i6
61DxX/pmbLyqbhhkTRa70HHD4ts0JDv4V2qJEGjyzGfFXnLSpaAaXqOj2YA7s7nS
VkltT5vkiSlbq/hPKTqlkhxpafS3M8AmfafrarzYCxBR8J/f/5Rlqp7ZPzJA1cnZ
GA/XuQQwmhnSEQjhDYUmYhf+YUtnzoXU31wviVGjjUhPNdBYayqxUJAssPENAQeQ
yb/6pdSfJV+2dypQPY9rGAXW+GdpzOKZ98RVEsjGrlNpHtpEtQj4n1B+GYwak50e
SCCXealxBV8YKHOY4aSf2vmt4J2aFAChxXcjXc8w824BzH/gX3tjt04jyrvy2vGi
eSKSpAiKKCpmL70OciTuH+8sS3MIFh5UrZ+yLxVe+3MwHLX/vfwoBvfFmfZDNk4l
9bVzjLeJH9ecLbmfnfkCy6cDCgOXXfhhuG6zW1ssHf+hXox7KSt23VyOmFIU6Jz7
jPY4r1zf2mm6gcLEgRGMTM9jh/O+iXxH/o5eznjtcWwk15e8KLnH4x2x/WDfLPRo
udJLri/qBczmD7Bk9SUMU4Z/6mFy27fStFQ2clhW1gJ+/yqFByq7Rq9hwwPhJPdO
9KoiQ9LA9YEzF8o/ahtpDQprmrEChUS9FzcB73d1GcyDmiPCvbraaxJ2bprFg4jC
LEMHgWurAibhOR63PRk4NdkaDUBHeMtdA37YTeWs1BemCiQdVZItM++TvC4SvNnn
j4uGPk2MqA37a5djH6khc7ooVUXje+XnLFzLT+VcUevv1ipD+QP9f5usCx7GxTNM
0cKqv5IMbCNgMYGUjHY/vDWTDXzWe/L1sCNainmPJuoj7I5L+/4cg1q4toupF6yM
ctqLMlBA/7PtOXdK/+meUO5+sI9iLlBYyRWuheYWDMvZLjhd2nK82pOD/O5kWREG
2qh1viH2gTmtgJCTchvdlr5pe4XGgCs6DgMZzXx+ki+jOVql0QuTIxpZRifTA3Sm
xEGtOMiCGLcotoxSiuOwMPPL3CSw2y+qOj4GY+PxVohhLNuAKs5g4+ZKlrUTrWoF
VeR1xBjCxsAjAXqYSbxgp9RWSbws0K5vMJ20nF7JEwEJsYrBvMD3odvuumrtS1Py
vpnmUP1PqnaRPp5HXRhuTFIHtiSItW+4es8RkDgigdo7m69IhKw7Yusq6GbcEH+M
gOG4tuY7WrLBQCOFvZiMydpIr0v0F0cUQDzfTKnZ/S/spnvJPbFl7oLc/7pAHVSI
vJe39MX4OF2ow0SCF15GCynRJNSr8XlgohpEhAIyQyKnzCzGoX9WYz7WPA5d4RYq
DHmBD2xM1I1BpyU6MrK6pG/K0VmMkKYV2qr4i/EQgJ3R6ljDrsWHwpPY3Z+HuUPF
izKvRW1vKlB4Bump+ABblbMjGPif5nr65xgDE0aIZaD5JBNL4kLJ6yuEu3PhLh8T
4XYLduiSa9RhGjCnlHYg5/mKbiPNdohcGs3l6k9/Q6DMS+x+lW76mliBXi6Al6Er
MBdvSWU9KR/0b1MSyl3ooC4sMvMj5eDHu/xBPARJQsgRjFkY1MDAdLVl6ZkQHyeE
SdlkMM+Y0vjhtb/PdXgkqSlbE1Qq17Tw0Ah2EhnbQACmqKrb8yIwvV+RlsR+G/I+
5D4REpfsrf4qb/xYfVY5n+VljsX2Q/t0xoz0Zu0F4Sx2S5sfvlCLByH7+fRCbx/+
L+m/8gUOE4BAGUbVRd9smz6CG4b/FbXjUG/xugYvE/9qop3uMkhKpfmhtaj0Ee4+
0xmKybcOU3K3Xs8aEsHf5VgLDZ2a0rHhrUQ7lYKRkgbPj0tGO4S5zTQplXrdmOS7
syAdZGOLaJ3pW+SG4yfxtsAw7Blvbpxop+AOHj/2k5LiZYynCSyXzG18hT+eX6g5
5h+gkYIhfE3mVagKX/PmR9r0dnxqokCqdtKROPgC5S6zdh1O7udGtFTU4lXO3ILE
nl3S62GM2uA/+Xg33AP4jyb/htFWyjJSGmurOSdDbCTWepTW2fVYtRZvv2s78xuy
FK9Y2jNm4zboeORNSqn/MXpaXjUvAn1+h5wrchCMJ29r06/CX3zWKhbq4vgtFCcW
bGMbcn50MtkBnYdOqh9B3FpnEE8vAZHZBBUy/SRVevuogTEe6InHgIFibvyWh6mK
7TUSR7xPyDaEY2YP+8qAaYaXz4QHooMQWOr4ilBm7KigYYDkFVTJu+wWJ8E4E3wr
jen2SC7pjjtGRAT4P+4yRLew8HHv8KpV5MepWhUKpXRM4SoqHhyxEn0I5DpvQSxc
68acC2+qV1rHdNRK20SvUQkY+3QcGclYUZeO6KV7aBwnG2AqM3u1Ae85ZACl005m
9PplzeMboA0XIW9/mrXvgqdt20Y470D5ek/mfBnnzj14JJ2rjwqfUtz0HKdQGaNu
ZIvngbpTZKk3tzb4rs4z8Fb29IytGauFz094CWsE6PsVBLMEVjsBzFqPUbFpplyR
XN+oaxQskZ52fILk6rsc096qCnxZXXCGjD8U3rodLBDEurhT3YnmX74jDm7N2Wkf
QwF6Ty2z5P0irEsuyZRV0xlByP6KCeTJVWw2ZWeNBhRb8AxkTnGOd/9gLIcb2vKF
721eeWHl+PERlUl1agzWSYrTwVoGU59LnieF5TdLI7lqxClj1Qhqtl8U/B/+KQHx
KwQKhuLRnMFBLCBOA6q2aIEtU1ktZlEet4g6G8LeZX0Yt/ayqgy7ZaJ+0DmZcQij
Gb9Kq5oBB2pgi5dixqjjtwANrLAIuGcQtD6EZpQ3u8yypCSIA/Xdp2b+PL8yi5tp
lcqYH4PP/cJ9iXji7pc/K7h2j6iwTO2Y83mtkfFbvXsXd8pQsaVMTcwk/jG+xufj
U3Ujj6m6EsCP307m5tlPVoVZyvR1yasp23dxpZDZIli3J9mxXt+uvJfzUc5kcdBu
POnwO10652/PLcbDjSBFOBXvwRDX2aUdBru6q8yqmWf+eyjc9srsMMBv6ms0WLSt
30kYncHYxyqGWinx0QWFjlfJLaz9Oe2jvOMyojj9wpbCzHjTOSFTzxlTqPKlid6p
AVKzLhYigM7tKR7v+8s5UejFu6VEjqT4Wio7wOGLCOzOWrtM0TuzVriXogKRAHSs
iTjjinwH1+5BKKYqHPJre4sdvuXHLm3Vs90cWB2+PVQa3nkh1seFmoDsaFZKxcZO
/dZn1HxmIpVL7v3LnDS2kTySAcU/AdB1duKh4HlyxDhxEmzVC2/5nX++OP+bpKPy
7DoXOj1oyXMoaxnp8BMLqDYvqZv0mvaipxGN8RPV2rRP0WVcJ48wPJLhSHJmmCVb
jgPjNlDwW7CY9gEsPbzFqf/n25ItZjHDzio8GM94X2hrpeySCTeY7cAOP3/+mnKk
5fx+/ckpNcmpP7gtv+Muv50zApdTDVoAy9xBXLnIUuMIlqwuZHKLiwzId0lB0NCp
TmjVdtv9ZA+wMHYw014PwDF/Nf9yJowUT3ZLObS5wejiVFm8yN7IHTYKezg0qdJW
OBeLrjp/sU9mQY7OAF/UIle8c7tAITXllo2zocEVqfCet4QMz+DSQGhXNsjwg/RX
FcPtlWC97zcaEN6LtdPBcv8+wM68ci3oGZDk3VjeJiwuNB8m7drgydyyplXqHc/c
k4oJFnj2pNhbVA7NytR//dkwJdsbXPXEwZ0X+qfZ8e3Fz8YGEuE6ZqqxY/rpBrQH
ZD60obgmMDKREiYS65PUfCcRcmjtWtBG03rPH1S3Bhpv7Nj3uapY3PlK2sd+m8KQ
ntHpsqf9Ub4IvjPyheMfSybVfPjRp/YGIkozIujCCw/XzVfT3V1Js+Wx0dFH7s5y
FsJL1UYUxXmEoSogU5zuwBIC4CtJzRi+JA7NXXGQwHvdAxlAsvARFHfv/6bcZ17Z
arfcXLMdJ4VuAnigq8G5Opzn2sQxXzSBs80v0nL2l50MMT+21EoRYhZoTJgYFkpp
jglD7XqPliQ2MU6QPVQIVtIVLECb3owDZPiTPbhyZZykggMzTnufJ8m5VxqvM6LS
3gmBoaBKT5TeMwIjK6uYDy/MoOqdvhWQLaH4RFbqHW9zfyk4D4IYTTaSf6Wzvqpi
9+7LMF7gufv6RR6DDKi+aTOCa3tLn+besHlLu6J6Va0V0QqjWjhxzcMUTPZ3W/+3
gCuPK3UyE29t7id+4uxZQISz/KoSgNqGxHBcg2nRkstadOn+CQKoolbVgt9Zt76l
P4fH9euq9P3J9w2Vv26QAIaB/cCb7IivzzpJSvKcRLAulqqrrsa5U4QMvXrhq3no
bnhjat3eXcV+DxzEPFIjR9qshy8ohihx8XSJD5pt+1du68mUFCIByeaQVJxylgZA
jit9GVb31tMF17GlqVG044mYO4o8qW6S3tjpd+CJ5d08FbcW4LzQAyPY2jGky10e
JomYGf4LOSBTnWrOPLquGZC2ZBEQJJdyovtqRyXWfxb9L5KW0SojKD6POAh1xlRS
TfyF97fJSr5esizacsh5HtzqcvwLeiqrlZfu8CnI8n/JWAKNt7d4vBixwPWI8It1
Eg+tm8jpDPvn7OoQHbOIqAOM2Qacr7fmD/ha3oyrGo9a9NDWwL0QbW+TQDRYhKvl
YZYkvdOhIcFTKlb0WViFw0/GDAzjD8/xZUYOSA9OovPcij4j1g/nXWh/kiJegmpg
Ew469g4YfOsQhHfnxIQWlJYM4s4SX3dyVAyu+HQUQ2ow90bbNT/QHTfVSk/KtfSG
nfVax1ueGZrznCfrZ1m5jpxpr4g+Dsp5yqwoav00a9gqKdKQrbgI6pvSQcPIkZPj
9dhiSkwKAAXvKaQzv/zDbzXFwphs1OGDyiS5UJc5qy2BrdI/L/a0A6MO2/bUvpZM
fAHX99aqkYF//PD423l1y7hXQp5F5cArnpk4M/mB2yel02ske6AmQ0NlN8YxSDag
bYgQl40ji1SVDISfhzLnnXGPBDRT28QFH3L5H+fKdg89eUU5NIHncg8OvEoe2peT
FIhn7WbvsjRtSYGgQRgHt4w90v1W0QoQfisyoy0wYtUb/uwfcJgMm2yGp1EqQ8fx
0kOyv92LJERtZa91He60jKujFyRWlE8tjZ2USReQ2E1Xb5tiYO6NZ2iFfWj19d1V
34TM4DkpnycX2psJP9UgY7asKWe5LuaqjGjVZo/wuGmzKh5a+Bv8MHoYSY957N+p
gFyoLBapF57B07/WPEJjNykhy0ANGatdXIXHHhdqZs1YQbNQgL+P4daBLTw7K/Y0
WvREJaer8SC/kwiwf7RmaNTHcHh5iDQsaN2am5zU05uY7nB1PDL0IB8+SwcSkayJ
XWbTGYVfqWfSTNSa3924/O4ceJ+fk66x6xRuTCwe6f7Y7Qq7Sbl7jazmlKRDkJ4k
oDBElm0ajvgM3xVfWLZ8YwJYEQmAjrc0Yf9L6oCMu3tETN/Ji9VWASv5uP/9O69U
L3m15vM4m3JOW+iBSeRgq97J/t4bJ7Y79eHe0/6KhjxIqy38+5c8sNmkjA8YZeZl
eSHXSfpykBFXSHUd9GQznbhLV7nOG19S3ZcBYcjscr7UR3sbrDQSjO7ToRIhyFNt
J80xZkgq9vTI+FIfON+HAUJT8MYlzP1gpwHmNkGoSPyO6EFSP2WYKFO8sYXXZxYz
sAvs/Spdk+Z8erxhqcEWufFCwT2cOjjwmtDf3T5nLZTcnJ0F+BCEsLVeUzQvLY/J
pnP0mk2gSr+OnYqnCLheB3uo/WHJBvSY0URpvuKotTQQSP4QXe7Rp0X4+1RTAZOx
yuR0D7ReLQsn9Vk6ff0kF4j9fb+NjJiPlNshI++7oRBcMRfM457AuZOUpveCOBFX
DbfknRi4cv7QPzkSdZisSPqvY5OLzORf2zm1tPtFmiNae1DARboVcN1vHW4LGKPn
hX1koU/k9CuedeqRZw25CPrQvFGO+8Mjjg+JSqNJHkkRXL1x8N7KiIi3XumTfS5L
Yogov85V5Yrz+PRVtvr+KQQIrOruxsTqiGsU/HbmlnodxPchIUd8hnfYA1nR7bI9
GtnI1yfutfF2XnqjV0vwHDQnnAwtDCx48zA6ptvQPKFbizESFdPtD3eQ/606Qnxu
oGcRwvVZHofQHB7NFqyOP+xChFW6qdG5dNNysYg7dFVv+tS8GWKRNcJ5S0wfrVzp
Qs5YKFIdUl9/ksc3utY7OXGwlL1wkxFOdCahmo9Kn2p0Hd4gVLcoAsCien/cBvbn
AI+NApc21eY42AcMrDUu+cQshDyr5Es6iZeaylDymoxUkH9QQ64XIGCL8PdlqQEg
mqM6QANngi1Ns7mlj8Om3EPy3icJXOHfDMZbkmvEkoxaAGJmzQeTGQnLIaEZYcdh
Z+AIS+RbM82fU4s1p1NZBWpjU1XjQkVbrDLxROHYGK3S+ZMAjAT12Trh7cnkoiFs
OSSsnsOWG5v2Z/RQMXCJ/8jW61YLO+lQN14TnPZTqFNwpYm8ebrDKLU0RC+4SNwj
7/M4mvvc7q5LRIzOg4nMxP4TBstUOHQ4jhz/+t9NEiVK0ezpAQyUrSBn7osyebd3
NQjZrySJQtxsa0VSa2xZJyQTsYachesoKrTd8B5ZBJvUR3XXnXTv6swJEZwOBg8w
FZBWe/rtmF8eNGh/eZSfwoUJMxoKmErJZcCSMILU3Dveo2l/BHk71edxQ6sULZ3+
O3eBqmlOqPNxsrOfJyShDH2BC0VsGKGlsvHWYk8GiQeQIKsRe0RqlPqnHlBGtxnP
h/thyRer4Tb8S9CSmw3a5wq/jepOSp/0XRQ90o2t8oM2GHBw0tXz3vGSoYYvbXD4
W0JoZmFa+ezcj/cGwub1uXbfNXsiLqD1WLMPP3ANI3Pm3KTQ8tWdWXKn42fZp+b1
2lWXZX/dI70TJYL704C7crwZp5LPmQz9ES+oE95jTWFbKS09IgLGiDXXpOu33W9e
dxJ8DzbYt7Lt6TPp8dpPFkbJZ2unZXhR15xcVEK2Hxndm5faHwOBVxuL8M3Vu4vI
DGGWJBYxeGKYCYRjw+24oF0D2AJBtbkcVcAiuz6GUkkC6cnakGP5Ns5OHXEWtXCx
ynTGoshzSFlc45UxNSkgI0j8Nyy93NyDX3OJcSs0GN0lKcCT63DPR3kiGlSMwl1c
eJIzyvH6WXxLH+/gF2QoTU5BM3LFVJQ09IN6AKSIrIWfd7gX6sG7R05VjWsMouPk
mbmGCMBgpGRkeHSODfdwaGO4XO5ME04ga+FSrDSDpzYeQJYYGX2AB/x6DBmmPa3e
X0l2pHBXeaG7Eepbl08X+RRovepx3femBlbEiuNwrh8Zwy3rBFLNUZg6Mp9o1vfD
/SS2d/DFCShYeadnqcOZB3iH8Xm8kB5PRn0fO5vzSnBjLRviCwqRpZD5oeFk7U0D
VBdb8zqLjFS9wDBqcE18n9w2bypFJ+6CTAU6CDaVwyBS1sppuO3Ob+m+26LHddgA
Sr9IJ9xIH8YvFd0MzH/0xXMV4zT5+F5JT1YEGz7D/St7stOqMjK/s0sLW/mmKgWQ
LXHlwfpX0wHQO3uxMAs7dvfnPWXh1LYdWz0NEZ5OHz73yVTkNdNQO/6t4AkKF4on
qtQRwTDelyUiE3xJa4JH35fdx9qyMHl+geyBqQP1+CZyTc8IMMqO4AGqnOaA1DO+
1qdVi9D2A/sxIHqIKuUsjJchB/35t+wXUT+Tf6Mq5SYGvDtCSs8i8L2Mu2+g2CFI
2NcQOaORUPDgvAZlOd24mF1UwOIFwOOjHo9ggC/2/yByvorZf5R0OzOn9Nfgw2bW
LU7A1WvXQlwqOKxJdLwM8Hv/by9lbijqef/5vtsmDwwBkhiCETF8NcmKs/gjlDUC
0ie682cBC2UmLWFszvMPv4BHB6Uv3Uo7iKmt4f9QINM+1mzaDWaOMt+If5pK0mme
p0d8zwWHxodpiGrvF/a0YQmQMZp05VKFsI+N403JnBauvOIMPzh7uijeb3YxT/GU
vseoZAZsG8YvzLDAyEjYW20FMZylR869cOVEoHsI1CJzSe9zEJM2nDQmF/IwfjK1
E2nemBcuDSAiMAd2+3DZyJgbq+X3bu/FKBeDyEH6116IYbHXWvbmCN9/51ZDZg89
oiX4Kw18CcIpXF/p25QzmRzTiVV1H3gA3IFv7wQt0UCY22PdfoLVo6w0lahiJVny
Nz1BBtJdelq/R7w+7a5hl0Ny61cXSBfhVKfgyW/2IV9rshSip4RCMKHjAQPjPQ9x
CUV5lIMl0UeXIpuVNoRHpINyExr1amLijlRXfISebuBKTV6AFAF4LdSEJ8Ktbu+E
e15c96M4bmsjON4XBDUzUPysd1gkXokhP9sbLSb2uPJiLrwFfyzDjDKdxdA9YhYU
YcPUx1XvrRiAeDeu2iHgD8tHJXmjlQ9MgWf8HnD6v5a7yAuvpqYLlxdLdU5YEy01
V8MGd4oLULgXc/sjBAEycXeCtIxdys6ww/0/drLTvdGWTGssu1nYkV8Sy2ZdlwUK
Xo+SUyEpXOe89ie2vM7GU/x9Iokc0WKEV54F2pKZD6sdofVihyhEisInRbi1aQYa
OGi00Qbf9Gxr/IrNh0ajQ1K79GWOAvmp60ohTnUeCDxFnv4IjZ2i3hwQJ+z8fg5P
TTxOrNBZ+Qt6cIAih1sAILawW+o0+wnuZvt6HWUhvv20BtmhVvIMLmuS2/C+HUez
S4v4t3znVTDisVHzX/LLxr2UGHSVWt7g99AkdyWQ+pKSDzep4y9DoAqmJhMQJ4ay
dWuIhNCIMakqyg2vWReivj+OnyLnp4pFdigoy3psd3cLBOYi4ox/ukWLJKgAnwGP
sYrsDsOZjiQX8AEpk56YV05U6f5gRH9R7JZO+tRbyf0RpJOvcMwr8h0CTnEk+jfm
Qq5wWaeABql7PhPu9zY59ZZ86wvPSDKrOxqpLtayJcraHzfwMXRPhRzO9FbhN0LR
KF/vfNlwLhEN9/xfJ8BAmqKXXBejJJrXUsfnbTzFaD2X2ERZhy5ot1GeTd9xB9xr
4lVdEUHlawoNlyXy2ai81iP4F+W4wVoDrMcdEso++erQbVlKdJgXlGrXQkp3L7jE
nBlMVragGZF3DG86Tymctw9+lAigGcnn4+YX7JJc2eOlWdVEiu4P3dlnGka1YAhR
komvIuSvWzXROhcoDBqYXLb2LfRxcfOO9x/oO7XwnQC4tKiBABF6h4+qJ6CHYgxa
9TNY6l7jHn8+TnAcjUDwLhe7mXs32d3VqN/zBB65HwLzCK6HnovTRNe1P1JQ0POZ
reOieJsmf94/8TxUS3uPWPzsCLMnin3XrH6wrP/cb+TMLQ7+hPN3gCR0jAWPmBFV
LHL5/iFSpvroEFMhgO6bAPjqVhouVpfjNdDLKeStsNpMA5CZlw40us42DR7hgWv2
MHV/JW8BD1YhFmLQ4cVS+aN9g4HEQZ7jVc4RfiFs52HDWz/h7AOy0uxm5kKFqg5l
Cerpr1xN9vWlCht1qlF1dKsSGH8jnsZG/GZ1AjypVCLB6kaSc0gT++5GU0svDCOA
/mDKNrNvTM0t8EdFlvZMb/JunSgK1bb8P3y0/sjTnStZuwV1Dsg2owv9jP/uGKPi
E5RFQmqNf/LySwbAgvBW4xf4iOhRzSwTF1khAwzcCZgMxhPVqiYzmuC2YRr/L/xU
3QhtXvYyemZxUmREwwIZS1BPkit5A+OULnrLk5PETcG5VNpSyIiztCgnHCRw4k21
oxnO6ZPLOgBRcBC6XGkHqNuTPZ2uQI2EL2CZRQ26SSUuN28cg90X8tldL9j5NObA
Fq95NUsq6TWSCrodXOPfcYvBa+XVQorUNUp9jWr+n17aZ5qMjwLSOPkRPrqkY9r6
ZjCg0nNlOjo85NvlILNZl5r6X1H7tIKmKmL/JkOc31IihhLs8BYynK7PypiCCf+0
AFNfubllmD8HT/NkVf62sxMrJG7R371E3+8c300o7dOtqU1sy8CGZ+biwJDmI5oQ
HVxlc/CDu0HGdkvy8egFJmKnwdK+8KK4tbfBcC0CRfkB9PDq4a1wYjj4y6oUk6F+
L5rJIaj+rRw/dIf1ii9JirsheM8PgMRF8PeVufQVvH0P1VTO5I3iqSd5VUxw4Ptl
q1oyo0kar8cLxnXFUO4cw03AN4gGDoVkGjfi4Zgn0zsWpDpAAJXblAklSPS8o8Kf
i/ih3r37nh2a28iC+xFSFBVLA6Behethwlo08VvkYBdyGINVl19uGfC0SxpQSXc+
YGQyyaFylSCKktNQ2O0uCBdvDmGggwVKj+JBLBgNvTs7TOPUvW1PKhI2FICA/GJ1
3vfVYjRzAvHO6FkqVUGwyyK7Okx8O29kReqaOqKbBz+nnyJmpmD7fwefDkSD0zDi
U6Fz8QJrLnvXYZebAkBTK8qrJOD5wESeZ/Tyg3DVm+G6h8Dk0UCcafLcJzBTAWW/
3QlupdClyYudDw2HETfqVBe7Rt4oTF74jrOKstfeNMELjr5aR1wtTWzjTqD2GUZK
1HqkTfjar1mOp39naCUHOmyJ3VT8ju/hvmBEfVDQLxy1b/RMbYybH6WnAr0iVCGt
pqr/gyvbLWznRdY8LTcItJUqoNlju/mbCrlgsgwiqom51fKRS1TwFtU8eWZEmB/o
/gBiC5T9eHUYgybzEsGwpAif8YcAgTPMyrrJ0kvOXqbVwSASLLjSIanKenl6Dalz
/DIxdNPUBTQtExfVTytnYS5oGHu3ragruz6nQXlFGmTpZRVhPtPPvNyOOLPm2jgA
XvU+YaPVCvtFSC5oAhC2yI2ghs/GZCYB+MLjulHzaqma/DX7XWH7cvqqoS1Rp94B
8sp/HwJ9uk1i36ftuREmk0WYRs+3cF9WZFlFU4umhetRevUjd7VhD5vFrrnETwMe
eMhD6ZKfqoIAzfCqQEocMBUXESa/YarVeX3mBoySS1b55InJh3fTzzHYHC+GFIcC
YUHOXSYrFwaWPG651eTmMdByZXZsaweAvzScXF7PzwPDvaY2MqPIEKbFuKKJ6jya
yWa0Diq04cLkNfnmat97lETMJAT0aabEHvW1e0zkWvIUnrXNuX+9nM/d4p5NjVgP
6XlfzR9F1kPbGr4IEJydm8A5QeziesQHjehuM/+YP9NWv3PQcFnKTUzQ7JeOJa4x
AYhVEuAm+U6BggxnH1afWD3nMb3ioztXGjps+TsDfk03URJdWQESDqwFkYW+W49Y
HEOQUsNXokQxCnBBHhQZJ2O616jDrCvJJeFPLd5eOWqHiHllZKsWOK3F3tPFlZ7E
N4r5Quf81PElzbiy7uvfQHpAg2XzH0tvUz4t5pqVxMCy6/GKFXyNdEnkrvZyRPoO
j5/oUpCHSxYX4/tEi62ZID/fbqTVUzLT+o31VLtk9nznbZfG64EfzyCXzDYh3Zds
CUQqYi+KbjX+S5YetT9pyv/1SnG++qOUIOFBbdVTlctVFhPormokQqTMhH1U0bN7
mwvPXnKmMAcx+8BIcIau51pYSmC1imA0srUVZs77BSoJ8q7AOkCFgj8GGE4BSHvh
Jq+KNdEPX8C9whKASgMGi2XYtJ9mBwu1YSJZWySj/cUlqMMdZ2iYdzj2NGSqspiH
jtaCbZQiw/AIEw/0J5v3OsWcesI6kOVNNqw4Gpl+hMMgVybekkdy3E36EX2apLly
6y2QBCtmcEByKPhS5bknGb59ye+AALl2dJrLfxj8r8T7LUDqExc+7lOCOU02kdD5
uEgMAPJrDXc8m28QKDp1d9Sc1M9txve7pVVVZqDAZEqh0JVFukDjMnKUsYfHSMY6
fG33ITct0qglT5Tc3aPjugT6rZ+xb0bX2Iyg0MQq5hn9+Cdv8k34bQ4pTR5R+PSV
JuBY7HNUWCL+35eNHqXzWy0t8OpNRjL8Bg42hkhcsC4UE4cgewVK5hozRjUULdEL
I2hTJJnnGXClW6gsqJlhP8T9YILzpuj15Ch6e7dNrvkzuL5wIl48jns6M9CNoOPG
dUFUlklp4dEEmjR6sWzpfB+29j1GdZscswE9lUsb+e8oIudYLF3GY4Bn/jY3leIz
iTBU2qdeOmyYdss4SoeJcxbu4xWnKb+XXzaEdA2vJywLIKCOSyq1gPyA13ymGv6c
jkBZCX3zeA01wZobvXdj8UYNfzDhYsBaT6kr2E4KWi2SK079jJVRdOYQhfbhONR+
LoCQdSNJqXcookN4ma/Lzby9BjfE+3xw057BptsUn7kaevZh8SQQq7vlRZlseREL
sUd8QfzEoT+56RMjhWEKI50EosUKEEIHWpvH5rhyPNu/GIkAHNZ1C5GNm/kR4NpT
Z1KYzk9aONig0bz7WMwnz1hnN23/AmBnW7BV9wGsT8TeXj/MxYzO1TqA/2cxpZD4
vdisqfErWKb1kmfuIwencsn7ubr2qhfaQ/bO5m7J4bwAsYO5p4y2tex72DycdgOS
nUIT+cWK1SBcq/HbTbgB/T8ujwp/QPlZsnyJ+OlAqeqC7DD25QaK2KE/m2HV57Kw
feCDbrwpTyOKizA3AT1je690L656XPvenjY5JM7+xcFHZe9DebzoZEc7cdfLnYLA
xxaxKwHqvUqbb7iispNUXrj4j3NmX4Yy3qyJ4rG01R88X3BPUl75OkappVFhiQe9
ZH5Q7VSaUW9Q8rbbv9hjztt5emajwAJqY/MyM+GPmC+0P7Mmq0ie9Ng1CSmaZwbt
UJz/+kKeurlbW8CrUWRUprbtv0QJWk2kb4NDbR8koU7mbdJr2mrY/3y1x/jV/ezs
E4sjpbpzVjuIxmo7rv1ScXFi5XRkrWYRxYQ90wOLrsXIdwhmsUpX5zyKMSdFKN/A
wqoBHpQzpIt0NmNQmz8oUmf2HZwtZOGZ13J9HDPdX4lhBCiFkn+pMQrNtd6Oq1Yg
TgDVBDiFR3d8Ep3nPkJNTaArYRH0YPS6EnUuZ0iqyxnri7YSiSVQ99dfC02OWfRa
iYkT+QVrMEgUATHsPf4mgAe5gyYegSRBHJANlO8BipHRlLHlQpm21x0m9F1Zhybn
ZHvcd6WAzbkEguLXbtxke1yy5eoOrecNjtc+S1izl1+uUc9ZW06WSUDURWzsr4Dl
16YcUPA0joYcLpnMnBREArIJVtreoG1fZ7H/+t/gDRPrALWB9KKDjnAwJU93TufI
waQEC0ZhD5xocp6tZX1uwUoIam18Qjj5f//tVV6VBiuaYoJHAUSUQ3dfpUzoeKuf
ky06dDyc/D/VA/0gfyYB0ujUsM/ggxY7nEyaGlW4T/LR7b7WWEzH0fpW55v4/ULB
PBHSwRhlpyb+T0U20MMBzs0H52AWC1oLfRWatQ5Yx8uv0yMReV+OvhfrpmxD7QMP
FrszfmTDv42N7JlEYSpTXJCNxMZkIbqul5qy1M5Ccjdv4lFLDoDgDH/Q2D99AUuE
8dnpln4Mwh+UGnphA+F2xFsQNMAayyI4xEb5NYI+A7TfcRAQ/L9U4/L9H7zweQPN
KRdoV912b04zqCal7EUaeSUJrQ7b63u3gkddfn8pzj3K/yyhhoVUi1ZynDt1dqJO
rGJJvLbbTV6Vsv0+IkzGzF0I5IKrlSMiKDGmZNvzA6SNAWnUHecN1l8l5fWYnTO8
A8R8FYlkHeSek8nn2uZmGL+oMMhdxfyH/45JkHN/yBmni9UW/uq9zTeb6BDRhuE8
bo/qRC+2leTWNfriJmPBcly0Mh88xP50amwtsUXqdmQirfXpxAxF3po6FT77qCMx
qy3U4pdoO8pTT7Bs0A7l4Ax6JyYlpavsprVDG/MhgO0MFiSQLT6qPtkPSSqQjGSj
BJxZ5iBo5XzJDu8f9/WL5vDplBclvJIMgXolsFJDMaNFA2TUjPWxZk2IijETON68
WnzlnzTVTNrf9e38Z41379wOt4J0yPkPMLguMNgSCZWxY+5PMizligp/syVhL5TV
yp0oHNIMXSXBaZ/JJUVuKI5Wk9AQUzJl23d6EDUxzwoMamKTPvXgc0KpQyWwpH+t
lJ/RIIuN/C6xHjlmD4VdTQ5pYfEfEau5JAHgqBxfEdNABsnXl2p6rbHiaD+4wsnQ
6JtJjCFd49EDKsBA8V60dCgcOqOo9paJnQUKYCor+Bjb9ZarqcUxSD2ZXl/DJkGP
ShcmZQkFs7U0oeENuru36E7Y7CftfUEIYj9CElDfO5M/TVPjoHSrnQ5D/KyVgPr0
SIrn3HvG9btONSiOzcQnnGLuBIjEePBBntxxTThR5ysQsVYFyOo6BfgwSN3iFTc0
59mzKQBA8pKnfAYumLLPKu6dJN0m7snwV/hbqOBlMLRjVRUs3RcMup/W9rGX5bCU
L0noZZLSAs6jULVTZ0pvyu0VeGqwqS1PwnAs6VmOKc2pqGxxoPhVN0cEgDLWsxgA
h581qiJi10dPCz5Ejf5ykoarB9428kk70fo6lEvQtog9xO4f+IByUvEf5hGMYxyH
71hho5Vo83eEEML76IPOpiWRxDglhEzrAmjUA5XpgCOgYPL5p74rbpOcN6tqK9IB
wAKH/YSM+aHr/ZsS4K6lckn+XWNaQ0zb+q9Wyzm4J5taev4DkM4OipXPJAN9eEww
m5irBCncCbckTuFAaV7iY6dPhjF/DG2RZqlwjHvoV3nAkAT9ZnycTSp9GwqiZ9vG
xNuIyjTHMKGFo52+VNM58P+6Ffg2KSqOk8d1/UoaM+WJ9OtpBfElmOWXyXZegPV3
4zYe9J4WBDu8Z6NXyVfZm4R+QxKLRlOpnU8gMapBeqhX+ipPdP3d5rdRv3w/929a
ZyTfnCG3SX2R/GKUjLARbdJNIJnZu75nEI78/z+2D9WBSS7RATp7y8H79pterGNU
QiRs1gYAwb07s2ErJRSNzRUnQ7t6zt5fsdBBcMkcmeyfp30NWn4y2/42NPZrpjHD
kkkvM1pQ5efoMLaMqsaX1+hQfTnBwJMIKRqhudQBkcE7Zxthk02mgtZWCmrvGUCu
aT20UC5EZDh0uiNuIZ85YVr8f6UTkFHqoBpZv50mfac5AE4WXCcSwzlD2gl1xFRS
YN9wQvXyUb5cqatx2TWOhvbTmyU5SvbvGa0Yov91WQdKasx4qzJBpauQk02dHpOc
X4VFhCMNHOP4rX9UQTRHpcHClsPzdQogxGoBKGY92m8+NCxPUbmcNCeeKGyFzllK
xqrQPMPilkcKzvAKQCKgP9fFIbNB0jDJuojS1P8IqkpiBZaj8jbgkDwzxECEg2bc
BzKW6xqzIENX+a+QGuzJ5qEZWLsSz0ThZDgPiM/u9dBSWJAvvi8lnFkKhqkhzF+y
uMmu712sjfcxNoxSSXLQINeHjjlQfEr7MzpXaOa+CF2mBYNutoDo7zPQs+E/RejL
8eybI4EX6pQdK/UQ0784hVJGllbcjzzfHZfrDlj9h5Nr1VTPKONHeyHDQ11Ehp1J
lK3cqKDraIRZkUn4pEDlggwyW8NXULA/JFJxjCovWhnr1GpCXpcF09xlxyYOWP/d
AW+nt7HgsEYEU+3CEj3tGF71I6ibH5kJNXhrBK+Xrn32hutkS/zIcSqwDhRpP0VQ
BHkdClx7R8M45sMM9z0aF2eQe67prncVioH3YkCUC5Xk4rONr7WN0dFUVTdX0HM7
qdX7f5Cor7oaNtE88TeynL2PWiS3xTvF8ch7PsopNAEMoclknZ1xOBa3IdgTsbzI
org+v9M82zT6ZwNPYz9HR8IuUfd8clEsvUouUl21wINdT/QSyFBHYl+womSwB/TX
UwVAx6h92GaJ7xfbwhQttxK2tP9jR4lgl6wYu4yh1R3GOF0Fr4AQXhThVDnwif0q
qmMYNjntMP9n6lfFPZznFyjVELmJk3FYo07gA5f80D2RAHodHpBNo7VncdnbmNUH
XQI2ZZ71iiTGWroFbz5jZKqG34sdbs3e/32HnODKteK+fyQU6Xu4ZMW5AaO+xO0i
0oHiHL1Ns9auffBJ1IbX8w8JNsJTuvKBTc4pLDZnpHH5q97KLHeepVlJcEFx8xZq
FgKsCf1BXJJ6XQZf1r4YV0z/CmF8Nx5QnRO8CMXMVCzP5CbgHgoLdhahpuzae0b+
BXUgda3G98wC2xXej6a7BAr12B1d+DDvvU0xuh7VxrWLJaM7bUXE+/UBoI38pdfm
f6cfhClcAzsi5dYsBugBC3f1oir9hFfOgVyMlRQdxHDrQu24wUqOGxeDMmqF4VIl
F6wF3hbISwf82Ckd1hxBkXHrdJeify6DtSF1ytlYINcrNXCidRVQgN14Z8EvXxta
yNuN4ogWpMdJhdDIuMH1Sp1KbctxsjA3qgZQj5gTYA/12a/DXpxpDV6LwqstKqgv
UfdDs5wg3eJ8rBGwk6Kwy4aAphJ7krRevSVaY0NmXrLpotsjCZqKXw35EP+82c6U
I5tSvRQbjB2z6hJBEjos3yrIxCcLA94nhbvF4kzdpQZsX4wRGGkKuV5Ykxqt13K0
GFvAc7G/7vx9PihO++yJiRu/lsCjXXDF3xxPALyHqOG5/j3gBZ6QvO3m0IBjq+F7
pAyJ0gme7gIZ8QHE1aKfG4a2X+PqDxN0iXd7M4FCTYmFA0+8Qj+eszpS3NScqbeE
t4zLgTPUh/N2qToCjKd25loo1B5YZRguFu/wshNTj6kOP7C9dXImR93j+2zMgEHu
zMXBM7SNO6M5FFCOqnj5fXG2OmMYBrHygX+xoxvt9BmvRG/i3SWx+d+yB7IA0ZQ9
V09sRTabIa0ljjWOyAXEqOgdCV94peNpN5Ol2h7XaOzvcy9jc8ShDqcXGklAneKv
ycKcmBr/aHA4i2iHXuiiYL2luNDtISEFfEIb27uYlD5AdUMb9fMvvZappCw2c3f5
0WRjP7w+hjEbRXYUyXFDimp70OUGCNRrsUBK0/nmUcRvjJejCOuE/m+WDC1c4cjG
L7mXeMSpSkPRpxJFstkVOtVrAzYoCInp9qIgYRKIKQS41F5dBTBcz4MFBcHRKUaK
3N665P2ZGsJpblmb6njd8UiGxDDrN8PJ34P77hRklCf2ym64QtSYQBG0T22l2pcD
LpVMH8hG9GkMLhw8+pjfigFPf4VVLMG9uNKANqJsoSBqwMDjQhcU5V41taLzLEVe
koTfC495n9TdNukO6kdbzac7WNtBXNLinqLgLg07sElNBj9hBd+IBpRnmFcuGwfJ
lJJWBy/E5AKjKxty6+sYX4k+IfMteXpw1zOULP389dUCYcu6iE/N2nQuZmf6V+3l
ugDyI6ciZaBKjquAFLFyRZUsY+2Oo9WnTDPY4jbrjRyIIUgPswBMnIzlEcqxjuU9
aMClBSP+LR1UI/V73/f3Qf6rhQ2ycBB96Nsvdcp3amQuZhbmcAImpYFNT7mjDnU8
OhIDmL1OLBDtZV8VAa0LNBBb9cX74kgFExKVMC06US1VYCCldRqTEJiaeZqDeppj
FvmOHJxwdk7sbEDJ2KLgMG0J5kFWGDwDJF4fRoDvzshup4K/VFQ4TzZDazf20AX1
0YNZG9Tiw20v4uwCTEdgX8PUruAgeNB+mS8fsn6VRnysIjL3NJFGFjyed780WilN
ofQ3eowjs3YQsI5V9IIgIfhtiMDmi+1u36qQWkH7c3ymYHybZ4/c4eNyr0CADe1l
XtEENlgyx+Au62gKy9wD5ola/9aAoqva6fJ8PbT3MjzabTdLYq5p2BqQE6I9/0Ro
AvAFmpBvGmMoGDI1aK1JceS240B/cNl+GeIKLyEJw7uhpEEp4IUg3F0UaZVEfgVv
/OH2Kkea2QrxGuCjfIQJMA/JRBBGGkVOkLzkYOIPBmN5KKTEZODXM/bmyXfS3RZZ
sljbxlWeRzs6t78g9DuIjpHYuaCxLZaf5KryAMgpYSAkOjlOiuMXxk6pikx4a3qb
d+UO0i3Vr7BrQ/Wd1+c9Uu/7m0ApfYUSsIT7KrzxEkfwSwqz36GQNrRcoKe2PzMF
7JYCkfE/KKNKK3DDWpxtuU+TvNhYTEJtY83gjycn23EQLxAYmYwzUwYXrtXLvCB2
RJqFarv3F+Xge1sH1qtyv0GSfsHrTpTNaeNDeHwfUqfKj65ZvJmAt41aC5sV0MNd
FE5vnJga669malNJfeSpQ2W76spged/hTvo1AF7GNtmPiINkS5J0d7axr4r7Z0Sw
kZoo4Wcof2tJU35ovWdRXqtJBLYWLhQvzqjtUlXLOjDPPVONmESsPC0HDf0dvix1
V3QmPVNjM9pV0OaVrA9jMAPpmmvQ1+Sn94H2kl9QWP13/Dsby/EYKOu2dRtokeVC
i1tQSa8XQHaiF9lPum6UELUdOzbHBdCTQCDyYaR99a9qf/zK4b0GepWyhp+naaZZ
Dc3+hmUkuAUyNA2yEOp3NUnknMYfafZit1POOpNiryWoTyESXXzRzKoMe0NHaauw
Ks0ZfZRL+lMNFbnU8vZpSPy5Gh30wtILs9QNPLzT9wcqF9k3qKVWdS72Gzjqrg0i
2lipP7ibTGUw939vZWKjOMQllbK7f8rorPSiBN6RLOTefkeVxl00slJacGYZHKQo
qoeYptwi1pymu8O45Vz9yIR4qX0xqK0TB9m6J3pEX+ZwPF2Xh05gVYNT9+HqNzPl
WQoBVgaiArNT9rI3rK5zJHWJ71oRKp330W5bKIDeivhK+y+tm877DbLcG59F1xoI
3U99PDmxaxGv0XEciDBJTXrvdNdxtutkZENqx2o1eglFBxEiehQ2Jqt2kYeSxQq8
jpl9BSVUKxjNWg8Jem9hw5/K4lsL8o2Z2BEkF4d4+Mj731NNWgPvbUEvP9L7A4Sa
EFuMwh0WJqYVnsM9X1Lj8VOUjqJB+Tu8/GhVYq3+sfabbOke7dw6CCz62NT5jXHW
P9M+TsnAu6fX1ETMQno+LACsUKD4xb/CuyODX7Jvl9sO+Xp7RngTUBDQHJEzIBTh
2GJrdO+uoTpMcg3muRMSHvbt+eO5a49p2tjAqkGPtOqvppKPOg5nuDuOHYrBoZzj
2kG4HhDmqJdEoj/5YyfUpd7I7egE2dqoQ0GclZpi8KHURWIzkIcMG/ISJBdrXfMq
8QQuWhXnidRYopyvRw1cMEqpn7w7T50TgSjsYrp1qfUWa3/cFzaS6kVn4BIqGNrX
Bp7JZSwew1brHDioG8jo/IUzagEYkRF+O6Jq0sHI+Fz8f+WV4Z3HDtvu8Dt1iK16
8I0hRtNgNQaepjlT9awgZ14m7ADxdnJzmGZi5UxPWWJt+pBfkzf8GKEd5ei8nh3e
skszLsOSwVen6Mzf3QDoxDNQhPrsdFpSAwYM0K9xlKkGpbUHliq8o84/Gf7q5lX5
j9UoBYPvyCY3enUqxaAf9HalqHXeMEr5XqkT8ng+pliQPzh2H9apy7lSmdiXRIw+
geYjOGIMcwbvxFajdKdfbWpVLneoTvjoh+dzJZLOf+WPNyBfXmKyUGSVTq2iOD8m
EeuuaPC0AArsKKVBMHN0OQTrvXAKfpGScfVbB/AZKUYaiXAwJOI8UMTR69skUoe5
aHYHXXb525NxA4uTdu8wT0i/FIcdzsy1d+pUJF3a9vYYrrBNtFVWMLSdGyVKF3U7
fMJzr2HupEyX2VlGS3rkjR82qVaHjVMLw8g1k0hx7hVf4nAexCdFBNIDhJR0F/6M
XBFp5ctgAQeXO2G4qwdp/JFWvYDDSOXbw4LzUhlW/DvpXUvMLcEv9zN+DIpgnvn9
FhBMzrIy8yrjFJvsm0ZsBYK1sd7tuWXhSxs+ofiGHWBDRhvYg1aBwGSbtSW+bomx
Jn2JY+2n1K7k9tWIHinETL6IyCu8260jqOa/XoQykoZTrX0/CwpMiIexmIeI1VJo
jaa4b07kQMNyblsApKHaTtGfhpQZ6Mpu/Uo92I75+jvuJsMpQ6uHr2Allsopxkxs
0vESsYtZg8QuzGjCMLCLIIwtNiP1yUD0TDu0FxHSrBsLqn6TvO3Q7Cg4Gs0gx2yP
7Yi9/MWVgRGhgSOr3M7OIBc+MGQ0KbZ/utMT0goJVbpn77xgQCfHPxY3l3k+zWtP
OBXtl4xmp82hT/ay0130GmGpizCZkI2symxpU0lLRRXsGVB2hrxNVDa/JCs/kH7a
xOEVeUeLQg0tRydV13bQrsAZcoKO5JD8wG0MrtBWz7UcUuciGzwobFJEbO9MPp4c
JOkAAOK/qg15cwbauzbb1sRQrJAUwXWGmdhL+UoBcd9cSlmtCV8QBC41T8EYPk11
9QhkPzlaZqRBVwP3LHF+ADTxvcIVmH9ZYmKwxI0rTLNl/mCDapoYYJv7tBwfktXU
o2V8zdHtUo5qUq5v3cvIEu28J/2tqi/49n53FOlKrAlP96/0Xbg0J4FfVUWQyJMe
639udhp63h/c+tgLelzUXG5dOEFU0dt9tloL3Id9iWg6Ag/bs4xfYZeNNciF9WB3
u07KacCgd0E9DzunaPvl/BJZr1lL2LBvPqNlo27X8m66fdjphdsVx4oBc4gIzgMB
uEI2OTY0WijVW1+hNtJDLHyashEmeOMfZO8JLqfg8mIDFBit6D1bAjTFMEI1MGCk
2HrypsHLppFdashpoTmo+f8ESvp1+iFCZfclHde+SZCLa0f6OW8paBUZoe2iqmOr
9wGAk4+RAFMmCDlcSHKbHMw7xDoKBJE/p57QXjqHdfuioInuZVDtIO+wuqrp5BXE
mqU0Azz4QoZFgakyDD3+YCn71GEOszZ3UKUB9WADhv7bgSYQ0NRR6tajg9Y8lSg5
kGOplVa7PmDCcdZbSxuAuhzREv48UpluAMJmtUJk4cajmXUYLTb0N5/KXHlA18R1
gXcFUqk1949DOX/1vfa52uKl82PnAwn5DhoH4nfLTvpbEshgFBrNdUP9tMDZirYm
Tz0PsJgdlWqu41lR3bS7sdI/qsQVzeAYX+JsQYC3oxfQXl5FEGzCctns3Y3J0KQr
GasQD4kNXezeVLCfIUi/jKDVOL1CcVdqJIc+8ShFlzRrswuqJjpXchSeGyJ0BlZ2
ruse1H2tXSz5+u2YdQn0ODc9JzS8ObCUYjbn+T0mPHKreenFwbFBNIl8x8oKycbj
fpDsfS+ifngZP/FGt2dHD7RlJVvAkGtyq4amFpoaowM2ILGLCSsfSswJpZw6FcRW
5UuQl4RkwyITvtDACqBizeDrbThs1WfGXNyBJhrAhF9stHt63t7dmXGIpIWiVfX2
4FKXhyOPjANCYBF1Xsd97PFdip/CP17SL8+9BoXPIjDg/cdFyBf2P7vfnzhgRrNn
uodkYYpbxqX4a1dVyG6HXYOyizSg3oR6nMAFsX1ntCdgEbbZhqixYcWfUbiLkzGF
SrDDWwtXLc3Rz4eEdyGa7RDbAmn0jsbrzLUJWDAt1pVlw9+xvjLG+xgQ6iNVVwjt
FUFfrQwbrf37tx8lzTx8qWsk0YVtAE1u/TDU1MF4BTJx5ePRPdbxlHUwuF5+MEkG
HpVpgPJs9UaJBmDOm7Ihg5KSYBX3xb48P/US1d7lHMjfbJyOHamerY/nhO5JvgHX
LPM0TWbCMD5qj6//QmEPRs7Z5sIQteD7jMwdDfdUEf9vPJwbBKhIdsZCs4CSJDpT
wiDR2fY24hAutPHNJaxTl4zXVdp3MzhpZkYx5j25Is2BCGEdJ4fj9AmcYWlyYwwM
3hN9CrlD4H9N4PXa8nXxrgX/MFtAEil8ZO9vxD86qZ7X/vZc54DiiLNkLfHSKv7m
Voh1TCsLcYxBO3vfVlEvCUY57ezNd+FI3F473OkIwnBp9s/nqI9hHhklG/6BNPW1
dNj2sihfXUoDPC01rdMGS3hb4/U03psrYQ0mLG5yPlr6laiTtXCQvCreaGRHPvH7
8XmlY5RcnfVveRITeEheTqRSJaAegKAYhy8bx/yc5YVaqYRHSYYiCDpATu/2t1GJ
X89Lwb+pKkW+op88QdN4iVJFjlf8TctF30rfsk4JOERhPrWrssMXB7mvHNGPWdPK
jQx/v/BgorfBvfW48PT0AbDkP4iKMIs2vlOE4dwwl+l9123oqA/YFSqAFjp5e7kR
qRMTNiV+K66GjxeQnDJUfpAnut/b1+oP3WmTB2JC+LX2pqMJsQGWukKrBNUE5MD+
wQSrURg0w14A91z71b2QPrM+rFnw7MpwPy0JYPb8WLIaHRC04YUWK878F0LM1qZD
hAtzLdcb5zDw+7KltiKp1Nsk+oqzuKpTKo+lgCpyThWhxoNfGmN/pu6u1l2U+opb
fhhgrz+OfnXZjUFkO2IBMrBKD3v5GQYI/tCbB+fGp5oJyIvIsZqoTcBnIPum9NpV
Vrm/qyEUjSL5rWwAol2CcqYRJRS9anT+FezDyw59S/DekAO1Yti2xJQiD75ilFGr
8I+oD1+xe9VA9X7sa056jMAJ8pGqsPQ6vpD7XJq7+kmIqvj7B3Lo8mk+g1DCdkaJ
0NdgwZPMcXjT8aQ9nkydT+a/hkXQbyXorCAvVrE15bNn/ee0naNyDjFG+/LkIIBI
DpQfgt78xpy8Pxd1d0ALa97rQYcZjS8zXq7AczZZS7fCM2pWCtPCfpZGU1sOOJwX
bKaeU5nu/bpzIkvb0UbJOQHlPobu/kBrp+vJPBfb4O+86LBhkOUuuuW/mrKBRGWh
8v7IYuDYbqbMgAJymu3ko0SvCA163c0JqsrH3ERpHxkx97ZzzK3ynHFtx5QfJpU5
fpl3O3ci3+9GYevlmR6fA+X27TA4lfynMCuChbkKxW2xXcWZN/6xDXwJAyj+7NmA
dujtfUD/gDc34sMdBso/VJdvgdTJ/k/1B8pSiBeaTLHjSQV6L0AyoXQvlLIskJuh
hHnBn26EL7n+gMvxWY/NkcDz2BvkkmPO6I2lbKxNDR3P7NXwXc3qNCeurhpSXStc
+IKnwluGdlv1k99gwcAQ2MiWTHzUKwQDULS7VjByZ4c8TDth3Qflx3LLOYpSxL8q
240o47yqfuDIEts5L8NMU4OEr0NlLvMBTfsU+w3b2XeEAMnuHzvWCu9OJYgKI2XY
2LB8J4Q/z4QIVwSjqim4+JxG6wc1/YQKDoLLSJ4ukvP9uwzvdpj1U20CgZdwQZ8S
AGzE+iHb1znmHXTaFWW/jPLKeSfwpAkD4JV9sMKQwKSED4LwKYWWMlEHTGFqCefS
JbYWBtmCbRooczBK2Y/YGnQfMaoBw6o/9emjp21ywnmNSmhNDRB62AwE+SLDcv01
CAE5Ppu470ByY/wQoYOivCen4IT52h+rthj55hQjvTx6c+dF8LHpjaIAsilf9YyO
s2YTyckhcIrqlDsXOii8VWb4ELoJooH+Hto2d7NflgBMNf1J5efg1/3bMWHIazrW
tKYop//Xp3IO1djs3CsEz+CHeYEtnZXaUrW2Odub6q037I7FLBeYgfnB4+irh2oH
V2Pv+AVmj255TgBQpU0k7zhNFVoypCoFU76bV784KWFNXLltOYuzSYdeNmCaIyHr
pKz98Z3wuKo+jvyYiepJQBqmGV5attXuRsdEXROHfWnAZH6iO+fMz8xd3Dm55LHP
YoQuiBVDUGgfLM2Zx8B/5gXzmW/M3p/403DX9VxfEx33oEToBtAhDhk3D43CBLOO
TbEtM1qGx2z80po16EqhvTyJRR10ZvItcWroX2o8aGPm46uIBPUHO6BNr4kgwIh0
FX3h+uTjQEp9rk4roIxnkQUOPr/9b/k0Tg1H1vo1avdZ/+xVV1ZOePVmOLGuGK0c
UfZU1AB6WTZa6xNPxI8zNCyVHAH3tm1jX1FRVmWc/oLBJJrnIevwR6aXhvFBcw0m
VVft1jco0UTCuwDTF167XVSEQ1BKG1QxA90ntuDQJ3qwog1QTQplBcEnMoAop4au
FP8E9U/x3c/WosvnPYWqxr16BEoAd9Js3R/brqHkHvNRmQIm1xE+unvLf6+G6O7D
WPXLn1G5CpJbtfZMZmuJ+Itii57qR5fkEvCxsLLsLqtezd0x4XAWQr/R15cM0C4E
dgM2HHdP5hifuMnL9C2nLqWgWCruYoEX2zKWTY/SJVoxjwDawI/0ksZ5vFt48I5Q
VHERJYgtq7nlpqSV5fUc0CGWU2wTlxzldjxo1oQ0H5CBUAh08rjaVCvNLkMEyWy7
0AzgJsWqhh/XCI9iiiElR9Pvymm+oyOeqM5jt9lvAf5OlEVKR21ogNwurWnD5Py5
fX/JsBfRVQebLkQKuZG0PUOZCoDaKCfUfQ2vz8VzCJbjotlsskMqnDnAmcBpFyeS
S86bSr41UBTLKJz3aY3rWeB+0o5cHaPZiVIxXhS871Lts+/nAUsNvx1N6h3jr0A4
nK2bTH0p4FfKswpKRd7x474gtvcuCvpUmSxOBirHm8DEip2W/ZXXLetiLWLyXmHP
EUuepdFTTHRmHfhJB9CMdWIA3ubhYtvOaj+p4cMeymDt9PzMo3f8amRuhQoHemPQ
xgIIvFYKsZ1Uq+17mumft/0zSwZTCIDa/hBO4cGPZ2MlaBGdYFAwwiPm0BLAanPt
iKeUjk58QemtEYOj62thUlYEfgVw2x8Lv/xziLzX72IwR5klmvBAx0JRyIcaK/ew
Q/ej7GM0fBgKSvfGFaAxvoRtswiCrDSeEYMnLKJgTqUtUN6kHSJ989u4AOmoWr07
OZw45xAXqMFEkMwLL+EiIodx3LtqyVV+KU4npBeP8ZdXE3Bryz04+nl/9ZZoJ5Rh
NLiY6CNjUqWVBNcIVy65yJjRWQv76mHK3OrO+ruVDE45Pso0d3K33CYwI66rtqzE
ANT+YWx1o5QMlMLohvOE07+zuTGRV389yqviAZy8I8RAYHNC5QAUbloGoc9fNueF
zi01VhqwyvK5pHXGYRfp023Yk1WzAF4F2B249zOODJF03LeOYwJIxfjTGWZu0y//
kau/YxiKoYu9sG8i/ANNP/7/Qq7QNSkSE5cmpzDK2Vc2ef2++ZwrO6cA0TwTUZDK
DYtHILbDsLwXSt8IHKGJb0EQulmr1CnczRtHM021F5F+fDyF6NZyNdKQOb65qct5
4SM2FQJgms5SZX4InaHMwkJkQLhDa5z5fDmjbcccPwQIiyyV/QPo+4qAgUCa1ksY
fGiuyXnAKxpFKXlBUiCreDkSWQqeFcOfyJ5cmx3mErSdpdD55+rNg3TYT36xig4f
VZAjjhbtRyARoXNTwmaV+02G19KE2Mqia+Z3IeoPijFhKwGRl6geiyZpVJMVmuZc
liVwLHKlqPYcMkS02n9Wr5JgZSeLoYTHcDgBJRFTErr3RwR0sUiZRL0JyQwXNQ3s
y5rlYwmb422IC7Hf2CrVg1MPISK27oK7rQVw19NaA/Afl5nlXigszChJ25g8jATZ
EMH5MMXtQHuxZM7dxVgwVqm82QK25IiGjN63A6/L51EuCYAiM2ku1NMXQnOtbUk2
JHqKIazaO5IZ9WJ1b2bPQWzYF5tOOxqmq2i9UEFYuCz483Rkl913jzEOQvLZ5yyy
R6hjF6aVYcfjBwd0tWG0Sigqg5efgNNWDqaJFrHYy1NE1nIlt4GA50DtUU3lsaON
wRWiAUTrz8nDP+8TbvlsVPB3OqjbSNDEX89LDerimf5XgJwg4ujEaq0Wm7OixM4f
4QUxVE153v26c0gOtyhjvhQdr1HHADngOCqqPgXAxPkZ2jfULWPTFvNtUW4WGt8O
nWLOgM4ubIy1fSfNXh6+YpLZvGvib1xnvX2gORM+O0HNVbDPMLr7tk0fONLvSkIN
YTVL/hU45ghm52xRQYDakYPg19O4E6G1woF6R05gvJn9OyPo/tk6RR5gQ9p20SU0
tkqDoxL1qtTDs1Qj2fM/+yInJXHqn15SY6379bDzGntGMFvXTIu4tjuMuml9pMWF
VP2SOw7SRm7leJsiuzGnzX8XQgPgPL31LH7khEVjTsUlM6BaxxT5RC8FJ0UCDOtH
StMsUk0I3TJt4MFgvsBKUtM+hju8HW9MSwjPHu27SO0oPdDIzNsaagJQI4j8Bc/I
5uoBt/M42YZjlqBjd+HaSzhU7o3ZXDWr/2HgNFLThvHE0xljl2ft0x4n81b7vPEi
8BfGMZwmLJi8na4PQJEyJ6KmhFW9fXNZoSOl8ihfF1UBnv4jWQ4AGPGIjldbgYmi
2PAFcQuzpkpR0GSRIdQt5/aMaLcWNeUfoybuwCnmjx2s7GTam7ZF/+Kli0QScep1
IMYhJh5hyP+uYCe4zAdE+D7P5wadKo74LSKTdtfm20uZh8ptuZO78HPRavyZDB4T
OpWrKIS0BviyuvSl1IPLf3kXvUY7ZGhoGgrH1MZhqEBMAdVBnn3SFBPIb8xltQr3
+Sn//7/q6lTXYP74NHz6Gf3ymylaPfe63f0/5RahWCFNOcrhGJaVftgtMI2M6zqj
bjdIWtpFjGCSZa1ijoGeHdNx5NiR2mc4gZW5vb6huqynQCQrIIT+jbPmvR30B7qp
xO14EHy7/h3rxvW21K7z3y7yY3qm4TK/flKfHndJIGPn/IxmQ4ULucHXn0RWxpt5
EaStF+AZI3w5d/nK+Qz2lJBmrQ4u+TTdbiP0cNYBsCAJ4JR3oZ6PseCBcRqWdyXH
ldqwP/N4OEPXe9Kamya/ssUlM4uRx6vMXsgYZC3HviED1gjWJAseWHQdkdsKUJGQ
IHHIivXZkf4TPmzImx8YPg9dGRLkWIkDZ0UtI8JiQcUzBYqEg7LwkpqkB7qg4iYZ
GQG276JDlvj0+JJ7g5y966jS8N54c1yVNcr97/E1w3Esog/91Jwuygf7QSbrDjam
rqwVhLPhgp44w4K1BdC5EEZBtgVJXt3/UuBBLfypMzvJa2j38fbvt4R+OB0Oht0r
WzIpVW1R8xZFMcecZGygQcL9sC5ibKB8Uz92dJIIqKErjkdrmJroDcn6/VfF8u7K
7MwsOQFrmmqBIp1H675LRknDi+kpnXvV7yL4FSIAcSxqa5ZHWSoNq1THJ8xUe0rN
AcEz1l7GcswIJwksK6boGtqbueMCk4aiOT/UeR/da3HABHydOg7/ZqwGIvXMZ7OF
uVIF7RVWJ/xaba151lhAxpckD4IlkYPvLzvXiZjoXHixffHVm08WmyfhVGk9GJaF
9W480WUHdgUWXTXr0cRvt21htObDCxWr2vMosHGv6a0gFv4Ey7bBlHlX1qOLbI5x
K8jgj6lPr05BHUTYgWTv4FKgnc3bmBPrqKiwIJQu1mOOIa+5UB4d/g0ddidUO1YG
8AZq+vPfj8+YfiojX1h9ClDYtw3w25QH0Hz1C6S0Wzz/rZWuF8B+hgOb0lSXgCQu
O+sOVyXKDdckN68TmfyrAEAg+Zf8x9iUszUtKN+7hcydve/wI/ffou1bM/LKLkpC
qdJzjYZ+3RDje24WWzl5wi63SVeUdrZq6TLpRLQCk9BslrMsM2LhB4UDvnh37bnf
cfU6T3yRf7u8f5badhW3E83OmiTBPWR8Aa/6EYUDucfV0pd0Tjk769ah57zNmOMb
n2K7tbynPRe56/U3X1Wg7qRrXWt82cR1P0W61nwCkK8O0BKqTJBalzMi7bMJQXLF
CBekwSe5tn55JLQWmAKWdNQAlDFF/nWEdqMvJaWsPCCYuUo0KELOhlZLc6CPh0wG
/gfuJ6J0pH+VofuepyMvM2xbjSK1DQDxZF0lxIgWCqeQJuNark0JjJd+9QjRSbqc
WfTBFKu/OttUo8e6BVVso9vYbP0W9DjY6uPP+fm5fYl77fiXMC0AWqZw0HZz17PC
CzmOIG9q6yUPBDlQU5alYvMS6CtYz/7yB3VV1bQxt4N/UCfkbJNqZq3zT26Plx80
YW31BOsBbi1CP6k3yT0+WZqZzKze7OeLHl495ewqQ+t+fuCJwIEFYf7OiTgvdEYQ
wX+eOi5cfV83q3fB2Tio3ci9qVu/8+FswXwfIFzoyGilto30YRq1HURwd0YS9DHl
4qP9XxGveGodsiT0+DaxLMO3k/YzR9T1AbR9cJvnKRTB4OggfS057USP2n//tZ4t
B94AQBnMCrNPhSjBeMZEnlu+6s9tUaUj1mn+u1hAd9Rof/PaFNMybu8Jf2HVVGN9
YDyrO1MVXeXSqTgWdtISXAZti/PobQym/QLsD4oM4B3izYc5oc7ardFUymJ0AUes
/u3F3GyyPew0CZ/SRmkGZxZUL+l6sFoxegCQ44RzJTFfTQ7UXr5oarn4T7QGYTxl
7ZoSsIWQ4T7Ia88MzQ8lcP6IbWaiFHR85U3ebs6SOiN9vwjNnS+vz98aMGkHBpjD
0fk+46vdH237vRJrCU3tbHQCZzXciwxh3o9JkWpd7EceJQM1to/nN0A2V6ZjSa9T
NDHXeg6MO0jg7LCpBHRb9d6jWda+2MJzYtNuGkAM/HNCVU0o2RF/DLj/imhReos1
pwl8bS1Ui5lE2WBB65owvigl3bgxSG+/wdT9hAIgiIHfZR03UhtVgz9dmIf0Msaq
4tfGya/BvmARniMKqNpgqXZDh17K4mWuAj/0TRuygJfozpj0OhqZASleFUCPxxO4
ZQMhJYAm1gg8OyV0EZ9WkZXXyZC91SEoSi447eEJj4d7TQaj4HpXjW2q6t6S8kEn
9Ea2YR478tWj3GLUCyBh3JMHVDUqKoIL1qS2iuNpXJqsJFoyp3fjmVZ4mDBi0uFX
u2LLIFPL12g++8JDU9mdNzJFxEmdh+LGvR87/Ud5IktejEzvZJeQPDDE86fijAP4
8xVjjfp3uNBPv8SIqcGrE3bHrwPDAhtyUbMWMHrDJvIs+AmD/jeb+yLGntFK0SOd
Hd/9W7DKgrV9xajRm4HFWcuJPgisblPr1aujR5oppV6BJGZ1qvhMgQmnzdqX34PV
XKP8rv8ze0u5uCddB7m/noexVIi11ZOfrvCfA6jnh2WjA6b56SKEmtLtLWm64chy
9m7S01P/iIiw0KA2Qr1Drr+yRhoxAeErMt4D9wDCdf5oEhDgJpOd1UbB0ZjoFT0v
qhKINUZ/CyC3UgIMLwJxQiI1be/MRvhDZOJ8uQeG5HboBoQq9beC1iCGRD9q9AhW
/Ch0Q1scm/ChNzxQUNCFPpan5Ryz6UiJgz/xoL+qA4kCCM1w+lJBrj1P9sTDwEmp
rLksStuJsJfWHyw1syA2o3y2YCUIaJFF47O7COPAlmLyKa/Ut9cOqHiFGIRJr89g
9MSOSlWsjuNcidNQZPN74H5MyOqwrBmtwxmxob3oZZMS5mObWh2n/b5Gd75heaFF
sq8XdYpwSNgW4rjE0Z8WsssSAJD3AGQM5mfHtbe0mKcFBZvbumFufK2dSxJPQWkT
qYJE/h8Kjv7IGCBBDX4F6K0kbQMDb+wjqHztVbW/8wNBUnNZvrkZ9CktAkhtgP8q
K5b+ChmKOtA156POnPMDTEc9SZ8yBB6Q5f1lwJsywI6rdDpcaHMlmgnSHn2HIj6b
FYrd4fjzZBCjjS5ahbi5lzqSyo3h0qjXynNBQs6+VTWH6rx8e8T2pHsBV+W2rL9y
Wcd0yKKEIwu/Nqr9fZ5cyRM87R0859AXValgK8fffY3QOL12UDgAJr2HmD6WE2OI
Yw/gxxt7HfzsOPPpoUSNrIvDDY+jIFaQXEABmsfmkJsfSKB4WELj74Fx1OgaIrrg
8WvRe1Hor7kG4ult0olWR/DsHoF/kEHTLHdh7Glh/mYBqNVFFs2q6juulQaqhpT6
XalRPwIHTkp7opkJFgCSBA939R8QEcFv8y1i3KYrvBGaCDClqek43MI91f+BmJUU
p8OOKVOx+7KXI3Z/OzyhME2fzOj1QsfLoxfy+LGiqhIQgdVX5Civ9NcoOgeohBES
ukiEtu28zWOw8zkKyN2Jwc8jV2zZS3ozeAk6btJaBJ9D8wO03h2EGUD+KosV8GVN
pz9y4YtCuofDEA09j38025O94zqyuS6QIqu6F9PPJqcrQUIeVD8Etv7eonjwma8d
95PHK+W7Zklgd0Xz07TsDfjM+6SduTlyTUcTolnCD02hsYvT5/abzHUFVsNmFqVy
V3pkKp0YQm/fGjf4zX42ukciWiVNUYEFmcgY59pAlAzUpotmjBrw9FqxPAL1HtL0
ElF9opC2xldq8SYE6RoBLO7ElaOtClP043xsYSb5BDc4GqDeIJdPA6Br/MoK/hnr
qCxgqVi1tPaFLBUwT3fLj/jOoBcza0JfRR0BEY5S5MGltX1ycfXFR96K1EgTCewe
DT8ke1IfmeB+TEYtTYgS5R4nS89bIASDaY6vNLqZVKmOKvprISnQPMWhqh6EkkHm
yjIlik+ShS6yyOmNM2YEqODkGojQOkSUZHPhUga0OFj1t4ESdL7GRkM3PJhG7+zZ
9RLyis9xbL6vkgd2o8lDX66mGNqdw7PRpiHmJyCAruX0h4v8I/CpV6zIElP3cjib
LP1ks0J/3UZlgdkgO0uaYdokQeQuS59P7MF7axJC1XXdu3oIwBuhkstfvEAoMpjM
23BQV2DZBZGbw+FRzax2H1CW8TZlWlb0Vkw3qM8clIn6hBRsnzjU0GBc+ULO4+l1
4nishFG9SEsAdSKlSuThfnKG5zJY1Oul59rgq+B/aNNp5xdTiFB1opBMfwmuZ5a0
yF1UTva92rtXn9RoK/rDZTSx3ov6bAGFVw/YLgRYOGdvuJUrh0xQDpOHFIu+/7uz
1kAokOTX5/WCV4+rtjSAiQyq8Y5+sx+vX0gcyhaTcraeaTWfq4xi1ugPc2kxmZQE
DfncUTngvBnTwiwbd/mcqwshTkYBxpvOvP5hQQowzgp4TM9q8fXv0vEL3rMWerEV
hMEXqP3zUIGs3LDEmD/oNW7Sf8FTKF+Ghzw7CyjDEbvqq0f9nV1S68VMKr2FvtGi
Mc0TIiVrzpCY4SlJk6IF5XwM4V+ihtPmi+HfzaAmJrG/cNdGaC2MTcwWaMkZ7Tx4
EpExOP4JQdjC7fACg1/z4oQFjEynFN3IZpLQLi/fjDBbG6kXKSmxcpEFNLi7dQGI
6v6BM6wvBigsWgX7lPEOpIIelwW24JJ7PcNO40zYpLd5ZihkcFhCQwu3muAUDjch
nlB4BnvtpKzm0Gj6EO08yvy7y+Kygsd+1EgLKj2jvyVXHi6Xd/WNa+OPaJV895El
9Srg+VlrGqJh7frl/9B1mz/FjHW2f3qr50zBXrBU+FigMY1P22ST3XDJk5BW4t22
YdQxljv5AazueYatetuUwpJmeGglzdr+p19rIAZ7IZxe4u0mrVk5V0gGSGG5ZW3f
FDHm9QZcnNnI/5PeFDs/JGL82n4TMIRcw+SpDWHT87qX68E9ytNh7ft9T+FuWBlg
9N+8Y5Z9whcl2fEe9XvyFlrhzZ9YFKF2uIka2bIQE7yHRAti3ttaFVkjrErneg0E
Uhi2l4HIOYQLGeDCeVEnzMphNBvg/4Mjl/cfENPTY6y579NEF2rxxtica//MlTfM
1tqP3rOtQlUnDAv1aHNfOcR/hSgNwYa6Mgdjt15WMTaiinuAuJRcuyVRN+xxk7PM
6AQMLB7xsoI0c3GehwjAqVIITYJyN/RZO8lPahfvJyM2pKcipTDP7YHtnlw+0cEl
fuUYOfdXkJZKkGldU5QQEv6W78n0XyzXA+VfjgndVrMx/LP0ZFTnPBR3PuwD/4VA
zevcFrsb2vOkhaoU5rQ3gBPK1Ec7M+uku1vPe6t9fv6sdA9CrkdmJqiEGRC191MI
XKjqlHY7m+s2L0qIcY07GFK8wvA4kbdSarYOwzzxptndJXdim+VMfJtiQI87ExW0
A6vmlJpDMmp+fdzy2Q7/it5xYfBk+gH3Bv4WhD7eTy3k+vrxpJWc+TEiqGFZ8OnK
p0sQbzHkWndWdv6JtR9V2S5HT06TppAtbYrYAfgz3owBa1IQP6cXEYTUJ//Hh9U5
UdWMmXlpOqc+PHOTCp2nhbtC+I7Hkvpsc+PKVdNiQ9Rh4aQhNv9W+sTwrgBNiYhq
h00Amef2D827TN16js9PBId8EOcKG1dJABW26uDBh1hMYebVQhGPcui1hAxWU4pn
k8V2ZlAcb/gwVjPDRLBX3EbKf3Wt6KJ9adv01gXZES5msFI7YjLbtXmn9AHp88Lo
bNf8mmcidfXo7bpLcNM7q9kBK8bEqRjih995ADoiIJh09oy14k+vBwwzTstWQKuS
XrsS5ide6x+Lla1SyTlumrugh5Hcw/jBsZ9LqNAXs5bvEitHK5xX/P0tOcScT0Gw
KruKatwL19HRGeZC4NjszfZ31PPElI/OaV7Kb9rRvlBut8ojSGx5MP3T0oGxwSQt
UTU2/PmFNgBpEDaZOgxhKv7cxScGbL+fWZs58EuqOYQSOti8NuMvGdnzM/TST+ph
ElILWqYQye35mr8ktnLQbeu9iyp4CbTOBETpxhW/PVEnPIQGmHQSVJVnVH7YvyfN
a9J234OI1fi0XF1BSM9Dz+8WYh8Hcu//d9ZKD1fxWWsVvhpH0osb3cvR8a0eiK8v
9mNNearnSO6xOqs8pmeDrt8xudPNROK95L5Lj/1+ZM5NcTgpnYbkWPiwfBK225MK
te+FBLNDvq/HCgkbno+rDVTKvlAlCsp4htvlxBc/ohuiF6/KE9bVZxbMy+5JUbcN
aBffiyiH46u3cqE9NdKtJ7/bPCLJdwB7ckV3SQez4e7FYvX+u3ej8N5+KEQe7Efy
YoWV8BnhaJfCr662pCK5VFFxkYJs4xmoQpxzC//BwEEc5VA6/V0SKS/fZUqC2laS
ocf6XcLrYgzk+udqn+qr4A2XWB2ueKhNQAyE9YCdbrwxAofllBenlyCUiymijQwe
tAETkmTQftBpZvK/x0f1C7py7LfYKns84gwGPkO2SeKhyPDQ0TGcl1L5uDvKmBno
cJhpo1HDPrqcm69gPiEyH2DGDZdVYRD5wZFuupEdVYCWHZsGerRjh5mXZ44ssUrW
fRUU+L0Zkife2T3V6GUBR0Y4I2oljgPaseMRyQuFd4jEW+U57tKaNJ60xZ1E2E1X
hgPEfe7/Wr7KynDq8YRKXzt7H16GBLZEwgLqu2PIT/tW0P8vZqmzEEmxLYUJrRsI
3fTy+Q/NuUOLdTLpnAZpH5aw1KFk0e+sTT8cQ1gT8kDCM2jERm7IEDkosFUp1JKM
Ry+1RcxGVMaOP8wyU3H4t3XcJd/sswIgokV9LosaC5W6Bz0ubHrA56LM4Jubmsie
IjxlB+3PsWM9u5XPPBzZJWP1uGte0K/qouV7nqOIbGwUHGfdIiCGutkEW+IzKXf4
KUwfwYuoaFpncqWLm5v9zckthClGxN5/T6GLpyAtRBWPBAqZt27Go4itkyYWaGbo
oONcvnyy3gpN6ZDTUgYcL0y+aykFWYTi8GUW7UdwfESUjaIaH7SBcZwpwwf2J9O9
ojoXAd/F9N2/ICXdRij1fnQysrOgT1uFGJ4XS7IWrwRfBbvi8r8Hz7WSNcpnBk7N
PWwxshxfyZgQvVbxSwDIT1Pw1YdGEIPWcfEcRLTlmQqDumMzCmlwXOZue6Bf5UAH
79xmilmndWj4sbhTvteDVaJ5EPeq+obb3zp9ljAMRq+5gl/PL7s4KaaJg82FG5lE
6hUH1TZV8QqhCnxkERLI2AcKNKOXb24Noj9EgbNLX7Jm7qnW4JUswC1kqa08cCwu
pJ2XzBLl0K22lmPC7+gvABKwm0Vxg3JyDhqS6ke6Q1Z3af9cHD/m/TDYYtUztGGI
bh5lGK3atL68CxfD9K4VykZ/ArcVcns7C1gYPJOPB9ylE7QQyb0nlQZr7Lr6ipaP
aU/ZfeXlHRXrrP+i5u2qmkoRFMc7SiDiYcvJWau0ACesbGuE+1IZViS+tj2Rl9X7
VYX418PfsNy7iCb01fcrptZYUuNueriGQSXNciIbB/VmPoRv6nKgOtSovPMM4TSf
0FyAaq+Nj6C4l8O0GN0P8dH6u7ILjbJk5ozuz7ImvQiPXR9cAqzT24AMTeAzYzSl
vwTuXmtAavdoRkYpMyLCTbYsE2gUU5tCzRhibjbUt1ewVnjoPlDvqbETWifI051R
JDvmctz2Z4+dTqfeMdeCmq3fOVl41pR3qcMN5/G8Jn6A1opbyuXqy1KMnjkpRQFD
Hc5jYmDqfEUcFRJzZC2RNdpdGcnNkI9KnV0lqoe4Z4/lE9jk4Fmzo3xwWOSitVLQ
mkcwueY6dtUogFcbes2n9QXGymY0UERPsScyUCOlaslyh0Vqw3QeZM2XAOxqgGm9
H5g9a2loBGOdGNS1sRMMCOhJCaRMp1lwTohsNXUex44keBQ6JcNB3R/YUCU0nNaz
zNCdQRXYPvSsL85ywVpC5OaKKSGB7Eu8qBdzEiQH5HeCUUOdfLM7OdxvShmaX2C+
fCEmLWgBa4FJD8ZFeqlfv9oLBXXTwJjtVcbf7ffgil090jPs47bi20rD8eu79ImK
M2N9MvfHSSemm2bxOp1oNgBvBLRc1/YuYksTUv9tr5kHj+V28caH3pN3ialxSjd0
Suk5aZOyDyDpsFsZ7QGHfTot5cKl4n4iYnJ5T9KeROdQ4eegCKejk1Snumvn0SuI
PIjaC5eGqVDTheTqz/hBgjuMJ6FfZYX3ujazMr6pN7sLmxFNPH6+ra8CpjwxNa53
JhzFk7FCSElRhmoyeC5RAcsurvHMBFnxhp41Oq91W/Z5i/yEl8RmUsOZxNxWJO+M
dlT7FnwG7Knyvff62FlmVjRWTpsos3kudt7ripOizcEnTVHkLk5UClYLbHqQZKqz
niF2IVl+22J2Gk1yl9Gl+4Z3ahtVAtgdG23HKgRyIzaVNVa/d/awjQQxwsrwgaGJ
dUoFtqAW1+tvgg1V2Q3GB7Wx4/cg2Cz5276oecVo0VOQdyocxNomRCk4Qiaxf+8E
qMgtKjdU7NOaPcqdzB/dSaugvtK/qNCIoVHY82Tid24tLfz0XhVNIq4vvReEetD6
YGLQXOPaWeuAaqaOBH8eND6sPg8USb/qTZRLUaZPHj7H/b4DRk7nEJziwN4Sgu2H
2JaxNdWfCcEf3A9vzdD0bRw10VbUSJeB75X7913uHPgYzSN983CpKH/r7J2lSAcl
xUTuqgrktCaIEKhaW3EPu8c6AdFxxluLV/2ra2ZlXqX6mxcwt5Ds4LB0rfZZXMjP
2RPpotTvzasY7Vi2SiQI1cShvWJ9tr0lSvKJ+Xqflav3dmUOJpJ/c4oECfdQpyQN
oRHI4FXAyk7SaEonMzxjVgvt/niUDcNGBAjn0IJ5SStnUa219VTQ/tPkUkWAxKfJ
yvyb4xDyXZdj3ZCpdIrhXgZ82MQfezxVPlWTiCsjiGY4ZTivC+ZbJmHFACh0zV0+
eRG2RQ6sO4RjgU9umfpvfYlY2DeVMYoPF7vF7B9DqH5+tgNANUzi4CMHW2FcV4rF
pC+yHQT25rnbQd5Mp2tloTOetGt00oI9VRtqC6ZuvF4OETmfmjLs5HFh0ygYij1E
jbe2I1kVwH7fJb3vtdZQz6Fg/UhV7YhbgOcipeJ7YNLQJrCsmBuMPBoxo6wD7rtR
DQWHH49HMWCFuew8LGh2pYkPyq2UJ84WhnkoIUqX84zkdunmP31eDCxYnOu6eXMr
NiLOnRnBqHEJUrxNqIxM84LO7zEKkQ8g73SmFBPV8A8f57rqPisqeSKdQhSUSp36
Qf4kvXjRXfeOhHph+THml1PgZe5M1vqRe9GV6/4B/yJoUBMSXAvXTEd4ux/r4HRl
eHUNKBTiUdCAfljLfxUgefo60vWwVW0avruV9bPxLVpoiIniXtZoQorEai+1FWrO
UunI+06qLJnj0fNgx5W7Oe1N6wF7NZ8MLRMqKqr0bhEHsKvQPVLpJDuipblVPkXK
rh1ZsjEfaz5jMhlZaKnuPBg1E7jiYTnBjkhWkgBxS5PIEGyYElY/St5qoSlqXjt6
6sY80IlNojcvHkcKPkAF1iPFqjUGCxDlx8Tfs6OMbxO02cw5ImKT/Fgxjl29rF47
2L+sEvxChZ2mqBre9CSSiH4byhVU/c+bnT2DS3K8n873Ke4sOIxdhQVGxs6zJTKH
94yZRPAEPpGnUYX+unMUqd8J3J0lhv2jGEiH+afELTTHSLHxIjvOx5E8+Oxgp84h
Yqf3oPYtgbUxM1RYMp0v6gd3+PR1DqJhXwEsIx9gaZxg5Ypf+RwIJE6Iwh6EyOJ6
lMjpGC/QheidMLuTSYOF3Le5MbDdVy6kNmMNpe4yMpXH06eqiZtjwdYh6Nta8CUZ
LQQBpXOhKtahjcoHt2Lbb/JkPQGurPVHKvDixI6hby5+381a6lTnZkaQdXU/bIQ3
65FL77eTMKrFiFh+unmSbgkKMHQDj1RfEHBGPsoYgnMffJTn/q3t9ieFylKcngYL
6JtKLaqhVfQRgEb5NFrz3tk+IrVK/wwT5//qDMGvALZYvBNC07mdWO2sC01VXXOU
9RHAjphVKSBy+0xRsVIgRcfd7vfUPQy8R3mrA0HaZ38qpNt8M4NFU8/bApqDBp04
XGwaqSF6uJVYD2HXzVP2+Y26BtowFaxjloL5jLx9YzWeiuZHwkKK+LzHbT82y5fG
y0/XcMECwkkw2iQRKavQbFx2ZTyX4nAtBcoHRD893svx+cvDi4lmA3VRcTvJ8KGg
OVz2YM4snFsi5Z9+E6QhJH5G57kd6uPZL/NWcuWNrFsMWkRobVRFXIdQ+wjep7RG
Au3mkrZvc8HFDD+yH8DQWdNaS2EPD52uJMQdYBErosgrIndVB9O0zmJsi5BA0wRy
Vonb8R84seGLED9u0Svfnx/KXMk2NnjhnY9H+SCwoa29qqtCUW4p/Rcfs4ISM/kP
za4Yz/S7N9/15rMjAF6LrPu9lNDBTPBKdmG5Kh4esdKLMBphn1XGifpfXTi0Ad9D
Fm41lRqo0PE4nmVdN5hiBSzAAPLSK7SUG60ZnbxSlHhzJLl7YWtjEm04v9J/lt0f
PIgIqeGDYTyH/8i3WEXR/MF9DCAbd9ZSU6NEpCiTvctXpicHmL7MF3xZbeOtyOYj
fUOUq5mXtNRxJfRO+BkCwEwphM2oAlRT9KTr5U32r/Nezt9Y2NuZuoB8vXUXDFUt
LnDGSx12Gt3NvZlOA30tpvOEmLFS1JdvmHJc2fzZKdmVT5J34IIIBK6ab4RnnJJ2
dmOcKiOUBIhkQVZ0vsHdl6KGeuW8EeA9bW/5rKdbiHGXBf91Zw3ymMYSsRaMi6u8
3mCCs+WuSMgvTYsSj8JQvb3QZQRsS7EIvJQCEyPU39EdcIyfERL9oe2Xd0Mu0y7k
6ogn3m9DXjn+5himfOoLF1pvwLw9aepEiuwWOCz56sDGUgs+4jMt51A4YHKlnyVf
KDS98WQetYDb/kPb5o3x4WofDCPcTtC/z1fEcFkEYoxuBOCM2R1kS3gt8aiFjSeX
l95k0y/viXAxvjmGDFBC6ztkZ5yzVwvKpgCNYJh84P9AoQnhoi5CzepDQoilhW3Q
y7argtyEJjpwd3gI3qINPtGyo+5q1A+QdH/kZe492hIDNHxibAhAqEe4OGts18tv
FPGEXB4wrY1SPHm/O6+VVxNIFUvA3P64Qg2fU5cfhbKTSKMyPHPMmAz49qPhmEOz
+s87e5Vttx8AWZZgtyDmNxUTam2GQsSQ2k8a8Ed/g7k2MdczGge5AlXjNGj5fbbF
cnB0BPp3cDtXcQonuFZ6AufDQDhaNOI/YU3V47BCOGksQ4kWgf4MCvpWZmsUFywd
vOGB317kE7SgI+DSWmnBjdqW9R/yVxuSx6P6wX7RmzdV5Yg1URR030nlc3DcP+rh
/r/sAA1+6QFYlVIzRgCb2axxYaBcCI/1fkwtRzXu8BkLI5KIaCvwa8tPHgu9eoPO
HoSKy2jz2g4pyr1QoPsSa3DcdyEr5Tn5XVf1SPkPc05JyWhSo+o1fXonZVa10KhN
XrhLrW3OIstC9r2BltzxtRmvfl5eIRt4XDy9ZYp1fZPXLFkibUsy8zPFwIk4rusE
SGUIFZVc7vQOSzrO0Qwv7+a63EoOe1RzhhA+CMtVMImQ10HU0rc0sAf2TuzQy1/U
nFapeTRwIIu9McCcDSKA51EJ+fK1clEuNCSe/18H27t/sVTB5xdbFN8HqWQGIQLW
0FYIHD39LgA40TZTDAwf4n6z/WvSOuJ1wIqygDR8jBpO6y2LZ05jDN3qPp17rSkq
DQ7uQF/ACXtTW5jl7rsbAIrkeAzVZIMhikvBxriU6+vNmQJEvCCNfUYCh+tgjEQt
qZ68fE0TbLtpP895GOg3fTEUES8yScs8RmeL083dThc0x11szbE1WxTH7U7rms7n
cKn6Szj0LK9QWEiUijNdZQn3sDGiUu78yQEMNKnN5ywiCH6S3bs1P29xEzrVeRwW
iKVH3coJC//Pcmwt0zQzRc4fmr0IGBffM0xr9waUPhhCmcPtLsle7EjZZwrQDgtu
/3BfAmLDMAG5H4bHgG9Dx/rLlSb9/yhlEJdgM5xhBsrehLxB578WhxYD3637xWes
fEvvYjFO9FlAO7WczA9Hb9D+Q2m7gP2FvlfEQEacMLWCuxk7kWDQLq8xBXK7m9QJ
Ba4V62COuwfCHq0v3/QnIQteKX/SkTOME7XusE4XXDhlB88oahMPLDn8fdNjlCRZ
x0toY/c2Ka20YdGNzbyuCM3M51OuySaoFvN3weXwiCRvaDL+OIFCGG/Pu7GlyqQv
2G7KKnMsdWsMk097pdwT+GFiHcZxVhBMKyD4wi+HmACCoMf354iFkgjW+j6ImRy9
7+UGUQDK4zf1hxtu2i3zwmnDz4c7VsTFfwkJ/gdsGCRV0L/VhOCaV+i5L1IsdYuW
cCRt2vx6+XJV+zEmFPXNzr8wxujwXw74ZDCCTh/1phXRoyqwcPcREMq5ef0LEZAU
TOTdNOmFuVWQTKqUHCevNjJOjPQ4hiuQgSicnAoel/6Ildi0w7wxK3Sj1FbOsDzU
+K7DY5oGRkDzXPJIpvqHSRMLZSDPyF39toqVtTP2o5SNg85uFbf7BeJcWMBGI1dU
rujvy+0TezHPd/otn7YhbF+JwzAMyiRm5YtfCkZIltz1rAYwgmM1BxYvtf+K+IEr
9M7NpaOwUWzgbLT5RyxPNISi6GDbcyhgRoUeCk+pmluYtHXkUCYqTrxNd+9DXg8K
hdX+Zpd2bZuvgDhITw12JyVQ3wz8+D1czSftAOKh6ClgqXHeOeqDpJCBGx+xsXyM
vj2feonTvuA/8kcP6AZtyY5eLUNlGLos5VUEtfTwbY+wc+Cs0c7ijFmL0CdNkAyF
KQJxpLmeZLJUJlkSCs+T+cEIIdMN8qvBsfDi81iL/n/MD8BPdfNpAf+b8zn8jgpn
IlmaeyjxCFrBKsObquLWdEyJSq67UNjYcOh74mqkNB5c1358P0kQMf88ikEGRoad
pRPxoTNFQ0XF+9ixcOqIXDuU+lIFCW/POKYWxZdoPpcWGCNtSIO/vuMZ+B11GD2q
er9nTcNqdNclC9um6f+gO6+wLRMvZIQmU8nRUT6HdHz05lA0eVX4rphJyhHELUIm
y0tFd5SvHl5vwFfXcvVL/uh1elkqIHvQnPLv3xhwjEGKCPK1ggDiVEIYUyQyuno3
GjGhyx1sbVrFxE0ovS56sMeOBuT54+jjgAwkOW62XjIfO7kr9zlcfkkLzLQI8X3T
Vl9QkG/xbWuQeIj3aZook5AliWvPXja4KNOs/aUVLtI9CenrkQf0Wwipno0ePl7h
cXz31tlArEbUb5jITAXiuZn3pu1AFf6O3K1GXhTwQN9rqjT3t8FoOThoAM9DtXJb
Fa3e8Y5t2VvdrzQDMdfDH3YALPrrOFGm/QwRmya1F+5EttA4dfqvCdNaflDvJ7pS
8KR0Btll/JCabTMR+w5RgBU+KlbX+hBeTy/j0Wobb7CV9m8g2A2g7A1b5uon1PWf
iwhUWB3RGvHMmEjdFwukpLCBmyUXSPKHi2Uy5GiLUJvhS+xJu/1fM0Bs3yazHqXr
xumMw3cTaGSseMeG4N2pw1N7ArN3vcIEdZW69S0utfdmEqEOTFnNkvtw6sMU112z
RMXMZqyagpp8nTYhGNncILWqciB2gdiRXw++cFieUQMj4CM/d2Ecmh+gfoURLDTD
Ip/a3mwgcYHasHDR98vfRVR5qtuXwAQ0QW+8zk/CSnau9lRfEKBe0TgiQaItTTZF
m6pkrJQurX0ZIf++STl1kOHaZXi5SwLgTbl/J6r0745oAH39hPxPZHvCdOHCiuCB
gzpV2WsQ9kfDfX+7vxhIUbg2G7qfobcwXQRWEAZ2cdJhEscM2rEuhzGQt4aaE5pj
7hX4BBspQHWmPczMN2PoBKv0hzjWHMd2RoK21wQFSmJ5dyKE01ZljyNOIMCcsoI1
ngpTLn0C183s//C+QblNvI6tAgTt5awMyKjs+RH2dQZD9XpjYbvmqKi/B8e/Tl7M
wbjXZtlWLIWkcLtWHQkCQUMzjEFIMc27Q7c3igIkT5PqLdyVC1N2vzz+ziPUNBNW
nw8306Za+nQmQ+FUq6PBh+muxLKrTvjDm3dz2Dph3h0iOY0IX9mW4CNc7EhjCIxz
mRew+x4Z1qu0/vKUhdse8pHJh4DuUzOBpBwA/HU9C69Pq3gmdaqZa0yLf2wDZwhz
d8aWUZnZsh92r7+uxvBRAdUAgjRgX8+XBqIwYTQpNjfspJHVavSjVab2DyYTwsPE
qK5ZFMix89tuxJZ7Mq77LYOHY5ADOspzBlqwpblHuc6FPMHzPGAxw6qssamuXJWC
5uDmrC4/69FSV9GZ0NL5lgoll7GBqklWWKy67JegkBSLROvkvTIndE2ClWNsOp7F
3bU6DCvfs1xIEwTBfIlx/xptpp7wtfS5fkMTVme7bymnJRMnj/U03qVP5ZAiP5Kp
usVcZ0+n1LlfjRQlkv8j6KoyPKYn0Y8TW1CbpkrDHGqmZXMM6+mzL98839Dv5uce
Q6rHzlmX3alnJfIFiKTAq/HRtKwxKic+f26FvLsZkkuF0xQuYxV8U+29SNIH9t0u
ubR56Nrt9CXkHemP4BHpyLsoCZfR2/l62BtCaseMbRONChOrGibYOhOHvBYFFvPD
ptp9jGbGtLJmrfHzJHm60OB7CA6ABD9f4vtfU9hwuENyTuIpTmKAWR6UvEh42oBN
9JbfU7Aujpuq9R4F1rLYVkcBOnsRX0dTn6qR6K18YZjSa34tNMRclQB3pf6djvie
o8Zj6Q6Khi2IBhysNo+FFrSaPGkMIMjjFSWT49b06p/0qWhfT5z5yclnghSOacsA
orT6mcXRA2XMQf1h94QmYT1YhrftneYZiIq9XA0UkyWuChuIRefkrqa4B5syqV3C
ZtYUFd4jFlKzZV4peJZIY2Jcr+vqEX4zy+F2GCsTmmt2uPvGvy4FdWqPmL4aGh6I
spHzGOCH5BaSc0Da89sWYF+6RHK4Gh+sUPh97VJaxqPhwy4LO2u3ULccDobBkSDK
crdVgZIHNTp7OuV0kSCsrGV056DMQQz4xSS49oIge1wTVb/0bQW+gCOdJycvtWOD
eoTfoXeAYkY8I0HOfnFdG1001UgPbpBWO+a5SWy/EORY7NWKjOrh/EESQB3nGQJP
E2pTEqxqKVxrwakk0QbQQ2xOJ3At+RKxqbkUc1/l7yil6sfHOqCfjYK7ODduieAR
YEpIcrs/fbcMdryMeK1V8qwMA5CCysqoptAIERSuRHxhxtSKt4GQRXoD9AgVQ9zd
ZyoxBfKjbotUUNZcC99EPgENAkOd8lotCYhTIci1sLzZZm33C0V/lWR57uSzllnc
Q4mwE50p/gzc9lH6ewClbndafXPm0wm/7IVI6zJFhi5XHrSwDdfjzDfirJeJqB2I
doksje/+knJ86JOLtYq5ANCparYQlp8igNXrCVwZw5eEktQw1SVuicMvzFmxgeW3
Fx90v1sK23X+MLWH/SzMnZMssLkpQ8AVLZKGgMDsXEN5fa0D2km4mrwkdFQ7U05X
GUlBwEeCVBX/q5xuHbO1VCtSBIdBjQ7PSrdVkCoQYTHeGOpA/C3jdqyK5jwrKEob
dJxKwSLWPjFsodulAtV7zjCKmf1a0XP38RE7GYRoDI7rPjgEC7ZQa4pbPUs5Q92l
c2EYD1NbGEnssVv+ZiB7daD65uQXq70k/x7qH7RoS6iHF5WJfWYjP0y8jzmPyBjE
PdWcYN61WJtuqj4DOJi9RbOjPg/PKQnl3yMDoegr8wGNEZmBoy0wjBW8FcDdsHXE
+PyUeQzh1dMtwNuPg4I4s0AgwTyOBupP7RzHIV8/YBryjFQVHdplE9DEBY5kH+c0
ngHzVgptnCgzDX/fvVNK8RNHJ2WEMP8ys+h14CuFNrImStAGLEpiIxI4CjhQXXiF
dGzieDidFFrIZXOEp7NQCjCUC+6GSHwygdIB9Nt/U7tu32rMLV41Mbfk+zfiZOZB
Ol+Oc/DE7XuQNM45lYMPlFd/+rghBe8N2TpG9yJ5q1cvFI5uFRxDvbHMhHwSOzJs
Bym/OS2N8bbDg2tRXV7jql9uJkZetFB7oQcpk3KX05lPGyqjNxjXss2W0JEx6iZe
y2EolmsAKdhOIcTI2bQeQyGCqVcqDZdB1N3tg0LVlVbGCOuAEiMXnp3kScea2umQ
Qcf8dn/cktrMy8x+mkJ+sd69SMAmkl/E+Ur0KVv5RlrY3QtiluGK5eRL1yKVwoov
UXp7NzAlIK/+G1Et5LbGb+DYiZ+1FKYFe6MeoWTDmk7PQUE+kcatEGPS/YxvchjA
xsiUwOntx3Rih2vdoNCbHPzxHdYeOfjnKpjiXxlDPEA/ckUX9iS3ONH2RB03MZJk
niVkvdmUrCMCLWjs6G1XC8RYU6Nxz+MAEmQfKL0gw1Ij/YPXZZXxEPhOP2BYbZLu
XDg9oxmnuASf+fo1QGOV2P7G/riBCUmHMRt9hz1+hd1lfTI7PElNpNJVDHJGsKP+
eaXoOay3hfxiHG3BTxqEKjEIOabjS2djD1SoUI3L0YBl+tPt2YKUvRx4mI8l7as8
ENT5fo7x38lHSoH2XRnl4gAquMyXX3/Rd0pt8E9FO81RLsvTLNa0p69l+uXP9bzr
DP2K++JDPXoSddOc8p39j7rIyyK6m+wyhSWL4FQ+aD/h+JBLEBomPe5OxLXHkTB1
K0pC1ekFdPkqSmfmDodmb5qfKet4rQyUeOR1mzmmeuYp7/Se5cXf/b1DZDsBEw+K
r1YUW2yZt4om/YbXseMlYS3N766rCzGNAyx7cLLhblVbylWCvCvt4Hu3kObfyPxE
1LyWDFJXZ0mglgF9dol75ejhG/yZo0QaY/x9l6QBLs3H42cPdEuYhu8hAle9jySf
Gz2hTejEig9K37v1xoSQaYriCOrTcpWHjdsJj7QNaMMCn8s0LrUMPmB+vb7orlJ5
UmrBSi2uEKMiC+nJGQekc7HHgl6v5gYfJ+Ag2uRKhZkDWpOdhOMr56l+jZOCh1SD
iki6Yf8UtDpJ2ZW6EywDGD7ipmB9rdFP2/RnKL+K/PvOiDtUIeXnmgOZJt4W/B0A
0xf5+lN+w0VnrpKcgkGFJ/GWQLZnXfyXhieMZ9HNCCyKFlWUsH14elqXsYcHwjjG
pHpYY6mTtgghw/GUNvEVoBuOt7yBBkVHMlMJSlg2pyo6foDoFsmbUd529aXoWTnC
99yu1EGD4jg/L06Ye5HqBEcjQiW0It+DeFVdPMMiCU3UGBasTz++veqa1JaMlK1N
4EPMgK0mizMdhIokS7IdwjlmrL6Leu26lKSCoXD5H/8aS3yTofgetTsuc/r6Z+Jw
bJTtVziZfK2LeMJAw4CBvqGb8GzYjqN341xdM7B6msaQy8LIYKgXOT+L+EJSkQAe
Ve5Biv1FfHfHdGviOZvir7Zs6APODtyA0qt+qDU2yLdrMY6PZJb0KwDa4mmuE/WQ
67P7FuyAscsU3fafxEaJ3PMj8GdGAcw9jTm8iY7Sa3B5JafmNK/3aOI2b8/jeRj6
+5WgAvMG5uAO0u7DKpoFcz+14fBQ+WD11htAOYRQuPsHIkSaFW7aRdF3Ct0Cs4ic
SVWoyxJo2/4ahJFhgGQd2b2gmc+6xMFP329cuBUkr74EH2kg7JwMZLIM0rLUtXLs
V6lOqRdT8KTHx5wYs+w8Qrl+jwzZRc3cFmay4tNej46P2hFN7RVHEXSt9NLZhefU
/cpuTbmPpoURuJPmfIEJSPP9m1jKicr1N7jj/wSyTEh2QmwIeh8yAX9ZMZloy1/p
6tCVtD4tWPlVfS7CeX8A9FoL+L4RD7RDXK6O5HJ+kHUX0Gq9X/TpOgFd3u+tKUtN
b6Ts97jnxxrRisjDTr9R7mrdcn676bJS8SBDmFeCGGFzUOKizkQInyOvBtXKrj0H
YtPGiRc9xRM0z0MQ01r4QFj6BsEcYP9DrTM1Gf0UpMxlt7aAzfs0Dc5SgG8oA1Sw
y3Dw+iGBA48hVrh939vV5NrK+x9vVhm7wGM65hMawT3oLLgqSkQIHRkUBWxthDO7
U4YnN/5Ar638yw+L5rWDouq5GO6QCrLR35nZ+RJKCIf//95FFmaiRpqrNgxQNzqZ
ma2zFVAKrMynCINCbNEXRZ7x+aY+FC7yfpi2uqruSSd54ZVq5RcGB6kVn282qDty
UMU1cpQIlRn5VsCc8lbakE4FAz0lvDhumRxMizRKuJLxACs7EqEETxagQS3vEHZ0
DTu6Tn0c+QGqqUtuMoNKtUgYA6SgkEvEwyfiVIyUR/gCkX2PMv4QlO26zk2WEdF5
9pn+QkIANqvZm7R0tG+F2NtlICECcwwjbuPE9RIloKrtVbRQZPhUbflMPIkgvTpY
fLM/nySzo/7GHSqvzD0MR+hcA44WtDCUaCUxlviGzLKwJSiC5RHdJ4zkX1km8+iT
OfML/VzEow8z7Ccb0oSocpDgAoViyUSFagy5xYO3OlZER0c0Axb5aJw7Q/Mb6QDT
b+VyfdE0GQqBXdci1clnhAvPC7KMkq4exxm0me5rMNeKIERb2c6HxSw4fvVeDfpG
pXk7JLZy0ajo59CPjtM0mevXH5VUq0l9GXfj0pVRLza/IKdB0mN8N6HVev9HIY3K
7UfCG/nPx6cbXu2n+u0n72erkf+KsHAxga7Vbu5ZLHkdGkapvUVaRd2jQ/LCYgtr
B5YGejb0jAdJmbJBCrao0ZwiM0wFZFxJ1ARML6+IrrkmAcqimz1IuwJpnO55jsVM
zI71o0tQA3ei+3jxJ2ypIy/wghBO18C9hg5RqjmV2OFoGbJuO8FTHHH9k8eQgS8E
xztHC26A6HpwVBi4jGfT6C5zOyaRI5bKX5xchvcN/lMzbMSBH7LxNnp+yjlTdV9b
wLW0zDQc2nc/s8FBVZ3u3RWJ+DIR4riVFUraPe05UTeECYr2YZyGTz8ZUZ5qLWvy
oIUeWdx9gAHFc2ICv5OVm9slTGQFaR7XK3n8qCn0DLwnvnr1NlPMF2nAwhrfi/YX
i42Hlez8yFpWsWdsWCZG4WN2hUP9q+65DztBEU9LJg2FHTOqdtlP+NLM5Vpskmp5
lRJE9eauY56dPootvrvdWbZG3b46hhbFzfjkXv5eE0XN3/cQWAhlwDT8HSareOWp
y4pRH14Ta9zsSSSoOC0RMsno1QiIKyDp8Z3aykwogKOTXyCLVlXWnEtJ+PAGSUEK
e4h2vc+leuKYkqcUB485e9wyyapEoqH1u4yC6beJJoP0HyRenho6v3yB2PJ7U/rk
qOpOGX/Lkt6moWiObsfiRuZdoTzQoUP+v9Dt+HWtREdKq05lgw5x/RRubzqPbL0z
/NRx+WT4e/pUsY/fDNMUIV6d/qJjvMwhL7/70p/Tz2dBt7xCA7OfTwBuq0HZwzFE
UDgaPS+BUZwQh2XFX5QbVkbxIy2D0u9ElFS/G8Ul8jl+cWNsc+e8iZ/CJZQOUIg/
GhVO85YQaY7QGrJNR3MSc4nUHQQuU331v4hGIVAdXl1Yt3TGQXQROgE2ERJzZwEE
i8yYcSGJRkwYvyBaLmuMDKt2F0FNSp0+2XCvdu7n96R6lnI4rNGoCwCvOw4I1dwx
wbyYJGckM9Lv3pCn+vFSa+DjlfTvCOS8YzjBNq9EZPnR3s53uCpSfXQIG/04Ts2h
zi+t/6gpL60p+JXkNgdxb0mb3PtYqE8PX+xhAD6ptsKg3DcbMulJ8ng9m7c7Zd8r
HCwpMwEwS8XWbaOa+dxeiQo93zaXCt2yATREgoN+HdiRok1I1j2836Md/FRFuqI2
Xw7W+03zNMoY2XVY+dJgcEDixcd/zLoY5j1JnPZwKJVAhwI3gSq2LoSJs0bNoNNx
EVpqTVk2o4DccJ6wNN+99JGdx87PMJefDSmmIuWT//s9zTGfTGjHXHL3XELLwwmk
cJgASs7WHAq3pzYQ8nu1HrQWV7qfO7wHrZxBn3d+N1qnVE1K8tAwXjmUnWuvlnT3
Vb5tCv/QkaVCVOszWZjxsA42BA33MUDS+dssrFBVhgC4kWnSIrslHuIgL1EpbOQl
O8fzPOn/BGr51Qj08n8sRG5br7zl5/3KG+WE8Zi+tV9Tv35JgRrtCvUAdYwg+Y9w
h0Zb/6Kzl2YgfF8ZF1sj+6W7Q/HaPe3VQvJLpMivpY65cikrgtBMIGm2gab1y/HT
/tOOneXmHVAAA9s/Kv85Pcn+zDrI6zgP0j4URH8aL3msf7aBozfsFbsKkL09d0JD
MCcMwpcsRKpIXljcTnjRd9F+eF6PjTadz4CRxil0V/QjKTA2gxuvP5wUk9g8X8kG
aQLWAxhgn9Xab6VRzvmkm+7TyW0QvJaa/Z0BnBook5i9n8jzCTuz5wA8ENGSoU38
9WQaxriKK7ABpmPqBDcmxJahO/tVV3EoM1OSl4v8asNJd5G4z3Jd8AKJCO3/DZWq
7uHe+u7Cz+rrPTEAWl3eBFyhW1LgDMEx/TXaje/L9O8eWTxSwsh1z0aBET0m/6YQ
2CCSkGSw0mrIBpwB8hMe/MNvB0Q1lL0GMzYVGMY+Phv+3+SKxgDNsmbqk/CLpmEe
NdLl4DjXi9AL9+w8Z6tsrqCGyKeeHEfA0FejX2DGtWANCqQfm39K77CMK6+/ApYN
v1MdAqKn1xBxnxZ0Lc8/3jpdBLB0D8jB/uo+xHV2mXJBZwXQt4iLj8oZz66iPawM
6Fkh47mqT8JTDY/wu512jX8sX3xY6ErfnSTCoyltHnC9YlhucHGb/GrNOjYLqsiz
GkZ9OkZq1xzvpTcETYIpr1GWLMDfkwtvWLKEZQsMQv/NjYcNFRwjXnqil8FufCfS
1cLzzLYXuIny7OiDRPTWpbCjwhNdOBVEcXnhoKUdRlmbPEPtloLvRpc38mAyCSet
cf58WawETmnqk70HkIpo0wvnKqWEH7BfXf2u727hbgbNnL87IrQNItYGKL8LbH4W
3pCNE+vBrpKw/igzmf7fRh5yw2a5epnA0jRoWqiMuGUHppenoAUTcKFZGsAyUwbv
L877uPJlLRXHLXuMpHroZqqX+qTOjfsstuX6VA1mtUTze0bccJX6bjgVsIoH6ljO
VozhjSqDyy99PO4X8OlyycpOXG1u7xvPTaQpCrV4zO3OvRkV/+rcA5KaGBA2Iqrb
VBRDGq3C9V25wUbXNfcE591ZeXy4G+tzCL8eANja61trInMGwJX7TLZiSHQ59+uh
p0W5risW9Z19WLaQN1y7qTquxQoy/mYLHyPztHG6pC6HhXgYpfTIS4KYeghe2ZBR
aIwV5/Si1Sv6u52WcCdwcuy/K4athE89pDMakF8IjmB+lOksvzi7/xoKUMihvPqQ
qPRbSaBmuQ2q8qAjAfGlrAM90zwBvr5+WUqhlgCVDP7RGmEQQRFFoWZ6BKfEwYnt
Cbci3oS0u6ynHsF0kr3F09zRczkNHyC+ZwJXtGqdoumBzfcj9KX62qBQGl8RiecI
ntCBhY76q4pGBVjEDed1ZZr1rBTC4gK/iZaUw9LaHrNliAbtEt/g3o/VU7V+Nb3Y
s48yj8V5dQzELxI7FTFmr5O4FD7TDxPhmMHuAsWkd5vKTafknp3yxi1SHEuLfZ6C
i1cVYNrQF9z3t0Wn1X4jzJmysxu5ODX/exBSWPecwICZ+6+do6YIrHy5rsxIf4n8
msi5COtOeklRFlrndTyskZxXuU+UpkSNEHB/pr1tyA7YPc+zpGWBrYVjvHaAbsZ6
aa66nKsGGcPpyXpUT1yXCuL/JGlAad2f2ESjEg5YB8itfRxtqeAvjU8Je4LsX/s7
+8ghmANtfksImj7IJerZkNYka+5QVci62NLQ4PkBmyuPD9TlOnVn13eLsDMp/HlT
5M1msN+5SyQInnpASPAc6a/GGGi4lpvlv2ztZL9vBVzB/cugwLl4zNBSmMZfchz4
s2bbULo7QwF+nkv52oYXDXqYwUb5+tVdQBbXxLnt0AXcCboIvmhfmtkMYbnuDO4T
dybnOXfnqa2xsorPTtGew70xaklIdx363ip0z6Csfyf6YTqjs9B6K0trVi7uvHdK
MZkpCfi7SQp93gU44GeTw9BQh/vIxGNWX37+zD4SxBe4QO+KPZRiLgF8A/PgPawo
cjTHJ4p34INNPje8Fz2ALMG0CGgw/mvurcrHTVYD1RfSrof3wRX8n1nXlI6Bio0E
BghZBAWAs5qolzCLkjCSjcfkpPCVV85FSne1wuyde3Y2hR3Eg6KIeL5yjo2qal5n
DXQVNFSs1o6iQY7lrRmOS2QJ07waakaWgqDFxamsNMAKcYrWLOkC78vCbsWYyHsw
ufV2bzsCJzMfVr4sU5ZqtqqwCSvmCPLtG6nKF2xG3umpV7S9wIp160xVwft1Wcb+
cDNfwmpn4ez2lX/6L6jEdnErBhqbL4ijigNXw3VOxXAw+LlAOnZJe7Qsip4Esnxs
mI8L82s2t6k4S8A3jl54fPxdEu//4DW5PrAo1inbn8H/MVh6W0xYlpHnZlSLgLCB
vxXVotalMKScsS4OQFDBXmWszNKalYKOtbZ3TsequDcJ2qNxfA/UXcve7gwOonjQ
ckygTnIHvgiZTT9Ds2l1Nrx7jfpOMaKwFwTbqo29q6x+rYJb9iObuja8Y+1owVId
r53dkyitJPXJXzzUEbU2zJWGFGN+qhmD5O6gOY4pc01H6m0hwuEKb+GB4cysbzAB
Jm4Utp0NFXzvdC2Muon4y9CMk5rigY7D6T+2HfcyKlfq3bOdc+/mn3jDGs5lf3cA
JGGZ6bP9HlorwQJ4R6Dx+gA91ZmbLNgoIsGQBlpKqIJgJHC/m0wJW+DGrPpKlCDi
Jrsza1gf2zYD3d0ReI4qiwTfxk7oYHyZ3UAMXb+qsWzVD4y+IwHx597PyubeW0yJ
xuWEf/ZIiFHpzLWZZxK+t6yoND0QTVYntV50MF+qE/sHh+QoiMC8PfWSsta49ZKy
bKa3AJ/lsu2X7t80Tq3yBkCDy0ClCclADU648uBqCohsPunc2siHR7wPPPXrvzZR
8PaMQ/9TfoyRuhARR0BkdpwuWBhxsSuvU2dHqtyLkLRNx9PzJshHaZLdTbU8wk3S
0aRjbHFMQpV4GxDjR0gVogVPQsaTc9/LQ457FQHm2UcIs7d1hhS7ATVa3xJVi9vi
taxb9/WV/WXHA9Io3N2NpiONT2w824wCOpBamfdRy2OEWQvLaclPvwSaOWoJI4Yo
vOcd65p0mmYHNY4VLURp/khHbU00ipJsUoXiMg+LsROeqyHIrhq1E3qm0CHrHuVr
bV/FHGzvEB9SKcF746PYgm8j1wx9qEGfXyXUe5EVSwVyTxN08Lor5m9M2GxLuhBC
QXxZLSk8cpN6XwyFQLMTSqwifPq98ru40bAO1S6SlhW6GxWUUT2DP51QrBwT/NHt
N7eh5M6HqkuM4wKDDG7OfNDAsBP60g9K8bv2Vit7mB24dpm7YaF5I6/tGlx2WtuH
PVmgan6WNg/uOW+ODBvl/4zv1R0+QALHYQpV6W4f4HUKfjSXMKd2huVvC2XIHcdO
F4oBpMDxapFV2Uom5Pyme7M0RC/opMkk+hZP9FEtCEpFwGsbxbGNED4KPlG0+lTk
wJ5FsNRkw3kzgH4fZF54lZIuoN7ze9YIYOqjmQDWb5dTUgW/ahCnlYlOrmA2DHix
MuL/WnW1n+d73kUszbvlrhyWze+WB5o03rKfQQ8hP12zqeOkJm0IHFAdyT59LMr+
vOLAq233VaAvUcKt+NpByPuK+Tqp5EuuXBRMHpZNBiMrLBbV8A+bHRd1QcSSQW3g
7kWWQkXohETLDGXEM+PLBojVn7QCPPqvJeYOO0O0/Y7lP22Fx2+K6DgKObW31z25
JPwLGEE5wV7HkZBrRXDYQwzTE202pErO3AujFBm0cZwyEMv7TmX5uYLEKHoaf59H
iXrqnVFZYLlCWqgkBKFk2j+//WPxEnZzotyLmLZql63wjfJumd5pH7oegwxiAagB
IoancrOhRaQxpp9WlcqG2cAuo8yJHpLBUGCps9NlDpwcsDJLhhcL/FIjKlz2m/rl
pbrXfh2bC54/YEnE1DGixhfwlML8KIN3iw6vH0yy/Oa0XmHYWhOnNcdbweM3Aj9P
kbIExZgAHufo3Sdk/JaHKD/1Th7mnj91Y9gF1NavVUovNbteTKzyKcw6R1pgzzpj
lEwq/mon67Ef+KDsHKKq2ItKjweHnmiP6ZH0YhPrV6VeIOKsFe/EE48nefy02yLa
iHqzKaZ/2MB7Nsz3pR0OgCjfZzy7wnRoXi8lTPAVL8+JO36nhTvolEf4IjSDTL/G
mWZsXF3G1Kgm7kPNBtIt+wRwQ1rPV+Ilj0DwdgtjpM6TTAT/G1Hkf7FPfIxqbF4A
1l3hZGpasEXDau+B7G7XFxdjJ0eISpNeeYsLphMKkcbnePULyfR7Tc1fb0Ed5tig
uHcIaxCUhfa4Y7L+HkMtbBtgMBVmWbzXlEfE+oRCXeysDb7ht6m49/BsDI3M1rmi
j9hhi+QU7U4q8szPyeEphqIffw7KPJGQ+EhP2mN+a8NamrAK0M2SWQ0MlHiheDvf
UrWvY49X6gQpFqPCADkYKi/na4uRGiqZ8YrcOYTxF7tI6VLcN4YqMqUlE5b2Pcbi
7U6GzRdbMdUKSuIHXAVMzx60rp143vwKrHCgDTS10BKxCOuTS4X2B0JOVAEoPUdm
37toCFRIq3z7kc9DrwoaYZ6TS5n36MTHHrWUPWN28zpkhXJvwLvVmXFsGpNI61/q
VswiVMyJ0PYMz9snOM/hVKoV15HAVyCTz9DRtlkWDT36mrYyk+5MFjpOKzUFhcbF
Qrt1Nj3pSVsmO1ESltThZQYcm7uYkwLrKXSjk0qHaGoBC/eWhq3kF1dsFVYI0lkS
MYdIQsvs7cM+3LHzRfzDmZOcAbsuNZrVWFniKqYUz4rdsG5oozT7UCvYPJ+zjpcn
K4UIFj5Un9igOLjs0BXBjZ/67XN6RJKdPgjBpYV2Wu9KWEuxHGC17aCIFvb4X6GE
cHqxYHEtrqp+kWV5Iespfw+VmfMu3CZv8hoTMBJ4S9kJBkH1HyxBshDrPviagxHo
4f2W4iTYMrYtzdHDdmfMwFC6H8FmdhXlbuFOukDiz35m2SXsUo2VoHHU5DcFn1TE
bIrlfIfSHf+u4MkPBgFXVLPU03p/OJA885twYq6bYsEW+KOzDrEbwQhUkWkuHBWj
03YWQlw35qZB2In3goOBUflmGlIqvR4CALPxEaQm/R9fzhurTqZGrUSQ6dURTtXx
j+fh5W8ffhh3/N5opMltZGxgTRE6rWWXtZcG56dvYhVKsG4+S2XQYz3lgoMSFT0s
aBnZqJ3K0z7F9l4TV1GYRDUuABQTiS4YYuQN5dqOvS2m8b5nBY0vdjgrTh3NjYYA
zh3rBC7oBopufzKyG6YpTcXU1+jR9/OFtjeBtG/u/jD/hdBeCz3RfLmG41YYwQW2
venCM5csy/c2o9FkBeLjvROcR02QnM4SGz63HhE0cW9L+x9R+u6+ppN8S+P/FVq4
n8X/XpcVKNSbT+iLg+Yv5DYPg5XQkUm1BlZjKifaULJlq+2+Jxf7s5ZM4PxI+/FT
HS8K3jG/ZqNV1/t3nSd63cg3FQp4mvqN9yBxOT9Ht5U4fmW1fEksi3dpr5O+auvi
GrzaQ5oDfIzXcZPbPR3aE85j8EGfTQyATXewUk2+YyEVXHcmOEFQbi776KWEJ8iU
+k9BBqha03rJoAadjQHP1q3xAEazHX+ChO92P5z2adiyI4lBm5bw1d9KCopHBg8C
STGfQ/BBVvyQLAVx+xzpaEIy8n9/ZEcd738ZOMDlc7oAGfpAPW4h0p4MhPskLB4z
UWr7Qkf3ryONp4kF8kUhJq8aIUh1ePNlrvYvaFUFNnGdsDUe8MnY629+Qc4sZRmU
Nv8EOtqzQ3+czg2umqbfecrgZTfnyk3019Sy5yhZULngq5A5oIhR163UMHO2iqyM
H83AMk4F7OdQiOAfIz9EVgel8Q8v5yPMq3xyaJlKX4s3byvRbK7PzG3u670208Tv
9hTCvaDqu88+tHLTm0BHIgqyWOYguscW3qYHcNBNKXNs+uzdCtIfmU7BpzNaiNTa
xuSZ4KSdGjpgLj34PMzPK1ZkDRxaNK3ZZH1nGkbdOP+Y1ShMTc6Ji/6FrmQHCAzE
Sgw2rEaUv9hLkaSFt6i/nfXXL4jVXOBY5I8aWF8arqJBCpfk/puVClN+llFM0Lh4
b9Lp72pAoBvfNBHpc0R2IbSEFhA34ACbwoqSbi/wXx5E3DpFHsKou8M1eEmAzTZ/
BUBZmyIzIpPyOIycl744zf58j6a58U3teuICf6heJznyEMdsgV0+1VZF6PRGfpN5
QZfWxnXofaDXDWRS55ZchjlXfIVLYT/3h2VYb3tOSkWKiy6KVnBXgdib12HJduup
LNoCufu+RIvJIqGkhXzsk6ee6CgkWtqvAV2nPdKKPuhtTNpwbXPj3WENf4XYGp81
8vh7D21K3Y5SR+XtEM3UDsoVtbRO+sr/XZnUqhO6RaXjZlRfpAFUeRbKYpM8Vd4U
ryl7fYYcP6p4xrEuZDPTdpUM44nvylXKDNjiT0nrwS/VTuAuV/YDbFzwbzeZFhf/
w2hBdWVC83ddHv9cRCDKh9XcuMLY/OWkZj+wgzLa1PCK9Ujfai42vr6KUli/SyYc
jZsATybgRpkho/ke8ETz3gUF6jzPDtTMeafVeiGeFHQ67YXo9y/sOKUULfk+p9bY
N6y1iIKMyCqEs/7P+fhzmnRxN3kJ4HxZE5s0ztR9C4PIj7Eu4Oar5IugDj7HKWNd
NZF7P0pl+iDWJaDi1PLuYm4psvspFKLGeFykUqdG5MiXiAVrFtCFyD0k6XqGIhGn
rWyxQBxW75krJG7sZ1q/CF7zEdmWY4ydtITUmk8KhrLw+sBO4tWdpI5xUanKv+WK
/w/NT4SavWDRFhGjGpSbxDubGksq78TwbP0K2hQcR7NFTBT+pdkQcTTTUX3TEPsK
8HSC4Fh1D3F+si7jTWTPaQ0blHYmHs0bLlCO4PmnL7qLhgFNpyVDi49FuiRKAW97
uz4S09cZzK7W0WrTofWtxLaOL6JG9zi2HQDZLZ9Y9wj/FKTj5ONoXKG2ye2BeJYE
KeRgCdvHxEypcr1ObojLg1KGlKmHtC0Z5Mal47NhKwgiePtUTTlCFAD07ggk9QHM
UdtQrdDCYKIXiN96V/uDgi9lFk1KhgSgJfoz8afLlgRA4ElOdqihO9DD/kLq6P06
NPypOzIQmO18FtzhATRrjiaiGLKoFZWMM8Xr2shYVUR3h8psXAOXzxehHzE+BeMr
aWL7zEYvG3v5Ps4RRVknAG/axdRiAoCzUNnS3NyQXlwOifDhlii8YYaD33S69DtD
ViYCdUmUOpXr9wolWMbQWXWvcu5d1iBQi1BaYF6PTEsfA9ybf0EqBCSENACTJg/u
3MfBijVqEiOw9IwhucPgNMDUya6mQc9sKwJMnbnFBoXOegtZ7WBfWzJpJ6eVA3kX
27Sue8JXvTrfys044LobDV7yH/hqXitXcNKQUKRB5OUq059TYbXb8KXVWWFfPS3X
1F3QXOxsLEyZ54pntLgjhrMKF+g8OvcCXm+8uASBMNDXvAabetlLOf7PPMWmb/x0
neczAfLlMyGwjzj4f8f0y4wxohhO2j1WGw3FXzA6D7D50KCi4XVpuuQknVRjnA5o
r65lWgr7/xjRbX4BwfrdbvuKzUo3rWM/MydsWw+Qmo2GgdfDAn20Uhx7uDV13HX8
AsSVbw+c3CLHqarEEKFD2bLR/4fwsgw4kqOMuS3A4nCtlNdWsGbKe0PTYFEbDUXm
rDbgN5O7aeqKc+lbWMarzBqSEeonCbnRKYyxPYNBOPob1rmvfYxXHZRxHn5ozNSi
y81Za/pjlLkqdd5m0pTwTI8k5QaFKZYChMJqCQJ0Xsn/Z4Imk+4nPeSvOIvukNWy
+pruBOIfvpPCVFxYg+qgUtW1em1lBvLwqeINx9ZsxCiMHr48tJ459VQPM3VcYYY/
EizakniMNFspfzDCkVInaRCZsMRUb0KJHBjes/Bh/PK649Aj0gXb8UnLHjEJAo5/
4bI3Thd7H98r5uBhj5F97SmuouICvKKw9epgqNIvTdTudybUkAuhDq3hP0Rvl5SX
5UGR0hhIOPXA+QnECHnPItSNXK4gZVz86cJcNsVvro8iX4Q7IAqnDs2AiTVnejDB
cGDqHes3M13rn1re1dOniWdwyRS3UvPOSa6CCG0tMVlKEY+ybBfFOFTU0WxluFjH
WyrAaIdYMbPiWNfkpXpIP6pSIfDH2pR0D/BpMx+v9mlG+mVTaAht34g0qVfH46Px
JcDt6RGBL4EiRIJ27VDoIAVjnWCpKK+v6ACTlURghEcxBDtWnFLNkWhgC0qTkoRK
xKlEPNtjbtCqJTDKt8XKGIP2CWH2x5KDivp1srerOqWtl49a1ueWhS6ypwOT2qcN
llGJaCB9dkTPp9UDso6dqS7JfwAWa+bg8k9pvocgvCzrQWjfq6Imb5qzyL8Imrdx
A1dnFC68BrAc5+Tmorz+Oo1N7JB4TfjqsCxw/JikSfxyXE2jGX0L0UAVXpCzptqT
AZnmT8610lJDFfJlLbJJuYspxoj3iaNOCHLrSDHLDJQDICrrB2TEo8gwUFuadrAf
UIqayikdbEj2hOipiVINm4Jiyy/hAlmzlP62unEs18xQzyssAGAEcyzFxDr121NB
9howbbV+QmfbPRdSfoyTw2TxjLAy8s/xjJX11MX1HOocBWU53GfmuNg9qUGYDIWj
wD8zz0XO/FAJI+dO8vSzHOw3T+z01c+dD+t3cnQMd0Gx7hSf44y814UdXLbhhOY/
sO0DSuOnuSV3+6yXwKwi/aqae+g9SwHGexBRcUWmA07m6P4KTj0OyZ1muSfAGoOT
JdyX+j9UJzUV+ytuoSHLH1Y9hNzKj18vz65aJKvCkgaUQVRL4hhshOxgor6+EmEw
XdHc0KHZhqM4YH5aYqU9pFieMuRL5O1G42tPr1UFYdQhGPOnwPM14OiZjCPcxsN1
9pnGMyD0/tc3YsX8jdZrVMQi/BbFrGmp60EUOCamF5DEjhTca6IKdI191wce+QT6
6BuPGYCgonXDUvw6D81YUPgtsbPdBQrUBG+v9lgIOq5cXJxDqmgqsdjtzGC6IduK
HjsVAcTOpo0prpuYNT2BlYmSHSWhFWBi6gvcIBnn3d5L3TjYrihcoowjuZuazbD9
MawCkdqumVxDPhlNFkgJ02vHygK9da8jVLGxJtjL9wBUKrnfNAcnViynj1u/TNFY
4lQ4t4rX7KjT10FWJrptoNoJIOrMUzlw19Af1LN+0/5dDqqAF0PgKHe9MCLUAhP8
Nr35Shpw8gkQepWIqJkv8R7QrQ1AJSXgWPXX+p8Hu2St3+BHNXMMmyfTUd3hIkL6
ZYoBpN9tbX40YwhErPqeXkVDWtv5FEnX1Lrb03yIHOw2xBOrukYtoane3x+ubOfw
PETL96SNRX5R1VYK0UKYovWwM5ekKb1e4Au3RcsHNvlrog8No4U2qw73SFdaXoL1
bvXC4I46YMMyZG4MTjVllxEUOKvzEbqARiDlh01rEsuu5FZVbtNqSCWQ7YNlV3OC
yEljny39TDG461vwotcyDU1zDG8bBE9chP7EJHdNIhBT/2F3DUn43FBi9y+YvYj+
U4APbu9BVa1aEhDMShZDnes518A6r1gOIuGjeJ+LF3v06c0LJdxczFhkNPz/0klb
C6a9m5GzywmeOhr8Pup9pv4F0gHxcnaHQEFRnNBxhji3dNIaE4fXNvVDQMZIUZwe
15loAQzRC9HoGEGSYON2CHPcaeDbeoLpiSVmxHKJOr2XwYsmzkgsaz7d6g+B/ThT
3eV6xIZYJtzsmsysJ6MPNfFwdDgb9xqEgXW70S7jtQh1RQMsckDm5kW5GAbDf4Kh
nubUUEmW+BCWmuwxaznzEK1odekrkUIcAHLUqOV6omofVGeCV+XRW1VdYbZto3of
hABk1hvaFwBVkyjA857A78YJsCVCDn8n8zuaOvxnoyYfdTZUnbzu8hOozkoaHzoM
l+UpKdmjJnLNsExMGdW8ltSKmJwUWQcrzoN+p6i/sEoO3YFr2LtqaMuWmw5N2P4u
9pyXIY3Xvk0uplSFMxhanzsHhpwdSQTNr31PX3MtukJ/73WlfZf36hiJEGPP36jH
VzQhK4hBc5EshwEhfL4wpHkzirGnv8uwhbsxpNlLjQijpfUzBWsoNliezKA34G+r
TtBkeOMYBRTLJAedSJyYEKfyefrzopEY7UK37E7UO2uUKowWef5SrKJUpAj6GKWM
h1yEzv4tDaFpbS1FV1FALxtivFSrx7jIZ/dz9cePULoguQyuTQv4PYI7kNmwNJeg
Tlb+MY0E+4WJy9JLwSfLiYDk0Yu7W7yqrcR+/Sw73eHMep1w5GzeVD444Mfw9/6v
Rt9PuAeubfUfzCvbh+8aa6FXaoXKf3vakeY3Dyn6xVQLzoDLirr3Nbbz3dIYQpLn
7DDmZg+cEWMP3qFQVYRTktfGvc1bZdKrya4R/EKSxojKxIeKY03wSqd+FyTOnJjq
l4HwMEyW0tImoqqA3r/+7jNNeRn6WI3EUVJ1oiG5JLDzgZlzW0K9dozD339N82dF
j+6TPlpSzRpuuY7KbXjicGEfhrXRZrHUmGgsT9CM7FHL5y7i7HIOpA0BZKcgUbfa
Hy0DNO5Le2x+Fiwjx4dFdqHnkgzhQt/oY8OpsvtQnv6X/av/wUYji+Eh+QsB1yOm
DeIpkJoPOiwowyYA49ylqD4NfmBtxws2KbBweTtf7W2TpyYzFZ/7nk07iOC02bsO
25Ea3EcmxhfSGUvsBsgPis24gLCdvsUT3aRbvY7donv6LYjpvk9pQ6LB70+wpbJv
lYa1OWSY+mh22PTSfCGLtE3sVHdwwh3YdznxXrR4VLJE1E/RezAhheubeUZRtpPh
wI/gISdaUmzvnjnuMfXOWAAY8EhpRdM2qIkN2FGXURj8/+VD3p1K8jjAAV32r+k2
Wt+cN+jyuH6KpYUqk3zCv57guHFgrtK9zbpxOAMm5afczN6TzWoNJluxWZGzeCS5
pAFCtynRQpdmsrhAHtwzUqyLIMVElayb6+A7FJvJRCtzqdn6toV+OyJ0CrPLf05t
kwFi2EVOt+oMl2UMpiA6zpaJghLU7DFtorP6Ev8lNFLP3uMiGv9E2q8qJf/3EwDD
ZLgu/xdBUZdUewTcRVHuWXKNumwZ+8+2FQle4Co5+7Bg8fSb2OZdosLUGytbuSbf
umiH2c0n9wEgtaTscCvb3ekKO5H/pfQuBM1UUbThG8FMzECJZuDTD9BZ06KhKv/x
bjCv+zXrMvLlVIZdkABuMOg/ud6rXtFgK22mBt73pmw8Xp+Tpegq2hL4SzK1gx2e
yGUK1PJEKhkKf0Q7K1u2WqL3ciYEqNiTgEk2Kx2kaOQNZPqsoTAe4kQoGVw40H9j
+5SjvicYWh3kyQgxtLDJWaf8Tu0keR0sKyXqjB3oa1UJ87bmy5rqAFNcBRp44Re+
xDhj+4UU9F6X2ibINovSNVm5JRkulcOIEwDWtLISSaYqrw12xuECzigwbglRcyE2
nc1SCeskiynElO2wMzhAAPPbhbIC4MuOHb38hNc25RWX2pgPDmWNJqCOsfq7Mb9+
j1wvoGfV45pCyHgYJC/Svz7oMs30WlSBswlb3kNaxbK2gqrbODAXvSN+VGYo5l9C
Pwp6kEOD+eVmq+Ns8BUycXY56a0CCrftwJefRkwIarDA5+Q6WRJVXNEunuWb1rIY
OxszVG75xTjXi4MIRCa/Uk/OzeB8V8Jmwwwm968pU2Rj1iQospsJXryFHz4cKjKW
bWbqNRHCOvaOhJNEnBwmzjnN+fqwGa2Z/ny1M0ilAeWdM4/sDdmqHFHH+9RXkfOO
Mw3ZsrqR2/fGYphQBPYMElfFExFvMDdgCvQ1GWrqepYbJKwqEc1/vqxkrnW/RWqB
UXKmN+uYmuA+TA0al+Nvgo6JWbNPCkFATe/3CRvfINQpLVXE1IulVI755r+CwVz/
Gxaa2w1azWcQn2ixPD1hogMuNmVA+8ZgZdrKAXv26APnt5EtM32O5iC0INbbpZpr
AoOeO8mNfp5BSJHj4p9IAiDAHnWQ0hIEAbrhbCR/6s15x6mLLm1vFKlvPewb2rr+
tufu1prU9Q2+g6vivaeepjFKqm+9lZckTrySRl8lrYF5GjjuhWSyKl5jhxIg2wdC
PUBqf81nKeD0fDP8I/i3Ij0A1wuSD3oOHf8QXTMz+C8r8uwlQGArZOKqkIuA2ER8
Y615ZYDDpMBdYSXMulSK/QH6I5oQOHgQLnSO5QFBUJig37cNbnRwCRqy9Ldd3yy+
Mzv8Z3rGm6HRqBvuhFPyj2f3mr7IVZtmnHzejDPuk8Jeo4o5EryOTzLX/Nj81129
h5IsB+vc3AloOF3djqPU3jshztiIRiMGWC4vzixOOtEO8kQrF3tSB6ELNYUkyJmO
JOznv63tTDW7BHJdeEZ1Wp9Kpl1xFe12L0jUnhS++dPBYn9EYVdz3bYGtWS4kC9Y
Po8HT7R0H1hn//OW+Tniff+ubXjDhNmEIarNcbPWxV0ZxtKSBSfkFdkgmS9VgH6T
tv6IZyG80Wmm5SQRydbCVtu4mPFNWgENwj+sveez5mTqPpNnQj4g597Vdjju/c0C
ERc7q70R71T3F79rEAZHQDiGINLgUelMiBiYjAxGv3UK5flfs5MAPb1stHtc5qTi
Kqg5/iMPH241tMwo2zcR85FWVk7rZMcqDo7hZ+jfpIWaWLaDjroTvIBZa7K/C70S
X7tXg4J8yzPd+d49d7YLxCNL+cTnd3ym8jESvPy1ezLkxwH3e9IipPnDWtecrkiF
PywkikVFv3gnVyaVHOJ75FiKiUJ2ygKjPz1oo/NImcAZj0I7jhooMUuDdaDOmU+P
m0VxlHctXKdfW0hpRiTMWCU/9PHzs/Vy4bEKfE5HnQHqx67kPA1Qn9shYL+Gnxy8
tSQdrnTGgvRuQwZ/xsNQQjXOmvMfkczJkoGNJrGROXo2tqzJSURayz1C0udOPgta
qNbjnD53i6xAAGRv2I9Prp7p2y2ro3sdRInACIYoDTCqrPZNOrRMZL6RttAyxLLy
TsVR5axKpJt1ljw1JfQoWis8G0eqNgdKf93hySfsrh+gA3aCV3UwC1llkZxVmFpZ
g+W2nB6zo1ksOSSlKieUvHm5xOI8sLG6ZBGAeu1EZwXod93LnMh9X6tBUZxu2zQ6
2ToWeHvIkKIm3w2tOwQrzb/GAw7OsCWWr4/J1qjTsPUvf1zeQX0e2gyDG2WtSBMN
FFNOW7lDL6Kkgtdys5NBW0PZjzsJ/L4qqWHc3UvYPWM86Zxfh6mR3Tg2WJ5bY5D/
mQclNaaTctAKeR2ir+hVwnJNh7gGUB8FHIjZ4lZz1EH1SFgdiVLdF8XeZLPAKn28
EarUkFMPmOyyPTV88lGZy+yaqHOKcEEA72lQtjYkpnQnVX2IZTQKhf6a8io555Bm
TT0o31FrEhRVnZ5+/m/QqBvzLLG3O0rvVFHmK4XFQEMp/88JoX/kovfFqZL/rdK1
61yXzN8hUQ7j2KBCHkTb2vQt5A/WkFkJa0V5dk95sJjR41mPc2pf1HkzCWUAW9dK
EY1Y9zMyOB40jMlwEmcO6bRF7qawRWWFwOU8ukcbvjj5u42uU5t8oxoGCyvMBnzn
VKnVE5VuTag63L00yw20QH3Sm9+5fGTWwMjIDWo3utTD9BGl9Z/BaL3/8eq5JzwR
yKaVO0mlUVm8TSUAZtyR2GHtq6Zv/mFvfxURYN7h46Urf+PE3ialetnfqm+R7WOt
Cnm2PgETTOweBP45ijt+JkJYCGxTsz7uCkaBeyCZZnHzoSh2Vzr6gMJleNWE9j0U
kiuHJVbFFg4U6c9UaakSw0JiDSLcUQkIDhnwWo3BbnXWtOpcy5+aasZ5WNi/hKj3
Don7qx7LiU864HAUJX9WLMwb2xiBAVHyRUs8mLHU3jTahVWkLDwLj8crb9Ay+dQo
aBmUoc9PsDpfMueg0sb+YBzqbnbgdOXcuNisJYpzE5FdXMufGnogbRtCEuef933W
X0tVr6uamEZQUlSuBsS5EeM1pScEjYl+qwcKl4dv537uboq0kG7nCAajXC/v0ONQ
VqwgntwZTVuBPD8AD0RzvVpMjYAc7f6grxR57vbP1zdiOGSx4+FlJZDradY6QQNB
c6QU78mbQ8SAzJQFIHKIMtMBPKAeImy7n+7GCuKslxiXp/kyKZEkcxLAs7UfUoSx
HMBqRBKaxOuler1NGSQLbSnVxH2JcBv56Vp4VSIFpC3c2mCF9mbZ8wEOYtVYEUai
shr7Z0ISVINhcFVu5bvge4d7Yy4jsu907NwPfVGxkmQcwC0igEj0cKQwFLY/dcI/
OpY41O8VvIantRu+V0hCbUsGcxqkxgR6nTA0WgbRmFSENeafRClTvcolNyx+UzRJ
ekao4YE75n4qVH/c90Wkgy5bbxNROA1/zfuy6MJgxAIHIE1MLkPa0JnrFRqfXCEy
li5XmkoE0K3WzEd2sdNI6Eswo+xxGTcE/aP3ENDfRUNBdjE/KFue1OKnCUVLzIUa
+XZXV03XVq4zWzbh1pe4q7o4Gh02H/FyJT7KoRR6CaLgABVtvHrMqDRnv7GWz8mN
OLzsKyNoh7K/CCneKOPQOVXM8Ec5DKRinSWkTbfcJKZMZpclHQV+GTOpKVwM9+hH
OGlbgy5zMjB9AfZOTRh+zggc+KUJwM9sx22sCpVzDlFvKAaQU71cUWZ3Qf2bG3+g
7tXR7rGJPUExVuBalT/A6CqiAwGydsWNWGTXpnG/6jvQh71/0xJEhQ4Jc4QXVS2h
rYqIu9LBvqwE3zpGYkneoJUn6pJyw7tZiMuis+M4r5eG0f/X6NEvHmcmmAvrwRpT
smK0fR48WXLjtocOX8TkCA5lShFQFhzzVKZmT3Xw/NORVS+pT+6pF1ATYldu6jZ3
fxMoml9MVvI4kQSSloVjXDNzIae84ycpGaFoXzqwfm3PXOKCJ90Tct8niVO7DjiB
XxZR0GDPjIP1w3pBL+xn16EiOZ43iNYFRdorscDFdn4Bv812fDLA6f6erfVjGK6w
22BSuCyyz5cR/KnB1jo4gs8TkjEHGvfD3xNaVLVW9VEzfOieHdfDmuqC2228quLt
SddtxZXSMlGitxlK4J11GqZSC6mvGyefRzRdWl4mPAPxf19RU1opUQr631x09QQl
oWZfIDycb4igIcfmRCSbaUdvgFQ2So3lUXR/RbKO6ce4Iav//kuUIlpt92PF5FQQ
oVxalRgJ2XaKOuwyFOechykFwDk2ESOpSR//lRI70QiQcsxzzv7RZ2k8xI54V31L
yFGbtjd0O+fG+gliROfw7oB3/0xroRQSUzKMNSDx7HNjUyeZW+dzaKnF5m/jwTul
imMNqMUdh2ssInsxiwPRD8mknMkcJ7ezkaL7VE5LOcTqNd3oMFQ8ZLxz4JWv24Oy
Wike3N5gnmcq7tnqToGJ0ygYVmFQn4sCoXSAmUMAAIEuD2V+JW40bWqb75RQYq8t
NbeF57R7Az8O188EVn7BrileP7V/WEQZElgd8VX2iAPyKzjktoNkpyPY++aghN3+
bMkv8DJfbQbo7ET6nwjuNNSZt5a4RGOLQGrVipJg3giRduVjhjkcOmOkrwrSYE9F
vKBM/C0DoKdS4pEKOVLGaY5oWQq/BLVbgoxOoTDOH/ENSdiib7YINmvvaDrblQs0
4S+p3sDDDsdIdKYfvwZiWJG8NQQ6FAWTb0dV1MkG8bc2kIF8Mfnh7RzDCuj82+zL
w+Hl4A9ap0lpP7yXvH5JekilfQOzqZMUyx7pHCHW1eYYb74znz3EEQK+1RfYm2Vw
a2pZ/L+2py4mUWnjPvVwwJ3uZx75B7JjoCidON2Xs/e4p46MT6X1lFQlPqH+YSbu
OJec0pSpgMGaJgdA4MpUDUZw3Vq7wcHmFSaOX1d3d5WDQ1chia8P7ckJCED37pMF
ht7Nq+f9i166GxI1WRLdYbH+iE32sOvmot6R8LWrVxNVBVd9vwth9N0zNp92c8Et
1IrHi5RCQIJ2wlwzJ4jPnD6ZIU3VeGiQAD7rW6M6FeZSnOYQzacPRnJCg2o7sJJY
Z2MzMYa7KV8Ty9ishZl3dS5lH/+1mP7F55M9OXiNKw/tfNU6qsAlf1gg2ttEIpnf
Vn2n1IvjEPygLuSA0C/LDgFUuiVUXe18S01S7s9PTgxinobx80sTDgWKUnHKSx5F
/LNkJ99tuUkg7xh3/bMVe0XdLWfAthoao/rqvX8REGerHnkFC1IXsWFjs9fB89kc
GQCGdfaSItsYKalBIhMD/htXRYcYQtEXC2LJdgLm7yhSb3EbbQKmsl1ziNmFlAVV
VkJU+9Nmjl2ob9j5QuIhgjb0aPWQ71Kr5AIoET8x8qycBLb7kX5oy4ofNAd8G7D/
VIJ3fqczeWukKppBbpSK/BxeJucOiky5rMflXwjno/DuIGI4zr1zVLewyuzi9nF4
ZHQD2u9WgY4QxXfTPWNIgbVRHA/HplSp1gzqoCYrWlbzMX0xLZP2DflPdz7IvlIZ
i649eAtF+MIL/SuRwaDCvb77E28qMcfaInlP0AyhoV0KEOHQToXBD0Xq0u9V5ocr
Dg1VTXjSKRyiDBw4gQ1h9wPYKr5B3H5yJOFbKnDs4FGho8MwBI+e3k8Qb5xLNYXK
qchs7W/x74LOuXPOJq1CByPIpZLDGB5VcZiahQinmNPFSD0nDg6xSYgTV8DGf8Q6
MIn9Gjykq9OpgqgIY5ROjXtYG5EXNGe7JI+CQ8q42CzbFaifoFNu1JylZ3dI9QjP
AEc17O5KWbsGZ9xyp4KKXHe+rT9E3Kq3WIOM+V1JQOgiQLgLxUwXieEOMcBPqs5N
KCuh8y7jA54QzuTZcPquG5fAvCty3EqEi70PVMJHBxd1BcIsiLhlL3iryXaoTXRm
Q+xVSqdbcaMVTzyokhAHcXaPB83To2GbHsmXB/0R7+E8MCM4LZz10+gSCXvnzUoN
ppGJXnWG7Ci2aFRsRicDPn01KAlwxr1jGEbpvxqFvI4xZ+3tYZGlMjEhcR/5WK8y
DEfwBYfeUT/eXiFefD0PxDgXVlW/X6RzfsXq8s2D9J3uB1eWZp0njj0fH2v+7gNQ
G5Bq/Q2kMV8N3imT8Jc4LIe4MVK06MsEdrqArqLqsfr+HwB9tiStvU1Nbam8f0BL
IOvcSnEZpMNdUgzehst2HAohZlgJujM/SCIYO3imHgZQnSvIYy6r2FsnbOKRjBrZ
ewaIs0oE1D9pMfhiHxVc/Al4PMrQ4idC5z3gsywRtY/u0wISXZebqs3iSW1JYC15
xJKhk+B1RcbD8bV3Sn+Cb66iRlSUmnRRlsY5Nx0iLThEVDEI7UK42uJgw28V2Y2T
MbsaDJiVs8gVQZHuHLNhiq6GVWwD34xPCqZ4mDnyTi6RMVEL2QsM2Q0KizBtN4wG
iP9etkP3E44IvprfaPyACM/G3AJyaLLskE0zX36hzZ+28Qm44vEYhxE8X9p5+GjM
uFiqmMQ7kLpbdPc03b2FrYBwTp8USoapYg+aB0N7JCQ5uoKNQ1raNgWmAPKnbXHZ
7GPrDesWpoy33fmMevXmtZJSnR4sEzfQmnFAvxxvRf7s6hzEoohK/5ETvDS4T+VM
d7NqItthZLAGuwup6GY/j2UAakB1+7OyQ3atK/gfUNLIsEVG/czi/sUEzI5xmiIQ
Jy0Z9NLn+1GUGRH2utEkpKgiztJMUv3JR1ZSZg5Sqq6EWmsy21DG0XbIoNffcc67
HGMfmke+g6yrjxy62Rz5gFs0E5HgW1Vmfg0qdPavSwdlRxhz64ogn2hEAEdNbHMK
qPC7QztSugDLeAi+pkXE5B6aivWWPK1UXyhas3fFssR/BPMjGBUNFYG4SBlprSP6
f6jZ0HT6t83P/8ldo70vhazUsoyjT9nwAegWJ89hHxt2+5HkHe8UGrzJHXAe8VOA
3LS9LPaKm/ij1gIDbXLurT2+TKxa9L73kqBK/JvIUtmvKE3heflda71ak+WGhHYh
jtcYQoVpnUev6gB8gw+CpajJkkAvZBX/0GrfxW9VYT2QlaXy24hN4stP7dcvgiGx
g2ir9tw6KmgoeXhjz/VW0Wow2b1NWHOkSDOA3fuAP2aDz7u6f3OQOEd/s+yp+oH/
LvdJqukb8elmyCCVHnaZ7mpGc6OU0TFdqX7IlwnStdlD3tQRxqAD+IElrKL0CFMe
2YddCHQH0c4pyyU9geReEEgODI+KQd3j89+RzHPNowispaWcMtVIWcHLYdHhUGxo
ne8zCke9iqXEf5eQdD2vTsaBX9BZhxa7PEps2zvS+aQTdbdiOJn6n55QhL+VeLAd
67oB2wqmoaSnKZt95l3D9I24ulNnfUFYPmAc9aB7WgUd7PQln6ABTbuFtEqFuwdz
1aaXSl4vngoZKpA0MQYvES0zNsx4DheZXE7oXg/YRmDj/Gp0LouFmcVb1+WSOPbh
3ZlrXAYtZFzsYisGGRNn1UlH49fPvxJYR/CD5Dy1taVWZym9kHJnMU/l3NTvEjtb
65hRNx1/G4iSqQHKg83CSK/FvcYjYYoB/gczobtuR7vzjKIpV0bHdPpsZUFQaWiH
NYH4UVYk416wBC/E/g0xshcgcAabP51KBLq4jXZn0cu11XIvlDz9K2AbtPj7z6C4
GdYIKpFbBCHmst3NQu7mQJrvjDpcXeq1s2VkbmdpMfKDpM0p2vKqJ4imLHX0nBxY
hlDrDSybHPhDb60FzkHsy5ZVgbf0O2kS5G8rYcvFh5wK3BC0wzT7LBo/jXTmiLCK
UFeJeL/VfbAhxR3wHfRdpaVOfy75+G7OzTTcvvSy6cZCms3dhPbYRqwkkkEfQ2X1
8tvjU5Neo3J58fhcVa/MZOx7gshmNOo3MC5+mIF4QOwE0hr1/rO9iA9TYuV3zLRN
NuCGefAFBvOQRxk1N9ejTKeVMx6TKH2sApfehMHLHsouhckd/CBoCMN4OgUb5S5d
qtiR/nr4i0sZFkOEGTTFNjRWlTzzyBB+P9r43akEjFArE+rz1CTR8GuY8dqoz4C3
Jd1JGSy/DdMCb0rekY/TPcCzCNhZP0zEWp8bet1j3lRk162GWPejw/Mj18kITwl5
QH8VW+5HcnbTJKypWPhfUqccNh6oYDrasJ0SOfBaJMF3m2ijQIgVejRO9/x5CAyY
WborXnhboY600ZDZ3AOGZOPm8MbtFuxFcIZlUW3Lf/P6qbFKNfh3OicPeY7WwyDH
iVTcHZQYGofndXB5bZzugFQi4VtLr4a8B6Ua30MIzBf5oCcQAoWYvy8Hr6fwJTha
nhREZd/Y388iQoW/iLFnMVPS2xpPom6CPW52MOfbkHxNyj/N/aEjax3Ew3tSjZm6
ajJ5q82H0k2UmZoFr58FJnFrOPa9gCx9F+6POmysYtvR3y9LfWg3uCb+gUoVUWm5
qZKosOl7pwEpl4BEHlzcpyAbqZl6Zbl6Q69YvYURV8xJzo+0Os624UyYWHtfIAjn
jjfmTlZdvwV4lvWnXJLcX6MBBRn+inLANHzUf4KvAP/G9BdET6V99v79KcGQEbK3
D167TfGZ6WiD/KH0u2g6E6ijrYdgVQptKbLjw7fK8zxuA2FfDyTDLHeCg/0bsMXS
RiBy/TZ+fjpWp3mzd9IWCMD3Eule5yKXSdyhwlqIbt6QVdHEdPw9ka2HZmBesztY
dRcK+s1UPhVDH71lUX1oy8fgrnMueaaNT39Ct/E9Ng/7qG5p3prMaiG59g6RGlie
8OX38iiQ5+BZkuvUhF40qQEKnShj1xhYdbpaMi8b+SlUkW5YBmmYu4HK3I90vDlS
LnZCAwwH47MjRKf7nBMfZQ2WJilw2ea6NgzkiUR8YAuQgL9xf9B2dpgN3pgNdnf/
vlakrnubXh7seMeFvVEkVq2acC7h6sazjKuBzW6Ywh321tu35SedfSeylShXXm6H
kkgsj5eqhoNChj77yE/r7BfFPRHY9lqGnV0DLJTi0Cyenog9bqSOVnQUGzx0KHCo
i6uZdSgkSMIb7ofTpbp1L07uDcqdyjazb0j5eGZFP/0UPEGJEcFAhmypLNQ0/Q6A
9Naw8URg4eyRZzkEJ0kyMT8S0we7CUDXB0ISR2mKMScRxNoKz2OorMZg+fK0lzpc
QYl0+fJOaH7GBheCbOk/OpbxvWilz6XdXhHhA9aOU4p7EccWO4SjP0XJcrVEFr6/
WjSHz7hLBrPy3/nSOhDA7ZT0HQhDSboldxajIB/ZZK5udQkiMnrMOvpoWDa207lZ
muLEK0XqohtRX5ttcoghQRkNHSocZyxcIWbfDdXA9NIwc2PGi4+QtsGw5+IOLUto
MHAf8mWOlsel3iMYPYn+IPV0APTlvGChYVJHlgSkHPp9SZOoj5K7Z7mpcwZSuMbz
265S7OcsfQi9IYiwKw5rXZ6OFtA/2xSo8tIMpuXMZrfoGJpdsyu+0v9u1DVvimrX
xYyW6WRd5apvie6xjmpG/RXk3fG4gyyWYYiipRzctyJmNita3vFcE49GfpJogBzw
q4KnA0Bv1nIZcU4/YXzxETiopPZNkb5Q6oJRgkYlcJh57U/l9gINfUDZfa7wrgkw
Y1eXf0N3SkGVkRDj1SkPZKT9BNeTBqYSuuOJUumIGtE9NpAU7WXvcg3uYzSjjDfM
u8gazF4/vOtXHvhu6BJNXs1TR/+6tU0WLhcP2tHZbiejcsJtUw8CsGJUrXwe7VDf
WKHDJnobnNKNMh1bFsG1Cg+3hpmVJyhnZ2B8rVTr8QtfV5CDpwUDVrZhc+D6U+6z
rvunZrh7R2kxluKU6eTS+zpqT1UxnLE/PjPsz9E5XYq+CrOoWgZMnO+ZVIYUf2Xp
6vCQm5l5QhEqBTl+8WgdDD4SAC/kYkybonw1hDdjSk0hGxVw59D2fXqHsjAokNBj
IZnfRtSQYLiwI2aSDe/0TLViEtTOme7p8aBf3374dxvVe0c/a+94g78Mxv6D6I3A
NMiAh+pgHbW9z939LVrLo5O8NfUVprHx5IZRaJUGNr102LmcAH+csHTKm+1cCMGH
2kmWQvMrxW2q/tz6gMv0+DklHorYUBGr/+A/uheZv/C0UNKEgc5U4gKEYz9KouGI
4RlIam8C0Wy0qdW+GS8Q0YIBDYS6BzoBW7liM03E9YziTlpQexMwWPF/LB4/xGSP
yBxKNnbvDbLman9EdwX3fxAPnHWV6XCXtcGNSNYAOYaTk3Ey67sq7X9YApW3DgXa
5s34LV7ereTO8bc0aRjNzwi+Mh9RAKQOseAJxR8N2FRbK9rbgvVHvyc3USUkmTO6
sF4j2UZK8Sn7Ts/WwGLJE/HXTdBKtZqFBHq440DaQewIkb72h0bDh6ZHVprdLULx
+EEBMMNFf/dZ66MWYruiySkhudgReN6HxOMGLtyowBDodea00o/MY6Qyw6WmU4zX
yQgsJxKq+g+6Y+/+hoYl6fUu2niuwGYjjAp7GoIZvtc4zca+Cokjjr++q9KmSIjK
ZMHngdPyKrD8zK2v6xabGP5GiEpASRSaJs5WYeKMzEOKsIfpWpeT4ieYO0lTcBlU
4oJ/WpOsvKHngGhzARUvG3p0fnM6Nr0fc/Sr1kwrP62ka4PYZDNnzUm3adn/VvWA
RpVtMNP2WEY20bnXpuSq8LD0zlpAymCUzuVuR1bj0GyE2oqS67zo7CP+oTyodm8G
vvPV+cOK72mX2oNxv4vpNl+gvkaMIikqetkVY2rjtHnGwWoLDRW1JAU05B5CCXLN
VhbFPsU3WqFM+uNqojUhhzKAnKk71N8KgpJGctnrkcEWtYWnu5H6GpNvZ7dp4GRX
V9z38vPOa6XBUa7bCJ+Tc05VUz1ZNb4oSnwTKbHBtvH+Rk35WQRGNWXPOo0cSQnS
y8S02ESMXANd1juqNIlUnDquyDqUhPzoiG9LgSio4g/sA7NpBvsEVeG2wHzjDYMd
HlfBtzWt7dULJ3e2y0dJh+75ciHIovxMW1v5d9RFYw0MP5TNMpaNLzb4Gj4fBoF6
AOiyk1uiV5jtXddi7MnaMBkUARbOuEZ1HddKgxumumJB2PNetn/BOxGa0O4c1ea+
Oc6D/tJr7+vRsJlqSiyUpcZk+V5BjYiaSKXauw3FfgCtBsDfyJmR3Qu6F/yus92l
ZuBFUrNk5XjVYh776ck1eEwvj+vv76vzKhjxRrrNuh3i18Pcg70QNTHHqXke2/uz
Xq5/RzBuz3d1HRyTF/dLzNDp2OSJ4YWCphZeac2tzfiddlFLN8YE9NWV7uVOlUmh
fgvXTxKZ8bYn8+TFXj9oyoqdnaLziWQbVtOzBVzH7y4dOY2Xj02zt8/kV780eX/H
XFpQ9JHAtv6WHlgVl/fISFuEfB2c5M1dJ86gYX9sLyDfUSD8cUFqUcKHcDxTYrE3
pw2FEdvpREHkqanCnpANAUHDhgap2J375bOuqcOozU45EyKgeEc/jQC46pyYwE+U
JabnPfdH5sYiD1yCd2GeQB0ym0/CT92J6GhgTmE/hiTU9lfuljKNkjFnzO3+HTw/
xu42gpSJrkESKXpxJ6/nvdQyWRrPPbxiOqYs6VbjgyESNRre3vPnaGZ980vaiNnD
3VkWCFqHF2Ix37Y9u3qomFKgMJIurS0QllAstovfiPC3FKsr7MJyxAxzSNH/AgEh
TzHMYOK2QL4qzNoGL3vpQ5SiQmmwmWnM3jLQxYL/QNMN/myGvX3XAOOPkqzbIa6W
T4y9OOaEbnnDbxaeg0SH0XL0/oc1n4AcbNFL7xEDCCi41isRgcdYGiX78rIFymy3
bo7rYTeJUCg4Zv+jow7XIsh8+rvSA4EChdMpOWu+Q8HMZqAK+q/b3MKEUvIiiTBx
6LfB7FH/YjM5gc1CY+1XNLU9qCdTsaKE2vYEh/MGoEeTFSfxiUYnhi3nsujWmh1r
tjLaob+bumGOUVQIdKiu0+8EsKumLXAfAWt860s5JhU0y+7hB0IMajwchbgoCBc/
mMp0W9uQniKJi+eeLlRc4KNb0r7YMEJMl+MYwygV9CWG8GXDb8IwKR/kJ91B6Ubg
eJ0KCvlWJkEmFtHpKo1/ArtCZ7YjC0AEDGGkIaIw0VRcA37gCxB52oQaosjtgfj1
EBjtXUWCyPXX7jpRZtkghvteBvj2ugFlbFBtBI54JttP/J2xOgC7q2mPK09/9k+u
mRwwOH3zn7ud+SpaHQi7TK+ogF7+S4eNoWVkR7khuu1pbwbumP27NZdYQJXa92Ku
1itBoShbnbNRX43dXZwJRa6SVHMOZTQbfYdQxw4o8bNh1toSf6qA76I3v5ENGrb1
9GLgOX4tgArcKRPse+5Jz33w9Y/USHwGaJVXPsJCkxFImDi2M5n4t1gM9P66rFpO
sgUCYFML5lq1unPH5j+M5K20mvnwVrQCPiyU3KXamcxjx/OfHcUJrEX/KTp/Yk/p
3LD9+wL9kY/Ci5YdmwSwQLLvBc4iUHh+AhHE9Owfgno2WprXwkeMUX/9kWSBiV7m
7abSZg8Po4+WjPsG8v/qq1zJhuEDEmZDUqK57+y/4GYLYkeCcmLy8Uw/nPUP4CNk
T2e89HKUlSldWDwKMb20R9+2JpnPcA5FkVlpxgKyLcz+ERP8DEMM+y7jNKuoH8jw
6D+uob+XM82GPjnQbuNwn10z2NYUYQ5x4YBzyFKthbCEwVW0fT2qBEhTXR+nDIwr
Zu+9a54rtDqO3oS4971Sy/gv72ul1JNeJEu0HvKA6MYmRf8mMSG67S0TLEDTKVE2
BZgj4Mb5uZkl9N8L672oM45Bh/FNgpnR7zij3WThTDp6hDuat5JyZpoNavq349ZL
LWOtpvpUGC+eQw3YRJ8dYtvjtzZ9vg0a7F7cCQWBeNALnsJmTRjcLF3Zc9oCddHg
iFtEMxBLj5ePShQBdF76zb1YvKaGIW8ejziNs9iyBqMz4xb8srLVFypuQ0H0R7qd
TgrwiysnlllaL0PHTgq3Jy7cBN+7LhN0O3SA9UnYtzbERf1zpaIZTuECEDMGtCz3
OlVdzapoAKzG9FjVT+BfG5I1Vc6Q1HiKE2tNL9dCBLPaZAByHWu9INH3x1sMlfpi
zW59VZl67cd+YLBzbn9Bpi9Rpf4KGN3lZuYujkmLY+D4VH8u/aibq2a+X+v8dDJz
XvgJ6nnnVIA/GDwgx7IWuu2vo0fKEa6S2ucoTwgRPPM/k9HmSIDyOfDdKDaf74oM
yrRIkvIk/fHZdCbAZG96Q6LBa9iYPy9d6YyMSf0Es8x48883QjZlV4eh0lYriaIk
bfdbtLU3oodOoY33Jd6nltdBnZYeJojmA82tE9MIadvLeQEQDD9SDLVxmWPSXvvS
SYB23hrUCAm1RUXLtF7QqSMs8KrhZ1x2mOaUSMNcZpIPrG8YMt3vovQnp1nvIXbV
4WVh0x1mB7rXsO1sQwLhouwqePUIvBNixz13/wfVqhkBp/5hCOIRq3OZyaB8UKoR
QrQ8dcFRGtO82hokcgw+vfe3KtR0G1BDyKnn8erqSrIeDlp3dKjLS78u/Bs8/lqq
f1qABQ80oWCfo5L41cvLbscZ5t0WuyzTw3+GiDPA9so=
`protect END_PROTECTED
