`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WtN1GMoC7NJ9ftVfQD8r15jSRnPiBlCLvok3DOArthBDCB+feEy14SthUxLpKYie
b+0zBkZR3gdTAS51mxS7+MAMRySLsTlxYupi+axgvEmTmEheJ0I9/1gQvqXbMLHQ
Wzq1oOmqZpJQs8hSyL5KSjvT/nt4j0ro8m+M3I6sQIeBiYmaaa51FSkaI8pOLowS
CP/aYHZhhtczVC0pQ5/+/Dm/wys5iBO+ucB8MUMfLPXYiesvquDhdfsgaeHOURFf
WeSYVCKA5gLnu7Gf5forEq/UaGZshfNnmzCmXhhXWPi77WiPg0cMj/McsRDIWgxw
CndcJSyhCvJQ9CL8dBnRcBW+VPFncJtk4sWXnK6VzzJU2Okip59GtvxZMmZeviCl
52AT5VKC2N32VN8yLd8HQx8xPGXWvqljiTu6T8YJwMQMBEp+zuV/4kwkFFLe1pH7
w7kItddzsVIk92hccz31QFw3BZKBkNxnPzLw/uFa9ydkpQxgP8pd9Vn0L1zGwKB+
DBnJeeMiI9JAtJvwnoiKU9X1ezL0BCMvr8tdgZPp+VlrXFSfDmFQs1YaPe/rbwLo
2EavKsUSetWUWiah+vW5tUAQqKlig/jM8R9XSGay+Hi73ytMrMv/glhJeAxtuIet
GTwccbBVH8BAmyQVrvdcufTWgeYhBplRsBRZcpfDEmaiIgkzX7RtWNPpKF69J35j
jRaNd78wzQLfT7H8fydcBJsuswsEz4XDnxBvGB41U/cD5/S+Di3OnWaQawxcMucD
rkA+d3SR7f3Lx/VlwgQ/9kVSX2d/aiCq6u7GxH01mM5SfmrdFBKiyxZgSw9qT1gm
0QNs6ZshmCsnkV54lO/8qjSnKyBGRTGlAevJ+374BgTd9i3V0Ixf3kQpwYXi8Z9b
MmR84xtQRrtZUs5XW3kEVQgpMgI7c6CClbVQoVCF7M57WjumKJZH5/542t7NUWp4
/HStzwcpZu8EpRC9Iy0dYjXx1SssC3ULJGlNqCfZ8kuGt4bBYNgJhk4NRrzNnrB4
yBvArocajODVQSKsIOrjiUP4be3MfkuF/W+p2sX8sOvIfGPMp20m+t8lYh++ly7g
r0Q8tEQD64EFVOEKnxSTBXRrFmiJKbOjF8BKzV1oND11oBOZUW6dKPdBaWTyhpKe
TEop+WfGduSETNGxQTGJgVdqE54su4vzV5o/NQ5nZaZ4gCyCs4br8Oovmjha4jC2
P+UoCB6yf/wQWvUXujNp/+zdVGgjpiAg2xM3DMPZpy2LJ6O3vtqnt4dSS4irAZqk
BYpR1BS736XzBzZyOw6/b0nmzjxqU7axkHtJEQyHDHypD73Eh4/YroRrbrDhuA7i
yFojh2YDPn/YKW9XKrcmKVH0a8Zk0r7VlgtcBB2Vtu4PnDTOF7uwh1Ul8ODXpXWz
`protect END_PROTECTED
