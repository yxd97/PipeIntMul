`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ckn1sGXbTHOJJKEdk53KopdLy9cOzNyB3MxXVN2Vl85V33IXQ4iFly9oOZ5lFBT
QtRQNrtm4XNWOtS/2iNKiB36BaIQMxgHOjSiWG1lnIzjw41fA0v8gjpdZVKMpfVI
VFOW8jdvbOYs/Au+kbvadqbhhUnj7lyooDUqdzVbc7hoNVHUTbD0wHmXbZsoXYcZ
9wVs/Ujk5Jt85atglq5Qlfitd1JywPovxtv5vzS38zvXDGZWQ6YY6kskpt4PVvEn
cY2kSQJnd4BA7zcT5FVisFajkbxyb8s5J/vlXLJyG9w5qjS0jC79D0MQk///bofB
LmDpPx/oQkkK9wEhPu36U1OMOKTtLLuW3vKJmxqAzI9t0RW8Mjb60hANZ2IvJoeh
DfB824Xb3UfQF+DkpPEFt5VMImehzw0vD3gHTrgscK3dox2VS9m8vvwqmKgzT5gL
6nrIWGH8J8SLMTr6SaWeu1qbptQEfeBBivUv+h3lyqnngX7FVwN85W4ykdPQC2W7
6bjFJVPovjg2vqRaXSQYYc0qLRuwb1w/QhOEEomRU4x9htOu72fG80lZpX/7THsW
tVI9PKySKCfszIZp9hZaqw==
`protect END_PROTECTED
