`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fTu9nEI9xOQatBjl5jqMFmgQhZNDeuR/kCFBhW4mzU26mptuROnyOmOw0N0SBo5
3i9CgzO+5lAG0FMOBrbyvEzC91ne4mYcM00qAHKsitl43WrCs9RjuVA7Ai9J9SAd
JZObpKHzTGa+pNeyhM7YAW2C7Yhi1fUmnfBHb8b1G3hTm/QYVFpM8+xXMieu77KF
bLhOHEI5oZiy+TUzk+77vmYgiUN9bUc8Y+5DyIqqqwP2td5VWj4jaZWYyhCq+lF1
L9CI7ZzZOMr1WWRZ4NHvdxQ7VLmhrx10WJQy4OQUeBrbTjI4OKAhsfMJ8qVFh4pR
fRqXPE4VFlDxl1rNz2z4o83XXsKCyW63rbIfikWbeuJqFGKTIn6naZGUxL20GDcj
QkmkINWE9b3NVhsT1KguEVQbB83BigIQSB1RRjjaxh9ZBemnX8ypM87J4vFRs2wv
lFsgBdeVOgNLWWR+9u6U0FAu37olQOkTyczTTz8achDc6zXE21YJlcmIqO92Rc7i
my+w068NfiCGluLusP5oOa1++UVCH/UaLwLehG8cQpOZvArXfTqIxEr8JnOuJFGP
Nk6+V2/U7bShK15cqb7L3lxcr38rYXGhAc8qMnp8/VW6Hs4hAI3v8uXD7hkZ4vD5
Y4HHUDj0uDvs9A131ZCFo4KdJq/s7L6ajhtiAfmgETAEJ61Tj4Jx8sIr6e7IQ+tP
mkElOAzyIeT9M+IMSyYPTcPDPQBe83IaqtwDitypjJOOBFTBYOmH9ZSyk4cL0H14
47J9XeScBf5M0zq0MUV46v8aAufPX4KoWVfKJAgI1AyIVfGB/gXyAiWaVLq1z74G
/V68ollVDE6ybAv7oN55B0gbSLCrvDbxCCAX5ev1CDpJJHpFLqkkwCQ6PC9KB+ZV
eE9gsRltqReHz8Fl0+dMue0c//1RFZ4Uml2POuQElyxr6VOq0xWafMqCLNd8mMmE
yQjnYgprx5J1aKtQKMYN83n+4+Y5bXrMbXWkKS86eRXr8P/wDNkgAle5nqXzBDNH
KFCB2P2JNE5uhXw5dZXlOu/+lH8qOGI14Kx+Es55umkfynpfeBObVUzoDaxw5cIi
789Vhw4LrI29/Kvun8pJe9mnD5V9in/eJhE/jSrmVSrQJ5Ko047fMbgPM6tv0Kku
v9lpIzwpk+HvYEuiv52FBSVyODwbeKZQx2a7LTqNQtXeAXBd+N/zE/0IJ+4XBZ6s
2tRprIys8bUAXQu5XMqGNR5yJPB2REZJXU4FeWaD03fJaxeWT6H0xKWm4qnm4TSV
qVvpjZN7vABnSjMwAUZC5/c7d7GIL2O8CbTxe3cRh51YHCK31JiSSJhiUHipPELL
EbFHEi6K/iLdQ8W/LgYVUm/kIKLEux1h/qMWdcbhaRzr5/3/zJJBg+dURWUIeDfa
ynQtUi3t39R+UotUZVKO8TdVvvg8aojnoTzf4R2mS9sN6+L7fpZXtAp24NZ1GHn1
+xpnMmrmHegR8tzY4SWv+j8kiIOHAm4rYcGoP8MOKQnhvOhidBfzas7Fi0mNuTHj
7I/Z6AK71/sWHWAw++/8q8NIFt8NuK8TFHShUyPWuA4PGM/0REi3x5NwUY9dTwIx
GHkyeWVyFeQcdTKyzik39ez9THdsY1+M4O/ma10dxmFC/MaISJ15RGqB/M2pmdlA
xFw4+wYI7mRDWnTUoWZa2fLrzZzPk29AdJYoJ3zEmGek70QcWoXFQi8xvLqUmYez
jQelfcZad6ikRw42EF+2uw==
`protect END_PROTECTED
