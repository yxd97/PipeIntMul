`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHU6+tlKSi3ZQCX/m2faD4kJQyM53WrF6Vxg11AH3LDeNYTiB/nTiMo/DTGVh1DU
SYMzmxehQiC1H6MCZr/LN9eCH15MLCTE6nsE2mEZFMom3f/6CeuHlcD3jCU94DHr
32ohqxgIxhd2XZmmCaMxq+IopXibjf59F6/hqh0aKwL+oMWbFYiww9swJ/IA2iAS
CeyiiRt8N7YmE3r5Y7Mj80ukNc1UgH39j6j8xbs2aGBnoABocT6z3nLZ0V3mzeeE
fMKbbOJENUN2kbIfbLAxeZ3t9XmsaXp/d36uR6MwgX1yyFltium1sANq+V9yyh8C
Vnkk9iAHVZ4kksey0sydyzbQ+tqKhoRquOdo1p+9kFiziQSUf58puXt7Z+MCRegm
q1pIxGvY1tFSoabC5xTQcdSe2bZCsTucdpg/vCIHvznIknkpp2HBcNbJh4ZcXY7I
EG/PFXjBd8gTQ+gL9V8zZtMtMusA3xgOMHzBbNNoI+A6UIaGVMIIfdz8tl6uSz2i
tB4PcA+ETBV5/ZHwKe9arx3F+PfRzkzwkwggBvKcHrpWbsOyZ2ggzdQ9uuAibe6V
WYekJ4idRVuWY+KHQpRZCX+8+/t8nNQsK7GVYTvdd/HEixQN2V13t6jgLkWq2eoc
Tt7bMunJpzASyhS5vge8mIKoRxvuC8hh00SCMQ+y00+zeVo+XoVxCoZhau6Rt6fK
Rd344UsW0XQC8wOilo7sQQpo5ciWY3loYmmo3ngdzaai4YdGh1j+HBBReIx4nGX+
rC4MJKhcwRw9vFE00g58OEY5ez9PtczLIf7ze9ZjqnztXSjKt2MyCwIkw+tYHe61
bUa62QnMMocPUk2+SEjI1Ac3N2B9UNGFjH7l16Qxqt5BRyXG2AppIcdEUfyd5yBO
vFuDHfUlzYZaohQme2kSJJtJuY48FdxifRMSTZd2pbBUfDSf2JuSadv4HsnpnIZe
WaZ5fDyY6CCrruE/TCMBe+m4mFNpQOgUrHd2eZCwfy5Ee4bKSuE5X6IAg/hzXkkJ
dP9T3+qsNDf2tVPDyGkFn3pscIUI4LI+f9scTMekFu8MLhQs6Ggu3Cwg1tnKOUAH
0/ZDddkhkSsd9/V+A0MelP/JdCauvxt3bI4yIQ+aoaeSwBgBuOeIqM9kvEyszY9A
8ut4iWGHo/EqxmJh+AqAoHeZZi4hd5IHGM0B0cm1/B1VjkrU2TqsKANZg6J3/TzP
rcP7nHIHwJZKm/J2n61q4HlBVUTt9IbcjgO5V3ubSjwZThD24yNjUmvvtrUo1bLr
DzwrYwUti/FMwPlZlNBpvCTtyy4CM+dw96YRKCPQRU6al0a1o6sjEx2Ff6LFk4/B
ssgECHocaERpyvsoQWGArlk5EHxR1H3odWoOGcfi9dGT7WDg5yRxJ2ao+1ZG0hlK
4nswGVuAPdXQp3nUfZud0B6PRdF9eQXN2NbZQJSGs5lYmsr2HOqOZIFm+ILXZ/gp
U4EIUnMQ2XzGvaaI9ZPTA6YkprvHOV9qv3mx87VoSvj3l9rLlR8bf0n0cFknjtdn
emXY61eLjoj7+OUyJOlS5jGbhGX3FaBXkjMqd4cpgPBv2DHHfl7NbPAm8+jRMtZW
rDqcM6g/vjLcgeAHR775sFeOVBG+uh2YGJGcX5ime+L0bYbe7kDffTU8NN7dvqi+
y0d3ek8vbrUep8vBm0sclc9OBsLfnFEpHnLAj9gkGiF4QPoisaKAiaLfr+NOOtp6
SW4csNFcI/NF5BpNwtu7eg/HOvkHbTsftxBgkoTTER8zAj5KzpSLJL94A62keavA
wfvRsOMq6C64XcnqWGCNdlah1vh0jmw3+JBhkH8Wu70jp9s4o/rjNo32bd7hgCpt
lUC7pqKV+FvRFFGNcZDG2R72/WJvywL5N3uLBaWm0dvxX5UNZyQShHQHp0ECxwTt
2hksa8bdZ/9qfYdZ2vlX3RrkQWcbxx/jdviih1n0HmbvimK8TcTQwsZaDYcu5sKE
KIB+zLmPFYgGe00Klz69l4foB8ewqgqobrqX5hRw7+kFSEnFknZ4dlKewR3WLUDZ
AbKdq4N/Mk8XRgi3zYHDANRzI5BVLtqr4Qsw6TkZdJBqJbCiMhIBM3lM6UzjA3iY
SDDs4cXxcd2h/PuVyElVZFnj09ggFb29rpu1FlykDAlNz2tCHPMuNY8kXiCrKT/6
g0/qzxlFJdONx/VSvioEdNzmWX1hMZlpWAytzG4bO6FO2WBbD+Ki2ZuqQJx7saJ9
1G0JXZwAZWEJiVNXzZu41/3EdvZH0X/7pijPTdUjTOvrCfkzOT2kqLcSLCxlr46W
lRkgPOa8O1glkGcyhWz8B2W/lIdQCII1teTK1rLcLDFagjMtNvvr535srkXvHUw8
xS+HCN9AoRyAOZqpdGeG8JhjVBJgBFBGkJsFQFCpQ3OGRk/exSzsAqDFeyrSryLW
URP5isteSXl7OiD6PvmVym9FFalKVl9w3JgiULS8wuiLtOLj2L7KztSX+IrTp1Qu
jMrgCrpQ1MOfK06DabbHiIcrI3mLYE37XCiY4AIUycJjjEuOwXrLFnlcDJDPGsfX
cfrsLbPTPTeQw9awno3XmjKOOJgj8bKAh7WvyJ/rW+oTV7z+aIyqwtssDGQrMluR
`protect END_PROTECTED
