`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ooaMYVtt56spFXj6xN06K7/9BixgLlVMWELdS+lUfv39Y7fec8LJ2M5cCYtBRoS9
eE+NKY/pF2QFqdkhB084vFvIQ6phtnG5DF0IMdpCygoe/Wd6mNciVvFYpzh9tg4u
t6Laxi/igNK//5XX1FGYt3cEESYwNS8lED/2QHnzt9ngbeCYU/0dKOi5bg3TV4p3
A4U16pXdJ5pb9etldBvbacVbkRN/+MsijKBayZhByUZaidLXelKyTYxnxiKSU4A0
9qBHIKBbkgK6DFCW7MxLN3ZOrz6MxaRmx+zXWP2ka9Z23X8fsz/M79vucx3/Yzks
mg6mTFUNrNrUrDI0p/WkFteAjcARyINESrf1AhU1xY4DrOfsvLxW37xqosfCMfT/
qVH9nMst0CeEVBbD5NMxn1t4zHypDGgfLcglh71RyCkEwOTG0WhumnICx42LGNfk
iFxVzWvmFIPv0BKd83LZco616Kzd8eYxOa73kr4wo7dHV+OqmQhRXTJzZ0u2zQKP
Iml8q+Rfaj5KbRVS2q+wi/ns4NZQoP5fRLOqfd2dX84lcO1BnRCNjuuMrF9qJzCq
u0Zk4PEzNveJc5qfwl9av1YzmfVqfweEgNEg6Pxa9icOWLQ9hEkjQSXwupoiSoPb
ELMe23f4tZec9gCzALz7Eqc+HKrS5MQjrXRK704khKaQ4CgMkSTXbnODWmYUaLf1
wbyOIOiwYJ+BWSZselnFkNIHbBPgRRqIlGAPqoLeXymFttX2mSSpJG3qlqFgzqcW
Jz+mnNzSI/pS4/IcHvl32CY0AkE6LvXnp+jjfs0J++OL9xP89Q7Rjhh8uAQ2x0wd
5u/uxu2SDpoQkL5daSRd6ESUT3f2RaerZwm5JOFy2C/hoAR554kesDor+4NwKQdO
zdJyRd4x8NPyh3ilKLyRSJjFV4spkzQkIVp8rsnwiqgYUTaBpxAibQbHVUZjj4rG
jh0ognfreSxl1CTjMUg8U/CLHeZAFt+hzHRZUujKTmJm29bkJC+vF47Z+tPrHVxv
+RQFL3GvTjRtMFyZAZpQyWYiROFFR67PsJZRzewAfzJoLx9KPjKp6JkVv1vrVSAG
jCU2SZVWVsops9JINML5MuZSCzBnBVy9YMmIeHOtTwcodEMiS0rC52Tqw0GplJad
phfdI3cdWi67e2MOJyxE5Z3ejGjQ7MIx7sXI9cte87gE2ZEa0xn0tprpbbCMaq4L
DnbGw8p/u/oB+d32RdXnz/KsIIIgkFf0vifNZEOTXa+2Lc5kMh1lj7mvG9nyVwng
OI3MSTLimH+z8hr3UoLLGR9uNKct7XVe9otFdEEykG8mk6Fh9jlWCci/efx6HkbG
61N5SG3ii0YnylqX1WwvcGi7rUWG9pehcZyIMZ2XbbAE51G+lvWUDhWkOY+uzFoE
K+Q5SoKhdrhB6abLk4+UtLQKO6EIOZscFrk2YyhRcSdkHL+2jD9A9l0Mk8wCQrIi
hlYKwkAR1vEVjYwxV+cRL4kTddlJ1Ij5K7UKsMhuzMg8OSe0OfPs8AjddATIfBOI
7uxCqZyXPyiO51rlx5mmi8lm6L5OHxA/LJ0bnnfzYIRMiG0ZsH74YiVxFL1xCuyp
yaSGd61dlbRoWv7MTH+V/VnB2TWPvJRgRWm5+Uz3Ef8F5lzy31SO7oZRVrjgxfVA
9upcZShryAPosY3SxwK5l1wVHwyednCrLHS2uL/FnALNagbvJxx7KMdDJ1ib+kps
quSXnO+u5fXGA5orIOZcEgwesaQTit1Kl+Md3+6sEfkGXQeHUvVu3HxLS47r1u+D
yO5y4Kky33v17BwDdj4ZlwY1g3iBuaftTqYe4BNGclwvBX7XFcghyINp41YbLXMd
exT+usLdc4NCMShmfl+/nvftNz9hL3XOcI4tnUCOB0IaNg/77ehNEglCHhYzgdeY
`protect END_PROTECTED
