`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L04r/yRq0sVGteOxftqcKW8es5g9Vq86PLRjMm4zuW47jvkTVL71+3GT/yyPlIfr
TLHf7weVMJldX+qguE0DbxRpaehqT+9VSeoeD0KK+jnvAEgaeWJ6jgqdfTBfWrO/
E+S0lcAcmYMiEgQ9rBlLQ6DGg32QXmN3QNLrD8GCWclU5Pfzf50P0P20C1HPVoUO
4nzmMm+oTKt8OFe832v4WwdayaeBThG6eUwe/KzfK8cHrfs9WGMR4z/8o030HJ23
rMafdl9EUEoO3SwxF2T5LLo5izF61QvHQIiDFKtK6Shuw3hMR8+Mt7+M8HMhARbH
tPTsxdsRLcqIl5csspWE7hsBmUWfFayMoIBDOTI4DyUUgJuMLe+bXrstBBBP7GJz
AuJ8EvEIX9ZXrSKTKAYRBYn7shDFkgPn6UBqwJ40Xv2rDUPBYvJzAcLGp66NjnB8
6Bzjv5Oxn0vwA78WxtA6HUY5xpDeo+ZR0rxvFpNk9wwdbU8m+qwcXc0u5WaD9ec7
i6iiN8Os4+bEVuLftxN5pihhS3nkrRNhkbugvzN+E7V/daSUEE3JL5BqNfOtgJrL
ooeL6Q0OUM6QXz6NDsdAX754YaXXSOt3iAtHwjbfxgFwVXdc5qDToPkZR9ByVBXV
4BTXTdTFZkShrih/pd4zShTzN7m6Z80B9cc0t8CmWAgF3OCDkwGDx6HLpTCDJYZ3
2hpkW85f1VGYxPU5bR0orPayXz0vfeBFk5EygTARaTCg00asWH9CzohQp0N6y9GX
QSe/QjEvT0wAVsbLbB0o81oh6easRC8oh0gu66ZdV/UFkwhZVuqU2Eg4VfugYMBm
YQy/6cmn1PnQXY6TWJK+gy09srYCZ9xTLgQ7lubqST1MfrWFTgh5OW+/ur3Sczam
jx2M85Urt0f4cwvFd5Z7xvfBFzMYM0sw72tXbL0p1Stcf6+B+3yIncxMlV3jPcT5
RgoXfwYJ7sGa4liRTHFe+OHqxI9muDYL5hhXIcolL3kWqm1MykwrkwfpOwWJYGlj
5MEzHFyGIcJXa2XOu6zb/To0YIxIqNDfOswK8hV1x5Bn+wlZOPcndHvwB8ZkQK9H
/p3r+XDmo0yuUHEJerXAaskXZZQMpm+SLgaGaUvW9Cx0mu9CIqdrqxU4csYV29xi
8hB5zD+6iU6UNXfoKZAgu8sqzFSRJibFpz/92DGCx16mWcU0PMQDEMpAnm/pV4MZ
NU4tUQkKmVB5nRscj12U1O7ojdNORBdUMD75youGD0+b187QsJkmU6cTheW+ZgyI
2anXt9nFwRyLyd48FbcekO6RGfE4v0qX55KUrGHIk2b1J5kkOy9RKmw4sYXy/U0A
TGwhnu0/kEgxF87vlz1E1+QfZEg4VC+K2xGYcyAvMBNAeAC8xuojiHm2a2vf2joK
lKZbcFFqp0MlNZXano+RwUGaa2SsEK9zlcT3JDaTnWCB1NHMsxOcCFBBKyr9H5fH
6lAMKvOwSM4YzTt0jRmfgcOIh8U7ye331PHYZe6LsWmTTFWeZgc2UKD14RthHlMM
QVLAdEoUJSy3fZQft51JMbTCiQrJ0Gl8YWa0yLGGXiQoaanu2aBXlMyZZqPky9LC
JrQlfz8k08r6iPvkZXvikuujnkeYSXvfbofg5eiC2EAJHgATKRGZkR8hwvh7fu9v
vGciWnf/gAb3I/V31Cl800KWXyNOrow/QtPEOFM/bj1laUo/dc6BtozBcPhHZ6sV
`protect END_PROTECTED
