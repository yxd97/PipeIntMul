`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+to/yhyWm9J1mKu3IB1D/jn96Yg3sNfPO9kqlR+E2T91j+10Cn1un3Ub4xOAlHS
TK8wYUAoEe3jpAIgNDq1dg4eCD2YqbKIlF7OaG2SSnDaBBAEVhnGs4bk3S0ZQlXT
sZE1s03Q1vaOinBXEAH2DF6rLfsX727x1jzIcY4GJHl64rbjHdPQBA6oyTsx42kD
pnE79ub3x1EjR3iT4qLLI2Zz1TWPI24iU5zerrXMV+V1J4puvEqDQLlLeBoATmgz
tk0Nks4bFX0De9AoYiWlUYGiCRRRgll8ZbpOPmZcpSwBLRyPIeHYgp2B88s85i9/
ZyGMGOu3WnEFItOJPd6ab0oJi7huRbQ2Egf7nI/f65O7Q6lR/Ws1gNjkFBwbbVyq
mq3HCOBmjpRrqEddvtGkb10jZqsC7+JWvf/ZM3OTMNOS/Euk7+JbThKNgpAVXmPA
TQIh1Nzu3ws4eQOU3O1thAiV271IgPvFJMhdPJ+ol9F7PdLE61yXg6dqnuonxzBB
eJRrOe9aqibQofOI0nu1L03sL6j4tz337g3XAdQlIkOoDjyBVF95o1AObHOwnrQz
`protect END_PROTECTED
