`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EyhCY0iJEYJTTZLZPLNNirLPvNnjJ8ln8ThRNGmHXiMwNmK3tm1I0Wmy14JWja/y
EcevFRNEF0+98qsiS55aEiqPVodtP1543zfMiayc85nIJL1YUt9IvIDl1QJ7ffS7
CbyFkyuFsx08GY9BQ0pQXgd7wt0FK1RrTaMRO7jxUEnYpuiZwQxeXHckV6z45kOW
zmqRX4G8oGXlP1f0Bce/0xSPJSrqYnHwN6FtPjldtxTIqJ8KvowNOQ6A7elh3Z0q
YfzLXDiHIjZaSBx7pQ1KajaHmOvVuYxxYPFDOWIzlN+MBtofLuQmEf0At6u2JsqN
C7IG7iArPRFxLJIqMVIghVaciCZoUKPCVR1CD4KbqHNVpfQHBzGAqHRGnYBsFfqv
bGh+9d3upfymAWpirNLFaGICTyVxMFK8suo6yz21WZZjYgXllnLDOSwBteDKFUFz
dleYA3zIsVERDIIzGcywuMacYRrm8K6Hlr/WpjZdg8UxS+vdJ9E6WdBG9pRWfEml
exUM+Se5hssIEEN00kiJIq4xk91sxGc6vyV7UwiTC3d7tmxBEwCyOV3IbVKf6AhH
8sX2WVKxOhwkKOaNG0ICDVhu8wtZcbgw5TyMC8fOvTW8aSJ0U8tXtL08UOfPMn+u
TsIjARrZ2n3pgYXJKtsEUbgWfbSZZ3PlfeKv6sLHCVVUrnevZzaPWY8O3zl+Kij+
mEw2YE1EafKheCIJSUu8RL0M6V5IQcZFqxfFKx3hpcO56waAuFT9hlnopn5yDWuJ
oFlGhGCjuWWcrHaYDfh9vHshu6Ysc4E00tIYotXQkzijwHWc5JGGwQAKTs4yl7Vq
FoAib8iQOW7mlchGt82TfyzpHGQoDs9zM3F31A3gu4UI//SL45ln6rPQMghVAwVI
LCxNjGy5GqZJdizgKOUwWBB5vjtqf4bXLocSpI+Tvo5rVFlSmcuMxCrnQHO5Vb++
VJ3wNeAJZ9ototUdFsRHNm7Zr95YGja1j1h/SCZMR1wfa7wAF9CnpuHOlkwvrpi8
6P9KuAdr06G8Pcqictt7oMw6MZqg1N6am2w6BkA86m9nC7uOd3KX91ZvFAF2zAW8
9hj7bTj5497suiX7DfpgQM1VdjYScnnDiOk3aXOKBuFMW08qg5nOWsh4b6dvuzJc
ORIXt6Kbtv5vk+cSKOPnIWEbYX2p42DX6Olp0ClFXxn38ytfYfHqS81sMXsTbB8P
QYcy4gbJE/2RTXB/uSvSuDVd1vJ1huVtub9Z6EAls4MF9pI6+wZarrHinHDgFkbj
fNRbnLYIwhf0cFaW5RHf9sQ128nkgajCnbMEYqKrFdo+AVBpXKsGS0M+yiM5XPnp
St3gjGKPbsadtvgx9kNEOKsHhJLLWhtvSgUhPkL3B3NdxIx01Ph35IqE8AYGlsAw
xTBCu0t62lI31H09anM2L/+aVua3wFuw5ATfYI9ksf+F/Hx6digrfvA5MuahRwGF
I0ZfkGekrwG2Ce9iZB1IWCbTG48l+cj/VW7KQOjI8A+t3NXfnHcV8Bo+uywlKFgd
d2CnfRiiw16bqeivo6Dd6gh7JZPMYdqMwlloUYq/55uZPLQqhUd8X5CdwRmQ9nnh
SuuVli5yUeARAdUTZ84NMbVUuDQpYRh0AmpBZ2vuSIzaW4QczHoOcJEpCqwGe3lr
JqdhrXJrV9XCXbEiSIFmW7ma6RZX7AtWhckmRzt7RERzKs+YrXrO52UwJv4zEzDk
1rwE7cyH8hW+pVEITrApN3l7yQr7aFzmQSKHfeJ3Gh0ocIpISL2w2OHqf6UTWVmq
VINv82siv1XVUpYa7MmO1tIzD3MKNWjbXnF1L7/Q9obVrM01zpGI7zhRCAUiRTPT
vXNjvpz/kXWZokIqo83Jf8/ijfhtP9RD9pISCWugRh4kq3StcoNt4+nZeGNyJYe8
`protect END_PROTECTED
