`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFs2PxTC13ChgYAOhjmQj3vvMdiXViQPOt41UYlw4WWb5U19uWbUlk4XIEEfQ0fi
RY1kYeGano+tdHcmxuFOQ4a/ZDx91ntXNDcvsMD/oqqbRQLaOl7bQ0Wbo6+OBbSO
gJzxdhtaQt2nLh78wWeIqwMeVdEUt8JAMS2PwI8O99hFAci0047DKQUtvTzoW1ez
mf/xXOo2FusG26YLEtI8o+VA0DIkoTKFEf8ZAXr+Diaa6JddiW1fAyDDOhjPyHKR
BbcCCw6TcIoKZ+cTznBRBpotNMpPt9KZQizUZ6j9lPtdSYfDlZUcZ42/wnAlE5lS
vpnB+w0Sr6MNxUAD2bFSbiLCY95gQBXvT5Z9a97HvRdeO4DRmix5E1wMpJT749vC
tzSwYjGGeL8sCBW3+5uoHfJEfVrNuWDlp+4dTLyWmPIWwiUQvRUSWKZcFSCqfTFS
twRWMZRXHQGx+A0mgtlIwu1ydA+CSLqjrnfgbu2SUGNGFqjPsoqFnAQJUrL+8El5
mzaqbEBeAIIkszPWrnfyq8vzMpke59oryqzoxU9uAfuDl9vfeGVFXBZxwhpNxENi
aWmezxYiYfGoCiHTX28fIhqSoxe8Pt8zR2TmKUVRdBqKmkczVjqjfbNgwPBV1FaT
QIyyXrHDe/K5LY/YrtltHQPO+3u1fAe9vfN/dUQESAwOhM5NCXz7vhOsghOS9HJ7
zWLisT41wmzhP9Vlkx3oJ1+J6cK659wMe1ToeXnHCZIi6H89dseRVbZwHDErod05
aaNtHCpAuxsDCHcho+P5+dQmkWuVjw324s4he/FXB4OmTRNyAvrDMkGbjqi7yTIE
D25lrAWzFQYcgscL22fnKV8+bk9G4sJlOMfnX/wmWDb5yovYlNf4+wsRKSIn/VrL
JP8Em1MuQPZ0CmHkgHQSyrxVja9zJXOB3An/rjm6B4F7cxaYRsMz2FAnlNnVY8gM
/XBmXBRUAdY9oJD9TvUQpggCkzLFmLrUZxvYNd9YGD7ZXDLzXwTaq0wwsXQKugxY
/IRzwK5EVQJSSdoPAwl/7JIN3MEFI9OBLko9iP4MgA2QmIzj5NpGc2idnc/vIOcI
WepIDcB+5FjkvWqy7YR3l9LrFeiOnlbPu1zEIVGscHHDVTk7v9EnvphWKwQNWID3
NwILvGuX5PclRkk9HgTBm4FgO171/II+j4iN9XeotEq5gnXEtx/tznG963CZo8HJ
1uDyWwEpwPLx4o9Po+frvhzn2RmGuPqy3/W7nWMzdE0LLvvS3eL9c+cQ+zyaKLCU
`protect END_PROTECTED
