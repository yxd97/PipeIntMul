`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KL0S5dpBe1WcvnLExFEh1Ry3qq+QtV3QZ59JRugmF6pE5aMOVuXcfFGAQmcYOJzj
eUOqjurr5XCZPXhViGLwzW9FyG0i7TppsZEJQ4B+p9MeoPekYV53oPTE3oE1yZ3b
F7bx/B7ldnams0kzBve8IEFR5HO4ksfVj3ONytErMP2YPyljIsZ+ZlhrTtaJ+FEn
G4pExG0fTjtefBJHzXF16Gwl70JNPgA+f+JppYd2TVu6eN/gATFCiOZvW/BVc5i0
NRvwQelTrQgcNIms5BC5WFpp9Y921o9KKg98yL4/u2jXdWFRmw+nzAT8YAZ6luIt
QBzjQN4M1e2/t9pT6Vj88PmQNF2KdemPwV9BxgBWDVZyjWKUTQxOT2N4eshu/9yf
lGquymsG87S03/3j3/W7c2N+EyHIwHB9VSV1b7uJkIQjFdcHv6TfmdeYllAkxK2y
jGxw9+001UK+D+ni3ywOsMaqWHo/Eu4b9ozpT40EkcMamIol5iLW4CgQezJpDuVP
KkV9wV+r4EeMRTh2VfK4fe+Lv5GkdecWK+Dd+GeI2bSK55sCFJ4DPm5ElmnaQ2lN
qUadrzpo52QTs7mwUHb7Vtl5Si0l+njpyy+2EglECmOqmXh3pQCW3NB24Jj21xVq
OroSvNr5Fu1EtiPQDmB1JyOZWDYBfToIhPYNpgNdQAPQ4+BJW9GZ9bm2tgRUOr6N
npY/tL7nMNyiR8cBs0zrfqxg5dWgKcd8ATECpEjn4YzfPZJmqxg53IwOTnTyLVe3
ht0QQfuTMSTBl13HeqjOfQ==
`protect END_PROTECTED
