`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0uUR4nP8IeVH3V2mfTVue95PwI0CbIZ+9BLpriOeF51szI3Ddj/6upW+5yG0prK
bBgvHHN1Twm1Oketcr8X9sMu+zsSS0JlTKROGU7dSaWenFOKT6daNPSn2JcRGeKv
D2mGQDffGXf8rFmLkIVoFoud9YuuInQqjShjeQfSNsMYXb1wvQupBQGNxzlQc3XM
L+ABvvkg54yjzJnI0Ct8/Zd8FssERUXNaYvjDNQz4mSN0fA0+fcTs64tjh1cVPa6
uYdWtYkKeOrWQL7BvxcXQw==
`protect END_PROTECTED
