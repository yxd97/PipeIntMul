`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fs49ywwNqF/50g4oxtf8Lkmog+9ivOIeL53CYcOH5OepyNlaThnvxEWOmkTp3m8p
NqzPgLp4LPhcU/2nfuKERLXE41rBloD+E4V+4ZMKsMciC1PLVLKdww5MnRg9JvKz
8SbFmQwQZqMKxfrcrxeeGFxKds46ffw3UyuY0vkWkhG6oyBLMHyvea03cp6qDsPH
CE/okpVc9cxcs0vUmqIBfn7GT6p8/rw21xcqP0jU1QDUf3IisAhHioWKWpR9sFvm
QBMm/NV1RZSyRT3KTqdOY4dYikgzZU3EkJWNfyksS33CUpqmscaXPXgg7qby0Bem
EjmatyBdf0m8rVcbmLiZOiwWy4AGYsVyp97jinTsPapZhpmBsHeyL7OgxioA98LL
jTcgNVmImQ87tkOl6fEDH9J4uSpWLrR5gg1MkpAPYsS5oAX7C7TR42Fuo6C3akF2
Glm9zeOHtt/6BcCQ1qt/MbYQCKHCEthZXwChs3R08Xrh27ddp1ohQaclJOi9ovuG
PSoVuev+LqNxO2/OHfdKrTw8FOR5pMbl49ghZTO2h0VG+CDMmsckBsYKmjoMKbDb
dPYpeJQ4g18HlhQZhmroK9KlkeDK2QtwNCQ8u0MjM2Hxa8THYdlS00bfhO5SZKbD
ks7eaa0QHYYZCUsc3K+vKlpVhyRLlCMBB8wdXqp4nx0=
`protect END_PROTECTED
