`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZD0aghEhSGFA2UDwCRmos8B4d8GPbRJ0czQnAztdiMhH2iG6qMBuPRCSH1FD0llb
nAcbG4/A+jQNwwiNYS7tB4EQLajY3xv+jpD2OAIaOT75tPIRGPhOcygmSmGoyIw5
FHGH3OVlE1tP4eII0in3YuxZkltgB0tcRYAEZSm0gfZKVDBi5NHUSOp6OwnoDSd6
X54R1VQMpExJShrcvlS+k3qEEjJzTd7U1AFUY0ZKyF7phT2nqXH94WYgZ4UNcGjI
q0/i4PuqGoTqoE+RFLJlSdPlr0uG6eDXoAkVNPt9QudxjAjHU4OOFMdSuoiOwjLr
Cxhd80LG6PZGIw0GwBAZdB2GrK9iNbSXgNd//F22vTjVZjFHuzR36PO4psawkAme
hozceRME6IeewoKnnKjhNfMCSlLWi8NJRwRKOVLr1K7rxhnzfMNj9aPw6Hf1smQg
8bvnk2L3K6Tb3nAQfCS7AFjflUYvSm+VMHmSE3oJAJXL6yvSDuyn8h7wMoZ7dkdL
77P+/6SXN2MQAcyrgXHIuqcr2LF1IJW45jLbtJpYgzSSEJI3BMrRzBWV1rzWstmQ
pwCxoqsiR/TR3a3twQhEfWReqBBS/wdTtsi8LdPxsOGcOH/KoJeUmUnRzIEodOlH
+UX+ggKogLstBzP0PDPz3I6YzLUR+ryKdedfYpmhfss=
`protect END_PROTECTED
