`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIAsya9rYXL3duUQx/XAMOi6fGKf9VJK7VJOLaVkBJVszbxy/e32ore4I4U4bVC3
28fHHb1RJ8/PXoMyQMAS1WOs0SieRkFExoAEbMfAbi6D+owBmKu67WGO31o/zyUl
T5b2l2s7IqQZBYx+ud/f6U3mktIb4/uqkddiQIoBSeAUSLh0ZPh//VRgifRff7GU
N3h3OeT7VpgvhxgNY1Y4mp04FpbmOrq4pyyMzHgltJvtJn/rW+zsVDdpPW3aHJUU
/K05KWheAJQwjobK/UHiwj46F1NjYBKJ/ApJZ0qXhs5oaXCNo1g8IdHy3E3RNWgY
Jyg1TBZejLei7VqvMFKxL92TDR56ahMQY/j/qSOsuVlrpBa7TE70UQBKT3fCLvIK
5fV1/eaP3HfCfGEEDgiLqQ==
`protect END_PROTECTED
