`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tgu8IXB5muAj/tX4twWoLn4FqVZm/6UJ0q6N+7pXVyPZgkdmj39JQz5ze8LPEX5I
g6397z5L57+HdQLKdNfQSnmH3pH5gqN4QwA+KUlBetjv92kRBHaeS9Z9AajI22J3
XPRzoU9Fc8pS1R9UY77yw+vSNiuZkRH40ouRjpw+1JrpifFdkaWbOWJ5Bgkhn8mB
R14MPAHfn5BDfrJGnfSpCjDZnKCPPJVWYa5jUzVD9TMUY4CpjPi31imbeaJ3g5RG
IfUD2Q1ZKZIE602JRpPFuH+yA5CnJ74tdr/HGmdjWtJH5rsE3Ws42sAzf5Uzd//y
hwRILp7FglC3k8Ii6+uuPiqNrGLa2AxStOFBqequWPD/y5NM5U2GsHz/w+dSQL3j
Z+ZfP2QzTNdA1g74VxhEkwdak4+2ZcFtJUYWFXssQkjgvix71bf1UXuVQgniDa2+
ZIey91tJhdUe1iz65qz9bZ483qZuLFqGb8lOOL35Tx66BQ6AZaZKdkV5S/WYkTsf
hynYroDdV/NTP/UwYoXK5dqqQWl+r2MxpUveSqlmwp9AGybya2E0oeBKTP19RRK9
AemTpZH3z2Lt6HMH25bfXA==
`protect END_PROTECTED
