`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DshHOhds6Tpx2ClUuSxZBjMVYYTNAOCMZee/Effu/0LLP1WHCL1o/ZhXb8BaGvNI
OSoyEqtt71GqHpWD9DbpQWckC3WPs+JTIDVY+h5O7PD+dV8FeckIo2UvowidRnua
ORSmDRECuKhuGQ5iMQznVZfM+qNtNeW8HL9jwVvS18PAswornKNMKi4p0S5vjxdL
iXA2875R9pBl1S2PQgDRDH394xzwqzKViT8KiU802VTRcHAFEm8YMfqUYSp3mcWR
qUgxHu+8x1upFp3AyqjR6MO49bZwQsNbbcjqLG8QiVny0k4HyoflUH48DBonCKYn
yPU9NPkfOkMk1cfbrZHcUhJAMM4guYKIYXs0bgpLMaD05nwKa9xCDv216EeCefI4
DzX8ZXVZvOJc6kga6I49Wg==
`protect END_PROTECTED
