`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKlg7lJE52e3Sheiio/9A4akAPe+JCm0Wv1shBU6ZX1zkEr5LkYASS0rPz0OAlfX
6w2Wk+oiYlpo1rJdct2qCX5jlTC6OEQatgaC2hO0qz40vj/h0IzifB9z/eOnIcUU
uWZ8bz9FoaIT8roLt4nHmtfxnQ/hKKbum7wHHTs3aAZQfEVs7BGXFAG715OHNsqb
V9wNNsFxY+m+pAqZgw9X7rkD0Bf3kDft5RuniqrrMqBsfAVnDd+CbJxBlNV0HYZF
BOD5SXH2xQDRGH/8QpKFxvlEOtsvth+QnQTjA+SuwS89IpcUUlw5UIHyaJL6p4uA
+xKuMeFloDY7dJXJHlo8/miqgeij2OaqKEq+0jm1vDqSrja3BWRHJkOw/WGYgfc+
ayC05N09gBLptRPkITjd3lfRtd+3ggHvj2pWNiuzApuSwn1CcKJFOoOhGVYEBsT5
pBB/jexQpHlxeZQxhtySFXd32GMP6ioyQwDpJwqk/2s=
`protect END_PROTECTED
