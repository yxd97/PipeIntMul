`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NBnW66CDNnpXvMXELIVtBdxUs2zNhFYmzqQ6mEjHfyzpLReo5CMT2TVXBX6MB1x+
Q2pbE3wKoGvmYttpsIHTeifk64tQhmhZKsP6wovaRPXQdMzWoWABhiVvAxQgrQuh
ghAr8XyIVD1/An9JnTz97EfukvVRuD79NsKMyrnW6zwUZRa80dJKJlQUcBQWShxm
Gt3WNauVzQlfijMf+4irIKbUGAc9Yq/kRcBDbVC/fAYCES4/TscGaC5xNUysxWFZ
9G3UYUKeRU3CJK8hY82bMp93o9fHocQoMyAcTbvBF5IMyqLcyBpK86qeJPkmmbCT
vhJtLu4W0yMIl/9ianB/y1TreiIBW7qJMvjDQTjSC1KzslYe4Dv4tDFDRtMVXxvj
FAuQCBcrCndeuJeo4QTf9ev2WoeqXCXSa6yXknNLRZl2qswiE60quvFCHlTwYixQ
tmJRr2wIoATnno8CUJWdgmVxwNyfsad0p6p4Vh0jrdLDYO0snn5VfEWvwDmpGOzQ
q0btqU39XYuUyhcDlAvbtBfWXf189WYdpYlfAj4/J2NTAo/n80o5yRpKdOIGKRvw
kZUrtbWRv0iRS+wcj+r8YWMVrKQWENkZa2nrFPCaSLxsdttS+HMQRE8divM1ExPt
a3Q3FTin/tJ3xDUqSHOyCsUDkxpSftO6txfLlQr+n3IioamXyRjUHMzm6n9BCLUJ
R1sJTpAyoOYl1AQhcR5K9voGOJTKuO6cyr+ofXt9sqOT6dkKabnX4Mcio0ZWuR7L
lAfMsiuFo0QCEm+w91rklO6abjicKgj8oxW1L+WE48OlnhTFuFXOWI2716tcXuB/
jdejQPlxwbV4UHyI6p0jZZoXbG7bR0M+8M0gxCX7Yo9wMtx1kBSbDBBw0Fkvk7Jg
kiPy0SSW6PAQUVfsvQsDGuymD7IwO120zicHCQmH5RrC1KnEVQsI84h1kW90D3r7
+X75EISSUZrXxd+L3uR+/lDKOK0RF0dUopC6bg0gAFZ/3KD3rGmkCVCOaeJvaL3z
t1pgeR1d3nQxctvCS477wdnLq8ZMP5mWmfZ39g3dFlhbJT3gu0+rNtn2O3ew3yzh
UXA/ArwqtMNiw/b8pVm98OJiNf2I1zh6Adp/MbZdhJNKAk7fuSEMms52TDMmh5Cx
jD7udDp0ua+c/P3eLlyIc567Jd6wTLclbQXMmMRtPXB8hXdmTdOCX0TOn/y+O5cv
AcUt96i0UJ7scsIE6NqkrV7jXTMltPEjP4MBFmmLdfSxhPDPBWmBvPzxBE6KcOd2
KWDdvY5WFMJl5IkQ7jtFI30egwfl6iOD8WVh1EZ4D5F/hc7jla+FQ5wUz/taZ+pk
BRPnX5Jz2wi+0Cq50dZ05+Hvk1zt/g79obmCCX0uw8/23hGqBvq6Z35odu7ydS2T
FBwtOLwrWJg+oKhQq5DrR9NVmCcLlZJ+J7Xu56hSkvJN5WH1rhdPruyiAC4TgU8E
L43aO2sPCsrZnAIkWt9jeUvh7SL8DmPtiG9cdHioYOn/WuqLoDXvla7HIbsM1gIg
lU2cq21p/Cm61kxon2rrdqgADMo4hzJG6FCs5RXcCEeAIiEYHG9f2Lo86r4dIl/Y
sX+zaQTdX2JAzpsMcV1B0B6fmxF7b78MQs93GVq3JkSoSA2UjRY40LhtlE0RfwtB
0XEsCRH0G8P7tRtUH4+4INTAgsEljsVinO8qJYugxNS/I1po8BLUaSXE/WbsBW/0
ONS1gMExRLXz/HirjEXhQsZj/B0fpY00WhNLaaaQB6YXyWbPD7ewyFD32m5KQP7k
ZRB6aZuI6UhgDtuSdL8HPI4aOrFnTstbEcyJQIM3oHvSRf9J/hLGueqB+jYqUC0t
dQtVAx3qocRtvO5JERZ7HtzxKUKXOaLZ+PXX9NwHqMnsoxJ8kVPUtGibECr6IUtk
3gzv+2ENN6XLMsQZOqMxfrak+f5lq2BqvF73x8wagJrQ19Rn+GQyMuDvnqkBFVVh
IH/OV+cHHEBSvPe1EKGZkGvqz9hoobmN7o6bsKuynhSdAPSA3/+syjsTsvLw5Txw
y6u1VECv+lKu4G9vOgjmEyzO7b4/rgRs6WaHhZxKKSQGLZkLzWoO1KI0qIHlDiY7
KcFRUYEyC4MioemEbo/MSNwB/vftTlkmcqbcN8IZmdsm1JavcPGx57W2mxBkl8uH
ZfKYcU7MUz2QlcUAQFSxmqjhlaZ+0lIjOZJPvNdYlB4Msft5kXe9tSa485QQvMMK
aUumdzJu7IJU8ZNR3OzpmsDdWDU8gS/Zo36+MZvXzkYR5f7+Cl2BxNQ6avmaPug9
mMf6ajDWGj+Y+yDQMGuUbWxRYZvEvoq/eEsns1L/ZgWs5AYeuFfdbOh6BWd6fY/4
IQAA7LCmzOBS1TJ18YZ6lQ42pq1T4mPyX2g0TK5mIuj7Q2dOpwPDcphexE/oNVLq
JXbrg3ArzBeywFM/bHfcsRu1ersIhsCpNUgBhGTvicKob6C3bsUn4TEknvbE8EI4
CXCB/ECT1w1iL+a30igFc/lpqAsrDJWamvZc3cPel0/Qn+bH5JTBre8r1ixYFHqN
4xiBy1+Pn2wQ5pb2JQ4c1qbXDxOhmpgCeF8dN3o4H5CAnYx9h4cWy6SDpPKganJ0
BaVfpzvIW3Nk2akwwZFSxQ+bDrxBfDqoqpOMTorXmcgynRm6MWD35T9A/IjAM5St
Qlz0IQVr3Q24TkCNXpzVxjc9U+BYY5Kc/V62vYw94vg=
`protect END_PROTECTED
