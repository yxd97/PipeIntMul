`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4KgtxBG0vyTDhu6DzjfVGTrSD0Z6kraJnJJzjzecLsyxwDA75Ppg6w9Zs77nBEX
vYEej5y5CHjykRC+gi3GYCSSU7EsKcat7TVG3732M5/EjfhINCFGTdpnwGSUUPUG
KAk/BzUKDMPqomx8/ANL2gZrBcJb9VtvQ9MqoX2KkY73WvdySa8LttNTwswGMuOT
HCcyTGzwIJUpmrDT9GmlWluLo16fU0DxvcwZSdpA3a1AnEG9t335umrgPWy2yzN0
+xYopKsravTIDf6aOU+Uz8XKghu5QA7NOKX03XVr7sMs3alC8b4f+DT9maMo7/5K
MJ6p/hGhRn2caNRqNHAjyXgZ1wVeIl5CsiSfK9AKrbug+JFylXCZiB+1ItiEbqTq
r5MWKqcu0lbOJpAVOZllKg==
`protect END_PROTECTED
