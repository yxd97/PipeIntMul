`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0xiLpxIv+Q3nCeOg0o5/tE/yFefW95I1fzpOFRobmYEtMkuIxUpwKXvB5Izy32/
x92HfE0aXm55HRqXob5bSIDp9CHPLEqvaQNcFwWGHkpcZooIaE/r/XjDs1wdsAAs
W9+2j5zMdJ1MYCo7QunpII9aYJJGvv5PmpBHM18GXD56cTjq3vzzHv1TtAqw493Y
/B778SwlbbnSjZaWGUKyuWxHLt209Wj2rK4TJ0Ea8QBslJ3uTUaeOFAbi7Mv+ORq
CxWf36Z0w4OtF91RvPqYQtaAOZHXMlVKPzQMYIioMeKl1Lh60grYQuRezPzK5zri
LMFTgJFvEP3ZJXHDC1BGLy846Fc9AQcVoTdQpevnxQHbwho1hpJrnZM2H1GPoNdC
+dFmioLMd2+O4dLuilfy3A==
`protect END_PROTECTED
