`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5LKJFD2+CT09ojyJOU1haAFqg3amwSpI69127Berf8JUL2P2lxJ3/klsodZzxBMH
jnOqc5HpEAtLk7icBwuGnimch2zdtapyrGWEQ4J/xcH6GM6Juv8LsTGB0k7KCfi8
5qu7CxEIRRXExYfRIK/nF4xvagDzHVgA02N0FcFXuZHPkGIKQUXlCerGuN1l1SFK
x8cXkpmxOVMl1OceVVokwiI5D4dSVvRezx3J5HZBeVG8g0zxq9W55A1XiP2hOe3r
8ZJaAWHKFZJ2tDHle687vMdosANJQYCSTSnaUcSYICp8r4UYpo2Ibdkik7B+jQx3
okQ58Bemlzl+4b6aFB0U7MWPTNe2xyr3IGAfc+y891ePeue/2uP9wIM0NWpA0wDG
pZn5vmC9nlPRNglvnOwsWCmEpaPCkJX9QenFm4w+hN22guTZrc4jkCUsDhYbi2ld
`protect END_PROTECTED
