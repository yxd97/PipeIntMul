`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c16LRnWsa4CCvjOUlmSzE4BkoiDXOrvBXER3kuLIqRAXtl0zLb36pOjW3UlZS+ea
MZVqA2R+fIehkerM0CLi3XJpOYJDybiY+icSiNpv/oEFkIuw90FgUxjbZCsTlYdI
PKQYYqjZEfBW3y8cq1sbjgXrwm93+FKXtbqe9CIdd0yLEsQyZN97AKFIqXOEzXjF
QvAyLsiXjHE9pDCUsLKLJ0dEYf4s+iqX7+BXKbaV/Leb30oSMnAVvceCjkNB0YaA
c4IjcSNW4tKjPXQpAsKGY3+gLVqJHkoRCm2BrftjcpANwofn6QLM+2LwGWU/jQlL
noA4hufz7jhXy6qh4CHIWRyFifJBkFfTYnJpg6uB5uXsR7g8JcAeVYb7IU4zHrK1
HIHiz9e2w6CuNy22xQoojCjVmTV5A74pIoJb/wR4P9aiH0SrX5qpaN4TKUMkEB0N
`protect END_PROTECTED
