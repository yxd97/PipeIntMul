`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E52vtYZt68srQ/rrl5zXVg05+PKik9aY9j5p2xbVwFoO2GrNdccdEoAHW3ZvxjQ+
3J5kfTritbjvwA33CEK0DvyPy0Y3GqwFGdAS2LHQSXWUDbf2nditidAiiatdvwjk
fWdTefSyAaCMD3/FRxQcIsxtBw9O9tWnuC7V6ZHugBvGTgSujoA/BQ35uZ6wmZmc
qjMWtNTUIYPud3mgQqzEWaPkcCCGIrNxQWQCFH+v8cjfofEcmb/BOXSib4fZchmP
b9i0g9rG4iKAM6YpKcnq309DAf87cKcWbjF/8DjwGQQwBu14cRvnxa5/qino71DA
FFq58YSION3xWyt1vwHpL3DG0qDJOB/cMjwy91oBj1aJpP3HgjPJSXjDoOgJFvdt
sAhlTdu2HS0tmjt7j84KU5Vogr+e5xyL97PoEOr+MD2+q2IiNVCoacGIMP14b1Br
`protect END_PROTECTED
