`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+XDbzCFj8u3rfsKeMQFYy/yQLM8Zyf3a9+P90hC7BU0xE0KA07vIWW/MVO5/oJ1
Ij8vrxx3sfqk9s+mJ7wycg27j4OJjSb4RppzvaWgq5Ku5fh5ydue8XbTj3jBmYJw
Ni9bb5jMVKaTUZZpHg+e/4DPhFMywGoSkrYKUmesGLwU5j0X4cuw5GvKxvGIzHD0
xRalDsIcZr/P7SmC1+21GO64RO1XR6yyScAFbmxJwem2F/EDHqPWol8Lb1LKl1Ff
DUkK/o4t6FTGRqt+Lh26Xj8PvRMuuzXNUJ/Owhw7HhI=
`protect END_PROTECTED
