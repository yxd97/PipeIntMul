`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkAk9VVhcaACSrIeKYxzvUUvzSY2zVNIWFN3BA8dY2JSxFt3tpy9xNgRz9nuHR3s
UrVlexMIRYtUDgAwPmjnFI/1ebye1nuY9BHto/NqusvTVGtPyCXWZf1T9xqlNlwe
p0Jv8Cksfp8eWx6um16Z/7wx4oTj1vkbxIZPRum7GhkKBbepYqkm/iWmcUM9opAY
Dnr6Pi8yVNa7QADfVluSXi+JW0ZL/rrkPg8aq6qy1ZUpjLr3sB41EoegDVVjH5a4
HYQvCHo3VyO/nfOTJ7/ThtQiRzstdq79YJygFGPhhfjkFxeHpUlKQ2OKuHH7i9hK
e30l4QxPfJy6ZkVvZEyKoQtBMP7YGx6LfI5k8wd78UbEsX5wKUFEQ74RXEOnEL6r
F6NtbFlsL1+JZs+xSvgHrJLN8d3qJHJcefpHNFtyeCpRPCHUR49PXuGaqMvyjA2H
ye3Q1L8Pw5Cnb+seg4/m72eYOR6LcCi+MyHDAaslLaf08TZ0e4HDapb3rQQaXL2h
Oocnil3Tfjckb/CwrogbnaNRTo+aEgEiplLerOwaWpxN7Pc4ZJzb6khGmrFDmmWZ
NsENfjbTcnMfOZGxfMGp/0Uy2JLhKILvY016/kHcACXA1V0kCciX/ABhzbKbwX9a
o/4JkuNGi3UftA0Ui61FWzzGmjR1TyeFi9BjmRjl82Yg+mVEUiqfczqkjsHrJD8w
wlFZZvza0GPld1+JQCcOueur9ZpVben3+zo5FEgsAlGk4LCr/CRv7MYaUH9UiaVU
Y4AdAcOcNr4gUsdUlrwZ0YSHgsp9Vib9TcuAUPuKpJ2fmGe4ESfI2sO2C09LP6zo
d4Iyaxb0y1/zshVbgbxW0+eJTMJa/kX/uhB/pgUeMrf8n68J9dXHQOOqMplAQ+BI
R5l7CcjwvqQoC1Onc4UqP3OPXeTUyMTvwFsDj+Vb4yWAY2cEKrEAVQQtmvJ5x6Yb
q5BYrBPENQq+jJGY21nmqrnzkN8ckOrFQR0UtyL+INAxXctTjaL9EsLUjGTn8Uou
h/B0Igir3dZ+k+C0+UtdMTW9x+G0RPd1wRMsmdtX8MXnqgSfP2X1rPPMMvBge3YQ
8RPRRomOqb74EfayGflxY+OgUuh9d69q7t9ODRXHrln4y02XlUaMLqD3DFFuEvKV
ZqaFlmYvD30peHfDS7UJDpGYOklKgxcdMUJQJhEmRdqiKna2vj5lDpmyHveykNYI
bbiXlnVnoFLHB6LejgTY5zdmBLvrWol9545WpH/7swYlSYD5C0BLlMMuYB0O93ud
`protect END_PROTECTED
