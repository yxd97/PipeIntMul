`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpNcJT73ARQWLYMfjddEb1vD0fMk/F5E4cFcra1ywbYN4PKZUlub9GuBoYiTyuMw
c1Orf4phzeUsnHDiAVERlFbtvt7ipvuyAqNMqFPmbzUi0k4JIU6H/TLc9L4l6nb/
/Hxpk8+xh/jeyKp48ShWwOb5ciPgpfZ2iYr0fUn1JKBIgacgnPKogsGPn+pOx5qX
yBQOMFcr0RJa4avm4KYuxpZP26L2HiLoYEz4SkeQrVcytocI/N2jcQoWocPEofXt
JgFnQZHwy7FXp3XiI2cbyGhkVq8uom3nv78NAIm/pZFfkenzoBXdhbTeusVpYxrH
AM3LhEZbhuM4Yd0CTJl9bgbBivyXyvMl7msxT1e46MZYpagj/G5sfTj6sUzXu2uz
rtWNQOs2FE9uYCYmF7wMpTSxi7aBhhRrY00ExKLRuURhB1Sy3cuQ1KmiX6xN2rnt
jb/IlG5LCx2Xh0bHxkZKIpWOcpNv+UNNaUt/CQTqew9NvrC3dtCzFgPP6/1y8qWc
yqflaV2tHpaiKnHFxQfF/M3LPXwZqleRqIOOpZBmDdF3dlpWkrDODWvmlTGXivw0
e6pfB3Creoc/6l57O0iNHQ98HIEMUmOeXqym0UQim0msdCudlpabUaVgf8mMSMp9
iVkKKmxlR9S/B/5dre+/t11EaVW0xs0L8UdJWBE8wDNdVG9htCyPYmhB9hoS5AI5
mzmpxXJUqfuleBlhhrkBzIJVRGqFBbR6ZpEX/tr8T22Eg2Lgj8QeTkqW8lmArFZ9
MeilpdXvOouz5he84UTbCjMbZwlYTil9vWIwZA43hnMUhGpKRX7v3MmOaKmJrNqj
BVigxOxrE/FadWfg5ccbi0ZXscEKrCgfkP/oxWMzADdxIxwJ8fvTPbfcaLaZKiJw
Zr+8d4DoOEk5WMuy8kLKWTqIkt03EAntBKpxdiiw6OawCvEJXplcT0FEX401Ohvb
e7uoGs1nJCIdWijsmF8y1CVH9hWvX/tmZ0ZzO0XjpKgG0+5ihypScKOj9G5V0wZ0
lfu7a18gtco3ExOy+KT7ImfXmd+CUDaA8VjmKtzM7uGImm1AmczErYvBf0wHMtoq
1NIkIihQFO5AxP3TG1i5Jo0sPtaUMJMbiZEB5kH6G2iGYpleAa09H9JibzvZySu/
V6I6ld85SYTQFwE90/pcGFarf4Zj1Jr+2R6hpP9jkWUM/5UST774Cg4KcybYP5PE
ECUkVSOCL+8tZ8VAXVNLTSJdJ5A4GyvRwt/JGPEvCj6iJGzvBBUXKSpUF3qcPgLc
`protect END_PROTECTED
