`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYTDKAnyWj2DhIGp0Rj/KAgkR2QNMSUqlEromvz00n16ogyedbEGTPXUuD4IrvCa
DL5exli1COFLH23ySO92vVdwKyXIfYrnyDSY6P5t4z4S00+IABLFypZLLX/X/vJR
rYSW60HqUQkCj+MSnVUiF0TjCembZWl7bl0OnL11z/m202k1QVmv1x6i/q9WQxQh
oMT+O7NdhPvTJ5bd8Ok9NEWS9bQUiIL48B1DvnccT1O/PwJMLFG+t3cFNpzr03Q4
3m6XSSvVRBHf1JrYLINoiTO1LnYtp8WZUb9V1wePdsN9SPeAq/c5VZWvZJ1jILBe
MacqAFx4wz1PCmysV6O/tX8Qj52v4hW5eM3pggxKeLw=
`protect END_PROTECTED
