`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6psh+q4Oh5gdNDRxQTygG+GlvxW4krw1zzB6aSjD1RN4OodNXEtwBbNlFlrLlHgX
0RuYVPYKIRKTIVLC6A/l1sdF1OG0LPRxMsPh/oZiiHN88yddIw6FX1xLnjvItuBB
0Kz9CaLPPm8C5cAFb3UUGvon0N/sGWfJQN2uK0ZZjcCgSL+xIkPbtY3PaeddBexd
AhPNQ0CxwX+ivNNtnwBA3jDi5FvG/3FoqjH+4Y542Or4D6RamS61sPOFhiwxBr3o
Z5z2FmbuimogSVrM2WyQy6EdbAlLm1MM04Z7kD/Jow8/cc+DU6rXdcUCOz0xBL+f
GEaKxboxB9ygp1Ef6NUxaokjr79YIXZY6Kn2SoN4NSdW269BUdP5WIjSiDmNTRBh
VaQ1EOI+qatF7hnzGMid/cuflNuv8798Eu7GFrqMD8kQO+QWLYGbqk++oxjDinnm
7RIPYAIgkHWwdDQ7m0UoVg==
`protect END_PROTECTED
