`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8VY+ganGSZcQa5E6Yx/Def2CemD+8uaDYRxldqXve3WQ7Q1m7YQTGAS76KEU6La6
2fJLHmqgAxPgSNdO15JcJYlEbO0evVcdhp6VoKbbdWYQR/6yLoLhQiw1Bfk8UEQA
S25zQ5dw0E+nRPSzcxbC+vCFqB5yBp3ayCV3+gsec0TMr2Kx+BizPj8sfNLpiIjk
g0xvBD2GnTi5C2Bj0CHqJtNDMEMqL+hBHjhTKoOk3rDcszcIgaCg2YrOxYvhwe2W
/wBON5sFhmOmN9PkHIDbQuEBCnQypx1sGjaAzEN1soJDpm0ZffNo4g8ekU6LrYeC
tmR5OIDBZhDYF+gLQDEYYDIF0NR3hXT14lyIrsQRjxMtgChpSXeDBlEvaEqAeeUw
tepO7wahND2+iK+mZnIJ4todfrEgfsj75WMBmiPotaI=
`protect END_PROTECTED
