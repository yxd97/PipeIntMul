`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NiI16IhGHiawuM4g5IFBb1zpJdMk1UELbpxJqhI+jaQ0fUYiaV3jYDnEhxfOIxiA
IGhM2eb05Moce7/fenFqh50bTUAXgxoEDg4xH1SzNu/jbPtHn5sDuPQV/Kv8UnO7
fKciF5R/9pgIYssAoCq6p/kye2Xvuu1cimTW9CZX0jJFz5lnSPNWAB8L+RXGaic7
O7EM5YteG35jFDsC84Z0hXcUGu1rEZz5ivoUDVDYwnm5gmXRW+OTi+J1rR7vvQ8g
hXsSfTPJj2vdejbu28vZq6l9uYmdjztByx1rYLyAyROXAvrE9BlSPLZgjRvh+kOQ
XsIdJD+wXnfGMKLNIQWXnIr4uV3NIkumjNDJ4pSM3hHDbN++m0k7JLxi+HhApnBn
XrHatFLbWUPyoDLWaxERR6bMQQUCdwHcOS9fM3nIp/bI1hGEdARKCgaL5RkGmpTK
UBJ9zrB3UJ+Rka8jKQ62NdC6P+P+bnPSzgAVX2PtHVcfYVSYbSFJUQYJNak/RKU3
`protect END_PROTECTED
