`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v2Kdut5q9AhV/IsMpsQv9qvLks4XEOiAxXWgi0d34wBZBOdYQA6o7Fe78J3M44hP
nB0i5X3ySCoTsdVkTW0nFwwpJ8/FkVg9vI0ZyAKTaPpA0/QjTywJqg+8Vrz/SPpY
GhKSxboqdLG+lq67g2T4YGY3w3+XwZZ0PmLz1AQ0XSqgkoefWzUn9PTCpIvFpZwr
U3bRJULyCRd5sDjnIrZ57KqjmopRVzy8OAh8nv3KgmV2qVIUmqYUvdR6vOW/hSZH
mDCxtdYQU5OTyY8p40hN6qJjoxWASD82cJtx3DU9JhEgXL+HAXKRSd93onfruWqW
jpN+jhUClBQhSO7Er5GYBu3VlUxV/MTDkR7NjWIf4grzzLYleagZOkQOsVNZDxwz
LQGMrdOvN9OKU23y8lZ24IAI3dXb+MyVsQkYhzEDdzE95hgzW0GpubV35cWuqq6A
mVu2yx+K+zW2HERhm2+rfv8tyX+s226LV/GjlqORYjo=
`protect END_PROTECTED
