`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GDLNTbnStPJJ+KIDrjIKt4hgZrw9Etac6BhyRFq2GhELfuTfXdU3UmL6/7iX5be
BqdPhQ1c8Q7NdbZEoMD0nB0y++bWHDNJfqWYUVRwS2umncMUXejfruai5aONETh6
j/VJT6X5X4T5taPXsKT6/VoPZoGQHtm4LYLqqp289ZnR07Jhze63kzKI9apwMuVi
DddDrVDGfsGz9rGFDC32CW2rIhpAvWuy1AlP2c/Oih0HcJZhishrpeKnHBCnXgUP
KqQfs/E5mxBc1JhrZZKSWLm/eydInZ5wT9ECMB2Ofimt/FeNVeA8Whz5jAlZqIem
p8RGEInOjxshnna0YflIio0XuuSSVIwItM1GRdc+4BOalNorcbS949ee0kkSyn/C
RE5hbKLCCDVlTTA3X8v7xPk7AyeNVL/cNxYz7tj/9yrrcLU0MXbOhh1jkm1UsdpM
cq0MHFC1Wq+KKKZy/W6Xu5xClq8AtqWqLskVkcIrZ1+ayDwVeZfFXM6a7qER/y07
`protect END_PROTECTED
