`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xujomy1lhU9EzPNJJPx+QlwUN+ldCI7zOMdjivhQnv4sI6z1EgzfAbVzQ8rIIflO
6kuIQU2nKVDkF0NG2ctZ2Ry27bQNQ+SDVu3Ck5pviqJNwe6fFWDCBo38tVEP1z9Z
Howx0DlDM6so0Nvm7QYpKWgFOmW0/yVcBo8Db5HVBYvY2lGInqJv/qwg/TabMPoB
l45nUe6npYejYvKhveRgpyUJFHqyaQJxQ0+JSHdrsXbx1oLimHApdC5hGliZWXLN
nRuD1aO3OV9YugOOOyzC6PbqoXZcH4irfabB3l4hvZeN4pEpUnpv7kt0lO7sHd7Y
2MsgbGIZVqu1ntLk3zNHQw==
`protect END_PROTECTED
