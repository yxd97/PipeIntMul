`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzhE8PvaIKbCYqtusCrSdA9s4G8I930j50Fxw0Yzj0Snr0SnENL5NbAsCoaifZBq
MN0kGrRtsl5CpKWoOOy23a9V041U0+3RRqAREhl4Ke93XZeO0N2wSqvA+NC4bud8
m96nKzBiLGzxeBgoU3k7ZhAY6gc1++T7SjeOYZq0JayhbHQIcRHaJ3zMyBPlbSak
nho2Q/cuDoJY5sZCK4hys0rPNJHoE3dcO24iXYyT/E3x2adCfBRK+8hrf9BPEyyv
E9YO33VbV9FxgK60/+WRNVF4qr610FPPwgPEfWxRfNxgVRagirxQMYJEHSr9p3U9
403NJ63S3zkLsTnAJsd0S9Yhv6ZUINxnCT2HGdpEjROAYFgijivi+zQhA4KecL+g
uBYoDv5ZqTclL7WJv3SwWJdPrLZLb37yYv0b5UuhH+aV2XBvgdFJPXoXhTbaiFES
OtBCsZJd7jCtmlcM0WugCYin67RwNxeOCaPwQvNdNhRaTE7DtqilO6tPsdsGd5qg
RZ1iUaFEOI4Ky0ia/FzO431+VpCuhwtBZQwmkfvOgREy/Hj01kJuIV4uPViPGU+6
4MHF2gf6YYs5Xmt9mkEmzKKUva7d9s3VNjf9E8sZwtsDM7g6GQer2wXYMpU4sHMU
Eszq/MpgEdmgkLH8954JaPvtCs32DIkLq4GovCXK9i2sEOze7XKEUSNRfWVrpSjN
jEbM20EbpBsdAwbBZ8hMBY38+v/ezCPTJR3E1WkyBmxFvA4aWBUJYITkuxQA/MRH
NOZNnLBHoNGAg00Ip+Ab4pqoTDBevj2jVCt0anlN85Q4SQjheDObP/rq5f3LXE3s
7epqlghClc+gCflXeaUe6fPjAYRusU7QFQaaADcK4g1g5VhTN9UP5YGqbNZR+PdI
zqE4K+jSNGEQ+boqheN5/i6CxHMKP0Dn3+uEhvtOmJlD6Q+NQxctVFOi1XzdwZN9
dqiscCERpZWOiuJlyq4RUgD+wszEEmJZdOl6YryMprTiXQzlyaFTJEFgFZths9a5
XABvxeHW8qDcmWYd2z4mtidMLI/cpXZlyusSVklhY8/V3e8xHW8UJzbJ7hSdmiMC
8xejo1iwui5TvtNzGg8vgzSH4ZUCipJCPCH2oLqdePro56BTuh2AuJdKxCbHsqdS
9hjyWzr54ciHVXuRBwqNjaUbdCfLsmBSqGzTCVAiMMuXrSmi5GVG3AYAqAejeMWx
MLXZ8lAaegcYoID4QBUtU4RAwlVrICKBEjqMcZAR8Fh2hmWSm7qIbFCsA2jnPix4
IIldvRf1XBYdH2u3VukALGJ4k20cNEuqowgCgYkevYCdlA3h7eiHM11Wj/dJC8T3
hmsFzC/ibzZKdu1aIniEsT/pCDfS5i9G3xq5ATxpJVb4eQzx49uRmbsSYQUMp7eP
RM9IsQLyaHAIbklUv4uz1HCNUQIt2GHjHcbKpOlo2YRQTpfgxQ8XQqP4hVE0qvTY
myAdnq2f/XxyuknF2C2hfLncX3JGcf6AjvSggJJU5+oA2hgErZZUSu4rfgbach6F
yGAkxl1xnqmtBYnxnVIR0DaQM52slj74wVMDPBGDudW/HJ8Nol+d/0eXGPRKPcCp
M5UWo6J0OR83IPFYBFj/MOWj2TUB6bn66nV8CTMRSrDqIQ7DCeJgGVPyFJhBiV1y
WwODss2SeDASQcS7xFthUielZGejzfcN31PURay0lcEwF4/n95CDwwLGleVlqIJV
C8wWqlcZpMLKQNtk75lQQSuEHFUuPE87cGY+vMNyTt1CqhVIkcAllqV+/sMPL+br
9mLFTqLYuweCWfLNF5AAWgyetx7IsiOnXK5vV79/i4J7ujobghovsFhBq8HOWsWX
fDzAuX0dxTpBeN8Uc+ENkboSRCUTnVRubAaokN+6TgYSYPFxdUgdSjLelqQsP2Dn
3RoCA5K+kP9VETA2m1RzjEtEdHYFSz/zn+UVabFJoNMWTRdO6pVTtp8tKudjr7ls
IX7nBaVdxgpa6vf/s5zRre22/ZDpwE7rg+6X6vaYd/8QeQslFV5MC57h7jm0vUj9
74QYxf6VU8Bx6JOX3hD0q5i7U292dl66Cm7HDbikCAXOHQIpojkZKrhpH2NQfoId
kdlhOw+XGICzHyJcWwtkgboSDcbCFZxtpGS8ICgJLQE405E6Xq2poe1J4qGrYS6j
fgeUOx2VK6O1NH8BHu3Xb1SE9pvsYtgP933Eh9igbnxfwt7dwCtxzusyMPX1GYVb
eYwTOusyWSSlngtABK9uqdYJp3gnsMx3qsWGF6Rwa4qd06cS8Gkcz00BF0QPz98H
c8HxCiLx/llOgdZiWfLiagVerqmL+lNd9sVzYyvdJi7+XL0hceatkBxvN6U2jKwz
DuQOiaqFUd5DjkNmcWyqzKX4/+i8viy7jxQoz5teRg0xwLqqH/glXg/iZYezIv5x
2hN8b4CmMwvQAs7Lx6HY22TVZGOQBmVKkcBGxI+VN1sZd6CnOYpsl8nmLXO/QQB7
gAVYvo6SMY+5P1Pje/7OHhBPIhjHrvZa9TCY+OtEkND6K9gR7e00g9UVZLsy6b9m
tDWRi7jrlUnUM08ohp86ctlvTZXcJ9CK68Lm2Kk6QQ3AjrLjYZo9TzuaGtrFK0gx
Qirt06EknmtczLbLoYl6B85jOyiYMNeYHrjMSJe81h51SGSUOQe0Knh9O+WweFKP
UhoiaY4KsamCYIM3G9bCqkEtG5RJkYQ5v683v8nc2m8YZOMJnJvjxhe82u7ww7AL
mOuS3jMHN6kDysbm4yMSn6KySAs4MbzenmEg9LugHQS6TXAkDIZbwUQrsFUOMrHB
Z88llEBo+co97hzyRcwaVFNIo39c6o6I5wT02gtbwWowYBdp1lrFoqGguIHKwG8e
fLv4iRg4QIPIQWYbTNTs4ulv7q5jyA/hU8rwzwPZ5xeLVjKOrlKnraRAGjyW/KL8
oj1J3iNYDBT//WqOvt+Ek2d4g5k/VocFS7t4+mUDILVm0vfKLHmP5kVu7iFQqKCb
`protect END_PROTECTED
