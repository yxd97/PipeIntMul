`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6X2pyeeaxwhmqPtTSmfjmf1boFabilH5T4FaJMD7UN1GIwAb5pJ2w19V4s1Zo6E
fhESqDRlraAy6T7NkRyeuc7XMaVKJgN1QRCAT+E9IQfg3IJvZTfBLWueg6Hj2Ho4
CC3G6s8EUdIXnGAVV7Y7oVf8fHct+Mu+8F4jeGATSuPPTaFsTG+o+uAsBTWJVXf6
jShgCQGS5TY+hr3JnI8MYhW4Kc9q8UrB8vgt2s2Cl2+a4RUsfN08p3SvXXpCZ9Qh
e/pL+nhugw217wHp1VSwqu71tkK2zRejuzaagKPavKMmBSUktvep9TTItNqdXwsU
QA30L1DSfUlfoQ02CZUIfaaB18JoxTsZfOuk1VZ2WnQtZWbkZ4toO8tDeRpUg1AL
5I+hsnpbgkEXtfWH/hKVCp/PMK2fStjH9I0WjC8sIGFiggbM66HUcp3/QZXpZHlO
/fuHpEVyjD3bzH4D1BcGv688GEiLV6/9Xs5EisuOxNaU1t0EB+hEBeqnsz5QQtqh
AO6vNxGkW/0ezesPOZVtcIA7/8IhLiBkb5f5IXhvhFPhhGerd6/c4pIqBFzJSXij
g8i+XKCCqGoJkWgrHLr5tJD2ugfFSHWVEZFY4agFno0=
`protect END_PROTECTED
