`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/xFErkmHjSA7dI2AbVjEBXcEr/4qFWXsw7ikEMYmLJdktijYBpZvSMZwC62WfsK
lBRAkjY6oeqvz6T1zJxeTh6YiWjY5tctrlAEgbfW036sqNssinLDzBzHalIZSIgo
l0ggCVQEChxV6n1fvyscJoaWHXeXgIOh2k6LjvugqAHQOFw9Kx1Q5ffV6Nk+svc/
2e2QZs+FdR8GDkfRupcSLV00hl0w5Utk2LEsQbJxe92uJjx4F/SjeMFEYGhpmJfA
sjGmLTWd/Geb1TUY9tX6wIRT2VE2BPXxRKG8m75YVFlYKmCKKy+sfhpvGu1WbzqU
TUNSZQbKbtTPXmLa6uiLVHWQg8Q8B5a+Z+Tpe/WT7dhJZVJabSPYUAfLlIQyiTWY
Ix1sL/wfAcK/zvHBEfD354YwU7Thdd7qrOR1y65/CJLpui0AUdHI07+ZAJoP4lfV
Z8XosbuD7W29dmuM/hD5kLKyYVaPMg0T48DSjV6OIFQ7OsYBTYrq1deP/4dDOPlr
PHoBCvrh8qcWbofmvh5X2PFI9EaJglIc2zAwzcMq6TDdLgtiiHmxUEHXQi8YLDow
llG9DN2mPF/UPBsUUaqvVpbSjnEh2cVCjg263GWoX8FzAZ6Zo3koQt/+UVjZd17K
P/0LFylUcBBZMlueOTYzmiyz18lj50QAopfM0v1shAHI9dtYVswJVhtp9Ue7+Z8Q
czCCr1iUP/D4Byuyb2pa0mnnE5ZHfgj+svDuyDSmDRXimtgyf6ruYN1WtAjkhMMf
TdM/bkJWWVV8Ka84dNXbFRPcC/IxQG0+D9kCwAXEpORiIq79z9ryMkLWhBIWTATZ
V8l1ZRhqOSxEOW9IXAKd+WJAO13Eomhks6C6vpS8bdOir2jqSx+Yq/vroaQZBeyQ
oiNj/rxJDcSB/B8/WG3tfMd63zdDlST7jgR3D6WdJ6ddMcrlDjJyr1pOTEH3QBYy
qH5lo1AkntfXCmQIhWu1dFu5RKxu2+xpuiufDugZaSL87vOC/D1aiwdOtgYJafen
4uGSQBwmbqziKgRxjaJjlANYag6KJitKUL7g0ttCuHFuUnrpBT9WKoAQTGSkYJQp
ZdLPIQZOR8TseAy2k/rGrYWeRl7TAqPL2UIxb8MDnPtBN/iqP93/yQamhITrNVkp
BKjXg2k737cD05s1Zf8wq71V0H0i1Adqo65w4PZ6pl/f8uA5H1cKINzymcY2bcNh
CEjbxgCkyvxtCu2Bwt51tkMMvMUK3nElldeSXw7MVLmTgkdss8N6nxR5bA3Q9Mb7
yVeS8f0QlWFUK63dljyXGaxc9dgeVsgs2Uh3UDO46uzE0zoeeJZnVnjeCyLiLuGg
slKAB9XcO784LGzb5FGooXcXiJpf3sD8AjdMSGT8nrPlLyCC29J6obdgDHj6Tbyq
aXf3OXl2ydyC0MvFntxexDtddWNfsjRlz2TFXNKHrwPLssdTqGh2ZERCDt6P0Dhr
FRXDQvIRqOVcTYGBbTIkdfmeqN+9GvBKo31FE3xtbKZNQnNcaZvHpVJmtMXSRAME
K2SQgi3mdxGK6fsbaJbpfSfn+4jJNtMYOyvj3ZRYytg4bu8gK6tpZ/muB3jnV7a5
hbx0zOCVr3jliIBSovNS3oyUqmPxejROdgkUbLm5sKG/iJNpgYkqEX6bHlWPafk5
MjdtUiY+uGNSyaP+xY4nSE0S5Q50XU1ni1VEFU6k70SYcX39wHo02NAZavAZO2mf
q5vgp9XCluD+Q0FbfwKwQUyhvPu1j3MP+4wrX4n0cXSBdzeegPv8i6fGgT8juFVG
WfYlTwY71suIbHnyAXN10Uv0GBSxBLVxDSXcY/W8Iqa9TyMj4RM21tN8ZVfwoonV
2V1LCJsX0r2xpIT9hy4PRq3w7o/uOeD0CPVxEC+m1ZOIAzhb52bAOFB8dP/dlPbM
QTl/jREhqNzkV864Mkiaw0MLb4nEjyRVfOqyGu5QXmgUzgQNFlsuYQwitDE0Gw4X
tcPlBBP7WWo+OSC9vRXshhHh1bqxPyz7BHW4n3RiT5E56jTBs1tOjo9zzA1uBKNa
XoZTSjjVnwC+1sPFLb/44ERCRRvOzu06/Sq7T1I6oMIedk6yV6RwiuU6WeWLQZKh
FhI1fTAJ3Ch8RTRataqleeiMImmZ8wIN9JRw0eUmJRqvwJq69P0zatKurHKY2YAk
Gkr8jj1fuMRyyRBsNlJ1nok3Ts/CBp9xdRrsfEnXWw1Lo6lbOfmYVF7wnWS9FVaG
UYT8IdB+V0oXhEy3gP/El61kDwJ6ZZ8gKOjXEaXQA/G6DpqYd6hw71J2ZSq5yy3K
9LfenOE+dvf3HYryHcnx/jWI4hIIvwdxOPf/Z6qLMVYfnYZMngSPHqMt4BLjrWXr
s5xBRP/fK+ghguA+31YIRWFmcgy6N4/aIEze0trHSRgLZBc0x3O359ZQl9yHd+Yp
lwi8PTaF9QNSrtbcIzea3B6PrjPVcHnZxgRMtqmilYkOhycHjocqQA9dJsD/7Wf3
8dMB9Bjjmt9Ht2Y/7hOr2tPJmbwHSBUr6nC3dj9kzPZk1gjg6JURKN4vkrgJDjHT
Lad1dO1ZGA87xiSzuReZ50OSXBPGWS2I06yErhjV5bY9t36X9UkvCGo2+Wqq/4Kk
bd0XCQPqra5FG5h4ZLYn/UiAf+wwkKVf8m/Up0+xvx4ZffEGX18QFYs+HTKlrrcq
cmaL2G7O70oMf41flcHU3iCobcBnIcpM5cAfrxczyhSll4QPwc8z/Ecpv6Za7+82
JcOU/3D+dVZCoXWW6ds02PGiihS9O7jof4MIGY/Uwi2uxTr5RxQpbbPo+K42yqDV
m/d0BL0rTNOqdc8/vLAHZ+SLCiyJpkqF+rnHMr6WXzY2V5/kdItBVxi9O/qCHQNq
MlTBeenYk6JHtZBGi31IugKRfjrFlotyx/kbcHe+OLv9w8u4NvmMPgfNt/IFaJz/
GIbRQnuyjYDVJfsX7jsgA+ut8w0s159NJ/YVHTGz/wZxx9UcNzn4dT9PhbOy9CHi
Xl0g40ONU4e2LIt1R64KYmWTWHsJjPwCl/pm37CYTAOEBgC8qWcyBPiEiM2haECs
b7badv96p9llR/oPpLhZ4yLIUoURx9e1TyN9cqft5SlxxfKCq9it5KOG/qZYq6ji
cDnD4jwjjBeEt/qs1jIOyujWTWqoOQrSw9raIjjpyMRFAef96rAzxh3K4ooJJcGE
d2Z37Q5ehbgdwBBEzqgvmTSuUdt15gaXBJl/itqywGzNmDgOqB/poO1OJaPBS59Y
3A0m/VhVzY1z8I5WhA1d6+yJoGV3A8g4hRUD5OWRLFVD3L2O0+WQI9cGcb+i45Zs
/IZPaBjX2MoGCvFaVu+RKsfRUODLVspMLenk474gJzG8sMXUT4LkQ1mo77DKLrnB
hUWOWSL2/ggaMF1MRAo835D4r91cjZTmol8gIyovYvUfQk0jlMyNZEBTWKM5G9Ds
2ZeYcNmjtIEBnHr1R+ZFPGlRkpC3vZ+JrrhCnasr9eXkAromLPyVQlLhkWe+20k6
M1lARlJvX8v/gLiqiqdrAdcIanHkFDE5LrL7HvyJd77q7YBDsocYnqO8wepaeYKH
rdgCZs/GQ56niMC8WWTbtK3Oq5GxNe+YDJiKgIFTsdZs+Vr0984Q1q+LCeDRjfd3
q2vys6mAg7WYwlhvqjbC72Jh+ipjyLRVsBmVK1iFKGMfKRAYQgjwaqlbGdMuiPTF
AEempZRFsH++Rp0NNN7TXkD0Wc6J/kRwppVgcLbOOFFQCd2ZAD++DZjVJVn9E4L8
aeqZ5DRgx/Py9Hjbk1nY7tD3sdwa9V+aj+HxT4Oh2m34ios96skix6WqAzolneKf
28z2vnXoVgbnnIJFPm0Uwaym1id8UCWm1LZeND2EU1Kt4syD1ujpCwigR1DxNU5e
kaTUerSOt92eMcMijftsn18EkcshrBSfHdJMCR61+475m2K2M4VS21gGhXPFGcxP
jWV2l1EWCHHjhRcLkCYsiVw3GcwZEdi1r5TEhgKbOD4DmLl67zhCvhOmpybT1v+0
ePGDcaxAVGSM174bddU9ApztH/YLnAQIOkejAcb4AmMjbNCXt8CNRMACQDs2LL61
EcbOhrihybZTQ76nOxg+SEzGaFi2syiMKznJOYSOYm/e8U2os43mrsBa+ZOQzw7e
pT1oAfbmX+ccgxPrGwXcDF+oJ75LthQQi+lEuZF0vtQ9UX69kJsQT4c96uiZYTXE
WvcpDDS2bqIIGTzPjQcqaf/5FXz/jRZ0kT4rb5HHIm5KAW6QMbj4fnyILlZHWgwQ
DcPk9UNC8dKLmoYdbKpZAEXYyy3TYHta/iWleIeARk3qjiQsVAzcobWWHf88dETL
Sp8kOyZdyNftE5k6bwp88ucLwhv1DwLMAgrlhFDoMI//nA04XUSHkURdnMMJJ/Zg
ywYiI+UdPoZG3wLagaeIVP2jLWlqGzD4HigcmFJ+Z6Z0vUDT6s3Ylo4kJYHdzGpI
QWVwjiiYyBYuLOWZ1feZkgbSy5bzaCbwyueSsL1blrIJQxVc5yfq4c6f34ckj6Tj
WjLd35V2gNtsmfveZBHPojMk1l7aKudP70i4HUvlSs9L8fnmMywi19sNvq+OFhtd
9TIX6pGPMVMZ9bGyohVmNr6J35KETtc3i5APtPQSBCYl9NoZYl9KZwpwPpjqkNaB
Yc/ib1twVCdWlBjlJIGjKNo03x8hw4y4t2GYuT/HXZYsbNjQK4AwS5HLhC0MQ7YL
RRg8qTq3STizV92CQVfsmhToSj3D4o/3U4jG8A2duWEf+I5C3U1stBajulGm+BCJ
sxuhJB/Rb9tKhdpc/n2U6GTUi1pLGUxi//v8rBOwPuU15cgKT5xEM/15RnypWeTq
I/Xvb0214ydfcMDyUAbOE/+J8voYgODpn3mHomvcmb0zBMBLfvHWEghS+3C2Ji+E
qiGCys87tyicsINMRJIGlb2zb3B+ikb6o3ii5xl4rRbKYwlu6l0TNjTHjgDs6NVc
oe7eDYxdLyviPfx7m6WFVC/YjodUUaPPFS7aL7Tc/HSl/I3aEwteaNtx8ssaEdwl
cU9eLmKZkDbb93L/vTm0owzTF9S/Kaax4jlZT8e+hF3uSEq/iA8Xw5ees3Th0nB4
gEDutEwP5+GOsyLCh7r7sbRHZysMNUm0WzF+CUBB22232ClvEPESlLRIizJA5bIq
vaga986q18equgxC+iL6DeRbbFNjNPA2OFd8/7V4IV9NRCOKJAnWnzCFm2ZobHN3
bhz2IvfXQe7DEzkNdAYBABRWSmIDEHSe/hnnULG6U7z326Cu4aehw4gWt+0hsHds
UGvTz2z/JBjc2MWRAXUuCtsGXGPMJNjeT5kDXqiGhRqNY4L9CUBoFUfIaIeHxkoc
6ZLpx1SYczQSDy3/YuSq1Gk7XAD7LxsB4sMiBQcHFZb/BNuV4zgdQDBLoKADj2s/
da3rW4vxOVZjMfxVw/v/0etKaT+PxT7UUt6i7kecsok=
`protect END_PROTECTED
