`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
idyrBWG9YEetSEX0MSxFH4AYSHVcVJdzjhuuGP5rzY15XqiCfWmPfgpkMCT3Pegm
5IQpmh9iLRXF4yTiW3diY9odQzX6TskYQdOsyC2iqaSrK3m+LYEClN8t3WDvn10Z
Ry5uyVaTlaY7nRUW2WbdUffR2Bj4G9oPrPXo9UnCIlRDF5+iwJTPAbCJeUKk6xWa
HMNFVgzUDT8dxcCsBL2epas5JByUWBodYxgc+b/zFAqxBI3gyclj9fzKO8QqpUL8
Wi2TNOJ8qIFeYBzXmgnW0exK2NcpweMT+uLSZePu8Q5WD4OI44nwosDB5DuHbJsq
JC2ZpP0YCyXNLfO/Zi2+bT0syhUYkSdycbp+9gHXAuwMGHRymC8TCQJ3rOYwf3WJ
W7kCRxLgdTMzvgGEXXqZq+Avug7Rpk8C4v9hPM3jQ26mz3VD9bonseMddhyu1bhF
bg6EgIEthZhQhOvRDr+i83Tr99YRE7h/bM6MI8BHJ8z/LX8PyckjmQb1nz5etSAf
hxBtD/eZVmkPV9oeexsMOuacIfG7hBtB84DnruUZvya0kDGNesrQ1anYTI+8v8DX
JpUyQaHbJ/nrd5zGojslpVrTyVxU0nKGwHpJEvRnGd2AXmKMlbf4qkN/Ny6IpoTM
E0aTH/W48rRCEcINT7mZw4KNS+o5SQUWEic/hxlsqVo4dV/6UisVoUIwx0jKJw9c
5+X8IYjApzT4Cc7vOWGlv6aHyONTPim5H+3J7EDNid7t8RJkBlKvP3MsR59eAT0v
gxWuq3nbUP5BfbSeU2J0wSY1V7gf/wReiCfSLYdHWoqEPv1FwjaPcT22ds9zTvCs
k90jzQGOOlvZtAHLKen3aGdYD0eRyvieqRYRn34IDI4=
`protect END_PROTECTED
