`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7gI9B1JbkWUp2t84l0jVjUNONMoA94uoTtKOtB9VLBuUdm06g20DeF4GYk7nbBah
zTwpfZmxYkxUQHNjogX5ox0e/hM8E1Y5igOuKWEuTEwb4wcSeXItAzqYSPwY3WR5
5oT4y6GbbfqN6bhoozcJhPCkXNHsANCrVnTfSwX7udcLgtEuI1/iamCyonZzMXN1
6n31KYQ6hZuWEkNIrR4iXig+TLP9BiHFHOXpg8gt5qcBU8GLxwPEPQIL9qCA1qGA
uNnUBh7u29EdAVPGwPGB5hAi/ehmwCDck+wM2oifYew9I7aCJqwrrwQEpLaA9YIW
K3r7aYyheKqzMs1m7D+yAMCQih8Psmx0laB6OHkfY80I/p8EPnzAHbSRq5CSnRfu
+O4N/uNG1P34OzbZDQtLtw==
`protect END_PROTECTED
