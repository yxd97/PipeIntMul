`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufnfMUoX2gnRctTUVVKRdGm2L4yM//zuHzCeoSMp1g+6KJYmdqNuzgCnXBZ72VLS
FHeHLJkO2uDxXVM1OVe+je0I4Lq7uRohxVa5UtVewa96ABP53IV3pQXvkJp8roOH
acq+R0t0Gw4zAKfPmM7GcT/ZzIOy2JKdygc1/v+mSYpi2jT5QJfLwVNPtXH7PTAM
ngOIa4Jxkv8O3f9gLTySqtk4kUE22LvymMD4UCsAGDq8dxtO67sinOpaU3NTpveq
CZ+wbuKbVRfJXVWDO55L4v9QRJk713Y9vV/UkNog08A+6ZKdnt1sOTVErcsDq6Tv
dS5ActU7vCbykcubS+mxx9JDjTrzIyrReiF3iPtvFXzEDViiAUaav/56BcDX8sb4
72X2x0gTMpm62He14s5+6q8e/wnC897mwqsA6oBi6JQYkz7BD1m8zKpU/38pC298
3KU/0/nO9j0bi/r9Ol9WHw==
`protect END_PROTECTED
