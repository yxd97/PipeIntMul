`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tlv6wFDdBKsQ2m90pjyscm9oJLvMOsWBu+BdXQhKgxZr6WpAToXlp3cBaBR3+Jg2
Qb97Hsiaf2XQlCqILPMw27Rs7+Y8zQ91naDPq9X1HXT38JOLcXq9kzu7THxFJrFu
n68x3IdypRL/8oWEJpGje2pUIRHDTARSVGwDFcgAS4d9r2xXj8OgpdX6iPGWKFuX
cXqGFCha7q5/re+6LMrjxOVM7ycqvrT6Jahlnu4DMoZqnevxxJq1gX8SKU2rRx3x
ybpV2hM9SqjyfaYJW3rUUU1M85eGJm1kB4JYzDCeT8CB3aYtV/OUUhlYsLmp5psN
l/RM5lggwMOGFnMOdpK7hcTsDntXmEloW527a91n4YcKLaIhXxGxN67EdBGlzHkA
06ugCDM8FX1XP+i2SlEwrZIEy0XQJDo/IUl4qFXZqqiLTFRCELM7i12/orpdOfmQ
3dwPcUdxPxmPR/Pfiv6Ho7CLIvb1pRGaOzCvxXh0d9B2pLlUaVj6fieQO0nqTwhC
Ea4xAvuddq4JAyqEfqHoOp56nMWbft6TEtVe5JYc6qM1iE17crmfocbWlwOXnfq7
TD8Xr5khoqBFdq5R108G2XiMLDrchRJCjrQSqVhg8NuWRvMRWAgY5sANXciWlaw8
gZv+IH3ycsk3e03jd5a32PDz95AvRsJSviHWmwwXuXgA0PGTbv4MIFG7W+szeqJ0
af5L3tN50hBXKNxG9FMHAnK6fR1UJCBTPgdzIHJT0XT5T7sQMA29wKMlBWMNjqpB
`protect END_PROTECTED
