`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJZs5q2TajofiimOPOqV67vvlU/27lKvBj+6Q3xaavk3o227am+5qU/Zpwrdasxx
owLjTQty4uyiaVEgvIkN//aBlBjQ9V0qGCQJ4o2z+KrGeaMBfSulliK8/HAWG0Cn
ars25o3mH3CvqIHWSOutxEsldw8pPvbrWJeS4i3gmhFOEL62OcQuRvd8EFAuRrIt
iXGK6n2XScR5TN/KJRgXIxJ0p7bHRjmwtBO1dz96wohehWsq8+wBCt//1om56rjp
N2rt62TQPP1ZYmD6rgCdvhQA3PyjTLb/CtdNeTBmN5jglPkBB3n9yQ+m3izzx9jP
2hWbUGoePYmyB/J8lCjae1o8dx+EQx7CJ0m+87PUqo38BGv455wb6vyOsmbLDpPf
mc8j3AEyqqLezgAj1Vtx3ieiBa21PFBXQ8ZBZbINtu69ZUwLtDbEPIlT7zYnmx21
WLdXsltXPycHlfQg+FR2WB1dt381u7JmURAAVhZ0gd2sQmEIlKglN6mJF9na7uzr
dZdOlPRhKwtrLkP6qwBNAliC7pikVUnNNaMPan1ioy9E8x41hNkhgOoKkXtxDkrn
54fzSwr2ruTHDjaG3JIxQwevhbY2q9NCoHznqi84oIrT5/0OviUR5YW5s8cpgQ1P
Zb1vH5P/b10FWerc+Hc20dr4xzKf+9oYEAtGNX2c4jshyX1PTRYBDPlgW5grAn8x
3gfK0iIRwzWpWQ6ZJDr/teEYe/LCJPY0SSdI5mnTcvro/681c4X7eiHW5Lonf1fj
5T3TrlPwEB2DctXTALEb4Q==
`protect END_PROTECTED
