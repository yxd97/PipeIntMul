`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C9E2SL7k9G1FjLILXsUWr1yYM99SpIAcWESE75teW83eU/JA2nlQbfDbDIFqc5+i
nvsMlrQB+4xDPmASEPpt+hqNeZWQXtJCKPuDNp6gPs/f+WIC842XiKeb2nCBsr8s
LYsZS2Oe8DvdrcH3lsR3ut59s1nxkxX589HjB9q5CtiPkUgBW5a6VnZsXbJsRkJB
j+CtCANgLfh/Ey0/uLjowe7LkVRelRIZPDfns5/Y9cAE/ygutH8f0UCKbqZx9IqM
swRh8d67K8Bv10LcJ6xcMA==
`protect END_PROTECTED
