`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eqo1a4Glz0jRGGmaLL9wHHMQJP185+bSc5CxS4RVbcGpVBSe2p6Z2tQ57nWdS7jU
b48TD/63fso2hjneuKLlf+95ZxZZ2CevebWQNVsjhSWqYP8QKXv0pCHaMzoGTlHp
3eCaNOA6/ReFvVXrMEfBlXcbt8devOIhJdgtzOKqrCiQWA6kX3CIPIHAWggJaf39
rJJOBCjvWW8TAjamSKluOykcotv8GiROG82iOnOB163qQm6eIv8VzSULoMXBy8zB
xqpBd9xkGUWyrMZFwdsXIigtP+xj+eL41g1qlFRmvMF+Mx/aoW32+GfTGvfT2YTF
tivUpLAyfJ3rLqRsP2xrkv1AnHqKKXmdCqV0XDkOwWtj03i9PN2sF0B7UDReaECZ
yIvKDOE8eo3qC0/nOteB6qiU9urWpGoHLeZuke4BpC/rIhXLRoI8aPF2yESBpW/Y
yb6kEUWd0IvBKvvQibWDNVONygQaHagWaIAJKk/Y1VothXhR1M8RMGxoMJ9IKh+d
2/K7UN9/9XEMz/D8eoNZPrjbD7up6qSCZTfrjcrlUY3EtHIYRHUdqpXNPWNrVj+m
geY4gp4JAP1Y8goYM4kPClZS/gY4CrczDVIm+DrJfWPDgI92ujbFfLMrlHm4Yaor
/Hp6dNwz/6lxjS7AvUusGA==
`protect END_PROTECTED
