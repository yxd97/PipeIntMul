`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDfsM33potV70IM+kX9xh86nqMrmFG6EBfxCpMg2RoyGtyilZbrpWe9ex96pJd9V
ak8hQVYkdIKzEraUz7h4nxELteBQuLnNlrEX2r88iMNziNMs6fMxZUPCJcteWMpX
RpAdOLlzAdMQgE4UflLIsjmfoDpzkzgkYjBa2rVDXXq0f6J3Bk3SgdvtS9RuTyi4
9QZHgALjXPUVX4QCrXAzk45aSCajF9e/S2cfmfRRzCaMm7QzNx01bK8uzb5METEI
zHdgCZ4JEBlm3XU/4PuFkT5HPghv6HV53Ujngff6r+Fj3cDWG5Ip65ajwiWJ8rsG
1t5VFtwdk+bAQEjYfm442Rb9RAdCbW5nA7IQv36TUtY6ZdQDZdF6Y7Ro0CAng669
J1Y1UbYMqgNPEA34V1ZoyHEXTjzNp6TnvlWMr4YwX8A8d3oDJCYShsHhPmHvNe1/
pN9tjJOAHwI7WzCa9y2IdxFj05/WRlh3lipoTne+MQ44QsYwXlQYrjA6eYpnT0sA
QGU1MjsafCOBaexPMHgT+9ZlFimeM+HAQqfsW//IF6+OgEiynMCNzKTH/K+tIoow
kezPOMZ+IUbSwF+qn0oj3MYSqRszHQCMBleFfp7PLgMdgQ8qjd5Ix9rCdoaJX9uP
FsJ6eqctOzg1/XcJagL5sQ==
`protect END_PROTECTED
