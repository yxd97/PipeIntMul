`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIgakqpXNUgx93tsslYCx2yQuLQQXWZEO4G130qHnfbfPg0Ndm6ok0N/abNpwkv8
q3o9AKe0voiXKpASOAiOjxO5YEmxOcOhgiW225vkSXnfLE7f/X29iJHLC9amm2oc
p0pWvrWDwqkvhcXM4ke2Wd8E1WN7eODkPc7gPUB2WKOJYSBpmuEyw2+wleUAYhaz
RFfqvnaqQe520DdX4rrkP88NXDBpyDzgXY7q8sdN4lm4OnOf4cR4k2GOgul421t1
ul67TZr/S/drC2XhkqwEdF/DcJA5vy8mSsaZGXeSQydpwMV6MsnHF9rwnFLWFUKh
twUuGjDYr61qB1j22XzL+ytom+Hy6TLqTja9aXLpGSRZnLz2yI9pLkeyq4PxHIjp
8fqZwomcoK7ia3fzvwnNzcwb4yACnaas5VZSe8egUNcv4xLkXqAqc0OEgyNOKLGJ
54AovU0YY1nqs9gbEDM4Px+/ygmUMDyIRAkj8h3fdHQF3fUKdSlaPFYXGo8YBI7H
KN6Veupg2O3iDQ0azgTHpnZs32DfPMjdJC4ryOp/gUHa6ud9FNgAmne7b14Gfc4f
2sIUE+jslllmLfBcT4+jr7ppI0aHzxCZ3/nNLG8zA9Y=
`protect END_PROTECTED
