`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4MG4TyeGukxrxtfuvumSBxhL9LwELvcMNZdic47G83b4zZPRyL75ZLyMKPPCWhtU
N7BBE8EblwjB+L72lcDoXQr+SqeozdON/IVVp1Uwt+8l1haKfgnjIYpT1zZK/7rY
FB96axQJBgkTL6g9awXy/moAX0Mtu4YBLZC/sUzR8sH1h7GnblXHEiKJRqc5Fp9Z
RjvuRliJPZMkW/DlxA7+W9a25NJbFcdcMyg3XnJkGwlXkxLK3Z5qhqI4g+bvdE9Q
vvoa4vAavwU8EcfagjN38Pqo4MCtmQ1QR/+4QvBPs8oa9mWBWhrZDB5mXIPmSk9C
+EkgNn1jyfLwXk9EHXILxAHuAuFWg6uAcNzLxmvjH2qFbLVForhAW9wgBMMObHjz
Aogua8A/CB6suRfKP24eusDg2zeIU1jlWuGb2dAau/pE7aXPdKbd4KggImxLBwUL
OgXFV9qMs3CAwy/2+B899hM54WyvN61B/Ut3Loar7UI=
`protect END_PROTECTED
