`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQJDN3u9FCKF6WWYZt68v0Pz6C3ym7TJa4jwb9yZdzIFY5QvavRZIMglFaDNdxMl
CPnTp9CCk301xrtxFW8uCJrvaemZog3t71y0d0khw+9NLtJ9862sP+EI9qNNwEbc
YBcdW+RfNo7u/g+gQ7/72Ar73z6u+2lfS1ejVhF7anFvMoR61+eiGbTNWh7HMmwu
678wqHt4thqyj1+haQzCUihUAfVMNwewqYZ0YNLewETTianGJ62NnxVR45aEdPe0
PgZeKTMcUQ1glsOy/+VIPzeI60jSKzMoqcTTpFUb+/LpF4++DKsUMC2hcq16GsG6
hhMSJ2c4Jle0Qd5GGdp1cYNysY+FpoPvdaZEEvHy/CTBDHV5o43z/hiuShFhhby7
Ur9LSTduRfO2WuFZgyZy0ffnDghlbEr+H7OPV/YjwGtCJ6lJUQTtOg4zq0X5C4EF
WRl8jgolgni/a+LyOht28XUTnrk7oV3uNPAUz16bsqxfVhZZIiykaZJpKaYi/wo4
`protect END_PROTECTED
