`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qd6q1xF5Ej3cKw/8qFagBOQ7FGvwPA7kX1w6C2MbxFV5XqSHhOtR9bDv5VnxXMiv
k0abm/vKZbVyDv9DornDC9pB6qCoED2WHek59K/9R/ZyzZYTfb7c2aM4aweM590t
mnnuBMrP+CcOwslfbJpK4/9KTAlS5NcJBwmUub7Q3XOVYuMMTYMwzK5/yM2VbCdi
a88U85/mgNx2mpu/KJKla2AKyIkmgsXSESI4HAQy8awfQOtYzQvGGhy2yUUVWhgW
n8gIjfaHdZLKiwbypRZj9QytAuaouuGHTxHcJIlwCrjpPeNT6GJE/3L/XMIjnxmD
LXxHoWUqIKTq1/Dd+I628KbHlSk6Erc3n7dJjErx+VrrcplDtxcbkqi8XuSoCyCZ
LMwJTrg9qzESQnnmQXas40zl0k4dy6sp9itUupy9tNjHjyvdcGwjILvUqq3UhQv+
HIYAh2DLovWWfH1znDvymw==
`protect END_PROTECTED
