`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kr3zzcDeCIhB1AYLpD/x7tT8XiOyKo7dxH+RaHUGafS1YS0wec1ohda2oYYfvG8I
Lbx/PzNu0pQO6SzPWye3I2gDBzkj1gnjtXGrvpWkpm0lm0g2ct4AwwMKs9WBPT/5
oHVmFtCAMmjhvh5j2AI7OggsGKQg++0Abs0pdKbcunW52fprMIMpro6gxZAcUwO3
HppNwvpXctaM5nqEi3ef3DG22uWTIKWWUfmzf3Bm8bd/Y4CcJLHXB9jxKOcLeKXj
JvF/v9yZhDv+X5v2dsSJcQLIGwOimmmsacpqZJ+P2BVbLUM9P6zJRhz70VuG2b+7
LA6qNHpX6xcyC2TX6tujGI4/OBEcirBYIKTQgVIFDX3uXbmech0kFQq2H9+Zh4z+
AeOWWs6XQWQNvIL26Oc0gA+xR5jDgxUHIoTh+MeawUE=
`protect END_PROTECTED
