`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQ4qx5kFl427dsCCv3peTqP1/MNDWIc8Pcz3ZaoDv/bXPQVHvL65OcnIcwyWNy0D
twyDeo4AU9TLzH4zeZFGpXoYp+S6762PEVYlpYjagtXOpaXvKRT9jueMaG6TWQm6
SZKZtPxSI8k/4+DN4lyW/te7BgJNUUkqTdOnnx1QaEZ1tEnHrZOHlm7iwv7y9FTP
s2e63pUmZ+unubohdxvJ5Ego3YweswjL555xvu5apOHsts5dSGylhW0qqKRhavYs
08RAUfqhTi4+iMTqqxNsqojWBAvY/zT9zfr10fRey8hX1eqKa2LMrZV5hZwVGo49
5SwGZXfN9tC4rpdVFor5mQyxBqiqg8u91zOdUYf37fg=
`protect END_PROTECTED
