`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0NzdVrBE2BxHIst6PEtXEQR/f+e/iRHItlZJ5oPzw09/mGBW2Q2CoHQAmdAQSzAv
/FT+g4579TLSMas6Gi++MUsPLHRihKU/+evLGegR9jfO/07+vpJqXq7yM1jYOdA0
n4FRWJkoSqVjNstcOD81EcogaX5PkyBigIUhpr8MIYq2ig2jV2enaLZ+JpL+6voL
Xt/P6C37vyU1gwit5sjfi584jJk1Cug8YA0MyBQOk3CcML5mFSsixAbma7JQsYXd
GBcEVGg1GYCrec4vvIQC0scPcuXAAoT3DIqa0aSgjaFhVIAOM4hHbbK4TXak7nkf
ZIXZkGL/xwezRcPPGYF69EnC0dUeKZCeNqt7ox3zrES0ysG5MqxlGN8i6pUjlFhr
QJKbBg3f3LgZJydlJyLqxTlsHB+swf24tiMKMdk7cRrPJzLyn8w53PQYiyx2DsHA
ZDZssJ62KI2Nh70tsfIEW1C/SkepUJJAwh/83Gd7BLIeK8oly//mJgsEDlqhRbFR
XaUtGGzkW4+T5wZcoBcll2kvlzP7sSlo6kkiMOIp4m2qGVWr01bfpVcxLdpzpDxH
j6gk6VBkoBhRMIB7P3CaMw==
`protect END_PROTECTED
