`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQB2dnUjJNPz16fzRIDniPFVJpZML+K23ORDeGIzQjh+IVdAG2lIwoSycRQTpYMq
y04GDRMXuHd/xnLu0t3wvqi18IE97XLvaaEFV/iZTSSL58j7eUhi4RElGjc5Ohqp
xOUwi5A7X8hg1Gqjo5odXwvifPj16GDKJSmRB3zrN0/quM/ZIDWLxI0tbspcI8Jb
GqSCbh0o9lefZQCT2fZFUOPlPU7vnoOVtCEQvEPYye2c+Kli1veeG0dKBddiibO2
bKN4uClYCLpi184x8OAks35dR3I4oT5PAGMLa+WZuP6FbLktOZ/k1FYCC03NDyCY
LjTTwRhQPfIyCqs3iUK8ZqGrgrmXabOiFpsXUuqNBUrr7+XbCnsfCIl5iz4nyW4V
9Zqf7ZLlv8b0lnqpD6RMXeOBbXr3+0WVzfKKZEqBY1gcayY6vryfwc0cygM8/4cd
SHWZI60ZzgIUGnwyCzixFFV6Q2sfqYtM1EV8Gp0VXtR5XEsMdHNbjS2uVym680Eb
`protect END_PROTECTED
