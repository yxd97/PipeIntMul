`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMa1kbAt6sd29u3fmOCborSvBNJJCdqXjbD2DN4VlExcWYvKlgecOt7EPQKtT5G+
EJ4ltdCfer/aaDYi3BX2g2zoqgWlBD/XPxt38iD59p0Y42BDO+iKIamhoop3HlZC
v8Y9r4QeCd/M02V3qZ+SN7XV8LOWT48L2h9LezzrjzTS3GtMufHXxj6h4RM5pD1b
GKBGKBxw+uogNfgAZmwuxesbzc2AlenvC6KaYUL0s8usaC/+GjVjL+ytKUb8FrTs
sQajuxVkBKmMlWp/D9NWV1AiliQaQ2J9TTPrx+vz6mg=
`protect END_PROTECTED
