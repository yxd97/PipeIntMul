`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IxAKQ2N0POyutdYCbiNu8UtVZQRTVIy7DTzeokJgT5+69TVjNP37FyMYgMlYRDhU
wgalubwpc4Wg7EdxJ99bjdHntcV8mxuUFiH5T2oho1PIxN/9VRPBAoAeGqLY/7Ip
vfUCIXzouJHvtoyDHLfUWPWygkXmv4cv/BcpiTtYSFiXaLWW7N5SOToAmWnqoXo/
Z8weRfkgg4XNpRGwSc7+0c2kfbqH9k7zrI7pxh257aglOo/YlIsVtXd76MuCejLY
OPE4I4vTKT95kDJJuYZdVDax0vgdYHgcVcqQHUPmJWFdMTI654BJjBLSjQF2PdHk
dHtjFhTH+9l+Az9m2KBPhBHeXy6U4cZF43mn3jwodUVISooCt+rtymAfzZOgupdW
LBe6ktrBKzU0XwJWqK3tV1mJhUMKTjQm6iJ1Hm3OhipUBbcWFXWEMTlTVumtGoSD
NCNn8HbSakfobsbFYAGOLFnMk+LMiUX1Z+0eW9C0THf6bsn8qg3iJi9von6+4n6n
ZxQOy/525+aK8ZUw1cmglS2iLgf4jzNj3ZIaImT8pz6lmKBP837v6NedxdPs3eKb
aPH4I6N+/I7vfEa5EobT+u2YnVQ1I2pwXUt/NMFcZfg1+MmuCusB3mHJpwNLM8w8
3/ezsu6aIwWEj9xM2ST/MtUimryJ2mw4CxNnukz9+EdQ3oDMHhWk4C0/zX8KFclH
Gyk4JS0QGhYV/PoajahrjfxjyRYWJUBeAywPlhwp9D1OvVH42VYSl3WrGMxi1vyM
zdBdNxBgizABGJtcvt2QBvTXJL/a/AdBVM0PipCbVfiblB7qE+pskcbkC7Lu7rNo
Q1MAJOYmh5K+QiW3IAIiczv09cpoTRs0FZw3JKor0hPGVp6KHTDreedr4eYkcSJG
5VwnchsJXETw1saOTQopg+YCfNbehJjqRaT/Ylb0C7nLIV3VwVRmhnSzY5roIeum
G2AO9/2msmqNnUasPMcRb/MStxSaF0sXtjxSe1Qylg/FP5tbRFCrL8xhGe48YQVe
res8G6JCGR6d5fXPHb7jUJ7/fXuN5GBtVdnLUSm4BJYRE5F0qXNNK/NZ0T6EvLRQ
1UYtCeHhltu8Ye+xoJYX2lEcRtpkIwGEagE+kdPDkLZL5LbETyGKCIm26rvgwHL+
urDjnQL8Ckk1RBFXz5UmyuwhX4+o8YcXO6lBhKaUhgZKeBd9zYpTBtgQheDzuicM
il2LftY2nGhGGU/OIlCbW430HBgxPYL8pZ44OVHTe/FNX9QqO/936up2dd7XAcqC
lSNdV7+SyzTeMGWqzBMNlFzTHz8ct12VExTKbZ5YyLla69EHE+FQe1q0nT357qh9
g1KsnDfT6crMDi98cTZKocTVwbZFQFudVQ7EU5rdLIbma8AlXa/xzcN93ItDOUqY
KU1yVCsM29W2DlL3qc5DJTNt6aD0Y6VpcmP61U/tfjY37I58eGzWAsnLRmdXjsiB
0fls22MXnbxh1z6D2xGOYfX3/yqWJ33I0Bnc/gb+MAqA3vkOXWENJ9N37XuLX9yQ
ojgZBXZhlgh6bw42Zh0nUoQc9znyxYy5UZwGdB36iY+P0mnTW3j7Tm1Smrokgbzz
pkwjdZPxd5TH5cXvy4R3rQg+ttlyj8AuUFYnDQrSQERSk/RAZsHr6BIvFJIujXYF
qepqEmwV3hutIRl0lLJdwEALS4zfNiBFrx158DmvxjDj2cCl0/xeT5rtleBKe++5
QOJxfP/UvTq62z8WZgdcM0Cihldr9GiSONS8JkPX6G54c2Pw9JPUwXCFBBU2dbK9
q/0LPwYjjl/E99+2LTh+EgR2FwD3OU9ttncWbCRko2OEc11o9trTt4H/WTIVXuqv
q69VMgjxu2zi43k18Ov1Dks79Hr2fWx4JxJiZ5jcvvk=
`protect END_PROTECTED
