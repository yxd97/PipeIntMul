`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cWKkzI+jNRinYz9OccYNgWCcMmkT1hJqBEvHnuux5SDSQAjEwdz39DMMBdegmPAv
U1QQkxTkht172TVysc7MwVsF4nJTbuvHB+PyVA9ee+YqHWrjFvbHZ6radic5X/q2
VuqZjjJ98vz45ipastfFEps6swc+X+VXcUV21zqe1sIPm2Uo2gwpd5pAJnT7jAQH
gDXbjh1G1rYRfqlsPu/AIGx30mw+zVVgkCrDMw4Bb7DbJl9PkSb5Gngkd5/2fKcU
M2bhQYTfZ5ylxqcSp+zSCpdfUl1yWeqjiH8zIGVXPstx1bTQugGoEW3psPc4vpGq
bayp5rlN3TZlMl/Pn2QTzxNoNywlslOw9vVRGXM/bnLy1Ty1EO+EMvTI+0R9MsUQ
+gKCYiz8GOmXrTA8CJXLqMt7530s3QmlUiwAxYAY2lvl1syYBSMtXUr7hOHOyb8z
ZlFyuAEqnKBDJb1/VrtmQ7dC10SBnAgBUMrm1HkzHe7uYplvEmceRM1sQJ8B5kvY
eRxcbU+TEgPVy2HESWQKKlMduMZ8CYe4+NVROMkV40n0wH4PyhqmDd7469wWkCFN
U1AX1CemOkFjulsmhdE8mDrg36rVPWtxd37DtEIc/IA=
`protect END_PROTECTED
