`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHExhAMQuYKSkxymY75wD74qebKKDCQgtmT3F6S2skjGDkX6XxrHomJN/u6A/C+l
QrOrGWZuETAJRhfwZjHdFrNqXzyRRn61OpBSRDjbfoorlyjg0Gr2pkvcWHyj0KVj
0AnwbVtaHJM6wlufCwUpRpdCQ6VkqLpBg8pCTbBgq0G1EU+EhRRfryKPPvc5HvWK
HwteW4e8DwwODIimgelzbDuuQ/PBn0hByTSWFzinChYWGilvYEn9U0rpAVwvhvUg
njSf4Zi1x5rZ3V7IPI39TL9YnN/3MjkxoZnzJ9V3aKtNWm9hUqj4sSyHVE6Kuz39
tu/mvt59kS3qSaWzwWbaLnNiFleXV6TqyzrSW/aTV9AbbpZ6XsWB41m6RG42sqOZ
9OfedrDjkDokOK7mG9QV4KobWs2wvkjOhvH6wqmRrM61CO6Zh8whd1UU87cUcryQ
gdfFsumZlxG/DwH0lMulRu0wyfahVGic0Zevr8xk4DTQmnqdl8heOxdrY0fGnzdd
k/2Be7T2vv6U66UhaQgGEiUUx39BnKMFd7n2b0c/ExnFO16opFNzXw8ufypcbyT8
mU3bQKR75pnpDKmtrSmkL435GkNZYbAExSZh548IJGJpfdp/hWMNQlmPjz3b9xsi
yqx0HvyBgEBgFAuwuOye4P0b/9nW+ypdSY/vaQFm+CYUpq21evA/pdU9KO9UqnSS
zvLDRt9+s9dTyayvb91czIhiWVyyLW16Y8koAKRrmAt7WANwPPqhEl8j+WD7f4Xr
hPjaAQQnfkCPhbyPUapDUKWPR/42LH+WAGVn0xbtimJX6nV3ASl5OP5P7yZrHprZ
vcvPR4WMlNP0+TlUfUGQal6UzRWdhciVgo1RIfOXM25Q/KyN3W5+cg0yG+Ttsjkf
HgD8kQa1sSAfFlN9IexyaoU+b+OHhcz/RcMoWInngtAPz5s5pw1wAfDupsh4glcb
K9h7eQDzi1Ks7hhFfoKu35HE5iaDTQgMkqWaRcd8msjjNAdOV8b/84r43HVNMz9r
U90CWR4t4SaCOsh8mcWbXNWdG+gdKDG8+zZRGPe22HnMPQFnArYw4N/fixJq0gmA
T4vI4Yu4Am4l5ulMAqjIbYXJwUAQON0ck10p669RJMFU/Pws3eFTfqNA9kgbfMd+
okU6OrvQm1m3THMGBudvlJBVnU6mx81OcmUpxRlF0ARM7Pe2EZngirFisM9ZCpwx
hRuUkzPx44jhvk8FYodmNZXWy6SUlxW2vEDJo7TetF/F0SXsWTvY4Zxk4Q1fUO66
LYCF8USX7okjkI1+T5o98CPX99TFbbJ01asAlkUNrMA2zvvGtvRHxslH2PlB0Znd
BbC1leFLuYUbSc8LNYsZqQ3TLofnklfqo8KRQcl38NmSDB8gBbweFnr6MvBbGgq9
2sEHUwcv5p056HkRxWf+bncTNQ7h3c+GP/w28m7o2wqsSyDpAS4ZA7epH909NzJG
MorZC9LD9Mhcx1eoU2YOgiBzaWEppav308UV/4ZJxZTTu5JYM+UWm6MZhxKiD8v9
6tMYPh45TPEIULpQ8khJdi2clARi5yV+hP2PubyxSVAy7c9fBHGRmspwHvREVFLO
vdknlHJzCQ/CQcPTZlZ6DGG2snWe5/egLUGThl+jykb1mCvLSJyf1TKVnL7cm3+y
FKetXOhYWH86pvDeY2haJOeceDgJLKyV42unmv8yOQ9lSL+C4h+UqZsLUk+cMjM6
Rq5F+UH1y/PqyVboWnfVqz5qi89+Sxbhr1vkagSTN0lI8xYwEdYOYBoBxSMiP6p9
GqGNCI+iR8caGYawjyNSHUrwhUMLr/86UrBP6H3gQKKs6CWK4PDememey5PDBvN0
pXC0T0iNKlPVOXzscD4hdkDhbXc5fe5H7rC40AdHjwer3KhkqNAvYwE3DRyjXcnT
TcE+gwe04H2632P8xO8maSHXbM8DMYYjKa72hOgMFymDJZC49+t+2hLNBYp89Gsg
Lc4CY2UqjkUPlxM9Q9IIen/S5vRG8+GW1oP/iVrWllooPggbYiscKPG3lQMfpxlS
O/kYysG9LJ/+JuIB5BfPfqVGSBBq9iPF2ZW7QRtjerv2+mqiIf/C0FdknR0RJs1T
SQZ0r7qJqNnaw86uXZ8+Z50lcKDoVz0VhcePjCt7f5X/LeFa38saojbuw+TnHgBN
4/iFNAjFAObpHQq3QAwPvoWoB226/8kl8ldguI3vjSDJefoIHErtt49CmtXgmXUI
cBpqeQHyhFr66gVpebK8cHB7FOLPpOg42diBwUb63gUZIroWWCMYxlBBQ/nzGthA
vL/6fskDQ6rdlGDdAqG8oHa8CSHfW9Ypde3XaE3CA9Cj3bQc0SFrnyIFR/r1X0DD
eM6EfdoJCwwzYERMtu2vxkhVcQgrwckiWbcvjhuhKRSVjSrMQ0BldL/SW3jivdag
7BSMKlWgN/mWVEK4Xd38UaPLhmoEHP+XPiV8XuYlA03iv6GJR5fIWOYNPbRYI77l
/yQDlZ+Iwbe48b7ylSUMlZx+iH5OY1Dbg0K7E+uJoaHLD9JmxH0ueiBLlOAfXpAl
iLtj/BEWX8cRGo/Texw0QpWrE8s7B7EPCmQ8NLlB9IRJaAj1109b7tAbpzzUlyTf
GGchQ6wY+8xGzxJ2ogLvm1XhLzTj91Nm4WxqJiwHqxHRFI3UPoyrJHkmE5di8odD
xn+6ngq7pvCsNfcNCA3THgHesFrqI0T20LAA7YFGkJftAO/UUIJINba1JTQv8Otl
gAEg9eDPn6K4JVrmB3eTmC7NsQO4RdsF+0Om9R34CkAAUCvoL4z7rDoTct6CqHVw
mye1FB9/VNcOpJJ425Z7B7IPvacc4DPG2AJdEwCcEABrrY0bepzsTqL/0Df6ElWg
mTEQjY6i08cz1JqVXGy7Uwre0uIrChXml+5W2Os6FFW9+yvjQ8YOl6PiaT38xeDc
FlTlHexI8nW1P9RJb40mS7d8NykcWWl8SDoZnhHQ8eRND4vdmd46q1sW8Y5FWccj
pNiFumCh7Q0WMxF9Ih0tcBmPL0k/I0BtPbh/yxpke7PyJ52+Wn7iUrG4B4rLX0Un
NdjVhK2DZu2pMhclLmxZEMPZnAWcUNqAlUbd3+E4WlTUqK1y23VaN/FriJFei6iu
Xgh9ccefgXWUfOvFYAAEhB8kr95bq+0TYPd1a0r/bikvxX/HQwLfQ5ZNiYyq0dbc
bxU5yCQPYSRpuzGdPv+1eyqJzz0JMpsaEy3i2U9wG4Cm18duTSBmtgd6CpUBQdfU
BXwR2njDtDt/ruBeSPcuHydDMGNW9R8rIF9qGe2O8oT7GytXndYoh+m+6T0o8Rlc
9VJzFv5p+ZNIk6JNTAnRPx7vSUewC5TkJ5/IqBay0DYE3wLaCaZWPM5G9FfLt1DH
6ixyDZnHRJ1Nz9j72MpBPpkNBEceN6OIIiomFFI/jWHWt5xEy4NbhDdESNnwKdP0
cbF9u1DrLd+OTOnAA9iDhnZ1B0eJA23fJjnhIE6Ren5VOGmTjKnxFjecPednd7RW
8na0BLE8LaULKonI1mhOQNGxliBHHctxWaaaODFZV6zfDM8nKOzF2n3495adUiaM
oIXP0TaPTPsFKHQ1f+dcWXkc0wyjK2ckc4WwBfHniUQoFVzzBP64+yDFrOGJA+09
p2XohANJO9Be6jWhCyQBAKUYwzOX0iujMkEQu2NMetD6oyvjYFhRh2rNi3U3i9fp
qs6hDJvBAevz2kALOxOmTWph7cL4dWjLP8nC3w4eMu1o7piiA1v7QX8ctCkw/1um
ZkMK3gI4X6SBUNkHJaLZdbYKmexijRg8sbAf+GvDEvdSYbefnjLLpDYv+PFD+ARk
qu+S1IIPeVOQjU84rZQ/qp9uFtA4+IDPROMPyl+1NepardG8t1PPKlcG6aJvc80q
Qh9voeXz1NGMa0vaozvnG3lYMrbh5Any0VYkZoamz8bgYLNvE+YxKtIWI83/rHqz
zoJwc4q5j7Cqt1kMNwhEtgZQCAy0xG1gjN+bca/BXYT0zit3WW9SiFR/duKgFiDT
jdPx7RCC0tPGsNutKcnCo6IzsWp/Pe8Oc06sPLQX9T9m78dNGIM4Y44ghxeUAlVl
NYSIwHZzpiwH4c2H9nsqPn+TJ8kFWKVh98sDVlB1mECskPTN036dRWO62m/CEvUF
ECKu3SrieqLzcUYV1b1B7Ot5mMcDB/wTOMz+8U7I5JUSvL0XW5GjnOmbRruqKdfn
c5YwNaFfeDmuCrehN8K3QsFI7vGYCKCSUU9X+xLToMEfmahnjiEMe1AwTlST8P2b
85bsBGlRklwDKA4uNyt36Y24S4bdMbbaQQyEWQz23Bzy0o8D+QwEIcQjstiglZCI
XY58T1gQwFBtpERWvGN9cuZOTuvJoh0rlLq7itRpFMJ6sJ4FdR6uGtcClEsjNnfi
tjA+QTKGf9feab0IDBZw8b3NfowFZwz0abKerpKfwW2YGcH9M0V+bNGdQ/nOT0gt
4OKVza9XCmF8HCV6U4YLy1J1WpUam3mE4DkorhOir9aTfvPq4CbWj3FDW70aJx44
fyg/WEAMLl20fdIWYWwTRN55JyeplLDfEefwZx/cxaCl1vbly5IBikUGAnKoBL1U
ZDpKACZvC9kVoFm0UWaG2k7js/v+JkbaMFI9DycHC1f5Mhu3H2PZsBizA0odT4UC
dccBOjI0QirPIbwxZJUkGOhVjjMK+B7fbczz2M1Hti5nHh+A5kyT738fj6i0OfCY
M4DTXsyA0jBLaF3c0Ak04DdysuLKWvglXDcdxpngtfdUKWQuCyA37TMAoHaJAicG
wLj3o1Vp/VWOq8yFwCXYyy73UEyQupXM0LpbfN0bySOU7J1Wcevz7kDV9f1U/WOB
vgH0ZWA8sXI1TKwrOLH+tyewa/826cZBi5pFRWKqzPIbS2HdliIo3QtRbI7fu4M7
GjwwIQNg2+7MUw+xTFQmR//sIyJTho1/DyEaRPjGrq/MBnu+8rpoEOcQbvJP5sZG
RV3w04XnftLc/lrPhXD5E5I6RbPcvZqPjFwtdc8M9h1wt2zLx98aJrOiHgIIy3rZ
WUhYmVqNEAfmuX9HUMatr0eoxAESIImj02aKduWq3iBkbSK9w3dvtockSdoAAvB9
AJqYwCkrpArRw3EUhNi8NSfYGaEioN+BQxkGsnhGmjxqX1EuPbDv+OIRBPLQS/uw
/xRaj0Dj1TnatcTfMzZufO2XCwLt9Z+96bmN5MS4JhvGX6uzYKQtSiBAMUmSvlaj
remcxim+R9SrzQUvV6QPmIokIw6/Id9HKqGDD4wnhzfz+9DfaPGraPrxPT5j4b66
MDt3j/L8xWz8n6PWtqnV8ozPGZ/qoB/sl/gDI2nQtn6MFzMHDMW3JGkp/KBFsW43
0qdIIl4KydmAhB/88JMOX1OVVjcE3nViyDsi/CYieV+EOo/PPULz/wl7WF2k1ZJy
LaHXKY0Yh2IZdMmEB4S9YljVPl2NX3JStlFU2bRUSlZ4hISDqcDkhF23nQc1SqnZ
W/QEY3L3HJ+zAwNeNJwZySDx1LlHnDGE7uwfKLHYTj/tzwT8GQulq2EYMYV+O6Rr
7ZUm5RggUXFNAZcq8p9XktwFSvt+PoXfBXZM8oplayWjsCcCLX3GCdiGLeBWJ+bl
qZJPcgvlFPDHjSVaLwU/tP/bk0no2AT+LKszvLvTLB8gOFv8TI9e9YLmrUZlBw3n
5DLIEY/e9wiUcgonukQADKWu4m3aVHUNHA88JMTMCsAW9sqyfXmpl4yp+dhUv3bH
hHvovzu3VnqNEYkQEfDgZA==
`protect END_PROTECTED
