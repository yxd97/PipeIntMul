`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
05dGSd3uukouk6n7yXaARfB0TWbtQj7tViss0b3XNPAXgGhs/lxnO0xNL/1c8biu
LwhBlO6fSubf5U1U4VUCrBtA+FJ04Mw14lx1iubxILT+hK4x0wZCGXdni9Y3hIj7
dObKTn9MQ+KsV2Pw/AWi0OQeAIVupZYUFdvqRLH2CDJLSgJTaRGz+o2v+jcvWNxA
KjUeG+vJsRUghnUbYWjhQOZ0YJv5JixxSnbshN6G2q5xa1bJaxXEqnZSTXCSMLhF
lX5/8E0zYXLLsuwFBMYDZLi02b/W5WfFCerO1ma6AYx5tIO8eYzNKHivQ+frDir6
HfPly1O39ZvsL0098nZetflqDqzyZYX1gfsmIa6enfptHLNRJqjFcGI0zGT+Alj5
MQkKnCom4+RfnrPyd2121LQOsW2t1m4VX4x4rnZAA3f0047hhXmp253jKqug+qBX
jQF8ZHvouMbYcwnUKtuIQmgBovUfWy5YkFmLW4Jqk9F4gdCbM/dfEUTNikV6uVMs
VhrTAbNUTeCVXYonTVm9XMlVJGdDedFxYrAAKNK9AK+0v2FChyj0TvyZx2/PysUn
07O5URiynwNPOzo2rxPCSGTsY3uhVPl9DeJ29ggsuagjNXj1ENXs+dpKKmRzW1m4
wq6+tUasl6US8CLk5FCcNj1MZNaovoLw08aT6gmDF9ayprUpiYINiWhuhoQDsjdI
UDzyYaTDZz9Xl8cO+FvX+ObIRIaofqchWZUK0uhO/i7LBDXaIhi0sJTkG9RdtFF7
f8svu/YcGw7H5RZ7SOJxH0B4V+/AKLbpPFZFtoBE0N2Gdj70Ne+M+I39u/G3MWxc
X+IfkzQIPolhO7EfEkgywpbsZYxPtYPPvMA2dJOKsc/BW11mJyE79XuIEh9ppqVz
yR/bDqI4uRmDI0zf5tHLMLI6XzSPP6BX4OYqfBOxiENV7jc3e09b75+NeFltwEwb
jpfzf8aa5hj/paTu4jjbxE9L6OibB5+Lqc8HO1WStc7fPQekHYK7S7YcHfs6NBMl
9B2pFK/eA6ux2fdu6lO5YwJc0mQrkSNskndwcE7OkXiP+JQJMEVrQINSgfkG3Vco
iGB29qrongCdiXcuGmaL+w==
`protect END_PROTECTED
