`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9IGDd6w9IC+DBakLCowQu8529eWx9hmF74PzKvy4f1Xh2AVNIOQ3hqpXl+HNxOZy
WUf/QMqOkhL2aOVs8yadWgP5XzxjgmSXroV93uBp6AJPkY7d50XASJeOf66hW8EP
mzwL8/okQXUq/UVkkenyGBlN2jeRTw0jsTwSFAsE/149AGz1wUc8+NMyNWkVIVXT
hORTbmH7njpgbs0xY4DtoEfBXrQFzGuGsBY0c8PcZoGbiHthYRHo96KOsE8MHVpJ
uXnRkJk7y3G0vdpEf/mWL5AhQeoNEcCl1E9MHsedO8uc7HcCU75X86YfTmSOgWXG
mbVms4vSZEc7kmTPe5zWvr5ifO0G/fZvJ4Ae2XMA2TWylhA1iYXst+ttgh8vl85x
`protect END_PROTECTED
