`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHOoRGwGX141p6rWzX+bMKyDTJapbYZByiDiS0CUrFOS+kb/DgcjOjWkHziwcka8
qI5v3vql3ik2I/M8PefAMxTEaRLp+ryV4/EBrwWgoWqRLTMn8Dkuhkddk20/geGW
837SKx1DHWrt4xfGvcWERbS7PFM00He5GpMsE9INQ7PrLxqe1kZYNMEAKoGoi+CX
3WRXV9S1zN4DqoqSWIqhSUyHnMTDAHM/bek3dEImfvIQAGyD2M5wWX8u78cbd4gB
9qmJvKTqIckkFWbuAd3aTaHuScduAX7N/Eh54ZU/wcf8Gdb5b5562yu+Wn6p9KAq
PH7vrewaoK+0btUgFTmabEMdqc5yzkVS7Hzfsr/8hlzlSx0V7wwcj/AWqXahGz0p
1hsPuryz3s1px7KxLfp6EJoqkUd/5Yfoa/7kHRXoK73gO6kZqpnvWjEEdhdlTWXC
`protect END_PROTECTED
