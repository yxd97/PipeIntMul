`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4R2Lm49pNUZrhZc0c2gne5whziylak2gCJskw08i5vo4ZU41nn4AkB+LN9WTvJ/o
nmHyHotdcnCP+0/zjJ318tCmSzlDvePrKRhzufuL2shVwfzqfElfC4SHnnIjNs+m
ZRzC6+2qkQB99q975g2rpjLBsRMdlA6LP/8k/mNUo9c8MP8QNzPHtY546n44fUZC
Ia7acpRkEXNp2HrYk6zSMLbnKpZGuv5NJLilm9vRp1DlwN00j3cM6AEFVpn4bNAA
AN91vnymUMsAuRK5IjHXyHCovXuiOtU/UiQa8ACey08zewl2Zc5AKsXxfi0e60WR
xn+/k4NzOkYNNrfahTCgzrbYAZr+rjdpZqkFD1C/Ah4Z5hs5LGkXuPRhxhof7exf
WpJ6dHQDHhf3GDyORqjxXsrV5OVtc4l9EfMvVBd0diLwCUuUYsEV/rODP2Vs6IoU
0a2af+5w+W+nTVNBrPDxH9MCfjL8hKkwTFfSW7RWMj0NuSdVoTvw7o3sFbDV27wV
7BqZCP9moJgRP91QZo9xQfML2TPHItOJt2peJaI+FFI4V1INGFRgTJ09Bagknm0A
PirZy3Ne+qhYZx/1/kUypx3E2RyhVyROLbSK+aimIn0C7No6j5xFHSvTsLchSIOQ
Qyq3nlnXii5oRWkAzraeb6RVUzz4z5MKaPl40I9lQcLtysvZFl59Pco3i2zSzbBD
Ye768WwOhD1o4hBrevX4Z/ZR1nzJqv/ORUq3G4KxQV/AxAcUSsWil92ybofO2wMT
jEVE7hA7wO8qgSl13By/zhISLiauv2/eyjeJA6cRq4CMpgl+Pp4CWCUUbeQstzz6
w1O3WqPndOyNYUBTODdGolGP5SITcyRcAHk1RwCUwDPKCghRWF714c3Bvvlo5Dbz
JVw+0RQKDGT2EnUxVhF2KTDtbjV2Fc39SUqQju8x8A2eP+LqYylXRi9qEwkZcz9Z
lPnbn1kWvBnKOgzzOsQzJFvf2Ds3/negMWl9rwyntYyqEBEW0hh18i/Jp02XGW8m
ftW9u4mKANpWbH5G3AMBamDx67IHUO7/jhQf+XTXMW3yJ0M0tGKVFVFq32+vMBQx
EjjyXPvcQowJa1d1phDe7pvQWftZ9aovIBd9/Wx9YNWP4bPOyW4YYqaszbSyaCU7
8YQ0W5O+3ngkLIAi/cu50tMK/HoXotV/NC1XMHTVhq0OvOG0kUj4nQhwecPWWiPZ
EFkuFEqvRUdAIhXVCzzuYPikvPfB7ANWefrLsyarg6MEUzSSYEMTIPL0ahCm1RW2
1NMHphXNAkvim4udtSQAyPr5Udsqx+ZhH7o/5z/mluBP5Tty40CurBPV7BtCHWfu
mX1QBhj4B3ISpfwyXcSCuIBaP8DyIblqmES49L2bSIepD2kFRyyG/dwvflOMyMjp
sCdoaYxiK6EabvE/KRx0FJbaypKQ4MzJj4ZkPPHOIiWNQNnaJdSPp95mlsFHJhOR
05eSgChGvjXpsBW2JfvP3FCRdj04OErZfHSbv5E7fn55F+KvYX6dJVeuDZp957mg
DrwbJ1jBXBR55JHwlR2aXY3cHClUVTjoKfxWLKiY3HIfH0rgBfUZID1oFhD7qRa8
XZL+gfaejkDOgnjFuSUHVAs+THwuKAPgg6hFn0iEOHyROae0zc8kLIwjiJbuQEKv
D8X74dD4whhyRd+EaEqpnGRkLxp2tfUIPlQrzzW2ri28ghL4zeQiAQKf0uM15tE0
awClYTCwuXHq+eY+CHUgbku3OjmjRHHOVPyH0WP9AycIM/C2M57eeZB7VRmBZk4n
rCge1k2PpXAkIVji33j9gJItWmIx8ZQKp7jR6HRK1uAGnscR3s5gKmJVsX1hQCcA
YYOiFY62WTs20jyv81qfijObMF3+nggVkup43ASmkMdR/d1ESHt0dtIxyIifd2kL
iB5LbPgXZDdfPPFHCG830kpPbmYFw0+CJkZYdEQSLX3EKhER2qmf5bMc/okOnlzc
h3VfNu0biPyNR+U+WscVXzKZXnImvZewGBDN5O0EXFrX8L4GJ6R6yCKs1+7cfrjo
xqtFLezyvPROO/NvHRQFXDFFzN4bHy+DwjJ6IF4dlaYgB1cPiiRP86N1RphnOdbX
H9Rjj6kuxax/KaIg/M5kzy0Tpp5sOSbLip5r2slu2Ti30O80ygbRS6yvOlGbdNcE
fgDN172twR2BZBDukKPfBopnJmCtRrgTdxN0LQqMP4r6k5LeiZgAA9A5xPqMJ1Ey
oCJNZJ9IOkTyPb6m27zVsfpcxbnWtFCG7xGxQK/chR4CFuJnk/XHtZgArv61HDcx
WRkzSEQf0+o5nNKumVNUlHK2RBpWBn3HDXTDhnPtenU/eHeliki5rNWbBmizWtd0
SAqwdVC6hN1HZwosUL1HEIGYmTpqEBQV+vJd4kcrLIXIothhWLvwpDGmkgoPx9dK
ldxuBcwJ8QfCVkgR7n3yQVaZ3CxYtu4DfhbUqYXYXh3MjxK5RN4haj527xgHRfxS
aTVo7DG6RhsHI5qrtFNmwnueepV+cCrRN6e8LMtmQhWvI3j/JsYxVMVk+fkFdfiv
oo/e2k71yNMYGnSc6NHh/CFaNyJncRmGkWSLN012jgUMX5RHXEWSWGTxMX4R6j/F
Ci24kV07SRqtKDWjYljWHLer0RHBsexaCWxGWneAAeZt8n1BixWKQVldpvbCwwi/
YYnga6wQE2XOzNw/yA1KzTyCwRJkzeHSaqZh1xTv8vjh8l4jO2yriumyFVsH29Dz
rJyYbKxq2djmMmmQeJ0l/nZ9GjowGElVhcHTnFnjauQsf4NNihwoAeov51PS/1kH
CdXTy4tSa+ugNzwwcpotqnLm+FYs0ljt8bTRMCcxbDVI8CDhS6PtcxvP5ebGkADw
SNgpHir2b67ufkKbc8nqH3igHucr56MW1BjRDy3GDMSFNVyzShyn1/YqMhsCgnLu
z9Xlt3nRy4wI/vSP3eg1Cjy13aXgGVbncHmO/ioS/SvWPKAPpCANvsXOKT2sNVrJ
/OVG7vZZm+2ojB+5WoW13G1tfukAowDmAXmsWlUy7tYD3kC72FTIXFudkfn7mg4y
KiKbfeRcAbWUKQ+81mxoQ8HYk0gUr3fbBwDuvddE/Z5whYEA7Yl88uVsOgGLsvuH
uxwU7mUDJaS2brScZfMqddvkt94D0BelcB3l6RZewGjntz2Lpeh9Q/G7XSFCH66k
mN4czym7oFsZF0X4ZGYM5ZAHVmq93JKM98xkzkQhOeXAHMgQFpw/Df6UOhu969s6
4ZCw5UJWELfV6BvW6/653ElSVdtX/TyKyQS2qrv2t/zwBcgrNiR2aPk1xdLkdCva
dhos7YW2YVEJJhAbAryvdDt81l+mMRmHVimUnh/POV6bq4a92S6+GZNxUrUoMnVs
Kmb3B7mW3xCucP41KGPwUHW8L/o+BM6XbGQLTRpKE29BfJYgifE+4wXj4FrsQfHV
mgEUDtp9e7mp4jt0gGw3myy0aEY3QAMEJlLRWwRHg+3PbbbaqrZK4a6vix6WHuH2
TAMUR7blnwwznJY6OQJMFhxgl0PWr0HalXzLJzMycS3rnnTFG4qDnXA0hjsGMZA4
L3UJkW7KyKv/s4t5AkYi1muJ09deQJKkoA7+JVsMq0xuXmg3MS4C0uhWFtaX1EKw
2cRduMp2glp00l2vusXMY+2FTuQlXPOR/tZFDIVCdfPiOvbJhpLzODv2JsVGsScC
Uhz7q+BrXWP4yFQI6+tPczO/jmNEZSZLu4OnkW9rNwRd58G6H1YudGKqQS12dydv
s/K2H+lEu9OpqW9iPW8ZR13k6C4vzRLE4gi0RVjoUsalY6wc8XpZE00G9ZcgCFVA
cx0zQ3gR9G3Wow3wz7nspA==
`protect END_PROTECTED
