`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJsahBYUo1VOLtizP+RIILhUgDJAIAypBxy8PZu4n86ooh0sjz2TxSruBJpZQgW9
vC4OtiSWMO4aCYUPvtZ1lj2m8UrPnggf1Z2Kl5tMvN1G4EuiYCzYj+zS2BMo2oRG
p9METMLTxdOktmBImcOKS+eBQ75mpwosmAptu/kBIXI3bjoTx082cDDmv/INt6s5
rwocSxlz1+TZpnwVyGaOe0GzNZE8Z9CJTnHQLSY4f2oS5H8otdowV6glKh8s6OtD
abpi4C95B7YYr5jfhxjDecqTWzgeKxcvEBz4+RqBS9is1qBx6KZ2KkY5tFj7boRj
49/zMp/GMp4alZqVnUL3KEMMcWgrYGPYnDfL0nMi1fbgl+sMUvvQIB69YJfJKidV
LGSLqeW4mX5pQBmkPQYMQrY2EGxy0qqBih3y4Rf72+K08lavnk45NJxkHOvSQj2d
EkcYEmPg0v6JTAhuZQfdDbm+t8quoGsSmGyPB4d56cot+G7PywD325SBEaAOOiqF
xOGjmIJtoBcUo+aNjlydF/0Yhatsr/oCCY8sDJ23/0p+M0Wwklo5yX01tC7Bw75l
+6iYwkXkAeiFicXBhLlwuuKldRJM6wQdRaAXpqmC1DLUD4Tibjyagwb+rKB8xmxZ
NEIFD0w1OXU3bg0kC8k57VdKsUemyuG+WSmk/lNEf7/ugI0zjvWpadXxYcsx45xK
XQS5VMB+Oiargw63+7GvLyHd9ryg657E6aetGbA46MbHz/JFmJboKImZssKQWjze
dIMwzvPF4eEhD15nZj7vZ5Ldi5bWoI7Vs/ALnAcPx47z51UOjALszgTUUxWa+Gqo
wHosh/g9KUzPoJ3/UqRvxq6YeULTsm5NLi+8W3LVXBDKGZtxXdRJDf2TnYt1ID1k
hx8BRNo1JxGs0Xd9LsbRLOyp+Xbb8aoS7MNIOvPgCBn2Bkxl3tionwNxuVgzcT0J
kV6s9GRDQxsBuWXzJJz1Ij5G3t73OWrXKShvzJj6pLz706lFkz6Uy5fhXzEU+piA
vjze1E/jXJ1tuqxNe5r328fSdXTdQEbZfcXv5cAr4Qq6g6Xv0g+4Jffo8Gfx3Xos
mIHYLJ6Q2AlRU8RmPBUh9OnCDUqGARTrMcSTx7MMIz4ZnHrbNzCx+nGvQXIBEJ3z
QWDc3jNNsKdekQ6EziILO0MultY9ML1L0a3h2NML0o/QdqNwnjM6vztSfCw8cLFp
QLIIlSHPYtnG9UiaS59VUPq0bRYZBIHRqyUGADumvXNEq0BQ11PoYmYBA3h2P2bt
k8TUAI9xaFEo0TNaxtc3LebHKPoD4Os6G1wnVbePF3coGAkfvm/B9cJomtPd1mG5
2OzZ9tfJx9VCKmZBfb8NxbC88iC8zx18vvJkeQhUn3A/71wEmwUJ1WdHZva1FRMf
wyyHBg0nrIv3Z9Hf2r39ehTxXJDmQfrdbV5clYTgNnf6o9VJp9UT5Qn/vyW+6X75
f69e0lpYr6sXl/EaWByHY0c4/J0X1eyr6ZK76BWsxl9mMgfSMkbjlrrkDnx2R8nm
8YARlwxjLUJMFvhvPYboNKzVLZVL+QhBLyYSU16umQruuIhmMhDBGHftSx1UOizB
dOJg3+ZkbsWA4dd1Y/PUffSGBFe5SEsz32u2SUaFkVf5UqxFj7c/NfBAFOEL009b
Yv+rREY/01gQ7od5V5r65CCZxxN3yHlLqS+mTHSlUM/BgEUoM4y9mdt0m4sh4mKP
GDykSLc45sMPWg8F2h0CpbshiGaL30fNtUB58Gr/pAbHaDTk4T+VQo1bUUdmqqa6
8Q2SDob64fHnbRZ21taJPGUxMJvXp5zasQN2pobkSaacIRxqa0H5LI1Gsl9DHnF/
/z4gjoVmCGHNvz3bB0TPc25hNQlzTtNS0w5HSYMz14GyZ/ZCIsTBGRuR4N7Ms/JO
JIhMWci6leEoCulZYHFPlX9QiFotzjQCrFN6j/2zPc+sDUvmk6uB39rXcZRLirOo
48KS02z19XZuX+4mUsiE7g1xlyryeI59FmijYO1g8ex5EvYxdyXqReVaKNucXro2
t4gBmzTvm9Nzau8MsE0+cRu7K5lXn8eTeRIVyqRIgg/0JCbmbCLuBTJ7GvH2RKFa
BScBC9I6jSPT4qfA0pI78VDsFkIBpYUVGEwCpoei6ahlihcjewELFbK6Sjmd56mc
6AnauzStR8ZWZ3HPAt/Ql62M3AE8CIFmCaPZc0yn4H4WY/QvGFWCafO7aQPqDGFd
WH2SUuPQGrvBRdgmjGJ2gG0kvdWZNp/kqZfikxBsI3m+OtLMvTOq6g70knlrFepF
Tkj5EL7uiD9rTp86s1tIjg3rpxGM0G3vaGU5vgTtsSYMkIa1NIi+gvp5rIIVvCeN
PBTbqrmDbE+LUNCT0YrvsKyaoMkQlmetpdt9kYATuVrvByfMpOYmi8bbDXqW+IiA
DAskw553kuiseMYP7KQzxSZe+sE3JOaLKbkewtyCfN909sClRSOm/YQ25XLCmLrI
kHQfIOxMvsP13Uq0NbFVW/wBcuC+4Kde9xoZrbYYej9G21CNAWQY4MD+7FGHtRJs
T/u4qEcnuhx2Og8IOVsmWz4Exmg/jVHqia1PIRAOtt90qkw3kxt5C8+sCbEQYOMz
vpTu/DxQltoEoVuSh6/mSBKG+dJ4NHNVpIZJ4DzFDRc=
`protect END_PROTECTED
