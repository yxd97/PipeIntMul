`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAtqLzpIyrPJWA+8gaTSFHNjEVif6TY5jvN+8W5tmv4d2qZq24IjspsuJJmfsd/8
eaz8j00UqOFkUef+q7YkhTvNbTz9JOHztOt70ORuBbLQUWSPOjsNCAwB5qjdgPZC
dRJlwDsyb/i5imxoamEB8iRXrZPgGVLTn8ZphK41Sz5GBDs8VXP3t456mVbOK4q7
wy+Tc9yHaGa45CL9jViKe3+coOfgvmKMxndkQOFXRO/viVNL5O2FFs+SvMK9iI+I
nBtSFS21vROHJ4wV8I36Og==
`protect END_PROTECTED
