`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kupj54XONG8FrUXmlKtivYHU9vwVjrYnlS30lAPPP8bPjBSF8ZCiLPjzWgnyWvmn
FWmjP8lv7aL3baYbLnELy+20WXM5YeUL9SsjuRm4v+HIgatvMFF5A7GnkOSG8E2K
ZObtCjDjwP4IjIpJM9WR6ceO5HoB5nBWqxTPvedayzv0psGuyM6R5epo0E5Rvq+i
nd3IrIVjUk6pdVYGmwddLtuVmeHoA8cnuvGqaEzWNFfbTE8GvBvZILHUmxF2pBos
rgvPkN7Xoe+tNAaEKVfSV01fZZxDRzQzvB8r60TVRMys1fG53DCiLqoE/HhPnFoU
iuLevQ1q92+FHCyl6LtrNg85I0E0+mMI643+GmNH6XUN9Iw7cH5M8ALgYtUlg1g2
r3Jmdj5uQfgdpMPUYt9wXjtDcAB3iNagWuxjng1q43fzSUQhpUhDbqwnj3qrP8ag
O03Fn8/jAApxyokNanbOjvccOkY0OnXN2l2XNEjGpMIN6KjvI6iICztq+FMbl6+d
UAu42lDv+mU6naUhSJJX5xOKDuGJVQaKrfl6Jb+fdc0PFetrUAL8wP86a3B3j8TB
R1VG+eOAViqIm90waD7MVFyA3t80Hx6T9vesDTJQLozLRIzA2yHL0/Dsaap65qLs
XMZODEMRsZMtwApu9pMIdOKKxDehu8YssHyUAzSRH4TN626qqmCOXNa8fvUbkBDw
jlUNWt2u8ptRKr2J4lAY4uO4uK3HKBQfNVtFGCdgmN0U1mFNso/Yt03Vl3kMJWOq
k6hCoUqq1Jt9zyszrSOEHaxjTZo9pmD8H4CSWem5gk6XnOU8ThXFJKMGe9c53LdK
EMDePWDgS/3+9MOFgG3ICcTLqR59z0dvsnmOyKHQTdgV9FuEgD6ADVGx+5vs5ofU
FtD2S5YteGY2K3YozuKYQzZrlJJw/V6bLx/4Q7c8VfrI1ZtUmh9JruarjoITembN
TpV2WiJyCjwA1NpHHIvFGRqoC2l1zPUZjJfrMWrPGCCTyu83Xkx2AI7c93zluQBY
4Eug1kmmR7bUWrXfEFeLoEDqgzZrcv8aPEVAUJMbTb/9XjHsq5zD4ZCawvW6F8pW
MJymvSj4F4H4GBX9sIID9hbdsu4hmEvNjxpFh99EMFTpj0FvNc8R73p/Y3/yScAn
3BnpAIK6MI6XpvKvnXhUzZtdOLo152o17ap4NRI8n+U9NXKU3oNIy4dt9qBj4U49
aKKI2GM1UaAI9sB8Vt1tG4zautwG9UnAeQso5TFgIQRPMmQZ/EV8y8vVdqcLfHQ4
HO2iofEpAOWQfnIkXkV1qe8RFMWCRueyCpkCsVwdWfeqJ6zzQmgKzl1mQOq15dKV
9kpnumGfOwfC2Vz/Jks20/IPK6CopAG0yl/ceGgYVqYlvSBs9HtI91b71aqdosrj
uK23pjmO2p22HY117np+6/Ax+FN0c5eXytqYSzqCDFl65RrF3dScw5tMVRzpuohn
Oq7gpJS5ybrh26EIy3+WNh2NM1NO4IuqRHiiisrQvc4YIcGSKFnaDPR85q1fpW6C
+wX/P6DGgLs/8Qpvw0gZv4vRrXDESjJ3lmx5Wt9WjlxTmhCRNRd184qbKKvWlipa
TiZWN92rZDYYtISJQLcL5GlaRN6c8TVO349U2To/F8xZBaYuA+Ih1L9IrbWcE0JR
R8/dEgDSX+XzOzGEWp2D39uW4Wz2jD13kEqTJgd5ne5B4I00OarRivLdL91gb3m/
oTpgLyX6bbpxoupQam7DlKoS9EOsBgjD5GlfY4Pug6k1T1iWWJFVYP76FUCpjfCP
GC95omfEZn9H5V6AqDquT+Vfb4FX+l4cVatVXdXj2aobl/9pX1creArcd5YUaEGr
NnBYcbf5ADBZhjfOsXli5/02Ku4USZ7dEt2r3du4FUGr6mqsYu3+S5nsvGmCT5O7
+K6TViLPGX2JHppKdQjktVvz2NW2PEYuGVun+rKr/xBseYUFGpC1V4NCsZagFDGb
FZS5TN811GVclYoyoMC29XwsfOuKb9hBXqr4ByKQyumEEXuveVKOuYsfEHa6k5c4
kVbB2XIT6Fpsa/lK2MTKl8imvsPRWtTfvda3e9CqEbVxeQDg7KfrTJ4xzoq9l0d5
jpiqBWxVGnG0+QOozL1MqNlQEdWkmbmCLhSo1vp8dSM7o7r1SVGlmNBHkUha0eRB
dP4kt9vPMXK5/eH6rW9RmFBGNycPrUKsgw2IMRELTiuYCwe5R+Prl0NqWijFHmV1
dXa1BykiBaLIR3imrIkXH0YWj92DJW5kH8+q0DAQLyGgpluQeN1dZ1MrK62krfhY
JX/Sv2X3BkHRq/bNcjVvzjGJNyLDTzWiLC6nVt4pF3e5Fqhdl0OQGhAcNaIBYgDZ
/F/ksBNhAEeB/FSo2ASG3wpnYGu/2H1bRxDTQfIB74z2+akHv+4eFpNiMOReh4CY
EF+z+L1amJDLZZJqNAU6huLtxUhlMyJqR3QLfK9qnHupMnaiuQw5hmFeW/6rfDUZ
CQY+3plGINLC/A239DcsOqLDK6l4YEmNzcgNNi9EaheeCEyvr7T6KMHzgCiihGuk
ENAVMICkfyFTHQu7Lh3K4A==
`protect END_PROTECTED
