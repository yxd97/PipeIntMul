`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oT2SR86ULLvjVWIk3Wi7n9oB6ySAE2ILOxqs9iLZrhYi1ZwmvzBW34cuVi7ozdq/
I0TDf9NW6R963L6mCwz2bDGEdr9NTmRE4fnD0d+KH/RxHoIly9sHWx0wAmHibIvB
//lsRhengD7QJWYzSv/a3pOjoeCySvtdI6nHkkA4n8nuMAkSY9WEPrDvbslnam2D
aNcGcLDJBcvgfLfkbBNXLwBa3eVshtfMrURtGWZcb0zr2cbAnrn0Up7JbrEYZNtN
3PXGkvjz66P2W4anAyQY5xQlIv8EQ0/1q63KntLGvQAYrTcuR9dRCveK9pe8BWby
LIiN5VrKM8Zeafi2P7GWaEmiyV13bakqAU255ZxMj3HOMLUbmVHR/0OMK4kHx0UC
dbFyPoW1kWcLOmCR6iPPVFpc8OBbr3ojUpOlhpgoBn0cCVhrLcsv3xPH3wveScQl
MWqbOWma1hC6QzDrTHthSNakU4wyku5L/MgxoIyQvtc=
`protect END_PROTECTED
