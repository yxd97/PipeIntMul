`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qbnNBaxhaGd5mR6w7Sqvupj34e8da7jc06qfRjBzdJ+qb19HEf9asOtUHWYzvpXh
5eTZEjqy2vNujapdTYvno6TxfhF5/CIiP7Xx92ABUtV40lVaBV3LXJjkEYp3gqAo
1yY1JTODHfcKr7qrN7a7+Sy4eHwJb5+G0tljHM4dWtUEDbL+W3m331coKOJiy1ij
w0RDac5Hea3b7d+EtbV0Hd0E75KoRoTCvu6w9zCMb9JWTAXS1FCh7WvRJPkvfKuP
EW52p2CfWargU18877s/024aUrDlqVieu8jMwHCKBvZVmOKsXjVwQk4v9ZMpEuLL
rXEgXIPpaqkJWg9eOZb6kUP1nvdyTYNb6/LpNd+ayx0OA9a9BTErhnWiSa0ugtQO
Ip5H2jcg/ssNu9F+mhbLwmIKhZtO5qJzMiK+Issr63q1DDvnLqp+PiCI/w5Kgo7Y
ocpGUK5HBeRsLFDPaYSq2THzDRCctsPlqjSPkoNmacSWkZmDXPdJh9JKVMlOGfe+
RlEjJb3IWvS3mwyqErRt9Fyp9bKqbBDS3t25dpgtR7i7T/58QCw2NNUypB8+6yjz
y+JPw3pZ68hjn4Od/pSHVq110nnGlnuYqnHkon9KFNeuQvBlQwnFPKJZzudXuMFy
4hJHz+/euUO+s2a6QVWtxGGAZmDzLn0goKqvHGOUjjQQVfudHaMcn20TcJWObHaN
GnGTctiBob9/pI2wc8mzP7xXA3hhw3E3+qkAtPAKvGo6ACpmbAVgM1vs3AcfT1gu
CL7mwjr2sR9cQgNZ828NFsIcKTwTqQvwVUef7J//9dGMkAOZZ/MZFh+HURSvAUH2
aSE9+p2YjM/+47rPN6KagGmPR6lyS2EP+zdrDnsHzKrnfHSv0rO53M31YxEITvka
sSOQFxbRrd5ChigL6sIwRihQT+WJupa3MPkMHkeiBDQH/lCx8QwRYomZKB5A7Chl
`protect END_PROTECTED
