`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CmNbXORC9H7ThyNPE4kXATSZuQLGIkDod0EdzsjMI3mOdSlHbXggVG5DSuqABWWL
o6/CD8zXt31V06bOe5jzx94HwvOGXY5sv7pcnJrlHpDt7+NWR5uWUTvIUhhzfi7F
+FV3wlyPyCF6aRZspWDOFtrrXlHWsXoZ3RxjaW3q7pPj9Rdccxs5hrq/nzjhUCKg
pcbeYdphOZj6zDvhelbYUSQxi6AM2tWoH4juWBwOada+B0WRzDcWO9yjCeHXocKX
1i+XROXtL+vO6OGUFo7fKK20ptAEcNZzj2SLmv71xu9IS1fRkTu23tprh8AoG9Vy
jnHpUCPQu/k8otAgXWlxjfFKZjJPxwmq8uKcoPvydTl846UepLsQacbAorBwTXlc
MqQVCpVaUvX3RCCB0PR+dH4PbgCgxoLVq0p+TJxSgC/tTZILB1gw5XLYIri1nkpF
`protect END_PROTECTED
