`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHLEe9Fx9hDDIBuLrtq9Autlw1EkgEI28BeLo2ywTSYJH1fv+7b2QcopC9fJv8MI
72pVuvXR5E9oR64xfrdFFtaGt8RD6Vx5rpRbYplD6pIISZyZOtpt77FTHmhTTs+T
4npJQ+sDa0lo2QXHb3gHFHzr3kTvbQr3MW3NAJ8c5eIxQgse94DoNJmfW1tJ1MpG
AElgLEAaOcA0+cfJ5EPLEFE0795lAL6kgUNgwGAxFIPcQGO6JxGOUrqlwx/RstIp
LaYlOJ1EUST0flJ87ireZFSz+hW3GTSDCqFu3GdBgtijK+VgtHiRtIuTUVpdrQC8
aAfgEBwPHHgfec4khywEYLn1M55Sgz3zwBQpoH48oDzT313nYpe8FlV+kwOi3zcf
kzxMoARqcb3kzCq9smpOOfb/d49eXhjdvNMiRjHYQqifVsDBx2RkorEX6WUgFY77
xY2TMWcmV5dOUpQGwXORwzG+4RcJstt7lsvTCt4KBhD/23TubK5wSSbYyDs+S62h
h8uSxhGeGNZUJJs6Lvet95ztBy0Mzy1WjotK9z049+pkaM/FRk2EFCI1tChGMsvC
`protect END_PROTECTED
