`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+XN7Fggt3KeShU0D5fExzoyrC9CTMOlOXm8rnMeXXlDr//JG31lc4CT4fTuzk1F
ec3u2Zf1uz6dmylpXWb9mUEZQBN/9nNcP1naUn/tvFTnaKHC9HTxF9r1iid23COG
PbU0dTKl8XdVcYqthRcUn7fAkNaqZu6v2uH5JMHPNZSC4M721dZRbpw/0E/e5yms
uTa5F86UjtuxV0GcYmGUb6Pqep/M/TnsJph2YhRfTLrIPETsboDRSCwx4tCr2kI1
tKOPl1QsZW0y4KpD1YXpKEo8DN6+R8EjaVjMQqmD/reJv9unqE+iLn8FpBomy4z9
4/tY5b5iv9JLnuz+IhtF5w==
`protect END_PROTECTED
