`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6E6ohAFPJCL8ZxJ/OdOOJGJ0U2U7sIR8fGNR0Cxg9xyraa3ow9SaR0KdRFrj47v
FmwqfkQdI0Nd7KGMVX+YS7/B5gmFP/F3alDFsMzK5iJtmV7cRy9mugk0s9C3Els1
NWTmg9xwSnS+2vBv3RRFQqSPizGr6+Zne9fpbuYkhJVh8EslDFjlnM5+p1fNNohQ
Vvdim8J1RQqj8vnJV3dD0DWm91ANTZQ+SrdIH9zJQ4DSYV6FRdde32aTq/CRe7fN
dFJBb456TZBwkxrzf8eY2rYyh+kt0IQM4hicC3o2zxszG+0WNy/BlfhbTcZHlQz9
SpDrKAlJWWHViqpbkRQi+5OPOoxv7mGYBuKmRHro2OT9y5qamBUdrLWZZ4jrqse1
iW4mxGOyitmU3Bux8Bwfa39fMGYAg7Mu1eaHoik7TKD75UG4kZP30FNsyXF1vyyX
l1nA/i4jlgwimpxBqFYN8SUYgHZ3qJTiJURz+2ZPRHxQhK/7q+nA469wZ6YshglM
TC8sJKG2GYcC0euXAnMDlK71JELJTKyqi5y1VyaizuM=
`protect END_PROTECTED
