library verilog;
use verilog.vl_types.all;
entity XADC is
    generic(
        INIT_40         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_41         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_42         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_43         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_44         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_45         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_46         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_47         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_48         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_49         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_4A         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_4B         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_4C         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_4D         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_4E         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_4F         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_50         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_51         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_52         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_53         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_54         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_55         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_56         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_57         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_58         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_59         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_5A         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_5B         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_5C         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_5D         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_5E         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_5F         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SIM_DEVICE      : string  := "7SERIES";
        SIM_MONITOR_FILE: string  := "design.txt"
    );
    port(
        ALM             : out    vl_logic_vector(7 downto 0);
        BUSY            : out    vl_logic;
        CHANNEL         : out    vl_logic_vector(4 downto 0);
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        EOC             : out    vl_logic;
        EOS             : out    vl_logic;
        JTAGBUSY        : out    vl_logic;
        JTAGLOCKED      : out    vl_logic;
        JTAGMODIFIED    : out    vl_logic;
        MUXADDR         : out    vl_logic_vector(4 downto 0);
        OT              : out    vl_logic;
        CONVST          : in     vl_logic;
        CONVSTCLK       : in     vl_logic;
        DADDR           : in     vl_logic_vector(6 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        RESET           : in     vl_logic;
        VAUXN           : in     vl_logic_vector(15 downto 0);
        VAUXP           : in     vl_logic_vector(15 downto 0);
        VN              : in     vl_logic;
        VP              : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of INIT_40 : constant is 2;
    attribute mti_svvh_generic_type of INIT_41 : constant is 2;
    attribute mti_svvh_generic_type of INIT_42 : constant is 2;
    attribute mti_svvh_generic_type of INIT_43 : constant is 2;
    attribute mti_svvh_generic_type of INIT_44 : constant is 2;
    attribute mti_svvh_generic_type of INIT_45 : constant is 2;
    attribute mti_svvh_generic_type of INIT_46 : constant is 2;
    attribute mti_svvh_generic_type of INIT_47 : constant is 2;
    attribute mti_svvh_generic_type of INIT_48 : constant is 2;
    attribute mti_svvh_generic_type of INIT_49 : constant is 2;
    attribute mti_svvh_generic_type of INIT_4A : constant is 2;
    attribute mti_svvh_generic_type of INIT_4B : constant is 2;
    attribute mti_svvh_generic_type of INIT_4C : constant is 2;
    attribute mti_svvh_generic_type of INIT_4D : constant is 2;
    attribute mti_svvh_generic_type of INIT_4E : constant is 2;
    attribute mti_svvh_generic_type of INIT_4F : constant is 2;
    attribute mti_svvh_generic_type of INIT_50 : constant is 2;
    attribute mti_svvh_generic_type of INIT_51 : constant is 2;
    attribute mti_svvh_generic_type of INIT_52 : constant is 2;
    attribute mti_svvh_generic_type of INIT_53 : constant is 2;
    attribute mti_svvh_generic_type of INIT_54 : constant is 2;
    attribute mti_svvh_generic_type of INIT_55 : constant is 2;
    attribute mti_svvh_generic_type of INIT_56 : constant is 2;
    attribute mti_svvh_generic_type of INIT_57 : constant is 2;
    attribute mti_svvh_generic_type of INIT_58 : constant is 2;
    attribute mti_svvh_generic_type of INIT_59 : constant is 2;
    attribute mti_svvh_generic_type of INIT_5A : constant is 2;
    attribute mti_svvh_generic_type of INIT_5B : constant is 2;
    attribute mti_svvh_generic_type of INIT_5C : constant is 2;
    attribute mti_svvh_generic_type of INIT_5D : constant is 2;
    attribute mti_svvh_generic_type of INIT_5E : constant is 2;
    attribute mti_svvh_generic_type of INIT_5F : constant is 2;
    attribute mti_svvh_generic_type of SIM_DEVICE : constant is 1;
    attribute mti_svvh_generic_type of SIM_MONITOR_FILE : constant is 1;
end XADC;
