`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dhrLEQrEgg3P5q8Pdnrd/ewgzpReJGNaCD49HAecdA/ozA959wtX5yuK8M7wbtfH
rfJQCzuS4IDeAOuTkli9mJJOI8IUinu90s9cXYAHhcsQUE4QwEqxXohjy5WwwTQJ
15cAvAZKCs+GA6/38t1yX4uJqJLq9QuKDnwoFwBgvXt5yb2Hb/spM/edD2RF2K23
6dnGUVsnU1PPkW+9jZGRV4sFLPwSJUp+iIsqY6g51VXyQtX+wUDBcnxUaxyTeYYr
Hl4a5GBa+fAkD/zG7Hj47Ns4a+CW2w4q4ZKdWA2a52aN0lmPr2FTFS0YxSsyjcTU
ODsa0aqRSwpo1Krdv/TWT5cwys+wiz8DNvyVTo4Z3Ayz1GVgmcnOoWxCewUilzJS
FtE3pFlIMXBx2zQLUIW6qx8RX3duasZi0KwUYiftEggYH7auqp9cjUUx8NhzObSM
qU3ljjsIC+K2CU6MUQqz4A==
`protect END_PROTECTED
