`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xIC1AOUefIVDmcRtvd57OidGXq4nVrwqPb903ga5u6WsSwm8Ly3hr0yNuGpkMkJe
GGT2v41pEDLPgA36SRSsKN9K68plBlqA3FZK+wOwOD+/UZIL38JpaF5ZaaTsurrN
MCStaiNzrkUntAL7+zpkRt18I0228NAPY7bTjMkSd5DTOxN5JhQs9zVVOpa+syZ8
RaQ1wTvlNUy8gWAZqX+SZxa7/6xAIGQNbqo50OMt9ZnvoHywao0KV/nml5VisQIk
VUIrnXd4ZyxnHRkw763fBhWzHvvHvmWr8emh1CDio3bbPcIzisUN3tq07MguTK50
xfdU9n+ySTbH0umqECiq4UGGumFb9DmriRu72FKSBA/6EIDMuZ8Ld8qJ8NLuJTN+
/v8eHdeZR96YW21IG8GiFl9sUDdblgwvuYqDsWMrIPofAzCdNYKG26xNqLjxPm0a
4N4/gXwmWilxHIReR569xklKx0TnCnPcIOk2eR0he4RO4cFaSorHV26qnGTOBTqm
b1QPXPMo5mIjxgUbO9w2QN80UEPyPTCuUACrJa8qqlT2UFZOCApzz4TIyTLLfc9P
5L/d6APLGIUMqDCAkWPwVI1EkVStnmmbyRk2HHf6Kz3/xcZGdh9Zl4h5/0TeCNDv
Vs5hdIvlx/atPULTcYkfuf8/rsdKqlf9v9B94KjjAnDxkwhFtZg/FUZ73I2FMmit
eQoSmHWX//7ndzr497PNOm8BeXhNFxyoOlywMpRfUnZWfJ4hXVHOHPMoQsVKY3dp
RhbQWc5FnBofsRHETbVNzfoi2NB1ks4UkNJuZp/4sUk2fJ9eJ+gGsF4nfO5uQVMY
92piCKqEVn4ppFK0o12nuw==
`protect END_PROTECTED
