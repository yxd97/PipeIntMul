`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+MmvrsIsQfJ7V0KW7Hpvq4jSKPM9Qe5nbmby0u0HUxM6EEIn23ZYeuj6SjWNXnZ
JAcd/r+b0qpCxSWMkvOcJx4IHXRO5x9CB/XBrxubDLZnM4/sHT9rD+R6j0dOtr2A
P64GLdztkpAFtsOmYFKI75+65VfZmME2slsOJu+U9BQo1dzqx6lZOttGTsJCebK5
uXesTp0li+TaeM0CbzCeA8uLj/Ag37oOFFM69zlRD33pwMgpdO/gIi7TVtbPCCjL
MNIouERlIVCc/fvXmp7kkWn/yPhG/LEhhSdchDKTfwMH14wPxdQRQMrds15tdCmj
zB/+uQduGBo/Ju7MPKwWJEoGlvDsGPqBlzOlGZipcibzrvD74/ysKjYqgDmUulAP
jwy/gp+Ii57wwZ5CWo8oPfRLo9uHE5/x1No9Ro8+tkix5jyRuZCtDLPC2Z/ODYiu
AMouWxGJohCuqQxX5FrPK/62tF/i3x7C1iN6V5Co5nJpbFJCvoi193YxJPtk9p83
bu6JMhzZDINywsg0ya812gHbEWaRnruClkjBnscInp2t/gbs9vfm+tReZzsBBWsZ
NQcvSMVv4Ubb1oaYePatkv6yFy6yLuAC+BvGyXFiyqrHg+PEva8dhJzkfjSiny6d
u9/aFI3UeyYkhCBYfC402PPxI4JdMbjKoYnKhgUAis9OvYehv2akIa3iWxAhGbs7
vziq3ZzB6GGUDEOERHcwhkM/yYHiTP7NVBd6R5tXHk736n+j08Iv2boOXqqbQJhX
PUR4obcK4xj5aswINAIkpBFh6tioDIRHlpwq0urxE7NluvlNsuTMN1bf/5b29YOr
4+917LDM0yp+EG7+/lIgmSLyJ2OyaL9g8u5Kw42Ndv+Iuzn0qO5WFVrPuAHDhYb0
sDiLde3aqjH2a7T4LgUACc8QOrnS5jn01e3fnvXzca3XVkEISGVpK0vpjTi+OTgK
hC/JuBJ/W1+6oVZr+UnhZAKJGL0aPe6BlMrifDaaSl1FKvOq6Rt+xPwc21HtnMcw
9N/Z2zd2+7yNse9BF6HohyVWAKxCc03tk9LT7THLn6PN34FB1daylFyTxAbmAuwV
27yoLMkvNebKPryUx3l8AXiPJfM6/SWsdYI8MQWaF4xZxGYRlx1J3ZRJLYWRp5l9
8z4gjYjQ0Aa0IftPmdk1Uw==
`protect END_PROTECTED
