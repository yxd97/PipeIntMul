`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QXmxEJflJMmMAMJDWfMvem7e1FTSJUF07382Gzwlq+jYfL/jaefszGTOH8HaxxtF
lSTNQt+0o31hNPNB7V/mea0KFX7SeV3GdutCXsf9D1BhiTjUohdCo72kMoZzrOYm
R0/R8dp9njq5wsAONHIvFNS0/CwIOWeS7pmZ7B/u8omeXgKT01RXW3Egsv+dtoes
rhGVjZkrdt+K0RflCkCqdkCtTlZHK+0lMNtSMHOuVKlSKLQ4QTWvLsmJpc15aZxR
zf6tnATPTgesN0ZHOJuNJ+m/23+sXCle8Z7FWTvXLsAoz/iJzpeymbxkY6aaPk3+
NlkW5Y2mSfbOWx9zdKlfKFNePFZWBtbKzvC9XmKxyAQkVUkj/OMXtHv2Lu7GznqJ
Ywyi+QWIeGFZ198G+p2Mey0IcjEvSXPRzBn8bQTTLNM77Z+n/yf55S9sFalFtDXp
mdjCiO8saZY+OduizMKtB2cr0MINSQ74CMEgXtvrQvOHpgC9fEJKZWgv06b4q39+
ku8CXSDX5xRDK97vR8iNz7QXn2CD0G4cux0vBCpSuKq8gqLkvEpAs3W46xxxVpsW
QkkZvpQD5Lg4Sci7NFRx0FyGUEsLRAHW0eUPDVNO8TLWN9M6lDbDUW1DcJbt2PXv
ktBzt8qBW8yaR/umUqBy5JfR/xBxUNhTSmoLWryDQzOAi8umqiV/ipjBsVtRgsEr
UA/bHhFHjLUef9t4VBx8WL3dmZQTULGJqUvva8pJvhv5t83tBN2xtjun1EaE+tVG
0n50GIU27dHDc7LzX6QTGDcH0TlPd18kwVk2c2eUFbYV7GbXVLzp/9QgParXzAyZ
F56nE3LnE0+OzXKLJEJlGpTqBNIbRX9qEm2tMDq/k8pBALIz+7Qe3jUc1ByKhzhX
jUesh19JYcFl/YytDBwseRAEreOeYFDkjWSb8ywKySfpbk5ahKljeeygtRbCuM+2
ydfAPflsyZ9NPu9AGW/kariv4dCFSRXEpHPfRP0UWtuAxIJSVWsSVgPslFOckfna
09908ZOeyd8q1yx86+BvEdkn/W7tcZNQS4pLWg9VDY0zb9PifUPEmIWfSMXMq+0K
mQfsLOky2+5W0HGiO3gylBhmTEAyRJYn3QKvViJxsUJt/FeFr2WeOomCJ743VPey
NTGKbebDJUMTzRbedaNbBBdHRAJBB/F3pdikGe+wfAO98X57VZLebU8U1PoKB+Z7
zCjhntROPRsukrqYF/UoHKUEJfG4aUDj2vcOEoCF2YR9ba4eicm9DVdqiTuIpwsz
hoVm1zVi3MmXGDqw7QKgFRyJfU+d/7EXKnqd6P5tREpoNljS2sFqUYboNKyDCuDs
VXKMY28fo0AfO4e7vrlwH7lFid0XY0g+7GJDfTCnvV2WNk3ZgAQnpxgfVeb/KVEd
ns+P6awm7EwXnU5U8bTevodKCK7xHV4Bb4j1SCMtZqyxSHCjqGw6LqbTrIzgBHWf
Yy9oWPl+CCUsOE05LLLDw9I9gKFStvUxXSh7nUyphAUr+IL2gmhWzN/9iLNM7kwb
ics+o8X+WiYqNvSqMKniacut798cCIMAjJgYDxb9EIa6nmgHrvUL/dJpYgv2cHh8
MeVzuhqA/CzJuxJGQj4eDRTMrIzgwf7d0f7jxR93MrvqAeTe+mxbt81fnhqF5YYn
MrhA51Zx0Zs7Fm/ZNdz7JFMNwE8qLSk/gfxsdWw0dwVP75ta0QwY/tt9Yq5UC78Y
mrgYdVW7Ra9a936crAwjO8XjrK18iOx9v7oF/nHWCufH/bKD2oQ+QoeTwRlXQ+6F
U4stnMfPUB3s5m2zIFLW/buS+o/aLvtvJ1B81YsK/9+fRCdpu7f284BCMB0HVc9g
/oy2kCqO0QmHO6fAZADhS40ee/sbji/mfPYtwQtwgKYXWcrfOTiM4WBC9Zqf9nDT
SxNcyL6ApbFGI6aDQNkKKjavwBgspTUBEsdM4LfVgfbRioLuyzxHq5gGteX/NlGO
Twur3/8lx3e1EJmbj3q/OA45ebdcEP9uwx3dpg1WC3AMDQSgNhB73W7cabDZIhuK
61JVFeBwr8QG8M/+j2sYISktiRJ09szzBwMMLb9tYHVp8mC8rlgQJ6050G+MSxXO
BnVqDMrvkVgIjEKV6PK1IHvL0yGOWB/iZG46V2jS7RNEsGVsO/x46KaST9RdmE2e
ccE2MVi7zFuK0V7j1ZfI0p8iRVKHXsmfbV2hTOjKi7XEcMd7RNEVsmXcfdBBF+SB
952Mee85KwUENlJqZLVHHVcoDintPxgAlgRpjeof6yTPdF51KIaK1BBVDuVg1Y32
djvcEVeBpoimAMDg2OFg/pkHcMIMSQHSu9izJPjdJzpk3qAK79/YgMCp+CwaIsDN
Ksyy9mqC+Wxg+vfTHmvMHounbHVvrNAOyupXYNhsjS3JYSjIAc+pcVMwKvjhTSbs
twVfBjwQIHiWIzfn0968Omm6r20ucirE+AvhzbC0DUdzgwvkxeXkiKDc/S6ikuVS
9oXk3eN7siDeiaJ4bfU7msMaG/eNgD9Nhw1h+3+AFoOIz7ULj/nFbRW5hp782ynU
pFgFHLeRArG5491Lbg1vcTBImgQA+UQDeSAnnE5bSxtcWE1RD44DUxFO1g3CvKZG
cM8w7tti/n2vJ7bsnW0PtIfYPkHRJIS5yTZiPBPoz1zt2NyNl8m/8VnvBLx0kK5m
oFTXABk/RGfXX0Ydyx73shARp5D61Lr3W5P3+HcLv9bgv2yGFfro4Eeh8CeN6DlB
CbbTgudI7x1+NikdnKwP/9Tigk1WU94I4P24j852rwb0tlFPc0Fx6dGuzZ+xsbWY
FUxU0KA4wy4K2AY0AhQxKcdl9s+CRuYV3HnmCziQPxAF9/reTnXvZNhrp353+e+W
Uto9/Uv1Ae9mUOODCDUM003txRN7XOjvOmYGT8IkKu//N4XTVQJwOI+h+dWFywAg
JKUUM8ge5yX7JRosPcy7RA7o8cnrwxyL1lbMsRqs+O7gEAy1Twl+QnfFRxJ/GK3u
gKu5KpBqM/HfywZQMAGLAFz1m0YIWW+lhc7OjXTVoGgnucS8R7Dx2HW1Hjv93S11
VMNMY+zkjuiEPLYsPxVdlyexZebvHPtXsfFDMaDrzDeo4lJ5AgtFUKrLs43puFMG
HKlROu/UUVCLDhxR10PBze5Yo+1rAm9O+ogdWcoKm5IdFSNc5t8RTC1ypIyBD2TS
U/HthEwR5eWSWHk2iqQGuzkA5S44g0cPEDxNrjytCI0S0VnKo8Bk0C+iiKa7Zo1L
O3hC/5jNPAC1Pgp3YwQqW+2muD6s2J3aCDrb0YfBCHSGG+OknLCDhCow7u5jmrLt
HMSS07rHVPLZUFzCvNK41uc9G66iyNvHx9OhqAj5v+8p8JI1j2jBXhBYi9Nog16J
8TR3q5+P80A1Oi5y4h+s2PEK5yE5Nre8cEIe66I4Io8UqLKXhRWRB+ILoS7Cs011
CL8P2krPfTd2GRKxrHXEZcP34EqYQyOt0vEyjpnYDlgGrcSe4c13ZYUD5rksGHCC
it0m2mIk8R+pgC9bPsW8V/Y6GqA/c4yqrcP+fFRK+Has/sX8mC9pjn8Q1nGfiQ9Y
KloJCn8i9H3FWCjBxxa8Eih6r7ZQ7PrIQhUhM4MRwW6K3S5kGsd9mFaSHZR69Lub
wr1hiAfYVJOArUhqpWhIxZLOjd7y9xt146wIIV7ASebta17W1WlTSQMel19+DNje
+gURkqDKDJ7OGU8JKZu1mH4c5POnDFGM1VTlzN555sMeN39UO4DfIwSIeLQTqSED
QSykuUKihtsJmUWbtWKrEhK6Pmay3mII4pRc0PyKtGAk9vvsUxw4YuKtzMxuHIx+
zOpwcNMy0kcjKDFPIBcoHcPfmtNYH0x0OKQWpEOPPlM9xhC38r79k8Q8nnElEklp
BvHCDSawT0bseV+H/D1j7mAHvdyQroIlcCM37kgfSpWkDcTJScS/Ddkvm4GD+n7v
/daonSuN21vBXtvMewmy9hq6G9YuPVEdM8wK9Lq9HFivqImfwak+ts8MiTAMId+c
EQeGvrl4/5+c0R/anju0LmYnO9nVkJ+bW3tcIFQAZNNy6DbdSsHJhr2sOVxN9Mva
3Z8R9ZYikshyqQ1QnTVZj8XUR8zsT2FDd9U2Z3HgrvVJ1agnFzKs4ENMb+k6O7h9
QaRVIqq+wz+GzQ3W7RdYGpJlRRDN5v3Kyn1E3eK/LJCyQFx1SH6FN7xU4BgK0YnS
/tbz1eljbYTn7+GaS4TXVC6P9fUi7Xgrtb4k3o1AzeVPT70N/JrOK9cMYNlWI7P+
ewNq43KvnyJQ5r4f/NrrHmhReFprvGRhYaNRt44E/S2Inu16aeMkdv1LS2Gj827J
z3/jzw9p3jTiWaQkzFdjRqIBLuIEpRcqxlmI9grAbclADzN3/CbVaIrD9u4/QA2F
GNZviG8EOHvowJw0m23IJEp3udmsIlYz9AzdQduncvQW0QBXd9KZbIibrehshjlH
uW8iwe5uXSJTkG1kaKW1ItcqnsnVzGuSmEopqQwKRK0XXRExj8rFo8UfEiaFZmpj
ZpYAQbDCSH2u0vsKoXrnlkN3/VtilHo76s89O0IY2Jd5gFIyhWgmlTARl5zu4s3T
4+sBa+uwo/8XSH36l7MBxIx/7TLhkHagaIGSNwkttWqQ3cvR8oBDvDTEmnSscsar
vg3i8P9LM003wqXTQ0FYvY2Oj4WL+jsdpgNa4WQMbouDtyrEAktbO5PYyWlxcL5W
6biQC4Kn+I1JoI6DHDYf/EXMhya72FwRDwUgI4nY2LqpDZTbZLg7ZjwGUDPOVAy/
5z3M+SlWeDZ1X4xsITcIEYFFEV83Mog6YfFTfkycarnYaeKORAcrNPnJ7cInYczb
pdzYS/CVrQSiALIDs0qmx3rN4vGBjSFFZaYQBktYLokT5e2i/bhBwTyYcNpuOnGq
nX0K/0qkQrtv3WeEYlJvW1ZEqX2sFQaV0P+KA6v0i/7hJV7sUh2t5CIWA4kJenhb
Vk3y9NVK6v5TEya3YC2MVjMhtnPhWgV8hFJDUTTK4N7s4oA7xhEo2akGCMsN4KbS
s7eaaHSDG0b1uB3KRJPHc456AjgSlu0o3N33xzfmnbOZ+tUxZu4nnzVNASeXCJOw
S+lbCa8km8XchZ3YIcu74NbkfRPx3uW2bst0onoVkgRrjADmlMH+JlxAwcAeCSWR
iSXT4PstIrlBdguithYlOuNKlTB755hsZeC0wZz5cGM3GnTKxcmjfQSFh3+yMqvd
TBPK5OL1PHB7VBl/1vRU2w0ac6wmiGr+KxQLw9YHkajuY++J4L6wy0UoHXSNe9iF
LKqUmiW2R3g1Rxa+2YTtwzLs1zmi7p57Yk7ODcY8paCJz4iiqdtanUXNRUCs04kc
Vv9tjm6eLQa3JmOJkqqBLJOg1WvWDUhMzI77RT64kVn6H31IMv3ouMzzn/z06c1e
TtuGypBaESP456Y+0evx4jQGxtp5DbLLiOJD7B6ad2f0kM0i81AuqXYGwlXUu/rr
JanJKhfWR68V/JPb261AarW2L175jyRRcxDsR429dqKKkieg4tw8aVm/ms1Ed0x6
aRFWK9klOAyfjWsF7SLk2ZIXUOs76wpwnN1k94V9e//2chHsH02O5HSLl3tegYGs
VXsbVMj8C0v9cSKbgXMmeLXjPEIMs8oCgMSeoLqFAVxn1jJ3S0k3Po3Uog/iozpz
j3toJ6kHRgaV9g4I9WI1CiQoi8HCTm/44wSZyowpriERUXGIFmLNBXQpBXAHy1el
TAHk6fTUsX84A0hUWX9YVrbZX2b7PAIo8zqe2/S6bUZPtmtpy+ev/FBXo8VqXYZc
IeDAOqjmw0mbMhTprxS2H2AWm9UbnB6Hw2ODRfpFmslFPV2VPtQzQjBqUDEFETig
m+UQKqZqSlxCn6HZRAzoxOFuPzz5rI7hFwmNk3mOCCBrE4qThE3tyxUsrvQzk/N/
wLMB8HNtGm68jHtMjXD7dNGkFGzl8Vy+RZtoKDrzvFF2FlSqbpFEhQFmcfUawTwm
hNCQapr9ZAbXdLp9b6xrT8K4EJNP2WJbO4JmK9t+HZmjNsRAlvpjWPv5Itq/GwX9
Q3J8XsSWgaCyU2j2Bnvs8xVkJa7G7BXEO1w9ngRSaB9MA/lrQJnrIPDS9OBtTHrq
pY4S00J0cuzfBmSAbzJ2fc1XY9HwZlm/qrycqHLBLrSWJvI7E9jYhPx5VSybEygm
VkgtEc1PT6dom46ZdXG0PT8nNYF6QkkI4SEH4av1HBq1vYeFB4SKl8uBPQi73oBk
UNstf0WJn5KoubdaSP90kAXaMVrpHoTD8dLc2A4m3Td6DQKPmiLhTvqCq8NFeXf3
GmIBPiPT1Odn6J9qT14t0P3eYdyOna5OJKaKM4o+hZ7jM/zot8z9Z8i4DF+3OQ9w
F8clC58oCRR8cIHdD78DVi187j29wjb3MyrLx55XQ228b3+Umng8j1cN62THThbm
qI/dBQgjUT8ZCj6Wapp57JwaHAGkuXaIfmoQIhAgKQuhrTKabwF8/C1N+IHkPMS1
Omtm2fI+yXk8VRf2uZf5MsUQG3eBc/cKRDr9Hv9VWLpvAtrOxFtNcYCcdG/Kjkl3
0FulTO8iVX8T9nAXxq//aKXYFSqvaF8ovkfODzW3xq6gIWiZThch7S91oJ0mRqxC
r/jhWJBL+9pVk8gwFkGt4AgHKCdU+pIR91eQMZpYwTD4RxJw95a58fcTB5+Ds6sV
NpaR7I9S1MYNkWOIbcfxFQ2U9iD2QaxUhrGbXxHDJ6fcxD39Nb135NWhYsr36FrY
/6HNXarTL2SMPVleW1vnjjBy1Uz39J4XXUt9l9pKRVIHDzSHAu72SOc8YcKHxbzY
llTQQA+EIGy6O1YXeKdvxGgDrdSjlKp7JH44N7W+jpeX7h6TRNycZUENr2tPdKiM
UMlrnjiY/97+YD2HZo7G6Fi8FA8Q6rnDBwejOelFX+bbxQn8yu9JdWm7H5baEnVR
rBYfWV2iGORM1BRKGyrtoeOUULymwz4mB1dYhfSb37jcVOQfmLnfZHDxSIZPPL6f
XTeresHA7NC0aV+32+cUWWojRFtD8QLkhvvqmumPxS4E7zpe3RzUfnhS0vTc+R7V
HcKjskV+m6Ti6rRIY7neeES4JVMSbcEjufJM3QsTqOHvf0OCCpYmT84dJolQTqfE
bHiMihvYw7r43tjVoFejhRlZorv/uadESUgjE0asUhqAJrOJZT6gfLxR1TMnuD6f
nMhZNTcX+nhzGOakE3l6bpeFPlq3qKcBPVxLn1wF+NRmRu5sLxIPkhuU3hotX9PF
VsmTVYiXTWHVAfAPVyRYgNzjXZAqIREvO1FgBXu4pEfRYt4o8TCMKtMosVslfIbn
mDe1Lt44ucPOYQBIxaHqc6mAuNkc6shUMsL/fxoJ1oebhvYZvjMBwe1UxJmoIP9D
JN+jUpf0sfT3dpoqTYbSCXTTMCQLQuivJk4kLQG8/9BnJr70/FQxr0zuWyMb2ozo
pnOJHZQsYygNjhKDIF04rcYphUY7HKw435YlUF9c5WHljm4aGmOaH13cD3wmAt4P
T6qPKA4Unwr49I78gzaoguIudg6WWB5Vrba7GHP8RaKk3EBpLB0rLdbmecXXwocZ
F+w6Nl8NZCDC8rF+TBQxk958gijL6uNHnmdxrv637dq54N5APWnt2V4Jop3cuz/1
4YMQ6puiUz3w/zAYLQ/4rXjOLdIivqnuQqr6B/ymHUYldJJ65x1Ow8b5idjb2RBY
9DegpsEtevA9FqfZi8kKExTodm1ks9QkPtTGY0zHQpytCZv6AiDmiasdVY6Py7g6
sGKsMMTpkv7yncbCKDcW1Tc3bXACWaAh1Y5RbG3+4WkWkkYSpMNJnSMJ+XGqQ03C
Qu7W6u+uoNlpQVn2IIiIWvkEx+7HJIKKh+cpcppEijHdHpnAL7nyYReFcUw5B2Gd
Am+Ht9kgNy8Z08acwu2V7L94Uw5f9Dm+z4Ag7BKM2RNwtweSXqDYAsz+4TEDng8P
tt/vHnkTEaUDCQ1n5qzNqZCxhL1JEMe0bwAv1tmRGNR80+cdGekHW5Y7K6lauX5e
ax6DQfNVTE6X/jnSDzFN3Z/zGxj2LeJFm5Xd5Nqheqe/ZVb4HR9k+qxFCbmcUNND
7vhbWNUtK4Obd9s/wkmstYj4cDwYi8An4p7NoljCepwKQ+ZYy+Uk9ASavtaSN0No
JEPGiT8p4m1h4oRlK9RRhtvld3l9+phqK82g3NRGMmiOf+a/WJZCcP8UA26benbv
cDKseIJEylakZZNIncwOPWsmC+jT0nc4WkrcqBFQQ4D2ROuQnX3lroOKTy2MIGTJ
qUH+4wCT73cLZf0/CWXCy6aMoaFwenpwqfVB2DHfhYUlFh9Aif0S7josMr7tZjvC
LS3Kw2gnWIHmE9IRloIADqAcvvMRW9zPSARCytl3hyAiQZ9lAUo68r6SW2de2bBY
VDUhcPRyyJ1m+CcawP3HX+WkYN88vLR4YFg7GL6khZe/RBotHwDlbEQqOzA2U5QE
qeShVJCzcq8Q0yozQ3LnB198O/iJro4WcoMVD6R6uKcAR/qa/EyPJrcu/7gSDhHK
/axlh71nceHfIIyUyWdcUEiW3W+1GNUrUTCdvRNx078lwg9pleN53m6Z1gt0XQIA
cEMSecveYcqkJRHriJVgDynU9F0tjdg0ntFjH1EpK3bz0Zxrx5ygjfQQhXndCz8e
f/CGZbMJjeBzHlVPM12vLoCxu9gM4qzykZXr0INmLHsLh4MtgEda0ft9Naj1PfNJ
ovZbemLj/s3B6vvbOu+TXY/WLeFuT3PUFNxzMxVNcuEdtnYp3HsS7jhYkv7GX5mE
6tGhOftfR9W0lzqu7fafscPbZl20JUF+kgzc9GuCJ6BIa2c1ttdERCYm8XGq+Rt8
Ahiif1Ryr802h9YAJw8w1AluwkYbBMY658AW/p0UpEY4t7HSpvNADfwvtXMUL/1M
Kd1ciqbu9C10CU6Wl3/4VFNN9iyvd8N09DygRr9Uz4YTJVrpCKMaSCXcwlsJOujJ
+OJ3sIBiHwwBHFibTG501YOVNAXGcqS58RC+dIcpAQAVNLueYHnthmxTDKw3vl58
Q8xLY/+OTgkIorBe8KNUhCHkczi+wuJCPqJEJ3R3U4edJxRMXoc8mnJkZ2smzVXB
YNFADxEpbQDMVokaxv6g1SL4pCk0vnt62amVyp6f8SDhkgs77FFaUl4BDdPMWMKS
D6EGT4meThRbyZyCbxwODv7U2RbmckPds4KjX+2ywV/P/jmlhjzWU0+z2B+FGl/j
0hrgjvEJQAptMdzpc/OA71jVWFtaHgpelhuUJCh5o8F+VLvObkkXAQv1W+mwTcQK
fPyTysdcHTsGJwS83gMa16kgnm1RqnBH8A3YMS41EDrXQghjyS+fGTlPldB3AeKo
QnyreCxe/6kKaXAxYZWrnXsDpXTWQBHETTX+goEACH5AAGBW4EM1/pPX6Dqy5vfT
snZNw7c2KNPPJ4yJKMWM1z1mKGdcgNhcUWFy4clEMHKWb6DaOhsUxLkUMgZcXOTy
0y5RjGoTrCglnbakLUdrZiNWUyR1K/aOCPAyBJL/KrDVgHE8pbmZTeh9L3n74uGV
L5LWT3C92YPzlFgxp+eP4iH/PK+TcYBIA8JOqR+Gtb/P+hDKHX9sOYqNEmhQwDEx
V3BDTYA1WL5SuKMDb6eWr9cpLcEbtz8VKw/BsSp7t7tFbml60WrfCr4Ab/9Z73nV
wDWsozW93dmbkvne+IDUZDP5vq0XrU0/XDe/LqK66ZnMhfCJKSHpBdrqk4V/VjhT
gET60CuzgC2SPYKW5+WNVVIaekqXYOSDfU0r88byPKTdqo1hWS0PLHGrwX+tsAeN
x9X4kDqAIvZL3Gnlrxe0orBvxfJA+RX2fJ6N1QoHprce/p2ztX0eY6MA3TCmUn47
KJqwfce2FkA8EorCNZkFm2ARPguZef++cyZNAizJGUld4Jb5Psag/mLagzmkzb66
xCfv6WH3Ru4to4zZtK+zcR8w15nwYKbOm61gvs23WXkqDJL4JLmIEUp/VeAAkj2q
NT0PxO8vVKcg+XX+FJ7KukOskIevhnLrF94E2Z1/fXt/rReE8b3N3BLyEcJI4vdZ
yof6PvHZS3S/fOLNAEwLCMZsuhBPvzakplb2t6eHl+z916WTfS2o/HMdE0jqU4lj
/74rtZlpkv3cWHpBurms9FooVdqkYWs0DXL7MnKDMZgCtPvgx5AcO0ybQZSfaUG1
O45I4Bh8aK/B4JenwQ6OL9hisN4dEjWzxKHPU7zFT0b6aVjnP0HiT+8LWmm8Ziqa
VviPve+UuzuwnnSN1T/5MPl6B0hdLzX2rZ1FYYemr3UlJDDhR7Rku5h7a6iHXOwq
APt2BmdFEqEvPz0R3ntqR4u3tr90fZMZa9MpRGsECToIAyepCyv9qZOfDXCg7flR
vsfb/qhEEdMNn+QS3ssxrlzI3kOoKkuJZawSP5brtI6c2qIiu+GZR1oeTKPExace
YnnBUKy2S6v/cE3DSW/oO2rYjdn1rh2jACxSbDc+sA6JiUiT/ytUgWxza0p396Uz
UJHXNpq+knO1yFDbHL/v3KAJUcg/bEmciCkikpk3Pd6bLOb5fJ9OMGk6r16cT48A
VUA2OEzB3XDsm5X52l5FCZdx/oK/j819mZxwoW5camljQXEr1KH4IFMMyukfgoF2
gzeL/uybrjCMci0bkdILb3Ax9z9lqHGZTD2PJzDOl2e+fTkv0eqflWqcQtIL5t3K
jUvhf+gemnw07ZjSB5EpKClrlwn50kZJNQmrYIPlFYBQcxrTq6VD5aGHv83xSohu
g64eCXjw6fN1KLRnDQ8MizYZDrolORNT8S2eEmS5QYVyfG4J0cKYhMYK+gZxkBh6
MFM0pbGuGamhDwOxCII7np6RdkPcxdJ/Hq+CTpc69cNexiXogmb18ASKFeZcxrlQ
WJ04KvpEHmWl+U5H5fCXamxlS1kjU/hWsO2CQrBQlbtSuuBA8TCST10wbeL8U8WS
2CqHHPSwa06xIZoqHxY3oV8zwRnC+8Ou5iZslX5b9VoBl5mCnU6olKEa38NLhkKP
vszW42y1mVa3OX/t8wYihsZnRVGJyr95+SWlLCnpz9V+lWNwH1nhPviZ1C5eWc6h
BX2DAI4duZU4E5i2/ebLwMz4BttBmGAAgFyiTt/kjW/UD2Md7vSPz1ckAcL2YRWx
VGYaEIiJa97DKEGfCc7OnW4i6nqkQmTu+H1dGcmKvIJKGwDTHGcn3WPmy7PQVhEZ
xJBbyLqu8mq3j1HhADgONBI4FFsDZlY3eiVgHzDYtWi2qi7ynNxMXpZbBLo0fdf2
bKEd5iaS1mNi6Puv4s+tP0Br3dh6j1tcmueN74ONZo27lpfBtsIDwiD5Z1NuQHKU
xglBBJBRMpma7tqQUS8TXSVRUVmBTHENQLJaDzl22yN7LBQZKlPlJI/5RJA8wtVY
Sa+bfnQe+UtSh0EgdiTxfszCYd0/DbV5aiZDk1GCs6mGTNGEPVN6forulqs9pQAK
uFn2argaDRhL7N98QvmOnuWkHqqb/3hDxESWOhMeLyyWnm410cGBA3keRmLc/0gp
u0XZMu0nPUoIu4nJe2+mM6ua1Gk21XCiVxyXOp1tZI0HB6mvEtYC9ifSOFaViBfI
LjgTO0pRULav+O4Xb2g4dDHc1mF28/ScrbvpnCAJ8mKtAEMYZkW8NZXvy0+f2ikj
SOE4486IrWDNwgGH8ElnzdUEdeQVBHyXRr4BY+6ZDEf18315Z5scTU5XvAd3/cB6
Jy7v443qhwbY63Eo2pAleml5OdHn3pzqyw5VD12s95PNl4QVMpHszXU0JvyWLNEY
S0piUQoSkf5tiigAFANzdtC+hkR0F+WYzvqYNB35AeKmKvWr76k3lgZ06ESchcBG
sHDleDymmiIKIW67HD1Ly8H3h9iUWRTjYxzvkk2ly7oLFHD9v/gudeMGpaK86OB8
EPe4zq/7EYC33zaCuBeno5l6tTlBlQZ+8/hUchVKo2vE8gmYBJ2jcB8pd3PUdeZx
iYwL/PT+I3NbFT/4515WSytJvwz9vuGrLVbzZ8uC5VGq2fzBjpok5EBb4GLZjIMz
XEk/q5hRqgcEx9mmBxCMEPJKaqbCwGNrWIjErc/EVMlZFjB7T1bo2g9d74XjEwhn
3IE3kozUkNo0lO0KX++aIlgdIpTPXjZoxgJ+4ov9WX7p1l4TNjSmMntOZeCUmxsR
vKSuJzHhyMyvMZCrJZHWwRV84/tbR9fdVNoXebhYs7LoBvj7UT73nlrbHe3P+G18
AmqFQc58vEvMwk9MiB7MSAQNSsTO3S4w6j9Gf2CIbw/mkVy0FmWbGGChjHPN/wvW
GmfVXf5f0UQGd6wRha9j+3atpFZQajWarJlvzGP6zKzhDiwNEJnSuaOZKsSKpQTR
Z2/KKen3kazV6NBeP0gYUz18i65jeprgJCn8vg0dQMsyr9PM69RGjVOj34dnadne
LyOjwx+OutakG8WVo1E5V3Jdij+0wHVIPEqjd4M3w4/O2kvRxr0Ck1oX4ttZu4e6
bQMgGPNgJ0sNEl/52C6qOlBOHU3NpLTy66Mxdu2254LLFObSM84/UhnyeAZUfY7Q
tGH7FplUpx5Cz59/MkUh9M/v7RmuQNlN9cAqL7PIDdz+E4CVxLY3h/FU61QWG5mS
1YuNFGD6IdIfe1ut3e1gAPn7Y0F8FPZoaZdCpxwIUya0gLGRnxdQhGCweUbfQ7m1
FTkK7M/lXOfAjrQvItZ/KxIehTjPR1LRMsObzffICSC8yXKC9zgawPTOKwdlUeEQ
vFdqk9o4sNz8Lil5d3NhDbimSgq7etnAyG/z5zjamkGXS6uvd+CZmIDEl8jFLOS8
kvnXJxSnxO6eTnxLYRuzVaCQ81p8158wueUW+kdvuqXhfX4LArl0hrV1IVVrlsyb
sOKXvEZ1xX29g1ngagZfYbinApVV5YE8fWlCZMVom0mRdNYqGX8fxeL145P72o5K
AuEjQsFiA7j2x41i+jaNKhJXcvKeDN/jBT1Mfsro4YKKXlPrNBwskrpc2zTnSRYf
XYMB8DjvmgQwm8ItA/AqqO4sg5guK6Os7bjP0xbQe+ICWb3vpfC5qt9ib+qQS85W
fj/iZefEEZHnTCaviEsi2NvLJWDkGgtH+asWmYGNccaa9QbKydj4KynE7ZkbR8yZ
hXVSaxZ1cyMt/ZUiHN466tkUFMwXRdlf9Q1XpU3dc5ZRM2qBluCCccs12TWlNGAR
pGWmw7aSYpWPSdQzV0oUAsgAvvK8OAvH1U5+eybE2ucLnBjEVbjDsUZG5T8D7kzo
56V/CgX02evlOEbB/IRU6vULb9eboW7bpzYgf+AFFAuWAD3bMypyvogjRExR9f5r
trAiiFqi3pXfVn87qlzj05ETXpXA9G5r1aRIljbsmAdPTS85AYZl41iUV/EJNRdm
Dh4pVsmQ8Tiv68H1VmzM12RgdNsm4e/fInu3nNn/cpJaGK3De46wvq19vIOJyGTA
UtGSOc293HQErjf1pm/keFG5/9OawXN59R+yQIBUh70qBywuphWC78F2lDRnzmT0
SAgrLKv9v9R0AZrNoShwRTpOZlzO1rIOGUbZ3NV8SUTQMNM1cJAvV40WtYmkVwBH
+zqFfqmOMXpJUJSRweGwZicFo3o0OJ0y3nlB2D+zCbJ3hW/EnLnxOkmYd0GK31I+
g0uvTjcdc2UgCFy4x6JHeo914Xyx/6zgA3DRhi2SJpobdhRexMAzls4vGJUDhTGN
QsATyOPbhaH01zPpv1+TRRt2SCmNxCQlBDVMTx/Y0nyjy0cBt0SzYrnwXYrVNcYy
M7XmjBuULoaNThJKWL0qJTGn/YJ9tqz4lR4DHgBxeR6LTuNnYDcVtJ2BiICqkswt
kAlms6munxGOK9GpiyVI/ji2G+SainHHiDZ82/pQBfOpO+ROYexGvja6fjVYINb1
VVlNN/9ZAL8dnKQbjjyiWurGJry9Sf56DiNm57+f8Yc1WDASD1q1FpPDoDKpzi7h
eetKHRCz88WT8x9QGVTIzYtgHUW6dDkHOxhfIaA5uxbvTf9s7YtBlHIPqwjLQIeF
hwvwMmiRehnZMJTcRM8+sDR+Qn8TI84ZCw6lYfIopC/va+2NtyX7tyF4J2HT6pXD
dlHvDWVg+reRCr9J3g5tWBafqsO6wePCiSjpnDgre94stmkAdGtNKQjGtmyhD+6A
CND9WmLrp/3P+p7AU9OLV3Au3ts+uE1P8tiDz+nsJvvILS8CtxzzEm76BR/rsUng
sIMJ+BKnioEjGF6qqARFOhc2XoT9LyP7IZSTP8gDKmGwQ9UEp6mXVxEzunar6VkV
3HQLVUSzSPHdG4jMzTyDoMpC3twds58h6St9EEWshyjZDaJxoZcwsS09yMuO5YJL
V6vxz1fFJ6XRVjv9YHIWYJDlLUeECERrOA1YGTtfBudz0zPUtJ/5xVopaps/jKpr
pylrsEOL+5EluEKCHFqW55k3hMdzVgk+741cyAg31eXwieYL3pSPF5vyylPvNDrI
P4aQ4OyxwIBLy0R0a5Fq11/k+NrGTRI82iVlg9DCUOSHEls/m+5cCXzGAcFZ4hqr
hYahT6y/ZYvq+zZCcK/RgZPnONFAw1QzKjR0t9mYMekXaAnzoiHZ5A6pX07Lh25y
NTUxu0TElEyDX/5H1tYEMWfC8dHv+G6T236ntAsbm75lSqFraI9n3TZbmZU7rp7/
hl/F9n9XcNclnbBBhw65k31fhB+4GAdqvvcjL8zZRzwmAf1zO+17zxiUIoBVkV0B
wtORXSRJN/np8CM63psziEPl4gFX+d71OVQ1ory4ONVLITrZVXSvZyS/rBAApyzD
iGaaOkixRm1YNd7Em5hA5pXvMtCWUfNCMCN6ns9XQ6UWL6svSTSE8nnW1nmucPZ8
E6F91yp/XOSYMkpwr4zZ1vdT7Ia1n+HT+i14TW8YVONkRFqRgM1d3v5ec+yghwAp
i8fRb+ERutptPMM46TiJgNBuxX6q2ifENIZ+JZ8QDbcY5SaeICiPV/THfMfNj9ib
PDdjLGajf20RkcjMtNJnQSeKuz2eA7TEvg2jHROy2RTkgWERKdExzEef+uwRgwu5
2E1qj2n8W2/qXyPD6tSlzv8mqALnlKRqnl28o6+WnTARIm3pxciiAqrAC0aPVST1
ruwKBoNb3+cSXz1M3ubC+lQfvggrqW8my2zW1VN+W/FADCqrfyIMh7nixyEYgLh3
RspzNmY3af/Zn9nnCcVVte6kC6DTuEzvKHz0gDiLUUixChG0u+YrlX4wwrRJRDnd
T7anKPLFyPYMktLoPKT9ayd8u4Y/wxX6p/8fyTZCdqIvUi6w7xs9tXfEiV1N5d+f
wxswCMMfDNDOry0OujZ8caZ5FG6RklVE5+WP4QvmKltb7RjqSWlmspY3cmvLp0Mj
rLyhnO8Rzs8zx4mLBK7fGV10hSovjPkMViqLv9sMUm9xndrzIr8HX8d0PygZ/wio
xKkWMhQKtO2zrEehih8PGgBIQQTZ5MLiYpNLj81cS+5hwzFnja/cR/dZ4zYDA65x
H2T0fXd3gDbBpMdOZ0XJYalnFnSXiP0kNBcFlq3a0bXuln+XIBcA8gWey1BrNSca
/qioAzLKO//KB+AI0V5l/g9E/CLsiPmvVReCqD0uPB6g89Xg9ojkRnaBQDm6JSoH
Ugh15lnbBM/5EQCvZb5+d6pd71pq7HGKRzQH1SRbqRR5ettEmk7ThVmilrWUn4hv
/KwhjKDiRSYA6J1+bbcpbNG3XlizEcNdjKzo6u7WeI43fH4a6JoKyHSsk7npyTxY
x2J0JAFLochK9CqpADHmTXz1pCKfuQjnC88ZM1frFdxYmyI0Ur+v0t+jx+agVd7F
z6aSUgr7IZMfcusQXwYidJaFfIc5bxvWTjXa9sl69F/Vv+yn3qFl4kYsq0TnbFOM
2SsACbIHjGot9uDESK3bkFprjpNuMI1LAV5WOeFfvDjg558P7hS/LLTs84NbUeBb
b308t1RD5afsfisyRdvkP36Rhi5y5rp1XOMqDsGl8lQ7xu2ym1mtPAO57ZXCcQxz
ab2EndJFAqQdzJFnfa2Bb5uqZrBcsSeFhSSME7zuAnTS/rkaC8BHT2baWFi/oUdq
T3LuvOLb8DCen2S/TxnzsYV1yi6S/CBuX4Yoeo+pnA7rONt3pno2QppZQBEviHlk
l8+7JQkQp/3O/sTq6p7W+oqlI/6HnZgfuzLSxrtHYLsJLSWapmoYYSagrADOv2MV
N6g+pnhaLmGOVwxoWkmUFEsdwxO1I71Y0C+xCuLiSTn5Iv2zmOZjaJzQU1Jbvg0B
XqEr8J7hB/RjV2ETOorMTCX+5l/z96AlUyU/zrYL/JRhnaGMW4FcRRzzp1FVTCvQ
VJcgAYrZx0WywkWZV0tH4hECIK8CLrDIULiB0KcdwHNv4Xh0nWcsGLGQ0/yNc90x
7sxNzQclQhtBlhEgHWJnbIoFGPzvmyhhHEsteV7IClGOii43xeMxEvSAPgFaFGZ2
5W8Trs2GvTaqlEefAmuBGPQTSN7wCr1ozY4bF/TopN6uVc5nVApzVp2//Gvte12M
5d774taFFaZrLVYaRO827mH8o6vnXNFzDxg2s7OkrCXsaVYzbByysU44juKaviqq
wBxtoj3iOGF/3pTwlJzQDHBd0vHtuh1bFUL2rkwHEHT6jL1KtVvbo/s8ZFiq/tDh
hsq9xT/RTWDQr2UN4cD6+UW7wy320yug9uDlzvQozhmb38/XXuvi8GWkOB1e4Oeb
mAo3PDzTfe5BLSH2TBWZLQ5qUSxEbNRR0+mRIpdfM1PemIuGos+fe4XmfV8t49tp
0WJSt6jT0h8HLbtdVu36Q6GM8lLAz90h7fSxeav9qc1J6h4af144LpTXfKIMY7eC
VvwtlVo21cPwsJo60dU+TUZIaq6W7fzvkIfveKeA6Unx3Cl2K9Cpth/HNWRDOvhj
IDvneI7p29elOBT6xxr/1Es4tM1dWkfwigRjHW81dJ2sQ1NVDgeWdZY8JHmOwERQ
qYyhjdJPNQR9dQi6qJhRRMyVb4CkqqIagoRxUSquSr+or87Nal6LJquTywfNsLxN
e8sV9QhZiSBYY6iUp3eIndpCepWBJsWBtfeRiiISJzN6w13AahQAIH0rihxM2gvY
GCnLvwfCwWTd8HfSNCtwFSLD92rDj7uklxmZePTDryaynUR9NR/AqA0vVQKA7gL/
ad+CE259ZtwRtajBdw8jpFXJla3nEoshLmK4ciBHeXwN9KD+oqCErm3fEacb3VE9
IRgcCOm3i1YxSkNNnsc1+mky+vr6RuA8Mq5mCnjN86pGtKKHyZrYjWQq7HEJr9vc
WBaugjeGLcBw6KO0ICIVMYVgr1p6yXUEbgNB+CYKNzJRf5DJ0wllcI02KAXk1Qx7
OgyLa4GBsMFtwbnmVb0V0QGg/V5UeamXNybpommnEXQE4tJu0/ICo+FL6wjvtc9l
99Q28ButyvgL/LDkQtZulEnOnoiSaCe0apUoNgc94dw7As7fXSfBvmq9M3p8EmNg
R1V6YtJMyAoFfUDDTd8V4hyFW2+bH+SSgblWWVnoZ70RdjTTIDZFvJfz83MX5ulv
f51ujw8OEfO/QBOzsUc/eIeEacLEzkaAGTlCoDIa+Ex5UAZAkSgMNeH0rY5ZhEkl
6sqgxpKHnKvFuDqSS0XrjX9A+oaQx6unc7WaM1vOUJbMQdBo2i4WpKLDfqJMphgk
KyJdbDxmUzsMbd5ab9h6yqxn3eCM8VVBINDkF6y2lXsdBgSuohA++/KkMHkmcXYd
kZ3muYmU7VKFqpbh9nTNQAwNadppp7tjtZkL0RMmBlAowH0Ow/G/23wKxGk8Ufv6
IxGAs3xYO4yX5UjDgNethSKY5d2oG/ir1S6Z94Yg7lQHsWJCQfoia3anUQtfq49I
sERTUo09udE/kqnMf42m9E4TtLjN4lpaJyl1m1ulWVTT67hm+xotwHNB9CbgmzpQ
xFO2Q7jNtxKbnGOR5xFYarZOaxcjWx/LiHsU7cstNF/eRIcLtKR36Xa/vRzUsfzs
sKJyOMtdGTg9jO24EWpMX184VQ3Egpa+IH9zbNXUtW+AW+msQ/BbCkbO1AkX7IPh
MM9nOKbqIiD+kJ9GwO4bDTrFgxliJbpdgLEZ3bS1O4p72sHjfw0xbLD/L/V62Hwd
JRT1gRqOyLKmj1DOwC3IUdbvvxPxXOkeKQ5kDSZ1wvxaaTD6umZJleFk0xWQcaul
fbNpe8midoTUnuZSYc3kHeFHb3CK/su4Ecbddm8nd/Of8qWBGkWdSjY7MCVMxEWl
w3Qs8nBv1xugWxLaxzQB/lLz6eLnNKkkB5NOB8Ell1u9LglJgqos+/Rr/3A6bjKL
dRMs6Gq2W/ukMJras+zUi157LUlCGIHEFIdDw9qRwF56ns3o2EPiVwXvzOUGxN+9
1MPdAii6BjtqBsvdneib5XZFaF+M0/n5px3s8tOeS7RAOmEzm8mL/OscXo4L5eMU
PlOEsvekSDFW3juqV3Ei49svIDFKMnl6mik/VWyKiUqzyyeVglpNM28RuC5Ktt6z
8EP6HfzEFsGIOQ6S14igQwoPTnzrPZh5cDyBGh1URPoOpC3jxpyuNIdAE+WaJOcH
1u1fX3nKF4wy8mujjlGyQkv+8H+VgJ8qSVrXremRRdGJMH+9pmTRNlp7pjEFSLgP
JUmkKs/U2aNrVoF09gD020wvQHwKWP1YU2zTSlwWz1MSfXV+qbM9jJUDPKwo8LfV
RoqOItcx5nC/p/iqZsEH6+XUEp/TQV+bEyH5n/9e+CD0RUTF0Ua9+T1gOfTGfOLv
dvJjLahrKoSh9KFa3hE1prHO3G09fPmvPbj2OBDiRAHNf/SAMEzaJNYxm7IFLfko
FnwfQicj9zDBS8LEuqM17qAA37kTkGeq6RqZ6PgUnHUgjL6gmUuAK0v1Tfpivsao
nmavK6ocMcOVQyY0wqEwH8ElshFGVqEogoaFi5/pvLBiDQRo08BYu8pb2qOxR7s1
g4BoJK78ikyGvWiQvTtFswpu+II0ykFSqEY0fA23Bai2T2oe0ZgJ0nvx4rrveoKw
MLN1V5dZbA2ZhqBJNHsb6mvPQPHeMEC0ZJ/hzLpfc9OEBLbxUNtkkvxJUQC6f5EU
zmTyRq2jZaBBvTSS/NhnniUz5/WvoffdaN0M7vP1JlZAP8+cao2sf8py8h8h037q
2Cl4nfAeOkWOznQgNe1TMNmDNc79RSvDzcos/5YBIgAMY5hpNVdecCs7YVE/5B8h
E06X1tchw/eV3E7QoZlpiLXGc6YaS46NOQ4b6hlLCodTmjFtbG1SnRADPVxm86/m
YxfQz0TCiWLh99CvHtrM1gx8hzburA9KmvRK5Hiwqt18o5ge5oiIpDp+IBHOMb+u
KP8feQ+BQqoArxvuBpZuzcxOpI3V6e2tmi3XxnIIAI6RTQrY2jgjNu6K4sJozjBW
oWB4yemTVaApvvk3vlKZ11R3OYo6lyo9IKZCk7LugXSkHi8S1GcRXKifSLGK6Ay0
j8NgbmRV2IzkDUbLEsod7rBfAOX1hrRriwE1ZmmlyhFh0ba0ahWT9hWXQESb98db
6jnBW/PZtfiezwyvFTEtobuIXPL5p4QmgcI8hAOoE53Q7bsOhVdQvneA39NqximR
YYqKzajktTnihY6v2QFDIGVks74/902CinM9kHj/5czngfVUuy55kKjTg/SeUEnx
PEvx29iakZe76FGnwzw7+38dfYFdCm5gS2mm+dBPekt88jddlnkoyq+Hc3dhbKGy
nMG9uUxQ5AzTbz2eV1YGpRnF6lclOtVMcV4K8pUpiAMf6tkCmZsW8fWpdaBCoy6a
hUgiFafRecnaYoFbKP8ynpZccMa6qWKBftd679wKoVQO2YbxF+Jzp/i7rY+lnlS+
i0HrEkuGsdeX8GieTUJ9hJILxTdRKetHePFuy2xGsbeUJVYH0LRWPNX7eY0SsoBv
XaXjFubxzFInvOowUmVxpwO/beLynQF+C3XWPJuBiJOXAlNJtCRZhS4XF7mBRQx7
Q9L41vm5Ze5cJFWlcoefEX+lv8RvQJ4pENevDBo4K5NkOxV6GEZHdSgtpUfgWXmR
kXVQ9lIhamOLHO0jsLq14GTz7WGEkicbzdmbJHYt9lZPHBLFi8zPtBpqdsGz4tuJ
TUjkg2pClK3zT4FZ5YxO/CCMzRNA0kXuvwvusxn6cfFWA491kd/4WNsTaZe8jeol
nAq7kX//RBPa2blix41NVEGX1Twd+1AE++eXktg6+YJXFrWEz7WoLoywcH1qMneL
KASl+4XcRuBgbfvF45v4I5I1TFX3Qs4cCaSmJDPpGKjoA51zDs87pf3RfCJe82bx
K9kzxFciDkqVliiL9GiCtPLy5N710mMSrkhHN/vTvclQfDYd7h9fcnEMy9RYME8R
2RAvxt+B4QjYYztNO4VI8+hJ+m0PvND/IXK7F+qeP3tLuq7iL3VnLgW0fqPS8bP0
eqMLm1gfCDrdCl2ArGCYOfOtR7i8Bje3Omu5ZHwM4MS7CfI6j8yUbnzyog5XjKWK
clqBcarR1gfYrhsMENef8ndmge7VnnCp7WPctAljWdfTfVRLKidmdyWFV/pSh6SX
EkG0cofGR12YwQkG7pfVQIXoLh/cv1VJjsKpfzPKq+3jFfDHApFKDJVRPtTooh4c
NFLgfrWIYJnfSo37qDSHddNy2m194HOn6SMPvS1xEAKkGiqMAw9mQw3MEfkSb9VI
a6C4kgvoPtxBGYkgaGlnc4Rq+3rFNMpBFFqojaxS47d4zGs6FhNAsSfGIwmaCsOF
VetJlxTDHZ4cfW+X9LwwaFq7hqEEh5knnS1Lp0DI5GUoScqnRdzymnro4FIOVIYQ
LwZnpOkTs6oYZdKMO2AbjnTdl+EjJseaSoitFWK5/GYpohyDAxZrfXLXngAcMutc
fGPWowc30y7BOr8E//SgzhWJjsbooEc/fK8Gob8iafAYiQcw1EIdcCmPoXP+LuHu
aP2LDpApvFOkEK2f6ANyU/HUQDFDk75bCFfRhn8hvrVMWI/vIP6Ra3G6ou9Sphoz
kXT2DfZVuFbnibUmA5fio/itCgF2oDqVOLeUX3qTeniPshWF5Q9hKGvXRuI1r5JH
vCepT6NlHSekfbxjBYDDVy4tNVelXND1jcuogxgpuF3tnX55pdFA3654mIMVS1+R
Lrb+9h230iUjqUsF2a3HzWVPbWbQOLX6RWACI8x8uuXivTltvEflSyRq4qX/HB1b
zhFFMN3o8+QCyJgZitJTWAnUdpRPQAqTcvL15ir1eKJX5BtLKeAizSUWDmxHj0m0
zjb8NIgDHdp3yYySnEWtihgWzPi+9l+FKlb6RprnNmbVcdQAMhC9+t9f0njcXVGb
OHJzbW/a0RomYw5UHICPg+qPH55p4HChzBRgt32Mzugof15yKJTJGx1boeFVv0Lq
piBNbhHj9hWsvG33KCaCuSHt15rJNbQX0DzGxIIStms8uYXOsWqBs+ZwMWkXlIP4
Esztlgu01wmfSXN6RkRVLgQoT5fhKUUJwwx0wBcKXSDFuJ5IKe8lJ74VTdborCrR
dKFG7YaXlOLrHS7Elp5ocxyxCUiyH6BVSgtj3iSEJNuLb09FNrGZ3EhGoBPEPiaA
jAjwnY5glhP6RdpBUO7IM/TO2HEA6YYuSXtlzZCRKQylDZ4++sWaevThqNKzOh55
c1z2Y0w//4Ci/FxmdTXqeexB63xmbj0zZ+D7/L4ZATGyrk86DrC4bCs8in87Rs3i
wabtT9tQQYhu3IHH9JBvqGQ6KmZIeLvzX0IYnruo9f6S1AZwB7iA5PzIEYSUU1mT
vN+ZDirjmAojPj4zi+kRDUiAtdkmnShCgww4WWLVwby3jujJfVWN9tTE7RpLlLrw
G40uDvA2eksKCGFzc/FQBNO3Dt5AvZYATubny0njoiy5eH9/JI01tybqeLAVOQwe
TXHHaM4aLfmFP1zDvzqhEtoTm7xLLhektHKZvbWz606gFKTdoFJTCNCi9jF3Wnfl
VfBN7+AIDGKSQVuYfSQlx2WfY/d6Qc5bgs5PiXSpV1PcMNDd0I5t0U4Mz0wC8Pko
ZggbTKR3mmhl0nBhaU2HEbVzwYpIIMen3xWd4UYJxzyAJdqK9emckCcgC/WU1zFS
vK5oDppBFnaOIEiCBHD+hCrjKGqO1OzvjnldXkqOi7FLheR5JqiTCnSpEp46Hk8e
TNxJv8vwStYlvaQOOxWIyqbxo0OdrJt7CTF/+L6RhzmIaJMQQlhCbD453Z9GvhVi
txuiOuXX81mGLrseWR2Fe+4jrIux9O0ogSIJ1PkKN0/NRzHh1AjCj2MrvkUcCMOE
Wa84UMyMcIEBsfQlWd/FGuz1U36tqxTzKprxjZ8wScif44NTwdiPyqsVQCOBWUFp
O/a3LbzSYu//knlT6NZMuQGGiDtY9nBV3g4nYvI5r35IwtN1+NO6q05G0R9tYC5B
RJ6Uf/sm/AFmxr8PiDSiNicCUnBXtS6mgJd3XYfjHWAkYapqfZqxTjCYxwSs5gzi
AHnLMGJP+zGMwDf+v5SvFp0aVw++8ePTw+1eQc1WyIOaI162JtDJGi5dey8hZ7/P
nWKxt3vH+eNTq5Bz+PFwtebvGTxXUiUJ3NlXrnn3YkTjjA+3fELArchNxzB8n0LZ
/zZqFHnyOU9I69AoXSrzCePtXbjBHDF7cwpoO3i3XOx0qltWsAEHvA04AmgI5Sgp
GGX2AdWN6BFak0LlKOeWeNdf75oUzvOFH1H/0w/+aXjjO6InAavn1WfruMARcEpq
/0SviRID7zBwS4zxhtkaioq4p/s3LYOku/srNPotwpf/xaR7C5nLbv1tFi/AltWy
xbTQolB8EnxHYKUfJADX9FE8hIzqLUCPqDmZy63SDg2X+OINdTsUTdsyzmLQg8d7
zD3eVBkV3HhqwS5v5ruvgeJDeLzinZyY/U7rHdmPdiQAz7z1JIE2bAel7ZG2EyR4
GwB+Zs9O2eyY6rwubDUN1P6R/X7IunaUtiEGtuL6ZJ+oBOgSvbHzlADsPUtu1rZc
uESfNdLWtnIzv35wQEY81pqnaF7FpSeE3kngAxyHT0c5NCbq74OWSV6omqJAg+3p
nN/VquyOs6vuN/Wm/amMMOzo6eAM/jrD0RKRz7WwZETbAPxDjJzhEAzgyGNEfLB2
uaiCrF1lm5DhbWbQ2whx1BhA7LUzp1Q639fmU8UZmVPMJP59Jdf3eR1508OGQHSc
pnZt3mERmpvI9E+kWBsOYHp8K/Ho7ZcHdgpeNWeKcpYlylS+j4+AxE/r4fd/SIzL
ltRLoDQhXvWO/9Qv/QBWl/09mdBp3WHdFl8hKFFfdusBl3Naz69hYg2qBRP2xRVi
5IXbj47VMqDVKlV1Ed4ynx3qIEzc9/bsTdyBOSt/AkckiyUiaucBitx+96zNfJK0
8riGv9iAvHSao5+cwDlfcQq9qJvcSTtTdkcc80AUKNiotvUZmRxC9bYmzW2Z75qo
tVb3UGXQpsblSzns2pXDKBTptE0XREVJ8mC9O7MkEAIiRu5tl2tKKd3thXfWDj91
UKV39UctF2sh5Hp5hkvAkZpBDoOYxu1yhsJVvXwmOGe4e1Pled0RS3Eqwi0jQdBd
bHOyxs6hmqXXs+TBU3YqYc1cNUamIe8yxwHUInkClX6xFgNaqKBYSJb+NMbx1Gtm
wuMoReFxhVbng+gOnuq4Wjun1lWQSpq7jT9vxbVukjZVdnDm/MOzSbvIv63OprG8
rwpRXAdCx8XFs2NPqmZzUKn6RgOK0tLkr3sApzd2CKl58iqS/8bB3mNniyhVtF51
uABfLumaENctQLOUfVzhrNBTe62GUmGjZpSSgzPsNKh3+SDZ/RhgYr1C+1m9BWOm
BRDvUaTYfzcC/mujUfSxJRc6/0i0kY/s6PWSLsf0icrJKZluq0jvuJ7H3H8Yi3JA
sTqJQOVcJ2lw6ujKxed9slC+w2V+pFhIOILzIYo05mHF5CuJB8YLkKoLzIYcTFnV
GQMtoWw4i2rjrdfdb9R+oHCbeFrbnWgNhxI07Af5G/4Ov+J2CU6lTgoMDxESVeVK
rzUJjU1d+WJPvx1DfHXa79SSxd5dB6JMd3DMzUzDbY/9yqyP0nA4KUi9llSlz6bN
+iZ+mTyLFls1MnOTXeCWfIbyVzNsOk7JpO2YO37ixTMdt7wdqw5PcnqwOlUvlVYX
pHyhQ0Mt/CH8TEaccpSULma+f0zEPlGhwQFf09v85IlSjdIobhTshO/eoak7ea27
Jfm6g9hwIYpb54F4wGupwHdapDz9CM8KBlh0jbA2+vKptry8gqSqJJRWf9EUoTrS
QnyuC6acs9G1XAZlITPDec7tOfqUodAbpa0VDHMTJ0EksD+zNSo9rNPgvLoTNwpB
TgTWMeadzflwLDytnLJnUXfQShUkVELYTonJB7Q79NLupM2M1j0EzyMv0UGiWUCV
ewUvL+/lZsqtxhapNORr8pKZja0xKjrE4PA9RvZJxQtJzya6kANBFq8C8qIzui4A
0kfXHQB+OK1r108lF3q75f5JEHfntckz0GOyqKqecJ4ag7Ebbp43qg5tCvk4v7YA
nV7eflbmRYI01ciGAwhvtIxlKmIev3VFTgmCXsqgQXwGg6eocwc9XQNIj9h0i3aK
RE933h68KKgUpGJh9H0siC+6LERTFKCF/AQGu7Mj7SbowN1p/XbH/y+mC0o0uGok
i+97zsNp9tsmxoHp5k0rFJYR5A5amNnrQ0YUGcbP86JKCK832kH1WW5kB5JvCmPM
kZyHCt8L6V7jIsUYgK1uPDrrGYo6dM9/3Im9gsDvhrva5TVmKrrDROapw/6msx92
OK8hlaA+PRFqJwM96E81HKHpy/GE+2b/KrmPAxS8V598VNhAGGt1rAmYYFuTaWY5
yCSdSyTwfx7+CokOxkpFGIVBXhY0n8pMhZcHA1HmuTX1l1ZUBSnWsyUggbp9ZQ9f
SgKzsOUF7dJbgrwLFW7RzORj/4Bma3riVd93sYE4om3zzqamTHftcxAhV6r9RBSp
p6cANcrBhCHj9xvrs+ex7FqejjlbI+Fu3iVpsFJSZg9gG7+hXxVL1JplsVR2UxDH
xHwt/muCcB7Ru3AWyJQt3SDdQ30Zwtd/3k4+txaSmIxba9HGiS0eU0I7VLUOCC1C
SiDMfn3lqztQLcEqDGE5R4OmmBFShglO9UJ7JRPsCJStZ1BFnClMs+kHSaaD/QYd
i9skDaeMrN5WjPwYRdK5XU3Df8taFmcvjCaEbQ9EgbhMrF2q/Ibp8R8MgCa0Ji5B
6cODIlg1B8rBGy5sUqGHEnsoE222/BWVfwU55nLxFC65KOi7L9bwaQz4zMr+UgWR
ifpfC9wjsdZeIXXEdk2ZiRJMO/7wKQeFN0PYPSaNySJ6qYdiKXSU3gOAKTvzfkM3
4FLfVhlLygH/ioujTWNlpfh0nlO3AK9ib7OdMy3qU4UQ7ddqRfm3jyEPcnZGrW37
gtiV/HwBZAVmxCZkrtFLtKeAv/qHgGmBphoIo58gSk+OWhYh5kGmG8AmDXZozlnP
dOtgFG7rnAXMiEtsyva4cjUCdkYGlp/Y4uZJKOp0iZ5ZewQwVfa4RN24D7l+BdQa
dmkhG70fTaM3pAWB+FUkT6VQPfiS81iLRJCC9mFd7ImwZElGlOOEFOJB4QoHFmtg
HCJnbQNuRnGQS/cuJEEvkkwsqG7yz/yyetXNeKKBBWZ7t+pB3TcKy2Wvj5lPArA8
ylkRk1E06ImDr7Ka4ZkdehyFL7Xg9za6CtOg2oBlCWe/Q+UPrzHBFjyrpiLK5H5t
KtqiuWJNIGifwx880FV1AQJw+VSB1IGHY15aiscOTEFxwNpXg8YbqYUog0X47rph
LWHJT+fLeIZHp/zXy+fZ/NUbpZfMlLb0D2sNTRIfUnWc+KCnjLuJAkbATjFBcHIP
F/1jNUAHu7rEZ/utwJUNbvKvIMvd0Bvui0KTBshacyI2hOIgVqCF+OarpZwnfUQ3
XTgHEerZTdTEOHW+w2AXssnCG77ZJRfmlRS/uiIyy8SBDKMX8GqNlhGS5qIIhxgy
TGG52E2eI5TlqtBxeADCC7KSCku7JZpYwaPFRNfW7nzgDwXYEAWBQY3iOboHNj0b
WuN4HYqWgVaT6td63vxZXQsONQSbh6S3fecR6/lCMKnfy5xRadhLLgdJHaMtIBW3
t1pINohzS3LavF+JLwKuEhoYzxhn3/gwDfTNZEUIvShiEnWTiKQo6qh/eg/hl+bB
StqhVK8GjOPRYyGB/K6TUrv9ZU+CAERlrLFXdXqYlU2QxnVJnw7oflSnDWSLOUeY
ETLLzuBH15F+hYUeP/RuOEmrrmPWptHgVWr3YShq2LOHoclwn5nwvNxwZh90RzX2
Zy0z/IHFBgbEXKbbvey+PzDlV7/suCcx6y8CkysvVCf7Dn3nvhPSMN2ZcT4Th1H9
1cNBEw3eURbEiAAusQ1VcRV6vLWFwLi+9Oqa5MZKK0mioG4WrYVD+V0sihkMGNHH
1aKe9WhQZOkavBXRlYVrh/H3rCEenWeKJn4hDTMXdHuxO/A68ra6H/fWQnhfOteW
Qrl6sGPpurg5QASTBHh/i8wZk46p9jrFLSHbJRs4UkNiCBXKAOf6E1U0VfeZhXXs
njRcFdrUQ8O1g6dkwPOZRxVLYoa/QrpWzLMd9ajr9Zwjp6WC0Nt15w4Fh6glGfFk
VepKAFswVNFQPwUNvOvztLIyh2tnE545/4XX2P+uFid0tnCRWi6T6OLbKT48uLsR
USTf8sc1pMhnlnvPnGZBFC2YFgYF3ckut0AEmRhRSiOu95vWxXoEJ2VUAgDeF3Xq
LvVCcheNT2rpK5YSF5s/ThJKUrPzsO8vKDd7NpuNmDn5BvPae+NU3AD8tMzHa71d
uIw4qzT99OGIl+Gj6ttwABKhO6ssrI/XUXV/MOR0lFP1cO2THM4cnlndDKyVQWIM
LWqsheCdgKvO4yX+hDrWfnz24s4iV6ts+BN2kGkJvLbM7vCjIhPq0GnsXsU2eyJ5
x0wkumB3nNOW+ne+8f968DRTmcUaz0hK//wyHcc+FrsV0WneY2Jbzmv7QjtERXH7
EiYzY3MqeGGHLH2l0L4EUbcl4XJiIyLuV3E/CpTzvl4GULAnGRS1jfxy2MTbMxT7
MLlO2IONl4asroig1PkfT8HWNeolx3v7CDgh+YWVajeLRPZGipxyyBzcSvS/0umm
EwqO0ytjqdVxAjElwGrsjllAsg+cBt+R0ITLEx4r1PeacojTt3H5yC3KbChuROyX
4qz4ht8MYNFn74xhtBNrGMOrT4Okfz49l5XQW75d/hN/BnIXWzPd0yFbAvyDnfHS
tbEgvfe9vnE90fNDiQSG79br+n1W1orG9BmHtwIFD7yCA/SidLzsgIlycHW32s4i
`protect END_PROTECTED
