`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWnZxjtbmFdWZpZ05C+Y8itbhgKlmK5r+NyDIdws/bK6qIpu4mc+1WGXBarvrbRI
M+ICVEupJ9yMZQlm7iaQiVCtGa3c2DK0uTCxNt305o6gi6GyMU84x9zcJCdUYrxp
YI0Wp379PYkCgWkoYAyvqJpKcu3qV9iRn0zFkXusbIL0zvauJsgmJtB4aO3egrAY
WISpzLB2wioe9FeecjQxQVVjLPdB7hx11I6wAxm8Pz/ZXSBs1jWhDjif8tTWh7x5
Uqdz2xiM5IxQo8fhBYMhx6N6W1d7nHNRr7F5fJv+/JUCL+nXZD0MXZJ7SQzHPjtj
IHmWyWrIUbU9DwCUnBZeVWfHDuf7okr+yPn5vEtIVVCabu8Av3hki0jTuo3KD5Dj
IMY21Uo3s12cXN72UdsjIstdRl8um/yBtv2DwtbLrpSByRnjbKew0/pOfD8CFcoS
B5MH+GOy9Pc8kSn101qFJOFzjs2N9/wwJh3uSIn8ttPmB19DHHlCEDHayMgsu8rT
SQq4e3e7oc1l+6ejRSWRQWiXmWZJ+e8UpT0+CBgodmmQ2l/pH8fflRM3hvKjxYwk
twP4I7VKim9VoSaA4uiDV/zgFCGmu5t289LtADtppR+UN0VPl6P6Pni/kPo08osN
XxTcRmJLFiSz7BIKlin7R/ipu9zJZHD9vuAtV/9FImxTh4Jd7cYM4/hEsd9FLLZr
83uTl8B9hITlud7q2jpkbW5E+PpVBqvV6ywYH6H13T3Y5/41yncKu9i+f9jNYQoZ
fbyKtgpZwPXdUOwMaWBJQhcON6NdwOtf/U5qtrjUA4oQkXau8snAnNpy/i6p9828
223Y+jCXcMRhh9ZbAOvuBHPWp/LbRC1T27SiqeLTr3CkkECzAile3nEToHnCEe41
HW3XmnwjXMZJCZxuyzPXVpQGngA5TxjI32CgOfcE0y028TFAP8LS08S7NKxrN5tz
XTvcM+ozatm9cWlEkbHKXFMlIjWoQH9zqhMkPRG9UNY8xWmMsI2WnPhxzT2K04xi
L9/hJ4b3+xvw+e9xCkgM6g8m/cs3VtMPxvqUPWrrgLFmr0GfcP2r+hYuT9ejhos5
GxxGQUKvdpInEjVpq8kpfR5twR3EZsnR4iaiy17bg9zov/prewbk0gAwE0NpJfhK
uxKINagzrTTHbHPQ0dLWaLvuoeOTnnpJlVqqKU5Wk1rnpDAeF5OeNqMc268YTwYj
YYq0KZFSrE4MUwXX0P7gZEd93JJBcJatDo6RKQ+lutmHIZea6uCG6nR112UYEOJH
q6f87XnPpwHdk2pZa0G4BhllLcjMWJWEQfefZbV7DZwGlggNtLP4+P/fzDUMyUck
c7RrWh4pxq0+yTEdHdvqocK/qUD7l6uNWHvY4nSRxNIuOGe//9MzwnJzb6LJYZ2y
7dPHzyXUJUL5JzpOx0v5gIIjc1h0OgiSqrfUrzlwXiSoAKZjT79AvP9wW7HY3eNy
sMx8vMfWDHa//mlo091OoRevj1clfnDS6hrg2ffA+SAH8FXBoxkPmDbnREW+rNKg
o1HNONsKceSZZ7dKNRRkE4cv8qjuSnLTnfqHSf9WDLGvSXvaHEeU+jWEP0Gg/kHr
own7Z0rXLMAbXNsDK2BzndcTlOWOLDmyOzxV7H0X0hgEgA2IMV/krWzKRem86VPM
e+bYmPXQMaKRbeBaWAhoC0/2vfnPQppJSt8MHCRUYPr53NRu939q8sMXGEKvXYyW
DW2tdvfOd90kwD1UAvk1hPHnWBc9siTqNe/Keg97eyYQr8CrKLujAnjryygko0qQ
CcPLZ6mwm1qFyuYlNUrvVPHRPu6gTanGIOy8xz2x5gkt5zFXBHqFY0ydKkIUIf1o
ndnALAWioOYl5isSF8DfQ7vc9wjDiFs4TBN1SxV7OlmIl7rmfSIauv9SjT+pc+LP
fntLlvZq+G2HVP13slkOYdcsYfSB/zfeiOAnBupr4fFarzae307j84wi9pef1Hpr
orUrunMfn7AzwEOUa1UtnjHG+l2pDhtcDFhp7c02zVrn3DDYfVsR2YqNa2xlOsVH
RmjWipHNHoXhh5WMCcNMeynqOy7SRUE/35yIZrMBasEF9Ag/58G1TQMsZYxsPye5
eMw4RR42YnOgHyw4KM87gChGvYnmchc1/UH6bIY87NfJyvI0N1rrPf3OLJwVVAl8
1kyhxLsPqnKGf5Pz2r3BqpYQJoi803OrYWZajx9ClzfhSyiCEfbIMCyxK8Dwik7G
8k2sGXAQNisLzJox5QifyJPaZEGahyCdtRLGG3hzZX7c8fYXPvzRaxKKGSGo3nWJ
OdsJiDTuBYK+gtC86H85zkRXqsMnCAZYdVWza5QjQ5anZu271RdLUs7U16nF+h8E
1huw2hkreItaHm9sUAqXsifQhPhDPgXz1Tf5uLMHfBSu8ZC2gv9IpDzXmGrtvP3n
WaoRRfM1hwmIJgw1jHm64+8rOAitnXeUybpOG53xKA1jvLMB7KLNDIrSm3P+rkM7
jHWHpzqVfCYk5Y7IoDcBsAKQBl5AI2T+DAbgI5AclsZU7nhLmwMNFgwyE1AjC8C2
+Xz8mvPcLYthIqjeX8NJZU+Ju59YEDXFcQRQP1wj4S5btrNwq4z3+d3rQNUgELRD
Zjpr/BEpo+iy5VolzjHw3guyN/Cm37jZbPMhzjXeDj6t8X8b38zdBqG2rPhOfs04
274nL3U0llXT+Fg8NHrxZCNFiLmkhXLO21f+M2xMewbYRsHv5CbiSsHnjEK8hxbg
y4FtmU6ZdruJ8uou+rsGecNHkBK7sVMP8u3hd7/kLxXNCDcSeWFZLtvlimezRMQ/
6vMG+jQiMhUrprQe0x7IcEqtiD8jDJKHSrGjxmnJpjJaD0sK2hmLuWsp+692JlXM
Godd6cW4nDx+kpQS5AjgJ7PCT4kIxNI2tUu/vF/oE5bVbLas0ZlB4xdBiA+hTRd6
stwFC4eheCtU/1ktt/W6kXe5xHEK57Pe9u06vzPGUPVoQHmHy7XuGxnCShsMScaV
SxhF2TAC4Btu5DTkswMNWN+z9YRHswKAWMukJToS+Bwr1F1qGVsZmmAGqV3tAKHx
8NgGg/bEQzh+VUXbAMt5jlJxdrUaVxfDkTgHHfea5j0lBhFMUbj2JnU6qGGJ460Y
NY43f7e7MHYIXy7DfWZQJPo2gGnK5IGlLsnNP+HckJxdkyTwCvm2zSUMTWodMb8H
zEDWZx1fOp1Nug5/8AjQu+96vEIGs7wo2+OgX4wLmTEwDw93ESXS8QfEfzf+d1fL
uGlcEwdI01jJ0xDlZIrdkVov+xyuYGew0NsBlMoqQS1NSPJrn/74ti1Z+Yriv1oK
v+DEdtO7OTFxuoRjbiofJ68N/niGBBHQZDOn6wZibBDVvihdJcluCIZsRJCGSyTw
FDjhZgE8Q9+GfzH0NcTJSCHdcehUjrOT9whV8piEOE2Bt2HODrBEM92xfKH+A3G5
cJKUUbjb7vdW/9FtW4AaLF5rv1ZAZaFwGjZ4W6QPu5fP9HhBtOnsrxORRygww0ZM
y20HnXZybRUAQ7DRjD1GmpQ2meTUtA3MjoicA35z8PQ=
`protect END_PROTECTED
