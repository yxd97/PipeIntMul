`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uj+bMcYdFJbDxRi/qfjthon0CKshTf+ZGemjMZ7YbDKy6Lo3BN2Ba0M2VwPWAhOc
Mg6sYLWsBFDynTKSSZrfYdPMTUTI9z+X5n/H4R+0QGRRk+vHyaaUfIYKU9yiMMuy
oo3Wzh9eYb1Em2C/7WTTiI4sVjVFQUkzJQkRlNh1uAaB7KTtykk0hdQv8FGcKxNa
UOG71XdEGEt7pGK4lCcK0yLWxJ6xg16Mb5CLEc/sSOueEJG5fvYRovCnYeoN8C3y
NVPhIKPN9J1LrANS7HnrjIume47BQkxcR7XHtONj5SXFc15Kijteg826jiZKA0zC
VLLYPCSGPWJjOsA9lcP1EplYw8VkRpcF8Ksd798h4gJFTLMyNWOZtBjqgl6Nmjww
zD0ZjqQSF1vGTHJ7rlRuVhYbXZXcR+HZJ6X14K6otFVXbo1lkfJU4OwwMktdMzTH
hkgo1pv66iVFKfzAZpSmkg+aXQ4lnCkAT75yIFIxkvB40kyLmhdOHgptLI7PrbrB
lIUyRKPP1g5vH/fAaEgVHnxGxtvcg4XShLkA5NE066gdcsestvmXi20NwEhsmBdC
NVLTIUdzQxe/fK3NorHsLTTSkTCLF1sZDLioAUbTh8FCwoumpLTT6n5ZoAYM/t0o
X8dS+0UIzq9Cx0xPIZYhOnnJ5RrrC51wftdi55jByhayCVetg7y+1tMEnxk3SlAv
6n4kuMYAB/9iZPqcXd5ZKO/pZ2sMTD+SkfeN3E+2vLJADCmrph8pgpLusG0QnHcr
ieyaUekE8Pua3xL93H6eKLkNyZs9ygIASV5NZGR0oylpVJBDFKjXe7pPQyay2CFn
VsVC90MhfW0a2on3uzswEg==
`protect END_PROTECTED
