`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8nWoaN1LNtP1aaqW5ua/thexcRPAL/o+nEQE/ohy2Cjz0elYEMtvnHa+WFatzM2
sSh1N25IS0ielkUe79UXuitFnw2KpjmwM6RmahxzQ8l/p9i1txvXNsg657t5lFNf
MFBj4BdJsYDPZRLcQRqWhA7JFth3QIWaEezcGNW6DC1d209XrxXuvkJkMrJLeIfA
BL/VMapetO+RztwJJLwZeq2qtzes07y/FsLdKaKpRBiwEmi11rxl+sQf5QXxnkHL
vR4roolgqwrLrOT7J9JtLipJcazkOyl0KA9BHrQF1/b7qNc+wjKf86FNIBCaPrrc
fW7KvdxlSOWNtzeImmcx7A==
`protect END_PROTECTED
