`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dd1stu1qhTxDffNyOp6ceof/ePCiEVHRG5W56ZTcHIyufsWUKbC8KDxFuSWDFMW9
zwjjKte3fONqya9+KqTTBVJmiIfGadiKbStUs4neUCXwyLBpnhrgk/mDS3DbSLRm
CAPA/7wglqR/L5sS/W+++uoSdaQ20NB/eUQNqBhOUOMHAHPYG6RfJPxzd2dnHRkV
YdRjPDI+aLPeXzdrscSKibRlxpkedqVXhXr+aSAK98YmEu78Bl3bamORyCZzzwVX
gczNSyNknyUOuhoQK/JBdpU7IPWlqFwe+j4yHg74GJwZOslZV04OpuDDAYx2f5vx
HW/TOWO/EaEnzgx8S/AOT2Wdoyu/eAlInkaw35org7hCVLflwCO9pFr03dooCAH3
3HM6OXQZsp5zm8ulWH0BuCItggaojAhe2+eOZpSuLAZgLH1DuXjt6HI5VQNaAa8S
03XtiI9Pqoigl2KRhchmhQKMfuL3ExvDzWxXCALpXu8=
`protect END_PROTECTED
