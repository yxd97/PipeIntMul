`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFL/L5KLo8cdoo0TXP1QRbegS4u2JkZfFLFq3FCdEb6azXY/CdIpZGhVh3xqD2TR
YnT/D2LDLzSJTMU9SeOOHI8QdmpIMhKE43TWQsrzMhnoZDBAyt3Sd9ctHhdtsqBw
wsAKNoIk2HbDeKmprYBQkvTe1eLY0LxaBGNj/t/t+rzDujNhWaZ7NJjPnB1L/ETm
OYFefIwAT26cx1cX3P1Yy5trgi92fUCsqWH6VeuocvyWpsp2wXGRNNwd+WRKRYtg
60j4Nu/g82TUxmnLHG4cIkiKhXraQT+4ZuTrUw8XXZrL6bZZVRq/qPCBXi+s0ZIQ
8TrydBHOHZJJpeZzMO/0ocvq1YU8Vi7OzZblSTTpw73nvq+c66guvoEGD0+LugPc
vkIa8UYzGLt1iunWU1EsPT3n6R/mM1fYVT4olkqhijAvVbDFvI1iDuyit4DHmRD+
cFfaDfyJiTlGpucVxWoPb17JDOB1oAUXWqLY5o8GDV34MjekCvCgR08dOUwkF6yD
`protect END_PROTECTED
