`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0uGQLb0aGCOKQysgU16E1naInmDOUDQVDD6ORcTYgtYNlZRE9e0DBDfXUPuVF3C
y9RuDM/9IaIga3kGurNGOzw8nh2ElbOpfY91eTmjRy1U2lGpiB9506t9Kyrl1jA0
dA4CTL8ghSJ8HrLSnWX6FAmnUCtmTEr/5cvdGWecNX/Vz7zo+sJdOANifbTPMGVL
xw0PEwBgdFwl3wz4GuWw36xjOw1Kfeh+mjhqHWBd5TFWm64P/hrhtSE0pDk/1K+R
E3g3jVR79HfPROfpIK6dn+ccIVFQfEyIgmnSiTsh7Vc=
`protect END_PROTECTED
