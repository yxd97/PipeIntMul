`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ED8aAsJyyh0c6Lf2w9xDvsdWCKC4clURgHxjQkr+9knFzDWF5wPZJDOC8kM2nMoW
7ZHT4iakXz4w979/YPNjJ+PAFEpqP0sXhtkKtZExiEtIZGDySAqAriWn5Z6rJepN
T6hOE58lR37EJvCr1nhqmmVh63bGxB0xJUSvjuGrYRkMo+7ObQqn8ATaZEg8IDv+
ZegVWhghKavRpLDFJCmx8pB+1aTiKYG0XpPEtaj51TTwcSAjMPWd0YxMTsvKPdPD
ltEtrxXbGB9anV9L6oqk1Fq4AVZB4XWTS9n+m6YijFwgnbLmN1V+A4M7XOIf2WAv
LeSMm/vJeCs5Z9bLflpTFNy+YLo5DPGMbiVX3di98TMxFpecLQO6D6shaok87WOg
`protect END_PROTECTED
