`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+tI5/l3i9Nu5yRVvdR6PONZ9f7edQSPwUyLbiMGB83aaJbXqTo5cPvRpAMcy48G
/1BC2iuswIhTcX2IFN4+sh0uQuNyFuJHC5X/NeT1P0th0Rs18oLv24FzRS7Ew08o
BHXEhlrU/sIehGrBAUiTkg7gv4CthAaWFSzHjb1hgbt0l1H8qUEVnKrI6S0SPob7
M8pis3Vt4c3QZ+MdGvgjG84n7qlOgVmG357M5RAxG4opY5k2EusLhVWOEOoQAc/K
q8jz/V8/5vIkuTOovQxEojsnvUzX82r9/ryvNwbIhkHGdWynAmAn/65sQ7SuYNzh
H9NP82pS8ewM1aHp/T8D/+lllUA6XLqDg2oamxwNcpLh8poYUjTqqQazPrq1ddWb
1O1uZVr9uMjJIFcXkbxOjqmOkyIrT6Vjw0MNXkxXyh9rbgzv7c9tcncYDoy1Xf37
remZx+3L6r+ezCkBWd4/AD3c4aWGPfCu/mUwaJIDuBfeSj3a7AdcALTWUBSLTSaL
ALFYZXEKIQAaorHPPESFng==
`protect END_PROTECTED
