`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHDkRhYYhsCikG31lK4dRbzhMSp9oua5+4fxOyYXcka1NsfJtlpzqvcasaJZf4iY
qFnlmWyty8TnzUDqr19mD0FtpCOrNys0CFnuOm6E+dzxHOJ3v/L8BDFn9EU4vitg
WibQ8mhXy/2Z6fAFlUBI2omRrT30PNzWk93PmdAJDXhoMwRhFOpiKZ98sksXqLFb
lFGDBfVcggbYz8oqPfLtieEgjo8doMrnHM1kVTUIhZwRdk4pda0rqDzj2D0Dh8Aw
OtRyBXQUBhf/H0OxHg8/+gqLFdmJAkr3m0bdE8NhOEtRoEvuRMEFNsUsTgH56K6X
KR819kZvLBnxNIVu6sSFI1W0xYKuRkfTDCfbIPv/zDRcQVa3tOnhnES6+Kn9yeu+
`protect END_PROTECTED
