`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3iY9J/3qJquAOsIt5ravpt93azK4F4gg3Ip72sH7vzRvpr6Ui8+vrdhR496K6E4X
By75XUtAx8Futtj4LnEHqomHZ999cKp7dCX07bAu+VTelwIROGWjbQk/ZDYJyHG0
EVzVwgf+egJYUwsEk1CBabNWCyIjhALiCa3BHyqcY8jyF4TYdnHzn1RCRRfb5/W6
WQjdYBjyTdLOHsUWdMeTZdW6F4Ku6ktbP7ptTdBskGxVnejQ6dzmIZLx/IhQidXH
CkWDhd8BOPgZEZXoAvwAmfz/XcMah5FJGbcyFl43aTGCrcWULeKunbuWCMj7LL83
CXJEGNiBPyZZUQtk8k9x3k7zril2G+FJAl5cjI3/UWj6tDuEcxGflIHs6nE6U2Mc
O94g9Wm0q+zy9Irba/vODW6Jtrtm5Yp++DFojkC5/1vU+6YgrF5vhInlIX39JsfV
PJLyVb2D10N6EuNLr+xWPdlMomwSV7ooKzaYGjygg4eVsiIapHhbG2FjsrkvwuOr
oPviTG4YjtmXPRTuD3dGDV27e18zj9gR7upAp9zvaa4rIRbUeIVYmTzSdDo4UKoI
/qPfMi0nOfvmBC1RXy7EZ9+UE5vi2nthb6CrIkjWQ4IXt9QqQJ6ikZM8Hg6zqfha
cGY2SHdkcFQZiY8haBcLkn061UWUkDqlwMMxbsqem0QJqIlPfPXIR+e0JBPT9pxX
ooQGjM6BVX7IuDPFVh1KyHhTVQBSNSP+eRVlynrpA9aNiRJhGlVExAw4XYe3CnEw
tWyrZVDxLhogJ8AjOKXgZA==
`protect END_PROTECTED
