`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzVq38++mdRqgXs9R8fO906k9gi8nsgTh3Av1H7vEa8QWeynEm1fk7BpIb7CikYn
glwQGEKykeXsaaBnmC9eBBeq9a5jvZUFoO/j/7ZD+GfIdiSM4fkHWyUHWnnmV3l/
/ihH3CNL7+3jrorfeZGaJ6b5WR+4JFGcrYKKlk8gakpQfBorBfCWHMMoMUPwx06m
6p9ypyFQQgI8UhXNRs7NJjg5+uZ8bCptvglhEqXWQ4uiX5G9uwfHLoSkFP6jnsP8
ORsnULONPJ++tMGFSpuEys0RwNab33dHahGkBGqG9Gjlx5VIj2D+IrCyMvUOZ6jg
Ok2xoio2bgVO+cqubNa/IA==
`protect END_PROTECTED
