`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NTPHpz+CPseJ2UruUDTkBbNfc1ComsWUzBpbs5qWHGZ32riRkOokuSMKyh1mlbrr
vKmsCO7d0emZM+CTej6Ocm1kVbWt3Ayr9UFsUmKJ9Qz5F7BRg3z88itYxNPT89Ol
Yncm2sbJGlgqCkLQ3tfwWDChpg6CVnTcru63S//wA9govFwd9PWH1VSOvBpIWaav
3FrKOuephhNcfP/15qNdxsE7W/NFycNJVCnoOHySShnVWdGrtwUdNs6fLH1KS+Bv
aK9YkvGUiK+kaI5dhd9cLgM91tAPsTCsbQ0HFJKFIlqQPfv0APpowHfJrp17xLbk
0dSqKb+JY0t5KWG/3ROfgHYjbCe1RxFwlD6Oosr+m61ya6p/3cssWZLcKNeTrm2x
N3owLgHw9wZK08susARfedup8BcaG7r5jAQ9TFf6jvvvqjcbIWURMghssuhzfweL
n7q6rb2+cTbo+bd7gYGxEY5q2V0v1TwbptecPG+pNgCzKA3kqU3DXjkhCSLkpk/E
1lGK0YcXM4JHV1kVp9rSXVzZeL0+EdYxg9Z9rc3guHGG9h2+t8g2N530WPzv9KsN
PM+9vStP7900icdQKNbEPQ==
`protect END_PROTECTED
