`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qja7j5DV8oNFRjI+KP82RlHkLdGwcpM/p5+AmCf3lbCTsMfnQ2we+Ee3O1K5ArtN
+9OvLkmvMMMDhrkXI3C6jf3P6v23d4/x/a5/vnugtJrXm3Pbo6LE39A0t4sEA7m3
UnLCGHzG+7OcySRyIHEBUETPV14tEeuHpPX4qX/hdbaO6hbKOfPgWdOZPmIT0XiO
LuDA6YSyozjghC22R6LLCDhBeYbWaQqMo8EVn/HcZ3hU4aWX5ZSln3phddds8dmI
`protect END_PROTECTED
