`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLp9OGjroBjGum5iebC0XZcEOsiaUADb5gn9W1IK+NMw4FY0y+2c4avseeFwJvti
wIgyqqwbjfoHxnfEWc7CRPfKHofcwMfKZpllXIMN9nCRd7g7MWpw26ZJZCPdUkNi
ag/S2neckAkL0FN04wKLQgtyOE82YKCz0O6Z9ms/zSfY+lZPxGq0HjpyiA1BDQ7U
sXtEr8iZkD/e2AUjkDyPVDTDzud/2K1Blg/ncZI8thN0NyGBn+X4SqjS5lOLcPbf
F/IQ4t1uIHCYaqGROhhogtrwKHGPqIJVGp6D25G6y/Ry/zay0vqgz7A56NvGpn6z
C3R8hEi4duFCoyvFHew49arrtVvtR6nDBOxyZ8b1RMOMRBX4QhaQkiO4gAGI4E81
Q6v8koATRz1WOLV/n2wooqAQB0Bm6rrNlQxzoDBAXAWzhDNz2CUfluFhEMly8VBK
moO/TRUD7qNNy80qNLSES4S1wkQp1GKbDnGvMSm5mKoE9gJCvUDb8zjZEz7BnGKc
vcLJ+qstnxUQhmogdvZKwcwQUk/TD6EZ9Xt5Sn0ePunccq2kfq0rs9SQGMsGzLYB
uKCRnACRF/ItalOe7ZigL2fkRtDC0I2BRwTNzJ97OQj75S13zcYkoQWPyOWD8enw
`protect END_PROTECTED
