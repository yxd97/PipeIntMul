`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0if7W+vgZOXpW/+eAzGoRfN+xgarVg72hiQOPghW/0bnIdPO3TGpejQDTG6WXK3e
CvhVh53zigEw/ux3EuOuRbjQpO3Ix9fGfEpFXlj7474sphJ3S3vo+4Sz5deon7lF
ja+M0MjffjKDVVPDeK0Oc9oL8Qzg5uhEtdbfnQDdxtcuekWB6VWvVM+0edMlGjuk
ahooq4g4tgtu5i/fNsZnwUuTaAkL5D4o1+1EWSIfsKUK6wowVdWus4Q/OgJ9ZrZ0
OInyBBQ81BdxhYDxtIZ630V7ThFBF9GCBkd0YQBzaMW8UlnLcZ5J4WN43W1FG2Ss
kXcR22Kyff1CLVS7EQL0uwuWvZlFPHXHRVo919lPE5iBopOnwwMaV7A3C3A/+sqj
WiQOwx7v/Y7TWuJdXz3eGk8peK8pbHIdWITn9IJMPQBrq8du0adksqC/Ix12Yfy8
uK/CNNBmEHNVpkzvbZ19uZKMSlv76jSQJfQnobC6QPz/aoGid8tZVFuHN8CYw81e
`protect END_PROTECTED
