`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2YEBD0bmuL0b+i+Um39FDxMUmr0vMTO7dSHPJstI1TelraNjJUQ624hQm38AOubM
pKTW05S0SuIvpfFuaMRV5W7rB8dYTMBYVpVYO1/KoquwPMtlp6MGuM4y+VTRzcer
U4XBVKcAqCJQgubFysPHoIzbIOsrFzaFeVBw8Rcqwyrdtm4uZi/BIapIZuaYtrA0
P2jIM+nSi1HmUlr3KMjTiAkvqK514oJenXIZE2kMveu3deR6aXL126a090VJQk51
dyxzoxtvsTdLH6oOnxBP2TW/HeHjXGQ6B0unykArpTi/r2WDbJzC95c2+g6y6a9e
2nmB391O2uZzxwOiUXzJ+iUShFZLihe7Q2MvpKOfkW565f8oJ9EKDwWCCwkhrVBW
uxJK1yS7S8skbn7aYzNIdNMdpsj+joMzWZ2jngP7piRzcHkDmWIcwI644Uley/w+
Fb1xRSoP36rHaDSiMQy32T5ro0DpFNETxaO/CPxQzPwfd2wqxRLEeg6i04kyVE2A
iBdrszb5kzT0NX2Q4mVk3P9O9GlDd2Tx8//Pz02IU0QIvbvtxGzMcSfjb8nmzZkP
`protect END_PROTECTED
