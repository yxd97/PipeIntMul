`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDGr5ZVP0xxvflPN50vXDZ2EE6XYoRtN3mHDG/AqQm6K9ZGjKTWb7GOiMCTXqSYk
kZsnxrYdUIATzcmDJsJwzWZ/uFCaiCx3yEGQAGsM4Cm3TOG+27CWaRSslQr4OO/+
LYcv6LQPgl2jdKKdCaYMi5f829rK1fYcd8HIf+OM8WS3CqFx5n3N7spMs9sIwnVn
NGjVKNM/6dKSZh3C7+UOKzstPAzBC9KDUuPPM6UHXHip3p6A2pXq3fPPClyqc9P2
xwCLnRymj2cLZhY0l2WgmrEKKg0kyP+UwYobAT5c50uHt8cbHEPiIAYpJrdm6sV5
wg51eriqQyuvwYEG4Zib8A==
`protect END_PROTECTED
