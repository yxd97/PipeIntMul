`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/UgnvJyy7RSmxpS3sW5dsDeNw3fdetHvXlq/leu5oLhUcKoztMaiHrDAr84qGX9f
qNa5AJdd9wCImINq1yNNz6d3jD/ldBut6CB7j4Ot0QaBarPdiMrHtN8EsPUIMq8N
yVHS/2Pmbe3/3MNxBlVn7nABAlC+6003UrlT+tXw/7UHsz37e9+PtM5GGHIffnL2
VVOoCPGb4ibES2EV3xpkQzij+6RDRVmOfhWv3a4YkESeVsjelaA9GeH4shvAtFeP
AffJUJ39x5o3xGKEF9eh6lzflQxJOwY5vqJ7zvHJjW7k+pR7kaOjV+qj3zwpUQus
uLnG1C+Jrtin783IrU0WFPVKiSC4eDG9UY6vmNwOU7vQNkAe6sSZIMsZ6rVyHV8S
VEWDmMz58wVm2EIg2jorJarsLY5Us/qPr2JLyqjcVUQ6T3ibpzW1ZE1Y/XTECUXm
BkfqTATzkjBSGsn9GE9kM4pWV8w7iipkYeWDigJS0ERcbB5i3OKKLYzJjOP1qFQ7
L9KoU5BJQBKu5gWkVrU0g5c/7kt2pID/5rHuRGqhr+yTe7safEhdMhcfaJhK/bpx
`protect END_PROTECTED
