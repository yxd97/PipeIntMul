`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oQRZVZ8BoZe/gg49TWK6o1yPfKKioJTsTZBtMNOlcba44S2jN87ZVaoCYcaWwFXW
h5vG64htDyESwZNmh7PD2D+nJfERHiDHyj7CPjpSZSWxEfzTV+vR9jocxuLPaHYn
0l4A0n7WMTLZNJzOZDr8h4VvYD2+BC1sNnHy9lobBbFqB7ja2J1acR79HJS/qq0G
U4CwGTH4Kxc2YtHT3TPzeUdipisMJ08aajOmlE+7xz6dgHNeH8x9PYLKqjRSTgZq
PWfLNwpsxbwRzI5ZOK9iaNAR3a3h7QffyzihJph2W6/7++fOOiX8hZkGd39vIDy1
92MJzHSc9/anpQfpAF0zBs6MsP9GBjKpDqZrmVovyOGqdLACe9N1e7bVe3noGJ97
E3bezOxn/rHq3rwXsTZ3Ti20BhBEs+w8ONVzeuz4bleYP4GYbXJ+yThJepBcMB2N
`protect END_PROTECTED
