`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n9VgbjHU65gUaZJ2vyTWY4H/y/z8DsS4nAhc0+hptMht2xu2vPLS6gU01TVNCS6q
NpoBs6M7gefvKxCLNjvt901jGaIJZDpjv1hwn/s6RcexrxA92aowulEj2TrnKsJQ
d7xH/jmjvkmDFHV0KtYNMPbBJ+1+/F7dK42gE0iC7qzJH8AK8O8/YEgxsfRlz82k
DajoB8jR+j8g1A8HoFcdTdBpPv2eKsTOj/LyTOrSPGOftIJhmgrYxuHGZra2jPXn
h5Uzh40xseCJR7qk4xe/81sFzBSEIT8VfP0tsNClmvx8YHmpDSNT44iqwFt+atct
tctVjV1qyt6q9rnMcJ26GA+IDXYl3c7XhTjDR3xBjdn++bdY/Ic58dUmAGF+zBRJ
w+/sqRpjVQdq8YbLPB9Nzmc12LmJn7QNYpPumZbS8LA=
`protect END_PROTECTED
