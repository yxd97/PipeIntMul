`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bxG/o9syH4ZAZQIS1YRzwLbaKva7L2DLa2ghtDW9ySIRPucj/bRcxw16GKYOMiT0
q0/PfdkHnkUuMeIDkN7NAry03xtl8zeqdKFwJBdGI6soueYrfSlsk9PlxomC8+7/
Vyh/DHjX5wrJGsmzlqqUDBjAkSzKhibbxnCChVRa27Z8YAQwAMRRKuKI6z6Gcggy
b9dAOdZhAgJiR66xHQhLcNkdt0MfujneWmcFp8BAqSrrBiXhvJvjr0gpydo20M0u
mH6+k86l1vX1GcunrUqc1bSjfJbx52QP50JuGuxI+0arVe9EM0/IqPiUWCF4PRDl
aQyLnE8kDCL+XWZHSMMCcddZ6UXoFNVoO4Z0Y6wMO47Q3ffuVjWM7pUvcx1Llien
`protect END_PROTECTED
