`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qfyg2snuC8NuFnyXoVnMqb2zJezzwyTiW/2ejFTyuPkK3a0iTV5JEUbheTaCN6y1
ZrOohVnK0dsxhLm7lJe/evRVJxFRNXm7SQhBXvUsifbIX2z3FMjhL0wlukZVIlIV
S2AI+WO79rMEzY9v8RiQZzbhAsOIvu5gSpNL87LU2opu+bijJeSeLuve3CN9cOvL
w+YUHRQuRaWY15CbpWprII1wEoJm5NcIreWwJrGReWRe5oNgnBjSe5jA2/Syf5oX
QuCrZJ+kG/CAqlJO9c/5qoDq1Xtdnx0QqYbI1gJ5VLwEeg1tDyPLcMjOgDtElWG1
R/kwFd63gwTq0hASmKapCKbAM5eWbiGflRs8L7Qg80E=
`protect END_PROTECTED
