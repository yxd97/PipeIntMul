`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/R2IKJYNssj2L9AOxYYePbaO290RJSZiDfJkvxhE2vJLBnf70xNt3bcDY3Gw1CnW
lcjMtQ/Bv5xk5/HB+lPFmITqHHge9CV8pqT4im6jA7tRFrEJnEWh7Vp2EQN0KSoG
Uyi/FJGxYAqYgA+FlF+MaMf3b0GNBhzqBXw4xq39E3y4C2ig9BYyXeesGCqlBrUa
HpRHhCPufjKaO60R1CoX+va8cUCqt91vb8IfTqqEKYlpJcSUDmuedYgwcpMr+LHm
ZvDuL/+B/qDhKSV2yNNLn0Whh3wUisWNlfDfzs2vO7ygUtOuwXkEfjsflp4HU6aK
M6zOg/2a9+PEVB56ydynR853RgC8GQLGp3+N36CcBQwcBxBgTqIy0D743edAdKfz
P6TWwXGJe3QnGPnLIKnHLBBj+stD6srBO/M6hekVUhjACmn1SyLPEBwQNQIYh4/h
`protect END_PROTECTED
