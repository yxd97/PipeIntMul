`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3t9kTaxYyMM49GnV0OExynM3NwTyNc2B1ogBQYgbqUmBoU3mPZifDWFJPx3E0Gy
SEi7BOn7rte9gd2xWbheGbd+Jv1wHE6ZRvGWtf1P/X2R8o2KTgVGIJrFkKgRYFrE
e983NJs/ES36Nphjy1vBt8oxyyiWVKGhXxRQWmsD/8+ck0Irr9yBxhbr6ZYET26c
U+DWT+J8Esgl9rUTsaLisEJv/NwVIOR04lEEjegx0buGts3AEyHjIkhVv/6qN4OI
vIjcjG6U5S5FZu+dHNdj1Xu8RBCfOYnxdH8QZ3pLQsMxUAZevo8/cVQqGNj/XrSJ
R75lXpcXbVxBe++ehaDZUqFPdKPhfAi/byHV/V/mmoAgfmp+7agMR4E35sNH6iST
SuaASlTeP7iQZ4T1Q1jq2H2uQ3cPRyYkdeEb2Eb9hDd+uzysvPsvh8U5dL3Xz2fq
IlGXJ2kr8L4PituyYDLO9ms5gY50HibfmkzjW7njQmLeMPHSz5ZtwxZKOi5jLpcK
eGPN7GDl6YL/+nxSAFrSbGNMqsFN70gLVquQFyG+IvLbrqzlkNPqTUvR4PY4htiy
yvV1n9LAg4gZq29KGzgOGmqcwAc2uRdf9ShfMYIQ9Rmh4niaQ5Cg2tbFH1VIPmQz
jDwbkttyq5tzd6HrbYTVODG36ygv2Tc5MKWaAGgeBgoulH46PG19TjHHlDI8yM0B
3IW73Xf4X7t9KVWhP/+x0ayiNpuaOx20iKiXNgPlDMCnZcdVsfDOY31V+dygdqXT
7psvFDzUz03skxzJwCLBn4jDwWKpZKsBZl+zgGaeJMxhCf9jAkhOvURPb0PYitVo
Vq1GUwCq9YtisewhsmdiFskEM40KHdqnP8IT8mHSJL4m+FZ1sujonlD1nCYOSpEY
v/oSFLWbT0GBd0kqN0qpL1KyRy2x3ts05SsTcvXmRT304xVsSyV70gDLZU8iux57
+9WbOrrpn0Pr4FkD/SF7XRbITGUy2Z2kFwRfIHG/GEgZZXFtMBhYn99mGFCbcE8T
yPjX5ckEpsRneNMNSP0bQrZsRlz1eOfsjIPapgEtxyswiS8sd0zfj5thdZ/1E6wh
k0VQUS24cgwk6C/n82mEwhIDrpljqr2TefcLXAwG/1OHNnuFWkGHc2EORfIAOu4V
JCKvhXZW7k4GyFXHwlk1rl+WMFNkI3Kk4F+Av7gc++xADhAZTpiwhnLSPqM8NAjl
+ecxK8S3o3v/yq86itZK7yvBIUGles94sKSRto7iMTVfzufTKibgzPnk/LNnOj//
p4Z3l8QXpCwyoUZtKeBYwJrvr54YWxTg5vPBaGmsO3HZxPjkqIBaJY2zRKwDAkis
J/PwhqsR5L+NVqqR1GrdAB4IlDRcAgbIQN3bH9BJs94R9rMLB6ZiiCtRyMMWDNUH
cK6ybUoJioQYgczxInxv6ttJlNOlghKXHmWSfqeyMHxnmVSO+xBr6LwG8CIBKi/A
bcpPTemTC5TUlx8XH2l//lmveQqCmOQxp+YhWACmieqPtgHKeAx/BjBUXOk9snaO
hiX55y3ek9GmbpTI0GTB5zTls63J3bO+j6kYLZNnW96RSDaedJUIbk9nuvP15+hE
ZY7wscalwC7ZxfAxSEUug8G59jQIrP9GneJW1Zl2soI6aS3Tl57ZXQmXlVfC9tE0
N2YSkx4JQ1aIoJBitLv7Ybr+6nRXrXh5nRxp8VV00F6E9eraoAXZsESR8Hr+xXCR
A4q+UtGibbyNbJILMqDX+EDl9TWrGTqINM8Fcn4litwS66wZF8bOziKAmtCzJD34
DCJBC0FU7G3loVct+MSvVvDlGhxViyMH/AO3b/VEZ2s52e1i7nZKUy9SEwrhbrbM
lSvzVBQZ3od7Z3rZVT/R7V4FPejjgVEhUybc22LW+AWrJEInf5BZzoadW86JJnYg
zn87h/9vSGGSxz+x7ShtZ4N4DUfunrSwxG3/0Q2RxkgUI+rteo4436NNO3HpfU9b
6HZ2aH8ZtOgnFae6xzSC8oUGNxQrhWyZmj9FZWtvf2Nl0Lb4JgsjmD4OVdNzUF0J
WawSMvU6OsoE+adtS6+PFE8reNqy9d6kw31pJRDFPL7m5eoxAzp77Sa7z0kULjQr
VZWFcGe/fw3yBASj9NEXVOXdEbMoUz6hctLMxQSw3d4j93nhJeYNUFvzupOKaHog
R2K1nhxFDzDt3Qo42jl5ktprseWi1KWnAuPL30BV6JB5XdnHbc61R319RDEZ7VzB
goeYPlzjh8jl36LbuFlrKHeePIEiWcwt04nCf+hlWobbtcy/o8o+YMDuJd+S3AmT
BXXvBD9nvXow47Lr21j/tzGlM479IV+OL04tqSR2EdwpeVLgYBeNb35cYIY4TO9o
CvcO3kTC49xzewVEaxCz3LEpv7MlDwulRMo8vLE7f+WbhSwTmUpUEN2EX3Q0wnCn
l3c0yVJC//MBeVV0yHX3xSu5pA8HnlRybNEYGf+Lxk4Jw1JaPP7IuflEZbpNGOPJ
OhHa4XdmFoT6VtommzeDBPzsLLq+X4YRUGPb+WXqLpJYGbi2KK8c9t46PxwAvg+9
eYm+UldHAJKjod9hb8DJTmONLAYaZRi0lSN4oZZYpKdqw8Rvfyq1aJnghxllYkoQ
7Sow/QBt2oXhNGE0lG2593iyPsQJLaAADe/UTxdYTuu0S4agGonQfV5BUQ9pfZsT
5xbunlweygu74l/09gNm7ly9eiUFdjLGV1jNqOTvOm7QwOEAKzXjc6OvOjfJDfzR
KQF2cBtl1FohSiHiGiNnJuD8M9/zQ5n9qZ0O07pb1DomSTx+Sqw0aBsC4pnH8mkf
KOqCq9mju+Uyfe4N++HeTFOYnEZ8V3fL7pM44Vvk344Q8yGlWEqlzqAGxMsQU2O0
y/XbZi+9fcUuL0HUhYCFrsdsAOVvoMIaTFvupuatbvk8xe1axB5PmTZUaHVM95q/
AS73g+UqioT4zIa3/NHowiy19envdwsNPcqI7cZ1HIa/xzfto/JVKt9bJlUR5tiV
EuWzWysBZs1kMYuDDOoNfgIqluhk4dtki5kEFfU9oPBqtKu1boTASCvjS4/Gm/ji
bp8bTr9I+7pG7wzfcsSyTCAYc8ht6Re/TlKKw2Ck46fIxoQbhlY5m7WUfxCDnq3T
O5YHTr5tcx8BTe4fj2K2+vImsfHHwCTqI8BfKW81BpG6S4SuCTzEgjFvZtCH/+6Z
UdaFsOUYlltHkY01l9Mz7bxxq4Zh6VTSM7D16WwkygFTQuyk9Utl1kBlh5cKxH5T
D+4Y1DanagI4NLPJ0od2cNetMc1EgGr8/jNAzM+HQm9fXtY2XQKRYJ18qwOnIjXl
Ito0olYNnzhNkol3KhlY+KkXUYYWcl9wyY65kXK3UAMM7JDSExCkHpBGl3oslNFz
YSa4n8bgYDHVFv+onqmw1207CSLcRfqAPVsMVhA8aBKbvtIXYZDSa01E/LbKZ03d
hR8f9Q1nKi04e0IjAfA01feHQPZoBiSKcMoMTTJ0niCvwkyJHHzjIElsfKySr4c3
zl/rG1R7gS60XpglTExHEpdg1/+22ayeWLoYj6glf5wPpbB4NkCwMoY+CnojeLpB
mKmZ1xtyCW3FsQyhppwvH23I8rPbEyAZEcfp7Efv3I5c1vcQ4sd4j3akjHhLqkcS
GDBW3YU35N2p4Qmh13lejG11Gv4nSaxBOciPu5ou+ewbVJ7kXD+tUxQaV/YEOddV
uRPtsgCs3JWkg62jGPMLeBBuuFdvm+sPeuF5Ylx77EuGyrR2LI1l1W1G83N3INpq
xR7JRYLsHCOFdnwW0ZhEv6r7qMZnhH6lepCH6T6GO3eMIM4CBs9QXUmID3sMkla4
E2VQ3L1IU6c5aufkr0ET3b0HKivS6qIFg/n3lY5x6yR/W/ZmZgPyCAHixqIDD6Gj
tlMnubit2YqC2Q27+HwlAE9hsjACHfg9+C1BJVB+dJclBvZ2CCRF4GIrJXyeAtU0
B6/+ER0mDmJL6eRaoB+NqCTOc1OwT34Mz7UczUkRK1hNhn0jT1v4hvwia2tAUmsw
SJR772bBXkO2FbGX4nHTB6NZEx5h+KmoM5tQEd51XLYasFsh1ytGifgdxZ3//oxN
i9Zi1gISUc1XJTw3docjaLKt9NgXYh9gyde1l01NVSJD2CsLHnqK4THjNdPP1oR1
tc9g2C1yob+9Iu18HWAtJG1J8s4uNUXkceAYqzzwdz/FR6jE2VgjydIaAjzuRD7D
2X9FqfkDc4WeaT4oRcFOjwZ1YqxNcDsj5hKLnuomhwEzKUvxuUuicM9gzQogKK0g
ppmwFmaPAppJ4HN8M3Ssduqrvr1Ns88c7K02Jn/PjlKeJzKAw4h+X+AfdDIn+fyr
d1Ng3fVFHQHOOAe2g3YiP6T7wNlDEQfaimWoTHM3N8Zmi/Z41t7g3IcTc3KjqUQh
Xh13BjpWswKuESycTEW08kOGdDIag9NL0J3DgCUwyad53rt1pcGBG5XQnBdIEw/J
YU2fmoyJarP+O7NNndpS8XjHiaTYYXxKtRbxn4gJXuNGb6yV53h1c3d+wcOwcBnZ
lCLMmgqWgCuexZj23TfRbLimnr9GKhqgJi1mIyGKLishmT5sNRKBar/cUU7hVh31
DqzrA4fP8sxycw3zIF48ynWPaweTF0AOFC9QOlVcuTNJC42thj/inyMYIDMoVq5J
3ZM+SVVpy5+xjk0QSrbP8f9cgIoDCAAUTJj3ngnDJ0jZsNWfUIB0kYYlvpaB3vzX
c8fZTzXNflcRWRZOWsSGjIJ74U+xZYroH5UVe0n3dgB+gVMWnhwJ3O4956BNVAl1
3LCJgKIx9pj+0YqM6QC7g4hnj/x3/Jvq2ed3P4hJnpcUp0HYayY4HGI3b23fwMI+
1jIWg5h3WeGZb3gkPfi3E+YvC6grbV3/ltuZ3nZWGJCAwPw3ZhqAvW5Wipg8aywR
37/aC9cnGctPeU0mp/NZxC+yGtlQQWS53oLvxRJGGQNpT7yhBVcntF9Qtunt17mj
H+Nd4umj0QMOxRHnNohR8UJlA9+1a4yAdgFrVK5R+gqNJwS4bdo9Tmzrh+HuGQV9
N/M1UEhd13cbkAtWF6QRCyUnglQcRJDSRnOo46f5akvWgRJ+dOqJ5ZGlm36LJsDJ
Z23kt3HFg6v/CctmGZDTyiHkI/OGBTOzBviQ6tn5yM2ShGtRrLU51GqZLYSm1T4d
X9I22uf0RgKJg1ClWDhifg==
`protect END_PROTECTED
