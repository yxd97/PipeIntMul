`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YItLDhOIBSF9oeqe+FQASLrHmzZLVMIXOTDQ8uXQBoPX8FoTSRbg7GmroowZ5u4V
7vVPR6DBIHj/PFquH0inuUPj/84oUKDwze7T36O3RrOtZ3Up4TMiYOCrboFUUqH/
CTpjh27WY7THxOQAb+rzXHYWDe+L88jWoseshm5oQc7hC6/sHBZcbmqMlgDiKTZ5
mDflFk0ldCzDc9OxfzMhTa7y45Q7yRcJ+dtgknmf+bbxoXw1V2OrDMmKqEOi90fl
8k2kYoGqGl30ugrOhH2jTCQwOJn49ucBerxxgFUJ16Wj6Ae9ZRVPeONsjEtcE/RA
BYRrwTbr8oA/P6d75dEFQWd76s4XkK4LMLZ+uDJ67Z7+4hQCr6iCEI0SZqwpCTDh
7UF0kP+5QfsfB5MQJCNzNT0h0xKf6YGeU5IE0OUsW8M3DgScBOWdL5TrCMIMvbJq
Ey0bYmzDUjQsfoNryZK34J8ZUUrCYSjBV2Vx9JCbJ6kYGSHmbTtOhbIf4Gt/rfGG
CvlBQPW1nSYO7D6JYdzVtTmVBd/rc6nq3MO1WZ5NMEJZkYnSqzUFa5HsAUfTlXjL
rbe4oNLlWhuMrMEmEIbhenRJIO2f3/EqU85LeEacQlHugvKANWSWXvhktcwSX7vF
k6DKRAcXN+IjjXHZviobzA/qE0kG+51d+uj0ji0EXCqeD566HjtaX6IFoLdBoXq/
Qd/ZVLt79VnGiPs87QqaqKaRfIYT+TYTjGJ83P5tRTZboJvTGvNYjrLfDn+6jYcQ
86avkqerEeWKz5urhNellLCzmBB3HP9+n0cyiq/Epcg=
`protect END_PROTECTED
