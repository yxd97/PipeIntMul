`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JwvVgFa2wvQ2vOm3vx+l8bRwCgdC3ogjJKs2zhl8WcrKT5MTyxIyEZEcqKgj5llZ
v6magiGfxgUvw3ZVH6gXHECBa+kUHAIHZ8tuZGDI+FMDC8P4VcMAiGL153OX0YFa
ZKbzze7XoExfEoYChje0fQ5wzEnGZTLZY2Sm7AjVF49QPQ6t6j3xsGj8SMvd2fs+
2GgVj+tIL01Z43hRSpo+PB3ua45aFQazoVSbsPrkSlyH+pOA4+Pk0S4vlK6WB9rG
/fI0CdgceMzPrxYR+sq5HlM84nGYot24M6rs7ZBZg7BNnyLrlytbON14nVqdnKYS
U79u3LjSmb5XxCd0jpDS27qrdhpONhbwPOPkoGOwZfc5oDZMjGVynBHmFiBPf/5t
qqwLTX2SSAJGNLWPmazID9Xtev1kwRvtbj6gdBMGH+JP2Wvwgj8e3dILvESbbKml
jwF7joLt/XfdlA0XULSYDGOCnf2tAuuHPLmNxiHLv31GKl9SzsJk1z0TOtIE2IJs
HIO0dIi0WevC3Oi4jE+3mcHr2SzYIthNekFa/aXUX/wrIwD4VwE/UMME22UciUey
/nDsQ1ZQyxSOu6NbF/Un5jo1H/0INNkltoEcUhpk7RF4VUNS5un9gQkJ7M2+sOlk
LFGyXqhld3EDSKfaSy3m77HvCVQzH5KNHtLB/eqDJa149AWyor5VvotC4cOsg11g
Osm+Vw2OtoFikLbeDdioOKHWVZdMqHOPW30tkEnuqCneZvDIznx1htf4j/fWlYyk
9ycvPnRaLjWykvFBpzE9gKx9mgcnk1Mky71cEh87BU1pp6yfhZnpggyzDsj8nqKq
pKeNY6clPVugQFi1q42jWbBTiJSOw+oEMjexPoqIg9NrfjiJ3R3T2rTm4KYrFGum
Z7LnzzKoL1+lNe1559XsIiFWOb+tTPxTbhHVqLrTKb0pDGo4l/5Tbtb4L1/qG0Qu
Hn9E5h9gTR8/jzorp60RI4vCFnlsugQWFEevxlJqLHl+2tc090a9yZtig9dyxLBP
58dbyr5Khsx5+cDbmzHgJmDGL6c72pj4ulIy2npQy4t8h4LrIhtRd1rBz+NXHG3Z
XmRgr9Uvymw/9xCAIWbwmwcVNL+9UuwLH7UvUBSz7go9/XC/5W4gGE7/KibcQ+/m
HxOV727I34NuUZ/D2L2h+6sCQXaVLmGnT6FEmsXljdJSu/htMwvviCB1DnSyG8BL
5imN8gBJBhZw9lumSR7NlxyhBwRF7JPxcoHPJtB5u2EdEmP8iYomYgjCZiMzp2C1
jmivJrDdMNT/YbSnl8avncSmMNvUiKKptKs1Yy1YBKJGQwnR6GhLPiYDFtnQZnN1
`protect END_PROTECTED
