`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9nu1iVP5zWMOy3H2PBzHM2jEykKeOXMQA1kOh24/o2Yf2tP92U5Ryge9Jd8ts54s
Kfzo+3uto7ERQOXl8mez1uICjr885EE3vHr6LePjZGPzwTiuxz5rgZv8SP/iVwSD
eVpIu+puxLlqE4fVCoKHXI6bDhDosgPL74vY7hlARYxind/C3Su7lofXW2a10dOs
aEEhQi1B4ZhTSjdKeeeVZlvMW/wGxixG2tuwZPFq0qG5G5O/0TXP7MCYsstzdL11
qTeZ7EBWoxUVjqHx5cbEH19B8FzqqQqGXwYntNrKATXOHWi4XS/ltWnsOi6gIrxQ
MEhdia7hImxWEcifze+4ZCBC/K/qO+axjddDNO7dS96S3iQIEvZ+7tfS+ZlzQSIr
B8s5wWZjlSZW3rf/8kAUhYet80shJfqZeUzbWmgc6Oobob1I2bZgKFnBuykEy03q
`protect END_PROTECTED
