`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TMqOpd3cPv9WgjZJ5vbCsdceYwIyJ7wZt37cv2jRmq7XhEphwhsL+S1yBYmeuR1B
zX2G+2q87GGKUXda8DXlp5Ood885Ksh238f1TuEjLu2vpqAd/4kGsu7vcJrRFNPH
7E4SroY4eYASkRl0lkWHdZsvobiNuIvTo+Ve2hcUADTrsywqRZtNYUqlqqe9SjJW
Tcd3T4XVVFlUJjCk+LbrSI0jQ52kY3eswqxV+ziMhWgqiiw3SA5PicG1wbn14b1Q
FCsLLHQqK7mWCPuWfaQ4kdeS0hML7KHsu00nN+j8pQEZs7ofNGzVChkXV1Zq0Rzn
x7umUWa+daLxZq05NvjxJKVOWN0Cehnx8B9MT4l3DNLSO2yGe94qLKTmsrVnCym1
XzMtZD8BMy8fS4VUneH8ll3IEuPmMsVMc+y/1r7NFEVVddR+4Vw0aiV3EKvZy1YT
JLt2ZhzjBn77JIrmh6oUSlx/MHndSOPKfstJTeFodPIOCstaHqc5srEWpKY8m7CL
`protect END_PROTECTED
