`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fWaW+7J7XUSZVhWZ96gAOVg1Y82qgQ12ntf5RXoGwBx6MvYvbJsjE6O7YYA/yUP7
rmpAb71YmpdzVoKDh7BT4OnSziYamn1tYrgheLkwh/XZJxtiwmqKhc8OrDBJMXYE
u/Yw05oIdx6k5K+3oLhtuhPJ2CEysVMaggbvQ/6CmaPOSfkHlrFoxu4GxfJL60bo
Xbzbos2RCYhEDxdJBx+Xgers47GVSUi5k/FL3IvMJ9tpxZQEV8clC/JRp6wCUq+/
SEVtnme5sw1I5ZT717mTqD1gXb2ATCh+/s1vpEVlPRYtTInvflmBddPrVvctUPY7
nIPCIRJVFFmVv/21g1S9J1jG17gfe/9PbEioMn5X7dqH0mN4zif0WMIFdNf9N5Z2
mnFNq7BRZfD9rVhnX4TwJ94X9U8hI/Qwh65sahjWCOplhQwV0WozN8yKRxFPIl3q
XXIon5afsIzNJavrEn9zNIsQXTALPv9I4euS708DBAufODdg4i2NAvifsdjNzXiX
lBETa5mW8TgTcWjGgdp0/973FY6jMvVBpC+i+qyQH4YOkci0ymyeQR+vlYkc7mqz
0buZqWFlfXIrBIXLl915CGbL4a7Gllq4NriSmIvALFLbrqj1HjsS/LvYixhyx8Pg
6xwvRkZWEq4VGBhJ0tRLhFiTmAcRjRyV2Onz+d9hmhzVdYi0VIXC9UoJp1YPxFn5
Wgli9+jZS/zw1hzs2BdP2IX0MbASkOvph7F4sQGWOPUXptkdlvocle+J4602EMwu
PsPW7Cl/bOZasXfV7iUHyEaWd5fi5GDKPaNZLfhsJ+AQbFzOheAOTfNFPtTaTfN6
VBfDyoAXz8rTE1qYaVV51rlynBxiFYFBltOntVYUMWkIZbXoNuXl+4ovX4prLyz4
g2AP0zxtapDjHtNE2PwbZatCTyDbmkeFtRryK+pIy7oi5YViyTSD7XmQk0rfCYje
HFD/uZgtKDYKNyOxYqC9oLDYmiPqTkxeSDQJZvTR9k6hb88+yhx3tR+dA9A1bDiR
2hfr5coxjzpPOLdQgMXJHNE+VKdLVE9cG/Q2/mFLDTg3+IJPJLC5+g+4nav2EIso
Co7n70b4vcTOs3kmKXlNPdrOyBaW87afDKoV1JVNW2bTRKqn1NZxdgd7EX6Q+nvY
rn238rm6J+/HK9O1AVunhat1cUtj/pykqrdmpyRJPJadAOiAPGtnCchNhVPCKvxg
yRTgA8Km2XtqRU+1IqKrtflyuyZtpwJmiPPRzMZ3/I/rYYKkRQpSVPmC5JxEzYI5
HmtaHnNjNMDg9Nxn5arMRXdcwQhqShAbKnLs5uNOCAu3lf4wKoaqkmDCUJ9xnbYV
+DureRhe78xn5oU9ldWFfaaVmANcfyhPi5kOuvDkhU0WBEPw0Uq34nqWSyXb9vrS
arIUXMP3l4lEKNna/hCyGeblVEFRyGoJyRhYawRmX/crs7KpFHmSVYNz80VLV6uV
yIWsT/bVyeqNUTO+YEa9YG9PkZW80eDl/zGXC0vRN565gfN0O+3yjJYWfNyFdF3B
rux3cAhzdXMrVme+GPwImZWUS/H7bM+xuazFFpHZmG4Ls6pEFG/VzZEkGGH/lAh6
m66WowuZHuRpprj1xrvuukD1BSEyLt1TpQKGFCQgCL9hWbOIshacrL6DKFqOpwcZ
Uqm8QqBmazbOtqAPi8cHwnupWN2fa3XULtAFEJf7IsZ42ZPyIDApUm7nwQlw0uxv
AKSpSrncSK1opZILKbX4u7Ohldj7Fr8ygzxzenNgLFMXFHHuqhcEEVSf6IpqGE2c
ubvULnHfGKZ/Ri7a/JvwIw==
`protect END_PROTECTED
