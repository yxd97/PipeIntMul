`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGPL2F5u4VzBxGn1+usTDhKkAofEVrp5YDTDgO1+M9Ru/oHQCw3RcwsJZPWYB/9x
nHWvY13L2S+JhWtxEe3xYPnvQfPDoh1X+BO7rKzBomnW8gtKhVE7w25bCRf2uFlX
aJGBJsbThaqrhbmnjiAvzEBZ6Lj4JF0acEzBwGY+ZLVO8z11vbnenYwP9XE2bXYx
pwG2P62Z3Eh61BoK52mSasNLY0s5KdYQur/mOOgt3uVoWtMFkmftIWSes17PZvFh
UujVvHWP3wRWt2coRMiwjFC4dDoIR3V8gMUblYgIOjrR3gr/EbY2fGXLg7TqVxpW
CPCvT6yZTwMYAzyz3ddZudZCiZtYQkoQ0aVSH6lxx3fdTGBsWjCFYeZVzVhLziZE
FHIAX4hpdFlsHaH38S2eB3NfHXryDI1GShQurW47nys/KC/1WiWqVRmi3B8B392E
hKQqBDdc6wHfeyY15wdfkczymUZgIomEiFUqE/4Bb1hUBdm0Tr6Da9145h1/o2G9
615gEsKtxCIDSZnSUk+BRT57l2HmOOVdqFeP6lB3n11KHDTUepXM+n799Z8XU+Xo
`protect END_PROTECTED
