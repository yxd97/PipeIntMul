`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m4afYht5pHJVu3YrL7PALw1PyNmT79+KuebqT9EJ3CoK1/qHRzbGfedx6ESlg9I1
uV0HWDxJhCDpN34uC6s972/16ajMPIzzunAnllxRWx1FthE0kgto/sBqlzc3R7Mc
/cK+4y4WH0ny/2b3ZD3EtZZ+K/nk1RUzRb1cxHNeo2FIOAzdwWDEIpF7c3GxpP0E
tel6l1/lGgn7NkoEUx+j4p7o5rCGByebSQ9TU91Qr3DZpqFPc64GepS1KyjOW1sv
5rT5sZpD3/8l24dNfMuwDUfyJqw+UbupH4he+HhN7mP/AQ71jVbkzY6T8Rw4hcSo
uxfMTL55Vwfrf1dMSSE0BG/yZWKDu6wnl6n2t761VAvnrrzFd1RlzPQkmz+OuTgY
zNXKBTPSgFNQ+heMEzz/jcgiB3teFlE1AMb7aVI+wexTrCn2r9TTRcluYiK3U+/H
l+G4FA0qbHHTUhAXokO+qJJTu7FmvYUncCvE5FTD75OY2dd1WJJMX+VkwuPs/f00
4+SgsdI5f46QsWxyq4G/GYdTdJ7fZINT9I6hr6ydVvOhMV0JunUKPgVzM4O5Ou/X
q9qYpolB+JnJmwwasqy0RQ1kVQEwLnOPQhwkWpWTAo4I1ZGX0RvbqkWrGupzUwT5
sa+8/0E53qZ3xpqgmGFCAM5BfLjkHjtJzXUxNZkucODlvTUWfsgFV2et4QHJhpPG
rdlqEnmpi37MPRYTZW/ZrMmlWMjuLew8ALk8BnKsnPVeDbUyxQVp5udAQDN6B3EN
LPOuJjichnzahyFPKrkKonCncznNrMcHrvKWt25o+IRWJ4AN34bKa2OcJzEWMIQj
i+W51yu/PyGwvjMdPHe6yBbDv7lKVsZ3K+gRnjn3/yEEkGGvmYUI5S03a0WbJ6iN
4E+Sxep8hgYFZIPabic1r9iPxScJhKtAJSCvQJrPbQw933PXX0Q4/zwcMWrceXk1
7I47jDTDqbkNHpgj1/xANJBm6M/089U7OqT6uuXxLho1E9296A4PiKETAS/XH2lG
h4/92nA08ZbvxR/4IK9q9J2EhD59YFruh9UaGKcop/7fz0wxHwuI4Ectjp3uFCxa
`protect END_PROTECTED
