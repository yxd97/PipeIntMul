`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k6X7BSxzl6xnnPGA12QMv/h5z1kgbbZ6hLU1TapTgul1RH7CWobKHhZ+/Bf01mch
zQpxlV33tcEByV+MRxiNty+xEuVYwx6HDV+24J0Tfwlk2pMi3hoR0zkF6A45M4po
0/xGYXGkT5a0GYb4dACfN7otCC7YpuqClynbv/h6+BSasWI7OwYiJHZz2XI7pWdb
Vr8A4miwyLIq97pFNptN7Tn/yp28tH5sr0lNjnXnP+HC2hsGh7KeHhHixur+tu39
PlPH/WaQ0p01m8uDvReRlXMTpWA4E3BlDfwmUuUCY3o4MMolz1pRNOHfgDVDWvkX
0omdZjfTPsPs7lgw0SoLly9YkMVEheKzfMPTdy1AAL6fd2epybgYqE2lXZ06Hd8Z
CDWzQwN6qAPqsfw8zhmxh+3yGcByofxwuMWfma5sWY01u4/1mZhEW+dZERHcEtaI
AL5pi8o4hP70noG8etai+kqzlK6VJqI6RfEG6DANXdGE8rKmRhej2eDiw0teeoU2
5+G3XBZCfhSTs4jZUc4DlLKv/SbewChNhPyD1hLnm4Bvu7lq5u5ENXXS1gC5RwGe
48fy+XPV9q3CMVktcQiT6Iyy+7o/cUs+N698r+qrXLvUC1aLBhVlSwx//TR6g/EN
gjewEqq0enFwvCAai9jdBTUdeIJy9+JlYZjmP9zjFKvFOGDayiSX67Yxtg138gHZ
gfrW1KOkoE27QIvUOojfpaLUeuoZY8E8s2WBdZhzh8q5RP3citly+sm+boOdC8d3
qBCS2mY2VDz3gvmRVYk8ns1k6RflWOh7236r/lRum5ZVoA85wQw0yFH7HLoZEGGC
W+q6c+qed5Q2dzEAz/eUfA==
`protect END_PROTECTED
