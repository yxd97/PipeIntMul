`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QL2USFLmbN7rVWR5J5tEbUkD6cRdw48ppqIoANGleoAf2ud7wJWHRwV7AXm02pVW
/Kd7setRbbbTN6bU5Ul62roNv1qcdtRgRrvU3AeZ2a9PyBPLdDm2sotpTjXbtFpZ
2/UmUcR2s0o18fq0g66tteKBoG/Erf5thgtN7y7ZGMgXdDAIh9x6Fo9CQJtZpNuE
AE2F4y+R4DdGCpngDA4b5Wd98CVbJ0N+fBHXKXBFWZL8opMUMikJqmAXvPGkw6uC
1tqGBu7vTqQJy6xrQMLqgl214rtMNNS6RdBbl+R0vbPy66gtl5YPQGLkNuj7qnYT
zlZVXh+2TZY1HyXv+dcnEtDIdZDgr3ZJIv34AERGM6Ae9VecIWckQgPFXht0lfeH
UfgzFbY1WKUB1M1bwc/m5XWZgts+sghVLJw0dqMqmysvOrSHkAixyq6g5jKEZEz9
EpMbpcE30AzVRZshRXRLQ6GR/TRZms3Fmu7/95SdTsCvsCi3U05b2mtKaA8+LGMY
HI9fCT7ED8jGjd2mb90egtTxQBIug+VfxNQI0CA92qoddNji2ms5gow3Stpf3kNn
GlfIEYVSq/b2F/h+kIXa9F1sPVEdkkhUlSQd7EL1Uu+P1Eh+RAhEAIt69Hb12mRK
/z0wXr1x0HzatvplME3wjonJWEZYAq1AQVi8XNPV5qG3/Yno1NSDQAwk7ZeY3+DH
F24OLQ1D0BqT6IXGj6HWM+pWxF/u9KDtjyF6UBO/Dxz6o7GiUTwajRpSb5Fs/MdG
2V9u432ZPEVuQFf+lm+keHsJdURGo/y+W9TNBSwi0+lcYve+Y/SjLgSU//5LA0kM
SBoClEFTmKslEZA2o8tyUNoKfjMKWjVSwV5HW1/4dW9iQItMn4ChI3zVSaZ5CuaJ
`protect END_PROTECTED
