`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rp1aDRzKnx8r6OuXP2YtQG0vvpY756FZ8eZOo+l7Zpuq1VwXfp/XiLBMACxJrfjx
ACNmWXWZGhfEjdUB30YqfW56UOtL95DOYCvgyoBUaiLe5DP3Khh5kmWehUiSByQA
S0uh0MmymSBen2w9/P99DQuANQX+DmsUkt/SNAo1mxPp19KWjilbst3O2SEuC5PS
uj0yHlrkf52m0I/rjwoCH9tH8z6T0Ms0qsooYxKylBLpo+NChx67+DbFqsVHB+xG
DIqRrS79G/sjTLy0fOYMhCyBeSus5CPrVttDUZ2o3ekE4z+UH1ZWjPE6T+0HGyS3
S9qqcQHKS7oSJBvFq333bx+jSwaQ8t5hNJ6DqiDChYr53slKwjfBnG3n1mmOqOnx
esRqKNCKWe3zgbMqQyG23xpVOpGStr+XhzZUUhPOE1FdBq/hN5fTzIHTN5f0golH
3SPPvCFTBn9z0c3Wqmj+DKKVMP+q3RoikTVXwu89XaAUeVqk8wLLTRv9bolI5bp+
dBJs55nb/RjcpU3V/AtpPV6aHj5x2F2tRhg13jjKw+FCUEgo0bzerti9abWnpm9y
SGeMF2Ex6YiLx/syJdjZJT/wlOs10koxhi6EBWydrIHaq4RyaTwStzn1h4GUitcu
oFlXoZdCIWEdQQUy+KSkr2EI/glZcI5nzveI1yjigc5ou5OkNNTAPogszGsUH03X
Zd+aa6v1NveWUYESZ9iqnVdD8ltZFiCiIjBI6s1nkfxABpekLmhAYCTcO5DrRwO+
2P6Qt9owR31J7dNu608qIpM2gHX/+qjV3u3nitQ6d7FmncA+KGriHyRgWUFNH/oJ
urkCEacJ8wOVdAROMIT9DgQ5H9nuhQqC1Er+NMhmcQ11kG3jMjbRkFUVn5ptRiHq
L/J0FhNtz2mIxmZm6dGs8ZTeaHqt3kc52eAz2PScNFbKUDIqWUVBqJOu9qVGJA7k
nvcZORj+lkr1pD/G2aQ/OlIFb8erQiOVkEyPvPCW2JFq1fEunF47Z1BCCDya7noz
VUzHoewub2mvsdo/Juy+raJqNb3Kw1fBbyuHrOyPD9cBg0lyVkBNlgM2109qGqVe
A3NTgYbaBgMGUWJdkXjFFqbcsM2WfYNWi+5ik05an+8yQ3gUa6tLJy2kdK0n1xSL
vjDy6WULxya7xakH+T0sZyGsKTYGIkG2m4dXidS/DdHdPFtx5ZSZ6cPwQLKJAfL6
rc7LOPK+wzON3Mdr5/ZAyyBWeNtnMpQQlIySSKN2bT36Jz5NGNMvi8sGdEyEfxPq
hjrlX1ZBw69bVvcfSl1NDvtbcJbTVnhsJMx8zB59/8qy+XRUxaLC6AHyHjwtAYnM
woz6P3dAGTqr014ALGCdhdON/w8kMTHV68OO95Y1+xav4/dkhKvyzmjMoJlecIes
aB6GBObHchB9NNSqg51LtTAJvPFDm60NMvoW2wQ5y2QoRhMKsCnpjy2+WpceRft/
AwnsFNjb7MWmpRWWbi2gHx5LI3JrurR0LKOJ7BM7822kLAtNxFCRwg/7BipsKCYk
OVej55l6Kzs7GmI0yN2HeWzhBhEVMMF0iUxWJBQLGMaQunwQXiydw5TtE6RA4J8M
/KfnF7LUJOzzY1dvSA/WI0Z5tktcJXPSn1DvEhDXwouySr4A0BEOVxP59DlScKF2
BX0l/ZlzbDszlwE7SU/FL0foc7VMimC2QZGs1WTu3AK+xb9bwoZmV/NaZJ5Uh7KD
WOd7CqA/o1oICtUR/1HBBhUR9SyKs1Sr1inxW2DRTfzoVHQPdy07iV8BpIs4QFj5
S9socuAxy8W91noyLPlejvOJyHLm+CIi3B0UrhLmQHmC9dTjir8Ay47guFIP0+RO
PgDq7tmhZRVZTnAdiV9itWIkrciopTe1hmakfbIgzgHdpffLRfajH5/3cI+1lpOy
IORPpU1FyquQHjg2VjY8rdb6/DwBKB/QGN/QN2io3+h+x3apiRWCrlAKxFtQZgQh
DQU9O86ZHmNE3vAGz8TziOFdZ/7+Cu6+nkSP/0CuBcBXP6+0gy9TJRcqju5XPc6H
9VDGSoMFpv01zIrudtFA+Gdu9t1DhdaYt6Wz7U1eDEl/1TLcP9RVOkPtC6NJ9HXT
g2z1ioyfMjJy7way2UQ13rQlk9yup0nYjVpZXbMID6EqDTM7/sseDP3EZSpryz9l
LkOZPAASquzxqh1BUj0nh5hvc4JQQI4Cccdnk2qawf+ii5NMNLT18MLJLN1uUQbw
FXmx5Z26GHndNRHSyUg8x9rmCeVEucbmkYgwOpkSS405b0FDu3GBlyMXo7U4OQk2
d04meTvBm768+ZoR7wLN59MR3DOxsGacLsAsxSvgfOV0n8B/wxLRf/0m+92CE9Q4
kbLcxcpOwpqvnfHt9wm3Eqj+M2w8Wu2XEyyqLqML7yGrBUrEkVa9NmW32ligTKe7
jf4rP0PbTUo5fPBT5eFFzNTwZJXUWmUZeW4WJInTCBTtSPsdWIVvU0jjKq0JAR3t
Oz3n0yZBSeSckM+/pRpp+BW2p4dNBfaovPWtGGvjPeUzGZMsS7G1eOAC28QFGLWd
hfblXExGVhVFp0gJpz+lLDU5mGeV1MUKC886az1l35Ad4zKlfqYitcFybtjhon0d
NcrmgU6PFgASXviLHNa4pHiUsk37KaiCg/8YfwdPHh4TwhEXodW0t4hzRah3B7PQ
kYjWNjZ20hvpANU4HBWUOHgAddp1NGTc9BcxCl2y7It8hznbOyOMLh6rdqOPGMlB
lK8dCUnx5oQWe1vugYyY9yUxxJGHV977gLhg4Kkeo+Q2pYywu7lWxaqa3YweCQL/
5OTGHhPMFgyzXF9NLUv4U7m7DijT+VcsPm5UbgkJ4rYMfA557S0qbd5JftqEphCC
y0PnmrmvOhTLMdQNDvZzhLmcehHyhWXRTj5FzB1xPLoHzJGxEXZ5VMN6OOKzbXev
ohJJpzvmL1/0peCxlxMvHkXPNDfrZdK9rEFOL33+JsoyhWbk/nI/9nweT7qTZ6aZ
5tVqUy8lz5zGInm+ExZ6QJcJv9KnDHaItZnfZdWKqZeKPL/fbdA7jb2AmdFU7nWy
MGQgejtG6plwqmmP6rRXK9ALwkMokHAn2fCwIkBBT//duo5dzOFjNUI6kbmuETRP
hNjFJVWQT3axmTdyBNx3oY/KWOR0W+wU0lCFgMRnj1sJttXi4qpRw5+VdRibdegv
CWb7SQu3KJrgvBnXqAg+QmL/IWmhZI9VzfyCDNBbQwgYdX4+WT9kS3PMc7kZLyoo
a6Lw/7+H7Ap4QR6hTcuiCdsohoa24R/a4BxN+jyn9Q5C9YrLdVg95Qr7ySl1lWNV
xD7IBCLU3lkN4jcSFoRjbRg1UQMNCL8CnMp7ycTL6COe7PuHTCY2iqsMmQ3CxEFP
xtCFcVU16M6p4jMpjorilg9XaGccWGGCmhHJQV3sbolYnZv4B5qX9H7J4R9m6hMA
QtBLUDXdSRv2/XHsSjoFzEcMnCSxJez5RZELf/Q309fCeqgv72ecaNHvWZfD83iM
uV57+xl2RVBzVPV/k3mOC4iB15lRDxSIdHTLPd/h6XfpLtwP37RwWeRbAmMKp4K9
f7x9FFBRsfEEwlVNawYS55HPOcgT/LL7rFjRacFMWbxTDQ8syAWajU1Fco6Dvj/n
eeTbG8tS6Ej9aoyxV72QkhOJFSibWsHVHfykWktuTFSiw93dKZ4cQLcngh0LqDqV
lE3YbFtLSRWJ6fowl5jt9ggyg97IyRyZSOkbkMxKokiybAIRIemeBPRaP+Ah+gFM
v8vLCGQwZUl2N7JZF+EA1FqPq9RJRQCHG4hkHfggCnQOCtM+SEwpUvdyisJHlF7z
FA1mBGXqR0OaNExj2SZIs7fz4aUFvhm9ho+qIHw7DqRV2daaVLr0L7iCtnj3A4sh
zaE9ZdpvexDNBCYr5bDnMcmld4LtoHqChpWc1SLSyYN3egmvqakIs7L629XHF0N9
4mc01l6AYxNvbxMTUA4W5uovzpfBNEnwgw2WeOLL04BaLfdp8slTbKRzkx+QOxMp
WMUQU0gi5XSWvED/504AAOPhPSZr7ECXgjX/w0oCMGCtkzRlHoz3611nZwRPmS8h
wfYl0nZVLh6w1AlXDwHOcYp9yTiLvLVVLlE07ETmUZm3s2wfL+GUzrAELLqQueKz
C2K8iw+YhZDxp8j9Im8ju2Gn4EQWwskfM78Kc/HRFwGRqEzMr/0rgyPhmuO4nKm9
KzUckt/vRRtTc+znIbJ6qGx/z32GNMHthWI8ncGjwCpn2k26KcsG5pdnXJ6/ATwu
4oPY7nnHwvvtD5aBDThtSjFmHChy7xZxTpxIohbxiq8ghCek2NFCQvdFT2MRvqbz
YDSBlKUWfi1hXLLhAqHqfhtgTQtBscHypW+EllM6OEIPZ7akMkE6+HVutCYoq3aq
8HnH31fpb9KQPt/Ly7HAW1DWC3AbA6UksZK9jJ/oXub17Ac2qO7/f7UqakWVQARf
LbvzokbpM/QcDepT45gzYpyCHbH+VRkjAZX+CUvRTA3t1QbiBCaF4EQ7v5KcDBAq
BnZJ7uWWlPqlFpBVRBHMNSMgHXHDhvZ9JNBCj1i0QsuARpwBvlBszgYLDHVntTy3
kRaJHlAiZvxqgANev0/cpSpBNW5nrK2VfdbFM5GNHGjcMa1taqtitMk5IukSan3o
7ub0WbPJHmEZPcWBwIBkLviN8dPD5lSxBMh9CUeOxLdvrl3cq78cjNNhTWNvvBcf
oBSS/tEZpXaLF0sEd0/nk55FuGmnz+KxRQTEyWqWQfHX/Irjuzrd/Php3X40pluR
3cBqzjwJGpPGfwGmpmsEWajjNVOlqqX19xiR3hImG9OTDkSzunqCh8AXUy6fLTNk
FfAKJT9v8/zlhu8EFPuuB4gVcGzgzaiOYZ2ItDmxGV2cOJEOVo5lg4ID74Q3fK7Q
bgJj8A7uQYrKADGD1FlMeKr69ykcyZJa/F5OIvgQOCW/BSykXjcsExVVhrqmWsq9
m9xbOtE6rM05be4RMLVl37oHwSGc07+gDaUQu3p0Ts9Rxpb8lssTSGwU5I08EEW5
ePj+e1vEC7sYw0aOAi0kDSLG0jM5HfFEIJN7YnZWnERr1MX3HaTK5A1pz3rx4ZeI
ydSGiCinNjnIeTC/ccVnl0hG9/YGakMsNqAnqv719aSYMB7dEgMaxuxRoAoqMjHS
hXIHE3zybmsUzSbo0jzeS/Tr9rnIzfJDDlIf05jI545BoJrTQJzhEqmSwoay5sWA
QOn2nfb6njQ0qLX8HOBFAxH1Ycz8eRHzDVit8ojZDnv9pzxA2gAidtBi7M1ki3o5
zNhCxVmRrfCvIQfmovqAn3IN7V2I7+Yi481ctXBulMrYwnjOSHQLMbwzBJb3knBd
y1iasNI3/3DaMgQ1Jp5sJRUIrQDDl7/Rdkhi6/vf04i8YBX6QTecLVHSv7UPsbRZ
FWRy5U6cZuvYD9ylFyfvVpeLleqKE9+buPn/dZMTaR534Db8A0dGxQzjyrQD3b4w
IGVSU2DkFlaPAtEOdKXSQsLxkjvx4mrlA7MAGhDU4MVRJylAxzh1Ijizk0lksqvQ
wTdiJERjVef/OshvSZJFvKdzClKIWk1yAfceVYwio1WvKkMFoNdVRoJy6lyMKfnR
MLRm/+u73pjYF3eWEm1v8h81V9L6pOnqK8ljQ3f0i1zdM58utxPjCjrlJOh0GGuN
zVm+WtsowawrsnpgCEY8X1NbdFnTpELTfDIiOcsDoX/SlAZcqqJMxAoFFNMiO0QM
CD8jsQ3w8KAbiBlhAIyWS/nEfCZT9EzvXZQJiGEWJXBBFVBR5uwegvvb6Emo1of1
4PMv9nTsxYlBppCrsqfl7yKvSui1ASmu2tUO5eF0BwBpZ+WQxTIZhhbaUZTInDjo
maDpBkiF4mssho56HGeFdf5fpEC4AByKVqqZeQvWYfGYHjLPUxSK0ztoxmoqxAKI
z3HAMzhbGkPYmUtqtJuRhq3/Ksmx/kv7K+DxUuYHvnJ7FMVBwLEJd+480x7BvY/+
c8jBkniYUjofKOZakuTRsfZxjsP6dc4pXY9/PUjHNBvrDVJQaMdx0tNeE6cirjGT
azbrQZ5Zju0aYT8cni3m6Kn+8xqJFcz6JzFq6JWI/zYEdDwVwx5ZzbU09bt8jY+e
GWTMRmnK2Bu5CIs9Uhv7orrUcOHC39Eebmer80Qhd9IDGY27foQHaxScBuny+h2u
lRYpAyPRS+rYf+paM1QKoAiiH2Enldl/hDzsRQlpfIdaiEl2ZLxX8clDY4vCCwp+
tuNFPSgB2OiPrQ+qNoytUITyCY+uZPvsmgRK68Vhnh3Tj0J6GLm5wTvGrekVsxNz
A/JPPDb6HdybLCOJwTof/Wl2wRJ09bdvMGuStsSmLijQv/XS++AmPmt6ndp7VLLm
n14WH8c1fS9wn6d3TxM8q4xkQQKCvQN22W/NcWKzTVg776xRcgLOEFulOsw7eEUx
12H7edGsW43ORYBRa5JKRsk4XUUwTuv1CB7rq1a9Jj72+jvY98n+uOdKNYzVqKU6
HPxx6Ysj7HTBIwk63gFkfSDT/nWBXdq2XqNvc0CejKCdqAGjv2jbe+SFzR5ZSa87
An/8eUsFR6da6i56CUJ3So6wltuepvQqt7OeDKgLEbePyj+91ideLDvVOTU32pBo
KBFM+ntzVyVXAI8mIUxtN2o9VFN68ulsfzd4EplKprAmEJeO6r181fNPgS9JS4fQ
fltK3Mf1g2+V0zTFV1WHs/Hy93pz+SbXLZSKsl1Ov+YrtjOH7DfyFGRA0edn7HwN
pueppIi8JYipDSamQFJy0wBI6FN25ltruzwYNPfTBaW6407Qu0k5XZS3/0HsQMJ7
h+RgGUdnsKqhfeAaKADBQP+gR8B6+Ac4NEdFUzbI/FNag+rM+CssNSFlHaOmIALe
bR1TZzdoIqCUS1SDKTwYAPzJ3gTBgGkEqUVfZQILIUAh3NE+hdDom5i1CUEQmBAD
jy+Sz290vtap7W6LBZS5jHLTGehEmRwQBHIy/us7HLVF3WjlNH9bNEcerdYXvL9Q
Cc6Ftu8yI/p6tjpRCMzztWPWlNDW39y3lXiMnF3goRT2Sg6g1M2VboRbO8i+5Dkn
PClASyPbppnx2r/f/AWmknja8dUsO8E2FNubafMDbPY5zmQ4IWwQUW6haunwPAr4
CuUbDql5emgXcyZ9qczgampklXngnkHNeiFTxAwq6ZgXBZUvuFh+5q0BiqFEUdnd
siIOtBRJTRR4XbXkAdynhbTbJJFRcJmtgDg3Upjkg5MkUyAD8tCZkAavemz1WH3F
l7meSjxtYd0wmfBGC7UVR1PjxfJlRwwFh2IDUylgOy5StRuWLhgCWNgHyHePUJDQ
SZKC4Gq5zC9nzeD+8m3DyE8M1POR6mFu1SyvZjL5PUDbXdPtFQZtpKh627pXE0Km
wuQqzx3Y+73vbWZ0bTdoEOtOdLG7q4nh0rxy0AomE4VjFFCpx0Knj6oiTh6BLC3R
1vG0J5buMt8VSleY7rTZf6QzPHQQ84AP0x8dOcaQZPvqzNtScwZ78E721vUOaH6a
T/gd9mYJnO4QN8UDDPdgC8dyj1tBpxrDqk3iasBfJyjRwBDezTKYBG6lKguPX1/v
hs7UFbq4fmDEtqJaLSC9iMxkNyokHQQWOPktm5ZEb6X+t6P3ckwC2nd9wO/eLHGQ
1WqmPj8ygImYP0v76luHDOUFkj7+zvqXdI+9JqMbtAM1u49xtNUNMvpN4gHQuVb2
CmW7RANMSL3NWRY+5zJ2q3ExkP8AzzS4SAaVpfNGWGb0fpFjh6MVFZZV3uV7u3rn
u6C87OH2BYME+VW2/AQbjtS43QFoE8Q8rUIkfqIFxa1wfhVuK3UopGDAPWWqaWLz
hlIs1N4FG7ucxm1YH62pMvUA3ut5hpxqWen0BH12uiV3U6RGVV+GGzVi0/dWt0Rq
mXJExynFZ0FqmNANznzB30w8XghUK8muyUn0lnH/PU8678G5UIu6VeOBM+ihKV+c
df9MJ/4BcttgtOPh0Uct9AePtBaAP0GILSvkPhIKNWjrMngI6Oo3vUZhffUUpYqQ
99L5RRpule+Qyrllq9r1AQm0R9hCTPnj/nHpf3OibudPxUc3zhOqbL7JhBakiPDF
vEY0RNF5epB0MqjWZU01n2IwWSSJSDrvF4wOC7mcrhD4h/uxQmP+jfx6Xk2UAndA
fQB9P2GXQHZnH0z1a5OrsvmDbGL6/ceL1uJxPQs+iaiigCh6EFmOEwGxKuQ8++i9
AM46OJfImLRyW/vF3F3KFwgsxe2KalaREAZdpQGPUx+tglUfTnXNX+6Yw2uEoqyM
iQccmmxXSaQEeQHPRs5dTAf8aEt7qKanVTcwWnk9ec6Y6+FTDU1o8BBVVGkHPUnV
01ZXdVVwkRoqwUXAmqHKpyPVBrHTa/AmqwzAvWZK0U6rWqo/eh8L7Vvl3gQTd1Gn
RfHnhHb6RFkId1tehimwKUNwdg9ehyizRxtaa8x6wt/omm3ENtXKiawUx5gv7SPT
U0THKvS2kH6i+KvOwwtb2pkl3AheUeQR8jbiYr1HWJZaDpAaZzS299bgmuu/WKeJ
lFwxUknwAlk5tlKWi7+wFxMYv6iVjJUX1jbYHQWKwBX2vownhmPjT0def8sp6+cQ
WYJ4t9ZTTmJUC/fHVKZsupcvGxcEcq4b0ctfq0gFRCSiHKZpNMvSJAHQwNvrPLuf
K0RJ/QaNqkdeL/dLEam2GjwQ0Nq5ybI3nErm903ot0CSV6y2JrH6w6AKFA6oxJzf
+zA84xbpDrAnlf5sGfKtsGF/tQRqG2MS48jOBADbvdlQETecOhgT/UA2sj7teJ0/
hYKmVNz6X/wJrQRgllit9m/00m3/qxmyytJ9Udrp5vwW8KRxSlbT3j5q3qLHNZkH
8w9VRgb0spByXxQfVXb9aECM7KzYgSISq9gDeBoc6+ABV1+A2M6zesCmae0yBiN/
KgBDiJgq0S9wcpkfSARBnWSzQlLAw3990nfn8q2RrrS3spn55LwtF9cxTe6rDhXR
s0U6QzC6V9abn/9BAwz5jNHjbqiEpELFnQZAFFi/vAYy1BmdllDuGBs+85kPFiQO
uCZAuXPalbn9dmt7FO9v8wp0WVhH46OZcRiKFwU57LGFjFxTPEugc5QH6QmZV4t7
KjCf4j52BL8nY8CYqWLLL21Pv6hTyQWKaQV4jiQFSUZHlHPJ6HT1V5pYFvj1XKjw
OpnaOFhMEV9vevYedZZvEGxi+Cgm+RNTDCGbhGjXCIkydhvHj4UxNXg3K2yZ2m1N
ECrfcdsGZl0Kwb+QGTCyQrUQRv7lgprT6k2ngsGO2VxS213ODqjc+JOh7MtvMu5w
iK7EejqdplFwQKjWJSpKe+lskPBhKqqRBifmGtyCIGdOJIWRxse3j2R/v0AzW78W
gGu0XlDh24kJmpCYEsdz/kJVcGe0Z6Kh8hitElBN3YSg15eDJQtCdz8Cy3UByKbN
6gXe0gAdQMFa0Hd4Tdd+EDuw0+aswej0vChNO3WL/+auaOmvJGV7bWTLPzEjLwsQ
0TOTppXQ3xmOoaH+HuKcl5YW38/bZgTVqpvG2etL2kC5ak3eBkjwIk/9Ep2JyBhj
NnSHS5UAsAkIJMR91NdT6D5MJZCedfXgkUX16XEHMSB3/h+ueeHyFLpilryd1I/z
oSvmDwVNG93LnMqD/jGgfLoO1aFlB/tpYN174M+6fsX3qE95cpWqyb/i3ZebLuwn
tbFTFsoMCqnPp/o3+8qmsYCFvHllrU+68un3EHx0asygMWbA9PRpirR+X9JUUbsi
7KFZ+yezBef6P4CtpkNCc5f1Gyoa9PkUmRI8s4DpNWqiw8R+YBSTqx3+8I60fJRh
7xmp6GdZNeSz/qyYhaBQFHMNGqB90mhvgrguKex/AbRYEa5dul3T34kdcQU9X/Jl
xw60ROSy0tdwupNDktlYyTW6PM0OupP66tJJQui3pSl0UE2tH2WLI/0QnmZgrzAM
qUWly/7Znj9UpQLC227cfvMlLyeRJ8IOeAfEQ83GJL2Vp1bRjZJJnWi/Z2nmK3ox
RY0ZoRZakkXQWI5U/eUdQrDUIDon3ifztNWy6PYchUIwOf539GI+yCZBO+vnzHbm
yvy19K3CNS+kCDZL2RieTL+sGTjmP5aRT4olg78jCpVNwS6pfogw8QzHA8b7VOZA
LAI7UL3hIUPl68UgIr9dvyT4h2AZJZHRkRxWts0cJ3F3Ql0syZ4AVksaU731rPFc
lgxk1gQaZd0WIi05fdLQxPwCw98FC21wvARtsLWU1clp7S4UZr1iJ1ny2AQdQ4Ni
ddfME3at7sLHhpCfKaZxjMcUILxgMW8TAE97RzcZIgSpBZsT8dgDbU/ugriuvhKZ
be3E6fHsQd70sVKcWEtrdTdxMnMT+2bzIvlltjkB0fE5Iy5tHug4xO02dqfKGdjl
K0I8iEq+DUIWlWBAZ5Tcvzzrg1tiqqYzPf1Y2eZeP3S9OLmUo5R4F19stAAo53NM
rT/W0gH2zzSxC74jnnVs1hfnIQ1wWu0U9KMcLsI3JjXmxMdIRCxCBfBW3ehrjyNs
3tXMHfE5xVyIG8r6ZFmnuUF8GrD+RSMxEkdioA55wpfVHHCVGmkl0FZaD33Z0L/L
6f+xhgYsJRN3+HJua+SWlAru0A5qOKviXzkoslrem1QpJgQ0w/MlG1sTKjzdBlBB
wA+1mtxe3O3/LdfDqfOBG0qcHV/mpC24NxU5s94o0qPD2VKf0pyKAx+bJYJ2fV9m
9mGyUgayIU7P45HCWS/qtg0DxOJOMRcgcb/SRl12/GuRQnx+HO9xBz/ltlBwmJ9q
vrxGBnOoOvjNrvbDTerhMmDVEMFJ5FUfL70eeOPGJMagLZwF/bmZ9SaLPFtREqfP
p/LrlV94aKN6UKan1tfo9oRoP5XwJmMBMA+zH2FhPaM2msIQaSxpfetonRIZSMqx
lPc5w7XBUi2dZKWI0evYxFF34f6tutDjJyThe6VV3l9TeJkwf9y9lGMKDneWEbKP
UO/yUsrOVEmoh8Gfcb0bsSECxw2DEHUek8KFV/21VjC0LkRpY2JCkCX291GFWKPG
QwOWydnB7XHnfk9f+TsHA3K2cjKq/xK6XOTcvAAuKwRsNuynBdRKiSBRVbPxjnMI
WehCAMbGTyIdOoY6wCH50pdvWHROZsKN9D+8njFMzx3fmRS5mRs8bpAuttMXwDhf
mJJ+UoAsD596YC6wqpPIkWA+/9BrU+oMCxAhhbbFqDQL74H/aemVJIsC/khdScGx
UHjGJqUugSJixSf1sxZqq6jeQRu9lVF0nS9xZzfzGFn7LYADOip5GdCr3MEuiRTK
Ln7zIhOi2KXsGAkL0MNfiN799hZwwFvsTjdTLXolZVFgWTmH87hizArK5QfJ4/Yx
OAY01PADh0P7dZGjic4KaA7yRanHbktWcaSDrESpTz9iKnzEu3hPXtoYK8tH4qtT
5Bv7jouaJye7tYgiQ8Huwci3SIMDCkvcMlPRNbofOyfEaNjB5dXUCGJBGHomHKGr
6TQvMcP7bD2k44nxY0nDR6LCU1sAGYMCVIxK+ADK+JE+EPbCCq/SXsE37hzH4ZVH
0oC4Jrz+5ZQQC2kue5N1/UfrT7srkdFdKULXLaUkNwHxFFlODeh6EN3xzqOmhba7
mn16Z6AmTUg23iIibb/Iynv7ij+BrsvmfLp54nU9KICL/4291NzpmPBU4QD6qSE1
7cj9gN8Po9IuhhuRrcKv/6osMkKXKqworEJq0wjbXEvDE5MF9G0FSt8OZ/lIrfmK
BSPuWUCFLlD6SotATflIxzy05OpLrLnQzwzHxFEe+qVbQfhVi5+kxoBaplypIi+f
goLDibqJj8O/wXZrFJHKrmEKiPdqXC406fcHHEiVXiVw7A6bChgwtRYdzxmqu/Wv
ZBiKI3xdQu6l9SleGDg/kE8YUBrdO4iXbaV5IlRE6PuMo438Yh1ek1PXGSqScsmJ
udkhyVmILuSOYyg6Dgq+z0a7FKtapqoFb5jvAUuzAXIOUHUkcAclei3fpJ82Biie
XhxYHk/KqyNDgpO8STDzoRkkXnHipwSDgK3CvDS9F4L1JR/mWPllBbQcbc1RuutB
NHt6nlw480T+rys8ulG8tscXSAR4LRy1ZO25Kru2xTwyHm8LeAUvAyT4wSouGRjN
e+7AIShEbGQyw2bLvx0Wjh472Hhi+BkxKPvcH0Gtd56SMTftlBkvs/K3xQ7IzPOo
NwQ5Y4tYMEnkt3YJPR5UBBTFMCvPoHzcmG13yWUaOJpCB5GbCNMZFsxy12256hXx
bkzIvQqQGH7KfnWVX1N7zpJH1DW94l2fpnPfHnLOVWzO5FtRha93CvgdsHa49lYt
UaiYVNCY8cQIrCV5mcEZuDrkcTeEfTGaO9JDmi6PF41RH2feQiNH3pMT8NJwQjEr
kqaJxt2REZoSxx/NN+/gR9ugvAyBNxj7e03Fjia5U2OQuU7JzgOGFBaiZyCXbDmf
5GSNC8AlzldH12p2bhmCsHZZKOYfCvIg3fRo4gv/7i1mQeQAURMWWGJLLeTrVcbb
MINk9wNmS6uJFrNHk8UPSVdDtAJf5AkDQu3Lie2Wub5pNX7ioA/ZG7Y08w46r1gY
sYDQ8OpJIEROXanPiuXLf2GzUhJvCRWNzCQS08H8qUt4XVWNaK0+LKCT8GePOg0P
he3jJF7eWbo8m8vS1ol1n49cBC4XYGBQvMZXQE/6zhq71QGfPr8GQMYyyrQ9fJkB
S90jAcFsoITQCKpxh5tckOA8ho6p5Slt3q8SYvsUKdyzkVDY2/7br7RGRUl76ctI
DpPT3znu6dXE6GPoChwUESQR7NOYSxQv8I7QL96eXIWMj29UBbGejmsYBuNiYc2M
ROiPEben85mUUIPzn4LwNNooAgPso3nFHKG0m8UqEn3X3ys/5NuMCdiLcyw1Pg1o
5CFmiAMgkAPtwCYL+oyEEDPQVkcqLWczBX9lxtg7aLkozIfuP/Hy67UvyiU/cyKf
BiuY/VDEVyJSgaVAtJltmp3NrHn4ABtPT7KMRw7UnTIB880EC6c7j6ethFjVVkS9
k5Pfp19WRoee0Qb2kNDxgH21wFHas358nDioAWRPk9jCvzEjKaDaKhnlraqXQBEJ
levawrf7YtQAjFhgozmJAshUZC9fRIa2KaX32+sSlQ4nbfurJZP+tnJgYhF135tP
W5g/jE0Oo2Ga9VUoQlDEmz59jDmIFDCZAau49/rbP/qrmmdoWjxiW/kbimXo+URd
SnKrWunmW+OsVUZWibHTxUeWqNow4KLnz1Ot08sOvSq54X/CUT1+jgMpVVIr90q5
gARCAsj5vll49bk+h+FGzrxCqqTTRkt++kBJ4k5PFaHO55dePVfm6u3JkMjXlMIw
kqkfmJgnzAhJHqIMXaeHGsbz+dHPO9s3128Tk3FcRLayO6tmo1HMZXXxvzZY423s
oTEg46N2TtzAMABv9MRwyJqztuOMsDe2dI/5ZAucRi+wSA3aXhrXCPkVPM5IgiL8
u8TrmL1ROOcLjoOlox9sb16edrmX8CtSp0CbQmWa4pBqLvl/MfI1VlMGzPfee42w
eTUEqkih6gwHoRCaUK1Im0nPGz/mkDqL7TgeMrn5lb0dRHYEn88oBNij+ETT9DuO
NQ66fNAPm6amjjuzK8LnDI0I592TYdxWWt5NbNZdY/Ndw/1B4JWttG19RuP9trwD
CbjAJ3z7vTpVo8i4Bq5+o9HGmrAzDL4uwRw6KZ0yuD1rs+Ldf9jhH4G1+hCGI7w5
RrDcY0BHfoYyre5Qie/Do1Pjf1B3O/1t1d0auQwgVQtAOUXLGFGa1Iv46hW3/6sV
0Nl/05k4ts63IPqyQXCflcgKCM+A+JR0T9jwJfbsOE0=
`protect END_PROTECTED
