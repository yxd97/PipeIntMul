`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Q46JDm2fsDkfnQheO1IaCQg4N85U4jfLB4FmrogAZHwciK9zScW2K4IXVqPhcWh
ejItlY/qcPKhUS1bwaRsjx9F0JpzjNJyVXZgSzlW6DHjve9f4dSuHCldVMfnlkVp
bdL4EB+ouLR4F0DLubiVibLISBCoNAup4XxPOkY/fwRbgvphN62x2Z/PkKfAqmTo
bMLRDLfzr1bNh2ClwlRW02IVIcEmLChLO6Ah7mpO9DXUg3H3RFnSYqiLJIvjNzPs
8/vzfNHW/Qn7aL0/UnuB4sMz9V+hnFAxSj0JgFvk25nRoA/L+wXOeo6xOT0b3u5F
E3DIA07cn+F+GJHQbORWmJsBsUYu7mBWOnB2co03YHG5vTVJx5sF8MWMGheToe2s
pSO4jC0g3tMwz8RkfyXeb17M4WZia/EWj5RNwXdMEJK0R/WhBt/A95aUPGmzL5oZ
C8RidUhiKZ7jYNIvYNdH7xlxhBUiuFtdew07SZCCdf3TNsQFJfKP/U8q2M38vhbY
X7F/mZLaC5GG7nRtsd2ZRIajJr5wwLGJwK0kvt827Si9Q77fP5iR+mukPRQXU2W2
Wq2iCpGYoW6Gq8vA0TkK9SfAqejASuI/8mmhFwU7S/PzXp2lbAYBAQDYq+1Wltfq
jd/cgkW6OifncbxNDmtqT/y5w77C2uEKaaB4eNU/VyC3FXdWAlOvpWLYl3sw1Szq
7zm6uG1Ner7fCX/L+2TDoyanN4UmMwbopnK4mtww2YPUnQ3K0mKjFBnwQvTi46ac
eMtgOOk8+C6WOY8MhZ0FLEbp3SBlNwGWovve+w9SoiZFYgDfWPIUAzc2tlgh447c
E62dF9Hyij+QW7/zUn8IT6ogXWGrXPZ6W96mqka7L2ou3qZ9Pz18q2JAIkRLIEte
p+S8RRpS9sg8I/eFtRjbbe3NROZrR028D/GuVyTnwBy4pzdCw0DqOnh+A07+pYtH
iJv0X2cH6X9+1M1v/wP4fyTwyRR+qenGAFAqyYy4+R+A7FP0X7uXPW5fM6xn2D3I
328iINsKS2OsjAIhO62wNVpdpw7sb/AGYQtOXZfP/MjKxk22/VmRLefKvO+ZUn/F
RBjBopvUhFzbuf3zxBRoZj3O5E1My1iXUIOIUYh5OU5x2tufNz0it8iLDjIoTAfp
RxMc7uDUWKk0eEy/mf2ZM0l6EmPwr8uSJcjCAPtce8gnA73sPIGsPTtl/u/K9bK9
630dNyskBL30GO5lPm3zcOcTIuNv9xnSBVmqByAuVNwTDbiXq/JUIogqO4vutpjA
0aPlDtJHe+RkJDBsDXj0t2l6p9oGER3Aruo1TcZAnoi0L8Ceu/OlVLuJeJw30h7s
jgqoCsXwWmmtPcWJsWmrODLDuWIDcjjFMaVx66RaVFaCgw5/wf2mpEJzynIvo+Wp
eWRI0rEOjODJ0Kb/brfX/LbOAh15focfmweYzj4zjhgC5FBIwwgnG76SsaKKV31y
n0sKP8lAVhqRbU1FWQY4/6k/k1x8oWCJ9OZal9DqRQzVrnvil4QWWQmr2GsQUz+c
UwEt/nrnMOH+LB0RrzVXuVqXhMjQ8xIEtlgnYGopPzTGC6pjBC4l5qsKYTLPnGNa
dzvBt8Lb1G355YK3Ufo9cEukg9HuL6S9q1EvZfZl07CamoTqDlCFppwDhcjx+Z+4
XZ8JPdBU+j/yXhUFyvJme3KPI20b9f3h66GVwPCwKfyeMEovyepogQIe9Lr4LyH/
T1YIu7HWzxTdkNfqESjPlo6rdrXOaB7Q6auNyhe+7YJArN+Z4rXy5rkG3GhiYt8H
Hju3RxmnWeRVtPZaW/ClCTL5wxL/8Ru/51MH8z+W7tWuBmqzVHAa8RKdWGKEB2pw
J66U3YsqTNxohj8On6j6BCe4AKXCO2IAtmQlAFS5T5hTyovbZteyYuDjRQ2iHgsk
r9/7klUMXJM6/qZbEp+O79Fm/CY5NQ7XrqJJ8P1AaxVerV3lqGF2DGw/UC6P1r82
k9a/Z2d7UnXU1+MIb92/o46advzClYCK3bwWcKXnchEJHBH6jSJH5gkrHAPJFCW2
yDrDSNmmjx66jqf+ZLozCdY5Wlqe/npIZwSxWKSkyW79WPG0K3BJcTaCStWoOXPG
as9RpfK6tYTZhM9bZSN2oC+IiqgYgB+PQWRDaoCwTR1kiG68QBrx8Fsl2UAVouyK
xpOIlcK4HqtQrT4zTHxy37yMtEmzvphE3y7Ae5jbPN3UMVH7d+RK6iykUa1izyDc
R6QrUShc7MQtN1b8XPnU5U8AQrw85MNxEA6LrGQwmkA5iGE6W9SbyECcae1ufqWX
+RMQmoNB4dx+dFXA5n64zSVhsMApPatlYf8vzjcm6Ce9wJMoBMLyH41Ha53ShcOD
93xbiR59DdzWln0aXybZVr1BnTWwD1zfREDFQHAtW8AO2oaNo0RHftLicegOrMpn
YwxBmPowEBrTGN0+PPucvhG5gaRbZu5bKWoc1USTCQ8gerA3d0U5gW0GQhz+Si69
eKu6MhQDtsxzNzAKpbSi2UTUe8DVyU1uVNSzOXPMYDloZwCL8YtskR/uJ+h3ppkZ
eGh0sR4jVLcT8BWqA3AyJZxqXEjZuNu4D93E3XgWkO7E7yxhC4muXzAMKRnLrjmg
+dZhCWOlJmAvVaWRFGO6/6B1ZE0DdyEWZ8MKH2zXsAlekCCDeCNvBxsd06Cdm0D9
84uJHxZUEG2iy/xOFiVu97X5jCVKqJSe0viFGvenik7Ns/2iU4JTP9xTTydt5kea
MVouKhS++TeMZfPJ5Dvmaizg3/2S/T6E/zYv5LUaEEXKVruLko7WvjJbC5wzclUo
y8wJ+9qnDbPax/J7CMK5gpR8XXoWgivfa6Culhly9a7mUJTwuKwUjIVvAcLEgDow
Wdo1V9fBLWQAkliFP70VNh4TBYNwg/hS3cLPHNLD9JH/TFxPVtrV168hbNi+N5hI
WpontmhCpB4AWZjZszLJURZhFALGgmJ7/mhKNnSJdPS8lYzGwjXjq0XMXV1I1cTo
+sl0pM3DVQolV4q3gUvVnWQCBXr8Wb0uQLu5GXWVzxP8smCBfTPJOI3scBvqbCxl
Kk0rwMspSodHeA1xaOChVfpkWUMJrqnVYPO/J4jGQ8gx2Kn0pTfYtFwAG+0lHJQM
FqtS4a09+r1OQc6DbKgNjEftdFETuzLlkr6dpjG8v7LzL1NKGfXKnmZuKqdRgLrB
mAIUtusr/6zMdIFAi7nC46M1SReH5pPJTnW812VNbvgoQ+hRIKJhMD9ozI9Jcrqo
tMG2lpBfo9iWAKIP2EV6nRJR4IhwoVOTYbY0PzCkNsEt7TxnAgj41ie9IdZPVF2T
Q+Q3Z5EWlpDwCea2oGtb3FMSYgSa8y1/hHhl5X8T1pPHoWn7O+ynP6gOG/U4qNEu
d5xKLZV4DRffAKp1Np7Yeoq+51ZvWlDdpWUeNzBGFTftcyKSvZj+GZIJ+EFu32iZ
+I4Z0L/DNkS7NDenv7oC6ZdbWXokZsY3IThPewq0LOPUEHrpNL8h9I9WQBiMsg1R
imcG8+uTZ4ON0BOECIZrg2LZ1qq1HdpGRDG0/0dAfG7qWCJL5OZEHwKphQa68Jsc
2D5IaHdPXxoBxOg235IJmhgEyGD9LpHRriZOB/PlrbMbEp0178BG24xg+2y70XHG
hlxjG0TQmrtf0T8XEU2aXAtL7dG5JFHaEb8g7i3/FGI=
`protect END_PROTECTED
