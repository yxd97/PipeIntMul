`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Qao6tM3YZnNeLwhYz5q3xauJElxLxeaNYio1DG/C4yTcjXUzSzgbN/YWUDGx9WW
5Exoxxq/sohNkCUKyanzvV7rA5Px9oFOiJPoWaZx3ZJbw2fbFM0WWzNt/AsmfF8P
uTgfNGAHFvwUW/bY2jT/4OrKbRejKsuvmupSczLSZ0EseLA5jVEJdM0Danb+A6Na
p23WYi5TCi2lpIUvg9t84O+J7N/mLcy3HAjtYRxspkaWrue5HDg9ySV572gvIAWK
I4FOHHVvy+fZESfpDnHJq/s1+ECzbVwAT1iSTEfodZscnhylYxmbcawuBdnxn3id
4U+b9F/zQ34RkqtrCmyS55XReViDGAsJcxPBqcyLk2N1+ovts9+uSgWUKKyAPqYH
4vIN+UC+NBD/rfmT3BthWxtCZo2Sx0LCrMUBkwo/+8HbHsv3S90BA1reVFPUqPPH
8C1x7s7T+jKVuItBymiNXBdSR31OdHbQVGk1L9fa75k=
`protect END_PROTECTED
