`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yVWm1KDZBU243hKvFbllkAG0xgpx8M2xzLj+PJ60cxvNBcwdi8KWyda/L3vqsCfk
PYGWEQEdli/W6KuBB3hmtsMsQEw1AAy+Ptdl/KHVJZcdcv2SIZKXhon3rn9D6ZcA
k+0Vgwh6RaeAlVYoediQ7e6ztgNsWAAsb4I8L8ZXh31R4nWW60FWwdu9meMzxSwe
B/dOOjhVZUQSkfg3JoUtMHo2QVgTB1M0hwHgUY8+MLomT23mWfHtMx4QcAaSvaIL
sjhcN+9CbE4Wl1lCBtzzqEwO2As/m1SijnW/MLjNUzA=
`protect END_PROTECTED
