`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehJafDGbjunLrt+oQHGm+M7kQHqu+nVvPEB3/6NejxF0mJ3BIYy3O9gqCrDV8YPv
wM9KXioO2SOKbJb7tU2QsR9rECESJE6tF+8oAhbzYrUL8h0rBHN+8U4CufuXYxGW
qc8uGLtcsrR5TGYVkbw+k+gOhWNbYvKT0EpI/r322WNDCoASdjC8+Bt0J7hh4+Sc
qxCG1ZBlTijJeJNfT6mI4ehH3cKCqun+Ktye41lXRFihxsrRhA9lTX+ojkE4M1is
RCuqAn43EQWQBU6s+iuxcJ99emWdLAKeIbszVqhQaDN+YglvZ+rP5ewcyntSsoit
l9UIeAKewRiv79gLUCtjIj/32gZeaMvltxA467G1fR+VzOgs9jQ5H1ElfX5KDleY
0QQj4bBykrlfHoE4qPMfDYh820Wt8H7mTwYx/emNMqk97WXljskU6HrlnjNg2/yu
alM14geKoyGNPPwQDyQC/wuvAJQ5g3ycKPJguL0qtl420wofoXq0hn4GQJZI9XeO
CvBxXMpnGqzEe1S34oE2uvpvAwcy+N1RNGnRclLhSJbMXOme+CSvFuRH1GDuPDGt
`protect END_PROTECTED
