`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OIRTlYLf5Aci+1j5vW4UnZnfxNL/a5ModUfb+aa4H617KfDXakLvphm6lmcH2KD4
sn9zJOTlRPSOaXVciKWkpO/YdTTrmjAna3gxHzB93xDyGfQAuLAcwW0iex+0tjl6
WFlc+Q0DC8XSB1C/Ag4RZMJRamRvlovLtrJ6QS0+l9R4nF5hyVmRPSWmCT3bGgO9
r/KpBQ0Uu3RTNhYAkjYKYns1V6HxOcZevBb7hnLUrWIycZRq1GbTtRqx8iqYbBJw
Cs29P1OtS6j+XwvL0z74gYv/AznNNy+w09ZJM5Z2Jl6i02YufA84wXGUZUjcHoFA
Sb8Q6oF1BaCyKIrcQpk6PKqo3m9pKzA8o1GEfzgKCtKv5el5JP9Gs1D5BbRbFGRQ
idDz1N829AzINmbdWssmLY2m3QeIpyJjek24YLLCAbpLvq1JlA6Rk2U61mUSjiNA
I2wa37jlb65Kwy4NomE1ioqt0Llor2PgIN9ASZsqcESZbqFSNrf28lsz8H5JrFzg
oYcR1LkUABft2y3Kcf1BZBtO6fgtu5J0nQRGf6s/bBAO7hog5IznVautUW2ScnfE
IAifaMBrN8cmzzF1gtRhnU2qMuHnteB03N8/DHRKODWOhL+QaJ7cjQnhN9uv5rC4
9gpXisa8xfypp6fsvw0bl3DSplZskZvUKXzrcPuQBuo=
`protect END_PROTECTED
