`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHYTcUN4AnqwyhtSQSfrf2ujhHgyW23EM8QwJXnFIAo4xRIM0/xtpMc+g+eOBHq6
6Pjn2yfzUsjOH+T4b/9R5Ke150Bf7uNFyAYMpxt6eoYZ9/OnwkKqMImIcKGCLHN+
Os9bo4PfPC8RKZq3y1UtuzxfHf97qrbfDSsOsEt8BDKx+gPITk0jXdfSKHO19qIX
voZkIzAyB1mCrCOV0WLx57xPHe6YsIXkOH6S0ZU3rV1/nAyBM02aBt20AD7emPjk
E8HLlPBscWfBaD7DwmWH1t7G4q/mPrn2osdoueDt26uUrC2IgbP7AYtaezos70r/
7A+1r7xX8L7ttXfQ/rqI5R91kne2GCitDoB2KzW9mxXbD0ej+fQnNTJCYuXCpCJ4
`protect END_PROTECTED
