`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6kFItrVIpz8CnI+kGNy+KcWckp7b8dL6cJktm6LoIcIp3XmxCi8ZXDZmFVvkGY4
ftbcWBzHxgYiHMPIYAtXBWb1CTdNVotlJd4YF/z1TBQ4aep1SMKRa54hUmfhiWvK
rEzgKhJQE7BlYGX44Z7tKtnUtNJ1wMfDVPNG9ZvCjc0Ww7PfGKVl48TUoUqir0Oo
VlLclFwBM/jgraJ6DtTu8KafQt8aJQE54dvkyTRZR+y/Yl8MthbYx3j7M4p5/cUv
euF47vPtCWgkS8cDSqmWpXOLpJYAEQggsi5I3cOrB2+olt4S918xShtd3JBnwDYh
WvWxjPtHa63esdpEoYfzRiceOBBCs71U0i7y2B3Q9qBZaPQWDBoqnpnqDKGOPcu7
PEaRd2HRS5+tSg4fLQskD7dNCau02SpAMlXEkS86S28UrPOtDt098BZ1k7EIt+sd
/umPwfQIN1ICeEirxnhZKBfgpB6nb+M+aopf5HGlemqabrZx0RJbpEKSv2jYtcfB
mTo9laOURNgoSlN7B2yjje+OdUvq3qAdI3sK9aZmc85rDjjt2GQs+woZXOxs/pWz
lEkN5RktcFj0+b2imx+IATLklx1t86VpPyFNtZqnl1wQRVSY5wOZPXMVswu2famy
Hu3hA9RjHV5Rj6k5t5O7Jwjz8msTcmFMXGrMuLoXAmPRtdDlKn3L6FD2jHficWEb
76/3x4/iGHw0EqD4Ne54TpMRPFoEnHGIM81bgh+2UubkXkHRIi1Xnuty9btbwY2W
eMGEprP634lSRt5MNasA33wtL567cRB/1ZC533s6lJJN/lyYnap3uWNQD6Cp33eW
`protect END_PROTECTED
