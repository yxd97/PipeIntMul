`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FAWN0WvqBt2sKtW8vqNUQXkfWe4beNhPoYO7nPvJ43iRPvjZrzhrLFYgIy7WFJeX
eHkP2yACP/XCSbN+pU/yZZ1ZXOq2x+SsWED0j2KrrIwChc18BEvQgge14bjr7ojA
+xynkKlfvIts2OQNYJGyBHmcQdz85Hy8PqGuO/B1eVQil9YHax64kPZm4bEpJBdi
Tvh+Bl8uwYu8YSTUKsxedsOcMoQsM+EiWvZI+HiqsS+Qc7nk1tSnsZOpXCqiuXsr
1Lut8r6Asm9zUp+WTl3Kf6AsQa/VqlTfb0HJ6bAhcJ84iQIlXhNM/KsHaGSoIDnH
gRtT3xn9p4/ECSCVLVdVLryl8XGzfRwFo5L4KbY4tv5NGhzjdIQLdLHUIhsJPZ/V
0IBJFOSQZ/JCqWk/oB2aElzu2vuDEw8GbwTYxuyogKj3ngu+aghvQWZv7HgW+30y
UBmOqxjLlIcMYqEJ5dco8rbgko4kvAA0Sfw8A0OzQWQn995MBbDoiGEVaumEcBEK
J3GkYuVvMFcYPeKGC2r6ioHlOrgKs2oGC/EVIUFfj217lKI5nel/KNzXQvpI/UeI
nshWIIyZd+RB5WvNIX9lEhX408ejM5wAWRit3p8O/vH5C2/NAcHjVLSbswObfOt0
vlg2EQ6VyzaJj8zEPA2ed7itYs9hVQymLfTjuzmeTuGnl+wmUCEjdqk0XLeiMx38
/arqOovh+MNSDQvjILh/+QEoDkvbGNTKR5Ic3FutOQqhYRMFTFdVQgxe5TGiPByy
ugwKR+grb+NqqYSqVcaLzHsfA6fT3izFKr/mKt6o/N17tP9+RLn17Mx6IC8lpzt3
Ac4WMj0IgGpHOLmmNXD8CwAp4y37cHRruytEaTDl2DrI6hSSD3fV1BLKHygcEPUN
7usF9NhOA137foeIBs3eIpWGX6APUiK4tJjjFKbjHTmWHSHRXi2xwCPRMb0g9Afp
17KOFWD1qsuh2ooqakz9kBTYr+FXgvw/6Hzq/pznaNhkdmjnT3Rw510jdXHOj3/w
Qtlk5eYCe57N2TDW/LeOYm27zb/fghNad6iKFHMy6ifAPKxJxhR5GbiL7pHfKr9K
PTekyLyZGARBgc1U2gWa5kcrzxKrFl5zVKFmeXKOT5A=
`protect END_PROTECTED
