`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cs/m1Z4HvKZdfVv7O0mpb/NWf61xptyu4OFhYKQYuV/VA/aCZbWZNV3WPPu8fzjr
UCuTLcKaUDK828Lujm/YZVC6pm/ZgdVJcffaJMzL6tKZAmw0YEK1EietBOvc8+sp
pJ6OMFSXnz8gnGwdt8gYLCIWGvXi8/sK/RJ2iiruHJlqOvV8RAU/RKw72tZpjgny
SvapnsiUJ1oz4CilKMkAAt6pjMAwB7ohhMlp0LA3pofpgCChz3aGnuAn5LuI4hcQ
zNL5WRE3Jytw+ZQ/bkFkq3LDxSGTLb+rGwgtEnPLl2c99vfIwb2lc9V6Sk6OJP3x
dRW4jp1q1XMdlEf+jmAYlsY4UymfdlSUIOCnTwZmP4+3KjBU1i/4wxhUQ37ruost
gUw+p4ZbARA+l8Ey6S4YK8kK+47mmjVE88Kntgq3u/K0R6Mx3Foxt0vVdNdtNeMF
ff2BK0DZbJhQoP44CZBCq1uQzn9g2ZWYVM/0tK/JwuiyClyRc5BHCe/ha6Dw9iP6
RApyKbiqUxbs6xLAi29p5CKdeUhcBKkD/iemGxY13xANvqv1IRaYc9tSdr/Yysl+
JW513+IWulzRGpbHeKHmnESXaE1bRFDiHiLkH+WRBisof7OsMxdLWcH6UzzHVoRP
m+lLErkDJQzgPLwWfGCKgirsD066ypz2PnpJKBpZ0pUvQAk3Pu5rnDBZXX463xGP
RBOds5/v4ogUeOKwnuKo/4I5jyuJSMJhkZ16upgPBRdFJjMk+0LeWmluQv4oQ2KP
xG4jPvMDvOWuznbeBLbJhcB0ixveYAEYvkbyT6/McN+ZlR0wT4C4QiSjfDvAsc2e
lf9/OAaqt+bDPTsroj0P0yWdxIJfhh4xCWDgRmH3bE2rWff3dCmAU0dcvrdA7geZ
XcWkOyCuXeniAg512XCVwANK4sckpPLqhaTmVRpNte0=
`protect END_PROTECTED
