`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHYMcl51qbngKmjVAmXOClagtAFhoBUUeZ4tmwxFSkmlB8oGqtTu8EuUlPbHFx3Z
bjUv1GIN9/9fYLv26YpMTI4voa5NuSz6dUmu1/qgN++6hK+dmCR8twQS6HH6mPQr
9btsu2loPh+0zXt1FPkzYBgbHXS2vbivvHpk3vm0PpuM2ipiZrqRBRZFZ1kVrG3V
ncCfn5uHxQabfzFyMaqKg+A5PdhCF4oKTYb2L68tvq7slnE48/XL6Y9pErW3oCrj
wA0NPlXEk/cksBNx+q3FUi+hkEZCLgfLdHXK/KdHNU+unk7h+BY2alOj8QLUTJy0
bJTURmSVvrJgyuDnbkdkUqIGAh9XUjcgjTAUUtCLmtBZOryGX73dM0l/f2p2Cwdl
99i5GXAB9gauwKHnqSWTShr+yVpEE2wXXgOTd7Ygj+cQ330GsE8x+U40kHScvkWI
lGv4mDjeJNRXgB/2ZQZ1w8wEOi7En6ASlDdNaUCG0cJBf3Iv3/jFyETxa7Z/4Bay
LdrQXr8Oya3v4dnT8Q9G4F2rkZY9FmowaH3xaMyi53xtr5Wj6B+JjkBZIzap52uO
1TdMNbJdykYPi6nPNBzdtDPegMsl7wivK3y2qYIpxXB21HEhXrfAw0rM9smbySG8
GqbZ2GVMymCUKEnR98nir2yGEv8BTQyvkDrOYIqKnR8inQWfCjuvqWf7lhoitvC7
cM/Vn75vgUc0sPflwa2eScOk7CTftEWPIVf4uwKWhYxyhaWaOqlEGaK/mEqpfQMk
jIYhzrZe9l/WA+WybOI0IYzJa5XcbViQkU8H+YVaLJGKHshw2ZVhhcIRySayGerb
jLoA2ypZQMUJfFSRoTVzJ0CtG/TG9BY/QdvwmcVwQD2Jhs8zZTT1yEnoz0QCZ4us
66eRkzlZ3scZwQOJHN5nGHWTQ21Dc9OJEYuFkw8oMP0u/jHBWm5rbjYmZzyV55vP
rlhGU0oahIkB2Ov7p3sH0Ssth/H6+7GQMWgtdpuYGXqGMWoyXiPrktSa0Hhz3tb5
ZI6b+JCFIAr/vMpyeNJqfXJtiuPB0zdU1DyacAe7c/sb9RUIaYETEtzd35j71M2z
5kN+uhMOtn02cv/WUJ3atjwXmj7rJlH5o+ZJDE5fYddrsrQCwvBi2rSBy3LCO7oZ
4SPpVJWtEc/oHuVrXVuUT/9Z13+gsC/dTz5cbhrOJho+oHUGRu/ycjEfQENlLhW4
HhMY+P4SHLa/LLFrxJY7hINkK4IQt9nB+qskvya/NwDgoHGX6VdnBx1tW/jyykax
Zvnvi1MFSSzXA3qB5TNM6i3QIZEg9I2nmxPX7DOO79F8C6w1CUaVmZoPmGGFNbas
eLCwC0ATpbUw16YdSrPUL5PaEcBFcjHKtzNmhIv9War+Yiln82qpXppYfLNBMs1U
0t2HPdkxTdxhCSJaQXMgX4hbXnLAJTFmVQknTuDINTgJOOx/NXtcCdCX3iZaB5Fg
RqcBIjUXavzl0NhQClsfT01pohE+KvVyTlNla/tzfRV2sMyWOgpMwNqW6I0hdWVV
7Q7XQljfM26fHovpZeEku8MpkPIRCXRueyugABvUmAVhCXAyudoGeyasqPZqmSC+
jTmQayJCUwOTKQ1BIiQXKdkNogZtcW85OBPcBGwJWe3ytExZ1dgwbT+IbWYLhb+x
AZRkO3od4AXZldooVKoSCSAbgS6eIkztyunJHUQtsypVMZ1ZoNLU1OcIpc2n6Uhu
Fn17hEUdfXg9gyWksvdFVhbWxeWLLMSWkE3PMgMefYvvVIsHm+YfPgHXQcfjTG+p
HB7LSbca4yeExFsJf/we/BIaXITQ7rlL/2DEDkQcnolx9d+aZ+CP55thLAiu3VNU
lkovD+AzR2JlBaSuPnqQSWRx18Rv+SsGpc9+YL6pOsjTVclXHD/+pvcJ4BO3GyvB
TVNMNW3P02lmeiyZec/cmmyRTSfc/EBfirZwgeJevEogVfe49yAPRQcgu/BuCC0I
rnbCI5qDGLthz2kY2WaEHhLDEjY/ylBSSKEznlAOxFzT4SQkvgFJIHv7m+HZO0o2
TxOFG9cPrFMt633AdfsG6pU9ULHqk5XLKM8dw9SLN6CroNA1XOpWLPJzPr5fDapM
+cOw/GPvj3cgdfi3kRKIvoBrB4ZnXaQSsQquPX5j4lM1paaYWuDQWF65DigMiE0O
OZgYcPw/BJ1rhhvhUABp1dni8+WK6IU2TneJ/UURXnqoRIPqWkoksh9FcnFGNHE0
yWTONxKfhEmxZRCuF5QzcoCa6lRSA+1tkQ/vNtztYZ9lVvA1ZGlIYZgrjoG+BEQg
SA/9wYv94KZ/MeY6yTRqXKGiDvmnD/T3oD1JT/j+5YJXp8iKQkmDJZRIONWvKNcZ
zTZIoknZ4hNkpA8Ajq1b8YBYkRzagfbFpQZkv4menyCR8abxoyAPopCMcYY70ZRb
+mRgJYwGY/E7MUrb1WEg/4Bsh0j5aEMf7OH7CljBxMavWdA+vrFaqym89Z8AePOs
H0Prm9lTZfPqDo1/OJmJv2QdVQuKX788FynNqVLXzZVo75fcDht5IW0XvwZIgW6+
RfnMHYDY/xAPfiLycEJM7fZoe8J3Ky6UAyuyBHwy7Xg=
`protect END_PROTECTED
