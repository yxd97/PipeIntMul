`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78D+z13a8bHCs8mO5pSJHjOkzSAmjS9bUClC1mB7Sw9K8Xg6CEFzfpuy2rcbycV5
aLda1AvHmLKbNx8v0Xfa/7f1lLgOBsYOkkh3ZQeHNS2ijK/Pa4BTFcROdS1fW4S0
kUAP7g7dEjG1J9vRtxht/4piXFNxxjAlrPc7niWCR15zILfk5l0DVdHdxgYLWWez
5903+8RlWy++4ctioIl//BCLxVgU+DyCwsEQvMAyjBUG8KA9+VDVjdLMubo2Soy3
KEMNu5XAjrSiaxo12PXlNdHxSOG6UblpNe9rT6L5SnF4l4Y7ycNO0WH5pLWL814j
jpxTp3/ZMMw7QR3S7ZFPQQ==
`protect END_PROTECTED
