`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/EXfV4SiDsoWqxiCC4guOmiuiNFcfrQflEHar66bcyxr4waKbnVyK3iot9s3M8Wi
wyNvTNm1TfiZWrp4KCbE+4agfHaMPwJEVtTf9Fb86TlofDc8Cavtsy3GYHt6vGcO
sFBCDG8mO927V+wGLIds1SCnSSmlAG2uogH3ZkiS4Pd8Dl1pbFCVrcnVvi3n972G
+ZP/fZShZSq82ZxIQ2F/HQSSTRK6QtBzQKjHxrJrD+n8N1e07yyzuS0seB6fS/52
ai7xoO+fde+VYX5xqqCfQoEpZAyfNPTHoccTcQpQEEgSP7dd672+d4aWjsOoAnwM
c7MUhE4QrgZWpbIEbjv5GQ==
`protect END_PROTECTED
