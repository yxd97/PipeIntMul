`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YC/V6FdNtEwBURm1rvJv90TgZnVIwsoDFGhZdgzA6NM9cB8Cn6BJAJ/hKkBz8zDO
uw+4eBQ2Utcl9hIS2jVHXPkWlCOjo7vX6udwELa5MQWWqRmgf5NeN/uvkm8HpDsx
p7oQ6JB2hLloSeYtZPcPa1a18BKkhS/eJt+EboHBXolFi6f5yE/RcC2+L8HiGs5a
UaCJeaiump41TRnLwjpHSZLzdrj8BL5/xF2CiYubNZkFohiXYfvnsKu6nBIP2dCw
p/2gr3LIZFb9rtDFpe8DGKOA2FewV1+FSQfJxbC8XfU36Uv+MBkklETdZdgTCfAs
ZPmBOhqmww6eOsViheYtBDc4j3FbDIdksf6zTLjfNiWazoDHfwf4eOyxSYSACRer
6RTm5LGFaSTT54eAyQnQncKzA2G4eK8+pYNJyX7Opu8laDSeglezLE8QtcNsyNz6
Eabk0PvLJ5FKbUC3Aaelpw==
`protect END_PROTECTED
