`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCB7tcJzSLjEQ1H/OeTh1KzgfyrWzfbQx1oMGc5+Ih0OhvKcA7exZIFRGiJ9bRhF
71vQ6s2vSwSXPJQJGmJB6LxAzvdC8YSpQNElRWqH0IPeqLA1gfBb4jmUQsLIbH7A
UybDTBDJ/5kvr2rKbgHUPsxb2UaCculglhE+n6DTEv0D2YmQO7j0EHEa+9JPJoUp
/w0A2pA+oEsrYezW2Flj4PxGxbuAYPI3NpAleo2IJeZf2u9GANz5s/nCJQ1qz5Uc
1TaMHU/tZZfro4/7djOFts4vs1wU9oFJoxlvhDeIdQZ4nHv8ZRUCRzAmhCLVn8js
yh5L/frHfm3VvsZ3j9nQ45YBK4Ep8nfw4X4oO4A+X/OG9f+WPZcPsm/JB2kLx2fO
+2dCQXSPQHT5S9fkieTYjy0gX23PAI0V9r6m796Dv919gdZldjgF/8RusRySWkey
4VwP7oDVePPZN7fcvf2oNA==
`protect END_PROTECTED
