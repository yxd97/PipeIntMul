`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsLb9WZKMkQu8t5+wgPAClRtKpdgr+sH5QdrGUAq5Nl1Kl4Axi8mftl+xgLWopT4
xSXedUEG3+LwUnegWYC+OKDpaSDk3a4sLJvjyXQhH5a4b9P07E7qajtK1u+Ia6Ix
y+QYCsMV/ADE1DSdGA4+4d4mkJUmajMulIQNcOA8kvBHM4OOPxggCNwO5Kh+Pv84
gPSuHEhnpcVkeB4BaRHIrvCiHsvZlDsTeyOCFtJNZr96qzTZSo6LypGumUl/LUyq
K1sBjtRv93RbLijd6pBYrGo4bDan9sdPCR/YQb54txlRadreQrODw3fSFICzY1ti
T+RvGrHwvE1sPVZgfrPT2OcCSn42wJdKjRlQzTM7+GsZ6fUQrY/w5l43ASmJbe7T
`protect END_PROTECTED
