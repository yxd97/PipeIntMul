`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B90a4lj1Ulx8uxCB7703TLiZhLrdGU7xyX1ImwL3h5cEJaq10hEIRDwr9i3zfQUV
t/2U+pGhwV4s2RSptk4uYR0tHA59LmveE6xLDMX+o0K736lM6Tf5//Ea+LvRj97t
q2yaj1YS1Bll0SygxwDGWMilr1rFf4VJQkPD9fQgGkPj6EuCn26WLPbZfRGliKcU
iUJqNFcy6VzplQ8/lkm+uptkMJFp8KdwEbVbmozGsF+uea60gpFXTWnziiEpIy2o
2NQGW+WKWlmrnXGuFrGxqCf1ch28Bt6Zr6+mglYWrqTY+8QZxjLJZiF0SnKGG3UZ
89ZnkjN5iHf2KnVgij+MgYJlsLcrd2xrU/O2fycIUlh4sVXE01pt5nqrs4bw/N1v
HThMGey7QL86A0ChGad+pBtzUz+Z2olL8WuvWJIHBg/LJrIYW5rGnNRj1rLaXPRv
uIcAPM+4L07PtRemJTPJG/UqnlkVl+7wbwVVrOju0teMj+4PDnQS1v990rp1PDSo
OpbNxbBJ4tGjUj0LPO25enm3V3WbPYHjmwi+KmTC8rOzWIUYg5B1Rfj/RJxHD91A
Q2mAG+pqikrquaCvEXsdwfaKPGmRdisqc3SH4wTWPW3hTRFDbOUPPiyPGn1UipPY
DT4XNalz5bY6gXBWEifVPgKfwzNlK5r9YGsOayHTlybTPaDg3x1MOrit2iL1i9y+
3V8fBmVPJQ3BL58MgjFsT15fp5OgWQIFZJwv5cQqHLw+vTaM6zuAxtB1OUneehO/
iDFk9NTSLv4jael1jJh2LNmnlUmj/U8fzqLwBhLNeHSYWERPfWoN6NzDtfgjd8GA
/XDfuE7FTMOe5TI41u6gDNmB4XNM9/JNMrwvarhIIusQVPzi+QIRw1MfMtBoxFyZ
tUyS9e61tr9/9CDznUFgl9i7tCv6feQKdA6f7061G5Q5hRm78xO2o7tY/nYZh+ud
f4/fAqkD/Sf82rGeDEQ5usstrddMcpNWTw2CabgiMVcolTdFBQBGfSYeyNyqHCUg
iFzGCDFN0btSYXH0bVzUQKJLZfVnvKbpH1jmg8hqbsX6njQ03nvUdFN/Swpq5ztn
r1o0wc7OE9F+mLsDkct0dvWe3avK5xJi2EI6Ax35FpC2VCOCJZT/MKzXeZZ0chtf
lbPlXLs4n+EQffrc/b91NV3T9GHV/X/Zm1CtXgdCqwsaqRqJ0OqB2dJsPx1L3O0U
A7Yef8UvIp6HLY0uMNaMCb07AfZc7FMvGhnRg3rvu1GfdNagCYV6CishGHBq3hi3
1wk23Aw+4bNsk6Tf7xNj1psSUyydD75FXUoK6Bx3muDThqL1KPl9hXdRJDye8Kcr
3d11qnXDhKGdoUo45h0Ih02MD/BZzwgJxgm+gluZ37lr52+p7u7h+bTAnE3/Gc2H
zjZws1FoIUnrfksMu/TFybHlA1ODrYlc4ag+xjkxghYqXM+1MMAcZUkoGbcYOPCY
9tdGSKtXocK8cZi1En8UbNuKIx/cNpwyuL0OyxcmAu0MbOmh7pZsjyYy2ekxncIg
GGraBFkHXqEnv1lhxnIZtWGXznVBr+DoXX4orNhHxABwoovHDPMhEzdiYzNhaT/C
X8MxKGQTS6Z3hWOpfBhJ6RfOoiIAhK5pvXkJeNJFs0bmVzPSNj+LBqwjITExD09j
amvmQQ0S3Xz7moy0pe9Mv9URPpcsUny9+IZXVpzUg7qodVz22MsOA4zrwxrERNR+
vb3GUZ1Pro7eWLPKNyg9lPjGfEuFSGzYq9f5X7N7x/GeF+Lc1J8Wja872e3yS0Gs
ZiiRtwIfqjFPDD2EQ7Mcc8cBI2zHGkhHEarThXxJ6bdu3iQxzXq+k5/JUcoJbrCO
UVBKsZdaqhYS/zYzfPAE+kc+EpbmYRRL7p47mbKNtU4RiemlppWt/GKc8oS0GZ85
QZ7zGNf9B8yaqAeSL4FRcBnpL19RwqVMgJbUCdz6QddP1ig6zWx/5QQpCdsO5fF4
ceEbDk1m1CyKgdB9rQqvfpqNUMNyufJcY+9WOQ0vdfzYxIPkDvIo5JPfawByI7HG
bhkPwkIHfQPF105fmv4KFAYRes9IStczF23rKZ3/hIvBVD5KvTiVO5Y3+87ODlge
w7lLpr71kQ9kBrapDPGGGpNDRQPiNiOdTUsTd44PRAfV+CtLTdGkAN7LX8NS5qRD
eDzuPh9+px+Y0MtaXB8PvM4y1aVs5VMM+YHnat2Z4Dzcg3LwKakxEQg1ldWLCBIF
GJwgUJDqbHs5m3jFNW3pjiotEgHoQkPT1YypAH3AaKT2mihgiMstk+G6+CzEQ0e0
26CdC9fjDqHBscnHVK466oHpDlxoNJxoZ/wma4z28kw4UXW6hYZI5S2WH9ToeGYo
1oXJqL+wONWH7qZnBOLNl73+UxUYWJ3fgsT4e7Mqs7vBzsMXx8YjFiYsgEePD/pO
h94hSzo++jp2TlQRJ/owZVPGNINXxBBPpq/zyTFstBzcBcMdQEc8Z815aZBUQQqx
CzYzhWfZSAdos00zglHrNwMNcELDoTcnXqUe+WfrrYACK3HbyiSNsWwYHAWxMZfe
BUgxL46qONmhEV0RWaKKkequF1RxZKVvrKOO+s1R1QDJffKSjSP+wp9/e0HLhHLE
1TE/5s4RZ5g2sgrtvsrLQVSEcWym1BbMS9bp/EvsZWQ+xWvd8cVMYGWDo7fLAHgT
GhnsXxI4Wu6CByuHKbzP7eH52wfY4I+dGXBJ27GKjx63zP0A5Pg0uXc0WbUdVoxG
2h277VBw65X+wuUACAANSp1oSuk39BHj91QKgllve/YpuzKCj1eWvQSj2Tb+/iq7
ug5pLz5amAoU6P39a2LjI8fgvZGLE8noHFMWsGGjwsxyVObjXt3An4I+epCWH65e
KR5HDTQliNUaqPiUIunAdezLBxq/FM4hNbv0dqDwcr0fmH4X4cEQZ2ofPGKDMS6W
KhF3Fe1kvMbjugPwHQsNlz+lV1lHQterlCAzUE8nZhcSzyn3odFoMjGkf5yWbXxi
oBRUviXk519J3DNu977A8x/e7zFKWmHHSIfViOEPzF+oYVg08Ehhnno4SrVF4wrj
afHsICyLSv/IEudgSMVftF+gs6gY/b/+vhGC9KhaGzu8eLkZ5FyrQQMOwzBO4KhJ
c88ufSrhve0wWmLAJIYybXoR5Lx5c5wyygOvSbzh+F2SUiCYHkh1mznRAmXwOHTe
CtUtJvvPu9xIRdHasNoO841y+0QjL3nH/CuNkKCWtzo=
`protect END_PROTECTED
