`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFNQ7WK4LY7nBeuwGCiKTUqSHH3I3Gucpa3PXk19s+84y7IfKUiREOZo6VjiGlRf
NO0YuhxManWKJcZCoi3BCqKWMvoZ8IT75rDzERDO+XlJCBBAuIzzEQ1UCZXiVN2q
sMpVGu5MuypSIdlNrxdwr+YyCKAKB3qENESohRXzpZuJ2nXvI4TIMJ0EZLgcTKE0
qBrQQdXl1KEokLdq9OIE7dATSJ53xAJmhvjJo8kdGSsMsWtUihEwnbyl3V+50v9z
zTV7rYBfhlIqUrGJy6vnWCivajEG0pAM3LMq5hKIuNQ9E9zsUIDBO96s2vIHqIUP
03a+sfNEJ5uy5+9nBZW6H1uN41mS7YnodAxAAmvR1QJzwqVc1AH8EI5gc2j3hKZK
BQLAp5Vm7/q/GVUxZ5My/PyKzS/sfIsdcN8iYc5dSk2YmJZ1gewFTSqHk6RGTVJQ
cUfKyGF5w5QQAqk6xaf7RGgNL26+RhDSpy3o1u11DDY980I204R2b07ixMzRbYNT
37utg0DW5znoaW5/vVtAcd5HulVW21EvtW8SXQKp4Z6mazd1RQtMNGAERiwVVGTe
T8TpLWDH+ZwS1sgBWX0vveJop6/iIufPeNU9LwqIXb+rBloh6xac7ZWsV/pAfF6z
`protect END_PROTECTED
