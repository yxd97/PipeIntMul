`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8YXaqjxkQXbv18r89XoMy6MM0Ev2JyYW0i6yHniPQqqwku6KrlIPdhNsb5eroWoT
9OykBJIF9kHJKC6lV+CQp96Od7qXoi2Vs+rgwfDUT3Mw7fbeoYLk2cQChum5m7PQ
QpYOPhUfU4W5CPtfqEdmv+jrVpFNy1ko/YjXgQ+IZsxcE3cI101Soe15/l42HKXr
8PYW455BO7XpPNF88LWqEhn1xalq+rA4pazqPs9DVrECkXSmJLxRZ7Gtk2Au9OYE
Rs5gzUoaHkFQ0xI0mYuofLykqRe8SHqKAHj/H48Anjelb88i8QvU3YzbH57pfncY
xw8IHc1mDNq24E4mqxM7QLjbR9iKvjvVUPBvK7tNoWY9/KSc1qtkqxjdTsbRlgNi
pMNEQoaoJk8BSYtvnu2UZG1gi+7hUFKkgZxCnz4bN3E=
`protect END_PROTECTED
