`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKvxrYk0dUSvaNJyWLbUFgSwRGvzS/7Vf26uOgFEGbsuOi6WNMLQe+Yi7CuwxZxF
GB4tcG9sAAUGfg80tMBKWQAAB9NxGSgN+/3J0wj/tQ/l4xCSxReZwsbeuaCzEADJ
dJG/rRqzcE6P4VQRekswvAAGsbD5rgj3AtZx4OgnlCHDobu0g30UkfnMMQgurkZu
cpvwwQvdkqxcaxSganDJCARqvlOGgLpDy3SKk1BfgaJO799J7JJYtRkhp9wjEROM
kpjH8q89TxEowwUoyneqlapowCVn5m8gXzvhIh7ROX0CmMg/QmLIXv/aAtfxSqBy
j5Rnp9YfjevSRFjlEbD0UNyTOhHBP0Ff/d/zLn1ep3M6NH3TvPL6NEj+73FzNNGo
wb7laXWomynJvWqVyRA9aKZjwyELN4ORb4+8+nkmFr6UwT61OfswPD93+Zf8NVmO
FePROcc7VttLNL+4TwVltlHvVFnbFQtMtTcMIAwCNZDAfdwMRDsucmNZ9HWrYhzd
`protect END_PROTECTED
