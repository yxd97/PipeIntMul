`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cm+8mYKmWTUznKcO8stC7ClZlia+XPeZv0xyPx73k5ycqYZY2oiHv7wH1ik+s51H
JNFJDnPspWccNQV8jQuVok7mERdNzm1WoOXPlhMnDb0Wtp2RtgvJCz5+4ar9HWDl
8dDv9SDEv0y/8nlNI8pmuqSB1iJrG1K8hDoccjJ1VOdjshM5M3hFap5rmtCuH4V6
UYwWqdHr0vkdcfCSYcX7a+SECpBg5IrYNu1yjg1drAMskr7EN4Y4z18AtwtqP6Bu
s7HOklAxrSmrrOKbWvhY9C5Oyx0rC3Xoh30XDypOKOq/RxvBlpnR7afh5tD9ir00
X+7UzLTrteRG9XEveu+1WdvpJW87jCDRme8AfTqEY2cpoNz97J2Ou2rIE5iS/4A1
mGGgmhKdFWXF6xpmGvQqgjvcv5u8umpqGt1EQ1OFY6lP0DH6H9NclhPSriwe420L
CYpemo9bGxH7rLQwbISk+HMiqRGvSjvbhkrdqFXTDOk2r3SxGqF50fvranoE5oVV
+8xjtChqxW9AJgQFX3aa0GnwppsLy/G5oE7gREPl/FIIK1KbydaoWsBTtbgTnwsF
j38k2oemuZ55Pv9tK2OVAnRpMy5OJNQIoH/tAQtlIhMSRNU6mHbpL+ytSl0wrs+o
JYEpVQKStI3UDiI3tcJV57hBJybBT5XMUqdHXMnfre3Awjf7owig59ijCMVoKlZd
gmfqU6raC5uwAu9zJllz2GrYQcjdxh4U17G1Bncjvka9IHHMb6yHWGX0UuVXz4A5
zgpF7i4YXWIOL19sReEn3o0yJuuSZpzxPKX9IoS8rPQXY+kU+PCOJsiY05MLOuWC
4Hdb20f9QALj98e454eIjDuPLMVHRk4M6aEbIlLNyneXZ29JUSZEPLs5yECsXoLj
BJpbjqb94h5z2fR6smTP5EugFR5hpofSNtXv5jGPwQogyE4WLG0U3oxSDKsYgNdk
jXDntqQgnDK52RuDIy+Xtt+Q+37aupJdrnW3XzG2MVSyYaPR09jFalsYlH2ouRpC
AxR8iXzD8PfelpU8WVf+cDwEAUdcmOpiVp/jO1sGJtmPICqBTTnnv3SVQBLvQmh/
ENyuvXYcDHP8PlZQQon/jEzhMeWTy5RP7FyxziP8hAkGkAD5OPPqVwlymxNHd4g5
de5ka4TO0gusLhbkJUGCaH3bpSXbyBcsP1YfKoC5AqHcFwdxX2rzIrIfbv0Go+7z
dB2oo9C1GHefd4jS+FJSJEgKyIsg9LEblI0oNGw+QwIc23lNGdWT6grZBUiyde4Y
2ip6Q9ymYeUT/k/ze72Cm3nAJRzhYS75q3OrY2tLYbSoCLuVZGhOLPvXl6Bih/t0
ffq9hIWqYzVpLCXmN4ePoJ4bgzsQuvJLErIvU8EOLUNvp1MnxaNOtXk8PfYTLCaz
Mu5sUgmb6zVfau0iGbP8/WWQeeb81VPB72raE6ot8mpzqYXsddH6QvIQ5uJWqhD9
tTVAIy6LJbQ/ouFPy4rLQaZjSHS5ZIqmsG89/YwRLzXWdtyBl07KD3tN9Ym5fJwG
PV516b2Xorq+uahZfvmHM5WFtxcRC6BEoBL/ufYGuuV/UVl00SG4gzUNlR7TLgQe
m3RjctoWt6OLPSIPcYANi5tIoSER5ASvAkQKsMJqdV4+AhEhPukcwaTxSA5t0Bvs
j/HQ8aj7bWkHly9ZunFet5DJ50scRsyYx9h9kAw/uQLvG7qUQ5AGFoVyQQWT366v
Rw7IttHPSyFzE2cJTomo2UOJyp6KHyg3LhfX8yw25WYyrPDENFT5Z9OYwFUvdxgE
L6Cz8XQcaLWowzkqLG7vskHo14Nnb5/giOj1N2/9iHsqdznZcDT77LYPsZZ4tA41
B2EWR5rQRRkfCSUQ4tieO60NazGF4GuaQbbg8bnP/kVUa//kRJACNXu5w9HBSSpn
k2J/ET5gJ2EejMZ0FMFd/f40NIsPL7VHCk3E0YjCrB+pDSmrtO/2k8B2BVYXBW2l
EovvBco3l+scQdwwKUewovkuLj4RE41pDr4jGmwguCGQlX6V1JbJ5xMc+X6R8S4d
NmnAZBiz2jRefP+X77V7dVTRvSpYIXfXOqcNhaBxTRbz3+44Aa9h0wq0/bIkDl5B
dmPhA3DgJ8v/rGAg1dm4utb5cjI7sBW+xLg8IhNPFyRtuJcmhhif+AOYQJgAUAeP
bN7mA1v/Ewrvy98sSm8yXu7KxAM32e70Hnh2lbPaGm529cHobfYGLb4DydxfsFVb
+VOe08RIMYVeubb/H70UEBOtasWeqcI4RYo6cMJSIdvYwaog2nVSysGRAqAW3YgF
qjCT9G26+5kKEDH5wy1UCQzTJ866Geb7NqQ1L4eJVSbReJjZRpMHrU0gcXVLBwt5
v6BlplNHLQw4/nUhcoL5Q0JfziRMkGyVlL/3xrNNVPsAHa6Cmjzl5ZkIjgQIWA/y
5i/iTkXIVcGsWlC8yxYq4fm+e1jH9BgozRgaMaGXWqrR15chlsi8LYcsJbPSDiHx
nOVXjlwww5QsSLag4weY+MQJicPILHnQ7XF0+APfh3NhmxEEU8cOxJ5pX3BgH4cz
eqY+iV6Y37RoBbCx8usoYtEfZDB1DkjPGesZUfwi4asHUa9zpLNYC5B3kzMGUqrx
uni7K8G9/1Bs3QWnt17hEJudi7P5jdjsChBcCkk0xeNLsIeMjFSrkUfr5UGrdaqe
cU40AZ9+QJQtzPhT68/Z/2D3sEwdCKD6TI9745OwVHslGxUdLIBV9iiXnPgo1ASX
U9nXaa1OLKyXO+zLEhhciiaOpU0FFe6035xKo3w6aiXElv/OOH1onsz77vtaVmhW
CHjVm5YA110YRhgpzyVpS+4STPcGN5OHq7v0Yra8GPuXWvsQeQ9Vi/u7eXwT2I01
euelcZz+Pew/BV1qDC6us58PznGGV/0/l6BOfWvrozL7oAwaFRufm8XsRTswRkvN
w8Nf69UBPe60UNu6kugSvJ4DtljoLR1blwqIaNIrwgXypnmTIR2wZUCT0pVxxl5V
rScckpWxIopqnC86w2Kqjf4tzuH7IsxvMPzHHNfLn7H4NlVDX2CDixYx9OR65Cne
fkUNSuSNCo5Au6/aCeDJy93s0gwgm2d4U8VEdvwqMSjoEcdP84+fiU3ITer874Iv
rYfh4JJ2P54u9NXOHbYAkur+Tog68tp29v4BIl5F/oZ3q/9HfGJc5pmMCaLiSzd2
6GrCDTn4bPFoPvkWBlCaPAWJhaLt5fYbncoQDoCCTrXNV+Du5oOk/YeUVXOy4qj2
otjglsj0b2htnPHJ4f8U2eN+znoWpQhVOdIiZxoMZ7s8Kg0zo9rObME2sqxIGgF9
VwZjcpf0T0rAMKyJsjHvpmEJ61orGnyhRaSRKpLtqBBPghWinW4UCtSiIBKDnaZL
btFdM1GnBEFbWwiW10ptAHXaYZoQNuDESIZh+jNuybljufv1E0H05rHLK18iyBm6
v2ye5EjxhRhxWwXPHta4vg1zAbF1qCsa7MLb+olKXPg9h+TmBYMVyk2hByRwAwmh
AItO1AUCDjqVvzqKOcTj/p4uLkSSczphtoVJ3+ri2yipBpnGETVtNA51DO+GRDz1
ZruMMB5qJckCiXDvbZ1gGefb8/aHUjk1p3+nKnShh+IFR6vpUALNLtAmIWzqMS0R
tcneIJ2yGTiIV11/Oj+h9xk1pkDtay/XMlYAag3N5JlauXZNgt4+pMNKoL7IcvTd
YRbvctVUm+mX7RRyvFXo7IjB7/Q6sNMCcHWqSfxFueOM2kX/FNsRF9eJ1owe4vib
8E8oEVIQt0u0l2qLsoQzzdCUqZo46f0P5GvtRLpC7KOdIdJXmt1fOiR0IzB5ZRqS
ueQjP4KXX08W3lnMafBFqB/kNKa9w58XVL/pkZcWa3sqQRAF/I3bHSf8I9wAoVKp
NZTE/Ki1hVV/5Ul2AzND2uediD0ZmgGatswAFoIhK6mfHJIQtu9MiL75nKaJEGKo
0DVg/6hMJnjEe1kz/HsKP7ZctzWG1cDDvGeJx3NuEiW+1ofjtOU+SADKdkbrpVaK
tFXjm6IxMbCQJoEGLEWEfUppoyp0iKGs5gTzAHgZRNpoXmC2VPf0ijuQ6wcF9wcJ
7a3yutcnBsZBkIa1vX6elXTM+ZolW0X4kMOtQ9W1DE8DVK51GoTnbmStV216W01+
m5nLbPqe2u4VSxDVcjmH/GU9vh5nrzy4Wk+io3fz5rKCccacsdveUBYrJLw+rjK7
1EayUpDU0V9HzAQ1t0AWPNMekMyaHffKxj384+biJqU=
`protect END_PROTECTED
