`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejpM3T7sd9/lfPqZLxjm10OnJhpL9rnYuDls0vHivB1PY5SbWkrOmwU+7IISKp7D
9KS/mZGqfVhZCx7XcrhjxfNiI5BHSliBveILEWDrc2dN+IAZpZLGprnD6nAKYXMS
g43oI0KFXflxwEZqKQL4DRcgGnSxNjUat6//K9bXeSJ89s53/4tNExCjQN4YIDDL
I3ee+4MsqJhNwH1wlGPx2CWGaY8ZxrsSUyU/QI+LpRsJbdstJqcyY+pcaAnaiBvD
m3FRsMbmrbBKcYPuxdSjQHg719MXBg6fptiNaLcrvuvZxmF6taP40QRpPwx5hSEP
Ovdyz7AEUn9+uRB2v/akW01S4gMeMtGWhQbb9R1ITd1R4+usz84kEXcd4APkeZcY
IH1iq6yOHZxwrDRhaObWnQ==
`protect END_PROTECTED
