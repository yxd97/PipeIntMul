`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhsRtLD+F2nz0O5Vc/KpulxR8hteQwawlu/Xyc8MW1VKWrB4DhekWaErx+a4FU8D
jcgTMAzjSMuWBVHmaNfnk16S/Mu0d1Ri2TrB+LKTPHW8qd62kpl23ksed2Hs3v/o
dphP7GkKNDVmXd/Esov3jla1Mx4bT0EZhWAn5F9kOzt056XBt1nIkdlOyRhtr+Fy
XtcpBHOI3a5NWPYZkSam5fBcePpaH4P9CrMDUWRZLFJO0tsJd/ak/r15UWfuqsJ5
uDvCYFsjIuXGtOCt2NzRI4qlx1xKa6+tkmNl2R+eRh7Qx7Cpkh/MIMdfjPoqqOlI
9uEL1v96R1/oU9EQpc9kfjpp0O982UvxviLj2x+0EHaoQxSrRLRiyiY1/HOsVjsQ
WOpg8xhWvjf3YZ7G/3th6kmIa/l9y2tKb1n4Wrrw1MLedXQrPkcV8oKZL3HGDdFf
OyZY14AWAAqImuDQRW/PW/ULHgps9K7t0+iS2jwohuxu8ZpPl8mfqwJPpvZ+C0rm
98UG7k8VQIdmIV07QGaKlNVbh3LNMDS4o5Yi0f4rEeW8MXG/y4GOitoxZKGiP+hd
k0Llh+EVtXLkUsQS8babStJmoq5sNsxM2BqWhbSLemCbMz1j0eob/W3TFVElA1Lb
M7DnLdz7T++uj0VfiPWXytrWxaKmuCj9ypMjRjIQcpkjt4+MPmanjkZp9jrTiH7l
U+3V6WP24Ik/zqU/RKGXhmz7fall4ntC+r7BoUZa5ivI0xKEWGeGYbisYtzb9N1O
6JkVnlqGGXRD4PtQrshUK/LiK7OBLS9gIJYCxNKYJ30uSsMfkbGiFSHzK8QOR4kM
D8ZvUwZoi4ZIXPaSapLoyy6ndpZjRfGqt9i9YqMEE/0=
`protect END_PROTECTED
