`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WQnDB2q64SXdEP02tD1j6fxtu2KwKX8loEMNadRqObkB61cv5ZZ6xXxR2IvoVLvh
6z03M23OMb3UD4xnThMY18PyfQl8g3h+4Z7LKZqgn64y9EtAS9upI6JsHaZZvx7F
7JHIwbkk8LQ/k90GnPkZpQfa2YiSSaqYyQDjSIvmkBrGueAEXTAMTO3DC1QlQp1X
n3zXQNxDMNNoAsLun5bmIsvu94kRf1bMT3auTAPeog/VebFvFr64DlGkX7lz+nk8
7V+j5k4g3vNHNC0NOg6mc7CHL8RdjogiiKKLY191Ei9ZVSjNMyM0MRe+6mGrlfin
kJQXz/EQbsq1E3KqEVhm+PnNjPYe3nQEP8Vk4M8am74C9VLlYk4d4S58BGR4QpH8
LRkd3Wb1Nz4R2BpEISEG99bm7QylqqurmvaM89pebVUVydKC3rg5rRr1+Gn3KAH+
WxqUn9P/8dch2oQA3UMuTrWeXg19V2BZk2IKJcZBtKpaVc630uMQuPwkUg6E1lMy
T5Uy55XmPfXdlf8/NP4/NMIg164wiCMjbM9Y0BThdyFqVTUlCYfOY7Pk9H687IhT
q5TxsgfFeRVK/pgVYymgwC4Aiabc8k1bSH3PRgbEIAtHrwCpptVJ/PE8v42d5ek9
9hKimGnQupBRh06uldziq3ym1tRMFJ8Y8EyVkh6qNN8sqf+GexP/vVAcfBXi/vig
+iKufGtB5DmNj4+ng9CTRA==
`protect END_PROTECTED
