`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uEYm6GOfT8jR3tbzW7XvJ+cgF77BvfB0Aw9fg2vGWQYmMcVRg3uF8L0pd2u+w5A1
JFf2mjOHAyLzbO73Jabq6Ywfq/KYZg53edZdmeuDo8f0UmPg/OMGp/37DVwQzCeb
U8URHoln4yc9sBRPfIT/y2w0UCZ0oY7XXNqfkvA4va8/OFZGqrhu0yqg3BNTiw4D
9VyzDN5PyEBQ6MaVJYNcTg+4BWygjup8NXcVfsfVzKcIXZTtzGVpSkpaMi2PjAtW
DefZ9G9QvdHW2tRa6Gub/BAVQ3+7dBVEwsEWxSRr37XHGvdnUPd7l6JZ/H4qXZsx
61gO1V/EX2RR0x758OdF+A==
`protect END_PROTECTED
