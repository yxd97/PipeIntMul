`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DK81GFPW5weVJjd8zaLTbGaGrgeG8U739FXEEN02GS00TjEwtxSKZ0LlBdARYExw
otpg2qVgfOaR5gBD5XMawNs2RMFDxeEfLfnB3qqn7AKHF+pTQUo1c5Espp38xFgO
K5+78u057wUaw8ZyGTd7Opf6ZQk+rgovuRouWV8Vb/T0LeU8PLQrzSrBf7NjjVYf
2I5EiZwEKO8wI7lEEp7did4yByVPfTGz7KzFnU5TI5h81wgpUJwk5cY9UDjPjETM
Ob72bz2jYSX8OgFwdYCjvsfw+xJ5IBF/AkIdtfnlSMTWYzTIR8vSIKoTa/Xeo/Od
Er4BKZh2Pve/WFA8kIxLNg==
`protect END_PROTECTED
