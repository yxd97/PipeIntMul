`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i95fTusZtKx0S3xrnJ/XRVVKYEPHPc2m2zOBdUYKLdP5pCEaooURBJqnOriGLq++
k0P2Ory9ImHDozE0zK5xU57v9A7UGKhRAjGbf3smDMX2CXesqTO/4QhQXVsx7H71
uZCf8SK4Ck4DQppkmORmEHJrzmgs4BzkrK41rBkNlphcWVSjMOS8tps/LrZVqJmH
NeXp2DGDV/H4srjRK1rN+CqcrmHo9s8ej3edij1T6oXhsU/LTSyOXf4/TJHkI5WF
BEMq4NYzrXJgkk1yU4DF2w==
`protect END_PROTECTED
