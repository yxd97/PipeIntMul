`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDpwfm6elvf/fbsWtrpm73nOfihCQj+/oJz9giNENLSR1/S1v5Lv6bDqjvnD4uIc
ALK8lDbEvcScBlWwlc7yeKuon4cxMoBrVZA951XcMceayGbALRjg6XKtN+b9ZS1L
AVIw5ZgeO9h8GhiZFEBFngFkqfnixdH1c7CKJK13IPrEyrRZ2F4NwWfVJ4ThJHC2
ge5Ao2pS2U4M+DnoQOnyOs+dXjD4canec0ArfNxND0T01WsP+2PunQCUylcQ0vFt
lm7Smr3LdF2aCNUjXnGeCQ==
`protect END_PROTECTED
