`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTuIYtJjRUkJODrwtynyMY8ooOo7vgkjspsGf8czHu6MPWR4TqQpax+htwdqY5O5
ac16o+8USfsEl2xAM4dYs0TiKToB0Rpo5jPqP8FmZa2X1kUkFjP8rY6uSgpwvVC5
xpmIiHpUW59Nrcp1c6t6KLZkwxNHHXzwmKX4GgXCZF3ADodczYHsaD1cS6FdirpY
JPO9x5cUZqyc0R6Ll1mE6UhxiG+V4t8Km+WCMv4OOY4ykWEyIsbe4AbLd/7NgY5n
m27ptgzVFNMaAexxcZD7ZeLfN38j5NTOUGkdMp0ljjM=
`protect END_PROTECTED
