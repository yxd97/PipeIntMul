`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
suMmVWstUUFlcMx0nDxhxEbFj+xKQl1WipdxB2P2pfE26YiU+DxjqzOg17w77zkH
+/ttrZ1hpCNa4knO2Yj5pXDDhiCTz0spXo7Fr+X5kNE0y5hPcaeq896zcneZYZBR
PP8ZG+iTH5NIIRXNTKQg2s+ugDIvKZ8dciprltobg2wHVi250on524fH65kiCML1
rhqVP7e/U2fyg9YZ115Yxa+AvuogTZz91MG9tRNdFG9NQ/63dRjbepfJsE3p8dcq
a0PQxurraD68GFchs/F9QKa0aG2uTMCpQiuuuAtbZVdSQp6xJOqXWlvg53tIFDzM
LQQbj2QxfBAZ8RPO9TTRgiqeFwdHAyyJ2ADGFtvMEY+gutvNfLOcTBzKm29lThAB
VK4km8h7iHkwXMx2y4hy6/Ned/kx/Y+jGy5OJQz0uhM1El3WXybTVTSS/aUKGhd0
a0hI+UK/97V10NdKJfj4PqfRuqn0w9JK4q/UiYKjdDdcS1so7cASQmJQ1LR1LABw
QVbx9D61Mlui9IOCHcxCGcJRwR3zrQ3d11iPzDiLip93GQG+XQh5nphm7aOc5IBH
rF3EEsyF2eVB3FRZ/EC+5RIvvRu49Hzg/51Kh3st9d0BTpaLmMKjA2CX61jl5T4U
aycRyBsd2IRd2hYdm5CkKyuSHFhcYauvsvhe9W3rNC+vBp/6DmIEMD0jUWGPKFlt
/VC1vQP7AoqyAoorvNDkqiNB5Kc6uuFAldMaT99sT7C+HwLQjam9eMhH/XqrZztt
HboFse3t43hWiEDvH0tsO2bo3p8YX/jPpeiRQfm2GnDZeq4YDOduOiZykfDIg0ZU
w7sV2vv9WoR1xB41FRx3poBBtO38wmF1VQe2vJjBzKkcvhLU/dUuVgd8JSE0YTxn
qB+Pezbo5yeaNS7RONGcTtNKQAukz7/PVmMp3smHpbu5cheSHFZZsX5NN9H43ZnU
SvPGty9gjqDh9CM42e4fZRZWsN2QmElr9PDepDlhYoRceC1WG7W+mF2um1xVElZh
HeqQn1a06DSQ3a/ALzoFhiZSrRtaNTuRSUsfK6nr+vNLxb9b+Pi/uFeE072lvgkE
/9e7p2gqQz+yXwVAlP+Qaxh957lBQi1ZC6XPr2CYIoF6Wbf8noRpJ67tPgb+97Zu
qVpRkkVgy4TlcFlmpT1zPpFoOfFbwFHDC529dMFsSs6uB5GYbHFbu5Y7b+olWuBS
TS3X6k452x/TnpR1+dNLKm+C2XuTw/+NvVlkTmknv43Wg3jqBXmKsKNczZ5yEWMZ
xTvGIW88znQFwwPy/o4cp2popAoC0Nc+VKfIZw4vR07VHoJSsWgeEif0lZLMdzDh
l5ya7JFc2R7pCwaZyxFRyTzUbDb5Q5DZBDpcNClPG5bsrB9VcmiO5An8oNRAqCDI
B/OV4UEw6xZlbdeJ0hYxrbo6NhiVKJT+stGfkA/0CcT9p5hq2kGalONLEzUvVTMh
UkxMJPE+40Wv7Wrl9iwJ7GaLYbwOEn3g0hl3rNELcrCRfjlJy1jEtnFNGhaTaFLI
pqP4J1M4WOrLj+IQ1jnkczZ+U+I2jJvdHOQbxw+WtJN/UN4ZhRNl01lE0KE3XgUJ
2CDHGV8+kjq5YJmTlygwWO2jrSAiswVlJooKob5kfHxPwEOevEU/hJ3MbyA/J7LD
Wxf0ZyzfDi/vCntnuYMrNaOuHtSuoK5JWCAue5IEp+o=
`protect END_PROTECTED
