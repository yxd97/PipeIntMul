`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NpSoSCc/M5bGNOTVGU8NsI/sbXjwtv//aVUGWtp4XE8O1Omk9cm4KD9Hf9rEzsq2
FPMxRUS5XeNypsJH/rZEtfh96DI4kyGMxxHiNJQ8rds554G5Y5Kf2fDoDkyHXYev
AsTFZ21orDijooqOTVFTotebGpMEi6XTuLYyQgADBjrLP0MOQx9tkXwI7v4xaQhc
HA2qf/aQCm0YE3HTJFPYFnqkEJuoVL1jfRFWtfPhhowW0KNUpuSlj9RstHCqHJxT
YOD/uuxW+L9RaTHK+IHkvPhbcDn0N6HOwGQi9QmxCXsag85kLiIQ9k1doKLJAjk5
W4XDFx66srZOyi5pyV6dmtnn+lVu5iC92BdLk9snUQKM8oUMw/r/HC0XTpN4xq3n
0U4PdkdPAbAsXVOYNS8Kq2o2s90tNpEWl2bHcmuU6GS6ZydQCSe/Jh6jhuZ7ronr
Ea7qxOZYNoSDE3UetkBiKUBkFRjsSLmf3cob3iE9LVyNb8VEPxTqMXLVeu47p/er
WC/2PwT5a8W7+fxN9Kyry+v3kI6iFcYvchQkygErKXWgXGbUQagsLgd+rcsBJGPU
IiCsbT1ZzTlYLj59WXeqzspzNJBNctjasuIICo3d2Vh0TyiJV+bKfzca2/41QDNI
WF3jSwpGP5rPkcVMiyGmyMVwlPi1ywwzTGXPqaWjzvRmLoTASbE9oV1L3jUygKG/
X5R2mg3DHcqapPPNPEf3H+Hge67mauwCt/yZhEjz2TZv0Ie9gUnxon8Wol3zqIjc
p139yd6V9CgD8EXc6SScopCPIXOzDVod9ok7NJlP7WuW54bzrGlzn0MWAjQrzCVo
/7dhullbvKxxpj3jnSxFYEBF6dLMjUs0WOasKfu2riHG+Dlsj58yOfwquxRNHeWb
3VhFdRBqNjzKvcGXX9lsebVFifd2ORcDWIyDCc/xw1+qontX2iRHMMoQf2Ul1D5Q
a83ldrPDqRuGVD6LziSYWPZX4Ehvqj0hwM8U1cpiQNEnC6YgCHD1LE02aQP9UJgy
Jm3XOkb04XOoaYw6PY11OeCpUutHCiKTXiHMykL3yjVk0aGC6Rj8a6zosLzkOnv9
V1uCnp2k+9P6qxTuJ/1/XKxmIf0zGmaK8CDJ78BL7gzQQreu+Jmq5BxvehiBGmKy
MegFg4H70eeF8p+CJV7527UMVOJqEevg0GFSpXXIy46EQWTfG7riUvbKHE9fetX/
rblq72ku1/BkzX1yC4aRSSanFiMnjaekEg+dh/KjDhpfGVPwfhMe2XE3ve1rZfLA
GzuTHyg3ky9f0DaqdI+C2bO/FQdYd6zzxPomyjt6QN24TqdWkF8YqnKiKAYGNQ6v
7pJ2pniGeoMbEbzvWVIx5Qcazee0amOgXeyKPPoCzdY5+1tkWT7wGf1RS0rzxUrb
3QcZ3tibZ1iwF/a1BLtNynNKdcanvCuwhoSyBQVYk5yMhING8MPweewJkeeEn6Oq
/nyQMWwk6o1AWbVeTiQxZiA1PDqs5q8DK7TOZXsLDG1uApmaTiz1R8OUJNCtp2sH
wY53OMNypGWmbN7sjfZrmm3wx8jBwiW3BfmtILfogUt5mt9WEu393VHCO2ZiXExB
7OBuurvmNo96ZpQTBnuj8B7y/P+Kh9Rr6FNUsGHc1Az+2WnFKyG6SfgGYM1IKU50
rfZTjO/mQ3TDLRYBYcjfYtdOgWu+10bLUsbRh199BtkeFsW2/FldEPr5ClVP46mW
C5AGfWztpDDnhVW2bhDb/g4tCHOs4WY039tItJN89ml04Jizy2YAKjT5761CeQML
mthPbyevxSEX4OirjnUCdUZPO7BgAuQAa9WQOIVDBzUaDbIoWOb3cxXgGnxFXHdo
aS6KCZcUZRQIWwc5k8f2YD88dIxueultj+ebCeZeTvKaJG+BqWe9zwTchfFdFG0a
r22rlqrDrH+8gjwvYkRmWSmNPJlqSYr93fa/5vDTjrdSlWpdtes1aCUJvW/4XKfP
7k2TMF1lL272DfswqAnjRshDNfqt0jbizCSINdkfA01JaMz2j7PUwIgXxJXPKCtK
S3PWL8f4vaDs1Gh8V21hiA==
`protect END_PROTECTED
