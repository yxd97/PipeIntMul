`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DSysUcRjrej9gVGgJP8uUGoiu5sI3Bj90rNl+Uujc10Iv2y/Wgc40HYi+Js1F1kV
ps8gQdDYUNGp8gwd4mQGFkvIfA+nuZkmb0jlr7szQyN9jvjvUn9R0oNkkLEz0OHA
dri7TFebZ7yakXqkVeLitjUMEUNNaqxOx4MI5BVYT9B9BzEqK4I4iiyrd64dVvfD
m6PIOP41h8KukNlIDYzQgqnGA8zwex/G/tSaAqDWshLqyeSVA+zr2/k+lTM1QmmW
1TI2zF0R9lRWcsf4Tr+gaIyuh0RBsuVywRajjyT55l19/C3r8zpi6eqo5gvDG5Hs
xeEhpCGaaZDSibbzRrg/Rw8/EDLN3IezJEfzYE4IGYwiP3xANIBgEcKt3ArtPPGd
9AuDkdiik7BqibLbClbCuEIZDRvvdl2ITojBOob2dEAevOo6WAFftnFWeZZ4aH+j
H+uck5u+BYVOu43iACYXVgU+UmoYG3a7yJ6F7wuVW+keRxHvmMKbY9HUHXoDR/kd
8mqwW8I2qUhNfYCT1/fN0F5q77jOr8FfC14op1eYz/uPvQSuxnN5sb9QyccOQ6GO
GTRqmwew1lUl//twdfPpEsqtmG0xdlW9V7NzZ1Xehl84ozGpYTnO3MGzwG6MnzLF
2W8/s9kgLaMVH10jaDWK+8buSKJEVo8GoR90vgn3xt1dDyjgL0tkKTbL//v0VkaR
AOcKIIhbN1oTIEf4T6ko7majRd1I37IKPyEpzw6vJ/Y2XJdvVF2Eom6FUm01tL+v
JjnVye7vjc3h75cPboAdEK5PnR9F/U6K4hxPP02wYRkF53xQoo+br46J+/9Ex1O3
Yut6Ly2hFD/hHEIctkATEV8OYigs7nSjik/rR75cHwivZ79kSVAKyJWEmaxWRZxo
WoMBTr3yrCWLiGeUS04zMutZlJJ3qZ9HyZ5vap/SlRNa8dv3M3HW2cj3f271wdmU
WDaI1IHlcK1s9KLPja4M2kRShlIT/it8BGhGtVf5mwkeHn6AkJw7OkjB0FlYi2ug
+VSgR7Cke7j7U6dpepnsCGX6EeVtD2LqV+PJiEnYbRtBhDil3HJlzaDCFQN+bI2s
v7kfmK4SHIiUUQ16bZLUqoH6DJYwOf9lJ/xJKTbt25P+sGrlW14O8yt4AjiEqeEN
+MHXSHHGdIxr6XDWBvwG4v92L/CTnNV5KLhTCHkTnI22JEDwFw1H/KCCWvApBn4n
nKXnt4ZJCSyNIs0pP1W00BfI3TOUH6r/3Vje6bCKG38C7wPSfx4PFbPb6EpZuMHV
mROopK4Jdzig8jRrmuqPErCFGPVP9QVpibJFK2AwqSw=
`protect END_PROTECTED
