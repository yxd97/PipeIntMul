`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5UvQjl5heWXiBLdZg7zINPnnNUGdc8D74jO1OJspi7e57N+2keyi4K3EsACCNA9
MJWyF+uPPFtRd1sZsOxqLMLjr8598vNJH/hUi1h75VJuWJle6S7DjCQgV/0lXf33
LawUCPf2Jxo8PFXyXgS6TkOLb+x8x7xrRwO8/b/3V01Nas8LpqGKbQp0WFRlJsaz
ugp0duGTrgVdZEunupzzKxHjWPjYipnnFEU7YnUBDPyk3++wwiK3S9x5YyUiKpRO
oF+d3irMwgN1Z5swHaV6a+kqAocX/BR0Zb7hpyk2PE+wHrCLc7a65LhopffqoqWz
KEf5tEo3738ifCEMLtkpUQ/RMgOSKxKfajvXie5y8GE9mv09+xKQu88bjEjR7aBl
gwPPIsBzxYhTyzYVSlT20w==
`protect END_PROTECTED
