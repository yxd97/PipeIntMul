`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWo3TqbL9+Um2JDotS5HrWktL9TqdNsaLygGjmGoFnBGC/FrKMXFmITXYrfdgBDT
gfsnA7uIQO0u15AYTRhfGGPir4iHNi4bGSULNhQNBPX3aS/aOZu+h6vjN/7ZvJcA
5dw1KBPY2eli4WWvuNPrZjtKQSm0eVabqvo/JDbm0H8up9enzRweph/CONp/LqhM
BaZy8fbDwROltYqy1bUWE++gW7DiDdGptVK2wuXH0oKPR7qheetaAmxUZAH1DTMD
pchW4WKYKQpzVsSwLZBw4LBMi0yC88xhR30hE6N51h7yWGLtxaklufqmHZnROR6C
qyM7Eo5S3re8jdBIGGf9jpMmU30ig02JNVL7lXPOnrRL5LxnSqVJGMdcOFtuHp7o
fs0KpLpJyeoZEa9xmi6Sd4rjVG/k4agvljTwZ80jwsMIy0hfLWnSKEshVO0/4rF1
2o+hy3f3mMDCr+l3JLYfPgvD30wTC8YnUPPQrGB8KiLvMIxprnZ4gtbEfs7BMtgA
+b9TkI99ZsnlXjcPR4slR9DsTgiPsst0vRr+ofAtcA5sVXep9QebiMBOzuPo3q38
/c9LROnwVvWUV+L+EpiU/xJfk+hP9rkmgHd9WXk+hta4xm/TQ4GgqFxu18yzxUe6
qbpgV6u09kekjGs3decfebpd+iFQ4/kLT7hRrMnFzQl77kq0Vz/LqMLcRlScbHQi
wSsiMQeLn6dcrknF8trbjiKDKu5v2R/3nwe3KjSbmDCKsGYWEA4F8a6NhQ5zEk1m
lex6uVmUAFk5UY9GO6n53fX+TcH1oyZ8pO9SiTFLEkQKwg5v09yJSDkKBMYiyFNG
jdGOKDCKO8v2ncf2H3XW5sXceRxPiRIvMmxSZEh5AGHcjfVfMeKX9AMtFbW+xZve
+nHUYYRmpr0xQ5VUyzUX40fDsRWLnEiCiXLgtBntIDTVhfg+q03CLLQI4+GODL5a
hYVlNoICU8SHkG5qt3RpHI71E4GmD9ChT5iYXlvEbfrPppvni6rYEQHUNaGzK1GD
XsbBH2rrsYEu84mu3yxOKDH0gOGzIwfodRgsP7ahcnVaOqFyw4gGpuP8TDG2i4Kl
hd8na5Yv39KkIGAjPgoi5vGkGAIuVDGfg0tWqdZ5qAjG0KEwM+gcgGvxIxrYLwYe
xeW7j4wiadgBLdXfVs5MhXVnNpHeslRzZcR7is8o3jgtqOy9lf8mQNJyPz+gyTx/
WlC9JtkyqR0cXlde4hJzXax+R3+dBu9TMpVGQZqIfhmNerymO4UVrFGhylnnlbEd
oPl2yC5xYyG3S8d04p4wnEIs5/9WqQHDPfd/gCGqYGT2M+YoKpigfTFpCliY9dZN
f/aCDiD0KuY9Wlm6o2debE5p8ppwFM1S+cQDdFGNYFHbpGslRfk89ypyFEO80WXL
qHYJAal/P5vCkYO8IyC1t/zIDcTR9XOI/gK9Zk1wEZLWRgCT8LJfQA4Ux2tg/lrR
3MVdYrM6ONaxtFxaZCtnMZav/AfKPPVx7bLbxkJul9u+3AVOIewoPTESNP1zHS9C
qj4vQksKy2qRJ5BVum6EWw+Q6vzd/9kWFObtexHSotIZOzOHqDcQ39yeHXwMKT0e
U8aZpJ6DpVdFp+VHq6Jl8tIeHYHgwnQHNNrC49vr7CAEc6cVlyB9EePrHmSZSUYH
MqrVo2G+R5xqgIDAaaCw06peU4jsWMesp8Rt7xKKDO1iALuFiXa9qJmk6SGH+DWR
+0H/JxKFi9Sx+9mWwa+U0OoAmncLlhINhZ4XQE2I1C1e/GHM/uIBvINCHnC0M+CL
713LCSnr63+UWlW4cSblYpAGBBWFP+p9UeEPh6pAhr5AHxslkiqxkqigPVmxSSBF
yVIpgWafuJ+TuVN/kiSbT61H8iYaLo+BBRPjo0w1kikGcgJezcb+C/qAq0KWsFkY
hONbkDtYRoVb2d5dhigEGFFtjOOekzn9W5agatVbs2g4j2+Xgkw6+42rCyJKWaoc
yjTgBJwvzCa0fe1OB1/3KIyXuiHnnoJSvpLwVRiDoDbCpQciLLdWHGHa9xhmiM6y
AooMZK7CQGu/8BnZYiyfWDbuDi9P4w+kU2zPHrofOdg=
`protect END_PROTECTED
