`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ep+qudANH2k81P3CzYnaLMUau5fPDvlO4ZyEBM69jfiCrID0NqXSX5WOKkkUF5U
w5ehMJVYkCkgd4NZSUTOH9+rRwhKOcH7lmdywnM2OzKW2vjEeqxeKmyWgfK6W13o
qI3c0ux1z5/D3YDc9f9aPDQgzoZgP8X43h3t1juQVfzglPiFxWbFya6mp3Sdvds+
dIfiHZ7lGEup6PiUc9Bg5tuystJyicOm+7zufC+3PMUgbjUTarzZw9BoJ/gOISaQ
cwPOwjauxVuphLfkwajUzHWY/5yes0ZhmdOe/upe2y2UzqUHVOqsfcd+HP7y9Lgd
jkj52Ud0eoqzMfSmHQAU2k3T7CsmZj3pHIuKoNLIwvVt4Q564wjUjPzQ/DrxpEL0
gpuwNWTP4gfZChYxVKL8jBowH3QUrFO3xK9IRyo4rAFhMO5fF2eZq+1C1Tlh2Dkr
Z1MJ42eAFLNeMC+KXIm5GtIjAZ10aCD5Khslgpu7yChGofW3vzEkEFcfO7y/SviC
w7Hd1ct0bDKGcQtcGnTi9nKC5ENVoOYWnD1JyjnVZqxHbzCp0XSe+HVyneK1mv5z
AMBw8qe8+kUjgdsJ7ZIAvw==
`protect END_PROTECTED
