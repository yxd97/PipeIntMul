`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WzSD3qTxhSvarQAA2gHSRAcsiC/eJxaUH9eMrYERppbRu7S2fbINluegrPgDHPIj
9meEXo++FwEF0w13K3VBFjep/mFh3DwEcJEQzRvs3EmtvqIC0K5tYFNC7bhANHfb
ByHgAJI2mDvM+d5HF+uVZvs6L/ILPX+s49cwtvQsTdEdehVJFLSSi1/9Uf3KXYEA
CakPGLVKt5Ye1BzVM3Y3/S+Z61w1HW5AmvPmko3e0upXSZ+ZVnXgiBpK7SLFXDVT
GnlPpEyRNw92NbVmkZwd8QzzW5mWDkwCcHKEwhCLrO42/wHNye3XYYZTUr4Pe5AO
AfbvSrNIC1wqPZ4v2QzbSHUO6l/mUa/KvWxsum4XfWZqPVQ3/QYX5hw9+6JiaiO1
bQ9pHpFRJK799tZh6USdDA==
`protect END_PROTECTED
