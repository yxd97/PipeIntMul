`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4mz1upozySjuXb+8oyRos4IcFJwyTTgi6V+NzwcR0mrx4GT20vALgTMwZGwcCBbw
EZ8hsM6mFfDdIEDZ/Nm7SLsXr0ipv6hUiTzSzm9AQxH406XPMVHpZ7gMixfdY0oM
VvKrscUIHOj701uJQZWx3ZQaYq7JCVlXxDQI66VOm6dAe/S5rHgCdOXrJwCxVukB
+Yh7h6nd192pOFOgXdQSjb+MdccUxy3MpGQ9KYtcypyeePTJe/W4mCCyS1TzaNQg
jGys9qkOqQG1RPZdIZ0/Dw==
`protect END_PROTECTED
