`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PWqE7euzn0l7dfm/1BenaozXmn0eJKIGxNewqf3Yq9AcTNByeIgkO2OaZvMbTEv
PnUwetADiFbP24ILyK7IJ8q1M5fKppJ1V8k8DNbQp9LhoXAej6dmdVEJDvwjFxYv
iKmZXlPziSI0NJgDmfj26MJvM0fGu93ZojjOrP7udCqkbUpXPXGDmrYQtQ0bOj6+
lF9qpp1SxFrYEKZ6Ub2QyKTWr25R9474IFZNA/utw8sQ/NNQnQ+NuZwtCgJtlx7w
xvl93wBQdQT4UYIPGNfLraOuYd3MMJDmyZnWBGntRu1XvbePCN64uSTiXYN/1Gu9
akd1+ZKkQjXYxRRoCL6s36+AHUC8ywekcXDsJSvv07ejwgbR6MKEpMIHJciDMw2x
mYxXP7l7EO7wU9XVJKbXYeeLFjqIYp9vCEdRNFK2DPtLJ292Py2j/grPSlXjzr1i
7fSEl5qqYRbkz17E18gw6NAQcCeo08KS3kXG22uDXJGdCsN2ZIygsg1/nJYlLhJk
uCyptt2MScbrsCDlFsyCsuzW0o/GhW1/PVTbr9b+Mww8hIyaHWW2rjC6csZ2d1Rd
17nGvZDFHnmzFk0d+Dd9yZMh7ja3sMe5zCF0BAclnIwpmAhBPy0CQUriJYu7zmTh
1zi9xQwKSbBo2lPHSFLPkBWpCsilpK8DXd+BzLlYlcAeEXWocq+LgGkrwteBpzcf
H/Ww9MOKsgDn+ktwvIoRbW3dxhfBbYfXgtYKJM1LlWIRIUqH+OHBHk3WAIH468vI
9k3GUyDZy8z+yUmqaB1wgg==
`protect END_PROTECTED
