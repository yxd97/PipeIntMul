`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wRja4yMO4FQ4J8yvBl6aeekEY/o9j0ZDO6OEBPsAJdB6mYfneKBqAPX4ZYdgtT7o
xlyFpzc5b7By5khCqZdD6Ngmj/7HalfuHxwr6co6bEBlyFzF8RzEflX7W0ayIQAd
NRGN6lnS2X1INN3KITmkQbCbDXWL2mkU1D254549g8soPyJ6OmNYtGbyx6O819md
SMzgTkFQVHovlalkPoPssYr4w6DjTurwAoMM5ixmrjaQPlej2M5dZU1md8Fzb7G+
ZHZYVVpXpZyzDzygcLtkCg==
`protect END_PROTECTED
