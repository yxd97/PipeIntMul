`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcHQ0dmVu/OFybjwPM2h5ZJTLpHvJuHaPnjfAMZ4cxMK8MNdBm+8+48VPvFi2crN
11hAOuNsS/nEPUdHsacTEsjGGyh0m+2vsqtpp570Cv44n5T17BIaIS84vYjd4sk3
5kYbZOGhzKJ2OpPPgtR/Uu0lDIU9evChbI6WNHdmnrKp1LDIxJcDHEsLap81N/Wb
go6lpdINnrCgTx8F1P6ukGXb7AQGFwxEZnH57tnBxudsYZZrH27nrNX18pZEtTD5
a/pZ6NcnhMpMjHQRfwMa/v/OwM5XhMhMWo0V7sAOv+YFD5WHR4t9qCzZaOI3yMhS
9EWsfEv5pTHJiukQOxEX2K+Ui8wSzhsPOvxTRgVENy2XKGEjZFhPxjgKfJgWp5f5
kwqlIy4KT0FSf1XDDkLqFLP8wXL6Sl6aJWTalnI+doLW+oBfU28GE2iyDTw2l8d6
uDTAO5oPqMYoyTud+xIM9Ld1J/iuG/Tfl3keHYmUA8N8/0Yz/0qcMoW2P684XGlP
UkFA4K4zzU1i+QRlvfYtpS4ebBgAmecDLlmm1tZ/5Gd+Mt1Rmkz1TiD34lbdtest
cfbueEzdJjS6Ra0o4+xh8RO/uave1Dq4r/BvsiLCHlkiNOgybzi+D18oGZj8lX9g
pv66z9dwrMQRx6AI+fCbICXMEtZWlhp99Cwqn7qeICg4JCMBCcysnFQWJFANTdwv
wGlayLRdm7zMnVMs6SR9jEOtyVBTtuC+M09gNVoqVSs=
`protect END_PROTECTED
