`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kfu3oC6W+gOlkHzHCXsEhlQQWKTCbbqcOXGg1xcMfxhoLhDrVSDxvzxG8NxSqnxs
k7vgC+iNlggnGcqA1jzkx7tYPXowe6nuRbrm/6RAVabYuLDPObJSDXTmTdb1OO3t
MrVW4khsa5/Ap7Xqy3fVXJTqszzP12iDXpo8jhNjCVZ7uwRQAv9hwuHXstQaj8bh
TsvomAoswdtmgPO6pzpcKD6rZarqklehlzQd77QGVLBj60Zt+wdW+943ljFwZ+v2
NMF+Op49zUJb+EEurKKUPwegFCprDS7mvqbbgwIwFHEgUUA/9dfRZVU+DbsGeGzE
9H92HqgIp89MzQt2s0cRISaejkSU9Nx49+X9YhSDVR2DWHhJOeY4DHs3ZvGcRSYj
yRJxQXF3sjr0YPWSW2cn9/ZRGSx4sld3LCxA3Pk7XEnWAWmqqkJknNdPd7FbC6og
0k8qT6QSXjQyrsN57IjDEIVqEEwN1xrkpaSjgUJNnNMzrirTHGNt1v90995Fd2Ll
BDKNPgX3XmtXYf92GDSXtMQ8JLWwaj2dcvYI4GSO8VJ51M3oetN1oAlJwp1I5WHs
pGnRhPB8bTeJH/aKqURpZ3L8hJAcsdgx7IeteJ2Z8+u02JsEbC0yUR6WYFaanid4
WDMLZhmAoxiX3v4nL387q9hpAKsn73dl6bVUMFc7gmslvQGfHSBIbmhHamNPRQce
qkfzb+afyBjeJhykT9O06GgATBOeSXJmiBWUNEXlZVV98FNJBwksvoe8Ppb/cUeR
3erBU89HDUxp5MRA30Q/WVgv4wXbU8yhUS10Tiih0m4=
`protect END_PROTECTED
