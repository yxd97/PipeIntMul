`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sLVCat3xgMH5uTwrK9+4QXA9+1jfjOFgE15gE6ZjiBLNxmzOjiQZUeP3PCXdk7GG
kApvJjyboJZwu9jXamYoKVQUeA5hVxM712BCUrmNIxATgMmPAjNDmgN/bh/lsDYc
ptK7sDVCBuj9xsNJRkjVV/RTnW8jYLTid7nhMYSJztXBsoy+N2soUEjtNAUlwaxu
jaFkcvIF+StGQTXF9JVCP+y+6WbbUQjAfBr2vASdhqYeAghL7Wdaj5x7lKE6OEVd
Wzaj67cn6FSIXAlUX/Xmu5GY009NXbt29eIbCORUpttIpAs3cmqARB3znqgPMqm2
3fQvehPjMZ9KIpdJQ4VJ17iTgTV5Rrbb3nF8rNAek68=
`protect END_PROTECTED
