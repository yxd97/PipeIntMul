`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q5voY2o15Ujgg3RMJvGOwKjBs88FN+kVSvHUN+5NpDmAmVRMDTBSKhHIyfePQwVR
3gXUGmx6f53wyPTEdXgpdhE+DC6dq7ESCN2Hw1ya+9IxgOMaWw7XsON2J2ld/45O
cWFfYspmkaq0AO4IRFLv9z8HGS1GEkmhzHsqHHQ5BZEDb4uResg4xZsVJFrPOEyZ
DhLpEx6zBYwcHf2kNsQBLixylA6NgmNRlDDLfKHJFjfkO378cYZa8DYo6S+vFJrf
F7CiWD+Nfs1jGnyW0Oi4sOGTMzty8UTpDK1asPnCcBgqn/+uI55FNqD0nzNJ5KBL
l33HfK8Q8fis15CXrXsXUgjYx273BNZVEYszctK/hUpllq9xVMjEYQ/F5C+RIVqW
ZEaz1D0qAGXX45wRvW+2IzxUDMXC8NytXMHfcBcTK3jFOTxexliMpS4bcpOHM4Ig
5Leic2CadfemH0KrWmxHHtI8ffN+e1f/S1Ramns0IjEPJ2DptWt8CaQFhcLzeQH3
dcOeTO2phmNEsax2sIOeKF37xMhDKUjy2lQ3inxRRdMGCDjgZm/HUSOzEDieeCzs
fGMDcWNeEDX5Sxnzjo+JkDfhdNThBa5Ug2kDduakLM5IWnFWxYYVcMI9tPo2DJvI
Xepue4yOcy9S8L9rYRa74yUbDg58tIpcJf014GgBRTstBfC5B2LXsJrBhmTmd5NK
SReI+9YeVPBxRFZLJs5/wDE3GGeOg9e9L2B+lHe9T/vtBaz/OoizG7z1uBq5WQaU
Hj6AwFwF8mD2OmTaSxlUAWWPId7XSk8NxZipvfuat+AXP9HYEWdRmiJPEnS9lL8P
r1J/+4qvN7RwibHOet4a+Mtb5xF8YtcF4VXHqqFah1Gh44/QiI1Ezr39uaNoXxOG
zPkQlHoYQsnm4B4i83yBt/NkGoCPVlshNfVvhLQC96urdZF82SMdclAjBnLH1v1N
6fbGEoG6cBzsS3k23i5PLVKfMOL8n8WFFMq+KyXgLpcRwBTSwgZNWNzNe2HRCzY3
DKKvdysuwCLJiBpU6d6vpd71kHjwaYX9B2jkDRfho65Icg16RkyESIdJU0mwKKD+
QShgAJ2zmkzJEJo9HBO5PUMzdoDXudYI/Yc5PgB7tg0CLy2b4AtVAdak2IIyEBPW
40uIlkAwwm07r9QIgiSIOS+bt/rIYDbDh48RgPQRebO+Ow6/dGUZ+5zSQNHE2Tgi
j6SkUhWQrmX5vjlCyAW3xrSnFi89V5W00nZxEd5S7d2uVWm5z/IdtV4n0LbhWd0g
aAxFvKMWv44Hux1IEGcg2SoIqGUjuuZh3lBSLbRGmmTkTc4nT+g4Cq9kHBJ14wbd
gPg9NpIFT8yUwAvwtFGoLbLezaXpO+n/6B8Jr+0b8M6jbVvY37kb3ki5jYjDiomY
IpOSykb8WbEwTvgpXiDKfzsvsSDf+j1hIWTv42El5SgYCBCCkpBaQ4X+qTv7ZKTl
C+rJmoxQ+ZnC/NnFOblunfxI9XDANRBwzGQYg1Jf8uba8oLtdRHBpR53rGrFa7J7
`protect END_PROTECTED
