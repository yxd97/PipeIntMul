`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIhqpsd4aZZMjvyfFakbUKSCpvGCd5cAeeAdoRj09qjbx9USLaP5rW8cOc3D8L+/
j1ps6lPDth1aED3kK5ccUbUwWXFxDMZByAm0D2phpQwhrV+KU9BvsHOabKVXILEn
tZ7SbMxB+Emy9DiFJZ9xmoy6ukb06sgTuvAkUQ40HLlRlkNxJeSZKXTOzs1j2LB9
IiR4RMadeZS29poh/pcLRx1181OeppT16SGhDJExKCVedzPYCyOXulm2Y9WKsvkC
OUDiNVyHcx9GYiO3JEPtvCqWKw5NPuXMIWav7cz7Ub14KOMiClxavnotlTzPlxhu
g1FaBkyMe/qiNWokz9GDKUkvFa7HZbWB8t3b/9Ueq+SGh/ho6b0qQygIHs1hB90a
qqLLitqWgulxaA6VdUN49A==
`protect END_PROTECTED
