`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gbbb8WNLiqVBsPXZ+m1HtVVQLPT1I7A5N5GHmrS5/DlpFm9XGoeAgpNSr7X4p36t
M9L19SjoQrT0ikj7DzYh2LFcBTcM7gLe3R58cojIv0ZWLkEEr7hVJRUT6aFcnruS
aJfDpHVuXpCFFgtd8NTI11rtdc+roGx/Wq3DBWHblwp4hogDy6FNTDfMbCJHsdGB
kxDYzso0ArnuQrZl7OFVrp56etBWvq+IVF+ov688s8FTB3L7TfNn8vwYSZO8btum
`protect END_PROTECTED
