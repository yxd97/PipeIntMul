`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3dPgYj7mXWe3iIKbbWSMWoHiICGlEJxPhen3eFdIZX8Puit74yzotcwkivzfIid
3FulTnef8P7dDw2IQIz2w/4GHYbQtFIMLZvgX7T+fKEpLQhL8e0MiLha7DCuabEN
v2WAZhnhZIYw3gSiIWIm5EYNUO2Z5fhAApDRCRWn16YGURY4OLl2fGAW3fKBE2wj
cNOGt1dKg53NKxuqcoDsWcCWT6cmR19OREbNk5LmSgtkz5KiPcgxrQ4kQDd7k7hX
raIZ0q/Cv9/8MiL/8JRvMqTUXesYlLQ/M9NrowJr21joSI7dyJuXmoUrphiCiCvI
sJngVNiI1u6IMR2uR0+dPWRc14jsVg8HN+34YMTz+PbtIOJ2CcI3bpxBzRw9kWh4
47yE+271N8pVre+Kykhv+Us+l6A3e0bmU5hmws8hv5L9fHTXzse6XI969SzQ9zO9
3/oBMDX2mDExm6Y8NMuEIbwGcjhy36tIq2OGDrVptc0EEhlbSdYOWLjwx2NsU9wE
Ehg1jmZ0l9afaKa5S+sZcEvpRnabEfRNFTgg0HHHqoiphcdETz824lpOLxR3Btge
b87UxwCX/OUXteZwFYtem7MpTFliwcPNEcZPRBt1kr8=
`protect END_PROTECTED
