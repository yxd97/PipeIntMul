`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I0tgHPXFJ7CREWButC+4cVTwuKAqlGLM9PLb8w6TKF8to96OejUrklDJToS0huwd
wr6u7PeXrRenzpXUR9If5m+h9RrUNEm+/tNmlH5LTX1IHn+vF7Ysdf4YULqOB8sw
DSXvC3k0aQB8fWaUGesQSS43/vvCLcjO87WojW28gZKSADoZsayK3OfyepgvGos/
isk7SjOK7uteArd6YegWHAjs6wU0p98iv2YMszR4nIpuCxsCLOjPxkTx8zRPm8RD
8eqzRTObKKpQmnnjzilloCnM2Hwp5DtmCy0XYIAaZJ56Xqh437yHbxB0LiJjO1LF
19RnxzhX3+acNXba3wFmFg==
`protect END_PROTECTED
