`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4G9xbS//s6iV4cjnM3S77XFj5CESja4qWkHwkZtqaumfWPXpII6ND0rsdyjrLUgM
x96J1PELy+B9+OpNuXBluja/7NINLhpIvUZlmzXrikgWwOo/2m8k+Yyjw3aGs5yi
ZWg9gl9xpZDyaN4dgOA0pCKAh7pqYR37ywlQueAlnz8TFPaYlN0FkskKvgdXD8ZZ
gGl4mc9T23pttFKBPgmiPiLMERmW5+L9W0572ZLXxUIrIuzvr8sf9zuIUjgLvGuO
OvRpAMqG5lj9M2WvD3wK/ngdL1WvmUlJvXoTSv0GInjlifqS6d2QeZ/JsxHzFZd1
fsmvDUW3Fe581DxzLPgN0RxWdCmGgmlyKx3OgHHepfPMDExnRSjJg121s0SzHpTC
RKqyaruHjbfBXr3/XiW6OiA3ubqzFFhYe7oBoieGffhbNTk2yG1zCph6kXyAFtyT
d697FksyhZ0H8nSbGrg7a5DyJhaQU5i6zUCc3sgyow8=
`protect END_PROTECTED
