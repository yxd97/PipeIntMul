`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dBz4NBzWZD4VyN49FOtU+4NfTdrSoynBuZrfcchEc3RJcth1vm5tBAfjhr6OslBq
KNfOfYKJM3Dwvd8XCshnQtAGwEOpa9AkdBWHxlvnWCCYueZJcfoM0Ow9/LO9a6Vc
91O3gsTLcvuQKAwHDdPY5kghHN+G0Vn9TflcmpVNt5Kc/jBSOf+s8VY3bee+CLfc
A9FmF0InFNSUFl2isHhtktD9R3QSlAaoJmBTWDSdLC+juypf2e5ExVOPv9u1h4Lp
hIOExBjEkTh/M2NdbaQjcNkQGtIvezAfrjejF5Dd+bUaBgei1+5/n0PEKRx3pvTS
bz69FNya7PL+wRX7CqDixTakJJ4rW0OQJwcP1u5Pep7rc+aJ59j273znTo9PpSDV
C8NJxu30ncmMpPcd6ATFg3sY989cWqbCjKkXDDsga8fiIAfi1K8Zx5rvFwSJhlz+
DeMxk3ceGqpflbaFHGdNVmlVn6oS35qSmYyCyAWULLLGCZ9ThmxZ3UuwjTbKLXkP
`protect END_PROTECTED
