`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OB3/8DciIYicl+x07GfMN5r+ixqNP805d3MX8bQxLWNMdPdPid5yCVQtY3J81gcX
idzgLwYeRYsHPR7KcVLbruUcoF33Zy9KfrqsRAH6qSs5V4Vvb29UyFFV4sDjmFzt
dDOaMIbzbS0Zft33jMaBmldY1juyyV2icMBGfYffpb+IYPRIgjInXaIoc/rKLsEF
EwNxsnhIexxJEWg30cEQEq729bnML9CLzY4qXgMBZV4jEZGSzake1StZ/B0EFqXj
XWKM8tLaeXGpv+gkwuxii5PMZth7jKij8T647ojR3ogR++x21BU/NkIVk3P/neYu
NrTRifv6kAcO6GjMDxFCIvVID4KnTziXNnvO3GXJggLxNNdDeGz5itfkeUFT7aP7
bzs4oQB/n2QdUFuzH0+jxEna7yaCaAD0mMErSj/oDpk52tGKR+hMahqEwir4FFYu
MpmFCvnGiQqoCgX3EexdrIcjs+8G93xM+id25XZ/AjVigTi9/VjRyIDdFC3KuqHa
z2VAHkwP3PEPSgIh8VuHA44ixT4VC3CN4fqjJyrxKrRBBsBveMeXIC54uQ6+pQ/r
2qZtgv7AmMX80cdvq8gwJA==
`protect END_PROTECTED
