`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wi4Kc0I4J1EH6yHotYbY9uTT5ih1bCevCbSG+04626JO73nkDU6xZ1b56lWOXEqi
OTeslFrzGLQ8tSAO9yS2w7xu/OSeuUI+A3urQfYwe8NMwfd1T4Q6QaeKk36jwj7G
y0wtAAbqRBvxlI43p+E5OhKNGkIJ2h6x2PWpZDQxQ1JJRA9sQnwCB81erL+jsb06
AYFTeKMQSBlwdcI0RhXsuk7bm1+lditfsTNnumWX5ebnb+OSDeowy3D6/vKc9pZ6
4UGe9vjUqpTtbdIGErXXC9q2AnTswOoEpL9LQ/Q+9+TDO/LeuwpRLDotuLlVGqPm
byGu1aHDnVpqwXsw/PfgEL1Sk7k6zMamB3O4Yf5JWjjOUjXaPrCrMS8CbuAFfnRA
C2PvRWZX+0qR4JW9zuEyYpRbn1UdvZeozieFaxrRGLnD0DoANf7cY2ksn27xgHd6
kDhdoRf6S9oadSKPpAvKpgh9a5WXXavGjrrPKWRj19960twiBLTiePVv0dPmfBNo
`protect END_PROTECTED
