`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCnyQFyFxEkjk7N68pBAAkP4al6XqVkYcT+s68LDlMRVUoWUhl7bfaROpV311bb/
gsjT9tnzYHZn7rW8ECsZMu86fsUlT4KbrG4sDE6TvUmhh4oFbtkn6ny5mj/7JshK
5FBX1c+5UtJikjG3NJCB20PWQ02LZ+n+XTxuSpgf7QSeeLX0aaVV1iElOpbQtCbh
QMOvxiCWz6yB2nY5EcEu7Bd2rWbpwfzviQlDrzAKmCBxfMk1tN6Ch5hJouZO9zgQ
ncZ8KCythuH7htP5fZDuQQEio+XEHnv1P9PVfRHcvhoAxS2FwK1jPTKho59D6DYh
HUghzXgrR5AQciLdVxMXEScocjJQy1hJLI7Wv89dX9svdMuOM3/w0YAnvvxvArKg
7zyqH+rTPiXDBkETl28fWsf/E7tWWRzN+61BX+HVnOmyAFl57y78qJi9ZV6NmM6Q
guqDWPCkFYFAhMOQkryyoZHI9Vyo3CXcjFBVL2s2ScQBbKL/f1B/ociw/l/6n8Wo
IOtGlnwMQkb0IyxJ+avEmDJiprtMzdieVHtEaHYa9MlDct1gD5/dHqRNTUhz1Xis
z3sTN2c40BolA7C4jA97YOqzE0kGIHQEqzmxuwaSKRa207yIBjCtEiPjGCxqbngq
KhitLDtBlrLsmn70KSbvV02ovjNP7McLnuNPwhRmewfcVWzkwqu2hUdqqzFzszIU
n7dpAlqJLDb2pijkVOR8b8o8M3sGPcA1TSat8g9qz05Ccexcknwy0irwRkLUDwzU
+AGYbik/g90QCYiuyUuvvxr/p3BcqYYGDuu8amPRLukk883OrCzLb5drZMvvoXrc
7g4naweGqa0L8F+s3WNSmvw8lJ6c6e49Q/r8+61EoyQ8pYlc1e7RzjgPHGel5f4U
H7G6rf/zcx/R7UrcYzR8rqURgSsUMm+BQvqa4vBIjOyh7ATJy45uT6hmGQCPX534
`protect END_PROTECTED
