`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzIy0wSIU9vSNbdDBRlnYcJ0Vr5QHhInSHHCdVocvnB6Wn0bm7R7kyCF7hXC5o8G
K/neA2Ti39ZV4AaQnGni7wNdOwtRvlMhYeDXqTkwxih98EeFFSES8lDX0kpkE9lI
KiJqanMdvnhDDWsjrTmA1NTKU6GbKtJvRGv8Y8R1qiM9/YB+W7rLnUqIi6wwfY2A
uenRJU4mKa6ZNvD8oDXus9XF58gFGNWa81FmAdq+Gsx6QKhcgDDRd+1MxHsSSms7
m4ztFwhkqbUD87NtBW4GKMdIiUnwadiI6frz0i04gtfDwUCbtu+gGiUQA+b7U4r9
hSaz/WL8pLGh5Hh8AYgaf3GJQ4tm+fgo+xlVYSOcmu5x7ddQxWDJXehFP/zLJ3yP
IHDwaqRDbrvVAHfT1CxOa0nGJH09pFSWUN+0fvLc88QlY8VSZ3ccTSOFvgck73IS
Wau6Dqbxt2xNu8AKYJwual4nYIZcdxjwXTpNOReB1GM9qX+nR4lyIQQbBHrvWitj
M+pUK1cn9du8CI72CjKbxW5r+otOs4AgSu47mCU8D3HuVyUsoUyTfHj6/Ik9oCoL
mWVzfNM8UkO5uOJZhoA7yuW1SpZ/eSuihhBGRpk1GUFU3dg1Nx1AAaI2mR9TkcQK
ROdjMcZ9DOCw2YQJq0krdQhzyme4rEkz+yK/3RlDMsbFGtKjRF4HZLzUNrnK+aGI
DUwacaMd9fNxcKZ5S0JM2qrhVMI3s4+U1ivQ7aA6cqL6QMsbqEwwFzoaFx3DK/4z
XtAm3DRQnhI8o9z14GwLpJqTLAGVdaNPyi9iPx+H4RyNaA/GBTu4Z1gphnb/WCVg
8yIM97VD3o1pJfXm7ny4kTb+8TS1jYiZ/KH1DVn2nloSQFMp7DP6v5bCUPACC2oo
koXceqF2NMbc7BMBHopWZLOAqlrLe2p1HYEIDTw69uoBA8Oygy2KgZXQiM+v/I6I
EZvMWsQVUWxjhMeacfyY7rCxjNAZOYRSwWMq7Y58JYabvYPE5yRv68uO2sDaFOFx
wjUnetUfn6lAOrvcknVbzMzZL65qLRndv23KFMfRajM9mAjHRnLQnyjtYLpBfuWW
z0e+IAiIWBSJX985CDzstO5hVKfPaM1ntQfvx9qPEnc3zZH3/5BqMn1Yd6PDqDWR
D9S+JSqW6ctDV0Rui4PeeTyhImPWpYYtRwbanpYyyRufQua8UwtOg2cIeW7bPUO8
A/BegDApH8bXSX/V10xu+rbyvUs7fgCN1luMOOXcEoXhs28OUqkcFTjG/VAhPFIY
pyb2x8UUp5oNHuPu9DoADopcLJAub2lzym7ZrIQq3IZAHeRbY/zQckiZpj27OBV0
RDVbjn9kg1cGJwjTlSEYRXISKETfvb9eWY2T4goQYju5wN045lue/TayuXe0MM/7
sQFyBJT2V4+BYDoISyCh4HLeJ+pX43f5aJnOLeatQqs1ZH8C8T49/hZXEaJBULKO
jK5+V4FdgeD33+pVhqywD54MU8wIZYEuvnuVzWN/CQ/g0QHh0CYLiEJHDLq6AKWC
SMsvHdLQJVxFgIPXUp+Amdab3ozHhFg8fXGSgznzE45ULzw6A3/OnkV4wdGcDWa5
36Y6EgcmbNELpoWnjc1QuD4lLPEby4tK0TfwLCd/TmxYAYbhLzF6Afks+kiDIYvk
jmFirMR/4qwvamd4rbLFqd+s3DEnmowZw/2HByqr+tY9BUMG9TSA1MeyHrC6uxjr
Db+JGjA55L6DHdATQI/58dmQcChUDb22av9hDytQla+J3o93barb26bs5uuVhzce
KAF/nebTIdHthivzKqWIv4PyJ6WHbgQcqZz+7Erute587z8+T6pfyfHq78ibBbCI
ehBF1fxCbdsZF7lcHOkp1mgB89+9a3KAHQbbdXtmpnswOAwfylrYBtk3lZfNbV1u
47qD2yX5vItz40l0VKhPYWgk069zGs6OPxeVWn5nVJZTmdtRWKX9ppIFfzitMkjV
IUGCjmd+7hDn3ARnrL9pCGBVgcicLMm7h5NnYfPee1MY2uGauek/185EOJ4iA3g8
yUMioqbNxHG5i0X1kBZQACo9UxQnu9o93bOlwTIbRw1P5YQIL38YXbw+Kh2jcrIT
YXqzvYYARKhJ2SZstChq++j8ExRicSs+8VbSZFPKo7Owfl2LgHRKw2+rr6CAAxLA
AzeoqljzlRNuJ/gfYUaz8u+OSm7LWecTfBf85NC7q7Kj7dVHcZfpW8I9KM0m4RmO
DcQQ+FlC6ciJdp8cxohhE3rU+ZCAR2uTLvBmp4WzIdrr9PF3rICrYlGp0/5FyLgr
hHutwEMQSXNXjaNcgLMLML+Pd8Fc1O//+pjt0JrFdurpQAiy2T0TfpaJvc9MbKSA
/n2GqkLT5t+IR1JFpZblJh46VwRsctEJQHILeEjwwEp6fDP3xv2LihH2e3Ia+OcG
XsQrjDWzqc5CaxPk8R9zBR660p+2ZU1a/xmO2rxz5syO/GxXCtVScgDF06E0qXl0
q8h+IsV3ca3QpTi2GeUATftc8P2uDOCJZ7QOqIQn9AAFa0Uw4l1/A/zHrybWv/3g
JDAbd+3HiAIS9ZIV4dtweLJMwcnuGSoH5gl5hg7OJLy5K/gTpA6bqh/BRiyqU2yV
DEAD/SBiBLggLllvFc7ShWffgO65GbgSK8VDXF97rynOOVBE1woc5YHdgs4TsqqH
wqr5XRAe1iDkYoTgnihTTLaM6ooM5F97CegCLtRydZgGc1ObSVygK1Oo1s7ugIxU
/6YUdooGkPlJebIIvwIN9lFtzXTdhQPi3v2skVGkgh5S3kv6zFQMyItFu4WjDnsv
cGo/vp2ruhNadoJeEthw5W79tgK4ors8cVX+yv5+PhfjyzyL73iKwQVO6lG9kVIY
kg6U6tNCpHPKwh+xVOs6iPXxXCJuixVnGqW9KFd+uDxGJX6pm3+RwwfoJNCAOib4
WFX/WBNUASS3VGArNQpa2lUAx5sur6NBH77yRJgdiNzIbsMbz16/2fLSlher4oVN
Ljq/XqiobnBLtCBBOZQ+ultukeqRnKRcl/IF5SYiMO/pPZO2Yx4a41Nb8zZuBP5t
QhrSgnIBOTUTCMsjcxr7s1Rw6SCOsP63K69T804wEs8=
`protect END_PROTECTED
