`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BP4ct3SYyBWR+Q5QV7Z0YrKRI1K65iIwHgxLMREfssc642xgwglr0mDD1OFaOKei
sMaWTHm4ecqWH0Iwxpi4EuP1yPyAMRmnXh4XerwO5Ayh6gnj00Dgb0u4NJ0fr3WF
FfDQ10Zd9Aciwnh41kKatC1hiSu76iolhWfnqHNNY7MAn7BfolTNbz+1dCSivf0L
WiPFa16gW3zs1rtKrSB05jJWwBe0YqHieZUbzVF/gvkRz0+/jbBd/WHjeTswu898
71yZoyXDIdQon36hGu5n1y30GOE9RkOqVTundfoEmTOrPh+m3/ZFSUgt63FO/5as
1SHKe0jcmTbgIXVGB1yHhBUKzf4RrX77ZTsvYMh/6EO1nS/Gs0G0Vyx6zXQzpiO0
YUQbKSYotIA/e7SjSv2oAPOo+9gik9+y9cIQg1zzf83gkJsPyIWTahfsy0KJEZ7G
XWH6s1jyhb3U7sApgVmMZ5bwibXjIxVuWGejQV9hyi+ULdvsfQ1jMel5Cdrf51u4
E1+RwX1iGmx06y5NRcWeJ1YGfVXtaSfr17evO2luF5z0v06FESr4pnRHzHYEdPOg
628uzX7beer67KdlzODRlxbpAEgHI5A+knKbPk0AiDc=
`protect END_PROTECTED
