`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8E3ZMolnOWWKGtHN1SdaEa2FXv1DgeF3vgYPpCsutrs+QyxBQRkssWSVDgOVj/yh
6j9iNxjpS2wgYH25Qs+tPavT+43ma1+q7NUIc0s2Uz5ttanOMmMwN9foNsJxE5jX
fy+R1EumORdJoN0GZHKa4rkj4MUGBRvjjxq5jMPxqPJxOXjrwwOJQATwvf6i/71Z
jZ+CJQvRudXY4imhM9EP8iKszlMbT2SKevW+WAjf9OAEU1TDnjdgxQ6vPx++Rt3/
cnJhzYZKBX2Xi322tWrVeufOPN8MAK0rRNDb6pbVbBwAziKbaXtf/snqenVlY/yH
hDpNYhAY3aUv8vXQXoHJcD7zehZMB8gLGLoVLm625SAveGnib7wKeG3w5TGKwp3D
PYsY3pRgLQrG8TU4L2LpXqkOUF+Y7YGy7JtYRNt2AuQGqDcctlPEuYrPjKpuiPkv
XYokSfdcDGf4EGDlwswfklsE1tUbjEW4i6+EYzNgHYe1NcMR97caN2lBM75pYLmm
3IDC+jZ6SvIXmHjZCH7uH+1dbbak3fdxeecz714Zt6+eM80wlQS0BtjAWjRAvsQ/
LuqHdqnIxMq+XIHZNJL7moYy4VF2l/R7Az8AOViUwONMsUNphTUbq1ubDoW/px2A
8CUfhISd1DVd2s7FqA3QME7uvHrOZEvGfNFAiCF5hqQ0bgGGsFHiHm48Q3Zxw9kW
7tK+et8a7rYQrcIrTm8sitxm3s8Qr5RwTD+U+0Mgj+I8XMRKHjhp1Fq/Sbgk7pr/
0B8z3eksdjBqjN9w+H+P1mGo4nndIxvoy7mpDWaldMhSLuvbf7fyX5viHFSEMnFh
`protect END_PROTECTED
