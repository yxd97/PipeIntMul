`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xft0aF9FvvgRltf2LXzTMc4wrdAUZNwqHbMUN1bTu22NgfBUPR6yPku9GyNyo6um
o5bxKhDVbYNhswHxlae6x5GaudWeKM2IFkG1J4LBSqIvu1t9cgySxY4ao0XwyMSP
Eq01IYC0qMwG5RIEKy0S0NBYUKZAyqQt4r//J/U8kK+JDYAGoBbRIO1EXkKsHg2D
ZH+Vl28kxczLKfqzHuPy+OluVHIrizqeOHbt8EdGHA2qQ5rUR+vHuvE48vpKWE3L
c5CMeYKj/B779Zrda2Hk6KCe12PTh0fwuvi46PkoVL/lqRxAGuAMqDI49suRHPpA
9eOZ4ErhhxywT5CR6DM8S4O3dRjnwqhVLXRxmfiVm0UcE8pCPk9PfLTcm6pPyE5c
oDvk5+8tX3uriYItl5Djenmg8PXb/hwXcjyFg+PqHq+1IROQ/+kqW32i9XuwUEy7
`protect END_PROTECTED
