`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOr+prWGMb/6AxdiD8mJ3eGsnd0TbWjyS7BS0Ra5NRuKVPz6RX7NJ5W8CU0SS2up
I+wyHg8BYGyvuk5GH4fCp/itLdwvRCMek/rv0JRecUkkyi02ImdLZAMaBeVtbrWX
fYIVxQU/rocT5wbxi37ltcD4ASQjY58TUNj8eXeKK+pl5mwuIoMhz3XzUDL4W9g5
2hoXML+0b1gi5LOvI1ZaYRcfOC+QeTNC12Cs1G3pL5yqdP73PUdz1AMqxL84Ts1b
hDWcCJrk693nGGx6VcGO5251a3ue/1N7vsn3hYryu8L+2iKMFPHvkwTYU6FgSXvH
pQDvFKM0MWDxAm1ILETnzDnACfWo7TaZ6XBP3LW4g1Ezk0xJkDROuPiHUSF8P1m4
noNi2N4PuuEgg/P9+yXBDZacgnUAJS6x7IamKy7mAETy+D5ijrJ13cxU7B89Osic
vcDHX6n3i0MYOilu71fPUHX6RwaIm3TH6PIUOjtHBxUYKihst7vaArm3d09pqKYV
Ld4pXM8WEMn+jxLREciLn5kKd9pIm0oRiLblBL7dv+IXTCE7SbBD9jLrNYVZ5Pup
W3W6aLb2SYgQ/8pWhVGXmxKGQdo7hRn7AUOLGXmvOCQ=
`protect END_PROTECTED
