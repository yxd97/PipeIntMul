`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c+C8EjhXGAQW/lGmfprmAdaWYAGkOg+k21DXoNsfuiRj8zwfpjw4vfg5njEZszfx
vvvJxGBOUG4JwcvE5ilFAYtBdc4iHSddyS/4p+Uj2IV9MD6FDKd5im/mMNIbjQCk
U95p4GT2ac5kGlXwd0lMUJAHQEzpPQYHLL0Ha8OpjeNFJBEtZksgO7E6zKIspkSW
QmgJXv866tUz4nq0P4fYUIuB3Ka25fZi54LigiWG4uWGRoS3TfN/dxhpSrlxy2VF
KfkL7ARBxROEKIx837HAhFj16bJQL3XhvEkJfCMvkxH4gv+PTygVy+jYRkQeA74i
dTDKBV5GAeq39jzhWB3V/YNDIsCatc5fLie1W0caYLBGWP5Iveog6FWFucVdD+Uj
GmmQWjGnV7ZDyNyTexF3SdjL4pguMkVzYluBdIWnHVfCr9Ev2hgtTjF+mQNH9euN
aTU+uOyik2YIOA33vOIiq/NsQHXliv+qzc6pL0/iebQIvMD2ZzLKb1a3llztHWLR
/BSQK0RJMLILF4Tv89vLwz6MMbjRCLROJucbkXIedDMY0MouMlYyJEYnj5ZRtRNO
RKsRx+GHp0EKGoYPB+NazrLmBAeMfaL4BOC3CFqN4Po=
`protect END_PROTECTED
