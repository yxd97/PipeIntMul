`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0u4vonzt5tWzfu7LS+Zx/kR84So5JPzDt7Lb6mZ71Ie1x/L2on5keIlPOj0V2vqJ
bKeUoD6yyFgGmUa+zeS3KLwC/5xohcFlz3RfazXD/f+37I1EyIRsDfhvys0muKtb
M40/sLGlWkAt10ZbvNrYR+LWrsmPWYr4TZzIxD1yKhNZW40QrAM1oP/89RHERbVM
k10fFT67pCuoBtrX4GYFOiFY/Y+u7Tm6Rua/i+AqX19VMwIXbjMrvVIzGAjB0ZDB
Pas733VsrFdduyp8n9WIwlIQS8pYWQ17ki6YP8uBzAf41q0Vf52mW+BpzeqxIRjd
0Mamy0Xtr38vOQThbAoldxFsBj8zpuVWa4ud0iKY9/ZGl/mq+ejWhlmcak/iyPZF
`protect END_PROTECTED
