`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNqniJ67e/LXc+oJmVwHjwt/KRQK08Artumey0r1we8itERhNtDsE7iAGbI72gp+
FumOfTXOtF18tnLGQcBuMc97oNd4+9bqhU8922jYlrKSHphXwNMUop5hNZcYibZT
fQ1GvzT9J1rXHW1kL3FbWq5MRVnMhtCiGdbyHpeXiLamZgk5LQVN1D94NEjjKJDy
JQYX7UfOg4Vqukd0luFxLG+DLfhtZFYdTglFOrU6nf+nbtm9UtXvT+PH6/gp9F+s
SUSzSFnHrnuD5G4S6pSSJtoK1mxTWPFAkYKsMMgNLdUzcQgfCbfWIcsmKO6HjTnD
DDFdYAxGSQGVZJ06567MiqPHVy2quVMFDvEz/cMkEhl/haFc4m34KkvM9JqOm0Sd
LgeUAyjxRPQTZkBQ8cJS7Q4dqi23zQsLxOQ6pmA6Pkjtc/8Y2WG+6fxLGSnYA9Ir
Ttk/3axYjBxKkdKHmD3AnTF4ThPUreux27Cq71y+i7EnhdemDwXUL32175nVXzTR
bnoehxGBJ4ENhcbuiHD5ZOXhHipBMteZfXEaHSaO1Eo=
`protect END_PROTECTED
