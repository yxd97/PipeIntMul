`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kRXqESgXMTxNIHUDf3SRxOHYpL+hIOp6NwaRYs2mZcpdnow3yGXY60X5cTzPiMJm
zeKfxRCfXQ8yRngMOdMKmYg1EWyY9c8jslvaz4zjSkBEvXOn5tqx5wDuJRUEgvCd
97VVICRuQHj1V/AditxCScgZ55s1/QGy9MQ/WZtiZV/7PcaiU6Y9fzD149r/sNrl
98ajtR8cnRaNDvfl9Mzxj8FrVXhLGecyOrqSMPkM3UiZkQlDwOyvkNiwefHP1exq
SeC5eiIAD5POV7f4Q9WexQEHYNxw6jyrIXI+/NWLQ93BNlz21Twb1wXaRDxHlt1P
DefAFR/LcrG3PUVMIch9wvExbJJVTiEuzNvvvEWbal0hUWgmFydov2Bfc87TZOzv
eE/iBwMVF58qBeta2OYo1Q==
`protect END_PROTECTED
