`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9u7WrljiKym3XIJLX6szv0o2xrm34ZtJ1PMAEcD6lezMWeC8Epi5l8bzxtRvsUz
64zkvLo8y0Yt9xQwaWVy34GFLJjpbSq3V6fkNvY8DTGGk9HuIGjTdyLvTAE2RRiv
sbAkdwQfbfOqjTwBvstUKqXbvgxRJE5jenDoL5xq9bXS3DNBNC5XkU2r56ZC/uTK
lD+7ZKtFHO8g+IGQYPUOdWwMfgY8tpksXphp4FX2AZzqzrKnhl1nI9BhFZOnVByf
UWTL5a0KTm+wRkaHKi6VGtA1vbvbvlokJCA8soRPRF4=
`protect END_PROTECTED
