`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LXHhLcrXFN9Z3JbD6UE0fMlEEfljGn/DGOAqtIbXAB87jA8y5wvxmIhCNJBw2GM3
8iEpB6ZtNhCGaWyUyrNS+4ZIBCtrDr07s4L0i1Fquf6vLs8Qdn7SYMrHhYX7wSnR
qQUNImfpaqnzzxBN8y2w6GXfwicaI7HzGOcnmXG+DCObQJNTkL8/83PBq63IlcHT
WjtXSgQiWfB86v2MqZR30ldVRfT2/Nv72lkUzVYccAOY5uiUgMDzl9MSPwIefRBL
lqdxEH7+ZlHY/FVp3gLB0pdGxtAG9Uwfw18rfxhvHnKFFbQqGU/To8LtlQxF2lmA
STXEfeeC3ZT6AQI9VevG9N3d46oQ9xfcFSVrJVmCquBKEEAVHBylU1HzkjaMpitH
oDTRTeuhIAhaz5rBiHQ/954wjEVAnTCFDJZ/Ut9k2wWfdiz2JDbgtM7EU4znZLCz
OIHNiyJOAYS9KBtE1Z8ncgCMyUkqh66l7pIiMBaJ5DL9QPV7FKVRzVBOTuk9+s+o
KIclWr3bQSnhO+/90uDTDT8fFHyCP/3Wt3zZZzq4XqfAmcsl1wLrDU9HFPwUi4nN
3eCok31W4Lttv2Dstv0NrQcvWuzNC1CQ5wd4rOyfwaQsl1jaEI/VWu3hJs7+3sDt
yu6IEmOZg2PZ1rQCambxw+awF17ju1ZTIxzK8LzZO9M5BHoKIxeidBjVSp5eGhh4
j3jIQIQesJLtw9klONakObFw2JRqF/lXC0BpHVNRLwi9OyaE4GvKEfPl0YT/qEWE
CD8GkZEyGYs9YQwen5gk2PXZD2WyWyOsv2aWJhtQZvXChLBELTRaFSg2VmuSticd
JspuwbLHlOK6iP+OGX2BbncKg3EY36QIPfcod2R2mXjE8G9DyhjHQiXTko5xREoJ
BbBuUTkqFzhsxGVs5n9CtxQUxvso+7EOlb7Fw+iZPaBYnVcl8nfvQzLVpz9pIhfN
pDrfv7Z9o9PHmlRFUTzVvQP9BviPky1EMv4v71QhSqacsaJo/QgssrRLHdwKy/Dd
k2c11P9g6dahahlcjbbP/1y7csM52cNJ1yU4UbsjSrrAg3XPHD2WlpvSiKoGpbO8
ymSGRkmJlFtI3xKx/FVK36hEcbH8VeBgHMy2MqWwXcd9QyhEbzvEIj2A9MKpibmg
cwsJR9srNqdd1P6gC0RQsa1LHXqXdkpEeCugnV7fq5mL1gZuGNdYA/Lhtpxii1+H
qZg5axrYmD5/MKDFNd5B3d7YuQQQ2SERycuTEB/EhhtlQq9799oYoHg/2ArL6BHk
3hTSnb8tkYH/n/O8GUFwUCtY/e1jpbak56IrerPssj2B2zKUECKrtm9Fyqyoy5w1
sbSJhSTeIIMOrGYhNKg4ZAed4cCw/Yx2tk+Kiz8gUCCEbAQPtiFj54k/DV/q1kv5
Mfh1tjlMRLcxYNDdHcRQXzomT5Oo3bfoU/mt+NH3m/BYqknUauqyWsnFeK02jwYu
pOI3pqRh5IBKteihSmCTghKAzzNYwhlYfmpQkDSEfaeb+NyYsVzP8HW4OlRwwJ27
DL/GT0BR7FyXkj2LWw+44HShl+xXdYSr/662UyjlOj+XJiNPw7Yx9QGGxlRhE52G
a2XJSs4b/PdLY/tp11f1run0BMeAjdxBZcOiZtNfZ+xcVv2edIhMP21z3UltEPme
DLu+kZOh9v0iN4UMdqBibHWBwKVg9Mf8ILNYsPbm4kujfKBds7aoUzM3m+eJVGXw
dU1lf3nIatQdJ3ruqUTXnRU2rl5r4iHKgaq4hE1oyTmy03jANGeBwj4TWL+UoNQn
GVtq22OaeIGLXOqkQieNEEH89aea8UKIF55o8FsCCMD5YzUT3OWGmBBvMxzkuHIs
rFO3nDfb4Yhs95O6ZCs1pLCnyTwFwbg8AHz5nSLxghzWrgqmO5qFyRDQqh4MGlZO
mq+o6xXhVfKnP2pJzrpX80P4mda33FMk2cJ8uWak3aeSV557XnhjovKazmvCBPcl
/WIwNyiZqQ7c4t12r6TxeZIJg/gBnkhnY6xi3UTRenz/uYGhPIHTaMuYhX+IRw4z
prV3Frh8tmkhnPdVLcOhNRQPOmYM5SA1ADxqJjryBJlIxwbUMt9c0+l46MPxmqZY
MVf0Txwp0p15LZer440z1E5X20rJHC24kwlUoYxG4v6h5CcwgnFDncYGAhwObzyd
t+0VOh1OrQP3Zlt1ehSYZH7bwuomm5jrxKcntfSZ7ZlIhzzaZl5EqFVREacm7OzN
OH2ctT8ZLfAe0zUd/kWiIJsHW9ayVlDZeSoTrCh0qInOmeAzbl7EQuHdWkqJdCid
fAd6+/2bTZjHG55gpS81YuRvsWzJb7DoTLYvvJICARITA4bE+HhClYGFw9uGbLKB
jSeH0F3G+/rwwPO57VjadPA0OQ+JGBPrFYyQ3qUESGV/XCopFB3YT7M94upRdLXn
Ik8/eVKj1fv/TKJ5P1hswBMu+mM2DXEVtpvAgD1G4bcDvz+UyNVFmdRAWc9D1Hga
FW0xM6xUpjFVTyn1OOB3G6Hth6gxwN1mobpGinhXzfbyeWorTj4AMKpTgkNSwiXZ
avegAAXC6SUrgQfqq6JjKNKoqja7BKsWmzBwVQKZhIe9w3yM9Nv3kQgFVEEgK2bH
FD/EYTVZ3zzY9HACgEve7rZ4hTHPFIpj+iog7ATuNUBjQOa3jos+sHs08gurxXQ3
21Kx/wmcEAgYMJPPmzCN3tlKCmJcyNE8CxtVvYu5ljlEyo0koNk+BmuscDACI7MB
36pz9U2jszPciVxuFcD0tjF69mK0Kd7g7uBEzhO4WxLs6VNM9U13pyciMr3WufDa
BBkgF2Wqa/FKoZ6CuOCOWA37wCuuJN/hXN/EcS/qM/UXTdNK9J8YNivYz2fxeXq4
Ma2VIelYbBO+D7C6p02ADADE//R0OK708iuZCjm7GDk4uMoySEMp3fUI/qbc8sWg
IWea943ouLsXr3ysP8JOnO4j49RFkYLC0JnpDWvHcVRNfh++B87BGSD/db9YEUdN
qxlK/jhIfpGuyT3kibxvzoZ3Sk1Z2RS68wCZbq1zmVXwMXdV7Lt+3aH+3815t4Qy
zIT5fGdGe8++divGZdS2IHAKilPUN7rXHSutX1nwLOekc6+uKtu/z3gIxtqbLoAO
WAaXctEek+BRuoW0UgPl36VzgRcidA8uwE42GsksvU+rYzVSWgIdtv1DGMY+c3E/
wFmCtVVEo3/D11IdEWG2pgJKfhy0q4g0kuuj6+Ml4izW3SqoeEZpQZJvZex8tubS
gkFPN0uf6+QaKUKA2sQCLG4elcRwsXgv4wLYbM+NKEq2Qy3OFTamH3JaH7d5Fe86
gHLQ9j1CXn44BWCLJa+iVqgjVPhRuGRWNM60LdoXLJEv1C9worYwRu6apDBsT8gc
yjo1LfrpjyDPMxUOlr/Vc7IigeN55ogoJEHvO9bH2w7GnIdvftHPgqMpXbDhRtvc
3ayW/K2dsto15cNcCtaVyKlt3Kze8BW3queFk/sWFq9CGKFrj5VYsmmV/uCJiYJG
nIo4658EM5aopXvxOGlQSpyVRRimXLaWu4QlPCRcj6D6A44IN+8Md7iaUSHExwcH
SPlCyWGTjSiKS/BRz0hHb8oGvjrHw9qbcmD2EK/2HJyJddHubkzkKt75qzHiVFMl
+cnryxXgLqv0VZmgK3GfJXqOolEfC2aIYAaW3Djsw6V0n4Q6JFk3c8lX3J2h+DbZ
z0T8bqh1OA9q9oRqCGqdbKTf7a7dwfoEkdGdofSwbX5ux1euy1PMxq8t/zmDzViM
HTdEneX/rpW7ncFSTRAksYSHRAPRjJz9sPLfuPhriImhy34s7w3u47w+siz0jdSC
F5o+xgjEWI9FZw+Rx5B9p2tFDTIMAzMwG+kxGhs0r22uKJNSY2dfApS6sYjXWCYk
jgnN6/xUegem5QLx6Qb7dykdTtZe0ykxlsOCjZ6g+wnHZD4INtCzo5cy+U3a7TbP
QTuFVvfi47lOLko6QlFwxuzTjOti983vKnjk7OusXwdPAwpCOHAX9ACbdJZrXtIm
YB7usqMY3AwI6gcP2Hi9bowi8vfl9nziQElp6V78u69hwYAt4r56M8r1KOOgCARp
WMhAtfJorU9HQ9QxtWNaZKMP2VPNAJAoenLYrdatlPeoE16QuA2dMj6FQ2g0ffXK
ioRnLdU7x/v1tsEY593x02CWu96H51jm7jMJJ2414bbtPFL6JsPmFDMmZY7t8opq
sV8h2JhB2alQyvsDGibrGlRmbRu5LfSHJAk/UOVCljdHT1KnXMp5HIF951O6OQWW
ivGOJIlpPaDziG3BnqkCuZf64OLVcz7pA0+tuwwPNz3T8piq7FUugxvKysJ2bJc6
8RD9AjNpyd0wCT6LizHZZ03patCVRIUjULfB1L2BUV3/tQLA8ikslOq+RC3nikHq
y/VMsTJJglP0Lh6CDP0yaq87+fLVFATCu9MkCnjtnikeLvcxcAadnnZc1l77jQEz
48sU9TLoJcb5gqfUKOYqYFFquFDpg903jiqpUjwcRDu49vSF4lc8ohTQKyiHfaTM
CeojbPwM4fSL7Yc+xXX3j4MIJlH6zk496CNqvQMxGkL8MLVGYa58PCO5CkA+rsN5
5eQ3lzL0+RqncIADXRFCZSeJdx9qOIHU9kbp6OevB+TJoCp5ReaXOCSNE2+L0VI+
G/nbURL7AbLthRrArlSImKWi4Ddy4hz8zn+WdyMEiy2mqfCz6vtwsTE6QUs0vhGm
8VU8rLKkkux4umbopTceQ+yrxyhlIUOoL7LZCflcEijqHU5yDLNBZ+Mk738UaV9n
h1xyCYMHn+0xiecO7xiFtcx5/8adBuWNX+97/EMt4IHr8g8+dtTvooqq1wGivAdv
87r+neC9nEVrykltEIsh4H+XOOucoZ0Cf+5S+FbclJBD1Y7ueRABKzO6HDUwi2Uu
Z2ZWSwSCITm2c2HPv7vWYSk69h6orZ9vJm7umo2/pSOZ7gIGnVQDpxgAWmskQBmJ
hjuv8YfqtnIZ05vcDnv2+NVVy7dfL0OA33FGXNwN73itDDimPWh1PRw/knf+buN5
dP9ARyQI1lyg8aHKw0fEs6mSrLvnfeEgLEI+6vBsKXkrx75UzUJO9NzLjO6JkFT/
D+rxZGZpiilVUXDVe/+w3mqcv9rAm9gprnFqvxOQzbPZ4hiwzvp+fFkcEiyHoNNO
8aSL0iVuYjcJ0HH8OIde8i7xjNzp1TIW7xOqGrQEi9ZtudRSYden882dXmCfmNJC
1QTzDyR+gs2PWZQ3Q+a4cjN44b/HoNZrzVTqyF+uJCqPLeY9rmalYZn2jCy4RrIY
+8QduAzxmWC0Wz8YwY1yu7VKdLowhGZEBdFXiK+S5L4nzd0etqAKvdLigv6HavqK
MouMvBrZESZvGFD+hH0NKQzhsdeHTpEc40dXMQoL18I5Dlm2lHRtFPo469p39SpP
SpgvjyO4kJbgq1+1Fra7bcrt1CrLhFNySBtnizwnA7lI1bCnyw088IrbVI6D317Y
nGii1xe0lMZjE/D1gA4csci7f6VQCh1EkMOSGJpJ1Uorxd2r/Zv7i1fVUnpQ1Orj
C7l/CBLF79WPZ5OuqYkLUvKyWo+Wq7OhHK8eqDOLaecYBsP6/8moeA10Z4AP4dft
O88FskmTpcoiqZmxvfvxhrGMRdBj0936KGP8VD0o04Y+/+uAKwShaTepJdYbsJHc
Gdmmz29KP44ZeS1gijfhpZoIe4HNDn+Gyidg3Yl8REQEFdLKGxFUjsjGeUCL5rKq
VYxhOkguMzI+kja0AT1lMIFMYEs8JZ0CKS4vwXnH2rdCkoMD5lYUBKUI/TIhzmbO
6lV1nxed0jjCLqFm//iF9q0u58gsDVkpfHwid+BRS1xOkTqRo48SA81kac0vj4PG
rvLN2Rov6+zRPdVsmhWReKrYj/GHRM4zMp23jHN0IV+mN4PIS2tS6JG6KX4gmQas
nlZU8z4yNmSsK9LazXBZ+BZrjGr/94P342NPx0hS5lFki019JdKjyWYIonVNMArr
6li3pF9uuh9ziIeUottUMI1YDorvENuUOiNuFOiYuTFo/KAg7ru4VtpE0KOXsZJJ
XI14V0W3iDtlXe5ZLbUnOmLhv2jeMcxQOKAVEy4uzrpf8NX8TolPYX7qObkMwaJE
a5oVBBLgIdZsV1jZxke9xKrPj9uaaIO72LXL3s0I2S+d/SoG1DfphS8PNafoGAqe
W8w5fcMmRY3B9lB3fCggr/4bXsVcVEIqaBSOYtZohr9eMP476aotCjE93W3A+gwT
DzUmXqtzzTfHuO1rZcamwK/v8B19U0TXnBkRzfsiswuB2fjBniJ8DiAk1yvRcQAA
bsT5P3BoGNIl6t/I8dJkcX4xUt9I+7UNXQ7kbm8k9dMRLI1QzeAXtxh6CEzJjs2t
zyB45Qi1KJDJo6T/P8C7U3eZaa14JLdO38gpFf7QGt9bzJl7phaRMndsfWeZqYiC
2zmry81bZVBX/EqSx2sBBtY8T0bvunWo4DilIPCTSNcmuxyKMn2JyB0hzmWC5on2
SvXy4EmDXTABT2vpOW/TzxGL2xzs8vk5YVHNFl5GtcRdAsK3F+VymyN1u7jLhWUH
U4ZOJOtrrx/inpFyfEfmhT+26jDm7FDpwnGmlRG0mCDXcx9vSXwkr5wiNl7Ow6je
2l7+dlDCddem67JiIUQJD1euo8JeYYgoewi+E38RtPCBydpokyos/xvdQTIXOTL4
lUaLA//+LgoScdzokR+v2+hZYPL2Ydu7KFBCb8eHmuwolX589+R8OPwt1a21OAdT
P31JjlUmj/YOS5AUz8E7vziUvpNbpOAMnCI4HYfAFdXVnq89MPcEATGnZhac2lNO
+pnMkF+1KMkbHt49XHOBcDBrAOx5mYn3eKINVl6XRcSaS2j6WU9919v4BzMsWJgL
/e0GYb4vdq1du0YyiISkRXtv8ulf6rfKuG3f6qhRhd6aT8u8zcXBSZ160CLxjp4c
dqdASiNyNLTrwSMTQwDDxe+wX1Qsh3oln+kuVhCgd9/doKhCN4GKbMowx972/jBt
KNvFSRYEQmrzhtxQkYmYoC9RbyxCaXoeb2upgutYWbmOZhl0Fkxcaynzi5BBxUUp
OJevgt/SHzx1zCS6rAs3tV+MbaWvju5nsQzcIG6FVClRIVDjzmHEXZeMc2uKJSBp
H0e9vyrUQUUbclSv4QBDxydEagWNdrS3wglMFRyR7EDP7hinROJOC+yIWdoKp7sO
TBjgXMsotISHK6X4NYmyU6AvxIQjhKUjPO0pMHos4/qG29osC6cGrr9NPDzo8iv3
v2kVOKC2hf/wd7Z2gqaYTiluB5DLr3+4mOBDzQdVbuqKAFxSRU42WibVblrLRDBY
hAIz4GMrztGSihj6cFd/q8X7sUcg+66iYtaOu2KzWfo9rp/ec+vyxXrvqz3Cp24o
0GSSCgwnxcPFdk7ncUMx0qdll7nRtYIacl6/KJsz7nVCpDtP/QEPw7IpcfKCf+rT
FJtWsEFxmaz2a9EM6zsNn85KgkOorgBSrnbvT5GIyFi6MuRmRA5ItfmBRLpQ8Y1Q
VJT3GZAFIntkYMOHCnKI6RosLH2uLmh5+MV15FAa2jPrcARODMJpim8QVyyWOCYo
Ai/y029B4CLy6JJzVcenKEFu1YK/Bm6OZkJu9jlpkPjzwpAgLJPFnVBSJUhDSWq0
DwNszVUEZEeWPXiznFcpAJfvfINvwp+L+GIP8F0+QMS/KC7D412NktebDIeH4Uuw
twweTQhmOhSxHz7UHcPJdja6qyYpUF/5IgqnoKZ8cFcHLHLQFRvguOvPDi2HACQE
IdyAzpatOxpb4NYv1mJdWIRmI6F2qRNaKVwHUzeDcVS9Xb7v58eKlNDWYP2/4pQ7
UwrvT/YAhzw6ZkRm6VBZqxYt1fwPA7otguPPWe82F1Tn9nqMi09IvUqI6c/PTsaI
v+9X934rK5JMm6sCwBONjF2Dk1QKeUNwh/ja364eY5KwURo/CXC5RkQlPmfq/TML
C5jQzpzTnRRvRy6vY1rZEs14e98Vu2bVUmlffQBW9Xw+KTYLBnnkNG8sBZ7TqaQe
pfHwp6mAqflZBf/4Md7xTmeQ14GQD8wVpwdlkPvTG+4TX16gqJEuQ621K8d4IfDe
78VTypp44doPelM2idLMrIl7wlQQQcdNgEauzoCogmyTxR63SoTzuhTHzRuYFKKS
1S+0jwKsidG5EUmdA1qKApmYSwBKKJq0W1w6nVzBmWPfPJKegX4EMIC2GAuXjjPl
GioP+KJtwJvKRmKVMmxXB5LTU0NfLS58PmmgkZmeoBaoA/ZbVYF6MOja/FE8/+EG
Qv3cZcutVn8ZH6eQnb6bvhKoonk2KKIxT2WcDSeEejm6r0loekgbmLR9OXcLEXqs
H+H4iMDQiv1AkL9JM4FG38Ey0p0/U7ynTOAxrEnrI7Y5rAopVV/Sq0ICIsyeeJne
gxPnhW7HVScrJGxAZ73AUzeTx6l2JxkCguW9VMpIMYBG2kdkyOjN5sBzWeFkZLLV
svNLUGfiNRrfx4IVNeRLuHydf0nbfLxiG1TWz79D1BjCTDOmxlJ4/RU7BQ79P+mf
fuVCPjuOpmtF8IFem2fWEvzsWqnJCZbY9mfLcmJNJqB3tyYyGCr6FrX7bvyNpj7N
nMIlqndP2NmDDrOlLSsAftKPutyaY2UeZG+tO2eq38U0mCacv6MqdNBtjuml9jN7
HCnsou1NoRH2WmzLoM6Q0D/B/MVFd5cjv3DXuzOkMDY5IWX00te3hKFYItrtkREx
cjae6jk3LVUhIY+aO3kegFonMk6OVMCQjj40YNfd1kKVOUaguK80pvC77FPjGjZF
SR8oqgLrWWe+zOj0NpjxJLrM8uegqk6z4LHanbQ77/uHaYsj0Z2v6GRchkNwkDkF
EpfLfGry5yxyz5I4WMcnjnHQF5ryt5RTIz8fxj17XLe3YPKfRi7CxMFlAw7bGPcl
ZOnx9hA30QSn+VBUtYBO4a2Jk+2Nd2joGdjBScxltrgSPQwDnv2pNaBZ1CNsdxE+
rb3zd6jlHWtsvS0gc8eLqBzNI9325rY6UqbD1gXxe+qs3/+MT23MEk2RsKAQJilm
EOQAzX1+kZhLvv1HOl6+HkaC4GwWqvyTOb5A+LVTr2BfbtfVsIi8bNI3K5u87/wI
AZ9TLfpuljyh4vMqMs0sQ3lIE0geDos2xLgk3/t4JeuhFLrOu1+uhALvlFOiQys7
PRqqlpW5wATJ7xNMAcZ23OaKUKvOcrE1mqIeY2b4bDakFp0MVxrr0YXwmao+7ZGX
UwPkYEHkJLcQeiKF0xN9HpVfnkQtsWOBU1kIKJV6/3rhYiB4LTvHzBteY+EEU3lu
+/dLfIMuX6Kac9HiUAGgiIU9q3/voe9cUZL69IrT2VMsaBSLjuC23V0W7hV5fzWg
VSSQmXuEBTbIX30ZEg1ywx+8D2izHqcqMHiSNbqIGiRtWUu67hPOu3pQH3lBj2Er
p3fCAVdizyhd75erJAP/8W94dX0z8G8BMiC8QuYhwHAJ+0ozEbnkQHkiZJm9Nqeb
TVC81GzpTUo6QB1pGXEFsA8syunqxqnoH87I7RCuV9Ll57ycJ7JAkxptQZr6fObv
TqWYAUBZ4KORnFMUUDPta6lxIBExUK8LQWiskGNsnwRdvK5JstURlGUYJS50njSF
UmblcOTpPLJ48GmgkwIg8E/XXME1o189jU/LWtUVn+zw6t6v40ttXcXJfPhphdG6
gtNVKUODoboXl4i1A4LxqyntiVAzICPTW+hq9qE201+/0hFzCJ9Fa5ZIxaLcRTUj
5BkQe2zPK6AjxL7DIk7OEyI1R+cyy2ppzC/QU4LiBvGq0mYmwSF61xo9AE4aRH/i
odbDbeoKSuAdnwahi4YpGVu4Hp7rKy7al2rhpDVKFJr0/wk1cKXoTAv+iuB55QSg
hNsJnFM1S9aMKTgsY/igL8Nip1FbDUp5vb/Dt8ZbIvWN1cJwzkU7G4VxyqvyCupn
03tYQxnt7UXr/b98alU3vnwDI00MauR9KoSUHiwImCmJEIgEQsUR3hPDbjGOk3/G
OGdfrBTOAmLabZhGAvTacoEvH0Y6UXv4WzxrwqraJPsR0+jpp0dC1Ej2+KLVKS2Q
Ov+W0ykvzQd3bii2Z+3WM63LyeOk9VDPhxjUuM7SDQ1m5wh94E20Z6qTU/XJd0jn
EDNst74Q0fSza88YsX1ryupHlR3D7qNarxUvlqUOOIiAIe4r31TJd9ALRS0MFhkN
BPlYRCbaUisdB8/9ahViG4zAFnuZoIRMR8S1BkPVt+BDc0R/qPXOZf9XmGiYRlLS
xW7t2sPmsvjBifMdIIP67exI8lwIV8BhVsnI8/RlAU70JGBiOGt/B1+GdRq1/GWN
yXXnkImBAVRAOqOcNrztm8Z00K+6sOoaPZI/gyarpOf29NGayS/J3+HKfR7uAH2F
O+RQJd7yvTAu1HXGtxwLR6cETuvAaPhI1cyJn7hDtsbB+qaTbRmG6fwLUCFQIRyy
2dEdf1W81BP5DoKsT4YfsTlmYv5tTtwKw2Kj+SHsf5TVZcCwHwWBmFzD+K5wHZQH
L23AoNEtEM+M81g1o+NGXr2JlQt3D5Jr2Q9T2zQQqHkWSE311xQQDl9skkYGd/gR
CxMyyVf78oO35bNbZ9+YUUYbED46Tc+pTE2hO1w0aZhrTJWxWvjwPQWLwoCn0kPV
Lt7smnI1yiY3BaNuVXzyp717Vvd//u+2eMrm8erKejsMYmvQTobD4vipZeb10Ki3
ljo7IHOx5lZZXT3Fz1m7Pa5TeWtV14QKNTKZ1VN49IpFjs/Qa68uUZZ4FsRQTVvL
Qa8ImYoJtAWyaCqGPSoBoBN5365hMkVez10ETeFz2lPk+xRz7x+eWvnlZxZrIXLJ
lfWJyYDplK1sI5+LfQvxrYJoiqNSx1ihH1ZHOMVi3yU0clem1dr9ZX2K8q6ZoV9g
r15suWDHwMnl0867gslI6NzdYsebXwSrviJGBi2FDFJR/AU0FTwbqAmLG/Nwh22U
6IB+3GOeJCCoL25madW9SBKp/yNYX8imn65URj7a44MOXKFtfU7HlPs+HlUP5Jzc
uKIOcvXw1mA2zJJzmsMpK9JeRupJ7LqIyFLTLQH8k1gwFlGsg9yjt9Mp+nMLAZ+N
JlVG+x226/GX3C9ERQglc80zc6fuM3IiJoKcZveWZhptn+5DuKBsjAdk/qI4063O
ZL1/trt1wtafoS5/JPLAw2Ufddj1xGpHvl78gY1y25g6R0tuYdpQZW5JLhHF1hfZ
uC45wPxWVF8tBDjKHAJ2AcbJMIk3Gz7zzIsgIkH4BKMQYNCf8+Po21MnxQjsRxI2
+9FB47t8lwV2JaSTRhh6dYSA6+hsrVvksxGXNig19ytfCj4bEkOeYyeJfjWJm60F
UnVr6cyTrYQQtErzkPZPXy8rzvX8UHUwy5NZF9Fcmt9CXfUr4xJPKNDTm4ZOeWRr
DdQP0U5JKVAE72eqvtZeP/4rsV8x78aovdy+GYt2g3ij/VcwfNiEPt+ewaWDfxTv
5K7v+ZO0g58DIIdNgMX9vE37SIQhosWx1WLoSj4veD1rTGOMsSIxrL1j/zszhdkc
B+7sXT3V4B7EZ8Ean9y66bhm0r4e/o/GP/RlCb6vOCZuYm14iLYgW2nVO6WGaGpx
7cBjGAzLgGxZVm7sHxhOp+zfS+Vcx8jfvL5Y+rUcFM55/2cUgykvoYdeMhNEsIUm
6dIW4DmIarTMFQCWLEg/T0Qieqm4vACdcmWFz0L7In1dtVlRmslNiKCkDXwEIYis
o2HlHZXEgB9zAXmz9mCFeBRJ2rRegYGVFb6QR25yPzIQe+4mX6Uas6GVbVcUHuAh
T4ILm7CdOFnudGVyakTg5P/EM1d3XeK/h0lB1/E20p1EvcwgWiskP2Jf66HbKDD5
zH/jhX9RkmUS+r66/3ptbyhrLoF4S/SJyT5TR8GRiU62JQX3PYwFsGZSobT7w92D
qu1j1uVvHXolwlAinxdqwrfNbsgyCRmEJUP0aB5ukCCz0MC0oWqA3hrGtx2jYzK2
SdX6Nvaq/6bseBd/vRuLMm95Pq7+ghk0EvhuywF1vs83b9zDlJ7GQPkLmTxYukPc
DqYTJ8EH4u+Uo1EiKzOKAVS207ba3iugYsi4HtuymMjLoHbdBnZqxyqB1MKKg61G
cf+DI9/Fz7o847vSF6h/kdAR6RHGhIWJKTsiBFT/OPlaJJUjoBY015wuI7TbZ9Jq
4LtWhMtHMJ8ZENniQQqx/yzkLsyGV2iQn2dDG9BwrxPM+qLq75LuaqJzlvIIXvRe
TgFUZk+7S+5/oDw0tGmn4S6OCSMNoG9yETUEN5IRNXxrEIPlAm1tfZ1GviTiZ9el
h8gp2EkWQYuU1cDPV0qlYzLEE0mvmDxcBtZT5E8690o8ylrh3+Uy7SThbwZ+PyzF
fiJIgWla7GsOxgFeKVJqlNgfqdxM4J9AqxYVUomPonFcJgiYp9RALXDuz/vdA7TL
Vrp4A1Gxc3dLMNAxyEJCpLYYqRGMzVj6ywirmbv8QQmvtupSSrd1xO2wj+y3q4gV
ruP0/POGtwnCBg/gdkTBEa9BOyM17a7PfazOsY5O3ZSlZ8FDCFlMtr+sPF7jTJ4c
ur1olmKQWywZC2cqzc88lgaMFN7RaMAgbVaYDgbIdzHLmR3aZDJg3DQegV9jcvT4
5NyfMjvHiWYN2tAgy/WaHvqI39f9GUue3hpZmCJEkum530+sQ9+g9fph8ePSegRJ
1liEWaV9ZuR6aRXyYbUT36EhYFYC1WE0v4keckTzcMoRAsfb0YGMecBcY+g8nTQU
NlOF+nlNr3cKaqOPJFpukx0qnHrEMkCOJJ/KIEG8Hy4FTP1FlCCd1tECLrA48Xiz
vtfgmVDUBdbbB5gQpNzjT955N2GaVZ3WJ3verkjqo47jNmEO0OZl0H9IIPrbDHxP
NCpYa1q7nkUOGBykOKNAgQHDr3VJL7axg7lpGd8ienOLQorALycOpLiecO6HL5Xr
Qh7KVljN8vtXMQDc5ZAJ83iUi9bF5BNwJWClYShMSxOyjUyLjUVKJuKPaDyFgeCk
jRJ8F/yjAhNb93/ALHEDcMnv0qjoDshNv/F6ZHBHrym9Yjbtbh3jqPJ9dDcjII+E
eaf2Vm40Co17Fy7X6UvNGUd+nSEO8XMJTao4v9Vtw6b6j+jgxJFYhJIHGqi4MFZI
NxYF2cz12vU9fks/1y0UU23WmFgqyVkOywF0nVgI8PnpzCoRfuXdUAYRB9E8+FLP
XKhXXVj4oNkwqwC+TmuBe1E+uAfuL5X3zs8zv3DMHL+X1AsssDkszVD02HhawDNV
1zyhnMe+XLf2Iro9R9c0l0/AFN5GqDIcoGpaZQuKoP4P1y7Vw3Po1/+nMNwq/CQu
PZdUnHsEJwm24CF1xC+B1qlK2wbzRIAU9V8J/yOrD5/LdyAgXHjjqzm8Hx+LvbpC
eJhD9buyHRVucLPyNECw3k6KV3xG4Z8exiFpAa8zyMbRx+35ujHUJg42rBOTD1Cp
ikJlaQBXdRK2cp3ePndFcBIEtD8mQpiZc+cRx+fUkxxsxgTwajloQhiiohYQ2kqR
cJVZyMZJOMoLI5nET7tqzGYIagjTq0jBqQIoXYoc9ntjRu6AFITuSuylBl7rOcY0
KWf/OxicIjtVlvhruoppIQa9Lu63slki31dMGjvOvxN0hVdbx0d1ydBPUQUnUjhn
2064643Q0oil82fxM+J+oPRjRHrHR1pSbboZKtilXrt9aWpM0IdKsYBVhNHJihJ7
XU3IMj1T92W5VQbIRJBjfl1iXGlW21m25beB/ZSeWdrDqiqV608u8k6jeBtTDzGz
V+4sCIBkExo1nnJWGkdEhIiOzqzxbOWOz50fXN8HABhohD0ZJ4EbYoZL7kXQzlxQ
7ghZtwe4/z7gNKveKFYgW/sLbzJU13WGJImaAnuU+H0TFyAH5dSLpxLMx6469rP0
DZA66lYxp3tQqTbQ9mVKxFgmtPB6Xw1zXB3JoxsFInu5mk5NeryPmftwZOihT8kI
o4wHUuoZEPLrFCIAQkZ8V8sqC2aHZd13hUY1gxRnH4GyuaoMEwePRuq/YyF3pbvm
uWU2P/iTGfaCdF3/wEEqycTJLf2pmNAm3l1BstYsvdZ0qEuPFvCBgtylBr3K/Sus
VvuEbAuhfZ9VwFXgZwWwbyItzK8ANLjfFNke1bAwlYMtWkjR1wQasn/5/y6vjz11
NaRu5JXCKDsiUXCI8/LA4w0Ui23dEF6mOCwT+rbKotgTTgmXviIwDaDifppPeB9k
fv9LkFhxnFeVBHcAYfPUhS8osVrQP+JfBg4ryk8EkNmOTb68CbQ8yUfFoAzh/Dn3
AGR/pLTzfmoj5smE8NdUIMIHP0S9qOYn12iwg7G1FcsXFXw8JWg8rB63H/7hk9cX
zsfL+NWfOcLMHULZH0sVAe6QlZeRQ3zpMAZ6WxlY1//XLzKlh4+3J//MJS69hsz2
+o/1DQOxqY5IPzr0HO+bGv3UcWGuXGpy/E/KoiSKCTizz8ktia+1zsrddI3tjwde
pVx0GB+XIvj5jDwNsCzuU1Eikho81FELp877CCUZBcf2OnAKChBjlqjB2sGR8alN
geScnsgzkvbqRKkskXabFN3mztkBVNPkEklq4AWlBU++iNLsrgurHXW9LOESEMzB
TPt0yYzlyvMLpF8YNmwnDWXT2sf5mbG5kHVTb0oO00IEBKjATcyiqtv1MQAEyVs8
Iv+U+uA7PoPCuGR3GnFKWJHBgdaOc8Img2cDULhvPO5yBlwi2czFFlKVGppWrdzT
wO6Rvkn5b7ayx9S97fz4YQK0gU/sgoHXKupzxmAnQOcqfVeR+d87B+SqkyBoCadr
8ZZY7wxdaI9cd4Iaik6gz3Z46AlL0hbnFXtJfAeQ/lZLNC8gyInqsqJNt9ejOt9E
W8+qYr3362rqebYDfA41ZOVAfch0pwUH0fNbKgXwZIxZuQYg9IQvvG16eCgifdgK
d6lu0gzFd8ipTP3/gCJeZob+ysq66+50hx3CM02HDWtmXBINSXRbNGS1boiqBcH/
OIt2YXmlwHKenSJFeAbJMOsr4Un70AbQeqwiVTGddgK9bi5z50GC/m9QKpU/qvFD
zRVbM/5v7Q5B/8cJ0De8R81dnW/dY74XrTdTAI84ErXQ1YFJ9wSlRC5LOcqoOlrA
buNzNOkDA3rPriTvxH4HsnXPlf/QhN9k1CCI6EaAEZA/6lUYqD43Yf3a9nmEnR0S
fB8W7timKiP5ej5oqxnZ03ZPXxRtzQkf/u8l9Vc84zzmUgAGyUwApS6grPhdyiEk
pvGuLSPvcTFUlGYBoXWmLC38R+uLdKblHBWloTmcZ5nb2btDagJ2Cm1hPgPEjap9
hZ9Qpl/hclPKgAe9SbVJinOcz9QNnFGOvu919rB6WUeZNQzZY0ALXo6YX+Z1wZjB
uXl1brzeuZp+yFB+gvP640P6TJwjqnBYL6n2WBAz9E7U1PJU0xokFrgGG/c+PCsf
GSj1O0syfenXvEDxEj8Tvf181WzESzmYp8LwimR54kuIM9T+Um7qwVqURrYx2n5I
VCsNZWIHvwTZ7xRm3/O+5ATyJR4EW/b8JxRYEoZLDdFm07/97PvyXMqTTtpV6PYM
aH9tzBEJEbc9Y0ymUOLFDUvATg32xhw33gIvsCY5wp4PewiEmcZ1mBBLIY+WylOJ
oGRf67q94qhLBvYwDz45n51jLoGM9FBKh/lSFGyws0QAe5gAZn3P49PYN/LJ8QrO
tcISEGWZEy+MGtOJX9wx6embNSnvvEWfGjGRM+6fTEVEdH5K0RIv6YgrRusr2SHu
DqAFD+SRjVRkn4YYx87oKmbd+qHnMRlwBIYF+TfBAQcZV5YYbyAXpocX4Y17QuuW
dHqw0U7/skgXTLp9ajvNg/tXMYpsmq300s8jsYuV2XfqNjKein6ZRGUFsOPDi1iY
l9mQU6oceurPLtViNMRUl8F5YMGVIMXzq+P7u5me/P/cX1HmGQvJxgg/47gZP6pj
h3GBbB3T+8XM4kV6bkNCb33JuV8brE5xkSVaC4V8dnJ4N8BMZE0AKc1v4FI0YSPn
IW5XjJa5/h/Mie5kndkelaBAURxOddWFocygZ5vcVPSzvuzjJecqXFj2PV/hgTjO
a2JKhe9eKUiZrMIbLRH3M4JqmYlB7fw+9TjV3QMjX1Lo4yTQVT/xXzYrp/meIdZV
RzHmyl8zdQWQ3hQ5De3rcsMvLEqIPR5yyo/iMWHDJBFGo9Cz5vbLGpvGRGga9B8i
sQhEcw7U0OaXNsePuLHhSDtxl/qkDvShm/XP5GgCSIbGvcArQpF3ANgOPrpeXUlc
mb9dxOEGdxNngffL0U7Ym3t8EpsP2MwI/46NS30yzf+L61kJElKp424DWWiNz8Ku
xr2DUiAHDz0sG4MaUFKvUPSzR1moGHcHnBuLQZ7iTmEJs7P00zf9A584W+Q475Zs
0m51WsgZiHXRK2Zk/BRzqSRWm++SF6X84BIXph459MchF3rcKAJpmwClkUZn9jtp
1sOZrkCVW5yztaL62yAfM+IQBHLonuhLb96TXmpjLX2AeHzwFDAcERHS1MsWc+nc
mGMrzkVDEoS1/FQ1Zl0W8cUFsiSeGvZGGM+pDP7Hs8IK5nx1lKUjQZGHa2LLcPco
2eARQFX1PaDnvgjO6bCY1K1RwDFpU4q+qcn0S5H28pOiwx5llJ6iqlNeo0gxG4jf
F3CLKYovIuDSuPTweg75FcQEhIxYoIeSTeSfHnNCCQXDLn9aW41q5UpSB5ENrGGr
Fp7hZlAGAM1J/Lep17dw9IzE6iYvgs76g/ZmFBiUGETMb55+aFHnR8Gf4IDrB6rI
ljK8H4XHu7Zi01kP94zU/qIc666zO7Ovj6qfc35wJMEddzGjcPxvccWWmoduzAYk
XP9qCxn6gPpfCNmzv2NQH1wVoGg8IP50trv/TUv3IYDWsS7b3W1/zGAM6kFwzAGD
PYxIujZcrrpPs+4GvLJxr6WjVyGyUZiflAbMQ1LKm353S7psmEypGd8gdoZ/gn57
Xph0l1HOBTHN04fqNMU6yjc7oMBtxCDS/kBZl4dEWxiRN3JrT+/fav7/419U3Fz5
STfPT4gJzRasCwcRIFH/WMCDjQ7TXRXARfd7fDK1azXJk76bzWVunT+mGGHZUNl/
OR6jShVfREc7YlskgjPDmMfmQokABCn7VJINSaMASFOdzfSYzNuGyLAqK0Ltc3JU
9FYffdwJiU4QUqRN1UzsHvCfAxzdJhWFc/rxN+BP/oeIPDkfGf6pzst517kV7MPY
6JxwT4x938Psb/g/KGf6dWN7IR/98QkGs7Nfg2/aMzohTHocK2jujDceqogQvgeO
VihiGmPS1sxAGeXF3981hiQKlx9e/8be528/m+0SF1Cr08ddxyc4KUZpvbu2Y84L
SAYhp7pzXVWGqHN31VzT4OL36VC1vbhoCVIknAb/BZZh4LzadgGMN/nQSATo5S92
IaZ5vZRNEvGllt5vSChGLQDMdLmSPEAFWDAGmkfGmIb/o7Tbw23EOPQyIlzSpD1v
ioYpcAJqtVe3U1ikbFU6Htqx2EZmoSgyDDCryz9BxuCq0XGnn3OzmuAN5G0YKvG+
moQ9e+dEG0h7g+IpQo11fYqU7Xq5mBD4ZvXro94RsCfD7dExwp6MpsQ1owkPVEdG
1BK8TAnEEpEID+xN9Qwstod5h4JVXUe9UtoixSXdS2PMqNvozJC7mZgvtlt7+zUS
Sa0qULbChXVBs+MmgBgu9GLq0+mAcrey1Om6dAJXpgl3iPqMHdcfuSkZ9LiBqW4s
DWS1y1fVeZsJtXgmftyIsCP2s8pMCJBbwZhL4fut/BEVr1kOscr3yegtzJg4NxC3
PHqFDm5m2iO6mLHKxbuov0mw8kROprZqy2G53MuT+KxtrOYqKj90BGOmSWCIzABz
8MCnhONXquAxLK8g6XR9tT4DEZulv9KhTg0zLAv0UCxASvyb8gp2siv3du57vnAG
NsPEMHWRSLybbPxujqvARHhQ9ydGtTPDy+Petei8KTbSPdQWo2kaMB/MjD/napVU
A+SVxm66MH2Rsj+fep4C2RZmWeLI04o+KTk7XX1xKaf9+/6S9pzVKXNNSOG0BHjH
rQ06jm7pxScdnOvVYCFvChORzbatcufLENd6cRLnmsAi3C9oloQc5+CtI5vL2t//
oKXCCYp+TGEy9aCbA+FdYSi90e4axbIqWPrKZs8xRW3ndE0FNgS0mA6AntHFsALH
ixT6PDKhAPjpwYudwCzbI7UKwowqxwCPjS1CCeX3+AYWCGE65dobW0+QsczXOrZo
wuCXPawkPo3EqfMOuBzbE1uUJMBwJt5QDXEtfldR6os/DQENhmLWfPd4BXbxat+y
DcIrB4/mrzbnqeB+ChXCkDLHf8pBM2OYOfGi4W55tW1tcjRxG9QUWqqk4/nUWvUQ
DN4EgDGbjUHkTU8b6uf5LRjgqAJ2kVxhxuKWxTyDUIp8AOTSa1oXfExHZV/Q7zdH
7irs4Vwog0DhgHq9YQ/QJhtAUYR8USsB/JiNsHsd9ZYUy2G2wZCJGxIZd8jCxZBo
GuCSZ0PI4y4H5nu+UA0FHKXQvpJZnOS0/glKZtiJ59leL431BkiVmwAvc5VpGqcH
6k4PIM4dW5Duui/42SFAdd5cawERGg/u2ogcNit+IyVASqy2snER7TKW/lQ6EWMj
Cx/0w6XMThjPOiOHX2NgciVrImp6M8AgWhnJwTtAbN1x37f0U5bPEpb8rnKCNix/
QbASVBGYr3F6i/Q0M3DVM+sH3T6aomqiz1HkyUaj/CLJnQObIFOdbDatpnlYJ5lZ
118Mh5Tk82S3DWAwZqAQDy+Dsbmj4w82PG1rlOKhPp1XAOr6PA2mnvHcn6c1rhsD
PY6mTSRQTyDvZjgzfVHWU8R59bjc3HyQtCxSqt6j3CnBFH0N6XuizDxyM7jP3vCU
z8opTYUuiD79GL7xjzQWg7922zRumtxm22dke8pwREZyrzSTUKYCFa6vBmvdOHhQ
3IUqEFW3qBIWYkvISUJ2NUbu1huRNRvm2M6h5k9520zrXR6NbNeRgrFpBjuvi21n
DQBd9tvmvLc0ewR5DiQn4r28wh34ZeBKGpfFL0wcsgzGlGSIn1/vokm+CrY9ZUwK
Oa0txSNjG9AFpMv1xQfIcrC3unH/SpVeBpGotMUBRh2yGxUf1DLKvgsz3Tzr/Ojr
QI8bViLhU6KYf+bmAocNwVhd2HGuf7OoztE2grGQ9aK8oCxMRoGsHbPMGdkct347
wTB4+G1pjWyhvl2hpXyYrzt/cROVEMzf8G9X4rn05DjIwUEEcbyV9ThbMD+3UXra
dXUc7qTg2L+ORZk69QwR/rG63dL3Xzjp0SisQXbrzPXshQjHuUoWSaCx+PTt2yMP
V+6vUYM56fdZ+UbUMPgo2SJW8Sh9wBVC0bCFEHL20PQrlO+P818B0SMX9XjiLKO5
B+WyhK/jqr9o1KyrBahe92q8UFvMhv7VIQu3T1kBSkCSzbM1qPfaYz+Sxs0YFT66
ELvQz2FypvLAc+eZ3sx4p7U2iCevTdWZs/wqxeMyCw402P55U5vd8ZK9jo99h1Ay
eFo2iTVRNu0y2+AkHQNJdJeAp6UZ75sPO0VoYtdscYnHeaZjzqMCb1kJqYFelORa
vlRg9t94fsY3FzUhl2AkwQH5MCnWSwdNOozNPL1fXjVFYLpvTL2akiEuwRVlLKn5
tEC4FvwJN4MeZu6tRg4JdIZcV2o9ZOfdNEXCnJkaagxipy9uiUhMqW94BtOsHasj
VQOSPTwUnvW4hmn5H+AIPgs11/rJcblVLFt5fw94BxGItSNs4uTRprGubVsEVuFJ
1Gplw+cVOyZsezczAdNS2381Y/3l95ivDRYT/cEjOYDDUxL7oUnkC1FNAKOfWRM7
T2zVIXu1QnNgXhEHzGcbR8PCLMR+cgOAY0IvOtziLh2AL4WnS9vHzaWHsZJUnp0O
S3QW1td4YroCE/0ADQ2Aa0yRYyH3ZGW5BxIEsd3A0E2KauluVfh18aGnlDWbL/MC
UafBU9K9TOljBfqMxN5DLyFsghBIL5DGZbzCBh7fDmnr2unn1keYSPBGsCQmL5zh
Zn6n2d7BayZgdj6wYp40EqQeKsF+XueToFZq9XjEYjHLkjLi1wNG+X1nQPlksMaw
mtBalMNokUiBA6aicLd6TX4Xm3sX+JHGIGs/8fAJclBgcqrccQXFMcje6ZpMrSBn
DRixm4/gNp5Knzv040h/KKmo8WEKOh9cZ6BnzbXtIcpg6ZFYsxeyiHByBlEXm0Ur
RQQVdoURZTlL36T4qe1IJI65oCge7igJoHXm4P5eN3pXoiEgPlpVHDPlToOFRCUl
xRz8DjRwUIZ3IZmWF8vq1Bim6WajTQoFC57aBXVHUzxDLIFyRnBBR3N4au6UEO76
24RfhlqrlDwAjUH7/KONLvwxumSofHxoz4upHrYFg8Xmjs7vUBHnIX8SbXPo74Dv
igEVeJ8XwGkY6NDNRxgg6v+T6fHbSGdueo0zlZV8wWoiWV0IvBArKIPCJTOBhrnO
z8ab0FUah/AUP6IYI/srdRs8f2GiCYvegi64PHOu7zYJdGG6aVTllxAjGiACozZQ
p0Mbp68CqO9N2Q5Ruy9Db693G+GTMogfKgH0FEPSUQOkI+vfe2ewnrOD0JmvcZCE
fQwUh3e0RGi9zsnFDet57XPgvk0AIvpyatx0fjJmQdmxySMJimDiIMVf11WXe0EL
ARJ6HPHYbPq6Fzav0kR16SMfNSMoSSdMe8gyGvv2DUomlWnVuxZyjcwvvBy0BX11
aAsJFgm2dmi2+pdpEr6Nz2rasDD+RYOBEqgEhsIthwcl7aKEZF8APaZyN16lE11Y
+1LUAgGR74wWZn/ADH1nw0/X4GkIS8nYdMY9RD44cuqtgmzUZzlXYH9OfSS9Uk++
HmIDe4IWZ2kUWYq0VJEHt2U7IgIkWXqq8+NkNLToSKOGu/5d06iLxOq8DPFQheCN
I0md5bIwplAqUSyseT2WVG2SdyemKJ0/QBO5ZOJT0/E4sMF7oWHGHXYXSACV1HCg
hhP2kcYPvKFm59dEhgHqXry+KVx/oOoyOsD9mmW+DEnvUfKGfYDQ3+frmlLFGnt3
9ynkTkHBBCj9OYvcunE64Ue42P950ieyAl+NlzmzgmlCCU+ALQtgNvjOpxA1drwa
IaQLvACyyBGss4Awx9RVRaBy23SiZ7vH5dFRRb80e9wY9omGQAcSyKwkjRTHKNsl
Yc/2H8Kycf5ZGSI/y7VRnLu5O/U3ngKbGWDTtXB9r6XSaFcWT7U9hq7GPOPct6xJ
oStmUJy043XA8UXUU7tib8/1FGLzLm9R0kpbG+BWQ1fk05U/4xDl1PBF5bIzV5S6
HBShCEBtgxyBrpu6tGXe7UWx5wBlqYCDkt7i9VOCRjRRtIlvzy2GLxTrJ6cUdEAK
Tip/rfp5y4xXIqCNMM6rGaiewC8UKEti/l7dTlQRU4K8exRm/Z3XxXSzjwc+ePh9
jQaPWLDMiEPBkDJ9rw3SIv+xQ6uDHdGxwONMiSczF7hmIuYKcCcWUbn0FuY4Zq5D
+ZCetLuOwfWma9NClLWREmAJUcaJOXpcqgaT1XFQ4QGEy7vw4qViU1BxWimX27Jr
Vm1IMpH1+ou9WDHCzKdwcXNRA5lI+AZG5cJzHMJQqg+jT6pGov5ZECTPKG5M6FMu
0/Dw5cmiPVHomK1cAW0d8Bq0NUUbgpD27b56PtcyNl8c7VyC42rnMh1eOJqn4JXL
Cir5zVEp4k1f6jb7ZsyD3Ia5CTz8P1D8yfaojUFtkS77TT2xRWMNaXVSul18jnp2
4pFd8FhBjalP/uULDhQfYi6tNWlIc/BiBCLLqCb67H/F61/DWBMIY/FClwdrcDzn
BHRe6/iG+GPe035W3RZ2Lzl+8gitBPHWbdi9oTQc7vuY4Svm4cAdJ+yy8dKz4iKX
zrDYa82SMKV5HQjyw5elmWVI2Md3IehVV8/jrSBWdNrxHygjRvGYMebMLZDT4Kvg
/A4VyMx45Umzi9WEjBr5u2WG4DPG5yqrtRPFJ8EdQknHtg8erE+pgywr7I1I0kz+
1cvNyD50plAthHbpjJbozGibzeOSFW3LtcUVLbIe8Ea9uSujvP2XiPuCbT+41brs
4qifBUUF/xV/k9YjdL3yokOGFbcP2oytG/wvDMmc0dh8DvZl1ErtK9816E0Y5duO
mmdIOzxR8E6E8JUj0u221C6bpXAeW5jrivM62QolkDB1ZiP4rRj9QqrrioTpdxTP
o8twrzf3iyzMswMK6S5J76IzahNK+EVumW0C29+vUTuYDD4TZxPQ13sRBkX+dgU+
8cdNyQyfaNslto0RVfJ87de5ZO8WJf6N5/OtTSJB/5AF05Eg2ekH9o3fYY6dtBiW
qL+L9n/KIU8DX+YVDGOdeXlrwHQZF+Ct/XQCEVPO+a89qRtvSvyVxGQXtzq47xfk
buZBRligx0V6AZn9p6w6K04BHF7tn9QxSWc8AMb6WqGKPvWRwoSna20OShtQXCT6
1LW45YWs/RdDVnIEbA5/0doN7iGlXzU/I8dno0BV2ViibdpDhQKt+XjYXbWll+3L
/8vvf0zBI2hMHTTQ4tamgWyWJUFf6G6+fU72ydXq/OBmocYm0WYSeUJkr6TvDcb6
/xv6SwN7HH6phYD1nLcpSWVkWVLDqzFJ0fLgnSE5cEHVatvdFQhZAvNlfL/OAmt5
aiyM+WChroulJ5iHSONNG+Jmuro9Sxe/oVnFT09o6+FRUq6Ii5ChlTy8/pWdfeMO
ZKHjS+kYRT+ZuUcCjl4ismk1/jN6trfuGzudbYKvYNUoh3ImD2qTWEANcZzhhiaj
Y/GYcRZaOlz30PFLUqxdkDS1JZJL04qUwhapvFNDaJlt3oSm0yPa5Ic1P6Ox7hFg
/3u941dafJNHk02aF30znLxNeKtY8AVoMH/TLBz0ef/6vULkJxGDmWEo0W/mt4nr
FZWT23a/6H8w4AHTwGZInsxgk+Vdrpu1fUoXvGXl4QrLIhj6YShW8nS93d0c4kxb
nhS+lRhhAPIlkC0CC2zFbfdwxAos/QsA2xTDHbx8+Uguad2VtHl+8JK4iw84OhNV
3dwikrBux+Bha//GdgSHFJ4WjnRRQsgB8wH/g7/yWSTZtXAEUDvkuJtQvX+oQE69
qW+7gfs5mzHSdZTGg2tqcmOpIE07uo5OlXI1EUPJquoUVG9ul8d5JmCRoP9NILSZ
9ifweItUsB1y8KSGDfJlWIFayGYZmdhCA7deydVnpQcUrtGGAcZWuCZqRRdknTj8
SbKPq0buu45dBTk+Pty1FqAKEuyJpBN7yDkqFzo3dnXHBaJw4NrrSIpaFOrCcx5h
7b1gMqdoqssLXtl5GtM4LEQw96t9WnOVXmarUaggWmj4JfgU0sX1lhuRIPEV2SjG
fmLPBcdD9ZMhxS58gR5dkPFdFEgRnSMCL1qo0OXKPlpXkb9Nx3GtrvLalOpJhxcg
fLdLLqIvVm8t6dS4ik3Bx68X2y0NurrLoahxq7Gcdfti5WXIlxD+0JbikUVEFF0u
HhimCFqdm2XKLPk9acQ9QtX81jdjkhzYfXZNL5jFhv0az2jfQdIGYXiX86X1Vd23
zDmCFQPeg5D/6PoCSWm7JKCw+bPRxQDG8oxn4+MHs0xcCexVXjCdteqtSbh3iUl3
FGTr4CU0mwdtzvACy9oLICF/t3PjszQiBtyVdbCJdciR1cEuu3W6TRaQD6UpK6xF
jKGjjyqZZdCJbVij9OHouySmqo7UXOUASf8AQsBN5v6+n4Uebabezg7Aw535MKVY
NI0dhRXZZlTn0YHhtP3YWfQavqvgR8zf3NplI8ZdeXE7ZT43MxYwH9Wny3aQMy9v
Lmo9SskyKd5LwRQO30KlVtaqI0wjYT/zpPK/qdLYescLZHPCNyvb8GmB8RvfztNz
gixYQZwYYCPg9WMeBjgxiaR5/NXTIekGWlQNi5IAOAJiY9OVfKwpF/gx1XwO05PS
8HTJ+AsIYBzbGl3rukNgoX4FCh34j9i3Q3LrRb0jaykLLQgavt8slx/tfGwkgvyO
5Fa93Qwx9bg8h02ilP0XrrAGZMJ4GfmB4PHTsTnBr1JoTLDjra7S5CHVJ5yPJVoA
I/3EYDDzbvAiW4rzZVl07Lf8I2hBZikSyT1EwKMaEtlP8OnfkIBihMwSIFFSCNEV
+T4eB0zTNZEG3VCzw2q9n7zQA4bN4Fc1pwUrsi5NJKkMG+dMEeIFcp3DNLmblpAq
v0gctOu5lxc5leILEODY/jawFpDrsdNnVt36jOF+Q6tD99gViHt3j8YMGbsDAZrm
hgb5KDNCb9hU8Q+cFYf79HtacCVNQS4115gq7ErZ+kddP/bfd13uf3NYKJ7ZryS2
ykV13Tu/h0Uqso+6v10tc9cX+ihLGbOi48jPmjIaFHfWJheEwnZtglBHGLre+PqX
+GpMn4rEP00WJI/9gZoeBehix4+hOXV68OhcWd1hqvWy8WDnd57v44v3zRtlIIgJ
EyJrwzVvLso5hxhSoKS1C2JhxK4scmVH7tAVO0bB93QcTmC4Md9BHzZ7Fqf1mqU4
JIdwQ4wIjS5jNbATvj1IXK3SLTzGZwsRqIpGp7tA1L31jCn0e68rqODPqT1n5cIk
ZSSNkV6vYJz2ifMVbjhsAIJ/XtHFx3V3N9tNwISGaVW/4AKNlpx7H+ElyhrV7iel
xhaKAIW+weQ0CnYweTZdFKpvNiau2JkVrvmAw6WERnMPKt3woQvB3eErMPkIipMr
zfXHA5aNS7mAe/W4I7Wel9e9xzU43245TAXhmCYpwoZVu1adF0/8dErOObjjtBnE
StKYH5uAoQjY7406/hTXF8kWUJjH0w/Fz+kB53tLqmMZEH5rG8UqoFZC8h+BAEBI
YyFV2WQgoiAocBhTHhkPEDB7uK9XQ35awsfobJL4ZNF05qtcUZhF+v2+42r8hOkj
qxc6+D4YlM2MZccIVwFosJ+/TkSeDhecYs+/jp8i3JMNH07gDzRtX1E3uTnmp4U1
6ci8pBYo4/ssJ07ICAz+qCtcpCywNNBG3uCV801Ct8scFmFYp8d5TEfSJ8+SJXuy
egTM0aWtv1X43/1yEkJEYJvD37sq9AG+k+sFeZHI7h2WLYlpPflxtnM5KQ8FEC39
n4zX8+GG79+L6ta2j/sAvWljafP3LRSSzw2LHJ8IFJ5ZsR4IbdSd9PTagLuVPR2p
d3bp7za3aPCe9t/Qrjn15EA/AP05fcTsFM3mwP+vOX90GyDbGmuumay15DsvZHcI
07bVvq6jrvdpvvBZ0JClCXWJlMMhUlAg9aNvZ/FpJZCEspP5mda6dWbK0AW06Y0N
h77brbibINn3Qhjnr6c9KU8mq+p2N7PmeXnCOwPq2DQsgnuoalzaYFl+fIxCqxI9
4+6C1K8BYogL0XW8sh702jMFcJkV0nvv5bF0IQGlD8aVGlFfVJw+KfXnz9sQb1NK
r5cdiVxbw6jGEJSiaG2UGRv4hsXOnncW+g+8DQQxgGoy+ROXGnIZckIE3YD+LUGp
xIR07abBm1aezaRslb1leK4pyyAOFs6U0ViB6PM0W3GbHGQzQ/YddlyvHlw2G/KO
td68W3kDomqHwa3yIlWXzcjItW7IksDzt6ey52Grq/DFaa87UcacncphujjibJNi
CVssjuFo4Cw/pEzPjt+3YG5XVlm+/6y9NO+EWLeEv7ZWWvCrcKhrkgMqLlGaUOcW
fkUm1RB3H+sLrqhTxkCYSoqezcUthKj4KTJwwpxiwknhvkAg8n9NBBh53p4saqXb
2RNX7Z37wWdfVXcuh1fl6YGqEXH6j0DEEN8VmqoYA1wmJscrt2yGqifps8eiVjBs
AXZlkN6IDJ/A25Q5EFePy/5JnZ5KPSztb75hMfJfDq7jFvRST/xTcEr/KZxL5bsi
4Qzvugkjso4l3m8svFF/MkubvdRpcl6a7afU/wel3jMFb7m0T3RQlIo0UGGPTPJ+
IYKEJa7zaBpffRrqYpu/7KhtdoJ2IwUq2v8LYrbGs/q1Z8lUNIcMNlWZUML6jBmL
sKdW7M5FJQZPgrYe/Nfu6nv7wBibqawOxVDrpy4qb4a1G4w9lhWHK7bOXxZAw3Ca
+Zs1A1zWUoMIjXQtZtRzMeTBcT2wAu/WSOLropiB+D5+9YVDlTS4DxnJtTrybqIr
nvpQHMja3wSr4UmNGsWyGzfnnxeeCEsQnKywMMc09gi67LoW73epssKAaJx/Xl+O
Jfh7jb3Bkif1sKrgr5Z9KfNBBw1+IUfz2YbdAVCeQ0zEfaC8vswJVN/yrEXlTiXa
YiW//CyDkj6xlM4ClEhc8AXTdrUoIteF2DGsOi61dMlYqEj1RyRK50l4KBVWJxcK
j9T/0O9xY5RQZY3fKEgnyeg6k4POcnen5dPpwYw0sIpg6eGKFisPf3u8VHU84cLy
z+CZQRFxiwEhhCiKadeuGdaYtco+fhke06sNbkx2XbnU0WGR3FjykwN1s+YxtAkx
ES7q/oCjAOKbK4290jxKrRJOulKEQSjbUPPFRbqV/iI0O2AJCUN4zFXD24tinnCf
CsT+aJMBiPSE19dPWlIMlaqxWLNRtIgAJpCgtAaelsvhYiUAxM3aOQxgUQJswmQJ
O9tj0CW5Z0o9TGV0frKWvIZggZROJg6ndHhzNF2Cz8pbknOOVc4k8MM5tXDwE2qD
fawxD7hgfkybCw1Tc1KmzG9KOWvoKM544JV1d7EfwTliX0RyhpITzcJL4CUsail4
kKbvFRLQxDuVQlK8AGN8V3MgRpK+1a3aEytxzL3KeTBOdKQk5v5n2k2Av3CbeY8+
Xa0PEgIBsEG5HypV+Ftn7Rz9PSXZGOm9fC9RIZyDsGSncWOJDUI0TsjysATOe1f7
ucUm/uxV2BDiDGJKQWDSFkYsFTNWKCpHHQXKqokKtcf9gVOE8/yx5i4YyV0AXP7Z
5pvGmKmdBs5JjoWLUQD6fA6PaI8e/YuvgY2BlkxExCOAUCVq3qtEyhttMxBYr/bz
bINl4eYkeYRMoudysgWh8aEkwsKuH4eNAhNoy0ZZWFeFNgTq5LT4EbbF7Qk6MPnX
Grr0TKb2qj3JRpnlMHsvz8Oj7mITmgrYGwzCvHP9xPKNclxaBZguzbMtS0VXyoq7
g/YMXTLPJcvbYeC28+zJ1uNemirDfKxhbmTbY0YNXqIYxeCEVTzEWQehql683v5F
24Ua7KNw/RNsYnfPSpX7pxvzcOz20988xOnbn94yyLfTBqAN/AAM0CTGP8wA2Qiv
1oAzrCbSYcnrVes5td1ayIaWyP73yTfxpvYN5mdI/D3GegXonCir92AQrZJo6MRM
Tz3bciokLudblcer/uVVwKjiitXaQHCY6ZCI/UbDwuYXYIm3L7jihhW9ZBFUql0X
SzFvOeqSY/lYV+4z+Uqag1/Wo1lS/mmUU5k470bqum3wMUGvlzhFieJw9zzmOQ1m
6o68xIPPVVud4J1265gPsUJDo8QcQfXT5IwCbbs7yt1nIh9hWhdFzOs/9NEQQ5UP
NDc4gi2x1iEBz1BYTw/XjFFvkN0JLlK4OcXB3t7DOCJfJq/cHYz9Q8ZXGJ+wYhCi
t3RTB6kdYMKLrm2VlirFxGfayc+5LmX5LZ9Rjzv9MHmY860O5ODwwl3FG/AdIie2
rPEGN7NOqEiWBJ7COoAeCOijTA0RMFOFNTGbZ1M8zwZ4ZcuaALxM2Sj9rUIpC13O
YxpBntvnaJv3LTQG3a0go0W2i+6k7w/q+2KdEDGr1KY50GGJzKmGhpTDnKS1fL8G
a73PTPaDWHvtqQRvgTwr2tZTi/Q2BWWO23/+kNQVA1LUIwl7VRAPm34zei6tRT4v
t6xxJre3ufyn1am/CsNWgFV7BnlnEJhtNPe98j/rymyC3tj0ZGTRVGRDAkylPwRK
jYCDT6wi+SUf46eGSLOZA82NvsQ6sJH4oDrWnNxnVs9v870bpfT9gucOY56/ez9e
TbwkuqkRPbomAj/LArin5ug5pxr9FjoOBnDN0OKl83PMYoH6SDm/PhYZHdSfMkrc
OgnWTDACrL/uPTSSL7R6+I4kvR+Qt5BRGT33JOXhlp72Tq+6uaOg6voqWs7IEHcU
gPLH4eRbYzNGe4x3p1thAplL07Zcr0CkWvIfOSd1yVu9uQALHleysGd9d9P0mh5U
bheAZ3Q29C5BZzdeHiG9sm/ehcevyKi/TwIs37wrLKH6YVHl4/dYOFWqsXNvrYoL
sdnuBhI7DNCDkHOCywLmXQEHE8LErNPTBNi/QbsrPJTaGIUiOzlAdUHSh8XinGEM
3D9afF5tBzKFIoIYxShlQxVWOcVhZmP5K/w8+LJT37dhB0Z7rvkxwdGeXXE56sva
3plqNWJ6xP7BIgTqxpvvFr/5U/wisTOldB0B+Dp2IRycxNlWdSD+Mb6HT/ggyouY
1Ar4420BBauQP9c322imlMEB7HHdRWIfZ6MkQtkj4VkBHszjsqDFrCUb0je7oPtC
HW76kR0UwOVNfNkpP/aetAc4W5pt5yLdU2n/LY83mLs8fbqIjjw+nrNl00VkkIMv
qkFwaML6rzg1sCp9AaPspIzQtyrC6RoYX6Ku/5KwaUTe4m1pD3amTggvdxFvZQnn
g/dn9Rtge5z6rhMV0reDXqNmsYFak8oovz1k8ENTbuVPzBW7XdZdg4L6j/WjAnQI
TUmxUJK3bFLk4IthVungScbzlzvSmvBS2h361JwEZ0RqiSJwl5MakqerhJh5zXKb
+FfJTV75b0+8w+M0bPgZODpq07bdwjjj757+fJDq5TWh/4M4nTRdY/rdq7fbuIO3
bJfcuspGwmfblhtMiWwBloqMyX725zIGYtzO21t6LbI1wly34tfqPIgQhswZWJxh
tKx2n/1VuQInl7kJD3Kuey5MGdXl/mR8JS4ody952S7Cy9V1r8F6WCKR6U1ftfK2
XMbKF8qszYZSsmQSrbfEoYjwFnQenrdr1uraTXpXaZGhzdbSOStBSHoD8PQWWNOu
Qr1n6uGy7QyZ0UAL+q18LYxLQyrYFlS5mbNpDThe0lGWmtP0WGNkovTIDFzjp5sA
3TxjOLWV03gUBq8lUAtnj8NwOOXt9A5NonJMmARTYYFnw3YbM8gUnpIyzuAcPnAB
Gih9defBWgeK7rc9flApBzu1ZGkW4FOhpOmEp1YC3SqmJH+JUNMl+CLxl/DHeW+V
qGKYqXDqbF0ZkP99Fb8Ah/DsnxpUQ5Z0+inpusdlbDvcaITRoiVOblYAMFOQ3wnE
VJr4QNTs3bhTwiZem9EanHNeqWs8Q7FmIpVP8cb/N5SKnK6UbhsptveXoQ4gQX8X
rYVPzbLI4eR8tfgBvTxXW/lpCBh1IOZj82WGhpf1zO5MO05LOCnqvcEDc+lcRLSV
Nf7XRohyrLBPnzNqsl05Fei0xNhFcKIXDn8pGljpH29mgFmO0dTIwlWCqrAUfiCV
Z+fKktkn71B55Mny7T4mayELyK7i0SDYZsyxEIQnmXLHdwj2sd4lpEq2S4pasXyX
vypK7gB+1XQrh1FlKSnJJTIIwG2sJcgFP16v5Mhbpuu9NF9SSYYeUbw49J64BcY8
1gQUJfd0XcvwjWItRg+DugeQZQCtxqViCgZQRyo8Qd1IhFWa4Ta9kv4+eyU2OI9A
ymSkdliJISfjDxSZF667NBI7TTNvd2OCLjDzW0LEeMzt/Os6KnQCoGW2d7WByoiU
W9DxgZfkNRoifPUPM6p8jyYxVVi4+CxABS65YzCJLe/Ew3eB5BlbIOkDs5Dh3c34
vApTWHveyGGs9jKeaqQ7w/Lory3xaO5XCnk6o72QG/xufugz9pgcUKeWVd++qPTE
xyzpeXDhxTdJQCRoS+ydGHfmIJFcT8SF294PVddwgKtF4k/PZ7FDk3Kuefp4Bntf
xb2hPksQm2S7B+bhSBSj/Fb8bNLAu831LDmetxDf3MlEdN2RixHNxPUBfvEzBMOQ
LsWOBnQrDbB4qQ2n7AsckCV7y0EEqDB6OdvUemAPQQLYpzD8/WOtsqDri7hi1xsZ
NHgmJKvZ2YHoytmaZzqZomxfrgtOtGaaPai1CbE8oxtp0tmZ0HdNWDixZp2V3Z2h
FXE+J+Wk7M3Cz9ob1ggLPBbinTS3mh4Wl9tQDstbaclhNBiHnap5lTxzJgvgO1Ij
VEDa/KqdUIaFXz3p+Sf6cdg7an2oKFIrbOwnY4mduHskD6OeEyMawj3vYz6AiUkd
Yq5cdYNw+bXNJXnxcDTCS0wE+EOb9W4Xc2ETgiM3dinTZuP7zKVBqTD6AtgzYihF
Up8sr2+y2BLKvcNmXRAVaBC0PecM+ss+6d7VDBeTVmdeIb/YJpQwHQsl9L+5+CEb
LEWvoh1qPeKcaMdl+qiMwSgW4d0zBp+ysSV3MFQE+r+lzHN1OOrCHcbABnumMQDT
cX2R5EC8Zhh7bDwpmrW8C/xNt3jnl6lhIkinb5pTGUHLvuuRcUSiTlT+3by42XWK
IgTgWjmTLvsth29ogQmUgSs+cpJPaiqQU9YZbHQSfDaXawqHthuTEcH/7mA74wke
d65wuQx3qpWtOA6xX8k+2tGH3U59JHJfB52/rqNaJxX45n7jvmw87INmx4NpjXP7
8Z9FA5u7oVHg4osJqTAO9E1+a0YqVcl082v4B1yWJRCKmZBbe03WRPNinwZVV3wG
ShLWzqgaXe7iQ5Hc00fBzpiI4bo/R95tsC092npRoNLol404qL224ULjUNusWdJI
0CzjPsFl6K386isg9CjXANNSvOaykh9X/HQ397hjDwns1rHnfydMXr/+7rel4TBI
M5QQYtK4bSxAqZZae1x0yHvqOpBG+OkbAVB2NN1sUKSKKxYU6AnUbdycPGu1esno
4SBdb2pgXEnjeS0wcPxI9I1c8TdwJcv7fWcAfwIsEpoVgsSxfR15/9n3nnb6Js+A
3VPm4gUOhobKabJwnAI6lysV5KjhVO3Pn6TjQhPYiRkjpXPa1l7xxNzxB0Vmto5D
YDmlLFJajYD1Aez9cYOSZdFhmFvCqVNKTZGS8YlCcbJGXlnraixB+Pom89Lq7Rg3
8crKnwj7QvhkgoojN4vQ4haTlYRlwlURYIu4x1dDv5LvCmpcCjD/MzyYOduuwIpf
VC6a6nC9QEJQpsvXVr9J+2AEK7GgysfYE223T8bAAa4lcz1dMDKacfXggoyxLz7r
T/mK4KAOoPm4rmAaZNRKMRnIuTs/zMu0IcBrK+a26f1bJAGjccnggpVPVQJpaNDU
CAiahsw1oIS22YOkHKTu/V7QLlpeB80Bp1diL5krJioxwGyrf1z+w21SuOjeS0t7
XUfOgCd7c1uhPix0XvLA50AA+v35jIC0NhrCcOdpe0Iq7oSk9Fdh0c+r+7Xwejg7
jQJWDM95Rsks7zpRviDIRPrVFtPzMVwKkgtCI76GxmSHWFk3sbPnLWOxcrt7eqfn
0U9VMBlz9mHfKjlPigFUdVXB6nhipFU4/xGVIM178mQj9OxJA2e3N50Eksp9hw/y
UNCFigbXJvNjFT5kwEPNPWlFZAiH7FEIPuIyIQkqSX3p5l/FZzp9p9dP8JGxQcId
egnSPDRfvl1dxXLyK9CA2v+R0IMY5nJg7EReEI5xSQ/s+TLeeePsi1iWvwWDtgzF
DBfwcAJw8ymgCeyMUFkuRPGauhr4cbqqwSCOWPlUtRLHn6ZJGgJ58tw7dzSlnjfO
805U9JKGs7857T/Tf3LsM+JKoxeOqZNP/+WY+yNvZP+8eFqeuy7bQsTBSzzlcBva
qGK6JhuDSQgbfZAMBPYzNnYaaUM/+Dgz7a7w5+MSQ7Mjjt/A1TV6oLg76R1jDCPd
QSBBHogbBKKCm56Lry3dSentilAOXn5ABrFFkGIZoMxH1+HeQfoRWYzHhnMHWXlO
SgQPKng+qcN+ffW0pco7k+QYH3hs7xQ7mOiA9G1mkJk2ZxtjJAsSzCKO8vRIuPol
KI3Fcogv0jF9/itNimyxNaAevw7KIJQOWuUtLcrUcaSn0tzueXV+EWgiWqfSLdKX
FM0sTTDSvd+5r6q9MwXP4QIkDFoBUcJBM2Lb6wdi+1iCRbHbl1puwPhoxKwkjS8v
Xr80V0abzludi+1pXkAI+BP5R3Los68N56ZAgCFbcFP7N/xQDe+cTU+va5QZOxW1
Sm9xEvB9etDP7hsXt2Wi+QIvVxJ2tU24+1yj0ruG1FP6tCdkMqSoUBWiMgoUe9U9
tJZAOd7SwuC3StIxUUGVYrDi5CTN4qw0TSkw8ceQ0AlhQqee35oGA234suq6Oo3a
fDrdYqJymjU3HfWJI+dlGBxcmJShQ4LhU4HX2QARN8bw6jGnjp2CVOiG/0wfXA3M
P5gTgKq+/Yz5yqyzu+B72bObyqmiKI9VJR9h1ssyv/peO2CMT1Zh4uh/MEaeq13l
fX8CsY5wMJxL3VwJFTrxcRtNwNSYKrq7/VhIC7giVTxszKratx405IA6ZakKWTDo
pySVwlMl4IOQs4d1dhEomwmcyETpopM9jgXNWwNiz1LNCLJUa24HJAwEif6QgejX
3nibmUbQBLxqSaWtPLG94BN+hJrG11c48i09h2bANSEDK8I+mwObrQ0fDDk6E8hD
YyLsHECQ/q0qo3UvjlPljsF4h9HcN2VFXPMUnUMrkUJn+qLm8AyWGBwJ9SmgZYnG
EoYnXvclJKL35W50me4B6TnXL1VcJ99tJy/cnJ5p/6YCto+8aFIFKDOSkADU93Ov
EsB/Y3ZjwYNvA1/eKKUFGwFF4qJRlNV9OurOI9bVnLzKlJja3T/n3+OldkkIqtd3
jUE0WtJ3sSkl2moSR+Rj6l8skwEf0iK9yASm5s030iDmkhtTS73OEtlLL9V0jfLs
2YTeMaL6pnyUQrlqcC+KGSd3SpZaFexpKJneEIIRvHKaJ+GLZYM947CKkYkD05QN
UPieOVBwMQVHJcKAXRnbzTHoejAq54LC70gDHngJpgIZdR/ZICNTDBYeibekyAde
QDqsmStSmk9GUEJvmjeVPA+0CYANBFoRvg+jZ48GbT7gHfAqhUM7Z4YpPms0OuiN
psiOCt+jfgVVF4R183/SQwe/RvM8Ea1HTLSckEOJNYxDnkoa8tB19pqT7lfmC7FL
lEvl4Mb6k2UbtiN0DyI9N9+/KZmqVk6LYkX1/GxuMAD7YS+0Nke2zl6OFAzdIPja
kYJOG/IMf+wt/DDqskVQeZEKTsRvDbBEL/uArMVX0KFWF2SCNKQPT1ejfyTGyNWh
dX+rMHOuTz9wBAmJ7xpgLioHCEVIXk7lQuZW73GHhVOxKKM6m+TI/aUFZFqlQBvg
RkhaF1A9vyCf8s52VXXU83119rMTdMqXLkY/vla+YdaZSV6M9VKyCzQJ2qvzySnx
GM+4MKRxjsxcA754UM/Gb+Gn6GKGTbFJs9iLr/5J50slVHgN6b9FkZqNyJXggAsd
NlbjA1yhWv5jlVjiV6ZS5D8YBFwlR4AtzCBluO4Wxe3rpzo0G1ZQCmGOd1P2f14t
fvNdyvMkpMtSRP6/N1YHGawbt+artULMd8qUJVvBxehToJ2ofV/hojBApMTeQxnR
DTRSSMp/NMQsZiARfMAQRIWScPF+x9uGxeVul2/nbXvGlr9LxFLCRMVcONGrARvZ
2c0PJ46nB7SGlsyRhGgv7xN8Hyvg3J72A/iDlpxFe15HIyMONFqykCeIdOUaBJ/i
NJKdpIEKnGDU+bcLDwp7yR8ggVZWcfSZXoOGqYb0VXiFlKrIjXEMTMIQx5jHeMD1
iJ1ylv5qRp/fklvq4T2SnQKsffRb7IprFtwe/5WoseBFSD3b46bVqBIn3ku4iOjn
H+iakNPO28Awu4ncKPDhiO8dfmAKe4eIx8t6N5hQGznuRZamn4UOUYaBOvY9ZLtt
WmOnuEfC3aSbf4zB/AVkgc0fb3XhB7z3GBzDAEnBl3ZU05oCbMkOL3ieMqAYE4f6
A+5WOIsusAGkbEBXFww6QTLDEPPebAgAug3k2clILu3KT8pJFpuAw1F5prgLIpaB
5amPcYtS5YPuTU8PynxvAvSwCo+QgotJjHs3iKMIn0ZR47XOVt+Cn3JWtXXBguUT
tE8/FATNiRrLJA7S04xwwxiUE2F5NeZ/2TjNyRpkMfxglfaBEwI0wIgL5DB5LaWI
BU4Q68bip9lrlUdT+P0YKa56fp52h3DT4w6hwB0BF4moENCD70Gj1jDnHRVM8swW
v2s9BKoBCzH/31uw7QOT2uFxyg5LrVYL8uQLKVUBfejc+IbA1XR0NpRp6EEtA6fN
3YaBGx93SFMNpafBr5tuHQUfP4ceeZ9Y6s0gztvDMXfSgLj/gYcNBEP82l3LTkXg
LfWEgfe7phSOctmf0pZYfotqXtiD7AYTiR5eOqCZ3TvKOqbb6KtT08/O6chh864R
6c6H7/z3na/VDwrJEMnbKw5RGdYsbJ4G6aN/22sl0IPpO/64xXipKDdf3lQVa/Ay
eHbRUSO17S8DyHO6ZAvrNNC7lCB5LCtQtM7H2bdxlXOfLxGh2AfObLQXaVuQDjVW
F1u2XseJ7+ctC/iFqE8sUCzKiSz999Fweu7bz39k95K37QmFMOXQUA8Z9NlMem7J
ZvwX20VjLsZHQIaeey9+qte/c4+fnYF9eRmus12IwWdyNY30MO918azUbxKMkiY7
qY4p6Cpe3SQUqgBDM3MzBYblwxdqqDpokkWlsuPO/Msk5myY8wO8ewaRhSMcaPuB
Cq4w6yVHpjaeEEwQvoElVqceqrr/3V/LO5m8h/juiLfJyYzla58k+b3lZGwBrGlq
1iwDO1ABPuDE1fnqBGsPaiczbgomQkdhjFDZjv5bb/mGyU8ExCKhgRTKQ88FxkFp
KXoBbevKAk/2B/Swx/r9g2g4O9x6BNDsTPnw2bAaZFPz8InIukKUdTpsdUf96D7Q
cbu7MlrcPhAPs1qLaRhAtRsQv0V26MPMtFzc0bo/VkB9gG08vxVsUmRvpuB26EQF
V5rq809lbn1Fr220WG7EcxYe/r3psu9dTHf6dKRjzq8+7i2ht+Mg+xIaoh7CVMQp
O8KHwtV1+mAT/7kgfn1Bqsu0UljVbbVAx/3M3yKPm1F0ZdPzzNId28p4rXh21/Qs
PrQY5vWFARk3gyGF94VHpJjDClZvFmBSFlPOKJFtII6Vltiqp169Oe5oneJgc0E3
Am72Ow5lx2rHESVt3VL0AdKaUX1IiVBDGLY8ED6tYV31kxx0Sa/1/ri31E0VZYuI
3Tzl/XW6YGyjpDnaXZN7iTEjiR1GRbzwG3JRjhcw4jtR3Zu/eoX2Q6V0Ll+ZTYfF
xQEbXITuAQgmyfyDmy3f7NIaT0jlK5gbtBzY4bweqCKLyQYbiJ7pob1OzLwW/AHR
Alc6VYEI4u4ArSbUo3NPDbJ9tvpOIX/gJ9tLiiMz2XaPC7HinZ3lsPPTy8Y9y1sQ
/Z2aNL1qwyVoqJSCiN/lryAPyFejoMgc9CsKQX50ibtnjr+kPojHb0qD1zW/RCT1
XT+/CsdrpZ4HkX86hCL5lMPmvdyg6ib/80RohrzWWNkzwvsT+7ERqpsRSpNHNmxX
rxL+b7tvOAKJag9D+w5xxbEPeta/EDhNXRUce0MTIyJnsOv+jbxS1sJ8h1uI8Bp4
xmoy7ccakkwDzyvrmi+sFqG3Mj1DPAJL42fAnyDHRAI/y4MPsylmRPKPXdRXlLWj
miHYCdLV8g9vK08zUwsNBlYjKDeywSdb4aLQzycH33/ZkLeo9UsW452eau57P9X7
KEogzXWKZM3uVJhBAIWKehz/W3hwnf2rlTZrWtkk8rjad+oz9ygjrbGJgyhcrNtX
53ksG+T3Rbgt03QQo1VM9sSKuSzzkqTPBw7c1TeSITBzFtPmYOUJeJzpRwMXqS7e
RxCStI6mNGeOkrlhB+XjEAhPLWnixUbV2ktoiqPTCMBXTxiLD5YMd86gGzo3fZED
E9yWWamzNcdnTfB2XJMd/hEZVPx72CTs7hJtk05SzOHV9nvfZYJGHuz6CmNU8HfP
R9eSAvl8EkWy5EqT523bhKHB0kYhiBLPcFLmswc1t64u1QRRNbidaI0K1mXnkHp2
uI/0P9nIOvT8DOHE9ZmC+KfUJFuJVYrPyE6Zd5SzLechgOAWgQ3f/uN8t7H5WkpP
s5cshApfiHbe++V0fIuc/y1gMaxhIc0jXqbD5Q+inLskDgc2XrIn1K5UdNDqfLnC
f7oGFz+WHkSmwctVA05UfVdKPyd5w/kkwWtGPBi8eyT8UGvi0ZPise3jhtnEpErh
9M/tVURMQgHhwLH6zsba71mA6S/e+kLbnCbs2w71NHFn4VEBOM4QW8QbzFqMP7Bn
vBVnzUgUqnADWE1HIdFTymuln2IeZirl7LvYCdPL9ZaJpb27WUqCe8IyDjl6iFG2
EFbgUQ67az1WqJybI2dpSfgpIOP9SAyc/IZ7JBmeork7cF9DXwIIOwApdVS+HaKl
Y7uM2bVYUgFFAB27QnJ7ANlOu8cV+AF+eiwoV+QdyDRKV7J0UbUvSurxvbvGZlVT
GuzEzdo7S2kbTlC38ooTXveUjvvwKsNlizqLuh5thziKOVWAilUAyFY2la1aXncv
ow5wfke7XVKKPqGZJGolX29r55+Xu//+gL4M1fV2azTz6b+fjjZ0KeyefvMA9BMW
e45/KOS01/emylvBO5mQUlVHf1IVBVD9k8Zb86mlkO6Mc5lNajdsrGXM9jFKh8W1
VU+WPn/CoDmrIjIfIv4WxUBSBS0vogr/UT5Xz1BelszwmJhKoa9vfckbOGr4k6Nl
2RTeA1Am36wzLlc2TzJjSlL1LtOZc4GIorU+BkvyVvzCzqIeONGAIX7T9AvcBDac
xt5YVPW2Z2c+Y75VQwGi87bQtIP0nv8ikuqXZwPm3XjIIDU+NTa2HtEf0dN+cteW
ObmrF8SqTzMz4stOnN0aloByqwxG5HpoSW4546H0vtB3tU6lms4d97JtH5qQOY0d
Xz1oANUleO/71lLwy4EYtvHStU9iJYp1xepDVY+xLw0BFqKyWtZuxG4bECiZT3wL
MCJobVQyFPl5nlTh0+17oYQ8Df+Yu8h55eVUi60n4C1Z8wgjIKvJoooTyeRstVNS
vv+FfXsHR5RHD/bZpS1RKZ/mBFGaosb6UwgKKM3c+vxaByCOv9FTtj2A2dOLxweE
go13TZpv/tTRX3iQ3EDhyYGF6sQWZYUjR7PXJ/YlRWKBISuyZV3XLVwmHvUcOFgN
Tv8OAbWMsJxgibvdmucGFiE39MfKHVrQmq3vToN0dwudvJR5r4wNoQCRp9WYxOBv
Is/vJUejVus4Fzzf9vH6YSVbur9tyPRAS/fVc/7NeMRM/XJa6sOWJclbqJKmvUDA
1ANOYTsjjJHCFzsmfeLyl0TAJod5k3kkB2ow5In0H9V7XtfFmdSAk9vlS53F4LFf
Ub45NpzUUghyN99Y1IBy0SGQ/l6xFyu8IeacCA2HBHYiFGsKqPLhmJybEWqH/as+
TJtM+T7Y0DWshHrTkX2OrA4cgufZUvsevNv9HaqWhHeKBzmsSgop+TIZBKlUKi0R
65LYQAgc+ZX4ONFZw4rDxNKs0RJ5NWHnjy9y5RafmjAZONgqmBfPheHIImE0+8Kg
8Iofx06K+JiMd9m/EKFf3ue3fhpTqxwmsKaT3lPjB8yW/plo9+mBZpsuyFqgmoIx
iXK2PmGTmzfa+y93OixX9Xr+vlkM4EWOiT8yB0Nvec+MsyHvc6o3QWTFjN2WEaG7
UEUd4r9xvUfl11NyOYw/vq5CkPblYReBNu0fodo4lXou5PsdO56svhXCjAxZUP4U
y495A7Gf5VAMj63DYpn/lNh+cEE9nSithuZqD8dW9b4Y5OsHRbl5hi/c34D5hOC5
9sEeu6wJZrewVTTJ2qJ6gP5D05rmYhr+YvgSdtX15zQRVjSqhrNAf2o+wUYivovo
pfAanY38RpDNipQjhVfZTCkoC5HBZDf5/8wCCPS2JdzFuFmH5/4T+TFsbMcqvnd2
jfxKoY9LISoqHo5WR08YKVp1DT/iMw8ciFV78s3mvha6kGBeVUjY7viAZrK8+flD
Fl/C0AnPIOQuYs+dy+cCGE4iHr9Te7FdDgxZTw3s2O+W0pjE4uD83oH8lvZzeQSG
+vn1TltWnbjw8wNooKPwCimAREgk/OdMx+BfEmM0wlwaHhaiXf3K6uOQdpfyypks
IJb58UVlo1NggS8gx1eHLWTIm/lIXM5il5hNpN/j3cHSnFJU+kd/Ldq/Is4OJsai
oNmHKfIQnIhKC7NucbmVDqC8VeqJR6/rSzkCLilVIj2lrSh6e48LJK1DwhUrQZDE
1HbbDZUJCVKvxRcwIRoll6m84Dfn9pZ40VKwMGhCaB2Z9DHS+CC9O8ooxICAIOIA
S2Jq6qc2NsO0WvluwBnEiYDE/zo4Z6NgSNAz6toTVwNfTa3q2llDo5w8VOxQdfpw
iHvUD1Sano5QHXtQD3/vm+x9AZlGaXo0qtsIEDojz6cxAd/JBi4Vphhy1uwl+PFm
ncnGI3/5+EKc4EO5VffORdt9cvGnX3xwf3Ua8w+JgAMFlVgEBdwSCbp7X3vRtjFC
G/NG9BzspRdDdIprCYQdpZ6+0mN/sGTIoH0Y9TPKpraQ7YR0u9uESC7cNeE+03b4
PJLmmN9GarL2Wzwoq+BdJjcq/Q9Ol3W9ZBOcb0/4cFudnJBxvbL9WsaVs7qOznmQ
icOSMC275VMAIicAD+ZrZF/yWXDmpHxQhPY9/1AN0EzVsLVeyY5V28dIlNoWok6F
S5paEBGJc4nBcwOEHgQpo7goSATNksAYK8123faDwzg20EPWC0ge7QwMSHxyWQOC
npI3LOuD3xgmRFAmW4ScS529rtlp90oHYWcDhkRQyuHMeIj/r5j5zg8DxjQRAWNI
KqkzPpS/d2kGX8fnwzyd7MzUwTGhrFs18v71N/NqWWydrmbLSlwAa0ckD38/r+Ce
DwfA5w3/s2Yd4g1uR2nYeMHhWjZXCKIaX90rafC1QQiRciHn1+9GKBRj8IEF9IXF
A1ZD7ldtKzOLmfu528A0w+ELRQrohYPz4/AktPTntDHfHyu4sJCmxON+2SI32bbd
uKEKgXdj+GBRqWvv4sa4SxojwlvLztzd4FMLSJjgInXowYXME5jkEFkk31HaBLBl
NC6p/rhKL4oZBGoaxTlIBb6mpmZeitWJAzjeJX8iQaZJKsy9ZXCiOdbbmgEPGOU7
Rg68UirJi/JyPBuG4iiB5CwSAhvjqDxxK2yVxJMlykat5U3WIA22n7u7GTmCVeWu
9lWjwbeB+O0DL86VVeOwRqWm6ZWfR884bNiQaRuzJBINqWceyxNplTULWB2faBgJ
sC5JGYFM7lRFraN0SysPdIkaBDi3bhdDkhsqZi6dmYJ8tul7A5CM/sHs8kERmPxF
Dv7fitXk2y2FmRNgI2Ki0zD/qoeQf5t/XR8NSjSmlDYhtyjiXZWmA5hCKLKk+SH7
EaNwKxslVzr7pyuPIcnvewcsOtjdWQb6P9G2MHdFlRtcCGEn+YWzbdJR0MCR8YXK
aHb7RTF57CWzx3bNlydv3hAJ9uvNdUefQWSwwkPr+0ircNbVjSZ/GfbPUFgQJ2NU
6i6EvdRsZBt5WGOmibEDTZLOtMIjEdhtpmCg7EgDgcokEMzhK5euyf+eyw66xAG+
v43EqAv9M2jkKN1TL3Te6xdfxpd9h5giCVNHBGd/lf54T+0QG0+U891rDPiO/bNL
C+LWi7aS53z9TPM3ntU6HQvYqREzy/HzzXleCaw2udPIzI0PkfzLVFJThcr8Leps
LBvuNxPQ/d1ldHnQwKK8OQrAZ3byDwa3p5DRm8T05o2WWwGSs+7Cyg3T7EY/JTBq
gqEn9H6Ar3ExkSjEWdKO886dfZOoIU0/x7jFc8IKwjojyYtUwiALaBe+Dr182DP0
rdXf1YFgdwKzE+H2ydVlNqm6oZPqexV05ttts6SexfiFqRyBlgrkahDV8an+Qhyg
R5exPg3nJ1leGYXOT16pBuF+6HSNEyX/ira2vv24NeGOBF+9vfhSMAsBg1Y8LOra
S+f5O+QAyWxestf4l8KnP1f/ovz58KwHO+ZjDuT7IUGgZnDWq1gb8oVSxA7vAI8G
IcDQliuQ9zHqX6Zs96wajzY7QIJo5Y6n8mEz7lSn1J/B6SBKFW/aiOCcwDJkzc9w
6oCCAP4Lul/P6LxKDGnuzr2igXefo8uGcdpkQ7J7aCANwRovTrsHDs3Nbsd6qsoe
edqfxh+rI0RHdCpQ62T1Zsv6r1b558vmrPOFWJ6vPWPxpg00J999zbBt2aG7CyTn
Uec8q3VsvtYpYmDkA7RURiZvDH7b0hGQHcd+3NiUzjaaat87AQKireDAVpciKHy+
aADHEr8EBs4h1TIYv0EE8RBtUdZ43vsMREpOJ18LxcRDHZlWJtXixLDjfENLdKKg
kQII/ikR74krh1+6KYslfyy8KZbKk86qX/KlI+jTd9apEEV7XY38FqMGeyfZsVFd
Gps0ua0MCBoS/hDBheP73rEAmnqVN5wm6EeehtJcyrDSO1Hnx/gVdG7dTdpP0xzg
HWw9AHDH2uxKm1USKvfwho0btjRyPOPcyHxB+hzuyWpfbAUi59M2/McXAvh7Vn4W
rigndX9pV2bGWrluzDQ09eTpVFZSwvnBxI24PCQZOzxPIkJ+YdVwgvX0WiSK64CZ
trjcrRUTIswyIc/94ANH26rjNzXeM6PbcXXjKZ43eFzT20kP1J8INbS4PjpHFKyu
4jt/vgYLDSPG4QQua157VR+YtLHS/i1RHLf7WyIu7oAPi/wxk6kWYOr7aEbwH5XJ
khgkiLk/CDtVEu8OvC2K85hYDZcX2DoReBAtB3liDU/4naJsgpCq9gheePrhSudO
mcnGF1RKcd42FbOXGboVXOpOgn3C5yDB25OYDJs/XYay4ReIn2/l+Xthp+GbKqNe
etXlMySuh4FgSQ8ufge6co9mIIEvQm2tdpjAgQ2JMlmPKMCpIWUxhK1uZngPKuPd
e0G9qkysQe4/PnNswtRN9Sp+ep6w9MFLLfNOsK2ynPCLEd1S89/T4Y34ja1ItOUT
F6cSyFsg+Kj+t8qwx0fNvevEC3TRsO5T5MKaEVbn8b2yEvubHJ5ZhB68O3q+ohNp
Zh03yNmdifTCCmijTdOPsCwh3ieeX9a+xpzscNl5HLqVta387bVzFXUvOWDxFCE/
skYVPg2HhzVsjiucJVbKr6V487xOHB1Ke3XJ5QYzA19GSODPljr1vishz4C7uI33
bN5aop+HG2F1FizCtb8bzjuNNO/TIzdIuZrVv3ZUymHvtQhBDf1tqk6PD33Gbk4/
iiW+NEwFwY9wQbmgJ1MmsyahWK07Siugy4CfcvGc8i3wFMh64ql/X1fYxZW95XdY
3DQOyrSbomnLiXKflicPTnnJw9VDUB1pY2uZj7mbHqNTPhl4vyD1q53ziK36vUli
YDpKNivWDVqEG9KWUAtzGGH1rKlEzfTLfWnbiG0zJ3yzrgWNn5SqVMlnl51qb03P
SLcakO/9JR/H/nn0aUeaGmfrzfH3DyQjAhP+kjrtzTDC9taZHW2W5CwToQDKJ8kr
msK0zeUbR+9E/QIMB64vz0q9o3tfl8kYwfeHQkTXn45k02J8iYrzZazWICP2b9mo
dkmGGbWmKtJcd/35noakXGxtxu+I5fQPgk8V2F0fbvrPnDdqqH88KTKVon0TuSd0
6/Ym8zWJ4SgqCiHh5p67V7jlC8BXSveG8M1ydzwITmu7SI1mRWCed/FTlIlK5exh
IwGJ1UaQhyxu1EkWjP5pKpKqry4AAF8bgtnw708Z2pOv+PblfjAWC2gwtSMlzqBn
Sf6/ST6h8kPU0M/IAbsK6wt5w4TmjQJJ6iuaZzpeYXF7E/uM+GofGEamtK/7JNpf
uQ52YMLxrv0bpAHNxQY+nTIA+D8grz1t50CxNojrLpDivKWnHB/1cb9R+C6ck4IL
77vX+j2ssTfOuW4F+EynJLdvIAvcLUTSlXgOF2Zk/7SL0jt37+RJPTFVH7ubTsQa
zhG009SjLEjNdaGFY+SbOVnktG09kgPJJSVgoeGSez/q4rTHOejA45ysuSEqIz5d
Cy7yuoDUa9joDudW7km/Jkn3EvsSwGd0biQCIpzmRpJkDGLCX2KOIAXr/Hw8+AQm
u2/mSuMFvvDW0BOcDwQcXSAq4rv7EqbFNiI9jjA80yIQIMYOSOiPmLUiSWK7gmK5
LDB5E2aNP2ns4lFk+masZFtl6lEJJ4ZaXVDWSEqyckUiYgVLHiSmiDX8pKD21eB0
uE9DIq1STU8SRrwYzyJJd7YNzf308Zs+38AGWqoTEqPXnmBq0/67pC0T2Lk4mJ7L
IDLRfxUB1MbnGc5s/oaYs6IxDFxUxCcpO07tqieBHHoPhdoGft1zsNs8M0szyo/B
W7AGurchuIg9Kjd6hZX8rYNxkvjWa5S5nXfhHUlCQbkkootLSIo0LNF1j/4+MnpV
VniHaW1d4JhRasU3MXSIXLEUUgDGhmN2gOS5UOJ0sczIiLUhLjfHuVRjycF6U6Tb
ojw2duMHswrIb3EeYxw7BipaL5KIycbb5rEtCg6An6TLuVdx9XsmeHtuQrEJPaMr
D05v9geH5xfmhmN86X32KIV7lUpYqLTAE0AMVXECVIipWGLig16tnNi/Vmb8Di4R
ESu4/o756b5kLWeqZm5kE7xY3dS+jjcyWBm2I05ecD0W95iVoByQXHqn28GN4cGO
I1FB4uLWQLPzD2fk6wbLJ1Jyh9rJsLEjMa3Lod7C5+8gsPWn0t8fCdmEM24zAzOn
qZRPXOPwTUuPQc1l2njjtxKmmn/FJOF1tk/a7vluy70B0h/jIvIOR5YaR7PNZ8Jy
W/5hiyhb1PYbG9UIUiXcBDvnp2GHZmZ/W9VvsakOgnhYfCh2EmHiCAfIJwDoZw9d
e0wAufxaLRboE0QdRNqSC9vCa4VgHrrUvdHVrCqFSqSVeNDcuAQhAYl6cAGoBtm0
bC6wq8dVxwfgzF3Ctg3OQhDt+Jl0f4ltXfuj2TJVlepHzgFUlI59elD2tPTvRj3A
jzxNBtOoyr/id/OvLezhSkPcDNbdOD+ibH9RfSGjZHQJ5wGRrtKdvDzAn9yFUY1f
9SE4OvT97TpfyX/2dTBdy82vPGoQGVEoY4B/Z0E3cixPu9bqobqqn88PKIgFdvoe
LQdrx4kVZR0Cj7ziaqyv6+lp0TPR1iIdHwVeMpZ51YmmbZIBZreCUjAH32iwUMtL
l86XIpaASwerEM5oJjtEC26zxbT1UQxLPbaIUodHomGH4GTR+7XLrHtsQ4k4/deQ
78ls2fLwuQsLsWhVXqBby8m2r22oiYGkts3cNPcFAnjHlABeSE4R3ez/IOx7//Kz
S6oWVwm5u+0Xtls8DtXW4+9ujBmHvWa9dpmqRsAzPH7EkWApNLWC2N9S5FKsTjwh
I8hMxgdvP6k4bLiIvX0M8VDcvkbLmmNARgZ0raqgV+rDewMs3MvrkyPvMDkF7l1a
+t5xx4pAfiVxDirXClOn33Zcepxd8ToQ3IxFD86eNOUtwtr8l6WxQ2xT63BBB9So
ZoBVhdObubXqR2ymsP0lWX7TdgCwoRUCm3cpgcRHlTH2QZyJAn73/c1hcEwukru5
j5VkQ2AKkX+2PprIP789f1H8Im4Mop/ZoWVPvP2mNUbjN9BOODSyH4eW6gfHrihZ
V4xKQXgUfV1Yf3bCjWWj7xpCw5sFXWyf331mEFX30U+4AkQRd7RS925uWj9O5ZGS
WSq5tiw+ba8EaIiOcfu4qEkAwQphQPNlhgtySoONJV4571trdHsumU8PIB722d92
EJ8M4/j/gg7+VpJ0Rgu7Ey/oTqO8WRO5F2au0L4GHPGwrlNrd+oIBgAUrR6HM5R6
6LO30DJnoXbNnAE3UDiUGQPvuRitLYtPeVAaAM5Ar8x/ika8EkcfLYHeRbZu7ABA
t8GEqpf5yP2QfO8zlu8kC21iqKmgwzaP/V8dXl+mcqV8prYhKmsi7Tt2jP7gk+jP
sueVwjBk70ZDuqELEh2QoOb84/qqWkg/1JV2fzD9iYvfjksqCpWhaGaFj+AyZXC1
ri0bdkfNUSQaUs8PjjHoLSTjmde1vTRU9Gl15cB3VEFy/u80hk0WoftuqpbH5Vkc
8Yq0BOmDmbY1aukmwdZiF4BQJW0lxzcKBVhfJqU+YXq6zO7bAJX4llBXCNu1vbub
tJWfb3FfNVKH9HQm+dqygGvLJ87tZhZiZ0/TI3IZxJkDLEjXWWFe3iQ64KvC46wC
rnD2+Zdnh5DZ1FqtsGcnuFb5jQWPhGRSMYy+ueE+xr9rpj+YfFO7WNZdnUpzmWvB
wybiCIVHfScRlEyu5+b2zdxas8MfBIKozGSp5AfG6JcHvv0wHg/t87ldqGf+esH7
4nTXTnppLEhk8yHn5qPnXXCwIj+O+ANyyN7NiF0m5jTO/EwdN6v3ltBuZ/0jkPjh
gL616h9/7TgO1f0DajJyCGZnj3IQladUxDLegFvTQyUNIDJafMM3/hjOudeaGnNp
D7YZurT1T3U44rKiSP1BmacxDJ3HU9cTZXsLCEEK4sHfAnAgQRkE/SO64VrmiVhL
lMTS9uhXrn1X5798NBk9zsxGxlBqclJ+HBkjj8uQCHyXpZa5g30xfn4cES5jfNzk
mBdGk99UOM3gwML2VtoOmYj8vRdlDjN8M5CDOzeC3yZgKC4QHGPx4hvS9nH1jV7l
9IvpmKFxLpbehcKLkvgCFcxymYmNqrShIj63y9jgHk05xicM4AZ72+1Is8Na+YUh
6pwJjsQ8TFyBdL9COOGJ9xqS1toopcHRjmyh7qiG0BN0DIvgWd1qtR5qVeE5I16m
fE3FBKxGytOS9coEYMmzzPOhXMJYJb6h1S8L1GuJKNC0Sg2Jjva0qM+MhCod7yeV
ciuP2dPe/4n9PAHKiRaCbwozxFl7Qk5ua5OgZkMDj9y3IIy9sOLY3ZHbBwNBWFei
U7oO4j0PbLPAH1ngx6EmdFg3WlGUBfGde8aZmcmC+ej8RS7WmMkwVy9mgTF28zxh
luM0nMjHcGvw3XYDKNTcKQJLYqXf/jhM2ZVioNL0v99+/eJ04McPaWr5cVEFm5bD
EqL23SHKk9ETJb1keOIjWZSJSmGKLOwwokPCX0vg+yL4v1geCLTmtEfIvHfj183A
ldivNQ5yEm4l6WrCRuly3wyr9ffOkx3gTBMibnCCWGO7LUWsssEasvTJ00L4991r
fhkYAm1uYDOsXgUzLg6E5vHaYnjLS06od3pnTL5Nd1z2Q4gmv51jAxZkhGZk15L3
NleQw1/W+ei1/LZw2/2GmXBNm6vKzQ761Xhy810v48mqpVJOIuwRqdUEE/WWlk8z
R746BgUqrHCl+CQkO007DS0yFywSQGZiLZdMFcHqfzxdLhBCOyHG+otkGzSpzu4u
IOCnuzoh95+SW525dQpDs9KS+m8lHEVvDnzOh2sbFHcpQmi4kIGPGIzD6xR5qPkp
65lbljE52Pw94RYjGYbEFAGEiOS3gJHB2oQL1nfhi4EjK9l9/bwCukYmZvaoToBw
d6bCDWvu5ETkoHQCre1vpYoQOfnrqUdFySAFLGScJRuhe9ll5/jLAPdEHCdJnZKL
vd4yffq2SVuyrJsBNLyR54Z0bUeNE2HijEsZTlCapYx+6OChlQAc7g8ait11yuET
kWMHORs0kv71pu+8nc6OdSEtsXArKvgINUqaL/gjuaDsNNUakh1VTkiUTO8Fv4G3
ltgMzn9r7W3dIwg5Lk2mEd2+3j10wDTKfL9M0ClIkeLVTL792BFNsd8mFWjv3/Zw
qH1V4xljeRjXnItiXQ+an9LqQYSdZA2wXoIs7Gk2wIwUYu2RKNy8N6kls9azMKhX
7/zAuDISlXtkbTaoeDCiT6ncNvFzloQlw7OioN4mfWrSvFSfvCG+hZ/2ecmqL9ZM
hKclvfd/TlsSiOwRKlQL/F8XIO/mBrC20udzhzmsInuTnkkMB5IVPXMA2ORZCMQa
BHLSmx55z9kf2AUqo1p52zDwPxPLyXXiBtyRDmHrF3ZlLiN/Oi3ilmEe5v+SvOig
UhWFUSbBqhg7A6QcPf5Wn1ffpypk455tTdu/CTGnu2RyIP/sulqgBH8hFOdG0vpS
b4pCzvlRB63soAZor8RVcFaOc/Gas6FUrQ0I4HAS7/Q/tQG34fKkkqIOWZzqSeif
0NhBPMDsnm/0KOSNggmyQFnO8eu7LC04Osy4ibkWoyJ81V2dVw8wKjZRv3qmXWq1
T0QOAGuMZ+uobQexeqdM3gLTYOHLpqHoIiiNX88MGVcf04DvQz8G1qWL1A7dpTzf
07eXCa+4p4UZ9H6CNHqOttaT/qQqFpRlQHSy9tcG14Mh7I4fzhN8q4PaiASOR0uO
sfmI6o+xnWSi+EbAdXvVz7/3QwDDRyOnkPy45HP4Oo/1Rhbhb3iGON6+lRyNdkXR
EpfAxr2jb2wA30PU1c9pbbRe1t7ptA4SLBLgdsQ3SKmrIz3QuhQorEgDSY9SeYrh
LVSO65KNTKFBZMvv4rrrzi8o8ynlFf8TvFvrw9ZlDPbI+5GaorIP1+c5Tq+5fkT3
Al449gGhltRcXiiDLHSCgvpnZW52OZQZ9mv9Oi1hvX5k2dnZK+uAeSz6SoHd/d+B
1oiRROPYM7mMnihnnFLqkQ8Qqsbw/4kofXDb+krbce4Z2HLWmOT/1demZuBaHoJZ
4SvtdLeUNszyUngpYz7b+XtvOWAsFMmNRjEab4JCaNIqhGFlMR7x7a6I+UJJgd1m
vPXcfZ1aXwNs+KbAUafYUfQGoJbDC2enFJurWAI66+elUunKW9W7PCEt9ShkJVKm
/Qa6VVSJHRiK5qVwqdzprLPaehpFNxvwpU/9HGPrIzdkfM0lfcO7FAYmwF4OM/8o
dLg+lf/ECjtr9TnVnLWi8gTsVefc8kBzDBAptrtejttCNA69lxinPTpBo0Au4G/y
iTw8RqPYTgFx2d0w8n5nII16HAnHzG6GqrLiUv7iRjv7sboyc1D454I5ZpHrpmL6
uyhtOk/y7LAiVeW5zoXdpvMMqodXbJlNj135j+0aGefKkULTlJCsBf6O4SZ052Bl
DOA8E2y5ZXLp/Lrz6AZ1IlAj/mtha8FCpXAN9LWTD1H7nHZduJc3ZozV14JQyiTo
Lewa5SvfCkbddjOQN0aMcI9ykavQfGJZwug53Z40LupWqZz6e+wiJHvzcUBOa0C+
h7JyH529UvCrrrFlHBnTwF24T2xED7jgzz8XBqjtIYhv4WmqUjz8o4bTwY2708uu
6wU5rcmRZpwbamDvPr0PHiMSCQpWHRW7e+4iGQmG/erS96bxVMQ8wjCyT3L2GyoA
FrL63IVWcEG9qr6fNcwZwz/jwrM0PYCKl8wes6FQQlyiq1wOIHMQgI4PuHxoREXT
uTITDf81xdppuHL6Tbzw977y/N2Zv88+QmLb93cQUv1s4IvfUyK5iaqtNwk80Fdq
sgLxiszpOi9jtivHgzmnSKwZ631jKcCXDB/oaB3mfeamn90m/mtE9wqiFIgjDBx+
5xWv+rQYmRM5usfL1LrunDKYa+z3tX5dZSdLRZBZ1wKnpsIsTFZ6e6i4ZuI74S1d
MoAvdpZMERJFB9pnWGlG5tmSlMr2jPrKUfnqVRcCrw+Hm1ee2ye+RXHWrPjLwY1P
gXmLzUyMk1C2VtX9MWaRoOU2u3kviLnCpb4t8bg+XAoGyiio9NUMmdJnda0JBEDR
/gGwutGe6/BfLOHhx3ATmHGJMiroIDeQIHvz5PGA6N9TA75eer3ox0a1cydJUNhe
gJl04C31l1IoLrywlcU2qZUVGjDi32+FRmEX0PKD7lnK7JTC0uRMgcOOXVxIvkYL
XJhkGXi46kcu59iPABzTruSrRDb+LESwjPzSd9vL8uwp3JF7Y681xvzHGHpLL2uL
ixxcfGC5/A9obZ++jIIxHAmqfgQKt9BNPAC0Y1IlEVTNjlP8gI8hMj7DkUZ9y4vA
RIWkgXtWMx7S6x9cYLXyF15cfDdFuWZJLaxFKDt8w9D37pNBjd4aPdcTwbidH048
U4a4E2jtOS9+bwNpHyskpYvFIY2nH3jwv3JUWOqFKuNuoV4bsAVWNq10vik6sQbc
QqsUGa2vDcnwxGyV5BmDmfU8UuAFNSr8+R5Al2I0n7K6P4yh5TVHdf39GT0P+1OO
Zo2nu1rTkxVJcjQ3OL4pEphIJNgTQ6bS0I+nGFXOBkveNB87Ek5TYFgVUB4uNyNc
h4EBX+xpfH/6UduVmrq63cugBedtNgUhG30ZiS2TGuxVxwU416gLC+z6YCStATZz
oto2Hvj7taqAXV/q3QTSh3Rds/QbLaZSpYl/nSwXtgLW8gsjry5TWHhWdFBjC3zW
3x/QbaW047Pia0R9sGR1+DhF9rqTY3jMt2cmqg65lmpYR+7rYdhZBJTBbkPuKSkh
DIBZDdz+CLpF1Y2XVlufofWaZUCFydBVO3WBTSo6N1+BQAtd+8Rd0pgVcnonWlge
UP4V9Vxxzw7YPBgjgmLg8TdmS4zkBbeG+mzxr4p0XgFUTP3oMLtGDK5cKNKRCava
xOdQ27X6EiBZj6Ep+pwRYOOJlUZ2Qt2wUm/LCREBuLJ7qCTFMqiC6I8BaVV4ph1t
9U/7J3HIPA6huzkbsbcQJBniYGlYvlCPIqRLeHzj5yCUNfohf07orZK8n63rmYmA
arzSQDvU0ZyzQA6BpOJW0m3p0gY3Db3Xj+mX8kNn0yUQsxuF9oFcJRxQR3OdRJ4f
i0V+3UgraqjVwjfC7rzngLXIRaA+7ctTVjZuVMawh8gp3pMDNFwQUVsO0OKUrEEG
SRGBKTvOIz4YMAffaanN5s7KSWcVLb9Gn+W1EGQgoY4RkGWatHvpf9L5RI/WTv+X
To1Uxyeuf+2u7mMxZCiTeJg7e0LARmR4jt5hPx/6cWncJsR4moZThIfci7pLUOew
+Gr8VCLo6PJGcc0ddwxdtAGAr3xhbDMNBdHl3iWInXrSRvNbPVtc7J3effx5qrEn
dBxUyfU2P1FAMELWLIRAvBeQcAtr/XPm1Z0Ox9T5KPM7e1oGotkM2DgTkCDsZqW2
eX4mrecAnVldUNrHYUucg7lUgB/fijZolcf1ruOdR9EZegGNtpSSpG8x64W/YQH+
heLGmiIp3piMqQWMup1DU4K5KWgwqPVAltK7phPax8NYYOgDwW8KEn8Qj4FoSnR1
bWK03yhBybVI4nJffuKVi7x9DnbV3xe1VDDPc8CQq0htlGsUP4PL8sKLULsMcX3P
FqPPt0qRXJG1msFSvLsfTByOHAab3gZOC88OUqDa03nn9Uc0xyls0rxvi7FQeL73
MM3FQVR+fBp802ijCp4XGzP3ByfZwBDJ8IK8j7pbdVNSXnKsf/U9nFW8cJNYFG3j
HGY9KR5yg8AoNacL9y54WgXEDagcA8g1q/zwBCNgLSKoTV9sAZJJ12ocfYPhvoKs
on2QOScDH+c5iSeSFWd41gGZgV3cwX0+VifNn/Suey8WpLSqK3lXUOZGcvQo/apC
tjvq3HkyhG8bg2+eYn2GLrZt6Jt3oZnC+JeOyX7XyjUBIHGjQUXogXA+TYgB9xMP
ITu3ryvmlz+69t5H2Xhd7QYFXwMv8nAhWObpLIF/FzhcHLVTI9gtLT2j7vTiU6uN
pozYVQu7ETnsxbdfIo1ETAxofoG9P/KR7Pe4D6hbnRM7tuews6+W2mWByqCDXRFc
u+D5dsJRsAxReOHh/VeBxO0ZMQgXDwSqiNVD8ypdLAhEMZUbIa94s9YKtIGE2kTJ
3eNOHLUdJCkfChmUHdQzwZ0Mf5UbzvzXN+gHlUqukyehXMSiBE/903MYfMY+bKeg
gloeKXnXJvpvGodqKuB+EsIJ5Rtv7jG66fCJugyBSzYuU/KlOyZBPjUQDepazLyC
lj1jsLZ702wAA1c8XMO4I6iCkKOyfj6PQiMUx5g1PqKx2enlV06zCos6wEPk3wFj
T8P4yUfDqVN2rcMArjgQyNI+6gcVNSfTK7Vu5PyGE2SU4HEX+xF7AZoBRPNLVe5N
gvqxPm5hsKZ+VS/Vf6pC4rot79OWWXe7pIyxT6wTd3YCpWPMX2nfQVK5bVtd50lI
Fz9v6ATrD3B3nqcgy5Jv70vu9UCx/mhB0jDvtlaxnYvMyBjBH2xp+KSQs4xILOf/
PJmrislo6DbzowTwSIU1HOAVEHqvMh5xAhtAtthiBDEFWlVFaNyXEMLER4WvzKA3
LVSsR2R33TTfsUD2bQMd7iRgZ90Kz89NOtpaykb9K0ezWzOcStBu0MepK5VnGPCv
QKWHags/qmuLZ9lEe4ryHgm+tP0DHYpgP7lO1AyzihpTlwjlmxpj3HKdioWimeWM
jhLg7IaPMiiazQrD1vyJLdYy5i51OkvK8lUI4dRfkR6HAJWPW0Uq0Nsk8Q1H+WWc
bNqR6DI43TPQcd2DaQHfej3h7vlCZo4vdyctJ4kRDgUsIMnjsf+587zuuX5Npxqi
n3g95XTIrftgAMjCO/NStFV7f34jv9AqhEb7MyvJ6iNdTJP/R7v/CEXL1nPGtYUq
X8pWxlsbRY1TWA8kEJkfuZVXc34aU1amRqQVms3/dR8zrx0uo/fG/zza5X685ECh
hsljNInWRNb214wrkxw2h8BSpTmVhQqwRoHOACX6KAPiRGMC1cfk52+0EakBjUI/
qAPBNUHF1sEfC8y88VtCIBLHv+3arhPvqt7AvIE0Ev7QvRoRpBhZmwZ2qqFmegLw
CQK7HGq0LlBaaqR96HAVW72wdIwel+fg2Vonyw2k2y7ofaKX+5UPTr37eb5W8qbk
1Eb4wNm/HC/TfGOX0ft4GuI72m0zm60b9LexJuR3w1QHYTX+z5kKh0WNZNdMwH7D
1Z02rSbUcNaEYg21KkTY5vAYb0GlpCEuR2Ti8jVSSwv2k9aVHr8S8rp+7fovXmL2
wx8TNpwfPefloLtthMislQnqVqWf+uciVXJ7ZIrudGq+56IXil4eAcJJ+jUalLDq
vJyAmlyYTjShmrJYZ1OOfBYPm3DH1Bb0Jbuz3zW1MH4Iib55TTb547uSbTT2q6vk
EPqcxdfQ+mqOaeGwmPNyWt16JpKnKmcfID5ofO6Bs5k6exwAGYefe9buKBmwS9U1
5lk7p7akIUYVLL4SQNe8yhSR89UT19Qtii9cnx0xVavkqezzN7vErl1NArXwg9Qg
4PlFHOb6r7CPw/1aL4pRhzj5l40ztmpDZO6nbpC6SZY107NGmFK7y/vg/kBFMMzi
QWjacFQzEeVXQt4JC4TpULlJs8kpAoa9nOiCxxRYUAJegoAdgMGZSPKxExNjcT8X
V4IwWBSKv4+tbWvpZRl5VMSiNGjK4EDrQfgPLWTh0lGDkFE3SR645wwiOnJFn/JM
KBdrA+OtWBOmj75tMxSdPjYuf6AJYoud0RezeFhnef5GvC8FKIP6LDAPQ5sSMNmd
ix0+3BBxoieTI51uhBFvKSMQE9U55PlyPy5FforyBCshXnb0BNmKUGUvwaO424Na
G43614WG2CskY7VYfujAdDWlpvSf9R8ckEjerGRVR7ba8lQhrkX4xlZ7OH9vhXIF
gCrojiTrsf23ljhSfsGld91bkRo+MjNYk/9VQpJuMTYoaIo8B085hKpYApx7fFhX
de1kJKfOPclWaH480aGERUPd+vgOlUqg9Umj5mDF4yEGQkd5zfInk4baKEOuvXtb
Nf5zWSerNRwcopFX99cwfxX3adCoTl72MbqPUrFiJXG3+8XBkOfFsZPjePckUzzY
/ba7/MfUpQ+MAWn/N0NoJRcE22enUoVULVVzEOKTRGuPF9UmBNF2itFM+oJXMJjf
KRopQnFpzVd7iETlYA0J/kw5ChSvuotk733DZyJoe3JZXWVAWa/uDBLFdCKhj1MU
/B/F/oHJHUYBYXU9cNOaLpRnDbRyu8FGj+vYNHYE9nuDqhPE+8yi9m0qrfJp+KDv
yPUDuy0GlKKU/7RWLoM0Bsl7wIxXu7s43o3g/trNPNM+KSTfCDRD9TvUEfNdcgsE
Xuhsaic3z8GzAGfyiaIDknkQAndPYFR6iUsaYk2emhSWAQXqYIgTVzyl4UQhOOdS
pOr/ubxEq5CaC2E/ZiXiLC2o0PnGMHI60K9o4Qo5dFZkNQFKnrC70EeRFfj9hd1J
P4mhC7IctLwt53537SdSi5JI4RInTS4KvpLx/dVHrrI3RkYO1B7venk+Gih5Y7RK
GTaV6ne4ie8rafFyKC9gELOTX4d3S4YDHxIMN1wEXofpDKohFeVCaEbt6EDekzgW
3cEbqsVwEwS4hA5nNFwkWCdHvqdspotar1tSsu4lsaCo+OQ4qXGcmMlaBmHCS3+F
wTccApM/2MskTdMrCCEPqBSG7Vy/vI2VxF1Rqt4grDQ34BZ5x6IxQhz4puvfJN8o
yeUFj3BlzhwmB/EzZFrN9eFo4+BH4I9RzkvMF1zvN6p4R/73/HvirqbzIS0Tf7pI
WiLR904tA/3wiVZ1NdE4CsRMaKcDdPHGqzyo/3bYHug3btSYQoNvemflAFjbut5O
mwNZa5obTJHyDb+9TLIe2chDr7skuCHrvEAk0K3f4mTVhsWo3Fx6wu15GG23T4JF
Yd8mTaWPMtZTDodtbyc8iHllLF3h2mC/TkOZK+SDEqP8QghQj54K47gWtISAi5w3
AqTzFb91m/WbGa0vFwybaXxvcIbeJRow7umARFeSjFoiWMNYNTq5UqWmVsihtHqf
Erm1Mr+cqRbc1RmlZXxDniNdNbBqC/5llkVBJR2qnRRXlvwQ/iZxNrAV+aFwNzYA
s5erCCk5h1jQsXildQI3ee6nP7+u1X7eK5HpSE2U9EGnRKHDlN5bV873n176z6tu
JMp3h9x1PPW/ZPywjtCe/bdzxBWqhrBqJyIpeKNJxH3dWwyg+Ahyayu9pbpW/4aa
Rn4p1IxX7H5qBrW0z9QCZxTEZACBQHmgW2kvQfnzXrAmdX+CwgckJPAi4kTKrHJC
7qNjDcxIiK/mXZynVf/GeAB9kDYqdIdki+H4WcOu4i1uOx2kOaP+UgcuFmzN0ah1
iFeIH9w/ybRJWxMrAjsdkZiPc/Zv8AQiX5D2PoMKWG521+6ENZTMwIYJmzDc3WC7
OUB2zNo382yiliMLAe/WzKo7zZhVCy0aLOvP9d1zTQZ/9vq0C9RgD91MuPnWav6M
R6wprwv5UDJeemKhRwkUHMcqBqefb+Hgule80FSQM9aNhkMAhanhgi/7Iksrlyuk
NvlOkn03o8G35PrTqCAabYAblaA88TiMufWsu5SV5dSqnSBusYCDKmlK1cEL0akW
Usnqnt1bNYF/qHsdxYRnJxKLd9Qyceo3YyJH0zATsEn+dYdnS6jayMeyNLpLZ9hn
PyIw+ru6GS77VIcAPgMMrJW5jnk36YlLn7AjCRKZqWcMBE6PYVMjA6tIOv8d5Z7Y
theNdU6upGl0sihyjxeDIa3KXw92tOwwkdXbjYuVWYC7gtzpAr9956BN9dCkzhTN
osYUM3nkjTZTqy4+qaMST9C8TUmUdk4M5I08sizxC570Aamuhw06hkkDQWBSfuTW
9h7LSrqvJgcGkQiZJVkkhpOJZkeTWyYhto4JwOPTg8ZYR/Q4BEJz8oppmUpopxzZ
YzreoQDUZorlaIXcWrjHXMWeUSmGHVGJp+H9BF7Qb8/hl1WjOuhawbKo01eVVeNw
Flvw2xgZMSoWM/+TbHFx6dTZaRUucRczLCcN0yTvcgNUcZRW4TqKgfTQnYUzd9T3
l5HjrdhEK+6WY+km8bpavU8GLCVjaBfM51Vayhzf5jCjMsLIUrkxtW0LxEyNlwHQ
kcyKLY/R4T625GvsYEugifvVxouBHntYPOPCbowCEQfhrvyzxkMyzJ4fFgPh4uzY
9ilS3pOQWlJzqPiKhDEjpYDxeWB2KnqT03ALEKGnC9SZ+qYtKQbSlX0rLHitIqyk
oU9aDSQMgwnirH8oXV9SJ0/4inUIJb79gn9qEaSJdHqOPQVZwD/E1WgHzlCvCzmH
RgtHQrHWF2VQSQSCpRZyTbXWK3gx8ZW4T2hQyIHg+g0DqaHuNpCAbyh8k9Nq+Xku
1M3D7xTypC8KW36h2Q95pXnGRz5Xk3gPr10qsP0j+vjrRqlT2WwlPA/4uqSCVeoV
hbrclKipNndEIuIYqE8EBhoITOI0rZCuJj5aFqafPFVyRvJ6loimf9IlSjBPSo21
Cgyj/FGMSea4hVoXa8c0sCTK2hDQnTzzQ6iKF/tYOYt+iOPexPuJWp9/QN9okWYT
KkC9rku82qyIjMs8SQiqutrvwUGvcu8vC1mk6Kmq3fKmLqssn3Ea+mdBV2vyphyu
FaVFLQguR2s4QGVWoKncp7BUvarq3GgeyCoSH2guZtZPVdfNM11UxrQVeYQSdFg9
B63HuqdAdbUzXVV7Ex6hWFp9sc1NrxH96cGc32nvoeZisavnc28wrKlcK9S34Ssj
R1gjbwOQ5BherNRWgeYBjDFu0D4CJnTAQx7Cp4+28dMyB+AJATwbXG/VOwyRLeGI
IS/7+5iv6214/UbG7Rhb2kf88AvTT+LHZG+mIVJHUce2DTk69q16u+FGCZd2NSvl
kwcfby3sz4lhlDaK+M+P71yoWOT2GPqHVa3UnfVwz8u8SZngCQCJwcyDdE8hIUlt
MSYM1wLzXFCsRLR+KyC/ZpS970h/heD8RZL94xHhIBL/n4Q2jakaB9haTDtsd1fH
IVIJp8tzFVrCgRcI2XkoL4MOM/3hX8x8PxbRole54UR+Ln6TpTJGrroy3Q6e21Xc
FZfQ/mhoWm5BqxqStjobSDLO70H0DpCK4SNBcEe7PKfmro6nUfVyWrWZJtee/qfK
JscK5DHvnHlwqwOyDpM0NCzcfsb9Gt6KrXCk5g86uswIsZN8NoaJziilmfmD+U1Q
l3wo2EOlfRvp8FO5/6EO7XeheksQQAQnHKv6+Uc4eUaiHItnK8nPT/AfSrceQun3
zKBtx4GtoLsZhCd45Zgz1+AU5PWTfNXGbRaw3T5a+2mL/l90s0CVcU1M/PBCvBTv
zjMEscC39NY0Pa+8gKxciDYsWDQY11G5DXIzvTDzgK2JYUgvoQZRvGhbizx3zxKo
XqbU/9lzpkjV/Jpx87i3fRYSNRu3VwPREtE4vgjwKpBS+ZQx3/XTEZDleywtrsa8
wudUAsI6gFy6NP9NvuwajUMpQI0x6Dua2mrgWjY+TGhuAQM81O4FmRd1upI08AOQ
adPOLT8HIPqwptOCVT9JFWYJ1UrGnJKGIbhNMbbpMGVJxvlSSU9srashDk7VOUv4
l9+Xx6mfAjqfbLuCPZb7jwZpWVczkN1lDN/prE5GdQ5OlMOYoTPwjx+rOQIPoDwi
tUdeb3viEm5sllt61fDRG3Dz/QqDfmn0ao+602Kc29PVGXLcJXSn6HZ8TJdwO63y
TCQVuQyE4KLtZ21qWovaJQ1JL0aefbx2O2z3g9qVT43xxSsspa8HzKDXiZdgLAux
wSB/C8tDqdV5/w7cxK+iPxcW7QqMGj0T8GrLGVVcyERrlCuIrYg8jW74TjHjtTKh
ZPGtx31eCeuOqNGCgURWujlJVURSKXqrrZ2HQjJVUl03c+XE5a5jyxmJBsJzzdmf
hV5JUN1zzeYba6GXjDqAyxefV1GBiwI2EzDqIABnMElmSgpuv1n4dF12ihGLQxA8
uhWsEWST4y6JOB8V/3WxnQMf8yiEy5RwlXsu+liFosW+EsMWQsMbnIRf6Jq1mOdZ
b7j4rM9zynS8uC+u4W6IYYz5ncyLwdCNizyFNh0ni3QbfDKYnBABbpwDc4PekIEm
Qy67E5JDsVoYDpG+6VbQoqaaa5oZUNKB9FZFx9KZqKPkUpO0K51E6mpG5pMDN6RL
RoPHV9M173wcJ1o64+jIBYbzmZS20DRLmGs/9ftcONZhOAmeiTqS4uBmrT848Mwq
/35pn1bW27xnwX8B7PzxoUa6UFi9v5CnEYhjtgT/WqIbjKbFgfRj9LQ9Kqux9W/O
blruEj0qlaRudnKVqaduLAr0x8/GKhvoR6ad2dEa9zAzJwXI35+pbK9xYCwzpSap
Od2SGiyUi8QnQnfPNWm5VtFGgIM63uHC+rxFGtA0GdQEg0TohfJXqSTdCFbNpB2G
b8U4LHcPUZ5nhh395GYECGuO8aX7S3JzRTJwcq7qqkekZkfLRbBiBhPuQTRFk0OL
irIZ0iuKWzXXRwzKzFiJj+yVPpwv1zdZoshj675WWfWNn/s7VZKt7L87p5Pl82V1
lpHKOp8Z3GISf1Nm5W7CY+zNtBfZRDoH/U6Mp+ccKB80sCDYyUdF2k+IFlL0mcYo
ucNqP7TzH1/jug9rEq1cNS5W2oSx619EYCJXbYw76UQfUa4l2WyWC8WunROMNz+w
DRTxPrLc+fdzoo97ruC3cNO7mRuHf1DE8+ssUaw59YE4yUlcAY8RD375D3wSuK3s
A276TywWoM58/gKEvXbvfA9H08Y/atfnnX0kMTc2x4SZCiz/sP42144QhrT34SOS
P3v97tN45BO4H7GVUo1mRe6dm+F3akWuH2Fi5NZVHGfWir72PEOh4aEMUXuUwoho
HSNplE0vlWJFD+11M0LRIp6MAkjCBYEQG1l3A2XmikPGKZVgmA5RddJ08z4Xeg5l
dQ4BItsImwgtJ0OqsN8KvewTvO95adsXVHakCO9TYXcxXiGBi13jEgEAaxmm0j+m
INLapjrLqmQZMKvtozz6TklTn3qLpTeDJVjtspoimVNciUKDUcyjdywAdkVvyiKD
O6a7JUqU3xrj/63C8lEdXzfcp5I644Ml9zUtiD7v99CCFy3m4Yub7MS9LrmLJxrh
pEnDhoCMtOE1MXpgMW5ewzPQKNTnnrXSq85qSW0WgaU0r6YOZ1qjssxupcE9V1ji
P9NakEvEk88OE741wwJYeK/g5bO4oKwXjDXJCNBoJ6dUdtCaov/2qdI3aJUgZgri
EMP55RPvw3JE30hygkWr8lQRl09M53SWfXZd9XK1SbBYo+aLBddZUQdqfnV2Cb1r
BJLw9CAjXJwJ02HiWcBzMFEyE5gYvnwPzNFQTQGekCiytknGLMAcR4CisG2lSPBv
IDSnixSPYWHNSpB8MZyVsTtnU+ZCINZtU/lo25pgFAmheBj3Z2eQ4uCR9Fkndu0l
xlNJlV++tt7PkPZWYKhU7CZQacE/MsjeSGlYwKrFNpvN8d1AEheWE9VQfg+U05tX
DeI3qg/JibjttBBRk5qbHCeChkpaaG69avcKg82nhytJdm6asNzfg4xHgljAR1VX
etTjXlSXbJxmZiGe8/2vkKZcEaxWeov6UF7SLXYdqRyOgR5eqMFHZFqpo17t+KKw
kkCoiVr1xZTx6+KFlGwLpcjYG49OwJhlJ8surrgz7vNM2Sfk0e8X7vjKCbeeRiOb
K3ovs+XoyeK6OCVAn3m5Pqqm75tb/JPPbQiw9GWEkMFCZmOt6NDwPazUA0tg2B3J
U5+B3nO2f1nBKjN+63sPYHlkMSZwy9ZsRvWiAsqTpXXv2EkJB/0gzsHvFcgytYpY
wVkXO4SsrRVFe5psBQpPKhlQ994UQN0l5cxw8wEsh4E+EZoHGSmyQAgP6ySuXDma
gX4Ki4uahtoaP8LYy3fibThM9nvaXB9Qx14yGYVR3PQ5LIEn0m6VLbmfWXbjojHb
kzBG4xojTV7qDfqD1hNsxkkEXR+4D3mbkceXhDQTGdD3Vt97g87knibFvp5q9xlo
zwIju/vyKC4NoxPE+alZMVneAjoIMWRDmHI0ph8e+AhdTpxlOVsy5Xi3mHOhISm9
vglimRKWb3ptNTY3SHILF/JEM6DZ6U/kAnLpLHuw0+WDNcmUCCCrcDWGDVJvYM3p
iRAVWzzqjDsxvQ7fVeb0nVJoomwBwbxISBg9LRBWedmP5TOW23mqWWRhnA8pZmBY
832WrGShf0P51uyYO+NIlb38B1U9A03s3wEeSFqO9KwfbtTzvkb6AAfKVvNhum4z
OM3Iz1p2VVJYAqzqH13fDsIwHXud9R6vuWRm5+j6+ata36sKz7i+KPhS0A4YOE7L
3YWfOmITRUXtTocMRfF5auYD/SPtdduhIVKKN8VfMU15fWXS5RIx1ciiuoSCgiv2
pLdBsrcyzWISxJ8kE8CYHs3n77v1mCT97Ux0Pu05MCLuWGVAbm+9N66u22RRXes2
2RRcn65R6DuCGc2/xNk5HjJsnwE14LZEKxaUX0A8kQBRLPgxax1wVcYEvSAVH82h
Cz1UYs+NZKTILFJ7RVVUvgh7fyFZrFWqjQzRuE2QfIYwbb8A7U6w3fBN5fXxhS/3
2LfS+Pdwwqsl64u2EWo2bqjWPVtPn1CojoXm5pU4nDClTDXilk0SdktcEP3a7e0M
+hVAi+3IRaKsUbSJ0GCFbGPQ+cWejfpL7y2/s6F0UAtQwTG9C2EKs/f3cZb4+B2w
knLyroZK5XocdA/bBxEOCtLF4+DXdqOlqMXrSRsnLPg+gVZ8EQSnDErXT2Zep/7p
E70HdqFXWEyhwgt1x7a9EHZ0JLR9bUDEvRDXi5bHcm5VxTm7qOPnF/xtSzKN2k0X
6EhzAAOh2sJcV5DTuluhvx+vOozPcOwIQ3wAubNKf2B/KFN8ClVflFRPAONKOGrg
sWFUy1uR/EFaqXahRla2QG0OLSx8P0sVk6merCzyvpDj0rv0R8gxGozb2AeTZUK+
IaVCndMiy0REfXysG5ZjCgd25g+FTacJstc2t9+ll+cHN6fG3PY6y1zLHy2MrWZ5
iwX6ZrhjhhAoDC6NSS2RIpQtuy/5cKuvutP0oq3NyQJXfLTvGXxWdW12atMPbsL8
iRS+Tz3S3T8rC1KarF/JrwPe6ANKJZ7SOY01MJ8RDsbWqmHhRJ6ngeW1X9SUPP93
88m5nKmKUqMLIIrt0T2rxQkxhTNnFHYFiJPFL7vjplOmj6BVNFxCprt6xJzJ47Ay
8DOVBLPOuEjrS2u9XbTdA7WI/JZXWzahIaRQshorMMkHAnoJ+Jz5JlNYwfWR2Xdb
TnQzzWgFl412Kh/DINses7IWjqmQVN/yI6Di+G7qjSMn0i1CE86ccez5dg9+7pBQ
dqConxA2AtzEXmb0VYbm/GpeYjhCokEYCXKIhDiqz1nhtICPxLI63D0aqEmINpLV
taMuxYyECqzUpn1CUtXUVXYCu+k9P0Q2cv9pHbdx5RFEK+fx2fNAbZW5WS8RhoMO
drFIjAaG8IJeHVMPM+q0D0KTrS3bPx/7zjE3KT3ipwBVCjZaGXaFgzDsqEUuH5Xc
NT/OGppQODLaMLh5MSr0Y/h7i/HFcA5bCZ/t8crMZYHMN/hrHKDPBvlhYdcw4s6a
dL2wKYHXDCO6hTnH+IgZ3KnmO+EM1+K61F+pD+hn4mmm6sB8meZXlFVSKt/McbCt
tniCS8zW/o6LNVjRDgLOQwAxCJCE+n/bzIkB9LWYR7M/1em6jh4p9diTt1MYJAFQ
mASkPxShpcdxehptKymRwhBSUNYNMUzcK3adem29kXjzSS0r8v2be0fxPG7s/M7b
s/hYMpK+BrqT1948oDAiwOUWRmpqyX8NLijlr1J/B0tV3ogYDRIqcFuyO2H86rMs
v+ZVU8ZMDN/yMJZbHJkmrl81m+6Ju01gOXfgXjcZRfrY56AjH46e4XDuKn8oOql9
MPBCBviOQDXlGKt0XQv80+9Wi4rJL0BOxLUIwgoSi6/UcgA4EoBJQnMM3Rm7v4nB
X+vzIT8SLLXcKvZCukCtyWsR8/cgBPwi79rxW36wXQyCa8G/hEJzfZ8hQ/MjRVOZ
sf92NsjdsTTPdCZLZjxvWM/EviVEJLmGVg6BlcpLTvkjm+p/Nni/alQR3qwB5sbW
Vfi3wwZvYWsAovzdnL0u4+JjyLm7XqSDrxrJhlS6pMhE2Tt1aEGKQJbjuCYrBvC3
m/u+yI6vJ3OIoH6mvwHP2fRRkxA3upTc5LMd14Lk/FAuVuxPt6uHyqOCIGSQLY0R
w0MAvW4UDlm+BtWgt5mp6rg/HDoyM2o6gnZ+3xRBT4k0ZMmtROxtxqudc2qzHpgG
R+NVkisxTJlJStXYH1+GaB3BmRdqJauB38cheBcllIuAdzk6l63uLxHs4ghVwtLC
wdO1UINveLcLhJIIL6JGFDqNTBjCnxEQzJGWWMYuu7u/K8FfBnbo0xYhx3qWM5B4
jkjCZbAc3JDSR2O/If4d9ZyukFyajb1Cm7qGdJBEe7Z6HfyrZIU3U8u7iZo1VXMq
yE6OhLb6WS2gNfMgkN43dLSDi6/ycnHea51VEV0XZB27Af5bJ/Affutw59iZpW0l
eC5uzPC8N+DVXgwQZWP+IUjP/s6ZzFCzDV8RFb2Py3FbCIZsw6MsIokuCAFctnfp
HvUBYTLt0nlx05DxeEw+W1H+gGcUFss3M0/+v3BSFzxTD66p+9BPMDeaSbNm1PNX
Xg3RjI4/VRMqLlU7QsY++O6oErrvclxzMtIPl8w6O8p1Tr6w4Kss1yFdIor9GLrA
FDor1y6QkYTx2eS3v9NTlJxMM6rB2fnjSNJjWpqDnPmu168vP7cRfawdR8llfUU/
uoUQKWfHGQa9yWBdUP6ecxPD/izRxIM6mWhJCm0JrxloU70PtDrA3qZofmPTpDAs
j4v/m+BuE3yHX6LiWQblST1dHi1YVImoSjF3kwxEfseZtEddqkY+qtt0Gfg6eyr9
OUFc6LDGN2zDxwkiNh1qB0Uh2i0Fqq4yd34Ve8QVgSh6iCIsCkw74oRwHxYcC5D5
FFOIxg0VfAb/n8lW5l0de33GMfB1A5UUtSAehZzbFmxh5SVz3UcTUhU6jQVPcPym
FY7Z+c1uLqWM0rUKk2iOB/SvC4DVQfGaxSGJmY4aUr2LwC9jSDlSTCUwpARS1/u0
UHQ0JRhZJrJgPH/HuUzU4oDl1NFlKbzXWrlMZYM7hQKUDHBYoxUaUcNbZtS3C7uN
ao/5GemyXDSPT3YNCf2ptQ1radnL0Zgxa7D+bEpa7rBbvHq6o+Nhfd31bLXaBld+
DM7egqNaAyiMrp3o7q6fr1+rwLUBIckRPl9xBqQs8jhvHcezaBfs/YFGyylq+eWp
fkW5twhkDz5WT1LylgOLAWNxkhsQ6CGvcO+QpQB+JZb/HHgB5aGuJsomrI5IrQxn
tAvnoQwCUj069utsEDQDMmPjB3slR8QMiexIvNsovtOVbeMMxdlLIQDlhK8pSF5Y
0RHf4hMnYP7vVL78YGnPt0HjxMQnamTZaXMnYWCDibpYFrE/VMeh7QPm2P4BQERF
qBPLOufVxD5fXxaDG0RxLxMk+L/UpdiXuPg403pmUh2HOgtanM3X4Vj6Nht1kQFz
tKoG1lrYUYp4eZKGV/7Hi2TZ+AUduhdP+XYYmbSKOYiZyPc6Ns8F6L04CLqSAiXu
f19zP1AsrT+w42v5nqDAvqxCtQCYqdHVggziHb7WUFzJUcyKnte+6X/slckAhJgH
Y2zaTK1nA1089+EFQO7dMcjNu5t9wixFZ4SDx/9XPN7ittDJkL5CRT4bRHYhmAll
ZkyRcOSyeDujQAVdCXs1ErCoPR3eI9wvdmv4JdqlAkq1XkuZS/3QRfjU184yLCws
BJM4sqQWMSA9etEgXz7KCLVEQlxvD3K7T3MAy7slzi/YapIbZvRcU4f45SjybF2e
G1rKBBIe9pFiS3VFcpedOxspcQi/G2PxBwyYk7LeOq85mahJ0dkGKmrSqt8kdEfZ
ZjPhDGgjxZLQ46b6c2P4TfgtGYUECOYCLfarD4qn1LOPlzJbfWKQpjAFdLmIGaHz
QclqVWgZL4hHE10YE+OOvdUDhIe8NVLN5awEouhFlVE8zdOnk7vl9RCIrl6IBZpZ
KBVv+bLq4Z3m1frX0JDDw+bBXqJvCz7Hi8tzZvSbM/Q+L5uNxiNdkanGyW4PwB79
PZJGiNWiQPJMKvbtZhBMC9jAk4mAJR/4ZVe/GKmW/xPNv89FOEiaRGgFCxMlWx5H
ur54Z1NAHMLqBRQYpzZnSQ1jyqc6MY4ldR+5l2M4+jCkbLl6PJy4Gx3ka6tqOxCo
fQp9wmIde/lyGUzKwgNn/O5VJUa4mf6juiKdHtO1tp6wbru+Q/cxvzaeuhu4RLQk
J1NfN+s1mxyjLE0l8f8yBZzQ3VaUq41pXPXQAwjxK8wBDaMEwifpMJAIE6Te0CIx
OaKwjSj4PTYDkZngcPIinzrqHvQaZLlfxA5zy1nbDQ2F8N6BBKY3E0CKUV8ZTaUV
qABw+s9v7gpjDCxqzIyVLjl4H3uvWHJK17P9szfQVk2S6vumaQj6Vb+hNLUkAa9h
Oiyr4OMiRaC8HewUuC7mS+4Kjn8MGYClFl/R7TcwTuaXcnUvt4JceRlzlI+oKMkH
qPGpf2Tv6XwmDfOad2agc+5Q01w3VIUbf6hd2EOrE4ffrYEf2iERnqr1NkjZui+X
8fDGSB5xiL6fVxVuvF/COTKl5fxvrV4xyIggZkJF7zvlpPl8r1S56evAqv7GvPiI
94FdNP10BM20re2AhNxeyd+S+a8kPop0k2WXQqlLWq7F46mHDI+6SPVW7TlUK9Ba
j5HLQcK9ZmQBopWHKHJGtBg4k7dhCCUR9UmFFFqqvwRn9LrLDk1SxliVJwmJCBuk
mN49rrijvqpsOUoEEE1gMKJtANvIHJFN1gmKh9GR9wAyuvX05OP5S3Ga/MJFH4jX
s7U42z2yHlBkiAlSNkteHM4iNBGzJ9TqNRdN4ef5NFeiaOTowsvAYV+E4Pv+q8Hz
1OEPLbpomUBhy9Hbq0FvuXTvzCc7LcYQyA4ppv7dlw8FT2gWpZsrYMt9c0bVqORR
lkaMOd6Fon2h6yHbc2eyy2J6nKGSDpoTVDN5hbtIgUee2O5QtRF/Xty7lkZmjoPU
gqDi6Wynp85qwM+N8mhrZDehj9TNj9a/6FAKWFYCv4zF5cx82v/YVEW0EOhEdBJk
fEfj87blo1T9BXRZmwp4hZdJVW2wnFXznmZLLQVCqhkKDhhTZ0zUo9/pwXC8ND/M
fYTm81tg/n/lcof4cPcQU10yR9Wle3G+Phnn0pm5TSez59vSrbjuUW4Kn2ZewWHB
a5x4D0xnMeYydRmP+BJH/rSSjT31wVfblm7338ZH3CryapEyMS4A2GwQxcaWesp9
nXNU28QSLSssKBpjUUwJClsvlgBJhZ2HQlJ5NIqX9GCtqULr5sMV4ZmPj6k9cMeI
Jy32LBsub8vrqL2ptuyx95PjmJ40e3jwzNZEB7eLYCh7YvlnQboQU5u0x+deywrC
rTt8yMOrae4T6FoLHYJpKjbS84XVo7CX8BmJc6Sjcli95bhPS6PCUC8KOQp9z6zD
gF8aacgPWP0Fq8HxXWfvxItf/EjW4pJ0W0pGe2GoT9AHoyvJUe4EmrLlQSQX712g
srWgYMAcLsvnPTdSFdJvcJQegZw3qOVdxsg0YhYiiIIFm6zyvUXmUAwjoCzeMzCw
DLDwACOUnMpeVUBYCQnf7sSzzF0AsdVwQsOcVj3BZwkAi1STHDrOo5gWV0E25vH1
eZgNDFKjm+d7jdHMe/di8GigrecwNAnP6BYXNKOSawMN2p3/r1fNCYDwNtNj9oh1
ASOXUNAQJ4Y8vwbHm1SlDzP9FCVooakmTBFqncqCb6jcIoFyXQag4AI0X5dyDNtK
W4i32GbPwMc/gZmhuX59ZjCmd9eS/VjBKPM44mfm5K3d+9zuKnGBn2aptls/mTqe
USXWajav7UWI3aK7ZMbfh9SCI5SndZAEv16ZKP2voEiTMUBFgTC2kBor2o+FVDqE
k8eRrGt369LHnIvkynDi9DvJDmsZ8wzSwCOa4KutJhJ6i/lLw5IvqaOp6NcAWBpx
LetvOxABnK+Q33fsKJR4gismVtrsSeFDgrfp21v3DyYq1viQwx5cfUGqnPCOiUVB
cxz4O2CNHPumapj7aBoO7mNsU32cyPunIMWq42qpfLq+ehg1RNNlqyi+Nb4h1Vww
0kNWVFMGeUfVGguv3u2jI3ax8xWScQcpzckQs3Cx5sODOWmWNDUd64PzuX9PTtGC
0fqZNAs9fg/LoFH5M1mf2jDos84wDUb1xZXvZBUGaued98Kx5MfGMgJaYLAfAhF3
+4wfUTblhYdMsE5bZW+yu0RWM80TOCHn0OaPOKuOaPxgEc7zw5oWGxYlIcmnUA0k
/11yEd11PoQVJhW10Ef5dqnOpGuRIpoTaiq9HEmUwzFl8uoMBMx+s8rCE9pmWK4M
/R0eGkHYYW/QUih2TlzLkEmy8OznMdCyoUcJy5cZkTaR1yRjiE2vcvOhZBLr6WBq
LPQnEy3d7cneywNVISI6T9L4kKOI67Cs8AKToludXQ6symWget1H2rRniP9/xKpa
pPLv0gY7nQAynBoaJ6PQ1tUVhHmO7HxmsG4o8Yk467Xjw69TlsoQeK2ayOLLiGc/
YlkBu+CXSKsi6xkHOXeyXCnHLzSenfcvEi7FDsR9+sXuCQMkOruRXoLGc/g5Kkj+
T1YjEQRZktPAN9Y0fPZgrvetYlrLAJk2cTl6TdnqSmah5WEk6i6IW2M2ITLm17z9
L2GHhX0xuWTR0PVBzppHlh+YDnDcet8yqOE9yBPk4EZDsSqXZud6AUGg8KqehLv3
bAfjlSJ3x1o57rvOByFy/lcEfdCnG5dZ5ecSViNI+hLJn1m3SW/ZqsbHCLuf7a2c
KP0hNvB1+sm01Fr/gPPqsf5jLmjSGSbK1IP4KgfJs946S3Fagx1GBHTJAiiXxJ8s
gjXWEXUUDxMuumOHJEnAVnHJ50AnQ0tckjAEY4sWxALTHQvFjOycoJOfMP+esEWn
bZT71bRqLueiJciy0GPmqUgxxmT1TtwrbWyK9XKkjxsQejYx9hWlKHHMp2ChxeUh
TSI/y/WwO/b0WpYsL5OOWMSJZkx0khD/Ld7ZLByjA4qPqHGszNzuyKo2P/a1Q4BI
zGnK3zsrBM1LgqUvJBlx5xD3JzePT1g+KbjkkPuNCkMTZgcXdFaXl18JwNMJsDsn
uUybCguPEtqFeLym45nXG3fgKRBQ/JKTY6+ghzaGyiWvfRTEOmkarZiXdaG9x1sz
OR9sif4q6K3qgw7AhBFVW5VQU9mSpox+P+qte4kQOhsAxZ0BhKBp3s420530R4XY
NLJK3k4SNzzKJ0HNJp50Gf2z4/jsSu1hYZqvhtFXVsuS2CAzQmvUJUXAiLWkWNP4
PO+3o/NpUJz9veaqRNhp3PNQm5PJC4sJMDIfcVHPzdwKKu9liRlz829sxKN1pxNM
KSOlb5qAA/qda5GTw1S1qfFrahluyKUXlSmqPjsCnzv6qZQcy2vFWVkVPQeSPSia
L5JxYsrEEgNieYZI8Lj9TYPSqry63l7CczvYAbPcyzpXq/olmnqyUzeV8Dx4lOyQ
NUiq/ENsBOqMl5sJ5Wbl8Ao8SaokVpnUnEdhbjspypOSTn+aPvw1I3ymrHVYhGgH
1YOyRCDhAlViRHjDjvPXmfZ6cvct2kvcHSpMDBBuhSefaLN4AtedCDM1/yS+Gv14
gCmm7yfOyXw+WSVjDZzQNnpCtcQw9y9ZT9OOkQmg01RKqGjCRgvI5ndfkedGXnYb
lybLZxBIQcOwRLOdW5d45bMs7xgtQNNjkzsY9xwL7zOMrCBuD8/OJXxHC2BjuVI3
43nkfjNAJLmpdfeTPj9aldjR6W1/PmzTH0XE5c9n7PHLHZopzY7kd6ty2FNvW1GG
ljOGzdLloW3C2ZxVD43MiwY3ESQM3FJaBHZvGxvQ8CQuLMivF919Zd3u/3K311AA
N/yj1xUknUqbqjEtnkm7WQ1nsBNgcXycDcEgHfhYcnkV43nfcI0IBGpcnwIwi05U
uZxdLW7+w2FxwYsOZQAPX0XifD3ovafLwulRGLYmP/7ERpysl/k+r1GsyJ9YaUOp
1xPEmo4ZJGlHS38flcvJTrMA5rQ/pKHd4iu6HfISCZwha/wHiOwMnl+y5+vbqkrk
CU2enhLmivXyqh02O/3IstyqYF2KFAku2XeLv2O+xqYzajUrPNTcgcSf6fYKymlY
X4TUoM69OwqL2w6RmI+DKW7nGQbPJmbwwxp+qg9huTaVw5Q81mMbb/kgsx1hUb2a
Ss9RODH/dybWmpWmdpWPuVwX3gr5hawHtMjTtc9MscBAcsscqfGmlHijH4AXBQHa
4fVxm0ujvcdTmWHmEOdqQuu7+fxBVr/9UycEZ8JkAC4pi9HS16foydhiKYIdccJe
ILK22trpO20UqrXiYZLI8Pz733XtUTQ4zBxj9oE4yDMa9HFlDmVhgbbVbILiHwyS
eCytj0Ma5lpMsF8remYJ2TUIrS6ZC28Cui8i9stEBZywX3LhUkkLkX+VJMfB03yL
ZtZDpEGl0MEgYRSPIe+kstD6kRj9bCxa2BaV/nyPJjyG326epREDmpnGWa2tJ3up
Bfs8gjcRqwnUZNuhp/MhnIQsQyWt56U5bj3UnO0Nurr9rW/taDAZplLnMR/V6jKP
pieVTWAmMxqCobhj8cp3mQWv3TZAuE2mkbLjJNhkPbgwUtKWOQp6q2PbYj+/8mjE
zws4Qn87/mXaZak4woSmIJ5z7Rxu8sjAhm4lLuAD/0xyQfRX3eFE+0Y0U80KF+m2
1cqO2KdmHqAI/DuwkABH3MwAn7RKlETysaWHHTK7omiux59n07XzemuGHTa0R00l
H8xkslUHRMh8oSDvV6ePvnxXkqgjsIGgMoftnT2LsoXfH9mG068kQKvLrs7zbA+u
t2g3MlJYJjpERsBSFqKH+8uq3ECbkEqyU03/B1JnoVgZuQOFrBaVKQfsHaPZv43s
5PSzAwYxMZtLPiQM47jBxW7Lur0aPyFyWrueO1bfiyWInnAZGnqqy0M7xiQN8dax
5tD1qHZ7ykIcDwCqsDXrruArxkM6s3rZRXlwmFqUWtzCfNZQIZjDJYUI9L1Yu1Nl
/Q/ISKUsA7080Jau+KYqV6Ij/L9CzwN88K8BFTsBUO/Al1qRplBTVg+shpae3Xvi
emuJDLB8+GBLH2d6w81ySMHCqPN5pfuJ2p6zqtpMSLO81Rc8VvyYKL4LVD8SMocq
9+y+nntILUxpZ2cFLKqDL+Bwxu43Tcs4OUtzrBA46oOqTBzdThU9Jjfw8bB4Gzrs
N+TfTUqN/BFTqLKoO0UrAxbfEMgAuH9PY5sWINdN9508lvBQunWKHBFv6dpND5Ly
AhJoHYitDlHUEOQQZgpZL17oVLfniHb+WRK0rnNftlFXSXVeRG5erRGdEuaeal/c
2MAbM/nsqK1FFQAaSSthTW0RP3hKEv7h3SZk05NMJirgNWGhsIWGGv8k9qSTEUv9
n41LtJ4oQrHEeLzVGbSLvQMZ97KoIpbdf5Yfz2lTjqFwLale7NDJTmLT5+7N8ZBJ
1Ij/p4slZSVerrugaSOFgiuMrzxypmPRZdmS0k/YpeBodQH8CXCgp6c37rj+6uoh
jaUUlk37LmBuWM2zhC6HJLLvE+anjg5+opvXQRTbKR9wppxwJ6jihYO7xlsuh+Zo
4AKvj4UwUsEaahVTLXPJukQJ91DzrM0oXFNlplYAzOWwYS+ZEyHGJiEi6QSZsziz
S/sS8GQ3lMD062YB4qtY3EChHmL7lym5ahddmBII/1hg4htq2w+WESx8db6HjEIY
DRq71FSmpZ03t0SWUe8Y1vOj+cXsxvxqmnk2yW2RkYPJEY74AMwYPesCjSnoYtrJ
kbpIb6xweDVWpxxRL+8ptLCW7Rr+wvNJj0BzQMJwhGInN3ZcMr2xtpCBVZtB3+hY
gkRnGEf/kGp5fcqIS1Px5ggl+l2ZzeOpGIMmEJJJeY7a+VfTtHzhxGYKf7hc1NFR
vf6AokD2euZy5IXlEYDs+va9wo2/W4ADyX+KxzpOOOyESy3lmLbmFpLxtLUo6u5x
W4hh62eYZMVYXqQOe0BAN8S+kXCJV/2sj1VLlY42KBgmWdu/Mz+bCoJkZzSCrX/M
ODBUeK53HU/KwrGje7IVBC77AeyiGRDtYAbz+rVE9coHJBoTNPfn+hU0CtJICYwN
tbF3vrR2qBCQnXQyggWxB4USnoY203/wE3nRESO/AcFm5DHxwmebuUzD6M/uMpMg
u4/ZiYfSqlC/rgC9U1EYQqHd8cYbCYm538dSoo0E1lYsTmJMWF/oGy4mydxYY4Mc
jgO78S1UEGZCRbHY99beoIX5t6KLdChfhcvNh/YZPCU0vJKAkqZ3WHofWcV6pdQy
6aUDI1gHczqxHNQzOCdV5y8Js7zthB0ptyehTNwmA4K2v0I4MzsHWRyyg5fG2ZQw
e1tAUF9XWecCP58+nN76JhitFB6Hg7BOcR+DeZ6fQ+Xn+DdW7f8iqbivBteanFH/
llVuhGSzPYykpAQBQ+FJzaVICuRxcDQnx5oILSLzxDIgYLmOIVhWKcgKmrFMTGMQ
60Cb4yAEY2pIGIyJc9MqVZvCG0rsyHV8toBXnoy4T6zlbo7rbpvKLkm+MYYv4W6G
F1jwvFXwaK8ORMewWKZNsKXQNvRXbdSPupZKzdGpe/AIhzb8m/kMzYkMrCdfZUy4
iT0Ialx/fVrZTViKFxCfK0rEcVQbBTSi+64fcgeSGXHeSDVDkeBKhXU2UXG75UTZ
6V/Y6MhYOMkvCCfyIJfCf/VYVjcO19Oh6YXNx2VK2/nQHBTMq0cXvY28EFZXtotU
GvEia6tjuRVz6YV8HsPS9TZfZmMuPAf96+8gmWbmAVA4pPCbaywLt4TmDVNcA/IW
Lm7WT5KbffmIbGMHQNuvtIomJN5M6RWVwpcCX+rj55jDZzjis/UTmbRf5qj7xo1D
0EdAZxjwXuBqroEYkJmilbAgX+EAdRO9qZVGSDbMkDpjfY8DbGDMA0wZpcc6zkSx
JrUShIJ/xiQiY7ecapi8/KHvBMFIgLjR2NyUnyWIdN2353wupANsMfP4n7lvVHhV
YvdQ50ed7qnwwZKae7zZo7iaTt4uaK9ef5MmBWQdxVR2Yddm/LvXKjAKfX7rJaV3
3wFW5NjL0U4rDQo9uRu4hgaWFySbe3DfPY62YfcxR7v/8nIiarIcCCaM0s4VKAvq
BF2PEsvK+OA9fa0+f7YYNfQ7G2lXsJ0oXQTMGmO3SsRiniJCaihVYaUNKl1TlAlH
Q6UVyxxI1au40ANAbmjAQzikc0fd7VGTwkfsRZH2UoRluZgkBMT3r5M9LvazUelr
oOyR3buLVbDI34AVKc/gvRXjvBraX4C67Tg9K69Wnt5OtPIEhbqXail1ipB/XGNw
8OC2tckEGjE6yvXIrcAHC3w6DbbaM4419a8v8yWRmdGBMMy9UrfczD+nthgZLYZ0
XA8hMSdP4h+h3Vb0ZTeexRZTqSEHacEnzZeWdfSEwi/Ye/ikSiKV0GrNvXkLTB4K
8walhpCmFofTc76Zg1nuqrBveO37ZYlUPdE8LUkAld1nl3Bp+YiC16DWT3aD6gv7
oEBw5n7MAeta/Qy2Zj8nNVoWKj6mmoH+IYTjzrps4c5yMHZ7dcMKmcOX1VdLNTnS
D2c1Gq8gixsGUBLMuBGwjjre0J4klzmhSVGOkE7B5ngp/A9kkIZeXhAvzqElAmaL
kLMdqSFP924Q4PBYvfBPrmicO7yM19h1KuHAKtgg0RHvSQrO1uLLau4Jz04rxwYx
H9M0hkJlZ7c24zq009oUNludKteNaTv4SvD/PNq6XD7ewmbyXaHSXVp0K8SM9q1c
ngCD2a+SU5HkByJwzTRHjzYce7MyNr7wjrThVldtJmtiu349aCQKRDWr4JJ/xqDD
pZg3tZigeRgvXIMLA1HyJiF+kkkVir63IOPTxCVGo922A+JXf0mcA4iDRbgSfqTY
vuGBquE0cNgs6crOpEbwwy9i7ZsvvToANJtKQ90xL9Kcr24QNI/3XMWLX0MLxgSE
sKVfFBhDzQZzfEPIaTUFwidy64ptx4e2gS7VUt29fnWH8Mchhs63I9VB7K48PlIB
40ZnUVggBUY6u9WLmQT1c/WcR5f/jhuxbxVGSoqGWBsWKYLRB+uS8YiftYqu9r58
igv4/niUFl6FGuHcdzfxLBEFQ/0hvz1X8HYJe/HLdHTub8dsYw2T9yFVS1WA1qIy
8JBiRjV0+jvjraLiUsTbELigDCl3kGSWzxHhFtSD4out2jBNZsOC/9lcL1/0rrrI
ArnUivlZnUtT9ibvdLwHUThjP0s9VwVQ6xRu43Pu/cLBL/NsW8XVC2IhN1Ok64mA
KqcbWO3jad6iTklaXA9UmPFL0gqemYhkZEY/+ETzwFk29aC4uxF66DbLoSsK6qn2
97zsxboJiZHR3ZPWQfe4SlrB5SsX4PjZkuKezF1ImbyZeeFhCq9dygaBgHMYlQvg
6IoksTglKkduIlk8fsv6FahyJI3RD0AHMIp7pzk1+Gl86ptRlvyODwWS5Rbxh7Ws
iEn/yxLuThJXMRdkwbdr+bnnMcpFa+vR2rkzVfWxuWOwy6LkZRJfbRyoz2AN+Znq
jDW39TX0pXJcCdHmp6rc09s3V3H7k/WIvLZOsOM5iVs5EgOZry1L3S3e3werLq99
XN9Cel+Mf9axgwESmrBDkFvxtr4ePl3/WoCB5VjXzPmZnmAPm/qeHuwhgumtAXAr
RZ0jXAkolmtjLD/z1C+dYniep6OwEUx4jBxL9d17NjB6+OpNWexi4vXi0LjOsk6x
0JBSaCVVXYty5UC6fl/8f5IIBsbmO1XJr4QycjzZflhwbbQx8SfCUsiUnpsEdU5N
1+QR9l5nH0nKxfRwNwjKd0P6uBGRs0jc71lfUllNstvw02Y2rhA/UronDEdAyuLA
wI/HWvnMovbkyXzObCUVjhQpkl1ahxTGdH4bUOBJtaIUgSbSXyQNxcMqfHdxiL2M
fSm1Ew2jJh3q8ZBo3sMJ6HJZbRWMOYccHvtNBs56pdtd05F02ARavS2Wc8T4O5QI
Vg74emO6OuTV1DrjcJJKuPxDjkxJyEhjf3ZGgZvaTT+9WW6gfurni7Q4y7ZtLDUp
JchtBN2uC/iduvT7c/osgXWISUBa0hCuHRDJe6Gj9tk4NVs/nU7hkvnYfGf6TMy/
+lE3+qZExwCz1yTUog/od52VLAKBlMosM9dGtB8qs2NEFpaLNaSpCNcUngJN/KFY
LD7P8+6TEWywm1RQH6WDwTcg6ibb9xGooKwelLmZ1shm4+bcG71me+iXhIz1UOgF
UFlCn9IEXneJt65+QKsDSAUlDTDN8lww5ZCeNEXwr10dxWPQOwinWwZrjFigZ8CT
Q08fBUDQ+Jy+ue5lhszGV+9VN1DSdYWNwJ/KAXWIROGIThHn0+4ZYhdnXO7Ez+xE
jTpAAQ6ayGYr6MC+KzsrAMUA0FcXgydpezFEFUpqbAzzafpXplhgAcz36JTOuBKc
62iChP25Vzjl7JUX3YkEiJ6KSQQQRQSYVyaCOqfs6jHvBJ4zWSxi6OejOcbhn68I
oZn95efV7vQsjC9l7j3Z8c/lkb587So/9f7tSwhBl2fxh658hZsWQbfWL4nrrXfF
imlUMda0An1yV2K52MQKWMWQUHejrw8Kwlktb6vXCZEV+arpcNLM4DxuwV8M2SGr
9A8uLR5VJ/SPfZUch9+5XvzLkS510iHavfnXiNX+F15bNnTLvojipTwquirgaPYX
KvXueJITJ7EcsM/bMBduhmsDicvwL4m+DI17WuMHr+cJqvzVYhPz0ZfK/bOfjkJN
Nziq6fIamftDWmlFOztx/8b9OEGwFosbnF9FdU9kSB8L9MkPG+AzHQUBMvBAcqGP
HddeysE6Mb3D5rSBdFBb4rsPaJyK9n/nPeUDtAEB4TQCzJEPvOLWhlGH5drcjivd
MilCUO5npXDCb0lyHoTiikbG3QPR0RVQmP+wTzqwWhoxFGQ/MZCQApC6rh7rRY6U
8hUE30JRPhPntAoCFiyXxoNXrojSvwf29YoS04kjV+dCDsbczJRJMq8u8XlMVEO0
vwTXfC9nMKUdJoio/i0IKZ4cAvDQTec6ahut9cLoOeFQyh1+2hhGnhSChd435RLI
b5RMudMIUexWQKd19Se5EGeIvr/IUUZ9G5w9FRZyjJXqpRJZVkclZJFnGDlehT+M
dgEF6NpuOV0w3s5BeGZFxGvesQ2672eG43wwRD0TgUASbFp9iV+OGp6mVVvbBRqM
8juWSCUiuH5gMxqQFM1Ll4XqWKJcNcL8x+jyX2VEcW4Balv3Dz00FxVNQgkUw/V1
6ST6LYEkEAtvegTWvmnOTwETocxs+5m59gdcC8bCtENqWKgNxBS+CHPIIV41P7lX
Cx3GIgoQE8hBGzn7Tmrf1J78pylAAVukBodJhFIefrKxQD8rNOu8w1dclN0JvoTH
MBKyi1wSXDsX7zGKDbNptLoy3UK0q2cHkuI4MMtVkrXSkeYrSRsU+naoG/nctrt8
mP4plPdl8e+A6QNzaerAtxQNDW5X2YsGx4n2jF8tp476kwRiHrPbNAdGWBUdtxzC
LuCAKm8mf/sFtGyRkwZBx9votX113ychPjgS6qZUKFYrjmX7+c5/Phz7PBsmAR8D
iktTxZZUsxfpLo473Z4JEcxOZPJVGeQOfohtDJ3dqAoLO99JCJrIOCnpe7ivd2Bx
FPxhQLg7qNHaucj5Saqagf+g/FlQQL7FnNvQvpntpl4rTGKo8EQMKIj9dK8rrJ3/
9qrAWic7MjanPO9Jpezm2XgA8xdj9I46je8H7lYBn26oGeD6iQ4rf7eCxz8qyJrW
d9b/CR6EySDFicaG/u33AvUa4AEaIruDvakEzFRTl7WT1L61BugjdXS4GesQcSeS
ozxMT2h8/4cJLsX2euxbccqgCtLS9JhOC3BBvlTb7jcTZkzbkh6NnU0F6PRQWMmv
AXpxY1VL2oGeLn4AQLk//Wp97PX7VTyw6rV+kTp72BoyVaYtsv35fnkDKbSRUkyM
izl7rvh3Z/DscmRwqsgUJqxbKta+EYhMh1sQx4mRTsD490N/ssgiFREXknQkDNYF
CusqrYqzNiFqXKekGCBtdOm2wQkaCGaIpb8rHOTuJ3Dqj7/rzN0EEwVFKRtmvhAK
pGPGwV625s6OON47yvA4XArxeQKlYagBHjvCA6rQ/A7q1+nYRL7DKWujypEacfkM
Vfpww+srLWvBkGCkgDdEgFgOjMcWVqf2mTM9elCyAq4acjWsI13S4BnyUFV0uVqT
uT5jncAs/Ll867b0lcAwLYthzAcsAoV8QBfLH+kNsNwr5l5G7FS+tGtAzS+/ymWj
r2GeyGArEwTEAqOQ09mVxSj77jPPPH5i2BP6oTXgFWn9AJ3Vg/CVhI48BQztgrGp
/zte4sd0iF+tVvdcTAsb0RlBhX6IBWOgCGJ3zcv8QkiO83sHqQXxNf8jSfQ24t/8
GKYcVMF6vCB22buPR4Zpx/WALZs57fFUX+NtbIfsX9MTmPrrru8QMwBGpwiwXmRu
UL3UARfv849PUXrMNPD3VRJ+6emZ+Wg0Rfk+gnK3C7hsjmUnKhIAz6/u1rGaaQ74
nZEfJwLlqQ3vNMwRCNZEUxMjLJPUAZpmshcvhHOYQiJ9mRQ4GMLfG+EU/64sQJJs
vIhm2jRpFgxQrOipvEBVqhRdOmOvSCQTDG+smrzKKqxLd8Tn2zM5KttryrLxlIB4
dfnsZofOoVHbV5/dChVkRKwd/tsDLMRYJKl4JeHAZ/wp5qFbUuSPGdDkC0OmNR9I
tCZAo7YY9RXPlnHDqmNYiu2mpRV/VTPV61uJRwHnYNY+YmwAq3r1Idc+J/OSs5BQ
GxjoiLxMxiOSs86/klJH9ajWY87JFjVu42HnFn1l6pr3jg/61YTh0ZadhazWXerO
mAmiwOF2+Ztx4aFrje0GjFdVD2lGnc3y1mFxIepO5ZtxcPbm9Fv0CTLX1SR/zJ2E
SE+a+l0FLp4Effli+Drru9beeVRLi0Q9W35X1t9X9QNXYDGKHMBq3SNTFZc23Cdi
tUp2U2GPFznVp+b2Slv3zUmRok104kPVdH/NTyQQ9jgLth6zepIx+wgdcvCop6Oz
6wD+68zrUUcvnPq8Xi4QDy/BFZyWJgG4KESNnRfTMPtn0+MgxGT4SxTtOSx4iHWS
a+Vi3klSzVurQfsnC5O6TKasD9vlv42zg3BMShJByPHNGclf4kDeVl4TECbrpRz6
YnWq3sYBuu69KEbYcnhO8bAUAqHGUMIGm4Zr0QcUfV5ZoNaTAtsilG94T9ULuy3/
gnAPWBMrkDpptBLmg/Otga5vK7x6jcCpykCv1KLwmmwkiol9pz73Uj8NUQa9TFY6
0PxNpeEzPZ1+IlW+v3NtGD9n/2E42CiGtKVuQ28QqVZFmunB8DM6EyC4NtY1X6BZ
dOe6ShaehGhPIRHCLYRhB8To3AbbgdA5iEScSNL0slyqtya5S9cL49+XwBUEbSkW
OfSP4zjzmy67oaNtY2kwu7YW4LdNBIxiO6s/VqeB9J/gruHiUenKeLd1bSZOmkqL
Cm2uNXJeWTDjw1ihcpvaW/BnDFXM0+xSJxXLtATijeNQzC7UX3ze1YjjGD9D90cD
lKKzf2RlYzXdFtFw20cdBQL4KZitBT8OcYwG9b+nnO+9h6yGoAe0tZUup1oQE7Ei
gPLqEbzZoXg5oscvgI5s02IM0q1CFzfgQGHLHiochz8YD6BemQu07IGhd2ooc4UW
iqVdo2MaWBhHblum62Grro9ponQO9Z1+o+WDLRytOtgc/KV4/YzqCXv5kSVCmyyx
OVkbWLxyw3pZtUC5pFs088DTChTCnCf2I7guXenZeRvhnfFHjme/sW9VJUDY6crJ
PkZ6H2Oq8hNsPUMZ8djjcJ9o2gEyfG/TqJzhuDhi+OVXlX5QdM3Ts8qrsl3DNeiq
F8o+IxbFOdP9gS1HDvK2vHddNXuf7oNHScaJspNm/M0/rLJ0Qz4Gs+Of/UvvFFmy
OybDaKBtXs1wWzzKL4nVA7sflf5mWgdYgXMnXk2mVV4xuOUClNiPLLCoNFiws/yk
ncHSQG/Rl4p5+ykOm5zps9xF7nkJbMsJM5fS++ZhuiyKjqjTNuZ6ZIKFIx1aIfge
323SpeGK7HgT5bVJrKjeMmYsCyQOFjZl1Nc32VZHpF1hKNgdSXhrJ4thFTczoc4C
ronQBIFvCquvwR92AHpNjV6hJAc/XvwR6xZP6XwAZMZFC90zAckJuszHy97bQKKT
lEDJZGAq7a3GAIsT7Ec3x0Futtlwop3kWWcI5dH6IzhouifeDmfvsjbQc7HIt6zs
bTQDueeRWJw/7CvVFo6JTWw3iqFmhWR1gi8H1r/aObFBzZiluyqrqfX5763Xw0qn
u33af2V5nlLLpGhy7cuIsqsmPD7lFgbNd5BMuFCf5//YZPmVsHv/syiIHw8KEsah
N3T88Bhj015Wi020atscgHiMdAbRtjDXGOU1suQUhH1xHSJ/tFE3ACLgVUPhskga
kYey6taziD6wWB1NfVWKDVnSWStYHs6V0FmD2b2fKCW9j/euIFtj0qOD6EczxC9C
eswic89kiQL7yOwiwG4eZEy7FCK6E+2RyW6QFtmLA8x1NH8tcDgop7HqIb+LwaLd
n4fV8ySxcyBgSOiwkPEnSnrvwsLoeWxcDb7Qzozp0mhx3vkBGKPZhYEGQkNrubOF
Z9OS08MiL8EFHuRrLnqYEp3UozxfjHw9CSCrT3HVvcabJd03lBSUf1F0pJo+Thzp
j719xRjQUi+cPdyhMh0on2s4G66SSKPU6h5kXo+HojjDGgIO94l3ROnZMNtDM3mW
Vs2xZDZBqpGjpEEy50B/Ecp4UqHdWSOKlvqjc8KC5k9QR7zTGDFIQ1CevbgFAM3p
C/rwvV3+/iNsXzoq33RdvCKx1ElB70GzPXwpTW50HoxknhbduM40oka/hVgIeynr
l40haA8MPHdGEuTkDWvzIn8hnAdv9EDbtnc/CU9TrDSbfAu3h7ZkYYXbRn6Xp8JA
tIKK9xZdRidINl2s+BaUiUDDuu+DNSzn2zHtueEa1eR6Ngv14ysm5PeFh6o2qDPA
eAK2zjaplbslDPNVL/QP8XyA2oF0WEBe/G3ecdYATBqji/zPeuHuqpwoYI6wXgy+
UvAt481OFcBliYi8jTvstw9jWKccFu/STCIIi5ry3l/XtKpZvIwQLE4yrpArP1+N
WvGvs5KfQ+SRPaSyeWBYH54ML1NRLMyLtpQEZ/aWkZAJtsakv5cKZV1Z8DjlUhai
uMWen5qPxoNwfBg0o/cBnPIhM3ADOhbmbtp/MXok2edQHvgDG5hGIhw3QMUPw/6X
JQmOAVS+zg4RmJaOAS5zVUZKZRYOMaaaL/1U8cVp42SwntZLkkEFu3sGwf1glTyp
ChKEf28CMX0YO7muT7jaQXo+sWrNqMWJAlQb7VeE1Ssh1AOIh8Qhle8+bli14TYf
Yooa6PzM6+zQxjy8LJKidIK+V9CApdZeHf9pRDiQfPrkTyRw9KHafvc24cq9x/d7
H0Lirh+pCyjZC2/FyeNs056dn4bVFWsfbTS2feAc4qsu8nzKKBbLYPYvpfQXeLwO
nRYHFL7w88RUXGT7jhSh9zAgwhvM6XOZxx+wh/Qy/wNF6815BGFN2NQ9drYrgsP5
uUSreBxHnaFqfOc2KO6p3JRl1rmqbGhkg6w1/wl5EZBPUnB+X6BACBe3t9aegIsl
J7HHyyApzYLOrkk+gyGulLsn/GbTGz+FRkR0Kqf+Ll3bB1PIPQlI0vwAZ89oR9BK
hA/ISv2izTJgZRpKYFlUTmlDW0Y+dk9amA8zag9keYHJHxidEqkqXmGBsdd3l7dJ
Gm2rp8GluprTvBr12V8k7JbWu02beXTvEwdyAKQwVl9e4zPEshBIL+K086JJwvR+
kCiPYNiLRL7kPPs3dUuxDmdt2aa2qCBTo+sHltKikiOl9mNQwyDsiaYXhmX1Tsqk
V0f2swjrgWvb1D3wfiJoCcmyvbf6sTq17dKwGmBfRamUbPx5mkzXU15WEuU60a5A
7XF+UYy4kD4vKuikXe8KZvB4wtECYWawVGZUzrqarblbfBMYN6p0v/W/VJ29+hyI
Ph5G1rYWcpysuBw8ifTbaviv9TXy9Zu61iFkdDME20UESoTpIdUBPR4rfZ7Gfl0S
pXPekTgIN05NAmrbBnEvpwf/atYaEO6DPrg4VqTeNLACb909sWONxh95zOXEZOrg
drWWT5SPvfEk97TuERMisK/fnVuDtwCK414wMa1p3M2ANDrUndvh66cJUAN2vR0I
THTWiEJI9ciQb1KtloSyJbORHlOFQbTCElpM+2yhDIgG/OThwSHQt68FTUHz8Hzv
bip4PZbi6BUPzgjbeq8YBLOTXglQIoYt89D5ihWapHYnvA14DtJZPHFQuAKzqNI5
J4S5aqLbl0yakp9pH6KXotUFnwXWml8gb3rGextVf+T0t/OScDVK2FaCw3ldXZ4z
ibCoUV5Sxzadx4d1A4GGPH5QnM82EdFBQ7xSc0uoak0G0RgFJj/RRl4x/i6atyXn
gf+FnbgU5tJRc/vKDRKvkMy+gA5PcTZE2tTSdy7HL7VDvZiXo24nV5RK7mQcuQ2/
BZ+qBkwc60xfWtef7AZZC3JKefIj2xfSRGp4xgoLCFNdKJnRN1fUvwsdmv+tQVH4
ryPxE2iuQC4wTMHwAdfPlInJYyrlXGOGUs2OFujyfgMNMXPxdEWvOfOEPXXVREyn
3gpkF4X4PXsIi/L6NDy22X8/BYbL5IyNHV7YaO6+3Y2QkOB/Xv/PGFhIlQ8P4XiX
1QUMBfgGU0YG7QqFoRHOOjvDTZNop5G7fc6K56ryc6/Tp+iASXVX5huc71emiOpW
W5ddsLDd46VvDCY1j6eM2H/D2QhTWRCJTd1wsS0XyO/HeysHMyUY95bNC+YFXPEh
KCmp17esKuxbBXnnuda3Q1pItLKDI/W+LoVUdJ+7yoTqegP4NoWU4dH0o/CVNOs8
648eKaNl/GHbwpnKCIT60omKzOly4MVaBQeoaTqzHzHlsPqXyki47Xtz8TwFY7xp
0cVtvXuJnnFQahJgEHZLKv5OQ6pPO6EwZvezO/ga0fdWtKQmvaUlpI57dpHm6Jy5
o1/3gNkQimTlySFuxOsRut4k1E3j1e8YHxYI23I1wNM4INDTy/BZ3ASLjEJVbJZm
IPh6BYu6Jf5MpDuag933GhiARQCdfy1Kvk8n38jOmA3lvLoAMIAS4pqvKqcldHLu
5eHzDPJ9Dph8QzAlukmxblQnpj0VsVKS4IE8AnTGr2nAWBa1dtPHGlfLjQo4H5/j
9X6J8iCDf2zaACdTtfR35WIJzDmGH+UL7pJTXJgydc250DzIPJOHx0HK8ppJ5BWA
YePRSQs0vLBKsqfBkqXTcvVDHSAE2w0Vn0NnqxB1pNmP+m/Xj86pEuTwU1LN9d5U
xu2l+6YT3wI+szSjDWCObNPQ9Cmb/BSgK2UHpi2wrh6f92rPY0FPCfgJRF3B9Lnn
3No0Y75yMxbx0SGHHs3AIALUXf+FUzQhxclrXTXfUKW91CXETpzY4Yq0TfqdtHak
0gLmaiD3iPA8L92GOBxFKzdobptv+ciiI6MjqLgpCddSWvMYyIcQlfCcRIgJEPdG
Mmt3Gm1NwfHKUHH9NA5vmhd9TRmpZug/75ccpi7MOQGr1mH+nwEH6zTP1jwfYmyb
yKZ2QQXMoP7qXEBtH4dkENReW/zZNt/mJ6f0Q5VMa5vReh/1+TpqKJJYJuvfoPXr
JV94BwOeNYK38i3viNnCOnU18xsZn8kg+paqeSZter9TAy5EKiu0DN4W2ffs32DI
YrAnEo9OXIztkvW73YpIVEy1J9N5vUy+nkftzThF7VsdklM+ZEUf69nLANVrNX5p
2CqPGjlWoXuHarreJwzsCOGMlIB/vxJkRgBPVSZi4dMsLBn7b9HrfuNWqwdyN0eZ
9J0/kAuZuhkzW9++lwWiqDuXUq+b46USPazyz2QRFNtqX3/jnU8A0h+UPcUAUCu9
LtK4jVH9+biMeHuyude3WmCe7EAvdFGCO7cXOuNOvhe+akykvPaIoiOrhLPYJ7HY
e+5zEpxNnnrB9wZqiTqVfQ2lTdq5ymXvhulgB3ltNlpjmFtwpo8em+9DTCeYa/ql
e2zzrOmwmqK7w1Gsq2ukw6YsckvA07MJ3SoIe3vMVLAl3ynhH6ppguTnDeMrFSdC
xLgDZkvrTiWb4Nl3U+LDL1YmZNa198Gi+FxEhPv88GDWltXauoc0PTozXy+opmws
OtPbHGV+XlH4a/NH1mslBEgYCxaA84Qhyy4v0NV9RwYeFNwHtEKS/3pAcG/Q7Wbo
2ZMFNmWExiDp4gdBPllEixP9wssYgDx/4farIIxEx7tOK/FteXT2/8NJkUfXC9ah
K2pUi/8H29yXXSlYfLEGHfb0RlZWMNgeKy/VQgbDZFFkBfzlAL38p94U5wb3wFt3
nJSmnwP2D8CxAomnBWqhmz3bXPLggdS9hPq+Twys/TcZjrDXkgvkK3rILxmYS2Ra
vCEsmbdhHhi1D+m8wLl7hrDsyXYsksHVScmWmRYl9fZevZcYu2iK6O6vgwBF0Ebw
LbX2VYNv0CZPbzJ19f6bYXTyq6+NvszCbmcwC7XNtHfNBZmSIIkJ53PqtQm1+Uan
sjlh+KYtuXroFGp37ZJnqyCs5pwxxxg471AgkMVFZVxSYlNfRdC3ClDNCaTddwfJ
ZO8wvmKDDe8iWPwtX4g76dGFXzZtG+TBN/ug2HDxZuQrRcmo8mDzFepALwyW3G1k
M6gm3pcYYyDEPInrat2yhcgnQD/Yr9L3OjBFEw+Ag9PVjqXWFdlofdE+8nS/IFDv
U/bSo1Thl59/1RdKKlMBsC9FzYuw4L4TpYiA0y6Iny0AFq71S8cEryoxY+0EXBDg
ybTaftKh/ZJVUuCa6OyhNPsKDFYV/By+5kt5QvxOk1SoZkg3O69QZddQqdHbQQoV
m+K/OioW+K+7jYMd5pzDtP0ei7gv6nBarbLi9bYcqrrTL8o7p2Pgp7+qVK2DXp5g
xP0xxTrN9aZbKu4kmljralqdmShJqwpXUSx5hKyeamu6KTkhAjYF/9KX2uKrBNS+
S1RmmS8A5DJg0s6wxhfFv35WPhRkuZPaIvh3Di/oE0mpTt7K94PPshSqxIN+eoxP
I4sq4uZLliA28MvNM/nFjUIHVd1J4AiYWdpaBSzOIq/1w6p95JrmSaYei9OS+Cou
+wSaUVHLKszeWAwBaHC5rY7/hBodGidN9IUov4ZrA+IARc91u1H7rwG8NWzXmrkx
NRWvjzY/wkXbxwYIthJ8EDkajuLxIeGigAO8pJiQ4Bfum337HAiu03wO5mpl0Siu
e6Od/fBtZTRl8ZrXWUMM//tnbv3xLfICNqo4HGT1+c2J5GPkUuny0aghwAlmWJ7J
IgU6RallFBLWOeSIdBIlrp4cyqNncayuCQKqmhqpku81JfHV6PtTBMQyuDnu7V3+
CeC/efB+WFAYaqP4Ljqy404YCaLhJNu++RgG4ahYbygPenKyW6v/zDwQ81Ze8NOi
op3P9N9Xs/D2qHzu6fjUxOmTGmiBmc2YB3bYfQ4RV+5JNnUoLu/vOnAtdJT8CXA5
AItdBq0vgdWx45MXgYopuAeu7LUHq390WKkqIge+EWLsZEQx2ciDXtnVaiwaskHI
aWkwqXCqARFUyHpJtJm17imIMVsIMZHZiTrLM/Hx5xyseRgVk1N7PPn7dPME7G/m
yzJMH3r4kFV9KILfFNF0SUNF4HRJxHKstMV0kDMkvuJELIwThfZiMCbZL0NWYIBr
ttI//g8NCDtpQC/7bORrWW3R5Xy6s82heZkUz7ZFm50YtaOwG3hfmWdCqNEKKxE5
x8iMIO7SHBnGXivBej8os1nGvZnhh0MG3Tt5bnBbh5U8/Qk37n1cv+EbYsYxVong
M1OMT+QW0nlECppFIZsZHQ/qbDQRok4Cxd9HgiPubTJq/rQDIQbK6BrL7PwyqlW0
wQJ0qCwL3nSvnWoTmX1AR9wgZ5KUJDXRTlxAEIZchtdO/XSKuBWfL/V/w6eVpLd6
sG39pnD4GT2ZgzyD/n7x0+Y5jL0IWhnfEYW8McWjKiAPQoqWReWY7ePOLu3Lrkj7
b8mjRgAIDkIc6f4k9AEJGjbxoN+i8xGp6cGuGLj65m4TSc6Jo4GcRzpsGrsz/VaX
YmdDyDzzcIpSnv/9Hqchh/7mD/Qogfqs1y1131p6V0DTf5AIzaqX2INC4OYKZA+7
yu2Qpv2rWuokwyFh/gZbtAZ25QX0UXBnfNt2mT5pNaX/jD6yPR2nTKjFI0nv2bh+
6VfnbhEVOX1nMNNK/e6Ydd/VX205nok8MyNcKdcJd6IeCK0rG5oIPZYkf0FxaXA0
tPLUg6PD6vCBx+4yR0UjuJTDCQOrYGROnNXOYt/HmJBCnD1yoRNlls0LgUq1RP8j
Aw+OD4fhsVta6v+clzTo6XKypC2hfEzttdCuHyC02l8uAeRMdszHR5oGa1D4LR9M
+cDfj5qIZCMAxL0eLUadANgTuOkspUKfca0hs7wOHRZ7cIdsfX8rg0T+v0Q8Ikjq
YSoLRKeVQvq0e2EXHCR9r/iwXBWbtWz4hr9JQKEOe/4ujW+kq4dF4fnLx3ExAXC+
ejPpwaYQ67RXteOn9s+haDoW3jlnlYrd9c33RczVcEMN/LineTeXyWbno44rTxh2
zKsYK0LYMjNdSxrdJUqG5zq4cwivz0mu8kFfYzX03Ugt6i6U0tJ6sfgekf3qsTXF
hnMzA756bekhIONsIUVzJNMr/VfNeiqOL/pyHXkkJxpVAkPwEMlJijeMKk65g2bS
3un4l+W49OBhgQRy7WzcX3/Qt7SRPaUyM55I0Hg/397i7LG+R+fj9/0+yudcpc5L
agkv86n0rAs5h9jjB/v3eyyM1+zPomV2HZF+qrZvoSS5PNyOTbshSLxM7rmVHTMN
YVt8EQJg8KuWyRH3bqf2w/Z70Un8ID6GE7joeiEJkrNEPpgbghO5wSvgWncRv8zE
rUK0IihZ9TFsIwjOXe056x4zUJksnIeoubnJ5AfQz1L5Erf3Bj3IYvXRja6vTvoh
+tx/fogw7bm7YS8z3Os+hYMmm2L+RGs8TxIcqfq7kl+iMJ/ot4tm8/4R6x3FGQBv
AlZ47WJn7zpNs/jwdhqAq6ciU2mKZtUFGwCCXPtTw4a0k/ZmKA++2XCpiovN4kvK
L5y0eAKxDiLFvs7eFHosb2/1Oy0o7nsYokE5viBjya/Cf6Ba/vQ0mA6PWQTpS2H7
SMjEKb219z2WBR32/gv3XuCAAHGELyqekSudiYJPI+AgkA7RSteBjvoxY1EJeAwf
r3bNqY9bip3e+5zoaD8g2foOF3YtQ7R2YTAotCgSwufnV+8V+o9bNLblvrXCwn6b
962ronXgc3811m8tnlUO1yW4OeK7RzijWJr1ZaOl3nsAXQ4S8qLChqexfqt7wcuQ
9G69i8OVuBwp/e21d0UfJfA15djkK6y0PkfjwHA14eUtZz4VegkBRqABSqrhHZnn
I+Pp3+RjoK/2in9nkEd5OScrSN7DVPF/0/eaEAWhbHtqNWAfBtmWWyQkgWPUBH2X
2ghO8cB0isJu0aM6/p9EkAESEmup/dmjgJLWykQNW9CgZyVkc63FkqC2y44/NpTp
eeXK7tdPl8nPX7mFy3PAP58knoBg53Qhik68oEU0RCv6I0Ny6AYDPi6cVYzaGWgk
dlGDifuoXIIX4s3bc8xPdjaQ/pkE8qJ+R5cJf9VI4h+yKtlRcj7AIduH7p1beb4C
gCZj+lHdNyhtRwToPV+vhkDR4uYA6SsAnpQc+AVRPPdLX2Wl4lZ5qJrTZZi+LJjJ
QYLSSKpuuK93f87oznvxkuWdMKZQK6d+FM23w3Nn5inCFNi72dqfZoDsV1Avhm9U
HByo48x/QUBxULlxbNdz6pjT8tmDxRf7+eSoP0ZRbhSqnRwjBARa6C3xpTLK1dGX
IbTrR+BZHfMjqu0yQ2qx7igljzM5m32T3ZSlzpih1KtrY6K2GpcsycaKW6ln5txl
P0rBMSwAoZIdgepKnUCUrHSiN23smOboRsAYpcJ1Zy3K7tPAOgFbNlpJzxBy5eju
6AavJbRKki+qPjQsFHzHmTTN9YsjK318kQccyWkGURfTW9A+U0B3tpBHFV0ZY91O
Ds9QO6FAnTZmT0PFj5P/t6uTM6Yd+GTSRT3FdsV3qcZSjwL3FMVBKC1R9nXTqOoI
O6YZd70a1gTICqhkpKZGWlChpz+LV9toL9h7SFjtkQu9rutLNFZxP27LFM29/txy
64LXuxaw7BOklLqeZ6JgKjuAgfYdMLnq/ih92p5UqQ6Bz6ASY3Yk8OoaZfvuEWFZ
a73WJAIiUk/r7pVS4CZOYA7Kxf7PkPRyaUxdrKsOrcfvMLzJBEXtYPkpLN7ZNGMB
horM9abvN5aPzyuNtiZficApD2UtUabjMz8tVCfjmd5I5wwq6ZBT2Z0h6KI14VAy
Ncmsz4LLxVTOk4u0+ehyrujK70e+22nxbLs1M7SUIu/VzAStht5T8Y3x12o//O9t
UCHxSs72/C/GcIrmD3MpJwlC8i4mIin04DcQDpVuDlTcfFmvQrZOAmio/vqoLaVi
RYO1AhGOZsj1UD3ruVu/atNiIZDP1P9tW6IcKEvDHeMHF4u1Yj5boZjsWmFa3ero
cigC+e/whbPthLIrxzmjxbxnCfRIbIvUYRBRWfR7VVoqdV8B3TdH/7pwoPhocmwE
Cqym/Bn1Va+snSz8Q+/cmAymtIPkWSe4esSKPMBRgEOHqO4vEai1GZ8myA1rUna7
84JGqkpoAMVmuW1BI2yRrd7xnqNaKAqg4MRBzshABG0xwifjyawEQ5LiAGQ6u9PU
3nDHT5LPipWFdpvzyP1zjWDzcok6uMzrs5v1PmpznjSxVRXiRWLrfBlfwEJd/YRb
YYCHLMwC/KYxsp+TvTG08SZY+CvgFdQzTh5E8AhEaZqVpLlO4famwRN9DCyoLamX
AuY0tU7jw07TX2m+vgq0d5iUhCGzafmgdD85FPB4ZCpKYdHotf1K4jHmQv8bFHwR
1niQeOQ0VoksDkHh1k4iwGFoQ3wZ6Mx0TbsbQny/48VjbAKsYSc8c3Q4Y3HArYzQ
xdUlt8xWbnr8lB05wcFM0M9lgWYtHvwB5Xg4pGZK41m28C+1zd6nMZQpw0gGyq4i
4dDc7gCaRmk8etlcFt0O4XHn5mAFTg5nmG1R5m3N2gQYrLzxy6k3guKqqqZH8E9H
stQKjms9FprxKImlLikI/aw/13bv263raGoHQBW7wsKLIgndBKIksKFAF1kZM1AY
8qZdkS4bi7Sw173hqeLYcPpo1BZ581lMwngy6YtWMp9Gy+GOYPSapq0md8dM59HW
6GIg2qqHilXfT9r34CEeshEKVA51LsoDghQc5soPMg59sVauglayxfgW528YvrSs
m/wNtKIrSrCv4EsjBQYjzWjIF02MQ+DEIjtFtnvnTtujlOOlQLpi7zHGuC3Po7sm
W5yY/0HNmr+18T9ObJlwqi50tkOnjLkYm0g/8Y/EdkdHHs33oXxZ6brRqEQBgjGJ
Cs4ap1C+LvdAGg8/zPv5jPqeHTMHL0eCHbvmEIdZj7fkNd/lZdDyIJQdaonU9DHP
kyUtqsmYSjde2mZgkc8ABDdT5A+UW1xE2Zf34FdzU+g8udwDTzqlEvUIpTNI98b2
eKDuIlXPWIRZJUSUcFaoYhox459tjOkrr2OyVb3nvyeE39J50zjpvj/WSc2NuX8o
tfcV8EEvwu1LXKiRxHgnMCgysSKyjegsWlhIfeErG+PQM5eZLVoHlX126RQpXfX3
bkTieHMlPJ+SwpbF5PLIATiPjwhzuuIGf1DBw5um+FCxWBuRZuE022IaCXH+aleJ
a63xQvJu+LOgRUM0wKequKTJbgYqXRe/aWyaDu/8KQSBPvugnwjRuqOOaZBwKsb0
Zs6ppU2Ph+G7W2SqUkD4/+wZiIJiouU+7oqNHhrG4uZBPrCTKvDSRAdJxuTxhQ9R
fecK88S/1ExYjzGBIiBP0YzQE1P2Vbd5ONhg543gtTBTw8OCoG3jlFKQlB/YWctv
s3VqGzDCaXEGjI1GsDLN1fcHH+/8vMQzFvOb6/Zdw+d9JEuRJJZeDN9h5GXPCdhI
XPq/IsvZXgHobB7DziuQDlHFY+KcA10yG9PF/toTCJvGPnILpOuuo+wgtYyf7KnJ
KFdGK76b54EetjL1l9FvaqQn45caJiorsORjS/00npPtHFvJUcITlKwfmC6/UCwz
CT2t4ex/eeL8cCXPOTn+lW0JzDgqdAAqOeI4LYEUmWLFtadhKFpPRdUS8P0HvDMz
PxdyvvRvBRhIZxa7RGglHEINqcZ4VTyzGtl+IR2BMHKkrSR7Be21coq/ji89/kQv
gds29Vb6B7GPbK/Yn3Kih6ztUEMmZrz15kHKtnUifnGpWMvh3v48TYn4crKUgEg+
BrO/JeczzAp3WLAv+F8E2f4evcaLMP7MWylD2dU7yp80tqxtFZqh05zH2YSl9uwo
jRJzwNK7mmp+tPZFJ1wyLV3JDbBmY09v9fU1i+d0k7I5xPPhuIIyylhPgLoADtB7
0MconfxKA/mvuVKiStpqXvpuUEGzDkWcZ0vZSStwc5ETiAXj/+VyAmR5/R70t2QZ
7CyT/BytW0i23hK/XzXgJpTieb7vXs+g6ynhfuwXBet2/m9Wz2sf83HMLrV9zyF6
SooJU6R7HSBYrSv/rwnAfvGpo00ShyFER9TeuksqbA+kjI87HgS26tAOI+Osdb79
QIunh50oR+31c+HmlTi/R6Ws8zgXAjStbKzl+pqW20+sAFYCqDq9QcarkDEXMA0V
jL2PpdANHvNcViKk+787NJPUvwEULY2PNZ1CscjVqyUbbvy3/lDEolLmNTNVzR7j
XZmbRTbLV4olIcqfYBjOTooM04u254ehdutFjjvK56jGX55EQE+rIELC6YINorba
3HmSFZUUpl/OnQF5heZtoyucFR4+3DK21hyd46g5Uy+c3kSG30g/I7Kskf/21Ys6
1M7cfNA4xv4rLOZe4bwtcUWc+tjj2EZDU8989OpBzwY/2JyTC3JCOnS8QKh0iIWM
wxwmu3LtCWMtj1flT06OCqGO1+IZOtPlkD/vmT6Woey9hd21hUHVtEGUG5JqEWJN
IAs48IO0F9sWNfO9LpyJWQ7pu14EdYW8FpnhbJGOpBdPtnIBj5XWvcrTzqWPToXo
D3R8oEv7PPk9jEnAubudzbp2ja+nnjjK1K7qTSETV7DYvnqX7y6/9zXV599BXNk7
1lyotp8IJjQq6dcl5QalfiE0bXKwUX/q4HkjZKBJQ5B6M3WFRAe9REQbbY4fublx
6evcVGaPMMGnPRiDEJqZ3wDvgLORfNGu3e7+xr/CLe1HJP6iTuPVRFFuu6/snDAK
YveIlLJ860Rh38mGUcFIUvDX4SKV9mLZhOAAsPfbuweYvKbWPZixIa5NYwJfmRm5
93RGpascGGPjW9rDWSZFxptOfpNa/uRX0r2tM7nHaNRTlptrjGeKIqKeFRAL/S+e
EpVvJgzaDebRsc1k8i69CpYkhZTHiN4Vicge9OLag5nZDBypjzfEETGDleABj1VX
++Fx4h+oCSxdtZrmahLCfu4645lpnaU1QFUH0lWpdGl0+4P7QhriLJx+727hrvU1
RCvt3xE6CyrlXy5arfdC3/jQjbr2fukb/w33nVVGl28DrfoGUBIxP6rRkSufM1Xp
xmTlgt+Dkd4Dcf3vgVNlk8WjEnmpscoZ6hLbIGLOYA+8Lo8HQAWTzMHCs4FOEvPA
l81lggxZg08rMS9jm/GmQVsCERxSpJrNxIploU4xxVlfCsl/UKOCEmT+pslR6iPH
nlrCQPbvlSbAX4Ljwmb7a2U96DbMAFsiXXBnGgPKaJ3eAN27MeWgPAIuBACIu331
cCSqj8ygt6hY40R5tMmeu3UL14EeqeL7dXLu0ijVm+DtTyAo3hj/d5byhHia8hsV
Yw5v3KwNGieFb1Izw55wNIFfDMScqkrzejDg9WMqnVkKp/om3HiZYMRZDJmIL/FE
LzHrW8BkDVRsb5sBcHbV8iSSzgy92gX2YoB4Sr7pEYzuF7f8VIKaImCdAQZi0tus
Yb6UwbThLmtFoGR0W8y5YL20XZe6FSx7cxcqcATmCFvGROBRxgsbdoIMHi5Y2B4I
ETX0CeK5ohSJd3YFX+LbTEZkRSU50gtYIp1AQyUPkgcApCypb+cwBBgdD5xS6ci8
L9AmaJvJGpkO3NbyxeqAHbi0S20QbxAV/0QUZON6OJMlScwSVBMPc93bnFGVLKLO
/LOwwBJFmOLjwCerK5RKhotSXzY1q3c9g+KvTkLM1mM4k5C/KzeRcE9KIOnh+O4F
JDzhDHjOOU/tNbDJR8gdpzohHlQ3JtlRHO22RvJwaY/JO78apKWOSOU2kFDfeT+o
pHFZiPgWC4OR600/IdvU8NiAU8Z6izWD8NgY1yPYudsQQKqXI14Nvgo6yVXDOY2C
fNJ0NjT7arNwZLDbBUAOAmS4fPyxrOdg7y8ZUD7Yi9gHxNZweJEMYCc+kTEblLyH
fwlQXSJayg3Avde456XJyqTX1ndSBbq2riLZXvV9BWcHXjGnNcLhAseAsNEbndak
7vCj1nQpSzyW3r0HdEh+qhELbWT91Smq7GHCpwm+AraQ4W8GV95h7decxj/IUnOS
EhT3yRXkjAUO/dUYljDVQc7zeFgyZGzUKxQQ5DmTqaLUvGm5V4Gxlu0/CDAmYcFc
yqZSke8uKUIoMTdQMexZ8gQQZyPeBzJV1WK5vzDByjIWmqHkVxZtxZW1wCyggS+a
4/VLyjt9KVYBlQbXuLLz/oeqauEEeoIEU8pa+hFNQ/lJbd5RUTIKYdKiwKH3ieu8
2Cb8AaIxbnQnFs1I05uolFcW3z4rPpcJnU5b3oHK2TVkcVoiBXhS+kWIOgj9noQw
QaWNFyeTFSIi4r97RaMjzCAeUoLwlMGTUleZQPpButGmd5lnzHLTlV5uofArZLCP
pIV0Had1NyzJ2RCbZpezjwsIAytJcRJBLQxmyGsZ82dVtLB3CBY81HZduFNVky7D
Z8rn3ZUtV0R/WrTBuLRdwEqzLkHd25VDvPmZ1CXfNYGmWh4zfT2xyCDjsYj4rz1U
KJnZCSFSkydvL0UOaxAZ8E9mA4ZKWbG3whCvvCWmctqg2qWYiNILrvqTRB6tnbsU
gqvC7ER4JDke070RFLqpa+COxZy19BjUrDLUYe7ce88cXnhJ21xj+eNW2X6CyyKI
8XJ7oqZGBa+V92U0m9t7hPSQBqGF0JLfUjrBJiiSZyDyMWjFmmX6DFpWQNSYrPd6
7pGHC8zGP/q6hCGGtbKNKc7zH5E6xKjwu5spBBvvUT7g7lC53/8+FOg91aacTFJG
MgIg4G3VdB3lg3mHEyFZakMVrCqQHdYMKwUVwly/Ogg8YGIRYD+xNYUORYN77Phf
6xII/YhTh09O0swl7q3NQoRjl1xnyhcpca30EEmneR3zQV7oZi/cVIHjNskUisBh
ILqjLKikmpQiJ6KCRNYPXctUSujin9IJUmAAPiE8NvK7mSdBy0BfNpv3sLplTbx4
O68MS1oQRe5LlWweL6eLJNZI1I1z0pQ4W9sKVN3eBZnjLbr+3jVo32A6Gn6YeBEo
k84EQP93vS8R/d578C42tek+7zlURLIzOZXtE3ePwl5TNVcbYye8A1IZx5AqqeLv
M3amMj0BAlvN0dYS7NO1tMPsxTspPvtkp13CmJQxeTNv7zwuGOne8C+LsAt7xUQK
VcGyxNRjrNyF5dBRyFnqmGQ7MDzAnPt+KuXtsKyp/Dv/5MykSYh+08W9lV9S9fMt
wvre0PKgSbfZ1FSlGzp/oOJgdrwEGPbfYV2epGGKqTAV58BeBHahZATYHWmPLE13
9UJ5WeYzcJUfUkeQTnMHx7pokOOJGVhiICY+CsxJWH0uyfQ9PRc81HgF2gK81GoB
ZNYwtCZQl2i2rGy58Yv3fTvAdw3uBqfvIsIjWEBpFepdVe9/QYXtV+QNdkkslHkO
Gu0hfdcr5UXVX/nHkXQo9xoMhLOex9+IgvA3O+7fWpt/G5k3+L27Nm/gjka5FGAk
FU08MGrFa/TlCgIXFehH8HSbZb/VDrSz1se3+9B6lXXBgNJd7ldwV6K995a9uEJ7
BQIO795cXOwKcSOiYujh6LvNR5B3cjdPfwNwCJlVCr38lIwNqzcxipVp7grYVR3f
TTDsiI1izm7D/9p36RMptxeyahZ00DdFCMtjGvHV4GB/8jh2axx1q2th6EKPnh63
+V/DP+EPg2xOAfsdrwXxFhthXAsTbWKuTfWNUULJEcnibHE9B5nfxzszGMpHukIr
KTeMdfFtAWVKsG8kcUVDp0fSLalmfSIKJs+onM7XXUBUREMYFmmlWi17vUM7gdj8
YTpkHN9AOas33XfO8DA5xWAc2DPokon3iJZiBGY+XxkXNX/oEfeSWWrWATHD4wA4
128u3MACexmciSGUoqGzJAZ/TlasTU3xIEXGvf/Ngtc0rY36yc5pOVwqYHw8gxWa
/jtxx0n3OHDG47LnwSyHg7CMM9WCt84R5rvQiwC7/dNhEZfrP1sUqS/zoYPvbvC9
c1zOjK7aEfy9afh/Ji8llaQmKKQp0sheIHqt55pReOu0vCDIuSNMo0yZBaZAlrAE
sUQHw/7IqYKngCRZpGX+NqwniRZCTYcAM2iuRr0SysFm4a3xlGuxWYb1/0HntjiC
UovKy57e46rkFBicTPd6pJfAYRZs5NRmT0b0EfNifiqkxxwMOrOB+ucfKxP5IEr6
bnF8aSsQXcXHOmrC6A4BAblW+reJSSXgoGZHHVB+60Oponu9onWduveNCjXEjS1h
XJnADx2+KTP5QqNqzlrVj3lbMmL8+IDe7nbHbw7nHSZ7302AC7pEIs5giYG2XxgE
mb291WL4KILRd9bdUs6+4Til/rvSvIMzVhNeoNw+/L8jpcNeNPe3OZMGIqU1NaX9
0BcTtTYmzTPBPm9nSui9V2shjMUP+DIFv4IpPKtSPzYrkg4MVNb5+iCTaCQ4n0Pg
7ZdxE8RQJD9L/MLLC1AFrtWHGiRicUsPkOcBvmhW+voJAhpks4m95G9LSrMRImWe
zUktzupofjndt00Jj4g9agqsQ9vvcOzPML0Fupgt74OHgSwqvVFvdPKnc7g2lGVP
bw/jRPbuelq16t49tp2T09EMyssmbkfaiJbEC60ILJRfqT2nSgiOvyO8pJhuS2oT
p9vnVUnLNVrsqDJLgoKaYAvgbjfqXxXrbpF4nB0UjFGZJppH+D57OyZfRiy7HWA8
AB6yHLTcWBsHV4CGfP2cEM72IPlf4qlXKXrrwaq3fNFhkbywza1uquF3HqcDWQ7/
CI1nywTfKTigOq34Sr4oVTlSJqO/nbmi6TXbh8PpciBDznTT9k9tRTLH0UGccP7h
hvcK6czxGmF38ThzlgWrlWZlWS1Q9PYmGerAMpnoZtyD/MvaE3dAZuPP2HSOZR8u
38kLLT/yUUwhFi7smr8+XmRgd4E/LMXh2dGMhxIDCzyBhQhWsrJ1uNcYXIyHm611
30TAutqgf9l+Q4g6gALzEbG1+oIKyxl/WVvdmeWtGaa1nPyw/G0Kv7qSYO6EWVMy
bF2K1IQhMRmwkJLHi2K8AA/qBsPZBCqnb9m4LO6uVk+nA/cV6N5SOuKAVzi8DO0o
9I5ZlGcnuG0DdsxunmsNFu9azolYk47DZv3GneFBfm8Ag3PZeL6evITO8VRfg+zy
LWBxRUtKem+NZfm1dWgUfOLCaQfncueVDCrhFQnNA7jMOyvBZAd7cQesbmf+K8wh
nVxR+MeCv2EgcTV9l72XuR+evceH3nciyeGINl7d4/diqdYpJbLMzOPmSkoK+fGl
V9G4d9c1LEw+0Og2wxyBxwdoddtoT87V5DXyBPlW0TQ8c2pwv8XCkIFMqCR5G//U
lVMPQ/INzXV+6W66IRZxPV/OMYdW/ArFHtdjrnPii0L7qn5vQZqxK6/FD2PR4vuH
X9I9AolbcX6m4eWW56l3/JrSHhGp6Ocd4v/6Bw88qjdCfnmwL0QRghb42/ajQztx
jyKtKfZup4cwniorLTlP5iQvz4pAc7JuMUtWr/r+vb6IQibQysU91lUcnRqkmj0o
zsc+/CCZ3rHZrIyDi+H+ZrlryGgZbEkHXH+a2gHHUc5StWwxBDAgMb4QlSSthZ9y
UrNE7/jyN5HiOkFMX99mlGYEfXgIrgB5gSRp+16+OrWBmYA+/6qWDVxPT3QxVwHj
nV9p4JMFIUxOn16qS6FFvQ07B1pOOWLcC+azAVWp+eAiwraZ4D81bicbsqfAGmJC
Uxb7rkVP6mkgJc/KryNDucVOt7MCAqfyXJYiDyX9nsorI6uOn0YIfoPp6mPNVTKj
w6YO4HiFwiJRDZKgLoF2QktHck+Sd4H1OPGhCUTTGwapK/Z3ldbHR28wSIXXmzDQ
XwUwAW1xdJkLLAeFJj17tzzWpfnNb2OdZIgpOQA8fnxU3GoZNdgYt/fpO+Vi7w6m
MAyA6QJtEnkw20h/S45TcyvoOJTqBm9F7B715j+JEuzrCyxRU5sWP3Y1nZpp36qA
h4CMPuKn4M1EbysfRHhbYiZjY8oittvZemnx1/LcUP6I335dj44MBFDguC79WnLR
5Sy7tSPYP84taTOBytY5oW1AM9+hW66qNO7O+LzUFuMHSiq4pxULZcVbMK9s6Hzz
ZMitkkmWLVYwEgsVLPgHJ9bu2oadDP2ptIQzG0WcBAaqoa4k6x7fUpILG5oMC+H3
CmKdGQcYXYnC/qBm+Du+VuFu45ew/WMznjfuQ331MBOUN9WdY4n3UKRTxnf6UQZD
vhx8c1Jb/HvWa95+ThfkVYwE3574rgTFVT9pZuaVAmVDyY0OwVhpk46CcMKrxB5E
y+our6GTM6UXHYm1ltI0aoeUL0jwECIuu4ZBa/BX8U3mXvk8Ib7ca1rcIJlnT5cy
RZxA5sMOWun4y/oVcfHkoqmEe9FSyKuE4vGLEFPC517loWsNL6LZRKRZlgfdvPu1
CF7sSoZyl6TjomaYRBi9LSYCQkoGv6eDZhWvqseY5fmY74zOgd/PIFDhnCZNC7Do
ghB+o2syXG7livLOHNtqT3qTYZS+NaHwgGHgT8oAAr+Fm/s92mH5u63krHTDqMFH
i+pOBNwvqTGacrZkFqr/IFc+WFcswoKSRgKwJheEMQofY3w0hVD6Uz4Kd3DECpL2
GHm591KtSApNWuy/Bxc5DmysCDxYX2P1QJgioz++D1/225C/rumwCYlDlPBFnFT4
mFzyEKwoc0fb6penGfudVujIksURSWZeoisUnan5AVYaEW+gzFimKigwZynf57PG
TqKBPQVOaeO923Wq8bXB5VR2D+7AqGGtA5QYuHTPcPiint8D8CpMvzPMEb6jHjWu
9sjutk3BfUqol7/9Q1Z0CUzxcocfmNXNR5O7nqs1k0k0UF0QAbTvnZvdr6/GatfU
EzFOzGq67rhV762/5GIDOLkqdapjI+fq7LjpvbgsfW+5z+8o1bv03tWF4wsZqE0K
rfpzLyviNzd+NdEuuaA9IHjE6d4QeGlQ0ndy3B70W2qo0iCroEiT8Eb/5UxFo0Jj
G1JtuC2hQO5crelAxwksfBP/p6zQSWeNvMvk8i3i3WDCQS07FJ+4zvtMfIUa3Ozd
HNdxJAqkhRuGas/axtGaoxkbcA7sAk7Js5mWH0FYQr+rgBcrja9g6KRUfSuRcMxX
qBtwdfK/TM+Cdm+DGb+9F63slAH5vWeuaBb0kOiLBK66L1KOcMJNny/LVmsyucP2
EkAW9CDuVO5Ft5N1xVz5I0SnLWy7+3u7UoA1rHf5BY1QE75t3FLNLqGEhrt9i+j6
ZDvwE3oEHuEih/0KjQplFZ3vVCqdNsWW2K/dqfAQ9OtxV9k2thJIR6tjfvjZP6h4
Ea7x5xiUHTvXpnJXwpDrgEzGkyRiFWLvpylWDxPMfDt6ApJSsc8obYnuIBI4c0yz
YEq7EirnngEZcE2bEwSClzmd2A9w0k2uYxCHzLk6eFdMGv/HDNBq7QWIbzS8K4Qi
0KR1kLCL8uN8xe7WTMuXhQt4Am46chi2XxnrDjDuLTelMe2qPfDXfJZGsvAbj0Nm
lOldCdBOae4YNSZhhe8ju/ryJvJLmHBW32/xX3wYfAstPdDChC3yJvwEkaQX/vpQ
cjUs1JUn0bJ8Js4zHGkcQccXyU3zWgPtHjvWLsRJ+jTIYNUQRubvZcywhm7p5uYh
R6GwMX1xrj7NypyXsY0h54L2VWL1hjHPKxplsn/iDZlu48qKiFYPRmk9ky5Q6D+W
7yz5gibY9htBd4+iyfdvY5J90Rde6ScGIAJGXPPZKiaIxsxc7DVst3ETbbKuR3rV
O+uVCYapgSd1Z8bbYjrgfXaCtrNhm5ZMXBqCquXwKiQMZt5QMdsxsMu0iaHieEfZ
vn1Wa232SFqX/fVEKRS4PG7sAZp/m6X6NDB9DaDVP/YVuAM1zD8Ak+uq+fRbMOns
+WvDtw3kiPR1BsOV17GjpmPd84MaBd+NmFFsdAIbNAka/BsAyB4BNJIcep0lyUo2
9BxK2xgPnSY7aEobjeVdWAw/Axl6qGeYDDTHFnrZB8BZ7lyGu5pA39fy7hALcmpK
anCD6KlsNqWyU4qmTpmChw10Vcy8HuqvRr7Il6zebZ348/gm+zL0y05rF7eAphk1
o2s9k6muLxjapJ7qnyZANmS11DL2wTEMscjXub2DcTNpASalgycYBoN2GzNEpXyp
qgl51IpKTPiiCiA6HV9oSD25EoJL1UoGxni9+x+7HNjnq38By+6tv9sBKk0x6Oth
g9fSK6+ODSstXIBToxTR+kjIzGdsaioQPRYV0pMq0U9Z7UAmTPJRYC0xBy+e+jVD
TGRdg0fyTbFt2ajKk3wMaxY+komdKW8cZMUgOceWsaNxt2f1uYM+rmxjs4FaZsNR
2dhcQGID7dFkW3I2H85Vg0nXRa2lW4q09KxFO6YlW9nqkNKjDz5/ECRbR5vIBl5M
cJYKN+29u5V8g2EQxVNlh4FC+j9WpUOp17tv0JxmEickmO4cbIsWzksb6o9AEF63
juw6Ze+Hw9Ae4FpI+dhvp/nDFswodWESEhA3OBHb7f/4ufFvPsqryxfF9bWB/NpE
0nI9jKjBh+eZ3E3NWxR60Yh5sa3WQ7mGjgwn10RwERK/cTweFL4xI1nfzmAF43J5
gjX/j5vYOqY9m8bvDZvE8SoC0DJTtOPnBtmLbNVdeaPw0gwzx6qCXOsyW4Ibo3ho
HSxCpCN4l9Fb9crd2tialRdMpFItag06ZiMS96bChQ+4AjY1udQNQaTFKSyOtodU
M1pPEiVwP+OnHPMc5Shb5ispQmqOJ8TDSRyPM3I5+O4vBT8lehJ+/MLRSS8zwSAw
7jBGpUB4ClyzkjITNhOjSCsTN12937gFErJbrkjGuDWpGEKnhcpAV1L6C/wK7CjO
1PmN9XoXGcMMEExDY2qmy/MrL1uGT2wsIf5T5ftw42mCPLh9wbDovnFEJ1/crAKh
qO29EhKXK9yv8mb17OB6kUSXZ0/SbD8zFQ34fM8e3ioENOfv1xjF2mRppAiLfsnn
FHDFiO0Czhg1/Cypa6blV2UqedqLwlAbFl5fdESrgfEccg/T+nHfOAWni9EIyNRL
nArNUjHO+bR7DtVJZX33YHD0UyQswuyFVd1XhEx/8nGZE4EDwobcQ4DbEgMf6I+u
Bob83WnqmlT+6WtYZtHO5rGXhdhw9SEZueLujCbb52I2hgH9bA+NV7vCzcul5VRD
7q6KkDRkCf8wJs6Pkmajw2jPzyvGgehiWlLHpXeF6ZLFwrg1nEY4oAOiFMAKBn9s
YgSEygVhbMwmhJfHyRorSEKt6A0avtb79fPw5FSalAfxWCLeEuXAFBl9FiTtu55W
9IEKWtHW/PHN/0oGgHD9If3pcwB9lvvLx7dRhZ/Gsr5Fuk2qzJVKtLd+MAnkR5uR
4t5+H8oE+GN/mq5JPo8SVdmciyLMSS1Jv4Hl9mrEDq/wVleRMeuTCbw1Xszm7rpC
Uq3wrfmXeHv3/oWp36CCC5C9GdBIHpYIDJes5+9y6vNlTKs9Rf4UePXBi7oPP40X
NKFSHUvcgBr7HpYaEaLYK41kMraKP8JiRv02LgfFLW8BZiWqxintZ9LrF3oJmgrk
t6yripsht6FxzZUxvZdrGQRhS4q6FcWa9WWm6Z3ReX3G7AdKfupADIFyPOvN5BBi
vCBnrKFacjdwzm1bYZWnAumZJujvAKDvWfrs/uK4EJdxHrJs5zeEXfufxHGmQpGG
xkE4S7HAiFpdcpcN+LDfR0RLEwXXwUGNKTbee1nmoWGTpeh6cmroAlz2O2us6UAe
XNpAiq37px/feoiQ37Uj7GaPMqW5FjEdYZeAFoXvgF0hWvFkuAsB1LQdEi3iOLIR
TZGVpO4tRlH0LyXg7nMnGwXgPz0O9LEnn0hiJU+aPFxf++2lTCX7600iOJo4cVvX
oB7ygDMUdzz73JewhlNi3VR96W2Rf3PdPhNxro6lgDsO3HsTnL43j5OQrDb33D28
UHcdYnQHNKVupBr6CBY5RlcSJ2IURX7mJmOHoxrH6SKQbF4wWqoIwVbC2C1CT0Ro
ruxL7XUxYR+NdnxZnN2WDfvmFGyT9iTdoRvfpNOKnJg94B3hGze/dpQtWmeEPre5
3fEZqmpgQ+vu0udXWywA9O10s+D5whb7Cfl11lLoTkx5MOGSSF5SpBOPdDl6rnhD
rw1MKXd9rwbkuZUV3And0lff57UFceoBaabh8inqFoFxAy5w5HbYSrpFVcgmBVi1
M56eSyjj56LV0vTg3VdQO6zTvSLq6E7nVmaN/LhGXv8u3vjxeFwjNr2BXfQKbxKw
cX+73D1G+NEmL6paY6QUUE0xwI7R6TOVcnzGfBRcTQPivHnA21yx+xdcQBhb7yaa
i9MTKXwKylG+hTDO2gq5FYtRrzRCTFHi4ujivImOWf+gT9cugZxaJhp2HG4buEEu
8ug0bo0wD82H5gztTj52B0UPjpB1oITKEB6unQudJDBPHtyMm83hWLtVh+RO3dU8
78TeqyG/K0vH/zSYyliMMRURSVV6MiPFC80poudWUno6RxXjJ/QrKRRgX2NapWlP
bI+5ibBlPZ7IwQjb3FGvDRkKTtCucT0Wr9KOCerLbhwV1/DVnNlwKEszVZAAS95w
5eBlHvkmwV8M0Zz2WRW9Yq/7OxeCuiZhkHb3+r6Gc2FJev99dszhkx8g3BcUcrRL
rjiPRMREUrBkOBugwt54a3/MfQyJeEixwQeOX2gRR376SYEbgEXVdGEKf0xxY/BO
kvI3MFoLwwd3setHhX+sMN8JqayLlVIdcDlqw9ZdpVeOC9ZlpgSU6LUdrOS14mhO
/FNkqvjxLoA3y9u/EDC7qm0ZHIEz4v5fFVQqspWvq8p0+CzUiLE3zh+UJ6ZZ0ii6
IGqH2nEots9vl3AjmxAA7KimJMsz8/IupZXfrYgvNMQgtIuS/NohpxUvSriSW46W
cchz11w/SZWS14EjN8y5rVNc5YOm4pET59ODg/4Ab+6xRxaHcXCGlQ6+t5zrs5Hq
HD1C3QEZZmUOetJF1rFtOiFoVc5vKqOnGQOlzvrkrnYs1QZC6y0OomN7EVa97dcG
h0zz5d6+NoyhXi6qF6ftzj7xGSW1BuCJnCqCdf9QJKSob4Qvm7ClA2Lg28xPFjkA
FT7BUpb+7qEckDkdXmcUia1vHyEFNAxKKHVwXQHJnRbYxfWmoyJ80l7A+9B6n318
nfuv44tz3bywuki6fIbgbZUFwgDI6KO6Lvn4KrqUHRel96ZxtLxjhVvgoibOHtez
0kjQo5ALOFX+nwh60MsrqN3+TK7FyDiQ033YgToznaSSo6cQdSEhdoORZnJNxAnF
vy/yprXYIoFE7AMVGX4Xv0+boPvsEMwop0zWvg731Pc90uHkHQdSNPfkDFtKRbh7
xpOKZ/wKmpVMrO2pwonx8jN/WpTJs7sgEHy8Isfv6V6WtVx1NcMBYKxgBi9dTdLf
xaCWKwtqSx4tnClP2ZQ8y66I+kyHIkOsBYN5JSA9Z7PVfXxsW/SQ3CCSDzGwl9DZ
YzO/JCqybi3bLOAC/DujbtO3XI/OhMz29MCsEYXqhmo9SPD7+8TzhVJkY4u5NtsR
9Bh92rzkTuFPkj1eo6NRRrCWkx30VuWaj7QjEhl+QLgQid2KN/4yb99tZIHMQyIA
LJA7c0spD0v9OoPoDIVhhaC4tvWh0oaOaYeCpAAGEiYpQEph4zwGK4Qs6IDq+iwM
mnGtPemxaUrXLYZV6TjruPvMowSjlb4sopwPthUhdmDdwiTW8nRRbebcCgIT8xDA
Sn1ECp7wF3Ut+KFSC+ynYkuDnbba27RTc9+8K22+qDLAmkh17sWJfT9XCpPnEwfS
1sE9Nj4SkgV0PriR2sCEw8B5PDwceCNOfz7kjsV6fHMvH3ewR54NDWr1s8/0yVH0
AChA3eCJzGxpY1ovynJJEs44ckMSH6XIuwKuAKlud04i+aSjH6FF9JvI9K8w0CEM
Uj1veJSsS4PRnXdo/FJAxDQzZ9KNJHq3ltk2Oq7HXJ84Pmz0ilJrPlHJNnfsjz71
CzHp6i2Z6nhP8NqmKeg0GTSZYdlDRZ/rCsAH2byOC5OB4poNdFnflhKRAPuID30m
DQzruOJJOofHiBD6c5bFqmCpL3vkSzjDUhilv5x2qP7cEaUoztzW8ecbdmUR4HQh
LuAC27eaBXLWYc/KP6Ljpq8s8nrEnu0U4/CrAtd/WJmwkDmXOhpcd+jyE5oumKJr
1wdvsWBXxHQMxZYhVwYTiHykuLEB4NllYNlMohqkbi4E0ZXD4qUbFqFYeArbe9tO
HQWcycjZtwvAZ0XP64WIeXt8tTbFPPEhIeINPd87/gv/ATqtFb+QSbufyP86u19H
qzUa393pUd0AEDzn3mdtPgzSS/X8PmL6eXHjbSmHjoCCh3Ggc91idmYu9Nw7HCRQ
0G3Gzb5nE9pVC0J2AqBhoBcuY4qj/hxbHOLEydq959OwQQ92S12ogS9ct6NfnCtE
vEewidoqagIqi/jp4OFcvk3aLmBoihmomBrv7C6Vx4cNvPDywMtxo9ct+G7RbTmf
uS/+vVmToNvCjPHttPq4gX3YZr8Jp52VG+jSIREFILSfL5L6LM0PoWlho4XOF0wv
Kol98OVPesSe+zYhVm+e9MtIFVA6zD9dK3cZuZdd1WVmzGK7ryH2m0TPU4yUX6+L
EHgydY8DUY+kz8KCqFTKd/48+GeE0VOmQ9G5kZNRvM4u2XTKFESsVIIm+CSOk+RO
q+S2pzx57HzD2AWVdeRHfQ6dh2D/7+JckBuiKCM1U+Qj6EAW/542DC/kzBmDzhVf
R3fURdYNknuzoPtOur7VFQsPUzjtQfaZG2pCWP+p/cd2bOxsnyOPECA+/Udfopm5
iullS/TYAm4K2XhuiCCYMeDuN5+WFuDRHfgngUUS0EDRmZd7sbhrx3tfQP/IOBQq
TRE+nMs7usEluTeiUIHTWFMGj9W6hFNWBFUQ+8TIKklobUU7UeAd0C4+kGOcb9Vs
KGHWazq/k9CJNbJvS8TzJCOnyyog/GKRz8feB9ZVwGQjSMlQq9KTbshcekFL6CEm
1n/EPOnmNWnRBtYq6X6X+GUMSk/9uvYiY4yXBVdN6Kj+Zj5nzg08sK4koSuVRKFD
xWUGI7465adFcEm8YHvq9pSCLrJxXjNyHcIMTenJHHDtzjXyRqKT+efXwXMtYPhA
0FkXFC0j4OuiTJ9EzR3VIhWFefH/ZUe9AJ6+3Qx6sC2t981UvKRHmhMPXd3z4ecP
l38Rf3GO3WnIPTqNL4ywyzccplEf03OFa3zSYWgiBn+k2N9QWNFSE6049xbA5VZ6
3yI5FJeSHdy/a4/+iZcyjgrKEu+tvmFJhRH1dzi5fUouUuUBp/XBjexZ7mjUDJ4y
akfitwEqMnWxQWQOByrt7TIgZ8XqhU/cXUDKbQXs2PcceZ4zIZKJh2ET81UcrABb
EKTDJVSDacpyd+q4QHviTRrxBB+i1Ueqa5WKYKrY5EO5H5EeZEiMtBbCm4g+gowy
XIBQ7n/QNhnAAKMuzjcyvlXZghnbDI+n+z7elBT9cU1/BlVgIypX5HyKlreW6bGn
MwdV36HE3/bKZUzRYvEF+JItiFdsHxmuRDIvGBZRICtZBZTeiJrzS6oaaNNoBOJ1
kNk5VrXjGYjhSQZYGpRm8qCexDFRAcxLP/Ko7i2oTUIU1rRIvTJcpvxFYPQaZwE3
6jcmquggzXAMR+gRfevRX4QawlSaw3GMpfH6rtwGzVA3ok5+eEo3mxLubitV1Qze
S4IGRJA6V4iP1a0op3YxG8FnOuV4H/423It2fpAmBUgwxNeWKJiKCjoRx/8J+My5
fIL2AhjPrMhq72C9KCUjkgvab+c8zngYUCaX+piFWbvXI2u3aHu+gX8IZ9laz/z/
A6m8ckapSfpbLfZ9erEMxmyimxL7BqRL41UTY35U7dDG8D4wrGJLIQM9aAPn/BZV
Jbxzp8LCKevg2+fr6TvgnrJSxLl8lMJ51Lax3nRBvZOTDkZVo/iDSDNW0J2Vy3o1
SWZvcVwtsyVVwidYmXv6d8as8fapADMOpO+gENGE8EjQEWHV2u6nBrcnsndg+Otm
RhQE+unHcA9vkbNtdj+viwiG13Uu58n5ZjZOTXuw4p0SlhT8EzM6//J+NcyDw6Yy
mqPxfLJ87XfC7LtuWy+O1CMqCUSgRge8v3kvoJDkV4m2Qudczej4++mKP+Ky5mZe
yukvF9FUfZZmackUAJmv/ugfGMLwRnKziAArp1XxAXV+oQt3gJRsWxweMZeoqWx9
ThSnxEXI8+n+FKp3PjkXQJ+LZcu+9wOI5Pt9l0HufkOwBQ0B4Pg3c5M1PdvSvidG
jvwceYZIP+unHrJo4KyxFf2JU/mssS/Jxjj0ZO7tmi/kv5CoMruKUpgPycLjGk7x
fEbHRsjSh1+Ex4nAZ/9mP9ggaOnNcuXoCDzx+aTJdYZSLhqhBAH8JoZYJF4G+KRE
nxGO3z5VTvBGTx5x2+GI/WLVs1nBNb9kwLDGnfU6FjzT6+JeNG8RfX2kqpMcU0li
/uOgyXnlzOi4hXv7W0huMkH29GC0onWD05ll7himMLDHkyHv9iF2T5WTQgD6Ec0X
HfCu9kJIYJnRER+D9hdzsOkS7VariKQdiazOc89iXmp73n8JhdRCmyCh2K4v87A5
JZFR5Jz4pbdoO/WYXzrUmHeRqtSTsGyZB6+EdG6r1TPhhqrKSb455Xipkc4M7yy2
H0jdBDlf6NVk5BWN0CMr72njAIoAbDtsHY3T4gY+cPW1CGqqXUa0ivdqRJhJcBlm
tqiRnP79U5lRQTz/jgAG6sUt24CeHadpAeAp0hdpDf5qzxG7vBLch2fwJct4OMxS
26OqDGE7w7BAOJUWBLtbwwcVE2CRs08X9Zyqhb5rK3qdAO1omjwp6HntW/RbFTrI
ndGBCZRyAwlnz2+eBTVI8cOpe/Pbm3xT8Z4XR4VoLiORg29lGpn7znGDDNpwSvNy
ZNJvvq4G5uYq1nRx1k2fqLWYLFVmoQrJKzk4Iut4/Hq8+Kp7/V7QPH9MxeYJlWsA
44YG5/gN1isD8x6nMJkb1pArOdzwNO9nqmxizvG8kmU5jcDZUxyeqkrr9rj31ess
tHpTGpZ9D48JV7rKtFHlUO17egvDzjezDPCihECPVG/KQ08mOIiWN8UetLltVZA9
h9Xx1YCgJwAiPOVLA3mMsLUyrFigRU5oURY3e3RVYhjXTupKbb61+l2+GqEgkTIf
l8Z7MkYrONeO6AtoWB8RamUzIYd7hLBME8jvUwNt84O5GZ3xhWISQRwi0bpGHaVn
2Shx/hP1Q0bjenG7Xazg2YIB7hesR+zuzb87XmZa0175PVElf1P+KcoI4jKRiC9A
6WWQuaWmHCLh1SkOeuTI/KUe78jTOZqRRU+iOA5cpkN2fQzLMIKTHCCbky5AJiQ4
Lv9XgtZ66FFplMuE3k68dLA/LXZ9oPuA6NYRz0mKdcqAyDm8Wb4at4Xl7UxzhXMf
Vq6A7NPt0nnkijVfPMHIVDAoOUf9DYj/prAdqZ1Fgan+CWVOu5V7vHC4cqgV8+df
MP6X4q5qybrs8+LaIcK8VeD3zo4Zne/zfDAxTeuoObbPGW5NbsxfUVYc3vmQny1n
vdgjptdVTdn0hKum2Zqrpw2TQi48/bak8I2h9UAt0Wm5jAEMx8H7nz48FQoKiI8y
//mrdm/7uAyYmiMgWW9CNyBDPMf3gPwVv6QotnOaFCfb+Z7P8qTqaZAI3v1jux2A
c5xEnq+xschXPcbKmCU/M9E8t2o152cxyifJb0vTx/AraJY5XL1fvkrskY1ZcjiW
uhQDNb6CFkdKeZcXl1fBaixJAeGO0CTh7dL5TqbAELk489SUnsgMT4QszIu/Z2lq
lf5noyL8FMa28NICw/PZ1Jee8BL0kSNaAgpkCNBIHIX5KRstMN9NWHl1BBMQElIA
W1kU9ZDiyJZzmCLOSB0CUuV8qdhLwZ7UYkqGnf8SSRWfEyfNAJ8ugkH3ZqhOkq/K
z3joS2L/nmbxw+uQr4VTro8PAnMRN8QL3g4+dzgkt7/cIO6+Qn8WP8e1jh+N1FOu
35JKShwJNPIRhCtLe1hkTXcxSdw4oP32V3U94WCLPXEfpWnzAShWSCdbOip9kCej
ASxlJ6QSfvx/4lBACuUbH5xGgDJH4xKvV9mF1/KeO5yfwnxcU2g+cPAlgmXDMMDv
/C4Ftqj6eOkwdup094RoGbZnaK4yqqpLTnFaa9bmMz7P2vgHMuTVL8pGuPPLD23u
jM9fHrXmDSwnLnvu+lRbsjMPxYd3L0RtvY0QGNPBWCiOxLktD6dkUqJ1l5Xmzkyz
N2rBHY6OwrFBD14x9cnczA+NKTRDdjKjrRUdTQYA/2Dlqz12rVA8I/ZdMCvZERHX
Uekq35dot6nj1QQ8YSdbJD+1PhU3P4BFsBjN5kV0sm0zSoJh5jLgMajGcFTADqfh
C13kdZOsPsfz7kYI+/yKxQoXYW5o4VXN+SC/McMAWnKuXdZcC72l5MeiY7Ik8LxB
r6w/vRblYXF3mRNHAR4JcDmcpEwnGLoRfxEC44rGyy//PIje+WnVPCINi1ovuB13
VMCY8P7PmrMLvsBMFcETVjMwLaFViV05AbF/aI3Pyg+fQs5XKTwrHetCxorDuxZ5
f/F4oNHqGn9/enL2BuC8xvv5H7IacctAN46KEgxK2JJ61HeNQWNT/LsnxjrL5qws
xIDPJqqRxGIj2PQ6//wmezz729I9omwx6eMNdZbGyw9I3U8Ld6Y+BNhdiLL+c3W5
VkfJNnbOuIkyxkHPbCRX7Jd+Spufamm/lKzeyk5ITKzkj7dqZokYb2kaj2iS47//
rX3gt6yr46a/pPFjEumsbNvhDSYwhxrbbSOrfaqcLjSQw7Wl9XT9cQQHymeFXxF0
J6oNR2uo54ukTW/buAf75YdAeQRFBuXwVxxcADrWgqB2YFe0ytf3ZaUtpyi4xYmH
QMuU2mdRBFTX7vjVfc/y5o97cvpgtDNvcGnx2S0xxC9IixFTLEGr2uNueP6piVM2
PfqTRwSyjN9PEYGk9lQ/6gGebFTV3lCB9NyIzcPXkwtLXVzJfeg5vCEXlZH02znu
I6gkR4BzrzxJEC+oaz7u2PoJX+bH64S41vUgaLjUU6DhiIzSskrOv36SaJRW18eI
0fxjhxWdP8+cg//Hwf4v36G9nDRfUlQgVeDamxlrYpW6ukp+o5aB0AsAVDARkdpf
g55FgFHHy5brcmFzmmt8PjNWJgy4nOiZ0BxYrceyOEOPdIADi+u26XHeGFhWldt6
/GNsndIcm2M00zcK24hI2TooKckg8HihJVtid+6k1BrSPOwqCfwiW7pPmDieUnQr
MPqQ9ndMksMqK++YkrfaWG3NBs3xDaGqouG0fiMH3Pv/eZHu3ppHRJC6ICvtHJVN
TjOpBpKJcxvHLw5vngJCcN95HZAXKANSqtGcCCuiYnH5KC/Tjd23oxUqNDGafgWG
jNpF4U+g5Gq43fQpSNQOQPZwUiOS3eb00UtA7ULmN+onsirR6FJj+NtX75g3k5Kp
c4n6EirUn7w3Znz+RFqPUKS62c66/ncVKSWUnQSfeivXx0JJDDTZtMJ9sRAdgf0k
OxaP4b7igliIRI1SrMaxdZvvYtFcFW9b04RB+bbzYzBqWdmKxMB6mnYMuSj3WJdP
F3ZnSde84878cQ25WVbNNQT8Dw3hEH6CRcMUtAoym218uq3XNAuOeM3pnr9hfcBt
BsOgb35uNyAX6FJFtoddzTI3htE51q3dwszpTWnn1MGyTgz9PLb67hpG3U4IGjQg
/+X7wXjSJAfJK4rsqErWOn20pjlPzErsXzfKe0udsSCReqmV8B9simhLl7Gqsl/B
TUwtx6LZDT0Z45qQwCbNyx/vTTJ0tkOp83RpRk19iHSTFOK0PGNPkDlMh3s+IKtj
pAJrscceQxMht+knFM+CyczWFRi2ufWrwdmJLq5C4jswRWHHO6ttpmhZ6nZxwNx9
dZJOUVAc5Jxr4eAUts2idPqTxT8009C46GLL6xVr0QLK2HXxDWW3rZq8PjMdc7TJ
vliH+4VfTyq9LVDUrxo8zTC1TEcSQLj7RZyLABbuKEl5iNa16k1kdPwbLZ3vFzNb
7/HkGinjraQg/Jk4izkd0Woo9+Vmee0vF19ta96B52tgpLs6OyEEbXt7feJMBPAT
EFyhwGgA4uNA5latZITQBGRe6Zs8dDwBO0uJwHxXqIGwqm21kZ1uQLHEhDiiswtP
C3YhkSNqFIGDJOABrFRlZGeFsHxaZjJ7FQwhjwYLBfe+9KYm61i4bUqfre/0rUhl
OOdO2nMYJ9O33BVpqD/cF8DHnco2sXBQNQi3TyXHgcRQbNGDGXtQDa5aXdepch8p
tWGxUdDxGnj0pdrrDmYEhGY2lBgm0WxklzNwLlI13k38atus7pCjy3u1/+b6iAy3
d7c9SOv9C9dpSN5UNan3fVoNGshTjONptvwI3l5K7xH9w/uaz3v5ijHdXbs8iAJR
OLo3b1vE07uH8BElmDys8t/dUCB9tii5g/A+BEjAZNuOqsIk9q9uQJi2t9FBq9R4
PE2i7PrPyRilXqEaSjGRdlIDwKwq8XPFNQQ9W/QkbDewPK25qBROWcHcJmZLHL3I
eDJi6jk8+BmR9yxURQ1M4thVkbpGD2C95iAOj9CVAFmDyfRnOIec8a+1o9Oa5oE2
uxoRLmN0F6YdgoUziA/A6qD11Q1vxg3LbO7Jalt70dxUzfMLT+QQ3FXFFEDRxjki
bSLIKmdepJbry5LzbQPFl9gSCegi/PQ5Im/X1fqQDUQAipyhqq8hBeVnf6GQD4dS
ePD0nbzlV+j5s1eIhcD6QfeLPOapos44+2gdtxr81dWJHRZLLPDJ/kFms8CX1VvP
RFCOkmq20YBqgBgIOHW5i5TEdiZoCjvQSz+OmD5Z5Ui6/Mycglh27J4ZfIz5yogn
Drx1jOw87GjyMVy+BrkJDXIy+cAQXj/RkmsxYOBKtzl7t1VvW+DoOU7/vV+0r230
Hveg0G1zWgavGdKFFrxy7qv6dhnFK4wRyfKIHBu3zmOOFI7/4cYvkiJtRdav593+
LD5tnLFu4nxNbF4Ld72OqC/9cSNJ/jE1fB1v0QAh3GFBw5Jhuh0B6IO1gqculWdw
W7MUQtWpcNWT3AsZJKPyFfkvbrZGatSq0kUkZtEbo6LhN9WYzVURWOyzL2tZgEXj
DURiApxWKgqLbZcNtSaBhbPfRDRQYBuViypA3W/yiKJJXVqbDI9zpsuqoCFThlRY
orS+u2PG9FYZF/KKjBkcO0NODXpuwzWryRxTlfgiG8OksWOyz9XH+jjL7agOXshw
suY4+O16icG3ytx17WJHXCBP21MITF8V3Ay5KpFCIbOgvLZXL5Mxgh8xsUbnWAoB
M8FY+I3dzDpy5XUcorWCLluhq2/JPtRKzJwq+O3KqCgn+4EFXIgD1nycDZRFrP/1
JuBh2LgEXUfmOzroCdEPRlAScwR2oMfsqbizl3PwtEre2qowt0WDn2n3hCClbnkl
Q4bclkglu+Bw8h0z5A0/es6E88K2TcYxD/Aeeda2PakAU3AijN7vzN2YctwQ4A6J
TZ/B5JxSpGM1YReiYEXH4PWLZIVumo/C37yrBMfyKGWCAcQEuMJGGj+9npypks14
Jw5pHp4+TiAQaLpWKwwg2NMc+WLZNHVymA31SIN0OiPFKFYTq8sqPOwyo6rMfuXb
/LUuJGrdSoyO0/xCUuvhPb1P3xalq/UlMZdVHVf1OeWk1lPGf/GdYEJp6SDgQunE
MopMcvuVcbZJN/Rzko82j3v4tfMp9ynemqETfuMoETGts8fWDa6H6x7ENmGo++8q
x58KDf+3usT/G0Tc3Trkl92sdMyyX3nNDSz1RqQlBVYM5P5PcE4VFHFX2He7rk1g
XAZE8jyKucN5yqhXDCMtHOIhOCFjvwtjpXS9OQlFOmVzD0zOh0oyQslEe6AmqpfT
LnT6z/POkNYr2pFwTi0IfyOJsDFe4PlxXKYdgodUndQVJxyndQCjMY4V/kIe8rGo
Ma1KiLG606Ofv3KIrmXMAuQ0ikg09yBuehY8XFUrEk4gwCUL8wrIwYP+8J/RJRHc
rw2DtmPkZp/NLmd81R6oigFTVcu4sH9kPk/WQzKxuMFa1t5aT3vSgaaI4uRuE/Qe
0bUewqaubD7046VAk1mY1wvS0Q07nacrlLvUBx8lp9XfTwV4ll/9Sq5zeAAPL7eb
/USm5bFEhcucWj22ndK5sNBs8Zl08UpRavJGOcN+uD8uu3jQFkeJP1/4tzPOJOab
EP/sv935Z46AkWOxxokeMPK6vPMgCu017Hv6FAFQdUSWeKJZLSoY2XzH7odokqzh
E7JrFnbUgN5ql/cIFfvOt6qTpGEDA8/ALa+XykguSFipb9Ls6lswaI/aa7gtRlLZ
L+710bS1DBqm7U3XBGUgXeJBaPW/Nf7AP+e/gqBRpM9Nde2KxHudgOBx1rZjG8+7
KzRQQ/kemWRUr28jeQ28alBM6wirl2W7J5MU14173utHxs8lLucKCTHx0lankBvO
uUPBHEShk2GpP/JhcAx0uJ3ZWTEZzN5ZJ32NjIQRW5RUKOhwZchhKiItR4jabIJk
qrcjZJUmIcJeAUaEk9nTpxazfV8Zp1acl8BFeQhBjpZp1tnjN7mRvcoLAQWxHoiD
sqg8e640Ki5nV7y8V5y9g/6arGC7x2IkVURiu1167Cl3pf3Lf+7gMgwmztbMaE4B
WvjPSi1XO5BB9s4eXNP2fZMVCgBw1CcaWnnpL9+oEnkDZtAy1ugl3VPsT8cuwITw
SvuUIa8TqBYjNtmiq1qJXjArL8dhlR5wA6/3WyzwDqF0x3vVuobcPlUQfL2vt9t/
uR6X+agpMY+LRWB9BdfN8W2Z6AJkXHmaubDaYPuJvcYZ5eYS+yK6jG/SrsGbdTH3
g1sanlOT+EBJIWpC4clOkth802R7GNKWMZL/H5kCKTJ26pQHGoPvO8j90FULhNKB
Mq3LQcn9Qv1b4kXdb5y8+vYWmNOIhRGAQyvi0c9s7RcARmJmKuhoG5gCCSjWhg5S
SadaVj/QFuyNSR0mrpm+OUQs2IQ18v2Kgxv5+zPYN3DulyUz6f7KAYQgPAOdxxT7
PFdv1o65ZGwmWmJLYgYZLX+aQxrKpXoOb32ThZM6+dk9uD+pc7u5dVQ5og2s4tH3
V/G5qzsiqz5ZpCixH94iZ03hBNIn34MZ/oXN5/QY6HvLrAhH2pB0iOCeL7PenFOq
0FYnu8f27YZO9KzbgFNV+bf3+3ypOLmrKpWmJf2IHoCylk45dLdTACbJKQbVKXwh
LgLFyqcHgx+PUKp6mRcQ0w3vs6psCBR/lX1zxcHtkDYH3UToCOtfzGXtMKwEfIGW
zSgaFiqulraYJaLE1nEodYGkkyyFnvRHqzct5icDXlu5+ZL1AhGA3n33Q0q0QOht
lgvoFEED/XGgzX+7fovMRSIDiXVMw45NvlZFVvttC37CrwYZqoWof66ujw5vSA6U
bma/Yb6O9HsIHqex+RDMsbxQb48SGQ+Swod7M1Oo2EsiClDXhfbyeAhXinwDaS/C
I/9nAvuX/IApmfcQZIW9bzHTD32X7tunXG+J30A+988pSFDi88A3ZyE17vBp/whq
R/yowTiKqt7ZRWUiS4ULi6OZuPSUQaBSb3YRPwFDnnqwijKuipyFUC6NVyURT3ZF
pp9WNUR7CTCGS+Mu4DIDd28ePxkLNzqzYdxGatlNLqk+ebpMTWInDkRH6KTuL4dU
67QEuHnqdXLPFHHM3fUoyxtz25tl0mj0In4hb7vNzBnpXXJsk5psDhMlZUOrmk+7
ryOL2CPYHt+l/U3gRph80+/7bsE3s/srVjGjeThCVxXNUWX6Tpw9heqkMHoBx4pl
QrEy8EP49lCIXEv4n3CpsEHEnUAmg9HIIz1Jtu6/ZUYqqFIEENfeQCbydw7yiAhT
45Hlvgxi2s+GL/i796vfrRYYtaM4ly1EAyPyMNc3jOe8TxPUBANiIcg6qWQuBRTQ
+PiLlVTmnZm/r+0lUsx+JIaGAz22sHrvkGkeXM0AEXPyPDR6iIfSFRAH/Cl3t+Uk
C4ibAXiIX435qrbxFnxd9tIxqrYStp0wQNcg4mADZYsljY/suST6RJSOv3HgOBUc
e6aiVhkmessYegXPooCvkewvUYm3/5sig2+ehOntpUv9AMMWrT+1WR+B6MnemSsq
4mELXu0gMC286nNYrjgdnfNhbMS9W7lPZL/8kZf1BobKK52vdaHpoPT6vJOlrLhB
PLILkbE+yDsQcwfH6N5MD6IFNI7oNi9JZ/uRDeaZfMCdVSUUskSPOf7XsYPZILA4
cWcrucXY28SgmJy9Qt2ncwRHT7TaPSKwqcS09iIFD+LokX8nL/RwhkgtHn3mqOJa
dWDJi3l6iVrs8uSo+Rf4lWJoB/eBUayQsUiZ1ABTxPxOmQBNiAOYjUzy/xygO3Kk
PmxPSm+DHx0s7kEV1zMWegeQUz+hMKMvPiEp9w5ewwOJuF12W7q9PSUy6aXqSWwt
RbsEXGfHvRUixvYFpt7IFOrNDs7W1T/pB9ft32d6fl4jMY1pkLfLGXWQXlX6IuqV
qVTo59PoavKdyQEEhwrWSQwZdLdolF1Z921AwEVISojtSIYyhWzvRcpTFVWck7yz
VCrX9JSRZfbBIEbv/ZTMhaBSofp0dgd/e8Cnj2zxMzjIS+6CvKeswWVjRDGuMRAE
+8eVZGXEGNKS/hGz595h3kedJib5wRUE5Zgy9OnXDADrd+mn6UgqqtVrO23mi02p
GJrH1w0uPZWDp3JfDm6cN1EIIpPPJ1aPP+9Nt7Sk3Co8BCVZIi4ODjN0x/BdxsDu
t/DpwwwkxkwWYfBoNTxJfFbJZzeOG4hhsMLV0qLa8T+RbX0m2+9c5KAHIMPkH7vC
Y6A5L7tgTlw/7BuhUI01nm1AqAmA0Qe/F9I+9/w+uztvUzFqyusMajg8Ntt3pxd5
5f8Nm6empUJsAQK5qItyT0NXUv2+htSTIWqYy6K4YpVVsTgpK5natz9VXwYv3t0Q
MoMBiYmy2gO8c9wZ92nvp6g1GVHKCQtZXzUfAr2c6KuRbPYPQEP/cCgcdqVTcvYo
ZD1UHhfWhachsFxvTYAbkvlXP2cHEw8cIfXOs9GWvcURHmooKWX1x5b4oURbP1gC
8ybx7ma7K4k1o1MvPXLYPR1FEA+9KqkllFLQ72M5x0vRGLNxBbSSx1nJcGo+6/dO
A3NtHuZrBLO0oRwPUqKqjJz99Sws2ypxILMf7Mf1vSOc14GJohXQV6ia64ilpmNY
sqXh6s6004/lmVguHJ10yIyPYPoDzYpRxwzoUTS0eVpCpx599ZppJ1MLAbEHItdT
NxAc0gyji3Bhpd4VM9mlslIq9KuDrFZ/1of6TL3vCqISt+9a9xQodxLnyXlRM7Op
zWITh+BUdL3v2YlBPBYcOrde+EIUYGr/k8AB36SDZLSIiYXjJ1mI2WETVkj5VEv8
hQmAgZvtaAn/yI3s3QY5jJythassKuGN5wz6HmRfQgLy/n6zl+kShU12CZNHw7ZM
Vq/I/bqM6mCs3+Y6YzVcVAJeWcjKnbfY2XpivY+DL22h4Pt4V82HC/AqnISoavV+
1M+B3ouWyVu+pVDrQ8H5WDRRrUQDuoOX8R3VHjTtCPOiFxaOsK7woZ+e1Az+9JHK
RzceRkK0gV08eL+9DtiwzPf2gM5NztdYb/7aIvElnVsKQUkaeqk3sbxVq9vOMnaD
NoZbzoG9uyrlPH5TCBAjtJcaU9OmjZ9GkqWP+FzMeA5Q0XBTQP8CIDBsGkvYXdLB
51wOfCCX1PF/bE4kik9NbpJj0z/kl1IZ2xj5aWcg33kC+l3yC0dNCnm7PqjEp+Xa
wo/TfKGWYinb60sE4p8iu69F8Vn2LDdQAqdhvFmYRW8Ec5p4cYnPUpqTwYoL4Ho4
Hh0nlN80XkTdPS23v/Hh76URx4tewJJOFQRK0i/099hKoJ5WmaitcdWKxeHhqaL0
E99vmB4EWwUltcqAekDSIZsbZM55qdJZkTjSyePnhFSXsLXmyuQqXfLEVJzspUJ7
9tGn761L9UXh4u+gbrp6njL5B7i5BJ4Gfm2MMmzE5ELEqUYfAxfW/iTtW3VNrbAP
ocmzA5c37ovFDavDuDFzXbKmXf9dYUJBYxxJNZa7PrHR24blFgSQrGWJ8XS2xBrz
Z/eeWkWYqhHsrb/6/HTAPaDAxhf3QE4yAhLTi9IMVv/hejuu2zmfp3RP/OqPzScG
WQZeaTHOqcKKy8fTrLnP85tjiPF1GweR+VbxjXsRCHAxo++bvAAwYrnZIp1Uuymi
HIEBcCpNUpXVAqjlWSg/0QaEPYmEnz7GNtin42thNzAi7JrSOGiNJ4IwnLHpfWxH
O4DfTa070rFUzuWxpYPKapbZ41sN4DbSiWtDzKQJX79E65TIC0s21LD+nKLXG+/G
fQCYqmFD+heQFt6rSq9JI/31gYeE+7QNyyM5bjGejp7JDrEbqRTiqq45sgJkYrGN
JkCNUfCwrWYfALeg3JTWFzC7hfF8rdV4knFKVcx5RjYw0wAQv2Xcdp9B234xmHLw
J68Fy3rHJGmEYkMunHVOBIWIxEwjILZCLctfnlpEim/JBfn2lZsZw2dXcs2qtyuW
aP5rKMDmzcFUulCF2S9TspQ+grm4tAmETh4aI2str9k+my204QHQWvwHOsL73dxK
8rdDmjKRAVp0WnXaROl2Lz1QbhD+vO3n2od9yHAScfUKDlDxhrRAtvXnilJjyKF4
kBOpy4meVv4DKoYdXE/fOB2///1e5fZrYMNL3wwwcN2lcZ+kdGWkz3FQ/a8/jrx0
otKTdQvRGcWlguSyo2jOnDuBdHZio8Qgogb7G7kS3Ks2GbgQtFXnVsuS3nGdcslf
D3W2wEg9QMzIK/Zd04WftMgYBjV/bgKACafdRexDhWpF+2HtwDhOAsVxNVRmsGzu
nnNfZrGhOewbZH49Ua/1bEnPPx70XFKM8GTCgIKXwHTQT70XMWayMDevZc7b+mrd
j5lsl5bGRrCZjVaxx1MNb5BS/sTyn7cl/jxHtJXUTPA/z85KbCOyZpp119HkO+14
MrL8zbiD4afKRZQCcR/ExI/nF+YKFwf9tb1bDA0PCfajSR4rqpCuwNAqDzGJENzg
CaY9Es4Im3FbhgIEZDIyIb+6rvakYlND3F0UdXVhrZw6ymaBSsl4eDQn90VPWvzU
/UtQny0dazEb/VNpe5gni1eSZ1MPgd4m6ILis5GQcWS6AJiaozjBwohEu6yfJCup
J8yhT6WSF/AtXyacU+r51oAPUSd7Mp6b4m4PV//O3taLTAfFVF3caahJ+2sqlPgA
4YR3BKryERzSqXTIvsWtelsMELubQe7GCIgg/AmEf0h+zViN8MJVbH8RoNwQYcyY
yTPeWCmuNGhr36NZzxRDjl/0IjO+qcz1H2pBkcEI318k1fc8bLpRu/6Db0WSETHb
yT2JCDdLQm1QSuM+m7ykqvChDCHSq2f3HlB+cu41QqQq6SGppR37nKgpby2q5gxj
MSzXX3048YpLI68aSD7tbq+fmnI2OIVtJQn7Da0dJwbOI+/OzIBeVrJuE2p+TwM3
xGLvH49TEyMyyNEsCZqlVgIfLkNVMt3nT3y44SzHx/s74dMiDYsG3rw85QWkLNBn
tXv/YTBjN0tr4G2kBoCihW29FZ9oPh5WnSLVGw75MKY5d9vfMEFE5T3M5UezbMqB
JICyTEPjDArVT2w1G7ZER19Vy2S0pA93HYBPSNaXlyVVToi4wYYHA4JW3zPafJBR
EtXxTm8MsS/uIDXhB7JojHPuEXg/0So2m2bWR4asyIY2oStOzwDoIlrojoAByB0m
iBcWhYVnsNtnlbDh+tvpRRMqBBEJ8IiGk59SXTi7NVSyYuLYlU5nYlRw1dCJ2+xY
be7pS65SseYxMSQTbND22d7pk3BYhBYMFtW1bPox8N04ifdZ5GIRJWkHMK510ohB
H004DL3y2nueD9rr3DlL4cWxfvta7kdgUfuImvO/BzWdY2ZOQHNU9R46g9KU5aYp
/85qtPvAsAS3HR9hzGn06opl971boEePvU66Mnus5FlF6hUvYCn5hvLwNLDobJEL
k4fAZXSWmdVks+lP2NNY+febPzvMEDMqrBpLm7lw1hjnReVKYMHkuE+duQ3wSC9h
7mq0fI8s9EODwF4rWJ2J7zKHQzpXN5pNEC8jwA7FsFpoKtKieCGd5jL8pcYAxAF1
9z2oPt0Knli+zJsMT7YhRy8o63JDxLI9hkdNeCXc4Q/Q204PESIskjC4Ha/j3tNV
BfMjeV2q6Dv9/kkbtavlFzDA4RMSGXxIlqBYY3ky5Eym+jZi9g5Uc624zKjQ/2Xy
6zf6JqQiRhTDSfBsALH0aOK0JmnqHAdZnguQTvzAXi+h10wYYvhrZDBX+C3DNK0E
UyEnomvxkE5Ys1NTwlB4+g1c58XNyOytkCQPaJ2um2F2KF8GQRUWndTePh6cLW7Q
ASABGSRzegRkUpgOVCNbL5dQNW6uJMPMUREX9tb9MPs0V7+RTAJTh1k2otfM7VNU
QxGn9ihxD3n1KO/CQloEpJz2nu8zjwaZnQPdHS2vJE420SSoOR29fDYcZZwdw9e0
Vwoc0n1pL30EllWpqcvG6nVrqYfqH00ySfO4w0Ik5P7vMYTgWpTUj+hJTfkD3Uzx
mIPmJHLPK3ZLoCLVx8xeX6nPRcbCR77EGww+JkOVROijwOnpu+oSGE9mc2ZifFLG
4agaGWmFBheePqyLwXVxROW5IC2iIgaXahuAuPzTxNqRoAzWoiAGhoC7btOgSnhz
MOQWkRgfydFTuDm3HWaDgBWVZNFJ+YIfn/Z2/P7ECbjA4dF8kb6Wg0XYFuSaMCUS
dODEGL5fjQbcTqJtYax6fcyMKSrmy324Ni24Yu7NebIUIJEJoL4AczUHbZCEu0VC
7MH7sBYY4vpHohtsXaF9d7LM0IqWIU9zk8EgVRZfi6Ncb+kSkSSYHL7WqCaEnE//
ks95Amh6/ijs8IJSTJO1kSlqHJd9P8V94GNAZTZu8WxZaYia/mMaVXlxZGBoGdFU
i2cBWnM8ySY7BvpnwDhyDFW0j1GeHZmBR6RRkEpHFiSlfk2ZBt1PNBT9FsDY+mma
o/vIRHBK3sJdY8UFy0/x4cYhOZvGXt2J6MgNNyVJ42JA8UEakkmRfkNmbU1UkqsW
cgGyAMi0/fwGxEZqlod8NnLbLJdbSnuYWpNRz79XlVjB4+kkeccsMijZyMLpc6HY
lb+zapDYrfWAnNnuXgVn0Vdtr12ACXcOqDn72KCPUQo77Jz2ScGkdp5rYVmQbmBN
kBfgGV63jPph8GAJFqMqdVqol/fRBN5tY9wvUYcLu92+Bl+/8pFnGMcDqG9jiLhI
cMagWCrpwt7yFL1QP04fUp5CLOezJ4drW89GCM28w51GqF9rUAda3QDNbGePvPgg
1cxY0qSASJkNjVsGV9KnTeVuPwsoN6qzPvcyWJxCq00/8pjL/v6QMfkmkZ2AAa7K
aC15+wP0di26+ipnN9EFC75fKXpJPF2quuP6XCZmmIWqXtEcVpWhJONlAeHq0J2C
YAz/gJm4/cT8dogThb68kZWexlNU0zNAEkyU6C6s53CZFbdPhjpaPigw5jv6V3Dn
U1B3r+W2jMFgRPyblRnDWoyjk+09kwm6vQjf1yI3BZF+n4XtxyvoXh0Fsu0BZ5d5
P+R01WGaim67J9GJqOLatUyYmGW8MLDM41eEuFHsNSOwhCM1lTrzSAVSU3mZHGI5
khNy26xsSIUOdDSRh424u0891r4sEEgG/UxbzOug3Gk7Pv7osrW0f8R8ziqZW3E3
qzq7RwcnP2vnXyiydwKV75+f0qfLojzQ/QjwvKQebb2voeACaAcX5bgyuqoqJXsa
UgPoeAKBMIEm1Eruef7MRdXZeh2+EYJXHINLnFLyBtGxrPd9tcoiqDq3bQ3tZPz3
ooMjcqxW/YwzqLMk/M8mpcYzv/l4EijKkaPHO1oMB8ybZ23pP9MzNRi9GjrsFzRn
N26k9bYzA6q7io0BgJ0gV00fyP2fzIEnp2YSbA8/3VUJVwF/T6Bz31NSNebHqY1a
M7MMQqMVsC/0sJQVGqNj4jNDrkxfDqJD7x7z4r2fIN7Ksbipn3cF3zrYnDoqCkwe
dJvTP2f1GB+cQhpLJ9n0QOQuCH2WRT5NtODXBH/P1SdEQdF8FgnV3HXnqhbCy9aE
UQvUEWnQA5OeQu3aw2LsH1JOjZlJxeQ+LFXf3kwK9dcqoRewAtFReYkTDPFJBTfm
Ldezt2iCSeUrPPCRGAhHa0QKi1zMf5MO/JXy+rIeAS5SIE3jMKdfyR86AhlcnIpF
k6RpwAUctGCgCdJjtZ5XeFXPtlU8BCjPD4x59TVFrKMDpS7UXjndS1zIg651ASEA
suRGwQpQJ1Qto82MXB/ITeuFPSO3OKcws/RtI3Hq47P3dNBUpaTGEbStlyhH7zP2
HubdcWvZt+E2/sdVI7QK6FgLEbWmAmLxQMa7TC8HACdkK9RoIGXa1h5bUCzBlASc
VZ/y8zRPFmRD6dIOIwqKwc4HR7eaUyzVPxtb9jXv7cQNJTMHlwUtJzhRWq3wQd4E
lNru/8+u/iI6JaHMX4lCmrpOnRMz+zFX6r+wjyp+R+hCMnqR9wrsgjWw/YGhfXbo
Z1/zWPtLjRaJ0efi4Fcoy4i5oprQHLoFKfQi2nGTj+jFwsYjaTcbblLZNRjTPk3M
THXbu15TzyZ4nU7kQSz19pssmhAJuUDXdQo5f616RqtZd9hmnrr9pco4EyGz/lQz
WxI/Fk1idQjPYrjUZDw+6EfT/r7SfxLdtsX7N8Xsz+pvZ07t2wZPqQV5dJRxWsF2
ZbeKwwRFohDltkuZ20zZ2iqtCA4+pwZT7j/QfBM6914dWOuuZgnjuCYXlLc32aXl
j30Qz4/Vuk4rn487aVyygh6YEvzkrNwy/DcSz3dbznFUft/7FGBXVcUyckXUsnKi
JduCBdRgenuhLFpnf2IFVnNuNiPAemswlyWidW2IhYYLWiIfbrUGo51UGCgq2FL1
EcYWN6Eu71RRSCMK4OVpWoqetz/RjIx1VRzv7MuWmx0dhu9W+SU35d4PLms5u4kR
WSMWmaeBwY1EPbw2WDES7wa++kACsISbGmyOBQTs2pX5dGwYCcZMcIe8PpaxUEEW
D32kQ2DlZTVeoMawSeD578nnzYzdU5camneIY00iH3V/n5JL3v0hvxvWBulP6+1O
K1I96QhgnZwt5Q5U/QkkzlFj00sec56h8lnT/usRKZyP9Sx7NlZaFGxz9xI93+25
h98yByiTe36eFqwW/h1H7JYq2J0XV0Q8N44hyZa6zZzmVekLyAKHK0aiACLFto1z
Ux40ndC2VCwsVFNKdB7lNID9I/EspydQ61X70XPKnq/9RvkYcSG9pw5lZUISDChC
hbwlOOHT3cPcfLv++JdAkUTZMZosg7h2XCYGWkLRH8brllzOiR5bmK4hFw2WsRM2
WJroUTWoOPlIlsIgdr3m/TTXeP9Z3UjSiGNBTyp0XP03262jpZSzoaobLKKaS061
DMzPcP5dVbGtMKE3lTx6ey1fMWqrhu1TKdLE7anO1erdnEPRMCW9cLo+1n5BJYsb
nRO98rktS+r1+1CQVhtcVX5AdxQ3l5vyaXaL/xfjRK0KmO6DllvqLPKHSnXbZjO4
FNT+qUmwZ9FwXDsMgKEVIhCeqN9hHIzSNNqfZhdRshn7x4WVygEg0TciU7ysSQ3G
/90dz9Ks3CY4P8yrNxp7MJfZKXSso1ndFPINrAb5M34n6LaHBEarGzIUZ0YSlzO4
OJnmR9ESd/S9xGNiyb2/S2jr40BA4ruwvCyFGKEtDwhlh1dj/jyG6bvkmWT2Vl2V
fJM5gnKde4+wDz+PM5Wzm2AdWeHj8Onprt3y/OssYFxCFxSPrszRDN4jlRNwHL90
0ytUPaFWV9pN+glJspdRyA286TmjeljkeAx2ZZObggVxyoP06q9YeMcro0TY3IV5
3Ck0NQGy4cS4zBs+Fe6pzwno2aOybAVnk8x/rGtuwoKtQ54OFDIuj1xFUQBXnjfX
6i/MQISAf20E8RWmzDhU0YAXo8Td3r+1dXgFNsXsfAKSv+5ifKUUIMD+ItZtc8L+
k/BfdLOqFMzv0jkg3OrqS4q1Z76i4skRq71KiE1Bo+csRqmEMMBaYR9bNTfZKvjB
FPQA+8sKEF05EXgDL60yUXSDyS/L7Mv1/iA4m/nZSE3RzYczc6qc+Qygi9YBMB1x
vNHZ400y+aDH675uMVw4qdPNFtQjI4MrlFVEpjo6uxWAnXCyjsQOK4kFZLpxRuq+
qEdqqs+hv+ovCgojEkbV1QAhA0U3ecNMUi2RkQgXnV8Mfy+aCUjN0np+HW3PWrHr
dXjm5H2fG7VMUV8DpmHPmL4Hz8ylyJQduwkoazrb2s7zPFcCBY091qAY7JEVqEzu
jBjpVKbKPqYskzIJgx4jNTzSNjwDLeQI+RytblmfRy0Oe2hvwc5UP5JWnjPSHplB
lDsun+57fVgILXhF4GzBmIvPkAeGvwxOnziuwIILQSNm339Ad80YeBevLRV2ZTGP
ssiQFOOEU1m8L9s+N9NmLkhetM4x4Ss2/N2+q8YReVUVRivCD3KOR0i4OG0w1w3W
0QRFznTPe7XxhUafKAS9rnCumbEoRicFGhdsT8AM2f2C/zSnnAoKUps+SuJdYtED
pZ8Mlc9kEWbowrf3kKVRtMt2Qa7LhsFS1ubMQTWBwsYu4WGkAAe9aHXDl/H93rm0
VzM5Utfaw3/3Eid7CdS2HTv+uo9g5QcrIvJK47Kltm6T3LqIEUFa1uLwQOooOcix
2Y+xxucnMPsfNeqKvQ3JwC8RVaobqtEY+8Udtt635k0xZ1pxZNYXVQAFtvNkH4AR
kr8NQy3FwUWizuyHxnUYGBrvHTKIuEn1nTcjm8VSzZXktFpKnZURSfpHQ9OAlTNH
joFuG7nj+zSrLkMv4Pa7jKHxyGMM20SCHkp/+IVxamfDO++zr/8SQaVZQQlSlv77
zLvU03yCi5E0+qdXMsnOKDfKgC+qMYx83DdbfbW0V0H69xsktcps1LUN3M46XMpg
dt/A6M/dEDVuCMn6n8vsqLhMY8zqSx9VrfoP906PcRYTH2Fvs6KnGSW/JOs9obxR
a2NPKHM9w34vN0h1npvpPY+A6gNt//JtghE8nN38gJdrWC/GV0pEEFUUErstg0/e
WH1PNsE2wKCdj0qZLxDzo5CzGVcqkNgrYla5WLWmqlr/MWqgVpTfwXG4dpPXCYWv
sQGZ7h4KtT+4Q2cOSsy8oRcOBZ7x0KBbc5vONc6VqjxSy+e8UERsv84jg4GanaOQ
63zXUCFLrqpFYWW9FXQv4QR8Lb6Rl+VuI+5VrEzAckqeiQgc/H19X+Fn0vWxW8BC
5RN4VvX1AJUzzK+1qADDlFgoGZvxADrk1XKXFYoW/aHXiBqgxLMGNUFbwZf8ZMni
QmH6aHGY0kyfN0GNCO3IQxoRnOX7PytHPxYrfQWgbqVqyIpXQsN3TDN2tYFogVVD
BXAyCHyFKp7nm9GTaeiRzPAi0JkR0LxhmVI0ByfUEGUGMOvXnvlIf35HvTg4oAG2
HAsZEfKkD4hL93QRfPRrBNrvKuMnAKmZVmftiisxQVfAgQUzMPRcItCu2oFMDY1O
8BS1WhU82hcky3/F1Aj4aXTydz6PJVicNOziXUSuKDVj2L3XJxGewHqm1WqiN8ZR
a2Vcp7PeVW43M4w58xoqEYeYDY5gXYzDGMxWOeyW48524+bXGjtfoaEBJbNvY1hC
uVmcqyL6oRFrRtbhNiS9gNFms87GwpWu9XN7ex5xBaGAk40Smu4voGtDTqtfjzOB
PvsrgmiaBjl9Yb+lFfbj6QNoRzusKmhEGARw+++Ly9vB1/oD5621lMBG0Avz80pd
U3pS2lNkLxJ3IUPNPvgEpWq8ODAmYgepYfBo1cP+VFwPQHCj4wRFsXajUJ6+AbcX
GnT1eTn5c0S3Q3RdgpNyJpGkDR4CIF98SRTBGDU1+A/IwZUoVKheyI+wZe8Wl5hJ
eFHcXlcMcffRc8mCrWyN7v7Auii1CAVcR0wW7dx6KZ3/7jUvayXTMpFnXkGRCSw6
+GkGCqGt0/r64mBeWNy+ls1mojfpo7fQLDRTV47NE4Q4TutlRUyPk1eqA1kTdAxA
m6cLlleaI/3v5vt3dysD8eYLwk0D17i7eMut6RavNQCN/JkruDXVXK18LjrVPL0M
W1PbJ4Y2O48UjXdmfLvLzonL0M1H/rYEkEFhdqMbMdvKrVvMdzoUo0VXdvkxwjhy
k2ntK04vrrYlxYeWMXRM70HLPeSi73yZK7zNZE/9vHXPUVkKB7HjFHhMVcDE69Cy
pEsvtQcvHMIbqDwQs5shRmy8Um1ihRC/t47D6mI4EiAnL4x27agVAo85zlkIymmC
gjWm17IfHUX41RBlvnLJOntcNYahQaRElIw714S5qjfRBe+DQBb7mq6wvgHYR+Lz
o6BoCokEj8Ma/Oi6bYKgruTfcsg4K+cJqsJLoquNAjfTdDNC2+9Jlnk5Whps4/Ci
vrcmydMav5DW9NjZk5gWJuzbx1xLO6j5r2dbHPbigyxFwMFBXx+6LHgp2aYmU16j
prMv8VVMEbvZPjumhWJMMPj8NpNBo1DVIdhhOhzmwJjSZgfc8Cn12/GJzzM944ut
MX3Hcvy5lTSbcNg54L3G7Ay/ZG1ZK6E2/cyawyLT9B69MF6u7sYSkExI6x9yvJdo
STY97TYoyT/uZifDnECjbys1qvoRVksECUlmOgQbpnhDcA4UiwJVfeJRFgQyeFh5
/wQG1W+uxH6mfewdgRX0TxBaRi0a2Y7qVAqyH22smdLmFTSg5Qw6A8vfqcy9jWnx
IFmcIWamOC7jNWDcvtUy0Rduu/yULMzXwV3go8w9jwfKjAXuPRMrEYzPxdthwRyq
f3JJGQ4z9TCfzDLxrvkvO+o0se0iLhixnDU7RJU2mySZnNIafcBrykGQEmVqL7gq
0Db5bGY6HAr7x/Pcf4hNfhjURGvK4KoEWuV162eJnokeyys8yseSVXpdsUELbC1m
3m8KH7iTvRHNcPn6sJ46dv3NeVPy5xKEKi3uzhjXhDfw8LkJKmTupHuednNVr/vj
9AGw4l2J7ZqLqYVjomCFJGgXlf3ENnG7PE0h3nqXAIcMjIuKi/c+j5xZgsF6YgRI
BbQcnqdp90lTPZtzHEHuIc+03+9BtEIvixhdWu14fJgbE+YPXF7DFqKwmeNyF9m+
5u/p5pvld4C3MNjuIKQLD9ghn1zztEmwj2/qjh2qP4Doo+4Sqx59A60ETM2TJyFI
0nr0j4tZsl95zYit2f2m4xHJNKdV8XJ7NKYKYG4V+f1DW7gpt4hAy8euOS1LosqE
bDvxKlyiRY85RcuFdircjkmvl/KE7/5kIG9sFSzcr8WBc/e2LmY/q95l07KMHH+a
kT6MJ9ZEYdgH2cqCg6oaBp4N4gtIjGEIHkkioVvJBYjfxF2er6+j97wSSxhDMu1i
dZFhToxhpPzgoske1KG1Sre17kOkhq/tfCqznhrHaBkuENy+apYispCoTnm7AA7g
z7Tk1rRLt1cpGqXfDIyv3zi1dtqdfn2pQYOCP6q7SUMZbreCETNJoPjuGyIb87ih
ZcnP6OrhM2/W1EdrpL2h3mvw1KKEDCo5H8nBWs+3HP+SxScifoV966rAO+lpkbRP
9zZ562QGoU54m5NKkj8L4bOVB2ypPy/QHfRE/JjhOTHx9RGZsOzRDWcxt37nerZi
b5le23olKghhamxYDA6eEwiGDVj3FPa++D5YMCi0iXPHWYcd4xIVovGAYUDYj/i7
l8nBL/hF9yDWgoav4hIvyk2gGsi59Hksg/KyrCYjUe+5vTjVf19SKeFqYsOXaEBU
dkercZ+1jZvKLx9G05uIYrGZc+VOksiJteR4mQCmcc0+Kq50crbqDLMMVIbdYbkN
ZSjevUjfyAtjc3huBlPRBTOU/V6k6+cl9KhTCOrj5uO/KqDivd1kV/nnPYaDraGG
zVgIn0+pGY0JdpkZJ3Sk1DkGawMh2tPuv9mmIVGyKNmp6zvdFRzhhu+np+TY3++/
FjEOaDUZQrPEYbm2iO9Pl7MWtPlAbBNpyNB0J5GBktMmZOp5xEwAKnLR8/nxDOGS
Q6v5FBTNT6LQZk2vPI1SMnXckntLNIcGJ+ZeKqIlMc2fafwPailrb0CPkXVCMnJd
VZrVKxJ/1JT1e5fJgqHeDQjAvtyQM/uSSv+Sf4KlzsbXLFiMRfBPhod9OOiy0S/A
sRJZ7beqPOIO69JnV+ohNcp0KR3eUOMP2Nmy61ZBik/yJtRs4OR6gQHp/eWr+OvM
Sg3zmAdKk11M4nRf97DHbUWqsIkO0JUZsFxheRV2f0unSxudVfkldN1/qVV0oSPj
l9PtoHlbnkeAhiMTYAtHf3pgi6yfoh2/TqwuuXFtxdJEFvBGB03Tq5n+/EwausuU
rm3AtxwKQwPNUZHS87ucwgvuvF3DIsMvg968/lBH/JB0pIu6mCRUqWRIlzSqV2bc
0i+Kg8DxZr+r+U6tGsW5luDcnv+VBpFxxUROzphmauZzNSAaOKVoP8sozp+V4vnD
iqAptKImIbffP5hHweVbjRnzhvpP8OISJuPSzodwUjMFw6eD6Jhi8wsx+XgK3Kei
joJmj1/U6vS1ImhLUHuT5WwcLvkPhmDq5dNMbW3HO+d8uSjD1bDxt3rPo6f8ESwy
9Lt/4vQ8a+6TdWd7/GY5Ek24jOBpdkKHOZb/cMlKzwDcEB6y624baD9G+vc8G9oF
MA37LcUoJOsbrjc3fz8IEE/Gvaqs5+DGwPOMR1FOJwgrqr4M0Nb0abk/HWpAm1TG
sOVd4xfbmjRnsF0C69mpNHeNpupsvPfqPyEOkj/3yx4vbKSpGVPCNpoz4ajmVQRA
n/jPNdWazPSRhdBzANi8A1MY8oXkLSaIApgFeFXjyuGrpHdNKWf30Acps/wjYDCc
7S9EgB+O/n3Uxg54tr6lk+gs3tbkspfUCED1UrXLEmKZTBd+aQr3+LKGevzbYDz7
Aui6bXt/nbISZv2NDb4VW/UAHnda5Hxhjl9kVQX6JvVM5+cWl6iIUED5hVHP7UkX
7V3BGvsc+iqPQSlpIsGNLEQOubWQsQXsPgFwRI9MVg1ftGKx6f3UyN/U4Y1Xpce3
wfSFTMV1nwvozXlER2WHXoKVsVTIv6wrHmI7jFeKidXlC+22LUFeHgIqfrRmJFt/
Wzy/FwLf24+oZoNsM6gs0xQv5zIBfw9BT3mzehxFwrTpot2/lgJueBpjstkDuHFG
MaFVdY6ZnhLyCRTsneKoj5w2KZ8d0gdxDoyzPZb8QdstSNEWNJT5mDbCTusFM9a1
gckv06W7eEc9NnGEOptLxx0rWUNZjSd6jyO6nq/vGxz6nLZEZ2+bA9lANe1KoS8k
clNfSCMN4to5xUfw/c6AscvKnAv93wq2xiv9KyFfNcXbSKTLzjNbKGlugZzU5yTI
iHccHDflllyJeDiKVCfWtLCe03Ub87knP7AiaPgyko043IhU0mIroU0553741aGL
/CcMmypQKYDI6WWC82nFbO/M/QZV0wdCSptoNAvdEQ1Wc3l8Me1LHSIWU+QTjhHc
r0QGUsBA4uAQrAoQgaKJNWfma+bAHPQW16L/8pa9e+4ujDwG6dJHKvOA0q864wCT
718fdIOOkTmjJAa339YcSgp7vR+WBixOYOlIgeN2X1AIcSgQUME+gnkMNaKmZNtd
lvKjkeROe9ExOCSKdj3hlnq7/XvYddgpiWVJN2Rwf32EEWFp9esA9qWRthYYuZI2
8+5+0i8IneOxg0as+EUhoM7bnVOSFzanXdgi44WRuChJVI+E4ev8SPoosy0raI6S
ux/unpYYPt2zo5PxBH93/gQLl6CeqZqVUyq3SaiPsGkNfQCK8AvgMIuNn/rMct7J
OacqQeEXW8d/zTWYIIOUSEWhwNhCjB5TunTyL+4bG0D9mVVILhhrQI9Wfsp073AP
mAN0vpJSHGFhPNEAxToa7XU4zuEP8OVMCiLKvqIKh4rp3v57W+jhv5W10XHg9kv9
B+brRkSgoIlNpd4wh9/5Mr7g8IWa5sHXYpOCVxckkZZja1sSDwmTy7nuG2+ra8OB
xyDNTjE9jlJTNGhMMv4PTFGF27mPBEEePiobYZiabiMH4wYEI5OsrfA2Gnxlk2kA
BeVyAbXgMm/zV37qgGbyrejTdAY59rVo3QL7yGfYSyE+wcMzjL81ApcFZscE56v9
8lt/u/8t+QOpfFJfvGU3bSVZhJ8Y5bdxQ52M7IbDyRTcqxYkAiBfq2qUeVhSoGlu
BCLph2yefyyB7qMp66DCJeQp3fQJg0HEyUPGiFpESmJbpO0pjmfvB6aSSIxt8a9w
9ZAUHJRjm7dlkUjiGD1QGqF7GgEsmA5l8etUvwBtft6jwOQDhbYssjg/kRmB0rno
ER+R+xsqLzl75+6UB5Pk//eesbWH6rKT+mv9ZshraS58BrrFKvvHfUMprO4SQNSL
EQXyfK2ZQKBXh5gELPIpnpRf0BSeC1mvtPVz6EI8eJmadWQAg5HsZwalMgZKXlDm
UYHc/0PTS2GZQv7by0HWibYolK71oA6cNKtGIM9+HcxmXT/OhlpGjG0Dnoefqm2J
zB/+D4VVYnIi03dQi75bYS8D0D9Fekok88MkIaBI5KUMhsnIJKgJY1aGT61gsj+L
soGPlKfyDiyyO/lQ+GMLctSxYiCXDkADDG+FXw3MjkP+8yByycPIUuy0+BmV1IZa
wTJ19kRSwkLCbGmihfHNFxLqRXIUIAEOHcQhhWK/j1Cnp4vxcURv+lx4IZDVd7R3
BcasfQcL9SuQrBChU7nOKXmA0q0kYv8LQ0TSqLvrzeqE0UVHHJvrHV0I/qpOsQGy
z8fHbxN7RAiJmmEIcgPHMjivcrWBJAm/O53o5lj41zbQx42pdUvVcaaKjB4Do0MW
bXryegZjUi7J3U2YN87RtvE5r5hC+5U0bIiEs2ngzJ+HUjJViRJ+dRKyD2j9ZSQy
XvQ/ZOYinNN/ALuokQxoo3JMrSnVGDskGX0tZLZB9FNkTgBZl4SSU9oouZnsrF2U
s1MDQQ4juYOGm+bwEHTHiEWB0qlpud0J32hXYx3FY7cOdLn0MzcwmVD8hA6EKuXj
CuxYqa4FDDyIotgVxNqO/oqClrHPhTXn/xxm4sd+WsKC0K9677zCoL5heiktqNyt
k3FaPGMxSI44doruW/OkwLEQ+jSQ+Q5Nhl0ZXUaQB3z8nAKAnKKqMipedptNCpOY
PgQBZvzn3MQOor50v2qWvofr6r1z+tKZXRaMLiamIUyhkEZQnx6i3ii9263Rp3Sn
IcyKjiGaqicldy0WTAW/dJf3R3A5rnXMA7hZ+4O/27CXp0qOd9FiDUftr8DzydkH
EO0DdYMrryATEUP2Z8Az2bk9AkSU2jJs/BRMaBopUOrXKkc4lk5evSfTBDEqde1G
p5zUy+7V6sbLevecwOFk9Tqy8jiNgokn7kxSqsIU/Puasy9x/bTOvQYt56cmynh3
CbYv0KRThijHixkvdLzzmnlrO/Z+vIk+hTvMebH7O8Vy41mGWvn2/+3lz2wJkvh4
vdVONB1YyBFr/oYuOo9XGkebmxvcI7DdP+/3ZqJZe0LgSV1QPOMhC4hd1qxRiNBu
6q4IkXSrCs+1tZ6dcw3fFVgs6+hwQSCIofEsOec5dPEkuq51GQS9+LQAa9zt8Upl
s63nMcFivkSQSeDu1TfUcQpu+QhQ70rWf5gg509SNBCJN1s3DYYRkogrwSOrdfkG
VfqMFlN1KmGREGKA9PCwG1XTsg0y+8NlGsQKBQCnh4Y/KOWLFQ5FFjs4Iw6pBb2O
xvMFHk3oyHoCVabBl69ZT9ri6sf9XFFOEZEwvuZkOp1HlbLQU/OY8BTzt0PlX1UW
jNmdGoYZkNAbsv5ARJhFqBUVOQk5THfbLGdXn17Umxo5hePxf1PZ4bWsMcJ9hESO
1w1zYWR2uu5HrCpoq9AYbuys+MGPQ7DERCkxOnkE97LrywzY/7xTKucPimdX3XDi
Xsm4PGMERh2br5NtLhO59RPWQqWq1fdcJR2lQbtDJ8kenlQGbNf97RQO2GOSvh8q
NzpCxumiKZgY3xWLF2TcdHcGT3eLUk/97zI0nkA6USaMkBkjDAdgmduHr0vurcSK
TirVkHqBTk3C93gx7Jo6l3MQt1ZTd2BWdCTHImCY8uUqMkE1ES22iNS57re4MSnY
ga53BrM56CUgpnpyXc6NUys74Bjv0pYOBZv//QCWsO3k7zkmjwNhQve1EAAfkRd6
4BUGJOqpzqKp35C0hTdZ/tem96zBLVxpupu5UQgqRlVdRc7ecgG0lgu/BHFqjbu3
4cL2Nn8A6gsv9K4TF+Ty9j+I6MfaOPo+z4ruXc6j+f6lVkgotqFOBF7c74ZcuLFJ
30Hi5BwZHbHHngjHoYUj/ENkXje0DOJFGazBICOrAkgG9RmEcOpwOlDDoMDoAqOd
1N1MhyHlSW90Vh7x5oXX2bKUBa1zV4TPW52FJRh+wD00squaOSIMpkCBy8b9MpIq
3OjKJAfDoBaAmrwTtv5NVKs9zYUUb2jfBA5FJ5llhaKoLMHjfMeY7gkx32+j93Ck
wL0rIGNVrFViDWiMCeDbLy1LjWhDJUza1rPHw6xhU3xGkLpBTNm4t+hy3szBUBWE
H028dVQescH7WpNzwNciaFGxRs+wj0rN38mpJjQCT0oYFpk4LGxf+ofti4NBqQRl
pxueH2S39e41fJ5h1/FI33qiACAte+UP4r0OzI/P8y7sFiRTNzKqkWQ7bFIa+tlG
YZ4xJ5mKtZfak5evMjS0wGg9lSPOcSXHacq9R1ERXWXfwDIj2ksSjpLTpeCpfC1H
Rj5FrxlTJyLiCwBeJvGSx6aj8X13K9lgpVGSHyunYwiEo8kdf64wXOS7Q0DqZ7tB
JtorVSKm9DzVnZwdU2vhWFP/3iUhgBjFLoabCoFZoufxW1cQwbHOr6XX64c1gZ0m
AwXCKpJaba7qIKAQ7HbkvB2ZLO+2wx3If6SyewPD86ExouaHDXFud+ZKGnsGXY3p
aGRKPfqweJTXVIt2Hhf9QxgkN8DDOGIKx8hudjk4dx+BChYYXt4RM8+br9kvtL4G
LM4dwW72j0TdKi7TCtdqhBQXXkLnJdUl+Il5yjtX/hhCzm96Q7RAee44f2LQYxlZ
OkI6Ar46Rj+PTGLZgHp0y6iUZPIrrt53hyViineLjhEVbcpNqoXPsY0i3wLvytM/
0IcSd3/LPj4rIu1sSnqRHcYhJdtM9TrrCHacaw6/hwfacftutnmJphEN7x3EuFff
78VbSK5aFBOaTSUizAdgaDuwHNgVJLTSIHWz/6s88j4Pe0zKcFf+1nV3EJsjvghB
jbRuS5IYHUkWexYDiuUNj1eZwR54vELwW2/gInEyHGYhj1m+ZUdWJuf6yp24yffA
LFjgOYq5Yez7/Ct7AVeuf/EIf9I0Fs4yDIIdqt4wa67fmA9uyTZVPqj/6CHLavDW
BykoJDS7iOZ5zU3SZejHbe031GHddrZyviwRY+ncMVaG68xoFaPFjQbvaVzJ7gSl
tJiBlUHsjA/NZS8QbvOY1KO/TYPP4Rx2LUdqAJ4NBQuzBxLiCA6ghjA/ZLKuUOIr
Ed/kIqWiOAx5uHfnuP3LQwghUxYHAwiIAfZyNg7IQCJsbL+49ArGd9/rJh7n1wm+
ihSFX9ZAQ5ICb8+5ug72JwkuZM4oabufCvb1sEVRIGHLykvSee39BKC0YIz/EpLv
ND0L3Go913B2f8pD+ZTMsHnyF3hu1UzvWhG0BYDSb+8eekPL7DlvA/+msIWcLX41
nP8kPxTfSdKKT/I8HuhDg4OWyBqYAfOuDR+6iivsPcRgIJ0P4jWmEDbwnuYZTmd5
5fH5xf74zODH+PFFEmlWAayYJtlCQ7TDWO/ESjr9PxxXFbGaJEXljFEKbCiI5b8Y
QC0+bFt8BJAo2rhQPB75dG+jFoRLVzGoEiMlGcyLu6JbT08aLr788TR0hYxsrgHY
lkbZBOwcdPSD6eiKBV/RmwFWq21AWKdjRAT0b3BXh7CE2baWcGn1p9kPj4rIYQp/
PQhFTyfK4qKtFuTn7ZApgGgza/HYEfVSDnJ13BP74Jiplnc/Gq9DFiXmd7jEg5uU
wX3sP9qfnImnFl91EWkmwm09yWJZDAiNFiukB4cToyCXbm2rRkj02uoUflEmbLo6
FNNU0Gku+sTdxEOvUu8rpKcmSh0hq9RwF2UqmrWwv9oKSF06yrwKcWerMBhL6MKW
fXCtppAEJ4id59GLV88/qdfzIs6PfO4rqIuBbl9L7yICB/4CYzwbvgjcUQwZH9Hb
hOhVKI295vZl0fjxu8GCHbY+ApKTCualEDBi3fPydjgqhoFXtx5fnlzQZ0FIora1
2ZxPxsKBXRHzepghPsdqGWWT/OG9yEl6ubmYpCcG7WRAAMBruNVUK/eROj+C3yss
eMbmTQNzBkl2EPkr+gMNR/cLo47zeTdDXzqWPOdTJTzugx03zlpUBbpA+3tIBdUw
xi2/y4KlX9N78aGMntVGNxX04lx3FH/54J1a+Aa/QBB3VeqJ6PlzWOvOe1rpP8iN
R92ZnZMb5OpIW8LGi7B4ik7CYJ8ePn84+cy63DcseXtBMwj5Ctk6okSGSaEg5xmC
IWxxZ1mrNgvMm3qdGRpuAOrKMJVixH/8ZTlUKA6icnFbw9PKduUYfI0aRjYd2Du4
ZunLySmlj/nf5LWtVLGdS4r7Y2AZIUXrr9WmqY7Iw8+tvH0Z6yRCy6K8Bzvne3KI
ydfxG1PztQpZ8oxA/dTW5U3ZRduaNPUffe7TND1vSEcBkK0C0HkHfCif1ObchVnd
7Chy3aGmVb8vxH+4oEjqqMxqnq2TuOMbKGRcBhl5gKFKMfRnXe9vCB/PDkNhivfu
sf8t2l22c0l9zYuQ0xPRK4mZi0oH5gOO7Sa/ysBNqQKQ4tEMbUvywOf5kyLRLamO
nhfyzqqQNf0gp91qo9CRVS1Yr0ikvXzu2CEDc1uMz19+LM01E+rZi8jvq0VjvbOO
27eouboiJ94s1ex64T6xbgTIC/Oj6Jq7zp7cpL/kN7uyRJf8ivQqfkH2A5JsVhe5
7po5ExLfQVHyKaT7ZbmTXBO+u5ckzYP1zGQnrfH9V9GIdQPpJZjzdyXMyo3wy9uZ
28ElhK0H0VAPE+cwNlTlysZUXOub32U8WvMMNZSr1iTnfR3yIFKYUmklwfc+HHcg
6p2oHcLchi9zE6FXcwgYg18N/0gip2nvYJZjlFwwKAwxpP84zX4viwjwMENrJkAS
/jR/4pM3IzuGycvZpza3pZWQrQB7BRiocYTWHBFuxYWYawhF5SKY0S1JPN3UKx5/
TkKouauPDijnWp7a550wrFZaFZW4nkA7gSbjbtDwIU4wU3WG8YSeRr9JrYhhC1aP
MURkz+7yA9lK5vITVuz/0EB7Zb+NB1KwtjyjM91/ODd1mX4y0YcBCIjmum0AycOh
93qnyNNZuE2CnYXjAhqZw0nZ3dHvXvroTox+wuKuXT/heXeyt1gOyNStDogwxwDK
cYD0AXvsqu12j3d1kKNwjNs8yaa6dUhC4iqRHhL7aGD/TMAsYnRIhbPNBJmohYl/
yTDf9LyI4i8jpjq9+rfTa41gbq/IaEbwqkQcAyWgN9xqgQGnXtjAsXEwmIVp6Ze6
9pdBzkEe6rWQJwJ3PtnaB1hSPZwMbhttYW7oRGtNfOpQ8enQeJW4zD3sww0aU5rv
7/7MKFJRSZUaugRsyExUW7EER0YLv4pX99lHhNGKK+QZuMpKhSh4yfl1/D3IwvCp
G8UodIAOYQIkyYRdVl6B4OTfq+izBjFYd5+6wlhk55MITGsoPusW1Wq0WFhRDmG+
DKrvqTzoqKY4fhGQVV1uCva9Iwjlp2AN9MmORhdGLY92wohSNF9C8jPzFDOwfxUS
v6EyhDtLJ7NXFQLLwzU86f5oFwudGSXzvZD1PfeNOW4PrEPlI8cEWs2q45MS/HlN
SawDLzUxIbk5zqtBq9Vw/iQQBzZmkza0O9QXwQlMuZQHwNFjMDkt8u0T58Yol45/
KFz3UraM9f1z+yxS8bQ0jBBLE2zT77Guk9um+QIQLIYTeBo9R/W/UEH8Y+5MZVWQ
XxKULhKecTNDloDpUibinPNogvYaqE4rUuTGRvnnWYm1xdQztxJ1TJZKx913Wo5n
k8PiOJoEnWYTwjNmxduEayF1cL1Ly8byoDpU4SY9qM7q4yCEmEoJxTIz7Vj74Eoh
VOeOTnJ8ltoFaSKP9QIHwfm3v4chqPW3dXeI80/xNwd29egmpKkcfJC+kKcY/f84
LIJB1Yzj+Y9kGVIWAF/otX5hU+8Iw+x8ERB84bQ0dPJkev9djnJ77uwIMev9HQTZ
r75OvFtLSNCuDoGRX0IRQT2s7ixqEGAFc6jv1O0wnv79WKfKqXsK+0NMqiSeYkns
4vMYeOde/gTBsgvehI+Ecclg5phwV4R+ri7XNP4slq6iRGakEjnaNwjE2cfysdfc
juErdvVn9Enayttf+YjLGDQ3/g9r8IyXoKy+qeAoYvmUFDRl5mw6S4l7TDa8dBwp
/bbf7eve20po4v3B2qWojmVpRUg6lzVsMuCfID8Y7PaURvEDpileqcvLHidbD53k
azQanr2XCyvCAEKQpQ9jB6PPdL3g4wbTZ/5ynX/vG6roevOkvQEuFaH6B5dWQ/dw
fdRq+R1NDYKL+pmg3XLLZdyhNK5WhYq1qDbrWUV3LLkSD9Dkyeo8008Sh5jqwOtW
Ag+enuwlO02hHkrzwK6XLP/L2X9Z0wn9o1k5twhiw1SungepPf/9mrtzE78CGSWs
odZr9lOdZuH+gJ6M6Vh9S7GPedRjZihKQ61t9ogLgu+BqVwbI9g8CN3LyAWBWEyl
3mvWaPNF1oNn2xgkO+Iu9z+x+Eqr/C0CqITG2Hifhb6sC0EdWYSzZuyX/2MiAenx
ZFXUXyB61gKYcqJt1tuVWkPObauK8eH0OjkqXN8Nf9O8TiKYY42oPkx5i5iVtGDL
3sr09yyf+S3pUlRnCqDFRqoK6GdJkDQ8QvbQa28NdqLG9H4ssZZ15h7x3FAPDBfz
YFM9/avUzN19TFEadDSn2LxiNZyyoyK0Y8XKC6Smr1/weU6LBA1dhHzgkXjLsuA7
rwLxRamnopRwYn32iPM6LuoALs+LzdRyqalBYlN+rIl3dcq94zp2ArSbDd1QEAw/
1jjTVEXEJHorYq/3x6XDEj9JvCKT/jKwUzsyzDV3dCUgiP/3cxcIUs1StXcd/jK1
oDo+ZhKQPgbp2ThqyidFQkTxF3KLwm7vHB5pDImh5A+OzuG90br+NFS5kzhekTpf
N34BXHF/X76++fgV+KwzfWir9drZG4n7josmNI06F9G9LXOMDZkwKMxOcnf3qr8/
kUVsxCRjjtXkdPtkeshF6l0dQk6qnMAsuFVfq15Zl9dbK47JpBtBds7eYvBFaQo+
HtMReeyq0cXVktVNm+s9qmPW4JjgeeCp3Y0azLafxj+qqqT/x5jAgT5eLgySllQr
79CIBUian+mUBZQyV/YVSdakmb1p+RgSV/Qe3cd4/mAoyk/qjkInwyQX07mx4AmI
YDSz08XfCHgXFsXYpvmUdF1MsFDSo1pfc/IR1PgJ/71MOTX0pFHpUMJyEeVK98Kk
c/MmSWYllGeSdkJ7rmzkm2csddwxbmFhBmQvUtk1VOtP2sQvVCFZ1DPNACztql66
odCwxoc9xSTQz4vL59Q+LrINE28g7cSB6c43tjFeaHj0Xb69GnGhOx5tu58AkO10
eFaIWU7jwKGo3w4sWUcwzc9eJMSisl5mm3YKDZ9wey87QkxY4CJi2bFXcnL61wy1
QlsKtr41kqZsUMHVIt0iWgAscbtSfWEaSrzqcWrYfDfJLoh5f1RrUc0K+ZkgrK+S
L2GyCFM/EMtKe8MppVpC0d+Y3qonXlpVoJ8fQQFxPLJjjxFHmqJPJYSnsZf79BI5
ZmwedCmpKnBB5FAppQhg9zrDrfwjFx/b6d5qpWYLnvtCgn7GP8CrRDWmix2QfRWk
zGNz77hM3c4R4gqm+Oe5tTvQERS8uCVUAvfXJ13ACdQirI2JUx97pGoD/8Y0qOIa
bTnuzmpZ7k1F/A/IXnPqZ5qbpkB37mMR2cbc+iEp2NY7f3NxMmZovoouppZPx75g
D7q8HyDM/cANfz8z4iAeYzoZMdvZOD6YV/9vCkEJPITSuIHESQd4E3z5zxeBSG75
Zv5cIfdd5zij+h1CHpjeIcg8Pyd6rNidtn2U1dUCW77MkRLjrUCcPYuWldidO8Mg
L5r1z9TmYsssas7oa6PlBcUe1/Yd0fSS39k9HhBRBZzRC5ccz+kkD7m2cxkQRk64
QJNcu4ozSWCVRa2+9dRJgNe9698iAL7nRTze8V+sfobvXPshhuCioz721tWzeEXD
31lrTD2pX0xAbg1HxDqmMYdNiV+hP2H5MJ8CxBqFtRVQEvUnQ0HI+bYjfAtdqXWj
6lmZUQhnfaBQvuHuNt3sNPiOCIJ/4EHoihC8kgplkN/1XsHht9YeMhfQCoIKlypJ
vlQzrY1nxIVAInsbB2+fcmBkzdWAGIrYNxE5XxnixowARstTOMOcCcuGX57sLbcD
lfyLrN3PsAwWBRO4jJrvLZ+IKW37JOutaNk5Tg0NGMUYCYaH7/OZsDnNysuZ0GAL
eg4swEyZtBSYIffUcxiKBtLOorITNIbInQUW2QEsWweT5U2SB7cKLnLPH3miCBxL
3+Ms1lPwPXm8ncsHI9BPNJZJmoYSrJ18oSn8vSYm38CGD8KtNPNvUkukXIBwHUvD
xNK+BierTSb0YY/jImkOD3B3c9nNewkoRhQxKGRc9WgTyDkLstweZwUXkUmM/Mvt
nuUN+zTS7wABd0/GhAQQtoclwcD9Z8d9IAqPcuWCTMGS/hifLUJFImVUxytU4L2d
fVKfOcOojAHnFh/qSPrb1NboQvzeoyekLenp5x126GzDkpVx+0EdMarYG03E3L3D
2uBcMVEq2kgu7DyINRwHiN48XBJ/FPSio8nT7YmmKt8Q7sIxwdkykKz2xLa5kmRx
xLRsDkoOkVOTDizCWa2kwpBiAUmM+3nZzAiZXeTz0dzhqEnazIJpyp+oVhFECxGv
51MXwnUSm82WbvXzEfutyEug9tihExD2MBizUIQLt7ZUcTdoBVq++iiLMubSaB4k
+1j8TqqVmllzDHG0nKV4MoyBThve3EsjM+1nHzWUrwewC+k4wYz+Zh5Y9llIAHLR
qj85ZsVKN7a9XbRZy5uNSyD9uUpYqFV0PFM4La0AYRScNZ0ByClAWvGoj/juFnA8
dL4FvghczgYvpt9Tt6PAJkxd9qJd1orhmXoFcjCtuDwcCfomvXk1blw2m3br9BD1
q8QC8vmT6SKzBqSpLvyIoCQ2wpPxSQ+/6FPpRtV+FWMnd1MYX2U2THKqG08qYJL9
PX6q7t7DyEInSvkGYjQFEOwo2yD7QyffkPgGZegUcA+u3hndJ74r4eBOl0lG2k4h
zsActVEQ3zR5UgnBgQSPbFHy+e4qp1Unwz2SIpuy6CZt/hv+1+DdH550ZJdGU8tV
LxS83iDK0kh2MxXJ5Zx9lu/DjWqndED5229dCGU80VFzeSYKUh79U54OA8MlrFqg
OVuFbiUeP4b9lnQr+b0hwEciiqAqlK0qRQPK++inB5i544lhnSI3+a5d3pP5tpcJ
C/IsZvEVKeUww5f1n9U+9f3lrR/EBDFJMTCioWan/ZfvlqKmjZwVwCO+n1LuTnfs
ZiWiynBSQHRE6zO4KlDcVUTcloMhzv31CPL5AQqwX0YHleJfDgo1GwFYqwSUhJC6
lZRbCpqohohmXeX0r6luI0JNSWc4Zka5MRzbYLPGk4VoZQ9GjHeoH/g76WVEm5jU
LoBnswvHhQURjqWVMCqBz2hyxfT1EpwOSQr4ruSlSUatV6N5mPnv5XpKHEyvnXgO
9LoxQYgqzL+Lp0xA79VZPl+sMazEZl0Hpl+lYwEdmAFbHkYa2g5bE9Lu3G2DdEVI
I8JjsIpJ1Dy+KejPkLErZybxK3k2LC6/CJrE/vtLD4S6iVIFa4hwINllFfwla6pA
fQrKANuAuzQqZMdNvouvudSgzUrjNYmdokMjiWi+BzDDuEtK4tIxqZoyBZZ9HIQF
9o/Wp598Eg++SfV6k5mEPn8NcRc4+x/Ezm54Tw0AwHIE7Cd9h/k6PvGCOUzZBxpF
y06eLAN6sSnnJz935Qq3VYtcm2OKyrlsMFrXWiKL0roLLErkN042BtNuhDuL6527
DJBVfB0m96tCQXnMyicGrNDqkqkkCHQ+nnBsHD3upG99Xga+MEOen40yhr4JI3zy
FSu3CeXSzd1HxAaKc2EZxqPVq3aaIMIj/xtbsdkLpgekKcp+LFn6Cy2HSLIs1sBA
Df0vte2OlazKRH57S6xUPQvPtl6x3QzXaflqTBNdL/eWpr3IC7SnDLppPXftqBV/
EMUukJT4zXeUkwKTLyHZwZiaziTAvP7I1xEDSQDXKr0ZH20BZNj+x3h4VUm16WQy
7tb9XF4rWDPCE3foOs0JAgHGCaaqUSFu3bIgfMXv5+CI0s8d9kk24U24tEx/g7ne
5BWMCZoaMlUT2XalfCJ3O5iPsmdJiFB2Ro5IHCPTNvUhzVSg6zbrER4AiaM8osds
OWBwHn5U87uwVi1kmC5JB/r5LlJpbqM7Wn2PL6apkyiQR9csWSq5patpy97ZeMWz
6jKF4TUW2FGd13QuLLaCvvBOKXS9LVceZ0IJhwnvwZkx1fSt6+Iqd+d+kiyaPTPJ
vl/oyD3HCpBGF8R47hWH77fSRaqxGqIkB7RYd45gk45qXdQuXODybgo54DXMXyIL
adoVTOAibDNGc2hj17uEFb6SDe0EVJkdnFpjsaKbJZ/Z+d3DqQfiWFcR8EpPGO+4
+1vJ5SaH0UZ+HjwRXH8XOPgLPZMvKlv38MftQWFpGEr2SNs3rJ2MCQhsX+70sfS5
lzWmp7SWA+6gXz2Zf65OltlaLU7lDVYTI+jWMhbvtsgG/pxyHfJbpXDp5zqS7C6Y
2S8MWoncls8fhv2TPmkYn4m1k+y/uPptM48cGlT9H/jExQNOWWIutlaFIAGtdJYG
w7M1OA6T8sVvVhsPLDYTnwLTl+OKW3jG6zja5kcc/qW+laNZWHFbqnzjp+9IUyx3
YoHyOCkTwUbOWZHt5bU6U9sQf1P3cIgOGtQzHAoHORP1qTJZE7SCrdmfEiRIBW/M
+keOGG8/dWruwlmIc6B+8vpOagCtN1fG0ApivebsVYmKA6/xa7s4QX/KFprT1XUl
tfzuLKC306Pflmxv0BCrsYnWfRY+c8ZklLLGRMciN8CFgan2TJUREBiu5fJqxj6G
Ge8nnAYkRX6mEyeqQNnxmsJmcGMB9k3uB4f6HQ4AHjIU6x+KVIFAbVshC9et/F07
7DylXcczOvsBes2PH/0pFaZLyoCP65OdnK4sZ4pD7Y7VKMvp8gDvfhilwRAUmEtP
rxFwKiF4UFV8JREoSv79TqBtiyRPPLMo6JInYKs2p/gPTmomukHk4uY6zS+j7WNG
ZqqzeKgE4bt8SBm2ypu48fIRnMu59nopATzqsAa0gNEovHfbZ3a5fHj5LMg7K20M
Ewx8nmNA7F8dRkV1+Xfk8jY7OWITscFQLqr1CfkvWSCN0s6orRcZZMRvCpEQPnL8
ChEsmH9tEnqHRGJM9Pc4c5POTZ9WIYNd4abTzwPTF9yz9fSFIQOTvL2C2ee9648d
KCBF0T4e8GXa+spsCSTF4MOuxJAGxRf79wBq3dhZPrjdPlGvlP9oWWgkscwphBBk
PmePbzOlfGZJkXAVJ5NmwyOGc9JUCdnm9GTXPgh2BUY0GJHy5V9qM6pAThuhYA5A
esrmGCgbencQbadHdjxblLaWCuCogmq/iBvia40DA695guCsa3Ww77EmkMNv3r90
Lrig1r77PHFfjnNSvbMtly25E9xePrPRTKz+mdtpF+LcTM93WpW30scwuUz4xWlS
mqrh4zqzj3eCk580et8eEWZe5bI/EX6mOOdzwZSOKTa6xYzUwv6flZwEfPHnBI7V
dYxh09VHfPUPQzwD9/8ocYFZwPwNA5bpcGtjGJMyKp976nS0H+7g7diQilDrxocj
/5/Gk40Fx9qFTkDjG/G9LAiMOWDMAicFl4lt4DnMUYqcDAWqorMEdhPvLL+DCBeo
Vj72NYt/tKryWpDdKTAcV85LfhYO7+Mxxf4U2XLe/hfgQXbrpB3ggVmWvhOpYw4J
qSyBxYmScN9VR7qfvjoW5I+QHque4CCTTDppDWJ5lw6xaQD6oyBGhTQ94o8/nhFA
O0tc3VOfExMY4df2ZqdRFeh1N2lpwL34dZyxwO8DCmJqo3N3JePlHPjeVtxuyjRw
D2Ouh5qXXeYGDyYYWl8gzNHlr7l3yRNgWsZR6ag4SezE+cpRssF7Lo+jzcOSWQYK
Hlcuk2KbXknL3SoNrMwxi4UBpXPvPLuUU6LVbgx9mRuLp4J9D+UffGCS27duEHNg
QreVU4Thl8hielZMvIbKCAVtNY0nb30SRlX4P7s8xIkyINUlevBFrn3j2Tm2n2fz
uCmvE0Inhv5JrPS0m05izzLAID2v3Vpj6vcr2gYPqxfOVcaMCTPek2Nt0KdYu7JO
bcZUlxanVNS6bUc4gzAoPoX8gDdNsexPAj3q+E8CsdRMrErvH4kpSQ4KogZ28YzM
8Of+9jQHQJI5yfNak7KdrbUQVoMBbI0N79tW2XsqaIKW7SigG9FePC/TmJkpZURK
quMdTXGaD8ob95pcJyEvwJVSuUlUbKD8xGpfW3hxm07Q+P7XAEB+fuk4riDQ2VUv
voOCE87CpSFXCLibncyN4NbER3s/KriubQlfMTHJtwBaQBU8u+8voX9pl9MaCb0F
ngDtD6VyuTuARf3j62D6ywGiq+yqT4nPOAFqJmlcf49fNIltDvcnGdglPUX9GebQ
L0yzfXmrusdnD8YUNaIkfx10plLFg30jEB3+ENLMkWyMBQre/HpYu+8TsPw6o7J8
9qt9bx1jj7Bb4Vjuqhe0e+tbq/aaBpTp5ZurNMbINf1fCobsddYlQgapmXSpTAGx
ka5pYgUzenR3eKoiXXAqSI/q1+YrOw+NSq0TMlG8WkDx0tf+1gtN414NkWnaZj+y
iw68fqrNHlp76KWcAMS/MfzRKjyBpoWxml72hfHHKCeKCtLYDupPjmodsGQVujX7
AmHxPnkWQO9SKOZLFDkQKBrWAJgVZOFra73r6y06Iuu7WRoRRESM8SpXBQAp2ORf
kxFcPXvi2/F19NLOzv4jf7/sC/xrR6ktNQDUkztvbs6oLnI4isebWAytFmtSIzW8
ca4m7AHETz1fcQriuDZEwXUtUfYk/g72S9cuoRmV635WJKkiDpHGMByAKwB/TXoq
BZwwuRk+0gwjEkLzTdPmfPnols3ybzlqr+90EPXeH6gYBNkzx4jz+ZcszSwyTAYn
1LxnhcRzAZRDc78TH7SWquYD0jkeAy/zPa7N74z1JpK7hPyQ+LCf0aLjyx1xbb9d
Z6nHjqXMu6ca7g7l5lNw+8Jw2FVgo8ww2SMFLL1KRzBexPnJyKtIcVi9MZSRmPhw
Yg8w+0ynzSqdNTarqgvmwkTLAjoN8ZTM2eumPkU69QEq4J8SxlY9GVUSO+ysn8jW
2UBOl5LLQPpRwEarGJ+03CdufuhQe9FGJdlyGmcaMzHc4nMbOMbLF9XN3OyWaV38
9Xihhjr5P/FHvp/GKvh5xP2wuVBhEtQfI+DRTXQtrMbBlibMNZmganV/ByuBXy++
o8AHHKiTalJyCuwXx6VYNt8OkvC/uSIm4o5frGq+kfEDMY6hwDHISd99XIDWs+qr
92NxSAyZuRvYPnrMgasHux0YMpwjrWeKjXPB8RPKwpXcXqf22z9GWbElaMz7XbUc
d7k5oc0ArOIrqD0vmXzK/nLo0+PdVba1aWZ/y5oRNHYCnfUc6NjKLQypmtJOHVh8
TOF0L7RdnyQk6f9fhqhmi+PgaRFKAMd3fD6BenDKxO3mVCAsC130tsiXgeN/LvTi
s5G0WQgJ0nZBj0WkUs8q1o3DbOSex2bQD8XX2Qm77t4jCBPrDA16mP5tS8/ngDzX
W0uis/cp7AqH3LM30eY02tRQj2DlwS86DUK8FsKO9vuUoMiFKO/F2MBFjkf4H8Zz
/A2xUxAdwRiaMu0aeUlLDQ1YxJ1Y4D0dYjg8iJVL/oE7nuQdeaMi1EhiolL87MBi
lEnzciIgQeRY5v8pv57w/5a0NfA3S3c0meUACnHnozYQSLT/YPyAWXX3nI5bqvjA
SdRdJLSSvyG3qHU9Uv8/wHPtNws6ni3SIk3EF38iJdJ7Ht29K8/IewLox8kZGiNC
YHp4QxEQnASPiW9mVQEfhrBXGYDU8mV8GEJZh/1mOWf0vQrw0Fbe2YDvlwDKe8Xi
R2kDgSgTE4q0qkARoKpTc61itW0hroYXhf+H/Xsaeyoe9YSvWfNccm0CYqkK99eX
VgaddM5plz2Hrq12UR6KfjOD+/SE6GUMKD2UXLpk2V0wFYYgjMygfDKoBtvuLS4K
Cp/i106vL54AHlIUC8UDkc0DTENZgOoirEp4UWTMzLA/x+WhKSeEv4PfoKm19GcR
ueYtKAyLZEeJ9LFfP4NI/+pbUTSiSjFXOCMIMrTCWzGSg5IzCPasoxhFucOQb12N
qGHIdY1rxOrpi3bWgiJ14ZelJ4Or4pHOy61iplMgF7t19e9w9WtIAde3SDNVzKDn
vKMRL/NxBr2XXOisLXvovsT7TSYRAgRtpWCfJ5DjrAysdSME4ANxDvWcqh5zZTEz
k+5XgLdtP/JPi5rUxhJZBUZ6dEUS/yX8O4m9c9zSFkxewUOG6umYXL/xQjEW7d+I
KIA9Hk6wufVToPRbRM4Di/gYwufO7DzDrbsz1Xc9pKS37dO6+bPZ//6WmX9Ig8uo
boHBx2cIYvytDJNvRi4xKvUHmQ3aDeHiwWT+CI5jS44/FSClzb8YGRoZ4Xjibqbv
f8mA1ZwXAyZBPysi3C4yVThxyfW/dvTBC7WWHbkdndM9ngKC6hCWz/bfWaqfHa5A
SWa5Mfj8xneu0ceQYLBKU6fWszAbcWwIZmBOVZzgE759fVJnCcC5+5NLQfCucV4Z
56Xr1eiUSJvkB2WoUCFBh6K6tpiwrr9kZitfjA/bB3ujO3X+uHeDw2BUtm+CS85N
Ivlx/RODDMcDD7vvsAjudYVpeJyg2PncjchsDTVtm5hZVghCsK60X4dQLRpp5wQr
Rfb9H0O0AqdKJNd786uY4jpj1zUN5i0fU+ZJhtFCjwyrIYZueBSHD/ETMY2U5SId
M5AU8oUYq5rCX/KNPeGr3iLGO1C8dtqGmf0RmiXjjWHRfTkmjqJiAFE7nLPGZJn0
CcA2yqPP13evvsIkWyOJsq4u2FgSKJBzK8zLCQuS/YafN6yazAnO7GAMMyaeYk4R
4dwG3NTQASkQjfSsk8eqIl7F+XaV37tMz+0vT7PAEqqqjjc4UgUssmcxIsKjCOh5
PkDGsVdVyNwzvfUee+KCW4crRAANHHC29f59V4pAjs+wDHWvnG5E+/ENuKChLoZO
kf7/gJDYAFHv8U3N790dkpHW/X6FRwLTCjI/yeXK5JXEJrfUO2jru5llid+FVc/K
mLuxR2fxviORLvjKbqrPmJSKchf2zsD3L87i+zJyjxn2uLCzuHRJJA+xY1trkFDi
MtGQ/cWvn/ufvxpO2CUixm/16c5DxnkKlUysJmEHJ5RkhnYulCuXDwyAOeRxnMBj
gTQZrLi602qhsa4SSG8Idrqa8PAOZYFYtvKBT/GvwaliM9ml00NRPYIBbcHsA66R
xDm5hwRg/02H1+rWyLiUYLW2xNjOWDRDwPJUCPeEqRIvOMm38Z3Lln5T/Ob9DMhi
Fs42/dEnDD1t13sPcOw6EbhSasxFJP+Zw0+KsQhja+d6pgBOVNpaSzNW77V+Fu8h
9sA3QAlsMuLzqBjRLPGVrsC1DnW3xmCbMcwJjsFbIjLbfZcLkCyGxkAvwu61UODQ
Yc/kG/JiHhVoqAeBHWY9LvuQUhdUpXwlrP36az8yAxVBKbTVUAkzggzMR8Ts91Dt
CyE9z2k3P7fLaVpo9A+gkluSK7WYIhSprJQAuBQQmTva+PMiv47r5qeb4ro0Oofs
/mHTygzEaQx24PL7JNlvd4goiVIkXzMC31G2U+QgD9fpiocRokXXu8QHRrTKL2yO
gYLSd3hQ6T8KFIgOhdc+ZtbWkEx39V8JqYHVPkUGCioYcSwFmfeez24i7bP1EKWY
JZNd8P8AygX0OtCgvo1SAQbL74QQSH9E2gVfcILUdNf+bqW27K9HDKfYKg0zqIcd
oDb3fri6vRDaBqARD7w7wf1glWJxYhMEM7DQAIZblnH9NmPgnBNKIMpT5sGDj0qS
+hZPzpjIqsCTryCK9rzPHSADnAnCiZfuYub8L7tvAgN7d7f7piIAqAcLc24923K0
gTFU9DRD8HaR1GPvplFM3cULcEOiNQBdIHoJBweHvtgS2YnkLMEjkh9RMDyuQOQh
Ew9iJyWmCnE4vnHNR+PR2Nm+crj9iJwQiDXoNOV2wiz+KfVrhaatm/CinZlIA6nf
RCcjcUnfoUfNYvDgFzkNfbxAUVA/tSKbdYQZBqaBS45TVjTJD7FfUObe8I2foWhl
FiVVTnPNVt4EN+Gg/hqCMaFgCDZyHyNas1CXqgShJc/xJ7QDK8Yak/ku3O6CLdBD
kulWJZ61Pzp64UJXVoyRD3O885Uku/IGPjvwhWfi6DrnfCXalQEswyNU0V8yfbAn
ED7PEK1CpzJTBQobMyLvV1oC5/Y2GqmMiQOM+rnPZPyB8GvopF/jLkiR4xh7J54y
Zl16/wo6/gkSOatj9OSVWjN8fjOCDSWn30HPGlGLvTBnsJ51A9+SYQql6qbCI5ua
XbUVg8Uj7DBTegFMPLHD3EqOJktTuLe+Tk2vp730VuFurswnNS8C5ikTZXTeZ+53
rfgOy4PBlb2e4GZdncF0SOnfWYABwmz9xgyPFZd191Px1InGS/rgal9/KgKgXGJg
sPamSAgpRF/P0GusHhORGiv0ISH6ZWh4Sjgvlff207bI77Ay3QGPwj4Qzs0+zOjn
zPGmqnHe0sP4yw6Ojy4rG+eO2IjGkSb0m6iEKKVLtpQUsuFB4ZI2voM4+sT1tLkP
cZVq2+wNQgi/TIlaDHa3mTGroiQX5B5h7dp9mivaqtaO2qtZZcWTcPyGEqhfRQ5U
LCWUa/gI3QoK7xsDWIscGeDMUw49TWHTgeG3BFSMI1PTD66olzSmWoNaAtKQA2Q5
Qc0197WweWXeBzsLPsSUevEKpePSDqt0GuY7Cj61XXym0MB16fiG65f4JhyB48N4
D6oEVp/66QLu3hktwF8bunHxnVzEe6phr5k/HuN3j0MRyywSEQi92mbRzUkbtKag
ip7GxkUvwuXLsPqu45pi9lDoQmfvr+Hij0cZOqPFtrxq7xsCmJZf2nYv/I1G8Ryu
MiTceZ7/EClt/Y6v7bZXqLbGdn1ob4YFQEEnRGMf5tsaDT91BvpZ0MN7J5E7RTXL
Bi5AiMASxALvzweSLNT41dCSqFhZVqfE+nBbgrFWkQuAe551ASn7BSI1ntKtmPC/
unN/EsFaOSku1HDPzgZoYSeP+xA8oKfoYs3k2rlKqaWc6v+12Ibb8huibc9CV3no
YURI5SdNWlhS8zW/kEv7rWQ7vnQALlmB7OMXmiALlWsUK4am5JgNCZGXdgepeo1r
9Y4zL/EhIOmGMegJuKC3vnF+fHM2bFl3COV+E6R7LgnyHnr8GGa2bLyv/DzEBVsl
pzEwhI6iGNbtIQUYFOwxuhNtZDBai81AMqvDoMyBVZz07Xb/X6L+GB1icfJlaSds
eV2wCG31wtARBeO7+vIuD3cVEGR+BqNqhS8zElJMw/IbT6hXdlVlxTBtz+R5dMiv
tRd7PKu0yJwbjkdiLin5PRqNL2HOl03P8bKhQQcq6qZNOyxc3eMd8c12z7m3u15C
KMEWKszAmzZROlXpMBAZx0rcBxuEdCKF029L8RFpsQ59jKgcIoAF6ja+QM2gXIu2
NlWTN4OR/xEut13yYcAnmCcMvbt0ckk2CV2jgvaIF7Tcc+IcyAItlnWlENzlgIxD
PXkFK5NeS/ff+ro3444a8QPBi8hokMjlwURtLk6lvSuhwxuY3rV5fJDfm2GFcxAH
+qE6eC9bd2NC+F/BK9uK47BOS/aUb7nPuIybnOwzTEy+nH0MmT7b/0Bo1T/x8+ow
yBTg4nI9dbt73jShcf8ilshwOacvg4CqdPZW4TqTnRG+wu+do3COslizN7cKelFx
FbghZUieyGsRgmIyV3+98NDdS8/KWhDzyBiPOWtH9uykluvRTA4wQoLpfnKReBD0
Fem1uCy3MYVAZL+1C5V5FkUj9mds/Xih27ICsXYUJu5XLWMw2WeH3SfQjTZfeEwv
UkXBT6Llu6wPe8vQ8YqV8Meleb+5lU/qmnN6Yu59q/ksn4nznOjKoVl/tFiIC6m3
WxR606qEcFR55eqxPHdVCQimiPJ+MV67Y1iJDMDgIEXXnIXqwb9VkCvdpU38xCLM
Mca5GvExW7hPXUzitaQ4b9Se9u5Pbb6JBQdrz42z5eequgicA4ZSIzD0vPMVERpq
iwYryvvREV6SqODBzctB+DCYXZwgigUUVw0b6DsK+zYkNI3aW3gzJfVcaE5QSihZ
L6TmVl96GAzPHnEh0HRQsIdAGuzRplTcdrp3JBk6qHoc28TNYw3s0DNhpVIxRIzm
OfmVp+Ihpf7uc8GF0cajYzCBoqcXfpSKY7WjKeiGaQUf3GzRYnnMYcXJukWig0oA
1KVQ6hYBRqFTxXQgj5u2LZb79wxIU2kEEjTFqYRyUxk8bnvV/hdFClIEBgQ1Hvi9
IliiV63f5nMTnaI1ByE5rUP3eIfAJsc//s8X/KC768qRRNNbq31dbMTQcSegG97w
aVPwL6iWHihohSZl+UgTWuhRqjNloHSykauaLYyAzc8tAUiRFc88JFQqoDPvXxjF
S+dpIYrKgG5aPUHxnH8pUKtE12QrFzm0sDbQpWoch+GTPPzjnz24WPefsHxlMOhS
cP+6BzgHmoGefZ9xiLWEKw80wYcLTwiHsf0ZCjGO9Z/eBv1vTlLolRmiuLW3HykK
50ugHKjQ4Hcj+/VPhOL+UpVaTBusMbJwFVzP20JEsXFeKFhY/mWSNMv+7ZIP3Ujd
fS3yKyZz5RuVqKeu5gU6s3tzEMYqGBPs1R7GV7tJne5GY7ZHX5PczPPa5SAnxX3j
6/WjI4D+mdt6dC1SIV5T8lx0/boN6Yi7g3vYR/ILLkabLAF0jk+M/k/qVw5L8EkM
y1F/CK6Xp3ad0sRTUuRWnZ4+OCoB3wgwb5+AGkKBRrV10yyODaAD6+856AzsqY9k
wqc4BDIEfrnEwbqpllPQBu+PGIR2hwkQT3mO/OFY6qmpcQcvsjSAqycYdtzJ4QrY
KWZjJKdA3/KZIN8W1Sg2McOAt47HxHXlgAewgNM4nO5KnHRrXTN/DGh3yAfi/Ugr
JRHYWGsxCbtNNoXU43RudL0YZnllECFIn6FJw6eYBRx0zx/H2q1uDtyDEwD2yEUR
bgtmY62ci2Pmt22aoJUoMMJj8VNKOeY3yWZl9zXSav1Ybfq/rmtv/faXCOT3w2js
aSUoLk8ebr6/F4LJZH46zzV63cyG72viPRYPfC6k0Kx9g3wk92ij0R/qd7/sehVF
uiJ2NzvZMlM8G7dFTpI+glhSlSXmojIQ4Zd4R6umfVDLDe7iVBgF++9eBjXJLZn5
72h1zjLZvEdUuLHzX6d4iU0KbqIiYO+ZNSKbu5mO5eD3fhrZJC78g6XGykpgdsa3
1FuqE6PAun5KU53fNAlAkz8X9UUPNU+iy31oM3hKkBn8svgvOgnkQQas0QQ2f4x2
LTXrFO/jq1hr4aP37Js+P2H0E1u3H9BH2QBQMBI7qK8cCrpGCi5jPP/ZoDvTdcac
2UymeRpenl6vEsmho7KqQ7IlLy8Nr0z5JQsbXSA435qk/tsdLlZzzuIe9eut+XCU
OkX2L5m0OfEYje5Yxz1BC9VtdegPlLqA3d4guuTVICa02SOfNYwBScFFKf8oGAG7
iUHR++uY4DHvwFOJocHVCE4NM0alg2wNGTC3NCkE3ubuvWYNFzfba0gj0n2f7uTe
ucP7k868fcMqQD2+NOG+8zc+s4su4zpuhuq6/MR2TjUp54xhgikHb845m6yfKJSo
c6Lkac6g+DJw4EJB3qUWdYD+0egFIxRfFmL97HJ9PBHeLrrC7PHxH4wvjF2+/7B3
P/CD/kMK5oSb7QENhqvtcrsFZnuig0KnX54mjwW2M23e1gCLEPrcQNawetvKHnSs
u+8pdP2glePkOrKKOfE3n6WTdWKJp6HNv3d8ZBn6u2Ndhh8KVRTbLppY2ZY9MCIH
PuTSpZP0CF0xtnUQBe/XdJeCLz6YROBQSS+ciaW/YpoEiOS+CvfbI/txb9iGyEZZ
/4Im2jcOn3Fa8VP55JQVIBcO/UXQaZIOgHLeMW9zGfEPEBTKDUU3jkx+N+tqCxOi
jL5/9qPPt2jtfuvmaIh/+EmbBRKs89xQG/zXe3wW6/v8Ni8EzRlPbcEUFRr/7Wlx
hBT3gAB7FSLLw8Lf404uGnF47IyIqeKyDr4cYj4/ZugMM7pVI+JD+QEYrHNAvAeG
gc/zHK5n+Q+r6pBt+sv1paJUQMPluiavMvldubzXNMcLxW07QGd1LKVN5koUvDyR
3KvDK54ZLzvSulQ6cs90+SoCsRMLVBjqXURZEQjWQcZuBcJHFibk2t+HE1hVuEaq
JQ3/J/iee8OBcIlgMS7uT/h9xvdUhqg+8g8Dy0Rff8bH+fJKZ0NUAp8zGX8rbKeq
1tBfR0tdrcOOthV5wpMcWkE2u5Kf4g7qf9AYt5Tg2jC530jWio75BdWUex4S2QoK
py8fz8nnP3Nd9sxCs329TkrrnZ6F9eIeb8CSk3hoHnFzb/CU6dcFzich5mMatPwE
TEtoFKSDf9Zd3RXdasGCxF+c6/l/P0RNeOfvkQ1MwWHWknoqq52baJYdXMATMCFJ
cnFavgrntYEObLpmxAFQSrrpByEbjo8MeNNREhxCm8bombPLNf2wBI1Q8YfFwofF
xxQtcUzA0G4AFVQommWqBSVwyKxIkE6XHr4eXKhFCKLcf58/O2YFHviyVCmJ0mA3
3pPdMuQQ8a2iGIpl1knO3jemOxjDNivggV2cjol7QJ1E7KUWcmJQwIpPl8H/bDGo
8/ZsqvmjzHBQ5W73L49iXoxTZAshQ7GgVDOoYLfRp9BlMCU3N4bW4HUzUvrmXqJG
PxtBaWGkJdVhsEmnjext/fAkyYZOutEMGdOQinHE7ihNF4Kk8Xdq+ROaEUXOPMfp
mLIL8+vVrzIEzI8VGIxt+lOV3/0InFQ5RnFRMvYe0W2zcOhFh9BXM6UJtDS7sfG6
QnFQxdZaELRROrc3aVulS8++EHlUMbwZcRvunQ3nT3NlERSLTHdABhj3sZqeKJZ8
/gNWqYuoa3DyD87gviMbL4JywSrfYv23JoriUgOUjlTJ/th19l7aXXLoHowknIBb
ZXngrpQmYZ0pNaTIWQqk9B30I7837GejkiMeWH3cGwvi2LkbacRVHZ649EOXq85p
MaGhOgzAShOciULs7z+tqTj8R3SfJunxIH/IozX/aulKLoOrFF9qkRIyUsZwIPyp
JYlSwKb/ayyrBl4hrpFrQK69FR/0lznZuk+U66wN3TlW+gi8d+vguxss3Ka/7Nxq
QBT4BqiFramwpjtnRggyfQ+Q2a2k+vGSZT0UfOqcIimTicBnNBRfv3/EFp4WkXM9
+8+X82RMXN/mzXH6QebFO2ZzSNJuEPLBULY7WfRtmIsrFf5W/GoxldAzrf4shD5+
ehrReWgV0RyWMe7fg9ESdewv19uYAa4Am9Xyw6f7s+7lTA+uR1dqIJDMjPhrE2ME
TQMXRQjOkn8HrYJqFIQgWBdNqCQ8ByzyZYfsEd5qapuX7V7jUvOU9FLtVgs7lpSV
DfWOYlAm+ggGRXZhQI4KuGrv0ftEu4rKJ3vHf7FgNM0tuIcwTUwWhpKifhOodjsR
iY+BlPkYkjxx02g1opu5gub9k0hXbyEOoqJVqKw5i64eJjAMo7AHyKYhmIUnCiwr
K6QAbd/xFiL/dd1CDE+hWEakgGpekzNcwe4OSq5bCGMPZ+CgDvyhc2OZOvTTvtLv
kVEHlbz8JSfjvPesMq485NwlTipSfU1lYfVLLe6w+yx6XTvlByYeB8bK4vRtf0gu
42zBBmt2jXazQ4M4QR4qtTOjZlsTJuu0CdbJux8P5RUJQaB8axb/K1p4oGLUGZc2
ulrPHlRq6DdUOxv7G3i0+P6tirdyjbkA8nsGlD8j/3Oznrd/KVTzNHtQ/TjAGdZI
ce0mfOJcDtw1YH1f02gGzPo4YqGcSREs8fyt2kIkttCDHFZpcYIHQljM23xKYOxk
fZpqt+Sbwdzot9RHyIh6cUQApJ9/V9XaC6FrJflsX1Wt8Xb/kz27SorjFe5aIdc+
qw1Wzwy5yrRxyehaIShifvJvGGaILVceLGS7gd2hckvErToE2i1ZVK/Qfw0di7Bm
FP5BsZldEV5it/HFF1qra2jI6bprMDQqpZOfpIGNdqv256DTYAjisM04Nj7WuZTI
0Y4zP7tmc7te8/tDj5O0MOMsb7eCWjzBztx1mWSJkI3fBeIKjAUlf6L2c3kpk7Qk
BEpdOq1+m9POVFROwHkOl44CwSXcTOzQ97IXHgO9zDDEt0Jde7CGslcpzx55kpAJ
P/ZOTYwVH9tDp7GPZQFbO5BGIYebed6n/Zu9oW8AOIKs9/i6CxdJLgS98OCYlKW9
OD0n8QCVlYEIWwCRYTSdxzHlgP1r00RtZZeTcibvrC08WYMJ1Iro4Dk1FNrOMJM1
01rHfsdH9w7pH3lW1KeezrLYtSs4pAgfD5MHu6r4wbPpLjRFB+DvtQEVO1bPlPOJ
ClTB+tnIpykPwrE9K7V3FHIioTHPhBLMwbEajlZ5xxru0sxvWuNR5t45bBcQAGlV
ONKMlrrDd1gHZg0ZXT1mLX/GQVyljdxPg0+V603p1/WvBY61wPQCJcDEuSHLBFaJ
yH2qp9Troh0Ce8YYsgoTRsK6NZ6LBBBY79FgB59lo2QlkBtDEdO7bhb2chYi5mpn
XxTeFm/Jht6yy57BeqRPbvU0iwbCBr5bgf2PbJszxJErVnQel+/QEt5VmgPydIFr
+Xi+8eHI4mn0ZKfHNOKp9z2SS4gXbc5541YwGXVFCXZl+NRoWwStOStEk/pdRPgy
x0GPJBXPUVfhbpFgsBzM1O93zd/+wBkeof23RWnkXIG9KCF7l6i7gIoaUEkTOUX7
idltzSu4RZ0e4qTWBCvTMO9Xx4fkcBVLOYmrTprio4VTuoJG3QMdFrbxoMvEdejV
0OJg784NOtu5nQLaiRv5dTA3LXOLGLoXShCWLdiZcMm/Hui9xxZO6CCbv3U4BonY
eErWvEdq6/EAq4DCTGqvLitT+eVPBrKIsRdmHJQkxbBY5f0mn0IOqXp33hnIirm9
7nPYot5vvf5Ga+jhT6qPFs9DXh9Dx0rzCtNRgpqTuuNXwT3uRY/TLeiH+jke1VKf
weaIO8Oc3VvvB0gpqV4EEhbkPk8wMRFFnTanaijLTlgw1ArczGZvNomGEblMcL+S
k4DV4sMSXw0WLS6w7c8pCqjXzjM3PCeHaHIu0Y/McV3sqhd3HlFr7V5NDujvJkru
FooEHsOgRtFq180BU5AGsMSUex1GAspcjq3vgiS0F31NwjsxMmW9PTt6qQqek1rX
LX21mJSMQWSDnqwXPxknh4CumG7XnkTrlJXRMJMi/6qeVtXQab8FBiX4U5HkYaVq
zvHaR9/6N+ueTpO0SlTk3rYGxE6VspftHdFlYpyYshHG8RNYL+92pyx+ULDot7vV
a1pqz1QaZ0mgJPWEHLHAq7CU5bVe7o6uEbDI8wvEszkEdBoiyfJg7iY0qTEmk75z
jjUKr7/x/4RAkeXKfUgWrXWVvFsr0QV+683mkcwiNppjUp5Qx3tWWTE57NYaxpcT
JZ8VziCaujm/CKUfuXNrXGazy32vW7EzYPhQduBu9W+RpYFhDoC+T5Y6tu3FVp+y
1qo3BnCQ9u5Mh+YGSCfv19hYtJMiDVWpoFu4Idiq5/AR+osd1VQEceaMyLRlKaV8
ASZCqkylY7R36YNzvHl9BOak5DPN5TtykZgr3bFUku74bsaQjvmzcBauSuxr4xH4
h3tscsu5i3fcIBjEl38OSaPKA75i4IL9Uh35f8B1XO4mS8MUkRLwcW0wxzNLs66k
9tquEvfhOasp3Qg7liRsJQ0Tewrorxeu4eq7YfcV/UUvK9wUdIS8qrk+XdPOOIVk
KMRr0rJlNtzcIjne1VdvPLfwjbvH3tOs3DYNvvioouXLWS5uBGLNh5MTZcRGZ1eu
ayk2usq1c73HWEN4DzslYeuWYNDl/MbzZs8Ip6aqSG+7eIUyD2lKBiTRQvkTChts
sESpQffawAgIbTYJssqbkAM2TZmi+8X72QamgkiCN3DDxI2x0fkplZW5Ef7qapL2
X0k5J2dDU61sfkvLSulKBJKKsvICLnnJbRiSOfre0rDCVlXxCbjZLnv7w/UfSdbn
4785UrY0e8bJG7X4+qQnthw9GlXZ1u9q0w77xlIYY1l3rlXREllsuLSmZ/3b8oFx
YC/fc1oWIGKPEN1UjLmc4EDH+5nKQUHZ0xQeMyOFlrdujAWGgkRegow7/gdy06AI
4E9clXM/c3PwHIOqxDYEAc1met9SLJ7ghycHwYEfK+BFTuFT3f8ukagb4S8FNrkL
yt2omLZPYt6Sc1KCBuxMfP6ngRDY9UYshNNjdLQZrlOLLW/9nxwfrGOprXu/dsDc
xF0wcyQkil+3A5bowV1GnIbWrXFI+sncOqsxEMPVn4G/aWLyiXd02HaIuFKx0ABd
fOPvCgbHaIpgbgEYR7qJPRYSGg3MnyOxQswJOR2cf07v8ui+CemEnrslZg53qBvc
fTgBqJ4ztUAjhBfGYEIcrQg9bhKrrGXxsPnc7GWYQCP6hf6OQ3kFMFp0suO2PQ1v
Nohq3LkctsPs7gDJgE6pe6S5GLz8g6sDLoxkixTYFCbHm9q/CBNMxQrHEbJ1N3bF
yoVa1yHWjYX9ZIQZWCCt7z7ZvdkWw7b+r2gb9L2KJE7L35OiK5q7YG+CX+1q3aUd
RJfOGTF3j88paHNuOnL7VqfrzoEM/PZwS139jYr8dFLnse54Oz52Nrl5ye9JORT5
Mon2dRSiqfyUDVvtxRWSP24v93r46ovD4+cFjFwB4zqAqSrmp+g/G/a0JsnCz+B/
Z9LF9GrBm0a7DbB3fgcH/LljGaAnjneHqhupDDmfhkMHURjAuXs1FbrQN8Ybx+FL
snVlDBjSAZuUdyjTRqbepBbRfwLbPmM9K4M+YzKjwhhQgg0qw7UFfuWHfPwLZ0zB
JuH8s7b1SvKJXJ4uxy7oKa/b0VwwjpTZ71owWYbUd773y/E2v4hteT05F3csHqU1
Rxe457x7zIsBzYsZuXahKR0j3nsQyn+SeVzPH2C9PUtWURvSQ7zsgpKdLhmscEVL
TCmj64HP3RZ/Pe1ypNhfJVGVEhNWJlili4gTmzwcifWduwvpJr4WbURzIwKgxoun
iWpAWA/sGytEqGPjxJ/oiZOJpuungo45LjIB7JFF6rj9co0m2Wh6xBIdmdOPxujF
joz5Ivwzjdl7WgGY4ln7XUV5CHR1AsMtyaMHowjCzdPppVg8vujab73gzFCBp3mX
PBWNHlhoblPdLPl7mziN/Mmd/+OZkaagqiiD12VZv6MxSQOWl/18YixbFWmGnnfp
04b4Pxmy9x/hanqv8GLfxtX7jZhe0z4Vx6mJ6FEUfkw4D8bZ/ghw84M2mbxTCl4M
W5Nqk23QRM0yD7Cd/0N8kJiw1uRt52/esJsrm2Iu0ikVuFTVPx1Wn6m44BLrKDwU
oIXC3Vt/wH/XAlVtIA8Hpip0a39cIuoIWLcsjUhaNghc+zJLBGadpTrJDwjlbJQo
mXCBu+ze7X0OkOmbKx3/svPtDFhMnMY06HinjTdliMlDRp/SY8iNiy8LSVkdjq6M
RCFblI9tLLtluflTjorBk7iGSsf95A7kG8+cYD/FeE7jrCDMVtr3cQyZy89eNt52
qC/+F4bQdaEU/RVVlsbMKpsWGVUPprpwjG5Vu/y9egoU7VaTq1R1thn0LeBlSkpq
4SiKmaKH+Vr85GVXIah5NI7V6V50Oljil25JleSxwqNv2A+ffD3QxQpD5bT3LQfQ
uBQQjfg+jxVLWazy5UKOwLqp9TPl1ruuv47uLtNeqr0OjBthjovuW0cQmJJsxAuw
qHR6bAR7QXSx6Lrd36GOrwwukhQhhnskgyYwVru4Kz40QNcSS27kz83pOSrduAGf
d7Ef1UvG3zm823C/eHMwqaYr8oy8arqRO7UX8Xj+ouceI8JAPdJhM9AdAfcibZDx
SCG+CFg3nyrxitwZsDWLJXoecKWbOg+2Zns2YmJ6FWUH5XVATQrZ5YME/y+gF6A4
GlUWPQsG8/MfASKu/K2SjV1fTDf9QpDgwIuQ0t455gdhn6L1DK+kple0uQszLYbh
CHVb2Nm7rfBzPNhBTnftFwYo6rmOCwhNTQifKNHER5Zyqd2uiMvbsFWZd8X4SK+5
mCogsQruAnRfZmv8whtVbfRtpyDNN6QYeUxCps5waPM/5aO82/T10tUopRrSDCCJ
YsRVAdc6Ud9N3fR+/lmo2eyFbnL//UBlPHhq5H+ZIh0ms5nzNUMTJnZviMGi6X96
jphcYs1vaIzAmuHmlBhqwYCZuF67Fknb2+GD2a6miVLkJVvvt198nFYUAcAGilus
6TtpnKQ4gqcapF5kvWB75hX+NlO5+/xv3glkrQau3z4MXkn2fCEhhZmmOsNFwM1+
yYcbaNQS2cHFHIbSydxoUx1+bVCX0N9esrOcovVD/uAP31fNFoApcpDBFGJ6sJzO
OIdTpu1+511hh63O2dtzNd8KHiTuHkfhwHlHuSVuiLAyTv+N00oZ8lpMPUiyiGf4
85DR4U6NBGgOqgFB+QPPGYLVHtfjPURwX43mH6tCPy5cNt4NEApdUpXwzIgrL5P1
mMBdxIID3Uj2FXDRfag9/pkNxLXwb8ALxDNDFgM7b+h2ZuZtzFfLn/vNbhXwLTeO
M2O7tAUIKTwGx+9fuSpB+V5CclLl3kcu2QYS9N+mWuoB/q4XSoSzkMpuLMr9Rnc0
x1alP0lX/d6VAOABWAduUFcw0sszWCzkoMckbcLBWjVGghBzkTZgzr0/HPndO+Fu
eHeiZ68DVCsnNAuLM/YBIjR0BuPjFJH4/ZKmbcWlTRz+Wu5BrNcI5EHQjJcVED+k
qFYmARrsTvAf/JqT2+wM64uwo/NQvIxYl9x7C1ncgxU3PsoQermlbDHCLgEs7DGr
65Pm0urgNFgRcBumJfsCAxWOdugtTxEM1LHNnaa1BKtrRZKy6KaJj7XldngKZHZe
sEhzFSS1TrMkF+rm/ieNs3F/AqxOnnX/ielAYPtAkSzJs4VN6girtEa38YKkEPac
j+tvfFSZBQJTIljDD6W+sO3aPlyJBRYEC23UrQizcr6FBoirn4tPrhm5263Ybl2B
LwG6p/4m18oNYPM5TPCrbkgM91lC6LgUtLwNuFxE6o8WHC1VKlKF63A+Yc3KUick
YUb7MnKcCjjKGWR8SQrCYvdOPDpEQS32ZbW9NhcnsTNuGN/5vg6klkwTxCiPjm2V
DzB9gHpLip26GtJRXjNGiTtzCAzPEj/6Q348NJ6T7CeV8TaXq52w0TAcyZrBqnco
+p1vcsYjt6dzC6gXC4Sqo3KGksJwzPZL0nEsWeCsnMgOGJA1ZZ4Q02wH5T9uS1S8
DZJyNmdbAWS9/WKDBeLeKVHJHF5SNRVWdufSCu5gp2OtdukbwXqLMezRjh96hW71
1D3LEixSaVzaz6cs2I7lQo+Mp0f/NfQtd1yco3o4Yv7rAUEqpArKxer0nmp2/z2w
F4jlrDqsAi6pKmTxv9JV3duqb6eM8siogymaIDwjs5hZmvl4eGl3I/z2EF0oujVG
1WWBhZwXFRR+kY7V1vR4jSSacEfCjaN0M33KbA/Y05a164HyytXoVhRjz3uxHVDv
FJDXql6dj/4IwZtktVlWnw3V0wTNRu/Fq7YLCCFesVErx8Nbr+ECj3mHJvvmnfwB
yJSQt63goEdTm+iAJO8V7zJpRI4f4SK2QOGVXW2yhiMy3wNwR/vee0uG978sDhJC
+86Wwdnbw13un4AvgAoIjTWkZ4e7ldOz0Tv9Pn6wV9lTm4Kb1r1onL2e5rKWKnA/
6rJOa+3lVcdZui8Y36KNDSuHPNhYUZ8N2sPLTqu0Uih2e6GDtps4TLBraTS3+p6w
eoXUmur4UF6rNDAHftemliD3gt+GtGnwl2iQV+TYTkeJY2xdll3xWtAPeoFsvahR
IFWRDPkYq08JhBcWpQXh7bS9gpo0qDdqHHsouWPBEQPNs9cEiGwzYSo9Flwq8bfy
xfXQtRW218NPW5z5EObiVEkHMVCXK0zvvTbofZvxsx5OthZUIN4I5cmGj0HGA7wG
w1EeyumJfyOpUlTDFNWydxw6akJeAMyhVVK7ZzZgW62O1kmFFh+ucqp2MT/uGsj+
cgZfeiw9dtil8OgASyTdRKXkJGT/l85VTH0lm5tMD85GmrIJ7Dzr8bpPe+KYh4uC
tl8yyqqIk/BxR8qewh9e+qjeZgUCH32iAmKSC75Bwe375rsGX3dDy4x0Ktg/1Jux
z3P8TxviHWLhSI4VdVhpPZdDXtidfozoIYja/VvPvj1BlZSLicprGiDyZ4ZYOPWU
0UbFzE8zOF+UIwvRL2A5P0MRD9XNCUxwwTGY5j17vJibtfSNKXA73xtxtHEixHmD
Lwe7kde9hE3fM3MlF60Fj0jKKZj6uLh93iWWH7e/yGncVAN5B4amrSoJfcigpwLw
ChAJ4qIs1HszweWGe8r8TAUrTYxtGwVRZ6By76CtZSYEPW1x5IsTdN54NuRvHNkz
k0BbThbYIzm4OmiBgiwuPfS/DPCVekks5I1h7wO9NfBH7wHBIfJsEydHWdui1uRK
W9qlaD7zqVDEGCn6rFDQGx1Hew5SabJdeEruBdyev55L2I7QvPAFOipvjQB+Uef7
BaLyngjKgK/xL/UT1yR952WSLeza2Yhj6bwKWyLmYIK+KDUrb0Q3flOBfG5kJ7Uo
uSLgNuatAKW7m1Ev6+LVanisv3V5FMUWOaLnSmlUf5BGBLqZPVxPQtqevI4ti7q7
/PFeE3WotUzFzQrsJjBI1BNW9DGV3OpZZVKM9NkICgt9nqUNQnlA37g/EMnUixH4
5rQkPCa9hFyqWvrTBmSpgYXalQt4rsS24AsjBwHJY65QbmnK23sAsEWYxf1qWQ3g
onPMinBlD02NiTKnnTdZS0hHpLbf/zkil03f9MmQmNSu3opEfdJjJ/EMkVUMAR3Q
wDzsusAxtwVVZP/YnjlOsQ0DkxQSEEAdUWyvdSwL0U4O20hyU28pWubNyFosd2ko
W/GcOfuy8CmltZm3oof3c78L+WH5Rxh9P6H3ZgqgCP3dzHmSiT8nl5wzZQtppH6O
DD4J42iwdJqeIQpsf84JSPHBVgVwBlzmhSMI2obLJwnI6nuje4MTkXzOK3uVbnEN
RwYyt+/2nBvzCUPrGHeUHXdRQ9YlKT4ursiOO7QdSc1Xaypg2VPRz7d6QElmp84x
jhxhYEUEC8hHSHJ8ZU0d62rRV7rscO7YK6vEM9mhEUtmAdjUMYxZ1aLQXPXhGrnR
4zJXdvJ3Ipa9NnejQFbMJqy2nvN31Z/HCz+GKkfIPfACnxBhGqBvLzkAzUQLlZQk
pYKPMB2kOuMuGSf0Vzq1t3xMJD38m8WGGV/q1FdGTIn+I1ERQ8N3WwlQ8WbYMIKS
Xay2zxBGzUVx+CbbY0igYFaJbFvvmg2nr5z0F1LJ+jPNY9kevKCAVm1HGOeNhcLE
vzSFKt1idEU3G/JOOT6/XBlPYxyQ6tv7JdJD1TYCNM+27N41c1wGgC9mILraL9Ap
WZdlXyAjQfQ+SWfuM/0c3i5YxYtQPM4OcIDIgfzVFJHYMjzJfe4n4MmR2XIKE1Au
PFR+gNWRQmEn7g+Ee0Q3koKxvUq73RD8E256lt6pINCGFmB8vT+w+y/v2OyNxwBH
RRYkA1J4Xm2PM/av7/zsh5fOwkIoGJ61k1tDKQW+tFgbFerrhLRNvNHWP6PPfKav
alkkKkF/y4bjGDNSwJhStK2QyAPE2iK6Sm/g/eRpkrszyyrp3ZYwgF3RqUWvy8lI
huCzkaA6mTi4PKLqHH7j5V/0jTluR8H7Q8OZKYsRNct2YTIMO4BaZpm7QpzBJ1hM
YjDeBU9dC+0xmOE0Zut3t9kQGyIeYwGTZ8ZawwqKpKZVtLdyJa7/G5IYZoaTTUou
gq/AO1fODU9YpTs2fOq2Jdt4p9z9+RnWKT/39R+nhGUGg3YYjH6OTWyuoXO4NWYi
dMKW1GjDUGW6kL7hbGxahUq9LnKO1OmUJfHMk1p7abhJLPLFuvvqvmnst9YDbzM/
cMAKJBE2RLghpqsIAhtPrdXgJvujx4DTrQ3NTTRzI/xhsxp2aS5aO9k7kbcSFsyp
6eE0oHTW+X4ZsEpBfbjw4rfkXEhm5cBTMsj3+RSUmoGNRR3OG+SwzDju2twO5Rl0
VWy0YUcFtDABCvrtgjUFWrjrNLdJA+wWGcBrYu6jbG/QeYGtERT7czA9haBuvZiO
sIzMgFLLHmTEBFnkQnWNgKmri0n5O8oP0HeyBuEmwnT5V8T9iUqYVNp+RZIF93wL
J5lB8meylEumRvrFrICDrrt4K1fxLxIKXEQJwXZbXZz4pPq1B5ALbSDxVtevxMdu
DDnK7+NS3fGPueeeRTgM9z5w2tufMevZhizWjZr8msIpK8KLOj30VtpkebTnfIQN
ULgi8Et+m4MQ2wgc3cGg+uBN0cBFMJ3za2ciIErZuf/R4kwHOllH4fEQWvdZOsXo
EEqOF3HKu1DNNCWayTWFxiloCXb/WxE3EAOgtnwLyCfDtnaWdIjQhfnhY65gJXyK
Zht41IzYhiNsPF2BWfL9LylcGDozgbDUy2VJ0WKwizLyHtGkQGo5j2w3kdfLlHxN
xW55Bt1Fn3HjlHa0vx1TFzxoGEFAVBhhZXBffkNAB6rKPE9IHm0SLDbnuCLUfrTV
8qsC9SPKJLCXM927MQTFAPhncwnoUxaongwyI2zjszMdrR/cPcygbKuzdZnNtGZ8
oXtvfKXIeVdXRkSFesAY56zKGYzv3Sb8pLMvdApP/0O2xYAtgA4e9rl39tL6vkZk
e32MYUFNRmmIWT7k0oY46tMcufDViTkfdFxT91Evj0zX/QtwixtV0vhqkEUQbqGY
ILgenouCqAP7GSdaL4p7dr+ggRFRLQ1CHXINNIuA3zFnt9ekhZ+5QJ+C+XJwo3T3
Q8WlVIZy/xlVA8FyGCElShPzfSs26pTfGWkJ3PE7O0Rr/gKpnkjF4JBEknUIBStm
6MPgl97Y4aqEKaXsaUnvs95A3BhunX2jXa57EHKhEj6vUevBfMzb9w68iFSC/vu2
tCDszIv/BBsMozOVfuzUPOsfdZM2HTgmrvaOT93F6vxD80m76evNcWBipxECPxCx
izj2jKfL6rj97lUTajvpnYdNulRm1dfG5ux9V/DQgTxlT3xGECOyMPOZL9RW5zqk
4YxTAFLP8/FByXwCczuNpTB7C3KGRAzzHBzP8He1QXABPiSHcdVWLwq7z9Njq42N
FBuQBvdHgdR/HTNYqjRHCr8pJICJW/LoJGIPKfpb48MdXCbovwfgiWdj+nMQtMGB
fmqz8lFTNV5q2+0NY0F7wTVwall5TLBnn9m/JZaGYP+w6fVuAhZQvIjgDB/2/YuK
vigek7MIRxZujZ7FhX6xuKiJR1rZ/m0dpYqAUTrvOBiUyoiIYBJYg0p5GyCblDxc
ehHPnyaiS3qmZO83Vz3mv2ltWJa6Y392wBvzhMHCPVZx7gHdPI/SJnP4ijjXh+dN
yJswPVflvBPSMnkeT8pKU3z+0i+2YRSnh5wgivJmCKk3pjoD3dmulmYE1CkUY1rH
MAz4CB7BYJfwz1acPq3HcQoFEGBxE2NyC8G4w90jMAapw+/X8Uqs0Cb4SVChgFBf
gtjqerdJUQaXIir0bQbBd80qAaXrPuwKDKLedQUHcL4+r19ro8pcLeenATC0l5Fq
ciKJx9NppWNE+aJu9LBFm1nylo8366SANmMIWnPqd9vw8Hl61Gf35r9CFFt+HcMK
Z4umRN2Qp8NE4co+od9s7WSoKjLrmCT9qgmQCDWW3g0yzfWgLtKpIwrZoJtN4vWk
DFG2+GmLhNd2t18es7GBm9soeE6IrcKm7AHFVXW7Km5zqHnPZD47itqXjrDlw1CD
Vc+sp+pl3I7223YJK3miGQ9H6QJvSTUB6X+sEppGJrHDpKw8PFrsaYKa/AVECOZo
keTL6zgZw3CSGnfFNQ00BiYz0uzuEQlfXJjgFC5uJSyfEwS/TIPBL8xaPbXQ75eN
0m3yer5t6a9S129vNbnqC/+h2NDohHJ/pzKyK+nWwZYOoJLAE9xWjvX/ehyIhaD9
2BnqZnipxIHy99B22Pbajc+c7VFzV7ylFjoGBUl7CDqdFWs/Tdq/p0yZouCcJS1M
aNsgOV/wt/ZKCSNzbjSeZvceF31rnHyFI0bYdzmTDytwrH16ruRBGDv2+z2q1UUQ
Ksf5zGQYfZKHpcn8ktMaokppmVWjIMAKX4fcKHUkMZYn7/Xn1WddOG+Yj0a1llTp
d3Ibb0B4J8D9yAPebyowPtNviOqwyZUivWErtkmPWcECIZ7Pe16Gf3cW/1wcDG6k
UM2YnZLXn+/DqVWyGuBwXNHwzaNXG0qZbY55JEuHwD92olzQrvi6e8Eq1JVQd+au
TBPk0Sx7CkS5bg0BNtAqYm3amGt6+6XrJwadwQCGIeppVMsaGpub5omUvDlgTw3k
U9BIe0BSp3O9eRGiT5ownbHMoipx0m30Extj2qtlcD7h2Kr9EAmymuPS7wVCMj1M
NDfXpBFs7AxNoZFwS1ga7jAruw0W63OdEO8WemyMU8kELGrX/rTVVi+prrmeb70s
A8y1PY80j4dTxyMrhSKtNoz57qHlTkMTjw1a/djUafKjX8Q7+zF2kGdhLwreoIoc
e0db3OHMX/VvwKh2Te621kAiREGVDqSO3ucbEwUW/kuOsyatU8HKmtB+JgIOaL1F
eXWoYxo9mKZQLAK3N6PcWQ38FVE+h2UCJNnOg3CxmNrmwGabYFPqxhM2uwEKgQRX
i68Fo2O7uo0zR15aEYqBT5kO0WT3RHPwPosEjTJzUb1l0KizJ8lJKk6+iOVnPoPX
IjugJ27g2lB4Yiu6ElJFhiFx9gcw2vO3djgHddSV2SK0ucO0Z5YUjOW71/w2TBQk
ZJSJ6bX+WK7ysZZ8u+UWfzQ/h1d3sdKOyD/0iWQQQCZaBLP9bhaFx9fymrL1w7pF
3A94iTJVbi9Cx455kBx8GdmN0ufiHkA5BPKs2z+HLEWTndK+EJrBOrwwT6SXjMJb
yGKhF8Q9ypCTQgcoZOyvABh04ocwI1u28zsj6w/5s7V5T5U7joAhEG7G1ybZ0GGp
/D7ZwCeutpDM5qsxDJ1A+60MwZeHxxAARYWiNGdBIMkF2qg0SB9BLLaCmdc84G4p
M19fWFxbghRTeX12nRyEqVkxShjqpucqI6tEFoS/Beopap7WuvADVH25IP03zu7F
9VGKu7WMvvltD0NiGZoOKBKt9RU1oPnKr2D4hGwSypAMnkRReTo6geQ52c1UhqCn
VgNa/OUxvFin+ggueNF/fVskVVDZ79XwRFxtNHjyZkxMYIQRM7RqDBxjvJKs0RQb
OLa2oirj0D4scaUumALzf3zy1bsb4ck/BCSkg0VK5uL5Q86W7wAS+flBDD7hU9rr
j4rR4MMKaNcUTMhSqbHyaV0Mw/3oXCtPuIZUrjrrtlXa0+2o4h88Wd3jEIapEkRR
hV/xlXH08iJmtLMnt5CD+/z6WzbViYOkzt44jBbKLBW/dyvikSeKGjPxl4AjcARQ
SnOFp9FJ0RNiQAYZ4J9PEZjTZsVti1rMc0DBOyGcrIbnbgIvWoOGp2Kth1hsssfg
+Btfs9E9dF6GUePTiGvZS07zYASIkxm3cOoVKsQZqBwgpDkQg/drrB2Rop4SRt5o
7INFz92/bwayJzFYA5E2orT31OLbShYTuPjGK3L97GG2zRmJVFoc0JPG0Xrn7Q7X
RPBM0QrgvpcZSB6d3rruxzARAnt3Bce8d/HWcM0wlG9ZEQQv+LodYmzOF33AsKeL
buu15cjEbtHDFWsX/AXmMuPZ/o4COoPcczCh2ELtd+uxjfDmfAVQA9YYo7bM4lk6
s5FRPbrMp2msiLr8xigRrg+qMf9stfN4DiLxQEa3fQpEGOy/cDJuOzRTZZJcyVb+
O6FrgVOXZnqJVt3TLDVYWVb8/PTb0+SRw/WCj8dEuo4q3jyifcptnKMfrbZe151f
04rISP35lzOd43KJEMS6Zgw7IBQ1ouhATOSRD9U8UWJwYhb8MLP6pMBqfP2ssb3Y
bZwXU8MredburdaFU6r5S+6jXQZO+4AhGe+eJCUIzYQrCSqKRCXUuxTju34z/GwZ
0pZy2XbH9zYkFjDiHY0AUygIwcKumNgpJEta3jC2huqsTkwJ2Jk+sABNX/SVHC1k
i53/nJlyqOlHsM5HSo14V1iXXq80tpaXnZubavvY0KeRvRnuJ5gQHFFly6Z27Ka4
+Ut497z0tJqy4MrJ3gSziTXIJqWPHmVn+EsaYvjup/vAAMo2IfbDRgaaqzQ/gQxG
NaFDxqs2mIaEplGX0olmnrW3Sua4ATdoi9eFtNs/ZBjHM9MZ/DhZ0A0Bwv5dgmql
hf/Pqy911wlvGbzHy4wGuEDHxOMakG/6JPF3C0Y2TjdT4qlMyOo1DJfjztJOyVCo
LMVBDxvOLXCvK6E51vQftxRf9T/bWpgMJx3dF7Lj+kl0hXLEoKiwLmYu0+k04lHv
N2i8I3uGmbQQqdrHbodx3ypv1R/UZjBv0JSeGCJDK4k6Wj9RW2LN0iM4t4YTCaN2
DYe9raeVGF8w/pn+d7k+ukn0rr7uFQ6kUvLEmjy3+KK6XoLmXRLfSf/+Gna/VUCV
6/sUXLKP7pXTGroXh2fBZcfisrGkPqGVSBIIOQK4nC4nq8WLyeouz1VcrVtjQ/DA
edhWFHGOb8T//zyuxuRMqykqnCP1SLA1L1hMW0Pl7Bc3/iizdH0U8jXQAAocIO9y
ozwEGbRW6ZK+ZIt1XIhv36ZHKX1APA7g25tGelIvqcUqQlbA7mS6I/AvDXpa5W61
UECk0WDN5ZGtZFQoAIu6KFHQPGxPmtmoVW8YerhNX7IzZ6Q2VsDBymkYoIAGOgvG
MoL1iMlnh2DmpA5aASjW9DrytxKJBw9AYSa2ifycpIo+Hcvz8AfCyE0K1wMfqKZl
oawV1FCk2DtGzxUIkTH/vLvuK6PlsTqoNXOyS7sMx5cQN8dK5gMPZNaY1HJTLsYU
0E4U0ojN38ZgGhZ4/KBoyocBQBpFfE2vG/pngQQ0HuZ3oyjxHMTqvjvaTJFPHjl/
jv01bHynQMq/w16dRPsiGb8s5oGbExgspVg0y5GPWnGeiFzKAKXcewONQehd4V/Y
VuhbhUpWqmbUFCVBqvOdrF0dPJuZ3CUozKWdGrBvBDQMZhFG1/Jd8rc1PhdQIVlr
0jBncn810qL2zA2g2bEzhh5gevYlmSUlOmqYiPBkWiKRZNMR3JLdz6ST+OOZ65QR
mce3zBX4Nbwj1rWqjPJGjXMPL0YkATseLFzSIQuhHXfBoA79JC3g1W8EfMFj+qnu
svfY5SXAtG4VJcDYbZ8DIZNOqe9Pv8KxfoLPkO3EA8ldWcUzS9Cy77pwDQgcOQtB
91Js5WzQ9r37dtXstkmGi1QMPJClB6SbhH7TeWqbpF4OfTi4VOBdoqWNyq9zM2lW
iLKAjV594+ABF2nu60KiZAmmOZGBVDnY6vQn9JoQqBsBbufzrsKPTF4OETk0i3cO
TLNG8inA+djcfmAWC/+1eSIHtbNarILSFOZvFYcQi11b9jtjZLtinqv58z/FrMPy
I4L/ZjaFN2+aFcyNIsrPRiGYwLip81I0UfuhEjaLfswY3vC4eID6/LSxOJkzivUB
clZgXBorIBLlB81hTn+UgViR4Ixf15FEyHAjGEsMYzd99d/PJjp/dl0r5RCu4Qwv
iqqdATlnUk79Y+okjaRYy9sM8uayJRKki4dPnzMPkuRDPDjk0d3+E8vhfwH0179C
zdCfyzy0NP2r+0ihnuC4jg9fQwvJuSTuyGqVaSZ2vuUf9U/wBnVGjbdryi9INDj/
HeInvXDLRlk5pFTSfcFHKp4OhVooqoiJWWS3U9dm8vxcPeU3h/Aj/rTC/YuzcyTD
Sv3jfNBYNrnVqg1OroweFtE/VpgR3aLm6B4RvvmPO4YauZaVa5TGu/iW/4LxQBHs
MCDO48/Xu6c5XMMtbUc63kZD8NhZRj9QPvncmcMgVhbFPeEie4VTV8dhTbkyViTE
vUGkQlWu9DnMW6aWkzpjyWMqEm8MMahfLnhYwsXIal6gOWpjq1ftntKnBnxp6aRz
IfpBtlg73mZy5jl2GkNeM5bt98Dph1LTn0aIxCSN4pO33n0R4jHk0Wiukva1JeLN
zz4nmmLOPh3ggOna9yGxPfmiLSKjxOVYUrq0KUL+XyrIQkDF4fCPKXQYIv+bdl6z
Bel7/11A58+5URUo3FQKQAz8hPz1TtsSxqfU1jmDl6QcgAKgPtKIVIhmgXMXFb1A
ck8bFybvL4vMF7CffHTBtq+4H3Q35S/0kFLTV+YHCEvM3jVDOtv9OhnQzz+A0qQ7
CGlPCOJmGnXK+CXbh0WuGIeLHI+6rB12sPBspDFmtO0gQaYyaU7lG6V0XQzuQwQP
tQdb0I0Kr3xJ22WY5k6GzpkgCOJphfpixIjH9oZxycz/gKrtMiIUf18uat2dQxkS
QAUmwW/P+d7OM8EjFU9L3CkoIPVCUAYs9/6vB/QBuk4TaVKy5MmEMA2bdW7jnHQW
jE1+yNMSa81MXZ/YghT8EjeeizO7UFgYbH20zpfzMcqxb19k/O/0jer5+vpDbZi+
Pyha0RwnCdi8T+UwJJHOFShppbI8MaCtzRTJ/UZTD6FwHorfxY9MTFXiDnKbivJn
9rIHHMln2XCNGT/Dkyx+NIi6IIPXlqjPIthYcj8D6c8Ydy8qVV+moPBuypuWf0b0
AOH1fK1QZYfgkUY7cnT8wfMrkRhg3xP10AlqB8ENkXzgznzNeL1WtIXS7sr6Qz2Q
XJAiL4DdhNzqFtqIPnfZVpFrVwcZ+5O2gv9IGEVUDC5rcglmcGfwEPFa06xfOc26
AW9rOL5ZK3zj7xBI297vyvte5eMzuWrCNnEfjaLjDOX/1tK6ezxJoYFq5lyJAU2/
d1ihI2+oSxNLhWDirXNeu/GwYXkJYFEntB8Y1uyUWjxBmrJZBEYcwi0/oCymq6Vv
/JW/9xJpRmTsFBmXeOGAxqmI12/CJvt9lxa4RqBgeP0mP2BQ/Tluicwf5kDVsDrM
Ho7qsz9b+phWPuZ7jUpL3k5v8i5qpGDHIybp5SHoE7qsdGQ966PPahN/xHoCifBS
aOzFuuq2kiOjI5A93Jx6BvqPbBh6iDg/HohMi001OCA81LY3OXnUOxJgkcmlvYzR
K3qD+P9F1UeuOy9AAEi1+isz3OdSN3VTpkoekHWag75G5niojkX7E37baHDgy8qL
jKeWG8FRnLlWHJhUZXcLcKU8Jg3qYgISRIV8Q0lXposqNu906EiYsI1eAHA5lVhv
pMjw/gAoiy5IVPLt+Tkk5q/sMV1DDK6gGZJwzq28VFlJICDLJQwV1NsWbPPz2+iN
NqGlyZRDATVrHYWxbeiPVi5OMrp2rUkRBRGlESjSCznGVZOLIzJ7oPL2ble6DeIs
6sw7j0SNWao5MA0xV0KpVnncVCB/zdPb50hzXRxZNaECfGA1Atr/EWKP3+dRWUiR
nL5PGZjiV8Zs7qufU0GWtpqgCj5rI3/FDwnedKQRb+nPh3ilSZuIu1pr/r7ihivw
x8zcR878LBIrjdeJJ1Lub9zVMKMeQcrjv5TV4RK3Sp8cign5dRyB0YK6XwZodP3P
6riulVeitJk5yTEJIPt6OIDMcq+YDEHmrypLgtLeLMaUJ3x44mM8tr0Qxf2VX49u
FaCkEGw17atLi95rEHpsHlTtNK/zAm7Nh8ODFYhhuG6nQ6bPbM/ymxPH162MMaTU
8m9wXKKXLTZuK/QWqmFo8MJiTP85/KbjNCrPHL9t4AYCAgc9++KDi2vJw6wr5DLl
eeFUvivLzmsTAoGyIUhlqF4tTInxbDwjGirONtNCWo2N3bEWWiYBVMdQl43DNUOg
s8nKAa6VIiUbCkSsGrvnf5kWIO8jYLgQ+rQi02oTn1U4apaZBi4H2j31F5zA4+vB
IGdn+meR2Y2XTyfntDxspkivoHKwsg+RhUIuPouDnO2ZzeNRdr/9p3BZeqNru2hM
5t9zd3JsIHv/AYintY/yp9czJjJjRzW9f25vRJ0UvE5qOnLL/YFUM2A9oaSdReqq
XTGtEbughiI3fcknC67yRC1NQjcXwFxAHOrDsZ3H6n0Iibx8ZkRAE3TcZmUMTSZI
RlmFA9MXVw75o52P4UXrAI75PWK4zRcchaw5aEBCs3d/ba9p8705XdoriLFMSgkh
4Uv1AuD+8LLegFOYDUB7VoLh6mmPVIsmfjCrfqSp5W42n+0fUeItiDNB/qGVmNeA
C03cfLpL018eLqzKMmPmEwCG2Lfpg5+SDoBSogwzv38QNVAdeV4xw+C2BaDALJUa
3Bsv8e/1Tu7/FR3b6/2srG5Qz46VAuPH64UUeSGa1DD+cyselY0owFxhYtMpaKs2
KQpo/HMWkeQHNwPLO4ui9X4vWr0lr/WQGhRVvS+LGNn5C4pqBlcJRyJraE1UfR5W
P2ViRvjuxZhln098EjpsLkPsyUJzOT9GDIvF2C0z5w5qVAre3VK55ZTiFO1Ph6CX
77IJQVx1gVGvFKOL42tlG2E2AGYrNTDg0BqLWdlPO475sYN+dH0aC8PDsLcnSc/E
CV0lM7XFVV5XwGTRYcSI9pGh8qaKwUL7dinvpPkk0nAl/gQVnRK8g91TNhlvG5xs
7u5SoIrMh5szjTh7aSgP19h8Mjnpiik9B74Nd/28+J1zmFhN60ABPBvOtAs9i+sw
MgXl+GbQbC4Gc83bTqfpFaQC6+s/nfViZ8al92Kn0PwwpvsBV7mcxI/OkvKiLpDe
8GxTzZqVowWE08e7F8tJ3CC8GSQKbiFnTmUo8Yiodosy8zD3A+7WDn7ffSFAnCsO
f424+qJnpm8jz3GUp0hWchyg6peNmWE37+SVh3ndC6MmxW+0BH26Go6QA6hNZ7sI
Y7gEHtTKA5Fyd9YcYUsgWsuiTrwO1r9GhL/GKjrXA2exEC45AOyWfDR/9MoUMUi2
zIYSYo2fhSnnGMhdvlRFw2hRBVe+WFHF19a3OG4a8/owsR6Vl5OTDZIZH8nLWN6y
p+xFa1nCHYRquxkSAop7d3Eqe647TPcnGWxp4IcBlFOiCnMWh9LxPsKvVEvUmpF1
cChcPWupUJiT5GXfWEAfoswN7p1cphHPo06H2BFioskKSF2GBJcfSqK9FTvw5CX5
R0twgbSZlDvlwGYMLKH3WgzjNAWKIMAhddYKzJNFL3OMoRJKs+UgD3pUBoILXeie
byF3Ia2tGlmhfJutSlPmtyEbsfWMgtiC6ZDAJdj9NuhXMT1tFkWf9S+LGPO8Uux3
uclSO6iuBsIuwTD/lpJi8ZgK7/AtunedIP4M2U43lhEGGePFN6a7RHcIVvu0lG2D
NRRJDwy1xuoeOi88oBHEFblkXYcv79VK++ppt3z9Wf9x6D+Cevyfs5DTAqc9JSMN
jE3T06KUUzoyqmy40u0IengDQtfaj2wO5kjo2WxZGDi6RXkFuUNNdZr8TwuuK645
WF1SqgV2VLZL3vKIfhY1RdvJQn4DReiAORNWEYc3HRfZ6zK7YOhyg80EenNvHzSa
9JyQG+ntCctgiGzUyYw7l6WQU8ZX4kzEhutbSiKWNjR8DzRCY4LeVg7MwnyWBv2T
8qGys98eVm1lNpVBLMJ/0lKEbzPAVNXw9/TE6Y+4yKP/sOGaN3k3PaIPPnNWHMSD
whg7IJze+8VYpzAQdg7TFU9O7oXXLEZY636NAjdlz6peMeb8+2IrTBpZIz8ApiPe
PSNU+K4dS0tIMYLoF0YvwTaf19+ytTbTYnKbGB+nzM2piV4FpcbnOoJeQuDz2VrY
rCW6LcAkxmJDeRKpc6SpfWEQeNWoKTkHyRo923qFfDI3OfGLpYuxBKo2JwcHCiNo
uvXIEYTtOSh1lmtXgbVQczRE3MAzMu2sYnIDm8i50/Jjlp8Q1Glxn6IcPGrGye8Q
si1Alvadx3od2D1/PCJOvlAfyr8Dx9JF+JUT4QeAeTDg19DWZu5tAgANiX0ZolQU
Rka1B7aE7g0b0PAZ8IsdU1DxFLuVJ6DC1kfTs0vX4eXtJgyU3mUXTtQDEDp2oTvl
YRYZT4hbE6CF9plnfimVisHPTjUrijvptjm/Gb1zOWmako3j/8IbZNTY77vnn90C
NknERHMPdz0xuZXTsYpVN9CvKP8856gKs75LVSQyGs0bkedkw+aPJK8BdddNSHKB
jijWzinV/1oEGcIhkh+lx8H5uvS5KEuYw/KMs4uItOY9bTsxazMCcTLMu0KOxdfz
iZdWrOUHM4WesmWp43V29cKHmiiZqGNs9lHD8KsHeE8WTDx9xMOV9qjSU8Kop/5Q
QUOHpWLasYAyHcSfKVLtTjvpH1K/PaMyF4R90tD6jEtpK87XGdCHU3ZUlMp5yqF1
EEIDZZ9nZkuq5M9ZLS8XClWYSqOd/oF3BwCc2Wlcvd24FQxCvStr3Jkz7iOhM6f6
JO6PtCVOkXHnCgeIRA0AQhf+OCKCOH7rFCIWDEOuBj4aP4JWE6MRw2QjTD+eUxH2
/RCMLM3iHWopFjNwblESEi56ENf4vvcbdAi7elfm5RJ4oGAGFnzDfEUtAjBKz09i
Endh3kcTsT/u4yW8lvScIx7jUqTVM/IkYTO/zyDm5O6R0bDyZWcCs+AciKbQqeB2
NXAPhnbPhjecKz8hMSaPK/2qXtAYjY4bCWdhmo3GtmdR5eF4PjeV7dvEyN/24LY8
ofeSjTEquFyLKyOE0zHH9+ZP7ZUjUoc4Q5qn9d0rGKLcdNRR2JE1634du0MZdY65
mh3yWq+uPNYUgNkg2wKZdO/daWvuekl/4WG/nBdHauPt5oESEUBbOCIdRqbKhfNg
3d6HI8mwtc4hlCKoBwe67KFB1dMqq2/GOG9q7kphoxhCCOtLQpsGBr1isU/BKMFe
exn/2su5JLhqvVlg41WbQTiIqtRP4NgSWo41w1Mb8wqGGKQDMqJUQHnKXgsiLJeU
C3fpB9+q7Rrq+lg3JYI6Zxw9B17IcIbB3x2Vi0VkWnDL5TSIeAEGD1pNyrM+c9dy
UwHX8dO+aX7zKcgNGuL2TVzIXqLQnpFN4eBL+edlSotlzd0PsfnbOsYEnW/hqsV7
EDIHOlOga/f6XjSxr96/C9CkezWC+9wTg3d3X8ezH6XgXbHb38T2jI1blXQTo1V4
HpKcqwjsrGyEZdGkJq7xMq2929EPXpx7Uqtq8dZz2MWsTNKLffY67uZRt/R8byCQ
At4IWPmmq7nwUfdqlNPrC8eglbsEhU8ijsWQkob1LvUs8WAH5kR/VGPkMWHIgCgB
C9ICa205wbq02VP+uFWKhSRyQ+6OGCPTGYgMyHBKyxk88WKNFzU67tJunFEAM4iI
Ox/ZK3Fy7tZeRj7aB3SToViH29LS14WhvaoeKk5gkTvri09KArYLKeN8NQdOqwiK
856epAk0RYukFhVWzJ1iwYRuEqnfhcVjKw/qfyy0MAuvRYU2eP5x4Ao++8I9IXQq
N7zyGla0FhtYfGwKjEEeEVFD3TzwMFoqibdsRBN+/ppGMepTJXyJ/nq5VQIEi9Wz
KBxZtKYyJB0yAfJbXmGIz8/yrjslT9fqQcoNqxIlCtuYw8WBS910MHaovrmFpn7D
iWgMr4yPQH8szUrd3JkLFS6YqQB5KOB7R1dZycYD2xJeZTxtZlS4r+gctMlD0Of9
dkNt+5lg/V/AopuSNn0BvArNXbTX9uTvMYISCIKIqhio5v/cn0600/r70pEZABvy
xK6bzeQDo/VfZBdfNKRGLP+DcVz6AvdNoeVJA4ZdHNupTw98gPAgnp4IFa2hVLEg
Wi76dfibCpumS0PJClXZm8zsT9TmlSH9KpudhCnUi/Plf1qBAhwnAiRugE7P86I2
UMQ4899TxBrEdDgL++2jMjpDgTsVvzcJg24WrKwKRLAiWwXFKk8KQXhs7/x8t9i4
hkLRlFIic8W/RQ3d7ztml+Lg9ckm8418xrXVOw3RW7HPWxophhmxW657nftLQHHT
KN7w+iMxmtpBUfWDi3GxhhuVhmo2EU/bAirawF0vrpDTiYSnCGOo3gG1lH8yjUu5
JQwRakOxDz0JZlceq5uK5NCJ5KSO4sOCpKC8UHCE8VruZ0Z+8cFnJBAbau3t3Kv7
sFHk31ATX9CcdrD6+rQQDNbrrIMNATDkf46p1slc2mcqxsetc7NwvnwZ2UNkNA15
V9xz6nvROCatVsJylbvMM6YL02jJpdv4u8c0ewWlKBxFtEeresznNAmpzJuuChJ6
WNbBlzlx2PTAyzYzSOQZ1JaIexrh2VAzuSAcWIKUQh1mI6NNcJxWVCo1tcGX8QxQ
En0RiU9hcboXQaIjEM6CQZOs65IarHHT/p5fhylb1ZxWjWNhf87BS0iX0CkCZMdT
7ayA1PA3T7Jp5R1TD7mzfYIQTYCRrk5/+X7Y4LoY/1SxOnF/0Fw0uKLrurHMT6+q
suX3m2ZEfYZIIv96zARrf2qu6/wIJZZwACYhpPUajukgVcztmRHjeH9S05A5S1dP
8B244wWUxW4Edf8fM4IYgVaxd/WC+b6fnAMRRRoOi/+LiGlbX7oZjKWhjY8tKPJe
D/4M+GTe1BNnHHk+sO0hj1dtz4PqPM8iCO6/yWXRNLNHxI5t9O2HM93O6f6nPW0f
8lAgi+ssQvE73QBuLS+C+sroMYY7+NbhLdh6i+j+cBapDUU2bTxCdSzu01SueMAP
BxdEc1qDvR0jB9dejziVPw/qr6zS247tm5gaixoWzZnHH4ffiNnmt8fKTeZeu7fR
oo5NgEb4JieHXpz+a57wzChu6onNHDn6iqLNusggfSlaMqjTJdlvUECHxixBxVjA
70ky5G6iiRCPEMdR6YOMwdwsHG3SLlMQs14L0FSGpD8ywMUDe3OtU9fPMyEMdAWU
k58V5XFqvvDVeFSqCMD+x5+MvqmID+W3VyPxwj5IJ2SwoC0NHyhNO/ZsNXKbtYq/
Nwf6r9ZmsXA6FTRd+dnm/qutmTu0EbHmzEgWaJPaaBpQi1p4lBiY3R0oSBt+JSBZ
cdAKO0zxmc1uubV+Cr8B80n0vmSHBlKMW8z3y4kY9DqvGd2PgUrR0ip4DwWlmDsm
Sof7XJ/0cgCcVTLkkuwEaOG2znoH2lx8i4xsaQrxQFspT7uhoZGC18ZVPPZVkZDN
x7+egLBUsFYb8vXmihtU77QFZyKE31AjQOAtkUn9BYvK37HbN2AZbOm3ND7GdyLK
noozvKfQH9YQdO0tSuUKCyWDS1THcLeHqSLnP3AjNyA9gCvOLiVJEXXa49YVjse+
OmhCh3hyoWJO2hwlbQtuTYwLK/6bHuno6IRK0ONC9Iwp69BzGYbkCwWXgDZ+/Wb6
SlxmyWBtDy7mTtYOrK7ARna/DbkxYLF0tHeg4y7fLP7Vrs+XTK6O4RIQ8DC2AvcZ
tCB9b7x3kAc12/aDFZg8kqPipQmohYiO+zNhD6B5LKzMDZMAA2jN74z7IuWGH/3A
U4ZbDpzgVvgsSyg1KZex593Ds7qPtQX4MWdPlNAudZh/sTfnR44sgLS969uj7QbA
5mYFLDtbvArt7q9VOJzOBdla2X3hyBNEhnAxnT9QsbEiRPfRUjqT3Fa3922b3z6R
/WtjyrGMLPo/ltokol4MKIsCbbmIZXw63na6+WXqRY47xPJLT/ke/cA2821gd/X+
O79kinzk85tLn/eRtN78uZO5uzJMFXHBDWvAJvVHDWY8opMiXcjfWL+L01uOBtUu
K8QnELYguC5EmmUkvUwZwjks0DFggSJDs6Or97WiAPTSUWDYvMRDHiiz3T0ygsdi
qmTtytXaLYPsLB1DuAUwDpwFEH36agmP8KvU4H90/DkS4rog+P/8nkuXW0bm9nL5
TCA5EM36NJm0DbZC5ZL2qefi57VGsTR5H1Y+RiRnMJHftrk0gBfDIT6SARhEEdcn
t7G+0CzhQsF749wJCnEvJlqQYosK9OlxJEfbSFGHgIwkNpCHmAsxuXTxp4toqggw
YrMpdRpKrUS6xWXg4BHoWYdX0AEfjtQduMZaPo8+KF/HECXG38UEgk2wahnJjnwP
E/Op7sl5K1UhumV1ZLMsPbVxOJ1r1/6Eo5c+RnxMuZ0eF+p/NAWsZluiujkzhqtM
7thm753CLkM6JEqneobUoiidinTRBXnK2lG4J3ufLtB1MdXcGwKrlAHAd1HArMIy
aQbR+lbQ9VfsJE/7Lq9Ok9HgIjKtWTDDJduYMiD7+0NhW6ZVt5auxpbbMbPmbJpg
/QuTElzme7dv7dfaW0QTe3vgOm4WVewwJ8rBA35elEbgBB8GI6msZk9BEjwYI5Qf
jUB0RIwnxKZU7LI2vME2e+U00BPDU4rKrs5EQjWOBJ0+Tm/1xZPkd5CbAgffXIdK
7aVcTGmWRBajtncicqDeNdwDgNYyzb38FF0CJt41rTJWLSl3w9bMDCHfEFgq3oA3
LSj2atzMtIIGOxj0bk+zUslxegl/kVzma8+Z7gCTguS/wNLCCGeEn9QiPu8EnUjt
aNq8mDy1Mj9hAlLy5PjKmj2epYiebREYR2w/HfUWq+Jq1zK2RFjOPT2qQx27VDsl
A9tPhFs3WjalbQHI9sz3svzsP+yNlzKGua4lr6Yhmkx72UVEmWd4YGmYiFixe8YJ
kcJQfEbY8OPtFdLyQwO+q8PUA74sUjjicJx8mV19m1k1s8yP8+ndQdvXt+wqNODB
VQsDW8MximoXMxvK0yuu4ybg4DVjmEFXPNHXpOUX0ypSkCpwYOPeqcwgEoXcyGfk
l5qBbA+Ki8GYpGPx8Wjr/K7jrNz8IMWQh0SiOVHNjO9C59YsZa0hKkrSXL5lndzt
ljb6XrqGzz9zM4faTkB7j0Op2LcSJasqk7+d8O4jmKak90/zvAX8C8ykCC5lBwsj
Gt9ial/ajEKm2s2GRDDMe7c92Xa/KmPRpG4EJ13S6dkBksNajg9kOvrGlFqDlulJ
9Z6kiurF6bm+MzvxaNN3NhV5LxfGugYDDJjjdEi4PIX/2SNyWxot7u+CPPTtO0qZ
Owqm/Zg1O++sS0/Q4081wSh15+aEDeFrx8185o9h3lvyGLI2U45pN8oSlen4qz7T
lX8NMUQSABkfpreX+OSlR1XNjWg28le0um2I4LQe+hJ4Gx9dW8smUiO7fwd6MmQ8
rO3D04RbTildGumhoKE5LXBLoOx1ydHWWV7Q9l+5gdwaifwxxcWHhFDKdNhWwUYd
s2059HykF7TRRogGDYgFKLMTdXPTh4ruSZYtB6enWs08ZxDQyiBsqU5vX4oKJHkC
IVSG/YLaYEP7KTG5uEWiq62IKRckCznD7X89qSE60dzhp+nO0tViuegfP8pJ1mqN
iLG1RHXf61oz9XCT5VN9O3kxl8LcxqMQngOg/1/VnQDp/R44IucHBfSj/rEwifzT
TAQRn7Oj0YTmXMgHuCSIBGWS3DJDSemQJDDqSzHJqWDDKLrL23xR5/xNasrSaISK
v7f3W42lQ6Z+PG6LZpjdebprkltrW8N/BYldjJxTNLCHlURGvORCgcYkk7qYrIra
iHFxOPUgokvtAIh0o3wOfmXt9MB1eo8Um1iCG5P3J7C3Q7ojanwb7UYMupW3h8Tu
lqNBZn7F/t7CGn7BaSDk72dIeBlmauWVm6IYaa0SAKsRS44dY8XwQSep0wY5PqKD
YtT7xvEgALYHMXmtIkVRA68EN97Gr7ybehEFp0mPmgLHfzK/+N5ZCqnH1DEvZSIE
71lmNynDBJgPTnf5PE9in6B1uSZXK2fdlsNXPHLS9HDTQUfs7eX2iwnYNcUPb9Di
0Uoyd44XTvjWI3XjJJ11mciZSLcwkPz1kkn1VFgP0Kpfq+xm0ND/G+tjLK8ndkPL
vIs2SBGjGDKqqyggTxNLr12V4aA1CReNbpTWSjJKXee61jyoU9ysJTXUgtdx8/W4
wY7idG7wOIcxchLT7RZsy9HTje0HFI2w5993SB+vcApWd+mMKEge+g+AY0FD4moW
rVTAxZ284mKJTSF/QZEQFas3Th6AcCbFvQ7asCkSgpfPcZ5CDLtykwP9ndzrMQLf
EUtNeXP7LnRdCukRRFQtot6esZNHalH4KmPD0Oav6hwRXVGqJTWTfDU6jQvVb6Ll
nI8toRSGfr32zZUmQtmd6N/ugTp2M4dgepUqZqKoC4ssMROZ4ttg5k0F5MAIai8U
kAv/qYXLt9EYVqp7AhWF7KGxp6J4k66Hli+ktN+VWF3efL7vzZB07NDLwGQLAh44
v9HCs2qmC09Il/gACxEex30pR+/m8P9u1+UIypmxaFHEMItqDBXC6wKeXaIzbb36
eC0OeTOcpqdhp0W/h+3AA0FM2LSNu6mhgnFGtcE+RB5XlC8X91GvybX6OEIHCkwK
/iUo2VbKty7JrcshNz0XgEth9hpk910ZdEspmbZQLALxPwungIVzrqIuDJ6T3hwz
s47/DYQTgbRTBQOJy6YfJevHXs3KOUBS15Q7WtZsli7mK8ut28mvBuueWVbE13ZZ
VghN6cqR0izvgju/+GvZ8GxaI4J9/+0sdhhJSq8K2g3dVU6xzln3WxUXV+W07bQj
8QW5YWENQj7yg7Xx3sXf+PsyMcz9spsd95JdDnJgZEEvp3ALWimouZnB7AL8GNJE
wGLyBUJqL+jEhW+xBW5L27+yWeqUgqV1/pyEVrNe4LT7w1bDCFcmrk3U6PqC1ChC
8axRNJPp42uemWxJJP+JG9H1/J5xZ8uBM6Nx8u8sILaecIhpoXYQGfvUVggqNXqM
6LnFre0lVKOVKrFT+MITmGZOk5sv2kNUW4t/z4dLrLzl38spQThcEynnOZONAArC
CSPvDQcRJvFr//j9y46ivlJZHsI/ywUf37dF+emVMvxjjS2v78F89rt06/6xDgUZ
YBtYOwlvoym4rP8yGAuXbk/ur358v9YKmALl33RIzGDp2mAD6CnnLLdg90SKJdQS
vRhsfvYIt9VbDpV6Jdg+4VR3giKUKAnfBgRf5YxPIszfDbKy4j7pqlXLrj/xWzvJ
DnldQBZlgOtq7jaIbbTQsIZzDQZZHyOo9waVJ4jTo1db2hQUCEDpFaHkQ8QM650o
uzJwDO2EI7rIQ2hFdgefN8k+lBoQldUVkfG+Dyu09rMRgSceXcF88DiBz0uzIOzB
AQFIvJ+wt8W/Br+mLFINHrtIWpV22D8IPZdNqHX2FvNUrCkOVYFJPmkVOHWVlE0F
UmfjqgAvue8qU6EfMTzzuHTlResVhX5W5DEQEPj8wukEYfcU4a8Q9uwkfg1dae6d
XzQINrAen1vYcBVgjmcCd6AM2YJA7zEyteNswVwaqLnQhEk/8H5pg6p5MEpSzaoq
MR8TY2lqZJ1UJMgO3aM1uCtJOb9Zkk64rl76xxwkDG87+jT8SvBKTtS+RIHedphb
kKUMo7vGZ8JqI/P39hzTngz2KnzSj/v90yLohBFZGEj5AbJg4X8wqwJbSyq3YYSb
BXK62GJ6L7mOEt+rptlEvCstT8vMmd1ub5Frr0f4SHcTTv01yEG5aP2jV5rXBIqx
3AUVIzJFYln6DkcNS3Sfc0UzCPaLIkKI3LxTMHNvuKC3bamCEpW9FvxTyq7iMW/B
/PEPhNvI1KSIQPiG93x8zc/loU7fog/QFdQ0aCEUdMS7y/UGA7urQ0lxlpIx+/0i
Jn11433ZrdSTwx5Eqr5Z4DmfoMkjgSCIfPoT1BWsCws9L+MYa+MuxCDRusBJ4OyJ
rMUM8zzGMlK+b0pQrpTMHo36vKsnvrE9eOYiNZeYWvSJePdcprariMgwSCrZsdhg
dh3mxo+jXVGrZGORi0lLKdp9diMh0VQ9XCpc4ngshl1RafqNIGur94UxH+uJEUT1
6L44OZZWdrAIvoSOtVVa/wPlTkARf6u3Fmb3gvT9wJ/EoOI93Iqg3RWnNCeEa1xb
rFo3lx1osS0vvKM0vye86GiBZn+m2Pr57FPYQcyjI/ohtLX24UChIkXa8BSIjEz8
Zy2Cp+jN52VXHhbC7iqt6PexaJazuCzKSm5mB8DDv/nylagSx8rLesrgk4jpBBYO
Rk8vbmMeGURR+pUNrKQZvY1RaSTWa+Z/ZimgfmvErILi2tbw1GuhcQ9RfcxSPfo5
rcJi7MOU92tz7mQTAx8iBSrq8s/0x4xEh14jC93zb9aUM3lgcd6gQBqs5XggVGQU
8RwiGf2r03vdfNsB5eylUrkWD2fl1j33zvzKZLrKSFhcdjYfNtGRsuG87wBx7eNW
dWdUtybrVQ/RImFpciI+4GW9BHkSEkjL4JtWbpg079lR6PjFwiis5P2EYseIAQiv
m31pYkO9DwscqI8LrW+vhEc9CuJOieT9Xd82n2mcYWc7z/1nAFPUKQ9Zw609kIQV
cO5DvvadpqWy8W4miTMcEzTDNm0VN29elOetMmNoK7BkqLTjvk+sv9/ZHgvAT0GY
u1InTmdDvXB97plWFckGggdkW24OWO0LRqUyj6MsugljYdP4HXRSIYwcCnZkfchP
Zr+S103JUqANeHSz5WtYlD0jjEdTGN/LNJZHBLWLEruH+OfDN08mzb7kVn6b9Pn3
HRUCh4hgJs+oY2kzuAWArAzLfjzkEd1NtWs2+1IYymQgF7iRCx2QJ/92dWXL0UFG
LHBWctJXl8wHW1MaZcIOwwcchbm6y2CvbUdhP1lMNUWcO7PvmX9cAXWZr8csyVwT
vl9kYvFbWQmzDywXBJ8SFvDLkn5JOxdYuQl00gcJcIfn1M4C4ZMqgpR1lux49dJ+
h1AL5O3KjAvpcijKPd+NsfkVCAfkQXecYP/k+6ovELpIGvhrXjtrdE/uTmAdwI/F
QqACiVN88rqYtK3b9ZhPGcQ8nhJarkfvjnrWxW+NWpWDzhZ6nVS10rJzA4jmopIw
oAD/W8SWnx0kLVqhAmay8GlZSP6TdhSuvdkFus5I7YpPbDJzOKCFYWMEGnPtiHdS
b6VXliLWwcGmHFUaffmGG7XDuQRv+DkskB+0tzZ+Lhciv2HfFPSEwW9M9unA0UKd
bT20vQKBIG0QPel1lL2fYD9XE2uUo9gdYYxbQZ3ZdpQRtSwy2dP25/61RahciTo3
zs4ZT4pI4nsFdaiTwidH/IhO3f/IEcDVjXrRWFKK63EPXLw2zSSOj4rrjTTMTagg
kIhdCSECHf9I4oDvA/WKAjDFXILK1r72OUeeAzmKvxpe6hBXf79dHf2yM3HAR+tx
NDctbYhffKqUWouSPq5Lfdf6unAN/1EHm7q/8kLlMxJn9a6wdcWACtkqCDKxBwS7
Gq+s7KMJ8OAoW77MAoU0gfbMgiWjIyhSKfdrVsTEHyyhPLpZy4VBxatEBB1h0wJH
F8FocJyjQ0x8ZdkfHTiVutcWgjb9LO7ZJ0oq+k0G0yaBKLdlUX+qsLjp1hslCJ4E
np83VarEWZqJlbE/8nnKsg7PFPHF9AIL0ussz9wtcXV06QBEqkTJKr6t4MWzs5x3
+4K3NzG88KY2TpreSTqf/xHXLVkMPKwYXFCAGS7yI6lG1gKrUm3CY99UOiq9Pv4T
LOBgU2kDFLWRhz9pgNUM1jG9DSU5pN0Ce/SrAXvmFoVS8X1TEhopa+drQ1qeWMbI
PIePJoEwbmvB+KIlCYgO00bJ2SYq1QuM99E+Es+2LhvJKbBZYua/7voUGMNiSSCa
9O02/PoAiDK51+LJSDG4Lqn8j/k7eCWC5PkX+UTIsfFwjTKuu8tc/Eu3Toyv7XDx
216+A7E+9A5Lo3XozoJbdO1qiwwZ34p10cz3aejjC/9VnDb1McWthFCpvWT1ie5r
98J57kHdGFU5DGWnVpuLpAZEoRqKu7NQp4IPQKkBXyh+FSa5+XSev2IeLJupWc5C
AsiXNeEDEWdLNMFb9ohQcIJss+GxFT/0lK9MX1b2BbDGjTQ0n/pTPMSBwp4d+XwO
JtMF5WcbCMrYpiz0Lo1CJVBDJmo0hfy6bY7e42ptLbvXYlvdP7/hixWTAcMRs3dQ
UUTZvWanjoHoATHWsNDhen3c47Ky/A0XpKOqMiiTQI4+p4UdLnlWhJEDB3TezAal
fwkXHONYteO5U43qx1BN5uCQsjMppNJjo5SN2F0Jr3CrsNscy9A6cP3ycHN2a4WU
25/nCzrdy26qT5inEorT+IvvQfDjhCHHFhtzJ6V2vBHIDfWF4ApjyXXUaY4jbPN7
jPJIe60LhOwQmry+6K4QSgjPQEmnyw4P181yaMZ+SQsBE2OiBj6WekiT1FkTV5mV
g61g7xWzJ2imEPm8WKYInyDMOQpkCxT/OYVXY87yNkZLmqi2U5zLNJ4fVm2MsDBS
NrJpJyTf+ktSywBRnlnJI82HpQ5jJBbpaKpwZyAvCTktuqPYGsONV+BAqZwtrqYQ
7oz5XjPINRcRqDwDkLqCAPf+MMvbuXc7nz3+4K0J5k7H1oAGZPJWdbcBk8PIqrIK
W8JpETvZMykg3E9r3ZwnhlQdZZjbr35Y9xK8HW/419Q1hZySOup1UdSra105kjpH
WfT49fFK+VNczgQwGBc1oYHUnHhh9H9dUx1ENGfnZoI/CaaxYtsdXLDElJJ3l5rL
tarvfgz6PhLXAK1SKpNeBotD9pg632TZzBSBTKZTn2qpGfK7nr9dASAgVz5gDjnR
PftjF/e696l2wNl1FuUzcySLCyP7TNWFFPs8MzR22hnHikN5rXK3VMvcLxyAQTjt
ogCW5upC1+dX+uP+W6JWmaLE3XAs/mQByBOp4kR5g4GLwq8EaSVT/S6JNiVsN2C+
83FtXlu17DfHg4fGpClntWcZT8fk0SytK3omE5HF5WHbyhKWD7IB6cWY5squgz+c
/JBdBTws2gmyrFw+725yQOxeh8mvrpYwxL/2t103UhFwDR/IYN1I2V60c7nSYc/w
WoGM5VprSUMVxM7vmfT3V14/fcJ4QhQ2hiioJMgmmvyntXXrJ1VDbUbKZkD6je7u
XtvHZj+QD+oFEcRWcFZzc2tDNKFyoTXjn5umR6ino6F9qtJU1uhc4Vs7+bxysd2G
EnPIrgkR9FLRX89snKrbUBCN2+N0NJOjgMJ63rNGSjx94hRuXHCO+1fPEfIyrIJM
ny6DWfAJcZmMovRykRwd3jEZ1nB6d6v7e/LvE4z8gD1FbXY61H3MY+lc5viB3lg6
CvH450zYYqXc0k+lcdtrlFXn98IbFJ5BPth0aIN7MbIYmL2Z37SkjJB/VmTTXZTM
2ujaEBfKRI0bKvZj0x9kcieLiDVHenPBES+ITa7csMRe6snMXTyiyY5Lc0W4y9VO
ff340srAXd8Wi8IWockXKsDgGh4cJfvFRGG2UdSb9JcJYlei+fYWJGLAdXs8hwRj
HFKd/61OGX6f8/fQc0dga5BcJod5RZwiupETaHBsDEeMxOo61XiyeeaxXlAScIdh
V080xoiKoIFFrZO4QfFDPV/8F1knp8vxkp4V43LA2H1a+3AeIC9tBZRwOKGIZq+g
jc1Kroi8+oIV2VuRDewHw21Y4Vdp/xQNBuwntXs6xgT1bWz4npMQ2rJOWk7qY9dy
81dW1qXZP34f5Wjs8vPZaXvXCGvkxmAcXb678ShimtPhp6MonizBfQk7g5pmgvr6
B1P1QOuMZArMTPRuRa+e4kPGtutkTPDAO7JuhQxEwo3wSJeQwIq+lW4oMKw4Vxxm
c1p1rNYsgEIphV4GtqAthv6PWSmabeIVbJHDTmDKgkQNex1w0pEpHfC4pD55eP9n
eop99IJg+fzYrThyGYosuL1HscD0yZXYvXMGPWOBRwuLbWCAJ7dh7gQDs90ddxOQ
TMwhwwT0w4EjusuJL3BMz0GYQHqJp9k6kG/ZTM+ccakQOV17W1lxft2fVO+hIR6C
c9krtr64lOiGfvNg6Ny2xf8/dMygn8FEVQU+kQjIo1oI4vqATJnsNimwDXUEd1rv
t72BfW3ijPT0wq/zZDr9ZNfy5bsYWPH+zKnoVNKhb9hUWmE5D9ZTjSA8hsDRkRaW
qiFHPQkyRyI8HWyzKEKEAq6BeNrXDlyaS/zdZdmS9Abyfv1YmpHudpH4w6rUEgK9
Z6Y1xmb1EtsSpFUCuOfMnhQb2kHZwx05789NwqMvLaZZbpUlln/iijt6NiVQ/SEm
qUBpk+r+Mmf2fkH5QoRfalmvQG+1yHLGiWT5qHLjb+A9JtFhnySz8/8/gw5I9FOk
mpKaJSN3EUQXyleQqytM9j0PubqVpDhLbPiZ/r6sd5H5ju9PbqrWf3jfXbZ40wWL
ECycnMgLn9ozNiiY3LJaN9TEFWWE3nhfHIGLpN0c4gnDQVgz4IXYQJ35RRPCO9NH
eBLQ7OIMOdTig0W8hbVaOR5epv1xnnfe4D2N8QbGthU8+xVAJPGmJzjTjq8CWuNu
lHc3gsR796hgjeDfgXUc/4lpE87pQ5KAwWsbFwFRXPRhXFHRjijW2hcOzh62QyNL
2BsOBjkxE3WxInMwkZ7LAagL2eKpT3ozdGIETU7IfVEwXrhJ2rqWanu3kY7wiyDj
aVkqpy6QsMUkD7ikMACulZWQuGyPU21aX27pqlyQ6U8uUHBRY5aiekV/yN7TWi+x
lj4YDuEGWe5fb74DZO6C+EFSUoI5eD2QjnDh5LCjSMbPiWIQkJgKv2BFttwmlBts
p0fSAgOMWOZAvZVE/mgFfEVova/E6pePea868kzKuLsOx57JYFcitBfHeiCxHX/x
yOGtwP6Ge8RawtI3JeCvZdqF6/BUw2YVVzn5fWamri2YTAK6ESdRpIAlQ5SdiMtS
ps+w1rAD0ahmuMo7LSrX1a+JwzIZ/U1/Vb8e3vaDgxOXqCviKYyr0XEvcT/7Jb/2
5oYWLfAki39M0RiDx8UILJ7NQ3KtnSnEjbHsaB4zfI2u/wjtVq3baz1tzRzpUetz
SCykCtjaySuLked2h0EuV9lWUyiwo1oGcQnS42o18+orpALc/s7lNWG52JCtg9M/
aLdihPsg5kWmwbfPfP27rCgqxObxZFXwOaeSBLbI+0uR5JVvGCy75ZVFyOfefl3V
FgjaeuKcGBSs9BG2yJs8/J/JVM/V8QFrTl3E6Vhs5fIZNZ7qiI1YCAnmpezaxEE0
+y0Xf5QR4WlcWnO5x39VkkNHPS5RK+72GmUx2HoyQ25AmWMjcbyLQPLV9Rjbah8H
weTSiBlfdQcoHkOB1clAQh6DEvaWeKtQng5Ggko6sp9NAlJIDTrEv4mQvaJGim/d
LYr63G4eO2AWU0Ea06gDUv/rwnko2zY5j+cik0Iwt4E5glyCnm/n42drm8fhcF0v
ateq6D0ZgfpdvthIY+0vvlVFN7+6nCuSZJ16/wPVHDGeRV+uzsuwTv7Pm9WYuYGp
F9sXEUVRngdBadprs/xD436HW67F3So5nWI9XFSdAE/jPQHuvww7oMQUCmFWwQ3/
iZGzkjvc3vb8onKw6RHjPAUC1zIu51gZOK5mJZe/EU9nFUbt+nTN9mFOOFIwvepi
INcHdVYNoiFYGUGoIuRmjTwa6FxZgBJ/TGLXNsZY14Cg4PoEPTD5gDA/ybNrJctn
o/CRbdAGHRvGMPIuAhyfM6HAV1476kB52FeGhn2C+MH0bmWTgq1HjL+VcYpqY35B
u7UV51S1HqiTCY5rMzQldLJc7bd9ldiiwzSqDq+WeKrvqGm6MvzInJ2nkI3tylxw
6NSlNmG97h/ojaQ8vIDthBbXQUnfqrU+nfDrhiSnY+MaCpHCjaL0PDyxLxxkTCyg
MZTCe1qEn66dCsSjZkqd3HVjrUaINDKkeLqKy8AU1PW8pL/c9EeeBdCIXcPZsmVy
IHwnadF3Azb/J2ak5q1wU95ixFx5G4Fe8tXoCdN5lk0IaJsBV/4jzjbewOFEiltS
oMOMIuSQhC51KkkXReL/zGTlkx2CbXEJhCdgRWqoHwVWXOToPXC4xrBaB5y0gkXE
RGAtyCVvey9Ye0M8+YStO7NKkq+x3K3kRDuQwCYc0paMn5Y7osRx98rJ+0K9BN8o
A000S3epPz4Cdut9WxqRIBb5JvYW/L2o/fFc2VY0juzxyvtEhNUukAgdPqoxMj9P
a1iy1RT4bnEopwoSc6cuYtvdBoQHDwwxbGO9RtKjC/dfkYRF8cfVyzueptd9Pd2/
cLKjUWajPE8FKOnDmQczGoN9oonTRhnLc/0ULrg1xpvTTVSTFRLqrlFFqHhlq/4f
Xo2UoFPaEHHudullvn6KftM+cLO/LrH9ERXz6PQz0ev3+J2FE1TBNHs6m+JG1TkP
Mh9Thwut73ARQlF3D6FB2aAFisnOAMJZX+wkCgUhMUILyRud8b+KZaWB5lKB9ceK
mRvu6DwNOU4yD4cdtH+r56fympqCG5r8IL7+gJTqbgwL5hMXo49bU3VNMvUZopfW
fitEfmdUJ7kKys68VFx/hXAgcSYmFhKxi6VhS3n0+2YC3BbkozmvHcVPLpPzAH+b
KjQeqUlVh3X7QO1SNsjFvH1MOfxcY8HvwSCmAymRrjGtkHSBJ0SX0i1oqk7NJ9vp
PcppF71fDsIRRKedf2lpoMfDk95GttRK1efPTEpbBJZUxQigTyKyY3sX9iZTx9II
H3AYIYyBSPWtYWuKIHMJCrsyCA/LcdzpTcj4zlLryGX+I9DsWpCORX6LT96JxBeh
ufKi7yofPXx+E4MUAdoBX1pRbjrJaArBeWUd96GHD582bztJGRYXMeugpDDNr7CW
opDbnAQWGzqUCQP7JZhmBwip5BBQq5MBq2QphObfsbTPzOWI3CMmxAvz+yQFDWmm
ai3j6EM+3QdMxQCxjSf/aRcUxn5yYOxh2g6aeJlNKOOg2gybsAL3+Vge7U3oAXil
MP547RArKEs1CZENFnpptxqXTNCJnLTJU468PwQ2QtEYQIHi19iy3lXCf0R1v3Om
qXnEAOP8X2KyFFUdyGNxQIkzbbtq3Genu7NIeI1nFRhcW6sFvct4NEA+jgCKUNM+
KNaIrs4407lx8KJeGkTLQ2LmnF8cu9tcFPtWsYbWGtMInufVh6NrQecuKsY6yvGr
6kgyQnQvUSDMJ4aeorq9gPaVdN5g7r5FwGtY6Jp1/S3TIPVWulFeecyiyN13Z8o9
iRV33BLDWrPKpuHiqiozblUic2uV19gzVV5Fo5Ja07HFmhV8naLitk0PcK9MdOro
duNwWv5ZtjQ5KaWxcpkheyq7T3uswGrXdleO6jVyXJqUMcwgWUfxpgQynM60laMe
N7v4pXqjtH5WXGPE3chEyneiGxuB9wrkykBJRtRnPnYo3dmyw9x92GykLxellLZ0
7mKW2Qme043rDZh0irDqrNgw+1p2rGb/k3nasgQfW0sOfG0XWl5314Nkn05M5HxE
y++u5IhdzdVter2sOPgpv7VVt2QPsuwyLo/EjjpSLHhB5kGPo673k89dagWt+E6L
hEfcbtYtQQvR0ZlQ6zSVXeedYYVw1N9YlQDNZ+ClVjGw3GlMOyNjQyHmyrP40mIq
xPMfu+864Y0nqt22X0ZZWtkdHRQ8+Hm7vtS/SkFdGrG+wiy4SgEeUBWjebYopjNJ
MEw5qVujjPkv5iFMsUsuXQoaiMxihdE5lzoUJOFG+UlCkpviA+6w+CgisxrEJTu8
73Wh99v6Qm60gku/qYX/nzKIGRQrsORvIFoA9jdKEWDNiwZk4Ha8s+wgrx1lcWp+
6xaR6ft152DqaZZNJYC0ixJN4IvkdXEkHV9IvQUK8QA9iu5ms3R+Q1SBgY7zjTFn
B9c0GqPi59CRgo1S6Vs2d8Q+PR5zOU1996Z0FWfyDJRTkUDNqhmpGTasFWuWycvB
AS7qXk36y5an6q3eHzhAdts1TUI6bepyQgZiSUuJaSL2gK/rMwf/aTNhwh+RYuWv
h12a/23KxP2uqdJpg3N6V3m+NZ7x6ItkAvmPTdfsB+rzMNrbuX6HebwhT2auchgt
8s/658s8zAu4EScUU1tQ5sMcWY7x3YX+hXlkXRahOxr0i+WSOMB14uyQZPYn+0oM
S297L5FOoqawTH9/mwKG2Ihu1lM9hopFk9EmH9xc2QQhmLYglhz2ZZxmz+/WsonA
MwcPSlV00U7JSqNrjX5fEHpxjb56spQ62ymHyZMkHxf3hc2biIiYaXhgQSr/f0B2
QgE1dw9EilqIBemfvGxIe7aS3i8K8BxEsClNrrprE2KdAud6xByLfQm+78AswJX0
mBqt4MIgSrsV8f5jjYqR1Uxz393D10Z7D/Es8Kvdb4VzyVVrIEsz14Z49nqe6kcL
lpi8yQLUQnn0tQHbs3I+4tie4NKBR3EbiLAGB3AdsZNkV/s4tVDGdeWlrYf0AbIQ
sZ6u+fp4M5CFhmMhX61tSxX76SCx37iD+RmsiS60i6eDN1eCv+UoD+92x3oDWCQ8
fXftCU+YrNDbAaTftR0y3Nhd3YZFF9mRxpJT1sn3epsI7q781ikRSanynjn29xwp
F8QVkPj2PJooV2L5pkKHIWMtxAMALC4e1aZPRl6HMTYfmnlGtoWBYOIrmZt/5a03
KlRgPN3fQXU3i45lisUUyYJK2oAZNxbBB3FwT7Iz3EJmC5UVQzrsunWk+3PLz2mb
kpTEQDmyYSuWZl0nuFcWmZjce1jv7Rkzl+cDZw5WWby7ZpSvkw78LUXmsGDHCl08
zqn+UE/Y5WZAhxyJw1vsqw1lQXl5ga8y1gaINL+zedSzn7Mo5v7YhXPWydrlQMQb
06soDU9SJMHe14nkQexHTKQhpt+QDX+KFBm356HSjXepw+r9K6EgfR47+7xjk87b
UbXDGMTM2azxn3Q0RDIc1Gv4zc9mI91kfdq9FV1U+z3WwtF8SFjueqPThZfKYgwZ
LbFW3wTWKxQ+G1O1sDa0rlFw3kU5ye4xGHg0iG5yrNzT6Zs9sYLJNlo3nWMwee/Q
JzNAyMqgiwxURb0WaeSS1mDpccAnjM6r7ZbKBfZ4+Ikp+gIFz3mVqULVm1zkxV9n
8AyIAracrruO9awUB2rm2LULBlBsMaqd5KGs/mFWfu/PViWPSB0RkHesL0xdLhqD
1hNAu+hJ1ysvdjrro0Ct2HMUjRnP27+ePYIa7HJ8RDi+5n+YTsBYjrViyFFN8RJy
3ah3t7xw9AvXd178VWWcKsioeCGsMBY+JorkPRgKNuz3fUAb8rtKDWf01vysrbCh
kJxG4CxYP1rvnhDiiEdWs2RG6QnIbilXZkHnNUsJZzJPBCmxAUV/PPGjzT79jzzC
TIajG+MS7Zfal3KOjLkcZGAVSbMwcVqlut+AUCwioQDDJ6rCi8GrsBxPV4hOr6i/
lvGutceIARMi7MMLDuBjam+HL5FI7Oq+ZNrJp677tu0SVNrualTHB6dnofYOJUGD
oMKJaTDUC5JzBX3u+typRQcI9v8bQ2eLs7C/9RlQVsTFQUITnVPNlhUcU7/0TxuS
mOEtDBhmbaQG09xTfJrNwQjxkOU4IllAnRcbJsEVaT9SSO88tZHV9n72Nui2J5cS
gKgyc+GkX31CgzyTzdSeJ2yyJEyl9L6JsB57tdRWY6wQqB+MNXk5GmmMVIO3Lvkc
vfhkAcd4/UFCRvaO2DasRK66EF9lrhVXavo9M2lvOJltldgKf+LlRUd/8CyaGJj/
xX6TGkc9uo0/S1yGfM1OQ1Zidp6Lo/p0smbmEuk2kvuB5Ipkm7ZVsRyaWdeynNKT
GmjqAWB8a9O1QJpi6mE8mtzjtiY5ySo3c6z8/BkuG7li3FjwW5jOjj/BpcWWdQE/
pEEO+2/NpnK53c73p+yjf5Bt1HcF6Ao2hFRk5wvj97d8+dvnh/GFUx0+KBco1Oo+
AFfUnlMnmDIKgr9XfIA5t2qdWyHUIl558NdCDrpyJmzPU2GFkXQuxh++S8cQAR20
7y2Rkkx3M3IKjSRn+qbgSX7XJXgza6iWSPeOCgJIbJ72rMLk8zs3KoN81fYp7+zB
EJdijYgri7sgi9Gq3TkiUQVjK9oEDZflW00qcSShLUQyBQK7ssEhRFathM8GYDCM
5ANV7Bp127S8MUPUfLGwOJdjt2oQzWZIWeTux1Wiv4u/8PxA+NjBLnYoWuMXFW1u
ArEPHghuLBGl2nd0qx89evNfP6t5tHBdy8mjWed6BsHOF5W/Ao9fjmrudZ5o3qOg
nuldRF2oAZ4WXOf5Wr+PVLvFEDVNUNnnRk42LZ1yfa49QbknKRI0ByPd+tg8RxZn
tZxFedvsd5ZrN3sWtsB2keXzqE4RaOyA0uJqJHsCG0LiDr1cCzjLZY9VZodHbic5
BpYc195DkBgIzFJb9BzqBBwZVE7QoEddaOipvHoqpFwMd4Id9ljGMEXdhRdZL/PR
IEzbYqoVi3A+YmGZoYN9jrXVTQi0uqqO5s93Va//i87O4tOtHDBucXo7pQ/763uc
durjdLZBBC6f9jr8um86U3IPSQ0AW5AJ3eh5mPfm8B4F3orteoXwtCSX0dD1xkW5
w7nP3TMfwINJu/LnNwrF7c2cpUsOjPefnABJ8lnD/bhUyTDEp57JZKXSiVXDAtZW
Un1xt4jvPAEwlH6fuzOXW8r3a9PQrscwygeujhNBOIr1p47RII21FtpIPiB+x/rl
rn89J9sjGJ1y02hCdFR9I0FYDEErqNFDsfj2Za8h2mv4z1O88kM19o4KSC6opHFH
aW5dhgWLfJD4k6iovTyDRE3gs0ONKkkoQbaQgjMjZwqVBLulImuCr+w5TnizLBdM
xIl+Zjzd0EUbQ8ffVKzr2fi5m9/cYJW0Mmx5G0vXadBbUs0zZGBLC5lJC0HVJ4Th
9HNCHj9hlkac2scbrop8PhYKjFUpRWkga3fQbxWLzTI8eISvh4Q2O8AxJffJDKs/
z0y1yh7aCaoVfQOubbn3HZXT3qcBwh1vJPRwLc4suVxnzeh3aggbdJqxfcm1PAVy
MgOexv9bmrAsy2cZvcoj4uIRjEDdh6d+KK/o8QajfEgnxtv4ncChYbSUC2Ib22hb
SfGPBmm1Os3Y2SktryqKRRGyk/GlY9ec4z6eI5znw2lzd4pfUtGIi12yBIxh1ran
6Hics7g9DwJIN5n/sll1uwTrg3hvxH8uPPEZIT/e/e8tziGkeKFgYxz+IcHSZXXj
6aIkaC0t63bgmDnZ0nIOpM31N8daGcJ6rUEwMzUdy1kmt0soI50mghxx/hah6kdq
UIp8Yy3mDjDVykRa/Xmrv6UT0G/FVTDbsr+G7oRnXLHXtLsYxY+MzTXxODytF9iS
IS/oKdGpq1ri4Ytn1HrVSA72eQCfIeOO7REzvxQSFIMCeaXqHZX8H7T+ckkvQTY5
pV3UGpaYZJyC2rJooSHK0Yjt6lGko7WqxO6qFj4YW4qxdkJgliFfHlvxcmD1DvE2
XFXmAMWIT2R6gvwv8LQBkt+UssQi76axrlT2ZMKIOIfPpHSbcysir6fvKJ3Qxs3n
Owgq55eJwQWyM/rgGEqYH2ItYpbpg7b/iZVGykutBunCl65uoCqFnP20jdzPfhjx
uHLJFdo7nis6mnCuPYM2gMuQ6qjwHLqSvUemx6xaRGmkvAOehzoX0cIWK5T9nwNh
BgvmwopEc1FPv2Po/lvG99MEuxDHGf5y2lSBWRHj0MutjaCbaYve3/RJCxCVlvea
jf/jo4CmGV3Mg9KsVtIrc9uDxzSB/VZg74URiFKymn//K2ecBrVBTsw4ZKxGBy3X
0s/N72oPYt6AW4BaWNf7GEN/OmoAsvA3JSubCSvdKudVUj6XMtFEOqvzjbeVKLl9
pgfD+dguwwpSj1Tic8chc2Hb3mImKjxUc4C+1tnuRoYN5Akpf7+Q2Dd1J3Sf1zA7
/9zvdSVf2t6x61pqL8tgDEQP/Go6K5L0qYAX9HHfxR/RNnz7s3jC6Mdwf8Gz0aCW
azZVhSD+x8li63rpfoTocxJThwvk2ne518B4PEPTMykmfbACY4Ad8zoBfREiVGry
WQS/Lv/fKfVSvl4/aasaHUL7/zdzlA7I+QD9YiKwfAeR2hGNi9sF38Aoe/w6ipjv
W2lfwnKGPoV8fU1t/FAbnmCTxDXWLZ7CHCBKkxCnPN3rz9VSsBVDcg9FnFV1PVex
0/ENIOUY64zsBSofss9vbfOpR0xlCEJUe6HhMtmTWA5t2X7BDyoJYaqoJ2xFDHsK
9gin0aocU2ck91/GZmZAMv02HukVN1hzBdyQP/KUsNifiRs2IPhKxb6oLA07JIda
prRZgqC/hqVc4BplmR2Dv8j5v037mpITMIJHnojawWJIpPEMeDI/12nin6iYZlsb
0Ic+34t1AUyLCA+eBuAvlRjIQAMQCjjMovwhOfNCg+gxCFQTXIVD9vfiBpGNQoJu
CeIZBUtcK2Efq8L01qvWzk46D06y9FwFygG3r/eD7yqXr9xBGpN1OFtRf0kWjJBG
fsbfxfsTrJsHV29aPbzUBO8TDymVHZ6ESHV+q4Awg5RAILmWyPFQa9jTnvZsCvhb
fPbEfQrcUV58pkstxEuMkg0EUFaltLE/H6fTHRa0zHhZPT2L1ToNmquXn5JNTVLJ
uPkrfxhn3vgomzIdl6ozFNY13doHsSZOAmIodfpVD/wDqejADNzSPvhp/PXsWzPO
z3WH1cUtgEO8gLK7eRrOMcIbO/7z3djec0qrQZ4SCE6JWawTUJVhOwXthvsTc7Er
w0rziC2oy6C448TlgHw/f2vSR3q9h4RC3dnQesKlMDR1Lm2BliUKTy7sqRDu/3r/
RAcxne01x34N/fkvMTp7Ujo7jbcCSCN8q1znA+1RN0NeM6D1ZLq3VMJhFGUgdPB+
3A7QJRdvkM8n0yPKTWGky5Bz4AP4V016UJq010z+4oVXFqcvVgZFJqsxOqHcHAEz
MtvvE3kULyl3yqgmvD960jfc2UK3xTNKmQHafg88hnnxgXldvcPJ97dBc732LFx7
Np3hZ+IPp9cZo4LvMNvzvwpOOAmmWoHdKI3ugZa0dPuLgEENlEEzWYIiBMaxY+WL
zjuE7ZntCyaKBnUcjaXni8kIhSAJLs+ZcjL11RNSeUiOF31OYY/dLaUom6CEdYgs
YuTn1ZOdW9Bgk4yeWfGVJBhH+NoCS1a1WVjhkWWk+YIw8+cIYXTr39/td44oDc+I
J/lbPAGXbDLY1woKNPaCAaiz5AIpqZH5WDW/qi2p9/afrt4An/yaBXHcdCseCPHP
0FGFPCnMqjE6F71wRQsU/r0R3O4g3j81rD/4zqYpJFterKw5v+R6qktQ+eihPEZQ
Qmg093HFMq0SrlS2wjLIN4Np5/PKXR2/9ySLz9L9v8Cm0/eDhPAh9hTyjh/KuEif
F1DHwdH5A2q+UjFykD4HY8gmMt/CTgJvvgRtP/znfyN1oC4h7BVGOvWWb5kME4Wh
NduM/T6EVPfGVVt0Gr21m9yRvCocAj0B+Oiv+iMzXj4vWavOGxyCgemziVZnEwNt
3hFVmqoRQSVnkVjnZ0/nyod4p6AcKqpudakvQUttJPKkg83JW/J9WVsbKr6uzO5X
5Zy6JD6BBlsntJiibajBdIQ6JBKBehP6O5Q7HcotsSdt2MRFJdM63A2IU5pRRiCm
8hKPBQNRPrdOxwFqOsbCPqn/XOe2EKcd+xQDFj1BZl6NjzrXqhh/HHgfOkUMlkT8
mEDcp4xH56WNOqRiMqvpmIlsS9+IH6yN0ftNZr5/Qe4FRLvtjZo3W9q3AMncMpH+
lfBELgFk/R2q8LwUYElDRhmnEDLVWxNEzmWscg0ZjOn9ofnc20OrMly38c2+Lujx
GV4Bgu6LVZSu4J9R+mYu/YQYTDozm2WB75It5Yxl7CVPMekSZpZWpAoOW5ZVGTnF
gTiceCAJUSKFoKH/lHWz2BVwxAAjXB9I9uFZ4xWSTgJrQv9OdwPFKp6IIy51zAsm
GRjYniqHSxuGezaEROBxg6PfFNsKvBJKjLM0qeF6znLmFlmiQjfAqnGVtzP/tdLG
U52da73iXK2XFkCXuuoUREDfgwA0b04lAO453lbgLNN/XHDw2cAfAfGoBlr85UsK
IsEQxtQliCbdfYOiH/4LUBfvSx4lOk0k9AFB/BPQvKn/8xasnhGDTq1YswzUkb9Y
miLyfSQsuCTASETUMtk+irOPrNiaAlC+W6fUorVsACZ5PB2ggE8O5fsiUgTqbHSZ
7ekNQrfU9RNkSJuM3AhUgeuywleGAzIzbyzEaH7kH9HyzgmY4s9kR1hCfwlRvciT
XqPvtytiHnTmaXUJNYLucVnE/TwoyOoDxlsLtX1Uhf6uUaxEkeL7sXPtDr513AaU
wt6pI4SO+KJZUmoVkk/JPT2cF0ZaB5hwj0GTeCydO1x4BpHf4//uTAKJz3sf7BcS
IvZnGmmNAWd9htiEA7ddue6zSL/9RS9i/jUWK7Vw50DpQSSaiWpDXxojrgVrEuNV
T1Z8/9uRxQeJrPJr4n/nknGyKRPoBWc/4uPgp/to5zsxrl40FAaIojunjXpY7HDV
8Sdtv1abrz4dhaDoiXBaTpxriJKnoVK3Nad136BgKhtB/qQv7KBCTiOdzycjaj0v
mQzpUP8bWChrggRuIzu6YVq2codqnrdKeL8uNHk5HSg7IUupeya/CEitOFdEsCAu
MlB96FYw8qKEvo6KiE6qPCGIARAapB7dNp6ONhanmAbB1bDocf/+aX34xOYaOkDh
0QghFmU9plEkw87Nx1n6e18ub3fkU7sf6vtxjBH4shuFyJ88dzqibXSEL1rhNh5d
I73KK0a7BUuOYwQrJ3tuqTabU+ct238i4W+WpOUIrnVgUupIFtp0J9fsCOJjN1Vp
106qPrC0IffZIulHW2NnkdB98H6Wmgj4YSJG3mqXsg2LjrYu0WQpxDadm34Vdgz+
JEHST4evPkf4jkKS503qeG8el+boV2Jq0UCbjeFY9lf6hVsvGZec8un54Szy7tpW
K49qe865OG3iGD4SNve6Cr4ayo1Sup/Z3X93hXjeyF6zoEwAi7qsHFqUW7e1whu5
rzXrKLF3LN67jFxBtUAAAJuUjXVf266Kia2OIBmXhnXchgNX/v4gh2ygNr0oL4te
UbEZTYNOrX7h3K6OfhHvS6wxdDLU6f4tE5R6UmbLt0fHA0F0gxr9B3GLS3CrjzbY
XOvjtSJIbUD/G9jQlME5g7pzhiPeD/4ISamIKMWsrKHqYrhtMiY9fuBYhh32Llck
uy8ayr7D+JmQwrkL01iExDBdgNvjpzeyMFiv/6qv8iFyA85w8bE+PZnhGoBzOWHJ
gBxEn76VYvDv2TL/FeEsSFiA47ONooHn9kI/bMdNbqYY/+FrQ6ZECOoFUvR2M9Wd
T+L62Y46eI5f9gc0tJTE1Nv9n8PT3MWhQUt3XWj5/fBTZrxqupbsO4Wa04/1BBZL
tCZevoHIuh9j+8w0kBMBoSgpuEM3oYvZCZmXW43AnEAlFmrV5ccoCGv+vGC9BuN9
r1QULrjywKnbPJ7VJas6/x8s0HeUXXANU7iIzziBTVBugFAEsr56rbKAdzj0Af6y
vYBBeI3ZCvEic4Ka5HSw3nhLrpzeEiTJi70QQeGpgt+n3k4mQpWlSaFL/nqRXh43
uJFcQYsEzGzDrZT4OAuu2suH19L9+OJ06H5DhCdD7LL7k1tL8BKaNauHohjhFN/h
HGlICqPu6MnNqtlPldmvOepQyqecwwx2wXMjNDz6BxHDo1ftJ0xTMthVWaU8BJR1
NkZJKWA+Fv7HpaMAEGrH+ZEUieQ9MH3itgiP6aXQdftXwiI9NmK64G7DSkQZWxLa
mzhgc/DnVSgA/iUskcpz5o8/DhiMUTIn2sNcieKJf1QqQZlIuJc/8N9ISM/xAXhU
OKpDo+MB/Q4JK3ZquSXG1lk7ZpKVETJzqs7Tz3BAL1OoGTDw2uNsqhvZujmd26Dq
gIA9yTSh2zjvwi+2ehphuJX+k5px6wHPmuOxfkrkVjy4kq6XhMQvwXSCVmf/v7Nx
UoJ26wiiB/ehZDD2GyIH0+TscDBgCwHadJ1b1/uCpgf4+j6K5rZhE22WP4xSw4x+
tMMCRRG0hBW6YybropkNcpbo2nmBg/zvbi6p1Mb7hXGdm/dmgJLGYB287jwxtZAM
B9UjnWWd9L49D4S2uguGd41l+Gza/vm1alOG1J3RMTrexnol3wkUYw9xCBjDHZlP
cRlbZdEitB0O/XL9+9zAZodR3y5dZF+tj3Q5hVp+P5s1nLHhCisLwMqqkYKJKw5C
czqTlO26n25+HRhbZf69AqznXhFNtHLxzW3Bv6A8Cy7lMpbPrzK3SVjN62jrcMaL
c/NaKT9PDQMWaNbhAHWS834MDqXDl1iIe5rG4LQU0TdNqKX4TIjQ2WW9SSeN/tYW
T2kG+Zr+HiCdEMwzZjZwbYYM+q98ASkqjGNgYPmQMPhcpjE04N3Ph6UxocEfzih3
4KndljTLhx/1so7/j+NWErpzHCvHa82cWE14nopknF46bzOnuUSg2MOH39f6lus+
zDOzwH1GTvQNUqUr49k51SwnaMkdDL1uQAPWhEpvYrFWdHSDidOhH5d6e3i/9D1/
jSDaj4BQXVPYzo/7xwOzDh3P/Q3u9f7pUr1Dty8abltczgqfvJmnjXY5y2l/vFFT
kHm2DLsarl/zeYl+ZahqXgzhtAXQlOaOHMtQlEXF2M9nxWKEwzeQ1JZ+nr8t3tyc
hB68vr576BhisWTEUF/3VnWccjHKSUs6QR7nac2TIMjF5gcWIT1+E+tkyEY09OuE
ejZ+Hic70+zvJt1g6bJPynXqJ57Bm1DbdQzcPOn9GXqbgamx96BC1dCHewu4TcSH
ugP2jlejikI77Rc4u4u9nR2PEcOLC2usK8D2m6Bj2yHRYwWjGL6qXTobQJjOafDw
axjePytFTgeEAg+ckF7BYA8OjiYIKwhNJrvoavZphGW0vxXQ6tJXanb0jbhCb0yy
WzO6tgNvTN404tBK4a6uTD1VV0Z1wfoI37fJadYhuVkIN4R1gRMqpA8qDYQhXkE8
JJ9QHIiezgmHyeCDKXZvYFItm9XEGxFiOo8dvhxyxRA/Hctyk+9H/R9zLG/fNxy9
3RkPbnHbj3w0aZGdSkPbWsan6ZG0yt5TZV6TKe1/L48PG/nZei+Ao2msmA/JycU3
JeovXND4fzB8hSqKUaashXLCEjliff0PHoUe23qpzXZ4/awp0thb/JDXALzljgpN
7Mc/MUUaI4JyUDHfoiLBHkBovEEtyPwdspC5oh51Fp2gauQJUOQiosVQMVPECndL
oqwkF0Sxqstc7E1Fs+BVYCVgcO+STTA9epE7iD0PvuOqavBOteGmEXGMoUmJu8La
c3cGCg3U6lavG0aC05IsXvf9OoQSFMTzDQEZedezxreN3TkKO9Q1YVUHb5ThiewN
KKXDHnuynv6S3QY1db43FceEmPxIGxPsMs/HQYfRoOt8624AHlBCpvV0lHlrsXVj
nkMT7eNXWnr2w8BF8X92s1KaF9CGKEWbgdbfgxnOqf+x94jfON34g1KfWyqphlwe
saD3cDPqT5h/r7hiEOCyWHKk3jcRBwZ6LDfMl/QTOGgQTnXoI709fIX3MT48aLW2
wdjPN5206Z0uMhCHwk/UkLseUu0Ep84QJR2qibx9Np2PIl8BK5ZOMWKDHVflvdj0
+GxewEYvVyVvJ2E045LRlr7xWRj4GXIfz2YZQ15keVh3zr2E4ehMprYYcd8CgHMp
IN8zNSPWjmoC5aAJDVtzyBmHf3KX/rXKi7EosrmsZK8U86WKzmyi0mJ4W8xY4Pw4
lsZBfDBJiu+XlKoWy2mFZs6tTMg/avvm9P6fWdUvzf8rpi5+RfIUKlxGnZllIeup
9pJoRh+R9HJRt3CoWq6ZrL0dgixK1hdRWzQ4W9A5D/acz20Dx/dPnRo3lWki/b41
XvHkFD6vZ9DZgiPWJjXfl+fUyPBYJOwLQ4oMjiKA1MKgfvHEvppxdY5pksaJ2QVb
uOVvnpUda5Jxq9NrhM8moBGE0QFspWtYnSQJREg8RlK0/mY4YSTbkS5mz5pg2qXR
1XvAVKl2eJ6NQ1QausFjGIssPWSD68A9cDeoAPjrRwLLjLatSE++teaV+7q6IliE
dx9Nqr8WL0U3jIQrdNcma04rxYggXK0kEy25XRbEKe8Xm6oeWVHHFV1HB4Udu2A+
rRzS4xBUgUjQmF3+FPzTnIRWaDXrNVWXfJc0Rsg6L7Kg2j9z2VwibWnQRTDbiwLg
wBdCJA7vkp+SNRihWoyWIF3BYL8IQz9RrTnWfr91Vh6udQ9yanLIO1TYrhlOBfIp
XnuHkZDpHPQ++OERPX0k2BryU3DDQvhqcoCrsOq/qluClSIxpDkLV7COveQ9xacZ
4lIP9/Z5vF8rECivgB7R2eaL1MJ4AYSU8/sl0LmWdWV6MSJqiJBibSanYLZ2G30G
tBY1Nzbh80rYszjEHWb11slvVorhOoBEacRPMf0eHAvaED9CyeEy45BF62pBfAwL
8oO6CgaNfJBr2nxA6NQgWlAJTg/xfaEKY5Q4G987fzv7cVUQwmD4i8WSyyprfuki
u4trkbYQr3PCjtAdOX20Ygl7iJx3yV67tD9y0LMDOq/NGS1Hmjl6YSxISFUX0qnx
uNPbWcMbcPoQZ5ez03nZukaYLfsxj8d5kNI6h2SgRE6LrHbYpWXRxvqpaPqlLBUX
VdczX5lopDdqVC9o9QcS4wQp2AYIwDMKXpre612R8dBeoP/eVFwFnh+mwITsg/gB
NVtX4EXj6dy2t3OhL1alT6kNDEg2sDP1sp4/AF9mypkWyjBHPajRLdYblYuUQJ0z
MmiSarK+MhRxjsA2mK1jEjS4KhfOwGkRTi2Qp1hN/aCNCQ9gotaYJrOUHIvlowAF
mDOpcVaCs4p0TTCMMx+NdQ1M2tIGxZWpJbQ8k95FkpTH8le2+y0oMIWzh289rSc+
cG4ytUuCE9SPtQAuXxHrsgPJTqa49qp+jvrk8Ac5DRLIMJJOhc7QTG8FDipSDYbB
zITW83YceMoqiGKRAVTm4eO2V+fqBNLhoztzrkiU24gDfuY80NPlCZTCdL+KGuoj
sJju3mFo9rY+e7nl/sdz2hn/nQ/9trzixcnum9mK6exWLUOTtqa5brHIUrd98Er1
ClfqateotW5ATMc0rDwrj9ZLZ6gm03ZizAe/dZ32KXlHxqWI5eGX97VPTO8G+bKg
3M2qURxhfJ4gOEO9m64n8cRwaXJsnFgT9bNLj/P9nqRKqwXNAHQs3fpPJhxLvCrE
wO5D7TXPDlG02ZYCB1UC0tnsjCSjw9H/pDQzzYxmTcdbCTI4H3Uq6EdqZz7EX4bZ
BdpkZI8LXIffF2k4JpDBxekmIWI5Q+SPkq5zPimU5HNrBial/nLxuAWkIAmEECcc
J2hSeJaN6B4ysPn05FBFyOIYxq7Au7LBOofAWx4uLiTfmPO+XlseEJ8NMvwGo9KR
jq4imay6/FWntoXHLCdO/oQbC9VBT9KhkNOm898aT5l2mUcKSFEDj5iRTkZNeGxm
DbZge4/IUZ45vV8G2Gv8O3erBUSLqV6pXNwAX4sKtx9bQJSueEBW8l79cQXxYDGt
vBnItE6mFu/iMnQHwcjvqzcK925Jbw9YrnPEFlNbhLQw0rWzIvRXkmBkauEckg1o
dlUHcS1ZSpF6kph3s7wJegMUgZg2w+KqPwkywkfgYYL22XMwfUKckw8EkBF2wLDs
MlUB+qDMLc9LYgqPvyzRgRW0U7ajJZMV4gRFu4j0f14ADvXkANaOWNmCtuthlMnn
Mx1G8mxjQTkuXJLIIzsqOIocRDRj+qH8AzhdnSokRigzB6EAf6SbmNPb5FxR2wF3
RfcZmPMFtSAR9pdFv3enun3AmkE1JBQZXN/Iys/CioRcX6WWhX5IUwY73BdCVbiq
nXr0rRsz+HxZlCOA3/Y1xwHaSG2mQnDAQuSOg7drfp1JAJxJEDIqM4Qp7zp+MEew
8ldoQ4aa47iq91FzGTOyDemXhl8JlthZMBeIAlmWIOjHaXPX/1mLhbYHz5t0AtOu
hOVTAA7XGpPGmmKNbWimXhK3NPxiCIL8qIGuMEdmyCE9o/0eWj9o6WNsmeKYUPM0
1pBfRPlOZHKDoe79ftfoIDK/+32sxmKGE/cv2TX/MvUpZ+T90ZdcVulh8RVihEyV
YSKJN6N5UiR5jarX8GyTAI1UJzK4s8nwFzQu9bIAQoLCpH/c+XUcoV4xESp+DOde
eGajT70yQcsuBN97AY1TiWaIRch5Azfpix5DHA7GHtjcRJZQVtWUNBdEs2y7OYOp
EtAV5qurweR5jsnFRkSdnlkuVKxUiLpE6eCssgrqrFGJYeUmBRfq3rwEp1rId6Fc
ADPcNpHEMP2iZ8eR5jiMv7QulT5v1IqzgsLrC3r8BKz12LTJhAcynjLFbIMtQoyC
9Qgtz74EUW3PEoIc0wlEL/DFaGgx2++JrEpxBBqr/otYHmvpXQBj0HU83car11Oh
05l/u07CC51roXKuMwywDR7wKRl1E1l4W+/hswFZQHyAh9hudzmI13VKrbaQ70+Z
RzORtCXsM3ccQNKQQVYHX6YeqYciDGHit3mad4bSsYq+pg9krq30rykQ+sQHDzdn
QfEvVIAF1sac7+tGtISr2o2jbQ7DQYtXoZMFG3Zi41ZA6FU/3zYj9L2fZd2X/SQ/
mo8IGhZAai2FDmIjfo+WJE9X1PcpRBSBJyfPVV4iyWMyxgcCGST/VxYqUXmicH3E
ved0V0kZHYN+c/rsJyDXEf3YYex2UHQWL4irqp1f1jUVPlTjpn4TMT8u9a2bwOou
tbOBh9ikJKbUzTAgl/rkiftrRg8Q+aWXcLMlrLH6Z5XmiQqQ4EgJVR9dO46NOhuO
pBLGN9ntFgIg6YAh6G4MPucCh94odFE1sR1fqTMX4dT6ZQ91vID6djw0PTFrpOHO
sI1bVzEB0kNlwfaEzhZmil6D0WT3Ja7dRpxGMYvyTpuaN/ExMJ6K5tPIK0gvBj5A
Z8lvFV4hLQS2AgEP5c6s9oLlHttHRPsYbpsI9oThsfaP02KqxtXtYuxDoSXzgiYf
xhlnCKttgwUAX9hBjO6mMqOVx5Y6iRZqK3zb/0QKn0Hq5noBKnjmOWakCodA+Xx4
ytlcRCZcC4VcW6edb2FxCjmGndPR/G+s1yQ+A1pOz/tv2GAThKQBUZLgiTEW1+ba
gXh4xv+4Ihv14cQZ34/JFC8xg+VWtezhB9Q3JRqHJAkI/iTOMwHKob9pgQrr1rWi
HG07BRCh51+63j5dkY5xXA/x232KCdfMk+lNNG+1XP0HPbcxKlxTryA0yhmnEBeY
Kx8pbaJ6ttdUSZpssUn6BCXVl2hIL347K3kRX33xtkkYoQvsXPeTFvnOgQnSf7Kd
0iVE7TTFz83VVsVZqe131tyucBvtZVpASDlvCff1/DK7I6jU3MXAzr8To7Dq4kpG
YUbxLNDm4WRitj0/pb0bFcWnsDMOPHxTDG6AW/kdkdf/f3gR2f2YC7Q9mLitzVBe
oMmyydF3CQ7AMGXC3SBJUBMS5wU2aJQ9v05DcZOX3GgJ4trfncYPw2J5d2FOLfup
4MJ1BKFuxAeLsrnCK9UjsjSAYMAcaqHhhnGMLdXXEbNE9wT/L9ThoADyeQsWiTco
5CQ0T8vbCs4D+pZG00CI9nnchx62UGu2bohBDX3jmbpKjB79dDCbBxW44giLOG/c
bbV2yU/lKTv62TgD19pmw4DS8lWpXZGiS0LL2eKJCFnMQjcv3SBtHoQa0fXlCHed
bh6gWZ7vfw7HX0tEANKKrY+Da1HG64ItcSwmyfOMp2C6NQKe87LIVRjzmcRqaIJC
nyO4ccaDgoj7OOGB07pbu/NKQ+YzbLbYO22e1fC/NQ7SlNdpa48AhlLxI4l7Rdi2
bX6YZB08sglW5u70sS768DDOsVWBCavjfayUuXK1rqCfq3fQUvuaLb1jfmqi+fD3
mvYES+1plLrqFjj6Hm2LNc6v89n3CBGlpt+la4nF713HeQxb/8BtkWKZzyd/TLy/
GSnRhjwGL5k9CMvu7srAMnwuT/+quA9TYktw5gbqET2iwwFuDQpCOyUZW0pbdT0v
3Bxuwr+qQgjx2l+BVmK0F9l+6CUiyBkuod36AarTreawJiA0aBXWbEl/I5IPNYtb
vn751M9pNV5a5C0H3yywg62YAGWUBuhUQAZwnK2KGZIiq3YrjM3zro5h/teoOh/y
wT1QcgP/J0zU4JYrQpSd9j5++jk0ebZuMKfnf3/T3M2mImMiqtTqaqMUQqReRI74
t4bWuoCGwBV/yMe8uHtDJZ+NU4tixkF3qLMl6QOHvg5wE4A5l5l+S00oFcxpPV99
VsXh1NGKXjnmn19k+ZwbWlnHrfkKq5gWrL/PtnNnGnlC/reVZS2v0o3v28qXKK/l
VJ5x6DqUBF1QNtJ77Vbz2T/qhC4WfVMEejoykf82jFRACFmSk2vNtCeAStfJUiQH
Pz3bDt3kdDKc3Bu+OqdcWzYYD2G0Fb3j0eAXCc6n2R6xXNz3fMIF36DTocPRR8kA
ZSgFFAT3zX78O8z+y5kStLBC1qMf7PaCPu4h2cfbt2VSjuubjRNhcNCZmYphQkoa
1XlNt6h/QSAXK+/EvCUce5DE/U3oLsQBJe/MbwWVOm/XTVKPeaSZoxj8FLTXZnyb
JwhMnpaYSwh5ShFQerOeniryil/1YYRsLzV5TQHDEEcAmnfoWgYmWeS1Ox2Szuy6
elJ2tgvTlu1TYRI0s0J5st5K01aWa3egi660jqQO0Fr5zVSwun9E5oPa37gG7PtK
82cw6XmNQWkjxvQudUegbWBomx0qVU1BvQ40hZInecb687zQSufZPbL+kenyo8IE
dVDhAWA8C4HhjFUqZ/dQO4AhlXsizc49KLfu/GTPiwHwluWEakvscC4x1NN7WX//
CaMNxtJhKtzD7F940fJqcI494tBnHXFW6SMGo0Ztv4P5VSHBUosDyWsrNHyOldqU
4Ds+CjIfUex+cxBwrdHpp6B4q0Z8lC/hUDBkS5k+Ejf6jyjeOccU0Td5yGzHybDX
1A3Od0QLEJeIzbCieJm3gwf3WKJ5uMXfJwqzWB+9RhuIZv9mwk3iBw2suz6xta3i
hOiU1lIzR6qCqLH0/dO7rc1SgRaUgyoDYd05qH3fnKVcEX5apK0ymrvpO2dIcpSk
JcxE59C8clGUIrBItGIi72rj1HUGPIu6/EWH6Br07plDTAl/l/jLgM9a8fxLcYyj
tB6c96W7D7yifdDZAu1ytU3Yqyz8DKuYxCj5mHpjjzCD+dCPyhm7zZad5+xvahhO
U34C/cxpxK+sA9wu+Z30woB1ItXXe2PTXZ9gvkPgDYAYpedikFTjnWZLpIxYqf2K
KIhx73pDyrDoLvZvYZWFRBUCAT0yxmRUt7RQoqZ2v8ZqR3ekBvYEKdVcXwmV68qM
MsHlybpknDn8I2UbL6HyuGJWVdrGY41/BcJ2/9xngMHs1tUbZQiMOKHRP9snChK8
0n35dbS2oGX4JBaikVQx3ydQ2SrATFdf3+FzjtmI5sSYU/LpBE40JWl1kSEzOXBH
i6tHdEO3mF/iqgVJrswKMF7u4yMBsLFsIUCNv8UJUSCkoqB9S/DrhYjnDL0H83bD
fa1ixkZcKBAqQkd78ofSOpgvN7IpE71la6/C6xGfvgfTkunPyNYkv7oOwpW2stXj
J3mAMYciVzvuoVBnG0DtmpHkqOSHuFaswM0Vddz/Uezxwq2T7a/6IeKDvP2pKF5T
FWObe3RMNawUbq81pQOj1fO4I4dW5zpJT2pVMBNI+YNPjpnVA9l6Z6M5fURRztXx
sSp38csScE/tzHLeXtLYwc/+cn/zqPdDigvhzA1A5snyB6yWBwd/lvZrpcPBtgL6
SAOqolWy1ulGgp59RoZDATZmYXwDXXvP9wZ9EBZJFZBvkUMGyV7eZlkJDiihRjWC
J5UocUm1NRJRVzXEt0T3t8FsouqZfN4h/pmm9QTtn9iEBCm/1ItcxCN9JYc4iFnu
1p4/mtXs9t7wSET4EeUALVxxQ0HASl7cBqqGvkqzaQGCvTmmWN5rOEAx5nSJDpgn
wPKvH766HCyaQJ/zkQeiDkz4oIzvKV35MG/xVVYD+h4+v4gFZq/SSn5PM//1Ra1L
//e+OFilFZHjTj/47g731Y0qusIX2G6TIgzmet0xu4Jninu9zm0A/stMqXXpyWJ5
q8BPs1WnHEXHqh88eVwGAwG9NpTyZmuCTSvVpjuM6WQYTK/lO9tkwMFUCtyGxNqi
wgyFnusGDS56qlkgPMoBDTWZl2NH9+Yi8nLTMrggvlvMzMjl6RDSCdyWDgZ78M5b
kY6jrAd0D8dnkv6M2qd5Oi/1mcR2CjKc8TdMLk9IGgCn7q/Zatuj5l/s73EDEHsG
BtSqyoV95rDjrzw0cCmh6Sc7h6Q79I2eJuRpAwW8t1bbR+p3/kZg28QC/80301I9
PxWWDUJEeNuUJh+ypH2J3lOTT58yk37d8RdeTsyHzvm4fid6Lbnzh682vhqXbUMp
O5wYBjD0LR4cf8mZpU9OcjGLgxc52NVIbxpVXAoA355mJjLJtDlK+jQgG39BJTaj
D9ZK3n9mcz1WCC2yXYO2ZRqOxDiPWpGdtrr1/413z2gHxZLMpzfDv/t5JayuOpfM
FbeNZiF+7uIX7kc2fNe0OFmUf1aZQEF+LkT3JBCFKKaFhEUIV9cA4Jhg0y7vC6jl
i4nA9yWTYmAfLZRfUfwuo/+i61X9zznbbxbpwUis2DAgG+X8IL9rBAjygZlJrVZW
iLJCBoEzlNNCmnacTSLPPmEJKoj4Rrn3sWYDKwQj3QZJxAffYM/dW20gC3xL0e2f
FNBNHN9CS/5uSndhL4mHK1GtVtMtrOqhEzT62B4eeeT0+W/qhg5YiNsLcT7NxOZZ
r9tAQXdpW2lQIArjsb6RcUgi8k29WcdA+3FwMIZMSF5SALpDkPqjA/YPnqvG3MvP
1am8FG3juAYcri5Oaz3ck/b4jAb7TcQlsKCIATXYfjOJ2y4D9TmYsP7xg+NIonwf
2NavpMHUv5tZXj+MEGxThNGJvl6VIiJdQFnB8a6TK1uUlLp9RKGvgYKuZquaaqHj
TTyqlxYV8D+A8R1yfvjDI1h1NXOKggNpPdPZvvJ7Kc8azPugfy/P/l6lTnt3phET
B9OFR9Q/SeAbmQA/YGLo2XWLUTp9hrLEt7smH3qRbd8z6/z1+z17nwvDORDVefuO
iSTwXOcfYpfMS2m5vlmms/LhtLsLri4P/ENrFCYPSYg0FMPjaSe3VWH13+WSTAH0
n+rLZmuUsYA5ByZliCH3IHQ5OBOasw0tTiVKnVLvHfBUjQiaT2aFI1PoppbJB4F5
+1lxuHlSCyR1cuG1j2r/TQfyQJkgBwz5aTVj3dl0hQU6zPlN78yRoh993JqeBdNy
WN3jnGu/NUQ4OOV4dbToeVtYgMPI3Dotjz+znFqfTic2u7JjdzqoehLZHMRO1yhG
dnD2MI5eyKKMHFD+Shc5b984zb47yIr50F9PHOUL2xVc6lWEs+HTq8J+sVU4SPb1
nj5Oc/IBN5Jqlq/JWmEUHMmURcf0yTA3N38hB2lMzaya0LYtI6eRF8Mup/8v5INw
jbjI0eu0XLEZbk5Mjgn6iKsHHNEG+cutqJwwi5ArO1poGCNZyleu8mB18shh85Gs
YNiueOame0XjDNq+GyL6C1AXDBRwQvvNG7Od/RUjL2766Rm180Xtyiei2b7Plo/e
Fy/9SK8SpqdOJuymdDka3CIZQNRr6KUGrrmcQcEqCY2cYj7Z1pdxiBLIbaybSEsv
9KfXCfIThK3UQYwRdjCwGEEGaIm4EBsJq5sBXnxz7NbPy4Y3jG/WK18eVw2GN9EH
qr91ue7UCRH+ARYMn8wmI1PtJ8nLBdoIVJuZ68jjAjBBPMIoD+CJQ5Ygek0CUmCR
FzQXCuBE3GINWZpqtC7FGjsze4TLZXMu1R93zIQmmEo3Zy40pm67zdSwmVYMp3/2
3/ZK1mH9q0TLfRTiQKmZQgO3LtfMSOwaEkmNdkOVqFMoICdOZLkCGKxXft+68TJx
dA29ogwiRorqbxSpaoTzDgfArIzfy878j4EtHF/WPGxHjwOaJomYGaiAr7of3AT4
lV/YhjfVJ4DsmoW6XvlAnpr8FIIsw1Odx2LkY6JgUTdJzv95ykY0jwggxMkp5Ssh
V9TeKqtGMs3oFDBrnIlu+yZXEPuvnCf/sj4jeD2zvFLfex3soqYANlRwXty9tnbi
n8x8A4N72UyI6RrZ8VNsdZW/o0MNKgaWeoj3MeozhT6WRJcoY/nHqYCsqpkL5xSs
zwgyZokT7Xm4OvyxiZ59Zas3wLy9S6tAJkQ4PftGZIUdozG6qFjTXqgAUaWbAukb
SFxp1RRQaLN/jKeJP147yZBthEsKmwy3xCnW2frXf2P/Pxpl4WsIw8E2iNJQKDvu
TZ8RY3xToqO7TYcKcathdJrU0pLd/OUjfIMHowa598TkzLQC64Fvn7cYddSeMQ89
/z/1sX3eubVVS1Y3U1qxh4dy5LihojM7BszFc/MDUGkwYZTiv2sY8loXqmwL2pMn
GzxsFxu7vXm8iYU881ceoUXCPmyp7ji9XHtCRZ7L9tef5tRAOZWUJVJMEsOsYjLr
7yl24miCaCytpB7/nCnPMkZ3p0gHjaVqPXFjZnUXEcgbi8j9jSKiXJLSlt2h7y81
c1op2r71VOccIMpT1qBxVQ4G4disJn1D6XWlrIcrY4szu7NYyl0rtaDQWpqjdhcH
sYoXqaLwEGbgZFhCJ2LkYCGTE+EYa5VZESPpDOWraofhHAp7j7nK2a7z8tg5BRre
ZD4Vp9L/UOtC+zuBnINMMoabwwWBXOJRsMFvOH/KNlzoTeRi1SxpPpb/FQO+9xt8
szSOMcAVokRyFH/h8Xg+tni2P/W6gB3XTjGzUWK+UdTDYjBGUnA8CYpQQGO8GPCz
0U90VRuETpSOaTAl5byUY2algL+N723rQtpI6eW1019Ka5Km4vn7i2S70L7ztBD3
jSwVE47/mFMA4YKB8Z8FNXGgArbVvwuxNbHUV40WQvE6PMRJGBsjpGV9YB8kaX4e
HDmNVaVP5CUd8kOnmDPC3wiQ/gdNa4cQB+Qjsc3ePT78rXxMXoSaIV2cHh8Zleuo
Bl7AEK9QnSZYeCa5QxclYZCEj1vA9cmLOm3GQDPuPNHs0sR94inh/jySKrOckHTh
aBzb3VA3611FrTiB4eANNeWQfZvZ2cT/gNOBm4Pc7tRIN40DP+jfq9mKvBk50Xq6
Oz0AnnzyJyIRg8p2hhiBqb6Qa22ZwX6OsWJt6k5+l5i9rls2ZjPOFm0yAhVu2a7O
LmCpw6VQI7vHIj65LA3Kp/xKSrbXSbmebBkvbTuNv2M6nnZnBa02SqtPFSIKtIiL
pQcqCeH0r3SR58JFdbaacySa+cSz6HAAbKrG8+wdSH0bGCY7UzPVvVbXp8kook48
/qWZVlMr5DflWqn6YJagH39yMc9b2l4eKw/fsxAz2zjzfTE6YCgMNyinVNoMvFfn
Dx2A6kAPZfLeqF+bhACmcZyr/4xAoFurpWXunxfeQN8=
`protect END_PROTECTED
