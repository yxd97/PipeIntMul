`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZOs2cs8btsX/J77c3Ps5a2bZmTX+t3C+5rDcmEZP/m5EilfL0pgtWL2G0lqsIBT
vwB3nOiPqdhH2yYZw8D0ZCQWefUzvsdQNx1ZUrpatGpd1ZRyo1CGlIbu4sCncnAx
GyAJT/RolBSfm3hUiHSJwuHMPCW6I+ZsG27z8ANhFMCec6Kq/OhK/fmjxsZvvHv/
wibzfeXiGqCmSY35oxRX6m1ynh0gZ2uTXsvjOcIzBN8VZt90ePc/VOTajci3+i6x
`protect END_PROTECTED
