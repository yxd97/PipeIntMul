`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWvwZOes5xLpHBmxIGfxNwwx6EzlGl4PCMCaTwEFSC5GfLCN8mSqMGKGqKJLTSLy
FBpfyfu9NkZQuIXO0SqvK9Lo8UrEv5TR/tucyUDZ4XQd0SFrbA0bds89Cbi5WgtJ
yYNf9BSyLZgrUd7rdhx5osQy0SaSAXY/qixwGLw1NYKMH1SHFvj4fsde//40klF0
+Luri9/PrWijTyW5+8YKLH9iG35Bk+2nnBX0L4fjXNZWMh7tjdlBmSZlNgH3EVqK
Ek1XQ56xwcjn6diUR2kz0zaLU1pNG8ZzTo2hqsEBdYZgRWccO3P/XZFeQ+3P2MN4
k0aL1opv59oNxcoCGyxsZ29n4+49QYb6ZcqE7t2XBYdTEs6EFE5p4gculoyXDuTc
jZxFquFKhiWJrRkejScNNRvEh6z89wt9ovdlEgc2bspelmX6ZqqAIuurGVnvIt3G
`protect END_PROTECTED
