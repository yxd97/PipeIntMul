`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmPzSTrHs7BtLTm4lWKmbc3hczoqZebCUsm8gZhmPrxE4u8BfxJB6Ph19I1O/x/Q
6k9hssTD1siS2PzSD7SVZFpqr2yUoMzxDJOqO45++uAHCSYzVUh5sWWWx3IQ0+HY
Dv8T1EGmYs1zcQUp6s2VbFlPupnjJuv9KPakoOAYmOrL+c+cWQYjXh2hbg6VmllK
39j0i52ZyqlhXDjj1E+P6MzQINIPIJm529DTpdPD4ywTjDW+5vK2cPqmrSHgKji0
lF0MEbh/MFAFUZoDLmLmp9w8y+7VVqmhJYbMY0jMmJy6tHXhpclbMhfixpMD0Du3
VOkZtQDteN50VptngWhkZILz9o7AIASwDscUdH2/V1JXbidXCAW8v5lSzkcUkPPU
0pO4dCPGH2w9//H1F6DIq6FgIn5DOtKi0lfM57DwalqPF9+W9QC3u64vDWhUN5ze
`protect END_PROTECTED
