`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YOy/JdjJSW/BCwGpyO9mStY3Ndubd6EdkEZsMWcVVxc7RIP7rTJNoxMDKUAuP7E5
JhSM3H5JexXJJvFv9kXNBLp2TF/JTVvNtgrf9E/zwnuisjQs5cK6lQvB3DRUG/X2
B8Rxl8gBLqxnF0MjwxVpj1kiu23UQ/taS4M0eqZ99Zb4gpjvbe2BnEtSpVYMOWxn
KFPnr56nhTqjBB/2GkSK4XyApBcAX5Pllk3AWf54wv6/kjTRovd+RMB6IOZIrGqu
Qc7CuHCnEGO1A4AsK6vwFu+pcrIb52BNnhCMxw8zcO9brJmkMZMFZt1j48SYljZ9
ZuYgMzkuKgDZxsih3kyYVUlvixpMqAKfdTSj6P0TyD/4ljscuqFPTuQeID0yknIJ
uvRmE91frrPnL1di5KgAxObxEp104AcIO/kpTxPef8Y=
`protect END_PROTECTED
