`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/P31YMZzLKeO7BH/d3l4fsRBV39Fny6ZssN1Lg2ArTguhl3SfFkCH8m9omS8ZON
5zx4B57Ywgl0MLd3up017lsnjFJ98vjdZcmxaDGp6qT/l/E71LHYE2SLEwbHlt3Z
jirTvxtADLaitjTDuoimHHIaRdaGn5CNroy2+k1ZQrv3IE6Q/A2rMnyNOrgDNf+X
Wa9KoswL9q6VFzPhrIIwE8x6yd64J9wkTZqVNnq/gX0GwkF1jZUIuLbYbNYwvBMA
0lQ7Tw84zotuq6LXRD/GLFRvYSYDP0EZ4Qtr9wtAcV6n3o89frJEwnIkK1J9JpJh
gNiSsmuxuJXM93cZCjnDu18fRKA93ICa74ERXG7alB+ehWQ2WWu2pM3Suegsj8B/
HQhSsWUvy6fUi05JlBAvpifImvm+VEJre6RcK+Tl4mUiF+LDi33HEkEz1nq2C+gz
Qwqboduoa1imUAI4Mo9dIAT+3lwkZOsErgqZibrmwLYyvOwH59boDraAnFsD4DfR
TIjFNj6Uufxxx5404yptFdk7UctXAufos5q1lDUICLlJ7Ao7sCT7GP1/ZUEia6Ze
ercn+JAqqvIFwNz8DXD3Nr1MEnVG21Kgg4KepaNyaxMMAis1jPMfsqkfB02tIBn4
yPZ+ZpXa3ouBiK7YvYX5oYTvBZ61UNUfhz+m413NlM+SyzELHZmWx+LYhm9ImJEl
cRPBD2u+OAYn9AJmG0TEMgxecPGlWFllWrFpnRWzkpY=
`protect END_PROTECTED
