`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RSV9AQDKphRTCsH8mdKft1Bl7bOoW7DYujt5XxKaqZA++Ng93bzKfaH5vp2oUi7S
jlTeAUOeYHD71zVsKafYj+uik73CSUzBcXlywxRJVWmXwAu1lUFzkotxgp+a+5Gd
k5iC4HnNgA5lhw8IotPWpx9CQH1cy3MlGya7ME3+pY+3hS46O+PB4x3Ojva0rZe1
iYHIPXANLAgZleHsC4eUHL0HRUyluq14bfZTB6Bx9/rckaXbDeYozv7NiFLYJy07
EyvBJrFGc14VOUFFb65Ca7hHDctF7XTfBvKi40FB02c=
`protect END_PROTECTED
