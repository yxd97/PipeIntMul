`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gsYdoENkW0jO7V6UNUdj/EFVmHS4XgKvf2suAGjg8P39Q5GZfe8ct9YdYOHpHBhu
M7OsvW3i3pcxybfygT0sviI00wFotkN61GvQecPe+PhschXu4uC5lum7jBgk3bQE
+6Aru1PBCUTPrT1pDd2TrzVOIK0h4838+ArpS+vrzCsxLIwRElC9/1Zme6Ji/ri9
fEbs1X1I48UhDXurY6rnLWO5n7ssKwWHSEECgEeDYkx4p/dja6udyiHd34spfA8x
McGhnUtw1E1dATV+iK57ReJxAWxVEZ+ISOCDfUhuKsDKTTE+0woIco7kfth1Ztoj
PwjzCBLHvR6ZC6E3dshN1IqVRzGQ8n/xK6a8Ut/dELLEMZYmN9/NE+22i2lmUdPI
hLkxlgtrKf2TYvIsIUlbaFR5qBRl2gyGG/wH2oOQ42X3p8ZAhNMSktGMTy3YE5+o
nz1vcmTy/VVdeqpA+6a4B0pBI6wfe0k4RprK3FjvL5Yb/dk9mFsV2EC3ZUCEwPA0
BuSJB1KJocaOUUeOwKhPNV1HsWXaoUpWoMv9Aa8KX9WzhvaImCU7ed0LDOv/jNG+
J9RBQGn9tlR5qayX1j1vc49AaRsppcmXbrbEfRotyD8X5vBFWbAPpZxHrKivSZtR
QR7AAtJQKrHwGLjx3Wzo/UAjaqbHSq1pisIn38mUlqqfvOnU3NAg3sKhXvdoukkq
ZTVUI2dj5QgDuCQ6xJon7SZnUol8Eobjxpx+I6dYDsg8QftiOPyywh6mxFAyUfYB
GvzrFFeBh20M/70GRXABKjcBMwbH2AkdyZ8MDHK0AuAG4rTR0z78Hz+LHCG1aY6+
Msdzi1Dau79pyxnWtygqCR/cywkhIyrfv0H9L6sZAPCA3wvwkRbyR8gaKwP2M+q4
GF6k2gHVRum16Iv96zcrKMc6738f9EvZE0lVhusckahS8wqh50n65xJcElEO/MOM
ZTH6a+EDvLT0U04/rs2Dx/KON+UKni1+EJG8mF4gYa6G7P+pnnCMNcRgbjM0pqgf
cAhmj42JIGtWHZVkvCgfWWq2480pI6gL2OY9PBER67LgsJqOHYHausLg6a/4cFnn
cLmWG2wycI3s+dUsjdOQoyvZjHSTERyZPgEHJTp7bsQBDOenkBUomH8y0Rp7nFse
C+AnpcjeHi3gBh2Qgoy512FyhgUQu1VN5lExlo6wmJt9kR4r4A7VWOHfQneUf0ho
yLzTiSrXayLFgVXao7piUbbKjOPArPcKtbCyPPY173psR8YzMW/0cCJSWFH349Fi
7fzuhu6hDTFh2+MkceUwGJrLqRxnIMzpOOO/MsatJufPq0ghoPQNKMBaMMpCrqm+
erCqr5raCIiVJ103Q0tGJkR5PqZFd7ypwDsmywe4mAxcW2lO0OqKxk2jppVylCZn
ckcT6sqqxMqrTHrKuB21bAcXVHMcEQVBElxjkDGkEo0mK4JPg2pkAcdRqeoAW3zy
9a9LrEB2daPTYPruvbV72spQsUVXKbQw2Tm3TugT7lU1tRD87X34qbhUnlk4Lz5e
+3rguHP15gxMIdoKw/BRnSATHSlIKexZWNdcjRzzGXp7sNE3qSU8Z3R6awkSBmVf
0cRjZ4rIipwJcZDM0d/ZL3ziljgJqEeh4Aewq8gLK1FiI0BiWQtyndjUV7lBHsy0
+J1AWLg57JZ8EggPrncvBEOIHRvYzlinzW9XiOLC6nAI8xPypA49UO35T4N9y3v+
PBwd8pXJJOTyX+39x+0FkIY3ZJX+fOJWksmE7ax9PyOk4pDPv1degHP3maq8iT+B
jbqYh1+O2KNhrW85NWgHNyiYS9KW/KIry8v8vF2B2qGqRLPqCJ6IyCFd7ey5dbiK
EyRext2XKRG9huDw7RpRckSYYy5MT40sAG/TwLb7nvg/J1RsCHFfFHqQKfN74mv4
O82Bj1uvX9AUAPv64upfUqU/ze0QcjKNOpVZIqcFFpm3wkIoIjWhytpZfMJdO6Oj
gSmHrlTaGA4JcwPset0cEDdtUDaml6b8sKUZjAbrrwIrcw+mJSFEdE4Tohmqt6/j
Vlk1f9K9Ta5qu+xy9P9/XK1VSI0GCGoRYbyw69CmSSd9v0LYE349e7rxaeZ0eIJS
0DxIx1O4NlexnqybJGvES4Q94Vqf7MrV06k8xwQ/RK06qi0DcxGKRLGmkQqZB7nF
2gw+hnsfxB4hYm1VwfjUAI02KCg5D2PxPlfDytHKEe53i6+n0Vskjmfe9H5iw/hi
z/vSN2DaK1uir83JcjlGsA8UDsaSvdQGnoLigE96Tkd4bvWgnCC+K12NN8Y1JIUV
EDfxnYmkEJb/Fu9kexkQI9SlXY0qLfaMRqS3dMPkR0pKoY8KcOuq3wfMI4Qds0fU
JwVbRmZBBhJmx7gFb1rJJx16jnQJBVOmoZfoEcUOBJ42LHO2zj5a9CIvU1q7M0ug
z5xEgpH/uBdsWDURBnllOu0+ofw1WjbGZn+qZgNTPb0JPgUyue90pyIMWdpoxkyi
ncMAbqQSDBL5WWHB44i0qcdkx/wk/c7K502wF+gPOu9bm6y9QGU4yzyjLz8bH8Ts
2rlbP2Oc70M8KuKNTGRtM6kx0YegwtUlmyWZ/z8xOZRpuolmwSmBe4jlomi0WFAD
3sQGNfoQi4uAiMwBZ5TY8yDXjyQH7Wkh1LZG2EQ+wAUgGJrxV8siNM2vYh3BwrSP
YUR4/IIdc5k4nOE1yxBZBr5nB65VJL04AeiqTvPoe2oPIq22m9A9YLk24mwVB5H3
Nwlj+i01SyxniLlZ+GnO32Fr8LQdi+LxmuhD37rbsoTw98vBKbVYMIHpaiketT3G
uIbiQOK81AerWGXJhpiVMMu8wY1lcGXuZjoL6vIklq5rc3giy9DsdPygl1t8xuvG
d9ZVNSAU8FOFz2cGFPhTKr3OyuX6UWQGmLGbRbEkcrG0dwMQlW4QQAg3ZXeSQOa9
gf/1bZRbi8JqqfBQU1TRmCzIptBYhGu76TvedhJOmDlQuxFCgnQZJ5CJel3JDDa0
R2oOool5wOWufWmz7ZEwesLmWuvzoCQWOl2cdAU1wQjWGJFFEyehgMwLFJYy0pFP
UAMKQ6M0LggPfnizgdswILy1CWogP2x/cobfSTKJSe3UjYAT/z5S9LW9xfO3CNzx
1CjUtVe8hdr0ABriCJQeH8YkAjwBsXo7TrLCFMn26aAmdqwnPiFyw1f++Fc8vMse
RLdeLh3Rp8gsoeRyCx9B99JzXDTHpHB0Hz0R7tGyhZGkpqgWDadwfcznRm8sqJXC
JwGh7tivmX7XVDZ6mZH9xE3ulzTliOxjpV6jfOkAD/nW+Y6EqmvWsutgzJOWb7jz
jmotyEabaBkuwZXQECCo+P+UUSMwVzgiVmKxg3s/dIbjIV9h+dCUdEvruFatHvcl
vss5oP6PoTiUWbd4M7rJypvAGA/1vZXsqCkpltKzHxw+M0lJPJqvp+s6ZSIOxQyi
Qa5e/tsLsEW13qlwk0kIvC+dA7h1z8Q1Lq7Tkey6jQYhR+bLkEgDXVS8QxgRIrFJ
fm8NCLkPYwM0J6aiAOW6qFUJwEDh8oJTzMOdL4DgxD4iusPxlqZSSeWo8Oh5/DML
FYkXYpdE7m1iEFDTwQVtAMqu/cmo6Ajejf35Auwgdny0bVqvs+wPDT9pf91fOAbu
12pqmromD1rtV6oP/g+qhOa+qbHALrRa7nq64cVD8JipADBuzM+xS55uokBGyjzr
/Zix0wOEi521pNKPEdLho7Cu6GgQdXM0/LuteKop3x5C8awbDivs07oA+1WR4rra
IrmiL8jSM8dhsRTrttgH3KVdXoCjV+YEV9FhrJ7ajP1vHj++xsWPKdWxZRu0wo2h
gxlWv1W5q0E6nRb24edECfYb52tC0a7oIU484rG79bhHzFnGc5OdcZYJ3aPZ8W6j
d+k11xvlQEMgDRDCJS/heHzPesnJEFWb/2e1XfKokXdLR4WBM4E+BhG/XAS/FEtu
haDtzTgsIU72XjN71FPhfDpcorqrsATenpHlD/2SBY0gpkGvXlH5h6Dut21kRzY5
XkP0QHqVfaooH+x6Hed4CMmWKlaWWLvBfvlKSd7BBTI=
`protect END_PROTECTED
