`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3tgSJ3cuq8kCR7Oue5bGlcUFrRTeurpoDlcVoM2C7D3qYYjLrJyLlewV0EnX1Oo5
Ia81AvKJ7L37Y4uRb4RrGNNiDTYKTKX8Kfu/DEfrBrkvaSWedmwBkDnObfz3jllL
1O9dPH4qigSrmWaCYEPb6f9SVSLyySrVULk4YvO0DfW4D5SVTMXuf5dk/05EgFUU
APLcn6v/lsiPrmMid60E6kkJUP0ighjqgOPIKuJllOBYziA+BfP2nyTKCQJwR3NW
iXsn0G2CyYQkrvWTfLZ3E4dIlDTeWMSh8ghji+9H8SmjK8d3QMSz+yuvn3cr5pUb
CIHYfaw2OEMMbM36mtcH+6vnCZ803YoP81ZZae89r2RsmmS7ydkkwYLk7t5zZcpx
J3Prz6DRCA6CHAOE7DuJJMJkhLFc3LPmp8BAj2JswY02c34Jp/HdiNMzWKUutJ0y
vV/JP/DHVa3mgOSyjYPg1Wut/Yh3iF55H1kCQWIDCJOxOPAiFSQPBXXDXzFpD0GP
bjgjck0rE5Q2UqfufYKDhg==
`protect END_PROTECTED
