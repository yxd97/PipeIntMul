`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhy+4hKL1joP7DHlp90FZe2G9sn777wOLUtjO7QrwJlCj8t2hbHFgVW9Q7LXgaF/
tXvdemp8NrzUkFgjAitAiqu9It1pa2Plwrw/8Hwlu8iMAqDy1dBG2+sqWCzqvp5P
D9jX77CjCTqgZXs7a6GKbAUZVI13diFhGxIiGQFxHu8urTyJxatw9ymBFCzvChux
wGmzVhTnK94lCZGV5dqPG2FGVOzLoQAXfAV/mGzUmTCb2P5qbEb4uknelDXHTWqH
`protect END_PROTECTED
