`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IYpORh5CcVk7wOV3Gtd1rCt/biwLf/LUNlIPd7apXjAL0I5VYdeRSqFgWcfaVwOY
1FU8YLCYBv8JcVoIQTRdvS/lBfxBRVIAwb09QKtk7c7KIuzm8WMw1rhKGrfAifH4
jNAqqk8qb28pUmVoV0dF23zLdx59XP+5XLXUpNl2jfeBx741W6Gzf50UKEnXLwcG
P+pY88/14QXDkrG9ZWYbNmmzhWEK6a/RNQjSYQDTFHmoRnugXQjEhkunZnr4nEeC
WH/0k2YhPx4YFIkb6RKnLJBxYysfkFJ+blLT0jv6QPyeOJyouSM0Hf8fQtYhaOxB
y3zCzgUBRZeCXqYdW0DIdD3/gnFj6rKB+nSpO0uQwi+OV568AY1n20/dV5sz4IAJ
HiFvzpe8w85j5gCOAszGVAhPQBZvX5v9qxUJn4IybFqYmdGLXWOmkPSE6Yi91acD
BIcDIvK7iRAnNxBw/7nY6/ynx1DV+D6KZQA8A0Jpa1/SlEYsuxyanrB1Bk9uWwQ2
MJ1Q52+f78XLcgtv5eSnBiSQof+Ow9HkBus5Ga/WFIocNnv7n6yhlZgvvFokr6yB
Z1OXEdQ61bbdtW/URF8iTUrTkt0sDXgiROf4v4E+Jv4b4BK9FiddYXo3Lt6T+WEI
uLNK+YK5+zpnvv+BIYkGuw==
`protect END_PROTECTED
