`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5wzcMWuzgDD/tMXarFfujAXQPKqht3cALK1/vjP5xx4X7Z8NwgdkGUqCscbbzXIU
oPM8CyFcz8pLt9d/PVYYa/1kDcKcMWhkHV79f/unKIgPXVJDcWW6V16tBNnS4rUc
jwqsn4AUoKGhwCxepWduWMJqUc/XGfVhYUEHnVnf7QlPwhheO1nP8XrR5oCkElNE
Tn8u1NxNEFhvFivoma9pMcyrcRiD9c+4YZY8K6UvCd8U/PbwmkLMrczeIBiVP9Wg
KcZfrkDhK0lPpd/9of7w8DcVQpzKQV5/VkqF2cQLBCVcuzMG9pki1TUWfIonl/jz
6KBXxON/Wkly74UneUTXGfXXAh4mKAu5UxUtosHQWlFUPYDMO/TXy/KwQInbTBlI
FDL/VzoSKPxLhUvMIVDZt/+1z/qG4JAZwEpgsFJAFWu4DUBVwQbw9+DD8PAjOngi
OsSkTlAnOpDgsYt5u8uMHC4FlHyBlcNfmVKKaCngk+Jzx1B6BpfekRierUS/Nsr/
`protect END_PROTECTED
