`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20cb2YGdZf8VUeb5RpTueKZHwjvsUd35B8859dN07V+LDnUEdMu0SVZB3tY2djlh
jlUKUzJ1KrB7OmSlp6XcSTB7GX6R/tkwbXTyWJWeKUI86yY3lbd5Wv6D6o00cPJA
3L19VDoCIXjOvMqjBSkUGEyNc0/TqogP+GZv3ClDY9r+yJV+MP9HPwhKHQyYjFMH
1MIfuIUplW8KDdGgU4xhK7oUu3/1qRl5LLsrgO+2YoesdYxOkmOkzZ25X53uNggV
bnBG5dsIBX4NgBBNdlPWIE0b1YAVY5Jtze7bcofP9OD9Ne5EKILVcKkGM+vW4OY0
ygIL4TDKS7p06WFvi+y1xNlacb8Mzrxg+uL+ELzkojrck+8yX2Gi30+gmgWLU35l
7TqW38tAVh+ECI+1ZHnV3ccP/3JNF6SO7CbkrVror+v0VNxex/W1DCt0aLwzRX/S
0V1N3dPmo8cNBsThns7wkNv1tU540wY7dthM+VeFoXUlsPgmfQ7glSnRctG9V5vg
RiY+BBjD0nJJNPzL2CaJWuMH5yrV2pW01INrNcsBWDg8yWJVA+Z05mBTpzvgLgmS
5pW5m0q7ORoxD1Ip7JuZew==
`protect END_PROTECTED
