`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r1f52F0UlmdOkU0fiIDgr1UEzc5l5H6E1TBMQkB/W8CFc9dSyOX7lrMe5B6cYXuE
2jW4jwTX2rd265ufLJVpdQsXgpWqPazG8LFI5Ha/BDLRX0UBC3qqDFdCKPX6/DFx
lL1PFzsGaX5iizBs9qT0FibZMScA7/oFxSPBNeAixydscAlUw/nlaIE5GL3JFk+F
03C4dTg3JlVmFtsvUIoqIc8HTxWqQf/n1kqgnXdKzJ+WqFuvYUZYqvLn34u38aYj
jV+HSz4sZFrVmyxYyOoZSnALUQ9nUsgUS/Jqz3ob5nfaCAuFuTaCL1QrhQz26G2d
VaIFwkvqIAm9PgJJFF62W2nla9gRWeyJziKdpNbpnLwvTQIWfkrxrTOs3X5qHtAu
YeX0n7TkzSQ3i2Ta407+SNRwAP177ZammaTYlB2DlOOd4kbLeQiyuxI54AKdMMSD
a3KKkN+QMtyNrxXOf3X43mFEda4L7wCPyuJEEftQtqIfKLPwVHVCE18tQEmkCZn7
TmGMNSXF9aWRzAMLuOQ/Y+snNjiGl/Ki+ainaTGEbhVVKEOYLmqEhkm/u0vxDyk6
B2aZP1npCRBqyYnCftFdVTmFNVm4mw0+ehuHH9X4S1c7EsszOgtYMsyqEGcl+ulU
OcbNIZtQeVIwc1OZ5aso93KLEmHUC7nht0M753mDZrJdq2cqd/cdbIWRnmrwtlm4
/s3NpWfIFUnRuffMRl96dO1fyJnUbbWIHA5UIRoIwMQoGY/RWhL3e0bzWbfQvSj1
hWcgtJoT8OamJ5zICXUmAg9QWA8NYnHV5CCBh7kn/gFNd/5mGmBT3sxQoxX55q+3
BMgzEajwcXKsLPLmiG5kC42r1YK5z4NGwoSGwP91e29rWjmqJRzfwM03q1E7meyq
PztlNJOizCUDVvsxDO3F4al3icnFh5vOi6dN0F1MlA7Qvj62FE7mhu32vPB2QXz2
V9qmFGaVt+LcY7osM5F7MoNMVtzPq3xgDuJ0FFpFbzE2qSWFkGAd90ntTIruWjBy
PPNcjM08OV5mAqCiHrpRBGYxk/3ZA4mAi08dbwzaMKeO3PJ0x5Zao8Dwq+M17hbJ
uHYbYVc7Rej9555Wz3kspQxkcDKKg/Wm5+6NPmsKAw4bKSZQR8EfBcPILWU6jiJN
Y5MgUDfcwtgt0L2tTiCWX2SX+Xf/8ndG8BuWbdVAYlwMjdFcYOPWYtXiKAECHN1W
DJQjFpBMEltqlPyriTOzfV9ZiA6SlDZPTvM6jbZGYsYhtjr3Iy9ZzRU3rHAzGKlR
8t31Xy/+cOD2BxjEVj2l2VFnh3QSjfGgFyy4uODKXD2htqNHzf7rqHKXhfsf8jpc
Xie5CWXU67mHS/eFiug/hXRaCLE9htcwijKng0mGmbTU3QZmowCPEuMSDW729a8o
5b3MlB4T7xWcLsDwBMjQDVBqlmtEkmn00sBrKCDSdmJ3SjG3So7b/AZ/9f5rEBmT
s4lVn3Nl9Uyd+/CWiBGqXE4mWlLzjxThwVN7xnAKEtooPJZgthJf/pv3qMSxTkRH
4vRVeKbHpguOuiqmME3iTgNLC3e76DCkfl8mtB1WW4wp0WdXN1AaW7DYwOeXwSnD
E1iin3vBz8B53TQoAf6+7nOZzOvpFb+RHpEEdNiEsWOTb3dPeq+ankQgW6Mz6XCD
5SqIlgiG2/y1eq9zz6vK/XS8lfo8jyiMTsRT6y7gi9Ubo/UrflkyYwy3GKPjtGph
hOym+AW1m+VNezOqDA7h9AQ89VkSbsjFF4ddTDbAcaNFBTVpXR45cv7gSy8tRp+s
b3DJgC+U2dFX9NzZ05YCuSGBMoPeP6BVCCTcnosNu7fk+TV5PMFOggPGobJk2/kN
9TZod83eP+AIUa2WpslHWsRSmskdI/X6fx4AnLb9JO51lPhzPcUkJwVG31C5wgSV
1jHrL9WQv/ZALJ4NhrKB40TZ+ErmYe2CJwGNEvryztETasiQeFcXTZFDnOQ/cg+n
O5YCQEizw6IZVUFh0BJFt9WVZ6GGK7RhVGgmWRjT28gNr0Fe4RxS9FKdeguUNHAj
rTPgqDFUK/yGQmuAyQ50nrtPgJmuUNt4sN/1vDxYf4XEi51pfn9QXABlWhgPmA3p
nSMEr1ZCd/k83tH4yZdZ9Psr611coPa7X0yzrljV0NBKTuOdxxGBoT/LmgAePWkJ
Kh05twPaFkRNraWsZNaidILu/tkGFWz4ha8lIdi9o6UqalDTs+6CVON3W1DxsD+f
KMh+/eExtxnCCZw89XAVA/nfQo1P7fV0+rgac3/yV3CJEAPI08SiZz8GEd8HSxOm
kuVfyDiOi3bYDYRluCHYgJ3m15AGYBCoZI6qszlNUxqEIgDYL7wnnX8ot+j8sSv2
u6Uc6g73ZzkkTus+Lds8BfL2uLLnVkqsSEpkyHRoXloxH/f58kRlrX17SSEn9Wtg
TjsL74w8LLllA+xbmsIFPAsO3wAUWeeYHyrHy03OQWMq23yk5vXKPfHo5mG3dg4i
GFC8yvQVCE5GOrw96LxqWUCVnsGwmbSnhmsxVl7Us73XkeSoq93yqOBgjcZ5H16S
BRdAzYhVpy74+20S0fWF1/MrikxIkqeAqJd3GU9azQnS5mnWLsb8H6ymkIw9c964
eCb6XL3w3iJjbrHWmbQTj8dJpgu0B38M44SgzWlc2krn58oV/UjMjOq3jqyvIxbv
mrprSilusp/tXCn/3ho9ArHC9UtSMu9wNqwC0zpByyEyqup7ckgfYjGjJSIxpEJ0
lw6u0dOwjVXTU+YZshWbkXUj7LqKW1MpF14620mRgXPJ7LsPqz80Lj9TfDa5hw6n
rF9sliqmzcTZRWJBA4qqb/VWoSCnlY14KoYHDd4gP2FgYlOOXReoA5SCrWGQ0x77
`protect END_PROTECTED
