`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
91TrNAcOOMKE2aYdQOwbcEasrcyBaCE2nDI+5auxZfTStS23wkVUe44Ii5lu3CEh
dX2HNJj2xzwTDnxNYiq3sV3ybhUeWNwFk2xzKimNDG6G5MMNgDxfuMNo3EzFmeQD
e7cWF/R7ovkUkcxg2tPalWaJ4ZxwbPpLkjEE98V5/Lhku+pIKlVBaYPqfLIqrhp0
W8c81hLE5pdGadLxb47Z20Ozdzl5n4Cr+/f2qrb2uiM21Ittx/2ZfTZd5dg8fQ8a
uBToWncfXgRY0uaHCKXTglKUudTqdqFYjy7wSX4YTX46dqhQ+tRhQnTuUsVV9tGS
AnPR1wMwpGQWQJWQB0olJCRmx6oJgGN/KI392L7I4Og9O2M8bgwZWWn4zUfKarMO
w3EipC8hw/kZells6LSNZhF4cw9SmlWo0eN5HmvcVu3D7GA3G9hb1XF3iRZ3F4tx
zaZdND2mDiOibANqF/BZi6D+kLzkKs0EyuqvFrFc4l6JAeayqHoR3iHFzKcuyDYq
RNetdmTgxuvMLcN4bzqRZrstFeOq5FGDJiBT/8bXyAvP2B2Pfc7/CutGKMaWRT7n
aiqytuSeGqa7U0rKpbl7PJC88Z3rohGH2O0pgp5E0Q6bdyXSdoJbITNE5DBzoG/B
SDTeyfB4fBuuFaHTYYZchj0Q+dbgRFUr3F61Ubb94Ombj2ywwA5Wk/Jl36GEueAg
t9Q5VcWy9cLejRcSR6qY89d7fyvOv8hf8+uOIIHzioVlkaA2xlNtBT8FGLcsZQBk
o7rFDbbW2rAgjLOBGVMrZQ==
`protect END_PROTECTED
