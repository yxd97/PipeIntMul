`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N90eD3kzjVEsG+ROpkVcuueEQRAVNdz/LHusJ5gEPlpAf9b573ok2wFK+vrkbGsQ
IIk1b59SnnC4lURPQUoL+ZRmkHynHUZuh9SLZBhQje4fIwXZXgg9ClS7Ct7Ldm5v
ozPodO1iFBPGm8V9NgGGaxVYJVlvPPWQRo9t4rKqjXaDikS1/G2XHocNnhwwA8s/
mv5vCC1exEqxsvnMZPWtaCtddObZyE1ysxqnCat2q2VcW5bmiafb/qL1Pr5K16jA
4tAJ7wn0WDW7qauZTL2cwQcsJN6PUcU6mrjT0qbEpTVWD4lOaVNlPpvPZVvD6HaQ
K5IjfHeBSHFEVCwQ44FHlFt6osR5Dw0/LSwVceqfTHM7X4WkvjBjXWV9Fab+ZFJK
bcP8zw5faLMgPbYUXHJEc7F+R1Ah2cFeQ0Ucq/bou1/u1jv3aQgF1m7/cZ4U1KUX
LTsQnfP2vKGXEgpx44++yUH1BbU+WLEe9nquJMcMNSTHRcFnjtMGuhKpAwXJIAhC
pzSByanQbYgx/rDkOWKe3rSVaZt4mZ0T2Qr9GRv7d4uF6mfr7a1zqzfbGEnOmoP3
xl1r8rnZ8oF6X2vgGqLBcRMYocU4+6F6Xyh7d4sT+BJjJpjY1PFkLrkvbHQ/Zc0g
8b37DPZj7rh8RQUftNCfrjZVW1xRscT9G7SjBsef4GSfW8b0F00Fj/8MyNAsFHrp
EWRKNmWmU1Pig8z3GYBcmG35f6pbJnH5DGMjCyVwNInMz+ZYkwRkNmaIhbm67XuI
Hg+QixBLjAHVFo/5tviJkhAsyBSqwcf93WKC2GIjVONIxuWWdkKhSEj7yQ6qURhC
j64jRLh+58DyyxEUmK6ZQafAs66VpsvXNJaq+YrqClbAl32N6aWgiGeDJrM7hats
9DmZyHcVG8csTqt7VC8F8C6l8t2/h3eHNt4zSr+uNax7cg2bF+VrhPXQDHtUK6Mb
LQ2pkLyLEoSshm1Kq+15dTGVjCJ+DfuK30K/zrFJFA27InaePuhP+TUvXWsTX2cU
oBLZlr8GgOUFWmaum/WZa5z8VRIE5btVk3w3kRTKkvoYir+3GJzojK/xwDK/a3TP
E061mRwNRHot9B2GO6oIA3TYVUrFb4Wxq/Rb1T9brKKjsj8O3DDj6AHzREV1p/1A
Q1B1kyq4HQeHCk+17CJKjGatrjojUGp5aiidrU0NNJXbHfFHiqqJhBAsbxR2kf04
Ldx9EysrgIKcR5cuS8HThwaln6Oo3mBcixvkLpsr+SAha/4wRafN0oCyVUx9G2jj
37+34rod5VDM6xR0P/wq26pa2GoGcqbJtJd94hhKIxOKIQTIeTopOt0mFPyq47f6
Ebr3llq1I8+xUxTyXI1IKz20RD3MMy4cUEIXh3eZpWnEs2tkPm7NF5ZlTb5JvJe6
XJJSaFIiklLhbAvuGPm8PzxabSyyuNNS7fDC723lDRKdVHMSgBPoa8rAmdSL2ORC
ULnPhJH0RzG5tvOfCk4H1cznfKXlypbTdDcUWN3oi7N0RaXZdSsO9AHnafogz3un
i05ZNod2e9iFOryYdrwEL6Bv9+2SBx+Mka4/VSleZmVzxfrOQs8YzND/R1gYnBWD
JDEb6nIMhOmtDdmY4iTXoB8ijeEOMf9pI90ORs01rVP2/FQdC9hq2T3NMEfp2dTm
KylsS8vqJz+0fYP6eZmZ2W3WhARkt73GqucqGXon9lxPQwYtjGZqp1we8VWXYS/Q
BUtufZUlEb11MGojp8lL0+lCsQoK0VwTjUAqCyWI7D58ebRMA5kpgk2WZuK9z2I0
qweG/E6oJ65d8UCpYd4E2y9VSckDPx96DSdB9+vECyGVuwjbZGKfHLvN7Jhhmc3L
55jl+BZWfg8qqm8NwjtedZZv+edtlhGG6oN7LtXZskAMXGlWJknS9GoEWVscBp5g
SZudZ2vK9/2WfuYRzEzQB6d33iLrz4S1+u90ZRWdEVn9fir+8vmrDPggQWxRTIXU
CKqZCsjZbrqz9Tz7vIthHsgFyNDf7/S7Y2KJ3OnKxjWkSiacrn6JYWCaRCDfO6KN
hm0aWBJN+hBXB/wEjNjK/Iq0GxF3LvJsj7iZoxxkDmOmFvl1fDi+mBRvOYu7hyAo
zHcr0qRV0SbpdeHZShMARPkji2bMSM4t0CX+ebkCd8zfc+8ohruXsQPLHpd7udPn
J/NO0dZ4yaF6BbyQ+hjenfYTE2c4U5ULoWLSNnslDWULb1yAKvvZ2jQhZ7r/4EQu
B+NI1oNAYF/oqost35m3kgXLpgYmdv2aQYj21htMuXlhS9WTbBVdQYGlSMtogPdo
UFy7Rf1Aum3U2fQpcef0/JLcOyK6KWsJ1zwhd91vghRNYlszXSK/e0kdYxkW/Nyy
CyWWizchrcUqqQVoR60rjKW0EUjWOdUEEOtdGcPZRrL9ZitW803scJ1bA2RCvixN
LnxK5R+xuO3yMu0WuXDMfHrg5xTSAVnol+DGA5E2gyS37fDPME0Q5CwarvEnhT3A
AHNT/jSSGP0uQrP0iQTaog==
`protect END_PROTECTED
