`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6NauM5z0LUqrgLZLG/XbD3FUMzAbuAnk2hj0x4LqgfpfQ16XU9mzq133dmbTYINE
euNKDnVDBs518ABpI4sQD2S34YW7f/626lmd7dIctplt5xqIwSk3B8VJSGWfSWQd
U7DFUciyKel9u0fy8i7LQs/MIvDaH2buULLQ33G57TlPfHxA/3mgdKkkaSKILwcb
yWoRRGTeU91n+UxCikR/8EtOYrXQYqENHsFMs9dY6KFnSGOrmMBfDXkZ4zA044XY
ERul44YonuwVSTbXSHkIvJ22ptYkUF/VXSGEV9T8QgaaUQnLSWcHqreLeXTCIHU4
lSbinLb/pQWpljgE6OnER0ZLbyhiTvqOSph99jg1dc+FkwqiNJtvWvxLKop0pyYI
rs2DxgWlwQohpE6TWPot9Jj2zDFyWF0sancWQcW1AnAXM4x6dV4jzidaA7MeNxSi
dCo5rt+SInTd0YRpS2PyboHxZ0fgUFqRL5O+EP45fiLOI2ZRgJnDIJUHVtiGX3UD
C5W1lSdAYg8/EcHxSChNIdbT5YvwiaxEWg5zKoRcET/WDo3ehjLPK4UccAgG3aGP
tcDHd3ztjZ4Saw1TiarPbDpVN7MwXtHD/gA/kYHK397kRN7gDJk2gMX61WeUlKUY
4YSLU0rsoHlFK257KRp2mtxvTpMY/43V2LnbsNv5+Sk=
`protect END_PROTECTED
