`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UTqoAgCQil55QDdJJEe7kJwmEbTvlrePG5e+bmFGOOhzVY3WdBzNl2aqVK0uFLKu
4eA+2B+oli9N+8c5y6HQC1LLyyM2zPcFwQ1CK9t7IrIzNNPwOmGouBNiq1f3OVUJ
gIiuTIClnaf+Qe/qufkZ9+B9e5ckZeTaF/Ri7glrFSoqMVGsmdgNQA1LZiFEhFut
ZFdIwpesdUJthXHbABwgbdyjb2oJB/hoViKp7ToMng3QO/qCFis3BtMeqURzlUtu
ltorY9vPk6xMHRNkxw/RbSlT7fgBb+LeZ56yfxCrBMGlusJElhlP53H/IJQkrIfk
LO/YS5A0Xj3InZHcPS+FdaiQxk5fykkbnA/P6QPfad43viUy2wVI5XFJZufFR+Vj
8DBsSqgNv+DBCMr5++t2qxKcW8fIJ5HZ4g2r0t/BWio=
`protect END_PROTECTED
