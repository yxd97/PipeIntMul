`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wc4O/IPgRmflbtCNp/EGd0xj35LEBL62A6HwVrnwWnXbgE/L+HdOoml1RNR83rbI
8ujC9LHhYEWNp3FxMOmi5W8ZfFKfWTH9sqS9SPp/2Cd+lTwGTdWUVJOF7QVcNUnQ
c7N4ngs0l1bDvmGUcCSGK88VEvJa/g5TjBmJ9s48AL63kO/a6b9bsCMEbwvhOpv7
oEG+HGQKRaPurv8D8nRA8V5k2Pa4bk4uJDrX9MbYPBID8CcP/RBbuWkcAvu+uQ1Z
rboo0K4K8oHjPH5UhK6APCS5Mk1phDjZv0ma6UFfTRXkfQSZcN3gnaMZgE2F9ONL
`protect END_PROTECTED
