`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPf3ucYG8fs2gRnccU3HJNs03PGgXpF0Su4CsVyaUM/cLUQmK2E63WfEwmEDKJMF
G1msmin4mUMkv2gWbA2LfmV4AU2IetB8aqWPf4mwFxkjZDQ93mb+44pWlTR7z6Xc
2z7Shwmgt/E2bbSDglhHjqfo59wP3Gai4j0p2Z8nsmcPOjrxl8a3/wlSb6/cVNIr
dZilGx5IdIPqxgf+DO3YSOo4u5cTuUx3X4TrdaczpIHQW3/yDMwdR5LqG6ev5D9C
YAE44YM356rpXlFeKlDuKDm7ZUPgAphJIkR0H5OSKSJ/N8Dlyq5R8zA69O6XYleJ
RiBzR6oeHLddol3H282f3nd2uAImjdfw0ZpRlzoFeTyR+fDNwH/mvV1RdfXj7fKh
XK2mEnRxkCd5fZSrSRuXOr14xDxn7HHzbmgtu74wGMUxsMNTbX6V9ke0w+74rhwW
fpsKBLA0U11IIbpX0N1F44LQi5LPBBn6z1J/greCKYYirV0dfwmao1kGWL/8vtDr
ZY8/TOzlcmJAWQPtmssl9goyumWU6i9zN7WiMvi6p0JrWzDEzacGdo9bBBxK5XHv
3GAek0RFTuPXNCIhsubcD675mBt/+gPCB3rL/c8CE7qELlXxrM++hzWhAVA+ou4I
iYEGpc6OueCjMvm20cUUmJJhyEcNTu1/GRvoX268JYaVkWzPlck6rrXPfc9OY29P
kKooqngf2f1n8vuy7cHYzBEgtuOn/CIzPOipVN/ahJLkHGkrM5LcubMgppFbBUL8
3AlDp9cK+jTyTVGIZcGb3xPYFJONtRWkAd/P9wNlqbQbWK7nB8AZJqP9n/5OgAGV
WjA8fM+/XqefIhcfJgvw+VUhgehs8gtys1jrHIl6xpjLwRE7ot/NlNfCTqknOOmM
TBG1Alk0QJPWesGa/s7GkrJFngJLRjxr7QL3VJtKD+JvNLGwzrQHWGQuRSTzt0fG
ImXS9BIyTcUVSSHfXClMZqBPp3Pfiq14qY6KO8we6vve8KVadMr5AqRhJx4jVB72
zO9C1MUuLlTdQwKG2uvs6JLCQgDQnV5s41FFUT3WV+E6UfuyrcQBZR0sUqMVj5wU
m6xma0PRyIQOjRDBI5yIIl+OLT4KAjCYzK7yNHUDSRhBX6jbqaAKW+XF+F8XUM5q
6HuZhwOghvyaqce2ATPMkElhSwIxSQuad3f+O0zpkCZLt+NU73r75swV6tHz7Kc1
WdaAVu75A+irnHsBGSCqn+9d+aLRw5AgU8vkWsTYh999xHRObEG54icGLxiXdDxt
v5yTCsmIlnc1Hoh63rMWnPmoSVvRUWP+fskuV/MDaIS7ppibPBmE+hlVmS20AiIr
8R/W9zG0DXcrWr3PIaMQMhX4yiXoN5d1kR8cGnFl9Ije0/pte3UR7HzXofyXF5g6
mfdMpEDU+Q8zOggbPFidNqKW63nt6trr8iCdFaI/RR/SMUwMIaozm/oaYFw1ICey
oXPlu7oQUFyixEjcgaGFSMTWquvxkRobqVlLOuippu8/sQyfMqBRji46i1R9rc83
abn+lQW6uSI385V/iHRn0+1Uzw6YbTUXC41jM0OnGecZzpVAg4KC/E/z7aNZmsN2
jIFozBVUjaCodWAA6pwzwEKAwiNUc6nLBTM/w2oX73AxKvHBq56Kwoh4HW5GRNDL
wRI/0Uewr1fWxV1Hk6Tl69q/ubqszYvMXvuZt58EoIvj5l7A7b5Gcjfr2L41Yx6S
ZuL2VaUsag5/6Oc08yOKF4x94qEJ8vj3EdkO7njFfI1iQWa83lCKhkSBUtSslfNs
NOnfYhBDOdW4rN0omRPjWl68HUHOYcnt3S8xQ9jU//AmVHk2OTYh1164i8Sn6eYP
lOWAwjnZASpe9Q70aj/XbZSDMBwrqA2jxaLriMqqPYjCLbThguDMFQql9qzjOLRc
BNg/X0U7oRHJ6DgvW1m+qvnjepNYB3L4SgnUz7QzdBR53NKqyoYic1hMq4w0jauO
WzKUmOOUKVb+tbfO1c603LlwsVmh/+KLlBHPtBH59XdxG08TtlkJ8ywYZyKI1kyA
nD9aFPUkxOAqHZE94SlHx93fNvbGariXcXz69xlpdK170gxXcRx3Sesk1lo6qhC+
3Rb9pk4BFN1WxgIMSnO7tli62xQ1C5l8RkCnFn75UIY=
`protect END_PROTECTED
