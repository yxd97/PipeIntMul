`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a2rRInN7infzyX40trrbAqJzYqYb4BgsiLNGjEiXvYrLQFC83M8jyTNKshXIsuB8
UWkCIbgjsUBM5/m1fVrSvxGxqeUoVbLXeSuHjJ+JzsofNkTl8GdIGHlLQ+li7Tks
72o5NpbCU0gqm668Qjgr1Y9sRmpjEftjrZI3ON0D7lTdhLAZqbcZ31OPnG6TWo74
YYYmWT3+TzfOfubrd9KIh4gQIx1fkpByhIBKk51L9lTF/mPEnyOMLBs06V2eWOS1
qWv4XstTqTi4cy2xmNf/7vMD3ewr55yhzJAplGwn0mgQhPqtpQUq9jlgaIXXLoSP
RCfWSqj4fs8cpDZYNRuQ3eaCawmt2tlxTLcRuwSodYzyxwhRhis+3lj6r98zFQMA
RDtWr45/adIPALcSKtlEmwaIq+IWliPL76SZHytKd12xqzLkJSIfIcutSjN8Elpb
`protect END_PROTECTED
