`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTmCsD58+XEd+3BkoBQifDh66YsKWNKFwg8efCAXKxgW7K7/DJ9ydmYVHEOBQBT6
E1/m1WAURbqV/0fOXQ0iWkCc9jPpMc8qq/iFYTnbzJf8hLoBdMIpHdL3oTLW2yWA
CqC4S1eGBoQ9shBd+8h2rzkw9JgC2X3ELHWTyH5IT6Rm3vxrQTJdodJY+sE9AAvy
M1zUDe8y0jhDVjxtFo84S7tpq5R498C/tN9KVnGfsXC+adFijLPdLosLGleiE/W4
907L00DpHO4SizKaIv6sWWP3ZU6NR5Fi2J3GZ7jNC5AP+shvnLrzPw7gW0ESY8py
k57pBZlBM2aMIGiebo6ze7tiXIY2kqq58Diibadwq7V9JztX4bfTWy8/PvqaDHRT
917Oo4Gry2Th0+xqerJ98YShfLB9FwsYEKvJNqp88Sd+6eX+vLdEOs8xyMg9x7pc
1pprtWdAl9b1ejI79UEL642X64HzRGXjuPKqaSLGsWh3KCdHZvr1wqgG+uloIFN/
0YM3cxp7lKAC/n3i1wC7Rhv7yJ1Tq8gQ6W43vN+aKypNjWnoYf8zhzfUJ9j2FdoL
p155nJvcX1rmdOUcaqnKOYn7Gxll03RHettA8jb5nXqpP6bcwZSBY+i//8KfBd1A
8cJCemJ2NUO96rf5/kogOj18nOsLkSm5nlL1f6SHBpCa/CVUKsI97GAQVqVO7rpn
`protect END_PROTECTED
