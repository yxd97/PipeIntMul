`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iUMuNhoVBzXiWqphqYj0+4vzf3FWQJs5PPBEN7WAh5Gpw3sJlekbupcCctYI88dG
9XXzhIxW3a8ZQA6R52DRb9mQmjV70jGt7cx1SPOAAEXmSMtkTHM5a0guhbJRMXtQ
szMrB+1HnUEB0Q+Fpy5AIpaYzCOMwfclUCj6d2Gsciww8ah5rdTfXCn1MBUadi02
KbMi3NQdRpjK8bZxxs7R2Wtz5dcSBKqgLSYi2JgCSjcPFJND/j/dhiSKvyXIM6ia
1X5dxClgBn+P4ARLGKbEHtYQYldyaWS14exezqm8TjxECKnu46CXUSjX5UhTuDY1
LHgR16a50P9QDxiaxKSRvg==
`protect END_PROTECTED
