`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfwyLjik5y5SrjMdoZMTxVTCjGuA4H8wSf3vdlm/9zEd/1BD4ji0UpqDkeeqY121
N1guIUQ/IvniMmkIVZUveIhyKUws3BqphkhfnimttJNNdaoQ6+Owkkxl/yFfC/Ak
aGuIai+851HMyIqCu2os/SPb7WFfFwGmZsg7OIpzMc+a6cxJZCI6bWg01M6k5itu
zq7JHDzA2SPr3/OGDz1U/eek5g3oc/TO6GfwnX6XtoXt9jfyQHtjxMH+oaHlIBv0
vetA1QHEubImFMKY7FYT9IR7dT3Jq5hDrB0rKcAou41NDP7GeSUpfV1ag0pH2D1G
EOG/nmB7tMwYjDc5LZ8FXnINifrGKo9utgQjKU5PC6BY6x0lpTh78Wf5/Gl4p2k5
etvtwh3ZUofigNfp8QhH1qF9q4k6RsWOaAhSuCaL2XwTVoDKN2yv0fZswZAx28BU
Pfq+NnyX0Xb0FQ5O9VYNTcqwWSzy8heT5ggFTaSoQLacjd0X0XQ4stIsCrPeEr6f
KNPh8M1zIoaRp/oaqjHdPPe3TXO+wrrmAXESzdXMURuC+lb58VYh1lhoExqslXtH
NDZRlb0b+mtp6zYTFq3WokQsGp2hFgWrZabGmFeBtkMZTTx4qBajoJko/tpmqBba
5a0HzGpG59UQoIlGWwOAgZdiDDFaqer+5Tty9DfH2tnjaYvDcuTSAe2/rAQ7Ehus
2aBsFVslep+s4pa/dfZV8PrY0oJ/i7MlGoJ269kf6a7vBo5R1qaIHtzOX2GKbwyx
bSqSTk6tm+g+LYPUDgARqHCKiWrJWoKV8KucnvKqJzPic1o4eQ2xu8uYt6ro3/YV
jTJQuvgej7bgKIvNWQdIwZeCUDB4uU+wW3ZzvAKTsYkkzcBenPl3MN6JPT8Cs0CG
II2A3pLxPIue+6d2ACH8xHlqiavn2RbfpnJNSzw44VPkw8wEk5VLlynHeTw9sHzg
8KU1Cpxg/nWF/fnqCMuyV6PNtRDDnfBDqKZLpeCvTx8XHf0ee96OfMMd2H6Z7Cw1
fzZ+RWyBZa2IRSoVJqodsumIDCIkmhataXXZRq8NLymL0M29byr73ZSyia9KKfzq
hP9F1nOXptukYKU8piwN+ZRAmkvHTNz2UqVouAgXpaWe67HzX9C2AjShCryh7mjU
mx1An/ry+BO7oHAU+d6EE0tbcjy6tQWYrlSuMz8MGTpu3KFMqXJV7hekJa1sQDEf
Mcd5dyfDLC09U/2UPWM0bWE1fgzSEQaFzyt7t8gavG1d87uJ6Mj9YNTrHfROCAfH
mt6nZ5vKLwnqEE7fQztMi9Qe4ubMECDrFJPy6vZczVzEfMgVqiOIt3cRgAP2YNsQ
XymQiyrtCBiGPR1qwSCAq9c4BDbnfOEszufWv8HG7I3NS+FLinue3wQq+FDs3Yfb
zj4KsJWRutmcx5P1V0KIzA==
`protect END_PROTECTED
