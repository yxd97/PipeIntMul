`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Won8Slh7uiT1eCuYBrRq2Lyp0L0nGJ/nzIc9ysZcmAA6D1r/EzDE4CwQ6po3HSMC
uT+Zf9gpoGn7eLE9TfTA44c22hTJY8VHh16zhI9EvicuFihBKbEsplnD/Ajqzefh
25yDmafEn6BX1U25Qx121XbmM7n+n+GYAYTWBS7xW25/HEb46XM6fqjwJiyBKmKg
jUnlJppzGWZyDcS59pQbrJJaw3NZQEINGUWNIGPKep20+5ER+bUUkggJQrCXa6JX
C0Ov9zc1FbZ3G4JOR+cNyO5hyqiV6vnXYRwMNuSKKpKTbQz6RbVJ6JdOL1yrxY6F
2TBVH+dKQVqjRs8LJfMIPLvePz9CwlJZDdSEhcN7iJaZMXMWhru1SRmo2AwSJkd8
eIDL3elHnrHYBdlGk7lXwhPa/5MEmfgh4ZZ22UQEYZTsP7ekMHRx4a1EJQxyeaqU
jsfUZYCJeb+WSm/HIz66MeT750Vweta7SMyRvNCnqcqhzqMQa5mjOaBIwwlAJG/c
`protect END_PROTECTED
