`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+cG5fzAIj36sNEVNAK828+xdfH5o1HM7d3DkUyVlY/YQQpsW2oHC7S4BEbEDuzZs
CrEq2jhIl8GJuMaK4lQGH7WxqSwh2/QS9G7DRE9yE+qTCDn8GCK0T3t5ZmUjuIJY
sKW0u7qlHa9EO9sfdFGjIsCk2k0vG6RXYUK1zWYtwoAgNaIWDu3mBCT52zT86GUz
hq5X7IRFXtGYvxkX7DNjmChuyrA7XW+jo0Tmy4WVRKu0MKtxROT9JyZ0zKIQFPVB
aQOYySFra8ZPFyoG7yNF4/Lq6LEsOfcfT7603OiphbMtUqPT8XwwBky2TSanwQSE
OmF08h0NTcH5ttLhhTlV3gsaHXNNal/wwMr9A1LWwYEqWubQ8YkoZS5OTbrR0LKx
8bv9IjN20obO1PfajMGSUE1d3+Bpv/aTmpvD3CwEJTLxg/Zcp1pi9m5XhtRcZW9a
HF48zJmjDTvEuLfAhTg1ZfrndejULcACzYm/4aTXQB5j695x5gIZ5tQ1JzTMHdW6
8J+FSz1n9EHp1hDL7uqYK+GO1pviVak2++U1Udjj1VsHdgD02cRhUBoBsRWP/jP/
nI7b3jl5jeWrtNkm3d8197AzJywojZg+6CNFmx4nl8FJxJYZ3N6S/NlCJnjxE8zW
v/mT7b3UTzqSp+0vOyNOgCbpQXLwOSs0/mEfV1m9jzJqlYlzVJdHRt80TdzUz5qS
46LsWtgpd3795IE0iTpPprYxxJgEiQ+ODumgEBoI4eoe7+k5Qvmm/Tzx7f3+nZEH
q+HDXtlH0owU6agTuW12rMX8ILGoMYJ2/oXPdr3D31L9ptpx5xsFfhY6cb/WoN71
9Nd+EG+EXvGjFWW1X9W3Ug==
`protect END_PROTECTED
