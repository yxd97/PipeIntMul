`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1V48qbH6AxpCxg7rd7Xs3vztu5YEv8reQkkQZqof/1KBw/CFWnn1cYgWv8M08aqz
0H/u8e3tJMB0lxF080b7/sn8Uz4wWMYzpqZF8pRlCYv6f348/fNLdZyyJLvtkL+a
9pESogfDnnSzN+sI5exedhx/zD/bBSEdEWxJZFmnj4dVsMO99htfkSbPBwC3iUSL
DT9AGQ33wHccqgNS3feJ5j+JbTI6y2kbNr2IKemqlbJA2GjsPfF/RnXgImRrZpdt
Cn6vHUiZfJRCWTyvTjZP6P+CbCm8YWsNmuou+PkCHdI=
`protect END_PROTECTED
