`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HS6FXf04wDBGU/KfsAL6F6A73kCT2r+HlSIFT+ukS/oqUr++JSRLyXEUPiKIQ0iG
phieKU4N+A8KL3bObdj/Jn79zSrXyVURDvhMBppCBubwoygV2b68L3W8OwOUxR5v
MegStXMCrvTu8scgIFNfb/r71AIX/RtKdNjxPcCNRDdK1X+7Vg/uggUWaftg2WcS
p1n++IaMgI3vpaJz6jHuyrwqvG1wrx318SkMqox6mVfgx1cnxH+2d94nGuyMbGNi
+NlSxWd9PvoNMUk6ZwffzJ9e+Kqu1XRcRmeMlsj3BVAK4hHr8/8GyZKADTHURIsL
xfVHWtt+uLPU+6aEwvFGe1sr84WdW91yfvBkTSF4QBwAshA83w2SGoQP61+IOzkZ
QQWgK9yBR41sC4dZc8+EcQ==
`protect END_PROTECTED
