`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6xiQd3sJ+E1+HZfv5v5ms7o9IkrYY05L7uhM5kWXuSa7d/Csh20IZkei58es9IH
69xP0P/utD/ypfkuCsi2+Ggy+d/m8Wn3XktIGyqLNcNswA9FPni4jVMulY2ipsHt
s/w9xp+MsAvGkUTFJfuonaZdwg0XFvkPNZk/YrKys9NYnwqakNkercK4FXS8mlKn
njh9zUEsru8fOZCgTqChV7x8mZr2bLPQ+ccssdR8nv/yL5PEgVN/SmYt8T8VMhts
qOcyh5wzRugkAhxZ4i48TYl7k9YQtg+dDqQk35rccIVzR0ZcPclgqGlW6YIMiT6Z
y+qA5yIpyynnN1WX0vc/sSYQuiP//TnY7c1hAnCV9mY5Gzzkff/Bc9IIjkczk417
FWcXzJgDSB/PQl3zckx2HIe/1ETZ6DDUiISRM1t5nkkec9h0RG1MidJz+o27vhF4
Um7J27Aonxexcf+0vJ6xv3x5wi3voAFXLY48nUAlqTAXr76vK69Svp2dcvPyZj39
PCErLytMUfOMI/l4JJNK1Cq86ZSyxqx0our37gcT5Gzb2pIgWCJgrvMRU+l79IXL
asx6SOzDYDG7FUfThqilSDROLjerMyWu0MoRYiJiSEnhhp1S3JF/itPkiV6nx2Qy
4LT0laJw1zkNhJfR9EoNCUNHvql0I1a/L/mix107eSYHf3Zlc60KvDsNetASfdRV
QUlE5agxjDQx39raA+anl+CXUiVCjuhm1eZio8TAXUz0vbwqUk45lJohTaZ1GvON
QUtGu0lI3VXDnNerECzqBqi5MB4buQ455Z2PsYx96nfk+sjcgW4HJ65lOp1Fv54P
Ho/XPrqx1SqbJNYMSsjHpwFzvNcjIwiNbYWA4YgrU8n7RkRmBY30zR5Ojpjhnvrt
ZFHgAk3zXtZ1PIkltXlgQBYUlYiWY34vFS9LTiyCUIKPwdeAqn2ixnaqbe9T4GMW
3gwayxbu50TC56UW4Pi5otBCJJ5E/IbzfCIqI78Xsb8qAE5mQ57/k4DSADB0Q+bp
RB5cCvuTiy5N//5XTPLQXA==
`protect END_PROTECTED
