`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JTq03ejNUqIQO9Y1qvKvJUgioaMk/0d8ttXpju5tsbynJZdYt1HO086UK1JGRQYu
drLRmT7sRbGOy3nxRHDjGWcNXUBLFXj5a+m4aeJgO6mi51OFYnnNQUzhZMRSmIw9
0eHL2Uw8o42nT7uSlRadr4ldZu8luY+O/hJjAGxul1w+FBOh9UhD75ICyoRoCGNe
VxQURhJSyFime9eoCHSfI+bbuQLmjhQQJvtbkLb126VtcXwxBlJCLhWCKSVKcly6
MrUH/8Yz+t5Spnmfn7RGz/IUcoOSBrcv8b49GyYaBoQVf2QdnwLe5fCVfPGTcKLc
99kgMjRd38nh4uj8AzP+adv2Lz4dQFPUMU7dVCQ6EtctjXJGakGaeFevgOR9+X+8
XKs/dGthmfF2cSH3pIcSOesrY36jBp2vSUXqSpSoAwSBIiRIKlPrjS92SoqZxa4M
zAtF3Iy+dxB/Aj91xq8eKNhkDniKbsAuBhqE+PFqCh3V+4JifTRnP2YdeElrD8K9
Yiu/wKfFTP1H3Pk18DPuUyMKcRwm49IJpDky8c2vBaiqQBbgehTSu4wbcXDNymoc
BKWJ2xenIYhZy/sE3aQNnenrKEQUkfejJ03mzdUvGY2fvkWq+3xcbcIDfaL3ny8s
XMpU3LyI8Xq9Kqz21EeihO4/HpndYppdgYSYkQN++NAgah5mMujzYm6gx/10rAO2
FjVm1ee6kpmZXFi1swfiRkI+lFfQsKrs5aOYi6BS0W0=
`protect END_PROTECTED
