`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PTpjJpsJLQtSuhPHW5m2lfMVhHpb9f2wZ5HS3bC+eJFIquQaYcnRTmQz3JHb6jm
i+9B3cjQYLABuXoifTgjMHfyMXBdyGgRZjebrCyqIk99VhOjZQde6OxNIwr5sgNR
h6L7h7JLBtacRVdjSNmt6/GC/hlriRf+ZAXCDvhQLVQxPu71J1/Z+6MurtNtS1DN
1lPg3tW5sKjsPVy31WVjOFallNSejhOL/ZLSi8cnYV9SdCfABkXOKjgUL6BXX25K
HGFWvkmrrJZ0ZM8MOZySAg0WQuy9gXAPb8ScYCoReUwl4nEKB5NIxMgGbA9eTGmo
`protect END_PROTECTED
