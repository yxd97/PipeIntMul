`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBKan8CUk4Ws/qG4X5KR80ilFpybIQqLxROEElNWQlzA7/HPKRwaLZWGQxKtruNR
FWffVaCHuaNtkCDW9L4yFiAe1UJJUOF4Q0vsgehEFoX6BlKbaSGAs1/4ZpeaJgfg
vdMobuP3m2uQ1szJMOAqLCXQkLfdcWpoMrAieS3lZg9165fGw7R0kMWIBNJ1uMSu
1POLvC1+gkXeHHlfuYG2r7wOOa7E3712UqJven7RPts6ZLQ/pON47ZihsVEbU578
uc9aEhy0vuCopoVaJKChb0cTturcS5vm5SoCC6mL5E4nAP3ulhbulkJikY0IqDWG
ckKtLAKDMQnSNDmEkGx+3anAHfolIrjUQySTL6EeoCivfn36i2B7QgSA9dlV5qAk
2NYiBSAXvyaE+N6/DrmoesRapBZh0k/mxZ3PqJyI81hWznFyzeYFwAAwzTYXUL11
K4i4Mpghx64bKbozImXwC2yxqcEFV21uS6gf+hguhFqLBml+1JvA8aIa0CtVef3u
`protect END_PROTECTED
