`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1+lvlMjQ2uTsegWhnNQDW6jFFzM6OzfZG6tMdUD8FPAlUkM4TEymDbZQdL4ZeWq
qU+Li/Grwm2e6yQPrdiY1WdTHYbjg+Z6aVw6Unj3LB+faJ269BPNABBvlUbSaBgZ
rr14xyY2O0U9lLoGy/mlDFWIe51P+nfJaTwxi6NjWSKm9HmsMzzguNAP9pNi7U6e
OUZ99syBzZFCpS4hmolbOaVGJmXPMXc1YW3Q6nmXQKbtvL85jBc0IblBt2Q7XHba
zblrv8aaoWRMFpncpuVhGqEPozRmPEHuKDZovR+TJwrZmlcdzSA+ELi6JS9IhtvP
6bvRGTurPtMYjngG2P0ypIVGpJ2gQZyWh7gIKOyr3SNZwQdNyK7zVm0WEcxbcbt6
grPHaoiYq40pDr3qmaVcXazLc6fNkIsfmnr30w3x0/rSdw6ZoNhPI5xn7PUXIz91
phrc4kgLWfheHCWzrJvvqdKdi5JcrCvtToZ2R78lTNmGIUZL2I4XVE8TxUpneBHB
1evOqXOgIfgXail76ADA57ETpUomt3dPp8DAuccEWAsCS4O40m8DJfDtpaTwNklV
bpaLyV30wxhfL1HCtNjvDrhaQ9Q42+sesHGuhK05kv/J6oXkGcihyDJuysW7vxpr
FYAogkh5n5Gk2h10aHGcpHsx9BKPdBnAm6uYSJ/m7Zaxk7yLf8HI6RGRi5YzGWOX
irEuvaHFv5Gu7qGP3qeriuUhl4yrtJApsblaNKpuXpMRUNrLjMIfnNIRTqrSSlI4
nHaHZx9QocyDxo+4eyJf1rjOscLNWewGPmro2TViik5DUW8c27z4iSxaPR2UqL16
/RkYvWFZCDsj/etFGnAnFMPLeCp2kiG5qYEomHQRndkmyRWOdxRbuydplJH6AQE0
SEfHhsXGffKPZpLMJ1cU+t7zvyK4CmlXAohNusjA7dSTIpZpPEgVhULfvWe/QBi5
pEhMoYoEoRmKk4pr1Xv1cJ+XXXwrKyB8pYVJb3TWZXx/9Kegd4vNDBAlZ2MdPw5V
djM+y8MTqaKNN8vEqXOI8sN0hUpKvPMqxqhJG9BpBXvSrxQAnU/GkVxHZAfAzqJT
/CDGLw5mwaUU3U6SvFnq9jEbpeNMEWZ5IrWnXcaUd5dY1iLTGj5dBX73B8p9BP1k
YMeZqQALCvSJONSMNE1Xg50wJKV/NRFjU9DCMztHy7j9uSaZd61kFQoXMmH3xWdR
NQ7U+F3HKKtqw9bIwUrDQ+khPAmkWYefru/EBySOS+9jPT/r8O4G5lA4uCSSQ9Cx
95bSTM/6jW7hLompbYAWsS2aR88THqkTcxuinC0o23oX5iv2BK48Xr+vxlrwISko
1Jpg54DwQb/ZCcBMcSDPuWvhaPILKPybmNl0DHolrcc9SnPsvcGg7xAcad/au+K6
hngpA3ODcdXvFrC72qSmngIwt+jfPv7/jknixR+RhnuNMROUByWzg+r87O8yR+6g
YreMxqBJj9djEdcnYRIX2TtJrhEbnqMd2fNTUX8IiuBTP8JJjUHuA+sSkXESgLOG
nhA8lWrbqCQnAK1b8/xGFlGAXSARneMtBUiRV/CxGrBQyAjoiRzPatAShI8pEdrR
Zk2fS7nha6iJAiTp6TswRhua7VJmdXEivOzg9mFy9y+or6HJxGSeNmrsuGaJmXm5
nx/ceoer+gUq3nmLVP/y9+q4VVJkv1TPjaMxG9T6wd/dneJJNf2flDSf2vUmUSjI
sKigmnzkgCmeyXTEmH/EUKlOrdC/lfdp1qSvhpKpx/C9KMd+4vkH85WZ6QL8OKYv
ZW+Hb14Pr4AkEFkDZAidB1TAlMEjT7oz9FREsUE2aHqvwvft07+g9BbmFGOvXxA8
Ju6rCXtYxDHBGpfiS8xVUVHzH8hGJS7z7DdHCHF0xaymGypTGFBqeUZYwlZiXzpS
bK8QTEIEic1UUHrUWgDoMFTrxO/Mqw7McucXhtnhAachub1TjEiisKPaEMamaSsB
fPNIhJ4n9EBQrCPITOZO3NQzzzm6I1Ip5XXW2pRE16hATmBviIWwO3RXMoQm+uaS
bFjme+ALR5T/hxZ+lS30MU0DKGho/FKEzIxcqvzNRODZwwIo+8QHWZ/31Ib4Kndx
IQsUdwzlrzGfPRe1k3kQWCaIjguoL5NuSe1572z9Ut75h1Q5h0kWyFN+VJHjwVHE
uD5VzR9Zem2TAm93BR+m4q4suCREohegFJlVAqu0vJfLD/wZ9WaPPLC4tiIl093k
6rTOj9iNTRjFQVfxQQu66WPBAAml5gdlD3pqKswO6dBnX8mlz+Op0cnZHWSeS1sv
OAGhCH3rXD3cyN5WdXazMtdczjQ4JPAM+VoNgF2Fo2zD7d3vJDcrUrDaX9lg83+S
AUa4hgD4nSYaQf/3UP2j91SLvMYi26FhstsHC1u07vtJ3rltI47NBecqcar4Q7VN
8UChXK5AGHwk5d6wTXvh+x2DfiE9TRvoCe99Yoes/XCRT3krytNLmAYXdVoaaBel
wKwqdKm9P1qyvVAtENFBbeN/6jKdyZyuO0h0gBWlJ7DTpwlR5nspB4S43Q+cVdS/
fwAMGLkRjHLPajYkxUUS86puuj0CirThT4hVUW6FPQbTee4feW5/hiMdopP54sHk
Iac0NXn5nfpwDg+zxREF90PTwsygujrm9rJnqrgIpxOFrzem+bgnn+rK5E0wbYfL
R6xcvIAAMI9VBBVlQ33lbJTiF2o/sRmqTquehk+YQoHvMGCdGooBNa+24xmAz21P
5aFnp6UDDu4OS2oyQPJCe/DzJR3qxrWWyXMll39o8yW/9/KBSmURmvALVX8iNnJo
M1qkcgR1dkCFKO8yqAT9WxTTLcX0TgYv8yx/lUw2axaK5r7a8Zo+65NLCZRjjXTX
onuVTL4wZN4iuuesf/Kc9GNDKjFxD2WxLJx9VwLywFd6gmZV44StHNWhu1Upg8a2
sOeMiJ9HseYWmrgxjs41ctvbWRibaX8ygCCzgObYtOQYVeXLn/D1MQ8S8gf2vaK1
`protect END_PROTECTED
