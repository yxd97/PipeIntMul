`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSDrb3zWBwL9ljiHAo/HdW/N2NAE/3BtUrpybHNozmItG8H6PHdJ+IZ9lhb9LtPe
CMq6L5kL4/8c/kbmmFa7xnRkDqL6EAPbKMRdS57W9PauH7Ph7Y1OoW9BbyCPnSYs
FBfpQkwlemHjTE4w/L8Gwz9es8dfUo4LXK0HKyj7ZW2D1zSwqy0GamjZNeZPth8j
LgSsUt8So6UUp7ErttwqS40Jtsv94D1BVG1L6foFJBfi9djzCPAcinaZCmBOcXOH
YBqqoc9oEC+8jP1EPYWuP/jGIYSd/KW+R+naTXm3cKBHKoz9uBeD1RkX3btWhgBN
gV7slKzDUzAJ+RGrsCkY7gxHVMSiILfidfd1CYzia/NEyq6dFKlidf7irkIFtDex
zmpzvUDGkEeByFm8ucQ8Mdd1O8g4mO98RDwMhC7VFdBTAqA21tsc0QQYPbExK6LV
x/FiIc3dCXN8Avk6MTiEZCYZ97wWTYdPt4+920WpjfFABoN9ooJCoFl/10DqAyjL
OCO9OBvqUVEvHA1bYPqOIDDkQdEftlUQzbde6+Ncom4exwcIUSlm7ccRvMmX+zXZ
lGz5rk19XM+G3j7e4FIqCC8AKDeJ8hpGd1OJtPmiQtwgK1yMO6u34pHXlNCZDDTS
oygPLzTozjRMKSLBTxAbRbRGdLz2duRhUSI4V9EOvt8gbuZ2EA1jKtamH3rD8tr0
uG7+1Kf3XiyHjNP4TodS13aI+WPylEd148J/TEeJXBSEGWjC8FMq3sryfN1xgpOR
Os6Rd2/4W9NC8VcQClgt/iRehx7IAVHMf5hCWVN0FE/oBoolHMPQW+yCMMHMo2t7
7juvXGqzwRcowSl9kBQr0OzAtcKmiZLy4URt97B9/+dOlBOOrYRjC25v4A0/BCPE
YI8rR49RDi6bW/HmmVapTWk/kpBeosPM3mmTqjON4DJCc4nqY/umqd0ocKjgpQer
TzYZcZA1Tl5Ix/L9rgkaAm2c8/DPzBjJJ8UBq0UkEtp0U5LmSH1HWDHPf3JRLebo
aW+Q4kwdqG96Daon1parWq/hIOt9qbWaVknUjk9saaNWMgW3g88JMcqPcWdkE3FG
5GaFHi89MWelIpgSqe3Kg8HysVWF0u6JdwI2xle77sfvRyhM7QYKZPp/bTPDuRsy
DPO1CVJK9RS0m0yPGNUGdx12JDbTbEMlyMMc8/JlxgIA7l1PofIDDuxMiaOX+RFT
/X6XxZ8/Df8PKmpZmWGtrbOfntVunMowmndR46aluKnYHMNyBvDSiIyxIEQg2Jac
srXhUOC0UqOy575UzxH117SkAB7DTRQP3CFwg5IUQFvEbXny+h3tB+6hiSip+tR9
D6p+6E7PavUatv0WS8MqEqCDTkUSAN/NSNenYD2Lq9TlW+ubzKvFvrPnm+tjekXZ
DW4+Pl+usO4CMn6RDgUy5Gq6VPSkNxreVxHvFa7lT4n2ypFMam8W5mc6QGX2z6cG
bkos2nuW4H9gfEVkuigOIiSLX2sQwcEHhznpDR4z0qp1YuNqiJlQO39LGtFUGVlv
N4e/6Kclygj7B1gvNPr6K6r6dy48+Ni5ipiW2R/VUd7kFTaRdQzopzeIBiXXK/He
r2MEx+gw2ICiJwkuHWP1DhDRUz5JmxgUfnQ/6C12Eo+CMbbnV+LbCo7pqZQYfADi
3DMfaov1kfdOm6/LXH9so5f2qzo0qyyiCTq3c3Refw8PPggyivFvuaWfepvaD3Yp
ARnjgAA+b6/H4KM7I8YCdqzGeM/v1u5Z21mfbJpHFp4NCHC8POp8UgHgB6M93MdY
cb6Hc2Fb2sQp8i9zUUqg3CeQljwHgga0Ni+0IX2OGh+feg+C55uQ9hs8ogOyw9EV
i/ijUYLpo9SzDS65Nl/JSwiSXavQoehypgpoiiXylDN43uhSKVRhorkzXSklL+YR
YcASHZw3YjaZd3KwkR3GGpnMaNEzqsIRKqVExrQvYCeQou8HmX86xlv9DjzCzqlT
XMAutwSEZmSolBZRAzE5D6gOen6WdbtQMKL3JWuagD1lxFUTdjhT2QVt4gX3/+7k
8VarQFiPRVQ2vl64WB7m1Ih6r/qmrKfvUcYFCV3mFSSb+ClaA30ZfDt6WSvDtG5i
VUsnmKQOFUau64OpbiUEAAigDg+5ftK0W2lXDWtDezfDF5dZSwhPv3ps6n4MJjdJ
YEgjLQUwUxm6DtoFDOPMTdHLX9aUWCXvXnYbIZP8xTIJm2YE7+Toc5Yt12Y1YccC
Qmo0TwU8wWgNdNm6OLGb7WkRU0KRj66J0wR78quwSHu4l+PGbNfuvTzewocqJB1E
pk5P7NksqU3J/rebsmlGtTEQjNWHIjPemxYLe/pi0E/Pjx+B0YBQKCGccKDCognI
ydSN70NEgHt7Q4Tdoro4IoC+TjX4ahb5O8Psf6ASIcFwI6oKXbtmb6dIKrevzInB
zDoNB71a/L+1/qxBodWGsm2deSGAAg80N2N1BvgzjsVDNuZ5JNXCd786Yw6xg3uL
UvXlG4M/tY2nlJPi3LX32GQhkaRAmeTWViZ7k5Q3AxdTwxqzxTM5o0/9C5XITo9H
R4Kt6thQgz13QJ9RZQ14rndgEoYQ9cOxE1NUUlWzqQJSPrp5YWpDTd/axXH+WYvB
ys9F9KHLLeavGiSoOH7jECBH3xR/hM5eH1anlU6sMC28kvmtxIM5b02Q90fHEk+W
PQ7JB6xtweV0MITGqOEGNft/ntqs9bC0FbgFTdQ8k+n4zab2fJvSqkUgmx92MDyo
nYtKF8biGTJ8H6smQ0mLdaJePMpVVy41eWxhbhha2KolTi9rRLbgUS5NDGREgMBP
GpJOtwWdMwRowxQddPaaQ+LmqYHcqOorBvJPgz8ZrByP+67V6WIyLHvieWd1nYJI
9ffYoc2QcIbFwsygDJyWQhK8fCiWrzLk6P0nzdqa8acAssMPHO6kron5gY/RgYOz
1sEfWGeNiDD6gMMzzO0Fq7E8tCJzVmznSTQxYK+G1Y/IbReT30i0S2Z3Dncys8T6
OE5awxTQbkJAvLTy+WA465YJ4sAAIixYOmGDRSCOTXX3PLVboJr+9J+jj4iL6LJr
K7wJzIerEbwSTtQWORUvW7iOBlDX8lzCPWY2QVh6Fs2KLDW1yUEj70fBb30i4Qb3
bQMfOL9VtEvov31mwHuplZsNqIe/O5xXmQzyuhjTUMK+apTmcGPQjZuYk9FfVs66
s8sFiM0YVMlSWOYzOuFIxp+NFqCtjEUvZDMHxDeAde5AOVMlBKo+nZhCvAwmu16Q
Gr3OwTgN6LuijatiQeGZHNlA6Qpia5wa9l+1ipePhmPqJlTlmj1W7dSUlHrSe82Y
r2ZHIf1etPjIoAYNz9xI5gN7ZL8iB4KtITlalZU48lO0dLmDHZ7NoF4V8A87+Jmj
6wKgY7YCaV7HpcSCBpX1g1fBhRbWbVifFL6HL4/n+NuTCNdQqnjSFsd2/gAcHafJ
YYPPLM2Xx129c9DMUeLT6nzKXIr7STU2pw43YVnnw6L7TMig7VbxSrXzfYT1Oobi
wRsF/Ij6e+ffg2p/Ev092CeQUw2qsTYVT8Un0z/KTfikAnR/nVx7xT8Olynj5hq+
EkSLbmYmZorThFXbxUmDWmnG97WwwsegjOCBtf9kHXlF5rCDyqkwx4KumcX5GPg6
RPF3ch8jxo1oUrAmSDBK1A54AluooqPDq7wBFbp3d54fzCpYPtfLwIMyOEJfLSG0
oX+wgNcq9wBfHlgHSSXbllRcLruzhCAaPj49+5UMaMj7incuoJtZWgir6IzUx4e2
w8QZMvl368x3KbDhg4v27MtNPdG6hz4D6JkNl/JUl2pBbVkNPa7RKt9NJbOj1CtI
4VdjtVVHz1040CC1IkC3214OXYc7Sfdd2fieGdjlgaldY/ysVjs2I0P9RvJcucHS
OZ/xl6Z+pMi8y17rMkRletk+8LY3zJZshyjMXV4wsmgxHhjjim9wqRDPAAbodQfG
75LX1iaa6UG2ajLmcO9iRQWxY1QuPFZIrNp1czWKT6m3ITZdVO/EG1BjboGpTBwb
WmLfE12QasATqLJuOsWeF1VupEIcv6R72TJ9rscpODbie1WFK54dtOhuSTRem+v2
UZZlLAvpPJYhbqJ6LYYUoe398YTs5Uv1BKeJEHNlgcUnEujmW+lnsvbDe1DQsWWm
eo65YmfhgcbXzSxcN4UkDH4zDAUBxAUwPNQD75t13M8ZoER30Su9+ezlls3i49i1
EHs/bWrZxJrOLwq8Ggzq2YEh7fq3CfOg38VxsAXK521E5KrmKDrUBjH+sY7fj3Fm
vBY7dq2Z/kl0OnM/hLQoISwRBIk9BD2WdZ06XGPdOtNXrSmPUoy5MpHJqVnLS/nH
l2QdeMCjt7wq/YtYbH8TDVK3UXDcKoxN6R2fQ4YL6EeQ3ZNikSF+4kPczICTU8r1
lE98JBxXsuF/LWUdIOYz6hP5o/IdL1EkqboBXl3VXMSsOUY4fTHRvwyyKkB4haP0
8sDDoTEaf/y9icedxcfhVKBTshV/bCOceUIaZHCIjq3Hx+fqn+Vo3/g9+yOFCoPP
0qU6tih3qqCeWQ7m9X7/QwsLEBxKXOgXL4wZLrmfPXTiv1ohspRl/j5O3ht/GjyJ
i0h3po1I+JxnttsGy9N3aHwOVpm7Y8dOI8/sEu7p8/dvADfyytQahrc2vqAgyFs+
P+mEQSGXf35nEWG65cKy652LLTwLNLo6/szy2FXWVpp2pAiyrW1K7Bgp1xUzARZb
+5mR5XsP4R1gpsd7MVz3d6THObrt531fDtPfddFmnU3UirT+MIYoa6yIABMalseI
GQKJ3gbXDpcVi9c6N+4HyMQY6pqRcYT5FBlh2A9TafDBKpFr/QnsTVLocubYHTt3
EDlainkWpYgbS01mDZOBZ+xG0Tl0LD+QZCfClNOfZo/EEuSgzLNJJhvv38/wO9z6
Z287jYJD28zrIaJbpUTqEiTh4M5h3tlo3EOizUjjanXiSbBdTi5qt0PYM7uh7leo
9gaWk29t7BiALBqzTxtMRS/7PR9ezCxz1CswXQVIIq7L+ZPMP2VFJviLzSiQ+Ytw
5bJScz1/ZAY/29ulB8UUCrNB/E3Q8PT9oi4dCdoOuoRwMC+G6F6Ixw9Bkm6y2LzV
0ejvtjTNu/WWmvhpjB3jx2f7FjK+MSTOuCFbwDCF517dm3jWfdvBh82qUly8y+Mx
m9ERXEzvastUd0qMrPi4sC01rboYi+O7mdcTskUVPF/0lBn/sc5UK06d7XbqiDj5
BZ8yeGEEYd0D3BtbWtLdD19qGRaX346oQwD+/OEg4yfW20vAlVV5CLR9VJ9bNq8P
YRqkZ6GFX1Y75wAiVJmyJn9vVT1S+Jj7Lq8f3MeyomLGpX+8THEoo+5aps93tdjs
FEX13BEzzoCVbWA5vlLMkkVLaUuHjObQK9H+9MyyJLPCCb1n3wuAwfpAKfEh/fJo
MS0/dKyfuaj5WdHo59TSvPxszzBOKYDr8MU1t/EX9UxCCngxVsLNGc4fMQB0HT8f
8IrWtxbPbtP6bzzfvzmwjbA0BAis04voWM0Tqi59pHjQpLkOUtWo7vaQ259YfQ0e
DJt0u4T9jtff0SnahNlJb5SUaaVtG/04XucjOrI2Sy6O2FAGj5uWeXyIVAq3Tk2/
uBGehS0IphgD9prmXNlAbFwN31bLWcX3igoICVH+BgI2kwknVtkEZUR8GfDRE9G7
0bjKdNKsAqK5V1HO9CnOPuK8nvpEZPWcnvGexcb0YD6CGSZYNIpo7I8Ac4CImt8G
g2CBgLngyS/8GXNebvD6hO3G0mymzsUDiMpyHNzpybL+URPnnmcWxIEbLtfKB1rb
f6YN4xoAUNLnAZ5SNvAlDR+xiRy7X2gq8BTKK+vXjryN866UvpLx44S48hI2gFTl
3sBZvcbEtGwPq14uruA922r57VHdB9ErkONHoa+dgTpSVBY8Iudk/pHAKbWqe1D0
9LZCCxbEEr+ztAShDVroU45ArQkYL9vR5xmN5LPHZrXLvOGwScPzkGgPGOCGwNZu
My+6lDZApcvMV+HLEi4oUMXkRonaxsHJDfzQtCrwDWuVjjsY4nOwP+KdXq3LMLCJ
P9n9PmoNzzq39vRw/oqScboRQXsrbZ/1ofgEyQKbcA4y9D9G6VkGZhocd9XEhjxq
n7gANTJ7areo2mb4Gqsbjx//c4K0emqCqLQ9swz5z0YMz1iVE0YKpSZ+gzoRkSmI
ajXPAvFfMe56C2Ae4i6PIuExHGrvZnUm3eKH6qAx3O8tH4+Zm0vGistJiqaqVaNn
PHSMjqsxtPx2U+CRudiomh0GegReBrwzOgPA07yd9vV1Nk0PErLaluQSCuDpRnml
7n/iymokmi6gvrE3ony24V3UzMnChruZuBWQ+pLXU8cd5tTdODeAsEanxGAEutd9
T9yAwwSxQYSkGJqSGKnjtwYGv65MKbfsV+lrnwwpcHLroVzxeVU72ifsj1keye4J
FQ8102IA0kS9vDO6nPG0Y4XrKcr/pDdTk+fFrBXZIf2vxTmGwIl6bak3RU7YPp6M
l5xqA41gX639wOmQWpFc9WLkZWI6a3rk4Y+YOX3EoEXkP8by5FUa+9P50GMvoFSW
O5OTCJS3nDaCqeQhOrQSdtajHvioE/hMnC9y7SF24k5whKc30HP8HAgMDHawbRyu
5fvEXhd/dOnSvW03CvaFlVFNnzg63llFvh/vbcAJRFKa90/RS7URN8N60PjqTK0+
3jaAt/dqqiEdQDybgNAv12eHilqBsNmFffnhp2dMk1uvJg7EQciZfqpgVAKYQr+p
OU7xcmbN+ksNdB1acBJp7f2q7lnyA+vTaqnG1sfd4aDeprNVGu6nUyrYhUb9y7HG
G4xaSb7Khp7882wJoZAKBxyPNHrSDmQaRzLCKUxDquzfvJWIdsDf8NeFJZZxx3pM
46cjM8TcJGps2Um4wPq3OXw6ivUK7D4xhujSgUjZcZS4TjOTUiiF2+EQyHX783nK
9K4jfolWjf0QCifGF0WfcTmIxdC97KgvdGQ85POVimufm12H9H7PzE5Eva0ob3vF
Ou0FiFvj3XgIH6gn6HtSEDEBoxT//qgfczY06XoX0LbIe9wsesAndL9bJXljo81s
cFgR7R/I08WSNUewVmk/2cFqfnjsJS283vUjuPEMJGOWEJ8v020qB3xo22BKMRng
/2GWhe1eFV1W5Kh8aaImHs6L8VaAJHfz4G2P146meltrvWuZsBdkQMu7nuY9VLoe
eHcn+ol9QPxgjeFuTvjixSRep4dR76NVw9ch9y63EUHhrPZufR6TIU6Kofv1DIZS
wwz5gTl8jBLu3fmMwAAwyz1pxOEHpHfq5Kayrr6iPKzLVJnUO0oqQbkPNPGGItuw
2JEvBoUjIO0YBwnUbAXW+szkqOrSPcGCG5wEqRVNQS+b/RVuGNqvHypvQr5S9Nnx
r6/EVQCRwi29imfTygrWLhM/3DuqqXxXspkpq+lXyEQg1V1UjV8gk5KRSqcd8wbE
YGzxTWRiE2/847CSl1m9ANNHfTfoFMlZikJTO8rVMaATZOWsjmv99ZPDD2FAOfKB
SgflJjySavZeMFAbQw8UAAnoHf7I25D4pjjSF5ONUrnh+1nQbRniVvdKSkqxI1DC
SbX96uw+c3QQpCCP8C2Kuk7rytWtSeSy7/OXuVCqNG6kNoPZuyJ64OCC3s/N06NH
mJqD/fQ9eagqokCK5Ky2wKFXk1vbVrb4/Vkkyk4r9fa17Fel5sCknyVNhDPKCNQO
auNnApyztpvIPIkmSE9rB6D7nPPxzdEiARHBEAHitA3BSnMrSyoCxqJVA/2G6mgh
UsfbSV+n9niZdZTysxTYX9YPpZT/I2E/mWkMHjEPc4E1L4LDfcKwLAFVYXzDEAp6
Dk+zezBPi3TUNOEQFyq5sCXqGqUFXKUedmtRq0Ua49iPDKAzzXHKXK8R7fKjNjSN
Uoh+Bq03pv+m8ERlOSLRImg46NtfG5RqpLTMrXFkyIyDj8uqU9fIwJbjlc64mGih
AfGrxgwYK7pkDnTt9Jr4haL92NfmWlZl6dHlboUTlmvLvvqZkw35wOZCfPHBO4oO
D+3ZnFYWyUe4xZs8S30N/2A5fiZ5poTPgmD4EfeUbiETjj3hyTI0zLDiBWq7QSuB
6ZJ3811HTzsR1waCbn1R0R92u9efNcDMCa9PkptE7ITvFhbPC6JnzpAehOSFT7XO
SxFAuutR5NkDpnUqZYxKK4L1hcOnVV6z+c9EUVGhlhjf/cgD6yGfC1QRFrxgH3JI
qcU2N7KUldQxs+RqbDLQpqlM1WyQxRBvItF9dGU2ttIHXHMKGUkU5h7DNnTf2I3H
eu0GFANC3iEHS4cXEzdEe6N1skEefsNuZc5VoIqgWzpGUADdTd0BjdM+rMb0r5qG
H2JhXHuVISvYT7Ka4oUvkRcnrceKb8jfUEEn7BeqqVtBzoU388bmKP76PfWrgZGE
tbEAJUtYbASE7yGI66VN7/KZk0KDSCM5Pspa8qrdo21TVuUb7R5YLmbNacDQlzMO
Cb88FEishxeHhKSxBVihJy0vDlhh79GYwxeVk1UgEecXj8+DOarulS9eerxDfGn3
tSx0IWOwv2QYetx954cavwcpGwb/bHI3TZdmj2R+5foNISG5CgEVMpM/kgLzOXHP
AS0kGJdJ5NOzN2zApxNg0hb93YGAODLA9LsRfbgkGzaNG4hS4mMkyRqJLNksRXl5
37nT+VNxSqhjSrVfhKgS//l0gXptgicMJqwuktkPejq7V2zi7Jo9Dp7/niuW8q8d
U44wlyqQZKSzoptV4niJ6XPaE3rvEcWS7Org5kD61V5qgWNx324VQFX9GJFAjp2v
BA4NIbblHA+sAO4pVbNjDmKcCXTodVrhukqk253M4vnTN4X/S4ZR22AgRuFi5uzV
SQPjrQGDOR/dvCcBFzkO1tNlrgVLjPd79PirpjgDjDTWf7+nKZqANSpDqsBw1/8i
KPfQjK8TKT2FVQCoVBPO+A1ga/CDc5IDt5mgB6R5YPwPnngBGCNc+2sqhdPQpZsV
FSBarJM3SXGRSFOcr12R8J8E/zHHxcqYkbM7Evgvbk0WXZqYZruNjlT0xyVLjMFn
ikfOZ7HEZh62mZvGyy1KmV2stQaFUmeGTn+fRPmFJAofGM2ByIavzUHtk55GmEud
/D4+owfJbPOD7wKN6vRBAAM6ZFkXUfQt1QpjkHN4yLaEZGfYZZ29wuHsvYEwh6Jp
I1orRrPdsnw162WfqM+ThWVZ+Po5zOI5ZFq0DwYpffJtMcy05cGZYitp3ticbCix
aApFWJVUoJ/Gtr0D6YsK2uAMl3USYaoFtCk6EkhKKet5H5OhTGiRkkGaWQyLIWjo
qZGveu7aP5tTyAlq7XmzG/z2cBoA3OJxqitYT8vMEfpAbeQuGzZnam5iVPfVyNuT
toLQpBhw6jh0OqOpsLkr4KG8/mu3EGQKTz63G5gWhzLE+815siK32z9xobm+LePM
kosWevrfemaotDxVngzWMZla+y8lSNHn/Egdww22B+EoC+a3F3xzWEQxBLZKX2zQ
/o7sRl9ao56lOEX/n5kZbxjrGSfStqIevrj+OUmptThFXxtdsL+m4PcrZ3SYxDrT
0Je6qjvwiQeL1QaMZK/itk0WBDcM0IYzgmcLxSUT/0SGTJs5mNySg7iWss9eTEyI
LPU7x9v3caBsU56wEUqIupcvsxPZixicaebRj/2xmipqZ2L7N60N8swDQ4C2WSO5
5WABYjHRAOUx3WSQaklsmswEhyItIyM0P+T/q9PP0+dYAitOlcNTX0OhmJmQr2OK
aypw1aHY0j7WbNw2I6K7dVG37f7hiu5aWgxOWqaV0AJVNu8mzGiKBNRbnVrRsqmi
Y9ieHFvGGY9tVzFVF6n/bdHw7XGUDv2gRISB2R1T89YAMtWxb4X2k25ya9rpxqDu
jWY+E2b1MeEmh3cOiTyl0zxAbtdNs5x48Mh7h7ofggogkuxu8iORX2yNt8qjNKX2
WlD4+Ftd8G957olntC3ejEXyd+boufFrm/NX2Z3rp0idU1E6QfWpPg2Ywcj7HfDA
oTG9bhi4vnPN4+bnQCHp7zcBWTCbX2d0S51gAN3NSvW8CZmBqC1V3oFf5+DYMKoC
YH8qwYDemU0Q298RbQVXkEL6m9DTj4jzzzslBoGAnkrZvYCF7hdLLVBVDNa3PNfk
dJcTkYlW+oOme2AM13HfnR/jIPm/idLt0PACeW5pqPzWf9nx3wcftoAHKKQvpbhs
Xys/lQPXpZmgiTIVVlAKQAV1zvBwX9hMhZDTITs9EL2ctMblu4f8Mh4/dPu/moLc
u10oFJ1lgH5/kb2NK412OATLayRerDgHcHMEk/rWVsRSdy1m/ynTM2RtLtgMcBS+
srsgYJ0WNv7nKGtaUtfVwYLXkQBlA+1dlsyETwhdq1nfxi7zucg+0l0+EBW+M2KE
+ACeNeNPHUh1rKhCinNHI2GGsm9URnApyyGMQXwbguwffhFnshoRsTGNziG3hDMe
jOXPhUHZ5IRZlYveJ2NvM1NdMYcnFYnQuy7MWcvXPxZDiLECepw6IgPhSrL7VZGj
/hICK3+WOc2WW6zidKhCvSjfBK0LM0iE+EKwGA55mMpr9kqKRGybi/hAZM44/pJn
msFkWRhyCl2rTsnlwz8lwbuLeykQK5eVlnY6csbnxk/b5hWEd4UDWA2TiV/2hh2H
Zfh0TA8CVnSiV4HDqmbHDs7BK6ZR2KUXOTSpvhkkHV5V0OuppWhfNKOiJzedSNyi
5hb61krPeb2ql4aNvPx2In99qHhYx5jKBXZE8ypH8+Z3+DrtXdKMvgxo0OAMhXcv
e5ZxseMsUOmrI7TALNWwGvy/BfhciaknNd4rSNl+S0Se8QU+6eguWS6Ig0IrOsy9
gHm639Kl39HE8qP5vy3tTH60nQd6+soxbRsLy/+rCjZrX9VEF88DiUjqYnYtwDL1
cqHV/SVC0Un8UhOx5HXZXl5peGSAZH5UuTcVd5AJ7iGWAvB2OfT+4vwI9UK85O/U
L3NmgaoBrNgg6pTF38UjuIvEMvIRNnKYwuQkJ51v8X8x+1yL/5Q8yELFRYmUmxtu
5iRNlGO9pM1RoSnrPbQoV30P16pcz2qhVs5r+UFTREzN7RQrKzoQiGQuE32y6F49
u9AZm+14obvhERxxqplDEpUlAhZYs0aeCkrjsxv4uqTCt3fY+HV8TJLsDQwtvdez
8yMoStrU32WyNbgrAAypYSzW2wJhWPc7xAtjuH1WlZGtdGv/jhiWNm8CQDbsM/Ev
lV4ayvze70aUYg/Uq8exwWVJtXL3Q3cw3Zzp78o8x6cq8rS6hZHSew8aTw2FbUXf
WAoLQbKqR4K8OZd525xWlRshyBtJCvhHkXjVDqAx2m7fL4xcJc6gaIqtW3AyAMA6
Ey2FHaQsmo3wnF2J7g3XSfPv/nBYJsH0R+WMPxVR/ylJ3dl0vVtjq29d4hCRpeek
cZUIC5d/cyY81B2MUbsD6DeoLwmZwV5jS3EPSz1nmi1GpKgVqQZ2JhhfQT2JKCT1
jIyQUaadh64l/+Vu26rCcpQg7iS0R7aRWbZTjGDTg0tax6zp0oJAGBFFgXIlAJFb
vG9DhDhuNrz+74T8WCwXEkl6atHXtFObn/ZkX8unnTE6sVqfmWAY0HdeSivd6GkG
TOPJlDKAS0v4Lrw5+m0giEG/ctOa+99D5JrH/cCUqsu0uL48JabbZATen9SG+GQP
SBpd31HSPBI5YjYk99RKT2Vq3S4m6bGWuZdDaYave0FtukjSvoUhug4ALjaauB0H
JxZ0DrQLtt91ivUh8GgmE8vzdfFlg4xleug98Nwm1eb0KZR6GGVChfb/v2ThM7Pf
0uFGZf6AafcVIMZlVQyhseFSP/YRDOwKTMfTVg9BLFHajkCt4gtYXxX8IyOUBoPq
wkfT7Y7sDAC1nmmqbJsfhnu8y7pFuREUwngD60CZMRLHsJ8RfBtsApTgEugNXpbl
M9PudCLzcmCq65N+zbqNT1qtTrJ4gTSUkk969mYOz/kzvUsHmrysgySBOEQKkkkt
dC+eK0ujWSzr7XwkujPppIJ/Ky9GEf9pedr+9zD44sb4mTfbYdzmZGQSKX6VFqDP
4W8mNtgdykm+7e/5WjRmqic8Z3Zc4k76QA7OKBAriWxZ4d3s3jxql2becK2le4+U
mmRcBNLctxsxbheAUzCI9Ysm2VrC7PYpwpi31xZhCFcryzvpDDnyglZ6KGX6CK6I
oBhjciyBzXAP+3rohtCx9CS9qpzrgRcM1kqipTfPLmNyxzpn+NZrz+mTp8ZreR+g
YwW6bRMLCDpMZrzU7clFmysjlS+Bc05KcCxn8rUIylaReeqpeZF347aZJC5tX4SK
U2oL14G/qG9ba/BsjEsnMsSGEArT42VraG23TJ1lgHQ24r00bYYyVkePocybDJdb
SWhHppBh5KyrypADSM+UpxUgZMShAVDch8nVrRH6hTZKDmUhwS7HT8WZL8E+65Hi
RHcaqX9OQBiVmD/kcP99Lf/VDcIbV/gw/kmbmhU7kpr1J1l8/GjgP9mQfEqDp4MC
k/z5Z6IRulVSYffgGPPUsbAU3eb0VICBPiQ46zGhr1Cz6Z/cO2X0LLbV69uOGtdo
6vHkoRDQbxALhvrhBZjDECQjnzWbAKGFMAh4Doqw7NoXAcPk09mDA0QOu0cHGZw3
B+FUfI3UCMeSRvVodJ/YHQduX1XXQgEql5QFCm1zcL3BcwqW4aF1V5UyOMmYKsYJ
92xhuKAMijBdwZTX4xpWniN9hC0UimFqEC9rdkBKVuGnwT5PRr4PJM6y3U0U0FAH
nXyDOKP7IXkAz+cO1AocU5twGhKdKPXtsvit5f8CXdWFBJ6AtPcUn0ba7mJqNw6D
AgcNjZLo8qXGjqKAQXMtpqirugpzdRgQEnlV/OEkaMDU1wMDTgm1H7bTNSdc/Zu9
hVKymPpI7scyN3OZC0Ee+7NwtM3h5z3s018GR98fyQChhZzfgDqw9IcA1+zawBrG
5Y+48ZQap5l/fZAmisd7HpUhXXMTcKB3s5sUb305LPk9mE20VU8sd+7uscqWPeHs
JD/O+BYGhezrib/NoN95mS6crUeAvJJZxVMXgVYM/JIFoI3JHfyBxR5ySdP3LlJl
suG7Y6lFXEDLWfIwOmJBQFMJyeqYONu622e6e5bvepDY61F9XIgS3EiBHJuvBA0R
tmtycZjo5ABgetKX3lfgVQdwEC7EnUEGud+MAycWfef8eLBVee16z85OTb+N/Nq1
GEEd952LopUTfpKGKVP2aqRhYgtRZjq06wYu1VCcwLVOPiavHHm8oCjCvcFZht32
kUZrEK4snLwyOipq+eZCNP1F2rf/Ofi0i5yyN9Hl1Q0zFxMMYyHTDsNTE5fSt5y2
3NOUokzx0WAkQH4yJdAhFzKTFDRyZ9cl93ULfz95hxZ/LQ/S3j+bw/WQqmpOEUi5
t3pvFzN6ZTMJ3WIqt7rNbu4dtmU+hTud0ttrBA1v5W7ZGucZTX/hdQXRY30UCTnu
abim0O6j1JQGR2mfxbYQJmNzUosnkQXifWbVIrF8JKGF4M0A87LhaYq76uxEM3lW
90DQw8B+CnGhcVKhQJiK8UgXj8r8yEOhzgwzRYMNFTH/xi2A1XaSkqC6GvBmfpJZ
AMTafz2l0CQVIc5AUq3VwYZz5BZyJv/HZqJcehIBxEipnWJMquwscuUmXZCbrd4Z
k4ba9WvXLQ04lAYNG4hayF3Mpf2cVZEjHFDoqPrxBYSMmoirJv07TSS+r0DcNSBA
EqECJHz7saGzL4I4lYMZuySrVNtCagdR1PE/lGQc3kvHeiPosAzw3gmicevG8w9q
LtrJezwil92XsWfr7f3ZiWlVrdRu4UorOD/rcC4g4DrYF9ZvNCohhrOOs9eKdDEo
17ukrNaaUVn4q5boulIU+auM747VuZ2TFfFZ/YMV+KEwYuORZo0KTXOcFKaBsUpS
ThYP9UxQSgJdTPXFgMBuAuEmhz8DCw+rDA4vUo8Atd+W7d5q0WW6L409OjJT2ATW
2Xfkq6rNVNpcWW7czqM/1U8cdlSUamw8X0+C7pSPvrB5sQeFVqIUyVi6uIK5+g1G
YCXneA7Vu0lFTp064ppELRT7Fj9DHUsxQQcYXrhb5jLAudK77ZYTNfTp5Q8NxlJT
gQ3aoR3DszTyvafzyHJeM/x518jQvFTUwJIoFRl7jx2ZYA7VHK9onuZGlZ1jJeXw
Pi5NM54fmFwJZEiKPxj5hI6RgczlZp3rBgsYGlq4GDWgB/6KljOuC0Fg10dVWbmc
aks3Pk89Dahp2/JGB5MNHVFSxIIQpL1e798abJG/QXGfdH5OdsDFA56bTBpiXbLg
CKlkm0Dj1uSPrh2y583t2WPHtq0X1hcuSNAQEHfU5bO+zzV9h06YAl0V19hGxCZC
JH5fbAlkbU8YHlubH7sqVmCHx5n2jDjxXLgNIaFllHcYlOKVhzqQEwBDfxQ9DAvb
pH0M9zhY8dXqjWlTNZLXFNvymXBeCKT9LcO9Sh8z21isjy+MCMVqhz6zCXrLSoAy
4ZXLYmx2dyCPOcKc+Z0zo4g1RKG2ZVXJU4uv3HZGzKncUs0aGt6f9loX600K14En
pugg2S6fbGyPJZoPvbyQ1ADtAKraa/w7b6dWCfi7r75Z/OmT1gqwLd5dlRgO7Kru
2wdO4I2/4t2eW4/iZB1zCoGTqcblDM56GZT1JkqSev4K3g9moZ9ZX1ayu+mOV0zX
6iBOAfw8iMvJnv5NmFh9f3og3V+kv0iRp0EDsrkCXBA9xzrweeMKoJb3S+FVVHa0
/4D1FBmLIxuKdxvv4QogpwjTIO2TJnv9ZyHor+Y5VFXJXWeN8mDPdTY6ZtjmbNd9
ft3QawOEJn3pxqjbQSpCIU75+2rkih04kCvblev4hmrkBfMYb7UWoN9gX4NbjDWS
dOMW7d0XCk+zxSfPQsE8znExyWko3hwpE7sbFs9ZvaiIsKtCeqUbQGSzbprTiBvf
uTkCFOY5l7sB0ESZl7ymcRUXKB6PhGgmIMHSgjhwe5UXQBu9gTbpPE4JujKucu1i
TzS+yfYMPxEyypnNu90w0wh0WIvI28LmCwwwjcXbAmDPdaeBU59G5834INdKwL1s
JfQ/6WOp2QNys04IYVst7VG1NIsJatfH3WmCn/FuGIUXC21XICHpoWmktLVyFddj
kVdZDtMS1JYz3W8u0PLCwKCIlSphAFLLAyNBZkSLE6b5ZOy7YQSEoF6UVlyqATMX
Em0CeXAXAkGIzKmt84VzSJQSMuakTTXsNdG2HPByNG/6miVntVZVUOwlLUEUJdGG
KrqzhzqN8O3VLqKhJ+6g2MtXwQcst141dw1KMDNDpLEhAcrRQtCoFXzuQvLd+v+W
aAuspspS29qpkB0GTphJ7TasZT/F0pjnOU2bZF/AvTKzE3ie9c2jVhVzreaG42Jr
MiykaMd8lOI8viN4BYuWj0YlEAznjOHOQJlLFBKYyn5srxEO2qT0EgvSocRVyMmX
1t487vlgdyc++8vMELon/DDnDG8xxYNcP1yUjFrQeookWo0cTuTSl0CE7zM0fVuZ
fFQ8SbyZRC7xAqhfs3G+ZOn+eiAB63QkUFT+Gb6R3MRUFGGYQImv4sY7cJxMFaBw
+hEjp54ELJ5O1/U7hojvTZ0U1heEe/1Rw6IJulz0Vrqbfnujc0HqlHhiM3YKmTP2
7afxWe9Y9LUx/eJeMMYIHzcKC5QzelYm1G2Yw/Xt05/dYDZq0ThLAXam1lHOuvhk
kz7df829bEC5d+xVDvXFsfm0dlSDYHoGn4Q7i/BPEAUVQwTO5gDM8Kmf0BsWqMPe
s6tHv1fFr7jw8xm57hDB1SfBx2d3iUwtWRjGdeha3eIdgVjqpwRALZ02RehWxmP1
R5h8hEYfFh+WdlD0weLXfloEPzF2jjr0lVjAFo6nqKDZSnYcnd5l5NMSI4WssNI2
kyN+VmEF889F6DIfShi4pb4hRMvVzDhRrmNNHwsqlLnSovD0LOWNs51D38tGG5AI
4WNa+wrLmXohYR6+/hnotHRdH2gl2OeV6AOwprjHxqRsVeRJ3guR9jZXsXPo3JR5
3bmf51XAnz4vc2gZDzbtlkKYchY/3vd8dWBEFxRkqWb9iFUu5GZ0r22Zb7fMKZlK
dGzjGLkMIRqrbIYq5odsmq1Jjzm/h2W7rS+JhwbFMwvc0H8baU3+3nYYtMonATXa
nddF4hVAWKoRM/WsNNHRDojlS7km2SE6OqGIoJUyiyiuSI0rXoBSZ4IJ2J9Iehpz
Uh7Bjw2rcq5f7xOeu4daAHj6qC5y4FNxdv4Q3jGn2Gnt61Dnyo4jFojjCrWB1dVK
klvmr9n8l30CaqoFDYY9eLcWVVJA1MWHUs/ScgyfxgleHRHjZ3FCtYhiaoLHb+EG
XjRTc+bM8JkjzzFtfhOm/AAScecyQyF0+KLNvbX5o6mFAyp54nuD00Zib5lpYlCF
E47zl72Cz7W5PEkKqUwIydjemZQf3n6W0s9tR+a2cmPV9qF+XBp4q3uceZWLiefU
eMpEP68iwjzU+J+l+eRdIYVkCDtE4MsfSkJso9EV8D8mXsO82doUK/gtu7WGOQoy
5GGWHhmomsWJGuoCDjFJ7L+X9eoj4V5CYbY2c2f1cmBeF0DzpR6DMWjSd+6BENcp
VgAIk8MaMcW9BRWu5yuTK/ttH14YVq0wAv5PiZ5tZh40JIqeK5pDFjRiF6VTH14T
anj8HqSQoehFeKjzr3CoMGoNy61L2dRhMawmnUc2z5rbQUqF0riZ+6pY6BEr3z0w
k2MLpdlteiabMVGw0X3T86xSOOkf4aiuvtLL7ELwwCxHT1KZ9WXzduJOQO0RKDm0
NGrAKpLKEabTuUxLo0pmB1XY5acmNFf/h2wyDfYX+5oBqiAkqPFJT5y7WGwlKBVI
NyXqdd+6vYdAsCK88Dmm87ADUDQpJ2bGoCLy24/kThK4H6k2j56iIREfE/VpwF0H
CKhTSJmDR8s6VZVM5qnvRV5scExEUmJkekI/GQ2McE8VjfAjExqPjXRqO5U/uc/F
lhw8j8ZeQ4NTaRSEM4Y3sDbRLGys8QkOECCpuHP6GLKDeN8epbpAef6Q9tpqpbz7
s+r8UeY0AWm3Mqe0tTEMA9+qqzly7ZbKdN6boCLBAZemHeid5BNWxTZK4v/mpcQC
1UPLoo+Y6bE+6HGWJClrKux9xHD/RMj92WZ6TDm5PMhsVmZuVIE+OxJ8zNBfayNm
LKnP6u2xXwuwQSkUXfBjn4v+fMPSunDfP6qc/JQ6AVIGOo2GYLHc3lnNbjJ3RKpb
QID+VuAeMjGrvtAxyAScySl0aGQhRhnajL6tmaEGnpqDDm9jRh0KMfJed1tr6OIq
X7zJOvo9npYtQeiempC5g3XUng++2h2WgubbR9P4qdvQhnvCM1//UPCxDjV5GS5r
hFlBA1WURqkU6K7FKz4MU587w1jTzvPshaI0eLDjh0d1hAMsmCv9Q37iT+NU/T7R
0+clDL2KW+vWPnEmPBjAhB0DACd2oWJvciaR3A3WkquNrcufrhF3dzB0f8bqRT+L
lbe4Kodw8oYzUa8Wq9soyKck0sD4hbM+C86GPPpCwt4y1tmIKxMpm/pcs/xeZwpP
9Jv6ldyL4MeUkPLy6/w2VF5+r4Zcm4pjLc/gO77VlVG1b9WScolG1um6VXXA/Kr2
6YDVJvU/K++SubjTnYEXhHg0K5ln17Q6fQ9ciTpnBcpe37f8aF2Zmh8A+QPd3vJs
r23XquGNe7FM+rJV0KicrTn+Gwttmw8nIWkv0FX+8hF24GkTnmpTKpK7Eq7StU58
nwNmSNi+aSLLDKhHh8ow//+LSt+ZAw9JKJPlorjvVJSYreHYCeR9R4SYwnRpznkj
9WT+u23JlWdacskCSuKzGsobi/IoCwnZLDwm/tDIJVANl+APxNCu/pGsaerDnQ2W
fjyV1wUIlierfzVSNajKAkwy/oqkH8IP57QELPcrWH03cmXsOAjjfQnWHQIUrvmt
ZPf77H0RdIjA1HZNgvz5SeGtgl7zSppv5P0grEQoL1fU/jEIHgmpsEJnItLFhGuF
Hlr1zjV0xMMC4AFEJqJWtketRz4GT7PEl/8M5VceURXhhqwIIA1etGPrehwyf4QD
cC4wUMj9LB6cdcztqSM+QLyVS7DUl03Ee6ihE/PXJCGDs52NpBaq3Ww7l4FoWdpR
YlTxMSF4WXnRKw1eYKPupK4TwHp410M/HeVYpTnsvIXdxl2NaFm7DSFZ5K5Ls4NI
5zSAoIPMonGEmWa41iZlNzTTGUbXzb09amjOicZhc9P1+wqEIkYh5aVObzWBoFiw
gbtQlPNm0HVWAU+tpXgL2d8BggFt39NE6f0n6ngyVH2FvZvi3IdCrT0lRUAaWLQj
vY3bsXRo5gja0Dlw2LSULCpfP5OAgCUvDMUINauv0apTx8ZOdFJWzAsyP4BRajCy
9tFBpZunUJyVtkOHw9Mv4OeB/yFpxIM9MhnAY7VHHWCcc2a2ExibG1WNXRpASJe4
q/jiZDI8JyOp+BVTYlgx9+DLE3+9QdS54+x7qvOGJlYb7w05n3I3YQz2hHzgGsLe
vJYlNgFHYXumGzXMMe627AmFRwjIoPOD05aARCnmVGUrm6CFe0K9fGRAcbuxF1x6
8kgCpy7nFjcrWHNECOSTlIBagg6RtG4Pai9Y4agXpDAYKrmhwRBtMcUvoRTaeJmV
dY+ixkcd3e3zgmJ2PRHtHEPfC7AGsiwOohhwVAvto359VvFv+IT0jA1PxVOg5CzS
+gMTfesEwLHbhAftLVwB0ILgZ656bL9JX9+Ckgdfdlzg1L8Vs9lAWnTaeam3KZrU
47GMC2TL0JTnyUoyTDRJomfD6/Nyy2AI1m/T7KTfQ7uqXuvTxSES0j04OHcYJLiw
oGPs3TnoJjKiPfVlk9dK7SpxYR2ZHm0P+KJ5HztuVoAgGYefjsF48M6vKqFTxyhC
UO4+qVSVaW+E1DWMFVZ1M3SFzFXDSWm5qWul6AH9aej5H1qyqaxsa7e6oWGy4Hoc
mMrxcKnpo3EpjuF0qyfAsV2FqM+nB6sGSRVGOGBytEqXsXQ2JhL4fmRfSgmClKUj
Ld7k4GifqKNStfnbnEiAZ4bvTPhw/PBKDTskHl46mslgF8Albf+T2HD10KpUXioy
RGM7JL72LzDEINHCTFnBahqXs4vhFoo4hWpVZREc19A84Zp+DJFmDGbUwZhnKclM
5M+ufZKFPz8nzrCXVjPzRBDhJvK0bAbjoLL1wPY0TIlDigPzNNS/X+PnKZZ+iVhg
XdeGCOUE0FH4p/OSIlqSSsL66TB2iQ2RLfG5h+M6wkHb0oQ2ozO0bMlRzN0fhSea
NdluF84zhAXdMbvso9jtkLsuTtz3YPVLeJKzI1MSfimflh4JmkjFNfDAuR5/pzOw
Q+dCE932OrT82k34gWR1TCL2zTPasKcFf5zYwEEyig2CB20n/icMrjroClBSJU9s
05iEkmw6+Iz1SFA1oPNmH8ykyrgl0zzSNxujqhjXJH72x5A9U1/lZAVhPPHBsAlq
zM76zDIbARhnMR52eX8ad6304OjGT97MUlqd+vSl5Pkt7zK53ABXndmreP1kZ1W8
+LLiQgYPfdfXZs9uGy+7KGjIDv93UlwP+I8GZocIm0Z2UKWSknUahtZgvW1P2bql
cOZwxH35+/Y5DqTr2cUl1olURm94QuOswp1KhH9npgEhZpDQ6cEr1D0JfzmkKmwZ
EEenpsOezQLhSm2n6HOAp6L6cXxpaXF2eLmUZMZfh5nKkaUAQzc5EV0ns4z2hRqn
6wbQ+TBR5tBYnJWMk84xplpgsUiohEa6ZEw5SB5uWr5RH3S5pPhOsJ33QkaKnBPq
xX23kEmYUp7hu2sqjIsM2OwI6i8KHpkjBACLI5R0i7INveL79GN75pmTrGogOA1s
VIRxOh5Wh2I45TMIIssyQgckyjtGS9Yshsom4lFmFor3SzueSbPFWIDqdhD3RtoZ
j8jBey0BSFh9vQJeohnrdepxSLDEmifcmKEpLINfdhrJBZqZCNtrpKFqzCZFjq+6
T12Lh+jECS6vdojvo7fzIp4cXT04fofqiUyYNSYvxgmpnfHaN9V6fI6+fQh13kxo
tjmQhrlmW6t37e1euEwmiu+eC4LGZ4q6OGiUvKCHn7P/9oGZO4WT5Jek4XWjVOkR
6zY5DAQZHqL/cZ5IOA4SFnS6sYrnjEU2dL+qEptWKBEgxuIQph0SjViU4heia72L
w6xeqMy2IScjwel/DLIxhhoLBciuesRDpRUGAlj3UQOYvoAPS491Fcf1Wyp3Wk2+
UN9NFOkiG5lRnhfiUP2f6E9DZa3hERG0uyjkzImWVVg9N3N6qYXrFpe1PWri/i4A
4xPm89xFNeUJh3tMAvVZfwIzrG3zbkhv+tubV9Y0MoBud5sQ9Piogz5/oBIgd6Ui
DpFaMDy24M0Fsw9vdm3lc8YwK9sqtXbu+4CC5vwkZQjNEO2A+FkZkW0InjWO6GzH
XweyTw8WyAceA7gWky28psXevtO991fXWoq/GxG/3CCaHFRDVTiRDENlqYHHYu7Y
EusvLxuwoL3+CsjFiFRjEibAA4/lduglc41hBj1eZ6XArIMJTm+FWw+u5hA+Fefh
rrBGWRc7LNgqGscJ9eLTsYmdyKQOtcJJiX4s26c69gqowRUG0ZRCwJ5F0wFzy00t
9oLa5+OiZbmamuqKqsaZZpVjEeLdYNCRuFCTC6GO3meUHF1o2kKsaJxUhXAD8GzE
Qt27/9rPsm+/CP6vzQm7CXVKQ0Cs0t4UhVfRRuExRCC7CXluoGxzMZjI9r2MEqu1
A2k3uzif4LJ8ir0Kt74VkrvGF4nIoqhXVhx9LIAK9y+/OveVWY3MW7g/77IFy6By
wiLjU0e3w+tpalClHTA2F+VfyteaByxIQ68DFr0aOn5MLMK1ILoKKHE/zzqtHzVx
jhAgeIkb4VMZzkbcKNOk2TfTNQnxeLz65IWacFcmtbyPf50KYFoYwNQ9UgP3uHgi
h9gK1e9f7xSBlqhbdt3wUQxiVJ7qLOaU5teNoR168pMQJdRQqBhbCHVLnaWMSTYk
KoKeU3nb1WiIBp63xjmlpjqa0q+Hm0ogcNhpRLf4pCD9GIdoEvySuQKPeigaegDA
mAmrDPrLMCaaFk7n9otwO8IAfZXvtsEzVtkBlx+r7SGq2yHCufrabOTEZIGWBL8G
/lvMbuMtM/rabBNJf3Rht2/L3+z6PeVEArKrswAddQAw1apHTEgMU0/Jusn5w0ep
Egs0YIxIr3MD0ywRzmvgJM7DatSgqwjM9BmUv54HNR7ZKK5kTVtwI0JexnYvvvY0
AY/ZxVphY8lscLp628PFdnFJ2LqHmlr0aYJNq1V6HuHE0kDP6Mz/N9pbI0JDY2u6
tmrANDBG/co6A9ba/Qx55+RKGxBQ3efxmEMugcxc86nujyJXd3xg2Pp7seD7MD94
DEyrl/ASjZ2sGHku0701xysRTmCYkZA2DeMXvY5G0B4giEVgxymLwv0sGEi8x3yX
3syXSmW7vZZJL7/3ZuUsCL3jQzGYughIfhg+s9NlKPxtLzu4b2gx/I9QSILaybPu
HJczDNqUdhh9sBG+TlMNJr+qvf2dqOZDpYtJTqap7qC0NSvPRarLGdDOI//151dE
Dmu0iL29P3ywrrkbwQ3EOWoCGR500K3CE7u76SiqIjiCQioF3F52FW9AeUGpRSuY
UDEBHyagohuJPknnLIftaHU8yzXjRG9LSxP3JYkAbSmZVj+Lt6atdNih8cWDyTTa
t4u0891bzEsoBXRCGf7eGyUd2b7yUSwaCn0cUP3BVDUKvmTq1ULM62yZoeBRHTYJ
TyV1mltw5fB3Wr/f2OpnSloardmiN3fjlKSJ5fpwQhSyDxVf2jF/XR+JWrlVugiO
AGGHtgB3hWW9XSeQz8mOTwJB3MjDPjkRriUIyVUSNeMze6Ht/7uPIy34SQMfyeIY
87AjJaI1l6ZzVwtSJ0tXtISFtC+aVNWnRgsl1RQOcfmj87ldV/YVlFLSGgPrSYZG
1PJYHP1h32KWKbjQbwnwZUvx1kUOrVtG5JT34Lhlh/MZMT5a0pHX9vUB/FjsC+ou
ncjNkTON5Ln8IPVXrzPnYYF7aQBIalOc3XpOrUlzUs7fjWKf80Klyol7wioCd8Lw
ogLygk+0uOsVpuFP2zq3+05k4cCCdXkVYg8XPzc5C6hMfObFgNKCFWxOWosCkMkR
sC3/GdYhRYyBfFOxvHf1Sot1Atq++gGA0Qs6mI2y1kq3xrW57JT6fvBEev39Jx51
vDGhn+1bUCP8MamWbP04ZYcTqGrPfiVEHhq2PljZoqGqw1R8iW1E67jJ8ZX0pJ2S
n80sWh0k0dnylBjSKxZIhOnaG0YSv49VRefso8rdVght7vbpDm9qJe500QZit9XW
Bq83U6tePjl9yWEkKefZrQu2Bzn7ISHj+9K0AzrwDjumHYdY2DAaw42pIRpgBuEN
0uuxb2kk21/KWVXbXBC2A9XMKeTE/hBOtsD94k8MbNh/JfMexduPhPoz6NMd8TEx
KRj9ml/zXn3SaI1KifxWCtgWJ9bml33gqWiHK9CA0h9ZgWLGpYjGTAQi2owohNyb
FDNurssBI2EBt1z7LbmdeYjFFXmlp/TWDnRNlu8aN0d32H25KlwxxJFbHBidAZTt
zbKV8bAdtL8gL0phuSdZ+Y2T8hTmsNTTXwfmtdnBOrKoPB01D/hsKSGDc6+4SBl+
/p/resUpuoBQ6Y7I9zzXfxAns/VoiDlcLVig3TfJwkcKbVd3lPOOoZSGiE1cBxHP
2nBvT+X0udJyjwK60AnP4z8/UDDJN5q8VhVwsXpbaJKaq+sirRcG98X+yaNADpbX
BpkyS3pK2qTcU3f59YN4VfZbQ0+1N7lKUptoaF7nSXnkIFVDFtcX1rsNNfl6DptS
FYR84jJk0X2SWVGHruxXC0HU50SbY6FsO81Tv9C2uiwX/wusaj9Epb8nnO/EDV5I
9Lhi0nSa3u7uCFqC6rIdqefigKWCSMbfZGB6QrbiuIUmpte3hpc7+Tlqn5W6xULP
zhVe+KZ1y/qmQSaBwmPPvZR5PRnAbETMDtxn/lJYp1o6tpm0+X9ILw9qialZLju/
HEWUYbUA+ArEKy7aQJ6JZy7cTdml97WNeP87C6SsXUaDE5FKfQr6J2IYN/5Vz+WK
moGLCAjHRtdwWwnSHvcAW4C8fiDKDIi1jsCVC5mp2oe8P+Zk0M5uhLuEMTSTQcKw
Xtw2xrMMhHvC5FBoCD2Yd/lBbVNXn4qG2axOhXumt0qPKnZbRUTtvuE2LF05ILMU
YDwO7RZyklESVt2aHUyFUpHh69qjfvdDjrHjtNdLAoNo46NLvrusvSm2mlxW0TRH
wqCaoYjb/gjfNeyMQ21DLl1/HiLNicFkW8qZmRuubKauEMNz1ZBjdNDHrZTWYpAZ
dSBhE84qNcQxiqIBUdXk/PK5Rk4XqC0PyqtaYPixyYg9SVR03I3SULS1L7hsYWHM
9XULtCcaqzkZ9FIhnK6AQVJiFdzcvW+IEdY9dISr4z72Yn+HMYh/dLBXSXtsTLmk
j93XymM7aw547mQvltICUxeeKc2Gd2ga/J1eAYCS/1hSRt0rG0P22I1Q4hmqYl1a
V6NFmjKLBKiN+agXeePLLJrE1Wff7ozvPfCM3dl83ldH/jo+EiYHeiG0R7fpMPUt
TT38+Q+VdX7kOpXFs2ZzRp2V2i+f/m69tFmFhCTHaane1qAgb0mzJI5WL0DXJbjE
fiRF7Zf88lSPm2vFWhtKzx6DElwvJsq2sMms3j0aGlxysc5l2lwTxoxk/6lGWtnt
EtANhn0EBg7FgAlmEhJ0bS17wKQGWeMu6EmG0HNzBsuyv9lOi5vC3aLm4/QrOhrc
2uxHWjfN+H688GI2FRpxD8EP/N9yYdOxKdhTSc9gg/TygDCkB8UeDKmI0v0ZN4cy
+hz+yZiwitQIKZddZOm5xLHnY9g95rxYMNn1H5oI+rBTTbqEx6jtQIGaheVfgcmn
mithWv9nmPtlhxiKcOjrRX82pL2sEfU0B/Mr8mDj9U9Rtgm+xwHgJcGohva/AmfY
ivIFyoL6t+MWCG+YSCVQuUBse4RJ2bKvYFe/9WGXbpib1tqBxUZDepw/LKv6WlLp
1ulgN3WKlPPrWjJ/u6rjgJe9eBGhnwgFzdNf75ONoadQZ+fB1PwnWe1bjLirSMsv
T5GXA6nc6KFjv8Zd6HwEoUe3gTldg2d+H9L3AYitVRAmCxMlKFZO4gRdEGwDfTHY
77WqLE/X+2IzThBqQs9mM4kAHuiRHsRLNe6fHh1VyI4dfjplF6cOE0L7Dcc/hxi8
THKq56MphMFQjtltyLJzLKCAJAs6JdFNHxzoehdDwfMg6PaN3i2Nx1owOlkBrw4/
INq+AV6guA7AOWGNGpuSdApXbDQaV/ZMfyP9JCO0AmPpkmCstyxXPRPNll5IvT2w
B04tCw9XS9lTvQOEPChzNWSVh/H3WVPxfk27V8TGeHScleHEIrAzsOz8PSAMAhHJ
F2+YjgpYuI4C7Wdkqn62yzNwCaxS5N2LciTlA70qrB67Cuc35nEP2b7943pjK1+W
LPZsh7PVfkRg8cGWUPP+ZdDRUzZ1XlGStjetMfN+ADXMlP+Ix6uNRoYHugqwgrrp
hYrOqaJTs28kBt+YROWJNoX4P6JgPdgYx9uffznG0kJjIZ7gwARiDs5sPB+fFw3M
ALhVDWZ2RUx7wpPk3QIQOZwnQgkgY4iI/k6qyvRpNdCxPLpZsP7HsoQ72wHaJh+D
ECRsdR4jBmE2L+wTG01XTiZ2EXFyj3JWF7vVeAOz4BzmdTw52LtCA7VBm1OJHIoV
gCFOYSFHG4jz9lW6rPjIlQf8S+B6IbFbW/uDU+CDB9/l7dpRPDO2DSV1zigC97Xh
hzegzfEK/arbhuPRe84XIy4DkzjGKO9N5yVrWr5Su/qXNDUDxCeLRTA11+ggF0aj
fUDEMPOyN9D7Jc07hFefNfdLDxAqW/EwFu0ImnvdCVCdwE7QgC/SD6XAqDKoLSiB
GTD4HMyb9RnDqzImieTj9Jg62+mEgIc4MOPENv0InV7JaZvMRE72G6yUcWx+QalA
+hZwg6HmhKOQ88I6u5moqq++gh79zhuxTnrhoI3NFsxzZC6ruZfgT93zXCQwAdQ0
6qZMtLmxBmnzfMUR73OCI5Y1PxiYpuMh2JZGpNjLYf34nBXNdP1JWy1YmAd8PcDk
DZzCqbLwHgi/Hq4sQngV7ZAbdLqsjL+6mbOxPH+PYxwwFxWxPhLWdRfmedXolB8Z
jwbd5IundmeoXDIMM5BqVFal7FUceAkKSY+gD0nnEQIMtO0oQ1FSSaJrsFpgf/VK
0vjJQrbwZZMAs060UStUVb+gKCAZIq95wzV/QkVpcNDzchMWs4uz00hD2EgKUFSS
e7ioagjQ7HVXPADWrLhQwtEt+63A1RHDbvhpMt6nuXszEZ9/aKKigBcF44PP+ou/
h5VX2P8QqadONVsP1k1sMVii00s/hj54uoO8xUpKi5+qD1F8///lf55absTIt3XY
bFZDzqQlzzFseAuzTSPAD8woQgo23E5StwFBV+3gfwl6OhzW9fnbJaTCBe8J/s70
XZSkZqbbas0LOON5sPDkjQz1RNNsN++5xNsAVAhEAcpPmAE9ZbNVFWvhkb5V/MKb
dwuDgLDpzWEKZ98/pqtEMZLqnxAPCzhJwoTxvIPkqu/ct16kplyIZDDmO6upMLUZ
LzlimsquS8SQ7kp8q73jb/60jPnHdSiJ9pyryo1V6CSx357DJ4hfVaM/oO0aOnCd
l1+7IH0azljLPbIHxJlIIqt3/7EScw//U+fYAvORD+SHzky0PiKInsn+Eodvss/Z
vib8B67uiO+RJpSM1QvjTH4mnIDmhQePjoKsncfrHDVu0K/uqD8vNvz/Paw+X6eR
k26mvWSCRAiXSVwvojbCJ0kEiTIk3HyQZk65VYhKRhw1WND57eUy4Zt7acU0I7uO
NG697S8LxykHPMew000W0+XjOSU4qK3hx3gCvIGeTXGJ7OPphjnJIYukBRNuG1y1
9Z6bgQYFg+nKfAY1PTeojOhmqHxjfuaKeMDNyGwt2tkQQWnkiDcAvZjwBDVas73c
ndztuZYvcEOCS1Kjjz5XQ1G1WBXHeFOq08w21i350cy2UhTy1ei/p4HwkHoPKO22
9CmyVFGtUkXZPJvUovCgd88ZNHWJDMciCIQRByUTG0yxR8gjZFv1e+a+uhaWliTc
suVg56GIkEb3Ho85mKnsXvxzZRv5FnpN3+sqVbCCPc3Bd2Tcwbbe7fYbObmhTvXu
ynW2/qmZx8ZOGY+nY8p2CldfsD4XnILLwYciMj1hJ0dk+TuHioY3J9LXqy9tBSiq
QY4evS5WTqHEZyI+z9H1l2ICjF5fYh1SgOwR+3bZQJPPPab/3vgGI8ldCxPnfU4G
JTQoPwHrLls+iQFMABlSCvhCJridG8tdU5Mt3c3slrjtavo19Ab9O1i6gIpr9KnH
HVLJe4FXCqPFl/ZGW6qwfJ913tHvDdWu3A0ZG8ytp1rmxc99XMJhUAbsrHv28hVg
Tt9SskYnNzi5hfFK5Ex5/1N0NeFRUXPA0A7AvS/AB6XkmPhEtrACwYTOMmScNefh
L09AVOag5AT+WTlnrnhYCeJbje6abJMHWVkTmuBMDn1GAHXKH4U8wYCbpXF9uwzT
HPwPVr/6vKnlqr5cdz/tWyTVjgfOLFl5GPMELQMUMUrnDONeIH7B1Jq8loaOi/HE
aPay6tSFLqBsNEPAEj8mW0UFbxGKhV65ifsiv7rtcxcQSJi3Tg4SeF23jStjYcdM
i4KfudDgfFVEunfYxZeGclV8xHRkcGLoKJh9KmZHaroOYRsuLYkhjFqLH8tYkr9N
PaE9TPL/gtuO9TbA4OfO86xDzpSlNJ1/e7++CwYGNT9QliTph/ujEG5FJ83PZhs3
aMsdTvjacMXRQOvp6kmYOOcgCFu74HUo5jkTxnF0U32YF3tycbgrQjF+1d2/ZZRQ
I/HJk5RAGDororAwkItODMziULDSyqwiKqTQBYHtlqqcwABY516wG5qW25xLsCmq
DGSTknrqJ6vVoPzLiWXwScgi8bJZHEf2ODbhifR2bpDGjCKVsj4uZd1PbnQyKrNB
F25rbNB6+g8tsZEj6X1CWA5CkYq3eGivQcjfBOpHt1BD9tH+VxfGPCn6JZYygvwL
0J4eKdKk+IwO/qt3N14bnGkRh0+I6TH2rIjhmrMCzeWnDp+gg8h1eFPPsI2PBMCc
2mRAgEcMEgCwwL9MpwIytooQnzo2zpa2PPSHqwh8J9nJvvibEVCMO77x5/sreG7/
ZR+gTkqKdpDQK53Ijq9ELhuuD3tKUuQcvI17k2Bqcjs/uyWclMhbIjgkRBkNS6MX
//TnwJAUJ/aaC5IamkBXD4tCCpOEQzLxcfKjLnxMszYpBg5WLqKUDn6ojGutt7vf
2FCNkUj5vHDRWwBBnPTwN6R95pF9hh38XJq2JjRtMWTmFLjKuhZo25DpDw68S9T4
htLJTeDeQvYIA+tZmN9Nu3P9LYz80xN+TFnJDbFDBkFohrxGuVE1t516/EjPlnTI
AQdGTzUEwrSs0aN1JYdI6wV3Li9iuV2YhTUlYi5xJIgQ/RZ2ujGRqNr6GlGiOfoM
zsVG6UV32qZZcE8x5HSHH+6I6T4+cUwJjnUavEBLjwJKadh6mUFZNigoqw5nzoGj
oYNvztu4SW6JdhSELN203RT8mlw3iP973AJ+J216yrexGFHqutHKRN7ZwyrbGwQR
xJcoGkr4mTymeLqG0XZbNH4fTKcMkwHrmWZrmqSU+KJSJFOjNgPYHvKfkRWP/zln
k+826p7gvPk2sRjM+fcfexzGXQ0lpsrladFWLcN7TZxm8tW5GY0V6rTudcehl8JQ
LhjZZeYoG6Dy7V80JCpsSCsjJLscRYv8/vc1eC4tWfdNMqMvbG5avhF8u2nfbFeo
TTe0MDGQEtlgYHsHg9jDFMdgljLabWRROaDFVa4MxADWrYIbeENjsB40hwaXq9Yz
mmiMlxjSQkMBYKohIRYN6XFN14gqFxQw+yHgX7jvelaBQTQQP27YZoj5T4z/2JcF
3brarNI776EXzNYROpViHQS3lwK3u7lLMbj9bCpdz6sA1BiWWDEDGpJMtCEXj+No
3BIsZV8knTCSWOsVSyaAon9ZoaCP1fRJRemv7V1tEsL0A56ptIL5sTGngDbzLRtF
9PflUXi6VOp8gGMHSrKbJ1UD7M8JSbPMhbL9b+f/oghs75ABpNtB/pezcyBrkPTx
tUA72Rv48CaLBlno/eOT2+wldtKkf+XEOtcfW33Av4NrgF1oX+2ZyT9/dvtNdG9q
R6e2OMbiT3UEYdRmVsNIVPACxreGP57yzeoH0Qj6w+hvtsJQrx26YFURQ0wn9aaj
Gz0KTyiqwfSjiJjuUexZmuoMyzrU+qOy4is9pzHzET8dAOwc7a0GHGLTw/j7rAon
mXhsN0llBH7dz4dswmsO2OrQ2wX5mUTO3f+I5fFGk9DndGydCRLGb/+XbuZU6pmY
CMeR59pKPKmnw8GOw5XycQQkgpJ8b542wnmWHw7+/yIxj54/DNxEYEL/cuSACY//
RdPLP2zeKLiEmYM0KgXGwxopZtfqGgax6vluJHGgnbYWqJc8KjteWVWiBfLrpxHz
Mt1biVDD37cRkSTXZfjZN22YnaVfljRnhjT/Upjo7QHCvod/6Ts+bmX+X7m60b9P
mfmXzjLbL8FifCQW+2CpIwfva41p78HJpo341X07lCeSK3xwvsQYk9q3ijTfuylx
07zwnkz1YtwJ+s6oU+TOIPrIofdbbAJj+hqklxFtWiFtHiM5Yr8gvXM7nbdZW4Hd
QDPyzDnixcrJSJAvHIwkhhuFfIk6/kDM5c251nBu45DZx0GnjMQWfWzNDwBHa4og
meZreBNL8NHxBShxvXOCHbUhKhmT+elRCJk93F0r0UrvjyUYXfoaGhe04ncwo1fR
edFniCBEQ9sT6vM3hbVhtdxWYqxrjavfVLLO0ofnLPIpkysuCx69p9RtVC2Svpjp
Y0xIzjYqwPaxsMlVXwa8PsZ+8+bvVn7r4SCMXL7r+mtm/RwUxZSMOXatL6k6KayK
C3ERHMeGbwgbGSUzGF0xBr32E744vHaBUzeF645j9Zb4cX31mYZLBOfILJeN/MTV
alNGIeisn7I0z31es/XlfKInYeSEOM4usfHh0a9TOS6SWhvOaBCQY6HLpK6A9Ksg
vm0EIL7LkMAQ0tjj3fREr8996pSszT4WfB++twdREgL1ub5k3Fy6spBSV4rNdhXQ
nP4EOlgz3waD6AdLjWL1+UGos3KXEo75vf/OqepLGOreCfOvFKGGB9iH8cgZChFG
W8yFS+TCo/i9eolaqbZ9NaEmXj9mLETkG6JOkJD0I874jEax4S/8tKR6S/fkGMbm
gM8bAVcd61ExVB9Q5YhrcYB3SWYj1wMYR03ukOPzujAXjDcPz+JA+lEmYWXCnlJz
bB06417aRv1xgcGivpuCwv/j2MuapjRBvb2+LF4EljcxPr3tQEm9Id4z2AhGCAHJ
8Wh59XqG8uV5YOTfn0oMxc88bDwo/1sw+j/FwTKqhNagA2pK/EQ/Tt92+OkSlWS+
7ldXFUJciJvSO1nxZCaFjzYknGvfSBPU+p3WNd2KKenGefLwSVdBzuJpRo4fE38c
K8N71A2dJfoJ81THHqwCvVdzl+3K/U7w9IdpHSohubmODfVPiAC5E40maf7pORAe
sZ6sJSvnx3HF/MUMB2z8RQWwAGEf2iZd9xxlhSYxKmPuH+A1pQgrbM7NtOBtSq29
QujuOCQ2jfVXxxGlJc3H7c8Ed+3C43sBE83QqE9rU7kM+fEjgsyK93T/HMv8ZnE8
UZVF3IRxFtHoM9o8z3gEuqracwNbbhGkw+41oGNeiP/u6mK182d1hP3WHPTUiSnM
xzU1HEspJ+iQ8IEHju/EpLeRuTLU+HSxOyQEaFdoDNVm6HjKKdeFNhQoJ2UM/ldS
CN/3lrwleJmXGk48MVQTucBeEpq26HshWpUsRQX6MVifyd8ngs9UHdi8WrtWT43m
vgFdgPE8sHU9/zapTDaKjnq48rYlA0ueU9h/xinzdcLc2XYJvIOYNRnuUnOk6tlJ
awO1XnzWex2RW2gXeNd5uIglCwSs6P2HjqmHASACzSnb/vILz3BhELSPc7i7T687
nWXot9w+VWhiyqz4bME0Q/uOZfNag4eU2Q2QudgyM5IZ9P1AEg+v3NNkCA7HQ10v
fROTCU6avWwk0gh8tlWTWaRLsxq0+nMZE2asQeiNDgWKHvj0X4HR+mPlS5y8zvmN
JVcXrWl9erDS1k7XANxNoWNArjmL3nmEk7GIys1/SleKGWV8oJmewThF+9LRp8QT
Y+VWV2cNr31sAbIminkSmOvIVX7SzzWIhuTlBGfgi/FVrjokPMAIc55Ue/Bi4Tca
D13EKO9Nx9ATdD7TifsVFr1dI6OoYCmWG7xzoYQMnFLMv8HCARI+g4jQfWRbolms
R5dkU1yYeR6uXDqbrKcgUWfitpuZiWiMSkRcpW6LIw0X7Z5Za5hEj8PT6u9GJ024
l0JKSWfwkBbeLRd+uIK07wLXwk/vSyXFaDny+xCfnubaisMZU+iEBN6WQIiO1z9n
oaSQR9WwnRv255yW+nujlOexYCQoZKzxHcqyIM8aQV32lZcyCHvX4BYWC2kEBfgN
LyAMSnpcnzDEZ/EA/Hh2bVNfJ00qtmjjnnkl3hSntkekRypZ6MN8gdzYRPomxIvT
IpwijgIq1wme+jneVhwMTUgs8UQPwKyChBSCVYrnhqrp5/aY+QE9NsciXWazlB5E
AnS9kD113c5C28o9kQE7u6LZCxQtAh+CauBLpwTF4Xq9rXP/IvrPFMtWNdioNkAF
Bb9hU0bXK0fWAZ+lgSil3HHIT1G1IhRsLphEudDEXahzreKf7OvJ5X9NXcchrfrL
UqocYb/WoRnEnd+9frl6DbsJgAyqVuUs+0WIuABurk9uNZttD8cTKVgetwAIcXIj
5h9jIJvyb77b+6jCciR6hIKtEpwdS5yt+pz8ep0i9QyLql1LjFEEo7anfN5BEFpU
Z5xv1GFm67ATV1oHURpKQMesvH3iZC91UPruEMDl4msQKTZz7Nd2TFlFfhnZEu12
IqP+sG0nycnnkpFS6n6gXerRp3tB7NSntUZMxsyRtUp3CxzBq3W5kSYWAMMCRwXU
LSMJLOxLQ5gryKo+r+EtABtKnqxlxxTkHPGfLPDpP+YCJm0Ha3h9+KLMDOcyNj/Z
b8+3abStxsE4Ggp7/Qi/Q6sTOut3AT06EMu7YP9Lqxr63PNGfF8I7DvztYfIMytC
YcfW1jGhLTINJHXWl8ryWJ2/ZY4JOb3K4wPCyuwKkrIcYfP/FS0pEN7DR+gclrDE
MbxzyXRao+fS/6LGCA/HNrxpy0aV+zhC/4Ee/2S3DhPApv667QiIWp438x64pYLp
ZcJThydQFfxSk6+0nng6fcRsGAit6dVnYLU9qmwo9wUYUJTiWy+OmYHuJJKn3DbF
0XlxQx52PL8ixBo22xWkQRUQ/XsasxlomZv5ggrggjRV3+lkkbY6jVE9rGbbHAou
5ARpX1FLqDLaA+IgAG0rz5L3fbsfgPVhNPdOrRlzM0TK2vVD5DnLVSEnjVK9FtWV
fJiMefbPGMfsqboSSM364KbYBYw8rb9+s+Cgdd1c3j2NKIctIstnEVOsTPgfwa8V
nUILUkVOQPTe4JFYhq6Ssjm09p6R8bKXqb2gmufkbW4whr7bF3GVASAK1tEIm/vD
zFcxbeACkREBNHoV1BJy52TgD2GeuRzgT5gCD7R/0ezmUS/GD5QctiKpCiaLtyru
XlkZC46G7DnnjuGi2nWU2TJK0BoI1ysOoZ4Tzunof3pis+oI6kA48Pt9ioDhsXJN
vvZb7XreSHZe9rTFrkCzKwaHeiuna1wHGNHDg8BfAIpSxa5mW5qLmc2iujfmS312
z+g0XYSZGWC5+D9LCDpZxDWDwf9Yp1XArOea6Ff6+nBaN4y/O4BlbdWZOOLf9fxA
sQd1uVBiF2539qq/187gNm0ldcdz1IGSmyGF7aAueb8hrAjeEA886XB57HHQtT5w
b7Gt44c0UDxKHOfbb/Ro/SB5Fcf0qhJl7eT5rtjnofVvVXdiG8Dkk6iA6aZdODOB
bZMzV7O61MrBw8XYblJnMNjchggspnJDRpid9gXyyZPSZ9FOf+7eui3sOBguekVT
iaBRvQSXKGsKJa+Qbxd3OcIFzTAqNMxauvvUVGVAqpcObe0LtzN9fKZ/8nWhCv3R
mrpOW1fy2hULaCqXwCMDcP7DC1CEmUlSScHO/0vBnX8tTCTPUE8zsq1tNRUkxtV1
uLAIapk6NDVThS5yAr1ZDPhVzQWIliQ0Mur5tdNKP68PXoVQGpvjb127EZxsSSC8
9bD4jwtMh8jnMTjzIjWVhXY9420E8UCsLZnKkmtPOUNmx8uU32zrHhcXT2WqufWF
QTh90HCuZUS6HhQXLTqTeMWL6tXWbP1TcwofKPx8EiGn3+rljUCYqvBj0orlB9Sv
jn6iq7h6PUJBZ80Nk74aO6DnysSrgB+B8MmUAvndsQuAKu18zgi64HMTmbNtrmXk
r9rrl/TBi194Kk2zbCV503HOiFZuKHLvCQZXzg4dZSLmvf14cwSjBsXty15z+acc
EDbGCwIAOpurCVoBLfCh5aYk7D3qaMJSNpZIpeGHWeXEK6irUv1r8/RXHIyW26iW
LH2UkJ3XndOgiGJPgEglkVuG5IL3KmLxeuGsCkiG89pfo3VR14neVrUb0prgrST+
x0fJ0QB3/HN8RDB2/KaIqQq0J9luSouDMSOwBExoYtrMLzuN80BUkuCEc15oh3TX
1+TbQPF8wGRQxzoWo6Avf+ZGcDEJV0yJCsbOF2bwWtYmXL3pihX7jjmHZpS9Q/Bq
UTmTV9BPuMTZfYS0xtoqdXSS5xHD4/mqqCgQySdy+6N+hPPuNiCijR1761NOWbEl
Z6VIUTV9w22TdVUDca1lrdaXADzeeRztdsJgGYmH6i4+42i5qs8rMmSlBJ/sdlxs
JzkXlqAJ1Fq/OgUXRHfKvSXzKxJXVDViQxOoe12t3lIZAr1rUIJFY7m4g0pMYi6z
z79u1zU3n5SdyposhRlofv5l8CSKy4WRA7kTytsQsfKchBAa1hb1C0B/X6/XeYTf
ALfcXBe3PV0+xk+9nYFKD0MtiEb66TEFp5noDUqRoNCTxtySzN/fTF8YywjyuD96
d7tBqaYgqifxwWr1Ebh1E+iXDLuTmgYhDUK3Y/U4XpAtPqfnHUajuhNJLn5MTdS2
M9dCwt95tYXoK5ym0f9iLXkiPesQZkbCteVqKmJ6TbGgZLJZv3rdZcakH/8Jh+aK
t3QZu36w92EXm5FYUmuMCjjm/yiaf/OGP2BOK9wnaM7P0156dyLYBND1IbOJh3Xh
kvGyvu/FeeQNWgmJ6rF6bB65govFLR5F33NM09TNUAxV/0SQ8O4x60Pmq0AIsQNM
4f13AhdempiUayx+HqpDdD3I50PFR+pxGMcj1cH8WehQ1HNmDiGnOcqT3l9jvllZ
7KVmr8lpj+lt6uv0HgArwmEw3Mw/AizElVRf6t7u+E1Bq8fHhFi8bUHUzBRZ4Tix
sQaQPA14N4Ae/gcg3095q6kGdOVv2KmnxC/VEnqbz2l8x561svK/OeM3MqSLcZSm
TN2mqkV3W3YUSv5QlJpIgo9NGOUzT9hyKJ7S3M/3CWa4M7pZnTHMH/fqqe2mAW9+
y5bvnsEwVN1Ba/p42RPHoNJvpgmtnQZkTiClsmpXVKj9a1A0zoARGOTeq+0REVKa
WgxWGowl8rXF8iYTpGzrX51186uqywxbmZ7v9VHChKUJC9hJpO9Um0ZxUZO7iH3k
fhstQbVwKnfLG9Zo4BJ84UVBrsdTKgjMBRpKKa84EunJ8ql2lV+1rvQRdFdn9QWb
AYk9Ebh7q5Nlxskhlcjmsq+WrQ5MJiQxNP1cM+zuNjyi5INd6LSNZiJd1RhJGfiG
FfEIUiVduNfIutKda0kaXLPJMmmc6HGtbQ6YnH4y/wLvssRpiOaORPJjIJKkoNzr
CkOfFDocbL5I17+oV/Eo6pDWEF04G7fP9NBCfU5r0/U7SemhWHg680DtRncRqhA9
MEij1GNdxzZOPdbFP36uNVGp7OmPyffk2fMSD54qFL4aD5oxZ2+R4IuLCMrljp2s
l19t6CtamW4+Jx/jAcihgvjob06bhWlDmYP6C59pUqctly3LsHU2qtSnaRSyxdUD
X9E9C4ddsyR1/nOsfT7cL1Fyf/f/OrGNYGPlt5lZeUw4LRkMgjNwLATpuNOtNSea
iC5dzYrtcAI6WCYj/BQxwTAtjimNRZGP/LMphdFxQ8uk9WLw90YZ4+GZ4hFfPuIp
Om9gRD1pD9UP69eGCxlrcMD9vrzSTef/Qqe/ni5o3tOAMfzXPYxHK6n+dcKXY7r8
BGsomMX5d6yIyykk8HjXz4xDRAw/7dNAX1gXMnzJmSLS6YiCHngfc3JlNjBPUpjt
2jrx1zNdBXqg9GWx5XHxxaamu4hTke3B84AnZeWgPRMizpf0+lEsbFGNOzRNTz8G
tBe/v/cZg3mzn9q9wtihO/a6/KgyXyyRvSrBgaaEHGjWfswvdg/zKs2QvfNrOR9P
vuMN3hRL8ncpq5QzAoAKKRzxdQo061uhgZyQ+N4dcrAhbq7MpHeqI6mfzFbK2x4D
SBf7Xu1hgaxLn3hn5ajAmZK6TgAKrDecG8asBfTDl3FuzLhFaGzxtagBgXXfexGT
UVVRGrH7sCa5mysJMgbf5T618spotf1URTjXeNp5phTClY0DluFgNGVqvKI0IJig
BRd4jgH7sdI/YgGM1XQ1B1PvyqZjVh+4hY1Y094KXYVyD3KIq7kUBEqHJBCBSdRu
LNdEP5y03ldAot+BFZ326FSfQwDYhS2SXsJM24JbpeTbh4VqndqwMrHBHJxRy8MK
q1gGEGRjD5MHgQdfNGpYzGTCDGGS1QPn3HVLnQZliZcsvda2F7irhWBM3joSLIcl
l6BfXzEN24KYJC5PrwU6/X9wtFLV1AzXR3BW5y36ZMHoqaCECnOAnM/1dVBPK2mo
2fojDWNhrIuU2GbqCQ9QOv+eLWhpmnVZy1h2vfKxZxVPTDtDEv4dUuPmyBOqcfow
lqxZ1pRk+WTYr3E9cXOURqVNwOM/cKG/Bf4dTBtannhnUI+fsT2xtt1L9qVEtuB/
jre8Offx692ZVFqavWd3UkYTAtZg/vzPIdEH2qAUSiR2CNi/0A3+VX/vkgVq2jj+
HbD5Ymna+uBLM5AdpybF2pe7fbTqZeu4hqh7flktmTBaPXkC+2jtP87NAZCoHUfT
yj51IEzDkhCIjy0KAPUJ2mLX0K08Da5mocQcfunhXh71DmACpzOGtEwmKQpz8SCO
VdQTWU4P1aXJosS7lm6VS4NaWLzcRt0YPi1zyfLNj2wEtTqjLA/BJsrnfNpBUuTS
9C71m1M0w6vNceAwhr+Rt3WlAzNBMgg1GTqC1coJYu/1MXV2J7Kta3zknEhOzvHy
TxeWs8aDQPhM8NcwA94Fy8Bxua8qNZCy4dJcg1LMr9TlA0ftX7aFr1XSAx5AJOQW
99vt9JwJhOByi2gR2VC81x3uuhZkchY+sCoDRXfRLJTI+yUUMOFRfVYUYLxvmm/Z
yxLustMnWt6N/UWa8EQDg7xaCldcMcOWqNXLVnLGZr796TgFe3ug/3rX79PXSecr
8/BvnqysX4GD3z1lyIGfEgUdwcm2Y1KvS/KSIJ9Kdi9lK9+9ea3x2QeGFRoJ0BJl
n+n6VLGvAnFlwi/ZulWHJjHP6luuq0lFZ4J9RLAswMg3s+J3PipPVjCvbGC6yEMV
bT7WMh4VV9m1TgImJS6Egpad2LJf23yfSDUqxic++bJ4U22Pdey+ezOqE+fi1qko
4p/OZc+FfA0tJA5FhrdQ4D92PjeGggyC7aLPUg+S0Mss2vZ/N7En2khTr8d7Hxk2
YfrEa7w8hCCk0EPdCBjPkr5S6B4EJDwb15b6KijpwAdD2qWeyUXn6kd+VEFSeiYI
SZUL1gjci0If6HU5Nb5jNOguWiAZgxGHbvv+TVop6CXrE+7HsRfYOrcK22vINZ2H
uCNEcU7BgpQxy/Ory2mXOdxczmEmKhxtUMgoti0blO/ZxdFvEsQuf/V4i0mgJ0m5
OqtrCL+dwuwFe0Pka/V3EMSKVVc0UvBA2bvVj3qHNbuuXJBdzy+izpCwHmJNNn0b
bgdANtpBcdul2SJx+BSuObXDQwjwR+TWCs0vDqfXK8K1JEYbQoDDL/fkfkXDtSXm
ySDXyF+J5aKKcqUDEOR//tXzOGtV5VlScOIRcgALnInEaKmAM4cGdRyKwQYNFOFM
V4QZ3RcBwEfE9tuMv3YwW1gx5Ps4NIBwSiEbrRFeMqZCRRShvRvPR5Mva9LoYnu9
J0mwRXZhC8eSWHC71ofztHalgTjFgKQYmtwDh5kxlfbKHDG620xumtZjPvIaUnIQ
z5kzi9lPgk49mhFndi8AK3yJcNmP8S4mgHYHetD0ZdMOSw9wZsMveWueXLsHYbpn
oQXvizY3JRlkBS8hZ/PnPsbLj6qZ1ILX8EKzXene8mygFIA0msgAEZcl9YAoyv1+
4aSdi8pbjLC8cniS8Bf8luXUFeJSi4LhwqPz004Z4uFbKNQp3xQsM9G8yf51XtPc
HZy/q4OrqN9pB9jhto/qIW2M8sktR2D55GFChlNXmZ+POY9OQf27eAgaHoj72heP
2I1bf3aBMVnCtdnW7i2VkNUCmXUywUAAUMK0k7WnKOUubfr5i8J2TowRtWb0T8UK
cXyrmakJdkP0xpepMa6cE0aQoNOE6ttQs7uLSHsPzYRXAbrO5bVBHwgp/mi0kJst
c+xx2Uk/w8qkyz15GiaN80QJr7fQc2GEXVfZkwHB9IoBxlw0F+sJ0fok4wFpZKVP
b5I5Ljc9sD8MyQlO8ZSfDOQnLbOQnlQ7cU916PT0DXrq1wzZKACdS3+etHZFxURm
NpgyWO1GTgC6PiUwf4nrLnRBEKKT/zBzwRftYmaoC/QeSnu4/3C9ZfNw8ReiKesy
cvp7yxwlulTDmYZu4NfAA5XagF6d5h4M4VSJI0Qmu/2Uq0kDC853dB1bdPAqOabw
vvPJyaf26Poy2OT9iDQo/NE6SZiS9adu9jGC4gplnBpF1JUBQPwHJMPr2VnJS0RX
GvwkZrYbzA5WxkDrZFiX/17zdUhZSSCLZ9cAb3RMroTRUgtE0ILNfQFdw49uTzws
awsr/bNAWN7M8ZNDAcaGZNztBfiZgu6kZir7laQCNzsYqfekx8VO0j8ObBYw7rMF
/I4Kb5ka4vLv9MLuOf1x7U/qqB4bJxGtEWrHjEUDqEcmPZAezDt9Zr8ywgWV711X
7T3fFOh9F0QxHQyCeHdh+U7jExz4m1ovkP+TEWdqLbXaqMyWxe7lnuuvH6Q9QyVQ
SnDqU+uxup5ld00m59/crr6mhf61zXmV2oNVvet9IrGrIyiqnSw8Gxlvz5GHYw76
VuQfvl+hF2rfEvdQbX14+PMvYrztyhUFE17I4Ah/1tnWZJvjUO1YFAUcKW3nIJqK
H3Zy5NPi9hbFce9Un59xBK4jDmNGWZJr93Ud4ijr8QRb7vaascWkbTs0fHg1yT9C
vya5pBu36TCUIFuVAOWTZUTr6LEs7b34a7Ek9aWqx1gct9X/n5pRTpOgG2N6Fafg
8Kg/SelRDhbgCzpnAkIBgwoaD37Cq/omTYm8wlE9hbU09u+VGwNfpMDFQ+T2jPXT
wFPGk+F/yyWtxnHsn+pJhoJ1xfVop/6rs0jlEbtC5m98AYM2kzc3Ocgw3CyFdC24
oDoHTmUz3gF16hj0wf3iAnILkPsFFPNvW6q9QaT1zzJ5xEra/mOwgzLmy7dVoLVP
x/h3OCdRwen2lo21sIgn4Pf2ay6rFztSQiID7HLH7Nnd7oBZF7lvHCMDRn+88ls8
AM9Mdf2y7oLb6/yn56dFdnA0SXGXd5Dnx6BvhXlSAbqjhq93qCovPLPsL1UhQofr
O/1Y6W/M8F/fmpOaQ5sys2slilHxYm/0XqbvFx2qMi2+AQgvs8FqHrDMUIP6nRce
PJl14pfChh6QE3SFR8QbdbrAb76C9paTuYYg63qfJa51A8FpsPpaV1K1kHwgxdGw
m5Mn2xJ3+ZxKUWmSI3KxoTbYLWQFh9Qwtv5BnT/MzDGyuyUEIxBnOJlAxQlA0L7V
8thC8Bam3JvMYYbGFsSWLb5XAdaLE8dM0K4G+agM+GSWZOWuzWBuetPjeyEeSyxc
YnsQ3XZIUPxP0qws06uWVeSyO6mhG7WfZ3Bkwd/nkUuFs+/fdP/I32mSUaR1h1Zk
pvcb5+TvG+SaJY+NLElu850w+BiIhL1Iz3c6+ywiTDuYrANyilKSY34jYR3lQlQm
G37dbitpU4eWhlh9pRz5uCbnGJNdlHAjAj7lGu5NN3MWkn6wVy2T2otzlhYoxrlb
x8Rz3dpciA1bWLN7+Aw/CCRzvhblPhYve1oibCAvXSLxSdNzKgk7p2aE/8XVUWU1
hjHUy7c59lbCTlqIRsuOWqHno1dEm4DIgqlINdi9OacWAQUqw511lKtvAMu9k2dv
J4fj8NXMu8A5+h87nA5G9QkE7haHB9750b+Abbo5v8THpqmtSGpMFBPEcx+H2CTv
ZQXZ1i+1J6FTgCeiDD7gO36k8IbvzNZ2mZwQiLFKiA9yjAAtg7AhrmSjk1DmPyMj
bzOvFMInkyGZtconuQWwg1ueQpvo1qWWEl7PkQdnIMFvzqkAo+YoncIEqm1Pyzww
oIOXBOgGQSZMdF9HL0tGMOsMQnQf3lz8ellgz4J/jPPXm3orkwAtlw3Hij5bmifO
D4+W+W8ogDKsce62s/6iQmd8MbXLIFbmw5k23up18lGTNn62/dtLDQ8RdtLOtRJw
c+3eeb+W0MPEIMHB/fCqljxz9lEylAWZEVuWhxUzD3Rx9rlqTgr5kAG6mtCBYOl+
kYrXRe9wiUtU654QKbpBMd9BNZNTJqz3tP7v030Sce2xcAJq4Zl5jYQQ1UKmwX7s
e5N3QdWxEyRB4Syt/OQoBjbzR3KUG+nm3nMO/qvtoFPwNXcNCA0w0PpOh3i1Zp4X
i9Ff7rC92jLMPweF+2eMyaNxFRFg3P6GP20Uo13ckmgvyyNR4OZ+H91DwJKFSJb0
rA284Q6Z6gYZntsp4gFtpW4NtwodZQ6eWRTSosb1LswgQrabAE9nkKpD13/tIlKb
MtttYps8FbQbp7r10Uzu8vgmuRKeVH1qIuwUONEPksNs9Ijod7GU91afj5XXiGGb
awPo4/FVOCZVmFOiQyJ8XjCAhJ8WFbvxBcrscBkqezlz5j4e2UkK7/DO3o9kntep
Gl3g7/0a4CTtNDWDYLZ97n7f2HGIom5bjFgqxd+4EtZV7TbotZ+zDxBFaKwi26c7
jJySvmFuhyRPIUf9OW/OHNEIVwHhNEAhHunpPZvpveFSaxyvJ4i3IEIewOKoNbI/
0QvjTqgD/JZk2JyhRe9lPJOyirgvjsqA7GRJmz23GHgQYyQlX+ZSIzDdLZux/Ml7
87m8Sjyb8uq3yE0lnmUqCqO4EhFp3SejzpR6uZrLzpYN3i/CT2HdzWmYg1ltf/Gf
NgH8/LvZgCFrawEbt6Kbhzl8vDO0TygeHgw7M7jGSjBnDBPX2OBUg4PdB5b7MRZA
PmcK0kAD2pK880MD3H0wZQhds9GhXw7nTMqQ8BZ4V9Fk4DBGWMJr/j1qnlBtRCDm
6KTUVMV33koe/jdX/b03IebkFZyU3la+8WtnUXPT6vCeAurnuu7F8hpG2hMBBkFJ
Ccawx57EMjUzG5cPR24TTBoRPiM/O7npRUQmPNzD9wIWmo2v/y616O5Bg2GKVd0g
3tW3W4s3UWcUTM390DSaO4eBQc4hmFeiP/JmJq9Rlz11BcpwBnhBScbMUwFjy3Oi
SoQj/mmfthEGvzoKaiBZTv2+4OQUTPVfzlgZ31Wuhn/AltjHzKqzBUz6xudqGzVW
1po5FgtdXVx2p06diz0idBlwZJX/VQycDgbx24+dhV6C0eWrJfa3V9SeKnOcTfdb
SjKF0MuqtKtTLEeYxbpjZV0XgyzhMdUzn7qevRFCNxOoAgkXsRW3ZsGKgVZgead2
AkHNTOK6tnaimfoxAHYeuSqIlxc/YX9a2PJDOYsUqNKAJeNN8xnBglIOaqxpHdxY
8AIPyF+j0dMJzpL0tY0tYh01eHmKaKfPUB9EcnluokeTzwwP60cG+lHbtDK8lVTd
EyESwthgKj2ZDzl6k7BT6zZZSQi9wF6sG3qAVSYyavQCtHnJ8bLShFDWOxlUNg0l
7U/Xlh2ppCEl04QH+SA3SptBaI8prfCsRrZ7cX5cdy/F+hkHhL18W1YKt83G0vMW
eZdX2myz6fX4stzo1SeSllOAx2nF+HQGbOKF91jAfj+oUQlZ4URkiWayNzmAV/wJ
gLh7C+Knaaamw4vTGMMS+xMdAvqfV/CfuxjPwUHI6ZIvl265VTwXOXneKAptmz/1
HYuTJEhvCbISOM7MdPV2KNWQEyOlb5uiHIDujjnllknAnAbdmNcQSIaPPlE0SgSL
SO8wqq9NOunDk7dVllCyFNH/SVm8tqtcli+sikJ7rlOg0Mr0GS7byMJ26RPdYMDT
ybfm0KvBtqtuR/x+pjTfaGurgmveNjD9+pDQF72p+kcC/YnMFtSzJNrX45a5VuLi
UYrV4oLoMvaPm8OMsekYTrZ5i61yMttIJumWJJv9WwL68u1MVYcZs3hKfKPLLoMU
urC7Bm8La4qPLMwrik9asaDcCHoJBEf8MpLBtYQgcCXad8gdVbV6kEi+wpr7+LCa
dMCTps7/p6H5yS4NbtHxaDmmeg6UZooJNrw1Mf2fUifxjF8OFimAwcsTX63ZyxZm
r0ZtDzxeAhNJ2Nc+2j58rZww3gIP3ljefiZEHZRnlOZveG988xv+MS6sot2u8dVj
q/tg+o33DqiYLABY0sQHb/VXy/CHi+0+OCAV5HeiLQJW4VWPKD+QRfQfTzyckAhp
2YYJ7lNW/leKqzHeyafI7r3Ocj2P71ia4x8gEBvoUKP/KFq0WVMJ5SKlB7HB6EiT
OZENsrFg57xEBh/cYV9Bz+oaxU2ow5nTo9/P2LRjHGK2bNnfGGe8FpAuO0QYD7OJ
ZlTFs60BZtEvu5ftMKjx+aOmq9DXc0B3dppo0jHd4yOq6aY8raPxZaPfroJDjonu
1r06Z/VZYnOd4l4qKfrZswOlf/FBU2gi68vW1IBU7/4NYSo0pyJkpiSauiE73L3N
efhsRWnWTNaUSjbOEsPUrLWksj/FaC/VcSBQBaaQyFdfn2cWv6BWEEcAhTO8454t
InlHlJmdFXQPgGoeVrA/SKluRpVZQUZucY0zkIkt7x5jrROWo+nPBUIl9RfQfh0M
neqQsR1gxoVtBj4+p/RzCz3JHOBxqL0GygLyJqSKLIyBJkqncR1Vblz9S2JpNrzy
X5QMPTpa7FyaQNi2dzwlvRVXKsQdeV3PgwunyjS8bzj/yGx3P5qBFNv6ghi7iL2W
WKYbPuyuQSoeSCXG3e/vjygvcFgVZJii3Vz1yFtr+oGBft2bCXqYHODufHl43e1N
sV/FV+mjAhv0K9C/qVxiJzeXxzMFaaAZXKxLoV1yok1jlzvcibt6q18PXMUTzYX3
kPWIxL/jPSyk6TEaxDvEGxDaLkFFpubPMkIUurM+IyKo5Qc2Sk7ttLm4EoEdR3Q7
W3cGpiw5RGUrINIeTse2k/CYgEAsYjLgk2iqo+JickNjZ06ysaS3bfDotOb8As+U
Lxs1GnuPAg+uHAFA6zxe+LpJoEBKhgSvn/AgerMxRvfBz6w+nO/4Vsi3QcEvSTFx
x7Y5s/PQcsOZfcWXBCOhP4K/4c1f536Fn0iL7JuvQ+eEXmCvMZOoZMs0V3f82hhx
c4vg4wt3xypr/q5B/MjR2T9jd3VcsKCs7vkDN4d0reKe0TU0qLZWgX/bNVWPb+cZ
T9eno1juJvj8dsvqU1I6Txw2iKINDgERJUKmDB1d+skXC9zqqMbX59sz6NDWTEDd
+WO0PQAiGtZ0sI0K3dP2amaJLMtRSTANW0HzLQewu+HrcrVT5gRq2HmOR6PMn/GF
4GRdOTL4I1MVu/mItbUdetzX0QeTK0vJ1XZubmijpNXqaJ943NWFehaUCVfbYhOE
OzTKm+YKnMjcxkLV/uFViKrY52kiskiNW8MI6VvB3sj4HeOgdoctqHa5NsV74Fug
q3dHwTKf0RMJBgUNpk5LH7E2WIgEX8Xf/pjXIT1x5iFGH2R/3IYGqfBHvkcXyzZg
jscxpkd6lkRXQmWupP4EtLXn2a+gGLid67ZRLDKAZ7vq2EQd0oe8SuVqmmAcSTc4
oT3LMq7lBxSifl2YT1Vd8pZqGSsfr9BppZZm5YhfTvvnQeeZvKGC5xvb82KBd/Mg
+ezosxuLhsnP/ZjVTtr9q/f7W47kOY05mMNvSZQ7k4JQBEvYW4nCyZZb4Xs4xt46
z8+2J+jcgEQl2loXOGuA0ZDP06o5PnROvtsa3iAhbnJ/2GToSbERDRBSexTqC4g2
pU6tO/685/gikp37wlMZQGO0sIiN1Sxz2Y6VnEis9g2DoU0RSNMXVOXxW21NSwtB
iTA2qNTucLvPD4NE5JkyF1yTtfDnnOTNrSVrmDDon0tAMCjcmV64Uj3UAW2pxDUo
IEvRonLz8P1wTnkb7KU89ih9m7wfdJBrFuu8rHCSov45yQMTJCfXI8FpcWy0LCQi
ftPS1DVVJ+FUlUD9YcEJ1CUrZk6Ls1l73IDkPqs2OK8pzz3+Y3wZYDyjIoUuWsRL
zUqfH98Iq8vB4MHbXulF/REGps7Evjgj9Ak2xfwIhXeCmbbyJ8qT9DHSkWzsbLit
8uH4XVBSSZDPUZUEJsZPX14yJ7NjNHDmMhHaFiM+eu0R1pc3oL6eeLGUydv2T9j9
EF3EVeNDgWarxry9uUx8lEwJ4Ggl61MPUBY7m8YGlJRiTyUcYJk6t6/cz7gDmjO6
j642frBU3fODfzJhgiEEL/ewpd5SvSIUHSK8J8455TF3K6WPjyRNpwPj2k0Q8v4p
t7WU7GAzcP23SLsCmuKuwzq2859YexOv8pqW/WhxGuTsnXM6nd0g6GrUOKMuMQ3u
zNepyIF867fx35Qg+jY8Xx0ygNF+3OGTdADOL7PAI6lnMB+Qz+BLo4P2Cn7xabA7
AY6yz2RWFJTuOR5ckIv9+yBwWIvVYb0bz/Ej2GDnItYCMBifw3EX1UgtYLAHH4Au
Q0/t893T0ERya0qVKqSbj0xzor2/uGRMXofbQ+q/cY8S/dDBmMK2FI5ho83LtRe7
t5K9jVAApHoKdIy4flo4TukOaGKDlucf15sCDz5MSfQWevF1YG2fqOk5uj5+LEnC
HD2eIQuFdccEwUmE/I8HBQSBaX875Q7/ili0VkbSbJbFBfBxet/hLf+RBtlOnEGc
CiaAyXJuEoqLRswxTP0R6rL0sg0NFFCCBGefQDQYx/OIs5ihuNe09c4oOpXT06Tl
mYhJUBMPWbNGgB83K8a+K6V6MHSsZc1Ak2Y8bsUa1iDhJerLlH/9x4hItbqKf0kN
/hriCLowc4k2gcHC5ZurdA0+dPDOiC6OgqFNtur7pDO0ruRcIGCt+XiCMMohaqtn
A7szQs8sFPWB3/QBMcAKfOIweleA16AjVssL6SagdXahuODGVxQErCvfK7+G3X7F
Vv/xUtuczBtM8yK+7vGjtv7P92dJkflY5Mw/e5V4637qmXzED/XqkZVB3uPmyzuO
5v5OTtSA84R8cTaRfdFYHNuOfpv2t0uLuxIQvTtUvQ3ZknuRswUMMcP8miVtP1Jd
npFVYVKrueOuUubvV8EETJcIzG7nA75fNkqaQF0U7pltU8ksqFALWWB0Ti4TgMy0
su2vwPCRzANe+9zZ0mBuZLqAm7rwH7G2AZOi12aZlXdBEtWuQij2ziDF9aV+DVte
642g89Dp29BtBVxB3STMUZY67Zz3CFVi+zL4JDyCG60HALFsl5XF1OLswco98hD4
29WiDXJlD89GEkq9gVtGvuwUmOedjDGPdCH/OTSt3D3534mcG+Ai0K+4DfqmT+yF
NN5lLZchITDmgSwoAwAWB4EGxlZrk1BQ5vjs3bJw0O1Yi5R1foXMADWV7YyNNufh
9n0e4Tc5xsYS7aPiOXT//pxp6GvfPuGOg7dA9yKk9I3M++hsucgTTvJVK3bv1I0o
tRlVWwK8elFTcTx9udVvHhjz15UAUpBevf8VOY8fS/Z4eYldP20F4ojNo6MQ5GQL
v9JSr8ExDHVhy0I1mcT2hvd2G69wi95cjudqSPJxxla2IzUrTWPM4bej0rj5DZtF
PPWFb1+7NGRjzqwHzqmU574gCrPGoc99JOdgT/F+vKcfDZPpRYKXmQO4JAeHDov1
5YnvuvzBT7RUxTPRdTIAooFokcb1o2RinNMJu2XUDQwQ5P7FcNaulzUAov/qQ33c
H0fOILq6YZYFzbLn/OL1uz336ZRbebs1Az7vDkuMP9WxMOrK916e9J5k6U7/aCzm
HTpH0O84yCp1PzTL5/MxBu59r/5DH464gt5bDyIQcxlG3fM2qna3W/HyabVP7mkp
CorEBnpAHzZxxpy9Aum+RXhgW24c3QcRQZlEreJ1Wufy2mlvn5WLoq4ju7oZApWy
6dKfhn2Wcjb22rL7scL/t/I5PNJJ3TTE4zbzqkbLm4k6+qITf9cnIDJbGwkqOAki
gJQNVAPeUau5tFKhrSD2k6yptevIsGUVu7PT38oz7aHMdxHfZCjmHiNIPBJD5iby
YB/f6B1ESrDt50if/goJBks8cGno4ZbFsbPfKNwY2c7W6O5wJDcaK7W4Jmhgz1XU
D2C6HhQA9s/srzXheQA0S8Zc6YatX4Wf5761QF8K69BN9rG4qa4Jm/cBjHDg0YNa
K5nnP9KbZilSQx8F8K9rtvcXZBkjuGqvvKofjmjihV7WJvFcw8GjP+fjUkj36l1T
azzPL4pFVVZR+sqzIS59uzmULW4AkkcoR+zJzynv3V4mdMibsYFP456vyntGoMfZ
NgMAxCUWkn8U29kmPQqad5Gth3mwA4ipzU04YzjQ/pZa8Xj0R3/UZ1ZiaiT52W1H
ymrmU9vbXBpbrAw7K3Vm0BPZo/IN0huV67BuZzN+Ni21mhUNj8v2JNgOU1sMCDuG
THOglvz0L2xldweG1MDfN9U/haoGs4McPGLLxvGKPwFDMH1wfERziS+sJMKB7hON
pYDaah1oO55b3wk9eHymgKYmfIjDMz5DJoqUuKSKE1WEYQviSiZdUBIfnFzMQgn+
yCg7sHscAmY6D2ustHhRCAQwzrrDXqUGW+Cljok4cvgP9FRwx6JNroBnj643LxIv
zlvHj+nijEp9xf/MA67ZY9G+wi7mCSKGlcmcKloHaKZHl3TDvKZsfq6zvOkXwL62
BBzADMrLyKCyad/Sj92xCYuKGV9hsD/tIYy6ycJNCXzrDU77+ZHatB6jvBrd+SXr
lcSS57bQT7hb13R8MZISTnqdnN8oXW2PN8Cwjme/D9o8XKTN782lS3JpY5KOfDsz
bwRLP/NWXC6oPBYHk6NuYMEYpK4FlxnHbnAMT9BpIOqI0ZnTVt11TQxcdaFDxVfq
Qs6F238MUWgxqP6j/32iYjxb1rFLL28/nkOLZS5d9wgnY7lElOxbLtmbtwSmF0cl
GYSatuodkQIz/VgAG/q/+dD0eGxC2hAraNsFsBxI/S4VJUoRUVocZrw9wfKU/bsy
POkZTozDCP1mf6Q1dj5VEyzITHSyNjQLssPDhj6f7vwQ+tU17SiuIjHNmi+BkZNY
yCyCDk8yb4A40l1ggaZUIKOiUlgBU4FfkNUPfFjHL2aN3KkY/Umq9ywPQnXZweC/
1qvZrBzQPhQsuTwJw+sClg6NwXHGgzlAGUhgdlpcncRlSPii/O9wR+TWQ/rj3kSn
iiX/9F3hVY9/dxSiB1dnT5BAWEKcLP0+8xXHxXQZijL+IBDpXcDeOctdiZz4wAGR
Jmx+MveWRoYUhaNY+xaG/IzBHebx0V9ykOt/XlZ3PpyGo3mJSvu6Qks2YTGLc7k7
iNdObtw78+wX3ySHkJi188rbsj6t2GAssFdq4ku0XyxEXHAegHrfc+y+y2PPUer2
npnchf+ISDOtFUCGbiOjW14NI89Ocquo7dtbTV6+Knm2D2dEwq52WoatpJsIUYSD
snvHyk+PFl6UDbrio/H0cpGCar+ik1YPS+fJbQVF94H5bnHOsPW1RZK5IWFGEntv
S7nJ/LwnUDOf64shpPAi7W/OqjA0gV7lBEpvR1e4xyJr+a1YRh9kY7a6nG6eEaWI
6lhVVoG3lotPfQPKr6IEB+gD/AbrCeKYHThavpnNYLzdJN7koJm4E5++3AY4JJAf
mEnepWXVuDrkb7UiYU5MBkLRMeom1lUnTCvuuJFY7X3lWt//IUcGJAoB4YTwC7Ap
Z0WHTjQOSh4rXuLBq6bd7lrdGNK5Wipe2dJJqK2dHb6D4uOExTKzOVpGjbr0APwQ
1wlzTvBqWbzcZTEoeiq4Ew23QHGCmjRwnFCtOMjE6dBAPBlgOmP2ZuZAmhvlcBHl
s5T9KJVC7C55+bV52EqvXcsLVfxkwWITJm4997GpmE/vg6Zi8bW+qLDegc5zYwk8
OQUTv8TrATIICqXdEV+sJ0s6gLD1nvwF5Cip20mD7LbK+GxxY0JVYO6yOP6G6PQD
gunA2qLTPyv9Q56PCcnf3a4yErBPO5jYkB4Lf8+yXSgUyCTtY5v9rds0YzYAkXNX
DfxD/1nLcRqbIKLaI86ye13bjZJul0OcMaPTgB9l6gVkSWuJcla+tyUqYKrosnvx
frxsr1ylbnkjTkiCB17hemG51o3IsjdUBvtc1hp5Jv9gr5PktiqJVGLStpRUAKzj
lGyMF+jvpqpwonB0z2XFWRpZptKNcNn5KjRzUqZwide4JWmCEdKbOMSAWtGXbVha
L9IICMwK7Nv0XlgsY5cH+oEt4YaFBiNLpGqdYsXbdjMVRSfrDVWaLKRO5i6lUaxS
s5OTzoPUtc5zQHMxwVL1OYOuNosvnt/nUQpF7nU0ruSR+dfH9daFezvt8vDkF58F
fVVMMdDMxgdwReS05eXMlic8WCgrPseJLTCvm5NJ6appKSLRClRyoMgqXYdQLFjz
G6t5+3kIezmtgIMiqC9WT9B77DCX/P8LLrkMMORep4Rg8JI7q53OPMoWwpV1wIkx
1Ir/sGLjbfwqp31FGqMOjz380on02GdH5jK6Fuv60n6LYGWNqr+aStROhWEYoJ3U
AXrfJrN4busIV9MB8gX7Zk5I48q61jq2hcGiyMwT1H91XFVBR440x+Qh60V2eT4B
NhPSxSdesu/N9huwTNPAIvmOjBa8nu1lq3PnVo8If6j3u05OVxu1E3AEQGScOHXp
+lQG2PQ+xBSVj8cfru2C1y1KB/f4/OpQ+MwbCp5tjJt2CPveIaYp0W6f8rOMJ1iu
w/Nn3xD/+z4dArwChPtt8nE7dCN7B62BPbxLgl/ECbmniZBgA79PLSJ8cgJYQseE
TVHWFFed13PO0U6mZtJu7yH0JKKHxmWJKlP4rIFceVoKhCKfuLfbho9EpN+18Jpc
akzgiaf1SUq2RYqxQOQrO0LiYGQBhVPRi1wwh/UG8qp7aIc0Gbw9xRw2OL+UPX1p
WER6iYETleXCWAgi0BBWN+F4KzGa0pnjeg+tx7RBPxnmYnwgRXcuQyREbEIUCwQh
6XeUcCzBVqWtrJNaNduuhW6vD+Fyt+aUzpJHkDN/UCs1IMaxrf0vL2ddjD+oG8MY
zccY6XqmpQMDmyZD+jUr9JUQG0mcspj7lsfQ7DCWnUMgI5JaDCmw8Er5WlQ4yhyT
sjKRJXrawL+MIme6EdUFtalz3efpXSvTzFbCmy2yB4hyOdUVRoDQEhjc1WMAC98U
1WlOit3VKBkZ76VK8USzSDuGMUCJ33aRvTvDRQrDv759VmgQUqJY1d3ver43eVXa
O0zOyLlQYKsTFzHnJIZMW4FYUnzISF/08P5FKOnzmV6vfaP3yYipXtlvbYQR/r4v
c3XTdDr8g8nIV653CI/CgS3otWjYGevI8V0LN3h1tMqvBpcIwkO1Sk9kO87KfXtY
s2EgUqC+uXUPZ8arOoNrqMYsMbxMo+t3CrRKyBqfyy+TYpOcjmCdFgcsLFzYQdN/
plAn0Aravik0mZ8teXzq0QF3Eh3urTNbpKAoIPH6d8PzbhlEFYGAP1X9iNek49C+
IXFcqGgR2o+ImklmVMme1jm4lii9zivQAIs/YlHO+7NFsS+leiW/B/bUQYxFzxKY
jJzAyBHMw80KTIiKYHKrR744vPY0tk6b3tKcYhMV1OOLcxosfdmTYbFvKwX6Wq+K
Q/o0xZ+A2gERojygRcPT3JB7YhL88Ur4ykYygAs0DJSoN2sJpTcqyPQeGB/jjNLc
864kLQP3gWIlxM3otweiCngC3zl/Msc0qjJHzu1Jrz7gfjoyUxWG/GZDzDV52yWF
wEek+Bo+Tlt2nWmMF38FexdPIASih+1IZosfhdLcoCEI+EkI82H0t83k0iZtUgly
fhCz5j5NrChDYtkIsRJxPuczDa0eAX92XG/D8toKQfac4i2kwKrsg3cFWTcHSn/q
/gotlmrc1GvgeMfiYtbM8wjT5mSK89wtJA7pWun5M4zlW+NnwGihYLDoLERPWXlB
VF9BgULJ+OCg5Jg+AI2n/BrBgd4CuATyoIqyI3vCVGVzp873AIR5O3HyM1rRfZ6F
Ktrf3tptw6Gtw+i+uMPfWACiDS/xgKO3EGwiUY7CS6/pHBC0K87ayizGXHrIsLPk
1KMCadjYo9hs+gb1gq/tGCiTeksutYY31XH9uFgKh4ChoGUF6S8PYAa/myPP7o9+
unOhAw4Te66JDxw9Vt9rssGEvowEjhNPDAhImHUlSXoWeKLb/v++6mMRjW234dxa
e+SjmnCxWGxvsXW2i2cSyFqxdX/3vQYKBG9rhuMRBmD2wXWwcMbll8K+FJX/FSoy
GmPSRUbMJLpnWxprSkjx1tRh4qcsLr8LB8Ghtr6hTYPoBZOfdEJ+YEpZr7uiMInp
0Wrq4xTDNYmLWIfriRVxtacFS6T9Hg27XckszRXZi1YdJMMG2/1lLE1Pg+/BosOh
x9jrjs11JhpQE3BrpGBa56krlHzHj8xRgv3193WCnMVtZmLsVt3AU3UrgAImaT20
+lOnNLh26+fvSXJCf9dODy7zmDxf8IsF7rcVG9i2oKmty7zV4PB39IVogEwL67oU
5dUepzPdyRMoCBHgnb8wapnSH2cPIcfPitHNgE6BKqBC1wBp1k5NjWw4i96K9OMY
yPNUhY5+AIDtIJtpoQVOrhC2YGXsAJDZ8+ZBGXZIqoxXaBbM5qaCcwjOZYdajmx0
ULX7WC1kFVdL0JgIt0CUQgmxhBIypIh3hEvQjIv51+9ttz90DUge9gpAmkVxBGbl
PrEryGZGXQT0hrdFjLivX7QLOiznDXIz3H5LUXtcVOPdbWv0jgJ3cNH4ijWtrz6Q
cjRme7KUNsWXxQnh82grdWaFRDCbpggr8eCz12aTzc13/d8k6s3pzJY7u8kfsToe
zmLaJVEOC2CzrxEyRjD4qqhbryLprMIJc56YsJ5fcskUsCHBJ59wG42EVkLTHzzv
0QiQz+4sw1hiYJgL0hpI534eopA5EBY8oN7bRUPlM3XO6IDw8TKBDfAwMIc4vhf0
IwznBtmKQnfkv1nzf3dp77LLwnCYDdw5h4ES02f15pxEkWpifRaK2GLj/XLSQdHh
6f4fTxvd5Qq+5Rc+MeguvH5kRE2abuKbfBrDxty+pQiZ4O+xjmTsq+iG6QjxPYyN
uhOma5J2MznL9iiaBKq3SFBTQGvM2sGouGoM7BJVqlNg/GGgTC/nOnA9CGXt9kHs
MlbSDfKc+p4QHRTHgqo1XMQlncEzfkf+ndlHBvHeYSlWh7Y+YOlxpxuVJQs3xDUA
aGjxM/NgjmYF9cePtllyZ+Ax55HEmslLvsvhFuxWr9mmCPuLRrtUhut2Dvn7JjkF
Bs2O8QTd61KnsenbJQUrOvWmKNG0yp9q5A77JM0wWaRZcbNXRmOHDHrcADn3wXpo
XBGk/ORJlqVeu8yRUtc6ScIjEcq+bsaVC2HSFBUgW0JTPUx9lvUGCaCFuE/thu6O
jvL6dAyIDmd7ndpkK8og/Wj6IPuL/nUY5L7CQQMNXuc13VzhpGR54byUqeyjoqXo
6YsQkfCEsgJd0Ap1hzlBTc+LKYg0FXd3aYXnI3a35b3My+DnQgmhhBRQwOqClXJK
0sANFsrPFwut4RyboQNas+PsFDbIxQ5Gr6vuoi+hVK+/WiCxj2JKgQKTSArEy6/n
LwEZHIl/lZHifslaSfjyoZe1R7po07JOYF5NhV3YVAhPicZ/xIQl9n4A8XsH7UXV
Rpv9WLhK8IwQh3snhtQbrVLyHWrBFENsT532cB4bYRIuOcjBnwoyxQ3fj41EDZwD
oag5QtpPjQodfdjE3A4xUcjD/b6/XjRzmKXLyycmOO6OXfFdoAoTJpE8NpRAdcEU
2DBAb2GNsen1m90Gsa4Lso+hnyQQFPT5nkwrCCT0qimRJnUL3gJWzc14W2z9lIsu
HD2ah3Id3tPkfCB3/hqhck8ZVbWOSHrT7f7/MKnAbNqm3Xy1WAnSjpKgd7pS6Q14
+v90I8lqnZ7ISFGGIdWVIYsrzb3Dwskup1P2w6hU+WCzaxTlX5ctp8ZmmbNfFBTY
im8Bm/PYVNZUodwxXAhm3x9hMzwLmR9iQV0rtOVQLcInPew/jvI25e79ch8aDLuA
aORnRbxqMtvD6zZCrwgBzXrbj/bvBYLyhRd3iU/rttygm6eLvZ5Kj2UgLJlP52RY
sljbA9M3f53PyzUc/FqZr+SCxvLOu8dAnOA5lSr/javrZ+FfnKJ90Sl+q+FthEIh
kAzc/P9JGk6fNGfy07XmgzVrRS5ZWtcN67f9dvD9YxtkipjK4ZMRt17ELvFajjK+
BPXym9vqE6I391VpaU/774x8rQhQbc77f2utPL1tnM6haLNZrIfzj8b1v1P14PqC
WqBqR4t/8ZncUKBLdLw0LnwDRpGLzqnpwWAEkcpB2k1dEWbnIigdEcfmy3iYIS0Z
pPCmn600cBNv0nW1GUo16YAzwlVlADARI2KmRfOdJMqHIThE3Wye28/dMUpH2s0S
DYAdnxc8CzxP/i/zaWzHfoBuAVGr0tfYRhYHGda7233WGBcfeHB5MCj9qKt83t1c
ysAzbx93TYDCDE6J6OYanzd40vShAYPYjas71VXhY7dERatMSQlM/nvQ6r4Gb2xg
3nb82Za8D8PAlyvmcTpIo5z7vZpqmuMb9qj9N6BcfEo17JH3tl9Ue6ytvNnALou2
UJWBTdEZylZWH8C2qhL8PgGRnHP3kx9I+O0k2Mg69xgJVbz6lRVK2gov5jG0fkDi
B3FDpQ06dLH8pu88SwrEJJlULVEAyALhOvXznXPAMaLJq8NoybSkPKxJs6ze6Fft
mBgEGjNj/SVEOf5i2hZPEctZqJ+Mrx+aLxRtc4oXUcbQIq0q1+YnRnsJnussDr8f
r0V6hGKO3+rotP3zzCkw0O2KA+iwzC9lCqdWkT3hWs/lwQG2H0jmCucyYOeCv/u/
9MbPrc/E903vV+GiHS1kd/8+uPUjM7CwvdJGKhcQGH6ClW98zPT5fg0hlDW8PcnD
kGbWpfzM9KLAI7SzRx5iL7bsY0XtZ/WTf2HRGcE1eND112okhIc/vtzJPk03AHNr
eV8I9bk+BjA7n4DCn+dZWMeRlE3HWp9aQ5G4RTHtqch13xR8OwZTxLhjuQKBhNBp
n0ZD1tmsBFSihI7BMiQGta14SBElIHZKFPIuMyxffLNZeidDaowcpJUM85Y4F07D
Bt+FDim+3yVKcFxsrsiXdd9TdszarYE/7+xXaTRqxYZlrsMkTbuEWkq13JsVspgf
ZisujeYJrcqqvxq6IGmcQrLJ8HYXlbxaa/SZYFBlJi4OafgE60yVEEOUBq01M5Ke
IAPQnVvyFJ2FTNAMa6Ef3Qhu6BPiOHqY6kLp0iB6M81wxV+XUwTQDHP70+sxCk3y
FHP7/rntAdyaOIy2AfGH8N8Ym+9LkDvQAUygIWzf9gzR8XxWKoWKXfP2eE75dyIV
fMJG84k5KvsOmdznKfiBzsI1PT7F3IqoBOQwUlGR7uRAUDWaAQBXOaC0589Y3wH4
4HWF63TXL2I6q4RihaqVgWWG3YGdZOnZKUKadwVCglWcf2F8p9Ld3aZJv5eeCjUJ
sF9X0F6KVtlHZ0Y/yvNtSOLr1ue9B7vXhCh4jC3/sTqaD/QPPUNpJ8Xw2pfjuPkX
+LgakxHrrjzxWKcBA7iCw96pqxo9sCcKv8a9Lng2wg+vRP4kKU3tKWhnkYjLeVUa
iA/P8EF+1PsFScCBdynitSpi5jKFldBWPiJ6BsJHe6tpz+q7YNGsoXo5FbuDWM6A
WN4+Dz8oI9C7X2bBSqq7FeOvx7bqNr3eLoajS5IPc+cVSru6Fg/Ukk3ab/l13qAP
tiHtRYrNKYeVxO0eNpGe0n6Im7jFluwXDgqY5oKskvVc5Xtxert1vjg/4ddQRCiG
QLMymeYkK57bsL8s8g/1cRlWlMejZOlsFRhelh0cB4GMxYJAz3KE+y73gP7eBnDs
Nq91zppJ/Rrqpc4Ds6nR2hTAxYHGn1nAWty/KthM6/ZgtNGhwLoWrJK5Hjfm2JH2
yJCOv0KNMJYmI1eTXz9GmPP0pDu6D0SIc5/mQieRnjL3h4Cvm8+daQsGjIAVJQxa
q17TrgPLnIY1b35vnKDZxkS2YKwkuhtoxBCr6NYu4dFpPfFZTdC2+u687P7bk6aI
LEFCNC0/45LY47VoaT1bzCsjb5G6M+aEnODMQ0uTFJflwsnz3P5n5tAChqdcn3Fv
GToc7S4MEop6fhuoykqUk64fvRPfztO9h2EzohjOZG+PEjlv1MY7Fwa6M8JpHRQL
S/IbRrRKTViTTGvuML/O+7OnYg5q0Wn9KNrVHyVJhGWUGz1BZNrfsoUwKLFDcX6W
5oI4IvDX46dMAwvzw15Z3dp1bvqhL1exP0Op0bJ73XwYwbj3M1AZzfVR5Hrz3P3+
J+2GZ+h/9B1GcE1b8eOez7lN4Kg6LvG6plY+qjMNTYdGIeboO4ErkIE/vHD5E3h5
iIq1ODLkCS3ilFrnDXYEW5M1XT8umFOH9dwE/niNTIKK97RCGRJilZhkHnZ7WK8O
ta481jeP4chGuBOIhGKzww4CE8XEIUHUZQttgPrPstHAAIZQxjKZiZg2e9zeuyfW
mpdKFEhzTGBDXRHZBzNPSSFPfrDdGbC9YF3WHGGlWVQvi4w9zwgr+LZLW+eQzdAZ
FIAypjXvr5fGlahd9TCQulyRcXyjuNP4168iNPeGfN7sq6FeawX8nE+8mFeFzcAl
ZFobZltBHnZJ/uThgaRKeyRnED8c+Sk9qibek6gck5i2JmLUcllHa1RbJuUToAPl
nZ8LxuAamyf1u9RQZcDd4VifZevLqgEMhNerhPyC77RixZqP46+xfcw7Y5iJzp6p
xsBptKcNqRn8t+1pvzOqCTY4WWNJzGw9WJZhw4HT5pfXWrApC289ALinX22bZwT6
QO+7J4CrTpMW9Yaa7+XSS8cGO5ORVJ+Druen4qrKL9wkiKyepk/yjhcMtbSt/wKU
MNULIGvPjA9gS2whMcYGbgJ04Hi6N5JDGwudVc94EuvKKK0UAZuidI5JcV0NwwPp
BrQM8UPjJWpt5p7v8ugnR/Y48zxHbLzPhpZjaExLdt+uEC/KbUEpqxk8QJoeol1Q
uNCXfJ1Sf3lQ9pwjSIe2xnx1C52f2AhnAY2sLrac5Ga2aeXwZMg1t1kxuwfsU3yU
6CzrINGPpi444dBKG/dnEAPmmEMr1yTGEAFWpsF1sK1LHfd8MzO0/hM7GoiHirX/
5aB0cbVzZqV/CotVOU3U9Ellb1PXrQPr05TtkK9g8nlQNUWFXmQkMi/uOpdB2iRe
dYvilso+WQouYep4CgQhYJa81l4ogvRjj5/kpq22Hmib8+MeEutZIn7ZkU8X2JiU
56gxypheLr4CcNqg3JvbYugfkS+WAKoedlqPlz+r2mvVhEQuJzsxsG1YTXKhzNs6
3GXV6EPUerFOEe0MYDxbNyOVzyOOvhf4iXch4MDRScPGebPjH7bOFJFUCz/1usyJ
W36Irq2G+xwv2xqApSE6DTOfVR6tE3W2OOI+9aHO4ORU+eibk3G8vEeNvddxrUfO
eziri0VMurne5XNBQasqV3YVqaEmAmdpy1rtah3HjcCB5eaex3rDuXt3S2+29gHY
IrJjYJouALBeqidHMVIlhuOJJ0vUlwpPYeOd7vMN91wW9fUQHfvFqD4gIhuyYGqg
4imX+sibU0UH3yzZJfRaOa6WnRm/DsxX8dNQQ9iylxonYSLzIDdYWWEVZW18FUrD
hYPtcXn01NkbSk4NLUHINP/jYeQ2Up33z9nGw2H0jUvNDbuU5s5f1ETQFW/r3Xvs
yzGcWW/HlpQ8QIgAa8+tyTqvayo9azky66McDBrNcn7UwA431xivaX24h4q3N1uG
+FLxep6ajoB52+6cNAdCS2HN6IalICahvn5Vs/mupnBROYaW8VQ6KiyxtQtV45Ea
TdFcBVRc02vOYXnTTDuNgYdAHND/l9TjzY+mxidkwZWQ9st5rq+RBsVfDjOMMMJD
Bl1ucNL8yUDLgtBPCS9NZ3kMYn81Eis9VKQCuNht7zcZW7iGGnA7raoCEzAidIkI
6MDVWviCgtCT7R4etdA54jIHpilwpScKZ7mfbR6Qm4SHkBGlpGmElh62E3iOnlFi
CQBWqRU7eBir1Hbm4oyjbRm65rfw6E7NUDrPzQRQPLKcsWrQBB5kDhqzX8SQYAs0
8nqT5qm3hgpb3KVT7Bx0yjiepXYpAuz2/uJX3xekzfzRLa5cay/1ye/ev+G6lrbb
9bpdc25DJFPzzYW30GfA9IePwILWQXnCAMV1Qge4yOgLeuZwPgflkynwkACn/BxH
4BlOhuvnUvNoQxO0LSyiCIN3tCQHkRRCRVC9qQL/dMOVuuNWV9tN3EY95mBqSWi7
54LBqF14gNaXjynLOvyI7koPhbdjGkoGDX2T3QDRZ7WaYL0uWZHBszShGZJWsXpV
xQdaSkozT3zpk7mYCoLp8CUJp/JImApm9beZRdYJRGCVcSCYCnuN/7ZxXaipEW1g
9kI8deHkBjKHoRs1sQgpIfFZlHi4T277cgJtGmUOlOIJPHv164EoT8582UnTXFZS
PMKqRxQYiqdvr1pXB5OlL3RfuYP1TRHIYSz2FVkBQ5rXmCfFGnd67RFec6hrhP6v
GA4/IsK0tb3d3TtYrmiVLWoL7tVC0olWxFtDC+jxWMb8g+klQ99KeOSLtz4E0pZV
vnk6/9YsqutD61n6iBugUUS7BgivzYeYhf8yaWMbdcWEpsiBHsUxdEIseDXrohRD
wBPrZcOT30BqG0xN/w9XdTAGYHprjM+VfbRHCMpQOv8ncgZ96Qc0sZ+atl4DjbpQ
KzdLw3aqLsJnOuib5xmog1Kfid9gw3izdAgCkv6ono8r8bA2bqg7CFyfIEen8axA
ieVcL9lG4vuwFcI59ZbFhzuDpzsGVyDhHXhyQ30WMMs+j1FDyWCuil4eseA1PUaT
FTdWuvkycntQ3+x5jCn8CwMN90wW2fPe9QLufoxq5xJ4aFIJYsDthYeAK+M76K5z
BMgn9l+cW2CsJSU8eyUhBV3WIXxqBDOb1RA9NJv4tqhTQgZF7dc/DBTRM1YQY7hh
l1/e75Wqyncs3q+ho1WvmB2QSolOf+u2B58/Z5VBL7idWWk35hOEJd/RZqhvI+DV
A1tpdKyX7vh1h0n/yoyQ/n07Vx8TjDKYyt69l3Ll0rMop/zH8UCdZt3jQPBLYbLE
SW0RVRcVs47UdISUbUHPRqgP0g+wXYYBkSvh23N/Jd+WkvbMuBhraRlNSP/+jj2Q
ND9B3RVdPPixfphHJI1N+4UV7nmGkzOgHfqggwqqANyvXcuB3XmB1xc5mskIrhZW
xuYTi6lIl0uzlJtXL3KJTP3xNAWExXwBQbm5jXO4xGAU0rJ5MOrMQgoGP1/meQ9l
2MoFqDoZzkxnFxdB2KLGLNvTuxeGl68i9icmImL+U0SFyhF3d52Jkf5gd2g/PV6V
2cLuk1WtvRPWFegEDPKMBlPK/gBjycvezdOzCT0XPVj0Ze8uZ35PU0fdx96oQp/m
e9Vtev5MtPUfQsZrVv3ybm4OYgCqLNhhemZ8xB73Nd/DrJ/J3CO2YdyY2ul72Wzm
1dwlmd8uYGYVdYfc6r4EB1mfLdu/rsj6sD+wAYLv3gVHK3LOZH1jmXsrvFioEEle
3Hs83hZx2Y63IWeFGxuH4HlWp5iFA4LaAMXR3c+4V26HxD91XdtFD112WMyh+M0s
fk01NWxhR45/FGQq8UkowgXJwXHltB0QXSGdGFvzbHXMIGBw6lXuWMAOOMCdnYdW
w9C814O6nZKxc+d6mKvNx0hrNHX1zAxuUJ9MeSGs395MCZou2FJu6W2XOEA8hAfg
Rju0LovWbnzWBgkjnzNLtaUCgI5dXiY0MBwoxh1MOyqYU8zfu2YmK9+M+o67GPK3
CVc++NuBcP3dv6NJ99ADBW0Tb84m5zFNkr68T3gzsg2gMZq4RIltYvZSmQ6t+oTJ
0iUuufgBRszoayggOnlmnbOhNKTg86aaBwEFi4503xja5MuZPQnDUcM0g5IPjWXw
zhCV0PCATXX2GeSKUjH9fFFG1eEMhUnwb1uu+4AlKqf0Henb8o2RxoeWv4YwWuDu
1FwQUqw3FWBp1pjxPpaX9QQ+J1qoW8Qm6bb2g9VI7mXODY0SD0hc+/GRlIsweBIm
/h+uVzkrY6EBGLsVnJKzyFNyY1RCxTX4QgUJPS2ca3mCOFE5UihfeZxvMAaCZSeJ
6oE3OfUZzyHWtFhvcw++265gICiakd2RNjecqwAp2b5GWIIaaaZr0XotbMX2BHRA
IFDjp+H27iGjhGUiY0MSXYUAdBURkHrsmMiTPKl7/a3/gtfqc8SLj/kZJPEKyjjB
kiuVEUP9toya091wafCNjXVkqchcBsYl6s+EmSh+T37XsxmE2qF+8qfdtLVthVMz
4iBw4F+xMdDPEEc68ourF+t3ZWdtqwtu2B+ddlcETv58XB5NZ+hmuRc5aT4v/RZF
DoZ3pYC4OAyJeJLXyuRN65h0nIvMOs24gRE3wlAre/e33MakBTuTVSXi+vaGWxj5
BUXH45ZC2afLG9plUXwUX9lijd+PXQDy1M20JysTMWxL1xj5OkY4AHvDgMTRwl7c
PyXYNUD2o1TnMyTr2hReVl2I7MpvemODf2rObwIRs/kgXvSp9k52YoA3/TaHSDFO
Sh6TLSC6v7z0gVVNDBO8aCUb2Q0k2FVqAkxre4OZuYVEh9Qeamy4jqeklBRKUGiI
ew3LcGXXjTD8eSj8qhC7vnvXSzv2FQvpjMYYwF3bsUqsZX9h2l8Bbmt+X0rUjTVW
ApbcwTZnfVw2Qc6O1/yxUDC4bmj+MDN9+xLS7nzdTLCN8otLa445YI/QsJZurCfp
V87VIpTuBBxd3glc+pJpNxC+0dLFxhcwuQaf/y9NabDGoQkUlKQF2vfKF40va2U3
lnsoH/Ea/RQqpF3FVpgAiGHg3DKmm9nugNi4o4FfvIInp0t3rGpD2ODfsVYap4VM
W4qRAZElwNrZawbz25IEt4jK4qkhivLSbbeIakXyldLm8cV4amo26Ze7C3f6tdhl
tp81eL8xqIGxiI9JSnAu3y1buOUstsWXXQDSE6G3sKUXV6cHVtZ19VfV3y8ddfvM
lYyYfOfua9BLdiA1xNX7jJXVXkl0nQIyz4YBtDJVyPgvw74U0s7psvFbZdr6GW5G
Lff6PYldlouQ6f2vPOgGDA/yWGBFpKJzwyckWFZ+C2XwFkLh+1V5fP8dCF7HkhQ3
+FfgsjIEWav/N2wODdNgU6mT2LrevUXMM+UdxUun47sp8m9eGIO2vcDYBeziCKIV
rK94bYKOoqnEgXR/z1versQLsKdyDBS+3Zy5ifnGIzI8iBmFbp3N58EHLod261E0
XISeZWSO6wrXprDVFUDVjgrrNy0YRFSbcty7en6lTUktAibDXu1dDq5ooZeETQis
9uN/bc/0GX53ITEpjIGCfoKFclhs/bvJLZ8VhuzlZipVpcj+fdUc4iYbrvc6oje6
y1gxfWpUejGN4Zf5+gs8Dxiwh77i2juVrdMacbQIWhccfMLK06RBlU0Th9wbqmTf
cp6l4K53s3Fm1bfXQqw595okA5fic7xS2xw9IcaqDgnSlZQDb8n4OUQzNcwTuBHN
amq4Y8sWWuyEjY3TR+6m45VfRSx3kdqAOzin800QhPeNUDaR0GE3y7UNebtcO9AA
Phljm0YnS6+bzi2qlFv/R3mkCca0BSzAMlHOQNQE8f28kMnyk5OgclojFjao/p6p
nlPY9qc27oU2r2D40BaPAMqU8b3Mj+RaUll0aKrHKAtYCDmRZxRI2r7zD22t4QF6
tjWoS3Jo9yF0VD02wtpQ0EUQRFElKZ9pzr6Fl12Hb0j9Cpn8gpSRLYAv5ACCV3UV
iTGMntx3IXWAmzVXG6xtUu5UGToFNcgidYnG50DZmYbsYIB+vsoC4bBui66eR8bg
5p2srt11hrD2mYufDAUvfoZGCEGVe9NxEdJ5H8et321ljts/saYJX0lW5xeAAl81
z+TE76/V1W9oSdQF9VEiDhz4KT6xzP5ulRgmxaCes8HJXz5ZMxstQ/okKzTvfjjG
R8iVnCWILwObXHOjqhjcrLwkl/x9dd0lEQbEYi8BWHRdLj2aRPRwTjwR2dRQ7ISD
oq+JPuo7j3Gp20OYIbE5L6yIVnJ6Tm5ypIZssCQvjV83hbmSPBK3flRCfHc0NRAy
4sqyOyveBbZ0MADwTHfLlLIEC0pWwe5QGSv4Caw7X0+BOsohsCVORT8oBcOMnPca
C4CT4WPEoJ6465Hir5WdJHmokcWbEBJPjTstMnZozj5bxYtuQPN0C0w9kRMoGWG9
R+WF9M9Ac3sKiMgYOhBZjNAAG85fYBVQmKqJQjAR1AkmijSjV5pULGFC4eg+mjNh
0QcG8gKF6WuRWVSnlPFWY7XEYRcrGn489roiQ+bAOT1wsQEXO03xxrSAv5l63iEH
Zs5rLuxcsWTrHOCvbJ2npVBLkt3bCXqEmtz9GQ6We1GkYoIOppQzudS8FLVHcwDn
f65doTM9FdjwSbrRIR7ad7YxWa5D+DTF9uKo5DK/WqzqikCw7HPdQ3qNKh3rBQ8L
oVr+MyXfckjXDz7PGSISq3xU7f+JTfPi0kLHDBNFezAFUXXObQd525DThQBo46q1
S6Msf0q3z7NwDMWDHSaJsuVhFj5lRNVPIMP/UCsNxe+iU+FHwGcuoBiB+b2UevsD
B05a4Hj+hqFoRA33/ormfCChoWlHUUu52DrcpUf5har0H/aolT1ZJq+4/kWWiUCb
qjFjJs3kiKgXIMFNPqpPw6VJl1r8q2X5Mg1GslXA21PVbnzBa5LXkRrWw9L4lIRQ
a8X7Yh5sSXD2ArQEU/YiMNdAzie9XRDTYD79ixkZkqVJuzdPYfjfTWVsO5DUXoBC
oeVlINe5u+j3LrBbkbpdpZJX6Vf3O52z8tFKoka17/sYN88eVk8ng/lO0qfnQ+yL
nFu09ivRDq9YxN0ZOAgZBgO0b3/qk163boQChnCaHTbL1paDGMCtgOVWqlIZF/HS
inVi5Q91b3w4HsznSIclgXHi+V2eFmIqCM/HnxCAiwDOwaz8/txCBGeHwjz7EsPg
r86lW04nTFBX3x0/o4lw7rDdkCS9cZ3cTh1x9WGnNcGI3j+cV5NOz/3eZsq/w8oR
a7F82Qt9pkuNoBZFPsA/LZJY+USZRiPcBoZlOL5td8Db29L6R8ubvPUl2eGHIjPV
uubbwem5gu5TxWYDcgQRnUYmyX9cvt4AftmlMSL74OEqdWqGv19VkW0g32Z/jvSo
skulUAlXOL1t4cRIdLr58kmqy0HHZCEe7eXADSaGakI5q660A6ukKQJBM1hBGByj
8B5+imQ+lfLobhPvxjTykuqMFfSug3N/CcC6CpUVFOKiIuIglr+mj23L9pmynH5o
IEgezuhj5wHMCLyfjOJusyyc+U96WgW2usxSw2XuRr5u5K6JHhrjoqvHPQKqrzot
jGnJQ+Dkih2GUhWviBPIuwl0DxUdbAqCprVDPHuqMb4rvENXgvh9mN45gfsOyRHP
r42ap80z1Gi/NKliomsiVxshf71ccL67ywQ6GJt3DqYRmymYD/JiSo+1m/rcvOL4
0Ku2VPuPWnoryzuPMyD8oGimXiKC9HQWeXZkTK9nJxJJd1s/k7IRlNNqXHIMl+wW
2s3C57GqwwV8JWIY8mNZUlW4WRKv/psLA1o26WDySlwSS6xsRPIkQ9iDiRbdGB7J
CyD6IvffYDS3yjoMalsQktyK194yOEXRJqRZtMhOTvjtHTZ3Ayxa92TqYSqondWW
5EH6K6eTZGrFsfnsQ7bysS0v4AW6pBC5mtZKt67BrdAwH4ozyxGUvFvRJoeN6Lmt
2YVpfm7GuAFfRrLpEbQaDrQo58PnHmNS5MamJ4ows+8eo+Mzfq42kDlHsSvGtujX
IRwWjQEp1ait+UPPXVupqbiuai4OtNA5yDfjzJCKhV9SoYInSXl8aB/8tIKr7vFs
0nEttU+zbQ41h8vJMGvBQStQSu9NTf9e6fMaeqlSt3pSx//C9ELGnfu428W/nMng
bhzlySYa3hyvbu/6AjMExh0tqJYndhLLYt30ba0plnPR2nvhxDYpZQGjlGBdfHoG
2sQcbaL6y89ndlL3JBTJZOuKSNDQWnWVjxnZGL1ehO/WABlgkfObUTYbxMkxVsib
MT/WQnOpMr6LoxY4Jm4jogGUVrWCoDNglVEsIDEtKQLAhgyWLJHMucCvQsGkaF7V
X13nxnyIT9IOInfhvBc1BuhFiuruMbbL+4g9m5nsJ9MgHnm1mRj3dZhbmgvNN2Pu
VDaxgJzuJPC2YA031T+aiYhHLi77kj7tkmzU445/v/9c29KLJ7D+3c06+Oy8fM+d
4FKRb246CbDDknRNQK2xbHaTqjV9PKHaPjq4V+9KUt+FIlNeHENHgGoJde2Ur5Ma
WmGTEYzJg6FcK4mWP389xFzI9oCyqD0Z8bYUS3An+a0gbfXCXDg/n1mMX6GKD5sl
rB789bSRzwc51DnAzCpgh0iRCkdC9tgm9opRW719wLx1YQs3am6Q3AnbvL6+7LvB
sQrRMkVnTwLpRwTcuU8rkyrf2uraDzG26VbB7gQcN716yFHtTl5iP0OrJE4BkJMi
d2/p0u+QXcuFqd2gbzPpFXiIhzRmOMNNONLQ1KO7WzBbMA4TPfXVimoGiGhOjEb9
FPCtsmd5C5xfSyHqCZOfy9Tnt7N0z3GWNpx5woSflBl87+M0Ig8S5OyN40NeHbcL
1x6JH9anLVWNK6dPEfTtfh6J4j9XEdUyU88WRQ4pTMu17JJxwwFtJuSY6gSBJREc
02zAJ9+ujOF5TmO4V2Q/jtOVaddJ/7JGekOfpXQNfCuRzRt+P2Ko4VIuCItEgDSq
SeYfvkBRMkn3yZJ4Z7XNX/sm1muIcBA7TP0oSiDpBtMCwWpQ3MCtzxUxgBIV7T3U
nHHyhmbOR9L+crsQIBZKXL6QEtzvQRaTXl/2WNysSP2uZPivzt0BLiqudzNdnvNB
8I3MADTdA3R4W0Jbi5AWRuvTyjK8P+MJITibq5qwNIJ6ym5lMSgwjUlItakxC26j
9EIlXPfPSXT+0DR7u8PzTV9FaZ7oMpgbh6GA9nB3rRbVtg8kfJi+XuSGkO7MxFgK
b70myODH8Gayvo4lQzD4rC20ZqrhWSgrb7GP9iWqf6BfYpEkdRie5n3ehgom13pt
PW2WfMfHmHWtK/7c6UOsVgAR9sJ7y7SPTbk+H4TF9VMxaAsX26HoPqTXGdeq+STh
BKFk9jXAxEVAimkaV39fcFlOs/1LWTXJ/gXJuJhTjZG0uX69d1V1RiN6+ngXhCfg
xk193nPWUD95+tRSFd/rPokF70HFkfTFfd+RAEzdXD7l78AKqrnAnpaEWeInmN2C
wuxFq2Jx7hMz8CJ1uBpQgnuWVC7P/fKeNt4rau5+1YyGQ7tYAyP551Zu6h0Y8xlH
AwlHBvESTP/Kr43feaiPnqm/GLLCvdqX8um/jlVPyu/1dJRj9RwNKgKMbQDQMVPA
JtySR8J7K9E9tVkFreaB8AzvOLNF/XA5zs3pqTPut7oTsAUXirnNx2Odv5Lqh2lR
hFyAr7+Z9teg18K4BiahOC3BsEiVossD1YLOgP5VB9MVQjUtVaAg4oza+DSIaTt0
snDCHWYdTPF4Vvkua+mUrjzon02EvNczdKP9A5XwATvXiUvIHYa2fLrzNdsOBmkp
zJdUCbxX50wrZtvLlTp5os8Px89GnLki7uE7g4lCHhBZ9AzPbvN/X7TiQqnaAFRL
CqJhM/74QO8di7QPl1AiQI1mV3ysX5/JtfP8mkBSCo3O6zDLlGmz23s3bb0y23eU
GZq1A3CRwnQYSHPMfyZNOA5+Av9urChBKSIgf2J4+yaMK/301R4DgibCWn3TP1BG
6gDsN8KrkGWMO2I74EdE+EpeORs39oXKpwJ1rhcAPIp02WlwsRKCFJpcboG3/7Wz
NyR/qilID7U9+ikPvmLJCUruAwqzHyXymc6jvtVvT73fxTgXGGXIfcV7YyZh2QQR
c6+SXOtcaNdvXzomgjtEhVTfECuzzNigWGIFbbpuGq1c95FYhEBvIX4YbaYDBgE9
KvhWDNGNxKcQbcv7z9snq73P53n4TEENYKckBhJk+2jLlwFHy0t15flGwVjr1JSU
aVn5/8rfBiEmZXPeiJj2p0j4Wrzci61u1usIAM2sfz8iUsZK9DivyIDycbx7BP+T
/vo1M46eIEqp59OOFXVCBLt6boZBn3ZfGsfxpJAf2pIdzJ9WnGn+/lomA6wcNKLx
A++ICBBeC3lzaGEOF1/ZAV7vsT2Hmz81016fbl4gahmCjQ+si0XaQU6nWF2MZCZO
7MitGmy5u1QRIZ791qQZj6siEg8Lv6MRbqfIVV1GDkSJdXemcPo5eSbKqfLSr+1H
VKekcLNn4dc5RZTRJ2kGkIdf7TmSsWP/S1Z0WFKj3LrzO/DGGNGznJwleJ2/m5hp
b6zXFggMae4n7IGwrQf50Ne1WZ/I15VoCVIGVZ0n68G04XmQ6OQBzsLSoebgTmIO
AfV5tvXLXmJ0W2U6z0MWNfm+Kf7P3eTJAtQEJvhGce/PXd1qC7/taCK6+D9RsOnL
82yrxyIzZ5vltdLu4vI0F3RuwfgbXC1d5lVxr6InvMJENHI5zXewdeJZGYX6l+tM
wxGc1IeyZb7s+2lbnuo6UN79Yyo2t4Sm4HEQZWrqkk4tbwbrdPQPsd9G2LSRYknb
H6yx44SmcGxnaiTC5/IjBnLUUzV3I53ouzkRkdjYDuOQxBJspW53WQ+H6TeMX7jR
5pEClkKkqwem6w/4jjuE1lRid200Sy7S751qnnl/GUMNlR7m+zMbRZlYKuzUFzsx
cc6Brv95mMCk0h/Ed1Cvg/L/3EerMe5EonfdEa73FekvnqHHa3hf6Ww5sA+x/67/
bsCx5o7ZejW4/Rnrf0xERG0ztW9u4ryDSgVwcEYhmKp5wxyYjeMSU0w/7rT/Envw
MhSFRknPKP70WwGuzLjs+M0l7/h/YKrAuqaVBdOSGFdKhaEW0KLvezTcnMc82Ej0
UMWHuWiYcE9/6GYlH8fKjxFZ6SvP9CoCcNHS6HjDVuM99LpFG/vGNs11WMITy2Ru
Qy4OoAHoKubKoMKS8fh17pnHffZnCfYAYMXOIQQn8h2vhlqw5c+aYwzv+gOyJtup
L0vdL56ruCpM+sNTXxl1fFS/StvtFb2iYISGXtF1PuAoTrNrZ5jQ/zNk1E/5QTSe
OoPW4xmhJomNSPXFiflcfEY8Vc0HlKVpTQQE0m6DqoqCD0JCz68fsbZY9TDSNqTu
XoiPxeLl8ZCyH7z0Bsv96A7F3s+FPkwrz+A+p9drXscIQYWMVa46eW8emSnCHFJ4
K3aW0q465miuBl2NWBxbECC4AMqU07ICcsUTAHiQ+gE0vjkMt1ci3Ta0tLGF7UWe
HaOTRS/1pJEbIEwSh3MWdXtIH0zZxAMPVmnSWeiUQ5HDbQOogfRFJ38JC5nXex2w
exPnbtkOEcYw+VKyUnpEPqp9+ubILQ/o4wjJ05S5yhGfWpROrdL14grFMIiMBwiQ
h/ev2SJRWGfkQsQ5dHdhQxaKdUil6x08za1An+XX+7OZCkdS/LdxZ12F0lM9mQnN
3wiMu5M5pKPhSfOZbJrBCYSemZd2EvzNcOyRAvPA4tF7H4zCm11glUyvrFc6113n
orYpda1xQwqgb39P0luMwwt91fxHwA3KNAKtWPBvbenybs7etE3vcXQNAVevXamc
nf+r8ZWhuE94T6yxLXtQy0GgA1tJVCHwVhQZV1QoUsjXXzwFJ/t1YQqPi7wAnkhz
Jzinrgn2xiEVIt5L6QJ/RhP0ha2HpdpECFcX2m44HP9vEv+TGcn8cafzjWxMUTP5
pldtmqFR5tAU/xodX4y7urnLm/jn1dEtCKr6qq9q+uJqjy5gIcOQXWyPZI97j6yf
0lnY7621t9IbNAPI7Gldy0kCeX8bOa+mCQZMhN2ZBMRM/W4H7mCwFeQeQ95w8XZl
WmQSQiSbamYgj4eOXuYesRlJAsvfCDcoRZaQvrua5O4OSsFW/NWA3ZXanXoTH1/5
N4BeTC+AGhvDFIfDj3GuMxnpbRy4aVv7JXBj4L0v8jRrgyHqo6FSYFFkYPHsoI9F
UEp0tOPtxPPuFYVAczHkR7XjvwuFUKdOP2pn4KJxMmNBAgH+OYp5XjQEsr8i2WBX
71PudZSSMLlqrdsMwnqpDYXZEEBFfvxIsmd3SiSU3K/VeFrCBHk0K1iUZEd+DcFC
Qm1FH92aE8Q1zXzXWz/Ze4LIlnOOwxBm6SoYKyercRul3ARn/o6/bmSxKOD4BD93
97AiA/ouDpo0JN7/em/a2FQe4qPp2/EeFXIvcViJLVBoZ8kXeq98Yj6/u7eZJKUL
ZD2xUWWlehztQLW72N6Gl/89Bd07aQ0Hsb0cRQE6u3SxTpAHqQCqvlblCfkWtuJx
fmmDUFwEZ/WHLzLlNXaWvIIobYgFtr35rsynXKi54S0KV6xs1i/g+5bpQMmHaNvO
SyOoKdZ64evu28Q4HOngCiUQ0iYYNsgYp6L6swSEA6B90UvHmAIZ8VgYL6pq6cs8
NGkWy31rwMA1lZkWnun5lqic3d3bVx+s/gX4MiicihL1G3vngoM7x6LAb3ZbgTQs
l2MmYZC3Rvwu8NRnaFaozCXHVi8LNOtJpuVQJFVfh03ApgtkBX8VsrAAxr9U+Nq+
Mbo7bN82N/PoWCOFu5l9QDddzeWXY9ebvNcJDAWyeZNJoZoTfVP68KC+zh2f6138
DIy0E6dYZPbovKixEjNNhkugHLv+pJUtTQnbGVDCIiMcJGaqznHOgXPn+vAiufHy
LL7J7nKO/hN2meyiMehRWlHnW5rmQwWC6w83KB1gtgST4MWes7jfsQFAlEwdORcv
uFt6LXsf5prIWwfeJGTkJRpEtfoDfF5ls+6ThFW73dAIWjxRuoA9LiKkr8fS7yM0
ZagVRutDh0TaX+A6LuoRs9JTlHxbxR3+bUIoc7WpehYbh+PMswS3zW8viF6SkRc1
AX5eLpTgkTMkwYH1tIr2avhHaxfSPLVp31av5zmLpId8ymgdASzLMoL67h3W2kEp
0I9NjyAY9+vBvkk7X00D2hO5xdPxm3A6xg42iBwF096vZTlvO8ZyBc1u+H0XFigi
fPGasQGK9ds9NyGCRqhIo8MZ0m3bDQl3Dyz5eJBJZMq99p25igYLMM5Sn84FCUCR
ob3A9rcMaauaiewe7zwoOxS6Xvy6ETP+7VhB6Rd7JP9YfGbBZVwkUH9ospxNjKTR
aHqXpZo9JmtYcf8+ZqdJ9Os2va2rqZWN5KExb6i+JSJHdKmvNNG8LTt5XqtTtqN7
pWt2iHLXHf8W/OOarsLQ8ujzxBY8azm1QpuXIn5GHyKie6re6BfgIccNa1qm7pax
th9JgyJmQiOcZwUJYaAApHj8ox8TluJDhCcJ7FR5j31mY8aXNUo3aUFz3V7sEYV/
quwnAGkn0Cq5XxID+yR9UKz6f2NmOkN8wQnDr0lIPgbvGMQj7J1Gq/Zdg2fMjRuk
zuT08yruzuzshFEkZL39wkW1l0JZTGp1fLQGEPz5iTdrO9fYvZOCoGK39n4rBn9/
0TNA6nO5Pc0B3Bu2laz3r+aUEAvffvAt84kHba5mSUQVB6cmvxGTBxaT2KT5bm14
eNY+LTztIM1QhmyuEZB2OLVykYcvrOUXx74eZ1gWOStI0ASI+h5HFCHweirWtmEo
+9ahcejMxab2M3xccGZsB39jFViGqPfpd5Vupe8aWsAsJk2XeSsr2ZtvzejtzcUR
j035eZ62XBeeOfRZ/r77tGIJPZ3VUSDOMD4dmfDKOeuznhPZbVamay84rcQy2UiE
yLPGFd3dI73MjeOTxpHJeFM2guBz4N16fFDRBqnEF2OdwCnbYwOMhK8H39UKnNqs
bGXzcRKFo2RK1SvBUiM6ESkVigoKSq454XmRREyIt3j9tcXwkwLiQe2BiaqigPkW
+PAxHHegUMIvzhXSt+PfUjjR133OHqzjAm7LSXadK28p2PW9XCOFX1vi65d0cuZZ
q0JynrXsH0JJ0yIVNMvYOi0eE3Lx8RmGK8UTVcZiJJdpIO7zf2vEPg7NxwCXNRfk
kKtsPv8z/CrVbiNbdG1stplR/4TMNlHeOqg35FhBqg+iC8GZkXPEnaPtg58U064t
pzuIK78Eldrbgd+C6b0afqTmE/YekP+k7nisEyw1TJHUV9HQSG+UaRrrhBmhAH7u
P8j4UgWrMHb0wv91V9M2TY8Dscny0bacFK/ml/69/U7AFKetKnNFwh+uYnMzpRi6
Gfs5IGNB82i+QXj67lll6LwlsWgJzjZ7ty6EBii3kyEJWNU0l6fIlsq2cx25Qqyl
hfZU1SdFg+n/9CgmI97+9nER3Z8ORk3/A5ZKfZmYEK7QJ8PkHIVMIbDTgFR4DBcU
XhD6lrGSIq9XiYIoqDnacM0+28tw8h0HSYlpGeLsIQnHc6WiVKEIyWpO96n17X9Z
BQC88zyJt2ndo/M0Y1e90NkxFRR0GPxsqoEpHinXGoJOFdWstrI9oBS5rcV+63hG
iQ8gkhUuaSq8/vvQU7GkIMsKiv+IKS3FrweULdVlvtWxKq0JiD8b4Gx0rQOwjq6l
ErAo5Eu8yNLaSJUjZxdMMI9TuJh6nxhNpnlbQTybriM9Vh3ehIXBRcO0yg05Y6lN
QXaKWW0v4X8U0Qn+DVOcjMsNiB6N+WGwob5kt3Xm4ov0kdChtdqGpsLDQNw1AEgI
0YL1NJFPAOcJZr0OIJeIWwVBN7F8Xi7Gu+UWxcuhgM5+8J91clDR8DlSyQQspJrp
/T+prL9zt7yJjlMfUIwF0oEsh8e8RaceTYXRMK5Js4Onw9Y8ufG/+6vdfSCcG44d
lW+L8H2tP1+eDQn8zSXGs9JvEw6uuGzvPJXWVCvkVmUx2cMQHiNhbX+cZLb8pGsr
A3aE1tidKR9WmemjVJj4Cw5YcNQwODY60U13h0DY9dVyemEIrrlJjf5NdDBkmFHs
AKMr+evUtApV1JuBymQLhNCeJ8FpQp6A1BDL4ARlkYlWhy3NtJjSI2wbvNIDQlZH
ifBWj4kmnZaYGxgnxZzdZROdkKynRdQtc5rscBWYlOL4D/Rr98CtwHptBYLW6ufa
YwCtEWjlJFnYH3g7hKlhx+OVgBhun198IWwO6qzHAGpqh8wVuioml2YEzwvg2dqY
/eOj49A0gphEpdlmeAxsgGPeBEUho2tPjpiwksAv5lWrwMu51yy+80W+DWuVBrHN
ryS7RfGYvOFcldmchXfiSDuxZmG3oHrA7IRm7nhSdktCim0rgJWnQ8VzwnO+bBa6
iXWc15ehf/cTr2qeD+bTLBRB+COtWFoE0uOnp963mLWmZEklCNHHKDAEMlD2hWO6
adNqnd+E5iAsVjE5ooM0ytYBojVZmgDDn94YohjEyRQtDpcWYksFCZQeKiBsH8lT
c/NZK0i734UeKZLnypigsyu/a+h8dB61vd5Ao2TbR7PlCj79UpVYJp+n1OhIz6bW
EOPLcxapr0HkOx6ibPhtdVfmq6rVweZFJVY2pfSrU44WQzEP1NknrbuFaaZN/pCE
DY6hk1y5vLIchetfzBlqki0yUqkwv6O+JFKxwWpKYUOt/KB80tRvDmF9Boy3DBb0
tHaAs8Vrli5+VPz+0ZjGdwilV22Ak472DPYWt6GcUmImbwKoYRaDznUummfj9dPG
/gIzKAtl8rIaWGQMn+vZYkmf6OkguU19RMx/C+/zFD16dICXMudzYqRIz0FVhPNR
7mLvI1Jb4e/MtZzC+mcCtySSY7ZPI6mTpd2GKPBPgA3GbYO0xAqv/N/KMcDrm9W6
/sCge5rNPIsSWG9m/yn8A2SQSKRbAigBE+OosDrDkh8s8YT4QWPjqXza5Niaa/9q
K+1j1D9+HrhdTKqj5RaeGSoH50L1dOjIJzoMuQAG440dw/UtXu+kfHbs8t0PGRsr
7FT2hh/Ueow3I9WVQVX5CygJix4Mutxb1vbwPbYCmXNC8Vry+/nnEdXO2vtvlmvG
HbhXiaXuvP7XI7PBGhVw9QYrkYZAPZ+n0tSIHrTCIqYy6r6/XmyyimQMRqyYv3G7
81+a/g4sCkfONfbkM/CUygGLsnX/RACphMe4SJi4Nn5rqrft9QfgQRsXWW7yAHO/
yZD0qdOt6aaa43RIUci8k5yTsLfEU4DPZ9t2hDjsBzsAqVhajFajA3fdfRTapFPV
V2g+aziKtfJEeSoDtEPjFaQ+dVXOWA69Yu/8Xe0nzYTFEXQ8w0i8r/HRU6ISbKMc
hwGbQ+kvQC311NA9K+Tb9z/CuyCbTMrIqcvnBNIZ3Qi6PXN2rd9rjJylKWkab3cd
NO1PtRSiNRXC8hWgAvocVUQslXYEd5jlrtq5ibJ37rvtUuwXoyzHg1MSk2ZyRpVx
QFekN1+iA4kD6P+/2DcWuO3+44R58T61kbyBBzA0EInV7ZhXtREvVRysVn6N4VCe
y9J/RU0UecE1e44eZ1DMWjGt8V4Yg5KJGRhb5FXURwSNBH2B6cBoTUtpRvBiDkNc
2QmUz1iuoQvV99v0pdbI13BKU9fcW/6qvNyl9JUSjF7vFX6dqf0mdUdW+xjlFW0K
LJn6U3ZiiNzztkSN3J3k8cYXIXGMiWqEkbbKMnopKV3ohcEOHl6rQc7h+U/u1C0C
Cu3dYBjgGX2My6qcPX6rizJMieSYNfW3V2uhdqLNoKV6ofsdi7pSCuIzcFpS8jxf
nNabDMs8ThFzqPyOcCKJdxNT2ijG3+bQ/WjrxU5EnWwqwZP7RHSzHsiXWtNoLDiJ
QKlAGlrYH7AEgTsGTT+LAexDJEODKAG15S33Q6XebjduixurEFUjUi/iVZANvGyg
Xatk5GiAJsWudMin1JfgS+9jnHr5JJ5/FIAlBkfmV6djI4zK75wN1bW5/BgqTRS3
vrz2fbOsZoxY7ylLy/eixCvNqtWjf9Ui3Mw3l9N7UD8i9r/LNpFzG9kG/gVGiJZg
nvZVHSWqlvaLiDIhln+mciWsdeCYdHhVhCmhd3R6P9Y3skGg+SPatr8i9k8S4QBd
UI60e37hrInZfGjh/KFUBfkTxLG5JdmXGERATw2mdFNtnZrme7Z11NIlAOaWYmWV
jePLO8Tst5BbO3Kihquef7Z2knJ0yXKGBCXrO5cC9rXsB/jTUH5JT0Ifc/8Zt7zD
AkoeoWpJL/FH2JlIpSOGUlmwu0KEqxn1rmUjp2rJV/ANlKIf8zVGnrRB6p05ThII
Vuap0g8YTN3OwookzoCTbOB8ntU0CE4vshRoXxp6uCqhaJ2tg0z84EjnyYE+VYSs
Y0yWeMUVTr/S5uLRZJaa2+Vy/Z2MzbI9jqP2dSrIjEYzYWpZ6sbD3AG9YXUiVb1v
iaIwtUGAgK0LhB7UFVxSOwMF/bdjZzryMl8Vbdj6gLcUDtHKMWPGxwdK3NFH3RtS
4oIJLCQAWrtM/inA0CuTQk0ALMlnLdxG1UXAPLO9kQXynKaollWSq9U5mCVlrSpT
D4LWOjqr6XcnUH37LSvfu5dfGL3r40tvPG1R3EXJevMBC1qW3YnNcZzBipX1RGTC
eANYnTJpusOCGhgOhrQP/5fngl6YSQH3uFYqZr7OkLjgtWZmB5yXYbI2o/HDLMqQ
2UIdTbK9Q4qv8eu00OQ1qjlYWeSA5S1sNn95Wght8/3UZ4P2yxuHxyfd4hrRdbxx
Ppgysy7OmSw6+aBy2Pd1DZJH3zL4PyGS4GCI+EFzuY4YhEoMbjfmJBBwHKpQcrIT
Fw1YXCoVbb5VmCQWkVpUNQb5g8FIHnx5dUWcKvgYQP1dTXYmwNrbO0z41/MWptP4
uHrBTQFlPZr12QfuLQahYGYbaVYNK1WpAf+M0lM0RjoWS70/Al5Za2B/goutTjjj
xxBlPBOG/gPsmWvzgHauOFeviDWhbr2OnD9yWil5qtYTqR9HAXzW0huPGHF6snfz
Tcgn19XQ4rEwLKelZV2JcT2ee3+I/+/aIbwFpHAGOQcze9C9ESmh8mRg9Sna2Rzc
gvbtHZCfumWYYime7dvvkwRzhD8MvR4mm2Pau3w/rgD7xaZ+eNDVacclWDe01NJ6
GsWSgI9ojxsiQLl/h6sFMn/WcJxZ0DpLYbccYSSifQTKUXiDPAIHuQXtCWAmfDjZ
x1qRQ0QBYW7WeJSpbtGtxWmYJlwM6/C9IA/uVkli05RxSaSoNAoE60g9YQlYkgna
7wTWX/S247qDXitBx9nJBcmwTBcCkSFtcu9ENPoFsnomMtX/RvIGgHF7DY8F8tT9
RpMu1ZpovsxBNebXxWtEKfo7yYnzCUTAAxYM9q7jTmMOSpJqImNAblbV7bgUK15t
COPT0vV3NUMTuCktaGOawtBNhPlk8sRUqNTwfQzTMXiXNzk04XBoNPHhjJZSEg0G
Tn7ZCbNSyRColag7QA3rixiExaw2OpZ1JrqWOrSaK66IcwS11KGZtn+ComXlJQAy
pHUi6JKDnZ/WwsedCj2424x0oWms12NkearJNEkibrEocoG0lcdI4EwxC8Bum8LP
FP1SXoE0P61aZBkkBWFFy14uUdPw3AWEwlkv3+swB/12iy7P0m0LAFTdv617qWB8
dX+SYXNE0ECY59TO/t1lQVN5J2Ofy39lVmkPczEBEK7/zamawDGkCkVFPROJ8fmq
g+Gz866DG0zQVKAYcoXahnX9oIOYXZKlWRHTatXith/xYlQzWEbfZWOTH0gYKaP9
0iPiVxa8IIzek01dvNjPPSvauqmy5kkbtvf1x7N4LRLUYs6s6Igw0f+yVYzFDlSS
R8n0jQtNRd88hftuW+MfaUJb5zv/Yc8g5I7rQTVu++e3RS/pMS0idUAnMMW2PEgd
lMvM6SHucI9CPbErfxOEEGBNlsgoOO/RSvJrKdyalfeew2KR6PN3xmSuQ9ztL1hl
+r9watFUXxiroKKAMitiu7jmiUwjrbE1TLKh9gAaC5D9R/cHeAcWcyInpBuBfE6C
WUzmtOr2pWuPhDK/9GnhWl6cIKn10I/8oTaYBMxrClLNPCN/3/1UclLOmcyWgTYE
CN5qi+6ZwzztCiafG5u3fWrndRLrUJWVefs68zXaVgQMJqs2rHL7s/FN0odGVCWM
wta7piv9O5XUOiUF628AMhqW980Og+K0Ympw55adBgm+w3OpXg8Pbf6Y+OwybSnV
EzUM8Co96jxsiNqrX1PNg41dBNL6hsbwBY3HQ0Ba8GVStDUMFEN4tAocVAY8qNDX
/jSH6uWw/Mij4epPTYko6iUDeaKlxZDwD8phzhPmvkoGOVMS6JJLEXqKnlBAFjGs
WlL3Z9diH2V4yxy6BX27yTPR4J6OyK4hl/1xxlFX/pIOQHVkN14BJ+L3XQiPjCKE
OpfxtmyeCnabTvOwCHqcmXu9ApdYXfFJA2VUQP39/MuCFBvl7iz/lUCU/6CyI/ic
yaiA3AuO5kABUdodiBKenWVpbA0rX3K7gEqKfuLMZXRJWRCIHICQGBM4uj0co1PW
Mdfd3NzfeE/rgEl+/fKkxqT3KoorhHqnsPoS7YYOwidaua/EcfMYi2yiv/VWxj3x
Hu/X0GgEcLSztDYSjkG8wA1/A31WrD+t+cEx3ac/wzVTfQ/g7IjDEfJsgipKXUsq
yPcKIdJr7WIm6SAnzmuvUd9KJSeqnWjJo1N3b1MFiilWOuHI+kv+7YdG9OCgi+56
DgVbpSOaXLBzDvWnVDqzifmqZlMzxvJY+5oHXtEpLyIZx1ZgvzrBGah2/cosP9+O
nMbMcJjobmOHeihD5dL4ZdJdN602nfygLuQXrOwkl9GxDgE6IutEtCe5xoy7IZEN
obP2ileA+j8xTlPYpNn5xhuYp0s2tL9MVvJNIsA2axuyy8k4wYC7cY1nIuiGKKB9
j1nW5U6bieGK2+8eptt3Lz0zwCrQUKKDB0bp1QmBaTUHj1orX0uwf0md3ebYMqsR
Yr9Ev1jkAHPjcb1bTM7ODqgqPXHHiCxFNpv5Vm/FOFVolz3/ZrEUf9PEXdo2Xum4
2t4y5ctjPRSyUS6T5Iop2BE4QMHUBy6OIUYmhOxNG5qARutfj68Hh1VZUGxLSzcp
b9rPCSUP1+gygc4MErnM1AwyV13fCIPCBaUqoyDBr0l5+MWUMurX+Qkqdv6urntR
GOLrhbclase7U12M4wYq1jj32tLvhc/tb2m+v1/0XD5vvxz4STRrx0/bxGyRM/lF
GphpKlz/dNzaJVCKQAwrPYV2KVlt8QIud+7Qb6j8VG7EmFuGLQPqJ7iFS6T9R9r5
ZffWsGGkocOzKPPRfiMzIEyNw/lO8QrV4LLoc3cdhBiJLPiNl6b4M21XQakuvj1x
06CAujDnfIDJWuFitu8afjN4u1s3HGFXG74CmZpQxx4/D/g6aJoTCAts1C4fY45M
cHz1CJh2DpnR38a/CweQinYcDaxGNvyXjUuYvanOTyp9Ic5VoOmE67S9Q854wFsm
Z6XuPmF13xiBCo82oiBzjGsw48rnINjxmaRCJldqxhpMCp7Om0B0zS5qWp80GDTK
bYk6Y2tvIZWiBLKQZ6Z4Pae9i4st0kw1N7Ye6ugo6E3seqXgpiaEWeTzGzCwEU8S
tO6hpPRhtKZ3+FBTvN+croIm4KBYO6wb3E9dLix+Zw5U64wwrQ2HaRbud8u8pDds
4Zz0ZhOp6FZupp5zxsvGsTdDdRhZH15mlB/aPwy+04wzgoI50DlzYGlaaKMfVE50
ifyGSIuiWvvW8v0hl21vblkb5qNlMN9aY05/5rd0Y06rOBYlD5zkUxRqXdabJ+ne
NWKMDI4WxKrPdmmFdZsS+wPiZOi4UqXmw/MXKDDNzHLEMAJCncPEat2oFHMXuxpU
/gicLATA++414LMW4KQClKr3tjPFLt/0twYsMYtPyj/6Sn+cxsVxx6rRnR0XfC3i
aOIFC80AQ4Tx4dyANzTCcI7Y4PQYA9dkgIjirdnLH5vMbELkJy/sqGriX5PUgmtn
5mwqsZ/48cOscoISdLcwKtK4Pz058SrIMbh1Gz4mOHEWwRHPZ818/psctCpuk4Mw
X1EEuD/D1OazzY8JbCaZc7KMP/h+If/yhkhCqTbKr503ytZA6pL7gv7sGsYXBsEj
tVW6RtJnTn0g9Nsdi3p52uX6UhT845JfWdlLF2B+Ea61eyJt0ifjLIPNJR8srbG/
5UloAsQ6OVDzKfUYt7qg5hbV8vpUeHoWh1WtoI5p8v3NoXEVc8uIYoryhJNzYFx8
8hsGp/Fe4mWHh5TWYcsqMrPA0SHMyiUoJgX02uxHNEVm09MFd3cw08sDuKsjy0v5
kb7eNxv+nsgh0cPlCe/rVYvxxLAORuM1UlmOV6UTxCvcegJqnFMMV1W5KmkXmoOi
dvIqZ00GmpXUunVTOrcSZc5nZ7eFjIvoXz/PUNdsPpB1o9urrMPv0G+RvvQriRBJ
b3fRb+E+VFAZ7jfWlql5Aj94wNrgkWBPAKBRiq13xehGNCADiV8Mj5O4x4OFbiZu
RAfOjQi/EQ71V5TR0a6RpJJzKKJkJufq1WQ1tjrwVCFjUVSIkIqvqr1O6qZeagEu
zulWgF3ghepJvJuYQ8j/UBemR1oPKv5pkDuTsCgOtbAv6MEDp967l871Muzn3nZY
V8Y3WOt890cRtlmqkLgJlk/Xv5gzvBVzEpp68R75UBBhzWpJeTefr/vu9fibCj5P
R2GJPGDYJCOpdiyDl3azRVX2StUx2PqUlaUStyS0daKkmPYWu+QuMhsxqDIn0j01
ZbygsU9sEfOtPw1FFCU+rffUwxo3vNkZwiLS/AYiDtFihd+wZNPguRdSTehWJBQo
VowWH5btZNQ73xry5RUMh36WpNRzYcI1uRcOpOKqS8KwBCRjY49tyeDZkFlHhQLt
P+woZuLj63PDdNPRNC1GALGWHtYff7/crl4/D7XgCyqN5ogzWx5wnG2lK5ulZZTr
rkzJIpsbzhigpwf5WQB8urY/wAyoNvcUyM21yILFRwYP+jYRms8FeatuzbtCqJox
CjoxYPRSByboH1MMLHBAjArwQWvw/Z0rLENABB4i41mHH6AebPTeKB1d6BYYt2Fi
zS7rCUmBroL87b8WtU4EyJnYKHyMKLqQAuoSsh6NUpvVBMvAUC+FB68/Crisy96i
I1uHGAq8en4eyrycwl1hJEx9G8ZU/9BwgA2LX/K5PmWUNYjGnX3E7MIMcBlpuU6C
Kx0cf6kpi3NFjU4kJUijmB7OPJ0UUeN+WlcYnbjYdC4svsBgbD7SG60AZLDWdQoD
W0OGthJ0/ogs2sdqmhqsz5MYTvZNnp5g6IirCLptV8ImgKelE5P2MUPACOBo4Fzb
cUV9u+U/3Q7SpYCs3Cq8yJXAbrV3m99k3gRiAisNMY6Te33Vcg2AuPnPCLmoI+xW
FbBfjEmjDvq3ltunFj0WIE6eLUHqU+ShUWQhFnJ+8Pre5NtlIiLHIqUIj6AWxKYu
4uRuJ99mt54iZF+ne6h7Sy+du49K4q2t07UkmEP+8SS8SuA7hfZbsjLuWPmR2N/h
oc3YoH+qK7uwEeCqRp6n6NuglGocWao2l+bFysqWfjsbX09RSvcHKhLwjhFxSzxB
BD9T8yl9kEMc5j/V8ehmLj5lyfsECReWU+JE58Ptc8cRjRHnlXdRzInTgl0JI1OE
fUA2TMTmNhBKsS9RnlABocUcBtgV/+XT6It6XwQxmMrPRdHG5bUiaVStf+pPeKxi
BMiCAQECeubQNTT2imO/Svz3LhVTgZ3eUtI5oXDjxTlB8MYXL0iXbTlMnvVbnv4D
Awx4UsI4MlWBR8xr/i0BwBRfg71aI4io/C6TPNOn8ILq+Fz9aTJkEsiSD3snMJtz
v08KbAApSL/9uksptvEvbrsvuYCksG5PI6cBPMgdJU949oTGAedx2oKea/t/nssN
NFzFr5TK975ix2AA3nxFsK6TtCF3O0GnmcL63YnUforhJ+gL+ItY7j7DURLXKM0K
SLRi0I5W4csoZydk0gF7t34epG/H+PehGQLC0IvGB3GED7oUFgAjrLE4jppQ2Gx0
0+sCITKrEeNDTY+dhU0B9vytL/et97nKl6foqfkiN8YsypCItMLLwp4yLBnioulZ
4+L4WGHkVh0U3TVykGbXwRdlYwEp9IeLjN7ntGXXXQZ4DAORwP1F3jC86ylQ5ORw
H4Mtn3oOhromzOZc9C7eQw0eeAsNw6x4g89+WqUI8Ny51dyJZTyqotqYFczCg6X5
1bvu0jCAa9hx9qKPRfhYOpYJBad5/P9rwAdILKausQNbP6rDa66rW1l0oO5sOS5t
E8m7m76OvGkc8NfeBOmOd8itJLEQ2zPDM4p7WZeaRx6JX0xRPCf2EPvRH/ittGdr
FFysmHBeZxDe3SbIhdqnAN42x+bRqbEr6Jb+0WsTIcj1Zz1gMu0h9Azr9UrfyH21
uzjAlfUtgsnrJfEy87/1qzMVDk/YIV83OaNequ7NmtojUr5yZANr/pYLdNaXOtwt
XUBOkX71t4if0tZgAUXD9p9YUWUtvYmmnprUHqNpkkAdvWaMbcjEywzj8u8RsNHk
TDS2I0KDGBtULrNfMyINIaru/Sy1b3FoQb2gX9zN1yNxpOxJjTR056ey/tvBTXV8
uCEt5XGzYEpJMps4j7dVAW5MzUTJHrBkVAY86vJ0p4fR2wC4CVZjKNDmcHPXB0uQ
/iajv7i6ONzlzdFlMbNofmy2kK6eUMtkoshZifsujQ39D7Z/thQZ1H4MMmEy5qS+
XWkiHw//FmGT/DqPv2UBWwhZ6NkM0+6yq23clwOx7XsT40/rT/NBmzCg6CMaSvfT
wEqyoNUm4/FTGlL3lRRdvCOJo/JrbR4eluoe5aaQo3qjpT2TKbARNLAiVBtyPJFR
3tN3wziQgeCpQNv78600wB7K9somTvGhzwYYySe9vMsqvwolWTq7xpEFF+Y5D7+o
EU5C/2OCmur55TMUFfBaqpZhTS14tDKF8eB38sPXp4Gdsec/b4E4GYfx6G6ai3oW
GDvYmT9S/Zkc0GAo8DTYIvPN/8mQ26G805r2kZSg8PpijF5I3y+C6ViF1Hq1rebI
EQlWR/7JeBlEpMuEyLztTGLMhGeQR/u7LMZaC1Rtk6yIDmG1VN6rR96r51Y0VLAE
gJwI1UqF5Tz0A9yqng5+W4aFr7WyV+/wZXX9bwNgA1dJ9prvqmUorpIXtowia+Ix
Sz8bE1ONARfxR4OIGv1qsiT+pQxaomsFi/QTwHU/L3Xvd9/P1jctAxJiGWpm0W/Q
QddGbJt9gyuofw3gWQ7jEbOxvl8nCivlrGTSKJkp6WNTGYNzXal6wj21OXguECtd
j/mH9dGJFQBfiwKUaL9HIlX3//IHlOZTXyVbjwc7oY7NCh9ZmD66BcQ32NdVi7WV
nG5t2Brgdyh9fJ0uOcNDTWO/mwjZ71DTyGwmlt74JgJHkvR85CU1bJiTF7vUi+nV
mb+KCv9iaDZn0eyBrMLJuw5sCh2tiRGxkAuFaNtGZ2pyREbuivwOilegVqvO/Dg6
ZhvWeSKl8jFz1V50w34ytSQqwfe06WQKNGsr+GjBjb4G0KKHwF+IqFtZo++fxyXf
ECIs64DgJHrggu5aLeq1iqvfrof5BgmrSou/hUvycWHxXHlAhMyJshosNvsXHKGH
nZlgxNiHw6KoOaQu70BccomiC5OqD+2mSwdQt52OdhfHtml8lD6bwk+S1mWeW7K0
khTACmbgH7/CjjFqv+lhepkd4cNIvT8+UIozf8zseg9mx+Ay9W8oXagbuPwcX2gw
nv1h2Euj0Sr+QWp3VfAUj4DoXteDPRaCJzqF80TeNHsJuN9wKhOy8SixLxLqog8m
c5QuRXlhvAbAMu712FyCxRZAOCHnnTpvMRlBZv4X1U5wlqWGuyjOgZUOZdYsw0uq
mSkdRsw07+mkK+gX3VnLaL4d8Ng7qUe2RCM+xA9/JGeUPUzC1apAs3b0k1KQPDV5
Vh49hi/sE3MDLaLuhWVk5qTC6QEeRXM6hQKm78u4XAffUBZnB5N4zYVSfBxdMokn
84L71Cy1VaRI/msIEjBsr4qRmSGYh3Lx/zOcU7QKqUoFaqPC46PNovCSiZZ8eyoa
uWay3UGnC1Ht9Bu4l/T/RbaWmdTiz4K3X38AOzNsM6yb7VnCBCo+ZQKCToPI7/Kt
8YU3cmygw7zQj6ziWKy/GO4t1Q9BMiibQZfw7w2jZz9cZM+mEccSHlxzD8Q7FHVE
zU0L+sVd8WJKluSyCEVhN46jNkiwxmVVosSCrKOzX39jrThEG4/jvf2uaWcRYWAs
/U/68zdAYUwoD8gz1WLuKmw8HGw5EB6SiGb6oOJ9/GQyPEapJAfQmwWlabpkQ4Tt
hyB05RgxbBWahHpVd12nFJbFhtF9zvOsBIkkAGRVFO0cmhI5U9t65LIAwEqunCoY
EG045tZG7WTAr3WBa7m7tO8zkt5jeYExXRmCehme3j4QMkY9NqbWwt6rkQ1AjO3y
+/yn4nyvyhQ4vBArO4drWqYcm5ZXTuSeZfr61SBCLek496azBtjhNqGmgggUiHj8
rEYIDZWd1sjsxrT1OL1bU4vDmVhqrSq+9M6moQEkR25jhD7UY6aDfDxgu/MoEBwD
a4q4rtpdXSPlEy+hCCpnZSpNxnt8lqkUlh85VYxoUVBpIeHEKxxsiYLJtBCoSg77
u61/dQ6KKZUh9JKBs0/BuRnXbsr1REMNES6TkX+3JjWx/9bzYoBg4mWR8eSNuGU+
BQVJf5bhrINburt/IUO83TeO7NVpmW6Wt62NawgiQwL3MMW9ogZKjVb+9K7e+AQj
o8P87k2Pe68txY11CW4eW1q7bRQ93hCtXDlPW5JzALNgXNiMR75KKuh9YXtSLk4H
TMSQ8Ga+w8nFL4/sSsAu833KCogmlj/xPH788FQKPVJw9cBeE+uOM6vNtGlkwtdm
iU2kNY/Pk3tqhnxJvedpd5PfzdEOtmc8EZ8MeTRgzxDnbISVUWfSvwMcMiZIIA0D
YG2YxsTUjSInmjjOUOcwP3Gn8RJFdcC8A/8nFBi2QmJ/AbHZieLbVN6UyCyA8jbF
m9FMW2K0zPnTuiEQCTSfLnnEB8npxoo151TvzEdLgBQRh5Ls2DEbPXUmxINv6s/n
S5pAiBZMD8iYv5kWIR0U1RXKgLu6DgFADomBt7fSbVxMxaqAVZ1HtKZG9uzCUz7Z
UvQI6f/B/mfx0L6uk1fZ/oPmE6ZdT+n4KE32lHkG1njFKIWJSyJc+bOl8c2eRf/e
PU89Zxp68ZZyv8y1/8V9HApeZYPnGqIsc3UjzqoCzJOH19UGBbCOq/NpRROoYy8n
XtqYjfqXPbrLXOOtdqWtPSwM2oWTtyZfYZaBMyGlRBWGh/DRSi2dz+XFT37Ch81m
wBqTv2OxlUwtlRJT4h7b30hY4u/OVBX+Og4MXfMBDuk30LKiv3T9haF/TTBKXy2x
aqVU0RLssgoFSqcqTqTl265jFFCb/6aWbGvecg02OMIvI1BdJMStq97JS7hJ1/gB
dNMupjBuMTIaUqnnXLRFQLGHHCdZY1vm04sndurJYmUxdyHOHwN3+Bdz34FOOEXe
d7Fyhchrkx8vVk8bq0ADqQpcid/4QQbWk9TSegT/rd/BANnWLeWv2VBSSUzGEdnq
Y8Js2Sk6ZSPROcs603WCawPJjSj3mlvZD3Q3E+MRREjBR8eBqHLGCI/51qzDfwrr
dK5d0V8kp6be4eY2uNHIYJjXlKlqZAwhTUh+/JD2KbCIISxoYPMvoSWw+uXQRo9S
o/aezJb+4EtwEIesW8PRQFDN8XMJhRbN/emBBEYtlYeIpfDQx2Xun4t5U2ojFIMt
xTHTmWbNO5dIJGZ3idTGa8n3IQ7VFf/QxMCt4cMGqKAVD2D9r6qhi2VWfvcGwJxn
vFb04SPGnJITCdz8ZDTCPazhaCxlRmp0XJXw2K5ucF3kPpscv+0laskKKQXXASIU
VRrwA8qJpy6zD/j0+SFkjrUli2arYfo8sQfLMEmb/gj710xxPMCsimx6NIodFR4g
IlXbYA/LFKhNtDiY9+MuPfdbWVZfyLCwljdgLZqza+mE/6tCnYSZA1hci7qQsNpl
vAVGMAKBihXB1OOh+i5mZfiBKPPQYuOm1tT5ivp0z+UKY8ePcCPBViSACKde+VC7
Yyo/S4NASM/42s7Za1BKa6otsD7OlpYbitj2VJk/Q5rvWX8w0Bej3d+CvGb9qMuB
/PwAEtwymmgNId/tkGz1Yjv95df+QPIq0NXqpwMeRf0YjvHtLI5w5N+Q7nSbJLJs
Nzl8sVamiBGhS2yA79zDafKJLBuemcLRGM0RVWhtmZ+eXhvV41rz+TEvTNdRxglg
rJGJszfZbXNwwqLKqnTA7fUl7/ySKoMckAr5Nf6Yvhgwrgzt5PsulM6qGxe37c2k
n4QTfBx8ICYC+BhIHGS+3kCOt6KsMVa5JlGKwIl6JdmHOVP7D5Ep2hdi4bVDJKeg
VYEmkwLZ2GYy9J1jjtlF0x4k1XO+eQgsLFy8aW3EP8RfQcNva5fm6Z1DV7y8UUAM
F/rJpGMFDczDFH9dlpvGlZolRkfy96jjWs62QW/CB29aSNNsvoPPVDgVvC3NJYnT
5IHJl7mSECZ2mIfCBLezdtIRPAiySZtdnrycyoIhP4jo03KqSlvQo8wiVDYmgjx3
JWXwibiLfR/bYOZPMq744PUsF6mZ3BhWoBCjCPVkCNwAd6fL83UrA/zq0Cj2pFks
nS/SqsVXI/mAWgbJZR2ncBHyOz4g/m5zami0pPzoHWrAkah4FboEgTFqOcNzokky
hRSIXsHRiMQKIiCL9KrcLiVy4LnufqLQjnrKXBYr8M16OrFuReLggx0YjmkHpIi6
q4sdGxg+eP01EV4XJjHu81Qg5JVfXiNSGfEWg33+azfl3wHMVuIaGtXnJdcPcrt8
OH41020CRMrObph8nUe8Jk9jONLT324HGyXhzi/d9aShziDY36ZfQ+z+qDr3Vweb
3yErLyVr7+fG3i9Z54vijcF2iQsxkj1xRUC8ywIRRxCOXN1QVYXKuz0bWuI7Fe89
4j7YXd8bPQiTVdEw0PHxc5qDWblxdeZXaW7HsyjQ75OG1kl05IztoJbqYql3Y3Am
POdk4dbQdUwgE+R0F5q1snsEQJT9hDKWq6Hrk1bMDmSAPLvClWKMbSn/rbY3rjN/
qJxKTlpDrbCL+KTrFhBSyFGeC+DHHCmuhZdC8h8eCcZRqJlBFT9EEyz98MwX+FAm
L+jP5pJwK6eh2r8ZpjmjxYZOOIkobSfor6N11+YYI/HCFtcr+GjaYDtXmDD/K88K
zuHvGiSK1mpHSIpC5luG1Y0SVt7H9nib4RjXYCeiWOnsiNdpvHGUcpwthUPOHfW+
JmAGH/eYKzu3Yxeq5A+NFjSuFK+HMQ0X5QzyAWDwC8jmcLqbcuOUK9US9t3lcoxC
gAC8JGR9J6K/tKHkcXmwDC2S6FjR2UgSpgr1y8y2rD2Qb06GqH74qUIchRF0LWf1
/1AySJov2MCC2HhEFTnW06yU0ovZVOvgHUGladkhr6Qw+XpBnxjs0KNTrHF/vBRK
VTlX0lB55m83qK9mQbOo5e6ekLphFqphi+F9ZTibbuqE+OzhfbULIXpD2fPVn7i5
CVpjFek8pNl80Gfjckc0do6+kuVyy7Zb2f/nz6O0vdAQewSruIQzdXJG5eGxu2Dp
RxIGOQSuHn/UsmoxqKkUMiy+inrlx4xZsTNayMdLNmPpMc7pbS8qRoqsGjs57SqG
iAlqpVIYqEtb2a5nUolUuPDt9feXJ0s2slKoCxC2v5UX1RE820WnM3w+YGzvAAUg
2hQqB5fkuLhTokWQgIDU6YWzwnqzRcLltU0TVDzpIzqnXp98GJRSnYFcn9hInmGX
n0vViKPWgw3gll5dU8wr0dOfw8vlsZEg5++L8NwZuBsZeuS+ntiA78/wc4IEKcMc
JGYcUYjrnrdFItgoaITWrtLTMgveXgTKX2Avoy+5l1eZ3Swn0SINJg0HTfSDMkuC
kx7mMTWzxyJoTwDhnynnf4Bayu5AEZ81Dg+RnTFM5ojt/x0mJCtWDcNal6pcDFye
fk63VPCUkELWDAwoEJhLAtZvgngytWa9tUD6lRydP5ksw0OcuBkqedG7R5c64H4p
tY8YtA+5OKp12sT1bJAIqz737U9Ym3hbdP6brt7lukp0Z/dCJ7d9NxFVXNvq6NgH
m7cNRTHJnkQ9KOm0NNURzGuwLDuoq1MwBVnYQziPZZxrwuJojnueDax+qQosDVnd
eyiuQbSdpSaQ9IKVFiLq+hDNGFKdpH6Oit2i/oESm92wFzs6Pk5wgCc907C2t9/K
fUb+qyim2Y4UArmH0XOADI6+iy45MEPHQNjbcC4M6qJrUcXhEjNNYVdJh0nJ4y/5
OC5BHg9+Ix/CLuXgmfXErlgH+0sIxiFsi66JPcChSZjPBQ+/5fx6Ay6GdMh729Zt
AIEBLAMuNuY2UCqC00yDjYhqPDhy1QfuWU0QYnORa++gif94ujeUDqW0ZVVIHn1U
G9lAXPbr2D4ZPx+pPzzf5bM6EXUKTXPAVNQkIRC3RipJ68HMFfTdnXNJ+HEnzNPc
o0YU+fXIDgaNoccPbEPqBTR2JuzSPwZGJSCI4P+ersBhla/HrB855+iryDwWLfC+
phrkxPnhjzKaoG+vdEH+BLbhYonDcnKBOnsRuZhwRcytg1INYXfP4z53I18mlO86
KRBGLeewYz3f21kJoujCjnvZLUNOr5ULNYUFmGoT874TGdONnTrus4ovd0BU71lb
ZueVHh/TIUtYToV6tLrWso7iZCKtdt1Y9z5S1MI2GbiA2uD85/GVuzm0wF1wtrD6
2Zz0EVGC63Xx7Yygma1Mf2L6GFGN+cXNIH4jwJsgBUX5FUg+zBj+pmNBWHUQ8tEm
llwWcPYBnZfQRb8jY0k1Qi+CRPvtXf7ad5dgwqbh9aZCW+Ugqop61OfNpTJYrp01
Ljp6+pI2GYfPUt9rv6C3PkDtfwSNyUnCOz0SvT4RRDcL/Nah8OCxE1bjFmciep83
M2NzQZZh86tIfzb6Fr3qzQapb6pMunQtqHmTPspZgof4zTWFldtOS4TxZQvaVQE7
WveEwrU4Ayt5+t38bjp4WJ0aokwrfIhBWFVRTw9IPFgPMZauFqqVg3LCwo7q4w1j
OLVi9sE9ah8CCDHpJkvTOX3PYH7B1QTVMc/jvMfM8LYqGCXfS3BneVSn48B1IXeH
sRMrUcikS4CICLDrJ5UPXDPLHvdsK9YUxBoYYcPjH7GIv2uFHQOMzDEhpxAhHmBq
xqGZTMPN3VuQ6I4lrD024SyiYmz3Jo4CRgMqlN+a+x5q1e6NI2h//16lElXJNIYz
cFbXvY7mv/e8ClES3dazMJ0eBLAphXwZXV4P6dhhHKUstuuO4dCd2FVv4xYzXWbt
Rjoz625VB5L0X+BtU37a/eS9xdJCh77bHwFA/vQbEhF5BC7VNw1jwBkoLO3aDEQf
j6/vIhKtRb1+7ZgkhKwrdncFXs49ecn1AY3fEZgH1U63AqaZOWeDiYEkTOIoKSeW
E1oR9yQ9tedY4t8CmIzy6h+ptsdmSb7DCGMUgh16LCBPgu/Y1bv+1rcGRP5o4B4K
FvpqUICYisOMb04240B42pAc01djBnB1hy2GCX4/7CTzDHh1g32N7r+wF6PordCp
GINh50NYODYCcV10z4zy4Tpr8gaCd2RdhxfESbtf2C6lqryLeGHKLU2iH4Z3SfO9
oGP/GB6gn9dmGBY4RKr1QLJjpCuRT8ampCgwzZ1plO1RuCC8yB3fMGeyhxuLKsA8
+Xd96YK2v1n3C5+TB0PrtlG/jrmGfJ8MCZzeckFptZCSgN5lB9KijRP5crfTGunj
qj2f0PhL8Fb2v5BMRkEZ+9k/6P+IEQMxvVvtPVDwYKdRHGhhde+pHXW92ZkyMS0U
P/+Q/s8ncZpM82M5LKriLbnS1ixZYyUveFpVVeXhKRTb4qMBvzJ56DqXOeQqQX0F
Y4G8O4WxhXGiOaHc2jWELLPEamwOHfkApPU8WGn3N/B4Y5TteEURYJI1ya/1treJ
6CNygU7SBZ46fSc668VWni1MoQkRhIyzpFKo8EVsCZvWjDPHIs03uPHKikP3oNpi
GakQFkoh1zlgNPt1OCAa+i757KWvY6+8lsPhgIl57Wlv18vOM3DuoaLsLbzDty2A
mwvnyhoZptxhMDvYT7TKF8wLSeB+BvCz1BnzevCfu7wqxYjP/6Bi6PtbWV75yARb
Uo/ZV4PJZtqw/QP4BBh8mYUrLx5fodX1HpIOke/Gmd3iSeNakoCLkREcJAAPLU7m
YlZTwvatTnRna9IAITru/BSvoZezcDCTo9VBPMkOboRA35QDMMVPCF+2u+rkWAdr
TU20geuseb2gLP1G0WrlHKyu+nXqrfgpDjv2JphjmYU0/FLD0SS9lRVkR1U/s+yt
tJ4Y+PFQPZqqKircVwoy4iu4I0jiyFKKrTDaBH5WAYSkFIJZunZ5Letj+VULQppy
Gd2n6B6zA2uKbdG4zVIent9SJ2DsFAc4nafvKQUlGRfSBxuC+733M+O4Htfa1db1
yBUU1Xvyak+YJj64U90wKcvS8PPc+xrFk0CRJC6V+wncujD/U9XrhiHGRCKaJZDH
i5lTOexog+gFRGYSYMoPw81UuQkg0dBMmDWkihd43QFm2mEVhr/ahUQ31zcbw9AV
B48rR5Nzzz+11QC2p+313hdPYFuL89aiqnNewUivNQkXpEaHDmzLB4RjyRCF/3k1
dzMuJz3Ok3SaiVPNAfbU+++r7m/sBXPa/qknHhYrtt97nsq3pTCMlJY2QpNa+XIu
ZB4ejKv1rjRilBH5fPUlHa2a3SIUBbPIBUPx6IgQLwGUpRiI+4EnTy6WPaNFHEU7
H9Bp/0pu6L5wuMsF05hbH7EHgnzGy7+FFdgik3sTnf1W7eNJcsUiSbRxbq2+khkU
de4DTJu+WtkGcXAJV0psrxyoCKt4Yx0zgWOqfWJ73soLjpF3+cfDpYUSvzkO2Maz
cz8pHdD81wXYtAgGOKTeRGn7dbH0zVZgHmHSzLacaIZGMxa4fcCEVY4s/pN4ZMgX
YaoqxoxvwcCDdVkqAKMk/wUIjm/7/DtNsQFGzuAZ0GjQyt326XjFabrZq0IeRNKi
o/UTEJLk5r3+T7dhPJzC1MsywgTC90qMURSpm1d0fd6vbHcaEA3GjLXmC2HLgi57
Ys/kdml7gwvdhJ4sxauHo7fJ60Nz+Og+Cv1lFY7AiRD9Jb9xnqRoMqAckJgJr6TK
BDZWt/UJa5qXwHkSDptdkWzuOoLAqHDlGE5A6Fo35+TNbxb/pCyg/8GyYO/3vejA
llA2dHmcvPvX0MZrp3jSHVre7tlGDv+CJLSy+Fr82gWMRSsdZntTqBMekqqc9HVH
G4gvvZtC1QWA37eebiBVwFIkiOmhWDOuQXPgGAxrFZlhj2wuUYaFAyGCr3KPZ5x1
QELHcYLez5H+qFyeGvHmcF/0krL3wN/1ZvaVT/LJ+9hj4g61Fb6YR+FTUMxBo7lU
0WvTAFuTosvXuTGBNiZ+/CO+OJW55A7Seh2xP07VNBoEl2syoXkt1PER/y47lWeS
zJK4ivqNXt9Azptt0BGWDoHPlXoMdBy10rHNVlXd0L9TNL8IPJXy0t9nl73vYjdE
3nKYPQmkGXpa881X9AMx2HlgvPkPcuEUVG82NeAffKCQ+qAnQPjzn3s5OeG1LjAB
Yp/In4I0a5rUx6PnyBulQ9XnjijRB6FumHkRavhT0o17HpaptJR43X+xceyP5WUl
RLfgOuxx4FMZ/fVRJrl7mV72Qc2WSuQe9rsS3IIdGCevoQWQGQqz88rGUlkz22IL
ZbjYlWENhg5DYUT3rZwDc3aWI94LZ6QzXBj0RD3ICqrOssZnAxmWpGh+YSuY6Jb8
3kRX5zp2keFYv9rnx/NjygdVeuzX1pvzY+/Vw9CoTGGd7V/R9M+vtnRNO98W7H37
MhinMxwILgeXSIbnzmiJgznblcmqIY+I+CLaY+z6UR6j5kh+ZhWes+3024q8VRXz
UMVBoIIqtjAA7yqxn++DaRJCvptNbZ1id59oan0yfukdFAFIQRXPN/v4NmYkl0em
A9D2NxNGKfdXQKqdJ5yWUBQM1XmqnJxI7aKAS46JRsCfXM4obzNedx/0XK9b6uKq
Rw0vTyTyzlj50iLlGsVEq8mj1skH+7yI+12CiUodByODQk1putwWEwVWKEGTNyEZ
Y84iNIBwNnU+XtuzIVf9o9QNPv2U421QnGjBt0iMvYx43RQSDRNYMahIBuHiHF34
ZCG9QPv3E/RLZrJo8HvPQaUOGayF8YW+Hv+jjXAqCbtp6/0YgcgeiBU+X34vNAbS
h2nfzXzHXEJ/pO7atvS9JEvdvaQbozfkZntR+SJkMHFMhKVAfjlytHj731+Lrmch
fsfomSgg84y6TvJXXID3JVbb3N7b8UnMxZCRt5w6j4BRfJFTRFJMmmkGPDwJ+8iO
sY8PVl1bUd9/Y1X17/DhDnBDDUbt1ADW0dPH1WaU/vo+KFRAq6fqtHHjUFCuxyTw
TUyD9gZnsZyMiyAgozYCyd5WImLH4iqlNvT7zWNwrae0x/SZ6HOO8rlIlwpm8CFg
e+lWt2tNYJYYh4JlghB4URivCbc+P5G/5NtDTaX7iGER4AJzc10Ci3tJF4wbKpes
NTcYlalqnk+Rq+pTH5IHMfWS7vUy+yERiTwYpYwLeU6gboWm4n+kBjuXF3fDmrCz
B1H94fygn9Xpr3yb52Uj1TG4iVul2UwXJbXK9qDY4dbAxYY1FXUXU3cPwsXppJ/s
aUwfKdr3VHbZbF1dnLNUD8iWYRPHlU5Ic1IzmFMUvYuA9AEAGT8qUqnYz5D4F++s
XhzEO3HS9xvDGF8796hwJkOCHTwA9YqUBFX1O6avzwrxgE7XlONYyPBBESkOMNac
s5qlFpyRVh60CAMoGSyQhPIe1rDa1Q53HFX3dsRRx55p/bTMah9pEv2mw+6aCYjI
go0zHGiGaGopWWqmLLW6OtgqFaS/ngqaD8iZgd5rBku2X4WeVdojpMtzjWb+Iha7
ZZ951uV1ZuBSLfK6Nb3vqizCqeFNjG2Hz316NNjOscZPS+9C/j9sHxce2dwfn688
ulxFUEtEJaHi2jQbKLk6/SM8lQK6IqbbJLsdZqnjQU8D0wvSNBh+Ckq2SqZWGQ4D
d4yOLzBQ1Z5NW58GL7uCqTfyXsB6n2Umev53vQnUJ2cUqVyLtzEW+r78itTpqwQy
rLKDjNKuzvuSUlYlOOqADqxm6Y9ril25Il6cLAcSsLBX64MBY7hvYCC/5t9J55H8
4XK6XrN4kjqaTiAPgWGMH1f0J642wB2QxjQBL2RJNBn9QDfEb6qPs+IBQufPEZS2
FR0cMKTud2XvBSmget9AY4ZeBEAMCdRyDw/UiFi5SBFOAHBAHO+pxLebCYWSbEMI
yUFOBfwN5h+TAuIlsv3BjVKZgBqBdsH4FiaULt4uHEHkJJvB6bvKZO3/E8VC9CNm
zjKbkZtZgpUXMeHc4ciXbFjF0ohrfU+qkIMpM+BeMhyaO4Aq3IsY8bkU0ok+U9sc
z0GdOGDaEjxTAP2nsEti4zymd8yFf/Dj8mLcxotJj4jVPhFVkeTbGyMGXYvfgJKW
unxVoniOAuIyltT8woBPphhF9nvz0uuUa1VOo5xl+gnDJ3BjUoNbJICaKbSIHjUM
iH5uFmL8VgAg00w+ObTyyDJvn1Y+uCh7SLEWgJl37uIfnUoqJFNHlx36hft4lYAf
C4DTRl2yPEWnOESRbukgn/vPbBQngNAcQktLqPnP5BX/Emu3gLD81PK4kfjGzYnJ
M12Ld35X2cbEiP5KnwHwNWOwJaDQEy0h81gXxzbixvPpQDFpHvYUjAcWtpsu9Tdz
L3CRqcGAqfmQg7Pu4Bjos0ICet3Vk2qvYx9I2sGVtn67RgvSdTeaeHAEcnzh+4Ys
bRrcZmi6uEFnahljHrGQBd4+Z3iK9f7JaF2rK8akxXrRSdhWXgi0XifC4t1Uaque
N8boM6GE+FjZhUtFCtbwilzFvTG6w4Db/mFrcnvIGQ1MXk1gkTNzl0PxeAuunJh6
lg/aejXC9vszn5xHtXg3bqHLZDKiG7hhrfvbOVcEizxY7h08znExrLe2dqJMo/fM
fyneOSVGVDcoql6Xyr0Rl4aQwIlkUvdeWAsRrwbmYvuBQSYPY1S9+ckHpomKCFul
aOioANFemAdz3usTNeWG5qXSIZbe1Rbmn9RIkj/nT3BVSq0H7ThwAhWyWqVVHXn5
4rEhegVToSOWmGpWwHuco0wA9gizGq1duhY9Tck5ARQ7q9lwXJnBJefKKV08dOLR
GY2WZf+oldnI00sEUJcpjD/8U1xjSQNcW50PyAdZW+8AlgtIp+u5bppJx64cJhJs
nOEJ5WoRCEkB1TjmZGxz9at3DzVmnrydyPkAeimPyvW8lqVq0jjl2+ZSl8eLjCFg
qQZW9EZEhzSarx5n9kWvZ0sgPp2nr8hsIcxktaJdUFzKebOyYBrHYO4rEcG1egJ3
TmHSgrBFrdueLhm37eYlbAxgtSkViT1PFd2XNs/cUv4weaSnCEnwUHJKwJ93YV7R
MOzbVfoN3cHiD8CJUYDcfmJlDoN6VJ0T3BOoXv6ZFeDt2IxzArBFGS2PNo/6C5bL
v+qHYZ30DBbgnU7XgoM9oaB4NG3LCskjjbQiBDKwiSelq2D3v53gf6G87DQiuQ+/
oXF2hKHmpkuuMFDXGy1ugTPsJTSO5qhtFnzfQ/B7Y0WeG4SBKSVdROjuXpkTd7vQ
zsLViKFUPpfNxN3Zc1t+uBmGFKB5XzxTcxxQdgdspgFWagZVxr4EMckbr7AuQnHq
n6u3gt4FkdbLzOzPaq33AC4ZDUkJl0VvT3pQqmHjNnK96WXyCCFr2uFk4uO5paGJ
fT0xM7sJHRgnAUFAg5P3WfwoHHUVtNFK8YpDD55UIifmaqRtexnoMeBs0uQeRYCO
DV29PVuYF9RKn9c8s+SSTqneekscOpQiGsvvEBfdoq7U0iP/LSYxaX0xsCEg0h3L
b4ifBVdNxzhKJQ+84I25WfTOPuozdpG4XSMyAbq69ZGZpTOBT/AxBjftTfWY5OeU
jtF1K3zC6qhQnwtT33pxnI4mfDq6QNollV46qQqovNoYmJF3eGcbvXAm60P1fvtM
0n3+oZXIhk1xA17lI5BlPB3FG37oAMd7ilAPkY3QJC8TiclwguxM6mTyi/mSo52I
IpzA/Rp5i1TtzvWiJo/zO+MWusMzOB0DF7I4sdN8QwrdCMvibJm5DrjjIquqAFHx
fa1OgIG1v+uweh0yTWUriTSfxQJ7Roo/z8tj7kPZLeSgcZA26/EENyhmt/6D4v3E
nW3aJeTmX6IH/n/ziHfdofF5NlYfTqUtBOB5tWdCDeu4GzN/c4lrnvqp+QJ/eUx/
CFacs5UwUk81XpJGD5GzUp0oNJudYG28y5CnsWOLNGD71MCQWKftn5sdhVjD3ggQ
UOTss1aI+HA0bPeWgOUZnjS1bW0oTlBjsioZi57c6WU7rWIF256ZdWi87judjKll
LTkegjk38zs3HTVRRTMWv0tXWnQA+rSwSzNWI25DNhemjd6BuqxmgyLE1NgBjlFb
rAGJW3T3EI1YJj7WEwttAfBFVZZt9ACKXFUrVXILe6ZGCxIp/INsyEfiXQXRruEp
ITvYffA21R4W0PJgSjz+J8nG007Dk/cW4TH9xJbwqWCfHQyo0hlPWknooboHID3i
VJE/Y4epePJbYqctgsamGcn10r8/dedSrPuPWw3jukkXZfS5NKnJdvCfTEwXdvHB
Ozj6TeZeyM6RgAKdK8uJnDULuj9dCReZzYAgK//oa2/hfDbLy2mbHbP9U+X/HHYH
cbljNxXEgBagolfMjPuxCxLFDCWbotD+Wd0szgxnHJiQVEqRikxzEmjjd27ZGUTv
sG/2eTCtgjHs4uN5HAcGDHQno7DxYzqQGoKSILzp1xKzppKHNaa5hKiJ/QMXG3kh
z8WgiQU0Yc0RsC93DPdDMrEAZ8WaTq8G/f/2tPxh+e6yeXyKwgyIHVbKhTdJRd3u
2HuBOO8qjNMcmE4sSxnXKWTfAuFp/6fNvxKuNc8mKsY0GXHJ4i0i/xw+bjjOCK1Y
/sSErX6frVB3R5z8PyUW8lC68dQ1tPsi7KTxKUgnIzGcv1B+aRwwc2QOfJIdnn8R
d15XRWyVo543TJRsNZhvP0toutZSzGWPJCwKWX5MlSAqZmzLMt38o7zdRlQrEdA9
TjrSpEy5qD4JGCEobo2KfT9F7uiplnPhHMevGZBnoPcllMtIddqqMVy7MT6FAU9t
NoYLFe+xev3NAq0U4JPr2GwWr5avCDMb9FPd3kzz48TzQolZPzfoQdZY8zKxX586
p//qELWdGDZgjnUL50JC4cYG3O2HVMQgvxGVJyS1E3x+EaI/EF6OoyeSlQHQWM7c
cuotQIUxY9QazRDthsZ3uesWaqkR8rmxtKJNURw5pqQ5NzcyYE8qQsgRXVyYQiFN
72fvJVpQ2aSnIE4w7TKAnQIFKf68xu6Tb+LKE+uC3tBecO/neyOWiChMqgzkjrOb
/wDQPO8MrFbCxk2sSEN35I+isk1hAOTkf9qtQ/KD3gSYWcNNGw88w/xj0gtjInc+
7i4FfabvQ/XxWXNz9ixqkrnJm40/floady0xBsLKhWi4+lndKP7Tswrmr3Ak8Quy
z45fcob9BQDw3DB7rmfdGzrHfZC97GwARgAchyw7klhNPWuXPy07s0ZQG+up0tQa
rc08iySVG1wYQw//Vxgqe9KVMwAvDZcmXZIY/r2qFaOswx85MDu835M4i7O5c/tn
mOwN4QtLCoL5VgaxLpI6e9E+80Coo+MsdsYseYX/Xig1I01Uu1jjl1c/wMT9hKvk
+nLmQAOS0LyBUOb9ahtSDx/e0CDtI0ShkTk7W//Y6KZogvejbGqovrfTFbnAlBUN
jJVqyI8n0PAb/WEXzmdyT+TaXaQsf9s2bDbRiFq2E8lHiQC2G+9knMSZDQ6+lLf4
XHryvt0CkC0Vhci1NPr5KbLQJ/psn5R8NX697uILDSAVsGj2TemVNvhhE+upVICW
oPD0OGc5Bi1W1sAMkAG0VZENGtvYvudsiX4pffQ8Cqjipk2tB6KmY7T7yDHvxfk9
ZbNa/cReBbvrmnvG9b2ZPswue3zAoV0RkpVvT8Vjlxix/0MPejlJFnTM/517X6vk
Hyt7L7AzLFBp2JB9xdv5ECsPHe5WiSGbUBpVlYXZ98a1Gk8aQwS7R9+AxH4S/L7q
mu1LKx2ddEPuMmB49VI+3S4KyxUyBtLGXhfHmrsuVmEQ4PpWOPwpQlNx6lyJRDKF
yOUbs5nXxXBPDsh7v9S1RrWCBALS6JThYj4r1IRf+NN0VGqkR7QnM6N9lgQ8w/qD
eM9X+EbRxg8szIRwuOuKKpkgPndftZhPyIvtgQt6wyuIel3IK+oJl9UB9RhVesbo
iblGfqKQfSLSYjPcP8uspqUL+aepsQ+0+4g7KPo6VgyYyBh85tuF6MoGIcKOZP/5
crewnTEku4JTuu05M5IiE+DwvjQp09XOfhtxjWPofrH3t9SrAVZGU6CepICLZzHD
U2r3o/Jw5It51YRR24yihB5iombYrV7DyUbfOw7JBTxiJOSGpb1yjZ27kpIRXcNb
4NC2niwLPTy+DECnkqveGLZPJKqooFxjot8a04yrviWZuQJ8RihlBsa+g/rMfhKH
XbucB+dRFldR60i3bWkI4Zsq7LNXtO27Nl5NewuPeIVnc+cO2P0NFQJeLWFrr60J
dnnUd9NQb8y40TYO1Vfih7/dUZ/uQrmdbmRMCtRJ7VTyR9sbsLNeIdJEYt8EE1qF
0XAMP2skWEr+lpTIsrPjHxRHkC7hbi7h6SgQgmxD3R6X+UPN+JBRTf7AZh1ToKke
/8eSTJhbgZgZyNSjopmjdxFK9c7geRSYsCHrjb/MU6ZpdbBakQwpakZrKOt37N1J
tN9Ph908so6RhbtExDW9ONuy/UCMcgK/9JoZHwN7jgvhJfJbs2XetMdpfER+ubYG
OWSznERL2HsdOuPGggGCohVseJLH5U6t0duuh03N9w7Ei7l9Iqavwj3MEdE5kFo7
204pZi9cFh5VftEERoVP4QCJZzEPTEMaNMfn7qXkRVU9YPsp675kvq4bhFSjJWjl
EPIJCHheZ3NJe044yV9Bhchzb6ioJL+jeRhf2fu1MWF4wB9CRqpNWWTjywocIfcu
liMY2DcCATzYPz4C+eE1AY8iKjRdySa7onBfhwKHu9ozc7Yeg6V3R1nFFguADZON
HbNq0AlnJUShglOTp2fQyFQvxG9jjLEdtYDXwHRrQ++uYT1ygJrjZ3ajdMVDaYGW
vYbaIo46kiZeDGwL15HsiHIhjKDdpoC/SyibPxDpeEqM9pZvveNGpdLG/rPOtror
hVrG0GuyWGJAJyXVFjWRqTKJR8WsHsRoxEOw6udX534dvWjr8l5hhjxlXOzDXfH3
erBk5OdsrhmDHhfCiyn3CJpsjaKtN3wf14Su0a1yHdhNIgAjDV0P3dI5HQVJuasq
tMt20lNPAAsgo55L6uctB+Hk1Jq4Va+ssy/8ml+4D4z9nSG8+x+S9etOBTL7Oox/
Rv9ybCT5siNPAtaEw7+gGVeo0EW7CUgyxs69fDPSHysw/8HPIQRfS10fysob8BOB
aQT2wztYXF9oiP8N35CkjupvmAQLliFqvKfXur2QGYPrFb0rvqRn2H4eFCxvdAd5
TMH1o/RbQyvxj7PBnOzwKzdIWyoC5Flp8fbrBRGA74uKiRvoS1lTjzPia2rreDR+
YypoIJcOvMmkYrVIsiW8fyKKHvXBVa0gjC9RsVQIuwLLI7voZCr+BOgSX4HQs6DX
ifK9XnYskL0ZDq2hcAafOABYFrxYm4X6F6EoJZLLCew4mLHEGgIvy/35+AuJTyGl
a8HuoQLc+XPDCxJxwldPKJULMpb2FbggDwDFZnSh8XTZEUzkE1UC2lr36NI0HEBN
GXiWl6jl24L3ziqsuwK7FCe7arrCsm4YJ68Pgc+n628c4HbHO/vYFxrsJP05sPI1
rfLtr1Zgn8bH4WCuDmf6UTvDUX2H8apkC/37DXD0m50CW5Y9HpPl4bYmBkf4+CWH
F+focGnxwZyEJkQsrB8e6a3NTDOjx9jmZwEsTD5/FM/sNc0fVMaGBvp8TNKgiuXh
0LnflaGkrnqJdskPKTEdDw5k7rcoUq8/vneSc9w+SwLV8ikXvHTHvoXHUenWYyot
TclRykUVNh7zf96zENtLZXAF40+JqCCpRBtyCSr3vpilyrK0dLr0hz215wBeSk2N
VuEcl7eBJjsEPHJX2k318Ue77gz4vc2UpnIjW5A+Rp2+JGFG/ID1nbnDT5/uL15f
O6o2qhq2LniscroFaOGygMhZovbqo5OH/fVMHH9YpGjWsZYwNEI1KHbETZzLP6FO
fFFJ2kZ+aaG+qYrZlN2nOgabCiiKncM44QlFPcCM+VLVz8MpT7XVayELeeXczLkI
pCyelqTrIbCCZlXvtq/anZf29xNhUk+1BiZ0Dlwpi1BQcVXYuI94N6quzJx/frvc
cvhKZ54LSknx3PYuZ1dmTDpMsrD1qmCTBTYczj7njFNd+lDWGGp3RBYPyhTHqPbD
HtUmMCKUMYPgMKr4DfIce1lBLfiqw41Ajf2mnmt5u9a9R3oQfBhKPY0yMObdBF3c
9Rw3U+b8WyA3CP9liD6LSS+nYBPZR5qI5Zz8KIp5bhmSd2+3mIvpJeXgcjtS2plQ
QT2BvC/zqn0CvQmzfNC/7ohF9Rs5NRGb9PHKzOcRRw+cE3lf/j5GEdZfDAqOKXkO
9krJHIYoHU6adRzUE99UUEc3+UIlASKFeZGKID7rI5H5nfzuYMbKKejyve2fH6kr
HI6UTLJAd3xbHHfaQqk2r1Sy3IeM99uamtP9WQrDeKZGywvibGtZSasdfMtZuMCO
plvfhRaRkJ74g4APtw4NauU9hde4hoohYY5bPy+Lm4TaappQIkPJBoLkwkGfaoOx
NJwtF1jiQZmuW6sjPQlsq7WGk3TRVy46v/hauHsMz+ByAheEEnIjwrmSak8TZqY7
eK2SLqUxkVzQ43OS0p3DXTaFPMHMeRloKdb7ChOkqsU91dsfElWiDze1QWtiCy47
I50JWYhPPgEoBgt9CYaPLE5KhpIX1YL4pm3F9fEOBKjCO1cZC+orVD4bs5MCPdeM
2Sc3luui9ObIZRkb3D4zzfc1vZTnYin9F36W5dsTNkz+pWaatHngYJbhiHqfbl8a
Ctpes6Pge1jndg/hYF1jcUwvVXesXfL1Fo3ACNvpt7AAP36XVtgWfnMFUIoIovmL
euqgP99gPEAhJJc0Uu/3tN/6E46WPtFn17Ak9b/UJ163tK4/ZAKbp7SMypYqaZiU
vzUoX7oS+00GD2n4RNPSKd5tb/6NRCwrJ/QHO7JmxYGv9aqncKHF9ukdJwLaBf4s
wMlwS+Kv07rMxkd7Mr8XdKOvMpjNXHP5ofJt5q7kRgTYXo4CVMs2hhr/zz4J/EPj
33lzKBlXn4pu9M47Li26pi56tClY+HV/wdevlVCX3QD2LJKM4i8mhENV0hipXe0Z
Irbs7xuVeZVhHNmYKWbQMj7wYiBpWz4TqmjmJdA3j9J/SUGxNX+gHidNwE51Piiv
LBMNiezDIECeibRGrvgBLfUdKfCb85ZvcZza/LEVuaGCFWZINKoonDHlkleYEROd
eX7umwurAgFQWHRqm9cFC9D1TAJlxHZw982G9AiENDM0ziDCbvOjtxiijq3zxatc
jVH2fQeoM9iqt7rcvohmsyQUZeDZII7RzylqvKvtqu++V16AGC1exsF4RUpE9Spl
zmnlyF3x0G3WJoJHabLHzj45VRyxyvqfBfv5es6xpTOKhKSPFdpZdPtD0kM5OIdj
fKj/X0olmp9r2KcdhqxulEQV00PLcj4+Mt7pQkcKyrejE+2775/QQnGwyERI7atf
5c6JQzvNybLGA6ciuWC2e/ieJUafjbpU7OLMSnqZpkoBwuldmqgWA8yyTxIYAhRf
mitODkKtQpaFRTS72YzwjtFngSoIxUlaeAColfY0vpxMOboT/WcRRXGR640GF+WA
e6J+fhZCe5RAFnv5PL+AhfEvwnD29q2xD31WVEkw7EYErvhfLGPqNMGTYEXaSlg4
IHSXXigJS/syWVSmbF2En0mJZpIYRFnQIgZwQan8PemYrf+yG/gap7+eIo328J8W
scnooPf3kLTiyRy8l34me3QDiVZF94eliaRzF5V3YWik78UCniFtbsXe0oFafv6o
lWcaQthlbmw1lGMH4aJ5ILmzpCJpkxo01/26SVfhk0sEs1K7UfRoI6M0KQb1ghK0
6jd8TorbxkXXu67Q0z2UTsfQziULG4b6y2dHo+K0vRbYneWiiYbImmkeWsnfNIEo
GOwAnIbwe136+2CG6ULulqy5NlWOP+uB2BWGAxp3W92CiYUtReebHn5dzRUtxTkN
VHKGJjA0c+1mkST1D7mZOggeAPLLv421rv3wMx9qPhcS3eVMJBXp7Ud5EFagW0cL
ROSEDb8Xf9Es8hlzSQq7/qjnALch3py+MSqj99CrKG5tGfks+UYdEXexmtdvAysW
W0xZUhaANc+rjT4R/eHuLjdxnhJQ2I8sqcSuoTnnmL5lWq0UvrlwbeTExgoe22X+
d2vXKr5dY5rAj419K55JZUj3brer/qSRm5z9drWFDy+V3QdPqwiV/D+oDK+RJkCk
iHTnuKw/7C7vIriPz0uEIlB+gEWeZBPC+HahrQrGEIQTOz4Q51VFqCbpreE337Vk
1rGBnWL/E1ziJVSgQncOXylgrSZgzN1cm9W3Yj9IVfkv8ioPQaWllQc0NMncTc7g
8ZAMoQNtQJdNQ+dHBDiUxpWNsF99qPeF62pJZyTqJ1lYjQdRfd6gjdB4rbDlp1qo
15mxKym7YZCHJSQwtlErGTfT7Ebd1fJOGasJjrX/+xq6emJWjhN9Ov7Q7wMQ/eUT
t0p1owdqG6C8HLzmferyKHWaWhpfypxtBCIilGS9jebGc77T4SiNLWwx8gVxUHgY
Muv0V+9NRDM1To6szxiuSl7dECTtQlQDDUokqZwGZOqmzvgZfMzf6vALAmOsl7vQ
9r+pQcjBbMfq8XqYiwz0tP+ri3Fcpb7YI4EhkcX0ROAVsDbmbrkYqkdsIokWlI0N
WLWDdvP9NRUJhsajgID80d4X3CDfCaQVEFIJRyuKmL+h0Voc2JzBkOfFGZGjvTOR
CiwkBIkCBeciPB+whTRDMOT48/LC34dJ0zxo6NbDJuyrTAdIB6BjGv7ARcSdXGgT
PL3D0QsdsQLXrBIQPCz1la3zrTYIPr1bSGN/FdGk3aA28cqa9YxijM5dTE7ASYq6
w9Ul7yG4DWp7r/RcgGv1IYkQQtk4GtUQOlOQJUWcGqJPcBlQTgplD9mm7z8zHT0T
kY2yt8Ndxzvy6OmSSYfXPRHYhGT51i/F3RmQ3qAb7yUUlpE/CxufSl3Ce428Naji
Ezp3IsNCwHgaGU0xp/M5VxtzEDsodzMTDvimg9IVksKd0LhvF+DSNd8kE9iF83qw
/uRiYrtQLNrmi7C93p/YKq1MDPS0DwL8QTTz4sxiiF4v16ul24wooA5KxAVuKptw
lfzq2n0NUwiWUE5pp5HmbCh6WWq7Fxk3G//pryKpkOtTeBlOB1bSXvop3f4ILsLO
V9Zpa80Y+4VIobScmEfzCE8MtyNAaS4IBqOi4KWwYjCEWwx16L82JSDUWiun7INd
nP2XLipLyt2JyWLFUVYZ4iBxdTblE1D1nel4HbC5l0ZQbFx2XGY4X31D9W3jMqXS
Qe9OLkRugXUhmLSpneRB/O6wSO+0Xi4rAsFR/ppgLWDc1Yg5TQyOU+nmKztl8lVU
CcK9v13Mgb2XjnTb9gVlWUeGer1lq/DK9X/N7ILRWaGq6uTJhojtZln4eosHojgL
YaRS8zgE6IWTqMNrgJ0rxKjv0/we5Rh/g7lXa/t/SCKSI+JfqCKdkQIrfDM14NKg
Vr1uK1Voy7+QOD/wYtI3ed879pAJsjU3i5xexETvDayRMDFQVqIhaasrZ6D2ry6Z
al8On7+7LbOa7c1FXgl+WB9weMQIkEVZ+E2Exo1Xw36Sr/3FrmGs34bARo2OtFLY
/MdcHlUucxIJA/WAWsWPauIJ/tsVdNpOKBs2j6gyJya+JggSNQN7xfr2Gnbn+rYM
/IsZQxToloaf9t1q9Cvru63YdJQw2wqVntJl1Inc+6qV+3wGvBuHsf62Uc9ezwIQ
jSfgk/jecr1uxY35cFSgzqXJYiKbMJkua8dXE60/EfDJMxm2/6RvYPlt1swoFEWp
ts9BZpmVKnH85PhqeeG7Ob5CsVZuXS0NY39xNro0CE31dw6bidZbraxCuGLxybVA
z50/7RVF5OdB6YTxfJq7ow5D2yKy24E5giDPgteJzX7vOoyipHiUnpx7xHRnpF4u
75I2/WZIPpj9mE5+xyzLfQXvJ4oCPCkmE5sjaQyp5AE9SOhO4b9iDTYNzVWyQPa9
3TBGKrgehIz4SZSrP8Xc6iuJYQ7nkE0oUKj6DNxW2z/dmx/IENRG48xDsoDLGyBG
sbtp+afQ213EFnhrIVGWK+dl2WqEnJNg7f/QSCag3vqF0ROiC9EOF+vt3a+xE6sU
sdm7tOarh9GzasgdPU7AEbDa3CA5TA3hol92WdaoQvQP2TPp0jphKRxNjWI693k9
jd+bzWJK4bWxkwd1pp7wj0btWeDYBzlY8HqACIcWhp05ViplaWNH615Ds6E+OzRM
t5LNmW8f/lMhOm6iJnJY281XeUiaJ49w/dlpicriDt88hCYlhPTaN2KJFaBcb+84
EFalPgiKFO/Izo5ylmLTL1j4ve6fw7czhRkdeAV3LzJpFB4Up4POtkV6qFnho6Mm
9f+g3/ObmNs/EmjKMAKOaJ7KzxrDQMyZkc3iAIOv3ExtvtYhHCr5We2rmgvJTcpV
5yep9dnLDBoqKBTEQqsRogI6fRv5kld5MbnIzFWel19hpBC1If7c3csE835l5HVS
kln380kLTy2MLl556gH1bWepTnbazhfrq/9T6WRPxzg1v7Y440cdi8obJMYHPOxA
sQIlphgWM9R/GES2CvuewAJOhBV00wJoxUVqRas3bTeszeQI6UjfcLkHydWqolCy
NCPm/g3pAKwgH5Nrdr8fECXgruqBrieEhLb60CSoOa+dp/e7pW3A3uzkS4jKHYLO
GNY2J9OVv8ileBNnhplnADRT/BsG7SUTCsEWFXenesTkIs4m1S2Ev38/Yu1XWWGm
BhaNUdyBKzKCGGH8112eAZ7UWS861vp35tjVFw0YDx5+h4P3lQHPzd6NGnaafh4E
lsgFgd/5CGZCZ7KQt7YDN4/fhIPjAVlyyiTS2iRvKi+y0tXRtjsAa74q5qFzsprd
Fbx5ulzXaPrZOfzDVFf6LQMMtAPZ7x1uAZCb/XntBlLKgQch0VeoTONBKW2Tu5m7
YaXJGBPAawsFkbh5zOkQr61PKo7lkO/4CuADKySJso35R294UYs10u4k/2NRLhMR
qamJ2HCeJEl9779ataJRX/arBW9KaJ9i2O4FdOu5Ek3n7f1QUbRw3O1gjantbkCo
lFo34FJAzWA7FqQepOg1YdANYa7XEFM2UstvdvXQUiGUm+QfwYN18qDapdPM0k4C
KEhSuS2NEdlj8hlmWPSvwA88h/FSGJG2SB9bRovPFMNSTLzf7bAV3FOat7exT4GP
1ou9nDxw/pJfsNdRQQkBk7xXS5I8qv/AfWKE7K2OJgnn9UIPM1Y27VdExivD0Aax
yctnQX4Is+K9A2FYUiw7hkngoU3xdeUlf4xllf428oeZTGo2QPIRq//OiRlBbFEk
J+AsBsqyGr8eHaSBvOEwcteLDta1I0ss9r+tgtu0mgYiJalxPWOKDKbCf7PU5F+c
NhbkOOpcPPNTLz3i5e+bDzLhnNQWv/3Lyt5khL2o6DaLYx7OdHn2n8mP8NSWDVWb
S7fuzs62QayFi8f0SNX/h6gR7i81MQcvP56CmBHjVMYJ/6S3xDPyH3qTFiXB+u+S
dQWk/b+cHqlhTmjh4dfS8EQuWXhoZs89sykWOzbxLGTRdR1UaRyUvPHvef83qx2i
zxJuPJkmYLmQqqpDYNO30jGZAyss4TfDJLOYDcyKN98+uEz/iInxKDY7fcSdFRX0
4iVIh9+7KOMwNDBVvggWVLcRKwZs6KDXlj/UFN1svN9jXVxoy5zp4RpTSa7nPC52
J3vMeJnSGYiobyxPTNM35782s/tIND8y+0QA+UwA23mNlMOJxorfS/bs2KnL+fYY
GoEnypd2wblnsGCHytuQQ95vSEiNWpsO5eOBcCLrvdxIkIjJCLRrDEWV5996QB6f
kiWIERKYOH3u9rDE2VqZjbavTvYpUwpAu4r99JUsUDhx7t3JYQSSAbK9lnoqs1dP
G8MVte01ndkfd6fObntVPCCD5BiEkXjZ8Unb1nrJEVScwTgJI7RgcMLyKHBIHXiX
iNINez0S8tf8CsZm6jEK4ToY5i95pPGy6oQaJf2ft9zMNz7pwbR5BPmEO2kO4xvW
Xho+KmG/KYiOF9vam851wTcts9sQViDSBV0lUJeRvjClXFZRI6uCO2xb0w+9CYvh
72A+AVkl1kRTuji15QzbcqmPDRgvqE/PX+4z9CSK3CgvM+/2FfheMcvfaqjLp7zn
yJ1AfePB2YPZceT5re4XSxfxaUYtSYWzlfUYtH8M0Dy4Uwi/9J8DGbcATT0VozpX
B1sRvZzH2mTKxpHmmmbI75JNdzDSP62znDvHO465QK1t98TAFXcO3YLz9GhodVuW
+ZzGxz4rjYeIlUec0D3mYPPCRNyAzJWOxoYPkldathxukPTK6hT+HhnWubPr2W/s
JXjv+qdXn9KeXuJ0XYWqMK9X7hbgGjv+Z8RvMP9uXKYYdiIUt6t2Yz7kzNOfYINy
G5Cod6TuaREK9kwhst9ZFd/AdrIeZMfTwOpevz7wGYz3vptDbuCMOjBbfVnvbq5C
UHeXtsGuZyyH8wQKR18QMHuq8FZ4oypGGXc6qOKhSaQ4Q3xaZclBkinWHwb92gC/
tNd3ijAWRlZfzvmd9lN/58vTi2J8bKZYYXogtHDpRAI3Exu9vpYBWHumehPcRiBX
/C1euGXz5SpdoONC2aLOTMc7nWd9gS0xIJEEGaYRbz0rBExn1zJ3GiZe5RVsyAzh
Kl3V+ppBbfrGmmScebT2jinvVbNi8sBNqB/SmVC/g9qUvWjSzEIj+ACWf4rqf79P
lr02sRv8YOOZm1jomwxnsphT5NrHrhKgvky8tfDmNlxRXtR0BlAINLJrJ5iNZuPO
oqL8zp0XGzemVkaDSoXYCW+SbULU6GN2Pka7CndxzXlr7dmnkdAcr6L3vGKrrNbB
ZaZ9NB8fPmyGhTympZE/4Kx8opfKDkkUlDHI0WZJyXtX+iVVNcPgbMPKU+3+nED6
03O0LGvxg8grUvg6FQD3ZXWmpfyVnVrTZ8+Ergxy851gF00DorowveC0irdae2OJ
MaWhYUGjK/RbpMeTxRUBhzh+VhT3i5wDAsVzTeUGbFA5XYmCrS0aUTaSASVQu6gE
Vv9XzIGRMlOFzVRB6yVxNCav0fO1p/Y9LJJSegwD2lavv95mGIt5K1p3YZm1Yjqz
cr6QOiscCzkuA3l2tsz/05GyFJXgnMkWnp8UixwdWqIz7Zt3YKfHeUkzEA+BX+eK
M9RkUsWweCHp/pPhCie8iQ0ZJISU2lrCh+Nr3SvkjzHOibSac/e1/nF/K135hKtt
Y+ArD6vZPy0e0r/NRlB4r4ThysYHDhQcv1Qo2K5T78x9czqKtLQthY/Q77qDoyCi
fLqWwrIHDlmqQMu32VHTpNnYPJYTsIPmJMhDKIMAPLZWI8BQAF8MrkRCVpt1FOGQ
gH4Qefky4ioUmkaQKw2icKF8q14jCVpWQ1wWK2jFtGGG0/BOJfZLXUgIRIPBZ7Uk
tXsUnmxiIOf2wzFwVMYzaPWZkSKJu5zgXgeEx7iYG1+x1SJsObHrlWP+OW8K5GRP
TfeHIgKpLUxCipVqM3s8nMg5zLv5/gMnIzDW/8xkWo0RoeFc52yTRnr+3vItqyWC
U4C1ZWwHNwKuAIkBG1NzbJD6W2gNHdU7yhqs3j9UHIK/APa8DnyfHPjlxctll18/
QMajSHz7PV/fLBGcS1TUS1LsFpMM7c1YZawCUQrUw5SN7tCojB/LM17k8ZzF5E9f
09xqAtj3Bu4hPlrR8LGRQ3XSm7IkmFHWle1bVBmnXIhe0SsdCuEmegQXt+hrZR2v
0sNnzynh8XL0rSNCDVxDj0lPTL63wPzENP9uy6UDZlk0ZUB/vD2AuWnzXzX8lU73
8p0CbJWvkcg6hrFgJ08OYPYbncBJADjDPha/QmmDAaTDzTqj/44mIrhFrVwSXDNt
gjd+dbbyvC6MuKyQtnqeT/z8aqNgLqItr6ek48vox66ZNPagXIMk+niWcCKJ+5Cp
1nghIfNlHz+OrnOaYqlnkN7Eu4k1BWz+PHR3MfMOnH0MBgXrGL/HSZ5499B7p5Jh
u0ASaA3YcN/hLJM7zBSqY/kKB+uEGhYfErPkK3hUyr4kn+ZAM1O36ZCZWhPnXie2
lP8k0/ZEOApFQOuHTm6jd9Pnc4NFTPqsbTh5AZdi97LXuPlYxZfDZQojqcFzijtb
KZwYGbARt6BEfMfLa+tEyrfmtz2R4sNJ40++HKxeW8hO3Akn7FfjYdlkzTqp+0ch
TzsCUNfJp3PvVEyzC/VsnkLEzPtc7+WMEyRym1DWN1twD2imtujdO78isZJCbafm
WtEmGSUIbMon6m3CDyK8rzTXDV9Vmk0+rhO00aodLh89eJjY6cMlDi2XPUj6z5FB
vQI+rHdNf4mU3oHNkifrE5qwwIYFnra9fFmtTmNYBMyvjhMXdnNpuQEquk/19R8v
8ly1Za1YY/EMAbecF0AAcfKyWIlDB5/ZGw+HTjGaVlOW4lErfZlrA6HK8dw7K4ua
34dA0/DU4XDSjn1UWJl3FNESF+TXmOAxtwmf7LsrOaV10HizUg7bqeWbnaXpiqGE
BkYFi2gxpU+8Hi6URxVlB+xaMv3ZA8bbqaM25hCIUomhhsBryf1FlT9/s6JR/zjo
uU12F1M3mY3hLrDI4zT8JnQz7nMrvCEFTtgE2ryRmuRnY8x3qyjsVbG0Elf2uXC3
vwgjjCyaa+EwNiznNZa7Riy0LxaAbgWdUgS7Dbc1XrJgJTdayp7v8dHD7Wk+7+E5
kgKWI4aVBLKSQOUvbGiwbFEgAwGpZURxDeRnuEubv80DMJSCfH8YfgWmDJ0x95xb
CctclHOu7Ql1f5Kg0qEp/B3zuxzeSAOZIOcBqV8btrxfz80feCNV7y8CdWRl5S2z
+s9EFlntPxEuqhP2IPbu2ocoxbFis5mULxtKWlUfGdxdJjSRzc/BH/X8QMh7xwVr
Z8U6NiQKI9wM55MZ6xSzOUQVzEveCVbB3IvdzGkgh1Xq9SPkblwMPwJLJOt+yu6i
ZBpCRsLQQmyaXLQ+cCGNHY6YdzRcS+fnGv5kxbn5Rugfzw7MW2ulc3rzwTkxwzXJ
1s0ehodtmq4X3vl/kIQjt5Il9iREUJfVLLYtWCx2SxOpfVae8KAQgPBqMt/WL4B6
fmLc1zG/3PLuIRWzVRJPedjZFWQCd24GnHcgu6E90Vd+oy3wFWI8BAoSY70ma0NX
OJA1IKBL0fZra1U9X5X4w/WYRnH7ec/sPT3u7907UfgBNlv4/1jUcfQTmWpw8PB9
BLo0o6SX8Jf1GVWuKmwghnFhtNzT+dO++LcDTRPnXtB2rvMA/Va9T1RrBN0944R8
VNqncvMtzYfIIlRXtY8tBSaC1/key7H0v8ERuTqy8bvXO+/EvKekx9rmIP2TH/Tw
bSo4ZYqQGoL/N6NVKHqqb0eZlBIkgwZfh0UJ5xSU8cyQqJZNmNdx0o4WBaxEfzyO
uHM+IRccarWLloT8WyamYP/2o3kit/BvstO2g5FZVMuMQUaj9kGivf/SZZ5oh4qB
79K7qyLiQxxGxIednqjmUHzAM0T4KFqHE9O3jQ2Iz3pp/rXrKx1duc6a8GS0fTf4
mEjVdgMq+kaP6OEUa7pDNIr6igB3lc9K503mJd3WkhYth/iGolFRfu7t8iTSByWT
Dq6yGRSkhn1u/a0S2std2owOuqd0Sfqr2IMg6RkGQL9/pcFLZulSCaFnIYxKzf8E
uBxDzPt0/Qjw/kVR3P5IZgjahY2vCSXVmY+vzmhiJxj82/sjYIRjhknGp+XgPZQA
qPK64aabH1uqFK1+HWidp6wghbyb1sg3NgdKt7HvV4Wtc4ucBnPbsePFwVxyzAxC
EViCn6jjsMdxlE2JucYbZpFYfziIFmhwd93NzloKFElt6hyoIJ0uv9LbNfy3tv1U
5zKuAShGW/+H9dsGoVk5wChFLh0Dp2ZTKi2tCj6QfJg98ackNkvBsZ+ebM69+X8N
zLL9i5Xakux8/Y5AEDqZnuCpFKut7G/Z6nKYwNutgbYK/rmN1OZ5g1cIL3nxYWQe
T3CDjOUX+HtDCZoorACLs4YizpF9miqtLasggjSHP8qhPJLNMs/qRXEBOPontuET
1daAUUxR96r24qMOhy+B+KTc6Z6nFLsIUraMMuNx8bRy8bKc4Es5/MORv4DeCo68
BU3Pss0UUpMZvd/zj4DDu+gtbZMmmsJf2qMHa2/NXnYAF/rG6cugouWK6LwWKyM1
3+GjRIqZZ/RWepHK3eVnVAE1/oMxFJTrvkfG1MJ3wArCg3CLSfr5TyHjPVfQN/eT
KBrFbSfw7owTyzjyRKJHrp58l3LZsS7rHgs9pT6alHx/b3cwPcV/BdwM4GzFMTEw
5pASkBgRtle3T69mrbHaQeMRalC0R/scp783Yxt7nrLyrpTQbinGf87O2A1sO7LC
26bOem9JUqvFqDOZMoOLIEFnZeN1epd7T7riYp3nYDqFwVt5CCE6k9xKwcblRgBw
3TYMy1zlK75dXeNqktDVBxsVcb2S2UBznyqY1ttmdojLXopSh2Yld8tFl4VBPNs1
CRZiTg67OJv758CM9NwmA2Z/ua//8+luLq+MkkmR27uDyHVlwgh8oLO7Z3OGNiqk
/ciyQ0XRhivTs3qYsnVWlLf4IBouCNS2eGEBn5weHg7HNWi//D93XOXVSDM7MS8Y
mPtTzxVDJME0zHgXUDGQte2NsCrwBdST32YvFW0gUu7v7gLd0Kkb3yhHRZM4WePU
1gDmQ4a0gNFFUBxgufn5MfkPGvwaUxydtXTzUqW97J3bA682fIkELersCbGLo6z8
iawZzCHPPLJJECIYZ37y/YERPB79ceZPVuc5Lk/zXcPnpaj2yrgdv2JV4Nx4q3iA
oqm7670wEsvDLOYRuY1qOJREEYavMknvoj0vjrkUu+85JnwwaosR5Z6NksxekhOw
S0zXWu0h1pFwhFBeHgAHBmaSK+31Tq3v6F4Z+hhlfrr12toFMsyU8IB7Be7t6A+Y
jJtKAaMNqPKI642X9dETFnI9AnbTastN7Ep7JCRxdxcGkx3hzZcQH/ny9D7M74mW
GdruGnV79KmsM6BHB2k25U5aj1Mgp6jKrQzfahZ24pVLD0M8gkiFJgp5K8OpQ7NO
mz6ml3QHpelFdb9gQSSw+ISJQVrhKCsrh/3YqByR+DM3mIGIPtt7+KrrTQQYS051
0IIQ6HAk75PRMbQmGFZR/ajO3jmvPjUfeVLGXCvcv8Hrd2uGqgIq3fCBfa+avHhw
bdi/n6Pg0Qv8ZssbdV6PDg25frqff2az2vdjziYsSo1NBtNoD7Pb/bBqqK4PMAT2
ojAd4sRnV7hDSdAz66eDrHznzlVKqeR3sCPzIJXq95pTp47Oq9JnQEK1streUept
DUWTUDUd7PZh4xbkP2TXQqg+SPwOPRiTVPpU5y2ZAPSCgzJYI/J+sWl376Ahgq5T
f4Vz2j/GIJto/5tqqZvmWqe9wzbtvcB7hmgc2/CdsWWxPgMfAGv/Yf/RjlYeNo7f
ACmsEumLQb34nhVBA7qwsGuQhy8VCGdm/3TDdO67ciuOnYGQq3GWWU6ur5WfF0BX
eal93+K/Mf+bl7rdhbJE4wYegG5rCglUBvqt4DSh7J7snZI8zrFJ2ZcdNTi/bNI9
uC8d5dKFjOoD1rgLq89J9/epRwd6rAYwl9rpkuWL1wDx8vcMWAd4BWga70PiXxbl
Rwn/Gi1KzQkekEWe+Jjk+rtUm8P01/CKpKxAROI6Z4tUbIXBNcK7mYIBJ7aHt/K8
3MP/vatj6uuk2KCiQMOlW1xk2SKI95rZlBsNerIC7Ls04AVZHUpurJ4faFE73BQw
KW6wqughOunOnSMlWlThk5hRsOUhIyj9bE7lDjR29o2As7jAFWvvvFgLjMY271z3
f37Tb3ljubaUNWrLnnSDy1A/TAjjAllEMD9VHUOWLAKJx3L8rqGPeCmu2uERKVlB
Vd+tYkI+fjbBaSqTRUr8r5UXuq71tgektT/9LCOaT/Zr9zsuK28xGivdzArj+sBM
onc+NzonD+cfQJgkOcxxmt2ZnovF3nVthvLyzA9PoFM+o2SRnT4RKyg5hlCcDbX5
NXKs1KlXbQAfqJ3e62RCzTUn/0BIkbXIEXuzr93KLIpMIRV5pMU7X9ICblLtT5Qp
ZqbG9rihFbKpceypiaPHZ9XiU6LZq33e/8S3hulIhGX0dgDwkapIRGqet7b2Z/ra
AWszXBNyt/6Xpm5LwvgDshSMd+1ROtpivNfCIbg9PSxFNdtQtlFXy6gi8ev1HiYo
Pnz+mUgkfiHPBljNNxT5e8IzZZ10GdJ4pEU7AWEr3kXv43GrTEOezOumK25SOqLX
Ce3JaGopZzCZKiVqVwj2lax0bbVow0wd5ekUiEH3+mqFM1DLwaUp6d30IMrHGQ/c
rXyZk3PNgTaWyU9M/bD+MoEdi21/558uHgdpkOknk6t0wfrwTUnCnhMb6LNvTFOT
Zw/jIrbVRccFJ7EMK599Kr9ad98o63LDxsAEUbranUKhczPLrRxIh3RuwCcCVQ1d
ZYN6Ie51sn7Gfw4XzU2maxTz7yT2egveYDp1DEGDhFf+1m+wnSKHuJ78PxJvGQ8R
7wdG4iw8AFKws1mhe4p0GuHw6qYTntbPn7WHXH4v6vTpPQo2Xt8Zyq7VJtjT/Gn+
p7Ec4JSGhH5a24xvtUUMz424q7XaMIvqSTlB0YabBykCevU3k2GChqbAAj9aRKx4
Frbj6OiHTcJ5tM1aYpPqkUdqhs2F4ZyJ6OzW1ZGDPA5qYGweTn7NYcAaAx7qnRnJ
b8jwbBmnhK+Q6vg9V+PC11OQq+GEjkaOkQwImfPEEp4U1NYNBsGwWeQBjdfHqpSM
ke/LXYw3kDFHgA6BmCLBFRf5jK59BLcvexML6DLZyk0kL7rAynXyeq8gUGzQEhAS
X31Rofxuqngx9dgK/8K7V8vDInBZaeFH6I7QocT+4hhBtlxx9EgTTMrVekIJJ9zh
L5AKmJBoLqosZ+yOOVExO/y6PoTyI3nDuWn6101oIcWlQRE5nRtIuTRFy6OX6NRT
H0JP74a7L2Tj87nTOzaF7zB+vUS6YwU5YZjq1LgUwp3MjycT8KCfZRud3xSMjBs5
G2h+OtbwB1EbNxyUwNUkhBThtzgWDLEsdq/vv42+XPRtoTqEl+9uRt27x3x2UyNY
euWcigQfyevNLVljN1zwLbjif3sYD+waigl5AbUrA59dwXKq68f5mgmuWAfJs3XU
CFg8LHtaidJouOwqU7gFXkrPFxYowNbv+oKgxmOsFi2fnostyOZC5x1X6zmNoqnz
6LneZAIV2Cd8MPtjihVS6OazFi3cZ6JnWxjvDfVOY68HI6AD5S2LwUqZFijRWkYh
v5qm7VeFdO/ckPD7t1wZveL05ld+HAvnQfzJ34/rToo7XA+/brmK9imTHg/vtv1V
y9FKed8cBTT2PKCiV5dwqWKMfzY2Ppbh9Qw2Iq1gSpg85uCZEY5aZ2Msqr3iJtdX
KpGsoAXET9ddKRoY5D7+U7tzsEsdEpYb0YrN85Oo4HImuOjCDu3kCE8FURTsKnnz
Yz9zidY1P10qOAPh7JLrvxPm0/6Q/GdiK6Jx5vngUfD7fxRZapmmkACwKrW9WlLd
bcq5qtT7Xyu3YtbuegocXofMVC8Kft5lzGl3N5gTwqCTVgtWl5y/zh3s0PNuTe4r
IlR3Odc1DYjtECcLmRbuqtNkyba5Yv1NAY9yV3ZIV1f0vgtAKTNeJ089MFTSQla8
h+fswHsd7dbE1r9VhFiAQRHLcZq79ffX96A+IjiRvesA2kMVFjiCvgkhHNcNZyCl
NCnJ0QhXgFxu6QqO9DMhl6xeBY8G1o7iGKDtyUNRfsa0NlGNoY0GGyWWi1Rh5aeO
VqJhRc5mxM38Gn391PlsT+1tZfl42PF4ZTMP/BY+JyJjdnQcGHQxY336SPwGqUQd
m4pNNGROUtPCLTMAO8tVxXx0xlLdkZUKnNLNLVZ7GDrVbW0qBJ45LvU4LerVzhXG
+BG9YepB3M0qt8uz4bgcNlQmxdviTtTAjXBXTONSMOfXIX9QGtuPfaTbrmmITzXG
ipxjPdQx56j2X7S9h6KSBNMlE3bZlYRjVj7BN2oUg74o63ScDX9aZWWw/ubAvc7q
wJHGQAmVEu79Ko2oS04fBFuqyXbUdovXAz5ZzxaRQ3bk1h+N5b3U3nlNPhH7OS80
Pusfyr70mWPONc8JWPW0rFeZIz2rwSqo/IrDcyCgOiboQPpaKtEYPgE0hUqaocEi
j2oakZftohdA+lsUodIF5G7dUPkfh6XnhT0UCrJVTaZRzeAE1DfLwPIoB1LgLYs2
Xj1oehwhgHLINVoqbjO6NMjC/5Xg3qKYQaUd492z7e2yuLYWJ1PGbhncQeKBc2g7
anStSKQn9CKCftb8kqspsKE5eDgmrx8bqtjz8pUYIbQgt6ztHVMgFdKwAylRFE0z
SY5LOTM/v+BhH7C4zLbd2V6ZxhNls44tnTOERsbnDfnmh4A6YH6/9s5fTVsvWlUI
j9Axz0FvSfdW6jQEJ7180FWKCPgZNXSlnrcHQgKl8GRYK31n8ccM7CTmAX17MDjU
HRqqyQiv0PGZHoUJQcW9K8Mou0OJbFQYwwVpUU3sffOG2uR6YZmoL0n/R2Tdvthk
E8KycTJlMWw7uvRSPkyW6remlPz/r2ctXN1/VrAAj6npn98k30wh3VIV0dfOZ8u4
V0zI4jF7NTtqdRr6N0aeywNy+R3C4OSo1VkXLt+v0wu7eWF75WuD4Fs3rWyF368Q
RJSk9iwFUNJQr1VLuvZ2yssWYs/YYu5q5zwyR81n+b+82SR2PZGUx7Abnz4GlXMv
P/uXvslDgrK34tYedWcIkjUndZLVXP91mt72edGr3Ato+/S6mNC+jwFpFjB7k0D0
m/pT3bTj4/Ip01Vj4pxFmQPVPZRHOvB/U4zVf63Vlq6XMk2qIHyJJ7tOfNz3jbeb
3JA4UrV03zN/k2RrJUHiRBinyR2J7/Pa5Fhz6s+KADSrQ6euitWStWQ2RNdvF3d1
BxDcyxTk/8WDo526wAJYTBZHXdn15dQHQl/AiBvWrVBOqopKu27o1d/wSc8Z6cnv
+Gr7dFjsUqASBQoGLcYwtKO2YWrs+Uqy73srRomHUQUS7Q0Po0SPZZj+9BSOx1La
cX414Y38YEGS4gi/3mzScuYZ6L06jbySCNRRI1l7YC35VQVLfae+AAu1U8OKZDON
plkcCwa+BESev0oa8q//iLs+ivjM55T+VR206C+zpQ9vuxkF5ATshjE6BsTq5GqJ
3rcojrr8ZysqJw3M27qFm0/uH3oOhwu2e1acZAeKqQVSeGCI2n6FuvEacMveRdBe
07hQOmQzdbRJR1JQFEBSoaY2ao5lUsRl3t9MsM+pfOhlqCQMexNSrwB/YoLPhOJ0
0K3qW7xFqiWA4JKJyYtoUwS3RBZ7CUaWl/OZqWfCPDyQLEgtJIRBt9DNxRPKfaCK
THzkhnKj2Cxj/01GJO5ujJkTuPQPy6cYxMFNS9ttyd/GskpVx07UBbvNnyNdO1Yw
N7xT1+uhK8kZYprzjsoNSkWXUdVn/23d5g2yBdjxMtIEMQJy4PizDFmR2UCf86Vg
iQeYvJyFIyNWO75oDuov/tNiWZrmLA520J2grjyg9cvawdH6dEnpXfbJ2JvE9jcT
YlOaVBYwmP0vcOCE4ytMt44xRvq4WasYTmT0hHxuvyEerQqwwCnPw5SiXTtR8Yk6
kn8Y9N9F778ibSD2AYa/lBMcsVhj8jbb9MzWJVvtovJbntsn6oIQVEsfwTaHxTkR
1UtIqxo/WNtimxuAe/Ro02NKB1Zat3rz0jbBoIfUAGWsIsOWGqxpheS72mqseN3j
EEzEeyqdd9fGzp3d6wz22jKdkqHPDwRo1e6b5qhaADYCPtIUOguTGN1MNizGA90w
VqxOby0BOGDaXpnaPjR8r/OfcbeJblJg1uB5eUHPa0R9os//PbQbycCEG0U/9xEP
H1QvHXPcZb8LlRpibG64Bnrr7xfTTtSmsZz12Y4XBByW6i5WeryS84LSxXaeGHKk
wyQMiz57xGt84MNYRoNtJIp5qftEtA5fAtSg2ylXm6Nd0ZDOV9VgqdDBkuUz89pI
4yRXeYFyzoycPVRJXiOgnF1mn0iysodVpPKxynz0T4gWCS8LI5ViJX2rY+/FW7iO
/E2NzsJ9jyqmfAa92MIO+rmZCZxoVii70tKhKDsz79r1GL+cXtF0xTzEPwOc1jSq
FcHs64KWQdXlyisXkX9cFae5G6uTNi4VnrmbOVwTpSRVk/DTANTZ2Qoyb37ecVFw
xIQNGCXMj1b4hTQzdkXRc/FzmXc3beOOgP42O+2hwOBU9Xhxs56mdDFPWovn2VNl
jcbZedWAx2awix04QCfpWB/w0WZmgYbxw2csigH/zMH2xS4ott8+7XuPNTOf6ha/
QNpwaxlEHxsP+NrLTFuPq0Vq5J5DCMjpH5+If8mfDEi+CwxSpr75OR66gh5Q6bwh
naSSKwdexJFW3aN9fxSLEWPAB4PUeruVmrvXC7a36Q1iaL0kjBFMRnAlLppUT+Iq
6C543D7cn7UQJtNfjqwlnVaMNhH3WULNXavUNdYcCluH7N6xL+CD5EgVbMc/T+pD
7gd2ktt+6X9Y+lwvxwga4lkoFaHMvtOghzo23wcdr+1CGyMcwLl+0xAU9GUzZ5Jo
ZXAl+u6HoZcxyWfggTTT9ZPeAXoJALdo0M+RYxWN+4rCYjaTtE+Zb+IAzxJ3Aqh2
w8oUverQ3Tqt0aKuqPepFfwnks2CoZUgB2reZMYQ6XEeQSp1iZbp4htUeIkw76Vy
jTRLVeC5DsD5GN/ly3xZMAjSOospKcW4oOqAjjBPY6PpEFMMEn6dO1TOIamPJ89n
Jh4jP64Ju/Q2kLcia048brnIkqJwXxNjTrbFvpMq5dNDsEaO6g40GpWmzYPb7WWZ
GTD1B60Y4TpWecL1M+CTTiOUkHUT+TReYSvlo8oS469NnARJJu4xgo9jtgusa9lP
0DvV9+SRMoXOK2XssMe9giOSeJlSiZlQ2Oiv6j+2wzQeYjZHeqSbp6cS4ruC7ijD
vnq/KHwFsS9mJwlE65HCT/TyuAvg3th10osot26VQlSYZx2BeCbPU10/Rdzwa/5c
XeoNBqXeUe8dsLTL/EklyDUu9fermf56zzbmHz8cQLZKzvWZ913fisDtIXTEG8G8
j8hjUJ7WfPeGAF/8KAn09T5F3tH7RCIhCF4rQ6g9tuzl+A4GYTZlC9GU4TRdbliU
twjiIaALv/WMcjs1wHIlSzx0pRMmkIcbCmcbElYHyPWB+MucMsTPHtkiBT9b8RJm
9xAFSUo2YztdduELx08LWqH4O3dPZx33ruSdkVHOyVBiL+u65RCYGSxR4JTvJvvD
TnMcLLBamJx2ypxFqjSLMNRdL611rBlmLE8sBwv9l/dr/6YewIK7eJfOloNSBV4x
6bFCDaGBaiu6wdfZfOaqyuXz6zUrYjYUIOE5QeviI6C7f7zqa69/ww8EP7FZyeSZ
GtxRaaDY2hlcku9eqz9qvc25EM3y0Xm5cPmyutsJX8JaiMqGuLqivA/SIHRsvJcI
r90DEO7MmPbbHaIrlpjb8JsmWQPikgesg2lbSUnwGoF0ICkLSqQ7AJkJ3AHMbS1y
I3VreSJN+mGBlc5xDNDRzKLWZ+reNuog1DjP9LGLGANydMjSJ0yNRwg4bdT0+kWt
eZ1U04m3oO1Zyw3Fij2SU1Tnz5u7V0G0G3T0ePP+n24tbr9pM+IFPBZdmELF1aW0
7t5YzrWO1/1DUOblw0OqFx798pkcK7j30dfoZDQM2IPgHXhkh7W8qoY4IypLfq+p
1QC276/qgThkEnSzbV2dlFeZOeSHSx/b9RIKtwm9HtS7fjeArUB9mcGC8uaqKZ8Z
m+Gj4W+0reb4h6W/zGBgZOQPJgjxesuaThHJb0r/deXpGVOpDjv6VnMpmCxEMupE
qrLshT8qDBmviFvlrAX1ISDdoiI043LPz/TmOs+OxpwnYAPIPeWqkqFzscoSu0gF
Qcla+gpy8v62fxqh+jsvEbmXsukWE8RordHyug8eY89fZRvv1iPbxHtkDZFWcx2H
dnWwSF4UQoFqIlr8NeWPCKdVUryABLuZ8EcK/n4GCZGWxm5Df/6YQGR4zjyBCC09
hq/HV5UCYQSqWz5x3BgRkmPvSxGoAXwArU3ERMatpIhjFbPF/ru7nB5NBXaBlXKL
NlrJHebY7poe04TgsZAHWrebO/+9TZRQgxe/g3Ra49Douxms2ZaicglRe7fu+bPe
3vuar4aNj5ASluSsCB9QdusBY+xhiE0cH/4tUaMu/+9rrbQg54AexhE5uvrdP7G4
hawTRfyOgeeDbwExvPj97TUGFO2nhf5KUJn2tsE3SvBU3YdHJKsGW5PtLI9bxyXY
EAj2YD/Gj5HzE0iesSpLdP1movm12ShfJU7+IGIgGjFg97GViEJpXa19bzVJ2VNZ
nY+HiU3eaXTn+R5APC7VpGJIQTrdj+7/TTZUY15ZZhW2Sx/VVJeYy32DFG9J7Ubp
gcKN0l94z1S8ZdgGWL8qnOMD0itvtlGvhoxFTeVO7wdU0eYitAMktnrTnLcy3MIS
w2aOO/2CHVOB/Qq4aVBotXWbwwTSC9FaAXxKN4xdrR/+mqarETPifXULIr6I+g5L
DoE97C6Boer7Rf/GjPjeflTkf7Sf4O9iOQF9a7oM9XYIUWnA2Dk31+At/tl48xP3
kkWjVfU9ajAVea4EvqLScUBhGiIBB7BFWT+P/OeA4mf2OnlUMsxOyXbWX+i/qlSF
uxzIJHnYjMabKRL9ogAJBUBPY0+wHqlZWxV/jc6CnxRFVaT5HPCDy10Oi8Ca0uN9
m9ZK4BKXofRic555zoMYu7O7dSpMAb0nloNlOlm5/fgDiYBgi5xA/RpoVuuD+xjp
dLB+inyMIde2V+4x6Rvh7ngbAyif3Q1zl4swyAkUf0+ZE2Lf4RYXePMN6e32Y66V
uEZxGdv7qoPjyxZ03rP+Qn19Zz/4jV/Tcwk12hqrL01gXROFxU8keZFiS+/zXX7+
vgMaZDOzoWbTS/G85FSYlI+ajAsb3/eUdVWqF1mabzNyV0MpVQ55toosHh02cmXz
dn7qBg1fOjxKe45KbXjAK8kmfWBm/UM75b5+RWcKriANKUz2ylWG6TSamDvFaBi6
D8rk6VACogvORx6qur2RzfM5StEapQr17LFGEJgEp2k8mrwuzMBD1LrxzKfopPWK
QYdQeRZktk+Pm5xNEtD2rPgO5o8ma8id6GhZMFsl+fascIti1jJftgPuWT7VEVTT
S6LwNXofjCiNyMJSNntPED6L1vgsSiLMsyPogVobZy0mfbsVr/e/pNnWHZ9mkCAM
5LfLRJNG+a2ZQn+SOHQu7O9r65JE4QDp3Hp1Ip9LBFXzRQwNic/d02I1jvakCawL
0+AxE7vaw3LDth5x3cPwXz5bbCIpVxXRf9AiWgl/B1XzZ54jOVuSecwz81yjzo7a
mK/AcZlQRmNVL+oS/VprLM95VK5dBBPXfeTvZ3y1T3Mv+IpqFaeBcry29U3DeGLp
Dqybebk4B3YzZq8lulnvkVsvw/+HcB6g4IYUKaIPiDJfpfkTocKJ4NP1lo8DINyL
Uv0iv3qWpvVU2oaBz+cmmk6/PBEJz1uGxfRfXzUg03SmvaERTRcVYIsFfEXwY1CS
2Gn/ybPcTyOzAt70bGPZL6xpiLj5KFpONunPRuyznR5nh57cINny65rDGfEDTdNn
Q4WVfDeHaaOn5EmT2JhAKIcNtZFSYCjRBwsAU0BWUkSlL3ZjJvMnxAG9HDctZJZ1
6iJ7FATs2gfD1XglpLgbx9yd8GVCEvpaOlqTxGyzQqBxTm1CFM0SK3ZgNmMKnze6
6JuIiYj1vz6jEf8yBv7qGCjM5ZNs1SCLxywCLb9IfJtzGmKCabGR6KKuFqwTsi5W
domDHjNj0+PwOcse/uiKnbyESM9ZPipTxYz++snsq/Ed2MUoZbMObInx9eXN/wUE
l2daEOXNwLPnUOEEzH1pqjrDxaKE5CHZo/w087Vf2Y4UJS2N08P1zZ5joLrJByWs
/x4Ga+NPfkExeTmeV0G21oj9YkJ/7vDZKHHrBb9xKU59E6I8hUIHevMlXumSp3hw
/0ecdDn7exR+hzTbfCNadkJwmZQSh3+kwqMgp1PDC3lqHGh/7V6HNrTTP7gO7H6W
FLERPlIzqinQCRBK4HkmHoCeA3nkPrhM35EKmRfKNhs8P9QsMwCLnqyWyObHLSjj
Tw6oX9yp1z5Ai+v1OY1LMOx+rbK2PHDNPuhWp4WbrwP4pgPcYkvxqH3XknK2v8ov
Il218oJBzpkDC5NtW1kus1+vhv3PzLMZz+2dEMjhAg9bUshN/D21eRndO0onsTuJ
vdJeYn3DEtm6ixTMIgsZlMiffMyQPbfAkoCw/Xkl9sS4A5XVN5NaLdF/D7Rq4Mm3
o3puP9qQwnecabiSn7v7XDSBcSGwzWXlzI1S/IBIt2AdfMAssyzDFm59sWZ3jRs0
yl8B5M2R4167ZAD7uDiZjs4MrjMDqjFbc6aAtBZpVn3m1Y8gphCokSZiUOHA/sRH
zkVkiWYNktDcW+p+IdAFm8u1tIZ0OkTAZZ2n13OiSs6PiDGNu6A7MbSsSAK948rE
77S0YHClbyQ3I2ACPNNfidi/JYhSJhTrXc7/tGTUf6yasvik7tgvA4evoQv+of9v
mnR2u05o+Yz72+Y59o1CLZMNmjaBMDSjx95AAITQ2WCXIDKVn1oi9dRw7Wk300IT
15Rp8C0ZBSanZlkDzoZKAuSKsfXIfHKyrpjYn0fNnKbIFKceQ7dh1ehCzHVb7Abu
hqADFnag7Inw7CX2i0JxN8FSVIsVZJftctHjE6SdsXGg3Zc39nWyfC7/ENycO6dj
BQalCUvSagrGmUwPZPeSiq/mmaZvLIZPPaexsb///4XeCk5nhyLrS8N2skNJHPuu
bAB8C04VWO844Y+MGpOTjqVC3DhntY7w2P+omquoh+aHCVCcJeWiEfDAerP5f7y0
R8GGBbqUc2aggjeWpBImkIvdkcoXWlNcyEAGhH+P4O232UadnCL3MwnzhtbnRuq4
R/1MByvQIEMdFvD4Kqk28gjoAbGEj3HJWqyTX+YV8JxQy0qWQ+MDyu2QUUOicZVq
86NUOVWcuOb5LLerIv1RpBjzSrdfuHTQCGJRTFXOrLaDFmVSPS2OQRyMgkjuD372
G/xOixTlKx2KLb8fJyUv/EDaA2CQq7IKtQy1o2c53eY+LSLmOE8e2Uz/a7iJuiMD
NlSgFzGlnIM07k9djUGzMVXlm6jpZ3EUTXRVOUNUJ2FitNipYnspZF52ipeKA0o9
yxOuVLnCnrT4qZMMWYiZv/Np1iPCn5wys4kMzbB0pHnga8WV+Sjdaxnk6zm1WmAW
s7xprBiU3JLCiCrn0wqdRzst35AP4fb9IQR+OxS+B//nRSfx6BrerwCdCLjm5oIg
RWoJSQf5s/4I720kmiHai5jSmbrSJQSpbczTCT5kiaekXZF1v2IojlyHFGUxZAUy
ZtTDU5cLQRhvsWb5b/65gRCr49WK/K5nApT5TDRvUSPZZmzrFKpJuTaU4TouNqg9
AMSipJxvzwvKlYjKGVWcPtkXLSmjxm8R7OufVuWzP/sfGz8PQYYZdq9Xr0MgQpWP
9n1pN3vTm1OSh5pZK9NSFs/k8n0izICJ/5Zsw7KsNXWISSTDAJml45blyVb9d528
IGp2R5/yZUFGJBitMjdr5tj41IVJPoROH32doI27+UFzQ1Mn9vNWb93Z2CN2HB3j
BhRQslUOW4evZ9m2/zsaVinC7aGj9cfOpvlS26xHhoJvP4Wecr1IbyfIhv7xA4og
jNQoOQI71w8OskPt49QqkBp53pIFus92+xMWj+XWKM27RwftEvU5FTrFnJvfHyar
IAuMlkaY5ng/T2/t72i4UhNz+DKrAkf7LyINfhQ67od0bZY5NqWxF7QEnq9kbSNW
dkwpDHzaH3NbTdJhOacjvkfOdUr6L5bulzYl+WsCOMToroiGGHo+Z0MdSfjSwD/4
MTQdZKIERnvS5dORp3kBWvbWOeyRVuzWmc5HoiwQSLq3K/zxDJDfEAu6znPbMMDA
hIK7x6tPsCs+6OTX83nPn/aqGmxyLwfovMbKgcM1ysSW875L5aKqYRut0Fp/uDlj
klBHyvG5UeHDy2B2djy32CMZdwICT39OcC2qtnJRGEXAjGhmCTKBPGpZkPiJNy3q
QWZ0UdM+VnZr0bbE86MH6xt6CGCuB/uVSqMODlS7gRCL1sTD3FbNQ46ck+z98iYh
dIC9/hMDhJN1+6TSKvEWAKWCitef4J7D59FpxShv+EN4bjmzKwu81iUUrOY43aEL
Dk26pa7gsCgI5bbajFprsDjFAYbVz2CcvNmSrpyB8dx/mLnDqDWqapuYjv0jiJtO
1Y4INbKqOPKiXU5Y3hMsxUMk4yZwVfqTi2v0IId4ye5xDQXEyvuTOR9ZLTZ+tH+1
+bUMFmOcoRPSjFBcQoFyCxRUi5/WTFdMxF68hSg1mkOuI1X38S8crt+tzPm6nFsB
2BkUYYT4fhieOdiRlwwqDqdJ3M+Q7WnxA0pVKdcGqc5D9qj7S7ZFi+Gtc/j976uM
nF9Csi4OJ+Gh7ELuvzlJpnvZC956LSn1I9B/65y+sbZE8rRW0p4Ea/uuRIk38GIU
aDdsJEvuOnLqlQyBmzgy3WM5CsGBkAaHAXts6SYfZUIIcZ1d6N0Innhnln+41Oh9
jIYkShJh0pJ5/StVcJB3ayWrsGtgMwh/oaY/91jBXUueVoB11+Bjou6ismptvQFP
5YW2PimSvysCZxScVek5L1PlhaVa8rrMJX2iQnXfBsOVgNPcvvKI3r0cN0Fi19sd
/eNAvQ/Qsj5ltIJp+MRwa1SH2bIHA3LLukLcHMjP6V00JQEhzfrVMTkhzCPYZCjk
7iP00ftHhsHlB8NiS9RhYarHs+VLvhrUXhu41BlXQ0KjINRirjiYA7WzSD/pVcUS
1j2288QcqywV7Yp2ZqRf4k1Q4OCy5WQ8sCLnH/ZHV7pdXhlwhb/NaXYpGaYDpwik
sChZxsoDuCuW9uQOwPDX10Ebe1qbYArfF/weI8PLSetGhh9JbjrEueOin4KJNwsh
K6P89qGL0S8RhvTWkOko85TlhkSNVpF2uTRziwuLGrlxiCYCbHWX7NNPcrcAsOln
/KAq4UGPT11/k/2YAgzoxBEFwaEWlQrCN2ct7SuK+dXTtWsx3LdTncEqZl0K+DB4
KtRWpJrDkeu0fkI7tOGf2AxYEPOXMF2BoxsZeVcWiUZuS/VwyQXc9wsZ2snszVQH
FxBkoO6CxGt5ynJm8XE5i3lKmfhZ5lpiztvUwNohXxVYK+2qvsccX/t3+u22J3uE
uKiY5fJW0k/PrFHSxjShd3dDzyWQRRCRvMBqJqGs+uveaie5kyTlU5CQGNRzVbeJ
Lp33ZBwsAc1PLo5/o1Z9WZFRHWkkOlvzh/8QQWjbHl9ndQWup+/gkWAZLvL0dwrp
6JCfc5HZw/wT3wDyK056f+tHGBVujEZCCd5nPpgN1IPguA/LswEcTqlhQUzBTtWJ
BvG51ukmsWBLCZQblfVCItoQ3uRhs7zV6vq17IQuPPv8YlVhU2Lq+a4Yw+tDYaLO
YQ1vZFbIiN2k8oY8aaLUeJi7mRbqfaziZ2ts4bcS4DwQls7yO4OtL4ilGvHX3Zcx
mvNg3BSjozC9YQKxiglEFcQNtiSNNWtYd9f8Aap/M+tnU7EpEW3L6IXRRdQTS96B
vkHG0I2ZJeM2AjIYH9GrRJIcRiS77g5fE1XPWLffnScxT9by/u/z/yPATyk0qLDU
mp9Fa6PpAyUL1d3xjg5XjfvYECenJIl6pUzTk65FiJV4uAypVqtgA98TgCdIOLr/
lD7py0KWv6pONjmZszwxyGi1elv+Ca82Fs7aZpQSf+b7t5B4s6pNH2JMazaM8dbG
r1sEmlXHqmMV1f0SEPQsl9Pq5w+xTH/llhVjVJn7pRxwAO+HD9e6r6/eUXyVcL8v
ITbWElawwi0dsjpobzfiKxLoGfBfYIQfFr7xjvZQOEE7GnH/Yy3AMO3WV2wpXqdJ
8DLqqE4G9NZuKjAHAf6LRlqPWy7BBQqS3vpSAOiwxVnRVRIyQNVP6lYbJVdJpX8J
3oBkD5EuBVr3bToieNY0Zd+k+GcJEpCLGPIE6CNPo3Zv4ihqTpkmwy46becn8Ch+
8N+pc/eoQuSUWZauF1Kfnke8Kwt2Jj9W3eqGi60udMpQw+rz8GuVzmQNDSelrPOx
+hF4Rjzu2Tm42IVNRXEksuJ73OHeLLZvZ+mQH10+M7HVm/4eb2M5iQ8ZQ0Lk4tQK
pekpVyT3jVYOPR+d0NOw+EfYHSpUvEG2uH87/WQZ+lcEQ9y/zObagHQmVtYlPXoI
66Pg0uHKrwOCuiG9TjxqOve3j/99Foeg8nK0HpxA72rwP+hs92oxR4q+TChaiSu3
t+kQ1Qg+SE+S2xM5GyLsVRuFm/+dQQl0soZyO6EzRCUpWmR9kPMQbF4Pt7xwqD/9
5vTQ3nwHATo6F3cxFDq6ObakW8Pk+qbcZMHgYuc3VuvicgFyPTIik71ZANsd4+qu
hSdjmsoi1+EF1u2DMjzcr7/CykiUz1LXgH7BmxtF02H7tHFtGCViQvBGMfoUGK6z
LrwbXxchvEpxUh1cgT0NHtR6wU0KnDwGKtfuIAoEqBILVLklhiHe+qh8eolMx7Jc
S4B5v84t++pzmO0uUMk+/ye5vz/zBttkVwc8GpUfvaqyEkJymvNe61E2cg4iPXGp
RsZfDymmelgzqDwDI8LzRV2BYmu8xCN/OOHJ6OMKIXmAKuQIBKS/fE7z4BpQhsEQ
DdVTKvF+vF1R7Ie9NaBca47o5TV8SbW3pEaooKk1nif7Hu8CTW3zj6mYWxuIlJEF
r9mkiFPyczyELMXzkOKma6M9wYTxskihWHrsjNMGo60BAmZT1KmssSaD8glNGsdj
BUb5GEN93Z4UCtklnqw5SrfOCj0V5ZbdaVS+8KLt7Sd9SjLG78OcWJrIMlOBmIc1
i8QHmIu4sNsCv08+ZEkhmm7EMU7iFzUSiaz42a3s1bVWoXnFNXNp36VERKqpbhWW
nQfD7IwAAb6LRxFjlBNksyHxyY+AfKtu/A2TbxiZ+z7TTTbLUnHuDCK4uQM8XTSt
6ARg/XU0csWwHN3IQP4v23h4fN7cyMHVtkgXuTWvQ7mnrqw4X20QWVBrnF+Wg/Xd
jWfK3InD2N95rQ1wal8zXn0uy5u4xzimWs2Qvd3uXNDoRs3LehbRi830th72jcMw
QAeOAieBODwim8wRa1h1I7ndBHU6B8j3/H67UMlTcAyFOXvz0SVtDwOGQhx+GdbG
gdenRbjNI+Miy2+1kG2JDCkJguJrl4WjTe/HdoBnaQznkiQ46fxtJp3EGem35gm9
qn/3P2+WHJa7c8icu7EZYHvw8scVuHgQwAUIEn/xmJgSMMhEAfTRzEtLBoifaSg9
+6YrUqYh1gtSor9VFkMzWkmMIq2xVJbADKADelPncalX6BgrmNrAzxnOvIkiiXOM
r7W101F69LyIDw8O+R/ARxdwktFxIkurnkAA+DY8u0Y4fbhVmXwO8h9F+8eDkwCT
sE+DaDB7M+9hczdL4CXodYW7M/1V0v7c5+EyG+tjzN2ek5q2MnqvAVblDzoRH/Bz
CmRr95ZVjaAsLItL3KeZ+SwvfEuOBXaeArXNkm0ey5cfTC9W5KyVz39u65rBGhho
ajUOPPp/Ik/CMmeC5AbtwsJv/TcZNLyH5Yuaazc/ExmoJmXc5aeR5hNhJy7LqyRo
0GehhEWGLbZCZlvj7/9pZEHXJf5xe0E8sSm3x92105F8jfFTMBNbLvv3iiY9uCJi
GPdDa6eBEcOO5PO9qI1TDxVvDNe03D9xE8SMNJSjaySeZ7T/Al3JLdf1tzob2itF
e8XTZCPGem0kmBuSh12z1076yTn7Vn+P2U+u2UVt3KhkhyfG5O/uk9ruDcRUdPxq
C3SmUowR7B5gXd29bV/K2qpDyUYZLeXhiFZzh3FYiX3dNKBPmdqELTWx274AJZSP
UzWSifeGVuyTJpyZZ0KhFhWW1RUTti02c76Wtt/fH+5aP1gUqPN9/n/S0z8JEAuC
2Jqz/mfMA1eTSxJXZ5EElNSs8oauMPNHUpvK3jBmeR6Wa21K9KvRNFxXQC3GZSEM
HmOR7al2jcFOdCoWGnfqffm53jRtdi5VHjsh8HqkI9yLGUFcNapy94FpOrsNLlJc
RrW27/Cg+h9Qm1drw0/7tfOLsdu9Mhp0ysVTxSIa/AufqwjeUqL9pl6L7VVQ20Ap
vBh+kfWFpgoFU2vpQyI7AmeCmB6aYJ9ncjvmFQJ3RF0t/NcyLiD7gstQdkqAgoub
E6yegja9tnBzd3YrqIwK53EgYV4e9g6sV/Uzn1qI3Hi2vTBB0+6t7JAYAr00Fu8o
I9iUHV+rBJhPEYsbbM6s29+8F51apvlLJbmX21kS2GuOp7U/97ZSaMWurUKlCwMy
QudhlcCKo8/5zWJyYAzRefK4aw4ervaV5hxmyNNrbIk/22EuQKuFs8e9Pkdoh1BN
0wb7lsTsA9WnRZuxj6xMFPYHHvx09Iak8veJxPtzKI7oqd7g12cmgXs9osaC028S
+AfEq0NyImMKEwIQTdzxtIrmg73qDq8V/SxBTQEVKe1o2GH4XMyKSNRH6NGDVZKb
lpUUptv0yokdvnX8Rgvii6IR+h2gUSHOShUv22Afxg1uze0ki99RpUZay/Qj3mpo
B8h7k3SOPZTHpLXoFLSjAIrlubQx9PYMhIcV9xtIPD6n+OdZC8Kjt23En3bHwtgX
iyn/+r0fGvXahzndo/N+ygh8fwe4qpw8D/GNrCtpVfway/nTj8ZrKg0iI/+WBqsH
cnahRW/e3gNjpZ1FVXzy2+dauw7sCQTcIvZNrXcWQ2OvJ0u7aaQmlAra7Bute5FI
fTZOoN1Ekp7dXLh4m1bF7OS9syhPjqDRQIflL2K3apzIyaaL4P3ZXrkoLTgzuMsO
m/IAo2Vcmcx+XfOS//j16wbq9BSPkVB6VFBJnLpde5oh8zI6WHzCBhLsxiwLo9Wm
YfOrOAQGEgeB8+TOi4XPOw6pRAjAwZO+bizS7DEV4q8SgWDXbT2/GA7YtAl5uPs5
kK6STHmAc6g/6TwZasYnFf/qr7NyzwVp56bKKRdWOWZbPZ5V9M5OOnZzTQoHYMjP
figr8K1phA4qAtQOFusFCKD+XVgFL89Vg+2OXECRg2asZY8rXoKYaAbJ3G9tUH0H
NXGG5BV95GXSZfip2soPwncFL90/ac4xCVLmY2VhJ0wBngw5Yx5H+xXBoW5ny8Uq
MPcEDjs95xw8q+3nqRNkNxtTkDIdBjowuimNQ20/fVor0+sNG/ka7z/JZoR1Y0kQ
hIBm8PzbqgX3Lz7FmxXGSNolNkKpdPQWSMbrwXanR+lZysvpJ+r1f5+7hJ8dL7+6
HA+LbFvS3YFztATPfBdrUvU7CVdRjGDO3agVaqMlADJTbq9i1lkV0HsSSurbZGQd
JdRjo/rUqSeGNGUBxhhziwYyb/knli6tusqgvTMrkzO/t5+o1cs3Prrme6cqMauD
WZQqjOVeGAUmh4rTDITvROqJeMHWZA7Lt9Wde1GZLqqE3Wox4uil6vQqPhd95Wbv
Fip6zNlo3oXCP9LqTSHRNW0U0cXMjv8Jw/KDh9PaXV0qU71A3ymPRIP9yl53xjVU
ZhiyCKov7K27BPLvMjcRv757ASNDj0NkFt4A2c4rq+nWaxKMWs+BmJF53uhbge7f
sd0j1jC0AQ7BLmCySleIhJJWu2Wd6ol3pkUxYs9EV4qlVL/a8WergYUpbShQWXKZ
B1jLwUb8ziWCrnPqqIrUfJ2rVJottt981IJJDuDZgmfbhURQtx16pPqWG2KGHycY
aNAPqhZhXTArt9fhE2kMfXEcss/HzMFPmNP3enrmOIyQwPkxnh0JaUPSwOt0cucF
tonnS3+Y33QwLFffnPX6hXXs0/aC9tBLG72SNPKk6aG/gzuWbzHK23KQy9FoVGaZ
wSR55Eb987FLO0JUNrd+8mjoPSBLL7wxmXQZCnFXSSAyDDp52A7YIL4PwC0aKs32
9Z3+sr9BIeePkTF/A+V7e98vBtLa0fZh1JWMUJzpsc93PruRk9bhS4d/AFJcF+07
B6Mo6rB2mvA3tIOtCrxpwvME4Ey5W3Rqbj+tLgiFvEhLsnIGTELDBew5U/kOmvhJ
lUyq8Ch9GA9RMih9aiak1H2Mn40m7iJQdQNW3SJtZqvjDbQf4iIrtauUwm/cR6VR
EuYOHtIGjhZJFuW3XcBF+09iPg7IiL7Q5LPsDPI52fADsqTDYNtWH1nUQ3hmcxHW
QtVHt2jY424IminUOI0EXjxLPkwzzpDdDGpTUBscheeSPdzYfBYZJlCD8CrTDCkh
3XByyJKM2P14TwGLHHmT2SABDVCJ3c+fjXTw6qekFhABFCQwmFyyOm7GMkGRg4Qj
WVttc9TEDiJOL9nhyKoYAIcOmrS5okEII6wZVCH6+vOqZmIWKl3ldkLJu3ZK699m
WVBOof+30FTtRnmQouhYYMzhWvivAFXDcArQvb2/DY0CK1gCJvMfOUTW/LhEY5kh
ed7enG87ldXU7k+BUZm81ZNvvSSUNgMVD5uXx6lWxIQEVkDzy5tpaibFNraMGjgb
7hkTtPArEz6WL+DDXqu2ebZRRHTjIvPe5bX6YC2aJNv/s4Rv5IwaYEB1PsMhVxtd
Ztfa/0o0DIVRdfANSfgi/kn08rqk5TpFtHRtPg/PBOj6mXIrrpihDrh5xex4C7fF
5hA6WN+Fz+NKvvVz8uYjbFMIhtqDXnStZJSBEPxgDYSDlzwqTVXF6Cpe0Ll8Nz3n
1Z9y+RhYa7VrJGV0jy64Sz05exFkyTpDLPvwbqbQLwKdmzF2O2ZNkFmqfdlA0MNv
1ZeV3abNH8BE5+ll5a0NI9ZOCItX3OTvh3sUmHoMKFBhUVP7UKrvQYe8JoiM5nZ8
V0Z3E1K0B6o34UD8WXm9/rg6PsyRPGhsphMFcHDKz37kf+wEQbWRCkRURK/VHKbS
/Bxy2unyGXghekUtUdSLLkCGI/LrOfVTEigIFL7KfMKt3C/dxCw5+tXcEaBzv+Tm
ciBx3EFlJJqLZvtJb3bIWByYiE6V5vx/1BuAO9SRr6jSa+n0SaljQ6BxzukbVCAn
LVhX8sBI/lmkUWTwGjYCw5YTj6nZpPem6wB7ca/DA/xpO8dFPC08oyJe346S5AQH
5L+TSBdZd347ZNe2tjaoXG5zKv30NTMNmRZlRX/47K7LDjHBAY+13SCfph6PyhZi
pRPVVBkaUfkznQHGk/Nyux7bhpADALJ71iJHuKhJxPM381KNG7tme73u/mWmytN6
66i7sg60w0KBnwII/kCxnDNsgJT+yOe94dETREfRiK6R1a72EkYHq4bshcOl4RfS
2OohcqQ20ojyCqRAesZogarsDGy59B5RzGL3ESbm68jwvMhiTm2oKihupRw4xaEL
DuYfF1mWJanLwAsL14uubA2XO/brTJFzJVFXYT/bCnbC3xvtzkhzcJPGs4LfYEpt
BbLut3IQ81yK6z4YoALRJwemwSv6Xdi2AWPXCq1B/GlrKwqw571ySkMj58H7o9Jp
RS9ZeqbLp2bJrf7ILoimzNDVv9DYWS8GnVvqPfqrXYwrbyNIgu6rHuBJlKh7k00Y
m+2ITSsDK/sx03b2rjMxK2RpxMfddpWbip+59pjQ+kUJFOOqsxWeeW1zj2Pm4PY2
IzhsN19ncMT6KBeE3M64f55aoNDmqDZeHGFoUWUpkg5pV4TgkoUQcFZm/wTVKZ3w
r5vDlGqcmqYppOAyE3tUFYpz+TtUvbedCSrtBQXkdRY1a941FbUuIPb+SANW5tau
FrcAxCC9+EhqP3Pzy3dLUbZkARVqM4FNTRfGSu7BPFp92yc95y1S9JTioRZrW3Z2
uaKj1Nc8Midqk2TM0xgUyPNvbTHtXWLu4EVt5dUu4aYMwrkKCsVKFYUYRsNDBuLb
nvb4DXuOmWRm8pp5Lhu+QPY/LJxvZecZznA/UWPzHb0KQFcwLXlTtDQaivL0nfdX
WwPid2ZQxZBj3VviR8atk4tbLF1nq8G1edTYaDV/EtVcjAdQOmU7LRTP4YrH38Dd
pg9erhFvCCWs3YGACNnf3HuinERdCBNXTAm0WC07MJojXIOFfD9YZuaFPk3DdiYK
VSwoUBJggT+I+hlVezNxkzOTw8Ozs7I/zAnb/iyqEBC93dn1je+Ah7tv8m4LLhg4
FtBQnSHoiYPkrN3b8hqOFqdcpV9mITogs96qFF2RhKDq4ISPQOaQAdrXc/oSpaxx
yxqnLW/yMuFFm4MHH5BoZGM3eL9Dx7eDSR0w5GXgbobbu8wTKFEKvUA5rOEH8T8T
VyVeQhn4vLXlZrt5bQOb5y4vq7irytknCmOJusmrEePvT49ECHo8PoSJML06d8E9
iRO56iWobfH5war/6fikZ89I8fIydsUFZ51Alk3nXaCSo0MxZSpS4SZA3MMW1OK5
Dov6+jj39cGj8o5/uSaJ63g+do1d4wfExeDSPpGOAp/TafWTChRz7vWfObM6NVZ8
zosgcxP1R8CsTpuwAJy1IUAXly/gQ/5iYLMMrBmUVL/5yPwm4HvDDZEQHWHB3fAK
pMRpDHyqgRJL97I62ljBrb/p33Cy2G8Kuquhsq9TdYfxz6JGmin62lcnLjGDL5hY
iw0qkO0gQEPFd4R/LHcSDHj3lbgR1qauxu1x22OGdMoubMUTiCm7DEiX0diWeRKr
rXhUdyqCf99M/3WTNcS1jdWBTtYRD0W2Oic8lRHIWZcc2dkXBP03L9TKMOwXbY3q
IMuYvjxGKhQdpX2hX/rbMjCDmWpjWeP6Pu0yUoCiPMYUUDCQJ09m3l2wW8U5VdF3
J8SjVxqBeh9Gf6j8ung/J4dWvJ8cva4ueYrugZjwRrdwNlMEMXJrQ98BTkPiRQjJ
+HfCfY5WUGKT/ClvsUEmtLOt0Yc0y+9gXZwJNrbAkD7B5E7TfgqxmVxwsGNRRu5T
RU9W8qbf8Z9a/8u25n1Bh1zORv2gK3YmhLdpRt++vwQXrDWrwP/a8nfKvhcPABSz
l7EjCvRykU+12F9w/q57zkDfIyaUl2wTM1E5k80TeYx02hAipOlLPhQcRTGbQViL
ZHRHhNYL6rGNhGPqVDyQlD9Y1gay9dixHE7NfIEJYwqo6NlSbRVMutHWOrTPfZnF
oHMVl1sUBDMEk/s5MlJzLMmLOiCF1dmp8oNHYPJkhpO5cVjN/BVAjDAlk9nBuEb5
4uhEh3HjE/9cQF89+JRUhfOVODfHHXy1CECFRenl+TXF0rxtpLnPEF5qJwrhiHNB
GhIqVwiRbFSfX4Ypd4KW6PYLggP7MEMuHi/RNASqbXz2DsLStfxvo/Q6SByUKqBN
LLDGhksxSPT0n+Zia9ykjy95P6rQy0mlyJ4EzWl9wm54LeWZoJWvuQWMIKjo6+ym
S6tVjYq/yVWQLyfZYUlFUpSYZMbjwKakrBA2CqPvLLgr2Ieh3mRTO2jmXhiEjgjm
gTzeCi4BMIL3oB3AobywREUtfRW2wLuVUtKB9/0EUPwCZLly9RSNIkxnLwdm0Ex4
dtABzcvUBJ8a0QzrSA1sTY3fGC9pdzXCmla0qoFe7a09ViYKKiFnAsZNRNVQyxbH
Bojx1QIWQUgcbDSazwqCPHNZ3NCU0HDMOODV9KfDYen8Md4K5vX3l/hQiP7UgdW2
5r1MDZ22WeDSw/Y8gGOOSJoK05wLqo4tldZSaBIyAPFWlVStU362yRawQwPJkMml
0iIaLT8vyjZx70vpI03xVaqQvpdjQSC4A/GEzd8IqpKBl68FaA8oSHyfoNVZelBV
p0MK2r9TDVM18MPYl3ZuR0haulagRg892l4n3sm/ka8rqqq6TILlZa8rXdWPvXTT
V/5LdEo2W6lbpmAGCEnqcXrY1WPnjm+IwlJ1z/jcC5+CRN0aT/P3U++0wolabuHy
zlZ5G6pLLkdQNFBPNc1o2CJP2+SBLViddxuwvZafSnw6RfAMMitDhx62ysCICcpQ
mlKkA3GlvkpPkVuETayiuXFpY0m6bbzx9QDjg2Lsk/NLj1+UgPdzE4i0OuyhISEH
LMSnIlvZXB5r5Ztz0xYGz5M4JjSJIwZvr7ePK56bbFAw8FOQccFC0BKUOOq5W/kx
QorjY1DqZnWGXne6se6Hw4E76Q4sJTbI8Ve2bdHU5DazRzQM5axBWyg/bpbhg9PK
YI+iq6JexIkSIRNnlW2vH0XOqQsvQoTxf78VWMUWauFhDrP1x5LQzj2htqr5h4/S
sPFIYVRAu1Txd5679fuwnytAxTS2pK3GNasBgPf95nn4xj3sQPrsfSVoKJOt0EG7
/ag+OoQC++WJFFCPn8XrpOWoQ97E90+g7pAMHOmj4wNkJadGesKVzHRCEoQ8Y9Lj
BZaISvewAnRdF3SMg4kvd94mrXJC9RYLF9SzH8r/xPjeBJ4yToJxK0vUzfx00bPr
bYlridSG1D2fd1o67+g91CcEpPJn505PHaladlSuzVJdn8srFloOB+WPb6upfXvU
oWMh9Ofol8LPC7OrwFqHKCFA3GyrYlsAUQxHsT6rrv86/xv3whTAL9iACisRHMT5
QtOiqyoCO7tDPqiV0AsF3BCT0CVit4IQSorUnIrjHGCB6NyuB7A0E0/FCeeiwmk7
JGHS834+0Zo+CXgr22hUE2JA37gxwlplyqV2s4/6jsBxiHl/TKYzikhD3yIynKpP
hJbOmt2R8N0afQDivCJhapO0qje/F2p2Zk0UPNOG6xGlwQp6frJ/Jr/czWQouIsH
1NqyXW199Y12xtm8eHbsRmTJKShEW9Gjccs0GyPBRfp/X6YLtZtsOjoLZuBYNuER
QJ831L4Ju4JjGRCL1JAvoY36UUSfjAXsiewfLAYNxC+TUZIG1sLj4NC+zG8h/eXP
4DY6VbZB+lzB0+YcotvEZZwFwPU/8FPXZUjR26g0wiZS6cyRb0o6S07VnRid/GOB
yIEotrdujQWqE3Dy3d/lm2U2Ge4ip8/YhYVYrap1VNsy6yqS+p0cplxz/VVBC5dc
4DtYKr/j5RuQHK7PiZoiDZTD/kL+OBP5HEo27qXdXFZxmmnpcZQEquhxwprKKlhd
VR1i5cQqDPNEtuVD/Ym8/v2yAeq9hcB74G99StLMaOFFMmw4uQzW77LPy1+ASlp2
GvO7HAp/uvcABbQKykuRIhgpPasPX2FKRysWGT0+dy7SmzWVKqf+rs0imL0vJ+fe
kA72BE02YY7dr/d6He9WpXj8OYYgDdTpfI2ikmEyqcOlNtB8J86wVxOTtl6F+oY6
FIj3SKAfS+lZUGbpuFeureCLN2kpWIzKuiFmVBv2gNAuT/ukrIFy1elJRfXN482u
w8FEW1X0VDWnnv18JQs+nMnvQl7Zll9cbwbhb/U8iFaZPb+LU0puSLe+KM8XYmD1
g3Wxad4zKQA/CbjydoF3Y5p/GUXViYvURW8TfBRQDW/c5cvNkuDLffhPTz/EjlJy
9S8B9zTqC3arwzkQrLwIqC4ffUdRu9bKJ4NqCmadJPut5Rk0X1ZeNtaMYda2DiPQ
Mwy8TuUtmtCRqE8dtSFuLr8rCojC5KpbRUjSCBBEqQf1kzMwtTg467lFdy8OQHN9
8cAc1PHK4in/9Lgv9yeI7hNXY/6ubLZjoZYi+jJAw7elLP0IdPwHUkYr3ZrYSRRl
aRaRMx94Za1YHs/pP0A9RjGGqx2Bcve1HNmb68z6Ctqa1ciUj8vHiZKAb+mJ89lk
IIgyr5Gl57zsRjO3+rOFUxJOEFjBdz/lZpyq9exWE5gBoBIc8BN/aE8JYTudfnzd
WM+QQzbCH1ojPQhDaOvpXNhnBIYy2xGfziQOT6hGhZqSyE2UET1Ax+Osk+X0V0AX
lTjRndTWJbTAsAyEIdrheaQ0w25ZewFHeTodYIc3xcZGRsg7Vwqe69+WuLEtrT5j
uBNYU5dI+eZTu/d6nYfo8RU27DDQCkNsZQvlUm5c8qfaJ4tYJbFwwuCc4wGOy20L
WtavbPTuGRJYsDaDnHxFvJ4RuuFYga2Jpl1Fkz27q+iFcxPNrSj4VnDtZTChBeo2
tNqfo2E1YYy8Pw+s3HFHOr7QMe0fK3Ce3n9wfJK2F242lVNK3LIqSSZ8bLi932ph
n7oR3zm/ACPPfrbN/lacaMKE/now+LZBYFBQJ0sgj9ImRf0lXFPhAqprQsd0ZzMu
8GhVZRekKa9dwmdjS1jxWnWStXnuRX6Y2GGoGAccRgKp8TJNTh96vQF0hp8VeveB
KixJZ3x5krVNjJ63DO0F5sgoIWdrC1y8PK1Smoy33TQL7TIkCo9cPqMUc8fyOHd0
ZlEgBtQ4uoqP+suSxOEnDyi5ziGqJgXC/xfN06CXAaLZwkpiF5OUr9FKQ2CJtKt8
oZfn/Brv/HPG647EUxM1+o2IhdxE2A17CYJ2ZbZlx7qNo8uQgYA6JLeF+fILJtmT
ousNXQQ74Y8gxZ3p+jVPIGo7VhV1OgCdTbdT29b43EHR31wAqI86XPd/pHIERRzn
UHukZYyWFNZ2xV3lLEk8+mYm0O5w9EAosLxiDsRWYOv0OWsIUywzAE9FmvRimOrx
/ALAKlT91td/QNBjEZ/uLxLyrbB2ru6ffPIwpAlsNVU3+fLbXAUmKTJ1htNU54A7
8ksdol02CAoekjnWminYclB8G2knCcckVvLBBEr+CRS7i+gMcp8QyMgJz5B56nnz
hfcv/RRQ9TfsZMjcL3oXtPlKel/NvlTUelilo2BJnjJamoLOftZJKcH6t9LwXgpW
zv1hPWP4nAPmeyrexSLFt8Ci+MFNvXFimtpSA+0GilG+L6b9m3ITQKMtunpuBFOY
7y/FzlcWnhpCmSN8uZuVZb3BMGPLTUDO7X+FpBFrFDZUeZvbFH+mAk57fQpjZt0e
GNfJJZSAzFYYibmCedyHQTqycwHLwUAN9GBfg7nOuaml20/qOh51axsj2YR4T9zT
ywfHPrPHu0THHiOQWDlBlpXI2SHGDJPuXcRYTb/tFcQuLV6r1omfaeJFE8nQYTTN
1yWUS2l9N9LCbE/rF8ons6ResBozmJvXGu0AGYzySsgKyE0p8CxVnTuscmXWaMMe
w8+mjXYrcC+9RchZisRVYBksJVtBFYaGBDAnqWMNvFSCtQEzqckGYcGdgXS+Z9dV
HVmY6stYGYE8xpuoeQwVnZl64eIYVhG6s9KId3Rt4Ie/pW+FIL+lR3CBBqdaYUga
Qwo9xLVDOZEFPT7RNshGlccTfpCV62pkIAmXARWuWa7pM2MuYHTza2fcqgLg/7Os
Za/B6X83PwFh8y4giezhblqXzGjKRt9aVx2z3NHldCHZRIPGEPZfYVUjfaMHVTn1
oA6ys4cc8o2HMPIkXVlsOWCuQ+EPIG23ESev7ZPeWJ2wezc0yMLIHZZdHJ2Q+jGf
zH75aWoNZVqUAjs19whVBMiRVn0u83ljmwpu1FHadgJTtz6RQb1T2SiV9dXL9WQq
iNGMp7iAu4BWe6fr0G30TeUede9kSsF7Us5wi2xL5lCyxEoxLQ3nYzWuExYDyTen
Ow+bPld0RtNzjLoeDTn8b69/ASsoZKRzruoiawxxSGGDqo6E8u1v9O5795EBHpw1
ErNVfCy69u92ImCx+Gjt4YgBLU+z4+KAp6ZQcdyCXGUFXdir6Li4VXQBxU9FHXpM
WUzB9c6cejY2Z/Y1yTwxmVmT2dtOzh/nIdScqnat6f2454HF1641kkojV9VzyuHa
j1kqIRWj/Yl0QiF18jM+cHmdzbL50iQAbFviDTJJgT3rd6pE//+/hfG4DBeT3hDy
IRWV/P+aMcMC1p+Q5xwIk6DEMdvt7gRMl5L+6qiIqMZXpdjIDZ/3pqD+rwYOOV7c
0rhZaM47l0FVicxd6hAJpt+At2k5EKRJoZtJNcloxP+CEqXlPPrlxq1V/BnCEOa/
eOtaIUhIpCzzD8nq2KY3b83sIcV/GZTABlzFDYUgremjfMFdN4p7wEUXTZizVqDd
DI/j2+VZ2qbXjQ++mWsL20azaGSIUVocLk6jqQjYw7+j6viZT/u92VQ6d0gyH02b
xQqYsFH2ukyDOCgBhUB5W5iZSptF2+96Dg4MrJifR0Poy1S+nHsLJwWwB1sfZgC7
Va6EnQqefN2l4b8UwvPlrhpsh3ZGnFmZtsxI72QvbWkuIfNvsVM/de4uMXjPMfxj
fQZ3NhW2Un96/Uw024/Iw6h91dYVozvVg4rW0YGMmAWtx2GAXOQUC3orra0heqgz
iA48/KXKH0Lel35EF5h3OF2KWLSLE88wQ9VD3TOohTRJT4zqGMnKnEN+oNa/4bxc
BmdmFq+9oT8inlpdtuaEZsJExIBmrVm6Lszflifz7vV1ZWjBnNY5a+MASuI1OXp+
PZZq9C0AEydccgyn2TZzhF2ZNjzEUmzTmtTwX8QadYzayDMUzW+/fEWAhZFZsp6R
qpnqR9x1nJiyNVN6BcWYMJ8lfGeYDEYZ9cwPTtGLVPkbfTqnajzRpF7xl5ihmpyj
A2aDMglHzzMMoX3bJDbXxbdNQXiHPATUcXWwwlzyGtrtv1F6wTpr4Smtwk5GUnAv
2rJMdv2FMULqade61TZZyXYEwsh6DumwADGQVrtrxFjRvrGvwoNXjxn2e1Bgc4Pw
HbQFfOn/4q/xnt7MZjj9q9LRtKaj80sgd630Jn0AWs3ZHlRq+04uEOTQnPX3o/Z7
3D5/CPfmm1TMDVqvLG7mB8t5zs/7MN/Pi90Z/Rpk19k1+7uAi9W8AUaunpTGsOcj
AGdMC7H0ou+VxXVd1FR4uVKNqX8EPqaKvpCXPhz2mEnrk2NsHMIBbGy17wN3o7ZS
ASAp4Ln14JPb0mZXxHPOSyrJK1/3Vk9Lz/KAOvdj5HHFbahH1SI+Wmoks9cvSpG5
ioL2RS6k7DRAnYJ/SzI8vHI+xOm6ayNbY5KIVOCIEQAYa+QhWcx3yrLEZB9/R7d0
r1yRUAOTtvzX+ZdauKNMVrgMixgdCeZaAuwGNfx5k7gTI2lrjAMUtUboK29aASSQ
wsxUPb9fX/43b46FBxi/cDe2xGTn4TkF5DESDz4PsBJJCZIKedocnD7SmkSEDIb/
C6n9/ta78YC+kMVAPQIu5ZrlcDqLsm9tg5cc0rGinzmXurwVkFTIyVi7kepXOlrQ
R7WOd8jvGtS8kA516itXwoq+Frccyw94Fa6Y+lkp/xe8IGHQpwMX3zJAbiFNAFBh
GsCoiAqz1+DPo02QPE5c4cEqwcVtER+CWpnMGlcygNY0ve/w+1cH9CpU+X3+h+UJ
sBfq4CHifD3Xxo+4JqjzOolf2SDLCE7jsMRVA2i4HKzTB/GTloPKtRfOTcq5aH7c
djiHUjBy3FF2tnnrkbSsjP5W6UIXYcA49YY8fVricZaeZRu7XH6mI1AMgE30+/lR
dEoaKq/nYx6tXkfkjoBUdrAIZNQMUVCcTDmrVM2f9UBZd8Qnls9qCbf3VcRntjHG
8reg7V7azOHHL7OX3U58g2Q6WYtyzoCI8uXp4TC17aqwNz5nB69tCw+IpkW4xnUd
v7/N32RZAy8z+MV3j0f/gZyVNZ5ux2lfzDcYBCZs0GR6EJyVL2djKxek2RXXiVct
egfFO6O1G8nz32UeDPn0kTg1aBtg1A51Sl5YEpFa3sT0s6tONCfHGYxDXa/RE0yt
AxwHIPRt34LEV/QBFEzHJodJdc2PrilxmZaP21QWlEQ38Yhui1nSYe4ZRJ0IGwoF
lkgqBngmV/KWIdnsCDgRJI2IuuRFhFZp0zACINnDdIdzLbHzu3q4NjKZwtW4vmXQ
k9k1amh48mDbZ32HTpqC6g121uR5QcMREK7X/o8TYEZXfjMLjobEYT0T+A3MUomF
ewI0wXgobZIXKUl1IK71WOc43zYC7AO/rG9l0F3xGwGa0Gnz+UXEvl+2+QtmK9dP
KeILRhtJaNfwVDWwRLv1eKgMcYDNSk29LoOgHwDxaDdVt4qncQeefs9socyNKTym
TxB0RPrNP+TdLyqd4Ee3N4Y0FYsmtl2l09IO7Dr8v1tDGmBB7xz4eQMclmykMH3g
mWL53fn4e/MB8FpqT9fbzZYbHQjltPsipy6e36wK7iB6povBCoKVz255oTlY2v8N
T4/RcDQuBjnK7zUI0LyC+W42BFeiKIOGPAX+3OqzY5t1HQzOLW9mTgo74We0Xekb
JTArPsZkboFzKTce70IK7vkGx7kx1R8dyT0jTSJib/yAfBYKhqVA5CNHP7vQ8ZZ2
3W9I1QzJUWauEieTWqZ6y5+phxh2uMHkMBatARRh21iyx1OvyfnxxnucjE7tZHow
jon1Sg8RXNjQVcGJgi56pD7ZVs203uRyiTiDhUG/A+3Q+JcH614LZGcNGwJymGlZ
Eh/AMUW99MNKqE7/qnOAGqFWWs0eqCk/0gJPsGJBWmGkZofUgQFgD+Ne8tBDEPa2
1PxZ5vuGj+TtO6Gwqc+ymqlS22ReRc4fg5WomJTiLnSfzkeBw5UfLqEL9gv74UIY
Ytp2oW93EQZrR0D3PjngbocfHG6a0bdgNqjC7i2z8R2lWnoXBUQgAm/Mx7/jIiIk
N3mlFEyjyuoA2Hp0DDb2H0yIlzQOwbOap33h5Io8v2zJxDC/r/s4fREDyGZZagZi
ug6EWO6+aTxcRrqKfQBZDpRkQE1s+x+p9SSrH+U7oUHFDO78RaBS9PEe1D77+xMB
TiwRwShfKnXVWsqh8iauBd+gfNgeogKm5UBOnkQC9/6/466mmp2i1uMYiouF2PxZ
gvQRydsOTIWzEoEratTQ//SzdzOtOvoZj+DvGwc/EYFSt2pj9Fu9ReH3+D1ZKiOQ
wwehGNcRSc1X8qubUsNviarc3v5bHDKYUG0uIkqbTMz0XgYv1+qFJ0A47MKMzbeq
gIV97en/MRwRj5hKjYGFuCq74kWSmXT0kjJT+2FZNXXvjKmqHUEpPqgQrItKjV0n
4ez/uCmz2yrdsjpO3RuCMASetaJ8Xq2Ni6MV7QFmHgK5mGGxwDN/mPbTgXjjNa2x
FuV1Vs/u3y0qxnkRi9mwA8cm8LueGyqR+8+HnZ3zaFy7FtxD2/oXoBnr6wCYPDJK
1UV8IQdVCyW7Vd1wjZj+cF5RulAm9SAVKmQVv53/STR0xSo76q/uVad+s9QT0bTa
HXRvVA3UXqbS76QeZLVHxKsNZTUM5fNRa4wgQuMFN1DzxdkHHDOeHZbASyZ1qrMh
SEK6YuqIHK7tW8f3h8lfNRhYkZFajkLRVcd3jLdLpfkBAJ7n66moeWZ21ETIU/D0
+UQz3PuFaQ77zPCoHeTzdW8T6Yrf8uMvBGPfjTuIjApFnMIuAJqQr0zYI/y0qA9a
CZumEOie3AXFVD6jmhVvKD110Kw3iEbEQOKyY/Fx3b6bywEjgvU6kWRXgle2G0ml
AshecXLO3+0i46kzz+w0kpsJ/b8tOLfMxZd6MSPpZ1enDu5rYQ4DVuaCG+SCBwQL
RWzZYomTqFYVR8Q953KkmkN4z1Ps5LdRt5NR4cJUHl2Ne5+1YRC9FtoFXN5IB4+s
0QH5Bn20JOF/wxdMI3KAEdxjFmUbC/4YuO/YiDI1leyL/rYRJI5DciGoKqqv0kSe
EeBcPIBK5gkxsOU8IpoRUML3GtwCB7yOboSOVOMCKhvy7jcmOHbp+M/TJErNvNaJ
Ny9lzXzFxwJyvqCZiJ0wYqzV1LbU5PJ8sBvyjIudYhz+/EziXDFsXdXgJZmgeiY0
BHl/S05dl5OkO7H4io4XL4o+TbUcWrVpsB3QQ5vkAFCkz9SC1GdauaNU7lYHyl+R
VCflwR9js44LAjc5E4eOWlovT+cqGC5V9T7wJtowljRT1voTK10WZW0OKeLqB0Hs
w4Y3mkZxmZeK1BQiMJiGx6NDdEDM9bxjR+s/8du9EQmKy8YLYOwQ1SC/np2JmQtO
MXKIjF0BzahZxJBIvTyG/pIkKVSpPfcpMGDAA9AL9GD+FIdfq+cD2ISZ2e0FkgjP
5ncIz5dApXs1qkAka8b585KZ/pgcU8sRVRcSbfP1ZUa6eFoinSzdNF0FLNcKOayw
PLX2ZO8Yvv2SfQePRP24dSvgvDPxroicc2FZvsz8CKTNyBM6HWxuTABRrDr82Y+0
S7l+So9tQAP9rk8Qu6VEj4OCV6vWDcUmGYGdcjBeixvYR9nCz34xFAtGpauC6Ld6
F2bMpprExwcxpBGCLz9ZImxaTYIX9Zvo0YZW0wU4xE/51bHVw5oO+jkNYvFD1ImS
yVID1E5VfoHpfvKrx/uHEN7CvFW3619R3fNQYb9HbJngh4vgNK1ADYM+nYXkz4KC
BsVlYuCSq7qII+vZHz4IBMkKsaTGFlpuY8Or100i19mMvvM79o7sj95sjbI6TsfI
xJqCzqmzaNBxtrAfqG5R1UMHBmhoXMOluqmytHfBVq/eDSU3m5lgXc83xdKT7CgF
cfXakOZvMawBNgxEFza4xqwhxmxN31cOI4Cwn70JKAZSNM6x7f5dW5WAiUAPgEqV
kQAxKE0j/ynC+bc2hUQiTtmvT3ClQ4MV3q5F+K8IGAmEBSSa6xyeo4raRMKia8lf
HZ3jeU8UXQQmf4nRQhhxfLf97rahOLzmXVuquzHKiF++vatbNrGp9fR475qFHJyy
f4zhk4t83G5FNda5PhFVKx+gVLqS9ANGxdFdzd0UpaIhrNdC5nsh7cErTndRqW4F
nFNI1OW8VX5cIT2Son0lWn6DXpn3azw45KulxXPc5EM+7J/v7GolesmBx1gSHtuM
bXWXhDjitiuJJwGqp8HeiCUj2bmMHhyEo/l5O0lwI8bqtCVcHqN1NhbKDlGwUQjG
VICa5rDWuNoecc6eVvfGi3gR5r2YD7XAjTigz78YQJC2Pk2lhHS235RzBRCiMTKK
z9BDvHYdsL32K2qbod1m8LxZhi/WtNluSO6GJcN4OuwBrIWelqoNnaphFIQpjpay
UAR4nywEdQLj/EjaerseWXrAWkdPpEBZBUsjtBBf+q90Nb/aSP5j41QBAJesXZ6z
sWSWeQDSWQ1luzhTVi4IRPGEnmhQTLKhjl8fzm4QzbOZ0Ei10ptLk4ng4/kDzfRF
bjtoBZM4P8TZlw5ClnG1RweW4x3O/7VQTqcK/mqCtImuazMkHljIa8D3jg2/z5wg
qFSDvvMlkvTGkIKpSlIkY3y0j93ul9TzrGY6eyZ6jx5Yf2OpvZhj1z2AccyheKtL
lkmQOMhQnxJQpCbKrgOwN6KFEN5VMYSqDStrKlIXVSpWo6Pa9Yh1c7A+6HGVdU5x
xoINtoTZ7+iCkq6l9QeB0kl9MN4ED8Vh/P2Gy0+xHSDX7qNwNHcizbMQf6GjxLTA
ReGKLCONjmb+gW20SyPMMHieI0HpeF+sndszR+zuGrnt8aeLWqZ8Y9mOqlpzCJro
QVzj87oN9hf4oas+8zfJCpNv4bRUaV60hIBGQFN9d0XBCGi3uzTO1npCBfb/eTPg
pA34KlZkBhoSEJ/3u/ar2uv1yk3MQDTsYMa3MRvFL08MJwsGpTonrJPq32m6tVSt
TnfJjiXCTKk8t6WmKZUZ5DkY1MS7SIY1PxqX0RaHg4WDd1jpFUqso98HG3wf76hh
PEq30HnXcQ8IC/R+DSLkxDyy+6+yHezpuG0cxqatvQTTuub2hk1Z+RX1yLMCEx3n
FBfQpKU4HclsWf2xULkOyFOef6Lq1+7yKQkIGIm2YNHVaCKi7Kt+Dqfs1fF1Hv1Q
OIZSIp6blS8NfhwkpPuVnXvKXLTYn3Nv4PemYdNZyn6zAJk4V6LDasgPf7cjBF+i
ptPDfTLYXCQ/wQORyVzM2G1fmHoL44Ydx8l/CZvbg9Gr0jwrWoinSnRscH6RPeWd
OphtULnO8yicuhaFUTTK6FB/4PPaduqsrTPUpnACTMsql6lID6SYrShzT84U3S73
6YgPv/izXANS6qFk0rae9zRSu+fJleVEuP61BlPQhI9aF1Hpu2P5ICEIhDBl+nYb
ilk2pz3ATXLY9jlagUfmJRAUz71TR+MLXpVDJE25ZTdk8Na6Cif5EfO8+SD4sWHv
pQI4OkKHCZINTourujlhZhCNInsZiXCm1PJsW4pegshEL6QNWYY2o8PP/l0Pg8vm
Lt/dGkTm0otrjNIV7rAn4Xm+gdi9bGzX0U9KJ+mGGg7pO/mUV7znEF348e99YKDi
2iKxullHEAAEymO18voB7qU3B7uyR3cqmORR0Z0Kdqghu/mGHbKGXEyAogsrmyhT
NaYW/ZfINmk0z1/e9vNKV0kWxgYzs6fNYdDimtSyV/Dw/p615PCPG2pb+gT39eEt
5VEER5J7Wv4HX8LCb6Jg3gdpya15VC624c2IihTFEK2lsb09fzO9492hZe+alNMd
RKnmg2TkKH1FSRHgCPfHFAb00amVMg49SjUkmVTkEk9KWLZVaCwUUuWCpVeBuuMO
4uq7Ckq0RqWV97aGuX8vvdUE40/Cdo7D+zoGJISqWkou0BKkX0pWI50hkKKPGSK4
bPefDj1Yovx1zn/UPH8GNzIVNvqvgPsOtU6dBeT2GvGTmt1CtDpZG2lQV/FnKfUz
4KW151d8+BsXrHc6wiZIwh3u79TuRPBZcwkNymleSKz8KlFmqhCST/NLixcFD6Tt
V1CmagZupY9rHNTsiCN+AduLhlxqcLX+QQtN5kLqWxYfy2WjhBdG2ll1qu5VSvLD
bUJSKhy3mBFde1a4dd0Trwnmua/nE4nzO9FfeEkPDdUNidvbLJBJ2ThEYlrnaYyM
/QeZlnuk/ZfWPgkvLqs7AjjBLSP0qAOGp8EOvQ8D4SqDKvqa1pOqhmYPJCQ/xjTa
dk/3ixvFgWXKv6qicuu6oKj8X4tJkTaTJwDMPAd40pEu6y57o19kgNRqRWI0iG1E
5Ji3zWkqBsyZn+dObAJ6l1OTRpkGNPNi2X8yOoBOKy1DOxj5mEbdeqGO6GWUVpP6
GJEC0CmjsVD/VuGpoI2CzSsbamcpB4BgDEuyOohWhY6HZyWn70XfhTQa2xPC0GDp
/yvD2yCe7VWY0ME1L3ONK6gaO9u06uXKJz5lLamtc2kV4BrgL0P4q7UoRqULUC96
CRymtZHclBfylzXfr58Qxks0sRRydRDy5J7iM+3K0cVV34qYWg5qRltw2qZHqEFr
GJL9Lku8aaNOx2Ped09PZbTcj1oGCByUrw808aa9VIZZHB/5YsbC6rNDoO3fw7UA
uu+HuhcOLp/BSxr+VJShSz20ev2Nnp+8SQUhBO/L1ZoJYJCp/Ti6O4PZIF4kQL1q
vhweUrmhn/3hMkAtAoyDLBhMC6kxSzUnObveObDG5l22kYBBHCwGfIExcn28bPNH
WPkkqT5TR0fmGzFqk0qF38z47d8UWa6p85xgeAmdWQEp/XzyJ3Ujf61yPNt0N9K1
QELvuPJVwwdZGT5DG13X966vF+AKa6kh0sMoQEzTl0HMfNLU6QLzupSVzyM5RKsE
ijjm4PjV43sbFV3a+kMTba8sFJH11tvpnolAi20eKMs4bB9DefLqlq21qBlP0iS7
MCJLtucc3hky459qGrwHzCU7Yo2uzRAkk4A/kMDOkLpRdiB+Xb/GOx+2oCKO/CyN
UK18W1rfEUF/plSLgVTAu11KnEhea5nv2G07EtRZBIeFhYRhnUzEtiqK0F1C57ii
SMuzhx5ZDsMLxVZrCsn+H1ZVaosCIWOBPsQBnZ1zPobWngNM/aVpux2GR1deWEZK
aQra6iwAzMDNLasAhDNrXXZrCkowqDZyuPqVbS91O2ryrsZjQTb/y5WfLpPpOEJt
au0gWjokXjrcRPUemLhDAnN+dspXjv7ghoe03+UfjJBckS30+tll2Dyge+h7AQUm
sedwTFi31o265aEY2DnSR9JcPWuUAvpsE0p+pZmRai+Jq9TTOXyy1kwkblhz7MM8
Ewz4FrPUslToXAVPrKUtoyYoaFmjrZ1pwBWmkcoToz0jU3PbXOgTvP+QoQJEdHsB
tqzEg9GpEui+tv4p2kMkYd9QF2Z9OHcsa1qin1nfqo8X06eWAwu4JuDTDmc9Gl2e
pxAJWaFBC7iiXkPniliyDq3yWxmj6NdOdWyOBl0ts18j8gwKgD0a/MxAw4OSmrvQ
SCFWVAuHl41nIQUTss6/V+askWFQ4zimvNRHwfiIm3gsseTeFna4acKF6dfxRzMa
HarvlGWdwkWiBoRZln3Hd9vBxbxnE80VKePbbxx+p98Aisrw7A+0EEkfafzXI97H
7ZtJ1JKLM7a2MRP/jUYtvRQf+WMpVuV/EfnVOtamsAAz2qEbHKbhvtJkuPyBHNuO
T6idgN0knbnvoP9bH8f1C3UDrNpB0342krOEwNHcd3St1lYgIOJxR7kFa9V8GtL3
Q6pdKTetfcw/W8c/TCsPtyjnq/bCdKu0cYIvHkaY5PZqeAmd1+gDa/AovVjecnkJ
oMcI+Z236tna6LhSRCRw1wpBZbmbSeIKkcCrTgbjpaNbHjENKz44wkj4VyGqxGpe
wuqABrLo+PEM9GvU6CXwZQX5jwxJ51Zwqaz4Rn7ZakkWG5rMJm0gb94Mk5mCYwBo
MwBbdxANPNWzWD1K5Q0VhC4sTnhFP8q+dToBDIrvLK76Fid81357qfwdeygJOaoh
OI8wZZCQj2iwHN4y08L/sjyvDTogpHr0umfpj6FPAXE1lIwHh4qBxmjAFMqv6OHR
l6ZNgx/RCY8WtN7k7FhoSF1iyObbv55oQ/nIMqplNOlxfpIQbEc+9m259LKbGwyF
D2r5uF5iaXMJeVLOlJ7+Mzh2qOgqmc/XAqIsPLLGg9FcmgYWvjRj7hvK/USH7Iox
bZJhOKCRyYZK+iXLtx22Ax2jhXOJ15wv/DKfa9uZWZ4Se0f/NV7GgSv+MzUheQI2
PublCeaB/QfiE5TzjCkltntOe9klEDJOnubw6eHBlugBvpn9rRegPSiqRWsYCdb9
A7Lyfp88aQSRyXUxq6ng9Y3UknNAFwyvjAYq9dd9/91LmH+8uamFY18g5vbgi7PD
vKkDkhKuIAdMONscQE4bQ1h2EFlpR/XsxsmijfKOrpAT+fdqCaor51fYbguLwnqe
rUhrcIosmZc+TIZ+8pb3hlmKdFXrp6WgCoc3gmeTbJAVNByIUj+f0Pc0XejUVQYF
YnqGauWUMeqq/XxFv7mJ5QIpk4yWcO427FDfyDlBwWeLuw7Oizws84bzbGI02GDN
02h6GcLbgAsOwE7KvvQxw2PnVDI4hhSWVevek37hAVbGuORXBgeRu+weZd11Vlvt
YiYe0VuuLM+qaYDs91WzYo446vtbVUAASMWpqn3neHm/g2GXEeHN8FBu4qJrGc9g
LJ6emRiIvIPsWwFJTm+HyOJJk0E2ocuFQAtlFdnzA+vzBOOfUPhn+YpcJOSSOEvA
PKJ5/7FjtNzcQ67zpoNQp8tIs6q4qOGJVAN5+zZ2KglWCct6TAFCjzkJ+MV8b83+
Q/XZnv+PkgkcoyVTHas7BcjFugknkDv8JE77o2wx2yLFnk0F/8v6CNumSPpuLgNm
lBzxcvJbJhzwREjm7oC/cgER5zjRUNFypuvs3GgWxhJSDBcp5fAI2IthdgHDAtAw
B6k+ey6UjAi+Bt6p7gaasQBsij1GnNTpLXXBdqXm7AxsBWwvaMrNRG8u0JJNOFYO
nlfC3GrC/BMUl7PZxauqOr6IPhL1PQ1mb9+KT/fsKOeVKuKteLX/YcPp9/YjiY1H
QW/DHogFmTwi4FYI/m75fvl5VHEjlY2d4qspDXBxd7dL0UieDEul2KJalc6zDbtH
z9fatPeZe8U+VuiysqcCaRmK4LCGrz8CqwPtTVVnITM3pMB7HVrtjz8x82VbGrFz
39x0Si8zzJUY4P7F6skITL9fWe9V5PSuSohFzKBpU2Lv6qTPJdj/Zje4DD2mTy2i
VoTWRa0S9iDEpxFyZGl47eeX2kbdDmHE5QHmIAwT95a14ABhXYgXEVb8p8aJhh+R
BzWsTHWcR8g8j+vHDOcnaFw80R1/6IUvCoWCH744Kc0yMCW9eUqm5ImqIT0qq8/E
6Ukf6HSomHTUlsWi5WCp6gJYxfRvwhu8tflAsEOfYPqC6BMTms03LreWWDI5TKcY
ijgOAc3KIWMG5GB1+KwvagVZ1QOjPvRfRSDNN2umjd8Ah5AI5mjKZ/9QrpLmuD5b
YhUDXvi4kgCdt+V1pJdQ9hRac5T02txGnnmWxJbGqMjntb+LLL3BvgLMyw1VeRNw
uw3PZV+yOetdwWWQTCT6xQUhP06gdlVQ64oYO0h4fOFrULglyR/qMReAVuGkiOUN
nIwBjzO/erOjoTb6BzoHOYjMH+ytWLcUGwPFo7FVUdd0A+CAfw5ljTkFs7agfg8r
VuK9RDYDg2STqVbpQ3Rhrr3k29krqjAealdRnOUykuQsKqaDbvfLeIz3+SlJh1m4
9RnF0GLro5fWsQCXoVeyYfUYPiehpD5ek0wV4v+5vbM4Mq0+VrSHVlWswJpP2NiZ
a23SuaegnI3gZbepmQ/CCbJ3wRp6o5PzOD+LG31LG0xIuJ22XrQv+TpJP/W7lPK4
RiAWLP7kxzBP8dOCS2nz4W1tBVYT3CLNKQo1Fi7b0n8tC9dRrfpiytsHlRIl4boK
c54jeuVMRR+vEGMoAXZ4H15QmgNPaziZ+zalv8d/DwXMo2gDRdCGElK3kemFzTfD
ueqRt2VRHRutQCZ0Mpblzx/2hmVvNjF3kNnF93h0/97QdpZiwXCZrqiKny22N/kB
rbT1NRvCWmX2you4R6RmBXg6nkEOf8kvOu8DJf7XHzXfSxMEDpy9VJE9ANw5bqOX
eVrIZEP9t/bjNDsr4cC6xUhddrkTKYWRWzfl7f6+tXsVeeGCR4xyLlmAq9Eh+zJb
nt6uMLdZFjC/gfbpcAYNa48HPsyWxwhOn5A9AXgCecdQf7KidmTFbEd4VEbspdgB
bi2GCv7ICBbL4UJIVJKyCias5HAUm4aAbDt9z7y8hKVKBwUa4EqNKpifiD39RtNE
HtoCT9pVV3sYMGN0pbpAzB7KyWHM05n1BhbY+CIiwsbK+AIoNF5HKrc4o7/+EDqE
090BFaWl+shx/gf9w7uPkpZxlawdotBizMrHJBje5nicNYRFp7UXbN1HUBnACbxs
UQWx4FlJLVRwJsyfr6HM6eDpRb95XgF1+pEm1cAxiNkLAXRs2SPHwCMFxCmh9no0
nSeXkfrVNiEd4qhNcJj1oeAX2FR/vDu/DPV4gD5EkcnlB6C14jATl2ouU+FDMRTv
WiJoch9FqsniV9ouZPJR8i/htBUAfqID2O/zvOhCUiN1117TRZO3SMybYdeJ85vU
mSgyeapI4IF8x0SAr4DZLNoNAr5eG3NkKlJVIrOfLOHH34f7XrQWFU1VXXcsT5rl
imLOkrcwiZPfAZEBuff/v2HepahYNuV1a0Z2W1XicYI8sDqh8HP2IMQIGkhZIhhD
wJph3XU83z8MVKo588e7PLLmt2cvhnrEjxiT/iCwQuJtk+t4bMFJznfJR/ZWjyHs
lmjwBsBZom7raBPxf91sPKLp69uPNidkBFa9fN1A57zeVm60BCtAzmlp/lvhdH8o
NWE3FaEnnDviC1C5lkrwhgYxmYichms8Cr745Eo791lj7yUpvsinEi0kqxpWjp3U
LCO9eFMRKXpLNWRh9xD0hfP5UaWIN1l+YtVGikcBbGrhpU8nzS47LNBefX3fEJFV
n6UGn0dVZQW/CKSBeEqebf+goVlSSaqvrpiGMZlD43uvMiYcK1kMMALg8BFO9v69
+M7s/z0lcQ/MPV2Gtl01fUk5+s//tqaVPCGkPloZpcWqpPsHu4QOm0Mvd9Ml7lYJ
wqoFkihY4nX9yO6Y1BzZNK6g6q8dm0zNImsDFun+LMH28wscSratjaC10aYkxLNN
hR6Jilbc+Jbxdnt3jwx5a0dzByretSzoiToN/n1lBW8fw3P8r/0uVEDuiJTh/inc
m1IW0LAV2ZLLBECCtF5HpWVlOOM+8nHgzfteZ8+Rq+gOxbagrOKTPKo/EPeezkzX
u7lCa5/Z7mbyOpcFu13Xs2xrVWqG0xRIVnYXb+aIO2vfyAn2/2aZdLqNHxPKolLn
SeoPTiHNqgg4mwRG7WF/npU0d6wl+tRn9vrfV+ciksDgyU9TSkkbmtWH6jh5dEih
fp+YR4dFmwMGAVGXbOId+bW4xtu0Pt15Puy5XqwutEqhDmHSIk2GrgUkGX7cxlu3
ML/m1l+FJyvWUf24T0Oi8A5nW8XghIsooTv5zuBrdw+aThNR18d6/6uvNS7rRRmf
yZbBa5WK1b5oFpfbgnEjHLTKL50gHBnY/+Ti7vjKx+fiDMMk/0lrN6bWjDSrTBLi
p8QqTJ5MDUEr60DPQ2hc7wDHmoBtcCx5rVb4iSWOaTIhy4ckNjjHVP8pKOd674Xs
LvF/eUB2mC9eTa+UECk6CXRELi4wzIOYJXgXgW8FRr74jZkBruUOnblwFSOg5RbH
51svWEgg2iuNBeEnoPpSyfikO0A82FpPiI93QgwT6tbdcfmHkRM3+fJIuALPT+HU
YY8ilRm6wTKnO1rB+HGEC0J9ZMCnuPTiN/W0yweIyYhwBKQJUFO8s6e/ItEGTx8m
i0fhlkrie+4m17g8xD+o7OGeYb1k/k8HoqQDsZB89py6Ro8O5EnU6eS8+pvzwb8K
FA+Qemg4vnzrM3c58mGNf9LlFfdOrlXzthmL6VOyd2ovBR2GU0isoPXrLhwGL8gI
hh/3RPJ0lZ7kiPPdzJpcNr9ECcebJw6GgE5KudxttOiTF5KfjfjzPwCnZ2CPqdAG
spYF5kKaVNqu7aus+2zM7UrDY2zuiTueiz084v8rzn9eTfYFnI9HJk34UR99sF0r
0vr2P3XUhJgN/X4mn5Xy59TjEKIgkRUXeJjWqoEekIjXx/pOrRNqwBBC9gaWLbCV
+y5WdWnrNp2GOBaeIFCcX5pRCNfB4a5JZJxFTitpEkm2OyXt+lsDa6g1F7QOLkIB
no93pkpGFaLhD2ex2Lo+RpM/b7c0RGAyzyvjkKzApmh3WnQZWN3M8e8gyqNuldiv
az6fk0Uq/fD6FGYZqj4T9b8Fa7LmK4mBIxGhAj0FLj+9StoT3/nk+I5JgQpsgWi8
jk+kg5khllKX8fxLwNryHnVtM+cd+OMU5hIRZBztZb6CHyqRlGVOnaql+c4cUr/m
rN4XD3DIU85cp962u5PKyDn4w5vKtIgp3mC5IUlf4BRveERV938bKxtv74nOSzbp
em5sVnoZUkd6e1udCl34x9hzD4SWJUVH+iotR5a/fgszLOR3ra9ulUakZAj8ALRA
tSq1UVjYC6XFs6fYuT8kxhpnsxts/ivlOr88EcnHZ7mqHPIKrJCtRG2E89dSphpy
OWpReS7GEtfOP+S1wgJJK8Dpw82eH1wPXdGeG7p39BCJyBvYpb0s5B7cwqsL+VhS
oGxfBhTnpyxaptf9wkgspj/6osLUdQr+RgeDgJ4zJtkbxXB2tXmSzIX8RKoI1UQN
yvt2JciOcF9XHlKFlwkO+OWiSxo0aq824K7nJAXvIUq5CDwW2bj7HoIus7r5F7Wz
6obJLCyo1slWdBVPntWCprQaXNfRpGoRJP8KNu/GGjX/TuV0l+SQ0Zg/ZgaeMybX
h06MES06n9IuIycMTSURmTMffDPpTIeLReEF9uwAXJy3FCuCl3wIBzO+5Owj+vpO
JEUltQM7pEDK0zqZOWGAHYuu73EGPt7SiO+NT68DBk/OpAHRAKqAeFqr5EO8tLzB
rV02ZNRd+isO8veCb6PK5qY7Lg1+sZUU8U3ciEkljSpHHIqr28yH1Bss5w90Gkch
fKsYsPLZ/wDfkdia32tDG2aIeh2jHgk273HfQI8fpvoefhUmHBXIdK6738F7COC9
2Hm5NuqkupGwd7OB1MlrYSsPbKv2gqpXlDyOzaMWH9MDsNjyXCXwAnkS0LAcSSZc
amWt+jRHSa6GP/kvOcRspuPllQAF3Cjn9c1opYy+xHTRZOT70netDSH03sklyzyu
e7r+APUR88vLlQ7ZxIH0zsG4ieYZTI4LdcMpNwOGPAua6BOsSiZTEZBZvKDoybfN
KmLSI3Yy568DQ1Dzs192H8Tm1XBR4sgevhtAln8EWW7GzKtpMl9YWO50ZeTBsgg2
E5z7Owftx1TYMod/QFyEDA3GsN995D6ITunlIWq/GgLddNYkdypFZOuzY1glFyb6
GHWpjBWmU+QS08gjH9nsej+o2ZeXKhjqnU56W/Xfp4iQd37gT0NlAoJhnpAsU37j
PgxfBIax0kyE0Onkzpv5vTbE8pa7ncPkQ43HIFH5YWBNqvaq3pX2dpjZgRzc5UWg
fmiKG86znRV7YNVgSdjb7RHJO+tHB1JkxSdMM7b+aG0z7/MaRkx/OFPQpAlGnRgh
PaoeMIm4TZzB6aF+7S+W5pbUOP3EKE3EbGtwHfx3utZbhB6bNCj4cuXhMVz2V61C
v/RzD5B6Sam0h80q7sF9JaHAvzjPG+cOUR35pNSrtyrFY/fZZb9XSsRPPYAiSOc6
Jy0allshuLCoPrTzkyWk0FNC0XqFEhm8xrqHEY0eldk69HFOz6opftuq14akJHca
Q9G9pY+aDoIXJ/Ro3jUgXuY6soGJSARTEoPAnTXyCbp6NsmjhJug7IMq51pi/vHf
tMyU0fiVFWWLPcUXCEufglefkgr3RxFIJHxsfoMmnkNMn772LSDL7tcyPdgUsmWs
LjCY055rfnfMeEt3d51+AWu90Uh9AGSm8m++dpvW6A8YGmQIjqRNTSQwJ7ut2xbW
yOm45tOLwqCgpecsMe98YQfb6hAQPRm9n/7AYZLPWLa1/U/ZC0hDwOwpfVc/Hj33
uRKPLKa135+nn1RaIsxmu7RfenoiHq0qF6MXU7hs7novC3pn1pfSHNTqjhk1PSyf
lfDq212kLeZYW+2Bpt4XIObGhhIVnYIQ+Lu2lFllTBgNkSF+1rgr9W75lgNiMdvd
l+pDY78IY7U5aKGPrB0ZzxZcCgFfdcXm7n6+dUFVJa+XJvIfdltgU5y0hOuCzm9n
jMlLfmr858GNVZey7jI19sbtFn1CQ7gxoFij50MTjqJdlUzwHMtRC9mj5XCBGApu
6OPvAFIaaY3Cde1r29eVe/0DhK0qV0WDUpeg5VqROH4bClg/flZ+hsMtY8e00F4K
TVWXnIID741f9pYYTh58vYb/LKLXwMeljkpjEmnkePMsJ9u9VbK6jsJkVgiTmhGN
NoW4EWtHArMKVV24LI3jTcHFpQy5xL1uYxgucF1j/jGDMn9LLUrQmIYcpO1ZMx2z
ktla4UPsIr8Bu29QcHwWyG9Gvax9UHFJpoHkzDoiSZtfvApsTaYW2NbA6h//a9bq
7MVf/fjYbv1sKlel4SGmyWS8+1l9tj/oQukqahB6iFzZDt9WG3S4Ghe6i3figVZY
FpQE90ukh1t6bCb0z7XcejEhdlOFns3YSzF10c4fZxMm0nq4mUvR8KF2KteQMzW/
SYJQOoR4JMNtC+r0p1RWDAI5lR8miOd+3szmwk7vaQRbgqofX+dL6mEM+5s5sIt9
GTNs+Y8jKe49Tv2BY4b8kDmTUn+v5CC/2dnNRSFAj97Lh6ZT3MGBI4MiTMxca4K1
t/o8NYBxSHRBpOOjMSvKfHh+P8KpAB2A5Dk/2tTkdh9Yn9nQSkjqY7hm0nE6gH8F
2Aua6koJk3WhEfYPRNOociIsXNTiOBggWuqjPVou+ifjNWOwB4MyMksA6zsgudEs
+hPzJGXL6ZkWGcCjWcmbdNVyN184/lOUvcJmqNlTevWsTAMKjiVESsAWrO9D0ZVQ
Jx8eCdwWF9CmfacQwwxH/AXcVvCizy76Q5nYgHH13NPFehVrieo3X9yQnmWh6o9x
OBr4baOsJdSA0AzAC0evj+U7Hh3zt2QiMxDdr9OlLYFC0bXSVc6WNfTqBhUhCumi
U5KPB43MHCugEzmpEyTZS/2CwXtKn+YXZJH+yeYWLbRK4i93Z4ZGgtHazu4ryovR
ofGvKkdCq6Uf78L3FMYjKCqQzjR7Vn8Fi/GQGueJzLdMCAU3MYk1Ay+95abotB2k
eFyVyHo2k4uOGxrf1OOcnEg5x+ULJFJM3lgWP5yu3qBTT0D8HLQ1QYDggDZVbtR9
QDvWWWil7Lm+Zl/N3Yt3BokJS0RblO6Dq31Q15AhNBvEXeuL6u0UJ3ZwznRk7r1M
UOwbBob4dMAKG5qdsG7zdGEbD55L4TAkbEqMidA9gGzQSgYlxC6SvRjfLx0YFed7
F3u0+ICRrYrAKvFOlRav7aey+qdoQTqv8lD9s0kMcfrvFIKZXdN7xPNm9kIp1LWv
T9b7Ousu1jCBwqCHLEN1W71YOzxp2X5cg6P+oVAxnmgbe0kst24/UWNTy2t6liP4
71jm2tm7a8aJ9VQNwqgZaGvKp7rhUrxdBn3DFEikB4e8Ftb78K9gotV6f1F7ZNt7
BUzR0y90oj3snRGz1ABdyNGfOXrspFDIWVdB/bf5BLzSJFNdznRS3j/huKzfcoH8
spTiIk7s3erkk8XzBoQjZ0CeGznRolF2aKGQY+rsdFiTaMJcRHAJrcNsfjtyRL4R
rorUPqlLQYkcKmpIj02rKZKiKu3KhFgpTT+hV7PUSHyEasuW7IRND4eIj66F3bT+
1FRblAePkVx/vERoSBARD7Xr7Gh64gm2bcZIdYXj6Q4rW5qolCbJMtaUDCBC4sUo
4mIRk0cEeUc3pwgGQsAE9OEAVMRfDY4duTX3Goxv2GVgaonxpLWcJmfjZvsCSBYZ
DemxYWi/WyQRgmXn1hIV3Jrmu6wTfclSdHBQent4gXkFY/nS5/3LwwknP0nRY3Cj
tZ7ynX7fZinddZ4uiOqXvibNHW0xVpjjiGlS3AOQD0MlcSf/MqmziYDdAu+4V1qC
26+5bP+CINrz9EUzLg2ZAzytkAozPYvn19KzXIqX7Ar1Phm2Kn0KlKfxryjCDEbp
WVnjKRDZ2pZyJqcnNxUAh+jT6sSX0rQf5fVcJQWBCR52tzaFoBGnLAZuRCAdwdh3
h1IPiUr0wd5/nUB017B2b/uAAqjCCCupd5tsUK/d2flUJyqe3cxhlW8tLM5VWpj4
irDoYetjFgLbOIbR0r+Nw7NjoKhPFgi0vBb9gYKDSw8w0m1Bt3wpMEXkGzJXlKgh
Pg6MflbGEwzPuRnDky5s8IgEzoldcvHQgN95gkyu6pQ+OQciB6N2QGcgoz55sUcM
EmwTmVZ8pEWQEHN4pYxQ7t6ewjjyu3CNu8x9lYNve055uZDUzwSGL5dAYDX/NqSq
u1b3vi3VAdjQkFRvXhgvCoJSfgmEeIyNXq1nOjqT0JpbvNetaMW+hLaRgspO1MGC
WV33to3+DAyoIpUeBTea8bA4V1iwhr0dd/JazBs/6tjK/UiaJ5sKKTB0/2h58EP+
aAtkxcdP1h0qvmoBgEOhfqjici3bVedqb06yvLieeVw0W+1s0ITzYSKuOzTd0drP
uTlJtBluBGfvM1ZDFAMb5iTtllPWmC6fpd/Iwy7RW6miFuRDdhDjK1Vz+vx8Ui38
M6Rwu4BYBmU0zlxADEKAJSVV2Bw9vxslrSQWaQF1S35+qvnX0A1M4Ifs32v3LtML
oi5V9ne2hN0uVwPDBq4Esvc/eds5Gsvl9q5IjyGLK//MTK9Uq2fCxKxvjiSbnRFd
iu6rB31VJ9TTbaMljIezLkdZRby3xSOxsAgalWZ53pKGXe3Hc5JuFZ3zQuoX1VXq
xSPmWEtovNco2jkzTbzSisC4N8uvFZc17/5ZTQ0mR3WrdjbegfVC4qMc3SQBPiHi
ZvVs948p/gJ0vfeHA7reQ+w/ukncceCo3wqpJKHXXJkf5RuFYTwrDkzN0ojF1BDn
blsDqbMuscZm1R6JOlCmAW82IcwF42Y95XGjLxBSp6dSEiwZ1aEae5DzFj8n2jmA
xTpEKcVlw1DI22yO4YbHm58obPr83iDWsNNEc1xfBij3L+EaynftWDqodPnX+Lx6
dMvSddz4tGDBbdV33Gu3KirqnbSvDaoOQ2vO9+vn1UjwGFl2lA6fDr2RwW2vVVAn
fXAVR4FbWCmfc/pwyPCP2yHVAZIVycq6Orf4aEKEzvaewgB1wNFLlZdUdd14Ez/E
DR3jfw+dLOUNYlc5+tGI+C/T/qf7haodUd7er/InUikAPa07IvDW1v6sYotgNctj
JV6lW7fHeoFT56JP8ks12xfw+0ACQ4CcQl5utzqde0tEWHXdmEj8ZA8NbXws0G4/
SUgKQwsUWepQd/wreZWbsjXNFh+wZ9hDTZlGE7chPtoK/r5TTNt/JRy/ZvCSi6Gg
4dqRjpkhpqW9xbJy0VYy9BWtqNDGsCAbh5IpRXcxiG3vOqp969inX4b1YwriosMs
2rcoLTgPsnz0U7uSW0MVaLmHfrZTiHaVcsDQV1EeEw6/jZ+wDakZWKcw9j/RUtor
z+HF+PmyxxavmeH/xR+SKz0vwlhTTEMPRrRzIAWDOngl85byo5S6vM+CJLGBH6Id
Uuh0kZO4LS9PjqRRyMPvRx1EQwi9n8cf1jmIZZ+ZthjpCFmLR7rg0mb5NTZnMRLW
sVbOPyVQ/xL79iWkmaolVXiQ9djrrBOfFSvWyZAse1eT9FMGMPmaLjWHB0GNNxPJ
OwnUSb/YVtz0DC2/v1vVsmr34UhFWKnEk5sAZm8dGar0WBhQCOAAJUyvH6w/x1WR
jW8tQcOL8fc/o8ywtcicqFvb+7o30ZvUe5k1CwWqWoO8+WtOu/Zz8JurgvjatCGE
bqqWXOj+XbbizZ0bwafKRPt9ciSNvRLgqXzCkaPzXBi+89NsHshK0k81HrdrYN+Y
w1OF6LiPKXNyB6v8gCLy1kZeWjar/udg0ywt4D8SAIhW9WJB2/NXZ5tC5Svpmxu2
PAyiuLxpDjL+c/3xPS2S3ArYctry8IASJwR6iE0yWLJ8ZAkTT/BaXLDN8Tx66E2p
DJptNK1KBpkihkRNdW8BLQfWQpTGK8tvOEhgxHLVkHdiUsY0Z6Hu0TQkNOvXSHnz
jkJZghPgVoYUMKUioag7aeYxh78EWwLuponAmyMKRjohw8Qwkwc6PrsXMb3FN4GY
iodKKU/5qSMj0fOSrVQuSpiWDs21w9xhGSPvXt3XmmzeN4fvjgcQLh9lj76Uu+Yc
Es+JQ9dLSbFa0r+okNee+LXEdZvwkhcI3VN4+S9EwdT/f771yuq38kJjSNl7qcgL
Lf89CL2+eBewOgyRYQV6HI2Y3gKCxVxNxwaFFJ6v1hZgoDla9tbzVez6Z9NlrDxv
/wDsLCRpdpo/lHEq5wud1LgNrF3QOI3X2KVt9L49deoOecZ3SlcJNIeCHMmONdrP
qpHZ1oRj4xQnzydpJeGD2uHeJ3w5P2hbJoVgt6oGSudcbWOJdQ+wmZRdQrzmqrtZ
JLPOx+QYr9a5seJl1tOSCdf5/dT2L9Ov/64kj9RbrsokLu5E+41Duti0U9MiZ7HC
xlH0t9RXVgAGfhfn7kiWJbdrM6is2Qs++eS0ZtE4IEUgc4OhPzXABrxkvdXcIQen
F1nhhc0IL0igmFh2UZaIbS2TQ6usuJHoZcJriabLUa99EIPI/OMqo763o+g7okt0
thtNiAmS8GHO92hsKYvaNoamqo21OwfVHWeA1Bhsi/UPef0GbKIebTCDcnOxj5YR
f0zE7FD1OBdhOWYBRZFMF/VG+DC1hVXyPc3H7wFiX6D8iQhyE6V4nPwg5P7IcTan
9wJ2UfCYUtKhwK9ikG+2u8Cm+O+ETeSGjKBfwspGZ69pwn6/7UXEQ6Sx+jCQjKXj
IO3bEZEPxRneW1vRFlRDPtUGxbutjtc5hwPGUXm4WdoittEGEEUKeMWQy4Io2wBk
YrBrV8BGQ1mgjN8mwn0mmeX/Nr2XF7UMrVcRkTpmAZgrCKtgKsqpKQAedu1GpXz+
wEvDVGCvdAdjXBqNC+TEmmloYr9vQCxaYH9CqwcwV9kRFDtJ1uQdRDOhs0wfb2A4
d6Mxyx08nQVzy74n1jNsDBLmyGEkXaKmviGyvhjCs5FiPW0TnXAdZk0ClF++ITry
Vxx5rxMmIk0wVvPLiUBbkpk3qPlK6pubobe2jI7REofBXHKiGJD8L52U8w6MRCzK
QwEF7JAd3DeFQgsSK2zAIYl86LQU6aI0SXHi1vy3FyZJg8mPEGuGgy7UEnBtlotm
BuiAh/8KDd75UTDAMK3KzCxEVbzjb5Gv7xOc841II6JhmV8SmmgxpkkwkBHdZDLd
sbQFZZyv1KlFQucS09S4VYOSr7bIgmLAeiOn9vSF1N+o3TZ2YLoaSW3UEZMn3kE3
Goa/zw7047o3PShZrtmsFv7pmYDLHHdgAREZrle8VQ5HvxSHr7sjIBist3ynjlbe
n9Af6On4CjBb3wxGC9LFrU4G3it0RZGPZuB8HIZLoxBvnMPdvPuxy5Wpp67jE/98
0Y05gsOZLoXTbuw7aS1APNOBl02J56Tzaz5XNq52sADvtYM4wfdKacI9KWoEPDTn
++ZZLe5k+0KiKs/lLHirM9XVKBhYHhhv3BB6uxJ6ET1WAqb3UNdShFIRn6h9Bpox
Dyboh/6RitzN5TOCABH5+Iq0yQFShmENna1FZ4Hph+KmiQVS+5jTqnizh5jQ0xX3
+t5BYb47Nac37HIKf6yPfgZhoBvEeBiFs1HlJNwUKFxA0k/bBr57pAzSgMouBcLc
gnba7k2aSuQVHIpk1ET1IVNnfyVykrkFXW0PNB2+k5Vos/eSDwnMrXe/Ikbv//D+
0EA1gon0ovcHIPszPCl5T0rBG/7aBS3YNo//ZEUSYxEd0gC0RHqsMibajn0yQDlJ
1T+4WFp1kdjbQLDzUAqU0mroIqpzyE/O0Qof1mfD6zu1ZcU5BTs6oFJc3/CFjcnF
7z1ws5hqPxBN5NxkGRGKPmyUZhs2lpIVBW3ocL5pGLpOCKAInSv0tv9aGvmHPq0F
0s9/ZOtqmEUQxyrdM3EN6MdY6VeZZI25FwThvSsxPlvCxGJ9kNYWWEPvIWVkcIe0
dvEm30woAe+htGMGD/DYYd7t57Pmkn7i2Pm2042Bs/QUbjznHhqSinfNo/vzyvMT
gqFguedFYJ9xypsAuAIGV8iwil101KKoXL4qRvpanSqjcNuNeQ0vqeFv9EkLNQrQ
qdatJgRYHS9MBRTvV5Dhsi5j1AqkcxiJW3jMHSPN+LH4c1XR1iSd7HMkQcwBaopC
G6oMLnH6dj4LCPihmqTwrjR6PqbzuzPgx2RQHVqpsHCbTVvkIaFZFrTUhuewyN6K
8K6fFyxH7/wPS+BadwO/merU1HpCnNnPEwpVC0rBhTOrtn1BT/lbki20uG2Kg+bD
5d74XEk4g6jSMGruR0ZPlMXZPPAYxJeiHJNIzFOR6ilbZfpEypk14IOg3dSlJFbx
Iyb+ASx5hvEg/0Hm7gOlkuy2eFV9DS84CZgZA0fCHdTjifFV5bHjlORQcmNs4lEw
iFmdi25PByos+6rFRNjhyo/Ny+TXaiPWduY4KTdHHibX17K21zvY2F0PIsulBJ/z
95qiOUc6gDY28YPwKM2dQt8zWMoZFVOYMFGubExyfcz3ojMmJU3HwQTkSh8leW/X
xgPoVzCbPn8muCIz0oy7Q5wpE3QusoL4p1VWkFpAlO2YPuxEdaO7YWnJBr8AUIQ7
CWFya3AmGuMPVmLZ0FE5CNtGNh9Kz6SSWNIJ9+QfLjlg3JzFPzU7YA99to5VSf0x
PW8vZ4A6u1EDeRjVxLo02FjdVusxTg1Aj4ZpbGsfQTr5BTnPUX+pzhtDLXgnBOMs
PW3fQWOfQgdvpc/kHZFaLf2oOUSyhh8IY8HupQhNPH/FBbzwQFR38TKDpG5+YfI4
BG5TQyIRIGFImb+mnGkqikYqcqZxvEB8CCPTaSRQyGvjTJmk6OLsy1N0or+urP4V
vUb8uJVcdrhYRcOsRDnGBHfi+LpsJMi6uL6KapU6DcfRC5nIDLzQ7c/X8HnUHE0q
Ar+y8ks6MmCwWLv+J6W/mfw/2ogDnG0PlsszQ9hIYuJ88DUVKGUmxu5a1aDbl+Oa
yM1i3iEMslCCQongAj7bCMYIVRN6x9dVmtWl01TAPiujOO2KBuyEI4C3L50Sma2j
pLwq2qc7cFJ1zWKxgHdD7AWESY3th7HAhFK3gnTmt0PbQqUVfxtVX4ICQASKd3gj
BQRlBkqyd01p4UPwZGnE3HLIIrdThVHKT+Ga3a0OHoQbbHhynbRq9gRxWN0X8oBn
3nBKDHu3I+GwnTlz4+d46nNSl/NT63jmgijd0MDoghCjFec4qokfffVsg+mJQmyF
HgeQRVyoD9pg/1hfd3hjQ/OfjflDZooMPWRR5Zd/n9p38tScxYxGTh3jWbFjeVOo
HKagTsgxuw3tpUEn99hdH7oB9BcGWBdx9wtqajis1JNrZ+bQ7An6myDD3Y3tlKuw
Ykkeeq8LERzekxhnMLZoe5/6IbWglKnENJSRBJHDDu6gQZ8FFoDXfY2QIJbh6Mwj
xJzNIFHpuCS0wH6kMCDpZg==
`protect END_PROTECTED
