`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BTeSyq+WZmS/0n7rh7IVgt42ak1JyN6yFctVHEqwzayguVgszLejZDCBtMGiGbDM
g0m2uT6w/AJrOoxgUmVgoV0BqRihxFzQLSGBtzpdORVOOshpSCuzwg5pL87QN6dj
Z4oQtciphNAgj3B/KrJDjwBVEzglF4SjHiqP87oes80mxz4aTL20562E0Lpl4yuV
noMayt1XbBDaK3dFdeOtoahdWRMxkOVnU4Hu+IzVHDJ+WoadEJ/foRE9kOota/+/
VLzdAQqR3H+E2Ai7ZADiOo0uqqsFjOdoFGd2BXm07A2siK5MZzb4rxDNb7IRId/K
/uhp6IuybRFKbCuKnF3WLw7mEIcmEl5NnWfTebUL4wvkhouCE9xLESxSmdtMCjoZ
H0WybkyiylkJZ47yg2MiwAUj/Ke1P36mnVqrScPYAOhrMC9H6fOa7Wca2zmAHZ/N
`protect END_PROTECTED
