`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
teYt2eIlt2xelB9HFy7NUedXQRLsW8Di8/wGB5+ugN3HH1QIVAeRXEnFS+rfZlZ9
Zwof6ZDJT5R88B7pQZVOWrZR6+LsA4elXCZ2JOCS3H7zMbrz1zRDpKLxOuAV2Drg
/XUFpp9SMjt/lwiRpeqwamehu/hnM8HBlacQ8gMmiJt9Peac7ESLJDv+ISkQoXUW
Gc+kuGJAVazz0HUtz7AIWqIFmHudfC6FzFyqQDhpfZ4HCxLGKtohBO7a4gUG+Ypl
YVeEcT6fhdwoExUBYpGTAvG4YRTEKmWnwVZqDwrxV8W9wfL7Tct1Z5IrPBtk6ztm
YB5PfB3N6F9lmpedlnixSGnJHnHd0WpIIRfuicFbcnvfimVPDgtGXk4RaOPfGLko
t3vCnvDYuU0Sl561vCzIXggCqLdiJSOezgvkqGjrhhE=
`protect END_PROTECTED
