`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v55bO8DBiYn4qNT4rcirIu0j2e+RH/4whJv+zj/K7BicMZIK+hSsLvyHKLigA2cC
zXa20b2u3/Ta58+PlqowT6IjHQGj0GS8G4Jz9/6Jk9JH4R5K6/Ngw0FVK4GGdEzM
9yNbDohUiZYbmqO0C+Xab/6mYD0RohxT5ixawmfTDwwzmMxG3Xd+so0VJvX0E7Ke
8PXcXH8QMtid3wtYumOl+9VgEoFBlnKTncI8RXht5kxw+8MLXQQMW73P2K2Mwtrs
6znGhuOiMag6lAX7hiibKuepAxeRJ7eyRN9S6hvV8bR5TFJcOlE0Lq+WqpBAeiMo
xuvWsJ5vYizi1Wnc2nZ93TKYWuuYWYuGR3+Q94HhMK03x4uW1GHQZW+vmNweLsIM
5nSM8mIjATQ/pJclqn2YWC868Bl4i/MhV9a104JlRFyp6lT2RZhKyuXGHaZLt+hN
5CWf6/VnrpM35pnKnfQwekGVdrfmf/V5FShX2FO+inQ=
`protect END_PROTECTED
