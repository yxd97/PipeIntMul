`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjOmhdFIMsV9r4WX5+V+ENAZgt6lWUJOzGuWrxVzIoOzEtBg+lVOhuo5C5KQHV9R
T4+/+CaQoqNa4uD7774TJeygTWN/t6C6oa4WGPZQhnaVLEmy3qUsKtzF3Q6/FRag
Gn8KISKWa3sStXjk0bxSRgUoZW6tCuiK0zuX69+GrdxH/BM5AJ0CPoh2GkJZaP7D
f15kPEWS2AmSbpRVoIfqvGALfz0o7fpGcyH1joFHF0kZUS9AyrIw1iJykjnaXkhF
OxU7bhc81Ghjw7gggcT11tcqx1a5tWxXqjRvBG9ZH9lh8b9x1I1GYK3VDVGLDBUe
AgZQfCcMrM9Sk2f/YFXKTdyXlw9EKC7t4Fm0X8ai5XW1tx6ekAMk5Zdes95ndmFp
AuNqbrFn+uhB4/mpX0alAKY7CmFiJBIMf74vA+svdRD2XJq3DA9Y4QZhh6awESVc
JpqhkGRoRpMg8kk8EfRLohWCoqLTUiT6FK2uo131QBJZJnaJFYa/f6ANXojpCOsY
`protect END_PROTECTED
