`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6tBsPPVV6fD9D+3D3xQuBwCiM/q3RQ9BRhhox9JSils9sAZvT2khNisWWfKDRTqB
wXidz3Gs0QDJ+KWYGgL9o8DM6UlkHKTb26Mzh3WP93KYp5+C2p/NqlM+bTVjZfWF
kmyvXREti+XpzJL+vqAqX5IZcx2D9v4paIcYGWI5RUE5sF7jIv7am7vWcHNgkk4u
jfCbv1tZRijiyatUy8PJaOX9l88kmCc7b+SsDpl/+7k=
`protect END_PROTECTED
