`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FdzqFR73hB9vBlLbhhX6ZoeMiAK+R2dNKNva74umZVxGftPn+oQoTiWXV1vjekh/
PZ4wHI3JL+EcRIg4Z10VqcQioS9a5ATXTlOUS03VAVAuWV/VmksYvO3e9ozolnBE
Q3HGwEDeylq7y80OdjcpEUVNma+OV7r3cMavx4OUEZHcEdpA87z93irFQKxpK6yj
yXTtkNUrek2IWxnHJVd6S9YNzxMKOx3DQSAtInhDZhEPkwjZS6FMHXy5mjpQz2gb
jsr5ifZT7LIcvJKfY6BSpAUgTKIQSedx0F8jLOSPjIcMkrcYQ5IPOMNphiLxqfMl
MUMELB8EhnxYVnLk3pwPha1eBs+4gzA5OjHejhJkx0/Pn7rahMLUPxvvBqMelO2c
PWP6+jWOTxvWBhmr7F5fAL/gKfw7MW3H/n10T/Zt/9hKo+ycJqKHhKYIjsyi4T1P
edlRyx02t0tTco7Dq7Gdg6HfMR5YEYtycvXnogC4qK5A9vgjcK9VkUFHHdPgsqLA
`protect END_PROTECTED
