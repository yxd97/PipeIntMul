`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3atT/lZK8epOTMvhyu78gvF6WBKkdV8j2RGvF2jgaOYlZQ4hQ+RPuJIGVvoqh6Ws
XqwfPrtvxc3vJEB9M+vT6SDznx18QQKsghTEaeoX/QWevds50eWvC2MGntcqoABp
RelgaW1vxJ/RLH5RD5AmnTpwI55MK1P1Il6FQRkYKCZDyOe+N1Py2KMu11zcFnFN
5Xw0EkUlUuZjLFETKZzx618Xy5mhtm0Ev45z0tm4UDCnnmwuSG5axV3AadMVVZHp
tYavf+cgoCc6e3/Zt+FqdZk8N8WjskOayM0h+lku2wyJfLJJPXwwK8VBBXW6BCvk
/j3Z/ioTLfhinAC0mQngjdkSCrT3q94T5UlPUHzx7wOYNLGGH39/zi/dFRA3RpcF
JUJBSXZP5WfE0V6HSKBq7nr0eTUceYvsLnZBcdue7BKgVPDMPoDaSMNJ4DsNtBH8
Gceh3278aYIVRSJlaR74iSLHDZtMziPR8wsblRv/fw95but2jNTolhTR9EGpZEft
7f8AMoPfYkkP8BpMg7Tbg0nAxPxMHkFQuRCzW9/jAczu0c00MUpk/yzRCDzQDvjD
mLMFDbef5mkRDGVtb/YLpIxsHZkqEtzoCj9yr4NSMQfl9pSkU8BAspA3Oh0jdnBq
D7EmCl3ynvSH/SZvkk1aKfxI79mXglZHvDpGJRv5gGOIwlPhUzMvaUiWoV+rJm2N
zJ4E+Jo7zeCUYWFiKkfoeVJLmKLrkBepRimMPvkyB2QPq1veNOwz4yLEXS9LzTro
8aLAj3TTRmo4IZqu7Z06bbxlkW5T1/3+aI7boSSsWTBZPw0FCoxQAIcdVlwETU8u
e2A/fWUYwz64ijcX4krv81tzt/045eIsHnR3etEiYw8qMpMwmPJsIkwMHNGdcNnZ
lrYwQRwe3aJzBZh0PThIX50XD9nH/H/8+mJcP++Oo7T9fMD7rwlTehiwc6q92xLX
HSMjk16H1tcv1Xisj9o7OPl4Rdp79CAJ871aRzaYmBVXghJ/5MkrOlhc8OeQiszQ
JD9+dA0DuJxCAeKu0xia7WASnxxKY3Divv606+Ne8AUEu0ElpPbqCjPiSMouwGdb
nEkn9dGRyFvpBZQe9sBYMsvR3XCE8wN8lG1Ferfo/tGpVRcXGiDSOvXxteXPqcZn
qQ+Ffsr5RrJ3Uvl40qVOZ7ZC1IXsPMCG/TRGjndHhZZDmnSVHN5Fp+t5rrv6G17C
8vY474V/iMJb8GR/orFSiRFvVsN+G8Kp1vGiNC8T33b3w8GQFV1Y2+zZH0aRqLrH
wy8QGho84iX+19crTlXIxs9t8dkUZntmogwjdQBOBAo+iE0EhU5HSBOMC/i4AXjd
eFL2JKaHQiXC2nEmvX2Fh9Wou1Nkt2UCEOnn10qbVjlTFuWSEaWfEV+BS583b7RN
akUdMAuR1G/5SMuTthldzShuPSPsqdxae7WnWUp/pnakTZ9zTYrAVCeFCqm+dcXe
VZNCA5cpIY8F/h1nSBqrAw8fzEq+aWxy0STsL7Y3ZX4SphNpyN1ma2dbJuNgCymS
32oXbUiwoV7yVo8M6oP2CvwJxUXIJONFKi2gSu1xqg5fcoiep4y5p3thdcQmSG+4
t6mCKZLS6RMTjEIreJi0c9e+RmFyJrsPIVkhdvMkyzxdek+0BVHGxFD18ZvOjrmn
S/2XhR8UJMS/i+u4YkiXbkxrsHXXdUHoKEMMMu3S1bPYvyPZO7PCQLl0cCBn/TuH
7odwP0Fl6R7DmcnyaG7feOVXAJFAcF/VO2CSFx3zXc33JtLvd+MmRKYg2TINz6S7
cM+hEG4wC5HjPh26CuE8iWyoAJw33K9FG6lt6QouQOatwBCy2iZS7qiboe8Dc0lq
BBLcSIGT8EP8Yqr1iK/lEntYweKpPXHMZMipUrFn0lPMtnNpLFSKh2dqjSN4ZnW3
nDVZiPWE7wUzBgZNJ7tbYEO6wM73YIpwmhfoc9QiK50+4I9QYSfhrjNjiSLbniqV
ivzjvwP1zAKbaxIXdP0SW4wlMjbOR2o0B1R7Q1QUB7ykQ0kltOKMtQIWmO+xDFEx
bZ2TnqFRMZ0u23+/Ziefx0ocivgV9G5iJYYzRs+qg8RaXhNM9Ya/PPI4qcz2Ay8j
NlWCETpHjCWcY/AzyuPH9QDp9w9eVTxbMH3NvjbonlXZwa5zxBKsFOpxDdy7uS8t
DdttQSnVeNvtKtvmiu4Vue1Kv5lUhhIB8xlFldIcWkhxHHCQQcnQaYSKEwgLUT4/
b0T9SQrbLIonb49Dvj/xjQHvCm7xiGIHTLe/LMAzodLMqUHMXQkOCqVlFxBSCSrf
LTLHZ+xGx+FtQRa0yX5a7NvNJ7JfZ3L844EBGvNk4M0TkGkHPEDqrUENZgR+zk1v
/Wy3y9RR7m7mjyMw2kcPHibbvdRIq/Y//6363ceM/HSedM0uP3clX4jzBamHmBBG
amMhdctlIiRDxHTo9IMTJnER9SvvL63HSiH8hVhBgmRxTMuuKiZG8InicMQTItVN
3yr83cLb6X43CzWmfBEVogBh9QNQR+lLSSAfHezfFb6EPBtExpKZ47yjQ8UzsUdl
nGO/tqF99aeYSsoAXIYWaQFG4ZtClstDIfWzSxQtN6pF60+h5CUHufkwoMg6r5GT
Cm5nPXBsIu87PNNiT7K3XjmxFa50/mFZ4Q8VrlBEisUStHPyyEtwtBbu5BnYQ+c+
Vp8sYPB1o5RAu8EoeMd/dUXkdZGkl+mKte5XHRckMQOOU2xKVnDH4lCi5tVB+Lsk
CE+Y6+RgbFBMWcY5UR9dBWvlaozwileSzubDEoJGDcTZ6UCGr2DhWNY33p/a4mGs
DIOjniBjJ3mN6iQ7cMDX/C5N5spt5fiOaKGA8OsD5aFgOqZ0AaHZ0llCASx4rg+F
BNJ3wdVCTGdHrx9SBs/Obm2m5iDEEpYU7/V8YosIWdIjTgcL1Jo5XOqXjHbPUOYg
KXbEz8rLi3toUb+MXgjjwhSyA/umQEKuhevcjIxK7oPOb1GsvsDcbf0TZjuuoY5g
O5mAFY6CAuXfdM/iWe3NEJNuK0pi2j1pcKqvuROdw83OqaXizRcJRsMEkGmr0i+d
4J6EUzOwJmR+g+nkAOji3yAHVr+297yCze6ZeEVJFPFiZHQrZIGb2t/03z4Y1uOd
il/5QhhbPY4D2wd3X35vD6k4KuuzoZKF4EgRM8eV0SntxF7f2u89cL+U8IkW7kIt
jMwIehp/wkVxUdPy5TI5SO8eqPv+Sbbgz/TVEpEe867vqT6OZNrTv5KADuBL1zn3
5KdHSmx22kOAkVJ+JOSIEyEp8O64dyBGxOrYbOdCwAxwzwixWW305abZF7YDigE4
nRhodhuq0ULcw01Yinw2IGiu1WKDKLftp7buym7INYesEOB11NdElZke3zWxFaDJ
d6V7mdUWXFnNJWHRjhsSSm8cAO459TPsVVekToIjzR/sRIK+HX1HX9KcfnwP8L+w
3AKdT6dfTlIIlZaiZ69tq3X+eToHOD5797IpBbOQO+28z9JAnO7uzy8W86GN+3Nd
Eu1CD9gJ4wFEzhXRnY2jbLhIC0k9iTf8+kX9JKJPBOcrtHtjVO3/jjfA1YTutZwg
hQsF9HjdpmV6X5YELnM6MnYI6CJ0FpySo/iShdD8Atj0oCSSIkZnHSJG4+JKD5PB
tDQBl7omYrCJUafj7maH/1Y7gQP8+4pGHeV52IpePVC7D59f27n+1xcfGWzs487b
DkELf1x1ATmwx3lIty6pReZPsRBFfjhXVGEGk4m4//11uy6vcJdciRU7HAKJvs1Y
UYaivsMLKoEdRwi9N5V8ibsR1gvwuHJUAACZ4TLqX5+TYR2jM2v5nL92+IBQcUK1
k03hxxPVGYkRvr3Kb13GUMNiKrdU6Gl5PyPGrx7vEl95pTnBQnYATrtwgRkv8XpM
kn9+ARrC2LMF5Zs2OR6clLRcHR3R19dXu5XtHrCX07qsv8jyH9NsXWGm0oTQgpOh
RI4IRbC0uhlBPLyD8bwsCq+BUeL9Fq2D5F17RUPc+hMHlEwNw2VUcGvmJu6j0JcF
LAaX2LzFv0w51id6tuIZWG8ns23dMuqlOq6dZ5PMbTy0swTenj/xCs6MGliAWjYg
vHMpMhEyA5xvCDNNFhVtU7x8SJNRmcD+WPgmi9mMD6Wj7rjiU4LhWR1dlAUqBmuL
aZrscVjCGVRAVusfgKI1SjuqgWTukUuvdpgbOvVgNT7o/FJ5T4xnlSWiaCmCl0I3
WO4LQXmaevdQRRl5/vpEX43QHHgschXKJqFZa/CHvmJm8PjmcWWI5QnOo4fb5DFJ
iVoBLwUF2gYSUTN3sBbxRGxqx4Hh9CjnfvG3MVoGBeJY9pUuChiPfj/HE/kmVYcd
fkEzHvf4SlujU8/8jVemp9S3vbdPUc+HwduGu3wiDZjYdBQOmHe7ZOL2Qipb/Em9
dBNqL5V7Sh4Lifw2UJ+dbhM+m5aw9USRZ56oj20uaSW5u3Auk+CmtyEeWk4PG/9O
haoEyDynWfZOqqbpEbf4kwF7BsJcKzbPF/8zSkfJRNbLM2GS9TVfyJzMj2lBGIAi
pqHGG4JgqojtHMLJlgRFQlcIC9GfWzVsHU0S6mpMR8dWF9Ad6tZhI4nbqYsd5f6i
rKT7uuVfAKhb6+7+02lLGhd9VjsDDda8sOR+UeHRim2ke/wlTutmiJKlab7mJ2z/
zL/go4avJXCgwhQ2bEFfxcL8MRySYIPfOxaeTw9Uq6oVUts56vryJn8rm0bBrAh5
svV89vsf8nJ8f8FNbsWgNSIMYtEsTmdTBZixVoO7Wfp3Vu2ouJxLVWLCmRuW+vXK
n035Zdk3Vlzirk/iYMxJv+8WBCQxZuAWc4y0iHyRK/zPdT1NAA3oPyHE3u1WJGRu
HnzpixGLlrwgp9vA62ZvzM+KxsIuhiI5SLDH46ZcCUX0ofcFfWOmO2nVsOs3FkUY
ICwyi1bPsC/ucCFy3Co/ezvQhxJFUzRMH7M1/t/+ZBBP0R0NYUTREiuzUTCbD+6P
u5YijR+uQb2nX2/5Y05LwKoBcKVnyhQvK+y3ZoL8iJ3oiY7TuCIOfPGrsjtYHgYn
tYbTBuPJC0QGCsVmdLMZCimkL8oMQj4P7xxCqoWj8IXVwwVgPZO8JF1tTpvzwQiT
AtYo5cOfVO/POqigR3OaLVfM6PtSlSebDKy9Or+AYRNOBtGmy5aCrZZamTN1UGh6
YDr/j59ixjpVrYg6isK8G6dUBMJVdWisM5jxQHHoBio0j8a0I76BOMRue9AsKn7I
ClrNkAKllwkHfmJGxAPvTqI9Ae1pUdGWf7JNaryju2Usv4TjCbTziUwr2TKCTHLz
lvuoObnmi1GeF7nkMmWTvgSGjbZ7bf/kwFZyuZrAZ3r2izOjiZ/wSC6ZSpx4Yfdj
1HFPLjo3wmmlFlFGd8cp9A1b31sUPgQYOygk+nTOkq+XpYJb6I0m8WSjjGuGiP3G
Engh1ekmPOxXpE0TfAdnvE5V/weu2XKsmkK20lE4WdcOr/BAMy2OtMtstz7U66Yt
r7F8wRFIFz4uyLPel3zuXAIDXic+a4HX9gHhNEbhZpKdgcXRNa3SmfulHfJeAfn7
KSSm+ZQxEZiMm0xEK2hnzxx8zT7d2t3gDXne8yTpcoWv1bUaJgkzqicVr5/NOH2O
D/ClshwLJlWywcVpYDBuHE7rJK8wJicHRB1XPznQjTdNEJ5e4wzVnfTDyxgtd1cD
pzvX+vpyX5ArLzCBkFpveb6w+gckefLf1HOKP7i53A/ed20N6KOBfiezNPJHEya+
4c3NZTnyYEbgVOBfPj+gW7trb/wLqDU5GSrfirKV770+muX6FaEcUPtRMWu1EM4g
xon1zY/JdcnijlRSPfPg/gXRTn3ub9SXa5omYUR3W8wKgrSF1HiF2ljYPtxDE4Uq
9ciWSzkwNGUY9J3oPeDFlwxeDA95Q6uziFXwUEzZqYtyeqmYFUatew1A9RuqUyMb
w4GiM6ePF5J+sFnm1iaM1n7Hc7mkoL+CG/i0apDk+nHJfUTDXwQm+fg8mhHh7A0T
Wi66P69v2OJJaAi95aW0TjDjvsWkrKMF2VFvNwcCxOxJ4FsQmgN+cwaMcIaeMHQN
RTezmHJcxVgSXzjUK3++6J7/67f9+WWchbaQgIJV3q07bU5OSWJUalaSVYmVFalA
H3NoeefEUobP6x8ajb+BXS3qsmOC1LnPUcI++F8DFxKMg8ToMhQv2TMvCb5Jq4Bi
trAkf4uSbsxy2e0Hkq6CVLkFGS0un9sFblSnHPTOx95iwWMSgLADw61nlZLgppfL
hHBUGa9TGlx7ixgXyL0eXpIKAAjZLbt/xQy4DR2pRRoBtwgflgHuiFkwxU41Ta2R
u6LP4RWbNo8YGFOMABi7U50R2UIub5qZi8b6zLBTWFVUNPV7hPvnwwQW+mhopYcE
K5nZh2SzR9Px2GTsENu5Bn03yqbuY1KAUY4cnuc4yxzGvZBcALsUt5tZr9a27avc
RhRwcmA1c3WBf3JhO+xkLztPhG5rN5+6gpS4UiRifgC6CMWcQlsBwVZw3iBGIgvU
WgwzjgCvn6K5lRAzQ8f57lFXNnuwCV9ALBX2iZOrvpUyEdzAeK5Y+k19OQOsxL4G
6Wcx262JKtbLhGszbfTdwqb+ef5T+R9FI01JpQEejG+VUP360gy+/CRf3eRVTBF6
u/847f2PjFtlb/n//g4C6tJeVFIB1EqFq7Kwrptfiig4Ag+cx/S7jpLQjN6AqwH6
+2vUhgIQcB1oUPiUBNOBkUQWGbsdUM91Z94GJCUg58Ezxtzw8ziBAHOTkmxPCYnf
xaBsIwAYVxtYovyA7g1/uPVa0yo4PE1z8JtkTzoKAKUhyVhb5qSI55LsSzbVgD45
e5lOAnj1NFGUzoWUqUz2r7/N9SKdPJjyipZOWQuJxTkhWM9XBHr0fNO4yBkemURs
sKHBdq28xinPmEiSS00rygMaaK0D9oljcMXckhtUJi0rysqEXvipeJvekdxcuf4O
XeUnoKn2JSBjEB4l+qhi3jf/F6uDD7yFEofW8M+cd8quICVEcBwCuNNq89QUPx68
KS1C3cGiRQYSO/nitPhO5qD7Ky429Yn1NlJQLBFggeK07MQjXp8FiJmmgVwI5/mw
gkNaiOvLSm0DtFcYjH7ipqiXXj0/nVv9WnCLIIfTqrxyei0ffBY1BFWkLeIZFgN7
XjoWBSOQkBufPhW8r7SWEZ54EyCn6ykxgiFywdp+3iOJpnCKQHp2Q2PkyGrKA3sz
0LwfMDcO8V2ykFsSqDiHqKUMacFb3fTTWt6RL8CIvUPhpdLOkAFhgqq+DKfp4mTc
MiZ/CqDFoacJvz98dhWldQxjPnSZkr7UwkE9TC9//8B5iNHa/CIYF5FKhhkGDGrv
WZTEqMpcqCQKzMdc60FBm7KTEznYvfViZ9oZ6UEwDfAe0ZI96EdUOQ3gEmUe8uzx
lSNC3bSSzC96WfxFr4ygWipXlWRFxVo9R6ZW8ABpE+XHGFVsM9GdRzrEz1ObUMAE
/PBF/9n7AME1RAaSI8OFTDtm6IXaJHDVQ2KtlDzE4Dwn2L5lLlnm5QyKmENeKMz1
pKFnEGJ/XYQOimiZLEvcc5C2eaUqMBve2Qa4p4yedtdfpQT7DSv+L6qPnUKIfIEb
djiWpuNAAY3dYtiFK37AHcVYeMd5HHp3qA8qokjal259mgX1ezyV0jvFGtJDo/iF
nahwWDwR2IgyNkh+WWpFVE6/4d60OVE3q8KAZAHigLU0IuM8rU5+fgQCmVgYvyFa
gsFHQKBdQtvmMzJREMWOolcV/4MMMcml1x6EBBXw/LL6tvLSqTn/4i8i91iU7MY5
FW6vwlvAkiZZO1iOLV1Bu7j/PvdK+qbdqBepZl4BUYpdtr3k533roV/HcZqI5ovV
b06RoWUVGeFwUfz3QORvcXg3DfXOuXQw32tcyIPDx4qzH0u9hhFpr4qWxs/wCgYN
HUdGg9tmdlL5jzhSU+bC+vkIDNKUjaHKENtpo0R7BO43TOFFZ0yo4C9t7czu6hjw
thuy8WF0WLrUv+3cHo3aHkHi3YoUJdM3eLCGBcVYM9ax/EinAJGuwjvQs5rdx9zz
6n7g44QK8HDpL1nEEjspt7yRxxqwMnxwYIGwwgU9jCknsr1Guqd9uVrH4xAwYyKP
6NcdA29gGJS1Pnp6t9+KjRpoRB3qSs75k59SsN0GAhrzEDC/IZt8oKvthlTtSvNI
2R+OnDO8bnWLLyN/yU8t2aL67agBVK73P+XkNp+Gsi0N2bytltai4+0+RfEAh1e7
q41AywbZhlkQiBZys+D/NzZOJAMcaxEwIYLhE31K0Ja1S41BSF70Be4U0rBBUOED
oufYVqkTL1waEZlJgWSpLMn3GJ+/ssZwWwpexks76DPWDd2KxQiQ7QFQ4P1PxTdL
0B8VpSKFiUDl1eyIMOXGmdWXOofLO6GFJEgTHxAXCdSHtyhBFiRJpdI6UfwN2A8n
JtOKevZHMN4xoKmZJ/fa88TFwfcpywsWjp/tUzJ5x0vVasRUxXoZCik8NTGQeRsI
C2sMg+WnBhXDHGKxujhzTCO/zHc+rSjDqwV1h6+HhwOHXjODZ1m1BM+BUmNv2P5V
U6X0080641MxCQ9mYI+QFJm7S3nwFrhoBEoHKyYunoUjMx4ZXguLKUdGrzD2u1QM
LHSzn8xnrGI8CH5Y6Ps9XraY6sycT4+SBDUSZLIdTWnNjAZhyEHBgErF7C4cdpP5
ksa4I8QlJyxLAIfU+0Uawglf9RbHzgd+yNfjiK5/ohP+/XpU2L+jQXpJzlhdfCV9
XB3WfaJ//QXD6vHcjIfzQcQkCnYGnMCUSX5GLnxpdg8MM5fTkvdAa6gImbzW95fn
4IOIwRFH5phfG2kTttNcwk1tuVBC3vz+ZCcEapJKbByaPWqHhDoCf+fU1n7gH8G5
w11xRuwh42pNZtQJiZwRUB2mGFMevils8PmvOoU69iffx/fSSqcn9BmoTZaEm7+Z
7lz0g1vkj8OPb0hTq6D+UDj77jAzmm+NvesFL3urgYOpPRF1VDWhBIK3GiiHEj1r
5VY4PistmXNPxuiCetizZGPcm6Gk2+W8k7DlphAl6zH9w6VwywbKqMd04QPhIVwy
0+XtU/D69Z3NtzSnJbd/vEFIHPParwLcEwnFhSN8huYRGeu6m12OU/5g7YHaT/db
trwd4CCdHR9uoMqMKoG2M1l794py9HgFdzox1fy5+srF+CiXGMNlKuZmrxeBIFyj
2QnzKCFGb9tn6AQx/JRlHZjR+rGDSDbN7g0V8GIYX2/5kmvlyiNa78+hE9+QL5ft
oVOF2mbs+6E5ROd6YDXAz31p+Fkq54u1alIWAaaRqFio9+m/pQ1i0Hdv3Ejcd2WH
LiQW1PAUFpfjbkxMx9DEUavCdkxKcFVCzmhluZIbj1GfUGyBhJbV7vVdYYVeT/jm
GABP+VGvjh+zuLYp00ZHWDdzyHNwoK5rS47vwhdLNa+MRqv4ghSARlvl/pKfe/0k
m9OvCdbx5AGx+A3QiEG9zl9Jtj2IETeiTVXeWbN5cDT6rD1nMmSydTK5oxiq04PH
9AqQGv44M3/gngWjOiTElSJUu0rZKE4tvLnL63Nc1GFREP4nY90DmnQ4UnErJIzS
2LQjY9npmYZaz413Z8cpycmwYkMb+3qkvV2Q6HnU/1+mmxCp7eY8apJh2FpF+MFi
v4v8XNx9OhUz/9pVPU/kyd/GVa17j5cM+Z4F1pePnG2kGjodL9zqSNWR8nrdViuR
aq4JEJtcFEQCojA1FQkIC9w8LyxJ+kMImAjzbyDINvQo3w5+MQyWhtIMZy3jxX2X
XGeddpiK56wwCz9n+DnggQIVYAN2oIDcyfhWly3PI3AIw5Q8yy55Xwo8YJ5jc4C4
cobxbgLo7ygvossdsc7t861MFYLkk2akymYMTbwFmdzCpE82em0ImFgLf/AxRHU9
QRxvSurX9IgBy7kqbIB/XY4SjOsexGoK1jZMR+OAlUeAjiJ4t4GnlQND0LtjXAM7
PErNDsgmO9M2ZwnybaYjl4JuJtJ+2IVIEokbW7g50NxaWwIl+vo89gIDqPxPlsos
tP7uB8AXqKGd8RcGwBqT+NkWph7i8899c1K5H09GD06KIHNfI97zJNOMfz9mX4ax
+ri9mh0sMPGv/E9WaIn3P/OKVA3Ab+pxvdRtY6/P/sP3f6MwEAB/SvHqg6oUENkH
j5caF2AJZ4RIhwQg0Pw9vBCri+lPSrL45v8SZqj0cgMVisoF8EBiglmwGlPwdJuZ
8S4n4h66pd+VyAEUV8BkhSvqffURy2apjPClWUMmELkKLYHw2AEVxoMCv6/Pv7jJ
mAPcdOv/JKTC06THlUdEzqtMmbpqhqIaY50UB64pAdZJRTPtLv4OnJOA34iOLnMu
ryCneSOIyAcuJFBsB5MDQZgG0f1ULgEGgIVKk+AYT9vagR/mFgYRDIiuFsx0mF/2
nsCo964mCiVdmzo92inUU5BsmUjwak+T47NMcM2AS8mfo/Ei7muQbvXcJ5HJMODD
U61WGoQohvSx5JQXxqLH4rtQghNp8Ijq9md41M2f8eZFfAPUB60byFECdPm1Ttrx
mmvFl4+QYcrzCZ+ON+GD4i3/3WjDhojkGoG6Xtz0LzlGkqPt6hZCS+5ful0iefEI
p0oQVcTVU4qp0mADRpWPn4LliA5iLi/tTcv/o6HEZ9IqqO5P6VD0eS+Fbzh+V9Ha
6R2d1mW5rLGjEqzhnWTcn5Z/ZWXNXBP5jtiUXiF2PFdIlsUjl3eG7eNtTAOG4Q7T
GCQKKBx7KzcPlaJ69CRMI9bvqaPZAjyavrmewiBZyaeR5/qjKdGenVooKTpep2bS
Wnzq49VvuOAwfVMKmEbQPOpGGTyWPxO+axpTAXl2QqYoxGWqX1uCApm/X/J2APIs
xZkp54Z+6e5lNRgG9GfruhuHm5vHeaLc08kxtW9d1vl6qAHK4XxutBYi0XqrnjQ6
lkNbBOZbix9BNLGwrpCIwdc27qwEs7rxyhSdkJaXNKovapxt38VMhmiMQS2eMC9u
TEcctWNOCirfbHD+P7ix6n8Y5DBHJnm4XShE/T/kDvrCscLhBetYO258obdBpTe3
de/B9CHlOHYt3C0W90DDbLp3euaACf/1LNF3+2FptalgQCBeNEOPAnHPg8a8u3Z/
P2k1rXrnOpxPBUjusSQ+NENbnpkIzb97O6Bc2J3Vz1IkZxrnZFjxdDwSeVdaWOlu
4FUMuGnuTLLKfR6P+AwKf9PzKnItxzr5KboHFL7QEFfLIpOVfIf02ZKBr63n7Zkg
Cbwy9zAWBFj7YgSzrdfq3FOL2jL9rtUBXx+/L4aTlKECkt8EX1xpJ3jap7feiEZx
AgnjRQ6CyGGQJchLr/+WIIUQWjlfyKVEiZmLtOB5yg50CGuOxk45yLAFWri0EBfb
EnmmR5q87Ck30z3zzAfCs0OfhCLA2SRS8l3IKFEY9ETJgHvsyRu06Z/d1y11Pgdn
eOLP5w8ktc1x6d5SAU2N2tDWPOT64q45fsl2bf6i/GVLghPGR7heTrzGBPHRtv81
jwpU5vcZllKpqxbuW6x2TAkFmJZhNsd4YYMM2g6Rgevwf7+nSJpDaiMvzQVfsKJj
04Ztpbc/LtaBjDxE26aIF2jvV9kD3976gq41g8gAxxZoieRY4ToAOAsUeWjlJl7W
+WJ8+SKdSoU/M8V7kNvkKLOVgsk56EFvcEAE7vLkShGnXSQPa5hcrNamAI1TN337
i2hqzzDxfagBeoWPdEVhVhG9jIptqQevCTlKCRa14opNXraptfzIS/T30J9gYJFM
RuxU/ezLBc77X8vacWxywFYMO6+sJdtUiAuJ8Qm96dF96eIfINGdNcFdQNLZNjWV
Y7fP8O4JzLAmvx/s5LEg76RUdbfWkS8YpWMEcGAhtZIhjpB7+SR/AfUgdHX/OuAn
ipMVMoEfc6Vnw+U5HTxOh8YIwJktY1kUhZ8GZn49ULAd2Qh3UIrmurYJGLUk/P25
qSXXQLPKfpUl9fpdI6NzgE0wTW/DRcYQjEk6d64ZbtDQKOjQwLT4EitNocfS1Cga
gOiHvPKfhl8We5T8DyBKGKDuc5l+MRNwuKgEmJLfPnpnJWUhXxCUVEIQVd/IECsG
viG/B/uKvctaD0h0s7QjENiFL+y1QbPd+Y1CIMvBdqCy83P6ADkyYHpkEsYimWuc
y27iSheP75/g2P5ZKqPnyQQb6/Tf77WT0UTUH4CVJcXhZWXgwhQ1/NhQRGR0gjmy
erabf1jxh6moGJ8yzCboY25iyyHUrVSmMl7OsrPr61XLid4dAlF56SjBWLxx6hAQ
Go6pupE/ps1kiQ68OY4YO62pm6RuFSAIANtQpgKkQhLmj3gvBuJJwdbEEnJD11pg
duPVHpi/lD9ZSYZFCgBinRX45zq6lXaBQRU0aOM1NsgkwrP6DAZIhU2farkbAVK3
NB/+InWctfazLW33c83Ld/J+Lgsxj4PwxF+v4cZ0kFZlB2gfz13Luxq60s7EDjFI
RwfAy+c3kNr57c1nEVOE8Yr5Vx5QHbodU8biIT7KlmMirWclNSUWnVo/ATCStqgZ
fFkWZ3ZewQlhnhCOyRT7oGcl79AM22pHkGylb4X3Y4J8Ri2vUWiQfCsUvlq4515I
kWCT3Suwkhk8LmY3rsqDU1Oamji5VldgAG/AnliEN5Senc975IxT8Yk11iHnw5uJ
AkY1bjaautZOxMJDb5cEcFFnXUv7Y/P2y4/2y6AsNqcF87SJ/i1SYnmFJD6vuKVL
0GwreHADKWunoOLsc90eqbz7hNaVEgp2VqlVObSEl8fa0Ksni/eiqHX0iMtIyzNK
roHG5Q3JNqBGTauGurXMIslFy16pOH8De/8XVc7McihVXLxIm2O3JBwNCXkvKFYV
EYPiYop2zVOy7Xk+oTmJELzHN9ZGuJZCD04ibJ0bTI7+GLEJAowYSpopRjzu5kR3
0WalMfchRbf7QDWNNWvJob2B52Kez1Y5/Slr2XcqF/+zQzX5NIeVdhD+cFXQik7w
cEuwBkIT1yza5UBl+ZG658W7s7tQaehrx6qE6LrychDHZwZaem9Anxxdqg+M0zLk
BsPi2I1XpoTjrSbpE0rmd9GbmnpGrhpUVfcwOHJaAPpsYQv/g4XLcqXSkDbQJkRm
+7kAEc6gJPIacQbKwchPpPYD1rlP+6jYCG5oLJ1Y5BJ37TCLbj/m4u3eCA+zGTxp
uJaTP/WvsEIjAGOJfaG2HjcMmaMObwSoJ/GyHFQBHv8i+EeMMrGNQGFlZy2IyTbM
vRwXDsVooX5m5kpUD2zBvkIGcQ1xWzxFQk+ZndzDSH0M3PeBDYg/6WAP0lBrUnum
j6Y5VGt0ItB+siyiepGpOVezABds3zTlRcCkBEMCgk8PCyjWe5fPnYk1qjA4gtMm
4OL0sCiWP95veiPPiUTO3mHYmIGm4ujdWjzwlGMCGI1PuPR3M3/eLllTKJHSvLuo
TCH32VOxoG0xniG+vogU0IDxbZ2el+FFnGqEef5x88mFNmQ1UfUbIdI9MtiA1DRP
I+Zit2UejRsZoh7Lz9uHw+eVuWapYW+0QBJgiqg8T6rvA3OFlxG2SSHzLz1a4B5P
NYCetlwJSXCeXVnNKaayEYwYm23gsBE+6F4XSWZrk6F9PpGLPhj+bvD6Km9IBOOO
XqbGnijfu3Zij3Y/7zNM8nB6QfLIbRRZZ0zgR+B2YG2fvO0AM4LRrr59MqdMMqjk
9PHY8hUqPWNy8nAN9OJSx9wHYNgeC+1i5QZE5+KfUo+AEjrMYu+IpLbek55H+Kpm
Z4jty37f4dATdE8FdJG9cnLgvVnQcOiB2jGzekM8M2BCOWYhxXh3nRwcEbhWS5O6
aQAuetpkv+PiB9cR7DoACYa+fi8p53nd/JvPYlKRX8+sZILzRE0FOjvhcY7f3SVK
UoceYAt7W6R0j9juaU0DJs4/8NiPVhuKn1+acFZgPZLycvAJNXAi4a1QvIWk13sZ
DlMLct0YK1gZWaAH1c5lUkPlX7+4/zeqSTmEH7rNFjqe9GduRjSSW66w3HMCgj1C
sCR9G5MmkB/r9iuSw3S/Y0ABCQl/6xT/ACGwG5RqPCzhYmk4e3egrDZd5qi83SW2
f5ZducGQLkSZMCz3c3UpVzc+KsDNi9dAs2RWpPjqjwB7noPtbJoV1eVMwtIsUt/c
fls5h6PkkFLZ4lwr0ttDiIp8gYfgCPmLKqxm3zknq5hyYeZbdGSm55PO+WX+6okC
4IcekpCIKE9od4X9lwqwVDnqMU8kybgvLaM2xfwWIvzdJDPdy+R+25kFq9HzxoTS
QZ04s5Z+BfLpfT1pz3vTpYMbTxPz9K3Zx1JBTUM2I+qM4tN9vla28lsHN9Jrq4au
loT661fUx4ne9wVXPV/dAQKiHIVTIY2eTjfh0Vfzb+r74dj+D/ce4VN5nsEsigPa
z+HUunApja8LmVHi/vHW543dBZ89Zq4HC5WTYTKMkIhTZhEbgD3NdIEHeLwgA8b4
/SDplDF1/FUA7RUG8aC5nOOl9lRH6B61bTEWjM3fgqcnenTPp2wZSwbBiNw7Ls5k
CHxrqUxUPY3KZFAdcKjbAYeq+rgbhgq27BEbgYmiFJiZXXC7t/nmYOcrbF7ySccO
KL9wPwrxP8UrHtJ1IjzI9lRhzSeOcB6Dx4KBKFBXGFfRzvJTl+14787f5vhyDPVT
4KT/wPn4Zgc6KbW+nEFLxplSkrkhAK1wVW4x8t9Kwe5H7rvvvaWPe3xfXH5chDvl
VKHz3g38SdNBuw9hY937yxcm4Qyugcu0x4Ivbmdur2KUU+RFxNyf3AkfIbxlM9UP
Fgfyr57Vn2WFCqi9RSdtN01XVUIcFPSgOweXnH1AxA3besqF6k6v2CPH2GF73dZ9
lS1W6onYIXmPbKdR+yV037FwqoSb+XfFU0cEHeNmz1NcswVME+Vmo6q/kPNQmhcG
6f6B2ZvGF0yvhh+XbHhQaegl0AAvROI8dsy008jk6HD60mgIHMBheXlEk7e+Fxy0
Sc+78h648Ps0Dpj9RcUPFv0IvIO6AIO3MwbimdaRLsO6mf8IdPiCqUYoijhHQjEq
ZeEWOCV+OI0Ln5EWrB7J5S21ZrzywX5XcIkr6psUO+TOPwmoAQteM5Ao3MXlz3h+
lG6YDAmSxayt7CBPQv6ozy3AZVPNORQBDordmnTMVRoogMKkxVUZd9p6mMqmo5Wj
yTTJat54oladrrDxri0M5xVqjK46/jKRgCDq9Pe/RDBqJ/5kT5pf7rwS5B9TZ7hp
6ZY14rtVURAcb9nkJthOIGeqZpxFrZEplGeSg+Nro0wcGpXMCo7EMSDwuCKvS1jt
5fvnM3rmvoFSMsh2vOodm7cXAUWp9h5Jk06nZYTQAAbsnGijoeXrHTh8Qwc06EqV
Vk/dCHVbZg4R8Rr+UhglxZYH/HgYhhgAPf4jRfNQBTsN3/23nxAMHk5NUVTbD4/K
gbFh800xb5CDaK/AsTXtawV6eBs1J4c78q8QGTCx6IWsy/nJtzIcgzdGm95ZPPr4
QqHS7tJ0tTy1ffkEnZR3SAxW9GRaWYgdOSVUu1g/tKQuTDf9dbpMBX5TkQWQrdX4
uqrDx41AvnpijnJbmSZhaKHUl+m0TUcPk7ieiVG9S00CHVMbkOz45kw/zOPYP7kF
TC4vf8EFszXftdXZ/wip12wnST1Y4aZ9kYp2wjD1sacH/NCRbp5YbKc0XiuFbKGK
e77AAQ5SLYUIgjeiajL7DLG5Kye6YjNCD71N0FzZia/DUJaPJKU/TpdUFPeihkFl
Hd8qXzPoTpfCDV+FUi565fm/S6WigUlCK9IcqEIvESQmp7bvfMV6TQno2YyEEUnO
TBTAOS/I7Ryl688LoT+tQ56duLu3haPdqOPsO1vTMyBY1ntvIVn/6xgZryuK/NO8
fQl6X3lyjnJt/FCXBOAUgYQDPrIBLnggiGn8no3A6SAlcomXd4EU2o1cXLbZXLaW
pNeNGefg87dl9ZSBFODTha+wSXGxBzEofVxMR0rgCXlqk1JDsgMBF4WlVhtm16dH
N94t2l7f9sJorlwSoH0jVJTJe4aXZ2+BFS08VpfFwM39X6kPxlXCb70e5xqG0DbG
nOvcaNXDKiC4ic2PviSgm2DSTXQt3++FHL5JdKRDY58yhvt/NnCjKEgnS79wvpUQ
PiUJuSDuPhWXF3ARRPxuXUVltas/XnDoqOJLOySRxmc3i5ocYvCpCjdJ4VAfjJdk
b5cqFBK42+jRuDuSR4aHf26rnkiZGoFhVmU5CRUhOMGJ3vwMo6BqKSR4rhCim3Z+
dbEceewYqgOUqC1u/G4mCPb5ktKiHQK+l/XKMYqbR4ozV8dMpHLgNujvtas2jj+S
fnFqR//+YAQElPXtFKeTM4M8iLPfPLkZSUbBXmiEuEKCmLO6oRNbwb0+HGGmA2NJ
25i+L+tAbxiaixRhMRSAq4VLHvWfcpYpoob3HB88vznqDvdjX2QYqQi8v0yazN5o
fnO3nxD2IzX8yqKjZGKDDnFEhbX09kDXLfHhAeq7h77NXssq8WIfdyfDgvBJXncD
lK+3h4yCIofPNNQXa/lj7s+TWzU3eGPX3WPylnOteyUPBFZVLwUx8CEhAKiRnPHv
p6NskwX1N7d8rwd/wX9iWutNLmvXlsmTjCquB+VOSpQ2Isf3KgPS+zZhneaxzDOe
Gq4FYa2ecVVSEJToa5jpumm/3nsfoJv3sYb/y4pA9OJffFS0rd2tdhCHAGnhMA3l
tH817+H9bVDIxm8fvirFhY/UAqMNBqNDyXGavUhIfoP+CsIiOn+PSh3QkUB4b+xC
1ySjDDHB0fzA4SzOLpw0YEj9pbd4oNUF5lisKe6ItyytGm9McZ3aKFJUVQx0KI5p
+/SV4EGayMrNCO6q0DTyUtTQHDqKEkzeDOY6DVYdWYTCeZcsM6TgH4z7VL0Ks1kh
qBYi7eA5jV4XSf18h1mk4xyJLuvxfNq348LmncLySfv5gnoYNcNNqb7HaAsWtj7Y
hKjHajdoAU9KiTbez/7gL8bE/KFyn7jFQBdk3upVrirlMv82VNxD58dCRb+JwEkT
Un6iKfZ7ATn8gB0NOdaF6Mw+qNEQl7eUtHQciwoN1H4YHVEHG6Agaavmq2Qvm9WY
le1L1kLl6kNoy7WaDFPeLmFvfHlvVU4Dkhq3l5wKAnJaIAb+hQYit8hjaF3EUD7s
f5wdwAXEs10LvcoRYOMoFMMP81jF6fSfy3lWoAN/IuZkn7InW3+/ECs/kI3UUDVZ
LwHOYDb3Ozg0xMIgt1hViNv+GwS5V2rroMyKGp+NX0jK3y+vzRqN8gmAmHRxdy3e
xvGYRJHU28a3L6iO6vFC4umKrEMVLw+q3+rV0WQPtlrlOOzbSznbVARqx0azewvl
KZMi2pheW2+FGMKjwmbBRtZ04tH+HX5YP0QHMfvJXt1n4RQq5iL9OH5zrJ7d/S23
iINg7dqHobqyX6J1OCNV184Q05Iw5/6xcYDBMX3+UpsZ2PX9NmXnRP4BSwO5qQcK
vjWkemOohtiWu2fO5u8BdR/ImcqEaaTMEvBzhzsv2C+c/HHnsXM7/F2PhKZi9V2r
kJ6jsOwDnXAOjx/39fxzDXheelpDgMBCkT595d6cy4Khe3k2VUXhSd1upxwrm8SS
w9WBgbDdq5wxPXkCQLFP1NEthEaaRBorxpt/gBtdVeGTI7UggJ8AjjRUPPBtCvG9
kMGJB9mde93PRPJVBd6vm8CV/RIgBVBHD4Ogx59qNTQ30OU6bmZql7EhHIHITaLM
tchXhruY/owFEzUJBCKiZ4yhdmGnpOAoxEo7qYePKMPei+MCL78pFAqL/fx8EZEl
URX9bc9PdvTt6zxPeI4PyTPSiP2d30y4CZ6aR7wQs04pzlUmfS4c4DvHDtdTJdEd
v+/7PVTCxYaImjc3RM6RSGnkiPNgOqgQTIZW7GtdY+ZSR/UVa7M4wuti4WcXzl6H
7wRS4W6edvD2zAD0C3WsvgIteUOyeeR8YES0La77Hvb/MVGSseeHuIuD3IyiQSpl
CSMDbGgeHDpsXSl04m7+BPwtofpRAvcZd1ClvBYW//7zoEhAh8spxwsCE0hnfawj
T4XA0VY6mRsIEKur+IuvzHXqrmXyIeKuo1OkHK5TbG92z3qlqrx0YbcE2IbHlHFH
ltS4ozyoelmn+26ABo3cZ7tv3O5qqSImZc/muABIScnvXIwZr41FvEoqGyvZ9kzz
hNQYS68k7RUfzkl7inHGAgmNK1ZoEJYtR0ehs16GgjaDBB20BRPZGqCj+6n4QZKN
0q5+Ox+gYMb38u4AQVlny7Ek7RcgqBEKSz9sD12OgTDqLFFL8n5ym/hsZUl/7oTy
Tn5kOwPP1m1UbV85ViWLrJ9ZUOQMEcvCNDz6hM0CaY872DHcspQ6GcuAH7MJcWCq
D5JVeJPpKmrqY9e11Avb3tCZOE3tnunSrW0Y5Wirl6M5XTMyouyV54MiCyqQwJEK
dSeuSR2in+58IxUynWobNp9idfKrcLec2XHAQ7V9K/ccRaESkUFlwrxWcxwJcij0
Op0JCDpflP/JjGn4vcE2HDRWzQgZ5lLy2vfvgnlF1jyZxWf4dPaz4xFPj1jARaCo
twzwaR2Ap95lz6781FTeMhMIkgGHNTAE9yvFXdsw1HwJUE+xUPRlsZ6vilxt2BeU
Q232DwKQhxHkKirj7WosRxF8LoCya2mqdsGiCF0Gf3SuQIj5e6oAdIpjkrW9AfLo
uSaxPmVSPpah04U3oSKxQ8iAsfFTHUZAY1Koly2uZzswbDv2zFG/xa1pgoDFj4Sh
pLfhY/kiUjtAjrxDfgdljk25su2UF05pUMJrsveEdWoHbbWozD4KuxvYK7tztHvK
46sC521wRxxOQT4D9fg47OODnJ+jW+oEmEKDykhW3Qiu4gKO2BfV5abfdIoF6fVM
/hoH0L4KHzT9vPVSoBtvpNTgqMdiNIlMQzDahNxZE/kzICYdYYBcHMT+gh5YmA6o
2bc1PHjRvhBwjRb6wkMh3NO99q6jJGp2a/6iPc4imOBOHHzQ1XF6ZsF9CjmHe2a0
zwlQdf+RP4WvvEJXslIwNfgeUnbtJ9CAZCX2WLkJZSCAyxpX1vOttpWX0iQZKMAv
Zkfk9dmQDA/heiUNsnA+PUv7A3wlI3PpGd9txlejNFyO9TPDxKEa9moXjRSYb4cV
JDYtbt0EPuY/S8/eapzAlXe7sBTLRlMEvZFn3+dEMyaHRTtvlILk0cJ26D0XxQf8
HDgz4hdTAPhddBMCEs+I/ds9tiKvQneZqGCZbH8bgh/RWaUcdg1S7i0phuGCd+vg
WGuOL1MSu7fT7wC/EH3UeTdSr4150MPtBrVrINAuFJ6Ng0qg+ZPe0QSmPHnPg1CA
Sc8LDM9wzJfB015EOf4VAS4h6d6lv0yYu+8kFtV4Kxl2z0SWhuN2aowWZJ5o9nNk
rAV68illel41OWzmLK1p70heuLGK7EFBQ0ByxWxxB8kaGnaMqfIIDY4dVMEswCUj
pM4b9RbL6tqZVdoOQ/C0DRanqp3bfmQQr563984tpqU67u44J7QRaKcQWLu7P76D
ykSbR/gxesBVadiFOQ1vMLQcvtR6G9Yf3T+aEGAk/5Px22Spohzn9c4jFa2/N7ry
gncqfqLDlg4uYzxTWt3OKhvj3GMagnGXDbOS9QNkNzSD168mh2Osn4A5Vv5MeWF8
SRPjm7Vh06VNBcJF1rXxK9TsWxnbaUD/1NGk7+iiqv/NnWrvLaCPdFO8jI4dKK/P
OPHc3/6e8y1K1/q1fEHUBw3frt7cUUaR48zdNkpxAqtgxxShI3X7mR3CmJqDjGAH
FCc6j4cLTZjGEWsRGP2ZM0sW3SqE3ViEzU3FRgVo7gEJqgsDWj5HxVPKc/dAN6pt
N/DHhmfjdWY8Frnf1lYN+kYitsFZ85uiRwuGDFw+bA771LBG0DzrSFsZ9AC/c722
HdjKYT3buaYHzQGi0Af7Ef/oqwUmxPqDzAsFp2jIh5k07eYQSn6KCy+yESCrGdhV
QTCXcqAvcEH2bJ1NoyHWRhARcU0qsVz7JFyxBl9q4dxzN0Wt32g9PXiGIgoO7+si
nftErrHRnJnEXOg+MAKaZJcQolkEUE2dBrvksrLoSWZBalR4W6/tNNfofi24PASE
yHDs6kD1AxydqRqRMbzj3ZR1EmZUpd9KXrLz2QMK712sAHA5Kji9RgNX+VfJeJoe
RyjAzLnSNvd2Jc5j9p6/2lgFRPN/A/6r2OdyuWfZx2oVDBxY4SILCSZ2kz6D53eS
oK1eFw+au9zmhKfgnh0uoT131voAPonWrZxje6i8/w8ssrlxk3T8qYHJwwtydC5d
/SD1CznmnerJgpJRkUN3uVO2UmP81Z2Qm0Wustx+4yUrekgnrZ3mwjrokhzY/arO
ZKitjOCI9/At7TBtapOaaH+13+s+FceRE2XHOEDpAcLj8pQXAOXm8cKc4hD0btiD
Z3dpSvv+zlN+h/fW4f4yPRpTOtCJ3O+jWB051RB6L5HQ1V8HXYyjOCWgqF/Kjitm
NasReGc+w2b/Pno7CeOt7qilUYvOwV6HoED+OEgZmV/3KtbM3D+FQRZ5K+laDQax
PlBH2rB9bQj7FhSlxivZWkcl6hQUwLFnsxA+FkGJGhlTrzctTufUn65e50vE5OMf
TJRfnOEzeMkauYcnVVOp+pcIZuVQPWh7K/aWlJ/WpbPucPN4g9UmJYAO5JkwcRfH
tZLQKglpUY2e4sjE9D/aygh5QyjdKhHF9Nd4DboNj+rnilve10foJyPJqH5n52sA
cxAtw6JzgVaB7r4sWChNd/Yi+w27r8+6XMuQ8BPlcAxIvBkhKOWMY388pYBaXMnw
VA+FeXAGPxGcbYkWrbkAqdo7f3bhbQ7tojby+ctOgmOOxFbLVlAU7ZZC0WZMEkn1
in4EzCHeZ0pA3KlreVoVZejx5CCl62wJcLBe6y78d9pcReAb+bLgrv6+7az1O68s
Rn3wDTcWUhHwLbl2Ixz3fygGXhuZ/qSUcWNUSJM7+su7Ed9KU6ddZixxcY0Kctwy
9bsLEtUgdnp2N7VpzJPxc/DBx6NYzAMK2ct4TwCID1fr/maXlbZ4geRVYKhyrxRy
5Z36p3lUDezpBbg7cFJ+Qk/ue9IyvePDAnFW2kA29oaK56fg40xH+SD2SwR3/9j8
hD6C4HTnLs/N+TXlHQTd++xN7P2Iiyix57++yNHODArK03gFToS8gWN42nCDbvAG
x+U9iXIVNZDOTq0/nCswTl11qc0R/ySi9ZS/NvrJke6WRLT/QPu5sqZt2wc3vzns
qezoDNSONV4UlIKs2mqiFB0k1ZM/UGngG0TagZEwJxH91x0QdZQOsiIJKh35QBET
4a3oXCRvpGrQJfqR79y1zxrwAtEQ8R7pboJFOCZzTyi3sXSZhlCJmnB0+xRfJcmg
IXZ9wH/A66khqXKMloWkc/TphDC7hujFstULYXlr7E6ylXm6ipL3JCT/XpAcxtxH
lzJZM2r6h85AW8VG39MaQJUyx/VUn3+yXJx44GTMIQ7+G9KP+dHY/0h361rIma3O
1zJNBB1FZTAEvpVJvL4zqXKqgsJpCV1ZTQGJz8zKViAhnuFfyFD3Vxncn17jKtr1
sOnn9kYBxJfASaMFFjnEJVoeyLNhKKhWxWmCBEDXHDUUld5ulREUbJnYlDnc8mrF
GwIp9cUWA937ALSP1kc7SOXvPH2g1K/9PE6xiu54kzIaW1VhRbMivmlhA19ooP3k
oN/1KR0oIrVAfRe+yw3IgSch9uIaoyysWlZamrZ/zLKKjYyvsd2+IXVoAbOtNm7n
1YP6rocpScMVI2MoYezfdRSFshlopzN0I3vPlSYIUaac1WNGHEG/rCezBOG9lTjO
YIKz6vA+QTvd+eAqxkVQIUYwMfOLYBhm671OGuZwd7arOUS3aryCvDg/aXqSvGpu
pYaDgGXvx2anGFqMHiPTC36Eg9AVw9yz3/1tK/tpG3DHtJloEPYcegB9ejTRvsNW
9LM8Ag18Wl6QsNDAO0ukNa6khENwVvZ+yFOX7vHrpMWWoBSFmmJysgnD1CPe2zHH
xUFJL5KIPeYPmeFZoeSvjb3ycQmvFXLwTWu+7dxTEFofr7jPiYw21/aOY3wLBo80
5GYXpxXw3/nhnXQ518SgDb+xpdRh0+luLaNbbcB0m3ePhVUWijBjfNxuKXJX1gnv
BtIm401e3NrxitxqWl9Bhieo13KcBzs1pC9W4mvVKSI6l6DrjZSACs+j3QRJcDQD
YZ+BsZbGLcEuNw+VMuR6//JggZLBp2JcumGfyl3a8+Q368zXsIac0G6BBd1nQEHC
b2HmhALtUa4fADjhT+j1qFisxbg2X05kljrnTj/WckKlaWRxb2/FrXxgmUA1XEh0
o5tU4zIdgdivPvU+gTW9akDw1yymVA1zd8zaOOMUJLHVps21m5+mJmgclpqEjB3M
xQm408HvYH2NlbIAQYFxCOZCXMw+88pCjWSOIeBjZ5z13iO5fsM16r2n5BfaWHYm
nDNYaQjq/lpk6YuDWgoOSmZuRNf9Pdrtb2PXNNX/fw/bwTBw4Vmvtly+j/JbD26H
Ztqg9E/9uWgolnFr2Pt9ymuNWW5HDKrVVUbGf1ZnzQLU8W+L02STqxj5sE46VYCr
TABVf2B+vFcXZ8nLNempdb7BoZQ77ON36OAe0aMm1Sg+XpdE6ifjtWM/HRD3zdfL
19yICEiZXIb58QLwg7jIELsXWaXD5Me/EhivlgphmVnB8k3tFMiUXKoV5fuEvWNs
Mr3FrM5+uR0vxlmIGhbyGrmH7aT1QIBZX54jZcd+Sq9sYVMSkJFfFS+JXKpqpsJj
UZB0Bl4tS3YwkuIig1wBoxb9RqQHw+gUydSxvNiNbI06tm1NzZpbKNsFcv5gCKMX
zXAaLnzmrZ01KbdUJ6zP3JrpVuOptwujtJZ7lIvDT/V6+loxdZvmKkwmceyyhZM3
bTDvtJm7/jOCj5DEhroCeTt6MnDWcuISTKug9OopElC6n5Ja+WXfRiiYlZ60phiR
ErRw3SknrG9BCnXO3VrLTdR/51Ou4IzQBXyY12EIuPWcnsGX3dkdbkSkOd+awHui
SSdsvq+3qpSTcNKOO2LjfhyjaO+EffwKzV/VGsUe4iomS54yP0oGzhaPi0MZ2mJ4
Quv+z7imICluS/SzArbpjl8hC3nXh8eeV/egG8lsWlYOS6hTkGQ1AyPaR+LUgBsr
GBIhmhll98Qs5lCvu6YXlxteNKPdnAZRXi6RiDbcAc3SvwdEIM71UW8Yd8O+9DF3
N4P6ntOflfqjaRZq/D17073G8VO3ooGoWb91BzAhAx0bk74jzzoDNkB7PHP+coSG
vKv6yCoe5d6s4LHNS6Ken9kH7TONGL9PTx5CIy5JlJxl6SZWGqAr9Hy7pJbidKxd
YMLnpKKcDLtB9/Y74nJMtW4HXib+X0nLoXSKiuVbcva9vtXMjUUfACCjXa17G0US
+S55NCIWyxHxhzV3wUtgSeJHVxGxiZobH6OuPnxHya6+mPASywhnVVqg4ZFYXEtN
2ujRSVitEq455yxZnwiFu/utSLsWj8NEKkYWcNOm9SboYuaSJ2JCrG+f25gpKAuG
LQ/OZS641kX+ZE74mYjJyg64y0yzlDvR7W5v8dGenaGE9v+eltoplR5y0soxpky0
YNCmCfifjJE8y4koxLlFaWXAb2sasr7yMsNxpJnlPnxpS6ZoB3gmR03GTPA035o/
9/ZBpJkcWcbxsjsXoVGp16s70jnqC+MaDoVmBXGe8CbqMo6Gr45GBfS1YM8mmUZv
uFfUGjQpWF4HVnEVtvD/PiBtxVbolcSLnBzIyB29swhuIc1+BTKCDpLdxLFVGY6x
atnr5MsJSKBTPq+ec1GrBnLBCOXk0ED14/ZcB1aklFAi9iy7WCYvV65aHQoPuI3A
aZN5Rn44gvOFy95cCtcm8DIXZF+AenioKivmD/9BkhdHJJOg9q6Pmo6lpFck8fKC
YtYdMj9hKMyG1UyJHAmDA6irYUhoUyunQR2p2w1FusQ7NvLpFaO8SmTebo31g884
54RJ2Yr7fZ2fWAAy9UHBxmh24kDT5Chndh1NlTH2oFm1BdokPOZpuL4G79hM3SMc
ET4euW8O8LmnR6o59IFcVuXuqAOuoCd/S4e1KUEE7H4XkgOdc1vkgvcLJZ9xq2DM
CV2hEhgWRJ1mbBQ6MtZ1g2ZvhUa+TSzllT5PmTYxq/BATKdjZNawKXnoLLLBCPqT
saXvbFFJSKziz0ZgnRBgAD1UlaK9SdFRdVaEAnbcqVPuBtUuq9Mu2GFOrwzu8Wkr
kGHaeNfIF68UPes490raiJQAsLa04O4Lmwxp2bj8da/gJMmPUvFVY7+/VJ4pjGwQ
Jsx2fDHuz42BeumZMQUrLi/i6C6gl8hbGq6N4qVNRpkUFFvRyNW9XYeIM6K1VMi2
6gNQu00D/Agyt4IdDxKHSLMON1nwR0KB/CcJNqULhunDd8nNuTnWPliJDOTVeI9V
OIr/9CQeJHK+f0/3Xd+48pl+yHW1oK3yOmqHwVh24IAvpmNwVd4BY1HKYtzBJ/jG
5aVtIltDpyc3FBK/0jmgPeSIeOat8AtB4+n2k4D2VCH5Z2GNrj8k16IGTZMuv9IN
uA7MgSuNorS4AvdDcGTPmapGEB5J6E+Zhs4CPTE3J+iQzv4mxBCoha2IDaQiEbnb
+cKKJGKv2Vwurx+bYEsjSDs1ua9bH/j1rEOKnyoSZ1TEQ5815cM7+h84oMn/Dh8V
xatmkIGoYIc3SdGzibjKEZOl2+t2Pdw0saisBk3mCh8d8gJSYP8vbYB8jevVGwOp
gEBMIECxFHKLb1spSLvnZL6bB1zmbdgf1xg93b1/G8p3TvBH6GKCmyxgbKi7QhUU
BoELwojqGYvqWbjBfssf8dUABFfGP/9CWqcSBGbMSn17NewjjgjJTsIJhrm4lAQ9
6hsNoc/kL5iNzvTR9WPQZrULoqp32xG0q1Nfv2t0DaQ/jAUJcOpmXkqjPMHvix/N
lQlvA77ba02d6lEjV1uaeJ/3s7T8LrFFFvjipHPXEhYBTtSc4yckMiWOa+6cOVBg
M4Iog33dzrbXV6briRZgCyCWjOgE/KwWELN1JqwBxtrw9Fz7ucm1C82/D2oXUWqR
iw2mkSVkcHUsCFHN5e3yf74s7BuBHhFSW0DS8HBu2mmUVSh0t7P2Uygmxjq5wpo1
RiELqsBXKBvFF0nHTOASt5/a7yHhTylyXK/nEN9sLhsjwKk0ioT5ydi9OK/7Au3x
v0SA9eHGohuwHLAJRJot0/bMw1E2ua2wl+hxbtooF1qtLrY43mbH446avltKIiHR
z1q9yLgjCjxqYXV2tVMfn2UNG8tG3EKloTu/1CZGNFO7CEKuQrphcs/pGok/ys9x
g4806EFbfLLm79f3Fcm6v4+7mDXWzABu2Qte2dR5ezc67TFzpWeZvHRloLAfeExB
u/tXDlxWih1UBgAqTUzNHIVGCbqD0GydHMIlNFjkMIqj3XbXnR+9KOWXrbuO+vqf
yUG1/d72sWt/0SHV5nBogjGkgTCpxhtHi17ilAVGGCQKGbj6bRuvqJ0nJ99dDPpW
XGlMIcEbV6FGCZWVdf+WpcwQxkEF9TuX6taHiy630lk9IPduFCpTyISR0Kl9WX7F
VEXZ2d5bbR+9F/jaihWT5UHmClYj4fuEj9PO58xACEIcatdGuHZs2e49jJZDSQAq
Xue90QOrn7EbUHZwgJmmrv973RztE+NM7QCNnM+CngrOO/eBVKQc82v9J7cKnjWl
uZ/6fRyZKOOouI1D+B5m6fHiijI5NeaBgNG+t19DRZMi3mqneZraJkiH3qxwesPu
H0Xzq9c8nx29vr0FuZ7LtZg8BknjDpKpmU8tnMcNjQXo9cvgN5sJ7A0o+BQYR3Xj
79d3CT3cUMj+K9PoMxXkoBk9iovLgc9rlocQfXJCCg7Sdwxh6yE9QZNuZqUTmbCa
wLBVQGPOlwjLYP/EcCpMwDl0Y1DD4/Lmtq3vvnNlXTOpDzOEX9H43FDL9xf3SIvr
XJbLtFg1+6hQcxKD1i9NqHaS5FQLVFZ8vueENHb4O3hL2CFc9SpZmgin+UahCcKx
BruUNry3rIWR5jdd7kahm7UKAUT26xftf3TsrzMYQcpI+wrZz4/K+rwz9V+wVLGq
mJLcKzDz1L9XZG9QH1sqMBFEqc2MXqX4K7Pbi8Y89Brhq6P3wFh4V/WB/Jn2POcB
OazsL/yDS1+LFBCp3023kfRxCtkBoTbXgWUP1Fxqb4bqB9had+H1qXpW2siunad7
vhyD7Xs5lLsyTNvTV1DBy7WR1rd4b9U6Ke7LbAHFs5pj+lbvZvHKXqsZGHKURoIs
3kzFNIOK9aeyh0cvsSGHmMExxpeSsFdqRFgdvPKI2Xo29UV7Mt78JiQdkggVKtD5
Oys/sGFsddranwGHdYZQxwjPvpUA+N8+NQa4jesnkiY3vPKpVqlkm75DdGirbbvP
pw7sD+tuJcMCW43CE61pqNMb2xzUY0zkwr2zSNh6HbdEddQpXiznCVmPK0z4BRkK
84waY+TrMHtJHl9JdYN4wtLTFkTEWUzuyVmOaYF6AdYtGeM3GZqAtkMnu5tccLSS
0xWVKrWaGnwK4PzvVmvc9zihP1e1Wubs4Je5jZOYQcrXE59oRbmiAlKk7XUTz8yE
/81/qoqcAYFUZrpuX7/P1oWu8NAGVIXJ69E7y1r6y9EMp4B9EYzhScr2WDkl2L2N
ESAjCqTiKVz+HWdBwSUuejbX1A4g5INncjkm87SMwqs1zsDrg8hWlsSrfOsmESf6
8YF1S5nX3+t2xesA7A/dD4b9krWe5gIWfiNvpb7cxtgXpOoO+yZfFhQt+W5yyk5R
/qnSaFqZz78/PDT1v4/Xyu0NFClUmhriM+Z6oAktOBOojVwPYh8AaQXyUtXmvpST
KLVTQxIu6CtXIOgZcQynb1jvppn9hywPpMsr0StmIqepwbAeI2/Y/2/Kz2TqoHYG
oq+91CkubxDARCSeRyD57wuLXDldKf29BKlahzRTl5ODWv1P1llbkfjhdACnhrYB
jZ4rb1HNKDGT9EWTPV5B0BAbiR/x/elDxAkaiRkGHUIVcnrHO3mTdsL+mHzVk+D5
/LZh6A62EIKtLYbVqmkwGPStyRuAHOsN7xOHxIvfUNWpopk2LoWbP6G1mavbPN9P
UrUJfUdiZwM+pCSaY6PCFTubLuIHj1usTx47W8jsjwm3EYBa+ZwZlIZ4CWGnEpTz
7QiPN4b800DqOJDGqulNZfbH2698EV4VQ4QBY4o4YBF3IRpZyAvWbr4k88TmrSoX
okhMkrHxHKAhRaDbcD6GX9B9RD4hYCO5UvGmgIH6jgvl3MXTCETNyBT8fxGNSXK0
Iz8xi/GJ6YXHtQXzW6RaTnvBsd0D+45NVI6WQoFtQJDQSPL3Ecwe9zyb2zzDvR/5
t6MwdbldozeA1qLl1RGvEp0F55rTZgwk6zLb5dGBy4lbvrYneMZ5THCGYc8wnjc5
dyXVB10f+SzTnWdGeksGH3u8/liasyVJE9p9X7ZVTrZRwfEQWc4ssY5ewT7vtlb5
M/CrDVHkXXYJMtJwzRmH61cbOtwfZ1+bGjzEX0+PX9ml2NQaWqMgtjlv0ugvTYKU
89BD6125yOVzCPoFBZ4/Gla3NZxB2NOb5xX1SYLnBIS/mfkoSBq7DigCfrtKdZeP
7M4MEyI0rRnLs6/v+pA5YHcMdk5XIO73KeEcQVuQ9wivtimUHrc68xk227ZmjwGc
GlS4jkH4DNVxCMoltSkUcjRPcV17yM/JKdQyPo1phSK02QXyiCJaB1SSVEXLhzHg
Yq3ernr6e4n8vpSehzyY7KGwCNgwszelOCWlJFXg6UE4XlqiuY+YYUTUqGujSMbx
35mRvS7HYz07OkdGT/fW1C3jH5CQdO3UxaSrC4wa8VssNBeSKKZUYMnnYZrVxYG2
dR8AKa0Luvs1MhiuZz2rLx/TkvOpQbcGYryodHDTu6CngIuyPPg2CuO5cwqo4gAN
gZM3OixZcS2AZ5FTPsVqs/cy67EDx1aAiwq0YksqYmmw0GznpYIR5XmtOSjBFFUi
1VAGP8O+CZ3NDie/D1fcO4bUsCdIIWX2dyenzYu4ZobFJGXAEGt6NxMamX+Ip2Ef
d4NJ9+jZH+laf56god8ihIWz70T664ZMMNF6fSQ4jxma6JKeYHm7C1S8yeWGuDAt
qUxgBeE0yflMUswItybKc5lGhUMdYQ/xDzFqrM+a4yZv7Wn58F902mJB/tfW+a6H
5xGccMLB/vhWfNpUFmRQKKweyXOKBmX7xLHo9NDZ8yaFrG/a5Z6DpN4RyEds7utd
k73F3vpgJSAzBG3+tDB2n1fqZtVRs8sESnwqyYT2ycbwNpiGXl3v6rrPO+rVAXIm
E63ebminPstFOXHN7I1TdhgaUcZ82hNvYWq8sIaGeu0AV3JnirUBay/SjTDq2V3B
byEEi7rNrgCLvY7doW/VMAIfLgOr54I+674gBVF7o5nXMPMcYScDS2PtmXKhpZ5A
TqrQO4HH4hD079IeFwDTObareWLUwPgII70lEAdnp9A8JAMJwqdkOJLpjJ7y47st
EvWa7JVqa33o6EwY6VloM8lUZLM3g4/BQJKTmgqglz2l62mU4NmcIv3k82776URS
BPB7hg8rDz0oGZE4rAjFATajhb7l6LGBCIO/5ODOJSZP5b5WkKP/kV4fZdkKteed
uDbnCp5wOgaiYF7N1CFyKSCPwlbKx3KI1sD9yrR9n13WNO0T2gDXKrjPAyRjO6pv
BfeIA68rm71nf0tVyYB2bqszrJa0GlelxMfoDBhXi3Z9HNUyu5tYC0q+14zZh1cG
AbXwUuZPyneIWZWYqmA96Oz5JsIAlowovANhO/4BYPLwvFV4c3ENY34yH8xSbmes
cva5zb/xnu6aujOSi+hnH1JbHWm9/0Sew6iFHnrFgDpq6qS59fsxEf5ZybmPzraK
hWRv4GLGxxpO9JYhvpQM7hPPKMtZRAqXbxMU6MH71EplXjO4Q/SkWMy+wM0XdRQB
Xchj/jNGnK7j14E+IG0KrNmHeUNE+r0XeDgJkc6j9oTt5AdnB5cQVdDTACbM96R2
HnVQyNCJ70ETpMns2BLATtsr9zN1Z+/l3V8V3GlKGY2NyCZuYRVkVHEjCdmkWBPI
z/x8PKFNexVlvg+/+sw8eQuYZgNFT0WKh14edcnPQ31ggqS2CaTrxPsicTkFGRog
8aqUTsGkyAq1KOd5q2JXGw1ft1h6A6x6s1pf4zqqHccLJG2/VjrHu6CR+Z/jNlEq
TrHW8fkZRKZW1DgimVDtxzDAZjbyWftAYCHmc/UCLv/SguxCiPf+gS6iENkJKHgR
3VWkCQ7M+BBGckD1P09EspaHJtPnUzvdwrTPDdi++fag4iDr8ZzdCWrOz6apD/H/
rDsWVq4mCBRwOFAuHUipyvl3/lLBoCzAZGFxVym+POcC45+9F6D1k1J6tY1QQw7f
Zs0zBAkgrmGn4Dc5Sr8g3MbYKYoUHO+vsKvEM2P/PQtScgyue9vDtnF8z4xUUDDQ
Pe6AVobjdJ6den6+6l8OaigJpumv4dvqzvuStTmbKL8gxFAh04gAsLkeYJDhvslN
J8G7r9S0czcgvvzKCYqVozrUldNOjT9Qyu3xQbPX7+53kK92vL7Ia+tddAoCytrr
ofgYAH3bXwWUGHlv+6RBzVohxHXyUUGyrtvgPxD1se31cyaNu8ngvPSuYExqc8dS
bx5pm7pVjFS/vRBGP3RkLJpVlM5fYAoKMDlL5CgxzPgd+ehvrOHH2uatrfjH2vle
Ac1BWEKp8ewo+9UQ/FDNr27e4WwL1TprrFmvgkeRrYLNHHVxaJyKV1fLagPqo0i0
FK7+xM3N4lAfsqTSBPiWKWlSrenGqUL7QoVS8MRKt1vlVWNRrB/03SxkIgOBGzpS
Qz754u8jKOVyEpOMeS9bNIUPeq0Sf0RYapoNkvngY1YGtSfh9/fKwn3IPL8DzPzx
MvQOQYhZAGaZH6EFdTpRzloDDCeEQ17L7P/dA302TZghs1mjKc2lWaSmszLXe++L
YHxQUy1E5JFlc6iiz3YM0CWh/geK3fE/sSUO3zFK1I6+Kx3rI/CvFa3xiGeXVnB8
sMlcCiRd7ju9HqiVAExITV3yxvV1zadreszwIu7rd803FtOgnymuP4u5FvAcB4UZ
ZbuP087KJ1UHIcKn1v6z5NhNT6e/+eEgBHSuoOE4IdP/2Hd/1sw+jdXIF9nXfuiv
NTsn5BFLJzEAPfT29nKVyCYbddUyEG3tEP1Xni+aFs4P+Rcc+EtHpKG9s9lbsDc/
9POAonKnP2fXopW/V6u9Z6HZhWyx+43zMhT/To3A10XF/zFold2OGMuFsJg4Zc0u
GSvGAedrOy+A6pRtW4VbrPEHLrKr0/vybgxPfaFV0AOQ1TznPDtc3/9YjkNrzwKS
GVzOtZddclZOXPdrq5X1j1wfwXMYoTC/vYeC3jCQDk3pyLmN3u3osB3WVpmaTnz5
tbwnlDBxdmnM+VuJAAvfq7GpHQWO2voHAdf7bFHdYDizDECiOfZkVXarritqFAgI
nkKi3vRmvu9Qa4pIl1wMwfxK53dspXbe/2dwCxBGbpQ/CrPQWb+MF4bVQRwXHD01
4LZoEvh5Ff6C5fgV5uAx/TEwKfcyyfAu7SMTS1rcrWO4Kcezy04aafpP1FsJ1oQq
ifz6AjAd+aJgzg6iM6UaAMv/C5BMqITzhfjLDW7+feGQvLKqGdHfsFC3Fv0FPc5J
pKFkDJ6dAWN/h0cBxYUhM/i92bPIJW3u3HZzj+CP2i/dWp4oJQabOEsD7GRGsE71
29GI7l9RX7fioNE126Uo4csYhDp9d0HoCGfEiVtjirBXk1giw1WZK9o71R+mPmlp
Kq3w52vRDLru7kW0ytFTybB8SPOEFmw3aDnKreNIM9fpXDCpSSXz8Q9Hq6pqT7EI
5HwRZGCv20kGM4WmtdHALs+vTf7wr6FAVSBLEwCZJsPesogbxTUPb1YWGAEd2FnB
EKmODz9ZH4nedhTxNEQGsFZrVlNaGO9Wz2uCE8bNo7cdX9fl1NamaeU08JqSJFx6
occbnvgWrE2LkaGrPT8NCb1g9pBRiivtocXWEBV/AsZDnB2ncR8dpcnD3FvjWt+1
86RnKVx7nZ2PURid1UrdexELEHuD9ovObTe25AWmD/fwP756bAsqw8+hKY5+muLo
keV3JcHFClZdfCKdJsE+1GccHE3jtsw+6KG1GqUABw/NSUy/6YdOxZA8t0BKwDFc
CtLqIFbnTCWvzSQYfjezaOgMcoyVG3rkee1tea+wiPbYopaBPsikCPdiXilnFAdU
WWI7stY5eEnFUhKqMQEWUJxz25+2L3jiRlqEocPczhPa91d95/6DOvJC+9LUAZ52
DxdYgvJTmMyKK2XX0WJ8YFA6DDYVZeAY5TeMw+u2BwXPApaf9HKbnw/34hcMK2QT
mrn0A6VPTVd29wPT7HPF+DC9s1kypWtqgoTG4gskziX8IHaoOVSxmbrk9QVMBviO
HrCSSpxMyTq3z9CAbKTgF8x69BvmKIbnl06IhyfRZ/FEb/GZExbwh61bm3GY1ccw
VBrUbOHlviIXtLdMd+84QY9cUKcUrYsb7Rb9YPkiA7a3e0sqmLKn0lbCEenafqD7
GQI9MGKBqOjwFzq1pJhyNlYROdcQbLXpx/2KRPlokdWsw5ULcx0GKMcUXIl2HHGJ
MIV42QSV2pBPXYtIO8p9Eko5/idMiCYGHsw7VszOPmMX0ogCg7eR+I+aNlOlENu/
KRH9DQC6BQ1Mdz7sjpLy7pNOZQTu4fqBzeELuNPuyFDq3Q/yWuR6lcAnL4DgCVmP
Eem98nXaglyx3fPmQzM0CzaQl8cDOD9bCrRStpifr2sRCt8vwWtakLSIdIy8TeHR
dbRkFFtiAEtuXreuVaoG1IwU2IhEaNgXM7TGAtgLl1F53jwEjjHIICGeWl9sqwwk
SfhBm8usPeCZFVobIN9WPdaNGw/D/RkXMLecnHUWXFHx8ZWAlRZQ5he/Sr/ORg9g
Gb5p+fyxP6oqvcDzDjEI9OI9wRA32m//UNVblOIenti7J1gmh/vyBuaLfJ+EhoJP
581l9uW9k1dHnkjO/v/D2jVMAnskEY0+swAtEbM6OgTrYF2Jk6bSwYxSve4d6lJn
sUNhdcajWUYeyHlCEuN9axCs0adrdMPtxEYn8QpnCzPgg0M3Z9siC3DS2ZCLte7n
qcXEX5jRAIFFC/RjbBQQp6Ol8cFx8YLRRdDmo/BC0rZbPbN60Goza2GkaCXdag/Q
k2LHMZqBFhEtrlyr8abzelQSDuloSDK6ge/JNLw739Cegmtfo7hVKzpRQRovegh3
EZ7S19oc9nd2fFPqgZcn6H3CrupjpOIDLUpARUh5E3e2ss0LjOFEfFy0j+8PEPDY
gaLQyWdSJxNCmIfx58pn38LzIJa1NJEE7XKcolhH1dkzdkR2HV7XXW61Dz7MVhR1
Bw54h7zOsIjxf0oDeb77HeZKYQTSO+0qnRzQ6O8kFZBbYR49V3QU8v9MncXZx8fd
+s4Z28u8xwJ+rmKCZ0HsbMa4CBI6tGvB3aJ8+8hL+Gjf6cuY3BOF0NfMORxy5ZCT
NVdDQPsCsx3Ir0BM2CEK2w9tkmRQF7YCscQgoqWWxRg01zxPw89ZfceNdLPL9qBh
/9ahCsF90zP2xNj3TJWh56C32Yf4s9LDumray04IJNGbSasgCUr3VU8j3Gar7deH
wdfDVEIV+OWRcSK1DMDhwrOfyo64ItKVFr47xugdSDT31pcrQXp7hrVE468lWacs
lcKyReQi2LyrSVtjkhVYMZpdOLRLS+KpRX4lydT062h4/xGD6rTyYQzvMjUWnZZX
1pAVuwyBFzf0JYrP1gYxCugrVxP3nWUWWKGQPp293qpNDKUD2vjEUXMyGu0qyZ0r
mTZ68xx9/wFVAtuynbQHg4wZVuA00hj+CU5+L4nmYPd6wj2w/1cD5bTBG/MhaFAP
ovaQwYpgnxgMKqCqlcGjF1KmsmcmtckSy9Gw37cxtrZG8cPa8TdsrBm+dD7b7fZA
X4F6QgKs7fd2ZBsRL5Qnq39sVaYIePpDvxrrW+noCZxrDxMm056gPtxmVXSWsSNz
jnnGi1FSEiOult80GR7OBFKyiUQKewA0uIbqICY/n8UMGkzDUM5Xq2dFoav2Ikkq
eipkBFF7BhngsEjowqbdUEOHJIg4RYL1zvWsXOcbBhs/KF6f96PjmBTWIiFvw6kO
iH98JSbJ7KivM7fV/FsmHEmOuuaEDG5iJpSlHPYUilTE6qrptQOk0wyw+5bx/i7C
6NWNXVK6JNivvDlOF2lgYNwXuZyP+RW7KMuAIOFXrDw6PRrxATNPGQ0GyKbhCPgz
KTJ2qZJhMn1KyYf8962jdfa2VhPoBowth2juwO3MZULqurGyRXtkjMANu1HPEGnw
ka9O6Bgtiq5Ag3m5GfwilnPXHzjK7+5xapVgMojIu+c/MxnSXKDfJivDERVJcSy9
PGY6Ta9orZENqObTVY8Y/pyQX5aRI6PHN++813qJ7XJu1N1VFJb5uuwQHTaxeP7q
fpdGddEUsMZWMEwEisqxFze4jQ1ndQMNF+1hVySspMBlbizlk6EgOQ/OFuACTyqG
mqiqZBSH/e+FQaIy/cTd2D8NPn7YCrRShE3kHFfr1aN35z5hcGkT20X1mWZcioH6
vCLRk35fLOXgUh747HM4pJ5wGrZM9ei8iO/0nRp0Xu/LJYA1U6jxaf2CuTo8hOwN
AchDtb5UlCBFU4PbiRcWVKymDUwMliu+JfxLxV2E+3SVUa+2eYWhcLwp9EFiHOqo
QU5qeNcS4F3xeA5BlMbw7ITrCB850KLnO+qcw8Z1gflRPvFDG7/oCJwHyogsLR/4
sawKoBZb5l1KkvQ54TZpFoXy9Mg6fXz7mlZmKx4GvksIq1N0Hf6jHPn281csH3GJ
W6Wn7QGqMQvtAfVXTWJF7seIVvuFhrvhZn0g4mCIUQrf0Zk0zcYNTeb7YpxM6bcL
GxSN75IvOKabza4RSTgIR5eG7xhAOsZIxZOKvNO2rIW2wOFK3EdiqHdmw3PaP7DA
fQRFNncPXx5hKiyRMWii94RzpE6IHZSRkhacm4NGeJL39vSp7doQqsUMvVEOmZZN
QEF/drFyJO8S9MCCNI5E6iilmfHTjorg28f0B159XWuebKxZS4lWL9WONRMivGFt
RB8teGyHPuhFeLeWB3XZWKpbKmKmFE/URIUI8pJbbu8BmmZktjG2n9EqDbQqZg5F
nK8wJMclUkwbr08Vhsvon2JrQWhrN/RfMz4AXHRzy4TPQpIDT+mU/W4eS8xjMCNL
YRrx2njEHbb7ZVOCNtKd33mkusxfBLBb4nHk00Uh1Jd1HNKr0S8cBwY9VcQp02lC
MN5XCdf0NxHAOKrj8cWEkijZQzrkQvzz2AMStYLz0ZVFmZfIcF4JWGfioXuBPmgE
vySMAghumS4l7GjSY7cZTTVurJcHX6mUUTrPntH7BsPQVw2wweEyZR6IrhpyCspm
+TDfqZ9r3CSC/uY6Lrl0u0OSjNGZjnjzLrS5NsSn95VyMTMBUb9yRk/R7Xcluomo
PT8mFNZbC9t17exV69m/wQSPw/6YZT9oGqdl9ddpp2JgTKf0uoy40KGFMy3SSxrQ
8x54+iiIrTz8xhdt9/uHQXhQXbncCJHqiO4AelM51942pn4dBg+gNmHXm9GKwYCH
XgH+eFCZWfpfBNzmMhcyZ5zhOLr+U/7I/kmtEe34gnf/XhfG26PsbK61A0IO/ZwA
HO300OVvtIIMNi11u7oSa1sHJekbtTvx2CXwhn5mQonfXXJDqJgMEomw2BeZDguY
IazMr26lfj506sMpuD5LO3bau19gu/wGPJyaxRa+RQmclSXqvmpkI05mjd2wK44p
utcQ7ap0y3q2WIhSmpg+4iNfXP1s8BnpZuCm3/dcl7Tr1za0i9jSox31Qe20Q4bW
QS/vIguVYP6Pg8+wwdYIL1GbJ6PKw/fsRFJ79Ubk/bhrd/HVAEIDJXDdus/7bpXA
D+/vUUC5fevg+Jnx0hOEQDsEqShmHATCH7mZfGOoVUaS8HF9qualm2bqTD1ooiXL
TeKH9ngld9g1iA5WFw0BL4IAlbOOXjp6KF040y8AxyXAtTdKJL/rlQe/dwZt6TD4
T1xEycBeVdSXFkkF3NxQTvetoZo6DBDq2Ox8/5fHILWVsbcsBygc9+D6PyDoiZXM
dVnUgrEa4dG7HClqtnFjsXfh4wfL1covN0L/xmOqKuDV1IuNj5Rq8Gf5qWwOhm4d
D2tLtru4iWxBbfVrlRtMfd1QgzX+uKAVww75PL4H2/db81bK9OTitlR+bZHDDuW8
Ezhcf2/Cuh48+U8MaV2vRK8daPPaJOorDfzntkvsjVB/cQeE+zdijnZqUnRDUquB
W92BMt6yfYzm6VqRGFelMc22cczBLrmTwTVPv50Pla87AcUjiK72Y+/zNtCBgCCc
ILF+wqbYF1SkiZ96vYiZwmZY6K2npUw1+iB6QV+rkkvsY/cqfZjjJwEYZUXdh9Gq
xon907TqaqHGGOFntjdGjQBi6buLf/YTOf4lQNc6xAzXc5hlOfclbjUG+9SlVOUw
8OYgwrj8Lzhjb8TSJBGTevPyCIan+QG9/Okp8EYmNSKdOOdtB5cUeu4JwHWTXhmi
d4z8BrkTvKwpRWKeYzVAlIsH+lb7IEI+5C+gsXOYe3Xjnl7/Cu4odOkiAt4BFnMS
o+ChzBh49YDzbJYnmWRSwvRNExTZbmpIEcTITUV8gTHnWPZfy+ZzTTw85Xds8nIH
+3GOVy0S+++skFLqBRXzAT+GQz0RHRkU1iaXWSC/90F4MSe0V6XzXgKCq2gT04Om
hL2HCtNd79KUUjw09NIRtxo6B1v8chWwfueNsrVx0jbV4iVUA+h/gvn1omDqtYSn
88JObIk2ePlqu607xP681Mc93MO0CbO+fc5hnFQ5Ff71LlRWhV/XEQuyNUILIJAQ
37TsMwOo7hjnNSiNeHJYex2onmAz+c4YvbF64RF9hr5b+CZUIVDWPtSN77Ql4Exu
wvDecce1YGFwaMyWXJ9WW3myZCGEcgxSxoGgFFIRbqAVV05xLGTEaCz5toGV4xKx
1/lK+Ntq1qMHsD3F1bAk/wE7AGXY9R66j+cG/un+6E1qhqdlo316IG1oYtuS5Amu
OvMAYf8amFe8BABXg8UbqGlTBdB5W63ze9SOlVvf+k4mEfjRcaVgZJFRlwaho4xN
jeG2mHFnhC8kQN84VvSsRD8Hxoq7ZjNkUYIVLw7pDMkjMozHjs0sUI18Bow64JAV
wgeajov/uhQtJVttr5XFneqHRXNG7fo1p/eWE1ryP91OQIeev2JjpRu8+K4e7xzy
UtRkLAGf5up5N/XpzHvc6Da6M3KFWqMs6BNzeuCDZC/8Th4XM46BT8RcXPSof8jm
rGKH3NHNe+54l3ZmniLac9oXkHIEdmISQH2AbwpHP8BWcJULidVSIiseGmyuXwBP
qrIMf0rsF2B4GR0GiHoU09N/mFNmN5SPddeVOVELhq5zgkg9x/RZVllOQStkYnet
O5ihEKRMbgpH/vIUqMIsvjv1ZPCHK4LahTreKKD0DtMxzXAgnvyRbHOFCZAjmzj+
e5gHuN0JcjY1z1pPL+AdW+3paP2K71b0AjAu+HqCA/2bvscqt2BoC6sqYRh8N8j/
/jrHAnNN9VTUXoKrqL3F/DTAvaUs8kzuJJukIxmy+bwhpdhpkMKiC9HNZaDfmWS0
IK3mX9ijbAIO+RmOPJlOVokqcwFNCAdmX+nsacL1c1Oj6D/MjlzIr0umYVyNd2ir
l2AchGWqD9VQCV1vCLH82UICLDkgTcd8B9+XRJQL/LbisZvNYX6/Z2FtZplS9KER
1H5mDz6O3mCLKjIJlN9JcIbPaQQVvs08QSXEnxn0UaFvwnPVDhmvzcIUyNHZf3+7
WktsJa3lS8TA1vdkJBAREoKqbZnFR22ASg6/4MpuL7mmEzNbTpeGlLc99oQW+ZiO
nerC/z1umPiYTErHiEtYAJgAQtQuCSnLhkIFhezKHCz004sBz5ukjqXXjroI/7wk
XqI90spIr5CkkEpY9lW3Kc2bNDhQalhJZTbu6Zok2y1WDRu1ISstvuqT5jMuw5/0
64J2UcBjfc5nmWlK/Y6v09IpR9jeQMEp64CctiHykpWd2x/YaRwj/vj74oRk0Ebe
DDc3lUkjkyBzCLSz+03nNZQX+fGft+dd3cY83MeFLJHsLKBDBxVDfEB0qKC8Es3l
Vx02H55eRV311AZkWeIyb0t50HIVZC2GmgRvk/8431lvVjl4bJG9OmGlp8YEN5MZ
YADF1Fjq8APgv62EbaLPq/4TzSK6x1MPhisXpuwxHFvsAzM7L9OGQCwRzKIHsFyi
7Pz0cN3tc9L5sNB8A23lC8jMDCWdgPPmaysKcDWMIgUPVQ+5EYgdOQLezZkH5OEq
NURdK/tmIigPWM3dUtkOi05nn7/3tRKjUto+cbjswF/988zWlX5+S7oOISXRpjF5
WOUvWTD8z27xIEqPnaeKvhJY/KRoGZI4ePyGPVUp6kHxVLodTr2rqb/iXJkzkexl
fL/Kv4es24TwShyvTCG4CorNCXwiqmj3/ndEk1P9hcE5bkQ1pPLIKKiv5ZFWP+y6
XKdlt363jq7+StWq6UjG4Aj1fuC59m1HdXvkn6e6bcc0BIkif1oQfIn/v49Wa7Dc
0NMaX5mwLbH6Zp0FVT0wVe22CZLV5MTU0BG3uLeR0fmKkT8yj5HNVkJUSVNud6h3
dkCGsN1rAkTbBORNfMkSs8e3NGEt/iHTRt7IrIgRKRxmN9VixbSbIfmNAiQc7Pu6
1vlNQIODbNaCBFlFWVhiQq33mFcIJ26we1dbVSMp2aElAnvm3WSkpvE2v+i5a7n3
jLrTe839Sw57j4WEvRmAVlUZ2dws94ECIQIWOHQe6kXOb3vLNnsT10hPXq89/kY3
B85YZNVYZmqqS/pYNKishF/BxuwtLXRtQnQkhGVOi0VlANDaK2BEVWCvrAHm4PV2
oaPYEWR1Tl/JNARrVoh9jlDUXnDvD45GWX1G4wLjHRvCwIjUt/YdB04/Pr8+1JQn
oNbOxN3OM4tXo5CUeoX0Cr7hKlNwGMWzL0WCPRla+gsDAEWwTYGs+42BpI4QyaBY
nla4kdMi2xpNvVldmiKTZPLWP8KtQXBnEPC4N2G/7kxk9q8na6Z3GR3ni/r22Kez
bW0XG27lQVAauq5fedx3uF0quKpwsa9E3yx/GpVuugJil6vsuWNyYjrQbMRRcfOa
XZfuN9HVSEaJSS93BTX4+0RW7UElup2P5nvdnsaaYSIowDF+NKrmdSP2BuAYnrac
qNSubHYgci91k/HPeto/tFU2oOsAHK483DQdBql1hLY1UJ6ZRUSQ44cvlV7HZHun
J6hmoeneaEvoH7eKBAWmFlb8/7zaog1HWPcFB3s+IMQBRtWIM7P4iuQIz/wP3bRP
9qMqC6yKCMhpV4sd0ilsVqsE09G4pn1J+Tuq3hG01M9fHr2rrFZF6VLL/JB82eOt
eUR34+TF0OatYAC4MZkL0FF8OCIFteJgyuK0FVgfjS87oxfOHPMkNYgyIbMZVHhT
Ak20QLHeFPnMDgLzeM5utRUR2CbzeAVx7djoa60zuyvobV1pgC8VRl8Cu7mqEEnb
j5vd/4TwLUyMseDQp8jNa8aNYddBuob9j81zLBCfszEdYRCd8MjEoo6jsMo1aQT9
y5Zjze0jHUtLNUNgFJzqIrw7qvI7f2NyuBxfNbAXZfj/xu7jGEKb7kGOhlYI3Xy5
YCjt7nIz62mB7Q4a5Hn/pBulANX6p8QsZfA5ETKCgNrq5ZUps2JP97zQHiOf8hob
nIGXVZWO5CjDA8NGMc86y0FV4Egi+ryWC8sgUjTAI5qH7tECHb1ayq39LEwoYvXH
puKT7asDyHwjZJEO7Tia/DxHu/kINSGEZpEsah8qKwy98S2Maxa6YY3mFY38W1tj
tpwY1O/eTVhg8jeXCsHCwNhCDCu9fuNlx5GUzKTB2IJgZfwULK0d0tuZrpnCX7TC
dXGe5rH0BPYTtwZx3SCVFwvGj84eMWSZqjL7Dlviu1xV9ur1qvw6bN9kOYtrDWnX
ymxxuVW/LuVnEvf0oApDOe6WM4KzeULNjErQ6h/HSzwCxt7rAA3wk8go2CQ4lB59
PNYX3J36Ac1KmZWvcWGisFNgMYSmNIQMe5iWDnSVBGVVe4TuaasdnSF/qeF9rjA5
mmRCwNP7N92ELJ6VQ3khHNXvQUTI1I0Ny2Hk5RglGHWUPLR5jtoPza1AVfDjXpBJ
2+ejeZdQpSeno1oP+qwFfL/Nwuuc16MXiQzHxF4GUNoAmUuHuhWP+1pfMTGALNLE
Jvtt8F6YjeYsBU9TYGaTa0/r4xfvF33rx//zSkwW1E8Qe9w9+tO28D0NLSPC/ra7
7tiyokOOH6OJf+TncGL4IX+DrXm5BC7b5rDIYImRhiwa2e4RBCX3GpQKzAIGBq0S
ps5b4gI9oLXSHh0geEiIP8vT5AOK7WDmMyWVa9Nc09RTwWzESKTfqoV6t4oSkYh0
aM5O2srq8rgxymowCXuZvpjrLLa5WW+SnyuZn1TGyjxmWY7yfTqxxNhoDCIe0XAj
sthl3mDgFsnXIFhqGNv+sASUVjD+O8xCfTkSn17I1i17SSEfGPJS7ROI4bMcuJTY
bwJLScFdrB7bws0t8pe7J0fPorBzozRI7Lqa6pgsVs/OqoC3Taqnu8WQy7fpAEts
ZgX1DW91Jy+2WYvTqCQMMnTC8DLDNjxlDdWUQntF+NiIJIDWW8YZgPPk2qCwbfBV
02e77nfve1jY/0WxcvK11x3XflIXqcqKyu6YVsStCjDxsYAL5Xza99Obk0aOR23H
6g6p0YJCbTxUTt3MtJ/e51+e/ESdZrzjfgH6nDSJyfJy8NQ3XQyNAQRazwz1uQiQ
LskjVfhI9kFHhat8gcBRfxorsmkTdPDc9FQDSKoL7+E7MBo1/mGI6VoV5pCCS2km
Z7HwWAsdNbGRg0JwnXxXBNZYEtdQIEyM9PxL2NGrviLC5uPoZGeBtbonsbBtngym
xkFFOj88vZQnxlFk4g+amu1gXPsLfIRjRRzTymEg9CjYY+/CWgo37WQV9Yi33Bvs
evD2ziDWQ0vEhwRF9uiD4oMibclstOt8Qp7mvgLNwdwHVqheAczCulHAYrVuQB+a
Ce85uT8tilxMLisuWJLbY0KhgqGuyZK3GIHKqx/rvRDDxesWj6MBB/r8PucW0fov
EsC6MxCkPhCJtQoib2layokNIDadVYPqxJeTIIlDavfZ0GTKLwVSd/1fKUXjN31e
AEia0tzrlnbJe5rhLZr8Gpnt+3soD1Ov5C2Ttopi+fCYqCI/ENWpZJNcH/GusX0X
CM9r4h0z5maXCFNuXd9LND2D/Bb9CZb5cYTpbNCslCqrK/qH7lEjl2ijTyJBqhOY
Jnfq4W6nTqEdDZj8ioO70NFd1wInJZ0DbNkzKKEqGjCRRrMHOaltPmxUzIUmZWaF
pEYWI2s/KyU4C9S18UoM+WHy8zPnoh+9o3GYB5lipjf5JG7XuN2KwIqvPii2oZ5J
Dt8z6DscuG8pgaJ4oSe4PQjq7HCXqH+33iBLSQhQo2C0v4nI22nOC5UxP/VEsZDO
NCJ4IxOnS4sJ8+iEL9GOfVSdz8McBWumMhGaZHyLGVGfACgf+H8qFr5Fdl9EilcF
EvUfpjoDKNiRlpOMB0t3JZUXq5p3bzT+rODgxyCxNfGvav0LfMmCyUb09uzXgn0m
rgec48EDddXKOtZrBC7GhUElQ9dZjQEUT8borKOM4cU7fATRiqEMF3xISOKOGDc5
F0NlRZwy3Oe3QDorEJIZa8Q4BpM+JEXLf4cWE3WoVeh9gqHSkkaYT1UTA9DPGWE6
69OUBM90ovxCkgxmEINrEbOpvxWdPhUksNsrBNhLezlqiEJ5iPdt56Oc1RT6ZM2h
BGftzFYSc4TrtXLpFEz12VMwIg+5s0Y4/rRTLJZVEysGSeTYArIBSnwaIhIKumlO
TifOaZrHjabfZ1hKhKlxiPyCO2XtuLz0r8UUJrnUtx0JQwEsHpfJdO3plybtyvbU
HalMzd3yYg7Gk/hhiXSn6wVgJYGy+wNP+w+Ef1cPWs/OeVTm+6xl2VME4O9KFvoG
o10fFycCjoTyTIbv/J7kPqH1UCn40BdbD2HGQxA18x1TJClHYWkiek7uUlZLDC2g
PhSJxGM7j2jj35joV9Rx9yO5Kw8JXGfV6yKtVjxTg1QMDmGu4X0elRVD3hAKujoZ
OZYpXzwszYTClNgcr6q9JuyNTcP3QRTyPwyYqVYSNs6VDEeUFAB/dqJH/4YUUZQt
anG6v9aQcPQPSuIRdfY/5n5jOfTSpg10O0nXxDBLBO9A3fHQajlEccxx7fQWI1if
txLlqeeicE3jmargKPyhr0W94I4eyY9V5Y6juRddq1f0XxzPqntQDI7RHh6K27EH
XECMG42VzaUOav2eIjiMnVpG2uhtStZHSQ4wdBYG3+oAkxs/oEDTTVxTSzjxTSHv
oRu9hRAHxLK1zZA0+ae3Er13IfR7rP9CbB5bnNohPsH1lHJL9L93f8EUsIrV6WPe
0Or4V4bX3H1Tv5FMZcNsX5DgleCbQPhVTqLjSYt0A+F1/9l1QSz2lSSJPgl/Pvy8
u8Mz+Ya12GpxemEe+tEkJ3mHRRPJdUSAU1bgcTRMrBlS7tDYfYYI9LMz4jnXxRoT
sgkV/f9L2cIEX0cQLW7GJg/nj+1Wgmlhyu9Mu+EIwkRoN510B6Nch2jlFxjvpreS
rRrbujOw9WPGAlfo91pCfI57lXh0rWsDYIt+gHC7j3BlcesljBTRhORhXz2WND5n
bLCilOWxF7n4tKHoptprtzzMgxg7rGEiZXx/vlVBLRHa47FcnraxEHCTRdGaSm8N
Kwu19XlX04apl6cwhGSk+NQ9k0q2IFrmsHlMsTU22FYK3YF4ZQtuqyMtwywS3yzk
9CfvKodea6Jm/NrKwW9o/eFaTqBvCmlmnXGfkyUgXuaAsXZKeNhwtFT8KFkdB9x4
pYncoKnqYCdGifpswTowAdTkXAg+vmY1WT2MIMjMGwkOhdKYp57kFXPVqRUyh6GF
JVKO/WAN8KYCFfuHlQSea/uujCge+MirDTSzvwytx7ElOpId/fQVxe1okk5U/7pm
li/o1ZwChskg92gwOnVJZPTL97kwi/ZG/9KIL3KHmizDPYDifH7q979xmvmDVO+V
9YNd+h+JoWnw4uhRzbWarB5OGU9EzwtjZ4R2o/xpJLr98xk72bavCXne1ZRbguX4
BdJvhy/P0z8qAclJitZt4M4TRrtp9yhvqfz2itFb9Ap/+Eft0U2Sa0molbN0dQYg
xLxZRlw4brzwrmjNpWTaY2pYK1+JDLjRMS3fIIEvlraTyskQSmDreXCvMLdH/os+
uQvHAarKhXmCsEJDRCK0bbVg4VLlGVamawfIrIwyrC1G2/CONC0Esjgux/0i1yPX
KhdAnQVQ/tvBTdD/GG2Eu987SfTpdshICHFhVuaZLih72Y/hY0aWsh6hv/PGEr25
EYJk/Js4EQlyUHPmOyjA55AoCGCdcXvN92HH7wTjk8jbhltTj1R8OjWaN2v2vnUu
BkIg4gUGxZfR1185p/eIctx+GBRmelSg2i8aUBQpGaZYzUFA4J4jBF4pavLnqT7k
sEKCGA/Q2IRSZufS/+LEdGO0NQmunvYQvRlc+77Apqoxgn9S5+swcRPyz6fQrmkJ
bZ4BQ3K2z5tvP+/Sj/XU0NkIgmjQ2g6pA7SVMV9mF3r2ztAYoAxmTzyTmV6NHrAE
GmQg0PmjJbJLuWUXzI9JLdSp6cAsu3O3O9yk7lcTVlcA+JG3GZf6fk4oR3r+rRns
NPmJaodVnJnDThNImKlU25WFztlMCZDIgQzE32JWgHLj4WjyaXfWcjWBhXgO0BJn
f/vA9cduZM27RuIBqCAp9qewkJeeCCu2DXgGYyJ6KNr0PbhPFTIkudAtHzOGO1bf
gPnEQDUkxiQgTHr8HQS4MqAXKNhsYtV/du3jf7cV8xH4tvyxv7coHITrsif4cmr3
uhB1HJyOQ2qMYmuDOhYi9Qv3GQFaFWZQdkGbjcLB5V5/t5yX17mNCfkieNNA21z5
roVHepPZEn1WKmu3D8vdWkxRo4xEhF0LMMG1Y3gE28GPmf5/wyiTJxuEohIAQQu4
X1a3PQg9h6CalKl+e7pm+fWcdc2EDcycwSrYjED7vtNxP8KTxRrQJM+oUowPjRuZ
A6PkVmQDoxzB1JqK8/tPL2SVDi9uA4++sgkjkP0vEYP9MWglQ3KiUmsZT1w48g7G
Wo3f/kW6E3y6n+tjs//EDJbbk9qkbjn61T0aZRRptFnAwBghPCRa0EXv0cRKUIpe
tCVkCA2HWsUEq5ooNrPVVP/IzWMhhYMDcTChA/g7FcIMyxBs4BTYWvVOl1lkjACk
1YA5M+aLOHBNLg3f1MBuZhc+Sost2HXCQ4Zz1IjRMB6e0C3WhTiiblVqnou+6MDq
Awwd9zBO12u5sTjAckwfVWyf0EeErXPlq3EWhuHNdIvJl5AOsuBDV5bDZ4I+cBYD
3PmaAx1j1LAeLSvsWdNqwnq/05pqXCBOAOs6tuBVqX/39L1yFSO6NbrWWWHG3d01
6ka2dZmaSK0nhB5F3o6/wsq6VSMN4UsEsRi0XglhnMU1CS6uJPVXugid6DFRjA4u
l+JGpz32g2/DIuwTmLtc2oeNowPKKYAE19PZlpeOdNLUCHY2GtWVHlshI30/5XpS
mf4n546AGkc1nfO1bhUWutBqOBsiPP+btaGjA05axCfD2d9N+JO3Z8vxH2MHG8j0
WPy9kd5nIsTqDk3mt1MWimHm/ZuXG2h7IjBeVX2+M/kRCtmsmYG2Eg2WZ8F8DQDa
b6PYCaJQsbjkspkcPOzVFKsGizXVjh9WBv3b7Eccg2mH3RQ3KK5tm2XGzNSbNNL+
WUTrM2Npx2jZxuOdNUDhdjfgWbaohqDpIpdnCZNTzZpfWS7punPtgbm42wV5gHjB
LNEI9v/pwsF8heA5dWOz1HqcfrCUZ18ukK7kJT3Kc3JNjhQ0A83BfWFPbkyqBTGW
8FwNz4mNNqeof5WC4fkUe5xhwUgkrA1ubDSIGQnnwo+facfsGU3Gtv5TWNgE1Vt0
RwN8qRlBo8oSUroRLdL2xmQ8CRNMVOk9LwnJI3QfJMCMceT6A35LLZ5PmWGY+vV4
ZZLbb/Pl2Hqm/73sepF7xImgopuQc2Kx3/waGaPi25/LweVuqjasXyq7X14RYR3w
kcHy5DARXa4UfmGKg+EO2jNfyniUAMnQs9mXgmE9INpGEzr+X1p/HpCz1upZ0zq3
Lqt2gX1UenMW+e1/JmJ2FgIPAPJwkMIKWuc9PZkXUM0UbLoiaxIhia8YuILIsq4q
W3HNeN+Q+mmP7SFxbHH2wuQD1OGI1jGZNXKpae+Ty0bi0e0v/6dfVJmm5nUjuf6K
r5clxLS6WHzMm3MklbU26LQyp/axRIKjUbC6u4wOvH0U5V08/eKapo7AI8YMePYL
WhWHjIgIz6JOXlrApihsAKVPB7PqzIuzpaRM+OpQdwhMpTEqxUNlNAi8w2Fe0knP
JVAw6c0hEADXcKdn3F1f6tMEV/maCDP+hHDYZzw17qu3SjJtu+A8IayNIaPpro4P
JUOCNXlaj3d0iYzKzxALC8Mfq7oV5Inwcf0dSb17GxAqLL4mXy9YBdjrXqaaRq6V
pRV+r1JBtKP0so1QpPBok+9lzBdJxfRrYtf/2rDTS2mLnMPUZ+J7dSj8sCRSBmds
SxaLAHJHClzgp1NAIaH3bENZp0XHTukRWU4HmWsBij6pFISQkIZvIlZwzAJPPIP2
XVvMSmgGmb2isVvQUSVssYHlq0DYY6Bh1tPfqZQ61o0LYJFLnIefM+oFRmFHpxPp
eZ6ys0EDxSAn0XVTHX1idAujc9mzAWoACccl61TmPoqb4Yz1COkCFAy+0b2wKoO0
2boJDuKPb5K5KTJNefIC0KvfXxm1IS9ALG/wBzIgpgtv/1Lhulthji32Czf3LYwf
KRJeWJ+Q9xwgsntjdVadF9Ox6Ju3Y3vb0VojSyDW7R594tygKD7M6C0Rk/kx8Axy
k1jGn3kDg/lqi6rLmOtaDuZRPCyAfGHmoja8fYfPhYxUoGLYSd9bK04Iw7QGOePX
800ogSAAR+V4Lk/FGMqQLnlrHYUb1KuWM3vFH1py0N1YdAInNJWDMeL+2Cn8yKjF
de2hoGQJOMH6QVxI5GhhTA0mtTrKJlf6ryMBG40/TWOb0nAXShGdQgLzHLwzmeNy
UXF5oPUjEVeHgyzcPLgAGKiuehYBVj9eKpY6l1oFFsfg435Nx3cbqljnV5TV6RiU
9yMKhBZasfMF0k6N5e1x8b5dqse69FG+dWO/38ob47MdHw3ExV7iRui61JVaH8tU
V3hao0MMK9syOtCfbm4P9CnhoRhjnJExGcyOM1IjBtS41VUPYkwZLj2/C4fkJzqp
VXX7OuSXfaKn5a6npK4WNxnHXUra17d5inRGe1ff3IR/O3bAOVdKlkGfdaVBDzsl
23loAEAgIzsiT0paiKbmvrSvpK/O9f3UmTsyD2pAl/vT4CogDQglBBoA8kW8F3hf
v9zLNms2RsS7jFvxoNX0QSE8WCGZTVUZOFHfezXK0TOBU7qUnK3HmqVHfA2eAPrU
HqM5rBUKzMfItbt6l2mgKEHmzSCcMY8uJLtf7evZ+K/2b9DUKb6ELoFPQ3d/a9W8
h5HnmTOghXr3IntiXXhgJQUk2kNP7reM/e0kP0fv3eFg0RIxllN7BIZ1C008ZM+8
EX4tJbmlN2nd3h+xolQlMFWYt//97S3mh5ru83F3azKtZ4lHug8EsDtKINunfWyE
92rpyncXEjCiT7vAG+XmNB7WixCWUu6s9bcJpjHXtP7mmxJ4r6hHekbTk8lIWc9Z
Nb3quIlNi+YkvxweX1X3de5q4JXBFLmcVlBL0QLceKDnCVGcWqCXfzOhUf1E4wH/
vMapTccFC+BgEal5hlhzuQDWz7/twLdK9GmDEeR/UgW3fNabAkx1HzevBUE70zN2
gjgcVqIf5cMduRXDciwfDps8qsRYYdLpr2PVSqC1NFDsnc/24k6U3w/uwmKxyXWn
d9SFKDOjpDWgqshX6gIR5NflkuSUJiK9+cYFtVC/MC0ExzuszMOo2FUE7jiWbc1B
95MfvkfjsxndOeK5DmbtDWwdq2Akg5hapQhpILSNKagQkp7nPj31jGr/Nf6EjcHZ
7stFdPTJWU8oVzkauPrF6hTzRTZ9xTTkbXRd8BkhcliwU8+BAtJ4pUjxT09VbK63
OFH9Fn97soWCOcH9FfkZUHvQHYX5yhH6TEhKH+weHbn8rd5GgIQcGXdKF3G2mxTi
kJHi1kcoHHDrkX73IFnynB78geG8aF9/CcwV3TPbt71yg86jPkBtXytx56hIDAxS
lwBFOH3mSxPHd0ZKWwlTJaRzvA/1UWc31VVihcqdRQH8S8jaW2gKv9yAGF6s9CSh
8v7s/QComVn3ws415q20UG32Ud7ou6BYv8j8Xm2IJDhGghpVT7i63ihARhuN7WBC
G4ndFRj1XbT4/3jOsjDxHrT0Sku/Jw1T12m7c0Qgf1XX35UG9QnL0ZagBIs8MmcF
MJvYcwfkk9M1X4wgFbpbi8X0cVnX5OenX3z/2lZxovz3KotozLQCkf+Du+OtNcC3
HkCSLu0ohm0JDBka/fqM/ayvkxBYjxOsP02avuWn9x2Tkd3+ZoUr8kTyMvrHsHdO
af5KFw90T//dTUP/D5waoR4sqiH4uQmUHX+eOFuBsB33g/xAUwSlcQav4aHLh03h
kHLvboQi6Y8jJquUuWINBHMWbOQQGpkYPbA9ybBdl2S5cxNQP3ePHRoIKgnKqjkK
FGtRm1nUz1JKi6B0zohPB2LQmRTG3DJ7ZdsbA1pY++aE2v7Xhs3DotGSG0T1waoX
vTiGxIRGO5tPFZx5IcPxWwt1rdN3Z5VkSXT9tfx3LGQkDDAI0/F9y1btdQnTQEn9
zxm5WRxP+VA7zorcC3tseQEhT4m/dRH3RuvSSm0lELALk1YpR9ef0kjAaJ8ab7Rm
lmVwM3mxGj2wFGKI3EBh9e6aiehESXwIVGfQLdQGOCau1bAFZj2ALLWlrkTT543I
ahEhM0J82f3tn+AtWoL71PuJrcOXXuLY8KR4Zzp9+iX/m1t3Ucp4CtgknWeIwyGG
lfBJaJD4m08sh9g4dxTjL3d9KMI+pC5ZMZAq7w7dbzC8G7CvopWOw6aoGL0OeUsf
o+evkgI5UexwzRdyCkEK7dQrtyg+NgkVmSXDbXd7fD881/ZJPaFGGWOProxnqE1i
4a3IZQ9jGnSDAgxPE5Ax4GoeihYV01pa9d+axPcsDZkp2sQGl+sJm0Gh5VbSBcjj
9N94izjHnQ1B/3E53k4kntwnjgvjWU0IfB32kipwZkAlwsD1OtJTbJK/zss4CKH+
GM+Enuo/i7m4lsvBwMcu0IvCVZypOdsLS1poXX6EbfhsUg3PKZXnKAsxsguwgu9I
JDCFIyuVdH0olC716P4MhBf9Pe5zUkmeb9c2vV7kaUqQo9JJb5wdOyPcgtLufUGi
ysTPR+tijJ3bSlIkh9yBRV7WvPudQABsg3WljRR6fA+HRixxRWGDr/ovyYai9yFU
xLED3/EO75GoUlyY0rxq01fWrxOZSfmt+HtRdzkw+h/+8Y0iDK9YYRq0OPnmoier
gaWfKHlLF4YmsMlSRB6QHfsXo2h8JxIZrZrR8srXzwZmth3BeOUL3USUmq7kU7jN
ZLuJGdaVcHSOFoz77KOTMIlIibqD05kjSF4h88xB/hSfWhP1mXaHZa3vkwFi+Ob3
rk1Du81gA106ZDxiGWVA735rVVhWf9eMN7jhnzWMLG6S/55ExBHYqTY5lkIQPBHh
bB6c/VzkkNbGiUdV1BvbJVGnxuSBWxjdg+UHGmLAxbMPw7uL52HM2nvVImF7lFLR
eBBGmQ/jZaeMnh1vC7GfuZqNfGwOVln3jpsF1Xi5H56u+YQtqAdDgCR4Nkpqy7wN
ZjE40YiEQ0MnF81O9+idxa8YVj71wxTcW1mazX7ZvJbbs9mNzGoyQB+7EPGyR0U8
/qWdgz7ygeNesRjUPiUn/nb18YbKbMeBLkIuph6ZHU1kB+uXI5lmTkWHnq+X64/F
h7Yfg2XHsG87wMJZryM1bB7NkFu+IYLS++s6BkzAqF1nB1ltjs84v1pW79ZR21Mo
8JS0VddtkiXmkG3KDIGHySW9zugGWhUQEnPeBRBiDOWpR3Oau/Jh/LzLB0ojOjoM
jw6RVoFnrmsljT1fbQPuQcOe5+oSuJ9ph6Jzcvk1xuUnb/r8TfVYi5HRm4RAvDY7
G9jTGRPdLZW+Y2icjZoKZntMkTqoCoLbjbno2Fit3XEi6idio4uD63xLGu8gfl7E
yYyM4W2HqmD4eVFRkgxuQqlBAfzzNo4NffgZ616UpMd+99xAlRgndk3Keh60iayK
tdTBoAh00kj7tDlMkorgJNH+JDWP+TZ+mn2JSEeVdfxXgmuFyqU6DQyU9vU8wTeB
QlR6e0nVU7yqk53a2TlTa8mClQI2WewF2wieF1tPg4OTgxJA8iLI89Vcskb/8emL
NfXFJo7Ie6C5owGBQUxDCcVzjeJAb0+ptJgv28RQ7LjDJ/jD/WAgXDFWMIQHH0jL
cWJDWY4Z+aOavrUKwKPfsHeRmS2x/9h+WaqNL+deqMlZZ3MaQJkhZJ5s2Q6/laIR
57dZ5bniLz5Hns8f+3xq7Men0AA7Mbdjz9bG0RTK6SUtqaJrbEVXnEFETWP1EGIe
fNh94Jxgw53Z4pZ4G00hzvmbl0LuklKHrn78W0WSC6MK11PEDa3jiia9GBMy7lpp
`protect END_PROTECTED
