`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g3u5X8bxYLWCrkaNQfQJfu9aJcdjL0XXefe15xcvaWNk3N6dwB7Zto6vcmtCz8F9
PX4JVn1cQ+tn7L0LBtXJkXPxTyr66HXJm4UGPsVbtTAkfhrQCV+FROt+hiG47VuQ
X8TUdFZLxS/JwMWNacX9N9Qxk68hU5aqxTBwN/L6QeqfW4xzVniUPeORQq7v5D6y
tMHyEeaG1l9drbSCyqkLow1ILz5BBHy3ygIRN7bfDtyMN+xngng5G7HIRRwfnpyJ
HbP/ekeifA8C2nvsGV6d1d9XWHhuT5E6alnxYLn0sclqan1yVC3195rknRSmuLbs
d6Pcdr7AqMZ3yeSimslL1XrSVBDbsZmuZWd1ZKY08vcoo6s6FxIbiHmgCxOZxOLS
wHYWsYkHxjewscSonf/kvm3kgN8llUmBKAIxpqnFD2o8yb6BDV+bwSSojVLobH8l
h7DiIU1bzE1W22+rNZQ1dejcOGoyeHMS52B3aDN1+toXoEE+eVsOGvivy1fWjsg7
ZhvTQNGmLFnQYR7vCp+FE5MYu0Wdt7xt0x47R3iQp8fMbKkZ749HsW7ih1TGXPR3
ihh0qQ8iKY/abcra3t+9EKNyna3qxZ3sdO4E+6PaIxz+/2xxA3PtLYQe8SG990OT
IFU2QPHZ96arzU2yvsUFvfJOYYZF6obVMYbD066iyWIS0edG1Fr5RVCtH/iUYHtL
KYJC6+M1kgYelcHF9NKhUUKWfL6JI1QfexSqhvpej/Mo8PrTd6jhzyL7s8wip0OU
FSfRal1tFQFNScWAamv7+C5/CjwOTzUHa+GJdMppvx80Rnk9mcOjUU5FWdmO9nbj
3E+Oo/AjWowh08F1jgJSQwTKYa04iizCjrtdDT00LmcAAfLcNNA6TNBc7pP9dUS0
eWXPg/xKBK/HNHoUq3EillNWb1jpFBtnIaTwlW3tq45u/rs5+0DJ1oHggthOpP5z
xfiwN3r+CQ8017jKT4opbUmUi+8/kQozGoXlVhCQccJSHSxr6LneQm5jEADoou6h
Vr2DYcYhWsOdyz2AdWuLdk03xYIAji68oL2jCnIfn1cMyWFA6D8jlw5tfhBopQJS
8M8BMC931kXnspX7YeY+uuCb1bmgDalcVfcvCHjoOL8rt8Ej5bxM0V4k+qdEvpWY
dmEpJTJaEmNRWK1r3Iz8KQ89IwK/UO4ByfLIhQiLC8j3dTptMsHXT9W071JA5Zbn
ByQ02fSR0fXTbKde9DgqkE92Yj30yfndx2ZVREXsYBiF1D+dYTFgCeFU5/I89Osx
fUl5TkLPkkd9+UMpwgqfCcgecorzwjsHn0CBcxe0EqVod8GfMsD7uWMWBXqlI3dA
XjtHYGC3yTrPm5K9cIj5p8bEEDqEG+FNbNpFfpslmZwmSt9nfV+df6oPGjF4ayXU
Qgu+OVuwdR9HG2R86xmScwdjMYZbzdWdiid05vdi+r8+MppSPcABJcbl9T7U1VGe
SGvicWGKWw6QaRymI3XfDXPj2MRB6a9FjSQKCfHnXT9g78wGkQadYhkeO5AAQ9Ik
WRqtMFCIf+zwqlEeQDqcqVgPe19m04aWwpQjKKMqFd9DFMZ2qzdhtmd0dA8QLzOu
J7LUZvhdz4zVLQUx5cOQ6seGVKgPsSVUtxsdnQ/y6hyNlIovP+dM0GvcggM8GxsN
V8JbfWkG5rLBZYsuTZ7IPUAwcCRqZvZa+7PAcRKKZkCgifjP4SzxCWO0ctZ/JZHo
F3OO19R2/CT1iy6zhTCou780V2jq4UgDmoT5h7/oLVM0JKFiQy6jdBE2enMs4saI
FWlmOz8CF3IeNU9l+7BTvsaWiFqgQkxHUr07WTPkGIoMbjUnP+75jQw5j/v/t5BJ
uKREZHaLPNTFzhGAvdkmYu9/kYAAKK7d5t8XZJk6lMVHSE4Ha8PVW2McMM5Ucggk
dJWLIBZ8Rct1J4obAfg5uUMSxPxzvyEbdc3IJSnCaMsCGf9nu+B+itgnULJvfl06
gqJxful+G/etPn34d58myuK8IL5NdQY+oRMVvv67BgCdTaRzzXZe5plPVuwN3oHv
atXPO4cQDQQznVZDDd8pNQrtWn23IR9t4gCw93Ya835eg6Fc4GzzmYoGhveA1GNO
Kqt+beyH/iDdg/AifF30CyLuoeXNdsozkqtyGjzK9rsxLOfAjgE41JVe2LZigDS0
2F/T0rCMetaN2rngaAMV/pB9QqKyV0mZV+A7zJaJrzsPxvjGnAPbTv44q/adFGOR
qj099x1a+mfiDq9rZU6h3SzgGDarmvt++/Wdb8ruqco/Wt5Xl4iv+/6TJuceP9Z4
NkdDofed0dXBKceicUW4mBNY3pnNLH7ZxcjtpnGYENqQF3+01ejx1JIqDa6A4bW9
F6CEsd711Lvs3zsVB20iiAhre/4yZcLN5IsowEYbmTKsOnN8/Y8sTKXQNewKAOQg
tMy0xNYjY9LPnOuKWFhPv75gNNXCww2eQjev5F+mepsEmZ3He66PJKsvVYTXxMFs
28MRJ+pUf7LVCInOezmLo/UnXCsXgHyrtxYWWro2TqNhqmGPW6fD/1BDN03bBkKb
xW5L/1dz9A5N9+51kby/jSHl+TTrKEeHkJeJsLq47PkiSPPTyGvMdyZXNS7r6bc2
hdrDJwm0OKvDGjHvBt/PFgsJVoZzpiGpI19FZYfxz2GC9wA4hJku7owq0WLwaVXN
AaLLDwvAbjc/Up2hJTzl2RHurCHlhe8hy66yYFlOQIHoO1hJ/I5Smyt59ziXudUG
Wr5QIHULQLQP0I34BmJ2EqH9FP9MC1yqyuxa9tBBfU69JbPGPYoupjzk27Yk/RQI
3RQk78GmJOoCedwApvnWQZk0ZpouhtzMlRA9HIf45F1OcFrWbbQwPCkykKA8zoer
yXHNEfgj4qjzY34bBO3ByJvYywRX/IXVhK3SUxXd0x6/DTBACYwh190eaKvfyEdr
5lTqXlgfJ5meRuab1KEyxQ+rQ/jH76AntQcFXgeinZjjvltoqJkfNR984nSlCkOb
2bbHWQm0RnYAD32LLDCS9ydwpSzMcOAo/xkyK5uR2s97zc1+9gCHd9vEBDbALlJJ
Fv8sm46uFGaDsZ2hNYYzfZul4QG6etIAKPlTI4/el/Q3t295pk2zKw8qVLpWdpXg
wlKZR+1kEmxwGj5C215Q2DeaiW41XAUk6wkoBx1/bcgt8F2RK+bqf6xWoGdVaalO
SfZaQpnOEa0rZW8qPVU1852g0LTZln88R8N71N37w1eCFHYejkCpdpwAJVCUQkKH
gITIZVtvR+bN4tVKP1u0Wy8G/59z7vkZJwVEmEjxvej7BmalCrqEHcem57Vb/AhH
tduA640UcTR41JhXhxCxwkCWvk75WLDFU8c2+RU8X5c9bWEHIYnkBA4D7cnl3CEL
jc84c0571UNpLkq2p2OreUBkvLDogzap95uX7zJ1SL4GTe05kCp2FPb5fZcMReOH
pO6ttCrC4GzrdzWK36jlIDYd80E1QFQCilI1ptUSTw0bAxR5W0bZ/SKHbVEmBOGt
wIiA8f69Jbs3AifyAXrJ4WPf12tiO8MXh4mnehuX4wEMtAklPwPGU8RKFNWj5Xu1
mfhQ1UUpXxOj0pj9QXftwxUNAR2gq5v21U5TXeoeIkrucmYbTOqUBHgYSCwwfIWN
C/Uek7aqXEJB3qYGYsCWjYkdE+IuFtGe88Wf5rCKZInlMSSABQZVoFlUnyKnCx5G
CFDTd34hiQPJLF1PSVXrGLQIWDxsAHMoykQY1SseXrQP7hNmqDn0sTOJFgXLAjaJ
wQQxqNU67lVr69Um/YkObOHIMS6JQAeqET1b8HMV6Lbx05/YsxkoZcf/rCDXctki
JvU/qm23kZFBzCa+/1hI+n/SK6s0kMjKpZ6k92IxUVZzFdqP3XOMXZzYzOBfJPiB
a9yboJyMMh5777soRjzeT5SwU1Cc6g7hE5Gj5aTxh+adI1qpvVQNcoV5KDZKgTbT
LyyM/mB9LPJSuKlaRSJBtCe+DSqvmxVK7ISYYMKp6iRUJuSqk1N4fZSj9NbNNpai
HTAqQBB97L1qeadeVKnkKbU5N5GIzCPHNPLEPyULOK1exwJnTCuYgssKZgFXVN/F
Xa8xIhyBq2fKAUyVPZoITLqfrSYXmq9Zh2uwzKFEsH0HQ0TAku5ysSzGgZLaeiSR
C42Yyq3TyirZxVUjOSDADcy6Rg0+i5nXiZMtK/iTUESksQFDYYyPn6jAfNUBbSWB
NL3tkmFIW086rytxnA6TRKMdcwwKxDJGdTpbQVm42zWH3zrxgPZYIaztdVqZ57fc
xLC+S4FSUVk8Y3vb3e1jLKYrWBJ2Mg9P6E5k08YBTmup6tZ2aYtXft89HPQdo6zu
dn4l0DMvJvsiWWvblvbQa0zBVwpiCxUS3cSlbqmF/OOiyVWpgJTRvk+U/QWloF0p
WGzWVhKHGDFgD0RuLTIQSHIXwvnguEflT1ZGoiItK9YBgwkSLwAzD3J9RVbZRMvH
OIx2SeBOv/VMogcY+ENI3CRsZRMKch2UDJENh/ZpjNnssyoeqHC07nLuVu3TJ+9j
`protect END_PROTECTED
