`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/WoBLP9Ipj/ZBVUmx7fJlWO5DnBzTYT2LCu7NTc11YOGIvYiSUP/7jrrZrBZI+O4
tGbHhmRWirH09x51rRUxuzQ2NhDqq8W+hkyiPPgQkPBiCeISx1h5DqPMr09oRupt
rNZBl1J5+T/QXaxmFPBjVbBgcY+J/Q68Q8u7HRHE3fre/l4iavuUIIHghGxvX7d2
KO6vYuK3e66C5RKhJS1kAVSWflk7kxXh1vcgUWRhz99szm/X15tfZbhuUS2k1v5U
aqUmqVwzG3FTIlvU+NDpqyp5B6EQ/MtDb18191gl2dOUmR0n0VQqVGxyrcDHtXz8
Vs2fTcjTEs+eP3T92BKB/9NgJeeHQxW7XZRDvgYfGPjGUOhJFQqRLPhc013zWY7o
L67dnG3yYz+RmYCLn3Ue9owwrcAyu2Ke3bj13bAj6AXqr0PiNQaUQ8qoT3rUSZSs
NrH3oKyCzQpunjAZI0UcPPSMC6rE+oDIw1XBmPyxWCgUl9gmDj3FMEO3SumYL/KC
HG/btYnhSDpKSw8gezVyCTCxlVmpbluBvRKwcW9X7090ILGqauGjUVNoDS+wayTn
iR6os72NyjKz5sYlqzSwHQ2pt0imcJrqo8ulE4C+Aho17ZOu5ADXxkWnHw9qGOhk
vP+H/FppQwQmaLgp4+IpLM9JhqWvJfJvLnt2J6U7bhU7ihxzcLzKIt9qZtlzgz3k
dg/8Eit72Xldi95JjkCkAF+PIqdFM3BrzKCf9dowaT4gGX5v9zR8Gw6aaocraOy3
BzAKzMOJE9ixhG3E0UQg5yKmlHEJIs+rMt875xBHcVCwD966hAoLvgo3WAOXKEt1
XhJiDOypy9/Apn7Q7LzyZWarSs3vLqEUyPSJsgoMUpcgbYmC/k07yXArr96XDwBh
/ZJOIsRC9OUkwdsPXad1hQ==
`protect END_PROTECTED
