`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBg6cYw5q54QFyhsS+L209qb+0dLtp+QyIJmzzXEKM4+EAo8idW54ukLC6+W5HBf
04DQuN/PTXqP3p7HLQtjFYWhoX+Yxspw0sqSWWoJvsLAX8d1qb1QVegzsB7HoTQ6
N7Fu1P9uHk+jO21+ytF5x4XylKTuO4EKLBEzytcevWJp0oSIiqgC5rVSyKGHFfhg
ZtbBAGtjA0NIPuJo5UKh1FzRsFntZvSMc282pkR4qY6voduG0fUiVoD3Va0dxEIu
+00e5AsZZ+mBUS/MEkZxPPFVY18rmxz83uiU+JLOlo3tFwlcgh27+PIoQvEGGGuU
5Ve5Sy1O96bELmyILa0LBwvWK08ylDHL0KpVIcdHt0H3NO3S4c25Fjl0nsBo0TQJ
qVtVz+/RbejVSDl7BIGkoTzH1qByGhmghJ5eKzXgtxkPDq3XFTze/MyONfqxaNjB
HsW+jtWorQ+9mo/57CAHRQEO1rf5rk9tbk6tY6NRS6EPDUl/zscCPmuNcChS5Ofq
HDFYfxqjr0k3L4I7HiNeZUOCqECKyvT0nVwts/QUaMuh8CkGwAFd4ZlWfYfngGap
`protect END_PROTECTED
