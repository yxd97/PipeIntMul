`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zl9F4WwQ9sXsoFbpJbwYkpwOZHCiMJZqCziAUfed9XJhENIxygJ+ifxgakMGIZw+
hyTeNlp5wbVgM20tF+u997CHs5fKJGmQHquumXg9oVIC2DkisMiHHy4+Cd9m9cKU
3m8dg6/6MkZrhajExV6OnSR3KXpUdjDODsnytOjA2SNzTPdjgWwhVTyq6MsLR7qX
hrMq2S+YdKmO46Wnx9d56eB1KqMhhZZAlxPaFsd3WMn2raQzhCDQwBYwIb+tWT9w
u9bYyx9mb+tGqqOFp4mkGWHvHPk1mz9ApZJ+5pFa7yWqq0kWt7IA+OgRdBcOjJzB
39eHsBT6Vt4qAsSsrgsCD+vxpIThakllJgX+9vckF0VcTR+t2nDtpSFWwPOdFA3f
8d6tH5aeOl5/a0AJfNOIfD4Z8QJOhKrTiUja6B/7+hTPKK4toH+1MB4fPe9Ncdr0
JNnJOQ9R+r3SUnuGLd2NBJU6U6DASnD2UxBAdB8MxiUnjMKDIoP0KCZPjedzOs7+
jWvNnp4SEcqIYMTa8G76YSlwXphYtzjlnDaQ3cp0NZGAe36A34dgUfIxi0wq5ctQ
uA07GLYriv5tK3BWu0Jy0k5gZyHxNseYKzrX/DPmzD4LkEs0aZK08j/79lQvX0rr
MvVNPHpuidffXmc/JbIHoh723Qtg5C5in+1UJpenY8wmXEzTlhOcdpUNBJqJFfOa
p2wuMDJxXaAmoCXjVsRO5gcMwcFgJ/tUULINS1FRpkpvNKJ9wfTn34QquXMCoE9f
pgVBmeKwpCwoQyDYjnbUdA6kgeIUCLCgd5zXXcy4PqFqTCeRefJqpD5nu5JPMG2L
tBkua7qoL6Jx0uVC/Rk5j99eBMNIsp/M0dijELFEW3XTkcJwsxMu8K914lQhGBvw
fWAWu2tvl5kmbSAbc/kJLzXFk5O+QCMLBN0xY9h+qoethpRwWqnfGaC4aIsyjIzD
SZAJNacpP7iLLgPgl5zaNv/NRiXs0zpzxIamDslTBhPi2A8UZCKiK1BPJf6N6+6D
ER2T5I4zPpKPVq4GshbuegGofbvbf3XgciOGztSsWMSSvcT3msxIz4YtF3+9+EWn
o6M6RSyRpVrFz61Y6TKmiuNdaKPPJB7gc+sztOt+bwEtQp2XD6dxgzaN+BkZll5n
jw5RoJocCQbLT5fxDLxhXa0wSuXvyMpuFATS65yQt4mH+yBJZx7sboKR3NKMOwFE
wZBgApzvfdlliQcFgr7tRhSgR5hV+i5htzgb/rtQsnsn33zo2YDrHjw4DNmATOaQ
hMLt0WEC5HfFT7BzQLMrMAkZOS2f7uPQOiu/AuS9CzhzQeWGuOggqa9Pb+fDJiWD
wHn9ojY0Y4GGZrqXWapwcXQcjxB2KUr566YuhWH87btGdGQ23ggusM2QFkHnncKV
O24y+TIYmMAen0kOvv9V5IiWkMNsMPxuLNFXswG4HwjE0bztvqUBIsdgdwLpr+Sq
OZDMfkaD8mRnWmtczhes0OxgekFtJhUXi7LOsydUmAWJ9yDhIBy4MX86cjAhdTIE
yF7TKrXcAbJ8gxr8NjPWw7UM/Gpe5rmzN2UCISs0EyUDSc8dpRUwYcX58gaD0Zec
5MomD/rFWa1xT5AA82IDjyzGDwsoRWtuxasSUD2FIBdnpe8OzF/sdeDQAIX7I0mD
LiUsjLRNbhPU6I9Vw/EE+qks5qA0RQ1KHQ4qE+eSKfg/J/3hkL+3qgTaWeCaIqZW
OyX97kSt3LS57wkhsnO1u1NkzcK2F3/pPSmQ00jIPnB6xpFPoCF1PhiPGkgyp1xH
vDOwHWf1spRgZsAEDsFRAQAZXj0XtDQqzplLp3HucQBaW5Mt6zpvUhBul4ByYUkp
dzAfd4RvmAIj2APo8OFZprKkLIYUmv3Zz1PLsXKqGtmeAaf09ijm+Gk2h4t56wDD
ZnAPMoLlnljmGusrsBDZWv0FrpTqZaj6ptaMCqCrg/WHVz2e9rCTxvvGpEmYClM9
qtWNfHLMJKuIHKRnXUSVKS/2WTYx3MJSnL3VwYbOWf1RcRp4QOd9Ko7JsfDyPk6X
nEHAPt59hmbxOw0Bqbab1p7etNvbNFki2vujLxAeW3lh06uabLvmimm7Vej5P9ZY
71tdCOApTq4C/Wmm2Ow2gwkvh9JE5aeIhNcPoS59S1W1xDbnWsQVf4O+2vlxF3yp
zsYjmNuF4RQYKHOaZKrpuD6jvt+Ay9u15bcp6JJXpvhF1l20IKeN+VmbDhAJipF5
KOz12un+TDThmEhuAnVm8qSJRH2ocF2P5z5axVkZ6LAh8oNccY42OxgOh4Gs2fN3
a3pK5gQOAbsxVK9f/bzecZWbGn7VR2rfrk8lRkqdN89QoiwbCGV1SLWyVWKlckeY
bqPZAXXmylCXjD9W8ah0tV+evI7bbRpigfh2RJBsR6byY+gn1a59mDWSHkiv3hKU
u4YncIK+aN1iISLB9jD/5OzC07JMweK7hkOIvbnMrCePBL2aq1yklYSFpfttFpKz
P1l1zskKRl2xepKgDB+Kgzot2JD/frbfU+hGJKPRyJsv1BRP7sKQ4oNDWPV+nEr5
jm0I3hZVIkFxRLND7EgttWIVKlVLXKxr9ZORPAa9k7+EBKwHnowvmbnm7NarGsMI
F/srckayni/9lDw6sFaW6ZMrS10SVckhOSZeowywfYyLNnuSA3HaN3fXtpsWkm11
B5iiX0QqSdwXGBo8InXhg5/bDtvfQHF64gcQ5lIY99dSEaeU/Ed9aSpc56BPiVjB
rpQfj+/Y52Oud0ch7ud0li/Il6FvHaJGJBegsLLIU8mOY0kiKR6HRh5NNqCgiEtf
q4gC2X70QgmviNxHyejnkzXPxQR8T5VhaZyO0bgr9PwHu3ZfUbiZCLW5MAdMJzZB
OaDeyKtndkfXOd1FEjZRpXDLKmCdTdrHWEpXItJwb3acJ2b9MVhplZSSyzNdq1EV
QFnMaQBSTmOZ6LXJ/3z1sPkykB0Nj2i0a3thEWFEo7FJbkYthW8k8fLwPEiKNnRG
35Ky7wsWR81RCMTcMFg0YhpYA+xOOBpL2z0rkayWxfA9zs+3d5qGm2PY/VnI7/8f
uXRR3zkscpHxo7slaTpaj2t10LspoTjlb0dsm+fqgoTHCN6ciHs95/uduRDTprkD
AvMA03I+xtYXwy2F40WvCvKe5RqzVxfXVvqPihngK1YAjvHHf4E5AgLLFQvucymf
HzpvV6hsFxOp60deWaGdYpQnohrKnWhgPPttUYktcoyQoKYRdE4VUwjYhxh9iuaM
7Bi0I1ZLWipzBoM7zhXQMoGqKBUOPMi85iq+YEw8FyJqI4e6kpNTZ7XPzxISUOzM
T6u1r5XRdD63o2no4poIboBiMG0k95re3CONI3IAqtQt2pOiWLjYH6diPSHaIZcr
1KzYJJhJPPuqS+CTY77u1PlSlrnXBarZ9tdoBzBkUXNqvLc4ps1Dm7FobbS0M+4L
9dVPH6DxBDd9NgiL7VtSi+zFk8UOHk+wfqRHU72ee4S9e3/Hhg8uUK3rnzFrEM8K
Xp+c+sTGYwBejHXbkW9AC19LLjTpcbf1eVSMAk/rXnkZGstam375dL2djv7QS//X
ir41mkmWSV0qa8IR5gYOB/nGXOlMozWMByMczw65XeJX82LEb246bR54B7R31Did
KkgqA2jgDivlkF9cGn9rvsOSqVmkoe6qRHf1NYqIHze0hl5Jl6he5CyG2E6F5JyH
ccFaHeQZ9n1yszySOKtwbhaKD+O6FVxqmcrRIQZ9ZRH/Ax6EJOd2/z/p8QStif/q
u57Aiyr/pAmRB7zOQEib32KV+pieNKF+TmdNC/9zUWPn6iGyjDP9vRyae39B7s6c
n7ecgXu6z1hENAvM7pY40k4sIg+qb7tiVQeTarfOlBprbhz4zmmcSJAET5oLgwKD
JvSEjQEE+OrmCyCc1ErhCa7z1BWuRVVhnPXw733V1VXH3JF00pt/TEtFSczW8SSf
0xH8AaxMP/CWr/H6cHaI3m7CWoGE0TTRWdVdP73PREuC2CVsqsgZDQqUs7IOCyfv
8q0XGugEi2vRQE+/Fx66CuaMca+a/fnEDetvsdViztnplo8OB/yWVErhQjY3qOCf
ym0kiTez/kX/OB4poli+7M6vBx3JRO8OPDo8Jv6qIGaLqQGui7Vl9mo9qoFD6QAl
9LW67S2Tar9/iSDgpho7+3bHQijCK9Xe2QXO8Ik4Y4LjC6DFI6aV1D8scdsH71eU
58fj7onLUQzESBE7Z0UAGci6weRnsQV4ccct+UMoqtVdf+Hetiwm5em2dBFOiw4u
WZX1m+lkrXRqU34LAG6OPzAC+ysbJQkKVOi1vxatfXtTFf33S7nmYMMFIV48+YH3
AiMetlTOq3rkA3EVmZVeaIxds2cSkvloqjscvQTJSKpGfu7xJ8tzMvoo7qVdfEDB
MdO6jMaP8SRbugMy/xfnzRhrRyil5GM38t3L3HpvudcHvj4DuM4lKrGJoy8uWAzm
MeEuusDlVjD1/XV03Z2tZ4s3OiyVosT8q6cObbKJg/YwKDuOof7IIH1Lw68ymkjI
VAZtwCQXG/jXaMN99ajDAa1KNy4CVlVIP0AnxWTwipEKBpSPNIKq5KbBad0R0QmW
5BnRaJcjZjs7CiYnciF8kkfD3onSH9SOZzM97Ja67dxWsneRJYF+dTXdjI1MRY5Z
vjyxjuPazqCWqk4K3RL6439LHYyRItymJGiuiCEIC8SIf4Wk5NiN65dVJL7LzYGs
IREO+ksqmVgiDovBHCNRT6e9QOsYd0xHm3p3zeJ12xrdNvyqjXT3AQbSx4zDg/Ny
PN85d4cKkefh6LgS8xdT40+kCUzHakoug49fifSkIT/1p0XwjaHFa1VluGXl4Ws6
S6kinVSd03r7L5BU9QGJPr6TtTlIOOfZ34pDGSph/CzfRaf0y8q58mkx2XvsHrVN
HYkEhjQxzD/vDrWD/uSgTHCqS9qCA/tt3lpKgSx7y48lSER2m5vxj1UkTC+AYsYa
2Y/eBq3gQQCzH5G1fIFcIyjNiUJEjeZ1kcPsWEqK1sBwcpT6C8n+OF03AhBkId3R
lqdJwYGM2OBS/jcAbP1JVIxEK31jkp0CCg0h18frWpJekM2jb3EanzIYSkvYaqvp
F5An8HOkQIubRlxuZlR7A503fDirMbQ5wJvC44fXAA/uR0UAX07zuRyxF31yqxRM
Y0M5zR4qaSoD+4ggaij+IEwYkevArZ/M8GA34lJTY+57tIzEmGpliUYz8MhBkuFk
LTy/F9Q+Rn+LtjG6/FkQPdA9PyKnwrvxBrpkZfc2GaNoUxjg+KP2mZbDWbI6SLpE
rQMYA44RpG9dCpL6HEdgKF2tEbb3Y3hVja0/8jADDSACfW+TgKvwEC+hlIETaowz
Mq4IxMZCEEX9v2kT/WftRtI3cM09VCOPyX1c8HFVzJeoQHnPPsxxkA2uCLW2SBeb
ElRyGMJW6APsTWFgC5i7XSUI206VK6a1fE+L5+qdvdL4WIJc66MKqDQgvMsYTN6w
T2WThW+Di3heqn4j0tmXZtm8k7r3rlJNZMvCR0xufZnHtYR+J02QiB6NjMpnIeJ8
jKmXpyF20Y6lJq1j+UagQY0lPJCby1snhFNixCwjilgRY7eZeGEglzpW18sGsZ4M
BjHxq52lIsE/JRHG+WizQ0IsVyVWRPiiZwEYhEh2Zn3pM+I5KDpdDxNly5psIqOv
z/a0yRrHASjK54eLpPPqu0NKuQ3i0KU5NrfijdpZLkH8y7eHOgP8SWoQoZiE+Dj7
t+TDDDWXYcrWCSTqEygxPSpP501Z9pPQDB1ghXlH/Me+qUGZCbqzOH+4bDkfldog
F1C3pxqDd1l8YTqRNZ0dw85Vo3B+HXrkvfG2a9C6VNCk86e4/Cq15iYzU/3a6b4E
vgnmliQvbMD6NWviI8JJktZD3Z8A4EO1jKe/3cDONhSxfdZ9lDQUOWkNRxzYZI5c
KOB202BomcSf3uG+cb95BeFDwJ7iUOr/XWWE8Fexn3CsqmjXB/GRmxZb69v8f5Fi
H0wDPJBFc1FWrqai56No9cuOtb7F3bRblabmItR+WXSJfTpRQAj3/1GdWv/BB306
aJ97+f9xiXCojZaEmVhYVPef8XxauEKhor1J/T5q7JJDTSBZ2+x5S1KtN7pkpOW6
WSHJQVhgPQOYwrN1xcgihUV+plu5kAcWsTvAQjvL7XBto0qF75q+AOeDNkiKBycR
SlhyGDfHeetr57/0wyrv50ZshV2xOA9LOPtCOabE8ajMM8N49Ko3dEABbUn+oitZ
OmlB2iylDByk69fO50farINxiPssUcPu9hVrgUSkHeNs1fdncRR3FknSahmZuT0F
guoADk7WTa2OxJ9hiWLewqc/gGjYmkTlJjITuEc7/h743RNlHSZTG/nR2vDLpr2Q
nc9+o11ZzPsIEJQsTSiZTZiw4FFfgQbudfNzIJSRx9GPk/rblMo2lcs9BV6WVAYy
huSJ6zBJ4t20KEaHzK8eWo7d+DQjZVXcq3BpHJEXfgCyo6kt+9g4h+nCE0fGI5k1
s8QxhjcM1CBjwednhZZlzw1ki7xwUbI4zoaeGTDNaRthH5VuRQhfVOvtsOvZ9Tte
z+sErAwYM2rgDMTKSGSS/tZs3BP/UvQkg1D5+jC7onvvEa5YcfsbCe3jbZJu/gfd
862hrhoOfenFJRpTTMzroDrxRyI9N3FWAkzr8twGVn8VeLXeL7Ka5kVdFs66ejpF
5+38lQKFKBsO5vf2zVF4AnQD7gPjLnu1/CjGnCIH6FEO3HMl6LCFKejvqMgObAYa
ten7t+1eWj27KekqPVmUm7JTwaWWeD9nx8B5bblVP5Id4hRcgww+KblTQp8f6UVW
iBnp9RzsP69b3sdGUxRfnY3f7TXjueOYGm/sm6PPbQ4udu7xSGEMTTNSMAHzK6vw
PpClGImh4vdjZrbVMcMBBKqWFdCmL0aRx7+Hve9WVPYjKZV5NIkeohr/UcMlDAfY
lclYcO2rKtBfwkn6W5Dc5ddsP+bnhaUPasW8u8+b+H7GB6+5r+OWWJmkJq5ZtdqU
qzw0+3Cf/BApizfdQW2fn/NJg5OoSfBPbbP/wGB+WRp+14yfew7BFx9h8YmIQHNn
m1JG7bUmLH8YfBRULz3IQV5QQPeETIsLs6NdeXHY+ix9ilDPOLQk8rmeLEvCps9a
z1+DT99g8lc4JSrnkiyE5N5Qa5pUmfdKRegPjYl3RGLUeCo7TomxIfSP83y8OSZV
EpvGOzZ63v2l6jHwgKvlyZR1B1cfoesE0tD6abmWzW5lrcUS9SB1y0EfPlyEm8PD
bnJURN8YjLyjETiQU7+SgMlR9NjG+GECC66GZlVPXdJkkTINL36dvQ4slP62muVy
i+OUzudOGIiSjxSumNSzPqv63Kbjk81R5zWCbhjZVP1x3q2/Zw5t/6wlvGqxSkA2
Ayaeg+DEzEuhtEamcNncpiI2AFDEjCr0ZMr89q6bifBLP7vfcVtip9RSTq4uOtYg
Yg5A7oeB7YUvd7pMeMczrJ385WM8kOPpZMnEGMpupiAhUw66PKmORn1SRC7vBIDg
cbIVMAWG8MyEZ51114360PTPUSG3r26NvmyVI7ZvrIHQIqOm+0aE8ctQfTw2B0eu
3hLub4CU+sJvzif8aNewuVyW/7/KFdPQukmh6UE5OBdTW7LuSQz76oMlhsXWcFTN
aJhbMlrnqgovAzb+TVw1D89KPtnHNzjAmfuoaXPicV6+NFKR+YW+P2FL7PXszpL6
UJEfEH6pTt+Cfnc6YCNzIfAC8gaHMDf3VU4cvdDuePt1TVEoLOIsurExbYtHtXkp
RjRmI03yYP/80/f2WrC4W9VJ46XLRDJM6tyfJFlgUAePoEtylqSxfcN89SsTSZw+
XpZtmeWOBkQznQcskCm+e2E30Vn6g/R8ADXM0dJWLtlrXZGSUSpv9ag5W9fGHXDo
iE4wSeu4UqSONAO13g/LGUD8pY93da1L5OyDTFQLx9ckFejURxgFkj6EM7xa/mnw
MiQtzBaAO1wXs+4budPXjHNzeMPpQGluRsE76jtkH0Kh6aADrXr2fW7PN0Dud2IN
FWiBcI2d8Zk5wtYZ2t7YMkhWbRQzScXCh2P2eSVCdW/gqeKx1f6vXAwcE2ZZwPP3
sl1hNRTEVd4n2Mu3yaRNrapCpoohU5MXURLGTMuORpx/rKnIi4lTFMZtsZjDnmGw
HIbYECnKqetXIml4kcLjcIMy25MDgVGubW6lT0dQ4F+ld3GQpz8kpHIMHiZb7Z0x
qCLTEY6fFoUpzHHWTM/m1/rsnqRE9i4KPHrb0dvKT8Z7PDUOdUhm4bvCum72r46t
fUd+L2M0jkfknEH6z5tORq6B+YeOB1sPP46YJyGJ5EhhDbs8Byabjs7ieUAoDIF0
Gck7xxK0FrEvwijVA0EjHlhyMhgsTVEmjX4/mz34QKUb/WQGcbrEQRQFt4X2KM97
ImPGCeiDoeL083f7k7EL6se0tcJSt4q0WXP+bJ5mhhXGcs55qttc6L24nW8Y/ZCy
MbAntzRtGOaY+YDWOI5fSGuIq9kO8nd16IVRzbZRvCOBAfRaxnhXyBu7niJR3Ojw
uT4lvpj+y2gBLfhfkm4L3ILG4KZVNLfZXDt8PfDa5bbt5geW8LWh2vLtjByC6Ksg
BnBd5cAK1yTL9isz1Up3RvFWLeEt3MzPW/JYn6onrFBTN+g+/WqKrmsjo5Dmh9AI
riHXruRunrr19JsLRU7zWCOpdV2hEUtOl59sZx3HiyevuRwZ+temhhu9K1gstcVR
iONrkAivJPZ5CU2cEnjqt0B+RzLb/P3FqU5tmZOnMd5KeYQGkbAx/SihevNbE9d7
ypgc6GPF9/sW6/1UsMA2z/R2/nZuYl+j87To0RxINav2ghaVH4LiKp4OJIt2BWDo
z9p8Yqwc5ZJBvwuLaLFZVOIurOVbUwtyNepj5TJ1+jpz7gfKZRoUdN+dxR5wooAB
QMP57NkbzsekClJxIcN7scPu6S6DQSuFHThS7iRnRU+LUrGBgJ3CbOTPybjMemqE
sUVDvBNleFXrOcYa2in9umvsbZtgttkWCRCAeG5VpjgQgLRube3v89u0sfjgY8Rp
2jpsxh+BVRmX46PtrRAExaKaESDK4jNgnSNMsknwxkvlQZ/Lk5ENTJQlQ3ZAF12n
KO2m5cS9+mZBjTmlTBVZ2OjuUCIokClzYJVgmg8kXV5e8HM8ORFgwGJYWBpclPOk
qt7SW1l1HSkURaj+maDdGVIr+UaXJA0V9sKthjsZ7fXlmyXjOXJPfDMRr8N/XeFt
TBRwb4ziJupG9e2QuTCBC5M/ZXGiI9tFbU9BB+usbX2eRcbqbfE3I15plaB1hHL7
jPq+BSCyWToyYlwtvBrFUA1u//4VlaeMTTD14QaMf+a8e1hSrfgZPaV63w+Uwnvo
O+r6KFqRVvDmjHdqTMi3545lPZNxkqIZOzSQhNQsiMXHzK/PwM8TZT5v9OmzMdQi
b4IYsRTJhJvsEqgfxatmW2Ni4qMei8B9u2y9bBWyHEO2Qz89wtO1+uHTS4jtjoK0
gd/jQHsR9FMYlC4LDeld9AIDUw4faouKdSr7/Jx6gpfZ6w/bCILDvU5ukdbvyTVv
B51O5LHw0i4lJDygHNWFqL+49n3N7LdzEGvw5FIczInKpWbGJqM5KHhL5UVUnmWx
fRwag+bX/x3t/dEuWItx5tDOj0u+TxWU9JI46fx1k1cU5ei5HY5rVCGpNEnCi1Fy
lmQ4LRHRiIdv8id6VWf8sHfmphapewwxbVXhZDkQkpV6iqhJ/4wwYmWTLwkVMRlq
RnCwoNrKLC53aJ1ka7q4tAO1LrslsZsl9VdrwmjSrWf0kFZoB0Yf9tE0wECwwjS4
cT8Ljzmip9eqQIrHO7RYPVbaD8jAUJNLQZBVZcTeC78xaDcHT0GFy6wXobBsaIhC
4mOWbnM+S/2XWJgmV7kR0+C9XkQpiGDGwODKyIvLtxCqA34WFMiunDcNAXrDY03P
y29Fah3vDFw6bYi9hQDovsCn7BosEdPudvuLzqUTgJpPxPd/eaUMGeiZGK44NDb5
izZAhmWKXz6KYw+VJcOAWlDLmIIuVp79qUMSdTIV4Pd3CjqlWgFOHp70B4pdlLUV
qrqCRgTwrTSGEoJLJR5oijSFL38jiSBo4xR1QVFL9TjQbA7lVpuM/+9KxPw7iyip
rHV2Udd/w2rX3Cz4tGHZjmk8esRcQ2MWRkS/DYNWMziyKfRAEvKDRJvkoAia9i3W
qDAZRhvWdtbwpQwxBBZJ6oCDB6KxBCp9pDPeMMyHmy4eEMUHAm4qRtaTUUanPar3
4Xa7dPXpYa3MaccECIolxf9Pk6biG54dlqfEywfii5VZE/wIctcrJGDl+dvGCcDu
HtepzHfQbSIaM3yS1J02/uahSM21ZolhOGJP4Fc3GwJJLLonINHmzLcv6K9WNeLE
JyOYHmqseE0K3NfoMVx8GFfMvxHTN0m5pqxLWaBOYWL84AoH4FGTmfreqvQJxPLX
5cR0CZQ6F7zN2rGQdef1Io/zdaM3LVL2+YMVhdeR5BUwhZXmjxPchxy1suoSsqFT
eSJj5R+6kGMYPKI5OnntZoAiMr7VuwKy/s6ev1qlW1m4QJ7EMbEPOGQBnmdJuMR5
fPYepAFZL/PKcgTndbuLoS3nZ1GQ8pn/dQkKDroloE+y19bm7sN+wTVQWuqFSvRt
yNcvgvati+99LW3x+cyr3IQ6B1LuFg44GaznajbM5HBCalikDmU1TKFMa03+VHsI
0gAMNysmHQ58/V+zVmvdPn2DR5TrSUEvLePpukTSRLflrjKPR3uVVwUMXIXc7poL
TmRFnbLCR2aYc5yQRfTZa6vJvQ/ftI8AiW0dx49bAoFJSzfq+f5B40LMH7XzNSzZ
Ev7q3pZ5mQA2Ijw5rwyosPc3tiS99P/TFDHsHx1aImiZOsVuUx0RqFfuKKJUyeEq
oOzK1+zy98LbiZH2FfJLMGh/8CP3J35p/aIwpn6sm02DpcUY6cGE165YMOHjf9uL
pp0Zm7/1upnGcT12ORd4z2JgaoAyPtRCHZ0VZbRx5kUHKePCbzsrbeoHd8MkdXb+
Jti5H34hrvoP1HCL+m1UnFxtiOtjQBzBBLUap5LC1+JFUT4x88AHDAa/zhuGy9u9
QEf3qPUl/h/ULVVDfKT00/i77vsz/C426g7939YI5DlXiTOoAcCd3Qr1oZHVAR1q
jq/gEp6Rn08lTupd8ZyADLt1QuvCszi5eVMyzF7PuQRngJXZD67bqSJNudRlYFKh
HIN0wU1cIBIVRbAND6scKFf92zuEnThtUUBsJhHaMoIteFXKQciPGY9o6OMhZiqK
l3WYGrA68q344G75hP4Xrr6CsJdKrzkJrI4E01C3lUV08bGoSHjQkpDL5xrlUavh
ycZN4EcbTgbJYB6qdzOgVe4OMUqQBwb8z1XqXA1DrQreV9g95qmcuqPvjoU2ZS2/
96aQ7EdGpo0eXDMbnBMqd2G8tMDsswPer5jiNZzztyZxDVYlDNjzZruTYOPiPPUu
Hq7sptorNPH9bhDs5UH/k2OPftT81jYl5t8ueAPqUKuUnDjzbXFMy+KqxuxS8Epr
NaAezTwhcNOqt+/SBYIXWsSRCx9Hnzzo9mlirr4sTy3py5PRXUFZcw9t/5im402E
5tW7+md0pmH2FJe7pYJDfHXVEU2XSo8yDOnXipzoC20uJWgSU4SoIZXndQXKBEFQ
kcxp64tLlDu06rIaT/s6XLMIVLAuQgCPRQWi3UQVUEs5/KWD4mujffMAs5FiA/AL
929UWMMwyBypArw3lR9s1wkUhEWg/bFLROZJ/GDuWL26qQlT7Jz0PzNK1SUaJIob
hs9W0pG3d+vsAw9I7kyzCcpUT6UnrLih33QbjAUx4Z8MX5DvgbePn2qjUHZLMvZG
KY6yqefQLcInfczcpwm77IgnCLeAn73u2jRwLK1e3UnLp5uztpyHCUeeFrrfbrYi
07t2bL44rYM2QabSQkrQfVcdIhJn9CaLkfcV9BnJBWSYPxsbDngEctmXunVDA7he
qgkbILS+6yLGblOGPk8kRpNVH3zaDX2YXTDBRXPPt97t7EDQicDZzfKUpd2eoB/C
YEOclwAosIJkWOIwOsOS+9UqSXzSxP6vlcfEpE1Q3n6GOL/CX+dBoxTmY9mOV0lz
bDQfqeQnZ4tMjhY7lw8hVOMd/S+qO7kv7HoZu+kWljFnsSivwMSJk5Vr6jNzpuW/
/WE9ulmnsk4ApitOq0qWZnhxUS9jv+LdkOIG+QuDdl45JmpS3XRFqtxQFbRxh+Po
ll7t5oskuEYdOijawWKVtlzbAi2DeerS0LqWVREFs+6mCIwywcLHsRktR3Ang5ye
C/jCV7WbCvpt4ir40YSrx5+o2s/sA0LerR6rMt0FpxJmDdfQ6/KCSdJLiSTaC59D
P2S6hcz5cc1NTXanVUQCsqAB9pBSaEfZvFyyTzDINFNKIV9+MMDpc5LgQBr5scZJ
K1g0Thr76eruLml6OIB5lkeZew+DU1QcnBIe1kE6CL7OcMPZj34Da1BLjTWyJcfs
eYnvI2LIHJS/j48NYvw5VNpXzl2hfZWMbLEsdDrqpEkWjq29sI4cYIcSASvLCphB
HYDk6XGzcxfEmf5Ol2z0lx6T9+52x4KKqEBKAcJu4hF1Y/Sh7sr1IcS4h43aDbHJ
7HMvO5jGhrxcqjvSH9jo6lXJtiJu1W2+rrJb7298wEGjkbdDpXq2WCADYDF5yz4J
ASQf1SE3ONUgvs6BvCVSvyREzN0VsB9sltPHZ4ZvmsCvACILsERxlHtjg+RMIrOl
MHoChQnT8CEyI/9qdNHhHXs6l0KxJUdYhMgMZh6KZuj2d6I7kNOORCqGBy4S0h5l
GZkC84TGM01ed1VD4C3ROCi2QXq5p/rKzI4ojPGnACsOBZj7YnKXbbqZvn5idL5T
G9w8lMqqhUq5zxelJ+WpPRW1L7FeG05dfUXjcaRG7VVO5Iqsxgz0OcUeel0km7mu
vvNStYTufBY8/OBmbnodxcjEthxsFvwvvCiyl+fTymBFnXZzlhKHzZZkGMRDabaO
cjREI8mPhpFTdHhjcC1JCAdE0WBwfmO6NIAVsbYAgSvbJ4K+ekroMSsH0zcA5/T+
Ug3xPebNOpJYr3f0TNHZjh8PB8/Es5jBtXRQAwClElWIzhwZ4YmE1mmXOFe0cxY/
RMbFj35DUbbMXhxajMV4eRZCVwpBS2Na230JlYFqELN9KwjKN0WykzcaWGbmckwh
Cny6Xmk8szkfrdtwHkoj1VEzpVz9lYrq1nbHb3afEpfLqWSJVz5kCwJib7+HeEwP
L/hx2AttIgNCyUsF3nJKjNlYQvBHJl+kezBa0yJoF3x4Ywa96+f+ic1xIiKWftSs
7Bndr5DSF3q0jfP8GiHx1PAy0ESEPT1hWcyR+mw5RiInBlWQK0EAOpNK8SdTB5HU
oB2S8BLsQz5L8ywwwBt9jWt0G4PBUzBOs19Cp8BCJdIQFmlxbQ7EOkbiBVUdfe0/
QjmgI2CZoOZMN3pAlVwVqO81cQaG2sO7xWGI9yZCjYNQ8AhZthf0JpI/GsW1gaXZ
bciI4kL0sDfGTE4fg2+B6LwW7b4E/hGjo7egy8sM7D+r28lJVYxk0Fh2j4E4ZoBB
5oPfB4gI2iTWM4WfTMOz9+3+S0Tofotvxyp1vTTjhGObN5Vs6+AS9UWFQjkGb7lr
Ah4swxRhQ+vu45leNc/6mximfEwKuXUhqdAGlJMuTQzTUkv0PjRE0qHN7cglzO2I
7ZMGngoIIQWQwj4rIKy2IoovmZNGv81nA9HAvARNMVp9pqnHJC1YOAvv2HSwknqg
YtEFZXCRmwFW4UOPqdNZlOlxdxKgY/aJnUaduqeEV9P7ClxZXgSZDAarlPvwViMV
GYqdSpJ+oCZR6DuHzuLBQkEuqFIIfHlTIo0PRfaVPnS75ZGchOMX7RxMmSmF2awL
j15EBgR9x5R/JtfGGo0ZBsNkj0dmtjd9YF6LTEN4wYZtXyTVzeZqlZTyCt95NYHn
L0aK+a2X2KjMbxBxZA7tZs02LdK1Z3hFHYNsJ0tEgDkn9QHer3sQt2vE2lAFj6oL
7WmXC72ubO8gtXa5BMFTGV8AScQnI5paCDexDBO3ZbUBxJCrht93HRRTbtdLjP+X
QhEXkF54SMUa6dWYAjBrMLzIMY+AkSozMvGQ8ruTBKP9LDnwble/VtEW5rq0e5jv
lw/GuSOQMqwePsIIAMYYZui2q4QchHgaI5q8i8RQ6Nuli2a03slgEJH7cBQYdfCg
G6znXX2SiXp8hWxlR9EmOKPfkH4TS/LgHqfkxet5Cbz9ZeITHXWcfe/L0lucqth0
ngCSwBhDy2G7EiKXsurpNM/NjkG/qVo9VSQxe2++VCGf74R0Pngm2Dp/piZd4lX0
2BzZVHT6X6JdG3+jXSSQcCsqI/SJn6ctdzxeZeDrqVxfoFVejs9bsBoCsA883r/T
`protect END_PROTECTED
