`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LB6M17Il5umG4OT4pnHLOZ6k44z7NrKvi18cPctAslDQ1yzOJF5JMB+3dAfH7Pkr
AgCu2ADoZi/Y1I5N06CnAIlUNg8dudlXN6izRYxr6OEmcxmBYuvgS2d9nLKMMkaD
iy82cQJKzzG68TYUqIGkFEkFfnDyjWsylK9H6zU7asTw36JEBfMipI+H67mGU/Mh
QF24pttPIF8JUKod4SaEIMCNddQgMDIhjWhKnEcq6zePQfaf8oxueXlRcks2ezSQ
roVkYJRu0ybno0lxsdkocQ6fUEmk2f96ZA8wdK8cMBJxzLpSBYDdY8A9qgr11845
QHOwUE2mYp/g17Fg+m4Law/Dad1YeEnoEYTpteypq/MCf7wg1J9Z6cj36lD5Grub
Ygx9PXx/Dl06GYpIAerCmGQclKUvZpgyUPpo69tq/4z3dTATx8psu1mSbtpNU8ld
5BPfO1Lz1jnvL2k7muhylz44f+fXIdw/zLOwAr7TTRNgehAK2KwKO9d9xLHb+e4l
rkVFe3DkGiRZbEYtSJSs6uWCPG071dAfCaUr7vzsmVqiXy7vHzmrr5r/dR4g/wDG
oZXEfHFdGClA8F2aLq+6ZfmThQyD50oBwSo2D3W5gJrH9K9lRq/IA0GPTRdi17dx
knrW015aiZUAIvLdkAKc/ZTlx3ThzV20f9lSKpNETqw0vWUZL/iCvMHK96x2luOq
BTMN8Is61JfhmWTAfKYe5A==
`protect END_PROTECTED
