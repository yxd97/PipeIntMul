`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mrNU9qmovtm5m4+jJmE4oAhjZ0rY072J9LBdOCTveTVrh7oXsbhC+YLJrlD63rYc
VI3UmoYp6YW+o+cvIgjKfhFcM4KqWsJBfeJ00t2jVkGffqM34xBIEM4GWaZAcGrv
M6WvtKqRWillsraZSdfHeyewnOe5JFrudLX38ZO7SAh9yWsoO0DS3h5F9gsOI57+
+CCrV9j0mrG0YRPD3rZtg6qWw3QBWtQo2OOuCMEwu0oBews4oQxNvAapFoV7FvWn
wrTR6tFm9612OHUFWacsUV/DM8E7wO70nzpmrAYzMf8WhWKdV3FelfhxygwWjo2U
sUy44Gr3GhfDBM+ggaLqFkWyQjhsJcFzWH/AKbkZry7cYtSIyu3izTmegZ0NGLir
0z2xS9veDQVZ6Cx81mJwZEYWrbEISK9kuFvd4vUCeOhU5qEs68Jxw0fKQLBvXejD
MAg00ECHDGk4BNw26tXziRZ5OKZvMKYShwjq64QqoqwmYeZOXVwQlZbWSmZBqma7
A4xvVNVeeLqZ/w4WEVhzNlDu9pix7D+c0/+aDlKr64wasyxGBGz7TBMq3j5vIivD
8/mDZ5L88bkf0SkJg9/BpXG6x4aMNq1YVu91IxAu5RA0Db2KnM0XFXzFfH+LEqhl
8JQ+KYq36e88y9m/hF9/wwNEZf5gJHie1xjnOAJCtl4FztRCTHMybo5CyBu0oyP1
1sbjm0aN0fV1Njjl7Rjj3BCFCMQ03JbsB+SiXDTX4NzWg7/oYOgS5K1mSwwm2zgG
gy/v1q+RP6PBpCSGVFawkpz0shjM1oTADCcL6J4mRb/m6uCGH/gRXR2ax+WyFRCU
Gd7Z8MQhwvl6Usms8ZcRROiG5xVTJqqiJg1g9jQs2iVlAONSLGWKyoj4q0uTcQ4h
`protect END_PROTECTED
