`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kq734eSj4Opxkp6OFBirDsKfMzDXYt7ix+FIEmov1tO2IEDrVydTAM0PRa5ncCC8
kSdJrjII6r21V6keFmcr25gTTx22I+7O4GfnKvmD85ZUoEkWYjOdP48qoQCiVis6
PWsq+7DujCHeD3IZWYGauQfUTTVU2o5t/feaL8dm2OFOs2LSIph1Kaw/KjZ750P1
gTnVc5zwqe8MyZ9GVKOgla5nhwqJDTQNaL77OaUyajdLDA5AorZJHoMXVp101Mjn
ONWwIfQvni3Lf29kojY8tfu0X5Gtc1Havbu6Sq/IacEcz/hH7PyO8wlrj1d36CMD
vVU3bEEJAFa/gGb4bTOkqTiuyNbR6R8ghSxAaK2NTMeSkpX/eIUkZNQqg02gCCFO
IJSzKtkLMlV7HlU/4RR7GWPdxuY8q+Le1Maf2uPhojWVeumZI5g5UMGui/xfzuN1
sKS+4WY+x+P2Crhem81BaPCV62pm6KJ/eSusTtssDbwc/Kq7Rhm1yrAc27Csoa7v
`protect END_PROTECTED
