`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gYNmUohtMOMlcjbzDNYZTgICShzWiNAtXwm/2VXycXFehQxiDxWAD3HOeh/sOD4r
FwvqZbbwl5QNWluqjyOO7Z/vjQ5ZxwtamywFsmKgoumtYPKAuRGoYEFJgK9VNk7z
lHEZHSyT/eIDGBht2IEEIg2/dpfwvg2pObtbSZVDKllESDgg8TslDgORYUV/JIdM
X1+fwiMNUtrpVqM7mPUK61FJTfFbRV/47mn7ak7G+IDchhhzvT9ahmrjW+SrTjqG
6XMfRRrkHHrhny8hcGpUee3jMzKtWoEuEU0ggQDoLkEOkVaQ5HAOp+ff7ho+xv9g
xH677ApUJ45J08BP7oXGWf5TyzDHtsq5mlLlMoTHm8A=
`protect END_PROTECTED
