`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pq05M7khrCuglLnn0z9cZnHjlEZj5gitvAOVLiERELdid/7T1h77n5OAn2dEdFlx
b/3MF2CqI4QHVlJnx6tvphiNI56j+s9rVbiOgZ5fkanehboTXuOFd4mlRfwSAoZ7
zwOnmE5q0IS73N4W0NhhUwG60Gaek/Mm9GHeY+c+kdD/QrgNgAOQscTTnK2UUZhF
oAQOK2KbyeBORtHcWNWVTOAERUEDUJSGuYaVIg3zXEyHhD2JPrU/1do1bea/725P
2hJYhHH5aecwv76I5KEI+w==
`protect END_PROTECTED
