`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hqGDMeHW6o9te7VNZsB5lPq3u68Q/8qaeGgGuweJbSeBzaIpiM2ZkoTyOmv9++9u
NRbk6tKzEJ48ssmE+ooey8zgQSC/4+damS0UdBJlXHlzY8Y9KzY6b4KjWBQZXvx3
j2nKfe8Y98eEevGyrxbR/xxzQM1mFMbRM6MAyBBWl7MQUg56whqqU61BItbScIvH
K9nVKb7lCmbafsYc9KQuWd8pmK+iLXnxfBplQSBAjocCK0iW5fKhxK4RIwkSnrdk
z6fcdYliLWw7bgUxVV8XUgHs+KKtnA+BLMdcCr/nT74tXKxD/7tt5UgkWnpMtwp5
x50KyF2tK7B+RT7MMsznyVVAGwElg4b3kgr1MmSnYaBWp0oREh0ox7JGyLOrKYDH
6UU2KTHsC9Xx5UD5/gk6gQ==
`protect END_PROTECTED
