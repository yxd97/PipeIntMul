`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T/2YY4jk7OiNmnCsfwlaK8KcEPONgkIAshcsU7zzGoAmJvM14afDBARjghVcGZU2
OTZBrJVgGzrFSOWDjctCg8kd8HkKNiTq8yW6qtB/LHK+KFFEdL+fB153EzRvkbYJ
Pf08vHFfxmxmyO13sHnegWPODipiCaIku/uCDqiGtGS/bewUSGEheusZRz/+8Jjr
1oHB68erNKiD8vD6Hv81AtZAIUP/g5rTh0L/wCpKoOq63++EVmzHuKMKWxAZT0ll
0fbAa3xZktGzL1BRWsIA1Bcz5pPLKepOdHAMRV5r2/R/AHBC5CvqiIrS2OzcL6+y
l1aksgqxDCLw953LSvPCpeJUnNhMBiKLc6b5vWbc5DBdt4kM8qtAOaJM6LCZEJ1d
dxlFWH2+YOP+GDl7RpR1X+M5fO8lTqn/IJ/VIV/exSWEcCMuC+QrR9wk6P5o5PZS
AQt4CEs/dHk3czY1gPwbPy6tOAOgLtcJ7YT6PyBRdkaigNyYH5kfaY7MBcEBF0y5
GRk9drHfi7RMoIaxQSGwLRpIAjOQusWB1dqRwDdeznRhl+unW+r1e6x3VgrBOmje
vtSmoJttjoFdhTaxV3+PoRmrGTNIbEnr7QcSR7YuJq1lsVs/DhXuO16/erumR00g
JAy3Ib2bsrpfct0/pwG/0A==
`protect END_PROTECTED
