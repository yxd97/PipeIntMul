`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOLfxIcEnhxSc6A/+SNhIrVCplaiqGomDO+OMj6cPaWgd8uAwhTYQ+0NHCNuKsmQ
s9FLJjAD4fPD9rIAvDpqhI0C1+qE/+kLH4w1b02GsqrYUFEn+KzQsK/7JR1re1Bb
jvplm83tWzqLlStQxC1QGXgPQYL/YwMR1Cv0EVTSDekUCLIOgIXkSOv9CVeSMj2O
o9jVjwMib7vLkzH0+PYBPsncCM+Oc5Qyu9L2b8NmBzYPbcLIL3rV5JJ9/9/KfgQN
RsaoudNgW4+Xez4T0AwOIqUHaqJePgJTMZ0qHTYoQxms8bUWvccdOQhNs0aGTstR
wb/oVZVPaoe1LpAnIl5trA4jB1QUAi2LSt2g8T4WHKQHTE+LSK3ekCkgele5F5rf
Es0Gb3OLNabNCJtpWelGpmIbarxzlExWPAQiFthMIwyhMHJp6kw4xhSBEX7KMi77
O49cBEpE0AABRbGiN6DN6kIrvtNkVCHX8akVczWZVTn8vQFfxM6bdImesoHCSEH6
1ZZt5ful8aCOw709Zsj38VZCVMCgFq9cy6sOgESad2+/kTasJ0uTS6sL18NDXzU7
9Vful9VrL2RVKrGJTNA7FYD1B5Cf4VREJAwE+UWTtxgWmkS0WcNvhZt6RCHBvMte
`protect END_PROTECTED
