`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFJC88ofjgA8P6mee2EcOOj6E0XCTmqz+QjEDhj1QSO9d7d9J86bEVxWa3IBFuAf
IVJBiEf7Q5QEgF+RUCF4kWrYND0+m2ULkvEbfm8aObK3m5mqYmQYpEvEhKpOzxph
49pAlnJFASqAx1w63WeMOrarH6LcL3C6IjpXo/vddmrFGskjXhVTZkcJzJ46ZB1H
whfOUX0C4Q/xsSmO/f17LguLqBvkDDt5q8TgJNz0calLbbjL+ShUDTV+Uo+Qq+b+
9uGdhabPg8XBVDC4z51TDqAqZ5OyaoU5B4smlY2nK8NkgsDw58+Fahu15xVTnjqR
qZ92e3GeiqQfUrHLnvjo6pK23cMtmq6VihzbbRyMXDrCyxB3kJIs/6mttY4EG07U
XJPyOnFU8EEVvnn8X07EmVu0VWcYclOJJ/DN1lvqMZwasCQwsE4wMIKBhxtqaoEJ
kJSh2CZtrmy48LZgMxcojFUXG2CI2P6NDpTatMGnHoEwMjkxwjj47CRXKFNrk3Zf
nYCfkX/W/qFI3X1KIvOu8x12jThfL95XKvb/v8kt8DP1fH1sIdL+lGyL3Aytfp+r
GxvmRZR3t8GS2Dt40Z62Wg==
`protect END_PROTECTED
