`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYMN/XfjPHy2xr2ASMxEjq/l8ZK6fEK8KfcjjeM2un4LAM9vU/fg2SNOVh3bPyyC
YN07/rzVWunVxmOiL6aPV2nvbsaOWuZjS8jwdHlo3U0lzzr9ms5OPLBa+fMtK3uF
3IffQxzWTSLLn+sJyc4ndirODLSRb7O0CuWOK4LJjcURRfJxTeavrz8AgF1NfagP
8ifvRcrGQIppO8fMfkuSuKdShngy019XXR/cetZCAuD134SeSXdFKz+IGMwunJb5
y3f7IMrqNiMOuDc2nwOF2bjoDVkrQi4z9t9ngBv5ZYStO/M+XhL8UG7OhnXTOKkV
q6mX/MUl/sqoJAbuJFEYLAHnNUHfiqLOhVOMUbrSaHqaw0ti+mufS5Fa8fBUmeLm
wRDxRn5fQGAyWD6OaB/IRovHZbyRfEEtXMItPY0QQLmjFl2V+LAl4ZcN+4FrO3uM
cyBOtipIw9auNol/VF+wIWUrPqigLX+z70apucxP8KVnzS7UMjGuLV1t7m4XnFu2
DcB8v7ogrTkp0GzDRULixfuLxhgYWJ7rWwbLESz4LQBcQP+23sv/JZ0pwzn/XR09
Wd+10A92SVlwJ0ZDBRZkwTzjLTYlPQI6MVlM1jann5q3zcbNpxGisHA5h4ZW/QEl
SMjt7C5Jwvxi4fXH76UQzROPzPUMD73ho1ioXGmDpYANgBqjCbU7AazQwoaD9hjG
l/eAPA68fPWy5+uzZNow1HrbeKI2Jdl3HfhivylJqzqPEc4ccDBI/qSDwg/vgHZ6
V8hAottLTEDIrDM0qBwD9UglTIzT/5S85GssuiWSa0B01O+uwb8IAcAu7g5atkRP
7pnn9EqDhpSuLqmW7vHt5aRFSRAChN06qJM1IFzbXRK0Ffk0O43CsUOtFpQbwDR2
OqSDLBtchDkU67JCc4UD+ogxXAqszVKFNpE8xQXSIdIlUEvfNAjzQZqglkx+UlLU
lAngwRkXcnRoFJ/H4huouUwwYUhXKXN8KolcLpxyQju72IZTO9xv0QCEq+bPXzs0
w97hfbpw/caZb28NhJQlqA3UYp9nQSsgnfvFsVU2DOkoyCT4HZQTvGVkqzXVAjFW
/pNt4Q7PDMfmdQv2jWlA1suvPs1iPj+ueEN9e/CAqOIDsFa+zhGEuOc5Ig42TMB3
q7iyM5mbwAbvjgcRZ7a0tvZVLI4Yu8T8T+GnjISKCKZ2aoaVJYrrxj6Fyh+bDem2
+Im33G77cFaXe2NVVqjH3zZKWolf+adNsgINu9zCx1w5u/SiAGICFEvwfyUFNfXP
i8i8ZggI37PE9WBlpe3OoqDrtdk6vrmFaWlC1oQ+bLec4wqsNZb2yWbbLKSWVRp2
li68Y5dCtMBY+/Ov6t4bTglrmdLty+Co8Y/WMoqEuFQUJG7AjfSYA5nV1wkIm+xF
U/AqINcIlUn5e3LeJ1M9jDt/zP875P+/Cw1aV/7Clr6sYSAchXSMVK3EPJIx6rkp
QQSOeJJN3a63u7hzuVw6fsp/OzLycpZhOa8ZzVDbyDcZjJWc3onORfjkOAE6Mz0c
qx7CjDOIWTl8la6V2+1v8LsDh9nGpRfB4wA2/vbnV2PZ/EqlWhzUI8vkUnLE7QBP
mhlxN0gPKJCAFBkkTTexh0kRZSN2IkokfOC4nISzrpPO3sNRdsWma1Mt+aS5Bone
v138dOM2Mcej+XMXUoNnn9UiJUrrXIYFWT0CjkpF2LLDvNoD1fck4DWqKA4jXVFI
7fEiIJNCJA6z4Wf2vS4oXZUp3RPTqSg/nudyvYKSA+cd+DD6w28mmtvXvBpwvxCx
co2gAuIqiRMuYmfwCQfQSUe0oHCy6siBpEdPvT27aI0LXF7bluGi7UBmyHPfjbQK
37CfUTWQ5/T/bfRzLWgK4s8+ILc2Tk8i18MZ0ulNhWOR0EAXyq0DqDsTpy7FpDKV
r7AUKlew4YURtxaEwiOUv/HQlpfHnhXyKm3RrQjxrTiAynMJLCLlR53+1kvBQgHP
w7do06l6n0AZkk6RD4aIZbJEQ4e208VvXHUXJNpYZjH7DnKzFmi3pChi5Lwuq6wP
mqhS3m4vxGiV7QIcztawg9t1DukBRzraGrbvk8oUeRMywy6xv83hhNw+OfrUWs4R
Jkzb9qxoyYZSrTeg8tBVKdV/ZOFBjxeSnVGhPmgDLLeDnaRgqZyQqk1gZ/wpCzN9
bQA1sTbVhBFl9mxqqjQy2dIFFacOmmsDsUUW/qyiVBpwF8IvPphWoDrekmETcxyh
GyTakbmsnVKF6FTPckVcnPqxktEQobBv9B/vSIs40uyei2x+wwEzfoC6IQToy4Da
35gejNXo1BQgmKlW21AUz/Q49YY9ZLBgehHC7CuxpuNzxl6/mP0kcr2ZzaexeOr9
UlHwgV4iOQJEy4KgmTIlsBbNLvpR/UDwA8rz6cTHo/cVP5omNvtDn3F4WvCJlKfg
NpPw1j2RICR2xbzdf2RJ5eVu7L44rZ4QsC9jy7HM5HWS7TdWzqxCrp0Y4b/WdvoP
gmjhZSob5ZYDHGfevEjFyDbUAvcJCg4iSSvSfT51Z+ETmGJNZu5sqThcB3dZ3K8S
Np8VjcuI/ZBswmkmhVdjf13Phb3H+gnZlRxapzttt7tTVspmdw0lKE6Nf3pz6blU
374Vrg0x6kYIV4vUyIWKCiI9mqG8DhOODjn75OVZcoF4GShrVDAFrcmfUisDo5dv
FxKf65+uC+1nSJNlIiDC23tpAeJb1m85fJxxp0bCnjfiAeevlBVyf+sGQgRLjFce
0ZwgXELXpFVkLrfGu3nTJfYH/oM9is0mkOWo2CWDGj428SdIbjMeZLGXuxuxLQbM
XK9HPb1OC2gXTFieyn+7MJerGgU/Th/6J9s5RF//E+4kKKViw2uckvUuRxTg7UuC
KiLbAn24P5XX2GAApyZFYzEO5zEMqkebvipe74Z2cRASwXB2tO2g4Aavg2dC5Cic
nDVbVHLFM7212oRn9Rmime99KrgYdGt4ow8znezd3ZSJ2eVubGD0Rk65cuB2Xgav
dhG2aWjxD0a1V6ZhXUpL16eERqAn0n/XOjNFaBnT3rpP0rdniKN3X5aCN9nISHjb
gjNH6hXjEi4lMKpuHg3UdGkTCGhuiWZGRo7yRzBB8jCx/hngU83lbOwSlX9kYgaX
tlz4BLoGa+/ZumMRCbYOTa+xZUC4ej2LewE7APBHxaFYtW0zFjys89FnmY+4NfbY
zdD3XwdqNaUbiwT0c2r9PTF+0Rd1XJJs4BwHjq03i3aFHXLeoxI4LKfH8UnbzaP2
6YySvxblbutlSZ9/ryoT4Rz1zuvV6YW5p4nR+NzU689XToQSAcXz40g3bVba22ls
IV5j5FWdLNEeqq0Wzr4wOBeNQUnMq3ZOr58p/eL+MWcjLGEmE2VO6Ala1Z636Kt4
vSsA32rpp+U4bu0He84r4cd5MRUZyMmMmKRozWt5USXqO+fzQ743kHXF63aywWCn
44newFBgrfCzJB4DlJDaDRNr99wXbw27elgRHM985o9jku42NSCX1bxGL477Br/W
o7X8EV9BvxmGh4VYyLfG54ZQ4ktBba0LRFYzpAkUz8jhxetVl36g3BkjuqzZ7jF4
t+JBVSyHaOfsO/E6A4Q+OaHKOGv4j2Oll5UDbAJ0K9Ag+DtBXSU+iVZuIIx5nDQ5
/WyrILc7yEFXnAnDZaig6cnKae9JuWzKJYKCD5kQJZGTHqVMM1+X/KA+Ide1KmW7
VnRLdMK4xlZk7kUS+j2+//Erw5lb5Z/qHPN28d/mfB3nkLcbukjDb1A45bp5NLKQ
NUEen7t1TLD5LpHHI0nmPJsu9QZ7X+CHyCoqTguxYJ4nBzRZhsAZZnassO9H60yM
tCgkotjfgqOmqe4jiduN/EBk8fEWNaFajKmj1Fpi7n6E2SitJ2IwxIfuzSpxl/lz
5wo7lwW1ihQxQVc5HZDT+YzfgXC6TaM9xmx2jkM7vc5MmNuQ9yxYaNxuq7gXwDk9
xOz2XlotL706piej9/bPL9aDeO5C3KIlNXTjktUBwWlkg2x6kPj5KDV4Ii1EBRwR
4zj1XBzJSHThhDj74ddoHaUW9pxENAqPD0c3HktKL4/cNmd/3shaPk5PJEp4IRJx
lSDyyjnCa8xMVxtyPZjYIAgqOehu7kKwPErrqdAo9slcx6fDHYdYoUalBagRf0yG
u/Zxsm1o5IrOkQbzs9DWQU3AuGJRgchCeDTjMUfW2TZKNYJp/scSw4yx8Ev10eX5
0fDXeC4eXxUdW8RY3HO6Q6rirAFTlapeSlO+PJKYsamSbwKcSCsjubpXjmhgawPA
IjH+/cj1Cf+V9miaUPNtt7tMUmmTZq/A64HZEHuKq7X59V2TQYMskZlTQq33z5TK
BuRW0mvvDLSjXRzDpz9JAZkyxZFYKyT2Sq8u24i00mI+/EA6HAfId4IMNogBtJHm
lzYl0PZx/f+qns0F3UXrgPkk3LI22AM7WxSJmtZefk48tpgIKqhmjJWOBGE5HKcQ
ABTpYUI3t+774b4gn8GcIqeawcgm7395baMZQ/VkBiv6Rc4BGamG7qterKDWSSaT
ANKVIayMv/LqO586qpGWSZKnGsH4if9dYkgV9O8t1fpNnJuFFYNF+EO8701dyQVG
fwWFLmldF3xp66MpYZk5hEjNrVIrk6Qp3S4I57tdbWvdWjb/RXsEAX4MoY8a+Y6p
3WZlq8NNIZ/mz7Jbnlc3LwxaejN0jYfzbX8hHratDzXuRk+UExDI8Cu8YFxPRFNx
oIdCpQ1vTUaeUa/C+qWEcnXueDcXJhdjOeppKlLfR+fjc/F8vwxsrMvzIaqUC0qz
D8KMj0G/vPxVxfxFQn5hEvhgPd59PJlywSxdOrnC3rrxLCFDY5e+UjhPnOXYu294
JH/rJZDsvaF9UDIJ7z1PoQhf/MiNT25Z2PtZQgG7+xbHYZAIKdzRnZC94fO6Ofcg
x9o9SvVL803Lo/mmL1FsaG6uUrCzOtR57yeSptDK+yvr8Gd/+/8AUClCAh7KQqsi
le6IxPu+6p/SVU5cwqrwwqINMtXx0IPcuYUBOXG9jov+IcGI0j36wDkRJhdjZGJ5
SPhD5lrFKOcev5t/f4J2dYR1eqaS2D+kUlYpOQ5SRC0diTLpWqjJTWyLy/19vt5s
WnJx40nX45El0/zzGf/S794WQyprD6izZSRkv9BDegublA+HAqE9dnXPpQe9vjCD
kBmTUmjUFb62fIRHdA84dqRwBJxnWQxq1Sp6rOgImTJ2qiEUnIiqRn8touaAjhTf
vq0YPj8urHCVTzMCWpar1HlTjFhYiHSSdDYObtUT39g/ClSU2tVhm8SAMDN4cL/w
Tg6uf+ZJ0wRq5SsCR7D7W36SZchAAmZ8SviCLumR+DZUW4TCfxSq28uA3pUr7FBe
lE4sEdANfPjHctXuABCtIi/SjhBuDfO1dVeqcmDj7/Q8emrr3KIUoqDTTVgA2xzk
+FIIccBSlfx5aFzuWaC2S4C5NOG56Tdn3fIf5D3CrXqQaun+I8VG0VHza4qRozJU
llOUPL1Ij/Pmn3VoE6EEEG1gD5YLnM2A8QhLHQa0u0WpiwBfpn7NV1+p/WqUwura
em8eLGsxzqznxfI/fb7Ky0tfEqnxWeMPqm9jPW27RI2phT6c+TsaMYaHBt3i2hnj
1pGo1YdYTr6JCKoZA9SGNDfwTmaViwNf7izn/dnVpa6j7IG9m4i2kT24bspq+vxX
Zz0wt5tM2Lh8KfJxVo5SGdoi11WUWoI4viajTajXp0KQC62Njdb+e6JEh0oE2Xzq
eJ/YP9RRZIoHJJDcB2Agkzv7zPJCbjocAkT9oWnBvWp9KiQd5AdOrCJQnVkq6qt4
uKzq7wxMMjKPV1Hmar+RBylurHrJuoC3RWu8Cydgbsrm1zZy0WPfTuqxjVoAQ7r4
RxNdA6R8cIDImRJaji1qvCbNkmCl58VsQ+9rdziSmumKznnIDUHrmgokrk2xCg89
DYdyXvRxnJ2HQoFH0/esiIL4OLBzMUUC45PFovVHM33P3gg5+Wpzu2fxEQisXbZ6
cydDV6X/u3yKZYEpa6/KDdkZi/sS/rp1I6nP3Zgve3LiuT32tF0KFgNwQfh0vvsH
OXrbyyUDI6O2esCzhIVxoNhsCYoBkadsHbO1znotg6WfVLohqhLt9kDAOykDOYIK
uEgSEu/bZlG58VEy6v/bZNo20Be4qxOUFXIzKZ//ce9/TdoObuvyAZCYgHqZevkg
4FKEK0c6ecU9b4QMssoMNh5fzE9UHUCnP8Vv6JsP8QCL+HtKYbpzaIZUqk26pM1G
UoZxQQZqJKYu+ltGeHxa1YuXI2NYKcOh7zh+gk7nputG/yNr4IRckahvxfXcCvUz
kogmk+j5sBw2tGgB8n4RR++w7O5D1wjrQLX2uyTl78HbSHJ7KAA+PqeZ/ptgWhk8
5+kBfl/jqOHmn0l3uB4twaJtbN5EN4pXoKvVL2bkOwZ9ipPooKmSom4RH5LbuhtF
CgjvvrFxwDjSPlpGthFcXo3Kkf+YRLAx66tTpGF9Gc66FU1P1uqwnVjQSBYiMMAP
/uwZ5NQ+DjHaJNTkyl6UoIEcfxWR7WukLFPkXE2SgT/EcAh3QBMbPDXweQP6qerA
sfTuYv0coMNGFDGpCvk+JElxCkTXAEXuSCDNZ3FuNbYTE0aWRE1yElrFnGJZ4b2r
Iyv6DgHNEAOmwo2uuL5afqSVg7eWOlo2+ZnX+uJ8Zz+Lh8yU+RW8+iAY5RvY0UHh
GYvZ3yx8BF+qyPupSGe5KhmCDCxVPVifpMKfwb+OYbopVBD6uzNZNzaGtf37ZYBv
UfamVY5bJRqNqjQMH6HcOzT3IaHxVX1QBIGVT5e5HV+Hr3gBuBQvMGMFw4KimayU
CxKCU+elVPBkxwMx92/DZhz8nNuLTz19gMMXnOGTTy5g7rZJS8JAFsKcIYarF/n8
frx/NRQS3PehPaX4Xnveh3jZgNI+DaVJLuvwJYrogPWSKhhOo8O3DX8bUSnMkFMY
iSS3gcYTioUK4aNXrV+W89rYPACQEirwsHR6K32Brne4eqLkaZBw62ii8jFNecsD
vEkqdCyBST2HH94CCKaLBFs8KsgLd2fQifCJrEvz0oWl1RrsqgiXl1tPIH3i5QVC
rC1Ighskjp1lS0kRNL4rhqbMg1gRM+im99InjQD4Pia2VNuv+h6gdt9pGtdZkvD8
X7HPC3TKHgC419IDNkpW1dFyBGzyjR87Zi0CQGXPc4/k4g6BoJTjajjvMY79ciay
nVfQ000wU/n8fqK5nAPweX7FRz9TYoJG90JCmcBq7UCA/iaa9fIK2z/M6bvm7h2V
28/eLj1WQSGyRIkUek+lEFYpHYlTLk8/dnfO+NweIvFjScGLfottA2uRj8HiLJzA
bePrkmm+KkIBDZrAXAyysbGqmnpFQlist5LUc69uN8IWOVL4pRCO2wcaytOIhV25
u+WjAO0WMMJ87AKz4ERtIS0zIcaYN0JFQsALTa1lglt6aLRc1IQ4lDuwU1upGpPu
ChMP0yfdtV7Ma7cGo8TvVvL3GK2G50U9mFSk+xS9YIjHrmesCgRXwipI4lFrQeNk
A/PBQqxb1ik2inWv7JyUrRLM4uJK5pUOpj7gzahQj4NU9VdBs+UcoOXryf1RHhJ7
zI/sR42kMlhkenrb0eVr3RXKrFTOeRAzeeBRacvI5Hg3unOeCXroEoYWWgq5kPso
Clkvh1v8LTjvqJliQMF+6OrS5EYfCRDRscE1BcdutCP905AgBfVfEdm8pjjm8j2v
qSeT/xBJ7L0BrLdC8biQbGKlrMAwafbLr8bDKZAO/0HaWJJQO0z29qukoNtEhenS
orydcus6woxg/MPeAfBHwCy3H3xHqmIsnKutB7xdVMCYbezncrzH56rF7j6qdl6k
1OUuAs0vS6Abn+p4NAAwbkvzIC8NJLfaI8VOFv6DOrhPP1b3qceT6dKhx/Zv8hHr
knZ3frfB4LuSwr4FG8lr+7qAS7HtksuVa1wMmv6y5iEynrPijn1vQtTBLHvjvQrj
6gf+yFvouqh8DGi3AtiWaFMpMWQuhxw85FmVApCVGXe6K7vN+UozoX4FdkGciW2s
OUeTw3LA3LI2Oq1Oww/CQXgb+XFt2r9oU6uu0qPn8pXNqHQJuYWqe9DzY7P/6l6W
/szgg0ScmSwlngacFH6twkBC8zRqKSYxEb1+QliiC57XX+Hz5Dh8E9w51utBrghy
nlykAVytmgcYN+lpSZ0k46w8zpIaO4W/WgLfFcxFy6i5GwOZq6TybRQrdEW9X2fR
TwdiVROMDvPZDYV0QJPacnyWmJrjH0NY8jGwq+4edVWzgtjo6CAP7u/FhIQtRacQ
FRvodTl3dd7Q9C9GeLbowDUfim6GxzgudK25mmat+KLiZYgAX8n53YFG0+WiYVHI
UDsXskODfbWQ4a51PAf2+w84A5NS79INXrxoYLPOT5bmqQOyXulK3YFaped9m+b5
LC68Ps4bCUnRx3C69WYxwqXTYF8MCSn3uvaZ/lcmMLU0KbStcPJmpK+YGoKXOW9v
UYinR4sGoLyM5wIS4JCGb6ADfnhoMeAiLXmB/WfNTXEHNl1vwcsXMWcRRB6MgMbQ
2GWOxIqeV57jGjuvuENXz/zAmlEDFXqpUG0jsgeTAqXmwmVXXM0I3JXniPioRZRJ
uySdmsHYDE1oK2WTIsz37Ucu6KJFSyXmRN2aSR9Ib7xGy/f9EQEpWy3/6lYdUdAA
Z3KHF9WgOozkqL9oOPrXnwpN3rRz0mltjILlqKd0iUPaYNLEwvncjT2qpKvfdp/T
UOVsMm7O9VQ0+7Zb7ZWtb8MSo0/xozWmD19ClVdtLHkW2BxnANNHEYomlUwre05F
4ZrFhLRrPCwDiSS3Rud17QYKHrgpcZxECkTu4UuNFFWcDkz6x75mf5XDhdPCG65h
eDFm6AQQlL7PYKXxXAqPP8NcQprkAt7yaNtPcqQYfgxRk4KJAWFBRnDvZ0t6ZJCj
7q0t20X5ZV7wouHSviEHzwoqVsUSFP3NfWbrnF9Ev9DTGSBiJla4t3/8YHzGsWcS
y8SQev4K4WRqsEWUWqAbAVfl+b4CNNxcq+hdtBjAC1dUQQMP1jgSwJqKX7TlpmJ+
AEfPG1+DqRmFH3d/mj/Gk6rkAQvJUwO4gqmbP7w0ydQ3cIeAa6TgJPYN8zNvFZ8I
nNtw2tmPoQIzs5EY8+HoztLp26eXR6NHybIp+mkpuCWXYQ9QMe8Z1+++pRh6ruVu
nvN3wE0sFSp19VEtRPwmi3Xev0CKTiyRTGilNxWd5sjuqPHrJFCKo9O7Rm2sO6L9
lc6XN6c/Q0JTTsXnEtpM8g==
`protect END_PROTECTED
