`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
igH4DeGPuBINe8dbhw7boMAFCld4Ikh8WeZjw5580jHBRMhqT923PDtR29cq7a4m
Oeb6OA0Y+hSFnUWNOEJs72PiK+t6SuwfO7i2EPtRZEaJNi/hhq6+UGqAXN4YIaiV
zYpOFzKInx2njHL4NSXWEJj8oLJk1rpBWYgpeTlCELaBNF1HeyOuYKcoh+u1mekA
sQSA/EWp8Z7ZwcCijaKpJZjC/AjTKZqlAE+v3Q2T2Q66m7xtoAjmPzMtMSqXcaaS
SWofMEzpwqc5XUg7dMVS/dw41krJBIZXGxYihsi+zy+a26+GaDDqfcp2PNcakGvk
N9Z/AcW7p36AzosuRtDCZBUIYS6smbH9BMdPGGy9Ll350DjFac+0DS29EmC+pCUo
/x4acMml73/bgQ3Fm5aPI32B+VAxc5MD7ZXehD4XSMLKPPPFE/w45I8zK6+kBfwZ
7GRYV2AvQrcT7RmmReqxDiXOaCNuw7i2SFqcCISw1Ljp1YIqoyUST5CiWWLdvhhg
S2MRGBTQ8ype0mr1UqL13/SqBKE3SPkzJyuyir9cgymKGiMRz118RNBR1izbhsmo
G/2bVpqrx97sGeC7hgxtMUGy/EUH81vwVmOSKF9MvKFuqj2sHNkTsu1U0+uLcLns
cdxWWhepCDQUd9b1MKrIKQ==
`protect END_PROTECTED
