`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sopiD58685FjY2Lrp8LlqOKwD1lw5WhDGBJeopV/Saj9tNcYFMV6f92HNQ101oFe
NyjPx+sCotVz/7I/2jnvSgtM21OJYP2rkZm51w5EvXSMEXFJmTGEUvJ5zWKqu70n
sHKtpvRX4+09rQh94LoR5kRZ7nrZeUDMGigUiP1Y/Nyd7a6JFcrZj0zGoHD+j4KK
cGDLtAPKLbnnNUuLKQu8ER3MheiDId+FU9O6W5VUtTQZ0U4G8QuBw7RGuEss16K5
Q3yCEzEkSpuhS2+OC4k5XY0SnHeVGnQ++KqhpMbRLtniy4NbbUeanSj0/Leic0WG
ASJZAlR7QyRFGg0sN04ldCuly0/BBhKVWlIDyfTfEdM=
`protect END_PROTECTED
