`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BijhpE7TUCFQJBmhRPgv9JZWILClnpMXq+3CQjsIyyF1rpn1JGQQjv2gX7Fuefif
OfSU5zddajMiLKkqsgSBoB2ZBxlFpaxKopvYwL+kzL/HlJNm99qwpxcogUN7eT/9
NOFI9Oed+JA44cwj64bHG3PcFTKiNB9jABKm47p0OyAEjg6jcAhcxhJS0hPXbp24
UXESiw7C1ExXxW27TtuWodOE4YoDLpsQc3VNvkVM05jhwvixv1Bmvs19HtuthMe/
3qNgcA8G9i1PIzOo5lUsqLCkDtGU0pjzKX8k9B0mkHvDCZya+cdgsID1hbfIA25O
aesM34ZTdLhoY38niNo/0j9BqR4Fridvgz1fq0UqfvbxDz/02CVMOf9GE5kArC9f
8rhA5huIvueqRPELCT46LClbmRB8FB/H7xFMfpGiDajjE6qUfN6jDCSAyRs3z5bF
z88pOrpxG9jz45A5oShDgCzEVCwUHbRm1nGonDjqHzQ1/MYMEfN270gSyHurxEDv
Ui/GbfyqqHNj3pt5VhaY1HNcdRfBUelHtC1okrFzz7IZh/84oe9Fk/5eg7nVVc4E
OS/gd3J2+IaM0EDE8FAryQk8ZADexhHmxS/2yCaS/MHjfrQhNs5MA9OArAipj4oe
15WRo+KJ546S3DTW+vMNf/AaxFkZ1xsobGE5VTd800BILU/Vk3izXqTf1TYyOX46
1BMiFpxyWCarHIQn5uXCDfv1o7MKdI2P/HCssBfQh1rbrR3i5moKeIOud3Ltz9IF
ZgUSH/df+TvnTYeMF3/6JNVtYrIyy2qhk6XSDSOxxUwlfLFFIn/Vxpk3Affo56ef
hPi2RbSRlJHO26xdAZnkNA==
`protect END_PROTECTED
