`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGVkSHrAPftKgkMXywfKe8pKfhVJ6n7qlKtyeeCZlhaK4oFaHiCgTWp2/4L7Klyo
iQhQhAln5uvvl9jkqsGo7ewF3vjpQfXlrexb3eu8+uWD3MKGNUm4ogRzMZi4h/nS
WKFhfzt9dXtsG8YQ9G9iV78e9Rimq5uPQucvBZM3akEcdhhQ1FsEHnPmb6dAeU+z
EMHawcXj4yia0AVxBaQifcwIa18m8mjTg3YsNXC5h00Z0t3AtSfe7T13hJ0YEZJV
jLMEPsBR22t0LHDb9Oe4/w==
`protect END_PROTECTED
