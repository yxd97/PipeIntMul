`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9JIHAQrI/U9NMIGM09lKEfXseWrfRWJmilplaYWrTt4wZeVc4hSEykupkFuzdN+C
5H3vs96HX4Dpwn/KmO2jO7eNsvbFFYaIHk/9JLTydViCkkaRQL32lYn15FolQFBk
FmW5wtmCoGM6cdR1BcDjuyeyw8EVs14nFcpAkY6kys9USBDa7hUVlsJDtt8eXwzz
9JOc2PvkhvqGIyXmxGp3wkrVzo9loUJHDSjgzQulZtVeKtZJd72ZSgn7yzOHXXaM
h90jO/ucn+170v6H5A2scV4JrFEI+VBUaiQo7anjgfFC0Lyt8zTam4DIXQ3tr8OT
G+bvC3CdwXOwWV35oWIKeo0Ak+w5q0EpX39gzV35mD1lrosvsmVMGOzwUsSas0U9
SeAAcoFPpcLkINHgdr/JXtJq8ebbmZxTuT8ZYtWVcFFqjX69LDx1Kgahzfq8YALi
ZKflXYW86t/PT+p4u6gMOx0CgjPGyRZyUswIz55IgKzfTYrUy1AX1BpxpqwLntrs
UKMhz1KkwhBVTMfAyhujMA==
`protect END_PROTECTED
