`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJj3oigjSeTMXV7q0+LuREreCosYyrcxD78KhWmaZ4M28PSBykmcgkSf1yKZvIib
/9MxANmPB4r/M/Y8RZ0TvTexaSbWNx1YeehnNwpXeZGMEiONR/1Pn9q1L7g01pzc
7R10qnQdz+2ACxbzqhyDjijijAdRzzsjpSukVOKgBVpZxR5QYaWJ9oBE3CgaSXJA
oWYpLItQoAaOeQCOUBgX6vY/IKY6N6EoF8VWDKcbpQU83bU+5Di8JXcOfIswu0wW
FWiFsKBe4lbQNor9+1fTKqv89gyqIKcn+8s1RU13s3w/NnQnbDmpWoEnko+oZl3C
bKOBEcObNGwvj2bhgXeGh18sRlMrrI9eYHRdF2lp75dmQDJh7Q/0gWM1+OOjH6jr
KzvzFKkJLZqBPNMvnfX3sX11B7wMBOCgybnX4svIWwDyKsNinT0sklb8IGeFIFyR
77Q26DZhCq0+7lAH633kVhPMi2Bb4Ryg5s3pjjvWMpnwMHQ/jERmss8pLJTEMtNt
S+aV4Te818wIGS4hnnjh7RDMY1P9E4MXonictBlZDEMde06HpLy0XflrEUIswPru
feO1GomRIcbMSl1+QPiOZi8O39x0XAEuSbXhDV7IXKqLluqHEVmVYEq5T2oJXgRx
Rc1G2Zj+1FdNExMd9NAtMouZVCLSMZl9uki28n9EFlc9khdiha5E1n/0cc4duv4b
A8sR2ahi0JVmoL2YpOp5eRM2G+nHIytdNNHs16vFqkvrVPW1c91Q7/3cRZIWk6oR
fgogOv5KPFipRtc+FsJSQA0n2oA2xMuBPDRyRkQErZ2ze6xoXl1hwEEKC7emE4aK
yHE5SnFWIUBY5XEBfEh6NJ/io715xzTQpWLBUthhop9y5l2zFJypK+PB4dNJGHSr
q1eEcczm25/HBdzGrTtbCcia12q5ncXFG79icHkxIgPCoCA8n8w+paMlcb2qf9wt
J8G7L4h0GTCnlIbssn1wTbBx1RHyQKDzEWPV3to3hSC1ypSUeyjJYWKGU4ObfPMg
UkO8IUb+cDpH2fUq1tF1vA==
`protect END_PROTECTED
