`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XHE+JsbB8VipukWnf5MoRUMQpOFRexuUM8NTA+sKo5yoH2cpgmOMjSDiXOXQ8P0O
D3nXwOsmRGKZUbNW0l31stzIyAfal0wzIjBGBG/DsrJ7LM9sMgA3HLzrQRvj86oY
QYrJhMuNzxzjile8t6CpqCHHKifmAZT5JjQZQprhB9CrGAZ3Gmk7OzBIMzTcTNEk
B3+psusCrWR5rFf7WHjCHsFgbg7Gc25PQR5UKjwrA59ylGmJ3hdtrdtCgAfo88Mc
H0h9zm43oRic1jvP6o8geP8/frqaTBx1UxM/G5egEw6ODwNLIllGYFvw5okcm/pr
cJbFsBXt+n3uHScNNwn7dKRnzThLl3dHFK0mSVjq6xn30TCUWONan3nwieoDScBc
7UaTvMFtLEtNZlQIkNbT202480eJSCa2VcXaJz8boFUG+xPKqvTUEnVMDg1TvfD4
`protect END_PROTECTED
