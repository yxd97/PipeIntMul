`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ENCOrEFnxdTNivqjeNPJxF96ykhbDnyZQwG8bDZyI6DP2kb9KT5fhlyJxDbNUmv
ZpMTVdF7by9125iEVOb3Eek9wcJxupJ3BPm4sRFfhd/RMfFedgBNpjBqBJ0ySXQe
r9EQjmIXlz/tWvgy+b9wmfDKSi08MeJKXZClRcDyU9VbJE4Iy5EjvB2k6tTlo4zx
Zaj8yPZrcHEXrUKcVnxf/gOPFbRAnJSaYUHmwwUdwXSFCuafQScqvveXT3P7IzM1
uLwx3DxCifNXWi0IXlmAEPJHGJUrli0KCErtm31AImvTgtd7libzEYkoZBh+qjrv
H99YETpc3HJjHU4Gre7kaB0Q4dr2VyQEelh1CNLGDk0iet5nOKLWOl8AomYy2Ei4
WrA028rK2zm6dmEY0ZzvFvVIc78Yz81zep6rmxgeHIhwZHCGPmv1OxR2fquBLz6D
`protect END_PROTECTED
