`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQcc53yEPc1KHvOTdbqdjkGHBbdV+oTZap/Pa0et8IkWeXce4Qs78nCDEgFg5kAp
Fc9dOUTuviBwPynB8FUUWh0oCG4zOyYLnSI+cDu2i0lzedUSL60AHxK3oUEactU1
B/hp6aVmS4nmPOk3Z4Jz+BUpSNmseMvUkIk9JH/YEcPWhENMyVFezZIjcJrd7hqQ
iz3bNZw9pLDp7BsaIJEPpAkn5kUD2WCDEYYMqQUUKWf3iQ2Gn4H22Pj492l8uT+E
jZ5svIDEPWyQrUvf78d33Ro1WqRZTs5hS/Efr4uw9HY=
`protect END_PROTECTED
