`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UsEPpmN2OMVHt7dul4iT6wWekU0KuREG5xpmMwoOIdsBcMoz35Olzyt35LYrtvoN
fetBpfeG09E22juOQ0a5IgDeRgQd8Z/NCKeFgEnTGaN4KfMTYRyn9EbXboPJEATs
BJ3OVHvMWD108VPNwJjxy/aZ6bp6odLVodRMq1V3Cd5PbDlOdvUR1qW7VBJXFyTx
iqjH7nHoPqCNv7kTRO5WjcYZbK6OdyrexqREXTQxGdwvk63PBmmA40uS8ArwibkO
Q+Ta+hEvfnBFOWNI8AMoYGKH5mG6M7WYC8fa7VCiU6JFeO2GzMr3HvoSOOSSrvSJ
PuUrEl8W5sRj8WDXiOujRHU5EzDV9psTz/pQ7+LAqyvJNuCFa1ekiEV2fXiByBQu
OyJO2g6EzZRXez5dmGoxDBkmz7Gf3xD2wnInCPI5sWd+rLkyaziCEnx1VN0UL63f
gjUPQj8DZl+eI570Ydg+jFU+m0AX4AMA40nNPj9lQ56ph7gSnIgriH4JqYtFo/aX
XvozMoCUIT40Ve8mhD/m2MVddtYFZArv0NffpKTsPX+QEOfKmIowXPR/8sEd/Ygk
mWlf62XgQQVbqDQ7oQa870kuheHh+BXV+PR1hGag9/SYOJqcn3njF9nBFns2p1GK
jo8HCU3ce4q5eEqcMsVvCPUvmnd9QFQel/x7QFXn88hrKzjhJuCHnGfFRwrOe9BE
pcOAh4DBn1yQyD2TNcCDqfSIQuLpzA8UINtxc5HWmLrGVadqESqo6BJscAm+YBaa
UUGykIXT5jXWAf3QmI9tEOVAJEr6kCFzj/RKbGsrDRwmBzFGb83vSzkdqEvkEFE5
MELDLxntl04HdQF/ZOl/3On2MR3SNx/H8Cs+nJAzesRat7WdfZ/uRR7tVwckXYqF
OPI5HM1Uo2Hp7cFj47W3JgPuxM/LcjdPG0hBRGQCb7mhAEfcPuFJ2YXvRxnV/Zfj
5OYGl4HQ5z2UwI+bvV7nTUJlMQYhM6YOtmUK+soEomx+VBcloq8Mc/kzCPzOZyai
SKpnZrcdWkNQMqV8JfEmOPh1jTFVuFq0ZPLZA5CmixYRNaUNoxO7DwGaTFNB+B2d
o1HffyTNbeSi7Pcriud9HeuX3diX1fxNfdO7HoqXVJbhIYFrreNIyRx98JzeEJRE
XXEHF/zcS84x+BFkjRzcHgfG8yPI6xGpFr8idsoMnQsALjM8dvi1QwAVUtW0SsiH
FI46qRn+SOvFffU2kUb6CBOY0HWXNOT0imw45p6a/gvLGXiJgs8NSS6bmOnFyNEX
nx1uDE3n7mYK2iQ0zyzL8pXugjNuk51yf3/zwiEdYXKj0OqFcg+wwMwLVkI4s+Jw
R0wyoZ3jK/yaj/rseyrXAqbyzYr5CduuQo1TbB6CJGHJzKRdWupxDWL/H8Qs1pJe
CmgbXNqOQXkwp9lzwH5CG5jB4XNiGO4Q8e5cqEXWEAAubGGluN158W8MK4g+tEKN
NnhAGyBPppIDvLbLqKQI3DNB6MPmDnwoIHECy4b8f8me2RqPDmyqCBTmEY17VvvB
wL5ysH8OOVPwCmIIEg2AFXFdixL4fKTybDKvtZ4Q817t/TlJ7a7ABWxVxq0jUhhe
wuf98LJa17AhL5AGURar05NGamF0K3lj2rgzDxmREcI=
`protect END_PROTECTED
