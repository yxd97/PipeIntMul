`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6f0WTvWOwUwVb8EtDXTmiyJXFA4tFct6Ycy2fMFYicOgIfJX7rZlHl5VIqMlJTd7
MH7NXX7v/iXn4h6dmcDmLJrppdcxLETZlgsSehYC4ZYwu5rK/MEh6wjmXt+UXt90
+LgiLSYbu1dUtxpNP3f5qnDhsqafyMwddKaUwyMzWEF74T7R8hVyX2bNrNzbvYHZ
J1hRJjrabga1QcEPPWs5puYh/dJ0vIUKBwETKm3Rrf+mBi2VMge6GDBbTTSilAcR
`protect END_PROTECTED
