library verilog;
use verilog.vl_types.all;
entity PLL_ADV is
    generic(
        BANDWIDTH       : string  := "OPTIMIZED";
        CLK_FEEDBACK    : string  := "CLKFBOUT";
        CLKFBOUT_DESKEW_ADJUST: string  := "NONE";
        CLKOUT0_DESKEW_ADJUST: string  := "NONE";
        CLKOUT1_DESKEW_ADJUST: string  := "NONE";
        CLKOUT2_DESKEW_ADJUST: string  := "NONE";
        CLKOUT3_DESKEW_ADJUST: string  := "NONE";
        CLKOUT4_DESKEW_ADJUST: string  := "NONE";
        CLKOUT5_DESKEW_ADJUST: string  := "NONE";
        CLKFBOUT_MULT   : integer := 1;
        CLKFBOUT_PHASE  : real    := 0.000000e+000;
        CLKIN1_PERIOD   : real    := 0.000000e+000;
        CLKIN2_PERIOD   : real    := 0.000000e+000;
        CLKOUT0_DIVIDE  : integer := 1;
        CLKOUT0_DUTY_CYCLE: real    := 5.000000e-001;
        CLKOUT0_PHASE   : real    := 0.000000e+000;
        CLKOUT1_DIVIDE  : integer := 1;
        CLKOUT1_DUTY_CYCLE: real    := 5.000000e-001;
        CLKOUT1_PHASE   : real    := 0.000000e+000;
        CLKOUT2_DIVIDE  : integer := 1;
        CLKOUT2_DUTY_CYCLE: real    := 5.000000e-001;
        CLKOUT2_PHASE   : real    := 0.000000e+000;
        CLKOUT3_DIVIDE  : integer := 1;
        CLKOUT3_DUTY_CYCLE: real    := 5.000000e-001;
        CLKOUT3_PHASE   : real    := 0.000000e+000;
        CLKOUT4_DIVIDE  : integer := 1;
        CLKOUT4_DUTY_CYCLE: real    := 5.000000e-001;
        CLKOUT4_PHASE   : real    := 0.000000e+000;
        CLKOUT5_DIVIDE  : integer := 1;
        CLKOUT5_DUTY_CYCLE: real    := 5.000000e-001;
        CLKOUT5_PHASE   : real    := 0.000000e+000;
        COMPENSATION    : string  := "SYSTEM_SYNCHRONOUS";
        DIVCLK_DIVIDE   : integer := 1;
        EN_REL          : string  := "FALSE";
        PLL_PMCD_MODE   : string  := "FALSE";
        REF_JITTER      : real    := 1.000000e-001;
        RESET_ON_LOSS_OF_LOCK: string  := "FALSE";
        RST_DEASSERT_CLK: string  := "CLKIN1";
        SIM_DEVICE      : string  := "VIRTEX5"
    );
    port(
        CLKFBDCM        : out    vl_logic;
        CLKFBOUT        : out    vl_logic;
        CLKOUT0         : out    vl_logic;
        CLKOUT1         : out    vl_logic;
        CLKOUT2         : out    vl_logic;
        CLKOUT3         : out    vl_logic;
        CLKOUT4         : out    vl_logic;
        CLKOUT5         : out    vl_logic;
        CLKOUTDCM0      : out    vl_logic;
        CLKOUTDCM1      : out    vl_logic;
        CLKOUTDCM2      : out    vl_logic;
        CLKOUTDCM3      : out    vl_logic;
        CLKOUTDCM4      : out    vl_logic;
        CLKOUTDCM5      : out    vl_logic;
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        LOCKED          : out    vl_logic;
        CLKFBIN         : in     vl_logic;
        CLKIN1          : in     vl_logic;
        CLKIN2          : in     vl_logic;
        CLKINSEL        : in     vl_logic;
        DADDR           : in     vl_logic_vector(4 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        REL             : in     vl_logic;
        RST             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BANDWIDTH : constant is 1;
    attribute mti_svvh_generic_type of CLK_FEEDBACK : constant is 1;
    attribute mti_svvh_generic_type of CLKFBOUT_DESKEW_ADJUST : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT0_DESKEW_ADJUST : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT1_DESKEW_ADJUST : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT2_DESKEW_ADJUST : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT3_DESKEW_ADJUST : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT4_DESKEW_ADJUST : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT5_DESKEW_ADJUST : constant is 1;
    attribute mti_svvh_generic_type of CLKFBOUT_MULT : constant is 2;
    attribute mti_svvh_generic_type of CLKFBOUT_PHASE : constant is 2;
    attribute mti_svvh_generic_type of CLKIN1_PERIOD : constant is 2;
    attribute mti_svvh_generic_type of CLKIN2_PERIOD : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT0_DIVIDE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT0_DUTY_CYCLE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT0_PHASE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT1_DIVIDE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT1_DUTY_CYCLE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT1_PHASE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT2_DIVIDE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT2_DUTY_CYCLE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT2_PHASE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT3_DIVIDE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT3_DUTY_CYCLE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT3_PHASE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT4_DIVIDE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT4_DUTY_CYCLE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT4_PHASE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT5_DIVIDE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT5_DUTY_CYCLE : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT5_PHASE : constant is 2;
    attribute mti_svvh_generic_type of COMPENSATION : constant is 1;
    attribute mti_svvh_generic_type of DIVCLK_DIVIDE : constant is 2;
    attribute mti_svvh_generic_type of EN_REL : constant is 1;
    attribute mti_svvh_generic_type of PLL_PMCD_MODE : constant is 1;
    attribute mti_svvh_generic_type of REF_JITTER : constant is 2;
    attribute mti_svvh_generic_type of RESET_ON_LOSS_OF_LOCK : constant is 1;
    attribute mti_svvh_generic_type of RST_DEASSERT_CLK : constant is 1;
    attribute mti_svvh_generic_type of SIM_DEVICE : constant is 1;
end PLL_ADV;
