`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y44vvl/C9jwCEO6FhqOv1DwMdc5PrAMQayT7jDn5kmZIHXiYDcPyc5dr5LzZA/zF
NbTV3Sygk2K+f7sjynckE0z1dvjlNtUUeuyIO86+ib27FLzTolKLYp7MfrGdS5ba
xA/rVpXzoXDzbON/q7yT2v3vN+a9aSaUm4qBDmxLhY1poUOAUfYGwGOF6NeX0oR9
DTIVvLhq1ki2VDMUb/iBfBZIRErJr6t9FXn0b2v0PtWKrxj3eP71eqcvQfr7iVQ9
53ZMbJRMMcftonv3zMZPqA==
`protect END_PROTECTED
