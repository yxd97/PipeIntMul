`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naFuc0+fZ2xy3L+F6VHUy9jOAwLOGUiNeSWl2lsBmgrvXt9TnktmnV5ZTa2flEnV
N/0/R+JMoL7s1H1Qc0EfPwQMCr6IZ3c99GotAhm6glJLwywScE+irjo4KGRZg8L4
Q1CHxgWhCgvyNgybCNiAjBGdaMp2IIyMKxAn5s3x7YuAWm+sDaR9+ScfAUH3Z0WX
1Fjql8+n8LLY/gxijfqLInQIOjCsR0BqVgiYm66jM+bm1tkvskfiLs6iDbfUisZZ
N3yFxqe3Vq15mbrbPw2xiljRH7UL8o8172kvp4GHTqdn8yZWNMaVWnaVJuQWoOca
sjM29QNUF4zjE5mo/IyfMhV+bWMGjuwXLAiEJ8KoBC2/zz125a2xGBwohWbildvc
52J9EVyRa+QgC6LdSdgPaDKiLyHwu1eqeoyO3omi3RjU0ZFtRmx6E3u1vqAnx/6+
YjoN3SzTf68ir3+pWDyF5BciVGdYpiPCpYmFjWE48CVM9qNVPwSx738Pu6n89ePF
WFld67oEGSJOKf5QVSOTfjOOFlXWxSp6xS6AVF50JijL6KyQGwnDTFNE8BYtCkkN
zwyjG1Gh3yTCrcodhjtMiQ==
`protect END_PROTECTED
