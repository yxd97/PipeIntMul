`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PFxUq9IaqHPLPxH9qbrV2PhcBMyl2b7Rxzp2am4szTtMVGpeiSpbduc2CrZSPDnj
6V2bLU8kWwmI9gBtQgtmEyZVIw+i9JOoRmAFqwxaQv3Y0BBUjJGfBU5fH6Kl2uPw
0DjuSIDNbJBpFDFgZIXdbZ5RGz4mKpZJn9O/rDQBNWcvOblGy0nxQAXbQeTeZ+Dg
Rx/fteJuLcoqxKUSkCQLVJUZz+/c0KWUq8G/JGjvgRtyhIj94Maw5CLsrZBQm5Jh
PsK094xoerKu394rBw4HD66n6stCi3BiQp84x6HHwooZBy08g2nj/Gm9pSqOEr/a
1DpILFJrCr5cOG3n6/MKt9B1VZx7aWzkqWKkEnULzek63Myimwot4zUYxC5Q6LGq
d46H0nVeBCf11b9wxO7sNwgFahTx1L0bmeCh0V/0LzeWK0kvHZl+s1edubkObTMs
ZEgA0BK85EZRXoZuXMuIAJsxHCd7XBM9cBW5dXUb3DnmVlvfUaf626N+Iqw0RWCN
CE+zoCg8SVGKoxh901vDoR/ThZqEMZbSrwog5UEj9gF7Ecqywak3DFvXHjkjalFD
V0V9zh02SpCCN45D859PliXhS/Gkmedd0IRF8K/30O3CakBpypfPLTuSAMmHqmGo
ovhDoE9zqk/4w+XKLh+K193vndGV5O11lOwkjcxiqGlpypKU8rMwejVhWP4VkVuL
XmPfBAEc4MbFntRIN2HE94Pnrf90EKd+mnNbsFBkr7KDc+Cf8CRMMnX+OjzLCXWA
XkK0ElpSHx9oberxJEpZo/cg1zmhgYqP9eTD+I6zvN/KmzvCwsxTrI0D0s+JqkDk
lKKsUvdgApG74bk8ydOe8NT5xc8wM7Fmh6IUBfJqhGGa1/NAZKy2wXdP0GflXp7w
mJ0NYlB1Cx+qNscQ5GR+R6HFYL/WAwSfhIEZn7rRT+sTUHLkYVAWHDHlM9vJTeCt
MqUYhLkXO6lyCsuR3AOc7eLvIL85bwvWWeegBbwH6fk8a+PtspLB8eqMwXwq3bM+
MaW/+REDsO640BEA4ME2rj/ah6E9n86O0IV3Z1Y0dX6OFXRPozpq9cNYDrU37HTl
pHY0LFSm0N+xviwlXwsjrUPPGMcI9rnaHlZTl0dpdayJGVIc93F7MlXXxjmkWpIn
P3uZBV9bXdeanyU+4CUv/SGSWG/dA+wSj9S9xypDAPsyl0XqFqyBnv1PFX/6+xDk
CmmKwhAQtz8EKZgFZemMmeWJTILhbvfWZwlA/MxOIT8=
`protect END_PROTECTED
