`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Wmnz+nE5tZOcMUWsGSLBm6Eu7hfjfnYvF899J7TDM504oHf7iS+KqhNnIY0E7NM
ZgFR66YZETxaseV3jPlLJMbaHaxHoiHO5VaASzHEG43gEg6S4hbYNXU3pZXLd8lR
Yz6jZXzPMdbu5jQeqVmFfXg/7j9D1gGoNlPQTB32ouHrKhnoLyLtp0Y6KImbGqlo
2Qk6V/femKXFnSIznyiANDsLWu80sN8360VtT2Q7k/wF/RRfK0nnIXYuD555uflO
gnt1iGYqAp/M+Ap3GAHWp8Qme0h6PWof3kkH9cEBexOjABJG58RAtDE7LXc8VDJT
e8h/XXddQwXsIdUsl/Qn8PDocwlra1sO0x0SQlOggSUKuddDjwGsj9wtqGm2dStU
0AoL4qGIBmE3WuHHGRbwwRZDYUkry5dANSdVCpIM+7RZjaUkSSvC6dJg8wBtIPIA
4VRwmVZwXkFOo+0Lx2gQKFIjjp3gLQpo1574mT7vGsP8NAzBEXCO82+xcGvgQz0e
VCiPEFI4w640xnHC79Fxn+I7ifUF3+G8oPZeT2zCOmJGC6R3Fcdm8S1tdZeeMrbq
0BhLmhWrO37HCULtm6R23PJNqZ+DEyGixGHXfpEpNYHZKgtZ04LkSDQrVERRoOf4
82hY3yUJRYfnkqXftYK6JP04pG/PPjwmMMtaSml+oZVk2+oZYPhmu4VeOLkAA0cL
azzOpQDkPrgZtOxg2paj+81mzIMg2H4CqDlV/RAtUZWXzx662rohrd8gDs1MRwXy
2pLLPA/S1ByfApIMqA+UKpXjzipLNwoj1M/pfL6B8mN+baLnoIpPS4FvD9hKRDs5
V/vHDePTbINrXddlnf+pdTvXtL0PXX9uHMjLraWCRkXmnIlwfi1oHCQmtsjCDaTt
G08IVFoza8SsRO8bhePWylBCGgqd3+TDKc3zd7qMpOqRfH+8dF1/qZepxg1SUp0E
fZx9YaTOg6JYZGvZJ9pOaE1LZFrkDH4j1rXmbpEyHMJZH1fBXNMxS5OHJjiNn4yQ
S+bYzd8WtjGY+kAK/dCRRXUpLB5/avWAXfOn81YwpkbLNKgbyFUqm5Lcnv3IECt/
PYiF9N4kyU7INQiiTY/ReSJwppCWezeSmS4LR/4hIizuezl/1G/JmK1wsgpzctij
AKndNHtBP75nBOgwKrfBJYb1J0nqS0e9brtMi00E2Z5jCTT0OSGfVrBDa3HoxzSB
RH0WaDPWu+vIxBV+2JpBl3WHWkOKHkthL03Hb4bjZc+ENQebTPttG1s58gl521AR
kjttQRYR9raOCswMnf3dwn2EAEqViv0Au+PqHdAwhCYqZL2dqLsMhrUhyhrDT5T+
Jl+nBasj4vZQx1ZBe5uWOXJOvAJeTv3st1vuqW5XKq8iy3tqTrrvc7QJio46lGNO
gkL1ASNzzKnSNMNSc3RGRtCYmWyFAxbK+JJGKd3ahGLtXHfA0lB5Np7K1LjSGDVD
VMGYBGK9noZvhyIe9sMOtzG4XuhSEqp/ObVd9dVKAlSOG3mG8lPvFHv8q/BlEepv
AQI05t2EESw6zcqAJgx19jKWjP6C3u4+O7PcBoi6h0ItsSn/yhw6QTeondqaN+FP
1hWYz2Lzf4O5LjsPI67bcZN/r/OFM683x4UqRFP85W+xiTWTKcU1OJ329JGjF38k
3kSKZbynFg+uPq97sPrRez2gj9huyxQ6cO43oWuS+NeoobTM370eMjztmyEt2eVv
2EKY3vvDh8dWVMDiPuKGrxOT5ztyPTpDMPBCuunnHHuBeB+Mk5HLIcwrYbFSB7Md
ZsyM9BrdWb3zRBekUiMu7zvlkBVlWA6cTUbu8/EhZFbt9mydXVAu7SoUjGNwanw+
cYWk1twMy+EF35SpXVMIpTtLEE7vZZEd8EPEGaLNL+AdZNLTUZTbzFknPlXjOUKA
gmfQfk5zHO675dxT9iRpT9Kl0WbG5e8X31+3lCWDV+3x5ZvFl7wAaL0J4aCD+4iW
Lca/4JNeDnBJHchHsSlcVz4a/4KU2PGeJyykk2G1RAd7OXCFHjH3WN8nud1ivOMr
d3h5rD4QaUX/127H4FWE5wSXTkpqT86rheHq8OazJCMjxZCg+v8PBPLCcscCQHZV
fHtwSFQm97b0AhMBcx6yUj7J/CpnEsy+1hCQ6QBLxEuL7x6AOaDyZyMLTXk6twfX
F+takELoYIo0JhsguFTTVJfKGAs+bMoEcRXnc/0OBD/nUGic/B22RdvBDT0RwgDK
ww1uqnwaN/0+bb+Tpfeur7zakkhmJELbf7wMghAjxS+m1Yv0+rXmPyBtTq2na2YM
xDC2MusMwPv3cDZQ4TUublzbhPpwyg44Ova/GcMQ49cz2PVn7ets/xOvmy41LnBp
b2hh+8YjeYPLxndvaipcXVCp8XUpgZQ4KCTUOndtEPsYLyghvtNqU8f5bJP4vwUL
HMzf0Bz8Mu+6grQ4MWKhqJz6Kmxbfu0N0o0qnkVu/jOQUvGEEDy42wlt47W7FaXR
DqE7HjnQ/al9GOJTn2Q58+OiA6E4nH0Tj3wlm3ekXMrNuFCOnGpsj1BZDw3JFJOt
i5SbiYLQppl1ie/jG8tTV0DQBwO82NfBolAvmQrWD/Qukgs+0J+ioa8RuQ7LazO4
/aQomE8R/lT/CCBvtKr/zyhYhx7Xvi+xHDHMHAjNbrNBanIl2ybJxmuSNiJG7rCU
M6F5lq2vCZ0f4Tahbp9spGOPMYR1jGcyUqDmsjfY2pY3uvP0nixfLRXR/MVHAmoM
4dn4DFpjdJShtjycIxZgR3j34WiOiYiCXedhSR1zNT5mXZH3hwR1g6V3AOu7mjgt
YZ2Zn+JxnU/Oz1F/LMP0pgzcxXfD4e9S7ksp3zB1kS0Hksq6/iuDXoiFcc2bimC/
5R64fSp0iu+NZzx+pOmrcTG4s5hqNIbBKbyLqY3+ZHp0iLvcYHmSkjxMd2OqBIPq
cqPChp5ltQyV9NPjUeHztbw/xQLBAjRO9BLxtW6FGIsweQmerlBKumdLFyn76bwf
V3ONN2M+lxs4tZd7l7Ogi02ZdP3Rdx8FWDUBUhNkflW7ePSZ3JkjGb/jO/bN+PA+
EYJ/VYw4Dq0lXxmUc/3+XSwXdfUaVoEcDJEq1aCC5bpIlyFlU7N+rN+yNNyvwoeP
IGhZ246o6MfY6uPXqfJhP8mLcSQzybFvWKZYcx8SVVxhZWP0i8mfLehhIxgOUHPm
NslXR+h3MgJPmQf0wHV6mB7H6AGrCXEXVBycTag2TTebDY+krRgXEKJK9lN1fk2L
pSl8E+s732xHhBpNbrx8tVVypbeO8+cPL7rd1LAVRym7Sll9mYtHB5inDKn5SeOj
WhIu0lgNsCNoGL7c2FfwUY07LuthCjdX2z+4g7boXLEVE/OaI12dCWCHvGy97rtn
1JyXhc8U+lXUT1HyYd1CX9WV72myR2nnnw+6D0Cr2P8OvjZywYW+a+wcRnM7H28s
XGEjtU92xnAkhRfeqgE1Wro740IEA0snVzrIHHtuuGFQMktT/pXK1jAP68D6i4T6
TTSphMPeM1rR5BIVMJWfkiQtrAr/GKmmWBatYHa0z5uJzI0+4UDhcLcIM9FuYt3q
9WCJJRYMAE75Ui3OT8/csRLdFwEy3tzEQF2M7FqnNxB4zXKnA6M/JwgSknHPBFqs
gl5pTYeXY2VXNBqX1Ts9CfrKvn0rO5J2PkovOcemFU79QUlXHzwvvfmAydFT56ot
iQTOEt4MsFHIzbs6tGV/MGBbPTVE416rKnt5Jw/w35ySeLpz2X7d2noSx3w2abYm
VqrzHOSWBPifCT40dhl34upFxADxvWBN5HDrcZdL5//M1e8evECh2U2nZXb0aZc/
YUNKYr2zQbA7eUmm3d80wk++69dWDkJBzfRSZT/nDlcntLQH2eDFbZcgFTNcIAZh
iay7r7l/QRee1OiOKEbd8sfgpP7SaMFNpXT1An95UkRaYEeJklvvHlUhVNzeL1s/
IEbxvPULdVZu9TFCdQY2DVyxYm6PgIZ59lDEPEIsEgwPO6GbqCKhfoYAzG9PUwgW
Z9B1f3/RuEN8dJ6w+wUiFMgc0pIibSW2KbtawszfCc29h1Y9C1twCaTJh0Yi9xnS
6mtQmvuWXEd+Z8sCAOcyRaO42F2XYLMel0TgCU/Tn34Uk/1Nhh/ntlDUiSE6sy/U
O98Ifzd1qk/yGF1iN5GjldXEG4eBlZ0scFeTf7WwwwPJJdVfYqhrpApz/IRfrNsB
sHIWlsz72nYPT5bcvqhcimny7rYAzbsxMck61s8/bCCV1VZmtGbDbOLawBawDUgo
wbX/33uPHMgnodHBlMOVn89DgWamRiOBodhRs8crpkyTFFak/GT5cN5QdwsWsC9V
nC8wJBQIfkIzRIqjlbCmn6x0URDBB+t+H5Sw7mQ1mfCNB64AtHp/HYZk1mlhqBF4
b6KBkCENf+jmzYekvdFlPSKsT1Iu8/UCNM5xsw3VRq4=
`protect END_PROTECTED
