`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+rKJwDk/YgZGnzMjjxzNvLFDi4VPeJOh+XunBVp6JehpjyBh7Qyt88eDn0Ude7E
IbFuY5tuJ1m8AbBCXIddmE6loayr1qYF6kSJZlvEQmoA9ZNnDWbdmypmC5xCKOXD
JZE/7q4WEMgqxrbFON9GUVRqgpE4qI+M6Q+k3cVj/9Sab8yZaY5sLAVpmTz2N3mo
fRQQo7x+PxegiTVWAxiRFoyfSX3nNBwZwq+K3eksRipqFmSuNg56XO4MA0Uwzqgm
TExY6s7LWBJtAxnxCNdGlhWmNSnXOES0cSyJQasi56PEbJF1TbBuIeNLoBwHP+Eq
9W7ZjTyDOJJKsmSBm79iCLMAckNfnwcHHETS8cwjNsmuJy+we/kGGjT4mbwNH0yO
oa2RjMx1+Cc3nJAh5CFFyoZjaFf6peiZF3XXqZB7/YbJwNyWUbEggxTtrObIsxsq
ppaAm8rg83U2ghIyHSVFq+71NsfL0rtplzRUBzyW4hnEgXNFwy5siUy70QS+PMvY
5ADcno0ogHCpZma3TrffP5wmXRHlHBNBQ+GftDaIiKocKu2+fU1fn0L4Cvi+oZqc
jUTJacDQbXIdmtCoKUc1UwkWtM9ZNx8QIev+H7RARZmPXXLUL/WBeHwDkTihf1LS
lObPsOv4vXcd2FNLtU9erum4aiE1nbUTq0hoxK8SbYTgOWE6kQoq43yjcjouvFJd
Vsx7qmTSPJJO6avjXA+q7KFEvNexusK3iIXjCN3J+x7KTIjBD8uyMeFeOn8Z8BY1
h643zGHNxbBIYx4sx0n0aL5Mf+zVygE7IOcqaz4JR0M/+4NQcvngb8hLdmVuLryj
9CuVZJIAEx8npf5gPM43do9mcJGjWmZexVU3lr0ZviLK36mnfYKiqbUMYtwAyL6Q
GN5rDY3vd3pHGGe4SltqfLSCJDOcu0wsPY5KqOdLuFBQHFxQXBmz39RldKYrRrlG
SlpAQUuQI8kYF6NMAmCizHyXnDdS7Fzb5aI1KiC38ZPX+TjfSIZy9PDLjoq95L+7
B2dmXrIxVM30vRnvh0iDQJ4BvG1wPHp2k+5u9RME4F1qOa8Bn6T+fPNC7xVzLsn9
P9CRTTENO6Tg42pw4USZWEn5OM8/rwqAm13AbiYXG6IEqKLW+6dr2ZYd4jyynzMR
af7KE65H5Yg063MS3v4ASgGjfqRXF+tO/3SG/nicgxlohnwojvWmyuyqQ3shZCcS
L74RA+GnAWqKyIrn+DWwU79RIW9fkiAkNxmM+l1VRQkkzTE5tP1xxGQPlTRXxeSj
UWkdWcF4ccOoVDPNnAzdOQpaYTrrEhv6rKslyoqezHd+eiwbUm9tgVjNcMFLg1R8
Ii3anzcWKt9UwRAgV4XfcpcgPEbEP6GytsNkSKZuRRC76uZTDl8n+21nyMPomVKy
B80+PpWGArEr23sYLq0kUbKlGv593FW++pXm7IF5ZgyAcfReXx7Lg3hbHHUskZdD
/zIdBDQgc0tTq4Fo2nXRJZyISXVnWHfONOwkNmqu33fYbsbUj8HzxRt1BFBPHMaK
BmXBDcpNxZwKQooBmHsi0J2ZAZiNXwhca/ziGLJS7T3KAccJdXNxfOWziPOo54JG
BVDbqDJDC+KKgjEk70UJmJ6HFvUpQJNNfyVGxVj46hd72XxKn+yo1glBABf9QUOG
pGU2jdGds+8OSqnHuBni/lWEOAeeIDsuoHKtxuPf2XT55XbXKx0BYRzgxOANJwlU
GU4sjFuOpUL4x3upGiaSg0oA8L2P+ldBJ9z9S9f08X3XTNDCJMeHmVz4I/9gjc7g
ivM1JrHT08EXZ3Y7CAldVXelGRISiR9sEpbZmzeunh+635zLCHB/UZMBle7A8Stq
Ie6HlN1B9UOEo2lWWLZnDPJ4hgfej7FB3Dl1CNWOQbV5ex8tYhSUMVj7/mXcUerX
Do31S9LZKvSZ6S+fD7MuNevom9FOFcPAWQwXdV8fGsf+ZgnwzeklxKnBXNQ1VjuX
0XKUVkDrQAF+F8W6A1Au7PPdqFiwpqs3hisQNnAx1B+rb9qKuSKDmbaK4a6XI068
GQ79/Y+fZWeFYZn0U5fD5xm4omoim/0C8b4ExrtR021E9F63ey6teDURklQzDw0n
HkWSyysFN+tMhWxEI6D9Y5MkyzUw1EaZSIAygfZAW92glXp9jivQS8yNnlmufdsj
x0unwENm6+dabY5PKUPMUSKT0y6SPljF/IMOVAx1peKhgLY3WMLBy5CwOq+Un9Hc
KE4JFkc9Iy7+PJ18RLFJ/Kls3t3MqIpnngwDTY11VN/5SKGXgqulcqFJpnxIThwo
RJBWRiacBAtRQVVwD7bORaV4GOMdm2KQM3xRiopwofaF8+0thLzVcp8e6MLtWLH4
rXvMs4D1yZUpQ5pge7s5nTS+40aAgz9mIxSbmMwhQcgztZan76Ews36NPwuGwd5X
0ry9ZeDIJFUlqzoZDxGpNIkqUMjtEbVu2U7rczvTQxX27rPz+Wcxpn/LkG541CxQ
sTd9Fr3vF7Np8eBEAVudK40hQxp5N3sTeGPBfZylbpMkOnqRiufGaS8DxyDM7Kvt
9JfK8ijqQ2RysI9bmfW+yZzYLM7CQSCHygaLgpx4v0L9XuboPAhtqw0J8oCgpT35
RAZKFLBjiikgN6oUzjW1LydeuRbxq4TXYl2H4Jg8DHh10j7J0ymvNFWpwHlhBFXY
bhkg9GrkCIqgqjAKXRRQLecopTLOYB+ZsU7ala1ok03MtLY/NxFPn8vxCFEL/+zW
Q1opCySlNU+bPLI+2Th1pTLJ2PQ6AQ/D3ogNaVAC55owOraHi0z6Ma+wpfrowu3m
pCJ6rrHgYCCkoFvzFx125gRWS0R5ZN0bW+TQjnLHnMviMeboXoQ41yn40/qO9lAY
GaAIZOGfQW0o2FloPBf4YQcc1JlNP3DpqnOQuurk3hJ8iS4FTpDFaJoIYUtk52Qy
0+Z2kFa2fP6AK53dGG9CnHLnxbYAFp60a5kGqLWbB+SWtSqPFSau5WEzb/Eo+tI3
Oo+XHPH9fwtzZbVI6SJC7Zfsz5a3qgmfoKf+7yml0r/hEwTqVZv/4cuV29YanVKC
8w+M6nz4SdgPyAIeZmU+ue54zf9r09y22Po47TwfbL9hDxyoGFpGNq0ATY38s6UE
gZvjc/MlhuiNx9kyIFBpS+t8+lfQVR85npuV8yb2Fsa7f+EBZvAkNYpwOsJNNy5Z
wNTJpfHjWZSky2jO6p+XEoAeO8LpIQSHOChbMRHRyCHGLsM5c790EVm006prSg6F
ai9X0Bja9Np1T4CVOlF+SYH6HpysFL3+X7BiSQJNhNEJlBXJfWEYNKEwGLNp96wb
Kk1/7khIe4pEMIgwLxsre464VKaB2eMOOOJ+yMisdbGw4OCje/rEkApGgDeOP7LN
kyMpUgM/8xygdxBQvDTf3wRb9cMoyYreOjNhJqhenA+UqCYOjrL48Bk+T0vGZAiV
N0zQtNMtk/nFefkxZJrMn8OnKW/9fESqEBgkO8GnaghvyNzMyfrtvm4SuJTWMCC2
k018hpC0lnGOv2OTs5sMtcZv2LYJukD4MgZnD0VpHpkh5wUMIjPyME0imigseBiQ
SOlH9iVS0BEyDJJEV8ESsqAkT4BmhNnIHNuhh6OC340nUgM63Bfyvr8NCPt3xSwb
J/vJ3l9/j59UcysUJs8lJuJyNDfCs597DSJx84j/0SIRrZdlV5SkTcwsxAktSiee
FMDoa3okp8RuMUSfNzB+gSNbtGI7XKo2nWMND4aMYH3MxhJ+CiejHJtW58Km9KMU
p9rk8dKB8jEHaw7ctlsPkFb0dY6qH+7NUzV7zwWovyYt1D2YhxdfGrx4UZ2oT9B3
HOjdrChNmOo9lZB1odnpsUkp5yYxbnCKBAIQHFjZ9iIZKylWiPqT4iYZ1YCBebBO
hW7tb6zNHHQnx1PlooRRnwqZIyMSBN2bzXS1C2c3R3m1X3G/hYhGRFNKTA+4oYkt
jT/7Rj1fYhOksyQxBUDfLhAg9yA3fJMulRxYtnObSWKdUEPtVw6fVDCF9RRcomJr
GiluHz8NkjH6ADLtXAAYSXaBHEGw9sNiurdtBwVkmO7k0Ui4SIq+b0A+sC8P+/1i
y7dl15W/fOhzq2ffPDETBRr7OOK/0JrijD5LFEWIB7Ua72DeD4ebMpR6Gcv/pvl5
01vX/vj/Qc0GuB4q4HLip/zQe82MPV5oc1O8EzO05UKYCY1dyoUoB/9EvwHhUSM9
96ls1dzPZPVq5ec37GYkO2uliTuzLkfPM0BNwPcCJarcn/IN4ImiVkO0ISjoM1vC
uBeRlJvNPK3rYIrhCtk5FtJvagql34pHJDUt97ZFziPalf0i1aDIa/kp424yauVC
uuR43JcF++NUENR9mUVKkC4etO9mV+eIADD5mZCKD+nNeoV5oFqIgPskcD4lFeV5
XTsCFm95NC1nj02a7JlRNm1kNaFBLGc2Tld9x1N6YY9Jvr1I2eoG0L4BJkWoaMTO
qwn+26qkTP8uXhrXBN7MVQ==
`protect END_PROTECTED
