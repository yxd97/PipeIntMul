`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mm9bpPi/ujmMQTNwGe9U56Bg/WlhpINdknLnUEXSwgXXrtpWn/maoAoa/9XD6D6D
XSdX9C5OriwFQKpnQCwFhREkrCUkgA1u0wob+qFXx7a/EEgXBZW75PtbF20cS3el
jnbxPXZJHHZQ3Y1cwIgdgKVq9fsCN+GOu0Gon4fL7dvwugNdLmaPf+kB8o7utGUn
lCIczL5q582PQmFEVa7GYUqICEOQUYtQKpyh83or3VWk4086cbTyQ6OwbibCbwg5
6c3V+NWXErk6YTzhq0r/ySMoiTIECjs46gT2klPy5shHcyEBERcZTVi8s4y93aua
eYBvNnVy2nrOiXCdWAWlBmI+6PL0wWgqsSdB3+BCkStMAPFxXuDWONO8nDroXgMC
p1qukugPNdHy5E3BoHsf0A==
`protect END_PROTECTED
