`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wpN2PA+uq1HrWigiwELoIs7X8X3+uPDGKaz+Wzzcj66JAkN8E2Iqgp7D1EcwQS8e
l1zvVhwCxO4Qibz+rFKD9MCq6M9sEcDpqxYL9Kq5BYlhuaNSQ15DYNdqBvel+T6f
/NYqfkgZGu08ekhYsdQJM/I+HZG00OV+lsA1OvoawAjRXAYAT1QqBDU5JdiHunFE
fsUlOl9ipBLo8UnvJjDkvf8wZce89HRji20c98HaARiI2LonJYAnwAzGcib13nPl
`protect END_PROTECTED
