`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/XgsA4jUV4E7oSWOY1nf0AKQaiDaljkErLp+sYrZQEuVjxHVj8xmymAl+eJKYdp
CTRGeFyEbzMZ9n2UhCz24ZIJCOdWYDyY9pwwYc8Euiy0DZkqtj2biNBNMY/rF5dy
04nK8vdS9BDvlz4rAkadOzWxmr+cRDCGyAGeJ7QAuFizZn7IRQPHvXKYm6/yTi7y
uoyQeEsx3f/EZc8veNwmQiYbux0KRH0pzHsAYbnFuDLw12JeYqGLu7i+KKPfFFnw
dmuIAhKXG7W3P94uBCaq3Z+csEMp35a1zRIF3C697tmIFIhO4ECc7kE5/xvgzP+I
mNK3FDkd66nl/TG5JMBPTFnhYc+zZT+tMjiPPU5dZSxZ5qPEtje9zwGVh05B9gEd
`protect END_PROTECTED
