`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n0PNrmNWGS9sPNjumk3gas5R73oQlCtmIyFO5/Q5yDN9vbAJ8MKXJbCqXesGY8cX
hFQnhDGujdOisJkqv9UjU2alVNzRv1Uus6NCtBZksmYfHskInsbLcTqk5jJkHIAJ
sI099w81mJ0YHigZ/CNGiOE2Ku/l+tKoK/geHWC9bl2TOKPfDO1VE+3XTZFg+O2S
2JD2pK0D7s6fg7QVXP+Uk0vuDVcz18iTi2cSqVJSgltgzYErfU0CChh2ZnYhvbxz
VpGXtob2d1bN6eFTvqO5i+vCeBfuoGhCMt+zt7nAHWI=
`protect END_PROTECTED
