`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/IyTW5HFfdcBUqk6zid+Ag6a3Juiq7EdOhpwEayRlieGtTvbszX031b3sQuSfZ+I
35za53BjDtvAbvB1YYssKdsS+BYM/V9wefemHvSYEcBjMba0nS6FfsLFiqITXwVG
x9y0kj2rKZU98oW1G9EDdc4N0toKKB9EIJd2ak0SXP/0u03AKXxetRz9F8hnuaTE
5PIDmEXd9V9ao47JiBJMoW1Z0fFEaMBZ9B7CExbdpE/RkWdzKa76IHLWnkRJtF7K
O/6buIGwMD2MMkhwRQocSH4jh58DWrojv7+z/1Lyg2U=
`protect END_PROTECTED
