`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXsvklBa89GLD65ydBUrmBK4LIVFcsYEOXkRD7W5n5Qr+8W1+U3oi/R6Hs304qab
NIOQKfPMlZhmEYHPO5GIEEXXC3y33mKAfwFse/UqOt/CkIpUGUP+xWuJ7VcDmqtu
UyCMse3ziAeVXbfmI4AQO4p1+/ldxu2gjWh3fu3kQRuJmuHoTHXgb8jsKnx0GPuT
YnrmWmwqsoO/GJu60J9tQGcVCT5EdLXGuSghnkh5SfT4d2dSlvJ+vH+OTf+sTFn7
GdX7ZB3GnI6PUkR0iel0Em2SiX7ITmsqpjDJdZFfI4654b3sKulCMQhp7KHiR6mW
1mgwOE5SGr90LmiH6lKtIhZnpdrTMvWA1PJLGqTshDA4OMCoSqLbdejw0GQk2i3y
7Cu39S6OxTKCPdCk5LsqxmAd8YuJR1G5Ao2xEP0oCxKNa6uYzGBdQKvbuBusz99q
C4alwGCM+QanuD+zTcEGXMUzAmZcW5LZ7eY3Vxv9otLc3wDvZ4gIUx1NwptVaSNM
cUPY3JM/41od77b6w/LXJEFVxyyObVZ05OyFA9eUN20PZ0RMLUwjyoWmLBAySz+v
dSesxL/aw3X9+x93OCEkAowwMAmWyMTUH7UEQmjmpia3BCupxgdFl1g7CfKz3td4
osmIGS09DQ6chJdn1daPzg==
`protect END_PROTECTED
