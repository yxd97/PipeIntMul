`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
48fOixvDKn2Yb+wHWK7/Obz6Z8vcR/BGAN0aZEkSGmQVKAWCmyfRwS8G/ikLNuF4
0Z528AD54UIYIR+ZmrPRWk45GonpkbFFLcuV4snyUu3xqANR8nhqSv3ooR8PWydF
t4U4tQi/lEva5ssFA7lzjrlS0BaT+fzd8d4Q8o1ll+43mEBEsn5vPrBdBBzTmZzn
yu7sJxk8w3pH0iHIDzX4rdYqty7GPUXmUQ43/qladEIdYf2ALeQNVVuwYJXD20cb
+uzUCLvWNeILg54S3N+3YKkAkuJHRxXrtf0VwMwUzi+CGDcUWeRvcOVMEMVFVjwx
m8WLS9Lnst25kxvVTBJQEv5IKki0oRlAWpjNQ2BrkmAa1vTr6c65n899AyuQ0Eh2
u16UTqAb8Md0tm1L/wj21/hG6DnIsIQR2EKeUssSojnpTSefKFy+PmrjrKs1c/xY
QGtfGZcz3hvsmZ/lGAu7oHomv+2wNKFJqjoCOLT2W+PvgJAW3ZYCKvGrzu6hNlCz
xNYPbqVSBQUcIDR3tagTEih7U6NEEsCEj7SOUrZnyIBOzhFqpb2xxKtRcbrdnAnk
u9uctsr9k8kgme0l6mPZW5i/9a4lsBmThMsw4n5PRSNFAOPeUpbzc1Alcc2BpSif
ZlBrcT7PJgNmYo0DLOXmSiGd99CyL8/46jHLHaUa4TovEfOqtMiIgwBubfs+IKBM
Zm1cRFJooV4nPoZagwVEhyi1Wfte6U21FFKOwqMgwTglP1BmNnOQ4jO0zU/t6nLV
ijHVAlV9Sk4qbXfnHaWz0vRwCQR6dLOZOJvWgs+PY6AuaZNPzV2M+Br6OaPxN5Le
U8Jsf+Cmfib5yQLXHxZu+RuKBillQuG+I647K6giJzdnSy+GgsCHd6CphrZfjc8z
PrkI0AfHaZz4hVYTdOr/BSR/kaFZj11hmsvCALCVW85pKbUpykgDXLtpohsM72gg
CAg8A5hV2+arBv+yTpC70+vNZEp0i/op71vMP37Nq+7Vog2Bme07mNqxX1G6XnGV
sQb9lhDZbTCpHqSInwv82StHbx9SwCWTe09YYgw4wKa+JStqbxyraRY8muuh9Pyv
NeIi9IEbL7sJq9mwBWU5wfxQ89b2d/YNgXC4qQyFBBiYkMwjod1pb6OItkZGvM3k
UKMM1b2uUfassUAZgUolwoZpMt+sIv35ric5YhCnJYc7jhUdzzLGgLcfWEmnFOnT
SJPuUw1lHcIHe/gOJedpXZG3CZ+7giQ5vVRuq7xObw0QRwwCibSkFsP43qqC4gS3
oGJT9r02pgBXAtVqmy0xh91f5ie8YIURqDvA+PV6AR96ltw0RGZTqtXRfMUnmX79
3vMmsXD/llnsasHjxTm862yaousQejJgEz5MNeD2vg+eS/heASVEavT1i/rf60GR
gn493T1niIzKxIqx1MMSeKni1PaqNh80O8rrZNRMoatXviSpYGGJdaZ+faajZ+bM
og/HP1s5eDjVoISbdqZAofe1XZl1Zb87sp2vMPAvoAgfNjQocE9WvvhHH39yjWKu
4KEQK0/0lcq1oX+X/CrnsDo2X7h6tRZQUzjxp8VD7LrT1bjvNaaRt+uK9sEFnTZT
jaouiCQvg0JSb97DScRL8KlEzU8ya1GrTQEY6t/i4qWK6cMZJE7JWUmrcUJx9y8+
gfdAMwo3WTeluuoRG8sxhmd4lv/mirvmU6KVXc2p93w3fuHCBx3WJ2OWuEf+A8RE
`protect END_PROTECTED
