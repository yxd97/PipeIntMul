`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ftkAsURVA39hzUkZrr71I5ZfFG2FnDWAkc3QZ4a1jMt4ILsIuUGZT/AN2xHl4hJn
sHRlQo4D5MlJLY0wPP/Sv2DvFxEAbWxDqFw8X2QdFlgybzTDFqIywZHpSEUGJ0Dx
VPE9QZYecqooUn3lptuTmvrzUhs3rGdUB1iLFFEbkthjkH0enaJFajtiY/d/F6PG
uBha8GGcaSEjW2vZFaiBBOx1IFrP6GcqXFAS08xURDHuF86b/tNgDSCplqiZs6/X
P9CBXirmuljP6y/RN3TuFECv5hj/ONiAwuuadNMgru726xiFN0b6e1dP3/ypM9bu
ADiuMqrLcoPQxPDkzj8FWDyc+Fwpl4bKba8h9eugzPV2Tk08VGzH7BA2gMuGSm0U
1Ly41Y0qPYMM2SAxDQT+pkftiRg0K+9SjFscmgn4y3s=
`protect END_PROTECTED
