`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hu+Ne2J6Fcr02I+w/KSaOCx0LDsRexMwPtjejRIIypcltLSQKjFPg4Afic2lSHID
Ls4Bg/Z11P3cWOkfYdPL+ROuCI4sl41mR+mujRAkvNSrKYIbbPfxM1xMQ9yBanB0
MFQe1m/ORq7OrnuQwYjW4PKM06vkOf+sa0yiC3mmfDzAgA3OODgz8lq58g34ZFww
VnJQTf69XJPAMDnB8jcRfa9abuS+WkRZYEpQI/MuBpgB/aogU9Tz/VDSA8K6LNiE
hnw0lXJEyz+d40nf76Jpa3HFIJxUd6zNJ/hGcXDRjnywIHQDad68FCqoNvIOEkCg
JRhcSy1qKMrsmzqo4ZuLSdhNvjjJ0CC6HZlvrUogKrVhMdlj072z68oXljMy0DUE
MD6bcxZ5t7irdev3DDh+ZsQwE6J+SIgnxfTCy3YN984tbfEHMLOeN9feVWaPZtox
IIr2394bspMWqvgKXF/1Ro1kOj70MtVB9SlHDV2M3Oe23Z8/+aanUcG3ZGuzWg4f
uDL8tg8a8/a//wlw2+t9r2NCsMADoG+8tlSm8v6EOCrU84idajwAj3HTRW/enZRR
KuVVKgrjf2BrXjKFtOx1USaWSysArkb6B4rpE3XtRoxrqGC1oPoOqEg55asc7QgC
9fDjLEM0v1+pE2l57TZqThMgAi+0H3zQOepIx2tUGRNoUMCrXIxN3cCaE6kjio/D
ZaKgPnfPU0PQC9LvJgkcPUfxrmUDugT1fexMlaJD2CCJZzUucLY4M0f2KAL5BTOa
+Q1dRtNir/anNmzPAczSMvzJA0RIsg6iHwwlGO7taX4PB6rFKrZbiaK1mbKVqbA5
ifvMbJtjrk/vzaAeWq8Z73JO8X8uKT+Kg2R5pa7WEcJE8jclc9hXSisHlSy2Dil1
1uz48pZaVZLpIUqudcpxAIjeE9HNJDloDWVNlIJH8MKoAmy+GtblSwksmylZSRP3
Tq3g7XFsMHKBbUTBbND8AZoGIevDG0OSMb64NHZBBx3/4R+jihxUNfw6/Pvsokt+
GYz50DRNrB1WVo+G2j2E0cdX6g3/rY/3J1AjYBemqNS/AHhwPMc/6mujDuLa7zdT
sbAsF/CkiPux4v+h3AMuYmBXRsqLrc43CKhjrZmqlOLdR+/j+WDjaRSrhXj5pM1h
BdPyQMQJd9Qk86Zu9S2fgcFMLNFMC6zLS+yI+aUO17kl6sQ4aOs+Ea0KNq8Nq2m6
2Db4Do+JWW8v/V5heBxTsK0LqRDygSm43pS/3vldiJ4Qj5N6GHqBwDLUxofO+1Hc
EIkXNyF1jKOn/sHHbNCkLg==
`protect END_PROTECTED
