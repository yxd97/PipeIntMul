`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ssom1Mhn4+DY5iyANWYBhtXjP6EnQxJf4FL0em2Skd7F3mz2eW0ThiGxCdUo0S5M
MgLUz4lJ02NoSFWJT7aD5lU+o/4SfrHf0Vo652go4FE70Q7B+RKNfuniUapkuBkw
UZshBcMkwkV0vdaD6w2tem0w2Z3LAFPri+I/dGaE+LXWKAy6mKgsTRY5mgyabwPo
89kDr0JEBWKkrYL1Vwad5JMkG4ffewNuqyt+eYnR6kxhIQbjkd37k8oXJuM+lORC
44H78fDm9hhJY6ha5STwzTU2iajyZ1+pzRis8G1RPA5YxtVgGjNo16ilbqPP8Zrk
vbTY3ayuZG84+2X0MXKAOyLXNzhmOhQvMyA9+QKFJMXpBityA2dr6XD7n79C+OWk
VfqZm/2vMgvmeqqwwJV7lNc8RxX+rksEeYvHTGlpP1brcNPJ3+PYF1OArzaw5l2D
eLfe24WQVefm7Zh606GXgWzmUojkUdwyRMzPbkeQj8Z7SC6vJDYbydzNgJbmnnRQ
gDDnEC+JavQIJTJQ/rVx8ntTi63EtSGQA+R55czUXiD3alwMA/A57HN/8TxJLnxf
12XVQc70HJqmlt8PB4Uvqm8h2i1qt8w9JXEKWIdnOqzNOsBQ9079cJ5bOAHZAuSR
DxnqK9NkZOUvpXOez3ReKtBfNOdj1yOBjr5f6k1EiU9s1bBY/zTU/TLc3xi/t35V
x90OiHagbMoJnIxVC9PCNfZARk8+mZ9TJ5RyxDoe31HST3+3nFsOorXdxUYZh9uU
nBA5EKVgUG8Vl1qqwal4BsxCXv4mYWOupWtYUytb79jbLE//LMlFCTp/uDYYMWYW
DwetGPn6N1DN1i0XgEA+0s6ujgAldxuK3hhIxGffGO7lFRvH58XcjFLUQd87xl15
hlGWm74HbIWFsduVPs//xJgUs4OEPJ0P+fUw5bhX0MM28X4wNkF4X02RSLH8vTcX
LJYl3rSs2m2CJBWGR6aosNFYr8PiOA6Z/t9QtegjQrQy2T9RM3suaiDfZtcXgXEc
QyH521c7jcHJJdlskpe+mt6S2LXu9WudQrLr9Wck4pbbVBLflPqnR5cthDafFSDl
7FjRiMBurRCF22mFublSgUvLJ33FTsy0BTg4Mxs3Dp+2NhJxMjfYO92zk4T+WrrC
SDIai3KiX2YeEGGy6SBn4T4y5Ud9adUBHgGwpbwFHbZ7C6X1eJlPnLQPnodBHPN/
el40uXhl8XFeatIWz4e/S8qCnlvE9ZxhLGTGjJC452vsm4rVbKiQ7amx9sDNFI4b
5v5+CeCdrltzwpCl0678lsShrQdz/4OdpZIldWXSE671lZzxOMxAaWhsLMtcyJOH
OmyYuUYMb6E0Yhfs95KVVIq3jy4yhaBUdi4y79xDJD134Uh/pclBYqdxaPmWDvM5
2b/q4knkShDmzlC1W75WPqu4zamj18ETE4fil0t5x/mEmpbBXpzSMcGGZ/Bu4yUn
FgR/ab9roga2AYvSmpawWcCKwDiUt1xslmArgDXVY4T95nKBD2VzDHL2NCcMCFnJ
NWZ44q21yS+FdBOQQqj79wxQaR1tCLYKa0bn2x/SPg329DgQNIxLol9Q6SP92+IZ
JLQQvEZ72XpOQ870D7F3mKXFBHQ1p68sOJFzFHnCxUbfblyp4UzI78EU4Cdgu/1k
qZqPRdeY3KZgb4CsDB2sNCEfxHA0Rpw2TjkUoZOqdgMNzwWWmCByWb290jiyhCej
nh5heBRbAO1lp0Jv3TNVsZcHaQmQ/lmlw6stnS4DBEwZ3exbqCqSBGl9SNCMTvOk
Iirma4Ub3eJbvJrtbCQcClZNbF4q+hua5PDZEbTbt+RXlo0IIawY/APLKBREQehz
aXxsAP3l/0pj0gLMHx8uMT2mRIaMgrQPWEjCpPSjz5+QMxs6DDXkWB++ASXAvh0h
uICnDPs3CYS/sUU1mZj6Jel9DRbk8FeS3m717C7T3wYMFVKSPAFKfCOK3YSI3h66
+MIR1TWOci/3DNnjzNKTsCyTVb0lr3xIQ4iBUQ949CcBgRMlb/uPGzduR/uCymjO
ipnmNNX3TrHBlfMAzgQtLyzqgYxmV0e2s7azcr2yMZ4=
`protect END_PROTECTED
