`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0JmQiieSUuDMdKJZSFTln6Wev18No/fOa1tv1WSPaP55zCPZhFLXK9NR8afo8lVZ
kOyZEq0c0l39LmoL7DKOCPypQYcyjYUz9zkH2ySVE/JSaeBCvr+eF8AOmF3g4YQ0
A+63yPO095g+TEbJ2YprTtvNccrrP4KpfpRp2fNzb8pxUrL88P9WzOtYwhY9WxSM
2mvKqIvjXf5tq7/d7c1lXE+HGbLxmXluWP4Jbx4+kKN8e5qL3/n4zsNtveBAmYJW
BS8EvO3KkIriu2lcZxpCmgAKbrop6/uynH9p70wUi+/NhHIuv9zLkvI53I+OCDax
YOxfPYu+aS6O9GTsHUzvFy3VyLKLAlp+Jy5Fl2Yf5Y3pQ+K+NSfSSYWbxY+Oj9vO
juG4FTrwnR2i09i22Yxrs3iYmAPz/ZV7wTh5Df9asPQZGShYZYiX3WVutT0ZpL+W
O4IFDB6PrjesNP/o9GRHw+Qrb3KyymuFXNHwu/eFlITmAxbVgXiQy/9M6PChr/MS
`protect END_PROTECTED
