`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TK4ZQBAq2qOQH73SLqb0NawIOkzo6DB9u9PFhpnfx+EHVmEIoKNkJiuj5zfeZZ+Q
6gdDaKJjmeQOOtAZ4gbvyis8x5zol6RyrGH+P6jmphseTfQWPLX4hHmETATljbF6
nEOhWohlGkfIPoslnsQXFFspj+WBf0NNi9PiYpaKy+3tLjS1lBvTeZ0ofsGzxWyW
iURzOEqIISuFUq/v/2UBwKsiZ9DlnMtbEhbMPGwOMesm7Dupy2k6C5B4mONpqY1N
5Hq0YhK4TKDhk+srGAk3v0AHGbcVCGn164tVU+vffZQhRtT2b+BZxtphnsSLDi5i
S7vFY0GLqYCI0lY3XNLt26JzLHwId2Hcq/3wiRnP2nJuXQ4AcaFP/dakMdvtBvRp
8PVbqhA0GzpMPM7Lr1vlqWi9TP0J+YsTGou0D5Szimz7YkGPqLQ32xp0IOR8cwwu
wgg4zPz5wOS86c3Yq8Jc0ynhP/MNtA2zYRf9Nhs5bDkluA1ie1QlZ8AtBzM0ZRSW
PiJ2tjOa7kLrIyD07hWaZ/BiSfSdN+tzqcqFY7sxjpcCfN0a+I5Dg1lY7E/TRShC
GOrMT9NkRVziOSfFlANWkw==
`protect END_PROTECTED
