`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uGsH169BsBA1/qDGmD3dZ+YBYTqkm/bDsovXOT9YBRrcCQlUU3xu7NAKXya0dY8
ZkVGxK9hfTaKAnBQQDMcOiq3y4AhFlmgWMTEIwTOvNIWJ9FMUhshdkdrGrfVnA3Q
6KWV9RgE/kPEDUvSBiGZOBnPzog8qgzwdYx28AlC20r76fKhLo//j0MxjPOtb54H
mCaOiOkF/MO96fEetygLcoyp/+IW2NwvqYE1Y/qmUi5XpwVD/0nCu+cQzFEOqlGq
Bdww958SJ47Im/l3tpjfv6m+ZlWpcO6AdX/AWviFlTP4oIrS++6lIed+eHFRER8z
n2NwpbViaQblfK7GGggFj9oFWVadx999QHOV2dECO69m3CNtk2t0B3kpIKZPrqT6
uxLvxyJCCOY2hecnWq5Bo6jX9SBoxyS8ZMVngARaT6aKiDfCAAnTdZrhztAnGXPZ
D4DXaQRk7hCEQo+Z43hD+Kv/kSyyolUoG79uSQzDpcqQ8au06dTuoHx1bTHkaXal
j05mrWwpZXhTrGZKAUsmavpXwbndsZe/I6sEIalTrkchKmTOJx1Rp7EuqrTD+CsC
rRRkBb2UxZcW4kjtXzvYYT7mhc6lNCsFnuwkjwBuL1RalMyT4g1QeJ31EoE1JUcv
ebnkck6ABSpkmQqiVnPynaQ7JTjYtwrf9ozyv2BYnCw=
`protect END_PROTECTED
