`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JZtImfq5I6gJMMK2bC/xQd23MDiIqznoXiT23FkmEDEL+kNAcWsPDawoqetww1G
QUiY/YXTgqQgfknILbM1wqlj3yPf1BAAr2g7q5SXPSEJnooDjf7gEoNpUeGG7Ny9
23fyn9U8Qj/VvxLCGPzivBYDJa95W/9NYR5fu4pKT0ElClTRP3FHJvsdIgvZSdwl
926Mg39W/k8IaHCTxUlwMQUeafSAgOKrJnEkV83xNMxEk9sZ5/RxwOxQpXVXQcuI
qMZNmC84iZ4U9BPddJctJThJEg89WB9oUaMhbq84WB16aiFJ4201Y/9S4zIpYgUt
D/v69Ms4Sy8Iaqh8QywK9ISN7P4j25VrBbG79ViKgP2NPYVD8F5JqR9BqA2ncA2s
lJ3LTINHdJDoi9y25sFqcqzS42+O3Fh8FTaj63n0Czg+R/7KhrcZEF+NHobY/rfI
UEXGNjYpJUACFCeXXNLlBksRvZArQ62ppZbqyvNPxxRM6fYryshXyb4LA6/8i3lq
EXTmuggFakEr+Q6jzt9Sg9BaeQDTi1eEBDOsGwEkfSYjJKX30iD3Ori+rOZ7cMrF
F7+mvhR1WqxUmfdS6bto3ktZYTQ9d7ZNBUW8paq5LMqsiI79mkGqPLS+dDoDPdzK
KHcEmL/eL5TLNzpgtI4Deg==
`protect END_PROTECTED
