`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
teSDt248L8o14tCnyogqgCM9+VJ7JaAmgWLGHKpCUU8Nc/3cjT8JPt0VtTg28gLF
CIm5dF4LMaYRSRGQibTBtSONQplML24Xte9JCiRvM5PClohsE3bP0/jo+7RoVLTb
AgqZA5OOaV6FMAk4im3rSW/y7C+9VSVAwCxYpaUbOB+3Xy+FubNofM4zy3IkEWP4
eiVAUdhRBzPMzu03v1qvelS77jDAxZpeSplGByZNu/OrWjNr+9mRUjzIEsFzQYJQ
zO22Q2G2zVTd76CF4J5t+ZsAhzEhYisFMykGitIa4eJV4k1Zx8bfioydwtBsPNBN
wWWeBvu9DI/+8BfQb2DW2jzD7MsAupjzHyAsU6IBkOFTWt3X05veUituYbpjyv00
iseIvysYaQhPDwsPyeGAReOgsd5Z4o7wiWpCqF4F2xvqpwjVmOOVvcjCvi35WpuE
SuZj0qMrjayh+2lKcmwecnLcJtuJHSWTMNgvisRjIbLADGUcsxnCtiky1xfyQDex
uyiftVdCLesbBi0uX6e/01kUMsR4cQnWu06cbsSs2RqC12Ql0H6qHd73vKa8h1lj
OcqZ3o18mzLsoFZOX82wP0sLXk43olPuzl453pkVtqBVQE023J6DXl7Rj3xffC9s
`protect END_PROTECTED
