`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2fx+O+xNvgj5sXkaBMsiPnQ3lynv3L3zCocl8BSAO4WHRXwdo2c1ZpflTAiswIQI
5bZDgjxBH/La6Ed5kRaOlpBphJi3Ggy/WopPyqpNtXhvtfZh+VxqG5cFc2B/5IYa
ycIuVLblTVjBGoO64zXP00QW8r1HT4i5cbszsLfz6q0j2FeK1JHAPBk4gpRlpFUk
Foxy5FQ2b2J2zRbFc16L4HCLCHK5m8nrjJ86s+JpayT88GFhPxcuMrfTvz13S4t5
2D2XNH2YjAmwQm8R+D1lNx+/e6nFd0yyiQi85t1ALySgcFKwHiX5ocMCZQ5EZyEa
BezY5UsIy4KN1dcw27qAiMnyuFfvkSXwCKn6PgLLeLSTU1X2HP7ou5TvHGwqjAVc
dv5WHpCfC9WRB8zc1t2XxjV5YMHvScdGmH+trf04p+qGKJ1oi6czVFhxL2aRm3cN
RSByszF22PCtzyWMj0FOuPSC7oU3Il/a90HViPzczIEZQ8Zg6rU1ic2YBmeIib2D
UyG9C3dkdn62pJptG3x6hYgL9s5DDoacqClyB6WX4nFX8ELMyT8i8GZ6MjoFS5/t
MG1N5xDcH1MPLTs3bCNbm2VU/9LjQM6yt1Z/xm1Mf1TFK7HTXLGQm6pDIVijvbLT
EsI6OhurJ+DSZppzrun6KKVNrHBFZhg66KqoQYLl8E7I0GTlp9d4o0Z25YIlK56G
heuoDM9pnrRx9YhLBi4g3D43ZL2eF1yWmQL1eeLF9tWuv0/c6F15KWhtKdhcAne5
N8C47SWBsfpNeu2BcM0jezVSBuM+400XVOw4Isg4G6HxAQLFlQYdPy8Tfpl4KJsm
M7Gcqcv3/nFjzPFzPG3II5Avli0Cmlli+S81KYPTRzFugvGBR/9aMoXpEY3q1rAQ
rA50Zf7AG0uG20uROq9+uuTCBW7GS1vteFzr/wybLSxLxDdGYHZi7snUhkAmWEmT
dtDBNbEqC28UQtUtC+r1GZJEgpXBFUMV74HdoRyuquFaMrsZ6ovbaoK+Z1qpCQU6
rJ9fiRMe164YuKRgulJU6/mdt6Uadc8XQBULl7kv/sx83RaRhlGy/QLTbONXvsW+
TMTua1aO46JdFHiT57wiGN2kulGXyIONoyV5Gcl4aMxooUuFUDYAhV9XDFkCpOCc
oi5EZ5fwxxXgkKllfJiBPnJmrQn6ZIqPqR1oCF/p3Bc9iE5rYsCJaTDkCc0ucZa1
cdLQOPRfU325FbigEGZO4kUq1E2qhlJ/fswhMzM72JTDzX0TKy7i0wbY0lFVyYKN
IyyMbEeCtHxlVmH3fMKijUeUWOTGfY0Y21lVLxkN7aH3dnZJMi1XiIwpZY0dEyCs
SC7AEJ/zH1LY0tMoEEtlakVbJHuVan/zYNfDsl3ez6+0eDMgd2mttqkHZ/iC1biI
csQeFnMaSPUUAxUzeTUHyYKWhq5IVzsRNf5x1nOVdarH6OZmTEy26YfNafS5dWJC
oC028W0zXJUUCQS/1VA5hNu3rlMgGC91Mb5FqLSpYFFFtQMMJZWnuYPDiNGwOKYK
j/47JYbiDMYSRn9EY5krp/aNAqEkYVwFg35pVLHeZhXEsfG3KyJbZDRLFuLhg5r5
3RylDlaNH/EQ+WbAmsR2eUFIDaeLOJ0RISE4MGf/oGEN4rafyLDeTdrQOX49oqnh
XJjEbtYl+zOgvjpsEknR0IfoEcHTRZYBQUpPdiKVsK0/pS1Z5UidGi6CI++vkWTj
drUsXTpvYYsv/5aT/RUqCf2QrMWEjoGiAnyQrk2bGJeQ6ZzvNgHvWWa63si9uccb
YMCsHFiw6YNtZb33DzIsEq2R7uoHYvtgf1FYUl/Z8J5EhAk+M1VklVteIfWzTXnR
iimEAcjyOUx3eKDvLlMUjRunA1RY4OqFbg/P1V4/YJ48CyFsdZRdGtSp51TIZaxY
LgjpCHu1mHdSM7h8xY0vPzk47K3x9CLor2SwIWB5AD/AL4t/Qd43e3AglbKkqHG9
n4t/86ZRyn+L7HCPg0aVBiWNv9pvFs43vyU5+vWzPVUdrnuKk41Gg+keZW4XpsKS
OdQiAnsIeO43YYtuYbyiFKr6MRfOYZD5C3ld+5rwSnNHcG6cJO3BGz2ljxdMFOMK
V8NS+BuM8qk1wTWIJG6H78jJV2k/f9g60fvd5clOQh2G0lUlhzUTzl4Cl8Wb9abn
r5l1hbSXsQbdXQ+LxAeAvdIGrO92ITCUBaG+QzIleRjGe6q4m1OQ8yRZQhAVrlEk
jUWTBCJC3yonjliBcUkytXrhHDiG52PAVkr499DGgH/JpvBoLRlFFJaZvnzWBV6S
NGBAzjj/tvoQ9Ras2R93uK+B9FtCFl48Lmwisx0C0BpNbusG0c4Su2z3IJzHD1wq
Hf+r090bP4d1HZn1kMaohkw04wuHYQgzNBOYRWaFDlTJJ7HMtexa492KwcU7paLv
zV6YDrhqStjiCrNXtPuXGpnLCqjxbxCQabJAOdUZLuVaZhdZof5uStS8E8wMjIWz
vaoEv7lht93/yKSzp2KotIQ6tBGDQNzmAJMhHCHFHShU2mqKEfOCZNgGb9rDXFqS
plcca5eXSl1PZ7W6uWFEDvlBpKP8vqmPmdFwFPlJQPOgfOQTRdxZ2531y0ZvlRHa
dQ6ZQPTFUUPQs0UOdmiH03UDhVbBJ+CbmWqJaFaFqhUv9d5CHiXmZtYwahpAWSMy
kwcklG0lI6jxOuBnomLXmJpV1UVOeBGJiVgmLaXqIjwpep7RQb0rabF4uCH5u1e4
S53Q5Dr6P3H1ms/LMBFHM/X5xvoZvCvGjgP0wAZhUceXO4DynTmHMWOrNemuy2Lw
3dFjA6DdlwvI6R6YRZkfvCrqvXScHY7jE9cI1BRJPN1zyBFtR5Jao8JwOtP6KgHl
hfLQglvhZXNHM1nldoZV7DtDbg2O5B+gi3UTcAIiVsBW4lFnqdZ8YkR08M/y1GB9
WkLsrJqy/8ZTb9A4AF/RGW+YnaFpSajYC5UlIqM+W+vdGLQhaoVjL1jpqxqwppwp
74NOlIsXtWqYZvas4BvhXWJJvuyUPb+VpVEey22LEAQYAetBzgZD1Do36hexUU8w
a0aE8kXdHDprAJN7Po2jx/qIE4obcC4rba3ay70N0NSQRhQmUj4ywNGorqKgcMza
2N/yf9T0+jNEanHRIWLq83iHmZ0Quf26ZKONGPRHEg0zO/DWo0JiVotcSQw82Y1i
+zwtgdd+wFjCt8T/RlQjFiqZGvW/0w247gxW1meymdDZ1RyIMmVIK7anjbX5QM4W
Jqt5XfLUsHbD7PqdZK6EiukQLYL6aP3ZYGuR7vO8ejOtJ1+H/cYZvDHLUKQyaGi8
4/AK2I9rbGhNG/WkZddcG6mNnCttwFdr/FgMSHN6OgLZeBQl9gxCmwrKKwQN666g
5U655hTFZgcyRkGg1AFIz+/Jv5vBh8ciNzI+11qQlmQL4LHZCa5knvHsgVy3eFq+
KFB1Wwna3P8h1cLZHE07nKLHuULUnyf0gaMNAwJ4b7of6PKbrNY4e4Hm3Y/B21Yx
9qZmvRhobGoNyvEDV9Q7K4Oyug+Gi8THWN+3tohiEaw4eCogrTqErAOeUjgAXd36
91OQGrZyNCT4tAhFk4RePIfGSi+X5N2wrs+pZVMrCrU1Hi35uCCOgQV2v9cReOA1
3uGHKahaqZo/814cjOUP2483Xj6gU78iJGArfF1BMVxLckC28Elk/B7p96YG9jas
DJPaCp1n0nLtT/z9A2UkqnQLwu1txDLmtgvRUvpUOBNeOJHV50a2l0ZFfr8gUgYG
tEINhumRJx7y9gzVg0W3cxMo6O0DeYqws3vlemVmiZHWlkzevKywJukJDRkmsfx6
tNMV6byff2FtunO7dZYdchcBzWtTcbWkEM7hSAegJ/0AV/hPtr6SGAUonA7WCfI6
0GGsCPrkGUO4yfeiqtkVD/GZcLjogAxFQBh6/QwY/VU14LdURpYfkJtPX6prdhH+
xZbf3wGkWooCFb/9lm7P67ROzgYgSrHhxE0msrapTFqAxR6oxgnq6rMEA5EfAIWN
zHt2CKKv+gI/Fc5/i/Oi7aLlvG4LiCPw0/xW72CNhAbAcDavRG+fEGT3HBcz0YwX
WrmZZPpz19R7ulI+W9RU3kMuQ74xM8ebA0OCE/JrPNmzPLoEJ36thSDFynZCQ+5v
yB3P01DSP0kaiNWxSzLCAOsiSPzWQdFZBWfBR6mmuNOBNUL2BfnRcGn4ILupMLBy
UL2SOKFE7wjJHf79rjV+GsejwZURkTzut2bKSK/XF0vsuYui0uT21JKShMrU8If5
1pGNUNZUWb0tppjHqanuqm3ivC0fMWrYir8AIUMgPGrfO7brRuiZF0l+e3l29Ymz
gTleCDH5JtVOqrhhBerhwE8pLym24QC6tC9Y64HM2yYKwqqnMjEpheFCMjdBXR6c
khPODr6eCEV6lRe/2pOtyIsrskHfyAWGbamWH3j0br+CSclhnJ5QqXx3fP1AUpNo
PFNvFZrv1xT7eRD4aTlDU2qJah8zyO1GURlHoAuaFAaKPYZS8lXvzWdtyN4Lx1xl
X85/3SSjstWLGYFJ4yHl0E4JHgxfQPAUkTAXN28c21Y893hS2fiyThyDpCcrlhs8
oRLJuLsfuroyOSjnU3SSePpjtVc6EV4+z7TT8crBFf80lkhH5UwrDuLJRq1HfWU1
lZ0YAN1huziaRwCzL1qYPRpSQcLI9nDG6no9VkjxRy548ywvsiQZiwYtm0F62PTA
GK3S3nm7SHn2ZX445ai7NekoRh5lNeLB5G8LWFNmFNSLuNEr+Uw1tEtPeyUStBlM
Cuz/eMky4vNvWqExBff89aLJwDy8JU7rn7nBk4SXdGFPPZ3vXee3f9A2hJE7eNtD
EIv8h+As9jst1GCuwIP8WQLL/DNY8s/VHy/zQFHZIvrKG4bT6rJAOMw8xzTYV5qh
Y1W+VM7DZmMozweRQxlHtcrUnbw+stU1rqHEDPYU0O1p6OPoMR130hjdoB7/C8h5
Rtn4GiEzNtECUtjN6g8tECsFHXLOtocj1BTtbZ+ZE8Pe1/JLE3jek3YM9CMXkGob
8UEisbgfTCXECkN5MDnXl8yTwwAOUkJWS2C1UN2vop3lHOr0h43VfPG0olBpMgKr
SDHE9PA7ItDZve8FEiMy2xOUnNRGuLRbZmqicTHl8TeUYKWYCZZ9ZWb+Yaa6LnSO
1GVV/h4Dh6PBcPCs7VJ5kiJcPF4YvFCXAdiD4AbOrS5PA7CnySnZPrhhu72KskU9
sHAKutKisoCfrPuTNwQAf7mJFzT6wbn2dTzX1SML5nr4fEl4U/Hdmk459aRYiZAz
4S1egbRX3WapElZNu+Ekc6GmbmbYi+a7nuIzCVyj7DMAFFiydyFDh3ZxdF9M/HBK
GRRhKCp3Hlt151/zn1433X6sQGyMw0ugQNeBpfMvc+h1ne4xe1FTAc+qoAg1ZO6x
xpbcYCY+PAtRzEC/WDplrku58tr7GeobSo7CzuKKk8eA3t9jhS86mYgzHZks2YN+
V02etk8b48yor22Ug98u5P3ipynVY8FBcVn6WnHDgdh+m/ZjbVgpTo8dzUJenNtt
wTjhqMvdbW3ZGyK6p3ba3ixhsdEaAX8ndjcNrVQ3tEpjU/mdaTZ1JZVia+wAT6Db
PQXIGds/5IPuWyJ7lp/JbnjUJ8tLBPTYhdZw+854PV8vrc4jME04Cc4OwYA0iuji
pf/tQcaLpKHdZcxwz1Ze2OqCgbkiWk+VtYMOqlyWPws4b3Lqe32TQSz/fQrikDBu
4LjxVZ3MymN9nKe1APAheETv9F863ivnzRSZ16QFFyfwQIl5vxfD6s3Q+c649uk/
VWJ0IiIKvGjMqfxG6EjU9qlEg9IM7LVQgtJmlQmY63pbq4kQEVhjUAyXby8xFPdd
u02rYcYmq9qVDHu10U/WXS2CnfwFzZSMezpclYLOeSA095UMXc6KPAfD101jY0BB
J4n70WbqJRY/DOUxGwmJN64zipidQH0Vt+AXeijZC4MFm4zc+rW0nypkdy7KB/bD
9iieW4EJZFcfZHHZnaQss0yzlL2u+YwIWVMiiKPAfBTzrsw2hQ5DpvcXF53ks7Kw
CiyYs4eBBTwRcilWNaaS5wYSASpmkP3mYmWc5YNx2EMzUIDBgYAeWjPvlCuGNW8b
9Mx8GLxssto9tXlwhiFoUcnAvc2O12pEdXx4Y6muiBhD13d8DGa4RPFYfOitPIWs
5b020mTAdgnWljGv8K8eO2Y8NUuHaP+PcgS9rXg/C2UVc2kXXmaTKipHwWRQvH26
49/OnOskalzhWlo0q+niAeoArQkoy3ogy1GYYZmnxTvMAT1AblEZsjhw6+rYHosT
nUOUPrK501GT4/PaAwvl5kSR6i3OgMDNmIhhPZxeRmQZzj6g1FTIZvrF04QTIiJZ
zEhqiyKMmm9qLC/Rp6OSY3LfF5tyP9F+wVmO2CsyCwWuFRhDfxsexM2owe68JcHC
scntZAnQS7ADxkqexmscAhI8i/cejicVwwCzxoS7Pb4ehciADrn/gyr789ltjTop
4DQssN2iA9G0gmKwKMuredfotfoG28f08cYbV+shzZ8h+Vj6nOtvWC1LWE9pnXtd
/zmauFEhEoUTq7/uQjXL8YZ8U7pwy2Bos4A0cy/K97Y2g3/xcLB9a+Gh1xsV/Zy3
bwq8XoVMX723prvwC6u1LnavdCGBBi3AGGuhyRoS/hbvZb1utqaqN7ve/UBEWl9x
ZTJZWAYOC2EoIljbpvnTDrSPo+jUCmdNibSSHSpoX2eVLw63yEWg8C36kFXDFYk+
F0CCtmwliagB5t8UCViCnFP83REikaHrJ26Sgb3TRSpG6U2d1L4DUZoglbbWlDuE
tHslYzoqQX+4HmVmPWIPqYxDb0lYX+HP06Pjq1/lZ+/hyqNr8GdZ/tO6jgpDSMVX
SRU6mRmRrQJwwl6SvBAmaP/pWm46td7xSHS0Q7ozYuReULTVsxKfuGw1mH4iWPJq
TTEJ3FqklA586NP2AIr6MEIJUwACs+VUO9lQXjBLfbyGHzSIZFlLewKMiAL3vrBD
xr9RbqV2E4XOs94Ya8iZ0BHfmaJJ37Y4nlQZZI/bj0MJ77W+taBM7LrVblZHf8Ty
z7IISVXoJ4LCZzTCQPKUW2whB+otvuGAeGMLX6ohZ1DEkEnUdGWAKdQf/GH0S6CW
Fj3qU+oE5OldvWizQovvR5On9pjDY/9yhRvZZUuHrWtELtwJWK+hMRubjKi2yIS5
mNAPvrEKNxy2sE18W4QynpDi0x1fSPloiSVo8iR11Umf21PJvPPCaBAMVHfL34/j
EMAdHjskofDNZqrgtkGnDhH9LRXHtqVeWtCIQPLA2ZSiYYrBYUFLTo1OTlA0+7G3
5XsQH+TvdT3ee305jN+DtItcJoNUY7Zh48GgDu2FBQosEQrbCsaIluKWpicLvpz8
hJrTmKf+b9k9+PebOPAi/gPF73ZYJJW8kfsXn8jCwzsi82MpjACfBa+rW/o9LkC2
vMuI92yFfved8HBWdV+nel28SnTGgjtf4omoec3ANlUfpNuCdsdY7Ellf2/p8bDT
aQlT9Zqb1AIOdp/KcAbigENmdvNIzPASYc1iwrQDmdOUZGrrpqMQssG3JeZ6vt+/
dbt7XOyXvYJVkoJJT31ewxZP56jOTISX5dLXR8/ZCLR4IGapoHFJxtPSfvstYZYh
x0vIGMEFg5kANC0LlMTnAybANw+8yyYhOVi8jQNB7d/kGM8N6fZ/jRJhUeRlr2ki
4eXWYpCk9yojs3R1tLV/lgZRikfNX5pkdDtT9lAKcZAqgjAFmyqJ2K69sfsJGOFW
KzyqP4wtWhkr8h4QHHZMSk2UBo7Gu4GzKE5AMgoaFHsGnGtRuSmaMgk+ZbBJTnr9
Y1GG4Nhqr27H4NEnJnUbgpzCWlGf6rlrzNTqMlHhO6mTlG06ZOTkpw32dxtZNNIm
a0uolOIcoKY6+nfICXBFYjhXA86+lkVeXceXDpBHdYy7KBqoL6ppcJ3EjMEb8FEz
Lb7Wy2oSAGRCOmjjpxMfyohwfLCgt+mZulYEdZ58KqgZRFpSu6rz4XN7MgaOVmSS
D0UkhuxKcK9GnUyLdYZWAmb+RnqW8QVENXOEbAWK3uMAnvPgiFHhXKDqauZ62LZN
ER00vcKLOq7HoTWugct6bFo0rnGSQQDCZlmO1ORytKmnFkX2J1rBgEP5TatKeYmO
ArRuL+cm/IEp0B0omCbz7BhCz4ZO46uOQR87NHhbwd89fSGuzBSdBe19JBFuzpFj
zdzvs7M9shf+vYQ3dC7+Kbmmy3RgiExW9T9FwkKfXtudt9xLT5v+I9izqjb+JqNn
w5ekpe7z9b2nRb0iq3/4w/hNO+usvo95AwRdrx6CsHUdSgScj4uo0gSqGj9nzO13
j/RKgOOlndjEBddZ3+Glc618OYOGeHAnJ+eyBxsXQghkPQwQzBHUrh6ffbTmo7wq
eaSXfwDeX1sVuHa2NytaLkVUSWU2fFZ/PCs7h3FqJG8U7+i9wC4YCRcbOmr9gB44
yrhrDvquVD6ZKN7Qjp3HCS0IGGzRQ7WQlf9xqysNkgKfpha3YSBlX5iUZeXwZvfX
hWn9XoxCedxkXkOMfdasAsfuPvrYdPmKg/RkUVZG2WLYqaFzLol5ygDw+fwfq4F6
KEx5Tg/PVvPi7r3E9FfRfRUKZiO5PUka4t3LMZUVXaQ1rwjUEhF8wTxPONMZLxVm
7EzxAYob/s31EWN9/fYwS1ScqUZd1cPmE4gwDnjkeHmGyPdefbKacAUg5l2db7eS
qztFjwiVlbmLLXa1KP4qhF4dY6p4jGgvS+FDca5pKhEijPV5CZxS09qWJMYUwPA4
3HwQ7ZYmwPtdXUPcot1uaCTcU8mi8Xj/mPwcM5BvWpWYUqf4ht/8pfj5buwcSZYS
5v4IkFveJ3G8Fe/RUg36gWrFwBu2nTMaAEn2o6lYy4PTyyrKWJfVRbaex1ljsy74
HYotClXaMqVLdpgCRxqvrwrqBano8qEhdr/K1RyI5a/PjglEHCxpsXh+9VVLOnCw
Z1t260+/YC/do1t1nvrV+0jGxp1XL9KO8qUoK3am0slj0BGeKyk+hl1yEfePULnC
h76X00YizwtZ2uaMnnIz8qFxiwVXQjQb0Lv4eBHY7uFR4X+TQpmJKCVa9ukG3JRe
9o8JhKMFKrhIL2XDEwnVb45pl+wJ8O9w1sHW1nL3zaqGMZNdbVm5dWYnn2s+Z2iu
doErGbi3ZbQHcqkif8oxDd3kSL60c4xNXESXrJOWoHCWWuVX6/jZnsyi/vsc5pdY
UKbJxktRCAA0NSI7/b/0T0FBaZrOp5pPQ+5NJZWj70a8gbvwtxbH1laECmn1mpPa
TrxgR/ttjWwO+cBFrvVMshsrQgua6TAUSFwFCgyKZdGk7WdRPwZZ5yzL8pdYCUe0
YdDVeWY4JhUCTAJo6F8nBL31PTOJ2vFWUl61ndmN810Q+RBNsE3dRu0ZcvyBvy95
/NOHBmCi+xOn6TemEJlCfze3ynPiezMKsGp/DR4kowDpVQUbPmrQ1EuuETGLZ9u4
W0N9Vnw+Ff6zqFEFXWwx2ZUPyedkEOkaAedeEavoEFwOW+FllpG/SAyFoyjW5Lhd
JAnDTjDx8AHlFmlZeUyyi9UkgOlbkEQl8PlVRCu+AS+1lRHlTLDqISUW4I0liDlD
EXHoXgG+aPm9Eq4RzkudzHC3NrFfwNzSO5rVcJh+9NOouzLDbFiCWyU06zSaTWp+
emI16UZZU8A1DqzSg7bgXWNRrtvVGNy6boql2lrKQUdY9vePTvTNoHMFyVcv/1Am
8Ij4aHOwnCvnsjQkeXNpjw0Ffz3OGfVwHanGQXL32cYuZ78rbS1C7+frSxSe4E/K
pCa2HC2M9XTc7u2enW+C8FRa+T6dXslHZUtEjFJodxz3ZjnDBQ5JSnpkRoZxf8Ct
iKrKy+h4CPLojDbZS/SAvrHdUKMCkRwpE5FqsOvYLLI3L+lLnrs2R0FR6ON0rovF
/ojlbAIp9tfXBumubXc1qyms3CCRtB8LuiGRgAA9E6b8tsAoYDCwBILsyzFb1k2H
hgqwmZ61RAFYFB1T3/iqyqRmfEd64/H5/m8I6rwgIgGjp6ptI76Zqc2ofT1Fd0vn
9u8YSaNOt8HtHFbyByOK39fiF+audoXFZIUfm3w8w1mNcz7C+EZn0rsoRvJH/gia
QUFfoM71z1J31kwPEx+UzwEPZLaJFEt4LGbwguQq5Q1+4ZivMIAFvrTe1yDVW8HW
I2+HHHHhU+R9X1fVtCQm3kd1nn33VIfB6dtU/SBeGwUuTWaSNy8wZc2Bcj/XJdWM
oG9ClfwXmZMwW9Y1nxUnA1fM5i1BHhiut/xnI1QG+leHUSY7ZEAi+dM9/WrVc0dz
C231+jKXy8mmYR2GIggpYhp1H0ul6tVwh3OZLKfVoVVQUuh2owmOZ3SGEzPvz7LV
D8oW2SPd78M6GcSuHtMk9ncw6Bbp6wctMYJtwG+JZ2U0lPlFAH8TCChvO4keDTFE
bg/WDoeB7lgLFA4CzQT1SKWlk7RsYIVDqNakkALJx80lI29EKjfEisv0qahx1/eM
5wQa8aXV1mT9f3q1r5pZ8DkFzDb2bjZ2mtgiwCTuhVOguMsg/qoRc2vxpmWaQmbw
siPAPtlzY9bjMAm8C46TWNMk5zA94tcq27ZDBOXrKfHY76bCF1WV/XcT1z4+D/KE
SkF90IOYaaEeJteOnC29f/M3sa19QjsqQL1whZ/kMixddxRa4dFVjHiugQPIApnE
GOe6Z8MWgX1HIZ4N1TwOIqz6YGYPV4+jVVO43lBN1GWPVkNSj4hXb2VjHgP994an
iIIGO3I1LaiJgKfZM1W7x3PAAwPw+3PJdlxrvtpFkj6YftmDo/ubN8BJ6+zekgMr
bg1U55Objg61QHSFfOZ6wD7V2lKQS217kHQ7/sYizyU2B06Xx3H4BDdesaGnQsWx
5ovJaKVuQyX6ohAQIiAgP6aPE3OJCWOBPZUICy7G3z5agbQFuILMlHtXtKiBQCOz
Qm/OgsAeM1tSBzq9rLRDxOS78SRddBa4wT1Yjeqgv5CWyuo1H/qulq1t1cgJ5iW8
1Pw+NY6T+pR7BQiF8nmwTp+Wz00cmvZio3kayVY7wgm0qfiDXqJWV/vy3HWcbZ+O
KGf+jMbsgWZeEoea64uVJ26Bff+mDSGCeP3/2s7cfNocZytWhQr9EeYoO7B8gPdn
8U64kOzgmwUtCvIZujWfCadY35WPgllD4mS+9FPf3MqzEmVX7vecUAmShLOV40Az
VtfCtgwXh11sFEmHACea9Hh/trUfHFlza3ScP7QwwAR6GvsBSAX+ZtRQoyuiJRYs
BRoWqWHFUv0xZIeK7CNXtA2pkyBDay4RRCtAswyF2xWt3N29DTkakFn+F/4LlvTf
IuS3iF9HsosFN557LS2UtpGnBWpWoBOO8wXvQPomX9clNKp+n0PW35CnNTmTkxDr
RNMLsKF0uLBr1kZZ1W3QOQHZd+v0HPWI1pWFu6EFe1ddYR7lh/v2WMv0MTB78s4j
fLdcJvKymEKTWbowYejHnNKbPOTjUB2ctsnsKSVukyFRi+FxM1gDRjEDZqzXkUGY
ZznfWx/b3X1Pl5uc9gF3iwaSLu1fQxgTL7oYDy61VucpzzAuQ0K82Mqoy8EFz+R7
8vQgYPOjZlaKCaE2BINFrRqPdnfL06jCgXcreRxVX0RNn9QgnrOg5eJi5yX7AI+u
2RBwUoWAzPggPQ3Htbko7SP9BWKg4IzKXQxpnOksN6F9EJ4ypqhoaQZ8UjFLjFyw
afd2H8Z2WD/DFBcC4VFhSoWSmsIqJ+ZbEuH6sVa/O1WqAQJAFKGKHiHR8GSH3X9Y
8S9Jh9ohBl4qJBY2UgCE/KPiEJe+WG7tbqG+go74PYfHDeuvspbK2KkK4lnlQ7mL
LsnB+nFCRj9osvYCCmjAG0a6Qs3R2wh46x28Ug5Gzqzp61g0YAIif97ZrGM84V04
65tGIflKw7UwqEckrdCfMSTJgJ+xOh7hj/m7NG7OABs4s5Ls2AQoPSrEwYPYqVFE
DMTEYxKy+PouBBN0PSpG97kgvszK2Ij0qegBwQirmzpZPOXjkxsdqU4FmOnYQLVf
v0wVBDOH8Evy6FwLQk9JZd073yM4ngD/EK9q+hHhXPkzE4rkezR3ep4QfRJbQZMa
hvZ0OzDvE0fXHFnpQ2GirUQ+CWRPHRqUQLcW/G/S7a9SkludbGboz80qbz9+dsSw
tKrq+RXJdtWcJa07TlCkSTXJqc5EzYjw52QiWfplzV/i6oEJ5QDAyoCcW4urOVZF
BgKzVYUbwZCR0aAWu9V7ZbTACypsnTQOd3vF42IKAsAEUZoln7ZD70lPqIi5aGSN
yBxYsTSFkp7Lfn8aWJ1NImd0RCgtpV4Oxr6b9tGZdt2VMWUzIN8CEB6Ys780lkEE
paT8TP3WIhjML1bo5s73s17DIAoun6lDTOAp6j/QXNayS7DL6p3sMpIWsbHkKX+8
Yk45iJpRdaccx4HtAv8f/HwIqtmqcytgEdmKF803ZVL9XAb/oxbprhHjWHvrmBWL
dRHBNO6bZ8t/9nHzflYLfz7OBJLE5a3AwweaiFRai/IKGG2SbTkHbCFCIHR9839O
MEKANuMXdXZDOYCEAsjAcvdipaa2zEH6UCZ6xu2UAhr/Tkt9Xl84X5V11ZzzbIDG
Dy12qgoN4X5FLtnKTG32BW/qieFffxKVG5Dz7kaOZvEcQAoy7x8ebrnDdaeIMOGG
gFrwkt4e3kwizA6qM4QR4XUIF6m3s43ydYMPxmkJEphNdYHgqdQF/BHs5/6bAyTG
Gf1fyV0yPl947b41GKUN0+2zjUCEd/WJbW9v2N/pDH3JKdbBWFQh4zJBoRUJRlQN
WaEnDDTWRxlKf1++UGztnxDAF5cp1JMlJsyCpqay2uyCSVfIt0e+guWXwcuBghCL
BBdLXu2sgPaflS0TPwJJl99U56+UpH5AXsIQXNStQ3kc/mViC7uNVOUpPL6XSm23
eV7GurRXCwJEanZqcsm5R5p/ATw4ezKGtbwsndDj4uUoDT3XOTLc1G1TfdONeIGP
xOMlMzRQOuEP5TQ7cSR0i1tLpE8CCPu9TfoA+dFD08jqFj5ZRxUAczFRpM3NnuYl
YKirqnw1WE1MMYlBHlvQNqq/PB6HDGxZrUb98xa2EhmuUKtlyeEYeSMqj4dNK4/d
sQCX2MumkxFJu4zRe3KJVb0uhX8AmooR4aqLTo6s4ELgigYR0r3Z8NnEfaJvgoS2
pHWen9V2q+hzOq7VePN+pJrz5HT/LXBC3nmdO93ZAamXw/qVCOJOpLri7u7bsLbM
erU9k61x/F7soHlu8hRnbhOjg9VOvKGCNU0gbXAtO10AjR12rvr6MRnX7lrcs2yD
jOS0IVCoeXhx3J9OmQqncUi0rL7gtBzXf38E07fxSly94Uv/cU/+dRQQ8uJgs7Wz
XAOxGFyMwwXfz6JJ+sagHnjI63XQn19QyALVR0h47IZtUtVqXT41jKracV5xVXRY
cTTEpyNCAwcyf5c/DosauX5STkfND162/G1BBvuRiagjGTENrX9u72xumbU8rWMs
hPPD2CUnILO4yJfDFp44zxIb84Euz4ypfAyIosHlFcafDfWWzFvLH7EhnEgAA02G
hBo9C6/e5D3z7Qg3JRPlTVmJ4t0/GQiLf0SCJikURz3LqK18nGp0wb6ZswT+gJVh
Ba502rTlA+ML+6egmNvxQjF8v8WRQNiVDtBe+KPYGQvSR2xNCFBLZb9apf+TG6dx
n7jueEKMIT7Aw6MjiOOpVevd4b6t1+fufdLWxWMlJsceAV2kwywAU5e8gg4Q2zeK
9Xeee7xri2MwiQF+0Fsxyztic9T6n+3L9lXZ1uymvqMpCpMTT949n3GOuIlX59fA
lfrLa7BD/zuHY3Ty8pB8VZzEexqyqKJZ1lSWNLdEKEn3lUYNTJMvbWbEV1vvyv5u
Byysnd1obHDW+x0LnzsjgsxBohHuN4EEzKi2eEWHfDaDBabVBMQfksA+xW3+3dRF
sGmEHZq/OWjotwQ4wCfmIKrnOpu7uggCtVMAxb9xHlQQg1zOMQ2Ltmq2ZFb4L96J
cxiIswYgogmnSXVEumSoOcqQz7yEVWUiCLYw986slqe1eUhTITy80qHtp3FgxkoC
muT8U1LLAVQUXPeZ9xBhb9iubrK+Ilk+nz4A7wmDGbeEC3GgY7E8TyPSsZtABPh1
aYelRjJ+U77qGwjm2MKhsP8jUESNTXWMtrwYgmqBM+N3xr6LvYa09JeyU0scnujh
qRe+JPRWwsUVTfgMZ9oIns68y1JGEuaLZ8B4PNWaTWuUsW4OCdenhBlBuQM+BwuA
jgv0lOsJ/icWrcbf7is5k8lncvx/AYaI1ulwAxkJMS3qTPg89imLjLoD0VOdsjUE
raPueTufDPrHPhJLkaSkuUzXw9QlqA5r89CZHXkfByYOIGSC8YAiZHA08gXZlo/m
shFoScl3IIXGd+EgoCgEP441Qf/JIP/nLeJjbQmH9uGXHpCeR10bkHoMfWsBWwq5
mp6WfEBeyFRAu0KO/0FiPLDjQjCUj7tSf0BQ2OPWiY5fKaH7uBukjS2zcDUofaOA
etaPpkTk/P6zmcJfhYU496Z4WpQ/+mG2weIW26vxtcFEzrNPdCiu+N1E0IupzKuw
/uZ2sAzNiozQJXfQ68xTyXGLZ6RBUdvHUlkg74FXbrjDY0KcGNQkO6nSzad6EqCl
PJRnq2czxfZwn6p5sZKSZ1dyOB94lG44VUZkW7YXFkI2pKFqjGKuITQl5cI7o8zl
yWnHndnVZFIeuf6EmsBuorVN+3fUJq0ZEbagLyFwirt0Y+S1/TMaMTsNrtWv8Uqi
cUvyf23opN5dU9a3Lc+P9tuBASpOdVhHcIOeGbgbeWvHI3FTCI4AtJMmbqhRIhdb
3+mo3rvThC8caL4unzFqbxo4+KHaBYL3BGJ/u+ypStcKzU2yBpg8HTunKpNQNdfa
zLsjylJu0m96vszpQWGaK1LHJm8wzxx3HosE2Kz/kYP9DDGv6mV5oscTZp6+SaoL
+VQo3Vrum4ilZ30aQGThSqvhX1CZtA3A2ph91p33UU97jcqzWF9jwjwjaSXMHhYB
/Edvtd7Ap/+TOojii+jHn06OMprzMtryitEO9evlpI1z3lHLSXxbkEeYn4I1Z3Hl
j1XITOuliN1LAxyBKqD5meE2CGfjDZ2zclObp2hQcXNdmS8E/pbNtsfUoaFhL6K5
umooBwjqrJlysxvs065jIklCrVCMw5XaG4MvbujxQ0eukhp+UGFgsv0TXP9Zl5x5
Kc+H1osFaLl6Ka3Bp/Ao4VpsJMelmZlHUJkoW5FoL9e1ZqNeorsEA4xLQ+8CGcFZ
oLw0DvvgTSMkUf5Ns/17uXp0XPXfLWfBfTO+Htqbe6HEC4s6plAEXA0bL/n8HRBH
+ywJTToXQNCdSU4v5P4BsQiNGdr9gKIJus2LyG4860OeLfOGqyQJY8SQsnu+BYq6
KcNuwjasFqepFyhEiIDueJAMZ7j948UXfoa4v/UUUNg+MdctxOrp8kpYpPe27m/n
xJmPNoKM7HSxsJCxMQGAadRWfFPrN98EwNZZXW12FzSrNa8K5fvvufhqMlBRz4Tx
+DBTpXn9ksx55LKhUq3NV9vQL6wShk/wxFBk6Wt2AQ8iNoGHVVC8bXgWc30kGDAZ
XTEzwqi3iK2QYWdX4WK3+6OL4sJ+UFS9vWQY2XdrZwzpHXXm8duD4ka127STat4i
A5vEL7h5LRwKaxTWOAQj+ZYstN1Ix8wD0iQ2EuwV6vbNwHfl6k4MLdPQwodrwcJK
qKnkvhpWYSZkaya9tv3gJKOC6mALLdlsntAwFRt+Qvv1+8/ujCyhc323Ni1FSmXc
vd/SGHCnijWBitmQ0BdP4mjhxgsIWCtPcUR1juaxhDMVimKIK+FXVSA+/vFbmMKT
81/aLyvOUdgGrjqx1fWc3zIQESsUE/5fneg//6ySjtGWiiM4B+gk8YuXbdMiznbM
DDAHKXAFXwElj4iKKxtb6OJ4cqvVa15BZIi5KIaXVb//3QBZNvSUcJqAeAyYF9Qm
KmYWnvsbk4daTOJ1V85MdwNya4ztpuLSTlge/0zRSIniVRBz5o/n4W9Fxa8DbFKh
dVrpLYCRpmBWe1T1lDc9yJdawEXKmnmUEMO4qoCSOR+ArZH7PSYh1cbpD/uYYdEs
xLb9qXbkovvIASdfCPEal6PM5I55OBUQXia9DEAwAVgtGX++xj+HOtrx7CeBNzPF
GMr6pN7sh5UoqBRashK/tfGGFUtLKq0JBl3dr1iXlTT+rrPr8TeqzcvtAUihGJpu
i9AhieG/wlHZm+iBha5wNI0y59N1YFx4iWm8dC2Z8q/EXkGghTx7c71avue7b4aB
PXfoJZQ0TfIv/hWBMWcZRF1S5bGF2iWTvUN5+MNAy0oi0DjmvUe6B4BeaJthCDaE
TtvjayzNtxji8OsZO+EDTPGVCRszyZ8ItCq2ihDOI+nryaVkDFjL+N0vbYcHNJRq
LiYJcWHX0H+S8hpI7Ih/LoEB00RxD6J8dvliUrSV7zaUice1UdJS3P4PgGxGUY1l
O/8kn+IvaNiyOAYPlGLPhwfJDK38YwEmt5H00mgqnacBq+8sOJwvEGIAhUDfdL8H
Rgx4hDWa1vuAaEUmig03G7xvNkyamGtwYygelWi6u1dHCX7+Sb5WJ/oBJeech/r8
WxVQFv+yaQ6TAo2HoMXJ1Ql0GFyIhLeDbBRv+lV5folWI79gPRYLMi0oA6DZyZVP
Cg0SCBPmcqJ4KIk3olv4y7cpndamvzJVyFIxXf2GLFOgrkeLI6Bj3dKTajW2wzrt
uO8f8QSksLlzcFQFc4wS06Bz1aKm410hhfuDdKgoSo30tb3bm6qhrt1rHWgZbQAe
/DR2MilWRC2GYTjHCBULR4ZQzVVYpcbhSoE2zvrqRDZQNjVG/BUvpyvVhQ75d/I5
dmQm3n7byNXVzQJdhYVw5oXC9hRae9eoOhSqWhCvklQ9fjcrPOttDH4Lf/cgc90E
WZYbNbY8DyLnYN/3JoeX4sKjZ2QZNxi+Xm9vtd/ifkttqH+8BI1knAqksCw8BKqd
Wg7lEWatqJ+jQw8MVEvwU7RAfZfYfRWGLS9/apzZznV0d5gfmCdeOB8Wup9+lUEO
igLYt2v/repYnGr8f9xM0BMchjE23GC29g0zZ9Ckoie6oSUCffkQ7bIc1RWbHy+s
mV1NWy8YtWq+vBreZBrVK3PfzfX8a+PZUbraD0eLq30lCCAxFN9S7gQM0mIf6kJe
C/8TmPL6zh+smeZRx/xtCOvZTll3bQ2pqEm8Tte/KcbMP59lBUcxVCiE3eQV53Vz
2z5b7Z8BEI5qtrbvaMf5uV7Wkf+LiRD0utHtk9GbI8bpsUHR79t7wHzolybrM/rD
nw6/AzohFsY5uQEhs+PthThs70o1D9NSs+b2WPpo4xgWkMsnujYKQPiG3BRveNpy
Bv+gZErQAkbwSNJNB3uheHLekutoekf75kE/GPM19qnVmuOwcUpSzTUkfmbRPgqE
+OCjiuAfuLbSOC1OO5F84FI297nvfdKtDdBmz1uQKZsXkTgWnKMO/iWL5tERwv7a
gQjPHg7bSaGPoRwZ3NJnKPm5LWXmRNE4F1JO59qrvpThKmD12b2pIuA/IkDbmZxI
sctgrdpPW/uX/7P8jwZothZ1kEcldcJgPsVQItvlZeuj+HDPc9T6f91Msc9KJiWs
PPdkCH+womlUdNl+taVkqJdwU68KdqrR7cFNNGYIncvPCMZb/jvfXSUIjsftS3dj
Rt4toSr9gQI8bgGkP1EUe54PZUqesjJU2jZOwr3jw3wwuXG5+kt0E2V7Wy5sJoU1
wohqgQVTwbyoXWeKTyKuY1tgrYbZDjH/jwfleCIVw3agkwxdlRAyFg4jaPp45kyF
+6VCzaSxpZvFpDfJa4rIl8ksOjxfzMFVC2Jk1KtRg1SkTVAIm7Wrah83iykSUu0k
WDhGUOeqXMX3iFBx5CKgkOOvanhs3E6jWIgnaWX1jwAwbjfZGd1QvItxmR9Ac8t+
5Hd5ZLNCu2+MKNQRMBwuku6DtflBnPVjggSGrV+UC2si/GvwGdF8iiUjf/oL5eLd
FYHvVriIzK0Jl52/B6Mtu2vpJFPJV3E4guDVIQmmSMc0GMNBM+5D3E1hm/1UiHii
iOo6K4Gv54xnKiIhbhajf0ruf8pYeQaUzqlYQrHYPgmnUMKjPh8MNOFZGYM1R7MP
DtuH3FzXQOQlFIGfG9n+d/osg82zbPgIrMWnBqEjnjfUOMB6aircDYewvXPADC0T
GTYj6e9oxpbxhWQ9FHzpgZY+C62OkwqKkd6bpxrdXc5GJNfONe8cqXqFlu9U7JSk
k9OVPMJUguWUch3bM76572OOZpxQ3Vf8rDR5EDQ4QLq+sQfVA3XGaU0KsnEv0CY/
yCh6D5m4IfGoD8AAG0/h0NynkKkWrOH41EZRMaBReEf2mPoH2b20/SHZ/9Ts0mKb
Z1Ehv83Kdn0ssJssS97GX8APANPB0AZ2QBLtT8BD1MR7hjtOeDeygsuy9vlh67PQ
ziEHW2UliPP/rapjyonyhAzBcnGloLKKfUfdNJuvDUpWUY6C3OUF05Q0NY10gs4M
eg9oHxJuIz44Zx9rVthZDk7UbIOrt8VeGQ6yzdn8AtM1DPo8pLpmMT1R2/VVRRjK
FFq6Wq5y23qB7vZHmRSoxiWGvXfwrxBjlyokpWtcbwal88If3xuDntwsdB82PQ2U
Ks83iuXtiQsOH96vEX9VZ7GnuSSG+iTba3CuuZTxkThD4T1x/zb7U7Oc9x1vzXU1
jfxW+zRslWwpqvvxEfkn8TJTOTS0zCA1YbI+K8uvI/jWC8TzqPcIhx6uchRZOpCQ
ncAWSCPxOSEv1bkyUqgXzGNj6spvjhAwbW5Xp7Nlb5KUcFV2NWIMF92H9ZZuDSDs
/Jqgd+d3Uht4NQKl2hm5JgjO2k2d1IeRHgSS9tFw5gFDbvdo3mfm/dtcQoCVWbfc
mBJ7joX9QhsMfRESasgd55AOX5kuKWUmCH9kMKXmiwGJLDlaHvEEU1tS+14ClEna
m1LAfbVa7BQo7FDr6KYpW/zsOOIunidpbwFlyh8VgiW9Mz4IVwT4/k14WeheYjKs
34HIqA2uLo675gXENYEosMI/KOOfTntvfpx7Zqy9Yk1Jy0zQxjHZL1AyPuVfPWb6
IjGOOD2HXQhC7h/6tXbX349Lbqe9u+hRf/8og3eua1CnXgZjGiffqW/3ya7qwesY
4YUKLUPY4uQxe+UNr/+ejn+1t1YuiCfmbbkb6dDu7MyOspJonuDyc9mNpNwpZ4D/
vfzHDtvb/dRyw5/3TY2ARNOFgARyg2iqGIwhF0YL4uDGWx2+V1CDdbgxPop8qiwc
guyDHsmsVrcgqNy8XNb7jcCgOFNZLB1fZxM1sjHnoZU4bfFAon3GA460hItTlL9I
cQrDbOmPSwoRg8lRo2EQj7QSHjYHVPDmxo4Kg/FVIRW8I1x9/TJ/im9yx80sDK4n
ZgqjYPrMeCmwcLjDfG+IBceImyFAX5oQrSfdMCxu41WyWLuPQAV4ocLipOnkU191
evthf4QcasQ8M4euiCPbnRb/ERRWeqK0TfNfMbz/kU5ECLSxFC7SIKGhW0hwY08o
LOXfVQYkXNjHpyn+BpgvhZZ32c0H8LFvD9WclwEHI03Fw1gR7Y3dNYw2YNIZ/zoZ
iaJyPCWwPt3sgFA9NXi6YbjAEVaopa/tsyFHIdvgx5VTMTtOtr/v4lQbL9OYjTg0
VcFPiJjKnnnMYS7tQ08WafWbmJFQBhI+Eqyk6W401THjzY/uk31oiXJ4Fnjlxkqo
XRKmAqVJ+zXnKYjCvY+AeZ2PWOqMo3EEAYOdemyx6QxWseeY+Fv8x5ptJUpr+9T7
erY6bcq6TDSoB5rJ9LCyClr2nsaDLmPyRV3aMVVDXizF2hSfpcB7zYpD/L1Wk99Y
m+xag3ejrGVrVM0Mj36nAzdQr6eve4fpRrP5a5djo96BzytnFONp0atV9MRj7OYL
b1w3tfUZUGRnlx9Hju5cOqi38Yh9KXC3p7CIyZY5CS/fu+M1jlE5X9TU86RGiPWZ
kXqY0jWTxh1q/1yQySuWZZg75f1H23oPeescTJg0vhcMEAJZ2BPoWVlUh9DeGE9B
HwBggH2Q/qUaqwNS19qSonATtdyMRR1KvkV2g/yFRIYweklQo8h42+uLtoPLgrHL
kExmSuwauDA/XtluoFp+7Fe0n31AyOh11G+Z5/w1m1EltOhr7tClHieV1KxMSLHz
miae/pExBSyPLigI4dtZB4xkvFGSkLGMIrJIxXqMVlV7+RcLwu3X6nscXuVDp80t
BdtOfcfS2iEejMlhrSnCVhmXV+5OsTi5p2BiSrB3lBp5kOl5eo8qMVH/yuXeL2pU
dLQlyEteg+uc91VAxYxrj48CKMHFEkQIhUpL+Z1VgeT3ycb7P4AqC6Sh4GxCyRea
dvIQzlWeXoGAR/nNelqqysnpYFSWu3d1Hg+YFkGxvzkIlw1I+URgiCR9xIPwytP+
bdFrQWxqyS+K4ipwmcoJ5zHcTbyWz/+NI1EonOaq7xuaIYOweTBXE5trZnZPPXg+
oEKTX5A9Ccb/ZeG0IWW43RRr/WFuMZFNWk34XcCIlPLiFUYpofyfPzJ+Z9XSSikh
7S7Tj+n0dnVa/Q6eSDF7k7qmimNQwhPYYOrthCYas29mnKjpRqQnWEPWlvs8BCkS
EDxB8VPijAxTNCnkTZpbsbfcp7V50n0yEYnABjRPMsWt8b54HDFvP/oCi9bipbai
lt/McXsEWNKiAl61jJ80oehntlrrGm3OzIsjq8zcxVXMfuanvkoTaiu35C2AAijY
VmDDPHYVfJT9pgwZZN2ruDecCnxkwJkzL8Evn3XZf3NFEzXeJI/phBurfnVA3U4G
8ct4NrkzArrIO5trtphXX3sq3ekLHE+dnjrfLSSGK/3yUaTjI7A5nLEmF1WyJsgT
/nGOblGzCkyFNZLKjo719e1UKTvuG5sSWTNS4OuE7Qy69NqW5p2YXsIwXjTTwX4U
r4dsnjv4qrET54fS4pAIZR0s2+6Hau340/Ajxq/NwnHGI0vrMnY7s9rhnev4LS93
0nEMwha6kmD9qpsY2KzjFKrZQCyL6hNuLyHhbQcQrwcJJPtePEVJ4efvLAQbBast
oPAxVTomUyidblUn2ZXhO8LRNHP6vLm2KCczGkTFYfhWwCJM7pLeOQ2Tjb1cxcss
IKpCcpRRhBVUrIVI8NweaPhb4oF7Qohtf/HryInh4FJsLufMi0xq8LOxSCGgfHfO
1gfbQGmV7yO195Ww/a3GvMCSHy33fWzmdYn0AbIN7kC0uNyEY9bG4p7FZa3g+fTf
J8tJEkYkqq5t7RQ/PrUATGY/NQ4XOmSsCmkD56VQ/wQZ6+kDYQEd21ZbY2mkG60T
AVP2cJUAXpgccBtNRm4IeBZLD66ehyfUdFCnx3+m9354AZT02HRkIgeka1sEXxoD
NVkuo5oRyEwm9CF8hedsBJdcFXBBXGYgRvgv6epxdhv4Y78W61VlHWaIFJ7XlijI
wIQmig6vDyj3R8V37i+3luSpQaNzdnWVZEI64Mbqt/QnPV24ArDPtZ703bE7ictk
hnuid/ZEZEAT1Amfes7B9E0VMNP5dIIM9K5HECYU0sQ9lc7iEUcrK9ZsBthnjFtM
8SmyK5AMMLLvimUEJppGGBNHUW2dqSSHSjSHvlBihVTegLekZULF/ngQ2Body15k
G8I1Hjvtu9xstbwcVz/5sSKV10lMCV2ZfxXNCeyL4p4DGrRwNVrdlmTVMhzSyg7y
q1VjqPEpWiuAzeVSiK/whMLji0ut9YF8UhVqH0HqXFIkfZ5H1hbXBP4QvFDzY3n+
iCzyQCk2J8rIMjGtDPty1Uv3eNtr0L8GKN10zrP5+ISak9PWM2hxHXRK8qn5CR8n
/CAOJjm3xpPDBvjYEkK2d3dFH3Z3IYcR2IFHbHdrL6jhUW+I+7lgBHWNClKXBe/i
9GDGmM2McTTQ5SEMcerneJD9HI6f91Sa7qCSnRMscEirzVno8a+8KPffipCtuxoE
Cvj9tSDXGq+H2rPNwCRHr7MSPtWGUgG5+jThGMTrFSj+50L/5gKIPF0amQh1ebBW
jY34H+zVgPpDwoVGcMaYmTO990nVLxS1q1Q5WgAgR0nRTki5XIxcUrDv+w72Q1YG
3+UcGPP/x4zUHs0+QxaQZ5o/d6McKewxA7XUULZLasZ1MDZj5GOXuKPFqrE5E3ua
wClmSw1DQcxHqNd2VHxapb4JPETNoHgSI+v79a5rPwCxpt9ccGqCafwf0nD1AXUx
4Vf9YC3ceKyR4oHrEpSMPFd5kCHEuXdW1IyltSgzBv2e0byM1p8r1QEQawjPTvHM
16NMCcT6kC24gFPSMJzy61NAsZ+TL1r6b+MZa64Cb8l4UjFArR+bz0bbTgRDE52H
gxvmt5ocMllFPpNg4KGGCzpgcKLRiSS9Km9Cp8y+mtaj6f3X3AatOgbEJtXeovUE
POtdAfgvR6JYIk1xjvjpEafwJXPLM9Q/SCr1v263/BT3Bq989FDtfuQJdcEom15T
tQDluLS4423kxT/YcFm7sQNpGThx2zV6wv6hsB5Gwqz3C3vbSU1lrzbocWzOfgcW
C/f95nKgrWrm/dQGKohMe3ISN/2dFqc/Zth3lPYNK9zE3oftToR27Bo7M9kz2g3C
Hwhn6AMOTo5f9PxqgHxrlFRPYxRxz3i/2v+0mUjgSTb2P04/f2UvXFxY91BjHEmX
okvcKWfjhrSEvI/twZXHvh4H8dihF+QvAun1H8LjGSo+gaN+MZRIWXz7j03uJM0w
mP4q9UvUYoYatfxK2Bw/7g==
`protect END_PROTECTED
