`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0fwtGQdTNJRD202S2KBHNVvI8cs/PqHIMQ1ZTCVcAIlgZ0q7Md/9WAMlaoU/usl2
Vij9cnNnsuGNtnd0hWFtyD/XhmiQLvU4yL9un/nj03ntvn23OaERPq1D+HJaW+2V
lWDFMvVBNF8GnS0EQi7L9Dl8Ugy4mPqaD9nlJjrsVvnHLeyQ9x+PnLWx823RCqnR
X9J8gMJreJS53Y2e8apKBWlwnwQcQFj98bz36YafcoIdWxb7ErXKdRsi1stE9WUs
tpGAq0QHOdgP5M9Vq1GVGpSbjMAf7mIW03TqFeltXs/4yBnjIxTf4n/etxp3JMFQ
ksGTR4+D1lXrSYKX2vPvdo2+JiJpXAKIQrM8DLCQQeyDOUqlTqaahL316tqdk8fX
XVnKu6zphp6j5h4rq8aHP61AzYIXcBPjVWZZAHCoB2W1n0Ax+j4Gq8udjr52RXdA
WsTX/jdtBS4rBd5SJCMuQLAgChACPw5ZQ67sbv+4E1QDYDRRHCi74GIZLw9c2q53
vC8AArRzrudGs1WNxA+uEkAVcd4OWWBfmE1xtP2mVfE89RXS5SaUryW2Vurht9fa
LzBzXaWlqF8pbCVJtlDdHP6cQ5oSAkakTV7vvaTErXqASSZIyMMzoRWy21zySIgN
picBNeOKQOi+R+QIpvWCg+t8gNgEN6XP4NVB0eCQRoMYXeozvXwn4yvjJS/FOSjI
km37rlerEzcg8IwCqk5cOtBSr1OE1rboyeGI526cgL8w5yDNXIqwToSFvld+2Jbv
SxKOKB7KKlxukraQCFod+9K/2plnODiTn/5D0VM3X3/PnWefcF7HSJroRCrtn6ez
t5vmY6Vq1nTXQOS+9dwnacWntFSQxJeuvaWuwJ7wRbdLby/I2QdDXk2q7lDndEFs
39KAo+HgtRp3QVleYwFv9PiK1eTbSegbKrMbusfYoieWvDbU+QqCtc6Q5ALz7yA5
freHildhXROLeErHHrIOUXbvV4QYzH6CKBRvLBI0IQdehAuG1Qii5x+26WiRTC7a
RyFDH0v+UwEykj7+ffvl0gcxnjJ/uUUjEcMrQia/F2Hn7XKS62ixAxfpg2VTrEL4
SkEtbsb3ImCOC9dulbfWMm3DRMhdIavogry5kwOpNG0J5hLvP5QXbfPPjmdXHaYQ
FJxmGEaMz74IKAj2j5S5thqfjY1t0a4lmnnO0lDEyodqDlW74VpZrvY0wYOhGS8z
dZasxGRImYn9lymTx2dcJZhRyycmEaENyyInCGaA/4Pqrq1s3aWGHBEWrPZZU3og
0QKfChpC4L4S7/jLceWW2XkPRRZU4wNYkTMJqvF/r5AtiM3t4d99X+owTv+/nCi8
SY5yA+CziHTuhZWPRuvGcEAAumZvWehIIygSTGhqIz8RmlJwEs0BH94AawxLaxEH
X7zkvBqw+YHb55GG9J48eGymgNc4CgIKmIi0t+OfmLVQJOoafVhSA3asWTvjN1cC
StDFhlMpksmH20jcY4cih3Zyk7CmLVxbWfYHSpwP98GJZEafbDi3u6e/wYY7DZsW
bgG0MTPjiGuCDLIlty32ReB3cE/G3ZnMoBvNArQMm8EXoLDt3S8xRyezs8BJKLOf
xp5WKB2whGdxhVWfNRWe+IhCa05fyeMhe13UnOmGImCOUH1k0249oVnPpI5yj2J1
3s3YtucqbIe8CC5Y7c6EYEtw9uiH1vGkhwFTatGBppOHbTqip2EBD72xnRUIMEbP
ij4Slg2JkhtKXOPVwwGZttuHUUSfER/YDVh7iYBzNYjrYcua9flAHsXNBxyFRwbI
jVH5jTy9k80KXogbPbo5/Q1y2pYbh2x7B/axOm3b6L+qTd7lZGpfsmTMnzBkCEgu
p8dqWeg3/4MJ5v3EulwrJFU/5LGwHyLNmp4xRErAgT4BMaFZ3lhBaUIABwfKECve
0mL8uRftVM/INuJCTD48HAdNSuRx234aJisgnIJXATmB+MoewI2bxRcv2e/m59cB
9kHKuZPbo4NR+05gdpGFlIpCj1npPrIW2TaRBCIZRewXjId0SqSomLC9DmeoX9h1
96C1Mxk8J9KGIQDtJWjz+Eo8lchM5DysTEx6TIjvM36IFZC9cWCQgJZ+Q8d/mTIn
2jsY1l2OQLEyVr6lD6y7x+ZalDVaYPWopn49czbmKC+Q9+6LaHsMxLEBV+4d1Yru
bZCBvQ3qibl3AhFKzWuYwOpKQO78Kbe1Rsx5m8EUQH7iKlBRyVUhGznTy5V5ytDK
RnK94UGpQ3ff8sZ5DaKcuXSDHCzPdDs16eg5WBnmlCbHhaDOxnWcvs+CkLrRXLso
14s6tYcKbFirXOvsznyMaKlutJf2AozRK8YXM5olpWvshamI5rKijLGXbAQyglZ8
5rD8lpqp6GfLj0I5fX6qD6rEv960BHicE+UTwQBTvFa4BEy7OIuD0scdp0xzEeNF
mxV4dFenjQXRPcfONylX7SLNpe5eGXnhKa2suI/k1dBjezSad/ZzseB/P7mGzvPV
Q/eU6y+LsOloOL6Go4Pgq8Q0x/71565LKbhOjEkn++iNY22wUCRx5VvOaxpt11mL
jNZwmYh3Dv/HhbvnWybb0p9VThOZ6sBjqR11h9goY3WTu+q1MdRXMEEFzn475uCL
jtEgIh82dGS1GVCAZQQzIg==
`protect END_PROTECTED
