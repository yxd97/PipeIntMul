`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GuITbmMpSVjDG57AtEqp7fZ7He+5nMHVvA/mnZLHDjxuMQPr7Lb/WEDCTbfdtWsg
gT4pTHGDMakdWzEVoVufzQeLDhIPLrST2ZCVsyh8JIsUrmiZy1u6pmlJLQ/UetLT
YVbSsb308a7rmPmQKRKAjswjtyZRAJVSuQQ+RhnW/T3lzyrop1km4KpIvlYqoI1F
zn56ltPs/Kq9N+iKVMmPPzl0yCvv4SccUsqXp1nTQLD9ZiWfdDWrsPg3qryop7JI
cQt5CwqV4gKOkp3M74h5YGMMuL1amJr59f57AWs/hAjD5BzxUd3635al9XSvB81G
i0QMOHXzUaRGjLEh1CUilYbqp3IcPUZvmEB8ZPsi7GpTC1tJAfdjnze8h581RBgZ
gzh+NsV5bTYGxbVD1OTDc4UTBMLPwHmzZ4h2+VTNQ17fvVuhwVyfko5nP4w6DvE/
cMmYcGrbqk1RZrKWHLSrQefYDB7v605mwSpg/AFJ5R9eJ0mBLGCrtSxnzFyRj85G
`protect END_PROTECTED
