`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ivq+8mqWM6DG+QBpQLmayAef9f8qTfI0jSmjLBZ57sEQ+s+S1xiBchpM3YXqFGSL
lJoESBGryohr962+aizObEXOGe0HdA41bUCcgT07Zxq9OXRIImu6AqHyR0fVZxZG
B2k1dAmcbA7psFL5mWLA2PoXbqGWMRQU8AqW30GjsGm5jx1zYD2PLwYilPVhgofj
Wvvzdqdx2/iD+hk2UeX720Bl91BlUm3VnSPev/iKWdnftxZBuVJccxzJygrPZxmE
s/gMWzmi3sMZp91toYQrB2KAQ+iu/2kdiWvWJJ+fzNM=
`protect END_PROTECTED
