`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n0o/RwWc9jjohzdtkqj7BTAX7cCW75MgCew4Ill0hNVCdMA9ZWM1JwD+B11To7eU
dW5o5LG69gFnJ1L67TUr9Q0KUHozuDKmzJAfLIxpCunZfPSJT8AS+5pqLd8uAVpQ
3cnAOleK/mQdvwtKaCKj1b5QyHaVDkJCXCIaCqg8I4M7BpyqUFys42wSXtA3eYQ4
dV0ake2ekCrG/45WvTZIApncQf8d9Xbwvf/s5X5X0mOblO1yjLsXZcoS+Rzp+Ui+
J/xX8ruBTFOIyvZ6VoNR9A==
`protect END_PROTECTED
