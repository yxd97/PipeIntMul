`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3sfblm6ZXKbrerse0yCBBhG8etgnPpVj8aEK7eRwuY/1mc9f+nxRRyXx3LcM3R30
x+X3YXFAzhquBX9UGBxgn/z9Y5AKy2LoHDofwH+Bsb+kGT3LSGRfIUA1MY2geSLq
owWeSWF+m8e//Um2Cd8J/j/nH7x5aESrWz4Wx21vxeZEDuS5P7SHHwW40I1YuZTL
hONV8OgNiRzURyk9UVHStnWS8tBaOIJ+OJj1NLlUJOpkkXRZIM3cbNDLJgkid1q1
CG3qn7/H7twnmE2ALaT5YkiI/pUqL9DbzwF8kJBEo2EuZIUR6wSP+pgieLEjquGA
fxXWl0RtmAGc5JTYpZuDVqmV621+TIDY9dAPuHhbhJF9774Pd+3GE/HWqcg2f8iX
tyHy7u2AnYSkUnq8div3rSqkoLunrGv/1MTFUbefeY8gqcjX9OCqYXM/lxe92WAj
S8rw99x2h6Hi0rkoY82Qf+U0iKk1r9qCOP7GzbV+D/BLJ+++pqLwjzs1JnOSmPVk
L7TR3sIBpNls2X3q6liHaINOGqypZC0H1CK16D0h5WyHcBbGfbLFeqdneuFsebDO
iG7MC31jxcKB5dZxBus/k66JjMfp1S7kJd7vr/mMFIMrLzKoaZDV9kndb69sDPrh
X1oTskVxIvBDycG5lSFWPC/HHROggyRUnCDTcW2u95oo1/Km84SoHVfftBjY+Nad
2kxp6f8fgVG+zbFLfE4XfHQbgqTPSbdSQIzX/jRXBIQY9VZbUr86MKuoOdWLF2Dv
j0FJS/rKZv6fC+2jAxfVMkPDAIfZ9U6zWAEx53rypUJk15jcOcuwCn56CyGdFuCC
IIhLKsCeYIkLbwxfmhYvTXYAMoorCrbEId07TqjZBJ/lI7G2CFUu3i58VodxB9xt
XWZpt+MOFZ/4S7cqi99Uz9zbnYfhXFHu2efA8KqPOS0=
`protect END_PROTECTED
