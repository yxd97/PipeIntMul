`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpN2IGg06CZyN+J/Em0DW8P3NeqLJZ5A/5sJEfk0SgIDJk+9AAmMEvkcPozS0I6x
YMCRARWMSmPQUF6is7AHrCr0OVRS8P13EvRXAtwFVjgk4uzTT9yCkjCXaqMJFEXv
HNjKhA8DEquaMbkA7y1iwmbrNDnfZNCWReMCnp39+qtHKu2QAoErh2ti+qUrSYfG
kRn/cnHIA6j+KI/5VeZ6xgT7NKrCvUGzJrcZTbQoSdv5jWGfKOVcTvY15vFusvv/
h2eNuYAs4HpD8ne40XlLnYtF+cTnRPpNa1nnKD0/nNsRJ8+jyrgx3f7SDgjYtxdS
Mg0opImn5iaDxoYE7Z+s8wTYFAmg46JX4ew/eyWh1rVSIvGoHmkDHbhG0LC/x6vL
/JF+hhq+IFsr0vj0D5eNpw==
`protect END_PROTECTED
