`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oL6CqRr9Q52BivuIjpGzeluk26goRa17A0FFpjV9YU++FDHqDoN+OZFnu08ExstB
JwSkJoMSWMifbLCGrWXXWpAcixpU4IzRcxDyEysUzli+RiJkV9yyDrWZTVNRqWRe
M6Wf2R4qypCfKHDstdOKdBhi8qt7pO+ReM9abxvrG1OFXFAKDxBbgWHbi6TQZHTa
4pssiIcwd4FYFlEewT7TvLGdzPXs8gP6FHuY7NdBEMg6KG33L1qE8thslbgQrwFt
4X+TVNvj6QjG44rZLc557DlIUV/xqSszptpmS53arXnXODU+ad5TV6wlExGwQ14N
6UDsIZLxIJxrNqE/jDdiktperCi2/NfEiwOTPCwpn3lSMneBFloyseHZ04zqko21
cCtR/obDtSJOfxaNavJkv+iwDdt67e/fgGfYzzxG5ZsxZelb43FrsfihsKEF3HLW
Mg8ywR6NajKvMidmXWdJ1+21hl1jcjIF2QLP5fjsrSi10ok0K07CEOYGKKsBWc0+
j8/Qp7BBerr8SuEJ/aZf5UuZOPoH8lndnKRxnLn3AwCbFftf+0Sii4BgrbgkNyXF
WMNKD+GJpiiFjwvPKL+Mr+ir2b+8ARNAQgm3WHcHG/MXxsoAI2R93IVbyuqDvGnb
iYj10s87/3IBIhBuWOsYQP0H0NkLxs6XpixZxlaC/t+mlkWc/eL+ZQoL8ub2ePbP
sI3IffLA8msG+gsoaONkQUvTMeLTCtHfbXpN/Gc+J6BiYsMDNt4RqYggP1qmLgXZ
zFFln7nu6kU3833t7dpcNz3Zsy4dDX1GprE623kDGr7uoJKaXyBED+9c2DPux4M6
riKbCV/yRTGI7+0AJcUVfqHKJDwKAnRv/GYnNF28OIr6Ro629pLEyPzPX5Qmf670
FJLIkaTWXtB2/EUnC29uPB5AaQmoGpO5RyV5bwtPAWfQoLkf962kwroL3DxUchBG
onE24Jh9aT44xKIVYta/8AYQk99HLfYQEik03amWL/h0RsPuuv8QjFegCodbPA5+
VKoaw5i5/AJ9n23MaFX54Fd9GUpCBOqKwxdCF8izxoKAAZxZSJ2yRWaZIzykMgF5
arqvraZkSsSRE7ZDWHGYmA0zs1/hUGWApf9X5VBBPGWAo37RJkUj2F2WGD63MXDD
deLEWBhuiWUoX5vJ1r72HrNp86usrqbxBRc1A0kOkuZhsEPyaflgjWAQJdaogMKd
XPwY8R27DzR0MGw5yfiZLcmlsbQ7Jjs+VkVWXZIw9uJ2N1CKXgDGTkZvr9fN0kck
LYpHvkrCPOfFe4wTa3ITV2tvH+Eic/RzLT5mv0kGrhbIaKStXn0KcXkHvoOO+WuS
+tweC7eEGKtfdW/d2KzkBLdycG6J1keMgAnVDCmk5u0QwW6KrgzmHOsVuboD3TAQ
ncfwRHcEBsA0Twtq5XsGOehh5B+/2UNjf3/zfXm3vzNBNDu+G9ZKYCfo8vRu5691
y0SKDt2fchUHAb9eKKT/AqlT441ImXdKffA/jexlr08j6XkuW+MfwWb9uoWVeRDT
pVY8QU/Z4kGgzJVaREi8VjLZC8QQyNmUbSt0O/0K3up1v/asjnJtQOYuFYKvZHgK
Jw0ePP0yhlrqYVlk1taL5hGSMEZ+qlgZ4lDfnknZE+2ftWwr208BwyNwXObJJwbv
YaAevMPBIJK2IJj38PaowmFKk4uLI/w1swnyfyoa4J6m61lkux+LZV4LiNJlTkW0
eY44rBHAr/bPgWfenD9boXvr4n8NR3D3Gn8Ey2+qhVhPu35YBsYBNE1xHSSiCG4M
e4PDfHGD3w4ieQ1q68hppK4DXMQcjK+4JMX1jgENF+4Ms9O5Cg5HK0tvEKHgVuWz
pSLh/VAVQO/r6x1CrJaDcXiGgvmICW751vQT/WmgK07FrpMsbIwXiPDGnOjdpzPU
hYWwkJPdYEv4M7XYQn3Uf1HrMjH88TpuddPdN9/RK9W0n6t1pyIBhvTps1Mp4Od5
jfyftB/yzIp9Y+cyTNJTQczEEVjZnnrFgBdz73MLxdKr0zAa2q9nsxPW0ZfZlNjB
bX5iKukG1OIUbyAENd12ORaSMgM4lRxRYNSOXv4fXu8RK03i5TRyR5rT0ygZ93YI
9fKSiVm4HkGkbdp3XMDvjsmM/PGscBNDhjmnSDCqa075TX72XSHHZHTSd8PcSjM9
jV3mZGUOtkjGZOnRahLIKaikWa2tm1XEpfdRbb5kOwCuV0V4e+kscP9vCpki/duZ
q3SUV1a78uG9q4YRpvhey/GoGZ3CY3uQoVzcwazMozEhfv5BwSfiXhW+t4PtVlP1
2EUx3K90mUKQ3YhhJBG0M2c2r2UU0sM6H1+C9VBRRFH97vQU8hlXgcLwvFWoKYu1
gtRGiG9vBXNFQorQaGE7k/P/SeTxQW0fXx6s5gNZxa0itTY6UYpCbHlnVWtY5qKH
tGPMTk9MzcALGonrLs1xlXrIjweItpFr/TIgmYSrU3jx+gTyK1hagvTvirhEI3+5
81idUW2AeRFh3AQggnAnZvAVYTnooV3yymKOIA4M+G4WI96mW4eRwVEo38apjvDY
cqQC2Z8cSJgroLvpC0fsZTvyshdo24DWMRkOx0hb7E9sF8K5NxOwzNFgC6SGNG+s
niqCoWztVeIVFDbnqNYNAXA6bYgbu+lU3tSRmwlvrQQFFioO2LXdM7KGcW/IBjqB
022xeNwYXbpxgzCJjFQMgqVI921rrEkM/Ic0+sd0PDR6TB4YAa3I3Qwqzo89pmlB
1vVCFNWUQ6wNM2Bgb4/WUk+m0YLcIUt/wVrsEGTPR0GkrZ1IHfZkBbj3vEuiYkab
EBKHkWrzmvtJBOuRlWrmlJwidh0ZDo4BKhMTfw+krYqG8PfZGi/KUAJ3exaejSvP
LJrNka82Kj5WObTLskaOgSXsPqFybMKX9PR8kxGLuh0GyH3ZKxN1820xONNPqm36
9+8iAIoAVajEr+BJG97D0vxUgLKo034y/yQK8tdd+ZL9ze1oXHDTsCtcg4o1ntFP
Q6opYoUua6W7eAmMw6K/2Sffl6QaRdyvC5ZGURJ/r/FwXVdaSJYbBmC5pc7UTFJ0
1VIza3OXHQDDGgHdE39BxKkqZYhmyZluGY4gGHWhBVHI/gF+5hCjkYLxzFc5AvHn
km28hUrjS1nC1jJyHnKwbBRlMszfm0USh0VF6HgVTlTMLY9ufshuytx3xocurdZU
hPQQfpX7WrI1etYFJ5ljdwYNPYy2h6CC3pxdoEnKc8nZs7l3QqrggyNIr7F2HZDe
EcFK8ZT1bc4fBIZvzC8KntLnVHl1sO9S9/Lf65M8+cQWQUcod1f9nFYYTlp/QIUU
oUHEe0hSNvsM9DYLS3p8RBK6f28QIh4OCMhyG4v3RGlmEDFcUEPp7XeptuxcLx1K
PQUrdxJBIdZ6PLbUSXeKLa7ra86SScKZk5pw9ZwdjgEkMmGVJRqMji/9oJjFJ7QB
bzzHUDeIH2DJG+8I8I4/L2hlFEEmsP87WFBXnJkOP832jeQka/HJuoyXIioIlked
e+519ANZwo9ynHbiUPzag/KE2MKILyz3yB1DqMCmQZesUnkHUxQ/r/ZMPvLupOHW
6ePWfQ2L+1/iCvcBf5Y6cLDu/ZyMBygkNWo9vp5lGqepKP1q6v55n390eBZ/41+q
`protect END_PROTECTED
