`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UHMtSOvylu33T/QXZcOH8e9u9KK45MBWnttWzrNSg+4uV+ktuNTWFlgJXUF6T0G2
bsBdzrih7yfbaYrkddw4J4sTRalBAkFg8tHrG5sw8Jf+RbbyFh3uUGdyc0SwIIu/
eb8DCTtCAcvfL0MDUEDg4kuobRtGgUtUxXR5BberBzrbInf2fBPzeDKkab1cuRiO
cJRN44VyJOyj8Y0UkZcszxAfbJoWuPR0QW3bZ0GnZFGLa7U3h+Nex9HXDvDqopZs
fSSh0BUmKNxmJJ7d+FXLw9jGuWrn0oYZC8B56W02g+IiTPl+B9UylQU71T4u05jU
wl49i5ZQPtNhb9sNqsW+D81xkIGcCw93Sak+j39/z9xeex6sam1C5YpE0HNH518J
mYsls0+Fm7+ZprIc+0LhenXlIbJp5WxjjO/pYpUEyRh6XMMwmGVKQxJFTr8kwbQU
A/YRRQIE4Ol7x9QSFUzC27AQ91fYFrHyb4HrZ4cQuAGwOJtkbhwqR0YfNUx4OTRm
kWaykSArHUkuJJ90412JCx6WBc659GGQPb3dUS4TK9zHPRvIgL7Oba0xDPVefThQ
/IuntekxZBwscxdNS8/1lt+Ik3jW3ySLEStKhVY1SZlPK0YAcjTUwgy0PWyEntcp
HUEqfaRLadEfANIlrLUarqu6gzDOJKPwaezGGo01g+TauixRxJmkBScC6QfEI8se
+wAeMIOCrCsa/b0zx7+SaWGto1ifPIjougLAEPvMlw6ZlWoeOg9hAUhIlN1bah4N
2ApvtePeFr25vkedEp38dvf1ZjpCcaeuleWhJ/BIlIRM1yT99H2FHY1Gqf5CuAfa
+X0epHE5mRKO1/+uyv+7rqutI2kL/nR+DKsT0QcNiT2M8FDc2FHCURGpswsu/J7E
GlnHglQn+USAo2uAXA2KDezQ8HuBc54suEh76TiD+MZLIcZiT0lQYjPwFh7yLcQu
vtmpfQHEBECVVV8MyvYY9WUd1kwHKJW2MyV8jbk4RFRXML6763DMpFXIwuXyak2n
wFOHAR95sX9HPF5jPv/Nu9gKkaKaQHb7cXUYU2QWlHxElziX4pYzjQoqVRTkGb74
Ev0/uvbNyjQ2Xbuk5f8QaobvsCVU7QGWi6QfvN0hbn6SztzTiZfs/uSQnTVusiGH
Q+2ox1zcIMEwYX/7g21JAEXGCpkVNPyJbPHeCLJm/9UvPz+Zaq3wd+kJ43YaVfr5
ebUdnqckLBY//xOGsXFkI+SJ7SycbTBYO0ilUsVtsRlBfaJ4PNkotWGVrKO4IY9x
AVgtQWqqtbn635zr7mhvF/Ogpew5uYKJLPHdnHL7JUcxiYwcqtwjxQKWiX9wtwq/
IxwFr6xu9FgGeLXtMKNbosuNkN6MaIi8Ro1pTBaG4g0=
`protect END_PROTECTED
