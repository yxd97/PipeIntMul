`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
stkERSL30Ur33Ntn/kMjLmf7luAmY8vgCL+ZbYUNtIQB6K4Wr/2uTvxlVTMJ3Pf3
zCfCqFL78ZuRSouJyZWoorJ2GYpzuCl5l7tvpajnIuHqUzvlYIKNe2YcDXRD/Ajr
E4kU1SXby3JjXxp2lpM4KvW8qZ6hrcg0Gw6MRRGG1myuIoCbXLwLIuqH/sZ2A0Py
NzpGZKmFFj4QbIMETWbAarOH5JTAEQwncLCpMOsjagJcpfCdUy8Yp9QK24D0TdSH
MEyXeK+z7utdJ5u1tEuA2LN3+FECVwUYxcUER9KW6ovBYEXeZ3SSsEU5L6wtskIt
r6yFAtlDv8ODlII2w1Pmzoz4jxkfn2JRxBqDmfw6Rmld4zqcsfP0ZHycwVdgjr6e
uYYYYqndsEbAxacJu9bCVvPqSNkjZ/f29XvL++JX4uRI97E2O5D1ld21YlHdJNBf
IZqD+XU/OlD/Pp1tI0l9beALXMm+wa6NRzm06jjCZ6OKfhsvvdXURwjQJfaBIk97
FH/36ZHzhr6K4xae/dIKH+DdNc2yYlq4vZfTgypXE12TdkrtUcMnewJYIjrnAC0e
dTDppttrk86+S2BRmOQXss8ZjmPe6SoSf4UA52H0iL7T5cwbgw7eN6cBItKIaQa9
MPI1A1Qa/GI0atB3C+oqUkQ7Tgk1JiK+ifD0ZJjkBoA+Zu0pxtXvI0JxnvkmrL1Z
ZpxPYTg0wrLvAXu20PGFscmkKedsdahoDD1B6z1ItQ5UnT1/8maw9OPIvxbXtgW8
8zsqkb5O6QsEmTP/rj91vLQOXE+G53E4XVQklcAL9cypdfUaZYOSK15H0CGNU3Ub
5BcDMRA1WtY9o3J4TGoKhjIXBZtxhz/u+1FQ5Agx77YUM70ioovSpO6aqUXR5hM7
aHZ47pqTW2kOn0H0TOLiTV6pViKyySgk6tT3gSELefzd3AlhwyIqWEHPVM7NMfAl
GIZ1y5Eu1T2iOtJWW1b8j0vykaccPJjsTiX7Pu939hs/cvB7rbHOQitzvCjt/5+H
I/+91tUjNHRw9xDyVGmCxhVGRv714pw0/jnhCs0Rd/qqaRRyi3UHiwbuQf90bqTp
vzoa1h6cu9utnDm4jn3v1NgaRDYLiFNqUpFzLK4hzl1k/UOm8KctuSl9wMMpVPl2
aHKZ4K9fvtGtl4R7M/xf+F9WpNQqNOUS0CyLTFzgsN82r8AsxOyPa0SYHPBQ15yr
8FkZ4fqktos8yTpofKwUZUaDhUBqMTW0Ctn9zijMe7Hxd0PfEfjYyBL/JciAtog6
y63ONcRigiE3cCt/Lueper+KRyabhKGuZN+di1XDeoBRge2PJR49s4Y7/NUhefIx
5pzQp2DABKo6EOqZpDjbV5LpMFSoeLthD7CTHHh/cuwGvV6haHO/RWx2yxsbsvil
QjgQSPqVfju4iRl9J10gMFoQMD8k66LraB/ibH83gXgqmw3wNG+ahZ6Jo25i49sA
0nhc88jebSOV8s6B90UAGVSgkDX5TbFXGn/5TXsad3mtSgIT5ZkqicSr/9xf/qTs
gjtZ639/brgeJGzAXbnGfr2SqipH4/mKk3etKEJ7Kf5Z3pkl2E50mdD7pogr4uOT
d+sVYwXgtCNBzE+Lko64F6YUudM+E3iTRs0O1zm7RvVAFhU/dtCceXEd7qdyvoll
UkfC3Zdby3VjLS6/Bv8Zbn80tcqNi5yf+FGyG+KNi71XU9f5yMxeOAr4HI5gBmn1
HRndhGs5xCBNmQ2FSJwCZcTTK+/w70z++bBx9CfqQZU=
`protect END_PROTECTED
