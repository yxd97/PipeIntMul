`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4bRqc3Ztoz6Euy9CbFKuJ+khDmyrnCJ6V7h3u/TvrnNHkCxzuWfJewR6s86V8SS
T1D421R0974vTItUYhOrSV3lEA6dugtOhQ4nKRnM8k+C6xG9ydZC7JV/EImaNLQ1
FiHpgP4j3A7QdIA6fQrjVKUFJmwWwVMmvjRPZ03/kGfXrEb85lJ89N4NG94ZDyev
OHQrIVIYNe5F5dAKNO0FJ9C5BYiVuuQt+FqDhvKYGziNpN0TI9w67GlVdW1NJ2zk
zdz7qm56Y9yTZZ5AjRb8nQnflVYgFwDNqkmUWXCAzBqwHKjiq61gt7V8uwqmrx9K
ah7SDcMrNGP1ychBLjWWJuIeSmLZNbltaYQVy6ejsbQ4K7HNkNsR/BsiTm9yOXJR
bxRb0kHr0FCLLKWOr5wSDQyUpATK+0BstPPKtp2hR1Gum+Z+PVgJ1Q7D6EL/Rx1Q
60V4NazNd05iY3ZiGdQn5Dn+oi6kFaiM/23NweaBuLbvF5Tc8uj2ONrTyg1SeXLy
yYBO9MWBR+ARmcvXV7iYSUX984kG7pgCq+/VHxdpdMRYxxd4v1fg5Qas7B0Za7ZI
O03BEsjKtsSm8JQ5hBHUSMNYJ7KP4Pri2M4xlJwtpWUQmXRm5xam8+N6hFWk3vqa
J8GzsIxrJsEfsAilCvHkhyI2uR6ZF7nyFEapDv/Pc1ZsZtP4WyCSatSqLk+y5ASF
pZOM0BKnoawZ/Lo7wboSdf0xk+PGS/Q9e+DtJMxiM6JEOAhzVpf1FeYaAwG0nZ6+
v5gXX/SUJn2jsaa0Ffq2SXojnVd0fqm8UAqsIv7zNtxtXDAjdsF1PUN7y5hTLMOv
dnmXyB4GhPBxKmRcy+OeCA==
`protect END_PROTECTED
