`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QzhoEfAmakNW2QGFR6/aSC0t0Hyz3MP9GbtwUEwVTwbv0X/OBjuXL+Meey1slP9g
OOC+/WSBQCLP8f2WnmpSlogIMKPHDUpLWDIiUocOap1yhwXjZlDWl1ip3/e2YGM0
cmx84uU1vWEe01HdWQZex29zkTCXetypgk7Rr1WOsdJc9W2QFJ0E9o6wLkJ5APaJ
uWaHDRlwNlpMj4u6SFMg0grL84E8tfm0kMfIp7ZB1RRSYjL+WHm4WI6qjTZiq55g
P5piImxOLUBe5rvPsGNKmmu6c6urpVg4mE4TkSUXgpvCO9qt0ycA3Ly6Kc7eF/qA
ipeIYJ8rwK2YzHJopg1OpZF6b1Xh/PYRYEuaVKQDJlYP+VLbHPg6205FyvJHrmG/
F7FNvSr7x7rQgT5o/Ee7IEZpfL9ktOoFUWu9LfjKRvoFMJDzaCLFdZrNdSq9Pnmo
1TFbDWd0Q637XHT6D/LoUu0F00MlxQhPRyKHg2ulC09PcIAg73UpkvUxRECJItMF
eWudlyzodqGwWuTB/KLom75PsbfFz8S8cUPLbFIyKeu2/DZMbFcziz/tT9nKDyQe
OdWfZ0SKXZAsqd0Cd27RZGTQS1N/EwwhOm2NY6HjIFFJlUYtXPHCZbpVtfRwbt4T
Az4KvfxcEd6uX31msYTAks45+bbx6CMfS4MUxgY2n01U2rRzjEZuoUbKmchz2l+t
1kbTQguKtshUuWlsJRAjN+qRFB4NbkT+OgsipLV2NC95ewaAV6x52XeWBf/Nb9Lf
KRrqCpUPl5i5rzbN5LEFPcFsa7uh1JGUNCOMZpM/+k81OLdIhupdrJwlo2+qGxhc
PNLu0RH/ujeej34XQIhdMZcfpok8dxl3NmmJEzdRDtfagCKWYEX6+13sxMSeSzyn
kETDUn1RidH6mJzJd1XJmf322XDM57RcKGYQ3UWbajzv94B5fHThAXKgG5SnEnm/
WYgHbW8Epv+IXjT3RkwgK5vAQSwOXpC/jmg43ICmKsQXUqipRRq7yNy1y8FtXKx/
768RQ37G1e5gdyPDeAVpcMv0giKXMisto+FBXO6XYNn1Bx8vL+phyQjwVBBGEzcB
9GMklUmqpffQcGdwOeCsT3M7dGYw0qwdenmbhC2e3ZLeaIkFUFCk5oyj1Uu6MUVW
wULxNb3zhFdSmYBQmC1KIScmu+WXN2hnAn+q7nlZEI9+InbY2/WVeJWe9LyldBgC
QLYgzKcGUQbnUrAIgv5IvGyw9Gj8PFEngqgkFYEsiaOdIhmy314BYpuzesFrhxy1
k0u3MmpOt2AfsqHuIHjkfy+HpFVv3xYr1z1mcb1n/RbFcnqdzz4SpYcgT1XISx7z
hI5o80sm/+RTGz+Z0vnVa0SXJ2VcKbCBR8CgEZw8Of1D267l9IUj7naMFRtS8FzU
dAO/JAzami/TWVJQOzi2M6dH65YBfp81ZS82d7ES68ubrKlIXl/szZ0no/fJJeSG
EvZdmEnJQOBUYuCFeRMVsubeKT2rr+VA4FO2V9nEnqlV7+vHW2JLAW+ahIqPegL6
YofwsG4NkC7vCvilAAHl+ZHeoXYgZu1PdJorMzt+pkgZaG3MrE8M6yYeQxl3T/Mq
pjx6IFgazLnIplbGyxb7V/Vt5umuX40+atSOHYbFZ6f50S4AoGk0tX61EBFxig+n
f35H/T3HqVhEuEInyrojRh2RTOhYkCT/NpCS5jc/CdiYrGSZfwonSwSDaF3iLx/y
scCk204VIVOYnGsQtZhafAtDothLr8pbwEGPxe36fn9UK3yNG+o6unWqM4NZwQLF
wzoyFa2wluYHk7x4zDyl8lSzCKw6vG71IVT+mhFvwc/rLPvNakYQJkgFI1lwv/Hi
brZ5UuyKs8z1scHlUNbKLwd5mO/+3h9MH9FFxWGusTE4rpOJjmPOH7i/H3J1mERW
Rg9JOS3wHDd9BKJ84z+7JLjGxwi+XD2TdEzcPsuLQVhV0J4SRn05zotycxJdqWN7
Y6mXVkmtA2m7SQIOz1BaOX8HBsS2wAfWokjVLnOiEflKJyqG8yhtF0GqGwOQOiny
w3P5tjqqgwROEVTEOpt3CuwpBTriiOl6n64aibHFnDhBojNYXsQWspFHD8vknjbU
v5hMsQ6qSopkBuxbUiKSTSAp2H7nMse8Wf716xh3P8T+iStsNZcli6sqjAfcTRee
1D48FbitOMqymAYyyPUi6E9NqmBfivAz6/SCsWPdkgCWXnyTIUDhVHKysvryKkqv
XxcL1YU+bUNtrfrwngy6Xyqnktat2RIrOvzlvgbbE2x6Rb7Qkf3IgQBxTiFifQ+A
ra35FXP05uVb4ObxWgR+7xnG/LvihxRcoQuO6SCUhQfV3X2Bshv728ar3qv/9YtZ
lJMpCpx2bI564iJCJHg0+A58vRlVNW+ky8evxXXeHF6WNpT6wYBl7X1YXHOphUrK
CtdFze1Vjf7IrLBn1aQVujIMjwNstEEm1TZpDku+U6LOEWtEo7T1clVj5fik9X4Q
QHbg7+5voqSzlRtzuWr8UfJ/RvuU1n13Fqwi5zp0oDZG3FWvROQQ/oYbAx/rgELI
ZDwPxQWeNvA4jlf+0zHA8uRcIzaobgPz9w6BajMzTGqpnzzKE7lpPJl7Yg1jbRn3
M1BMs/HPcZ2FYig76k1bEKe1XWTHxYKTzd7KuOhJEk6RRgTDdmtvnbEkrlul7rQK
FWDmpz+dpZ+s0HojOv/kS6XOZfLPiaw6OMf9MrYMyykoKtebyg/QC6nUZUnjkElN
4uEmkrKJAKw9ogGkKgGUARQRTMd08NkQZyQIWngPmFj/Sos23J4xZAtUxBJH3ME5
diZs+BGD+f88Ed4AhudWYvdciDRwqwKhYzI0HLdoq/2nkJFL6TM+gKBac1us1Jv2
Dj2PzlPPLfg0cnK17kAnAnv7Vg306r+uevZEm22ICSJwnTdPrzhHLwAjDQQ+rR/k
JQfUsEDoM++29perjfBM+/yn7CnV2wXqFgW3TaS2FjHxQclbpfgIayC5Q/FMLH55
5eVZ6xqxzkcRBHVrftvMGUaVb29QYE3d0/zOAgAQBWCGxr5WZaxzpZAyZrQtSLYd
ybBHqMXm2CSdfbVy05G5POA/Lv5NR8kLL18r0bPwBYz7ETgIBIoQYpCYKfXQvbcF
AokjOSo2CXJi2q9KzQLGNxl6lruZofm6YV29jywwCcOkclggziXyRDQfyT1a7siM
huAqf466iuGmjUoqp0+doM4YckGPMweY6pedHj+NAnsP4iQjnk0jCFmyo20zqnYO
fDl4q4/sPVUIXhxcMlGdDNZI1ojjs4vsd9BUJnkxo86asAaMSApSKN0uphkqYBld
Bi7sT8wGVyIVNIoSYvXjelrTEI4SRjOA1SnbAzFlIPBQW505o/HXO8C+8DHqTxxK
VedBrIP8e7GrDeT2biqMrMJDM49zcSnj1bFPEhtpLvBl3e3x8ZgvbCcYi40du1NC
4AqZyp4OBJ2OhbD5ppty/j6vGUI1ooVgSdM7cCO49fCiMpPXipKXGYVy5IVLSIa7
VyG/aN+yMpA9GHRW1aZOb1KzMSBuZIoikQ4vurSaGlBtOwSYm5glEy3NmvvNWIkV
BLaVGoWu6HcSFitMyvZkCWwXnqrR22Gw6ly6qZT7CicAZxFuLhC1KxX++v3U1ZQw
RNAsB8DGRcZDFbTmp+acdOdtraxAuKnOc17xZpbOJ3xKOjVF6s2e3lq5BjLsgmGy
P/0WuoufuL77i6PGCZ+4GB381mfxAVEPQsdVh35QbsCCIXDzo1+KDkkw3Sk1ERer
rd3KfHFDuZQ5HYUPkzDeftBGdUkxmwoqUa7SKNwSWYibAQMjtwxc6UCp+1VNZyHf
/TwgS5loG5l6dRwm/2+KhlZCjeKljm3c3EHpSKXTHHogglBdjgCAUUR2KTWDbxWL
PCyB8BSSxOTUueifC4PxCFuqBV6nHXEMpHWO46zJ72A89kpVEmhnqqFJmIXl7m7S
zjrf9uvrjUBlMSdnjGcONTa2DMjI60Cb66dBdoUEeOVEKM+aIbDpan8S6mSmsZjx
XRYEwhEU8e1RQh/qRIlwMsIrdBT4beXZ0gIoZO65bev0VhKcweWpjWR7k8ZQMnxJ
TBdsx/R1WhnX/wQjELv0NGRpP8vKGCGzbGz4goYMomIpZrmjtDB6wTc5FJvICKZ3
P8l1PiUm7QyoCJJO23sAUvEdPd1dA4PgIHfjMZ9cMI72yWsRgeJXyy9jJ4KMtnWy
LTRkWBP/wXUChUN2iGvrjZ4MnDg5XsPgfQw/YxU3iFu3o622ICWW739jx/YzT+P+
JI3kcZus8OvhJqbSu/IfPD6vSQgWWSB9lV38onuYAfUWz0NHJgXey4Z2y1wwf3SY
QbIJHfxt4PEhwq9pmHmAuYoRPliB45hGwBGnsdtiGAqb3WVZCUs+mUKh9EBTjvBV
5epR0tRSy0kpUgDveTWCFn4qxV6EBqko4Rjr6FOhVgHyG90i68zmOJo1pTlqCj0G
3XbTJx996hLxO3YNdF/zqHCw/93ew1X0nZg8hrLSrvgyecenjg9ux3FkMcRr0vFh
rdcTpULi1FHSEPLpQQ/II7CbOlwUc9xVz87Bp1UVxGJi4ZU4cNj3/7Myvi2YnJDE
bJkZn5i4G8OS3fRPtzJPPziemNuMlHZangEGLSXD7+UczheZ5S4QY7y5s6S8rnSa
WJaGiN3aJwTqvq1VlXwz94HfjJMrsgC+vh7aAWnQ+cXRKvEXiclbu2ah//beD5OK
N5sV2TUrzeG4CPv0l1qDO5gAiv1kNi2cw2fXbBwzjsYVuLH5oDp2LVp4syUjg23r
eDRLoQYuOXEGI9rdBePRuQZ/wV+8s/lYbjZ4Zg09a4A5Zs+oThYE8JgfhBsCd7X/
tqZfhQ/1ATlC48GIzskGMS9T8Df4MFQb6v3jyAd4ehLqhMRlsTDScljPrJm59fRX
e2uHgKL1pRnW0/k2tcx+VZhrL6ABM8CxlWDulGkgBALrPZWZs1njpRshW4NJbwkl
v+HfHPyFL+zqpmsXorS+hcI8PdC4z/QjZbFhO+XbFohPGonKYXFjc6cblykEDziV
bvTDAv75TKkT9jW3eUk5FQ6YTEhkzik+DnaqIbnFXYWlkukTc3KB8oGrsR0hvcpM
y3aTnVnss7BYCzc1i3XiP3+6dq5vNiRt2s0StGAirfsKBP1z6PfxYCarYlWL52OC
LlEj2LGuPZkspZZQMmaBvgGKs6SryVb6hrhzZwNkFTZDTLOEhXNKGjFymYi0CTq5
tonrx/Xjj+//rh8xEer3S70VTRfsBdWcOvZ9zZWhsXq8mds0ZpnfqFjhBkYLXl4P
EZkcish4D08qa+8CCpWhASI8keaHSzsDDYKMCSzU5Vg0tmPqEK8kG2ENoj8XmhXL
7+rZgoMEbmVcyQVS4D+Sbtf2o+81SjbHr1iVKmqQl4p4nWh8qMa2Y2xElhugjjz+
8FfNTct2GkVxVqMvXzDHYnE1dzLQ6Bb4ZkBf/M+DqLmgtQvKAmhSQDnl4zvWhb0k
PDCKNWP37rYYuIztjRmX1N/0h6saWSNF6lBQNv38WYcdJRaEIPqAkhBqcvIX0wwy
3ypVy3Uc9Q3xCyP1likm+QPAksUjJEnVeziYc73wfxn5k3XHi9DhU5OIncp+HYd9
gtBDMMe8h1nf8zyhqRlWPHvvJj5WvR6fkwWAeAhdmr0FJHt5YRrB2wPw8zHrWU8R
h9/p11/hHGXAQj+kZGuVQGpF56X7fH88OpLBVTCWCw6iSYDdMfHyAogOQHbhR4e/
LzGgkHvcwPcTWCb+6r9awEWN+6P13Z9BYHGSCfc3kWtjNB6AxEC+wIHce2p/E4sI
5sOsGSdUBZI1H4ZFd5c01ZCUgbHoCQe7rKaTNg5F7wzi/umZoxOd6z424XyuOuPB
QE034e/iXp+OLDLZ8m9N30ee/P9bF3PcvnmTeT8r+GvaP2Of3wJKlRM1Rcvft4Qk
DaIfW01FJqm2Ya3voTX7NFLdBwbicqxmXY6xZxe2Qejq0Lg2xnHge3bi98tOZtBK
ncuw29n+sa/SOuxwOYxH5Z+pWzgCUk+16wIzrjNOaWPxsRQZMqp1EBuLgQyqQx4Z
JV52qYhEypMWb7dS7hYD03WCWIClmqoD7sLYfT76ZGibRkZqVbtSoLI+6B7ofLjK
+hPzzXMdotJ1++b/z61m/RkdJ3OW3UjERLEPV+PI6rqtZc8iC40NkTeSHy9qK328
H4gnQW20WWdXn4MPV+QrgMnsWCHIbeztjR6IOnHh6i7iV05pzTUCmo3AVsTEx46s
/mW1nXSheg7ti0AqmCnYR8RhsGghATj/iper80sJoPeIuYW5ljrd0Q+jYWQY0A5u
ekVaUa8XSvEw6oJ/vKm7+IGAe8efLe3MCp9KwuKhw365KPlGPd5x2dxoHIrgKNW9
xAAsgrvkWa+ZDJCxDmnLhCYV5G0y06TxP1zBjqM1etYaxq1tw6s2l5eFlVnb/7sV
tGA5J1yiANIUPdN0xpMgKmQjmtxEzmLuBnlc1xtzVMugHmVNvfhOUBJgp2lCKqrK
cB4l22+GEe7hdcxlQq7/jDCmgUeeVU0oySTTM9PL7wRblOZiFdarkYGQB6F5XUWD
t9RFln8e/udhlRGbAccJpkUFDNcB5cVjmdr8gtErX1c85BCRxWWno2V0Xvz8L1hC
L30l5aU9HcyvWhoXSEQn3dRXkzg7ssjQH1rjFsJvzc62nlmkhN6tM3C6KKD5I9BG
XLpzkItFmrvoacSmxgkNukAPTVyb4tzhmO2jQZJHeRK+OdYvOgueQfRtvwQjfSKb
BJLSIAVmfe504VAahrqk5GDzKMVycTNAmYetERYd6kErCEcII9WkyhziD+HENXtW
+bX6JmPNGpXTyYNzcl/wavB8tmVHaBEc4PnO+lqaCR1ySD/rFrFVtzZ1C+2ra4S0
lqQoGnsgGFOxeeo7d268moxTST9D+TMaebap5XT48ZrL8QJMDIzvDwgfRx8ERIXj
omymE2Pkb/Mms46RiHWfD2GFqEVbQMId+5OyG6A5hWLEIuPOPnGFRTs6KFamFr1G
8DMdnMeW5Tdi01cwLuOuI8bWDCBj9l6CEbeKlHDnDJ/oGr7pdxFMW0tluzOvduPJ
f9bp5OTFlfKw2/a96/uATRCI5wfgXcrw55LN7C4zffcv8ct+F/yfxjYrXSDKh6lp
DJZzahzsgymvwXczhqOp3BjvQVQzBHTRffBpeyQRF0Bk/aSOdpg8MYKKFhaIeFQp
jT2yzRXc5NUxh0QAoZXH9yQ8ivwsj09zyKwGFsk9+Llv9hlnzxkyQr1Qs3Q7dCyz
Fg+vHgHjBRrnmvPRTidVTRnjQIvlFgYIF8yzO8THWsehuoXKfaOIsAbkOMSHgHrS
nFbW0Q930x/LLaCRZ30P3DPjOq3rf9ZhHHu5ubRV4eLA524WrZ6Z5xiR0Rd0Gx9h
pbnFZEMnJx57OcqIX0bs8kx3T8WU+nAsIdvm9rqQQtBc3B8qHehcLeiV6c9u+tVt
VD9uiFPfyd1XrqJDcFsdY81WhR+GVP1yXuAU1fxA7UNLpeKxxkp8xr8TCYEK13ON
HBTScXR7wQiVWz2sKhCTaQEywa22MJVZta61WsvaqWUGLLxz46ishTwLpyoOmabX
ejqbbGH9aiyIyXynp3SiQCcjiqyrgskL4M+ndzMigZ7Z8Ug1QBNlD3+wybvF1llc
Ot5RclykmeDEQHG+4szHTq2ue2TTO1iEV7tzPbKGwuwF6EK+BStvSW2i4cqt9Yby
jhXyjaXVz+iqXKhnvX2D5RpVFilYxIXYTTec273RZX+Cs31eK5gaK7r+jSAQTcya
FXwSADpsD5Sb1LKNpa1LeI7EFDJOVuCqeBJWcpw3p8qZ6EwRFMwOet/2A5/A+kSY
vKAxKoKCb2w0bPJq7xJyV/eg3R0dcEBQWEITzLzPxvNk+wmy6Khm1ix5ZaFvxBrQ
ZzzLx4LZr3a/nIIX7dBEwHmZmXEF4Lc5fO64Iwn/oOyebmMSenlXuZAETS0eQ4pJ
mi6/iKEpiokm12sWRa4H1cED/8O4cKMCSTaituGA9GXLXt0zkrWTCg4AMnKG8p4Z
teAxL0VQ9NV1US/KrW1e6yW8fgfdzwnTxno5mLPxYFFsXZ9CGSOgnxM3cQI/eQVt
tB0ujoD7AMLsU0ZIJR/MnjDz/0oxjtn9MKGEYEbhkOOtBkMTO9/Wws22gWwy8Yt5
kDz0PTqiaK+4e6LBbexS8NYui4TUioAxmKdAvar5KOhMQX5MT1x9+L1rUS3vkARS
Ih545YkRmoDHzZ5N7EzDEf3WxmFnkQlYLh3sS3wjsjdyIDAZjlJZwbv5HbW6UyCe
w363BcrTfIBaTBfjHHpEHb3Z0Z36NObJpmGa9/Le9ScZWdDUPno4Xxu25xeve6ar
tSIdHJikq1ojk9GH6EfdBCwgMvkq+y3Rlr2MUbSQFJBFNI7X04jIjuY6THBfw5H4
AB4RBJFwQb7i/8JpF4GS5mWpY8dryFakiwlojSvZYPyX9WXfGflHU+wIGO3Gwl2Y
NyQEdXpryrR8D+qpbWPRmjvdu1eb9bwGERW7jV8ULG8ZmF+UVvJoRoLerXBSCRqC
ibhQjyAAvtFFKM4u5qFN8gtd075GMGur+dC/V6Yzl/yCnfl85/ownVlklDk70HC8
o/wyPeWaaqvaodF/ml0pkawGMMOJuWoBXMtt9pV7jOurkhqNEV2vj0tBtb1hvlRZ
xalHhK9neb96VBQGuRUbcW67ryVdP/bux2csj4Xt9IQgJyGs/g8i+54Cqjipg3e6
mtDx8FjgVIoQFkuZcyGBMS2Y74auJNVfqKtucR7eqfS6719/xOezt2Qotia6QCda
/thJZeqvulhwUcAWs2g1BpURXm/ss9ECCRhszkCyMwXYzReHeVu1oE/zQlw3KqXO
F6d3qTwcCbleHQCPI8yPivNfaZ1hN/lt8LVWQhMM9WAijWYSZtGG3T73/jf/3HIc
XLJ7XunNSgdfGZLsNLUHhsA5dec0M0mz8O6cJdgKEsGXG7WPuQk4HLmTopAfd8LX
fa91oHKuXeDsbILE+DyTjlTVJm715mjh8aSkSaO61xfO1d8vNvQ1/xfy7gbpeftd
07ADFdojdheoeFCV8ZPOcSJBxS0pOU1Ei4uI30edNPg9r9rXAKPkHQP0rsoipmex
E4Xaw+Arqe9ZOer5vxp+ugFA65MlSEkze0Bxmi52khNzBpHxpv4hTx8UWhpWgcUR
h//yLFlVDrl538bsm5tHL4YObW2p66QdoXYxnfNp6Iv+T/AcDMJPv/klwe2x7OXK
h9UErtVk+OI0jhWh5i/p5kPx1K+KerW5XJxvacvTYSaTP2YuJHlpWG2dUcTaRQIa
NTeLkcuXYrH+MQvR5nGDd98j7WN0yCHNUzbgP+HuzsPICTpbptbVrGgGPfNvbr6Y
GsMUBf59frfUBs3oDbe7TpDkqrLIyk7VEskRgBiyctJnz945r6HLV4cX4ahE61v1
tP8tzLGsgrM5ap27es69xa2ap0KQn8f+0pDkqsxXYjRSUwjxYcDqBRwkwxXFucQe
DcnVQXRMh5Wi0yXwgcww0zqFZsjAxx8N17vi+FtW3+DZ6AZYsTpe4HAWsfC9cgQ+
Oq9OBY0SQKfYhpBh6PqEZcQbhngeJ6kGLkQgM65CAi634eRonjyC4TFcvNqogf9/
9eLQ1+avytJtIyFjzBh2COGM2KCufw9OsAocfCCWDPeGO90sXOoQwI/AOY+wQrMz
XHQakP1XIyYmNkbqZW27PeAbPu2NMnRbZb2sln+4NTCw7RsUpW9mbpoOxqKn4rP3
WjmGsVsweRkDRxzzV/EG45H1b6INAyDmgfn1xjglMw/5B6p8/PDKCWhw3PiGO5lV
wdjLcdk/hxIIJb5kveRzQ7S+HnmEH4G9bA0t6w24A1SLHN83cpgg3VNZ1/D2DTjG
bp2DrVT2k9neKnTHMAhMkQQEZgRG5+EB5iw+lPv5dEZxflw8LGgYdB/n7kLhNd4+
bNNEy1odBt/5hJBWgxzkG7Ao6y2lEqiX5gJiTsjWbelNP9TIBhfr7bZwIccJjc5/
aNy0Fu62FaKA3HY460PjR1Sj6UBk/pL3eERtCJS1U+x5Z6HkR4BAMDBMJ7mrrJ05
CvWvFLPSZBd3yu9oSMzt85jYqP7OSOf3L+W4QoJG2og1/TX9IIhODTa3indLJ3ve
ga5Fc7OInPm68kj5OSPcHTC4qwKo3NQ3ylB03WqzYj8Ivf/vAnPJYg0+prusraEX
QHjc8YBHApYN2PgHObhRB/9m5Gc/PujDQtsLgffEQI9wtpBaYdSxTLZied36QztV
usNWV3Dashg9yEfKNOVEL2aoH7chhTKCBWTPqQ4TJ4US/+RbftNKck2Vf0haFrmc
CwKFUOag6Yxb9NiCkfX9pIIAF2No7MmSHD9DTLBcInhxPwD7EtMS9IzliiZ+ZsTU
MKgi/YALfsi2RTCDQeKudrpvbw8tucjwOWA5HxjUxnToAzA8sg+0idiDSo4rhF5e
VSMmvk/IK36aw7c/lHK7ou36GX5zG4rCOtfyNnh3F/ujA2j7jPGwEbF9nii8p5Pi
B7yqBkeycmYgOyY119Pj1YVBgpAv7tCWzU6TdLh71Fej1cptvSTlJrZtbNjjWB//
qOAFbowlsoo7IX0d/q8yoVux8VGroiX+UnVXfi9482OszzVlm7LnufY0eqNQmjE2
Q+EUtVjM0LIvPV6A7czxlefz0fmxjk2PwtaqGGvfDKe6Dz6GE7oiHywG2qxzzEKT
C7VK25jNeCXHURfHIaE7vdkV8KtFSPLqzEJrzeZ8Ch4+Pk1d06JKu6W0IH8dO0/8
b8yIlTBd59aScYbmunZ1kqDHNB87RXyOYhhyKCM/4qVU6Do9MbGy8y3sBx22rxgy
nZY0kQomWD93L2ls4U21GbbTjuZzSrc9tCPRm0lphWLwnaM46WSVpekjIT/dqpf5
ukPRP0nW/MR1bPnT+w+amfPlY5p4MVohja/7ib5Wq5fmXlSm+ADi2IN2sxiVATTk
G/1BpQXhJ6ros1Bl4vg1n+S3OBuS45bHr3sK+YIu6/tIlyVETORYoYZqd14r7OM3
45Psyg9/1tScbE0uq7x5PEsIdcX7t+7eLVHjfcGwZo+b28cjTaR2F1s614Pmx8bp
fpHNQsE2kKIjem4fRVGbhoH8228Cd5xUVb/FbfItqZO1ou9w+SP+VGuomRrNayfy
T4Ri3mAAALJKSCB3BPQYiOCww95rCSGfOZE/7UinDyxRpJHiZehue5LQl/PzzXmy
PjIVF0+qitzdZyNvrSDOWshR7OfUS1p6afY04DBZa239rDu7NIAAINWT7BRQtYW2
kaX3WE2pjpjCLBmHfML2c+4BxM779QdqH+fz/Dt0zQIXu4g1sD9XDqa3ZUdM0nkK
ggyjZf2XgBfcggfQ42oIeLfSaag6f+YuU+JjQbLKzgKbiPn7xJfeRROkwJMZJ+U3
UREMb2PCCY5hXi/9JLc6hHTUpzqIRYoq0gK01iOEphbe6Gm7YBv1nnUunaEdtoA2
aBUAkCCg1urVclo89CZPa+x4QXFj062+lXjTDYDHablCAD9FIXfcEEgaQ6ZaWUoj
rS59S5w1KRYxxwVOnib0bZ1/m/cO9ieJhI61vlRggX72SGEGb6h0K7C3Jnwcb1Fd
28S2teInRT1x3gup+YQDWeusBlvwFCIWW7LLqSmQ2ZGUPrP3nt41glClp9L4HTcg
MBbRkIVviXKjEHYtFrSA5SkqUbH8g8kY4b5w/WfTA925SUKnbnheMZdguA2PME95
1ljx0gQrw7M0n4EaFK2H2ycm20aKQB9XS+0d89Vt0TX64h/etD9omrBGR+WDEczh
1huwx1ktxAfiia8e0q3H01u0rhDjY5ByvxRXW6LdJTjJgrgJXVtRtIm6naxnU9nG
JRIaRYHhMsoDWi4fIWaXgau3v5ccT1veHihASK/sEZ4zg65w9VFO8wR/n163wHfu
ssFRkToAGmxrMIDCtMox5tIYte9MQ7FzTFPV7qb6aXJuq56ywe5Cj5gtGktN3+gv
eFVrOFUp0PF/SfhuLd8cI67wsK/qy6xA21sz2XkpgY1WQ0rvPRlKbajBAZFaFxhb
ovI1lW0aIH2u72AOxLpyDosNtsXC7UTUjAfER+EGrCHZd/q6LfDmst46VAtOxpla
ICXOAYsbhv+r5slv1Umn5SAPQJeifh52a9OeGjgZtn2cDwJelnIoAPfkUXEm5ovZ
zXOUeiDs4NrpdcoJirLA+g6rIn+RDYC+JD2Ar+2Ywbyy0RXqfIzIU4frpxnyEapa
RS+DghKWW/HfUqT/NwYp2hokoNjEds4oUeTD3TuXIC/sk0pwS9auMyJBTrlscg7w
wD1n3Z43GkexINsCsWzCCeeKxRCY2LgtrDEQXczdwq5XeSLkx6yYkbUh4xTvxhik
2peBRcc+S5zOrupibl9OsML/vn5+VILJ7ypxdlpVUIn0nzAZAswUZ/yYlFpHUeFg
ZtUZAVX0ICTI3YvDfozdSf9A88r4TPRKjZQPaufNaqIN5RaHSPYtDI1mXXQ6Ii1Y
+EXSugovU58Ty0oelrFyf5s9cX7ON8sSubvFogHMzovplK9qZCYOFNHIx14K8S6e
KSq3mSA02zdBuMIxAG7ldtaIFzGeCjxYixK8QL9ELnofMgLFtpVKdw11JMmQlPZT
VXZxE8i3gwP/il+UgddTTRlTsI35YEKypi1TCqpf+QLYawu1yhJtmDabwPUMDW5a
T+lmWE5idVYiHWM1FeUkx6GguOEs9pHfjZy4R7dq9QuPxJSiIlrDru1rpfcCMcnV
/PBDv/WCgN5gWCizRp+Zqqb7qU6BPvMb6t9fFgFV7DrUnrU1deX9Dq9npYCq1lfs
Jz9z4CMRTPK/h87L0KE9/P8QL5kNhPx3CHK0L+8LNDteYRrn3e0sHSkv4XwvBgMW
xK0930aKE++2ELA27pF0YKhlAwwKPuRCchc67pSNSkjqQdLaAKe0b5kwhOdN1zp+
RZyJwNNQ2IEsbxRjHINpAmK9ZzIIynRH0lEeoGmgZQWEd9vsdnU0XXYd1UK5JNn2
PWKt87+PJ6rHThZdkQK2PSZ2cIdUmXNGWC2OTHuor+xB4Xz9hdB78ZmSJGOtjdiw
grn6s6yRP1CMqFP9QA56ghwDsp4egpEQOR9qodaM0P7rl71pjOFMviKqaN5f2DFR
aGH1ulD4QQRHHMSFE4v0R5xgyz6TcfJdqUA4++GDbczLIdDh2riChEniXWQXKSus
wSzdkr9lah9GcL6Bb2M1ma9d8oX7kleN2ZXXajZgqffzf9lLTIL/VCNtlT9xHO6M
74UfPgB8g8tlyWe2vPbEOfle1xB6eXDM/ZMj1Jg+K4tsCSgsANHhRKun6bEUjSpd
wOu31J2OkaaTXI6n6P3gpJ2JqQTWB+EhzoyQ3N94UAmBPYhE1oqeCc0VttgG62nV
9Zi6zuJifrROhFkQLysmOc1GkzuvX2geOZf0v6f8tZ5XnH3ZmvJ4hV8jKx2Qf+k6
T/lWxxQHsDjIMlUL9HrxTyFEavGF6ZX2h8I3z2kFcA89jMYczyVafXr1rAGOb7GO
E75riNjpNC3jkRqBkij0yKXpp27A2R2/c4s3GPLapREVleyUPmA0YT0yFgyW4FZj
6BvUugv3wCD1IQbEiaj/recrgD/PGxIG4jSpVW6nRV44NQbcUo4MvLaJpT9WbsrO
X/nnu+/kMT3ntJq65HjO5G4uE51X9vtCYBYPPNRYYP9/r2ke+l6b4UGl7sN+FmKj
+idfJJ5RoQ8UpgPux4Yv7PqGcmSb7wvLeuPIZksb+XGSW2yqdg7o07NAMQu2rj2F
nolL95CLqc8cagZecOB74Qh9Fj0U6z987e0U2/64dMYMi781hkJd7tLzP5CycA5h
7eUEEDToOzyl+mhb6HRNNUjPr1N8kBQ3evjheAkjqCECfxP1na5vMkbybYE7YguM
cILA7yTZlctnTs9Jv0BQMGbFn0LoSXYHNGxETVwVx4V9CCpccYce67YkIiJxTsmJ
FEN722TKQbHjlwqklDYd+Y0v5UWS6boyAZgc8HcM3YLBjOP8B+dqVe3ZkpaTkvQ6
3JnLLArl9POY+Md/QBT9TgJl5aJxboksvup6aE5D/fsYTwNBrGWEVkJZ/hhlFU/f
R+nN5h2QHbzt2laFofQcXEchaLsbaP1PZMSxRWC0oBNRN7EtxbgMHxx971K8Yhmy
yGoCTTWRpKDZwIabQ7Pb5EabGslmGJ1JOXHKEu2NKgXuul+I2KrtR4G1D2ToHWyX
vtZdu9WmZE/fVFf/8YUIaUCZRMoQ+uv/AxYd3fhunPkRwcVVLGJEMMiWdRwkF5dq
Y/39JFBe7fM1brksvMhq5mp/DKG7Ed+ZTK5wwllcW54xdHg7tBIl3P7v6bC7NUZ8
ZYdopuNt1YsdogpaJqZLEqy7HT7ocIdGXOBG6YRvC2UWL91l3+8/dk0ZU23/oqWH
2zUBtJOjAy0RKxdsrorwq1Snil1i8o+3mVcxl5P4cOOHV5cM/fgQKj+1o3FM++Sk
lbqe0RlCY5DF0wvcHf0rQ4EiadGPj+LZXR5yrRQMm1Fi0JpqNvJxqyNJvsPqV0l5
xV1JIsvKlIldt6OyXcZjgeDJXpWsrae2WLFGQDRRAhZtuyrKa45weIHi73J2JKMd
Klp33fQA8B8EEf3SX/U2DN/xkaZ4YBKyjWQYS3ZGM3L29zo+8xHaJu52DWv4WIuW
BJ6DnNZq2TJbbXpXZAgRqUe5bXO3M9cSKjE7uKYlZ/aFStXgbY+GbUI9x/GrDKAn
BtkCOcXoQZNcAFafBTFODsr6R4vu4vYzOx42qmXHlacIZwg4D2JU3dwkqbQzBiKJ
sRfZoDM4hZ7G7mYTXVh17XnE2QY4pr7NjXzxIv426q1ECHrEVMwVvRxOA6P9yWBz
84iG5T23BygTiQISjMTmqoKwvyq6mNqJPSNE3CB9j5wdGk3v94/spH5+hZ8384kk
IZFhpTqC54Za85f4LKQnCrEFbmKjflcqFLVb0Zj3VX6WZoJEzUe2HypmSq+gOQfP
iiDn5XDKVRBI8vyPvOdeNIt+kRm72ca948jR7WNWTz8Ctu26rimZyyPVRYdF1j/4
EUC+a744NAB0J690KrIa/DwbBx00mzEfao+gcF2SVvnuIBrzhmFqVTyZQUd+okkZ
f/nooMkpqX6AHfa61TyIGZFebyIgeOoE1pDSkGfRXjt/WGr93PmdKYJlT4Z7aSag
l6dJtJW3rKsXah5nKqcjkyRhg9ETyW8FPGU5d/ePhRkObYXWFXpct8n0aAAJ0s5P
xVdVNKx4uSdLi/JmiahIiyBroioV+Pvw2w1uGzQQPaHXbmIG7CXvPnGjZ1IlEi3s
xi7XZPSLCAi4+OrmWAcOnqN1F6BKBVRRn9A8iidZI7RnELycRwbTUeBJCgy9WkMX
EOksTI+a80Ng0cUJHism+aARHkRR7GCaWg4AiqEbpGiK4n3tZSNOb/U6cDYB1g4e
kd0flDYZLfOrQ3SVqxY65ddt/MDMDZYWHAFXmXjNvKS4CVgcZBljxQgPwvxCZSUu
NoibHjp+T5F5vCTez4QddPn7fNoiAQytZuB/610OEqEv+JbRunQpKay8Syilqq9f
vaH8e9aGegzZwXnsAkSdL7s9HI4y3lhYmMFWOkdoO8i4p7QNAXgJIPEgQTKlq/Q5
FnF5xmP+FvJz9UtwRf7sMPkj6PKjvyGlvcL2bgMz40P0wmyqrsLFcJKHm4mzmLbU
d0wjvRsWP9xQRlNP1o2RyRt0KT7fwlXJYVpc0Z2CXaJTDAEoY4n64iQjeRe9ePYl
SVFcpor2lHbj0PL7O6AMvVB4BCM3ePd5XDZw7JUwS+raaViTCDjG2x3ivXyTWg5H
+VCIwqRl5vk+DfWm/u8QFpr1ZY5/4gqMkRqRNwUaXkUmnhvJagT4lckK/DfpNz9+
qSdPhP5h3FxcC8HvYIqgKf52d1QDf1zLTIvKDFMiwq1n9Q+TI7qSlS5Y2x8NQEp1
j2PgB7l/fOLPgPlmphaq8C8oITnT1LHgjVp8gqf3bwAkCfwaTyH0EIGC7wLGCv5N
YWRePL5AXp+SEt/pa7R132r71mPdxzMLQH57qf3dlme85tOrjPOE60usn1eTqTWU
NtSBjUHODzpT007ASfBGZtqqFQUvhxaMIhhcdcd/A6Lg9phZZnr7K3f+RImXvaZU
oKoR9hTqQTyV41TKtmAmI5yWmlk656BSBO60yI2S3OwtkgYp8Iot9jbT4bjgddqG
/YmX2uikQ+nlqZ/HqHCbi91dRO+kE/xfUsh9hl9uV1buvoGyaD6mpxvqVk497haq
3F9VezuAhreuWhYq61qYN4t46GAVxbxwVBt6tUoph4zl65rbMrrTuwVZe+uGWiNn
SPbhoccCQpG+EE/p49taA2TJuKVvZClEAjHqsAqqcMNHjtiRvZrppcH7QzLhD54M
6qedxgTum2c7k8fI3pD5+zys4nF6kmphrxRMVYHzJsirKjDsIN14p4h4KuEyC4Ep
KKXySMCle2NjTCMvYyFWSJg53niulyrNxA/IzJ1ux3YcJTcGGa+d9BD165nsaZ1u
JcOVdw6pL+t8NvCXyAvQRPkDWfjCTiqLDHKAPaN3fiInDkYlscK10SHPmRe8UEdC
yFW1FpVC7bAJ9AQSDAj/JUJiq/XHj6MDbvvhX/WS8zYa9H/LACqR32Eb5SDnH6Y1
0ix5YzKY3RcjVWW5bmDZFJXtMOSTDjvw50N4u0S6lNzfhKYREpf9G7nKK3A4vA++
sKXXeyHrBi/5NT+VG0fQ6ZTTaIJTkojmGDG5W9pn7FvKHJYA3KeWyo3x3/SQ7PD7
7k7AYcBSuu4EJODJ4HJHSoOMMw6o0BZYPtqcWD6Ru9cWVUtRVmnswOjWPtIRVxzn
mC7zGI7N/YtNBA8A7qRFD/X3YRIEVuFTMY0bSIyeLet8OR96T1CUeeYZsQha9a9r
jOC5XtldknrlG7wOp4fJCbxDd0hXIp0FXvc86CMz9Spbj82ZjAGIcnkCrsuQhzOv
YnJrvbTV8n9cv9ouPr6RNWGhJlaB9BJoGYP5s48CFI5dfV0UQye5dnC/UxCReSEU
VKDft7JFhbNwjRTA3A2A8517Py+RUEmrSzoLCbQiALlYiKyQF+9LKGlrqSZB6jPA
uMO7n/7V4czJQ24cKupNnYbqu63Nl0/rutPDmFcAjJXhC7LodXw4ABW/233MRoCp
dYjSiNy+6HLRhebVmMG2i+UamJQv5uMS1U9qLuUPq1ppxrF15XeMzD/nJVDZvM2Q
aU4I3ZhjIWLuaM/XDMOtGkm2WdhvLeBhT6I588LImn0KuneMrHd7sLRrdO7bEwii
ja6FOqnpMiCz6fB9DYDYReFD39UXa4VV4fljQb6+swu5/SX714yp2wYuJDxsHMA/
EYcB1eQB8z2WKOGEL86KKcm1AOEt5DpPP8GtHK7/3pgULNYdBdRIregtJO1og4L+
Dgfts7/0k4ZGmXMdObgGuZ02gyhqW7qqzjxlQvAdsXlKBFdj4JTV5AP/laflgX3n
MGwIQ9zhYppexIr/9XeG0Q6VofGfHMCaZE3z14Lj53dE9pn3nmKwZYDPjpfREV8d
029V5mhTbGXOiQ4rLJrj8w38xD7XkCzpqZm5Etab9FtbdZxbVaCpiIXdoGfXB6ke
8zM6I1pGAUOAeZbLXTDV0IKxc7Y7wM5U3crWu6W8ntkIw8o4+RO5vjb9A/47WyPY
HHcrC298YxyjTLZ7LzBbu8KH8p4bgfa8ISEa5N4DIaSiga0E34xu9yDt2ZYfaMEL
dkbbNbUQD+sg5Y0IOfUbV5K4Iqb7r1lTfXFjepJXWMii3w9ArU+n536PvN+xAFK2
59VFjfdeT45jjaatEw8XWBMXpJwpvZWPOX+njugxCY1ALrLYdbltVydWZMnFzI5X
TxQIrMIEzrWrdtRApMERZGugAW3BQ8sW5X4ZsIzH3T40KmvieQY3aLZLuUE3kFqV
WajnAPQfKWUIIs2wOB7d4mTWNqxMFfxJcNQbxXMeCFDOJKLB/D/c/8RlNcXNDMpV
EAiTDghRmhnzRrJUUvXVbVafaIjkmRoSLnG6JUXfkGC7v0ATOB0WB+lUoZMDH6hG
TtpBkikqd8darFlBrP6z7RNqizRr1MelDMAGsieKhZLoXRJIWRBqk1LeQVN+oWJx
6z36cvGXwDvflUib3/D5ZG8Y694QBcV9j8bzFFKq4uAZqMdzw0zGeiCAG4QGORhF
sLxK8Huty/SVUU1KvbP88Wx4QA0esW/hnIDBrlhke+mdWiqYQZ+VGskvbdcy2QLc
l/rAtuhJduKNf5cvZ40BGGe17C6LSE2GXvE66dLob65PTPxhYqlqRjDJY47ZOfFg
bIQzwdbfH3cMa2hiHQcrKtRpRfECCZdG1HrzBL7w+NXiYSY/AlgMqpNZ83Rcxice
eqMMZ88fjU08xfU7b27bp8AJbVOEgG4mounQtgMQm1FWzGBveBbthmvyo+qQIpaG
GXYnNAjIHdGVDovTWb/CDYcl7OdWu3iN7Hvx4QyUHn0egei7TXBomBPJa36lxXPn
ktFOwT+2vxf1KV1lESdJSMzO0o+A1Y2spEadcQlg09JofgTgYxP+M1b6Z+iRlGF3
1XQnDvrx4PPUXmhqWKApz+sbUM/9uoXdY4sOyHdZE2qhZ6uhDmWGUt/ChlQhcDZC
ntexlXh0wyD073aGzF2d6LOBjKy3uwETpUy7C13xHxJ69TNFe/B3DYWe6pzuAB8B
hLNql7ZMy2/t+fz9RTkOo3nGZog6CwTafbgD4xccbxHxwiZeijaMiRrths0hc+Vw
ABfAoEYIZGwTwc8MPu6t+jIP/iS+1+pvnCA7wbSvqMgPRU94dnKK38BXWiswfEzx
KAH1YG3of2tPw6kPmnvbjygU2wRReDerrHWAcXpcJsV5vmP5k1p5tP5ir6i3+ZdW
PNZu4dpv82ZjrDBgrsiZBjKCfMigz9QeaOJLG4d/oRNNy+jNHy0vgGlAoxAH8m9i
imgdbK5+ZlECXb7HT1CaijrAcog7iWpD4RxZ7sfzyqP6YYVF711aNDmf6e1Ms47M
P6PEc4O3lXfDxoMFkZhNIhq9x+baTREn+qvgI04LgKbidEKo5pmiT9pUjuzP/DgF
1BvUe3E1bHBrZayqvE1FNaE87Pym9stdC+XjCEOjaUveFJYq3lKE0GtNMiXX+Xsh
rKPpPsXJkUdDg3Babj7bWx4xgyvdhwaYAzxDjKsj1ep7cxTHCEwdmDiHks7ZPX8t
SaN7NVeRr7qvl1Ek6Gj6iuP4bifiZTGKwnypTxpvabbytmSEgkIelZCucrxORf48
TAaAkCv/GipfY6/DlzeBsiH/vG825qYIr7LEkNrACbLpNDFjyKOKvU1FlAe9ApdF
8ZmtWX+SiZUGAhLYUChlKz0hTiLBaUlhgA+/Z/ur2bCVWN8TyAoesv+Ns7+sUl0a
tEDLAaj7JRUa+824FO+5B7/iBKkdGhcgiwz2K2L0xMY/yoq1yfsV+wPPBqiGes7z
hmmPcs1jU2btJMOcDA6wkIrRkMdV4SpAMrJ+0Nz/pAYVxLSS72PZd59u7fKKvxoN
LjUg3PKUa15+wlBNu/nJZudvqUgWe0AltCLRrLkaV4aft4Vjof5djH2fbKBPAxBU
HOMjG+Kc6cy8HBoxur1b/7gmL5w2nu9mz3l/GJ2EftfhlzBEEoNHEobHTUfxRkN4
6w7nUtRphkDjwvh+WWw/3NbPPOJXAU+P1wjQR3e+gDBy3yiizu7RIqVFV0alcZsd
p+HVfVEdxeiRik/zgfxXwkS8LlLKQGTHE+6UP2OEmNXRowX26MJRiXwA9F9prHyF
3jt7RWmfaiMkS0uZ2YZQabMWXrBe/ReiVZmOhSlL+qmVBJQSGCMm8gIQvME2M+Id
aDKj3QIMV0owXvi9JsgWYyxdogaif8ztpiM12BK3o2omaygcdK1w0CLqNn7nJ8sD
Lw9LFrcqjTHzbeJZ2QZJisufH92lQGbe0Ra6w8km6/aT2OAeolKNam8hWSi/zGfZ
LnZYvtGzYVar0k7xgt+9JrJhltxSqOovsCJx63SxH7HKS+niZEfl9LiseNElu36A
aQmOUfvB4UFeJ6fr4VbJ/qGRRlfZQfjKY3YfiIGhzzuGHpFIVv9HIjWXYHW+Jr9j
q/ecPulejcIOgbVjUbepM6TBWOrwPbS3OtZY8QPagfJ7ZFCx2BxRxwlBW2t7HjFN
nalMijVrMLR+Ni6jG3ko+9dEDsf6vNEyvYWOvTKlz6BMQHINliJKvp6cdWv1WPsi
RxxQ3xnmo8Uu05ujwGn6EyVb7MNAvKUdnLVLBWRSc9gXsA+8i67ygAI/Op3Ym2By
+44xESgsQW80tAjXe0w1vmkdxM0qq+cIuxWikGQSXMpr923bzaXPhkFPBokHT7u7
6L/TZlxSMfA8pBzDuuJKS1RfNleX214ReAlQvfKsCjDxgt/ZlaIlAnffP7bZbgms
xSevxkVL/wwvR2G7Mu6S9YmWfl+yOGnq4vIXfmZxM6bZ/QkQm8O5IDWnwhvr+0HP
dTBKNvVdg2w0CQwU/Ow6ashDEa7ghqTtnGhVhdEeiUFAw5WzbkMDiox5SSPjAUjX
DolROfcX6qqQPfOhGMiJw2SQiE7+q/U1D3kpCGG3NVp/vjKq2wJjIQGRQWdGDyqL
3Pd/EeOognTisI7oSa7nW3jsMKOWqEdZjTKSqRSeYGNNmcJF4gzwiSb32a0ZGYbl
zqe5CRCfScrzMCymTSI4yq7pw3EzaP/hbnceEZXOQgF/WrYNjnAWPFMjf1puA7Nf
SwBZgJbZti3hOCfzSnzDdA+aqeh/7o/c6rHT29ugWAgf98nDD2KyeNe+VEGV3N50
qyjf7AhOsgp7V09iXFZWBSjqCGYdWumoRcDYPnDCGan9HNCsZdUR1VwVyDXd/4AB
2Au8d+Ok4xpkoO9xbcQoDTOwAOzFoa4HIq7bBay2mFnF+zVi4HybtGQbG9c13zO6
QHhLXhQjdW8gnixsnNnzAlrNSLES3KBkikh8TVMip7up0TXo4cM8YQVgGnU4JPmL
ND8/h5t0XgOB3LzysJHqedRanTt+Zm9eOoZMLj+CLpm90aISCOeYKzMmmcpooei9
/UzOgKN4N1xh9S8rIdkf4QwjEERA55J+seegdEe473TBuaNaCPYdR6WEv6S+spHm
iCYwmgDfuEpAeMBsM9UAbBknYoga7JquZR7qY3dHGoeNO5Zk1MpWF1QxGH7/wX5O
tty9Djx3CV9KfkyzcSeG77RbjoQmY3l+Dld4jUrUss5aIA2R8/EjMQdHG1JNjO86
IN+lxOKK2aMtii8RmhYNmKMPrbhfnJOyVZ1zTIRJUW0jBwC1S9UmljXjUWzKI68t
FnvV+XzN/DZFBhlEkxLUZj4G8kEGz1AhCiNQFpQeiwIchQfEXg20gkfLvGEjBJz6
M4qzjCTVqxl40oSFsWj3odv205nQiRB4WfJBg7jqY1QTXTY86j7/QXnzKSwXJLoG
Zk/5f0JaxH1/XLr1/W+3kS1Z7LZ2QL7HCCY/pmWOU9yVMn4CFXzGgRKlLp0EZLrl
tOdqIq8nqlmFz35ZHPCGe4BYN9ko8WY9z/MO7yGKH5b2GMWHzSAH3lYzvremp8gO
qslMF/lsOb/n76CborAsf3fZm+u2dfeHTTrWMGkxji8fdwYvNA+mu709tX2PG3pH
XPdnOpkK1gt8fesnnmkcw1BJ/E6N8iYA7N/QRXU9aZKzAcvhuJKUsrjucTSw3W4S
s+n147nJMG+8wmWebGeViJsvF7UksjCyFMwMZReerNF8d+EuIOxa+wim5V23zDSv
eL89LfKe9C3TnYrlIhAGqXVpYchx/pT5pZZ5wy8pXXAgbc8JJHoFra6larL4jL2O
KgIPszpvaxzYHk0MA7hDJXvQmRtfjxlaJs5s6KhwaMABTyeR6iI5rOLO/YR7FsDf
sk8Mt8SSiqJ9PjxWnN43QnaJWytHcDAUwHTExUAztUrhrw/bELxZDIjWPuclbvbB
/gfKpuzL4s/UuhcUYi8ZuseR4nVgMgt7CiyhiotQep/BnpAyG5Furbeg7fNRzrxk
SDIr+DABMzbQuDOQEkDwUqDZ2aSI6XojBj4wTbiKOruvZbgoXSWgoZOylOGnW443
lxul/AVUrhqiYLdd6Nr/+sL+I83wEesBzHe71GjwGPXoSTr37xAjlARicG8TTIOp
BQVUYwY1Ij6L9No4SMUURtJcXSGi+0+g1AIZcCCdLIPsf9b3umgCc1ccZrTqyj8G
q/5L+qoiBOUoNAv0qQO1iVEK679x9t8ERcuQinYUCoxF+NSVM1Qd8wRqSfbv+erY
yL5p3zYd9doXhmxPA0T5ROt4WuwHUu5gUVwilzQUWcAhTzqBadsY6/+OFZcL42Rn
2p0xiVQysw3cm1BNo4Zb62NgEAV5n+GxCupQn3Mab8WBU4n5PnzRpczkagilrRag
87I2dQaumOVEIgHm+1Gf4k0Z00YIR2D8AV3bJm04tb4tyAwxh37dBfcWTv2vfbMg
05Uol2E+IDgiCi8VlUUS7upV32i9JS41sy0ytzNy5MmiH+QuI9ae+clpQO5iWsaw
J3fjQpqN5E8+QlKtsdK5PMHw+HA81ZMabMNSGi+rBBtQe/RjoZtfoCBibkVvBwiZ
O+f34GLC+PDeRkd6QyCk+2A66ShZX9LYqYhp2v3lWF9pzqVCHnsXrmkIpt8PELqa
bi5p57zysKPKMDJNNeC9PcN7Xr9nYffdgwjxUILPHX4LOWDq82MXLTbH7F5u+CuE
nZEyBwCrPo/I4OBwmdT8dB/p00MuSwaev7Bu4tcVi1DTdSyyXiZCmYhnTEqbYJjH
pJgncY5CHocXvwttMF9JmyTvt1K+PalfCm5XYioFpPrSCzrCTta/MURVbyikXqpd
iWp00lN3DcKvJR8JV69cu12oXCw5I+2iX4JipVNlUsq9GOIDyWeswQhX0w+oLlTS
br3zAXVMF9DuFEWMsBImfARXPzMU+9SfchWp2BC3ftpsyxyCJXLhK/qefHf+7cz9
3nG5AnQuNzrSgczjrb30QZ/lhMGzQ2560ViCYeKzV+NGVpmCmI9qVgpnBbzqlMiE
8bwdQpazL3ZL1sC0SOy3kfMwoa0flj45dNZfK+iyj8Cwfws/OIRpb2LP87AB9AS6
aQP2o2UXO2qgpsPSXlZBJTvE1kfITWDO62dwf6tfRdVyEjisD3dbxa4jp02ULxPw
WfEK1SRtZ2dXimU9RJ+Wu1TeGWUbvf6/bmstrZ+zsmFU+NRqtrtuGMUQ69lpBxHa
iGflVMB/BfbIgxBcsZj9TUvgIbTcNx2JqABco7+RHEvPoqWJWfKgUYMfEDLsHcnb
zQekjXvDpkARqL/fenQSeI11fMLcpPr5fvhDzuHQvPq+L7kqLV5Cp2w29RMos9tW
3aO35OHk7aEdFhXeideiOLeUN2PWYknURXQYCuxGUkScej/n/JYf82gghvw6UxsO
HKgFPiBkGQCWqgkLufHdZYxP8VFt4bXK5mkgDRMOfIZbL4+opoBPCVyX8FCxZi4e
s5WzGjvW8u3oG0EMoiXfacTVeaPauVM9VS03lLVM6Jj0BITQeSL6tQuR0sUMm9Te
U96eunw0eBpmqbBLHpb7+VyQ8hm6v76Eq0SRghQJ6RIUKDldtxxwCUGWFz/NolvW
Ac2kmI1diFmCsOKJAZzLMuLUEw6yB7IN6OWdMmjnTlffezRJ1Y1wSBeZJCLm3A7o
FS9XsxzDiU9/ySY3b0WC+BGwD7L+XF8NOYbAcmbXeSr7l18PV/uYWwy4yr3M9zyH
aBF9gPhI+LDEXl2VbVPeCArSMqyma6nPD0M4Q9ETArOKCSnnZ6pdkrK7ntlsBgl3
f9auSfCtB7tsEEmFNr8Q/B5gG1NeGvRKlWd8IDfu28oDd39RQG/g87gi1rET/dlg
wHtCu3Bw/ayOlb8rhYB3RW8A6WMgjM3zJOl+toxxY73rg6if1qgeveLDXodAOtYF
2Yi6ebM9UCweNdosjMfU/fJRLAKBYHQQdermTGMSAxuJrSjPxctB8p2Pyg0cUuo7
zpqVgNwGOuUPJl8UgT4goTCJ6sgyDypJXpuwLMOFvWO4p606Nkka68jcOz5/LeJh
JkIl3IsAdEffAoRqHAcjp8mk0PSJH7MI0w739OKI7GVw5HYKSy6ydb5FE6ZvhALj
NrfQMZ/L1hjljGgjg40v7ww7tXc9kw8XArHmZPIybMw63m4Z48t+97MdeJlBkRgh
iPyLZIuuPErMChXWVejDuTyAWp06t8brYyVqTI2lpeDFUgBJ6eKIlUJcGjgYc7eq
Fy9M/Byi9Ut5lng5hd5zHJGhyHJMLmMJLumCRWiPo1ySHuZzPkl5aGjuWt244jqK
m0cou3aTpWmIzD+DUu6TXxk0Ue1iaqx1j+cVtM0Lr27i5PXL9V4AcjnUaT6WuHc7
FOoFdQ0HbplCjJcV0doVjKiO7iFaOLRalzSNUs24mi76rcJgLMXWDJxkDOjnoquF
bJbeqcRegZHUs6s3JCh/iNlIpco25RZpBOIcKHSZXc9qWWtmCThz66jUIJkhjvGA
YqZaIxbwRr5ssp9hIdmzHrUIP0CfY1hKs3azIxygXVgMp0m+fZHkuD8uL3nbzDxx
6jUYZdyJH+G70qQds6pFOsJ8Osljf602FPEHm+GoiwP/ywKTiod3JFr3dwMfJ0Ua
xIQPXwojiDT6gQ6IM58eqQF69BbmrNDivE3+ON4BqMQcKO0oyva8bISGQkbJQgcy
8HtEPCAMep1YYmntNZquFhAwB5US3HOArVk1efkjafk5YS9PuWwg+5utNZVrCN+F
SHAmAT0okutNBs/r6CAfUSe8MaBtHznpc3xTK7otyxgMoQcVHsamrs0QiuBxkJXO
wUWOJf505HcI0Q6guLpUBw9UWD9Nwa06YoUNQXR1KgBMXGBlFEY5wBn+JiRUyeiA
O03JmZwz4r9ViGB0Jjh7D1LmSnGXtOPxqVMOxx7pwdnET+WWqKL4xw87JQIZUkUW
NXuIP0kvL+aY9g7L/lOu+YNZ+b6tzqDEaIzsCT9RYLeJuN+FoSlXk1aLrLrfhRqM
sorWULuDd1OFI7JRNXPlCJF+mHz6EVF/lzOEvIWz8b/nIZ4WmuQSyRj2Gq+ixO9p
AY5WHOM935KJbEOkOFwJbkrrAo7WXi6MRfnfKQU0Ns+E9Ag8PQ6NbCITwFAW9g7B
smyFVT4OzGzP/enrrwiyJnB7r+ThbhUcBccMWOwHiLWPWqjNbsLvzUpuI2+3s1iR
C5aG59WbzNsEcB/C89yhTEXzRSh+dYx9lyh3AbRLdbENPZjMgCtZE/jUPFxHkF2F
/cs8y0LPZBV+z6fRV8YTwCuyKFR8d9GewNNN3KWgr5tSi3YPN3FqnaX2+iDS2UUm
C32P/xEbJlnNMxjumMaPuUmRONyTY1CiDYrwalLuBFxVwPtujZFET35ATNQ6//ad
u9NbwRod3Z3gDJcckxqkWUPp0QgDEqw4T626nnFQOsnFBjUiZegIXElYXwiLLe2s
YbSy584XoVRHfU9xBqOiTsehTJRkUd1wcMUnMkWHDB9o8LUG1G7sQK/hzFiZkTgS
cEBr56sCcPScE6y4LXeJ9tcb2XbCq0n8SjBBfBVcW6SlGoWv0yEGc+Tn9tu+PUYv
jzau1sRtNrKfqjxpU+lmJT8a86SFUyrH4SzykvlJdkQ84d6cbt8+BSdkpTv5Xp5f
YkYiqnE1hUHiQBJr5Z41zjuDQG+hnknJmzi5FWqheoC7fCVUkP6imLj/7YwamWRw
/NvD/iZGMgs9F6A6PbIeEewlcSNGmyBGlzhykcY94tO8K8KGCpFii3k4XGMXNAmm
Fl+zaz1tROuRBZJkr4GhBCOJlxA/wYkyVK4q150zyI4gG1pX/bLQWooft/+LIJex
hAx55IdU9i/VIY0WQoa+DiS+GZHGxgpHPRA/cOgiEa+9PBEuULL8RKus8534CD6/
ENKAMH6IfblK1cL9mwJSzD4rhdB1/TO+5DRSMoHvh6Wdg6DXHa6LP0HRScGaaw7L
Duy1IBUWTMzLRNnU9yzjDqe9+G0XU9Hy1l39pB+17euyCSZuh39MT13fGnAQs/o2
18LuGxTjS+l6sGc3Mwg1TvpvR7NyITdCoJixCkbER6SQ5vkcdwcqDU45mWz0ESQQ
8OzzAz36/kbqtKBxRfl6024K+T2qeZfdBE1mDLZm8udnCfWN17Fl/IJhcDXiyZp+
LwvodJdcGEHQYI3g5zRtPi8ytyDwOinRGGoLgUCc1eAcQ8RgSxtBPY1T+txhxtc2
vYbF1YZosyWcGSgJXPvQTE4fmkIf6eMpAlcaSo9HdcBtD6kJ+yFgNpPIZK61Vms8
/6qmpv6nEhEeEcHgkdpAqZl5FMtXFsShz6xsAkNDOhDuctvyHINwdKqnMO4bZiPA
HR2TbpnDzff6vHmnfMIthKnqmgZi04g9ZwEk/JdMh3J0tRRzR/vxeZOCR1dbTOsW
mkWCy3CyUFac32T+7uGnwVfhgoAi2+NAySs2RccUszw6xd3Tm3GNXmOehMc0dz/b
5utojAjAH9YzMCCWtP8FnucZfX5yhhG+KAOs/AAxrldjjZfdzYvbgyXcMe1W3iNg
UYsg0wFOjuLDTOzcVvbcr1V2BNhLxSYVUEDnn3PT8+U7oYoykUlx8SUlQyJnKvYa
I/QRCDNbtW6fVzUcTRp0+XzUCwwjAoohMTjalf/+4IMdqu2L7h1fRhMvc5TmAFx+
lyHLjRDV/Jd+/ZWN6RcnK4yuSMaWTNyP9W8iEX93Yx4ctHfOu4Oo0hh0xE1zEglF
HIYLV1S/9w3Lqx/+hEMUOGnjumjDnztql1w2VVXMQcSmS4C/SRSdXs2mdwVhaa5b
SIHKvzS+f8avZydDjj2wyrIv/rxWk4YZpF6aREGeNbn4cjWXYQkqcn4MMydlm89C
beTurMr8gyCAftK/df8jJxVpwAeML6OVBbObsPIvHulvoKj2ek21RXi2OqBGLZju
SqskSAgw5ZWD7mNXk207AbVSbhKGaZLBB+qBYikdTG26QEuSBu2Z5Pl2tw0da0dL
SpgjfBQSNslra7XWtnicNFfiY78ktY32mqHg85pML6XtW0s5R0YJ/wm0K4IjsPzY
nZB2dfAS9JTJzwd7UMcOIA8cRTloLzeL/6v63s1uqS84r1lw1TNMrtYzN3IWmmta
j7Ez58FgJQfbaMZ2wzJwutwh5aUr0M7TYRnjrTDXnAel6ptVQFJ32x+qDjG5Kirh
ijqyFkya9cXkJT43t/hOQw47SbCAk6pdrMdfCiLVvy3dRioc0qqKz5OFXRfoWsgg
sHvdqECGXSkKcBWjCsiVT3nUirZkZOaLL+0mVCmX6GC+JfG7bVOoTLJu2Uee3KIj
773aPBTQmuNRSzU780gkEww/C6BuQxO0CIOEM0h5VIYZyDfZFBlbXPe4JTYcpG9R
L2sl2gdC9hAQqaGSzH196LWJFKMSQbsy9sVmIC+av1PZihYyTEVXDJimDbDd/8GH
GKI4gGniYziBSsyBTYyTou07zTHABR10fsujt9WMNSB9DyVYnoDVJwD8BpzwguFa
J0pyB8JOZYd00GRhyscAqfjp81f61V8FHYJ6/8fIkpChXrNep1OUSmvRbGDJEfsa
Y+ty+rm0f/k7MKeyw7lNpX/5WQ3xrA0Ps3JYHnO3Nr1x9hp95+lpAvhvFtJDNDpG
vX9dEzOhzCYu86tz7J8H3j1AuR5CMrUQJW2TgCVG7v9t2dGBtm4VmCg3Tgfowgum
0Lk3AE6ZJkln4zksgdhiQgQ4f9z8rISIVufY43LrpN4jV7BA2GgxQTIFlfYXAq2n
k5JWF+7BFMPw5O4fKUCvadJbRuw0V0nu+zqU257iP9m1ZRLrG3Rq6tpS0fa+ti5D
kMMysMXB/UutBh4t02E5odzuFWYirReVIpRpSjpfKfTKD6NgBVw7l5XylOWoGMxH
K6cqVLiSciHBd2gtaTL2fzihf53oo+4XYYXCON8BbzyB1Z9//UPzMqI4/y8CvS4d
VmPS+9qEEHLfnxIUix/18xGLrRBYEB/d2x4jeNZeCRrf/pByPxHLO16xCII7Q53M
/vmCq5hCQY/8JOEFwg84pxll0fwnqRRxh5SSTDnyEzhCu4y++atuWECAKIrTfxlU
3NAqUkfDG2aoVFE8UdQqUnP42oZVg880A1ITqKkhNwRZcFnepuENePkagNQXWfi/
twCPj4a2ibtRpe0BmWWajch+CuRRRbPVJl+v+Pav2CgtssBOMOqlbpJwrZh18LNF
vVraAx1+86mXLBq62QehRuDLEl7CnFcfWsahPuweUImKR5JLT/J3SwfP/QGV9blb
+8wDOLqW4HDx/hiwqS7ZLRZODDT7SbAUhNAM8EcspBYz9ZT52OZyTL+1aX7dB4ir
hq2E2TRixnaKzbYucLU5p6GU+nFI+FFS/WmxXe0NUCFCKld969U8+48JI25FEnH3
Gn634fGAPY543zMkvPWxPpWt+zc28erBpsgzeIXVAytxeyP1Q/97Lzfczvl3DmEQ
KA69wrqgHtVIdIElXjvhAaoafkAeI4jMp+3WrqRpw5BgrIIkZUQHts6HD2pzhpIE
cHvnaBrTYcP+whWsFyugmfcslu7ipH+yRrZKyg7wiKf1qX+8UX9xHQj/h5DP5YI/
vMvlnrEb3pELkyk0nWIiLekbmFa0B3/kY9rM6NsYK1Cgs1da3zJxA4salk0bX2m/
sO0TdXon9PZI/xLptw4R3g0n7A9pDsB9Ma+PxYw0DaWsn0dYowOZnUTaUi4WneuB
lkyLwZroVDVKYFPsx+5ui9Jq3tQ668QYllno1rlbp1MYh7Kjo5/Ww+3XoxyZuqWX
lCdMhPSbzAPZKJuKp0KgUQvN6TnKg3nsmP/RR72xY1OWkU8wO/iqYR1Oz7c11X+a
YQZhKM40IExTAY5GlvzjWsiLfXg0IqZm47V9ErhVsweI/Q/EX9Qr0Sb2YX1ysl9B
MUhJrOLc1oEyINwoZRwXTnM2RMIyo6xMx9x+9MgTviKRnsSm+UyOWWP5QxwCdncR
hm0dcwfoi0KiyBykKwc4z9H7ZZebDvc4b3ofiNdozcjBM4kWUVb27TKMkag+cYDA
1qzSrvP8P1GfluJBD6TgDk4IBfHjJIZkhzUBCym8TwhM27Hw9ht8Unoj9PW+dru9
g8MdsXHkiR0r3uAie7Q7A8XmO8yWe2HjrMHFyx/BwS3bgl9NG5yjoBtDI40ATWk4
nrq8AXJpv6GFQEDO0pDyVrD5pY1kNeAbI0rLnatmitCAJQ7sKBIBdkgIR4U3K2pr
4UO+MwvOn7Qs25oAowE+mx0cjxl6w560lptxHLUZMvCt2pcB0vSmu1I+TnxLU9FT
T4ymXQ2VUl//lORdAONxghqoLxdOAYCjVWmlp3SWXAKmhhdSSe3b9QzV7mQ5pNL/
DhDp/efcFk4F7BZUUiTPRk75VCgX+UudH/thW5LvEL1lq2F74G0TatyvUQUAcFe5
F+e3bUBvf6T+PzdYhiUWEaKQ2P8GX8kVFoo6qCZ11IWt4IKswyUJPgcNNZ3MYyyd
guWBYoBnBZ3gwUf3Jb9f5vQypdaf5JIkKcNoDWcrf3bi+6Y0jjR83AtUv+za+ypY
qvLtfL53u7XeVe4Gd+dQgcpbnxc6rEz3u8s7DgMP3sI4GZDqWbBHW96e+GVPrzZN
F/N+mwzAiFcY854J7x5ije7wuxC5CW6bWq6/t0+R7dM5PMZXXapzB/Z2SVV2Q1oH
LMxNXoyFzs32Wh4Wm+0T1UfTWq7DPPKpNQd2xlYKck+q/yhuogCr1+97m3kDNbxq
Zrg2rWcq/PCNdpMWdT5XxmSNu4wx6pHF1yGqKbXiQVN9UeVpeicVbYFVJ2ys/Nnk
ByP93o4a0HPVCFTFx3ymYtcczRf/HcAtgn4PJ6gbkICaYBC1OG78UHgCIe91iAKd
eHLkOURv/CAKiAc3RIC1TLJAq7h96DNybBxN+3QnijRUk16uuaqWlhMGySwZ9BG+
X3HNXw7z2L1MbZeo8xMTmknsLBhw0oqhUE99ywdpmptEXj4BNOSf29sSpwK1hlWj
qPD4qKwFGsY7RdQuLv+ux5dzPBeVKeFygmrj+/PDveFY9omgDN/1Tr5BGbvfvcEG
4+/lfgHzeIO/ufpB+H9Ca6X6sIcxSi9PNNCtp6ofwIkj5a/fUkacNhT4EZeyKcH6
5X4NO9Gj0wt973RE4ck8DqPk0JcSlwV9TJT/AAB1PbrVeqJePic5x8eelWTwQL+O
ivpBF95kIbZG61V5tjP1YfJAcmF3a7IsI3v9ucBpl8BfuR4c0be1VbVcFUQVemWY
OEnC608KWXbP9p4jWw7jrokmg3Wh5KWAfJgtAbDKu7UtQbotMmmvggee/xaGP7r4
BV6tCEHUXVl7y1jNMq/cXzGP5lhy9DgkKqyM/SzbJ9zR6kHRpVs20uBlKbEq0O7H
O5TlvmrBchTwIM7BjWiDHcgqS7FIH5vQyVQdbAQPZaj5DCci8vIFDaD/9jMlKaTX
9L4OMhZWYFbwTho72KNotUJ8eZRwVHooDcKd47YrkCiTF3O0s/Rh4qbv0KbwTCGr
egoDGXiANUJ6m/vG9I7GJUerBEUPvtH5Ch0cY3yVrSmfcJeVvDGPIgUiCBr9Gtp5
Xg3QaoS5cY7HMG/p16TlaG6QVWCKOo4DHZQN9sGR8LzvxF0ZTsTzUEw7zayaMUDE
FCpAMNq/BNJ8jtDstq8IaSJ0GVkhsRG0auUoTN6YH2n0hKtkRJG1+25C5BfTJt1n
ua3y72wgPdmE4GbOxLOl/96QdGcZDpbrZmkVi8tIqQW3B/vQM8BHXiz+EXClXzNB
RErJKHGJW+8UZ+967i+B1fKmZ+VEN8aGeo4jE8ek4c58Wkfi246ZPCSD6/Qx4V+M
lbCpT8EFwM5iUdLrxTLn5LuO+7JxKLwFqluJ/ITAlCVewxD+QRKLe9u9ejIq+Xup
/Y9wl6SHb37UITm60lmLkc+8LQypIzQUF5uyDO8pWrvs2R7JL4J7rM9/RbecPWvQ
vVfCNHeGZNBRZTPyrqw6YVgWyDppV0bbvYSCU+7IoPAWOxVdHffwch/nVjbMTktr
dZP94v8QrRsn9pumcFQH/tCjzOpr+oytZS6dvQua5ZUZUHiomjRHKnRG+pcpJ0aI
XtBz9W8B+6uZRmedUtqiXG4Qq+dh4uQ1L52BJSaQcGnZpmFN84ZANv0rJzuEOhT9
UtQYJJNettUwTnncwtEjJSkLxyZwoPRJBrXPr8/QXp8zID5ZwafC7i/V/RfUX/CI
bNcR6eljwZELByquIUYn5WrnZoMP8gaY/yu6WOrd70ArPrlyLVZscZTgxYxkT55A
PhPsq+58uwzxv7KE/VEk+clOrzraSSiqrpPR0maATyBvyEPTEmTYqEhwUREOKBdu
wIjdp7QXTJ2Xi3zLVx4n5pircxcfRIz6ASMhPrfO2OB+ENiD2KJgiQrju7jaE0/k
MgluScxt4KxoukUp27BWiLWDOHRGfP3e2nCrRVIQL4oQOAApby2Ch2mcTCIrbGpL
Ghcft6jHSOFjHd36xactNytDXHL9PyX6F3LOCnMTihNL+6vsSbEYMpi5pStYO5uD
sUd+KZ9jBq5kG7d1i6OfMFi4ipjTYJ4dT5ZBFu0WDu76wz4mer24SJZWNmnuAIhf
e5TL/MLNrmTL4jxmdb8sAAowvHPZXm+HuDTk+UapDyLsQLY51iIfTRLPafJsNkUt
CSnauSnsQ+1b2bTzAUX0KRZb3YcoZDhML8+O9/YHbMxgNTlOaLwUfVladB3Tzi89
9T1AWv9pMLsZkZGx8k0D/sS1qz2yzms8d0X9rX8APCOSDQaBbiFOwWJT3iShANTU
KdxVtBbmiyXk4K7o0lL2TRHcaB+RG5OtrGax0Wogtpeb9HrevL5gcUUC3UYPDtVM
UyYT7GK+iJTz7M3Sz8X4JPSA0I6XeeJPRhiFESa5GeRHFxg/bDaKugJAsM9eLMw/
/+aGHR5gogwqttQoJYe35YE+hSaxHMDzzSnHLR5ky2UzuD71Wui4Dog80If8nJw0
fnSrA+W+d941fz5mXqex/PNQXOqclBWw7XZ5SVtgyJk0P1VOCu7BD+1QuOgwbi5F
D9kDVry0QsYOB9A9mr92SLDB5CV2yd8+gxj1h8ED8U5FfZgpYpgkqvhGNzQODWwm
qw+jbGSEVH83i/1CRnAGF3mAKHr9ALr5xIpZmUmtIDnhVHe/vac60umr25FXfL4z
KfgBRubbyVg9NobDPMZyvCXQXDvFjrtyNx8MxE20P+iYzTUoLOQ0PKwr7gZT8sya
zgw3LfeN05GeDcFXcP1P9bVwM6h2FHpYVSLkIfnRsRzyiwwyQUbCFstux2iCvnrQ
G+PqPMHfhgfe3sElAlE5cUIrAtR+4bnL5kvMLRrHplV0uA4d9nqefXrZiGDfgow4
uSzo9+GUqtMOQW68UdLFWCmsGF6F4Q/CQffN17Jw2na79jijHslFC4aohBK4C9Un
lvDshrqfGFnvOQEpiB7ZDvxqLH3Hctxz13l1fu5+zO5vUnsmSZi8Xs4J9bfeET6Z
8PZF81xWGcAhaQ0pUzVubsGKduBwQ/RekZJoTKdrSVXGwN3ZLXH/fUvkDrv6619X
455VUOk5L4LdV9/2MaXGMtEoFK/wySleoKeOCGWHohefEZB/OTKDrYjkp2LXr8VI
QQbOJe0obnu5Wfu7d+RrUrL3Mc9X1c7t+Ti/nzxlCGVTatRO8bMeXZncmQ5DvM8D
URHvZYqpM2JcQm4NHI7ijFzJtWDu/Ua/K9c44y3A3RNDbTrbGLKqdDea74q+Sgsg
TcerfUNe8x0pO634b3fXirU+K6dz2gicNkkO229O9wYT3AJRUs8i41S4QUJsl5er
xs+cm7osi7vSVsZ6KJUEb181GovnCVlu0IYRVzN40vQJsHcF+DQXavo7p8E7PX1d
voC4TLgeyu/35WAxabJG9nW68aBUirl7ytr4sC7FCLSxus8lZDwr7xfpvX5KV95M
WtO73/xxNcU/2Lt+IUmLp7o5suh2uOYK/w9wdok5STmOZHqPsDeJp7Xl2Ag9bIYk
EfBrYvuMPh26rvgbgnhHhJWSFDV7/Fmr4yKZnr5IopPpSTqwdWogDoK9yH/FaHXq
oOYAga4tt/5p5N3AAGenkuqvQb/jNiW2fz5GgPBopxypMX3jamVTBg2gtav4IhoE
1WZgx7DgHnCQkrLeURcwbuh9r6TZUqoryWF3R3MjL9toGuduh1QYEXQtUBCj1rIL
JGjyJpbme8Kzx9Db2o4ZlelN1x/YGPy67a7YVsUCyZgAuOtXjlE73cdntm7lZEiZ
Dz+btfAOadUeJIWToUjuzpd8+lPSwg9tTmcFkgtCQCDmUPt73b0qH8gV5i9xk+Qu
WvRuCT4dGY3JvbXN1goHKUgMKVFtt6EhDJKqTxrohcRr8l9k0bj6MAIGVy03xuLK
NxQ5rh+JM5OpkuOZWMa3ls9IcmskRU70oZH6pIHNRMJxPii8nLvpAYlNyiCKDjnQ
A1Rppk6h9wrn5R/+9sMQw5D7tn8GV9WjvZ8wzAStPh3yGf4cF7A02hAdr4krt8e4
cZKqm9hoZreWCmOQwuoasFzRKEZxuCXZ+OLpj3G1AVXi9FOncYnNmsicQmzE9ny0
8xVsT0vugL7rTZofCc3DqcZyKNnG5MhW2hW7EQt7zc/kQHUFCIptdt0ilwrq9dbP
uEkLTt+lj9Y9lvP7t4DXKlmHpLEF7WUBuPlNpndFlILJaqhhgFfE9RIG2Yfumbl9
dd4fvDHPrOG4bUolKZ6eM23Bm9EWNyD0ftwk7GLmkGnkZF0EW5c5SLG24JOWRunw
xaXTT4WwKOTajBPh3DGb9fzNDl61lKT8ZshacCCOS3iFjba0BDFL4NLo0AgGeh8U
X8cIv1z7omAUaDXSD3Lydc82i5TpC2a3lXDSddsV8Jt5wsT2++I99iXRagkgBU0+
iTw7QDa2k1W3hEw8AUexRlB3R1NqJO3ekF3YnZy6rCRNizT5pMTYPLToIbwLoeSE
29oeSChDce0f63BkeyEcHbwN6yi4QZ85N26iBCUFOi4Y5grIwkoV3AFUVtujDdnn
/2CmOMyIwFU/fkd7Q/3SwPvSwQRKd9ZO0BS8utU9Lnsqx4lA5FXDE3M9uBRzzF+m
kdeZtE5OKmsOX3iF2zgmNi1rzsmaK5+eAKldT0v87p+GtGYSsXnLYqcl7EkDAkF3
wLlxwFQ+eXQu/wzt1zupKTbsuSyyHcS1K5Qp6t933rWRLuTxu11QUAj8FiZYS2vT
DWLxddKjgLZabyp7mS2XqkvVK1Huh4xekCflmGlhJFgyMeJg5HF9nsWcVwQ9tlne
cVPE3cIBQf1l6VYBC0NGzecJNucXC+T+uU1HSSKHFZwiR5u5SAY1hUPIFj65eWDh
tNekrq3YmhKTNJSKrpaaaksef9XCvadqshJMjS7gjVbcP38JZcnq3K1AKzKCkxBB
xF+rq0BESSV+5BbWj6NJETU+HZfEYT+SKJsC8IiDbeJaPMVnA0r8vQdwsbAznFlM
P0t51xZ+TNym/Nok35V05Ab2Z6pVn5iNIZb+Eo4gRWmmy0ri6VUKvAN9LsITSPgx
Vy+q5eGuljz1C/spwpnOrgHl8XjeUzbSXDng6irQ14FourWVFaQBvqD2Wq3OcuXI
ArsxpDJ/2+QVskx6S3FFd9A7t0e5b0Dxlfy33MwXrcKIksIIvlPYyMO6+lSD/bJc
J6DNAlaGfuXJscqRbheLsDuNOeu2eEkCDvyf8v7iXofyPz+DMT0JeJCyW6BF5KEI
L6/JTkVa4IAm9BMx4pzdRSlmjWe9wC1dpE6c1Cvvi2g+lQJHvxWpkev51NuDAx7D
xttBhRQV8pg2xaQjSiA4Nfmo5TGRdEaQrdHz8wg2aCZ52TQSFLJJsdsnOFLKANF8
BcpGsgZrylHXTSPrClUomBBQqKs/ilJ2kqhfwMDG+5/Jvl4KADDAQnQW8lbqAXLH
Ag5XZJmyKPGxpVRv/hPMY6uDSSiku6z0NwNXmlQUWXNrqmOX3nFvqfWe5PzJSsfr
3XPnAp5UNTm4o05HoaaxH00at2ZvFEjL29sBJy11BhZt7xA68Qq0HZfdrBgjgMYZ
zLdsydcnV11MevH43KUL4zbLV5sU5CsgZNboeLUNM8YPddBYJkwWoQpdchKIDAkb
eICWKZ/23OPBENLOhnFrmCaEAF/rsR9nIOmVMIOg6yEyEs9e+R1UKi/GXyE3OcbR
eqaOpSlMC6Ix3GdI7RCrLtkSKW/rE2qcRw0XBd4RQ2Mkk/2RnllrwKMnSzriG+9U
1EEG4fwAkjhdQ44hq+evadWDXUMfC8nXuFxlaKOCjMwRwl/cjqEE8anDSKiDdr8X
p2RWXynQa1mZZsevABBmkXQX20/Nd2DLkOnGuY76L9BCzcP6QiPwCL86L2e13j0I
q9wBz+o8nkETEYSUb8eZ2Y/wkR+uuL8M48xL4/4Zs6v53CDDjMRnBXelrge9CRv8
v1UP3S3bZJW2mTCZAXtdKza6mYtPzVQ4nEbhB4u1rnZBsSYvP12TQsC+kWbLvG8Z
5gTIjoddqB+M+kK8qNhYvsRlIuXaENU1imNGPwmWbGyqgZuoIxULsy8PWQNsZpZZ
cH3bvbCHkH2YHMfzveOjmwq0bJBtlVjcTQ5WtnkE+UWFDQPj/CjM0qNoeMMUeTLj
tX8sIhOXOwm0M6sernu30aCVZZuRkRAiT2IJhSfWZbwhqd1OqFlk8UwwCmNB0Qro
nPJ4By6EhTLfYTqMtdysYpJKY8FnRTsKtUdbpZdEMWLv3l/TSi6JZD0xrQmmaUcB
rfrJg6QSUXzbXcXbOr1lD+A1VjptiDfSdF2JjrxHQDCAG4Nkrb2D0nCJQl395bbT
xljSm0LmCRuBXZxirPQXukSatDXgtWUf2T1lVcp9/y+jgxu4ocVsaSQwiO/M45FD
kQfZevif/Ln9tv8Ozmv3B5RpX3mE5IEfeOBGFW+pNfmANkMlpXJkGLRgxaozwpGC
nJU3Ay8/RdR1O3W5BPhHhDeuy4IlhtTgmJWnp2z/v6bZLM0uaLzTvH/LGrj4JCqk
zR+xchS1crm0aT53NHpEXhFJ+hGbTuB/8kGBLB4tM11vueAnbPjkvNcykOyLEGYN
xsz1GAmR6O5O99EeEfbt9dyfN/GbIiFDazbezM0HldgdNbVccEbaFzxQEKi5ZLhL
29oldwQWGH7UkIC5LJhT+vXwkedtIPrYP3Tt4CB0yiuqpd7+uXXuXlwm6+nHr6VT
+SJe6JJ3ueRDIvV/c07IUnQNA6EjhUtYk6wd92P7YsSiBHHbHTX5xfPOVGIwOCVk
8f8/TvIvPhsD6Jzzs+WRHzFTkKOtGjxx/BhF5sO4tElKMSuzDXIk7po4yn6V0mTR
5U+kHcAtqkfPLbGh6pSLOWm7gQwMlNLNgDsmvW0B1LUFpbh0aY3UPS7jPTxk5dIf
i/Z8hITFDhb/Wqtb+wl1qxnDSh200pDB/UUAeP29vQtUpNWC6s8h3b3Rioap4itN
V4LLz3JPNtNOIrRZmC3KTX/QHLJQNDeqMjbul3CtDdlAUh0lu5anpawIepQpjz2Z
Mz4o7Dl1AgTlzFCyX/sqq0ERLtsXcnTnYGzur4Bpt6mKujz4gKntT1UMp6uYBbc+
9TF8F03ZG90EES7LOxaVZDT1HNQkRTlfCDL1Ac7hXdrazJTpjKFEHvc8GkC8jH70
Euavx0bfHTopaAXFculp/OcWFA+VpqyUJOg+ZxTEqH8Q5GXYx+euHGsULBKqEqMr
2uhiz7xILOBXZ39+v7S5RvLOs43cdIFbT14pUrz2+Cd+T2qBJ9I2u/d5cgxcJ7UB
I6HUFc24GHzLw5PQCeOUSiAiDWo6lAJYQaLTBzktV8FQmzRdQuuXAkiNHaUtCtGn
vq8hb8+92OEDXn43VVtbYKIA2uJyKIyM3PT0l4er9B4+0iWBx0MG0867f1SivgAv
9w99qwDWz3CKrs339jQvrj58cAWEP46+arvRx6ND9tnUxLl8G6pvigLYOx/zLv5L
fCdusaI/FdM5JlzqHAEFqpi06fqEIsAIB0R/+/1K/L9nMbYWPHuHtWrW38BI+1VW
B3QbbU32h4xJB62U1Ef3Mc+DaGC9CUWZfyLHXD3xF+WbSzcOhzjO9Aye9o0pxHAU
NNkXUUIPYSDM/ncAxGkow8FLi1vuCDev9FsUjBKNVbXejKm3QEQC740UmDicRVCV
u6oMsD1SecMhfX6mPmWO8+sPSbE3Pl1bdYNvanoDWnOlBLrRzceFkMxyf+4LSua3
yxrWzvWkV0CRqqi4jjLb1FybHVRl7n4a7h4PREVFpTh+Wgyd23cppCSNmtgccJmc
XoXXjaAbQbQ1ELVr/aMuLP4beMnMd61gXQvYP5wnKYi/EV+HiAHNY0vih8QeK6E7
zL7CZEyu0hV0mm+/geY18veQpeYvcWXiwSLqa0RnWNqN9ftgVflX85FTnHY2UIpC
Hw8eak26vDSBkonQxxYV/tsmskp4aU+bUdT4BIltUsTB/NervchZsgY1J4vQz3zo
vLVuRa3gT54YFIyIIpZ1aZohM/5Wi271SnzK53ZqcZCYozx4NoXj4nOSrvesJhuT
2jbN1HBi/Vb2x8bV6DUON568vavSC2Hj1W0dtRDg3gnFA2dmr3iPnF1vCsFSF8xm
LydIuhAwA3jjjKPch7FvmOyPp37W8OIi/ybSHct/VF9vWBKINWewd2CtP9t1pAeU
rFbFKHaQE8Y8foPiyVDTTw5dtNRSNyw7JTeQlwGoD7pD+ne9qYcKannD7n5vrP/v
P8nkMYEAu6+zIWeLPhaD6bohTWFdLa5TJesRcVXPiZpsEZXhIV344WuWGeGcVgs/
zU+YZkiN5F5rqHzqXDh7IMIEGpGhLVTQ2KI/TQCPWU5y7SSMErCyPS8pa/AAFBQZ
1NUg3GXqzWiUdsmBax6r3UIxUa5zCxoTYqwiWVu79sMape/6WsOh+x1pWYvQFjlM
3gdEY3zE4kEPoI0fCHZYwLxa5AuB+Shits7qUuubGrm+11v2Jdghd0DeFAT4CRv2
1+i3Ns9RLsiL1ZiR0fmHghRJ1zjCsb8GXJswMSmgfKiA89MOn2Gi/XsjQACkJAMO
yHR2hvZpANyeCNy9UZHZWJnZmJ+xIHX40+z5cShBGNncaYcvHO42PB5uQ7PKg81F
po9WDvANb93oIr8qmUbVTBWxpYpMhos9AsUgNnnUh0fHFJ/mnuhJSF3iZkJ5Kfxp
+5gQkFzN0tg36rB9Qh33sq03N/za0+rTSFXUQmRt5tMsaeEy1oy94nDh4oplb8nQ
w8T49kFXkEOZpXjDI+vLAf9DUQYFI2/VXaeuveoEyzSV8Oe/THVDUlveKtjmx9Jl
zXrlnQhOBzXeR9SqIKuYOWpT/sPufO73ciMMIYqvDVvi4dUze+13zupt3BkvO1IT
3VEfBKM1sOcqsJML4/bpPbiKHZ+7R2+JoIow6Y2VbHeoanKMaV9yOszKLKIRg6aJ
KxdQT9esl0XUZ+JtWnL1IFX/W927WBGGO/AfmgKnlChaRrauAgWd0aHX+PCFvvId
3uAQi87D02GPvrjls6If3eOOZqEoUKaoOxDExTfOPJTeIb8zgWAj5aYLqtM++ekH
fQK9j/9/2yI+2GQpkIzTaBbDkjThzyywuk+efSReGyR74l/Mdq9U7cndi+g0tmdn
0++IRZA6J52K52z1qR3aUEZAT9R1uJB5muiTzENlSS1zv0byXffTmgdVthxwqH4P
AHFsIh1ZabRP7+1NyJ5D+BvHn45E8eq8ki0OTm5d20zZdLAO3NnSH1DIVLreI+6e
O+RslMPDpyFxjfB+hNuTYJdboePmo9dyuQP5h1Uy1ZzpuKUKKA4FsE9YK49XENOW
ffsmTKBLC1BTpX9dSfa9DNJCG7YYQCI8rWnAGjEkps8YUouCR1J75zIyifIBkcFP
yq64L6fQYpdHMiDdRoLbWjtrQeYBU5f5Ih9w8kiWCvc/IXNxIoheqniKbwM6xCK+
Rmq6V/W67FywSv3/ie2rct+zAbtGK2keJzlE/wCcQaCG0DxnNIjTyYiilNeGdbnX
ppttnkCACyFSV4sH4jeeE55zL+SFk3erUagwX1RM1bAXWaIYIWWtggHJLkQ1UNk2
zfL1qBZq7u+1VRcH2yrSmKaFbCd/+TDibNSDSpoTceb2VpeJy7hIvtRfntgQVCM1
OaVZ9CV74bPFC5fAF9UWLglE9iElDoDycs+LR+I+hxaqtqu8y68XDZ4hFeDu3x9x
v4reDT+8u6c3wQIhuR5hx4FWa7JexMt0gKEzJ+DHHfa/Cp/6CTkFi1OXDDgjQ+Td
pkunAlTN7k3vanC/cTNYVPdQWTiXM+lhjs8RorSl4KQVY2htP27OgaooxJD4m4xl
4Ggh7f5rgEeHCWsnaSHUHikdnG1VvE6fnPMoAr0GMMVnrF0PhzIIuNJIQAKZLuez
ZQPWgSHgYheNVQu+vgNl+2lHZxcI90HqJgzdrJahdn9LUQf2ZEywQbWM/izDIJbw
VP9FzPgsniQDk8JdqGMP0ThZDFB637RmB4L2X9YdVDbvPFQyOvkjbV+PbfZth97R
Fjvkt1VNv0goYzjRcIxR/ImwJtL2Yuzv0O46HduYBzXGCbMppXFl7R+lJoJEECZY
Df+myoxDi4PNmJJUe6j1OuG8C/XFXBi3dfTfRk66jFfT2tG0oQeU0AWB90OSFz4Q
M2DED7nqBfGrhCw1qooEbaHsbMYoQG1VnkFSxfB6EtnUudo6ksx0U8wiBO+MROgt
RrZXHaimuZaKPbK5AUNjrx0rx5HA2lVp7QnX8NN3+LxmUIdVNH+Dp1UdJwRaAfs/
EyDZW62w/nbU55Su645OX+rkNWdV3j3rp08Id6e7q9gtWjxGpNPTQOcM5Uxj/D+1
fVx5Oh9YUeWptDQ6CysnFFTOvG9CAdk56xZapYWD8GU5R/ZsTN4EaAWekovY8/f2
xCcdit4w8LDEkS3kmjSwGCNP+naDEMRtchzm/0pNGVMTBEAAmKxlmiPONVwXuuX3
UerMaVIIpf2+ay1Y+A92VhGEYXvoug3n7LqzRtK8wrZrIDoGFjoIv7yx0EvSZWYT
y5yJ6x/WHdvJCHe6XyXcreI1ugLQogzAkWwubEusx8LLMvA6XPMdNd+OjXVFUHiu
uWO+qISJI/I/8tYA3PbNVObbzBao1ADIgx9HgCFHxFsT7wMMMO80kMqwX/Kq4GmG
EGCh62ME+/RnxPAedZGuKPOH6pRNsGmngfOan6n7o+m2Y71WChCAUqn0Dd3AjDIO
ciQCjdi8YoYxn8o64lpapLBwpIb2+op1j4a6ggzUl8rLOOWbm7KXLXuP4PhKUzHb
ciKS9DsmnIhIjuy3iJTHU00Xg6bJuf2JuGx40VH01MGSnsMQ/f2w93WUp+Ll5jw2
UdRAD+mSCmTiPGxEDX4rjRNEugVXvQ+BCbUEtlfBHSAH4H0aoby76xf3sDDbyGwY
WgaPYHRbtWfNFA1sg3xlLl57i39JOyVVOOVAa3kla3A9fGKO87xJwp8jKetKLIQe
Fn7dgvIJ/6RxhphCZanFksWXjMQstGQzJK0giW8KdqJkgjTFQZOa63nLHaFrKFAN
JoiR26F1cpaak7qKFrvvDr7WLudZ80y7rra6Q5YGHdRX7mo1qX2xpcz6uWVzz2BJ
w7pyr4nzXx/n+1WCBgKP3XJUoSzSk5bfJhwrvbEUNQdK6+GDaGq9QoYnw/Sh6FhV
AMZLOZ1+gSALhO4xn3aFQ0xVmhXnEBtDsNMposBi1EhsUN1F8XqR1LCpo57rW1Bg
aWF/WtdlhDpTQWFP4GTzqlis/tTTH/oX4x5kCybsyyKr6CDis/cM1CpUVrxBNAlQ
R5MvUCmnQ0Avz8jDP8/EBehzTI5aWQ4ZWrMY7W58Oru40H85ITPy3n7W1El90w6K
v4vADxlNDNw4y1nuCXfozkdESWTxfkC17MXGcF0n4T9ExIfCRQlacSkhsaCzBZk8
gjVQY5ZDVcvm7RW4mf2ZuWPd61S2OelBtAy5sB3BnNwtXkeOUkB7vsNFPEQsP7xt
HtOGmJONoQis6lYvtup24SBfHDpc2mqUDMgyzefXtZID2Y5ey1MqSsMBLJLK4bcr
KZBjPwzVkVqTz8RmZIoYcB3Y1jFW4k2n6vIW5aoSvwi2tQzrOd2dhcN8/JB53QEy
/BPfFw52f0HOL2qxOs4kTA8BP9ZMTluLQnlKslElTimRdzK4cs9mVnA/1RvU1WxZ
3CM8e9uK9J3RPm1btbuME+FkxFw31WVEJNC9Rl2EmfhuZ3KjINoOFBlVIDuN1Bh0
+bnYah/bCKJbtq5xMke0L0Mb5nORaHP/WdEWEaNUVCsgiJLTLczV6HkWTXEbo0ej
bjjiZ26hIj477Ili7cfcxYQeUK0MgQO7aUWu7B5PGXR6ZiGWxpbb5hE5EwBtdRxh
Fa+I10cEpp8B9va2Ko+VZ6mDmDzUBknNGkxjbm+p+tZ6pPBVC5vmWBfvCprfJPtr
kFEvWN9mWe0j+ZGzG3LvlOwo/qGOD6Bl5ydowQZ0OCuAfr8gC68s2e5pUEhFwQPy
sod6N3e/NFVERmyPLC5pk86VEPBVOlb9AFO8K8xkYYu4OqnfgSNkdWqxTY6UYHca
+5Om4dUeFH4UakrgMdA8tEo4kBR+8IU0GT6PQC3Ax4/x6YM3PLsYaBhRS0bBlZ1Z
nD5tUp/BK+QgBGhKMOKYts3gznXZTJQ7ILTPIItn58G9EfiVLvlbgUxmF0FSmPHf
/ULpjjWBoaFWx30mwGZcudA6EcigSLHz57VD3PSdEh7YxSg/8nXQ6NVuxPU+z/m5
9Alt8bEe/A+FUGiAfMhoZSJb0qcDxjQ9ntjQ6GGP++S3jMd5+I/JwR++G7cDBi+n
R/5vRFna+DVbQQpTz9jkHMRKhb4lGTZ533pck4sRtV62Khz/Mm7bnFiw+F3uoEbc
7tHkgmUiXYmcnQ8HCnygA0ThgvVqapioLWrpHi3kU7FrTpfh4H0SLLZt+B9cRo3M
Slep/j0QSfH07/hpzFexm3c85RJ/QA3/TfLIKwH7hBY3aAHbKdXgfBf2qtrjtByu
PZBcE5YB+7Xe70evRB3MxLl6vtRQAL3eV//YhqXzGfn8KqlwfTpMPqjOlgo2WO9s
vS4nOzK0RVnVU7Lc6l6ul4rBWPNKO/V7cjFp/Jhtd1wENKJtcOkuLnyrEyoZsxaI
8jprMw3Z5WSfyq0Fpk2wr7zZvDYVycpskTSoA5VpCnmyGtrJJNEsdR6OFD13cVR/
VIuh6iB6nuOmGzw3PmSJGTo2sRpyL6uZNiSAfqHLsBiO2aS9v7Cn1r5IlXf7jrew
QeF7ucfa39fpsYBk4kFDJvnBp6BXCzDgioZuR6unzgWn8aZtCtOQvtnPE5xWrLm8
z30dhewwTiBQHxByhP4NhXovxxp5PPW5pvKW9lypvuU26kY7Cljp7xf/ABrTR6V3
VYGB7u5Se3dTzjhfAdlJazpavGNPIxxTdpq13S+xtayfSvDtiGUsbaRCUl/rGh8p
ApgOo7+VmPuCM32NDomSgys8efgSHf7oB3Yhss6K1/Occnu4I8I5MbtaK3d1sXp7
uNyyttFSmlCEyZUvM444nACqm7w6344DeP7Akw1SymgjQ1Uq6i0Um1h0B7KLgFmW
6c8pgkMBLbFSZionl86xkUlYWPUCBmgb8iRnwt2fa0QJQe6Wcyrgf1INaeKFBqyH
dR66Rmr7xx6u21K2u/c7geZA5yVTUT2sAAUYDvKxsJn7Rq6ICgCrvLDzqU9Ny92A
k+Jz9jAV7bbYITPXHBsIgfu3EuaFzs8h9IjUOuN+JmVXDdNBHSE7MXFzHaHZJa1x
F4R5NQid/rHHyVp3UhVGoysjaGTN7cGRBcCP37iEG8R8DkH9jaexDoLWtqdsm1ji
tU2UsHzkxA+TH37o/nFUHQvqSZAnBucwnBksyhm4D4TMn/zs0CXfN3su2uYdYvFe
N+ZmaoBJHR6CLzfmXvxzvRx5O3rx1k3HI5aYWdYt/4ylk8YBNeQIhEbvsGoBEbLl
mJNIjAvIfQIQ7we37IwC1nFMGWazBGDjhlmFwv0umO9qF7GnuVjL5G8+GkdwgXdO
Me8keq44ypM+g0Jqu3FrHt99CESwowK/en3VRVUUvDM/WRwsX1CkdwGgBFD+8ZTL
m0w5t0Zenvwpr+LxlPko6RYk8E8pXY2Y1cNVHTILBRJ7xwdsOsi7UXHWmutp+0H1
KqETNDdqwrOxrXKvXqQgmSP+DJSHNniFrJfdjr/CmxmBlsjuMA1kqzXoTs2GCNd4
izwQkSDcMZxGQ2PLXe3seayqHTG1/xa1WGx6Gy4E6icbQJhxwjwm3BSYeqBBz5m7
JXHfaXs3LoyhmEuQmBh1+w6LSw6WrXncGsrjZ8k1TrfZFa4e4FQUYR19mWggS5q6
VWi8u0kMvegzrrOXaaUWx12DiEbCuGnjHf93OP+lBk1+i9MvWs7iej/uG9FlXL5s
3+Xy0lAYSg4d5UsiTFrWuavUXMFgk9qDKTWt3MvLogO35B0fWGtwzfneBgrTc/Nk
MRFFfWle9+onmLaFpQ8TWImLc8grlylOpJAYYFYNHlPnmFa2KiUcs427naybeQdX
2KPkT/qVab1x7r0gmoI7WXTlh61GAEOHrTdD5Aw4td5pJZTcBK0Iv88ftYBCWjrp
rVWuszXo6CnRdjz/dn71bMtvtdle0hoTIVpyTBG4/G7fLcwEwuOPfqYUcl3oXzNS
YVHdd2XKMuNmky89S/IS+It17ED4VT2JbQ+7GdtS5DBIjTtzsZUfA/OkhJnjepm0
IvsJJ2oTAJVMQBYn2u6mt5P1W1kHtyTRMbaMO3SH5KJC9sb9py0ZaAF5z2YPVGCl
ldkHZo+rFzHPUSsigERxZlzvWN98DfbZXJYV8rIxf/Ybe4aZI+oL3caixNz4yIus
UeQlcVdxeh5txI6vIEL5WePOKZtbULvpB8Ou+ZztBER+lTV8cDWJLW7wiWYomdPi
QHDlrCyhUzWZ35OVmMhu8i9j2XpD0rY7RWzm07pG7dFCbTEzEWqgpLctnfwKBm4w
2HrjABgnBy2c3m+8RH3u0r7YZd6fB2UKVjEgWlQ2V0tN8eA3rb/7j5w1UTjpYfQm
CGFYKkaYk93PWI4f39WaQ4OSsUxhAf5UK05babVvAuYPIeHoXvNo8z4WUg9MPjkD
XTzoioRJxM5G3Onme16qrr+8FJ1nmt1x32bzKDXWvt+u3tX7WKgk21r/cL1hb7fI
OXRo00FOtdAF8wBBnDMTpiShMvo814RsQtsuPKYfj2ROuTxI18UaFsokvRIJrpYK
MDkQZFN6/+jAPoKPdKgF30CcJxwOzbVLHs+S9/eWu/dRZ2+ks3V70AU6p3bIOvMU
aAvxj5bipsJIchW8SDgrP1H14b5V3YE7BKqE/13aQZm6xdMRHo2sLLfrlV+v6c4R
6Uh+M9Lpq2sIwJ+AWchEqzVNcgEteHoVJTppQ3grUg2Z/5vxc2n7ezIbCrVmZQpI
LNxeCRa37AO25bqeyzIBR4Qrov3GVApVvOZwUm5wy8icBWHQoI3vZ2+t2jutjjWh
PXmMNhjWn+k7wRRxZ42GrFIcb2X0dqHNL7+1JXtbQqlWCjuEfjcHUHfLJuCAhA+3
HY56r2I1uP2Pcm9gpEU0uz9eorK+QRaaScJcly0KaSK4UID6XajOCur5W/fEWlrC
EBUGXHOQLD5OARF81uRcHR7gS/akUtM5R5hMz2KHHcMyJCPeZJY8qUuiHvNcDZAG
XIpHrlcmS8BAnjmmay6zZgKB1KFGFqcjaS4CTWf19akK6k8tHQtg6IWn51d2o6lB
WW4kJ+BPvbQzTJER8ImgHHJPcD1112gqX05A9sJLRh2cWmcTmYiRUvm+ZVOQrDGf
R5ssvap3iYqI6DSAqoVxbh+TXTp1SglxxbgUGRWa4Gkjyo/0iJ3JmtWXdM7tkALs
2FqFEKSZKw8EyTHm17CGPI0dhvaqw3N5IcLXQkMVpoq5MsoNAwQE8exusoWO5Wqq
22/3cot4zrp38Hz0Bg9VyxFQvEtN+N1jmF5ATpzmPOHUFlG3cn0yBbUu9yCPVDGW
+2smugb2l+3MasD559VV1YeGU8Y3xQsXiLxKONCH28kwFvkqTeGLycXgVbJ3nOyU
gfAYHIomTX/6DqmZWyGmi3SH9ICl0DrRmtEbljpLBbwBmdLPCaDW1RvicwDDJi77
N6Jqczvj838g9ITUw9grbxLE3gyvY3fNr2FRgoQ50E0axaIh+zIP4ftBTS3HibQL
sSjsMoAAqlzU2z3gn9oZfsHIih9X/jIfiIP3/yQgNgnvvhitMVOIlElCZ/hUFtnQ
Xz2LTOMLY5+tkqHMwvBkUodKYbaoC1AZ+k0bPvpdhLnHufm+R+rWaI/hJY6l80LF
wcfvjUbaZJOfJ88OZUT7fwF9sXwgCzPSN3UTxmIgZjnNzBA6+oH3cf35Z6Ct2Kzg
ryWtxn3FYGvrPvG2R3fcPZxi3xMUqzhscY+H7uLZZ2sjA+RmWpyS+VxfSCwXuiYJ
VtBL4dD5qmdtTP45ICTRfJXvwquDESd30U+x35MhF7Qw9XTr+SYqa+VoJDf3HrUw
21+t47vdEjyqeoy/2ygDYHJusfMa+Yngzuf3TUg/SBNzOUvH+4Xy/H1bBgkrkmeK
85KdYkY+miFvtHhwlxylGQrORHJYr/nFU4MHMkkxEjpbxZjJjJW806wZ1yUHnvQ3
/ZwJc9dRDtupU8wEEX0V6yUjS5oDA/sI62BREF0MLK1Q5mbhrCSY/5zv8EtV6TW7
fdbaXx7ShijL+5PIacABACKmiWDVy7frXuAqHpFspQyU+46trK0XvJcPvgUfIrKa
FJpHTWXZcg0gS+YbgZwP+NfzW5HMAXRb0Xrclu7ToXpRkPFBbhQ6gmI82W+x//og
rjtbeFAIifFjV0W95X90svE+m3NhQbITbBo+W33cb+/5oqT/t58N5+qx2ufNjBNN
DO0SLJi9V15gGwv04lx4Z5FyPtjo1aRBrtg+sIMD6MaZRqbYKVAfJBniN5XtPPy+
R9WYrodjG+2Sg6tb27HBf+TnL64R9qhKfXUZ/FAQCop9xBQ4OMXBvG9R5hM+lJ5j
hHENkYLydVPYUkxR2AtL8rytd6foTgFPiYCWHJyzciAVZjob/AbIwwQlYvvZBNJQ
ZLtYwdYUepzlS4nLMqYO2+MoKibB7OBpcjUaU6pkb+T5xEQ3jBddgN2FciVt48rU
7vK/OrlJPO8xtRCh1Q861xtWszGjglXe2pFBMJo5d7grvR6IRCdXVWyQ1HPLA7py
JXCiqZUMFE4IMVuMX9N/XKLbkIo+Sy6SBy20WlCan2V93gnfrqdJr+3My5xrzdPP
qxx+7IMRV/iFFPaJ02GIYsQeHiMV21vMpgmZ58WNeNfQR+ElYWhEKNQx/7H40vNL
W1sgcoDnO2NUs/0T9GZ7AM0sEb0YjLnM0aVVP+a4kBuwBH5PbRHdk2URCxSGPSem
aAjIfBFpazGi8P0YjRZfRZ3OCr8cHVW02A8U+XmDLJVtz30x9Ndzwmx/ivh2M0SS
92S7U1H0JeVdlfM5NkHK3By8e3dOHWVnWPDNI7El5dlubCNGsZG6fmJ5b1H9wJLE
iJzMHg3R4jb7WHKve2SdeJlEszABrVujuxTboxfn0CQ87Z/DbeY+2KUv1sfJR5Gp
Ok013qR+mw3TOGWKlEU/8qAr57T8roUGc9ASLKLOXkfL06vcuJwHydPPgl/szdt6
taBODu58WkP+aqUMlJcTCRya1Z2fRWqm0GLPvKawu30qhOp3Iphm8xzsl5wtR1H2
oTKMhrHyFl0Rwv+inOg0c2M5CbOM2Blq0XmDiqbPWcfhdRF+LYmUB5ioMntyzUC1
NUwmeDY4gSnsaJfdE7goQ/RH2tLrr349BB1JGQkFKdj1TyG8ZFxw2qmFz69MZ1O7
KQlxMUXrLMzkWahX4Xl7ZojZM8mKwhCKxjifNY5z4497i51qHGX6fl3+XGZ1HycU
DrBm/b92reO/xg03YNULWvwU+1irVm94vO9WVeFpPygFyNOd5Np6cjfmubzMouKB
MuIZUkcunhUMXcUZ/I/AM4dZM/uBqFet5nabQBUUT4WFKMbCSSVnvTeF3mohQ/ax
xWdEn2UHlvIkgze7Riq7mLE/1GF+jXXFnn7VtHiAFZJ3yQa6EyUQwzr4YE8JA4Db
bT9wf5k3c71wXPGyfywXERKsJbivlVlHHL9HT/8+kNeD3+XDMNmqzCatA80FbwzY
vncznTfojERgG/wW5uCwm1vxHWJqJgsJUZHj+AM2594npnu6HzTbUeIaMc+L3ytC
wlC0voodD1LtFUJzXfJ/8Y1C12WkbATK4+uiY0eFU6/5TUOeq0S4qG+nznmGazNj
f6ACFKbPg6Uul3MhLYb9YvXqAdXvnEeYJiGxooVaWX541g+kfm+xdO3vnMf+9REO
fxsLYd0Om/HU9uB2MuMZmWpnudMVt0g9Z5tvetjanwr2H2WuMVGJdAGudL28OpJG
vyxJ0Oh6n7Su9f7E3pIbe9AwIJkL/HPAIuo/tuIXlKJFirKqMRNR5Kql4HdO5gtv
H7ZcP2M/LKRoWcDa3YlXDmPjrz8iEFAOP8UlUGNh3wwd6K6YOC5D/EtcUHDZp0wx
HSMVrZGDBNXfH9omVCyA0h02t94jYO0Fwv2IpjxtBwKznEXz8ufNUREAvOYHQ2Ib
VgOP+ru/hczzJ3MkfIQAiPASAj+RB44/T5H7J0UUdrmEl1TEP/5BHAWnDKt3wP2b
4lkEJn7mnCUBW+sbLxwXJgupUBBC53PJyqoQ7sN9ZAc7nSD2vWrRTYrhvrDT1Bci
I6/fLE26gBfwD7uw0RiPwXTUc4uOQJlAcTamihCp2vhMFniYTUs+DqTvlM9hzwyR
hZRnAaJkj0cYx3/FVefpyzHo5ZISw8iIOKC5vNzO+SHTAFtNyuI2HlwIfErUW/Iz
hNsjweQNnEPsYeNUFKfvDwPuYsOjJJe8+1Rbo7nbMhwCpZP0e4zTX4JjAYCfY9hh
gupqlOf5jpD5Mhr76K8PTyEy3Qiie+m8S5tzSycpZLV7RqrmK6dlewiCEMN5ffiB
xF+NCO0H19eGS7x1XqDsV0H+GNlvFlVf/v2lWKBfimWDegcjHu3ETNLiaPdRCSaE
VHfI+NyPZtc3FTvuUgbwVRpqm27/mEqZfK4G5w2SqLJ/sFgiiu+P0JAJKLRep86V
rRh6ABcTD4EWz/qJ+TghwBKLkGhAcP8BSmKh8KzJVyVLYVsb4n7rs8llx+aT5FRT
W/E1mLLnBD3TbJJBTHOyyWXCJZhI0pNRx2w60J9GORF8ZTjkaffRfWq/Pu7G9RcO
bMpQuVE+tQuvuhcritW0j8fYtickA7OkUoZLeum2Fug05Lg4U+dxp93ocH/lycuR
BSrVaS2f/GN4q2qqLZSnYLuv8fFk0wk776ws0wlhwn08xRGn+QXGY+45Q92aJ8Qh
xD9B89PRVwSBi7ocsx3p1/46f0PCOC98YMpvqloF/GDzsbq0tffU7tSw8h4McQbG
XJIy1Q95G7i2LtXuTZt+w3Wm2qtKW9UW0DETAFLMtDpVi00XyKNXrvUolMhQo+EM
Ae/HqYy/S/DQWdfkBWbqPUonhXxJx5OSFwOb65+5CEpS6PDdliUSpy9eMgG22fP+
PYlzh63xNZ97J7tx1s4BI3Yc3JelEjyPW8z94f14GcV1kjr94hUFYDMKPamWDmoL
GXlMe0zp6lsbuwBYbzgkgPLdlrNwFC883zBbJNkqBBGs2coNVTYpVQtZxc2Kh6a1
wks9lHlGHniHT2PA0B6kqxhnBFmE77ipBisGyhOuLJXMCpFw+ZQZv3jo3GsaGk13
CDWnhL6+YyRWkOEWX2hgYwpZA0nNdWO3nuBpopnmFNqdEovR+Itwuz50QHHcyvcb
bcRpKNRpWh2ucKPk+unQOwRb0p/Laj4rZKtz18RqOXLW4ziAZxbhzTBRveO7Kj98
+M1Cm4eUqhD9ufSeg2Rb/VQKoi27e/8bB54OGfRkXHG+UBQxoVp03/oTuc7kvkVN
4ByaEZtvwRJpwzlIZatmpfHmVbzObfy1nSSd2tHrfbUW5hQY8bRTP6xM1FnQORuo
kONohS1+UxmSLKWEXv0/F+BZ319IJXAYVrvtc9R2kqEek5MgZ8yw7w2GFPHVDDcX
M1XY8s+L/f0kLiv0eOxKsmIgDsO9Wy8TPvi0T/fSNJ+EG5iKcNvgUR/C16IXRxgB
MaLzTYx4jXbIOFv6CUvy+eKhkhbVCMvok4DoUlqPLbxDYL4Snb4fbfBfAe5TaQUx
/Y7k6p7aVMoL/burfl0Zu7Itwfe5bc4q12jHVa+8syQ+sBY7RlZfghtuJOhScyC/
j54atUX5nHPQsbdiiuuEyvHZ2WcCuEkqu1JIT9lNi9t24K0qo0N0SUTT5Dw0MDvC
OiReiu1xEKKeOnMOvkLYUZYsV0EB68e7wYGmZFj56FPHcT8YU4J2a58GyfYhZu47
SSh/1KKbPjoSIGXQjdml7x3MxoNjgDyOpJ8EBGp7TFpADK7/NKkq/FZtwi3hkI+W
n0C+qJKgOLHA8aGa2+UNOeerGdudMkroFK8hhAkQQ3SW6i7kL1/ejQYJm9hpsq21
2RQe0iPj461dFnK1XEi0Iw/9vpSwZvhVQsZPlUZroZbpMgxyCrVxZJTtC0r0ndeF
E36vykefQ/pJ3qJ3lcL/ffV7Kh9XaY+BAXNZTsANtOy6Hha6vPMz9ZuBjjUOj35y
N+3PSlt0qUrmBHaxSSV2G5FIfuome4fuPEBu5swOAKMF/w7QhNjiZTxQoh81/4e9
dJDITvOWqWIPkauM4iIUMsiS9T34SuSmIwTrFp2pYd3qc8dcuNrv5VF/xzjleXN6
BlEzSZL+XR1Kxt9aq8Zm7csGZTLnhSm2DKiUyHVtLc8uIm+bKyopZMR9fRpUqQos
PopJT5K2913fH6WiwQxyopIt/25yMaNBf4A6UdfaFRA3zTJTLLKiT3HHXjRfNcRo
lagkrvsibnJg2YUd08MSXZBf/bYoGccilT/RIJ25OMAfB6ujflqfnxtpqkTIP672
vsnHpbJ0jK4z5pDA33dGA7+1mjFImfnlBEV9CgqxMDL1a0+vXNvamaThmP3gyHnc
1+YNGES4JSAiWko1hzPswEA9IV0we9LuHEeLHvLvgAILdLEPbPzyJD7q25vMcPy0
JvxBpo2V4s5/mB6Ix6TFRHpYGWmc4OMYhbCOhqa1480/n55USHYkqrCZNrpBnPkk
MT1GrsI7LI8Ju4lcLlhnQHo/Ida5XuPNMrwA9x5336umGuGfIQLltELwHldNwadT
vfXcZmAPxQ50l63wSB/LTxS9A5wOYuoRPEObYRdWpjcohJL5gmTw5IHFmKiGZHMw
bHijXVS5Bz1h3sQ+IKSAtV/CdqWknDK0KKaSSsZgWS8x3X5f4H5l5viOWX/U4DJu
ompUWAAlQMer1QL+9BcJlC3p8q+EEo3C/X6A5vLhtXLMKsg7yOEElDv0AlE06zQB
ckcP/O4uB6j0tBeSJjQxcAt2J0LUcRstpjprGXZXtyqilnaBNePxp1JDofy4h0cD
DD828LdjlySNV/IuWvYyUW5Duj93Orm8yMFw2xTxcgMGWR8Hi885GDubKaGPnh5t
Ym+rhiHbnUPsuDUqutlKLjFPASyMdBMXE/DWNSYoz7EMY0AHkSSOTgKfw4ttG+X6
XEF22U4r7AwcFbk3Wc4H9AZd2fWvAZlAgry6CtSLtDoDoROTJbDdAIsZTOiu6P6U
FuzwUSBKK03MPAnuvGBXx8ScdZzX8xAM/uaANL7FyEYMwjGTfmCRkZuodWwWjPj8
hExcMG19GARrG0UpzK/WsnsDr5TEO71AtB94S4iDcPsOE+wZVSMVWysG4XKc1URj
X5IXqCZ+vfFrbJc6n0oeOHEh/4Lnyg9a1e5qIGNovuYL4ZJ9h+L5JWNl7niVzk5u
v54F1PQbZr1XBnjpA6qlGjSYzOOzHRMZKSY0OiF0m1SyJ5ew1LL3z/mQZ/hJcfjU
y7R/dfPpEJhkbeQkrGCAzkAhzoSrN8PGyN645g4fWw2eBMYERAyCtpCtTykABGBT
i4VPZ8YNhp6VcI5Pr0u6X/3dv1scK3IJaHLa2TiMa15+ZzZAs1lWuYWZF9Sxb/Lk
p7Jypq1DhHlfbbGx4hNGxUlXBj2n6cgcqp7UZGUH0FSS+iFpbPeXdUuoGU/PDjrr
NS84O8NWcm6JWukBse3UTbYr5PgYfCT/ylSZcx7PH4L6dvy1pjd/G++774GMFbeC
AH+ZQpnbfbo28qjHRKyuQkNic1dcDXE9yRELYqM4LwOTE7/9yu+JKSLCv5dJU+jg
QY9NAwAtJgH8J5KgB/AaZdDRUlIhcjxTenKJlsQ/FtQ/QnzRnVfflZfjGcwdebYN
rsI8l120lrEZTF/aqm2uzYVBEJUsPF02TgE23vxUo7RXyl9brCgz7XqvOC73x8pW
dFOVqLe+FcvLGH+nOY9+4qcoD16bii1LYM3drhz8YPBfGQLFopzYF01GgWOPGBvu
z9cIKFX/CNqB1BcI7/qrs8DuVQgJPNGrs1284xYKw8ayuwbJpbO23jTPcwClo1Y+
5kwIUjzChRY16u7U5a/FKmWwL1fdPmidoMWKbb15urDhgAki/otQfI9iIkMvUOVr
1qDm5gUfwyQpn3+/eZRuQep5JGsai73so7kvO1uJmH2+UMRWVQHyX6fpvCdqPl+0
7EaFiOLiaSRYM9nlkm72PaOjQqVVPE1y5KK2I7O1rnqAN1dayWRh7omp2FI1jMIM
rbU9OrYfBuk1qqUqslL1ISs0JhkMNImQRnL3U7qznmlr3eZQ1SmdGcoXy3PuCPD3
jdSB8lQpSsH5ewcmxxfU6OABsh84sOMDksMZA6u49n7KO616Tdtw5CGwVrt0wTkM
UP3LwGzSZt7+wmPnLMF+E/VGXPBS6ivLMG5v6YId8sJCCgNA63Vi6JkgVkeMoyol
Runp3p8jw1TvEr9wTS1kSrxNex/EXNFdLymn0E/ENJ1Qqgbg3xzhC05H0hE3ia5G
7zCayw8R46yGvHP2Uix3cDUZUDNZkOBFoJo9D1NgIsfxmUzMpwI9Wu+khKgIUh1F
HqnrXrnrg/i4jopT5VSkvwe7xTi3yznyePSQErL2+72RNtoi+VwN6TFd0cuOtU+k
`protect END_PROTECTED
