`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U267bZ3OG2ligmn3YzVO48yOCoYiyUTsFDX+nU9QRcAiULBssJw4tQev/MrUSMkX
SDk19fDEAlpEbR/gzeN3YTymbF+mDCC76rF8Wq/Vpt3vsDmA2YMdbYQJHCDddwHK
QipTFihOBI+jKD0JDmC6jTpfdRWnU6L+YHgZyhzyMK7mN2inOf921o4WI13yDlMx
6qK6xWKApKSM/Z7OXWtPoWox+/bYOhQI4iBSG0xgIa35GizPL0CZlI2vxPCaboOv
G8J5skg/MbnFalUSBmLdPQEJUrNw5A518XGgknJ6MFQvMsDQfGJ2HLFV3Cstm4I2
IX/gdKVxgIu/zp0mmcv7kfHU0vQVUIreZuy8WlZij1IAvgWCbfFsSwUU7nvxj+lG
GFYVrPXDZPuIdtEnBjIzDxH8aFLK1ioXZNjIvrFdQEBQyGFABcKqX3GZt63Po/lI
V3OB8GRjrUH6zG+jeI0cpA2x9eC2tRtpj8iFn+AkP6h31GBopGjYyTlhyISOSCKg
ecn8YjRtMLhGJtZWb0s/Ppj5XEMZnz+eklIVdcIN05SC45RivImGw+1CXMrEyx4D
DNT3MtaxgKr/xv42PnnHuM9K1W6R4wUtWfISZp7M/AGCuIt7xAyS2PmuYfmVcC2J
jFrtVKvlWaKD3EpGkURLxfsr2Rl4CuMSqdZopeVmhQM/jJoOMn6tqUIq2OxdfPyJ
v6xOSHyi3m1+EteTJfeGAO4TcViNvhJVK2Zblp3KQNf9sa6LB2IuTXYaX9dxuk+2
yIbsavka2yTTWH53xZnFbLB+LPtg4SfVfOxOsTVwMUUyJThqDelQN+tB2Lm7tIop
dn2A8fupGhN7DzC8nCrCz+LX3gpnmk++99YCUmsAuA+67Rs1z7SPaW3fechGNBCl
5lSzxxwfH5woZl8TblWMdDIRxB0O3lxeVUhuTejz31SCBHPTYAytPs3F2/KmxyBJ
q+AMOS0sXUCn7IYc6+0dDDT08/geuhD+QhqNAw++GxQwZtU08BT2PHYLv+P6nKnS
2lwLYgd55i7EDejib8fvRxthUdUJ3TwyEDyIp5lRZxPa9kWTDshXV4fWQDOHeCw+
FPkTrdRB4ejG7B/yQ95XrUIu0/CCx+s28G8rIJDPQQNVJeseu1238wae0zu1Vm93
ErS+o8LZxQ6Uk4eRi3UToduRjovW2nNk1GsiXoQ6FzaRjPZS7u0UpGQx5t4ynrNs
GFn/S2Fxtop2rmWNkO48Tjcsczl0S60sTwC32s5NYnP5nKrku5/1LmlYFjNteKkc
+coBm3hggd2dQFHnvq53zHXJXY8PvqLG1gE0usc0PC/ZP3y3I3HJowk6Z5aM5JGh
oXQnQTdCRT4kOIXmITYU/bEcxG3lppxHAdPf+XGZjuLpeR0jVyneuqWAe2qc6KgA
JEoN8LlLOChPK+JVvdw5BzPnzF6qlU2aH0YZppDhxmpz1UC9EkqQzEISoeYfMDfZ
WXxjZEDjSPuE0gUsjrjiIZNJLEF5nu/HxxBjjDPa2BsfloJrMXnbwNVrnxogPsab
6icxVaQjE0OqPkKlmWjZF2D3UnGVrKOlhBeoLSABg4Gb0Ramdqwvx0L+MYDAg871
zzBi0sCB8POAqM/cia5Ahnon3NWykOEpJqp7UPMVznW9o4+bmBVjycXNQ6k8JSeo
PFRkMJpPHzaeh8VGFj++840UmRqEaeHo94pfgGFCxIhe7AIeRpy7E3R34Q0vq38T
gUGx6JG01rNWz+jKywP+VYEH1htONDnyucRMkOPvC2qFQhGmmwXeUUkokIkQhu/2
injg6mLkNwJ1aA4w3OQV/+AfFEqJQml6rXmswQUTPUmd2iTZtZiUvKtOYCgBuN+H
rr6FiLtk4ZLkNhXRavNLpETWzaBmjc7vR82IMFN1TSfTdsFkZWe25YnCPKgHjVaL
V80Ccwzm7dKpRwV02i+ctWR2mVT8mK27DI9CvziIYv/A0Ic5aFkx/rZi85DZUxPt
urlEdx9aaaXotyTaoM0RMDSlAS7sZcNgbEtZe570o32x2DyS0547A9WVv7DHIVjV
Vq7DRjVga0+5ccFX8TFNPs9Y4wopJj+Tkz2FU5mx7LvTsr/QptECzCMw9EWyu8dA
hjblUBxWzvrqlo4PkUwJ+/q6Vnat3vfrNRYwXeprxtB7lEsMCpnqUfbNXezDuDM0
NdcYVW7TpNEq9YMfYtHqo473bwz+CnkxbNOCc5oKVpJRnmBwmpgrrs8JIemC4R5G
LmvlLyw/tsK+mMQmYOKwf6ucVzh7ugVVS5sqo3KeljZPH3SkhZqI1Ca9g22I8Nx3
gLfQ2zoGJMDZwmarLVdVJgE8bJU+lytUC7ITdwy1oSOTtf7NMxtG9mmrmLNxUUyr
qEJ/hfAe81+kh9gSEuLy2d2FTLUs4CUaSKiidnKFX+grTQoivBwzZpPaF7+DE890
bDylUKnfyUdBZJnVrgQDfQqw/EFEp15hRPtx+W42Ol2p5Rxq8jNqdupfbWJEJd8I
e+QiMxgPZjWPEAHdBhc+24chOU25shVchVNhY63gMq3aZEV3ku2XxrNPPpR6Ipzz
wexW/eh+TGhxaBsAyjmLXBxle1pu/PCH9RKBCj4ECI9JhLN4JCN91JY3E17zZyIg
QITk6ZuzPJacIJ6RtEfYRe2OFpQDPnYZfAMMDCq+xkHDTDoPSlspOZay8U2eFIug
8qV1h61Tt0qFCJ98fZyfIJ+aYWWgEsQuSD/zNq3Pv4SXtN8601AQWO4YglPiktGM
aPiYTTyBINO4W6FE1EtcDeYKS1t2IGMFYWbK6Xsb77PhkktD8jAA86CtNurVrWu3
5QzGqvp6ub8iVn0ZMPbJiZTjlwwCuKuDoaTPI72xovPA1PtRqyB5dsDCs4zjWAs7
k0rr/wuUnwf5B8QDqxIcUeM8QYjy7APACxlVXFwnSr8suVG5NOTC0KJZXoGWG6Lg
cVdaB75AgUixylLg+9AXuTDTZFt2pKq6x0zLPznF8nm3AAlpmVK0onCX8etH+RnC
zxEaaO/2pVjagU5VKUiFHSDGDUNJkblyIXfTTdsk52o776klH2nasxBsy90odbk+
+8/LaeOXgYQMcl3TdUTktCaXMFEouwxcrBPwGqRBHRNr23VX4x5EnyVXoRertyrC
NrjfMhEPd9chGdG8qaB+9hSmlkZwayH9r8PRuNNNs5oTQ6/m5VlF+WCCJuuMFw38
Pq6ZP/IO+3NirJqvElF/cPJcRl4zKUmOud6J1fSgUyFBHwkKqENNpzTUg29P7DQN
OTyKOvJRuHjNYIHOUpLNiEEgnqXT6B/4STwjlKYs6beJWO0wEfKG7EeP8PtBdLx6
ia7TXf4B3x55PfzVXnAHiWwxH8x0LKRD0yqUOsTe1rFwgfepBFXUbEXGkixrHmKs
qY9ecTODWasbQiUU79cwnnvLAv/L/6H+RvvEtq5FlaDXibUlWCquUY2OoHXcXk+j
8ANsuQ7sWpLEMRFOi9gogLvMffmEbKBSpGHD7Do1xHXY2jSpfQdkcbXY/40F/R8H
9ATalMtFOHW9z+DATeJ7UZpmL1gvgqiAwa/uNPxLoQWf9M5EGG3+USyMNlYXv7Hp
XXe+vco2idwmdl9JOh+J+bIZVjvAVrVYey8236D8uBuVyMbYtY1KuODb+aWLUWr3
iLGo0kwXsQK68A6viiyCY38w6CqDDZG1yHnZfvUKuNg7ttPRJuAQQGpMMWBVl2wj
b67xouY0qV4eFHls6WCDMnApGiO47SG4Gh0ILsUY8UpHpfm58VgqclB/2XsVZpwP
QIyMokAJbOh6FOLWbdPE0/NU02GICWMxlzHTXe4Ns1te7yGMkjm5XRIS4uokW3Fo
7i6k/hYYhuMhDKo6ZbcEXNubBkRiTUzcBPmtZ1MhNG4nW4v6YatDyYsXyvzpU0FW
3TsNalT4802SaDJN1bJO943+AfKTsBhdkxRBO5MuYn0rWsLl8b4qCmAejBJ5MxgV
AUVqWD3SIJK1reyY4fk/9I7y7l0U5kfngjaDlZo/wVMHDiF5NZP499kfJOvZvBVt
SOPeadrrECoFYxGXhDy4L+NOQrsdzdJicIlvR7qKZEB4FUma95sqcpGhCAgqFYr+
DuH5zDJoJTaH90WIZQ6c+DDmOttIdETsYAhncndx+80nprmLXMrmE13YKInpVYwX
lB1KEGE6EUfaOfRuwcts5etr/b1mB74L6ux8XWbQptxcN32EukyOhUuiNsZ4FbgV
NRP2osaQmR35iv29YczxPEtYNW6NWoVtNx4XPEYgOZNwnge01bSuauzLKRixpfMa
C6t6+H+inFdAJ7c1KTznFiuwxwU2Y6wtddaQXfb8dFQJmEOWM1li7WmNxZJykob1
ISsShQ9SdKL03Vc7q2eTxQllVqL1b8QPxicyvsmi+k83n3rnHYnkuhgcvZSO9he8
oSAKngQoJoklWo/bOzr/yR13tAbwzv+PRkooWqiJFZzjqMwnoJt99wyjhcRBMKc4
dRdGD80vCHGjnmXyiSHs9rZDaHc+EsMxPVCqdQpjsPBz/9UfK5XdaYWGjvG79E1X
sPpXt/cjueKjOy4KixcHgO6xC1Nhiye/uhE2YlJvEV9hfhdLvZmihJ36r4Mz7FSq
kj2li7djdkQlDIJyN/quu0q2C/rPgxG7YLJ+Po/H23SzQoELYEmP5RJML12+hED2
EgLt1ouT1G4asBull/yEGn/12DV7CFUZMDDS0OtIp6/5IfER6vlquJtZWqaf4v8C
uXGkNsddL/2KlqU+BpAGs8V+IBfipT94q3z/j4TIRNTzcuzeXzzHw8H7ttdiEs5B
ZWBDJXQ/zB2c4HYUK3pxopMSTV1Yay+vqLhNj8zhDJkBG+8mIJ+DjCclt/WVg7tB
mQOtwKEPXEwcPZdYNO2r6KE2yt/DY2NCNja6uyxpTHb8xIGESPC0l//OHPpmIs0H
+1RtECpWhavKimw4vw2kE2F8RLEuQjU9gQASEo2PYM5wVXFVzLjitA9uofqpipMn
TyOucVBcoGn0P6OY6ZSvCA==
`protect END_PROTECTED
