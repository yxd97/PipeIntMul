`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLpVXgyQCRwjy0CIbniKCjDbTrwZxBnovxdCQKDw6fPPKQ3xsvq6CL3qxdK95y/6
wAiD47MCWfpWpns4c/DYnku9xNbAFPY5IegiSpA5UwiV7FCZl6rFeKtvFtVz3IGZ
2zADsSgVOOYf0hbtbHFOHAElfkJU0WmjmE+2Wba+lRNYnjNCycLHhG/XYPKuHRwr
KEXO4Jv2GYI36KQMuCjnN6Q6S3Cvck5sEIXSxP2FA7k9AbChG2IvUAu9q1U2sdJl
rANbv/pfqKA1HU4TFbT37BFxEPtqOWAy/v6LJAqUonn2yq0s3E2uei/1qFHnVu25
w0ZzBrwBixNFg/v9/crvRbkXqUeNV1i+BgJP7z7aUp129PnKPqLwez0TmMY5ZonL
lTJEWzJcxnNmlETnQCBG7+Z9XLs2PGyYN34Dr7avklIjZJZoBFC04MlcJI7QIOBI
`protect END_PROTECTED
