`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzJtJh4n+2PjsOzKXjNJvyzu6how0tJ6pV6KCmqViPxDh3rZVg5cJvbGdxqn1jd9
5cp0VvbMr6Ksj1na6RKdbzC7Od2zs/NQDzpOKRKcjwLk6KH7IQLYdbCX6YpID7Rs
la9qdceAdTVfdGdh2D8FksJrQbDKKfKgmMlpQf+Wxy/lyBi2BPxTdSW8QbvYv/iM
a1Rp0stinmy+W7M2zisW6IsuUE/oEsAPdKP8q6hPMC8OZk8gnLeAOSf6o5ChELWT
V2Imyoh+zq8VGKQan28dqtnn2YtiMtKNUxzYZngE88Ai8KfT1iQkUyDUdqv/gtmL
iprhoUnQwHFs5iPgFF+s3QtMtC/WP7fvpdySmK/xaBtOX7jU5rsJNzai9II7qHu4
ZtNgqzs85vAoU1EPx+rPdDDRrFe4RBsdnnYVs1Eg+HNYNvdoav717w4DxmfGzZN4
ObzpQF2UgLkxhB3o1C+uB47J8RK/wXzBtF+s/U40KVq9FaJJQTdnezMOpUVX6sfr
nw7UDf738p3ds1jasgiD0QuOw/NvpBsEmINgJMFxlcW+bPW4cYDPxEOFW7Vnj2Rf
ctsB2ty0ngOzRpQq6LnF/3s6u+nndOFyX/pd1fJNWAaPbTDLH0QbiPCCzgdVwZHH
NwKezyj0h7K8Q4yWsVrPXh/8J1Mv/PgX5X/vCUcDbctPce1T2JOhtH+bvgC3nEbW
RfvtTq8e8KnpNC93iOt/YIV4/5094wtL0dgHxdAByI8=
`protect END_PROTECTED
