`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k1mqAN7T3HsQas56EZMK3PbK+uh7BZ1sfba33kNwYm8xtlV1HVPQomQA755JCZK4
5beTUPPHr+EX9XE/oOlm8MyIf/eaEd7JZHun3HOaT+MFGEdMofAo2J02kw+rDbLC
hLz+8I6w3lPjqzYVHQhyfrd9o7twhUuQ6eVfFSGFEdaW+RAL6CuMcz/cZaQO4D/u
Ut++A7WdW6Zd4DBVibY5GYvAs/xicpV5lWK1xRksc1RksVAbN/hzvoBeX/uJEf61
E429Pj5WFPkOt7uS1WlAC+guZT8mintUR9w8KUYvzOu0lIJv5yqsN19w1fdw/Us/
jMHEXvZ1GVFiVeUTh2jAdDVTT3VEP/HTsuSsTX+pIDLVALUSYm+iUwTLtXQYTGkg
UTYZ8+r1Oed3SH3F7Qen7D9axabmNKDDGvEV7cUDJOWLijNkpeQdvv/of/sgQLB2
9Ub93tedrs+8aMj/OqUWxzwSkT8dNnuwmgTAwYrO5whJb78zxXJftWM/pt+SxSIb
0WW+UkI9FAzWWhAiUEsxlZcRc1Y98N7V0xnM2t+PQhUUCtUgHZo85l0gHgYaguLn
UMKoQFzNEzEYAWl+/jQ0jUBtW81yqNBzGo/s6XChhNJCd1HppMF3K1eJea3ObU+A
JETyJcpczwVO39GQsyZ+LmeUprTozM2TDFI2ARTKpY/iEKkbAzMrCZNSAfvmGepL
PiyAV3dvRC3r5QRmnfA46qnFjJYTQaY2djH95gnoMVOGetV0NeW4cIRFQUaP3Ugu
YCepdqEtmAxgrj7vsuyAeTdcew6G6iQMDDQcE080Yfsd7ZodgYRjDjnyPyDAife2
3gDEjkRsPcg7tEqR2Y7GEQ0aWCufV/ba7wEphkGmmxk7JfY+A8DY55B70Lt2GwUB
ZEULU/hL3m4YMnKsRwt1P33u3OUK7vNBXdgi+lMEWT6P0d9vQEEV/hak8iV2eNqL
lzroRCOEpXiwVM0j/RFl09RDRbuBniwaNwnaGQhiNDHwSd/TNDDcShFUwcDFy8Y5
i87UMfUcO/PEcfSSI6cFHtUV4DngKRjslhy1ZJiGQF12IVCIAcA2htHBSyCKmNnP
StJkK5xPzPxay5RAdOHshKN2pjIsiFMMWD8011+CVx1sV8UkHpgc9wiOuDNArOPD
SFMNJYajF2NlgvZo+lOpRl8Wa4c9qo/qbHoLMBkoMMSub/PZDRzu6MO6WX/O8dk+
iJWXA62z5w5/+EJkCFykaXaTyNYW58rDITMFJl2t2xevkwZU8irmmQthD2JTBdsg
eNiY6FKAFKtL292EAgwgQUWpnZJAkhbWfO/8yNbw5DBkYDvLUCYL8U8G8Nevgy5D
7bvGazilbG5MO9Hz0LXbB9BoWHV17PjM0hIH0RDToKcmeHInTis/JmAEOhB6fr/u
5toaLgvW+Akp9opaoIoTdaku7chKV8G2nefEoGw03Ks+bHiH6LM5hM933lgzQjwk
GFX5zCxXM5P/BYK0qY9c7b7PuIpbZ08HXQesxXy26CHbMzXcgHrfuRpYrPDyP6ST
DohD6fEVxoFz4dUCxSwSQHTcxfBjdK1dHbaiSYsdd8z/HpTsIHv2YlD4+lymRJJX
Gp6LQV2BmIy+quhpkj1hCgfi0pUpWBYfCsUcx2NWlKLqAdjMcynEqtwdCuOp3bdh
DJdqj91JdEhYgZXl319d8fBiDI89JjSzpjchBZfK8l9SJGXZ7oLxNOjJLFsl6HqS
G64oWsuf8UghrkKj6xd7n10tv5mN3P0VJs1yZeX0OSamiqtp8TKOn/n86bJpzUod
dHbDocwPf6AXx1r5ce9UFMBdfrQYpJU/iY3uqRqVD0/8+aHzPGV54j0FQQwDH7oT
LDIy4xc69J2SzmnUK4rrY+psrw3PT6S/RNIRPEwyRgWAfWOX2KyzEVweoj9b1RXO
/sD41fiz24HFuluMqZ1mAw==
`protect END_PROTECTED
