`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QhOSUZLH3yG0NF61iYCvG/hGhGJDUlh4mAiwMmIg5E6kN9w68UseUY4IcD+85RyT
vRsOsEQAdJ1tHLuCnskN8hiUL3nMvZolEk5JbavvxbSM3EGcCS+gY55fN27mXzyh
C2Jyyryyvx+TP5DMOQFfIDlixJ3BwfZFJNOBDZDS6GMAaFGxRnEpiIgwQ4M5Dp6I
mUpEDuZAxtXQQue1zJHXM95YYwFx4wm8NAKsWfeFWL9pbagtZHOn/+35BB00DD9B
OmF8CrzcBa3bX8uhqh9MBw==
`protect END_PROTECTED
