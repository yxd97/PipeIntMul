`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/DlVVMrNomK2BFyvgg6Xo35gTo+R8I5r90zPIUfLsOoLVE6ira7JaqIvWi0jdn0X
c52at1Nr4bDlD0Kzu7zRp9vnwZ/aW8G7smCuxwxJv0ayZrS547UYxOYWr2twkmCO
cqKH3VtVIUyYY/xP6hOeO1iFXpoulA23wTP8vg8Cq9N33N/WiaqPq+Y1ukorN2L1
ncrIh3edjgLbic5zMF0qLrntXA1FyD5BMCCFm25XwHOV3rG+oEblFfb+ZHwQgCZv
qAWXmnOEwxRs8TTcCUsnHA==
`protect END_PROTECTED
