`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2oA30Oa6gfzF19Z21qgjad+Gng5YSDgXO6+UBO0EquDyyMexVccZJhpmVQcnXBz
MectHmMWCRftAekVgC5p5gUTgd3nRLIEmNoBAIexOe8Wj6hAPrcy0wOt2FK5N14n
hcEFGnde9WbgYoUcTodI/CSUZ/QCW7M9nEz2kP7wU0zbTP1xOtBuyyo40dKs8/O5
iD0/mvkvF+RfJCdAsZrO/UrMZK6oFrERWZbsQgE01BSg78RpN5r7E7QCJoDqvucs
DhhQF1lkwv0Q6v4Bt2KQuO+sYaBp4FAQC2ecbFCBH3Ose5MrxhAEhlk6WjQWLrlZ
3sQ+cnlVVP9+DoFkDO+zU2zxnFWNUYMhttXF3R/ptjZ6Yc1ASh7hE0Vk21Q3y13X
F+hk4LM1QDurAE+puTMf47bTsKVW5shKZrQNzN5wba6lOYU1FIXcJkTZT9OCrbmt
`protect END_PROTECTED
