`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JNoGp+JE5/LlDQ/okfcAobd7ulF5OJnDDs9zVAjtT9EBEY1fKHIyuhCUWhPxWOdF
xRSuZLSwabLOxNwO64YKfDIFWT3FBqoQ5FSGLSK3MEljr0Y7jvO0o2dO58XIDPpZ
dUaO2hjQnDJWL7HdAEgdkm1UPo1d4lkfAgcGrQUtC/vRgniS8U7WmLEQ5aXZvoYF
bwG9xKtBKVVt0S3wQ49zW5P/XdR3WE60K0pGA0OCF60HWSihl8gaIkav5zzqWpd0
sigUB+BRVQqddYojql9cMbt6Leptg5oAruAHxpngbk+OicnSXJK2+xPzrMN6yaCw
+Fq337WzWEWkX4McvslzSyKyRi18TttKMEFigHFgiasSS40m98WuCHwON2nKm9DS
vDRBDgwTSuo91thzzUVMJch+Rdfd7HCx45v+uKYg+1A=
`protect END_PROTECTED
