`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jtvPFIoIS08yqFmYd3aCDQhIYJTW0ic+yJWA6oJ4LpUEjZ+HcaeXKM5HgMXa77mB
wVmDohU6A1jz64OCK+i2KS9CdsQZxUkzQnj7bTXFmGU/Vv4wTHpjzCy6HZU/InqV
ly9BYnjBV8ZewTMAS7pwy9NNy8OFKi6GIKHnMSSXp49cjqRdt0UsHgf+N2R9F6NK
EmNVPM/0HQ9zCawVahdiYXy9AS1X1+PBEX2Ck+n2mzJqqKWcefydJKFZe5hiehqS
a3heGHc7hs4Alj2xWgBSNAVw19b9kTotFNUJwUj+I2LmmBxJHY+hFpj/S94ORaZX
j4XBcPA7WBUJocUmh8yM6jaQLRGPIwlTP31pCFulvuyv8ijLbW4wmtMwq8xEruzc
73ZCnUM6iUapZEKN5vULpx5AXZh9vZ/Vj/uuSVXsf0JJoj0chE1cZJJjR3CBDkAJ
KZgPJGi9gMcO10/P/3QZN3MsZkX+XDna3kofgu2lnoHjemG33R3DrYdgevFirkL4
`protect END_PROTECTED
