`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGQkiXk9BfYQ59c5IsqSP/OGre2MC8s7aUBUiMegCivc6sOzU++foTTMcdrAcnVt
aVnySHnuI3SPoD83Q3ZEFpeE+PQ/fV9rt6t0aBDVOCapV9xpbLsROI0h2EkFuOm4
ogMhwwLTdpi9W5LjBVKGXq6t98gWLcOBbf470r1GIT97s9XNY+HiROlMnNid8p9y
cfNtR9QlAzbkYgwynT09aP4WqnmuMh73O3ouWH3lNUpCMRdljg9EYg5Dw8xe9BWh
uIeOv8r6sz6yLzJjY62G03CpVW7jRlt9mKYgZ1PGZevLARiUi4dElHbFGBgYOeID
wqfDYyYtsVWIuN6SY66cjBd/8ZsvnenFim6jbBG4Fx74HLGNk7LHSKyPbqYMfQHy
eAidIzNh8TYBRhUxpSRv0FbEV9+vU2P0McJQblNoLk6Cc0R+BTD/tcwQyeKwf8/I
`protect END_PROTECTED
