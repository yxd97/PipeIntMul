`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TcI84ghEqTQjKzNuQBAQULB22/9ImdsViXoBpXX3UDYNzdJFmQYfKeR8Pbrt37BW
Nusf1uM5Ldhpkw3SymjEKzy0dBUb3kwWm4tBZ63nCPHZ12qwswy/DNeLwgr7Snmi
ZYZpFvCjKbqVA4gOkTEYgKzkhr6sPa6ex55WCdeBMV5o2aTGKUCQp75xT4ILuxzV
59Yn8Vb8YKfi/j31/HXf5TH1EowTKVZwB/kpFmmft8BGj8o+DBzCQqqfVEkg8ZiN
rd73kMV8MBG5jkEjKPbPsl+TnHY6eeVTOwn6bLBiBkZ+tvbxdHyIUc+eluwELzM2
YrRHhBveOHpe1j53ieTfe0GsDGeUvYace5Wx/luCFaz31tLfFABS2vjZSTQE0INT
Q2JaDVNtYhJdGGHIUr7UeX9k4Q6uenbHS29N1EA5ogHLWH288vfXAP1PyB+23Syo
Q4KYtm+SCh+TG5xWYTuUXpa6/CLgW/FWqKe+2FsMckxe+L22N5WFPsMCcjmK1x2e
XNx8XMUeMlR9HhJFooA5PPWbKwkwJTdHpaIgTJKsE+YPihm++CgvNorqDwTayAsE
BdNVuKP0JGPXI0bPM+j4CoPWJ6WeAlTCLJrD2R0nx+8/BSKm2mQ6LulYIBWCi0ak
yW3zc6ycTNbJ6WZogms3PaSUd0FnEGhrlmTD6E3rz5An6Gt7r7DrqgZdACbmeOfN
jjVP4ZZhoxZjQM6elbGlX8HCo+4EIKVy0pZ6JP7YL1q10C52ppBjO07c8V+alhne
6bf6pvbINjtA+gTCfdcIqjBs/gmU3K1rw7yAj51L9MAo9/uzZl7Vf3A117lTQV4L
UyAOjuPg6H8yq2zEJKLdiSpnJgpqD6AnSVk4IUBMh3UQIEtqh9llw+J2W7v5FFkf
dm7Gi32UubVAy3BSj84Q5Q==
`protect END_PROTECTED
