`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUeEJXF7IBBY2Qzb9gtzow2YnrYgefMcOE4A68t3PFu1q//hNPV2M8VtnMprgsuZ
mYBBe3tMDNYC96f9t637aqqYc4erdMuDxGUB3/ukZ8oVnafdZNL74lsomuMcFWPT
4e7b1NAD6CRCBQe9uuEVQVam3Yzey2a7ibtEd0z0HN7wgbRNHfZBDJHfy+BB9UcE
U1WOlmhU4O+OXLvPMsEKEjH2A0Io47Jn4yP2JDDylxkvfu851MszA9Vqh0wdWExy
J3HeXYySeXhJqQiRRtq6KSI+jCN4AF+7KMXVfvG8CGw=
`protect END_PROTECTED
