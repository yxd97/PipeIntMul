`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFlgZw0YURDRqoz4L5wyX/znu2U5MyvgQhUyzTKooimk+XCszZLzLUxlas2T1zYV
6Y2P5RhnBkuirxYHCohvEToGl92N+GBpgHS86za0444M6pigke2oXwxmu+Q+RvzE
tg2a2FlkbYpPyo0lIwcHv8VKbSkAsvsWihGNMKJHb/NHNP/b68veZaAbq8yxjqO9
jApnYcrEnzcMGXGL/5zd5PDAchpWnLJ8G9Kp2Pm3/mpPx3KWI66Ho6Q3uziY7dwW
WQG4JQVta1v5Zq1UWM5ZF5Inss+GOiHyHb788CTt7yWzgp2tZh1bWIOHAkrrf1fk
aLeTrgFDsKQWWbDhSIqzew==
`protect END_PROTECTED
