`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LegOTOhat3swMAWjKw0tyCPlSAAEi3fYRXFtyJ1I3bd3idz3exmrryd/7S9iWUvE
/WGTktqO+sYrWwiX3WsUFW4yZ3ytKazvfH6YvRa6TE644imChbLhb2ulF+Awsjjl
TFFpeIJjjgMSolKhGfF5J3oYDvbNeAa945RO+hxCiUfSugqTE6R3NnkDeQ1Tb2H/
+0ghwF7UhdEriS+0WwWTnyUZKejfmtNCq4wL8bTXPXPz4Z59f/UPpJARkdHvUvQr
iCWi6VRez0ICTNahbTkgo619rsWn84z+55zDqN5wwOfW0DVJHmqcv1ZH8LCDqR8Q
SQOOU5LriSl5Pfv8gkAhL/c2Jyg4AqKHfnX9B3NLZ1nc/a45j0IOINO8FfL/2gGF
RH51Ic53zwdHzV0cT36NVpkQjTDREKvk06g05I0VCL6Qe1IwQj7VsSlGBQWrCoWk
/cW5Go+MpD4hCTK4d9Tm8T1lH0LM1aiVtMnHU0AyvFP0giQmaR6zRCxmmWaiqd22
OlqXWGocqisSKO5M0+hwQfbZwqJOezrHLqSCjXNppY8YFWeHJh6T35FVKTFoplWm
Xw9J+/smHIICL3kl4yvaEHpEDWhJ6P27VIZDmr9zrwJ2aF498ToPZOoUaCAuPAgT
3hCGC7ofsJOJGjdiWdgBTd1uJ3BoTF9XWYsgLhIVahU=
`protect END_PROTECTED
