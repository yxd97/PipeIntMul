`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3QM5b08Sd/7jd8vv1OOsVPH7d+huAQNKIrfItzTgLTVmJ/dH+Rprc+QwYYxql7Oq
FpRKr3QqJrjvX3Cj6SvpspQUEyu7uiucWCLjBoOEf1MU0jJuldA5L8Ofsj9WV2/P
EWoZl2Yeyk39XkO10XQ4qHvjRO6Z+5vKU6h2sxAsNXA82IBxiIfLYtw+Wfmyw0uL
lwO4/SCtT0zEAGtt2+vzI67O8b5KoJQK93X6jUZP0DbMmBbl5eyKLM46x+VtY2O5
gTHVU0LIMyjqgEcoJj8JdWuIlf37gxylQpHf3qMgJHxNneAQz9XVW3mpQV3/+oIy
5e7ebJeSLTrpyOksiUNREiGmUW1M/znCzjI1L6EZxwe3PLq3CoZyC6CtFr1yqFqt
SXaC84z0yBqUA+IanSo/iZx7ALV7LDtn61wFBWhhX9MEobg/f2ot7CICu0mP05g/
2AzPTCSlM9PXng5m8UdBsyKvdQpHU7GRhqIap/uAe321p5I/GL3CjSdENSGRkUIK
r886ft8PGT9a3Tq7ljhvLLTz7PW7pAAQoqwzko8uACITv+lNiou/x5sBmZJSYPeh
CF+ADQE4Pi+n+o8eqfVA4dL6y4hEqsOliqh8RasggPGJTcMWA3sJMx9ilBlOR/lF
nGxYQx9YGoAeNLQ4RBaUqRn71Q0wflIE2yQQ+9mYJHctxy6BapBlpoFsm8Gb7+e9
f932Hoq8ZLtYYLVRiuxNDxfQbSzxRXkfkoni/01i8rax6tpH5e55lE+eAhiA3gQS
8i98UIkvPnTGJKjTTmjmNtoDUiqKXmhzG6Cuq4+LdOhptaz0Cq4BjUYjt0sdyekk
pMJBtPB+tDwKQGvfxysL5V3M/aHekxDz7BbibxEm8bemJ+KVxK2tcwKxq/hos07B
KpAwmKCRvsWSLdtHg87NigxVwTwNptI9U7f/JYhYjOyFEx+jyJQLsvjoXxrbzebI
KKn34Gt0iQ0P77a9P/bh3Slnc8s7XZiqEqXplp/ubyCK3Ux0Hr9BLyJSnqH+YNs2
C3ZMv4i1QkRuBNiY27OfilBBCUS7YFGqABVUHc57mywpvqZ3ZHaW0r7q6TZaPi/7
waqfYRSaQYebo90GlJCQwgkx5jvP65BMdTkxAP3R92gE5e/ezTjduRS0JRzD9sRi
scc1U0JHlTcjzZPA8D41QV7AZBmAqBW5wWlnNBEnfJTccn164jh0QJGfhEwe4egK
nYB2f31sflpLrhNQCxRyHBHtc5ANEKBoXl5RpcJ9uhOCu8xx0mjdx4KdXH792N8o
OiX0loJK72HH39yrRaYEMJnPNn3pJC++yDx0NMURJBMEPFfm42K/rbmFsNg+5Bov
CjNgHQpUVTgDAyWBxY2Wm/zJQIFk9nV8eAeA8BAJ/mj9xLWE2BQSJdwhUmarn/R1
FJXmcoZukLO1/x2FY+brjzn9ZjXJxKYbU7F01gDJkMTlusxDHRgDP/POD6bwhklX
l5NT7Ij3sMm4gPaaCYvwhxPDVRLF5YvZVWNaQJdgkUcYi6hpUC+u9mzjxYWxSirk
CzdO+o9ekqxoA1ERIxP84df6ZIFZfaz6VBD/QSAJXrUBHKnDlHkodjWk0tUj3wlS
RMmk1WJAN7ijjmqhCRTE0NzmjZno5cw1SlQGEe6DgDNhjBqK+Mrk3HrRvVyG8qpC
556OqxSz0zYF2Bk+pbruL6GED8pnOLbW3/EuNFauROLxKG+sFVBJkkTdwLerBo5t
5F8L2hJQ1HVxujyK1vs4sJqAO7SABMnCZ4vVPhcQLkl1kS1X00B+H9ofNv5GnP/Y
wIg5+J+GLTK8aJ1/tFO+7nK+5POT1aVosc6bdeSyJjmnw0MR7L55/ryxa7gM1Xgv
nVl9HaB5Xr1Kx2uUEN4xV0U7OpiUR7A+QkUz48o3aTsm0EpYJW5Y0QV+kVdPMgvD
Up8U6vaFKRmLwKpVamdvsbcE6z6+8J+6EOd5tYiD5fGCJtiTim10JS+ZPUEVP0J5
0QvsB1iTZAPqqJJHV9G4YXYhN9sOYpb4+DKjBGwlK/iOwW2Ihr9mZpdUTKFXSmNq
k/7yMMuhvHrED92OCgwNflVk/KsMuqAHcmSMK9HhOz5honz3sbsgKilyjMA/oyAm
LMy43Yj3oidhki00kdPazSs8LtXhaz28F9mKReDp+j1vVivoUSR5W4E6T1Nl+vMO
NbkS+VnBcmN4YvLVKq12ZXwYSZaHtCTeUbwofd7CGRZeDw+JJ4lkVX3Ft21f7eS9
6Bfxi7wNe9fNzps1UjH9BJ4QI4SiBDMAd66N+bkohHzzJFKqyqx9v5ppjPshOfmH
nk8ccXV5z5gsgptdurRBxraT0jpGEmdqva9y51tpy5XZ3bNQmgIbrD7bL4XyPJX1
/7C2TpdVApPq6PlGAsQ7xB1GVb+ivuQn5/L1zyTP9Nx08sDF/ls70nZErv2m4T74
0kxXx9w60T85hUnljXmbi40BHWWUpSj1VB+gN2/T2/KdYjFgQH6evPK4AxeBWZ/S
YcH/V3p5HT+bdF7TRCFih6SoR3+fKQqG0iAL4nPT8xnfGv5QHn8in5UB2pAyeb0L
ovFN/rKJfx9qDgtA8+/TCCdIFxy7PmTrR2UvpY0v4xN1N8tPzMLndYivpNjTgf6P
eR1vbZcyOW2WDW8mp6Jpl/ozeNNHsXu/dg74p+oDvDTVfZaXr0nEd8ESioTcTPMC
14TcPYA7ZSd91ONPwNYI9C8XzIDaIsqWOJ0Q53rKdo/IDmqipyLrgTJhaJIGqCzp
3S/ID2z1gbyYtLAi8Y/tb4rixeydQUzvKRRWsoXjsMWCdISQnt556nLgYQjt3sUZ
7G2Tmdej1oF6enK8clOz0WUtNiyqFnCHI4cfM2ZsNVOJTgI9f/xed7J8vNUJGAWH
L2ONJ4fyS4mIRlNU7NPW4Q1BLjlJdb3nulGxdbp6qvFW5aGD+Cc1eBSqQPFF4N3m
I5N3Pd0MWV9YH4BQZYB6nrH3Ueqlh+CnhEL0K6TZlmspCx/PqYaZaw9JcIE9nen9
858Oz32o4MWV/Z3feO14zVIpUCZBJ36hHp9A7qGXVXZHYe9V5I7gCPn7Ei7bS1rz
Leu6NFTXRPe+L0ZmR/PMWFqpjKM7+KK2yk9lrTMeWqBHRx1n2q5ol+suXZJ7/mRZ
sE3zhlEHErNFKQCWOH/G3Oswyq0mwreqUFlzP/SySUIxuhWM7b+P6nbwYr6d6Lwz
sORRiYau8fCVr26bUQda+SvyWbTG3iFqZe/bxy7snguwibrUHaSxUk4yDkj0hCbH
yeqVJW6l/zN1jFzXRbEaemx+42cA9W6eUnCwo9bZzegdkdFwCZYfDvlsaRoVJVci
OhwZffRzKI7hKYV8hEM+RlgGA1bI9pSXS+rtXh1FmGOpuseUYTd/Ntp86As6qkeY
GThFtQgghI9H+7ClHZessw/+2sSY9L+8hfZCuP3m53UkJLlJ+b5M55WohA13nyJD
NKymnYwAAd2+57ql2TgkZ7wXtdtN9CQCZqric5sOYQMZNXKl/ITWrgOoYLHmgGvj
dvhlponFpyFDt0ILJP9vJmlW1JfoIVsqvc+/sCs+P6KoQZ4GPoJVSj5xXkS/C8T2
NINA8rEubtw56RZE5bNsgyC9U5L4C8LETuuUjhtb2bXHOaxZjsot17CKSrXyeC5k
XGfR053FEsqArkUS3wSLn4V/pAmVoSH4fKXOn50pKjF1jOqGEz0zBSSGTjLO/APD
x0dI9RL+OdcoAPSn7CLDW9Q4h07WIl/A7KsQ5TDe6xGS5vd1HKR6Ty5JWgbjfZFf
rRhUfXsyMI3G9WTX13+1XI0N9hQtFcCxINIdtAZRlmTPTUcAgejjYW952FFWHHBN
4CH+ab9b5U3pMTyMc60mlYYB1Vs8vcDnNC9TpqJBm8x7dxAMSSjjFKSQOQkRWhVQ
Ow0rduoGJ7a4d5V3CoWFVL7lxN5aR+jYI8rgcAAkeg+LJHSjbeaBFOVq+H5810Xl
BKam6QQvHmICy4wW29HdILaJZ13Ev2/7+G0mcLpiNWPMkQb9L6sOkW7WGqZsQCOh
iAXqnyBBlBgUH95iXKvQDUIwAm0dtotU4JrDxdil/vRdp3OZET6muz6A5f493Nqh
st85QwXkUqeTPEa+L6kODmgdwIADgaD7MKF6vQB8OvpG9cWiuFC853q6Lj9BKcaN
UJtMQ5pFarYUAOaDUi4n3ExwsepliRtAH7H/5Ofxw3Qg1LVzpcOTf7G9hVF4XwBs
T543bQfvqwo5h0VCljPlOJUk9lxRuc9qcqNZ/PmgbvFjXidVGEM80kA7dqKfm8fH
vY0SOhM2U+xgqMWIqXs0QnOnIFqWUjVQYRhVHngeKSm3TXlu5BvmN7AaRAgsPskT
AHFwadSfItEJfRfZVVazSAF8RydbS4vIFzZXJaRxcWcFVWrYMqIlSIFKzHonDXmz
CwaIOcW2jOAUh9+UTLCjt7feOLK6VQkAO0+fXi8xMqubSudum8HVV/woONrUfpdZ
jtYNNgfcT3Da5u6f0ZskcyRfvYiZAvT97pcEx97jyICPCIn5HKp/QbFzfJe6GuN4
g6dple/vPGJ5J4P0iu0AIQYHs18lJXnFsVTPYFZGevrSJ15wsJT+GS6ZRK4qZgq0
R4FLGByZi6AoRFZ3wqC30ocwUuJ4l26rr2lJIvUfbPyhx9/Bt17wUFAcvQ1pk3QD
6WH0fIGIzpVgkNE+/Y0SY5w4y/Lvo8V+wlvTCCZNGdXsxzroiNJUyCn//VJoipKL
kpChbZhGgDQW6eUDmptdZ7uwyMzvBbOsvcYEjtt9M/xbAgbugDXPGuBDFkvQDe4J
+Kkmyk9xdygltcC04uNz5aBbPc9NG7npwnqo3mmoRyTb5YXI2DuvrFhzZbXhtYki
j86hlehsNu+YqeARzsCmmpzy4KGpL74VPIZmUAhIuG0Hi3302y2y3HS/wnUHs20U
ruNWPa93YRrVOGsew00sg+m6nbqBTSU7LlosY4fyKmjfdRgsaVFwN6u8nAxs/3sA
IGUwqCMaQiST6H0DdarSoAR7SNt8edpixRURPgh1t5HLBJFJX/McTzccpmyiJm9e
1fkzToAFsWMAUQbbrdeH0ZuPF9EayKNj4Fzz19t2C0ghr+PaMuichSPW62HMRT2y
bFjoPA4O4P2bjRPH/maoCAi8wygcMcKxxIsbQ8dX8mFzUFHj/ZR0O0WmJtb1C48I
nycDnFdmGHSESqUpvD/WYi6/DTQ5bFdWx3PR3loz2GAJIJhPo1ckuJn0A9VpRqEA
LHeFmYhYta/NAWp/DEOUcjcd3GPryGOVjGfxVvIzJZA2h3dTZgnYdH2rOmw1/MIf
gSAD/RvK6hULEHxWw6pYpjkHbnkvGYK3Hd+9Gj4R0/U/rT1VFpJYA2PDxgRKqGzm
PlhUII545j8YIgaSEbxdD7i1BMtfcxCmk8aVudYVSy5nqHPY4vpYHZmOYASNfBRH
RXruGEsiwTChMgTVrU/H5SiFpf80EynxAT3C77wKeK21xVg7cfa/UZVpFg2DbE8A
V+4TYCIsXKdeIPxus+nl7KbXkTcgorFryrGdxA61ZGEWeD3Xsrap0Ejkb21eidXr
NPMYp1j81FQt9X9//hnzBDEApxCe1qAkLTUCyN73KT0zxT03j8rb8uNwGX9vWLwD
XEa7GA7qstriISZUoWifMHlMMW0LSmEWhY6C7pfShXd0yutEk1SVGvEEohrcYP9y
gWw5/1Ojm5m5/WdonbAxSaZaaCbrzT3sAX2pXB0Lpsyh5yjihp/ViEOEOQFmh/ae
+9uqz4s6E+ClMKi9+dlDX5zDpceMs9swrRHawxAZQL3WX0ZzNYj9MBgLNHd+5Mh0
+/lLgNFa8nApeMVYgv+nqxQxXEpilYzOkcWUAQq04kbmjSRX8bn8wsp18nc2WyEW
ytIcbHu06jPyzG1+qq++QX9lUPJ1f2C+aUT4w75QYYM=
`protect END_PROTECTED
