`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sUnTK9yzvloFaGzZ0M1/ebu45GuqyZVVWjZ/gf71cOndtNDBB3RHJ8+iuNJuIgo1
p81JvRBhbEAoTRn2zfHe+WciE4x2//dlw2rUIpI1rr6XNGrb+t/D5Czw7F3xGnFT
1URmdrdQlNV29bUDisWoA1iBuMghd64qQBsNV/2Bw13SHMYzBsCWD2IdDMQzPfZb
xjiUqYg9lLfrwBaADtboXyXc71BWxBYkc38rYUb0A40rFOr8YQ+q4yqMf0QyvPeB
+bjrz9q+nVTdLTvPp5kWtRs9bOBApYGnAIL0FMl6opJRauHx832zWfCcY53x9WC8
F5qxCnnuyzCw0LB4QkFMNhRLDVqhPSODwgDUjE4F8pKLA441ijxL7nDrPemyvMK0
luavvxD3Cb7L3Q2J2GMQfVMU4sqXlJs3zSjtA9d7cJqrYz9inIk8eEgcw/DJ5FFr
oYgtc+sOq+3EcqXqACc3taQ4CNAXMdV8HSYvuaMFhJmgmo2dpao7lQVHE1CN12YJ
veo+AVbaBx1AsQ/Xg9cHZcNiS0i/xvi2H7C4PYfnKliV+t6kuaflbPwssavWn6X9
C//srJKE8U8SSMPnysVZQd9eMbN/a9W08APlRKz6IpL65bgiB/wTOi3q1+ko8jT/
LA0RgbCVhTqx29rG5kVrPcDhUSKzB0vSCdVQ6c4Js+U=
`protect END_PROTECTED
