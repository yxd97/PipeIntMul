`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x8b8cT/+AXEDlE93G/cjmxpDzR2oiCsBRBwN2SN0cQ4OzewT84eFmyJeyZ0OPROG
FU4rp+LRLoIkNAQGyttLiK2+T1z3513Itr+BsWmk5AtoL9cEuJNUxe9Nz9bo9dyT
Cwst9Oo7Nv3RQ8rUHFM/4DCzydGNOEej8ReOzfVWkfvXayAKWJzDblcXZw90GVYB
iJ4GWgu0JnWKiJDEgfQ4M9kWuOPnm6WZY8oAIXHAFgWHpQrXxiGVNuLNZxCc+z7H
1+XVAi1Q+hmIEj5pPAjg/fPDH5B24Ktm3LSMtXXQ82G9YmMZK1ovpVg38AwYpFYl
VFOQKYpPXztiZBLRQMZ16ZRUemvUzrhhC1ACXBuvx3IXdM5FrqfsbuFT71QbLQBg
b6XnYXCCJxmh3enOv0ovNZB198HlBBFj9egaXNkhIjyoiLerL/IlZD0A52DDuOwg
Tf7WH0IOc5QOsNK6cbovg//Lq6g2qe4vKOfkKOcum3709Q2Z14yP3GTpwuH3Du89
63yneudmZw20Kji8X2b6DRjMOl63PfHM9vtbshGbJvg=
`protect END_PROTECTED
