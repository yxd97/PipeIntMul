`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jsPxgzJnC6nZ5gB2Z9cE1b9z76NeixksUAtAjS/EpiEtDvFd8WtWBnONATatzFik
NQV26uW7H/03rV9PKZa41N4BXRcXBkaQnFtfKv2SzciuDnc4MhQN6TFnbmHDczew
P4feUIccs7Ddf2+7Bh40hYhujrRBgK4JMSbdRaI4i/N+mgNlAftJwTHGUzfd3oe4
YNMa9ZGdOU8D19EB4z5GxL7rHuaBpfUWCGVgZgRvwcUHDEFWrHeCHQapvNYvxCBi
zgDXeHr8aYwpgkyeKkKHvsZwLSGLFTZjoXNv9XE/0uWgi9EdC5yA9DHJseSyNoO9
HbD11GBk0MXpRTVv2WnHqEL/I34E1XuPEI+vIGcaHIyfBNcDaEJzuhNX5HgyvDA7
0WC+l8BMjavVDjcYq4TOfwqoJCh9MEj3q4+8CcxqvkZAWYA8CrH2hFdirGCH9AoT
By3HmXBLqgmKRbnGVx5odv6L3K/2hMnJidV6plZU6HFH7BwzO0k/RzaDWT9/jLq6
+YfxylJmtxK+iAE8MAqE0dfHHnEhNHMJdxqNdjbWU2N3CePwXN+RfdRGVEfFy98R
XHVb14CWlm99n/m9FavhMQ==
`protect END_PROTECTED
