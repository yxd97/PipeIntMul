`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6G9eR5+A1OBtBlFwWe4xh08SSSO/HD1AHbenmB0jizLMChhnvHe7niFO0HNsS+aG
KKJJd0jeq6Chf50EDEKV7eP1p5GAeSdO/oye+mGvO/9fLj1h9JhosDy0jZ/98A+D
xsw2X/TTzUFix7Ll8QnQlycb2b3ZdWH6K3p7Q+5ScYsvS8ZYmYKn07jvckJmQNkw
8PiemhaBMdELJeFz+/FYaCq9Tmbhljc7EmNSrlnTuoFqhOGm3MuWkTxwQ0ftgaPB
MsIdxw3Q7nxmwiC6GrhaVXq7j4TI4BHAM3WHhZJqUUEj1tuKtuO7ePb95UL5wpNU
hdaqkEmTCIUf7zQa0OmjXl4xu3uZ5TXPtCJjTkbnw/TGTv2uLM6/Ykk3qzaL7NZR
1bf4syThV32N70hgg6RItDV3RPhnJ7n1+10C3OGI4Ca5/wyVOclvbR/pOmD6wNjT
yQfSRgCnmMc6R3nMJcKeHO9hvEzNymJWPaBqkYFpvmu4A4hSS7E1VFnmVbHydbH2
hVBLuHzE5Svi1iH5n9+/5jkNHPOe+hGbdD+hM3HC9C2M6foCwRDS4o4v4ZWjkfYa
zDbHDJhdQq45Hw6lfOemUYWBRGAPT5S4sctmU9II3aEmVctieXZdETJiQCajlCxg
FQIGuW4O364ZynIGgX5RzWywzS2aUBJmUI3yf/fJNOUfhZHgpbOfWjZXrwTjzagy
S9IraTnS+jjxkMnclZAfoUVP8W0x7rjzPG9+zQkIm+H/x+aMcSqp2pLrdaxhd1pv
5XJvuBb3dUFo+3kqve3GIxZU2SooE9qW/8RdFJwxE+ZMoD4uXFM/a6LBi9mb+Qn/
ylfPVHKHOqkOh7ptov2IJHzM5uYgSYJUIz8gTE0lcr5okasbyF1/lbdVyYSCnF+z
Kh5l83PxAB+F3M1NaAFr2JXk4x9GIYHB1VLoCf0fONIp4vhhHmQrLCifvi3EWuI3
KHm0wtbFUMK5pKFojbNgxfkmqU2XepL4RwiynLulFTQq27h6eLoAWllgLZl3/cX5
hdeMh1tjM2F5UdskPj+iqy9lYcM4K2KPGDR3P85UQ5OePsB/1CwBpYn/IzsXlCe4
o5Zxqap3y+pxcruEi137+bT3A+zmz8mTJHGO4hntAgBglvTwqPXDiM8hGCilT910
TJnC5vC2gQkwuMiKhMzcpf37o0y7VgQRTUZZfBrg0o7HqV3mar3C2le91u2EnrxA
JhZDFNH69wwg4vWX4YQqMRhlCEjz3KqsrwZJTfKPKSm6w0UcVp5/0WsKFxwZ70LI
BxzxlgIHNJzEDwYHZ++uEM18JoZAfcfV/FWamH2hCkuL/xmr6RIyaW6gd2K/8Zte
B1y2w0LB5SJUvMAN6iOZYS9+edH8qd+nluhRzC8ZP8EJEEFX1LHF+Abk6y9gbYAJ
ny3StZ2F1uRLjGEThNLM3AXJTtNqPe6mb3CpLX0bFHCaH76PWSy+PhundX/jQ27R
mRrjUdWuTIV53gdVvZBh6bFPWyiqPe+S913QoO5LXx4vyJSnH5k5x4Re6iPqMfoQ
Opn1cesC3qg6qQxuzP1Q34f+HgeS0Gxj6CeGxhoYxJhfP2P+P5mJ2Tzt/cExARlE
P1blkz6SCL0xMOPsH96Nq/wQGTzgI+8UgAvVqpVlA2FGruj/iBNsQHJmmf01RdD5
pRmI5odxjaW2QllkzsPxVMD/rMsbBlgmtTLd9RVyvK+cp+PGW8sXCjO4uBpIli9U
OGdYcH1ogd7SyYKghfvFkk8zyXktfa0v1D9tTEQWXhpVL5dBugn6WzfIbBhEyYgo
sJAnpp6HEyodnnshTIaKNX1chXtoq4l/yV1CFE+OM5U2/2kabX2Qz8p2bTM2lo8W
1njTwIj+SPdS3Zb1Ahq1hqlVw2ms/ViUG4Bch0P0NRczwMmtag3ZaA7sAYB+ijGp
OE0PPGm8jp/J0Zisw82CKPQAQwecCbTc02Mm+zb/++CiIjfixk74i2t7DO353/4W
ZDc+3QVgFyJx3CIhi+zuL0X75ZBLrwVzGkmEQBjgXhWxMRYUBg19kEsH6By+MUBV
GjiQJi7F/HgeSs6pKj1KK+AmoBjKRYykcSukJuehatO0GtFIjq+F2h1wEBBBr9Bt
BYwMFbV3zDUVFKLTQbF02R6xsym3Q3w7fQv7nagkd97v11eEgPF5NNfrELwqxd3j
Dk6lfJhHueL7b4G8YYyYHYdsMcHz8KGvHpPtDiq8xCtNkFArmHOvP8GcMl8xNR1w
jzjaVbSKgBlJAnqwCODtUSxlcPwlrEtScS/kB2uYw+U=
`protect END_PROTECTED
