`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JD8/heAyqJnMEM6tP0qawRryqrFZCDwvSRZfsnJz+qa+Mu3antqBwvB6M9vBI0ck
H3WJJBX+bRGIVHNN6S5bAfi4hGubsVGOhtqZTPJOwbF7rp/ZeRXZIHrkEHeS21di
skURz/I9vUa3NWXh2gf4P3tMEzvAq6iH93wSgvnEijLgWDVj9bNMFMDrYT3gTE5e
vUkTMdXiEKBb4B2ZXM6GthYSrVzVRnIOqTsKebj0scAkJo3YS1afLWCKQHNsCYr3
jKyDn5t/G2JSPaKO3SJygEKNrNIt5M1oYUoi5QAJMD9SbLRutGphl9YdKOEBZQhK
u6jVgI0wxjBit6ylb+EIb0jY1DJIW62EzD3fowkjsHwoWitZEDbWaswzJmaOM81I
wB9E148ViX6TcQvha1omMV5Yodk6dUYVZRXgO/kzoFAu00tQPUCWKlYqhtI46NmO
uTu7FDodNm7008Dov4Dxs3fqPXrEvY5yVMAneDV3UQsuJZtJMUPFqPG9t4xupGWY
f/prSE0f9mmhQCKEIqoz6olhq+RQoJYD3WvKA4mTFF7yAKzLFrmPX4WJf0J3LHzE
jGTLD5+ekRI1XNVyeRrmgGoFd4BJhjceFggEoXQtHpSPQQkrR3kk7oB1Ep63vncR
/QN5ivJFM4se8uzH98P8O03KC3kJL3j83vDXoEK+F4oMV/Z+6aqoJz9OoZFS7HoK
u/RaTFV3ANA/MgAfaIHcH62ibeDjkopl9/ji7UgaeH7xcqevvo0I365+lXTNlBH3
uyQl43ra6YC9As7uOz7HyZ9gbUDRYgPGMBrNTXa/XGiyDT78vqAXyIMqcnMmpJIN
QlDO06b6Vr4M7ngyor5bGvBY0rOgzfBg0Am2NqZGOicM1RW0Vg5e91b9sR2jl7Uv
aOxHViZp/c2gcTe5re9udN0hxJAbvppHP9HdIE4W+i1cfelWkgrQscsbddylY3y9
UxraqTLemgdoNOmaSSMsvOz6j4WFQKfpIVS0/OH7k7jq5y3jrOwJb3xlt/Vy5HGM
bGMxM4t+CUfY1PxK/6Qw3efGu/ljKUljGQlnTx1JwjMPpPPXe1tiNSFNjHF/YE7Y
esdM4q51mGC/W5zd9VexFAfY/lTxtWMjqhO+Xu6p078USSIJcQ1kn4nAInXq/MFx
jDi3C9HulzW5gupizpJFWi2qMytgiskY8sqe0xiVCX7+a+q+oIR42/f9moHwUduS
6sRrWWUpNIglnh1uzSxfYZMgIQIwcJl/uln9qUyb1REbrwnNTao3iw0Ok393tFFN
IdAPw00ENgmuh1FZ2GFdfTRSy0kV3tXfiGxRwtwuqe0NLPfDZxmRHXAfLLegbo9e
gIwz23wl9UER+90miwhxVdPB+A2Hn9f7yE+g2l6SL+noy6t1G2HdV7YAxEdb9sU+
X4izyL9nEXr1N5Hd8fHXxdsLCJZlrsyY+a9kFWtdVGrAtCHZ7eHGZ6GoLrbQ8gPr
f/rbVjgocz4506v+VqKzBTEhsWgHbFGH08zZ0EPZKav9JUet4zXFnZeJ8JazUBop
j+i9WMufDEoWyTmu2ouol79sBibuwABFCfoBTNSrlGwiOd0Vlg8mvAi/QhLxgmdz
DwanhDhBqaMKceJwj7MqC9bjgVAb4cLwvcqHwdCOgWb0IEk8cWPVsEL/2rszjkfR
UKhS0R2CUuFp4YDLxEF1MWosPxKkNLLATBjjUjYpSzS7ilT6S+u0iH3ReTYL4gIJ
slYVUFJCLmp2GVRa/Z5MxX8NTTGnExx5qiDkVMTcG+MPOox8t9zYY/DUaVnUKKfL
ae4wzEb2EQkpxhI9ecXwCB5wcYzgtRwzCcLhggRhXSNw1Gnndcq/VXH/pTsMZaPc
NkNtqxmqw/r8sxsS6bboe31JpOLpjjOEaPNCBj48MGzRxgQMDhkqBc46eTOnST46
N6yj/4n19fzNhRYRoI9M7GevxPfrw5HAmdjJ4Wu9oMq3pHp5RJlDud2Uu3Gyjt8E
OuHQGd1qdHSB3t7bArQobLToiZbwMUQPxE1E0+/z18K6wu+Ddj/HQcWUEqcKs71F
4f9HuSqRpkCWRKvlyis7N40ZNNErU7UCkvdeVUsR5PRWbGVAtaWMpRZic8UDI+Xe
QfaIqUqY+h3RoPqJirxnV2yYwHuVeo9h5H2vWHiwLASZQmtXwUAE8aau7Un+7ebp
9FBlXrG4+D+N2TjaObinzC5z195qM5IztkSX3ILn9CJ6RT3C/5VXjqBP7cJwGoN2
UbppQR8zaTIkLjdCjJ2ra4UcXBE4wKbUYXFnX4V6Hz7Y5W/EMbvvv3NZt7b4gnwq
iDYRl7KHCHO3ArCE9sxDoa6fXhG2u/Vzncw/Tdnd/lPwBSP/ni/aQook+92hBWKO
zr19ZUaGuaGZmx0BQg2EIjcxyIX0NcuAdKpwWwVnR+LZ1yu2EO90sMc/eKRwdXPR
aXW6NLewVOvlxUKsJVNtKSLdAjyhDA5HscjDKa2DQeQekEitgbzogHZmdqhSUxPq
lQq1Pl7Wux5ax2NTZZKBuOLSTY45DxbFhLNFEuruFxkeeAR/HSZ63VUeM1pAkd1X
X0N2vWLGqDCwMuSMTw7yzLjPit4PTTRS6af/WYVZlsF9Dn+7mTsmwMsq6rWIh6eX
BSicAl0FdGHceZO7ZRL2nmh0cfF4TBTXdmFaenSixCRlAy0Bjgs6RUO955/dvl2u
+Q5rpXKxX15YkZ2g4W3LvrySdsWoeGk2DI5NCTDafB9CoO6pmxlI9e7sim3VIlex
fUuiPWFRiDJCdmAcyfqQKqHmsE+tnt16k+2rC/eXWndjr76CRmg5O2xiMtNXWs2b
UuUZelbZCW+IPnewjO2D4prg6czbXApnd0VfcSWdFxvZcMF3+MXgE8sYMgM4P4zL
jJGghe+IHiqDax3WQqpDVKU3ZUmG5K6kbkJ7gm/cb42JnRyM2D0TVSDDNIiinqr/
iEjCAXfWV1fdKHTiwEf5W0LOJIzVcCeHFUKMn+cS7o1eVRNmmTW+ENFXzIWabE+X
WKpg+x//Jv2DX+DugYSoh21/ctjS8t5rV6Hf3t/A8c74gIs6K7R83sBHwGzxXko/
NgIl7p3jkvYGZUegKwz+h4M/WleAJYd3KXDav3kWVo0NOgLHqBZDRvxsdRpT5Wrj
G0bGpaVwxvA7k0Oqy9Qau2nwXab96oB7pajzB79+6Yo3Z315QzFs4FuAybdlpLOb
x3An6R7qNZWiBMnaoGSDrA9Nwxm/6D5KcwV8ZSRczORyWFOPcTBnpjOS2sm3T9Dk
C7oTIRRWEiDf0JREGkMCDqamgQX6wlSLGy9tj49SoRKZBwdMBoNX/CZQe8qeNqt+
iOeUJ1CO5m5CPKLUjSPiKwNIkAioDfoFagCitjWr3uq1vSCbSPxcQCJnKODyS367
YZvyfQvh33OvUsbbi8sUuUpZxKjDNS+OT+WbkSALHQLKbOsp6hJlFon2GcEtxDHs
o6m+YLE6AbMnJeADgcDy9/5Q4WlB2HT4vmCJUmkc7BDhgefAs5LzyqwQ4n+0doyH
yuZ6GMSLLvP+rE1YNsTV9gRssENbgJjNmzG8eAbpGuf2LWXxZxXfFXp//6pBIl1R
STfDzqzSo9nlIsvvbmkDKEWxsSL2UPDk/0hfT+UGCHZKtJ/iB7DuH2zcIBy5E2tv
5Mf1q32f9wEmj5lJoaVVHEByRDeeSWsin0rrVQKVQGos0IiKJhoOwaXE9mThf9gJ
soT9SdRDXTp13bsw4FC0cb/5tyxC4PavJpKdhZrWLt+s889LSJWKubxTI/SeKGRw
Nlpp2AMtRrFO9NLvb14YK+95T3U5+HpdMIJ7MM87YQmhxTOB1x0wa8sVYOMzeAEf
uFMNk28YzqKXVivg6KcU2sVgFpnBrxNwz+1KdP1OXFwIePWOITmC4yDNvpfLXpiz
T4/swFDABzaS0ueosTFkKj3TRVVppBeBzigLux3qJ1nP6CsKWMnGGfwPbf4yH4Ev
8qbBzhrLHBrgrK1gTMKQgwhkO3chTWZUrSIyjGA5qlKyYgo6n7B0zTHHv+SSp4A7
v4BDbu8nKl7NHAvTqJI4yiWucE5H+QNh+M4+MBqwDm4ZkfvKJZC/zFfftnDd8RDB
7jNXAZKJ44qUi5qwWB+5TsZp9OxhrBuAU3/UMBkdKojN3gXhVAYCV16yVElCCLZ4
W/mPzv7VCgnHqXQoySijqgTMJyBxKBamSTsCYv1E7QhJbluAZ1CLHY7Xik37U2a5
8al7VQIBhypkViABp1VYTIkDzMrfjGAY0W1+EmSp64Uw/gVd4zcGfxMukL/bJ1/I
kdSqcjbx2GVgxB9ho/iWk2KnsIPsLM2m4vOwSLXsjXR3on8u71zO1gKbTz0OyDl9
X37PeXDEKEk4ITokJU2zboWy/bcXhbYt6Y4ujeAsvhB1SkX8sRQwVZcmGi2ouOBb
rRToesRKDm5RBD2jhNHNwjAxNYlJdMu/svoRlxxB+fys7GfIQomo2Z7iZ34Prf0L
UaUpkYw+UbbAjHBOvZiMbfDILzYUFgRu2bJ6BvF89NMR7jK6flgvb2WWitgC2tVC
YAGT6A+eloDkxIIwIqkw7iYF/ZcmnYOwuCNl/gpx0Bown9ua27fSdj77rP6zQkXg
/0S+W4WsACmkA9Rx+/9cE9ZkTH7NBToZ5zLEsYIZHsqt61gbGQ4nGdLbbfrWGJKm
Fk1u0QfH9w8ie/i8vsI9bExySVot83VWECBXGDzH4aEBTSGY+JzDgHZsyiTP6Dab
Mu72tItNZTB+SLzQMD0ZlKHiEKkT2oz8j9SDvus9kzjuIzDu7lJWV3jwZSpY6ss4
xtzl586dtmzYD9PCPJmFdmj6cvsvU0ypZbUYamr+JxigcjA/EKMB1hhDMG0Ir5P1
BEHyCrnUa6QH72PRDlqRHsfMeMgFs9SYMa0iDXozKv+Ity/27E2dM0RfsvIwLHOl
bnaclFS436fDNp93Wjv0h0lllf5FKlhOcg/H4FlgFkjoQsWV+BBP67pjxRwI1y0r
FtREkqzF4cWOVZdwLWcrC0PaUrk5QbnUpicoyQ09oyXkqSSq9Re/sbJ/0ccEQKh8
Cu29trOeWK2r3yroGNeHrv/09kFWEqZVUZMLJeN9QGA1X4kiIMiWE683WCC3z2dx
VMuEjy7LhM9NkdnlFCtOGFn7FKAPbd5ePcVE+U25EVm/GvRkt/UATR99tIhi0k92
fnOhE1Qj/SQo96/AZbuILBQWplQHAIH9yTT5iqqiijWPR679SsEwH2MGDOu9mVsg
fGtoqi52GFz61+jIafZWSWmtjR9lUVyo2/vkLKSpOEJJHXeKdPeb7CH+cTdeSgOY
bi29b8Zzugz8lPge8KZIOsIwc7L0ihHGcjAKyW7DEkjyuPokv4fSEq1KoFgwpRfQ
d0L52SSeYNDJhPCbxeBh9he0m4Ds9TPJmGSiVUVwZ7lucnum0/JniGHHBKA339rv
cu3hyWOSY8stcnfZdBCm+duRRBa8fzrBadnBuWeH2n/NtnyjrS+cVBQ2wbhbtASX
nPYro0sDzVYqgF4V9BFLCS9cP/6LzKw5SeAUoun+bQTQPY4gJNS2cyyih9ggShhf
NQsmQg6jQ6SQ8i1nuJc4BUDJKXfQvhaYbX4geoLFU2HkVB9ZAiqie9cQjCIPWeGK
XOHPhAX89kJr7sb8eV1Dm3RGQtrwe8M8+hB0cupamdzvQ/zar7shPq36CnIHqLF2
98PVkoWGEod/2VJUoorSeM6a87snO6BF8n561Cw0KjXemq6Nd2a9LLPN26Ri63gd
WXqFfzUbK1CCkL47aO9FE+KDEvEzzGiJRNg9F/9oRNeyo3h557euLp3yv1JRj4Ib
5FgTavOCcBBWBBBkAtjZ8PMFWoxZtvalYIsVqdpIoCIaRf5D849s4lSOpTz6i6bO
T3+Pp41qKQP6VND/eC2xWgbZBqWC6Sw55HPBuey9AhfBlzk1c2MMtxanQjCNc2Wn
MmxhXBIdPiIuX0XVs+rAygKKmHcq5+2fBYyvy0pXCxipLebbqlzeVSq67ScKmBbh
yKlqNWQLBqgnZP9564Njo5ZJf1D621S5d6iJPul1GgDny6Ju4z5WR8hWHmaah6VI
1YcWliypv09dag54bKXLusI3RxsaMxd+X9KkRjGCjswWKdgoUEEQyMmMAi/zq/pN
bMG4qSkCX/rx8025AIQCwIjWbWVdlHremjVo1QSzzJTFR0MxJQRwbxyiek8hlSPr
afUo1jdhfPMog3Rp9eTxVRbZhZ9gH/yosrOstt2HZOGVutSxgvklg55UJY1DWjGs
EnNf5ovqgACM+5CHtXRoNUH49DjLvgHHGRISrJJQOBxAb1qrAn51Lz2v6TvWctmt
xikdXUyVbkrk9TlLdWpyAYI/9D4fw6sDMoIum3ypfs/6IsKE0TDAJnG9Kq7zoxVh
LqNZulSAEVFmDEo5GsALI0cmW4XNvdte26hSiV5eRMunYVXzrsDVcZF79iNwcoYZ
MVQtMjUZOJs7BpfsTdtKXN+IdW7bbivt9Y9UZuBP2qdTscxtfxth907SmdAkPvc3
RaI1vLC2O54xZFxEoT70P5EhI2XBt2/YxKKTkQH+ILHsTFr4wtgILOKERFbIFVEC
EcycagDzYiPr9AJ//ECsRQiOjtTXJ1sEfTg0r/hEKewB7yAo3G0rPrBfZrGAV5kG
IWXVYMoz3LTZj7W1BPtu87Iv3NnPJk3yrLihinr0z/qr2h/EJZy5Qr5msxXNHGXE
ogNM4zoY1KwbQaOHaZ5nI2I4IyJNGqlGxvpb+rRmQk4bfH4ZYHkpBQzZdMJaihRz
kskn5x0+XtU5+M7LFVRgWQZsk4vjjcpLmuzXeNypJa+apytD11XZppvgttDIadNr
SfSm+qcKeIZ34vaGHoTj4EIj7wQ0SxzPhxMiz9CWuKPqC0JOgB9/HN+RlbDyPSHc
YqvRr4agxftTzhjsf3l9zD1IuMegiQZgn7K3ZFXPot/JaKWTH0fCph33+WNDXYbX
qSPEGN9umFi0T3n8MnltMU0E9xXeRPV1UMTXQzlMoTuiT7D5sF47lVGLFxfw0gcg
lGrlyF1PFmtB0mNhFFGIY6skvXmnZFGJzV2REaO+ZzkMC46QoSX8pSPBMPDEkCjc
W6QiBAOni+EwgvamafEVsS49VgY8YK65v6nQpU5HTb29bvQPzNsqCS48L4SEwWYD
FklexTqglJdQEPp5GPXvh/AUw59P3CpB8qsybnceQKhClu59hIYaEraL87lt6rQN
NfzEofJNNZ6OI+kEWLcUkUJJm9vGpTGdh0+1WZ9Ld8/Nde+a7/QKJOVbO01CZlxp
pGjIajhfDUCU3b2kEAfzhUOeBSE81/H3fdODHeOffsrh3hntRdAr33IL0NB1l7eM
iGi19uEnAwbb4DmmXdpkghQwxD2796UNtk9JKGtlPPMP45o3bbqMxThoY2RfXukA
tgcptfT4S/1wwWhStOLhE+SZ4Y8uK7KcujM1gVZi3weq+uU5TlGJttYZx/Yf1lNu
W0+dZie9fxOhtS+QsoixRG8erW1YB2mT6RXQB3LcdAAFuyD2jnmURqKhQ9jA8brJ
Yca/kRCUCSO0RNrz0cA7jXmTHxRlV4x+jcHQfr5AAi92nMMorkMYwCUnyOsn66Du
7C9MkfIVlYaMvcpxAyffMgqHEB+hGB2n/nWUmXYVd8xAu5he7MTGhh6bvdlXW4nK
aZhb0iFnySGuaqxFRNUA8+n6MlTPHbUiO5QUJHE397VO0JroCBQM+W/8SMHekXkL
aeVSEMLz0/0HMaW+3NRML4PwxMDNmEhZhmKhB+fAEW4xswzTlIvdNllzBCoRiT9x
h4IKGH1b2yy6GFh85ybQRP2JDlZfrMvDlkVSpuQBKRANYhSNhMAlxA17pvaOIVtO
pXg+Znbj6mq2GJMktphkF2Ypch3Twkgfce62elylEVWocoqYXDfJiJfameTgz1Mw
IjVZtOlMhjqyrXoMUPx4+wMkmvvWjjojOoXyCPQhlzcCftChKJuRgGNVRFCAb0ZX
ugA70iPrlPDKPzlePKJq9IrUoaj7XU4puomB7RgiXJGqlQUMIavJXGiQ1Sx4CvEP
EloWtpSdCNUaOFxUJjVTdrJtOgOIXeQxjjENVrJNcUegO96r8S0vTgG41S2V8egD
m8e+ShrdrQnKWfr5z3F5vgBbLAa6Wx0bYHqWgzMaimlIGPxFtGSjvUq5dWkHqXXm
pnbY+soJkSOIyREaz/uFFR/CxHLHiPp9x8BwAhpryr9x42kCDBAY8dl8x5+TazRl
hWOIU6aYRIqQgxI8heHatdF5nXL6T3acG+NTz6qaapG0s301BoL6+fxBVfJfuscA
29wmn01dCJfVBodCz7eR/ILA1q/2y/IQLPAumthFitdH6AgldFkdt9BqGPBrm2Rm
f7qYe651GcgjH/0TMTW96OfNM1BAsYmUBtnnQ5oHLHXm3ECVLrz3s+TgPfUkSR5K
gR0tj9YDfHpUhPsgMt9RG7wnnObi6/Ia4EAO50bXN1HlAK7gmiQFUMfy+3029WrI
uPFe4maKp9tresgaBjDPoiP8zp98LTCFP7ee2beq485pJD2BU1+U541IA12aZ4CT
PryLqK85t7n9dT+9jLZI3/7DKvXSTEJO2/r8Pk7TOaR/m0xxHucnAaFt/f8KwiiW
bGk0jKFsvBcveM3H/WF5vLSTwUlRhHObRsytdTEou+G7cMWmcaX5MdXKt+BVONAA
lBpwous1PUPzhX5dRCYiSzDbxfxbU+8ut4ll49lHxQvoDhqdRvcTRuZqHGaHPZp3
RNvz9Lyc/xriGEOkvel32X7tBAac9FFRYJbiO/xOC42WQ5i0qme4rW+dex5HbOaQ
7nTpat3K0+Vq1DmVVnGvhR+DH/W1hcGe31TS6E2VSureqFVp0Zf2aJJvmWO1ANQu
d+IsBJn5n97NftQfXzXeMxX4Wmn8vOvoqJZI/f+1kUHOjHePrdktaWVF72yKdgcs
BPn94jdK44PjYVDkAUlcphmlwxL9zNioB7dvWWLBrtA+jGw7gmTIHtwh0kRHvURN
ZrW3CWr7NRnEyyF2isIyXTTeqZltYHPUOar78w+vZg+rXUfaP9XuFW9LwjzbzKYx
sK7T6mXuYs3/LReMbuMazF9+YcX4siSlEONlxtvBs4ghFLPRUZzypup0kg/kvyh3
xyKJ4hm8ZAiXZEiUk/VCh+m93I9xRASzB+Fq0o+3sne46G9hS7m6Yq/XWO2P9CD8
FB62dXpp1Yjm6k4+0Npoxw==
`protect END_PROTECTED
