`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7tGJlJ9j++EZUJOzC02NIlrl8ffaKI3XVrCog7K6d45Z3vyoceVpIzBi+SQtBcWh
6FzAGNmdV/Ivk38+gLjjQvxscbsla5RuqTPyYhBEt+ZXhRE5JwDSf3xI66gNzUEv
vFftmk/xsjTAu1rDmPIKy4nCzShYoosphfZ91pO4YW8hR1VUz/kTnYaUrxAEpBaQ
1Rtho4FC/2JkMcj4CVZUciJ5/lPymn1eERPVCm+GTO9g6LE3K0vwMMCDKn9VZnK2
LDPV25TJGJCE+DpmUtymJlkTiqEYer63FexwZfWtx9V/G0qrNQhAcMEp0TXxbKTA
XUP5SbqgbBP61pPX8panX8hh9VnFuYDueZLSyMUEl4QEwaNSeDifVj9NZZExrsdq
65wVkyrSpOcZU+981C3B9FxNJ1DW5cKszdDKbDYVBqUL4COW85G3yxQ5pehloLka
mVkyyIU7kxqXuKinogOCmfcggSJtZUc5ZgvuBMGl8wr15e/lU/vfeWu1uGbpOvpg
0fqtnU9yurnV168byB/2hC9HP4ki58u0mHhhvT95KEnEQ8pqJ9eKTJlEnGtNf3ri
BR4puD8FB4NUNEfTs2HJG1MEVxjxSZO2ad49bRe9uQQetVACxN5T3h4/l/UFXam/
k4+KwtYZ48fwsqg3HKptRS90Av+bU0AkCtxlF6mTO8fhvPdmtKSrtsk4eTP0LQRr
0jj7p2BzsfePIHJC+h2VJBVVeOTTWSFVRGUDiRzd14Qmige2HjyUSovnclyrmmn3
YZhyaNU7U5IoM/klXcMhyS2ilMMDbhnn6q1BdPE1ARVyhLoCnwo2Ubim5Qg4mpQf
/6pyHXo+PnSGbIkyfNAsz2wZEPAz1zKo3WRE+OcACeE/JqM8znzKZVpGQ2z2cnPx
M6/HJpscUOdky/ohQWU98jhaNV0mh8CkOk0lfmO0gR1T2TAinW6M0HRMkI3Auxr7
hiqKwFqJcvUzXVpHiL22rXT/Dk6DlXI0JfJbmZBqx36QclW5c8wOlwBI45H0R8lc
YkfDtx/FXYX1psrbeqAfKI7JYHIe6k0Cftz91HXyYn+xZHQmb8h9ESrO6q4j3JHC
wuJueZ2s+hoHs337Zpj285s0CxlocR3w/Pxbk9eKdPQjYWPoF2PVX/8L3HcFpKMm
OKBbdKZZSWLIlJyOzfsy2QW7bEucsT8LCMIP1OzRnMcRMeQDk1GJSlE4msvLM0aj
aVILB/df+oM41pMIGtQjpjHPNJQdxDf5jRY6Vtcg3k+nlbXmfCy7ycPpBtv8nLmF
WbmC00y4/ioZHIn7Eu+r0TJ0wf0xdso8FhjH849sBYJbusoosmE377ZD0FDa4t7N
nvZxjPVA10sW4NjS+kQBhKQrPb/+1dGk8wS/HCM5R/3T6E+D+TCGJdU33j/n9g6n
/pLNnizEP4s+VZd6cIHtwPnQgTf7QhuoWW8nFy6IniqqBLLRnkX8w6zfEjhd0qJZ
2bWlFPDgpuKopm/tYnxGbnI3JmdQcezGbVVCXxrc3avjA1uvEEYTUntmthAsmrAo
9Aq9QBnvfbh7M+qDOSO+WOmqnRbgaQ7irzMKpeq61xGLWQHIj4AXhWnabqZnz0C6
dcPjdnwQVLAEMdkXMQoQCGgZZjvdf1INDor8IHVFWjcfwY4ftZOzDxP+Fvuex9fa
yF/7jcq6M+5xp6vfS78bODQu7X8YDsIT9BOBnoFnNf7MjzMTnrfRMYL8oaYslzeZ
V1W/azF6uT38je85+Hx1kWu793EQKdkyojN6f+tcxIaZLcvBjzXAdBtTEDbcrimq
zqcgzAipdHPu63UBw7HXF5d+x+L+cyeUBb1raOE1lyQ/1qpST4Q2J8oXAe/rWmmD
CAs6M2q5/p01pzznjQTTI2WHbCTSZtzFJOIWAa87lqQSoRXkfM6rdNCfuKxxEmjg
wlwAZPtFHgNOFdauXFrJFUMCq4GallsruUb3KK8uENb296IVrcpHa1LL1K3XGrHm
h+7AyKWK5neeuEMFQCaIKcR50A9vxMOu4JgwuhKZTZmsS3VWphjiXIvUzXxSzItr
OTfehaHyGvz4RF4dgTedBBMzX7HhWsqXrSma67bKbChDyegf4TxCQ5U5kWqxHZOv
rpIM3Otb4YsvqQOrahcaDEzsFJw2hZdaje8KvpDcL4+euxoc6QHr/j57U944/+wj
8jV2q/lqjo7RTT0p57k7TATmv7S1+rUhJp5DRiDleK/tt82cThm9LxmF7nKX4PqQ
sLWCpmLGBSSDWg/P7C2stZgJHuC9D4dNPlHjSzCPFprwPBEuLgWymLIdwIVZPnMc
hx4VhBh5Q575jj3hgxgtDvoNHPf3u7nVhkLNSFSlnJSDWW0PvJEXKaEXCWTaREXj
dIjMshW3gPJo10SXnLtGCX4F32BivwkIxtrb780gLT1n6MDZ5PXcNPQlOnJDs0tu
gfcIPhjJiqYdFZxxD08Ig2GyWS7fUX1f2Q651lf2E0k3kw0Rmgv60yNGkF6lmgls
8N7Bhk1Uuz35r7kxM8JLmKF6VNTWRfdgCJyJQAxLGOL2A0Eb7Mfp+0PCaX8z3WbD
03iDs61c/Ifrv+lFs6VyImA9DpqjRJ+gSDLa/AjG7qRkAhls0UHAw+Qx5PA3gsWX
vgbrzCjeeSs7Hj/gACXkXNgsb9KBOxrnX0CayWZBxhq238TJdXZ3oOieJaYP7JHw
BNO9EmhIflyY0e0SNGdNQp8LYkbiaJRzWzdv1BXKvLt5WgaQdjeDEyAKza4j5w+o
QSDN7FnlT3JZmLNqt3e1atfhqytvXChnKic3G7UlTyXEoNXmNI9zzz6RJkfjxQ+G
Eh2B2EUmiJNgIRRDXfCie1K5M76qyoHwoSca21NbVD8ur+Rynby5RXtLEvNejQ2F
tRBU3aS22p7eRuaBylPePFR1vv8Yq31/E34hyWnJ4LCfNgHRE2WpU3aHVg0vnjkJ
MEBUBK6QrWV/ZpNS6uO+aVUKNFw2qZDwOgSRziEcQ9ae15m80ITeVXPpRI31tvta
RDoabu549dFVOkI1GwaBlFnyhucAlGxq0WPD0cZkBKIXaeVQEczIbXT6rEREDrxq
gauzMdy3AMDoogO62IXlCi5WI3bRUWHigJRa1T/p8sBFiUQlny2hPEOxXfUYmfrb
h7xH6ZZ+sUatiz+ozp08rWMYfYhW+rnWw4oNA9N40ZXzVhmHNbzlN+2/gPAvnWQm
+2oWSg+E9aTqY0cqzKrUVuzjnSPXAqkZNtH8EhYQP5yenkbxwOEL8EmxMqB2Ec0d
OlAWX2GRSdmWavyLwARBq6+p9dpJFJ/ZK1wQ4l102iXXBMqH+Otxop/IDhAi5XF1
bQMdQ/WwAODy5h8ZH6ywmEpiWlc07izvZnkBoTZ1AjaTujmvY5SNcBpdMTGzHGYe
V5pm4EkD/3sl/tqjpF4U5pW9z8l/h8syyYs3kOURgUVCcvgzhxbgvspnmZ8Gqap+
Z+8MrR0N4PZp7rKZHWastl+WCDM/Y377yauC98fIgiO5wx3WRBpuUgHTssDYOGPU
pcD//DnZrg2r97FEjtJZWubgIpvTPLFnk9WI5crmvHVOhXVplqD+lhBZ5FiOK2FE
Zz8qTv9VDTylFj35yMEXtbKCTVhcl1nlUoIRssqCTyqh99i0R+TgU3kdKGU97SqH
EIDCppXwF6fmgRUn0ASztyvz03OI7TMQQ17oqQ4eAADNq/Qju/1zT5jkBw/5kZsC
PaZYAIfRoNrFLEvOkAAc0bqvb0f2JFPBfOmRsaOVu7w2wI91h0S4WZNbLNG+T3DW
zNa/KRyDMB645LVtdafjxUZOiI9FXvBrbW+aHi/rHvJxgnvOwJLwKwPzCr0yOKyN
OMLSS4pnfUT8ansj7+SdrjOME38Omz3bP8FvjVBzXNZiG8d1WI1olb1BObctYA/G
xyiPFgYij7t3e/+sPwcMgA3pnZzTucx2/KyFfDjJdAY+GHFj6aNSJkO0IWzpTo2c
E9RLyUEu8jKt0Ff2rjn7tfGwi0XYj6BCMd15YaztcuZ0IJNQnmfNQcHNaMTuMTNB
AB7y48qcAOaeoLdSWIp/VhNVX8LlBelE5nzdSmYvrd123/4+pGLTjqyOknzUdwRU
fxdc5vX1kAcrM3p/pQe7mFINhbocSZZ5tP6X5quyccd0NqpdOL1T0/d0TPthS/sw
vm/wB6xLpOO116duhaSopkAVbPZAXrgVfxbDbLPNsa7QkXbA4avHn5jXRmYFdMhN
IU8hZsMhb7YBiGZD60V7Ho1ZxgRRb89dvq5RU1kuoRKwC1TNcqAip1xXQDKiO1p9
jPr6eN81r55Lq/+/yRgkvq51GdO/rFChiW1g3YTgPtMvliNvRqARsZuYvLg+bZAx
otREi2aKSmuBvXEJUVapw9pONax93sleNT5F8ApFYO4=
`protect END_PROTECTED
