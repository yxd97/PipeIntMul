`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Ah4wOI1jpkst9Ezw/oRwF/eBDFnKCO1hXSu8naG0gdbWrqX1dL0j1OKGSw7qY9g
btLesAvfSyIlks4lyKqDPykOJo1cLSNYNVwgTMotC2AEg74nbHvSvYfoXr5DjHkm
aqvycacClhG9ngbpBIa6gcbSTF8Tzyn8R5Mimk3lDYonqvlcdF+mxIy7OWYHWLSf
hxBMtCqMt5fv9q2+WOxOoc9a5XlKfHC8D10scpoqPlCuBbeWTLfIS6d1WslNA1ET
Z7npxiYo0tL1zwZAJJ5Fzw==
`protect END_PROTECTED
