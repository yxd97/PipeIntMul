`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fbcHHNjBwSgs+mT68MhsEk3Gb7ym2akkn0ti5B7BHw5qG690ZRuygZtcb2/nIsQ9
Vc4v4NTkfdLRpil9ehjk+a2eGG7D5une3KoWXBHP2Jft/SBdPg4kIrz86YD9Hzh2
nFG+iRuFombUZxLTor8+5MLHwWfCxVtNaWOY2SdALLe1Eg0A9Ur6VNEuLZO9K5Sd
ghmbZUEkHPLAz+veG/Yhm1cXPf9pU0MxhUOxEEe2k+5+FRqVOKwaMF0DMxs+LdZ3
V+ixOTOUounsJWCBNhhYn27llL7m34yIOc2f3DhlhwpP+VGUFiPb7ceiK1fJeX5A
/ZGkMbKG4frqe11SwsOu2Y7S+LdRdadRMDURZumr/ZNKl5XZK9CgCCqB9OcgAb/M
De85gkRYOBeDoNuKif0MpMsvt/8Ftc//zF5AON+47m8SVGN7c7aXC19kZJck+5sA
t4lZpYZoXu4hhjZIOjRACGIIf51JTue5ahhO0gHovAqPM4ed0RIzowt4nkLJtb+W
KOvA5LnDa2g4f9tL2fZHvpv+BVbOX9u7v3sxAENWC+bEGj0Hxz7CqJsfDfNzPznm
XztZv30+Lbr9xMPdXmnsPQ==
`protect END_PROTECTED
