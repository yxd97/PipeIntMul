`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zGwookOkRfHUDpYKw+i7wDGG6ca1MEdpYU4RlWEf8RzNXyD1DOVfmzhlTEB9qgOM
jr2yo5/51vEWrGyNOouXTbvmfNfWrtd2lkufD4fWNUOuIqAVGL5FcJAMknrXFicT
rlJq9f3M8f9lx8Un+qouKqsbRIvoJDuLIP1dMF6x6LHFuYmtqJA20UDYSmhE9aRr
DwQYzRek2+8NB8Takg5z+M20Qhfh0EjyCEiyCsJAv0cyngqKivvN9A7EzikPg++P
YM8TLZIgTgarHNC9uUUZ7mLEJ01TWDELdtMm+2PFMlmuKrAue6pk7jdVblQZSYn9
oShEGwZVX0q7Br/rKj8Osc9W2w5w87N7QGu1JpvQ9a7Cx3hAqt54OOnV6v5kZ/G2
lDLE1+7i5HxHD2l4EUVVpNVqCoNayZXcgtfPD0XAYTbAa9rmTHNJ4eX8HS5+LGdA
RYPzKXgHf5c92U9bIAVrcoxJVSV5JDOcw42qkyoU0Cq5ENU6Fjagb3bNa/o1vAnC
dYWzeg1pJlKH9rRTV+n7VCgTjCLbCXRuW5QXIRKWuqB4iaVk2vScj1+EXmCxcMrn
tNRg3C0klJBTtbgISEjvcsPIyp+QLnhPQj3oIuqGQRppaxmQ5+GvInoAgR4kj+75
pPHN1KeiqQ0UEtXX24tXziYzWLAvUINPhTC+XIBZd1BuueLispNoS9afdO7zB6yf
S5iE8ACs/9ZSde6kNP3UVdEVz0pT2H/+gwh1ADvwRqoIQsTscaBZst71AXnWJGgF
XVZMIkF7ufDqd0eHG58SDmi7cqXadCI5BX2/M58vT0NlicceP7DEc6stmhad6kdg
RA2wMX8acH5uJHxWZPCW8Lze2PiyQZKbChM5Ncrbx6T5eGrATA5152zDBZ898xMg
JgKlkNGHDLVlbonC2ffeIeLKTGhiQ2scBV3KnEbncGA8K6YLQLPJJJQqpq5NCYNy
`protect END_PROTECTED
