`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkTNoYRM6q2Ji5PyOAQta1/SHbRIlaOd9LtYZHLS/5IEyziessjDL1/WrkRBYkQJ
LcNpAD1WThXmAkTJ+b5W2/mdittBe7jLAnzvp1/cp1B8t/E0yUJ6s/jqZ47m80rt
IQhxpzykCZPa3YtLPl/Jqm68bZL4EQ2sTgrYhk5+6y5+jzpMnhPKjBAap8W6lIg+
FFSlVxNwh43o5WUXV50uW7kbGqwcQV9MbchdOfbpQrEaqEflffm8NnE/skq7PeH0
UxXHAcmMjD/lzwbbn3ZH5swwd4qPDpbDqy1oiU6BrbeEOMENH8RR9zDZqk95+28h
uQ0Rx60vwEYrmu7dWxF4ih7AI/JjDAEqpwSCqlspHiP7A/vg8dQCwFt9xpnpsGZd
dvgNFBJq79XGdil119FaprvT+nXfl0VDRcB43Azgz0zXPH0DqT8qXWpPH/5ibNhy
aHBeKBmldWXdUODInf4F1Tww5EIAOCPerGQ4cubkc/Enr4i2DIrghfv2+2N80Oc2
DFxUiIBbV2mSvVUVvqzLQigTWabhKIMdP/dfHwBsgdA3OhykyRkikT+7CSKYBu5C
CfSUs4ezlaoADKTAagKjAHQI0v8g1oastzP+Uo1UrsNdcNAXRe86fZG8HjHElPsn
cJQzwE0Qk1qZRxGYVFUjgE4csDJoBR6ZTm0ms8e5nW3NqMbgm3nv3IxhCk9HLlFb
ykrdM1s8wEPvdAUJbn3I1OawluIDxa9OtXejcGae2kIFANh7eQaWoX2zkmmkx5zt
GdO83BJsbYXKGn6iEKD7z11qtbp6FNfzCX/FZTEXJ3egWl1eNSyzE6/mKo2Fyx8W
WtCSuiDKxIB8KoID+HB1Crz6o7Qwj4ZFJAbjn/q31YmAZ97ShpePIGFLm/mbAKnv
E8iw9Wp596b/3wtQm8DjLo8ynzQB0vbAsLedJVMeZHuK0o1k9IYmn++meY0a4eFF
g7kxOWvn3e9cwRZPdqHDAcy9JauOS1bG9jkFE9OkEEYIIdF9nEm5lEjneAEKsvbm
xx1n+lk9U9d8D81t4m9eblw53fO1oOIg5lOfoyuI1h5A3oyH+hS7KoBR3xwJilrX
EzsrnqRv5kesTqN0m35puAZvngxRbbc3mm947vvmJLtoqeVCP+1nDdg2Etv4npue
yDL/Zj8Ktg9auwot2rFsGsbLOHR4ZP1qjWKFrEvYXzGTeEQrWE2hjhHFiqcLneeC
27800yuc+q+Gy6JkbI51tHemHIkMJ26+3E2tgrhc7Dy7gc7zj6lfa2kpT9fzAU9Y
++NjJoDwuz0ZoTi+FKnyf+Jn3wZOLkivsYHmm6lZosR6ajSfVyxLYotlqsYlh4tt
Ox90SEFMNuysc4xNrmi8w5Efe30Na8jT2W64ju07MxtDDVz3qnD+H/ZvpnlqSH7O
h0pvDBE0dz7/jK0K6EwZje/IxrZ20MyQENi/KWN32oTNQaj14J3dkQNMBX9H9+57
vlZAe6o0Vn7AjGxfpkk9z0vClXQ+q47QaxDgrCdfWcxUI+ZP9rmMAK2qIuHNUnPu
c8mRyQ8C+cup4NxO9VKjMH+kEZyGPOn7Qb1xa4DQ0+RTOOqgmrliTyZVXpqhpXxW
ylhVKHvNzc0PCls2QuIqtQC12iZ3ehWABrVyM5oCoSSznNBkg9V3Ni8PwDF5LZVP
KuIjF4OROhI8JZiNg5gOf71rFpHJYCYdWquPkXs2PtKaCLFLZMxkwyRNLSagyAba
NH2BcSaq+C22D1tRVlLx4w==
`protect END_PROTECTED
