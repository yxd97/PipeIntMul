`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EY6yzOvQt8ppisx8wm/CM0dcmD9LOTojahlCXqYW+vv4oCX3F2wuniE2n6DaTUME
6TZZY4gRdDt5miQPH1h3frAzpD2pqWnPv8NXdHMZ8/jf2rjNJRRW9p5g5MLJyur7
zEH5wpkPL8pTTnNI7tOqeRL3PAEupBe4RRDb+CQVg9LeTWZOBu0bwHELhmNut2nI
Sco9DDzlXJ935sIDUKh28csygc3K9nEJTW1wSekg9lc/71JdZ7YcgKLqS8srBSOk
rj5OcVR0sP150rn7S2YLWHGFyAz6bGSr4oVGgjWoGFfJzsdbL2AyEMp1ipXznBl+
Jf/yhsv3Vftm8M8tVEOCncooYlDhUSTcqKX+YtUREApcaMPUXBABlG9AyYlj2bom
IuX24MhU9ozeb10bXYT/B57vxSmhGcN5fJvP/s7K409ZCxLiWwEWOGx7u9/mB71E
TNUqTHpwqSfBFa0IajQ+qsWQpmnNuVxzknCSfW7lkDtq0dFnHG2mPEZoFWD258Vm
J6EFap/2ZqaKm28iovqDWFbYFNb+b1cwk/bQrZuG0JF81T2tSicpz51MlX6cyGGm
C3jFd8JqNbbreibPisF7hYMi0uhU1lRwU57ndTSd/+x5aENRuuwhMFcz0M4+6vaI
OagfxwebiXIqkeHLhwk2ag8RqzEPA5MMWMhKL8s2/QoG8fYAnCDxoqHc1BQJMN5p
8pemEOYnsdfuodTORiMDXmn175GIoIH096LZ0/JF3NH+PsNs3+Z5TOuG5FAh2MqH
VazUnHUisICWVo++zbDvzsonV7eBSS3PHIuLHmRQSAUPePAyREw6mUC3CVd5+F9S
cvjmYeMdJ27DDtTzLsTLSspg7Mt4j8sR1wr+zeasXCLnT2qwu56J6jm4Mzrzr3RI
6Wf2U25lIRnNdG8bFadOYfS29d2A/myawVGll0suGA71GSeh+i+oTNMObb5XInWl
UMVK1Tb67ypGmDL/kv2FirY2+DLKAWZ1s0UrFIJ2HeQvIzxUElXyQ3/M5QZMgol+
nIwbcUW2IOsmHXmfzzyFaNjNDq1JMDMtZvQ2XCGOiImWT2JNh1cZH1g0Kw3wRPuT
MM4S7PCMGZn5odPbaO11CcoSvmuMn3ltn37kO53qGrZ4XUfBZrY/iGBxn0LVjU2L
P2/li54FIZGd2S8HZjvBG3R/k5gQwsOOvR8odVXShLx7Lpnys7FpCp652o27MTwP
3G7iTeXjGdSfDB56pUuxhuTUqvmcox1Hkgijv7zQ25jsiqQDDEKyA/sUsOpnfeKa
ZhUERTXdvziwhu/sQpdRojKei3pynDumt7vQacD5bBz7My5DQCHxwaxOIE/9uuk7
4o80DR7Lp2ds5xSQeSpSv0MSvPSFi5SAayJmyARjiIkFAJ/JbDpScReDryNzmGom
K0vJrpWGRn9eOU/mszOcaAKPaHFyt02l919gaYlcuBxdLd017IqyRMT89x77v2ee
d2MsVNnMwiP7dJyDGgQxaYnOtJoPvIft1WH7kAO7ISDrk3JSzQ0eh0v5cRBVm78F
AT7Lo81yWFwakZcuxjqzYRTI7lyJdEunVdf8mkFEyChlfK1TguVhntn7v3azdgtz
2o+BVpe+wQwlpTn5MbCoY/Dw6En+J3SYfbAcA5gzVsUC+/CYujjHIPCYrWCXAK3Y
F5yAJSVacOHucQwws86TG+uktYLWb5kREu6khACBrTjiGoTXhZcb6A9vUjdw3/TQ
JYzy54Qloob/yyjSHFDetuYdEgp2Gm1f7Q5kASJQ5G61KNUQj2Qt7pIqi3xMnofN
FoKBnQPOClMRa3W1TWyBtK4VdcKr1WIZT5t/wqaRnpCuhI4A1mokoYsNm2bJvgQv
d81DpFAzU+Z3PmA7735hIR9wdAEzHoXKdJF7v+DBFNyNxsbu+phJerlobxXbbUO1
DkZVSxH3d8Fbe0SvRV/bQevZO06wO/JuIRkPbMEGCafwCkoh7C8HIWVObi2b6Gv4
wGinBeYnMsbBGhVjPqIFymHtb29+/LHH5yCRmG8u9YDv6IYzGHMTxsaCYXUAR5FL
E7QzbqWMcWdhfImN8wOZ6mx+aa8HpPzLPDRUW8IwJPZO0TuEO5p948iLU98ACz8D
x1sC/0axsEWY+8rwhmTc27teA/co2i4kIp3F0LVy5GinAivQy7zdDDOO4CIfm4XH
nQDFkiNQ3R7+stNiLXUE0uX50Ia1WbGv0sftx5Iqu5ZaenYXnofT2POS8xSL1PIk
VhRtg+33ka1fECYibhZYYKeAacwE4ymc3GnBm2EL7UcqNlK9I7qDtbb78m6Nx/Qx
Jc0GwGVfDUYG+QPQfLqDYGkB+U8SVcRAAhumy4r/g5LiOBBMC7PNXBVWOxkR87pw
S93pn0U/qIUFGFAwQc+kXlSmQXCLj/64D9nq9A6gsFsx6Ko2YgOxZoWra2AnvJLQ
4K/yYqRj8xDre1g2hu3k+OVwoqhWVOHmrMb6yZhfo29+mpuhGz3Xb4mL+qKHutX4
R0IlhzbFDFIDw9I1JSqXg5UxAIihsHDuSwgXbEypPpSSeUrZ8GWm8ZeRALecJL7X
Eb6cDq27sxZx3QgHOm5vom1xyzGYittZidwYDgZ09pzKxSGKYclqjnUQPICw/WtD
Oj8JN2Ndwn/majblWAOjUDr9F0ou3Kob5GcfeiE2/9SiaJtaXsP8kmlTq68pxcd3
UtEW4BGC5Ln1leK0/TuwUyIZQIQhQwHBUIsT8xCtIPzf6TOk1sjJ9a+jRoj90jV5
ABlNEe2Xmec/2/nqhzPC8ClBQCRw9MEVSbM/nlYTkpb09MEYCGJAubAkPqV5rssF
FDdYcjfIjxCkXt/nLjJF0T45u45Kgj/A14fijSRntlGN53TD+8SgKQAH8E2aKnqw
kJGFHjAz/XTQlsWUUtca7SJEcQmVO/fpo/9kYQ6rmWDzEpANX8QQRzJM6JqmGY3t
qEDzkdLsJnzfdigkvmFzrvlMFsayGaS8ark0QpeolBZVh4/lec2+DMMmCOitIzBE
Rh4qLcXtXSO7xRMfLWn+bNuRaofik7f+LuOGnd12ayfwNjrPoz3pBLfyKZ+HH0Ra
pkM1X3qJjOZi8RC6/lDK9eCXlMNY3RzVDoahbce61OLT9ZK7rpFcLBtPE9h5saT5
FxIFHAGloCiG0fjxUPPmGWJM53aJTE5cLUvh7/4PVTA7O3wfEcO6imQVT/2Kw4vp
9u40C9IvU150cErK1ZLKpRaYXX7E9t7VCPIpVN1s4xYqguQZqbJRbe8SoCIJbMo9
jYD7QSCoBkj/OSVrGsloV1eshorWGTA7CwW84GEDD9JqWjksTyP6tPwOxHE7XgDl
NAsSfpdtmSFzFq62Pzy/cpDVosUEZfgBx6BioIuqJT2IC0498C95QQ503eKM2caF
mtohWUXMun7Dssx20xNisz6e7Avyi5hHw2iBkKytA+wz9QNjELqDVh7F0ny6cYhL
E0Lnem5EiWtIku9fAAOUSfAsdjmoZP11nh6ZmbLFciAiYkAMA8dkheU5kx9CNbFS
6mIeSleJTk0vXBmybQisyMPyWpATwrJdkFrniVZLeUj0ZArWx6wAHpptwtwfAPFi
h5zXLtjmEB0AtCiZsFaMYqP2jj23RhAR+P15tKhL9z3CzoCB0EaSWjLOQmSddKt6
`protect END_PROTECTED
