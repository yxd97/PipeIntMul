`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rPVimZpblknEYIfPIuiOE1g4dMmhwqdbSK8Dd7uoz2cqO0PDQPsUNO9IOyAVuqs0
dG/lrEIFwwYb3F4x2QTnd4N3VIwNyYZn/FbTYon7fst9djlS3ZPFqQvLAPIKpbgm
2IVEwZEk/VbvdYLPRnm7jZZm5AskF72sFBxbIVSIFoIhRPmcuZq04xasXp0HleaZ
ZsixGOzJHCqLqcG9LpeKscFBt4DbBoNmqJXm7+YR1YOV/FyHPmVDvgc9lfjtnI4q
NXgikQZMSdsR4bOQxgl3cGN2Kqk/ilhSy6SrXQ9iw0CU3MG6s3upNjRSKWmJcsvj
8r0svMRnxsQpTVRgjMMlB9wup3wJ2+BVmViCXjHbvxHYRsCrfD3gKe7nPl8yAAO8
eSFRwGnDgTB6Hjhro31bb1kTx/OVkJREf7imcUso6ng2MGWKwcbeNXRiJfkOP4NT
K8/WIzmCrYV6LFdjlEJJdKtDrL1p98kBs55r/j0cXih37LjbBCk06DMZIpoO1LX/
aEf1KSYaw4I3pVEdCWXGqiXdq6CvH87nQSqtX9WORXB5wSrcUAWPiUJ3DR1cEEct
nvA2wHB+/uqGD+FiDxGRq24hmlM031HpgGa2y1rEyy9FRh+U71CqndTcXtXgNUd1
i9vBOYFmzLqDcpAe9KAza3JsdRM2pFHhFyE2H2oyEZDiNvHx1Au1QFHLnOnhJB5b
N/XQWzkrrBjHS2IVxi6xRvyCplpG1rdM7miueSm9D8gwTEUkZmG+Zgb5Qh5i1u6S
d9aOlCXL82yXXRBsugUWZLx71qpR/mVSI3mGsF8URlu6S+oWMoqncdi02ulh3+f+
VEIrvyVXlGe6HcKtJLOYrl2ofsD7mwaFJn2Dug8avp48/lz9PUv9viB+jvUFKzGV
rxutZN6r/CRqbx8armTjmmtH3pbey6dHYkoC10Z9M2yG4GeyvEaeiTOCwdi9pktf
9IuJcfqUSqqENQt8JImPCMgumCCqIguyp/iEOGoYkFC3gA1q/FNh6CvEEHKDqNOq
ATmZf5ojtk8Fb6JJ6qvZFqxlwu52pXJ3zQmvVNizXTjS9VHU8F+mFdUTlHKVt53D
fP3vvpFXdqjidcCXopzGMIzwtNTWGX6PFQ0Vlk6+Nl8l2992NaEm4lshS7TJTRtB
WZDz/5uL5m7OWMczV6OTItynrdjNEiFFVuVr4dqsqcIV0+qwVnALrHB+hYZPCkR2
B46kuuImJf9jLQfUcONqDKnHi3qjmMdGyqE3BrfniEP0nfNJeQ1e7d+DypH2lIiE
qtQMM2xU44XZIXL3FhG/DCFbaCVQ8RwQg+mqogAr5lw=
`protect END_PROTECTED
