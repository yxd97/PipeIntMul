`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jalpe3DVpaS07Y5btJdwdb5eoVF5S/aLjy37PISlzRikGkU0ErPFh7PSp7fNDfd5
xpCLDBz4HM9yn23oeiXACLxyuv0H8xTkambgdn6urVR5AVLy+65z9SqruTdlBM/0
wL7ox6iGH9qCWbsyZojR8MFKI/JDAJKon9qJ4W2HiRLGWiAV9UajVvqxDi9h1Crz
fV0RjyjsLcqjZrTuKDAFh2vGXBn41aKxwxe3v/NG9Gw6J/36XxIelk7VugOifLyB
NgTqWueMh6TkcmI6lB7GcdYCtz645jEJB6euleYRoYJHUbzjwMKx/ke6wFDxSLLX
ERi7+BR5YWRYxNDJlNPZLlQelsE2YkC+CS4WefyVkjCdp4dqvtTS67puniOwnM6i
N5UpLs4Ury4SW48l57whcw==
`protect END_PROTECTED
