`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RG1ZRZUBV31E1QukgE4nPVzM8VQu0Ijv23y4sPFWBTEBSyTmh094fz66VR6ffEAB
IeaKdnhB2zHsGOItegMyg4Ay6JilmJsRfr+Ha3isU0T+0K47b6McbbymDORnP/3y
jJAFNCuCORCtCO4r93cRu9vAGn3q4e3sQDo6Z2zEtul6jAOT8OkUj7086Z30Nc3w
EGuKr8tVRguPdqcNdFN2F5mi1jnX96t7fpjKJMKMfUBbMw+KAz36c/cqJZEx3kLk
DiIn/KzLLhbPkI5jcFhuq6DWjcIsUxk7metDfcLGu2SlgXGX2pZfaPPygEDG1Tqh
WUx7CAClXxo/k1TgMKplHJyMEzUmMb6B+inet4U9J2n3L2WT3dKty6XsTu8Ho1PA
Qmqf31BWivPL8DN1xqSXEw5sC4XDLNJlj7BBaffgtTUEg0UNUYpvklvFcjBAwtt2
F4BZM2Vra6uxu1jL0fZxzTcD7Kl0Gm7QmcIsSkW0aBiDTfFLeq0FneeNUXAippWK
mIjNpaW+DkaHPob0zh0LQmwz3w5VkgEX5FSTaq2jY2FQ26gzOCNJUOCp2DJNSH8s
r3TcO5nQj3Z0goCk6S0lYuwjtxQ3jI00PzJBRpy3gZkUwVjg3goF8FPA0rPTcs7J
Zb7fQwglqtNmBX5byXwpLWWGcTRYDcY+Bi2vT6XxSPma5nt4hHW5wnItmAx+aJYg
6LvQkKFLB5fz/8IqLPSsME1UC7hDEHiqrrXUypXUnUxILGnoY9eNCVApYtB0UuSV
HziRQb16m5KUJThvLrrlb8/oPFDCSe7eZ2c2nChnMc5gNYo18QHYJJYO3kkgZ469
fFdOVKv5xjXM3BLiOUv3ex+FvFyUFv6kzZwbWD2WrC2uBd8mxt1BO781EFbvBnzG
UCXkCwkfU+hhu2rMy4GJFB3qSO1/pmVoHOjPsCba1P0M++guyVqyGGE15/1bRicK
9N7DSKTGb9YZ0Ewv/5ey0Yx1qwuFE175oaoU6FwwJb93lIceMChh2ZUtMQ4wbpTj
PNCsjzdgcajon+xv8+Ssq3rzDgUt2YNgCc9y7Oo3MZ6yHqhen68NCWPp3LL4Ecq1
5zVQ6AJGck0F8/kG36JERhXpz0zy1I7RRGTCcLC6xGob3UOD4pT2YVsJkTU3zGtR
l0/JNGuMI7b2sG9F/CgZSa4j+dG6DkOihf0Wb889rtPgjoGFE5f3mSRMDX7WNmCA
O6WD+HN1aNLSSj4ZbX/G1anzrYfL2/u8kiYpJnBEaH06utvNjLpOLJfhSK2DioU2
hMJjx99U/7Btfeg77raXu1sotZiUsbtlisdkIT5fhKS5AeCBwNpsyIZsYlcdou3E
+/qbCFbT1D38umNgTdJHEyPBDsjPGQvft0D7/r1+K28vcP3dPcEwcg0KwtqAArBW
QsncNwyldxX2cHmFTT8lnwTNoYjsXEMNaWNWq5kND95Xb8uVsue/V8Adz5mDlI3D
uEGA12j6zhgpXiethURnuOBafOY60XfViju2yUj/DSmNETFrsG3MHO4f05yLsS0H
6ied49q9II1EuwK3nohpEH3c+SR3L3XH6jWimfvA8Bgcl11WmCjUTcQaCRnoMst/
0MMnQEM+p+BtdQ6XuvsPWaGlaI54WcUeTZYPFRXMl8LUMMQeoXYiLbdwDAJWUlNx
sJVF+E+9lDadObwbbSiVqpFfi8EPnrueCNm/8qvhRv5twQ9KHSkRbCbIhPyFGsQw
6wrBBptdfOBuclQdKQrQxgN8GttHm7jm2dTuUsphFOrv90r2dynq6KRKBA10QKku
r5SHXdj+VXvkIjIxSs9ANJ+FTIQKmms+GXcuiPbpulbAXGAkyC7o8pAd6TCgslQe
R0AciFsGKsBAQz2BTkYcrrjjyLxs636m+mXMN0VMdwtEblRCYNUr1Ee4qY0sHTBC
hhNRzi0w//trsXKR2LgcTfCxWuf60GEinObj8y7ga6TMRXcmlY4vGNuPyaqE7tvi
qJhkXz4MumiLkTPE4q93FLbZLQpKfR/u6oAS8bSUDaMbgx5LMxky/pcP6lN9cJiW
lXKNOEtBHJAcR1YvLrUulJ3AXtMnWr10N7LqO6VV9YU=
`protect END_PROTECTED
