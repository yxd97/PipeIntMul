`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtYs2NCbnH7gNoR3z8u23QFflVMbgrDd+W9hiAlGlDnjVUM9kKx8TwUy++Z6tIQo
FCbtS3yAlKsUeMtHOMKal0VfdSs/VGs7nwyygAne3Eb7LePjKGTCUoy8hcFLaDZj
MkvuCW6yJ1wdyG8tfc/q7TcwoLRjT+ZSFW+wFTPK2URfnW0yZ2U3Ymcrf7srp4e+
RBAuKPDlAGj1LSeqXEXf0Ue81lzKoP22xjqo9rghPo33ofjidmSSJcpcIig2KTVw
a/3AM8k8hJXdBvOeL8o3Q/XO24lbIIQ9mpFbBtL5K0ZTEGNlbSAcPPRgJmqh6G1c
K80lLYmWTGizzMnk8D/A71XUYv31vqt86ZabOS5M1QpETRutRrZLJiaU7aus2AjF
eR0AEZrCjNnZegTCzJWndA==
`protect END_PROTECTED
