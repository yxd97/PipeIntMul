`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ksZ6qlHGUP0iP+nzykbWgQltWKtIJDOMr70ni81lF89GWE1TEppfGcOf1IkU8QLj
d0S/k66k7h3yA+UScnBslE+F1pKcbaM3SSUYyaaQKtdKCPRiRPdzsJUvdBUgmAWu
lCZPzPg4f0XCUtl4V8Ey2bWS9eNetabe1m388Cd+X/MSSiylBmgF1mLpO33wNUm9
k/maqUTbWEGjvcAyDoKTOf6pxUwMq/QNfgiiVNClw0Isw+e7RCuFYAwfRlW99kXX
WdB3Wwf6wOYSkqtWovkV/U+EvuSge7knZ4UgemFCRX/nyDtoAX0oMAqj7EO5frlb
VotXmrmnVcPWm2v1TavWz1N1ObmohOomYk8KqNb5BGlBI+s9I76yG4x1kPes3gP3
bzff9A6q4TJ7U2aS/2JlSXYkV8Nt7L6+T4JSihAPF5+dNTc4YZVGKFMnIMo9MsPH
0ascM6XMknTsBm9HcuNIQUzt7ogEYP+KpTiJORuVYd67vjsSX8ZJv10Y/TGjX5BU
NWUfotnGOP2BBENXTWBDW3n3HZjyfwaskFHCVJQWmaA=
`protect END_PROTECTED
