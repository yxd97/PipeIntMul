`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RRyvbHBFFva4WPM/boZ8D+bzEwl8Pten8+wtrosUIk6sUlZoKyL1Abfxs0pLUvsQ
/Kt8kx+jbzD7L4JHX79J2Tv957o773h5U96MBxh2eFN4TIGvkAkRWOvc+yYPVmTq
7IdRh1P5GzIPvxa6OEz9UXLqwEyTRyDVN1Z9auE/VCHre+rEYPnrqLn4ST1ZcvmR
tVK1ep+R7qwAucErQpzujwoIAao/Vl3okTuT6dce98m3g5teX6kB9C4j2BOUNmFG
wXmANMuSljvTcfelFAWJ2jZnp7iWztP/GxPd8XppGCu35CoKu5s1/un0Js2YLm7P
FdpS8/1LDE3vW0VbIYcEF2Sp1Vwq9XEhp9Ww9fE6ls3lyEsOH08QByUkwvsaX5Wj
2vT2Fiy9J5RkrqCwHiDVlQ==
`protect END_PROTECTED
