`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YETNAHnLDmnCQFg6JLPVESUqk/dNm8JM10021gIlfxOnL6SEqrn+okDlO3c5KuDE
aUOVSFo/Z0G2LcTFWZypIrhgvjSfWVZUux420cIFSPs1FfsYZ3kWjDawnbydtTaf
voYw0IoTfFfgcaalCts2LvgDR/NFa/a4jUZF1na0y+ncIebUZGEyJHIoE+lXVm2I
4b+dLBjP5K0Z/OqimJpoELI9Qq3i7l3vGnYU6nxLXqbY8FyB6OnE1G44BKfmRKqt
Ls+0PoVG8QZioz6sxLoYEMkIoYzkauW04C4WzIZTBTkNCCksxf8VcoxUxUe1UKNP
Zhi5egmTDPVIB14QYMMNixjtapUsyw6JAn2kKlsqkN63Ouljh2MF6SsYB+971KiS
NwuSXGk8JfigC//tlorcwiE0c0DtEQ1ZYEqrGwdjjeqSQiEge3JLqt3eoHnN0/M2
iXirXrIxL29dTSQUHvweOoG6cTtjjHg0bh2WMWrA0SyAS21Neoz7dBr8BKF0ZYU7
PSZQke+ETueNU6cYAjQj3J7I9gbDjfB1MPH/v7zoQZTXYcqOpLfu+HC4PX0TNScP
j+NLHgAWiQzy3dnz5+22hLNNeAQzOvGl7SxTk/c+ASjYufEULG0WDF+L/8kuszwo
`protect END_PROTECTED
