`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iqrXaWf6/06T6SaK/QgV+2W8nd45nys/FMW1A4OJMbdpGLUbWI2GXc3Y3VVTxWp
21YcV+tE5Fw0UHfgAhbO4p+8Ws0HvUtXNz0jQ/YUPvd1mFbkwTJXu8P4QRPWWUb+
JeUFSm3m4RkPXEXLo/USMck5UnMGZ7FW0SUhYPbdagC3dKVCZ+wPQ6DEu9KLCRxG
79Cd3U64R+juXBOac4MnSbXMrXQ295e2ocaAaWQz28QTmX8Fk1obHJKLAAVqyDen
6TuiyY2Vd8VZst9+P6end1Bh8Wehh6F6cIQwqkMzK8yvOV2Qrh08I370/gs1Rwz5
jx0+YHHdrJQ9Rj8MnImHqWIpzXXoRx/5xmxl+a45btoS+DPv2eyNCS0z0zITA5SG
wiVT2CjJjYX/xwEWNj4VCeN2n9fq9g/Zl/DrEXtLIVdQt5vyeL+zzmBHB5HNIH10
hWaTaJl2t4odJ8ZmRZ2QmyL4ky/lJD+Bpf8aMcbBCQMW/3bEthZ1cTZQSK2Pxgw4
iKPTpjT/6tf8ual0y6K5Gm9oASjYJ9jEGZIEy+GEHWfkgyVYLsVfiMNuNTLz91zR
CmKM4kq6lXeYy4Q6aAY2KRD3AnCv13XXIMOIupf1zizHsA031RNRq7rCWYygxmmK
Epie9xp/fWWjND7kPtICMERGD+GUgspUhKxOJNbgZD18wc8Dx+4ZPquLBzQ1kMEo
5OJjob08PJtzz8M90krYa4WCaRaRyggyThNrVLWUpo+dW3wnndC8V/bjjDcPbh2S
xE/lKrohhNf+PhLSHTo2IXDcyILudRhaG/L8bfYeNcOtW6I4kLzos3/QIIsUCi8f
hqXyvHz70rdLtXOja6Gsygqq1dR5vRVFpB72rsBAAsSa+BTpbGdiUiZOHjr0Oev6
+K/HDpEtCqs65a7i256LTgDx2hJPTwXu1mxsIlWqT7tS8lSezEsFBdWgCRqMYElW
WbBObZ0Oh0wrv4zoSULrxW3NLzqWHdku92K6+9nEl7Mgvm9n87DpmJao4wOdG1nf
vwPY3kd9CIwNRzx0VAj7Yw==
`protect END_PROTECTED
