`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiqWbzTbU8A0MCVbCYj62IQlPRurFNhCNHqdkkf4QNwo6WeuNytQfEdshEqOu2O+
S+s2Da5nnEeRCxXmeAeUoU1IS7UcDisT47ZH2inhMpBoPK4nITJrSpwavB9ZkF1X
DC+AxACB2kMyDj3b663oQDFvt56N3bVvyoE1SqcNAxUp5BzPz68LnjEUBc4uK+YP
ttzjLF52yDVZV1MdVy8FXJwRu6VoO0sB0FdIx+wF14gLieaO6G42qGwsXUqvXKTm
Ik/fP4TMuO61NpUHOSaBCmnIBiXleWiryHuHMWe0FFxCNRrFksUEkzF6cdOvpDi1
UNKl2WDlu9gii9FsPXmftZ+iXyrkZ2CbbeaVbHgZc8S0KwsnKShZ6P92FK+7Zs40
hpV9wQCIXxsT7CDNZCRGVjlNpSN78fRj9eMuai1sZDb4wru0mEt+8tdk3qJeRar4
q04BPYx2zAmT4BdRiX2WCJm46zEwkRDY6IBCQQcWKVh0S2V1gCFMWtXTaG5TnUkJ
umkyvbNeaG73djMlXAQZQqYwZeP2njF0+JMMEkjyOf4RzSpo4t/WCUyc8W56V/74
KgzfkSUTuukDbl5saYJawsvHCnXGXHs9PxAV3l1CGqbo3wor5FwAiJkpgYPya9xg
AeVw8UddXRingKCxWx+BJ49yrPLg7CO2ATT0avum7PDC+rXg9jdJssuVlHm+thGL
7LtGlRkf4LiBLErdYf9NMzmueagxSO8kZw/ZwkVISHvXyXKFPVtQ8i3gz2AKKYSP
dHhNK8Cj8Wyh3iS33iNcvn7WXxpKgjd06qR8fM41BlMdzZZIWdN7Iq/3ozxck5WG
coWd9mRWY/aKLgILzUSBOx7V3BdAMyOXBvgBA4ZJCSmUSGGtKuzOqBDLSoeHDcFJ
wx2kbU1w8DkB9mlY+iOaRFjvzJPdHXhemh5lKbfiJb70ZwbcQBotyPI//KICdw8T
lv4dT8Fq9i0IAa3R48GlPCNkRzEkflgqOXeeOi+K8f2uAT9BsOhTMCfnSCKcFLvo
dRS/k/SplJLYn8J7mQPIi1ol9AOt2rYzRsqCg+3bNMwdDjGntKj4VP2Jzvqu5Egk
mqX9PgiNd6E7HZGRddmbDCaofkJ6UkB/SKfQrtbwQ+Jgbx+cLKeBIE/isXLpC3GC
9LaGdtuYR8bkFbql4PmTG6zruVqfXB7lMi65Rov6WAD4osjo9jj+t+VSj4Wp7ylZ
qujqTTxpQ8m9OId7TLbMHolDuEB9F7ErmmGe6GKOrC86bdGAF27+HOUu05TYUH/a
523QTYOt/PXUG7QxrFm/3H3PASZ499SAfSRcHiYBlMzkMeGasJnLkc30r932JarV
c2XVpGcGKWIlIOkffhpDoY6E2FBT/DDtU398vz3j5bOArJC7pnkvoxYqcBb50o2q
42K6jm2pSI52Q/WMjMkDAWAY/e6T5RtbIu6r5SXYWHZ5VRxIK1Wxfo9xhDNoJTYj
22qU8Qq966gGY5oI4fuulJ1pzq8W4H6cuJ/l0pCyVGAx57PD7/NgS4FgA7d4og0K
DYJjm7aBIwo9Mty1KJAO2iTHvkUAKQN/cQR08ja9Cvtlc5rlfa+vSBLMWuaozjl6
XGIuZWP4hNuEFczW4uUaeOOc5BTzHKlZ+Cr3TBsS7r7CsQsYSf+zEYRqh107PvKC
4Ib5GPh5AGBLey6KAEt2lNJviiWGeu8Xck6weN8/mZD8KirYl4GcfZN9NIu+jFb8
hiIRAR4w9KivqNZZhlJbqb5gfDCDRwAFMhk2BO3WcAIY/qykFc2kEBhHDlZkWWhk
c9vvNg3Ek+sIhAZurRxWPPdcmNDoVE9FGTYByepYVRfVjp/DVgaEMZ/2XytRqTur
5YCvBuOit6MKiohZHcgXQH9qtv9wDlDrufYZYrmEreq+IL0WDZd2xDvLmCph5fBc
zYlKXOyOdum79CP3Kkun1ROVCDY3/PwJW/RlO9tE7OU4rSwe5BsYCxT8MT6qjKeM
5QulWdMQAsKHDvUsu31Nr44MhkKi5FLDwmw6K2Oi7Q4PbSh9XuKvjv7zOt5OHmU+
AQulPYnKAMXUIyUxTMuogG/7D/wMwd5Jo4ygAfz+WkPjGyYKSA2waU4EzhvJbExI
WY0bBBJCGWW4QTZMvWsR2KZfelCT2KoICOhPv7rKJysNfpBmiVZ2n6UG5mbt2F9T
SEK6IrJL5rjXhwMKHgYp0gGCxHE5tDAJc7vUdwUQKL5NX6gL8v42djqvdDSG2XQu
H4QVSggBq6Zx6qNUVegSM3lhWDprpXz4RJplaUAgbtn/DHgRDrWNA9gb7ujMF0v6
DXaR9JjB/JQlX+FtA6MpKKEX9vSwmORiP2XGQBQaAnmT9LxAOefySCEhpUa1ffuv
rJnZF7m1dEvOEvGAYBi9HRHd23x80KHmhdWzlnH1/VVcU8+HIPz6kjQCvjkqzV1/
6FFoiFXBl1vcdTnoDTwEymTBobqSm3qrt/xPMNVz7CltvBbGUttUpFqK2BTCqGfQ
Uy6+3O8JxJg0HK6+8M3hGsmeaNRhhDY9t3naakeSX0VHS7PiVqsXw4s90nYVHjYk
lVwa6oQFOXHtu/do5sHzQk2s5gvuauEipzg0yVGjFBO18hh73f+Wdlk8tr1sykr/
W82HWGJjaxzWitzkU8gz6QVJILUI0KZtgb7PEu+Id8l7/TLYL8ByBw6nCdpNN/lJ
7vak70s/xh8iJ/2k0xiL6KylKcO771vBsGAlEChrSGN0kzZ6sPLAcxV+C7zTdzt/
m3MFEjNOvs/jnLMWVxSdE2DbZY0XMuiQ/vdhvfqXqGb5/pygLAp8dkGP+nxctEqw
qzqYYkYtJEU/K7QxmQQENGI7uMjMtWF2regHXzANgosqjySJ8ZBW7ZJyK4SoJuUA
r4oOde82k7TA9amQm8LdEEjQZPe4MLC6BcQIn54OlWMOV5Z+yCTAsaq3n2zAaJyu
`protect END_PROTECTED
