`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kD/l+3nRzgd1vr4/v/17dhQijvBtkprgWub/rtgrhQ6f8Mqw7Cq6QSGOYLX0lYEL
DK2RZWOZ5bj93MaNKcHVV/g2DxxozwWHL1VrFWEA8El0EAqDbSYGNqefNVyu9NN2
JzFfAW2b2xJt+WF2Zqvme7YAoFa/O5gHGm/Fvjkq/uKu08rz26uv58fjPkatDn+D
JXAddBqPytwXzs1VPa9Ch4GOfi0bD1X2gGuyOyxs+9Qy0wyY7cUKz2ijfQAdU5VB
ekgcPqJ9H+nFqgcvk8s48L/lbLTCNRJBiYC2TiCt+YMuqL6p+eASH+PpPehqOKE3
VFoC8AcN5GbC3txSknsIhIq7YIHR047w2bYgrBUbJmPApQitmUIdijfq+B+OexMm
xVI5LwwJX28RkzgN3bqjT7fiNe2W0r0kMk+ASI4uJmpKUhYIxi1MsqUd+aFRUHU7
xWTPvFuEEi+evME6Ci8wQspXN2jialqRsCTZrl3BKdk=
`protect END_PROTECTED
