`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypXBu3o5sxHeTd2KtzEarA8bGr7l7aZdaNyWwAO/j9927LfqNkEp3DTlB+dvlf7F
M3nJGbWc5MCWtyFggNztNE2okYM+4aBC9vA8qotePS3mmVeJjWo2pQUKQ9BIqJgu
fo2vqh2hM8s9RLpUckUyghQTUsWDlkWzGAM6e5TImYEupwHQ/QNRPUM0XQkWlcHs
DRY8XyKlDQfZBvvzQGkGRacOnqCeBbf2LwHE7ORLslJVuNJ1Yc5C/Bboh0HMdYPa
9n9g6zcRhWXVlyKiWcqt13sgIECyGVGZNJt3LV8ZRBsYAue3K4l5cZtIpPTv7Qu7
syaXP7Mjd0hgijFLkiIZP4X4a0oYq9RJ0pEuX/UOz6LHAYGfcBgwN5j030+3vcZK
hX2pFD/GyHC3XeUEXD1RLFbJKZDQGkaTEBHozhzZtBkb0LKNZv/35KWq24ZYEbtM
gz6MPWuSqn5YS+GD+hdvV8yK9/dpQQ5dhAAoY1kcD4RejeL2vP5vjp63AzGjGGdp
`protect END_PROTECTED
