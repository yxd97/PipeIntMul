`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ti2mtCnjI94IP6lJqK7qeMeZirj/E0uXeM5/0QfQE4P60y9TBtr4I+4O0z16Hdw2
Gcyd8f+81kBCjkoUzuixh4XXNFTRrrbU1Pv2FkqPTjU6afZC9a4V9TnQ7SJ/kkj9
0XJZ4VNVdPrxM2B+dlLQDk1+8wg8owD9qOvoa9F8xpc58XAh8Dh0UwosjJxG2NmX
Z9AAbRK5ffLdZflQPQefIzTmCL/o98PAWdOM0kzX/JRE2uP8b1H4+JJVpXVlpUER
B4G0TeRKs//cOjnaaJ5Z7m8uZfhUxQVACdz10Cr9eFtVrgY1auQHbBaPnGxdhlPl
1995a4HZ87z3I8j9IYmMSNDiWmSA9QYz8S8t+z9l6aM=
`protect END_PROTECTED
