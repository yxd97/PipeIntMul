`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OhP1n3fFbtnOeNFbuThkXbWT+kmli8kEqHj71Bka99DGQ5NeRpCuNWCqR31sTKp
RuAmOhvZgOYKEutyh+8pS5g3QyLK6iTXLWmBX3l6C0GUdcH+hdAlVDLlmkXInhMB
cZzmijnLZmMS3CaY9sfHGO3yxbbl4BHU6jo2a2dQ2AyKpP+dSFln8QcGClNNMe8F
64AFqJCSYmuCHCTnV4IccmYyBwKb/3fneDnfRlDJO8yDitH9nonbPhQf+BsQ3a4b
ZgQO29Udp7ae4qIyVJCrYCJVxkoP5bqKp64M1SXjDwJLDvs9BHuv9UbpplyhDYkt
pXOLSaHimEe4YdUI883gRZBUp+JcnG9Wsyw4htxRfqmmfTbtevls5VmmDhirapuF
dP74nuhrfGWuktpv/DEoG88YZZKvC5QXBOCA/0Wu2LKtKmnld9TfFbI6dPRT3s68
XDyo9viAsvuA5N5jo8+wkgzm687e4zVyP/sHR/iEpY2CCOGkMCbZkJw8y8Tmk4O6
fasYp3+Wr2T06l4Pwdexl1T10/aRE0oEPH7e0e+Vf5Nxby3Cpe8Fc71cg3fqqCBp
LcDGqt4VZvPwLMuRVj1UAJ3FEq1OAPdJaafRVWeRrWRAbX3y+PvXjGEEN0Xt5Wqq
VdD/6Gs9CIlbIxLhZaY3Vs9o/6oXD4DC81pP+ZVAuXvmqeo6OPLh8qnY7nIggqW7
7JgFToBgx/TKqeVxONOYa2Fy9Hk4wNyfoYd4/d21m4EEHH2litLameHNwnh8L4Do
T12MAfPpuPJo9fR8GHRrskQhpouJixLsorlyYf0AHJF/gm8UwZ64yfbD2hdX5Mk5
3Ekcp04h6WZ4oF34eLkAngfTX1sb72MG9E4Tv6jyIttokZMY7AJxNXwzgZoARCdb
LXI8KP1iHlBBVJ3Y+H8cWcVa4hvto6c7OP9hPgr9aiJzigT7Z0ruMaJwZFa23in9
RLGfnjp9+KlJNigD4la4wfo6QGtkBkCzjkY26l6iXWbKsEfdXprof2K0lYujDM+9
D3VFizETKn6VfSmg88HhOVwNotYRkA8/KB3OwhZR9JT6xUUWcQJ2aT1cy3UzjPOP
aZFuA6Q/B2F+NzGm2mefyuyrBez7mYme823e2lNsTVoTTIdfwdV2oT4OhrLQuUrl
NFwLtdnWMn0ibgJUmk0Qt/EF5RRRuij5Acydyd/sCofcXrLwksdD89UWD5s4YGSJ
TtGW/WbcL+GZDUD7HqO6cr6Pb/w0ldaL3y8nxafdodrRxmjZ2sV+5FTbBIcsXjDy
Qo8h5FZs7u0UlBoGnCPDCKkwzUQ/EUsy3wPGMx2Qs91yrvY4g9j2iFTBauFiVahr
y9R7/IOV3I2MP20SSlyigxUItYqVt6GevnzpTQOqoDy0Ii8FrAjVXc01CbzdF1pa
ZE+bEIpAMIx1nBMlhkE8zIjRGZKvS8Nh2i6L17VyxWJQVKyGAaenucu/+6J1wzBy
T51LfQpqDm/dg3F9/aKGWwokKYt9zniL1FQSxoVKxdvcvhukGiQbyvaZN7CobSsW
y3vdH3NWa187Cp05RMgarqgoOn2noRnCDHi0yKhdAn4zxY1jshVWcLzW9YSypHhV
L+NIzPPiboHTQKazqs3FZQCo/YqVbexYdvO3W5UDx43iUayKUB4VnIClxJ3uFhYL
JGUX8O6AEbW6zb65ocwxxEHnX7UW4rsUUYT3g2iG5Pm9bSPrJSN5v7GX9+uZW5Ke
+DfcPesbffJOm1sDbocSvfoYR49U97qdZptiR7AQvU3qC8r30e8dnmaOxeZ/7OqJ
OAjn9XB8WC3UMmShZGG/bpDOuQU2mW3jYQm9xeaMUzBJu9NTpaUZJHej1L9th9p/
LvbkzXQHAEAY9nX/BI6tMxisN9ry20YyA2xQcXl/Uzdxxav6MEch7hwBeoZfzXt5
yz9WTAIUCM3tcfxhXX+Yy3L4LQdG7Dm8JRLNY8q6oMAJ9YTxKhILvPnXLf4CBomu
ttPmbIoD5vin/ZzNM+uOaNiBRGLKUDnecpZ88574WGpSP4T3QUD4Qu3xF3f9Awx5
QOnFvTcYGLPgYKzqYq79h6Jul8x136ylgx14IwmMmklj/mvP4qhqxSSNagU7bwq+
y0Y42aiQt6+HSxiKLbrsZWfwWEXZcAjB1/7Ejp+MkLfjOdEyunwmbQ1mx6is8zFz
cjYZF/BGXxC49ASfrf7ze2Jmzqxij7syKkpdhytSYHveP0BpsR8/Ww3NJNnGnrcT
1VDT+gmoCksXozluMPhhZj9GoJ65bwyF6/RWi1GEO/NmnNQyvMP7tzTLSkVUmwef
UmOMX+ZLAvK34/XKvbnY1+n1wuXLZDGNrIxx3gXUSt1ACScdL5xbOSzUUZ2S49wH
rOTlENA70+v8KQC1tGP9BA7MG/JsA0Bg9gGKFXDJXJBsnWaZh5xRP9LXMn1Myh/l
TmdSkkwX/5kyMAiouImIyLkLePTm1SEMn8ccBwQIOGNqIs0Eyy7D6sGr46LIdBqD
Qp0N39d1SDzz9F1JlRpi5zw72nhSNLmbTNJ6m00E5rBOLa6gNCnsmlQ6HIUHZ+Qc
WFS9w4LDhMPQAmx5ISkqBn2JbLRUViCnRHdyp8oufsMWJxGkeYjOTUijVwE58404
Qy6doiw3z6et2d6iD/sNx1AqUgoAdAhxAzCV2FHeutuXZWBSJuDuuSfbgr3XyxB1
EXi/IW6zq/b7uCu16jVn3NXt1j84dp/+bcsKAqv7HAx9sTb7KBPiDW2fqMRXDrA6
IwE04kyyfHxuwHHuEfzO4ieepJoI/SmULi/w/dqYBXbCPOMgT0j0dl3oLG1RgjUr
dJ3Vf6mfzk1zEbQ1oeCqRAmZ0ehdJ3UW+1vkDpX+E0ycMLcQdgTyQsrWBc3RQYYW
gz/7itiickxhORseEggkqACwr308J+v/9p2KqdQssoqm97FJtxlvV1X5/Fg3do+6
+pKFjXTPWZlfmGP9sx09Z+TlElAlQ1pR3qoKntOKJTFd5BcaLXa7hZfiOV2st14z
w2h/uC9RoSt3sO+uHS5oL5mgmYV3RFe1G2Wzt0OAM3GyWfE0M9GoFtshMIvcii4o
gF7c59hFOysRBmZ2SKIF98oVh3pvTlX6kCyqHa4I9zMQBJosbsJ01k2lR73o15jf
I5t8xbtxoSPYOZzshvSdG6vCwDZWAWTV9cIDugAUDKVaTZZnlbBCX2RQjRohp/EM
WNPWRfRGT7BnWknMi04GqGw8WlwgjezNPWtnuLHUDDaQXTYfyxBO4z5xUhRmlndy
+D760Sy609ha7Huo0Tk0qQK0Izmi/tBl4YPuJXgSuy6UYeMcefzrRsbme+WKfhN2
g6s5d57hTiEHUMoveoc/zcEC3AWvoFb7bZwv7ypbQqXCNeAdpL+wwFH83trumrGu
jIHbWwy0KieOyFY9UMxd9avBh6EoCqzPnKGB2EeADmmWQUl81VQQKcCwh+jP3qb/
vGnwlkfcB1ARDuRNIE1h9/TuAGFlIQYtQsHn1Pk20w3/QRtoExTurtXVkAy5zu0D
Cezpgq05qp+V0tKhWZt6LmCIgvaT7Z/jovuPbjxtiQhpaL04DZPwn8Fgi5b5ABlZ
ef2t0K34hyoIuYax1GZ0NJj9vKIDlM7+iCchEiT59UTIiEK6Cm83YDwbRWNFA79f
/2t117DaHTmBk9ffZvXCVWqakMNSMAkbHoVc1R8fLcIqgtR6dcTezXiw7uVQwZ2c
GiaH/MiCOzGeHjFzW1UbAmgLoTxY6adjyk4S3G0dC9Ol1mfe/jG+Ij7YStvPROrY
JRqE3qcsGfPy6UbMj9U9Cp9ceeDSr664kppDbgklRPicWUU+i4qKVCFSxokXVgB6
IJIJKXcKIQc/0WVOjQmX9H6jq8W0IBvDcx7RbG/OPnkamSRpoMtMFtPJxcgHvFMI
1hpgD0Jpw7Rq6sw43UvB5EzCJ43Sjr2hMAm4IKl4TTVThDdO67B4m/TCR2eSKqg/
1guz71qITI1jE3N24lo7oPMExDPCTO0lROH3Ek6Y3eatLPxQQ21sRF6db0A5+odg
WfGHKOcjhgoo+4LTv4+OcSOqdCG1N5chSbqP30jlQXkpaENShh8yRhgOQT1GUv5R
gnmBcw3U6VXSmBlP6HXeRVb1dV9Jx7UEhEIaegXg+zHMGkoNF1CxN1m+kH3t78sh
pvXGaQRCPFAMBg/8HKCc1eScDOJIN9jlfGjrC0YBgxd+M5/0/3tjpGX6DcJ4YZid
/hmbHQQyokqrc5X/EnJhEG1/J8jjf/l3lpwbQsofYAKyXqedlwwN3W837/5BslIE
Xcip2JGlkf4cUiTrbhTnwIso8KxH4/5DMFCiU6YAP7cpVmuOFGo6P21iOGiU3N/8
RLF2MzGNV9zE3zdzHdgmRNCg3zJ+46HkZm6O3ViBGVCrguqErF6iTHbyBUUEHR1N
qbcB20gs0ADCBJDDsq1xHZTQY0v1w9eP8Z1QuVkZORtot799ZSdJSkfOn7d4uWEQ
Rz4g2Yl31/ay+2NqU9uSJDXfM97QGSjMm0jcT7pkvmtRkrtuSXKOy6x9+opCEKdA
sdjChNwwHbgrJapU3BYPuQ8Hewfh9448sq9u4TqRXiQM2J3xej3RwWIfYEXpVkWZ
+zPufpSLJyqBSXAWPk8wU1G4KX5BSrRLM8kX60ZdzzQkiLmgjHysU0iUQsz7imH8
UuBn0pihp8QeypcxKUJ6azSaEOAMd/jB1iYEP7uYisIRxnLcmQPrmhgRlSC9BnNz
GtXcgxpkreXnxQFE+DqombBHCgBcGou1MuHCWjRqd9+csMED3qL4+yZsx+cjU3m3
06ZYyEZNnn2ebWsds+WTBTLBRpYiA7Mw0K7779vWVC/OuAHf6lNR4wkq4MbXiM8N
Tk3UupKz4agRoxXxxW8jiGX7d84vHfYi4QsfgKrPgW836HAO77enXVLgGpXkeciZ
3MDCLgn/+Rcq3ml1VE0Rvl6zPsKSwmCmyxhtJi4NmPBorfyRJhlxgnhUjclCzLO0
C9ByTWpKh1bSylRmiXDponsXRNdazcm6NQHn7jVOydIfjhVrPn+ZA7HCEaKM6zCv
rRcJffbV2/ipiVKSvlUVgAnP2Xy09Y+FjiIg8DvmC0dwLd60ej7QLF9HSBPyGNco
hH6TyuIkERfxnvJTFdCz2Aa/IcsoFgb0JHDXlbqY6+V7cz4nSbeXFRyJUFS6eeSw
2p+lwEpVullysQMXVzEvOYnQi4hoUY/XPhsHVR+UDHhqr/sAWCgGSMgaQUJk7sth
sX7QHOJ0+7D0/Geiy8y2+a23RDK4EmlhrgzRdm1xM2M9JyeQgrTkeHGxB56hDg+y
I6SOcgo7b6Swfl+3iONcki9v8zTaw5gHlG1lSkiIbk9AeZaaT/ycre5o9umdJpxR
QrYGoB7M4UfTvg1nQkuSHc4bp7KR79IW8i1gMTX7XCw77AYP0gJhZ2DqriVRw7go
HSNWiQyAuuPTGh9Sww2kvZ6UjAbCBxuCKPQNPVWfmapLOjfkS9nRcEKrV1AuGQh6
uy+jysnUgDrEdy28ZYQwz6SCEheOJU5wfOVKoSuywS9WTgFZGugh3lJA2/23p1tQ
Fmsw1A/I4kPAW/u9Kdrsu/kIcAyGw5Joe2mLOuu/p/nt2KAj7okI1xNFvM6qRO8r
PMnzpw6t06IYdGOrtnBzsJelzx8LpP8g4S8qFnG1zPUfcaOnEPUFPfpD5NhVoRhp
8fgslYevthagkEHLYKbjoiY2NJ6LDLWm8G3yN6qLrklnJt0lroI+bqWufLjmmAtl
QjVB+nxoytpLpq/Ft509pM4vjl7XFDEPSIDOMnKFxDWXfsVfFUngs9pSAjSos2xZ
2fkfiec/7Sw/M77y3PPFHx2ub3NFa/UmVDzT7Xp7L639Cv5viww2Ujg6/T0ZDvwt
/Wz7TY2ILjcQBf1C6mdR/Z49mJn2o2HgaAM1X13cwfDZo+4PPJhQi4uHpowLgrYc
cEI6kcBxguQPuvPWJv6lzpTknQKE1hszYhNWT8MavkKeZX7dnlAR58zF6vyMzSxc
Mj+vmLl9N1c2p5yFuhvH7m090LBpGudNydDyo8tErVqjsVPtCFPMTFiOdffdWCpz
d7Tr9Y8yjaCM0kMfsW42aa1+rxX/Tv9UhaIqtrY8yQIigGorYqCNTLo5OxGrDji5
xbeyUM4qt5+PMxeVo+6D0GsMEsD7Lwn3OWvt9totRPvDzuvQrbdaaoiiSDiPq8pf
uUJ3FYH3VarUIQf3OmO8EDUM/YXWR3aqgU2fzWH63fECckinnKUmFmCYVnnEy5Qf
KclAkOUdhr1HzfzyKjsIDK7FBFBZov9Autmg1cOO2u+kMiGQ46AZ+Ic4MqPE/rws
Z5k70ZtknSkyKFF6uaPqYl/JZInZlYzMZfBEqVmbMPVPejbBD8OSKo/cjxA4/3js
Vz53PkumUq/t8Up/MY5/8/D08mjTAQSSoCP+6rCBbIrdU06bYhmKBqIr+GeesTXh
zlo0E9Ybz/l3aSARC1QJo4YDH4hp8pGFTcnp6mc6AE/jadwNaJu19HueXqD0suwq
5+0NYZ2TbH4OvEQ9+rxLxaJWsNSgc7KOmUDpSpySMyFs11QnhLIO0EzySfjLSxyo
ldrbZC2spQR4Ev2Nw6TcoEJaMxtWn8ms1tK81xE6B7LTjLv4CA4xqNsF/jthHGLo
fSoog4p45lG0mYHEpA6ipgypr9hC7V6JAlYKGvmrs3XEqF5RDuEwILq2YsBo6wQT
+JXfxnDKf2RebxNnb5/gbb4F0b9BLlJKMwKFjgim0k4KzMLXdGoE6cp5FngzbZAx
j0DhZCWwC7V2ApAwjLM7J/y3rm5fdTwSFkkFB/7Zhg1hEmP3ex/0D1HDQtiQNRkJ
czK69t3regY0V/fP6vFr20P5JEwrOn4/tW3XPySfG2ieqR0o8FPb+zZUHs0Wklmu
+WFDAGIPQKf7kPgvapn8Xjnw8AlOj+5lJ3qbFCQZfJBVsGp3gviEaQCp0K/EhiDp
ICN6wa4FmfVSyaK0y/ZkatVD/o5Og9M+cvjVWxaJswnPG6ITnpdlVM47ocfzSHnC
yBhUTx6FmxHSNY8HhMhsALeSEBwt7qxzb0z6mAmwZvMDfo/CtBe59j5Xg7KFHk0j
VQAJZ6JnH9jenidewCSKXK5oHM5PqtoRriiDlnrGkpXlDKFE9REjzh1NTzzA66KF
rmVMmLWnuYvmIiHpn3Sl/9tRPChvpIq84MM0pXU+Zm2aj5ND50aFRkz1h4gdo37n
iTYeJKDdQthQNW3fKykxl5PoNsPSZ2kYPpNI+DRzK5zmc/rJG0aFlp8ztlm7Dcqw
fargP1CCVwUr6DadByUuUsYf8vSZFeO//yPMdV3Vmw1wqPfVfzMQM7Y0rffJ+42c
DLocdwEtFLm2bdSL87u1Py+MbSQYoXWpCu9ioDhXRodEK2hNbyM3ODHiKFEOd5s7
gChDE4bQEiNnvEoKMhRDZHfUwl1qks71fURcZ8HR+EFpGVjFmmxKGn6Eg7bUVepD
oVvPbH6Wppbt2CmEeQ7J7Y0sYr420mySoYgJdLYwvrba4QpmoybPdk0c5t3Bwt4E
WohozIwehx2ZBhGibl9m5plhX84i/t82+SAo7b+9nV/3tFRdoE4VA5cqGmeCPdvf
mdmJGvt5ex98Ph0Ee0ZmLuACcuZ/9r9NdR0N44Tf4Y4d/1kxDy4FqRKhs1/SlOew
Gh2s96QRkLVbTBkQem3GB6MyPTh6zYIbLa4zd+obrUnepIjPC7GYJ2T/D9gTOKEI
jor9zF03I0YUGMefB6Iq92GdFfTp3STJXy9BPlPcOxE6vIDJGRVDvQDq52SUR4G+
uYHK+3ZOYcNBltIcw8PBszs2jOaQpzZuOOhW/h1tyWhM9Gqa2N8/VctDN3U1VLxc
IfgwdlfWai4UCx2NhIl8M5pzwP3EOAjp0WuhzpYHY829FVZ6iFyCZ6EI5lpsw2iJ
wDCgdUisWCeGmKluQrwQOtYUsX25ZMBpb9Zgj/NLHdu74dzIXpDYm2UL8jcsWEhV
iZfxoBc6RzpTwhjkDHECEDUgnB2vq4zDlmVrgW3gu3N5iLXcMu1Zzbo4aSCsEwma
pH1U7vt7oPFll+lwYMR4Ir/iMpu+EtDGO9uGCi36df04ZUniEt1KgbnTK3kDYPzc
JwPr91tYDSAMrbK6524e4Iyr3k4dxvRYjvjrzd64nn3pv6h9B+rk3xVG2uEmivzD
pG7ZvRWNKhOWXiBMN8Nc/BOWuBrXNYteP2WKOcR8jfy0LcK5L3ekn0Y1GHhehE5V
LJujWih8pwpHpTfk09AvMOQZmY2dFVrQDZysuHqHXwrobWiDWSX2/DuezoP+gDxD
r1xNuxtm3FpABTlErngkuW1sRLis99Rd+GJiWB+D7auhUY11juNMvmMYpXcR/uXf
BTucPnz3nCD7105iTjPEgYoh6WqTqYdlqdiWsVVPYBcw/kAIi6J+ayXiYpfFHAUV
yFLX/GBkah/fWE5uPVXitRnxBd5fJLC746le8hJPM4+wsAl3seCmwCrjuu2SenoT
9Ztsaua+2rJNyYDQerRfCr38tCfpdyIABOTs74e13AeJB8Cl1cYTKFRfgz8lU1c2
/LCRKumfBbcsJOxjXL5MPhclhDUgmDPkqrku7gZ3UOelJX05qXrlHumxugmly9RB
tEPCaDCqP7rjflewARSmvjT3tfgB8bH/nUaTiH3cnNrwwJuAB7XEvjetsJ1g/57b
aLIC7vft05qw1Cq6FVSexyQm16Nu25BsbdWz483gBfoljgBVEtTN/113rM87DI1o
8gGYHhnpFcduXxfZT7LjjfJfrdTxbj++9ot9t8SfmxQ3SvDI8jBPJxgbezC5wxrW
KNmmey8/DuIBn6di0aQvVYWxPxlTFn13YVdnkBv/xcLI1kO+WoxtX3OjHacjYmUO
4C6ues5lNnu1eD3uvFyvjbyvK+0BC3uqf4AnxbOFYnDq5XyaKz1PLZe+d5JtaBEx
8hEdAWtQY29OXzNbz+l+OeJC7Ysx9/sglxG4xCgQhlmrsd7q3PYWk53vSzf59Qkc
b7G+bMbhXgT69uKOvCd7eS0AG7fF5OD424Ge59/gbOop9Y7fl3fZTOyM2PECCMaJ
lNmBGqisB7m54N6JE6gCB4DIvL/PoofuQQl+9cfo6uAKeRnjCY9+hSSRpVBC/j0d
wmleN7InynLZsbiSLMoi6Iv+HbJnQPLtYL2urX/ypbiWBDaNaY4RKJsDKvxDuAQM
JvoBhiG5YOnXKvFcYxUetT2LNZQfybYBr7HmMEeno74bLQVYriDjDcQD4G3jwfsa
20RpEDiXUC030exODO14zhCF48+LgCFUTVJ+6vTQ6388dWxCbG8fX/GN78DAT3A5
WOR7eRoQgyKcuOpUFPXJMmdbI3ijI2F0Eo1a4tgA8nhR36+W/7LKgqarm0REglfl
Vdme3UMZwnYHpvF5MC5lrCLHcyYwe9o9ZWDzSX/Fl2FIaS3JO3r02WC6GrVN0v4j
9UBuArDxLI0S1JFnZ9UPMyxSzhbkY2dFEOPIgW4wK4jU4Fo4H0KW2PgW5h24OkW9
0OO9lATDVhYF7gkcP8/mD2k08ELxU6U8KSic2q4UFXxy7c7s25mIRGl2t98FzOYs
7UDexVrzbS8eQVukSDE6uYzzoB7Ud88k7kHbiyfDerE5vRfL7Ye64UgQX6Cg7zAE
WHAsHXMzqH4UalFB0ol4zcCgiaN5o4KHNTafAyGf/NDrcY8YzJPf6pPgrIMrlXUy
nL6HvGal2ED46AJwXA2o+S3Gr9Sm/crCu+mSVpYD7f9v3G6Jvrh1GH7uIV2aFoqw
WduHYbbbKNc5tQrYJJmRL/yAQ+wdiptL7n4LGsB5jvtR55dqbpYtpqkh1YdM/1kd
HgjRHcA14r570CouIRVMlc87XIwSrUahfP8U1bQVTDligthJYFuvqiUg1X86/vJb
7r37uN0gy8kv0C7msqTu99kPNgGU2ur3n1bbdQ5j+9wRqItT7AnH6Jg0wFNRFovj
myaZOGVzeKvrL9XKDvph9wqiQw9GOswunHA1a+VZJUxfrsIZs9ZGHYAf0wRgL13b
6oxJdpgdFTBZLiY6UAy55jCKYHzNpjnhc/jiB7cD7GqxRPHPAJ6W90SfXLQpJelO
opKTlaNv6mCjGvMI44+T6Q+F0a9wdrRcMY/FZ+wwKqt8MPTZLUILAafjkD9GNHsd
pBBNzeo9i9zE7Ake/4I2/+G/UEZVQp9ZYBLMKqMv7us8v9GvK+CydxrcS/WTCBNA
AO7+v6yYUzXcP5SBb0Pf5SHNvPAIoWWq5TR/4lgdAZGpTqX+pK93/4esUuAbyWb7
KWH9aZBPVkIyWXzKUqx5yezgMOA+hyR+FKRgEf4NRZ6vdBIajRhq2GeR1PJSybcE
YTIGjaqnAzHdV6cYWVriwVIKzn+/wuxFw9aRkazMzxxmJLTEyeYtlgOQ1URZ1nmN
VFlcdqwr3G+p3T12sr9Q5mmAO3caaW11j1nQsVW5C9J9xcAyeBMyiCw/Yqimohxx
UaXnZUnTi4PfeTqkVNBVZcH5wLumF5xkfySYZBMHhGFVrvZCL60IxmPf5DbU2mF0
kblOjQIxOAL+Va537OR8WUqPTictLlCk61tVhhJPgKK4ciNyEVN80Q5juvlTJ5Fq
Y0r7G8yw9INVzYtFINmGyfVoNMLfeD4+KpNsCd812ASK1Gsjc/KGLrvi0CV1qEYI
nABQoabfble7GWD9WFJ66kSgTwLZkvjW8QGmVPgJwAYCARcArh+fybh0+p8Gp8yC
BkeUwo/YLltbouwFvrPW71aQ3kYj2pbyyZLuNv8sRA86kSrliGRGacMQr1rLE1HU
84i/wyAX0j/SmF/SpSMPpUwUV0kluLg9UNCwpTdoDMQwwoQY52SBn9IUdlu59EYQ
C4bJv3McaxgRXOS2/AGT+gy+s++h/O7ylnfOzGSRaLQaqyQGClxFZrlLzo49e+Yv
wxqEtlembcQ0kePMw+nTRxBMYbLwXigvWg92dsSzDM8xBezfnMaRVMFRqs7AKat6
bdVT7e19IqW9axTXsf72t6QsM3i/4iIw/4cjDYle2RXVnBziF7HCR3FYdchqfF/U
XDME9m+Sh1Mdtf1nfAZ/ei8OhvAHFzIbeWqCwglfbMCuY4KDmyNvS13UKJ32nzBc
+6q4pDYNkxsoe9sxjQzLQEsDQ5mKjfq/mnAZj2xWoXLKb46widqFRLlaVWJFGsEQ
KQU8sqnFO9X5baGUIex34yKGIDLvk47I+MlHf1amX3dIIiZDqYugAq/4pM68hcSK
EBKBIevVpkQFFCEd64PyvNSjrJFdsFJrXn5ZXE8MQdW1QwX0Qwjb0t7tMXdqsDnm
YOcWiKemNt1spn20iPunqnOowHbQzIO92rRXFsuyyNPzjks70eO90xswiLI6/66x
dvu6hPqCiEXymeGwobpByAtqKeDpV0E4BlzeQo9dL7G3OfsLFPn37tta1Zpj6m9C
lmCrJGF3I17DA9Fxmw9eUGZ/BVuNQBcWRS7lcTnCR18Bw8M8hpGqOnukkDCZisCo
gWs5OvlV1sxOS7kxE14edskCWH/Lg49TqdC5FB3xI+X4/FPPh4cFEdH3v3bmP+ai
+s1m6ExGzy2uB/f3yD7e3ApFybXBhAXRzSpYo0WBAJZJ9TFeW0epL22DSuMR+9fT
K/VVO+myCubgl7xBUAK8U4qew7AE8ASuqu1PpR2EjlwT+ajVeD/pk2RXlvLbkMTC
3OIL4oGGtsiqDincr5We/0eXH0y8ueIYOaHSFOEsP1JlqUe7FtBEdPIFuBqltIvL
LKz0E1NLOR/PkjUwXTRcWoVA6m1Z+PAqIDLbcpPDlg60+Ap49YK3p/hHX4y+Xdls
PCP+JNOzaaP3m2idHRob3npKZLYhnJ7gcvs4MHkaiSMFn90Zd3CDZh39jbzruYEp
koa5JpyfJ5qlNqPH5Pv7xmmm1w9tYH4qPipfwcO+44gxyY8nT+NhZ9Xp/qp7PRn2
2ovTWBbeFwlcHVUTMGoqAK47L2qqpeK/uN0oU2cbyCI26YpC6fpqza/Hq//mISNw
ye5HJwrLMzDUYfxMUIAoaP83daV3dd9t4jC0rlPQhyZ2kZccGrQkg2/NPSKAIFfd
dR/7hzhe5M/WVGzu3iFv9qAQxWjzWQdabFkMu6ybNiuhF66wifW1B1AxptntN0Ub
Ta709pSVTQLc/oWutxBjhKhZ5rsMns8P8uAF10qO2C3Y5Ks58WxpTZspnE64uPlV
7Ply44QPsGuv0PdoCxl4DZvIXgBZV8T6Dly1LXNg0o3dpgH6BI7rcHVqObc89jTm
nXM076NbHZcteetRgvjgX8PkCb4NDM+31q2G1AoFS/IpehXqwpdZ5ci0PdoYh9eU
sIirwtYE6AJepdTyTDxZRqtApG9kB7Xq/2+Zy7wDUU3LGGMIrJXVCa+WC9eKtLy0
SwSFbMwf32IVWhV188jjTqJUNB6yPldJOi7tasK6051py+TETv9U7Hp1i86GsovK
HNxKNIqBk36Nc1dBpGhl8C9xZcG5vH1QPUsp1CBlhwj5MrKbhzaepqaBM/olEUMV
C8dR1/8q9a4hgKy6KhsQ5XXDrNk1NbM1YVUs2gJAbHgBeI8T+HBzTnwFOPsItpw6
DWIPPnQwV51tXm/T0YJ/mgGUb3fgd7thdP2qvzndJjvj6xMzeaZ7NoszotRLGUlr
uTMO1pFBewDhoQn8cmW4C6gx175Zm5EUn23MP/3FqAFhuNTZqvydz1pUW1CZdJWb
nux4StMquYY05juOhPIiYVbXQ4v+1o0qt2ZT4Vqv+XHcHHZ8X3O6Q58M3oylXd9n
MtBJzHi2+XZ6GL7l6gZxUUzgAX+Ye3AMqpYMpCYTtDoZAQHldA6ArIxjOQ1m5TO2
R2dDKZ6vyVR/qig+HOzcRK7q793t9S8o/Icp5SVc908bIbrxsAYUzk084lKl2o8W
SMwXjEigl46v9IU9UabhhhfT4CQ3ehfLRz4NNjLkZGl/s/m2btfpqSPsxhK659uR
9HuAfxK25iXIcNR4gQVpb7OyMQiNX9yk5FRtXckmi/sislebmKy1LEl+Nc3VXv7/
7ZBDf4Nm6h3khSuf8r5C6h5bpFSHerxu68C+4m8NbA/P0gzLA8g8ifefwBgYwEtG
Q1yhGDkvZGxd8grzK/x28Twv4Xa58vwacYd/ApD7A7tYznSW3xU0CN7A0bdpysYf
mnz0SrMwiS1s807ssNFS5cpUTlaMU2Nbpc4id7O+7sVHMS4HDWfLTXdLCKv6K623
mM7TimOZI3q1r8r4OLFCJfo77H//53qsJLHGhJ183UY9+x+FJ3/z7ffD9vrCWRhS
Jx3KyBBZBLz4j6veSeauQkM7x0MIGhtRdKe5P77zUtnxAXBxkugTXkkRE/6d+LJa
4kxCuOdkbXLzSoKid8jHFkhrwspy/hRvJEXP8YNDUjAJZCS+ZKTMSocNk1laHzia
wdBcpe2oXQKK8Y0ExYusABlKYnn6+9Eu2wEo4ck2hNOa28MuQmUPzdaXJsGMGWnt
SKn9NHm6gxZYjl/myXNT/oCRXZvVqY4zHIjxC+QMlncw0VLJn+qGbsk6dnK1HHG/
lm4nYXegSnB4Uy2lbLvh7e5R/UyeUPE94TwChUjPxXPTyNUVjDknyuWp6r5tb0bc
zlX7WbTzQSoRQf5ibIpSxdq1w/OsbsDMngueQpQZrhEJez2GWeK4UvDLfS/p6lK8
PeyTTkjqsOgZrnX+Yfb5Y0cRzj2nQcMUH3gk8RkgLdImbHSp+YBTLJSciqUK89k8
wrhtELI0qBhFXenftqdcV4LaiKU/AE/2DckW4NbfM9JNUqdVg81tiuWCA/K1J3zJ
2LHOoEle/ijOyuXFCtZ4lR8y015YTJ69WvhBqBtAGSnE7k+DR3zbeFVx1R6yS1qH
3zxEfbk8KMqk2bPSjS49y9M18tVjW+CHae6WCj234f8ijwQ6EwsjrlvYJp2f+COF
L5f/UbWotZhpW/3l4pXrg8zO9HnqqaLBqg9rBbp0Hh9xuEg2hpGK7JMJrym+ObQI
KocForliezfrLXKuh2XA5qHLsil2qwtdjLcBK9umvWwD4lm8gSnr7j5Ezq1ZxUVP
YijZLT5MdAREhSJTxld1cmDszjo4xxd9icCzMzvOmbTASCnkWys26UjPbi6h3cLI
HpQ3B/9DVXluboxW8REqnTFEikqsL3NFhX0SwC3HiE0qvU2LFXg1kjbpUDim+M77
crDdHQxPHng9GO6/SK4ti0cwru2n1uPkpzc72x5eKFblwJuJA5JnaUrzlBU37oo+
RrQ7C69II23SeIL3TXOUoo1fHd9MgiQutfQSl50W8LphjPMjDOaxFyAguvDTktMb
3mVja+accGdlecbvmrwJLnJHc8euTH9PkJpizDuoWhgctUt8T7uxeho8OOxDv/OB
eTHm9a2LEuD1P2G/RFWmLQEpvD6jsGd/UzlnnKKKLq9DtX+FWEDBtAZxghfxM3kp
ghOf4pH7cf/ecnnk9kqWRa0RWietbhu6G/C927qc7Hp/UUG27FAwW2Sijn9vI12/
piu/P8JfdvPMFtYDd9SidCKhemYuKQ574HFMC9M7lFJBn9JYXyZc+IZrtDiO0qd9
UjlRsKS/q9olXzbh7y7e2jKNf3YO1pvSkEhUKGSzdzcsn/PTA1CsNDPuxHAiSSBl
b9zGvlZCt5DPMwR6yvecWl4VcTBF26CeUB1iDT52XUxayLH2e6UcietgAhDCipOS
0pvsECe77cGluUQA5LMRcDaWc9JWNptI/ewAH0Usk0DyMINh5WTh1DZUfnGKTad1
2rr5VE3G4UVziZwBDFT3HYts1LwT/iAbUyWtO9hSdaohpVD1Hfc80dtjmCR2oqSh
UBwjETFDqA+5h5DDmsdVRLHOhZUKY8pWXCCUE2UzSOwCbdpVJYsET+7E9kAUEyIV
JfZlr86Gd+gNbEQTRdqaco13v6voVf814U9XynXZEUoCFqqQzQvy145pChKpfLsp
pkQyvM6+J34Fn4wg9doUtxbo71h1QJMmYg8+GbDftEybzKOOhdY5jMpPPZ7Mov9D
A8lBCGz6RESKKbblaz1ofdiRhj9T5YzOUXLptAXwV1LwJPS8aU7AF+i1Ln9LlLrS
rOA4vqoN9WvErClIRWZ3GpSioc4Ky6h4o9l4YFfxsGE9ZEggSG8aXsL9u3N7y1p9
PxQJdGuLAECNpvdybfXK3nafQn0j4YSrIKZ1EmMO+AG9XKuQ2SRVqD/N0UL9nWqq
Uil5lsqG7JIpF/leM6lNIr+taE11qABU6kvpHyKHAqJQlIFct71S8DWDb2y15+d0
4fm7OyqfduVAz0xEeHkw4ssproEml8xiF8/8yY2QAbV0IbDHGk3hcY8UcEH93A3b
ZQSEYdupvFeeIplaJW+jYkQ/6p/6BaW4mIORS9kzZ3AGxaowgLHmiGuy+bjkOPwI
H7fKjuksLv7w9/twMv4SUQ0n18jT1Ems/Wcaev3E4q/UR9hE6i4D5zqv8Qy3uBvl
vJ+aocACrpeW0ynlz59oYgOPQx9w7pPPsD0MjrnLqnKa11BpWRd57jsCmcvHP0SD
U29FTLW0qcZawxVko8y4e5BYtqW8TMdvJuzOCUOzLG2hgSzvcr9uOcydgHunvf9f
qP0nTIvnU2g32F8ePUINwilaKcLdmoc+oiYM5h1R46cGMRfjNW/28MRemUAbU8YS
Zzvx678O5LqsDDWTKMsr5ryagmNOCGnafM7ysTVXn1mYUQLCGJ3WPsO+QEwA5hOc
kfzy4Hx97aH42O/YaryLEWMsSl884dlrOf+O0p9LRj86HjqnAQudgNI+I6KvsOj+
s76gIe0hhNTj+A3NpLEBLgA+3an/5ipY0paHOWp8On4U4S66AGI0NDzRbfgzlqD/
TcPHCAYJb2XJ9JV6L14j9NGTAJjdj87OjnGgb1blaD6Qz/MZy5r3YnjlZeer0Nrt
Q+N9WNnysHXq2MoYzdfGdyC5tQphntwMlH8zOQDG32sKZyAyDX2dc1B38X4j1Ken
EcfjknUu6dYOZ1qM/wRxKrGUwsEozTVIJakx3iPPQTJTRxa8SdhKTLM9JEj42x/v
rfQkA2BQj2wyH0hSrcv9TUwCg5J/vvLf/sQxyJqlzAFoe96EaRLmCKCBYPP3VhTl
j5N0SJn1Be44H2sAQ11ybK55WCYL56mNntpTskVm33lraDiFsIfWPPlcIAVCmy0Y
Rq/YUkRfbVhKQeoILAjdanygED75vTMw6T+U+Y5UL1QouP+Q8TjtvceevvIiPMP+
hN52AMRdQPC/Vf5HvpVzOr66DWAZJ7z98U6oFfc2bb9NoStzhMfNjybPlLdKhpvN
vOrc8eBujc8CZbd6vXHgmsk4mB5BW8aBw0rsKqdmx80472ZnWe/6Wh9M+H7TKy+A
SEDdANTLkBQr8U1b6NdJV3ePVDmK3v4EmFjsig4HJyanLy+egJGVdlk53ZfO7KZU
KJ5fVhu/gFqJ7QWOHZ5C3bELFcnTGmgLfxsWMqDeFKCUddT3QHdGR5eFAzf9yF5J
6AgR6KF7urdp6oGbA/P7p1mDDZYZtTRpOM1bhJKcwdvEgRSCd/W26Qlj0MJM1lco
67rXR5S4I+0+N/QsM6o7sTqi8VM8f3WgzA8juzzig+VaDacjtrw840w6pfpSmzUy
PAsdr9vUGzenxp0g4SAnJQR6T7LAArkRGotPrJVkrZ7Vn1yxPhboq0Bxz7V962pq
t4zgqOBFTR6GYtdsmQGHxcrEpW86+mxmnaDmm70SAt4MprKsKyO11gx0miwCx969
Bw9O5t6qCY2V9HJtxEe7TxQg7BxHrRzfRZ+eK0eKsDd4DzPhxGvquJGIaMg7TJrR
iOqg8hxy4dFyYKBFDCHEBMT0dCnl9ENTZ0U8uEbmj1CIbTJW8S+LBPljE03cAfrA
igI9pdOW3YNOzOtzdVg3R3QNRjC4CdonWUeL+XP9zjwW2WODySW0NLFQVsjFczAp
Z5XEkC8wYvWM1bSSDQ+s23tu00YMPAgzotedpf68iSaaK4ZvCgAz8NMB/IVPufMO
F5fmUKRBC4uuXew0qH+PmPc6a8xCry8TjuOujRsY7BVLH9OZpJLyPnIVPWrzGcIl
nnOpgK3cqH4JSvlJWjdgWMThjzC1Dh+yp0JSHK9O5p5VDcSM3A5unqETccQcekHG
AKEqVGOxv0uBG+i4FH23ncTVKgIfisol7GAD1q4OU1T8S93jf0cRSlD86tmVBEdj
1C7ITJtNePRhVtSmD4uoqLuJAghIREYPUQiLxQ/4pxO8FfyzRyK8xQkJDImc9/hP
XuNG/G9Ppwtyp2q43eK8XZJSpqJe4p/Ni43IZv9es3kAUvwTR+Rj5MLryU5cM6xm
nyVHy/5YUS234Tn7htfzNp7qGUuYGi2kriEdR5NnBdrxs0thEnntSbhIBqp17I8i
5T0fb+03SHCAB5/iGbgOoBAwUXneJKAKxZLw2ud0C0WfzdyMpQaKDzatFu6RgcMT
NqKkJt1Ezx3fGtHnA8+et5wauBvZIT+mfxSbNWzwUz/OZSLAhXLXRHnzIZt7T/mv
+58u2wvCQcwoNXgtjiZVmz6OQBmSO03+Tmx1kXMUNCLzkr9jKdN2znoifGcG87rx
Z1WBWi9fIJjNvWfEmtLoNs+a6xBAnFCaBv+M4rbx4CxU5lNbGIs/2CyhaxlYFsjS
fXGFQkpSat+BJ/K3jXl5TKTMheKM4xkktUqJOfve60J8lcBqFYgpieyxlSfYKt/m
5cjrOkDkuvjep1cIZr/CdEdni297WrXeMUOWhnJCmzEOd406RD+UlFpfPg9AFdIZ
NUbSouhyKv1J13Xuqud2i2+AbwEgCeqGjn//vLKOVUkORuOMgOo6P/tM0XB98imQ
uPHm4nl/cRu7Z0oH0rhWiKaFd4fZl3+rmeMdxl6c1DI3/AH8eO9KfW8P/ErDJSEw
3g3zDJtd583VP6Ln/4zn5ygORlbfoSBrRxnylph5IkAj0jWkXkK4w7s+W3VtWnCM
pzlauOBB0Z2brm7CwpsUk3MuAs+LejOdDo2ozKQdcN9US6e3X9bR/CK+eiUHpY01
oKOA1MIYoClD+JFpbI/YmkP+IdoEWeiM9pz/AORGs4eFKbG0LDUXQkz7gQLcTBgx
sFQyJraD6NbhF7qIBLP59I5DOWVZHYbG5id29FEz6tPtuzEW8oyjF0ry4PGysEL7
+eMIVRs0Mxqh6kX4uX/atWxSL9VxSGM12dmuYVyQAufbtH4vJpNf1PIeqq7DJhbR
J0z0umAJJBl84dKpeI7XsZD9aZFb/ORlogyWJMsVE4hbzEbtt4w2F63wfh95qjsa
RPlQyDnQyiJN5QnE9BZcMWBH8MimAkQM6Ud9BhkM8kGEYyGiddcUhzs5ey20gwTN
2GOp/L0gCeFvTdFzL125CsurtlgTCyRp2chtDGHnWaOibPqj3LNxRfCn0h5tWNOK
/UqVtxcHHwu7+AA88HHodh/jx/eX/hDbM3itMz/exg6ylQIgXuMpHaL8muN3KS7l
jC+4JHaiJ1TnbvbftbO9vj2ChppmBuPaKRRyrxNwAOQ2xO39zvbgW57Tgs0Egfj8
dcy4H4NE506j4WYzE07zO7JBzi9DE0PqqyqvsQ9E7OtNCH0yqvlief8oYrmVLydT
ekvwG3zxsUiWqhLwTkAMOd7BWjiV8SUlI68+Cy60ZcmtoKY5TMYYxmIbxNIdfNa7
KT2MCRqsS82cgKmL7VqPyit0QVD+SExDYVxP5jRRB3PhOeAWrqegW940fjY3E9l+
iuEXty7IbzjJ3Ul7j15++TNHbpuDNqtsZCP75rCrBV17ZM10YokLqoAcx1LsmQCo
Zs+MSFQ6BpTKEMnjudE0QbhvsznXFLcsJ54w3CXywjIcEHcRA0dqVJ9CJIE/Nsk4
/DkXZI6OmlM9k5n+u9aXpksAj8T4KPxyOy0Kgii0LghrNnHAEpJhlKNS2pAqxmQ6
XEky7FSmqHbIioLqTCHjuVI1tnmCvERTqiYkb9O20Ms8mWG0mFnnKDWVuqRG5r9N
W3eVyOZquuLacyNCrYtK/H87xN/qy2Sm7aCN1pjq8xFXmvjlTqPjSZ/uXf6AB40z
C/+rCB4LnJTSdex0SchsKXlPCJ8+8EdM8Hhm9vvHr34Ff2J4Tdxw+Rn3Gl1b+egN
CYLP8EO+vL+RJ7pl0CL9mHBHFdY8tMGujVuanvHf3r9m28rLb3Tlyq/jVtpGy5dt
9zg7d4uZ7c1B3BoxPK1/iXuqkBtkfZbpPTuNNWDbifCuubsOKbz1WlMJxQQORkp7
LV+o5AX5X/wcjuAQGUm9f5DtnHWCLCcW4iuknBPe3u9n2S5+5r7OFoFQa86MQ5l/
BkXLdNMFJIhix5FbmYTBC5i41CCGLoO7UiKQ0LuUf0OcXRxkwZ22sAjdvm5UPW5r
uHOpvtZ6DIV4HWQ7VU99/3emGxId/Kna8K30KMSijG5acYAi0G/DzdesFtLNhmWj
vdyPusL2A2MP3KVfTRh+lny4Fh6z7E6+R+zaA3TYctKzSPXp7vqC2A4zZwHKo4UH
ovdx6RHWdBSOPrnwvrkIOlLcmaG+DnO+vcO/4yY+ACVs7GbXSZL/G+iMy5nOkCpi
N+85Lc94ltqQi145LP4EqGKnv4PIJPiS8iCYvFs6XZBbCfcukCvuM1eVgHq5ANNx
5jp+Ln6WVBQ4oDUpUsawD5Hp9n8Re8ZI8iTWPP/W0K6nvElD3GgvpmkPVpCP1m5L
TjT4VuAR22/F2EdKFv56AwCCxoBMShRm5tcErvV00rs7mQaf3QqE/Q2ksDvcdsJb
Fo+fV3ju2hLnuN+k0SGYVNB9P5/yCqoOrWq0vCx93qmyk8ygJmFl5i4ulmTeBRtv
HHByf6ibQ+new0XgUZHdvQgSn3nNJbbneEmIbfRSPdR7njgH5lti0h7CroXZN79n
RIlwuUaH6THofZbIHm2g0Su9jR7QWiDw0iSdenRgZc2MGDYtAb/I4mJc0K3PtgSQ
e9rOcD0RlsweJDUtU531+J7AzJvuGfL5K+LHfifytoVxfevTtA9nl79JLuNEpae8
FcqUmgWo8Fznb5eEieQ6a4HgxwfN0lwq992IHt37KE6NAk7XObTZntfUeHz9ciR4
0X9eBK6BTIeZk0Sv6Pa2viTnTfTzE8zbo1dufj4Dx4W8cBU+EF/ZTHh57+87pYKG
pXrQ+vccHX3hscHFIYOXHmRWKfvR8N7kYuk48xtHIGw6X6qlH/lScle4Yba4cV9O
Sj9r21iSX/5qAis+8FAle7o1L/xeVa3eJX2UjC5I76ZSXiupRPTOVjFQPaqejXY4
kjRG3ubnx2jvuU5Qt+f4SmRcz4LtMeqM6OhSC5E6CPkT8cDbIEn0O4cxtXr5+Zff
X9mPpUuyBgjEhGsU2FaWUnrMCRHBBGg+SqzDBVO21HLRM2ccc9xn6rATTaUOGRih
u0XjDgo/3hLdz6fOh7y6UwCCQ33UPf1MMMJIBIf6Ua8/zEIcm9v3hNaeMJO4tPkG
UHMOwXGIncUmhyLEN4kaJHSkYyyE3ClZuKtVZ3uhGlCYdZW28S/oYUqP1v1ibC0r
hNHzadxZ2mOmUHrw8Z1dtr6JbBwlZxzwot3Zk1nyfg/9va/zuMLRk9mn/8yFp+Ut
W5hoMMLbCZjnA1wiHI4oDqz0KAD8i/HOxG6hiNcdGedBUqobBromQFEpbsQkUobi
z5Ag8keVTSS53W5q7O5aoPHs4qvP0uvP9B2zT5bTP+ynV7kjW/5HrYnbu0nnoGZQ
SL1R02pB/B/lLVWxJypwk10a3Fm2J+R9SnYEeSTPpjdrXmexataiShpVLpl/y5BT
L3uRa2fyWdX8CMLdfjHIryvvT38jxr+N1xDrIrcypGxjCo10ZlmF5uDerl5iwgma
ZvuKzDVKen7iMRTOpwB1mbdOQrWZa1vbq79hC9N749ct8lxE6ioW7GsS/XqIw6Qy
8xPpA7Q6XCDPfmtBqUe3al5Z0LeYe4BHrwW64QnH7PS0ybs4rHl/Do32sOmsViI4
Nwl3zyULwD2klHW/Lzp6gasBj2a979SpgRH3uiNA8+HzUHkIiKlka/zpYLGCIXHA
zXaVUd/IyDPlcT8e0xLsDog7a6pRQWcMgDnMvrO6h4UMKB++AH8e0Y2xSD8SrOZc
kZ5PjzAykYLAfPBWy3GeR2n2Szv1nUe5y55kPeJ7Xs57TzYSy0VKVnY8QKHpIqNu
rQKeUPnvyaJ3QUDeZTDZH8PrZQeYfJi0DQYMpuydxejYHMlspf6CHUy/UdRW5n1D
XasEFRCDiK30wM8Qve/fuuH/IkQTzPHW2g8f5tM858R6rlqVQp8zwbm+xKI1ff6V
db4BkQeRnvKflxZmfesrnjKFQm1jUFr4K+rsBuFgwzh9nJwFRrEwfq/KW6OLEi0M
cgmlIKTTf5cI6iBkldKBn+/ouEcz17Z5MGpKO5mIIDaovcoGG17GMSDF5eGWLYJl
oxAcy1nINBkjLFAYoVwaoIev1vxz8PwawDCCTEdkZLCSCXMHf7mWeVOXEcPs7XAm
yGKdDPzggCJ2BO8AIyjoZy/3gp48fDr+HUCKli8TqRiamoC702swS6AkWw6sMFbO
nRfYFY+Fp/+0d9MZg/eO87CUUGyjstvk0SVbvBvPI3gQMxgC9n0eXwa4qiD4DCOX
bwIZRuTUQO5QxtwGWkRHAS3PBXCqOdK5K+PF26OkzKcn09y6VcUmOtFD+/Ymszol
mAHSv2hMsW5EmItx6gDtfNTNZs+Sl0ejSK3hl9aYSJGQXXTiEi5KUz13YyC77HHR
LuiXRh7lo6JqW456BVB8pStuftSEGPhmAgYwlaJ+g8fwIdSfv/GizfxQ2lEyW8Rt
NHq/qnX7CVTLdJokSsei+NfoDNcKHrkNBqzww557UHeG8ogD2R+rxSsRSSKqlp4U
egcujeQ8m2Ke4QGeGrp/eSDwgJj1OjKK/kl/aibJsGsaW75UH+z5qZr/wQc72lW8
b1gc7A7oVLDcHYXw3gfihYkxaI7fCy6zD7ZY9aktbDAN6LhnHTPxsRP5htE3n5KX
8QdM9tt7pxak+q5flSeS4Vrxt8jeod+38Q8UzSxP8yHpiiGiqwko6nzp0IszxMG7
8ogju9JozSCVnKUzIz64Cv/xn6MS2QpoFFP0IFmHwRvoZcv9tXbZ4XMEXUUZdAui
IvyUSVTv5oVToZnxaiv+CnSLW6gTiSTk/nDvvTFYbl6D/SEQ4nhBK4TDhHwbyOBZ
ok0WcBzj1+j9NnbXVVGzw8uSMMj/7fuYEv2i3Q3Fq2BpG1NcqpBtZseLgTX0SJh6
fIz9C1qh9L3l3b5W+Jny+3eAOro6kwZ+wwcd+kRNhw5v0FbWc9W2sHkvG8SF1LTw
apTs87Xs3Akatthmy9kH5Exmaewgz9HS78bPrEUhMJH4Mx9pViU+10+aB6MkYG2X
KBisaYW4/Xa/bi6quRJpKNkoHYNAd9QnAYsZAoMA7nQJMPd8qRd+JwVRqD+R8v6T
v1UxXGiXfBsbWz5L07CF+HYgixxDqCWLU2aVfjzuqsG9Wa6W1DUjEOCK3HuFtHcK
2reL7atUzRSjkoRQzBqseKtIehxf225FVf7/ajrSF7l2QYlyPmJAJvQ4X8NDJ7tX
trZKvk6OGptwhp0YlDfcNWixfd0Ycj96u+9VC1VfG9Jco9Wru8fnuP6C+yIM8oVO
qQj/cNU+0E/QARHUTRA5t5ohfCCNwqIyjxrOJOjtaU1OjtKxvZOOEq1A9e7mN5od
LjLXXuYGvz50HxcPEHSCm88L2fU1uyRx5pkOih65V/wWaEtFSVOllnDk+cNarWBs
UIWDELob5KS9zUf5yyDxuuVFVpxjtBWH8HM6CabGx6B3ok9IocfL9+lfw/P/vgK0
tSPgocW/GnPFmKKHGqlo8kGUJbQiRdsSM8FClLf5llvoeWsTivQoBiTWJyDu4u2a
mWBWSlPfu7RlZm7szpl/lH4DWdelGHE+Vh9dWNmLpFTdTEzg1CQHfubKcT+N9aVG
nnSBjnVNO83wJoHZahzWNnsjFGtEsTwHvVvCTebC95SpKZkKwjllvc9n66oJnRk/
Eb7kEN7SZPqEhXn37/wZkwo7ZoHH1O5I0HkdwzQzmfce2oKVDd77QWARUtLWMFDx
kbz5pJRqHoeV/0SApQOsbW1HIrbARydlXdRUqGagFg3PjMVjA8B7gvixKLPhVjzx
Qj615s1yEe3jeFrSC9NbF+wRY8GKmV0bPw5c/qZJ9kU/soQyrDrkXx9Xsq2dJ7og
q62ab0PiP53vQ2+tiysU9aQ5VTzrH+aoYtplyw6bVIpbnr+0Qb+bITHCvbiop04G
TQmwDP7g10WgqDlcUyQc9Oww0rryjOXEP9lyWRBP9t/zckmsDCH09RCXl5t+ICBc
1pYZuRtRRbLNG6KUojERp3aHRHTPmIielaDtbWopvHhn32u7nNoOHLa5ArujL5Qf
GYkSm1pdYAqs2kAEBNoLoKop6+HUUHXBSeHzdV+U8pOLFhWjpKHFTtXj2RvVU1w0
K4L6pG6rxwhthJ4/9FozVFuJpMV4ZOWamQcV0qrxXUtCLkrxDIpzbfth+2+CYr9q
GCHy0//szW4SyvUIBUEdYfkJeNkjdBd6v1cOC1BC9gSShKpLEsZXZJDuvPOQn8RV
u8LodAeH9Utj51CR8z+LEekQP237G4aIFnfeEWuhRxtOmffA4GBWrHYzX5UhqSnF
G4XtRbos66Yw6YjLERhDa9fb3QQ4Mv820WjflPB9tSe6aoUjtUruLNqQx7wEBtwP
B+/4Otuv1yFrgo9CcGwpaafolNqvjRSnoSs//Z3hc7d/RWXJsXwne5BVp/gVsKR3
82fi6jNiQPYxiUgm2r1OyyIwnMLcCNXZSDTEPEAgSE2cAe2nrn7CfvYM8R0A2i1j
fY3z/0hESlqHiK6WLCC0Solgoguvp6qPHM47WdPtG6Ofv51f1UtJBhUHtCj9TRTZ
b5XgZQ1vvKjc7hPgqnFVBvLMuB6b0D0pbiuZCw24at2XNjWiz4pGx+/dmUmpZ+zZ
SeR0SsDbyz5eOXF/Od+mkbFBa7dSrYH9ovnCrTTIJ0UNrR5eoKgfc4DwCdPITDFu
pxddWSgJB+Dv3r7T/vqXCQEq2ddDGagXPvA/jcg/4haPmLut7WgYnH2gE6+8lpyW
u+lqrMnAoFw+kdpTqYx4YVs1DEHm73Ja9POvPdi+lftHEDqpa1nqjLknCca6KFjv
Y429GX8zrgmdC7LNlC6VWpCl/EXn4eXHkyO2RvSniF9taDT0tV54zAYwt7tg+Wxu
MlKxgjqEykK32YuHjm4pIMco5df9tuwYiATOay7zotGMtwl5X7VZwVSETWIelYas
re9kF5N9TNnM2lB+bVvetW+BuayfhHgJk8sOoJ7tTTm7Y7iU5ayHmUJ5xhHKZu7Y
var4AnuuAl6pkFtCzfo2l5zH5pKXboolz+ZVInfipAzVUDM7udDXcNOFnwi+kvnh
DIZxfsY2XC6vXyQvhhw/FbGw+cg4teDo8wriZxVCH9UYTREAmxB99pHPi9i4UYwW
exPsgLVQqVyhekJqTI4AJR4ev81iNOi15CgqCSavO8zha5JZrTzet3leUft/cdUd
lQxlef0ip6hannwFYAUVY1ZRM0PJHaeyEfynV5IOiVY7LfEU+9KHydduPdBSauiI
pj4jF6uVaensfupt2pVMRTNeC/EtEMurq8cPsj4AWboKXjUt2r9IqfwrltoYHspr
VR2QgGnhVUtDrDiesUTZb1PMCMVPQhNYtnSxdryTM0dSOHuaiOa0AdWSWCnh4dFn
lIKoPCZXFx6+lfaiGoC8+frRCMLI3UOYbxKc5p/QI8iMFxOBCCAbM2qtCIHSUYRs
54nfXwTBbMkWFD4HtIE1FPmkYDV8GT8wn0Q0wXsMqFMnRK6VpE1JRIA5AenSq65f
QFbhUngpeq6pwnknXCDYz5QgQ5WBcTGL1GkqlVIi1dKs2MQPm9LZ8GmhvY6e4+rq
BVVhzdrWoFFfmYeMBYJnQyA7YwTl81QQSQqNJhJX3MNX98MhUEdu4i7XR0+r8EwQ
DLyj6Rf6cYhEMifQQltzhRX67GCqpqOlBVE6GjpR54CX3Zd7yEISV0EYKLwbBUSX
biMDFCYDewGgK/WvwrEFRiJwLEDT3Ky7BJcqD91b+uG/YgohNKUcZ15Ei8g2SD0H
7k1/BCMvq3JI6ryQkjeSQkm2hSAdVHTgUN3mr/rmBGG/C02TFo0Lm5rpGfiE0Btt
6GZ/3F43Vlm1BgNYM75FUyvWPs0C1Is6i7BzZR2Gjqgn/A1eKUbVIpoFSkZNqnPu
nmuZGPCYwUElO8WBtrdow2wfckdQJDt1fDOKo82kQW1PaH2axts5A2I6IA3ufZ9E
woiliT9EArzHEpSkMs6p8QwGG3athzJ8PuRrDHKtS0LaY/vaJoGC5ZNMywpHv4r2
31gyUMMuJF2Moln35er10EBO42ieRDzf88NJ3w2X0uYQDUk/B7VVJIXaoSu074dE
T1EzMPeWEfDivvDfCPI4c0FlhVpY9ww3MW9oJllfaAlHJj4hkrZxlBgH3qAApMM/
u57ncGghCNmh6lVZq8sY27Vtx6injPOqDUOAKhOmltpjHapp9iOl92+q3kQltjz4
G4cOoN+52J7Qp4cjl6PEihTEJLr1miYT8mw4lkT/3WeXjbLO4UEA+z59i5Z1Kw1r
S4dinD/5Ohnmrze5tm/PKoTHPeo3lB3zglg2OzG1Yfaad2DRO7tll+jgLKN3smn1
z1WtaCFSBPPZ+sK+uXzYsv0kH00wBEvZGcGUhUiJkVn8ZySVWjYDy3e/XPm4QKi7
u0d1lTHary2OxCdqfjNW3pJ8XiDYFUD/UPQAxbts3s0xN6onLxcg6yuBP9D8ac9r
EWZ1KwxqzGyY03hmqXIkYeOn6hoIW2izCFGIQ0VvT8SvjpCUZmlzhfk9uEeKGwcs
2HIdUhABiW51RA2xZFUx2SOoYZFVTRk49F3X+sAkNKZhrbCKoCwwZ6Ek2eW1fUVR
mU4YjTrkobXn2U5ZNqsPlBwVmoKUpoN9V4YrVK6Ka4FMAedbYQQAyA4597e36/ze
lM/lRpmHCAk2tg/PGP2mrW//egNFCKnYWq+FKslffEzcjH9DVGKJj0vJDf6reo4K
GvDo6WYJ/8BAcdHb9kmLGsQJ7qvcitYOj6v8YAEB3+nr2eP7Ja3n3iyRf/1QvtNF
mPn1IcTWr86XhBRwjSDmPiaQb/7L12lm240Crp/pC6q1zBQaW9DElBxIthkTgnWi
LrfPJpmlzGxTPkpgfw6SuKVbJJm67cjmO1ZJy+2IviHQrsU0fnJIL03zSzftPYiA
U9bANI2MMgmEeJkbKweb4h564VVhex9uKcnECsnWz5+lwZl9HfJSgc5XwwrTy1QU
pVagSCJYqHf/lR8msbRiNUTzyntowaD710wXS/dfwiSkstHlJWpqysufrKrvaukD
Sk8lefzAWIR721uUUp1P9zguT7RDEbqUbngzcMXfB9GTxCDieCD6Ib+KNS/wYWl1
Moq82P2txhfpwweq48SrnNnU6zSPrrOy9SnkFdqNggjnTMdB27FUryvaP8HttDpm
oX4E2xfveR7tvBuEELkLhUpqzYYby+L9Ryp6XbGdU506yf+aPlXftzUT4/bjwJrF
XRq6st8+E2HpikP302E53K5G+QCn2xp++vl6sjaGa+HB7a96su99AEChdE88FRPH
beXCh4NQe1JTgH5ogF/ho7d3jc8Ryhu0E+nbrPe1Oh3ONklSrYCFl4O6QFsUtt+2
sFh+ygAaaLPVFYBCl3xZRADaBwY2pJbKNQDNzsruDq3f/QB1mRP6ZBnhRKEDeYRc
pZmbLzHEWKVzBtiT5yOnoOzLA5Hoyj7QfhW2xdmNx9TAfgQGw5feQTptS/eLOMda
xtFSyJKJxzME9vyVh5GUOi91rKoiFNBm0eRbqze3YB16S0yjWSY0k6v734S3hN8q
W2N/0pmQDs33Bf7FoVMhIA5pTAEuPkV/UIi3JPznrSAMh2ZdC++KrDRMWpnlqQFI
ckWw8h+YkdXJ0GsPB1cIrBVKTvj2oH/A+I2snIrQ2ZMmJaeSrTkr4kXeGPgLkiJx
Tml5kRKYy82tyEs4euA7mk8WOeXj0vimitEcW1b+QeOEVOW3u64rGusMf82/YREf
GaSI5HJ+Wdq7QseUII/fqTyrlrIeQTvcNFmy8XhlsSoxbkS2d94mTkZTzRCE5VYk
OIvZec9KaOm5z2HvrlrCcFr+PIJ79ubqjzLM6Nd6q5oDnNktl+snFzyJUApfFsFy
eOFRydr50ronfNiuI6ZO1RaCtFXmdWXkCkj6ChCl04d26HVfGT2M39CJ0iaqCl0w
l8jZPeFAZe5JA/Lgwd62ieLzpfeSbP8fv8z+RO5mkYJWagiMQn9PVs0vlI1bSfx7
aaYAA0jJBbkb9TWYDnoiv1XKboelnKbc8mhjIPtXi7C8kXP0/mQFq5HYHagsG7Yz
bD5ktEGTVXvBaAtE0BcWs6uNUYSv9lkElfX4Cq6GVduzvq2MbPoSxOfYk+k8JvWl
SV8yC9E/2X2L7U6DVMDzaIhDmmpPWveD8wR5RgomvDKOoMmlDPfHHFEg5Ag0tlC+
sYyTY+gc7s76jB4fa9XfcyUGj/f/CqcGPcTvu/VCxPK/Dg7szvDgmG4B1+JZfU3U
OaA//MgdByxTd7nKnNZ2UV9ijTAR32WwKFWLHVdHa0aZZSGOcZac0pga+DcnQbML
bxEn2wOn1oxG+ZNd1ynx1hNSyY7KHY1fHWBS0j7nI2TZfOA7sHU9GOxjf1yYrxb9
3L7aF1WPWImwFB9yaptqSPfECvastjZ8EWOmtIXHrkL7S972cSCuXX67hfd2+z39
i2q8xNAPT7TRQtVLF7XYb4Z2eOwEnP8CzCbEibv4AONGXqp29FJuDVmrGe/O+YtO
v7s2Qzi1iFIHqO2tQu7gQpDo3Gmn+51IaAIUbuWicYDtGypGnVhkUExVxIq8FyiL
pQhZ6d7lI+1pNQztS0PPH7V/Iut8mRWRsKGHsVVVJM297gv1OV6KPdY5450TTuWl
XkKlDYkFSuVv3LWYS7ny+O2ucvos8faz3GTCkLdrV2UvcDSRk9pP5nvPa1E1XWBC
2d9KK0iIHwGRktSPS0nUx3LUNQbCeyIU/CVXyDQi9JqEpbzSoUEGqUnRiVYWLst7
75FNP1cIRePRZ6wiT0Ll5wv30JQcnaG4JqyYNlPMsxB1PGFiIKnbWxrHNfTda/q7
U7awbqlfRYSPmf7lKw9wicaiIIw//7rEVQcjTYzCjLqe2dsCoPrDPCJEiRSn3F+k
WTC/WppVQY02Qss80datM2PfTHN7c4j6K9azBfFy2ttUExcf6Aj89s7VOuPBxBin
gIsupxmdpp9QoUJRT/PWw0qQx5AWeBOalidYubkbDsu6FxtHo/82TBM38dad6ypB
S/Umwav85qq6rrOmBdUF0Mk6juhMAU/61RPFoGDKO3Gpr+7U6+7cpa6lK5XxDGMt
28lwFR3nUuk28klDOmYhMxsU+EQ46FElxZe1rAGw9Y66SecqomR4LlzSImokQBYd
y+QmSCMHHwSfSi4EMyRhi7AYVD0xLUPvNnEwO6id/cxkuQLdkIDOvMpbUiEuK4YV
QhTBdT1EMnc3W67WbBCNpkUJTHj9fOhj5guDwEtvIf3Ycgd2Lj0C1K+rw88JRT/y
Q6gVAQJrTpTLPG32rwUm71dCq81T9oDMPctzdGEkP7KgZmG0Z1boaWQ0PuCqRqFA
nSb+0vZLngDnXz8qTvdsaSq3DThteVC/WewmPJ3XRl8VbDcCiY6hdqXrwRqaVXor
5EjnQjyGvmEWVnBx7tIoSGwVLOc8xsviVC7r3WaF4MaakCJR/bkwc5hqDsCXBzAg
IPvTr5oA8mIYKaxHxHnOgCGFXujQ7Jz80fiFzsF6nth5ObpbFdxNMPvX42zKxmHt
j/+IspcklXoxRziaQ5opEL0AJ35ZgwV8rNLA3p7U1VhfvhxnZ6ggCItYDdyRzDP9
OYEw1cB5YqIDKmXfMWiEHAH1eNHeM7BlUZ6EQC/yGZVXk34W3WiJ8r+Y2QV8y0c7
PDyHVY4YWgimZOgnuND9x0TN6+D2n7HQwHLAsnEjeTTVYyLP9Q57Sz48MCrQCs1u
hyNjXRQFCwCpqxfmgx5u/ZNlUvDg7rTMQMSxE8u6xZBlsLGfhhbrgkCXzcjbY7B7
+iGwt71K2n570U0YTVY5fiGN7SRlXNeekHz4PafOx0JalXm5KyfCP7mYROyYQ/6L
CZrNU2z29uKQGwmjaUTVn0LPZ8413xKQHYJUOaNQJxbE5rX4uBB50oZfmjLHqyHS
LKvh3u9xzxAdif8/gZW82JZdrqUlYz6pWQBT7aLhoXBThdwFMoEe2gqzoWI1IFYj
0tPdCs+5x2VBoi5RGhKxyVo7USFPXEq7RHXiKzd/mbAydYIKaynicq7wX4VvnQSh
XSQgMKFQedWSy9o3RqjYiqFIgtOsubq2tDnfeb8bPBPe4gjfWqWWDPyS5r0h7bBw
Igu0zr/X0rKQh4h9wFlxVaHKdwVX52mhErD4E5+M8ZKyb+FGLEEWrmXrTXyxtTvh
LDda2/YFPVHDBp7yEEsXLpxQj4SaaKIKiDEr1AQ8cSUl3K7UNsAtjG/FUrd9wzED
qHT6fileiwwEB9XliTuT2yOQl28q3uKLQMmFZqYQFU/VQ7jEChfCUQf2kVI/Q+9x
ajRCO+ZX4Cut1Cc4c7WeIAprUPTTRZLsEfNEE9I4z5wJM0Pb0drcVlMDzEe5KKNn
72rc0CBCioMUrQbO0uif77K9bKDkAYbRPZOeaFmDxp+GygyvRvrdefMSFn5iLfpl
4C+gNlvFPyWPSMN2b3MMSzLgtEqX8PxGo3frifVGDplOWeWmC6HYcuAX3H9oHkdn
z1eWlxNVqt1KJUh1XAURWJG10ht8CX1Imohh5oQTGJBV5mI/00DIo5359u9NKqXL
mljjXxnMl2s+Zkr4czXUfz/qanbRJlGapRAi3JLy0n/ecFcdIh6MW/o9FsRqZ1lg
8CLbLhoPzOBfhHWgWQnB8LrAz/loxpvZRmToA1y5THZMp3qMKgfCG2cpJ3E4/dbp
b8sQDO5gUuBNgn8ZGwVqjdlijtI7jBPz5IU/z0DZke0DhZxh9bYKmEjNzIGr+/1R
75G2rVV2ZUJGxsdb12Ai65Q98kkohSoIUWU6roLXk9NFKIMOELk8hvL1jOD5BLxi
IRb8fWOxoEaYSANuqAkeqTsQ92oJCpFwG8OcgV6gYyZeX6Z2OJWcqWJHf3ox53+w
tTFHFCoyj4cJqGbn8W6wDyf7zuzbs/j3mK9yL6j3szvPe29KMRWjgg/nDnlXdluo
mHcnyEHd5dble+cq9GDmRgw/PHRS3tEbbhgc8/QJWnE6LglD6FiRsJqRMMelAhq/
2sAbsf/vGIFkqpV3wJlhJTRkVDbwQXWjYukOXHtnnBeWnalfIxXXNgE3PnG6d9g+
etv6m6R9DgPEhbDHqF6Z+vO7Pg/vePPhs4p+WDt4SxGKq2r7SGMxXrSOQC1YVXUh
DjfFRz3svstSHZmEm0F2pFAU2Ch+U42Qwz4YO8onkLO8iQgZclJc2Pgqf5gHDelw
mUN/qbqYQ6qLtPwKbSqgbPsSQlkyae0mbX3powu+JIHAgq5y/yjqITWrCOJWq4dd
5paKOS6jsiGU3EfaZd9V2DgtL32Zq/hCQyxO+ZS3JKVNVqqwix9tCNpJ/WpOqXZv
Vl2d+cGGvtDa5PPkiZmtO1S8sxuoYv2/g0/jrwEo2uokM9UcVIA4CxjgOYMxatt1
jH1cEeuS4tUGQOcRaVysmi7Qu9HNbiJ7FhwfystL+ckZI0WJ+E8/z2LhOCQ3kB9x
nIWYjSj6FJ7eNcuNVcpJ5mY/sxdIGnOpj4Lik4e/+//Ck1WSvZXoILmFjZcyezLt
9FSKQkpVlCdvfs8NrNzMQM8Ki/NpcD+Yqivtu910TO1HJHrxrnE8E/jUYqBF9efZ
vOw7cE+yghn0LMft0vvY7JQ81rW94sn4obTEJsqtt4KZEo1C9tYlcvMIewy2BAnZ
gcnPazl1KyCchODhHy4g6vZwX8w76HGoxUNipNWe31E9NgFS/QIMWhqfxCiT2FHa
2jmj/CoUmtBdlxDoDmJjdzhc+BAO4aIxHyqrhHzORcKqbQfgfBHa6PKHnsH1uMY/
4j2JLQ43aNjVh1CrQHjwQj7OZdB8xSsTf+szBhLi+JFNztf+VVCOp2lTsVzSB3lp
a/J00GNDG8fLnLDdvV4ZHr6TaFg6q9GHfHR0tXOthNf4yne+rMLGyHPAmeDfsKui
q63I4KurgIi//sr66vxmZkTFTRy39YYkW8NimomfG4s24ne6aPZrP/g8vbSmdLjw
/6ZPxPDsLjnJupRfH7FRQcC6my7coIl2bzLoFqL9REMFU6Z1hWCxiXFKFYZO9h4i
QXtsS1CtwbE2sFCtccn6jH8Sm96janaI/OA5FJSS4trKQ91vw6j7h3v1nnCUpg5I
4+NrH9iJxf0gQJnILgN1PIQlr6d/4Ztw8HHoq7lxJJs7QrpTOEpzJOj73rAU2KPM
bD/PQM3adgfrEiSqnNAsdZaumO/EdS8ijsr+J7FILRMYLCQ3iDQVdMczkLnGmroK
WEJxyuB59UkKkVhJerPne03yx5t4X5lQt+TD5r2ElrL79w3gnVf49WAFo5RptPxY
q/uV4Hz6QVXY82ZIJMzr+bKu4KN3X3B6k2l36MVCFVi90+1KjXyqUm8YsB6WQ8wV
cRuVCjuc7QnOzLHt7xq1pDMVfRbK/Ck18JpwV95mVKMRCUA3rJJXwkgu1y2DbKkC
IAoCphVFeROlKSI6DPfIXFOcrk1O8zULibqlPBRc8+mQoMQEYsAjO8nUIlMWFrlR
nCpvHeMvBS6uvO+WNaK/rsG/UXPvuwJ19zMp15ex5FrU58sjTzFqPoI3r1wREjHg
wQTwnG6EVYREuBoahwbvtqYNuZLGHEMSc3nSrophb8m6Ax5hYmd2vG3yuji0A5Wf
d4Jfc3zHVDhaNT7b+S21EFO1PgFHxqaobqCLajvPWvrubaMVl43ntxzQ1rjM6yIi
Wed5DmCaTgDAFN/uumlH9TrO0X46azKG1+H4eQe/DnOtbVTd0FXosRMvEm72C6m8
E0BBe/3CALdXOM7BARilj9D9ogN6dMZH3sBS4QXmt+2uKzXQJfmsED9bNPoorhKk
bbMWFZnfZcSZMonH85ZLPeygmERdW8wDKULUHXuzyinQVAAVQ/rv31s9So+QXhzp
WQ3pENgLw4WSRAhF7tlY4PZlDKBvb9sLj/Kz31c6AdtX1Esb1lNubDtB06nXqM9k
DEzgypIDwESvq/7sFIJ5MBw2zDMeAbbZT7+2wZp3bRiz/DLpPhEtezGSOJQva7g6
n5HtdM+UwOJ0ZGMowjB+Z+DWyzEbQBBHWyT5M4vDzKAWIWlILxobqsdm7Hz1Z4XB
TavTmX2i6ho+6y+JMhmWVmgrHbgYtfUjHy0ju3V5tW7lqrfmEFbgVJvmiTEkcmt+
S+P0I81QTknd29QWY1MKiTIT/P/BWrWCc44cF9zHfJI9p/PVEuJIOsCQSRmHmFOX
CqkrdLm2WXJdjzRCCBufaLq5xFQN/ufHApo0sZK9mPOpaBVfWXnAr8DzF1SjioJg
zEHT7+V0y9WZum9UW0wPtjSETFfJdmgyyJ9oeKGiUd1HDEm5Ur7c1gu8X8eAOBuI
U1eDUW0vKWW2+yBZKywfuM+uxfQJBRPGZzIHMDFLfu6rFfBmwRSS7yfdm+JrpI8j
BluwGAdWiTatjkHjtsoJSaNaBnCqLZIn3UHUkuaS9Bui7ARMYpJa1aKuzFKd9nbk
sEBjqFDSProHi2ExCUe5wF+od9If5griILzRCS3bhFdoSSfunr87TkaDdTk+tz+K
cmIkEmo5GBLpM3UbPRmwdcbmIwhY/zdOa8gm4HfNZLHjV+aV/DOE+PZpGLnbKKkQ
JtQ/G0tmEKhDKR9shptUdmDELFItN3mwpnTFw61dfIMe4a3uEQDONk+SJqNT97+E
6Tmzpo+JoZtUBojPONlaIVI+tDTHZ5RC3Wkc3O9g/47G7pcprfYwg9D6k5qLmejE
uAJhPQ9RrSEaMr3q3RELlJbgiwULQfnvO8FVPfl7y67a4fLPRUWuBNUmYaKYl0Yg
43xgR38m78foJWdpJLQ843bkm8/5mTqd1eofEQstd0LHC5BhluZWcTljEP6ubo4L
Kz47YiTJSQ9ARanjOcIkekDQGOoLhC2PExQ1Jk5fyLp5XLU2mvQLNilHSLOVhfcA
z+Trm4hjpmS4hihn2kgHWlgwfmU5nT/Vj8Y4Xr0FpCFkyUdh84I0yDEP/ukgjL47
wuFELB1xxbCnEk4U4tw609ERoJMAnKwhPxvrCmZHDp84akGfV5RcQJgDUKn+scYl
hHjP8eWHNStFjV+FnjGMojIBUTnQlgG5zhE0uPczTnYsdb98z3JpgY8E3CXpuxhu
xyEKiBFcuQgSSRGjItaQgES1lGNEY5/+3LUtMzg2stkVKo0Bgfok9Ov4z2IW1Kw2
TzA3ypWhk7dQrSOgpSadS/Evj0zPoLJX1Xj+Y5xDMoYNRHDl3ODh6xCYSGTB/9jH
jZiB7nk10V6aFZNMq3v/RfmmYDN7lq37R102ooJlNklxZzaO8gh7ZRdAOR7ZQAkJ
51ePfpqi1zXXgFpVMp2GcTeZvvDD6fEq4uXKToTIiy9j2yGcfnIM2a4ELYmqkZOh
luaTILm7f41AzkIyu4dOzFmt2ElwN10ENp2bWUpSKvnCAdtExnavnYduBdZ0nJYa
IEGrwUzKSiFgndjizCMbexYP5ElrjFhyG1VPT2vJjmLyUnWkGjL1i4GGKB+nBhIy
0JS3/SAYA2mCGdq8rXA04IgKw9/gc4/aKJOwGV+xcZCTib+oo7oFTtQs7Bb+zajq
SDd+JlBINoslegNqKwZEpxbH+SEJx2MGUZaEqL+6vbpq9MS2YkocCXo0lSJyGH5L
NQz7lM8pczEN5AtXIWJQfnznyKokFYSIaBp2UiZUBs1xtEGrwj8rQanWIQaeM47r
3AvdARR0ay6LVrIhlKsW7wVkhDAYyigez6DvATAr70+KkGX/yYT8IKZiNeT1aoKw
RzHK4DxdLXM/eNxm+MBUeqHcFsZveSUys3bqSP4gPL1TDfmoMss2iHcdxLGmNQzg
kg0NGPgA7TaRTvhymqZ4DYLBnya37ce9EDkH6nIhtqN0eooTuvAx9Yq86ZMLqYUb
iqSDp62yuBJt4SF9AYs6zvcAHEV0XOjAnbTCjiRR133p2yRTsEBiFtwYGi3d06sE
CfkGQumRriPwFoORZICFxWBfWYbRa/VMh05zF7YKqNKnVpE33Vg/PzNBSxRlbBIC
UiOzE0C+RzKqom2mlcD0YRgOtfr78iiCqkNusdWQVM1sODU0RHx24p07dlQNaDD8
wSr25oIWsfc73TgaP+6i3gxqsfr8Uwnv2TTYzkEZKuFxfZw9J15V+576orcgmm3U
PeZzgE77WeZ83PVwCbTR0ddaU6FpECaINpbZNPMXTAh8FXTHHpQBKan5duI7ALIO
TiiQ0XDAeYtxmenPhzYgUkfO1XIbDzKxQ3J/yus/1DhtSGndy+mVCduk47Pl1UbW
zLcSKc2YXj3gUb+uya2y9eju3hM02Uwu1REGiuZTNrC7zG/sknhhZ054xWmnNTqK
JFrD9Z1JfxYZ9aZoqVJ39Updvf+DBwbI0pmoqC5xbdVOsj6xAEgwxxibqx4h2m3k
8uXOZ7C+QPFuDDjPjWu23kvy3xFQH30umAPmEoVUf75HjWR7eHsgLhgICwXl5A7q
E+0N7nKV4GLiMEZ7rk9GaSpoCdDrPv8D1oPA2ZkTY9Z5TN/cLoQWSfe7IjAVQbzS
qgZtO3CcYnu7wzPQcRSCW0UWeUTzSejKoP1uav1QjUyfgItmxP+A6btiN4pY3NoY
0WOpMRJsCvxniGDSimclqI60oYZL5wTKEpTNPGL8olAc/soqxyJ7mmHvNwQt1oxE
QPLuzT2yvB+COFzl1kjpLhlxJzyffTC5OcelcH0TkNpJz3q53CL1uafGSVUMA9QW
Pr7+eXXVdoAOvbbff5+qXiYz1og5dLqJikTDA0xLWF70GVTeCajQRe6Kb+Pxkgoq
vUig89DcOCQ9cHXOvmB2Lc6pulIN1NLoI5nYKYVhhD5bVK9nkvJcJ68DurHf0DHu
WDqSZtKtPRCOo3mU2mhDCEf/gPMg8toZzo493/ri2GfnLwdxDUSoGruxc9pH9wgp
PDBvAOdEbfbrPl7V/7TjY0eUjND51Ptrqq9OiD8s17oZLNAjm7rsrKIxXT8+DzuA
gp+clCjvQ3YqykBM+Wx88IE+Zods/tQsJJgeakf12ErPG4wDExSn+4EjTNYGFwGk
ThjARUhDWdup5BpCI1V3zZqKGSGt3VjXSteGXviZvdOJEkmYFvCIJgET/YNGFQNs
5WPOplbfQeyyMkpg6+a2oZ2xSLSvExb3J1Wb55LTmlZLfMICb4LzRXEG4urax4IV
lZM9IYnMmM7DOdXhp9mfujYfRGHG3Io1+KaehPDIT475EC35K5yNcd1wFjAMs7DO
E7l9q4SCwG9lOj+XqzDPm5UvnoS5ee7To9fZ86Dt/Bzb4UtVhN2VIYPMXmdb6zdE
7004cYBnfcWntOHWjnhYblXNWZAWyQI9T/DyGUN791n0eZW6zlaHJgUu00n9+HdM
kiJ1jET1Xp1IOFDB/q4XQeWUftbsFm8+3i94yO9HcurBQUxFV1Hj7AFc3jj+U7Yq
+P2GTJezKT2Ptzpr4KCl54kiOoOVcwlAY5wkRglleVHyzZrgVLpy6XaSj4aSTCRh
4felYqRZI5mgwPwKkTvplGIQb1vxGZzOmCHkTXQfYyVGzLr1Lf72W0m813s+E6tz
rZwFxgethVwsM4GVo5+1FA8sNlSibMxgQ0K48zIjrW5DnwiuNe9XMOA//nCRuizm
N+1+fPaX1Oo/Jk9OywU6VrHbPx+SMJXPZ7QCjSRq0HFaV4MWN8s10GtKNKRntdrH
f+MA7BAr+OfO/RNYHRsfkhQtAfdTJMTWMk+SwKbz9655wCC+MRLYKb0YMvkHySOk
TxyDwbFrnmWARzZ+gTfAi70gffxXTsPYuPCiNU+OQQXwwPjHcApLJPyEGnptz8gW
MHORqKeEMZZ7KPoYN0ILjJDBr34uD6aSTQ7jN6mB9czRfFHSM4dMEpR0TeyXvx/L
+NO94c1hgPWkUVXLujfU/M2jtOkN5H4rBFJV8+jSmlA0xW6nCgkhemFObyGpZk+U
QpY2iRTpDnj/jO8AcTw0oL17HARkdiLO1vUZLmOd0szUxHemzb0L9F+XEJiQyQhH
rUAC578Dcw7X+0RVPCCZ3NkXaWEq6b3mfW1bK8h917yjbn3UPA4lwVIPzBiWOWot
0X9N8u8ZnuvSIJXNSrlKRdxii4O2o5i5iqzqV4tTMxSMWPts+KQiupvzVhBKndpw
4ii6ySWqm3dk9ycQC0lzPSXt3Z19N44LpuNYjx3nPUmtAadHHQXcMKz68OZ7urgx
QpKCmTf5CSbwdb4OVRvRR3FntBVDq8ymCfQ2YAJAGfzgP27ubIIxLjyXUtRoO9Ca
9S8PQog/xOeguyphNrO7Tz28efjGZqI5tA0VuwuuD3KLowOrqFsVNOi8ie8DXuY/
xyEaa64eKDGlY3pd4075RS8bJdxN7Is7s6lNzgkcvAieLQVt0u5uMfoxI5fbHgiT
Vezls4Drvb0KXcuof32lmgK6cSDMez5KJLP3kyJFIcEJpESF0Tf5Oc9fM58PQ1MX
4HR+tIftMzHHsLzijYTRZ0hGYF63wsjO48yvPtAHzO+DuR/lbdRYEAlkrRh78J8n
xJzjAkQZ/gupid234BRpaTuNG0w2FAIfaextyOUnGAd4P8IUiulYb0+WB1n6Jte4
dUPN6NfppZMEBE5JFOssMPpDTXWAn1d1yY2J1xrylTvP1QcVhJMISMykwM2ezYvE
L31HLwessLdC4KewLrTQzgUlfdYf5ueB7BUYTUtRiwG5Gm95m+FWy7uQ45Mpltqi
oaQn+TfXoU5iMDEkJkjMwYUZ1QDZL/SDjELw/+eJkpql018oTX5VlgPIWLG6lM4i
2rGf4KqQuuGDOclzAVTHSzKB8vvsE4Bsr9n9MIZ3iHoZXJWHzY4SZ5eJzFhvIW+W
SU660ZDbjAxm2cBedQTW5zA/jAud6Y30aiQRnLup6siOWXAVyRTJqRPeLZpBPcUK
HCEbHP8KcZ+v9fKpNCkHeyBhFZEi22ajX4y5STH2v+2KBjyrv0WAtOT4zoNKYCiN
ro4mOKHTcrUCTl/MUWxl7SK9tmsCCbiDl0+S1qoyWY5euDOq0U3yu66QOUotTKH1
Qd4WLpJjaeq7UV2Z/i0ML1/uDcgmvj9vmHwJdSokpne1kPHIL89wn/myMdRj2g/9
6EXLcsHxFAQJP+S4Aka/Mqfpg/c/WI2dotoV052T7SgIdGPozEj+lC1DuIXm0hhh
i52fcbTe5qaGRp2wLEOa+6MgbEezz69ItIqxRLJPwXAwnugprwDEXVlH+HUvxeRt
qkfQ6gdkfBowdFJappbyMIdOApU38o7pv3XdUEkyMg+CZNzQeqTSHdDHMWoMrmX9
3hXzCGv3iQXoOX9jf53nm8Pzm0tvDVa8T8i5nKBdYPi6zfp9/ejc+5g8CMYUiQJh
Esd2W87iS+imX6K+TZqRJaV2PMO+ZEXrv6PWnioyiu0uJ+fj6RRIr/PUw2+2XbvO
82hUdRvx+inXXdV5fo+/UHc5DVRDEymW761qebckYZ4VjPOGpIc4Fp7jXC/NACB+
QuE60AGRuNIenrlZg90q1e2kn7QUec5azY1TJeS2a3lSD23ywH2sO5yuMO9XNYS8
NMkx0dM/TpczeFFwR4neIa81Cq5jc+T42mLEy9ss74ZXpVXj7lNhN0l7cOLykcGr
0z80v46313bf8Xu2yksmVJqxK4y9CSBI7plxrFHfI0VT6xM5GCjO6Vj1T1R2yNQd
DcrRhySPKqY5Ulq0iDUsfgeRu+B5H6fGcD/MTsRqyUJcV84rO2B3zZIqV3J3Ruqp
lUhm9VbDES1D+pZbV4Xg9pAoOumPcMeMp9bvcKUJQ+q0iUvmF89xBhkOMoIO5Cx1
Tu2nH1QSnor6ETUHOTr1jPgp0Jn9NHIxqOfdUnEs70T2xuZi7bsZ/uFi/m9M77tW
IEDI7sIOR3Ldq4JcO7VVpyYl2hr5fpWzb8l9hW/+OC8fFtwVOhv6n7lvEh+ftWJ/
jzVk0nP8k7YZ27eJz8DvgB9oaa5dlFjkxxoSAN3ttAP3pGkAEgWaQkWwQf2tKCU3
Zh5rJrB8K0P0SXNuw3swpbd1WegoWsINTxNR/xNf5Ix3LJb3ubRnmBjE+y7Suyc9
ca9b9U3Yj7mBhOXQYLPYDFFMW4xcRG6ooZado0YPQswbn5grE5KtzujK4dAcKCJK
TUXGu3HXh0rBtzPE7sJf527OA2NMVfKocfPxdJIccIZtHLVASLE067vqblzbjt3n
+/hFV/OX3HtQ30zUDkUojfYR7l3qjQMbXj+sMN44+T1xfjVp6U+m/zGQQfsVI1om
Wg0X+xJ0QN5VjMyhdJNidqk7qmPXeq0/s1fgQMuB59dqItm6uY8/Mx/z94wVPg4i
Y6nmhD772Z/Ys6oBtHReIuAwjpbd07EpIXQYJxK0wFlRLLTNB53z4vd+G633XMrG
MHZOzrPL+mby+3AAExcS1m8KBYLTntyjMQqNLyeSlANFdImFRLEFwPksjusndR2c
KaXbVd0YqSPDRQ7nQbKfsABh2m+G/63p7M5hKE+6+U8jJoRBoA+QJLtfffMw3Zba
J2mPnSHf5HJL3uJcPFJJc6ReHURcQ1Car03JL/AxhyH4RP+I5OHfPxCy1y/u/ADs
SLhntzXT1D0CnIASmcP/7bb7PoVyW9VGEI/iF4nLR0PKM2KkkHhF3jpcWEDAiR0W
gNGDv7hJmwj9FCNhM5TSmsYzHVyB/OztTQzXcp8y4JdfFzWHxU3likYJqXWMH/Az
gBuZkO3Bv07EozE5loErQKh+tB2GpYeiBrFvwb+JudAJ9fYZcAe8c6ASCHr6E/GL
ja8LTdZigxyWtcrrS/huDKvbNO3K6v0XPIa3L7B8npNXXslbi1LIQanNH1fA3Lfj
5cyyQKDE0aOwWiIDzThMDH+61fsaSO7vAMBa1JP+vGxS77ywU51xxbph8l9RhzLE
iA6NzTRBsUnEfc93t53995DUKk4INK8rDg8Hbde7uLeU8KPOeoq613rUMRPNOYq5
m9uRKwiTvTl/6Lak8DjpiXpHuwU7sAQtEOoiq0elVEPvpJJ47pv+UOdtCzfeIJkH
ipuCOJMQA63vljKMmb/JEZBU4WlnvI3bsSD7htxhZHq4ohC6EMholmP32kKpuMIn
9m/P+LPyXZzbR+fpIaA/Vcob1nM+Qd/0+9bFMc/pWPBhkjIFzwlGbjLk5HJ16Laa
dNDzPrhUdzmicLdORvvRK0l3PROFBgOYfSfGHCEu/JxKjaGMtMJaRNJQsSf+MFM/
dXc4J9Z//SlA9exPos45PqmMM0djy/J8olVD+6AzoInGBtoXh5pB4jIzs2+PfhqI
Owsm0XLa3yRXkLXFq1I20C1rxKWdIMDC5eay/WyOJAn1mmZ2BMZdx8bC11eIqYnE
JV8e9AoFNCtlFAXCN3l6OMI+QOuNmU4IvonzUdLiSE5ly7dQXGCzjnL46OhVzPYF
OzA1AXd1Qx4FcDNgZCFlGBOpHf+RglPqLkCb76ClZwVvXLoZpVAg6/7hhQWZQGyI
UgjfLd0LQhy6xxZfTd7EIzrUDeLM/RjXSB82fuSRPF6avz9eJEuFKr1PCLoV6/QD
56jUNbXq0o7HXG7xkmaX80rblvpyV0vtikQ0YCJP2KDMGVkgbeIMwjNAmZi7Yboj
75ZObjj+cXP3Oeq0DaX5nIdklRChj/cMnACwxHf5Cyk02FHpIJS9gFxaKikG1A5I
sL8q/bPRnL6f2oaqB7mZZo2qsuYvFFGtDXafBPvTwAH3tXbQZXImKg2TO2jpD3PO
lRjsPT+rO98f88+8KXoe10J26/+xVgIvvfeko2e34rr+h/8lCZJtStpRpr/J1Ay0
Boc+NLJjDfgT4AItp8IhMu36605ZpqE4aBEbjxN9XN2zix9+4il4V6dj3D7odqVO
F6zmdhGIU8lt7rm8v4o271S9hCv5jaacU6jeM1tsOiCtF+71Z1avaCQaYuKNAa6B
55SuIKGOYrWm7NsxOgwikvO4qsGKSePMOxw17WpnARW5tV7hSOGzFjsrzPicNj3d
oipKhPksqGpQSbYab76CpNxcVCEgZTnU2z3Rjkd054jDoj93hGHtd8himaD+UVYs
qhyqtxKorbCBLV7e/LLcGqDxD0tZ2gu/1msvxzz0TumnsDXKWq4ZIIwNlnEi8fX7
hvtmn1D9wJmMPaE767//k+VFwpXT3IDGnRMrLsA4wJsvfRQvb/zfxdTGxF49Mjgg
ta+AMHX7NGe0sJh1pfWBxVUV16ezUXQmrp9Op4mSEsgXrQwmU/M3K6r8eVskqNbX
qCaN5oxz98pkH4iC8Db0dYMrY/RPV9ypr9mZK5gyCqs3eTTQJbmvLnKdX3HrGhit
CNf0c0aiVPSJCnJhiUAD65KkMGVi0YNL9VHYVbiw6D2KikGzrjSFSle9SOeO78Jd
+Zw0/K4XpW8u5OFiSQBCrOsGUwn4O92BOoWkZZKdNv80nVac7LEKX58kz8BW7BAX
pXBqfnaM2IZ0bT3MD8070gDP09Us/jRDHXQtLejys6ErWQXjor+fyU+6alMamhxc
a15Aeasv2e8KIYLsIX/IBrPbTOkTpfk5q+eWkvX+8uHwlI24ONEmixTjC6mreVov
76ZEyQ4l2WFt4Hxf5W7dEe/PP1xeUkJlNKLrhAy598Jk6QVh4mq4d3f8gJVqIWR7
tuKdYP3VS7SbWj7OEuq7oEzXfOuX4+rocm3DMSMcBWD48A8xGbA1aArWVi8ZDqaZ
B/pDYAB0WTznY83SeKwR3PVMHEpWgDsEx/4SrRSr7LuCfsZIeNAmbXSX7JOG63cD
z9LIzTDhw23FndWdEvzIevAtXJsv3Y9CP3H0s6dnq49PC+tzq/KejcwF/kpHU5SJ
Nnq+P7oRpyiG9sC4Ecsrm/x3/90gVW+LMH5kX+8abSLebIQnRryK8EwsirzrGcCY
oBCPrpkHoiz4lj4hcsTtYxSblcPLDZUNx3asxJWgg+JAj5bBjkClLuswJvDNUJh9
utBh3oef1T6z32m5BGxZfBO0sVjB/iSJGmsBnr+nkcVsY2tDRBcdoDWq9ifXu/SV
v+RZyHVpLTxSjgTMjF3d8Fg68WkdcfMfpAtwP3dE5vsWJAflUn7aT9i1KlOBH+9O
Isl6KiLLbToDMuWyUvqVCUCpDUyZbb1Q95fm/xuyEA4+zNCwX62R37QjEd/RHLKN
TZpU4bkTRpYBPn1iuNwL5dr5XWKlGyclfkJ+dgiRNcP5MyGgdouFWEcS9gw9qcuW
H2tjmxyoCV4Ad4DLyhe4av+UZMtNvxmPhRB9F3vXj9/qRCVtX34BcbGBLG5bpCU3
A9JzE+ubw9N7ghsPuc8OdeRcF3J7m58uf/5H2A75x5tpP3HY5ZMLqixG1euP5GV1
gq0P+xeXyx4rGUMBcZWp9eNUE0dly3e/rdW+oDMFkL6HwuIA5ABp7Ap8z0Y6bKa0
uyOox5G5va8/Sw3db9V0ujkMZDLFIAMcaJh6x4oiZdWtEeVOzk7IrByGa+nqRSJq
MdMoKN7uLf9Vg00brrVo6g8BhCYhFA3vdmZYSXh/xBBozSSyeBYG7jAY5qVRh2kR
+XZfJvHWKbq4L+hJLb0BLm9PYT6ldIr4Tvb0/gF3DAxNBrRQi40ka4UjvVmGb0vA
JF3Ctl3SxF3BHmjaENidreHLUmrlJo+AKu+upx6u0JO2nKvqTtsELAnl6OYYZ0Ah
6mMJjTyPGJzm1WIvF/Nkurk+Am3yQY3YbzumTuAlQoxnleAre4B2WpbhjfJBtcaD
zcGQWAoFehhLAmqDViuIybfOp489Xex6kx43GQJ29ZI02lIO5sHyVvjE95RWJ8k2
B8Y8LKcJjHl7bdaSKdxu/XhjWbv4/gpUfAriiVxAxslc3jcaRvpNe7IsOERSraCy
5LDcSNmMTIPlLxjHRY1WIrvVLwZwF5ih+BVuhovP5RaefE59ADReWhrYqBcGVm7A
+YjHUxVvkAzMon3/4aOSlkTDVmEz9NqqaicnbgojQGFWSRd1Y0NfgTf2wf4bQJYp
BvGcQgGD+VZnfwT2rjW2sa8hBq0AFe18AqqfEYWuT8SqRW1KZadE513rDaE7E92N
tc0tQ2ii9dItfp7dizsU+oTQQdDf4aZg+tJ56p18cubVe7fW+OvHZRkdFeQNb9od
g7biJK6mNi7j6DJrOYcCdXFkldB2BsBoda30lDYNCJLQdFOkntei2U82CsPmdxZT
w90oHcguxGWwkdwXGYbBSA+WTyMnXw3RgqVE/Gcg8eGCB676RpVxpjCw6qsT/Ukx
h8ZepmN0vc1RRndJ4pJA4GN6aSPdwrIklM3Ucu7d3e0DhbybKOMnl2Y4tTA2U6oy
5K2zJa3ukgP8eEu6g7JcU9pn3VDNOf4l7CFL+yuDoeXDG9XmKV5pxSKTbvtwJ92W
K9G3UBsuEI4bpVel8iepzu2gsd4ZG/uPg3IA/sCsIP+wxel7a/p8PT7i6fEjMydc
5iNSKs+rbkRopZ2tlIgRi0un79WP21chBrJpRGCE8e5x8vmX91hG7EVGNps37Ikd
FIu2j8shwKHAWJgdJX2E1Flk/76sA7Ms9VwaA1GzPXYXyTFTX7YNmBjawqGMZ0i3
UIqpQCI3GIhxyrG31MP15J5toBXHKsf+Xct8qVBgsTuWnxN/adDKSKm11y/R+wk4
zs4fbl+ogFZ5puTUg6c5FDVsFb3Gua6jXUNO7TW6wCYNKpdsAPAI5dQanwFquo13
Wm+l8Y6F//Ude0h+gcylVoNiJYXxdqNvXDjPgF4tjyaKtGWtlIBNomkvBqy7cMS+
YlvEug8bzxXHZHQ8OW3xfsbUqlrB5WPiR6lozABaCBZV3vs9YNtEXGuX4sN2jArO
4+pRKusSp1MSgbivHt4DENenD49kvJLmkFxr7xGXEkrGPLdPhGmjRfIkG57Mu8Oy
rluqwsKRCdtoyh2uoSaKjMQEvT6Ci4eaEB27ieHHRrOydRgjQEN3herfJUmL0COx
IAeESpi9j4sdF45t/GuM8I2MHYAM7jJBcxxPl9LMKi7fMZPcralBEBESNC8hrz2P
XvzTJhocB9a6g8TY9gm4IvIqYpzAUu6RTsN1MmWob3L43qddkg3+VZBfTolEHCBo
sTn+1tYq0GInckrAs1V4zUnEqR1DOgGS4K0ztShGiNL3czusegyTN7jG3IVMjj32
dKmc0owQpZCWXCqSajKGvyXvBcsS3HLuCCmCU0aHMRJSysLzSYgjdGzKMqATN1+p
EdjpBFocgDOnlSC10x/cBn+bIBrVE7cKkWB6UGRhOybB/1zIFcjrC4Df95tIcpHX
zYvRBWnOMDeu+DL9lcA358/yWnFIiRX6OvlsPuTH2aq1nwYV2BdctCaW3tQo5aQh
p1E6ww5x14u9Tfi+8G09q2O6AHwuCMzVsay12Epu/EFusW/DCe5OF32boM8EoPKR
KjWrDMwASygLlTagjUVMC4oMc3A6QBQA6EHxUP/acwqyufpHRuHm2/JbvGZv+dxM
SkQqqf+m2kmV7DVQvQPk7T4H/miBZhPIeNIEkNa6fRoZnzeT3NflWKjQKkTgPj1q
5welWMtO9pV3fq7R6EipUf3HI8p5Dd9A3ORjyq40ETi7uzAGIfwX67plpvGAzCOI
gRJ8uP3g9p4Y5xYPydihlXk4q7wLXtWrzuhGLdEogox5yll9YIHV1dEpQOSP5rtF
F0pYU5as0eNrWyE2v+jJnEtbGI+m2Vf+JT7S0W0maAM1I2q5OZyIntf+m+J1FqWG
2h1mp+pWHPgRJdpkgzCcYtNGiMjGZtENEEsd2ODgzXTl+dHuikpKGSiYd9hPLk3k
qC6zxfAfHXWWBJGb1GlkKyOha3zHkwI0eoUxIEwww2Gjf0+lDdmkfKj1P3HPvdsV
4x+M9fBWSSg/ANU5ucPM1MJJUnlUEPkQcP08oJm7zKZTw3IyLGpKKrC5Zy/56+Na
gdxf37G3C3MWfjFbRgABzQMxLPSrvbzBcJltc/8OQEBsuGFdzRfIoKOT/dd26ziE
wTrepnbZoirC0Sad7BO6mp5YS0vZAPWQPgdqbxk/EKIVzsdmB2cXExQGt995u2LJ
gVYAmjqto42H60U0PBPG1DP+csSyTItfHnoe6h53ZZfAyZcMWmrhHSXgwTMWD9Lo
xY8o3MVN6RNIgcsR3Vmjp0FkLvNfWgxuJYpMQ/tId5b6ANPw7X5o90VQIq0oCUUm
i89eu5gVlS0ZvMfGf7/AoBAxdpgBnxebiUcGUBVpwdTKwBX5fQl1PaNIx4Ze7PvI
QOL4LJ3MEodDIlQgQpbf27RHV5Pw1Kg3b3kjJCFjOiwcWpHvicJOlCaQaOsZ+GyG
+wKg8QyfR9e8a6Lasi+uGOw+3IrZd3v2wIYbP22Sczw2/39IjpaLVngZtPOnaDMm
Fsg9y6D2RyDGIafBBCbaN+wsGzJg9lPyhCc60kZ/PUf3qtYpcVB+VEwAgeIGC//f
jqoat/8wMvvXynxCCvOx40Qm2J9wFUfDjInLBZ1H+6XA9LxkW95y6x0H/YsJKZ6J
9LPT5gvZOpgKtw/iGhhEajjdvKMH9mYC4ht3SQ2UtLqKg7R1cjiweVhEb81esbh8
q94fIAWht3wTCwcmiADxMmmiy6toBULYPg3eQREUVXFo7et3H1OJMo2TpEZfVvIR
g1y/J+P3GSXP9PDMBPrkGWgz5EyVdKMIX1uP3ENANB2gXe0g3yZOhtsi1xf4PizF
0dXErkSgS0B4XouB1FxXjmqT7CsK9uB1n2BNbhdoH+4EfUxZMYRydfVDUCW0H92Z
tgl0TuT01dox5vask1B7DiXQi/LLdSzwPd4hdsG+/9FaeKBnoGcmnbs/FnqnP/m4
ZJEYWebAnOB1ymansDzqPApQFryuLBoyab3kkw/IHvi2jDKOfHzRBqfd+6cNgwBU
6w55N+DjXZvKw+IEcAOlGM28/rS/9FhBDFCiElwbnH/rfaa20okSTl1PAkzh1qH+
jkO8pTyHNcAuxIwWjIpa1qw4A4HoFtWfzKLjsjpZJFhNsSzTrXAqoczp9XjpIwbR
dNneUtj2Wnh/0Naa+QxiYgc5eoNFCVDnGC/OkO1vaHt6d7Cjw0WS/l9GZ/S7cTUB
cyp5xUIq6ndF5737YhgtEDC/ux6HS5p/yfMOCh3yYRaKOQOIJuetcYIETKQh9g9h
rMpdvxllyHkCI9tTDy6cgahUDIzoY50HO/UHeKQjOJkD9v5ZbmJDwa95bej/0Jcv
7kXQzWK+fCVjEduedku9M6RAX63zibnYEpDXV0ETLADcc5eEL2wI+ZrjnMG50DRE
1dxkb3LybsJP3+3JBwH3yKPQXxLRRVaKKpSXqQHFA0TSr8sYXgKltxl+CrrMXLsC
fW9qbecjnE4PBN3DH0pPI0f8/7iJJ2GIlCHH3gL9FQa7GJcg1bwzsIUKyCZ2Lz2S
MotWsAQcQu48fv09FQcAjSfcy0VA0QgqOJbLXEyyKE7hsBnrs4y9K7703tec7k6u
8WWSp2oJzjKdxUo1oFM7L8oywHskqcu7qNAUOkyM/+w7cQAWCHfltZl+b5AU930W
+wrnQvKJxvk9Mm0WHJUAvmJEf0YuDGa/+myGpGLwIQactTDZk6IZ3DdD9D0VUVf0
4PQJZbnFztDlihC7iz42SZBysaM1CSSyZSkeEbzobR2bUlwRQQOGJRoeKdfOGWZr
Z+fG5xqDNvy7L4TEIH9RL2iyLnMk5G6/zqal7+BuFtv3PrpHCao41jh8WDaZH6AJ
6Q+Z8BatlGuRuRKvghgIQf0Jc7Uw9DpVHX8ykFnk8Om5h9fPU1KLQk4YFjWYXcCA
nz/QcJcFCLMnvhib+w7CWShMG3xyMjvhcsSn/atiOMow/oNLIB50a4O1tLFyShxu
PD/biStllCjJZsQVVB5RNC4jCel2Mb//shJkcKtnhg3JI5TpdMLMk6GyodCn8vnV
jt6y9nbjjRB3aPnbDARhi32qUwDtjKkqKFYnswM9njYrcCp6D0gvi++T4PSX948R
mOePkhnx/n12Mw9GVZw0lKkCtTE04RFqX9Odf2BXSJLhZZ8517+K+K3ICAOHCpVT
Ry431pQcElH0MEmfiVITdJcXPLHgNlmy1De+nuVVYRaoyVroicBv2nNszoMXHnw7
WBxZpxsHQ2AuyfN/IfWlHc+IIBFXArd3cVePl+I2+6OERlQ06XIqOrk1Od7JvpX0
o5xv2o2AZf3VFuSZktVAiS/lnWW0g5BEb6HQE/YRIiWefKyk7Iccm5/5+DmUWL37
s0L6PIrr+9gJpXG64WEO+MzKMyhxLzhIay/SyfKhelIlyFLUB+Sr5hMjjmBHHhXp
+hjjfgvUeGbj0hRcxFH6p10GAqX3R2bWLc2MAhmY+B3AyrxtYu525zwjxPlgN5gZ
XhK8AlCuaMdM+kXTwXcItx//YopG5lOZJFE2qZ+PG1J53546EQlEqt/1A6AHtnSy
5F0GHQHifVUI3pwgJLIh4LKCuCvF+G2WK4R+8+OEjds9RVe8xgZiga5ut+O5Ixum
V4qoNXGeLPkA7uFVJJSmwAZgg+nIHaMXE27omZ2tFEsoxlEXFXDmnp3G3Pd/n541
ExYB20qLm+tnjern6dxJDE8W0/3xqwak7c77mFjPqJwcqeCfW+hv4wPFmRqKHP/5
l6Y6gs3FbG5rWxij1aY3YC+Py7r8zAKjURAyrnrDFlMOgZ4yrSTXXs2pVr6fDC/Y
XFAMUFkTQ544f1UQaO1Q2YHE9tTalnn1F6ne4cG5WlhDUC/lZobgPQaDGJe3TomO
6bA4c/Q8mCiHYMhsndTKN81/hF69nyCQo2Da7ntjnhIbunV8L8GeXOy62f6VLqhv
/DcGM1JE6mrNViX+OSD/fQ1cKNBnNh6C8p38iaARJ0OBh0o463WvYGzyjkmSThus
sLy74EgxD/tEnlpq3bmMHIND05IDNcNVQs40HfJCfDmY0GoUfsxzGipAtpM1wyjK
Hw7gPXm5dSzTnaPY43/0OjXjGGxOWydQa2o8A2ziXZy2GRWJml3JfCdCnQNL7n8F
ihFxZlayhV9tfUC23QJomMZ/KE6SkC8SH1PXWIHy0yfTQCOdd1Irv+Rcn3caffdH
MlPo0BBwztCXlURFwbSDUTffY0sD1xHktaKdMnv/797rAxEaDL9vftw88TpwM8L+
53d+CB/bW2lFEm8nJMmxjYHd8WndrJJecnVAWvfc6Et0obQgncslHkUv7n//7Bg9
ydR7nEj9Osm+vDIrFMitPLEt+OgZ0whH2pgsr5jzAfjo+0eYYZ3HB3Wf5SVQuGrw
jnktHQ75906dnkng4KrEgdMsAMNo0+yTl9PSEHSLXWLsSpDsvsu1uaiV8ZotTEdG
v8FKvSlMsSK5v/deu95TTi5LUZCo8EWph9zOuC5D3W8pzH0hrrlb45PFMfO1IzUW
BBenZ5ZhFESVbrCff83UsZxBHS+Q2KdHPbeKnCgUnPnU8j/jB43ffgqflGCjlH3X
v4ASeJJaGoRM8v+j/RzaUcRDZjfp2N5YIEue0DonN4qgk8xIC1j/5YEFmhBbo8JC
nVnhTZV64UiV1VQ8nTfwMEninHZswz0Sj0uBMSPXVpWzWYail+lTJMCf0sX4LtRt
/F/OvKY8uuYZ9Y72D6VdmTaXlp3RriF5o3uVCRbu9BrHwmmOiZa6Kfe2L5bqpB6t
dfoikTaFaWds/Cutzmm6JtWP5j/JK8nNMH8/fS6KjvTZemZb0Hld008z+om+Yyaq
jwwXlV202b5RXa47bIu8sdW9cvM3Gf8t5A0pt/9eel95XqJEUbB8a5NTJGDQl6+0
qCifzbAdMe9mp9uNt3vQfzFgcd1bfrhZx3rjng9wLVld/IuzeP9Popr1EIR7eOaS
/beU+A7+XQ+G0s4LSWxLBktsTrmYbV1IT48aExB7x5x/NAvaZ6EwhrdZ2DZa59eQ
Y4V7s3P/cKlxStcsHV5ETS0yjOXzyoKWdPz9g94gUkrwswf+85MKO8iHLA0nFaGS
IiJLm5jz/WkVJHh58CJzzmJEmdtADLpz2/GmoUsWN6haAsPyHomJ//pTSzYd3Q3t
NyLFJaOijOy0KOaC1rS6lpNUI60LKwdy9u2ejoDD3S0PvJAB7qipcuwWjOb11zGx
x2EHOHSiDZyFkfZGKi8M43SyalZn5zrYejIjJET7GocYRANvVAuMyGaSZaYHHIol
JS1RgdFT+IXG0THg+G6vFO4XTa8p8xAeWV+kAJj6PZknHaQE9V7qg7jgNz2XGqVV
JhO1bCv85SLJBGCYXnwIpU23z68KnPw6AyJ1ORRECyZ5HYVeXMNaf+UodkD7F++d
8/xQNE13fbCtAazB2o4H4cc2y84fyL354RsXwDOU3ldlKelNYXhoNeVbcaNHB3ch
vt+JzUH7XpUA+9UQEXiWTSArLVPgZwVDtK6KPql+MUWxv9Mt+jcFsJbsw9+gGvQ8
ddm7puEFJ/6VnQbR8+yK9RCnncLQ/2pFdBUvtK/lgwuSzBuIOMKZF8lJMOD2qu9/
kKLwqa+5rk+d8hYIE6nl9XQyShFJCtfPBjq4Y+KE5YotY8ITHLJEybgCr2/lTkrZ
ke4AwqA9/Oxy73euf33GIrNIoGQQUqwOzwhst2pULX4gepC51v6CXkT7cNbAIvPR
vQoyGYuVn3D9g21ipKSC5bGZWCpM/3DNagHy8RfHw96SigrRFOwhrrp46E6ic7Nn
qXUyxNPsGQwTDca8tFx/HLDT1G3ojYtpz+m/ywHiQLANxZ/qRSzIL4jDBOBmilW8
oneV0MQaR+q6qYmM9/H+7Gg8uEi8suNFefowW/o9hBVZXwNd7+xYkQ8TQn7YwnHJ
2iAxZ2jjXTT/wRaL1ShOiOtTq3SOGqZ5Lqfcy2/Q1/eznKxJDjFtgXeAvPh9ykUN
fxsuEb5etU+uncWdod3IXwe++2X0FsFPpZ4Mfo/Rh4OF0JZIQguYGsbqUqfXrfBU
DC+bnXcN3wZAxUoWitmei2OrMVuVdpC0o+kkINWSg2aXrxWL7Hxqf10LDRht/Fdw
eZHx/EpnhjAJrts483MN53V2lH2vHjtognghCFpI+dHX3mBV7a5B9UC51OKMdFwA
OJ3MOfN/iGRW7KuVU0OMb56w0weIgzM57huGJEE4X03tw4choCmN/VjoLjKPlzCg
kUR7mTBHJFGuCS+nwJs9PPA/xbyk1D43YAwUiXpvyu/hjT4Myj6ZIwyRa5xoUKRs
ldlfGxNybOkyDIqV3goYAa/V4njmcHar01lw9bT/atqhj4k3D9UNgGWiTThN3BaH
+u3IEwUr5vuEfyWxGZi1/ozpgpPzZCLcCbWjbm180Ng4H8lbF0Hp3t0i7MRBIla4
528S8QgqZQ2BHzu4qIhZt7oF8iSjmEyZobEJijqMi6CV+KPI7qZqLB3tBuJhfi0P
I3NwvWeF4tZuoLbv1gPzrKpDo9emND0YutEGk9AWOZUvuDtinDe27MsomZ+aOaR6
rGnifAOcJiMTzZBds0nVFl8QN1NbLU3xIqtPvw8G2Supq0wGlZ1ehPO7P6j/I2/3
BP/NmVJo3yuQiesNzYX5RbqBcW02rpjXkx+JlNK2bicdX5ubYmUtXq7kvSSERlwq
KZm6QDq81bDiSsRzhB1vEYd5elDlTw2DiBqm/x3J8zOgWplT5sgM9zH1pIilxAgY
obn7fKSJZhVeyPmm06r0C5rU78XyRuYXe1uKGJxf2X+wl7JGmitmhDzkI4nrm+tR
8V8FpBycGBhSAM/YyvrqjBdqGlmv9Gi556rCmjk2q0Z4M3dfi8zW5S4OW2MWoPqI
CeZMxy4nqcTD6/EdKB/jpb7p4Ra/Aibp9l0Mij/USSnUpuKtJGuGtsiX6y2Z3Teg
JAWK2UnCIqmE2SQyX7SumjRq4pkWhtfYKKS7syrN6kLLLkUSDWFI55Qrr6ZFAZ0W
7ozWmMFdmIXDNwy4PqwspDUyY3+ViuO7KDyIh8M25gYrLP61+OZ33iA7ITLooA6+
hs9aKfgCoI3Fs0XhxYCrABuku3PWlvps00QDgW4eFfXwKD1M4IU8rFlnmKcTJDIo
ETuypoi1e2xsuf5DYSW0UnIh+HnHnzg6iY0ti5hy/hny6Kt+5CErsD11WPI190UW
dihPCcx3pL+PNgjg9+l70BJrhBK55GrY862/cAD0s7ApdoF7SnqT8K23i+4ID0jQ
PmhEiGssMb1rVEL8zjM80r3BkEKBHymmIupXnmQtdEanLB7DUuFbFmDKLjsPoxPa
771nnqu1x0mgsoRUy9CE2hb9WFm2B33scpvhNYG9GWLZys15DXpxOGb9l2GFclWH
CP0U4FXRO7R2eq6kDTD3t+WDe7P1+n4NktcGSqoRfuZfNdH/rjeMtvL3BE1D3ZTj
Wz6ibteEAkMqq5A312WjtexYse7sWiy1a9OvbhGD0kwE6ylmFp5rl900+Kp4i5CA
H1UYqiKkp/nNFJmKHpKeE0fFZ90YQC5DC/hgl7PgXMJFPlYDKCPeQltDud92SnMm
XqAQJzohJxKuzxxZ5mUMORmF6t5zt8/H8UDpWlLP+CE+FH+eLONaIci+5HW3dcWN
hdY0+N+hNyKZKUks74hybsVRVMhSzAMLEOrsD2Zelmi5fJSKIS4SDYm0Vy4G7MCz
I/dWcGW5pZbaZdw34eXu2xh7Xsy1Gkm149oiNQVHI3TLHRS+E09p34Da7Ur3FbCM
d/2GkHAZgdpwdq9k5IiOunJsclcDDQvm+HQTjD9bgSYOEc6iP6B1wHTFsOZuIpax
zo7+PBV7Fl3ScCW7Jh8fxs8OQ/lE5RI5s/WDU9Cwam3bl2Rq21sXpIe8iDNJ5NoJ
lJt7wZDK/mqBBwXk5DiveI1BLwS7tGzc6F2je3ohD1fpx3+2xJHnAMReBOOaCkLc
UuOSeifeTjI4yPvXT885nckNBU1tC0eMJPqWXG5+yeNCkMV5slrPYTcxJsObQlxJ
XjeoMpOW+5/3FFmKEeru0kiz3BELq6NFCh7szKb738KTu7RIaN8a5stJVB+Doh7A
VCxm/91M0cQhz8RjGXdT4+7aAULTprIFZP5QuFfg7DM+JtDlXanQc7wbjNsSkC4j
GRrhnnYfRd2YdOl1E85DgvYA8IiLLNlAGIVsOHDqfFDgznTHq208X6A5SILoZ7Vb
Gk+Z/nU2S3M/9e/tc9L5jDooMVhoc/XrTgN2jMVrEYCbLpO4c/bxo7daxICTDTBv
/wSkG7iR/AlXHhV99CMKR12T1lUWKmO3Jw3EltM0G/p4KPu21lrP7Ck0qHJGs3M1
MqYb9h74Ta5fCrtDZLXiKWYVKyGjbCM59Npk+yWGcAIzDz8I/mfzTmLBb1UXlZlO
awRFoZeQJD2DPqwDsWuFzu6cwx6lB+DUHy6vseZ3SXroWg/zfISXGUIpBR35hJeh
x/QhEFbBhxDGn0ypQNzXoz7YI8VOowUhF7TJfJZVzrmgLpVoWUqMr8EoG0iINbOY
8VMGYe2aU2+q6p30Ty/r77LXcBld+Ez23Ln3NWTN3hUNm51IO2uLIAgsLHHdZWN2
3CrEiIuw/aFW1zMyxyLjjuQiqhJ7kediSH4Y+NqHRacVLbaobl94YUac+yV03LMm
bbiU3bDoBDe1754Ah9h1erx/NI9YUfWgJ1rWiC4PRuzOc2cFo8HxoJG/23U3ECkP
g/bAm8yPOGRUbOQAmaOba6qa+/PmYwsvHbXB8mPTnotZgYQwEhxqsCX4HBDkUHCV
Xzf5splXEPFl6xr3e9+DnIb5AEgFLp2vqJSH70HKKWkLgeaSE38EWbyGhiPLyZLL
1R0lBjrNexPG1XwCuWDuomRynoSiPQ72hNIRuLOoXPb4ZV9u+QTzStOXI+E3I+o4
KvgkdfCB70wZqmn7JQNreKN3LSOVzXArkVOwB1mnWCGvtyFZbKvzY//e+vtHQFvH
WHaj4UFq1o+zt1XiBWgwFtSR8ShRZinEnhhT2tFdBoPjIpjqevS/vJ/lqzPzarHe
KekR8PqBGfHFM1B4djAwnkMKDRcMEmql7uwGb2R0/8yboOBjieLK2EJYct8dR/si
micZm0lYKzUClg5ehxIgPBl8Dhf2u6DHyxyLKwp92AGrhIqsx88fIojcP4eQDJ7w
0n9IPJmRWbls23hORnxtRsgR/eJCVpK55oU7my3UiJF97BDbDm6ty7njbC68mK7f
f7aKxVAC6TF5Tpog9warg0GloEt1/1sKLNLAbtJc0LRwK2U6y+U2J+6sLye1B04M
lXMhMGLwvPuyCwsNX0wC0bgLkWNOpPKkeITD6xBt+Pv1cNwXVMEEdRxt95zArkAa
v3mlvm702dYfBeIJKXwDXIoxbRmrXsCaxWuwHvMIoU3IFox6bx3gwpG4+PEKB1yF
+WD8jVpcIkpBS9GhVAbT/eG8MW3G6879DOjceTLJWdZyhv8yjrZy6bsde07YGFnI
RowIdRMJzW+ZgCH6cc998aAIdFVetjEbzGzIPD06WPIpDpOIacHcicygt7qzRm1a
5wbPA2kQn3Rjw0+MfewH0GFxSWTi/WceuWh2CIf6+xSWcBNyDhwW8asDxde+5XLe
RIAn+j1Hh35tiqDwpgo6+BVRUttPtYtAaDP080GeWlMD1LtM2WAj7lfXtxQ6Oxhp
+vFI5TNtvvCh0T9sxXRdQCKyIUMzxaMIWsehWCy78rGHU0agaRBzuwNnF4QBV38u
gppiHZYZ4zzCmE8DSU+ibm/IvhqsLN68jHtQFOXJxXgCnGFYRbPMItPUb7LFPTPG
gtFapD95pbPQwvN3Jh0L+Oa5ile6u5a4Nb4t5Nm6+e26K1g983UafDg0KAOYk2Td
TAaImQpk885r//WP8GCi5TsjV38iCrYVdgNPTRm8j/+pZZJah/dOkTpCmZMYx2fY
3XnFlFV9jnoxjiAgcEInFRBMfWGa0WVin6WERyibps0uP3x0AX61voSc/k5UQEFr
GMnAVUnzFYExqA9lcxqwo34t7QrisASCmxZggJ0u53JmjGSaIm6p4dQ9We6jpnNc
zunTlePxuQWfl5WFXCaXibt03dfIaTBfc5tz2jN5GRknnOwyN4TQUflzWoIWirre
8Eq0X9A9hz9UfMHq/E5+oDw3tgH9iG2FwGtqOYzp66h80Q9EtA6gUsVJFtWjOsKi
lm9kuKatcozbo62NC0oXZ2vLjYOaNKQxRtjS83GZ//0uZbNuecc9T7mTytoHsVwW
5F/dXA6brHUptavlgpNU9XV+WY647eUghqw6TYpal2Fewmw3fD6shcBcgfjN4tiJ
EQO78Q4xGnwFjvhuNFX/pbC7znt2OQTGG4OFk7YPgPhDHMvUI2GqYVFRoyvJ+n1H
ZDwrpH+qXPXkQbv8Ii4jkkj+PQAnUN55BknMdF0uehnwbkq4KLomyQOsv2EpNKSW
oN9esK52Fb8lFd4HDkiBMtkzqFxcjXJGrLXPzXHYLRVA4ZDodiP6e2tjitri7QcP
S993e/Fgz9v6eAx8+S4qTfcKnPsDbzQSRT55DnrEAHr3w+Q5IhRiUoAGPZteTNC0
F9tMXruNHdTtKL+Hz0ZjrVP8c8PnAiFM5oOH+AiOWuLZhMDd4fzghQX8SLkjdJMV
z8KcUNcNUIQfRIRfRvop9kAyPfa2+nyzMD2FAU7wRiKBEaay+GNADSFE+Py8o1g/
Mf2e8ZS2d04IDheFUMceqedUOLV+VoLYsSfLmr4Wdi6pBr6F952He5XdVMsoKeiq
OS7DpSmv2G3eWPUYdHSFdZODcZf3kvyQG8kdah30PMAkJDUaEgXY5beg4yQfAIPI
yYT/jSSVtnO0sNJZIHrgMQ/Z7i55Rn7N/1oa5MwhiClf1yXcqsZOhVs4SqdDE6qQ
U4RFx11eGlBfaA7/Of36WTVN8veJvBcuT/IdH5a6s+Hqd2r2uW3KrW+hZDG10/bM
g8YKJ62llesW821+dISZpHff25sEkD2mrYoD5ZCWFYZbGvvjfLb9VEqXOmXR8h5m
RLRn0tF7AvduH8fCUBX0UteVXNFFzvMxLcerD9Tax/bLLWBwfHusW1TdnLO741O9
FRzr5jo9AHDjUsQ/SLzrWbyqGEp7A++eIQq1R3MymqvAspzUfi6G9qAUjpzSRDAn
0y2DXa57DAZXjJRbKnKd5ruXEQrxjwP4XNz6oFlQbktlEPEOzfwFX9+ixM6e3ccH
uIGHarny7u5HeHGvTz0NaD/pw1qAQJnT5TcIKvWdez7Se0q5UrANdaFQ1MKbnIKM
htltJpxAwsCTRcNl/fU1bqjOyOjF46An1W8eJHchTgGP1uZTVX4TJcajFKdHnbGC
ueMFqEKtMq8h0ji488RmHVRSDuD++Yz2AyQ5w0CZwtLty+x/rYEszPEoSxe4v/xf
JfUVPRsj0thHEEr4mL93qdyN+OGdbztJLJxBvxjhDRV6sNUJS8ljs3rwfYrxoVVV
aDddT3CUQ5Km6wZPa8oJqBUJ3XvwVbB8jotAWKAvv8Omy7f6/isjJCoLHNIO4XuW
XCt0a16T44ss3MqdZRtI1entvemFRIHVSGT7QObhZtflmHjDniGTf4yVphqNh7Yi
nChnkevUwoMrfMoHHOrqG1qZUGiYXMfRhMhTM5ZCVyjmmNKSwfEpCNQULQIMIkd4
ERCk4FLdsw0l5/nWWe85UgzdJUU3U8a/13MMQoHLUX2fCNmYicwN3P780YdihWsj
PIOvuxfnE+vN48Y3zaHdoJXXrHyWoDpWfKW7GP6DpDW+0cadOwUVwkcJmizN4JBa
6yera9Fi3WYm3XH8j5rC88r7Q200zWuxp7RxZ9rNam1WVnYOuAitcW11tksYFd2o
vm05FjoJ1bzP/fGDfIn5CoWUftJPg3iJjLhQp990i63+N81wEK/0FhrynfFLKEpw
nmMqBIvgw6YKgOKmVitu3bx8ix+dsmVyUIefZ4tVf4ZmENjBnDjjzgNeMw/DnRf9
WOWFR0FAetv7wTzK/tvpWrgl0DwmHyTBZ99Pnhb7Zm7UmmJLt2Ri5ruN8AFatzVF
qDOj9ZKZKStupJV/duZ8F4wuabCY6DxBY9SuzOp8OzTOI/C9994CWnxkbrE+f8hx
5eZcu81diVrZW3mfjNcxgEYJYPasSMjwXzXQVD0/c4uy8A4rG2QguFIgODNxuArT
YyrC2UUyGDIlhq9ChRTs2/izhIKjKnV6MOD+VaDBfM9jZAhkVxYnpcmFynZrMzzG
QteZZVN8kd7Ag0nZJaxS0kmtvvXBZUYaPNq7+THzO8ajjJHCfa4B8m2cIeLK4Xqp
VsQS2/pddrhL6f2+DRg3AKmqKV7sau203hc2iIkIjWbCxpfenQyQ2kHZ2InrYa2w
xWW34dr8OzHOmmTDDxyPNX7fJ+Q79F7DRtiqT28PmGFXZ8wlL2S+BGg/YVvV8v2p
YjOkDwKEByr6RrPcB9j0og3BRGHLN9qfQ1mvKhZqIM6QapLo7Tg8OkkdprgJ7mm/
0mO2nXXdXFtkEmuoC2Ql8oSyQE4TRra0rDUlRo6QbbZMptFhQpWE/vIGrQz+AW4e
/UbhgJm4ANjEtCIeYrVbDFpK1l6J5Z1jAN8pp85Risgnrq4FQcXgfJh7LBEYo6vA
sABKRTQZz5INEqb2pNR9duAkT/PeyzqcgRfRlLX6qrNftLA3DXDUcRGkSqLighk+
pl6zNcKEH0LiSpH2x9eSaAXkwlmT4H0XHYrKdMr/w8KCwBaTwpdx23XKhndtY6jk
dKx0EvUq9QpkkjtHAyXYtIZco8Nc/9FHjJXaptc7VuYtCN/WCjJSYZaLmMlsU5MP
AlCCA4fopVfEJuIpg6Uzva1xcXhnolBD4NPqh2Cjofh6WKdbHky34YknAciUp6I5
q0FStcdzQel9oKvrWBcB617aBnKWKCIl7PIoF1d22IWJL/4nVsVZcYhOUVjEWu9D
vzK0odJaoBkD3Fne2de1tUK8ivP0jg+U5LBKATqOfc3EWgZXktgslHqIoetMFvp7
FsBsaChCe2Hz71UBDh4r5izYr+vooPIyfRaLyW4L+hEH5z++QFzddO3MLtg6B6Nm
IbmLAhSRDz7xNsEdZleynLwqJN6x7Szc9zwYPY/5oIrMELUfu4XRZdTbcrPgBW/o
ZbOyFHqPuS9nLQSWjysq3O41BH+X9zBsV60KnEZyjyQ/JQxKnTYP2FI18NEgYrdz
YTtFX/IhwQE9YPGno2y05Hg56Pfk8xwPL3n8m9qjMltMhZVU2suqkyYYjONdjjNe
bmFMrs+Cwyb+f+0EYTchHSvtDwLHSD64ug+LLKbH7WaqEO79X03NwibR+AcBvdvg
5WNaadVCBJg+K4TDGVaXcqM98allEYny6Vryl1W3c0UpBNwsblrnew7ljOVlxLcD
iZE+2PjIHxkPaLFJf2Sy48L4mn6T9hnrKCTDMUDIvcmirEqSuA0IMxWnTJt2dsvp
Z2q7plODzd3XJLUS2oYAzew4Ri4rvzA4m7cTCNoWgoyhFpjS+cz+bWCM+/BqkR/A
0hf7DKaTeZ6g2UHJRZSpKXpdYe9Yi4V+wA/1M0HC7sIfMR+pd6mQilgngz5oJtMb
faxWzIu0V6yDgLVJ/QRbefxpMDyEGcxdtElhFgZdmK1uX0FXkZRZ6a+df1P0MejC
hgwZMptXWO+vDWLkJxBbtYs+Uop66RBnMtoHZLXcilV2of3AGRNxxvccB7FuXpqI
AiudqK2aqWf7AOMUlvTMFoLflztVRiIZ+8NJwwozkLoW3AUzdCEJYks72Ybv/0Tq
Kqh9DS9PByYE19OgCJGMRTpieEsIyllB3nVmDBVjB3LAYh/TZKRDBz+eb+Jnc/bq
mCKe35F1C36A/iqVFMOaV5EiX6V8d6LWI4L32XVvdU38v0WhWd4rWBX+g7MwLZ59
oFE/rUy5Q8MaHkHKfa+rPzXq2maEVAh/3AifYjDbqQ4jxtlka3mge04fsvPfmarC
gWR/Znj9mUpSsv+WEQMJ7wSh3RnhMxekDlKyi/cJKYvJq0yu/RtJEKri4bLhLZyD
el+BJ210350OjL/zJ07uHXFza8PazeNWnTB+ooawRn4YbZfGvOnBklpuqfiABxv8
dVxllhclDUCi9UYFUTGf33g7xd8s4u6X7yo857iMGcnBigJJftuYuPIVQg2DsZ2h
Nce4vpgrKnsV3gZNp4QmJ4Vh9nTPHrFiASVkO9Ma/IGvgEthMgsutgJ6L2U6qIJw
lzZvGEaCqEMjuNVwiVeUv7cMPxJ7smO4Bk8p5sNcIdulbOEMK6kzYmGJqBomzGl/
826zPyj7EisnfaiucwVfgbWW8KI9iVEZ0zxuzHIY8Q3WpCwN2clJgIr2I7pvRhYZ
mfjW5DrD+LAvJohujTpl6U68ShmuALm1tCFOYKR4r9n0ooM2I/ZPfSWCF9w5Dl/g
bOO6wMNU+jUum9GEBE4yOo4kwLLIKSFSSdrh608fESZDNCEjIShs3r1G8GdW2qbx
iN6E5XUSX2cWNILgiTRSiJJuMqIArmG9yNGUFxhQ8NebzUCiCe2HgxyCO/Vd4oMu
JRaD/qlEiWYjuj6UNQai5+m2l9GtBZg2UCXUONLNGPZnmWGcIibZKZ/01GoC0E4C
yODpne1SORHUOfs+inD97+fs/0mw0MMPuyB+VztYXLRL0+caPHBf2DHZpkU0Q2FO
eO3CFBPOEfeIRCEBHxNPb0A9U21YmFYjiLqZmDzxbUIE3igvOd4UzzSihg9I8FnT
KRbV9W9lGe8cxFTzyl3C1WTJebVd4ctYF9Wc0FjRhwEX0EaF6dePSeTqxo9opX7I
caN79PFFdYAYVaOTIuJfUMbJYGUbcKG+YxqxjgT9TaBrSisnEs12DswWtXtReDFi
t5DkUjl4mRaYETnOpVA3/KrttkY8OefF5l0Jg5YPopPFaDchEuZduduAKzNWlj1j
/4+VvrxrJ2mUilEFPK04VLF1piV+tTjlME8/mY8IaYxXzKj4bRP1mNbGIa42q+Ql
upMvYdoukgYCFLt5/y9w1jprLQOAzi1eHQYefzWIma41bsRayeewrOB1Xl1NqU4l
65wTIOphgrvRM7gwocgJDyDWaFYaYnk6tz9cn/ryunqNZfCB00HPaRi/6GAPdTON
zPwX6OyYq7xy7d9CgLYPXQEu4UFGf/k0jXQ/aG6jokJys5MSJgvPuWidg/7BYu5D
zZ/pEa26wRlsJF7tPTFQgOM4qlyivnLhSVc8X/Hwl5AVDY9ZabSiNrncrwRtvz5q
hlpkln5iVWk11aPdx8QoTl2Kv7w9L1cXS6brrLt6JkWDIPZwRtOLysTY++DTKBya
ehZkBs6quGA7+PvzraEe1HnsGwFh/qOsSkTp9ttqE+D0Mc4qk6qra+QghiJcQ3FJ
LxutefnPvlFgQXAa+2JUwfWYL425+t/x0MlfxU5BpTj+jq3xojuET3JnEklucP93
Xr7lSAnuMkf2bq2ypHhDWaLp6hP3i+Hjki6TFl4hE6De0afC6uwtEpBRiFABS2mQ
t478RcRc4o/EBZ+5Yc5zS7P6Ij70PlrS168wY9gbMJ1E7WnWm0hjdEouTHIxbACV
8BaYjqsE6hBWB2IuhOnZcKMbuPb+LU7MMSbA6fjHpfwJq6Fn37o3Ts5vLiouU7UE
HHjTz1ZOfw4FpJmZQsLdAiaZoZSD5+NJr2jXrF7e0pnEdEv26/5LT2cXHZ4PLkLl
gn44hSF+FjcvzQPZe8kgLJpK/O/lD1FD3jXacz0TGEDPjn4VYPcVYNAV8HY9kpsG
6eB/DxpOphm2QM3Z4mooKQuV7RF9ehX+ccc+4HmADU0ZobY3XnkaA/GEhYBbTwjg
L8HhFJgkDRjC0C1lDiDt9/QlB7/NsXVKtCOknt2oRxEdjgE+M2y2WuzkeeOm87OZ
1eBIYD4kroJa9zntYXocfmS0w2KIndi8ASyqzU2SiX0xwrfsES9et5TzisT+3dj7
Jqb52Zm6ZICKf4v0+1Mp5iJtjnBRCQ6/EbdK0kLiFLSllKdaFd4texREWIoIV7/i
RqAcHx0JxD0m6JkIeKPfgY5YfgDuMgM+TVVt256dE2BdayOaq6voizMOFtDRVeyj
sWpd8kn4t+LBYDpK00E/sRVQ01MAvtxATuCmTSA9dTaearF6RRWPgE69ku37IJHX
W92R8SBOf2HilwFrch77hv/x7d2DyvYExdI3ZJFoOiAQvQcfRPWBcmK0G60lgR1y
3kBolGkL7T77wtC+dfn+9n1H77pQDf0HaESvlKMxKCMg7u7T2GCZBe8hzEeFPq2N
wFUobmsvIjiDUSDG3L3Om4I7bSYTX6ObS8YTY5/hLDjwRqT+ySDT8NiyKB2Q3D0c
4Bbjzu9nxmmhsr/ae5PF0ApO1Tz9rslwDE09RjDrdPtWzuN9xwJYrkNC9PvxuZm7
TF8nb7jGxlBM/wDjLzA0DVoGRzzu6GdOxKhC1hgkgz9DTdrVA3vYoIQ6F/CbPecq
h9vBEQDPB7D0w6+BNGKziFGOYKbGwkn39sUdevabAps+AD4y825cHaeG7aqACX15
asySozs0UaxllTHyuzZ4RJyrBPuCum7GmrwdcMBUI7plp3tMzrw4jtjp7Rulyxz3
jwrWYo0QSUW4NJ4ndMTr5HL8VgaJ1TH5CSLfcmzroGopqNCBsn3HmcZGtYxdXwK0
Wtjh+2Y4xWinYUYlndguiRey8hSc0rzepYbo8ld0F5sek3QWM0hMdQREGWcTbi77
2MF+xI0ZMZSVXLxQtnXzLfO3/yzu1PGtMvlq2xuXom+nzzPZwPr3zGKekMAYxxyk
UkKB52mgRdXBa12VaFxzg4vFQq6sZS8VMicilfnmm6WfeSJvgGpVR4N36vJbiR/a
0EOJsyTtS0EkVj8OXtqhccWqmUQ5VCuEBN9rClmqSJhPP7mVe4BFaczTF/60FcGn
hpNHAATcf9Qa6xVtkUeGyya81029PdlKjYRdaJISyoo6P11828uH6FUvvKYtASPz
ex48ry0gFybpgYIwgtd23OCL9Y/ZJu3t1OID88upBSpXT4IgTSENQJePEEQ23KII
FEZYG6EPCGzz6h/qNXa2mc/+bVudAbRYWK+6Q935qCtBsbG6nypUmAWiCr8KEaWm
qHhlhaX/X7yIURRVUHcNCMHzDWgW0y/7LzF+F1nM486TEIn7jo6md27q73573waS
JG9AprdnbWSZldrN18Zgpk4WimUr4E4oS9tC9LezKlNW2yrufkGgbZbEJSdKDpkl
nsoBhUK9Ee6+21Iioc2A37Vt8LdOyjMNbkQrtTYcjFGsO2Km+2vQB5h11WxouNYc
wSKp8Xmpwl929pe/Vt8lo8+hSbtrI9QBlhH2frp9BOGC0UpGyVJ0IqkkwPKD2Diz
QbbbCKE0fKIZ2154fbEiWA75NfwBzw+PHlajP6KPC0+Ua0sRE+fWLdDAd8lJ6dgj
jYt7mwSty/pqQCIqszeGX18DmZEtjUd+xhi532hCJ83p0c1ceS5yHccON8lL19a8
jGWqlpC3AxY2WYEvdqDSmhprVhMAhk0Y8eD/5bEY9QxX3U7Xtb/3VN72Cc0LWJxK
OhyANmbbtM0I8NFwlQkO+GytLgrcQjvnQBui6Sp0KaUdJp/c2wAxdUHTV3OZaXzZ
h8YEjnawzsND3u4Eawvx+kn3wkf0YwkwydvAdiG0yEYXX14BwMvj17CQMyDhmbqD
Id3N1sIKdNOUVfq5MwDp3975jQoFtBHHi/XZNbHk0aZMasKLFVG9qJvnBV6aLJAR
BrkB+IB72J6rpoytfay7DuoAeTiUwbtWg9VlGOClI+jlz7BqrZ8FOfAhHpHz96ph
Hzz2H+dtQkB6Na7nqCjtg4JK5NSrOFJnT6t3gl8EODs2DUa1vi6dfDMlAxr5kRFg
dlneHQOeFO/aUPSh6h96o4/xeCO52z8y5eMS+QATZZl8ORKZF/e+6EAkf8Oyh2Pu
QjX/PFkRecco3plFxOrIL8GTBbtWxuJn/Y7eOL949I2HlWrHlOtb5dz7EBUAh42c
VYYFnHx8X5JmV6s98G/w27WFc/mDySc5oJo2omOlTZDtuMLuYDLSdlDhw8YdYHlv
/n/xvDbJmGfTWPggwhzIytY52RLGY8VZL0p6R6xobV+QARZ/5xXCMr0fiq5MlPOg
7Q5JxV4envfCoSi72Gr8Scjfzg3VD3ua4gtAS7F8jXOKiU3Ijdb/zFesmFaNPKZe
KbGf7f1GAHALDIjSqhTOqoVOji3IXzkpOMk+nSNgvKiqUWTaaCvUcVfQ/vIA1jHj
GKCf44o0GOl6ONjJvE9kMvdD/Ubveibgab29IXUoT5olhYRwKVhCl54zqmNhdb9w
pW4CXYsM8hXB16aNhu2oiEtk5nYSHLb01JywiBhKQ0riUM+MSXr/9H0AjNHSS3tJ
7LGiM1a1cSTYHO9/RpNaD6ECgHjh4og1cw/4ZfHT4KdPL2DayKWij6tmTIyuAZSI
XRzHsg3zMAIY72qo+NOEoWZFX9ZDdZmCsWxukngbaAlzoeXosojGr+w9frdk7uTQ
eUhUP9RPXOMAnabTgwlh0Jr0552ukOL+hwciX/JcHp3g8WDUvahHtPalfpzP+gSE
Wlp7zpBsFFemTkdravDtoG+HtDsh/o7HoSoEOROshMiMzR5Bu96eBGo3+yv0sx7z
cDT8eRKB18ZSZa4FkIwdWQuQ1CfK5/4AnpcfAh3KojOdEUW5fM4vCh1fkG85oOom
lFhnC3diRiDEbh4OPoCNbUxuVTomJm5LLH9QCnvHmnj6twezQ2JpExesHyKuCTDW
gkeFGG+zrnydUqrsbG+LJvhG/+DJ9k9ezzdsuJFwAxwlkG1PUnoez+msHGhl4YXZ
o0nflSybXYlAQ8z2Nv+Eu5LsMoRgZN9URFTUVbL+KRtCA4Dv1Dr8bwg8O+NwZzle
fowwbiq0U93o7L7zH3KIK4oVUZQWqFsPLc2hDCTwJGIdq5/iQWpRUaE1iwMCRxOA
70BE7o55bPtLmNGuZIcBspmgesQbStTkA/F5ktI/4Z/2NNzfxZYEgKXi5S37zgqN
/tBE83eVBQOdKHrnUQP0NE6REno+x/OyEE1NwebfVGWYqEPQQeUdtOipngcpI7bB
XT9W6F2+fgn3HQEGXFCZrwul3tCyMFGkQ4DE6l5fRdJKmiFZoVA1UFRsUdg3sand
Y2LGSJFzbbSyspwAKNPfXgk8nJqUqg5u+4CVk+irWpAqBnKWytHNNaCEEAvRObQp
Yso4BwZLpBOFcrhe/XGnO7gTrFHwAjr8HI3Zpo3sSG4EobcmD+niSIxXeFVS+rmB
ksiedfSqKQwIG5L+gGok+knpSThyX1TnxnEpVvsvovvgpy9k9WLixy4/SZsPW4D0
8bC3JJQ6dRYgQh3pv2/JzOg+SO8WUqUcS5d0wuuf60C2pZCAZoBJ63b7uL/62GsC
D5YF7nOmcMbKWGRz5P5A0x5B9rt1F7gkIFGk6xuYHG5Zwzm1QADEU2o8lR4mj8vY
PusNrbN53WAMQptHiJ9YD2s0kGpk0Jp+BAHiPRSiuw3YQwp4z7BplyjlEPJSSd9z
uQLH7KiJfg6PWQtlNu2vtdj7pCY6Q0Nf4eDUvOa1aE1P4UBMMC3Qpe4HUgdkA57H
5/+YtTbk7EzF2yD1xWC+yYvEctVfOc2omZdrG8QXQicFz9783UG/2XB4FuVBfA2s
bi590G7iUZ4hdDzq6POrqBWU5ncMqgcyjfsnP5R9lkM8IjAPAOti72oH43kKAaB+
vcYkryrXHsj1hl0d6Equ0vzobwShAINtYRiyhb7J8SOLiOMKBF5znjcHbzV9ZwFj
KGI7XUpiA69NQW9m35xodDiXwS66qest9tDmkenNKXo/veCwbqAjWa2PHBZqHuLH
buF5qJwz3i1DWv6s8DeoqMBWgB9HfKNpnCXpdu6EKOHrXQLRCWSvID/bwrluwNjS
GlOFYA62i0IKXCYSATIu8DXTtkmgKT848GJs4d10uOl4NacgwqUGIb/cAJPb3vkm
2pFe4r/P9B5Pvd8MafkOjt+ZESDj4BGnRJmF/ahm4+TFzmWvl+JA+V3M24JNRukw
pcDqB5ti/9Y8SiU/FdEsOCcmOJMVO2/9A/0xIU6Qh9TElqw4lyZNcWYiG5VLytoF
RwK0coc8466U/eG7VPZ1U5J6/KFSva6Z/yGtK9mi5UtboQnx9K8TGBg4+Z+hH4i9
/1Aqp112cBG44gqq7lkYNBXFPld1wP1SPGp6R4FPZt2Eleum5VnkTt13aHSm9zCE
cU92Iyr1iWTH56z0/bhil+3XbNa2z3cMS3xlUXRsmhSyCE60s4k23FeBCi29wIAy
Z8SxtFMy+y5nT1DVRcE6l9N2a4BKKn8fyV5qyyivSyNfKpRnhZ67ma2Vj42z9jr9
ZefRUHSnnlMiJAju72E2jVNiGdIV1a2AGzeGXtXSyvyfXD8fnuV+YGfCDbhiKzfG
v0+aw5QS9g39yJDMDjkmbCN/B1GSzwxzFzBdNXiIgRoIb2TEEXuER0mB8pZRZrAV
e8+z96IDVnjU1g1SaXiQnlbekRnHqRVQiknCTetzJ0zHViNOCL/ZbgDcwbyi1ypD
DM9/BQrZaca1517rKk6tsAGwBN+9A4oQwe7PuSuvOpWmJVW0e9P5eQw3vYpbVljd
ToyVpMdxByn1h9wXZ7Sl7nNdb9J2xbfu467kOo3aItbNleTUrk5cFY4YBPJ7zq3n
/hNB+XS9zC1WVQbSVNU8BLy/WaBHE+eN7uL1/sCTxvnFr0npPgZNF9izNEubrESq
pYoJsfQsfmHVgF3GicnmJ3GWceiiZPZt/ZLA2adM7zo7hVm/X1fwx5Dr/9w54JTb
+mDK9lS3G4X/YcrWZIJ1iCGEGtx/2ALXYI2H3iPPae4/uE4kbuhMEHX7oojpH61I
j8MdO44SXtlR7hkQ4zQJQ0jLSNzDjTtw2pMjwUId++5I8VYEASwyemEl02E26Klm
84EHPp8+zsJ65Iim5+qgPRNUR89K/RIxxC/xKdnvlgGeuoemJH8xXO00I8GVeLNA
8fdMY1WQ5gfkSWH0MiuAIyanCxWzoo2ZGv/APxzX1gxD8Eq74dtjBH7zwgOx8qyz
tw2N+cN/LVafDZhMhBLZF4mGXo8ZkN0igO/6tNlDmGU9F6dHjTlNvC2lNhTp/y1e
`protect END_PROTECTED
