`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H112RhV+zEZt1NetGVyl0h9Lo1HmLvgKpdxup5Vet1oh4CIcAMKuEvqGk1VsBpY9
N0KIGxbXtSrDZJbrp3djSSq7AE9/8IkmKovBxPFJawteyi42+TBfT13wF+Vvkjnv
N2avf00OCb2rltSFggPUhqHm5TkkHIT9FJ5NtJbUn9egHX30nnIkLCLVXdNuYTJn
+T8YD9Dt+3nL7zY+jiANv/63sT+40PAcuOSkbwKVOUlF8eKDeAssEUnuU4WwIOur
25Fh2FcD7cU/x2kKknCdujLC/yUCuz/kEh4GWSI70RoFAB5HAkuZAJnoeEELAom8
jbAspero2F1fSrOSIvQ5tfWkMRMDlXp0HeKb3uGSB+vmrT1KnL0KIL/KkwY8ZYfG
ZOJ3JkKm3CemAzBIaZ3emEStuISTkInyHkAyBij3PeyTBjonrTQatE5nYjaDqpvi
inwVwIN8znPKLIhZejiHFmth2PrUADM1LE6pNHESRvJHYsz/AiNhkOxbqsMaMIEb
6kGQu3OyjaJH5b6c19Hq6LeeFy4n0JJOmxak1hFP83p3t2swt8/JO7/YUH30LQOA
zGb4WQrj0Zbyn8884SZQtmeodXEYlrNSzLEUvfZ9VzI=
`protect END_PROTECTED
