`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UpEHGGHXJDvK4YueE8M7v1I2lvmMkbbXvbBS8L7HaDuBFK8poPDbgcpw4ZhAA5d2
enQJ1ZG4oUVurbFdgM/oYvqfHe8HJ7DLMsk807H2phmRw8Lr1sK4sThPt14Hctsk
6ZbNEQ+dzU+GvG/0tilPXZVF2xFqIS910bgWDvnw15K7Wt6HrXJ8FDAfGz76WQKR
NFQtQnuP5eyt7sR3YCljEiVKJsvzKUSy+ZpSwxkuUD+jIs8mhEBhIyHgellTf4xX
jUMBYj02UdE6+FJDddsIDaOpJU3L/k5aPYcfGM25K58iwEQ/+BlrztNLPNZUNqp2
2r+TvCZQqx9EdaQ9Xu1PbHioruB0HhKYDLzUT9ZjEi4AZ+03eiU29MLweWCSm7UC
BK9pvHOE6cL3syN3AU6LzAzivxEVLLJMRjsi6BJxY/Td2rX9Ba6UKDkaHiKdY1IF
LD+NoaAP9opJsCKzT4wLXk3WxKD8xHXUbSfX5YLAHevPPSkCvZhVcsR8zJAsYxPY
`protect END_PROTECTED
