`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDYOJ2NVK4vGqpDhp47BLWkvtD47tZoz7HKk2ISa05bL9Ro13vxYmgYqIA9Lp8TQ
QooM3GGA63dKpxDspDJIuMaQ6LJ0sz/C7eEbsVlC5ozgPjD22soeEnxvAXkI+Lt/
2hTt8SgS9uWmYrAvdb4TtTOyO4ASMLJaYUjrJGCeGLHE5+GgCHT4q8N8RKvW9JZm
XtwCkyIN0A4ZaHDGMGjV3YNkvDgsjWCrke//Y04UZfAu7fPlpiaja7a1sQwlPjKl
5ypGV4ttfTadaCpxFTHV2hIQdNvlFYzwIAPLhtUsKUkzcom3RWLjaMP7wPKb0hGK
qEq4bd9/mXkRNAygnMmd7V4IwDNpae7vPXs8q9K0W6oWcmPGoicQHkYe7o2kHVGG
cA1gkZt6C5Z+29gLPRbPytlZBpqL2UvKLog0VCc/WacGnsZgNxbShx5oLElqTiHa
R3/3271NKwolP5wFWEe0nujJCcgILq2n0bpk6Yg1i2mjNxpelOFafIDxHILgnFhX
Br8iIU2Xvz/nhPLMm5duLoOfdtALNQ9zpn8e10cwyHwyiAG27/0EGpa6IsH2uMzs
dSKvzAWLCBDwmSeAdG0wxEcERPoN86TX89oBCT4rL0SmLzroNWSLu7pgLeXAmxhg
brT+vWnuYHZWggTSjmutL3+r0n06NCr45TughzcRE0ViegBubSBO3zJUuJ4A2hjM
efWGtzsCq/xmZezybFOsz8WWadbHBxe7pdouLcDqF4n9Nwb2DvY00wM/KQhQ6UER
CRwp9i6v5IC3+5q8C2P7CDFouPtQo0oQjZiJLU7uXxIYZ7AICqtkubFfjVEoTY89
APbYbtieHLNZvN/YSj6Y2sOGBucOa4aHiCWDLF+UkootdQKdqSUNoGKlg6x5yhyE
/+Lfaz1MIhDZIDtVMDHK1tlf2E0jHNioHAhN5+k23tlXn6FZzC5eXG1u46Y9vFQu
32Ro6ThWizmrQ3zrVKv6IoQcCw5o9KTVlTy3Wdzi0eHJq6abD9jceGRScokLlaoP
/zGtw9LvP31Z4WOXPKNaCOEY9JwyUgsWlGd0MxC++QfPSxvAY6e4myP5H2+SC8Bp
8mXMpJSVi+SQ5L6okfwCEC+FJOeLqnH7J8mbVYkGJtKeGzpKX/9+WuGO15rfqB59
wpNaWjaQ4jeYCX1+EUdkBfw29k5j4OHTLHO5i2Ghoh2uEzlhSRlg2u8SO8R8jc8J
MekcFn8GCKdI+8pZ+HN9w7xCqwGyCCeiXn/lorGXUVf4CkEYZ6hfPz+AtQQPGOxz
X2CKph7YvTOwcgHaoU4jtAxD48an+xwHqURjXuii8Lvum9RBa23/eac1xI3jtzJ7
T++3D3FUTkPw7RnO6copBPduJgtKogoZotjO50ARoFKfiwncS9z28fAriiYBT816
LjqKjQ1jHyMEDWO0c8Y7xmxuSHsKZf5O50ypUvypLlXBFtD8icXnYuXX+dwUIXL4
V+OTkC1QcKFnUXgLc66lkCoe0FxM71v8PhHaF6d6dno/aTV68yezF8CBIVkqwoWD
`protect END_PROTECTED
