`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6NczNxK1jD4JRNvhEyNsrvotCTqqoVYP198X4WEOK5+TDzK/dxHJZuAbbW/O5QS
1dmcg5H+q4pwJP5/8Tarh83gqnS7IXxBX5rn5Sw6IDdv1anPOckif/oQC5wB24YH
ilrMNQhBwpA/a626eoBqCfEHIW80z2f7La/DU2i/3Hbr2xd+TOXbCZI09Qx0cUTJ
xyekb6eWtTpdphK6T9w3h/9pINqoS4ikMkDklOcPTAcVK2HaEKLU/fGC1woOPoc0
vED9woKopXB/1t0H08rHiqO3MuwrLkSGHjA2WSyUz4CDIz7qe5MeWdb4xhUKwCFe
jKkn3KBqfi9xtmpeQ3qv1rNbB2O06r9X/tEmljGv7XETQZTcqAcDvNqdm/Gjyo1E
kdSeOtVJYRbV+Th3Lz4uc4s7NvNL8V2JNtylvmRjYSZos0jU1xWJQLXFJkR/+V5P
uIrQ98Ot/LeksgPQ1WHlA1VHHTc3g2kW+M4SiCsfeTU1mg6sPSV9dfMjEke9kXFn
ASP1ziVBQIH9dm/KuXwcfiQL2ghfqNXAFfFF3TC/6am+znXFvx1hnAi2VB4Kxn6G
oJhmThYhARPuP0U/SLM3IyjU26ystOGLgyklNrjBRXnSk2vkTx3g3ixOS/+L0Gqd
gG9gDwotycWgCoJX6dAQl+4VDIXcKCcTyedhS+ETETIB2bCruqtSTn1w31oBllX5
U7sOYDI3yMzNLJUTWXgZ8fGhX2euEBRuK8tDvDClXQpBSRPdnY4ul6di6c8fWnOk
oXw1rDrqIm094L8sKN8fPqXjzGdVVxK9MXBYKgiiJY7upU0MOqKrLm55Z4zodqBC
jjUdRswBMdnU+EpEVODqLakzJVffhJ1ASOI7JPwsSp8HJE/pRaMXp/m2XFjT6vrK
QPp7cAShBBA4pPQEULLPt0xBTo3Vr5Qe9KIt80Vctt9OzOXH2FuG8jLKkbYzFPSF
`protect END_PROTECTED
