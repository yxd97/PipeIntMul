`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjxOIp3/mOjquO6bIoC27l+2+wM4DAhN7SXtglkKdqtwwyBcUSXpB/sBeJsfJOEP
g9hA06lp+e80PW8PlQQMpQpj6QkwFB38syVJlx98jNqh8P8eE6NOMWd8scnh0GNU
PNZX6jsZ+dE87n07B8Ci9o8GeaXsIKD6HlXzfI/klR1j1LRXY0IHBK5dZSEwnesK
FRNlaXnU3y3PamslP/zI2C2AFgT7cSEkvX465Q0QexnlW2oZBrHaKp9pBPE6/AnC
gUf+AEu++MLQuati8tL/7jmMGJwVKLW3PgRTpwlJOfuxofdPM2sIolTNligUyg5P
K32HnOaiZidbM6rEGz2VrkdN8B6hl1Se42unIwX1GUdjXAAxaNowvueDwTpxzyiI
b4UYYoiPVCxUWzyuaDa4JqL6iBLkrswGlt+d/YEArxw=
`protect END_PROTECTED
