`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x36EztH5VaEeMRqZNqnn/V2lechHGLPy9uz0CIH3t/+q1V5OnkwU1OwCshG6o6DJ
BoJUvnXXuefUQDPEmlvuCZigfLEs5L8C/PB46tpO7tyXSenUwnmRiOtrZukrmsCR
AUxMy2rD/4Z/lTBxAtVtDoVMMcd7UqEnlXFLxyfiS7kl6UfAefCaxznyB8VQ6d3Q
wVJubBwW6vFU1Q99kIWeQ4rQpBUJp1wLgFlq8mDFa69b/DWcN2neFyL9z3dHk+Xl
ytnBV2prboyeurhMBtpGeHByfZFCV7H6GYZyu8NFGtUWKEkDh2NoWF0DW3Rc/1Df
wZn+0sHCSS2cX9MvcEal6A==
`protect END_PROTECTED
