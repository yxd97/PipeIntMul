`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tKfnRLhRzTF6dWyIExnO0TIAnVbc0a4ZGjwd90SMVpOHNFHhlLtQKKZFVZxnJANY
BCrvHjuOn0aqoWSR+HzsTK20SpffaPptW9MO5Z4VLFK7DsLigUpYOpESQuPZ9BN4
y4TrAQ97eo7l6owTyZuynG+A1aITR/DvhHTuIHfr54qvLPra4wVyJtjNAdrWxruY
n1MjRXeQ0PJPHuF1wsQ4dnyIymh1tZuXqIP4F80pYPvz+X9Gkc7mYARfOiiize0M
CUG79gvr6ARLYwRktlAUI/CR6UfCnsLvRhfNfRzg4eNOsuDpDVKs0Pls9INKiA5N
t44PmC1q6f4co7iaphfuk4OtmoSAy4k3jwouTLJAWjXRExqZDty/gW9ev1xrAaZC
6TUX5wKv8jd0mLetL/sp1R58JnOngJcL4WV+PCWexY0xaTZ0dL4f81x44JD1j9zJ
opxPtWpd9BuO+LfkVf7xTtAa946Qii7bqcKLz/S+O/Lk/fqIYaQ8ohPntSDfcTdl
`protect END_PROTECTED
