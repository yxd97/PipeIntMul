`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xTsdyedwmSq78U3SWCX3F5TS6qxR0SJvoagVLM/FYL/blR5eGG4Xce7Ck1QyX0fG
b5vv1q2iFC058M7b7LDd/K9f8iiHmrABJw5YHYao43P/HQOG/EV2qXTH1s0zZhxk
QJ5xvmoMWghuwzf3dTjHW0UT0mGcLPeuuAMyCnFJqjjYcFnrd5fiAgC/mdi/+bdS
sSQsnniv7yaxZ+VCzPVv8CJlg0wNmceAa1j7jver9K53PWQtcr1nrj/H7RITTUTg
tYZoimbPMrwxrEJHn1sRoy5ZMVmnG2TqDvfWzRVvPiE=
`protect END_PROTECTED
