`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kW8tCQDfec46y/b9n3JLufRldjk4cfGnSqcCtF9gJeBEu601Y8WIjZCOfT0ARD/Q
WkVmuRdchvRcQRJPX076A5Wy1ljAGkoRtkhQWyKWk9LgQaB0dY6GF1FWPOVmOimv
DsEw4UD0+yrPm6akQpDflA9Lgu262D8SLOKiwm4VksI5nQpiOWEctmILdeGCbBK5
b7IZWRjf8s8kw0g0WwNXKszcM46gI4gh8qDjmMc2neRAh22S+nDymhXBgcO7sKC4
GwtZ6rfX7PUX/AqnOFaLujBl/iH5MUTTANA7TpGhqnqMVq8gVVRjDILRVOt/jhJU
hmEQS4WjPCJfDBvtn14o4w+0QfsJLYGqdv+ugk/1abkCsdWSjsnu84WVH9EQnDQ1
ByLYOMLBmg1TxS3MxsIu/P/uE018dSoH6IRLZ80aoctNhmSDYlTZ7qXKsbOXKb7B
xmB6hIoQjb325ti5AITZeKDNHUsEzD1dnEaVQbzr88yDNgmB3OgMtBAfBzhufAOs
QRugd9f4Uorb9T8VQXrwvOT8049qRhjlysJ+kULcobgmGqBWUHzU+m/L3qrn5iGe
Tb4+Aq1sJrlZA5phSYELE++mItx78/eG3n0y+KtbwYZuiybE++jU4sCp4NCx17PT
7LN4G6L56Yi6LSJMMjgD8UEGqAvAg2ne+zE/7I0yVR923HoynOOIVXESebqy8OiD
t5DfYtUtwTe2Dp5s8O6wa6w04MNrnz2wjIVcZy37Q4yjnLnTeocU7grR3/zyU7IS
tLB7CdjEAXWwhoVNLRrP/B2H7HgrjmrAoIHpuVTBra+pRqfKcATG/InVb4LWJt4Q
4L0rUQ0iD2/h33NbEi4tyiSTImI0YWFpFGoHUXX4OUo=
`protect END_PROTECTED
