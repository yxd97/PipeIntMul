`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41qF6lnJPXv8CTMX5V8EyL9g3Mc3nx6r8Cc+FORdIRwxWD9X5UQlhLVu+5ATiuf4
AAj2LWqUaTn/D9YGY161+/vn2gA/rPYaSStv23rFg1+o+nKKnxyLwsVhlQzDAQpo
rTrzYKZZJhqUTVUnJiUMAZ9zuIOS9EHKxubwet6H8uhYl6DvxxiYo8AABvfHozg2
N1YcsVSD6IJ3H4BgMr1nuzxHKovs8Ld8tAA9P5RLakjMbYI2rZ+WQUACiCp6wo9O
OTDcFajBqDgEdBzMz0Ft+lUks1XNt19nlRazLUQJ871pWxoe04IVkv9keu8jsSqS
cMABum4qfKMGclTLTXj6dPr2Wgx9PvcNBAtCMP/lg7v7B0L1mfrqXApVUWZYnwfa
zSGg/DkSehT9Fw+MaUBdaTw8RIt+yBjIMyoJYtSU2GGf+0kp3sWY09cdmqi4leCv
5/pHCYhrAuVZVHm+w125MQ==
`protect END_PROTECTED
