`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HkUiAUbtIE2WzS7+ehyO4KslUKBXW/1W5dUSvf0VTMf5PJP6snNUNBWsZililG2
yiRocYrkFcfH/ud4xTYdU8djnvP8/325T4z8oO7Uq0S+lxfE6JkqftezzsD4IDGk
Hg4lzHmSTUJz4245021MoFJsVgQbMq4nLNLAlkavG0tQZmozefJpXrG/3rN6Rfk0
AhoV/1rCrslK7NqpRqDOi/L9ayUySjYnqUGFRW/dC2SHe68rIwRJcAdOpseqRrLB
wk+lbFNo5DaGwmgEO7A7bPYD9/EbKbGp1RZsFnSVg8eSCZDDwTFb9QZuCHKuxVtk
OcUs1EjGUAlyXAHoIgl9gd58SJeRl5UEiKSXgLuVzZAetjFmMmhXwevB/lPQlgtH
pHSvc77PSTchmqowU90buhR6UlugANFykacmWolPye9kK0J0eAytae7kkK7gougz
p6MMGPz9DIVOReYbE7mqO50yft22YdpwQ9ANooPycfGUBSayzw3nVb8nA0Q+ZMj+
OEs3KHMVPR11FTLTwqkdIf4TOeL6DuaTNToxEmi1PXmuAATOqVY4/tgBTBguTafa
66FH1MONRWzqEKZtliEd/oXqbcGE2YuU7FpcWotkj/oA3XvuNLdcCIya2uptzfKK
+wjUmctZkj8M6DoYe14HGtc288fzDxIok0x95NpVwMaUPsOHBqcqUoLrxOtmrGol
CMhx263+PzmpF7v8Mo6HLyTsNOtlVkn9QkHR8Q2q7UBmpUNpQZHJ12ZYWJ2vBTpE
OFBQOKuc4PyHT/Ql8uu7dtdrfk4krX76T79NzjVh92JEfiW0uFCR15xIgWYwtY0y
3X8woh/dxMzITzQtv5JJpldKoV05j9WstmbNU0BzV9XboaL0cXWt7oVemNGGJTJQ
FIK7/psp8c0XOdF0zZiRE5VY+vFJ8GD5NtfS9LJI4BctfbJ99ARVrNHb9VyKlq1R
UwVe4c4DCyUTsdbsjrxCkhrfqMC17d06T7GXjyKpqM8jQTxCPEGsLLT7qjoIE11k
C7if/25LrMnCrrJS3d6AiEDLi4lH237PzV1ZPx3//0+FiukuoeGcvJ6kQLrjDqI5
nJAJdP0OfYwXmuTE42NZ5zgFmhD0UzmZMXLS54mAGG1A0/qJNLdS2XMMLl2ABdfd
Y3MO8JiVJlorcv804b6Fa/3zv2RpXwyrOERVHisGCOFeDqfNtxmIRKdV+mYfsILv
pdbD5t9+wgPvPkzVNKV3K7oHdkiPG8u/3RY+wK8nLsfFr6EhhxQRXuz7RWIXCej6
JBXANYZYrf4/uY8qoJEMpwRGrjG2ZHLpy5yUIIY2E5yAFB7sepxOvuseq77AsjWg
F9sxdEqbyN9Jvil83CeiWsf6bu8w/+IfH6kazc50ScEFf6AKO18pUxns4bHUqWVm
7GYEsVgF1DaABpnbzDCfEz4vUMNyqenhv2rqqGCb++g2483OlCcKUhxJM1scZ77p
FYMUHn2jHSqV3DRS3By2wXhrs0TU+J1bgQLkdcgKFpd0MA3LWVBTS5SlVdRnHMjI
CaC4+wq1lD1pTa2pXNJDOeUDKwLiDaj7E8s4ilFLdLHP/5QUr0wdbPynOF92bd8M
yauVNnAQesW1me8E1V2JLQUBAQkb10/pReyQCYX6brcMWzrcFLebjyqCxTwS5/vO
SUrJlTyfSLJmo/TYPkIQBXpNy280AHOjorygjuKNaFkdv1zACh/K8BFgJrnrCJsT
zBrFdDlQIq0w1ePdlU9B+cqGzFkBHnK30kZvAI+b3fzLaLOz7Piwhn7r1yH53iPh
m6tpjpNY9fh/LIhroY77yhnKvVNGxQQhwT+5crWswPp/zOpiMMYYSwDPv2NoRSZs
p5F4TGhuiciefSILAW3CVCoGTc0n0ihin/9qwkXUa1M3HQyYsTRFKHso0paJkvU1
dQOa9OVL/iaSQSEXnp5uqqg5H0mOWflDqGjChZ8X+e1Hof/Y3Vf18smbzDmmfiAl
TAO6MGaJhZihpTwhfqBL1pQDRLPosbEJH1dutQXzMen+aY9HftT3F820/TAB1vFj
GGYwc7TpVpQbD+XAiNy4MR2s6skn0/Dfj1wkKHo74BMgBl0ePHNkl804e4+3Clzm
jZUfW5+IK9++Uhz74fxind2KBkBD6EJvjDw5nOpPc8hwUs/FouflGDHfyg9RbKHP
/zolk6G1RNr1WrGdIpqCki1tSgls1KriP+E6u2skH/5WW5NYMCLCB7gbEbMnlabg
EOWDEg95pbsUAiLCifa/QMFdLSwQkBpnbr1QGRJdLJZCo8FcbHmP3/KXAwktQb2l
5eNQ2q6RmknJV8d9VBh22qtmfIwYWA2X1O4EHeSOggoHQHR7uj/7uo4axDbXKyqO
JMLFSZfksL7jc+hWMTPWum2NNVPw9Am/QAonzIFeWACyBlulyUk39GpuxXtksMhC
W59L9nsCg/jx9hjDcK+1zwZmmZbK94cwH4Akn2QZ9dePuIdlyak6f4BJQffy5Nck
VrcrLc6WR1R8XpoxOhY62MUqN2+NPQhl414jPL8kleaM9YhSY+SNxXyi6obIQQdR
aCzkVWQ7O7WW7VwlTBuUuSR5YHsx6axjLPnDTVD6aXTLjPRKM8fT2876S3XqVTPh
K/yz1QUvo/XZWCA5657V5/RFsj1n2bedxElHd0QcrP3ZGiX2dpxGZTE+cF4PZsLX
IUpxYuM5OVZsJ7cJlWPPKF06M6yggz9fs4/0Uf0Tp25f1Nu9nZk0Yt+uuTyc2bnF
cfnlQbA/sUtnqA2jvY6ocPqV0YGKjsKBjke6qyAWT+zxg0cZIM6YZhSjp7WfXruY
E4JMXIa/iWDJcGaGDfVjw7n0XhERfJ+FuAAcxxdSMR6mz+/09IQlFgoWKLEGKlse
XBNi//IV0Q+cPvntWvm5a6ReW3jOLXrYk8rYkYwjSUI2Z/jxp7jNtnb5ZwFu+isV
nPwI4RxUcSAQvaXwmbr6mKDozqnoxpgM+nfHl8c/uompzBEDJSPUNBuGAsbJIyCU
MrDdIElBjGJFOeblbRlTx/q59uPtU5SxwKFQRHaoakHKB25GIQt28xdgGbY4XtHt
7rsXyQ47yrp2oufmfBJG9wi6+BrZY94PCAFBsWYkiz/96T4RrSHEjzgpg54wzmeu
EVqJX0ffCwEBjgjGtrPelxDxMWn1qhm8iuSCSuNf23w5zMiJvX3D9GXbxRdCKzYR
QEa6hvF3PwgUInzJnw1IvAxxiomE9jDboVfvlQC409cC8TGkcMcmzdBYvYp5HMp2
Ld0D24gmf56Yh2A+ChmBs5GTEEO9GvXAhIMadGAtb1wBw1ptb/GBE63ul9Lm600q
VEvbZ6821jlGvLZp6NUdZuS91e9nsCLrFfQTuc/Kx2oO6qC/gm3We01CrNwTr03A
HyQ7qzbY1GnMu9Ux9M3NtWAHYpqv2QGgERLMPK40U4Q2nlstXlurgguUEsSwcSGq
xzFlr1PPc5W8ondSaHNl8hwNXXVm2S5OaYsw5argz7AlqDkEHTVY8ADuoYpIJ8WT
mqs1vq1YXA7GsMgtEP5h8Lzug/UQq47E+akIOH8YLttYQ5VAGSBsMQkIOeK/CH9q
RDq5RDI0lJYB8sjCXO7T7eW22TJzSnjsjsji5tCGZloVNDuep7Xo6V83C375KvB+
vEteocgH+wOdc2r+umEIgw==
`protect END_PROTECTED
