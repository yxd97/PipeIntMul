`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5PQmWhFtDeU96wZAUPYhbyi9JQzvnDYd4wkFPzLweYkanfyL37hG38fihB1h3r1+
avd219CCBIVG4lI/lgQItc7NZ2fFNXOAt2qaplprjbjCChuHQWV/3pwJQ8YD5j3e
jI4olkfTe6Oe635g+IBRRif/idQ6BZt7AHOiUOmEK9HG42wZvJMFYiYZq9bT6rv9
IomguGw5otH2176nfQX8TPll5TPZrGLNO80naH8CQoMLk2f5Uwz3AF4jwy9/0kRv
jfRmfY9EyZ5AUkg0bBymIlfsHsMy8tmppJJhHmVkJfzj7Ht6qC2TaxNziqfUYnMI
A3xAEPW0iD5sQX8vI77VEoilFnoJGsesZIhrnL3Ic8nuyxwEoI4Q0RPwFMqeLTRC
+jwD1iTddNnsr0jzBJO8QHl/E3LzJw4vd2YsJ7RdSDEfgqNUYGazJFyRSy6+Zk62
7VKjy7t/7LKv6DcqvPO5Zea9sjocQT70kiZAoyFVhC25q5Ggm87zULmH6cNNsLaI
wggChiEuWUv9Os4EU9E1yQ==
`protect END_PROTECTED
