`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvChiKWX6wAI7hb84aN1gkBvjFZG1U5V5YhuGzhUKVerlcam3cPhGQ+cN13i1GzU
UGBHd8OWOOUqEuQVRVtJauVj9ppT29wNJWaUTQeQbdFziPA1qoPOInpQyXdImfWU
LpZB6oZ6zJMdFU12M/5cyNCRsDqOfJkSVRX/DsGOae18Zhb8JyF+qMQPewPX6+Y6
8Z9R8RHAQLGxb/bI/mB9Yr24S8Tq5z1Myn4KHTe6QnLIOJG2sCs1IIZdKLlFbpvV
1Y560whWZusjJO5xerE/08yqKLuXkR9T6VdktOXqBLWBHmr7F6ccFTjK+C2lwZ8h
ORmPyDDp96/fF1mUKnYo/liW7PXmv3IZB/2IINHSBXOw5eOAVUr+nl9O88Acgnpk
1nH9BF9tg4QKIG7TZt3qby/07JpqM1SO29LXqS+IOFA=
`protect END_PROTECTED
