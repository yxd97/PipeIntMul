`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19Asz+2WEFGG0ijX/7rRFSx6NrSQTozXvpZuf0Mn0u7SYbRYKhkdIFwee7KFza1R
Oe+WA1oZ7gRjvsb8H6LEC51Ah4z2RZqIJLA7AFgND2hor4QTuOj4/rjpk6bampgx
1jQITWikxxSEbu7tp+vmHcC7er7K7YyhqqEg7ktX9I+dTE0tIkRFCcuCsfYcc61m
5Rlq3TVpBzxeg4w7gT8EE3lUehifU7XNBrKtyAcQVYYJLmueNzSVlD8rTonAGQY0
NAuHh6+SXMXQ25IV0MJvhCOE6mpLKJoDgQTgM3DEZ4VWG8cLcSy8MMqp1TYl4/TS
B2azBR6P8gwpnSM4EegM4TuhPzc8QTIs3Y5nD7EWkYkmbrhTyTc0qBmKWv/S19sV
22ug+xk5EZOxzyBdJL7nbQUD3s29CShfCJyN3kodQ0ByrnhtN12BkGnyvD4dX7Sl
oRxrsZycQ16bzyfvohGRgkoAHDxlilNGU/lBO1QD6Z9wZzfS7rhZmqBQU+iOtV+Y
Itkk49wD7mo+xSp5fBTuAsYEd2wY2XuNJ6Ouf43PkklIY36pEeGGtBiEHyiH2ykG
7GkVCyWgfh6ZInzKnU3xfOJQoeEmuwlE0nejD2hpflMYyNsLvWguNma18u71K2xv
WIxlkCgzMj3KJvxbTvo5uQYDjYMfi/gpPxdk9LRpUyuCaX+u2MS1xVNxKiEbzCyv
P+woEh6mUQ+68sx3p/rev4XVS248mDXks1x9CsEIUBOyJ8h9sz2jH9ASbsuaNi0D
YxXc2Crttzibg2pZpg+CotQMc7k6+RcOHQwj0lyWwU9o6ZiCaHJWjcqUjVQ5kCVk
aksq1kHMRtVCTuSJI51cGKwERTl7As8qnt/1TxUirkEQbMOVQk460di1YyjUvc1v
1AkewSCkUX8q7QRC+o2wLsKVwfruwKYwdndW1pA6jKfqwqDtrQCF7xt0slttCDk7
xnCwAa2z2DIrWuDFEz/65bPU3g4NWDd7BstKniwdVEKwy/MK2yeuzYBl5RlbU1JW
SbDlKb3NGbsvYkkrfhzkEhsbfFvuRKwJmHSXCKUstT6IBoz2HXjkNmgmfkHrG9Hq
gmvnaPOuE8EioeszBGAi7AkMvB3F4WazX4XolpPJV3A=
`protect END_PROTECTED
