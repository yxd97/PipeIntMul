`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrOnNk8kA2aV0WMFWaQbApIeqTEdHbg3h85nJAKgXktM6Z01mrKhJDZmSlO9Gwja
lkEqyhKmJBg4ber2/YypjUFdSelnkpngMj1oq/+wlJHLaX/mdOakY4U5pzTihP65
kcP7/5rUrmNqjL20Vs7s8p2zYW0y8xw/VT1JF5B7suqlPqC1WeNfnSS5oOI0Yy4H
YIE87EzU6T6doOv9Z2bvY3KUjyA1vG9Zef+5VdwqXr7PJLW/Vn5Iq+jdeAAMHCME
gSgBKJ6n5k72sw2XyuPAQeiWs1/obhtKHu4wC+HlwNdhGE0M6Bn97ggVa1Ee5vZv
YdItm7tz0nWz1F12sahl69lols8DC+K16janRS01Pbu7pxuvng1R7xfDRJi5oz5I
CTpgmGoWyEjcwqAmt42O91mSy5ogAlT9PH0vQP/aG1OSFy7PJ4yuoiDqcIyUaLQx
/R3A5007c2DKmezHziEZTxEtoYsrsDNVS3yrdJe1I48qSpztWbMa0VtIcTlmouut
ET7JEcgjsTIVaZx5uCaDKHoF4Y3dbJ/PQX4/BrrLEGlyYR3TX0pHUxIvzT2E8COf
v1ZjGqctv3atu5YrRoIZWZZu6CWrWKjCjnkgArARu4cXqoIT746VUlmh0e0kjYxu
Ufr6zsNVQ8w+97ly3Se0d9m0RuoZy645UpNUvsxuCnJEYAUmtZEIvcnivWlaFoka
rOTsjIuhRilhUwbVh2I5la5/jwptnVJOiWXu7+zBqdX9ypKpZdbaTSFmg3TQL73k
tWZb2mBERkxVWpjEdx9DCknve9jY0heig63rdVScp1nHtwp5NlJRraeKxrXWLjtO
3okxDHsWEgashQPdD1kDzsQm5qXLVxv0p8Bfd0VQ6Z3Qqsm67J51AzIddiYePKWt
5W9KVl02fL4TMpKr49fuINbViR6GT8T9p0Eed5sF7N+3hNdT3GUtHHck/lj1xNF4
HiVlpOo2Ml5fDGsC8WmP5X0Yjx8KHyChz/HSwfH941KMxFUNAYiyhDa6+j9JCNpA
/ce1Z5z1s8VPdvCEi/NoxzMhugnELpXqHNMrwy76Iqw0rZb22lz4UrF/8yuz/LcM
QUrPB9O5yxIMGq+Dnx8Ti+N78IOFN2IOmxJELf8PbMsD8+cko5F4T6xN3jl03JH4
CjgtUxA0pPPefcARoNdBAmKBqe69sVi6Hqvbj7b4R8gVVZAvwLZWcCynz0rg5OIe
wbbrmfVZKlSFgqcg14jUfqTDNrGk+kb0cizVjRggkJfQXUzfWh7Xh6MgPKEfIr5m
yWZdVIa8xjUWH90lBvVODxj4qW0mE9VJq5OwpEKmgaaNm6tZ4WAI4qH8seCABkw1
7aBc1BIYP8DEoH59b0xpRTACfBgeztZB5roUhB0xGmxXBJrqProA41m9shpxGeCa
vb7O04+LzOXx5IErw8bQxoAYzv2hKvBpW6SZ37SvmgcnzjZS7I1xm/Lk53qsqurK
jxoNq3xOnYTr7aiLSSyLoUfdx2z3VI8pAy/ht53san9WkohpDOyk+L0Iwcb42YiN
plEiABvK6ydtN8wij6rE9Urqa2jCOCGeykzBkoPaQFWdu/fSi8voVenSRFQcoZUY
lxN8ytfMQy24X2U+XLie77ZsWQLGaHO6OPpJmGKOvQVaewP1Ny2txmKGPaf9Ykwt
/2vD4mPhoQZfoiuBe/85tVV8jTvKOpGPn7mdozCqiCSAN5BzF40xxlf/tRGGo0Rr
sL5nod90UJQI/kA9Tfu5eLPcRCJRGht8CnwFvU1o4CVGDLoE54pyYnSw6KBL51GA
US5cy5c+BFyBQoY6P5DS21B+MTNbvSdv9eOTxlp6/8WHLHeO51pAGM5+Y3jU5m6l
t0qJ7vUmdlnydpg+Zs2vM0nWm+1k6ykKWk2Zr5Qa3PKxO7ohJpX9Eb/e1rm1rOcY
2AxhaUKwXt6HcSRdJYuK9bVWbtExLoICGhz7NCadcfilDzql7QTurkN2luYKWfV7
7im0RS5cPT1p69fD08C7nJgYOUvfjsTv4m7PQsx7ijEI9J1wLmfsLOnr6PO9sHw0
s+Pg/3oxOreg0NKJ2G/C0x20r13MkAzkTwEGGIwiXQ/EcGNm/EyAw0fzE0yL72gz
rKkCC/L9js8lP5gqx01q8E6CXQsLquiQGMtQeOIFhALftjtM0nub3p+F3hOnSCGb
V+PnaVlTR7p8/Pb5Pl8O92dg6sZ/0l8ee1QkY01W6AFCC+xVGwdXLyayHUiZwsln
LCCtTziRrca3C6Zk3x/dQPgptzEfqaP6YHlYt8KnfFrCe10itGG3gon50Mox8i0+
/2mtDmPBqwJ6yTNh5MisUF9APG0cj7X+pSh4iw2ESTcRtqm+RjAn9jNFMyGNsPil
nGOKzvHN54EtUuG/h7ce81ZfpBYUCAlZvQduokXTpKp2YVXDPMcjIgOfs6+Jnb71
2gp4ecJ7yYa1rJBuvoXPcfwFMsxf/9DnWtNvIG7rwXdK1hMwu2fFiBKFVKhaAMsw
+Wy7xnBb8DLhpl0KvkoRdcx1w5i2FfYtw0+eYVCYJMHzVD7nuESo0LNbWbSmbMaF
1vii2gXPGYLo7kQet6C11OrwJ6dek4Mu68mKJcqh2gYceIvKAzY2YhzlIYI8ANSA
2k2T2m/YFf0NTZTvsRX37l0ttgorG45HgGc2YC0octcz3O7soPHs0gOx72BhY7Wk
AiHaSuG6LbOVoZCkYizzCfpVWU01/76q5cbLCpkU0RKPttWCxojV9fdDOxj0v/Xs
gX87iDGxVu/tepgxSYxwkOv89Ii9VeYq4DI7K48zvmzWGGiyxhdCEjpUozv5NgFf
tXxVUXRplnZOOVnMGMrPOHjVAfnNM0h+eKCIDjL3GYtii7Z+oG9JakmRgmnP4H62
N/5rhm7YrwSUei4vTi3ftNBklA+v3LnspnnuJqf76pTUTohjEMqdpxWHS8YyncML
zTi7iY9WE2n84Ky/o/y4L0H7wSVh4DK1KKMYTKTNQfrgGWuO1SgXtOUnJJrLMCtk
bPeFarmgCDIgE3i3Ty2xSGTxdjCJw7FNe6URVzCvxvdbXuZGgjE63tsUJ+iqBW3g
Cz3c6llXZ7e8+GN+Sqks7mzHeKMVPEzpWHw+KuwVRpxSKtd1RZU6ycI1TZilXem+
kFURFbd90sHKZFf23W2QBNZhRQnIjfb7b2+5vaFijD0+9FFMfJsQTqCoViWRhUew
uqvcSeJ9i68sjgRmvD06r3Ec7XXfP8EgrRLzvuF27MVClIUF+/H4oq6XvVE6twoW
dB49zF8ipcpFnXE3VyOMNFYRFQcdGEXaOFc+otgyFMN47BBewdpfqUNN7X6lWWdG
A0Mrg5hzblhJmPR6RzpDrth7X6Gl90DlLq9rxiLBUeG86VNEuVsqKf01C0y9zx6y
OEirsVrJO77Jw0tDuLXMvm8ULFmNMMuzjgyhd9AgBLyJ/mKW/AVQ5oyN/eeYfQoI
7119uyK72r650H1uwxlT5QbC7dEloH8CbzkoeY5rJrlfrhtXIuk3UqjJye9ngFje
mp+LXECFPFSPFBj6pxAp0mjGVKqzj6EDyr+YxrK4EuhLc0N9pJQb3iSBSKY5dz5n
vjK8Ih2cNQ7bFNEHpRxjFC4gXA6vABFdLQQErl7YViuBpq11VlgSEgJbGYU4/civ
un+o/uVQfQcXrER59qpmiVWp6XI5FKtAAxtwfyOaQ2yKYqhr8XJMTkj6FdgaktbG
1NYDNyFSDiB6wvCe/CsfHdThitJ+eKBR7F55hhhmY2YTo3S8RcXZeeVTSEowHwsl
rHURKkqpv+viYfY09OLKsRIIrQQNuju5YOlNFQWfIGVGo1fa1Gkja43ID7cT4F3D
aCvoOsSJHrUG+HR39VvjUlsOOC1q+3d9x5uFshKcNvd3hm4zRyDapjX/JpdSoYRT
nXkV4qcbnuIDOg0vabo5769qBZKB/x3JzYDVs+QoXxicKB751wc4e1tKQJyCAwJz
OvL9tNTVmq0B9XPe6LAMLk7fCSa5ZgSdXgfovZaCK/kjP25kQgIwvyvoQwdje1Em
IjP+TIfk2kJHFrFt48h/YhjoN45kuNxmTiDa+DwPuuLkuwO/3V5sMQULu5m/IcrO
XzxsZ83fL4SDzaY1KuLZwSieKKLVsP0/PMReZ40tZM+zOX+CQBJD4OJMo7DLTHz8
RI4GmbhuokyYaellwnlemDCiUiYr3OMflD6SrpMRoU2ORKdkW+ExLlGV5zsm/lAO
MFiDOHJZ7aDVJXzZ3/L168oAHtVrnTlwyxhlz7pMAzjZ2ecj8lzc1lTB42VCvcsV
3FbzbDq6uw2aSxHpaLMdoUMgIqfa2emBHRDeHRiL4xKVDowvqG53lz8KPxYeidFw
dBleMK+y/vk+PXnm9xsFRySAFzAxx2WIU58t64p2AwAAS8OQkIl0HeGbB6ip3YhF
lWh1/syfRdWwh28FXY1SmqZp1VXHRI3IZm11SljWoAk/Xw3k7eZntAuLuTMHV7CY
2hED1w0TpQzIDakEWWNq4Ia4FYGRwSw+/8YsFQhHEWw6r2IRTbMMm6DMIt8UTx70
vKQ52GNLJp9o1Zrodcg6yM2Fs19idLEROsEgBlqpRTAePPj30zwYoNENgpug3aJg
tkHFQkGVTO4TSLx32PvUU24bbrZzYwv0h+xH01F4h4I0VEXIJENK8hPaacDJkAvZ
VXjNWNPbb4HrQyo661FqPukWPMPLxf6praYDtVw9c1ybx8mtkyP6deE9T0KvTnWq
+0cuDP9o9dMMoecU8RkcWC9pyLYon4EtExg6trlbix1+G3q33p8MwUcshzeR+2D2
sH3h2Ms4xzQV1uxxx2ijcc8nciN9i4A/+261kxfIn3rQyZXkuaLd4ADYTcGyfBSJ
SSsUfuCPv6vIS8/JyPxhuXWqPVGTssreLX/IzsHB1RbzCjB0T6q+tuOsfH+kOYeC
/z0sRxxHZjGY3ZQ+QEZZAHKBgW1jAjmrcgCa513mPLkvbekgL/ExYy0LvE//MgOh
pV8PlY5pB59+49Nj0MnR9ZDGJIL4nNqIDpkmBY6nnbPk3eNv8wyChQcYz9pNUVDa
EJ1g39oPtg1JGMMYuYXnrlIuSWBqTIC1hR2SnW8Jm2iiOVK8/iboo9egaB65iQkS
F95+KPKSWJmI+5eRwisIgANOzFsSFpfNtzymUhb4YW7vVghL0BwgG5f0swDJ3qYR
Kd84/LHKRT/FkeCwbzNF9nVGGgCvP9ZV3/1TCk+Z6r3zwtwRWxGJgjA8SHFAAZrQ
iBfinfhlv7iOkWjSEyDkO7JrLUDt46/UFGaDEJvafQnjpTn9S7bZFI3EcyE5FYj5
PnUra+TgJwQpDkKzsn5++MXfq1QNKN+LGOUCzarIscYzKm10WsCtQf9J86cUyp7k
0yrJdWGTWiX4M+l5wJheOo9hYLY3mJNJPwooGTDC0KFaqapuQmy648D5hJY/qC51
t4N/MVeDDovTivttcGaeXi9cGSgVvVYEVVgHgmx6L8MrdsrZEO4G7sTdP3EO0Xnw
S0+WYrli/Nj6nPwdb5pFYn4p4JS+6iWsRDsZeyqH4OLm+OUAryCIrv9beb6CE8xq
txf5UVYrwqB4N+dUXMDNCK2hQ9H+8YtCKKEYSs+a4FKd2uymR0wMH0HYjhI3m8uD
nyI2YKCYWZtpLtb3bbRZiOeq8pHy3vezkeBt7oLYNtmvvkjDwptzIwwF8XKQwVmq
qd1yTXiERbfWKoF68uLlPgSsRZs4slqisCswX4voKRnNNs3JziWzlK76EzcHbtYm
DFrB9PFA0vPRcTxhqxLcesVfJEufpaYfc/HNPpJA/RYdLdmx+uevEzQx9cJ6BraB
cR8Z+jcc+YJlPdRJZ05iiXdSxVgoy4bLLQS8oHbaXO/mAmeWYLPt+SKWaahorcdY
fnbRCXw9HVw8lSCzfdOd5xP2cIGfsuYPcIJ5k/ukeA7udR4glD/3ApC50vVK/Jhz
UOIp6okxXmaaEc0ZF9LsoZ0F3SoVc1rNV+UmLuLbQJ6TgC0Lw5kEzib4syp0LVb9
eEv5aLFERLfiCP8s80+A1DMXuA4GL0W1qHtNFjXsxuVELoM0o+ZwaF2aGOhUWIgd
HhKw8/Dznf/KJAsjzXEb8wFtVItss/RGecFnna0tnzYLAWnF8m0ZtxtxSOJja1OR
wCgm2eQ414kjtZEhaB0c2mXfxiWe1ffcjQkPN9ugV9Ejh3e7uuofmuMEKMKaP/xI
0Cx/mb6cxZj8JUp5d6PkzSOjaDCPaD1lgKcJTP803t3QwF6zxvoj3/WKBU/UDu2T
l0KABXQoEcsewJuhMTwr/FAOz+ES1kPBFdO0fOHjkFtuWXB0R19/lAqitW07kZV4
ZR5LN/j/GBvyAwX0GCphf227bKtk6fmn5qWN8bgVTEOxugwR2B7REoDb9sWLxUT8
g1pIv11q8PPPK5B8MW+yk5P9c3KcqMWV88jJipNssR56Nw9d8r2ye5LJMjHjc/9C
RTu3oIJhpM02/c48VakrztVV/LQVhQQ6q12zxyVCdoRIYszsw1cV7vo0xLqnJb4t
CtcKR9vyalmXjgVdCSJh6/1Sk1QvVzHfbs+OXIXB2nNiEn+ZXIyR9KHHBOWnRZQt
c5ZvhxFUC+vMJXZ9ERRU8fVVrbM9RoZG/gyugrBLgMQm8DIweH5uXaIXIHTo3de8
NctzgBwWNn+mZC6iumJ7ISKGFefJ8Hzs4NO9DaOHAEAnJtOpTi3GsYGxWKtdbAKc
foxgfFj5IjRlAEpar/KMc73tVRPWWLSe0H/pOFU5zzq0mc2XGY8yZ/yRs9WQ3VoP
HfMf6FMeKGh5jif8E1n60KUdHfsfq9X27Xi9zEz1jciQVF8IxRdwwiMGoERcb/ed
Bh8wf/iEUvYtPjpHC89O4bTCR34cPOpR5g3E2JaWaDZm2PS6IB75E0wNTJ8dr9Xs
7EXspWROP/A/Lu1LdlSfk1aLDaSHRq0+TA/e6DOZgspzojmZHaB+wYVD9Rmpcb4v
Oz0yPej6I7XN4f2Km3Ikw/4KqI4KlA3MI2YuLN0sNTctic4iVpMx75aC2HlYLjBE
yWvXZkEbTbT9LAJSfOy3BspB1Shh/an84GDKHAIdpG6ysXnI6o6l3B4wj9CyV1Dr
hnYF/22+QyE+x/sByZmb1tpDVg6VWKbEjXf8IEGvLIrufXxkay+CJaM7wBJ0qd+l
tQVGfOk6XGGkPLuADsv+2UQjD5CsO/4aB00c+b7xMADlZgJoplYwyp9qf+NIQ+32
+oitI0YALkqzusUIib0qrXpnz3aTRwzV1TczeOkuifIR7xocyK8dOSmXmNb+A34t
XWCpA4bctcW8tRoWNw7Jc2Ar1XfS6fpgebGLqAmdNyRmrGd1sWXHET/AmH1WQHZa
pd3QL+zZW1NGcDqZgRAEizJNWSnJ/9BHeIntheM91LiJkbQgEPUe6AN+wH6TuwcH
fhsuedC2bnnuvpaRdKc9xi0vIimaVbPH8a77ekSG5sTN/1MAH3/LLeNp16ij3r6s
XyKWatDRGagowMIx3ntVKuDOvEMO+TFXIlj4k7S8saFvi+H99IXjh3iN+eJvJrNn
4GuIHWuZDEIJ4mh0fH65Ouq7PETO+q3GHOmUXFuysYYP4fiOU98y507xyGfeyJy8
z2+cGQFSmcYa6sLSJ7elw0ndT1Ixn+jZThd+5caUpO7ShEVk/4oTaRu5LTqgD5w8
CbraGYzICS3vLh2t5exO7rWCTpjqimG2/oKgU9aNu1/pey9E1r9xZvuPMuRmW4jH
5eX+CUHmulXgt7ft6AbTLZ8DoKHQPAsJDREB/cG8pJFwRZOZtTT/NnRlRNiJyU9B
AnhV1lxBRM7mUPq/w3e/WYDeKHGWeFqFNW1nok2keClKa3E9cw1lliIm2JHZXDlO
r/9ZFcR72yDOSbOr9DDXoy1w1zoASNPzuJ+dkIh8+VK7inu0PxslUH75fjAQABd+
B4KjGApU4VGlE54n84eOynlifHL1cOkpSVifr6UBwLw2fi1nGSZFVMMYN5u5VL/F
V/t1ox7WJYY6k0aoECl+A7b8NQxQkhX1OxRW9Dilc+qU6cIyuUOyMt0R7CotrklC
fSKXTzzRE3KYRNqAHWK5Z5EYvxTgwoaEglOdwZk4HIv15NQkwKaLxDiqoCegC17I
OjRwBdy502hPLi6w6wG0kxaUhQydLiZHf29UJgoY5wivLNsFPbfYkDaSSZb85Kj8
qXmMI/m2vsnLKV7gcBG17mTuuI59J4GCNb9Rh4bq8L09RM2u1vNCxolUXjq4Epla
fyKAaHCfkbK6SHy7Px6M9/Isj2EMukbdevmjCS57mUQlRGmKOoZ0D+CSNNea5Uki
iUXyJLPdFOC03+caMMPj7AmYxoJOQBs21umTUEPZEToKuSXHB9Rajoc3ar4UqMs9
qnOWkH5t9xG+cn7nZybQntBLjgAY2wGNK1loT+3Iax17EeQ+bLJ5iea7kkQY/iA8
zNexULIiaRjhAeX5/V5119ePGlG47AIEUAMSgIRAhpTIcXN1raflILkDNTL8hyaA
QoVxkOEbICPf0B60bS0JdoQ7zEquQ97eykTThlZBliL7ig7uygLUF9vYmO6Iy9cZ
weF7FCRLu6smTyFpcS8jg44zVQ/096Wv3+r+Gn2AE1rfwopvztz5uZKxiAhnaVnc
uT4TQz+Vjbxb6anYAOq2TOkfOfnFFTHRCV1xfYZ7fnJ7HwMHHpmZVK/OpK62mNZu
Phib9auR4Jp8SOK+rXIx85yq2p2AqyD53X0ya0qVYX9hTsdkn7aWFvDkW2K2wQMo
VwvKtBCWMjbwlURYcmtS5EeaOB9o9d7xcO+IiZsxEa6jOAx0dbRGeIptdMr/gzb5
+ATIYaWHr0iSGYKtG5Ta+RTdQ4MTcIT3Zxg0NDZsi2XRL5RhlkWIecxZQbXR1gMV
GO6QmgXtmJNVZVO+o01rqYkJqKhmtmBFGLWxel5+9umFUcWa1wGfqwEw99ayibXK
PF0ZGbTgysWJ5TQbFEBHLuhmwikODEngVqvKelNvUM21q8AX4UDHFHNUZUk3GcW9
krxBxjdZYrxg2oBKxBGP49i35jr8u70YsUUJaMwSbMiL7tQ+lnVF0SmGSV/mA4CT
Ah33XyAOKTkY8u1P5ieJY+fAe2OIKUsLJ6+WrxbgXLWYHYAD2HzrlsOj6jujqVDF
4W2gpeZl8V1ijTpNdhDn1PSdMqlywAkmkF17y15vtgsA0pQN0O45qXfMuTcbC4uE
sDwzoAI9K3mFp4PGk22+Woy4f0X9gniYbOqYourhDuYZ7Ao0Gr1W03A4dGcwIX/U
7MyVAfgoiXRMxh2vlm3kFsapGD3gB7NE+fqlBpIcauZSyyTraUFCoQtJm44bivmd
8Wth1/SfFEXaFS07KaZu1g4lBGC800YQKCzJ9tkXJJOu5Dr6n9IygCRCkaEKyXZ2
OyJdOiBBkreQ1610HpXXRaGhUiGp0RPXjhfakoYLrwZaA+ebyX7fb/HauHgWlnN0
kl7Fmcqm9cq8GvfOJ+Q10+w7nrubjUHKXYWC0sIb8hhtkzwejQQX3ZROzAVs8437
jSMRb/G8l18AGCaYcmOCGZeI3gXLJ7MCh3WP3k4kPV8jxshU9D7Nv24qDsl1bz+X
/+QxJPy9WCQNtvES/DYb+FULD9Yb3Vi2HK3wXdF7QaOg/SKVq6D7lfK5KXOMjIeB
kbFXrBZYQMwCeJdu54uZQIzyNVE7++WF3fVc1HY4iADcGVF3THLpQEEY4meUWwTX
xGV5LxjZTBP9uuVBybSqrUJ37/uk+g7ZF/MMpxmO9us4BXBf4wgRpyeJ2rfdseqg
63Gfcwr6DQdpPaSJkUyoo6QFvEoNPTxSjZZNFzmbIpP676WfnItAPQRmINC80CwN
9DORWZKztErvKEWULnRHkOjVIve6gsgfTZJ/7v/ivHtWELLrlnPkgVG1K/Xdtex/
P467jy4C3k5a+nEu2Qonpf2voPb4JI2hj0Qx5q2y+oAMfXTwKOzofeyQEDFDyquv
LTyOliWV0GgaXIi+Y/7ala/Wo4paZnXTY6eiQp7q3QXB24B4mjC46Mu0B27N4O3S
arPzze4+Bnr9gn9oFJWTgMZal2CEyTt3jQtXTW9O+0qd+lkOZRF3UkVrjqFhWkzp
KbGbirDhp8spPsp/G99MwAfMefsr7iCDDTW6KQ/jv2VmB64FHB/H1wniKVAUqz2v
JVrxAQVPrCpPzDHKTnud/H/m2JpxllMLt4/XsQ9GLveOnhBr/1x8Iq8tmRMoivc5
T7zzk3UntCd/13NslWfWIzLkSVAlcoxR35omvYn9W0yWq5uKCLp7qC8cVwNNbxBv
gv+udoB3jKV1vVNMrlud1AK5o1NMR9SsQaoC/1Cw0KIGs01u6OzRReOp8lsvq7Iu
BnWpzeKKxPy5sAa1KX8wkSHA+9IAgpU1QLzmJSxqng5tC6HPsz3X1lTWr3uAxoSf
N8PaVK0rYWt/+GjOqNCBGJzR5dTVWWEHN1XAH2//HSFCRNuSiOE3c6W+gSbHGQvU
IYzArYpx70+zGTnR/L6LGkQ5eeH4KGRJySu0JvNRkTAhkNwZ3n7gnovZLnDXbbAb
KrQ+uOSkXVR/sXjAFRjL1GQl/Ae2kbbo9jsDwYr26DstYPm0lDdvg86QicTHabny
V4Oxe6zugrMIwUtgFO0p9NhpC30U2mN1r8si4Lqh36Z1KVs1FeYXPH//zI99yu1I
7SpiIbhNfaTvV4h2J7og92rB6jMlegn1JddrcJofYn5GtuUn2htXruPft+Gl4wcN
GD52Mr2NrYyy5W/SCdCt9CbHWhfdCwsWCx+V3E+hmEYpyMhEThUYa9EPDFJq3st/
hbnOefhdzWUPBXDnu7+uKp/ZekCA5PrS5z1UcQZ8y0TwaifPvKK6sbVjOrB5S5gb
Cdz855VrM/INf/6yjSJ6FjL85qc9hWSKr2j3hqXvtetVXqCOe+byovSCSevFKrqE
Pg2+JalV5fGtMOz/T6gnhM5TNByDTtmA7QDjKyccKpM12bSgbYsPSNQCJFSQaWRY
ZXcYZtVn/Yv9EpyPOOLZjIsNRLherdc5JbWkO5+KmGZAGvmbqrl2e2MPZp7Lf6Qg
ZnEUm9HI8TcvaThCLHQU67IS6V7L2m34Sy+z0F6hIQWhHX1M599tw9d1uxKXdVqY
T5snt/ITDz9oSf1TlRJfQsKJZyp4nQ23qDfA6Ewh2tcIVJF3ixjG7CiAm4/s20aQ
2iw2mQqkNFN9ni7vvar1ZJwxFPo9NlFLJL6RUghIJQfXZCgjW0zXN80Rbh7+EaDV
fzwXek7+7b6fnLmL8FUCXuuGskEHm8gTBHmkSJehquYbyiaMdHWrXwg81vPk+Zad
5F7i7XGH9jOrPNYyQj3HXDU7g2ngaHcvCiDp0ZpZZ4aBiR4SvV1wMa+y+fe5giXg
VniSQ9S6vKbm3mcXdw4pjlLCm2qVRFnhc5EVwnkkykb++kj91+YxKJ24BrRJle3U
koA/yKUSzgA3NYLcCyv0uMkhBG0hR+cIk3MtJ9kfCQ8+xy7XHGk9DmnX5ghkk9re
9H7gB2KxpHQRR0v1VEpLTmR0TLweEOeNdq5QpFigzQicxdaKe5lsC4vWRW3sjI4G
P60gHxmZbfHu0AtZc7jATyjeMcA/Y45PIYljmSF2kndLK/iwP45C+t4Zy+NVaj96
2yWhlWAVvmK2GAuCsIKSjRJLRFVrEBRhCHJGPTY/nijSLl5SjUrZY/qC4sMYXiKf
3dCKwLHpwS9uBZjKMK62QZiWZE+xFIiSyso2sgKO9lWnNuH0UE7rZUs4TqSFWpCb
BKVjMwQ9UITBAr4WSk/0IvOxS2kTPQTmi7YL9i7wHk4vCV3stmHqMfaoNjJ1JX9t
1CUsbvib6xXtqNBchUcN2vD6NAxR2oBfTRehIl1e0MoqNXE+qBnOR6J9ImCfhm4s
kiT9h/ftFl4XmiE8AH+Ua4fH7gVzmmphmaeY/z4s+Atru6aGbkNdEF6sWQcQTOt/
jc84IEPWT1bGEsU5c8qngPtGAMApBjci+2wajwBiDgIp4htBuYA3AdsZWVnNksTH
MD9F1DGlsdsLQLkRdU7p+xLPf5Bs/TUD4WxhPg68imHsbCiv0pNwIgdsz2qbXrfm
Dr9mwjCMqknw5TM8vPI4Z/eT0gt03PWq0ZzxhvXFEu5/1S/p5I98CWyXGJRSL0ug
IXh8CbcL+JFyvE5Sq9CFOEniVaTCi0WBJQzJto1DTU5G+aItn7PwCY7fSgR9WCol
9YLZ5fPgMiwrV9ttaGVOFwzgFzxh8yZHnlvfnVwN9td/Mq0/S9zOUAn7d7F2q76x
+HJ4mIqN9ON2STN5ZirfAdL5y295MoYPw+MbKlVuEz1wgmrFRRTB8PyboHeMB1d1
X3O1ixNst3t1ZVu/Gfdr+HJM4hujWMpqaLit1PjjlwV9vGOuZbACevUIXirkBuyi
QYKPGpAbOJrhaJJMoKtv2TyNUN4g1FWG7eoIwVD3wh3BqX4FACXEl3T4J5Et7KOR
BlsIpMxVnWuj5Mp66QRZ9vMExClGcFg4XvqgHQ+Vol4FFdj74oOef4Fh34sw4YPc
/wsez++PY3+5twQYGAGbFOlFNaZJz1gsPt2rfPuQQfJw6q6cqJoWKPZwzbM9ei14
LV+/PhtCWiAXky4RNeTdViSFtoMy7TRlr/6xC64lkTbWP17jWhwm0glqXGm9t8Cq
Y81OM/Msu2AUUWno0SNzy47cI66DxTD9HbrJoDg5u8Buz9u1iFvrpfHlf06NToXH
zUOUiur2Jw+/n6zFpfinBTJYUF2TGwVnteFtQKi+4byRn2T/ea2UBN+RY0K7BYfi
TlYUPUBBu9j0d3zZOQQTZsvYZjFHXPGs8COX3cle4VaOYUdOhkPgFAOS2pvAXWZt
l09+MC11GodBdbksugOIEA5ixL9TKSlPi5ino7K+VaivsBt43NlDAwli5+O0K1lS
G0lIIhP40+pn+Jm87oozRRfmzSt0SqSIYnGDkcvgfMqU0188doy4vJ23pXRMnTqH
bIcfedJCSRi4FCZ9JKMU7/JMEQkh4jG237WKE8QDbFDs0YkipmGfNLvG+YrWh7/2
mw2rH3x4mh7dX4CXZUhQfQzn2KAuuR+ngRRZeiZv/ZIjOEl1TrIFxAPCnLMtYZcL
Nns4PNFZpwKA53XWeME4QKZGGmU27iRwsUOoBAdyAIxhiGfd8Ig/56BAJ8nVm6uP
56f/+RT33NWhYDxUXa4vJ+MxgTrOXgVTH4mSKS8LewGAa1O3VQdRv6MDvHQ7POav
NGUTNCP6N0hj66wVqQSkHmy75qlmPswXcsW8y1ydaxUdZiFZ2I7yaGDHkIT31xJn
qxJvFefkUMw/jSP7wHKW2NzWdGzp80mSEBH687o/mXX+eajmCnjvIWP2PuEnB8Vq
YFZq0MQtJuaXIGCNv14VROkD2Zdp1Yn9EsHQYOqN6s3hlMdSYmmtlTFHk+f8uOMd
8hC3tLgOpCGDnLlikfqDYMy/5Jc3Cj5TtFDB0fD6i5tJarIIbJUiiqQFO1OWl6du
kqkA0LFipuxmyhYR5+i5ijgdVw1sYozCQIhTVCf4YmrOkPWw6oTfkrvCQZqNMgX6
roYyQe+2/Hqm8SNZg6SDMYIXnQajFoMU/Vjoyo3BXZEFPBciVxQlga6jw/bv49ID
aHqUNNup9lQifRvRupHdkVaGah3PYZ404tPOsswLR77Kj8shzv/aa2BBavFNbL93
BsZkEalzzbDYn0LlrZON9vfLkoR04Ws5rLhzmVGX54csSz5rCXG5btYRHbP44twN
BrZqS9EHAQSDSRUerU+RFYtBvyZVs+LCfzbcMu59wKOL2xm66iNPf3MmnPrcn75p
m7EWKyaU2Eta5vmVnpNH8+pi2lnDPF2bEUwXUJT0ohNqosLesLLvhZRCIlGcK6mv
VqhxLhe18C1YUqCQsec/3Pa+7RrjMfwXAn1RB4UlYVzMc0HWygLmjXTlqmXN7KSa
TejhFnF/WFLGo/YB8p4ypEQiikkJEZkP4Z/d7H+uKeU21uBWrUor6R9iTHMd7aUm
zh5YNblS6J/eDyd9WX/h+W2zvhe27ynMbEA+RG9Uq2rca6dwvmaR/oeKHTuRMqMD
D/obeVSYwxHrHqN/lo5exHrwdyqENZEnjXZkQspLm9B2UJOugEaRFx15PVbeu64o
pawZug9Qefit+ic1js7cW6v7h2c6TzcuhVSLszbcqVbY+3iEBMb81blgotCxIP8b
tqesj52swvnomG/k0Rtg79tShx6jqExWaVMqjz5wBjsg81BRyebyRdMwopD9jxhz
O2TUnEZsPseE6K+sE6Q55bK+YPAgD/fpa6s2uuinKEWJ8r/ePmoawPquaX/J/j+z
Lg4F/sH6BqSjAoTwK6mOglnnr/UjdyuXlZsNRrg2ymA9uTkPA2x19IoReuOQKkTr
vVudSGgUPE+dg2nWg99T7FYwcvANSTDaiW0ztSNDml8rau03qp6wBSvAMUvlj4rA
AbItkSO8hfiarYse1aayhx74dszCQQGCGoTcIvbKVUJCeQfXzayMWbDiKX+/h1aG
Ow2QdnMc10AjfbuG0hXHreD72e6xvj5yudGfoBUN4OG5gscAx6pV8wJPESpQ2GK5
6fIJyLqWvu9iWaaRxSa2uzq7FOdRGanJ8a+3ELlkN497FHHNgLZfD6XeAYcvlV8j
Ktbn2Um/qADGD6US5rucoQKgiMGPk4XY6c0nzb4DpnNS5mDOZSN2+3eZ/uphCWXJ
g4S7WhVKHvztJEOWcXH+JZ0DZpT/MmVHcvoWzQdrW541NBk48JYZzIUaJk8ThGOw
kDWH5waOwt9igvzOnoCupr0Q2QSGawozcy2uVBbgRKvAUXeMqu5OEwwfjGMz9NPA
edMM/DNjqqIHeEI/iBtNGJrsbc9BnXzqgbWWINxfJc9BGdqHVEkr8Pr6MNykdA0D
jjlQIwVzDI/qRcbUhFZiaQ57fFnr7+KWQwVl5XuEIDlWYfL+z1UXTlawkOQs+gSp
kUtJrB1sh98OFvqTfcav7ZeK2xsNAyQ9+zEynS1oMscWtD6wqmJowtTvFP/yfer0
ao8nHoohpSgA6QV9NYp1wY1rG5LnNaPHf1sS2N9rUz4jlbDyG4Xa6j40cUK5BQCu
edFbGr6vX3M2jX4PXusG0t0saLCuN8xZBWT3adehki0JUrxldsYnnVmGJAHXNevc
63PRccS17RRIcjMxfluLVZVgYTgde3RPcIWSQivncEVCzsxWHGD3rkj24kMbmbSB
FMUW7Wj51ujzTy6+OvXLjfl6B1fOXSFpnmEC1gSxn+ylt7LTJr680M3nOhvFJdJ/
9u2INyQn+cAXJRnM0SRAbL9Jk7nQZPjU4L9dncgISZld4mpVpGeANv3wRmgi4dOw
pIFsTEksdeXsKaJNIQjFxvrUUTLiMJoYJX+t5ufmfAG9Wyx3sNKB+TlWpB2bYYOg
Wj1oyd9SfPuQWFf3XfhJZWHGO56HxMjPBOBc1PfDFyGBeAxGQk52pIv+yXskFuV2
oKHegcmhpIHK5y/wW1KaLiSu0qe7QUHKJhBVGv40vPBqUfTrsPZuH4VY6Kr82Yuh
GxOdgJPJDWlhNILaGgkFJxN9saHAZO4HMrW2usA6+IPgcIZMyHayYPN1Rl0tfgB9
Xi27msuqMexcNsRwve8wzKM1JMXLIeMXNnpbzNDVita9+Ht3OBqp2Q2J1pGNS8cb
RavPatCQyE/M+e3chuMst9g/luWUIC8RJ9XMz/7W7bsH0tf8ectZmf5QiZNekd28
JsNyeRWWm+mtujwRot6EQVuDbSJgW1X1wFESDLwj/eLPiCdTp0F6feUhUQDKW5qd
c2lnldk2zIKz3Z886tOK94XFR3UWcO3EZTaNxphNuHmUQR2WokrsNvoHxeToEtn6
xUBSr6bBfObaFcmqft1zaQeutydo9Rbt00Zy8/ZleFX5BRfJo52u76gz3qmjAXyD
nuSAeK2CRyg8xhiV4AV06O37NYJkBPEKFBhQpg3RohrcW8kJpVVIwT9LvdTVokk2
diAO19GDBTiHR59l1QNjKSxBZJbFDQQE62YvLpqIO9ZFpyfXPUfpTX6nutf/Jzwm
SVg4FwwIDcIbYNFLv1+iFodtuP03FwRdCy9qL/u5RJeJwkNETjicOeuSbf1UjQn/
4Ff+zaogY7L20rL5kXar+8iM47pB4bCwPu6ARp3zbHsh0OTNSYIkAygUVVVXnz93
O44bT1Lr7nBLrR42qeeAk1Tpi901D1n+wZMw2D16JYWq3UGPTspeoVi96/hoBRdG
sMwQIqQtdm7fkxfOasT9lsAQhzoMGUAxYNYxJNiuO+ZLfSMOyeo/Iv2AoeqNrxM5
bLRDE0J7HAQWOMFr6kALHHL2KokjMLyVAhyNnusbvgNHIGaR8CwTG7Wzxr5FTa6Y
8llP0MFXlFaDFJ9g1cxCQzPJWEXInlpXEWKOjaunl4DxWR7PB4rZ40cEQnE1bfvQ
lsQ3ZkTAqEncfzv4LANY+NuH3j8OerHHHcBBBfPUJ9O2vbZAFnwhwlUugh4vxPNP
ZNARQELPQDy1AY8TPCLrUtk3kLwr4l/aSSVlyC5MAY0CAPjl6wpYqgoe4o3wH5ux
1EOms8T67Gjw4JnOsTEsKOK/Xlh9kivZjFeKPG6E8ASb90snEu9LUdPJYlYd5Lhn
Yt7Q40n4Zg7y1G0hnX7nfyfKHHn3ToMoCKe0bFQIwtXa3mlWciOqvk59Yl/20Xm/
DVfbzlhTgl+OnSvt/xOS9mIS0krxlWg3/ter1N2BDvcxbCE6eDy7iJSQCt4PHuh5
9JMxQowpNnfWdj9Vm86ZIGXK90wUtYR+0K+aZTLRMZE+wS64+GJXPnVzMLEyDI5J
0zbcUg6NZVCRh79oDBK70IeADAtnEYf+ElpzHmb9Z5yP7bnUAWr1/Q1WXYLS71Gg
xwGLGO2kGMFgGVcm2eP8ay5toVLCACN/Q4MpCouVFJrfVjRjQn3BKihxjMJF8naR
CDNew1MKprAJzlG1YDvxW93xTmF75qZkB3kOfwJAuovEzLoizYJ2Es8dzfTtZFSQ
Gt/V13PV2PrX9QiG2FldACBjcl2ZuAav1dEnSTdZb/ZMtKu27oOopSQ2wIXEhK3O
xJAO320Ujha2BjBrnXTPW15V/00h6M9BPv574lluKNICvJ6g1WceIGuYBlnTjGQJ
WfWBpRIMwzfs0OSxYAjhOHvz77AxQLxDrrnIz69hMd6DVLSxaw9hg/XiOPealwBo
LLVRiSAVEkSezGl7mECNLiQYSmgjl+G5CWpkH0+kTGfhS2l5UzlEL5Qr6tuYBvEm
Q54JHuDJs5xbaFtkZdJZyS6HOiQyKPnwPEirbaFnbhGK9mT8wdJkhaVYX2PlKmyr
u20DMJjERgA5d1Mkg2StMABEyGzK91CGUyWdE96UXmcmHOBaetHbDgqfBOm4P9QG
DMvnoZ3Knvz55XhHRhcKGza4eKKFbrFnjk6HYIbbcQa1q2netl/HBnWld2P9KfQ+
6PONmBH0+N8qs8bvIR6EgTY+70SMSd9SO7D2FalFGasiGAyXoK8CpgD6yE2S9ksX
RbwUaVKERU+s9O5sJeDJuPOH9vuLf6zABUTKk3FMuJa7/eMWm1BV0st/9TX4zQmT
0Enkw2uOysIdifjT4bRI0XH/wffilKoRPH3vCxbTcxNgok6dV1zgAaUpXC/JAY/Y
Vsqu4nsyq48hnoLaRmuadrr8azAqIYp8zY7wTk962nTY7Oe0Md6khCq65/ualy7S
KKze6GO8QV/+Bbi5xLEQEd6m1G6WoR4T4qydV0QG5v9K6wyB8x6V9UHJjFg+huYB
jfN647U3nA0hwL3NTWpqgOSICd2lmmOVYnIdJKIW9/3K1Yo330HYL8hq3RFYYPFc
L+YyLWS5ItROnKq+E9O4GGjRDKfmhB+p9Qls0ufP1dYBd9Fh3VElRUe6OBS4M4yk
rEmXbTRNw1MoI2GAVB8C9CtrzQn9NAg2MJRhz1CsE9m6H6bAGmRJV4sAhGVA2Voi
upojkCDjESbPrMzQFFBGSkZ2+4XI3RP7TjPqtbn2aQB1Byu36EGZ97umyqgRvwdq
v9aEpSoFWBk341sWEqGNlA5YiW+OhHEsZrrMNsas6OUrZXUNiPKqynpikQGXVE+6
I7ApSdMafbqwx+AyLcEr4Oh2T42k0PWgoTzyccyHpi0MX6QQpJv4H7EKL5DM908w
IsiHyJiPN3tMDFw2KnP+jeUJXoZ9C2ufaVeo2YBKRfIUQnbR4DknI3HUXNyku2Ny
QimvxRugVJueV/zVoeYwotTGrzyC3vYb6P4uTckubVxd5jNbkpH6mwrq20/n2hCf
1HUHZUIZFYBEznnG1W6jNNm7wsD0/DPhYsw49NbvFAEGzyvc6RLjm6GvvC4eXVLi
VPeB+8DNDVNj8toeqg+1ABhnE7fyCXkofZLgx29ugl4LKNXmitElTfVopDvlX3yY
WD8lpDyxdty81h2UjnlBlx9n/A+Ydhh4Z15PDYYZISNz7/i6iS65EVc49zsM+g/I
sAgj9ty5sbs5n/FZFjeCSrBU8d/5p4i0cD3UA9vlzzq7qGjJuZJAt9IbwQz1Tgsf
xWIR8J47JDYe7SEEyt2gn4QTibTkFDMwDec/5Sk45yNDhsBjImjwC3NXjgZcmOrn
rpG8enez4N+8/6gP4iPJzjunrKve5he/O37UbVMv6LI3PrGM1mAdzMDEg0ogZht3
btKh5u3APBPgzUB4Ec0MjISTUFS2nnikmKOkGAxdncjuBiSja/c/8RUYo7jV+IFO
iQ2wfTjn20Sh8TyLYiCj4l4/qa7H8WTnlWrFbErjSXCMe5hMyCCw9EDBeHmImFF/
tDYX2cO+v7m3hO9l197tsIGQ0pBrd+GVbmLAvYcRiDmQAZpemwh+aqlqO1Kax6QR
/HagP1JBqmDmO1cAYBDHAI8xxqHSq4XHUiBlMTt/GI2DsKpC4bAdq5a4E32dOhZB
aiDgyZ7hw6qiZ2P1MDur9J7+dbXaHxKIhC/h9a3CvYDRpFARCu1vPY6PgSdUIl4A
OmG4mM1wjLq1Fk/TYATGIwBNOJEBIncELLQiAFzxNXIbr7zzfyMUXiNIDPIqXvCv
v+chg5vmAVA5uV0IJj8hVEB6MD5XAvqZrDaTu4o12zRQ+2nt/Eqn/gTX7XjxU7TF
9H7wFIW3Ht6LVDuSo3iqoOpSWRpiAMCF5ePmzZOwsBkKhhOIsl6ts/ajpW3+haw0
wEVz2w/r7feVBIA2B0+HGfCxULRdVNZNBoLJiQherFacpl+UttTSq94Fm+xtQU37
JiU5EX9ApwDUOBRh2dTVyEOk8kFGKpWNFMjZ3X3+jk4Im/2Ea9L3cnf8SYB1wXyD
+TBDBsHgXzvszr7vuXLrQBKWrq60Mz9Rfq1R4NBLnLh/IiPLGjwvv/Ae1Y2eGzGk
P7IcJ2mWgNO52V+68NP1p8lWcF7MsCXz1dlh1Jgmm6232EK5Da8gMJH03sJBdbcm
C35T54xGJJiip8STnQsnEshK93kzas/JwoEwhB2DVaNMkl9MqxuIeBzuCPwsSIz1
y5ZvFwEA1zvcm4SUhCPNJeAq7tze3WofxwhMTz6dZXUGdQjiN9hJe10j83hPhqB8
9uANgNJBmnFX0vQhlUDZtDlTTd1UC1HGF07H2CqWnNazgpx3QGIsrOjEWWSKGGh0
B9KVnssZ56b1NsLrMNOJH/gJP8bkDZFtJltIOtFloCTfY3BeHpeYUmyA8PyPER3n
9Gr0Z2kMoqdExqgFOdlSmTSH6zBhu2kCNWK94DbD83I1s6F4fHxm0lqF0TJRyeBG
msMlMsnmY8FKLUTIzo+lyXGzNv48DdOoYNsmZfM+B8KDcUgrH2KqDClkMfuD2AgY
3IpEg/Oidw1/6oFe0B3mAqjBsFIzURP8eu1/MHUjCTJwX763mY3ymanqcJXBdFF5
m5V4Xls6iyvzQBtZPEGKm7lw8BzhtRKz5VHXpZZUaRKrvqv974W0SUUqy986G84W
3vXBOhwQySwbbLNePjJUztIAL2OOUg4CqrP2T5ACB6/z1VynxsN4IKg9Fy5sPC+4
s6jEOglbP4jWUmTSLEUJca5I/LR48vGGg0nlQ7E9NNedg3EWMtz1lFfl2K3skpYC
3+7KWIKMTKM75/oBdmJfIwd3676vD7aQ3H5sBveynBuKN/szMM600N99Hx3PLKTC
cBi3JccmOSqUESoB6KOArg4YAzijWJZv3LRZymEB2TPJgqFe0xyM+XCYIejTtK+r
BehCM4dqyDE8Co/R6MUSUmGt1x/JwREIS5LAK0BA+SOWEHYvMQojzjkXAafNKwhd
xgonnrp+kN77KjdKXKtnD999touQvxpESAaJNkFcDqTjS4lrbQORUt9J26M3CRpd
dUeWUHuDOnKp19d7xNxqP3Op/kgc9taq89z8D1Yo68ChoEY87KRmiKcmTgVToqVK
GotI/iz7JjPGp8RzMiVM5Ha2pRxb3jvLI8Anyw9omALwGVJGqthOrHnGJuBdAWxK
KqmYvGK545lVttEudSbHdS2l9TArrUCAS2Klg3JLsVDJm+1fhPTp6nauSlmbhtAb
HfqwBITzPIJttu/oinTBDQgKuBOhxZTBqkFZs5Pmy0y+WxSx3C6qI9PUawkrNynk
7SsFERqHVOyEi6XOK1oR0AY32tiexjdOEl1/t1pWoFbq4h6g6oB4BDP6dvVjINLQ
cJJegKRpPW6lcxhQWwrjLqdZRxLjfYH3iosBdPdUEJLq4rPXjxaftS2DYffS3hOk
6vfYw5HBamYVjioewFa+RRvJdOe2FXMvpPOVc13vqYK4TRZb5GyfRtcxkjFkwMUt
wLAymqhp+01r9Q5a98B1EJPD3ltcZzkTPAzuz3/eQZiKj7L7cjcPWY37rlWj8ETJ
DURAenxNnQ4RyEThEvzs9CjU+itzPD0x9HlUXlOv72IrcgWtc5NckWt2ItmkdawS
kxmX3cBIMp2yuIRI26Wb6f8psy2MPQck+2f09IEOiEgrAc9Ozs9tUi40f8OGhZ7H
GxRZZjaCPTIV9TxzhRmmtsDyZ+JmQbxnKaAKfW6BxOwtTQCTJyL0fzQsXSnG+ZLC
AysrGQ9ZIqiBeWHO0KFTTSl/ZWbEFKIEpdfJAZhe/FrOZA38RoVP6QCgr2gZJvtY
SdvboxiiRhNsDDT3+IWSxSVccxxnFQZHqV8Tp6TQPPZ11f2GtcZSm9LaSqQMeyyv
MzqUdJ/VUcl6IiJvAC/7Q2XNQW6Hs3jEBM3rdd0W4Oi9vrge+jils2GzywjUE/4o
oHEw8EVlHgR2cVgS6hoG4IDWxsISx7imSkroBAYUPILhesq+2fEaWmBBM56a7mAU
TFy6QMxeKDlsounbIGdyhRxbzcbpiEZnBzc/8UIawCn6d6nhNg+/XPqcBdV1ch+g
3267RrbehLWEnAkFvkclR9FiAWXM9EH8TlDXMM1tZqixAl3KNDLfnOQW1vhLlB5z
7H+YfrBF+zES9r+STmkch6Syx6xjPNCP4idPSTgEq68McM0n/1/mpzn5lpU0uf+q
lTUqRy2k2TrE1o4nFK5Mq/FpzpRB53fit+RLQNE8VU3iboxyDSMu+N5/tQ1uKUQV
JiP22HP7Mu6cHi2/7r+nqoLlE3SyARfsUFkVVV333D9/32j0DrcgFoDSLQsVPrYH
/QLj7VRoAD9uhel/kIiN1KZav390c/tpCG5D34PCjTQa5zN333xuLXgJMqwlNH9G
gySbQ+9LhHcqg1sFDU1iinJIm0mgYy9cMypeLdSocTHnHX1ghbJQVAATsv4tG5sX
YvnDHd8lhzKWZ6CQSI5+jhYGW37n1IUjLpH8+3zlaW5IyyiM3upcNNnrRgvpEEr6
WrSk8VkjGw4p25muWr3xt8m5n5g3iguOu0FxkQAyECdV3Z16B+4lnhICZLAnYZ0H
qMUxaSK4saguDnUavRW6/oydLmzH9OE0V5CE1GOdpVGHcu9bQcGRI3bXDQnnrpBp
ua4t93jjea9DGyj/FXU6nPBF1XD4Bqa7sqm1smoKqQ3gkUVBuNp8MDtZm7JR6Gnb
lKUN5TnP4t0dCJot/h5zZ0SEHc8SJS08CxJo3mGtqyvjvMdmQCXnv4jEDnXIe3sg
/tb5FUymvfpJdTQUsiDxEmsOFeCnHwfuobrSFDla9BV1xGXxrk3yD8eyVij9vqhj
Sj7dyfSZXINcVJmQDi0TVmOQVYj05COyTfnSpT0XRn6ZQzLoP0PjK2zC6tgMNoz6
mlOduY0Sw7LF66j1DSeeGCz+PtkNp7266CyId0WugwqnptHAqv1sH/UrL6vo+JAK
q1L/Rz1F4fgu++/BmZMwhPGo67IwVcESjcgIr3DkNSlvcfR+Hc1uDQPQtYMBPonw
PzXn1ObVvcrxap5bcheKRmTgapvgo8RJ52mdWOpkH+I0bGcZdj40iTBJTtbDxqtN
juhw1lvsd0TtnCEAevmXK0UqdaOCZ6jAZixU1x1MZ3ssVUnIpifGreVAWoniAiU1
CBH3OHvCB3jfy4mERMC8iFwlvqZGgyVyr96zLNMJJOkYFDM0ABNsLf5BFgltMybE
J9IcTrZyqoPlaPWI139v6y8vXhbCcg2/6fPZRTCe3oFM5pwYreOR9knZ4kaBbeCR
/a9+kK4lvaYmJS0oBj0IUoDYSPomC03POIzRRgVA9RdxuZwfn+lOFITDPJWM+e9u
zy9pmo0C1poqKn4rvbmNvxjBHvaKPTAnh8jhQ5lESbi6zz3VpXroZXyX0sDJbqzt
ZKfmVbSwJwyjSLrQl2vfbJ3vijYJ6uSOnd51umutYDNesBchg62Jhd9sUwAjGk8r
+Q/L6XUqji+H6vI2F2i4TQL/qMUmg9J4khR/9nUpcrIfKBclJfwfkgvK6DtNqaiC
IbDRXxHq4ZV/XwI2eNhq75/2eu9uOQlNWgtLz/7e3lgrMYVpqrGft8WAiv680Zmf
L92BLk4ebcEAILFYU6F8UpEtQmxboGC0m+Ia+i1fcVKYk7HoIN4MVBzisNJ194Xc
1ZRFzu5KCx/nOyO3e5tdBnKQIbtZBYUcdrYCz1EwerA9fpOUezAlRo55YjBSxag5
Ty4oTUq/q3QxYGgBBlYqg9ewGsJZh/EdRyvXAWf7fRilePzjB+kawNL4+k7DwxB+
Afk3UVb7AbUkiLi6otSbuNKlxOVeeZsl1GCGEx4OhdgwcNx1RPY8GYCZNqSbJR4z
ad5zOmIN3oGnUyGcCmUlslk7zpSCRih0A3ruhCn9cJYz+EYnhK81unM/qbn3VFWM
sXPmUgboslWbYRDpwctn8m+AismqsfTuS8s9hJrh4AjK1K3fpTFfKfpQXk1As+/F
Q/3Z71LAvRX8YaVdkAyuXfzsBDIy9l2pZ1aDEcygoZTALLk6OjxUpeUWZQ15l5K/
g0V0A8RycjfcSshQT0eFbzyCCg37MbiqeYvJ45ws2BndYsaMKAbFvdCMiUh3oa2T
90geUIR1nS8acXKKXnEPZruoxCaZAoYS5GUgby6FoAHO7Zw9yejLZbasw0WEa8UD
kQkHlGr7HBnPupWiMFnLf/8LyipFsmbkNOJ7kIBK3N8z45JX4HLOzHZOIN51hhie
KMdz42P3EzcjJVWoDmctdoOHLlYNNkN/m6ban+a11Agu+f9I4qBxIVS12wjoZLCF
26Fo1Ux7C08cfDUcmwmtiF3ChruBGX6zof4eLsF3VroL19BH1a+9SZpKr88p4rOx
Of7hsSLRAFBxVW3JliTeC4YzBDmLXzQGIwFhOWrPj4BKGMhMkdlPDAopJOaTpzav
57MzB6sWgVi2p4W6/NjZ3iyC3FX5WwsnYPEdeMEPHPyU+x0zw4Pf/HFISefNkwuI
0A+T6q00WSpv4fEDCv89X1AlzLDgLW2Dt7QruHXWaKViRZazagNfp5I4y0pE+Dfu
/vjceDVyYGV4HX/VxszVuPH5cdNCR26pwQ4ApOr7eUob+48/6Uzxx0VzoQMtZrMj
B56n2s1+NxXES3vQwrELdfFtuVCH61nJUTtCmKLx+A1I37b4u4K/RORV16Nt3MUh
ZJct7tx0yJNHBR73pdsT0lGeSVhZ37ZHfysq5ZigTHzBxKQ4XzzuI5nOQI0qeKOk
KgwmQ0ffjRbZ4c13FvhXr6K0Xco872324ikG7RMG+RKusS608WAD1y8flD3l0Z1M
m6C5MTsv/IUzkXIq5ERNQ5MODbyVCQ7/fzHtVFZZ5TY76bNp2f0ce0t1huuGyqS9
vy/4t7AWRlcd/TkP+9UrYJX1USg57CrwJxKj/83fli+fDrA81RfNZ2BcLhvMOquM
wqsMznJA3SUedV2PWTQWzGvYIe7uRB7DgP/cBwZe+1XoAkHI86diWAXaEfyTrJX0
pxYaghhZip7iFWcLl9h1LT9VA970NR3wtPrOFclabIBB3u6Dl533lvqUmAXbfdbz
PFbQKdKgH5lKCaeBs35WktYyki/MCJIZBz6NT678FuNkNzasYfV3OH0xM/AhgBVp
2E+Q65Sy6klFmGTPRAcgAcx4GTH8vY/ViCl0lVt5IR/En8wCSn5t7SvsNkbI+wEx
fPiUPZpritsoWb1Rg/kkEgQeZESeQl622tv+62wFBcGLFlwONpVmd8yJAjvKb+6O
zLJF1sc4BeXV6sKiX340XQhcstMTzjictjAyC9snRH87MzsE6kPwLo1T59JpCm8M
Pl4S/5GHIJYigBjGwDkfU4P5mkv+BgwwJfS7QYz7x4S3iVQwYS46iQqExIAF6LA1
3oRC4I7u7fTEYzcpkRWhfO/DKT5D7CWSpRy5I1MHY6am8/lhpKVJnTE73Tm+mfsf
iMJ786fOV6KwIAqMthPw8A78BamcZk9XIL110l6KJ/LvL/DZgRjY3zkn8WgkgCZW
yz13zOKpjutLdJX5aHoeKuqNgmf6Ar+V7v4xwfFWBFgAVNJ2eVq2evRvDC2fGgvS
9n2e6oTVm0il40PM5ECQH4LA1fmeRMzM2S5IYKuRge3s/1LDKe8xbuxeXKU0Hu/Y
9QxQSXxx69day2jb8w8DlgGSksjccOXsrmR1p6ysDfAzR+bF0a/bwmgu1gntr8IW
OKime6kugXRh+IbXS1ciqgZ3heIw2Ysofzo5q1IVLyM8Pyk47xJkGnI2roj/5uDo
g5TKFnzGct4GweWajg8VcRMpAUHDPnBqqVBRYnA9HaSIzGslGwi6O7NxcuaIwbgk
Bef3dtiTFfCnB2SQQPTgdnhObcQV5zRQpLsyzvfdUk1zn/6Lx7xcXEN+eQGgpG7B
pmPb02VrjbzOqVn67CRmI17y42uTRUSS0Ds85pfRSaMQ1mNO803u5nDMemwRh/TD
C4beaoX8dFuogutURv7MjnQPoDpVDFbQ96afO9pxET6yHgpNONuQA8fgn9GkTdd4
YR0eTsEdNRCOLc/hgl5yAzFRNWMTuW+f5cA+ATlNau/YAunrQMBxnQiL8ZAIjqWt
IpNUuHN0NRI6V4T6rJnVCEA+eroEp93YrwXjIYOFdwc8TNLT7uXHk8e4AMul/pLH
9QPfFja97LjTSTOiGh9zAfVQWNzpax6pXixOBcFJ9AynfvhTDJf36uFuiUAlPBjL
7ifuuzssbAJR0Zn7DGRzrAp3mJtm6N9mE1umGqyk5NR6qqyBmK5UFUvfAqWVUMPb
PrwO1qN2D2nRqQ8ewxQPJXxMgI45x7ihU0d1pl2Z5KRaUamOqrxlXxBLbIFBsaTG
S7ARIbmpT9i2ihq5D+33kx2yJmk3D/fRY5igCmvbYkFGUM2mVMW8izV2AYAcDmMs
7TZdChgppjKe5KBEu7DNOheat4+jt5NAJuAX0YdOzZc3m3NlJ0RUq6GoKUp++hkw
EfNhBA8M+/jdGd/eFk8s7EdJluPl4/sgQ5VcdC5GZNvD+2zeJpLHCkQzAoohRfpj
sJJGQFWs4AohTgtVWvOWgLboIC8Frn5fmqBL5JWKEhyKPI69AaXtjPPRiM18587n
MIKCMu1g4n8J6DbUczRRuLg02TIMtrNG1goLqPO6X/IJzaOAagORwBgDSmRdlrpq
5FhurSn2u3Mwq6wG29DlKDCxBvT4NSN7EBy0u0kpkrZh3g++1cl0KPNLqQLwIdGN
k9DLn20RE4ZoWRRR294vD7Csg9voA9canOqwe1mmYGWGNEdqY/gtjm6/MxSMsLop
qKbjK6z8SPlWpvle2SCl8bcmC94QN8sG9u4Y15CyLbwSW/xMTgLbxw4Aj07meyxT
8vfZnjWBbhEO2CGtajRw1XZfil0azmjHTJGAwNH2YBoOmy8zK8dLnrYXkTDxfeTW
BAwY9P3uc37dsUbVn5AFu6HspOKCzVkfG92aSZUp15ZKEMJfafsCjd3+Z7F8Aagi
1caH4G/6cZlgn/1gVh5gvTnvKsUzLgdXVu/AQisd6Y/MoCuC/aXmtwqcrNL3nGug
hJLh5ZeEWGmbU3Z9/0u0S/ZWwL1+SFG5d9o0irJAC+/ewr8IURa+p8tRqwgVDGUC
2Tsrpmc7vXdWg31goo87auGv2drdR3VtHYwTe6pMbvU0az04Vn/Ty6HH+gIYoGi4
QlcSTljeq8GKA5v77YaFXYSEn34neaOIIdzeH3v7DY38v7MvwUKgDyZaZ1apedyb
xINKpmDE0GugrcreGf88CGuwhqIfncn0gYvg3mMT93BbZxof/IWdWFEIM0NmCBkk
xAcSzpbVSeHNTKo6uZt2MIeqxkh+nAba2HHfRMVB6/3cxKxDPOCNQckkbNqxQSAC
4OzhkWAV22IDjlWxcJaz565pDDcAjvOIRiJ4u06UKsLd4BrhBGoJlVFG14t8pRKI
thz3HoswnERXnbAyDgV9ve99MTxKAqbhP8/c3Zxf2DJ1QXvH66m36Obb0rMWiYpZ
as5Cc6EBKCUk8krq3PPt4y7RhH2ru/Vmi4rag0xc5FFmm+9LvrmygW/zufbo/9zc
5pjkZsj8B7qVxhwJGqDomAz4tyflGBS8e+Eq3TRvgaljmVRX0NDk192K3vXKDfiB
64kQAvZA6dOBAgvOfzl+jl1VF2d6qLDH8dXgYuxlwkljMgFVnRtJCBTB0AWM4nGe
gy7qBNVhsOSIBwmSJUs3aQpgfVY2NzemPabIOploFtEC9BuERKYfPOfBQk9Nq8Hf
122TaEC38bvZa5eeAIWUOUMNzQ3viXCXxK2skSvGyRkaaP272Y0Y+MyRoLQKN4L0
WT8jo52RTuBR7fGlR1YXZE58fMk2VGiYVu2bJiE4QZ3g0cgxuFzqsGFtzT/VjL6V
SAjU+EsYlXlWtyE5AEkaxp7w4reSN3jLWD9OKTMvQkk1fYZy1ZsdxxbVu1AdTFPq
QgHeWZHPosTniy7oKqrJ7r0WrU48BJuHYTS2c9fENKgypKABxeR5Nd9IlEWHf1ep
aw7GeNNqGcOziE1tp8ynTSmYk1b40dpdU4ZDTi+jj08Jvkuu4xcVR2EANAns6k5I
WcB+m3PjdL60sJ5hq8kyWCxybkGGE0wFmpFJuX4xwZZrcedKgb0ijDIiHO5uawcl
cxaotOW7A4kPJcibnTvY16H51JrgWSjJmZMFfHXkDPmwW/ANL+xx/b8u15eV7apX
QDsbylvhTD0/8hM5DNZVy162vUsOYmSRY31Tw3LlFB3oYyDXGI1cL24fu4CspLQk
0SIcuPSEUT7zNTP9AZm6Q1eQGZxKdWNW8kjMP/pJhVnCBMU/LERR1B3eNyN+BeqO
p1Z7/J7ZlzrlfRbyb5RuWLAg4Uxq85zOY3aLaJhbCxND1nPBn15To50ODaJ5YRFw
QLE1InxVZoVxqUyaEu+8yN70Htj6JOF7ypwx7PeTwY7cKkC/BYn0JTT29lO2o1mc
QJmq3gkYjhMonLxL7qJ0N0QN6enwcCZlKJOiMCWsWAHrDxP5T7i8Wwnti7OkkoqA
CUNMAsxp79Av2GVxaWERJFOsNjwRBnhEIEpJWR0rOaElbh6TXXzrQNNllWXmmzbb
1UB1j1E7nJ+sH3NmsHdATtCkrkjKhnpMcbMUj/ZnVqvTBHu2zAwcFr3mREu0ya70
/cYpyED6b0mflDMNyXY43EQqZcGjeXXyWrDcoEW4OkwkrX3dR3N6odXwG+vs+/Hs
JLx6fKJD89Nq1eMcyb8PrIYgvkD9JGz/kKM1mUJmdLMEYnoJ8vYBWnOpnSBjyiqU
n718qCW7cDT8FzruNnpneiDk0PH3JYFnz6+68g7YfUhPkudvXEoMSaWPuH4e3UPg
G+hBXpgsH+CbpbQsz7AZ41g3lWH3kLEG5pPURNFoiLsn8BGPB6mbuXhBBc9mN35F
9tVbQqmf1zc5wlztTzcHdBxf+EwLHXK/hHX8AnIL3wNhyeuXetaRcITUOZDcaB3d
4stnhuVWu4yk2h+6pN+KeNVu8vC11v2roFKn0B4LmQPePyOdWLpQD0Gi9IquEc/K
91wNWqnqN0Utthu6FO1sPPlT+6E+Suz6q0S+3A+mvVKTPfdQoixHfJpbbM5rSBGu
5MCPN4g0SJrJNkAO37vd2K6yzQayI9mcgxnYsJNPTrOdywRDO+zLY6T1gxfvesrM
ukPNsMfVFK2fyI/q5m9WqjYxtTxqi4c8cD7NMic5v2c2xsxksx4mVDUWMAss2Oev
lj8kDglTri8aO5RSzxcgIsdZFNOom2F5+/ORN5b0CHUVf/tL68RSE9RCCou3Gw1i
4V8TcwDS+8JR51YUStrF3XpgctfeIuvGCBUE+B4sLIkk79Caz5ePZF1dX8ZN5eXD
TXEJoC7GwcO+do9O252VR5Nuce7yKOtPkFvasm4RScXKpmV6IJPvJ/Y54hGKwrQQ
ZGKlPeZenU2efgjx3OnGs3xOmrzphLR97RW2w6lblmdIObCf4vXpqsC++9zGPyEQ
lwP36AeUaDSzWrJ6ugCAU7fFvQhT1GOdvzy1/5xafjKYLnxx1S6b8LavTUKaXVv7
ojGczTrtKGUUQ63g4zSJBvtZg3I44JtfG841xdz5br06oHJm0sx+3PODej5s1gMD
S9tzuU41WhEPDF0/4NnRYbjJVrB7CKv/oJ6/hRkcRvlydC/nB5C/iJmJHaklYOiE
AJCVYZz8ZDgD2T0JL+VpkSICNfOCfQhj3deZc6sWetvib91CC3BIkcxb+QxcSvsN
R2TLOvG6LX/+g7AE7hLYtAyc9L3UgkTWfnB+o2pCyk1QlRyA9Z8EH6YWImgGjl0p
a9fWdzQD5eHwDwXRHQBNqD3T0mbrLADZV7/n9o/2iEvHHTsTT78DqdOHazQkSNsa
rEjOhT0zepoEQrJkfno/WcMAw8ZEf0yo1F/mp4yEX3CgkKwTYSrBjvU33FbRbYYb
YsJ+acEdWr+Pn91Q+Jbp3oFB5ltmjLiqmfjXavzUSTaF8co5udO/pBz+oP8Tj48k
gl/L/17GZXMPn6/mvoB3m4GqkFW8lDJnAcniYIGm+K2l7wh0ayaHtxBVVgTKOzKA
zPUpykSQ70UqjPnEpgP5RA==
`protect END_PROTECTED
