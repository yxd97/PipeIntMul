`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AsJkIDU2WxU554s8vrt0c14l+iJCl5NpfvMGflj04x/2w0kfz6/eCOjQFPGOTI50
OArXn3B8hCYuf1Mtl4d29aYhmz/JiNivq8NpvonDFjzYv49br22jBdRVmoWddwV1
LSaw1zDBVBfp/7ZKpCRCNZ41nF2wglatONoMd4YRdbyyU/OAl7u6K/k/KntuL6k3
GUkO7pKd3vDfvOKgA34jMwEtrgFlMLwaoCswgO51IgpuGS4gKm9X9zH2YG9IFW3z
7Ms3t08bgg18bkdIrWQGnac+44M5KC2XDUD21dYeYhwk+9Gq5sptRM0t9WllgLwV
MGxid98/69a8DyqXlD427B/+LxceOvCkXiculeqQKj726keA2ep+UbcCU8MFXkRv
h8fBJAePLzMlIz+Pl89q1t36eMTXDiZo4+UjZKaaJWtjPtXKhSDuFxUNcZTcV8YK
It5gRy/UYvgxyo1AdL0a+iOx07eM/9eA4U82q1Z/vHWaDNlwy18Llux6bHIGW+1M
6DrHDcs0ZMRvHBT8zGjvwSFK2Dhi8BYbnmTJ4pZqbMB1IbUgK9OuPh6NSawJdYTG
7GNQ2+aKtwP545M1Bndx4hWJdAZB5nJMFmapFBFWd3OPmmGxz1QLK+vHf5mH9bZ7
ekA+Bb5tqLWCHAVqBD2tUs95J11vj+I0X4bzIl3pyXMOYq4zbTChrc5GS0iIKYEm
u3ZcbnvmppqP5d6jE6xgZh1RzOT/5LlS1QAbiu61RZGl5E6VVxB6MsRnIcCNN0ne
FVLGmm1GJAKLY4QfDiZM6Xu3ZdK3vz6twzttk7AkSPEF3yVeTgJozgPm7erBMS5J
JU0liG5pYBcIN2Rx2uzN9YaoYDYov5ercZ2vKpOWyh6MS16ZPC6Lr05J/KkXs2eP
jb2m9gVM2VDVJhzurGTXpcvl2ojXUu45b5tGHl+bGz1uZtigF8d31OI5nSuBnULx
0621m0F/zYmp7JqB7qevzZTa0lmf1mrbLUU+OCVTP88oq7j+1LNjABtmjIIY+FPs
erwbf3LuTWegwuIXvFiRZjfS+iQQdbWY3c2yzkxsMM/3Wr6r45BpV3fxkoRDXVSE
7hhlhhedkzhbJhiFmnEK5xVFV2w8wpgSci+Rx7iP5IFofq88jcu8Fge8UEd1l2oB
ZElTJyXJ7+n7PKt2y8pus3Y+zwTC+2i3FwtMO0QLOtC+xjgT+bOxbWrkujiMTd0B
Urf4b6PAkOlt6iWZYc2YnFFRZtx/co9V7lXnEhPoRbOk3WDI4cQ3MzO6EAFpHeIv
LL8a/cKzwr6yPwP2hb94HTuFFvkDUTfk1ehdaRMHAfVEju5BQRFnGKZ9pWjl0tcM
2d5l3RfYeth26HRnd1Xl05IiKSGMThrdJ1a8tSxVOiOqwr2IP22UejjkG8D9e7QF
CuwJbxWEJW86XpGaPlRzLTTBH93fVorkOQABfGvk1KsuDSIv2PrBK29pu4U7JVFc
Nsl2cdC+aXA7NCY0J4Loi/45NF4CXUXxcdYaZwE94zrbNB3Z3eLQjYHTop6QL86V
e39BxVc4SbPoeM3nhUkbgTUkho1QQiBa2U3eHjT6tdvKwK9lny6lwh+NSequFba0
dll4tu4PP4zP5f5AeqN9jYn5cbipQnr6ZFIilFpXLp4k0fS7lHl90pSQnyCkvgAH
mBPFGLPZWy3Ie26tQ4LyV0mCXfTst10B/SlSgDIb8Mm6EUphaI2N6HPJYaIiKd87
g3SDqZv4tlfZ8HDnU3d9qYOMqtLfSmZaaldrM7cgGqzzczOc3s3Ldxqv1kx2tgHH
2cLWGyMQcODfOuMmz4cR8/0Hlijd8OKXaNzSUdNpiQPBszRofBrJrEEFkmeHPsin
H7YmZ2gT5hCfmVz0LwlMB3TcHtdpRLwLFh9n0KzS6MhhIIOnTZpsQHJ9+FocPIDF
hwtISFZN3tBjC7aatF4HwgGRABoq6jeT9ntRYSVvdOZUliYm+g6RtUaVIIsrez7u
t0iYyxScbKQxz7fzlHehNjkgYFmzhkXSFmoIRgZVM9H059pnYrmX/B1A3Jb+qoU2
o3j7eZmyKvt9aUJq1lxsIHc2IA94Ov+CEJXA7yiSSTFCmBFYdJ3U1Qe4Kjyefcxy
4x933LXXoKMY1T7XJTU2fj1bDzRA7lMLWiudfR40PvnJii/ECKQIXLRNHQ347l5D
co6VajRS/gLlLRpxwzDCTzkAtAZ+IZ8HXfBwLsZwy0TWdnj/+tDAhfIAQ9XD6NTP
HMSNVewySzovJ8cUGgMggft0/FGYuYrInvc6GvM83t76NpBCJSvb0sy1wqLOzkMI
W1+c9+cfrfwpMM3IqoDOlSDQfARHr10Gnl9O8DNjlphgFP51H7n9JZqjOtm/ySK+
ry+Pg0RrU2Aecp655Za4o4N1qyXTr47ggJhPKFQTJ8kG/86Az76BcEAjlmPbsgcA
qLaVR/k3yx0v8fOYsLuzHOdS1baUe5r3Qf3Zxdai/oIZJAwstrvPVtYg5ckr5C/3
/bFvnMI0vhkjXWWQdjP60dc9KLtNTGLIcDtZRi17QLI5EUo5gCn5ZbCr2OVv49Uk
DPWROZWEb60RjmEm2UjpMz2hildAaRuFeUiwG5XK6Dg5K4T1/HpiBUv/mc0DXno2
StjnlaMwnpdsnAqwuKGlBYkreWHvjubcszwlF2zNkH7xLhP3EHjCZwUvd4orHyrP
l7/kuMU5FScHMbCmJo4U4Hh7BfLGaAL9SuWBW0AM2unZyQ9xaD1MS498SRcKjFIK
3db8tB3ii4nYSU7pRfvcmx+GuCK96VqGbkgJqrzIwfGSwy8u/ObHNvB+Yvi00H34
P8SZ/XB6KThr5khDZxM79eBFMplOEyL/kcTjBW8s0mqVdTWL42XIkjEcLZnHPdY4
6uKGCjePry0GDAc61gZd6tkht7/gGryvDHHxFt7xHpsT9q/wat1BgA0pqawraZSM
yCDspZayBvFHhH1hXgF2fE2JrhUXrXkmk9tLZBCttJlgqut+LDwlhGTMDqOAwHnp
UcuHvWRQAJyJgr4qwHQYeWYnrkJCFKEyNC5KcYaKY/X0OUmPF3sp2PRt0hHXwHD0
paFwjyvxgiW0BdLVNbN7r5HFQ9jHkbYmiT/bcJLwbitE5q4m9vVMUnUhzsRjhJmN
90tnXCf0iYHF++zDwdWxMprAGGaG5w1JxZcLw37qaSLPg+r6iCGviWLkyeI7zlcx
SvcOu8mnEIbC3f5R/p0DlpkfL3Wx3i+xzVeVSW+60m2gJSuh9OVWJKAnrdss9QFG
cZ4FVQvBopW6nV9JfKmBb7D0s1bD1/01F0+z1ZQXTKKheKFaUm4DMLw9NAOuLWtH
QtmA9OuSXzk/HxaM4163/2WD2rw/1tX4zXCt3TofjYLpmU3YeabYFxd5qAaOBlZn
lBKAWVymSF94ZcAkKN1ckbQ9YibswFd2b43URepW1DygwTH0nKATF34X7sxSV8ge
DdcXeJfinjzhSRz/cFg7KFKMSu18GPU1hEor/uCved8=
`protect END_PROTECTED
