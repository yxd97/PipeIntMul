`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j3WKLi5z8MVR+W0KR08CR86hKkS8nWl3u1E+h5Obrs53zTb7LRlmFKawtlhFVURB
ZVbQllienXnxIfpQf/M5BE33HrR4fntVnFCRDkcOk47ivZL7wePQOmWVQ41+TquW
FmP/S6HvsSZ1EGtDNUspon3mhG+Bky4B5SsgQow7argEnNLCcuB3b+WoRzXA1Uvp
XtiQC7RiVT2dQvDSlhc+SQwV5ab3HalgcHY1DeBGh8I8qQfm0RVfKLGXesWo1T1q
ssEUCU0U28QynDk6F20VLWAhaYyEoww89yiiRYda5xhX+gvh4alexM3wSElGNNzw
evkUxat2uBjXS9gAA47TTUZBk5G25HZwIeGz8T/jHf4rRBlpBPrySqRFfaokovFP
rdnt4QiO9cC62nmk8z8nuWqbSLCrKn38e6mOngI/am7vtYf9f+9hj3n3bbq5izlO
dxWtlmquJCw3/T9hm+o9vzmP3kYwyKKkxiTWFjn2ZAlthJc8B1Nd94cCIOGMM2es
+4DoqP+AXvnkPDdYLWQQY48KCedUbAVUo9vc+0dQY7A39XdoEIQvXYnc9T9zqBfy
dgUE+1hMl2E+KXkOaGVAuM/z1PwR8XLFF7E1Malf9uCKKlaooPTfq8kU29LZoOxu
w8LN86Y/isASjIIWJWAGLATrAcFsyQgNwdkSo2yhrOpf/i72CRaLNOyy0SxuXP2w
5TRmvHvxL4uZmmEzBb4uivM/jggkv+fx+w03AtwPt6F53JFSK3IXKoO04zG2AHXz
BqydxThY/db+LD0a1BTqO0TuA12xrmQh5e320TWxySdFou/+nDYYbxpObBzTwOwg
nGhapJyidsX15/58iS9gNj5nR1artJMIMNJ171NT0O7+RWVyC6DIcH1eKs0dKlGV
LZdcPet4ZtFhNyRKbtTl+wGWmsP+dKBRYM3lJWmPtbSvtHE7I/IhQZ6a5fcJFMwc
7+UOGNHer3MKtLBWDVzxYaC1LiTKW4zXo6KXfI6ZvGOFfgXeps5ZDlgCUA9Gzm6d
DT68MdyRQbz1PqAOj8eftqFKtuBhFipGOXVgJdGRgRyAvVdjHfkZ76kNs71n56L6
ecBz1YfBLFNboicmQd2KYx6VwK2+FwEMWh/UYBwzx9RGnpNPkf0OmKJeLVthhSS7
3oU9+g7+BlxBcUk1ZzDsoxNzDyFPZWbJC9JFU0FEFC4DCgmlbUSiMR8v2yM14rJ7
lG8pYq6laOIE3A3PihVtODJlH5yj+ZZYE4Fr+QQ+rbLRpADuy4mRLTVSe8zqmMNf
Ap2wuOqzDWjJC0Kg0XbjH57JrXVl58qG+daPTJD4jzNqLsluSr1D7+rWuK75KhcY
z6ygwwkBEaDz+E+8+tWsDC8Guhufb88tYeml8Q5YQVi2RoBpLjvH0wFLhednqh+p
ZqIG7NZwkSHk1K9YoabVfef6Ziv00MWm6GJNG93uPh0rDSUai/LwXVqQrH9NTnzo
0iexIeARC6+8hd/QdaEZVVUy6uH+QDJ+NjcOEDv8/IacBLq23cekX+4kr6cs6Vdy
mwVhb9OBldbLS4fFa/MdQgMYBI4Tk9NKyXeh8q3qoLMdyo5KqZX9CW1hOXoYsAJV
Vk6V82Nx0vSZRlIuDqtf5mvtmhKyUkaZnktCh6Ew05X3yHSPfdUc+2Ymmok9cvQJ
zDPZOdgerWxUds3btr/3MAPOU5tF6FTNVqauxX30HSHZMVubCfsG1w642ZFVFBgw
f8SwgG7yC8tJS2mBwGez+k3CSMQ8gb0hQ4x7qNq8Xl/JruJVIy8uMmbJcBRA6bgU
9EZRCScf6J0Ev8/DZTP/ut01cxEsk9tn3/+6KpcV6KNSIchonlOJsWWcar2eTatT
u1sx0YpE0BsXRb901aAOwqd8IVRIjz7r/Bz+hhU5fSW29I8DADpuPT7bPRvzrlxD
OkMcTtc/B0ijhuOypqfU6zHHxrpNei/n3WYavuagGUXQL2hgE4VxEFZWR2kb1Rji
GLaYKkv8HMg/qDPX+FmoMKsRc5YTYs8LhypnyNFEykytP0LJwOETGqx32KFFvROk
yXdUUNh9U2HRXXLLeaoYOv26lxU1b6nfvms5RRIn960MEujEHqz/TRfQndkACE6f
lD0eplLItW5vEay6SAJ/+JGfIXjmm5IdPXn2UTpvG5w8u5aaxfbYI3d9nqeJ0UaZ
/+64S0cM8KELu0fk2dabMDldt8LFMSMCCvJDbyDZY2iIu4WklhpcH61jRNZ85n/I
t9emWRvZvRxCzkAFvyF74cBHks5azRAxVYcNRAghGJGCyhDYD1p5C7kt++5PffUF
/IpuT/9HuSKQ6OSkCQrPNGQU7Ai2GSmP5qTMx9FSUyNo8FrIjb4+Rckc5hncDLC5
TYlNcw/cVWrIKmzEmltiWiWR3SUiHPEcu4A1tkWkOo40OKLDYCL+EZYH67S0E292
SbutGPLespXxJrdubV7K9yqHhwZdnjzfA7+v3P9Ohe1Mf4dDjO8fiB0RF1Bik9xE
3lR78x8+dQIXAdKrwQDRowBJW08+kyTnc0aHEpSF3OWLsTISWgY7Q9eLsdBKTqkN
uRSOWcJYwv6HTlOXTrp08JyRrxV5mQHpWABWcHI6jDaQK1dkNqyRT5dlm79/rpQ2
wGw7A3v1yg8fcrEdvKnez4IxGDl1aZ8I03DGgULRlVZMmKaZL1+nQU6a60rVDBSJ
yboRzUBhWn6mPWDE98B/W5AcDPKaucr/zKnLHgF0BeZTpE/JduiXEuVVF8FRL4i/
gN/zP4/zXF6tiz4SLlaCLpvlJT2Vwzx22G1+77ELGnWkB8KI9McuaBrHoHEjA+K9
0o+oJ7sUn/uz7gyFbr6radHaISi/VyU6OsFku1gZkq21pISFiEZ2DQ7Vl/MPCQRF
lm/JHb1MLbtPoU7JgmCvms5WZvQtxiatilU9I/m/tZiN+qwinKWA9JOdi371VBzE
LLlgksxhRXQ6CgtKdJ7zWRit83W5WZPIrXXWLRDMrVJJc1pvDumQtgDCRG91eVzl
CfKY1ocwkKsDy+nZYBdbyK9vHYr+KE1LjmgUmn9LH7F4S1smBkjdnLC+XlZQGP7Y
B3uGEi1WGl8EI+T7IkeRg6O/nMI2sc/bSqFodx2fpNSi2kH1bES/Ib93o7JWoJdw
CLmLJU8ziBI0hcojfrQYlINfZysEvAGNfMPX4bkhc6E7prMfOXyyyg/NQUsGymyF
2SlK9I274W9u3TeGTvW/UEfelO+TN3NQqbE8267+Dx90eQdbWBa5PEGL5pDqkWdi
eG8Kf8cbPg0MAfnyf9jmB1SjnVVSciosYrbulwOT+hlVy7+E7mHGJZm1LX8XlT9u
IhukOfY/t4IkQmbWAaD43TgUU4I9AvLKsNHn1XrhLXmYBJOCwF0OjpmfqvXp3JEQ
i/VeTscpN1LsiDldmP43R+Aq+mAtJMKM+Pcz6r7DJErFlhA4uh5j9T+7UH3at+6x
GWz5jnCeQaJq9trf49WvlFxVQpgeMznHnbs2ymPJwkfC9Mq7SpcoRqMncfC7Zl8R
lKQe6gSBZKyg+FPqu7rz1FcuNBY0DBV1v7tl3rdQbM0EcCNilAze0ZeGsfxhWL/m
ARKUI61Q++24MTflB41m41pZw5CIxaf6HmkKPE4fiQwKxTbtIew7Ag5/1ZrvLO9t
LKOzhQd3VVdWFEELpwXKwWXkkJYiIGs8oEcjd6kpmN5OSICDtjV868BZ9Mj9NLnM
mwqfO0WBAwlgRPJ1+zG5O5PrNrOBjekmekbZSEP3mZ/mpF8VV1svNf7KP32dBeZW
wDTfP3Eca/h4Q8NEFj8ZSqgnzocpbzY7GBP039ZRwCwYodr6SlGn8cWOozI2jIsY
ur7SDekSIUMmgAvo3VerYDXCC9+XeIOpZx0Q7jhP4E9YNOEaa1tuALPdyWVDX9uz
w66Hddw4ndzutUd9252spujKWPMciGYq01Rdt3DJlgP+oXVRQEdmB2lB19brM5Xp
FF/Rru57X4+dDo2YBAijJCnwLF2y/2BaQQzEybXmuCzwCOtrAkVOsxkyzToNKTMr
6kcuX42ztxkGgcY6Xd1Vl+sc4bDxerjhfaQ7gNiUosUSUn02mEVNOWslQ6p1C+pV
Zd0Sg5DuGDg3/UGsdmP0t98pO1/e6XstloCdg7S6EyMfkAnz/gm3JKvudwgp3MCD
/0mVCQ1mG8G3L3lu5I+gzlO19CNb1osEUieEe4Q1d6wpPdCYXjX6dxkVU1bE7xq3
Sif8RWjIc9f1oy7htAMTWgh12wTYdGg8QKXE/IVCexsOjWLQoVK5HEX1Q5nFdsq9
G2BvT+jx6mbGz66REwlqlg56/roBY/5G/KszN9JdV/C/CH4SBvJAVB4ioYr3Fltd
bZOfbVJWzwQZTq2qN+tlGUkW2oBEHi/bNppZZrpAbUG2XXoFTXwmMbJ0NK3xAHBw
tBSFr539pKWOFhX4SvvuxHW0v4LOfQ8myiduzI4f34zpUo1wu96Wcctn+xL7aPTq
IONAygax2DngHhNKfRHaodsUEA5maUbHAIuUmgvtGhsZwIHYblNZajh25riPrrQ0
scTRpxyqRLOLfhtBtMEb3ZgYfZDTKtVNP1c2GgxsFeScHt+6Ue7pJ4aRRMfEdjxc
AgWsRvaQZq5bmUFdmOS/hW7TCh8l/UdUE6Meey+LrEiDvbcVh+c+/e4vsP+m9XUG
r6KfVa7jIoeH/IZUPZfnuN+vrriSY6pcHmpM4dLHpvD9Yxu5z0pOGVAc3RhV9NOw
qLttJz1pWDpTlfSS+wktcCqakMSRcImxvM+NXuahgA/hOcRyCj3FDyweGxKMY4va
y/kEIzPPFjhn3qcMMBp9k6gdwsun9o86jFxqJj8COI0jBCnEHevXFLMtRTXX/pl3
J+o24tyduE4/PwG6dXzVUR9peYIqD22MSkI9wibM+hwd9gs/WZ1xQ2x65OECyQm4
eRHO6U/rtmPGW0xksqKQ7IASzzjYkeIvte6wF0DSOqphDhw5qEKDrDT6zPvNYLPF
PvcQQW6JJwDYKser7fjqHe+3b9FV/rWWgxmptiT0RTFv/SF99wgaAxb/yEldkK8V
oR/BuQUGpNltf1lb/Q6AfddEwOvIf586+qu3L02FapZDjPcbKoF0+SKeAXb3aOWl
Tq7+XOIES1gl3AojoS2V5Bp1Zsqf8ZOPat7F0EqFIr9SDwLj3NBcVNn+4bnJRNbi
xmWNKRsg4GwJJC3oZQD/foP2oN/Lspw4qChdePd2bKdIbnFzWo/UFf36XbWVzTY3
NlN/PJt5RoxpOSlhJN13Lw9mbYPEbvXDwmR0ayf0H3LZhrlNVjb6NLmVJc6bAGl1
Fw+EvtgDJD5AS8UGUpg6qcFk0wQ+BG4PnFymaMuwdrCkjootn+CV+ZV22tspQugP
LfR1xC2ggOfoMqZy7JdRi2kdcjQWOSaYcTqw8r5lzAIWlah07GYHnzBRTPz3dfrS
sXWG5zsOjYz86wIS3w1QoekJWhTSyx2xUWU5NwLcKZorZKY5kxP6xZiIa/xiyRqw
Bp+5PJSYTy8FkjtxRUC2pnjEFLS+dXZW3LrKv0Nm8Pbpny0/2JjcSOeTAYxS+G82
fSaa5tYgL2IRfZFieHVpeY7bftiwb2TOdmekdSL2Pc3zhHOOmkZ1U/YyJCsREiG7
3gctSNRUJLlv7d4lPS6MZRBGcZJncGxUPt/mmbFIEUGxyOMuxclSqopvKEUgKaZ7
GQlNL/MnEhtMdFnQJBdZ9e8IeIo03ehDHLfe0F1t6YTkld2OWd0m6vMKDE5DwOv7
hmUJlxnH6gXp1Kp4NDHxzAoRrRaItTL/0gkdNLG6YJn+itHbJyCZczkgGyiEfmb3
9xlWqaSW7/EVAwo1ooKZiC057M0dvmwD6FnjaRpSwmwjxY/OVqE0e5qcO5kgokN7
TIoDPrfPtbCGyN25In0UM6MWxq1X4eqqxN1yyeBINk12arc6pno5DmMWDGgjAuG2
Vw2Y2vaD1zxbSxL/zULhM/DDRzRg1cihytPXqPc412McmivY+Lvx638IacoCKL/u
yvJwau5SKFQ4smpxDh76Gyb6qr/1VyIp9BfwDmJWuxeCNSQSAkT2NQX1Q39yctMC
NjbluqKxhs1Tc7wOC7zIqFukXUUZkG2khk6+hBtdeXtFDLP+r5WzQ0ii0ton54D9
PUZNLUY9mcfGDxxDFITerQFbS0VU/vXhB5kcM9RS1gZQVV+XKata258uKsbcJKIP
cxmJrCR76Pvr+ykhlnMrtbjBrx8wBvRDWeaXcxYZp/3TB+UCBopcKYUlf7jiC6Ur
6+oO/UHvG7XBWiIEZP/0dMV/7+d9/5nGhOPYILpLBip2DmlcyiDskVDYR7sBOJ5U
n1nEpuVUSI7u6N+mbWwDGqBya0YLqA5Li89zAF/NOqtAeKFE19qfN6CjD0jawjQ3
qShaZ6et6jp3SnCRyIIDXkOILQjQ1Vi96R5SwU2HWbx37ZbFy61RShdQrIDT1+1G
YtJJ+zk7JaqG3oaPJy3BYsW2WZh3FX91McEGMw/2k8h7w4aH1tpbTXBaxOi7DAAu
aETBCEc+uhXu1WOFRCzePr4/vCUjrYmLHvyQoXIRx5I3i5gVk7e2lBMQmMlFeEDq
AiyC6i8l43HcnxCxGwP83mIYFcySSaNhRjMfKCrHddxctNxHMe+RTMx6wrng00ra
7Hnwkcv0q/w9PZ5IoK5Vkg==
`protect END_PROTECTED
