`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jI6zSLBm0hTqihjHmfJHJgdXgaGZvlYDITUtovwLKPJiGGSQaEWYJjHleyhY0R/0
Hr8tg/meiG9hN4G2rzcxiBahoYnU+7rVmwAzMQZAvuHpcLifoEi2DiDsGqw8ll5g
84HVU4TaN0X/Uif9oQl4r9gK4T8kLi4CW+VfIghWuG5jpBoQ2uRXVBI0v1bDRHWI
Q6W1TUcQtGnpB4EqtKsirCt8IstETu7I4H1mcxoIuRxCc/+JMLClINF/5PxdHGQS
vNuodoPxXeEMp120KYE4wt/INuyhitzAcmRbeNoXmcbMJmDybzrv7gLcO7Ow1b0L
vc5A4kktg+hwDNmLxKYLjPx7KwaR1x/Pxw+Ahw6gSbtWQ5VW3rDv/hwk1PHWB92/
EeVd5+og8OmHFMCtcRa7uf29wE7PNBp1Ktj6c6FmNhp3nfXYL0xK2ikeey3Z5prY
lWrzRTT/dsKcM+eoPZOyF+SkQGTUEi2O8iO53A6hnvX54rIKOvfOiZbC4F509auD
GCvwWwXtJHohB5CxAy+N6JAWxT2gSNmzOl8VGIiQDQqlBZQrs7NxYJRZ8FM1YFc8
gh0Q0aWrTA2s4I/8U/jbnIKinxAYwKK+Ywfdonsed4hUdANavzki08ScEQvUmifz
FuU1hdjD1+hZa46g545JHnUvH7rV9pgbimQMtxnxV/8=
`protect END_PROTECTED
