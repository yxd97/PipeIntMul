`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zH+QeIlcadSGFpcnEbSp4le7q5Aof3dCGXxXmWsq69x/lexxmmRxDozQB/Ics3p
Pkq30vOHulMU79z2MDS7pg8B7zB65TAkeb7dsNGcz4S7E1is2KorloWv6I/yVbBP
m0RYiqJHiOsXmwNqypuRo/7Q3KpqrAIgzCW6h3Mw2r/DMKwNBb3b2mNjUgezDuTp
sEzgOdA2gRUslKVlDqOhKhx3jGP1QOYt4h2ZGqWNj1EJ7eHj8FSe13Y/YEqhyA6g
ZEw90dRox252xxuxF4KEzGPtNW5gaJ3zkCQz4KtRrvYWJKSqvAU5hv5E6L5nJ5eM
BKJS+ZciyaS6cL7/HgS8Bf0kH43RTQg0SgRtosc7vm6uJcMws6YyuZJvKQkX9g61
jztDakftVEpcV+SdBs2HoWfrXv4TiriCaScedrgwC77zODHM2+pu3x0ZG1GPqrxy
QPkMWdckPaepeZ/aONUe8b14HHebfMSH+MxyhwsCqWcBKVohkJYrA1SUdKODBozZ
NeSdnhbXH5yYvQvoioq116GFBs41EBakmmgrvKg240TtdGS9orfO3zrGgNY4I4rU
2V+GlxKXlqWkYhfD49gyxrpSvcdwd1MRx4Zm1Fur8X7nRwvIpfkYBt9/ozFb2Zt1
CfUwTVhQ6x+kx47bUtPpJuwINBP4QbTAD9ugQwzzcykWNliZfFhJBOJJpObvCxM5
mC4EpZ+lyS66QHpxIfMk95s/5lY57Af5mPKr7JhVVfxQqxMylgPJl2PRPLleo0Uu
TRRQHKQTDH5BugR5K5gP2SxilehPycygmvfnMn6l32J5MSEWHkm94j2CAMYQIPZC
uzB7SCVfvfAAi8vQtCWfc3Sw+hxCa4ai8B9T6RVAAeQ/SEtuAwFofykMvln/Udsu
A3hvlAYuTCLklGz0AwxNaA==
`protect END_PROTECTED
