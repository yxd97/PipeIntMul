`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9wN7W0IKFUj8yGgMy9iOKvw4YWx3bEjQRyWLnXv37ZNY/ZeyrEQ5gJlStiqP3VJ
Ca2RE/Z3dQW3p5Dr1EBJ5Pkq43q1VY+0Lqz55ZO4TMcTrdLnljlq/l3UL9SJrF7Y
TOHSOay1fioH6PArSXMHuwZW+xLefuYi7/ADltZn6DqpwJNU9OeM6W+eOAK3gRUg
56fQSk3VTyZ/odDfRKb2UrLjtkZntUolsatExktwhCnMbcrjspPNb3cseaLQP7mA
a1NVMfucubb6hJjhpcvR6Q==
`protect END_PROTECTED
