`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YL64Hu92aYwAedJ5DFjz05Zt5ynbTF0f/hTrSWP7V6AQc0c+cxHFv3KV5+8gkzhL
MnVAbbm13Os/VGAhRpIvWjjveHgdTaZ3xoYMD38lLxsY4+fkH6swa8FMF1Ekkdnd
vcVmel9Re4bEwQvm8L143z/0CT2XfoOvvEN4mPul9ZJsgoMCF910Bt28jGvI0Ek5
rmdo0zOhTYxlPjwOdQOhFTLTVMfZBBrHQb8WPtljmndiHxwXAm9uSVER623ZzTa/
iy0DukpzArdlIUE0tfRm3xjiL8c/zoQCIeBN8kem8l7IHLqXu3s1wnv8RsqvS8At
9EJXP3LkdcwmSaayj0+Q75WLQ5E6RfHefGN3GmqtLtr7SvN2yH/H1ciZ6W+jdeIl
4XljgKEiDvFMAVqh42ZUjOeWOPV+FCHwGnUJRf2UtpmWg4/Ov0DCQ5LZubmAMF/v
LVn3sTphKjnIYcojZHRp6wnC/aUtJtJIT5DpGWcB9dO3ZKfOkArNxo0t6jsxPNlU
VteNw+nZDv/5kFulhu1gNMO/pzxkcJ4eyUmpU4F/sbAvUkvyy0xlOfRkRBj5cpmP
UgN8tI7tyADBzDAfasjBryTjXV4xc7PqD3cGQelpcT80+vQOsXSYC8rrS1vdm0H9
Br3n74LXqWWgzm+7YL6XzE2iJIfjf6fL5s0M/Fe2bCLfpX8pUMYYwMWQ1kGH8qgL
Qaa+Fs7A5LX1bfDpIz4mrl7w8n4p2T63Nuh01jcqoh9MXbG5JTNpZtRtxWuKYwH/
hAj1EtFy+OM4E/rUABS4eXtl2KkH0axoj5MMfHvJyHsIpx3X9HTAxgqMnewPV10X
ImLF4vqQelMlwKugqUryVI3o+5LO9dhy4+UUKwtgTQltVjZEWaJnTx1ljwh4aGsd
8OluFwl4mAVEp5IOzEET7sUC0VyQ9Xc2Vu+tQwzfaNmfex/t0WShmfTpNur/6sCn
2QmpkKNB2o23V9ueBThKzpXqYY5kqruDkRWON4CdzP3dQOnn8DPjiOh5woRNSM7d
3Q2glHZyFYtg9tWIpJLNDioEHQRvVAOJFfjSKIRrgdbzKbnPmnCek9VjPrATMWmN
m5ak76DIz8AgHySl1aGlNqd8ie5da9i6ENSKHlNeMJ1sBnH0f9kVbvQPuRNYnAoI
IIalT4tfPZhI10C6VXgfP/HQHxyB0ADMF/BLRAYAHPYRbPbsz8HiyiYE/rA7cvP3
LgGp+ZxV8BnupaUYt47EbRLyA6p9PnRm/2PSN/tEtO3hOiJaldGV0DOJMZqrQnEa
EcXvCv1zdVYxsCU6GiGLFGUCh9qUqn08FFvtZmU7JvtG5TBlSI5FOP3nhY13u6Gz
`protect END_PROTECTED
