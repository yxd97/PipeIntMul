`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64vUplLSRp5p56gwSNtkkpt3kG4xvVIcJufXLkPaHd4IbRpqyR1kibYQ4tP8moed
aVvrLMICMnmIqhnzRnIhrTj8MSVxKwQx7uxFHDIO77gnJ1n/1qMDb5k1BytYuWhb
hELzDwhBJS6hnFldDvTQS4VZL9rK0H99wKw/hqXbe9B7E84ISW275UzbjIUpbsOZ
Njw5/F/8WO8MKab0qq708+aehMnLR+7QJLaXeFBxiTqjjtvFXu+Ku8UiY5BQBrIj
8fydDfzvdunZo0b7T9m+26u09oY9y+Iuefe2KHHLMKVMukqB4roHhyfwadeVuZ5E
k7KgWNHWSv3xylJ+e8R8UkJhOvSMmASBCmxNIKxQJlYlda4+VLDfbYJL9acYSnZx
rT1f0CvWKsZLOoOF364Mb+ZpC/NS6EOwNTPtDJ266rCVdBaYr6KHx2fXP8oTF5ol
oqtyDjnQaUlYjPBxgKtAoq0fFMM3PNPZuNpphdHF0Cm2DP/Ye81LbnFOvYAGd2IH
+AHRGnZf/MYyCqQ0HLspFoTOayyIjFNu+Y2VdG2pLQtwG2vSFXsjrIQ6ib1NWAV7
kQC+QcoTUShBQDs3mZs2GGv0PBwWYoR6TuIApqos5rMIpDg/PnG3jW+DTrpvZBlA
OB4NmbZlK455R4DoIHXJ9A==
`protect END_PROTECTED
