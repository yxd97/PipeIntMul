`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
klML11uRDNECMcWb+xc5gabPAdfOix1wS+x/EWojpi5k02NWx62D/qqKyFnZXuS7
sZIlKSdPnX2SL7KFGWNgtU3p4gDlqUS2RwX8OlgPlNy107sczcFgOij7TrUIq+0V
+uU8ffTccnPk0Gdljq+mdrVu5t8Yg7T3OohmLkLahG1QE/x/Xy80OQnAM5B/jguT
3vvzNi0vitKDZ6iPwvQdFPGg+TKS+OwW/WKt+d0YPkeY7XY51zFzBvzuNHVegVlz
vtw5EvxE+gyQZsEWRI3wnbp+PMFwlKTc/s/CsFfKCHmS4bZ58ZWfGEZ3S2OEDLzR
8YWmgLU9HwL0yTzdbQgoEQGT35iG1IjR3w0egxB6+9IdX/i7yw3eeVp1pKI6AG9U
cHUlwc4ixE69+E1xLmMG9mXvxg5+WFH0Hl3DoEYn6MM51b6fLiVWyAsqAAnZXtcl
Pw6cnJm8AIMTPp1C0kwcO+AMqWFIqrqQ7YOuDxoGhlgKCFP0LXOIqMSpke8LHzZS
ecfz6fDu3vE5gttBvK1roZk99aQ+uqB0oRZ1t2C51+0UML7EFscck0cL7wCeN3nc
6CtBxCh7/Y7L18i/PaEmxsXljQ4NRNz1ednwHBVkrFu9VpkBFjo4pt8xGpJeg9Yw
ioLA/PyY8f6d58NBm7/kWSzMBQmsWbuon1FKwCGgNleuM1rWBPFEQRzKD6wIDKUc
4m0FWwJox2dXw8Fvl+Tu5wsCWU50U8LxEo/ONss0e/2fvxRPbhnN96UQ5Z/cxptj
kJxyIPeqPC46nEK+oVwFC8g+mpUS9ypJfHy9g8hPZPAUo2mdoT0eBUubhV0XsyjW
RlSgJp7E5eZpx4v7S0rBKg==
`protect END_PROTECTED
