`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ifrqu9zuhQsfdy2WgqFeChCXpf8sklIbJREeoMkHeTWrzICiOFODtE2YEuPZZRFo
ic4WJJlENztDXxDOUL3jYOGUFAGskSRP0ja+tNB5GVIINxeK1lp2oty2B3HEV0xc
22/dY0w0bZTAPwHtBwb3ZMhguAL5YnzOJqN7efMydq4AzZ08N/ZnyIQc8J41lQPV
WKhENXnmzhID5r96nBhp5OmllyVNJh7OBFLjNkLQTrUye7UM3Nl2U1fGtkEmM0Qp
JuyRhsqj935dvYOtetm9hcLSKOkU2Kc2n04/XhgbDOqsDNV31E9M6+56mdRTcnI2
cUef5vHN3d2SMPfdWaxp4ID0B9YNddLfFdp6DkYqt8Nbh1daZfrDQWVNkYnfPIqP
cG/Ua6FbW84erFtn91Zei5P2ammEX+lpyURmVNBqB+W/KKqinienUNZzbGHnPvto
2giLJLLeyZPkKOq96v6gXKlTcgmgJ9aveGruGhxt7lGJeM+Pwai72mhVcGFuU45i
`protect END_PROTECTED
