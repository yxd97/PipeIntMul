`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8VBjPnGy9xljv9+LlrMfVktq4bMnadwbEGP2AF2cm7PcNjnMEHPvMptHTxCxGvr2
AorlxDk/kvCU1wDuX+cfQSSueZ3vEZh4Y8Dn4OHRcxCGAZ/iDQsBavlj6H8Era7/
vuF/BLNc9AloeX0aAnaFf28fSKruQeF2z+Pt41E6KfWmH6A1YMatjln9U9Lkux7a
LULQ2QmcxP0y0bO2cThpj8pGEuIqXJUcXQtyOAktm83qoqQBnCmbg0TuojVXpzSw
zKq/CthWR3TugJV6raHr+k9eciSsDD0ylxMoDy/N3qgnqYc1a/T1cuHPoNZYXPEr
dPgglG3NJu/plMG3yzF7huaMarRzkZ/6CyHUQxnuv0lt7iGBlzB7NPppI0w/1j0K
DHkiFKMvH8+Huz7BtNHG0vxRKlbdBSdHkJdDFcwQ8v0=
`protect END_PROTECTED
