`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rfDiQGmxXyF4hyw9bTugHfYO5fz42SHbWCj7lfvm4SakA1xP7j0zbCTHjHlI0oZk
m6CqsX7bqvVkdU92bwn0xos87Gf84Ku3HaTog7FIFOJWiXSSCclcozeLE+W+oDUz
+/NLAlG9UfXW4wUbOJCMhDwBrTAxFE2Tx+xt89TvbckSnp7rUFYED+v+lIek9LT1
xZNIYmv2vdx0uoSKim5QG/jzSwZJMuq7KXF9A5ZlqyoXPP+OVxEgm97ybviDKvqW
LZ6n3rCIDFSuwBKIYtTZLBr3kN84vcJz+R0RGGJ/4FMoBMm2jQeryTCZdpgDGxlm
3MeUoBAwZ9O08eIKzfqvqOSoj+d+iu8n4Nofi2X8Hy57ON4vRKNLgoGRc/PBSJKi
xRpeREiiU3tEUGTmcQVKN5V2krmSbm80ku3PYq1/eW4=
`protect END_PROTECTED
