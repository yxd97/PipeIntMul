`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9nRc3fBYlvZAAQ76lz+oUe6pAWJpOe7ysmFNdEdSveGrljdB4rHyH9Cr4IWO0rkX
iA4lFceFeli/qrpMkyIAOp3MIkLp5V4z0vqrZQyd5ype4wUH0r6irZrQbbMHjxI4
AXwZt3MpUHq6eHI919kBd5H010/vSNY25IoaOoXBYdPyeXlHykIsEzUC0hsgdErL
gEsdXTrdRtgAUbXMcreuSLA/xIbmhaUFPpK5mk/blOGHpmSYAFlbj9eid3MrPFAE
rjzjbFXnSphyTvM2egYMpw==
`protect END_PROTECTED
