`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSI/EDjkjExDxjQP0I8tcwP0aawDytFo2Z1+ZUNOpFBnHs7o/FaMLMQOSsUCST0s
dvg11nA/01XCoKbpyibZPwgOX9gLV6vOZKkVwZEjF3sEdqVW5WcdBeIuaEMDiFfO
61KbesPhWQIk1CpfrPyBMeGL6Lh2CR5i69GiEv6+4egtG28GiS9J3WhlR2iKwqIi
oB+KUv8ibI4vpIHfx/Px9UQ6JeN0aCLOBk1nT3grg4fbQN3VkLAVzm5m+bvgEFJQ
9pT4gh+lF1peqC3+uHeU2Nx3/+XhkZ/F0DZPgzeJBGZCH7WlIVFSO0l+XF2G+VBv
Ss/CS9lCxS+Gwk56wh2FAY5P0Ua+9ppppj5gMh3Kp3TXRgU0adhh4qAduAC9uhLT
uQFPW1IqUeoCLhF1NY3jh3esqqEvdYAi8UMzgaBl7Rmnw1qCK/+gEFsDur0Xvnjq
KaZF9saE6ccyr7rlg05yRmC+podgB2rX2g+MJ4A2UEmmw/akDmJS33e4/ws0btd0
epn1Z49DvFK5AsQtGJZ/nnCWEp3GwcjbwKzN9IZp2NcWXOLkwqvpqdWVjA5fIfFR
`protect END_PROTECTED
