`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCeY1SM9NAU0LpeUp+H/KQAo0xdiLPdbA3BlV/sKVDDEusACvziAlafrA08cy4oe
c2OPMB1pNSninOIZxitXFFQUA8pbSy4iEWKCrZvinxLpjJ9uQcvA3KNODS3R0MKx
KeiOSyKoOVR9tAZZyHAO1bAE6K0ouVg+dCOWjxxjBcSSSKwzK/2g6fWHkl9uwAIG
ogU9Ln06tFqaAeHPO59PHxsj4gqKNaHKysUhvL5gNwE7eJpNMcT0a34HkHx8sJWI
q5vRt0soVy9Lq8WlUEvrVgslp2JVLF7ZpJ0UGFx82+gNapwcY+ehAmIEOQ9CzJQI
uQL+XSGXHesvVPIyVKmNjlgCEIROD9apejV+JEQbloJfdtWc21u7InyFlJuuAGlX
wMnZWzVeXUSNRshm1272z8TK7YQsPocEdIQwkHdi14aDdt5j7J1nmmG/9QRjj2iV
`protect END_PROTECTED
