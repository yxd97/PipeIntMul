`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hiPYXztcmEqGqtvHz2vMFzqA2XujJTjZhyozx8TrUy4Mye7WLgN6sa+/yEAXnkjl
7zsJ/I6g7dcOMyFzujQf/JwfXv/aUCb1mGXM/r8SAHSZL0WQtaoZl/ifvA3apUQF
sLGnZ5VK6KFur/hHveApGbI8cTNO30lwyY4jF614neJWOyakxV0BxI9r2GWhGvRb
pvK3h9k9n3/X1ZJGUEMVs6ysDn2eYD3pGWEHfKlZsQUcghJkfzhVjtJIPyPVfmA+
aQlfwu2FPseDzaafH8FN62XEwsAhzqgUHCZmVcBnuT5k9jOGH1xJpYi5rXjAit/k
t4/uTkinpiouk3SP98dhznP5qieOY7+3WYiOZI77GTpUn8QIa3GxuQwkECW7ouQQ
L6tilB858xWwlkc1IqdhWwlJ1IooBBvhmlPCy6R4XSSKkgq+WJ/SPksMWAidilSF
`protect END_PROTECTED
