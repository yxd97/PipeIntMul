`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4Pr4hh0t5bxH4/Yf1UjGeU7irxsFEJHxVlzUKZU+4fezXC53sUw0BONnR86hsUw
whgVhmiOGxcsH1Jc0iKZf9T4eswNdKJSysJNmJJqJLwLI05vR7f0pCEtwaYckZM1
4q1O9vmMCqh3zATnklCr6gXQGj/bclIqB2v6gT2OwdElMeRuXkJW09rB2wKrwGLv
BWaXaJGfAacG0x46M/3FYmSJsYoVz/26HS0mgJ2CsAI//d/njvCaG7VFjgFiUMzv
3Ho+29OpICeqeQs2F84fST6DboyW/9WO2wESjke1q98uRZ8VmJU313Li/JrB3Bpq
Z9pfMksibmSi+w5SJge0ectAVT7CiBc6AsupzLKQFpzWYnccB50dp+a14gqUsRcl
mvxO2PpEwRc1EqM39LfOD2FPB9qkvLNy5UIcfMAy1hnWRadfTMCpZa/pVE3G4/kb
rLc8wWNMA0I2y+4SoEvfzw6tjRm8EnFTEynletSLtQxL1iAhSrZhlizOW4NMTi95
4jVWnfJLu2G4D6/YEWfMz6yteyuBVxvagf0ILlQpKSA=
`protect END_PROTECTED
