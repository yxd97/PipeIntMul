`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0zx3tzYri1Uyzkm2sf3g/Gxy5hPnt2D9GA/AMpfnEYJGPdXx9XC0sbwWKyWGR3WG
3Z/x7D0KNiX8c4/K68JbX2ArE2ami8sPoMZcO79n4uwE4Xj5G9sMWEb2pugpfL5m
B7Xx6KGhgeZ5pz+l4ZS9sicGvmMe4EU5E61S8NxkNxuRPMM06bxK65E91oD3/th0
TkCmz+HEzrmESN9cADGP8xLxDjSx+fLYzTbsr9NZEOedZC3lyVfFf3p/celCDXHt
Tdk8vHb8RwGDRm7awZvPxpX0dTFS99NdmJGtnwDGFL5iQ8pdWRorutUAPSzES99k
lcBSw1B5m7jiVaB7lipPV7R1FXlbrrEMcevU1Nkuhx5UmcYkaAgoT0rcTB9PYAeH
CVMc3RY+G0FN726k6VHJjD2VooX3zL4HckZheRNuW9GR+Dgl0NBYxpdOi6FBCUgN
SIBK90+gsjVw8kOvjJlo2IyCewdC0m3qYo2QP+d6r8XZFWb2adEszsuM1IBHd05T
QvSeN2zffEBKCoCrUvyzHafWg7UoHM2PwP7RTzuxJrTyAo+gD9jVtRBU/lNfMphr
VXV1mnE7qvhZVDyNb9LXXRLdIxEF2SsbfIeF4eQD2kYDGm8sSB1leggmzapaAhWr
/VSZhDSTnvEpC92GGIgWbgAJ743JenwxCkWB6g/WVns0jG/RrnANQgAkHF2FBRQG
ppE3gMF7OtGek4ayjiKM5khk+nKRCbg5AJi+TaHwzw+W5uWLlR8aeMH54yz9tiDJ
WFmsWmenrAtCvAEt4RhQxg3MnQ5C3U4trFNiMaq64XWNdRQMcm9vf/dqcEbGK8j+
FK0fScWeni8rZ/jHsg0UhxipwB40dHJgdlGapPiFuViKZbOK/nvm8WxIA0/hcpuK
JRXJNUGNNyNqcVQknatKDkN+Jcr/KcfaPJ3jvbZW1Y8K0iLrS0zs/Ix72SVeeyqZ
VTWVbYKxOC5oQ8L/stDHTSjHo2jj+iAkE2n3cWICMUbgUXYShCpQoguv80wCuwuE
BnJ/h57je+U/UejPWU4Iy8+9dXqpOLLivKtJN1XpHyoMpTMaWqHSzlpZEATjahfp
lptl/lIBVITiRh6C8qx6hRCHgX4aWvRtPCsxpVsQ1g/+0QgxJEos7Aqjwnt/kIbP
28TJcWVPMCSyBE5Wde9vO0l582IpoLd3SRMTLAHH70nqbP1vuCqhHd9L77fvK3vg
M+CIt6Sh8yXftVNsrrHcvw0/986ZQfKrHwEdckKhE3IMW17gDxYQOy2vvY4ymY6g
rYwX/Yj5tk8goomLnHDGd6zPVS13ff9NpSCJoKcZNXdj4xxbDvDcFl8bLsQuMY/2
dohvQBuj/V56aVecu5LNpg3zKs0F+R38XHoCapwFiGXkJnSKL4eg/MMPIa/sIgPW
J+jHymPCvrWRlqGwluiWHxK0KUa0yiFFv5kbFA/0/38YsxIAtqeWlSUIIgnMVzQ2
Dyf4GY9lmbmRSLevfUPD1w6JRACYK0/n3OjyXJrKix1YXUtnNpJfsbRtRXdKn0IX
ARofnNQ1JqDyCzlDBLmS8dcAh7DbtX4teXpMG8Pcpd6scDQBCOq/7zysveHIDm5k
0gORZ0ftEFrCjsyARoC3xvCKFa5toLAEo+rM4nXQS75IgH/UYzmZqsMfEHLzv8Ps
KTwsqw/TszoNOTSY9RRZiMeLauC4q9QBCFELPPYhtUHP+8CuUZgeTzu1Rhm3UKfP
GTPu9MhXuQyq+e5ySD6KM41nfTCgl3GeyT1GaF2Y8n4rVfC0iq60g/UhDg7aXYwm
8dgPTbNVEml3qPAERsn3rvZj5Y6dAFO/x5SUiv+KiTJYriuzcNcN9VGGuzupjM7c
Uj3NvAFPFBDmhC52El2HYc0R1S5qVnGF7IBJh5vQsNwuhPJzXqYyrw62Z83JUKhh
5E37+otz9bDwrAIs+CrjpoLXQRj7IfEJRS2Ky4XOjQzJqsqRXKPWMz6t9rCYevfy
eGFesTtSc7062nc36PM6n7pKyZUv6/qCydPfApH/gUBfcV3QQ7mlKe206Rv9mV8x
VQLP8Rdk/PWs3rA/e0+RuukSGDAAB85Y3NSQjc2wEvET+piLZZiGEm7PEhLA8kQG
+wiYchQOEkE77i5yS6GhIS57SjyBVnpGcoE8u3PVMuVFQEGrHz3fTHOAFSvuyUbu
ob6wfxd6XMKjorumUOcUaE7GDCYrd4eJfOkZuXQcD7TIClFMm+90qHIancIra0Qu
huOwHJKbqsVbLeEFks/1tPsGVLiFLIJUM95AvX7R059PvEX8i7RDb61bBnIE39Ad
YQAnopmyHocMwL/tS0BkYzitR7D6m8T2wH0PRsHEl84kW/fT6Y6y6Li4CRGpgZxQ
tlda8feFItVEmpQPNaiWfqjyyZz5J7q2DU8S1hMpgdI0YLb2xHG6cLNCmQa2RcWg
62L0xEDlNrkFkRytahlUGRK8tEFzKwGlOoXRAo4PkW4Y5fy5/7S4Prvm3/YMddb8
2X7LYkOM2/8/WTnt4yp/uuFT2lTlj9hEFhBmbbgzBlwcE4DgYycbKDCM6AO+DqTx
bNuEaOigiZl/pMTmFHt5BCyGbsu5kyt2en0riBR9ZD8/7K3MqnGtz1Y5mkgVfQRE
U37wRvoMmo7xTT/D4fjfW/gz/cmX2cJmFV+QftMubMYRnwUkHAxOn8YaqaITsWaj
py6+6nmadl6lYCFvPHOe//y5Sl5bnIT+dW3CcYuVWyo98njJkHFT+rh9Zair/eBv
sgpQ1Vve70HN3i8EiEdRCMkw2Ks3havQkt+P+gmy9oigQ+89xq3DuRK2EbhvO+7B
QAMVyMiOqWDrlKni8rTImbYpSlbbymnU1ZH+Bmh6wmT9/aq9gamoYL/mxi2awyVX
Ym4jXdJ6ckwdU7yOIauBgXTCHkAAXuZAn6ZhW4dEM70q62MrwhYKq2y+bt6Qpndq
1MxEnNGb6adc1lGOg1mF17XRkB9IwKigbzGnDy4guY7rNUWlgQ2YvTKbVNBGT408
p9XSO02x2pODYEyGHwKfKb737YMgM5k/qnNHLPrHi5mqJVH9nnPXh30flfZ0qklK
gw3p0qJ0lG+Ib4mJoepqXrKMixNyze5Qa9Gh2QEzTRmfc4ElHBi6Rm6gUeK/B/2S
LtSqsSBZJhDCD9ax15uvZaeeNB79h/mnWCYu1+eELhcDpY5s21zZ7lHTU66735et
XUT/vGC+Ggwd2a+GR64PVNosClEUJKyjLE9eyoyHB3/Fi4y73a8bQJodX9MecWWh
Pyt2XJnDXpUqEYAZ+tj+fgcGxqAKDw06T16SApq3WlyEWdFNs25VjTgMSHedk669
DOsOYKb6EMRdmVePnUlOtHPeObVbP7UEx3YDpCw4+ewp+gDi+AHaA0mOXEFnBsx5
iQdixrN4ZRHcKVUyz+tZREqazvXmyevntLQ8aY2Z0wdEety6gN2/6znlmaJCO2eP
IORzRxDIZB+AygDvffI2EDvrOFkHDXK40X5V2hO3wRsny3rgVbv3y8i1ExsIMCKS
sAuR+9m9UE1DPtklaIywoZogUm/cbVJAeJxt1J8l+haSDBNU26VbEBKrZiYND1uH
0+6/yWoPhfyzeklXJjPF46D+/s/qkEGY6tHAIsaObmLXkazLBTKH/zdpk5lgPAtG
PEhX9XZHpU8/X5T1JM1vIfGEchThSX7rr1nzOXZBE7R8ieC8GawuKNhHX89lXTvy
CL1VM/AH1iaU9y+Cd2THHrdwNlkLjty3c7QN+CgtDazzwXP2quz+U5oEcg9sJqvp
liaMqrBX8wXjibpafFjrc3bHzeTp6XD/dIGvDkbeCbO5vUpTY2wa3xkP0j2dTRmN
PIw+ncEoUEjNR04qg6ZPIwjPshZr6AzHLTz2ucYawg2bOpuXxhSM3TAYsi41Xn2r
tOEzHIltDpGo6ubYQaIP2C3O/qhj4wagLlgF+SwV5RCubCh3eeJPxpf9oCQ46JAg
VW2PFqNfujGokvyrpEQkcqV1jIBsDrBacrgBpQl4496LqcSsCz9EDtuk04y8wtuE
LQ9NRDELN/fM0wwA4eF45XR1SOfk3FzXJoByM0st/Z8EbcoNzTuuy7aQ1+R0TJpg
hMh5g2SEFJCR9HquczSTpt6JtglUO1o7HoJ/Hzj6vnQKFAzPcRxKeFHS3GyrFfzZ
DXjoH1lfgcyM1TylBjYkO2g7C9ib5fothW78ujYSyp9Bakft+Zb+LdEqo173v04o
EZBEDS5bJ9Q857cTuwZloUXLQPQoEsMQf1BH1DkVyXeIXLdggU+sf+1JVxr1NJNH
C9CvvDNN9+Z4eUQmHe+pJYeVSPvgSEgDZiim5Bm2LPpEUVytPYhSF9w5V/sdlhCC
gjM4Z/84fQ4uxrHkdv38b9QCGs/hq1ll23IuO7uN0HrA8ZYAI7dur5Kv4lgqKmU9
wdwT7HUNzx3Yjcvp9AAA/sZL+XNo7rbGqxOIp22Wnd27K0EoDeIcR39WDSuUS5nX
IeE0AIudhjc5mtrxo9AvLeTvzzCmUVQ7n1vfWZglIJQ9xY7kx+HcRglxdrB2NGKs
kYoaA+Bphuqm99D0dxjhn3Z9xDkcYgnKNOtTQ/E8mMqniro2p6a3s/pDBc2txE7T
BP7v9G4GLlf8qTgFz+6zCf57fPtO7F1s02hoauI7SZUi+FZsfrwJNsfMaCN5ZjP/
L+vLs6TG1RsQgOIgMe5/XeoYcu6+9IXXPH4PExVvj09N/L0SYAC0GC9ly8vBjG5R
FZDL9jzutJxwpAKKnyo3FPs9Y8eJNXKtUZr2Tkhyp+AC8by2om67gwtbZFvVMIld
AYqRnKJSNZBWlH/L8Qlff0ywiosI8+od7dANubAs9u9pdsJDdbjqU2pLuJUz3duw
hoxtypKlBqadWMsIcMVdu66w3Fez7TgA5FadbEDC9VqpRWTJ+sSRuwBPrSFTnRVw
gg7S81rcXbjd99SUqJc1G4RJpiMwwvWhpdBfgrk1VrmRBKNVQLlYkD77NOUfpa5Q
wZRpyvo2j7orIGrtfv/2pUtbJEOV9sUCn6AxlcUfewmHjtTJERQCk+5JTZp/kt22
rmDzzexL1baRf2vG2TWa9//0lgCEQvvAV2ldhr127XjTcMaT/nTu4DUWQIJn556T
/+9DbBHIoeLFXwTA7AFT7lIsWzGWmOFL2GvR6gXS8tPOrPLwQwNRPMZGkpzZLEjW
rZuNV31kIrugVmoOfIBVGDPYalUo79X2c4ht0G3Ba1cICT46WbqSX81zT4wEM48n
q3qGMYwGq5f3oyL6c+fp8tNaxX4xSp+JULapFHuWWrqPVo0gtKNE0pq2c/ycEqgh
EExQCQ4lNZPgRzaL/+DLybGL/laNuE8lhLpEWVuQIuSuYNpm4QWdprJqJPhjvndj
GsF1sfpFJ5b3LWW/RD/sMgAWA74py75lOjynJA03nh5b8W+NXv/wK+dq9M1JOdrm
fdicGM36jdCYdxFhvbEfOXHNzifNRbGmoZOQMn1qQfaw4TGJDOq0SunsNMR23jng
dz3RXF2CwZpheWhgK5jq/DTmlshpdTfN+R4oQiFsXrQWRAbYKDAnOV63cvPrwVww
+ZjMhOFQf8qr597S+0YoE9vog5s0PSHFPX/E5lJ2YS1sHlB5gIHZJscw0UAAj5f2
OYcRqwQ6BZoI40BcK6vOKyPJWHbShEefs0IDcj5Xkw37NUAKRwXqbxqJtTNvQd6L
cvawuhhdfUl3IAb0fUFa4cNkfTFEBPNE/dWyfB77lhJXM5Hdrv1dVcY/bQRrNe3t
gjImZpcq6CtZldFVedIrjJzn6CuuLMM0BQ7uaquZMOVMTgqF4DqwvWEHd9ySdgKW
3Ntvf+mO5Nkl/jhz2+NTjtLK7pcHIDu/T/zFtaHSydhqx4efd/vwFohMXq4dABpL
BI41a5ELooQ0SLwpBvF2j9XYy3+eLjp5dtlkxl0Ig7rt4M1MW1byJXQHEfvqphWU
7e+OfftTZqfh8Uvlr1bywKiRho6J/gwsqoqu6V9r8Ywf87Cpe2Ggk5rfnoESKoeG
AtZm+IcudE1BuuPPWQNxuxk+lMkUwfG5oGrN3M4YdTyjUepGU6EI84yK8v9L6BTy
F+0soZYqNGJGNpWMApxh9X+tzbVuOO0jqK6AkhEKm57VAm94ZjWJ42lgziHQ+Thv
RO31lfsVhMO4VH8Rg/ZOQIySn9EEU1ZeSkeOTvFkitdVvx6i9Z/eyl5DRnfZe71V
4L5OllSHzccK1z04mG7poq+v5ftwOc5jJExsQpXu2Y4jXPiCrrYalnqoZiT3O7wt
tm9pg47c30uDqQv4XxD//UakFMAmEbvNc1rAtwtb3ISK5q7WrIvf0Jlfpvb79DSC
N1w0T6dhNCaZmiygZCGnZGRKVXBvbIVQoCV1yYslYW7aLh1Suvxayt2VQSNlxFqE
D8XpJuTKTou1ED5Si/SGKjxdGJr6S63aV/7A40flSsfqJVeYfIo/A4zTQEYwxWhd
VHNuUFN1LaFmrBiYolvURwfxChX34nu/YgrNps6pHq9pJ2dRfSzRftk8LnX80smF
9mMIitWHRDB8TL904sQUKKBR/72kRPLbDkOk92DE8/YzkhPUZIlroSMEungzP+aJ
Xzqzp8kgLcpzRE0i49bhZt587oFyr+5zWrdYIPus4OXYyPVGAxaBJVMvMsxcjKqe
GlH5Ac6dbx7VBvgMyCgPYO7lMW2dCUgOWkRSiLM3Im7SDKIn50AIOGcw2s1I4cyv
pnLVdLpcqn4ESAdlKOVlHgcWbsKYMp1c2pssAbh1nCZ1pTc74yFsrJAPjWQXM1yd
/hItkPvY6DaQcafZBuTQWZisuebq4J6GC/yZcEzQVJqDdR6ybgj/pV/U3qX0Dy8h
NjgaSnaUT9jO3YktfDXrnsdGnaaA9PVA6Qvgbm71teugOlj5Sl4wazt+glfk/RsF
y9nzl0Rk2IB2HlqP6ZFbOYR2sD3KzgvuC1hlW+ZY3XEDuB+2UdlYVSI4DApJuM1t
PaYXCbdC/R/PB0wl0vnADbRzRinGtdExnn/Y+GjmEWtKfK+ABhY8oubJxSAJSOxa
unfVPAfJwU/gtqokb38F4201NlrhEv+spY/H2G0SYT6Xjv3I9loXdnNKwd4kDgbr
I630tKXBlWT8jIPnWZHa3DQ92qt2qV5IgIrA46jCj482eJBvi3AhLHB0PpnbVo8W
Cc5Xebx5JeSt49tDs/7aW7qKi8vk8XUaqlDGx6wSBrlp6VH8xLfynR6nS6w8YApJ
67hJfoCpBkG+zp70gAr2HwpvYluXj9JFsEfJgGtHYSJd55cXXcjmSsjipdQUXZki
+6nlqXfYDr75t3T5dfAwLmgRvO2nkAYgJGl+DRFnt0sVZxlfcbSp//+eBjhw9ZYv
S0KEU8ZnSKuans2XffsIEYDJAELhMlhBN/0jWC8XRcQnQIW4kN4XSMiuO0Ay33gP
xGP19wSPxASA4Zvrf9alJffxADfhH4Kf5Erebuy3idJEk/2cSLuDF/xzgFg0sO+0
Hoouj7PbCdf0fr3UEScjQBGBAJvz4Uq5E4+cTaaMVCRDv6kD1btgzrb9R3mKYSIy
TPjv6g9AbOlLjHDOGMY46KG1uXPnM5fVL9Z+sGAEG8vGanoHmGgzUzWyg6vSKEVE
rUQuLYR4ZkeA170eStHEae64Gq2SpNf91I0S4629K/q9XlliiIUTMeITIs59/wRX
7bZ08AueuhjO6evUdVr3MRqzr+cj9HxBPurTr4VuTbLsHhG0JF3gHw2tMaHaf/k6
ibnxK3QMIBcfEAa9GNp3mluCRrKcelduhLx//X3A9MoWqfilkoKr9LntM8CIT212
cTfB3H+E2DSKUmiRSJmTzNrftKgx7i/amX0lYxsc5Wk9kKBSgASiQY64R7rQ3uLH
mFACjGDEbMUT1O1sAjCBamwvaw5BjcF6AF5nksRASWXxTBe0dQfZcqVAix5nnwYD
ApaGL4t+pHxc7pmOVu9USTQTbhRXV6RwvhBr0Dq7KQl7QECu0+nfD1szikmFmRqA
VcsR1xx5BhaM2eFO/de0yg6wFf1WATUCmZvA6ksUyzcnJNPxNE6Y3V/i4hmyyjeY
q3GwZEl6ZJ0fVYvoIKP3I4ZgIjZFd70MzIs9USCxTUmmCPA8vYBrTBey9LKoQ/0G
TpU30rtMcKP7Mm9jHoliWkXQ+4Fh+rXJBA2rUKfyGvYWgAN8aPPK6JPOD3AECNk8
Ogtt1E68mQHUHy+7UGvvpRuQquVnJ/BjXutEt4Bs46vbqZMFsiRLlAwvmxM1HP8L
rF0EiXmH+z8hapsjOaXQ4xGq74CH8klQgG1XxbimNoYWNKthNO7vJARVaHrStnNB
PUhgtC+ipTrXg/T5xN1hNYGltADulBdZxfSAGoFd1aCmKgm554b28RO8JHnPL0au
kEI0bBdooOF2MAPgxA6IA24xYSsFY95i6zfK8cSBsgzQS+BQ2/XBn6N2+ywpmBkO
SnFmoFOgTpF3qoQ7Awp7npK5tXtUFoJiEwgHpB+0tZPdyFYbuuCcW9K1k92kUyWz
+X1F0t5vByD78LyFU9OXoqGNdw6FdEOYDwH8ZkzZ4tC7ZVJyiS/634ADr+pUNczw
vueMCcCLHF4PAVV90b+nI1iF6W4mjtJAqNYvXpXZ05FZ/GWOfY5ukJpERX50L73t
X13PlS2JHWgkx/xuU/iEhnZXkRoD5ugxiejn2ud37NkOq3+YvlUVuK6l2WiPuQCa
wZsYroXzbG+E9U6wDsZNgB++crWDvRWo8BugmfHMOLAp86OkFY4Dt4UHwOIZKeeV
TDMOv0afapyRyOpxj5yaevUsPAnh8m7eysSTskcrztISj07SvVOxFyvUmOO447CV
vXPqPjBarloeFQbf9cUqqKPVYNhgGVSNW5yALEW++RQ9efIhsbuatmmzzSiOEH04
bARM9cLiTjhdnIGmQ5NP79g2gCt3HQMD6F4arQMEXDYsxwdxX1j0Y1hSfxIPFIqv
FD0g6OxI3ws72K1yUafrHgvv8oWoztF9azjFPXe+LBCQBrvR8YlN1YQ6gjxVkxQL
1nI1aCaSthz/XBG5UgVTqkpAK3pe7Yyj90M62jMUKMVLtnK9dHXqCdISFMcdV9/E
zhDN7Tg/UGz1i6JgA96OYvbP78bG6/3AtftUdnV0SZJBKopDBG1yqKqMK4Umy+hF
eLjEz7w5WHKMZ4xo793+qUOjPjE6KS6tvlCS52HXjz/12gGZKVMy1ZxBR7+t9cwp
y9NtuCs5D36U7OSe8sHV+NQCXcgALmFLz2XUH00L13v4R9sTcIVYv70rZLg+WgnD
zXeKlpmlZA5ZsGnv5n6/wbXyNOp58AZ/nY7zjTBvrPlr0z337IEwbOABTjTOlPws
pRR5swxEUrU6bQFwor2iiGx3WYDS8pR4HtWkusNmpQ79j9UVkDGXMgxrYMdcR0Nk
qXrXyk4NOg9X4DUKhpSY2imgxlNRiV5D88CYIEy2ue1VmU2FqN4M1UlJlAzareKU
6Ep6ZQIMMiWQROOfNjCPxkbzAl3ZJzL2POyeRVu4iQCA9+W2b10Rx/b5sRN2eaHc
6IWujUtPQr0pbouQKtQKJ3i2JfvM4Q+k+lqNo/E8fIEYLyckqGkqZ+ci2PztVcaa
7booDWSIvtIOLiklE6Wx9UAI8J1nBHmZaj07Vu17y4b6QryiIJmaUkh9lSr7FmXr
PdEibxOrOgnP841cUB0Z0cQLuUqylaXdAzAeLkUxu4RsV3Hy94rGsRvg0LTK4t8q
qKQkBokyb3+QEiaO/4tVIoVEruYz2o/ftHzrUnSuAq88QiiTSLI7IcvhaMsbVuJQ
mIWEqbQ1aFx2l0zL52XoO79I629axEmUhvzGS9RjXLwaf2kj2ewkqo50V/1Et9fK
KnW/BkEyU7IN26x7akgbAS0GGT/Z2IBjhjf+ujG+TXX2MQGY1cOLT5gKt9KCd7+q
YAgDzpw14y3yxVtKSHc+7Pih7Hmc/D7UkprcQtch4v/hpAOoCXAiVLIJUoOPAS6+
C1Kjcdo285UCxPQLoGS+ssxgOXc9tm1Mv1EwfoToJFFALXLtcOvGDZlyGvBWFJCA
gDB7VWXvLJDgmqKRmrMAn3uvfqQ4SLftmRf97jLStsETpJy6i2fQikkv2uFzMJKA
YHJwJ8udX4lKC+y/mqqmUkmOA1asaqxl2hSHnSI4jsijnGlsdt3t/AoZ55oD6aMq
IMHlBQNHCaDvoFjXCgxGK7CYauICq18Rqdp7gmymQKdvn/+icedmAx+LJTZzUdGo
kp4JWg4kLbmJbYnS5tpQF1MYZrRnwMdbjl3hVQaEbmSph4LBoVJOy1ovFxxVW7du
rwJOz+gIGcVS0zlPXgwqg4h4mUqMbZysYUBNVm0It57Ffaab8n4b17HXV/t/kyiG
Ue5oBXBVm/+57xpzTuxfZTgC5MUNDzJWUzm5RhvyOZiUt9rdYIWUNT6d335EdeiB
nIc7suSHLbcrkzf4TPFN3u+ZsJpj9/FxqJPlhnICwjE40qKQY/wFNHuz8EFU20ge
I2BTiJ89LbvVj6a4xzCZJsWuKHAWp8/oVau2wZ5IblGRZpuBw3Khdq6O/HzOd9Lc
u976dpTbi13M2zen+FuFcQGz/leCs4Xg75N72CZMosXTmliO4lN+FkOlTo5kcfOA
gCjGGH2nKTWMuOCjfwSGCFoNy1RWS1YrvLBMqhtrpLTr3yDm6DNbDaT8jFy5Qg81
YTLEjN/lvDzv7EOg0ZP4HM2JOy5L8bXfKo6zWoAw9hrChH11U5rewXo/iRFJrE1j
Lvz0sabEmD+KB5ztg7ii9C/kAdA8I4in404c2ZC9wQz3Ct7adJ7fCDIW7VIT1Z2n
XgINdg5Bwg6Zq0IXUs3onmi+79TmnmE7Bto3PGGw3Bc0Puq/dh/jfIBuATq/O/Ui
ZOGEcJtIUgXUhO2eEw4Hand4nckl+0jfvlIVtFc21wzyuqqx9VIZPjI43EYKR9ja
KNTNYKW7/S6KsFL8RlxEHJ5AoGeTSuuQ63f2kiUJxXu/Fn0JZPOPUGTZPbaPNhmU
gclGo0S8aAe//w4kCHAgPNSwBRYS90ZATalYkZSLM6N1rryIl+hP5s6n/tZ4DOMG
L6A3pC5JrqYWNSfKz50krHj9oNBsVZgxp9TbLpMthArAuQKwYbXN+zJAJaUBXLA3
4VvQOe19ybRRgn9KYcxKCTLGaWJGNVY84COq0BP2v4xdh+xnBT6iedU1/9zp8pXF
CXOPojp7B0S/IruttRDlf3gfVZP45cZpKsx6cXrkAXe+ORoEDMCjeZXBj71LhWQ9
3Rt0whXL1Bep7GmkGpNevFFx99xyOZ4r1NG6le3EvxHT/rogsw7VYOJe+c2zPLAR
ZDy6AUIH5dfBNhmBkvlgYosCFtthb9emIy/Ffcf14rL3sjQ9tpjU8QU6O81Ux9EX
yGClLEhkYQeumpUtLJmWPZuFuwbyKBasunPsnQgnX5PpaExCN+LTZRVRnQ0yBZcC
EAMF3e4gFs3dj0cIZl2GUkUZEWZCCFiXI7OBPAipWIgpoDl2CLvWFPnqiPlVLldA
IQPJX2sarequPc1Ri30QOvnIWpHpD5YnjHiG+S97jsrPL/0zwMEeUp1bC+uPxsyn
ILUTGjHXZ5qWTZMs+so5/Q2PTbr+LJrijnG3nxaAWU1F4YzTSLFwyCyYyNmiJR2U
D6s5e/bN7c7OsPr2KyohOOcE3MDvVbY+zaM36v7cprXGYVbEiLoNzt81Gcz1NUAb
CZYgucWoioX+L5vb2Q935U2iP0bSuDL5tCHIS5QTMcBXZmQnTNExVNZMHISjaCMx
Ug3UYrC8zdJPL6gxe5xSVljks1umyBzX1sEtEhvrpLeth3YdZoxP4gnTUjyXMph/
rYiLrhfUKAgfkf+XSuc1akyS2oObMBkwAfUDfzbMhb/2xgklTmtRQ3AGJbyTmwWQ
Pkatz0ODc08GrRgnjHc+meSXBQcWwMqlIBMqHy/MHFDrw7QVolVsERtRcyuEfmYd
SPP2dJYecW1Le5NTsq4+O39vh9QXagO0N46alUpURYb8mQfKGD7WjX+fVdmRSUos
nRQMMGqQg0Ytfz2EnqXfGnHhyGnFWMi3w8vq22us9G1u8wVq4WNa1UgthenqcMfT
eYCR+cIzlVt4PJ6zOOCfHxsROlMBDMv4nRfgrc66KyqbR8yHS7CVUC4CgHWh6NC7
086Bbh7iFkuGQz+ps9sGTX9aBHEm502p2jcTe7wXY5zcD1g9RlszOvw7iS5qgJyi
js4de4UctTC0kRcRyLxdRYOPsjqLH8fra5FSLBhF+5KyBWq8Hmff+ooSrJ4MUCq+
yE8kRq8L5cxCmzafk9Y6f6ZpAwjRENZbDTbwGIR9ZtSWcQfMwUYSxOLl795iFdkU
OsRY96GyMJPpISiFK7zwsb2JyfT9XR2q7ILeD/OH0m3vKz/09EqMBNIMW+ZgIdpj
xf1Lc0XBeiUiGfKkiIkdyuxdxXhB+i96nYHQAXpN922YS3qkkoJDrA1GFRnKUZzo
vVhStTrrJ/EFUwqb/iPE5zsR17rk+oSzI10r4Ij0k62l+VF9Fou2o1KXEOVvndhW
SdS9hcvXDXEykMqSpwxfoifaGp11Q9y/P4MVCYLEn8OSYLSdY102GdDd2wk+P+rk
SpKErzXe241TMX/FCurVWWnvatycBlPuSeM7lSKpiGhcDgiByO2Kti5sVHvoCElE
jNfFetgW2PdCjQb7sxnUerwof6lPw2nak9NgWRU8OwvtdiveopuYY58AQRrw7ejZ
lsbL2YVSFu4rj7Eof5LHOChvKnX4knCKqOdEV9mnUVt3grN041VZ+5i3EYiIBaFj
mfv8YtBuvW5WLdEXvfjlw8ud/FwUsMLLz220pcC06ZqsTGyk5SemN6AYQV8CoJSG
t1uKF82H7ebMZZWWuLeVcvWd8ZQhDsGSIyDv0xXOaL6LwD/lFMdGn9gkoiaofe2m
s8Ez1t744SDPAmzU/4qsHn21wXHnwMQ4jF0VrQb3+81VBlofzI+WWkMnZm3b1JW/
marecL0MatWIPEY4AdvABtHj2Wkhxe92Cak/09Y0vHlJPF/272Gxna0bJgYNKfKG
rPwj/qTeQ8Vw4rPvhB+QnRcqn+uImBf/nC6W7NSOf4n9Nm8GnJ8AK6IiDWAGitYS
VCnV9VY4jlygbOL+w1n1kwxXaJWlNr2CExWm0XaKZOQUL5aCcA5de3jL0btvKqKU
cX+vf5plZBb401EInf/FP/MHT2z5WMjdcAt0oLmLQ625ifXxDwZU4PdmKOntuYpU
YtDaif1AbRXZwtN0xG4yDS4s4oH1uMWv5SvQkBMVN9zds/fK+tyd3w+GEJ3/i/Lj
By6ffAq4E/YgtPyTRdnvUfycAVyPWM3CGQI1feQPu+/fBMhWcmbtIzZTeYMC8yCP
4UTwCrESPl91aUOwtu6NWE7B8OCePFD+Oa2dNPLHSdT1xCxIY/lDfjIxOx74H5LP
fRKDE7pTEhe9LazaoQxMCoTgFa1Q/a6v7tTJVfoGnqNMgABpq2cmVgCyxIwOrPkW
3iww9y0aO9263j+fvWE6n+J8l6yEZosF4103MAg4KLUP+CYpPN5fnIz5PGjXbfYi
8ZZdj0pwXrgT/QoLxaV1lDebawrMXQRnPMZG3WFeY0rQr8Rd668C7wSQ4VnDFQ+W
FUCs/BgH7Zv5S1i88EERWFD3KKm09FAEKBlDxE4pu0B82a1AkHT4rFHSeuTVxrWt
oVjShyvVDbLSUriRQyLfeomYl5IzDASDElBWmC7xDkHmIHciZALUqKVP9yT/z/3V
+oYq7s0UpuWu5wy4xYsIMgpYPYPw7He/iNC2DusodAsTUP84AYAi2UWnvHNnurKL
lYu3iXk6jQn0mp2sl+008IO0tXsXB7kg3l/YwfSyuX3BIMHACFn5gR2MufrELNVG
03dTATxIHQIdvZRTa+ImNTIbCI6cyRt8xUgrdLfLJyU7ApKW+80YNtpxSARSKskW
uGxWkkgJYmgfDezjrPe1zaApw2TPDE3zzTXfgjf/Mj5rLTu5AQ/A657dt7GnSRm7
ly+NSX5q5cavqGnwsOxtDcNCZu/swmTg5Ur90rVTtb/Zul0nIdASGR1+cGdm9GDt
nzYJ2fRPNin6Rf3j5XJVs/x2eZcUZdQkqpCCnT4O8s/s9RGuOCkYXTgRz3i2AudT
fBYNb5YewdKMVsoqPk77A7dvEBoSrcWsP7DH+8pxs5ehmyZIB05heRxro8OXRpei
O9gmPJ77bCKMC859wyjeoNJ8kmiUAn1QwLq2dlTYcMTjjJQteTkFYT8sA8I+z+m3
O3Zvq9RlIOaburJ1KqbQN7ZzMq96B5saaEuBecJilzuJmhVItIfDny4YfpJ4xV6m
RzpRtjvZPPXn9MMxBlBtakUCFKpKwNJmzPUTZTTOc+p5d7IWzbVVkXkZ05z4oRZ9
/YR5S04xKZlNpczRE118w2bRZGeJKWPGoB/Q/whzrTIgoN+pP9UmYS1wl79i/VxR
iEvjmsDZMgyxSn3O6bmYafWVbWzobVzzgDIxAw3H0EsWIrdYUCLNdNoszOcQK+wy
QADEzWkCK4/nSVhc/lHL9O0mUxQ7g5MOP+0w+6HpGSLqL1yPMBMHnP9zkKFsrX/X
9tK3IJrly67MlqRvHTn3Fepc5vN8IHo2RcZQS4m3a/VOoOjcU5RCaABXmkwnx1wi
/sk5cyTRlynlAkfGkE//Y5iSH7IoS5y5F5lxrURSENDdTxJULXAItmEWkxXfDnXF
HxJ7mCDAFAgoBUO8+jRQmh8KqGQI/5qNMINRIgce1pZqRYAjjlZD+GrKVhIpXYg0
Sh7DONPvQFhuGumeUeiNaZMa+wQZaTaAaZhtYkbSodcABTIi+oHeYExxYLDvubOI
ZlDObbTUGZXgPENi/pL6qs+l3dV6r4AqDPCoHihUW58DvN1Pzn3iozGe3GNf5iuB
eLMb6Hd6AfZMhW827aM5nlxnJBQteYU58MVe6/z/sA/r5EdQpqnx/KH+HPHI8up2
a0xVg4ISMX9NM2tPi8MkWLzpV9UEsXoRKnQKhl+ggt5kkER4KPpq4BUztbtIWp5b
9+uUGEcVpL5QrZ8pf4pdFK9ttUrNaTcN3UY2h5EHph5Uco2SqnVtp3k632YbXKQJ
JK8PSS1xIvAvlkSes+0j1pk2bLgasjxGVe2dSWwI3nf/KidygNLEM6HdtY4odNf2
2tZw+7N+AGgRBlBsBWt0cjMt4S3PshbtKpKvMBoGhhT081906K3T0IMb/DFtIUZL
M44g6xTSfSsFz5Q2hBhVCFi2GM81kHR1QlezY7vMZdAAR44LQqhrhy/NGe9hRQBC
A912X/jX2R+LYDNeXFE+r7ugtyVBPK/SzQ5hkCThbbCe5G9kyXup5M4shlK7KKaq
q+9kqcMN5GERQlwCCDSZriAyjTPEXjqQs/QNvULzgKWKduQuwOD6Keg17cwD8Aqs
Re97vGopsX/lHlyUziAVKLUwJmg4Z9U0rt5UJVEEKFA5NJpzMdvUJOevctIStPpp
XCe2VwDDPltjBFGBkqKT25sMmXYHICNfScY9UjlDEBYhhxvvEUY600xw1/b5ZRl4
1CBq/oPHid4M0zy3vNdp1kOcA6hVQg2jHItL1T4ln8ZEGQxH8eqCExCTUwg2/6M8
tr46UIKLxgBGnlX4TSZ32nNLmKJWv2voqJJe/1DVWDZaxHiVp7fE9cJu/0mBF/RH
FDD6BEyaWDYCqAe2mad0aZxb/1IBaGM2Yo3PBUO0FVojiLeo6NeENDptinALAKxJ
qS8oAa6JzmxnvKEemSvQfM6J5pEgS5UCcGKAyqsxWFtp1IwvxlXDA5ujkoxa3/Jn
nBxTgfO4dRU1o/QP7pZSLiqqHp5C1KqrdwPvd+GYfJ9E9yXcyueF2yMxB2GM8Tda
2Ljw/ZtfyMSCr4KYnDtSgU0n11AO9Z5LJmgU0SYx4QcBJ1Rfg7Y0dct91mKFJBnm
XGr6f9iY6MTG27OOUoVU7eNeS2y9iZ+thCAvUpOR+5zzPN0X/oFAuY+SG66lNYjz
15mUAeOmWrqllgc5AzMitT3y30nNJusEB2ksaaXzJ0GBFELEhCrYVzDYGQr5MsU9
7xzHrwZbL3Rn/K68FjUm6vNuBl6uxiYg2mtZDCJXZjH59u1hQz8oJSXf6CFfaahr
H/fl+w1vkpl6QGyXx/Dn4qiZk2JNmJurWGsn2v7yfSWTCWL82dHmpQ0rk7dJfYqr
libKKkSGJ+Cm4weqT+E2wR3mrV9g3hXCMAhn1VcWppyit04rGYGfzgTZbyVBEig3
Ext1nwicYpOgBa7a37jJzPuaQJjB3HQ66rhOFWQLBCNHZCUpGD4WNVig3/rUqTNW
5Lt9UN35uCuZoVX+qNdxBP/bp4rl2jdUuNI9zfjVtwW8auOtNh0CMPiNM3ammg3m
kRtSzUR8jTH5aJI95gPxJx34MtDO1uXGLMKknSg/o8nXy/h0dluRVUQFbdu1YhAr
rrW2No/CV24GOBNP2fdEKp78v+Hp5ZFTZVTTbSk0wpoQKJbHR5vtOt4bM6aNyTQL
4L8kyliKce/tyoHVc50QjFVphclxrMVcFsJn3H0t7XOT6pcFgD6cId/0WWP9K6kX
olDVOctGRIzA4ofbkN6FNjYMgqNkoU+pw4Ov5ZxKqaMN1CZEY0gTdRWoYl7j+ARL
3+m3dqIXvLL2c1Czyvv2X1eAAcT/mmHopHMGtxgvzT2q6HG7lC+WUoPEsJ4IXuUe
/2iiz1AoaW4Gw7IwVIYEHgWzkLg4fntFuf3G5DJSwGVR6sazmDQJ3IATt8sEzSF1
VhClMnnlql8ZVlU513u5HgZvk2j2FZE6aggsSYqhCX1Wg/BEixIXAUXyywHq3ph0
US3JXLoOT5IO4CbzPEdUr1hM80vxrxg8f9n9PEr+Qy4O3q3zb1PmjxIvWQgKNz9t
vhVRD5Qo7ODx1w4AV4It8WLxlpmI/fqKqx82sXYAz92tRQzVXtx9UoqQ8uS+1Ivx
0i41evg1/jRPp1AE+3mq6udlngX673tEY3NgoH6P8aQ2VmHMCr+EWa8EC58bvhiS
VqsyzZp9GaToSBQZd4ue+E+djke+xRVDtJYBdbmnmowGCcOXyYEVtqe9KWAgCK5+
xFP4XEt7Ak7F8mwkQmbkXIPlAmobUL6rycaESKhwpanK4+hjn0o3PNNDw7cIBkQH
zHQjGa8yxSYXZqPojhMKPKVyWXAyyDN2rGx8YtRwsbRe48Ayv/yQ9xIIkNhEV3jJ
NLm5zh5j2d7+yBIHHurR2iNp2St2i5LMBy9JSyCqpI2cgRfizDsrJBVZJ671jHlo
sN4gxV7/GyNiivo2eg3ciMiZB28wAWVfllnwasrqWkJMVSCdHb0ARYXcwJNUNgCA
PJkNXwo2PgGDfnO+mha2ZpKSjIDThirojEa9gyLTKZ+0GPq15sP/IcWAAIPdz60i
Cyu6Kw6pHicEuFbtY1Vda2eybIRIn7tTvA3mk/l5Kiwiojfo+8+6zYVEJ+v2PvPF
6zjNUlj1S+sUW5/5U3Fyoh492o+YsOEvt5b9Q6zaBYXoOGRyzcT/j1MJMkMiyncj
Vne6A2ux98aaTdNIItNAsO1bmUGI4zSskOqqoZdixd/5d0/dNQ0X9mQnsjhRZKhu
nEdbENLzhPrW2haao3rw4K8V6Ey5Va8bX39hBVWH850O9bsp8bOczF7bcw4nut1f
ej3p0FQdxZjKfJDaNZ1Um+EPfY3vWi5oYtgAZ8loqUM5e0cb9io3w1NpDo/4rBjA
trpV8T3uFp7vnHIrufI/MSEZRqS7F+4/l+0X0UmqL1CTmty2aCwuaTKN4rhKtnM8
dIOe3TW0H0d95NhVTtjNa8M1yXzQsZnMKd201P4yJRMVadhkXOFl4eb5tqpXhRXq
8rWyctyyyqJSy0EUjWbvXNr+p+VTuwjIihauGtz4Egs5RXjMUtr2UTB2jr8NjX7Q
W8X91RPh/CDu10hN5+NPGH5yiHcv6uEyzee1mCgJ4cYZtwUY3CNvBCdLy5A18nkj
RasqQ0kQzwRoSrYFqKroOvQP1N7kPyv2HHe8v51+kuDCc9DOp1P1CQ7BBZTMX6qQ
wOckPUaH95TwnK1GO68e6tLCw3zUFZHs/taZM2oa93YqOj8seeERZRXkAe/BOtqL
l644qdBSD/1i9QqUFfDtRY8DBQHTwaCRUHUgOUtSKlC5H7I2l01PBEPXeTgcoesd
Sn18M2lDGJ4Q4gBZcA8wye9+xNKtSpbwHsuAG6753SQYceNo58+cNyobehAA/5SZ
FPlx5yZIcL1tr5VhXNwv5q5OvruMNj31swjcCEkUMRX/eN0SC39JxV9SN97iGAhF
qXtW2PPAEBE9qatRmKP9gdWBji83bKWaeEGK+2M0CnXGQZS0SrMMBzuxCJv96tSM
kRC/t42Vmq34nbcwQxmqaySYkVEzq2Tf1QOpVUqKnGm2ZIlqhUUltTuVNMdxYDJQ
+Nv9cdV+sCMAJPuADsIgMi9AaUmHPFhnCklvCX6aMfzYnzIZrdPfiUY2wGt7gEfU
z9CqE2pfc7riAcCwFa2wDtkn+poQgIen0WWWmyfsRr6iZUyl2gAk2ZkdLCcZtYmZ
ZCs4Ynv1WrWlnUsDhByO53mOZjEpy9/L9995cTmQYK5gZrUUkglYwd0/186JwJTP
JdP26BV/3sIjeIpmiavO8b8FhEYV/jZZ1UFbXEu+YM2Tj9hhrl2HlXfaoWMtT1Pe
0eNixRtboBITwEeuCwXNRUuV0hPKdKJVisF9Xp08GfkXDgvbV2nYZZIEZuUKiDuI
v3gdND8xvC2aN5YI17vCxGa/tjje92A5zSRIpccVHv08/5h5pif+MvaFcpCHpVtD
HrchBrAiQ7pbvtpEw8yoGhgNOgfHk/NdVdQsxX1Z5ZIk0PKfO2wcV2B6dR/yIxT6
HK/7FumJE8Soi/tFW8JstIlMTQBROsYtEFZf8NU5XS18h0tVOIv5se43JP9g0/Zq
VXl+k/I/eZADGj3bm0Fwogo4RHdSCFUHqGIVNNY2bqpQFHikWePhoD2jDyARFK/T
kWiT8TTDwmDmFbyKbT6FoZr0H9KZPua1put2I4N+jdZFqkj4TgSeJmUCB0zVjBRV
juRAKafGdYEi1Be1/j6hCFl8ct16CLoIwTus2p6FmaMeMuFooBJM0CRq2SwTMJaS
cdGhg5juPthWyPuY/vQzXDPl4Y9VuDgIXWWPjZuc3hILvPsqRYM9hd2LO8AuLXaQ
V7OxwLJzx6p7m4+B6LdplU0OqLsYxc8cSTvJZROpnJvruEm3H9x9QVxJ6ycher7G
yzzpGGboMGXeMUdFySXm9a7aC73r8Fdmls0i3KMHoCr0aVEHfhVnnGhsvi/oK/rh
ym3alduUWN+9lh4dXCgm4M5uEvwN80VznajLMgvc1IJwUl+e9i9ZzrFnXbDO18zZ
cvkZiOx28UnxEMk/whCEXBiJJN4+A59J/ar1Wjknm2mS4jORDMiZvY1e8heAbvUb
St2VcH1FjJXT/yAyEwSWwXHIQw3SDoQ0GA6zfeOf9vu3McsEgP4c5JPGqLBS4MUz
G9SUMTp6XexF0/EMeMqzDBZ1N8JoqYgIFly6qdPZy51T5a5NibYQlW8ZU5EteBGU
7BdsFHJRDhi8oWwcPTf4B36x//MlGmCVGXJgYSjNfYcyHaMTAqlEAybUlBYpOdq3
IC42P8UE50ppFAhieVhh9bT+tHGuPIo2abw+Re6lzyp1DhwpDJ/gL12W4zjLYuON
mZ1jrVwmzQdUZh4OUJKLzmBwQOUNgHxIJppdNweUkfxXhyc+LBG4rU7+JD0KeE62
odX1C7opsOutaDAlpcsq7E6uOlvWT5EwSg5k0QU6TzQPwUEBhe8FBFgsyNVUKYNw
Ci7dTmO4grCWVOXhDKzyVV/u9aXCrg2LYnYtrpExIrfwSgHxYtcHL7m86Bs+m9Sb
TW+P/5tYNYG34D+Buso7s4VXFiqd7vXWdYhePONrCgRHpbCgrFSbGSgwvbUmmSjP
HVGi1NWDorG6MeY/bZav1xxb99XXgt1zQ0DJ+8OnE4gvEk7PvlfnkwHjW83719ze
0hj50lpsJaM6hiZe+gf5By2SMrdwKQuJuaq0C/8nOE+zDamDeAixVK2dOqyRCvxK
0WXLvEgt2uzGvM8X6wylXLeWX9VJiF93YmFTkW0PkZY99y6uDz0CVRT9GsOAQdwo
S/18gS5nwi+teEQ7hmoEYFMqJwHEFB6gatHo0G/SREQRNQ3qMaFRU1J9bGPlAkRV
uWSr1PxvgeMgd6FUK1ZQYa7kP1kgDl1q0ouip6jyGoT0626byIgaf3NLxRyYTX7p
eajg1lS8cc46MiPrRtXpLTnhlPamiCtlUShhPpczPkNx6OOJuKt/Q3EUKvca4MIe
rqtnSAW+AjaH1BkwFsdiz60c8ZQ8x+24fbud7RqGNtqy1o5iSstiVa4GXSORLZ6T
Lf027NYHaNnM+3/tr9zmVN4IMp5ic8fqkkoyQPb+kL9Eq/e7Ejxz6YuTagigMLIM
ubOmCHYT8Ins1W2rmnP07OTB48aVyQkWPfnkUQuyQ4PLLJYaKr9mIXRcKjs2CYrz
ChAjSgOrz8fdm5f9Sgp/WnSLbmtA+HQHOdJQ/eSARySuD6KKsTycNGGUV3D/zVwf
JPsyYO2a5L6jJ3y72qnGs4Ib8xBRcB8pyDnzp48BRNvqwi0yWj5M1BBapi5xfAyM
ugmJCVwhDyeNWeKgo5uXHGN4PYJo06oa+6SnBt9aSoVsXeWHRXksrWlWtmKJJ5f8
ID0JvM57lzomj9Forge9P1geDtiX36kE6rp21wlUrxcjgl4eYG/MjGNDD0uImx93
tGbxDt7xA6leIY318dntzHFdaUdnzBo0wd91vwNdEld0fhDbHcgvSUTZgz37+PGA
8svKofLxRKFgK0hJ13tbFxT5iBraoE5v7TzZ/KtWg6i+M1jEZHchOU+/GJvENCKV
jlTBwTK5YUzBy6miyR+EQ9voE5jOUkUlPelpgRiH2mNdVKkxIa7Ajkh3AMfJPJ0O
v0YQ++eaDDrTbRkwwi5G564G+xzaWMZz356ughRIifAoMtGldGlXeZjxzTLqRbkm
GA/6bSptoR9nVCj+/ToDVn+B0fhhJ0D02jCigxc+Voe+wQxDwGbu0ZK54a+vKkcO
olxHBBO93gWsqdlnw9a5DqqMCtlvFwOdrGnXuRylXLRBO60feA/FLIQZo6p894Ew
BN/f93zOVBaGmf7i2ZHUOm2YNJB+vUL/3Ui8KoxeNvh+2oEkvSAvlNnMZev/50OC
o6pvBf9tNRRwjFRN1zZ3x/xAhrABbrlSAXm8613CYuULIP7nRo7Yxc/cP7GZzhN8
42N6i8UBT9puxKQQc9ClepiIbkDeGOWtwU58tygeCMkquhqYq1zx5ROCYh76D7yS
k8pzpv/ukAOyEJepoNtfNp/x/GZsfNHkvD3b20BkkF6GZ3JJXM7zYlEqkH0eRYdZ
+cxxLmBixLYIEdiPGvjxqteVtlkJLTK7pCBi0zEnNGvRD6kdmTGrRX+4ic6Cu3e9
Igg7hV1sXOsu2SPHa+RX9eYibZgYd3DM68gArUBtp1wSRgG24GYODDZ3w7h5fmXU
1MCm/4OUAxmepngmkyDgJLonM2Qxdcwb6tt+s9PlqDmSv7Mrbl0i7/5xsReU6E9J
CUN1rg4HtGx55SgT9Fk2k8IzZlCy5AXCBD4iPRJtv0VjW15dX0pB/4WabXfqsvc4
qLFeZ3xkACpljdfhYq6TSa2dK2m2cwb6o7g8K7LyRbY+3OmA4NqwA9F91ySvQStf
XJdB5bh0sA69CALAlhkk88CLZ4Keh1mUMHYxfiXhO8+8NY2jIrJ1NEZv1ev3JQE/
ENWGYl0PDw4VsR4vswHDfRMNgMpGL5GhD3m2Of48yp+WRo9RYgWHPnfLL7w6tBw0
bajYaiBodTWgJvuQysegXh5koJ7cpU/jsT8NiavwXPeZQsuewTwehO5P/JpWfIJt
FV//wLulI7fsVF4RUmZipneF6xHu6FCZGoy9kwqC8TIwjdbbtjMsvID2BMBNJeZW
Vl7oVakfLAiAhCX55O7HnI4iqQUYimXTTnwHOqgFTPIu1afBOG1jAu0cIKxHv8cn
SXSGyhtbh6KbfOBaaoOtLajgBB6fJWQx5zoR5YUogG5VJQJOKSvffn0GaVFw3+ec
FpORvX5zDrCw5s6uSxuyQr4UQYt6VqldrUxZ/puKK4iJEGq0ap88siWcaWVSODe9
LAeV32Q9rZDiyb4qBz6feGv4ttP249qQB2ggPfHiYuSQ9fRa3A82p7wDbIiHYmb8
vBLecm6NDJp3TL7NnBgvBawfhlZHgqxuHuBlE+zYXWzFY2PE0aJB6AVgo+2xlqXu
kpuaaKUpyejzZjPr7RQHSa6QUyBOo8SdEDQEmKvlgm4CWkVBltPiViM+vv8ZDZ2x
jDtnNGPvD7kBg5f+SqX15AoLsx28LjZNFsENGT7EnTfYhtY37ZAMnbYuzUv5Jy9x
wgZ4MEksX1RqiZM1FktpMJz3DN4/PZPAN6qaQ9FthO8aXFoMCd31WagWMmrryzXE
oxKWYaEEDAm+O5BCOkQad9Nfac8bW/id4RGADe3DgnZO4LFC2SbWlHY4G5PPKoyq
e3793E3XF/kmQ5Vo3PTRQfd/msITzo8RrzmHD0KvYh7VCJPp2GPAjD1yNx5KCZn9
bIN1ULqs30wYbaYV+Dz2PsdDQtd9wu5z2nqSR0DGiKBqVrGAaNTAPyMwxl/n4OWH
TKl5HL8/2EChkZqA7Wc91Tb/TWXgs67KN62Ikj0BDlSZVpPAfDI7yoY54MNt15iv
SKZVuXIWppXwVed4S9H8pwnUTW5TkcVbu19wxqDrHBp6wS0u8BWjK9xA+UXRR1GZ
BGgeE9lrEquIB6WnKWL9ICsG0aqfgfIdOqyiCJfIPioj3jeizmLm/RALWqEbrGz7
YXLzCfNvM5nakwqaB+XyMVN2FKFaMnWt3JftN5O2x3RNS0baMkEgsHHhi30/xdro
KC6gXh+eFBnF7Z5yf+vFyZoTOkJkw0HSbKmB1QpfO04vY0rPtQh7p6H4ryo1dnRM
T6PHTZ3k/laAYTOSkw2cQhx8Jy8AlGvOtp4b8Ji/CXCQZJblQYgcKAfqd2SaIY4I
OETSCgggwgT0/THAudpmBhY96gQxzrhvYq3LOKbdoBOBa07QZdWw57pVUp5tOgKG
wR/GYEPbZKsZ2NRa0FsKkgADvUbHhBAYjDDrwebWNI2FMpAi4CJ5ezmzozKDJJFE
YkGevc2rbiS7fLdNkleFoRIYgyWW9EgfTEcU4KUUim8PowDY5PKN7wqKXFWEv6Zl
BrHOBqLDsdghSvXBnCpYXG88DtvQkdSHI/AGBaTnnYy8SekpLxYtH3ih6V1IMx5i
WZZ1y6P4MyholorXwlmAagKoPa5azYkPjjJ0hgHxAP1EsP/8u9qmOE2zR4/k2xA5
R5lANpvePpZEOVa8Ob1wLwphkNW/9E5w0gjgqewO4HiqoGXV5PjaMOVTpGMZ1YrJ
x2xFwrYosVwDwycDGpRkEybBy6E09oBdkTJlEWBI9PlzGPIqJgx6Jt0oji6yBBBK
zJj+ypnPE/zcTTHcymmfNwBU5GLs8K0LWui3JWsAybT1uFFdbNZzTd2S7BM5WWIT
COoupeK+zhRYUPQplvRCZxXN+zpPHz11fq9t4grs+5OpzRVqMsrxTZSmejsPjsI7
ufWHtKvyhX+MxkzCbLoQ+lSGpzBJ5cGZAHwWWoBJ1qMPdOiQ9rADWoKx879hO3I9
V8foMK3cMtKvO1CA6vORCIDg25/1izqZm5R8oWx4riGV/OC/p9D3ceMKpAiS6Ytx
vo27yK3N55x8pjEppJg2ssPMZ6TGt55GWNxdRlYVtbUvwZtKdwfCG/F9klz2OtCE
J6t+Y1j1lGhgymyQBavJudZ7Iuoe795zegl2d667042wMrJnUViUynDfppEgy4NA
+Cv6kftjK/zc4Ju5LrUHItuWLeGqc4UQ4NLcq+Lustqmmyj6NXf4TIPo8wj/pLET
OHPw4s4SyMLB5382XGxMDL2pR4gMhAdog/KwhUt0Xz5wZVU5jRaxHJMxL5wB1uDu
TUDl04t6KqKyx3PNIGaXPCC24bOtgx99/bNO3URU7RDBzBacDLzO9Q8OqREbZOjf
nmUpvTdx6zbDig6pwNhCkU42+iIIFUSQgsU61V4tAw3YmQBwtDGhYm51ZPndAQq0
4XBy1IVnUK4DhWitM5h9Rb0GqSfTiwCgzZpblsJQTyDGb9Yl2wWWi825zIPccg9d
8TVWQJtYj/ZkSRx2JGQfD84eNpl39o43uw/KGPx+x9rkWP+c0fKd6o7tmG1hGYhr
CBDPWgQ6ph3EQwnb2/9BdSIt5OpN89z2q6TxCVl15GLqggviZqqDg+9byolkeish
jsEL/EF+AaHOPXwfqYYup8CnIVqJiaNoI4VhsFhKX7p0UYM0PSeqhUPjgK4/ZYF/
sOK+cDOoalvrLWD8VKI1cSXBI6zdlBzKpXuHJiSTSc5UAcFbj58sGrJhxMiY5Xo6
L505YqLLdZOsrufW/ygn2jxH+P/GMt/onJQTeSLLj1u8F3Y0xDm7jBlqBrL7Gwmi
WgroJdugewAGy2zrN2fGFbmi99Tp23N5M/wYo+dfA5Vh06XUu7cKgZkNUoB9w5Fs
t0fmXSRG8LnyWMVqwBgeCFQ3cI4X+0ObA1i22f7B6/s5fTEMEqrs+XXX0d0+xHsF
rAdPdTJhoB+HRRfLo206ndxmboaS0xIJXnhbhF0nLxI0jPPdHlavI7EwAYI4AHPT
BqjpRnVQAS8qPXqZxnM5FJRxF0gNEQUs7olH1bKi2Vegy3wtQImsVsRJIg6JE98J
tgz+LQ+QaX4QSUy73lsUoQfgVy+p+6C0kwmMiet9+P+u/zyE8mhT1zfthC/fEARF
zUWPq7yXnTa6kP8ChJY+1Fppt7ytE/CZozXSMXjk3XnuauZ5zjpOR5ry0AMhqAEU
JASzjcEjTmO5zotr8hlvGjaXU80sEW0Nv7pPIkvUy32wTd2Bh1Zd+WruUZkTOC8e
97KSVD6PfLkor9ZicCR/zoDf+P55XdvmSwNeNamfOIup0NEyiIPVNMYLSd3m86bY
M7OJLF155QArNroZT55GhxxXpiLLBkqncD1y5M7aMb9kRxE64uxDn0I8CmG2U6Ib
2bp7QsoLVr+UI7A+T18ZOGHTGUFnpZeVh7FRQ9n7rHKHxIF521CPjLRfqV1dDTWb
IU7zlF/JgZ2690of1hAqSUhtgjN+0av52Ev4BVRv2me2M6vVxpVnfInmP82sLb/X
7Hcm1ls1yKGHd554FBoLm/Pb/vvKseGBwf4JFXOfsrOsnNP2zzFyOB+REXnVxHR2
aZCiTqlyDYfwfSviQ38JmFB2D+I0Plvh4s2Uf5BshowjhNg2b1Vtl1eMlivbjp2Q
rxc6Vzu+igtFXPotqMWPPP6V9u+S+L4zl6ESu/5GMLq+o/4MdcEeA3q4pU1q8Rfj
7z7iFJym5wJwLwvU6YPee4SVe5YEqKUF1Gk6yic+PAw+O1q9T0NMPFVsLAFbE9+U
1c0gwp0yw58XgqNaJVNMPqUunPanYOifDKtJm9OWqKIUPVbv5rVA4Q7zpX4gdBwU
bE/L2Aa4qWz36vjN3ZT1Yfe+ZNMzgaixhAEAcI/VSMOMdlWqGLyhKJzXsvupr3eY
93Pr256d08jj874iAuVukx7Zj0CHhdfHy4CVtpirkv+8IC6SRpE71qTKyOqc1hDP
JETC9QCY/mEelCrnTeVcDdvQcA+cDj5UrWq0zRZ8Dc/k8Rr9tAjMBPbvTvp2bpiI
yRtE2BEXiK2qlUxgTDBgahne1fJeVpZtEy8lhurjdhxRlUGc3UUCm7U0LrJdfhRt
Vsg0wSNEVDv93ypcW0I0H1YpXME9kw4jyzNqjahWUVea4EBFTAOm0Qr4d4KIPMhY
XAqpAj7UJ1cUlor10bS0dx+tg4QZY7q9XYfmX5njJVL3gCSzhmc8brt+HqU5A6ic
EO1h32boKcv01kt9W3V6MV4NS5UA2MTfUxbHybEdkVZnCg9sDAF94v+2eTKAc+FY
fDGUXi1C0+AM6QTIoGr6p1IcRPisONV1b8QmLX3D/SPgaeS9PL9mWfXGYxyCaeUH
n/AefStsz1IlFNSWt7r6zraf3FSFUsU2al2V5f39OPYeGg8JxLV5fmwzTQDU+dzm
LSrZJS0ynIsqVPi3O1GvifrHBJKZ5FWLSKd1wWURBSHqAZCFKKTKOOysNcMhbjjU
SYchX/NnWQBZRtr0njNakRUDE9kP1vwiPgTDJvZWO3n8qlxRLwhHx+dFXHP0r3Yq
gUs1bGaIVXzAJGhJsfh670065gAKbir4WYbnn+SvRboqSfKSL4SJkqGQP4Q/kfNC
XXZWmWy6ublogbwOGTXLnLhuJpe9m3cc6tYh8Eji2+G8IwFBh7y+U4d194JLLQdt
EykyMJ7kZ72jXE5zYiXyNBNSnuLOQjlOzgQnD/DLTUBGFEf4avhDgxZAsQIJKI7k
moNw0qx06DBTlID5hY7K2LJ7BN2kDHz40IFtt7I3UufDUlCEnGT2we7o4GwY2Mhh
GKPwPrDMMCbMJYv7UracUi400OIhd13j01SIxfnX2mAguZkuiuM2mWSXcfd2sDih
rLDPzKLRNBC2CqXllJKzQ3s0/gDO5WtLfkmDlGfgles9FUC+5joBgF1o/kFrO/CB
VFw+oco4ZSfNrnidEEUuTfPUXhi89sh6bULIIGiC02kpTICZE7mzue2SLGGvCw03
TETkdORImXBcWGrTCaqP8HzmwPpOy7XXptFGiYHf+MqvCDqFh7R8p0qd8m8xVU3c
/j2BdwPhWlesLGv4lPsRuBmRQw0hAkFsv/n5zn9tCLRDERe10500bFGBJ8nlP70H
DklWntnpmm1iZsU9VBahBgGik+WIf8UlVuZD3xk/Ncl+gcXPIQGxoMGsFWL3OINP
03iFZRYePpFs7tkgy7HXGIdRPTyvlGcQC2Zy29B4hCyXa7VP1b5ku0HHMoQ8JHEm
fsGfUYv9FhyXv+YHfLu9NMvKQTb664FVWsMBbZI4UwN/V/zo61bG19LruFauQQPe
1v4s4bXiYRf7mBLxb9OV2TLihD73iesHcjYBpgGae3qBAgtA09Wj6V6D81XF/JCE
ARCgBP+6mZr7A1CI4Lqr/6Ek7pnw+YnRam0Iv5CeinqX0GrQknq0e9+jeicKQss/
m9nIUdvRu+k2rzu+bj7rOM9+zaChCg4gOSkO+TrEry1RE/C4veP1udcymr0/jOey
ItxnhWMLh47zcFQIHp+VBHr4eflBiy3jkFE2DvSSamOtqWqbqY2soStW7e6rXMNh
n79ON55hBK17961O0Q7RkjUq7R+sWl4bDjO6sfFJh0kbLPrOzlolXpAhpOCWW9Yq
BnJ9rhOPTZil8Q6RjIWRQIU3ZApKdwAIgSLlyBidUJ3InuvwcIBneuxI53BKZh5T
EjO/z4hP4Eu3pwzDqIr3WY593tXM7ixlzZcWcaOIAWiAuSzPqBdFS0htzRWoDhr9
CXZOD1K4mnG3ptt1zba8gociFqQzTWUFRdzCL3Q50lLQFIyi1512Ke8qGaHiiZP2
S+pp2prhpiBPUo8NTpKzaXsNhNlTKT2xOBuy+GNHjHbPPGTsxVKPTUinBO61Spmy
ghKnkWGaZkvzNTSUDDCM4SAM+Ln+B370UaD4Lo4zLFz+47AXpa0/AVbqER/S6+v1
9irDtiQYXjWoX+UcdwQsi7bfYhizInLVOWcTYJu4bHtgS1WGIY1pI6386HnNVCAZ
KMaFZ6oPU8zGQxbkpXc2cJAk3AdplO0mWV5ElwZ6mt7b/+nooUN7KYfEDF55npdG
0tUKJGAUnK2AStaiJb1UeZlrmjVe2OMbhf4hZ1bUCsW/J/+rIba95RGtjVcroofW
mOInXTT+wadhgOovzJsNm2KPP4u9BYyo5cXJkU13/WnMQJvZ+n2EBDuCOWBeG0vQ
+b2vorsV/tSnRwOMEEEueQfr3yB5z82EFhyqo3viEg0C7mvqTji9Kdd3SWxJJB2/
KBJcb22FNyAtD+HbyVOoLqoXgTDVfxxosudD2vSxhfWHwM81YCcuhQ6qk8DSYJ2d
o+xaVrlQuTJ54HZTMWxGf0lUqDNrR62rgvvtIoVIac7To6sA0lDDLfrWwSd6LJus
LyNpGyB/F5TvJyEK4eCH0zsiFqFWBY/0iocQND6h7IOwzzzRx5yWkWZtlSTJjMVn
dCbbMFdlkR055o13aTLU45pzBQCIYKqLvt7F0CMMowBd61PZqe1NY/ipLlXUmII2
Z8KY4u4fp0pe/rWV6KVmU+DBfVmF8aRV7CwxjL1tz37oUqHOct0BrNj9raAot3kd
23Dq55Ym5P9iDDemoCox4o/gPDNMmtW07jYWL3MR6EVtWvxbLwr0elUTijfvfwX6
2vJNPzkK/8sUXysOHQT/Y5dN2s3Vv4lp3ZsFWLP1NjqfVpjk9zTFSfu/8D7RsKw3
sLGaI2DLm3kIQt2kjX2JyD57xFS8mb/sT0AWjfkjW5GXNYyn2dy5hHaEDJDCZghH
eGNoI2CEOaH5Sabmk8zwsd3hBnZLrsefYNOmICoSO69Mmph3TG07eenKsYb7L4XX
l3Cv8+6iNb+6vpDdBRod6Ksln0JEFsHszDPAhyIZmxfs3kXzu1i5VO3JmbVThcjX
I1GbcgkPp+kFWP+OI9iqqADmoVh5PfIbBV6tBDfvMKjJuffm9rQHEHD28QbPcMDX
TFx23VUwnvNB8mWTHU0rAkcuJpc+ydH3ATEQK9bTdWekR71aBssLt4kVF28G2JMu
PxxGp0TtjDxkeCwJXAK2lZqMZj57rYfJ9DWC+9KJ2JWvcb+GT7d45vCu6BT7GPt9
0uJCf6lHXDhETDSsAASpc1oTRJinHSz+UUAPt6ejL2mO+4r72jMdvB/8po0y3cqt
lpa6dQ5srphPG57K5qVj804YrbKITmakSLbaVXL1USaDJOaO/hE9liCW5dEV7oRE
Fu9NQ8L7NTGXUrD+EMGZoIZ6ZFAE2FhtAOUAqt/4/t2d3Gjxd62FmblmN37YX2Yp
VmeYhtYIIh8dYFhbzlezihEcEYP4tv3Tt0hGgSKVnPmIHC8lYzDu4AaV3adjJYwR
6p3K6BCu2pHEYY3lHodA8PfvH89K8P5h3h3thh+1awTbJ9WBhCm02IcJ1OtLly7y
nZjP59bMoAD7o9l+rI9+eMFIh5qyvEKQlI4UCwPu7D/zYuzjo8hXRXcL/BINInni
ItDPjFObth3+LMwVFGHP8B5cBYuCCnVdr+y3doZ27+TIU8FaK3+VNLrRl3Zqvow3
xRRzP1ZNWP1RdOP0MHEtbOI/3A3Z2MGwvh4XC2lq5JX54Hg+pvFEXXSNaMHZhlqZ
2Hs1wPeBpYXOw3UWvvENSD27TvbGUduXCJoFNSmYg3prbU+NhDxnfy7cvXBSDhIl
QTVV2E1KmKQ9kYduMkcqarlTnxd/ifhyAeCr/xzlMQeoDPLw8alcfyn1z2FkbCtz
9hhZgmf8qT5IqAXFWgkIAmTC/UKWiR/QLbW95cOylJBO4I5XxDy5omsfsQYVhp/w
9Bkp2xteiBJ22YGyhjJWlvjfUbrBy+GQrDAsueNTM6kqIWdAmhBgPZEGD8puweyA
bg8TJQcSKI2Vs7/3tGhFbkIp3xx0HywJZS3IyxQAhGFdOnxF9lTVePmm136RLU8/
15GT+36JSYD3Qd7Ejr4e/qYHHnfMUdRmN2idKtPVx80xnQgZGnhCwINNDsitDqJE
y5IgOu9fmEsLih9z28NpNdCpfFyt3QG5oHycQnX6hjC5PU5Qk6kgnauB1P/sQ2mf
rAg6fwhVevWevrXvGVavszw2ZqvVKDl1RzkU+z47uIz0GR0mUSwKPo9S4vFCWrbS
xC0yoDCzBee9+bIxEYh4KkhaNDDtIlKqOyX3/RSNze+jDXflCelBlVJk48xcBnQ3
nB5dzut9BNthlzhnFVXbZYIAHCTHaDEufeemDPGQ2kBn8TeFcxZs3yuihXlnErDI
Pz64zfxCS+1VXE76cWkuBCcOniS2YQAme5Oytrz5fFZaTcW28zIRMvX+/uQr25eH
w9Tre0lrN0bNhUeR5oSwQAd64HD0O3tNH+2fdvmh7iu5dngKWJ7w+bviwWfAaNdo
iY5umSYw/6zJIIxt8ib2O4c57Opl/0KGAG1qK24uyIiGsAyuHMNMOWTnnjlu4APr
W3G/QxBMuFz9cmhi5C5GRXPyNR8boZwQfpUodR+7bffixa25csgUVdRciOi7VrV4
lR1GJEQL+2t8ZdKl3hqvvqQzvWenkjaF5BJ4kLxZotGnGdg16ejqdB9DrFlQDyGA
lA1qb/wxhAn43G3ez3qCh43eZJP04Uyivm1dOERyD/p3H+d1NNXYV9Zr1fFYhILe
4vjnSRQLQN7aXlOeQHBMg17MmXquV6yDjZpU2+RIwUNHAq/plE3Z9KTQbt+zDers
M0koLINsYuIy//h0zLzDts9VnDUeo2dchPbISTaRT1kj8l0U48N6XBCRZDNLBglX
cflI7x39/P5S37or/k1qsxi2nUp13Cr3D+iqJZUuKPmyz8d2qVTD73yYOiJMmIpj
4WbspgK1KO2pwcGzGhzN2Rn0G9iF0ySSn81kMCZCp0bw2ID7U9aynGlp/LPP1nqT
rwszQfJ/l6X+g1u4EiQtt5zeREGzuhf0BuhgkS7Znsou4eNBO8ApzDCSH2A4HUsE
mNG/PR4sOV+ac0l1ugX3NKunB+ndrqveFUWhxhGRSvAeSVaGBsF7f82QUdiizETR
HJpoJpX3nS5BJHZ2bNaVrMeDYhd3oyqWf8i22KaD5Y06GEmUqxtNYy0iNOLJh2kd
js4OHwEtcfaIR/N2rI/vxR23HuSCjz3asgnVA05xR7Y+g+fXVLxMS2WqultIRXYR
JNY9JRcEOaq2SR6AC4D2KZVsCarE40CdEJMLnUSVLYsbB9zEOM2juYV0HpmB6qp9
4ieNSGe+BrqW2muPL3FlpXzSkiI+WOC+zzXF6I0g7vbgGC4kP21Ih31K3zcIEVb6
rmblmSSsu7ifOlCz7QLr88nNfJTHjdRuUB0wrWHltl/yVUWMO+TMYs+fKRY8AVVb
Hu8wOlUbg0cAHYWcuLNaUssV0N/hN2T97WPhxnkOEZ/2HIn1mDaovn8cGOmPY+Nv
Aj0k+R35VQ8ja4jseyXA20BhLhDtRLgt1awcczmGcGqNOiXZpigI4dFu/pq5Y5DJ
bnj5tsLrTtkejY1ODUVFpRqvkaEdOHyl5FAvlhd0yuZgoZSmRfhiB27e514+9FPG
l/2skwTehHbJCZ+49lmrvp3f/uEVzejv0mOv89SXH6X1xipjDryTtX6Ad5NE6/uP
cKsu6nwKcuuDB4pOSD7qdXVidZkfu3uVDn3wZoAOE2EGJQ9lzS4psxOWGjWicSNo
Wp0IDZmrx6uae6RsVvt3oKNsk8e2X9L/H9fXxZIbe8jDr2WPJDhs7CH2HOS/e0lF
T49fKQLi/YY5lNZ/wHBS0ZRoaoJn72ep5rCuGMfvoqbqbbIWXK3eyGyVbjz9Fc5z
aZMAatHYA/kbZSHsogd8PJkEekdfkW3YDVQhoTHH5zjOmpsFNtdMyvHqueLYyM01
zHomifrEq7BzBtpTRgmRUXhLaCCAhAJIYIxviLhYGQIQlyc1IdeelHjpk3WxfkgD
5Ydyw4g/zj9pVVwgBQ7gf2TMRjaT46mVczVE01KubJIIs42kc71fATyYUif5B3ek
F2moRwbL9gvXf6IjQCNpGdbwwHhcnO72HcSaW/pTQHQctYeNhKMdO8ZgkNLznlGW
fJmzIp9AWN1USIrnH3cXlxMhc324ANQ3riheiabx8BYKOT1KtCoEUPqpDMC3dVI2
Pd2s2A5VWojluGWNQQcS+QOh/MrszsmrlWg2gHFeRAmJjjS0+ZF/t3gAAo73SvV4
UqP0FgpYprRcejfEoijvT7eer9n38ChagcciM2et6LBo5LVr1p+RyD07YjLvUoQP
YjSH6DjM0v26pDpPONK+3+krEM+VukivoEtmnzOEKIkouFQPmdf3jMBvrK5Dvnd3
+ytyqHrHPELLzQ7IS4jnNUtUxUx2FEZ0Zi9eckKXBmIZJBpJeLjzf+oYLhr5I3Hz
URUDXuzuhwcMPZT/24/Jfdi5VlVqNH9TJLiyzjizS/EqSLbLExU7qzEO0PtEdXEb
imVGTWPQLh6i/q+7/9RYryBT1Y0/w80We/9dBcl96O3D9in/sxixVN3vaIvKSaFC
5zFIA0jG2NNt4AT9ttgDjw3MyzyxRSs3xy2+J0T5qfIxaMSmycfl7mqPbm4R1PNG
bMz7Zh9dfIfgrl9YO7AswN5zMfxR7gNWdWyuexVdGUU+ldEik3j0qtqpA+RycTMD
IpJwWZsivtBZgy/ftvyCoKd2G4LGtXc/k56dsReb8OUCdfwPgVS64Sl63J1dHht7
ZGTZ5DrgZd3hPNHociqZRDjQQSjmbw8Eyssd6ifRrC2T7I+rmmQaqVRG7tHsxrsU
/1+O1+CEvc/QdC5TwcjqjD1kjjx1qSxxINuur5Ztj2RQOGjLAtUcQxqFIfde0z9C
BrlSa2u8qdwRU6meFLBAIDoXjeLpqt7FeRssdftYG+mwhQYT1eruapfrgqUlw7Wn
W6ILAcAvOZcy4x51396D+WQzFHmLBgT/iFDADIercAPrlhHz8ViVP8M++21ffVGb
w8hbcxoN33Aa3uqOkahS7kdQm6OVi3aWePfNioe2pzd2zFgoYSIMPIRRC6tsYrZe
RCQJ9SWRDUa9h8Njy3Z1PzoTSp7yYOiay8P0q8DEdCZNdK9Ys8cJnRGiQQaF7L+7
wp2uzScl09NHnAS2rAFIPVE3l7bW9xikRTfVrV4PaS68zA8eOMl33Ep/LBv2uX4y
rkVJOyiURv6ZJ9aOF+cW5/a7B3/0hjjrrTZ756ujEeMxFw6tKKSEFTLKFjuGrnBL
lRBjVGI8Ha1JARy6b7HOB9gVy5jXLxcApfIYgeTJeFl9Ot0Ot5lElmpfNZHEj4Xq
H5yqH91/bt5tducdQt2n+G10ZaGVcdDMSiZv9PXSYts4cvZXNNU0phhX0Wn9IYAE
S/zaRaNvPW7L2puKH5P6G1gFUrOz8x8OOi3wLGzDtz/skNkRN2gSscxWtmVS136H
/cuOVWqGFXMqXTEo6F794Q2bWHGPx378FNkz0pzbn1+MH88PewXzZUBbGsKPJBdN
Ka81MbGH4Br2Vpfzpi/uM6aepkS5HSyLQTD5NYElFS15Aud0sbax8vLCW7FwqYXk
P6NeFxE6HK6JciFZVRuCAZ5ytgquoZxoeqS5XiU38UYKqCFYlKzU4kGD5t7//NFq
SqLh3BLQGAPz9EqL2rTZI1/DCAVXTdF/S2Gom9LthfXDIfA+0z3RLjTlvkasWDoj
ZtDj5NnSRMmLSMK52QD+SEjtnyFbwFM5VmCF8eLRUOsOoRQkNVm3Tr7LP3fphphe
JklA1K6U/+Munxp/Bl1ODXTDTywc0oUMIRcX6pdl9QC9b9MloRjS1NGd2WObkgwj
dX9WK3uipEYVG1giOa8NAZgDnsQ0fZkGINgGi2qCjAO/HZXlmCO4Y1ORL4vmmdkV
XVuRdD01nb7s3Tr/vuZDHoAknNHRUJl6K9/JsVWaD18tU0FZFP0cWqZ57RfyXi76
Sbpk9zQCCOoIQD1sMTr9ht6v6ey6jd3m9N+QbGXa6rOyn7KKErgSgEUhzshOYXA/
s1+ko5QB2UlXehqmq1GCL8BRcyzLwHkkPH9aNBzhHo19JJwBj6yecdupxeadIpor
Vy1t/GQXyzaRMW3Kd+k+lOCPv1Q9I74ZzK7hg4dQinIDjsKazMVi+GmPcUAoOAKM
RpDeoSLpVBmQTFpVp5Gy0x+OqZFRcMt9B/pORg/KZqHOxYBjecD2OPbdt+tXPq2w
4EMFrkNF0rj4DX+m/OUuLOkvu85toObW+aIEoO5kpQpc5N9CHrWHwg3lJt1bcBJo
mRkyWx9gyQbYNxVXMr+kGlPO29OZ8ra/DnP+lkx1w0jM8kQdkoLWW2cr61cBa2Sm
uMh5GbXkB8LLjnJS9SCpCK/UxcOzbQHYmb8NviUeAEkj3r4PpffeqCBfaMrZI/x5
X9LcFxIg0i+5f0s8d7UGAdW7gd7+92rYtHXAzByErTDAgeLO9YybJ4Jmg8n3rs/F
VBz0W08wcvJ/t63jDaTIBo0/woC4BEHDQYRIBveOFVaBYILIZEeQ9P5IcrvoRb1N
zRC6NR822dvKoAkIGNzprA5ZolHcWUu47+ucIEOyITXTaH/j0Yxk3DtiRxpBBv9H
QHVtndJbwA81WoUhdrWGjKcTREYFZksF7HlJtl1EZ8PPyW3Yp9TRP+CUS1qn+A8s
X4O7At9jwqpRUe/VNbUgt/ZoboGXwxA7k4yDIQ6QQfnVKSWaQ1CKsiM4uwEYpXdX
34Q6VWKdxvejuG34VdrUULICO7YsNPB63kDb/sx1nI36lEkyskTrA4vrYkAuKJ3Q
fMbM4ltbZj5mTLEtOcqNM907ZmU3SNx7IUYp+QpVMArM8fA+Q9u3VCOs/Avsp/L+
KQoy+WzDy6P/llilmcesSFyJNkV5pbsVLvPTcBGdk216MGBbMFarh476DJk65KG1
4q9yVrUn69tZYrJiJT0KOnxd+IgyUPzwO6dw4tnPUmTelMdiUKjHzumXXSi/UCUx
emcr4t0tCrNX+1B/xXYoQbckEWhNn4xkuTnXSDjOXGzJo0hU/BArZ9tlXSrXvwS5
9+v9d35KDrbEAuCp2+ri3dL8UKrBbIb7t5HaLY4wb0/BSFm2u6xBd/2L/f2/NRTH
wIxZTJHwzAjHQLBTVJoHPjq2vXT/QAJU5qJXeCXMip6Pn0wuGbwDSKD4mGot62di
81XROz/H9o+EDQi0EYHvWfud1bebNa5CfZCusIrsFLski9QeShIKsUwdmKURfbIQ
3gHyCw7VvdCQhF+Zhz1nMOcZkINzbpW3S1QhjnztJeLiEl/uTk/haX4pSeviP281
soKeYYao8m0oRS3wNJpUbD11jBrWsoo0/L9S80Kr6knTm/cuWM0SC2xG/ifR9cb8
BTrZiT5cuBCObXNiHxrlPWSrTqAWxen0qCq2/FSN6o2Fy2NC7SunjMVLfe4auaWS
lXAZ5EzUJGvgN3dx06+kfDLPgmO/4kJk6A3VdbAOcRR2ASOmEm/ge2tiiVuzLvdF
wYuPDI4wcMdgnSz396ElNSylXaACxVKrjthy0K381RLqRU7FK1bcbLMbJ3CV6MOR
Ia20yBHy3pOH54unGoz6rgocym5FIidcmFrq3lOmJ/UxXLIp+3dozbA143QkOplD
wlUfksvgJ4tQOv+HNM9ivqjnNOvdTc8Ln8GCuhwRVT7Dq1pgR1HHJdONm3T4Fc+R
A4pId2ySFribQ74eYZbrEd7XTB5TRTEkVFLPRbkvAD0uexcLGnrWsU7zm5p4e5zD
tZOlDWMXP5uOAefd17Au7YfkOomufsQDU3KY1/CDeBCs2SujF97iQD+q1Lcv6Cbc
WFlMVsPlk0+cc5OyqS38qlsmrQdKaMGPaL7l7wjnGmTZfQCrc156RDnHegxP3BDY
Ui46OzIu6TiIVCwpIOZEDGfOCrGEP/QDhQjlO5xzIgivuWxafqjENHTJW3jHm/xS
2n4bcku2CXbJtq71Z7gjHVeIhz75SnVJqtagkHV7kv2I3O9XK1WNMkuYp+UMPi0R
/kWdAUsPcY6AS8dLZLKJ0n6fN/ICNos5FtctV1rJeje5yPc1mSf16Gogg6Za6Heq
+uOzvpnVvR8gmyRCGyG6jICyDpmtDXjwhyROzLyQzYThhdbV/cPNZmWWK0acAiZO
goRkurrFDTidkyMl1+HWNVZ6bRHt9WLz74B4cl2J0DJEPq+1BOe4Wkz5RngouLT6
oefCUc9iOnMNsy3QrBLvi09IixfoagaKLe+JmOEo+x8zQtWlm38X3MSgWEmLDkIJ
E5tOAnsCXrCQMEIwMaKNdmcNSQTt9+X4lf+0CVQejBOdU1Pl3/Csyhx4LiIzzvTo
rYsrnaLNP8iltiIxFsdDZnvSvtn1ZRJb3HNPM2hcB8yNIf3IOvY6bLBnHdGVazBi
zepTm4Io+aUjqNb9r+ausLqvBci1EEXvMcpiBTGu+mrCYSX/yUX/hMzky9Frsu8F
soBU1qe7JrkSE9EpmhxiVMmezv356qSa83QkCIaiw6tCqkk1LeYJS6RfdGvNB4BR
3ArNdF5bMi8BgIh8yOkgQd/70VLH7YiUGFjYKRpt8tJiz0Y1Y90PgEt3FSdlIzML
mCW0rWU4EJPuMvU4fUkwQwbdY5IZSgY4SOaIKaBRQj6KM3EQNq93UxrZ26A4znjG
30aw1ORC/Zbs3EeJrTTXePXLmGGU8vi9+LNm3n00eWTTxhvRV1E67/gPoEFcWrQG
UMF0rLrdOxoKOKVjPqIO5AkfVgF9Zw6raeUhmexcFFta1b30lE3J5EUwffukn5gq
VX3RGNPgagSaxg8RecjGkeC9QUrYTdEhXCHNPYIzlsxkj8bubkDIy2NKx/n7HYrC
CxcA39iBNzGHjMVPBgJI/qWqgL5oO1kkF6XlMycBjVwGNCZLr1TEWzxY6ijp3YCN
keAEG/ZPgW+HfVQMTiVhJcbGKf9/h1jDDmf1hQRzzObZF+Og0jryB6TjgRA5ZsnC
DpZqR8W31cAFUc9MTsJjbZQIwH38zBXPetFLGju6O5E/IvQ9ziZ4W53oLX5ceQyR
jfLYR4SGpmqb1D0cfxPgYh86zu9fEl3f6wMBKWDWuV82xyYFbwuTQF5av26z4D0U
zpND8tSKQ7+d3KGCLAq7Z4AXjF1ojj5XvHsA+L11NLIX/c0ksNHwSF4QMNYmyDwk
+vyCkaM0XPu8OJBF5Fjj1GY2qfVuzriI3e/4+2W416DnwhIBMezy0H/giI97FXiU
d51VVOi4xje7TBQT+2woW5tBxEMvwTIYWNu033H5HtAdSaenMCduixyZc7OdL2fm
GgEhrXCRfdxZfbvty8TA15l+dTB8+P/XPe9vj7G4s0HIP9WxGBavnLzu10TABKnb
+3wEbiHUG5T62gskiI/FadEQSbMTNyIzLocq3kPBQsf+Yh1WIOQOmmAgRXXdZ9I/
A0OZCmHWLruK6uKQBZbd6NHRmTLhXN3BabX5u99NEjGhON5OUGM1Bkuymip5nI5i
8W/MbjkVgtw2cv/4XT9xPguNBqCO5FRMnrVpjJgWI+Ff74WNcnFu/kAPQszrPyrC
cGX/8scaoNlTfOZ1Y/W80Kz2tLfg2/nRYPdr/xobsV7tyAjNGn0uP22ZE803LZiv
PWC2M124j4cxElghO0/vMxENkP/6KDbKrKzz8z3IT/UUnl+/GI8XMiYQVgasxihU
HpSWQWaVLvflSPcH3yzEVv/OCQ2CUlTaujv3Wz0UIz88ARzwe6Sapm+85vWWNZ28
rUzTNlA0sYRx77pzjbVwTaeLJhcJySz/bjRrEQ0O6EdXNX7BLTILbbO8lWwRNkNC
fuhew6iQ1YgpH4uKL+XjwwGtchI4PKmTsEnu9HiV1MDanZyIyW1Aljx/8g0oKFnv
Sa9LdOMphaRMoJgc7/PkH6G8FEMoynBFuDM5OgQyANGv5ZL1k0wXu9EMUti1FBWt
ACThoJeBVFAkVQshraajqGfXJtjVsMrAGW4//7cAKsz/nm+l1aZBl0Thp1O6/0Kp
UYKoombbV5e0J9XI+1aTcLOPnxictgfqDi46u9U/6fVGizDGgkrzKa6gyGSjkY/Y
fjSVSuV4Z1XLg2zsvXEoW1kpLP/7RJMuDkhlZ1cd0TbPxWVOackPig9G4l3kaNck
RYnHeiysB0kOvSI2Jo0WZxDt9m61bAqaJvywWpCMaCmSAniWH2QCYSuu8OqaKl3F
S19aUbKQgn8AghJcRWrzEyW62fvr/ZX/6PJBEBTo25f4mNyrzTWW7JWsoYhl4Bbq
V8CLPsnCt3e3ONACX7QZV+0wwTTLh4LYY6ufzp8vNqn0AHHdaE3NbdgD+y66+iMY
HvIb+msRABF21ESu+TRq54XrjE6vFCStf+3I03DqkY4tKwa2UMzFF1n8q2NSqJ4b
n3fWbjbZMpB4rextkvk58Oocd4dBX0cM78Q6ZI54X3v1Q0hw6GfwEy3EEuijRvR7
jxLZe/YYwAmpKFVEerv2K43e7opAz4NvGkV8qyLO9Xj+E5sTNpH1UkleC9av1j9e
E7hI6Mhe5Ydqsgq4waWeapSiayI4/j/F2I/bqgeHXlfTvWI/Xqek+O7Zoy5MYAD3
YJ+F7QngCyKCv6N+F1nlbzqojovVGQpie5uSdiePMWKmExe109f9T1kWsLadIM6e
DT6++YoPsziyzew3332f4KK5hWQYe2XSqXFw4n7SYJbKaoUhtjD3awqVjWDLp+yF
/eixPV0/tjS+GQQ3g154qHT+9zbfLTmpBtcbAeIiv4UG3Rq6mXlsuR70Ce1KFJh+
fElqdF6KVdZGtfq6FxEYIwW5351fxr9jwkYb7Ia5bD48f8N2OubDgJKI16Wm8aEG
MDQKez4dk5pizR2ZEoXHpu82Kbj8WHJH6/iqf0BI/6nUTQZ5g779S2ahu68RpqtM
vIyxOe8+igx5cZH/heWnA69oDtuLLq+Yj+UHzL/vgMqyotf0auJ7p4UpQUlapH2p
BRZiU905hrRX0s9QuEdBh7gaiN9zZi8TqqYb+viUq5V1BphJqXGyKD4IdJYyL72W
pIEbrIXn2IbAMbRYMuPphDdeYGhSuv1+zNLbctU54ffGFizBM4c49ntzq+I4PeWE
XAwRUrf2DcFZ1dY5pEUTfxMvMj6ylGpoRnsqbGAss/UcPekVPFloof/u4GMEVDL9
exuB9vRyol/Yg2IwUq16vRwYIxJGfbv0WYYNrCkk4BFBmVRX1B3gQm6GtwA99ICg
DAY8ngvplnsquAizA7JpwiXfYsDe+DKr8EjxwFLgCtC16uRVSvmD44ERyldOa8++
Horyg7CWaV5Psnh2WAVL2vhw8aURKWBtglnrGDoXyCmFdT0CDL24G1l4e1l861hF
qx2dfGDu/4xTFKhuYGW1jNQImstcgNvZmwFOQEBxLxquqXag0mYm8tzT1LtFTVQT
a/+nUMrXrMYq/JB7LGQGB6mmL1CZLPDY3JmeHi3BALjPNDZm55QnwCpHjddy8Xjv
Vqc26y+z21b5HFCf8lGIjCXm+6aKuYBuKMBOVh0tcXyiSsDzITg7NP1LrLzBrOP9
xadNzpEH9GqTosIdcvmIPXPK3RsoZs7Ct8fBCVOOF9lccuHuHhWo8OCeDWsQjues
KgHLpwy26dmpXS/fwFQjtWwC+FqXeiJuYa50fnEWewrwU1Lf0LfUT8Ld//zzvAM7
tuHTobm3YzErzQ7U2F2QOyYi45lvdPKUiSMf5Y30prhLQWxXcHUtvIbrTtXIIRs1
1HYwW7Oeqn02gB14etPhclOln5x6h6fM0wYNgvljo0Qd4Irnf+ida2JdsWrX11Ss
WUUkcfvG5EaKVrJF02tjLpaMZznZKrgQzp5D2+4nY67IQ/cmz+hbbERaBe6HppwU
hMSZ4vzW8TgL2KhTd32k6amz2R8Y1o0BUfVGYayD3v6Zxryg0yjGrrF8woU7vRt/
EfYJGxRE7n3IePvwKsPSjvvMu80mYYfin7E34KSCD4DsGRiPcSyCl4+iO78gNDIZ
SoBOhkaTpkN45K4VZYPBwHsx/07YiXmN57fQsTsEddUlavgvJGWaNmd6ER5jJiNa
FkPv6pBzGbuwEeuVuAZhx0HtnutPhBiJYNVLIhihMdKJHr3b+aJxpRbpOEY1qjVd
Y+hr+qu8JFFO0Y3+pWrjYsIHjtn0VuNiTch7vF43z/eBhv4fDEujDFrE/Dqw1223
THa5NlZ7ePzxf0lT/EPLiZiJKrsVsPhSrnmxE0YLRYeQuw9zMk0CnWq0XKnU9NH5
RaYw60nqhRtiOX6wQTaCN4X7yaetx5XjR7J2hBElr+W4TAGXGbc3N4nWuoy2tZ+0
A3mwI+dTE5iF/QdX6wnw39v3YkalSHAwEIWZNFaaIHcFsv7K+YIRAbSFxRJdM7Dn
gRLUM/aNktNEDDAvkHoCimPPyL+PNmVxxhK9FhDFTtVNHPKU/d62rXlPxcHqMYBD
LzpeSRZMKMqRiXUdGrpjj+xdTOuJFlo3u7KdvNGinc1XW89y3OrAgvoBrUcfKU1g
qKI2c5DErOwcS0nYRPTyhq1bzLkvgY9kdRyVz1ELy6siUPep78CI+OhM1Tz1hQNA
wD/YO+/ip5A81Qu1OhT6ULhlq2R0wPvfW8Dmm2Kjl0BNZzW04OoGN/SbxG3Eu0z0
KZ3nlYww1QKMhiXHKKPA8o5omxWb5ZIQfu9mk1ivpdB+A9tkhMLcNjDelBhsUaBT
IzL1gfx6TqhIXwucYtQxr4GGnkk638REejW308XhW3UL+sTsXAriKDcFt953c3el
iwd046P1WBA2l+Xc1JfwMNGCBDPg8r6WU9ascGqV1wzg/n3gRG5XH0CVhmdKbqK5
C+TcLQcKJlNp4cwG4bh98mgRaP0w6dlIVr2q1gs6w0b3DTTvWlrH7AZNBUy2Rcym
Fw3SI3HzgwY32kJYc3FpG1JdMn0PDb9RLcdVndqRkEbUi9Gp56E5AvhUhQidVfdv
qX9PPUEm8/2jR0PP6mi8/hKQzDkUB5FsqY5rXAHtjfNefyGDGdbE5N8nAKU7JMmm
r3zER64xiks8f+A7A9Fb8hDFZlTxPBjedbfHoGljFOhTbZRl8g+CcEJF0F81kWRR
j//Gz7HYqCfbK9XL8BCg/vkXJMACF2HXbMvYwcwSzNeMv8zscTzmVhlN2yXYpB0k
SrNBlrP7FlK0OHZ91+KcRxzX7bhpnBIjC29gRaXwAz8MOT4CGXaGHPV8N003rXok
WCpAKYEoXdXszbeJRTSqeGss+21/qkg7DG4LjDbHUtFMYCl/pAlY3wmJsGEAcL6R
+BfCZr+omuDjgL4Puh2mZujAaWPRuw3tGCjMEuBezHd5Zx/Rymqol5xUk4KNwPGK
gHo3nNdk6T9+QOkcUrgH92MWF+4AZKj34MC/kZw4NFE2KJBOevx4uQA8/JmMgvUG
E8YyWqMKOdaKbxCUJ2fxLg9l/PTwDWh/QmH8AJL7J5kDm90YJpQhTtwdGCMcyGm/
oN8cSzRkFTGjVySBzQ1tGOx4cTZO9H1JETCisDG74WPL1z2EYGa0FFHhGjLv/6WM
daUDdNAEHel38wO96q5/+rBaLiclc4b8HRtMilE4gQS0gza8xNC0Zj81peLCL/XU
0lQDlAwH/u6nyWHEOHMOQzxkx39MYDw9r+TMxwlAL7GfihcoaJBiaEaa4XsyEpDC
DGRAF2ojf+Fi7TTm3bMK1bNFolc+LgdyBFX20YOImIkm5mkg+ZiiwOLEEkTa2sCO
c3pSl40OcSW9xX+1JVXpa8A3Y0hybToDeNX3xXe59TrhaoL6idKWTzwEiPqtXb4z
AW+rLDnmHNmGc4pXglUaTvXUt4hO7CBmBojUna1s+gnPqKKu7Q/RXG6y3pYgNLLp
vwjVZz7b62jh7e5huDatgJIBR2lAD9ogET8K59jglgXz8fiLQKNCnrxht6kab4M8
O6AfWPdR72lVlXua/iQC3XUy0ekLwJ+GwmRRzEoxB4XoJ0YzIZndE++ztszi+yID
WjYdGnCS/NmwU15SLUXgXVgOOTptnq2/frUB2682C5gpIHVgMguNFDiFOgDVo9gK
Lp6vZfFsUD0sa/cDOMcSRoWver/z43c9aF7bg3klAymNIgChpZlpVNwhp61FRV+C
HrjAzD8MSBxDxkBkdedtS8PgRYeG2ahrdy5vJJYASAIQK/2xS0Poko0bBthe9GKd
PueljZdOxFk1X8UWBXwvCHKkbu/1lYx+tFUJGwZ/6xwjOzy7lpN8sMLyOrOQkePa
r1SMhn0qLMGvPjBBFZgBSNL6TYpdeHP09NgkpkZv+QGRqdNeRJDcGYjZ1YJMLxKj
HmPzOJlDtL//KY4wGMGhIKksZ1oI5hyxA3vf+NVSU1qv179JYJhpIXtYJlkZWc89
BAt2YdhU2Aby9rnoJ3yxdSxWVf2WLjhpl0198RJ0R33/+fzlyc/pYek/omz227Ed
7FVTQ7USN5fLJviqcEQIqsf8C88trx7s4mJj+UQe2zl21HkT5AmxDPvO5o/1oiIX
ISwfufl5lW2I5gMHCIFQWQzGSfbhI2JnCHKXEhwLnQpejdt9vpGs9GoXaA2A7MFP
xNJzNsqjztbihF2mHzlE9J4G+CD/+ibnABL7lOyHOx9O6ZLvUma633B5rU7tcWPU
tYsuvVAD2uzGt7/5/NsT/WeEzpWFfrvT0QECqoLAFDqGd4hJlG+0W09P2P1OPj0t
kyyWe1DpmgSFdiVJQCbCBnpcsjkh2DJA0dlBQ3URLDdVppgCwqUqnpvbs2pM8KXa
avGsqu0+EU/NeVBSFTAv910IKv4TjcNXKQTalAbQqcyVmKIE6ZXTOMlvhH31IHyF
Fkx6KpcQEpbzC52Lp2yk6XX+NQmm6/yKrMAkgFy7XmDFJlm/yczFHEvritfcxpKt
T+IYch1ooFQTt6WXJuxqlQkH+YtlxQKm5OcczFvesIAXu4DkHRJS8SEUbk/woCSQ
LxQn1zOpm7Tw19eaSiHzDRO1piLm8++jp/R+WS2e2WhxwePY0gAiacII3pPVmSGq
hKTlPbh5g1XgBAvIK27wMRspKZ1eWqWQrIuXJeaDE8j2Mi2kl+6hvpwdc5Qq4vXL
6+S3TMaR80GeylamJTd2HOYsw59b895EpS28IBjUuWXh3eal+biUQrsko84nEAim
OdoCro/LmWI4EGYhu9YrfnHPTyxkBWy9j/tKhVIx/3FKKrU2iB/DogQ+GvKfJ48S
lfPW5i9MVmBcide52reNFsL61FqwoSSpRoB/Oj7EUwP+/+w4qaAHGAtnudmI3BjK
kI+ORfVwZ1YqJKW2vfLvnmv9kC3Q7y0XCFE7UtWzivRVlJH4hUoxeSPSt/As05+i
ciz3Xpy3nA3VITAmEah+Pce23CTi+B2OilnwUsdjBCEjl5D+hPUv9/G7rtT6At8f
oJEAwZ6x1t35BIdsFaAnBOOKl63Xmf4Fi/QjcWxWNxpNqg+xxuHt3WPqmhJylPFD
IefZBJIWdhp/s5H4F2k/nlSURSmcOhZM1wkUAWCE85vZgAjIvh9XAkOfjas5DTPJ
LIfSj8OhkBjmqDPmxjO82x6Ah7L0/3pxqUVhrxMzaFJHzxvQ7qCbaW1lXI7ihfsj
3bB0I0yq/84Lip4WRJQpwRkP0YGv9EO8zMYc0tOJq69hbELxzOIP5FvsoyIN++5e
ZpmWmdTDmnmX0su084U/SP2FlOyKeTyzTQbMNrn41hT6GitcSMWkm6nPfh1qbHh2
vIDWKpw/BpeyuE/m+jSYAhT+rKy12VrXPk1EZ6K6xQhAx4oJ07FhqACVh7lHVbWd
92ZWd58TTR8BYGUbVCBisAsXEiUgMJwucQ0bwk/ktQcyKQr/Soa5njADkc+IvqrX
uVMNWsbHJI5+5cH1+kzbdAKouoaAzI2yxuBSXh1rhb8HCmgul6iJpTWUJRU1/Mmy
UBVsNbMVjos9DN1y6RiNuf4WRgWRejg6x+r2Drx0/MWxogFAHdy9Pp59W3Lm00i8
mM75pT1NHg+jMuIcP7iT2M5xZolkzarApzij0YF8TmRbLcf6BxNrtmwVr15bLvwT
L8xeJbc71dxfwUZgPcuYYhJQzWLrHO8J7wWMx6qCj9Uso6dQ3hl35R8clAn5V9no
v2U3nsry+g+vsR30hqHAyhCL64XzlNDtsNLGsIMKBn8LIdygsE/4pjSPpzpfH9vZ
gjgaAd5q1gJ9YkeI2sX9u8xZI//t+V1m0F8L7C7A6TS/UeGKI+FYct1l8RhYpSHO
8LnVodxNo48wzTmRVmRVIVn3UKQvHhpsge50MOcqYm+GS94QczitIFWv0AHcMyHG
7sdIzIURzFTwGdWPJ+xQNBXFYJdUSnPanxKpR7uW1FUyeutEVWaNTT6fqXy7JtHY
OVrRzS6G8ogE7zLfkdI87ViDw6rYi2I8/Wz9i7w58D/xtTArOTL1o7o8qrJhT6O3
1DeRCifaAWAX+XmoO/z9xcmwCJR+srsh1GMGo+5s0Cf/w1YLShjpFxRheUf6D1j3
+KLdTWkICSLg4KhhSjcuVPSNoBch9AB0GRN4FzFh8PaAX9BI+DS3dxE+WrUzbWnp
xtMC+/wehIgJwXTasocpuonlwAW+we2J0yqIwHg48HVU7R2Xwn6K0ub6gqbUrWpE
fSFemCoOQYOMgJkM+SE0EOqJPBwwO0l2+dMGuxi1MzN4ir0fMpRVurqm9c8/ZGQN
VXDwDAvNXOsaqk56wsy4HfaIjPfhrAjBPHpeCeIOkvLC4TvVChgZk7NNFeRG1n7V
UVkPVl/fo2oA8f25rwIrcrRsAUVk/+QovjWmnnLvM9JDVdhPSwrQfBmMxdyU+6Jf
JR6SvHqEDjnFCVcxcTkWjPN6Kxb4gi8eKrScKEOapL80+BM4cF5FWm/v/Okyuras
J67d8xfOBFZzUuIyfQrXKGfj4lIKMQEYae6pFpNNpz3DEB67o+vBHJovX7Stq6/c
ig5gi1hgTU+UxKpchIhcB2dUk4diwayetI8LC4zd5fhMfj0ATSJ0sSzDw0YMAyC6
UvPUvU1f6EPKyAZCP4iZ61tIjUtcSrVTwuXcCTYy4s1ZCdZ5P5DwukDySqpkBYcs
y/HgQdiDcWbK0b9/RDbNjkXDj1tnlm8lCehMpjV0ghpHS8l9mWWAYhqItK2PVpV4
PIL/o7Momhb9l/yo+JXbz6NOs4aif46iPjm0MSY4f1Yx2s8Ibq00kfElzisZ1cDC
ZmlyqWirIVQCD5LNX68PkjO2/ytU7DBIzLOO1N4yR4tWjPTB4zb29Nj24kMal1vq
XoeS3VGzsfPFSaQqzN5UrAyxjapzZhPmQAur6Cp1iag+JBVhr1sYGwLCI9cwyDGk
PLbSaNtE0Cx/YjNVMe0ZYZJrKnmd/fnL9fnZBtke/yiS849kVNrzpPJOLrNeu/yA
gClpWBltP4DuEt2Hej3ickdUMzXT7/kWMJbB6nRHP0uvnSfhHVAx5Wz7Mb2Wnyec
F76c7C0DNquYCpfQAYC3XEUvjFFGPC1AAHkkjY2si6o6VWPS6E2HXh8DLpbO2fEj
faxjjHpLmbMT/eVUNI3AaUl32AnHhajSrYohfV4NUvM/d9+vpGbyTaNWVQzT80AR
YlyQ8bw8wkcgGvmmkqCHIhLi+orxCf1QkjgxscD/DN+sLTSATbEAzTf07KueLLfo
ZK9WbKUVrp/LLte9mbJFpEuSUoVNVEhHCnrjK30X7mc9kws4cQsHyFFu7DbU6n4f
koP5vNzHk6BeL+46eLg1I8cHJbsD0pBS/gmSwm7UpbzBownaHq/n2m0UqBaQ/cUT
Hq8l2SCcTVv+LuND70ggkvbZ8kEUD01nG7YAyyCIJoIySwv6vsSrsxBx+E3xam/G
LmWAeM9VnlPeLBdpYrVmobMAD7zVQIi9TIIp/xUV4Zecwt70o1P/xQfFa+WI5B86
5cMBabZmZBPtsHfDGFW/mpLDVWU4Zxan/50YVzzuFWGLTZUanMcHOdxk5xsbc6E4
z94npEX4MWu9B0kSd4ZZbQjIe+siI5Eq2mYpPB9tITHvSmfKJpv/5e8i3wlYTkcH
9+S7ZYzekiOQCaEH6+m6PqdK2EWBqWhfYEwbInRMBWEO3bzp0Ob4a+ibbXHT8Hxl
UjzcD8tFUB48aFK2fIOQ3mUr92n9dFcYrwd8l8wqcfIKQmP52w7psQnMVROcBF3L
5yYtIfbFjUjmJ/3Vql2tLGfVqcJ8AB6swN4FKHozLHJYkxCaWGYcTKvumV+EY/a9
OJi/iICVuDJF6H0rjFp1OeQUkUk/W6WLsYpu2ED74niu+tY8Y+hEy+DNa4uhpZ6E
O7ud9IUMyJeWTOTlauOa98eO2T0fe3+jiCw/iXIFiCLYcjrAnzGRb53tVctmXm91
Qhif6q1OuM8BXfg3Mf5MoH7oGyKM4dW8d4oobQmLcHj4rqaLgAw+00/Skv2Q8O0z
5FPMrSRyqNMCNKw5iw8Fw6eXZ9twi+TYO9+5pyhRimhKkM4+hK7DSO6esnmpJA1E
MUnMqS3tulJKOEergxxfCTQl7q00F3j5W3sKKPp9Zr5V1Ra+tmE/pQ9vM96mHfuN
rg+qWpcVfePpOy8YII8Ito1qyLE7wqzQ5TZShyY2zcptQxwlgE98K8kNeRByMVF5
rT/jFCBLAhc6PV3hBCuCEPseUhurWBgKEEegOAK+27PCo+7btok+xAyjhalcmEdp
YoDPnZHQIKM+XghJ1sEAfbj9618ekGaiWo2CA1lJBE8S5Nj8ujCRq2olxBNfxsRi
hYVarEV3ASim4/6PmVAdsSUu+nmFfwIw+CMuqbrkHjx1JiS92WQkkGXS+y5GzLmc
6ZJEppngvuZXLTmpewYNgWXClMt0Q7saYWTTIPRBISqFOJj2vSJjXY0fkl5LEuvH
E8bR3iZvjydmf3b7SgtadRUQIQAKo1obXdBsQgHwYXjFwgKJzGwDDHwBL8nAqXMA
HEruX2TKk47oEDq9j83+OVM6NBRIBonUWVsYIlwBYOdwbfCqnDJbqekk9dy1GdBD
iFBSDf1iou7Snl6NTW6FOoYk0mFPhrOqDRC06VWXwnnuPo3ouDGD3O/+KAgfm2Qu
3KFf+wt+9/jOsph4EQblWoRjIFErjaan6FzpiPQio5TURdO/KAr5nOpZjDIzNj6b
4l5SQu5OorGS79KU6cPsyi+b33pV5hssvHAJDSuh+JWi0Uu61qirbDW0Q3I0xHM1
uPrlSqmlA8LdoHMFe6BRcs0qWRgRdnfoBZmmnJY0u1SRQhXm1ftSnC8KWDwQVTNv
VN+gYcMkQm2omg3bKbE/7rMcd32fZy/OMfIuAy7SijgcxR9kEA7ybQj982X6C7cx
SJ7sz/fo2EmYSGxQC556LvDu/q6e6CCiniaF9O16fgQEsiOfCd0ora1paAPj0dHV
Sb5qH5PsJm6kbjUBRA9IUjbxcztPNomj4xVaMz1som1gxKOTogP56XeUTyj0ACGY
mq/wANswH63HAlMhlV2AlP+IpiVLOfZarf5m6iYSvm9IiFJYRru1Eb3YMCFeN2jj
a71ZYmsvpOjmKliaqNozI5f219FcOo+1OaHqwSinvNgMPscZXEVnXiQX/kNSWZLf
e83pvmRpV3H9UJAIlMQDfnfX06ifjpRAj5MWT9MBJmqe3CzRr91zSzwZpOrsGfaR
dRg6bQClHgZ4xS3MHJs3f+dPhf8qY39HNkJw0pzb1NfEySjn51AEb2GHIKqvON6V
Vq1UnYFxkXDne/WhEm7qUBXLVy6qjWOctQS40dvndB3xulcSYZLnEeIFuQzPSWBO
Zbpi7HjpuYWdTjqps5IaK7XaYJxmVu11isUL2DN9xYasPNY0T6bxJaUKGT1YZa+7
gMQ0GwacDmghlHq7KDf1LxzJiaQLsj5hDqUtRDPDi9Alq2CInlVs10L5xBKWEj6d
44M1djT1TJAYr+fbodOLdBaFoG2AHecAIf/g4mbaFUmtIBDsOu6S/HWvU8s9htaU
diAf1avljy20RQBScSq6OPUHKwab26xh8AYsSVl2W5aoao01Rjc9XEgqIb/Imj3W
Ch1rtgvtiaox0ZDrv4WmDUJ6jDk/a9la52nVicVXAIqSyBOIqwGRs4S6KdQK6nKr
mWe1+X2vjiJYmJm7XPtUG0/s1TVRBp4q44/Q+c6eamZxwDZ48En2uhYrFVwlR82P
ShoG51/UDy4cQMeGD4nitLZdoKduoYgT6ElmW9PZBuzZ/AfqtOxb32piIKeWL1GZ
yuD5D/9v34TmokOfVE786qhZqIQed77a30IXDUzYPAvb53isF1fvSPKGCvjOjpDT
AVL5WN7koHy/rt1Cjnfnis1V3rTCi05yKEpZiDVNK4m9JDQJuQx1biFUO88XB1Te
hmuokfvtapTSMkf4odm/WfXoRcWuM0NWweQXuQs+h4T1su7yU6wbZ0F/mRbsCuz0
waL6wkUSkuXoXwSihVHrBO/acCbhWX5zdwuZRFXprZtaxnsFX3oKOa85p6/yEA+d
3ZG21xEqQxXH0zOlA+/FJUU6fRFDttDL9FuKF1skfRydhn5xNZ3XvOOnlvEf82bZ
tWsxvjNij16TV8/gQqHuMtt+s3466ZxF5pq3CnGyPAr86UOEGrjvmeRAkCuRf0EN
F1KwNV5GncLylWcHSFbR3MJIz7ZAZ5mb/Cq3oQ1GjGHposWaZtS8AMyFtNio3+dH
U41Bx3iMAZjqMAJf/EsIIN5qXb7NMLS7kbRIkWcfE4xhmP7rADHPtLv1ZkOrPmGM
Tmk/opSNIJTs3oiYw/SzNCjiszgROxueUUtmuu7HaX4lUpxWmSWibHS7ou0GhMh0
TytKFsjQkeqD1+Ymoeh1JnEfteVM8DxC5q1h6Fan6F6YcqOU6yT14mvFdrEhKUXC
SIbNcRLoCiG2yRHebEzA64HddTSqkZgZnB2HiPpsA1LlLZ1Xr87tLus1rqBqwbqD
4GI3IZJbfbTTI6cvNyLFrBl1zB4wPiD/jCA+wKeP+/vSbPj9QuypzQM7CuntO0hs
0nYBLolLLInFmVDzCiN0wZ4oPqXxP9ZpOxsKDPNP/r/xRsypGjfGXtinn9Kp/nxM
/Tl5K3y+uzS2IqfhJowBz2ZLpQTqoucWmaXaGYcyPtHi0NMw8hAyhGK/TWMbeJQ4
SeyPPHdqDNvCCiHAoZ5lzi2EK8evpWU0L+8AYnGQY8ziEafFr3DaxwUZb3Oeg5WA
HRfUYGt81k9zOsRdXNToWyts5IGUbBGqoOokLVHKIf/FAzfXFeEuzEt6kg4LD+Yi
U2j1cfhyoUoLucFG+lqEKGYDbv0r4hNtAkrLLE8H0sVkhTpOQmP2LD8FtFFfiKEG
VrsU4M0fD0fYcRY3cvdQ4RO9+WELcmcEqbo8ySzVGjGqAkWHvc6HXTAKgiG1pklT
JMsL4F31MkeS0IdCg1mWPNhq2wWX/ZNJfK1sRd9MtfcqIhlJWnU+lFWzbibAqFJl
PajAIzpHDrYXSqcW+uVdX8zTlO4SYWaUYYREKl0gijO5D90bqNXg3KBj5uIvIlUp
ONGbmc6EIsIkQmb6uCpAiVvpv9AncDHZPSn2MFSoE2qhsyr3cvTHvaEJr9Qf6mnq
DuokvUOLUcqq2iCPulrf4KEs5F0LonrlslsoXfSTTxDj0UXgGrsSyfWjnhj/Oak8
yPEPhB5w6JYp4qpOUjMAeSHPYJbPt2xjVs9XB1P7zTaodm01VJikrTEX0LWmioYK
QHUeFk0cUrv2B8oL0Tb3LyN03IAeKdsdwcU1X53btHHJ/2sRnwQ8jtHrGfv3AzmT
67qW8icd0m0alfx5W7W9A1KJFKYVOmmsbbLtvbNqgRj10ndzbMM8JqsIJBNKRDZa
7FHR9uKwrb62qDCP96IERSP9TNltnuaZEjZDXozvCDjHCB736Aa2czkn9ObNz1io
m1a+cldCSwpCBubDW2ZO3KRH6a0sg/r7Rk0ARiXaesMd62W2RIPopmyjkSI7vM1O
rm4uqsrIx9hu8w9uGY0toWDJ5a5/u4ComnazKpXzoK9uzbOo8/uywNlzCA3R0kki
aMHn2K5lL5MPTKuIFO+t5iFVAdTDvx9JFc/5RJa+HFMnS37h0kCilbpDIbp3EcmR
qpZcOiYt5nvJvr1ZsD+GxWiOGiuxPoaMqspNNiL+Y06vQPXFQOUf4spMM1z+bc6d
/cz8C36Onw22oz+Lkjq/SPqosIgaT6xERXolWlT8GIXjTJduUrh9r7IozIxsRO3A
E1TTbGhM5wsMWFJTu99VucIZTeV5iPdXpjdnZmESnjn7KX/RrntMRDL/sJz2+Ter
W/Xf6BxSDV1GP+/vQaGR+wOVeDgprZWpxyFNKxxXaElVf9XjGRQ+o1N1Yp4GwkGK
qOnUxbBDzkOmhD/wDurIadBeyIJE1/BVd/Bv/qSq7UU35x2mck/pcWjkZKvn+hW5
Dfk0KIuN/79D0Aqu5sF3b+TIkmiLRAK2TpHIeQkHcnfXC4LvWSCDdCGXBgvVelin
phMNvl6aeU33w/hydTLZmb+anv6gQ21XJO1X0P5JxLppBGgHfaLfSAKVC+AJkqed
XeoWwQ8e5HMuSsHZ1ig4fbvv2YeUMEEJtn685nQmg0rw7kaOdRbcB6vQZ3mWSKQj
gthPX7TVe636RxHZnZvA1hPSZ+ZmRL5uGkEKnCBEVs/Z9Af3eUwtu/vnNYhU3qMF
kEfBZAVDbIHbC6cdBHgpp5iBXNdZ5cdX6+/Uof5O7XxuxmInnaD7xelevSrFX297
Lz5AOzQdqnkTcUPd8SNJ8IgtarCkSvFmwzkZwmzGS8I5GZbeqjKmFg/opPWbOCF3
+800Il3UzASFRk6alSUIjl5FD9354lOtBQusRLJNiy4gRVP2fdnj217zb3UGN06k
mO1chG4MwuZFtsw/wJt6zcE3Nkh0UkHftmsoH0AtGoOWbg9zouvKS5oaa//bu/hG
RsAdcgrHGpIOSR5/sKgIWqGYcejb3Ul9d6TLBRxEXYJNWiRvuugcRoPP/zmOBOcu
v/QVQSxua7tX9R0maiiVRvDZS5CIY+Zzh/MDUeIf3vZwjP8wHQloIxjvtBumCfI6
3q8hSUPKqgds+mpwj7lFDNTX8T6B4sAYP1ovO5XUz19nzPNz8xson88QTlJ5MzKX
eBGcYI+kqRJdLjpODAzrtk/WMxBhQ7o/Sd6O1hAwchz96apNI4dYkqEc4K0oOteU
f36PfV7EES3fCGQw6hqXvVnFWiMq8X3jzNj43oGk1tZtY6HvwjivB6k2T3fjiJS1
LJX4/83ZO5zTT2iNFxh30Of3OmMe7iUMQ/4hE2bWanBgoJBO/ib/FkrxnYPVBHJZ
d1R3OHATn56O7xNardee0bjgnEVlfBC3IEoms32Y2tLnEkux0upBwQZkXjSM248D
SMc7WZJx6CQS3jDzW5wLDlbIRGVbssLAe5rHdZQf6JRZ7yvj9ndT2jKQeH8BLWZ0
AMKZQcLdhNoLtZN0vDNnShjJ0cw1HPvYdwX54eTET19jgZpz1Yo5BtbsqN+78MB+
fB6/1d10r11EOpiNSKR5Wb3ztemf4WfRL9z9JC0RrKcrRbiXRLa5goPrn/oZs640
RZh19xn81QT1Ldqdq0iygOxpgppIXpHTYb+axVlr266z3GTGTy0bCm7iHH0JOPit
o1qUPYOHfIWMKMpmMEx8mvVhqN6vuHTD5NRs8U5XwbL0n3ewMfVwtepFS6eNDoBR
3LmOv+LDY6PdV/FAkw28GiPrzwuUr+8dVREl0DchQRRDM7UpSItvmUaUS8FxtI1W
wARNOOyqKYBui/1gd0Bj/2PK+kmcQ9R6vpDRx4+YeSlQMV8iZ5PB+wF9cor1AWeH
YAcaPJhQojxDXnsR4U51HsSGuQoxvUxZYfb9rH5n3DPlWnSS75BiTsfN+PI60im0
wtMX9KMvjXhqhutL6UzTJrE8Bp7xFGzckNHGuUQPREiCTTkpqxKMRK5JR6HtAuT5
fPlcn31Dk9psBp72LwycPvSaUd0jibuDGILM+8TLYWKkPKNZUGBiF+wuL3RDQiIN
rh/72BsUb16bZtz766sXepCnvoFW5eBfJanCEVUwZ6W8h9WbpyTY/2x6P5IrErA1
wZ4cbOtcC/MX/8MEFZft8PoJq1aQ6KP5t0tXHiFE78j9lfrhXbhgmp2i01Qi27TZ
uTFt6BpEUiAfl7RedMi1ioovStzcpMZ09UuiT5nHjvXXyE+CsxnPgJlbQF4o7l44
OpLnrCbta8F8r4C9WTUu6aiFvTjoobJ8xfKNnCVljCL5GXihGY6ZIrFttoXtm5+n
6nLh1CXaVPZPsqRVpacWsZHWlJYpP9sIqfnWkOSmWD24hIhgVB5Wulue16BTYV8l
EaNwT0vEaQtYCDyGbSX5y3UjZk4jdjs9oKSuujqjb7zTQy1/AogQdYX+Q5BRvQE5
GubLTBuNcsatIzcta/E9rtCpJk22fhc02CTOneG78UFjsVVu8f4ljAxKKD+wPHnm
rc+WlHwUCGKPH0YsNxwfk5nT6niyR7qPcyfgbREQiacgoE1qWTFA2sEMF/X5CHgv
QY/FUHam8+J+E8ktmLiVD8CBdVknDzrkUb3/CR8gu0btigrGiF1IdRhaPVqMJodg
wsZtzO3JGxNwLdVz4bI8C7BEt7OET4THRm7jMXR//BjPMfLSh8vNT0vanReEILUr
+8EnIlp/srWTUepb04o06A/sqtlel3zcTiqgqsyeNRIajllNPge3LS3TdT4ktqBq
l8MgDkThES9nF/ooAv3yCIGSR8UtNnvZzWomzTnmQJqtkrQBXz0g3L/DUt9hggQz
Fqgd4sae1NyeHwFVeI2vgswY4b9ryJd2A1pjydNXZFWWBOT3ZKipYYCiFPDVYkwh
8dhobIpNRP8A4tWN6NVwGcQ7wv1/JxrEWh6nu71FGxCoP0Bn7y89/CAcmvRpk6ga
X21zDmVzsEElHZY+u5uNSMos+JjCPLHZQtlkOfZZ0+8kDZWAw0bZAN6H0dMrJ5qG
SQYvMuMqslVMDYFmyblyZH3up41H+eJv5JBSGOFmaKGilPnNeGceCVprIu5DAZB+
gF/YXE4CYtmfEb0Ml+WyQ+GWoqVf5d9G57smDoQ3cq/gKiBjjtOEdRvWKguEYlSe
rbgCtb8DwmxgoN29GyezV+H0grrNVlTY5TKAPxA/XNsyoRVspi7HYdYnpmPgRRnL
OdoF1xohK6njxbTDGQbk8RQ7I8sk0lv/uMfrQm+BVYDwV6c/m14qUkh5cZ+Jx05x
CmvTsbwW479Y7NPq8JOSjMYAFbWcobfdEuAl04kFOEnAbCBcc02/ZRwRH/I4SS01
O2dwxcJUH1ZHrKM613rb2GQ6m+YhGsRDCHLfQ5DaElvy3qGCkvq/pLM+gu/+xnOL
LRx3XnZshGkKrJCPHwUvxmwAH2DwkGlZj4c3G5AwdonRd7swA7UI388UPQlv81Fk
tpInB0H8VvjqPXQekvF7QOhoilgnHZW4xf8KLDlzGIZ2NVSHeRe9q9IZvhLjwYg4
e4ifNrhQnETd9fBZwn7IVQ/ndn5EmVL+bO6R25wmFzU5MUT1YAuO0B1BQjmIT5rr
7SaM8st+2kodyL99dHk6X99en/GtKOT5PS9bzQPSPWxZu2B7NYhs4wUN1f+y/N1T
gtL2rMeZfA5l98XvFzT6oxnmVCXkp9TlLb0WcX+drqWjz9yVS2Lru7JJ1sljRWOF
1uFebwsJXeJ2/igqt1tnsjstGP90xmvM53GdmI/VOyOC6CYIYjuqC/PpH/y/BMge
IeywrvWSsTUUhiVZwYPEtz9TZZn+ziHETXoiRc4nf5KsCNOZztEEFQLsYbRLHLwG
mDsKP3RFiXifM7BYIZbcU+a+UDus4/MaE89AvH5xLL6WES48YNHn3yRLDRKiL2ws
D8oXqBEYZfJvrhiy52nZoMkTAGBc+ZyMliGFaRs/8nSOETJpJVWfy+hH7fKU+t1r
sAaBzQVhzA3ekytaGQCbtNDmyJdmAbvpp3ciVd3/sGJviH5kyzKMABkPZJt5cpyR
qWbG99oCcRZG35qQJ3FYOS0tWLTh40JinUVp4CIciUKc7cuhmOyiS3Fz8MFIoI3r
NwAoeYXmA1saq4ZMC0JrYyEMTgSwbv9Yg7zgXYO0Hwf/IUkwmlh0SQpRMnoD3lOW
CKvbUUihf2WFJwAfBfryJY7WSxP41Abl8zoeKfCOkOwkRlDoQ7sKlMzaGgld44G1
Jlw1fDrMcMDyccqQBZyw0kQ1Plu9XfD836HeA/n3yx9jGn3NkhqbW0oKvcoEA2lt
032MXESL1Q4DjmWlTGojWauYBT7CvxL2h0lQD0MCttxyOx994Zfy8KWJ0Pm10Zaj
B9AsCm0jsxoNbPmmJvSAR8BRZ2a4aja9wKBBJkshWEoARJdFKvn0vJDpHPDqlsD/
ZL0waReDRxJ2YSipEXFWPqT/rl65ANQmehx5k8AcuPLJjJ5ch6/IjR+QCxtfQ0Kh
tenRDRD03cguNS9ZjaZYyL7RzZToGnqZSPlUbQ8SnYVYMNc+9KnZJg6/EKcIR+pb
plgU/ySI89ypdnt+LtcUb11aDXP9Gc+w2jnSrBWg0PqxUcwRvrUrRv9ETlHa58wU
CqmVclV07ZoGCK7FCtvVO4EK/0n3tpjLQ1khdmFt5e9Imn7uJ1NYuFY7GeLTPzZv
2c9f5G2iRcrsVnnQopVR06ZKsQv1hVBfP1FpBBUh4mJG9i966oKLqO5ZVXbGAFwO
T7IbGaF3VQy03ng7qNKYr5/YgJdWnED5MH+E/ifoRQ5OprtpLwzAOj1tjtDbMF6A
wsaTXTa/XcrwK4kSVD6tgj6gUbxqwwFSgVENH+H1pU792UT0iRid47k2y7N0M+gw
GEUiRxgSgVwG0NgeUhyBXGENtQqk7SVnhHzWqQNSFeGAnQDetYtBBUrJZdFLoEuY
rH3SOdUnE4ZZptPWkmGTbwsMqzx8YXUzvbJtq+jquE6cvoUHPNjqN5nMhrln5ze+
FXFENwvMN+46v2ez7zeE7VPt4Xe+MAjGYQBbV2LxOPW5RK2tvz6ICRFQFRC1XgA8
OVAdxQFsZx8vgfha5JkruAJ7RBj9F2gk77YJUh/hJnZNrlBLzp0MOFT6RIbTSczq
m+Gn7JG6vaXM/Gbef8KRSJxmMQAEb99FO7yToDjkPq67+wajopAp/4MLNQMLbjOv
JKROysbG82mGOldns++m9B4VEWVRc08X1WntA0YgvW8eP8wWH2RyYPfIZ0mJ4iuW
xIzcghBIKCMqEeFvQBbLt+wRkvJzahJq08dIpz57C7cElBM8zkVegIofunyJbPlk
pq9pyBR077EEVDr1GS+eT/WgeWrjOrQzB/zs/Td8ZCwikDDCAd9i2P2Dtx3w1OOR
RHh2Xfj00ZEgDZzQ+5I7yA==
`protect END_PROTECTED
