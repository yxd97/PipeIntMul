`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hwv4iF4/UTUz4SWO8WuvCt4Y6NeW9YQuMJqKiY2EMq0kzDpTXEtNovWshje+R7e8
RkTIF0lNRnVwO3TtDYcng7kf+7wMMGUoFg4dXYH0Gg9g2hGPn3BgcX7yQqjbsCPk
n/7PQ4cKeIZhf2d4Pk8NmqoCcC1O6xyarVfQNRWuaTd0LJX6MiM2T5a7c1sMdrvz
ITNA/BC8msfH9UudRkXu/EBe7yQnakcpopMvxyYQH3bEbtxTWOuWoCTZfFjnyymT
GjJiCV27ahiX5vL14NYAs+EhSvtnw6M478BvjwFPnz3Hg3dvi0C3ZQUPWOmKThE6
`protect END_PROTECTED
