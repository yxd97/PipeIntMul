`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5t7rMFfohcr4eiMFRf7zw56H/zFY3v0a4lxpvofttOcMPFM6+eFT+vry5nECHFi
Il44hFKiXfoLVhNHJjnTfK9tt7zqblSHMnVCjLCfGvpULn3V4daqH8N94woHd6oz
fKj1mSOveA9vv/Vg21GATRueJbXswOe4pdoOpY16msQVeZCZxTOW789gWBHBtKbN
nfzTFYtehzSDNOLA0SgWTYsG4Fd6QNbmrOEinWT+xW4sFXv6lOySauobNvMjdkLo
n+Vtl4tsJiUO0M8Ed8yWSPQxRUdUwcOfddMxDP4ltHcIZX126OMdD7YQQDtLQDn4
w80inwZnQn12LShSt/r5Y0XTw9X7Q9rtMvw12tUSvWNEdlfZSMqJ0WDilfrxjWLr
jjVVdDvmU8WSUHLLVeuWqEDX55g7l7wx7ELnx4lI1lE1pI8HzNw0B0ynHW0jQYJ+
ELm7/pVR0R0cVlfAbFMW6W6ZQOQ8R8/sBMGWBTGEwO0bB9RlRPanuLFN43CXzKko
457+mVQeKZk05EATkLAmlfHI/8mFRxKX6aeOiKE0KwRATy0NYpHbd8FDv17VWEX+
EQCo6tUMjvP8IvCTb4DLmnkBOaw/oclDkhiFZZyfvXMT1YT4YgBYca+C2ElEZ0G/
xUUNEJZ+wDjCVDgShcb/9ZxntW2MahCWuXJCukZt02M=
`protect END_PROTECTED
