`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TljJGCTUZfqhYPuRdFvZKLXzYJUw0Q/4sUyFMbjfG5ClGHZxcJmUrQYfiNjOTsgv
73xStdws8f5og3I3WSNaP5G1khN3FpEocSO2lvatjzECxFNbAPmLd674KZyo3Wuv
9maQ34vhwn06etSsQN2oJIC9XUVyDnS9T+8BIaERTkzgYrZv3eGazZM5YExuvbY2
wxmSAg4oJnpjXl7d82oFcB8FTbifA9yT9c9W1mTa5j9zqynsD/Xl8wz0MCRpYCFQ
`protect END_PROTECTED
