`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eeh2cfoVYrQZn8tLHMm6/T7u+CNlJpxoUk9lDijK+1azu18+VWpQStGZm/N73oKl
SICEAGli5Ro0+OzGSJ3wxZYnaBN3hdkU9/vxNWhjd6GKAWyTiR62pd6SYs7HXY+N
ZwlCZhjUBsmoTUlvWz6ZZdpakVfU7Hv3E4rVqOgAo70WHN6hKYW+t/q1o2+H6kSv
DtWgXk/FtG7PcMvW4Cp634QtT2fc7u8yx7VkG6g0Bjo1v0GezEDHstg6rd3J1ExD
hGy9QM7OVgU6NxYezTbPd/0Z0OfVqGe2g5CS4YNS1GwzwMqfPvFMYIw+fWrdGZGW
5csOkhcnyoNUX8w6V3D1zdWRm34aqMeYMoemEhjFPx/V82cCrq+lpSJnA9/H2Hxf
hXnSY7Sjw8keomMOZNr0jJCPPtGt+7db626fh25ColXjXNfNMiKUUg0ZaKbzCHMG
NIZUOFqonmEqewbO5koeFb0pfeMBokLuv18iySZMh2+yYt4vlPsuDAYFcJ1dX/YJ
uKhSC/hGwNpY1hwuO4jvbpps7LfeyNdgCbsP2EF2wE7dUhZlryjQdvDU3R3x73Bd
vmP1urVpTV16FsGLKd4OkBtr5zHWMJRWpJ5UhirD3x7KJ8HplEVb7H1cA+BDIbtt
+UCSTf8ofE5Fx0jA84n/apjXiRqkMnvbOQvoWisQYynkF0jRGcLthjt4Tw0Ksbe0
VBRnIvJAPmDrZZN1wgGgpa3EPi2kFIyOW9pRzgtJru0XADLKGEQtbvBdVvZhlpB5
6TTIJHIomvtZuCAxEZROKiJA91X0ChYO+iEgSIK+zrPjmE8tWrWK34zugCDfwk4x
Vgrtd1c9RS+lagUbnxtpHO1QMaRqek/N0eizLjAt8GbCS/L4pV8XLxC19dwChNTc
5AtGYuAB0atL4iyln8weqnik3mg1YwtRCp+nffUTX1ur7Kixty2t63F+TBdM4KWf
Yt1Mopgd2TVySrjU0xP91384Q8GcER5a9i0AiijCMT0J5FxeW91J1DjbA5KOMVGL
7cLdFs11+7KCl4AabXOZ5IcfuwDQEYfCa9dsjEKrpdTSq8O/GMb7/GEEtTcKLoCa
PwyIyou0NsLzjHBQBRUTvX2JZ8gQmNODlCMvgmxH6fsOYqLUld5tcrKCHWtrilJK
QYVHJSF8XvH+26viMbbRfoXAQxcwnHqHycaAC0rjiV3q6uVbwju6PVm944vlfHvr
4OZDOTl716ixnkWMg0L7vW3GgBqLIJW/nWVnHlBKtPRX6LMSnZKuEP0CM4wbhHCW
GqtpyJNVdtvdiEp5IhHux/TsnJn0CaKtCoIsgWDSVo2xdlzRaadcnIW5Cz5rHloJ
6PabjTOPy56JapLnCpXjzw0c8CnvOevZjTuueTJ9LZIHiNhJOy6JZOfEnMGWyQvr
KK3nxIpGmkVSjFLdTo+xKmQ2dT6lTQJU5bLOHBP9eNiSGmOPBc1BbHM1THSDn90F
kqseVM4gJ5jTglOiX1RQ2A==
`protect END_PROTECTED
