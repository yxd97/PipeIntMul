`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuJ3NbOHSaj6Tsks5tTf0MNPAuobrXoWKJ+aKp7w8Gsf2q/x1cDgmEMB9McpcVXA
F8uQXkMT3kvCZ/yS1qmrIruvltmyKqw3o0mHVcQkmfM5R9YjjGVRiAqI67P0zMwv
uPa7bkKYJZ2NWVE8VscMy9uu64TvRFNMemLRKtFxdtos9dmN7vp2Y7rXr7i1fJdX
kNOoDW+jZ0tH53rS0AurElqIYhLo4zVVbMEOLdcWfrA/j64LUzr0jCAJcVHBCD+y
OzD9t6+aJl4wBqvnShAdx2DytNC/PN7M+JqPqGk78IRPqch9wUjeByOYBckakrUT
JbqMf1GTNxHNBKbELGMd9OBUOa4RFOPbOSgC+/js5LjH2vvI5hu1FgbM0Fm05uXA
MLhO5uOMjmB+QJPDffGCN5oZ0aWf2eJrKB2n95WSD4/JQgD58T0RvLhrynkJsEFd
8twNV8Ok89sGRZGsz+xau8xsB1EKqgkVLakt4VKMmssJz76JRBtPTnbYtCptGOEm
EDRKH5uyIsIJgapYJSJdRq4xBRI5ddsxeDITIhvSSTx2OFRJP8eVLPZVNZE52LOX
50r/kf6CNGnjuIAhr3lDRENOlOQD4SL5P3/MH4I7VOHCmlphaubvM0sXWVUKYe1p
r5yMaam4MdnYWBU93tccCcvryWxdVurbosmZEKng7Z9XlDQaT9hxcLxH0gdBHIgd
U0YTLstH/vITH65DGVKsbjsQemZV1LftKmZCA2aKQikROdUOF7ZVZ2mGJqvzt6AM
Bd9kwRXbkXTG5mtkUXuVlB38QD5T5yGXprzqi79OF4lrJkCiN+1mNEIk7P3RTsRq
5kmtPcQFx45bmZM+AzcgmQkP7heLwuqgjLhSrBsQO+baLik99ZyNQluEZNuLAUGA
1Y8hCFVgsObkti0l9DwcwFsRvg4h3bxoD27U4EbcW2HEYzmUjmgCPghGROQE4GRS
fNEKKFFXBrH2Zatt4Sj9WZ7fqspL50TsMqh1AHzjvlBgoCtBQ+Bq11gmOgYCQvvf
SmwmWZh20Zz1a4VRVdzQl6OeSIfoazAwE5nscEc0FAJ61OYjdU9XCXsnthYCA+yl
vn94Y8DlGd4HPHz5iP02bMyqeOpmoW2fm4vuHEvLWgcK8+uvyRWl9DF7L7ZDExFo
T3uCrghLJmPFnBrRhydxCdl0ouMKHgWfctOCQET7phkDlIEHvVRP/gAJTHHdxUMj
5jKWcJNZqEcl2HvrgNx0iF90+ddwj9uJzdDp0j8gqgk=
`protect END_PROTECTED
