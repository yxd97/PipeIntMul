`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bKv2hAiIsqCQVwK8MxTGc2+toxCmA5NcY/Vd7VUO8WKxapzHqie2OWI/QpNw6rg+
BeY0Z24Btz2AfbRvBiCGlxi/urJCr+cdSM9oY14m9TZ6Q+MZ7JTHJG14jouuoVG1
S5TLL+ierK8QWLOoSPTzFCvXhK2hx5WndBO3RKi+4m9amfDpnNbLBkqOIzuZGJkR
3YBaJyc0qEY3QM8vBI4jHEl884xUmp0bCDMSS+Hd0hvvLIrhvuRe2mmMvDUBNxU2
mvnNVvlldHLE6YHpWZzjYl/z9WlXcbJRTqm8qbV38sTIhSjD21serMU/ilEvxf9M
J0GND212nqt40V/ISZ+COZuPCD+S9yJhC6znOiWEWS9JATFiurfD0uzZNpfxQ+HP
Pkyl3h+yp8ze/ixACzRjloVAaE37ZWkuPGxj8WpknwPf+vsEPZFNa6CbFtFmGYj2
cQBpStxjwsYw5Lj/qSYbJDqSbOw0KgSPemzFWqHM0wjJF4s2xf8M+YF7m9R4zpQY
OviKJErcjgAdEezjS/9onbzpmBNru8nJufsX0KDTUkdWwk3vJCDEohOViOezjfOt
3y0jCS51KMURuV9/g7a8ow==
`protect END_PROTECTED
