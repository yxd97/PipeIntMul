`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L3h4XHvq0S8MfoBcuzzR2icyraaeHPJUP+LrlE1dwZzMsifBkN2sY3saZKzMfys8
fVk7b3kkdwRaPJqHfyysA0VGKYLQwW3EnoheacAIaTheaiZYi0XahNWKcngvmHPR
DZbZL/D2U9MoBFE6Xxp6vDVczPaBvjdFrbKRXNRaDkVLyFJPpj77KL6vde6EDt/r
ZAYwOybwuCgG0gTMqGwlsbN+cOibeVpGx1QaGzrKWovLhmu+S5aLemdZ73sujka2
`protect END_PROTECTED
