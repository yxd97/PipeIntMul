`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhmGA02Qi6MPBTO69tVlT8HIXt4QzkEryeNZS5keWpUzXtEnHheKLBq699FtXMgr
BsuwfpXNFmpWDy+37sKBgoQ3IPSd8FsVWVCdgKuOU4mmxd1JA33UJf03soycDkU+
pJJam2Ool7qkEhsybpToyvUuyTYIR4hKAbcZmamKfEQIbvs9HXlDTpyj1vZVgWdx
uU+S3UqilTbobQzA1Vz/ylUanSnV75O0KQzITgGiHnMFxlHAxTOj8G1B9abab1By
Uh6Hu0c7GxBOYE7dL/14vqcwJxV5aXGzxdNkXYbS3Zo7mNILfuyBbLCB1//N3HVm
9DlBGcZ9p//vyCRlWvVjy/SIG1Wd3hnBFFrA+ODWyydr+0EFN5SZ9KHPH+WKW+Uy
ff7bThv61LMn/afPlwxEP2/VPHnnR3m8cXSEOICZnktosmCWWgqlJocCFpkgpVSg
iOZiaVRr3lU9kzao+HDRcIu9209mcpFAKbIlB/AF4m2g2bIsNyhbQDROccKQgE4Y
7PyhRaZSc9zgMifBflLVXdBb9G/HWxp2jbnzjZ51yeTeZ2ZYLdmqliMjMB9NJRbR
ihAGjzzULtnNEWWkynOOrcJEGDyBUMzE5f71FVvpS0FVuuQO+Ph4JVbq0OoA5bol
`protect END_PROTECTED
