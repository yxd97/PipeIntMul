`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U+6t1NFMISNiZsRFNylEycR8JlUkcFKp2ClydWCUq9Gr3AmeTGUeExe8f5ABIpi6
5b8IyM0E+X+OPeagI3Fvm+30nnPOAPNJpLPfPy9ixT0HQSUUz/MeWdXcsaLq2Wzm
23PDwIIEq8gy98yHRZsS49a2MLUaCVe4sb8bfK9qedSjl7j+c0ysOEsnUE9LX9eA
88rL8m3Drkpm5l5tDj1CfpVVFBBTZT14zf5vRK13NDifTZKNoQQaqnZWF4Fs8ErV
AHTRySq91wBtUqwydno0dmd6wY6vxxw2KeHYsVTSLXHZU2cSOpoG3cAiQNOBRC0C
CYfOXpTwOYo2KqybKHLIKjbjCqndA6sCTFPBdA+iV/sASjUICWhjM9Kd0Vny3SsH
o0cbevGt0DeNAubZ5AGGuZjd1/wuU1II1xkukNgtkfY=
`protect END_PROTECTED
