`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/SKMxNY6TvFBPpnJLrDs9hLXrxTNLbCUNP5LDi7xu0sRwdmQe8neXFusIn9bWss
miL5tKf3gEGc29aifoXNwTlHDaY5OaDkLUpk9zcovoEqmMlGFcoIUhIkJBeiaHV/
gP72rkOB8WBzrSUvctuNcn8Rer50GIgYC9Zj0uS3cp32s4hdUtevx0U29fJrw+kQ
nhD4Gr2QWNhWFuUt6TwIO07EchfDKqbhWUIbqz6lKj2sHyq38WG14pY6Q+aVsRx/
BZHgp+OCAgHr2EhklRq5ETyTBM60k9ZcEO6eeMLz5p9vnsX8vliAfx4TpYvUYjW1
yJrs9C4vxOO4b2vZHwaqz2VRG17FDvGKn/wbtS7gkKiNnT5n4qTiWWACHJslvMIS
A6fvWWZzSLIAmE5QbTZCC+smeNzpP1S///3s9ltlk6jI9VIIyp6LGg/o5kDYNA/z
6x+uQsgyNE8/AW34fGeD5ukkpzjsBxMPyqB+uh1nkkS6L6+RKiMwe94X28FwQdVc
ORIfwozQAzXLBqcjRisLtuUo/mhdu0gSbodG2Z4Y8aPd/yvTNA6ZmjH1m9f2W9sU
aaVgFPDezBeOFMyUcn03XJDqTZMFQbSxA2aU7pn3TeFpchtD+uWoLUWIHyYa+8Qj
DqHZzLz24i/DrJmuCQrwfHXtuRZXNDV4/Nl7OYlPVUszeb+8t2H2H6t+KXtXluiF
zxodj90oQH6+jgGoWSVl5ePzQznU6LocJtzq+RBaXGFJyNrVrDiaar1DtVyPfJpq
D+4PwomeKa2yXfQCL0Rg8wzAkVkKiNE9DTaFNjUT7843A+pwD+SQNwamL7xaAl/U
lq7oXNTeQmLIksBazCwCfWz8hfEKG2FrqOZ/hdh85MpuLoH7K2vE6kFRKQQwMej2
qQ+PG0e6KAcf73Mtwt2W+W4tKJcWmKUIGYN+dOtm4m4WzIhgObRNNMk8rasTAGWu
JTArUbuoCti8lF4pekzhQMKxFQeaYN7FtTjyb0QDgEOrXckC6J/53L7pl7NuiRAK
lNkp1NeOT4Gop1/ihvWwOkO9Rods6Gg5GJ9gSxTWmJ7rKh/Z/dJnYB7pEQoeOwyi
aGGXF4PpT/6BRuDrvZO5f62mdGWKV02TjPIgTedTlOfknGWLVU+fg48zp1kQ7knj
BU1751aGzmamV+VqDgVm9EITtMy6jXaq6oaeylqcXnOXSxSz6G8MSJo0JUPiK8Up
hPUjQdKCBvq69ZSMkq67xSAj+YSFSyZyB8DnWe5rceLZeyl5S5yGK8P+EGuhKlQM
NvGlqWjv9dkDZh7BjrY4XFTudAy9diQgdH7w8hOW5CPWYLga+NBn/itmnLojoVbO
tG0DhXAP+xtwtMckJmvEA531WIlzxQpKAfr3CaXrXCXRWhdPlE9Vy+zMjud19t0K
HJHfU8MWyJxeBa1jz5NSUW/CGkK5Zbj42tymqIKxN+GQmp5MZek7xHKJLonx9/ob
27mk6UuykfITL9RUHN4NMbqx9dVuTE/knjYIjYUmkun9Nc66wayjN7nlBGEm0GKa
CtGSg6Iz0m1MXTAD9zBqieE2b9mJ+Celz+n2aq/Y+PPziMQ1S9fnFbdx/XxoNL2j
CePDa3kCghR0ZcoQ1IXfC6n1KPUYuLzWJ0sAimtl67EE+luJZomvy4gz+8AZWG2/
aLRZu4eg2W/jXhq8FL+FnvAeph7kY4/RIzWWjT4I7l6SFT+01RX1x0k0h5S3LBse
gwxpSyAbT/YHYJifpi8cg5FMKYAN1mdvC1xC+Uw9/8ygwMk5hJpJYOVAhWUAzy62
qFVP4f/G06obiHQ3tChgfeYQ7ppY3Pv2P08d6WegkBPU4DpajlsBqIFCCQzWvQ0o
FuL5KTSxziRxw/w6JHnJdbeRtpguyQyq3Z6HoodvdF2HNK5N/cYuKNcWSjy9xkqc
2SNObzTDwx5Gerq5mBm8Yl1IADKoOpVxFHiSsHNCZ3oPSwNnM2wIx+ahznZvTbB4
oApEHS32ZY+CWh2DFFgQBsCyJoLQ3m47QCxw/rH88+1rZKTvBCvcYFOdNBpy7J1c
DOKIt+WgW231ky8vHdk7SKINYVZlCSiD5/HvYKs/kicGVY1HFcfbQdSkQTLmPsxI
7pt8Kcq8nj5uFPyqTkKUpv5C5VTS7tsmkuuhp3JSCD6k1e1IQFXHjF1Ogdq8ipsV
L5V5dIesjEww00QFamQgE000hq6/us4HYFPwswlVZeCrE6xq9ejwdQui4TmRP8Au
eaN3UsYi2maK83cPaXjJhDLRnkmYW+4d5QqN4qFPhVTEDFWKzLkv3CQu9VwJ11d7
/o3DQnYHSx3U0sIg2ICODkD9161rX5K04AtQ0CuXSiwzs9PIrD3+/yPmIZ2ZguDe
l/Tbgma1PbHlOqAfsPCmwcpaFiRKeLrg6XS4GOZ6YSeCz8CYwvLCySb/7CQ6g7LN
4gfrGHJLYB5dnn+HukmOtY2wu8iuGtXsmhuJymSQDR8v7CwtfauE4L2AuP8D3YJy
P9wGsWp8WKETM8UmxcgvdHx6sEes/2I/akftgOAk0g4/Jp6ro04ksYh/Elv3VWSi
WzEJybh2Zljc8z1HUGF9Pn0v7PgvGx7nDa81wwBslrBSwIqQ8bpxY5I8oZ3gJEv4
5kt3cDOH39s5EGuXVTmDE6w4FF/SC85px6AyXWbH5eBGoZjh3rQG0BH509K2pJiF
/baq8Ozkeh2NX2yxD84M9QE6eKE2JFvdpv+BNB7Jt7Z1/ceuPR0Tfouwfzi9sCNQ
fU5xkhAeiESKox/cSA5LXvS0fDmTlC08ZEXEM6vRA5oi+f2vXzR2R8/ZwjOIdrnm
SiMVB9++b701NnTtfp+ou4xO8RSsLnViFyLuZsoTOu9pBI8a7P8LpNVof8pLaxkW
EXU4tE11WGrfhu3EIZRCISfhq4IFKypxLweHWjQlwr3mhbInHYn9t+74LyYF3HyT
PE4nE8ydaAQFx7NWJYYCQZtUbxvlSldeNwOPKNvoUtXMzMFI+HegEFaWkSyJ93xq
Hbsr1vKaa2OpgBoLN+eN4pqcSTQy586fdP8l5e5iChtJenQ0CiDKVIZudzOMz8Ni
lLpRKJTX4NWEUyqeEt79Vo3SI4gq3z+Qr6kgk6EXs0afof03jlxkxAaKB+f0ihJh
iPxGXof42eYv7Nf98VGRw6EOdaOh+e0xxL2KDZD1gw4Ve726Oa5eBKLlxukHwab8
T0M8xzeRqSJM4n2S/nFXVnnnjMGJLThZSJyqzUPpvKJT+AGp2yWlaPWpnj7B9D72
MlWEsN7H07i8OJIyul+JtfARrEAMuL7PhFRtWB0VR2egFaMjCul3Fi2m5EmQZF6M
78GZtpxCVrt9MuQr7LVovQ3CL9lkLk77Jq+QNd0Ds9OP9i2flw2xrZJNxqLm0vW/
BM5s0ErJvITFTWkrv0dU4WLR3Pl/bm2EYV3vwinx2PyeRbV7Cr3LNpyrRdGgW+CS
7z0sLPZiuhmOCEgXO2FKlEzBaC6dcUSSnZCqKLfox9Dv5kVMlSl1SCNs8UZU++Oq
D8boECor4Amn84UO+2mxrtA11nnfZnErTJ5BJP67arIN/JhVahOAeLlweYBtto8B
4J2sWdPNrgsJ6WaJFmTefeMS0Fcl3clPmRLbrJLXHHRkkVXkKTdkS5ML7V3aOrJE
RFzbYrINBYTwG3UL8ZmPoIVodQMKbP/UGBQQzpb5gMqua51RC0Fk/L7jSzjuAE12
ef+j3KdRC0YnOUsGwpH4OmZxupgViQQ9mqu1hs965m5LvjA37/2PEpF9g3CXU382
yS4hTPZ5IlN4xObj7bJxmWVGPRFMxxoGBwWRBuCFdvbNChC8uzRi3TMNCksgePYb
S9xfQuLBkCj/I7iLV4aiyFRtSNW7qg5U+AeqUu1rxFSDg3OH5V6TIw+hJzNz0zRW
XTimeuyduj1hxyCwtt5SEBDA3Z11/+vI5btab+ViyftWocFEZXoqdQvdiRW5b9OU
yTjveTxgPykrsQdr92quECDL5+Lopa5NPHQfCqVNNUqsVpRJ0LBCsgsqAVzKmchR
VF7WjwGiiaL0Rj/BeYYTjdeutkbu+gdqomF/bM+Y0WDDZPwsFvnc11Y1o7nOjPE9
w6kq8Zx4c002kn2yipS0kzyASDmyG7Jcimg8KrDRMUDfnMLcqHKL2M5yv8I0xRrh
GQOONBpSfqYRmmfxWIJDqtZ4X4IAyOj92D3QupAFcd2je/E/cE/gsMf78IAOG1c6
WgLBqymv51QW72EcQEODz+Ew4DFeQaIkWhyH9Rs/JwUO8ht+PUNUu/ADiQ+jUygx
iHA3HLt0Cg/xhxIBsUE0fV8+PjuGxELG0TXseXg/Qf7HSbNm3Ef/sLkGZ+T8SoZm
m3YZ1LlryNk+WCZk+rdRl4DdopWR+oGLWO+yNrcOVNr864vuT2C8NSFEeLWrwt/v
638ZyXk0VW7PA4sZlqOiq8ivLSSIykU4Bi3a4LUUXTe/suEJj9YoNNMFqrEpLyc1
17jzeMWSm30dHaqfqKrLGj5NJzZkSBj8/mS4rE5nbPk+sMTP7ZWozJ49MZdwE3oS
M3IWFdus6Zcwt/yUP9lRHFY1U8UbyHfOsHprQMiWD+HaBYd0joHJdKMD/Wllv98D
4oheIz996s5Dk0h6QxibVeLdbwShfCFHxjbm0p7s2s28jNQLfxxc7J2LooMuHCBO
RVpLnCEIFmAPxcfBxa7GZ8fJmEsZOjHwP44AuawaSL52zpwF5dpStkdOTcivExzg
ui2OQYCRjRUdQbm2NS1bykA18HRA7W6H2Ah7qM0II7uUiS8WoqcaM5EHei9Lnhpu
kMFpjvTS4SdLAVIcxOTxvYVC2wgeauPrC68K16FNzbpH0QBeWIbMXB6hu+ab8u/y
NrJfj2ulvgSBHyIelOHWMNQwEs9E6v8nu9irBBazvCANJOTknjPmSW/mCLXAoHfR
VajRDLjXRSKtKb3fDuqYbQVldHRMYZpI4YOnazOPO7zVlB+mEb1S/5znxVCZcKln
J2yw2UPVWTwq6RpYhVo3pwr/7EIWYFlPEo+UI8Dhq5BzL3IHvkrENNCLeqDOT/yB
UTyfzj007X8mo5QlI1vDgak/uwfSMQSvcu1PiVUwKenVyjJ34vAkhvIvyhqSeP2n
Qy5y4GKEkxwe/Ho+fzr/dwXoloG4dtYR60NNbnyaCvbbiXABMWRgknp87gWkRiLo
AT1Njq7yS6CsUh6m6W5gqlvV9znOeYbbV1yb5zF9Cvle0UcWgByRPTfSOt+yhR8q
+zky3kE1NTaHT4ZyLLR0UYeLW7IM7LGe3KIvQN6DqTl3kC16mPRq7jD6a9aZLleo
HDGhfMD0+P/kqvBzWHiv+X7GU9+yozyLSstZxeFuhhplAbvbLfx/CpiMCHM2tLec
lhAywjLSARKtWexeN5KMt0h0AJZnTaJh3AZZtn+luA72VNNkg4BOWld8HUHwj10F
f9BXyUDyOgXjRdbmsqNFbr8JW0T9/SLqrHZL9zrpqx3UnEBogTHcfcX6qY18H+yQ
9Mr6D5MGCBpD39wp494cWHcVkCiS5LXe9LdspG5XFMMtmHeIvPS1l15CAjqnZ/TG
4i3WJmJT/u/WrlPi/SdccNOrekOoDNI4BteOTTDA2K9GmCeyy5xZywj6bxA+OG35
XwDDbjTmvWo+fvrBYhZIQb+8y31ak9LJ7SVquBs0Tp5ubtPkJhxBw8O+3v5MzKKE
e16DjdkzxCK2AEwafcKP5pslwixlAVZhm0DnfKvgoYxulnAOMwhdSKuqnnmLvM9E
r3r1S8zuyr6u66yl7uA8BMoBFZp1XZEWE8yZOxno4SfsLKvSN7N5GU76ts5WqAQl
3HoU/hKQPfVe3qJ6AI5OJNVtvhh3FVdGTtaOYc1AKzgAd/DU1jnOPE8WMfwgHTUM
j8jkQaSTU3Mpr44P7PcL5DXOzY1zEwTQlfsT5R1d12iPLVA5VrlGQDY+DfufGZzt
lCo+wELNPHhSKfOmvWbkbNox0vUNDDQbnc9SkR96+lU1Dww+KiC4tMVbbQOrytqq
FxxumJDt0fjGxOJ5sv+tj6xxd5lVqsp1HTNj6Qu57/Etz3EDNFoV4f/hG3dtkBO4
kkFDd4h8GJ8E7wrSateE/UmT/FSw/6argAAo3fd+yDTYTIUmWSxc9yasazoDv8RC
Tty1j2/QiXwvwtptRJphKh/b3LwlbQrR45Tun7SmI6gkFTJsszBVnwtZyllFllZG
NtbQo8FmSTEMywmdJXqNJceaF2Ep5tmFsnTPDDvMoHboWoz3XzRj0ScMjEJBWEI/
hIt6uJ5dh5ygXmtsoT9t4jAHmgWfVVgp6hqPWF6KmA9gqWsIwxO1cpzcYUUmflhi
3/cIAGWZKybm5++EhrZbfyJS8mUpFw/kcmR97b72N2+BQ5Ou58zYGUbhkQM16PNh
iPJNbAX1YZEp08YeYi0dhghTLBkrNsw/s7S7qT3MsGLl5/jH2eDZFe9+inav49pr
6Ce4U05IYRaQtWjhePAey+ERCMeF/DSoBGfmVxMkAjfn2hlaIDUIVQ7NsaHEBz5M
y68qhxbVTLFj4CmWpOjwoG6f2o6bLUqKIoX/yh08h8kjH/7F7TD3iAleolVwHR4w
5AHeIpWOK46ELrGAV8tkQDY+OqKX/Xb3mxb57QLp1rGN0YeF+QRJ8WePE8mZmdY6
Rv67Xw7KsN2aMIwia7zVYf/FJzxRsMaSnHeZXN3OMuSPQUufZUQAfKes9sd+Urb7
LtF6A3mq9iOALsDB+78frA6era5heBGli1/VXljp0R8SteKfXsGYtgNRHwktilIG
16sE+wVMOjsjfLImLo+ePesgryLgB9kTBHv82vD3Gw99xguwrDP5Feu+wj1Dp1Gc
EAmcCchvqBeGNk6vaJhH4nUn8JYWdG/1IAqwjbL/vARwrDW8Nvz0QqiNFa7eQDsj
oOuMzhwOgtXAIG59YaZIZ3dV/myTKpJJ+QG685I090wlpoE7k0qRXXmSUZey+VEb
CzCH/IVm19AbKVKKv3myAmwq5JUWmhPHKPCENUe/ThMZGi07cDQeWKiOkyPMTxWy
vGPkbqAwwbbRNR05dSgVL3ICOdr1ByMjbGrAnqOgdcEbhcb25YTGBDm6ZL0IIWBk
1CdarCymduz4qKQYGeQCDYxaWe3YTpFnKPXNVsrNIXi2tRKbONHVYwarxcl/L8C2
FL1dP06gfH2QU2NNrrN/+VhTrXcjLCrTheiwdrmQ20Gax7L33OgqdfYn84mbKco8
ggY782NXD11MebYFdWT6wbksK7sAcXuGqVCXANf3fbz49aCYhPzU0I861os3iN8d
bxZu/udWTw5yLwo9MC1RToXVmDlo3jZiScRs6s4FIGLYidKrBY+HofY/D7eZQscT
PUhKsX8a/bvnUzYW1cjjgpne1OdZPorbB/BysJeH+IN4CezewAn2CLnf90DXNG/u
kHnWpk0NzACdDALrKeIG4lJBEtMF/rOYPtIpXy2tJuqhMI/mZNO2OL6ODdXgFCvk
eujtN5W7AeBPKgKIuOK1ErvUL/vx6N2tQbsYseQ6vRyTgkMhCP0DqjZPYUfHEG89
l4nD6ZyAH0W48A+/tEuAlgivRBA2nePAvcK3ylw9ML/gx+YoArPdngK0W+xy9fva
sScAPaycOC38haYm6fzmHE9Sh/ijjTI9IohGQOHFG+mIhblKZpqUgLgbqDYPLQ4S
mS9AsSz/JjLqV8PFvvj0VIhuLckOZydmKdDGugVEP8QU1FDaaXcRZgQckIbtPkMR
mQ3JKmkrl/j8WDG394rA4GLHN4PoeX4F/y4zCNjlsodyRLo1Ac1A/+R+iqfuumSQ
gHylwycUQfka1/t1EyLPibASeT1ucl6Spn2bC4ApkcyaCtFLaqQoCADbhu10iJka
11n9F768vhUBMZzXlQkvOhEGFC5nRRSMI3zVnUtXie9N2CLHOUeZ96Cstrk2jOGW
dTRe8xBU7l22UjdYrohk1M7aLkCFu7wfujgi/48w3yAB4S3SlKrLRqgNzQwN2+DT
E9eqmKxE5MF3H7hG2f/Rk6eHn9G96MhzIe97H2jCoQr4Jf+O44bIbT2tMpqLBBWS
oUYvv5hTac/vxD4sbYlhXwIpmOnvS4ql51HBZ5QDVFpf/ucy2h4PbCOnKAgXCedA
PFfKgDCf+csD1ij+ijBnXEav8EPDXr+k0YmxQ5nw6wCdVoW4xh3xNuI0Tkg4gXTq
MRK3od12OOH4vJu8OEtq3wYhDs1697B9bGcgR2HT+YPsOIgJcQdeG1g/BELECXwS
w0GyB0WTaRFLwXAiWMNCSrDFLtpHG/vGpTXpfoUkfvSdXawuMB/aUSpMabsYId0D
3Y/IOwon4ATThhgOE0ejZ/VRFtp8e7BRsyED5phr5N/k6+HWYk19+jkuNHF8Uy6U
x+ZEFq0b20iwFADS7ylfbe7Kwb60qd9+OK7bVUywQY57s1GeFYM+lNNT4+cHcGqd
oamvhUVuB88ddIrfWHBqdKxMtmtsbTQPuzSA1HnKjQzUTx0X+VsZGw5dJinrKVvK
hGkRMl+/V5VKmCsnPM5WVRKQxeUob2eu2OlJwBu8Z1ZtFAaj2kbhumFJZCpXOWoq
B536HAf2GuPISPsSzCI7RNxgSDqWXiYsfIjRiZXyqJ8FByN5Jl31RsVI5jusLDnX
18g0y3YOeqK0i2KBUYRwmqBMlNA5lGJn6lXYB3AYDlQRZ6kn2NLnPUm5YadKttXg
g8hW7ksfaRy6X105FPfLHxJEVCwFbuAT4xmudDooy2EhadSunFKo1mCZKm1R2mBI
YuUI7FXDpUqPuXM1kAsWLF/ZN/92TODI+q412CpMQ8bfd8zR6H3RuFtl5jsVAjSb
E948KhjNC1TBtaq0Z4sH8t1DdlYDKErE/JbI2/Dtx+3zNVwwVLOulTwMkVPVNWqS
mDdrQY2yZsYWaDeSwSDUGeNtFmOpAtKYFd4YSIS7tyMjL0foRVaVRMTdOSsW9QYw
oOkchQcRZ3i/exf/0qSWyEmhPVlJkhJeX/B+Hid+3dmqe2I3j2NgsYKV2sGvl9EZ
2z4h0igr9HpoLD+G9FQc7W0xzCN8kxPRB1oNFA8kEo3x7XAXaJzisGPY7uQa5ZZt
6Dbt03dYA8wgv5N2n7NfAaUqfAeVUGZrG0FFQ+Ax41yU6wIUXVmEZIUXAzr8bl5x
/AHCu2lOEbFEH8vKzGweN9jqfp0XN1pL+qkDpbgxTuO0MCTMyX3DpXznsZkVR2fX
9u7kxkFIQSTe7q2U2lj6FOC1XnoKjIeBogCbLKAtX0hwsW+GvySYHeO73H5MNPf9
JRV3uHhlVFp+j7n0OZf05hz0/m8JdIq4XCSLJWp1Pb0cJ+/Ed+srPZwGNz3Njkiz
2zDzmQcIaX3/ZwkKIqO7+FpY401gGHMz6eC2xP3qaJ4wlioPF7nTQ6Gwm9gkINEk
6hX4HOd4EALScdhRLQM9JBMEMO3QwDJYuWT3vojssHQgNHnhESq+s9jdI2c1QOyf
edvVa8gz3ErWoHHyMOBDUMcNLtoVmt5psa3EMmKW4qFVcIi4Tq50W1U08tA3kt6i
xYBrwWhXUvyMdE2v6jEJTCf0nQWR4BnNbiKizCh101K9slvZXnXbBAG4XmPYYfTn
jEbd2yxUoTiQnceZZRtjeb4QeIIo1jXlONO+wLapDM8bbGTQvRB3IawFTqu01ZX+
r71iwIVhMnie+1lYq1p9wF/w9vbPW/fChG4cUfPJVN7N25u/7MGF9Gk3RL3KVAic
Iixa85oJPMgXGjij7o8fuUqbMORRHlQLNwNvGOMO0gRCI+7Fyd71n3Aj5dzSdoYG
9IGiXub3X4qokEExH87dNvOw6m07m2xsBWxqVS8x4Nn5eBWbz081s6xj+ytM6lSy
RusjQ8f9w06HqkCU9Y+Oy3f0lhcQLG53pGsrjFWNbTnnRzjK18gSXr0lAxKCWWX3
40SP2ysw8BLSORbLo7egs+3LigiGIMhIOA0XkztoPRH6dgg8PQ0J8TdH/6AmEPz3
9ZbEW0BhnrhBL9S39OhcHrq/mdTKUqxx6UmGRtPMsddHnaqF43uhZZPfh6tNrdPr
l9eLb3dlGT25AB6+78Yb4Ks7W/si9LEYegoNmgqUPCT9v6pZiLTTOeI0qz8wM+jX
0hPeDWs4ujeo4SKqlQRr4A==
`protect END_PROTECTED
