`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xxr59Ph4F111LLxuDu1Hpvg0eUslYFWf2iaSRp0qxpbeyd68GQWV/A+6jTZlnbF3
ROp8XcOcx908b841KtGGPeNx5lWfnOkwUZw+bxhBolkomLvQgn7MBVrJj7F9dKao
b0t+smxcT6nJKNaNkL40DFt6PLVclGSZENaGeKx5JdfgeYzx6Y/2Mx5E/5NNnoHj
IgYrayzB/d0MI0LT4kcKOT8R6SXv5FZfuH/jlICvVDXXRxCWzHz0wXakesyeKUbc
zxYDqJ4EW9j0b66Bq4q8G+ICs5ME014b78U7AQomzfVQwwRySFqxpj25JS/soHik
Ydk1DiwsP96qK9Dm3LQsD/wsJRnzNprVTBQwPwk5chbl0KIYUaN3wdrLxQrsH0LT
5985ZBSge84rDsK9ihh2f8g6zzAWWdXkevf76WGDt3ez0jDl9KnT4ugUiZDIpUg1
NvqcWStgZYEVtjkPgOVHb8ZDMySb+/vXWjlljbRmRk+xbY7jyPI6h+DSjh4XCOq0
qIn7xuPZMIOGlcgobkHGQd1CrnQ2/BJFZcxeDJQ5WDo0eaTd9zc6Ez8U2pCW0121
+XZ0kZCvsfs4TcNZEqdZSvDfJO+cMRpK6YM3eeZZGVim2idELQ++Oa+x934cPGNH
5e3juZRTB1MmUlX9s34pYRJbRbs/0vMqXRmxc+7FFsHvOqoj95t74jXjmJDGi1R3
`protect END_PROTECTED
