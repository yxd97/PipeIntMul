`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8I8d1/2MsdB/wdbxNwfS5Xt+iK6XMhZ/UaP1ywuds3Lj5aRpMdLscJdg9z753R5K
2OKffJjD8J2a9bTf2iiMfQNMyoF0FJNIslOWG0T2Juxsj77B5st7zsn5607BkBFN
Yqn3kvBuCmHm1S6vKFqhsboHrGo8rwaBscpjYBHEF9D3HFSpMjYUPHpe4AwqgvpM
jegQIDZxTMSyo84RbnJFeSDm2eCrhgYERpRQU3J1Hty0LFIpWtQeF59mhld2qMyp
8VUfkB7wDWouTzsBeVRNORZivMsFkosHNiSqhlneZ76HHWNH7zWEhnaN22Stn+vm
WvkChkw2AsOQCFM3mz7tcZ1wk5wn4vwUDS+bWmNQlQz2g4XbMeTyqxDzfw1lxDgf
wmdi7nu2sLcUxCn/PNDCf6TC9Qgi1A5lZsyXBztuLCcvVL+MwmyNwz+NQ54YKosO
5LLuUjsf1wQEfLF5Us7/79jW2U8FjbS6i3gd4Zb0zxO5q4snqE7ORfhbpiMFtO/v
iohgXtlu8313wAQo+qJXGOOMfZeSTm4ZJN8PTmyj1nhQQP402SH9ya+yj/WcmVNq
DsBwLRpAfq9uCfzgiMojUVssziL5MlyGQktsy7BZcHgXk1bEy8L6UAp3RC/rqEbk
/u++YAk65OHe8ZOi58iU49bGqRHEn7QIdxGE9WoQSqmUvHe2gAU0r0f2N2KcBk/z
TRhNTRG8Ej9tyn4kS5LjBdc3pc0btwocOpYIUX/mr8/pchVbBijkPeUw0Evnq02J
b3KAp7tX3cQ4H54LtQVTBvsLpSF6jyNF4W2A7pOCKA010qQCD00MGJpwBQM8i3TS
+ZYvYxgsLCGfexZVwykEKAHlHzLdCFQtON15rqGqiGNPT7/x9FYX0rr+bdtkAk0N
IKc7pRqNVzhQfkhHrlHF+i+lcHHowd4nPa0sjhbKAndpSQhJT6u/mOzsQSK75PAH
T9xZqhZZfCaqCdO8OiOR7AMhLes7pbBYP8blsSJDh93UEhpPPISPRiPcXlyFOn7M
NRfyVeQq06tuPP3ga2cqyqo0glp0mpaDVMk7MG7lLkk8LdelIz/5Paepkn5gvkO0
H0nmA0ZmPFyPOzM9i7ECJQ==
`protect END_PROTECTED
