`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/t+OUKPLlJBm4Jlkn9CyW9sRZWPkxpbO3OXwWFhcs+mgtQXtB8n3vz2nRku8flFs
KZLbjb1fI+xdVaRMOlnb3jOzYyzTsSfUaob3wA1ElmOLPjGgCSl19++kKDKogiEh
mWge4sJBFB8GQ2moSwsggL9F1EWxCz6mkcqTfLvhQInhPp/a+L+q3VgxcBwXu4rY
SH0YNKNxobupIUoSKkeVOtWA2O+y4A/2G/ZCNF0zEJaQneC6ll1Qf1ZiVF+Ah4di
Y7VVTCTuiU4OOXIOYUyNUbWRH7eoH78HY+HrSOz5hdJpgwGgmVk11PUMw15BsfVd
udOs0dzJhSCQkcx6GEW3ulPuhpqc/asmrBwtm3Kk7qcNCRrnCWyw1wY8h93e/JVw
4hqbJNqrIv+uRB3pk+OaARnjTx6lZmK7/NgipuTeyDKEahz3nlcAh+SE0G2Ti/hy
xkiIqaT14ilrrolTf2d3sfJzX/e89r3oEA0hDjy9xNBmnLVqLNudZ4cxfJCGNaky
GZCNwkWoKcWl+Fs3ZEC8dHmWpR0VVaPt7z6WkyvEL0k1eB9XkhSewY6hCdTJ9EUI
C5QW/OkFSjg8slh0oKxy5TpyGaAj3ivNixKQClnFZ80X9VZNCKxne7Ka+M2UvmO+
ejWIeWK/MFE7h5z4gfAtCZl1rQPYPqO1n8DO4ZbLgSJa9TWP70pK4JJ4Y0EgfISJ
66toMYHia0ysCrHAT4lZbYhYHQIDBjhKSJwz7LEhgRee4TIhV5suTgAg6f+XjnDl
P0D4BPEkJZ4jXyt3xiO8yM7XvjHc+psFFKaOaDUZFJZr2DR+nmoURU5RfuVkY93N
iIahIigokmx3nVtXPJV82apfmpIy+OdS6Hcd5u6rE3zunf5KHM+rnzAvFhe42Tqu
o1QuQ79lCDugQwNUPvKE5HzZS9f5xbybBz1bpcyjxItTSTQPUR16LfnQ1sxhSto8
OxIivghrN0J/V0nY/WcQCP0UgaumgrlHHpplXYziqlLZOgr+GQiT1d82hfXq94xU
KlP3b0Qn3KwazM4GUMEJ9cloWEfpkLCvbjlDF1oObxI3MWxKGskhamlrukk2yX/L
T7VyUtHRxlM17GB0qfMgtdVmwzhozxaHhIOd3zAIpbW301z1HdznSpmMOrJs6AlR
4HkjJDVV355mzQ9ghSPiZP44x9K79iuZ3eG81fNecIMXwo5sLrjmOjLKej8650mn
L0/4i6Rr3ncavliGWjr00NvlOhPsf2PRmNf+aG4JCwiN77mdmRnIrFAPwIQmeDbV
dadro5ebTGCRzekV0r3kuEvqLdPjqbIkUhc0mv4m7mdC4m8fn9083FvIh7prf+1k
zAKu+SWiVDPVOCHWrEAaDa5YJNu02zxSE1PrqEF6WZXlRuTTSNC3F5LJZ/zR9pi4
JT0gF7pc+6qIDLtl4Y78HXhiq0LIs2mD1jYJhT9v4OO9Npo1fC2KD3XitrLNKgc5
l1tlE/8LBud+w4thwVqyDyeb0QWq8P7GEOPQI4CS8GJAWngY1/rD5HW85xLxGX9v
Wik4BxAfOfa7oMNL0pV43O6JI+67ThThVrpAAHH1Dria3deKfL2/IZq8S2NZ4Bbi
hdmA0NiB5M85Fi+kFX9r8agTlAt7wJGLVGC+xfueb1H6kO/4LDbQ+9ieWnz/ohmR
vv5i9g+7WX3CQVz3fhlkaQsvsbDFu5xIvc0fWK7/LVEKenDjZLQGgOyuQoyFCnVT
nZ3yRiOK9MLBpJUSgJkDOzWTJLTQwwaIIt3KqBscUkb0EERuwH8uJ7LV5SqXngFC
Hc8eKFiqoya/XR//p4iXDf/mAaUuiFXfWwYVOGiTwLmnIhRl8tQpNKJxyiqOIMJR
B9iNVB4msrs9C+35UagFtl7tUsG5JzL1QTtqVqQRlk5yPwmpEgKbIAqL3USr9InV
x/lnwjxODzNnIS6A3rQLU3BpFKGBl52MMp+wypVyqmz1Tpx7kF5R+9iTcVWzQbjg
VKjWkisdzP3s49unbwuEE1YXQX5zTtuWxyRAQPviGOSYSLSjFlzkl1EM/vOxHRQf
sbtpJyTPp76+5qaOLEHKXVRDRIZLPAMppKHsBDejwv6YY92e5Npk/ca9sDJ/6UsH
s459cQ4DjVIf6rcxcucnBqmuJXTqfJ7BlqnQ0SzCK4AtkGKbu9kE2hjs+7oqpkbw
l6/FAElKkk/cnI95/sZjRMT8h5DtVkE8R4wm11XErFO0Q47U9vtim4Se/rH3400N
M71IeyPIl0G0Bl+UivwYKVx4IwV4r+yiKJFYwwa5zdfQdSSjoV05r4co219IJCLf
yGFjyq2e/9x6VSFAup/TzOCEfFx3ckU4aA1PXbuith+Nx71wXsq4cnAqMZdl/Dmg
rfIMp3AeWWN76bgdvDLBisoPUewDX7dfKwxAx/2An47kayX1xyYh06T9cVXfQQgm
P7MqS/N5Tvg/xoR2ufilILrsRX9eAGt+LrBx1KvQ9z3ZYUqWsR36iDuuT1fUlEed
zuAr+L85LUjugQDo6AExgLPmPHRvPOx1cG94slbe9W/bAUGONEEB4mmZhhi83Etn
6RHt2VhhqAwKVFz2QXOEAXH2XRI3SVgOaiVI4V8teGHkJ67ciyFm6+tZi64eJ7b0
TVFQILmMEIH5E/V2DDIy4v/feklINHv8vVK2HXkBeLj1QDYSRVut4RbP3WlkaTmN
8+4sA49TKVYpPEl3NXMhrlLrNkn1TICSiTAf4cIIF0H4DTd2iQS6PBBrG+oBmPz1
enHA1hKk8woeyOsYso0S84k0fd5OQ8bM+CQTDmoEGF9hp8vKPblSnK+tczzSAnE6
89I5HI/FqCCjXy3IxHMEjbu9iFT0azlBgcyiiBCzxZsDg55YvRFqOJYAqdlB9xSg
kNini68joNy2TUz8RXhg1IyB5Ct3/dczLyXPWsN7zEuUzKVGIKJZPKwmgWckA/LU
/cAJ5QbX1oZvyEpZBzGNM+7ocz2nL/Q040EDDyRVNCtnFoLaJuEgba1/rodooI/7
DHw9JkUSeNDQ9JutJq0uGYvaJO9lh38lQw2irQ3/Ku6ZXXz1LsgzpORCT6wRLslA
mr0QN+B7DA/9ChdmwFLevzdPf36doxdKvO7UNC+geg2FdBL/SusbqUtPy2r7t3nE
Ha2+d+1634oc4xLQCf9TWXUITUM9BakuEjUfpxkBPzW3ZhEjN7wfrWOxrYz8dYcl
FIj9DwcAZnSt9qDgbzV9XRH/fP+VQp1Q/gkNuuKbg6wXvc1TFI246l1UoNAe0jox
GzluM6bOlbjI041LMbpZ7YwWdalbCGErn7xBmoqdW4JVv82w2/HBto9bgKpvbArT
RawfF24SzycK9kDaBbTXMaNHMthRTGsueT1dXdoWZDNhxLGqQl/RNNZmCd0Cavrh
jB956AqzuPXnBDQOtGtHU2r82ssIe2U9nIjrTwZTr8HeCE/cmWXC3zEw0guP1zlL
5O+yFBEVSyJ2XkOSTnIvr3fgTw2Y4+U4+vEwTQISEWi56YaXwqAUaw54F/WmnVay
T1Nn1UboifMpUVHfnbtC1VriOg+lsNRNxFDdcuCbvxhISacW7OrI7ibipKGEH0Cb
cPxDL+q6jjSTJ77slPWiApAoKohQmkeMI9vDwqFsdfCJGQA3TB2nOtLJmthfFW0b
cDJVD0whASLpLiHILR493FYNZGSjrpx98/Jjfew/7y+bof8+j/68G1Ec7IVMNxgp
YkWOr/lEhEXdgKrVH3sKU1bdBSQDJzWcPGTI24lEwBecj8pAr/szJwzVIkbMEYCK
9oHvEiOXgljrSQhCb6W6QELMZr4jB0MNdXtCakLOyZ4v2hIDMaVC3zGpJYRbcVIU
L4v60K7LUGkWyCJ1cq0rGNmnMxQYyk/9NlDDUkoq7e1fxkxR2ST1Y9SXwcf2Ln1R
RMI60RpoGPB1yZdxPj3DgkCl6VHhVyG/MxQfcBYg3bfJsKRBxorNx37jzqrWuPeP
SGxAUj7aBomCVgDLNoQWjHJxyaeUaDc0P8tww2WPoV5AIJZCjPnqpiXPKAQyfq8P
DF0swTKsETCe5ezMV7UlAr5LkGVxGnPRXqSbZcQ/gDgRM2pC13oQsfJFU/nExPCk
fhVEtHk5SHKuN/r1/1o3Hzw/3U6UELlUw1/bJsSlsqXS+LwP25/hBiVrLd/vWItf
bfxZMvWpsJ8LuxfYMxNgi2R6Q4LqFHkWt/ATPNZOirXfm0ZDJPsgZX3PN+H3wysX
2l+fZkpW/vxWK6TiJ4/mfpOE9Osps3a29PpRWpN/YOrlAhlQjkzofnuGSWXu5QD3
06elrIqQYwt+gNDcZ1BncqFM+qaXexKIjaBJOcY1gq1seJIiNEhUMX4k+fHZoAeN
JYJPQSE1W8x66nKutsCgi1Nm2f3JgXI6fz8DwbQAeIeRVVQHPmRqwqWNrav9EgSO
H1MLCDXbyX62sUctRwmtW186EYh8jlSY6PKFhf3KK5nWy5I3Xf5JSPVmGi1Hg1C4
OetM7Cxj4bkIor89u+fj6USNKI3n5JK168PIijPTeuPpRHMxF9Vz/lBLGpQriXpH
GcjKkohmppb6RgJ8E3j45Yvf3I1A4UpwlgZL1nSYC+y/XW5CesMss5aJhhjA+M9P
sKpU8LbF+vTeETuHefUh9sofyRxrlTaew+f8VeeSxeqcRG2uIH+cdXY3XfVYn22B
ChJe6eFm5VtZj3fy/GKdA2xmSl9sS1qZz8ESZWMzeI/tEiMiRITD41+GyGpgXj53
tXfQaUNrJInAq3UFjUO425GUJzPkVTzXPsA0ZNee6/DCfHDQnqFHbaEgMp0h1SVn
7bbMu4E6dvmCMbz/ZnAC06kVOJHWtOycmwE05CwhM9frDS8V7/3iFcNXkSiuiQJZ
rCC7YHS3ch666sBJTxOMd6Lj6qTxCXEYSwO/J+7L/cBRBYIcYGCpEcDyCN16QcOY
lMW2Ax93PBNSvt+R2JBh9Nnq4dXB4YTN/Ue7HKGldxttMRMK0quAZ2qY2BcHcBk8
SZIvN6kh0rFTbVMVignAy35iS5NhNx4KQablU91fVbg8yq6V3jcyNiw13gdBkUyf
q6qunQz+1+RWwCHOAvO563iyZTJBtSbT2cN3PKF4Rt1c1M9t/k9pFoz8tjus5eyj
Cb6rZw/8t5oIyIrTF66OWMIgXHfbtpRswI8SUj90QfkjTRxB6Ifaki9FkKTCWsE0
XGsqYPtEIUs5ajmEhxrAYMW40WH1Yyv8pGN6FO+2hGKdUdw1puMTf3nKwQVkUxRl
b266WKI0vppFmtUxNQls6BCG5M3GvKhYHtHtx5l5J3gHgdNiKd9sImA3PK2nxUJS
3e9IkWgacgJ9pWjnj1e58bkdiEBMCzo+tgWfUP+JRz3VQrci/6rlvdbV9ojS6SGS
q8S2ShW6+f2f35jSelZR1SC0mAYkaV/7RxepJTIjxfnmjZqFxJbcrpDOJsKNrsNa
JC25amgEtFlFhzvA21XqzWLKCyPdFStPNjxX371/tV5Hirz4msvwHhYcAhs7Vgfn
JBKWYKjP+PnfC1Ise0TyBrmtmCHYwA9nb9rn6DaEvLkl5jIDs5QCgIKaT4Tw5gL2
BtQ5xKi4GVtllnADtQLY6b94tEBwKqXWBYC0yklMVqMoEFJa2MTpQtN6v3jvYqc+
9ae3MtCh1liY830rg6a4exr2v9EcbGIq6n6VEld5kkumZi/5Dwuo3ibqrVYclHUS
QdoGXoVxXxz6EuEFyYKTIdfXCEfklcCfdNvxyUbcweiqR1PmEkSA6g8Agw8SkUd1
S8Am67NYbv4EpFt9HxDrbgqaCX6w8rgzRXIjrxP3jqbJp246tDlF4/WjA0vRUGja
/HbU2ofhkSrpBWSeHuAwkwat1kndRsUnp1rW5Ln4FYu2oal9+2nqraYRJJavMJA9
9vhapRzVX6LZC2kLCp2Y2lxEbfy9Kc31oevPxrgHVdGPeBighfV6yDYQo/QpuJaN
/8Kx5waxc80Mw71RdMHpQJGfyFLahaMDiMMoxuxoX807naUYmCWvQJ07m2+RvYu/
S4oWLTgfhc6ZQLhA6bP0xFrqrYJ0LNyGE0i5sTgZcZpkj6YGkwQb0lsWR/ERHuQ0
QGjnTuyRV/qjc4MYXlUdcdSeoCUPuBsOpSvt90XqLEPyK41N6ifSxJPeVCvJ2pZI
/1hZRs2yHYEsDschIFwE9aTeTfQI1X5cCnB8lNqlxLPZqWd9spuQCsVqZ+MOAE59
iFC8aGjRPaxfdmy4L6o/OcqBi+PrsE2QrPgOme0bIL4CdJBCcT0eKlOO5HAkkXrg
QvH0UyOEcc3enzWY32gJlbQHKKOutDO5joJHlBTL8b5/6QPxZfNh9PMANiQEOcRB
Etb/x5/0/NOvAeCkRMCeQhjpodyVz/6fbhqgVTbS75oSjJstD0yG9mSXb+kXI9b2
S2VchR8EevYJm6jYI9zOLVGwJszG5E3/nF5AWvUPkUwc9X6WFXjs1JwF1yZvo1Sx
EGEvMWaKXeqEYOBHCCTPWluudwOGCI5LtL6hzjwgJVyuaftVsUFwr4Pblzplg/Ew
JFJ9tYeLB3ZZzQZ3I8rzywKfZg49w4t/cTMihyIDQVwd4gF3o8Gl3TlvTOSrR9/G
qKySBlC7RC6A6/bgxQZsZ+6ZxMm+0btm408DD++qaHEhxcyLMqm83GEbbzv0RmtL
UGh7vieB7FYtNsHofwxU+CEaB+o8+5WLwbWL1hOcUYsJZYQqBZW3dkFWofZXdTvE
L+5jL/QtkunJFvJEOArJ60+F9N97aBcZ/fYKttaM8w7S2y+MdDJrLGeqwisFoXoo
p0ALwtlcCKGP/Km4AnOw6ptBqRWKFD36j3FNpHeYsGaqYpAr5t5twslwkALN8SwV
9QdQoLkYgRVYC/rLtin3kciMVhO1SeiChortM9FtwmQx30tmV62JBD7IWUhuWWIl
mGrDXo3BWPlBtBX7cJNQ5C60tADWm541aHFC9ag6krZPShchypXSkhGxSAQyeILG
Kv+QGml1P0BAcjZf+Kb0swdCRhOmT/FvORU1jY/R2yHiK07pFXtfT7rh4vUjnc4l
0Ixn8JVmCO+rggGy2/Ks/3X8K2jwwW9vRgFAAUL+YulWtu+FcWsbcUpynhGUug9y
UCr48n9UMdbazv499L0f6XUWQU6dFFaZPmYLTnB6z2Y4CzmdVBqWnQyP33KkoVc/
GTVvZQ+XLRkY/TVYtpQRDQvyweJYnVd4mK9NmlPxtQK/LIIAGZseIA821HLUcWI5
BaQexPgIWsP3ss7O+hYOTC6ZGy0Qul2Oes7HkmKN3HILu38vaOig5TkjOXJPg4i8
b5ALTsoNRyb9hTARG17MK7YVYOcWJsK1tXk9hnuABcWO4UsknAXVVMBnVRLHSMjN
qeCzqceBDD2KAJBXiFNq/wVtk0V9hcQyw3iwsDofrUoZrP25/nrfURIXyiZkTFLh
JA4/R/JAkDhhiryUuAnDFCkHOcn0sVk5Zqm1WmK6dvRZ1EuDOES7A9qZeAvOGns0
QqvJGOK+uQHk4rynQeFD4G/itYAbRL/yT+wts/DaifFXoxCZXq/WFbBzyPwUxrMq
twlyXfSuXNwjCRiBg0Dbr34BIdDndUimRlh308ORjiZVRaeyALJHy4BIl8TakJD9
qKcXxEpFIYGs027KUkFZo5JQibPSmSG1zc64MP/kvEQOB0w48l+u4z0w0GexxgmR
V4mOkluBquiPMmdgqR41zwvTis8J102u1ChDzHLndPo89rmcFnfrQz0j9TOKYVUq
C+DY/RYSH+xQ7xb2QTOG3McfmmdE65JGXx8j2KFkdNY453N48thjy6H0i7P7qoYy
Y6/iqfADL+AE2U28bHCJdwOqugVnAT+9khM18tj60qx9QIBLpuwUBIFKCRhoL7M6
VRz+rwoVztyfjPCCJkU3DvN82TbQ/aYGxPzLXVeT68SqzGEp/WQaLYycl+u1mxuI
EcgfMdWNohToFvVslIDBIGnxMjKgK5L0OitVTbi9W1TFHXkY8J95fTe0rCSdVArC
z1RTy2n712eqSkkAsNiuDklmTBhdReXEzT6Vgt8a24zIHl7MYyIJ6KvsSGUdLQ/N
HglyB/JbSeczu8MT4AHLAT5tplHZIlOkNnbILt8qVbqEZOCGHxiKxNwZF9BGt89D
VC6bBnWkNg2t8SkXwCoFSz2TTEcy8jLEYhBG4gxDLJzcy135M7v+n/d6TBCeK3Bx
vKIMA8TmKUntbHpZjozvecupUngHCSTImQKrBO+i3OqFOyCcL4FLLwgLn+65F9iU
RqnCF2wg48QB3f7TFwvZ+ub5IafzKTxCMMhFUNKqRU6tQJIOFzt0K//nUvqdyR8B
QRcZK8FvNxvUJPzgZcQj9SVvLBHKu8bDTe3OvJL6myxHt9JDLHu3CejJS3hUZMuQ
ROIFNDWQAckRkFnLQE90rhAIsy2YwLhopdGGJScBK0C9DZ3AyLsii416BM9KpF4/
KsY1zQEGe2gITVfhxKOE9Xp0b3Qm5PR0bjRssXXSB/rKgL2dSieI6L4OieXTooqL
eoH2kwAjVMnb4vG9SPJkfe7X8lcPAWImHVXv8Uo/sEH+d9szz+d7gby3+/WzdZ9q
jelHI8hTqGq7QAxQSW0tp0131rjUW22fp0sKAimJzRVw43ASil6nUkoYGDJfiMej
56nnec35t+7JAPDTbjpfYLlds9LlUZDefuxNcK+MX3rYLOpssFjgughzrHAyQN6P
tmESFqGSVYflJOmk34rR8Iu1Gb5F+SJqAObvvIhKY80yIbA9zX0MAmsKOKSbEG3V
H8x8W2aWdxNap/CnQFrG08a4F/NB9bYVpht0RRJVuOYKqFKHB1NQ9yPuMtFriNok
7oTftt3uBeT/L2uBJ6AviDpRuF8vzRaNBOqy97JcpfSQUbOkMDSrnG5IwMS8vcpq
9lJwbKPfZF4ENFicY4UDyCk9mmnPTjEIyY+B310Noo4tkuv1kGaogabWdl4AgAdv
b1zHRBw8bfNT1WQnyQEvh5NDZsdWrFqyoRBh0mN4mxj2XaE6jMIIxG3BqfrkK8eY
FE3v6nkLG04BoJ0iu2jXjv7mVxtLlvqqZa3jdh0d716iX3sVnO7nRvH6sToDhQX+
DGV2OkVXObEJ1R+LtmcbpNvIFOcXtLwQe/ohDn1FFrfT4KBULtDD401ezXZZmtyV
SQn4H8aV8YJklMzpSBo6mrrgWtLmNeAV3kiGHBi5IRw7oGy4DWP043ogHvtp8wWW
Vz4OZYN/W0BioDQ+y4kqLqOIW6+NVsHm1qYlFgAIANzTwdF6ddXwhIo/DO1W9A+k
eWkM2aO70WYYAk6J/9yDLlAMeRU/Abv4j5g8Z6GzkRreNfHaiSWtEgM9Pn5z5vtO
yD0buvj/S7Vb0a24OjxaAHIKu6dSPT1kPqPTklhU6Fn82mEiWQKF/R51Q7Du45EE
xpdNZ0/nTazECXV0SxJBCgD6azn1D5Y6/gwQwGjwYZsx2lq5c1ImprfjYb5pEPvd
VQ/7lptFkbunhrNR5kuBLeu/EstFSe9ZzO7yrF1MZt/BYg/08aFGcggpdLKotFtw
FIgmqrEEmgaWNGsQMC1onqRe0G2pSPDK7a9rl8NuupHkh6ep5L0jiEKAc42/EHso
jecYomc6HQf8nUSSXTpEbHuweG+XN8vSJu8K7eFe5I+ABU940TQyTy+1SOsP7lLT
PLRsSq4F4tI4O47bQkJxGc7rqvZ3j75VYTzPwFR3QpAqsv4xdvInkLn5KKIuuEqt
LU5NP+y5qPOxKATdUpuM5Sd9yFqjBAMcBaxlEbaiuMnqnyntqs+i1WFKsB0FY/+G
5ppOykdjLrKs9TPM4kLBByMmZQ/9hmmmazjLxWOnyuXhecLcFQn+2V3C/Hg6V344
Duz7ngn9I++z9SoIHwemNDwQB0lahOCr3aOFb8jVpgdg1yrKE5PDUnIA1aDuAD9K
ZWEiODT4RmOS27hMcLm3FQCvBHsOGcO0HCP6+8hMpn3c2Qnp1t9luw9xrOFusO9I
DJtjpJ/YuwnsknLmsVhCsUWFsa7OFXkgFlXpz4cdD8Q2jlbnyGmVogKWsc/1s5lR
BKZFuBW0vz4gMKc4B4pteNntD/RkyIm7pLqjDNmQ4ui1lTaOICgnMNrd5EZmYy6h
01A1Hxj2phXdlXC1d25Nnpqza3L5Cc/nLuQ7bGoCI5UXvnj9u9Q5aXBccHe8lcJK
f5LDu7hZ0O79v2be/v2uaVgWvZHsXB+tMsWJJO0rmNhGKDJINdk/ei7BHHkJuJpC
I/fKGz78QQTwYpxBcOvyTlMWI8NGa6tVVXUrtQFrGPgklO0BmU9W2ejX8g2n1Hw0
hYkx1Cizdl6AGD/GHAEjR5f9FQxVhW2IefNpuS9y/Mv/HSasrqa5FeFtMPxPwTF5
2Brqw+Uc6hRXb0HoXd0QJP600SKbLfVGsC6M09tlD3Z/UczZsNGZ1nF1YKDL1yIm
wMuhSkMc9OZydXiq4uzS13Uxg2JNuFuHl7TylK4WVqaEtufnOw/0y+mA5uceiF24
CZ8FuVQ4JLDRueNyLRWiFNBiIyMuv7JMagWwbuPHf52Eey/kUSS+lTpYoJYBRGzH
rJgqyAlXyljqDGhaslbnOmj9/uhSbn8A3CNowuN5RbiYmuAqjN0G3kDwmvNimscn
Pg5iVxcggYm3GQ9lekfa5roM0I8AmFC8Q3yVK2ezNt/ab1fmE2Ri5qOItR5qIQim
CbHRuKwhJbDw0FqguDh6z914v2nIXiwygy5MPguZ6KCjoHW2uxop9l7mEvHT6Jzd
SBK9bwR0QRSFuymiQTvRW6lY9qnBJBalYdE7s/dUtZz/H8dY8smiVf6FjamQ9WTR
Vd4cxjijwm4YZTTg4pQxF9g2cKCDRhozJLqAmV0eZtWOGUVmtmyaFg3SeOhMmvA3
hd7MKY3zE0YuzTfv71f+Vx90xrqJfMWDDclhZpYUA2UJUd3x0hAbjqxsHb00g0dT
sikmiEEIdf/7L8bMSz/8FURJE3i4C0WyOi/WjLM0sHyJPVZiR9qRsimvxMKqv02a
sY93YNHyW9aUNK00sYJ5jtbr525p/zw1cxz4EFDYYUJ4F1W3HTxPXkcWlKPSxI7L
FU0466dheabPMLBBCg5UMgZgiy7B6+PCMBc4AYzvg6qEBcEaAAJ7zCGdauprPQNb
Bxo3MTTAM5So7txRWvU/B168jsHUscCam79oPImF2hSg2GAPt3BCEhFis/cOE4ld
vxiAhxipWSFk/Y2tk65eH8P1mtvzaDnmUBkaUhCOriLy5Ub9iqYDt0Qho2NWidCj
BBWjQdqka3nr/y63lJIuOrLxhGTd1Kt8fBr6vX6AszS/dGr842xPA9swo3z7UbQy
T0qq63H9n8dHKfm8ZtyQ5XJsJSiKcC1MxiR+WqzI9RYrSG5JeQ2uiuojMvB2n84U
sYfbiNQvfLOHsAUPJzpQzVgE/7vEK/oGrd8mH7QZfnFNv2gi3kIA8cpcMVx8f9k9
F40hC/Ta9qrxaQrQxZxIM4ja3GdNqMGxMsIMYrwoXwVNqdNJBtKJ2EFjs3bDmaCl
TGHC3bzjpLX7s+lumtpLsDPfAj9A6TIK93CBDtagwZCW3aqnHVhGif2jl0oVkzDX
oFLrJjUA/Dz9x7aU84Q8iNLWBowkbucWtUHt450lP68iCwJwHmW71byScpismjhB
DIpcOj88OpFrGof5ztCAo9Q0HpvbqyiRpsiiUTzje+ovOUwJhy2trDt2SYZNn3TF
NN5VmopeBS434PhEPrJNusuyba6n9mVjAEGi3muIxptzHVUB6q9yQsvuyLPFnYJS
UNRjOGohwVIgEN7L5Z7hrQxMcpKKT1x9/v04s9v9c5jM8fr5MnmU3DhL2hbyw6XL
pdzZa06amO5+BoQ1sXvBXxMhU8JGAgrQa/2KDHc5wZk8jH35ejNjyRCd+OPdrJDl
DKEO9I5BpucydhfHsqRfDSPFRdm6uWw/k/5Al7GKFe48kwvxzruBqKoJfz3AHeyM
ArUOQFoNXunWoHNlcgN7TyM1Y1DhlonyZX+PQLSAg/o7EVKdpbrAQsP3ZsWMJib/
EHPiJurO16DEiNxFoFHmmHZ2mY7vibMe/g7+D57EfsqWJuMtIiMRuwfPKzZabiXy
pg9CKGiH8gfJKO6Q43YFrlUDbxXb2pNWO09Jch3HCO8+bvuBZwSJ3SHZ6NwMkhBU
lmml8wbxSDGwLnCT4/X4zCWnM+jWhkuXZZ/pXJlHsfReHhbPcuM0GKcELu4aGt8C
WsChixcm+jYg786WoL95qG51I7zE3YXj0I0rgn8C14zkwV/4a0P73B0aXt4ip9ou
hM5bJfqAXaV+9DrYUtrProqpHvcoPLclRWlAWb97DxSVLKpatOGni68V9R0bwidG
0bK73MIzJSdj3ckMjtKjCu4t4MTsLsYF5O2dOsM1jGLkVN5a0XrlI/W2qO7jI8fn
iUR5vN4nRtrh87TlnSDpZLcqeO4KptQeWWUzyi3vLS/RrWngcRc+HEP1gZYgH1Cb
FrRCS8iPDAZkm//4qPAmI6MAj8dTQFtGTvPkFDZmLqxEA6374Ck6qQUd4v5P+Y45
hSlCSEdCvS324sSiXNExyPSGpJ8le3/rVSjHhedUMErif51nx3vrO5chI8pahGX6
YdOkgaQiX45ZICkuTAvzDgw5OoV9dda0PzQEBaq2wuthV+dujsuLww895R2Z8TPP
T75lAo+QClg1AVfvUoIlZ1tEFIBEfmQAiS4gfhpMpDvWm/qhzBIT1aNgB6G5SD6f
2E23D6wpgtyF0B5mXgOuCTcoOdnVGOHtVNpRR/p2+rjVzfI02oGExe/AKSwqEA3j
P9rc3GEt8vz9HpES9JqDK3f87KGXNwMZx10KJrUhUZTMR6t4XTvLErue1ZjrFabH
QPdfI6Ab/mGG8TKVkTxvvVCuFWPoGrYAX+KcHcDhN9WHNIOPComr5G/fa5a43VnP
sORSwRd2v4+aoWjSRiVg7TmLdq3/qBA2EwaC3Z3spP5ZjXnMAcdUpV04C2ZKNUEt
Vm/lmuTNjMNmgI3LqkI7ywaFHNFqrOXZ16Q0k2sVbi6AMv67wubmbvpV+lKbVhkF
lQ/leCjY97DxPzMB488x/rpJPEst4ETS//M7kyuNVtI42ylZy+6nnzzwPyQdJpkr
PYHe6AGI7weJgkTGeKQ6my6B/Bc7N4138yKHmGFNw2dKfd1QmRmU2dw2nzxqINhN
uVMUr58G6JlowtZRknG27X5C2peCmScGo3ECDcs7BdrGDc5xd5SVQLZH3ILAIN8y
+R4KSjJlZjEUGHjL9ymbdMqB2TKVEzNr4Xq9xAzlCMmY7YqmeQivfIveKyXvB6xS
mNNlYlUB8NovmIV7RY1OW14xmOVT2qJLT17eh98M1NaqiBD9RQknPhimIaWV7giE
`protect END_PROTECTED
