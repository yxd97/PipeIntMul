`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zEkRgZ4g5lWBnwMcIchGBOp853/ctiZOua5YGYx89zk3PR8XQKGxC1wiagBGxyyO
WhZMGb4P4h47urfLB5dVaH1tJ/LuaRucbd68Vz92dFTtdQ0JeIDDR65/LDZ/QJHK
gRO/YtGiN5qxPV4OFcBHUg2bfBqFVWWlx5i2Ia4iU4VSYL+61A8uZYOsP5TwLsMv
yo5VafsxyI4WFVLwXBmdK08+Zj1LFUGq2x8r6H8vL7fJltiebcPJIAOjru+GLZUL
iavsTXNApkGwi+mujZdnozXi0llXiCUSKRUsNlVoB3veVZXF67h6Zh0tF3pl+dfQ
qb/MyhGqDpBN+nTzVxfyc+5bWH/CLfACv2wNpk1m1L5ru9sCJZ6/zsVxtd92xDGM
S/3ilMdn4pvGvqI8yml4HzUzWDs68grV6q50I07OoRjLVm2JCRN9vQ+cu2/CN0BG
aRa01qNwb9//bQEYztewSJtDFwv+aDgQoV3m3WNacFgCefwhlVPMGgO9ra9oRH2i
g6btaw/qsb2pgHYh7wyRbWhVw3uo9BTMx3CyL26h30Gw7RAjJRRM5uqc9n+5ldb4
mNEKlC1ZmzWMRV6buCreIYLA5LxaYtWArtPoITqymzFTHmCtHrsr9ExklTrhPR5a
Cm7yrp2a8tEkkoHTiG967uCD3EwAhDQNH3d5MGZx22kxMwR3WtpBOwJqg347hzPL
4EBjh86rU9uZcDv2TiOfuCIricBzSSEVG726rh3Qt2+iG9Gi/SbYx9X9kjdDA3j5
nKLdKf4QenLO1tjGkg4jbOXk39upIKn2T9I+Eqtp5cZOhhi1U0kQuignHcbbFIVL
bwjemJ128p9n2dXsav4OfFV5fIHZ7OebmD5vrMTQzK7OmgxcHI78yzyssuAhYJE3
Kj2WUwgZL3Hmi0reH40h+Tv76hrZFkkmtDRxqLz3bWatpv4CP3rfdEpayjQy/gMB
QRijlvW32c1S4P4IRFChrdAaEDsUGm1yWYO3SNl9HciZqX9p+A/uNddvrNf25Jnf
`protect END_PROTECTED
