`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
shQh1acs8fm0WgcwAYcYGNTpV5f5Fr4HwGUp2ibi7m2KVv4rgmM+fw6V+Lwe/qeH
c6P5871XXGQObgiXagFBRNfYfSLg2HGwWuoaHaYoq5RG7Kn7V4LTbhG2r8B6JC+R
IA7NDowZs94yWaX6rQptqGZvRcQA9gYigBTAoT/Y67NIXxgTNcF0M5yS855WTrhi
IWkd/urJAUV6RruOq13km2LlUyLcVNnMJrFU6+RcM7BlBb/8QdtwlQXXVFHTaWF9
`protect END_PROTECTED
