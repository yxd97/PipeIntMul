`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+d+7AVPjMwGQPmgV7WviCM5vdMFn4PZq3uh9InLJsrtj/qiveK1NYKhBp3JXOxo
lr0IsB478heKbqz+6jFp9o8N7gleDf+QBrRHMFh953egBkKTxdF8OpGKRCRD0XvY
hoqHCxal4XjY4N3z/9LhahE4oI2mMvQ4fJ05MuDxNUNuqStzZj2e7aXaLniKKKXa
MdRn3DVurDgqWtYwa6l90+aQHAfI1P1lILLYecydjqoU0zmYVClpv4euWPYCHt6q
Ur2hj57SC8tKfEoaVDBe04XGW/lQuQQt+ywtAbh4T4H01fF1g6h4yyobxUW7abQV
j5sqtBcqajR9Bk0NW6iryyQZ7vUXQg4mUKsem21Wd8apUz5IVQOMjBgARBorToxS
4kXcreybTmkW19dCUqvppRMsIyM+UMQk7uxo83FfskLa23lghH+3ydD54XHZqC64
De8e19IkxyD+If4Zp4ZPyRhWwqMRJDVhrbEcE3Peo6P1QcsLeJhzFsz6OyQmDyMM
EPmLzWaS+XOiFWYnw0NQfzkQFqEJR8RpmJ8pQYmrefRlhSU0IToLExy7VsNyXNsR
Q0RLiOH/nhXOhwSEF1Om3VS6/GX9j1MlbQb2VVO4OK0I6lrBr4zxbovEbWFsohzc
QdLmGTo73MvTwNg7Eumw0Pd1drSDIBcIZ98xijkyQwQEK0mfeIow3T/zEidqElGu
EErhkRULQ6X7nnQBBRS5TIX7nZQVIBp+goAAWu5Vt+LldIgzOewmMM4a7fuenlAd
01CThyccS992l3ZyASDFCLomPGh6webfNO7daMd9PEo6T1okABVOtA/VZs35O8Eu
PdWphTAhPlA1AR76BC/r38SrxutqZmZXc/gRL7pDInYu57lWHiHvIUpYTFKO3Cyd
ljCmuL+PhOputNjaEaKUFPWL/9DY8JK6A0wTIq5wJYtMuGf5jXA6Sc2FpE93kzgM
EmxvTPTSQt6sihSwpeur8FruNvsWvs7ZYoyCRLQ3HG+pIBbN8fn1+cy8ZBUOWFUt
cperQQEQlbJ+z7SVyzV+e+zC/llEaZyC8oYSZ/Z4BRzquDYpHLqGpOKIbpAVqI2m
3Mz0Q0syQ5cBXt5aDtINM8rhvIrqjZFA0GHAW4R3u9Gi3YBmMReqlVU4ZTCXhiCi
Zw7uHZmTW5YQUVgBitiu1L3hrMeE/9+Yjvpuyl54BRiaMoiIgECSXotWUwFbSOW3
GAP02I9qvlhBls5fRWNm04oaqwshgMU5VLCZq4RiA0ugftwaMrgVHAn3FXqbWYFs
rSoSgBwERmuiC2Ts+bSgZYTLedF2T1mhnd0GLhseXwdpZwoZipE1OXA/J2Y6bfdO
uapL37zt6qs52t7xvppIsmN/2W78NyZ8GCdwoEDSERJif3PjhTOBTdofWLzKem4u
sNZ/j8YlysBrIpoZgDiFtH/r7Xoj/bPgR2rPpKCHrjcDc8w0Heqvw2dvaNXwXKfC
zR5M/jvPbI/DL5OGnr94HKFRwuU8dy1yVMvUex7w1FYJtbwCDaHRjnNTNSKBB711
o6RW9fE/+rk2fwA415IwP9hZzxLp0bbeNR/u+3ZfXvJu0lNkdDGl0rYZV5xPV+AL
l+baGbIl1ms+B4PG3xZkCaGQG1zD1R21sudElcfjA+G9UWF4ihcP1H0evc4vQQsL
V38RKSInbfES+oang0jAiPVTOEj6RB5Hffn3iwFexMXKSzRBYj4fWWwzFfzmeFlv
9tZ1sBekrS5HRe9xunoM++ei3lrH6xnHjZaM+GrEQLDLkH5tMQqPZkRkg9R7xZsZ
iGz9X7hJPOyDFzThuNj7Qgia3RyFKZFOCn9R10p8IErhmJWR7tTARMy8rKegAyPm
FvMhJZdIrw3C3KXnst3D0MyF3udv4AJP09sTk4iaeUeDhB2Ac5tUvtuqP0hjcf2d
WcscpGkni3FA+KOaQaHm7uTdWlvUprsPFuAjeCTHz7xq2qSEkIqBQagFEttxj8H4
bFGd54ay/Ii8YwzBvQudtEK9XMNCeHsu0ion0hW3vV1PjfJ8k9Xu0H9mAdSQs9qU
I2VNeDVUKCIQTMP4qBbkU9yXRq0nfuIoU2YgPZg+ekioQ01edHv6Ocy4XWneRUQ7
K+BZeDAHkLC2Z8Em7DEapgiTyD/PwDzB/eUZzDkeZgaR90y922QEdN8DvOQBvBjB
26GSnhVqWdhr579dyqK+zZXY48TlfRv2taLcFoBmYWoExcEj/8AC5Tqz6i80xAoO
iRjhe32p4ZnCsanPV03pFwFRyv+cb7GNqt8V2/IK14zMY4Qwfb9sQlq/bxUABBcT
YD8wDAsp97ezhdtB+HX52EYTTy4LC7XseyoxLLs5DOhbZnQco/+tz8WTBtaCaw4L
V3SOQYLGqVj2X9R5HB1N7+TGwn98s/y/l4PjJVwx1mqA+nvLiqQClNaNYvY8r5bV
Lm1ji6Z9Jl/ASaynbFlKQcJ3r33fC86pasmgjTbGH6nm6PWA5ScB6dimQtzSqT4g
LzfZim7giVTyY4YswhJHjxGTWPINkMgBxrgl55S8t5qD5lXH3jPADHEuBFz642gA
GZjGgtuX+tQ4cVL2gPe4ONk1ueZXpQ5gCFIFhC55I1FFq5WIGjuz3mu4m3nFOLOo
qfix6hK+aw/gUuv3b128HF7ghP7BUnSRJ7W937/nWLxVq5PGcoZ/JIWSXyT4mAut
kETom7biuuqyTKAppjrW+cYKTLAu68IN+pGlemqMNxggdPGx1hDeYHcYB5GRmoFQ
w+8D8Xo2pIoa8qeiZXTRGEa5FvJ96SCcX9oDM5kj8fQPE5wxaimCB20e51ltOZcm
r8P0nUF8GzfYMjTiXTVvSslZAt697ufF7wtu/sbCt4JSdb0Qt3PDlWDh4/HQ4m9W
FN86FmKRKBYO4tpz2yi9dT29EX01k/PUOVPmK2TXAisZ5SMEL7FB82T7o3HV4/z6
F7HynjlvSvM12ep7HMzBN0j10NyeuFNYB0C1llofiwiV6GuJxHWAgW1Yc26qhRJo
ibNAuSuhR6WJYSUnW+PueygAoKAdlz/XKDwt4ZTVEmuRK+yBVdF5EwW2Kb5Os+ZY
DDe80A91ADb6c3gcA9asOrWUnssMnA1wACnpX3RqAOs+7Yn1f/ZTAPxXSMlLZ4ro
WJyaEWBsZ+9xpP6UgMiTFU7g6uHhmyhF5iGqCnNMsBQVgkafF9msQ3XMULtTVj0W
fZ7+GXgV3bNm6KqRyMYuMG9tp69nzYCXvk8s09giKL9a66ppqfmiA4/zICTBiZY4
zPtqf6FcrPMGu2IdnmyvZ78XYZiv3PMCctdPxqoecBXpdoOApVuLid9nDpU+5vxH
cwQBBFaqy/by4M1EvMLqMkLt3K4c9ZAeipl3m4KobAEHIdZUlDOgvL/X4GsMB//4
tXd1KfnP63SjdNydk3b5uhh2lQraoS3oD59ZMH58/m0UEbXCTn3Hv/IqtE6nDqhx
6YVvjjBtBkOQGI3HH7kWryviFSfAKYfuNmNm9+GqRl8=
`protect END_PROTECTED
