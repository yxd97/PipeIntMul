`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
og6f7xS1CdK9hzeWLFbRnASCxAPegzUvtWcav1F+xKqxPWYraLqm1eSzaHoOx1a3
KrvmbFpBhvB285sPZsVthTQBuJXJXiFMmnvhaJo8JsL9DuUWWrKsATsAz4YC2Gyk
CcmOBK0JB5j02UiBxnAR5PGloOO/UGvdAzz2h7Tscfuv7HX6m5SVfWtBhlbfbkhE
aYtj1hLdx05ssxs8fPKiyas9FX6pnpc12W+iyQeKZ9mSoYfUFhIWwQ1myI0E8uYT
vtpb+xIJ6COvw4lP7VvT36GaQUP8rqE2OJf6Se3ERzmbMxOluQ10sBrZRu9UdI9b
/cgh5WziSu+fxS2n20WCDXPd9/ZxdsJXE7hocGl/BfTlwA4jiUNB7Tqu2J9yXsPp
W8ysjugk3/ycl2xMKBD4GKuh57uRCoy/6wLmpCveuvHrob/+5wkfOPgYoo8FCAKO
`protect END_PROTECTED
