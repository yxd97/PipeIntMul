`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGr7WPX9rrCs3sQbbuGhof0fBDRcTB8axIN7hyXy1xNeWXpJOGjZMKXO0CYRORqx
EDWHo++iIaWUIIK6Mt94U4F2iI7DE4Q9avKfSqJTH1AxgPdSCjXinLsZlbJ9pFkz
xtD9fRbxDOJePRUA0QuJOW3TeUW3oWUSZCZAUK5tN/z6x7ex3BouzFbMb1NKPkEw
tYWbFqg4E5+bZRwCG5bzORi756QAeTSwVqlU3H4OqDRCY6V8shxZAOSh6hS1+UEA
hdhNANo2H7IO5NdXz5wDOrr/OWSnB9T42PUfFNMi1EV3ie7IUU3fV29+dEMmGnIy
0SWsFQr7XRyw6cZKF8AYnw==
`protect END_PROTECTED
