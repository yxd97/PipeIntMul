`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+cApK4V9i3sz6mrOXvkNrHhRitgvWJ+b/r2rziIl02EDa/MleDTSgU5AJNJmnYp
ZlQ2xh4SJmuZKwQpsiT1/Y1T6ttcMNGvXIDJ78yRovX6YxTL+hafJY5CPZ0SwFPL
Y0yh5pkqSdbFshd+48nPCJ6JGbeYcdqqhMahE2BTpG6vc7ntqQh3YR89PbPUiwE6
xT7Baoq3STlKUf+7Cgh9a09ddixqbkD4GTYkL5LB9HSrnX9cbifDdEB3+JV/Alxt
cwJAxgGu1IZeWryzujt524v8rbftAyxcgXlNc/9mHpv8l5u9NZLWAaNX27u6RJ2n
x8itJLNX0raRok9MuBqzqAUimW/gin53oHytkG/y6zFtAPV/jrglJogrn/7mjeRf
d0m/wnzzbfaDCWYUeVgHZupj18ICYoGtygU6MX0IBPRk1+X5HF7FEOUahAGzNqzM
KDmeDRoK/8zbHK7b/5DYkJ+MWyDHjOfZCS1kIY99Gl7MVivU0PEXMPaMzWQnCMa9
Ydba5dB1OG1FNS7Gyu38+cP7emOp2cEoPyFjPLKQ9/bd6vHIZkL57Oy8J9Ph+hl0
8akiZENPkoodXvVILotqGMC21nlWj5a4VCVqMRj4E0U2bw0AZ+4jv9GnsR9ktQL/
McELFIj92c5hrTKkSQPXNkrm1ijs4UnSC5nh8dmWmAr5BrFUqi6m6ATKpiqSZ8Kv
XGkZKe9UWaEbAerdCNa/1iIyHROHrbJP49whefWd+3LgsktsRno77SgZokr7RqUS
Mnwwk6ov7pYFrIJM1GBp0ze2NfgRlnZyGVpitt5bFwG4FxROv0fk1sQeIKUvutGJ
VNtM5rm/8LANyVdyFyuBikYKCCOrdy5VMCTFd4osv5Hn1xofvi5hF5LQn/IlFhMp
t+d77lFalWxvalkNEVN38lRNkyqN1Z9MuZZEkZ5GSymCW4rrcR+vf2fdyOBjn3aT
FGU5hXDN5sBln7ji+L51fuOu38kz65l61KcT82TjkL0/lioUArlYXcwxWpAhKcd/
TzO6JpBekZ7KDTzbma+bmg==
`protect END_PROTECTED
