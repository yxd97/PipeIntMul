`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OkOqK8sp2/b3xjwNNTPZOufH7dtvDziKS6YaXawpJHxRGo5DWIjn4ghdissFGjii
h7Nme1SZ0KKq8drYKuBP+klvdkhwcxrNFryU0NeeGaCauwsgkh6Vo/GpSfO7n1cd
gb8PSyMAE+ig6szR9k0/Zb8a70+xhSUYtW1AZneYhEwXQoZ/94XbwaT+82ceomjv
tUVsP+E9QX7w9a0p3LExnzzER0XJSv7qCZNyq+rUu3yYmfPi24f3MtiUe9UT8FzL
ngkw6Nwm6oFUaX58Xy5RLQyxcyyVvNr1FokVC1gGtrbK1sTvbkSRP7lByKLfnpe7
advjKpJwPDsFSciUBsyjAx51vlJZkh6Nv4ft3rWGIfPcQk1O0bBCxgsgZLQoN7n5
sIV4K59Ozg2CNx+hPmv6mNjjBM6hSWaB1cYRB0UUEq3gKy+fveXyaJtXHoLiH07K
qpS4irK/OkF5KaGPz/3www==
`protect END_PROTECTED
