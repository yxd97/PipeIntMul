`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3mcgvEJNUlJBPtof8tuDdGDmztdUPMJ39G9c5gReWa1viy/c1uu9PuHRTVbLZLe9
PdxUKH3V1dCgVfIhmxXdn4hSX5GHNAOv2kqZ4NBA2OlDyCHsagXTVwWYZ1xiBl6H
TAQGVRDlE+ekoUuiei8jmfciXf/K1Ad4kk+Hmzw5BebJDiBgB9IDSUbETh4+riUZ
T2t8vbHYAzy43CEy9QbXRNpVPV7Tq37RIHSqLjQaiUeA+VXLLtRE5UqWvFDq1uzb
Dj7NNKkSsSFsfm3pNybov4TZNJkKrq6A7PeVXJ9Qm7JrYvEHsQtKUy2lzoRkK3LJ
KbNYQkCsgtSB/CL61AtLtjvoU4A4R/VT7aGnK9ov9gPWMVDcGRIvSS/KFocRmV86
hHdcNy0noqqtaiAGeuTBoBEPLWxJFrWjyNu3ZIf+CS2proQdTO9P+a/lN3+pCK4P
qbVGD+C+UaPHY0X/mKTsBBUxXHVK4w2WnmW3P6ULt8gMEqvqi6CVWPvaXC1uiX0r
sa0TetXgFs8MwaX5lkrRp3n266a8uP4+AHfWawjAWrW01kHZKJ+gdFlzTh3OlDzj
HM1Zen1JzU/uFCkMLIblty88v61btPTwlAv3CtRYlMFt8Leb+iK7eDpyms1iGBXE
efsUJWBqGkX/UKjh20WaHz22az8EjDLLm7H7whbSc2KA8BxA37hTFZSojGBnmPtH
lcePKTGiGAt3VHWDx0hXigSwheC+j5k7XsYr4Il6dfM=
`protect END_PROTECTED
