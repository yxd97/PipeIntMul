`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XKumRXcvzZW/wdQ0O69jQiZS6ONnVzTred8tyHw/Ltj2bQNROT9FChRTGt0csVQ6
VTOLfXDYx8byuDaC5GYR05SuM74ksoAh6KssOlfzoS0IUIedf52IQY/U89a1r87J
WfMqXhcENjPMzCK3ue5fvJEL9DKoRY3oNg5IPd3aLVa4oJBm8YzDjXn8JSdxwd58
iaxDgb6oqvFxNRV1KfV/jupca1Roq3IZ1jKuYpORM+DjMyEkBGfwAjyGvPx64J6J
1KkWFnLFMQsweUT0zJ70Whi9eEhG2cZlj65CiOeLI8EMATM9czPCs7bjd9DtJhTi
DvqnOHdnROQ09vpQuis+bp3Ish1DZukdxqsQmZaDfm85+NgaMdj6fpRGudJZiPHX
8tBmVscwl9nOd2A3dZr3IXXaV3xaDfe/ibDzrQRGedFqfI8NcLUyQ7ZUF9rUk1GX
dIeEDYEPaYKyF+BZ3G6LKgLj0VhUJAPDx2svyTBB7Xcee3Y18CGsPNxgY8+B5eL7
BLeKdzhXdG7zxNCJ+ubn2YJYHJgcTD+Uuz0JsRbq64QoyhDjxD8Swq388jBgoqnv
GQ7H5BP/oe88yVuTS8XKYDcZmgr4B5VvoZKaqSTJXvo0WiYDtA0J1XEXD9j/pUwD
1/J5gvP33dhoeIpdGn8k6NxJtODsAwUf3Xhs/OBrT1yURiQ45mmprFT+oVgXXLy5
tJZzqnYrHz4uhS7n3GxCOQmOkmDj+GzbIENMatrwhHXGwUKEXlZWykydSIewjWDR
n2vIJBqZMRHfwltto5rf1moQKcEaLgwAE6pRLYhsbG5KdOuo9//HTcwUJmXmCnOM
jI3QTxnEiKSvFNZydNH3itndPbNTzAx4YKFve3+mkaq8jkDHNuX0Qbk49zDX833R
jNuaRUsU/BLSq7fR5b9cAkdUhd0/NJIdAD4Bkiwy/TzFMMLskqkWyxZxllA1l9zu
q7ulSu+7eGyeYBqKRi2JhQ==
`protect END_PROTECTED
