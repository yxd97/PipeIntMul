`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+WuyDDmnILGY+S20RkpepQbhhH3c73gW42cksqu215gxVjND9+Qw6bmtAmHRP65q
dW8Hb9KuNGpkB0LGVecsL/1O4IHMXrxoR71fQ2snxdhRp6gS3nDM2PH8tJ1D2PRJ
QUpMq8rnDa85QuuqHYiC38URsYbbBG6YwkErmfvhSQT+XzTx9qRzUCsah/jx9IOL
dR8H3BNW1XJldQmQyWhnXMOoDgWZ1SEMmNcMk0C5Rc5mAhFVaWbAkS9npfbpAV8S
yMmusc791sXeIPVzL5OcBVztGIUoxEiw3BG+zCulh+YqK52pL1kbJm6T/fhOXtrG
sKvALrf0ShnJMvZ0HCilKo45XLDly3hygKbrmpdGZeeo7cBhnWUyUSuIoNOHQcwk
QtClWPAIAan3HXZwyfqOx+lmSo16xI3q2hNTQTIIpvWMZHvAiyxHnp1IFTlixg3A
eGxJrO5EdsPliZ5/4M/DQjunE83q5ilMdr5MNx34pjqo17HIA5GQfyWOvyCEz62u
l22Z2CFuMXNWtY6jofGXCSkbl1KC8BbBYF+kt6LsM9J22aqDNbSFxnBWxztBIQpJ
QyfBi78P9rwxAE9a3uoFP5IdAOBDHOHE/FXzE8hcZ84rs4KIUbcXuMAU+VOJMho4
sDMhb5RPx0M2O5c/NaEqKg==
`protect END_PROTECTED
