`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MC5b/XeLgF8tVwM5NihM/6cnovmeg3jfBSCCKAiZ4BVBMUAQ6jseriikwGTlFEaQ
03U2o3RFkLgF2KEt9t3bKXi1RrBRA0WUosWQViAeiIqSnGaqsnIJQkpU053du1ud
yNLRKIlfmR7xfJPykGRmis7mfwi3expO5ZeEfRPGaC9PlsSUlFxEXGD0qdMocHHI
ujiiBBeEnt+wogNdE6LNByK7BksI88BcNgraQEoSiIUTTDuNXpAlyJssFsN/iKUK
Y9Sf4nwwIqhxZ4yE10Mn91ghD+FSKT3vUMJ4bTGJFeT/0QciJzpoxm3sAM6a0Gpp
I2TAnF5fag6/ghl4I/Mwhm1aAwsaFTNm3q35WVHzvBXiXMz/yPVuExPYl5HNqRNn
mvlTeP3GBcqMUINZbUz1AA==
`protect END_PROTECTED
