`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tRS+iTWos/K3/F018emO1O7V6+KdrB67ksJ3gln4TzlQM9k5ouMJSfBWv0uv4AQQ
9RKWt6eJiRuA0w+BbCUoHY+LtF2JcIwT2cqA9UqhfufVJSss9/nghSD7otHr7yvc
IbN43ugPIPDzxT0hF647opXg214vw6+plBKlIDAmMRhaG2wytMw2MQ9astGZ3thX
7sG3GycFr3qwMTe0GiWlt+B7neh+hIRUpfytdetgYvnGFsf1oX4BCyXPUS/vT9jc
30+WHcseBJzp7M4flgFkzvNAhni+Vo7mQJcBICoNuGBVqtSX65EUJ1tMeqt7WKnH
2enTc++RM8t+0VxUv1rtALwRuzu6dFsNXKKUTQaiMoqTliGlU/WyFFPjOsournkd
RIOeXGy88i2ZSkz4jDsFA7k3cU0+tivs4QubT8fWJ2kPvt8f4m3x99CITTAUxb+9
6Qiw2X326GYbeI3CwU5v8wW2doQNPzFbFyxyP09u2pLjZx8ClhlOzS/7MQO07twp
z2iinRPly973UGKBTaOmEscftRsmDmOvP7GEQFUf/lYye2BjuUVxAmgF6OMVfjoH
8/NykoW2FPmxvsiz0fIHhXwflcv4Bb1fHvJb8BxoO7dlf1a1kNGXM3h3EmAkmegX
QZXgQOi3nV0RgDCFnKsNdxhnNR9JmqBRTj58hqbYbPy1unsDraRsgnnw16mnpnqx
LP5l139DPUi6AebFJzdY4Q==
`protect END_PROTECTED
