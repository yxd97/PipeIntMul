`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mva+bBzHSnenlqMpHuQ2NLUtOL9gcLAfbuGl2LzERZaFlqPFQ5sBqjQXOh36hkV6
7uKj8dIUOyByEqo8lRVyL+KxbIsUPNc695OMBT1V1tvjTC1N5PkftO2IgXLrJ2BN
arzOcfM3fgUWJM0jjrsxYK1nNI5tj8gWmScXF5QTumx45jkCtmF3yP9UIdut+qBF
a+oPlDSrqwteKWcTkVglwgIpN/LfQkCA1zif2I6japfwRtvJRe8F4JPJuXWa4VIF
rduZxq1WD9z91QXQXE8bRNLrSxMOtYKVnSlMRQPCZxYu/A19Siocs7r+2JYRdlif
zJpo8397B17q8bS5y4PapLycmEJrS8n26/8q0P3cNgCqoHi624fCfyA9LcDAiKHy
XqmAmb9nVQeH/566HFHCYne44GUdl9QKFaaiEaYDaN4dyhMhi1EMK1wzguGocD6y
PBdfqYPtGlv8InVV7Oeyq+4tijfHnifU1pb32/vIbmsLZL91mwZR2AU8OjKagKW0
ynh+7u4t8eg/GMpJU07p0VSbnnwwx++YHHzQMLnTTa++s0UmNuCiVlMPkFAukJYl
EQJ2dATXMcSW9YwjxejDU3oAJURFxYKDCN/G8hfl36SJWvvRtXFidz2HpQNhc7fn
`protect END_PROTECTED
