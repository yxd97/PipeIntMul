`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zK9spREtB9UzOjBDQ86DU6bLvsaTMyABSDcELCcDxGEhgDn9dwv9cz7fdGnwAB1
FmFlEFxKjuPC+YnQZ/A6ewoVipVUfrSI3dwPC7FxlrOtlKPtO+dWyFReA3yNYmpt
pb5JcweMg0i+MciWZ8TWiHeNlZ8frp3g7OaMhjD2qcyzWOcKh4A38uO+DImZ8Yi0
f79x5D/H1fIzTpfPD87JY01x7nmn9LPxkiroBcfVyXXI++zlx3e9qeYe5RZncw/g
Mt/idztFKRkwS/XonuZUI3ouboQxeld+qBAvYuw5hweqLgy4s9mRlDkv8m8KgoD0
oJ9kiwIp6na3nWsyir4csYqFsVqidPk6mygOC7h3EEhCtMyfzkMSShz0bb46V3kH
yLlSTVzN6FYWtRnOgraOrlqASj5mMzgZvGZlhOcTCxyp/pPNqwvv+w04XhXHhtEv
zbxpLe8BE/CJUfjgB+MktwlN++sCOkyGKThB2to1DLM/PHJ7LXPH43W7/K2LS/Jp
`protect END_PROTECTED
