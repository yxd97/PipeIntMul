`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zs+n4kkuYZY93gli/ZG7zZrLAslBTzze9IyTGypix3rsV16jHgfY9aZjDu/+ag4m
QBinoERbbGX3ZCoeE87aAR82UWM+AZmv1Y+sicOFxm1HWU0XDT1ueYkQJuDRA96y
GzsWU7Zqz2kTWwItMXz9PUe+bb1Pe0AW/8O1wB6cvVJEduDpGgwXR/zevt87AvC6
BJj5sDW0b9LUHHn06xrAvpfmNVSPrFNSkjwTRB0WhqVnvGVFxGFsPv+sQ4U8acIc
757+3Jih6Zg7c+3Bu4FxDZNsQsHqxy01HSZkn14S77s=
`protect END_PROTECTED
