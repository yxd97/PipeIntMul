`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/ixFfTXCNTApyMJ8sc4quFTyfXGhHnT6DuTI+9KgUvwY16AoGFaiPWeLgTXfGwB
HaXvDYY/DysXRDFUOHS5BP/AViQzHEgBLhb+jSsyxAfU29SBOdsrr8oe1jfkTzgJ
TZUgm8JHudgpThC3Tqs3exvkmKGVIZBuFb1V+wwTUSjVzSA1oIRvLdyUDwK0TMin
3Hk1ScQTApHbleZewOTO+QwwDMGk8BCP3E02LJrbBmnkp1mcck7fQCOC97WvOR3D
Dgi17MVRgX+NFi47jiTxG7LF1G+W1eROSSj7ZMWRXdpsJlM7PF3TOG06YuqezDnn
72BLykaUG4GlPuFhJo8wpGj+F51v/Q2PJoNkLco+jKdGNaQst3HFSKw4p9WzAjLE
oRNDe0NVqR/wREkeN6FjVvs9sEeQxlFyL5AMlcAiQnZulL8BFCe0qNUoxl6oTRdS
3Z3hEyGxve791HiOKOjg8Duh9K0EaOXvyN5PkpCWN35JGGnsukfLLHzQ3fOdTKQm
eXSoXaDDx4pmGPcmPI9tBjj/d7zRLxZm5Hl6o+y+aLxsjANdLZdsZgO40cGV4h7b
nztVrHcJ8qHh3/vR11rq7NIu2d4BV0LveLDCAJZb368ITAESAR5HOvihjVBxIV1/
WoT6iCHcPWjkIYyryp1JIZM5GUf7Q+Pk348qxd0YiNDSFyMGpkeTdBXkitaY01Yd
qhERuSWKJk98pYtkLTOyahfQnHktw0+XrT9asLXdtZbN6Yfj9J3tKFA8idqfWGbj
p4EqtP50F0KHYpBpTqEgqg==
`protect END_PROTECTED
