`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQ0IDaLW2R159x0LcyBSIhy6GVIDcLjeQuGbEHoRmXw32NQ+M0wGSWB3onJBxxdI
iqb9Ih+453qrPwrwL7NroOjn7zQyZ38yY+yOUahnt+TPJdG6Pf7ds0uf+JQTmtkq
6ijvKv7e/kiG7rKLuGo7fnwaTCzcyeqb7Vh9HxaFbI4xwRNFqp/V/ditfaeqRudK
OkF1UBvpl+crZvaXUJUPgbYhlts/WAtzlaU0MocbpGTSfx9X9aE827dFtHqr6szI
Syj1q0bgH8bOPOhogJwpFDiO+OSzbRpp84u5t0J9MG/B3BLiR68oKfEWTKROusQY
15FWi/cBFRQMINFKLKTm6LMiba58phHIQiaAXO+9P5Wn3DeY7WjmZxGPUoOi6WSD
rbUsf/xZgqfp9x0Pk5inw1Gg+OskFOH8ZkkgVfVfgBTjc1K4zCBM7g4sbwZWUcEX
Kue3Drudlk2/dHduiGwA5boaEGB7z5V1ab0V/yleJR+lNuX1O+vx0l1Xq5McoKGp
`protect END_PROTECTED
