`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqMW2F2AgUZ7xL+HA0sfiksNdGyXp8me2E2spInoV44w86ZqaKdFbKfBPU3QrCwc
AFSh70uC4FNSQyC3AXrMhpKmdNVKvui9GrzygsTWRQToYpMbeAFzzA5bL1W2saD1
m42hD5IMmqBWwfcxEUfIe64TNTBQNCL5n0Ji0G8i3R/TI7ZUxh36bXXqlx9dyxsW
u8Q3TsMuWbB7hmRYlNjzsAbYCgxPYGg+GiocilJBxU9bKhQEXYj8Jl25vFEHWqTp
kG1g3VYp2f5Jjd3EuG8+IIdtDZaSFQdVdmDjaMQ8KmNuRmO+Fk35UBjTA5G2n7yx
xZnF+bkJPOLAbiRMB6nJ8kbpxhhP1ial1ziZasZZQnbRV5AcNKXHCHzEmQ/wjlAX
exEKHMYcuKrpDIYhGirz5dq9gMOMWhKn2Axlzpfcy/GZTVijg+JPWPvfPEKq6VdF
wICmzOFNl2+tnyak9+uSRHsNckNGfMf713sdxx+kWBXgy+KNF53NuyAHXyW4xQbn
fDBMzO/W4wW6/CGLGXZAwIzDOQpWxowo7ip5bRENkW7XKRQG9fbYbckfizOctdMk
vB0AH8oVzZNsrG5c53SCK6VKjFI/dPLXen+DoE8OLsFZdvhoWCiFR/FvnAUzekZ0
UaOOX4aZJEpBKHiDoTFMi3ITDXlNlErE/d0yk0oHoE9r82F+sLeg4ZcpCUVcjGbK
Z9KhCGPET44n8af3m8j+/9d8ZwLQBCC2d+d3ep2e8Y3Gu9bkKj2hfHZvBFoCn82D
04zpEtfGisnDGqPCj1zu83NfYdTkPnN6Htq6go7TPf36Z1M+dKS17M/dT3uBtiaR
PCTZpOJ4wRQ+ni4TBOkERMuNw3u56DjQZw4vieO4K72YC6jHCLGKZDuvnH0nhIEn
yiby3WZnct/CHs3PeqAQCRyCmRoj8mmwlGBlIJDKoS7+8oP2QVUsx2X6n1X4sDwi
xjoR8QWewNQzNi79u4TXFugHmE7ytxoGEl5AOjTSzKcHdwduODmlvA+7jCsnIfL3
f4Ardm0Li7ZoKy4Lwrmd58B00RB0Nmqw5BR/H5NkIyba42r+xp0Drr3fuzOra2Gi
gKrRGKieqiOAbnFA0GykBeoehHQQLEfHYyAzyXnUpoWo5Avj9YDJQ7RUHunHO00Y
jur1KZPFYLUb5LeMm7RfG144bVoXd/zuZ3tiCAAMPg9r34imo9MvNEyW/7qI82hp
Q4yEN9BXVd3q9LRxz4c3Qg6hHxaClzXy667C0JyIlZXSp1VxKtZZGHCwAEyVBwLR
+swyU0idL/m3gJYAfYUjY8WfNBSNOZ+rvsatUWM6DSaalnIADmIAKkPgn6AY+YKY
cwADbpvCR/7FBPkG+Az3/lwutKPcBjfo8jci8/ut1jcirrmzGWHhtpDcaIeKWe36
+9rIPi8cHu0EYsuRJJEm6KHK/DFJCVYUE+oRc1MFmaoG0PVmYV6VITsijrBdSO8B
NISDTnM8J68jMxNr5XjaGffl/bCjy8UZSwdchcxSfq/edqJ7HBSvX6/zVC9vjw4N
bwDkrNYNun17a2+YhqStrIGSykj9clVOu1kVIYlkWaRc1lCZP/wmwicWQaqn0pTr
MTvaPlGt30PWjAo9GEF2WNHFNr/y2IiGXcvEFvuayArPm8md0FL/T44yZWrvNQ68
G4qobyL6wp8f0+ObJaFDPFvDBKbaE4Kia2Cjjfx0j/aX+jANl4ko3doaMde3M/rI
8PZm1lVWcxG/GNYJH8IGJIXkUc7I6HT4Dkofo7m/Tpqn+iohYeqLdIMt4jF36BvZ
6jsI5kDV3dIOsFOaxXzxQuZO7ckERAzhGFMqsc6Q4vAgMzdYtxKw/mYV1rOktTlP
YBukJxguERIPcw9l6q331/n/eeOKoX4OeVVQw8z05u4HrJXwAysrMJFic0JKCdxQ
aQEwEbAgGzX6I6eZ7ranXNBSOSQaZp3h8mIO7jBb2DBxCT5/pyaV6CZHlXBVMzgZ
H46FHgFMvmUmjuYJQ1CIi+nb0xE5YC2Hei55dUO2G8xmoK8UCyK7uE0XLv7N7SGV
1qmKeQ+Zy6NyMm0ycFuvajP+mx4eQcfIA3kcOru5sjlbieoO/p6kVsXD1ZVuqWJS
CFoJfrgfkUEEGymmJOfl8fgsbeao+6HqCxdJAo3qaJWD9NzMksh+ih82+ASoPbmx
rA4GnLAXYqNssOyrRgqhuzldOj5oGLrRK97bDicOPUABFBlvoVeqhRN30i1ItqAF
hP7NIj5ArKRlmBNKPiUOzO1axTyqaOLeC5clAQWFtvlKzIJTPOBa1eOI3H4fiO4N
pRTqao2Kl2bme1M1Daiy2A==
`protect END_PROTECTED
