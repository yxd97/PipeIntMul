`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vz/3FRQigktyHnXG3NXnl788jqYM0oo6krGg/DF5JYmVPKVM1LsTMhtU6VHxElRV
/jV+R0IkXUthzTWP5Ent/B4xkkjm1O4ItxReUbmm34/AeRlMvfsx+132nt/8yj8T
V61T21truYaKZrINEDbZpfp20Hrp8CAo0Uj6jCkhQMj8gp3PFZT0yVOjli7GsQbA
cqAFpwG3Lm+sl3QeP1/YzjA4JnHS1YZIQ2Az2vnEha3VCpZ2e6bdSu6xe2IUz5iz
Jrfxn4AzfKadcpUOv1wYjywWd1fmrvPFKH2uV6yGT7tA0OD9J2CF+j94hxitaABJ
lmxuL2dSncxG/BmxRCBnpiHy5oXJk7HuO/t2RftZr98tgY19w3rbC1o1F9TrUtRC
1Jlc9jITO9I42vjcotOy/bbCRDDL+VEkBDRGRpTJzshUlX3uWkt3g8RdP4Yj6EJ/
6bmv5skFh1DGrc97FxMi0ows7S9M+VuyUGmya4y5zvKEAbIRGUJyQSCRwa/d4c0e
0pRwT9LSW9j5anF/nYydCLMPhYuHdU397hfYMuUV9Tiv5ROwrE60Nf/9IAepa/eI
pWChO41ksaGPQlNXf63MufW78EjMklb49PBh75fbRdtVZ3fX+f9LsH7iPs7M2f25
cqJ10VDVeD23mLzg1SzlsxV688Bb1UY+nHbGngdRPg3vMZPHrrCsx2t3o0/v04ee
MtUL/dq5RszDujMPX6pId43tGODMkPmgOas57VrVYXN2+Zcwi59Ginr4sIg6aJhu
SgUtGMzPxbEYYG8uW7pSDbQo4wiU1vvm3Ry0eaPHTHA8xiIV5rqMwbaf2WSnkoKi
hh5oDCIQDr7us6YhZICkRyzm+w24lu3Z0cg12NHs+jIUU5GBsdtcPAGSfCwBrQaO
0wisCmTwGXkByV80UbnNkqUsq+AGuepAw/tEOnEweGXWUASrZi6RFK5L76bFiUgU
2kVDO6BKO4oYH7qAEXGGA4D9p+NheAppXoz6bMyCV472VglTFQaQdTho86Hs2SBt
vfxVmpSNz/id/PF3ozmkuPX+Nc6XOkJUQAABL35DLO6Fk8L+92bgREdoGg08vP+o
pSe2obGoqTBSH6n4DppXfR0lzBNMUzKDRzDeumlM4ahShnxNQn5ve65baj19rSbb
6AAa0JPVDyWe0yytGpr82u1k+MygBFmxFHvxY1N30vNV5H7cGwPywyYACqwOBrhe
JTu9uA0dd1x5m1kqp7NA7E4GUwujuSrRniVjA856pqlWTkSQXWYTVsLjeakV6iQw
RxehZOFDetHybZC58rGtEfuIH68azTDZSApmnyPqFJiX2/jsloJBNUX5zafTbLrX
+Xxci4H7QaadxbY9hI8dodcTqabz1qjHVwkfEGEfBQIe5/2z2MsBx6DRAEoi8f8Y
QxGuP1Q9yfrc0kRjKTEU9q8GfGV3I2MIYsqQ9bB1yTbOY+4tN/cnPUR8pgAEAOfO
qcT9ozHtu5lAyREERL+04licjj3X6zu9vlJrVxiWS3Iz0YfXffdHY7VqhvtKcZ9d
o35wtIuYpF7u6fHvQNnuEuXvC0Czr12eUYTCEY4oqQVAdRzgxIFi0AxAOLsahUMw
k0huKyCQmaA6DYxNuSvYCRoLpL1Gvh0ZMASLAYWytUmH9tin7t28q9ye/5C5CAWw
SDY8SKkLj4lKBULuMvKLApASGcR3psdEETny/Jyh4cHj3hzqnum0CgXy1j+JwIxs
/pTux/FTU0eNuHeIrG7Hl/nB0c1jP8zppOXSMG2fZMl+Qxgl/chMqfomLpWTRzDa
POIj3lwrSgSJuEzaKm+hMRTcnyVYJOVaTZz8s33keDCc0IfGzROxvq+7loHI1gAW
ebp8GTQ6AFXRsQW+LXuVsYm72j9bmCIlBRnByW6wigNx89WFq75yzzeokQYekP2z
D3m+bYEuT5A9Y11Uj2fpZc4k93VuUMuCyAIB89zlRJiXqbqEDHZJ9nwZDsB9oQgr
PWASOcWJ0pUMrdWDVFMktTIwTvrtQ0cmA/uVmCs0RXQLgzfDFIIwHFLqjHz6RsJ3
qq7wMr2cF5+6RATkdnVQQtN4y+r5N1PccXGVVNdGkV3UVsNfcPviEcULddAMrtb4
YFB865QDuDBbH2JHaF3dC9NAFYHN3OAgqbtP7fNg0vS9oShf1r9CkY6GnbBq7B0n
vzHcecUGFE+ITfwND0WzIxk9JokLtwtB/ZNdSq+TU7mKrMhPzLxEsUMLb58CMPRW
uhFExkzqLjz3ZWHDYhRwSOq1yHHu0ADGgD8dZcMUowHexgFky/QqeH2DRz3dxmTR
m1Nr6xrUXw5p3DBKbDAmFHzTZKdq7Wjs0aY/z69pnw0GbGT6+pFgrhoDdxSgkaK7
Cpy6+D06wZ4QhIIa8Pd+LsthI1wTHWGa5KE0P43mT4CYh58D0zqk9nlmOltHVYr2
5r2BQOVRZDZv1WMRQZVRoUwTtIQZAWntctknyvYJOZPK31oycOQ2PAvWvHyCoJwG
HSPqn/K3ko4BPNeSCO3V2uWK+M2OwRzXKTNftcRatYNJwsnhnBMYLyR00hsnjF43
HXAJVXkRm1zz8b3lP34ViNn0BtOa6+7wRCVsiAI5m8z6duc3leGNKVYMUF4PGuNi
ReIiJQ0IkX3oXD5ED/oene79f/xDJavMU3TSGG0tF3UDfIpFP50Dmh8z7tGVTCiT
jC4H2vRpxR2gO4EiiqBchckh3lvdZNDCKiQvk5BdB3JWcCQjJHsiAISEt0+pWYK+
10xPLhRJEmIyGfYlxJbq9MBtGy+465tlGcl3nCnwChaWVDwfyZRX4LrzaTgQGbsu
hiWS95nRcCNWHbkfdtc/02A2+fVqM2SFFqQFltsKIBkGOP3a99oytQzHuHZNesxf
Cm74KKGP9fhQRWnDbwU3bBcSc/A2JFydUhYeqowtbHhMSbKgVc3O1TVyHeFBwtmW
Uu+P1et/HmjWj3DxxYLX4q4yU6/WuGx00BX9G62XbXA=
`protect END_PROTECTED
