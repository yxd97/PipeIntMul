`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XBNcWwAwjcCUJ2cz8twvdmQey/g3YoC9Ax3filUldBR1mr7kv2oxBoRrX9r3sd9Z
YJM8+N71fdxaK1tzDJK/ET0WydwKFLPgexO69FfGtF2yQ+eU87IeD5U01EDi54qI
HOaPeOhxqfXPlH8FWv4r6R2sPV1gHQSw48JnKhr9pHOfw53KmhLTYmsXUUeCy2bF
78XuH7OWcXx2z0Ydey50WbndYkQkvARbUnRqtAlTyrm5EH8cj+gzvcnrwx/yur7I
aNVEPu/iuLjJu2NiCY7vjOmfPkekzMeV9EpKQ4yGG6Y9pGrGILsPcio9dGwORACE
0SJAFq2urWGft0B0JN48peLe16uF2fviE7guIXCnxoygjnDxMWh0nwonnH0zVoW/
zGTdZEW4P/5uIA11KeHv+v769A9i5kilg+fmUHBijyqAB1v5zaI5POiKF/NX4Is1
QQuW5MAqbCTlTdtSuALg9atBIXVcKavYes0Gx1HzS5LogWs5VT0exG8KD2l2Uo0q
uPmGcmsLayQfPcVCOOx81T86n8XeJyglcUDCnzyWLBexMlEKAOwXT8KriLwgAhPm
F0wzEI7kdmTyfvS557np0vmE4tIcMc4L+IFMmgmls10J8aqPNHWKoVXuYWf8zomg
zoE3fYhg0zS92+d0rfPg30Rtg6n30agGAJ5rMkaVEi2OrHxCbUU0Iwg7VoM6wnyd
Q9Zy5xzUOd2kxI714YuogDzlNnQlqye8gZOJFvZEnHgubBTSO7ZIt4M0VRD9i9hR
RsSr+LVctF96N7huryoji7ivNdLmgPlkRMTRdnpAd+N758bzS6ktdr7x5epaehDw
sBk7yPFbqPGD2QHvn021KWyJn7zGN9c3a/s9rfF/USOG7avltK536iEOvpQ+6AIk
EQY8PZUgi/MBph4tngyO3w2Ortz/n5KF1IR77o5yORAHrfxuARohf7KFWcfs8wFw
ipbVrJTWuL0cSt5Sj/20oITIrUrN1UMyG5vlwD1m92pzKlpzQYL9EDg7SbQuqJk7
2z3kJvtFDHxp/DYUJ4Ohyw==
`protect END_PROTECTED
