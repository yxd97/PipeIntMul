`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4oO3hMn7Tj0vOSfx6CBqg3qYt07bCokr+J+6J/4pQFZP+z57ymU0ftD7Kn81Te4
CJqvsBQcW1EJps6oQvu9/H87xc21fqoRWRYe2NtpAx7ewGC2oWyEbog/DKa6lS1v
XKMjllQJjIYj1P/jOAykI5vgJGpGgnbT8qOO5718Vt2aKpVRZ4cvb75DPWzxGyGb
5V3TjNIPYQAiphAlbK2fGXx0TkJK84ZOoXVyGjuzt0RZFV5+OTjK81SJcwLqVcLL
h/F4VfLFvr9qs/9cGAguz/xxP3zftYs74f16XedVkaWKjevKR7hULDBTO0HS4JUQ
GQHKcbPFpTMhfEcZR6/D3b9lejqNQeT3CRhylCRxJhlJJySjsx56F3BwkVTqohkh
XYjEzHxkT7CyidsDZe8XMPFBQ/qRASXyVNmFhvkJdMcoMCXhfBoJ+C6Lc5wZ8lZq
T3GBCDTvOEnF7XmrEkKPGf1jBhOu10gZDi4WQZ9J2KansvXj5DAplFZfPQ5kWfRg
xRS7XqxVdYkMC0E3ttCuvkUsYf7CcGjIW9ya5ypBqGgEo8ed6cKSIVVMsRus4qXd
bE7mjBg8KS8qwPbbjkEKBv5cYkgMlzObx+cPsCfKuLhgman7nDCGzhxtBi9Hl6Z/
oEUuQ7OJE9hTv3gpSiz0CPJ3bSXrdqtnBp67HFL2tr+t+qTx5A75lTKHQ7Spbqfp
zX1VfZXhOlqoFJ0rX0eGyu9X7pdYT6vvi52vUAYiM4O1OdW+y8tX8ou87S+GZOSO
WAl0MY6Magc+nYyLl79+YWIm4l+4s2y0nItLyAj2FIN0LMBuWsoDYtGcrgFWWMJv
KjwG7PEW4zdfzYRpYNBzOgPKOykQZY3uMsY23u/MOvEfbRPQzPS+2SFwUzwQxuFW
VyxrauwCH2T0vx8j5+njzBWfaRzFz1NhF+WPhLfqT5VS6kHMjXHUoulsgiqMn4SH
YksBeF4tHdeWl7fKPIgzLYqVu2ua0eFCG9tEOphe84xkzkIRVhePQK0pMfjYORmY
boX8sDTAEU3klteofQP3Ya4hmDeHjVyRxbYo8AUS0ew1w6WqS3GxpTxo+DzK7Qrs
kJglWSx69SuAK9tR+4qDb63m7eHV89idPlYY8mW30zcMvzCrL6xB03QfTQOIE4qz
16F0lfKeZFNTCzCigpuRIVvVvsuSlsC3XF+xSQxqdaKghLJ82KSJNKAGM4iZyqFU
Ma8QT3+JiiTpz+Q34JTnYmdbXCR9GZfIwc7HIoxjShmGcFtSjV0tV+Eb6DZyQjT0
qI/gf50D3Z5iU+DKW3hSxQhHoucPd6XKPGlD6hTS3SNb5eMRQyMv4PopCsm/sY8+
L4a8yu1LBsy6HR+DVxZCSL7hGkI3KqX8rUCOf4dX9vxGKpgq9Uo8ZBfQh9FgNecg
ex67+7d8ekATcuVQmYrUtVvOR20qdJqBCFbE5dGRVvfn/EXQeSJ85/5v6yUw9oqB
Id62My8+w5zSwk+vopmT46bZACm8srapdwp2N7RtW01Bm+aWxXHxOdqGvMI1OgdI
VpT7ZVuC439T8oQN4X5R9+892gDtmvywrZAQ0Z3MA1V3KSQKPCRjcjfMbIgDaidZ
7l5FscayVY7kK0w+/rXGleiSEJkdlnVaxFWBn7zfIibYcNn2B+uLNbJe9RvbuV7O
BeKZxw7VrBxVv53OmOaeSbAGX0bKzq4YLeEqc+rrUFgclrWwA4oI3LDMLt8EYzLT
Ec0ofIPya9YsZZVQfhWyxKs6plaw9QldwCSy4kRdx3eFQrE7I4SnED2lZMbGXTIg
VDzVcTOB/9PRq/mxurSJb7+u+nBe1Nr/rOC69RDQ+a8lMwCFCK8VeToRH3zawMy2
VIp1xfOa/m5CzhLhXFAcRInOQr9tlG9Y0U9k0bXFosmtJI9YkrwnVdcq7ZsnWp1B
Yl+SHgLzv6bbk1vYjAuFpX6DiKiykpkXPMxWKmz46BXcxeGBEsKWLU74KhnP9tY4
xUdc8Za52+FKLPkMW7IT3T8kYm2P9KpO5e5+S9g50lPuR5RpH1AX4xKVseaC2/YM
48goXozBsW+bMrwyq2tUXDBpVc6ILwdaYfGjktpTgB+Mo63czMD4asgRcHnDg1yF
bjB8u4t1r7caX2QiX4eowbmASfWPyJYsCfZCzfGY/1SYCcUkOQeO8G3cTDdMMVnf
eCG5KtZDZ/1FbZPUp3v+QGLlCrGuUdlvskG+MPsB73c48NLq8c+4ZahoKFNI2qBs
PqsBjtInB4ADeZWADX8mBlQcLC7qXpiqOnKlcuj2AFyFAW54Xtp1gRvk6FjnopdC
sSJSiLfY4k7HdUJUqJHiRszbcUayvbG2KG3wOsUxvry5f0IhHn+xxjSylv0qQZZJ
RZlIkdCHakope4tjCX8GTTSNJ0aEa4MJQet/iqGEiGrXL2eMdNGxXUnVFZ02C78y
`protect END_PROTECTED
