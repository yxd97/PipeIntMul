`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOoAymX9NhtYppb7FUqRQlnBIj9Rhqmw6diM6uNx3ZG/oqFcVSoQyewsr+xm5qq7
6MpysfvahUr1rStpoBTFqSV5wr+pN/jw2B4pioNjDRM9NkKv7zkuG9XeX6CJ8Uwg
WvBfQTZpCm/rehFOXvpAkxnzoEt4AYcaCHPAMTy9UItyaIgd4NBWXfmRwLGn/WdJ
Tqmff9yC2AzWRSCiikRYi4QPi90fEJ9iB0NpycOuwzORVuZxTYh3O88uyU1jX4LO
ZuGlsPqL7a+soNPZVbubwZ7xZoqd01o877AHK9RoOX5aWpCamBc1ITrFNe04GPDw
l85moVO8feHWRQgPdKmIzDn4A/FAWpZSl8jHGzOzFJAucFzgiGv8SsWPwnHGpkCm
m1kW1U5OCvn/Hu5XFybdcmCK0v4S7EfF6pEPKvQLCKC2RYEq23cmf6+CFISxQ6QS
urrQSZUFMdt8OfU5+I3KO7r5K9jECpx9sYTdRdK0EUznctLWgZT5FOaXN+6i8ntx
HDUxKyyVF3gr5M/w7L4lUz69d7USKJXBCVeIF7+B46gS6SwJsVrMDkQVFSRdLq82
/PoihrZ2Iyvj1teWC2QxpbQMMEpiJX0deMeLzAvFUGA0qYQHnr93es1ZJZkyVv/t
WX1NMDrii26JV1gVwBG+t4LhrcuML5TmoW3p1Y7V7UuUtM9yIFwXi5QK+VHlxPOL
ewpKXqDTHO3dmcx3ptPYzxWC1Yaa7u9zr7ukppIxRNYN5oWxl6+8V72EdUh37FSL
3HSfcxetOdOr2DM0QPhWd8RNYdiEbJnGmUo7ZzcAruxgMwYnlq/ZBPdr+SUS1GRj
HPbOHpPoK7FsA4Ys+LgrgPFp6hko4dSf9sYtwHac4LET4p+fKGhI/usk9nFl8BIm
4PIJ7scRaSuAzvcpTv7UggqN/Fdh6xt/lE+3qZUOreYHPhg4mRnO7EpyBFzu0Iri
cmxjZYrQp2mFLP5GWVwEWLLJ+19tYgW409NT+mqfsAtvelH0OqVXaVqfHDRW+ikt
9RIVfvTZsR2ocvwxnhN0zGKeDFNixhXO5128RJabQ2DH7ozQ183kQY6vBT7dg+yd
`protect END_PROTECTED
