`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4A26yS6di29lsDhVIZr7tL6nJhWbMZtKvmaSQna0wIKRpli1p3yZpj5vZzHVWmv
8X0rp6tTW6eAWLw6C8S3OxK/rS/qGsYmvzkoA/EhnreKQhkXizRK9RoIJiXoykvq
2/6AZpOX/f2NBm0b54Trj8LWHMCTkKltdNTXBzPAzjbCXJsKNW/69XWIIY18fwCV
VIKuyEcqwi+PMdO6pT0dQ+vu3ndX7riQeG+RS/vKKdnqQbSIlPEZKVkcORXkVyWv
0+wd05e/l1McGY94iQ+8xew/30bQqEMGv69YKv1hTGDknjheaRnCyTp7C2UfWUCy
QutIrNJvXO5741X/my/96H3eeEk57ntm1rUuywz0Rp76t+1xCujuFwFe86uIoxIx
8Bbrq/bA9ZPzEZ37qQ78lRgTUYqp/Lja8svew5fed+D8T0a5glpdoxKwmOIm8Jml
Q/vDgc5yTqhTXCtgrKPBXGNBb/XRSbsYEu8qNa32ouCEVbTFP48jdBrVyhGtJsuy
5oraqVvOdlYedRi1qRhWxvjPJ725gacwa9hIdGWcc2kdEUC/HaDIusreeBRJ9gkW
S3a4hPySUO1SagrpZDjfuY4AIivAxIob8iMxuKnGRRYmLUXODpMShWTdYTVt6iPq
giQE4WBesTTrqahQotoCpdL+QxP095zqWPx2rWMMS3Y=
`protect END_PROTECTED
