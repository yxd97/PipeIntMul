`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1SRLN/ivcaMyfWe1RieLJBcf6r5rzoEPiCxfAxsoO4SoUCc9Jvi6cWmXBZcdRWoe
VGu2uE0qMfA0JT1czX9sdfmTO+Dt5AjDgs3jjWGFkFu1UBWMAKigjDWhmGKHwCF9
hZFlPgy8UTWVyE4xekWpKPJ3VUpQyNtWanJT5uQMHJSruHa2pBFPgRvoho0joOl9
ump6UdE/B1zAXtnonG/ugC7DQDthI3CoYN8sX+LPmu335BcfE4sA2DhXhEoPOKPc
YhOrzRgMYmcxKLlsRe/og/kCjGYDsq2YikLDFaoaCJlvwde0JKvgwLVHxiGLT+Hk
DSaNxQbkZG0Hj4927zhCkbl9gW4FkhecqgEPfzRAfIKGpKR8+b7NMwIT4Ow4qq9E
B5fMOO7Wwp6RQ8n7Z+rTbHd5SMT66TQqhkdkvnG7MgvTj8aFLDnPETiqDC7ZQ1MR
oW3Grw4g+/u8bYH4u9H5Vo5QlZ/2liHTLVPe6w+8dajz+WthZN0CfvqIr8YyAVug
xVTrj2c4emUgKENcI+pyDfkX1LagShOmBTasopiNsJXSGuYsIkl507HieNLuT5x8
Fwp8MzhnY/ndW3siDqkDWvuenAUHN/f929pakS9tAHW45oWsJR8V5UrRJ/SoWx+j
gjUOdgiTrDIKpobCK9Ud27vlfqcmaiBtdUgZIa8brfqYvAVkxesgSa2ySnaMMr0V
qxx5opDUn6+7LlJTTnDSpHyvGV/Cu4M9m/jF0VD7iS3J3CFXsjAIgdvN3uDOI7cW
lvikT6a0f1bgCQRsPtiaGA==
`protect END_PROTECTED
