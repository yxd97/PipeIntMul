`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRJMoG1fhtf14lguFCyuZiM05oWyYjc/I+Gwh5jh1Avqxkk/R87cAmtnHZYT/Yj5
XIAwMSfgShGx1Xpjqay4Aympx9GmotI4bKAIPzD1fBNoufUV2sUQsYapyujtnGAW
YsiVPj+zR0aywHZRfcOJePJAwv2ISWGeW4u6Dq/fNdchh4o4sMfOxYnH0LvF6CNl
EEet/HNPDbGxE5Tn6LwPsJE4AKCkdxGIzCf4ma+q2YUONqPP+BMXvQWztrH/fVxI
E2UVjy93OgSXUFX3Gxz7UCsM/53H4vA265motJRsVTatCws1DPU98GUpRHPskIrE
TD+8+qS9qf0GxjwIktu2X9pR1AICL9jbY9/ONNUaQV4RSolYGTiGdQ10OjuxiPm2
fjYyEyoIdngMRDInTss2CHM0a/mulpeg+odJW+Uv0m2hZbtxz81FTsvQEcQdNS27
3bMfn1ay+w5ni7vqUBKvJvOBGb5f8eMoxqG+meEwXOFFIe3p3Q9wyirBxAX+HoeT
M17UuwP3/lqvIbbsAIZGqhKRoYVBmCvl446lIJ4uVV88ggdt0LtJw2hsPWuH+4Kc
99IziJSdpdHy6dbLcT1l6IuRq9Bunq5D0/lHJ/jmyV5sCfxcfZ8FGtuZdfuRunVb
G9YQwxMwvCB/xpcjeATTbQIZZ2tW2sTCPTfvl/ZvVIygaj+EiRhDIYmyKjZ+8+R6
kaYuuzvPYesvtm+l8eigq2jdrPm/jA3aciHNRGMDh3wYSC7f7GVhawPy2cFTxvMr
yjT4yzAfetoIhxJf7BdOkXr7YUQArn4KjdKYFv/SsrfLPK6+eECzWQpdQ67fDiIY
nPQsXf574ax1zdUfCbzxEFLC0qMkzeTqsB6iti2DqJ/ylEhagVKRSRNZbdY0G0if
zIfRDAbFauqC3Qee38aA8w==
`protect END_PROTECTED
