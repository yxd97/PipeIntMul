`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3ZNbawoH1KANfKyq8KL4IUM3byjuq7RSygRp3KOm/CfDmjusIQUId2iUZoXWleX
1ZfFKJvp+G8AFveWkjTpnAnZ3htuwjTsTN3/hRUm1F5E8MAzR6/lC6Imcp+URqjk
+aGr76HoQrHi5sdNCIPcOtlHOjTgoPqTppiYBrkqzy36sNN8LO5Bp39Wit8Tnxyt
1VP10oa9N8gA3mqpvH05N7R1GZPIA+SFm1iz3bUzipAXKqEcwFOdoOWKEdrkjOHC
5UAjwmvb/n0VCCgF12Q67R/S2/BuYfbeRN1TyapALLga+JNL42Cts07mV1BFowa+
YO41ZkSraRLVlFyehtXppejWyotzJcQQpY4uGWy2vhEZ7brnghFvFqQsxRKdqysm
BaYFXOcSsZUUaaJUMLyS8Nm+aoMRnpAFOoojGzUBzv/8UISNN+isuq13kz/61Q4j
TqiSgIskoLtElzHIM0uYebhZ8+VSft7Qpkh8+VAUc6+PSN1REfOdTGUBLXJK7MUs
9qv27FKqcU3Rxmf3cLCRxi8/r9Bpf1sncB+YNpKO58snHeq9egS556wgZh4Fs/7q
kdMPNnxbfp8I1TukBlhgTEyYWQvR2GJzq49f2sUM0cewzPbNAGO8fCoQsXDLPWe7
sTVIlyX79E8fYIE/TWpCxWlIeo/mnCNsMdIiEGQ64zgDNJ3oKEVD2KyoOsfKHSPG
XDksSWRz3gy5y/JLmMDQwN0D1hth/WbblaNt5hQLFui9x8LCFet+pCjfkY/7AlvS
gYzmRwnlTHBGIZejVEEPKlyMpKGPP5Z8kPFPUwvvTa/EicEHkCEtICPopOrLKU28
MWD6Kvy1tEDYYk4VDPv8vdsi3R4+gA7FnE3gVdgb6e13W/9TMdmkignO31LByDV7
BQIqy8mVLU9y4Q7CtU94gGGRywdV3BFrBhGWwUkpR/MhMC+GAFn4/Otnx7xgYoGO
4eRz7MZKEclzKqcn0GqJnOtSW+vt8OmFGz6XVMcga1FPlhKe/MzM2lgeznTdlfY4
6IroNpZij4/tzhSomoq2Py3kE2Ygga/Co9PNJcK1er07+dYjW4hTueuplgW3AdJS
4Ne66MURVRtMVzisiAv4sQ==
`protect END_PROTECTED
