`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bX+ipTst5C50CidOfcvRb9UakEp6Mg5tr9pO9fnSPKpHGzOmg9Z2j7KHwRitYk8n
ukYfeofpNGm2gWAYxaK9F+vumerKCUfoWvL4Quecu3UAWz9HWxtBGAxfIAtMTK4p
cbrVzIez8Xj9dwB+9LtmF2/+8pRNsSRLsVDB3GqL4538k3/rVMCjWdRBLOOgO9Rc
7wlRriwe5YGbM9gtktwAvfecouLHkmlqMVg3o5ws4HXQf9g5Ki/vxqjaiZGTq1sh
j1aMqydTsE1pbq39QLV6KU4BVNxCv6VKR+Q5GyAwlN8idMYhdncUMtHtWEtlkvfo
GfzPglfhgp3s8UTYa0hhodg5qo0h/gGVMJ+z2GnP70GE+GX2HKH1kz01jx0QKkwt
V2nJXyBgkhcE5qLO9lM6mwua3xY7KOcpEUNk9x/0l3PZIZibiqY2xPXaLffGWmjK
uPXfl/HdYwj+8EMp5BShDdpZvvIvGPiMMHPTm+be3DQwyfE+RTlknwYzTrEkIL0Z
On1pFfxjPWpkYKlaYpaaf7OBoAwwPna5OZ1gcBJIcBIoloXbAfmAORrmkoE3urIn
KShL+9tVghQ2XZQwtQuMnAq9x0BwCXApA0lS/k+IBzmHdxHajw+maEpJd2N62lYh
puzg2OQQOI3BLQEwFqlrYSg39nRvMyZtD7S2R5qwIO6F8tf72Bb2OYnaJReTM9fW
cPnfgp5l9gHYfwDD1VOEhW3BSB4MtHY9beYMItCc/9hhLErIGJfzGA4IxNzDUmRl
BAT6ljmP49f2XuQ7zNz80jKWSBj4w8KpKgTjVYnx3Ocji6flGiZrDGiu2z2FYnVB
R6XJtk90/NvN8G96Jb45bM9JT1yyI5enQZkXnR92p8FPJSN7ay1kOBemBooE9KO6
ktvYhzzswmQV6JZMvttz3i3Wv3AYefBvOQvV735uf4kdj563tvTyMIA+R/lgLkNb
OgORMnd/LO2kKAs6MyfocLV1kEki7uuMgoOfql+YtYZShHrXow5e+0rY3I4LhWRo
pFLt04j79ha6Fivq040PDo2NthzeO1KBrzoIKrlJMF5W3elS6O4IvtcGmIhfnvaf
f9NR9do4f2xcD6e+CbDavilBlL7H8u2HGB3CZM8yksKPc+EYpXtbpOgNHiihqD7d
z/aIZaz+OAU/iaHJB9NwNaDoWYW5DDp6b6O5eXc7Ms4GYxP7Doiaru01qcfoKOzK
nLRt2gCyWxt0mdhv47Dm8oSPeQDuoCcvLgDRx4sPvrWOJSZk1D0B2Ij44D1QbSR0
oh9jyhuXpDkYuCY89F2kuoTrUstZAPpET8Nyr62A1lE34tc2z5+jr9ZVAgT5wjiL
RyUYseu2LyaRfELCXi7koRbEo+hpvwJfmmqk44tTvsE6CZARp1Wex1wRQBF9TlHY
+GFbYDJ2AXUSc55Cvi42IA==
`protect END_PROTECTED
