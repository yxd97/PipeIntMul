`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sg9sBWXrKVRVqW/B9sg1qYJVks0W5djhyedsMLFoQ38msMlOHBSw0OqRFtqSkqYs
pb33Fn2l+sF4wAScM6/fcbYplFlNay72ycJfvbDTnpNtG35kkH+cCwoyKId59tBk
o4PCw8loW2w5134UC7UKZlJqhU+rdwhXxk2FwgWTrWQRjx3tXhpFXvZD11VUJZ5B
AMvOmtM/JBzlt4dP7tYtihVMGAQvXCPiXyt2tqmZRK8aZUMIRK7yuc4Tz1l+g76S
Djx0X2Ukz7atM0yOqAqwcjHUY3rBrZZj6H59B3Q70JLk5t6zdVqcUXk0xeC1mbO+
jMytxQBwQZsBz8TVOUiGcrnvR47Irb8R+cClQ5RllX+hr6rsPr3wpkl86cwAcjPE
RvBj0viCjMtnyMcfpjqdb2+AIkKLI2PMaHfNev9DQ8mOlsqRLZahvkviCdtvpqVo
q7zB9y+ioEmIwXsxjIUsMmpaP1sgBPqZ7RXP5pZWDx4=
`protect END_PROTECTED
