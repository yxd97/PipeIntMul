`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdaP1C/i7f7e35gh+7WztNZu0cgT53UInUg+JIDmFNqcNDwcWjYafESOCPvE4rv4
XR3gnt49urYbF0kykpQuiIeK2CRtDIV007YXY77H/ORqS6puiY7V9LQmhLca4WEQ
SEulWKotM4B+H0xsBWc3IHEQOF1xhHqmPjDNhrvJ9V6Xa1nyplnhqJCeLKo8Js8q
f6TNHmZZUJz4ScpyVo85/cEh2P1zU+JvXZRXfApailTQXP3dreEHQwQsXToS/P2x
MtZTeKIlQ4o4ITT7evbArytwwU+7/NuoJNGLmmcT+40RnMbkHhoyfy38UX8j8Vyt
QM9ehVyyGdhmHyEQ8DQLa9PyZwa/4TdXQglWgqSERWjjs9MPWPNv/iCMD4CXWJYy
WmwQ/IQ+U4JOyOre0lgc/D9Zkg+qt2rC6CMDMqi+KCmn1ougmZVKcdtsEmRrElbZ
2R/KWgshWVQx75p6hC24pQie4CbMt2BJoNCfxxA6UksGdY8HkGG2SZPelsfz+pWs
lZkwLnabuOlnF88ahlrKGdFg6L7zejCnz1w9Pbky6AH6Cvz7fYIajKl+7BObofIC
ETS2Qm44AwI2OasOCINzIjqLlKbJdNY/aELjqW1iCNO2KWyrN8ySIDtOfAReqsSK
FPLbEtORdy2sPi7OAAfMEwZn6SiVREiy8198heyR1imhv+kpFzxrPoEU9kT1IVn3
Qr8VP3bnr3d+1LU6DCXm4yLOX4ObAL1mYOB8vGtSV0pnqAg1uD+rZoxCPrmdq4sQ
n/iy9WIDnJIos9cGEMgRmS7FJxHaTTVojV8xw01/8xrTvFLFW/XGQ7NC5MYO7vwf
PW0NCUuqT7AmHYCbX6X6Xmq4/+oWhyAOzeMSte4GGzeaC4NasvbVXaPu0lStt+mG
seDO9c6hPr4SgXBTFWpd1LyjogdOZnjvI5yTrJ2+fsNVpittGArExYw2YY67hcGR
er1Z7BpPQzorfNPI0g2Vl3idi+qurAc5t49KIbU9vHFxSznKbY4fjnB8avWMEdfx
sdMJx2nQ5+BbCdKZ682rUsMkhmehKVRHqbN1fy5LTPAf+Cn18vxzRCE3hICySDcU
02BEuTzB8tvH21EEb4tfK8YuXhyuOw/LbOaGFgpdUlTsNIb0yM43O6E17nqMN/ps
gtT2iYCjgrFOQBT/geYoUeWxiEPXSWe5Jh7kLuTBDCsto/G3LESmC/H/6KJj7c4W
aciHjlpAGHEDdgzqsUa0xk6/HxiW7Bl2QqpYpe54i3nLDgd4uw3qKYV5HrW9uD1S
4qEFjkj8G+xFTwOddThHt9GYYgCQ5ZyajhgAp1VqootFMOQ+yOylP8jBPo67cyQf
sdFZ1kNfOJnAIG8NaKhCT0oq9ZeIPTqyz3/H1EHmEL+OAxJuH4eME7QmPIdt7CgC
yhoYrSO68g8ywCj9mA7dmYU8XWRUuqWvLz7S8qTZKhE+gLTZR/f9F5JY/mr9aTpf
qmkddPqi1BmesDDOmJzEM8Bz3s9uApnCc9Pgh6zjrlhIFmAwQfKZB1WsZWhOXhSR
FMXpx97M0Mc/DRKdmVQy4ghtmm436A9UsvCkUnEnsyYdi1c4hD6RIcSq6GqwS2I7
h5ZA/ne6gsgNT2su1W10OPMVs6qu5qXCE43q72/OwIOib5N80iWk4+TrKrQ0Is0c
5ir5d3PN9XEsXxYfgGI771MdGXcFFJ1ZQiXFZbMDnKO+/dE8WZWv6dADA3wswN9b
rvC25yn+enHK3kSkYVc3pa2PzUaxOx0v7IiaYJZF4YEhYhVLkf2YSHtq961Y8gNg
ZrIRtYLjNEutfYLBhwNbNz51U6ZS48YaXEeefAAauVWAgCA5vN0mmDlN20r1vZPK
y1jaLfNsO+7QH71Ncjr7s0IxvF+3ErQCifs1VDcMY6J0B2f0+hodbyc/qHWzOSPr
521LLSOIo/3pFcyVDKMFgvgRCwJCqGTTfruFvtPJMDRs8C86jm1G5QQLCC2lK1cc
fHZvz4ytvlAwAqDTxZy/H9mxMRUq30+heA9YT2dvS0CN1HoaNUi/xljhH1CYuA5z
D4YMz1PGdjHj/bXOmKdRd/9S5BXgCM4vBCRdFE1Qm7ZO0DjrTNraEDAwZ8Yhwtzx
bg88JqMnrWo4YXcW3t+zeFy7vJoOQSROHBvA/CBzp5i44jmKM7tdQgmRj0HyagfI
tJfsvHTuav1bi3rbMAeJovVvOqe5dPA+kEQmp06jX1I=
`protect END_PROTECTED
