`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l9GmBe3RHoBnln0Nl/7/59JClEsOFt/vlhOFuGWZxfBku4TQz1SrMLC8/HoCWz3v
7uwowtu84PlCtjcVfR1ouEPukmiCbz5Fo+32Ilesq36BRh3TG2MDAu4xz4uIgwfV
I4YkA8gpDs0bz7UMgCasK1L0kywssL4j1fy25zlnXVhZQ6r1VEhIOWWw1jGfdqtZ
HZpk304wm5+nh4m3EH5feeeZ4oWbdAXxvdlXzX+EJ4qWUl/HPf7taexwHaAC1ygd
`protect END_PROTECTED
