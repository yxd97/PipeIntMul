`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogSXis5TQre/BhosU4kpcMwFhAmZsE7b5pjqoh/iBPf2oHSQgXjvqwKKkhcXVbvT
xnHzHpM4FQ1HznHsVBZCF7BgOn0z1FRQ/bGXrf/bB6qQHTQN2nq+NYkbuxxVREjJ
o4g7BdzeYYKrz+WQC0KfG26t6csAYR+oYc6ExZJLLU2HWcib5B5D5qKE+3V/jZiu
gAeeIuCGK+V6F2Yyha5OmUeP382lsMQy+Wb8Qk6iu/9NGgu00wFi/7pX6VMbwnOm
eZKtGvKMaHngT3h6WdNdos4Ou1GzdDQRNsvYLiNuiKK6FD4DU/Gp1sj9iD445shO
cx85E+nW8ulwNsnwEVNhy7I/aahmmI5hGR6l+z06ABVtE9k5GUpPpMIM4RCr4P04
IUoY55EQP7Qwlrk73eOh8Kogk0DGnPbxRYE+lUMUxa7JDBj0WcmJk711eBoD94xh
Af3ouL6CjPsn+jaVLU4fv27MuqxdYz5vaCQNF3MJ+J0=
`protect END_PROTECTED
