`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLcPYZQbCduF3Yy+wJ6cSrfAOUWj0AK75fJoOp3sngQwiTcYpqR7y3hgydWeHkGW
QQpxCBhZkoBlySBT3+qGAHRiOzijXWxYNQd2dDEipH9177tVtTJ3E7AMlOkbM8NS
e9Hh+BZrl8no1E9WkeHlbIlB10PKCeRdqSYuo/OZbW23DLvq0yVXhrMQ+NooFXAM
LZLTH5hg3gPBodhZFRHmFjxHnI5BSPZ9x2tpb9+YGX3WlLGBWDHtYXF9vgqDtYT3
6LS4w1F3U223ZzRgQpSDHwzSsF1LGkliD3u8a4PIpjEQg424eBj9+9w6FBkQiAt9
mJmsVeFG6agNPBl/bS45VHtej+rv8rVFGSDafwkrhUqrkgej6qM+GRO6ISZ/mYKT
U3j566i0MAfwbvJBTgPyinugCx+3blcmwuJ9jwtNxE6pWThzDh1HVgDZ+XJRmZBJ
kMy/RjEx0Pyr8e8qspl4gseWJ8EpRUOQPubbpeHZy9m7EhNcLwZF+dtxKrgWFQmn
PwMEAaMmCCiJqwuIc4lNPNzUGuyQ1WF9//6rG2a3gDneJWydJK7cJKwllPiNUD59
96JSKQ+upHxcW0YuJGi4vg==
`protect END_PROTECTED
