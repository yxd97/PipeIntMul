`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tm8HlibYgEhon5iW5wkkQd4Sbw1a4aqYaLwCrMzoL4bg+5o6hWW+o/TZXOdjOCNu
/O18fdtFhezi+i68ZR86rZJwKkg4va8qJWJhgq7LQ8CHFcPeULrAy+I3VRXDK/H9
Nsnn4C9KaoiRoox6NbXfv6dEi7AqSoB3iUuoQUqWgqa2if1J2ZNkPaoxCR3w9QJz
s76dSyMnVhh8YQ8upsO+VNHQfk6LaEdf3IHERN8guBbZLCbuCu46N1Fjqh4y+lx/
3gzlGeDPa8z/aRWdHG5C27ofTGNu4jeWZTrRQMMxsZMol5+Q6ttKoPl9EJBFnYp8
7R7DQlsNqJssf0/msq/MLEI7YcOJTZhbqFATOSP8OUN6YvBnckqwGywnvnI5q6v1
i76v2O4QfYYLX/riWAfrzQyuBhkb+hMDqU6kEK+p86uR0Mue1VWu7PjS3vcPB8lN
tVYzKc5SNuUtUaOcow/sZCVoEWVwagcz+lF/e9rCofCRVSkqKaZqpETdr/ADT0Ms
AtTi8wkcUSXBnP6lL683YbrgcoBSmotERA9z/49EVHIhKq8O/7wnz0mMMjkq8IDW
Hrl9X12ThvZn3Qu2JCj0JxswT14HrcKSAXIC7B+7mj8sbe3P+slD/zapRnKp3D28
Ndt0eCIWXI60ET43cCAv/DfmxFs5sa3z9kaOeFXK3auCnULDTmbw3SdX7QX16SXW
2gLIolJBxSl1qw+J6RS9mUbDILVqzyKv18CYN7PfZv12y0nsU3wlDn9n5GG1wSMD
I1kbs9R9XcQ0Ysr1pv0B8g==
`protect END_PROTECTED
