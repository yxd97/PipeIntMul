`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HyKnwCUm60p6v7qalSSRL0AQeVx9rsXz1Bgn/Jrok00wbunJYw6+bCPKc3tpOZPv
JCA66zsQiYeSpFWtUflwjwHk/TM3EfYpoF/SSLFlQPGCTF41LoOSWVRQv5yuCFBd
vEQ+ShPSBhC+kiAKLR5z8knSRZnU98wNK6RzaXPBFbfjL6ZJte1+FWg1MLTfu+6O
e7uvoWdAZH967FLXvKpcXCcHIrpe9XTFRK53l2mOIWWNPNU7BgmEhI0xtx9GDzh1
jLLkeDGJFP2DR9h7NkvSDXa1iUEsEsfKXdQwmj5/VRbahMFKNcn3wE4iV+kjCMBJ
Zg1td7zJPo/oxFrnYUpVu5eEtWdmaQGj7sHGHdAKWZHZ7TIsQcQVHxY7BRrJVYw+
0JBgDmZrNR+wLuzqwi6Wwa2ygd8Aeo3XnJ6N+8gofrvm+qMRJI+L3+uFBFdYYNCX
DBL7RW9Kj975+5HabJifDw==
`protect END_PROTECTED
