`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjhrdW7iH8qMkLLsOxAX2FvYqNnSUwOwVcKw0h9IMtgJ8ZIf6YcW+kxw6q8xw5qI
yuuKQi6HggCf9LwUPKRxJQFBkJt199rNZJp2TxRbpnAc9v8WH4/pqezCMx/19pYJ
Mlu8T3IlLv1c79s6+S5YM1iGIFKIle/rBsqGnMBJXCyBe0+4rLt/0u2dqMT4O1Mw
yLUZBqQoM6MFEC/Cq8uN1CuQ1AyOYAuyqqk1b6fLZl2AR88qrcauBbQ/XozGoerT
C5UwLqTt7JR4nGfmVGVv/XRA4CuCPXMiTkpCpCHy8srb5fPHh4Yh7lAFrrWrCMpk
A0tLGX9YgMMvqpbeVKWc8wf2kP3sMv+J/sJl0rFMuO9yrflIKPgzRhBikFkrb5J9
tmpw6oEahlJM/CMlpZ7DFu0Q76AycqamHHxP9qXBwv8khbRXnRTGGvaEAeK3cAIo
4U+US/W7RnkGW3NxyGE2Y8u5fZgufta1WDoo8jLOkWDbSfwEcM1S7F0sWQEl/QZN
+Vaio/hguUwIm2eKsfsV0Tl5mu4kWb+lbb4OTZdyiKRdjxy+4w0h7xuW+oxOn31Y
3fO4YCVa1zJ9dsSVFyhuQz6IzRY+mpGPDvS7BxMi26YBCNkNRvrfDqjKtdDRLz4t
NdmZspIQVwmViwWcKMAp6tJoRO5s6uFyW5uiH3HBE/pIJwdgq0+JCVf8FZnCYd+q
N3IwhEeq7j2OnpU6doFIuIDlp/l3cjRBBaKzDtyMaUDWGwaTIPbTYLPV+0uXtTDW
NOvwBj8H8HLOxGoKs50Fs9jjcetE0yMDHF8eEBcTz6xG2IyNuXI8CRSQaM3WMad2
FunpYgIOJ92Eamzh5NahADQ2k+nPsLZZEppuJD8QDVnDbQQ2ioqFaQvTsCH0MqcI
rZNGqYowzTFVsojZ5cmpecoNQLPc6qD8pujb3nCMGIu/e+3JGN3st/WbnekXyTId
gbz+6SptVdPuTznWRmadRzm1hXdiTjDeYl+fdxZNXIHejcC6tRFmRWrEhJMZ5E95
x9MGjlS+9GEteu3GroDm9n0muBH6l/YKvt88x8Vol5NOg41B79p4FScwimp10JVy
qP07AOLaWUb23fxFqc5N9wQxkwNwI4io3Bua6ZUa6ftq4FOBnG3knKSc1NCklq2s
zYIjoOvD/+lO8LPNV+0omJPtgsVxLdlwIi8eLRP1jrDk6RDG+maKT21eLHmKMDoW
B6HDOFHRhnrnQmlAVhv6ZbRKIeBe5QNt3z0cXvj3WG5DiJtbboqll8+CHMkUnVRX
w7E/l1z8/YHKwhLCNA64rQ0eJctE9jvqhrcjkCd9jJmaD1fd25PH0ECTmbS3Mx6a
ocEoyIW2pLmmJtJAKGf6dZTch5KFw37HFMYrsC85O5CBVzUQs9x3ZLny1YMmOvpo
r74KTjEMJhiYyNvBGU40Tg==
`protect END_PROTECTED
