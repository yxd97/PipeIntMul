`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HiuJCJk/aCpioSYaftw1W+tKUOznsvqgj+jQe/cte/HuC48AaR89mbWY9H8CYM5b
7tVSxnStYT2QAleNzp4hhFu5wv7Mx30Qw86yqHdhCFSQ1Ri/NF1/OdMYHDxsii6z
B8/sftcthsUHOdKtStsUVuXSIhKvgpnMiHiFA+TnFmkOwjr83Cw44dT9i4E5NlAt
HnG2gEl5Sv19+PmmHep5oMbUkkrSrn1i1EjK6ON0VPkghCLwtjbIKyenDfQSmCbd
Mu4fuYQybnLBrua0nk3iBfoLTvoT3UH9+ZPiVAZlZZ2JQEkcmZXd6g7p2GPMgaGT
VFFZ93invB9lZ+4sVOJx1Zj4xlXvDW5uKTAZB4Eg7zuKfuaeDUWApvf+cD/y4nY6
ztp7HZ7DPii5FyOmmO9EpW1hYTAg0xNYHpf4ninzoXYORqADKX79nOct6kdEYwFX
QD5zfvZ1Hw9ecSa54xHu6Z21zD+dzjX+GILZvXChFUhdAgX/S4GIu0qy/8MebMIV
yrolfNbK8FG6nIap5CsdTcelhH7pu2ubCT09eeuLOsrbvGQ7NJW0rb+atVRRc5Zb
wUl5xAbLv6G5k2JgC4Yfw5ZlOvLHdJ7+CabpM50jY4EmC/gKFY5D01/3CdUGRJCf
Y7Ok9TsP21IlZqQs4dUDFsw/6bh032NIlKSIm2PtkrvpPBrzns5HQjRz3EBOjE1L
Q4582RJ29nP3nbMjg0kBnX9kb5ze2RQ236Nnk2ou9E+DYYYL0OBVzMwXs2VUY445
iEHisVAwVG4Te1dY/c0ug9fwx/BraL7yiX/2y9sFeeiYiuTjp3Ybx3G9m/S7v/VC
kRX+K7FusSHIboInrzArOeeCugRS72V8YmbzSkiVj9CWqhQbJEM+62U6cJ5HwdKk
hVIAiM5aI1k0TDpKXIULSRZqng1N1sBp0iBhxb9mceX0jg79DSMCPjyMACReKWtk
FpzKeKOcGeIWjLLNWDt6rhod3qD+Jk26W7oZ/Q9Q/9GMOQkvCVMXq0oqGB/8tXac
yW9/R1EjahxvFNsB8j3DbAULxXAesTaSiimb3s21mI1cp1n0lA6KcwkMIZSAQp2W
TM444dAEomn1x1l8JI9BqarrClv7yg3JfeElfa+mt8+P4O7VwtCyRmX0D/fK5RVZ
59rgvzuaWXsdg8270yOQDR7AuzPAMpEAwzOjC5Uc05YHWeHSe+yETn2D+pp2n53i
9Bd8ybtcQ87T3uGFwsv3d8JUnivcd/7Wmz3eVaf5P8Qppq68qOT4igkQPIEbiegs
HeUf9hNMvn/LkdlybID1vKntue2vl9LbbtWFnbpQyy2qzg0fEmBHspgVT77lAEoz
g5ntVsLKDjhZJOPOa95d4Si0RvwTvETAyAZK9IHBHcR7l+mLaFy/5hULCZg5fCk4
4IvDd5DCNJBuifQICOdSApLDlBzNY4CS0Buz3oVrB0UOd5D9OAayiUjMzXfpPijH
nEvaYVYjNER/Cw9HgSH/8xHMj4OyypSfgrys/3189VqzjHv7F1L4/NwM0MxNCBT1
Fi+anHYPkLWB1znqZaW2ksGT6FPnzmnyXRYJAgZEQ2thEwJBhR4DW5hAPhtlz1WB
6hsS5D6q+sh0RYeTX0c8G68QMCE9TWJ+d/liT4gCxq5UQl9/6AzVAmFKTQ/oU9r8
j18K/DhIhvwAto72tEunzOW3h0Ffrgi+qd1dcl1HbdmW7xHknN1mt/+QV67ksZGl
GWvQC7NDDUsQ/ZZXO5RqZw==
`protect END_PROTECTED
