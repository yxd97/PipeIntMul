`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olTQG5uhL1rUJmzuwytDyWblxLrtbeTtsmFxh1vp15TPg3ZqjuOM7CCA8qsfR9M0
QbaXwk8jvNknYuiQmQZvz8s/AQjlBLIYkZ3ReYZH9PNu5CZRyQ/JzRQHByJLf2VE
epY9UgpPjUMqQLCZRrMFk3qSQCZze7VMa9CF29yPXBZ7AqI88de33IarMtnjzo0A
Web3eAQvPV1C3xeUC2/ER/GKxdWAjktf3XXvP8vLbYndpbgxDRkzWGrJc4Q0ShqU
eESp9KGilskp8WS+yn70m5rHYdnevjLJFITZgGSaQYSstyN8H3bDM0WHgQCTnIFC
b6h4bCCHtnFbZF7yaBzf123Z+pdYFU00QJLxdrrnuVQ4KgRtH3OG3ydL26CXnIIf
VNpdA4wgAowlRcHg8iQgEcuEnvDH7/IRxIt0dw4lD1x5eph6UXI5aWvCvpoJ0Cif
6Z5fjSe3nS8i/YUFlnep2tLgiIF3hGnEngNLL42HDhYZGwVL3WNyUBLbQVe7cyPi
iwD8axuYo3Rzf7tufEcJmVVPwL8o2Hfck26cgMOM5wHK2gteXXw2RRMsdX1uZa27
5zryvTEDKZAWn8RMLKxECARoUS3jZGrqzVS7Mj6Q4U+kNEkXCiqvlLeeQDEf+qJV
SozsUvPP2zn9y2rOWX8jxBH17pzLnlG7K0NIuNVRcInNzvksPMNv2LHXvkIERFTd
RJiH2TD2s9MUyFEUVnCsF4J60o4x3+nBIrAexmVlCTSrHgqQ1Heb6R9px9EZmfXV
siTu/u1RTDFpdOq6qkJbygBCi6i9KEc073Cp537c5BlzbPMVqvXFIlM+f0q0sbrc
01CvW0OqDg25P+bkXXEI8Uz8sPhF85P2quCr9qcrpisntGFD5Q9LmcrYYzFH0P5M
8p+/daCDSH23CuLev0jStHGUUeLJcZIx72r8qE9a2lLcXCs0lqv8SpG4J3vwk8wm
wv7Tfmkv4RKmNqdwczwolQbNKvdnzR2OpC0QyRtFija4nPyMZ+jIEtFJuaX5bYVC
RbDW3KeZD3TZGhAISmrzF6RLd4ypfotL1BLE01yQq3L1Mb+fV9gXCKfeXbwdPKbx
HkIdWimpzL1qqI8cRDQzTWW+wQVhnJeqo8+z+S9+KybEWOHI7/ENcAE+Kdm1JwNu
5x3HebwbBe04itodoTIYQmFo7o5wEV75ibw0S8ZGU36eNspr5FXgjdj+1NwPYR0C
SnZwHkpdCSROMNNPnUx8hnni8HR9GUvwEc/iSFR1181rvc0S6iqOhVQqdGVUsEmE
gyps/o7ISN6EyeRUGdtqNiAIGeUZaZQ2ixNu2fJuC2DCb1DWwoV8+nmHDhb0EYlF
QuLKeL/8ikqSi3fkSMo+wJkuHYPOwi7NlB8TIpjrayv8ubuY3Im9yxMfhu5SZeaN
0q5v7xJnunZNHPr3SxD0C/nnBe6+CsfpbGmJ5NY43jPkH3/pioM/5yVmoqFePbeo
/Xk+chPCSIqbYBLR66uKwDbfPP0pYJAUi6dPU6y9T7wf7vDvcHMHqr6Az/4rSmYW
CTXjywENS20zQ6Apca6s8aYyU6Bh229W/nTw5hw3Wz1/cw+DLdagdg3htRiuNOsw
KVFK3MOekttTCJpm7V7lK1ubjtm+TkIvlawpmhVTqurnWS+Kzks7IBj9c1L/UrKZ
0tZI4gl9YcI9/hbAhG1VcdWcLVFODksFucmLkYJekOCbhrn1uZvUIAkbH5NdeTR6
CAjGHSy5/e6/fgL04j4Sg/O7GbTchpNte1HDsxClXscHT1nm6/p/uMeSrz6lFNWV
561D/Xi/cIRcuPJthNg5rBDsTb46dxDaNQnrhGl0IP6gkz4jxBO93V8lhrRDBicm
4P7ojoRegJw+V3CiASXAsf8Rd8op3Xt+XWATNHvgLoEE08Ylp0TX6pqePB5rq4ZI
MQmrfDfp/AsCZSJmftw71V9+rE/t5X4EnnfZQc/Dk35ubOFF9b/FT8F8zhCJyVDx
tcSigeHgltiF8OdLM/jx1yYpLzr1JVOV5mR/EzEtga7pC/SVQyh6JzwLaN9rXhoO
CPHSKO/AEhzTcUOtZQwu8KY9O4CJBLSWnJIYKd0DyagS9dqu5gHwYXGFhdmUE0DA
D0lhLGiaPVmXZHmkdEec74eVVJrdvXJBgrMf4CSvuAZlpaOtRoj82zMIzW/Q2qWQ
IAc7tv7Ib7Ir8LFDPDC1+0VmawpE4La/Bp4XqtDyg9QkD7l/GZVdR9NFckqjEIXN
TbWj32YEHxTzHK2ZDdrZu1SFQiEvzQqMjyqWT505OIOnD/Dqf5Pg5v4SAGUfdax4
UIZfMME/9JxVBicTj3lZe9N6bL0EEHDAwhrmxPhAi9m4Gkxj47P1b0PO1BsnMoMC
pRG4jgDM8PML9vM9hse6rHTyhpm8xl0MsnhCKF4PQLhUdAgKtXT0XBPgOlMc25/v
OfObmSRXUmefu5qGL3/YWau1eLUd/7W7NFg7GV32i2RwL/LXx4fAMq/ROy4wxPd2
P1nKG1JgIIlx2HZKz9ElnfrEfsdPcWmnG9unpqYOQlNgla3rT0kovFaJYUCWLAJK
th2QQWyFUazaDctlwHYCAQVgMU745GYAq0JWVRSBsqI+aUXPGTacyM6Kt5LJuGQ5
jzIVFou2EiGyQGpc7xedSAg0iATqT1aC1PQ7fXx5kx/5nlJ+TFlAPgEIcznS8Mg8
heYVKpVm5T9p0oUNvdZCnPiDYRnf30nrxaqFcej/0K7EweXKzE3peCNTQiV4It+F
y9RxIHZGDg5Nm+y/D8XNuKwHg1qMCh6H7UZZ+LoJEquqjaoHcBH4YMnvEVKsQxPT
F3Qr3cOi5O7JWXrTxCuB5oxMfViCp4CMSXrurizsjRUl+/iA9/nX0oUND2NF1vr8
GZ7l1H8xViPEPFrZ+dtvnh5+ZlZIhyQhl2Z5AFzwuT+/7mRunZmS0PUIHZxmCsBj
4vPX1QPBSBgbpPRpBb/Dlg9zuXyXK8W+U8ga6IfGfE6f3o6Xtssix1uKTnyd3Gep
Z0kJA1jaQFRxGH18gMb8PxmB3qYZ0a6ZC0VzmBmeZVeSbMwZqpxFg1Ymvm6CL5IU
4OJKcdTAkaG+3WPT8q9QZjLcGOPk05N0/CTncJ/Ze4dClp6/9trxUzW3/anSSQdC
1VFD+BGmgJ7AR4IU1J9VDQlut7ZwCj33SYcZub1qvvMqvD/2ANRdRWqb2ntcnBxU
aNnYOzeO0ZBXaJehDlaaLIiCZRj+fpJ+80OAf0Of10vgI0Chb6Recy+lrWL0gm/n
4pUgq9D1e637EZPYTnN7izXL06xRlwaweQAYc1UkKqhORzjQjBYIfz9czKEI+WRx
DzQKsHaa4wffO17Tp34DEiGO8tbnD61K9pSh9kDsz50p0TEi6iiWsAAAVKbCTNrd
VXqmGs/bTOmw+Vw9rXPBXJDmUWe5oM/a6ggsysNGkNAFR+tTL/T00h+ZehJ3dDux
tWWjumDBquu3mcq5JPQr1ouOzA1Z1siTpY9LIvGBUrmvXMhrh4bi2/p90DX/DvXe
h3wRCgbxl/pHejE4MxcOZzVLu0Znbrb7sdcR9hVPMIGzEVEmnQJKSUOJPYOZfKim
fA/PYKRo7OmWEzqpIzjZRrydt9eOh6Plc0b+qoBABTdn49GrDR7JJ5zhlVYizNdt
ElP6eoITZaM+MQ9i+HvqpFXx/s0BMwPFrz6a8oTObxpsSleiw8xYd5X16ggKRU57
FkJa7jnOqIOe51OJVfb82tuCuukq5k4gmdT9cK2f+YpU9AD6x3DHkYjKVneCuGmd
lFuSo/vWvaRmlE739fPJvxURbYjmcRqv6lp04q8VQiYdgOCXHSRUkFmgdspU8C94
HXPxQRYRGt3+YvoxEOBDbr15xM0Bs/kgw3Y/4clyqjamU1K4bNFP5VHQ4QuQYcGL
OwdmwPRMfmDU3AvD6KaYz9rOyH/HRonXAbHCqvYkeLeHPXhUzmbx6WqRTiqsG+z7
XWL8TN1IJQ4gcPf6ttRMnP6EBaRXnbdWW7HsRuUmVveIInktSr4zf9+pdL/trBvO
nxp/4CMy6XyL0Lfapluyrl37Izk/w4fWh5Hry8ncG8vSycOm9fNJXTHaGCOuOx2Z
ZWNZqE8dfLKy239avXwOFWX6GTYdam32LhNlCl9mzY92s484tZb+qKqbiTvM2VlN
xU8guUVd8EISapbKu5ZeeTbcz7HBzIRtGfTdkmEWJOBJuTX/co1wO4Wcnz7m4YyO
aIGNiweM/f2htPznx/qfJJKDHwmsh8a7DyDSCKuJOvwv/2olW3PKF/fYtzF+OHkj
k8YOfJRBNFWl6I+J3jL7wJhOHJUeW9fy4e/pvUCNTA6dYRwO2WY2S1FbrkrlG4g9
kEWAaqSH7b32P5xulGHi9pj5U1YglMfVOBBg5u3qYzuTmVVog9AUVFFHmtIdQHiM
UV78EQwoJFi1vqyoDTm9uLmd9PLvjA+R5LRwLyvY3rTl14CHUMdXRuY5otLkiyy9
UYMBUismC5umrAlLULr8sDG46EujLPEegLIuhEmwaWN804BvDguJXZzOO+077HQ9
Kr9QZmq2csDGuZxjiD6YMi2kTeTqIuWCo2KRxH64gf0cDJwGImBP2x8DoFXe79ho
dI0xD+j892ikN+BVppIAVYlxgIooYMoKnzRLBIRyyj4loQhatJ3I/lR1KAnB5QzH
76VoXyK89H2FFAQ/M8fpqzObXcY3gH0bRNVnMScYe6CLK6+th2v0vlRI6xZnzrMH
rY53IT9Kh/h2gkitE+IAiURgUfxZO0j/EDR/VKNB9dQHl259eqRxf/c6rZ2yEbyk
nRxX2AnMTO4hVbHKjAk76mSdwmxtlT0KBo85J3Duf6BFJI+AzZLhFeusBMDXF/e+
xzHIxvbrx/CMUiSuoB4vZ2E1AYEYURf/JFzK7EgXaUYTBg1PzcqwqIdyyH4fso2r
P2WsBuqAyL5wdtEsLc55rvcaa02m+BJ8Y+A0ia4DTmuO4OxgFdOtbHKp8oO7vKkW
t2ZL1UOf7mmKzo+b5nircuY2f4kCa/6KcXvbOnYOjXMHrLbdyc4+jyswsaj0ITFg
AMXa5EYXA9ReIlzVmU0hz8Fggw0PMRujSNbxXX+HhORX2qfRMdxJjYgHtUhHK0Mw
up9B28vSxgA5DjEpIInHye/vF8JwpYXqpyHiij/XbbVxb6AEKLsHydINxpAtMffG
EVtnn1J49YjUtsdKiAK8IOwXgbjWJtZ3ASLT7fplA1eEJemdzj6Lyz02yww3m2gd
IdzuaPAZWOceMu6KhRk5sH19VcijWbbn4elv8gLHUu8bvFJf6p3gVYnBG85OcXcP
Vo48554fxFXux4txgM0+OGJRiyv8b6luItZ78QQ8T18KU9kgA/zD6lpIqwGf+uwJ
2pk+AjVlPdjIDRKg+10Hfxx3BpmhmPb3UGXKzzv3CMkMPYZYjKH7b/JggDjCoRc8
zf3kkE1zk8hVU6oPtgVe/72Blo4mMS8Ub1IBqfrIGEbEe31BwetTQG11OxArYJ8v
5/LU+nJlFBs6UmvZ5IO+hkAhex1U0DkLsx+35zZS793k3pBQs9mN6gO04Y2VS/z0
2qs77Ec5c0rbjfJfHT1kr+hXv9yUQNs8HajKh1pZZQyUt1Lf3c2rhk3WqLZ5EsE6
kVBi634y3pYdwhKjWjegVoV5gM7v42arRBJr+Chyz/f5Qqsmt6qcH7HB2D7k/kbh
EWZVJS/DIZVQvSIY2KDl9pqs3o2SmCA3w4PXOKoQULsbvcJpLKD7fAXEQGW6d78f
aqQ4HFxusEgqRU/lJ6mdsPjn+dlqidm7fZoTp6ViRou7fSkUQjatty/dgjEQzL/l
x74yLAs8EYwGsgsxa0mV8rKLkIRzqw5DmzLEXPheKpaKW3vPESPJNvchtqQY23TC
T0MR7A1axtx/0JcytECg2MhgoABFZi65s+WiAtzu9tya2xfZc3L5PYop5yDY4Keg
`protect END_PROTECTED
