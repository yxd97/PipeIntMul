`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pWFy570LX4frGvdgEZdJE1jC1+CqT2A9PxSbxenItMN4TPjz5GxxBN3MVdVsrQZ
VXvcezUSVDm7+2j0D/4CbPdXeKz+wGqFLebaoKzZwN1RaozouoX25dZ9Y1tjq5Ax
SxGxM5TKgG4/guTKA/dnsWyiimtGkaLqrf8v4Mic3jAvCYc4nsIcHsFyDNoOmV0c
rfkw2xJpe4KkooU5HlD4LhFjPnxtAl8EyKN1R7PspVL16UOmCRwzPQQBfbvttNej
d7ooK+suY2H2TPjEUKOOw/YLldMfQwYrpOLNFBNiaB3DCfl/3tjqe4sKAc5ywDqZ
ktDR1SThN8G9H4d4RGwUyXPzDqZME6403Dyvdsx9ga/HcoWjivQlvkLj5GiEJHyx
Wus1RUzOUVG4WjhaLtYMCzJAlHM2V28AAXb4jODir3EMgCZdF4D7i9JqetMZ2Z4j
w2bPqwVa8rx8mFOTmd0tKLjlqTPUp94X+oi8v/1Lb0fD3o/sYKS8hi5OFutwIM5d
Jc3MN1inBKkwX2ZU4WxlHvmIiaubU5TaDI06FkM9NvObAx/4QFWXZghuGfrZfm1/
R+3mSXgkNHN68GOgWA2r2SGRumDbo0b+efqy63mjEA8=
`protect END_PROTECTED
