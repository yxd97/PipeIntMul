`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrKiMWIc12kCHBShq0jSPM2uzEuIV2k17rcTXxMdTuBff2ieh85+7IE8tyk1/cpU
XUnAh9eJixpLGJhIzqS5GIm5NlYLrYexjeYtZJqjnVyX0o5/WcS1NbikJu+juGP1
JIp2kmuAkx6F4SFVVPtHiwRdg6xFORYo1MdHM6efE5IwNciTau0Xy5Q2Tiunq5ch
zd2IEblhLI4BSWgZ21StBBx/1OZ3YGKidw0EU4KrdpgR3rxcyQ/1SbCz7PV3shR8
TbNoMengWt/+DRSYAifCx+GG/c+rFfjEDO+dYAzuyBj7c4CcjV0pdZIt9v+2Ief0
2blkD1Ai011ofuoFrJPlaFY9gui9QB9ugCE1excDRPSgIQLCbpZoHJOP90mYERQv
JqnC1rx6NLjzmpWUDV3GUJgPixZOlHGotFyuj6UQi8gVUuWumXBr13zLc0JJSETW
zW0Dw2r0wZ3wwnJa/nQLi8cUQ7rM4P1U9ptTl6yetaSQrX/5lTJL18eRx484isnA
loc3KtgQTFSshTMPRuXgaMrKMCOCMKNWytv9JTgovnXzs83+gAmXdDhieCJcHuAX
3gztEOKU3+44SG1Jy0SNI3vKbt8wR8hb1+PaDWqpVaEjFgSr8Ja8XG5RzJjelwQi
fhCj/w5n/FUu/5S3Wu1eR1Yr9i8WLM+/JInLpGNX89vNR3pgXe21AzQ2R6v/Mlkw
43IK8vm4QaIPU6exGIqSPSjd2FOL+B+oMspx9OUXbg64QblE9YMBlp9ZslvwhCtr
fF8JShUdptnCTFs8fEAOSDFmxO/rXbTGPrn441l2ef77KAL7q8/IqqabvYfCGgKv
ilTILEAYK/r7e78CfbITniemi7gyYoxvrrgQ0OawMFH2/UKqUbKBpy4bvN4k7tRs
cuhYDN1MMmqHVRmhszQa2orB2Z0hxI7HvvqSZlhOjPrRagLNKGaTuTXqeHLeq0nh
7909gSNYqDSXJoU8R8jj4N9TDvfIZygkFQtttEUj4QB9lHN7q0oUDY/SjuqjTSz+
YGCASsjEj3QRs7hovstItQuZvV8pDMD1gSOmsuf237mcaTKN6/LN2Y7wtnunqcuL
u2+9GLOAZHD2QhUA9VRDa7KzaD+8Utu8S7ebGwlCKbr8GMzPYiknQ/Z4QWHjRcKE
TEjoy1Opmai1E0WrS8tsATIYjDXUZ5x9fcFaF5lZ0+XXcTfZaW6WPyBxxoIAre9Z
aKfuUgO2nZdjUjEdSVA+hThT93a0RcHGmapm1iv1UQYgD/lASmRxrSnA9D6HFcCr
U3lv8devRO2IooD9CPA4PpU4xQzKxQBKld03HV0K0PGRLbebsrGP6ezH3adNu2a2
4w3DK/bjjSxBZ2AUqtxasIJZq51cSlBpeFp35hqm95L65jk8BEiAzB3g+Sm3bIFd
iucZqFV16NdtiY6jwGy7k5byw7143+6VbJm1jfpROos5oQOjhHSgQfDkzX4+D9zC
aRQpl4YsWuQM/DIwqnQn/d5M6B4ol5S5Wr6sncCJRZqyQAFIitZiktWvv9QFntRR
HCqGZ5bGnigqEMxpqcUZ4LVHLegKd33/aVBmNa+/Losq6z+PLSFnFGzaPMvBpoLI
lk7oRBysknZFsVx/75T8KvD7NWk/SjSvHeVTB2JFc0myAQQ7dmwTL7kotaVAftm5
fG56kENM93znwbS3ACGo+WQy8vts0uIIlkME/DOLUgvpnHXfMRCPa2VzP7Akzik0
w4QVvfc3zgHUg5/LAGRGY+g4U843ocN8G1Ci1D9gh8/NupsdOV1ePCx3bRWpN96g
dbdZntGDq1WngYVjVdpCve0a60MV1SpE25Dlv+Szg7EuFTTdtOk2zaynf6vGmmHB
AVcpOjQVpMVa89uUnFEY54HxZtft4JA4gquDWQXoESUDWX9sgoxOHL+YnA4CEEjF
KI3uH8RX0YotY8MLv1XuV8ddquZAMTC1swFMMJ6asVOjnM4xl6JhvjCi2a0KUm1Z
/+Yrrq9RdFCOeoYoycnbQHoNMSLOYyn1Y1TuEZP+AXAKKfguWzx7XcDoYZVP4a49
7/Gzy0M0oMOn6CY7hAkKsKYetRxg8qG+IocK2vHTLXey5p+g3kSt6WjdOLuhCX8H
0QAbICO/Fp3Z8f2Q2iJbZ2tsLjPKNlkMEwNYXzCBNUfBjAEeczXuYgibPLpIHrKW
LQmNeS3vaKbmAqkxn83JhEvZF2rTzW/s27uchMhyx/tWiBVDMwUrMrArbzlwxEaZ
mJ9d/U985SMRwPH0zl/Hp339FBfe+EWm7OAKTYYyZIBiKHGiSnITJsKR3JbDUNUm
LKwDMpLiJXMUGuoCsAobgnc/nIvt3ZkxZBwZ3eARqNTs7cekTsrqRmIv3S8At4wU
QUVoCYyBT85iImZHbpS/JMSRmrY5LiE00VwkbnZ9uvUR8o6aS6X44wToO4SFaq8D
HVEzMxdIylyi5rachzcP8lE1QIFaIvrqEOVwxUAX2kIEZW7FmDFz91TURy/Hv4Uk
1g/yzR4FvVOmpa/W0H+7uYiuv2C4R0azc/qeYzVUMJevDdFfO14LPyUzKy557LBR
NeS/a1GeeVKNMTY5FlOMBCBA1a9hgv6rcAUDf3smD/D4dJGyion+WYhv3Txv56d4
p0WdIqx+ClVg6SKU7CyltTtytwDWw9fxb0GUbUhvdj8PrMIsN5YLzwvDGjXjhvgR
juMXsiSB7e5pO3MeTj0/mbqUv1a/lYFcNEbdM6DvyuJGSsHudnUV80euKZIeXjmI
3RvwJcuqBtncoBmWwQ+aRFFaYrWAXKt7kGg5YSnQyWJ5q1PwstHpVH/xa2VxKvkv
j3EWoc8CBQv2mok13xmFUui90tMX3JE8efAmc7HnyMrAWLmyQEyO/wIbNvk1TGID
IQ77JBSj3dQrhjY0Tv4h3V4qKKYul2H1bq188OXq3Pe1M99rl95m/R9gvdqJ0/Mw
f9mfo4uMa2NyedUAsj6cqsPPkOM+8rxxw93WdcOj2jXY91+f0MPmD+D2y8/Kh9KD
NkwBYxX1xnawWK5HRBVIuByiEv7YAZltvaSpI6oqXKW/octOy4cche2N5DtUXUHZ
Op30nSExpqirZwA0RPBTsmNp+zEVMohMHA/Dk9fQb2Ovj09CuHBEH3W0axx8Lgh9
7POKJz+CfMJsYGuEwMYLrBjF0XnYnOsXn/aHKGA2m9poJCuERQ0wbZ1lSW1zo3fk
P3E8uMkbHMlqkXBk23rYt7gNDgh6chdula+yDba3OcWl5DrCmWtai0mRassixnFL
SGB7B9DskxG1ipnBj5O9578+uA7p43kNCI6NK88Xo/tiTZcY9Mj2VtFmRFKrR0Aq
EJJmei773wNeNybtFBK33UTyn3raNJbiSJFh9OUjfnxB67xsENT382NOJKLLOT0b
BhF/qGUPM5U4yqpwN88rSAXjwJzwKcpqBrqWmZzrTq3ORGRTy7ukOT8xHYs8KH2f
cBoT9R5I0nn91n2qBu3zJoDbvEr8XGi6Bb8jb5o2NFCtfFD/u35JX93Ht0HqpXz+
kivLfOfgXdwOI8wW5JCdeGnX+9laMSOGBE1qTyRblKoZY2dTaVtgvUhuIHHrL6M7
SCHhtIwZzKMA2hNdnC0ZCX3AHj7UIhecn3GFKF8JVcdiNrsuWz/AwMfg7iKmMWNx
K/48mgjtDJiTJS40RkDpWLZalqFkn3RAAhkEKybNWjNy+tdZR5CYYV18uUW8pyrm
T68fdITOMZx6L3UrdEszK0XLmKODQvIQcP88qVFTtQNpBGZAKYG4jEEplJC+9Q/B
xdxIdq5rgeCIx/f9qHFPoB3zHqh6LtfLJ4iHw6WprGVnt5bXSWwt5JrpbcVZK+gJ
s/xDyW8D2+9ZfbwfHAlvHBc3VXWh1DiUlbPycTo7eQfBijHWa2Q81n0a5FjFTqy5
lnxBm8yPtdath2mIXWI135ym19AX5nV7lIlLx938Tz9ZtbC52Q/kobrHhBENur6l
bf3KRcDwRVWEOUGRgOS+OEyPiqwskqdJVMusnabn7782X3l1+oakR4twLW1N7RvF
k8QRivRGLJDJ7SEkoO8sP7Z8sA499+Hyj6vajm/Z/NvOMkdcoPvTmGnIcgGqpL7o
xcRWsYL7QVhERvto9DjsaznThcU+6NMcKkVfDQFYmgh0GT04nH2+4t4OluQIHgeu
sqJ8jAusZja+8Vh84KO7gKyrq3otkltRzUDjmqCqEWcqfxTZXBoj0X2VjdQBKQES
cFzDE6yYUpX+iFLLEbBsQp2o5mgoC6u5cRO/w8jZ5FrZ3aZ6xKl3TTGQDg6kdWqy
vrBK7MxS3SnHZU1aVVe9p1iaX992+GG5/LKKrEt/hXVlY2+mS/lZEXe0AHDGPvWt
UnI3nJMR0PTMsGNF6LBlkyZI27LHuftEw3bwegb5iKFbODwjkBXMr1H/q7Kvkjv8
6/0RwduWpXv/yMW06DPmd+kkguVmvhWw9ix9Q6uL9wvj4O1+QKFVW0bkNHurLu2K
0PHOWk+hJ+59O9auwaacEqMKRaHR4TICzwd8miylfBsa/QF9Jk5N1BH8NaWINoZS
TChy45yYZCGxMcWDx8ONBjtv79DpPt5LMhv94/AOMitqbhlzZcsflySwV1WF4Rd6
idGEucsyMV0z0Q4TmEurwLpz8/R/RCjuIrC6boOzla4vT966TREgzd1kvTFkUnbz
DTqKL0TvjDurVyE2WVI0TeC/01/KbNUpNCZhPk7yE+RMAjC48YynKhDATn85+G3a
EhcezcQZmN2DOI5ADqweuH9IWYX/yThcCgnQa4q8c02+h9h6LZ0s72ddlKsI7SXI
1pJyO3em6W514EJtzLMRo+MAYqZmKYvbwm1uhUCqmY9Ajq7cch+6wNfl7zvkPtAN
ePnf/rCrCLlxgi4aLxqkgv2wo31wVlorEgorRTsgeUsqOIfzfvdtP46rw+IgoABi
CrblIEtb0DdFBiM6PtgYde0o/SIXYUwxs0/pxuO0ioUuKS7h2U3LMO50GvsxoBlu
WqBcLJngPHKUTedaOgh3HhdwcauW0k6whxmfAKL5UWmeavhHwRf2wi6ocY74AEGf
UJEVQVOokijWC/V7PJKBpE5YsejIRXwIApJCiXJWDDHiq4MZK84+oGFGYmDOxhlK
IUueL393qatd7Pi9a39/4VDIN5mjHGoGtd5Xlq622QKx5BAUXOVrSHWuY6KgpSIG
Gka7D6mUaI7a0DObN8ug0e8JYehtd6TLFYKjEgtREHMTE1Wox4P3Q0k+of/xlbkz
KHUfwMh4kVU3vvl215X6J9OT76FVWfgEbRsf8KlNLT4yFSS4cX3fb0PacPhJ2RNO
2ML/xbhWygHC4w3BGOlrX2D+9+Yoc1Tf1341eKhvwdCX3e+qsQFzxxxdFw1N+YcG
ahSDOX3bDLQBAEYW4tel8eWakgha4EQl1vc87UmP60gJA2SWNe/mWsZLSd7SkSrX
dh2Bu1lBt6/B/RLbc0W6rOkjIpIVZ+0yJQXyu74PPU5p2VV/5nPzGdiEK2MPitHC
oyQYk1Ca48e8zEJbWyfTD3C3RshqxdWNOv39FMzK8UavzczKC6QR4cGZ7tIaCAD4
etwlDFlQY8rgdEMjyreqO8gGdvsEktfXtpHEDv6lfCfk4JKQrBg/Dh+XdI2VOxli
ITcV9F8XQZBbtipkij7mbQjZSl8uJTZ1Lb0aQ6unBVI=
`protect END_PROTECTED
