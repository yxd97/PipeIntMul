`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C99+0Y+o7c1lXfoXMGoNuPNp61sZdUnouQ5a/ilZZw6nRFLU5ARcSWqNTpYk1FrI
iG0CmZ7fcrFuAVfP4lSu/v1tHn/Z7N7TzM8+PJXVo//FHFdvEzQzbamb9tFAjYCs
P/5Z37j3LUI2LYtTp5SOODsmtzVAmrcpTM5w1dT2k0s68K/hkMWbPzYCKYK929Tc
qgDjLTqneRdZL0JR8czPEJIFiUh8BuCNLW9jcKa6pW8m9BvAr/mjuXQmRCWVLjMe
EOgRMHGnEdex6zdveA7phpBJLYGmSUwG0c4DBf2CFA50MaAlzBtV/viU9JUiG6Fb
l5ljsUihm3PMJh5fdfIV3IcYbVBfJKcxBWDxywvJmKrSGkQd3toYuKIkinawIWqp
3kqA5tBDZKEBd6dMu2IdznFM0s1OtsTDme29HEmSrqghkiu6yJiZjfFj+5/9GfSq
fb3CzGPLGsJnh54YNMEVjT7ntTiTF2vg2R+wW5yYJJgyafp2epvizLwbga5eg3QG
xpshb3mSCjnG8r3lgm/YhyxZQU+2YTEpEToBSYKVnlATckPPpd/nzoxbt8JrKk4v
kUKgABoetfskm/I6RGbFvW0QpMsUE3AM2uKzX76SbWEIZpmdKy9lH4K4jBHaFzep
fQRedX5FrU+obEffbRuca+IUhY7c8kR/+qWppga1nExsJkgrPEUUKD7gMgF9OH21
GrTrJGy+dW13NnfN/wJ0DkuX7TY9Ij0/CxepMrvnnIhGg8RiNcyv2Ng4GIfD2bik
GiYujMc7VzgyvBRpKsn3B1sJXURmiiLQCJ2CMB25oB0XwII2XbF8rju7EzGzYKeh
0XtDhmXx2OhGrli9kej31SbehUP4eIktyvtY7BT2Skj61GoGOudHhIR3zUJn6CMD
6Zu9Tn/WHpkWmrd9rZwZ7iVEnz3kMfefGoF424b+vK0F4I8ByIBQvc0rFekcerOe
ymHIgI28HfmgCkDUy9jjvI5MoI31FNYam2MBnBoF6goVhIdRnlH4uZ2w4aq8TchS
SKBUg1OfToSa9vQp0qLjhV1f8OSPwEAx8p+mSL14wrMFzgZ63+6nKZWJcxl6bHZs
xofRm320/Ufm3fEBn+oC5fyNe4kDB8heOdsdsQ2A+WRhleKyNzQpohC1ub/PV8qh
SQctgOrxk0Qoavje8p/k4ZfeavfoHk4bUYIC7GY56ClSGJIKlRg/8T001Ay/pVOa
SpmdUEZrbZIBSU0M/4Dqr857U4JHfuXFq7B1EAueOpCjZXNZ3OI1ADRZrScaAovW
GnHTuo/tROu2EcQe3sbDLfvsq2HJ1tIllzOKFm9WmNYachbbEu898DH6wSvwl0ds
JOfXKvC8hIitstOSUE2Mkoi0VnhJxO/iIyyluoIx7bhIZSYLXv/9wB6/fsVDMLyc
Dc+p2yH5c5PXTeVhhb59hoGzxUoGJ3yo+TsQUr+37KTEc+/zNumanVDD8FxX9nTb
GEuoCmCxnyD/4uP55ps7GOtBUcgC6BAKFsm7fbe8lSi/KwT421+z8xYwElSKXSIM
t845ukUd96YyFkD/C/zwNm0v+VMvuDFSw/OP7Mgh4RRS//VvzS17oiuewgqH2oIE
c2ihJL5pvBv4cEGUpHaEAZTLws5hC9OSVq2PFnMCt6CONNXyrWK6dvDbAFT5YQUb
iXHX+H7tjUmwBk320MPtt2OzBw67ImLJVcOGUV90uq6vdah5N61dlK5JHlFv8DEE
U3gF22nOWRpq47su2ErdGk1p2SJI+K7EcOXnpEtyjbpTLS7ALX92g3ApyHETgCEe
79fvRAXjs6ntSacFn1+kTZ4UemOpDj5KzW7pJRgqjOV7l0bOE6eKSRW8NBB1YDsz
skc5w7IraBsG3rTftfA+v+vwztsrwBOLy3stLB/0NbzYyjoR34ZILl5YaTNhmOZR
N9UKS4ZiFlpKfcNSEVOoPQCr3ddaGSgpF7u48G8dQsw1YAkMk2P7Ktiw6JtM/GXG
bkIKu6QYHgewjYkojjvjmri+6WBY3wtMvnw99W0lKnJ//dK2uLyZtmVLfcK8wzw7
w6gf09XBWPtDAcTu0zUDoFjZCCEmkDQjAe8Lx/ZosZuit/DdTyCo/18uqOBk6eYq
v2lFITuoWP6v0nY14yw/xyvGzB23my3gUmzOKuVC1RoKq5QWA4jArKJiQB27s21L
aKVIo9wsbCRD1je9uLd4fR1kcZBE7/6TxhOOVZUumopJ1ndKkgw7AtC3WPLYkDXI
5pNxZpur3I8F/3HQ0V5rHH65XK2zunrINs9YmSjko7aDe1O1LQCfwN1jhU8UDSvg
vbekjuqNS1nPBz8OlEmJIXmn/5kljlxSpMEml5LyI845kLRSEjesnrJiHTebbI3l
VcgE+k9rvDNe+CH7puaHWONYPbDVldfMymGs7LFX9JMrYghIwzP4ApSm6Ec61d6G
cLPubSqroM8efWDcYx2OMxcTIEaZ3G23yQlbXvqMsX+92FPxzYT1CwqltgQ4061E
qNTfP7YNNfv/7pL7JaVP4gmJrgRpHE59cp7PAthXdWCB9g9Wa0zBTo9dGQlc3kTc
X9DXr+rKxKjCj3B3S49BBjvepU6mpobG56oBDBgrF5XyMZ5LSrwljj2FREBwuywA
Gw0Iukso2//z1aIuG62116FK978MCa8vMN1/PFeJYdzJeeG0TCi3EFgDAT0v7rzB
GhN9cYdvham4V2bkQCEpg3gzpOhRnIWKbCvFV5y2NbY8MX3rROgHZ0qfzB8NCYoB
JgAEsU+1pt/sMoxEM9R//ultoIxLIKqxYiUrB80L5VZ2K/cOzGMjJI1yHgoYoLWq
kiiVQ2uEzxW8AgUQqWVUI6xYgyUm5zkSjMXatQ0sPDpCHURxGXxo9PzHuBT8axEq
M4a1HidzTIrbmDLua+hCRQRA7NKys9S4H7s0piGT1gixIcUFqG7C65ljzTQRbsia
eJCHrYA5hpAdVRiPXWBCcrcdwKhnmGABVnh1tQJUoZkgXNxPGXIw6jRzvqw60fA6
ss4BLVtRXXchoCkJtPvcqJtsAhEs2dUOsQ1Jf3NEc4enCTJr98lAbZQMiGuNj4uD
`protect END_PROTECTED
