`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6dABKNdZsHsbgPgUD5JuR3oQ5HLPT4wPOFM4+n1zCc3ZeI103ypYsOhQAppNfkz
jXb71P9t36kIc+dRKO2P51FYEdwHtkhlP6lR6DhK9aHoH/yjNDS3xMnrJXOt9Kkz
BjjhhgqlnGARWeWh261H8D3APva708AuDBHKOEn+ptdLe7G03Ve5r2dXsVefXCCa
0eWc+IaZknDI37ylzGWu0BhfWWLjp0xD8SBuXDdQQjcOjhL66iUHnMUC0Q5xt1/Q
wmOSB9sSohWwqG2MZNzG8njlD6aF3ow0Jl20mjOU6fo3PP6F4C61/4thMPhK9hL/
dtqtUbilPebWnbosq/EY1ZOtQFSkOkrqPFiuJiS/9hZpfkt7iHL0cqYKPDi6xb2a
3XsAtuVsLAA6RbUdxjhZYLS3cNKtOOvAbPD0YpKHpdvCHq6vR5hMTJoDT76omvUo
4exleCi46MOSjMeUjxAOcGBfVsbRywTj17HAnnXz8/ohcT2DHyy6dXGjmufCckc0
h4Mb7kAko3AZhuRsoPmjRh3MoGhKhqWWdjVeBGsUyBD2kEEds7YgW1Z+22yEtgmV
x3+KNAql8K9NxEtm+Qunf0PlRBhMf5gIjHHb1usTnAhpXshFN2325t7cQ/1RmiIV
/kVFVyMLXzXN8HxeqKqQNopCbLodivLyUbVqYnkIWpQ1igvp8EZdHFuAcxLouGhR
rX/3yxrN8VQ5p6egYFhTCP9SXcouBQnGYw5KQTQmwdyr8GVF1Yn8/fTck9wh9bIH
x4JxyTPamG78dUc/nrc9gEQQNelLuT4oX+FjH8BjZlgPQSeXdHDNwl6mqMqRcHWG
LnFqToFvauaNq/cSsrCWdgLY7CiYUT3SJfKHbyVws7lqkFfr4FJYX0l1lXZ6ACrH
armmB9m+eVMO4VvucbOafrH8pZd1q9wtQAqk9kSDT19hMG95TtWPBxHFjDvGAaVG
6W2gLcdfRToUfdMIetEdMBDTir8HXnSF0gn7foOxePzgYcW4Ti+0PHcQExibFfoh
gBR2j3j4ZRGB9my4qIJiHNHMa5EeOcoKPvRfhNGT34CQSDaqMyOaOZ1dsdOUKd5b
muEKeZ5H5Qp01K7TMUTC0YgIqrek0vO9m0SvR0FOBPGSXkxGjx0vwiopI9hau7y+
Rz/+HylURCNIOaqOv+lG64sltvbnMfkFq/gs3RWiDwlcVXp6w3n5o/zR+/OW8Ugp
LZiCPfUw0uEQ3pKdL9Fls5PKPfv82G/PJG+KFUXE4+YVe386N8Q2lQdkkA3+J4Sq
`protect END_PROTECTED
