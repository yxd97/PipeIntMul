`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdoDokaZapY7BizBkNxd8auRA2WUigkz3bM+MtXwKPFBWF5wEZCYU0GqAGmPHccc
IEZE06Z6ZBBrUWvxq6ilI/VptaNP3lqGClYrt5bdZtTsj5/zkxPjiNmmVJCorKDl
6vrSDZWhTbt8AGBK8IM30TUAk9omdbZ3EtPIwAxiOED1RrSe2z3/4LD30zsPRbAj
+j0lJx+gIIlRJNEWpwogx1n+PGOTVWUyns2z5qIHArQuSeIWgOdG/3+Lx+n+2qOb
7IRP5siL38N9Xf7pYdXWsqUxWYHwy66Z/Ij3Y7FoM1+aovNTzMX4RnYFjn2jLVGf
coMmOJYWg7y6ygTkQw3D+n1g6pz8KVy2JehrCqBQF9/A3kykUnqAjw1WWQ8EedJt
CYWZzdncspfUFXDeZ7CPsg==
`protect END_PROTECTED
