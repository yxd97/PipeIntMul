`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZodAUXF0GONfmz+gtOb8eRFoW1d/xP0CY8lsMu4uLrNNRwXnfpYWSY+Xnc7oi4NN
zfIeGcZGDblQAcOLdilYFYKF0eirfmBvoP5PuSqrsL/f+9Rfl6kEng6A7KJlZxa1
PwtiHmSMaaleiBArut/7DRvKGIw/7a9zr796lCyIAEJAQjHo+RCtgmgsZjGPuzs6
IStyo4UF+wf2SNE4e1nx9gcT3AO7HzVSBbN8Ey4lwC3zyiu76jWWSXTpynvy8E2t
po2FP8IgJ2V5ZIVG5W6fBBBlDwaGf3c/EjqtYjJ4bW/1g8Q0c3GOw1dRaJtL269A
bYWWsGnHuar071XkLDupxc1qhhtaJmz7nRdiRJkqM2ZyH86L6hTMgz8rBp1LzFSl
alVtZyN/FDK9J8Ys0sN5muVEvmFYSU3enXqXRXlREvXGsoJQxo5+f5dNkEKYbjCc
`protect END_PROTECTED
