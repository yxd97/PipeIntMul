`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fpApj5v+2KYLMiSpy/m2qPWA+3ISgMJYmJ0OXowjP5+zO39Sk5q0MEa4KLNJcuVc
KgLVVnWq50PIXAQ3+NjOrEBZAVoA6wHNJ9gAZSJw0XxkXqdlW/QmzaoKY/Bb5bJf
zQAG85vvdVsEcaSPK8do+InGLL9CXpfa3VrQS8B6gIsew9NHZ+vqBGXiqL7BJDpJ
acpIITJlJHtPQrrL9Sd9WvdiahStmLZXfI2LCggk7n21ZKvuGKRWb+DYfB9oW/Zs
9A40gfCG1bSH27Tk2zGWzv/GXWp+GQuNYWCUtRUSOybmky1xk3U76bIeKNnoPvN4
7J4OinwR5RviavfZrAZ81roU6R9SvOlan9SZzebiGqQc6PIC4ASFE1dawZOOGxZy
spDxeAp3U165bO+2p5iMeA==
`protect END_PROTECTED
