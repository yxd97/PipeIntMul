`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dTfEx1H3P/dnofqRc8UHVCQew4dTPd3TCSxDOGZeqVIiGJmL4MFfQEkC0Kd3O0U9
fAFrMcwNDSbEmssqYJLIAoYy+Xt65Nn2IH09kkFEQq0v6oVUNn4O4z6uNYhKVdL8
t5QY9sKdi4PyKDc948lK4EbqgIFN2sSeIJT0UBydnjlYODPuw0bqomDR8mAycQrQ
wWv9EDMLWuHzM+Unfe4/D8Fr5jWZgBtUY/y3mppa3Xqr2SA3RyRkmR1xmyVBPa89
k702F9OfBYrU8nafDWphrpWqcGaJgZt92S7HkEaD+1QqYhL2qZ0e/HVw9ObQPqCy
2iAqLbn42LGZJ2WIyCnKeWP/YhbD/XgTl+wrewfiw2QCxL707/4Z7lTk6IE+Lkam
ysb2kUEiA/0cXWBaPIwlC7zxVjqRT6mOBoOifRiQqH9N0YIu7rNCOx0ZJygd4bvj
Qfi0rA4QkNb7wtW4eGqzEN1KZILxmOT1XXks0q71bSE=
`protect END_PROTECTED
