`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+KKD/jm4UjNLqJcrAoFzHKq+vgEVLRqF/nfvLOQXVn4hwrNd4U7rTzAZs0DwqCD4
Q4yJ/7wu6sgGz66DUGj3mfXN9z1P0AN8XMHJ2hT8VSbp/lFo7ez3SfRIYD5cdzdn
Ksl18ytE0d03vS/FO/3/wTVE/kVEy926gJhn4TulUStbYxpXfsFO5hP5RHcVQdNH
RfMCPJzGUCK4dXdyLy6Fwdcx6dh91U9Dfum4EvHt9zFiXdYsNGgGNjXMLekwys+U
+sfyeHWnHmxNg8cHyJ8RdpmE0JK5DjYcuI/XDkCfji4d6eK3gVUonr3kXEh0MRsL
SUItmy7/0OS9+/yEg4Ij+sys1huSJLMrnQIcg7VTS+BndqcgwdAwlu66TYuaHpVT
sQqZNUVtoDeGt0T5ZSUeUylYhz1slu9l0uOcMxIO2x/VIyUkvTmIirXKdoMgIY4S
YUyWo2KM5CjzZUu+dDtbpI0y9D+C9Tncrn64Otuoh1Qmj4N8B96FwoVCWeGXUrws
sdSN2/gR8Mw2JCXKwrJ2rSQ8YRcX83qr6bJ3V+9edaRFOwZZ/dzjLrECdW1upPkT
VTl8uzS8CMCV289aY6byvs5eEFwpi0WsiDt4HRdFa8Te34SKkceVB4x0yk37SaBF
CFbWUeqqltSIPj414BfOhfU6cUrvlQNZio97jiW9psT3KFg45rVSXRE6p4ZIiRnW
lkejxngBGf7NOCdJFBMESBCaLPjL9Oz1ljmHNrhqFDs=
`protect END_PROTECTED
