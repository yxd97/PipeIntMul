`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IL1D5tpl48vMzBTkYZ4X+CK/ONWdKap1p8Si8D/193iD8ORv26J4MtUdnMb4OX6
dMxKPHtJ/exkUTkrCD/kw72R2iq2FdnGr2ElhD1LVnbSmWWu4krnAq6gGUqOU2oZ
37Im2wvLcx8CRCDNxl1xCX2sObZPeqi+LUN4AoDU9zrm982ICUgRsQCEWshs4mqQ
cyzjw3FEkWLNvk0IH18zrhN2TT0l01ajcuPxoneyAjC0h41F4LbfDlKhRvHd6wPB
yerXucfhO+u/IlnOgLm9erkCen96Nbr12UK+Z30aLHonpsF1o7F4HzxSB5zZjngr
cHwwe+DhWrg3q5wrRXD2XCj2dCUHkH7QLt3QnAlsDvxYIIOcdoY00EYVy8ETUab4
3ji+eXWDlGZrlnPT+QKja5+mR98JwnW9t0qm5d+N0sltwoZGYPVzkMAzc7XhrB8f
5RxUKXyHYbTa+fVcPknkmPW7dKEbZ/QEH0D623dfotMgrid2PP6/Aok82LqFRZXO
HB/7L0yc7Al2MhygFMxbWzFF/gm9xxJEi73nQtN2mVQVlFall0AYWbs8Xmauoesn
uBLeuiJXyhujzM6zrNajnRmxzRvIFUVWRDw/+ED16BQ=
`protect END_PROTECTED
