`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3weJhiG+f6uOAy49olCTtxKIadD21wk6Ki4Lnz27u7fT4zITjgtg4fkNyl+Z+AaO
/6DsxYeRXWWA62cAGppf6i50g8W/CWjHL2+Q7wwTK6nZQjCDbWQwTHymcm/Tl2Bd
PGxZXEnLmtnBuYEjpnYULAi+CRAZ5at9SKv38RyocsiJgwGsjcUO02VUvfnXvHdq
i1kUcUo2boAkE47s0Ugfbc113QM+2Fdqt/mYUoyhhDHMIWMGiLWbbt1j0RXu34eG
l26u/Bo/hvSG9uvVGwvjY1lR8tbUm57hVdeNzl5Qyq2IDRa8I07CBpsTcH3CvCFh
JfHC8b9a2VtBeTGnjw7QgbgwjIISFmIG2AksA5wiakqaFX6nDDTNELQrt66UC36n
rk4/4rpQONxjT3YFYuSuOA==
`protect END_PROTECTED
