`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eJYTAVxSM2LMLFc1PMgpcLbMdixKwmxpugvlv7apdywLk9VJC61eKxwXvvFDbLb9
xiSkS8UUGV+2vQcqgSD3v0xGcPXwZaae1lKTx/NIfWKOnoOj1qOhBwtccQzaOTtm
Ad3txUhEzxHWBPvd2R+ZXZqGcPrex72tRhSIYPodsrv0Uo/PhBwajJqC2CrNjJ7y
2E6dBckuXVs/dsBIX0glFZEjaDGOekC7YNK+YDkVLZ4gRVeBmen4ky2axpyebrVL
DDoU5Hxhi7DVutwILaG4nJ+5BjL65DdorUerq0jbIHvrt3BjX3heXqMDEHsM1YEK
gfHQbnoLiUvxeLr5aMPvoeRAGSNwITRW1FYa55mSGcDRVEq3DFzLRLEi9oUoRtJA
kWLY6FagdihqYLDgoqJKStiTnuuxIH45plIzzG8fDqz1NpXHV7Zm/g+C/UJ/flAe
uF4RAziU+ZlUTF2qM+WqiFaFShJSS7HIianGeg6Ud5UKkekpH+Gi3I0yu1zgohxZ
I8RkLqFVFA8Ec6GG+qdlH5+3AeIa91qocNcGp8tzWKAe75plllE1YuW92oYnjB+a
zXLGNpfKQUIRMfPicJe2w1SAcoxuSLPviamqXoJ0BVIivYmbYFXwS5Sdz56JuZvq
lGlyacOHXqThOeQrvUEvTFn29nXs5+pieNWgNDoBxcTeBKhJGlBFdurruDvTr/jC
VOEkqXQ1YZG+lO9Q8fF8mw==
`protect END_PROTECTED
