`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
93hqr0uGYOS4nagnk6m5wEIIegArLu3WXqwlTInc8aSwIa6s2xu240d6+/mxa4A8
g3tRfE+Yq3Gx2s9nd2EJpYTQRFSa7klFSCyYfL/53bMURX1VgIU16s8ze8YRLRq9
cL55EADfQ3gfbDCC4kcTYvI9Oay0PSrQ/Dxhq4+JS/YOVZaO6G9Qqam7Nzy+Zgr0
7LG+yrJDlsl/mLKmAAt3kX07PoO7zUY4EJPRba0XoKTKnmwwdo0+Y2xMaMFHBvry
IaguMYjgOXEW6CCTKMQhEe1X3gmqf1AENxGUEsMUOPk=
`protect END_PROTECTED
