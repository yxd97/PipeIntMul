`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dbDphjIXelJ1B1pVxcECjNaYkx+fwySfjLDrHoM08T1r/ibmyt6O13aDY2uh1xGu
PyO71exDiUScqQZsAZ0xEyof8fWirsS5OrvChgKN6NELQxtCy7MVzyM/zjrGK69R
1+YqHxo5r6CjEQFCk9E3Ck9i1CfK+6UduGXxUe7GcbtAjc/+NwGTkOGOZ4wXXaqX
2k/Wj95djJ8Ru6V4V5A19+AJtEhvkKkQy9En7nbm/2xmvF2TBYvOy/le4MZkQyIu
ViJ6A8nomuzbKlbg+hq5kBYNClLDMUYxvyAs8Kx9WBB0qB2YfjC6YDy2te+R64YB
YCNxV1w3pM6iylsJciAfKHlZfjyqy8BykSwIrFeTIw3DU89EZHt7CPeSLInSkpeL
+SP1LKbM8ccb+v/q4En8DQcYpKyjE9jSYqSQ5mJfUUZaqzOE4pK7VVd2mN7PAoIB
QbwOaVE5GFACpB46497aP+tAayJfU9UdPKdRxzNmvkeYed/kx+CeZ7XxX8LcFp0n
VgIDQ4WbnflDLsoYJA3r63puDOINDz5gX+ZaUED6Txg=
`protect END_PROTECTED
