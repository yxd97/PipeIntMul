`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OenceEv5war/PZHDA72UAIexlEiPZgt3QSPtcZXiW58MC8lORnAn5ve2klug2maQ
45wQqupJiNlB1nS+jS+5hLiN9xBRJRfAn3HTfIlCQnLTtBGraSarZTv1Gwf4LN/z
hJ7gWAZz18EsbDMnMI1QCZM71HDz3pF52NMPN1yzFKcHH/um0/c5UJ+lQ0Lnt/Hh
33ThvCTYzXXVazlVZ3H1zfwTQQnuT4zy/vv6hHxRM2hNwoOcj9RCrxOtzLGC/92b
NPLBwGMfGQWmcvbCzs390xxyIsnt/nRo7JNzuyHRnbLMhsDyuwRr6MdnUQxPMv4i
Cb/H4eH/tByReIooSw0w4hETFICkHPCE9GPUo9WvCFwNSllkM1D9lCgdBCL9NYbs
G90KvIHWeXD2qVhq9/Ycq/PfTMv793m9xGhdwl79oME/qNLnKusj1miaBIaKvmP0
g5wiJLoappJGK/XTrGpBbXeWC2FxSCd84KEtFgJIGBpU+Vd5+7uixQTWYJlQdEKO
L2RR5vIiokelA3n5cz0wZkDyDIe8k15Rqp3nPgETQWWyWh5+KHQuWtDKudfGo67q
0O4raKgmbKpRGzgX/gf5i9g+hRiSh7amVhVn5N17juIhpT1Bc2BMUe/3Z3/4l03r
q1b10IRFqAbsys/5N7wjUgUZOehArNGW6y7Y1JJG6syX1edI59Vntqq9bCNOetWY
arS7j/WpdBYs/X7pkBOkoCW70/IXvdN8tLYHDBWlfdGfj20jpG0OoTvFPnra8hAx
XBqlI1zMepqrBTr8hxayhyUP4lPsdlcypHTBH36Yp+8aOTHeuErf0a6hiIiNvi1c
wgjS/a41LNULwSZisFBK8LFekxTOQicy1NSCVXaeyOWx3+TrU8K1Iwr+jMDOKE8B
47nrXJNih+IA3CbVTCvz433myHsyDTd+pqSccFKxoG4o3YNNAHipcDfPjpn4u173
BvblxWCMHbmIpXQss1E4+2jHd7An/EGMfMuzo4sY/uCTy63HyjElIsVGE2LCbHYj
QzqiV6EdIArw8sMBCly0oT9L1LNR+Oy0QzKwiJDaoIikvDt8Zbg6h3wf2TT2DKkQ
hxbDK8lo34c8h6imOB1FPO5eqdY70kruIUFzXtFXSNB2eirbtkGElxF74U+0m4dl
UcRJabvfTstkkYlqZWSrRJpxHMA+hTmIHcJugcAmssAhcWC4cKmfC/Vrz/LdTvUw
X+IN3Mu2SQl6XF4kx/h0CssGZnY6/86jKbpqlsq2AHLKOVTboLJKMe5G/P+nVmMv
lAhxWXlCJB1NMxvan9Gks3djVdzMAJN2rwAeRiu0KFu/cn+qCSKJYGF/XnfqBBem
7hl69Yb47Sh5rRJ1dDdON87oF/YqLdBh2iH3r51mAnIYykjwq5aLq26+46AH7qGb
DbvNIDcszOJRojR4KvUR3kPqAbySTXTciI7HyN6m5GIRkk8ycGckLSaGHmuTfPxM
kVRo6wcJsyh0qSfAHhxXFBDLyekZG31Cddmr9plSjVRcVb7yNt6iJNCwwFRAyxUf
/BnCqwwZMtcuIRzZPeuA3G9fN2fAtblRSIlVzy9M9jckd8rJp98gZ8bfltqRTMgM
BYBRVnmpSDzrLrryqkriuI6CmfqvhQHVYHoCfj4ZRGfc5GmgV1UhUgRhZn6ff8yl
/29v1CYISAws1bhBUPAPs5MoJEBXqZeoS2+t6Wsditif71sdSh0JrUwZlGl38YqM
VJY7oEPZTXqb2CpMb3GmM1nYl5dgoZn6dW0r3vn0IbFRprxZb7qn68e0KmFsMDDA
lVHwghRbzHiIrrMABxAvn+Td+ojeQAtHyEDYvXgGISyQNDL0xbWzDzW3A/XnARDg
eD4erBdx2e0ZQ9Jt+U2Ivl86CQ2NwZVzYZq0LwqvwXID91Q1FBZtiGsci21w+Dwh
aLDtYcqMuVm90yQ04RXXmiQpDDc+i+KBZUAaJe27aXIbnwlKP9Xt25YB7VBKJZqK
GgvOpUTbKTs1NA8J0z0QjE2Dx9pBnJppuE4AxlQ62WYwzDKo25zT8bX5k1xWyMyo
hkOEJLBGE5n31HD9g6avBg==
`protect END_PROTECTED
