`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09Fj/wYhMF6mIi5e9zJYatt6WmMzLJplX4zBOdppFeU7OAob+Z14+uWDZSTZ+EqO
lerq+8i9BU3mFbdDO+A4gjwALtYNUGk7evCAbS75iXQEdl3bstnpsBddkixInIib
OSR2nmG46xugk4FRnly21jfnhHmQuE/mX9Yg4y3Y8thqG8+F6Q6r3z2IOkxUKblK
N92WxcT1GAh5lPqAQ8heo5vlT6TvQrhw6UEMEW6AhcW956lwr8Lc545US2ruKM8A
WHzzch0uEtd23+fQ44OTdnu/h0sdSWdqIiZabiv5KI0a88Zu/bysiahFNFqzik1G
PGl5xOVUWnlbH9LFm/kCds/eH1vM35jgnRGwKsTB3EbxiJQKK+FM9fjjHhNKUS1n
j+OMA3r69e54hx4vhz7hAaDARTBaehGxbYIZ+/uU9moHUUIWBhcnLGXuLSBetaZ/
TOXNWVEOvGncjISGtysvpjBUnejrs4KYMCmdI8pbKaiGd+XRYbThHoiohyxMtoOC
q7DvBRQ3ifdJIuQ1MQWPgTWclpwOLVHnFPQjKhXhFceeNq7i+o2c5mTgi1CHdu7V
pXh0EQYu5Evt5WWLGzCylcZ83Im8plhMh4pcbTSYyXbdOsQYpPe3+3foAL3i0UWH
569VexQRUu9hxwS9AT+2URGRs/VIlM0CT5djW2GewKTBoPvLC/beHezBC/InmvNm
/jM7YGOSoKteGFlam56EJHk+U+BTLCxSOK3ZTDDCK+8pYdiTQguxbBBbEGv1o4jR
7WYApQtimwhUVwyrfJoLRBSFEvHKZNTBPw8/BZ4AxpFDhqYFhTUpVJk6+LaVxsgF
HZquUXG5cMaODnFVvTaeID22psW1Mpr56dJB0V6iwh/s6iM77JErlt/Mg53xh67+
z5TDrdSVyNh9QY7z8BevYJzuoQqP+xSjCiwQeDlYgFUWe2TY+ZpeOhNEGmGc6F1N
U8UT04NnBIH9jWhhIWvL9OhZwNYpOHRdTFPm/IElw3Dtu97/Wf/VQ2r18RdjKDTo
jIdjYBi5cu2LIBTLIGvoeb/ykqjkbgGo3pFjiyEx7brTw2S3VHP5NDx/bkMmGTqV
F1kFvz6vRrf3QKQqonkUNO6pehwRqjnT+S9nTBh0fws9mcjH1fVL8f82s9chUo8s
yrN+I05u+kQvdnD742++LZ1fsKk/kSRTrJ6UI3uElTNwJZUZLGdSiqetovNCS5hy
9T1u6GqkLqQqyiriNUV3M4+aC2cOJVq4Gq8roUxs6Z5nzBujd16YawZy/aENbF4M
uCaUr1WN/tPMHiQSzMi+Gh7MwnT0D2IJ7E0zWLMp408muLtJha70ycrmA64WNPuO
XiV+Tx0tE9K236yQPUs4vO08Km4eWvK0jC1rS9f08vwejEs7cKwIEk/91uRfpm+g
WDlLb2G64sj55Po7fyVRZ9dF+tiYsZH3X6oatGVA3kMk7wvuOaYoyB+BaEphucgx
Odw+cy2Qy03UWlBGZNki4E4et3MG/l1Qr2Gh/VyAXWclX1tgW0LqP9Cfb2sT38t3
c2pZLdKHJ+w0EvME3X9ilIZlj2cpKXnlUW4tdTQLQ3OBhFq86qLhMTbhPh7/pu/0
Z7SXFFcdqjwdaZkDZk3m1Lv/N/sKhesixXHXCn7gr2CPKdeDh/MNmp0vhTkOce2Q
m95mvTC5VMAzQhPIG2ELGy4c3ierFZdTQw2cXGf9lpg3pdfcTJlPFV+EnTR5w4lR
Asf8IBti5T7/gtgdDj02oaSoBpv31gp8p+hk8xkG+isiQLiyt1PLMsfmr8fdDSN9
gKim/uO6eRc3R4g1yeKvC80bFb+SIoGVj6h6BU87ha6RAae2ctKuI0prBMMHcGTR
YxrYfRY9CKqLXkR0skncUkM9StOWTGhgbe5PEEI5MXXIZJ5EAce50ab14N/7hAiE
oJN7ihXcnnD5PoYW4muugb0yNsqQC8J7DAbSr9viNH2/2Yshcp+7myvBo/ta3pMd
epcXL7MLfzkSE9UJUlgBHba6yzZ5jdG6LfDI/Ea4W9x/SBPhzj1THDGCMbPyvph5
9WFO8YxOsVOpiLrPCBX2ZudIZFAQEdyIVPUSP7jslUnkNe2rhAuG94J47igzEA89
6w1UzXJNCn0L9UiMqiex55MCoAcCAbJ+yLfWKKKLpIul6XPbr+o/L7KZxDtcqQLQ
BVYiXtwwRIutZ9a38BmHeS0fIJYBPN4hjRRqHZo7JAwSdrEsXgj+p5A3KxaqmAqP
gWZjbu64OT1KKm9LwMuGsQXcDvMPGdd6+60KnH8ZL7sOuvtbFbDFUu4LfsiYUy4Y
9W4kqzMz6/gFOYhBVFkVG3w4lmDrBb/kwhdHX8GmCFERazz9K4huWeLe66N1nEtp
TNJWy1bN1pCi7LOXOdWQkR4+bx++VAJURIuV0tWiE03Lj0gKYsepmo5HfNesxWqg
qujzzHPqdNcHCEDsWV8k3jBgPv/6dAj2b2mxxhHjojDMUR1bK6adnkHRqjlCjjWB
QywSk5K43yIeUonjpClj6thgF8A6isFIVgb/kp5ky/gNq9Hs9N9M1Au676O0utam
9ebkerzTweHsK7g8CIUlcpyXxqsRpsuIyt8jL7BO8Dc7pkIHrGN6L1jxeq6DiciJ
a1P1d8wEygRSMCd456862MU55tcgmRWE/Ro2LMvTzmPlZo7xH/DqzqfzVBnLHmoD
ndW75Dwpmr+rS8J/96MBiOZaJZhAmwHZfUrliiMCon2cA+XZp2OLSJF1Kbf8lH/v
8Du2wiQfZ2j1XOlkhStJT2sXbYOQmxJmghQEuPsWKPkrQVVlcld4XylM9Hj7PB57
ppyFUFSzJFcjAn663MOOBKQsOAUJBXBU8yU/YPKp/WcuQcdjhUTYNWTfIPYnydG1
GnGjxLFPrIf9H0ZTwMh5oNif8iMWOgLb8UM84bh9/q+PjXiVOYwd/FKNZrJK1jdy
aJ4+fPtSZIRTKay79mCA1IXEKHlLfK7+EQflRgHSFkuMedvMLneHQ4wQuOJD+k7l
pe/hiYGF8YLmtNmNnYtsXnBhVkZd1UqoHrg/2POV/cN6J1izBH0xoHb+PQfN4U4w
8Czd+rb7QyZnPOm9G+YNqrrH2ErSUoLqZFa6u4GLNMVArdhL5RTfTlEvR0JQKwE+
kDxU0I1hAHTXy+t4VFORKDYB+M2mnt3nNLCqbDXXRXdl1CMHEzXxh7bB2pkK6y/j
CQKXO2dtyxdViwjpa1cLPgUG4O7nw5nCIrA8UCPAwV20vtrQlzyL64CDQQftKyfO
tEgpvJd3FILiPsYLxeJpvbcHM6niB6noXfyLcs88mPNB/+MYJmUxOWKqmEZrOTVu
y6UQQQY6CQRleZC7sDUpM+9vuxDFeQEv2Q+OoaW7CzZG74kYrHRDQdHfISU4eoly
fCcBAsAxJ3NTWuenJeij5u3f/C4Wg8JHqoc8uH9OxUC6zgx+ZPILZj6tetzD4Cv2
+CymbHGq3ZqbR0AUqWHoio2TWVwO+olCdOTmmnljxjLqYTApeNWRqUNDXBnhOV2F
8StkjW6jXe8LYiM2Q7eF/nyrfL8ahPVmS/CBXky5yW08HM4+nOL7PbmnzOEFOrUH
T/j5UYtVTKl+e5KhQUBeDuzDc1YvQoU/hBRBBQ4eeQrIxVnP1EY3s2fUprOF9JYv
wV8kBPW+eR92HFHTVcE3vhBVd6W6rW2zdoIMMluFYf3DGdwrBacCr9L1Sl/7pt7E
ytO4B4snst02F9E2gRBTZM8QsVti27acxvymyykxOrrK4jP5r6O20zVGNCbyyuHv
yqwZcPxrvvYibUA4vm03ZXxmYljzdO5fyh705gcNJ/gMwXHBpEFQl3nNdCWh9yHZ
kcKS8vRU1VJHP5VhuQbJWB3vg/JKoLoaVcVErynF3nQHdtL7EODGBqLOIIjeD4MD
dsCOtcrPH6zu2GVjMUyJa0AoXuuSa+cAxsKESbWlUMLRs5OSlOoFuHDMFGi8b180
/4WJm+DxIa9zY7kvULHsTp0hT7H+oWeQ8JMAv4A6G76J23uDFPSWPVHLV4XiBWnA
gaOzbIPYl+1yUw53nmxs9GFKxSq2TrSApVTB4jjVY2VyCDHweFYE2+x6fr+FQm5K
IAIBiZsBDvrAOcd8vUGYamIHE2MiyY6lU4tXRTrZu6LzTfxWAvYMqq2U/NSLc5sn
siXGm5+n5XWY/bJ6QwHghYgvoIwjLkqTIzpP7AetPYy9xJc9pR5gYB8RiB7d/uzb
FyWCUCTE7N3tlfe8FWWXI/7yDLUiAJiF3ursZyApdQvS6i1w4vBuxAA9P8d/K+vl
N4Dm6uBla8RkpF+1oMhJ2EvYTKXCKCHgnFoDYq8uQv0iHESnqpF1+fePnq4zB09k
OW4BnpnyFdT5kUbKAyQlGOmiWVo/eHyjoM4I+1VFLi9CbKOkt7XH3fIt8tsMcmS4
PDaIWH3TgGK7uBWwRWzmlB6/jlsacm5Qe/mT/HH+Sv1WgFCCyPJ0OWFSyRR+Jx02
dTEbDnCBZ6JfufEpVVETDO4lxevnuipwVT9WZtE/nimjtNR5TTcuEWVgVrrgKhPL
KQx7tHOGTReTqPanzqW5wImOK1RKz+L4g992NNNyZM1za/IR80w7BgAH9yNP3+2F
U0yTzapTnQ21/06bs03XEy1Urqf9SrKPs+4mOKUmLZPHvYFc5APOw9ZLIuQuy4hD
R7jCIRj4wxFqvLrnUkepOR5N24cCIqP4znj+l3IuapRceD7J4YyoROpKTJzH4R0T
LQeI15UETypqXaMnoGE5mDrd71iQZ8AfhvoWM/VDW6elp0nBm8m7Zr/kxIM7vZA3
FnwQW3FnR7YJ9dyxJrEC+C8K41WvqMcTmvf42Erh8yGvCHaA54BSHebNfbyBo89H
BGwAOC+0mKqHoAeqVpMjE6P6uf8Xb1SiS4SdRticXkAtONgVwUnoncR4FEwAODYi
uNpvyBMsPC4DNeVKvxMBMTnYb+6D7eiM+T1mj7wTmNZPhTISeLOAH7+obzOFr9Hk
fKhbmNGVH72AK+TNV9YSLQY2g5ueAr9OBVa8r4z0iIJokxAX5GTtXQAhkE+pff/C
DhoKWZGCbgW1CZIqBDIRUg==
`protect END_PROTECTED
