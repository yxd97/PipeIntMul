`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OrfhtLBx0iqhYPphJiTuQk3jt57ub68kqQZA5Nv01qhsgyvMc/72p9/o2RSfd+8V
KjSJxbqMNGXQTBAUl7RrEdXQ9lj/bMIgUWXUKhwfxIE8GPimk1TvlySQWfOxWk4f
3deyvThHULEFbGqYtdqtU6XapC/gQ7IA/UsD1fP0HNiyiKKalfpNjQikeE7x6vjg
WuMxhcyRz2yRbzgom6CJ52it6x9iMiu6eBxSHT8rTWACFwQSssHCAssjPuI7x0Gx
HjYAnC4wE287S4FTiydCWzRpe2XMOV5lu6ttjM0+uG9wWwFwYML4Ln9ZPtnyAIcy
3x16tco6lgBc3w/XVxVcSoSzVq81LmZ15s/aBzkfXEy0vOYd5vlz0WlzsjhWJHD4
IuRGRBjgSHR1atU2X1MUMf7eMVZIDCxWpkB3z6rsMlcBZ0RbK8f0WliHCFQIofIf
`protect END_PROTECTED
