`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
prQcDd9ibdg2OVUQU4NBQuzkR8IuCRy+LvgBDtZgYo/qQiwTs9pYMf92z3oSly2O
2xqdz2naofAT31J7B9mPkjvfiJBsJ4kNf3yM5Nr8rG8dDH4y81KJHYTwcl15VH0Z
9RoasqwS9cJ0t2ZmjJq8f5SdlJeVniFzt3GX+MuzfYDItheVq+3Nr2IHyC4g6foz
FcQg4a+JlLaIw15lpw9xF32vmJk1Xraurau8eV+jAEdDP39tekJjNi0z6Frdn+cB
b2ucw1EkE4kX4kbusx+b3Q==
`protect END_PROTECTED
