`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5z5K1EUKvy/BamU3COlXyFz0If+UsahP221MigeRAdWhatJjYmC26uooRYrkIuaA
SEj2VqRo0c61Nxi21WEbq7yXyTlYRRMBtzvNkD7/PpVdUOz/6r4XhroTkkqhMeJ1
snhgiTiBm0mILZ0O3T4W8D6UipdAxBedfeX5NsHKURTVew1yKzUogj0/u8LEgHQA
7WQ6fthPNT8/SaZXGCFU8kkcEuz+k9dtwMn+jp8YpN1RpNmaayDE9AtDMxD2+aeg
WgnfyRNd7xBc9pZqC1gs7DvxIwdERQ238ecWsdC1Bhnx7/fY9vmRaS8VuwMA+bha
rONssj2wujNiwiA7QUPXiNqNNwx/fskXatNCBw19j5tqPRGhHXPGHQBh7pVAzd8r
MnuHLiIvVxbNguNph6R7hxd8IJv9GGPV5PRVHmLlRujiqt1Ru8xvOa3+Jg0tByzI
JiemktVvGNe2vJsErzvQ/DSqnCEbCJVWIyyMrvyoTQUEGjuh12uIrQVyPqgOvyZf
qJASF25Tp97h7CD7lJQoK6NB/x7EeJfJvEt1FbT9KZIf+pmfm6Vj6lD8OSzaRS23
35DnNValn3cqWFTLMl3RQzze5j/aIOSK26FcArYKR8v0d1GeE8S4ulTAEb4uHE1K
QQ2NkwxA8bKC4CUW4xxFCxmsOED9n2rgzzSPStORAcobQAUIgtcE9lpuxPYMcH5A
bcl7DRPlKhnThuYFWXHKIwUf/v7vgY4YN4F2vo6zg+G+/Sry0GsR6KrIst686T6Y
fInz47txcm0/bL5uB7gpU/Y/pGItnpeZjM1h2rcvqtpy2E0Z0CExSnk3+5pDFCZY
yA8whwTa/hxyEVwhLZ4cq502uBYgCKsMIQ0tUkBbmq/rQ00wpn1XGLpv2lMxsv/J
L/OxjQai+2qJ4apEaTInX/vWZ092B+y0WMfw5pAvyLYTZOBYLQ1gPEJ1JAHvYx9V
4MuOlZXG2vGfrtFqhDlwXntteNf4Ci35nEA+iT0Fj6+129WpSqV5OKjpGUp22q2q
uFL8dJz0L7G+UN+mBEiPZnClviYdvdt0GeH0nTfFUrKOQRjUO+mCHxweaukyrCG6
SvNn4q4JbWFzc6YQipalBaxGg9rFVWHGbqrrD4KG3xyfCSxWLs/1yPxFODA1/3xo
RKZ8tY71ZVV5ul0djsTDU7bOPpFfLpoCU67DStc1XcjLocPp35dk0+K9bjxH/qUO
jL+s/jPBZOOMGcwiTWupNQ==
`protect END_PROTECTED
