`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WBi1c0YHXwBs5S4fEQ4vu9zJnUQaz1DuE60F/nv6Ty7onockqWiIhVUj8l4QxCHr
UD/KVY9e7y7qIRTrRif0vC0rPpNY7/2ohAaqKdM3tDPT3ucRmFDdHTWlSe6LCdlP
vJeLdH6iuwfdKBB+LxEVjn4yL9Xc65tfvSalscS8rZPk4HASe6qprDglMqGq1C55
9FUm+jhQBqquwI+7ZkgE0pp/DSwSomJBrbPtClNqW8V/xd2CDa8WRiWvE08prKGI
DWuXL8/ga/G9K1YOvAyML/wGw9xR0PvQUfmxEU5RG/0h0Fiy9g7m7ALygEFUjfTG
sILTLRLmYzXPhMPS3V61iyl1PI034xWAj5wfTR7E1R7pvxzizpi1KScddLBy/0K2
5Ubb4NGMv3RSB08fxQdM2l0Tmy9tQ3j8dIBIosVrgOBbORul0NpYDLCsNm4TtVCX
276sMFa1yp0MlnuxRLyReTprrVGtYYPy8R39jLLFABhErSV3Zcar0BVkiVlWuBDi
LUa7tHq5XVZnLFZprbo/kkUay5+BF5C4jI/syRVPCHbqIejXLBfi9Ah4PpkHZ9YF
cX6rGUncHErwkN2rYYECJ4YrQmuBfH1dsttNRpcdgJQlumDX17nKhal7ZyRsovgf
r0fNV6zKMJaSN5nnWeTxzMQTL4c0BDK58tlnJB1kl0v+bpK561ebl3hx49otEUrG
AGGGXIcNmiaEKjStXv2Z77QjX1eBA2cs9vUkXEE4wNtKtSb7OWT0O6JML3jiIuTy
IDU0NWShTKXgFx9kHoefJw==
`protect END_PROTECTED
