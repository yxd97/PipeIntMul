`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZL2lcWbm+cQ9RSkp0JWzGrBjO3tUKuBamQk1r8/IE/jH27yHldvuwOOUaoB1qom
9QsG+ByeUQNsvF/hBfIoLFHCUthsiCLmI/XpAddSPJxtwCcKdRA7CPMdxQR2SyPK
qS76zE99zEySeT2Qq1iqdYiF+CsdsZCYxnxU+pen24n0uzREr/1RwXbVrK6ZteuE
7mydMyeZD/k2vftx2QUOxXyNN9A+ZaA8SB7ffUhzbH9hWobFuMwWitL6tiK8GR8X
eLywk3Z2woU5S+yitdfUVsqQvgI06sVwGRKNtl2p/Vwe/pveLBWnzGYQt5mXLjE1
UHbNCgWAaOL3U6wWcTrKRA==
`protect END_PROTECTED
