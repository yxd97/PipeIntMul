`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jG0bqbx1eZHbNpkkCFmGg6p6nCTnyAwHq3fDalbjaMgrFQPK9mKDPheW1+88iLxt
l5DMdqSVYbvtaQK3PT5bPj6lpqPph8uQR4bMV8G+6PctY1ukaEx48hM8PSzT/bjD
zAEWThyCNcLPFbS2wQcMlp8hzawR7uyQA2UMKQLii5KN5sLfR21qLC1LC/Wwnw6D
aY2d2AoqPuoizdvTZVEq+b/jVTG/utOUaZ4xPk83/8Ngl87M04L9Qa1+qa2Gw1tk
kqk8YRQvxKdyXGLNxfuYnyiz0/76xYw/uFxdKRQVwDQOhkMN1y1UK6DrB/M3Q2OR
eB4cCF5M7BFJ6X1ISzIP/K2O2QgbCMJFA9SWPI/utYENMFfXlyriyNmz/qdCsl1O
upYSsHUN8AauWmFvrWZMg/Zyq4N+C0Czd6ozsYmu3xM=
`protect END_PROTECTED
