`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TzvDUgb8XzOOhS9lo2vPrS/o6bnCtURS+Gglpyz60Bov8VLp0vDEMxjtjdeG0oY0
aRWANFPddVXutdVe1Uv4q88N5fVeD+zk7c7H+Jb5QeZa4J1Vt/rZmmlFAfWsQsCT
aMsyTBfULKxrlVfIVIvNjP2DUsbSstG5ANSflLoDrZrcpOQobxrD/nk2GZgaMWwh
cvZMsLH1RHY1ohY6JtxNtc9XGkliuIfO3ngBIZpu9B8+5c58C6rqjee1oPEN6PQW
B1NIG9dBDfeR7S0tuGaLcZ2yIfNe25Gycfgb0Ec6p+GYlk/LxH3Pu7OFtTXdTAqm
v42eUntX7+OQgPNG789rtA9Z1+ff/bzkgfb45JgphUwk1MYA58OQG4cNV0KFjL7u
PjfMfEI6bpFQcNt3KVAPsg==
`protect END_PROTECTED
