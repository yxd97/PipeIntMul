`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FItJzsle+2YIiIEDnMNtLHBNwxmEM+olnXDUYINu4FODSE7jn9ml9G7Yuy10kg9K
dbk14F3AALAEsUKEGji1cG5IVjlAf/rv7WpCJTN2+C1ok1TBIM3fpPMFw//sU2iD
wEPNP+5qbz/a1c0wv+mT9Dv4MgNgZDOmaBLV03KhD5nPvuHYLxBpKSExgtKWZwOC
wR5Fj+UB07dNHezAxSzYMC7CRBnA2d28uGY7ICF0WIT6hn1EhnU0PxoNkpFyDW3/
x5WPDtvQPNn+hMuZ6o43yw==
`protect END_PROTECTED
