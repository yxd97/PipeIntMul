`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rQn+DCEVaS7JUN1ZL9xtBoQ5XrcCBURHMIqENsDe5GJAbjDt7oCP7YXpKcPM2Gc
VJwWtmMCGAu5ZCN60TxsEpjuSPdzs/Y3jmy5VLjXSthiQde0Ia79AxNQrGtjaK0c
Km0nPLJun4gNIpo8OXgD8p0U3VvJDWHH20pWEzeNwCRY/h7gJMEbDASjUHlwirrF
Yfpk7TFqleZI/6FPMOlQm1xhg75ac+uHuc3wIDK/+h7+JB6rK7+NhEymhN2/J7zg
Xb06KZKeB0wxDKR3Vqk6c5sJj15NMIW4ojH6pLoR8+nmMR7KyKX4Q7g76mH7J6MB
k4eKMX8oL87HcXdIhp2iNVayZCh9XQEyafmQ7+AQvekQIcj8uDtd3YTTZcLNvemY
X1KrG5ycnHny/4EOawzzQsa24g6qoOpOCzV1waclyFs5NB2gWW6UOy0UIgnzmE5y
DOhr4eXHljj2SFn3G9q6iPzd/3zo7JrMXbPnb0v3Wwh9p1C25uXT6v/JdK4oPbt5
fN+HNanI6ZKMCpKK2F1m+ASZZoOeGAUoSz3SGJySWLmBqzr2eUWt+fa4S4L3ua73
6J0tJTz8VR+xBtQV2S8jr/IKJt+jZ4XIzgk2A89nc1LAyPLII1UfSrEA/SG5n1st
luqqYLUYTmMiBNHlXsOgIIdO15E+hbwcKcg/EMWs9xJg1vUNuFr2wxKC3ubfG6ua
OUxD7uT/MY/pPndX+y1q866CZgixbtrwWDzdYRJCi2jUUAdck/nzPhDvhXC/ae/M
Qn7DagSQhfums7VvYQhGRXb9JsUfoa2c1O6C6rNWXRiXqFxu8yxeMz3IpFxRqQrU
c2JCH5R00TuqY09JuudAy+N34/ej0RNhTj+v6u7wpU5gQKJwZXKd8vR/kzPz+eAK
mQiykygGlm9BYPrvF3oT4UrODssASTH1dxYqmK1+rC3lhQ8NCwnUu6LbpGmYmMGD
MQghhHi2E7j1fKYCnCa+oKt0Epv03yUQUWphU0IQiGlVVWz5HNhC5K5AjhnaXXfd
pQQ1X4270TZBYk+1GVwxU++i0tGFmUtx41WhDaBlVcpcy58QAomA8IYvlZ4mPiWF
30W4JQcaE/itjfX5wDmGK/Ef8xicqw8DMVEf9am4WaxyL+p1EGuftL8IM6SIYefQ
4OmB/KGwZQI1zq5VR0Lv5I1V4G6yx1Tks+2PPQf45yNdgXNsIlbx7QYQZc60PtEc
7bTD6G8GXacvdWdC00ragUP+KaeykXWNtCFzuYwp7pZRtfAWx3+purd9yfxxwvdJ
htunFRhElZSMtC2y8dl6ppuJ5f9/LBRsl4KDnqZuWN63Uy0iQdc+Pybfh79D+vz9
UxAhHaRDClxtK3eY2LBOdRT+0TH1iY/4Zbb0c9XyWvZ8zVTRojcbZVOEkI+6AJdR
wyG7lN/yPc/CaKP5KSQ2OqM9cbZL7bypy+OmVwp2b99uFVBxQPrPSH3MYnx+xau4
aguKe1EcI7nwxGjp4qpIMiKAMO8Nb6XvGIdeRjYh/MofC3kGPEa0FFqLC9GE8UhH
BEOp4K0FMCLRMTKtOwxUJ719ajClQNUilvJcgYYAmHZvGFJRWawYGx7YO0lLSt/Z
dG2VUHPqS0TGlybyzdQ73rwp6wZLuCP5K0H+JNDRm2pZuEVnuELtaRWiU0gLfy2b
uqUCnN1Gz3lbQAzvISXs/m23vViYPAAiTIoEUE856iGWh85fYhjcYsGNPoJo3b5k
503WOrZi9TTDixTp4QIGCygEoOP3FjQ1AEkw3MdWsf5vRa+YteXEUnOz7Xax8NUK
llHJtsXXPvwLXfqzgh5o0FYPHtENrjOJjMJRJ+ej5qSc1OOZebXEAFlBSKGl2Ta6
2h/ObIbPVJWw9skgtlXFJCnAHslkHQgo+1D5t/MOZPap5wDhqpuHPOft4DqeRHRP
z2Vw12vvqtzCoD+G/dP87MeknSlu1FVtHb8jWAIUwD5SqlmU06SNtaiG0kgJXB+M
/2rq1dhOADJKJeimmLP5gewH0cGLLQivsQsyWXI8YhyELllv/e41xjIY+1ACBkO5
7iRxm/cyvWiOLIrJA/UlMDwgR2DLyCqoMleREWYnXzrYv5o4Fn4IIa/x58iM2/QE
YXh4YbX+KWhIEfD4Ur7XXnE7m7XKNsTExjzITbXUAsOIybnITUFBb2GQSndoYDAZ
JwKmuqIIbEfmTeZcpbdNS3ldy9n9F11JS/V+ZpzIyvuObx71nvaTIZ1cZDCBsTGM
I5vfVS59wb14t4NGkgz6Dq38c60bt/3dB6X8W6TIebOrgKZULLbQhND+nDAh1peH
1NvgYje8TWGt7/Y1KxzDM8wqFrsEjUxjKhP+hSjbN9nR2tf8LlZV1TXVUxM/VO9a
YEG6Uu+seUp/vRvlPsLBS7I9YWKITezBGwMEp0jL/DkeNoJCY2QLIWufG4PnIqNf
pNS5IBX3HOFrq5f+5Ot+p5pT3GK8k810XGHs/AfP8sGhdQyOhaXzSi9EPfr1FnHx
Dvj72o8mAlixyaBla0tUFRsr8Gken3Sstc1Yzs/HBsYrwq2VkxqG45il6y+iIHG7
I2xyDHgtef7UCExmgVtUCDezDa+qtws8fRAchkwfCcl7r7PtOHzKD8N3bdm888cV
eDGjF1uu9nTCuqk2yZEB81IDgSvGbKUrm4fYD30PuvWNsqERbtoVebnZFLSeYnui
OJNMR/Y6XAnl+mOhyyyQVFw6nM7Cxe7BkJ62o04Gh9vVYA2blivzmUrUqaN3VQsT
TyJ5NipnqSRoT+0mkha5ApK8GpkdiYBD8ilOQGD8iFcUaCDAHIY/JQUdX4MJQPA6
`protect END_PROTECTED
