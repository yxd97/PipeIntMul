`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41SAPj+TS4MVpomjafMuTraqyCWtHlaS9pW6DFyqGMtiTq1MIzc6CpOnJYwM/WVu
d+9xcJQLp2Ls099UvxETVhPn0lfjEKKp3HLTy2EVubw7EWImb3Q+vADLXmn9o2Jx
vD6HLtJdIl87Mk3kvWmR4wMPdpb7isPY9FWrLDui9lFyQkxkHFLvBQXuYVRO9t64
GDODi5oJrv+hdwoNUvmUhxOovVGI9kWbZVlbYniTFcBMVv7xfQhCxZf95JWtC+qg
`protect END_PROTECTED
