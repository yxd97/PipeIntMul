`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1G5NDu+0uDzbu6Ks7ypYNzpDQZrZFlC2ZsigybJiRIxbUfonii4K1rD78m7pJlVx
SdDqR6YV8rNBF8zPjfUTnBMJmrhpNE3rz7ox7WSG8tcFRsOBB+yGmUKfFmM0nYeU
QYPYFM+NV7pBFA0m76ub/BrWtIurP5ozS519UiBbDnQdhjo3VMhHvKSx62qXI7ZD
2GxzyjyIm7fJsQQR2gtd6T965TkK2FRb9VWISqKPgWgUPrVKIyq9ky70WqD6IjEg
+InAClcUvGBWz+E7SwQK+v2Rg+naLtS5anPkO+D0E9X0VuXijVPCi5Pnrjesy6F7
UfGhWjI0i5i9RFTvinpW5w==
`protect END_PROTECTED
