`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQCkFXTWTXC2x/r0EBmxJ+L0sgE595/DQ0QLsHDUbF/YJ3yb87dMoCq0zxRCo0dY
xPQkyCagzKWnXW+TXLr7071CW+evFTEeeOYM4XQ0gTNfTVZChb8CD/0kzqhns4dR
INFB275StFGKEK0RFEDh+OzuvQ9c99Auq9e7N2mq5c5cPUa/5K2Wfd9Fr0MERGnx
Z5xZABvYwZPkr15OxmZOVAgiyYPA/POUMZStxrHjq9yvvOH/AdCV8TyDAIetYT9C
1sQtWP9IYlWQRexCxy+P0PL+2VyOYEIEKSKV6jSVuTfW/iKG8uryt5ACjzYCl6g1
iHVLyxlrexyUktp0/jal1SGw3dc5tOmlkxhKzzNJLE1odjz+pCzGSjBhuOgvInvN
0zB6OPA9+ieYcTgGasMa3g==
`protect END_PROTECTED
