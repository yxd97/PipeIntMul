`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HgRNTqSSDEK4YCSuDRD2mFzb4O6bIWKpkIWVc3uLbr14joqHWqjqEqmrNnyX0KDG
LfGA7WKQJfQ92vHGmJ9QGMrI0xoRJs9IstS+PIHNMIDVl9GGJQGxS7nA+PCsaLdm
q5vWktB5XylVWyg4TqpzbHyTpElbz/atDWwvjd0wGg44oVhfNOfagz69MpoOkHVr
XJ4qVoJflBGPX7i1x0nOiOJ6MGRslwddLJK2/KoN0w6d3C3RWnG1GAb8orC7Lsku
VdLSYKIc+W4+eHS6bsP6Ripn+LTe04tCrJYRTNbhL0F/5RseE2Nms+fKGMIVJRz7
sdNvQ6//trQyR4+MBI7RE+gWjdM+0dSzJsA4aJuyTXU1sOoQkpPJ+x4SYi/UvFxv
eFrjPQwVNw+OF1sfQopjNuVoZnxozNh1xy/qMyeloRfeYPI5pGnY9qTyW9nPPknP
p5i13p/e0H2Ck5Qup9Ke+j72UzzVIvcEbLI0oMNhAu9cBypslEduSxldnS84trpf
V1iFWXW7C03r0L1YpcjT1KQYKrj1MRUoLKnNN2mb7Hl21n38yqRtRI5ls72+IoIN
OUaHUuuqPoBZZfaaGmatP+7SOUcWHaV+eWcqJTE+cNg=
`protect END_PROTECTED
