`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
186lpmq2lkmvEhE2oF+8rTnlZdLyrHkyj2I1S2Ddt6dPmOMWfkPIEejc5PDHeVPT
2w2sPvyJN9smmOVwufmVXNMNu1CywJb/ZXO7stJUhdOb81c8I8ApJABoWO/b0RGS
IO/o0pbwV6XxjkFPePrv2UR+Kl5WgfJ/w96klF91x2eqEQvyX+zCAdjp/2xkbOUK
Fh/8gGMQyyiPecq/cDFsue27v4lbcZYaQ6REtNesNFaKFieVLBzpEY72IwH+ht/p
svEu/Eoss23qadUvm3w6h6rMSQM8XZhOdFwopuE/9hblR0eqy4AoIKGdB3mTdQOo
ZPha7I/m42zUNUBnX8a71rhFheC4Mm8LQp5AhdAuAy9KexAcmfziENZJsb2Wf1ks
BQPegy7wi9lP9pK5nkappro6tQ9/g7OrxkPkO/69H0LxLs9RZIu9kWboZF1kJhVL
pT7NodPLY7868O50At97Bdutx/VCeXHnPFzkYcIVDiSJVGA40FYzfzRNVqp1yIlM
Hb1wdE3D9a+HT6/Au2ianCyszGkYUWUlmNjVlSLl32QNYVrgcFQAzeD8L41zTdmq
//Qhag71jw408pfIsqcIOQ6qNI3FrEKsXj3nGA4nMY6lr6JYGq8Sxi3NbgkM6hdf
3IHzH17RjGDwK2efQNveVi/HLsWd4dL4jAJoTYZ81vY=
`protect END_PROTECTED
