`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4VS+EeQbPj4I1cw9Fqq0kL123zZimFVnYvFnszPX3Guj0u/Bcoc2QNsFXqUDi/b
D+tnWB1j2mfFkRk3Wm8/0P6dCZrvvGtGI3gYhEmiRoKevRGOv3i0R4DWsZk+Dneg
B4GvdnDBXtFJB9YfvsEuDn7p8HIvJO2NMXENRpdoJ3odHRmrKd9JxKqDwt7sqOjB
GCaHzWrUA4o8O2noP8ICL9Jf3lyHTmReJ+6/WAFnSsyOSZJ6p0ok6ZgGBmuioyq2
84MhOkgh5STnyj1j0gDDh1HlRJ9+waannRP+mpPSddGzqcKeiGDyT4QL8WVPNWbW
D4kQ3oUHMwZkhw2bRjdAzQgJjmCSU/ZdP2EuufcEPF89i/kpBs09CqXnJm8RaafU
cZsrFluy7fI2uJ9W3YLDlyydLQFMBVIaapbwYRA4/IV63z9BXAG+N0+nfwLymn1G
5r/EU5WzE6WaHq2XM+TxnDJ6J4b13e/3XlFyH4ytxNJ38vHTIN5LUVgXlP2sdCXg
1sVS3x5Ubvj2uLoI0oW18oQczpNf0QsbAHx1BOK8EBP0DfZZHPmjfzkdQ1QaIeuo
FbjHnHLmUwIrgnpr089br76zLLfjUC3y0xefDG0i7GlmG/4xkuNWfVszdIhWO7TO
s6OiwGIQDcbbAOnzfQVY3g3WVBTMkRyeXjFdXNRPHigwEYHCxFnfkiL18jjLRZ6U
QWV3V+8ssTJ3uMncTQXuu2LYCTN2fi/zBdgq0sRwvxaCEJXOfQjWvyOJjl4/T91U
b7tR6fYp0W1u+n5ClWHabgcywzNTsbmpooQ5HPM9myFm4ZXt+inmXGoK2/re5NAg
KYXplo088wRqQ7sV319Rpw++7+q2nZZCVGf0zVUZSBpCLVOvBsgWygOo33XbcsUe
IL9Xu0gZJYnsN7V/m3H+dSkXS7w8gU0W8t0gN8Z8K6xVOKXN3eC3URip/YYX1Ldt
TwMBbkergSVQ94B1w6ZDf7HJV/FbxA63OocbVF9Fjbjva+OB72gL1tU+fUqLJUy2
N6wGo41+LZsjeBc92M8Gn36RfzDA1ZssA3pdhITOOVLUEICN5rx+KRfr2Ud3IN15
duQ/QjfokJVenwcKkC3BrsHZjS5N3WHQqq1JBuwx6gE=
`protect END_PROTECTED
