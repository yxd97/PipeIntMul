`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iC+2KlGcvIMJWCEkZztbiDMIG8D6ChA/C66GljkpMez9ovv7dZynOaBWaAh0COTt
wxXzKxzEjEgSngKrTm5SnBLX+tG3EqfNeyrgLXL+G/I6J9+IEOte2S3TaBShiVo5
r016TjVAr71wCRf41+vapTQaRjWqiJb/LSQwwzA0EQPeV4vIDX/KWiJ5gaCF/Qe2
SSxEHKqmL38SbdLi7rmXnxKrvRdU1DjDTPBJME1DQxR+XeAkA7FrtxBqVBDcEp6x
T7Y+DyRD+AQXq2IoRMeMbG+LQpa00BfY/okbtJISRYZwoWMtyLDdF7BelS1GdYwX
GJ+H8AWDKx7PBoYBmMMRGN7C6Sy6xrS/QiSy2MAt2FMVXful7yB8LzdSe96u10fy
8NNKUsyPMdEO4zHJDv2diXNmGXBqQuP/7vfjcnmXR69kZ6BTTIn6NrE65iFOcuWC
cjeqnt9Tfx8ptg8zy9FvTSugw2cF1Sa0JH09livMhcdelP4xHRXihMVXJS1PLE7v
SM5j+Z9nPHSSfxNeYG/OzxxmZK2OWO5kNY4dXJN34jZJ3RpsOM7wWQGr8Stq0A38
`protect END_PROTECTED
