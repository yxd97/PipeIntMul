`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glQ2zv59EkBnaZ7da1D0GjTCV9FCO/q5DYas2xchAJCsHbcULxSeIFRxFZq3uqCr
HvTPHrbtvWcUaNjZyNDP/2/eSx5qwwRgImBETaMGk/cqm/q64QGcQP7uPSdzeJnK
xqPPbuWOl9aOWTzZSNZR9Wq9j9b31cHC7RyKYAD6D8qYGoB7LIEeCqZi6RRKxoGy
2GZkLBdtZ6X7fR5Yi3Z1u/4WLHP835tgG1+VJUpGsiCYuIjma8m4lnjdXH8MM4xe
1rEzCdwW92RnB7HSNJeN8arFu0nhhKKRhJ+X7EzR108aQkoz9pCfkVE5RfY+WtB/
FaLdOtdma8ZzCgF35T/4AQnZxy5rBQxhjyF4n/hqQ8tUKuap5wntsgQfou15gIaG
4mpGmKMzJIZ9BsTddn5eYT3wSro/4XtgiyUxNJu1Q/ik4xETqSNEZeoRj4WSqem1
`protect END_PROTECTED
