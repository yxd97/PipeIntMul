`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gGMWHqFnNS7aM6Mqoze0wee6kXYgb9gl4dwxm5TlMVRn2jo5r179jXQ6asV2Q5lv
w+iE+X3g6IyrY2xI5IdqApRzRQJZAleR2ujyTd1quBTaD5J6romslT3FXIHOb1KX
e0eKCe8YySZlRAPZZHwadL9Bx3TYzV1zZJOSEufpp5Al6DvSLrJ7iLbv8vFpqztA
Z8vVvQH6cPGgG/bijxrq8u3ver5YnoZNGWvFMY1q+auYefC5QDvA/c9GWXBZ61UY
hSxs9+dmpQvew5Xwj6h6cvRShwrlOmCSWkleL0O8mNcEoilkyE8zd5OYdHIKP+6q
eTauPtOeE2mcTXS+qvb4oaMbiKL8f4QcLoox4T+GGjl7oBOJfe9J4YZf1MiSlKbL
nOQfSMWta3vqqydAM6tUx+stcdnUBiLM2Xkc9sBn421Vm7AU7Hr4J7ZW9brxGOqD
aU9b75l8hOAesK22KhQIvg==
`protect END_PROTECTED
