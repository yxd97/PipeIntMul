`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9XKePGckKAXUciBhBRWytqSSSQKf3hMzLiZTLbIy2LYQtb72DCyvfsDSInxzXZkb
c8Yz+7QqxWb3l0CH64qQbnZbM18nbUnQ+nSctaXZJDNuAJ/8pZyRZcNoAP08TgXn
o04XTXL87YZBDMRHTrg4dHcpN0/0keCBuESaPINm1j7MUcRp2uH918Oche7fy8GZ
L1HP6vusFgcISNQhNfeSiIX4mzCitI/6xLJ2KygwT/qsEmKm7sFTYbKWvddXzZkX
J5A/RFfZpLWGaNxW98whoOtNde3Mn0jQnyUeE7ecP46P36JNqmD289h+0sG/st8+
6pZ3dRxC2n9kdIjsr0mTygeTJJ/MV9IL7bRFDO+EAzHZ+7dCVzq1iZkfwjJzQfIZ
Cj0UIEjvmZAnGbN5JVmGNQHdaxTfZ3TTLP9tMI2WuX8GJHAkXqF69uBUzGQgK1/K
`protect END_PROTECTED
