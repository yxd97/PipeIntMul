`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcyYpgduGC7o9LNBi0VqkLGzcU1akrrU412dEfF6jhioBpQhTR8Gha6XIlSvsfdX
MXfp2qazFj3t6mIRGQ5X0N5tmk1J6XBJ/J1qxYPJQlh1LXV66fRpkEPKR0vqZGRT
rEQbrOaIeFqCbc8Qmly78OJaGFIPAqDJrZ+GqHvl30l4yT7EueHXYtTpILRfg7NF
TAA4iQAMMzT55P7sXeU1pcKlZEkaatTdLcmD548nyJh0TpgXxVbrK41yErT0gSXf
bal2LpborijFnClGpqXMWjbLXj87H44c6juCu07Q+qdSpRqvGqoU9JlH3L5FLmHN
77PopMPuvkBuX+Gi4lsEZTH1fNjFHTEXSizSvsHiSxpQ54lFpbhyBiq67NqZ99De
`protect END_PROTECTED
