`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i6JXMy0EgRMU5vO9/AQkJ5P+Q7+hp6YZCDFJrGTD5bjRb7PVvsMV91DELnnmf+xa
I6tTzmeMX0iKgLJGGxDxIyq27fufAmSyBJYL+i43uPJXtozH0RRPDOx2E8VaSSRd
gpYQ9KIhzZXcDylF5PyOZ55uNXi+D7O6LAuO95WOtJn14j9xmC4HrwWenBuTBfG/
ovAUdE5NFO+TMbVT4wiScjrs2V2XLFe2m//tpc2PC1z1jQW9XoKO48bdV8umsBmy
CVM0Jt3JOXm+fYq3AvWfF9ZZuPkx1kR9rlG/JgI6/dPgivBqsn+nw2NQn+GZcaxH
1v6zEwS7/0vZx2rQo4RWpa+1HEjHpwBJg5sCt2UJw0tF/J52/FCfJSW6uAHlEY9d
mK2X1IJgTilcl0FO868ZPdWgrprtQf9FzUUYhr7DxUfOA7AY1HYpWYskSJpcg4pg
QlMHKfhFQibkNKb/1MGwnx1iU2T1nBgslUbkTaxPf62LsOwNDPAdVgKy0gjGks3E
rqmD2c0Bh82B8cmfnjcPvT5PINhEITHgtGxB7DDEgG5Wnya0WhvbY2P5mFVBVMd8
Zj3wndM0E3SSNXW4mu9iIRxLpgNujNfd3xJNF5DBsOW1rhAGD5G11FRxggPcGX5G
Y1NE4Tk6SmEvehoOtHGMsl8aJJM72KeOCwfxvYNW4JbRyVD/sG47OesRxlniFXGb
+w3G4oAG6jLQPd8pRskSBQ==
`protect END_PROTECTED
