`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b3RwCtN2L2B1NUzlHtrVIX6yXZQvHufrcvxwqnSJbKS5unElBBRzVs+a1bT76pTw
oMRyIKjxdRNTH/X/W7SQgT/2cs9BwBf3tbNujQxgAvcF5I8klOkjUhf1axzJ+Gyw
OBVIqJ7Ym4Qp/Q20tkrsnNEaluqs8IhfKYXjwF9JSIRkYUwqKNR5ig3D5qbuBMxm
sRIHeK8eL9IUBE355tMAz7d63GuHMCi42bHHK6mpuf2Khx+3ZtjQPJZ47iUu+jNE
H1lZUeTz+veFfZDh+hPSMAwqwHsCWalC9QMBZduCWP3drGI3JVD/VF20vt9H5t4P
oFKNuxzLj5ZBwkZODLQy7kpcMKoVch8+ARDmkU0IGYLz6WHCkD6K/C3201BUn8Cr
dJzlxDnjg8gBfpBxdY3J1g==
`protect END_PROTECTED
