`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EVy6cfJZWo7CObERkZVzYvyJjG6oMh+8kH3a7caBxdkN7LvoJ7OW0ia4gI2plp8o
UDZMDVsr2d1l3323jDzBiBGbDoT1/3VJYwvwIHPRup2k8edkGSe6tTXHguFDuG3h
xAA16wKy+ceC4O93Iy5HgbrfIi36EfopcDX/8Eu/x1jHhObudVxAeYBOLQ5N1UV/
DGsPwGyfXouH3tYADfdSu25LTCYa8WkzOn/ymSTTQS/KWITVG6hVR2T/BTcgCBu5
pBKKMXgrmQLwzwq1lZlF0uP50247FP+V4TsKY3El72o=
`protect END_PROTECTED
