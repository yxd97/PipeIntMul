`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e8Y8xqc+be3yxLcija/pGl0/SksgItyG4D4FYqXVmam12f7P4JuMWwYvWnrgj9rv
Ch97DGQUUF4e9JAmguz+Me/rxwhENrW5D4L2Q9Js0HMC8yQURY1ol3s2Bprs7Hlq
1uv17lyB8/h5Px3DOGp/HwRg8JrucVVt15gO7vRrfK+LQ9yAFgY7eXekUq9F9IeS
wzZ/tifqfIxc36Srq6DhtLcpxIQYr6JN+7ZPcmHAFgQIcBucZy1D0sVv/qgnW1fR
sL9gWckr1IBSSDh4bOen4FKnI6QbjNAnoC7GiXxg51tmJC6xP7pwDV7CO50SB1y1
HaC8jfJ0W4kEpLlA7IbDoHbMAMAKjIo1l3iFuHbb3H84yf8Xu4tk4UTYU+GaEdww
aZ6pIAyj2IFjmW0oZj5ZhkWzELgwcOSmOXZG29zIFKk=
`protect END_PROTECTED
