`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFwP8jK67wIO6BHFCYwNuh66XEPxugdks13psnx2/F698MCb6HYSGKvqUZoSN9qQ
krxP9UrWn5cGXhwB497sQOuq4+5pDmrNTBeXuiueBZx/+k5ocCmfIWTz+dI8tRQ+
zvNRDvtGtU95hyITnZIH59ILGqLDUO19WNET67e5XDRWkRm17s8wthplZlrP4p2U
/tJtaRdUhmSetYuK/dsGgrg+bbUGeKRDgD3Yn8zNJnx4xMyZoKutNnHx+PwsFrTC
yxBXCQ5InGdSS4J7AttS1YJurTg6pv7ApZQMatEFByWr6R09MRBhPkFH6W2NhYhY
Pl7ErXVArmjOsShCraTNoH9zP3oS9f+d/7969LISenO7IxeXZ29me/FmLXRZvJTx
HcLX6+a3ah/OMcyBZy2FN5pMFgw7PKrTQbnKDoT4/O6eyhIBBxati3U0XWJkIdP6
TPvm0nSEiMa8a1SS0deX8P0qHUwM58fwNR8SDkFAi8L7Wh7+nwSTSg3MEQOiB3Z1
KucX/2BMQQZh9AZ4y/63h9nmpONh/HPKYjckskwusJi5d/clLtioZmXNb/SsdrpB
wGVP+pR96o8A0Kn03QyOZYnzHbkLbKDXHMbZ5VLDcnUWUbjAftyfzttr6KGsWqOU
awgLGkoaBQtUtxFV8RKLSWI7gKPXMintly4QhVfuzidb8H+TsYRPJ8iEduxRjJNG
+fy041Ehc7OFxNct24/wABbj8aIp3HyYO1cm90/XX9oHwyFMw7n1wDOXqr9F56Jf
XIoLVcj9XnAlLx9bKT+H4A==
`protect END_PROTECTED
