`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38EKXpkqja+BKUFAA9xXnGcpa/O49zaoMtPPDEPk3KWn2GPDLvSwI7UeXInamYIx
4Sjkx+Fy2rHdGQDC3Br2xMqZ2OjY4bxxKwImfeHI6uY84CMuRsWZ+qWc+3YdLUCN
z3gCzS3+/gYpsT9/58sRW/JrgHiD4TECIKoAD4Ry3fkstF1KOyN1jGHIz9guKtnv
nSTNwtDkiNfK4kDn9R73WnK0qfZWsWifXzXgsCN68i4hH4xl0Dv7uOGkY9GjDnbp
ORv18wGKJ1pK3v+TmjHL7bAFo1fU8ikOLWQ/oPKql3JM/joRebxkKhsojbIcoEPg
kjTmemToocIf82Cf9XIiN9eR+fomaq0pEMxYjUCl7RDYK2CfZ8F5VtbLrhgWyYMD
OyKuumQBXu0qs74NkGp+2GkJOqdcRz03M9G+54RHI66hp6DHxGnXXfUESFLZ1Nrf
cs38CUhfnDy2l/OBMc6BzkHQWxVu/N7ykQJCQArJAPW+HfG1NKqE6AgVP5wfl7YB
2rJz2em/0oZ4kway1g1e0/pq6og7Xc4rYSOlSkO/Zh1xcWx5Fvf0+CLfpOyBmQk1
kv6B/nHhok0TSLh6Y3P9Y9oWiWy8cMnpKP1Q/nW0uhm6rRz3UHubf8nWvHH9mW8R
wD3hUmyk4ywW9jk4JomB4w==
`protect END_PROTECTED
