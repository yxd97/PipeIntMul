`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Jbdra+kjLs81LWuA1o8A9WraAAPjV5Z+uYS3gC2XG5qu3egirNe2oeJCwh6fCC5
ss8YSvmnuXchJvM68mAsHc9DAfp2acOAFyRH9XJZCB9Y1jXNa6IfW5POYP3MxRnf
5yRk5xZB4tB2dSaMj2hS0zuu4jK1RbMN4Ke+KPx7RLZG4vbhszOF1Il+p5WtyK12
ExnqcHaav7at9PLAnVqZ4xnbgYQW5TYUhHCynVdSHbjUe1XHRrq7UCrLrFJ0/y0+
2h4IXyj7OqY2XWlrHHzaDr8TfzXZfLSNS5FnvQUCR/yOODOeQtx9SgGlRj60ysZE
mZ8GBgKU/g/Of+cVmui9FfB/vb6q3JcBi4En6YSZdY3zUepjYq+OwIwY0FIkD3wE
j+ZlVg7bSpFU8+hCnNkbb3VALr19+5hD4MVGFU1+KZQxUzg01hSBlqMSLD331zqS
lAPYvSbSXUW2RIcDG3tmdWfKUpwYylCZn8IQtWQd3d0aXTrZ8slTTLX+/OunyuI1
xBmmLqQE273Vn9mhpGPPBPt0BG81R9sOI3u/NdTJBfM1vbXkmXOLPedh6ULjXLjY
uT+c0Vm+UGh6IN1Wc3CZQ4n0gHZq+mAPsqdsnsM9eT0a2WJ+VGHoMO+PG6v5NQjs
MQc9BXiVqIaAYLALs+wQnhHIswvX0uxTV8HU8MlYmr3RtUQx+da2QF5/FSeQP4Xi
LWI5Ku7QJDpspthnPJPOJGWqJQTqfqyvRau0ikcqsa8snxhHvpkQrxeTeSaekU0l
WJAAKbwn2iXRiKrmotpsqvLMjLSSy0CZgiZG5f+mfGTqM4KBmys2jtp3DWd9LZfZ
3QlWybmIgH8jSPvqAo65yl593kNoS9O8AImytygZuW8B/8G9rIbwr54lu9zo9khw
WIZqTMY8lbsN2AXIc94qzb2G4mhdaJi46FmXL/KBkVpx9rFaP3v2XnMRIQg3mKRi
8iTW27cfNZW6yzQTUV9v/i7ff5AiUxvCJHoP2qsHPVQkyWkRhdKaGJV2ERFMDBNz
ZL96jE826NlpJwpeN7h7DO9wtylZsTojmnNssK7/IPxF78DYfRjJRhfR4nyXqxbL
m2XzOAaRwZDhUK2Fe5qnN1r8EirUjodDe3FrZW+UcwqqZsZNM18TM6IvKo1bh1FH
+e8ZDBVJWFmiGzkKFnGtoBvJEqgXZ6jUuZNIcv00a/EBIZqrkfP+zMBds+vb4AYM
K6KxbqdXCDlqIoBja5YZu7pusxLJYuZCfZkxzmu0q3i8uXQVct/PKXSRAaZ0wOrJ
iDqSyFX5emqcOc/RbVEOiG1Crf6f2lqKAYfSq6qu0eGGNxYAAfQNqwLoIPRAFyDy
K5d9STDFhiK/6H0Nc/cH/29A/f6UY4Ao4M9vlTFeskaKit3TKhJ+Mg26GdbEABhP
dYlqgAWb1EduaLyybjiePdDUIvuqbQUjPB0Rx7MPri6UZRiz5Jm/oaOCCk8RsBkd
SD5hPYHXnSDIuutc85DT+/qXR+UUzMn6EUIf3VZxITyDmdVZrdN2lYIF1N1FCe/V
kltlY2t245sU/MVe6r5FFSu/T/u+POYlTtbNHcsmn2dqR1nC1lQaPfevwpCHjk8a
tBlmLKplxs5Tc6SPxHFNa8i/OURBV7dR78VDW3KSnScGn3w2c46fsrCwkIWTzPhG
rxALPC2OGCnIdaFwr1H9IIF/H2Aep8wmsi2c6ATLVtXNAuQdiW3XXlYoyGKIXHyr
bv16mKjleo3caV2h0vTBr5luKTsMa/ZiuIJXlIG/5xl3fB+CrGbacbmcOz20/pu4
lqEelYtNXl5puLEVqc3POjCd8UzOcU1odVZUorBaads=
`protect END_PROTECTED
