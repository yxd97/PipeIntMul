`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eHrZOKt8xSMLiJ4yY5n5wVCBykxfTGDJMORzbQMPcU1S+vDyyYaqJIEYWH3xVxGB
wQPRsoD0yhXgXX4mYm9gFPvFvjOdTznw4tIkGCO29lnQg12617lQiukrBswGG5+p
dd6YUoje9howbZ0bRegindh0cdVut/2ImPYZ/cPBt0cyEnvofiFW7Up+npxGB7bG
jT9EnQUrCMdpCNZl8ZHOoUebOxBjYjUsawn1a6PSruFLvq6B5F9Vf8t7WAOcmId3
TExBsK2LoSFKgv0arW8P5miA07lmbWRGcmJ33kcu4vaI8F/hxa8/WmqjGHdo19KF
EIzGscs9y2XnzPy9+GMJf1qWVPT/D0J8AGyzLMo4ZvCM8jeeu/DmJSlkJpHXlMWR
`protect END_PROTECTED
