`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1i73KkRIS0Bk3ZS6rwjdj3NCT0anlUbYh7M2yzrvGX+l1Vblul3OZi8kKCwtSomS
odQAFbI1Slc6EX4dnKyaOpozyU1EYZKkGZ9b/08MZ+gw3ikMSzLg29w958PYP34M
sJ2ydSI7Tgt22So4qnjLgRb9yGjIC4kJOw6XktOrTu0Wlp3sZVXCKHKpMqZsgdqv
7CHiB5kdxp3s5WkeANOxJRCj6I0R47EmUjXLm6w+vjz41ZFqOMUGfXHBeIVwrQrb
AEHGh0WPyMmlNqPk5bEDVsUhFAKUaohuNuJ0hSDxKqyFFWNKNftFWZTPwU5V0wxT
ArJKz35sC3F/ZPWxNSb1QFPBUM65raqOKXsuZ+xWGir/lu2jCzebv7qjwT0fTEaX
KKcGb2ifR9Ok1TkK5Pw+nrqbpS70Xpq0bHNyOKAEqzc73GsIovEcL+8rSGDGRWzW
qpyxw+L53tjtbnzu/FChkV4arkz2swORxqzwGyhiZWEji1Oe+YiXS/avrjQ92MJg
GIqQmFM58oJTbN35sCPILq0jTM4pAy6HWEpdR4bCLYvLLzgJbh8RvZ3LlIviCzNX
2iVmrslvmLcgRTGbnHMR+wyyGQHi0Z90AsaIMXp4c358P4cokiSrH8gA/9c4j3sK
89g38HeU5aXznceN93j3Sua4JR3gwQ9yjF1e53psCAOfSEiz0peH/k/1efboSI//
vYfuPzLXEL3FAHum1GGUyomeWiLy5ac+dQuimH/zIPbcppK8ezFiBqPBPqG+vpt6
8UswxsomdJ7AhPbwyapWjM0bqU5B9YDp65ZyE5ppA9OTSCQPEVXBYz/0eVyRjlDT
Iq5Sgg1V04p7qUDHGcp5t9kbSAOmkSa2Oj1bFstXxd1ZFsOgNrH18XPJp7Lqy6mz
5jqNQOmIAo9Uqel0n2/8Va92XST9xDJ5MRxBrmGPmIUXssxL1+YmA/pdgwxpmYU9
9kug/7p/5GUG4ylQ2Su6Ww/q7VrkE2P9bQ4cGUcW9Fidq4fHKkUVwSHQqfz6WqMA
oV3uSk+Xi57irEvQKMCOr2wpWWAlUH05qt3YKKNKEPovmeus6bFJjbuUntHmsoWN
T4cTQZYLL/nzgCjg8HWZwmx9MNFGpl+o+WuPSdL/1GMvV5jESAEcyIizfcBIvoFy
TF6xjgRrcQL85FvDenaVlbiywwpOt6+JVRfuf8E+CcONl7j1QvX5W5/puVFU4Krw
+XXJyIMQhK4Ydg+JWfFGh58I33yAo+x6XnyOWGyFIpxQ8wWsqQDDsa4+cNhvphfD
Yg3tNyeQpYPy5yyHoR+pBINehm7GnQR4JOgkGdPGj84+E7cGnoEdFP4IYjas+7UR
sn3khy+7sqyis6tzFTPgFM4k0bddgffDwsZDJdaZTLeq1ha/GlMetrVb+WGGxLfg
`protect END_PROTECTED
