`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/LJJExYLcUzVtHEErOn5V8Omtj6JW54SBtyjJQjwtUJ8fL5aCLTpY3Nrxno/p1c
ZvjPc+UbldcmRtihoNv2IlmMdTGAbZgsjwIrA4GbFMl3YHDrNjyuu+hbNX0lQEVk
vxYvn1+OORZBfBsYbeplskQu7h7y++EINasc/BGL85Pvne3xvRpu7DRXyBgrUGwT
NR9DSFVt4yqraT+LfyzvRHywvLfFPrPfyC0W861QcAvmeJT2ZEKv9MTnbrcTXaSl
JkgtuCxcVcSmhoCchxNGTZFQedcmA0woAqs6AYhy0S4Lwcrld1PG/goC0dkVZmqe
vGhTZAmtOmnJPYkQUJsVK++4XuapFgutwOB3EtcXtjY4ZtGb3uVvpgGdQ6DvHrtS
heqI1sNwocl9QI0lfhp1oQR92ByOZNuPd3hxzUy2AC6XTPGLLfaa20GEpcUJwSEg
o1vZQi7EIuaUJ/WUWX6Ul4/DSOJLmtMl7Lvyg80PCVeohuYVvRQpPdNDYHpRpKeM
nsPpxwsFd7UgLGv8MTDF71JPlT+/kb/wx+pNH5DOKJx8y5MnMOSe4KtbRL0ZT/Ew
ScI94N1aMfy/7e3VKAhjIgyi+dJr5iBsI/U90fJ+qANq4hfEoMrz5xR8RoHJPz/F
K1HhMrbfKgevh0BLGlJTnZaiEsEcyEKEEcz5ZyulBsjcPu6a2XWys8CVF4/m6e5i
b5T5/wL/eJw9Z5li7CMeKbjdJfq5qKpVR/1hXRUMUYHex1wWI40a9ucVKNyGeQ3c
CEUuEr8Qr7ZWCaf+abLcZ4IjzSZwffQchR1pALsIzDUIxZS2TTSPlnj8TFi9vfEB
L66MvBuLVie9jUgCFPykaYzLW4dzKQyWwsPL3VUdKR7hXpvyIexw1/gHQp9gOgms
DLRYukaZHLqIDTx4CdHT6zDDVZdktqFjNurK38XLBO10ybnNPVYx0++/IJfme2z2
KQ6JZtfMTphOp6hhcU65kkCbAhseaPvbKt0VxTgHuvgu5a4p7Hcep+rNnH3yldrT
l3FVGqECCtvjbx1K70D7bSVSDiN3IGjNKOtsfoImd5Cup0zTbOvKHAv4Md0TWk6v
k8ode0MTtZ6gx2aYi1Vx5/a0awxjv4UP86QhmBMfTTKiu3fi6LRFgrsSoBsOhBhG
NfBrnjNI4n0kujhruMRYblyeFx27Z2RVZFX2jZUyh3K6tNqSmoALH2i5g+c3EBw5
10W/bRkkUiVZtfgpZ1lPkjBFsFnDniNKQieFkD4iEjCF7D6y1rCXAaXERUUgF7Tz
2v/8xvZqklQiEZ2isYKWUecfbS7lMu/LyvXbXJUV6vfHURifkM/o4Mp/1T36Wf9X
l/6FHjT7eFczzQdDOVN4Milvqtp+PkOOcxTfEd36GX+YDPFwWHupZQLVjmdYnk6Y
YauF4PvcI1TETlAKbi07sU67iV4cx3MDA11WD1XkV6INeppsSttuSIaqcj7eTT5T
l9Dx1lai9bkvdbH56jg+fYWqG/eoLauadfGImu39O7Wyp1LO/3QLSPAZaRS9cF0B
9CPV8EydfEckfdoNIPuwgMj1AYwqJkpbVyMlJgHuOQ4BavXO7QFJOMkCyWkmi54T
J6drZDb3SXZkE993PRq/alwqn1Jg5XTMKjBXd0UYdWEQ4z43UzFk3S5S2t9RYQsN
6puApcJZjddc9PuKmYHn6baWVCIHJWOI8MjyEmN2b79kgjrIoyWIa6NlsiS2ShnN
Y+UoHAqavqcQyTbhd7oBfKHJP3gkQ5MorT9LLOXbs3TZW9NXXxtw0JFXz0f2+HFg
eJtROBqI5S17SaGagtQGCV+1sluR+hQw9/sxbSvZ9HCrd7DzArTXk2l2DBkeBXtZ
76ybw5I/X211FNX/R5i2ESqRwWAUirlVf2a2L7Kh4/29Y+2ZAHaiFhAVkT8gKKEr
Sr45vP+uNf1/XpeH3FZ99ikJb8SUbE0z75m2hNfAG8bmDEA6/3lrXop7XCC3hr0N
xTKRxUB1FFZNVDwEeMsS8r70MeY8IkIvj+i6PLkhW3DeTI/9P9Jc3IrF0pmBXtAt
PUt5vB39gM/HBQZpVxZtdcZcAm1pv/qKDPNAf66jiO4zUKvNJlwl/wbgDpFvqFXh
GsIuuXGdP5oYqH3lLZ92Fz4045rYsO3mAVhbRQwotFwdRX+yLZkdev1EMzyFD0Sm
gMqe7QFgZWLpqhHxFu7xPJ5Y2udnp6A8Da/hZqoiKg+dKIXnB7EXKc7zTex2q11Z
aKJ13Ytm8p9In7OtMU4i+Or6EFfeTYIgFriW07XpwwaOKph0nmE0eBkr5OaazqbW
Swld1aYsLnqwcqD5mLlkLG1O0woIffcyj3iGI/1vesxlZxBBqwpV7rjljvHV6QzA
HDUT9l1AWsejr5SEOfMe3pmj3bZyGo0G9s9VvbmHVdfMlxSDXoPWJN/EIGoXIbvc
pbHtYHBKyItUiRwaI2hVvWto40187N13wghP/UW9O1m+zmZk1saTXOTNYNs+sUMO
UkhA9cvgJubCNlwiarKFvEs0COh6B/l4IWu+K/Hm/vZEBqIoLW5QLdyDxtjCjfrM
/oiT9tBPC3Q5OOYvpYf5XIJ0Oj5/xGWt+ZPZ9U9ikCdHyzZNdExP1GKG5uj0vLqd
NyWtL6pGuYnmqLcRg3/gty025cd/G5ORVD+/AQR2z5pHM/G8wHXvT9cSoNgTxNt0
P8hiT+q4IdVnPY6CgTPDegaKuUx7rcIZGaJzJZZUT2ihE8vCcFdAjuDon3au+Wdn
`protect END_PROTECTED
