`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oY5wnJg8w4zTyl528oHBNETrlLOMoj0U5srUWJ5O6p0AtWimM5j6yMmZiwUqKypL
0bmPLB/FjrLoUMqpINBa4XV4AJXLBVqw4u4+SPVDCMcnLXhYwJX4nr7K5ao1gQZ8
vQetx1m5iyj2CTniQSPD8YBtwtxEaNGvUCawcOyDCpIXfVYU8lsRc5FgE3Zwyre8
M6wt80z464sk061J7khj7xO+NKn/o88smEGn462R5y0hBJn1gK6DL+9O943skkuo
y4Dcd782vV2pCYM8pbX2e8OqjA1ncDJCiy9MprWe4Y1y5tzIO9YV6T0Nlw8Q9ssy
X/vos8NguGYLk+JQYpdufF57PaZcsEiCCxzCc/IO9hssUqzEbCMgaCBSyHyH0n26
wSg+RgzyayOO8ooZFKm79PY2FP0rIaB7hvFZNmFUsjZeXGPAq9pV7JliP3mfdDOu
XgPYIFHQ9gdqzQH4wDhAe61qQHxEhYZun4aGXUqVfSpJlkXsvprRzWSf9UOeQ/oz
Jw5dPsHj6iM3d/1Tw1mUhgQGETOHIBXacTPHS4WSAOY0ZJQ0vY8N0WjXWGqtHXqT
QXpmR1WGxOmxXZIgul+8Q2uiGSjI7J919AJzXFQ0Az7any6IgSWQb10U+B93yn77
SeAXSoJ1hD7oMmDwQsnLnchynEF8kS/G0HqTgzFjo3xDqAtqvjNCgQ6Va85QsCYD
OuyQcy1NI+lPRRsEJFzlukhTf6ar0bLX5zME8h+hFg2YWIlqsSL0gt9iVCbAJCEx
sD6f/U3Fk6gOoXdplDwTsA==
`protect END_PROTECTED
