`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGH7jsIivM846gYfVQAd89hSBcUgyatlhs1lgfFFbBecLDNy7UD4oHoNOYCcMBJi
kMjgzsWkN/ng9we+OCdIzIVd932cUt1G+D28TutG0xOgXsv5T26y7PiktaD31ouB
qIT74kCT4GvJrB1dRW1D2XyTHfaviaSljgvskKyVRQYYF/TxIowB1O1VnLaAkH9+
V/P/8JyV6NI3SflHIek2xkM455Ye8gAUpCxt7oyJrGzoJPE1cxUhss19S4aJCK2w
EGekSqCIj/qE+k5qA/4VTo0NHHM7Fmwb/XLNOng94FgNu1i06If4DwRoh0KmArxb
CsEcU14VWh+lYzSxdjvkLUCsYJwat9V4jPRxfQRD2w+12PGyw8CDCLJ+868kBIad
HnHN3BCGTQ1uqT9f9/TAEVEgd47/62dBLdHonyAnmxi0y7VCjrWX0jBXlrd83CnW
ZWLovz2j4m95ig4dIx1zhMC9VoUrxgFlD10CTFtwfinck5HbDLIBcx5oEq/nyv/0
prQnlEbmXoUBSTECoGdw4dXBs7BAGYkp7F+I+EKJvClvjtrBwWP1FlLzV2KpPOG9
FYi/4JVkIaud015MsOrfmCX1pjQP13Bz9mxhESl7HGM63miYhYF6Bif8B1Q3sWVk
vxP4o0gcqtl0NrgADQTj+HZMVwvyfwwrbgVaxnFfC6qR6pr+imJ4Q4lwWMpBF0r0
nvCfH/TDYhsmjCcSaMqAjkz6XsAH0npEapessor3hZ2s56K2erdhIpzYiXVuZ53o
WdhCqpBixSbF0Obgfe1Yay6ThF6yrHyeHrpACClfXHargU6gCRM4qhPLO2E+tuVv
lV3oaWxAUJvm9ZJXIX2ZzR/wBjHlN6Z92Z5QUwN1DKKojLkJ/nLHqrWoGXG0mfDp
/zYBvVxCjaPpQDNF09C2NJ1DM6zlrO+LzzXfEoeH2u5zXphfmb7LjybIftzV7x5M
kEyaDms6bNyWurBExleiFyWfTvBYy2nIPyOi/7EEDuysbsollT2idIaEmjZMmsbI
i0vONtMZLPJhT+QdpmlahPEh+5MqKTZYqP83iQVwEXZ2UsjWAphQVPPGBfW+UnW3
sW8pIq0OJp0aAmVXxSJxIZuofT3ewm6sAKz78YFzszHBgAli6UbSBkZcUNJ3Zngn
wO3aJD7U7ZNY+ts8le5VpR1hQr9spRairc+q4GoNmg7X3eKDHf7h4U09rtUrah72
URExjm8kFrMOztDGNI/0iw+ASYBWoL1GwsgvXMIYad/R4u5Z8Mt6cRrc3wFAvnNj
sK+F/aYVVKO6okSExUWXa1BEY3PjJzgSpkEPlGFb3zfVCKXxWJirAZIu0909FAhh
XVoA/Tb8ccQ1y9XdtS6mLZ96jfJo/kwBZzNjKb+bvqz8p8fUThvAvTa7dXITj+Jw
fIv2I+to7CsvohHGXEKmfvhV1Sluu1ogCSLbAfEXr1NuoeVDCjgUcTgHhQxxckWj
mV5kszCd+AwpnSXHEkn7yO6cme3C5jncE3YNKqW2h+9hqp1wqTUktCAcsbZaNOuG
6pKHfjS6aGcIJOPV1zhwJ0p4jNYhky4khZbgTeHAiX6OsheboptDQVP5e49VuxYE
SoUFqtynfZbQRDySKVadcexAtPuj3vzVF7osTMxs0CYih3MPC3NKjCatJZQtCXvU
f/i60TYeqvQ5Tam/75zZo8/jmNmQkYLKNuSUpnwf1V/6p/7JmvqQlWHmuQjp8kvx
1vBzGpT+FOdpcdCsjfZnBvRbgqYr47ulJSrdt0dUGfWBnvoHr2i4owLRr2XQGE5F
J3dg81owaW3cDoLsumT0VUIP7uYktKyGeJlX2AKxxVhzyd2N8SrDKYd/CJSKPeVB
/TM/OhG6cYGxLlV/N5r13RGEvsb4sIjnu3S45oS4dhnudzdRmEiwQ0jIsDAuZEd8
tEIt2uqHjnuCU2Wa9oJU+55mNO9Br/md4QCSZy2r4IK5lY4ZYeXufeTWuzGJQWIg
guntK0KkC3n5WGjVpm1Am1NaaETuX5cdF9hQHRw+iaRVKz9McT2FX8t1fzgWKMv+
vr6dQjs2WXpYqa5vAWGvBoMsAOk3eJ4sWpVplQuaFuJD2pzo2J6tkiTO15HTz9eD
AqkZzSXt07cjcE4e88aSic6T0J582irbYGe+kNGhnfn5DRcio5G4ms49MQLljmAr
TO6Ig9NXHffRUpuZdFDQ2WJiw9Azuj4IbqxxEcbY1VRfbWTdTcme7q8sDid7d6Ug
zQInKmuv0bPmphBd2AaAgvQp3WQ7EGVTt2AcVpuOzCoqOHQEfh9H3HOAxxKqdurb
wD7jrKqM47sM3r1vxhbqh5vjZL3GX48pXsOgZY6oPOFmk1Hb0LgQAHuEHwPNEmTa
cNZ8DUF6//GhJtP8bGlleWuU6iOVXRPMGEgC/XbocDRPszytksXH7FPzvpaHpMJ+
0w9VPGHpzx3mbG7ZYjRi5t/ajhRb+zT+NnMWPtFcwF3vBYd8ahLnK+UjDtEPpzD4
zktQp+P4qLzQR6NeQppoLWoISu6L0t7KJTk96RwtdzZuiPHrdG32U57e7Lodg5TN
uIbl9dPPDnhprjk9SPVX5GeQD+GjR2q6rWh99VectKWdP5ObuFsVYZcJlu3mYvYP
Yggau3sEQJYMrZDYQjkAcoNL6UvZiDQMN5EbdCMnmUN6AXy57XONPsscWapjEjR+
7hmkH7q11StT9L94a+4HO+wrSQqLE/H2h6WKXrxf6DA7FFfCSXB2MK+28n++cFgj
hYn8DhPuTMeMO+GaMmg56BigfDjou8rZRCxn5MUyMhi8hXX5zk7Y6PGZzKals+CB
zdwaCnqcCEg8eUENgdsc5c8fqtijbn5egUGUcUIqC2q9ynjcOMK/xlLIS6myhT/W
wUB0F43CF0UCpEPqU2CUT+Fs9RZWF47eKzTygoowbHHNDddjhfMfTXI/fs95YgR2
xM4rx2OiXE3jdPEhCyX6kh2ilScyt7/HkNWLVeru+BE4tpNcgo3U+rLOsDEu+xFN
oxm/EQxTYc0GG70B5uc0cHtlAHiTSsDIuQPe37lTbzf7whLRmzhFs6NYURGMfe4j
U0maU1WGFOVEE17qfsFCGt7U1seuucArXYxEHtUCKE6oCrdblWl5M4vaNUmyGUmT
`protect END_PROTECTED
