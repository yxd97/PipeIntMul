`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OBI16hi5Pw93ewGNDvD5edgmERe/RKujvQJdzfzGE0qPVhfIGmQWHvbRa8YhDRfk
wEjWfxkvBbNbq31Ycp+XC5mA6lvJXgcSwqfcCrkzm9zV2g85kJBuBYY/l3DyM5tR
Scp5M1UkB2useebcwDB4d3gGa9p7Di2eRcwptiGv5Zy9CGg/IMqEi/rpiQik06vD
9knBXHFij1CthMXYVOzwsbsaMAEubq1mk/Y4bSIr1p0uZGZ6CbPppRsXRWFmfsz9
ly/WicR8MkMejiPc89n/cPxC4rLZqZMaQyhahfMVpMOLtnHDFoldok5IkWohbsVk
`protect END_PROTECTED
