`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oRzZRNsE8Ys6uSl0vtPq7mWnWqjzGeo+ttYRVThrDf9PM7ZzPlnNOBi7W5UNkPDT
bmXuMKYTlFlDM1Zsbv8M+K4L8EhsIaa5JVIF+yuRGgb7JMWLpsSXv8HZhzSoMwNR
d3wfDYWN2kh6DZ0UapsXWdkeKdNHMRo/aAcN0tgKZW9vNvNkrg2Y9jnV2j1ZIQaD
YPUEi/TVTxeeRVW3Ky2tTazb2Pf8F6eXFsb2r/XlW/aWnGntwENEvo+PmS39+tfk
LVfMPS6Qa8R/Ijd3xQGbb6/ETicdOlBKGJZ6g5YfJfP35mRQeK/iCPXhwbmOI4zz
W1YWBHeAzMIpkVN0uvxsYf4KEdKm+JqHiqAoosaifmFy48A8Y+WShJZMfMyOdgkU
wNl+IZyIEH1UUmOi+cxFuG6S7XL3PerUSaoKuHwDa3RsvKRY2MpDb+PewdznIpjj
D1LIHmiH5BSwdVQo0tvhv0GZ1wjeIuekAqjGQxZEZuDKn5p1dJ0VOHmQOArGmkg5
16dxRfb93SxXuKmzZlTBaIAhfel3PDuMjIm5c73/WDYFq8NgSXzyLdSl1L6Uhjjq
OeOaDGdokfkMoXkDIxyWNWID12bcW3xJ/VMWJKF0MatHv3byq88nD1gNAHMuncw6
x9SJXDLuISpcKjUkRLWndMVBoFKYb4BabTXm13NdjI/SQLf7If2dzxpk3g90iW/y
4CcxiGBS2DLpkC7HstKWcdOS5jys9uuXDEJfp3YJQKhG+m6aDKwBR/T8ijS7DDFj
21U/FKjDVkxZtch+8XdLBsRtd8smf1Qppiu3A+m3e/80POpo/WTJQwZlUIhR0ne9
wG5/P31QDjJ/oW4uBwnoMrhsGRBwR8BCxJdJJujb+7qV5oFre2xKP9+x7c7F2gCe
wiXYz3JY+bWbSATs2JtjkJAxC/1l9KUqt+mkjc7xISK/urzJ0Zc/l94OwuPZ62ZE
bI4FWiAfPd20jLPLbAG4ltr/cCNZ8zc/rXHctsCcoKh8uU5oioGjvC3OX/iCRKEM
g7ml1ScEYImYGSxJpfxCrAMx7sRFiHf3NiD/vMEjIzdKZuet248CuCiSzqrDZPJf
VhStr7+Vhejrbvadq1CDlPsMEBLen7N0AvxTGRHDnkVv0WQ5yGXpD0JetZIZK0zc
tnnPxc/RKetdSNGRe4+qldi4GLLbOCGca4ySmNLlSmlB5g+okJzUBjAt3Jeu/Rkr
dQdbM6V2tIAh97D1jgIbHwE+sjIeJ2RS5ChNAsRfPX2/OyMs9RrPrz4Y095TdoKf
NOCURISaRcoiW/JyCdSQ+GM8ubctNcG83eusZsrYuZcjxy8Cl+ZvysTIJgaWEga0
RuNlV0yQhxA1ZAE+i959U4WuK8yuo/uKaM8FrEYb16qw9i/VVgvbYuJlfkn/xzqA
8LfF5Dlvueb7tCbkBtRWS7YvHvHik6YPfGvlbBlTaa9Ndne7Dpx2klr6un6qYu0r
O/ZBlmN0jPygbfkWM/+Y8uj8Uu0Lucy5CZYXlRRwV8uCHhcKSYPwPbYFJqh553Vv
qW7+DfON6z2FdDhrQVIaR42idB8J4A0lkjZABzhglW5iOPJOAWCCCVW4j+m5CEgK
42JNPnfIw2Q2OMeF4xIIKh+kSVVBkXNKNVzgccAW4tdrjyMI0fHesG4n5Y0YpWxE
jXm6B+IN9i7mxarPv99JPUEJr+C6o2TKFGgB3cFUHSja7H08rr1YXtT8b8mkFprB
LB6funoJA4n2J5zB+8s1javXEyPojoJfpQKi+Hw630/Le2eSW8dgfP66bj0QFYJb
mjsQ1lHUjWbxaL4vH9bcm3WBbrK0wmqNs+weW/X2Hhpe3AcAXB9NCKoiin6tvCL7
ZcOwwj1NNqytAxjxsb1Q+uCC/Vgy4mjcY+7ERYU+uwDHysJigljD/vyrb+SBlMS2
aLV6R/Q4QXlamuIV7UZyAlCfuUvOkuzPqeqfS5i8XpqhxASCZ5jkj3MC1xGj28gC
cEvyDLWdGQ1dHwqE4HCq7Rm+lVj4HmXqM/fbfUH/iWkhmM1bltwMmUzLiCIhp+jK
stxErRJESoy2wTpdcuenh6CbOUpVabEitxlxNJABRvHOewCY+VLUaoEmz0tCOtwt
4MQf+a8ds5pWqCj+2Z+jixEcjY3vpdQKtvMGSzwsYJtTWZe7jbmKrI0ZnpTGWUEs
+P2RQ/3rPh4KBifPbZQGVKHblzDKsy1Fub+o0R6gfOkRI+X7vi66n0KPsfKpfGtK
Q9jb0WG+U+WcvoL9eEJVA4bB2QJuc/J/XZCfhpfKdN37iC0wODKowdeTGk/MkKOu
ASLd6uchpsm+DuF+S+rmRoFwQkCKRjzc6GEJXN2zw1FVWvF8epQt58X+8AtAWmhU
LL3Lvt0bdJg7YsexUTi5dQJuXnrqR9hx35hn7BleB6m35KyVmPoFkPBpjkU6MBgo
DZDCc/Z8rXITrUfmCtwa+xjMW7snofnUa4rswHyovpf7L92cPqZ2AFAJcPrK1SKs
xwbNZDZIDoqecw6xaDW/aFvICvgQ8ATWoEPiUh+78TUqYp2Qtqg70ZsNFjdZzVc4
Q/9uRaJFhimKkr8wSPpKktutbkpF4Jy+QXflod+tTuZjMdUgB1l93bhG2rF5f/1i
OoYhmBw4oT8sdowJyBVl2VAbjME+0YYyafZrxt8MweCQxhn30nx8O0nfHt0gReI5
8KXXheszC6raHej7G/tnFVO9WYL+cpYq9ypbcCdh4eXPenb33563EoH/jfLihwaG
ETskgpFYrQCvEmEaQ+XYliHQidueYq9BaV5/x5omLxOGqx5RPZh7a/hANf0FJ/Jx
OMNIyng6PINV50fj/x5PM7uhUN4j9FQzlZWw+dqeN2VNVSmJx9O0Z+q6wQE0ifAc
d8Twax/lL8hV9Zp8f5eyC4I8webDE1hQwpJeFHpoHgW0jKOmIanUPdG+2K2uc5WH
08BbpGNs3yOQsWtiU5y2RtAyWQ1tOIbIZF4b8EZjjs/zpo4FprRTM/FQ/k67c0Bh
aumUWOJlEk+WEzOG/CBNKfVhQom20mDKEOiwGtH/hoQZ8M8866lIS45dDDSNCgtn
OxPkiTK7Ad14GG8+LnX1fPt/XI/oeUx0x4soTKifg+8oiZiMyohqY6G7xXfnNdp/
zSFdH1ZP9Ch5Ik+9hd/jiThVov4DEw2t5do1kBtw5VDZ3Yvpmos3QKRqrjzfp880
wJ/eLchNpVR++Ld346Syd6MplFPrcVbOA5tGNpbEXDwHLTAwww8C169eSbK9eC2V
3voSGA/TwiQwy8fgTULxD72quRvSJZFbB2j8MI2t8LIpKUUrl9MmlkhDDH6JE2X7
rYWgVGaoguKMsf4n/8wAMfy1RA57KC1FHp9teDibLLfD3waJPSume0x68x66Dept
cfLlyrejtGO02Xik5O3e/pQUi4oH/OYA9LgPKnIf7N5M9pOpIvPKA49pqzEsrP1H
wVGYu2U79ha/hF1CfEVn9Q4pHvMSzh5HDFsbc5Q3V3uTXmGvo64hIPNz2AKgplXS
xQO8VzeiGMlYA5PE5+tELCHxkglelSAIy+dJrL4RHnqkyVT/AX9sE61hsgMSlHwK
J7bWWcxqKhH+U2b4cZoXnzyZoZLF2yWjSBTMRSrc5d/cdzOeKgIMM1qUZ2RK85XB
tUMd8A7R/DRfspy62x872MBjSELSikYmkZsfRTiPRRSUDbxNEX37aIMBtH1LZWaa
FUW17yhZo8mPaUTxHchRrEjrmtLRKcWSBmlxF8PhOttdnpReEsvAkdMEYEnS06lD
Z4i2uFC/QoZILwjN54j2PxBGRtw/ymWAkLZ8malFlAawMiySJRmk1crV5pnkmI5N
P5KLhLMJZoD3jhSRZ8pCe0LEwWPt2Y8FgL6B74lC/YznGMoUMRcFo89jxYT82a4P
iBKwWR0aDJy+sizXuNtsELk/ui4NJ4oAR3SNhUNz5m7iFulvU+DcvfWG7omLJ1rQ
qDCyDcXgkcYwpRc0nZOYdoIMzB090ZHoQ7OPkvpfQ0aH0ExA1Z3KczD6xQ8dbZZK
0N7BOtqWqFdOGUElLpaAsZrEjH0yyXTw8JYd9BHAYpIYiieIiN3uUKoX4S7l5DlG
/EdDOE1stuuWBHKhZpwiMoeBg4JpgDiLCcXihwSTV+XqP8sj0IMyduqOq0b9Qalz
YOHOi7xp8dVB0tciPT69YhPcGtwQhGmvM7q8xY50+x3GTeU5dHpAJXfeDlJZzvm+
EB0LOdfdv377g2eJOSnOg7XyNNLZBPVWEoFLjzquQSkwUw0Nh+6f5yahRaUb7UAD
8l4jl6qSsjreJGrwJC2jNElF93uposEZ9Ahdo4Up/UgI4xXgzXLCdvM5jkziE0rk
83Qn2QF9lqao+4DB7+JH5gGAa/hmQWzuLXcW9+HyGjTwnPouUpkN3BQl0oI6UV4J
ItolT6Hd4+F6qUWvIKEdF8GI8OXTTnvJOIceRYCr2gAlaLqqbwQ54hH/DCfNABJf
KdKhtTv5BJjhO/zBzqgXbjceQXWaGmlojcmywn20/2Up+BMUDz1WWOZd00rxrBgn
WlrNTxv1TBnR2sVjb5R4pw5cGsGsUEKj2DAIc2mKGSQzglTqTdb7e3pPCQWN0zrp
jh1LbmRHUwCG7T7dCApJTJqw41YqglyA7lCvdhKRMK8uAwFZLavGeQBr4MbwThE8
xis0HCTi6fSroQsrNvaOhECZiHICUT98L/XHBmj5HGQl473ye4m7TzcN3cKD4xZg
UhbwZBPwvCXz8R2TIHLSdUfZTOZto3oe9pBRf3YUbzPt0pZ0cilwx4TZTbaiSLu7
vGbrIVOpD6XWwP2+ksy0w+zU5ivcZun+dFRZJcgtzb1Q2WHwKLNLNtJrsRJUvIrY
LZag9oTJ2eCLOpUEk7zYIcXBgWQTBZ5S7uoAwbfAmRsvVfyoOfFmcdEU31QJHJ0+
GLSlBLYDrn6JbZBaQW347ORD6xiKDiNGRlcUqnfltuvknbxo0FBa1bWGmCyZcAUB
RWeaqYdWAVJTpfEs1Lsd9nwvS/nPHoBulyFoeEIapGoL6Kn1q7p21GFr3aN086Ri
GU7uFJXvpSwG+LUiEaRYPooFfet3YVgiQxHmV0xMvM23JGGB+gncw1OzODo3vkQm
1Gn3b+LpTwzCBb1jLcjI+dRM61vRHRFYXk9HPG9vvvGhiiia7LMY/HExEAjmcZZb
th650rJ2mR6n4u8NaXYtwo51gadUWSlKf4C+wH/Yny0gJ54GTLs+a3lUg5ULlwuH
UkersuDlv/jCQCkb6uNtJtXQk0+h3GCa1BZEewXax5qpQJnCmTT7+6g7gjO3MTrF
PRIxFdf0TIX5dXgKylGWU4aEyOKKdX1YrtkwwvIAIOZ5zExEmq8ZP5c9CBBUaTu2
xHta/lEIIk9SAXLszH1gSBpkIN9D2XW3fDCCu53zju5gfh82kaWTh+8IY1/mLqZM
red5RkrWX13xU9rs4VkZgb1eHU1BoVhyBrWv8kt1nz3BI7e/qq78hF3PBUfaWD18
d9luE7oBOFAo6Z4R661gKC1hkCn6ErGzAJQH11p7Qmt+pjCn0vAOpExE1kBh5rAM
rgWuEyS+5xxN1fAFN8cblp0gbo+6PsY26PmZpM3PkdbWv9SZgpHb+1CGIQtlWRhX
zjxFodGAAYJnllRckTFBlKBeCsIJB2wurdqRHn2mi128rR4T7YXLq0kS77oh4bhN
sOvOHwUkv2BGaabPqgVEbGBPyFG6tpyeN/y7F3uBuNC87kmNM6pGlctc9W653nPD
UdZjT+JQowGoNmxvvZQumbft0qpRSGdjHZaMUcbcWJTqUA7Mx+/Jj9n5GA1n75Mv
T5sMfDsp3uaAU8pyQeEAWOj+jCsjNPNRTbu9HBk9x5eHT3crcu4rncxhL/JjxpyM
Oj5nf7JGqqbkzpwTJEPoQM2ZIRr9g2HqZOVNwK8DlQUq02XSl7JVdA1LZ9sEAjAu
qSJ5q1byDUDtSrRyzEx44dc9C1Lwy9ZyUJanjFTQspvLMaCHIu7WJmlUafwGT/z1
aGvXmdCLg21373xWMbutb+4S3T9exUyL49aBBqd7ufiTE1Qxnc3L+FIDzNjR0UR9
cV5fFgHjEb06bBqpGDZnlkthJrzcnabCEHuwt0i9fmu4pK/fipVt5zYJBYwmCLIO
en2GZYT7lslBM6n8i1kGnwJbMpKkKfmM1gGmh3boVxF6jxkbu0HEqXLH22xWvHdV
uviM2i7CROJnYqt6fDSL9sty1K55Asp37YGkwm61c21E087bq7MvhkiT1pDJtcHK
u593ytYW3E9mQLiGWOLxcBwfAwrTRVQN4vesllAXqLlk1XfhyQykyIIEYSrZdQDr
rbzhJY/z/j13jk4JE2uRD9D2aKaZgoUQM4XLsK7jUdAyMWwTE+lvmW1upCIFMybR
FHTVPtkeQmOLtcV7+M1hPrMRqfEIpH1rUI7T4pGmmsaqU0HBFCeUn1io8KQWwo5F
NhblQ8Z2bPAl7OBEpXM1MaJD5xhTDd4WnR/tp8CEkeupj/oAVMtdH/fNlDj5oFpJ
Pmgl4MXG/OA49v1mGRi9xCdMdW31Yt2C/IVw99lOv8+HoZvIGWMN2XwKkYXphcil
QXZD+U+UDlj1LDohSkdTbYqq9w/EebC2jocmHHDvFXakhXas4QR0XWzWnGw7PwaN
WOKdqgkxpILLgakffd/ewwGyitjZ6e1AWz4aohJzdCmaX3ABkSqkjXe8fR961Hvb
80gaI0eHCOZsZwHZBOFhDpzsNfkyH8zxoB4mpm+9J4baTXSr/d/o8bpDEQal48AQ
khts03fFOBpNwVi/JcpJ561R3TboRm5fxStxYoGBLsg2W8a8AhYwQFMeshmYngA2
QUIUk3B2PjWY06sRdnIOGjVr6zqNLRDsQdaVxdN0SYzrHAMy0bk1CoVGXrf1KBsj
jhx3U4qNR95Yh46htcgGERWv1lRhzmL2atG9ZdiWP2cnH6RH9MsYiU/tX/675HJx
gvCAJDKxugoOVG+gMU+OYTeu2JhI1Y5p8B7xAQZh/ZwdWhfg+bKjjJ6dMI1Zwp+Y
XajOdz2YFGnpXyfmgLcPmz2ACKRXIMvZpLWW22BsgeedXZ1xI1lr0S6pizZ1fTZC
WxyEHfCVh69jUtym2TAXc8srSfdkB2RpO2ZSEKbbldyrYS6xMs+ARHkxqEGt7QNZ
49eCy5eyiGI0jKaLtn4sDO/jsge3nKRjmDFZ+i3iUpybF5RicGK62q8ZHbiNzijG
v0TDmdl1qYrZRQ/jLJZzT7d2WvJbDbGWnlBqltht/8+2/UHNgtAsKFwGPpO1WpBS
2eq2biYopTnXCTru68FSIjayHtUaHoQWWKL/luDqqxT1kdTUxPK3GZBRo2UW2qh9
rtIeTQTLbb9FDKx26YoSBUjKE0fVVLuwiSEBhMP9mKCP8XPZ9Es3d/Ggc1al8xEN
VP/mI0+m65VP6cbrJwPcM9WcHQb1ylDaYm7omSB1wRt7POZokYYytPqFFJ/UnCmP
0PahzRQgtP5El9EszDEYsxnfmSGp286ydfyQae3XUoKQ5jVbpBkxWYr9Ikq0vWV/
uwrLxr0PW5piiosVJdcSxoZzIkEZ1t8ecQP02Yxqr4BYzX0q2HimJeiw2Pp/bXKr
xAbrOWdP22tSc/rfp1qn/mPp6QlHtyjwPdGslKbEYuZ5kZ/iX9irnAG24C5+FR4N
a4NE8lRTK6aykfj9MQkQfWa8wBokZ4aa7CE8pRd100oIExbrGZNKCXGZFPmFldBr
KM0yZDOardJQJJQFv9awT0KWvWfxnFz8zpHhVgXBxOVRWXIO/uS9ZioNTHL3MmA1
jQPszc3QK5OIc0zLQrnDUsDd8i/R7GMjMyrGOKrk6d/3NHpSou8QNOIBOmYE7aCX
e16qE3KbL0OoLcGNAoyI1Xll6NyHC4Z7mswRiJdu03BfJkewnempWMymKTVqjcTc
i5STenIiRKGVWr33yTP/B2aFiVKjrFF2ZJ+Rj+i+ANguW3SfOSDG5uvc+NFPI5lt
QpdfJIaXTtYg3syIR6Kn7qS0zGu3nM77+2s2wuR3UCzOqVYot6sAo1x52K2ZiK/0
tViTWtYR7iadKlJ2elMgZvII6U5hC+Mfph5km+S1dA6DsfRximbzV8UBq4BTwNYz
ySZeYVLp7YHQIzaVto4RqqFCJnxlTO2WXlvrmHP6XFzO8UoedA1d+uEIE5OIQAyr
/sPc0SWsfgtguCE4bROrmi6+LPT/1996aEGdGVqZ7xhPh0afdiFBh7yU0VnX5EaY
Zw5chBdf/SeMt5LWCiV1Kuiv01v6YCx5ofUFaiVV6dvs4et0PQKoZiMnAtp4/vxV
yDjjRs8td1tRV9KpKhowB0SBu4q5yOeeUmPP95xyvnVNOR0PYSlZ1O+Jv5YV7lOZ
SiNEtJEujrPTCwHDTrhTWB8HYeYLLZVbmm/ePiiADLNHRhsriQZZmN2EO2sCUD9T
0eEOimW54MJAmdGDxNRJHNvqRL0rga+YrgTiG5OP/wBRqmw/3prKiqSoGoaGPVNy
fkcN3igHC8T72UkkYpFk0s72aEb7OOfr97Z8f89rG4pFf6CMAhDQvtKxXYXaA3Dn
hYVHNUQyW1UCxc4OYdbSPR116wiXMhJN1Til3cjd/TTQjF8dwO+ZLu2F8b8L3api
W1caIatc/LDfHrlvpi1kdhVc1irx4jdhHVsHAMWMvlmw4C1ivvWogceG7rpVlPXm
7B0Xl4Ke+I3rNy4XZoG41jOBnlLinK2pldn4v1hSPWzI7bxOAC2VBRqqLJMQzims
JoBgcgVWErAMPTjxDLeu5UF7PYEPR/33qIhc/+VWrObwZEswVHKIE8Y8lfJjT5Ih
QnjMbOp5s/hkXBu7Zbf11uVumZapWBu39s3QDmsYCzBLX+pxhmV26+8R4ZMg/j5u
wTXif0n60qsV6MHIBjTeZHkhBEZ2ImvPov7XV3cPdr2ZQpH0PkHS0VJEr7A96fm5
nwPiZd/eVCBZcpVRZkuFFD8yq9nSfU96En0KFPLOk3K3xh9SKBcXjOGqo9XaPgp+
6V/xei9AyhtfrGP1lC4mT8cpFnGX3M28zBVd1NGobZHqYkuURX0PQwP2soQSV+lV
ru4SkGLxbZs41mDok8k8kCfSgIlOg82yIA/TFieYlVeBQ+cyzXPYabZUkz54TjEB
xcLpA9UpPGmS6RYKAdColvc3Cc1s9SzaQAE5VyP/u5h9bzAEZfsw00kDYEo3xpf8
s+OQBez7o2RL0AD4A9YdL591ykUME+if3hy4YLeJ0YZtYkh/dGKS/HFjdtxoyp43
+YY1fyLORMrHZsZQpjz02CPjYetXbZ9Tx0rBuKMaVl8zlL8obJ6PXIThbabifwx5
5tNjNONG1u9NBIsaJV52b9McH/Cur9CMdkpVnbmJDgpQQhVFWYzI2APQJe5wq/VD
jnVk/441KfCg/KFhcGJ0Lz/w7PBSeHICxBAEJOsfIkNMVB2YBDhVu7OWysmTtnXs
n3jMcwvMcGzsscCOzNj0uLdODwV1RfI8spYgGUz64gW6HumEujvIMAIAZA3qVXc1
MOFB2T0sXQOs9YYFdT7c37ZYJlftEliFBe2K7XrfrZYAjbtSzowRtubExRP7Oz76
nnarGZM0ho4uzByswqHi1Jwuk1P5vraUtrW+iKaFsjXTuEzjCnLDd6m9EcbRIJPw
T220FbTH56i8rXBwk3ApvGEV1GnP9HYjabVx+Ac9LLy41HAJt1uU7iMsq4Mn8Jzo
g6cwPbC8d711redQwfNQxgoZfdou5jrWGsIsU4s9a5+Z1s9crX4XoKaIAmliA/qx
Ol5XRaFEZ1VyYJHoozczjmZ2tTFS7wlDu+qHefXj3ANaqDC+U5xNy0BjOuKR/zpQ
MyV+rEjAVHMLi3FE0ZCBM4r7tc62wTiOUADfLQi48PPWSW1CSxP+n2UM/Sh3SKGc
BjCtTJgxgggU1G2lKptwj3SMWE9Xce5dnxrjEDDNr7SsBM+m3MDI8EtDQ5VEKKMr
t82+7WrIsfCp2ZAxsxzj88Y+X3RkYVB4NgDmtchC9XruLCn3CSEdrfGO+e04p5Dz
dBDk5Dy6CA2IrzQ+k9p5U18IpJVPkjPffC9zQtdIZ8fAcdwNBFHcYp7vGZZ/4SmX
uBKHBThYaCfXznlmvWagk4QmPNNIfkicyBGbBtj6TIh7IGANHq/IMF8geSmh83YL
+mVvib0MDs0OfOqILwUoxUoWj9zk35zM58A9LunapX+xyKzrnlsUVa7cdps8ZeQB
tbPl8Lja5VtAQskS1lU8ATMgdFJaXGhrMl6TL3l7AD6/uGEXhM3xvIdVGKFZK/JT
n5+UiL2kEdmR9Vf9xPEuX3g+W78WRspTsKs8d8vNaAGhbyo4n96tQWK7dC+6NcUo
DLUJ5Mwq8wp8tSi325nCAw9RKaqvqBTV1oBZvHeJnBs7ra2ovsMq2I5qupWdt33C
VRdefF05kPlzqNr4x2+au5zUeDUixkLrVgJ8UQqeKn6h4n5wI4ZORLJEaKMyUrZb
QQpDxYH4qisImUVqnu8C1ff8KBVuHpQrI2H+AnRJCrrXGVLCKG8TYbzydejC9zNe
EyFTdJjCNQjPF9dfzizNBo9X+X/dYsGhi74+7B0JwW+4wWKgZwUw69KBZCOtO1ws
zxjDMKw3QQgq0UyKSjvk0bdlet7RvlCxzBnnhbNpENi33ZuAbzaK4ndrHiIDRJcD
2EVuSE00CVmV9b7BP05tG0GzSBO5QPtIo2ffyRn+E4mV4AzKp1XeQlUctHqVnBC3
mVwE9RaH4EDDJbKw9nQMYRsx7Xi4KTmFnkizzXrf/e0EctZxElb7u5MqPcF5K8Hv
V5nRlrxP9HQOMmK4UpUdbFZFW0eO3dIoRfbe5Vviucxw5dVSH8TVAA+Kr5U6/pSY
2HkD71UFNBWRzYF/u1pqXkfyW45An129T7j2HmkKBKo58zauRnLlFxY/JiFO7A4i
yVXhjhtOh46vK7lx2/8hOOgbxdl+GP11quBu5tNhUVITOoJOqg1gazq7RdFLdpP3
m+IK/rD6S7mn69PmlDFWalafYMVYCi7kRA12mSxknKFHd+mk0zYqSkhmiBykKIyb
mGiRdeMWnm5ZOx2PjWMxP4lbE6IeW+b+/p9h19S1x4/Y1WO1MQSgyaPWMJ5LQw2Y
Sm39p8JQgs+MnabOixDaaLRdrif9sE9MmtrXF2c/fu/q3iuUI2ZylT4J4hQ6pBmO
9AiQVK50aJ9jyAru3kNbx53Z2zlGGnNHjaLruuvYtDzgDYBk/751f43ZGLNqFcHb
lM/Y5afd49GENesSOe8433gR46+17VECIF3ru0+afFmNbeJD1lSFzGvvn7LyRikg
PLQ2VnI5x/XW4ljVQmfii5wMrO/hAvWFHPp8Iz/UAuD9mg8jXGAtV6MsDjr+pHei
91Gx4+8Xf9EsYW8tQQnGJce3MdTMt2QD00auzr2KAnh2/DNtkZ3qn6q3rBo4RNQ8
8rCRaw76+CG73FeCF1ng07aUkDjwziTa9au6izEyo94bROS+YchmlVXvrrlXpXY7
NRtmBKVWgDpqg79bft3DEry0miStVXkYk6A2ydH442cAz3DP/7TQ5OSxCLBnbk3J
weYM0aYVP9kafn0aJTJ8NyyVzxsxNJ6X7eQg9K5MpHRg9VVNgRq/WbWX+DZl1F9K
KABYOg4Z3xBaeOe1/0h4Cb3NhIH1fBFiJ06NV1Fv6jSDGB4lw1/4uplPTS4MmqX9
baUWo2DtZ9c0IEn0D274W5WXNFHmw9I62I7GE/oAt921xgFhiLGXkhBWHayc96KR
oxEJgV2vw7S19JE6LLGv1BmQmsGtGsUNnRKKkCupq/jn4u7MG+nnjle30CFmPBTG
0Wl+knRSWJFxF1Fr7BgagFIt4BHR3M4aSDm0vqDPJmCDEULy61Zm2Gk5SXsRtxyx
1PeXPGMrNDc/O1G8OyTAR83kYrYrny9nZlg6NPlz5JYhGmmuXGcNqqlkDRjHwBLn
RXRIXlxU9itPXLrCi6s7Zt+FMu26Nvfg3HAooh5xZMzAE7ZkBQ4DBVu80n2O2Hft
Ti9o/mDayQc+pcIkYWmNXQkNoZWtpzt0+dIGE02XQ5h/L3i34vtQ7Z88CX+uo2HA
bhbyouNA++XLOpdjSAlfvLdLdfVQT6VP10XAxS7iJwGuLYnmqxi4iJVBmm+8pLvb
glt3+t3OvgEhC8IoO1ZA+f6bsClbGEY5frC5++TEQ2B0PQuioj9AVb6pMc5UpF1K
Az7xCEkfIVGRFdgF3RMDM2s1dhlBULANTccjqEO9q6U4xbtxSypWQo4gSOhOuMC6
4mo6119M8oYZCPPEPgkvS4yJN4zqoIryvUP7IC37ky7z4mbgA8bTOsSdfinTJyCl
cPNriMFcwxMUDZ6ay+mRlU5DqrS7X4MSFDkGu5ydorPdiKyyWfRNK9xY+j3MPwBy
JMA1AjUDX5ToMjoGcyInm9jOgmG2nXsv0WSjHbOwxhmj5Sq60w138pX/zTJFirtN
bj3mqHoH6MU/EvWgmEtUld4gyyHbIP4suScDsEZkAEiL21bKLR9iotBfh9mQb+RU
rHUDUsBGEb6kk3tguUAFgGYdOzOvemilw3Qgx3AytkeokV+FR1stkH/oV2uUX0Ag
oClZZwnon5zg0zYFooUyIN4oKfyGTkwyGdu8Lxgw4CIfIC6xEziSX/77FDRO3Ig9
k8rVlTL6xGuDbq2g7nKaKLUcuYFJEDmb1G96jGWBHnszDUjO+QXJyL0Qg8dgdk8s
6HM8AnAtnbh44gp9+HvGdn/lBHBVocXGOCsksPctu+GQxFepQY8fRIthfA7NAroI
QitbrQN3ajsuXeYe5CmNy8KqN3hdbZVXMw4dcsuYDqFJmGTPPOwFYiKsL7Zt47nI
E5HDIH1eTGMXabbET6xAnM8gYvOPfipq5v6nksoHNnm2/xh55YP7NhpLZOJKbVMI
T6CGu8tnNgJW1WWiN/g58zIs2uj14cZYm5+7iUxNqgTNc1kDz6MgjcghUHrtb2ka
xTZkKiL48gqz3fF4wSqZQfJysnDyr3oQg2EeTqWJoYjlHOZCFG6/hk7xIARW/+rC
C/1iXBwvL7IyEO7GXZagO4+fmB2VDVCi6YSU0f64P0YvPMTLDIpeILiZrnBU+rBA
8rbjSuMocgPKWnDiz5dCu0TWXkY9Br0fA07rC6QmJWhoa6bdIxo5Yx3327nL+YNr
r58BnWYWL/uhrNFXiDgR7lnShRU/zMMSoZCeNsffXQVveZketT2eKL/2AwoWiN3e
z0r7xmPkvgmC5/c2Hnc2eWv86dg1sG/tBh650mboXh5LnHktKlLhUQEYhBkg8bvi
G6Q82w8StpvSl+PtLynRcKxETkOfnEKlkR/MMIJ3yijj2SZLv94vnAOBP7fGAUO5
FN3cHgc+Bz7/Vbg5H+cAsLO0Oe5YBKe9CsHGfDV1CbB5oGPNuN7S/gydti8Z0cKk
cotk4CvvGniwgL5VQ54oFJMUzTuzJQlreDYgPvCqWzZEVj9s9v4cb1kg3Ism/+M/
Skngl0svJl7sKM4sNJhHTfzP7MLHn03DHynF9s03a4Y212YmPPG7be87TQRw/ewt
vnokRKsyVu1W+dqfGjBj2oTdTM9JJJBQwWPr+2+wTtKBqPQYUFNLONZruehWhLrj
fXB4QWgamzw2nn50oFYXlgXRJaQBOPw8dhDYQqw6Y9CirObZAL85mDYaMkJYjPc+
S3QMHhdGa1vt4vQ3nX02vsT2/Q6XY1W6bclUVO389ERAm57g1xJYSeWG1woe7NsN
tftOQdujbIbTdwLbDlgfVdl88vSxB+ncXSIbdWskgm+I/xtBXxASQUHMpjaDE/iX
Hf0OOGG+G22zWvKxnHMIYedBhHf25h08b5cH5iQuzIE+Qd0rKuETrQAkcJbhUnPR
PsVlfN9YcxpHlO92uB5sPuouMloaPtPStpLgjgi85Gd2hl1XqL7VgX88SfXDGFRw
8E3IicfalaJycXNUN3auaHwsNCHsQU00GtwtrM9eO6VB4WRuIhRNZL1KPU51uFkH
jMU4loqaONtPWbKtPsoJq6v9R0OIU6DQZaCui0w61oOHJopxjceCOhMWfbp3bflU
SX7WtLQy0hcYkLeEDpIkdsOxoezlwDarQ4/hSy+1WjgEP8jBwiEWqwiI2tSbVgYW
LfYXUT+/OsPu39t/4JhJb+kkk5X5ZwmhSvHfpbdllg2+r+rXGoRjkKn1OtXXRHYP
1aBqA/4RLA6HOxr3XvGWN8HJb9+Lqo5KCwObBQfycxn2Xxff6NwZysAlIFu4debo
gQxfEZ6+nO437y+3Ow31P9v6jFvIIk2UrIBuVl9IWoYP1e6w4pXhhNXTq+x9d3fk
q6beYmox0Ie9ELEKI3Ol4rvmGesn2oaNEagYL7E9+OZQKA/j0VS4K4r9KrQQQB+z
lXqSiCEfGrsaPyp8LddAWmZJ0ejWxy2Ceasoried0gXE+VDDWRvOiUutKbjcjz+w
3OIBNhsy5s0+0yI9nzDegW/q/aII+G4hVd7yTs62U2G7wzhwJrE5Ma0gLYtdBk0V
1Lh56di6H2XBQ281WZgECAvEQEgrWsK7KxsDLLCOjk/8qx2zN7J/4sY8ACau7fnx
nqmzXnYOEDMN1cxtmV2tMcLVI/EO6Z6aXsU4IwQX5xJXTcDoKQp58JdzuwIaD2RV
n4Lhs++xuP5VEMgkwZ2sfxXPm5f5gE1XH/ssrCuzeEJKNwDtiqDEJ8ea5/fU3Bhx
4KU+uplsSX+0UyBzL0oMb+R8+4ILT4B4tzrnuY/uoz5qR3njUp00C+sOkUPy2rpA
nXOnHYwGvP11cFzSbabcQVLeUDlBdLhTkFkYLWIZIB6jDclRIQ527qcPjdkPJfp4
b6qdy2D0HE5tltlresxnETF1Mda3On0ogyHEVghGvY4mbV+9I/W1MB0VnfxMLg84
wzQjTL+zTfYDNm0tzp7tlxwfYFCHD27cQGQjRLq5I61BwaV1U5h4u3558jj8pO1l
mQ9BLO0YjdvB5YZZf9xES0QnyxLsHUw5N22AveOGX3YuaLXH/UJv4W4ElY5AQjVS
e59kU8+51MHAUJ8e6ljk7tqnLfWe+HZMUlhLOgZzSo3P+8cfJ4h12rMgunCzAtem
Bl0v53gXpPEqsADEXvwddAVaMK+t7sihhUFNNMBRS619enf0ifg/v6cvuAZ4qkDy
Lb7GOkcz7PMIPs9ulZd10Z5sslqgZp1m7DIdH7RavrDUs9uRIAaYugHRxFXE4tPO
SBiR3NbT3xMuTAdvHYw0iKqD+yL7FBjqfGRn8janSpVsiQ9xcSaiqiDXRQWQ7hpx
KiNE1+0CUdSEPGElvapKkmsaa63Fv7RDLC0vt3Y2Zv96ZpLrHXs8qpBU4jsKcgmN
oU40GS5LVND7cvcmYq4ZHja2KucGmCdfvVMq3KPun6LgoLToRNz8s3tatVDu4Pzv
iiETBeGn7Czxf82OiRf3tVvRDCU3LFVDJ4u+vjPomSX1ADpqNxWU4t3G6yiiWOxn
SmnFwdr2F2PAq7QCF+pDHUBHBHOcf4tPW1nzxCf6HB7A35rqGrAv5xyS/aGIfQJ9
2Dh+tB3WU7URSbTTa067YsAeuEpS5rsA1D1DU7NOtV8Gsn6keKILO7tDd1uT/6BJ
X+zPQOwGhdnCL9+gOWtZIeXEIhGH0yfK0i1UyHxao6h8qnQUFBECYR0gw0JfLRld
X/IgaRalGMo1i3Xz3wpPb8wI4qsjdTc0G3J4xA2J4sa7sc2xhi0dSeRCFJAkoud9
cdzwoSbcFsdSJ/CH+SOwqRekuLANfWrwzMjg42psGGY7e0xaN4MOQS7xAsrYzm0N
gmEHnk3gZdVamsekizHRb2CnJQqcatgDlGfp4sl58b/GdnfuOtsIjLggfhfUdSe2
jZJ+dX2Pp9BAsY76gtxDcFz/4k4+6ZtLlUqVONgCPwdNeCwK/H1hSy/DvYoTqZop
FisA6OdChkuEJBKXVulgNgI9GWiGHT0lFN8cgQ9cVgdE/0sMBB6raarQJ2Jd4W6c
FYBeuHSbHUTw2wHIOMdIqWOQdK/hOZOvL9qSq7j+xR/iFZGKlPJgwG4rFM753EFw
H72zXCK4fp5DC7R4J2hGU16u8ILAz3x/3WkJllgcq/W3RRQdUa6E1F0l2J5H/qKq
L+mYP1J9BvKPpUlrLOiCdb+hEl827hJFEGC0gh67dXNDK9SEu7BDmIgYAhVd7ONt
iFTSYDOV74dR1j13kuZGuCSTkP1AV5G6RodaPAod8uYPScuobKtDEQFbudNH3za1
wnDIlzpJQMPbc9hOCyugJSGqmNelrUL72V5pfr15NKptNG06gNmhOQTG1cUcIP7D
F1ePHpr5Mf3gpTfS/Zz6FXag2xNF0e3fuDmbiVQmm2AZuxtTyYIBge0bmPNvDHT3
5dQDYDe3/Cv5OOcekWw4+TQejf6aRUm1QkaCNhL62FJIteLioswxGcaYq4bOZGgm
mquGdr3Y6v6Xxi8b8rV72GhmGj00/ch4uq6pRhNxBEZOL5mGrgIFrWYOqUSFIYvD
wQAj6ugStTK0oEiS0e3mX+Fup6/hxEV7Cf1ShNQq7ucFYiXh7uys/NfHykn0QGYJ
qceTVCV3SGkS6fNDZHm27icBsrazdU8/V+WHs6WtN1jujoZx3u2C7TbzyfeRez5b
FzNBaDmBc4Z4iPrYZqmVKIHi7Je4dS1kwR498r7e03oes/M4ZcH+m9Vl2YBJJpZH
STtOoD1roNY0z3s6TEAo46VV7BHdrbJ8u9SaqH3MbR+H/7KWkY/XjEwXMRfJEWQ+
+oLJc6oePHqHLWPAj6TRori1Q8NYJDgCMsDNY2piWAVSDJTk5XgSOgwukZydF+A+
faKs1rhvi9fbo1YNIeF2EYmF2KsPk8stIa64gYS2L/8zcmAPbLk/8ASEn2iTY08U
oyaaBU9rq+xQ0rmnh8HDlWdg7+j4mJw+FdiJO13HLCCQf6Z2O7P1S0G0BB9LMCZ1
nJU4ICC0EZs6Jsp2Fi+ha3VMkEJSC/Y3Ut6nLERjfMENHBPC4wMi/md80amwlWx0
dUretxYzrzdFO3yIeZemVt9HSRxaeN+2jKCnsaopERb4ORGQQruwZrIzo0maXU/m
P1n0GX5gsnjuq2QPza6hQlQ7+Qwfv1RlkgRxPto5oThzv8oGnpbJHjkuxc4P0dqu
dyXiy4s8B6WirotCmzL1/JI8pGzSxOFHyVr3EvsuPHETD+FD5fGBdZrZyQjt+JB3
w2naefZ1enU+E6CUlE1P5V4qjgrF+GbAFkb/ryrEwAGmG5R89/od0Gqx3I8Ity+R
0FUgiLP7DUfpmmI0Gub4lCnLeaGKSh67AOi443Mj2TFQOn/Lb50vFIDeg3jGtU05
zYqjtCUGgVwpabKwRjNFjophPwQtv/f8fnGPi9wTTECEQfFjpbbTfg4cIqcY1itl
uFGAw2lUoORYsJl+Wf8SPCduq9cPBkFpuVWv8VvrF5FZWDGi/9hJjWUMw+sBHI4V
4J5/0kPbiOlO+bx5HS58Mbbijczg+aMeLQhesJc3h8wjwZbC98jK0j0Uvs5NwAyj
dWOCcx2Dvvqhew2666luZBQQAxfgdFeW9Jxc2mNX7+z8f5WG2hMOIVY1VTeBml4b
4DRD0/v5BxamqneR4aExayC3VVr029GvCqmB8jOTiJqVvKiSE/c1feMZpEaGA3Mv
74OF7Pg8pr6qJOSeSNZtj8drUzvL7IcOEDYJX1S8oOXgUTBn5QHeC4agfQUca11r
i2ekH45tzXI4w8W/Fs3iP5oycyarkkyryoF8UFClD8zSho1/uADCzo8R9NgcfhsK
3SMnCwVFz5M1avPnfN9TD3dIfWBlus/76jxHHm+I03x1yIL93kjqRYkbx4j2xsGW
MOSvIbtbTkzFa+bC9HpjbtKjQR0AdWr+jVhvdFAM/m3PNKL6h09rkTSMP2b8xgxE
/rI4at64hhbYgjB2+R9FfwahWwtqSNWAYvSscu9IxlPSfcgdzYdH4HNYFD84sriP
l6O5FlP/lwMCTQJa0WWRyPJeT65ATTAaq0J9FqMtayuTMErAte2X0DskRaHHrONW
qTxz9zDnj84r9tEU4Mb4gNmBTIiG4gOBvqaW1wE8nj+PrT2Hq9DJzLC3vs7Tdir+
oYEwduzinkXhwBAQSpgV64jtOjlaVpuFJR8yQb6cHBzh1czxOKroDPfMdh3Q9C5Z
83TRcHHDSUuH23iC1jh3YoCtGaEo7RF47Uo8O1b6ehYVaPXnm7OAZIa6THFbyzr6
zTdT7h3aZ1JtEBgpG4kUUgf+NU0SPm54+lpkCjD4eIOZVZoqo7J/3WYyHbxXVrvx
C29xv0uFQx/eBmSbvxhs3Tfd+Z5eEHGhFRSXPnVY6JdmBFnHRhjtP3IAIn0tvdAq
OBGtjuLEb/g02lrMyKGcemPmHCLzw4A6rV8Xdt/YU66QWFKqQcqUVfBUr2NQIIro
Ulp6DVLzKLO3lMoNUA1cKB2D1cN+jiR72nXwBZI/yXpj4CTGsIJZHEolh6RzgZhJ
/O6O7FlzCa38ayzqCxuwDuddqWdNLIIYVHMYMXM+wcxKRv/Rn9fHzg7/AKsRVKFG
U10nPFUH+o6/7O6DQnjFWeWGPAnUXUBRRmeFxpphrMoUAWLC4+gqKeiVmdd3qlOc
Y+nY23Vn50z+PyN3/pb8G52ylYaWuZJnXlvQTmsDfONlirJEBk9sx4nzyg8TIRV2
EdNzigajSXQSIE2zgorJGLO2y7YB0aW4LQ34kBrop1KP5R1rVLw/jU5r47UNYOIR
SBL3e3JyOaj8Jp2d7UBFIbxDJLVpSp+o4Z5idrNymPDpdXWSf4Z/jQzzmKIAOpd0
+691skOPHxsiJ2rn1S0oKu9xScy1SGwa5/wX/ECZoWEPsS63HYTecTtTHnQf+Y8Z
MSeziQEMVSOvR1lXQqzehZ6dRAE9Lcu6iALBGQw9SrFGfNNWXFVwZovA1/+fn7xO
AjuP7rWebi8nASUbLOVyRYAmLlJNw7eYfq55wwsTVf2gNIn3fJXxRJaUOFIBjxzU
TvaAWSmUioWxz34QZMCNrP5BxdyvqM/am3mpgj9mWb8IVroTmDydiQ7mHOwj2NEj
mlIbiswqM1EkLuTa96aJhGTnDeHSyniP/beCE3t40L7HFYZTo9zfqzogpDDlDf1i
wk2sR8eH6O/ekbDCtwVnJPAHVvGHOWddcee827aWgCa6B4WwFAxk+HxijcQr1yRb
7s1QUgI+AUkHbLc9yYSJnGM1YqodDu7w56WvHgPAJTTc9nzMNvZAaxVqoZHlRzaz
DV+uqmYC4MfFpDxWyQra8qRGLLJNyIJlB0FrycO3KKua9nGww9XSXEklWxEU+i9d
/PDeUl+qSqgltX6KL6Cx4P5wovpjlA/rp6nItTb/cK7dZ+K1NTnU0JUHF+ooLXfg
1XaOjtCoOcoBBTvqZK3iqOCwOEaMt8lqLjuurmdvQnLf0mpmKqzz6ofLKV6nYD+0
MCAF35DF3Ypcf1z0YJNygFACVRau0MHK2UrmMBZEgfcW+7Nxj78iFVEMEWqqfYZ7
Vjzj4NozyZO0YMhATZNR212ebDlZf++45UE7BBbVh2q6mNgemArAOJ2jx3CfuvNx
1iqtbUzBHnp4GR0Atf2DYuz2LF3CjjXKZf1GNHNlhvlYKxHmdRmcYTmHNkBLESBF
DK2TH3Si37ro8hyCaNsZQOAMD4XqhzaNp+zkf5XX/TxoU7v3JGVfx1tRA5si1+G1
odMKB/DiP+D62aoF8RqMe0sYRFDKg0lDdEBLxyLcvyT5WY8zTKytCtY8fan8RCmy
+FN7fqd88OrPKaBzpWvw+AvKi5imJNa/5eM6SzzTZn0Ih8V2pklxj6LLxrHmpxhs
tWz8o4ghlFwQnjOGz8RzcURhadh3JmbyNLbfmPf73eY6t8mHodCAkOntDNVj8dPy
Lat2vFiMffwW6osQK5vIyW5Ek0X5jmFHy+gWgSkkLbeRJ8KoboApI9AWKSfALriY
bY/wWuCneyf4FKIJRVSF6tjwCa0LPOAaGg1PTONW6siTWO9+mJF9tTN1XvM2mPJx
0bHPCbbY9fAYLaOY2WMkEEEp8s4GEQLm91seJeNTbCYp15JQqqSMbzkDjWfaRTzN
PM3a71n+57Kicp+OQx5ToonJcuGsaAObSsf2EuBHNKM2IlFp9tp6Wi2N7bfjzwWx
vRs/I0iKMWfUMrDv9I8Bry6KDXPl5FqN0MphFwVHR7mLGHbuDa37wBV8gzHYyB0c
b8e8YyymvJ7ydpRsE+CJxaAtz/ToLi+uInJeA+p+TK2tHHANrmH52Ac4e3nzFbxR
UUtQQLPXltHwC7df9PzlJgwuah4ohbGgmyRlm6WDHMtP+sIuDVpUsmTDL3szCmCN
CjBswi8HzZ7x4kVOnRFmYSSsROTwU807j6UQQXJNpXYIG8TblAmCvz0qomggs6ie
u7KtBRx9tXOy23AaT5/bEY2OxSs5o+5H3+rWGhu+xxGAiSWmrV4Rmtg858Kg+xi1
VcvXnLIOF83Qr+P0PlEtulv7tAmy+i1U58WME90RFgZuNyRi7QeMHbhepe3iY6Q+
KEz+kxZtwdl9YO64wwxN3ABa2xLeYUjG8h9Ebgs8CUEUYk8A/5YIffJhKktX7sbg
52t5ItW8HT1Ihg0VPt9PbHZju9yaPraHiNxqHpPjmYHJLZbbOgt85YDxFy65zTR4
A+6WotcNsH+dsRYG+WEIOoSX2Epf4SYsoJ59VdNVSCdLEjz2oop0C6SWTcf/pv7I
kQ6pbkh0yZf1CXhA53QOMyXaH2gAlAAKzGaqW3iEeDIJiZ3kbke4YKJbEorwotAa
DJHfE3ZiuU/8UVYyR5tfPGd1SqxlvDYZlg2TOjlZdESdYZ+hMrL487e3VoX8VG2v
8Kzexn4htuL3nH4B5TJAYFBZVftzmkL67fG+SIoSawkwYbTiw7Gu/9fYuM55c69O
6gTuCM26RgoEdb+NerdIFyaJB3XbTjIGTNZ07vda/XgY4324L3ZRw0d1PpHeRKvu
C2J2fEq6VOzF4szI0/UIc9Ho/RJV8TG485Is2+3yCudpyPzgtYLhyXrQXBg2euwL
4/KWciINGFRYhuGkQ1A8rPAXywHYYbjGoqGIb+ai1Yxp2RoFdES6VVk1O6YQ4+fO
4v0lW4ikHQBhg/oYuSQEtbiUE+8EEWEfX7gZn2R5TlScv39cjHC/TywoXuMnAYZM
VdXwkh/i80lKsYzzJmHrhyaaBX5oLZZZyIVtLlZ9L8CCZ6WRQVjbQTsBnOsill+F
t+ykAZ1PAHh6fj6855DX8mapkTUISmV21nc/4l4fxxy0rujfWKDxHk7dDslz+JuK
C+o19ZY/tErN7lIVAuIs/VSRUWNZQb1BGmDbXCPlV/AEVgJwTYhdsjMMwzxCsXbY
OqLBZ3x6qBUFh3KIA7SKTmZc97oGyUQ++3aWOypTR5+bxzMPgLynD16W3pslG5Ky
0DprOyYwLPRGj73e7JbwFBDTXjjBgfc0hNZ/FgNEx313NnWdIZNjMcXqVVTBJIQj
kcsFQyIpyp8dTYZD3GsOT6wV2nqiEJ7Au4a7vdpotr9mTo6Xudp3RAImnXgVcS5g
kPU95VV9C6jtpBWyyyidEBhrtKYuN+oDyH4ev504N1LLhqfwXd3qZ0ccFusREbsG
CjyLAkgxpQMtIXVEQgRcKnmDLAFw1UQfKfwbCoPcLGPorMrGy3C+Xfo30nBoEE4p
iZVxelLPssvfXlnCG+4gZRGFb1igKEgjtw2QwbZ6GMZpkzjkk2lW0F8dwbOaXb2m
yoq04LzbOCfBSZ8ZB+9MmMpJCg1bTtXGuoWQWh5YH2/P/vlXooejyn3yNWvw0nek
6pkLI29JcTltWvvqBcjr34putp6UYZ85kjjypca/QPiiFbM+jG3c9vpbn6lDcorq
flGvAvc7ULJHEDJ3QLA/6uYEimYzCU6bPNmB4Cl+pQu4PyA1HPoHQp47gJILbKsK
gbTPTuF8ATrylXHkMSdkVSVp9BNMJnPiyw1HfYSW7OWLjlW+z3yBNpgUaGpL+tyx
ubiFc4kAaSPngmabg8Df8s27NZgS5tf6b38+BLHRJQFeT8dpBxDhcWWof0zIdjIQ
UuznqM6vZI5pVeXPjN0ZmqKYi5+Ry1prixurgnL2ARTPFAGIGA7GXu4/3LfaokNQ
RzehYBDIlvZ08IYHrYTB/oQAcjYm8C/sskbiMlMZfxphfq5XklvboAo7F1oGIm4T
41LuklS/lb5PciUMZcDn+ZXkTqvi0vnYBJ/59khDRkdfvucXNhReyzD81qcdlrAC
xjSRLrXt+bm2ZGFCMIc7pUn/XB9jNGNR/TmiCtlQmWaRa3xQ0eci6AsLBR3iSfaq
VH/WK4kKIHRv0FgJhIP5k2uVayyhbxpsZg3ed+pDOPCjx+7GjueyqRGMVV+JsXuA
kk6grEyssvD62U3qAv2EFOphn2e9xpSMzFZDMaDWbX2yAWn2YCPuGfwqY2nTh084
qMK+2AaFnweGjtpIO65Wtl2UZ9GhMO3sKIYYOdbHyE+PgP3Pm+dEwLaKtkZQOwGm
ucHgqnZ+9hPYsC/ZU4LSGiy+zQSYCM8khD5Oe73yBNp3sQp+VddAvZOp9mW4YU+z
lxDY+1n2mbIsS0amLsYZvmNaAbI3Vd2DrdfBFT6NQ7NY983wlgfbhFyzzsVp0/53
6lsbV0bKIVAPKlLAtdj7XQA9Z/MhnuNCevNYelnVxRjUnXCtkwv+y1uRnVDggJXc
yK6hA7v/mY2gwIOMKz0ppc0Ivle8a3GRggLYbRV2MdKPXr6jZaaFfcUjJvu9yX3G
3mgW4Vw8bWNEGjqzocvP4tl6+KGD6CGEETMwVfvL4KqVpdyDbRWhPczfXICuDCA+
VoXP4UNbNKayOSk16tUkDPEECFawlFjh4Le+7I61UlOTdyq2bliTQXDc5+SSOnjj
964gNNOZr3WCYlJznkkNzp0ar3F9pgb/yVp/4bVJcZdqCmhrQcjlR9pNiDJJDZdI
WEkVsdbgrff0Rpkz6FC1i/h+9bKWkC7s8yD66mUgXvE/XWnynXebbh8MZoLdQu3S
TJi7vrXyrRaG9nIh1mSwqCBSEsLa29JuvqTeD2gPu93DfLJ/IXpUYJgCjNdByqC/
yIr701R1+YClOwq3/jAUHTLTIWmXcp/OGVbePOq3sqrIZZ0hhh0AbaNy6ETfG4h4
Mj6mYLdLIl7tcI+mbg2dQWeJT1adgSHxbQkjB2M/ICNKmBstaVXvTBJeNA2Gi3Vv
kNIM4oVYS4sOxIpzFFguRvc8Wa7vojwCrEqithPfjk4612q82nv9LqeGjUOAdaIz
YhpIE0DT2xb7aAnayXjXfOkvOjITpsCuyFvmEX7UOGrqkUHYElH3O5xfM4g2bGvF
Z665DlNXLXbWF3SsapTWr0IkPQoxLUCreyLnYZQLLwoCHrZu+DEbHg7KZJSUn7SZ
qLwZJdm6hmeSz793CoSNMpEnsyxruiq9h2cYuBYOnXTqkO+rXOkS4GwR12yX787y
R71+rl74JnvVq1Juw1pvZUOV4b1STAWRRgyx3HV8NXNuEKqSjuqFtDOjXk89qDwF
F8Ym6A+6/mA+Uzv3VTaALSi3vTvXmU+ht2BHLzgM4yEVNZwUU7xYcC7G+QoGTlls
YeuE//eXGsNTRRrRMamO8powQG25wffVePViHrvbLoGMLhphvVFrSPCSXVtk7NIp
yUYJX4W2LSrDDirvDgOFWq3rj/brnr0AJ1e5hY4CDF+emN8SjWLiR+12jTGnsP8G
wKh2qgKiv7a4oJWpfVcLJMKZqjZNC4lk2uW44Hv0bgP29IwjI09KAZfBL6DWF9E/
/Z6Pz4GpMduSleuvla4KyACJGAWuELl+JWaoKLJCuHD9fK4Ou4zlL52Voke3ptIJ
g5wE2KpEhdegyz35ulAq+NnI2sC1D/e51cNfb5uG3rB1FBZ65zrr5mxmlG+2ed4Y
kA5UCDxOVMqi33PcvXwrFG5x2xy9EfBkvVLKnlwDRvesqIxHstvhgaxxbkx+mRQX
y3DdOwXn6P95GIRr6Ho9wRRyFbcOocwtSHR2yJQxLZEYLGf3j9j4ACDlpSbfoEwr
ihLv1vGsCqTHJECZA7wesXPHT4YLAEi4tSlvNWgatY8+nP5b6q/6NPo4lvcjBp2N
v4EJDkgdmJvSVL0fRgtzsUTRra4YAWDKrxHvihwaurGkD0ZKctk5413Yu22V7It9
OOGMA6Da1pyHusSZg34SpJwxQDI/5b7wDT2mLX52X9gi8hVhx0sn4buengZSTFCD
e6iKZvQAr1Foi+92bmv8cERE8Sa6aCehyXB24IXRwVFC7uhqpS852/BaUEsjw9a7
5j1WCgcpXUK9uphxmLG8qOFCd8Rh24JkxwnWmaAJHr+o0XbBsXMRp6ZPjFTFD/ov
cmNUs3660jCqBp+B00Zm2SUzVleBiXNcp7z+mg3RmfLFx62HLskeJKruK7IT/M0+
GwXLdKh0gdbmmVTo3nDiExCMtI0zlB/kePbHWnpjqVJSWgHbd1snnhlIpRDtsnUz
TWbzuhea2HISvqggydnDFd0Nnjzyv71Ml5ImkgfrWUaBQtw5ueDywBYmvzdt42Ab
KVA0O96+NI48srVmAZIMVDPEfm8ymnUMkrJ4MoqWV46HPfILDbf9Fc/UT/GWYRfr
kmEGi4e3hlQ1r9x/8pOJG1OENkM4DMIVHfhKYsTvNJK+l3dd3Rcc869UytYKEbhl
CPt+IJVpHU923TsnTxE/SfSS+dK8DxXcza0VQQ5rNc+HpS1UO2GU6R8WuAfN+C2t
CStU4kkmEXMqllJwDIkHNjaEQQhNVFWxjfK0g1AmO02Ti6+WCqsQIw6CmjoZwveO
QnnBiggbelvFYTePtJ8mDrqFxy8ohndCJTiCAqFOg330SkYp6sWnh9HxX+rFU9sn
38S23DFCbkLp2VHNboVbJ7N1Tq/t3umAvDyofJDItNT9srqjMGyVItXW5bSm6u8p
w/X3W2VEha65mbF4cYE84uvaKUJmnXvShGilEtIDaaS2KpGrZmUYap5/s70Mn20H
uQO1dl8O9vSHp1lk16lZsiFiSGu6a8Nhn3N4xNqIgvUrMlLaZ+IMIYpPxsb8jLvv
qt/rIkH1fj/1FyXuxasYSy6mbIejPm7jHKChZcXPtxWLKBwo3oYXJuT0eMx2qA4u
dZ4Hg8UoKN514iYzEzZQ1MIIcoZwujnGjOhQ2MZZ9MBVXQCrWycA/giETfYhRZZv
OXcrcejeKxQ6C69JCtpJGwPi7EriwMIbBzvr+PHhWillE+Y0owFsgMsfjMIRROQo
sTU5mAgBVKHJfz7mjFkycsiKLWIKI4315ryiEnQg/UYjPHaS/FDoZby5N1l7qlKX
pQ5RXamAiNqztEzv6jrb3kHQNC6SR+TWS7flOnoz34ZcY2JE1hJZ4B++FcLO8A2s
rAZhgqdT/8WknmZTDxGu3UORnPSRGs2ZGiwMyySGf/4TWHLqvWcUHhnMwHfPQjG5
59BrxlPk7Xcav9n8QtadvhLwlPQ2DFyj4gXnGBiZkf5XJXjlTGwUG2zTQyQJ2vJ3
G9FNGmRXtK7Uc9ZTz9uLcrlSZV4iUSvwU1g/uvc/6amNBpwBmObZK0RItF8NO4aL
pRgDYAc5Yzv1PMvpik0Gwp3SUn/pYT889yB79e10AmynkjmBL+9ujGmpNmaUOtx+
XIjVkuNvXoEq5ZigQMrvOXlAgIoFVBjH0rSjZHf6Eya4ZyIyzWBd2JHcFTAZwOOp
DnNt24GtqbmuBq/ewSqvEyS5KUG9IYP5M5Rd34RuProiVxFtY8zT1E6jRhnP9+u4
NjYJ0cOIhC2/opwzCYT4FVUDQEoyZscOmcSTRhVJYRxV1mwIkqkkxT2Bcj7n11A2
k/40PFtVxK5wpphb/SEYUvgsJTvWyH5tY5UpuT5xbXTCIvI1EyscQaQgtKrehLP+
Q858tN20+ubANxHvxF164yDbaoNcoDRnyv9i+tp++kealOyNUiiRAxXqn0+gFxN6
DzB2otVzYbe76IMgwej/DCqbzwJEk1B3cK6qPAXXDYJCjyeZs6FklxjQFAMAf2Nv
Brafzp6BHvSicuf9kzRdiH7O/GXDjlT9BBhBrjhpPYW2OxIQ2Sv0ZI/kmNPapK6P
t0CHlj88YyhaKJKzBRUo8l6E2+jmW8TlZHYhN2zvJPMb2+lrGpPAPtviEr8VxYOA
vYEZ9oQeZ7//dANbYh7FV/r1Wzwwwcb0Mdv3rzbwBXC93J/xHt6z2yhB7AheVY0z
knt3Eq7UhV/bVmYl874cCWQgEFpbs2zKMvOCDSvslqIsNfzGJ1DJleV8hCoub3i7
+EunoxQSrZPVvvBd7tWHpFA27sUvOxnbVGNo5n5xXfg3Jv45iShlkXnCiHCEnj9P
D36c3eT6Oaj8O02NSnBn7zX/O85vDXl7zcHODYMxkcqhZxCl/MbxlSge1NHZ/0y3
dLZCicF2gkDKDa7GgcwK2bKX+7vAqflUeZ1DhvUp52rifwnGsQcvryZukkEVLsV7
XCirNdOMZDnOCFMAjA6VVJAq1h4yzRuZHES3sGMkJg0TIzWSk5g5jQxRqf0ZFtQZ
sQzgqQf47eyl3m50Y3239o80jZotsrSHHSwyx4jvgKdkbnqEeA8KieJo3C2tuMDc
Dm3Ca5EnNYCDHOF1+yUXMRyzyBv7LJmPA4FD9GsB/0e9rX2r7II1NS+WIjSZjOcI
nXAfOXoli+HX2/w1HR56FYGh2P1676oI98R97kexfvG8I069aP1OrzYQ67kk4VfT
Tda30O2oGakopIljKFjuJ1j8+KM7qjYVq9nodBHL8eDW9NoUALMMWkW9DEtZmVWF
uuhGzyddVgfeT63Dg3ZUfXnZzm81iDldETlauYkflYLwJUeBoyWcZawJuwjmrevC
3zn+ES6xnYRvO4vltON1yeuMWwXCnxSWCbNnKBd7SMinRF55vKM9LOJwqxqL576+
V/+VzNEkU7iyAl6b6z9Fbv2f5HGoifgAbnRs0/j6b4cZy8wfA+CISxMxhBm6MfdO
k2dF47qIsk05QilfXPs+NH2RutPIw75bbrQAYSFBaM635EMrvHiHEjN3DyCAL/Rd
RebY0m6ZBqmT37cjejzO9oSXmm0cUsniN81stj7UBjUrrRzZhG9dE9Gqpm5PCdFV
jJcPsuCoDqQvoKBbhcdVRXZFJ5EFXAfi96RLayCQcgZmhsqlpASsxEcpnwSMbX2M
yj5iyyerLcI96ukekdNXWeLJY7YbjlNyK0mYhVDdRIaX09GzMRxOInEEyMWL5y1Y
8n3VFClgaRKcseVbl50C8Ta5ftddIHCP+3FgszKeeAVvyNw5b6+z1NKvtjC4292H
HAIUimekCo1gYaliHRZX0OozCFwkmhybFe7HAVcXbcq/Ue7vJk0o3BomUAd29RCV
9VOx+TCzpCcT4Tx2bJWVkIHpsL+GimK2G1k7BfauLPJw5YmhK1gAqBkmrDw0ZM+S
CXCv90alGR4tE+Sqdrhe+6ICaxqIPCoCIfLgVNIu4Uwjb1kY73/JyVWLkrQTDdBi
AkVDqmOI8pdhIkck5kPw6aZ4gFlpEfB6zxIMOTDZYbbX5ZWHGgWQQ+FC0BOta1yl
HB0/Fv0P8O23v7rzaGuHpIuTQL2xSh8DRqym+ydwi8UNdH1x60HQSFIMyBhrLo/n
R3ipq1OUSv3kENOvApf62fEi2LrtF2owDN5rZWmIDRapqvDDTCMcTYnomR0SxP/G
nYvvtYq69rpwBtBv3S+bGxYhUUDpMyBDM3LMTKGTKasQlF12xyj88c2eXknkKQmZ
xpFs61WcWef4bLRdafEp7swwrXi0T9SXQQv/NMt/o/b6ped4ICeBt9wfNDIH5l0X
sRGrs66bRghs6m06lUcjKbEHf3b8sYIFf3XRMNlx9BxImSuPvqISPHSKzFYxH4zP
5xW6P/G+AyYMTwnOi5Hd6lPfJ8341fyxYZOBiTT8D3EJBJTc1G4qLBzJN3ayFoON
GOxkSqB8Ad2tHyq9IJBZvSQpHjGDfQeNpKiJrf+sZcSnh1gESfLlOZFQS1ALbaZz
jaDW3CzqdFS3DoAiBan6X/pNx3zztu54VjsnLnDXYwoPwg0WZiodqzEKS9XChxFF
f38Phx0AF4J0hBYRRA3AJ7fX9uhJOWMWN+R1IyIbHRYdS5HaTQfRIWEIjHR+vjSK
C7LabwTQOLqeOBp2Ndhw/L8UnzDneygwN6TfUWVITkJzUzNIsLXzsoBUGO0rPCcZ
iUwcz+lmT4g8v4LsdXyYqsXoWgDWUr45d7QeJsow6KGifYfVmHS/q2ECGcBPmdqn
5YPFs+ve6NqPNKu3Kkb30aFDDzG5jkckT1CcAzEn/mRv60JeZUcZUWLj2Zn1FhbC
E6G9J2lKot0Kv9raznc0XfAubqA+TmXw3pn5MTHr4OWCuoYrh6e+UfegHYZR7ERd
Rx2bn/I8L6IxgbszQNELLjQAk/1pKqpDGcsWaonrAPyl7BwIv4YWjQrYoKuhf/fS
GI2y0Ssd/hAPYpUWLGqAof0klUUln/xIhaa0KAPuFpF5wFhGTb1XEVj69lUir4Fu
7nqlwSNeNwiMWy66UhK9QjgmJBuZ1IFRRMedkhr0dGJrkqh6h8Ajx/HmnJxKe9YE
smdlc6iD1PZZerUmrmEfMUhBAzR6+K4Dg8O5DWfN3Qua5cxJnHIpKTRHIjdmHxUf
IhETNZDqwvkiP0ubmI4y4FdUi3JoG0PtW9RV4y3V1OxmSciUu+2bSANUMBLE4fHa
O7t7jxg3bCGYBx1jTyCboP9Dk+nCNOuZP/Cu1NH8Eu60vT/x67olS1JUy5qSH7yp
gdNg2+u+MoQ3GcEJm/zz+HK0+ehAPy95j3IHl4KbfM9HSKy01TIw/YeNTp9nGvme
pci6twlGFJH6UFlXf9scoj8Pw5YIgfJiPSKy3VoCIEmvli6WrlhY3GgJs6g9wUX+
gFnpJzQNGozbdcVvTwoBhaoegFKkOsZL8KN1YUX+Kxyk2BLDXR6mcrWSYDJu49L6
0VKOPb1QUVY3CcInwwvxmgC9TA43T0g7IyyE19FxxvlhaZ9hUiO9EE7ZqgDUqSD4
0f0IRw7FyoG/3ME/it6mqPWFEDq0IzcPGR3/+FtwIAF6I5F7u/AK5QM4xlc9ek0F
bD3w44BM6uc7nMxfBkuIEnfhrSaLTeyVr7hORe3XfCyaeyP7XTHRF6evOEnnXANH
AHrEekBJrKl9q0bJiEX0q/WtgzIpPiH3xHmdUk8UoHqqrXDBpIDqzrJjTBjrgaFt
zUYuUweAKfqIc0UkQz5wJSK11waXQWrYPK4vi8sWyUWSiYjJylEFsQnWLTj1qPI8
F12tWJYuCvgD9xUYV2j6URhwc3DgItP3CrXpdwsFcKz9RTTaAj8p0EdlM4EAT2BV
yvVvlqbL5UcMydmoAXTKC800tgULDbDH0v+EP1x1yY+UbIPgOApwO8Gw4itL6njT
3vVsHMOTfALISHb4b0KgDM201J9lpPGiqIi5PQPuY3kSJRr3F+hNmrO9Kk1GxEu1
aBG4aYW11Pz9hnMjT5aqRSWA4uu6JvjUyWD+LXuBNrUH1NGQtaTiffKZOR/aT2v3
OrbVtvX+ixWn0/HMsqpzzQUrd3cpS/60Ie8o1VadBRLnfc40T3zAkRS/ehW4wer2
6+H31WeuMZkQDQWyGiHYXruD26RbXWCsGH2HP7ie11nTJktEFw1wYX39nSz0pyRS
ZlgE4LO8NPhau+0hkBSMIbOEoz8DwjIDWS3cXzLsSJPxvGoaTCcORcfx6ZafoGY4
6iO8McFWqIOejWNayPH6gBfmS/5jbYmXM5B4Zys0KP8=
`protect END_PROTECTED
