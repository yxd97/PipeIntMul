`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ua+JB1riCnv6jG+6Rr+jyfYXKns4Z/UTQOcgezFggF021f5P87g6d78cYtjbLT3X
I3dMJMEW1fPpRFhSzZKnydDWnrCyoN4S0VLVANdhf83ZPh+l2xgoeYz3xxL4IQOH
pt9VmCQbrr8D38qlTOBBK7MdZZpQO684PeXLfNf6yzOysncdN9V5ryEGFG1GkZ/a
VJFALuLrTS5yuI9fN/4ACIMfRj0DPkVCTeo3BJUi4QFNxcP33V5dJsOJnvCrBq5d
+PQpb06qiWiOFbcekBxM3h5OIs8vIqAPgK/i96nhQIFCBvTVoVRtdbq6TgVXbGRb
Uktp3UnzZxlMFur6OYU7CITmJ171gtdJto2y7RIqKrjX3HrLs10ZT2OobqMYPONC
PTJEOo/YDuFuJjVS7Zvoh1azlKFu9D4+7f3O3/N4I8iuRYvindvC62lxSNwkvh0a
uxEBDgXhE59IBXSP4BCZRI+lCB2fnJWsJmEXDV0NtokiZvGRC1Xd5gmMokJP7LSw
iD0ZF28tvIEtX3tngeTkowPGbrPPgV8nykg3SlqkR58W34+aDwQxxd1CeeNXqyfc
iiZEikEKYwPglVS2TcbUKpym+3TPEC0gsZqxBtBjM94TqwLXIWYIFtXQrNp7IiwZ
NiUx5DjxQKQxzCK/lccqqz7jXIxDG+eLYzhD+QgrrJFLM+uUVXAmKfxN3uGVAE4G
A3i6U3xJ6kIK0MQBbDpdzXIAHE9LudCWzKoXUj0JaTbFok51/bf2pVkOrVpDkPYi
N8LIy0OIzVSVvvhWZYCzWqv5IU/94sL/69hzHRXeuTM=
`protect END_PROTECTED
