`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHpw2xCfuWgDlyMfmeM1L9dPCoys2+FQvy2AdSz+bLV9pXf0W5pgnf4rW4P5AACf
Kxqo2ZahUIt212GmvbfJOqa6Mq+EuA41qksv0cfulskEuWQEMrkwbVBNPdo4sa4w
IDOq3QcPCxW3h46X6ilPCDbmar7/ImSdb0WO7Mcw1s+cn80XDFkfPjJiGetfDSJJ
bMNa1nIAfyLccWVBjbu0HsC4DVI8hRGKIeTknhSmM501o58BYIq1B8TBJCdqinL4
FIs8MMKImuwPy0mBSzsw71E2+VS33BnujE/c3BxmZQCKwplMuRgur6iK6+47HGDi
6atzGbWvdxjeLnPDwOLOI1ZEDcHJlLxtzT+kZlXeApcFEDUutyAnJq2ex12pXtOX
t7aJCEN/M5TyQt4/lKkcp1LvCk2zGig6xOvwI3Rblj5j8BCaplNiB0aaN8iVAIfK
dnoZmW2H955QpI67TUAJA1PirQbIAu4DDJXFJwP0a9flH/jYohaoCVMute86aD+W
NhL2lxhS4S1FlwD2SFd0DjtkyiLcmmi1SoJF5UgzWfUEJXu4KVqbgsKOj/ZnkbMJ
4XFi5s1p45QJ+GM4k4iZaqp7L97MuIgLy43O/1LJMDLot10DQSKfbvcIidiL9DAv
ISdqim09FA4HBko6gU7Mz3Xciw9C+1K6ynk0TCLMtSDKF63mkVRS7GB8DJJdU+KV
E2jBgTMCb5f8skG4FPTMlGPLClPTIVtAsV8BBJ13w8rq1nWvIcf4RuWD7KbTy59V
gzFx0GFFrYf2ALpdSKPBSQb2p8DBLsp9EsbHCYJlqjnrh55HbleTPXTBPBSSeF9Q
B1lfof9a8uRP+LngswW1okVCYsOBMWWQbeyPMMg2RSo5Me8O0/2Hgtndsm2q5UYg
Vz8qBQqSEBCl5ktNs1Spt9mGMcrdyRwV95413f71Wc00aExEG6LzJDTdd2MKgnfA
yI/lKK2QYa/2EnaBCoebOR6JlRvMz3pcT547bFftYSqfteGyopQXuPbyjRPlhHQP
0zVbKqHsXm5N/a+2HOmpgNKLFKeI4wVwe4n6Be54bJBTIAeuOdWAXEW68HlPhTOj
8gK6Q/yJ7zj6ajU1lpl+zAZv+k6E5Yu3P+ZblzcQEKn9qeaK1lzxlDtpnfaYU8+a
62hbhRpMQPkObL1M5Q0cGm6XEoKbdOLFB0r7NaNu4LzIEEyZkPNRcqoQskhq0tmd
DmmIbk0ebd+cY9lgtYG9eNB46QmlRlryN0HRSKIh0F3ZpNknWyX8X2wM59AQAunV
ryz7s+6dVcixGL4dJZiVrA==
`protect END_PROTECTED
