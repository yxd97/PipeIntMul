`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Htwxn9UDWjZJMyQJ3+Rsh1PYXO+a0gQXh4/S9vMpfSdsZm7mJrv2ZHEqQT8q+5zO
i2DRh4bCBEshrzP3jBfyLlDJB5o0/TNE1mSvnUOyo0bZdYYumZ5nv3c+wQEQcSU6
O5nR5Faap9G3o93LjGE6v/eYu9fHCxoHVIRwPY+Og44XkXGYTS8CqdCy1VMHqLAF
JugCtBS3F79xgJ53uK3cedFab0vDePvr/IAeY9iErVwK6hDmeFrko4gEjgENVfOY
6ei10W6XvWSd2rxTA5FVydpDqnoLLztYI93NEBvXAuLTeR99gaFQd4666Tq6TA82
Na/EZwkRdkaj74Mm6vgqcA==
`protect END_PROTECTED
