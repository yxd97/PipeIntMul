`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b85O4sEIkiMnBSx66/O7sU+DczQUVjIozjNtLryFqqKkgGcQ4WB8+tSAMXT1xrbM
MQZ5r2Sq1IczZDQ+Fs5ZukTsnL3prakijBpjdbaJ3Gkbgknkg/kPGa+iotOZVQ7a
vEEYUJCbPRY/ERmZ3SN3i4KsXUoD3iProGGECMdJAzodLt9DNAyNZPLVNvtZtbPx
nCpsAgx25b5cCDuJRZOjv1RTWBSDLsHlXbbcNPmcqEPRp8nFUUd+de+RwEVT3JxX
+PCrJZN2pUqQ8yEUZRjskujExHWC0g1MzovTSF6R6Y9lk00TPNizgR/6T/u6r1Y9
bl9Q7PEzBTGakHk7Ds2icgqMKQWl9lLIzOBKfWWSrN1vFuiZFLAwgsarUmZywnAW
iKIRCj4uE9lWzWUiOXMpobp51TsI0En//9wQSe62K5tYWCd7n1eEJ/Q/ec3gU++F
7khQzdphnaOG09XM4vIIVL3x3dUs9Q4Y1MmE6Qoh/GqrGskMgHD617+56tlZAM2l
dem7j0CtqJ6pnDT+T9iHDmU2+WbTQwGmRDL3POF3N+fyB8bWEOmNmGcJFO69I4kG
eHH4VYzfBCPXvrUa33HyBpjjfgMp6MMQE1Cg5LNn2LTtarD9aBJ4Sf596o6FDIuI
B2cTlO+prdSJvipqny8ceraMnUVpHnI0BKRhKdrqxu4=
`protect END_PROTECTED
