`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oee8HcnYOiWrBD8VS7wzP9zj+OuICILCfnADYZTTJUwklxu2qZrRW0BIIzGMWSmv
S6NWYYKNDIgFFviV1zikseR982Rt/0eKIraUC/66Uc2+zumuAYRb7tqtyegNR9F+
MOvOhJTIA3dHmT8sWpncDEYqoOytc39wqqSZk3DIsuDlfLadps1PWQrs5DD/Xvtc
OCUPpbKlbFSlNXWxL4dAKY1vi3NJbqeBZ8LNW3kDRBMEAS+qGEafiUWBlyFNiw2O
PwZczjyPW1NbObW1cPUJSt3gK2J9uKUoCCOVHxwPdWd50lgtMZCA2NhiaGSHhksx
`protect END_PROTECTED
