`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F3a2Is8ldMHBe9/PxxZaEYgOzkY5Jkql7RdPcMEM5wrZAUmIUekbKIGxZ9gcs8sC
7QYszFfo77Rayus0cPR2AjruCi0cfOzdn65RGru+lZ3465lCvn8NMrv5bJG1m7rb
iatwGbNUBwZC+fcckqAhXqH/IKOpvB3rsfRKDBxCcYrYT+JvE5u6LWLLb8inRRqm
o/VwnzIDEiwbBYZ7pzC2UL9oGEfK/TApQc40iv4SGHVRPgYQ8vHZ+15RU1CTG78A
0BBOOU7WXCq1fMcyl5M1gRZFJuApA9tjmPGY7stXrAOX1Y+qkpa86yo6AphlAeGr
zOL0LhDLzN7Sz3uQ4ed1JJNZrrj1AAiIpmOHrFD/ncRciM4B40b6p9ddKILCKx54
/ah0dsqCPTcFNs3TQRX2gK50vu1lr7/PGpisi6uttzNPZWrmUuEXvpCJjDwl3+Lc
cYh9VAgiv9gouo6+Vf/ySqOEAupd9NChnIeG6uYQiMld28woEEeE/ltcJd1fhmJU
GWXSUqxrqPflO6P09oNAlsOQwIdC2i0lr6lAI4P4arYwK/vwPppiVmDkWYVXrRyQ
R77LY+5gZVZ0LdtXPCbgL7IddHqBSlQN1+p6b5meo4aRf6L/MULRoBM1TpKY6qD/
i3UApoOYFCRgpztBm4APpeF3FaKmHObkydkEYOHhCNgpK4telUFcLlwEEp4+M51Z
Wml/WiWA2M3BWQnIqHlXX6iljrLjMW1zfCPlXRLaD5EbocCokMp8G+f2WWZ/+Y1H
T0IlHHugEv3cyUDCfiAU7n10q9Z4qySrfekm74aWZp07ZcloRwKA4fn4pHZwUlhB
6M70Pf4rd4hqqm72O72vIhs86kO58KfLMvG6ZBWtgK2yXk/qZVjo4yQizsw9DK+2
lQI+p1fG40LmZAXKe+PiBlicPg71Y4XU8ouxwNLTjkku5RreuMnmRxpi6DYzo3tW
LDL5hOCwzNL3okCjlQ8xIJq/Pk+NRtU28j8wgKwOA9jG9Yk2FG2x/YMiEHHv2Wbx
WYDK6Cw5cB5/fmG+zpa305MyAED0b+QJVi2L9UwKNB65YksvVKork9Ht8Khd3VKx
3zntLmFz3RikTQwFgPylhjHzaxr+xMQoU4IynBo2f33/Y1n/hynaSM3JkZlm0Jjo
vatcFDycLOO+0R1QisHhE05WDziXS4ld2Zx68FToBJ2YQNBINNsslGPBi4dpU/qI
Em34rGMZtfsxAW/2VjVrSir1BxC4p1rRdY+dIBBPoRiCEXaI3DFgJcaJnrsZDEnC
794qKXxKYt8SP/FajnhoZNqqTsBonXdwa/ITfTlr+36T81r5HYzea+RxNIlknZgs
MrcPEM6kj7rIzSTqrDcgq36TIHPE8lEA9N60UgelOVDAZrLEgIN4wvIJgQtKBrYy
OHkxuuYavURl26OG5ajHKkSPmHUVMBRCXAJiUzWHYrpKTNR3a9tG3faC1mM4MadS
d82yN0LaQc0AdmpvG9QdRdkrl3mCWb7heLtHYL3xUuoeuhJ/PB5E98MNi7dDGKKK
CSfe9kkp1sWcHrMFaYnhTClmqj7W+OmeHO8hKWZVmCPMc6Mwima13iiRV+X7SeMV
Grlr0p5RrIHVW6qzkO/j85KTHXPuWf0lN8/fUjfGNDuPdRxzdnLnlzmlD3UivmB1
HGzGtiBfpagVRvpNIXf6UIYBOm7mDU3vZuJW/4Nj6esFiZP+UnotC9rM8d/QroI2
OQkS+5/AMiJYQfa+RBcN9BFjv85526j1FpkIaNfqGpvI9ogbHjoy6/L8bV6DZX1K
aFM9qnQOMVThx65sqW59ykdeEsF2oemjqA5TVZ0KFKWaSrTFE47R+n+yY3299e+w
l9Ied46YKSV06S+KCOwtmiqmr/NKtke12zo1bqClfPGTp4MmtgZjjGLef5KKjAAq
ENXr/jyqNaOnGr7hYHvsrNC2LRqZNq66a+Qf6pWpoMtLOKrdBVt7NvSkpSBQJmZN
Cej7AlpuHeJlDI0rGk1g/NxtJsFrvoSlwcwslt/fL7smQzD+BWvP9ZJIQFKC4ks3
Az4uEj7HbZntdwRRgLBSmeP5NmEdzmKdNTzgmDBZgwDjF5oppG9htn4x5Hgv93EM
p8mlwO3TRiYBA1F7KzBaz+iaI2fDQ642QsDYQluJ7V3bFNxazJjgWI2aA+PxkXYl
KlKP+v2zv5c5Jbp/cDLJQUmvQiMNj/Uy2hd+xCZ9+ttqf+qyggvxxbgyeuGguWeI
O6oPlyKOlYdUl1h5OBX1dNmOWnr8mkAd2s4RyFR/libVrL5jL5poRF3b50l8ULTk
o0Jr8vTklLN2Gdrn+Ie1s3mBzfmCOpaLPfd7e9eSb7ULn9mu4J6+aRywpy40htl7
vNe2o47De58cSmQ3jgXrwvxe2ocU+HU7mQvdTVj55+KgCJbtdCDTlzlmHlu8eyuv
fA8WckTsqFB2OJQ5JkiNfYW+TudB30IG6KbHGIUby+dEm10nItEwBuPkTupY94KA
tReSHTDu9aZUmgcEmsgHphjUy4357S51DjkAIZOWGwixbM7jJlOoVAaNlnjnvyrg
amYpPXiboez2/H09/4YnBkGwHrewePNd5UQixz5NKltRoenZKJCrdRudN7Fc85Nd
Eqn9M29JZga0i7RVT9FLYcBjGRN6l6pMz6yGKwnmR1fTdz76dQ8WT6E6uTzLsLbM
y8KmCy/hs900Ssz/oAEfvBJlHeEchgg8rirLrUiOI3FMkd6sM+tb5nDAEwH8qXM2
qqgL8CNODcc9hZd36r4R4BY0GLdX8MdWtNCZ6DaauRQQCuiKPGp5nFYywq4W6rSE
sCBifhyj1oyk/tlSN/zq7gAdmOl6IWNSCS751JyeMWeJ/BfBZ7j6FKKiLEOXdLcx
NbgBrzSSCnwaRTWZYnEsgDb02mtethgfINFuqH3yGNULw7GvI4diRFO5MMCbXe+d
isPxJiKESFkD4Vgid1CSEak2Py/TbZwDoRooVgksjQE7D9a6Hd7usfnnnHzuad9h
0S2wmOEab8prNZe0Xptrq/cHW08N3VDvm1T634oyWp24kHCzKUReH7QUqXZ6VrfH
kH9R7F/F2PPTEzwHYA6KuL98uL76uxn8pGP2RS6inE2sAApIBgNKxt9urFYEmjkL
NSKGjedG8eSSazCh4PA7q1N+gqDYrB79c1BJQgWg5jjmyWfEGiW1rzUIxsE/gXpp
QbmduwscMJbT+Gbt6XmxZYwGP1ubgAFk0j5ZlyoalcIW2C/5isXrt8rPIcUbq0Fm
3ca9HqkkANtBvQs+N5pL5A86H5jHuvsOYHmIU50vzweyH0jg0/KoW3hPyfoa11o2
POzOyK2w7nveMtdkAmdmR/SYAu+Y6gfJkPRzDdccDeRlmGVG1/h6+3X1wqJTaEEd
8dLQHh0iwiaJftWHeXr3NU3kuQVRhjmPHwMZ8Dr+Qim/0Q5RmVDQC4dr3cf12DAp
uhc/GQULcGVbE+gwfvYGotfQSgT+8qhnbKUcTDS4Sp3tajeOVic8x8HBN4Bqh4Fa
UdlkxS0dDJBsZuV1I8JoV3/0SCiuvl+JpA3zdDi+Ch8Ui2fi9IDWBl7UCG3Aqq/c
m5sh+nJ+TqnU4Hr8sYC59QV5J/GcWvqzUwC6R0lt5M0R9JGrLU6mw3F4iENJCr3K
KBe+qG/DyBHU0hOjPDCXD4xPbKbrvg5B/yqCpllroh/sWEtmaLwqLUpLB0QDZEef
FTt6iP2fiQJlS+GCHlcQ1Hdj585NCLlMCnH+b/cTGr3IKY5L6wHu/VUTDKaWmLC7
KeBbWJBwSdUZUhC8dU92pgaVxKJUF1SNLwKuYzP1HugcRTeidI9+sFFbxiYH+Mr8
QKuE1h+zF/4GfyOiFhaOkYkzHqm+qMHqbCUkNJAhH4tJ51vjCKh8O/QPx9bqu6Fs
XpnKr3R+ptY39GfjfNctsYm8+tx8+mqCOmO5403xkqj3awI16XLWM+f9qkaBqFEt
k042d9llXkarME7zXpbBNZcMM0bpINtaHVTejnD9yaKtAr1oKCsFy1DmSRI57BTq
BwrYYNxaTrUehnV4JTsX9Td9cNdYw99m7y8bhB+7tI9MVK8e4spE7S92FR4f19J4
p9iQP/VNMd42PYBRjd63UaGv7cqm2HLlqPgXSZSACydmAwz+nWYmjkzLOwTHwGme
SwWqLPBPh24+yQ604+HabBIntBi5giqEKoBMsbc1nDXTEnAXJPYqksLqV8JmK7D1
8mnl06Pwy/p0nWW2xE6RUZRQUsFkxaat5eZ82kMV8SNKKB9Qdat3wPNjfvQFtDjn
cAFw801waf5oE7wey842GfMbr7msgF1bsODy2bRU6w4RdDIh3c/RJvgoHp0e1bVG
U4tzrmDkMd1l3PvtyTleHZ1mdfUeP2gGJeR+dH56LK5GZQuBBJOy4O6rT8FKk+Dn
8ofRc8D46byjS3mq4uGxoXoJRzD5nLfGbl8SJeVDhPE1VNO+uXYOfBHiobX33rV4
jsgpUcXODjXtXiMMcTVsr8eFteb7kWMzqKc0wtY14Jt6Bn9MBE2rkW7gV981DnVt
cm6ma8jEGDzsZL3+a8XGm76eeCwqE9WS+ocu5AeTn3WFSuQw5WuCczJU7ObysqcZ
A+k+JGV0sLyGzMgbCWTthIRl4l135c+2uQsStue67SNAgETGrUAF3sjDWaVYe25C
orOE2SVlU79Q3PDQtj89kFcNhFB1Gpj1v6Fh2I9e9ctA9a3GClmszmJgs1b4Jegg
4o5xR27TV8ze1nDR9rwV0oj11hvLS78coKRZbSjm6tmAhexDBqKPnkI9NBEYPCtd
+H1hbzKNez9l4xuNwdjPGR1iXK592Gg1XkN9o5ovgrPuocCv4IZfOOnTBaoBmVAe
42ibkL1GVW2HQ5R4MTeUOYxJNY4xzuL8n5zKjWzyUCRh+CW8eOOKeP/ZYCucxt96
QIlKn+oVmaLzAbgWMjvhXteVPjbI7tM5zDHReY+tRx9TyVn2nBeaD5B8RXqPJ2Dq
//xAko42u86VJIvdhtXT73d1HrrRzRyqvL66v6YN8wRzR9SPAE2GUq7cOJcSWey3
5SqnbRCrVF+w4Wcjv9vhGQhfeGNL7LSv9/cKfiRyFCiBgix0ZK7eSCCTUhGQmMFw
Sh+GOy/fKMPcMNDA1E0OwiN4DzZsXmbxgORDTm7Nd/OMEqOKHS3GHRw/qyYg9YZa
lmHBTUA8fwTBuUTAquuaMMsjhWenblqalvhyF1cQ9zZN295XS0/FFV7eZ9GdvC7m
bXJMWjjkq0Qn6uDTaMmdLA7ug3gMMSPCxOJcqe7whWM6A8RyVfx+XE7Hm/ynrmh5
VRhcJylkelggJYNdmqYJJbsgMrcVvwolrcgrsYFSPSoezQj96FjAnxe3IFzdyGPp
SFiuohNSfE0XUIG8qt/FpmCV9ghu2D2XqfgwahbL4b8cGHUcfRsHM9FC2NcYEEsR
2aZWCWXVWt4YHjkoqj/HzGyJ9wBi3+c+kN6rN/hUamJeHOgrcNF2EKdoxZW5mpR3
J3qxKtqdnHA5vmXtNByOPX9vPYWJ+UC99n4vD5+YZk9BEBzIW28vVY602zVk+R/S
D9w7nXTaXOqv+0j13nFbvfe3WkHL/D45EySvKcsHs7XBSsXEsK+O8THgrudYdfJU
mXz8MZInxCBxdADxJ8C2r/OL2s/lkRvhKS4bLf2Ck2qrL5ZaHtpL5zsaEgZXM9pD
+jzN6jEUh/Gj0Xl6p3858AdeL6BSpMnruYYF6Hz/m6Xivuz3nCatvKoaQ5H5hnyR
xzvUWr0879/5S9U81MVhC4Bq1vxk2k8SHlTQYjamBnrNpxxcC6blPPpc7UpGgiwP
YNKG3QzorovbNbTCn1coYVmPz1bbyb4KifyeZA09PQ8kraWhvik0gR/40uW83QkY
6rpDhBhEiqsD3CWrY44vAly7SpqNpVXGIqEdLb0a2JLSHDaYvULL8iB5MGqK3PG8
M2EnH9vdb2zha9MD5ViQb3A+cFUlxK+TZ9nytOCZNptQ78cTXKRWMOMp8zOpzky6
VZ0HVk3f2Ux922kskuFLqfbDaL3IsRKMvl7SwiFjpLYoMeaVaMnqhfgB96dEqrH5
RimhY6u20aPwXumnmHRF6fjrayiNye59bDmWgr0jhk9dBX7/osw1qroKV9l9dQ37
3mQjJ22K3y/2CjqnJemFt5JG95JRiNlGTGeGWpHeg+vLtxKaETyV48paHdGz/pEP
ynYYkA3n1caHDmmbJLq6ky/lHE19lqGThnw83PHwOxUJklVnqLe819JrA7z3jf7m
TxtVWzrv+mI2YJ5nC7oWvTVR0ZH7/gr7vfOaRJ6TycUViRxAq3FPNv2wLgFrRFtZ
UV8kmG72PFPt/JgLbWiW1OOcKcfeS7y/ifCjtEW6dBxzvlxazV8T4B51JduY5Xj0
jYgAm+YUnMwTwQsgY/QBwIQf9d6apeeMjUCmJYBchr2Mo8nF6CX/3cHAwCi4LsdC
kWcvs4f0G6KjpkSNbNKjaf7LdmeeMVqKsJKmQAP3Hf0porSDRG2ikBmkXiCTLhRv
jNs0zb9Byp6t7TUksC1Z8cpdZXMyR70TqlU32NN8Ta2CLEVNfCtybX5J0dAF4Ygy
ht0fxVo36mujmfFUmKcMYJhBHyAZ/E6ObS04V/sMEvQAJiG2roxkWMqxeYgMrlTd
+Awz0qEhyfnlilAnetY9mMTNx438ZVXEqchZVuYSr6/NpnVQtDmWjvQaD09plVNH
a/i/h2ZGPkAA+oGZDDRS8aDkJcBn8lx0r2Q6IK/WUWTh52HSAarAdejowrHiu6U+
4fFCZRHQMahGpS20rtj6yaHFYOXod2TVragoam7SuR6Q++tNHEziPgaVDDbbXU3c
7KDDpiztp4w5xwdUB4jjcXhwPVxwEoQ2CSuBcRLXvFmc3ZOvuYeRYxoReUMkSiXu
qZqTEp7uTBP5EZoySPGURT67xg6wUOxaODa2PjhcGC25U7YPd/B9ilXe1jRolqlL
x2mk/FW7iacZZ4GmMSuYyF6UPr27BZfWxaH4EJEp+l/+1NkP1gsFyjCophMqgKep
/pTaqP736v5dAJ5r+OFLX2/cbqlhXT/epSWImJWZFmI4LvDO1I6xJwyOr2Ds/HAj
8Fl1FmMDQwJCQgprMPu5SPf1L+fEsnKtx3BQbB47lL5L070mc2viNfPhu+uNdt6D
Vx9+SkA3SQlUBdHYmcsJ7BXekHRFqGXrBINLLnqSTAskTNjGGnfWd++QlAN6lWMt
gRQf4NI1/f7xSX0moF+dpdE8H8MvRHFrjM1Nsb3dAPpETEuCYD0JPcidyXHwbhCp
7gW565dLGskINIyBJ85WUjOoYmW1dYBWBiusvk2NnkhEoZ41iF5LudDaAapWtVD/
3JgVPJ/UvRLq7lxlMG9W1MIJ66SMf5Vz1rRGr6aryQYofkeLErFFAY0SYl7MOiGe
fRiKi6N4tbxnEO2tMj8ybRC/T3+feWdRlKGJvul2yteOGF/MIykebq51Ww/d4rWj
vVkbV5hleieNFPMzJET6uKzI6DsaP/bYhwTUqdt76ey2PAjnnJiHwog7XBGPlIQA
pp3n0iXyKQfVlYh4iijBBdRECczpdnpsKZandxfPv7nGd5vYKWpWM11GEbGPvg89
wih1ErpSdWcJNWIAvsYk2/7xuplXMnKyrpgRahFMcdgVmgB5zI1Dbrd/HKDaEAkb
6LOXvZiQwfGdrw4FUDJaJYwefykDTKCORsjjVP8NfP7VdlTgXrUnC/f3AZ77adqp
3QXgQ/esbhhfuqqRZp/Vra+/4HLlsIrWY/5Ik2qmfsVL38r8INsjsCdQRg1M0QnO
hypIc+6OTMU1V+ds1yyjX8XqEH6LRy/E/EY/7/X2Q+xIxR3q31+pze+2U//nl7Yw
FK5X3MI8SR06doL5t4YzHRLUG9FOxkbQLAVXOD3p47JJMVK/2x7sfjbTnMZg+1Zn
90UIleBzJP6UVz2hfcfmXTCiAzhPQCeX/EYcoantd3JGeX83HA/QO8Qe+hA6h0so
eK3CdQODzWRYr+ggJmASP7ex31KlZuliVoIbu5hbU4WzF2DmkjxetYfNTPGLrELb
i1ATUPEvu8zgv2dbNZ651qIjFTUmzzk+uSMJLmY7lVzlkj51l167eLL1n27p1FxM
1BNwR3l8IO4GRWMDuasOhAihaGH75M3UBeFJSEX20ZfEDTqE8O9AT5SEQAWTgCuD
JKvfbh85pAfyjidWTcCIRGuPua4WhhSC4e/OMl0LtyVhKGXcvHWWRwfN2+xtn8bJ
xndK68y0DKjluOoF8HbCWADyf0LmgvwSEeKSJknDlT6oeu7o32ncKVid3uA4ae4+
T3XxAimanQCPHWHdlmpWSXK9gQIa7OhNNd/iZRsFl9fLZeYMptM2UW6Q91GrWSir
Y0slnJO2bc1bt0v+5sSPTdZkSAOWVzL046YTe0FeFEGM/WbIhPPifboy4iPUnFld
pVSxAd27fawQUZ2gqkPuH/XnWU2JYi3bvGmyq6ryzKiLFs9AOOVdanGdwc2WBC9r
kpV77Pz7j0Ofx8mOY1yV0T6/r+3tylPH6SOUAaGEuUJroiGhQUDITLJHTWz7gBuj
OkH8pHCQ4jV9DDXiNyWg/Uzysrt9bE3Opp9D700t91Y3HY60nR/Wn7d0pqTgj5ic
hCXfZmNorb3fTR5euNi88htNJZ6QpWcd176EPE1GQGMratXN28QgLVRO8oIxyOFs
NNJtRoSTP4wG1jFYYodqqQfQNjZJU4QJ5KW0i3nbjPSm0RVTvSsQbCngc7GYyFpM
nZKWbsT7x34FNKmwdKB9qlbHTw9qq3BOeOww+MuX8g1XwdpST3pqNeyK4SjLfGVV
fNqi73c5vm4LfrnWw9c3+emF8zWKjbfpWW9A+B7SeQz7bOcf7oyTx4/ffG0sVDIA
wnkrLryi2AHSCHYwD38HpODLi7cnl6ogEcdGTY/sQ/YDkK/6dRky8/ooQrI3KB3c
Jxrd/OVnRL0b8K/61+bvQ5sH/pJbS843q6Nz1f+c2Z5F6qW0F7uNv9Utz7G60E8d
3E4bzmgbWahLhF9WhpuL/uPsNxQbLgYdJtE9KT7nm+dlJbcDMWF2ZtO0CEBqM6Mz
8ZqBIRFn3cRh8GtAmkUPsHBkB0hTqDzUTn9cmknDM6jXyzczYGsNviCwKAOb3PJS
NabMRM/9pMgKgxxbJWy0Oa2QqdyKDSQBgaq9bmdAdvwDyHU/thUDCCd3t310eKGQ
70jCxA/sBuoFmyV6NL3GJlsneIuBlN8GqZk1ifqJ9je3eZDC5i6sIjFqPBXVq7nX
TB4Mf8I1tD9sBFFWoz3xuHDoUMUfhcBHqJwgjDWsZMTyxTyzotYL/hPg9U3yxf+M
WYzmiuVl3SRL6bBgXTEjTfaBbHvcqvdlWDKklC9pfsenlinSmYFWd5qP4f/Xw1E4
rHqJm/pzM4g8jFg5wll8jVqHugK6ilYTABUXWoOCyKK1v9HJXiKwp7JJn6GuzD7V
OsJXTe1BfXIZB/0N3G2oMpgnx0HU7bjY8Yn8DzieofRUwhRZ21rjcbLo6VY7Kow1
8fVJuusdAZEzTuQ/P2/9Mf+iXXEnEO1toexEGAGgJCa9rLzgdyfv43qxmSxmZ8AZ
NaTkj2Mm1SinHAE84RTIbqMei4bbjf+j/SrUh6Iyhx/I3pmjkr7X+S6ceJElranp
zYzHTcjhgjrUTIkwhZk8Q+TQEomJaMDHDQ1IzJiRS5gzTy5a1eesK0ulFrHxhC3o
Zf4UfaYZrrdQdI7A0y6iBeIcQrleGee0eEmXnzkf/9Fj/2pd53JjhpDK28rEscgg
Cr4AHrLsyYuBsB0Efb5z0GaB/C7lKH6skwKOK0mJDPSsZA4LHMmpFIXyT9XfDtmK
Ykvsl0NW3lSfCSvt/5hBxIjvUkgtAtqCUu6AJI3NFCZ4u2AEEq+4Xp7U8WNzjbZE
ajAjdPThcVxF42VoeBvEo1idYFdYAQk/kS48Ogcho2C8G6LnrhcMeo83b3In22eV
WS4h7ocQ48Q9lk/7FRZw+sfM7OLsol49884uRVO7+vnFwqkmeQLpRnQRCbCZXoy3
VGoAjDdhiQoY4DcWHq57f0VqqBO8Xny1IONqtglUpc/d87XCTaUb3QbjNOOYZU2H
aAexDhFMPOKWClKswBMFreClyirQDRxbOsiD+SjFlz5cdFEB9Kwy1IGayC/xelnw
p7ZIYpMt9DJf3CB5vduEp1wCb0lVpmMfFF0iyWl4bvGSxfoLXCp5l6u6qi6ZFvvk
Xl8+M/FegQPws1pV8AMO3TuV28YdsrZURcb9YFB/5h91HLRJcnS/9Aoq9UgiybwT
wuwRpPWnYZxzGgPIU+JWbhRXtlX7mWuqFCKgbYbaIDBe4peKyluwKT8NUeN6Q0Kh
Tk0CwFi2prgVpuqHX8pw/JEagh94dGSio/RVvUDrFNzigG6RwQ1d3MPDdcrUuhXL
s03QzgJFxDH6XZkG2VyLvHZjLzQW+AOltB06n6sJeuqCTUXo9dY6HimZKGQOpcxB
unZqXtv6S5xi9boRfCmU5ZCMmwQGTgV63NoIB3Lo/8QnCi5tS3uetmC6jQPrgXP1
3HC9Cr0lTR2pMHzu2KIUBVs+XpDe8vPMzsoOsbDjuutn8ElunCjvFWZ3QPLSbdpg
z+as82K0uySqJz/jZRq+9HMdD56UFOuiKtWwc6nA56Czduj/C/d+u77EW3IZHN2S
nWdaJ5Lp9unqfy4RpYf4n7/B+R6VSx8faK23pV5v9LUtj1fJKRBKEFaQCSHVS3z2
7ftM5QLyawAPLK5rjCQCQ/IVvbVmwecCP8gtxkVNgTMkUtOHv+uIvOJFGlCcamtl
aX79PozWpfQkMNZ2GszjhZq+omsE9zKmIs2UgtO3alu5P8VtXhQEX+Y32YcknK3B
yQM3REK2/d7Oba+o6I0l48RbiqgGB9AIk7l12ceEx/LalYTRTaQSztt0GJyt/jas
Zmm8SSjp1on/HG3R0BJiDCyowzKuc4NGSXxlB8bm0b6gmOoN81bsPhMwkQ3r6CRw
1Gmic06E0lxHmknux/y9Sflzx5oyNbJhxf7qb7gS2HqNS7mjNe/J017rx/hITRGc
e5Zza1jd7iuigNmMiRgFJBsb6TXH/OPFvAkhn7yO1MSaBJ8cXNeT9kMc3poB2S/w
cVIvZoWrEN0+lCW2CPPl9PG9SU5omd+7jWkq9OSKgGwJHCNHciBsiooHjULn7C7L
9k6X/gFTRw5RVdKZH2wPoXeGWagg7rokbE15DSy7JXJN+Dr1Y5yrP9w0pjkv5/G2
lTRGFO571p63mZ+y1UDPTlIFsYBaj7wjucxydH7okU8zp4kPo11KuBkHHdqq8ZvC
xHsnVn+g3mM/wL3hDiN6J2mNfuS0G7rQtBdR3y0uRNSP8hLHSsAm1O/nOgS4YFwn
yvbWyRIbV0vGv3vZVm2HiAiwH3wYLdgipKPHcEzBCw4qvWC/KC+e+fT1lovbf5Y3
NZ5UeR3FltdLlUvaPUHKfKZGA6G1aAP9e54TtuLIZh3tBDaj6dYgvNkIZXV+s5tF
vK6xL6J3YD1iRdCj5dsjO+zbSyhyzCBgS1xIJ/U4JZ8g9AjnyGkqKFF7onrkLxLw
nh4utGmXV+LvaDhXaYG49PeMqS3ar7qPyBt9oWTPdDG/jBVRgCpzWN9qpPcFjWgE
/yr5lmH3pX0987u/9sezD5q/XH1udqS3WFCL64tT4fIoU0mojXMoA/s7qr8WWIyS
vBnDEErTlQm75LbvPYPeom2y13s9o3TF8hVo/WQX5eg+x+FLD/dKd2dRyLnMgvc/
CtvZR7q0cFZ7KPUa0LrerJ1bZ05UQpipaV0ztl8ofx8p6uZn4kG3xqx9ak4I3yxa
usfb+KffaL65IHHUiRgVzsH2pIKH9irOmvdlThu7luFT6brAhAHgmmhIaFzbxJcc
UDNx4IoqfJw9g7vBCT9tIfnp0wDYAJuGnXAYPHcHIx6oOYJc6PkQXIRQLZv6EYfw
o2pgA8ET0vRf3GEWYQu5WNZ5jkktldQ8ImixuvTPyFpYaOoPM6YvvIvitoen6oHQ
0QlFyM2ulJyP7ed1KfCgPwPk/d+I/otYXRRntKBtyeBdr57A4qhRnw5hWn96k8py
1sfQTGFvvyEL6d+nAzfIsyxVWqSuVEAigXWfrmKI68pvozAh/ghBRoI2K/2T55HP
kDpNTtA+9ImBc1LtIqgc4zNBTqC/iSrgSpViC74+fVtb2D0SoOGxcuboRT2V5owe
6FANlmYuPpMMH0qnk20TphZkO9OUyTKJvmYtuwpFhx3JkpB67zSQDmcjpj2UtbY1
abgm+eKwoWSqhIzYrn8tW1H71BtI3nVMbR5Vz8tgU9Y0KAQ6B03QWkLduA3cs05Z
NZJUwpmk59YWA4+lMSEWjfMSzKnnHFEw2pTNPQ6PpcOkD371YkW2vb/+iM8bN64X
M8egZvPXItHAHOR+KBW2oVXeVTVQbsI91rr0PpbelQx5MuXsdeQx2SPsfuYZ4Peb
OUDc5ZcKmgLTfVWt81m1fiDonCw8Z2GeFcuYoT1ZWp0oO2HrDzUTSdDYADqU1a2e
/i17y24Ie/Jem3u+5nWmiVn8z8KcHLthkU4RiDLZcA/abaOzPni5f2H6/ls6kzxv
QNCthL5+qtsUz08UqLpYNL+qowdAB3qf9ROMC2hqgmC5RKIguOVB+ZAXmM6yLTR0
G2Q9c/gYTAtu7SkC7IdUqaOxKLfCd+e11SDS4muNP6o+xtYz/1ikQal+3eQ/2BEg
Ia+ooRbnVldsDdHoSCtEtFrVLmyj5OiawEf9lNa4ZhKZzjmWOjp0P6e0syuO8Niz
EG/QiEpZApNghHFH7qfKZGuNEHa1Edc5KJOxrgSvTVV1RICRWqXWYevSocr2K0ne
xqu4pZbAsvqEn3kspaJA1gHY4TOOys4entRFMCkPma27q3BBrKnGnjNWy+7aKt2a
PmOGwwOIDUe9BB5/AAGWszoEfpEaEBbetYlyLDT9UbedgMkplCTfCby+8dgp/N8P
5mA7AYx7L5bDsP1fHpLRPxuzUmxyjGoSWVxWiuGob0c2iKdd5NyNFQDZGdPRe4au
eAeBwRICULv/M4PAbOPgRM7xIiNHxyxgc6QaPL3vH81dWMSdK27pLiqOdGiitvQ9
FewwS3dZwL6NF23SG5FKqXuIq1Y1QhVt2Tz3B2sD5pnsCUqSdzPfjOEdko5BaYoL
tVjSgKH954PmlLhkjkOC8PhF+gyRMm3qYd0Lq91JoQT807b+xsxU23ttQhydpQ33
9XLv0A2sle1JGRduDcXXo1i295d/TgOkhvQkGDa2dZEaABUFc7BBs3A97E2k9nMo
KBnX5IlkYyoDOzmhLZgyK4b3m9oX8v3LZlT2bFL02C/elKQm+yzJu9Cd+miFbI8s
QqOmVOP3DMNXLM2mkdKCBrg6uaJw64HSoOG4GTO6YQ49tl8D0KXnNnWdLlUPdP30
Bi2/mZGssyuU8NSZz8rrxRR3wNVv6Yo7U7Qu5Sq3NDml1JLcbCHBa7LuPM6IFaDt
ElP6ZTzk6crfrYedOB87fKU8YfkQ3AUZoei2HuWH5DSMm8/X7ZpYRPX7DGhu0cSc
LvQchSdMXMGUsS/a2KgitB812ppZ42HddCD71Vg34chL3YKsDf/WfDQmNRE+Hkg8
fNnMW++s9HSNur8VuWRuVLODBkV+bNVy08txLj6vPDFrh3q93JMQTre4vWSlhbZE
4Fr5j9DM98VI13mEYkhSJNyHxx+Tjzj8z+H2P/lJQE55mdPzoO8SoIibSfGVwjpU
1qWTitihf/QvDlIiyk3EwpH0fjDKeL13/1G2kBcP9xH2TdJL3nJAmrMo+WWnoBKc
NjJ0VpQ8de3/MbZfggpz5BB7wztK3z6WXp4UutO43YcWVuWYdZbQUW7heJ45Hcdh
O04ah+L2t1Lf5Z2QF9kVS7W8Mb++oQ8LWxP9sK8zvIyC7Y/kikvTL70xNXAsGrhO
0AjcMJJfCuSvsW8D2FWiR+bvQjR3o5MpKsD/CYi77S9+2wttXVrdBe+0V+O3A7z4
LLRj2PdKHX58leAYsjow4/fOBMelXFMho0jON++EKOitY2yVVUBLAUwEhslYVyiq
5QrmWLyrXtTU3OXXgifkkcte/Ho0jsFf3NEsA0hAffQ2DaWnEGdJc4zcSjW9R6dr
vJntqAi4Kn421cfWwwsoiVI+4n6VATMSCmgxEzd75hntsaZ2hTMIMIolfWnQlUn6
PoeBjpqX/PjjG077x5ZukYM1XDRPkzLX6xQnAqB3H96zhbC8cwQW5jpwWO+qR5Tp
Fk3jkq275q9Hb7ncSx3XThKvAM0DmDP7XWUbr5PrkYA1Z1xcl88NAP31ICC/D+S3
jQ2wP0MVXWgAloiuL+QG3Ot+BcdgGUKVcQODyyvG3RwGqmLaMjjA2yY5xAjetfl3
NcDHzROISuPQ8AS2eWRSOiBSVDS3T6J6ndXCo0yFpERH3yKHYEl+JWGpAbMAnDqz
aeUzYdKitTjyxFoISjjYdobImhm06/d0Cxkqb/to7aVLyH+/5OCRLhG/tTYMwGqb
6lt7vJPFB1Fmh6Zpu5O+x27vNMONqOeIU9sEAy/bCoM8vGeDncc93G/KMdmc6y5g
Wwbv0h3j5QPvNVJnG33+tK6QrIdVVHGBXw1FyT2Fn0wCo9DmCTzWgqqPO4VyiJ08
YK7qcL9Yl73qgVQRZI/57HzaauIM7yF2zfnRn/7/hZ8JOyiJgvvAuAhChpVy6OXB
9AiKwzfBoMnumHupkTSa96tP+mtjbFyb4eLvvXDCLr4w9YV6eb6Yo6v/ArVguoxR
nucvLpy7FLyU4cKPW+zXy+6KU8AZJ31hpBe3fNE1QFAk626jchoAd8oNfNJGr1DC
QEcywqrYfbtdQwEhwu+BZuTd8r7U9wVOkGjJFXwc4dsCYRZaLBeTEla9eW1lfVYe
7Gfr4HX3Ic4Qtw7sejcVEv0G+y04Qp17uuEU38+FI/OTP+0POROZSRYtYcnClKdK
9oyTjS9AKEbuo4bPqVHqa0Ei0z0PbM3p8+H7P70x60Ld9e7xUWyBvS5Dszf+CMLJ
7T5h7PeHTdJXikC9TW4eHCWSUcTW0xCkC6nWEWZw2VBaauMdfMjtWz++/Ya5O4Ip
YUCr4OdRPLUPhqIxabddj6+47LqLmTfOUbLCUfgdFLLKRxngSEMKHGfrpmB7KLU/
q+V3Sv+4G3kPCUm+US3OqJpI7F/2SkumrkDL4apqM1uZKZcrudZ6mgjO6Jom1lvk
S8row6KtDlgqXJdqJlj3KxvRclKyBJHiQa3oPtrHfTDvpT8h+5FCgR+8dE6jxbwK
+zoYuSkwyQNJtIaWcUuMnMb/WBCdARB1uU1HbM7/iF7FP4W9pGK+QYtlTMtJRETv
T7b0+WZQrCZ4t/Don1T5qSO3mvdbQnUTnMtaElDfeun14NrNdDehJB02vD6EQ03k
TjK7uhtbO4z5Vv5c/ByFN7TQ76X9q3id2E7R83t2eOR5acXLJTQk0+0MiYOPGp0l
9SwaAeCYSlxsSDJRNdnijW/XJUWguy+3w4EXCacy33X0MNtxuZ+iwx2p3r67Dji2
yFOY25/ff6xyOBQx9D429UoHHyo2SUOQ4f8MdT69UNTspfiY+4eyoWLff52siUrf
Tr1LKVqd8GNl3Xuik47pw3eA2ySkH1P4maDWbiXuRf86rlhr9WeonIpynbv996Np
ECix2YwsPJosqpjv7ag5t5WgzbAb+TthtJXvHnNeV8NwE4SfN0FwzIj2YsyDFA1V
m6ijZxIWibqW26dmvT1x1X+ZCE8RKyC6awe+H7E5Zj0Ed9ty7cYaXDe7NG05K6Nt
0o+2plHfFU/mqinM7ASOPFC1tqaK0aTXxASe7O++t981w4AK9KdxSD2/EBklOYMk
+/xsK1AU1jL0Bd9sYyDIVo7NBY3t4jDjzRRuF2yCzQ1dYc94++ATgL3KIipZ27Ff
MXJ56V4fGXr2v2IHfEpHid4opZ2zStloEog09otd+/S59Gd8TXgtoTK/lHExLhUF
INxM61t0Sm1mmLZBxGPC7emNOO1nk/tYQHmKazKji3v13RiqqGH9yAUO57R3oqxV
puQsilU2n83NzFEO0vddZke7D792uzsKbpMHVYSPEcHD7uHrToRJ6GfXobG02nHJ
gpb6RS3H6BaE+EZK8NvkFIY3GA9HDtvXjhgvNJQ0nsc0iiB8olgLSvkA5S0A0AAc
75b3wz6tzNCfGK9Q/XozFJjgMn435RbvfPQkJIBSOu1Mlnlxe112CGrhLY3D5NNy
Bk1DjvB00W3Xoh52n9DOT4qjsWs8iE4LjnPh2Q6lY3hBO/WYtmQdjB4QAU77dZxU
ObZGFneofjdw+RvB0XgizGdUcUZaeVZY1bK4njKAlE6bJ8kFPcZojVxzQ6Yimjkm
qXTqJrhzNcLHHB7oALLXFIJVqKEOmeWPCQzPyuhi3yBtuAFRBJjKBaUGtM3+R6HD
2AVTpo7ADDo9Fv8CmDao9/H0p2oYEJxFpwZPemoyt64x2vxeV0ySQm9JUUVVVHrm
O6wrUHWBJ3CxX5tDmyUn9Q4vN3zr6ZCZvDsCxDMdWvQArBNJrA10rteDSOnczedY
Ce6aLAgMz1v6B6n6I+RoZCIixZqExW2Jq12gqMv9Rf7Atrg8SeEmmYg2kskOALFy
Y41oR6buFXqq3Y0bL2bWyKgcoDvnmqynrVYyDyE4Q7BPOJhrCX39/Byk6F3prTjb
3/IAKMyU7097ioTjwHGMJ0/K05mpiPM9UXNl2wObGX7RHgb9UC5zWsAId8yBJzad
KTCVkp5AZoOEwy9E0Kwk9S/uLx1U2Ik99pSeLbLPNHbj8riVGLkTkmgrwX9sJTHQ
Yqqlr75wrZRIq3D1D+rtC9QvQFwWts/+tXK5yX4PqkoVWO3THjc9gnsATuc4Y5N4
RKm9fEbmq4w8580fo5cznKKjEEVn2HbIWcGl6F22AveJjjql/lfGQLupBHtSTnQH
A/LjFrmQwMu9qFB60WrtJHqIhGJGRslC+UToV5ZPRsasYwRoGZu/DN5qsITuFsbo
EwCgryNpZb6EuBrWCoPK+w6panJJXS2saLDZt9AtjGVyVCCxl2IW04SjneS7TJi3
cGJXrxXtLMiCJKdOcRP8QeAwil0yx9xHiIIxF66Vhjyag0pTXiPRzaHGSNIBa4WX
Rh3gORfcZbsMrAz+oOXH8mkr0eQ8YiOQ5tMNyaj4RQlHE2Fpa4ZqD76ediN1p3G9
Bl4GuGsx0gXCpFqNmbsrJ6SDxcX2EpyWaioOXAU7r3uKDHJA5rYxOqdHjRq/qVA/
emimtRu19Wye4Vkxi8u0ZBjyG2VdqGv0q+MZaZvO0wc/P3m6Bm8xutWxsoU4231W
8NrNhrc9Zok9BG8F0ocGjRdBNuH3H2C2HI8V/T2kRopBW0LuLKZfxV3jI9cXRBbX
svkTWU2RsGI6+x6lMYg8FHVV6ifmi35GMBbH26U9jE+OSedpgNwGxKZywZvW1+x3
WAqxlo/YLrNVEE6qWbsfNoj/5v60XyDH6C5oM6eTpI0giRn5t8vKdQtB93oTapjP
/vkIVnQcqQAJ8bn/gbk99sU85YguvCnULLLlwhXquY5R1ag/Z7n1NSwgd40TtOE6
nZvq0eti7XyLdf8racIizWl3OhXlJ+Ne+qWLxDf3LEueJvdOUblP1DY538FA80iP
J9CaCDuEDovhYJ7teQOsuL/351hE39T+mTH5/nXF1N7QpvF4PeK/umHP+qpSiizT
AvjjvB1jduHOSEXiELe0q2OH3orp9RQl2ejPs6eFOnbD7b6pHF3mLvPvnpT8Hu8k
1SE8Oe6mQLBxgIi+WOCNcOchBivAdDz4Hr+Mtw2zhsCQFpLbu22n4ieXG7rdd49b
G731eBWfsGfslTXU1RSIV79kRZ+34bOv1lBW0PFqlC482k1d45b1r55GXbSk6hrm
NSNUEg2Qc6plf53Zo9EAsxOxFKJbC886sGTxVKuxCx7h4gBKH+1It+itGOPqt7Qt
5S251mHXyWsa8BJt9/tCnNJJ3NhH1CjA81JPTIwLkreG6axeIoUZ/iCCyqxTrTzP
YyLEF3HkeMRSSKxRVOVq9PPQ9k7VFLZ3n2TdMg/DF3Yg5/x0cK7P8EcupqhRNndA
uD2u0SIdUqSs1VI1sdueGmUM4NY2EZjd8Cs+egtSlDlFcd0BBw1z0mGndqEsb/IP
pcdU3Cw606WUaAO7HeYKm5LDGVeR+TIQnPvzSxj3qaORj95ClZP7vg/KUyBhn2gU
+Fp+iPylGOvKfnD94XMDV5lnOdlqTRmAYY+8E4MxLsQk+gOjLGqRK7Mj68gDTCus
fknHrMjG1jHPwjeGl3yyBYjug0ubbT1VuSFhKFMJXdFkaJx3HJesDY+BRR3ERSej
VH1PWNlnd50lmcEwPCm0aZpnKkHnianZNkOvpnEi47vLuwEwt90Rwr3m/2K8Kunp
ipQ8C7sxkZ9OheRL5DEFKHAJNdolLigRNIIFI0s66XUcpdRVvViAuubKEdBEY+yQ
5oKjzkGhLApmIXOpmyll5H8CEb0grl/4fBChzuYTshyD6JDnozafS//IfmWX3uSF
RYtgd8J/5/YtQKl9JpQ+vRPGI2gLD3KVty5a5WcaNHct/1nvbsnbgO02L+9oy3PF
xgvlJmtxnXQVX37NaDGcZETBfA8HDg+Ov2/Y2Pp2MaqcWYXtBzCDwkTBUMsfOWT8
/yn9ir0RVTxnr3fMatvF9pobIypSO+Wr28WnQIHR9bT+KSTVYfL6m2tXPcVZyodX
pf3ERnHBfzYWgmu/nTpmGYKCfATS2SdGRVIycFkO1abjoYrQtrJCLQfh8b9b1gcd
xL5aDeS7O/5ZvzTKfxK1BMbwuGNwyJNsJICoF0n0ZmFGjwStaVb+1VIrtSp7A8Ay
1CnpKSYAWs/3+j5S8EbHe9uqRCqbv5GFrT9SnIF9bcItemwemEPw+fnuKEaRJyCd
/A1cEaA/2njyc0+O9BE4AXMju/IqOqL6SZuWQh9AJqeNsEe+fpChaRpIj/gvsxD2
kaHkrwWhog/BdDN+9tvg6ojYzliFIbW+vwu9o2pGlXifGhNMe4y0+CmNkRL1SkhC
7I16eBxX0axfMjn5A26Ig0A+9tVt0qwJpsS9aM1uSB3ZLpOxTn6NF37xlcq4MJ+z
gtT1r8jBexQJyp1igIcpEz8GQ7b+7wf3xFUB3s/FXNx0E9Bq/QbMKdEM4vZVRhNT
4d+cvU/XcbWvrzfnFKgcaH3IdlxPNYHyKH2a4EZmDpVJRC4pDctnON+OPbFG0ek8
GXXBVdLiKiaGPAG3+88vd/u31/Ohnfm7JRyEoK/JdUnYu2klxCqPlxcjN40LVAjP
MMhLxoUMVXgEd8UugBZg3vkjl01CwLfWRvf55L0EsASN1Yj8U8dIYBT2bJ7RhwwJ
eDO86jLz9zu6aEujLNeOZ1vp0U0sbUWoz9NbsdUfH2xeCTNfnFk7hZ+uVSX5CU1M
12T0BoAE4x+9DtQm3XoOgI73XcteA6rPpkwRepjNFgEVVOGoscQY8pAyoKXV783o
lzv/Ew77ITthlT/3wpOq/DM3nj+PR3xQ9znIsg87+0oPBIcipEiZt4lXzSO3wFZq
OJ/FtBzL1X/7QBdSmdKfKqNGzpklheh2lcbyd0jt9OYnOEp7nubLLMEK+9dQ2N6B
5VkZ+8BNOZRcUgfDfg7neujfU+frJ6RNUu+R/LRf1wr4AkIBJ8j9L7e8+1dLythl
NURjpx+7Ct0/XnvY3HN9AO+n9JfpYvSdRjHv19dJjd60eJbYXFO3/PJtgW4W1IsT
76aX9jsE/wMEZTFoIWG/CSD0z8zLefp0tYqHCBPazsRtx/VLEBfzNcRsJHJao1gd
tuwLdywCs6hnm7OnpC/cqSHfH7ynfOMtC8Don+ZeZkPb62YWwBSwKoIb20rfG3CP
lz6/xbyTcQi6WjIou1dq/W8LJX6CPh3h4dFrl3FpPC4BU9mN2J+ePkuVgjfcP7GG
PUPYQdLJBmja6Mi0kEC0MfGIjDvNZkUSarGIaH4SxjjngatFJuG9ohKXIfo4UgTN
1LiaXBZUSOO0Wzha+opg277eCR1B6Ifm6k5jgxI0v0xjBxycbQvWOE/6H0bYGHyU
BHvIdVg7m7/CNzYbn87FvUzHMYTuiIimE+mxrTdDVucIhn59LLDzYU0HvftpJvwp
4JosTAMRdxbC8Dx6j6JFnGs6VRuCkEo4HpULyiQYVPetFgPGLdJVx8XVz4NdklnH
r5Xg+i0w4jK7dT+M3F0NhqAgzgHt0e07UXPsFxlNsOfC6GwpgBkPtUiXMAO0XxFq
FH531dX/ErnSTmOKVnHEtKb4XBrPgBOUikLVXWhV1jkVsk8fPzUV69bvBGiE846D
fVf8wjjDOPPdmYbFs4PkMG8e+j0pARZxdaGk0Hg56kjglUSiiLL62bLS6l+bb1Nl
Zafcgx0aJ6HH/vv7tS+B00U6Sj9wlNOx+1r9/wbTt01q+hlk5fr7nKj8RDHokQUO
rWba7uERazLp6nCkCq/1yyqv6mYyzaKru6ITir/beh18sLcOEoeMvtMIJbNCeEvz
CusdDFnl26+r1SZsZ+ZCTG2T97SK53gs2Tk0npE3hzYoLgFYnuYHLxCAJgxTZO06
0ayJAkKrJcX+Dt2HkDE4zR1NwBEjfPIjf5xET8+Q8boa4oyvoIvWp2wyg3Pv6iu7
qxn+cZ9GoJmNpbPlwl7JYAhHhRdRYdgvXxjKKO/kwyYlyKWaRN6GRGJhyl1vUdw1
61KGXgJzXq0TkDHRnuC9FK+vryhbXCn+tdpUFSPD2gTXGsoLrz4BmJfuvr/tmUCG
NzL7Iow5PH/HICq5yx1LNFcTSepEvHX8KRrG1bPd4JLSl3bDxF6fUTdHoHA75sX8
HvrjpItWUKIgHSRGz4ebgRbs6aMhngWOFz3/NW67Jy+4m4H02Sa60eiwpw/fWb1b
dtAqT97W0LIVLC4rVAmY7r7cW+Pm7BNe+hdehAR8mAaZBj+guznpIhYYPMgqFbxW
fAF3sXTWtowWS04PnMGy61t0ZOdd/r+p2WwP2xlMCcKTXINGMKnn89czAktPcJ6h
hQW9gy7kzuIkqPRNdkbkm/qQiM4TNu+6TqPr8bFfdpWhjtaI47gS2caV7AJ7BSbl
/2svvA52ueSQ1PXGt0JfprLpOkN+1YJ4I4FD7VH970tociwNyiN6X1Db3tH/mo00
/ts1Bti2zPQD+lZG1ItKwLHLEq3+14MymXBGI+8cJktFFSLBoICcyLMDn9pP1QXh
rV9XVoNHWGyFzqe1WHL/fnq7ELOZW0Jk8dDe8EggDRojgcI+Iski9wwhlBfOF5W2
wwV1kfPSnqqu9BgLTfY/IL/UiA6MLarVujlQLQPt04aFujOjnS+SWk4L8PlWLKe1
zdWZzfWJntO0t3VBU5EAau/8aZFbUT4dj+d93oYHdTc7yPwXsUpm7IDyXKu1/vMT
bog9W0PNYWCEr7ZPQJBGUhdkXV4IWIfBYZ/2Sf9a6qE9fz/0jhOdoRlvfFb6GaZJ
YFqWcAnxzYPNNw2PMCuYd5grvl1Wk+dty9sdS8HspZJpN7vFfbSfF/0n+I4hYtQT
8Ph07KsaOlWXbytrZ/bJE4oPD65l8SzfA9MEzBIDREb+Mm/6X0UTa0SgX/a3hpkI
zybchind7lzGWk5skCmaCBtWARIoX3KBAodCkymZeVMyyiyGyVNqJMZYvkzboHod
z1Ky3rBftlhjPa+NSNxZgx7VJwoKnLpcyzlXdlWrCiiHjm9ZZ5eOUAL5127Ai7Ts
DtRQq+MH5SihmHpvD917VG6a9d7wFF5Ve6vJwDhP4GE46qItquAvzAA6DnS2FOvL
i+6sgKd91f+0NrjHWEmvnwaEf3dYacassyzW771HxV5zOTn3RM8Sv5a3zXu3boXM
Rbv4gILA/bMBeDMaITZNPSQtwyYTiSESsGTTroOwh4R7DTvQHVG8JUq7wL2TFim2
9IO+qB8GiJDrn7GDxHSNvQfnVJcMQSEi44ozTjNeJctEpnt2q2iiGO0467ZcbYlV
Q6pqdsBM0n0IyG3MElJf4d0Lhb7irpeGtai5eyJ2udbBH3IxPDNJaOR96ntroLV9
SeanvHaNBuuJfbpzpqwtV/jCJflpMkARHkcQtN2/LgeTYQXBpDYq2fQYaE2y8J6/
4j9p2bmI3QzH9cZ8D8C4BFi3zhTKT4/H/824pIFNCXdWufFLmyuKzbMGW5n1HN+v
FlMhRlpy4zMrV5ZADbqY3v4RK68N2tlp1zhoHZ6lRWordv/lEKYDuNBKN5yedLKJ
6RM1DMdrtkPoF8ExAbVjFZQXRS9+qmjPjByWbBsjODrzWQlrKBKGoBBI3hUpkVA2
jDMulGfmbL9A0rHK1U+7XMjtqETM11qj1Kki7VtFHMCQGQa3HFQxHmDVVwYeMD9K
iNm88r0pjTT9GXrp4q1qlwxOj3O4rbqraKzt7Yk2kRjJhTCO08fKk6kbpAgdhMR6
Yhhlm8zVPtHRHmdqE7ffw1a5sUC8xfAn4tryn1hey3TzezsJr1xXIDQH7qMy01Ge
ceb10r/r+wcpOp7e7Ac7S9/1LqKfjHaE40UqwrK0wBhE24stNWWujODzerXjDxY/
2wv8Kt+6d7yidx5iqAFqJNdXaDidsLxDJFTNb6xDID2Qk4E0Q6N8mwv4pHWio2D1
dKI9xEZvQQtor9c3OH+/BuNPpI1+3AJs6nsK5hsAPNPaZSdIzr43+90n82ZmlLEt
QbZsf5z7AsxBE0yS4RC5wotBG0HPFf4xCziYwJzBrqfCHJIpdRywGQfj4L2fkbnY
p/kV/zK9xmEbv7WotIXy1WFhsiLjQGVVLdO9se78TxBYHnYKZew0e7khle5j2H+p
6Ge/yucCZrZA0alUGJiW+t6ujvf8TTZCJbMIwRkYt387dV1eyM9AWIvDmvBoFMcw
Wey7IdFgtesJ2nQhUC4SmAIZY1hwsjc6QOLZZdFNWzFbWj5z6dA0XEwQW97Un6E3
vdEhDJ4VjobzWIRw5s/Ar01nPTj74bwHTLARWPVy1uoSlsU3CJ9L1cQKPE2Admab
/zD6YrdSh0iBXZq3EpeZtm7YP9o70+cuJmnZXaMmqz3hitarEx6dIto4yVRHW0SS
Ota3EfVFrpomqB9ehDHGud31Rxz6m2+YtE2hRL3OXr+BM/H4VcqVvzgfZMrtYHKn
AxVzUkaDZT/jGRZSaR7YMUvTS7bD9IZ2CbsoGvlV9q4k4Lg3pEiV7iMFkIc7NURK
yaY96+xt4bn7Wd75shCt1mgMSfRYWKIq4dv2K4HKd0KhFY2l7wY1XNIBNJn1LGSd
sfN9Zw6JOFZvs6YZzdqpjLCtoofj+vvGdFGlRaN3jO91jsyg0jERMJO7zrUpbPcI
5VzP4rmvCRj5BUIRdY4LyQIcKWVeCzYNxjEgVLR1/905GYf4nnY13MaMmAyxy8i3
yswIczd9WxLkeer+a9EAQ1X2x+8VmBir1ciWyvoTRLrCDJiIGtE84yPVI3B6DZXH
QT3Op2QJytx3lAGsH5dLerbSE90jEwFw+lscp4W/iuZ+LWUCnNJOYcYVlaGwPutH
/FByA+nn+cPy7YO9yo1DyrrGTwi7bDuLJ2qPcyd/svE3/vfVjnXz7CcUxB8F7/pL
J5Jg8OChRsG0lFtXA2UdEaMiUWhlKGqDKNiQf57WboQsD5T+4TQ5Zd8ZWLthATiP
r+m2A/Jsj4P0gQC8MrgNUtPVG38cGmxHMT6MJ74BUjhHBADEru4aczSL1hxE56Oz
Ig1mOeR3XI6TMlSxHL6jCeQpiFt1eBNoA2TOSbzb+/2qF1c8A8hQ8owYiRwterYq
VsgUNGQuBH1JrV8pctANlC5BsoY7Go5LMTcf7VL/BPZ9Uqp1YtALfjFYGfachoK4
tWTWs3MbjR/3KVyW2zcZv1jriBDpm6nfC71f/44qG3xnnh760UJqnUIdn8zUHeCW
R2C1gaOo0FEvRLl9G0/wE3g4E9tzkRAzE27J0/miWhnh+xXdRkrWGHy94g5FSitT
CHmg4Ck4vN1TLVQg8kBEiRNqGhyJeffRWH1gDDgSCYKPI0yXCDkj9CqiUC41QjXM
KUjfSiIegdG3WnTE+MVDW0WvA0PNa37+maYkm3PK3/XLEjfhvG3pfHPvFZkoZkcy
10PPpek1ft/DnINk5FrB9RSVoxc07h8q1p3CHLmbwuCJj/r7Ea3gWCmAodS//d9Y
bNKOJPCk+U9OHUm8mJwKHGFF8tx/fiPsVHLPbMlDXle+vxhL8WFESFhV3j1hU87m
9c3kcNA1mf1vZGYmZHk/pgt5h5kA1arY9ib3dFMPXRJvVKx8VenNZe5yPwVGKP2n
t52MHkYuf3crgDLBYeCFMwYx6asWnA0A9wsGHN1JzI98ZIXNGLQ7pVF2PlxeLXJi
SB+WC5MGq3BvackJJmWQkgMMZb9YYrRkBM1aQESJUMKobmX67/C1/wFgrl+JVzY/
1dD5HTv6dG/JEEA5mHGT+CHPf9LLyYmheUNyOLY5XHrbpN9qWlQ4pfzr1XiSdLqx
gYDx0ZfhZcb8FqrBdNOqF9gLVS85Ed6TBctVAnulEEsJE0iy0RkIzgioaLLAXyaE
EaBTiswtoqyXwzNL+0XAGXPwP+XYlhoX7yolkXZEFQXwkyVOfdV3wizWQD5OLTRZ
zdRpm0Htb7wh6EVNQcwv1SFxY1x1FiG/3BC9utoy/XnVMjmLS3hf3/bf5H8PWWhP
F2T289RGyEb2huqQyr/UW/4H6iXEyHRqNGurGWykG7C2+JpjD86VAX6dEX7NiHyV
CEWGv/Z/kQgDAOfkXH7PET6MFxnEzR8bvvq4LwfKHrOAtcXHhgGXICah6B3G//we
1Pj78u7jPmOoYWvm6E1NUqsqdtIu0/LSRR6qrTT8YWAXzDPLjB8l2zs1nm4Blz38
WiZrXuksSSB03BBUn3oROxssS4FYUBX1Lus+ZH7G45EtcLhUax+R8K69hw68ME8u
T6QjaU3ILQrYkBstbj9SmKPQx+o/IdIDw9i6LokGQv0X6b6SoRU7sviCPTz0zbFn
dSibKHNO+kIvg+4xotZ0qN4ININpZ7RJ2bZApicyiUrwdaJ8MCW1yH+Oq8ZGQ/xn
Dcq/9YJT4GODyyr7CPQCZ/9nJFsz+91EAXHGQgjcXWE5OUOrY5A+ojFNtYV9Zj2/
kuSLDyQFsu2cRVrgELrRv1X5GksBn32eQK7716MusARWXp4S8J3Ae4SGZbLru1Hd
1EtuObOC7ETOo03ga52gGoRkEMcI7kUKSue/HS+imTbUDxzCo+YOz4k23o31pWkn
8UE7uOwyqNSZbVjyCvMoDO/IDcQxRrSdd3tnLdCADLj9CmZvL/I3sgf9t2SplOsd
glImW5bZ5D5PcOsswR/Od7hpMuSS+9UCa/GHWj2l2lHhztvOdGU75n7/FIAt8j7j
xF474noD6TR34k8mBNiz0VW4k/vqyhPiPr29x5RnMoVus/ckMC8zo6Mq6jz1oG+V
Box8cHHOdAZQjon6te1JBBvq8wRnQZI248z2LuUueXcLQysoXROpzxK47k+3LB5f
V/K6TU84fajWeDwe8EwZkSYEYSoKzIVB8Q+Wm2tPtfkN+3KdVVpzjpMkGJTLL9X0
iZfEooo8XSgZ0BZsM+9zfHWNmZoRBpmpBrb5/Kg+GPXJDEv0CYYxunPmuWSbndhT
z+ULarTTKFUcKWMSP03PwurTZ0ODb1ysMI3i+yCrUQRL6pVQ4psBliWruXUnkRbh
AmECBJaJ9HKCfkUrJ23bk3+daKMUCmRJW2Nh/yA8rgEuqRWiTBHrcqJ1MjIHe9eL
oVDJqEJA+RqkZq2R74duq6LuOR7By/nETD/PEieI0eU2eILG03jT5QTHqaH2H1bn
pa91psCtW4Q+M50hgnmPAr0tzC+Hxx3J+5v2g5YD7iSXq2wluZUsURpRjCAJv35Z
VjAhMONh1/Hm2bfllkZNO0PqEnHctcVfKrCX6XitCJABDeIxFnV+bXgq5LPKbs62
ZNvv87Yd0pznDsIj8qDaf38zSXEgAhjFIkgIhkoPzI/Hb73W4JeWXRM9Xf2X35Bt
0MdCXVTLb1VFeOm/ssm1Fcd58QDYeYxDtfZu+RU8ZaU4N+Ongh63dV5cZGcAZ6kE
sHjKoQqWnyGy35uEufKI9SsLQ0f7tJ5lFaXY62o4OL82lrWFG09bO8dXaKOgTp34
eCi/95GHfkGM1wGEbWzDk/iA2aVBcDX0Vv0yelMjsCfgh9iSdw9s0RJCENKKQOuh
D6SFYTlMwFNKgG4OKYv1JMRPR9jD7PSNoBsb2ET+96RLT64KHjIn9P4Is+LWfZs4
C3aMll5qqE3VInLl5jBsitXjhf0eeX1j2Vwt3Mx5XgYyGBax2RKNuALqkLOLWYE8
/RSiNRpg4bVxhxAJwBH4Gek3zSDPigXd0NKdgvG+d2LaWw7Eag6InHbbhqDP3jqL
Gb5+HCyh0vWIkH3b3htj+M2+3u3nlX5l2u0ITb7gcpj7qrTwjd6kn+IixOdKT1ee
ucC5mwdiCx/X+zX8/pn/SH9jvahrB3PeCNWlLe4giyd1B7DLH20hDJVP0xXbkgxM
b/P16dApcjLB6Jwj7g0ZmXgAv84jaBCEb0JZicrsnA59/dSW5VIKJHkw+YXW3dIA
JC2NlIpSrdrvFGzAvpft6suhn8L1JLBgtf4/F2kIQi6hF/si3ER6FOek0YnyISih
0QUczY0exYhdjZyGQgp8oaPt7ODC0WdIaFCzyQMriQ3M46440aNGsMalFRzqPp3h
cBCrWJ2tpAwjuwlzFGm16Wky/xOOJML8E7F5btn5Nb9q2V3HIjVBCnAosrpYhxI0
bWPDRXEKLKCf08F01LJB6q7X8NflcfdeNHn3Wt5c5UFTqqHbOl7bivo8uf+Re0KB
XUClsZXqptua+8TEhpQ9YYu6abh+a+jkcPIHilGL386VOfEWXN+D0XacL0IGGriZ
rgLq7PneSZsia+F2QyYk74EqlMl9XZ+D9hsJu/x0r7bxD7I9G2bU7wKprZICCfii
ydO7AqOpVn2dxKqOnRfEzNdZVUXy06WZSp5J/0SwEnqFk0auMUwzStWSEiG5tTm4
Q7Tvku//uQgpEsfgQRCiOS+LQdUqIOoEb2IdEHtyT1HAs/zCc1JYycWMhZcKgEul
RWVYU86N1NitYvu7yRz9viIoPS5fQTC3gI2VSF5nJVHMab2aFyN6UF5h+ic7bpNG
aoXY/SgRQlKOY4iraWETx46ftY0GPTY5J1A/0wtRgAyYE0bQy4s5R1WfwWS2qcS4
igldtZgqUvKAwHG5613lWo7zZwd7IRYfpofLbeKy0Et4u2DkwtJxnT6pjcbHqZHL
SZg3YB9g1Mt/bNLTIq7rjOMaLiRyZbIsMrjozfOGI/L98caK8Ix94x2Wl+Qh70VJ
7dIwC7agJovLR5zs+mrI2HTCvcajiYUIPYpPgyKt6BTecfO0QgLqNiDIq+qlvCVP
bSQeCRS8UakSUG+mBxCOMDK2uodpqcInBIwa+QdOqHjUHsTBSzLNsfbgxRFmMr/Y
w4HM6mgQ7Mubz0yYdOMrA2yiwpMTxfZlkoUOUPEqstvxEbkHxMuWQV2sISU55NSd
yHdXM+flkWrtQETxxlyqtDTzlnUmEVogrM0ydsdPMlH9Rj6yeXZDjkF1nInEgLzN
3nSuHpHyKv71qEm2qytGX8ynpoyFVYPmEbqJAjn7QWG7fmh+phSCZz1c3jKKNSot
OikqtX4LSsdf/jJwh0R1/GTjHAJS+3b4KmHYrk7gGQx424vUvGsHZdITKQSt85MV
evn47wCu4sRT7WZC4EFVUHqdHFlcSP7U23+hBl8CpMV8wN1ZXc9L36d/iKrPPtJD
R0RBW7HiheZRnn/Bagzc184u81j6ELMZYih2guBND3Yo/hB3WMh8hrVg3EcJdPqC
W4oDqRDsr0rb/ii7WpV5CswHGxRH7tBWkIyUzahd946E4ziEFpmoqZNGjVPsaDM9
dT78h+M+FcsZjh3JoPD1/wYAXpcHMAeAhlUtj/0IYxEu9Tb0iAm3Bb2mhM1OoPb9
V0HeuIfY204Y1dUiWr+jxl3nzKnfv6wz1c/wbayO6GX8i7t7lfDs1X+4uV1JI3HA
Ceq0taS5BtMYmuBeSyQeLx8AuT8VenUTM71ngPUmtzINwHLZHwU9S9YSxRoRe+7n
fU76FTx7ni39UQFqNB49C7ieM3wj3ccRDl6dIc9FwbhAe1XDHWzcIGQeLCEuwuT0
1nF0VBbqWjl/D30bEaDB8NnCELflHWOtl9Pipj0vZ5sWNJYIcgpETMBd/zcEJu7O
ml9MzbN5u/B6mX6C5nmdgTt2rSCRi/IEuJU7iaI5zzNPzs7QbhR5UFBhM9yW2GPc
CGV5GcVW05QmBnngpgqLg6sQ6WBRsu8Q+cOBrqFaFNsWLMIlwwGEp9qjRuBNkaHj
xQMTUp8bF0q3Fx/+ToS54IjI76jrf+X7wP1ok6m9KKrZf606emp3y7o8r0VeyH8J
mAlK0NWX1EalBV7CGAzuB86wKW49A4bKAE/H3dix3tyQudb2QWe9Ur0zm5srTv7f
YCY2UDqJaVDWpeDC0+JiLtTh9+2moL+6XgF89UCB0IwcKYk3QbhWosS2gz+slyir
U/Yc9s2q/OIm44TlHIehLGoTZxizG7TmHyb2yP958lA1Y8woCSx0427rNrTER+9f
S7z/BKWjTwV44Qokk773YUILqO7JUcjnwTs/gZXOU1HauTo6sltzigUjSUzoGFqe
mdSYPn/1h4A+5vGiZeye+LKQ4jxTH6EMtnrJSgH4G0wYEB1V8HdEDES+qobC50hr
3D6hsS7Lu0Fjchicukr9N46qSP2PU2ucMnxXaqFoLLXnxfb3V4ckZmXLBrEK7AHP
3dqZEeUmI8dC8eVP13mmq4jwS/ztHUpuTIcgnfUPlkE0MwbbZ0Evxi5/lnqqzGiX
C7ijNbycnBxtpJNQvuvOagk4utXeYaqJJPmqpSPJJSBtaRPPYC0VXgxzyDocH/23
Nxr87028hc5lF485Komla/xNPzpIgNVzeeafhZC0kzq+XjhLRhP3j7QEoHV3B4b+
96+awEolpvtPYvEjdDmOC6BE2uhZ8gnRLJeUd/Y7sK3JbW3nb4yaF2hTYqcHtTqL
mj58H0m8wBl0TQO0BTiC/pAMB8ZLtq41vZYL53NUrC0xfLpLzoB1ThocvU6Bca1F
Bk79khQcHTkR83MdzSiA9h39/NDY3i5A3cNTrlEBS7ygRC0Ky8G9sW73kITuk41S
IxbxicH2dNeSAoEmX8kNsFTYQJWt59L/abbMZaDIZYX6NcTpw8ZtpyJxXlaOYK5N
wYyg8TuMT1pMKopiCPTlV8oSYnkus0tH1pjcdnqco6IE9Bvk6GAHLq056r9lZzbV
ojLPRTwXqsT8JNGVLEooMifWOS/d3Yu0YRCAOOMQ52zQOO0f4iEjhPTPsrtC2e0z
+6NOKBBySPxNGt3SKdT3nsaRRk/MRSanJonkyXog3evPodKY0GH38seJpCAcFprC
QIUj+TvJAEnQS5TBOtk4dg+n7V33VdlHw7T3haG/yvOdyxiL3LWf0mcxibr5A3bY
3wUZZRzvwjXBDOUfjyBcNaPraMYTgEgV8vc8riXDjQJKev9jpcTLkVd1ZBroKS+u
ZbPfLEtNnxvHOz9zatjEBDJX6lADe/Mob8oWVpz47tN+MXmmeinyFLqxgYtmW/t1
pOl2p3IplVizlKb0aObYYqNcy7nY5XM1hfbDXtU7GfGstjyMFhmaBoVNK3nj324p
MQUNeKhImqGBh85xumE5Bg7OING/cHxJcWOiIopigP1puMtraCMqgoT+QGdHT+NW
R98UkhdDtFKild8m0Gl0L8QuJnz7pYHyIUj1i5hGQtERABx+jPdTHbm+I4raGm7l
5OyAO8p8Se4woV3O0mqPTpY25eP2HXLJQJ4qd/jQu53mOc6WAhyMK5p8cPymetKz
M73d2wHfnB6iOODVSgaKNVSWl8m238LEXxisBPauIYax9gbsxmVYbcAqEmXOs7JH
/tqwYkJO40FqCdIK0boG3WeXSeALECweDg89YgZFAqtfsZHfRYLJXd8uEvzQke2X
jSTmBxRtj0tER3it99lp1mEU4tCNKaeJu/HxXDB9m0O/3PKPcsY7q51/xOhxW8ZW
BOxQbTpV5/lGKe4Wca5qxrx9BAtnU0Vq9Oo+U9SXstmdBNERsuA4/CJjVrhtL/uE
Mm//qm5o1G9pxHh1JjcHsEYDgda1QLUiLz0HONyRgvWej76RmSnFWr5ba+CE2ggZ
aFXwvFFfeHfsFcf7HGC0m+4ATupTIlxlNrtE9IT/UyVzBjMquVWgwXlJq4ep13Ft
vbqtyPUbE0QPhOXtRxlbUpAoaGtbncPjZLHb11wfxHMTINv/RBlt4e18cF3+RyOk
vZXR3MU246HzJAYzkgVPHfwN3ocxBzvDC+pewzQz2Cy4Os618yCn8i1IwhAmXij+
H08gDGd9Ohe6T3uFGYSEGylW+AO1er/k0+RYhP+/Pj5XYTXw4YRMWvECp31fWuXe
SF3FvON+VunplIhcgTghuyJN8vTb59aqeePY6Y3z7nx2iybOKklRz8VfbKTT/seI
vYCuL0a+C3ZdciF4evwUzEYHQ7kU9fDwhF2Vq2TiTjP3ZO4i5o94pvy0PsReEIuo
x5R/Qz70DdBPTYx3YEJ8II1g0uQVbR9eESRM9Q3VXTkw4445HrDohoovaFmeEDPb
nmo6QZlqzVpTZCyzG6DlmRtpKwNmBxJKbSmHZ1MwX/EcLrfkgvVy92BJZoJPK1x/
LOiDCyloM/WJrL9AAlaloKdT1s3OdJdfL0LbrhjrwemD29YGbTuyOa3Vg29qadDH
tKtaOy3n+R0k4tXSkIXeUKJLMFb1tp0tsqMYkZZwR/aBpgoUAHjaM4RKGQyqFJzS
/wd7khO3gPjKhNUcVTXNDnmfG4ZeaxnlbYey4ZkOVf9kMD9+/IXUw9w12hA9osAu
N2y1SmWf+KfFoYFdMOY5rz4ba8nqaB4G+BExF01PFJMz6LdKsyJbJDjwO6oA1qOg
b0ZuIISYqkqeRNDzdnDXBxETJbcGrqPA7XTkEdfzdr6Q9uOWS0qfxzrDKvna43fZ
tCrzLNTGmpLjzI8JNANokNPL/osDEr/dlkirfsVJZBIrDzAYP9OEncuXS/8rs0DQ
XTzHW69fcTjhAV4fD7vGzHUMeLXijmBLFk94RXxu3p8j+LHbh8orz5CnF2UXZ7CS
2NwtfNqw2bNVWSbBeBP2A9CTAI7EtY4VrKO4tkZBM3x9PDzENJcYYVgSk45LNUGa
PFPGMRUWVGvR9IXg38BD4lYN0G0RwGb6SY5O9c78kuSlGL8LwsgYvEJk99XvE32W
j10XzVaLOXCcje3zt3a6XOW6DWoYPBbyHxhKOPfp2opCC1wr+1S06N96PCAuiFoh
ESqCMSBJTFnFeOEBtUg76g/tg06c4IEFOZoOCotKhZVid0v2Z/RUE5CdMQo+aHIe
tNzMuyaLJIo1KwO6hKY3xVZUnZb1LdDui0G3COx+N+AxHXfdxUkzXI+xjrQVAcTE
+WDq+OjnQlve6NytFS07qGYOXEVaBrc0gj9zBmT9Aaa4igDd8bCiXUuV6ugojSRl
kAbss7F7iYOm5zXNVnJK0SMs0cKhv2pqxI6Ya6aT6vREVypAzWjzJ/ReSanxrNz6
qCVSFTEQK1DKueseBeCS2jFmrlTNrdxrDw1g2yXIIPQXsbapsAfXqzdpGjvGhoZk
5YcxzL2EdSSvay5GR1krV41O8/jbPhDGTOLm5o6gOVvDs7H4vyHuRL2yLQ2EOFCD
V4ADhbZsl2vQpKa9Mzf5ZfohlHj0FFBX5KzzammF22yPC7HqlNvCEcEAfBm8RgOY
cfiEiFClM516k5UedrxsLJI38CtoNsj8XhBGiEWKGfCLqSaSlaWKwZYKwhfylwjN
z246A5VZzFMNZnBIKXFID2SZAgEWHEgczLDj3TDNOPSroRgrK1PRIgAjaQkOvyX9
Qpqo2kOKBKBMtI9SYdCniNUzerB4Ee2OjOquTkAqM2NHqPAZo/NOVsj5XM3Q4oOk
Eo16FnkV2MAUp6qONuHRhViEKInQGN+6uz7yZlDRd7uPVly035tPRTB/67P3/rXC
iPgbC+tTZjJuLkCyz8UEYvmusrAdRNcER/7IP7ZssBjfsgzJAbKSE83pbDQt9SaJ
B5MVthKzQhIAX9j4hVpH4eg75fHObjEoPIoIiAw6OObhlCdErkLIdvjdI0Q+spdx
ZTFtkh3dgF07FEIzPre3BioBPGobdtYb5IxxYCcg/vO5sfDHGXTznp9qSHk7srK3
l1uWI635YUG5h7p9QcqWcSQo/V7HFvonA+Pk5EjARmvjc8okyyR0Q2j9eKNC44di
b6UdXQpuu/BSE4ZJfh04oH6bS2/hz5sgX6TAnO8haSdltjC24Ywu3Q+zThu29FdR
/OlJlka06noV4B9juL2cZj705v4zxRs6CyCbsXHZGUYS0QqMnBPakD25iEUYYw6P
T/uzpfrloaigwp0m1xlk6qmEcsGVoLmsY/7+LdbFbmVDKH4xs7m3Djp++qIYhbvx
BsBdRbTdjd6jttCgD2LILtiO7SbNIcbHJeDchCcQ7Qdu8mQiR5aF75JSUII+L8qT
j1SgPyV+0tAmeniZCDuMiZO6RrHyt9x1BRpXyWWhGhOZhAzPpaiQiKKXB2nYvIxP
v10/XJS0VC6xV3a/Cn3wDtIpZnWFtS+ljcS1fmejd9ICWcjPd2Iy0aTvSLdv5G9x
yRGJ5AGTxx1iDwUAvZcNYTS6xbqG4uTrcaEv1DtreIeRMgheqMyINHDbyP6uNfmu
QIxaGZ5asw5660+KJSWNBsJATvJmWCNyIHWo/+/KuHV+JZkSQqjUM/InX585tGOd
R0u0r1xwCCc2JX9kOY26tW88rcDOQmCpvP8U0FF1lx7bFkGe+nBuGStNI1DTSMxR
pU/dR63+u24qCmSsR8zCsOAuFDRJIXnN3VbGYa7FXfH51Id5+lUZyEF4T9gm6C6S
uBalSEQP7WFK2qkX3bu9SF/5HFyHbZWSHaVm/JlhBzrgZ8o9Dbq8CVYNi7wvN6qt
DdPhDotYSNpK0IkaFkjhtzcal61+bjDt8qgsQFdPZJePSTZ2BH8702iI0plzEINI
Y/w4vMLlLBUJrGIAj6kuGUj//w3wja2MFa56uKfctHL45/J2azVkjKHl/khX8ePM
Ax/XqoRUIzS2Z2SSuIvXLzvRCVIkQecXVCp+SvhoxtCZ1f9MtgbTkhSSJuR152dE
FkarJA7Tj1VPzCenDNxTuxViH/mBqEP0VSKjYQeviLPr2g4V01gu38t8fgJ62x7E
3Kxn2lWTcb199YTi9qsRU+ms11jvgpUm62uH6kbw3AVNh2z7pXWGIDsZ62fqqddL
pRbm7p7PUos5I8rWoG0uyStF3HPBWtnXzcu3eaWrEsxT4TORbKWT6+H24tpW+NEp
eN7diDWctyQJeHFJ+dl8aElbVn08OZcoAIAYU/eXPDd70sW1cqZCV2GdtTzP69je
lt8gTs8fMLvDpfe3yYDpLvZyf1E1PsbxKJOklC3aY5T+2WtnJdbh5dY5gpGHh4mS
Bw72C4RQJZUJsFkJmE0cKXHFYD3xVxedZ0E6DdIFWPh7v+KnQbpGPtULw7QWeg32
XTn9FnkDfDea+kiamsTz8CYeVHpJkezSzNQmuC2xWNUK4AoHsqJaC3qRe0HDAQPk
3qCLDKRMrudPOIVUjl503yyPJmHeibOxHF4Nzk/hdWL0mwO/lWtVMVCmOeFz3HXh
OzF0agwGq/w+5NbA8i+SGApQ8MctAyJ6O2LKSNA0o22Mu5p57dyXhcxIqnt5LLIH
9fVaUzxlCcpe22XU+DOSV8ZBO0Ooa4LtzgzTX5ACc5/WRwpCKan8xYfj+5ygu9pg
jazpBynrBok02GBe66n9syybQmJg++e5R+9vxoZrEoxj5SznLIWsR6ophTWygGPc
J1VgwosLOWZ8yNkHCtR56ufOgmHCqXte1fj8EN9y2DsmtvWAAlo/vh04DZS9CYKE
LXh1MHDk21BNOnqOyGaVvAuqWwDJbMx/0HFYrVyrmA10UyzdXq9hBnewPcIDVinG
DePtodt2nWWnUeCBdh0TqL2Q1CFygYukrqPn3TwysPy9U1hab/V78gIe465+5sNR
LjO1lpTPeiLgx5fbszaI//CW+uO8Qn9CqrkD2lt+QAQzip4tL5ojXW95E4Hbukpr
Tfr62sQFjowBTywNWUkCRqIrXve6xh+xHatvX7AcOODeIHrShIJ8xKASfMmWFcg/
+0Tgnoxz7pyQT7VX6fG8FxE7hhTaNt9wgb4GoTi2bGn3s7mn5s4Jokon8A2u4eQd
ONG1ylC9FD7UHlQtqVUGsE0IJGMx4WjjCLpJnHNTa0qdxs75BrQhUFLu3OzLmAGr
+r832UrJEd8VkVpySnUrFvoGSZoGR71Uv5EJl2y3BzgtZmH724j7MOMEdJOXKn3S
btOO0TXrRHtWgeL02uoLzUw84abmokRMEj+MY4AGQMH2rVEN1JPfpA0QXu1aVczo
VBg/VhOg46+G/iPBl5hGIo5WA5V9kanQa8Lgb6tJDyOvUuoKEbfDWHCpJSqFKf8u
aeJTnpU0f13nBjNhPHAgTCftfQgYzF+umKsj210ZCQRzomcHe/liKkiQHm8anAi5
bQhTYfS4EzoXwYAiJRpXB0RcT/dhpcAqb7vV4iVADHXoV2obej5QcZdX+jq76QbV
A101vXijbsb1v5KoPjVvP0kxXHTrhEPK9S8UCEK194z3WlqEiVFbP8t9OXS33yB6
2XrNZ8j9l8BWRVFYiZ+ZcZ53HcUWN+aWHxA1G1+2n2UMv8fvGBs/usmK+ObFkXkO
cC3Bnw0lYBdzteabXJwxgcPUXI7cOtwyeyYBpdKiVkH+4bG/YnmEXsXm456ULk+O
Rcwiwi458DFf8bHTSdyaXOXC07uDaQdSDdV7D2t/EHrfE+sLHxRUxPc+ybJtSI7N
gw3oIh26DCsItD1FpnehUVjnonfp5c1P/rXcTu4pAR/BlupuJUxiUTII0kmfXINN
rVxl41gIwbo5mY+yDuLafLuMUcLy4qFkLIRMTlZBtfpp8tIFWEcuJjARtAl1k9gr
U3R/CzcsyLA5dcXIQpUoA89S4NXOFi6RNMBiyPsKAHFDBH6i0qKp+r+HBkWPIYFo
ncOqwtmamAfC+LECCTA1+15MVNKZrheEAye3iCEmdHol0asRw0O41QYbuWyYk97B
9vqpSIWEKeO27NX+srIIMJArJ8r4lj3mK2ZQhBqUzu1Ga6IgqwHDfh6zwlhdpN5O
/GE+6oqFsyF1U94hcnf/PDyW7VbS0+6Aq8NkJR0i134pOf7Wcta6GxCzhVUtH+Fk
rf5Ul92CZF1mlQ1jsZm6JGxtTq4MnH75n7QWR5thnxR0esOb2vltN/bHvjsHUDG5
XP9+VaGfAXL6RazuefnhnCDTDDB8eNu+KM4kjuMFtWItsRRKkmk15FtaPbUQ5Eg9
xcGn3g+9swlLJR4gI6DeO6LG49mxSanY06Orj+Zw9bhfltC4xmSgo6UGCODQAYMo
mUlZ3bmIjWYthKeOE2rr2YOhrG+6fL6qkWcU9AJxr9yzelIGH2zdXE1y3ugG4o4x
PzkBK+YwmuRXYEX7KIymQere604DmpuW/9Tw5yiIDCe8utX73fSMG9OIL01dj2dx
MtlStLhN/Q9LsJAIosX9vafcRjjPDQAXE2GlZHgOtqMG496IE+4POUtxmN1UEDXi
Mb5ZxGiMX6LA8ZEjMPsCmae9Bf6D9+iwvytIefvSCWyES2dq+BG9j3R3FCnpTsEi
MgiDDzp4OVuxfNPjKfW9zfKKP6+NzLcbpHZgaWMhHbMUQzHM48RDrCt7XmgYR1eb
l5Ssfy8SODdZqbh9j14hbHSJcCZLYHF1wV3B9M51iHe+1KKlzuVbzpYQv1t1n1sN
+Am4hp1IuES5sjxJhmtD3f8b8rwFBjUoFGgM1tJGT8ViUFXpQMdMrY5yXJ5atO1A
sd/eTcHu5IyEhiS/6zfpSSbi7UNm9XZEgHXgwO7bu0u9rDQyGSEnmnzB5cV43PPJ
NAlsUbK6L3tKzT4Ekh9TpZlfokU/KQ2byk4Zw+8TCaaX+ZT2fSFE1OHiyu78dSp8
Jb4YUVtlaB+7rt9IKTuJlYolleQuU9tAVgduISr9JTo5eRKABdzHlKgrddAaC7sA
cstDNb2y4F/fPYSttGo2eWgOaXQfyMnCRyI4vQkh23fFuBugeFSLT2hEFHp8pKaP
V6IOSTVOpx+YbcdroYMhPriEQWryC96/ikRtntecQDiEFiQ3koOI70XN6iCfKIAk
+v6rSEC/P3LRjRR5bkSr2lm4CfPgapfleiEAGJ1E15JDqbuBmOI6nDjLs47AhQyr
2o2704pBBUsWHVsjvm9gzwA6/Fvmzr3OBjaslC+S7XmAIQuTSFVj6NcGnwhdb6nw
jqu/mGHBnjnn6od5sje2AkT/7JfC+xWjiQ2/0AnjmdIOZeIpQ3+WI5PqEcG1pbo+
IV3LIIa3P2u4f3z+Fe6bpF60WFqztbu5ubWE92GRzwpawOLFps7OWcKrUY7w+KFQ
BHgf43k9a5pRE04L+g0kFzWv42GRyQ66w1uNbK7nh5GYmdOLYlBsXxqu9SjOKj3n
zIAd6KUoY6MDiTfRWsR0al0hdxSCBcUNPz59IQKq/oOVFZx/6LlZrDmILaddltCj
jf/hMwpmCzF6JlQZQ6ObHjAjJz+O7aYs957LYG6YYxQLHwwgsi7fcQ9Moao4TAYs
WasqtuMXmP5D4Q/5nFRoUpLdp0KIgngiFNezux8vR00irkCQh/QEHKYbEQ0b/4lt
qfe1CL77V4jIVyZbGFENFTbuqu634um1da62wLPE8tXy91KErxi8K3jgMh+rTvlU
A1pDQFA8vMiS18VdnO0OnmTB8rKt+aUR8WYSGQiFWqx3ze/WH2dE7PbZfWCBWbI2
ql/WZsMSf4Phbgam2u9O9gTr5mo1RTpq6y+caUhvinrKqcI68x2bhwwbQTe5vx06
Vd9eW/nnlEp+izUpP8WOmRanGoMJ8ei4FamFQdIr4baPtwh2pcvgnt6QYV46puRU
0hwPfYoJ37ao/o+Hsm4+Yxt4qQedc5hZgWabBYhv1eSHWjjawQfhY/l8+LY/YsRR
6Cg7bfZZnhp479gp4fvxkW8I7MnuZPQa6R59KB4m47a1qAFajgszeWYiVXVzbJ0Z
J4WrD/uCIFK3uJAd/psOzaBy3TPIZLtE0oWTswH8cTiHoC7swTUABzgBDY/EdGFF
IGTSqaGj0c4HAva6XjwEdAgVlA7YZ0UB2rNJCyr54IPDKbkRR1XaDHR9s+o3mwD4
kb967Fz2obvE4wUJgR/ylrnD2kdJgcUXx2/ABR++mi2yJ62EuqQtn72DgKsoXCp+
nQgVGRin2iWvnHfq9mz+s3y5IAVyrvqFPWYD58LKjiXvr3Xs4a01gFRRR/I6Z5YD
1mNBPQ4sG1QeE72MCPvF4pGcASfhPgR7Uagxn7zkH2Wb9oo2kgPty1/VXRjFTRlj
USvOYdvr8ORSAlV9m60fYALAygVysWQuCw669GGLkNRJal5Ao6e33YWQR/QhU37j
pBk4/HuFC4AqZw5z6qGWGxQcwYlWWMt14glUHvbl2tkltm+lD+0P/949zwT2TOCm
pqMnnduLhTjYmXuWOk0Qm5Y0Gy17ekWSarmwU3K2Qn0ed6sVHLFwB09N+GGLjPYI
4yXLvpdMK/I90KBQi3FB4QOIfKOiIO7dcaH48DdXU3yZBeer25Mzx+E3hMC5C5wV
5tlhoVFiXL/2a4GTTbu8NzaHzFg1yjBsRPVK/7XrpJ+0muO50+l4Q5hJ/MD/mqXN
x6LkpFFOsvOTkOu4bauAukozK+HbF0IFhRyziJTixi//QM6vckePoeeXEQOz6/ft
2d5sRkhDZSzAsCpPZmNMAoU4m2CrFpcCL6LKCmI2BPsUM4x6gpw8a6U1TmwRwlbX
/GyNdiQpBQcyL6CIySB34tsYUsLPsm98/w2dmmTDdAAr323N57DFZeMqf+lQh2FQ
iNcmuq6i25mnAxeW5j8et7eD9+uNmN6CU72tdsKhxl0jsR6XMsL4ZVAyZCNRU9da
sitezpD7r0/GRGUfwVQhgn9nSjCLLQAdeKrF++mx7fRObXmY1HUwFXN5LP9rdmlO
YaCjnwCOTUwnL/pkQgksn1V+LEAbYrSK2MuC3I6/GYZ0E0feN79S8j0BiX6PSVxv
5TGVqGSiSlTCvHvYtBwUVTGC8B9y8BzYgPpXYtpDiEk55Svwg1yDMC2f1A4it/Tm
Hf+gn+GFu0F1KetG0f+Koh0cijZCsxwwbzuPRfFgX5+KygmY43pAvVy4NWrg9Izt
ssikaIjzymJxNlZLPjCjGUHP2wFpY/bJd1qPgBj/cAup4J/GJSR+l37abncbFJ/k
hl94DEG/fnUpwtc8b9mlmVqY4xc2agA7w1ylU8gtEQpCk4ly1+St6ms8NaGteCbb
hKcMkDQnaZyECvJmXqrgu+qTnMkJvlprzU4CtQoLTMUTHKilUNUi22u5PC/Vl5zD
cHwnej/egG8cit2BvmeiIE6ek+3x/wuj7mY7JtURfaQOijOONqlPUv4TzCL3TyH7
ZXXfYv9lwp+uHgzySLVwuHfYAJNKoNy53R3tSgalkv+m5dQwgRtQqTsAzbunuarz
usGv1Wo6LyUXKLg12TOTqr7T0fSZxnbxpGAMjMcH61V6xOAQ0mwvGX+ECSDUSqHR
1oymLZvg1/lH1wBNTvabAdrtgAevDA8fQSgQKZV3jzdTUJoOKCQoqt6lH2YD6mzz
YdKqhHEvVOpFs1NqRLsViRPprd0/tDBr0ED5Yx9R4xIkP7sOY+Yegiu1oNltikJp
PXOIBCvTdOJl2wnEZ5OjHwnmg8wITwwOaGPSRyCIRc/0Gp/SuBuY1xmPq/+GhHqD
KcKpu14S5od8Z+8kORDvonYm9H5dlNSsOEA3PFRPzne71+/GE8coj/a5djLbjSVO
+ruHDpgEKNKOnhdpYn+50hvYifpYzYkO9HZzKUhY54TfG9A1x4gFxB87/YHjXZd4
tLnQkshxG/3JohuIuQxGcSjbEWKX2RbQ2go5u4OS2WNpKenEzB+x6NyxaTT9XXK1
ESCC4l1j/f0mb0Uiecq+fC4TqW+G6cFj+QCFMHe9RTEwMG4XrDWVuERJd33L/Ucd
f6fKQ/gD9416hbME77cwY2tBB5QvFgW3D5q/oR33NVZ1aBuIyRbM8zyaH5CiZMqF
mAueBufyMeMbVn3iEf5MrtArtl7CrIKXaUDsqPRHpB4HG5FM9Yh8a0rGlRcUnGQ7
kLrl1FzAz9+hGuF91Tc7pWYgA+hra6+IGYNeCeZvHurIjJri2BThd0OWIyTYmCPb
u2vzxxt71z4ztxtNDRPiUvJE5dn9i4JC8pMRh7RtOs2sP4+EmyeoK5iJscU5KUhf
0DOmWD9R4vWPXtK010yhJ77IXFIRjUP8/EDvHPGaIG0Ndq6vVYsDXx4+gD0Mbacs
VlcF8CsheqE6HDQ901thz0SZ5+P7Sz3DR15Bon2n79gxaB5envZg3SeT6j05zPwQ
wRUS8H9YajRlEPUEGlZGITJJoQCntdkXzFgHqDjdkvPVvWZy9wA3jjVUPjufROWM
UZDTN96NbWYmYX2y6LRdlXHknEMY7tOBZmMTz1y1SFlfUEiNvW+jGwA1poPjaksA
b0L6YknLy9Gfdu1rd3OLmvCfUZVvTdoUr01trE4sDoUKG0E1AGOqtFCEXP9OYoE8
qx0MXFWTT6YFgR28l+i49wygKrmLEGY3FZS2BsPyWOzuiQqy7V949vj+JjOEqFCm
DJZVyw8l237oEN2xc6QLkhODuWecU9zi95KjNDJdjZehiWOJW6CKTFWcG7ffazh3
p31vagi9CD/uqB/Np32taS3U0ofMir4BhInTghQoM5/Ju4QvjdlEEZ3HpE2cZc4g
AcQeezd2ld0SUszGeYDK1z+Jnsa3hlf6D63x1/aM8lzU7+wjNVvm+xZxRQuiotUu
cA9PlXUxx2LNK11fzmoMygV0sERVUKNmy9bPs3OfPrIYU2DAmTatjhELynzgi3/p
dDdiflGq3KYHi3xJcMhlrAts7nLgS/586YJayXsV8qUPq6P1FFMKAK4U3hIFe8bH
WxA+NfGE3sZ1Wrl4np/BvLvH+VD7OefHkZia6OBQmWOCNUKEieJSRm15/WCKwPmp
yw6FyT81LNkRNyiBOA9wQWdXeDZqfPJobNMOZPm3qIaR6JnMSf/Su941D+9xa+nZ
xGpoleDNw/yZg2+kEW8AE5oyAKugw5VZ/OnSH7nsKdoF/zqanSpVUVhwZFKyoMOy
c6k94ZQDpP+AEdEfbcsc3paJGyg3du3kcF68dubzl08HyvBSrRkZj3uWpr75TCcN
8aH+i694vE6c+L4pLASM+Y1Dg9Te3sbtaD74LYVABuguHyrI/knB5sTev9MvUqKk
aMdhTNJRVDonaQ6phU1kQFCDIg2O1DkFdado9sIkQh9JyI3OrCmgwJyw6Aj59A0P
bsylRcuYqlNtLbSEThbHMXtRNfgevnH6/gUq7CVGdhW1RmH9Z+tT3I7dkBAPYcSz
2OyOLjhNDzs7/6L5pCouXc1I0oMJIRjkyBz4LsX9o/ybd6/J1VElk19zC8voa6+L
AJKejEq5XD9AoOBKJrKIpyvABagGph32lpt9ELTwT57OGJhoKMGXZO9iw9NxiDTs
u2St8Jgp+vrNuB2MZ2ss5VucXmFqW3zqMVKDPiDHEnpq1XrBbfDfZtfGxgT27I6D
Av5ec45SL8Uwb1LmipBnmzPdZrO9rfB54Cyd9ItuV11TTrfAHKPa5OZ81cIYuQVO
+iRimjW42mPGK5QvJ6wvnzloqe8O2tzsH9QAmYR0iWGobOiaGdg3XQHJOVY20afF
uVnC0wvfGnqHF2//YXS7UGkwrQnJlouqxbUaBsTqKrbuxRjxh1sDqPb25dJkWyyV
B32T2M/Zly+KS7Jer2yH44JfZ5PFVVMWkaZZV3+hyWuHhglW2cHghJYNrEhOGE1L
kRGPfnLTDWbESWVQZDmHS8fKW6kUiua/b+DLT/P1vpRpVEy/Ma8QrpSU4umeZMnB
PNhLRFnzgmpPXpMncNASZh7X4k0uRR3uxdOO/+pXHZJMMiN0wGiWZFPXrm6K8C0C
oSjx8AaO0OQhtq58SMn7NBb1n53fxjo1hfKLO91EQYsm11dkt29/9jR4/MY+kUdJ
FsYglMS2QpEaSjZgeN8SqqzAx1WPRJX7wbWkKsH1pJMQwTGGAP4eWoxlI4yKQ8YV
o+5VeJ+9kmm5d342/Wzf6BtPpoqrENH9/uXobGDU3EEqSQ1TaTz+v6AtJ7MA/cO6
c+JVOlBq58NpIv+b6oKahgKgKFsMuKJ+hvP5nK5JLQbnxA/ICq1/5mxJV76UTzSK
6kpNYSWxA5c2opJWJdcwSrNOWVYz3dSDoNqVnHxA+2XopfLQ5J+4Lq9JfKVRT0Vw
4aXFwshAlrKUIlmvdoiF9WFD9CtOqdqDMIwBhTx4XrHPoJd5AOusUwz5X/qjSxIc
o/KG2L2E1P97FGCj0cocvXdUZm/PsgaCKHXyzSmK0so1shHx27rKFneAtyIQ1ZI9
ho4A6FYPQMy2bjj3lZh3taFAaD9VS0I/M2z4VTTyBoufqvw5dwKvJyMaPrAjEPkq
R+DWQ6g6ZiqMPEsNRus3R0SKRahDaqfiQxV/l6gNWWZCAVKfSxEF3CHNOXan57i0
XAcJokJcw4yRK8RTcMFQsjOrdp5QSsER0eOAey92z6q/DIusfWucCUrxSMJOhBRs
4OY5KrIqJtSFEU1/4g7RTztwiAbVNC0/+uFi3Kr+h8XWjrq9u0cLsyqy1T6In59e
JAHiKPWVfnaIGoNbn/A/VEJQ20UYwmAmk8KHPYCVxLNUXHJwy+zGkWJYxVriyjKj
ysOseoTcKATuv9qMHVNMhXL+P1JblSHpxKJxq7wwWgUgVUp9uIP+8eazjkDoF3c+
FTfGt+MDCc2zMwKelsUlyQ+d8KVs+jVA/wzhw1fChu2EhGxmfHMuirTibsbzmmYT
7dgb/Mn8D76vYo8zKzA6NVnzTO9IuD6z2DcCKcsKEHLhZiv0MOuV3XvhXxOoRfVM
R3nvMoP/1/qTLsY02yPcpGPeGuyMokx2/jngBoThdQ/iL/9DEya/J3TGh96jJQwG
E8cNh2+/qgML6EGK1mS7lh/mBJ4/FFY17gLlMXBQHemANWM4NkryknivUIhORG1M
DdI+Mc4guXF6TFVuPuIzlBa7IcKcfLGSe5OpjtrCaPEd3mj5GspZDxxSwV5O9+ds
qvZ83xdQqWi7TCdpLVsvnjm+MeDm48h+RsclBKTfPky3wmM+TdS1NmLcPx6nr4jy
5mNR0qAqnxkcceDUQOvWfirJ5MUXUhIAifrvT7POp6tXi08NhcemI9pUG97N47xa
t2Or2zqN809yx20i4PitDlRO6tz0ptgzgO0/oMKFxjxOV7F+3ixbioi1wOcJw2ZF
doy+i/I5/vwDlEzNKTE0ae7DdQUqR9PtOZJUGsypBP1iTKLDr0gZv0snrJNo6sYP
p2Waf/9FnCE5eMDKIy4o5j1583IfNFht6ZmZXcv+sOsEERycG5vGfH1lJrvjYoTn
mAbStC+tzKquGTnNH+HZKrS8PU0kTztrcz/xamLE3aT6iJZ6A89VTh+q3FiMwBv5
u+foEIRo5Tbmf3lpA67t3NzW8N5JEe2RfQXluKp13Xh8eaX0ByVH5vmcVEzQvmUe
L+sdRJ3VizakKzulv/LrQcz5vdOm1Sm0ixQjJRcN96aXK/HLv/AV8KVTuGqwMPO3
6dg5wHqy8wrrJ+x+/1PJK6IiIiSMGIsKQcxeg4dJ32gZ0pRUJp0pYKFLwJPTPDYu
+g9oOrtN0amJxqtFhDF1zyZmMGeq2ahuwU3w5wIggBfwHDbu9jaCCfdEzZSTUwsX
rtNUReA5aJQGNrnw/QW5oFIcL5O8WXTPGuOyBSoYljFz/4tRzKH9chQBoiCR+6RY
tjgZ8nLdZeRKbDz8BP7jyGmnnk3NlkdxY42803VP4LuhSI1u4cDajIIwrUDCp38W
rkAti4jeUEilyUD1+DE1IhvHvMyu0NjBTjj+EHXzqt3kHOTNY9DgtRQdNtvpy1es
ch4bCuVfWeneSscXbcy+SsQreeeGt5vcdpAGk0TtQ5GdtRpYTJiI/4tXTxF2OVT5
As/40VYKkAts4slfKHuwIOkJSH9iq+2fLUrlI/FgrrGuifnSxy31Ng1Sl0fEnPDj
JWA7KiaFLev9dF1lmeAoNL63K9ZFPcmHsFAjbtPenwTDBjPLfGNWOdJ37qXWM1cU
1/+BCczV8KKR8X0JXl+Z9h5qE2XuIs+L6FFIlGxIvguZ63M9F/gRjCidITk5gCsL
rGO3Pz2zwrz6BFO6vcrdgGv3YGPlw8SYJj9cc4lAsnaLFDYf7yrA5TacqMAiZDJu
oJqPnk61QQW3ImKHJ3d5Or11IzKxwxuvck6IbIj3lrmBGwA/P39AmeTZ3E8QxMaY
DVTRutp4G+C5j0h0sSoLANcunAMMXlUX2E3r0attIRyfhaJ0XAH5e2pOVIL6V0W0
/H8IWKyjpOCeSv579GTA/1u9NZMtGtdHmtaodg3h78QS3hzqGHcuNMseQmz/g9ij
cafesgLBtV3w+BwoXoFHM1W02lki6mfkM39v5LyGGtHJRSduGXfrpwAux0+CnsZO
Thintd+IabvnpYX6SsQQmt2g34WjOx1yXMZNFIlsDqpgTtFBLGmoAmS5YsUkg+OO
KfUEXMsRwWaKCLEIAkflRItBxnz+NjAzfY8If0VArFhRuvwu9ZesJDyFlqGzkxU4
xjYrkvLjrnT8NYG507r6zyTBz4rzs4vfUJZ9WsWrN2IazppGyXEAhdUGlWPIVvzf
uYcoC5wLHCrJ74GX+rZEvZbIEYNjXlcCSuqwzFmHiIUysGXhXPeplQVPUG7wIWGM
7+TY2gGOerK3PARsIiiLq+6wxin9knDz9d2gEDdbRMGXB6G2zD/4j/MvVHWMX/kd
XOvDo9c30LiNX5Cd/pNgY7dCgYOMp9zWf7u0xLMehZrFPHU5pDqGZyP5xdAq11AV
f6sH2fzGdv/CdHt/P3B6Fc8MJl/jzdBPKIhr2ruv5Vw6RmeweWyumztlsKV1NlQl
40bPJU1/L2aba5v4nCuk9hmd2VEZYtGVvIjCzHGQVvwwiQY7I5CYpuBxD/t5Nnhy
R4e7kTrWzu/xXC5IVpibvXllPEFsNLqE6tXqZbitd1dUEEjytdJO1bQr3ioztYRj
AtESoG/Bg9xijNbfFZCO+RM6p4FbrEHGz8xcIsgEZxQSVwkX35ND8PfT6QISr64P
QgFUC/f/FTznd2Q3rfOChL4h6xZJyKw4ddiEKAK6Pevc802p3D+NndOIeOXL9Aw/
1Utdovo10Jrd5dicmnKISsf+mpgiYk7d38DzOyHz/NTWpNOj96j0M3hFLL8LnYBu
PS49oPOE8diNZgNhvpwmUb5Z1TZOSIHcwTn95AKf2Fe+ibPSED8SpJd/xCjJg5z1
jr9RXRTzLUMc9fHOXMkBBU1TUp8Wni38rDE+pZpVFxR+Fgu8aiy38x5j+vmR9bZX
tQV7dugVMHBxTy4k/6jUra+BrLTEm+I0EQ/WratkMhxjSDA14stvm3PpbDuAVBn/
aCmx/K9fUNlWVOGI4th1TPrydk7clfbB+DJZx+qHY1uoQ1bYL8fk221d+NGUtoYS
NOtUANcOZEJgikadPGfYSSRu6O9v5Fjn/IAe4/x3skKF0vFheuBniJXjuDBGM/n/
8g8xwYw/n+RIjqs7qL1Tb1rkZIGlIiXtcV+9nHJIxRafgn56r9c3J/30a1MmlyEQ
AoRFS1iin+Z55d9/IVQOyWs1yMUjeLKJGJdoPx2OAclKc2OJAIBZuC+XmM/uk5gL
pUi0nlxrJkUOHre20rXzWiPpb7NnsM1AWBZ640ISoEbaRjW/58PlzNK+O/1Vq7qn
dMPLTA1Rjs3sT35urWsJOGDFLm6ur/2JHJWZY+WsYfkx3gmnHUkgPiWn2dgmB8Ku
+eToxyugDtDTY0Wl6ii06zcQFrbvIEF/yeB31ZioFENhaNSCLJEbTj+eedbxZZGb
L5VO8loxh+i+Cnlm7DDNFi5vKgCeYKB0mZRK58vh+yE54PTgliJGq8A4rFCylhoP
6GsIYuHNojll6lUqLxHByroBYcN7JQz00O7SuvVDxX8j3Js1ZhOwUk73AcxHLkTU
o1BwADKfRg3qzv898+GJXkkE6fO5+HqXn5e8p6p/YmdSNsmKhREPKQYojxm99jdf
rM0Ij99eNJyaxg/u2rATXOtr5VIR4pkNsQkU5ERhaoGG6ng16wMGfe5WXPYeW7Vx
YneHAc2fAq0qzt5tHOxl88LsE+I2JZiKG+5L+FpTWvEa0JYU3HLBLVUiCN6x7vju
EsdhW4igVedzcFYGVQUSl74vR5a8kpeDxisBQCAQkSKnK115S6kejHLNTjPFRGxa
jFIhIETXZXHRukUcFPMlDnxoHJrv6ZD3oT7Oybtq/raZsO6U0M79rcQgB+ywDiNc
RDwZddRmvF8IX1Co03eg0mpZe2jOulAYaliIZ8TUAvJR4hg4icTLT3SvMit2e2uT
BTh6s6W0xedCxYaK99zE6WG2/tPEQZhzwyQhTCZeml4CGTo0RgQKH4cL4PBj6iM+
8+xhQ+btMLQ4CI8pO57fbJYZjCMB2fBVSW+9LAo22FPVzy/NHJjg74dsbXPx0BVE
SVX80kJ+JywbT2lpIPcqCNXzyEmcLs2Z8+VEYkbOX5xSN2QpIWStN7zDbvUR/J1e
0CJgBgO4pFvr70iyp+9kgR3YrzCFZRq+GeS03lYyngo8GC7ynFRtBDCG/ghuoPdJ
ouhkLesDlduYslww1iSX3RddEpO7Wr/nn2TpYQdV726AjTg/zpSPJ9Ee9dMfDEQh
14C1tmMWf52qeCA/B5voTT/jzj0hSOtwucqPVVvl0Eave/4Re+O0KEmq/qJd5kxN
Jj9lmD/h8JiHWf3F6q9RzC+OwK9lcICjwIwYlWYQ4z2v8oBvyd9qi5OpNu8qUGKx
CXBDpAKenOtG56gE5YzQ2nBCyimk+OdQLvPdholE7Bwwh0vH5wTog4PQLB/QFEdX
iKLQ2XIxe3TLfCZpWnJsEOHcyRRNQsdWKKkaY0GY7jT5xIa+jq6KC9drJqHZTlQ0
pcAEtzuSTTyGFNQMnrAIyEsGQzWqevXVmnXwmOoLjtYKJHkgY8Kn5Xz3dDaY/XBG
mMuekakREd6o446syf7tGfQMp8yqD0qJ1A6V7HPe7w9K1bLfd7A5ooybs9wkFKcb
uMIYTGeGW4Hc9yff5u30zUrVS3IebNhGqHMYqB4qtOfoaqrRfHmjs0OrP+V9L8lA
98pfqt7FgVRkXzeWQ4DDLtFSy37YBqFm5qgwf5cT76ijpXgRloZl3ppHPTXy3d2E
oDxNUe1mxwsJU+z/759ekUo6Rbj3rHcGh9Qa/5lmfYdOVHOTZftrsZPe78oGEW++
Vg4a3urbJ+DMMKgSN4o93dGNt4csx1EGhO455hd3X7fFD6enH5c4vH+h2Rwhk0qv
M+dH70q5AVrACsJKujIEzmdgwzfnDchBTZrxb3oZtZYBQoIScSOjiTS9pelsoTUJ
F+lXzA2gxy592QRBDpwQyMzGPVWU+VvZAhqI+Ps64GlEiUhh2Xwcl0Mq+JAI0jBF
YcebSycnL1zNYfTWJY/rLLyk8v/OxQP5TcDfF/dl1PpAZLE3+jozrt4mpYsU3Rig
HIYEfQeG5J1rFcxwXjH6pR/0m2qYiV7GQkTdciH+FVIY9kMQ4UZXkmAFceySexNA
qsI0Zlv24A/5g2jgp9ZIt3+ll9IOMABbgDGqucdB3pq5JPJeNY7FRAV60ml5JUAG
BPsNzghkzqpkCO7blYIPktaIcEpWB9gdukseUYTpOHvqbT0ijSmXv3js2Splh4Hl
+ampK9kGP9htExj1kcyBPhe6yxw5x2iptehsSXl3avCGUg0aoU1qXUXUNCAwKaoq
1qIzS2M6IJ3yvfB+zkjb7RWpfeeukGCGf8cQfs1cwbmksBG8K6Bamefv3FZdbxVi
vlqHp3C8etWtxEAqNroRmScXE/whFqyDqvcXOWgOQg33BA4gj0S4s6mMV872kHZi
j6TukloXEVtVdtDQQnPhAbxuj7EcWdJYwbWjFNFT2EqNfKxDDie92qwqdFTbF8Qz
EQEVhjSAAdzBvuzqCPIA1D/ksuemGqS7IRF09CKy/kMgEyFO/pqLUMgE+zRjLI9j
1WE8Cbo6qbxc46u/jL5fNNJgw4M3GvwVs0dfL2YxHD8GSQ2MCQJCoWrMYQVjUHQk
EGKYrkK6kWu/aduLf12NCu+SVeELEY/y71jh1Lp2vD300pshuQjpGlkbqbA/Km4v
Mb/DQBFtUrfcvC1UFM83xMEoYkWVGS/qLDh9EBZ0EwauKxVXBTOTWHD2P8z2ySuy
B8LvSk1AzN9mDpH/phK34zH+zH/3F4SoG6dFWrPb0cfJzV8zmr//9PuBP1GFvzaw
ICviJ/rJS7NucrNNPiVU/erCgpZD4VFH4E4MfxCL/uF0/0S5LxmBgd8cTlBP6NQZ
Lpk+ibCiZiVUZzOmYfLi3Aq8fm7UNIFLJWzv/ewklb0NhUsUVg1EJJMW4Zy+/kNk
3pSooxSr/X7CaFgboiMSlLokaGneqm1ZzPEsoNujNGxELgiVKVbml6lRZACbPfqX
mcj3cLfHzoJn6T2I/Nq9drwFcwPG0SciaKFnOoO2NRHavvNYJPr5zu1Y+M+yBBha
pglq3QyQ7xxPH5AckuYHL2yj5hKvgsA01Z6fvC/3tfjpjUcfsQyuqn9k5c9+J9+h
fFwU3HUTXdJkr6fdPZBvtnmasrJrX9rsDfzwh//iSgMoU/QDfjpEEu6ftZ9/b9Lp
2wF573+4QFGMp8/VpM/Azjr1T42QEx72HGe7/yRT5yehhI2GgFt/3B6a4RigwFl/
1uAAVX1IglEZljHdw3hpJunUHLEXrtG8z0T9EpuWuuh1wkhxQj98BA81EhWUea00
7bXdDL190yeOzgmezSi5Ryu7nLzJQFcTSS4B7oOvbDqLDBYcrk/7HQBXohCdz3Xc
0eGaBJBoZW3LCl74H+LeyI/Fgzw6wKKfYFwlZ8wc/liThX7Ol3fH+339wZHsPGLZ
R414C1u8H/IGGdJemz8Ygb4tRwx7GXOwdZzeJaxMvlZkvHrAaP5p4LStzv+JtyLn
lBoF6iGrV2GO81Hw/uCtMDVh/6cSBARQuPLJi4c3KqvufKL5q5ZN4glVdMCf0fKc
fdinyI1fyoyNhJJuHAYy6ubJiRAIjsQtmsJUviJ6uGuwR5BUgOV0SQYWLR0YYcWD
cXSLLujif46kcazmk5R1nlmdPEIUvs53gAGryBdQuwC9gd+vvFHqsCgEli0oEiW8
jn/werG7v4qH0vYX7HlkudXcrx0d6GAguMMGtDx6dmLI+2+k6P94EbTsuCMsSFWG
tzvN5eE7ya7s46X/IlCjRvVcJyzL7hZU8an+bkLgg8jmzsEwkhg3u2el5nVXQwT4
zyxCqkO/xIIKkjmm698h4GU748qUP1SeGJE5bERUh/ODcLKJMUqVMNSPLvnw2ubt
EH+TBeYym4yryd3omFE4FRzLWC3cUZBBxOSlIsM+FfEIMkGO17bKDX4nW5OsxGr6
q81ugVqVPdFrAORmfW+ttbIM2q6T0UNpjggSBRBlGvvGArEZogpelDMb23xHFjkk
Pbkk8flaZU7W3Y6qex7bv4bAEdAYQoglrDiqTEOBjqzc8HOVQd8F4FOO9r9+RnAl
x4qKILQ0H1sh1A4i9a6RK8PaL3PGttIaiwJb7bZtG9LEYUB4kqUqD5rWDgSJyQiq
LbEQoCE8tiIqtjDwicDpa/tiS2L0qPOgxN/FUpvgMWqe2mAhQ9/xSFIKmqMDYvkD
UxsgmggDJflyKBadfyxmB6SzUGht//+0VszaZhyKrxgX8VPeBw3qdQM7MMcgiCVF
YXv/gRCrT84QYbVtL3IbmoK+uiuyHAfol83bdgvAKXgd5OTgHeE9izyvLJhDCXWM
M0JefGh8QNfecPN4m5sUBQUGSTN3xx4Q/X7ADUvAb3XKdef9w0QqM+I4H2cHEcR9
nin2nLM5eEyRjl/uIL5N2np+GWVshzGJkfUDv1n0PcqBW+Yx759d6m0rb69WG0Ul
0IKHVbM3ViXfAt5XXiUCJBggI3R6it4Ri9H7p5CvfuzHpaIZB6hdREnRMCFOBQfh
yuo2UwFIEdShPsmqMFnG6e0aKONMHGmOjdE3Cn8Y5ryKl+i+PpEBttUiccupI5nm
sPLd167ui8T5jGhovc64XbGibqFQUMrrL1YlK6EJDVrwvNQUj23TZVRiqUb4DGdN
OvhdRrbX5C39K8YMsmaPEIqoqUiiu2qsiuhXztzcQ54BNcThXkUU5UkOkO+aV3i/
ygNuIR46gDuL4dYYk27Ls1QIJeIItpNBV/Zj5dpa9M0GFqYhZa5Ywr3pqPy4AFLJ
rRT8N4fhE/IjtrNF2rMxPa2/WOAcpQXDoTORt1QDBvPK/YnA6Op7KBz6H/+bAkH3
4W/5zrY/RUxsLsYVWeH8Xah7SLBZ4Wemo0BeQqOjkwHnPGWbaZu7RMd+kHJ1PgOL
dXgyFIKS+8V6nG0SNMHaQOIGIY4pbda1Xu8ayDGepCb5e3yKl7MmfjfHGG9CFm7J
PQbA6y+Z8FPDnCn3/arw8b6tR8w7qRyV2xs8Tectt6Hgn5UqorY6tscT6VeFaXO9
GJ+4QKTKk7nUozRoC3AIvCq1soWKBO/5ZN2EfNlsMNvGyzwYLR6rYp+Tjfo9ghnC
2Q1aub6ycFAzWABv8uRFSC+tEdzKMSLb+2ZzBB3MToxtxBsD8v2eyusha2VsbtEz
WdHcyw4Vxu2jzN+7DSh2L+vTmgVhyOmBoNhzcba6O+Q83rNnqZ0/OcTHWiYyozIC
l8v2EqYsAaqrYHBdmB3tMhCSd17hBMAiBS+1+VzY2mVYyOPfachwc35OSA5kmV6W
BsStpTul50fgui2GOhZ64bp5ZfTS/YoE2Op2X47M9HkIwfREmSJS3v7JiZjtqpDa
kz5UV2bIMVM4RQWK36eUSR4W4fMpt68YijYbxArudInVT1IaIjJbf0jrW7MnBXs6
JtejWKBL6D555cy1yxOUN2XzaFDSs5D4adgXdxKANpjYkuvtqM2ybWKr10HIHvqq
AiWqh1Oltu1QUUUjyyGfXIoKipCfOOQsrOEm59qCazWM4mhPrnelyjVCLXfmIPDW
knXR6sTsXvU8bi0XoVo5OM/KebSnR8tkBsp6tWoipP+aToEjJBc+4najiOP66Zg/
jxK3uPpahJAKT7tY5COfrz9/xTJ3mVlCIpahNwEYPYUZfJRytfTX9z+0o7qnQ+wI
rLwZZfmr0pjOWJ7DDbD+77NVOmZACG5+6WBwjLbtbaWqSENsa+sNrxozNabxpd8Q
/9r0jz67pEd6OduomsoMt98xfX+VTUeFz66U70RfedvpkSNxsUvjwe8Avxdcfchk
sk9Ml/mdyACi5jgK1u/VhVO45VlaMYlrbbtgEhaIwQp5K9FGvgJnw3C989ly6RIo
PtXSGh4gzy0dg9KTPCnTptfcaplq1LZUcG3KrczZAoNu0sQ9whYyX3POoKItyi50
56BHGG2FA+5lmaFe+FDamWnUDERaJl9O0vRRApLarU/O9529VEQiK0nlo9w494rV
eY6PF9ckT8K8GWc7Ts90MwmD5SnKXhmoko7mAEYterlbbCV1K4EMy0cKYos604b8
eKt0zJagfw4ySTOxEwpMjj7+6QVDBkeebiv7XTG8R1r3xJ1oSxKRXyWhs/YKH75h
w54j2coet54STQpIsa38NdySr2KbQlCNlFKWyBf2kVd2+pSq5OJ7qt8+nt0Nwr62
fljjMMJQd8nJCXW5aNLBtyaxSgnBd2orknIsZeHczLH2uhXLhNI9XKc/MtFiEYZk
XcbeWuKM6q6ipijeDcb/U9359jTyiQhym2XYMr8UgrMO0WANq8F9vmO+zMVYYzbH
vDgLSA/wxYW4vPNhNaw43ytAX3BRZfE19dmlePAmWyTs10EFYNCeiCULTHq6rUpQ
jJXGTzrYYqkVd2nmbAxS0e5lHU8WL+C7EbRYWt1/z6PtSs3JdAdhqIki4/KWx6Jh
QP34XumKMGmMxI1Rt/YoASWkQBxZq3Z9l7NW9Yc/nDTJNxqa0/qGKQ63370F09DN
Xo7OuQ/ThJwVgqGoa30+Si2SONmS8BWnX0EGjnxcR3K7iO/rzP02jXQH/+cHBZof
prVibIoHrOiel+3Jvh3LDteXj6H9Yc6SyxoWqcf9aLjFUaAu32ieY8rK8F1pWcuX
Q163FlG3tl0R4Rk0GY0jPU6nPqPnME1uDVQ/BJqMzsAh2LpHMNqyet4MTdkdY046
kMcDz8c0v0rhjiNaBxKOfeEYfZv/ixgANioMngg6WeD4yNE4+4V4aDZPBfbnQF/U
BFLP2SiewUbvVCkowDuKaJ5225eooW1ybQCASEyWuRhabhl2N5/llCZXbRl+aRMs
fvTQqpDYsNeiDaLjPl8rv3wWuQ+HaLIfunhg4Vkn+8h5Z6cT/qIouFEC4nUxNU4H
vjeXyZCJ/7fcEQe+KMc2hGy5qRwvQlYcIRngCezaeqcnXuuqOBV9N1R+bKd2l+hz
WCOYKrtxkdGNA7eO3NUtpWLDI6bp7gQqXNRJtKATVkvqHKwKXH6ivUF9eMY3aJBe
gBrCMBZvXMY6oni7yap1/uPwuXLDgELg8gszOMcw5Igs5tfId5g6icoq9wpZ4+Nq
zX2o9mMpLuchlX3NX2CN/iOJVuMH6Ra6x4LL4Ag8n+XPQ5zsEZdxlLcXjiVcVuB1
W4GpO1zJd27EjKuJhcuAl3mvFt4HLvP5MaFYKjZt0UoAEju06x05skAP7Jls6Ya9
8V5SiuOaL0UQXVdVBWKO+M3QCT72QVeh89uv2yIesVy6H4yePKB5HGDHll2CoTyk
dtd8DyC2nNkHfQTBn9VmFN83RIDoMkZQX8t6FQUJ/+/1htqnKEDZ11umXbJfWS9t
CX8yU/jjFQ1b05r6Xqg/eaYUjErzmHO5xdQ4wHoSdwKgfcAgZ2OxxDOtQtRG5r1j
daIl7p4wzEFJCLhqoFt4lXMYOUJEsJzpxEU4096oF4GROgc5ALKViEchDajDCPMM
jsOqti32QHxEB4+gb3tGzNm05iklAKpQ/LVaU5TPoHIEkNtROarPFidHSMRCvbON
OAAE1iVsstLIK3MvSn06KMQtSu0+IdemmxBLKSjEotZfuiqRVJPPdXmwWNSyUG2c
lPgiTvK0RuSDKh//D0sYiCxe1ks3zhfX+8KL+se4hCLnqXD/GnAwKiUBRY3qdjYy
knmfRX1Rw96MkRm3s4yfG53ka6ltAkdX1/pFKlB2zjv/HvmAvEU96oNM6E4XFPz+
f+WZdMocQ7dEnv6D0DPsghg/I1xRCu8kDWAE3XXE/n4QFvg1Q4hL5sDBsGUdNlGE
SnwRIDxEt1dA28u7yltHqmXfnRurDtGP0iZ5QlshPqLo8BCc6uZJkvpmTvwm0VWo
uW26KHfDAEVIUOXcBWm552RulJNwMpx9iHwpe9oKaFcwtvdW4ZSlQCtisPjgESo3
o6MSPKtGXh8X4jOaO46XLcoNlBcc28aMiWBUpGsCAwaYf9jzoG3dw+7p2Ux251QK
wmrBG/ghe7NasjQQNLk9xUguInFV8IIxxCRA9Hi4DbXFT9z31m8md28vFkfZ3nOG
66sLiZAggaRZ7Wd5bGFpH3Gx5i0V0CcRaSFTsyEbxbcwr3Vfpb00VeU5o+h30J23
fyzDyOjQo78Pesq6DCVkxPZjru3gat79/ZLQf0zeKwLBzdypAcgxWQQXrHNZVhQV
EtNdtZ6k4hHnMDetuJXaLM6DOYTi9KBbWzRZva1Bc+/EZkVWiiTP4STwU92YVWrw
dvAp/aGjALEXyQKncgfhhJgJEJoEoNQMmBXUyPIKu+Zaphj6Mxs0PnoCp5yHI8vq
Bp/r1cRIh+2ldhoSIg8Zp/13SL26r6w1S5pPVDG38Q+dZy7GmRYajtgtOYngz3g0
GBe8KXNaWxSq2n4j5U6Uawe+gH6yhoQlhBCLbiQ5NeQpHiYo2VVTNw4JWIUBEhOS
qsGPTqFNhH1HTGaQ7dlz6qTWHh/nmbYRXVvQJ5MAqtdq1higteJIqIbk47H4ShRF
xE9yHfE6sm+g9h8Nqf4h6SRb88UbUsNLexblGmCZCU1ASqA6IFMTyZue5r1MYscE
4vsy/7RPD3uBLey2P5aV/zzO1lGYehCbA1LD6mflycswa5oJuUiyEeiKKP/GRPBx
eWg3Ca5PQDPhL0LGuVOW0OhyXX+GW3BUQkvr2lnSF46Ty8FO1HCKIvM36OxHcTYk
13Z43meO19khs/xPsdh9q57KXV4yA9QdYcWV/O3IlJNdCOe1T74TRC2IbexS/Eo7
F5SjkU03G3eiPj6Kvn0y9yY9eyoec3yV29GOWIrgnOyDHjiDpvrwrBBH2s/jDJnx
35Ro9L5Va4Puj4dtejjs6wxd8ORW1cYBmzpPOEK9pfQlqsPwaRCiDG2vNbre1iZK
2CEXKn7JWUWWPh1mNyqauZcOz0ZPpA85w7kbmNphqzGOStMU/BDq9g1HVgj8w0Mb
5ATpmwV6Om0dEJvkCzwa8zAR1d0v7b0Y51FHSzhfvu2LtF4I5kCbIHZneCwU2V1Q
C/naLBC3tEtFPIlPtcufT0ESAjksckJbZz3qUIUNdZWVOkXXkQiZR9BG/HzijMg6
rO8Ucn8zChrVObrqXbKrgcAcGc4tMbmlzlN0ORnkFe1VoTfwHgcvmesl2WZCaqgI
qqqPp1RhkZr0pArn/mYEeoug2OoF1v829Q/2ucNLkdQkAS5u456WKrQ6pir5O94N
hqPB32tJugyRbzyQEcgfp6u7Sj7AtaquGI3a9LrfZLhDZhxeAXz0svwDzRo+9i8+
DtOq81Y8KN+J+8uCx+Hbb/Ea/32dx9GIWtEBChSZEjsskePx/zfz545KbcuWujtH
TVTyHlrgI5BjYQ/nkwR7zaBu/gJJ3pxoEYH2IDRCCFiZLUYJyD0NxQK1iNtHfeHj
ZnwBYhOl8Ag9XlklP+stHGJo3jfIlmcME6yIwKcnLcYf2JbH3s2LkEPfhHOYQUlx
JKQmu7ZlaqQAZcw298oXnJsYyAMuDXAyYLVOr2muuaiJ0orbpgkOY2iklgPmhKz6
nnLsgCk59C4NYJICOc2VzrywoSekLf1S1ybDYw49XkVFz+QCxPoi1RlZs3HqeICd
6/BOiUX2MjuIFKG66ncS8wZtJCxEvnPrGWVeOfWJrPWYG3nIZyZkwHodspMzNaL6
BuBAbSZSVhRVcwDwSdZTrWJjveNsJ1aAp4I9MNRmySlJJ3sVrrO2oPWYj3xNN+GD
ZrM9dpJmIs70m+Ek2/yJ8ppXx4p1FwlW0DViEGtOBEacYtuENtPSPfM1/avOk8rQ
HtNOWUdb4ZUP8wHzqGQ0OIMwNsfEtqyDlbqrHj+O5WUkLWvTscEtAEuSRU9u83EH
sfAbI72dPV0hTct7sWfsTeLrqFfdV5NOEjTERnzfX+juN1YjmW2iWGLMALupkCKd
6jLyOvfAb8F4PktqAVUtq2/BzTBS0WbybUVp4zmdYovBySr9tBnseFN4RcapXZr/
/6CzNQNz4H3YRbZjIWrZncItjomKLnv77oOhto/SqnkK3fUsmp0MCJHtOIIORV+G
5p/11JudpyF9rWBDKpI7H8bHTKRdKfZrpHWiFkFqqpW+7QoXIDEk+eGxGP32QKz5
X53368N3lt9mGReQpzDLs6YlUR1WPW/DVaRWLcZCNZkbCnRD0N1rGAB1iKup14dI
BEDmVWAr+mZOoFfXg2UHidZdsa0B4BbCCIHzHctmfucAY8PGB1N8/Q9ZVxb7g9bJ
fi62DhchFrvuBHydfaliVe3ibHm3owXpWH9kzV1C/gfPxeWuWO28Ocwqfg9NAwFM
SDd3f4AyZU8TqRxikbhRH9XfTShmC7YyC4tkUTjE1smrgMu8RVQt0dXARArswIde
IWZWn7TZDDx59OuSiEm8gefvPkvL/YZjM9j7Fgf2W7zJRRIkHfm2h/j3GxyS0l1E
QyaaO9ry5202M9No9ej6xiTZNIBMYbeQE7z6vXlI4Nwexq5j5uf9jTzs3f5L5Rw+
0QoELtGxtOEidoFk3PWKkIJVYz3+Aeul3Ocd9Xm1xXZqqJ59ZXkkkhJan43MVWrQ
KQEvy38Xyc7Wa/+YrOvzDGR1zM8+VRGwAAEDZzPP/EcSfQIKs6A4+a/sxYO3F9JH
LiQDnLMkL0Ul0ISVCSLRNQBnuZ68WuXp74i4mCCqbnfUvtS4jMpT75kaZtSVkppN
lCMiPb/F5mE6lGHgw7SLvIullJf0N7Efg6aGyf4n/NJ+xJl+4UucWJC8N8V0u3kl
KwMnJDdBqrhtd1GF4GgNW0YeiR+2lzU4vFSmVrVpKGfgse/JhyEczQe6TJWZv2v/
jEADPZOMh/GkjJnL+N+mTlkvrtoFPTdDZB1+ewWn6WB7/UFRPYMDl5gkpkC4vwkC
mAroJpG9EXYeYyECt7MuXF9ZTHyxtcPd3Y4vozlAwTAZWToodc/Uv641ErbgAwy9
tJiAJZomr3fz8H1qvB94vvyQvU+bdMkO7ZX/GANaFJh2Dhu9kjORUmTRc/yBfpF9
syisqlEgJQy3/hZmtFt6giQrQsEiyWvjnQUlPE2sEW1FvRvaCW38jBsU1nucpxdd
3eSxor73uvfOTjZzWY6IQN2u++MmtliUoApco5BnxkCkeNVttXMvH9rg9Si87vRk
gs7r2z300reNsngLSQD7iBNcfTF3YCb7fkJnbRrUN+1bFu/HaOT7Dqb2bkGoUWQb
XuX7xI80DcLelwYu01NsilcnARM4JppMz1//UfqlkTfgyj0UepkPtlLWKJ2UCXdc
0pIt/bXIYkKww3Df2x9ACU/MMtuCgbNHg78PhUXIY0ruZz0xN6w67vDjaPfOaykb
P7jWElE7/B3uxXtuXwPO67HweKIArUvM6tOdTNy8+dnPZLBXLQu88Uob4yBlubTT
b/sph134WrlvA58jqug47YIfHVBLdDQt1DKQ14dipJH4GeXyBlUF+lle/TOPnn7n
8Dyzd9fQdb2TrQHyE+5eyngfv+GO3QRNXEqqgiKyL3ALBoM2Aa88NA3dpMoniz7J
CcYeoNyr7lc/lV63t3xRg9BRyqD2U5rcCRxAZIpirzMm4G/iO+e36hJXqBXllgwu
rEldLs70+Yoio+agZcf6EJyqE2t8CVaMZuRAjSCYTXEJL66Fix67rLGdYzWsd+I2
ksMcb7N7m/gp6DiVk1gi/nE94sV+2gVFOQTIz0VIdusDEcBlvWwMgEQOeZ20WP7c
dQDvHeW0KmQ8W3z77Ux3P2TcrFQKAS63maytWfNg1c2cI6TFiOKy1Rkt6/GgawiQ
A4Dv7NrWYVEjuUcUjXpoB6xMWLjfkzCyTNFJhvpa1VkrTyjrjuMlxNYwzd5PJVGM
rzCDErrll2JC5XCuV86A0EI364JGTPULqGAsphTPwT/WKxbu70SRTSQV07MY4Sel
zxtLlFfUCGy3ulAxnxDll8FZXvjSi/dlm0F0B/VFpUmC8cHXKrasunq0oYLvZdDO
nSdYCNAeHmHbCEchCT7aVTPN1EdarfWwrSD3ashwomYK5UYrWoAwwe2vhX/MQrdO
HzVe6mVLtrLk1PYLgbbZp0VgvPiLKaEYxv1tYvnPqgO5RH8pYuN5CQmset0e4XHd
L2dGdd5KCcyAkNuZ+uQUW1lfMNxNeCtrwGpWk1BojYbXRGE6Vt4ESkVw8SJtodT2
d+7u6Et3HFi8ugkxWIufKjg5IED/HU+lB14bzUWGpNdu+w/2hrU3hpLaRWrqHbr+
dDQt3obBCnKPOoALlfMJjTmpwkDX3JkYAmjtogZygv3YC9av0onCNCDd88CQiaYn
L/yQkq31+Lk6kmkYzmXEph6lapD8mJU2krnICHSuOzjkrzqKrPEbu9H7EsM3xlTQ
yR5fOi9u4uaQ1d5P5VBoasCrOdAlaRriumTi9eoEY71B30pp8SbZCacRekeE0aN9
vDiMc5vNk9nQUH+qXjZOSQbHZr1dzZsr+Qcj/l8EpQoToG2c5ILUlbQ/Ye4a/55e
3GR/P/8ZFp8u8ajQ9UitgS7Llm2WrBboWqXXa933NE37+/8g2e9otTZlg8FKpeQ2
67+QXa+f8sZHFUAoxxfnh7o6y0N4bUT48SVlBwSHXc2xb/hoqCLNx2gwN75qcW4L
0F+1P9yKp3sOrBGZGBaGyMfAdz6QGVy0WG8VtZ3/AOKUiCUm6xXb0SkTb6uZL+u0
Y9R6M9m9ZDDAfuWdRuCCMXHJVvVBi8gDJthRAlMafRDGK4aaUU9KtixBWj1Dat/x
EgVRiEVlF/pwJsvfhQt+N33twvbf5R4mPxw9092uz2VPNOSO6gy7WSrx+Zbie/9w
7e6nfasMbl632mO1QL90PtxWJ+PJz5NMd3WtDXfM7nefuGZ0hDJlwg8QUR2/shTf
sM0/s7CqJmJlDOHGiBL8wlRuuZUFOocR1IHBBosS0ocoIS7KErEVHWEDW44hzCKI
C8Pc/oinZK/HjwVxSrro/gNNBX999FZZhit3zeVQOJhUQy/874ICSIU5V6zrmq3g
xQwhOMFvUwpz5VgnCGu+5vBZ2GgJDfJYp4mgFpWDs6Mfilfv2psEjPAd9f+ttpEE
pMdeQy99po+jT40cjP6t/qm0ntxqK3Rn0vK8xpgLI5rbOCZ3wQ71BhzMdbuIRitc
MuTgfkpz9ynSND76xqR8RT/+1tn64Hx+isdV6Gw9jDh1fM0FXKreW2LBDnraEHHp
uCMI6e/keQ7BX4gCKlrs9ct7P8kNLppUbvxuyLNpGWwao9+IwgsY7iNpXjy9CtxA
i80f0GlytA6bvL2LH47HJenDxIIK8edmNNtYbBctC1XQVTOH+B0CDCX6Gr+yO3Y/
ld8+kVECjc4l6pnCqjP0vMG20j59H+Yrnp17mkUVZDaQZ5BEwRC60Sw25UnWzJhd
1xFZr0poCZbamLtiginclh7RkfgfoL1h1KiU4nLTHfu7Knq2kPALRqFR3WM/zhXG
+Cu4CjjLc8CJ1tiazcdm2OWV4jV80rYwt9NCr6ZHu0qiv9lxRFOGOFYRzFG6bbC4
ujJ1JgSPDe7g0ozNkhmaeVLAPSPVeRXwF1gCAO4tOmIWJOauv1QHXInxMYTUSGcV
6Rlgl7tuyajzTCELCMfsS/Xj2H77vWuW+uL1T+oODs7/LM66VNsSoGiYsZYi6SZ0
3I85pRLFKiRFRIMYOlJPFy4f/pgTQ4zleNgYmn0Ic3MoDC1yOQPnNcjHS5NQ90km
5+Ry5Ab2EG+m7dMr0Kv1PQS68AnOPhk9DQBPuXo6BvKJtIQCPEjMTDuJZDBqlwXo
HFdBqNLLOs3JUtFVWAeimiUH3ST3Zvv5eh91FCoNA+j6h3UirMz7EyBPKQ5gd5+R
kJ5nW1bDKy7oR+5oRkCzz/MxfBy8VhvUIv8wEodTr33nIwPJDkQGDbJE2qzz5Itd
lgFu1vXAb3XIbQpcNan74JLpTUgwC5mS96qgk3wNF3cjZGvCFAweEuUFGB2Y/dFS
YN4kIeAm3e8whqakMeIrW3SyRX42ajWdXBQINIWuLMvlq8j5WBXYWB2eFQofHaEO
imgfeAhHJPvzNBaNQorIqCztH7Yi3x3s6JAnXB2hQPu9N4AlVSIdcZz7mSF5GSt8
+gaiftCa7z9wBvIxquAuym+AjvOPhd/M/t9KtSyQh4FA8gJ9kNb4TvCAFC6GJfI9
LExYZG5tiUXwSv9vx9zQrJ6tIQ9ALPUtBdMvxiDhcUhZGwLPP+aPt3xpKYkvsM7V
V5OIfJhbWZru8mx6aFrUtrg+s6H8pRTO3HrYDvvq4M0ZjlBMsPXcIm1h9Jdg/NII
f9k1484unLF4A955Iq4Cf/Zkk+YhwjasXdF6tPekB4xEr6cpGeQyuvjS0YVNRsWH
/QOSoiVK03qoknU7GyKk3NHYIZKjKX0AkutBZPHHQ4t9+rgUC6iOXQY4QrWsz+20
4HEkAbQb6r4++iTGwb4A5lZxKzdsoQrt2b3/hGa/MDLAUsWfBcEouF3oXWYH02U7
oWoMJx0UTR5hHoTv+ha5zCpkByi36tXbPlcK7pxX2UlSeddkdW6WjodJgqvJiz4I
eKVSObXZ5up/ddeCiYqgQ6LBK2HTtrjdelcJk2NMrsPB5ObKipAJuWNPSI/PfIEB
mRqUscDFpxjBu4xhgqsXWoxekN4z/+ljQM+srFNWv9aDYOZpUSJUa5a6Nww2MHNn
zCT8v8cA5dAh3olCUN7nKXcVdD15g4T5BGpojH9c/yLoUlz8N2DxssstNp6/xI3P
cuNcziaZY4Aydpsc28xS9kXveEAz6SXs8wN2wC2Vrqw74OPZ0eYCIQM1OV5GtM6k
EALfjxRpB5XStMckUufbcIyvYGSq/VlCAKg6I1LHQ/R3SvrckMHknWopZxDfNSUM
bSUT96oxfNT7zjg4G3s/7kWGuii2rgZiSAWAcENn5bV3VH9SINCH8p+uIzx1n42c
rDI93fxAbBFarlKPzz6+Vtlm6zzZDfowRtsRrx4kV4g75CjLF+TilY7yuFtH7nVF
/e83vgkUuQCpuARY+5EgE2m6lK+GOmN0Zv0i4mFCvd2nrga3/joCx/lkE/vREAFY
DH9ntznLydD72jffgYHCZ6GBXyl+AzRSm+jHdDLlOOqSU5mjYMTuDeXJedCNhZJd
AmVUFRG2BKEjQZ1p0tmoZ9cQz7pnJTDnIC7iVC4EFB9WuhstC8XpE9KthQg8XzIv
hPcEQZtuNN73tQXN7g/Q67vmIGDCKSFz51KCj6KFQ2fcrTOePwpP2yOhwQhRYq0x
KPlPblmXtLx0vfPhKs0bwQRTDn0xdIMqw3SZ55yGyqMlnRzImZlvRVdck+/CdIuG
npsWlj/5TeZ1k44g3dl11BEzyqWhJZCn+XxA6pjQrpP69Sx7x04k9hc+8dcyI+Io
GEKINWiudlN4s0Nk/mVjRsdv1EeedUM4wsZ/jfas6s98AjUQL6CKKAtL+NUwPA+C
QqUhh+eZ2vswEb1U1MpStM7U4h0HWtuexKX6Tiw/RQGuUISRxHk0KJFM3xN/cYyN
DqezgkWMPP6EMoTtCdnp3C4Sfc+tYd3u9Mox+W0Ia6JJUkuGvEEpTL0srefVd0H3
8OBDpGM/Yjb2kvkcYgjerAD4jJe9sUoYQj4VtsON1pxyhdtUDy0Gvy7vnNHcIKhe
OWsTMqOWns63Q5ryOqZDFS+Qxy2OsJxBkiEjezzFhMXl3/22IZ8XDkRRAVxYEifY
wU5snfFMa9aQGFoSWc7v3lCN+3o9DgO8wfv+XzWvHAgavkVAnK+8WRIuauZDY5De
Zojq5AwnPOQ/yFGFt71YINJtaTy73szKyqIZvUfbfOnyD9aKFmkEXvqvXkq/NSqQ
LUYBJlTvU6sKnbxt5ifKJeYNyYQ3h1SvvL9S9XpGZ6elZEYYBP61ZJYY+akyet4p
ZdQ0mCxyAfyIhB/VYT0AOlLP7fYzSYKU8jljG4zr1FZiB9bXYM4xuFRYb/Mt5Tan
fMloffRvxATFlk0DkTSR6z3IltO7vAF71Bk3MuOyMBv4FqW5+pICuGfwcqGqQqpN
IbePJI2rJJV/Jv84+dRVNAA6Q+9bdXx/d9PVsRms3U+fu1hIga4hVYRyux+NZhFU
54YjJZVUNeNc8BHMHnskNwp+2uwTyQL706s7Ds9ExyW+GJK0fA6bL21xhnyzPywu
7t6AxUhjRL5lN+2saomQkpIn+2PAU72lz/IeLnqa3GMaay0jLV5tIHTRc76fRYAz
3iUeCMl99px8IXtIEwyPQEFKECU7HxgH2tMoIxM2h7/UUJ8+UfP7DIKOXIuioC3k
kh+EdanK6IYre1jBS3pwtcV3iFUBPx2AKvXSrmHVOW9N/t4o62ryfFF0groGhmJ6
Mqb4lmSzdHpUw+WVuoHgs38dBs35WSXKOr3MDdu+OikQ/8fUETW3x/MFIJgJiiJ+
1XK4h+A+3YA4yeG++4L4BdlGXe7mU/WX7aYfn77bnui7BNXbciQbk+dFjiDBhvHo
V7N0fgE95oPhB6rxAm7lhJri7ED17wR/NpBLyglswIjATClAINkaLLLhjUaphNBQ
8DsKXQZeWjWtBu2qV6NCotSTSNIepx5tGsvDSYi+nukVgFrE9J+Ngy8HjuGgLtuf
tgovd8nz92cov9tORsoNhJ5mcNiWL1ezPMXVbzU22sOk3ACfmO0uLf3ccuMZKFFJ
bi9ikfQL1l06Ir3EZde09it0x5hcBxdQqET9Kouu1/ATxl7TDH7QhKFLoUZi6h0J
9xsebFq881BHesMEdcTqbymdauOYRgAoMUeiq+XKqPq31VSTVubbSLCF4ngKUUhD
kjFhttrSRp15yo91hhayL393huSP9UTW0/yfCivL288k1iz+x8xJ4i8EFrHg0ZhS
4f3GuZWVEPuX1Y6qiDGs1KNylRUXEQsPAA130DbXiHFWw9wwmfjSs6IsfkB0cEBC
+O62FFNCWfJjjRp7Fy6jlx+6/pMz3mkGNIaLCjUgbFE+irM07M3PxHkDyP03VefB
dAiWB1t91qZwucM+d1Uh/2D1P02x1wmK9ZUVXp7ruX+8EQGyJrJnEBNaf8XBVc5Q
TYIK9LmyNlV0iip9EGwkPdYhIA9yaXQfYQRir1vX5iNrknkMCqP/oyYwh9XL6cBO
4gPARS7VI87wmZMN9LbErfpis4ks5RpE8SK/cPDSlGm1/2S2ko15Ikjpki6N+1Yr
G1ZgCXRnNvfU+EokyJodhswT8evsBkOjUNq3KtbtIqQODkKWOj9BK3pVhpiOthUT
3JDqBJ0U/he1zNN+0OiTuapPf11n1CAeGoGrIbmvtbYzExgdq5i3tDqAhNyvVtkz
BcE/4jIzvpq5CghQz59nLZEqDsZ8rOZqn7hfpXBlug35y5UxEayLbtS2/Z/4fG4d
wQwGopcaYLtTBvh9WdVsPxeCt8+fk0sVxAIpkknaoCqY3eLinv2hO6Fm3JTRX3Mt
R6wqSW2aT7Tgn67mM+CuNTCdVdrddYkQEZvxyBIAedZTy1SUNt4xwnK+Qx/lPwpI
3/zdeiOOd7DfagnL6FF/vRn+tlB/eqmCvzux8srhaaEVaTr7mThrBa/AwX98d/fc
taY8VumjNGUAMmmerJp34gwiOtN7X0E/9IekseTvD7Lxi0Yoan8AZUsfptV4fNjW
QJ/NjinzpSlWZs9BLS7Ie9HnFTXtDzoYUq0/SiaOoKvLU6aAS2iU/8UphjaVIPaN
993N9tCPErNissL1iPN8KulHhN07a+J7zCown8VjNoPyUuVVQDKBegCwhEFVHUWb
mJAjJi47xOVUPOWgxfAiMSZHuiwH/cHeHlR/p324bN3UWN9QfaLYNh4bPpqBd9WR
5ufm7tEcgrNCWftJuUvKhbtCx5EZ528JkR2ZWq1PhsbvbTMmjuuumZl8F749fRSN
5cHskfr8J5+ltmIiVXOf0x8ezTd5z8Nr86IYixpfw9ugsWIky30qOmrvptG2tajJ
Ii0JGqWCk4jG4goVKR47oyjoI5j5YQiCFD0iLkR4IgMdjAbctakBjA0iH1CPY8iL
qrewQpFMvLD5yYfLOe64i4nMcvWpEB0anjroK/ws8nK9YNj6SSH+GkSPXcgKxNxZ
7TsTgZ8vHzKTG+EX0Cztsa/6wNLZCStjvDRmwyajYU4/69NDy9RNsB2wTkgq45Td
xyJA7G7nGFARNcgyx4U7WVsm8+hAE37csie7GaMh6OdeS2l2Brw1at06pYIfqNbf
ZTkeuLiLNKgXTZv1wGMcRbIJ+yrEOh6k2KncRaqrh7rI2+Xuzwc5GajleFuEUVQS
C3B4etWUXXmVsY7zFGm/j9I5x/wNoIXGpHytotyVe2THIP+aebbUg0iNMraYSNkU
yEto2Yba2AbtNQpE3pWckMVGi+RW0R/qr92hQovhwaLUvmFr2NHpzHVxgbvDBAbu
P6itzr8X1MiZ7Wn7gM9XrvPujJbR0e4o99LAD/7g8t864bQ1+uZOYTBgnFQIAIHS
+BOv4SBJrJH0tMdjsEjq5dRVLVNkUHxqB9sQVp4ljHE/DjGivmdVYwPlnGzxJdx1
SsTiWkSBOk/8rsu2AvhHEZsr+/Lfwqvx7Wo+dZqEih1s+KNjCasqccCPQLQMK1b9
l3DN/a63Ldsa51qOntuP65M1fPK1+t+4AuHfB+PBLhMRlUU6dFbpCb1//sDrUNcA
Wf+rPN9Dh9MXGZe4FcfP+pl5DB/j1q8Z+jLJayqoXbs4dGpRBWgq8KzS0vpUfAIS
YGpretv/zUkEPkcpb4uk1E/EIgP/qN+LTFiEBZwYpJEJWzUlOrhYZDWYfW13I6xO
xOj81EBw2OcmX9gKSWb45yYGFh1+C9rd9+ad4y9C1Tg7igxT3Z7je2gLVjfW7npE
kkNz+4bZ6KHF6D4PgOeBjuKFR0elIQ8wbFO4DhyNubDe4N3fokY1bHBg72uwEziU
icdP2hvjuou6lwMhbWGZ7hR2Xwep40bK8NlpbFahGQHwxnnoY/uFIP8TviNVuzZ/
K/uaWtsqperU9DT6bKrFjepYovRJtbF6WfPk2WrkE951m2YDGcAvi4KikBjbAJwR
8GdIRl3y5fazsTUJz4mi9wkOTdkm/JeBX7E3nLOkp2MeZB4lS+8fIFJQTW1jjV8J
s1iD4novIXvvIaRTzOx6QX6IA+J1Cb6l3jVO6xC1n1ZDNdwzEgvmGqfwOoflZr2J
me5lE6Q+j7GYEkDviTjO7i71fGc0ciHSztnUSQ+66iVHyPRfSTz/JZAk28sKewhc
hDWbXsmaKRybml1W7//+47xigugX3KByd8dKimmMMh/MsFDMuofRZLomLPp6Vvas
F1xOjCTfbiZ7ikuLv+FTXcqTMS/XGmYQkHPKW9Ms0l6k3CGYcVYPatagb/hUAwZa
45xvhV8IGY79FFdQ8KsjYuXRFI/GZFTXSxpsqFBVBBLDbBhYyo7+TQ+XxTXMzTjq
s6Kvjtv/ZFPbQ6wXY7sBs9/IAYSWXy/8smLQ6rymW0PxIkSXXmOGJyxhClwYFyfv
asIftXBhmfFSwiV74D5Gvnrc2r6ffnZeG/g6gltwYYJZrgZSQlVXyUB//DGt060t
7D+3QXV2SrrcqUqJDBbjYAYcEXKEQcduQHt9n3ZuIDvRf+3WW5/UMj4odYuRdc8i
4hKdiRJZ2I9RPlkQ0zH6vbtshDkfQwCEpttHfrmXFvY6rXPaPJXiTFZnCtEulaRF
hxcWLNoetAWbs9NFN7UsS+WiIUeHgM/9B5I/Je/knY+tqlR29K4YMT2rzXwHaKi6
8SCM/t0bpqyitcWPfs7kAYk1DXWr7TRK9ZOmO3Moqwjxx/M7LNqxDiBxBoT5ZZUk
IeaIeyBfSj1Uv22kK367VaVrvt8FgE7XGVUKW5Uw/lLImSPFPoR+xt/c3+hRQ6t2
0//fGt5VzDnPkq/81HZRRjmAMdBNXmlB0axKXv4zt7KyHmHsyQ385AF7Sr8BJGLc
iVDVSbZVDD00kU39NoVHrwM7Kj5ECQmNrKyNpmoIMaDEtS0f7BQuqNxlHb9cfilW
PWv0ftow3b5+AqtQ865jj7/K0AnJcuuhW5OyV+QThnb2Y5mI4ZK0cQXPDRr2TEAu
JekMrpqp/qr2/o6KqUOKBeL0hAJwt23UVQ8q/eUpz+7vtCZ5jnw3w093EKH1kdYu
PSUfzvP/a82+T6ZxxUi9CDxgg72FwOS7Kr0Z5aXlxlTY9qUL0VP620UIDTVkhc2p
a690JGIhy/tSKBJI6Z0mY2Pda4IUphGDR54+cLgrJxFFuS2Wf9dfKqg6Feennbhd
+L4VY9C7uPpUtrfjpWXTixTeP269zuchXAtqPotyGJFEzaQ9DNNDctME7RxI+93q
husBXXzuX7w0o8dO2pHdnFe1TCKn2VLVKvDO8zf/x3X4K8j0AJPT7MdIF5KeQq/n
9DKmO3ZkkbwPAJiaEKc4VRivnRbRBI3PawreKjWy2tn5RwQwF1aiCo6Oj6P0qnGV
nqrKYgoT2gqfoMgovRWd3JQFshrjrr1SknHYXNWAlMDpu+GM2tcXpJTB4iDftVQ4
zXS5sRrtj+SrIHGnZRjZaF8JhZB5ArEbrc22q8ETmrxIeOy1Vkd94qserWqcGr0p
YTAChva2MsHCD8V9hPMWPjqhXG8jTmPbPrFydjO1Se0QmM30Z0IH3Ggkvas7w2Sc
9P8/i4eXX3D4UgSRc6g4MFxyEXvZJGtuUb+itslYWss3i4levuuA9s2EtEeqcXZ3
nLmPb4IjeJJxL0pgpEtv9o3TDwmQqwO/94EO5uHbljpgjwWc7pEra7jvSUIHb6+q
vlsdt2vPbcgsXbU7cHEfQ1174ixSxFChzAVN7jqhp4MekerLZwRJ1BfEiX4kn2Z5
2FySV97l5slLjZntAzMJmsZIxIKOzabuaqjCEh1aKnohhesYNZeG96S0ABGC2GKv
XOjuK8VwRpSCkkIZg4H8OzpMHWWsqjosJ10dPKAz9B2zkjzbv5Apngc9lmo27l+s
ypP8rbeOEpGcS3cZisf8nILN44qBHS4mFRz/KMRGgphu/x5krxnFIThqFl60PnBW
WZ9AvD/oDYqIpuDwwg2rujamzO8eNRsDUeM5Vg3HU7arAL+VzYyxlNsIvu51cbsI
76RNVGlUHOHK/+Ka/uTwmgbQhY6E1t9RchDZXr/FbhWjUQ5o6iNX/1/s9f6j+wFu
qmeRhL5ftuo99rHf8JfZ5DI9KV/N75Jj67Ok/z7Qve+OCtfwoV8wShI4uC79x5iu
Gi8+DSlru3LHhN9hSEiI3IA0AmUThl5g2N+Isn0J0e/nCXkmwm8pbUFU1WDp8Prr
udVgZoXTOP+X9KzIQ0v06lhu09r/3VTeApzUAWACYfDWh5kiF7R/+QtwR4oBkMt6
lF9uJMTtfCZMTC6sXGQXFJw3ZJoJ9WNjJliLhgxXWXnKTk0gbaDRShAzQyBTsDXs
vTUlURpkl0WqxmzdViqsYTnK1POESPbUb7+Wo+DXQceFqp1/Wqq9EdrKGRhVqYB+
YcAx+cj/ELB7WjNqdvZp6lzLGSTZN5FfGNFUKX7QUR1gSTR7T+uGnNfv/G0EiAkJ
SaMHGtrCdAJAxh7+2Z+ztcz81wzRCUQl5CaJFY0wDNdpZGozoCQiHoPuZ5Q2wqZj
KD97tEVV3tcUuqza94tW6sXUP2K5dbskDnjkb/IQDUgpSq6WLt3NOujRxs9LXq8l
p/MK8DV7JK2HMsjFzn+H0vKRvExMgrXXKohfCcLQVhxTEwdVdtpkUrZO47cUO34R
ZHCVmCKwu2XffEbwl5SP5dDqVo8c7O3AZ3TVpf5tiIGANdHcdaqK8xApSLXrtCbV
/o+ZMg+CcsJZsUkSbEBwSVGEunUy0O3mE4YG9mqtmR9eJShB4/mRpRpDkkWdPWd/
/VaJ7g6K+KLgHxxK/I6/jtMD09U0OhL6fXEs83WIKILGmGdZkrcYF4CffQJccsTP
lHHBTz+SSB3BWQS++KnaRzrcfXEfwpawDFd6Ta7ZYtJimRuYholH1HdcqoC1j0L8
wItS9mfWaayph9EAjbyWq2Vtm4ly4Ubm5vyPPrcJ/8trY0cN+jupkvIsrjKd/OhK
WsWwDfJUGSUV2qrcrICfWyDHPJU/dq0Q2Zbapm17LbJDIRO8xvnYb9s3rNynUJ+M
gIGCAGxf2pLxYlr565wmOnxVkROZKnz8An+XKzKhcWDjfTLxWiPEY2Gn7/8LYWGX
EEsw1gU+4tlysY0keEnkRubSgGhLqwJz3vEyz8ibGbvJjQDuHiMvW/xjO9AVuXwD
a/1h+Cd7EwV9jZXhQ7TQMD1bzcdF+1+lZ1ZpoeLnKmaA95evxjCzJvIf22qmYoks
44SGEKTkyCrDfAA4OFbL/VcB1NQc+r+GbuIYXxPk3jK0Wvrce+KKqUgsRu+iUeYO
Bm47tNCsaTE1EnlonUnU445iD5FgASzghf8zmCgV5sb2G/2OLN1HqKHfO0VdWDCb
bpUDq2sNjR4qLBEXL5fRP76FQImEWpw218XYk44N1wgK6V/XpVpWGgAcx4VnmOcs
Sdt94Iyfi03S2S/xHBNcpQpjn5JR/sqkW5TE8JtdV8c6tfAipAcl6vMnJilke+wf
/SJSQYWOhgMzb4vmZM4qdI49SJmRMcZ20tXMqgf3Qpyy1CbKE3Xw/2WCo9kPHUoV
jgeodXUJgiwTB9/AI6iDI0urp/0NlVJxzYtdeQDQoz4PS5inFCNCpHECdBR/9dYf
y/NbUOTX2KjMtxvmRR2KLcD+N0fH/qyHNLTcaaBrS1o22oBAwtBYw84ErgUE8OR7
jG6UZ8qIjjDTWcF48hFvQ40PmxVYaIbDt676dXklb7aWC9IdcFFsGNyB5XQFkdNF
TShER4DJRo01O0Wf7oR6GPIYS9+QJbKCmuVgh0WSMG5OvI7lUUUvM/MYSL0/d41n
2S4fvhFIpVXitQKh5HJH4HOvHg80k6S06aI+YX1ni7zHw1U4tbhuokF72TqSXwO3
R/0qoh1jgja0IVfr3GfuNL0HDHyoDbbki9o/5TVWp3jr5zD7YGs+X9RS2dj3PZP4
3eV9F/vlKdEf5wK0+ItFfx5DrMSffCXbm6/k9KLP3G0B33atyjr9rrM+3jvp8D/i
F8tEAYRe8/xYsDnTtmMA8ZX7v+lr6NNROroK14LU3MrqpvqGanVbJ8OWzVGWy8Pn
aqGDjhIO3NzFWQtiIV7YwZVNJoEdtWF5plr0qyXPH1qaiocO0HLwMUWP32+WwiJA
YSK92qt7L3kmNUgm/CCgZKe5EAv6Y/1WVAMDaBRkECubHBkRsHVYLjRic+WWKpVN
uSlAAyliv7OEhmPGOIToIpTB1j15uy1VVBvB4wF+chSKxgf0HGMt+J2qMX0HM+pt
tqNyFpM5TzFPo0CLtUzI3ap6+otx2ao8kkwGLu+lmlIMc5R8TmjNEIbW0rN4qeVn
ht1b1U4Qwr/bnrqFg4UWaRKIEaxsF63AvG19Svdgga+lfTcypPJ6QzXD3QtiMiHv
zkOrHlEB6QZaoyO0Up9jvSI/7qTzI4g0l83c8MA0juSb1+TlV/zpt9oHANm6Bvbt
sYI+dpeaHRi9dP6ofW2KZh3RR4TnzKBTlV7SYaClY9cqzgYghXv4lC9Edp7AKoxS
LVyVDlhZesYyoM47W+UHak1MKJYHv6oMpzLOAumEkicuClsDbzqgloaquYFLmLIN
OVEDLjGvdSH9fa3c6d/GiPJT06jRZ6ltmFewAAsEs1efbnoJ/17TD/Rq1VFxbcJa
Z2msYpN/MRRZ5k6MBm0StNTBUWoiJ0vDECL8ywZyJ6oDUOA65CJRtHz5snhwPuDr
fL6RvDmpaRFY0yVsXm9Dn6H60wPICE+laM4FqAvsOsOmWD/FWHr0uo9NTsHThzG7
be85gj0ng1EbTotlmXYFac479zH+K9NDAd5lDwrbqycubmrybjbDcixt40q1BhDE
fyceXaE5zmnuFEuEEeh5z7YqjUewThQzZIqMRhZIgzQnolqCiUSgaorD8CxIbTSv
qXth+XjmgnPLH6M8rqrC+nkmsv00Dh1GaqSzH4nR9dI7S7nygfdnQ/n6fIGyI/95
IC9yZZG3Gzul1RmnPq0R830NVKdjMGoHJZTm7Q4BAqc7EfQEX7YFEyGmHKxNMvT/
gvXRIE+d2jWGja8XtEMptBD65HjpX2aHhagPvWbdCmRWAbKlp6+yrk9HErbQTTlf
iXggIjc/aQH0ifx8SvaE3Ka3MNcvFPuRjwMa1j/t8LCR+p8Os/UpbI0FJ6UrJWas
qxpnzWKmWMvaBquFun9JtwR0K8qur/y7WcGsb4adOpO2RVz/fw/R8houSkO/YMIi
MrHsLKIXCbsdOCe2c+3fVbE39O2KA0hfLZYdBmOaLniTQdoj6du6w4YP98GU1iGv
KOPyG1qSndM29t8xGx84AtZVbIEmu/yALs2meMGuN+fzQa9PyJ3ILFA4o3zlT5Az
Ewg8QxaeHIyZAcW0WDs4SMVb8CrxQhZgAK/5sd8JQuH3ieL96+CC7KJ4CPde+eWa
ctQp4MxYeIsxUrUnwSpmREZEujILvsZH/ISvcyU15lq3WO/TC5ZpUyuU7VRHV7jY
GxaFdMoPEBF28U2YZY+L2hAk0DtVbtkKhV3DOwbb9jILIAo0147b7UBIemPzXeyL
Dl0hlHYl3QOG+V7k1aa2GSGAwr3n5if3+5S+iviKBVBiuJ00ZiwuSWE6SwDqo0Xd
ttyWS9ryDwJ4Zwc6bhLdx9k/7g4pTcHJLqgu4P1c5Gn3UwN6slSNLJ84xOYCg1Ol
DoALgVuOaqfJVrzxT2w/Ty2Nqvf4WanT6AfOfKU3KPZAIGZNjOuP+ORmHNssEAgr
MxWVU2tOUqUXT4H9uf8rgkqWJErytfqnD514cTzm2lc1m/0IW6fkmEvNCHTqkSCd
LSMVrD2EmQvrWKkUPQ9hO/AhzByxdOzdNgwFxlCtijp6hhZ19CKNWhB+U5EQwF8b
jG0OhoBTJMI4FbzBq4UVwNS0JLiMre8gJDd6E0g5rPB+aCWnkxrsC83tOWfnoNKh
1/m5F4EDwtCQKFOtCJpRWKE719UyAo4CS77hsHObyva2B+uuNl3oxtPauNUDMhsh
7fmkRieGwovNbXcu0lR3mcv1mIQSYxq012TvZ9ZErUUPAaSdE0Q5KwuMU2qC1XNP
F3UZKGa5ZF+aKnQfXH0+9ODqMlpfyRm3EZglpmm0sf3qJ3LPHzT2Cda2enpVtaA3
cdbhv8mhipAy7bhs/wrhFM7V6PaDwjIaYnSVvlhyFsJR85t8ytE4LXdUOuSf3gaF
GQKPWKkfXuXJqwFzPj2hT4TcWZ4RlMQlsFjgS4psZfg/FEvswe+/3QhPvE2EVV93
incltFassacGu32z9LWe2k5ZRNlffST7rNioXz62XJger2bWjDTuF2S2FLiRaFyu
6b/wO95uew2Jv/Z9ovjA0cVo2ZCZhdgJakqAqEQZZEdugWfT+BFvxRpiBusM3tzH
meF4O3I08fnxynY+Ec17Q+enqgF6nZOAIpxTgpuCZGSvBmNn0rLSyFkzPHcNYmlg
k6odfk+ECw3Uw/N3YBtOkJULI9ECEfK8hDrIBWVA3hrPxqjBAbVfmfkubOyhfZNT
9FXnFyCgNFNSZMu4ypS8LAvpC9efPCkxYWI8gtmPrB1fPgPAXHIzt4YQNf2ripQf
hMmO9ePJ8HpCvq1N5S9W915A6wWOuTPQrX8titr6RJhemrAUv2jhYE58uovR4orB
cVyWFa+jaI4JhbZ9Ojzx3JbeDm0qSO8ON8j6ePwvh56KAQALg2Zx++nQJYHgHy5Y
IK/L6lHuVneMZxUf2+hz5+YPP4HiQtUgYQGx+z2+l7bJyQQSbCcgDhQj5VbS3/7B
B7fvNUYHF1sSh8sMaEBOxKbP/iBUL1B4eY+eNt9rQN5Mh5Ry1d+2qqCGguWQiDyE
Nil7DaYvcbRPq0zJy/lSJpOOwZU/8Qbb6b8LYWd+y5zMpTvdD6Qu8t2D7hQ+neN/
KEwZwQOKFtCAlGk0Q1+qMFkr4hsUBN59TfgTkqFZkXHYdRPidkPNu1b8FUjNObFe
22kmLoogEj713RtUlBG2AknaejDd9lTQ5QMEmmqLKvfcJbrKbRqhuXEBMWTy4JfR
/AwH05y3JmQGw7S+ajTCRfJ1Y4LtfVspZhMrFOahUF6bhvaj9lQJhGUwcy7LbWw5
ce0V/DayTF53NQPWy6Coq0e7aMNCKXpW+QKNcaSM6Se+KGx5Dj+epwOLjn1JaQgZ
EEIqDWMb0zqAMt6srHvjsiDhSwi2n9/uSofDNNICbrWfNte0EXTMqF3hOxEVNfk3
VQRFIm0lSZxzvt3oliNczl0l6zVsqfB/mDZuu7Oikul3gaqZ8y2pC/59fStvPPiG
zDpfubNm9rpctNt9C2CEBZGGl6ZYg3gfqFdBUDfsy2EydikakPmOU9VtJB9zsI91
VC0q+TmN4zWv4uTGc4dan+F3kM8Nn18u3FFXgjQ65fF41QiV/LX8piw4jbDh6pYx
gn8KgQcNOOLA/pPxDWryKifIa2QX1WEGotjky9wzKef5oII7jPAs2PVsq+YzG8Z9
ENP7q8/BSaFvEtysMvl47qFhlLTQ0f84UaJWv7zJ6gZTUHX7Ts4dAHcnY0xWmoGk
s4IIHXuY9+khGyHBQXjy3hnwulUwMrN8jfB2bIOXSFO6Mg21K4+C7GIRIJv25sgg
O3CHnyEf99I9CLkE/j7WIgBnP61SSlbQavd5enBNq8db04OXJiz/Rf8tPfvYaocM
MsWch83mf8CA1STIAYHyL+91yPGZcQ1+g9iczB50uhbTnJEmohEa0Bdum+sa7FUk
J8qju+bgcGG1o6d7OBWg+vYnQNi6HdzuyRaWkZOMZNj0NRzqFoMx7hVvmzcL4Q75
+j+XsTLbw5H5lmds3YnOHc9vGJfBTCBLD0MJ6zL3NVh95YZOn6fN9wJdhVddPxKA
OjMqpE3r9PVVtzF+1/6xCPIyjtBI9WIJK0WQcXhQgevLqXUQAd1HldR6gGoV8ycW
nuCAac3iTWevjY8FTEGRWHhDKmJGkvKjIqUlPgGswh2JZrqslifB4QFcjK6YR9v5
5jkbp+FOmvCctXBCHAY36wk+HGPTJo6qY23kiFwrDanpATdTuAX3AudzZWUa7Wgi
5Y2+AWjIlGEyw/1r6DPvPzVfJdNIVOL5f/8EXKS950dHXprf/7b3fycNdqA4DsfG
+TYQx3MTMSIRmmyFuTZy4v3hou07BwFhLpLJwob73NCbOd9/AqgWhIhtUYDBj0Pk
1U1F+6jnrX66nYyatZP9dSKKLQw/POuTiB/fQz/dkoGCgDTo/s/Pg+gfEaSGlYr3
QBBc74UpLMASwJxjCdYOfcJTKZSSD0IHAi3s6mkA7Za7VQlVyrSsIBOrO9HTw/Lb
goVNxsQfjNKK3ayTNaZuQmhBCstM4At6HAPGnoOrh3eexBoMM+UvCOxaQI4+12JE
Xk/LghEcdaeAvAL8CbWlj/GkOCNODbc0tl8EwqXPWl6DBhX8xzd7wrcbmJhDUR3C
3ePamrvux2IznKzsoaUWKgHus1vaEk36ojpGE8AY3jS1hel1Yb4Z4YlqJKiuR34a
N3DFF3XhH4GCRxV7646uMMmBpuDZl/hcwvk6dcufawquB6wjfCUhTS+H5Eg0WuL6
rAHd0B8l8b/HBAyyykW14KBjENf49N6TnPKuiSeB3tgAbLGYCITFAmb8toSESxn3
LYceh5xmW/dWCmhP8KukVMI/G0HmsXsQzLGszGNnXGMnIvh1zQ5RHFfEieAZP/67
MBp91RtyuwA+Unfo0ieEvA4f5twPjbFC6cm01+DenrCg+In1/AWfF9t0rrN4+MwQ
463MfYc4TScDI4HNPyojtEgi8ZYZ8/fQLKGITnBr04JTpcsfL+BfuFWJEkBxupuy
7vaCJWF5Y+4JqcMI46+hJCP3TI1l7m6UANwtR5/FQLcbN76EVOwoe0qWvHxtj7Xu
XpNK8JpuX9zIyBQT4GWeQiLDt0JJCYnZXBU01atFe3WLYbnkfTSYM7IpjB5/2Mve
ogdUJ62k/LWpfcimV1rIqS4GlaNm/Zx5f4kEyn40LPc58CZM9nnZjhQ3vvN2NoeL
blnxcUyzHSKebnArEutlqLSFFTfguqP0nYtBHqGi1/s6N/BfFOJlrO6yiCqVfGh6
/X2rVygOIuuP6g1XiGVEk4rhu27T88auzTHv28AYa13f+kwLH+oHUL0FnPCqHx8E
w/zc8YjM75WiJIov5c4JBiHn7Q+qNqC3zdQqdMtj+GcS50o7i+sTNkjA9tKyfnaT
p9kTqoWSqwkdgMXbC5CFQgaxHe5Pvx+sz6/xa7T8B3E98EoBDNE8j3qupqEOJ9wr
8RHA7kYa59Pu5CtBNVAu5HHL82oFEYApQGoHMUVBpO61eB4+L9kP7b2AQbyNnNEi
6LZDDsZpXkKVEPGS66/QNcoPJHLIICP6litr9/vXRPMyIyR4B2TEYg2nqQ13v1uq
qS5DHN/tLyiqp2cd76e00CcOF8JebvLnhRQ5CnLmcN8+l3lHaALgFSdg61OkDRoj
Sdb8YeFPgr11OoAsRjQlMJSNYGtSYNR43WXp3qomZSipwUqEeavX11A9fs35NQaB
n53UycocMelTyaGSdlf5FKDTA17VhWq/X5XqEQGKOV7lyZP/P+SLC+LT1CeZOZt8
xQRYu2sYNU0567eI+kTs/D/mnZqTkkBTe5CstD7LwtwTbub6zyOWWLxrzONLlc1R
cL4z1L657WeZUsZcZis9aSfwp5bICOWf90ZdqffOOl6Cwh9ZI+d4tuONJkhDDxbf
kfbShr/azJmUHYs+8sDEYJKKYKRA/Azh3XSUmWkp/RdSdLGhPOD/Hu2LB3RyWZw2
+ADUyt3vXcZwsuNk+mUiVBfHaUh8PooXy33M+Exyew2bkUH3Tlz7Z1LLVPKVTs3N
y4yM+dcUlM+ycxWRiQuJZ9PyPDvSkLeDIRnKbS5k6QhELfpazO5x+YGREw//V5mf
jjsD8ibRRIUkBNUfiK+1tgCiDPOdsXR7LY3McCH6ZbZnqnkWj4rrJ0Gn+LU2FYhI
oybaOu/abGh3g5ouE4zKy8gdN703v4Os+0uNRs25if/alV263uVst1F36S4H+r+y
zWhCk4yrsTjdl0IFw/S6APWwRPY5OPxpEep9rkh9w/und8VAWMLG8V9GZrYGrLce
EXRMd3c30vPrqsJ19gikRQ/4k+/Cfs8+7Bi3A2F6dE3KizAJAEGdfxIQOKr5xqLB
2AgcGAvt3Z49CryYKpSeu7WJRQ04BKDNO7bmzD6QqWMzGASdYInh3I3cyqa469o1
FCbObwpiY2qBVTwkheg29X7MOeGw5LRdSqYBDX4Gq6EiuKw/a4NocEDXKok9StOV
FdJqkYNQajIgET1HeKNHU+0qm/Rszf36E5/D1/6TFw0T40RansImD4CVgruvabY/
v2h0JRw2eCyXe0twKhb4Y3FfIeIc9320ugSIEjW49cxoVSBBKl2uyPBXBTDLbxqQ
muORVVfipDYbw0TtMoPi4oBBNBdEXfstIhTWrzDcmaMbtFocacGPPRUTgcZQ7IkQ
I9s2kAECdo0cz2ugEsP7798w/CK87Ufgt0zRiiI3r3Ihj676T0Xjj/FR5Wqi3hVm
IPyoPS30pw3jEyJWYEPHZgY5JRR+2akANrXBUzb8P4KYBKJO/5l41vjH+JN99lsZ
9FEVSq6VJTW1WG412vQ8l98UcJPbVHo6c18W7z++IQUWqF75ixA9B+N8N7RkJFKl
9jMU8uEwY2+6zTVjl10ar9EJZfyBEz2pVs9zeK9wBG9ZrKNoz5c+yTkUVxH8UADC
QlHCzJWrwYVX3CwbNgD/1zz9XLZdLs0oF4I46D4U4XSpk7NuS6n27w94XYDZtkib
cGGfGcQOHmbAqTImczDHu34B2tzk/RbxFvxfjEKRiwHs00WR/UWRkEfJJzr64GwT
BvOv9f1xxsZIClggynfLo2nbl27/C4TOPXt69ZY3j2fLOcyr6SsbRPwRAJ19TZ0d
nmK1/UrIw585U9nR3CXNdE5ORv4iaTWMS7mp6qEvJ2Fy9Cgbo0xebtPiUGutZxcO
bA1AbtnwAaKCKJveW13rNLpR9rnvFOzQJ8UVwn0hwVUVB3RXOlCbcKC5ReWZlkwI
3wSAtJDYsZM6dM3QBL81kWz7Jhala/Ec+yD0sUUYIo7wAE32a3WE+jCLa+V16R+B
lBvqxsOOjLGBwKBqKtQ2vncoIvbnsCjgLknqSkLbIlZwUJ5A7jrjF4Xj8TtrJPN7
PYIV26qh004LaZSgslYqFq60/4Vrivro1VwBi4av/UaJRCPdfkt+huZ5E1u7JMPE
AvPkQgGs8pLtVoVafwgBQllMdyyA3Zg79IWlH+HulhvyYsoD3Tp991HUIhBgz38b
zhljeywkf4Or0tVq6M10m6evovh2nKIh5T1f6IRNBOYsrylAldXulHmhHCuYQOMG
Rxjngji66g2sZyessHJilSoIGXGAJ9jRc+p5gdC4uV/NgfxxduVnn4W9FrxRHtJG
bJqCjy1RXP9SaC62+gaVG7CftHhD6mLSB7MQhTIG6mB9aNaOC/eQyrKUYTfo+FNk
PUtLJ4nAP/0eJLkHJK0EEmT+mlZT7Zq2Z7JSRmMRZp4x/LJjpIGEFf59XD6PB9YQ
p1TMCVlSKbjEnhbFxIF3OoOjRlAuFQ+uuBDDNho87Vn+ByvcekQMXNv1wvynmGiy
SqrmcqiFlIZFaRINzp3JOvabVbGXUt22Gthe28lCmHdYXTIqLWO0c44dcYD0gh2v
xuRKEac5x4s4QgbyfXyMEdxXsNS5MVP+eGJE5ehQnli8DnxczubCfS1stpnK+mDk
n+E4si7UtCloJHRBU13poYl0lD9IWOdEq/FFJEu0MLnm9GZXittwA5Rj1MdP9Sgo
dVHGx+IMJ16vAe/pA6e2661hFikSLOM6Ipa4O2rfZQ6VdB+2jep7uAAh6LKqUsI8
HaJEF2j980wIf+/ybcqrlppFyr75F9lK0pCsi1gmPraIKnKFugRh0zEkaRl1ZeWl
2lkmRpFS4wZVJLm+I0q4iUFRCIvsJ+5jXQiD+UJuSs5947hexHP0ZPay6lbwVwKk
ZcCw2Dc95SorAU3N9MKE+pTJtWbwGWa/PCr+4ChUZPhX5ft6VWO+tmeVdWdcJJYJ
wMY0MfhUUVWJA7/X5b1dgnjpJY4Od9ciyDPadtt1d3YD2fuzueyfzaoUrDRvnyHJ
TjQr1O5fj/p1bNMFRfsshTl8qk7TdkytY6X62QIT+v6cyGd76FCmY1cXQ2IBBEf9
PrfXIzkAL2t8t8V3r/+CPzKTaLqvB3LIPQRY9PI/S8oeprOjVVnNHpZFcPDuSV5w
+HJUzSDwHFAStcDaYNN80iWWEtphsC/COWIWWJEmMXFZhGducqbtyIPiQ5qrD1A6
9/MHfB/tSjBMFaZGKc+bEYYRwOgAq1+ZaVyvH+7crQq/iYaswb+WKa8XxpCc9nOY
AgNDmxmecA3vOzzcbevwOUaWhR73RQLYBYTcV+sJVLsEYA7q9KHR0OrP9hFMyAkv
HGsrShAbVqSvHv7DeMOlyyUndy2L1ELUgs955BBoM4NuJtv2xj6JApBWCgRzG3F6
wgr/bi84yMk46KiP4WW1UAi5Jnh/wWGHeSnJrdD690/BhAeWuEqBwzgk388gssDU
C9iI1vwTTPicFY7e8j4aDNReWTO6j6TrAA010Sk25F4adXuvZGf7ri2qTDD2ZYB9
GhJlRVFN5zWyz0Aqjm2jLVc4dgfhiRSQQoeS9QPuww2je9eFmeUnpdnaXIFApWyx
36zq5cc/Z1g9GI3ehnJwZy/lLSoTlUoGbSvAuhWd8QawRA+nqXZ6rVZSR5289suD
JFZ4zb7KsFaygPWDp6st6Y5znZkGEiUdDt7hN6Q8qfwHmhfSVfyAzICgnjD4EC3m
/tXpmQr+2oGuwFwc9etsBR9KqaB68pSuYTwk4EA1rnAFIMqJ6FZNMQq/8w/oG1X7
QrjuEfj+8hMI1UZ875GP+3bzzeyXngUBHUWAk6u019+fqWB9LQ2UjlrWHlZbsnzc
IRVfWW19SMdB9GoTjB4HUZSs2Qy0IF+88bgDdFvtAg7P/3TgekIkAl01tyZk3DEF
w8E9vkNoseR7byyKXZqEAqQqjQzlenFKNVKBkjw0c+7RlrhFvjxc1tv0V3vfLtDg
TQ3ZdJzaMS8/9TnsCoEnvOPw3mv3e9xLpxW2c6svIz9Ar8yoHlM1zRdMwXS4wEsB
8Jzex7MAURV0/vPaIJGGYIzuNxXWU8LVEiA0vb7E2awgwQeArLxXd9vimArdFinX
03N2YkETqvG3n+pKq3jMaWzxjcFnRezcYVKvev4nm2wZ/JTCnZHnKnl2GyYX9shI
QY2RBmWF5wBewzxdScIECheisFza26d83iaOlzc1jNyRc4JjZFT/vihyyHbiRS2f
h//mfKJLa4vXzu1cGWl3Dh/wC9VMQA9OjgsJYvgzT9dGyGbM1L4rdcwcgz/N1vVl
lxOEmDCdiKtAxEzEkeGKE3D2ZygfeikQwY2AhKoYh4gvB6MlXuItyXgZJE/raWNW
y5bSzbJwa3cViwn+FwBUZP0JEA8X3v9oC/y533mwBwZEBu3W80ShUY9eOXfnqYzg
8KIWFYLEqdnMC7Tah55i/wvwJ6yJN5sNT2QMv7Mmb7l5UfbfwhIuiQenYKIdGR2D
yyllsXu6MmUg4NKkqz+Z8sRwZvUX3leHZG5KY43OwGpjGTKt+pzvB6vyuJ1uBDtQ
52QvW1uGNMDefDxaQfkwYYzxBM6iLf4t47RctWGokoGJaopI86nh64LIBlbjd7rz
s0fN6um+B/EXotdEB0XcYvh7vJWyE+gR/vf63HdeHwy8sJCubVF5RHDr78fv+hCP
LNBEM+BleQ6Yrq0XPdQ3h/WcXpQyyfa2azZPGDdSmzujQaQjh2NT/hWGhhcGPTHx
Yd3SVBKIwp528+mvYX0s5av791RPrs1RKhEqjQAbU1F09tXPnqkJz5fX9viwoDXf
K5ufp8NCUxEnfuNU70ExURL9ZKb18pNZoiz5bh9mGEXRubK8jmGC24OlREftyqRz
fV2IolcFwy3ctHNumOEME3GWYha2il5aPKW+xmkkuXayaKo+m2UcahGda8Mslb4B
2ExDg4oggKkEZALaWjgHGIRxsy2TrwpTXa4rZHOL3G6LuE11QFxHMlCrahl4EAQG
IUMdlidbrfP0+aCRTg6AwRzioSYrHYhZO1qBqqgvSN6mndoQ1VE03w9E9RCzrwHl
ubttXtqbKO8Fx3icbf00v1lIDw9Cm/YIRHrkGHb0yVUwXyj4e39adbp64YNwXsoD
OwLgz3BY594zR5He/lECPpevNoZZvrhDvgxOdG0VhRaNKPl3xI0V1DpCBVaRr/qy
HLkbh+3kYUkdX8/z3hq2Gxbt95pqgoRv6RzdAQMJniqdH64rrRTpPDFLuVGdd+RV
PhZ8WeHKjigAnrkNZeYrjUlWuzFEhSTE3L+Q5xnuw0DrDZ5se9NYUMoJ4VuQOyhb
0P9PvDB+e5LUlWD95iDVAUHzheZgbaOgdWtp0vExOiXODYSUxkr7hMSUEj5Dybir
XBTg/O7jNzGLf465yRyzW70DMVjGLqKj9e21JJPSdchGaJ2PfE3XrM7Z6ZAYLpXR
Yi9NCzex1zP6/gYnpbM77J6iivqqaFd4FLW2Cn3x/tQFBbfX56odSUxL56ZgKh0o
N4bWa/pwOZKShHCLXrRSUSPezlmGLVZgAcc6x0ZMGzEab6PKvismxE24R33AIN6t
PEaLIm25yLrRP9xq/Qsq6Q8NprCarbIxoqP+7gO5ZvI3DMbx2LlWE0YOIDWcI5E4
0s2/HU4qH+EeIRfeW3TEEQ4tmScrZCreFflpJiYnQKjEJIEADY7fHVR2tIJdadku
HTZTZXaFa04i/bjeWsH3R6fjxEwdnTJGGT5Twredfa3Wao+IQHvhEY7QaqjOrWNT
EjwbavzmOLvz81bFc8OTxDCBvpBzt7uRATuCO5x4sTbEqWBxHdpjwc+jNnwfqS6c
w/MBHMGBcNdtU6iy9q80Fc+C/ITnHGRZzxE9v2YMyXvfMLf2iBxsYvfI7bSPJZVT
duds/ObFPz/lMil4bToeLCNGYlY8NPI60vsFWv/HZCQHdFc+IEZc5r3vB9rPoBTQ
3B10bpgIZzEHIPJDITYX7OaW9JQZ+0wh4whpP8H6uxM8X3njIOKcmwZ3TULjRtbo
kARVc/yFwK+m049rOFIgx13z1o1L42qYU6tBCxAGx+8I7L/Dyzx7e8eGrQxdq/gO
F6JSQbdB9nz/mwyEE0t4wExmKpy8eRSLqM6T5uQluNLDMazGhiO+c8CVo2Lm5/0H
hGSPo/IIptZvbmg9jOGn1LeSgIvXBt56tS5FsE9VkGM4zfzrE4uTH68HKhq5EYWT
CF4ue/064yUMVYyzrfFREjen2PgTHBEYvKIn89yoPmvy9V5JjWHTETz33NKhwcpM
n+Al05EG53iQkmpDLnM6+5eIfGBJCe/Z5ZfNdmRlJDo/mgEyh/2rvrlV5D928GHg
RCX89/15CvoxkG7ZnRhh8lgoneafhIYMN5+bHvDTsXaTwrHqbTSnAQqRk/zkAy3V
bQgiwkjCbYqGusXW9y7RMIgsQMcltHXguruwbApJrdhy18c8qOfDNNCzcTURpVi0
Yj+RE+FTv/BvZfypxq0npccZc/GO+e5z7EkCL9GZpWVuEjGUFso0Z+oHmAFMfM/F
N5GiLtAzfeFj2g2VYpaVm0Hs/Cy+MNtP4K9IrlXe5nxgv0vBrpoB4TkCzpdjtUF0
dqDH5gxLuP0vsokBRnT7Rwv5qTWiUJkIOzWOFexR7bRNYRFHWevYKa5hDJW29HX4
eeG7J4P9nIv4sWVyLUPk8+C7+wZJuNOxRACE21xlIBb/CddyRw1GL3yJP/oJd//s
V55vSYOgptLodfnH7pB+9PpPOjQfDVwTImIXdnXZBs+bCoWPGrORoSrAXufETjsp
C5G0XE1cqqsY7771INwacPIitE8DCzY+qRIALvQnx+cz7kbtM2rHtTCEAgnuZEsf
gQJ7Uimpfav6Qcb2KRN21nshhwBLhvK/WRImkoG4I2LeHY9NXI9kVffbPDYiMW3P
Zfg52rcBNtGUfbAZDuv7lUIHyiyQBra0HPpPBVDd+SQfeXmbG+4+LQog8gCfo3mV
0WYevHkhTf3vxT5VccR+h8dA+o0hHFVT+9YdgZgSTVSBgdvr1edyau/45Z4Ws3gp
avm+azWYRCi9c2xsJnRGjbcYbulOIOA9BKzXAmKGlz7nrpsQqpi4FB1yq0rNr7df
8TJ5p5zrFW8H6o+t6cxwrR2bIKXO+RwVU05wN7rw9nZwcOsBzMBnW/ZDQv6Xhqv8
DWyNnmyBUXZu2OajTaffMVsqhiKW5FA3sjEYrsOyIfTlb05MUquApF9ya0ryuxBE
n5+0TPjyri/AH5paMKXi/bgVrM8fdOz1AYng4hLl+VkovdAAG4MDuANH70UUyArE
yCEmZdftvqnGionHKoHSnQYpUBgYhGxTMK9IHls33yFHLd7BNDKmzPLmfhGbLWtt
n24N7RUH6xq4gTsfxYdmrAkHvxeMQph7vFKJ4v0jW1K9et08J87xxDD5LTNP80xz
qJCscRQpTyyiXMc9tkS2/C5XgX3I33lucXvXcqNghxprIi4CByUGXWndNEAQoKm+
I6STBysbGtqbe5neGatFZi+beQ899wQWW0uLU+CT18k8hxMN9TngKsuN/sder9Yt
WD2SoIBQE0cnyGW4BbO0MQlz3sLAvnfzTQ6ZbD41ITA2RGeYadRg02vR2KTwpG/F
OVkcHHawPzJGNAMto2wzdRanFUX68Z7AMsirPTNC3vmuLyl316D4WGnzS8zXx1f3
GEjfBMqs9roa4BQ6OGOYDACs0m0tg3ycEBxWbAzA/nYdkKk1hiQSLKLL8D/KD6Zl
ozO3pagT6tMlwnGkjcUQrCNeC2MrRgTnpv+4xmYqB+jZbcIT8XgIO7lhwv3mqtcp
7OQypyQ96Rk2Mya3MjYAE1ERQd9sALcsgWr8Sik4iPx7ByvNSvs9q50FxcPma5Hv
QxPYf8dW9725+aISQKXdKJEylSRWlyMiRdeEo/E7wB1ZaUEOHvG9eM1ODIZ2RCTq
xvCcAowMOysFX8OcSwRoJg9D/e4DoyHS52xyWia2UeaKmqQHhO+h+2/pQT9c3nKj
WvWq2VmkfRnxjZij5HY7brN0web4sY2LbrlSg2hIQ5tKJ2lsagsJy4VrBZwVOUOZ
1h+GzWpcSLDDoxKNDn7ttulYMCSL0oH6vHT2ynSO805n1x4iP02avpk+16QkiLHw
h9pJpoQQg7iWYfhpYFtgrH0zdNjYYUjrACBC9NV+HT4FtuYRWbmZXmTRCK0icvuu
pIEnWDS95KJiMFimnm8DvyvlotcUb1/cwWN03yTzxkPtx8YX+5kpll5GgoszUCe7
uPMWMQAcvGrrl5DQcBV9gII+uGtzdXDjBMoZD+ZRXH0BXVAna8VdFCP1WOC4LWPE
lHGDa9Hn9zdiMc0sWnDnnzPhiP1MRIr+4g7A4z1tayLzWGw8dOvzS4u/VPNlUx1J
XVryAV3Ucg4CSHDYzcDWd1UB1MmBc5cKUaQfF5U0K5PfRKX785ZoN6fKpNCi2HUh
WDrpJp3Sw3vt01sPTNkT3QDSDfa/wtVU2wDRn0t9Zd3ZEJAVzFSfMoePic/ru5kO
Y4agQBoqLz3DDSVFNYGV9zfLtU1fYgEtXSr2wbGu6BNXkf7HlxbUjmbbVLuh9j+0
ui6BRSnWRrOjmJR1WhKRnMYKTQ12F+AxHOf2smkaW7TprCzfhTkzMfRtkHSBMaq5
nADCLcZHtnlg6lAy+qyAM+GKTGf+zdBscOuUk4ZynNLX52apwUHraScSeVxZmReH
ukbr39+FHn+3iUVh4v7+VLXuX8sGmOl3DS9br+S3cZAiLMztOPgMaj92yob+cFH2
+kt8NJU6vqBPgVGp+ZJqD79B5L4wWDnyEkw/v7qDTG3Gr4NX0I2XrtPZkyjZtXsP
F2rvhIhrmNAulPIyZMlxBdH+p48VCTS88Ns7RNBkamxaOdrAmw2z5cLeKtB2q98Q
AHwLETovsYEJgZ2Afg8A1FV0jPpBZlaI9vtCWfRA7GH+srM6M1q6mbCdOZjBTgff
IkmB8XJCLlfaY2CjmoVigoDi4+3I70mjD6LtGPTlD65CiaUp2uND/UJCGftntb5G
aDZmrlwo2eHCfQII1eSs00y8h5uhu6k0fVFOzjemDD8L7zwx8UC1zmVSZNM57vSP
nDmQzz2is3qvq5D8Yh7L3VB1EwOXJiA/IIEfild/Ov5CItl/AKlzKbE8UxU2hwFK
gun5rB6koYW0LPN2hS+Kn/9/m3PKfMhLq9CGcGy++R5o5UVdnIbp12pXfNZ4SAQA
JmNErVanOUsZwEmDTO+wLLir9Nkxt4I0cYBBEsTY9E/cm5GAjh3Bxsj3jobXs7lJ
0LSz2JUHtUbNhv7Pf/c7Q7WViseDD0mKvpcrSCzuKSbCdJMEslA36/vcRiTN3Lzt
kD3ZOIM3mZKkByIz8kNK8G6GXaKiK6QQbthEXCQR01y7Lrdht3y3FJJmCcXoaOzy
WEjoZV2/uE5RLLjfjdKzZo8XC7jcEb+88bsW3ZXY2uSCC8Ub3sOr/osdJ85TXB7T
CIehV78q7IXbdc7A+O+p0wQKF/xpLhQKR4enTMe7rUgrQ4aVF3eVe7cwpdCwNxv4
HXkBSE2VbZ9q8xNEMM7jnOFrw+XO25czQ63FRdMhatxfp5DKc4IwRi20vS0ZqyQd
epQwST47BmA3FZ0Gm9pyOBkCz0OGMoSNl6SYFO/YG2E+VhH8F+9WXjnDrmShEZoW
cYyb6Ivw4dOGZeOMXaxvwwz/tN8N4DTLQ4q2gbhl180R0vmXq/E5RPQqUZ4vIJDK
rLtxEvfPUbvrVf/bPn6jTj14LI/WaG9HUGRqFrn1O/sGGW7ccTIs8E473WcUBCaR
j/d0JWBBiUsfu6RHyapidvtWZ3Ryw7sulUrvIub/O/wD0daIzzs8CGujQH1dBIXf
nZH4osjGygAZAH/KPl8drubCCXisSHl+hM17SSQZ0o9aZ5NtFP5Vl92Ff0WXJuI0
odOr4+WTGW0yoT/rSrsl/wCpNBwNN1Y6tiez4IM7mgFWCdkpfBZH/IYCB4cKDYGp
JYkIxxTGRfK+DQOYTP5x1u0f+Wkn13fiwwmDEcNSbdg4ra40rdiCZKZixaLesVJf
zZ46Qf5vCbfVaOHFymgZy3Q8XzHffNlZ8d18RD5f+CmRMVZVTnJ9VGDZG0PINpRw
OCeUWjAS8ll+ECWT28Y5b4I0KqYeyAdwSGaQhBtiTFNpdBc1zq3B2IkoUmEAV7Vj
ipJBMBEynqg04GflM7crf/mb3ujcupGJQOzDjhTogEPFt5UloAOwcKnr6mBu7zNk
a3gTCOzAtV029mrWSCZAU9MPfS07zOuFYMM6i4HzCMyvTpKrhxDiLVEN1NDm+Fsh
xXtSz4AkZzsShZyfFc4x5QvP3SkrdwHfIl7VNmAhcWl7ojL5y+DnFY+T5oHkSb0q
SYqxdY1X0RrbJIBeX6IuTqX/DVfrXqS7TRuXRKm+WXLS1AEjdmI+PvxGORtgotus
gJmxOngfd6WDsay3lWOGerYKUYZNx+lvWj2Exer+/I5dWl3XQ305MCUEyamDo/hw
SDaboGv6nghSuMAeUT70ZFM7jY2HadGbM90Clz4C4AVA94u3fNgdhAQmRwmJGpBn
Nreksf9Q8hAq5z2rscnWOyI91lwR59hIq90TFcy8RFc0Xi+uM9mY857Xz5PKglx1
dPNvFnMUUZBj90qu8HXNIHtFr0X4JjF0ScY+4VrLmv+WweZ6jUvfYFA+nJe0/pIp
ppyJFe0bLPh24H0b8tbyzqw34qH09v5I18NDiURrotL+t6JEVg4lpfDx4Jj8YEEC
VeiFXWlpZ+231iQTgrP6z26V8ZotRtz4YgIPt83rLrwZ/a4TzTBxxKZUHsN/w72p
y++IIUqCiOrUSSRSHykzER9szrlRroI4P+SXhrg6a0/6fFFLQQ5UCIK8/pztXCzK
ZWuBSyigu04AIdpgRR57jAIHqCXIgiWKOvwtTn+HCOX6a2rbxXUFKmBY1LOcMr7w
Vu6pOkRNTQjBcZ/PEEPMV3GUGDVlKU5RzKVlR0vssDaloSMIuT3dZEKTNlsvzpjI
nYFJbWzIDyo0EHn2YUZYLdSMJxtnQgIhhUnLhDbWVrZC+GctwKHg8R1pDR4b5X1p
s677lLp1HTmkij/oVw84vc/KTqSkxU7oK8J4U7eMRMj6lUH1dSzSGO/vs2dTlsdl
wRnGpdifAFnRcuHiE/m/mcEkZ9p0PHoZ7cWwEjMKHAXQRwNhqZHL8B8DB032+HFQ
oIuL4YorpU+5ag0ldJNQq7IStdxKwH+Gf89VbcC0phzNw1eX8iaOvXYFtwpUx2Xz
74cgKjOUU07D+S5Q5yIl8ahGKIJ26nvH8SNoLJyrX5aQUfxBZLzXuDdxV+aSJQmb
j/fUfUwqaV4uc//Aj3GB9sLFhXiWAogQRlg120cnvGxcs+K9ORtAzS8FQAjmgXf6
cT42KiYo4GefFTJg8/UqDFhWl7rLIGHDvh4EZx8TISuwnoPzkF7htGmYVybh0LUK
QVBUtzmU2a7Rwn1Kpddco+Abw+jYRKvSKlfXT5xOsX7XeYLxUWwQRglkp3AeG7PK
TNxtLLd5D2PIEQZ3Sb5MiKerS0HSLKSkDqwSUfAtsDmS7G9kgGeyGoVysDCngAW4
3QYLUf020MD8/tl6ip1ZjhrK//dvm9csCyhUzAzJy5sl3cIhn92smREs1HBrYhKC
1239bX4xuA3nJciXzJV1j5z4IMLFdRYcJkhRzxhFRXfmWbyN7AvM3omzePl/vUNC
LxvXjyuOmzMzS/i53Ej+zLLaTpFfQcYeyrOdPmPwjFqmFrk6YXNg95EzsisfGEYM
F6R74/GQz8DbNOWicqH1OTAdqkDxzBdTbkNSamLqNihs6vyBonuCiFIloeCw9pCr
tG01+WyZxthNBWNEqZEY3cbS022Fq7kDQNmt+EsLyHn7EJkSjCGSr9VQxYv9t9vy
7AiTNnaZWUgWI5Fim4Y9sRR8bdm6s8obxRH3qX28ul4ENLjNdgQ3LWcYMY8A7lDc
bDLLaCXDKZ5Jpx4WSRba319tgmMjkY+qQS2e6xwRvIRdIzyjeBMOfDnZKZFY8MsD
Ay3bBeD6Jgixmw1PfhydzzcFtXqKaCWH7u1V7duW/KTsY+prPj6q2uJdPhkzeWOP
NqZOgmsq8tcJx9CGL36Q8zVDd/Lp8x9MEDY4YpmqOiE+661FH/dMK2fjUP532YTq
aWdvzU6eHbeYUpaS0go0lrtmhESotaQUvQxXH4B5lsMqb3NdcXCTH1Qu/h9Hode2
22VKVmsL7g3zv6J6tP1cxDuAz7ggc5rc5Oxrsk+k+J4NQ1lszfoYMSTgBRUfZrtY
La9VkzGu/JCs9YjoWd70lNUrEFp/UTGVIFIqRnhu9mZT5a2XVrzbVP41RsY8Dn7N
CIZSb6V3lxJgNdyoj1YcT/26eGYH9ArWXzMKmPD0Jxd07mCz+A+3mGh6zZlxKTo8
YQ1rlB3sQD7xJJ+ZNyS6eZNGM7f4ZmHMMek0XUKd1/H8wS4rvVA/lWAo4nIM9y2K
Wn3og17ydtgpkfbZl6P/09FMVXOIhEtiIlrIbB7si23oWelFCa0CdYQ3PEFJbA9e
PDm/SwhvX7CoEwhs0rLHDMTE6x1fNpoMljlJ6i7RKkbuGq3Q7+zsuK/4eFoeAbHT
kx1LNRPKjVa4tvC3jvUK2C+SpQ+pjK7YzaoRavhJ3CTzz6CLLCgEDfhgcAqx0qif
krIfkOiSOMH/INH63xFYcE2aKsrqkV+9Comb60YpHqX4MZV3/4Hhya5pbDlGbXy7
rw9yAdnQORRtoPvWPWm+pMxMjfQQ67kIrzW636tArAMLll2z33RJlSPlt9t+ytml
yny7w5rZpOKY8tJbJMd/cFoQrCuQa/pJJCeZ2zrIan2DCDWRca13vZsNIOzeKMvc
3vEHjhHp542y6KSVTL3ZkIV4beh2lIglKh2omf4lJBfFUFNV+/T4VotUElLTPzhC
z7ZPxPzidGLu2h/+Kfn4ETvSRKqJULY0/DM/9AGVwnDEUDkkXArSAB+hTkqGqB9O
F54aVv98OSBIhBBVyuLhZCYUtWn/yj7T82a1/Bp71uVA+u5oa3fyeds+xloFcJMG
`protect END_PROTECTED
