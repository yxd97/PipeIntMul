`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
edin3jjuXk7PA4aq7hfjRRrw9kOC8Z2S8gFTVtzBX9zxL1bRVZ8diHGYDYqwTsZg
gDP8g9qDUpq+Qd09kjp/70BlMyWjqolXW/tcwg21gfomvT1R8Uj3jWHrM7jQSTOW
7tf+gPMGtChz3faQ7uHFfzQSM8mJ/n/CrxiSDi8d2Hyil2joTxBgDlp5oSQmQwK8
2kxRitMEQ5AHJHIFy25Zn6+f2MEY0KceWElAdIVBFaoCKkl8p1Lmegp4UI29PO8g
pnxcHMeCzUitlqjV0zor0w==
`protect END_PROTECTED
