`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LME5m6+K7DpPNh2NpYlfP8FwbnWCr1wm/5dDESXCSIUDrzpI8EWpLdf94nzPNtG7
/lU+nS4SgRlQVDSZixyON0XW4NDwDOdiSQcwStt+A1vcMKHsCFH46pjJmQuzIbmb
RXxfcOR5XI193alTuH430+RyR858V8fRCRmH+StxXI1KZl67Oi0tYo8yV3iMxMat
Qh78LHGL2UvPB5VrKDjVGfp6eB/JgLA5FpXZekwaMi+vBQ/Sf2CjJMRB8AJnDNTc
lCqG93fL+tWyzt14Bhv9FB499oE5NoG9PKKjXRhUdDHJz/LTcgWwobuf1hbwfn28
2XsIvbkzbKRRuJaat/T16g==
`protect END_PROTECTED
