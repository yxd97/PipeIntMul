`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZkquswG8hrAfR+/yz15JFekQkTskycNLTRG9Pf+SzliXsM0eWKnU0OzlaK/4Uq5X
SuNCPYSaBy0I8lnOTfqJ48lPJhRF3zdN1p4TVtYNy118SqT2fys6SaHBVSBv6ten
bGG7/UhbcnKac6elvdEpPE/WTdmLGHE7rq5Gt5E6wMwVtJT0MX8/AnwuVMWwRYV9
pi5gWvLhomQM2w5t/5ysi7Py/NSkENrmTxORR8VwPuapThh0oeG3/WFCYQkFC5V/
dwNiBP1JLkMlmXDF4+/lGDHNgm3gAjNynoqMIxML84+3DCCuZlG5WG0j0wdq2Jfp
mcNDWTwggMLfKzDaCP0ptJue0X7y8SzPLwgXlSYh4AkbtTrpyRbL5Ssw/Je0rCAZ
+1m+8BiWzBRYn3FbqKPZ4Z7KQsPbd57Ea+bt8/Va2VQ=
`protect END_PROTECTED
