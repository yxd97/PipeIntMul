`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bRk+gpAM766HWow1JF/PyDPHoCiTvS4c091HnT9KQiFYVYNcibY8zjwxR65AndMy
+mgAGef0K8eiAUNMN41H6MqBXrhzq48uuyViJThZ3QQJyjK05eoirqlthnJLFBHz
WwOX7Qga4y8FVQNcIRehHd5AoEJ0ImNtvh9e+7SlPPFg+hMzCTjrYvCaDFZXgXz4
M6vyA8c4lS3ucHC0AhoHprI50NtALjOsM91knsl02J1vMiQwAoxZYkXSr5OmiFcv
UkmhC1TyeYl9W+sFjknIhd0r2mpNn5jFw1xYwFbziY9o2L1iho/7Owhu+Jm9hiF2
clKxkv9NjdN6FrEywumVyQQh1VkVTc2M81RamNuvsKZO79/EjuVN7xv9HNDflQtb
FZ5f1G6YwRaj3lSnkNExbH8fddAZy0k9/JRk9/KXfhbxMzx37F65X0CsRB11iTvo
HDezxjL8FIU9wAcwHsweWA==
`protect END_PROTECTED
