`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDqSESD9uwhN37Ob1Igax1L2Ba7gsuxQFdsEJp6Of92gcqMddiu+agB41pSfM7ee
GkzwdOPeUCtQ/4A9oy4G0mMI5VZaRmjRGE0X2rhKYP7vOT7pL+UjV2P05ybz79l4
Bcoy0kWdm/qxJ6xnqKFsp+1ZIhrLZeUvATSVwZCh3Wv7yLsa6lDdbSsBvAkVm7lY
evOKr1EkJRaAaq4HmtmAztjLZRvbfgXwn1drM8MDpruaw1eQva5PBMXMC5bA6ODS
TuF0UqLqN6Fwb25EDar6OKfHP+lnq/K0s6/Q38/pTfkU3YTQ040e9aauZwmrN5N2
HQW6i11gJHJpwfv29KcEfnSka0NhGWOzOe/SgbJRfME9FKyBexD9V04NQh7KbTz9
Q2Ju+AZolkFgII/xa73ZPj5LjS7l15yBPWFzJNy+gEBZJmltIP35hGf5275OQEyp
9aMXd439Crg5WQvXvhejWiFrtl8aOKuPoo9fCo9rSJ8q+blKonkpyuVA8vsUl5ki
6E7CF1LNrjSIIZS+x0UZx1O7avf3mHNBqzYVTW4VciVt/yF9Q7edQovQZxlcTtqG
Ibrq5lT6wCB5G7OZ9CoURYW+3ROQxCjc3Ut4jcGCLrxeVvFHaMETPc6q1lblDTal
mautaqKqvZ6PLlysXvS36/U7BPvaG1YfKioQtZRQ4O8=
`protect END_PROTECTED
