`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9skrQOEGPzT7FdTaWjbxa9Qc0ps6OgSjIRaw1QitViCKcBpJZG2X83sB+xAPnXpn
SFUiP1+TmWO2BzoK/6OA5ne4YKsl49jW+Fh49FHtUSXNlQu3plVvoLIhR64/r6er
CNl2wPpHi8NLkWy5kYDq5kGBcyBu3cVlG84dvOid//VNZO1USG7hhVllJV7f78tB
NhonnUPdYYRAtRRsjCWKloYIlF+OytsPuC595PCsiUt6yyqjIE+Wiz08//zvtfgL
+iRJf1LDznSczTt8WXYfW+wxx6PAOkPG51nKQnhu2VzP9BAp6GDivsTD41cKpV2H
IdbQhXlp10+QpKcr157cdp7w6fo9DTjfXMrvgZx/D2I+BVcPYNNkpepkMMNfUbr6
Y45tWj+Ww/PfYEKsqgSPp9aUkD4B4MfyXdYGOKoLCjTSr4B+osoY9+ELHmR3noCw
cbCzL6ob1p3trvKjwSaPGA==
`protect END_PROTECTED
