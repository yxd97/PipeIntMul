`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fM6nWw74TekthrdaZs/U8ET5hxdo/7EACWjRnLR2FKsEQ/qXy8lH3Q4Pu+cLgb8d
7AJyJ8McNzTgVog6oCpx8Jj86G3X+p9cXUhNHjZdwj/4jM2vktokATeiF/1jh4SP
olwbHzNHncyuZ5138yxLgSG/09KDEPbSvuq1EXCJLGNpwzBAKe2K03lQjcQ1kUL6
aDjtgCLuhwc+ScjGCRYHYyJwHlcDKJf5ydBCQS58lX6s0Bih70iSeHiAR8aVfQSX
2OxFsHr0tkA1vijq0KQcZxtpp+PegZde5u8rVSsj9amOq+QgIbP1d+2Y3h14pLxv
qgl6DF6JsW9+D8Okj1EHKwUkXX9XwzvQLZ60IvO+DSc=
`protect END_PROTECTED
