`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5LtmBiFX8RWpHfDPMkP+WHHVLbh1/BDGPZJPjcG1tqvHNw5uGDffuZRHVu/IMzKy
dbsK2xaYegojnn6cuGNwC0WxVzOXa+VnOf/6hlEHQaRK/5lF/dmgNNT3T07UAIwv
pKQNOfP1s6KTwDETeSELU19Z8zxx2Uk351t5goz0NN2DlxHl+dVMtooe/X16dpfz
ugrlcwUO2qOAtty6FMvS/FjO1UAo8xWvHOuf3cPOciE2xy3nWbLPRtJVFZ+m9w5Z
BHL1rvvQn03cwsOcqRqBew0Nugc3kuTkktYNzr3ITyardjwQLzPMPrvNaRWPZxsp
uscEk/8Uxxwg+4girlHqI9t72LgSNnIHu9gOlyYqiLK/2w5Mnv1T+ZrB1TcUV772
+4DaCCHjnGoZllVRfr1oo2D+oI0RLEPtsIJ5Rk+oFCUKOiGEi89Z03s0Z38z1S2p
HJHdJp1QXmKufPR965cJO2v1Ll+JMeY0bdizRisLD89LTWcsolqWot/xVc3boy13
JJZhd/1IZsUTIZhBtu9l365PBPk+bSrhOix+kXunMMtRP0qab90kCbvQ4o9l3liR
ALu58b/I7V1QmhZunRyKc7Hdvzf9fATsZj4/IshKEgsEJRIX2Yk5mIMTjIRQj0nU
QSM0wYTixwavoz8X74e3SmZ8T/sZNxPbralWYGAWHl5HSdizt2t2pCDmi52zIRZV
giXkDngMYi2AGXNtnav8t+ia7DyNP143t1uum0aEURTGBc3N9vZgKs42jCL315SA
zZXYC+mdp+UOvkaGlgV/4+vfR0ADYpIYhzIZQ7yBc5LidO1Yc77pVRy/87KJqPJy
yJFzxAm5G3Fw10e9/fQ0l00eq2Dv6uVLEvURBZfjPf0gkr+e/dYSasdYL7Zf5G0m
/usbtV8lfbUwW/EFShmVgmb8VLPG3TVsn6fP3VgNccYyJiWculGFmbSC7h4Y5HRq
kIJ/FRBog7GVJnRIziH9SkZTd13ivHdtkWwlCk89sEv/KHG/XNvgvHheu2O16bwa
Sa9YM3hYq8SMmhL7KjPfoiz5Ycr52DEZakVSwlXpTcUu3ZV++rKEfuHFSQD3b1mg
Pv76MtgPNIwpEy1JN1AzTwz1aayjncLRrbkyeB6LpHShzQOkLhTw03xeIqVaJmBo
DakPfEe1sSqGXva6aFDcZOD6KtYULhPrnyQC5fiHMeZbgphV7TYe/xDNvLz5SIVw
wK42KLbs9EPDB0b0TWqrr/lrUBfx6I4a+ZgDETj7AElBcHuZPjRkqYnAuKycjWUd
B7VA3bO1lLAXsk4TkwBunfbWe0dj8MjDN7A5ivKhD+7mJdN2aNaFpmZDwUxmKIMT
N2XkaSJQbN3hf2cfcsCJtwLneVXLQNQW8Q2FxujLKtIybkpMqvvJmnroHw/jm1uH
vEPiTdQzrD7t9haGCFEQEB7H0auDTlwxfXtDP76nbPDBt2cVjQJOzFb6FG0+TvB6
Luu5cms9Z/donZcSYhCR8BkDz6frydzW+2SEFtbnbpL9a2I1Uun9umLw26rAntLI
hSJNupGE2pX2Eo6H2lz+KARGr0vZMk2Ld00zuaEvS3ht7PWrZ1C40xa6AT8TqwDi
hyqYo1mRD6sqbDlAkiz3NTKKtPT2X00c1WV/hTQkLwvNCNwY97O91sHyZd0yHL6F
9VO2KAp0KbqmMEi4vrhzcTc6JMF1eOeT4p8P9Dh91mP5wP1AtW9sjAwlvGLzPUI9
NHYlZ7WvOaTNncaHiroYV/oY6MQd3aRXga1CqPJIYWmv4XbCt8P6SSp0GLvIqQvF
LWaYcWepA1aqfNZvf/s1nKvfnYi406ML8PW0MNtYlWJtmOVXMFR4R/jXaLpvKUBf
kvYo8arMj+V0TM5td1SpMRu9gOemzY6jkcTDWhXtuPVeQvjsxqYSdRpJgSFOFPJT
Kubt2eDjuZdRu9uX47xIkhYfr5Bey3Wc2a/D79yVY4Bo8ko0XYEuB4LngVXzqQdb
gE6SZZbz1jU+MT/T+/95jHyB31XWuSsNsVYgSlJ4Ea8U3j/CLjFDWRxj+Ou/QMVL
XWhTJtLGjLSWKeYz7QM27g==
`protect END_PROTECTED
