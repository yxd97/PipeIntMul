`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5UM9KV7YNic9x9tJy7lKUVKPRsh9wi22dhbCu24d9Mk/zQcQVY754fmeG8Hrnc4
VNaWNBfffzpfASv6CmaTEFZK0XxjNtQLwi6blAvrK9n9t6JjfEDBOC5ccoxr5XWx
mvJ+7uaRugS/DuSLD+EkP4gMZRkbbcayR4B0WTM+MqaX+DdS7NegSydU/CoKKpi3
yxsJXGkCVHX0FVv1VkU6Semfu70OiWwz+gVUZMHNk8fYH+JgNPS9es3RazjGcYxH
NTuabqcO9bB3e0n/QxXk1axSeUW5U/SAfoBLVDYDH9tkEpvUuUIh/5fWWxO/tdZP
WnQFE3dFGG9cpR6S0x+M+iAVbi63i65A3Xdc7yI006qzVPD3OgjQRCc+cuRwK2AE
oNYktDZJ7LJmaijdmZ3okeGeBdXe3cJ4V2AgBuJfZiqB35UTKypJw86j68g99ydN
Wu+7qLwXZyy5Mqq4ZVCVNUBAC/PcCpP6Ov6vBPGGSzA=
`protect END_PROTECTED
