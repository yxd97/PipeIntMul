`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CuPx3f4y2td04ZrEY+VAjqHI6WIMPl46FI3WSKq9hiXZlTMEYLrxXLljNr/abTnK
mpHvlCIvTs1X/qfEr4VuQvcpgLzV6hrHCrEDS2AIdH5+8hK1WP5eZ4tb/osuHeMS
W/Ca/Syc+Vyt9MR8IaLHK6IDOMbMYmr84N+MK54omi3/l0RVKLRNlmXkRoDZ4umm
bXPmxX6gmKAC9LX8I1nxATheBr4crLd4KxP4KTlQZ8OwLBzi7tvgUeU+ezxkl5F8
gbhZ8MYa7Z5WYv4p0j2dTY+wTNZWvxg/jZu5FVxpWEp6YyaA3a3DRFcL7A0veyjP
n2ItWu96z6ouHnxsediDDqHmIPRMh5UPXoqRzbkcBfRYpwx++jnPorKfXl0Eabh5
C1QYweh2seiwKurBZqT5JjyM/z7DmcayW0vxnOPiLYYpRarcHpP2osBg2DDN7nWC
MgB8ZsQjQ2b0nlB9BCDqAbs+3fJVP4AlzuEiYgHcc38=
`protect END_PROTECTED
