`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KELkQlsiDkUngBXP6L10sI7IlJr6lxYSRkljyWqNGz+8oOgWnhmheogrrcd8FAaM
f2Ln/4IjHYhMkBarZrgMbXGiiATv4UTrp7qgeKo55hiK4Y6pQoT6nlXDH1eYR2HO
jFb54G/KkaIU8qp1hSl4lkkr7MrJPpKNhzsxj8RjP9Ph+vZoOaZjLToHtJhyk7Fi
PSk3z5DkyBbbpi1YwygtnYF7l+IAFiJvr2IKxwkLDrUKV3mLI6bVCmj8qmUvh51i
tCOkZhsX3zJ20dZCL6wdKKFrL80ysLzH6b9eQtA2d2w2aFsZqQyezCJekhkENNKq
SwLyokGQw9Rqx0nnridwZJ1UPdWGyLdHCiWH3b7mfZaVsFE3VbsQgR4v8aKvUFlu
PdXNyCEbKoN86vENbfQjMWktCvpmT2VpLKro6T1DDTaPpTTxNUEfLHBVWZ2e0vIF
uxSkbPGA4O3lA7ZOtf6ns7CbMWHjD0rUwW/FvlHc8Ku2wjiL+GyzOJ0SLXbuHGkd
/c3vDNhyV773ZpV4KlDVv7ZWDHGo5KLOa4IGOpUxJznRjlOWL9YLgl1/6MNUmEue
UBwzeGzAw5gtVAugXFq9TlXkvbtNA/7t14WkIXwb9MKyZREZyfFMs0byfhl5DNTH
sG5pWLkl3SoDrhQymOoD75ZZXpnXxumllTbB9vrPQKxJmGd7aAhD1Fw/FZONfRyf
/rJHX3s0A3cFIq2fk98roTWJp+fpynA959Re//sDH1UzlxlYKqXW0ZSxkG1V3Ryn
VcSWqkoN6mWxCn0SlzF2RLA/EDRRQrS0T/UQHizsFcvYXWnphppj0fI0mhEQq/At
njsquatvPExO3ceigxHb5DmQTWlOM/ZnjGxby8Lvb49hL1gGXt54+XMu3J76HELm
EKuSHvI84Jeb5GuXJampxF1b/zIRbqhXBCCCSUfqP96RwXbOBE/sAfvb5UM+ekGR
2lhZ/R1E2on435pWSw5TMA==
`protect END_PROTECTED
