`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XkUXJ03jmf5cL6L8H765bb9L8XOat9etVazTgJJmV8ek/qOUcn33hiq9DAXtbW9P
49jVoj1pJP0VLlTv4QZ3O3zscCchxJwd/Luv6kTekJ9puCCrvyn5MPhpdV0cErAM
VlQ0yCYhjxcCqW3B/g79pNA7OirvxAYPHtQvqu/Ijv3k+RpX9UOrSaJeGybXBjtk
nNFkmuWTEoHJ257P51NMn5wXcCfKAKaHggacMMllvH4Nq6Z3QEfOKEHidReTjRzt
OCBsW6Xb2th/D/hHMyMdXnG/gEe8PqGdDT0uDS6rn4Gh/yzm5SNnIFrx8k38ybPC
AnMNz9uEtgnGeTBy7KYi2r4a7ZB3pJ+81UuipmMYKO1DkarsSvEqZNUYN/oV4B2r
MP5y3ncsgYR9d3gLRCYF94HUzK1aqT3HXhKM2ao+ees=
`protect END_PROTECTED
