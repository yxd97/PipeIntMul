`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ysj0NFQ9wRKpZyEhx63cijl9qcicT86oHL/FijDQhGU0ERUKI2mDmjgQ+DJlGLxv
L0K2KBSe2upyqBC8FykT5pgRKw+tBSQaSS+OfmNJmzr/vQdnNQ/kqHcH801IEfPn
ADxplJAxlx1WYmB1POKXReXQHyfH+ecGDlsdqkKWgVniD3xWjNYPUci7doYPkQik
C/lx96Z+S8so8D4tRAAW8w/Pl6ACRch7aoHM7TagMwfSFhSefj3Lw1b7NIfV4YZR
lA5hdVrqws3ugLjLO+dEvOO6Yw3SdIMi3XZg4IgqwrOa/w/OIMk4hfG2DleO+Yww
iW+btVVvYEr3URk+uTkX2yhLVPfC9WBk8I5nVEujFGablHO0D+CnVbNuz4KcY//+
mMrm/OZ1E1xlJp6R8z3kt/hqeZTWGxl3uJt8xRU7BLwAlVe28DJy8Rc3ShV3OPip
gHpG8BM6wqieE41+bNmcLoNlQTK2YjROdAyAtyW6rh23LbujnWlAJrhv9ypky/GF
F1K/vn7xIzIfzR1HE0YlEwYu6zOyaw7msTCcsyS9ZoU=
`protect END_PROTECTED
