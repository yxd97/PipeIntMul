`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jG3y5rLjafVCTBURauIPc1o5MrmRABn73fCZb/bEuZTSLtyEHePdANXiHKiYbj/j
1+bc+T2f7AGG/bV9/XkYPIuXUM+iaXy4RWtZ5uK4i1QO3MD9i3xoE70MscMl8ivI
4qjUYwHEWGF/Mc7c6H62LrScsCHDUdkDcEKLTGVDdfljhfsgdrcM4Hrln6ZT7Qct
Crm9MTmD+O1sJIPajoo5jSjJCme5a3e548FFGcBukQfDZ+4ZASU50xw5vARYumw4
KTX86pRi0lcQyBW42p92CIyGs6NWq1Qc5YavmrusHUqYwRD0ZLPeFBiZaJKcAmou
42nfYJ0oeufS4zDVRSnz1rVrTWCHhahB1pdoslNuq6WY5M5MtDEUASvZoEomToZW
rEfg34/l2/ofz9UbKvXSoLcvi1WUEJGMgzrtmlDciL4=
`protect END_PROTECTED
