`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0tZGEedjvHIKVx8uc9c0wlu5/WGOvh4nTbF5cyI8W5izTIl9i+kmUJB50U31iniT
2UVE2yqUdW5WFHaNeSRhNBPg0+srSgfmifWWQMjWk2fAd7OCqfZif8RXAf/qM9HA
sKDAy0K2sTa+pQwI3jdiCVnkPId7zgIHW1+Odddkq5OJZF69xVvsaShhnw8Tup+J
cF/96jaqf3w2DJH66LKgZTHwxESgpJUgP0Q41z2ZDnA1aafF9H7csC0JDqgLmYUm
0yl0Rokke+J00PQ8hfuKgQZD3czqRTTlZbDm5KIYnxyPR8CNUr9MGbTlDaBOLyap
Bi5hGBRgJrr1dXXNK9Nbigpve016KADSvzwJhCMn4Z2KRl5zPPgbJ3t2ANnffunz
Gwm+6ifKYieJffTcBRMlluwxhPlor+ufir+IiQmOAKbgVxd+CVuicaWc2qnrkMRb
uXfDjQk3DKg+pXYHDU36YGZPvE/V4WW1pb0RsLnYEpOuSdzxpHetC82GYMiCtd0a
`protect END_PROTECTED
