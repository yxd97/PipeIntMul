`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJGOBlrYWhJ7pTJX7s6JQtUSU0/mzze8Gtetyw6rIL4r71qe48TwnCNPW1xxklMS
xt+7p5j01U6ZWylrJ2nEZ7JHDsJdo7ftUSt8XlTwT+gFUc5HzAnI050yprnmTeOK
REbnS+r5HQ1O02YUg878OrL0mcCFXAS/lxu5SkljZ1EhpfdqLLTGcmDsNtEFM3TK
gdDTc0hxqRzL++5lYAIG9IngPA1emLMZV1c1WtB44CAsLQ5edlGBG9B79YMRlfXn
FwBjSIJsuIqdWj6s3Ca2cc/mWyv2TrNLaE0yvM6C8AYI0rlZ8EVhd9ZgAT9by938
rwRrH4yb8zEFg53k5S1Dwav7aFeTL+iR8zpZVWmgXVz2BvMXZIUyEXjZNaU13Fxx
xicTg8SJb4Cdg6qFSNnGJMZgS1bpoj3uxZoHd/yRQ1ghEj17jK9k6CwsICLPpDw3
y/FQzvZcF/RRJcPTIn0Tdiu048VyCgko1AuJ2zppf5T06pDLCCu+5LGU6NxURmne
mtqDRNOSMuXC/SjQDsp84KxUJsvALgkT3X0kFXGNOfY1nhGOs1puJ7n7dVm0WBQY
VH8sAyl1wZuPPx2VcIW+QJFuTS/5Df5jCz5ljZziWBfKV1O6Yugi8sEQ4DTbto8x
cRfZ1BqGMDKDzaR1K9vAli2uZdk6TL6gqfq817pDIhCdSGq9KlfOoY1rfh1Aqn1G
RSbrscXROcN1vANZIfXr+RNYosgIkwEsJyusgfg1WVUJFtTaOTHxTlUekhvSSZ8W
qoFYpkdPYnMqZQblnVobqqr8Vu3Hjt863KaVx+Pa3dcDUcRsG/J8fDTtTv4Yreik
sE3VKG6Q3Avr4b5lgiTctI7kN3SCdl/XG/yaPVZlSV3QCD7A4kXTtZEG1uDxzPNV
xtZoHClYy81lhzplK4bx5U2UV5bQP5XGqt2XYEhmKt1zEqD/M7P2WSg78mAj2/pF
CK1M1NVPJe5NvQp32PY0IiR444FDjumdyF0AnwANamt6x/xekxpaqSx8xkoghMDs
4vYUEhhoH3r9ZNpwDxroOhauBjDcvr75ibZ5dtdOfLyQpyB5wr41vZzJZg8OxyUR
4D4iUgJXPw6ZODfycC2yM0FoCnIxy7Fj3bNepMpyB2gAokps/+k3FAyjJRcvVTqq
FFcrrvfSEBKTU0s4MdXTwPA2LyHMeH2+XgP3iITOz1U/Q/doSFaGMe0JdEkmNU7b
1Cz6NuZVEmXgZz7x/5WGzFcSp6vujzaQjPvlyLVbSSy6XHrx9cnboGMzQkP9A+eN
0OiFak6hV7beuV8lA3BHEdyrjCUs9O/8BWpHMr2gr5UtoDCym4gKmgshd/cTG0R5
jEKU3FVA9G1pL80LVXi+r+0LDPhoZ38jOC9Ux5sTDOcUh2J15Dv2ZsIffVoo3p71
MUYb+lAiM50iolXUYbxnzz8EU3ruju36Nrm0cgEXtwWKQKLqiGzm4u/LoZ0501Mw
58/pt3CZ3PUiCsx6IUdMVL3kfuJHBlT26opK+n+YBEPAVW2Z+P5hhKu8rGVlTj1A
yNJf0K2ddLb2dfEFgQYS6ddnxWpdVCG/D/9CcOCjg+r9oeio0QzanIEzPhwMCzWY
9V6Jn+yeSg5XSTFxygOFaGmuwBQ+YQfCNAaRj2B3Z+W2MUaEeSa63MbIa/71FZ6A
bj3ozJfiwpdTOOzIsyQnMjjF9fj6pcAaaEwwVrTZ+j5DxiHxrTE7IL/eou035wDT
jOXSOK4RpWQb8l2tim4meLVeO2As/rorv7lgjw0jENUK1aICG6R4Qf5Vo2Mic7T9
9qrCE0YzcaoHvjpdchPPR7PyGzI/6hPWTUWTQ5bCV8iFKlPAFlScfzBS42p4vF5W
Wdg3s8tArd/nKb2cLeP5SggdYBnvaBROSOP4O9a6lc5SOHONMrq5FvDctz65C9va
6+Z3MMgE48iXUvYgfGf0ghPs3R69Emn7bB42okDQSpmQRcIOsAZr0rxMu08eUpHs
cPZpVmpTR5z8DMtCZqvMuF/V+mQ6/y9C9a2WLDcUjpCbWg3WR88LnfKXcGnj/4PI
bJ204WgHK/mPbPR7JF8GD9JjQZ0WoocpaX5TybeJNvE/BqL+wWr+MsaEx4lcrmMo
VTmUxnKVrQ69qT/W1IZpdSuZn7m3ugBLQzBwaCLu+URz7p3hBeVcJO9m9Ni7mVed
auwtduaZ8+EfqJtNBSUBibtSgoqKozVeLB0GFxfJ2jaBVVFyHPnu5UOPqYkx8CbX
4a9qQyXToD7d0D+KseL3HKLTjZx5KNs8a0g9BRGrDGKN/8wjzbqyCt0iZmcxnBLz
sHUDSqg08ivBhWc6QlduVKoW2mgZM3uB8A4DJ86Mhc8ts0u8k5v0OoIU95zaOYCM
1BSYgV8pojKDj25DRz6L6rJPCVTcFa/lyI61jhbx4ZdNhxso0lLit5PYe2HbBSh6
FANJnI87jVa13WgVJXTs25HZVmbB/HxLVPKoWkcJbYRXi+jSdfgcluUsO8Zii8+a
DaoFq1W4l608L7NyMnlifbUAuw/G8rlq+HItud9Ucyf9aoK+NyLP5HXBFlcq/Z0y
HtUghGaYbWfMQOTJzaGw66xoXj2K1p7kgbwGZQ2t6JR2Rj2jTx9IWyfKftmc36dA
X2rAr0XF5hqT53go7tuJbFEngbXPR3zG0O5LsdU6h3K3fkWAJ6+tXkENosuTeORB
Ak+a0Kc90X4bb7vpMwKcmbTmqeEfBYT09qNfrzlaLJvOuG6PqV0b/Wr0j2XzG7Ph
/UpdxItCsPfX72RGqJy5XDSaIild9rxJ8LBt/EGQMKpVqmBM9cVfI2NOaBkVj9s0
kcdeNw3YzXW2t2GVDUdXRHixsMu569HOIU+9GASNQguZsjiXlX1KOHBPgXwtIVm/
cmJRQO71dSx+k1HuysWpMfvfIRY20lRp2r4bn0jOM+EeknoDl7gufvAOYvC7oNKC
2BHhFAbLXbIZ1+1ipwD7C4NJLJ3pbiKyLjCxSdUVwzbtLAlLE+F9Qfw725ei9K2D
coc1TbMuGc3uoA69Yq6DpruIA0g06cczFAyHwiEzE5mLrYARpTczM7HXgpjoJFGq
2sxvCM7+LQczEX4jcBXmkXSmHw6cOJdulSKHgncWktAtMzWnml2GQvERophGsNIZ
zB2hVeN9ax/GTyoZjoDaZ+hSpl0pMLX+fqQnetyzdX1uW3FzdZ/ySpRm7zTzO7bq
ux/GZ2rg1sdX6WluEoMiR3jB1W7TQ7IVBgR5v2MHKf7oIZEnzG128pmi9+l5JXWi
0g3i3gkhN3aorhc9GP+8T5qfbO+3m95qtrwCpeohD2AuiPfAXg36laPjRzjS1pvS
B6kZ2Jx/yKrI3GdFvYoi9/xcaM2/x3UwfqDOzhzrzsVwgPEPKpwECSVsqi6poqAL
0GiSeyYNV6anAUyeVs/T+zpH9vft6inGZrI1Ark+PZm9pWjUR2VWzxb7Nw4z1n/J
fUjMEZL8fSXL6npPpfwG3idhc32kFr+wJHvIvSVaTKhEPvrJvKI5D/mefA35MHFP
QIgv4lDD3eawJZIOf7w1w+Oxy7lEk2fnMs7vdJ+p1YQOczLBq7lAK0JLlmM/PyLn
JlJwxjYo1U3JOqENLd+GkNeyOBgI9wQgdW4JdL4HCPl2fyNUQrgyWIkHFrhFibUV
9Qh+y21h7m1v2O80vtMcW1fInEMKDdYiKO/pc/3oY6bTqyWEju8pE6HPp4eOr/uF
BvRVJRqfKmOZvhIEng6r4q6qRDCtH6J1BdMZn3CXjx55FotLH1y8OZt2GSUTOgWD
IeRs90EXh9pGTO37+NRMSN5kFGgA5mkkTjeX2X+Osz+Qn4eCf/pDblz5n4pzKvfE
hw8O0pdolQzBpfV2+M8EWTE591xyo2jgAEFMUDlXqEW5CkkD84LCjU60edS0sIvO
eId2vSU9eLcqsZeyMPP0znkruEmwimsUc5liCR2x6OBx/Qau91uZpH5JkmJwuffF
P7Ht/qfX+07WZSJCOqhbGnt2aQ5X07A/6ap3qFWwk5uxXNlLjEzNzNYQTJrqhueN
kVdT1Dno6M7DAMFDQlr+5eT9qWcUsKz1M8oRW1YDSdQGvfVeazVCNYaF5vBFS252
ktR3l8VfZkwDBI4IULCKN6/rAXxYIqsA6LlFtfxCa/4VocfDSHI70wFFMnz7hpCR
hGHG5++fJZ/JPhvVlIvck9RMHhmdlvCupaJ96OPFs1aNtjwMACLiFW23PLnxKCPS
LnZVNHE9Mk3SeyYW58YYww8CVYlGL9LFg1wSIvmF/KARTQ4NMTMjY0rbfM4kC9DC
IDvgGNc7cnD8iGhmbSYzQfwU2rYWlFyk06uzy+l4a9z3yQ398ooeo/GL9DZfLrUl
3zEyt2JvRwtIACaZyRyVbUj7QvTdpEsYjmPfaQSxLZs=
`protect END_PROTECTED
