`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9pxNITY13vkD2XAmpgEBHnH5qiGTWMhGn1rxeheQAQlryCADIe+ZXFk4nv7N8lb
S3NxdRm8ju7YVAO0cgh99w5k9ezr27BrhUuNxF2ax5p12bYgdbDdVahAgTWusoCD
eKqIbV9T+DYDWf1WLHkQLPRfkc3SJcj49mRTjq0K4vCZdGXIdRz8xwl12gyUac0L
Q2eJ/UT9iKdfSbEfSCfMocVazott7dR1F549M2Aa9FmKmY4LGwc+0h9aRmwjRhdF
ce7WX279O50pKDozYXZ1SZfC+gyEM5J4qPy/nnlT1s/ISdsPOddPVd8stjSjuTKF
455ViL5NR7iuc2GJ4Hf+Kc1VFk+pYfhjnpdwMakb6Bwq2gcSLmrp7RdoX+EaBxWk
eeH5I54zHGqCr0xbgUIWm5jSe4FHNMHWiERUE54L/t5wpgxWxU8t7rOYpKpnjawC
MDT5tMaOCeK8F65rhIv4+zZlCp9ahYpykRXu6snv4lA=
`protect END_PROTECTED
