`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7mgQzDUe8gkqz3SGp0L7brBZPoA0wOPYrvoq5D8Fmt3qo7u3626BMT9LsJpCbgl
O4+UzUcYpOBbSZdEpfCWJT1neQ61M//00/dTmMBc3R9bpKFWqwzMaKhyWaEUSID1
GrI3AtCEBwUT92n4gH7AbqyI5PrQZ719LkDGNv0j4oNZ3byQsvjnA8RToBCwKaqn
8yiulZLx7NwTbumHcPPqzgH67pW3SJsvRoLx8yZRchSxgITlVZHAdVwm7iu1c9db
76pTCcdQx3igwPwemiK6/HR7RiNkiZgNqGEGkGvXJqaZOt2buqJkwAc+4aGMiikj
6uVF1StUWOcUqrtYswuMRTtk+QLgWwT8KOAnproHrmv3YASgae+zflYaUzVBHYSR
JCSjaxX/To/XUm4qMxUl8cwxHi8pwBTpZvCkm3eBO+5M0DIos2W+bKYEpXybJNua
4zBk50ulcmOYJ++VX/ZkGVWZV+C7vPzJkJprS4k9OONkqN+IyfqROB8DCxavAi3Q
y14uY6d/UX4HfG+IFVgYXXRIzPAwGhVlg4E//Or4ldkdMLkeB340wGRf0NNHVzh2
aLAVxsPN65MbqIHjiwNcP8GP3R1VXTlQs4blQddvmCbEbGm3ckH6/Yk+xc8mIaq0
rZPYbTZluJcFzf4XsIE0kZ1893bFaPlrvsBKxl3UbTW/p86KMoewdBCaecBRFNIK
`protect END_PROTECTED
