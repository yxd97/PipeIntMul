`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyCvmYDBrkC9gF0U4IiB413+DIoCbwEbI9j4+E+C/mv7zxnK9rGaOrNbHtWsYoU3
MQ4fVgChEA0c5zO6vCL+IS9fieOsfaSLbRipGZyZneqO55yv/JZ4QEL4mg/xfJEq
9ljHw2BKouloVFP310redIXFZitTxl4dkUSki/JGpAPgZ4hcXtgip8kPqhm1Fp3C
i9Qd21qAWlw0OcA/AeIeMpErJg4eq3xDBGkj5oydJck0uopK7lJW9Np5ixGNFHKK
9LxM32gvSMi2zBHikkSYkZFT/mQrcsArSGyJ3v7IGaYHGPwohltbq1oHYHj3fKSE
QidXLWHzTUw+kzr7BBG88ezMkJN3Up9qoE2lV6JEZMggxePRCzFkB5QWMqJCN0N7
Z3hY8DqFwZv4NOQ1/cZbW075sByz/eN1vQ2hvkko+WYIEqxp+2wwtW1t3Xhdo9tA
LmvAQC2Hs/aKzrhbU2q16b+kQEpdOkNe2UnHJmQ7cBmLtUwOJKHVh2hkSv1GqVW0
`protect END_PROTECTED
