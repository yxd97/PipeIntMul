`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIyHCGO2+1kH503wEO1/NE+OouDZXZc7yaSg+/fVsH36NmfFA5xVPAXk0NJ8D1hp
2mAXZK5c4F76JlWnc09qNHohsVcSK853meV7b5Hc/xZfC+rnzsDD+P0TDnO+3AMh
7ceRn+9vc3N8qofLtwLG9XHE7NGbf8eZ4y04xFGVHfqSkpuSxev51ZajJmAxX+0Q
n4XFUOXaX6k2Fj1eTWQwxUT0Xw0apSY0ACdcLAMM964vJYQN2ejD3ItM4r4y7w46
QXRMdgbxPFJGQDX9FERBqaPtClKY5QVCjeyfRG9s24UXqj8mFu/8Cqg7Uk94Fpf1
1laifLc/9F31mAZ/eQN/mXF2B0y5+D+tsFU95R8Yjzci8HLf8jfcpfVY2Z+ugAEP
+3HPaFYN4yuqMj0ob8EN3oxqJvtGiHf2xNQ/32TJGuQqqJLkn8BUj/aThUixmTbm
EAZgXAH+8s8D8ugSgWjA4dotnrp9NYOPnOP1a5UNkEiLR83x2ciWrDociaEFy0MM
bxenzD4iBAj3IWCSdV67OD2iEjMAIhkpZ8J2HpmvbaT0dBOmDAp73auJPAsngnsj
GQT9w8rwdEIzAWvQ4b+MhNjNtuZh/ocvK9RORG9AIjCwT2Biop/gkr0sfuKKBwHL
m8vME7lffqI6AGW81NQuvMaaKR02+LhV0dWfhd6id4ny9TlTU0odQN3lVZyUfcWo
eijvhXPKwOS3H94mGOHt5fzBYkrkBWOzjkuGQiwuW9iGNgQoeeXTHjKmEjNbdFZa
iIuhq+EwyfHC48xCOixcqO8scWZbL6yxu8fhv2EtE+SgLKkBVK6MNEAFYhsdXsh3
R0YFMU4155aUu5jJ+m23t7ENVVoFWGBsO5s+7PGIdCmFVYZ51Parzej9Enp9NPp8
T2qDatB8zrIOuFhO9VET42/MGso32tqCPkWP+st9DqfOFXdtByqlQss/eT2c583M
W7unJUbLaAkb/gc1/4cazt6Pc7TmQSYo9+q+XvYaVrhjWY5/z9i80ibbnCtbHJ+b
OsRuqSzkao88QLkwF7K4EDLx2VH1j3HwsHYKhIrRH2EJVzlRU6R9jP0dmF4xfaNk
1m/pcJSP+nlxzpbP66dc6FDagFzhrTQM/zRpHHx3+nWQl4TuRrp6Yd0wOYasvGcX
1hy7rMXGuMzmIEO4eUCxVdTNpRSYecabT6Q47OBo2lBS7h55TzP5v0Y9596GNHDx
S/UocQrdGWU3Zhn2KBQ2BuScHIpXlBHs5rjCteYEITF7uxB8xwfkAuV1/pwzX/Sl
ZnZ2N9GzgZquLLAQpidj0SrifzVDiG3oe5jf2KHQTF2XtkkuGqhgBeAQv8tyELBv
qTdxabZiv/F4yinkHM7j2pMLjXldl4YyiUeeyyQbFjVQ6/XWRMFjfXEge4/W84DR
Z55/CUHK24zhqtGDw2U747+yvX8DDCWH7hmFbUDQMhyFNEAqph5kf8urm7EQGDPZ
wFQOGKfkGYU4we7U4MXRhmBUj0rmRV1rrXe/VIaPh4IMEbHRZvUNV2ABXugX+Vjb
o+cfCI9AE7rPA30pGgfOoJWutclvDDuEvkvnEmlOwGidB/zjnMlUt0BKv/Sw+Vfo
`protect END_PROTECTED
