`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4MGJLpOgu6EC1N2b441GdYFKQk5tX84KvJC+ukWU6f87JmPGehh4HqZPfI4nGjAt
+63Kgg899FMlcTHhCnEtWiMWcok9L7wxTziFQVbLsqTTc5jCo/f4vxW65OTEaBx8
goYK+bTh27SHvzpSvXhMaRfSQPKJeDiLNO2NNZjKbgzt8cRS571EUVO7Ak/AwC9+
qprWA+wuEisdm3nH74ZbnRKRbRmmCnGjiRUnCYYgtf0PeLGInKsznaKMSmFWqVKc
xSq6rnyPqk4kyfjmqi/fSSeokf/hLOZw5RfSdlABLQ53WfC4gRtRCAbYMHvwFJT4
wEBeX7/QJnDYM1xUMcb28IKFo4y9s6+cyrCxjIOZ/75L1HW+4ed2in0gnq9gwvSP
ni9sUu/vb0FnWuDiD/MNuyiBSkWKKLrV9KZWniMXVpaQDLGpmdiuVLd1FP3C+4dr
0vpLHUkFoFnmOnkzZpkatq252FVPrc0FQDLEzHr3dFZw9n3tzGOvY4az5oE6oYjG
j7LSbFGropxpkmI7FR6i0wRlL5cmaUzR7+AZgPc3elxV3aspzfohB/roa/McTyZc
QaZWCnfDXR4MFQ3Q1mFhPCczdHXw5+smQXjU8jN7YN0=
`protect END_PROTECTED
