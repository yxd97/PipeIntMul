`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Balttgw4Uhy1tD5KZ7Ur+aZR4UeOUCgX6e56i7EazsIv4d2wLEmflveasHBnV1UH
m7IfYjOz6x40stjo9cDd39LxS1aj9u3CGLbc85glsXTVwVxs7KlmPiIk7OUGNz5o
KRJFpyS8xfgyUEagV8oEFt+mSJV1HzP7YVfIEbXdo8TbqMtRFTZJ/mXQr+tKd2CD
AA2XXIfp13idx4ZuUV4DPcWa1ocCfAF6rOHn1TUv5bkj4pWkjRFG86pp/fCxvU6U
CvlbPlR15ksMrheWrPHE5012e6cBAP1vZsVL0lXcDTGUUIMs4HQff3X1bsAlJAl7
NyAy/aD94cMHnKeK02j8RrvFk+DzOPn4pCEzeMeikLwA+Ke6hdUotVTGRh7VJD7H
HTjgKDLkyC+FMzvNkGTNDL3x3zw3FM4EPxPVCdM7wCw2sLEP+AJHqu+Wvv/aTUrR
bxZ6tIkLSWKjIrjPoMRz6NYebUgXV0A1W3T2AwzZ5bQDxF+dUMk644QPa1/UIlMG
1M7OTcWfTuqhhtqiHU7M7oMDnYH1/gEiGbllgXZ7C3OkN5ZQ349lFPurRiRjkNN2
F07P7fVXFp1ajCUrwXURUFZz832JRYQRR2aynTyBkfAYOm5il/Is7Qwkpyu6JbR5
yqNs/BAEE9Du+x82+vMMHgUIS09i9M2gaE/RbrMdxlxDYNJtvpsuXSE3zrBPMpVu
NnYxG5DdRbwSLFERHi0JuVl0tlhdRTjs+SB6dm/WONWRGYCb5uoFFx3YLeaJ2WMj
FGWw0NTnaBqfLr4cIh8mSmINpWtmEO/yuL9oApsOhncPU76fhsCK3+SVmxK0E4oC
pdcYoTpM7b9Pep3Fd/TB7uLWK5IhIHV7Ac846U+yzjg=
`protect END_PROTECTED
