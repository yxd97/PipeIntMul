`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oOG0jUDGsP2u92tzWlDpKduebCSIVUEabIlSJDQvbuDXf+gjtlvi+pZn+pYqMPb/
ukZsKkfKKejTxlbl/IozIzNyPuWkAK7oCGPIhNgIYimp3B+0q0+vAXjIqnigNBUW
fliCZcsAJTw74sTBpmFweg1u0bPHZmesTf2aGhVuwgqd8GK+sOmSrVCFn0faID7W
Ph+oJZk27MyoISGCLWSU01Xr0dNkdwwOrnaWFKm2sMv1UwUiR7bKA+YgsQdbf6eS
I4oToHexWOthCKzw35uT2ZF8lc/6Xkemc9oIhvLLXCi/Do1D71xMt7sDJcgOy9Jf
KEfno22+H584tJsZsyFUkyGjL5JWhgUUkuTKXel6vfADbRiwUDNxv37fD+NlRKlX
ECQY9tR8nNRoLtUfJ52ZCEe+m3ulWYqo9sDNhVCEhgwPRV9tKXk+k2sRvmiYBewN
n5a4bYjmwWlzTGpIpUQSYQ==
`protect END_PROTECTED
