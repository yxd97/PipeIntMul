`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8z/qyUeHW6sLho2mGsWSe5JjQUoSRLDvIsp8k7EWfb8ivYE8LEVz0hVKNTlNyx5v
ZK7SJojOm8mfXz7sQDUaqXdd5GOb+fYC0JkSVsU+PnBd0MPhkEmrwwCEYFWQtIIn
ITYuvIsVHiqKK3Aj+GSiRiOnirHPlKMFfLe7O10U4eH6Q7OWwOy85Dh7emHe3dmp
NeF4nIkhseg0L4eF2NPMhFf3Nexcwuhhef0qcinQVphpM+3huJuL1NvoMn/l7Zc8
zeHifXSQxi7SOE6FVzsNNjy4veaVzamEU885jHVWESCCe9NE25WTgtRmfUF9ouPP
eqRnuzWnUqiewK74dYv7NX8lC6KA1OiinYv+q82faFNX6TACO4vfwl0bXj2P5r6I
ly6qPAKpKAfok9eLxCKe0GncCdnH5UYf9jZp+MhAHwXy/sGoByZhfoZhPZGRtFPS
R1rBjZOapQXPghlx/L1NE2ZePWxd9WVu4uTRWeJig//W74nr0OV4anovo4oRp7k9
`protect END_PROTECTED
