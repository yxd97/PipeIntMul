`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epj0S6+nAkwQxOfbRoX3oiFhexZieIsXok6MAuS8mtqp7zufnIVipIq5voFqB0Bu
cMIy3RMRI1uUMDtTOcNKSw6UZ/DBe0zWF4FJSfMYQcdcZTJlSd9/z5+pGyIv2ek7
wW0ipmIo2TtUiiQi8fuQs1QmYU3kOjatR6eANKv/DcnV3YUR+eAFgfrFMcd8Zhw6
GWbxJsEuCZvLqSeVQoeqqYH+mTkeV6z/gBZYRA9/wnVR4S+hzFf02i2QduD5iebw
+NJqXIBxD2H9gn4e2guS3UWoCev9qzSQCoH4xNewUS7rq/BqZqXtaw+Cew3xXGUC
enltq0XmayItCC0sybYbVf+DUCYgvd/wGICPS5PIrRZghv1oJqFzMRvrvqdt7k9G
qHo73ge230mmwRPBvekt3Kairh5reKoFQkqpA2oiOmRAwqhy9MBXIO1LJEgnIm4y
hv31B7/uC8+tOgx2MC7I+Td+M2drf+YT65EKUQAwg1NiqzrO/7ijPUtjJ9HHowQh
pLGAjtuqwF02SBCAsQc1+dNat5thKsPx/BSbeSgldwK64tPDW6o8Ne0mW8aNFV91
KDuVaxlURU3q7FwLgwI3WjykOObhYAoWdHaEjZUGVqzzG2PPU1BaKgnPqZOXpn4q
T2w873KtSqiQ34Z5Ftet2oKO2TXMO1HDpA7w+Nnq4uHK56mG3DBOfWy2nmXHPUf9
dTTNCkavc9/hnnr6kZUxe/Y8aIWqI4GHkHXfL6ZARebugrMHn7I/3iTIJ2gSK/ar
R9vqdhbCS7hzMjKiaefPjv6gVhP/UOPN7Eah7zvXpxMDvUoDP9qgdLozPPn6QWp+
Xrso84Bq7lZC/0uTlSZbXpOzenT7H+s6R8g2Qo+t4H9UxOUMfUZbNW5qZ9gISoPC
86XX9LvHU9Rwuky6fQ3Abbvm2Hzdp8Q7ERqLQN8rJzVBRpzG6uwank+hbxG+ThFD
/pUhjJ5pPKTZOXQOvGv6ZHyvggkxFW/4k2YlLEzp6fCfjoYYgfHBJiiXILaVFlE6
l863Z1Y/9WccWQYRnUD6wtA+1/7uhnO2rKFkZSjuBOnzmLVX2nPtCgZtDThx2toh
7g3c31J39Niz6MJHI0tevRwRkscfAeSqZAPvPU6NRI2imn1xV7JR+Y5ymC3tOP10
kzAZrZSQX2gaW7GLneQjKgZzd9YqRo2uJzknAufUYA0+9werAgG6GSDxPKhgtV9R
llMPyedStHqS9OyIaFkSl7ROMJ6gcgxLUyQWTFvCNFGX8G84qnZWQh/6fE7IsaMR
+vE6/SGq6yNmQKMLYQNwfjN1MA+vZpwszEKZDspEBNCutJ7UBhqigAsYFBYCBAvb
9ULee71fPMiKSPKAwvsOE1li/kd1bCycajIK+Wj1VGQ+nXxkPt5Do6P/ITrkqa5p
RRQLheNQdEioYCzjErt98ICW+dNOkNqgJY6g0aReNYpXmh2AlXrTYL1VfZpXpiGb
sRmkZNm8TT193Kr0DUjm2Zu53ZpWmIAympGQoDi0KNC8AR+fQA2waHdJML+Z5Nwy
`protect END_PROTECTED
