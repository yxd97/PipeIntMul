`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Us73gVBvRJ+DAqkIxxY+igm6jrpULbL/eKvMyyptlzPokD/xcAv8kqD78RUCJnUD
w6nvA3Ev2TdcUKuzvXif89BircZizmLsZxgt1JXD4GEVA/+bAE+D5m9xRR6GHiza
eBqusrEV+f1x/nFvzWesFUV4d9wcL7lYmBfOA3PG8QI/WWBiRtzxR3YNi5fRwFSi
P/1OecxH5ErbJAIn0P58dKmyYEEfkyWbthwBS+EMUll8rCxfAciw2QvTbUL4Kzcy
FzlTiD7902Z8H1y0ZO+fzkBf72dthqEeK5Y6VmhmwMh7cHALc+CD4emnFEmIrtoL
Q2KLoNqhBltNXQxqukp/AnXWOZGlsO+VBqNHyiLkOGH4GQAAQFNkrKWJI9YS/+T8
VjTxOJTe4E/f8nnOp8TpRHgpgNahUkE2ixDXBHUFgqNjWllLGCVVRGKcF5ziEkyz
3UHDiBxb1Ev/IsV0NoXxdTyIdtYfAv5A4+8/1GcYIEbdGg9RH4JaTTig/35CwAMb
HjRx4CR1SJSU+0WGgwsYUt1yGvHUi7CcRygxCU7/cdUGIyWFNqV/T3IVZtQ29FpD
MwuuTXqd/ZDaMnTDhaQQiRIF/9qCgxJoW3xN/P9JF5v1DM6x4fe1b2Lti7yGNgc0
DKM8NLlrjyiTCSNyc3YSAvkcmyCeB2Pj7Rfh/UznXvsY5sjfkIDE6ZRQ34zc2RO/
zcFf6MXRPRgstdvcP4k+QKm1rW3kRVlWwIRrtleVRYNx/9TEWGgFlH0/KGwOBU0i
qWkF0a2segkRGCsvt+/25uhcOrz3/Um3J8h1gjbBs3xpQNDeD7oRM6rk8XqppwVi
h6hTbUUC6TEgnQF51eoZrHPfbdiDDnI4ppl5jZmJ3H/vWzMCwR6qAB0cwRyN2mzA
`protect END_PROTECTED
