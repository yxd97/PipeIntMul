`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BG7CseguKRK0O8EShGt34GJWTTYwHkL5zHu14IWvAldH0pO1Ov6dXZiGZj4sshEH
X6zNXjnBBVM9kTll5uDtqSjZAT9SSdIFUYr5PqHKET2PjCVwwDCv5ZuP+jMj65d7
uj4tOVfgTMDU+lf5suD59cvNWPoAlOyo8S/PeOyvsFIwj42Wk7gTYvHv7wRMBtQM
KqyI9nb/ovzx3QjgodIG4oiMA3zZBQCIfiWgtuAKhZh3e/sIjA5pkLnRRnoz4QGv
1/mslA4zAkCUDjEYFRvU3GEjUP+J4NMKoZrJ67VS72T+IwV4jgzApKFst0Jo/dKD
yxYydSimP7MeTI54PXQiA+21+llTTFfgxN740HrbVbUjL3Di3+G4jHq/OIs1zwG6
AeStqLWM1gPtcneU9Ii3nHE7RgyD+PlYRC4dhxWyWmJkspIpySMCLemEd12ncoF1
XogWWQXtSP6Ygk+UJyZtgrNIqUOIjjcgRjCRC4dtkwmE89HGgIZd3+/cVs/fueGM
`protect END_PROTECTED
