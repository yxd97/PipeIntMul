`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nnHx7wXn3u1kqA9PVPpX80RBUtuJcpjpF5wgqwzI+KbPescYWdnvT9E2gO4BSvKd
B54EFL32MGJVCepaWaPPOB12Xoq+XQMc2auUvDI826g/iaMKYZxK8Eab2cvJJKz+
MdzCglT+NlLu+61M/Lj/XIGN9qDaiKuopz2eVOoZr7NBBO0Z/8rdG774En+DAkpV
zq5YfDixLooMhOM0t4nK+H2EnDNdHyrPB9zu96OhXnEUPbSyHX99EV785/yI/Y0Z
sfMAgjrgYUaJ6GNnfizaU1iqU4c2J80EpyiIboGFfyGtZSgyR/5crA0yIUkqslJv
nlQUw/nwcoWH3KcF+MtV2T//9C1/H9LYdaspOc7pBc7fEkM6e6WmIhtfNhn3ifxB
JO6+aUyxxdpYHdy432eZ03C19k70U4a3xnfmLfv06a9dHcxVwEbOZvZ+oBW613J3
`protect END_PROTECTED
