`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZVmch6lXsD3p5hmxuqChpnfGz/CaDbr1oFOX+5Y45Nchoj6ujLQqyExSU1pvtsab
kZDFL0QdNxsQ6Y3dGcuDkMCCVQVF5RpylmeTAHEBmiXSmJ6er1DntPT3tLv3LyH8
QHKFfR9t0Wz0tjJ6oBVZUlTjNlGmF8RRqdG3BpBEGpAvN2CgIzdXBj0pg+kwSbRT
Z6+vJG+FigLHftlSB1lr1NlL8GgXx9iDZlf3e4ydmsrysjA2kdEo8Z6u9+1wz90v
er1E5nGXcsA0IT5IFONOvx3puvtL1/ECLFND6NNTuseQEfd4bICVecfLsYNU0En/
tSNkhIiwwtGjRR5SQU8HKQ==
`protect END_PROTECTED
