`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lXsre0D6vworxfLRqxmW7maSFGvOS6X1XN2hZmFgLQxA9OGYLJspvkMxNSVqREy/
QRnAvg5BNvapyf38C8/A3zzWVpwZ8CFwPO6V4ql/DVvbxweqJlIIAe+txvPWrPoz
9jbi3I5MvnH9783RXdqKqaNzr0AHhRrwyytX/8tpLeUGdVLKUnijaDNijU8p6jaC
Y7gwNXmd2cBCjgPuG0chK4+TXZUbY0utPV6cNV0WjVpWVmCXd0eifpfZ5olQZcMq
6WNvA8AQ6s/0vwwNrx9O6oPz4JN4+OwVoelN1DDxt6ny5F+nFhV+BSsDN5DqtwVh
Q3GuTe6OK8ISN57TaxwNJw==
`protect END_PROTECTED
