library verilog;
use verilog.vl_types.all;
entity PCIE_EP is
    generic(
        BAR0EXIST       : string  := "TRUE";
        BAR0PREFETCHABLE: string  := "TRUE";
        BAR1EXIST       : string  := "FALSE";
        BAR1PREFETCHABLE: string  := "FALSE";
        BAR2EXIST       : string  := "FALSE";
        BAR2PREFETCHABLE: string  := "FALSE";
        BAR3EXIST       : string  := "FALSE";
        BAR3PREFETCHABLE: string  := "FALSE";
        BAR4EXIST       : string  := "FALSE";
        BAR4PREFETCHABLE: string  := "FALSE";
        BAR5EXIST       : string  := "FALSE";
        BAR5PREFETCHABLE: string  := "FALSE";
        CLKDIVIDED      : string  := "FALSE";
        INFINITECOMPLETIONS: string  := "TRUE";
        LINKSTATUSSLOTCLOCKCONFIG: string  := "FALSE";
        PBCAPABILITYSYSTEMALLOCATED: string  := "FALSE";
        PMCAPABILITYD1SUPPORT: string  := "FALSE";
        PMCAPABILITYD2SUPPORT: string  := "FALSE";
        PMCAPABILITYDSI : string  := "TRUE";
        RESETMODE       : string  := "FALSE";
        VC0TOTALCREDITSCD: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC0TOTALCREDITSPD: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        VC1TOTALCREDITSCD: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC1TOTALCREDITSPD: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AERBASEPTR      : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        AERCAPABILITYNEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        DSNBASEPTR      : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        DSNCAPABILITYNEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        MSIBASEPTR      : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        PBBASEPTR       : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        PBCAPABILITYNEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        PMBASEPTR       : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RETRYRAMSIZE    : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        VCBASEPTR       : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        VCCAPABILITYNEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC0RXFIFOBASEC  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC0RXFIFOBASENP : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC0RXFIFOBASEP  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC0RXFIFOLIMITC : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        VC0RXFIFOLIMITNP: vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        VC0RXFIFOLIMITP : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        VC0TXFIFOBASEC  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC0TXFIFOBASENP : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC0TXFIFOBASEP  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC0TXFIFOLIMITC : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        VC0TXFIFOLIMITNP: vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        VC0TXFIFOLIMITP : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        VC1RXFIFOBASEC  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1RXFIFOBASENP : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1RXFIFOBASEP  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1RXFIFOLIMITC : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1RXFIFOLIMITNP: vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1RXFIFOLIMITP : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1TXFIFOBASEC  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1TXFIFOBASENP : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1TXFIFOBASEP  : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1TXFIFOLIMITC : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1TXFIFOLIMITNP: vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VC1TXFIFOLIMITP : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        DEVICEID        : vl_logic_vector(15 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        SUBSYSTEMID     : vl_logic_vector(15 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        SUBSYSTEMVENDORID: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        VENDORID        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        LINKCAPABILITYASPMSUPPORT: vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PBCAPABILITYDW0DATASCALE: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PBCAPABILITYDW0PMSTATE: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PBCAPABILITYDW1DATASCALE: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PBCAPABILITYDW1PMSTATE: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PBCAPABILITYDW2DATASCALE: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PBCAPABILITYDW2PMSTATE: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PBCAPABILITYDW3DATASCALE: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PBCAPABILITYDW3PMSTATE: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        CLASSCODE       : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DEVICECAPABILITYENDPOINTL0SLATENCY: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        DEVICECAPABILITYENDPOINTL1LATENCY: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        MSICAPABILITYMULTIMSGCAP: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW0PMSUBSTATE: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW0POWERRAIL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW0TYPE: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW1PMSUBSTATE: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW1POWERRAIL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW1TYPE: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW2PMSUBSTATE: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW2POWERRAIL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW2TYPE: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW3PMSUBSTATE: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW3POWERRAIL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PBCAPABILITYDW3TYPE: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PMCAPABILITYAUXCURRENT: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PORTVCCAPABILITYEXTENDEDVCCOUNT: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        CARDBUSCISPOINTER: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        XPDEVICEPORTTYPE: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        PMCAPABILITYPMESUPPORT: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR0MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        BAR1MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR2MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR3MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR4MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR5MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LINKCAPABILITYMAXLINKWIDTH: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        DEVICESERIALNUMBER: vl_logic_vector(63 downto 0) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        VC0TOTALCREDITSCH: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC0TOTALCREDITSNPH: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        VC0TOTALCREDITSPH: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        VC1TOTALCREDITSCH: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC1TOTALCREDITSNPH: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC1TOTALCREDITSPH: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ACTIVELANESIN   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        CAPABILITIESPOINTER: vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INTERRUPTPIN    : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MSICAPABILITYNEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        PBCAPABILITYDW0BASEPOWER: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PBCAPABILITYDW1BASEPOWER: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PBCAPABILITYDW2BASEPOWER: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PBCAPABILITYDW3BASEPOWER: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PCIECAPABILITYNEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMCAPABILITYNEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMDATA0         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMDATA1         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMDATA2         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMDATA3         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMDATA4         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMDATA5         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMDATA6         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMDATA7         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PORTVCCAPABILITYVCARBCAP: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PORTVCCAPABILITYVCARBTABLEOFFSET: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        REVISIONID      : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        XPBASEPTR       : vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR0ADDRWIDTH   : integer := 0;
        BAR0IOMEMN      : integer := 0;
        BAR1ADDRWIDTH   : integer := 0;
        BAR1IOMEMN      : integer := 0;
        BAR2ADDRWIDTH   : integer := 0;
        BAR2IOMEMN      : integer := 0;
        BAR3ADDRWIDTH   : integer := 0;
        BAR3IOMEMN      : integer := 0;
        BAR4ADDRWIDTH   : integer := 0;
        BAR4IOMEMN      : integer := 0;
        BAR5IOMEMN      : integer := 0;
        L0SEXITLATENCY  : integer := 7;
        L0SEXITLATENCYCOMCLK: integer := 7;
        L1EXITLATENCY   : integer := 7;
        L1EXITLATENCYCOMCLK: integer := 7;
        LOWPRIORITYVCCOUNT: integer := 0;
        PMDATASCALE0    : integer := 0;
        PMDATASCALE1    : integer := 0;
        PMDATASCALE2    : integer := 0;
        PMDATASCALE3    : integer := 0;
        PMDATASCALE4    : integer := 0;
        PMDATASCALE5    : integer := 0;
        PMDATASCALE6    : integer := 0;
        PMDATASCALE7    : integer := 0;
        RETRYRAMREADLATENCY: integer := 3;
        RETRYRAMWRITELATENCY: integer := 1;
        TLRAMREADLATENCY: integer := 3;
        TLRAMWRITELATENCY: integer := 1;
        TXTSNFTS        : integer := 255;
        TXTSNFTSCOMCLK  : integer := 255;
        XPMAXPAYLOAD    : integer := 0
    );
    port(
        BUSMASTERENABLE : out    vl_logic;
        CRMDOHOTRESETN  : out    vl_logic;
        CRMPWRSOFTRESETN: out    vl_logic;
        DLLTXPMDLLPOUTSTANDING: out    vl_logic;
        INTERRUPTDISABLE: out    vl_logic;
        IOSPACEENABLE   : out    vl_logic;
        L0CFGLOOPBACKACK: out    vl_logic;
        L0COMPLETERID   : out    vl_logic_vector(12 downto 0);
        L0DLLERRORVECTOR: out    vl_logic_vector(6 downto 0);
        L0DLLRXACKOUTSTANDING: out    vl_logic;
        L0DLLTXNONFCOUTSTANDING: out    vl_logic;
        L0DLLTXOUTSTANDING: out    vl_logic;
        L0DLLVCSTATUS   : out    vl_logic_vector(7 downto 0);
        L0DLUPDOWN      : out    vl_logic_vector(7 downto 0);
        L0FIRSTCFGWRITEOCCURRED: out    vl_logic;
        L0LTSSMSTATE    : out    vl_logic_vector(3 downto 0);
        L0MACENTEREDL0  : out    vl_logic;
        L0MACLINKTRAINING: out    vl_logic;
        L0MACLINKUP     : out    vl_logic;
        L0MACNEGOTIATEDLINKWIDTH: out    vl_logic_vector(3 downto 0);
        L0MACNEWSTATEACK: out    vl_logic;
        L0MACRXL0SSTATE : out    vl_logic;
        L0MSIENABLE0    : out    vl_logic;
        L0MULTIMSGEN0   : out    vl_logic_vector(2 downto 0);
        L0PMEACK        : out    vl_logic;
        L0PMEEN         : out    vl_logic;
        L0PMEREQOUT     : out    vl_logic;
        L0PWRL1STATE    : out    vl_logic;
        L0PWRL23READYSTATE: out    vl_logic;
        L0PWRSTATE0     : out    vl_logic_vector(1 downto 0);
        L0PWRTURNOFFREQ : out    vl_logic;
        L0PWRTXL0SSTATE : out    vl_logic;
        L0RXDLLPM       : out    vl_logic;
        L0RXDLLPMTYPE   : out    vl_logic_vector(2 downto 0);
        L0RXMACLINKERROR: out    vl_logic_vector(1 downto 0);
        L0STATSCFGOTHERRECEIVED: out    vl_logic;
        L0STATSCFGOTHERTRANSMITTED: out    vl_logic;
        L0STATSCFGRECEIVED: out    vl_logic;
        L0STATSCFGTRANSMITTED: out    vl_logic;
        L0STATSDLLPRECEIVED: out    vl_logic;
        L0STATSDLLPTRANSMITTED: out    vl_logic;
        L0STATSOSRECEIVED: out    vl_logic;
        L0STATSOSTRANSMITTED: out    vl_logic;
        L0STATSTLPRECEIVED: out    vl_logic;
        L0STATSTLPTRANSMITTED: out    vl_logic;
        L0UNLOCKRECEIVED: out    vl_logic;
        LLKRXCHCOMPLETIONAVAILABLEN: out    vl_logic_vector(7 downto 0);
        LLKRXCHNONPOSTEDAVAILABLEN: out    vl_logic_vector(7 downto 0);
        LLKRXCHPOSTEDAVAILABLEN: out    vl_logic_vector(7 downto 0);
        LLKRXDATA       : out    vl_logic_vector(63 downto 0);
        LLKRXEOFN       : out    vl_logic;
        LLKRXEOPN       : out    vl_logic;
        LLKRXPREFERREDTYPE: out    vl_logic_vector(15 downto 0);
        LLKRXSOFN       : out    vl_logic;
        LLKRXSOPN       : out    vl_logic;
        LLKRXSRCLASTREQN: out    vl_logic;
        LLKRXSRCRDYN    : out    vl_logic;
        LLKRXVALIDN     : out    vl_logic_vector(1 downto 0);
        LLKTCSTATUS     : out    vl_logic_vector(7 downto 0);
        LLKTXCHANSPACE  : out    vl_logic_vector(9 downto 0);
        LLKTXCHCOMPLETIONREADYN: out    vl_logic_vector(7 downto 0);
        LLKTXCHNONPOSTEDREADYN: out    vl_logic_vector(7 downto 0);
        LLKTXCHPOSTEDREADYN: out    vl_logic_vector(7 downto 0);
        LLKTXCONFIGREADYN: out    vl_logic;
        LLKTXDSTRDYN    : out    vl_logic;
        MAXPAYLOADSIZE  : out    vl_logic_vector(2 downto 0);
        MAXREADREQUESTSIZE: out    vl_logic_vector(2 downto 0);
        MEMSPACEENABLE  : out    vl_logic;
        MGMTPSO         : out    vl_logic_vector(16 downto 0);
        MGMTRDATA       : out    vl_logic_vector(31 downto 0);
        MGMTSTATSCREDIT : out    vl_logic_vector(11 downto 0);
        MIMDLLBRADD     : out    vl_logic_vector(11 downto 0);
        MIMDLLBREN      : out    vl_logic;
        MIMDLLBWADD     : out    vl_logic_vector(11 downto 0);
        MIMDLLBWDATA    : out    vl_logic_vector(63 downto 0);
        MIMDLLBWEN      : out    vl_logic;
        MIMRXBRADD      : out    vl_logic_vector(12 downto 0);
        MIMRXBREN       : out    vl_logic;
        MIMRXBWADD      : out    vl_logic_vector(12 downto 0);
        MIMRXBWDATA     : out    vl_logic_vector(63 downto 0);
        MIMRXBWEN       : out    vl_logic;
        MIMTXBRADD      : out    vl_logic_vector(12 downto 0);
        MIMTXBREN       : out    vl_logic;
        MIMTXBWADD      : out    vl_logic_vector(12 downto 0);
        MIMTXBWDATA     : out    vl_logic_vector(63 downto 0);
        MIMTXBWEN       : out    vl_logic;
        PARITYERRORRESPONSE: out    vl_logic;
        PIPEDESKEWLANESL0: out    vl_logic;
        PIPEDESKEWLANESL1: out    vl_logic;
        PIPEDESKEWLANESL2: out    vl_logic;
        PIPEDESKEWLANESL3: out    vl_logic;
        PIPEDESKEWLANESL4: out    vl_logic;
        PIPEDESKEWLANESL5: out    vl_logic;
        PIPEDESKEWLANESL6: out    vl_logic;
        PIPEDESKEWLANESL7: out    vl_logic;
        PIPEPOWERDOWNL0 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL1 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL2 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL3 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL4 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL5 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL6 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL7 : out    vl_logic_vector(1 downto 0);
        PIPERESETL0     : out    vl_logic;
        PIPERESETL1     : out    vl_logic;
        PIPERESETL2     : out    vl_logic;
        PIPERESETL3     : out    vl_logic;
        PIPERESETL4     : out    vl_logic;
        PIPERESETL5     : out    vl_logic;
        PIPERESETL6     : out    vl_logic;
        PIPERESETL7     : out    vl_logic;
        PIPERXPOLARITYL0: out    vl_logic;
        PIPERXPOLARITYL1: out    vl_logic;
        PIPERXPOLARITYL2: out    vl_logic;
        PIPERXPOLARITYL3: out    vl_logic;
        PIPERXPOLARITYL4: out    vl_logic;
        PIPERXPOLARITYL5: out    vl_logic;
        PIPERXPOLARITYL6: out    vl_logic;
        PIPERXPOLARITYL7: out    vl_logic;
        PIPETXCOMPLIANCEL0: out    vl_logic;
        PIPETXCOMPLIANCEL1: out    vl_logic;
        PIPETXCOMPLIANCEL2: out    vl_logic;
        PIPETXCOMPLIANCEL3: out    vl_logic;
        PIPETXCOMPLIANCEL4: out    vl_logic;
        PIPETXCOMPLIANCEL5: out    vl_logic;
        PIPETXCOMPLIANCEL6: out    vl_logic;
        PIPETXCOMPLIANCEL7: out    vl_logic;
        PIPETXDATAKL0   : out    vl_logic;
        PIPETXDATAKL1   : out    vl_logic;
        PIPETXDATAKL2   : out    vl_logic;
        PIPETXDATAKL3   : out    vl_logic;
        PIPETXDATAKL4   : out    vl_logic;
        PIPETXDATAKL5   : out    vl_logic;
        PIPETXDATAKL6   : out    vl_logic;
        PIPETXDATAKL7   : out    vl_logic;
        PIPETXDATAL0    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL1    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL2    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL3    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL4    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL5    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL6    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL7    : out    vl_logic_vector(7 downto 0);
        PIPETXDETECTRXLOOPBACKL0: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL1: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL2: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL3: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL4: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL5: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL6: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL7: out    vl_logic;
        PIPETXELECIDLEL0: out    vl_logic;
        PIPETXELECIDLEL1: out    vl_logic;
        PIPETXELECIDLEL2: out    vl_logic;
        PIPETXELECIDLEL3: out    vl_logic;
        PIPETXELECIDLEL4: out    vl_logic;
        PIPETXELECIDLEL5: out    vl_logic;
        PIPETXELECIDLEL6: out    vl_logic;
        PIPETXELECIDLEL7: out    vl_logic;
        SERRENABLE      : out    vl_logic;
        URREPORTINGENABLE: out    vl_logic;
        AUXPOWER        : in     vl_logic;
        COMPLIANCEAVOID : in     vl_logic;
        CRMCORECLK      : in     vl_logic;
        CRMCORECLKDLO   : in     vl_logic;
        CRMCORECLKRXO   : in     vl_logic;
        CRMCORECLKTXO   : in     vl_logic;
        CRMLINKRSTN     : in     vl_logic;
        CRMMACRSTN      : in     vl_logic;
        CRMMGMTRSTN     : in     vl_logic;
        CRMNVRSTN       : in     vl_logic;
        CRMURSTN        : in     vl_logic;
        CRMUSERCFGRSTN  : in     vl_logic;
        CRMUSERCLK      : in     vl_logic;
        CRMUSERCLKRXO   : in     vl_logic;
        CRMUSERCLKTXO   : in     vl_logic;
        L0CFGDISABLESCRAMBLE: in     vl_logic;
        L0CFGLOOPBACKMASTER: in     vl_logic;
        L0LEGACYINTFUNCT0: in     vl_logic;
        L0MSIREQUEST0   : in     vl_logic_vector(3 downto 0);
        L0PACKETHEADERFROMUSER: in     vl_logic_vector(127 downto 0);
        L0PMEREQIN      : in     vl_logic;
        L0SETCOMPLETERABORTERROR: in     vl_logic;
        L0SETCOMPLETIONTIMEOUTCORRERROR: in     vl_logic;
        L0SETCOMPLETIONTIMEOUTUNCORRERROR: in     vl_logic;
        L0SETDETECTEDCORRERROR: in     vl_logic;
        L0SETDETECTEDFATALERROR: in     vl_logic;
        L0SETDETECTEDNONFATALERROR: in     vl_logic;
        L0SETUNEXPECTEDCOMPLETIONCORRERROR: in     vl_logic;
        L0SETUNEXPECTEDCOMPLETIONUNCORRERROR: in     vl_logic;
        L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR: in     vl_logic;
        L0SETUNSUPPORTEDREQUESTOTHERERROR: in     vl_logic;
        L0SETUSERDETECTEDPARITYERROR: in     vl_logic;
        L0SETUSERMASTERDATAPARITY: in     vl_logic;
        L0SETUSERRECEIVEDMASTERABORT: in     vl_logic;
        L0SETUSERRECEIVEDTARGETABORT: in     vl_logic;
        L0SETUSERSIGNALLEDTARGETABORT: in     vl_logic;
        L0SETUSERSYSTEMERROR: in     vl_logic;
        L0TRANSACTIONSPENDING: in     vl_logic;
        LLKRXCHFIFO     : in     vl_logic_vector(1 downto 0);
        LLKRXCHTC       : in     vl_logic_vector(2 downto 0);
        LLKRXDSTCONTREQN: in     vl_logic;
        LLKRXDSTREQN    : in     vl_logic;
        LLKTXCHFIFO     : in     vl_logic_vector(1 downto 0);
        LLKTXCHTC       : in     vl_logic_vector(2 downto 0);
        LLKTXDATA       : in     vl_logic_vector(63 downto 0);
        LLKTXENABLEN    : in     vl_logic_vector(1 downto 0);
        LLKTXEOFN       : in     vl_logic;
        LLKTXEOPN       : in     vl_logic;
        LLKTXSOFN       : in     vl_logic;
        LLKTXSOPN       : in     vl_logic;
        LLKTXSRCDSCN    : in     vl_logic;
        LLKTXSRCRDYN    : in     vl_logic;
        MGMTADDR        : in     vl_logic_vector(10 downto 0);
        MGMTBWREN       : in     vl_logic_vector(3 downto 0);
        MGMTRDEN        : in     vl_logic;
        MGMTSTATSCREDITSEL: in     vl_logic_vector(6 downto 0);
        MGMTWDATA       : in     vl_logic_vector(31 downto 0);
        MGMTWREN        : in     vl_logic;
        MIMDLLBRDATA    : in     vl_logic_vector(63 downto 0);
        MIMRXBRDATA     : in     vl_logic_vector(63 downto 0);
        MIMTXBRDATA     : in     vl_logic_vector(63 downto 0);
        PIPEPHYSTATUSL0 : in     vl_logic;
        PIPEPHYSTATUSL1 : in     vl_logic;
        PIPEPHYSTATUSL2 : in     vl_logic;
        PIPEPHYSTATUSL3 : in     vl_logic;
        PIPEPHYSTATUSL4 : in     vl_logic;
        PIPEPHYSTATUSL5 : in     vl_logic;
        PIPEPHYSTATUSL6 : in     vl_logic;
        PIPEPHYSTATUSL7 : in     vl_logic;
        PIPERXCHANISALIGNEDL0: in     vl_logic;
        PIPERXCHANISALIGNEDL1: in     vl_logic;
        PIPERXCHANISALIGNEDL2: in     vl_logic;
        PIPERXCHANISALIGNEDL3: in     vl_logic;
        PIPERXCHANISALIGNEDL4: in     vl_logic;
        PIPERXCHANISALIGNEDL5: in     vl_logic;
        PIPERXCHANISALIGNEDL6: in     vl_logic;
        PIPERXCHANISALIGNEDL7: in     vl_logic;
        PIPERXDATAKL0   : in     vl_logic;
        PIPERXDATAKL1   : in     vl_logic;
        PIPERXDATAKL2   : in     vl_logic;
        PIPERXDATAKL3   : in     vl_logic;
        PIPERXDATAKL4   : in     vl_logic;
        PIPERXDATAKL5   : in     vl_logic;
        PIPERXDATAKL6   : in     vl_logic;
        PIPERXDATAKL7   : in     vl_logic;
        PIPERXDATAL0    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL1    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL2    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL3    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL4    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL5    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL6    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL7    : in     vl_logic_vector(7 downto 0);
        PIPERXELECIDLEL0: in     vl_logic;
        PIPERXELECIDLEL1: in     vl_logic;
        PIPERXELECIDLEL2: in     vl_logic;
        PIPERXELECIDLEL3: in     vl_logic;
        PIPERXELECIDLEL4: in     vl_logic;
        PIPERXELECIDLEL5: in     vl_logic;
        PIPERXELECIDLEL6: in     vl_logic;
        PIPERXELECIDLEL7: in     vl_logic;
        PIPERXSTATUSL0  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL1  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL2  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL3  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL4  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL5  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL6  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL7  : in     vl_logic_vector(2 downto 0);
        PIPERXVALIDL0   : in     vl_logic;
        PIPERXVALIDL1   : in     vl_logic;
        PIPERXVALIDL2   : in     vl_logic;
        PIPERXVALIDL3   : in     vl_logic;
        PIPERXVALIDL4   : in     vl_logic;
        PIPERXVALIDL5   : in     vl_logic;
        PIPERXVALIDL6   : in     vl_logic;
        PIPERXVALIDL7   : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BAR0EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR0PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR1EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR1PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR2EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR2PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR3EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR3PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR4EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR4PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR5EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR5PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of CLKDIVIDED : constant is 1;
    attribute mti_svvh_generic_type of INFINITECOMPLETIONS : constant is 1;
    attribute mti_svvh_generic_type of LINKSTATUSSLOTCLOCKCONFIG : constant is 1;
    attribute mti_svvh_generic_type of PBCAPABILITYSYSTEMALLOCATED : constant is 1;
    attribute mti_svvh_generic_type of PMCAPABILITYD1SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PMCAPABILITYD2SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PMCAPABILITYDSI : constant is 1;
    attribute mti_svvh_generic_type of RESETMODE : constant is 1;
    attribute mti_svvh_generic_type of VC0TOTALCREDITSCD : constant is 2;
    attribute mti_svvh_generic_type of VC0TOTALCREDITSPD : constant is 2;
    attribute mti_svvh_generic_type of VC1TOTALCREDITSCD : constant is 2;
    attribute mti_svvh_generic_type of VC1TOTALCREDITSPD : constant is 2;
    attribute mti_svvh_generic_type of AERBASEPTR : constant is 2;
    attribute mti_svvh_generic_type of AERCAPABILITYNEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of DSNBASEPTR : constant is 2;
    attribute mti_svvh_generic_type of DSNCAPABILITYNEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of MSIBASEPTR : constant is 2;
    attribute mti_svvh_generic_type of PBBASEPTR : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYNEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PMBASEPTR : constant is 2;
    attribute mti_svvh_generic_type of RETRYRAMSIZE : constant is 2;
    attribute mti_svvh_generic_type of VCBASEPTR : constant is 2;
    attribute mti_svvh_generic_type of VCCAPABILITYNEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VC0RXFIFOBASEC : constant is 2;
    attribute mti_svvh_generic_type of VC0RXFIFOBASENP : constant is 2;
    attribute mti_svvh_generic_type of VC0RXFIFOBASEP : constant is 2;
    attribute mti_svvh_generic_type of VC0RXFIFOLIMITC : constant is 2;
    attribute mti_svvh_generic_type of VC0RXFIFOLIMITNP : constant is 2;
    attribute mti_svvh_generic_type of VC0RXFIFOLIMITP : constant is 2;
    attribute mti_svvh_generic_type of VC0TXFIFOBASEC : constant is 2;
    attribute mti_svvh_generic_type of VC0TXFIFOBASENP : constant is 2;
    attribute mti_svvh_generic_type of VC0TXFIFOBASEP : constant is 2;
    attribute mti_svvh_generic_type of VC0TXFIFOLIMITC : constant is 2;
    attribute mti_svvh_generic_type of VC0TXFIFOLIMITNP : constant is 2;
    attribute mti_svvh_generic_type of VC0TXFIFOLIMITP : constant is 2;
    attribute mti_svvh_generic_type of VC1RXFIFOBASEC : constant is 2;
    attribute mti_svvh_generic_type of VC1RXFIFOBASENP : constant is 2;
    attribute mti_svvh_generic_type of VC1RXFIFOBASEP : constant is 2;
    attribute mti_svvh_generic_type of VC1RXFIFOLIMITC : constant is 2;
    attribute mti_svvh_generic_type of VC1RXFIFOLIMITNP : constant is 2;
    attribute mti_svvh_generic_type of VC1RXFIFOLIMITP : constant is 2;
    attribute mti_svvh_generic_type of VC1TXFIFOBASEC : constant is 2;
    attribute mti_svvh_generic_type of VC1TXFIFOBASENP : constant is 2;
    attribute mti_svvh_generic_type of VC1TXFIFOBASEP : constant is 2;
    attribute mti_svvh_generic_type of VC1TXFIFOLIMITC : constant is 2;
    attribute mti_svvh_generic_type of VC1TXFIFOLIMITNP : constant is 2;
    attribute mti_svvh_generic_type of VC1TXFIFOLIMITP : constant is 2;
    attribute mti_svvh_generic_type of DEVICEID : constant is 2;
    attribute mti_svvh_generic_type of SUBSYSTEMID : constant is 2;
    attribute mti_svvh_generic_type of SUBSYSTEMVENDORID : constant is 2;
    attribute mti_svvh_generic_type of VENDORID : constant is 2;
    attribute mti_svvh_generic_type of LINKCAPABILITYASPMSUPPORT : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW0DATASCALE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW0PMSTATE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW1DATASCALE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW1PMSTATE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW2DATASCALE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW2PMSTATE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW3DATASCALE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW3PMSTATE : constant is 2;
    attribute mti_svvh_generic_type of CLASSCODE : constant is 2;
    attribute mti_svvh_generic_type of DEVICECAPABILITYENDPOINTL0SLATENCY : constant is 2;
    attribute mti_svvh_generic_type of DEVICECAPABILITYENDPOINTL1LATENCY : constant is 2;
    attribute mti_svvh_generic_type of MSICAPABILITYMULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW0PMSUBSTATE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW0POWERRAIL : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW0TYPE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW1PMSUBSTATE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW1POWERRAIL : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW1TYPE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW2PMSUBSTATE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW2POWERRAIL : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW2TYPE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW3PMSUBSTATE : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW3POWERRAIL : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW3TYPE : constant is 2;
    attribute mti_svvh_generic_type of PMCAPABILITYAUXCURRENT : constant is 2;
    attribute mti_svvh_generic_type of PORTVCCAPABILITYEXTENDEDVCCOUNT : constant is 2;
    attribute mti_svvh_generic_type of CARDBUSCISPOINTER : constant is 2;
    attribute mti_svvh_generic_type of XPDEVICEPORTTYPE : constant is 2;
    attribute mti_svvh_generic_type of PMCAPABILITYPMESUPPORT : constant is 2;
    attribute mti_svvh_generic_type of BAR0MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR1MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR2MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR3MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR4MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR5MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of LINKCAPABILITYMAXLINKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of DEVICESERIALNUMBER : constant is 2;
    attribute mti_svvh_generic_type of VC0TOTALCREDITSCH : constant is 2;
    attribute mti_svvh_generic_type of VC0TOTALCREDITSNPH : constant is 2;
    attribute mti_svvh_generic_type of VC0TOTALCREDITSPH : constant is 2;
    attribute mti_svvh_generic_type of VC1TOTALCREDITSCH : constant is 2;
    attribute mti_svvh_generic_type of VC1TOTALCREDITSNPH : constant is 2;
    attribute mti_svvh_generic_type of VC1TOTALCREDITSPH : constant is 2;
    attribute mti_svvh_generic_type of ACTIVELANESIN : constant is 2;
    attribute mti_svvh_generic_type of CAPABILITIESPOINTER : constant is 2;
    attribute mti_svvh_generic_type of INTERRUPTPIN : constant is 2;
    attribute mti_svvh_generic_type of MSICAPABILITYNEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW0BASEPOWER : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW1BASEPOWER : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW2BASEPOWER : constant is 2;
    attribute mti_svvh_generic_type of PBCAPABILITYDW3BASEPOWER : constant is 2;
    attribute mti_svvh_generic_type of PCIECAPABILITYNEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PMCAPABILITYNEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PMDATA0 : constant is 2;
    attribute mti_svvh_generic_type of PMDATA1 : constant is 2;
    attribute mti_svvh_generic_type of PMDATA2 : constant is 2;
    attribute mti_svvh_generic_type of PMDATA3 : constant is 2;
    attribute mti_svvh_generic_type of PMDATA4 : constant is 2;
    attribute mti_svvh_generic_type of PMDATA5 : constant is 2;
    attribute mti_svvh_generic_type of PMDATA6 : constant is 2;
    attribute mti_svvh_generic_type of PMDATA7 : constant is 2;
    attribute mti_svvh_generic_type of PORTVCCAPABILITYVCARBCAP : constant is 2;
    attribute mti_svvh_generic_type of PORTVCCAPABILITYVCARBTABLEOFFSET : constant is 2;
    attribute mti_svvh_generic_type of REVISIONID : constant is 2;
    attribute mti_svvh_generic_type of XPBASEPTR : constant is 2;
    attribute mti_svvh_generic_type of BAR0ADDRWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR0IOMEMN : constant is 2;
    attribute mti_svvh_generic_type of BAR1ADDRWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR1IOMEMN : constant is 2;
    attribute mti_svvh_generic_type of BAR2ADDRWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR2IOMEMN : constant is 2;
    attribute mti_svvh_generic_type of BAR3ADDRWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR3IOMEMN : constant is 2;
    attribute mti_svvh_generic_type of BAR4ADDRWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR4IOMEMN : constant is 2;
    attribute mti_svvh_generic_type of BAR5IOMEMN : constant is 2;
    attribute mti_svvh_generic_type of L0SEXITLATENCY : constant is 2;
    attribute mti_svvh_generic_type of L0SEXITLATENCYCOMCLK : constant is 2;
    attribute mti_svvh_generic_type of L1EXITLATENCY : constant is 2;
    attribute mti_svvh_generic_type of L1EXITLATENCYCOMCLK : constant is 2;
    attribute mti_svvh_generic_type of LOWPRIORITYVCCOUNT : constant is 2;
    attribute mti_svvh_generic_type of PMDATASCALE0 : constant is 2;
    attribute mti_svvh_generic_type of PMDATASCALE1 : constant is 2;
    attribute mti_svvh_generic_type of PMDATASCALE2 : constant is 2;
    attribute mti_svvh_generic_type of PMDATASCALE3 : constant is 2;
    attribute mti_svvh_generic_type of PMDATASCALE4 : constant is 2;
    attribute mti_svvh_generic_type of PMDATASCALE5 : constant is 2;
    attribute mti_svvh_generic_type of PMDATASCALE6 : constant is 2;
    attribute mti_svvh_generic_type of PMDATASCALE7 : constant is 2;
    attribute mti_svvh_generic_type of RETRYRAMREADLATENCY : constant is 2;
    attribute mti_svvh_generic_type of RETRYRAMWRITELATENCY : constant is 2;
    attribute mti_svvh_generic_type of TLRAMREADLATENCY : constant is 2;
    attribute mti_svvh_generic_type of TLRAMWRITELATENCY : constant is 2;
    attribute mti_svvh_generic_type of TXTSNFTS : constant is 2;
    attribute mti_svvh_generic_type of TXTSNFTSCOMCLK : constant is 2;
    attribute mti_svvh_generic_type of XPMAXPAYLOAD : constant is 2;
end PCIE_EP;
