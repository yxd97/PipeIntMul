`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UcPnACFcqLzxhaX6EPMRaDuCuYoNjE8aXJ/qY+ksqUi2i78qEl+ejET1TVViZbXn
NHqnof/nhQ2sfhbupTtR3MXO5UBk2nPjTlLgueeSAGq5gs1LUrOqDfrrc1zUpvFa
QwcAY6n6x8AqJZmUdkV9tke7V9IpGJGFs+XW6EWHEQ9ykunPLVWuQwkAU+esFd4I
/PnjvNVdzdOQxYbF49xc7vkHkfIQkq3kzSqLgRtEUAWzz9DcqzuA8tIQtNjpAa1S
1a2aO2ez1cJbcacp1fUuRA==
`protect END_PROTECTED
