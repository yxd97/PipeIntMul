`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X8vUjW7i0k5QOk7UgRq4zqOjZOCIEfbSogIKgXL+I4mPySvHxeUUWrP8mY36WyV5
IUg0CnMH7G5Ed8p4sBXsCnaLQbL7mFw++WJ6RNdfiWcfKUP+PmTBAgToRzEOPNAb
oU8o0ytl3Yyd2Q0uEnCq13YQVX4FXh9mHO8T5Lzt1IgM3nO4pN1STl0fkwK03bPr
gAc9xzA9eOooFXeKUAvo7dxfiRrLlqPO5w3xKLOFhfnWEhslljvtEx1fdck9jN+Z
s0ANCKCBDfg/EA2FEoPLmFP1t4qyjmClzyQrkCiKp0TZbNMd9P8eXO75UMWdemRU
XfLCeDdEL11/YZkC+27rLq9JJ4Uv6DVSZw8Ha6tsFEyC/e6OiRzTY11MuFLORO15
SrLPX6Y0CTYLJQNiSo8VQSUZPM9Z6tfjWUH4BRE9Sr8=
`protect END_PROTECTED
