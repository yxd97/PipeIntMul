`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yxRO9d6CNkCDQhUi6FONVr3vPoh50IdK7IZT/K+cQJM/Dc/ohIcRxMHxMRTYFHCa
MOH1GpnOQ8QyWEF9+t+rycWHKQ82t5z8KEEorVJjqAQTz1dREMf8JYOvvLSCCVsu
VjdRSGJKt1Fm/X2t2abT8Wih4gY4qDyCzvpDMKDbzQtmYJCnKe0Y7CtK+HVQ+HwR
81aUX38ZpFkJm3fiX925KXX7ebxXwHm7WzYIstBGDxqNyNr22L+xYw6pVWCfpa8P
UJa6vgR7dE5YcTMPxpZBjx7Uynfy7yfmMemmILG+fTprVFXv3EZ+Gi/2KHi2USp4
vU40kA/v/n7tYAFf4Usb600yYimSCBZ9r3c1StKFsBevihKgZj2iYG/xbXx4sacs
O+8EGFjPm9uu0IpMr6TB3hCkWWPiwuD3NWShODUrDLa4Zp+4Mpux1iD3t1SU00SU
S5UWlCGk9AR0pVL8ThXb5PPb0HkZju6UIJ69G1yphl2IlauM4nIUfxEm+CgLrcIv
k8gsu++A9xpL1q7Siu0ftklWvKUpnD6efshx69E5UKh4s5qc35x9lxHGHiyZ7Atn
f6cjCmwowrEY/8yUQ9C5xLrJCFt+XkKvbzBto2aZ2VWLp8B8dBv5X/Xmgn1TIckL
uTCLVlfcRGzRqHIaNdRaMA==
`protect END_PROTECTED
