`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ieG7oYlFXMb0A1j30ke3qjaL/VhbDvdc6u1grr4AML9woh7GifpXoro68zZJJnP
OwVL7CByZ7CowLFrHOJz7OrPiuYPEsnB9HTQijypn91jeqZsgGEsllTe11lfd3Dw
AkeP5znYi+E6SLkBJK+ECEMGNu3zokQ4PngKxjUeU83MfLvaQDHcP2m+6ywpIM4P
6nH0UqdOng6UPtdy+Mqw5Bhrttu2ZHelxdNnQFiH0w0CCLgAF1LzgQrYXg91jqTh
coGOO1iy5ZBm2/7Eiw4GmijQq90MDjiM3ef6XZKZFj9/RzhMKh/Egsnj/Jy2EQJD
c6m2ds9nNO/aMCIWnPqi4ZOZ40KxCq74y49l0DPYSjSrL34y7FXWGxZcUyYSZIbI
hgnNPF8nHOQM6T46IEKulVQbd/gZ8SgcNvOVHUHALYEiHDd94W+4BMkidioDyDHS
UyvGg5qtp6Sax0nBeh8R0wm7K0ER/wzeaa3MLt1aLlCIvNv7ztf9Rz8Dnq9BZ6rm
7wk32UpOcoObN+xX9wfSlTyqSIzV0fnFp41QWfzsJ1enXq7K4/KP+or/dABhPP9x
q9V550xUxCCySB8Ky3UaXeXvlsiopcyCiwEGx2Hz7LkG5Hi6sR9bgD/buHVodONu
FsxZfyKYuEFnX/Z927yzvV3KGgnuOYl8gA+voo0ruQR4kA98iQ4iRTKo7Bkzd+Gu
1Y8seMPiB7C5cq8wL3QabevnC59K11tkABUoYP+1sGNtAYPwFNe+2u1yNXgrYbA5
i7QcOdpiRMfTBKc9NRCgWoKy0/o38jIqVjrQkCV8c38tGONcGFz68C3sxO8Pf5Df
+TNfi7nqOPp/sIA/Yb5T50A8JC/bMjQIbPOIRnl8pIV6N7xQMxTzt9c4TBEU3WPO
grE3W8co2KFzP/U4H9mvzOeXtVKyXSriZSYgX5dNe+PYOx1mymvfWbcemJ6bg/Nc
GN01OlobPfJtjxYw1b16mPlLe1mnKKj2wwcpwdZ4qwLe/ZWXHc7spya4cDEkvIIQ
6NPY+GkGcR4yn9Nxr+cs6FtNC0L+dyw889Q0JWh7NGbU57qm86HLXXjMyBpAE/P+
nLr1Kt22U+oSJjtLu0WMdNwS6GJZb9uZ3CKp9rMqWLSRGt0jS1hkwVgsvLywQk+L
3T3H8MyOsd7sthvm8lC1zARj9Ebxfceo5Pma+0ljOC/+nbwDG6kIkCUktBtxM45s
UKf/zDBY07JwAHMuV3xYOoWReiINjrf/yhHt+yWkBnwK1yCi5aDsaadlgHe4Qinz
`protect END_PROTECTED
