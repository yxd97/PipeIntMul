`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TmJxnW5RgH+RUdmPXXkuNbNUTUj59IzDLmUVesia3rs0Z9czxrqJqd51VlRzYDwh
Wmqq8s8KW3Y6IvELenUxt+CA++QTjNnkyJJ8Wj/D6g5NKTKQjcGocltKkFNkzuWp
RUO4itrI3fXSOITyO5bApkokDsdR3hHk4DHECKJ3dc5Jrp9TOPs3bDTDu3BYGWEN
JCNTAV1OlasC8DwU4W9YSVhPKenlQz4yFhQ1UD7v7UAtFAu3A75mKraifrVgCM2i
lRhIH7JN3aesxu8/C6uGFw==
`protect END_PROTECTED
