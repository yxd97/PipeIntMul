`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bq+gzCoXU3l4j224eRc6B3qrD7KFqkeT09TWmXNQwvsdUmc3z+I+GwJRlmnMD9dU
mFIj2HSiamCksnQ4foyPtIoRjxGzTtqVxq5KMUx6sjRzvln/h7x2tydZlhGxTzk6
aDGvG1CZOlnMEqImwhBFPuT+Ku3jB/Won8SQFkh0mu5ryHTDnrpv//Tr2ogjKUFc
ybpfKWkSOY/My28xLcR/R4fzJav7LAtmISqkA5QMXhpk6vs9qVc/IRWpkYJvmU+a
oekPGwkdRun0DPSpos7eFcS1ViWOH2/cQOOXPh2Om9nnP/nW6PJ6h1N9Ep6285ZO
5bQxCrKHNDiJmSSi2pBZguJ0YD3peLVEjctN4YA8dntzBoR0Q2Zefy671dWnGWvD
At2oVTujYzpxC0c2uBOmzWG7LPEHs0P2ntOMMAUxUPHLG0my0ydTgxlTxV+T84Rp
1owI1z+cXjeco44nkiG4xY7yg2gg7dxY5gBT0QD0moVDO6ZhHT4C/9mfehlHxXac
XFt64MPCFH0rG5+4dzPR/Fwiwajvbnb0RsQu2zWUYcOLYDsoCKWX3TrHUA2thq4k
nTedcJSlmkROe6pcJ+BcSdClffUCnW02HS23iJzE7AbqlyOLCjAAXf6wxCr1MAYk
vxo1SeT+1/CeaPwBpQVMpcQcHbBIfZvnn9f/aTBv4gga2lQA5KPu7KAH2UEhVMTq
r35ES/hdAh94mrTMHHf1MT9Z3JZJcj/5v565dnOsttb+9GCXL+iGLhraU8oftCIM
IlpYpX9bn8fH2KfVfuNnpqrMkJmPKgBYiKqR2HCR6DxqrbaTtgtQSfXlp6VaRMQl
9pO7U8FufcMnTcjPzbKDqYm+MmnA6zX6kufF3NUCUhv9zc/27BnycWcKSEPAjnx7
o3o+JRHBqjqlhkz7OyC7S189UEB3DYRM5wAwgvyGL4P5fvTlWWuY7VPinPLorLWZ
bHlTTdMdbet3+3TnGtLurCTwYJ2wV4xczviXOuzEcTCOxBOOnMUrb09uTBC+3xRW
vkV91s/7xtAUhUZqW/bUgCZdTR3P4qs57GH2S1oBpTMwQWoI6aqcvtSbIq9xIRX7
dDVPUTixR+/lydhL+Cjq/lHZeOCTo8QyG4Es9CldRv5yZZiFwDkJwxzKCz9VtNj5
+kxRUSa01/GBhboi6mr4BNLkhzVApkHKd0VO0p7uwPM77kdJaRvCkc4sT6x1wGf/
THgqnZwcq5GAiWF4OaB1ijePhGaE7sVoDbmW9F2cU+IHAMMTWVpACDEWRHkQWb+Z
QjHPD/a7kmZ+na1cFBBSeFh6mn0CiHWwQUE1lUDeQ/0urpgj0hn6JqcLoYaiyCva
9NFVec3M2oOaovyBzbAer4epGA11P6vwQKfSkS8UV4l+rxEccFkN8fXttTb9ywHK
RsyLtqvr8Zlw7gFwUWAcQ456Ci+8auE8UyDU/MrpTK0oVnO7XzRfVGOhL++m8Rsz
2XOeetocXttqSl3J+pRAN4PQb69kpdkDPIeipi5HBN58ys8GTXE+gVEM8H4IOxbP
aOgDP5YAZUzqW23sNw8kTopgLQMo2aYmJQjhhAKXDmYJh2xMNmj7az7QiqgPfw5J
+vZxT5iQMHppR/sbGdSKwVDJO7LqFYJQdFAbJIQH7Ya6MOm+O66Y8SCm4gdNUHM/
OPnWnBIv18H1WFX0jXPnFfmza++8xmJcP2AX5ZFepHWmOh6KcSyGt3r1OICHkf4Z
uDRinHUop18Qgvx8jpemryh4IE6MiizuGCwCdVpFJMRsM33GeYgyff2ndROoNWvS
3bwfwnXBSSTsHEcD0gWjXlpJDx0F7AFk89jR0UtEuHcJgKdKNvJOSGLLdPOMWWTd
Fk68dw8bRhpatT9G4sYzPgtH2kCllnIkaIYxGf3yVhX5LMeueb3QsCzTQwjkHOKh
SCYtfYDxn45pMv6CssfX3IG/rCKaVLNnj7Hd3NOQ3PnhNTCSo2u9MUQQMpNiGn4n
nblI/wqfdsyHxvovmeubj8aNd849Fzz8YZgiAXWNb8aSgW/pmwsSDsR5DP3yxfVW
kbjmAr05Ijo5vm9nrWZwXIzR/iokq/2+Mdlcp/aig9vpo3ZrOrvEeMfnvJLgQn+L
TST1tAB7UFM8ZDYOzsmlGUhDVITksXJJx0yU16iFoCPq9/aqsuGZ90rRETgb8k/A
ZPlxWoGsBvSLAK0tM1eBl6OSYpeQt4vXzZHqceJg13c0d7LH5pFElrAfZkGHATv9
D7lInt/oBSo2KsATTaYA3/O4n2ZWmY6ItAmsNuHUxB97d2aHA+gXfiSgwjypISCv
4BiCy9YlhPssz8jyGeFy+4Ox4XssnXQ4dq9JqrlyIsRq0xTe7apj9gnFX5GppU2N
Lv1SgeobK+5ciyDRuxW8n6Vih/V8Fr/OgTvWvqpWuN/ccQMXVk64872KRnwja3lp
04WJLMsKagwYGboM7IFgelYLqhhZ6MEehTdahLXrnYtG13z2S+jSYek/sudH1pz1
r+MLRaUVj2HbAIeISZ52XgtLfIf4MFcUxA1lPlnj0d9R7MWMmUBjJG47dz87Agym
wnxqBHTi38A8xMHmbLT/kwTGicokBn5l9JT7RtxRmteY9hiuUF0IALjWXdshP42e
wRDaBxMd7rbGuUa4ZRq0OKmoJBcCMaLna/ChEGLuMRMEz2X4AmbIDqmOP0trqPwk
e9pmRvQ+w9vt182D1YNA0/nCk94Kk3Ol0tlM2fZVD98Q3jhGW5ElLE3TjRmmVWmb
M4neOyqGMIVBQmlEZ3WEn3HCPHj31IrISFvnfUvZ2N7GcPOJjXKTA12D729V5Y8t
baFRbhBu4NZlEvWFxh+002z4QAkA87lJjguU7wyHmo1414WzTC0SSNY0u2nl3dl7
JqjPvpChBQ1T/48I7dOjKOGE9w0jpMINnDypKlMPy3Om5Ca5FTPsiYYAD7Fk3NZO
SNlYJKLff3nJjpOt1qVVdiFB1iFPCO4yowHXLqfVymGCNLqSW+LunMVveUgR69vc
S6j8OnrBFYvNZK9LfUrtihByuwpqjgkXGQsH1KOeoAxzXmJaQkDMbTb7gIDzg+3y
3fkl8gMs7GFO4h8VBxsylWFY0/eU6N2SWOjuE/vUF3Ag0NPtAcxl3KEObmqhB/lg
VTR1hqzzcsfXh4VMIfuOw/M8I7zYNKLiFJEwxQvXyP5SJdM8s+0ML1kdalcOWRAj
8p8DFax90xC7FcNNeMkoScWTRU/W9IA/seZV+dcJOK/Oqx9yJQ6CcIOghP9U2cGO
K7+rk7USdvAvZHFjMryqsJXQ/874u9Agww/eXnwOVDa55HNjv3Zi0Fe1AM40NzR6
m5v92tWWq8/zPCvs/jv7cGsbWPAoIIgbZ2jbvCnUZ5kQ0IKa+28Sfru2cnpB4QlW
y3GXgftcNRGN/i3nbS62aOiaxfgtJc2G4IpOYX971y1ykWaXbkUzVzFqKM0QRQjR
h7D1GvoYU9Bl38HHD1/CZfTfLzOljvwlerqqOiNU6HfNySc1ecCyco/V7+xdIuRj
WaMVbGyeWqliLwLe4Dt5+JZi+RmSJmpsGU5F3qeXI5J+ka/K1ykc+egHOdBPuWca
I2wV1PAJYVN+XdAf3KEmowR8UDc8SUlTQ0V41Yviho0SFMJYS8vDNW1Uzk1va8ja
oxwwPDpIoCgLqG31ILmO1/CH9RKY+rjh3fsXLEgIg2gl1Uj1CwYBJub/iua1E0Q8
CthDZjBqjD9qBmYDJWhp7nlIkhT23hWJLlS0kqxAXxSsjmen0JshQ8x2Ba2Zmr21
FbZi/IXRWBktOqNZ0ODsmqhhu6fAjSz6mru8H72VnfVInmGbKL72Ima7qrOe4tZN
4e2lBEVH7jo03x3fnhOeApv9av09TQ1dUKT1+5pUT1VXH3CIkxh56yJWqSRd3t1M
FB5U7viojY/wrVtxHQ08dY5YW3R0nYFlcGKKnFi31g6mizR5VUsyC4IE6e5eHUr1
dd4ltoGpadulPaz7Gqw5N9aUWryVGFmNTH5SoOn7GaQ678Xkamqb031knNLsjTT1
u1jJNTLM2/L06sTI9h9Kq1i1VgLJ5pDQrStJpkxkLHxmErhgEsSMFfd85WDcm1NG
KrsStCUWqYJ7cS5u2PVoqPZsXSYgxww6Z2oxyUhXQoT9mgsvqyVnEnyNJTQRyOiI
lP2fd41kaAw7MbXhd6YIJzw3SzdOHg8rR8xMFlDCE1VmmnpZPcyCw3KMsqBtHjRE
u38uefg/hx8DKaacNCS20nb1ResPT8MGEtJ3BFnHnh7i04bhpHyovN/YbrSQ2Lfr
I9VOCbkvG2VATgeTv39Jtpfb1DVZ0ZftufQ34gpj2CvcjH4NzuvephcrMDE2BMmv
hDnHnF6hR1G1tQMfT+MURuMsGv2nWB87SmLEaUiDnEozelHDSJaUHCUyqka4tFJ6
w31m9/JjKrjqwogXbKYiod52aOhBKPl4RicQ2SORhUw1H/fBG3yDFrcaxy6GfP3a
xOhbS/9jmNinlJ60uPzoLtCg/sP2YoeII93AXtCuwK0dqmHHwz2jGL/qVtCQcGEF
8C4b1JoMVudXxPRxB1PcVzwq2pxxnGRoA5gEGc1ICSeTA5WAyJmxH7aKSTgFgoPK
AS+Fp8cDw5C5sKWsK2HmMpIqdMHy+MY6VSWIAXN8abkB48Zkls3qGBjOj4mLgV88
qhBilzqFg5mlPdmMpNorctG7kNTkJfxKqrl6iym2g2585ygvFzwfVeVtbq1GOtqi
YBHClB5Q4ngJ0cLn/lLG5v5AO0RigzDGmzI42f2ZuLvAa6omeN21YJ5MEoc/h5P5
rp89kwCyJLKeBGhAVPV04Mw2Q+M9IbnsaeX+ZUqWV9yRcglMkJoGBf3L0WD+A2us
fTaRJW91NpaOqQiNbNl++bp4tWOp3xEqO9rF8bizmqbeTahPvK4kaII6PJ4Pdb/c
iD7WruGnxJRXDud55zVOCNHzJCiEZopFsZJo0KpFuw52gDZClaqwKu/MpUK7y0O/
kdpDZboLwOtJO2djgBtjC1tIF9kutQm0HbAlIs5Xq9Foya+N3XulAk5BDVfx6IBv
QEI8/Ej9JZibPGzbXBG319L7yoSgz2BJpZjgRopkopw0EEQd1oOa98rTKzC2+6d3
VQcm1EARECyfs9SHEIcDYjcVfgKMqrScKhyjcyROftoTFFN6dxjzZ7VgFq0CY8vA
qe/hYhEFPmPf1ln33qccwUCdZfI5GBlluGVn8Ej8Bid3jjaNj8LmXgCfkUDGDW/5
71UdD2L7CPeGw6YlAFZUe32Lq0L0Y90XGc/kYhOkHFMvX2kU/LiGEeQmp0MKV7tx
hGoqfNkBVb04Cb7YCQYFjnPfTz/Q9JIVSxP/kDC/gfFwokOXD9fa8vjFanbC/wPK
VjVmN1e6FsF2Ys6J9YyAcSl6wEaae4YfeMCaSWMhEu0r/Aa5DpYIgSJK8iIomUUZ
c5uPDg4/CKftKHdp1t+d8fwiiROk4XWLRrhsWYxkxRDgtpN+MvLadwi/Dzse/1Q0
GKaOzt68AAsHn7St8eiNjxbTGsjxW8fJdjZCLL/H2TwkFpihmNd1+iVa5UosHvt2
InyX3vyPZjwTGyVOBEy+r/HkkUj0Iqs7YaEGjx2KJh2rC5PavM3IlRGtxlLFpgOz
wV3H0jJ66Q9dYTFiz7itJohbfefya/8ULliVqyDrs0ZhYr9YafLnmdmf2XeRJAdE
FoI2fx9M6necatsJtpQXXWRGICyxe7qr9q+LJt9C0IcUtMuGrxGyayWZeKrN9BK8
trK0XQQNGBy1tPxizxTjgKQhsoQ+yKSmiwZ95Hx9XSACbWHtFEox+5BPxFbbIYR6
jK8Y9piRUWGgLu23dgMshcvdn37yCw4irgEEOFQjs4gz1PF/4sgDRPx2Y4SmcVIY
jkWp1Bxvzsk9VrZA12+OtoJZlqeNRor3i/CVTIwafTIb6suvyGckuuxr1eUP4PXg
CyePf7fpxt0QnOUBvooWLZOsgb3cJqvdhpMbW8IAT/QQNApSYgMBIG4RJy6b55CN
XeLC8HfCf6mAxwYBgH2dXUQ6ikMphOYVS7aK5NTYDAwyNwFYrRCaPdvrCzT2np3n
rACqqr8Q3FMRpB6vzVsgsBMdonNP9IMog3ZjrHYiwa0qkG5eEbekBz/TSzNKUOOt
hbVXvyeJh8pIcAZRCbdocUe9y1o1Bs1otMaFAbPva6TCXVnATeoDXk+yjiZ1AfDg
skb9wAESigP28Kl0l4nmQ1wIKVb0+EYMGz2vHwC7rVV2ragXkTp1dnd9VCNfYXPt
OjvGCXSKukEXaK4YHS4Cn1xtA4q2yNEfDPktldxTe1nF2s4dztDdJJF8cHp+njpH
8qzp4+lsw9gGmdQcxe+wHTUnKi0Mc/fJG1xnWiXT5nS/rdomx5e26ZXXxVyc2x7J
RjtAnBFfygFiJP2lt2kHbKE9/0RB5QdfqChWGofDOvViK1h8BnLawTFXo/OLDDHd
5enIpBhyhwDDQSywbhXdj+bmMhi7hNRMh+oWSBv9SIdi+IqxBKdjcDr5ivECZFs1
4D9wQ9DQCuWQjKKXTXZZwzLuiTLlwibFcT3ZXBEHQPer0zGlYfdD+dIwzMKm4khT
JzMeP4TsNlXnAP4Ig//147GHaG8qT2mhjTZi/OxroXf/WAkEc2JYbs8rWZ6GAwKU
orW7D9KZY+/WzkLWDnZ5bPSCcB7As6R5X6VE3IQWktAizV4tynAOe9TJ7vHsO19N
EyHYTUus91R2uccrO9F+jYbYdRN9u0JFwalCoWSh66IPwYyF7ZS8t32waHbNAzxQ
55skjBVbCbCCXwy3xxsH9nn1B7TUFIk7aS9W84RQ6Q1lpKLvx3cz+tL0snXyFzXl
dmrzindaITiJHr6xstPZHQDf3i5+8Vwysu6khkbVK+F/KD89QdnB6s4V02lsyFIR
1npMPKnOGwBznzqRDujCAlqYuPuw6fl5p6eo/toowj4mq7kVumYfjsOzf7buRk0m
/VJOSEoSYbO7YrpOXCl5Iy2YDUJicJXzIH5uOgzBIb8+PEsbUDCxJeuTLtg99GoT
5+jY1aedncQ/E3FzUo0fj4eA1kdRHQaeDc9fN5oZmlgONi9heHH1TfiH1r7J3hl2
Lru2O2HY6Q6KS/A+5d46lDNY+jOs7ioifBmlqflmHIa47RKFkY7eb43Ty0f6OaX9
ORyMVaaPI6N37aVNq5BdMbQI229wRPOHqHMJTH8fv9n2vB+ibngAdb8ILysnh4AA
AtIWG8sL0715wvYjxcoRTjmL0WgrfioQNl4OVzosUKI2HY7zBeNFxmjo2ohSU2OG
XpJYWVxkglqvs4tkmXUIi3JeVJ9F6ziEA9BCU4b3z/A2Xnillq18GwpvUD0AHjnD
BLjnt0CIKl2eTNnQoPxLGthvpo+LAkJF451zXJroZ1JS0hf3FzE6faWpXTiClZC+
IH9UwguirTHUlbONn/zfV7CDyDkklnOPejPV2KihoRZQEjeZX9xOCYH522q1VquI
hsjZdd0QvRmWK8TrLsXrGxamUQqSN3L1pQ4HRrdhn9bfYtwDKPPePjspBNhP448/
ED9Vst0cLLk473ZHGH6sTGkY2oTX0cG6lh58C/1BAduTKRAP95dv0gdrAkYMCH0G
2kZbRPk+VI06yFTMcHJSTMgxOgovuHF6HPDFjQ49yRpbiIkKJXhpmTmtkXXqvuNr
pFq1mS8WABE81i4rhlPEZNB5QSt0455zNXvsau20ws9dRtEN9MiEQoSSxXI5bmSR
GT+Y02rlq6nxLFtvCDbyGn58KWzAaZijcRNVlaZbIAqglQfBGog9huWxjvw8K4gK
0wP+r2LhbZ7LHlix0LYGTsLdPyGT5PqRZetOI5i474ICKfFyqKMBjbnkPnQAs4Zl
Pv2gps9itOXrrnUwjZQ1HgXw5H0M+EmzlVZdebxBcqrKA0YOk2cVRjcMAPyaq070
P/5z4+7Q3hkF0ZM9sGzipW2OQXDUgeAPCyds4b+qj6yXmo5uWX+xpeHBazisnOXC
ANtrzEJ/lcNj8kRkbtfhmtTBEY3B5CMRibmxpzCKSQuyvkM8oKOpmmBhZ05Yb5oG
VDZZtBGpAhmTEUgnk7melUbXp4bBaG+wpTfhLEPP9bHhgKXwLSyFSXqx8VT3vkDk
0tVU2BHvIjE2wWKNEkiJbzso6U6l15Mf8zACX0yeAO+2jppclTfL6paGBCYUMvi4
LttMaxR7pyQQ/bPq5MoyPKhZ3WjTWnwW6fp+gQ6evhIbSLqwGBSfIoIfWHo+uHO1
vzi1hiz5lz/ho559ivK44TtqXoHTflesGbgQwqJgKVdazbhuWdGrZgwCfnLfH5Hc
9iqVbpn4ScwokcX64PLqyb1zqpDGsIJmbj6mRe9Kh3Goyurg8qrrNtV3aGvuqG8i
TSiijyw6MUtyeRGUVRFnHGi5fZvuDtCjJVa1xsfsOVjGoRnZNAR9RViErhRm/RJS
Ar/2Z9uNuBTfcaCdtDWJwHm148j2wdz9v9oheJh8lLTq8PYXz7XlEhfr4QQ3itjM
4Ge42RqAl76/NleiKxBql420hLpGAQ5S0Z6Btq1z7PFXg4o5csmu+Fiw1AWZYnAF
15DViTL58kC5QaidwDvemsTH7RVn7Iz6AnXivxg4PIq1B7TDy8OLIAyCJGDPzPsZ
Auw5gxXZIIp4VGLmM3u80SEm9matV00O/KRndKRfqhnxhAmw28zi+jlWaP5s2Cx5
zw/mRFwpah79Sd9vQOtTNzncX8PiyKdp3wAhzKGB/Aod9wdRIRsnTISUx74A62Wu
LoT5vKnuBPkRu2829DAPkWxLU7pxcgDYwe+o3V5LSJjwFn1cTBfEcOwW8NvuksBx
vX7zeTN76qmA7QhcFQ+QclSP2tKeY0oVQDTPOJCL7tzH7Hmnu8SL/VQNfSyHK3Wl
i5HSCMJRlT54K/E4XumEKgfkNwVE6TVcqp5RDFA1KSi8LU20yzmdHRjZdH6o8/Pv
QtwGBLiyxBFai21lCgL/sCuVDXxrtP38pM3WHAte1PrSxnUqnA6q3kSYlRCzI15C
KEQGuS04xd2gG6huRrf1Pp9A661wiClKiVWDdpaGzDArvA9iWZ9tEx+U17XTzzSz
z2T9cdnC/0qDzj3REaWfK9VPjchXPeoVC+TGwRKBq0lW6ljjXD4kuyDjgArxoSdC
++y4R2SR6IMQxyJbo7o2UHWriPR7k2XrWNuf0GRg0CMmFVO/V1wCWwFUq8DO+vZC
p/D10KZDNn/JlYFU6pB1Ufwbd39zTLDF2Puey2oKlmNZTp3auyPkxyoEu+H6dq2q
T2v+ciH4rllsNZgbRHDEK6422kFXyxoHMZrslwi26Hspmpd25mfiIUjj1lOLhqHm
luDbvQRSv1GBa0TsqDQHZIeCED/dnmVEuuNgoaDlY+xnBiIciEG2fe3H3Cweyrtd
OIzMyBOtzcsM9/B/Z0tGyj0GIQz/YPcHy3xUCudtryoN3sIvK9obtasg2BloWf4i
Xc+ptkt+c+q7FK9z+RGHmyAA1Qq3sMVi/ddZLiJtwvKKD9JW/6Nc60nbNtt6g5oZ
0IHd2Ef8l8bC+nkm3o7rRMIpSvcS3XHahME4EPXUwyrECChfY3afoQyQSHYMIRaa
hECTMpdlZKgaf/e08WlEUYj3Qstqm17APKe6spIpNZJFLfgH8qH+3u6xK5Zx3A8z
5msKH3NkzvFTRjiVeY/3L18XBpGBbgdCEk6l2AYkEt6tua0CYgGYo2cfmCev12H8
q24J8R4Spqx6tGju0pR1Fj53njNQ0gdkxb2Rexdaz3orUmHzfWSOYWPE85IR3rbx
ih0qs39v7yd3vaXMzQlHhXGfdbB2jaNA+bc3eng/DRw+5I28NAwS139KP5ju4W6/
4x5GGFJVzPx4mWm3JNyelhTwRKB3kv33Q9Jlg0WSqWaspI5Geh9vnmbwGxQCH5Xp
qviaW6vJ5IDoe8lURGcf8WnRWje8kHu1qV/rpQxcFO1kTTgxguvWhTDd0FUIs+C/
Fs+0MY8BExOaLkfS7dB74nvHPOCe3Nm014wlkEjWob24isLFpqF+iyq/4hx0tQ/e
sWTsz67MWeigiWrSFiFutqqLmzTPh99u+4XFVfydg+yqAIBOKpzymxoE4HUttA8d
22ygrFmJKJMRs70WiXYDRkB9aH52BOXClQi+oenR4guBrHHaAHwzdeCaeuVKXUDz
onhs7duZAbKgppojDZxLmSvVfOpQStFNpGVZ3Rn7BSIMmdaTREpoF57OAKtpd66Q
5dEw2jen6SAM+DRyUgfjfmyJK2WpMyEvj8kClE457fvKAopVi16z4cuSgMUt0oX0
fscn89ZIid6Iyx2p0ym05QidLALM4h17WxOIDHsnmf0TgjKqa/tQCLBnm9iyrqh5
DSluEUVRoV1WUR+ybTgId3/dvCACZm7tpCJUFpJKXIeuaolCdzvd07MWBQaqaXj8
r3eosS0ucI7XxDqPWStRSrK8EoVnLL5hAGsfWAgmxuLBUKumLHyoQEXsNq6bbBZh
HMnBM70mYoUjAU7YehBL+HFK++N2XaVH2bNfoisjo8SUS8epEogqEk4qikEWSmlv
ZbfSJh1W/G5AUN38ZMbse7yAGpTia0na0TWY/0FK3a9S31e++hnofYeDmOSVMjpB
iYTTpiOPONecNp2Jqepf1T3CZFKEEV92rYcdcwu134dupsBCIY2NwiFzXTALRlwm
hhXeLuoUPQqdGb4s9AqaCaVp29020EnhZ2KzmFokLLW7b7/qzCFJf00NmXgNbX56
NMY2tvlXpIl8vJ9P6/yNfo9W/9HNd2SyddzH3KvqUmlaNlgHnqQx5IUqnRUkt6Ag
n6wIdp9ufCrSsJOckkJEMimNDefctlgYKVJnp1JW663Dn2VXmJdAqOfldXzpE3zT
m+NmDFx+Hlblvd9ORd5J72kFgFe6gVSLVGloekH6T1yXN4Dnw63K4C96477TfjwT
t2ln/dnbq27UGYyLky//eUsg1HjU4XKEsF48nxzs8Anqp0CBM/qWHpQAlM+IBeJD
3vL1toEAmWvls2EHwPuAac/i5P9KrZXDTuNIU+6lWbl/T0TzGSZ9AP+1cQolPRsv
7kw/IOz48kir/+MyxtpEUs4atJXpS1l71mALbD7sqfgAbayMcyynOyaiX5cMJ8fr
O7ySH/WGkNdDic8GhRaobIPfg7OELv6QXFDbn94K1ReJriG4km0GwBde60p6nQu8
DqjULqKkgH3Sv9HYjREuxhbibKWw6XqGXczhfHh0NdTLgd4ZKbBQM6rCubF2tWe9
c/LCdkn4komVEGkc2ppf5IPGWIGXJD7lVzXgL0D8SQ0MvhgZgoQdNj6pVXDIDPDM
8/A9bOR/Bk7XcR6MPawE7lHBmAeqHpyZ6H+rpCF1ueRjDLSgFtMedtC9+AAjISdC
cdXlO8bQjO6lXoJwI3mjXp6F9VHJKA5R2PyFeNEIEvtcqhdC7MQmT5RkGfFOVZ0W
2CXGFgW5rOanv20u/Fv3sR6FsVzlE8NI1n7fzrdEBrRWKgeskZ9LtURJPeZqb/pO
JARBhMCN7wBHcvkMwMWbbuCo0YauFY2E7IldA5eiZPXTWlPKJu0gcvkE/KIpOv/x
ljJPwrD11EQ7Sqnm2BIikFZdb4HEFj0/Y9aGKCp/RIwjmNq3D/rN6PWtle2SrLfg
OIwhTIxRw49bFR3G1fWIK/E8U4oPd4Zb4IR26nc+m3C5Pdu4AH77OL4D5n7ShpQY
fptajdQ7VJ41cD++OQ8dxIiUkD3a/PwuGwKJkYNJ+4GS3hv7VrVFA45/Pauotds+
iYrSaMt2ZyB9ARJd65HbntVLe5bZyOOn8bYgttvb1oICesqXSEi53hML1Q/mpVbK
a+hEBA08s7FEAX3ejlqE1gfdX8VYqvtgP90sd/kssRzJc/AOvDFkhKRWvJMOJjum
B8Uifvrcg39cLm/J4zMzCcyPAwg3/aEWNrzFAxBr8ZcQd9ZEvx+zzGY9YUgXUCYt
ptZMv838gHvSMcKUg1RCeREsu4cx1SYWux7+wsABFMep1IKVNG7vJr+SPf89Hf4M
YbejxLs6eSlUL/l8zYmnkPwCU4nPQtInFVzjKs8ok3EDQPWWT/PLr8TLGwX+i//i
xGoDVu0Tr2Zrlzy4v7oy2EISv65gfJYSVb1p4xS0iN1xWb5rYr29yT28sDJO1LMv
/3YnvikPEYG4QtFsVSYnVtGvEkEz+H41jL1aCOYwOx8glGZasEG6Dts9k7/8DHDR
dogtZ7ZVt1+5BCR4YyNFn+Io113RalVCpBmThMLW2pQ87gG9qQ8gN8zyry5bNk5U
KPJIzZDdJ/rC3AmxfaxC4P3PYWsrKOja2eh8YdxeMU7tpdOfJQR/qEW0Fi4XdfNL
oetBRsOa0HiSEu1geY0tFjDjeFQva5CBxRNphKfMB+KbHbIAf2pBLf9OtS/Dw4uk
amvu4AlakmahVOk8Mz5Z4xipV4W6DYVOKtdu+rwCfCNEDC/cOhK6hBNi2yyVn/ne
9sYhQWk8vLKKPqfMCM+YjrXD26j62dsYyQ6OGmH5yhkOuvke0U0C8sjBBHM38BIS
/fTREm7/29MhvjYtr0YFs1QEeA0SmTl4llBc3Zr3R1Yi7yRcBMVShETavU6rlqOZ
K/o734VvpdMrRWtBaZpHly70IRPSgX95eXUrhhobdLLZgiLFKLrgscD+FYVPgzcG
G76rLSfmBoDL5i8RzZZ+1HaL0H+p4EklSgUPzUS7xYPZNbeHrwymrNTmXy/rhkUz
UkpJE1kSdZVWIRlG0QAN0hH1NZPGdiD54oz68Q5AiVLPtYSdIcFxoqfxVMy7HBKz
vDNR14Vf45mGAPT8+BUVbehFvkG1AK2N1hBvQv4ADcbWeuSOgORbA6l3yt8ONrqw
PknECptuwY9C0hUhNId3WPYkF8Me1bV4shEVGZcXhl9dGQCGokFvqrKDnXn/vDcO
iuSxRTO+4xkWEK3V5O/HA3okVGJg1NwLLDTVL8EhwTmPYtd5rk4bmnrHCA3pSrVO
REOTK+2vZSpT2sDX4tzcVkoafkLUwQauQILYegfkmAnizz94N1lR9tvABDJmQ0Bx
M8a+VmckY3oz3jV+0JY1DktazUIJlJpTG8DrLQnD7HhZdm5GuDq2lb8bF4w8E4Aq
vhl5+C14YUtH9VKNqAu06AbE1r+k0kTZQG2CN2f6fo+gyfgU9Sr4lfNKeJx/DCEo
GImBESVNWUOWWg7js2+skAXNzazrqSqVyaFSa9ivI74n9zAbg3trBlxLZnDaPv+m
zET/JgZY0xnYjqnHPibRezxKg97ZO0BHHPA0ZyLRdNUdQnNBrzSSdWADMZF/OYEi
5VSZG1hj4hrKGl36YGrjgdJx2XKlOQ+5tbyw7r055eH0rF9iI3+5DkRBpsMRePNB
jhecnvZD1Rwi8r3hOzQB4zwOp3XmgWWc0eftloL6asiDkmdLenD6LYVlvaall0Z2
m+PCQvbwgrEppHGoJcNuvwh6UT0TG0aZd6WBLjYif6SqLKzr4cpEE7p73vlwzBPg
ES1d2jzfETwpd8EpQ2vd7vCYztmab3bw0AYmeu2wSIlDUVlgUjMk3NC9KSBRo49f
QZ6AQGRRleayOrLvw9ISL2eeyXE4fCgKLY+qSExj6mIqAsYqM9s096PzgzY0Vsdc
/PQTiDS0aXUll3/xwKFJawWZf4HJXIb4ZCtTmIQp6SuJsz/tavjN9tqVcHlZZt+C
Wxfw+m2n+D+4IaZkSxOYgk0RfH3IIWwQjK5IB6OloGnKwoDs/+l/PD1VYwdEwjwK
0tBcB7zRO9GL9fPGxbTrsQxLuLIchL1InK3/RwMmfMWFxQwxEi0lJyzz7JQyYs05
fham8Bb93Ere5goddjv3T9hYKC6bqUUBe2BrIuleaSkmoCAH/PCF/HlbAGbqkXd3
nUdYfQ2Sj9DAOZ/f/QMBhtFfOs9Fckpl69MO0FfCuE1LscpYfFHXICjkza4PEeVg
Z+OugVdQlzcFsyNyPlI4C7V/xeAek0QGdKAAmc1DT4AiqgyRTCzm5KsKrKFsFFLW
b9/bRgWrbf5h5ND9ev5jZUD4f3V7Z2jRGETKNLZJ+s1v0Q9unNbAoOiYgxmqXlbl
osJxwVWQ0AOD2a308zcMAohjZMoz8vFtVk7CRRFaopc1cWdPwVBmd4YqjGDKFnuB
WYRNF2bt2Dg4luacdg8sZmU8JtwEfGTRKcQEg1GlUjb4/kWXeKvpgAAvqzC+1NL/
/99Tqd8iRLi03n8mk66frfYEK1BSpNVGp4YdLDvXgVu+RVZowezex9nZ7kTUtjv3
OLZqejXxXdthi2+iPfykrZ1taVb82Jh7gaTTDF9atrUuiF/IKpEVOXwg4IdPz0UJ
nFPfo4cjNyuo8IEpNa6GKn6ng0RKjrW/O8jDarKm5qZZGYIeqXAvatUgmIy5tP86
iREipBlhwWUdcNCAJEghwAGXbny5jqtS1r9qXFWO0XI2dx33IReHNrDA0BQLeqOx
unqxMC6uQNHi40tlpjx3a4XYsS13LGURn1lIKdKlGGbvHM35OIQDZUDecLhAG/xX
4hhBYIa1LMciL5vGORn2kAibrXYPSgwbD8zEALjOhnLlqqLRqC6mpcIjrd5ErQSh
8sFgNuYp3eB0HP/xKdQwyzwnlMw/Q90xA8zRR5l75dZLNedUfWp5Vy7nXiEDQ1aY
KLDe13bnjGFKUOpSpq82VcHCiv9Nl8EheWUN3ldwTUv9TwDVXTWqPC5+A0zC07r4
5+4gOmoov3OGWo/W2MUiX1kvk1j3maykilKkNTceH5Vs+zou64Kw4j9R60ykbAGm
FrYKfu/09pdDODVWL86ipsxKmYI9I8ROcNg+VGB5+4YXhHVacHphOY051Y52yvpW
C0VGJ1kNNGZ7Yis/Z5p+kpvXiKHE/oJIHJuCw0YpGyNWjltvpCnHgzKrGdUlia6/
s5SxUu0gHG0ksugGA2ONdQwAIoUeYwu789OkPQPUE7VGnEY68MgxEl3q8mKRn+zg
rbruIeo0K4MW/wkovpTNA6u3r776qgpX+HKrXX/HtzE6RN9jY2uPN0KzgqOCkl0/
Vpy8Q7155FOBdcT0gNQ+be7Rs9BBWzb/LJh2JvbgCXPWVg9kLXxgVvyTvE6WNaph
up9LQ5VQxbcc5p1IJma30CF+cFM474PIlvzz4IjkXN4m81R3f/GH1N1yHUSeZisF
ns4CQ9xEo5tfKhisrlYgm7k/mCM3qkpHUJu2PvVNHRQOC6OTAungSuDVPIsJh+B1
GAoZhXfLYUay3j4Z4ZTG1X+zb6r8Nq/7mooq2S88YooUCY/dp0leL5Z1gr1j46ti
eelwqM0c/GlYC1vCUI3C92ADomtmXKl0B1W5Xw64/Qm+mpI05CvjyGOUqftWNtXI
zEXzrqQaEH1X8fCQXZp6M/pqXY/k1Hs05FEe15eipvAiyfy9oBSNUgDZqCd3DcZx
d/ES5x6Q159L/Gaya2MNfcd2tOqXw6cclXKtngiFI7myKEQl0tvg45fZm8sxBYkH
2rnXhJrkvVGquIDgSjHJJ1hFwQFNjpfeW28/ZCgHXsVeXMYUq1a8QQVLPgeIajbm
hyaynf/Y1JTbanjg27n91UK65b3couMOV2FdaPi+VB4ny6w7wW/dmEuON+3F1s4a
U8waMz6SrvPnEFS0n6f/2R/KAsOZv6QiSD0Vo8HmR8B25dmDwvbG1z7KrKtangp8
4/PzgSqe7vvPkDljyLP07dGebEJ9VOHMvF9SoKrzOQl1ICtrjksrgs6kzix1Uk3N
BQTCXyrMgFPBEEL3FpX4Brqpm8jTgFpuKCH7SN5ycR0DTBeG1zmrotLEq7LV/FWu
1rTFXph9JnnDq6OqXaHDrsbw2+piEMnPZxuUaud01pL1nEnuxfuO4OTcjgDDgS8o
6fVHV8rVkr8QUEgZuREu78ga0K3WH1TyEJUIn6nI7DYXgIxsWVLl05VIv9r/dDx3
hq4w0R4c+uL+riGzWJEPyXR65XYqyRiV5cbdp7VY1WfaxH3NYgbvaTzV5eaFG7dp
lwGpSVf5Tfk/h2PzUmwSb7cG9JA8yAUQX/2b3+VYe4UWeuioOeQbuQOaP/3xb4qR
l0LMCYAztDfVdcIj1U1MqNxb9vmW4j4RL/hng6BKCHJgiFqaEATTiw6Auy1I2qZf
PfG7SrIlpGsL57TxwV5j6P2B3HOu4x2MM35w/mvYEcIDYqqDc6C8mcdUUEFf3H+p
/PZWiOfIczdy6zDhvjGdVdJU1L9DFggqWJxEJStUwYX+Jo1LwMdIkBeC/oxyA3SL
8bIFSOv20IeDpjvGztbPyi4zFCOd/xF5wmtyhTfblQwhYgXPwexXve/SqGe7ZYdu
j0dlukjiF+I6+cjYI/Hus3nGG0ALbuDQkoLwABHUXGf8xxuFUFj9HQcn/Ff9BZhF
mCzkxi2TiIE5eJuVBSceRJnVVXcWiBof6ddcnejws0NFNh3Xej4Em90sTDu/dhhs
1UytKEUCaa0JECht9s3Lu5TpZj+UpeQcB09hxklHcVuvBDxgbGejmP2ZEAOVmXWs
G3ZHX5rbClcqMiNamjEz9CnfiXnbcaAnKXm4+T07k8RoyUoPSXuvLg5mlJcNJq2G
zOl2hX3oB4Prbu9KQxJNVR/DJMbBKOfx8TStibqSUun4tyn7WfDX7ja054ExL68v
2RVAy+d2Fi7tMsV0CQG7cZAZJF3YwGydAkQTcqmC9/HbHSeoJmYIfZQAW8woYZy5
gM46Ov9lYI1T/uY27B4daNjJ3QpXMB2eV/EGOs0oNA+4BD5NbInE1lpe8EGctoIj
xlAbn3/lHI1WREGBfHYwfGi0Ba4nRwuus4exFsqQlj5Ch6rdREHFrkWfAnh+EJ6K
CafR3TlWfdbRuAQScCFGpu297040PYQTV+/gdlDmGTVxXLKyqP6YW+50uR8oXA6V
T6m3itLq8yvVANi1N44xWAMgok+plsU6sFp9RlbDnUOyG6pT+NPOE0+Y3whHQpDd
GxClfdhqALGPELjuy+N/MiZ1wmMk4hgwpLJfX5HVscN1r6WYvBKP/iz0S/9TFMWj
hotHdSCOx5p7PfIhj4Ug88P+VCFD/EcQz8nPjSRbb9P3k+mtCWs5fIwJ9hoLNZZX
U/8MyP5rz9IbkkfQWzkmwVCgg9/YdxO4q0o1L96FciLLjjTIP0hKeUiUhzF736wT
3X1Wlx/FiGVd0ByuUQgUtHMYFBVwSOOn/EuNQmxVQ1J3BJIVSMG8Mwge+LAcM5Gu
Get4mO1Ae0i8XnbUqmFOjsuECl8GDqFEVH9ksxh0JyiDl0TDTgYxTgz/Adzp0Qp5
LL1BNbFmF8aTVUDAwJnMbUO296oAELSH3w81GUQGgySIXjWvfu64fnEQJJUaN3fT
rjv83t1qQVIrQgoyJiodYaSL408PvLgD/lXyo4tCHgTJuDy/wYPVZR7Dn2oCe2vX
CyoVhF35S6kD4/VysNiUAYnySes4UP/GfVo8JOnqjrR6RTsj1SyAkdZI/L3nR2SR
EVvqjx+yp2S19/mca5SxKAkXnnMY3ogMsKhFFAobB3Ab96rUZ4DK4ZiPVmVJ75mE
pJSRyK3umBR+scbp4RJfiyNRq+qXM7+l2jq9Tq8dQbEz1rKQLd3Cfoxjpu8qnmyg
dbErAkWVMkT3XX08kkXfUAvNekbIjUr9dg6KX03O/ILbAnscfAK69Z/RtXPgQ6f6
VasMaJrfYoOdzJTAwWPl32e/oQaDiTXHBgoGQBHtIZO+UvbF00/ZXHtjtwMixadl
V1vnDhJafezimmA9aHrgGgDnDBfj74KbkyhRokyrOjPi4Y357SEgLdAjhJYTJdjl
kmX0ZGXZIDoC9jTn1zzPT7GNk4yfi9FJK16DqdCwFOcynB/sQL9lWtfNSBICVkFX
4Oj/9wOhTXf5+91NoXChKfIFYDkzXvx7rUe2QbmXR0g28XwgSFcc68idPL8lMvL3
Z9f8eZBJMqxEIJy8wE7YAF91Z1w4Knkk47Dp3z1JNgS6q/mCskdS+DWGmclDmrfe
T+2f5fIkTqJvtEStC/G7fHH4XBxq0hXNyhwiAr5DSmh3kDZLKxAs0LYLPbjIO71r
fsSWGEWrjJv5FLFYmqNi/H3lZrTyzsUXj4mKOMp3Gp/1P7a2C1p+YmyjNFB2Mwse
91rYPYiJUXKOC6mDO9pqnGZf4v8vVHDYv9OfyYKkpzIZvrTszt/XfKHV8Ahrn7su
/Rvb1gNaYJKknWht5lpUaT7RWnB50YUfAMa84bUEbGiwa+LiXCjGA3s/zN/XOACn
Ph4gYgyD1MO7ChFdzmfFCTEJI15PrAM569aEXrosF1zhTW3gsmgQY+sx/iLVOZ7K
Mly1Nms9W+LUXtyTeYeraN4YyytMun0u02KgJzlVmY/cVq1HpTyiEDb2Wvav7Ex9
GmACD1KalAkwtt/HnEUOfpigbk1AtoSr5SONYwAe0V4ug7+xiApyeEz5NI84lh3Q
O0ZEkTLEyGwQZfZt8InDIPD23ZlBTT5AldpACra7qFlOOITpFQFBS6svhdstp7Xp
8cRCAk9csyGdqJCqQk5xLC22FMbsIRUDsXBGc0N9fv8tuWvl3Kcyb03/qOvJ+7lz
K1/qhMn/Y1n3FPR8rLeGd0j++h0mNzA6GA+jkUnvwN0zhmGP/X7iea9dBbj1Mkg6
Ws5GpIETnTnIgV+0BWfmF9rSklvmlb3lAsghDCNkS0C1N1DTc8eukQFd0n1xEE0m
dCxem7Piigz+DFORs1xgWGSILaNa+lN0oB6+oF9JvU3CUHzU5BmW05R+ZFgWIOYh
HGiZWsBIyPvV4v6MSmB7H7ekvyic1SxHqfFChUi4fIKxeVXDl21groskDZGnR3/1
9T8NC67NXXLe1mc2G6nn33xt6YANfAN6fhrsyKTx3sTZUQDxAVVOb+v856kKQ2zj
wLCc/WUsUAoC7z1YEnPmIvhhfBCiztSM7DERRPDVK18qRXrS2brGscZ4EhJA2KiM
2+qtRnzwGjxAFngXdHktPZfYkpBDZYJuqoYv2NgiYPibOBAZsUavErGC7YBlqldu
munKOTSeigwkpbCPDbStY/7ASrxD6wac8R1NdUlQc/KJp4pq3WZrkh+s6uP8h71B
UJkdawfssgJU86BgDwppod54Bnnb6QGsDsM8scrieF6u84yri899jwl4hTog03Fy
U+NI9aC2a7SFxAo9dFiwVecX9nX6nrSMttu25LKpcZF6fou+lmxiO3CCJ/WPbX23
xWuxQYgS0QB4lII9QPTK3oI/C29GW4G2bZt6Bm0vD4PGO+OADTA0mB7RUJaUamil
ZcJNjNVZuldSF/TjO58bJ7v3LrErW3qiXZFrZOZb4GKvAh4q9UpNp8F3b6YBi28X
b5eHzBpY55AWhj2c98RFTtL7QYQvzF1ey0olRuUHteFOno16IaRqEEl0xnWM1n29
86mlRCzG8KrRaIMciy1Xw9vQ/Y7HuqCVcgkEFbUe7NWS78fbncVyYKTnA8KeIRDS
7JBBNEgOQLUc5YD4nRd90xE8oxwh/53vqviuD+VbEyN+cZ2JfWf2/pFPfDErocFl
HztBO6Q6joeSn3cCf5rrbXw+h6ezFYUpce+/DFTAgOPEhX/yVkAFvOmXR7YC6XeX
50B1avpOW66JnBzWyJ4q1ejuqPQLPiahp4s0sNSjJi8PSl27MT0MbiHRwM5Gv3Wk
XisOvJhAyhMvFDD87CIVprQCaP2PyROITQpEdI2w+NS0wP7w1f/bOzbGBHcnxigw
ady8yLr4sJlRBy0x4oh1QmQ8MgbraNYCkOCrGegN9e/uSKcCgpAqUTy69SClaBrX
zcy5sgqtzEz1DhDmLqAncsK7GyBoJUr9uFe2H3MDDPo4yA9L1npyOtUwCNAq1FXL
uIR1ZlZXW5ppd7NTiZ4s72+oegp/bFY3nMyxMS2m2anG8+SGJyU+d72Uro5iIEJs
OhwzT6OoS3CXcIYuSg52fYIWULRlP8OGtX6u8QunjDDdbx3qoILBP6+939w9V5Yg
v6yh/Jo4FywW0G9I9xMkz46nADJw/vziEj3vhdRSipsf+u3uo2JyKWPdH96e9Oc+
iuY1bMI6mxeqPYxI9NlhZ1Q9E7l/pJf9jtx0cB9lz4itpiyoeje/Pqd66WhQk2lv
CXdR4m6iIVFVylZsbAepf+VcAlIGc4VOmLs0I1KATtBt8t9ly6MofaU9+C0gEKAB
t4L4cL5WxdJGgfYy1qmeNOR9HylfJQkvnzHagT9NHeUEItnC5F4di8hpQfSu5z/9
HfuCsM86yJJFN/b+dz0zVLMqBMd+lkVzEMuzqjzK3CLbcXj/ovW10o3xrAx3gySX
W6btfcsAjNAlhKYRQ0479AQI61p/ni1uDCpssxGEHEkGmKUzGEDXX5W2rXUbChfS
CYhnckuaf5oKm1j00UBvrSczbcup8HxhW5ios7EAspUAjXQA2MXU7Uzmwq3TQK1/
dzbwv9+QYw6unuWjNcUKsIYPgFBt+CcK1LbVGN12aR9X+iDQyFcWe7rpHLZHPxnW
qNynCOjGsRVObr5Yo2GZaIm4EITAWkTCMMtF+k8ubeB9oUbEiwzPk5OJFn5Q/sBz
J2r5axq535DVBT8qfWPjGp5N1rILAKJoHtdr2YZCZ7eX97rOUQ5czCpBpDXJImZS
YSzLH1mDM8Ynh2Q4ges+NE9wnYt+294kiOzWa30kS6HUgBtlAydL3Eh+Nk0Bfqil
8+xUIsIHR0FFbr9qQyjYi2jDU5ZzvBjFxXdqVferybSTBHiMA5XYF/OR041JzNbY
K3AzDKthKdQzF5zWYQuvax/kYw1qXwwDWM4fsHFiChn839l58QzYR03b/gl/TSYu
Lz7pvtttPnJs4P4I8aWfLUvOVXmlFfROPodnsIa0uoKklAdkjiGbQfWDE2BeIaR0
0aXCf8c2prEg0k75vw9FACBcf15/41zYLI1mQjvXIFFTd/iQ1u6c7axLhDDF/lov
DG/EjyRQ4V54oIVGNBJAhDWOKUkCD/fdZucnuXvwsi1L3N/q34ETrCw/VL332HFa
VfXvDm6jUNUCqT+X4QEhMdXJ10UeCzxdy2c0Daq4EH88D2E1GOblD7lR0wUKQupL
BHZCQm+9m6c9SSY8pUT4VgOUqPFUy6p9nat5yJ4t8zplYNSzVgqb+Xgl9k6F+yQf
x+I0D84BtWqAzcKgKSpWJINksgVUQASXcCqwAI/4/GflF050OWGnaoICMAIcaUaI
W9tiO10TzPYilqwmVmsAcDjmVpLpYnR0e6eQ5NGlI84nRLBqd/j1MsHZqXbFvsvG
ekFvk4V2/JbUMgsMoXfNhIb5CEKcqXhJyf88Lrmj+Ur7XV/bq8kce70obOxa/N8j
ScWD2bFrS2jpqs34MMqZCQ57r1CaCROHmuA9aw749oR1Sk6w6O3vD6pYUe2nb4jp
/Ve42SKygtvPsdaHWAHY4Zi5tgElI9pKUOaoLvmSrgiACB8CJ7BxOk2fkNNfoTbs
qM3RCd67aDQ0sPN4Nu39j+lqkRNSE/NBNFKQpar1z6yRijlz30IBGHUjotSXqJj9
4yD8uJCTsGq2ja8jkVCpjldalpUQU29HVXvztrRjljjF0UOhSzo6MiL0fJXY4OwO
GpQ8u3tjnw3EiXUmOuPkEKGd7khGejHiWQ3PRzO003zb6ZT9oNHHlMAlX9+4xIRG
ozyvqXQXp01grtDPPuJOhx5ISjl0V5hXPzWEtuENKF1p3PwTKypt1F68zN5TZ43s
35+8FXeOiWT/mnRs/jtHbt+gcfwNN4Lk2eyrNfoowPNM/tUzbswblmT3vrV3iLLQ
HKAqMfzy4kiKiSNGCy1ZND1D7o/1BZM3NjzRs1Ms7YOT00CRlXARI3ASjDQKpfQC
CTkpXKs9owbuJVJjwevu4Q3pYYTrHMRUSu4u16TDbhZstrNp/JdCHPYOJWN8KLRS
RvDybHxz5XPKAgPYCgtb5zui2vWRDHzKYPXy+VtEQHRSpqUhmye1L1j0rySo3GiQ
RUSw0xlcVsSBgq3vMcCdUa0ZiY3pPx4++w89Ate1dEHhi//ufTCJe/R3oCKnzCFb
vg7ZcMna+18dnK1wI5JzD+aAfH4XFl1lLbsAjx+u8BrZK5M7er3D3555NsFHdBCL
0skc2EyyyUinm6TwubxvnqTkvgOV7YCzLnAKp80HFlCe2kZX0yhh8thAfjbCiIaH
5bZLtP66QPN+tyUeS9T7SFZf+0BQVOr1D3AeN0/w82MdL0IDxWVRPOv9PjBeaEFP
G1bC62tlO2RlXKjorKDsy3A6xKT2TcoRmbwt6Di7V8LVOt3EJ3KMTJbgesFC5Q3N
b19yeCqwLkPx46ymsMbB+K5kkl+xJhAUfHO9B6DUbFELoAzVHPbKbirI2xqIJCFs
Nbln/EvA0Gt+6r8zJKtXlW611/woh/hBV3A3oVmtXuTttPhjcpMVAXfPyPijq6xL
ABYUAUYbFrGPn595g/Eqa56LOAy+0jLxqAMPBU54FdEqfWdlEV5tQfClWuBOwDLD
TapmBiB2JvMLbNiDFtAwf+XdoZG21NT7xiRbXxnsLcMWBhd1Sgqxa5s0T8FlUzOt
bFEfbKkhuDvE7t2MbU9bX61iOeE5kkb6omOtwSTN983h2IrXIIZWiOLDhfk20wgc
Mk7TuHc9m5PhnWeSMGSuZ1h0UuXwMVxQoIzJjuJ8rieo9zjU9bG8AVVfk+mMkVfy
dEHjaK+h06Z7biKCJHCeWawyw4I76LblZdxbohf6mq+FcXl0PLhqLMOpBrmpe9Md
N3czDkJuvJbUDtaGBBwOIYS/Dl44PRZXc+IT0ffdje7bhkdBk8+0N9r6W4k07cFf
1eyF4NGNaQcxldTTB6xvX3rJNUIpa+/zbdK9ueQ92ssogiCi6SxRbjyyYnZjF6yD
mp6+yuoSQ1+5L5KFAolqIUdbRwYsVJLInTrH7cR58yPZPIGL7nStiNRkHP2EvYiY
tbbh0seKRtGfCiuCrsIVoHB4lFSInfuMSlFEtXWxl5aeaY+6pwu80ZSpKPpxy3lt
DzsBsHw8wmixNNBu6M298Aw1YRcun70UIo2iN0mXEx8rkB7O3LgsdbFqyQgvtj/i
RfjZNGyqz/ZHGEd8Okqmy06RcVPjo8BM+lq1ht0Hs4WxXEKVrzvTfFgYY5zYbJ8O
RFo5mcgFWwhJ7sthQn9/COWKTtOcpobIOEEnUNZ+PH4KnlZCxxuWahoLP8W1no1Z
9HNuwd4BgfL11RuGCUBJkGf3lb+uirfboG+v3gQgqFs/HF5bxVdxM72KEqIeAh04
o8hcnvyVIcCVt42GZFYtskPdSaPnb957pshiZ4am8SMM9nE7Hs7tX7a/Y2xW3JDq
owFszWxJdC328/OCHItlBzMld9SVYwbwvnPxNZem76lKxKIkOs0juJFeneTdwdQ6
YzXRxgaU1ntDjocJTx2cYkvDM4YivCEm7ulSIJ6xx32PpFLK7cQUHXTkwI3lg3vU
/67XFXhtp12jHHd3/iNf4lyntb7PssDh3U8wJAfDMj/mTrbDLX3xOaDU1n7QBDAD
YumNh/ZzE3zJ4ikOAGvWFKmjoi3jVW56WOsi4K+I+65HT5mRi4BX2G8Cb6HLxl+r
4L0lyo0ZEpDtUdRDHNgUaV6S1YUICuOsqAxqHZrPVeaEnC9P4SomoXqFF0QGCi1i
zKrkxsbo1A2+1vptGhGb/zVDFWlXxDiCGjp4074OzV0QcSmsbImPQWrB5PV4Y04r
3usiMSjqKB9GmfpbTaSgTRRKxjVJWgJCRANf4IWA8w0a9Q6PgTYplPwwO2RPWIPl
91xukyPMEOSk8rMpkltbsahXqHo7RG7uw9GE/Vc2SBo9w6KkJAFSH9PHAuel++1h
QHYYvOvcF8smUF7iPOsuFXnW5HP+TKsRSoyody7Hy+/kJioejJ4cn37ZyuYkdH3W
pCj3GyX6PYtIdtQOpnOaO/PRDIL2TU4xXIXcHlYUM+PJD386shC83Iqud2XiAjXq
B+l2BfGOV+7oao1UbfxFI+FzCM9co/XHozy2XmXFOTJD2NHguH5QI0EV0bf2PzXD
ya0xrhwrzUw0wrxTch7ayR5+vGDD/iSUmuFoTTWbXM0UodydnLYm7fSseprKFnvj
lClSPuMS7AJC9PJMc1puXsOwgLvwjD09nvrklh2YPEdEQgTDpJLdSFNMRlK5NPDx
wxpe6gHLqfPgRY0zsF/DgmkkQwoq6nrwXq3Ftv8/PRJ1WgGItY8dpCqfmsJPxfIY
nCCnMp4lwioVTI9AKE8w6Nzyonm56rh5HCu/4BJk2fu7w6hUDCSnbd6s+fJ+1G6O
dG5r2PTWCkRhN4HPZSKfGir6dHzh5aWSol6O56rjlSnlzpImzcc7O7Yc1WkczAEJ
EhnpjGE2ABRwXlsSMCHL9K0EtP/6IWqutx1Rds7KYz0pENIIZMNgbqJgOkw4wE6l
7hxQ1U6M1alEYb+UKMGBX5AwzGTrU+JuHgFlwEoAF4e3btDThENNg4+dxhgdVVMB
8r0qcXeorzeTXJgKjRwWSHgf6RRZoVmU5Tn0lWE4CLUqT2XUvyINeOf2yLbefb9U
P2RPfxN1MMe9mutqPdQdiXQ8VxKrsfO0spomHKJOmkt8Bf614ctpKD4PnGFm1nF6
0xeicDeI9ZIE5YFYRFTdnFH4dE8lhIyvWu0rZPfYwfHeVW19JzFbj46P9t8Vp6I1
i0VrqZFnYJH38CqW+e9yJgeOMVWdNnUe2TmBuURuy/q2prwFRgmscGEfhcQQvYYq
SxWVMkKhWyHBjwcXGNBy/BsdEUFdM2tERjit8kgST7DDmiq3U3AJfoK3CG1MempN
m3wH3prMv7oqFCeMRtI1/MZWK+T5YXjN4pDNrsKaMDcSU6G5rBot8hyu8uIodcZf
s5uG46b6litMrifLFAjnyKFUedrVGa+bkLqxXaHKH/iWPfDj+uG3OEpANkhFhW49
5EGbbghfDfEUuIVFwL0qMx50IeH4ALUEVKIeRZnEy4rlJVGq2RIApOGwjiGBULek
+EkYsqkqY9VRYPbqvvvyAIwG8JZiSRO7hPYNVnC/LPuSQXyP1MBEHuuLS1PNjCHp
c2IqKRtOYs8/NirZleN0ZQnJ9nU5LRbED9hBVwj1kNE8gEl1eZGEpXsbyxSkVZvE
9kBgXCSMOu+Sgcgew8rk36BIMgytUvvlAhxFeubazsytDv5vK4q4RM6HH18rCQKz
GZUTKcgfAtQU+XvGsyEs/KtIBNbDAPStcW3mjEUFOZ+XBmLjyhfru7IP2fSG1U6E
jbPwVlVe861xKEn3aoDDsnqimTgofix/eDHDqWYowZgJxSpXIZUlOjLi0PSb0aMC
RYOeCaHJ1XYuvHZTWE55wgy/asaUVcZ+UGwXQIRSbXpO9tOhXIfy+yCyK89CllBp
UFlOtvJBvHTvf++dfb4g5Yz0AXqz8jWkDhmT3N4SBYsgRzykY46TZCQZkUgsDjhz
VFHSY5ObUTVTssXcZpV6PpbJnAgAkhkdasKiORxnKHv5J6GOgpJYg0x3QJZK84rh
jzejz1Sf5o27NeIr1N01wTd4O4XzH2GZoFGh3aA+L3kKSsy61G9BPHJbfPalw6if
HM7DiSURhmrk8CjXy9h2C63J+2K1KVVKGN0MAHxF6RJkLYoxgrw8Mw96w20TEkZ5
/10iUClEngENs9t0dYrihSlFkpmnMaTbniB1jc17UKyVpIHo+aYt+tWszHvxkAyp
JAxc6TyK01EkV93wHUbnDXKzc7a8C2TuNU96umuX53RcOsx6uuGx8X9pcxQJ7RID
GE6svz+N44951fnnHh7CTWcDSonjSRKFQK/BAT+1Y9F0PeKrWLGCXWMNfj5flJhh
6Eq1r7yQ3QONzu/UctNaM0r0kqWmwGAIMp/hSwSoUAqOHtoGmBhZeWxV3RXc8gTZ
64HnUI2S2Dm/Mp7W87BGtY9EMlJ6KAkI74FMm9T0ojlzmaAT9m66LM71TSdHzTFS
yZEM4sEtOYcyXNrAcMUc/2xJcgFj+IUwS+XQvDUqtHECycqG3LItQugtzaEqcvSI
fFS408EOJ81/jK0y5CakQuh0LYHQGVrJLB3IdWPO6P+jjYTz8G7rOqBFUWacoYSf
5yK/jW57XamaTaA0BnoDDZl2NJ7syMa4EE5BhDs2fcd2wY5PBFUMv6pYt545LLmx
xHKmPoc8R8Af8NBAQjchvkYxwZQ6z9Rj9hcTFc4tq0/RmvGuRTAa7DI0Si7dadvx
edXpGeRSwKlgFqH9DcVI4W7s0/NLgGq8lPSFh81BhMigVtvL+lptccbz4JGhTm57
I8Oi/v7GLVePSuolooMKi11OFJqpXUmUQ3HnPjZz8Es7jEjcm3NJGJWZuT5Oc4A7
uoSnM233m6ScSLKEq1JPm9cUSBt+BkCN8StLg7RU7kbVJyR6scnYvQMG918mC+59
6MGsptY6fsO1DQJ09xJ0AJt9ydT7bRujPD4047Q37pLElRf6zZqbO19Ps4yYUMdg
akpm+JG17hRrMhVfrTjJ4meh/Dw49uGe1HOCchr6u1c6rJbDNfMZet+M649zcj10
/yqPE7WlSYHjDDNDHD5E3Vym8yUpaCjLcjzpKW4xeXabPHmbU2+kr9DUlOFvK6iR
qxHr1My83+9nMDPToOCpdnWyv2MxN2tzDaZQDTXJhEZzJ0es+iWQpvN8zNSgfwXG
SdPwFXs/1SPKkVESU2dydxeVDgR+I+OVmub2HBh8qW0V/vfJLEHr9a31ldD68Kpf
L1/JMj775BICpWDjr6h4QqykBr3W9R8KUUopWo4GFvWUUQCbT6+K5g6FBVmfTthC
/87M937iclkLfQjL5BvoTdEqvurGxEoj93tGQOnAyIAOvM3nGpbP6+0CFgsPvaRT
EC0BVRXiBOxCR3R/f6lyTSpmMz9TfBNhM8scU6tVE52vQj7yxmH9BaZP4FMzKZX/
N5VuoFd8x68HeQzZpS7ndzc4BdlGYyj5Hhyyvc+ITyjNyju5vij3S6p6+k/3165M
IJWu8JSADinCSwfxq/8nwKxoX/YNe6DR8aqzHu6/FrmHQgr2k2t7mKfkgbRa2MoX
InBa0EISADEupzgUw/ee7rL0f9HS96eBEPBOhRuF8L1dt6Cd5V8q+RiuFGOWmJr3
jdXjUbITZ9evwHz1PopUJPMRmgASrG2Prg4p+CsuFNnUbIkzpDA38161GIVKfssf
56nTJs4negh+zWDxJBNZDn8VNO4CMMDef/dQOE3UUAEf8NNyn/mAlLmaHevcp2v5
VhW75eL6IQATJDSXlORxgkFLuifp1Pozm2Wn5t5DjRfMGl4RLQrptehL2mejZ5MA
wNfJ1FhrS5+4X9c6yAbXy95oqsJEVvJGqDVroMo0oH2EvSBNwmubdQxIOz2P0xd6
fJ+yg0mmngaqEk+AxMSi7VwzRar82xZlLECxO/DXRhXRz8rbnabMuyPz5u2YsxCy
l8eg56RpMQnDB8ltYtfRzgkcmyfNr+v94FpDkusBgYpA/FgYQum4XH4Z3dIQ3Lyh
fwRpCdKj0mqpJZo2Uzq6opx06+scqHOqI41qfF3xkOdhRUzpO5lFN7T++HexBIsA
lAWY2lm/CJWGnc5oeiNkdbSoMoed1+3gi64nTcJvN5GhDlNn6BBUEK2HiCTpc4Ub
nMLNhq3CafHwTFgn2+ipa267ADddRDgZFFw2i0Vq5KYsjqnT0liWuBGoIJYgjk+q
hUsNdWE5dzcgZbDt5NR33ily69mmujH8uBFDVi19OZHmx9HOAG/rCpMwMhchrJZ7
tqwyTwJxGymR5GhYoA5t2S7J01x2lv02YUHbzauUWAMsYmRsLM6KV3htyrYAeyxN
SEnUm6Wqr+0ZsTygmxgacxjkZzpXx1rqSYESrXUYovFQctONICrotx4kfvDq4h2u
7jFNqoJEGnM/Qql2gcdKlEbL5Nl6mtswfc5xFgeuB/UK53Uma1k3dhuiImxj9EDW
hFep+vvt5w5j+1T35b9mhEm2OfAD7YaX8Q9eYSi7oN5sxDNeb+giWt8dfEQ7mHD6
asHaVaa4qaUFJkK0N8z7ryawATcWcTGWmrZdsQBXvEGoxvry9C6DvEdoXRQVu77W
dWQq9/Nm61IeM/8MvjrhXlwb955gX+hEGhfHU11LQ39qmi3vOzzJzdKbqrZli/4k
zB60ADbaMBIej2NFzNWObMrNL4rVqLFb2cZXkaBG4e1FnIj88ALjKtVN4bPMtEfN
y1JvTpW03xCVVmMJ9ebs4MMxQIKSkNosZhz5csCrGAt5Fp+HIGeZq5TCRv57U1qO
jGBElk07hBjQkBElENoiVxgMAqD2MIh6JUsfTUvhbim90rVL3bB2ecvdxLoi0fE+
yNeTvn490orJsIBWIs7mem0X9acPvo3niykY2jgz9uRceoGEwGiByGhAapB8v/Io
J9/V9F0UwALHcf0BR8UHYx8ONUKyDxzC5QyRR0z9fGrWkldusKRG8uJ22hk2PmYx
dGReuGjCocCWFzMMYRUhzq55PAqsCVNzjJpbfoeYn7dV5UcufDgQ5mZptcG0Z7Ms
vU99LaRz5OavwmR8eXGuZSWRjgKUVYxNZ/xoUVhGkQapADQZyAR/QalMoHOG+Kt4
8BFb5ziSfb5coyUh/ExfLR3ESQ6vqXlMESKIHlwQmFWP/8r+06XEzdMsObzPdgft
1ECYLEaQPAU7zXxM4UlKoXWvkC/VLEtrYuxIqgCIcflv4rn0BZCSC3PKarJUNCMP
up4DjzqBW5n4g5phXi/ZrpS6iDra9FqP/yTHSJEKV3nJb7PNlZHYNkRWTliy7lbj
8tiX561Pt5Qvzfo3nXkmgZnHotMUML32QZR3XMKSUzU0LTKoTJ1AITs/cz4w6FwV
tnNkVGH/0FoBVD1w6SSI8jfXgTF2xcEjkFlqSEck5EuagpFSeVOxK8BBz4m1zCno
rfwVqRR/OJYpQX4CB+Bn0+CQTAkj6o6jprz5sT4Ul8/ylEMIHBR9PND/bc/RWoWE
Ocl+GHfRNeEGbzBNGtLpDRRaGEv8R3W3+CMQGOBt71ERdU/oT/iEabBs70edqIWX
c3lD9bBbHoxDlzIH6qU5KvCYVkrFGVtvHn0AMmPk6fArSbMRpePpmuE9H+XlAp8l
oEzZfDY8+ET3FJWQjihNTEW8NZwxUir55f8sA8niHS2/sapTESsoarUpEvSfaOLf
H7BvBV/DM1BNToCjuGClMUHXGHTQrREZg3bQz51NauId2Lg16Z3Rw8qSH9S0nq1/
oFaX5NGvHew8DXtOg4tnND35cJudxTRQ6MiUYfsxF1CEIqUIzq1PM2IN/zJfLJE1
utBJADvmVRlpeiQ+E8Z0Eu0/IjDGyvTDQF4n6rpjHX9+pF8PVicGH8T39wxUFcjg
IcYTRk/7+pgRi1qIgxLwy2TEIKn9oPfBrS2YKEycdSs4qBKmoKNoguDnHbGWaBzl
kVyDiULp/Ah1+TCAXa8Z9yMySXQqN797EXJQkHGS/idDRzaPl3DCystZ/J3/VXAa
p3icvWpfXm9GqzX+YEPChfMnLmCgfvsbxN1h/36f9QBK8WCqeGAbRUKHBYZP59pb
327CmmoMjBRVLuDWLx/Jn6UzSQBlhphCSgPjcAEWJy6KPvExe6QTa3ogb041qmeo
Zfz4e+mkgjSqAUV3NzcwBfpVKTP+jymWZF24m+GMYgCopMOaDK0lQEUZphTa/ZhV
yV3ntQy8IXwYsaxMAbcJwkqK5r6X5JLGZUBDBQ81sf68k1ke6pZFfTh7Y8m5p2XF
6P1zX9QQK60wrXtpjmk0TYZakNNjF8EoImq/dndnn1VdyDUzfX+ScHKXxbXym5ZZ
8sYZJedrp0ia7Hqs9/si0sJycZFbAMW3BARgtb60rbBe4d1/m+L83d6yK+qVZOHe
/LifF91hRvEILKJCFQfkfdtH70kXj12tgaC/5qF5XzKYKMckYVbhwW0MOvZ91KVt
9b8aBjqSJiqKi8sDNg4i0uESzhxUK2qu7YczkLbhpx5rDCZNAK/ZDgSnlerykN6L
iAUE/i7C+nCqRkAXGxHmHZ2pg9ykvg5fzLkc63ZtYlMq+eQhOL1PKgWRimyoKkl4
aAUQCfStGTPWXaazF9AubJaG1b0/Nlg+oDvVLUUAUzmkOpdt6AVs0Apu5FcU8fiZ
OHrmyJRTYMdT9LJwE7kzdq6SRHnuPFnXAsTAw5+yZeYBhO14kQkjTeWsszxgQ1Ig
EQZ262qOYCNzTdSHI0FdmKDXnB6dpkUH31atINMJr185MfL/TWwWLdqOV9nNaxaw
MWVqyXza3CiU/uYC8k3XIljUMIkmID2wBVplOdyn4KMyydRp/2KxyKZUJQqMBgUL
ZWd0cNM9alSuD74Y9MeVYwoKr3HV0tgvYYsoZ9bhz55lvi6vVDH1a6mJK8p1jgOM
br1TxxBXF4nuPyYS6MuLVXAa1LzTtcShiD0l66PGHhcRxOFRzxaOGykspmOIiK+5
f1j1u3o07LN4t/mJYH52YxfX0NFNyF3gVPTrpye8O13o+6G4+OHS7HsAe+1c8M6r
eS9oI0VxVvKcfVgy0R3HGfXVHyumgCI4iVimTZyquAzjcaUa8E9QYQFLQR+Y8Vc3
ebAVwmUigU+5KNa5MZ6tyObaZfEx5XbdNfD8j/Za4pAFUnrLL9S2I2iMxvm3cFJd
pr7tlfG/q/uAnTISeG6RLlHQsOud0/6zE5BqalHGXIhgkakxX9gRDBZoZqvbcAQC
iMNImu1hjTVNBOseBVMfcp3EVNK3ToXG5TV19upe1Jf8NHQsaX+4OxlttHct1rSf
DSVDNFQaWnERl+8KLhg4DEue9BGG/0cljoDOen40ypOHi7JRT9hJ3RSxje9yW58+
WqP9t32PoTM2fF4pUkpQPeK+nobdtDWb9c34Rp1rV5+aAPMHD3oeLp80EBbBJX6s
Wo2blJhTcCUpOep/IjdD5DmhTgglfM0jncTVgPQDfsjrBVP+9bnc9HWsnJyNZkCi
wW+8t9Wh8NaSULROD0SSPGqUYhbrC4NV18QitzgC592wfHndbStf6MpR2WHh8SSz
/b+xfc/Ot5ZpFl9b1d6CKkFZYeopESYHow0c/VOxtF/SjELEzED2XxDURAR+mxdn
C7PTmV2PSGhetBksQ8UyMdIhd1JrmJpO8F8G25wlupPSDjQ7YRI1SYZzTfkUn24d
8n/Fbxac6F4aS3z/tBWRp2ee5kWmoRu2k1fJCaglPnXDPw1kcLITmKgHg32z3fHa
UIm2zzQkUgC1RxKILXojwFXHbPTYfxJgi/zXOmUWxUm29JwvBekzJYOPXYN44Ves
HvVD6cG060Zn1B1Yku7xk0UUI7Sh2W5U2Ysdb9lcBUJOmw9sTAQbEQOAUyoFOwgr
yAfklXhu1UnDC6RjW2UGtWOA7JyNm2xn95KtfX4qM7wse0Ar/dsugbOGAsjl71EL
tKzkPAs96A9Sz6TwqsNTBGjK0Fwkr7eaZJhf3GDgDom12g7F03yReeVpVrymj4Y2
VIxxn0EdGoKvRXBdAxLe68gagD86WoD1cmdULZKowzoCSzH3cddvgXWCM2l6oUvQ
fRrtDdjvd30MyDfKuNd7+bsKj90H0qQ1HDbaiJFDzJRHn/EQRX3pCNebajT5WXRg
7VvCN7DOb2Wb307pA10yIEkOam1I31mipO1EdFr8JvVd0dRAXOr4PGxlqwb4WCX5
GKhHJWNZrdkoLBSekOhY9ON9nrhowGwsQFEGQrqn8TTCGuxEQcFVQ9lwLrFW07w9
OLsvrTLiMIzsV8YCn6J6UBPXivxgrrI99eQ7Vp/s7I+jyJdKbf0psVx/ieOJl0i5
QWifWt0KMO45OVbco4PndNkR+NVI1e95JGNUB8h7sY5yheCY36Sn9mktsPdbiRY/
/Y8TNoa+du4gf7iZ5RyhJfWd2XTsNoNsZVwRAu96TvRr/dqcUkUuRQ1jF6u4C8wv
kPM4Trh89yLv9zhUkncXPPen+OjFOrtF7KIrBfi3xz4Q4T8WnbIgnHwMgvW3Kbow
pAtvft8TQuh9+VhmW2xQRtacrEuC/DQc+XcWrB63dxoUiEY2cFwELoYKd+nvLw2m
Bo7CHQIFudeMp5ZA/zbDVHB652Q2mwjnQ0d1jKJelkCPodZdLrDQjFg8EXi+1+pT
e8T9S9+VN6F3dcpj29KFhrCPaw2SPXAmoSETUqmaDH8hNB9mPW0L8EqfGo2jM5gS
jNX+DUMgJt3J9fY71De9a+Mi90Oe6tlugUwI755Sh1NvB6GEveXCCLEsxor67DZH
Z9PznVV/jQI6m7m1aNFno+od1Js8f5kF8LwUoHHK5iuuIhLi/mLP7eDVf/uJ/hBV
Xg1xVvM61Sd+8LCi94LN0t+wyM8iCxKOwPsQwYd0nOi9A3Y5Dr1rhiopcXpm5Ygv
3bwSE+/3rTZy6HrkcJRFsBgjv2pjOzx1uD0he6AIxUEUPzwxqG5w4Pwq7sXHvaQj
MwQJF/C0OyOCEqEVCjc9W62zrv2slqH65Kl2PAgTprlHGGMRWTVroe9/fQePOb7N
T7kcdqofvmrzxgJcJy+2eLqzu0EmYyVeShUzrbkGMakiArjuV+o5TncUoWC5Za5U
/PcuLXh3j7qX0OIpqqkfAy4vJNzPlgjFUMWhzKOGqQAhus4zXwGgsy56/WBZCotr
TwAloVPOW7rfhIbCGXHd98lVbrELYOIqM84yDKdx6ZBJ1j/r/YSK18oHmzCQ+O8d
fVwyWFztQpKL+vrZE2ey7V4yNkggmRci+2BOazkhqf5wLkF2B+5OXxMHPfx9a6gO
7FG2TyjwQFeANuXFViNrS9dxe8JquqnmYhK0oWPLIPrye1PGsPdyTwerRnAPdiGC
aBYZ1oEwyEghaBBGg3BDGAS7nobQVQALqYzadyNrVTfQI+aTNXshhtPPVD21dXcw
agv6hVxw2k+kBiB7Wly1RbUB+FSygy5ikzpSVI1dMiaZfzf/rd33wguCRSCmsdvQ
vXqU0C9a0atRg37/v14xjJ1iEaWqjFdPzcMmyAFYuWr7xdWcGsP3fPhzBkr1BGkk
kPax7kTlB1sMkDA0uhvHgoN5JuGLFfWhgR2cR1H97DQNY2ul1zCwQWFZi+zkd/on
AG5IMcPgVnuj568E3Q1D5DSrriSLou8zrT+7vexqi7j5cuULd2tUK8HPSnsooxAZ
i/uTVq6/1hVJOtY/ie3ou0Ih8PVC/vaE3gqEOb3LEaVNc0Yqa0uoU4oFFfPN07lx
2pMem8+oHL4SdDulj4Ktjb9J3bADBM9EXlXV9KMZU7Xa8d+rVhjEFChNtA8DIBqL
z/txU13d7jfVwhy1TWnBLWlqq4U7QQnMFAgbsb7GM2y8UTT0WnHuHARs/iz6LMnv
DqUm8T8ZbUmKMyznZfHo/E1mX/ICU/erDSpSLXaCsrzUxETC+UQcSXolob/9C0fu
EGP8QWDH6QgYMPvE9GjGdZOGSIOK96sNRNwPAKNuUwGREWL8jcWOKd+V/h1XPvG+
yeVuErDgeIbnuUq+PTgLd71NQtqcKDyvqqVKcUzVl1B+xZW/optOEIFbYCLfO5rW
Sq1mjY4ymg5AfOTDx5pkXA+JWTbafgvAOFulE/XZTU/ay4sCi0K1dHtPpLx33kag
A9ZOzJJrjJgySiziptwhyBmuUhGO/hnT4EjH7IHCDcjvRbXZhL74g9oxUTuQ1Qx1
8tTKdrLWgGrLB7YzLlTx6X4ikj5m3dlZO5aJzRD36VZGVjF8KJ0OvuqKCIsyHe5F
KTnWBc97qqfwunCj9v2/OUIlkZ6uLGoBAFR1O3VZwEPi6HoMjq8B+slMfPvPGtk+
QtgourLgg3Tme/Oo/xp/gHiflmlZNyXYtn+BMQLCHsQuwLNNNh34UBTnOVK0MyV2
jfnKE19LGwfll4Rcx4vIaW+X1wYwkU7iwUDudMORIEYoS9Is80MwB19XHshYdm9z
dx5Q9JkDb3musVBbQW4oVHDTVlSlF3YGZbYvDxLEv94=
`protect END_PROTECTED
