`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RJ06bkH1gQbuX9gP4qAei28+44vuwnFLVYblkx589w4mSSIBzkHX3WnbavXe7eBv
3a7TPdf/zbBkQOMN7n1Ib1bd6/2svgeSAcdo0dZIgdiTuvB6szp9fdyhASrr91I3
lfLTMq2wvoZGOyOoFMw+bjeS+frS/tsaYISO4Ca3t3gxgvBN3MNLoHSQCKSQzWJe
fBD6DyDstHhuOYZErajKIn8Nu3yKM/oU1P+Qgk0hq10F2qjebudz6oPN7XR1xu0d
Mtd521ytvjG4padPuY3LQnXUHqf7tZT1ye+VaGX7WxLBCtZRvZaRHMNdlAo/+coO
33xlK/uS9BlS0CxHPV57Z32xJClwUvnwvo6VkBVHlf50+9FTXK10zZwIvFv1IuM9
FgphqObKA+7NsX8cXxVEdtpH3tpfirIr4VFLHYq6AZQvUzsdQ6Op/iwncIVgW7Ad
AHanjqsfkGc2Fj0SC603Y32NCzPAOY6SSObLcr85FAU1x+i28NMMac7RMKKeH8IP
`protect END_PROTECTED
