`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6VSjnffQdQK0lQB4Kg+7Abc72V3NAQQjm0wRTW3dbyNKLgRnC9R7QuLB0USuaVO
e3CDfOAHTNj2MjcGA8H3hvx04QIRpelrogaamF9+W5ubw9xMvXPyucseH9GFkr/n
WhoO24BRlC0zYwkHj8tuLAslXvIeXi67C1cJmSjdU54nGBIAfaQt5+zqcUYDIi3M
WjOE73831RniePp+uqCPOyFcOpaabIGDHBP68QUfV0PH5C70mU+2YV8o7N9z6Qqq
p3QpbLuqfoS9RyAet9vOwIdmHIQa5Nrw/JyNPv1KZcGYM2qNtWObEBGAi1lB4k2r
NMY7ldnUWDZ45ujxBfZ1mA==
`protect END_PROTECTED
