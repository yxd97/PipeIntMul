`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sscy+KkM/H2iggQNaOjoligC8YsSJFmV4ThBIhKJAtw7F7rrl8UuR01nmD6HNgYv
R5VOmFutiTFQAz6DGAYriv9prklC/5VD8qUBt+r/JwRfEh2K+noOn+2xvTm6Q+lc
FH+PcdMJu/WoWsJGGy8dCdbN562M8cl0MXKoIsCsCcjXKfHIGMUrrQN9f7wg7s5p
+ymz69tfpwZdvQZLrjxLkt/W6VQN56BJuNVeSb3GIgqTQQV6XE23km0k1lsNIp9t
4kY7Q1JZKe1+5/6oSvxOc+rii+jBg+XugRKf4Q09GyYxXa/vHw09CGnde/f47DwN
oR1+tHROKdxm2pomsVyIBblfiPUI+nTNQ1LqvXHzY+kZ2CfO1RrBQuHbU1zBlJKb
aHUhi06TS33MYEVJgxY0fCiWxt6G7CNmSI3WynnYuNnKJVuy/aNNU07rkja5q8fW
jmop+gJESpt4uOegSanHZh/rR/mMNnTFzPwCw3WtCeORmXQdKRXAsvs1ob/RMYsP
`protect END_PROTECTED
