`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DFHP0QwNEzss1pmF53VaU2U8kwhTKyryRaFjM5R3mHFOc/fcf7kqkmwlGuZu1PAU
CY22ZpAQDPz1G7FH2kwCs6/G7hs4Q11dH2N7f5TiOQcZOGMuHVCuGkCBshfUPVmW
rC/PJN9nXJ0lgJBxj6TalOhDwBeTiDExxyo8BGOM5tSnlinbjHjdj4pmPYKYNoBV
nFFct2obVMlWz8sZ6w9oOw==
`protect END_PROTECTED
