`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gi06gQ8LmxxN0/Si2nP/mNUxRj+PYq8d8blYNR1fyhXMVz7jpRBhLSckwaCNWnI3
6PYwa8lqwd4t7tVNZqNfeUWcnT/sPL7iDOXsPNU0Ngc9pM4i0ShJSiBWkTbMguCY
TXmTe31okJydaBEySZlnhUliGm4atpuUTbDHrLW310JTcNjHCqV19cH0zVnpOPIE
WXVJWAWHDPaIwQJgooVebtw85Gt+QMD6tppIQkvYWUF/gDSW+0fukZqAw5ePcEap
ipVgkmrstAlIs+/4hlUS3j70uJKxqlUVMcrQji17jFTMpXHJ2ID6T/JkGFRrO/e7
sxx/2RlMKLu+Sr/eKrs+WcGm54twzKAGVbBiV/wYgVsbFSglH/JspfkQnR1ac4ZL
d/yDi3/0usVyVPqUR9oOWzoQoHvmdO/0WaQakXITstfxW+8pNCxgzRFyHDx+4hjM
B4vGW3123eArxH24fGGn3Z1eDEIkhsN7t+9HacrVPws=
`protect END_PROTECTED
