`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0S5JYxkUIzITqWIr3c/+IWTdCV1tT8DXolhaIs6UUfrYe8jLiLRguTeMI0C9mkY
MVRJqaCTKEbn0IdyL4kLA6Jgu0n6rJOSiXf5iXi/kzmxJlC5KPkJi72jGIZ5g7j2
L7hejSpLQ0K1Q7xH0rNUltjm6NKRcZoFDUQt1jYGmiYlF+oZ3lit2ZW14fq1yO4c
QCXf162hz/65QQg1FJnHMyw8M2Y/8keAYSyyEJSZ+19/SsQMzTOy+m0c3cLXux7b
EsCQN/iH6p3j5SSLvULspjklo+mLc1EU8fPwxElHxsp7fuMPKYUSFGs4Czew/eK2
2Qz7z5hNGnbTPEvA1OMVuGx+qFvyMwdBV4S+kM4OeujSRv19dR81DQunrbaxZDtm
z+Ia/d21O1oawsdsWHu4vg==
`protect END_PROTECTED
