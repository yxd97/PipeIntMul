`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I6yQ4RyqiEr/Eb5lbQWeSBiAgd7CEiVYNo0p4UaoMqlFltDkheVnw7TTrfoP3fd4
cTFFDdYJtnDxgFfd/ZuqLZs7LotEiv4rrkWhSIK499cwCz4Soxr6LvYyKwsyKgpH
AI4kpDW6tAlG5JEZMpU12IdloTGDSp3fP8W/+hplad1VH3DYJ5d6HUTdOkPxNd6c
pBOqg3jR1aZDpwbd8QDEjLWmB/KDY7BlDDV1VtM8ZBr4gErkgZGoEGfGuByCI+L/
Llk7ycJ+vIMSAYwqteD84A==
`protect END_PROTECTED
