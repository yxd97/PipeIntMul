`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ij/EH9B6e1+IE/zbEiVPVCloK4aL5j8SWnrsQHtytuvxPtYv7v93UF8IztVUjbDU
VSt59NpuI4TGCXCcX0sGXdmwqLlJ+MLykm08/N+aCDAF3pKyg6vrbEzE7Wyutbyb
+1PAonIkJRdJFQFgY7IyHkFm5WSVIKxclkQ8wghQI+hRWoXTJinOlyKpqBMdzk4q
ksBN0DGZHcwrDOGqu4OXshhyJPKNctmW5IiXKSd0Ft7uy4PJxOUCQIxI3uBYBY+w
fqCwsGjACID8TfbGk9dTJlrWClUThqcQEHMVjZY5g21Tpi3fmlQH0EgOprvY82bW
JjxHciAshImLjKTs7fgn/qEkWlPbEHdYuAhy+g/3bnGePeny8W/Ho6hW5sykVCuY
8b5+w+C/+dmJZT5tEs4QqLoy7z8JKPNSyOluqMQP3srdCEgoFmqsrpxgcUZXL5bt
DD/71NL9I5TH9eXfoH6N9JO89KQOeLUWxPI/Sc88xelTuHzMxwz0HAmlXIuNQsUy
pLuRQwGoqDElV3hONqkSn/rDLKXML55bbUzGrIyHknQfVKNwzvD3bIgVg+j0gkNF
NquMb/oosLM8F45ry628gY5L+KwO2qx4BZS/K4ffbnEtGU1aNAAIH7OX+rp0qnt1
/BPzaBDfNiQ2t0Pg7KoqkVjdm0I98dY/8Wwyy0bogKI=
`protect END_PROTECTED
