`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q8fAksZC+CLnZ8JzURH9RHgY4ufpG5RlvUb+Qw/CYDCFYUUqc3+vgnXKrc/2MHhz
bIzj/N71bJi/Z6IvBtP6gyjLk4ijV1ozksukcHYuxaPAieuO20mm7UrEFeJTEW+b
bWi9D+Ju8tKdX1kJAn/u/u0GBS8Ym4fHL85iCRIOSjVEJmqDFtKUC1qxuewaCk7M
0nE1sOGE6QfgMXxSQrVqBl7Nm+vy1u91gYbGDRJVnYsU+5MzVxUzLYdY7L9wUT/u
FqRha1bhNgFrszQUjzR/P8B64E0cK7Zyj851wtw3w0FBKtcy8BnESkzPf6O60I1W
+bmPDwrj98vUnwRg1I7rl62ljs4+CXTo2cqZnfilw2aHoh0iuoJ3t/bP6ONWSCva
AxLnt5IKwWF80T55BdIoM/1ujS1Bstg26LMSUhw38gd+wQVfKR09IL5KZ7i1DN+h
obbkGwKiI3TgJyKjOM/LUZvVDCayWCU4AnTFU/zLAfM=
`protect END_PROTECTED
