`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZoIjB4ITcz4Z9UUkA2Ztd963SYiUozwEDKZjnSST1mpeZh+S6jH4CsTLJU/SJ0I
IZm2f13oq/T8CBINnCHesgnWwKQnO47xsdZDNOXTk8cknn45Jx/C/3KCHM/V1AtQ
lMVTfCgSnoVQpQadB2ol5yF1j2vZsKw5fn3dkdV++BCEYxwBEojs8NromSv2F59h
lYYHn0LZDuaX16R0pSt2C4aL2kDVgQG1Npj9IpkWskT6wkBBX/kE3aEyeCE4R5qW
6L76X/wa4cKyajoKqbrrNscnlp14gTPUhpZPztHfxD5TVnDVVjOmXUM0/OIilm/3
dvs9Genhac1A+CQTwIW1VHzoi0LJhUfYO4+KPpRLcCtss6pgVQSiUe+IYm4RWDXW
ltudexoN0IGl1jjqrIgQyA3zmkM91xEvqJtet4y7OjFh5ht8de3okyAZJZcxpCQr
fiSdBdwpU/MmSpvMqdfRYxl433ps1Jun/qP8SXsTKk8kKwl2wvHyJEDYuZSS8djD
GB53kMLCPVY0Iky1Z0pivsjYjb7Ikb0u6yybqOebBu8qWRXvoq4VpDWJef2v795x
P0Gq+aXg13PUMM4E7MhTp7NttfwkyvZgNfuI9pCCd0P+TK9/Hh+P2X/ZpbNFHlWt
d7QlPSmGGq6VMd+bzNx/yuP/pbEWZ2u0ZS4IltcCyE/zBJte4CZHl+CeGPvVXSwH
kYJC9clHOyp86sJSCgS9/1OV/+uzbjP7X0XlOr5bjGVh5TjOvkjpBph91dhAk3Cj
EjgVbzc4Cvtjv8d2c8IFQol1d7IulFFxet3QhphJpKcSwJql5QZZjsEIxeD5KuXR
31v391uWprQTTRH3RHvrk01nThw5fqDMqyRVX3LWv96MQ8KUMraiBOjpvYrYm4SR
vTamiwCxgGdxK0ApFJIitO2Kt2w2FfKn1zOaxY29J6nW+C82gJ43fSmwFwqFkdjK
aZpn2L3EbueecYOedDCmCgs4sUocKkjzezb91Io0uyjmfZqD0pIkpbuO4OmNrVoO
7Ts7XEuFiJzcb0TuXVaE1hYNl+7/qtiI96v9UW4DLm8ZVHKvrDqBaHwAnl7h6BLa
WykuQxoSzWmSNxisaqWY+3Rs8sp2T9pcfl0Bw2X/7PrTBr9HnczDBuPUBXm8SMrO
+YRP1+Rb+wWgg5hDq0zJZykI1g89ASV3flFpfZQxyoprnpc9WJhU3gTePhOBV6zj
aI45627yYj6WgBlO/YRJdmcIST/FKbrxPK/7VU+rhM+gEHhPpiGw0Q9XNEvNu0fp
zDlamOujA+5iN81pc4QwFMwfbfDwBgfB5geNEOdCunpSTXgsAA+GhE3Ex3147GWR
T/bJeasQh/NS+9A9wywCdKvXZTU4lwtLckOmYpEqi/VZEWTwsi2uAvgvJiq6kV1B
f47f+34puamLptBCM/vpTXM1d9lWjK8S0D7JCOGpZb8HXl3LPw84tjIvAeQ2pIr6
7gytbrTm3u5IQ/u7C5fCx9BN9esx2+EI9htTrJQtHWvy1Ywb+9cVdW8BRauNWTCB
VNrN3RrCMnCNoJVRq2ydRUCdHntRbwyRq9akT6dArdaVJsVSjN5GLa8JAOv3pOB6
QHE9EsiptU9wEqk5au2NJIw1cK+Yb2GIxCc6412kSaNnv+HSCF6uePDEDVszp7G1
K5x5TDel0Uo6FsA98oKbJAdwNY1q9/50Hb+j2cZpd0dqJ58lPZ6dZYIXZ6/zv4uC
BuUiqReJ+pkbnifj32Nc1o2fA7xO3xmk8RKSI0Lr67WkazGFHTdCZexJn2GWA93M
Fdin+0OZe90qbLmaa5iHB1BxM9p9TleylckgIAL7gtM2w8ewTa2+zvAfMfbj4/py
YGiobF0pJ3nc5s+ZqqCsWek5jJVZDqbn9xCtFRr4Ofy6oWIq8ejSYoxoLkVZlTB/
Uy6ofcuTrZdqnL1biaq8aBgvXnpING9zUZTSlHgCcSmWOUgrGUjBRyyw2j9RVbtU
e3q+QFJJGH7AzpDGw0cZhbHnVdmESnBrcEyjAJVoNikEVdH3vr3m0VwtzX/k86I7
pcsXl3nuGX1L1Lt7Q2hSbFvQTKE6bJS63yM7zwCxdULchT4FonEzDeEqdGvckSLv
P0xT+W5UvLLe82k4AFxv4iBMmD9D3QOodMibTOpmEF3n0kZrgxFNumu8U8jiixCu
86b0ei/jq1Lckmdma/viftdat+xKlG8T9qaAshlvYmk8gSIlbyBaX6tL29/GxQjc
ZsUTLuN3Nnql0xQpooGrVGWEhelGDaLnFlKqjuSyTNZrQkdnuM0pVavMXjqRR2nM
4ohEJhiALj2abwiaBWlR+LajGBU76kkOamg6E04vIF70eoXYKPrBUQ18pnmjCc0t
s/mGpEoPtYq7sTbkVhq+IETJvNCZnqGrGOnsq1LktbM=
`protect END_PROTECTED
