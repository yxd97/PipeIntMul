`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+swN0LwtRmrjI3AXTVY/m9MHFaBoElPilu6DVV3gNo3Kfq7rENUkLp5g2Y3FgRx0
cSievc6sFo0TAT8gEk4zvPO1mMiP+tPUI7yegqm/RiYlzCoiqbANyrgOX/ahvdpO
tXBDN+clk+wJKOLFoeI5kp+lmqxKxU+ZLfNG5a3ZPHpDZr8xhzdCUicoLssQ+fQi
SyZe1ggaRlr8QBC4he3OCn0PFuprep1ze5gQSHVkb+muRsdLyA04v10JkJxFtk5W
lk9kq6kKN+n6iCkZ65+NOPZk7Z9U/iVNyTkGPKDLLB0=
`protect END_PROTECTED
