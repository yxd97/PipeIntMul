`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kRZ8v4CAjOe/nN8JPsA4zNgLSzafxjZE8LDh9Kbdi6Pyq0fzjTJDiLJGRXTBrsRy
6IOpEQJm+nXJnc050ROsqiTwv5fHax+YYrMM/jtZs7utBooUUYkvtTdH6ABSBgbL
kg9ZlR56RWoAAuUneNrmcmUtTd3uyWJ3zhJo2kit2fnJECIXTzvXeMDrUPY6n7qr
vQrQED2J0ewnbBYSYJZo+JSvFXvoZIdQLCteXH8YFwsDjxddL4sRc9rJl0+kNoSp
PQDfBVK5V84ZeNp08H3g5Apxjuc68I31TgFM5VaT0/XtuaFTFqHnOPLL1YzRYTEL
8RExWIn65jkpN9hcvQ28IFApSB8arGfh9yByJrvvbSVTBNBoieHQ4/xkACr6IzkD
34/si4NE2GkAxfuvkSgouuO0Vsz93+1omuovOvdWxUWjj9bSzwaRMv4Nb+IYTilc
`protect END_PROTECTED
