`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7nCGhtccR+RX/RL3HwltQa1pYEYePlShjTJxH/Xco0UYijjrCNJH5vZ5P7cQh7pZ
3O1FMrJ4x7Ve6+Fb3ZLfHSm8uP0G1vD9NogT9ZxIAxlMft5JtrVfVEQkaj/G2xAL
0ooTOUknQkk+bil+j0PF9wz2WHDcpF1u2KvXZ9n0uEI6X1EGvY5uXYTwM4TtXU8s
eHiP11PAMMcBoOgMy3a1ZpMqSsOFsAD7w8E8FpNhdJ2dxucA/K1Oji/R9kZGmg7a
jLsqeeUFDaUbdX5BECUg97TJq1gYXUQIYuWQahxt2qmKjszfvJclX6lHJLl47joS
7E4EZB7+RO0Nn6N34PfKyxExPr3UxLJQxaKjj64nkOPddxfSyByn99ROfI2iBXbA
L1/GiVodHw6ychhiexeYAGHWfIei+xHFIBlJ9vHIXHl3II2fjq8L8eb/tc4Dwc9C
V2uFWlsHuKmXKKgt75Teh10q4fujI5YPwePAFH20V6iIK8BVUyQ7JDWOObgB188g
WSDe9s+BrGS/0m9a5XI7wFWDRWKudWDQGD9kGfWbG1i219mJKNUamts2DBZkELNE
19kEcEXTzUA72HfSdV/cqw==
`protect END_PROTECTED
