`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mj4ylhfyjdVZ+RLSWypoZUsWe4Go8y+WqMrT316MSni7uqnaMlh8utvtyeDO7DfB
87CSNw98M2Oj0FMenO8y90uIwa/IEbRLfU0OLmj3CX2KLOsXQzpyNmCyG0N67lwN
8doXxRztLsEDUdMilMNBa32v8DC6K5afJtKdLPk2l18bj3dPr70PR7fqIarKSnur
R6Xx8CYOC+7wEbiccEbolKq+LlvvixaXqkXUBk3GRh+0MKN+XsI4lk6iHUE/ae6S
XLlYuwg5Y2h1f+asaUSB+LA+awYUstuaLS+nPFkTC4QfQMMHSCixUBg/MB/U1XjW
TUw+QXJm2VaYrN8l1w0tAg==
`protect END_PROTECTED
