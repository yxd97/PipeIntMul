`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rN9hwclT+d5n+dsL8eS00phw0enWyZbk1gYspsfotp5gQpGGlMhP76bIknfT8WD
oxab5KDI2EgVY9ejwpmwV16YOWwqajUDPntaJqCQMQZPSTS+3XkgrraRRSiWlui4
8MMixuCv9JOBkur4UVtShXq9RKiwHJOTGXy7DU1XwAozhi6xnWlHsF/bhRtdfH4n
mB3DNk7GG9wtq5ZpiNMTwEjDduPzeMy5GTC6z+v1N1qJhSsfWwuwi3CanvllhQw3
3hHGbce+iQ+eG1a2QVeXvy667oL+8v9hgzDhYjPnuHgb0o29/ReYWGC8ozIiPz+x
fiWBJDRVPbGAmgv3CCAOH4urKGVc8eSLuwBK0liRUWq7/+EPY7dxzmXjhZhAUgpA
rR9NEuKx1B6Zk2o9UdICizc0fHL8Sv+hh+G26dCCtSuAVCKC+L0OxTai8/ZmqAz3
+3lUQo6Wbyjw0nftEk0/REauYUNo3IoXfKQNJif8gZOQbHdVvdhgXV7kYTQlFVIj
1Z10YvHWzd17EM1TmsiIpwHjE5nGzMhE08P2lgmjpla4/JtkkNICYaAI1fYzEns3
f37cm/n/OeZBpy0HrxQ/eK4LdetQz5Xq5wBBLa13Z+oeP5Pb/y7cE8tfejJYmRk/
947/U/OyplXET5T+ETOQCFNs26HoDQd+ISkWgIcPsYmNZgjmXWYrNd2bs9axERwG
ksrOS0EJ+smsCA5cX/Pkmi1UzPy250Q4Qn4M+NDcYHoZCnGyuQPPwL0jRCTDJ3XP
+LAb5cioZuv5EHh+ryUIBzs0kGExGFRS1vEIl7zmhgrCM8yCbClR2ONq2JrMZ0RS
53zA4UmdMT9M65Anw7Ju7xzEzlIayKk75BU8h3f+Hs7cpDrW0XN+M0tPq7IZ3Gc2
3FW1QbNZu0PxfcnroTjyx/DM78R7PgDGBGFLHr+74o43JjX6UYoK7BUQpLaTGS3F
qMiJvow0GOQ8ml//P4PEIAhM8mh372QRRmaVNLz4YVIh3RQgpqjbaxMJuYLnmEJS
lrZgJYN1liaJRdFtTRPPcHTbZ6l2tFoWKgcX+TAS5SHLdIKvivg5W2LCLNs7FT7q
hYoGs4cHNu50RBYrq8CYSW2iI67pTTUjuOYNc5cC8bf5WooQNBl40Iv/78UGo9Xw
qv2/l/1N2CXIWGq2DAo5EkO+MNtsf0hdjB/OpUYL3+vDR7PyEjjVrPpSaVx/e2j5
ruszHzBGOWcrILIx/vHOEmSvob0OKI1i5twF9x1k17dRIqZL/b3M4F+7H+kfDZwk
zgQSjIHvWRKcoxwhUWupDxRHlwsimLr/iN78zfPTi1Cq6VjwXwoq8H8BNiyYck6d
8RDI/aoWoEj+7jfOugliAiTuM6RqGHi7UeZ/m+RoA15LGiDWSTouDoCt98Sr6crs
uhmFnBAldf8KyzOkXP3GmBRyUwN1GrLq4df1KURSp8kNSnZbJGZtwZzhxC2QOnkm
bVGvbjagHx7Zx1qkNSkLlakaU40DYl6ynEPUT2tfNyuF8oL6F3jzuITNWgb4SE/i
vottgoHNVNyTHB2QrzwoQzoyTi2t5x1JnunIVU/VhiqtOs23UosCHNvJTUv+VP+A
BXyqhnvWSouWhPKsz54kNt9r0WZHoy6jqu6ZVujELvJhGfZIKk9ana6X1+m7+Fzk
5KLrxHsyihUINfpukJRerRJLdvWiEdfp8ywbNBPHKRq+bGVk/LGwF/Q+ejqj4RDk
+6+LotBA3Kye8YkNJHg5+mYXjsxOfrR6bUFlJKkQA5cp4Bl1K8xMGYriBZhLxr6k
nVFT04D83HwZjG6JiTvHnbD2m2F6NqKBET5TxBobRdf1zO3UJ2DJd+TqiY7Mt+9P
clZ9VNqSnFh0I00Av+eK166j2/B5DFQ3DQ4KS2tVL0p4gxNEpQ1QmldFAx4xDjIF
bM4BrVO46WCQS0o+IFaxmnv5WcfkP/HjrHP5t0H24GGokbaPGR0QAtNmvVhL3t3x
6jk1YTw7N+mIqtzu/JGaLvpkQCPWn9SwDWu4REIZXDX06QS4k5Vj/X7qe4dwIr9d
RHLa92sqs4plcdM5zvdvcGP7olmqwroFZ7KVQd2eu8A6elUCnGsIRlenTahToqFm
aMA1mdBWdXgZ4Y0ecG/aN1r6q82M9SkwN7cXtsrl6DnwOgI3JJev/dec1VhmQmr6
rCYwYqzR6UEH+yf782PO5KSqrzsA6b35QzNqDlH3N5cmv8HduUQjotmOIFC+dAzH
GmCrmLhoV8+EIvh6YVCaK/0EBVFPDassSVAaUPY+uCaMiOhlX9d3JUIzyLoo64JN
HfFsjwts3gXZ/ycU4kxAymrhBaQoer8TTGZLijC8riSu0RJyHnm9+Sh8ImGqr/qL
L5rAljIEsP0znrKJHi4VSCIqdJvvQsP1jS3lyTfwBFQ9duximzA53MwrYc/DDou7
lQQg21KfyLupSI97W4bCir5bhnDDyuzTq3YnK4BlLUDJUrbIWCd03lj3AJY9SJSZ
Vrznli0zgSLksXXnKnCODzjuy8NZVECzDuZ8HO6iHdurNmSuVYSPK0uGnIGBPQLX
EfMdq4wSGps8ghKveAd05N4xQf2LbiVGlWQLxKhcgyatYe2ngvn9maAr9TB4DzoU
0Z+WK3QyGUqyo4mbn+TzbMNEi107Xrg9fT4xMbcyZcxJrrzfJ+FsqA01hKdAFC9C
ZlIt6ACMsqdsVLCttlaV5fG1ieBrjZNlezqr+ylAjg0X1UcD49jP0nc1RVMCcmEO
F9whoDCeqfz+PCnY6LZem4tAyxVFGcy2ivD2Js5asd5eCKHjOczPrj/ucDN/lfye
2s3S7RL8F1T4RfBN+BP8ldSDV4PHBgObwyLBmEkArCsGy7LitGlZ85ulV6+YV6O8
w6nk8Pgx48Tzok34m6zddMGBTCZeWY5ib4b06YnUO00KwVkyP9IG2LpumC3F101/
uUAC6pAb1OuT88Ct2fU/rmnqQOYKz93zh/TRtWh+a01ZwmiTYYTMd7PPj780MWew
n1tFnaquREcl4Dz5AQU71KHRdVG5nm7Q46bnz5ibgTqhVki6lH8KaIbGG6w4NDL8
i7lbyGQJbINk1yPDcUOHt8SB0+t+IidX3RWc/f8hDQ5eVzC8JVxTuNfOprEpHK2W
x6/hV5Eybwa66LApMH/s2MDm8m2M1nAX2Gc0z2lbfYurG/ok8+SbDH1eiiGUs6f3
qHO/Eu1C/jzt2cCgVxNBqUN0jvlcYdRvp/Ko+zFq2n592GxsMQsi1o0kAeSBUSjm
bcEFsNa6iMt3uNJgc4UJG3KXGf0yIDfLM/qbUCnpIhB8Mw6ZPShM+/OEm1EftTbV
wJTWf0+B70jTD/aNR1AOR3RD8dg1Jrnt9lD0ekXOVriv0+wlsCQ98SDQF/gJefEK
FyhB9JA4VmDFNCDyeCFrFkGxAYuQRVdB2TW/ymRxwThn1VEJeEacO0JHBuUWWEBp
KvAkYsaJH3IoZW3jmrIdboMeBz9T4Txxjn19QlwI5seSmRtWld0GrR7c3wquLvqW
ZSZObVeVpLjSdm06P5ruY1YbG79+4sL5dcYb58YzODEfXbKpBFgtbkNALNCx5y/2
KluAGdl7sQacFY7UvjC9bkCArZwE0VncE0AkHHUbcbF22p+q4Jb62NckS/LUitwL
/OIDEw9r6WRz1GnmHf6gZrDweC8mTjA5cgnt3l2auILGdyBb1DQQyCVGG2TCBild
f9U3Cnqg/II8k2LFkGMprRuNaGrBDalJlqD6lxlrg/R95JCKPGcoVemIKMVzIrDn
6yvIqaXq9Rw3w+Oxkr7Ucw==
`protect END_PROTECTED
