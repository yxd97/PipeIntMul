`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DimR2DUilVsSx7OdFkVEFLnPslMGqHpvWn69XFK7XIVBNPWXBnx3BYFPmumcN+vT
yvY0DGsAq0a1Lqu/4RkDy2+8LnZs8J0pRPgSvkThTwp1ct9hMJ5SaTsJ1m98OG0c
2oLf2KFnNxZG/Pr49ia+k5UcO6/tje59MKHtxXlGgoU9+CkTMwB5l0fHvq/w6lUG
JsfRGwLZ6vIIoosDivLvphe74ZFFUTM0mTiSUUx9LLvo7gdf+Iar6Pd0AU7zb6se
efClH9B5vQK5/xiOoMEczAw5ZN6MqVq9t4c+LcsFXhcMwlbaeq/v3zzV3X7s0bEa
pTgNsGUuh/nbL9NDplMgAZzf48z0J4fgCmfsAAISqgn+1xnNXM6ayRIB9YH5Esw3
b8qhoZgtbq3isxdmZ1SzTsyEKHKHR1tIHB1WWwqW3/q+m2BTASD6imJD38g6AI4m
6ES0ZkJ9w2XEyn4WLB+YE35aMnCL8PKN/w+Sk1wm8563MLbSSBq//Q5BNL4g/FwA
laqkkpr3Vl4DfVOXYALq183H++yT7SlyvBSKAEzsAiOYSd+McQCzVjLL6wLtGIqC
En79vOuTiqGItMS2sBVI6QEBCvfDVRh3zau9TGZUQd4D9dyT1C742ZLVHlxM4E7p
8x+WusRuiSEL+lJ2S9aMeWb5h1lhPcUAKlTPTU2cbd6ZI4OYrzhFlSYHtVkNYMh2
5zrMmj0WOG5erCvUgGYwF4Sd+dko4HUqr8T1foI9zvj03HFJFJMer4RiJZ+FJK+r
IeJY+T02N6bZp8H2LDb3PnEnvHYrRGYNYQv787PyBJA=
`protect END_PROTECTED
