`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/kSWZMrkl5AU8yuvlqZpCzJ2uMTFbYA9bv6bwGz6+yyNqQ0OVVLPBtlyqwdRbie
YPLMMWt7kD0AZPOYDC4H0n8OdPuCIgjwC8c0oUD/1u4dH51jhsFaLbHx3B10RDTv
qvtpOcsflN9u8K247fksdoqhpAdQHvWzI8BVTjBBMr451eafoI8chuEAvO3UZmhy
43b5oA8C1PkH+/37FSqiVFxYru+W/tLmg5UaTUZZx8uo3SVYZxxe0dhwjfPkFayD
lfMOJGuf6mzWe5tVZXEztCLYShVXO8nwmnpB2wYURCo=
`protect END_PROTECTED
