`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nT+gZqiucCrEPgKVs99S+ThJ0ZRDzh2up7V/kPSITyX4zEBT57VUkRGeBpe1ZfU8
GEBcznHFIffu0U4ZM0bb5eKjLgzATbkeIeru6HceGhcQo3dntHPJNDtDyTIs+HK0
Kl/c4UB/vhKNt2LwcWDB+I/kPw8y2laoXZi34VN/uF2vupLMdZGbWFi49vtGGBzU
cpZFurXsxK9ih1/EMh3Pp4A3SvML/Wbhp1t3KD5IcD6cLWna//YnjqFCdw3lQ9U+
SrEw/o+ZvW2Mw55Cp7aaa7g3TdhjAthN/V23kc0wDfS+jCa4nKUhlWWw/XnkOyNU
+Nb4aT52MHlURsg5+xtVHXfwozKX9xnFC2XDuLgG0gZ733Y4KUkHTSofMcvd4d/9
p8FylowBN8Q2g/cT5h963PAWhmlYKTOBvBxtAVF4NSS1DG5XXtUVQAQSHHdP+y1Y
hb6tnDYEIiGeVyjUcJUY4AxgG7K5FgKD4x4AWv6dtzXUTo+Na12tn2fDgNgEDq+F
5+xXHcc1uZyBc5fYhXd2yA==
`protect END_PROTECTED
