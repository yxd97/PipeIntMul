`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
22TbrHDaFRxfxpBmtAOhCAIEug7H4mSSDFvky/enb9ehEWZFM7tzVfS2SoqVURJp
vk1d8xenGqRTPGRPUb+NpP2LghtR1Q2XQdSC1MwwQKeV6SiofQqaBi8BAbR5Zwk9
hSBxVW2L4CCknpfscz2UtO7UD/fbWM73aq/v2bWlbYry732gXfLjqroVkm8G0vwF
aMcu29MEokgQIN+ErPhDV5m36PNpSuAx7W63411RQW16WBfrS262WjnTP0Bjr8gi
JDNAXuYgYad48trOJsT3DoCos1VfJNb7KfYJvlHKcvm+WO7n8k+veU/bXZjK3Fok
eA7Gzi8inDollHRfb30XGPWm4HUyuwaIbKQJvpnR364q+ZvWWDzBO+EkkiZwDSEh
RzCzmxXZUkqLXAPVBqmelq5C4d/qbHQeIzF4zZksRQNg3wFOt/4x0aQaXRh/fuuO
VMWPdI4TqkjSS5x/L2UXINOAY31mRlI0SAQGeCq17X2jrGTr66Oj/Fmoylhj5OPe
+KPA2rZtkdWA4w+i7H2T4IuzdA5JK6PkCu75I2Q5PdfEfD90Cv35hxBIAGlW0/VG
`protect END_PROTECTED
