`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJWT2bwGaEOB2GuN/+9pit1P5jnGAojW2DQZUxCBqWwa2Qp2RapJXUfKkCoqJYr9
7pOHS0GXWgtXl1gZLx+ZW/jySmKrKzvZY9dSXJFKcAVMVjqlDnBHrlz+hjK3xJb7
8rWB4S1a5tuChPJJhi7GTsZT4/ZFi3Kv/HFUTUiGIjByWEBYZAInHL7hjuCXvndM
Hm0KZseEMJOmh1qKvoryFsLpBwBOOh0KUUq2xwCmo6az4+v38TS5V02BJRToMgCG
FZIOSH65l3Xo5Erx3d3jRoXV+BSJQLKyy//HUa7QIasRvlNjF+SNvrX8xSA5r381
VgU8LKTbBlHj1hdF6iJYREMPk2e77av/+H/wOLVc6kaK8pm4YwjzXDkxc5pdhMHh
i0O6g1zqV9EypUp5Qx9AZJps5WEr5MrMdP1vDlfrSYjTZI6KwNFVkG/+BhaLiunE
90B+3YW944v8gXbkgZSWdWATwlcsZsLo4sjipNE4Yx+xON3vpBPjaV0Zg9wfCaga
+YkcdILU/EH8zjGWQEkplA==
`protect END_PROTECTED
