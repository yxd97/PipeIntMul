`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQZRkOZWd3B+o+QYKVGoe+NGCueTKPUJkqHJWN6nF6l9UUDlCd74gXpsy4CmfU8U
WqbYQUWOs66fpvsFcx99AuzYUqWjcHxgD/rSTbHIk+1Gc5mGCnGg7uw+zhjmZ93w
iEkpYrWSCVRcW80VJyv0qv7PQKzVB+AuEicgKy1o6i7qoIn5xvYtojU1zsQoms/3
GEm3rBt1Cu/g/6Att3DersNnxl2sDj/ohS28dqqbpe73QbQZiDuOoNCZPw4mT6vH
kU0kUMUcUtoQC5sjm5QaPaPnhwDEI133V3TTAYs+XSFrDKUY1pDRsxHpW6CAvYO1
0dH5mrMUE9kcWOBZFJfK5W7Nu9GtmVQonxB0psAcs1pNHfqEBnwJJZxF+CxWvUa1
J7GjCGyZl+1FSJHkzJN+ub5OyrhgTvp2wNvbqNg6qs/jLWhVxvqgjZfWf3aqlsK/
w4jFCVRrbUeKT5pYH7gxOeUwqRFJNzk97GoTWsmKZngXpVwdUA9tpCE/qIqAJxHJ
nx25Q5Pmp4CJfUtomJBZiH/8QRipzQ8hvR9TAXaABWsCwT9qrBYaEemWP+fUWYa5
WW+5ShiJBl8HQEHPgwmTwps++/lbpmj2pDlEdZrcOzhXN9AY0tEncb1U1jaNsmnI
ZmRoJKNGrL7mgzRUJByJHQ11daYzXiGmF9SaludBku8c61CRIxujXnghGTRoo4iE
iaJ4ULXlndGKdFZd4XlK7G30Cjn0t7chueZRNhJKTHM+M2hxwwUs20M5AJ1HQibA
`protect END_PROTECTED
