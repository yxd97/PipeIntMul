`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UbBrAi7lUbxn6/j9QM8T6q54VRXurjv1ZPnDmVk9bzUQ89Y4nDsNylFWit2jP4WF
1hURUko5gzWzhwoRH1zQdyEjEDy3gceBHBUn5qsbIq6jYe1r4AZa0fnVR5VOLUOT
JSArW/oRBT7AaNL4tTzCAM5uAmWOAzvdVc0mAmOdX3udJ8xDx3tH3Pt/QH12FHt9
oEGVUSx4zPx4TyjwfxSw/50Ul65QbxZZSWyMYJYZceUjW43ncH3nQBVVNDWQX1f7
4m0TL/e3jtWZH1slQFmShIUib/AWG4hzP69BtBmatN70HwWX38RynxizpmfojrNy
PWppwEarNoS4GnTrlLWC7XPw/XK7mJC9p1rJPgS8xBVzTqR4RnqvE/XeMj0Dvn6I
RoeSqUR6HLyaz88yELMksxfdfUHkvZMoYrXL4EgKZKVqii30zppDGvsJokDxoU98
DzS6OatwWi0FzYykChrXLwQvQUp34927Chg1gYpNf8MrWWtZowjpPMMcL6YkFR6q
EXJiwdMXoJZFUa5xh2h9pMA8nCAysIQV7ZhNJxJoU5J/Wz3CSSaKwn34FPQ59G4r
4VB3IpZuNdQ0928kmeKYTKfzrNFWv+cl8jsZ8+FX+Jw=
`protect END_PROTECTED
