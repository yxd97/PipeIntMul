`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CbKZc058SGKvoP/9Zkae6xZw8qgnPz7nGv5V/IAu9w488QuuO0e4KAdXpeYiIfUv
YWD2oEL2QZnUBAx9nxAuW2akQWfU3vVu9ro+uHH9p2rD/I4y/LeScZa0s2tgHeym
qjQe8QHUMCVx8r8N0pSCe8bDwZIQUqBOkTBD6TgHmz0bXXQwGgJ4E5f/Gv6ME4fp
mmAWOFxx5ymppkVCsll5OySZnYk1eSxssIoXI59+NliidIMgDWUThQMDZwp2ndDl
shrA9zoTK2vRYB4Bw4yhurCFP1cR7tZwJd8fmk4CXlmOEFN8cPmRvnTlx1q0vql0
Y6LPGAvYYGqLSAPykcmgiS/4DH8GuyoWXeEftU6HHZ4=
`protect END_PROTECTED
