`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZY9WVaC5x/m+FmqT4usiWzjHX/rSGuQujWb6HQ2FWC6DQpaPFgxux5PIfqOqOGiW
7Id03IU3ycwkRtfmcHgtJWhSRI5ktfES9vYY5gkbFbzhSDgEbanysed7brcBqSGv
/EVub8LzKwVCGkmRWPhX0HpuyGsqmXW70U+sh0OYj/t0JsIgPHJltyf7Ojang8L1
kGgl/MTO7z9eQTTcil0WpPolB6Dc9+MDUsrBbrA3h5o4nV4G2g7FsJIGZoXX+N/h
22GeoyHzjPpwW+Mjn06udYaim9X2hnqwt+PixS4KByHkPNYXP0073WBmwzplrZu/
cNI+ol+MNCn3j7a0vRP+1Rs704EVxZQhPgxWm3doLoSF6bQRpieAq686PvTTVkY7
+uBulliKAGsKuA+r7rpKbg==
`protect END_PROTECTED
