`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPjRgC5cy/U4O9v2RGyEl3mYp33t06sqX2DBHsYBXajgkibYsxouGPmaEDeJdVdF
TpclmVRf0BlGc9BlB4Q6nPeS8CHC+TE8kaIYihatMeystNoQLFhkvW7VSiM3/TyG
WjdXu1ceS2q3EvC2hkdE2b3SGczXa+jl6iEcHiCfvD0ZyKstDrxbdNaKi/biOiMx
Nl5KeqlCFcj2Fu+c7F4x7FwgMNPZJhC+W+ozm+nQZolWbWsC6aizuhhObLghr2eJ
gxyfhEsjq2rq1eYEL7VpevD29wB+VWiKVf7YjIgqFB0=
`protect END_PROTECTED
