`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TlaWhc0eDUSjONp39Dy+QHDneQLyn1j3eXN4EeNfxTMGFq4MPABmIV0P0lPRLzIt
++cYYkWBPOeoJt5SCO+BoEldgMbOdyNHhCO/eecrm1UNKjcewVZA+sewhFuPew0h
1JkaTNolFydNArraES17Psl/ln0h+HsKkQ9ZuIyczsyH6titWxX4P3DIr/CIkS5S
5VYPAhuchDhGILb6RIBeSEjoEfffDqA4qrlgK2z3b29TWkikXfJdaqK4HOL4Bl/h
BamANz0oYugbEujwwIC0BXAHSr+EScwaMfuYh852G74u8GG7Sn0SvrGHkOOjsFSA
yMZ5WFnPMjJV1BIwJeU787QNn82Dw6zVmOdsM+0BVP0cvgUPl/oPVRCj2thCDzn4
LePqWDfNl63IHmgffulBd9LQ8R+zq3UzjPkIyXyv42Ze3nPAHa4X86JV+0I0stAC
prlm8/iXE3+PKzkRkCab4A/aMuELEWQCcLlOqGzkKvnEdlB7MOK+655WFgpt8IeA
HhzibvLEXOkpnMiZXEMAZM+VzGQ/yyBIDtnGaHFkV9h6+7l3/BjRLUrPE/wSD34+
T/Yt9luAa5PXzILuEqdFMY1b1meILLMZuVc790mqH9DVmZHqvqDWmDMS2nAxolop
siymhJhVYU79LLeF4EcgLakaEIa76nN2Z9MdwGb+o6D76vfR7oRtqsHv86PsgQLY
eJs2HArzI9Nr/KjQgAA/5DvGKoCdgppZqsZcSrStFu89suWn3H9GZLrikH3p9xlA
3NIfs0I/08MUJ3Zoh8u2bymnBgQ3Onhtl32aa1uLRg8HrlWYxxje0DHmc9GnSx4s
9mzGup8fBD4TFt+C8SZukZfRnU9WERyx4fCTKNvI4IuzDeJFOflhTqkflhyKi14q
vO6iOG12rG/bNt50LbG+DRLfhnOC+473EUaAdNkzZehnvBmAc/INlTR2YuIHungq
XCNoLGCD5qGaSrR4iSuQWPLmqojSiZxbeHXKbWOTlRm9PWRiXo1Vr6fn+tlbFHCh
+1qdOYbtrELN8lcsS+YMBEs5HG++/KdTDRrvVdmt/xltwEa/F0tQlJmtnPUbrT1w
/UO4zODUOmWoV76L5pMPEfRd1bbKZUJ0KRVoqFKRqLlG/0taXYpdSJkZGzjt/Zd4
grtdwqG55Q8FVVX6NlKt2tEMO1xOQNT20BquNmREM6K6ljDfDl9OeEYJyb10RRFm
yAujCuzAseMWXahJQSqZtTAoaa2GjRmtK3DletSIKkh70AZD+ZC9o1GM06xmuRAG
lMeHxb/cTenq+v71U9y7dHoVQWe0cc0J+ykAbwA7aRyY8vpzrC/3EpOPzD/nXwZ2
uWN08dEo9DaWvu+K+9KJqsqJXLiN5pLOubRitg8FC8ikqs4RRi1gUYZYGS5EVjGB
BWX0jlRYBZ0ukRSWJPpA8B6Z0jBvS/Z2/QTfVEmE03w8Eks9noZKf+LDubHDJmIQ
e4D9YhhIrGkQZYB698P6MpjXV2jYDzqJCjXE0mMm6PYccGNVDDbPiRGLL3sw5MPF
Z74UvAS2Xg7uwrCoJsr/wPN7I7F+Of3uGvG5HvL4qfunhHGG6YVxqHoF786L+vPf
3UT3crWReUqvJOgW9KeifKozlkCEod91L9+fTiddWMIKeZDaHj/PK/YSyPjiI/Pw
TSVL2MO3SxVKwyVCzqM3oGMNkqNrnGFEXbIyunG7d4ipGRajlTc1lAKjYkYENnbf
CKBAcwfQCPciYtJYLswBAaKgiOfK3mBCu4dQ5v3xyoWya5fRp3kyvs8lNAEbaCwF
8HCc8VGrBrxPs1GGvxAoRbHyErW0rQPmeiHNG8M3a+03dtqmloTCNKJfp3fSfpzn
ORX8uGgJoNnndBshYA2x4K+RPVqatOx5kAE6l4C41gEXIWUMNpiF8PVd3yEpx46S
hG8ArKLcjMCVB80yiwkfE/+zhpQJRG/8NQ03cpvuFPPTYswFXPBISQFuJDFD6pqc
2BPbQvfOHuEAV1/vKX1TxQBxWmT9Wgibl/jng6tI74eORPxTOmP/KrLyHA34xaGX
mazSGdSN52vJrD3Y6V46KziouhRRIcMLKTTXvKPRrp4J4TVX8t4mItwRxDxoj4O2
INuTvYkgyiSABevDUrUsgEDAyyxne7o9jDc8z9CNtZ6/JGFgwwT2OURUQLimhZZm
WMDtoIUmUCxdANnmwAT5G5nonqIsRUxwoPYsfmwkAW4M0V8Po2UaTa7VNs5g92Tf
LjWQT/H7Ctcsa+/EKYod8hayPhlPT9XvvLF2Cp+ZdQnvTapNzBrULpnv1xZxl1U/
WhLCUHWeZP/V7djtv7rKiUkddpdY+yFK9Z2cVXJGU3RBkUVDRbt1WWsEBLAjhPlN
lKSJKrgYaXTBQdNmOMSF6auyKG3TrTlZJRcpTh1uTIk8B5EFerpDugjHn4nE+74x
rEdWdDCsSK9rTSwgjt6tZ83/b1nujhG36xf0/0AkUioCxAFgbycZeSJz3Jg1p6X5
5i9X9Z5naURpej6qZmEnnzGBWREvBCC2BAzKAS7bfzLfKxmmZg4sFk31IfCXVY0D
Y6B9bVJaXPa5KOnew23B+LDfkO27+0dzmDb8V7FI7swNGKkVXuNT5Apj0JSwhXuI
va2a6N2aAqgFratbIsR+LOwJ1AxjvxsC/6j4FTJiqhz95jRk35efuwudy2qKhbGH
L3aGE3XX0NVllrs/+5iAl9Z4NFZMtv3xg9naoV9o+UXFQUdfV8oMGz5l0JlMlEsY
bZiCiKnNWUJ6K0zO2xDLrO+YNS3K9wbt/SjBcxVszxKISPowVKTi0m7eKz4SHAcE
hZtCh8gl/1JW+xCy0d4F9dxOfG2N8Us0UYAX3ipECybd0loC5wgtZayTOVvy7nWG
VXqxIO2dl6bOyVAycQSuABbCmUVWxrjDIJXVSXUy+OH9rBhn60WYu+3bMpnwCftE
E3e8j6mEhewn4sbXJoJms4CiRJu19mqI1euotnU7rz5AiwZvjzPhlOQ4v6mWo0jE
11223HCNVh4/jD9HCqLLsgwz5ZDT25yZkkXan8eTL11xAsqg054ywouVS9Kx3PB/
qW7EAjz80XSTj0SeninWlyvE6mpWA4lbK+yt8MKsMPU=
`protect END_PROTECTED
