`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFNTpeMS1mWr1bOLwgy9R/yJKsRUDPGqJT0SeoarD0dUDx6XTYWKF6v1ISA+JH5q
BMSyHpwTj+UeF9idEfx5ra7swZBWuXQn7G+yFmsrz1x4Jip2czBQC2qvTaj7ugfh
U5/y3uK3TrJ+XJMuq57Xl6Tnv67c7upbI/VKrQV/xIrPx0AtgU4fdlHvxNkQD1qu
9vdiYFDez2WA95kKkHCDbAL1gQ+h32s1HefYyHYB/jtHVed08VLkl4V3R250mGEn
sNDekcLFeTpwd3//RbyMuPp1VEGbo6RIA3YIXVI/Xz8qLOyPDKM8BdUFj6bigp69
3fpRnZVsWXxdzcAvKYuvTy0d4qFHGg+Evwpt8pL5UyLsCJVUKlMvabIrozGspjYZ
mS1w0irdi1cpWffI5PP4WSrM0tAk4u1yrQg5ba0QpS5+jk0RptxCGU5wgkMuFcc4
VKTBqwH0na7SnIBrhe8npGvs3X4MCNZEwOyMQKeHy7SZKtzAFUxEX4FkCnrv+OIL
5LMoad0PZjuktVKqcFYWICzapxNTr+VTC2NDMNfLtH32Z2SkJxhvYUZKMTuTHNxm
7P0x2MZ3Oacrg8lj+ahS0+yVtg9H2AMA7lDgBZ9m5Kd8LOkYAqji2sLjsFLwvnt7
u3+ZTjxqO6hz5kloSv7R7tJRmqK5LQVwSLLdWBKghvZTRGReh8omoCSACKs2OHiB
/+Pr2HQwMfE1M6pRlWchiB+Vxyh9JuuqG3fiJo3hQOdquuJ8ZvclfKgKX6e9Ig7R
cyCSNss58DKgdsxoycjsnKlUYdDTT58KEd1ziDnv13FmCEUwGzOul8eH7SmZFltu
LBEzIUqSCisxmmvG4zRO1nke8fPvSNpshHbihEz1sckkUABCXhb3kJfZAQtZsl9o
C1Nbk0pTtKG3/Bi7M/3GK0odCVY9XWWUhxp0v2qY7LPl67g1U6q+bhlUvah3x/OJ
0BDCSYMzvOWEqKrl5z1pb0z1paM+m//1uCxa2l0PjKPwGjQslpdD74MeyoDKNvjX
vVEqV7sTgvH85jVYgfkcuXHLhTLXe3NY31m6h3w6rRPpW5QAaUAxwt79N9hf1ts1
jtieinLcW/0PZ/PuMirb9hn8qhsgwWYZhUrtpKxxUQ/FsWLqfOxoUFmvfr+lf1Vi
ZZxBwHHFZp/lzwZyrz6FJ+E72heksVhAXL/5fGo0IxtNqJggrsW6fv/m6qo9yi18
bl4pI4kGYQm+/rOzzYEw/A==
`protect END_PROTECTED
