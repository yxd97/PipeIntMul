`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DdKVBSpfw69ahMuWG4tHW3r5ZvFnj0tQ+U0P3lxhcWNQnU7svELHP+FfNr7tRvv
+qWpSCkJpnpf8PdqSnx0s0MZGpr5uWV+Db8tgAdpnej/kYFSQO0PBMGQBhOkdMhf
amaDF3gvAmSRH/k0Hnq7j9ssBOPLG20AstWs1cwRqsH1bW+0xYgztQuqXZh4cBFG
urP9+dokAwpvM/4+s2HSO7Xwok7yOCyHpYgVV+uze9HviXGe0RouDLEc5wBvoG4C
GOXtiyUMGjYq1mD6OZLOV7/tML3kYUNPDPjHOdpPVfQAOC9CFn0rjSNQ1s8rib2e
Z2YFBz6pq0mKqooOvp0J0Gd9SCos9qWd77qGfObsBpuMuhKBpO4Wa0SJWcGzCwD/
wl//k8GQoz90bewcNPMsEaUJIj4GIEhV1llea2tPgRICsAA2TKDBsEdo9FTN//LB
`protect END_PROTECTED
