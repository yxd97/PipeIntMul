`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwWBXX3kXpTh6GGeJ1NNjnvnEalnzDciIVm+h5TDzK/uEhxEwF6gRFTOlggt5+oo
9XOOOQQDS2a2l06rJLLSBUX7DDOH1ta05YgRChyWDX2VQIUguGpr1sisdYtO0YqC
cB7bvC+VCH8u/RKCWbrfLY0wS/GlPdaxsm6l9wOLhzgHwvJ7XrOQIyN5I2g2eQcp
meI4czNzJR8bRJpw+lnKzgJADbSCDHPT+tZ5cFyP6j/Fcr2z6zCB9s8xaCb0H4rT
G8P+uVSmWy7pZS90v8/W+SlNUtmNkTZh+K6HPyTvZrzOQrlcnk4O5OQvc31mbtqP
x2tfBb2hthkBYgfKRctd3WJUd7AhPrtWLdmtyjq6FaVLZ7rxagBDD8a1bOViaD2j
jps+ws86UbeDu+mwnvEKWg==
`protect END_PROTECTED
