`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVZiS17PD6xVlEpMgA5AI2NPMn2pxq6erN4PMYgeTL8lT5Yn/oT1Va4u8GRZmx3Y
nYRUVKTx9inGAW9mLtHb3QuSlwolZS0JF5nV/wgzUr/nA/bj5QfBLRohsnIyZrj+
Yd4fTQ8ohe2AQtePvAA+ozWHVRaUkfJHx0D+cZ+xbfHSIovKLPSJAAnajDap19P+
Tw8eBOaWo5tZC9/YtCe7l/0N9ONbdP5kjgJEIPl0jUH231qtklJug+YLR/hrKUJx
pkDlIgjsP/6uyPhjg6Zt5p/wfHLRZmqkIRBXT310tVed3fVpJZkUCIsjVqnocgA/
fW6NDrR4NBCxrjlY+Eg6FkA8ZgL/iUrlKOcS98GfS2g8Jbj1FyEiNoFqb7HpM2ws
wiPSggLSbQv62L6Zfoqjp14gru/O3f8AcESdohocsRJwTTSZjLWQXjrglo9t/snp
76sSvA9SspW2pIY/E//EV6R5hsuL8VzuPDWtBYpM3Qdy4F8zbZe35zsUomiD0aY7
FeQyNhQif5+8l19AWOd5D4Sk9kKxw6UgcAE8a/UmcnTJQ4cWx5mq0BYKsWlFLDmb
fS0NkZq1U+79F8jIM5gXQqOQiFdNNEdpJW2A7uYFfiTkit+Cazchgh/RZkQQKtjw
Ff/K6vwtBmXUjQ2l04h0JFHhzRIwGpnqVMZfiQVpuIm8JvlvHilsoTLXnrqBK0AZ
iHdFtEZ03etsOI3rcnt8KjqUmWtHBmMzytulpFApMT/bHc9qbDwLLWPd9y0BRH95
VKG+GwzDxiVWVlytpAMsBm5j1uQwVqEWGhM2T/9NNkpvEMvosayuU6SWo51Nl03+
D5nyVORVZAo/GnWHe8WhjlgHAOaDMzcVs6syiLEhCeCrh7CyHPWGZar+5exQJOgV
bIFHVmxVgwrlY6CvG7Zg4vXrkYYawXjgHRY6udZMhNGsg3K0uGf6JRMrzz+tS7ie
uxn6QF6FRrmBdvzAeYYiTuV1h2kzEAkC0s5vp5UE2hUPJldDCzti8yDCJETLwbVB
lfVNf4gSiAHd9zVeU5NKfvNp15Xh2L0OAqB7woTEyFffWuUSgZkuhdeJYIv1ebhi
B1kthHeSJkiBMbcItAGk6f2An/Lby3gGQUMjk3WmRtrbm6YDblZCtbbWO0V726hy
va5NCcypTK87AbpgFgNnzDUsdF6qONe45Oo08h6yC+Gsbb1UNBtTz/NFY/edI0QH
+QYLVRxhWA3GRXQfn7CUAM907pL9zX5feU0vmtaxRuf9cXzsSglANAWihR5zvfH/
eavB1sp/d9PGzHmznsZU7AkAF/cxk8b1rxAMOq8+qwcpRHnoGA21MCOkEli2PnqU
7kGO9Xb4PXcht6FEiicIWDC/qQuvJw2LqzB4C18Zh0zIz/fEJmfObRvQr5jVYb+h
c4O+Lq3DtsHqrgH+SKUgyPBSoEfoJWwwdegs3LNOxfZ03iF5rqOX3/nrpVNBvyv7
DOb5gOq0Km5V9B/trICJmE+anGz9b9KxEo3SBAREfg3m6vTt1eJRdzoCseba3DCB
GHfJXbP10R2O9T3TkQv+pNxrObOGkbmcimZGl+fGgsA/SCKzn4MIMSs+/mejRwUV
OcJCik6cWJMemOKT0yqXZwLm3bx9dhzxa7Bhe6F+w6cyBbv8Osijy9yI4US8mSTs
BnnZDLEF8Yn0qTTmK2o2chrEHrecilJ86ERz1xVlzn1Sb8sO6OSbdT33piTvPL+U
H4aoXbh0IkT9pIdZ5yrp8vHZZ2av8E0dbgRfOCwKPzB4Er3sJfhV8k8hKDoQl4h0
fLg1vzvcERHlEx8E/KsRybKm2KHFdNhz+V7EY1mOEPhut+yCcWx3WmKWazNy31TZ
p4b88NlU9EtFUCEkzY5pR/wUqaxlMnI5Y0uNyjTPmrvXcV0C+7OjaZIXu7f3yzGZ
xf4mequxYqXTQ8Epxqe+PwgOxgZFa5xVweipaCMGLHstMhies5/P3h81rpGC49i6
TpgJQRdTWwLrlEFo1leKgDWp+qWmkmZy+aUG6N70HLmko/mSimP+ad1b4JX7KGNX
cP20a+qGaUw5h/8RIiiclMCawaILzHAxy57QLNFq7vPWbN6KR56ej/bA49cM1AAv
7QZIrBFsx5t8vCe8N3GiGDTRSKzgR2bS/eNht+Cy5I0+RSw7rE+b9Mqb+5CzSO3c
sz0T3B+RO3N73ZdBeVx3ZWLybFF47TcYBsbISyLJmE4Ycjey01HUEziULwVP4Pw8
c2audx3zQFh8LgMg9y62B+QcNhljcnFtf8hnfYdF0DtJU2i3gnXKkuoaPryh8OUA
8sllbmqQqAiyuqPURtZu7IabIH2KOJqfzoB0cUgE2iufH1vN3ZoKRT6vI3N/XN0F
jsWQUqb4D1CIxfvgFGFPwiyBjDN2tT9dNEFd/iAA2iRyNNJl8X56op087VGHVQoq
saf/DBOLRZnVyZ0N9NQ1Ho0YZl1qwNjO7nLbW+yMSznF0mK1kcy6jGNfAyPW7s+q
Bl6UUthLgsYlhMiqAi8h/7FNZ5fMcNSM7M00taOt6seoAIB5F9HidL6VXf87pWSO
kZl2o//aIh9308jAQ/S8SQybXV2hU/FVk3Nt9VpW4GmWKdOkd/eIN+0QyMtHnhuX
2fLbEcR3hWrz6e0i6Iq7gnRDWcKF0TO0XicSQ3pkEZWbuBy4K813eIYM/BuYX/iW
r/Vz7snQzFfYpgGPAsKIPvkzdx0OYR6fmom+qR+xrwF9SUvoT82Km/6tPiuxFCWW
XBx1tRgvOqV56wVF6iIchTNs39K7guxCrksOoW6SskCM23rWF7p1NucVZ8gLIKbg
wLvzLm6npUiXdykMPJEKniUY39VchlGKQUW1AC/G0rISnDKiEbIlYnQKYdyuauRf
jHRjfAMBnv7r3xYUyEODHsQPJmfsHFa9a8nAcnT4yMYDhT9I0m8K12IRRMk8qdbq
93m63Vw0XmsxHkh7mcEa5cK1ojMKm/VqFx+v1Gk98a3MJHhtbWgzFRvTDPph8aot
Vrb9GVTDUUI7SJ4bYIkSdWqf5JVicaJRcPJ4bAkfwfjli38eXwgLa9NNxpbpEQ11
qTh8maGYVdcONFGB3uqjU3zaIAf48YTHfdTjCM1r+8mQCxobu20y1lmataZjgV76
QeyxtYmNQvz7MmU4NYKITSt1qyKuIK/T/w4SJMG3yURKwV7s/HbK9qxDzlWxfMdg
puLFUx0chpI78RTkl4XDDxhV0wXiQObkDtSIH6Na6hL4ljRn4qQedhsoBY9jVPVX
7nTJBKQ7H6nSmtbaz4smobF/B4oWt0OpcXW5W4QFGB8LJpB4ekH90ZP88NxT2Mog
z4PMld7vAhRGW5FNJqJq236hM9yhGzwJIfv+MESa1yeqJTtdoYdbhd/rZx0M7Wyy
jz7jE5SH76ekBOtIWOo3oQoz1V0DHpK75JgGoD1lSAli87PUy2wPKt+kWzNGNMdt
V/rChhl3sM6oQH5JUamTN6imUMkiP3XrPDtPSPfipAJM/ukFVsnqI37u6xfi7+xS
XGZda7DEYUfZPwqBw26YDOXhlefMnFEFT3oU4ayf3lskFkUkuUt4/lef7KEfO0rn
Vkdovk+BAwGQrYk4vSqt9QY9Mpqk0oQdtQqqr6KLTcOAn8Ky0FwjgsZWrjPCOYmI
zMFE4723Nf99OtuE6hu26WzdGNhMLdt6hsOy/xGc2dxn+KEyq+VRpxjfsUxn5Hs9
yLbfc0SdRQrPjIE6JpNjxEXTeTjOOhU0Sk96LrdI/nYqxvgZO6DAMwe+cAKQeZLU
lJLsZaZPZ4c49LDiJi8SzyHEoMZdIscskbAmLBsDv9KTsxy5ENjcBCn3wbYVSPHS
38Nhn6BQwo+F56m5UpklHoq2f/9a5WSEmX6ef71OU422kbutQbT7P0n+lG1DJH/1
Bj4gWL3N17nbDu4YMY3lBrJz/YVpVYmMkPTVn7mCjyPy9mRjctLAayq0laOdXFS+
YEcr92/VL3nRlMGf0XcAwtDQHu1iZ90g9hkqSOThLptysop7J6tFRwKKZD1d8OFk
rYStSdcWgiJSMEbo5oRSyxcspUJVFmFNFMBWc78aFgklIYy2sZQTYsZGzJpNmcrf
isSDPjnO+3bffRzkrQxJMkwSWx5S/Esv+aln4k+S6nqX9i3DywyciQF3Siebi5YZ
ub9ieGf2IUvxdr8UIzvOIGZrRdmYgrKTl+00LAr+NW9J8JKcs5dNtAPGGKnPHsaS
xf2R7DiqPkzrBCZge2CLER4JrE1oSOiGR8FkwT1gLHTVyheqIvM97OElt2lmIAHw
rgoUftK7uyDhLBFxK1fg/3Sv2+j+TBl/SjzVlYpQSR3Q7swmXT7hUlL29Z8V6+gf
Rk0dOnmnSCdvI0D60mA0HN+Zfm/YBicEJTV/IFpHaTBI/BKMcP9MJn4zixTc9ydX
Of/RzpN3Bxp/O2RWfjX734WWnrxoH6iWoXGoLRgJsyg71vFgjBfx7qEpiFuDz4CH
MvOa0luetNV/6Bt7/l284A==
`protect END_PROTECTED
