`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gm0MkPzPB3KYEFFDLe45cP0L1wuhDcq72uXi3Z4Ngew401BMFkow+KLnA6gud3Zf
OOocPCfQtTqTpXmESMSM8xzUXc6YS6tgBBZytAbYPfARFNwoGPFl/p9++RZ/BsSa
yFPZ2E9K0TFIB54ALlyFs4LYnkXcHCIeccNHfjLDi43jGxLsn0y7f5rK9UUy4aHN
/ZNLdYM4n18LpA78a7tElLQwFcJqRCnsRCBqZag0WMokYagdK62wo8YRkGcvArs7
UkeAD2Jhp2iFEZjXXPP2yjLB7Mnnm/yMvUq8rCUHTULiLm2Hd+pEExZEs+MM6vtg
mlnagDkOlJKcPvJ0Mzk7jg==
`protect END_PROTECTED
