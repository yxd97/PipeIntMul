`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1ziD43dxOxgPca0rJK8ejTFe3hzIE1lpE47toV6jMU+ex1JQ5M0Ukck+jQCzpok
OSIkPrvUVW9UBrcuO+p2Asug5tMwc/IUufWU8lRmtNSP6mr7mvUJ50JW/6FkXh8V
GJ4vNrgUfSoPVHOXdi3S83ZEOqg8p/WEfAuNARLIDAZRHiTf6aUcGbdOPaounf7/
OA99J00dS0OGFYnq+U0FZwb1oZ1NUgYXKLzJv3LBYr7+C0If0u4GyWojs6gaGdrL
BwStjVl+vrm9oiuOgnUj4cSy9zhDE2BqpzbM4V4ydSH341DGaZkQcLSUSmJKQKZJ
8Zax6kOriNt02m11h56BsRWM1QZvw0dha4PAl8YC36kNy0VqwFKl78D0OaHBAjuW
vc3fiTUSNoWUTAi0MvCMSOdzyW1xaMxWF45C3hzyNwS7Vb3hQgfWdWmMnaey1QHd
377nRI+oTlAYo5l8ox+RfG0t5VKrLzYjjvCTzfs34+tv9L7UMC5bQJrXV/twJ3eW
VQ5kAELQW3Ou9SG7bZ+kJtNAa6E3hS07mtu2Z6y6r6QFghWoQZX++Ouz/L1BYPF1
UzrVBwHPQRL5mlqty6FCc4Vqsl24xU+u8ByHwudJCXrQuWyQrQ3cfB7QsPKOrmpD
gLCgqS7Bj5J6oK6oWgtEuOUS6873k6rFr62tJY47UVwIImdeAsS89PVbtmys4tY9
0olWbx7KNF6FJ1XPK8wzvwRI4E+KP+8lZ0QujBZaN2pLt2536rXCH6FwvOcIio/G
/f9Ii6Bd3lAc2ZCog5/HmjZzuFbOTsCn6OL1nTgaVBqtz1/p1Z2WUvDPJ2SnCzeJ
QYGdQvHVKEQ5xn70O3wiE4Jb74uIOMzmZn2MR0JqscZvo5cKQfeL976X1UrTB4HQ
rkAFuBeStr12spwjXgdFsSrdAgo5zG03IpFa+we28WMTWPy3soha+ifqkFP6Fvq1
BtBCuPA2KCuDU6jt6Xwq21/eCB6LRaFlUsPoS1RDVFicIP+r7OrTm2B/fFppz4l5
nL+UhQbFlLDFBZPgx6xOKFvC9b0VqGnngdDwd0Z4hq0DQOI7iliHkogAnmu/nnZI
lbD7HZsGAeEVNrIwCxuUUM54gZWsAU0+zHMRaaIA02dI634eujokXpfGX85iCWmc
9tTqvoN+bPKyd1VfyU5DVYXIHCfjoXqFMm8vIemnFzx8qjO2SZOAysrb7n29TM4j
KDw56LW5v/cEarOrhM9LwZaIez4WwzHMSEzKwc4O6q0zZ/Q/9LPepGd1CyDdkFST
Im0fw0gGKf8JvCPGZCjY1YDD/WAJcU95fd5XWi0Dhdc+kyfIuGg5Y8gJmLFcuREB
W4599GeP5i2cGxHq8nmq31pLyQFIXHKMqTIMHCbqP8m4D26HhMU1S42oG785cq8B
U9S8K7DSo7v6rp0/39Fgkf/0eueyQmd+4zcGGyhEYyMlrIrGJ1pnqwnSKVKScezL
vk1UadMvnAXtBIxC1EgQej/QD9Hv9U2B/Uhw1bU97in28ppUNAuU9aaPmZero8AJ
7JBrk+nxN1Y9js3upPbn98XiTQtLdQ7gsPtQAivB2TfiI2EBxZdTXWi9wLF5+2zy
vvg1TFvHu5cqeA5Jsslmueqoy6G+HdGw1bNu1VFMmL6YaoinPoeXCjEwWwN7GS9k
pen1ag72U5kwj6NIibPptWkc6ntgMcFvGbc+sYa/Ehx+G8Oa2p34ydz06Znay/Z1
NDJ8ewo6NK6meuFM0EAgRg/EmjLLfdSqiUiPhJH5PLzjZOKC1n77+02qsGM93ol0
wGAZZq99HIr5aAE7hqDELRzS/RvCAVHhkojtj1YQami7TjUqirY7bDnTt+39GgGZ
2QdkRP6nuPgtfVeVXvZ0JfODF42ZXxvV8moGbjzU9pCMkFUofMuIbFMprAm7QyaA
/nY07IGEq22EKjivE+iItwVZQHo/6Y6jmosCSTww35TelQhRCe1z5hhdj1RpUfCG
+JOxnluc2ZAa60daBYHTA8Pc+uZ9YcC2MiHVNNNwugkr8K3vBlZTKommbvGXWG0y
/meiZoqeeqUr4HRpivkkt0vgr2WoZrpgmtHqtyJcioNqaS7CW+vduZGvzvEFJmYQ
NSBVPqOzONNDYaJeRihZiZV/KChb+aDab1uwcmBiUINY883+tprvuQy7C0Sqddd9
MP5NKaOXp50HuyrXzdza5LCR/uho2qsnWWkc5JhMYNoSDRSB4GERO0hFw948dMF9
hSmRKk7T4vCK1oMiaDH1oPzodqTVt5cmreDAU1IpabmQYZf0VhUDuJEr+Ap3okfI
B3igrtPeA+0vIN7rzKbUuDneyVAsc36GMHmY73a1tD5pxkMhu3DJF0GZ76uNsD+k
NzLY49VGhmni6D2pw2OMIqUiewEN7dbGsn2uXSGTcDs5I2h+Yu431D3+mUM7mBg5
LGM1ntjYukkxSnWhQmdbKVPjqckceTsZtwv4Z60htr7pIHQxvBQo1fDTpzMyLlzm
C3uy2AJXULy+D7Xq8MIUQ3pcOL/C/iLlcl7pMY8FaZRE73p1k7Sbr5cgAb1JYo+B
lMe6zQ8pSlCclR6lnnOOWTMyZ5ZCtNp7YcAEGujWOgbHbHFUTqJNWwRR4Ep3x82p
etxQUL+oKD4Z4HS1EqhwTqFL6y3yCbv9sNDpQRtGwddO6+qLy4ArymmDtKzL9Jk1
DvJtft6tHFxo0RHUbrcS0g==
`protect END_PROTECTED
