`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfyRYiu9snhOfWX47dh+s2rfLnlRe/y/+oVukpaMft89thm0vNFEK0UlqLpMDR+5
pMbKnLK+1zEvZcx4ZVl4wexvheb+6pMIe5KoumHXgzWMaP+nUxMvHT+UYyUKwCCM
6fis4xuS8i0iLFUlhCPxCi9/ufHxC0iyIT5qirpW2FgMgIYOXxWHdaH1dy2m1Tx2
TiznIDN2uPoJIhVts87gV3m/A+kSihK5+SdB9+4Bt8D1JBv1Pk+dFQVpXPiyvI1U
3sj2R9n+1DzrDBAdsEgLYSCVyXFSJb/FxoLr+6f41mLuU4DeDMxnSuEEispRhR46
8z0XQGywcIsVdydyIl04nF0HHBKtJ2xMCM6es95Ofk6bsD+iB3UrNR2ebYIE0JOV
OyqurNjV4TXtf8TonGeQJhzucZUzFiRLGdssSE11rRUuNSbm1W/+fIfinUc2oRnS
nlovzjCxuERApuHR+z8lVCWQhvlPXbX17ODTJjr3vksbPdJ5wjOOWf2QeS8Vqnop
exyoJwR0io+RD+k5A50E1C6MONTG0GyGtdCdloXX2KwVAQL4NXnv21BmZOR1mLc/
EJumUtze9YKZfp5LSCSY71aCxo7TV+grYOTgZ8tnRIhebZRQ3vNmMvLfh6I4paDX
98pd4AusamMCZ+CMd2mVxJg+IwGXWk6qz+C4/Wd+BHLzoLVIRQuu8NP/2eXfhMLJ
2pPHYoHR5jMguYouWVPlXMjylgoswy/UiYmEZPhlRIImx7b/GVxYf6awbg7Gcd2i
g0se3oMgdHQ2T41kw7FLtJhbHXl1M8pkzHZNg9C7cMrpp46QGkNQYBeMslYG9mxl
di9tmhpeqwdvFv4kFK0Gbwbm/UjWT+ncNqh3AnvTlJ4=
`protect END_PROTECTED
