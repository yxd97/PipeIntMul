`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/QRJN/WlDGkDmAPeODbh6TQVIxOfEcDIGHmpudPLArlRD9mwJlj0Kme6yVbhQ5wt
fbgytvsDqFogsbt1yvzDGJMOD+Y4moJaSvd40HaVlaPgqsIVMoJ8/2J+KaTV2alC
4HTRbMqyVeTyM20Pc6RpEAZ9fjS60DfIXw2FtcPTZuDbIiSnQMJwyA+Jbv8XGM4A
dfzCOXCExfrsObxYh7kFkSJfk+dzY/hVJc0uM5Evg9YU2DqAD997OtoMZEBiTxUq
tjl14TtzRVWnWM1MOkp/SJ0mWmlRz5naglS4Ghnv1Xpymo68b9oiZfvfrs95N/Oa
UDPh65+YndZxSCKbXPth66cpGQyTGLDzAL9OtrfOjyGV+kbALKSReoG9QXtN+sVa
bTJdNx8p9oPYBvrAHziGjqCUOr3S4CWm7fbgIP6AJCvrzmyQ/Cy3K1cQT+0p5Hsd
tDszn4odRALEbOyzst96i9fCpSh+CI6oWxcC32CUy4a4deB/q6kTP3tQ8CRDJlqJ
vnwBPHIbmq1skiUUXnZTjfEeUSMeQ3foAi5Amo/uWTr7KJnUgMFVOqLLOd4gVTKL
`protect END_PROTECTED
