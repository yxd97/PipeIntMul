`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YBPzm4gfcA2nrnwX7Lpq4E1k6qisgjwzLEnuMYBjDl81HfVBAFd4LYoLbZp5b3L
y9eRsgafWUIz67as+I7adoSRVhujsUbgimawJvM4u7tcIoal4bMC5ttCulznCrmv
d1luupRsXkH5HB+aCEqiHy31tiBRZ+pCsJIyIQEL5WjpvzWLSxIHWCzCE4iFuOKB
majx/AlTs0pgI0ymXpCHUFXlb0A4TDDD7utGPn69RxasRNWCA2Gb/inFx2xK4iPF
K3Shf7PQ27Ysa68gFrrBJn7w5dVHMt6NQ/5G/+yjkNTa1BM6FDPJ7vzhF2sfGpqN
803ggWcC6QNKZ8Zojx0FuspdSgd07zhontWlV2PP2gzgxE+r4SF/gGnsIb6wOZkg
7GdsqB2CPv7oKg/CwWRdSGY1eHyJXGebB3D+yu0iXAjh/Us9U86JII7eBNJ6StAN
VriilsXIpRJYx18VXeWoWGb7KvTQUzy6yokJ6xM8PiWTOlaI7UBNhHZ/CfQeyQ5T
AXsPjjU7aGfP95EWD/DP7mbsCTErfSqDipMZMzlgwZhAvufnKSAMktXWFbbVnmGf
rTiX0xFmmBPL8YwaoF2vrJ3l/rF2ov6i9Otb0dyVXjHvZpHFv6jk6gPQFgf97pdw
X+o5qIgYkZFKTxxqecGEEofM0zYrXsZjg6QFVF6ygsJPb8OPfa+SDs0T2CCFtL1x
5SHIMsy1fFAY9p43A8pTJ6L9Nd/28fcXQUqJyXqwe8GTAgXUmf3oZQ2xPYidyt1G
QortHwiXrJMkkEEbQcUnmviqXGJATg4+ihOHNmtNxY5rCIedrGlY/ZQ9kw0Sf2kI
1PnOlTPTOATM1s+dH6ZQfwByq/MWOa3NOPPAttRpPr+5niuGpNPntezLvWBP3D4P
5nq5ANXgqOVYn/h/kPSWUC+bkNu//vWhZ37ukc0wsFdZihqwUPPxa49xYi012/fv
Tno8GHSG6gxFGuYODMmHmhN/K0KKK+p1JpDpTjLNGxT+MRWz6OHljPzphoVcyOkQ
6y2hkoGRdt9yfSMcyOyfyEjjuu2Sh4xcMOInSr10P7lFnT01JanJltnXyrvAYa33
QokyVEXNkjwhZ6q6xEGz/EFAiPEb7w04UI1YSX0NlyCb1mFLDCDQt6hY8TBw2Mqy
CGnYpCosxUkxm2WOxmM50WAGquY48d15T5dRyA96mAFkFgd3ewPKB34wev7ewU9G
A3F/szzxzn6FSZPSfQGWGRtmtM+LD7bb1L3fbDMC6HI04u8TatTG0ulich9vO9y4
dQBPKRnxtTsM8AokLOkXIXsNlFOMwXm1I/VqYXgRGexMbiDqie/hfnBoRQ0ImE1r
pUN/2m37GqGRD3YSzwJhiFXMBaqwrDc4mVZmxeVwAbBtdWroNOCjU1mnct5G8tGC
5LCgtxCvziGDZI+nqv7+Ql5FrX4PqxJcTBPb4HZrbWnzdU+R2WrcaSgdtmFSm0by
Y7vVA3gWjAZUUUTSkCFBonVwcMV+6W2/RI1s/QmsMHmoYRyPLiHNP4WraSNROlyf
+MJcV6oLwP6py6cyqOGgLePDL/dgFGJ9ayDggkn/QslmN0wlOtJ6L17EZBEgDnk1
7bxJZy0Fl+ncBOItIPHlzZxqSbsbQwduDcJMwiAs7APqjtrw2vu9KG40Ct+2stPw
JElisjcdpw9F6jfDtgYCBZihnIgDHldhdrk/X4Pp2HEr8jw5UG1MAO9uynw8o9FL
s4JaQ4T/TvreDXff1haATfUZnKhYWQKcKxZetUJH2FTCjg8+CL2NSoabCFjaHCDI
u7Vqn7PJBpwqkINLkKPdywD7R05hJJfUAnJEsiQezZCSV+hSwfY8vwvLwyFi5XNS
xRLdbgUgJokf585U0Sfv2xpMrBSqgC6k7zo1WczD2KTp/kAUB8AXE9lmG9cx6CJ0
DMhSkr9Txyb8ezadjVGy/Fn1z9WBjjIRKBhUhfBaLgKZb7pyMK4QutZSqsGelXHg
UuGH/hMdWTQVe5H33Oxm0NFSDltQFuU6NEifM/UxVY3x6MFOi49SwnPAjrELqLya
Cp62vVdp7tJH7Qf1Eh3rDOiQ1vq53SYYhQDmzjed8iWbgGDlIGfp+HXAoCeCxIbp
Ks0yfzvfJ4+TNmZbUbomPQwAhYOt9bRiqDV771kgoRXan/Jz3y7oBnv5VpUMbtfY
mJEYRCg+eDDVp401AjdUm6YNXc6d0Z26iMnAwGIzRf1gThgK6wjMy+Yyuj0SOa5F
3GvUpIgpXNVAUlY2Kd/tJ5mmQf87Lef92CRUhyzp893uxGORrnwABuHMq4r9lfIA
q+C8LbS3etkFvIifEKNYjqajcrxbuLu2uYhXxzW3FWVv/OPdLJo+WkyCIUhMHIhk
VuICWJmeGRv9jCeFgzxZusHWxAfM0rBt+MleMRHg6aucWvjBt3I9rWwl3t2dabsQ
5haZgUxSUAHm7vAI6Tcpo7SyaT2IvESBojInCoiDPuYkyV+NrFzOZlFEbhhl3d0B
5RuhJoLeAbBx8M0pKgfHRT8s/m+KWZcaKz/C84ljhrR4wgHsG1dUQUN7snOQfVLA
8LhWE4z7V6kAC2KNGrvF27/vAJcxzQWb0RaqNXtDwyZqxZQi9sL7MnPMvk6h19QO
dkzrH0i5U0Bukt9jE/WGfgHUW1HcgA8z19sWvPelRrS0hl8/Covz4KbFmpAPupwA
uIc2UO+CRBuZ5Wgqc4kMgX1zl9CaLIigXoxLPxdr2Vly144YL8gV9H/IfhCVT1XM
JvxVwPncc3avfbiwtK4txDmKh65dh3KrfGz2lP8Td3+A/L/TpI8bAMH9ES1Yapvf
YvXxZ4Ch8xhHFBF9GSw7Ip1Hina5btTRBoHKMiXg7MueMihzSYGAkgdXy2fne0sB
aTuJp9f9IEsjujwnVltUpyFssMRhxXHlWSH/YgnT2Pb6tpM46FpuK09fqdtEhnlE
HRdqEQPxYU59nXL5D8z/U/Adn/aaFyrhXflfhdGNx3wc4hQlt01mnNRqT3E0uccx
qIGEMc4dMTlwnBxaqBlYiosq8sVlYQUAHz3gSdeWqZnvxRBssq1IwUxR3jLrz/6V
L7anAIFNuZ8pi7rUQWlkNBfyNmxPjFQv1U0NP9NLQ8dqbPvFXTepr0pjlhDkAy+6
XHsH9VxoxqJqDkILLENacmbbVqOMHJfnvtnpBC1EW/Ep431uyB87p0EI36eEaib8
MLfZkEWAuYwhiMBSu987Ox9aGpsSoRsYVxcgEio+oxXpKZZPw6At08JhH16mepFr
QgBn9TWWR5/5pCgYArMFKsj+irfZ2PTo+HMt7tbddYWSXHPLYPrDZYdImpEXbC68
qZw3NmWBthmVZyMo85/tcQ0E2CEiAyBLULx6kFN0HaG846BIZHs8OYnlrtTNTe6J
uSnsCU0/2ESM86M61838Dl6t/CUbyRWuii1G5PD6BS1ttnQd4kzJpX3ivRBGo092
g6JQHI20E4bxl2YxPnPUAufwxKrSoyYTvBTWGNBcfB+K81ldcXFa7/95LkMB6bef
YGAFfX0h2WOzkuHnjSto+Y01zKwYtp3Bx3Muwn7ic+80rQ2Obn832nU9CCCPa5YY
WkTS7pzSSP8JpT2iOvCiePNIB5Lb5Izh+RKtO5CdW79DfBS7dD9CrJ2r1Opb1BV1
Pkc3HYMyKC+9sFc2f8xpgFBl3yBKKNXL7fLgrhJJfmpqWCJCRggCP/Tefd3ehRPu
bxIF92d/zO/Izc5sYqNPuvZHEt5jHDtK/AfmLVOidVJkKcWmcRxkWc/kK/K1juIj
BRZDNfaZqV1Nv9r+3dNTs7Ecd2WHPaEoEdGsFXqRKEmX8gStB0aNThJCmFxJnOLp
U096fsv54ToAENj7gWjDIVCuRymIvXx2j4b/7xvDZrq8FhduKm0fWZ3nIxGe6O+z
pFBaDY8ShtOq7vlwObr7XCztnDp1H7BGAct+eItIWaoTuWKDum0rY7IAnPUyZiqp
ycLLKE/DgDPvNgvUu17EPyTPvDsr+hq18afIkTsONnjP3AX/CipEOeif6ZUqkQlX
9TZNNJLdcUsmvaxaMYY6jJu4pDq+N5FJfxl/bKtfjJKUrZZ9fRrBcRatOhq0NOHO
ZIbzYX2nO4CLkOxrKqamIA9Bra9jbv7WalUGAcXde/XfODHhpma4KhfxSzShvUB7
0ylv6mPpUfux+Dsr6w45mrMc+3Nso5Q4zQ7Pydcyg/pkPgkZhJHBCh93lHLhyVo3
jWUvbMkaIONBMdBBvnGjBHtoSvLU/oDb6KFY8wqo5rcu/v8fn6Ctr8m7PsZTpBPF
NzbNQH2B0IusiXjXAJ5a+YlqyjONinzXi2083ZaKjBc=
`protect END_PROTECTED
