`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DAw9zDcPDWkTzukx2gFVpgczR3TvLRtpqPzkiXFKt6uCRE8WkGQri5ZckcTJFXed
BFpKWJqTW5HzpPrDcSyiy4uJIIuqICMlbv23W4HzCLZK+v1bytrdeJC6s3jcjUzU
j4F4plKhbKYhEwKPv7qkJiCbMBopMZj9REVhmjKaQrqehcLnPbWJ8T7O0CRpj5vv
oeUAp6luOKTfcsYUYhqOE7Ci3SiWDBmnNgoVcdpdbV4RN029Lj0GVhtnwytgciil
iQrHTRT6Asrw3LA02jl7ya9cB0PRlc7FJz7w00t32Q1ibLkan+Usf/YFu8LFH3vp
x06mpknANZWWaKi7Bp5W4KcJMkHmpN8kLTSHvDKjMPwvBTiJ8OZGi3/elLiZuXU3
7q38HAh98+dDGrwta5AlYAqh1JlEaaw5ndP3L6IZDsw+ofLPF4HXEDLtvzmy0XSe
SIpN0ZSTwMVXTFaujjbTwKfA9oCHr5eUKUXc4OwRNCdpkvR+TuF8AdNle/++ojBx
TdENK+/2DclI1hPh9xEu3w7cE3MLqXq+T91o1UWL9edIc2VbewomxQxrpn01LKPk
z+BIZ1RQ0mJEzn/mbuNjEG4gwsMY8oT0Dvnab1crD341p/pejYAHfrpBnkTmbM7Y
VIthhneOjHz7gkvq4K3kBwOTGPPX6VRXjQ8vVQGh744=
`protect END_PROTECTED
