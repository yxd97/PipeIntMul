`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e1icslhshxL16kqXn1ZOtyuh/6uyQ/K0qONJk8KHukhout9k6whSE86O/mEocYob
arWOzc6RL/n/oMIGdUBaKfjKgz6qX40CuBS56+uPw0fNdaFVbZOOMYibSK/60zzE
XRG8HsEN93RxfnHXIw5Zk2qroSRUawepsU6J4p2FupiXP0f7rTITog4qR9Qh/Ec4
eoxzsGqPx4XmNsNbP3fFOUfK/GNwFeg0ROGAGsDJwTGyRl/+gDAsnk1Y6AxybKvS
MkmS8F3wALacfTNbo9gc/WYQeFEPhTXrHncgtH501zPkFXAJfIN6ibL44QczboZi
kZWxBznP8ib88Xdck1lmGuVIxlcl0TQziy8Z1BeehHLz+VA4hv57NnDpuSntELFr
/V/gMMEwYzshE9fbuvJKQtkfYGEIjFbOc1lT12Vz2op6WLY4Uz11+xbqMXpVIz60
yJhlZb6EhcJaQb/JyN6Eqrc5UNdfgrrPad6FgPTkExYpeeeEKyDS1ZoOF60xyTuX
`protect END_PROTECTED
