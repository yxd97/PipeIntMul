`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJCQhYLf70FulTTIgkyhwwtbdlfWzVaWIHzmIouZpqVaEJQRTH1uSG5hjrrac+26
NmTkppCqy36j+R6UrFWm1KxYMmJ+OUz49pz2MdxOOFfm6kwNbAvB9MEDD+gCYoey
hvzssSOodTkVN5Xxh+8fuOnXlst05YhoaUEsRGqvGuGUlyGskvmhdHvK9PYoxqdJ
eiMVB3jqwek/swoATpT0Agu4eaEWcQErxBLwiGac4H1FhyGstdfr2iuJ765+Hi13
oe/GQkBHTl21BO7ZbW0GSZVJbndWJD+1o7UmGEvapPhkNZ7ppMkhRBiPOvbaXg43
zp0VOsVSqyaSx807T13e7Fd7C44oVzCVw0psrDT9lzKnHN/xtna0vrGH5iLBgkIZ
Lb+C2zIW0ZigviGusROeFlmJ5mWvyirxMXRt+3wiELGT1oWwgDaR7t/WJ4Lx3jY1
WoC1AwMDBos/Hit65yNYo4mVPhnFWkTa2S8n4ORdyKMaNNKOJ5BKBOafLsvbbFxv
31yDVSTXt8upHRDcHrkVXDOUV46Ej4wURz40EjAvujY+Vg0aksY8cH8uUETphBvY
3HsgAFrfDDBWBucc1HwNIBMmHSeoGamrwkG4M8+6Ughhokvi6/ik9xVIhV1ukNs2
vqsnchyiUeKSsIuNxy6o8D3p1ZYQx16wiIl2A/MyaewM7E8fg6yuoKrx4Rzi6rv7
VOftJtHwdnefF88RxQQ1bNWHl6ohwE2hm2ejANhh0rYVEt1GxX3nYlq6inJ7AvYx
0oPGsB3VhmrVree0UhyNspdWXkJJCKwu8Z/s+sbo0PvUL7nUIbtK2Q0xZaEhoYAw
i42T0tlqpmqmKx7O/C8t4COlbOjwKyYNdTSSgop/AbkP6vEtD3m694fp1o8aStOV
iyhJT+prfM/3ySSWANibDLgtzBrR9S8hB9WwwjeldSeGDTUX2F7P+1Ec/+CqivtZ
y6jr/qapYMBeDuPXdzkX1QUYGgsagbHvYhXV4FeyQeuTqv4uewjl7a9oSHwJbBsN
iUw2SzSxhLv+yaEq0YcbsbI0C88Z+UHt3WapTLauWEDlXYJhOQ6DanepTDIDsV9G
EzV0PBHFX0FiLMAzg1sk7lwjPkKAXT902BLINBVStVcwG+QXn7qXHkbtYiV7K+82
cMG76YVMaHYqlKSuJZgwbI8S5Cq9xnIhdK4NLfTUUpUDzZtf72z0ucGho+L6Nec/
KAQE1WcgorVfvjpEXtycmXR+twBy0jRdzOzIleAgE7I3Z62tE2iP68VEqkoxeQKc
/bzBZsSu/T86l8D+nWysr/MqJRgzA3rPBM/gjvYX09W4Aj/7lUxaJgEsnR2/8Hwm
+snz6URUQqh6WCpSAr2uzHJNXLhBEOzRRiXMj9OxpiLFcMr+ksEBxnt2IzvUZQYN
+KpJvEaiHpM8zMVPP8T3qZ5yncmEFAko++wQnAeCIi0+MJbyfZGV3UJJdjrzJ7ED
b8XFbA4FoOe3AAFmqYzcDF3pvWgAhaQ2I/mXFkIyMkAUmSfSI3uU+nnj1PvULDww
ocEXFwoHaJZDEejnI+cR7tjZfgHtJz2aXm7xKrWwYjxbKN4e4dOyrixGFAofIs6e
lNZmhvO1EzsrijDIkXQAd2WmcHkxIz5pQt9ssZX0a832JLVQVkhuXsC315MadF0H
WyZszKjsFI+Cp4kbvPz9AaniGHmvKk71k55W8BhUJUDqWNuCzy+psyj1354UCEU+
IDopnrPlyIKuldeqBl7ZKjyg9ytaemHy+9IOyGCr9x++iT0Gkn5jsU/nFF953Mqn
n1UmL/l3gRZAoVgnzADK4t2OW4fbdcgm/yvwD/gPayfnNwJqtfmq+nbL/L6t0IPL
x4OHUllwVQIf7Ja618dslVCdTH5DbsraI+SFmAJRSlf/DPWY+q8186gHhrEuPsH8
u+6g6s4G0XTTScyqRf1StDhZdJZ0qaQ7o/TuThhagQxfK8yf6FPTN0uW+dAejfAc
hu4MC6WyAOMqN4GJY4CX7XqAUipiVS7elKwidKkCbvrnqDRHJAJNndqmyM7+t5oN
e3u8/KWLjy0coIcT1yYViQ==
`protect END_PROTECTED
