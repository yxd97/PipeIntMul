`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqAzaH8+4RpiaMWDVNn+XO/SRmqpvPCbIc3DD93CaRtFesQFVy6zFmjJkubzy8fX
PP6DzRVRd70GC4b3j0PptrQb6BAcnmGDLntYZU0KlCDggN5n4iwi8Hmym4PdKWNR
JCt1Az2IIv40aqArcRAbKeSuP3tKelf1zl4HyPfksoltFutJrkCBs/dZBq/KTlIO
RhI8iwFtDFMIP+pbPV0gzFwzzdxKHA3VAGIfe778nOv1vv0Wek9CevFP7v0HwSCq
yTQBgoCuYYxunQUlb+9YyQHPTdcNJ7BxQ92zAf/dmdPzK7foPaDMU0t52Q/RLSSk
r71hoWZgpkuwk4A69hyXFwPgOii8tOYK4hhfMAfF+HWhh7r3BGWAxpODKadha3X8
teNC9ztJG0PerkvpNg1G9/nrLNDdh7Xj3WeoH7IYVHiUkOyc7D1nJ61pOYaWZI+I
lh++FKjTW9Iy29wSzTQTl8hgNnh2MG5Ibnk/fAD0+/TnXD7kmOvi888KOyalt0aP
wK+53m3ckaNR+2qfQJ7rIFFW+20y7op5vsbL42LcuGMj45BjVN7jJ/wPXXnWApHV
Jqng1Sl7YOyrem4oS5Lp28iJbtI0btgdrzI7fSORvPc6OITvBUL8C0ENxQciJlB0
hcW3LuGosTzBPk3wnjxRHyOXqWF2Ey4dIdgAenITmNiSJ3MbbvzegoyiT6arMbYI
YdoBVvrA0tJuvh2mfCPVC9ANz9d/QbtOHP8dNZX3b9vK27CzuYhqqr/00Pm+1R5n
+tMq6VgtJRcNdDpvr0gT/16r7k+4ZL8DkQmMt/5kaAZ5EGDtlI8bQAjKcnkhALGL
r5SKX+BwWQtNnyOBMf4JbA8yXDz3pDsu44jYnof4MxlC2M5Heaa3+jK3fJsVqeQX
Fk0BkHSfpsFByzkhSUBBGM2TevqvIqkVjTadJ/625egPMbvtrOk4sGa2uSmvnDIH
Q9H36Nd+sAy5BgS7kBKc6f0eRymJ4w54Wml7cqPKoW1tIiXUuVIg+W7bawA/p8Wn
34PpeZwjnpVIReGjB0RIumPVVZVeR8guG+EtBEBqPvkEIps94iGJdmm4fEjipyHs
zm+FBb+m6ziJiQFRBdR3p1rN1bNK/P8QeWYSZb/E7w8ktu/WWXccgFrN8g3Hptu7
N4ZWZ8kmfmtbwchVQIb6x/B0YtUPLh6N9dV/Hd/Saj3auA6ZEFQzOeW9PFjuFObR
Fem0Pwdl3nK/ILarvhHua0ZRjZ3tKgnYMgXouuRCK1ieI505T1yHUV6udkDCJZ61
ppDvEPIyj0bo2Kq9hB+xNGPsX7gs8a1Eapg+3kPcWo+S0WeNjEUexP9iS4Afh5dO
OADeFH8AjmVSG9xGh7ArrHqwtVZxVPrtBcw+NjpMB2KF6+kUi4Gg0En5IUtN++YV
o+2+SfoabEtrIG2Tmzccd2C9RF4R/QqDkadVLQJmKaB9m3/YKCPStunWou+nQlJE
Pap9/xBnQCCjHkzLrsCq357QRiL5Um6ZplMmAkCCP082bgzpoF/mSWqLvRbER/DI
sanqBapnE//oNBJynikFMpC8BGzjVqF3yw+IwvRvU8PCyfX3rXVw3LhTEkfbS13M
O8Fvl8Ox5xwew+KirV3w92EkO4ZId6UJjxOq+8dCAH4xPq+570sqRsD309tKtH9q
oab1mZF6HJlLXynGYl3wLfrPguBCXdB+cTKzD03crYSU/0Su0OmSocBaIm6ohZLo
e6f9t5dsOyBx/SiXxX0KPR8gDa+2EZQa6EOLL7HjoYH8Pc4LPpZpEP4wQk0oVUOm
TdzXnZfsN7su3DcozCXKz78XyNre1W8T8NF6zHQemH1p0IKlvX6cyosox5KB9t4j
B7ikQxfVr+13pz1lnbRsIf90XxgblrE06Y6nARyrCAYm0TWckIdsuPEoPQcBnN1e
viTr3z6x0HZTypv5dPKb3HnkNaHZ1qNQwL+IhvukCtmRbgvOMJ8EmFvy/yI56H3w
EdLf9o3W1p0nIee+ycUNv9TeMRGOAhEL2GFRaQYk204IuYFxrgbAhPUyRpGz2+p4
wGUlrSNbpM9BTkQC7VLpVxJXwNrmIdLMT4d53N9DF89JvBqTdyOX8orAKK3eiSva
87HxYyewoPZZYZ6y9RBDbPearfYauT79o9CtMaLduzGRUaGAlHSaWPR3PoZ4eBBj
zJtRnIo+envGVMlQAjlwsPkSLj2OgbnmPv38X/yYxQcNS2h5TuMG2wpFxjT82BaQ
MDIWyHsKGDR6RewKMEywD3VuOdcdvvDQWt91tey28S43G/5jJdCfOa8HHTX1PMLN
Cw4a6IgdHZ1vb7R+/9XUWE/4VefnsULnMKoRFlOlO0+pNX7oKm8C/Iye98DPKFA+
Y/QIzfRrYf8UeZj/eOdFNdLEJEKBvii/aWIjGPFmiDf8XIQIam0pDZdHb3We7pSc
rQfePmWV3tV+XvrNSvFXVpnW4aBn4d4QAxEQb1OvKD6/NZs2Fk9FPCAnPdxwXq9m
ZxWEyaM7fU+vZq7KHGjzb3PHzHPssbBySsHRTJ8DZP8jNaXcyakVPiXf+UwvNbPO
kVoJBTDj1cPBdT4uOuLKaHHYoRmMcz7mRRVcPEPLtPa7ccN5xPOO3mtznr3FhqwY
EicLGAXAOF292R/Ut1L6ntDUkSDfsImwn1h2jV+lxpGujNB/rbBsA54Q9KM9dGD/
zPlmaTIyER+pam+3DQT927zH8UpiBNQHXE/YlAXP5syYv+NvgcVc4xMrJuK/IPTn
AS9tNTz3mTJd8c6a9pL0Pln+pGZ/Wv5987iMsDRIhLfY52ngcZjpDSPEtADwm0DT
3g9L2QPP82/jNr9b7VVFFZmZIzp8YjpjtVSlmVNgHG8sGDfluegnDEJlX/vsufw9
gjnkiKqfgiz12dr7yHNzEhxdCrXEa97BBYwO1FLycl+M0L1wA1TgwWyoRG9cFWfq
KVg7IHREuzTvh7A7+nMFCuzaCWH4RDj7RtBTez7QtLuNiA++eDKiGCw8s8Piy4aK
zZr0+vJ9T1R1jG6JLpZIXFMX17tzRR/OEK9xvoKA05/WP++wkf9snZ1Q36DIN0Ml
bjKZNoqZJ4xcEN1R0Lb4waVmVy1wT1H2UDhUxjgQ1ef91U2erbFnnXW4uLQCJYdO
gNkiqOAhFXULP0Mckjg2dk494mP82fpKJAVlpHzObVITxyq0/EhtoQU73D7OLbBR
xsD0B/dTxb1LdRlmMxcriTSYQYSFitMQKDQ9Hoy5E6mUrW51AnOtYXawcAXPkMwy
Ft8g0J2M0Ru9vz7uSZ7zhdraI0J+U12eTQU9DTr3zcyBtmk4lHvAAfBW6VndKFIf
3WOHutQH/FRLivFG4kD4/jf12crFkiKpDCZfBQhB4eOpbFLtWCLH/4xFhVn3csze
eNEkmvkS+DU6Gf+D/d4n8vdzwWnYCvK85fcY6Rk/lZen5LD6wZ0nM5e3ETeHPbi3
5jjkwIqkuiLt3zHQPHx9ErwbZAHudCj3Vr61cGUr2Qc=
`protect END_PROTECTED
