`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b+DfrJE+xFcdtSGbJJ8c44UUbjZX2c96CtsDzdw2zIBe8O16IBYaQfGxoOe7cMgU
vr3wGzHM5jxl9jMnfFM2coy5eOG4vh+121FxAfcHI1iGdLev0PqoIFp2XVHHlwpS
n41T5te7oObaq2NcCPiZ+uXX3WInqGcZE+pjRDFpFKhzEG64Pn7Y7a1Hi3PYLG+A
ik6vX5pgbqx8FS3rJFCVCRKlqzW4S55t0d12k5IJjk6G5NktDZ2YJYZt1N0Pjv6W
XauaUHHzy0zyKh4jDgle8LP3nDEpI1mHX1FnXS/rN1Y9eyjNVmUcyRMiHmn6a81a
TZssGqJ1NUnR//lT+CyrL7WPH/ECNjDhLivs9qBgtlqpVKSWsSpm/agZ0mUU/kkD
GpyiU6ogsa8FDs2+1DIezw9zwLc54EtPW458tZR7MDNO7rUmpijoMy2HnwKvjZ3O
`protect END_PROTECTED
