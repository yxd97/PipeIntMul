`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuPAtYAYAnJ9AjFVsDuWKdgiEWQPK+sHDgc+I0aJYDQWNo7V8tlRu4Ig49IXwpLg
zH8oAcOZIFLaaMlENIxVc4/9OT0zl3Yy3FVEPf9N0/mxm/US8ZwJ7FU95J9/nDBI
O66CTdCMMOaVDokNt1ALzQpCclO8+hbdjcDes9WBirlb3PU6hqxNWPEt6sp0H8L1
2c+pIEC71JuuzO8cmaOoJUKlGOrjDeqlT0rp3SukXQQ4nPOFR16L47W8QZyNJnXy
p6GMW82F90WeE/cohm8eQWxpSUoRr/VQLulqNuPjobgFdXml4QTLe8EeFwJjQhZ7
6gqb5God9yrabQhjPnNKcK+q37jvKn3H/OjbZjOJgfVI1aRNBHg9QBTsLjmnJvTQ
tbxAR5n5YxtcuhzZwlWHhRb4BohYwwTYHd1fysbnvXvHakumXVVir5f9BjZvF26m
Nx363pLXyCjazxqi2YbrFZ8g4ZWvizVvZ0RuEnivcfZbWf5TKDJiGwnSDN0HPiHj
H3+N69Pch5jVTcTQZjLT75B1vy5IDG4Zsmr0qBBCp2PNvae/5hBtJXJb/Qe8Okie
VCn9Fwyk8OaHdygIXN6x7a2T5PRR+uT14HwGV+W4tQg1meQkZXUlKYd23Lz2kudV
ok/Qm3UWdWH9NklKxfUucSThIsODr/5uQ4xSl8Yxqhk=
`protect END_PROTECTED
