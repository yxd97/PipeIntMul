`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2wDYjKxpJg1226XgoZUkjrKhVcVeK5q/izYP/eHLE2qt1UAuXyhRrtEPrYyiRy4A
OwD2oBR2VWyV2wpEZM/INvtHg3EOGr+SC6wTTRGBBNeWkGN20LK4DUegKrZQ1BOH
ybIZXk9+Qihp/20zXZvgmHOAOTnK51XkaB6pU0i8HSLX7OxieyHVAkB3NAAwR9c6
iyE+dmrZqC2FN2irm8rvYFO9zUChYQpQUQPY5ZWKfoddN5jROaH/1ZSYxenjIur3
9T6Rj+8GLuvXznefC9SIDPUSiiESTktbePsa9x7/VyrqjmUAgdj4+coFiv/SdUBa
VWo+sxMR1gW+PI7jbjIj9vp6VFe8zWN63TlBFO96YwqTAoUqGJKBBthhCT2SJnVy
CZjNeWIdUmnYfv9TaHjDXZAc8Qda2rzbdpPtpVmF9vrM9MgFvb/d/QEQt03FoCfE
XTf58bHf4FYYLzHRBcy9qCrO4wwYqv3JPvT8gwigsW0nr2HuzOxO2V/mDie+bwsl
baOvU5vlGpIchr2VaVmSFbiWFs+Bt0gnFEW0ZGwlb14tQCXnXAF9JwIAvimUDJ7X
T5xXbHBrYO80dYNJtEX6fyNE36HSC9lGzwcHeH+o4728wCXhaNSdHaU5ySGG35Kg
Tzs1xJdh/T93qmtZLm2Tmyk4mnX7O/wqPinflgTnvc+cjWHMuoGpPm6BpYHMz79g
eSyV2W3wdCsAmx5c4egTWFVa0P6raAJLKD/ct6APPyonaROvMbr4Gf79N4XPxVVR
3bOF2L3zjpWG1r0U9s5tj5E/Y54ZyBV15Iv7muXul/p6XtiI+hDeFZsJ9UCe7cbd
QrmZESq0HgYNVj8Z4/JjvlKihRutKLaVnha/0bUpGljHuvjRLdQRGrLwG+GuZMKv
HsNJ30a/hmTWxdpsATTD5+B+dlw81nCEM4N5DeWtEXUJRlqUiaLE3wjyPoaa0TSa
5H+iWzc0TqvxMGHU6XbZxg==
`protect END_PROTECTED
