`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZNiuh8mLAY+7+owiamxWZX3+ZWiIyi1Voyq05NKB4e1k01TJW4jmg4BaYJX+IQ/n
X6mScGOvaPaK/HOUqzavi/y+sLc7zSdTuMybQMWz7/MWNOTVvwyNSxIcePRZb1W1
qoiswyFmHTqOqr+Sxr2BVSaXlxl85zW0xRD3zSY7x04nUSV5Gw6g4jg3YBZArSmA
NSCWJR8ltn00XKoODeSoCu9xdWTZzoSCLxrCK9fLXK+zx6a06spDHHatSMzG6iq9
t0cVSdSY4eh+cOzFjAzJ9V6VPJtoiNnoeTtaHPVgEnkvDebN947Lj5llxxzTzBbK
9K/S8vnajS3ss/0y6GfgslkZj5lXlf0xXbUE1IA6eMTY0bhim00grrV1sHeat1CZ
fyz2FErD+FZPXUTex5pci63pOAIitJwOWXUEeHtWt/fZlkbOUo5Hlgev9+MLtVEp
aCcjNSUpsx0at3jc4YoeUCyMCXVv+qzJkXIw35tut/CNtErsF8CQ0iKe3/iDqHw2
wUD3UNciJ41GdA/3vpF3+HNebCIYmaJRdxzx4R3rJoZ8CL0qBN7cNCETxbaMdNDq
ZCe6zL2DIyTStzMUpSsUU+wXOKKYv2x8H8fitRCV9+k=
`protect END_PROTECTED
