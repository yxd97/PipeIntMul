`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/v010dgWCf4La/CwRxGjD4GTaWxZRw+MwzdhrM1ZKZCDsFIrAAl4YqupM37e8jwT
G/DXpqTeT2PeEDaFC1lycBp7F0acVYQGUZ6Ww1M2DNvarxh29GjIxFXhvrsQM3yA
AxCqE/Se/Gux+tziwfQlVq9dvNTpsX+xntC8Gy8yaa8OoFat7Oi/7H3/5xYM+4H+
hDZ4bcTFKfyZBxCW9vJQRaUoAxl2uTylf6BdMFxVnVjfhO+kGxnAkI8zXWrPtd3o
8LinVA0tMIWSdIedIrgV/wUJ//u9XvX/NKok/A8CGjrnyNzBD3qz/pgZ8sKx26tc
ZnutzB0AIa5Qur7h1o9yg1oYlVl4Kg2VnduXGvfm0UOi53axiW/Xujn3JKSd+Dlz
2hzwwHayY161fAGpceYRmdwAxnmXfBRe1MiuR0Iyc55b5N+TsUfeWL+j+4SPrnqQ
LFLsPSlB7Hqijvru+JVCmbcquu6VbXY9d0BdqhJZlRGnSmrvxJ5fBApdl2t4lQUS
tyW3ApTfdF3RewRRnHfN0qmEBzq3fFLeB7/ZTEfJp3m8dxioXvmCiSN3o00x2dUZ
XJebCkgsR1OJucV6QXGDDJF9tIsY1DMf+fXng3zQHnx13w4LAGdyXod5q/MPuEGg
doCivyUOivmp157ILOnwyEJdoOsMufUwyDWLZi36oU4dzQ/i3Z/sLNDHD+ZfAjNE
pXQCgzt7J6x1gxQz/A8B+E3i0yt2sE1WERkZyHaaIBJFlBhiObYIuN34LHGqzjtF
Fe3kSO9CksFXqTAMjm9jb0SkivGEBeJN8qEY4ohtm+vo9Og8Jxih8ldoeIY/RFrl
NUtOJmXCr158OcaYTi8t6Kzsye15UgtgeAtO/JKO2io+U7Ompi4jQzzff/zHiWVO
GCPCilhHoAeXO2LILWdutqH7kG2IB2/Gce3Mc4hAp1dxMjnjSsPbwfc/+8nevQzv
rxTzOhu8uUvGh9Dp7LbE2sEfhew+uvDhwjBGQPSBuMFFeyDJ4ePflYd/s2Ey88+d
bt/Ix0AeIlvmq98Jzd2sYlHAxPowzurCpCZpf0BJo2idqq3uPO08lmWyYEaIcAQS
Om9JskxvJVn+TmSozhmFJpMJ0fZvhZGT2/2BTi+YSjo7Y4RuPsi6/Ddrfg4sxhdm
HZAko6YB2PfRgixFl6G68wndalPoWKSa5ipFkM8Ni327M4MLKsPQw2Qax9KmFo4N
iuuOwQT/mcFaSBSDCuOHqOV/5uwejSYTz3y7DYDhlXXBy0K/DqiQO8kG3R18u/Fm
SYtrlw+52MRcegc8rkgxquAJ1cK+ImcLJwnsfnoG2RfkU46xYnENnzGmUqZFc6d5
emKuPmGUtwWPmal19D7GJk1wh9Po0ubQnIg3Mt16TEmWlPD9C9Rq+T6bXshbNZud
V1754wIOWuA24Yv3+UDrBaXWZa310M0zY7QZKf5GZsd6wRJxzuFaNH1Eq+XbAujA
BHhTQ+/oQn6eHpm5c08iO+PPDabGsweH5A60jn/2YttJflExBPNa+8HdKJGXPn6e
2pivzs8TyTVbQz52IYgC5M1Oiq3mUtMTlK0c2Mdnn3Mw21TlY4YsJNDQvrmZdyFH
5rB1Ujlm8CNt8W2CoRx4Sw3d5QEZBzdYXFuGS+LqlWkDItifWmcX9+jh2USAotWy
w7uf/d1JURwE1c03oryZiWJU0swzHp2zefAHkwhrLghQTaMHfUbSPT4RfrXaKTC1
9jxX0MlXP64M3XFQUymHLfdTjaMlwNhlHQT4XC/2JK8XaAveng7/ZI6klsuJ/Uwj
zamS98C6431US0YQ1U42GOfil1dXtTFbh52Z2/CAau573wbd/shfiUJLhb6rR0/k
S/bpx0SpN6oguqsa2/F8SNmu8bXAW+jWan5+bVKm/U/mQFCnZlJ1FyhT33bTsII1
Bvc/0xkpLE1qzDB9okOopinQy8+e4gWksVQlpjhpVj5v+bIahpbCirbrQsc8XfYL
i5WxZUKHzxOdL0PpRgAcgYgVKRnYbNncY9sSER/vmeaex/K5Esx5RX3u6JCtTOmG
yUZm2VWI/R+/PcgXQCzUgaG3dIvVNvyldtTEACWwrW6GwkeTWdrT/3xrVlAlH486
WyS1hSeR/n7qed2KI8PFykehfJLJ6y8ujommoSnLFsiC//LLRdpEMbvFJHgQXHAG
pHk+wTwCXSrAOBFsd/8jbCkIyoAg8/RoCEK5Lwg9rEtNQhT6zaC1meAVUHzt6QlB
wmcx7oz7MjTk3DpICqKKiL/CQB2OVM+a6PIVSgXL7U2t3VkDS6Te2i+ZXrsi1o2F
4HP257UJocBN11F5xlkYS9g1Rng4EXmxgU4sCQ+BbHQWz6vyEDv2xNfnT3QNPc8P
/SnWLSL47Hry7IG90avokc08jAQ09/jkauetYZwLve6r8wmmCCeGG8FdzXlo55R+
qCUjnY3+vbcwpdoc4AcdOttRO40Mx9yhrfDsmeCUm1uNNmfijJSzL43Almp7ktKR
yu19vElX5rL4PH6JHNZkzK6CCxFdQ2AQJJCNyFnvnVj75/xthmIyNToJOEzMLnSf
9XbJn02/laUPDj/5zqVkW6I4/DxF/B490351hkSXcYeu9pozF46fSSOBIYdtIDJK
zb3o/E44vPrExORjE9fdOwzsXbftP0Cgrwd/kXxRwQ1YEUH+HxIkDz7sbMWNJXMV
UeRY7dgPRqPDr10rZSXQKu8nUjFGyu+Xe9zYm9yWq2+yZSs2QAdcTJX5k6dFEvtm
lLC6ZMQqvXKBEsoWP692jVz0o5b6w13KTn8w+JAZE6bdsje+7nJLABYXI/UPQ44e
Y3R4Vq4PDJAyAPlw6Tl1460k9SInd5rnVJ1V8poYSpd6RAJTfEHAss7pTgB/Vzd7
i4TfO+IfbPqAaEOTOYHJ5lSARwEarw0EGWl5wHTJblC4s8AmevCN03ooO2jIbx90
k/7frcRdp5s26I4PEtiWx/khJrfPYJopABRGh15fWJfyZaqcpoYueAkmlEmLKqs5
ToYo9iHOp08HgmxPYdaJyACIkJuJLZDCLdYIsuhXzxzt1LTWiThyI9VCoHNz05tm
SyL4mcTgMKnC8Is4TDYiZcF7xlVUo78ecjcA4s2UQe1as4r8+Hi4S2W8KkYvLKJl
z3aKdSqEcU8IiZ69NSaun1j91/jzQ4kz3IUUhkawXPaS5FsPsHIlp/iG9BF1McY3
kvFdIwm43rYhdaRg3ctk4yFv46jr93uLMpcFLj64Y8Kj4GPkPfFxquMakDPXXT2P
cnLXdzmlxzffOVHdwiVm1+nGYMICeNOTgHCIIMl8bIF7cDR0soCCb6dT9Z5Jk9Wl
ouWoLR0hl10/AmQZcs3BJmqivNHEqjPYTv6paH+7jqnBIf7Wo9S3YVnMkW0N51Bz
cY88Cip/tpzVsdwPA9tiBoAydwzm1tlV5igb7b1D9Xeoduj+DHAsdvB3aUGAUSfj
S2t3fWceR8mIAFGx6/qaEKnOrFWra7wXEiZYj5561GpYxkg3uEGdCO+jGez79+PG
bfAHhMRfHW7E8wpJzR21q4MXz+qZBl9oAnCY1VvOjIF92qy2od5pbVOyFzNerpcF
vlmBdQyIGTZ6qTIihNhK8BaqDTzFx5VsulOfHiQsf5+V8DQufXbQygQSovUywJbF
DmlwgN0NyLaahuWThQw4KXqerffl0JXFHahEtz4SF7nvUgXjzjV/LPjqLyO61SG2
6n/A32Z7BnelGkZbLuP7ftoj6iYuLAKXH85/JcuJwoo6bDAJgrK5Q1u6WVx9Grwo
TlXxYc4sNi0NPnJINybyzue++E6LMo5vQt3nJ4KllS4fz5bgC/dtEPXBX2vSC+B7
yVAdjZ+p3hTW+ZKkC28c+fWbh5AKAFNZ7r9ZXbqtIA+xIyxE4n2IzUlxnyqICDEe
lPizqm8h1y4SFbuQNdDN9Vr2FIlzZiChwEphajqA3r5hksR+3YUhBN+/GHQ1xWl2
p5ZKG56Qsv1uTABOHNjRjnpHnXx5L1wjKAlWGNidBxDPeMVfMwDlXsF649VpUZsb
7W3dn6kjnHrO4T9zqwOy1hvty+qdhLjw4/jbjMnyUad8Mb9yMJzH96EgXIrVQMcR
0AgrKm/zjZ97+C9h7egBpfFhGqj/9a78X21QRpP6qlecqvqyOXTrbWVRTOoGoHBT
jWSlhvhbuVb6tmuCmctkF4A0enn4Wv0+qzC7aVgGY4C/rl2mSTzMEf5n5zDe/RHd
e5A30Jd25t+roV6cU5yk2yZ3JcCQ+Jetx1ca96gu5J1axxNSnqP0bRs2AEcdg5OS
Pv3TVLB7dq4UP53Y2q+aOmgB36ImpIl3q4htcW0tCn3HHeKz0uyfkLPuj94VSrSo
j+ASlhg/TUbidc/QDO+UH7/eR8stHuybD2ZKRYiIXWsnRNsdOF5P79Kw1ODv5a11
bCp/KjgRGNfbh3VjeQ2U7Av491LxfhLDSRPZNFsQQ+KRj/0TODxkzJ9SiwxNwlUo
VYuARqZJaQn7a5+C2/QPPrGrOy2L2EIewFidoUVkBIL64a3pPD0K3BdTkG4K6sn9
P5hqOkx9/zRyGTtCXmFzdR0ULr9IVagZU15C6v9wCZlgFxCIqMjdLrMuCA+VR06A
3tdI0iit9dybRkJYwrZL+QFt7mSYqwNnorLdAwLYIzymdABx6QrcimP0R/bNFzBL
k8WOjgRZHO0YJGOY9pen57jVM3s6FO1eFI5UYj+6BZqRNw14wzFZO7KrEQRxGlUp
pUNCQtV6QinHzhrsneLnOxxHSYvo5AIV6dVBktLHisxvzxeRVm7cUw3M2Fk4jCeU
eydkC+z2YkvqmgOIunSro2V9qi7UtIjoYGi3+vk2aTvzMECt5Rh3YFP0+INPifnM
PZI05EIN3AVoZ31yowogx3qpvIgtl60c8JZ/xdoJS2Jnzd5LtNcorcmDtKLpIqCf
1qeQykyFNyVuQ7YQD7AgEOKkj9ljDAm1BN1x+BSDJZ9YibnxGutrtaBTcalP+nj2
osJHDhLd6NWMWzP0BY7w8j+xbt0p1F1mUx2R5PVgaDJYBmm1c+WABCBk/lt5HIVm
z+JO/XZ7A6YvlidlkTF+8uXDMclZI4lrj2kchrezFh4/hIVJv8UHOd+dTDi2I++i
btCG5T1vw0/PrVQ/41S9r+zboRKOQTwTleH5SyVUMBevbw/oyc/JwSyPUa//YapZ
ZCVXMzR6B+AMid4jcz3MReSafPsq98Lbbsr2uvKjTiKElrrmPcVF8RiveVKHoqEA
aymJ/Qs1IaZ6fUTJ7gEpHhr9OreQiEeeG2GFEhHKSDLOwcepr/QGRdkHbD+VH5dm
y3BrFHYHPpJG9485yE2p+c/iEeL2Eu0Kt5i6dsXcKIcx+R8fYDINiXuHwxZrJYpa
lVTCgB3juhhWzyqRWT2rc7N3Aty8M0PAqoeliZW+YZw0X35jeTXvf/Gbwlesvk9e
3zsoRfITbHFzH3/7zZMshmXwbTZUJcDs5kp5ZNtTWjsMlfbfU1iSaCOR83OBT3Xd
6/L3sGjN8Y/6ZsjWi7wbB4h6komj7Lw+SuskJ//KqiuUYat/H8r0LssHBJLDSd/f
Nx6wZp5uUjzbz4Laj2PMwFlua6dMnJP3NfpckZhgcqOL+EYNPs1pLaJ12lACiTev
17ebClobfVcZeMRsxtLuw10pagjdncy9X1rrB8N8pzzIz+v7rcrqcpNau+0uKZbQ
bvOKJ+CxWqbtvopeQreB0mi9Zql1bBi1LvVtTPmbLHBJh6Ind1m54hx8eu7gQlVS
VHegc5YqUG4+eY89+HWTLwxmati5YaVPEb5HRrluCaH4uoBeq4zPt3gMkxdrbEsQ
JrrJ2HLGTtEl6rrkUKI4FJ9PjxpxmjxnpgWQ20mXD6XOEIwTHImZAHqX2FE94t3z
80Na7YL45hhmOfTAP9NLfhfRKa6oBz8YKEUGNk1N9M0WImEE1VgurNCQD7ifgIG4
kexzMXZx3m1AKSL0/T1emew8T2bN2elJmcXE8YDR91tY//fW1Nyp9xpoT6huLJ9X
kmbV7c7Vwe7oBMKyiwYLoHE2vVDV06rGb0LHYgRWYmECBuQgzXPzd57EsPJr2XZO
0ncfZ6fI/nKgxsUKignATW1+LUhqx33Bj8jx3u6S+6AjqHM1bs3JsrhXCNL6db+5
HiQHQW/bqilxjKhyvHAifq3hJem2TXEwLIy7Zn1OsvG4xrveLwgDkpS6mU2OmFbS
SI8bO3kJR0RvAkQVe2D1UKWNA3SK6BYBGoeeh3k8BbCHKD3IVjzxvVgTqoL95O1L
dGyeWqGzNhs/lhHds5TczDwTZLafdkK5isH6wsVrhrpZHlGdTuDkzXAi6dU/QvPc
8+0hyINjPiS27sGlRy1VfFN/cqTTMrsX7jTSrpVlfEpLfYUnMQ1Lk1mM6z4T50bi
rIDksP5blAYo4Egoqt2dgs31L2LHDgX96XbXJfMddvszEDzLtxcC6HikXZVUE/R6
3hjlXYsSV4HbRkMaquf3yKD/dmokPUdZAxgvpXDxgYcGhmuiLiay0m1QlIkAGSKI
hZpYsOQsqCOyKa9ITArS3DWtEwf8krGjbmzDTnzbYbj/7BUhgn93wKtxb724rGFW
M6xlApR8U6x6cZMzqacuIt6vWz5jSDBgxCjX9AzezlY+pO2nboqFEsgKJMkfKXul
dXcEXzUXud2/crPEb/fcFCC5e3wk+bOgQXHiD1U1yPkY4/7ouV6CEdOt2rqhBZKS
Ssdz+dQ3BAeUiCfKpR/o66wStzFV52YVpkTI0tADFrV3/bULXSeLI1rvdvaLmQnR
zFEifqtHljW3UAmrh6M0//YQupK6zmAInv2gUF7tOSkV9ng36qgD8RMebfbLsFvj
Vt60aYxpj+BwHPFfo00P9ngrYuWSx+NDVT2WaYSRmSH+Fn8G947ene0siqlRxU5p
t/5geHR2KcFaUSHrUx+FQRA6lwtXuhv44MyIjVjsLDzb3ZGtFjr6vMu3jqXGz1e0
YDwVNhCFtROi10hFzBCro+4MjgAXw/aKyP9FVMTKdmsIdQgRMhS1NoHLnh4rwZ1+
YAsMN4/UwMeZZ9xP5X+dpIN8rdNYliKHLvvEs6iVGC5IqwD0/Q+bsppSKGEY46yB
buD+2u0tvNdT/f1nIZMEtXwz+b2IG5OkzcHmFz/OKbkGsSWGuXnBP2Lyd3VWK+Ei
sGWob9BVDkIA34MpXoocGBPzLrTI9lTB5uoTcT64/KymESsTgVYtJ5ctlJJhrKfo
o4BtyDavmawZ+FMqqiX1PXbDCt9kUyN3K2XQ656ijrx7xLb/wp7QJCw0xlstyH7w
C1ce082s1OCVzPT434R/esmvyg7xxV3WOUogf+2BowlPHriYKwM7hCph77lT+pQp
hyzEWWFYkPCnn+rJlj44+N+CVDuC6YtVh/V6hejQtYzL5UkdlZqf0CbYq7TAisfY
E94ADAMEtPtCx174yL5nxd5KPIRVdrrjZkEXn6dApuIwCSe1rQa79RRBK6/4C1Rk
gyQ8aaTUtG/Hxskc0Onb3NCYAzE19pQ6XJ9SEQBLOPgnFL+S0d/BeSCm+UXqPHxq
PmKH106KRP42J/ySI0yNh1s0H0iQ+ncrkyANd9egzhOv8pPVfboTv0qVODG/6Ot+
5I0h+lnkHNacIbeyJtTdRIqyte57EoVEcBp2Mx6CpwOrDjXJ/RQj++08a/2eWZsW
+29DE08EPoCu8gR9AAWOtRX91OiLqNPygo1wg2DIIU3rhRB2rcmxQN6KR0I8WGw2
aNzuUNaltSDBCrBZRYV6qKK0It7tQP4ihsiIymzaiBUrurw3MB3lHGeQ3hk+Aa4p
otb+f68fAzG+wYTO9PRvGOA7Uy38shp+kggXSNTTw3hb4fBjSjCBGx4FHRgc1JQX
3W96G7PBI+5UfxMJWLBPrboB/FKkZ1NXO229z4RvgOsKCJGDqVA1uRuU/j1mT9Fo
o4/l4qWOrcc8maoomUcSo3r2gi2llXcVrjuHpnhMVNw+s0K77sRlDXUlQYIhl/Ub
HMxPKEAOkUwrIWGlFDdVyxa9Ster1i7t19XA5KJO+VKMUQlKYvVNZTg/Enmf1GV3
XgK4Di/V4eRknpLwI0AjrY4gZFCsUaDlKotWSDFAuB9tQnP+3FAknwckgngrT2JZ
jZUrVz4Oii4jo684eaWF5j7CktSCwAEFfHZz09IUB5QNWUMgRPS0Z1mtVu7aPQzR
/1b+UX7gEVfcj5lv8//JdJrB7Ie9XWgVelEHuS5k7LMKCQVIzDfQLJmEns4y6Fkt
j+3zXrFgRNMOR33eQwAfjyd+bhuu+b/BF1JzNO+oTrG9yaoCArkzOFX+qZBcY6Fb
llBMCoZOETUf6b7ek5msngC8j+qaDmT1ukErkVCV0i+WjJXst7KxGZ9PZh0VHQOW
w3KiJnbEyBdq5shu43nVHXi7ykKGZBk2sk6212HpwceTVE4WRsaaSPdWuBFLzxn+
/sF5xCaDIgyLba9aX1z03M6D1G2Fgrs33dk5Yp/6ibR1VYcKfewr1BU7IIiXkuzV
FXbGwjGUEcJyMfB+N4q7Jyhx52JTjzR8RIt2Vdr/EpNcUbIaIr2rPK8E2YbpIlI5
EPK4HRJnRQmKZGhfad9Sc24l8s8bFTgfpzPqV4zfljkvim00JxfEcwsnmZVq6DNz
r15v+wGoLEUb9l3iUgqIHfJtwJJeTijwBeE/cnkoefrp9TuNGa1B8mODSA0AHN6v
Yr3Nfld7dHTLSOdgD87kaWX4J+Dplhis9b45qAUI5P4wogSHr++N70kWXEhULjjX
BWfX25jFDTeswGEZtqQfEYrZB5Jj4M7/5JGtXs2nocLC2onCRE9MKofbNqrqgYwQ
900QVF0ep5okO/qgf1AVsZbvMuYesGwSCYMIaigCiZCO5oVno77UmR7fwGwIsTep
ILyK0qEJ55ReXZVaxLiAw1Z6NrckvMBCSiQaN85AfcXrfGkZ/Y1oWpc3MfFD+SJm
NGZUvc1r/74S8O00al2cjHQB7SPAS7dvMcePuq9ofKh/d7FT0WlKgCrwNcbtG/2x
4JTg1xKHAv3at98TRwETkRXMc0gdVebx6X4+EmC4qzYnWWiB7A15fV8TSxTj89pp
IzM7bxXhn2SZV5jcWqLyPvQepMxflfbhctKOa+j5T7oYDlIxEPkZgqkumHq08Jh7
OYPBK7YsxrORP+dtmzweoirmfF0VsNNImt8kgA//Qu/+Fj8SzLsrRoRy4J5DSH5l
YpolQeJSvUsLNdVMVE8dHN3LY302cUPGAkhZMhS4xdjxS9Se2VJeEejHIlF4m0Vx
/psZFGKYemmcU5a+0Wsp4Auy8GvvDtTAaBV/aDQopEsehifoJ0vfgQrd4NxBkJpB
YEhgRtc2RBZs8AlyGOIws8FMW2WeTZiHcLGFn7TUBxXQ08BXANhmuHLjvvLH4dBp
sJ76pys1nlSy9lWw10p+VGPMEFfN/6r/ZcqnHSKANhg3alTnBL6XBrBhvgDa1SYY
Sv+HQLVWK5AV+ufmM6zq2X84jbk4TZSvadFeFCdgRW5uGTPj0AfWj0B1eTHW+lqM
bo71xQw2tR1Sbb4WHIT670SkCKyq+8Zr14NC5VHYsWvSX0atp++3AYHEwnGaRN5z
lJNO7Q8sGc0Su3GnGnmvGb0K0eF+7Kak6zt8tW3Bgc3PkVWiRW5HD2JICxydcy9C
h4N/pyE3FS0ijVzIOnWERLLj324yk5W/RlTQUzZyQ89pHR5tCB0nrfIO84gFOoFK
M+g9/nNUt2bQ4Ns+cg+GB949U334kmyYqC2+kyHhWvK7o0GcF+JuVJJZfkeRWysr
NbfNNrTNqGWwFtv+w2QT2DgH0YxXJzKfiV/LkD61T7gae4cu90tZUyPQxrQjFdYW
ApyBCyBJ/XDmmvyZNDbabWN1ormLpwVHaB99w85TNPifWHkfA8Q3u7p0n4TMzSlI
PmOSYNAo54mojHRgyfAAfWVRHoHqOCPcMB0Ni9QZHk8CbQoHfrBT/VlHTTnr43aK
VIYa2fzV5MQUC3Ldh5IkESszSn+yF7CCX+X2zradd2M1Nwi5JvoLxaLNaznE54lg
2vqH3zx31YfrLNfIV7BJNzplLzJ4FqRXvtkT+w8WavnBhRblqHNeG3RItVzkYC2q
ZpsISPFA87tVhXK54FIfGUB0WSnkaTYAcmoKbIjF14yL79MD1NSEpShF9a04A+b/
0giGHoAyFsQtl0HKsHD8jmxCVCkOGcikzSCu219x6Z7S9ODtKEgzU7WVTFt1/gtj
Rc7HL1ucrTRgO1LL41LKNtlEWfXufowL7Hn1v8BPUzTODn7k+rdf8YpSjDHPcVwJ
aKIJRU3tGmBbeXk/iATSZxEcFGi4FYuKccC+LvuhoXu3AHTjX22j4AIzDlg3hXNI
sFSU8pY1c9X2GD08jiI4ar2g8/4MJSFgofqW3b60LuB2PnDokWP4DzYflzZmZByu
VaF4GzBG+x1OsgKKULnsD5Cd5JiDzti8d5kxo43fMnX55NijoE1I+8aPagvCoyVw
xLn3hHWG36D/waOPS6zIcVdbRd4v0NXgT5Ik6xTG4D1Jgr2nXvkRUZDe1XPb13Cc
v5Mrli63tZLXy1kblCSDQCIy/aL8UADEXaJGsN1FpLeyLtTCRcgs3iaw2zEQEPpw
uALo76kZFtpfU8BrqRrmDOCDZlfNZk49pCjw72qCDP7eSNTdBEeyjheWB3VxUrr9
jdXmzv3w1tGorLCyKBT2SHEiDY0HlivO0qrBAH5PVF2zCyPn/nXCWkNSWVpOSDpo
ACoC4RTmr7R+mPDwMhdGh4beYaHzlEEvBgowDfaYtljOQxdIEWpU377x13dk93Vi
D0MMDgfLIHpYy4fEkbRIH3TbmGtmbEgyzsAuuVzZ4fygq5cEwcC7de+J2Ovh8onG
q7MzN9JkSHum7sigxNS/1F415a/fUScRR3HhtlA3AnzbnjEaCQ4bj+WyMgiKz1iy
BsqZ/eG4afLI4HO8JtyhDGCkRQU2Hao3U/nMY9sR+vbbWNbNrkbNc56ypnygoC/U
ohkijQVxNiqmJWLS9DTIsO4+VIGiFO/tGbYwfNmeYcTYO/dSMNaCR88VeNHnwzwr
GFyMZ01JCeEC9wRwu4jC6kBy0B1WKYE0RB+wWghX3nIXgYViXuvp44CmhrZFaDVB
O9CeGao4bneKIFG198FpF8atxVvMZqo/Nm8BNrUukkCGf4OWK/nnkKNqCz7fAAA2
61lbSr9I1cA2qRRBBJSvm6gKr9PQ5KLk+HeGHpbfLKZqbY78z8EG4n54/ps++HrZ
4dXAseJBPYtc8ta3r+8Pwtg9USlNrytKvNgTOo6TwzsxA6TAIQBEyZ1xK3OR4ydY
X/m2OIB29RcLNGsh4ZgIwAqT8A7tfzmVWD0ujReS4HUwlAo5KXfUyr3Ed7zFAoZx
6sS4u+M2TeT9RnVib09uYkYTflAZ3Y4kg6U7lfrBCbEPY+CE9glyaKgL63Nx8Rrz
yBC+EtB5iKAWiWBTF1D//wTJYOBaoe0/42cSXG3r1AMHdRw/NMlY0WLwtBd8sgGY
GA1r5zIdmxXMaY+eWhRLEkpAgEnzE/THatmMB2e75Li4Y+k0JDtyCO38mDjCb9AW
dxGwrT/sR7BBhbUmAOUUZCm+mF79lGbG5zLoLMTaocrGnVcc794g9b6qnZENXOFJ
gDo1gZGgBZRvjJka8AiR3qKpLHaDgL2xJyAw7ur3CG4=
`protect END_PROTECTED
