`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6JcD1w3mTtebA3Hx/pc2/eVayuAE3ndB4xbhOiAOoxXAQAVTMklHrLS9CZAYQ4PR
Flj5UHZL1bnbtxZapMLX54jdYCxKv0V0PWx7X7/bleZnhMUHO42byZk2SrGUHOiA
jWpcDkNsu5rgqVVL91mQ1iWlmQjYp5MZOnW1htZAXb9yuODp2kX48jlL/QYasl7R
mWgjUM/bgxqf0f7cfXJy49XgLo+I8u80HP7wxKqRuR7MWjZkZmEVcCajm/7eglSs
ZOefo0rXWt+lAvHTSChis2k9DvZcbQyAkAu/GFPC8lwepJySYcBYJ/ONOi9N1bTL
2mjq7PUkTCRQpHpZ/0CwtA==
`protect END_PROTECTED
