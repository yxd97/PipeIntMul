`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WoZHJZKmrWiHY6eTDjODOnPccys7HVBpG5ZdufZv3w1nnZRGgB6RolFsMEJq/Re+
3bDAVy7Qm63vc5Q/5JidWKTU0jrro7i9CGevCj+k+diYmCRDQ+D48bhRndDIeFh/
OXhNPz54/zJmDaVFm2ASD+mUa90LU8qrn88s22d56AQ1UVnLb16f30JonQoSBm/w
/ZRev9d16DOi1LlFkD1Y4BvAESgpXOMIOBIIJx9dLl5LVy6umiVgBYpCD2chj8L5
lUpkfMxOvjMsO9JzZadxluYglc8/O18rYs0fg02abqkZtpntOB4Bjjw+eCJloqQm
ulg1AEA+UF0ZUNJTjETeRKXMYNAs3NsWzY0hBV+FAhiAaIedPQGMnDB/mfb9yn5a
AWSGBWVSHF97WWmKgeHyeiNz4umGXtHD4GJZ+iYcXkdh8Mz6wjnbU4hCMa47GCYr
ORliM9dwsxoP/V6H3g0l6Mhq29fI/2d3TeRXQEy3jU9BpBtlfTEXzcPpUp4pHbs4
`protect END_PROTECTED
