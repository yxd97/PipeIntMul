`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xNxpzMFqDYgTATccnwRWI/WJmyG7NxJe67T3tEl880+t1XTo5u03jKX54mnvHvv
w1/WyOHpXgeipV3KkCEsqs9CeYRe4yqXpSKWr1nTWJpE3MgANcZwW4NN7wBd/Cpx
dd6X7FvKvfkYEukaHSlkq6JRWm1qiPDpqt9lA/CzQu3t205iJkLNT5/XUmFb8qCx
uCqa2lPIVlVfP5JYtuHlwAxFLhGSA4gNqaEMpYAWDNARTD2TCovW+zIcYsk4dQN1
SdFIkG3oyx6dGbjnsfOUP/Sc9vEMACpcdGBrhBqenNZwfMoFdRkGsoz+SGzI432m
N49s7/kcb/G3NojRHk4pMbMXlinyfWs0OydEftPHn0+9D3fRAWOeTbIO4qBD5iT/
IgPEwi0LeiZ4w8i8XrUYwwCQ3bzq0Z28U0f+5BP6K60=
`protect END_PROTECTED
