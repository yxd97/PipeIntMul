`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97wR5Y2/gvsGoHn1VAlcNVifn+BQU5EVh4B6R1AQVTgxJgj+FVLAccagJab2uuVR
xYuiisdc/INa8fk2sk4/8BO/XtWMIWZzuNY0OZefJmM0gIGjsTM/1wBplJi0tIlV
wqtlEgdn7BQnaMl8/5S608apgJ5d/9LxjNSirEBKvHQwvdSIPSKt5VzSpufkLits
gYckmrYych61yUMjwswKmT94H3FXKxi0Ee+Eb3ithJBW+kpXsOeU8FigOz+yWqm7
z/T55tAEmJ6UR3yq2A5nSiMdfte2xPLDF3xldSH/OGlmaXa8vSQ5mbZaapqk1Xh6
`protect END_PROTECTED
