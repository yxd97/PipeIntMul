`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1mIJGnNg2X5eLjmMOJH0h5RIGFvAx2XHKckV729tAmDtDbwlSQD6bUJpanbwX2a
KglOD4KZf0o78nGeW0bGjvXCxn/aew9R+85c09A7bFyjeNO9KxW2SUaCY8UrLptI
nzbVrPLsdYkJ0Su64m+nxwdFnpr9oHGcvYBYEk551slEwWaOkdLop7hEUVwSnZfY
jberFZGogPhzG7UHjWgu0hlyxOojfDG8Zggx4jB3T2ZCaOaZOfquEGXkKbr6ZDe3
Xkdsb/UOjcUG/gZCOsDYW+n+zR199dpbNKSisfVQa5+dIrmXcreEvSSM+G2SXvtY
Hjuy/hvPr9OQkF2Z2aFsrQSzbSL8Kf1HmT/eqjC4MuEY0QDPVPV/vl9afYM4lxll
FwRTSK2ndIYX4G94lNGqu/Y4/rmUcU+4Wtq2f8ldpdH4nIHfmxUvPltuyRTNLQOZ
UdiPjhVXoukStmuEokDVTKq7jPrOvODDH3RPPJyE2acF4o0PQAV4RV1mXmwqhKP5
NuMe087A43HfJ6BYM0Gst49PKcx5xjylaqM06quAVVzGCxZ312ja9M3nWnAvkQHe
pdq702VkMh93jOEuzWKCLRjO7nNp5M5aWurMz9NIt7NLca5UAsyWBfGgo8ZtJ96O
kMULBRaD3NWhVFYoLQy3zYbKlor/R5joCatxD6FAliHHtyVHADfy8tgsa36IQjdE
0St0v4/gXHAhCzZgVEVKgCC5E7Itn21yCQhD3HzPSILkr2DXefHaGghmToS7yX0p
h50u8bxm7JXbxmg12l+TK0/9ELkAsYKW6uP8s3V43Q5Zb9yilrFBYTMnyRCjj5Ef
ewnG+x0FKqqSUaDx9XsX7XyFGybiT8IEyptMeBTpxuTQuEwy9KLyHAANfId10qG3
RaLnkDN4O3W71WXt7uRfNRzMRRxOUhDnvVviAJ9FO4SKVnNp9cyb/SsMFnSQUOfv
TzhNej62rNAD1LoNV6rDym+mWDAtUJhZcnBoy/UfQV213ziW7sVNzpm50viFsN9A
aDqioWZudBl2WlYJHEkOzYCcnbv0OwJTz61habNs9lDVcjDXYLl+AEiYupBk6bHG
1YeWl6Yb3swtKhUaf4yUhjEvQDKuA1TIA+4Ymb3qUN000rt9CEpIq8VG4UD/lAPJ
UlEfJPyUi25/jLgzWUZYhWtTxazR0sBYB4iWaZv1oqg4U8eSion9fejwp4HSzq6w
ytR8ZojjvOna3XBgzxgALDIPYubsdKhxblrT/6DGpLHmAie1gEqn8GtiFk6qLWOO
efwmL6D7eSYibC6QWwtQP7Jb4WgHJsEe7HccPGQN3dp9sMFZXaorF76C0QM1mvGH
t7yHuWUhvCrkayO0EqI6cjFVhp+4E9DE0gFCQbJfcFG+vs1ClNzrKrDaEINCOosi
HfCxF3nkOkBRuJvqh7fupkIT4s5siaAx2G3KkNNfZb+cUh+Jcj2mqmxgTN+ruF+4
7fFqWemJxsFkt2iIRtWeTgB0ceZrayCZsk6Rj+ykzex6wCvRa6ljJx5nsGgr9bFO
bGKufT1JmyoHu8PDdJIE4Urdw9+v7TCvipsi1c1lVGoTLlwRLFBwp4wJuuhoWybp
6AdR/Dty3fc1ZEch4CMXgzgCzV7Wc/sy2QD6LHkn8Hl069bVHTG+OOoNsZWe4Dpe
sQkYSyLQW5/eslRyEvsvHySb3Rp2/osGrIhMEZk/9X7eZefKGXusea7C+ass4gjD
22TM77eIgUgdmjY9uonNLw==
`protect END_PROTECTED
