`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jxdl1uutbv2rnpXuCG4yvjEPsGEL/+1Vz6IbUSf//Ojd+QmW7iEQytMa1XQSyDxS
qB97NeexcqUnPpvccQllw7Begym41E+a2Hk0xJYxezHhC8VGogNGJ31bRY/LcMH0
Spr5OzjFiA6oBUZ1e1FofKkXlvFP8MNKPE4i+G/yqIsiq4RNUwxkk+UPzKV7efoU
Jlb6TkzhM4GE/PYCqBZ0JyF4LGqzZDb7GiIPFvZQuM/Ym/V1hDoo2GZFvKtrjLRE
enpZwI/TL04KOUcrNyf48wtKnjteMI/uD1W+CJVZDa5SpkSokA+zt6UeaspOYUzK
Pm3S/hN3tyS+81HrBPoY2C2Z5QtiIlekMOwPjfXmg0FkOpH2WUw59LMyHLvdobfp
tUJzAgTBrqvR0SlvT3K7T9/8BzedpwwW2Bhz1VW8lEbOwqPTreNWZaOgePVo7gkO
`protect END_PROTECTED
