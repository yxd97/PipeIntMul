`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I+WftnTJ75qDdmQOq5MZlDXYWsPLRbhb+S/kJ7c2M5J7SJl6FoLFOlCFcpiblzFL
HjIIT900N2YHKa2O9Bn8Vl0bfFAPpvhKaS6hgzFngnDOhFXkzdUiIVWbCczbmlHL
FuQEwbFk/B4lAB3xD4gfpRxURhuD09ShWIwOc09z/DSfd/kZBXguh2s+Cj1G5ioQ
sqGuVDOXtAF/d6ww6LmK3PdsckctIs3YHBJ9EW/w089a8ZHoVGcHNMVMTHqRlR28
m2c4sLIM94SJSB9oAWV4EkXrUD2zxr4aJjI8ZXDpUy+Ih0MAVt2cPJ02CXkBe7Mm
fkzLRPdOZYGfQH0niKCKJmxCcV2gobbT7TWfB0i3fml+qwvW4luH3CbUBu2S/TF5
nEBVcke3RnDL7FRxqdWp7e1dGCEZpGNy9cqL+y7XbGi7LrekYLkazYgWCVbCj7GA
8Pcnn0XDHKCIwVf32cSGaufULqyXHfjs5qfDVeuXGP6Cf7L3SLCB3w8b39zrItgA
tK2sQwSqcEwmeLUcDGCrI0VUToQJ8k0dFbqNJV2cwrLRMkNiB5OtJr4dr9ewNUY5
7/y2VromFg300JmVUboEY0TjxEovebL6PxSXq5O4o7qEuoYUH9qPhlzKRZQUn14f
cIbVqK2ug0QDWlurPeurEAevLBrJ7ZSrkInm1OMMyLzyPAxCNlg0BI1V3SuwEilk
dGwMr1VuCjlZAjJtnw/pwCLha7fz99VkSFYdvX6DyaiIJpfVJ9hRAMlyp3eIGzCJ
s+LAXlnEREmCNkHUxraPzOAylqhfJmS37V+j+tot9QG1lGGRCl7D8gon7sXjWDFM
SQIpjKhrTRiiCF1ML8SDdYufO9O8QhKDJdAhztgYvRQxRBatk0pazu5mY68VNgyH
pwV2A/Wj4tR1f94VJeKOk7wYf/Fk4YjEEfO5l+wYzpagTa6sVhyenUOgenjs/7iB
cSQkgfUk6/2Mw1q2IpB714yVpVNK6oPeKnxkYutFFFmeHXWBCTJAfEFtjV4Cnd33
Qr+5htX4hWHXlshy8rCMdwLtvWrsWhGkC/tgSbOuokQ=
`protect END_PROTECTED
