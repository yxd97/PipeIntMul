`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dBQhU1LFtZE2Nn9KUkUfFuph+VmuA3RCwmwHJVPZ/W/ThuNLRuh7Iw4rl4Rfz7BD
0+LZZmW93+2XeQXxoF3ehjrjKl5mtnOKssjcijGLfdAgl7r7AmQN5f2L6LC+sM9A
bOeKYKiYRcJA4NbKBKEk0PTOwtNBWyBnBXgq3qE9ZFCTqn5dEJyZMKdAirnDZHSp
z5BQGBl1Rlw0qDt+BrYd3YXqkr0CHP6v4ZataEXH2hVwdL6gbKOG7/C9+b+p2Pnj
DzZMPf9gSxro+ROU+QpN5D//g+nEmevBpl+2kVRMF2Fy/ykH9IV1QvfBNkb/q7vJ
u0AcMtm9hNcfUqyIjsR1zTc1lmYtTCaFf4QSxkQFrKIiym8j82HGUETSTlc5LjsH
PD4YWTLue/02NVCKHdA+TfFAYI5fZ9LNJgjnz4BVxcIP1viLQNR42J1udxajv64X
wBF0DzrW0T2gkEiR4vVb6kz0a8XyYtUi0YRm0SP445VCKf8GNkRkFaKv00XFwohU
vBWVfWsrGf9qOW0KzpXdkXhIxNdFKiXUswVjLQ2Rt72tLqqj/QcYXucbzDWhoolb
v6Od9pEMBkvMDz6T2lRqO2g40sxOihl8gaZu5ilOaO2VxIpAw877NmSUI3Y2VjQH
HpF9RN6f+P7YZs6mdrnB9Sda+wF0ePRH/3/ozXoVLXrAMZmC4Daa/h/qvuOTt+lQ
wQYeBFPaGl7rIWknhM3TpOkfZqwz7koKUNo7ZZNDg0aremI0SG1dmsH4OiYLhHp+
2ckHgM9epaDMIZzBzYifefQ9eTqw9JWQPU/DnBqYIU9rPqltZdVCZqZfbOrkPz1H
Tv3XyiNJJtCDVBZohGYZJ2Tmv3iAE9vXPHBRr1xrW1ub9PD+ZDMNAHtFmBIeoRXQ
OHfoAa/Xg0XBEX691a1Nay45hQPzRFrLF1dgcE5e7rsa6kxyQ6d+JpmTBiuXm0e9
uk3Kx2UAYQA7GPdliPRPSpf/IVVWbT+DlDyKImvrCxuMBchDWLzytrkvzIgeiQI8
`protect END_PROTECTED
