`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sJ1nCPGQRmkErWspZTDlHW3SL1O5PGpCBmYggRDAnsDOQNqsva+pX9S5mKihVLCT
MfnfhUUZ7EXlG4N/YfCxIWvf6dou82mgLdObOsic39KONqLcXtgBTiQjE6HkYPBN
r6oYlQUgqzrD8dgCxwGiZlw+XFC9Z4PUJvscUD4hRIbNhOleF03RtjTt+12UJkXX
5im76jioddaxiVWNbLp+LlfbfZticiK2UWTsSDMyZu2ABFfYasQaTtveF/qyK1KU
emuPwHrVtY9smWS+FCXgGKDRwg4rZ9XSMchiPzu74i31B0M3N025IEmkiHoGZVUl
zr1Mq4LkBjz0/BiB5tpFGRQsDBq92IyZNQCYZ1UFck7Ae62CEh1llvNzEWy3Lo5B
8lMIMSrcOBwjvUGNXYEo0D37KxPXA6OoLGcNe4x+eFmp7dckxYmrL54GdURv1I4v
qvgk3gmyvEYWrG/jBvmubfGWYNujEW6ZY0mp0RuxCls1C8Y/L8FfYvE3Yxv7/68B
2jxmE69tlKszk7IAqaqrBKuNK6pvXN+QVmHPOcGcbgqLc64nTG4ut/RD0XwT4l8i
McdupSyp2VGWltN2E2LmNuDgmFV6Iot/dAG2XNVsHJTSinUATeXG9sDpewudVh41
vkqD4OR797vYgCmm4VxTGiFyZgjzMO++efSGpD6CBNXQ5JII2M1MTxMweyizsQqa
WyUyKMA+rPunVlC3i/bfLT6QNnMJWiQlFR3vzlVS8NTpFDlYZrFOwR+nqHdOIp/R
OPsYuaSYTHDI9IzTjwN1lPxKkSyCfVFbd2RHouLYn5IIlsoEr28WZ1WHWnvrANtZ
ZxaHvOA+CYuaKQM2u+csnxhnrO+pGkSNgO5YIZnSUnZKJSlqCekMOwfzv/BmXZZu
7YxNt8Q5jtXJBlYL4bdNCDyRRluNRgA1wZi0SSm0OAyTPIDCaUk7ebJG+ZE83/Wg
jcIwRIjdZqzKYMzVljq5jsdzjUFJYyZln5qPC4KbMBAJxxGsezsaSZWDt59xJiwv
rGqV6rnfiolaBz9TWzKx73tgi0hiMxG1tJpQ5SYyOyMgUMAWzDDHvjEjGmW3FmzC
FVIPDt52dTEiq/BYf1k5p96bL1onCUYcp3NVzk+thwLloL6+R4V5SSFA+8U+iLtU
v7NEtrED5G/kNljsF3cxDmH6UrpyF/JwjQIyeH2WzvtKRSy3zPTy9wZ6uYj88Fmu
8djKz9xsOupLx7ukLF+RJWd6h3XYgzUssmYNEoTNCQp73iL7dXrhfbOYfh3NwFj+
3KY8w0MRfmhCYdaagM687QiiLRNlbJQgI5HTTogwCaEoQY4bPxf/FZiJ4xza/sT0
hm6qFrmj1OV3nOIGvygzA6jDuqMDMik0k1QClUU1DD3MEdvIAfIyr0pXv9VH+TtO
bwaTV0nNSowSsU4ZD/hX9kOFwIY2hxB2n/B6aIvvNY5XxDjucsRrtw5Rg93LXSXF
fe01meOwWcE5bnfpX2i8WZPc03PqvEtKAEaStWRvYUaXvW53T9si8N8j/bYmllvi
KWZThq8j2yux67X2uqYYD/cjERdQPAbGB/gOZxQGA7wmomyx8BdzmwiVdHvTH+LZ
gYs95CMUTjogFgFYZaK7eTdgLG0iuLkJIhWl+T49PIOQPInG6wbafEZEfbomT5e+
TANVDh1FlQj6ZrXQQUmU7GY/1EbVrITUZZUH8fxwhEmd63wvCQBm41oE4r6jtuWV
8gb1GCBZsKVeTSO6xGeiyVNhG/mG/0GKZFLQM4q5YaPUWYHBgkqicQ4jCIPOB6bg
zr51hr4EwfFXpgYPD818LNYcXxBOSfCm9q2xd9eNL6oF2e1lHBav0vfVHQNi0lgG
N9FIg32MtdFRd2DsmhixCvwki+uEg7F89zpITq7kjh6oVzTL/IhK1F+jPSPEvpzQ
JMKJAXml/UiqwgWvmJg2i1D6Lo5nK3gAgLMCVHm2x1B0Ds7v6sXhonnXbUMM39Yb
sR20G7WqFYL4OaBeOjNgR8mxEoHhXy3VBGSDBBmXPyQhuO9TGZc9j1I9tJrSmlyQ
/s2jpda5fOnBsCmPVgbZc7UMW7B1bGSw99+AmVQYUZIPpVDtsWJvhvUMVgP3qC1g
Xib1STzuAg+dIUw4bGdLPM9xHliaPcJuGhNhZw609A4x36JcTrFkPJGPQ/K4Z01U
doLyk19sVV3SL1+lWzQjofU8P81h55BrcaSnrc8z6TlgbtxwJHYMNgn8ol8G2t8i
yNcsauEK/0w8ClTu6tYgMpxiMBviWivQp24AH7wox2Z50FYrZY1ea13u7jTFgkDT
M5xSznfy7J/y8EmJ20NxSo/vQ23VXOE08JmnexSnaPs1Ho2K/GxsS7m6Nyzt3r+f
3UZt/ygrZaoMBslIEBJRnfKolWrdIs2cgxnUJoQ4RWHQpvTN0RROMA4UR0jjKJB3
KZFj0GAO8sKq3Nd6lLiHj8XOruAunvruPbEdUgoD3d0cLMuAHJUkudK1xqWPf8oQ
cpOPIq4kLdY7I10liyV1GaqYsqlPXspICObrln8fznX4skegziJbSKa4Bq5RTYsm
rOVFRe0md3Lj+qoptC07y7B5ocL/jGmv4onSWHK7tDnYOdH0NGOyh/+naYRRRrAg
G9tFxYN52Hw0ZJmT9ffnXGFHrUkfUuSMu8hE6rgph5lrxGS8oARdjb32oQnGm1t9
1caUcndQvlpH8iMIqhfJ8E4Fh29USlXVBhKgwlie7X0ZQonGnQsYctvPFuOwCVP/
i6S6igCIgA6u7I6D6ntQNyM/SLs4uxVUTVlsHKl3LI95zMnOvSJ/OXZh4laddjS2
OZeFBSNbLUPyVkamvFT1dDByXKkEeE9TT/fFPeF+mBWbgPpRZmG7SyKSFUNkPrkb
09Q7jadDdfHuPXY4ChJvhwVOcMSj55Wa9RvM7M30LMzYNchqeqEO8vaamMXhL7s5
bfw0e6YftCfBft2sm4tc8UAHVePvltkW4gZHrq23nbdweGsq3wF+oZDXoF1cmyY5
i4ZrV62S1lfBLvxVSvaT40gCFHZdMyXrKubAQOjfAJkoMwaM3cfwW9+xkGEOE6bS
GzTeCk6fkOIO334vySG1SRnqQBk4ouyWdi2LuSYrIcbFR8rwKFKceNcUryGAH1RS
xK9rGjdDP9rXwxahRqCUFxFKJq9bIVufWIVUrRtUizopF3HWfCU8+ksoh+fJz5Ru
XuuPangvp/tewOjdZ1wbdHli56APqwpBx6wT2m9jlqLQJMahJK5h/SIPJgJ6KP/v
w+0MDtjCwEwnTfxRaVgoi7e/oXHSCg931wc90WOQFW0l/EcWz6sadrHUUXAlHxf0
0bDTb7O3/zTuAigG7z3wEt2bDo/f7yI7GnTkdCLMj2TkQP/E6e6CH3y3MtXYd3W3
oToLHHsIOsnt2inVPsHIr0i+TYYhITxr3r5Q0rynUtYf2IeZqoVZAh9ut1nT2KyN
/3kGN0i2CvAxmWHOcUOtqpbSQczo3hAnRH2ImEr0CCXWTvx7ae7Tc5O39HPZFK2C
3G9Q1YD/VncfpVv7gnEjxJQJaSkAIK38/VtyRrBhA5GZ78rjkJUYBppe2fBmz3lq
8/KSy0ZLRUTLleUTQtDvnsbJWUBfiLAgFjL5mCBXKgpYxEgW5NubQ4U+Oi96EtNE
pteuV09DAfsNAcr301ZaIniHIxQ2fNapCgtBab1MtHQrh8t048i0CK40RkjzvlLO
fn9a0pYguU83+pi2jEHuMaBwdM0GzaSnBSe3e2kK+YBKhf11dQNba9T4pl3aUSmd
Nm2wu9E3YUYkuPnUx/JBHTrryCGM3T2bH/fke2MaZ1NGKB/1PE3ji/dNX+qC2qdn
thmj8pMaFXeIRO5e8A4lqF6WRBJBnbWzsIoakydYe0ZWnIlP8p8ygsk6RkWvrl9E
JE0XCxskjTsFaCiT43yYldJJcFVYT3r9RPBTqJ/J3MmR/WjvlAg8tJzl60hW95Vw
axNfOY8SJrpU9c58kFxg251zS7YiS5lVYggL7ryHfJS6jceEyax7CetR29G/knWX
hAH98YtjosrYolSdSrgendoqqiS/ys6U5L8ITPRDnIlm8sWHKhhm82Hn7h0DCe0v
YwOlaEvSCG28ZQmz2N4LgrpywwtQHyDIfURpbPJuFU4S6vnu54dfnOdICXIrsMFv
vZxFlpFlY5jiVyfzfKO37oTFx4byuWs6cSXAH6zqXNyDPNAYh9BGKVyyuLfK6r6U
VVu8z4Iwelmv4AwkMx9KzUntbR2ZCq7mR/gz/iGF25R3b4mQrs3Ohutts8IMB8pG
MfMowmLNcijLBME2z2VN5FDOP5qkRNmt9t8T1Lo+5lc+lMH1thJbYDamFwpt1c1e
P+ESNN7f9BcuQHdYGfnCVzcZjHKCC9bwkD7aQWMgVLMpYGU0VzFZi2zK39UnJhFC
dNY7A7pirIjVT72XqXdp5+R34zrNhsZlqhj+EcTrEFrpdq0zSLjwAPEyPZUOrlx9
yfHPq8jUWxmS2WiuEYueZRCo1qIqY5IxTjNONMGZzDTN/poHyTUnx4YzOqaSOFTf
mi1bUNFVXDRXA4Cnv0GcjIvfL02rz9r4BF8ctm+YqeYRp1wqMdzfA19qwwpunhIt
fzT6i+5H3XTWXn/ZB/7RyUsQ0HQiDCyBSnZtZJFlzwrHwRuC7j3ngBYnHsQZVJu+
zYn/okOto86iUKon+fDIIVhxH4gmrUo3bG0E42p3T0bUJNqyvVCCf9+DLtztjdxY
AmQx167ZyHb/HSTR8E3MyInwxL3V+s7ZLYnTEhbdDeu22OwY8VW+/LsF3OpCirwr
+mWVWWK1WIk8uqzEG3Rhu74NVaAoKi2yOupdgTnDqz99UHf62WYtIrG7x8FXz/AU
XFE04pJAPAp1L/Q7uZdXw+0GWrfqrUKZQot55NV/GlagszcfFjKjaTGnhgoiyefc
mfm0oWnG7LJcRJ2BGflnfTclXzouLMZo4BqEvTmtz81l75FntTLFzMSTqeKPLux7
Ksvl2/SFDWbInmkhcTbumxf45qJnUQOdeR5K7Fk+ICKZW6F32A710H386m0p3tz1
VXGVtKV+ld4CFDfP+FGBes1EOHxAcpNkgLWvbBCH4vYw/94M7PUYMe8wy7XWLxfu
VZdR1IcM+MHkIZ7iLHQ5kLuYNWhbJQu55zhUYmhg5skHjHUpbXhpvJHr7gC1vi9v
nC5lOsYxQdkOAMfXwVESr4UuAg0O+1zwjnIXDHG3YuE5uoUWkDh3aknN76ikUIsE
7GTPDKD2+lVNqmrL7IVXUIeU5VABS4QntmgBsZxRSdHy6dRlvYVzwzFmDlI/PKEk
1JN3I4WQAcVN8zxiBRiSTyEAv3iKm4M77x41hCmN+5CE7ZmME24L+Ifrt0xpYwug
0PI361wrSfBQxxf5oEjVcUKNtZkJ2bTEQTXgOjw6YgqJ+tObv/GPQI9gKVEF76+V
lRFHa/2CzN8eNUb9nPBgqzD+fcRHvymZ1FQnQ1+7gkpj9fVaKuWDLMdftPZQUOzN
3zDlWWJxjdKfUVzIYmSCtV9V6fy5ZHMUTCimda8RQMwaPeGyVsMoDKliF9wznDeL
KBPCaAWCjv943MwZUCJ9vK6e3nE/nHukmbJ1e1/KHXjxYHlfOxO0BNffjxQIRJNG
F+iz/xrPdAUdXa7o9hRtz84YU/CBYZnOpKCrvC7lovp3NyYJfF9CjORSaSBG1Y28
OnJ6ShkzinYalG4//HEX59oU/YWp27pIoUJjT3QvsoT0LKJJhBVqzPb+w4kquiAe
p6GWRhZqRkE9VCfZrcRv5EZYpU1h7iphFZfLzRQvNtOBQO8jVlLx8QWGiZcNJAXJ
kzxrsoCTRAT1U2tu2alrmhJ/9ZRW0Vl3EPhzOe8B6w0WTw+AZ9MK0Gky7P4OCwGq
6Ok6meVM9X0WZL0trp57632MNPr/0HMTPy5b21XpLq2MCwT+rDK0yQq8yv/hBOQK
FTmc34a2ZY0GMKFeH6lHTJMNI2IhJ9L1xtVSMiQeqbWcfgcJMU+k9kIwsnM1g34w
8Xdx7kg0CeAneH1/srz9yrQWJsHLpoL5pMHLxH6gTNXsWlXQzNAv6kOEbFpzdVA0
nYg/XwuUCIhmzejr1d/TtVpOt7uPZy6a+P6gcOLnjHP6ZWE1c/TVDUkWMdjwXEkV
Fm8udkp1M16Zc9RMdqu8QA+HwcQ94RRONGVj6fhZmvWb8x2Q1obMSf0jVmj8RTT7
RR1pFgbfTONeCkIxrYUiGJiBksSyMStxfxopKQ9bqdYWLPHiXgR3ex5gwiy1fpsa
35L7PWqPSQG2c2Db5ddFsFvhm+R3ngC+xGe/Uiue7o+39DbkwYpqR56KiUvLBpIO
mpSZFdkfHUaWSlkMgZjKTXETjzuCGxGcRPxrQFKfjkxPfyhyE3G3SI8iybjjszir
m4M/cYKBZapqzYQe9VplctvnLo1dUJQwZvcmEQzKJHlBWNL9pHm8WcnAcKk5OVeR
AjfTuelXYnJC4KPfoQKCQZlBwzAGO19v1cMv4aggXCvVTGMQKW0mJRCW2Ss8NXsK
gqQSy+2Ci6HrpvN/xFwG9fbMh/GO40FB6W6JqMpkqBL/4OkVO7HEoqWgLBBJOznF
qlMirqZbCngLUyaYinTUO47S9HZn2eAqYtTvNR3laFtB90aem/15v/TCSvfdnbw9
cjvj9OISe0GF04AGVLrtkI7nr1v340X43UqYsSeQYWhZVkm5Xi0Mx01oqdnZEy1y
p8YsczCU8h+u1+gAEWWkYHQgAJZ/oCGePr9VjfVW04N0em40w1qniBHAwY40Qnpv
iypjKw/H/ZYQOgqfPLToiZlUDpebFW0AXSq5ohzNH/Q8h1Jvm9MDd6WrBmXS3dce
RuVEM+Vt+cvHT53TZJUqWbAUtfFTla7Bw42Cc/LUgdo9uYYCIAPv7MU4j9DinUty
tIBEcmk7CG2q3jQLgx9pf7ZL5Jr7YOeFyhDk/P+nLEJhhvSWwHHpP3vvItZY1idn
hSb1oc/9HnElQZdxtZitZqW3s5xKTjTLLz7UmPFMTFpHyySgdvj3fj9K6YCaZB8n
BBxnBFHkq39iTwq94Hy9iSheFyXshV9aWF2AmSJC2En+cJhrKdFFMar5GQC/MQ/H
Y0x4kExaXFKOnx6Y+2mEEPbpm3EbPNkT5C8tqvz3oSkSARHnCVF6sklJWtqRAX1f
+9W8PoFjJU9JsO4UAXFdA4/vJ3qrFPEUEGuYUy6+I2yF1ku+oaTHXecOqNd3eqSH
Obi+T9IgKvTaOnwThYzflU4NUEV3cA2WKWHUjm7tkcNI8gOERdijuVNv4KXChyIg
s250Ya+xtlv5HFG1KZZoOqSOhg5FBKdiRNoNKvw2Oisb7axjDSFryjCjSC9m/85N
h2OAzm+ztAHGf60+GQJoO8hkk1aqxiL9aIHhkhOlRT9RuhQb+PogYd7n5f3+gAAu
cwzrH2IJ0mI6EYnCJNhtd1KhR66y2Nqgpd/4fsVnaxQGnT/9B/Jg+5qR+OT2I6ni
5fsFYpSqu09r9+PGW7F3XIKJYTonHDj+QDh3ixOdHVwrDXpg/5/LGitbyYDappkv
INKAv9EghECuJp3yyM3HrNFgcM+0Tga9d0+lUbncHwmHcXeMaXHz5OkUmVrDN6xA
xxGn3pSBhg4bymkWYN8Dx+mWCq+r76hufHVnEmrmlh4lctPL7KcgV67wJ0BiI0G4
yAiLK4yT2orHbgsW70BUr/Y2kVmy4gtfyd8C4FySviKTwDg0uajGK9HIbmQTvu8M
5eyX4TEi0KJrgqTBVc3l1iBK2RT7umqsra4e38yJe8bzkp5aUtae5xHqdWUiXxNU
6I9B7rjMxNwDK+w/YbIGogFzwGxlpunQny3cmzUQ0lBYni1IiZiMi8zAzHnqIwt+
i94o74fLu5yj/TYcOrNxDU+/hISfz2e7XNKD/qGdt03jLfgW9SwGowNQow/vjpDT
qCymLADWOip7gXQnltYklNfu5R8UI17oL+++lqRXCrKEuHGeNY/Tfteua2TWV5Xl
WQ33BNHjpcdv0IHVT9NGrFxAtQ/tq7DL5wqCbSNnur8ZQfAsE0kGjE7u12DUrayK
5VVjgwEvRhnxKMxAF6jOdk2fU9597V9ErqS9pIzfRNvw6I+73mblggqf718WcCxF
BuWTTPDTsimpSdRLlFcrlJKoaoxH47vcIqcYH/tvE9U6oPJOO21hd6FcDi+q+SJ7
r7LBwoVlJkO5c7yf3xWBCaNDVJT/7moMMr7Ibd0N+ombtuYUEBTBvX6AXnJ5V4IH
Q3PzL9yxk19WL+d4IupYEydA5TUWyruTROUffFYcd1lhxbbC7rh9W8td2vulWw8Y
oclTL2/T/vYfFzXNhJMXJ4AaavfyVzORVMIUJZpRlZl0R77mBKwbET58rfoiN7My
Cwz+WJVm7BaTmgLYKpbMbXvfwFlflqCKRSWWbeTBWgTh+Sar1W6EVw4qy43plPUP
gIHw1nHQACayknpDBNlcYwtlWBMHxLnQpD+a6wDgXNVcjl/R+RCA/zh9GScodudO
Mpl7Yk5FpKlQEkYe78Nk+vvlXyySff4NLLSjWVLV0mNRI3W9yvgY+hy0Ozfwp4J6
vWKZPhJX+P/A7t5I6wQhPXWNleLMlRYQsEcY7YNGJ8zoZpNgUFTtS6GsA6kMalAX
mjWqN3M0g7CcCovIit+RPKtwp+Eod18QoxqCXLQzCDF3/vBFoUVCW0M1agSi3X1J
eL+gleuvkHPTqhgR17TW0ufUcHeK5is64sKCFtJvcdnw47ttarftUs+Ov75GmQN5
75yxwQ3LLxnIDZ3BOmElh6hB/mAysXNBJjHJDilS3zni+nwVGge8zuDGCqfm4e2F
cS7cIdSzuupyFzUUw9yGSEltjwYyxWrRWQ0TjKkcSn/9XjsnUy8fk5ETL8Hk8C8p
k4T0dA9YZy5axoLA4a1WPEnKDgKEf0RxWPq6ZL2mPZbOsfp7gFklVBWo5/Ybpmna
sHZvAZa1M+aLen8MghrAKNAgaaAzFhmmQbPJchV0yHxeAeF3/3hwn3Z+Tki7gtPv
xkgGiDpSQEFoo5yvi254uekDKO8cgfsZaoo9jyyHuREOwtTiYxuoN7Mt2gj86nnY
DdfZee5nL0ZwZKG3/x1cW1r5E4uMMnaBp6++NHGqaEZlFnrHB+3xvnp2bZdHPCCd
V8qP7BZjF83qpNXJIIV2v6+02jRz6mK4tbl3XRYoYAKx+aqvmQxd70vSeszfxazr
XvQyQVoob2hjHWjlrR0fKR5ik6ETypumZ9q+nmduxj64K4lyv2T4IO13Of6FXPmk
nN6xmYV5HI/ntGfrKhbhch8fry+IFDzRvAJSBD2DcqV5c9DwWR5PRwhh9a375qrF
+oS/ltwiTFEVH/A3ZmvIMxMmStg3uR0mKgGJMKAxb5bLBSxqx6mVbSeSxUK63l8k
NC6a+dWLAfboKGBSbGrElij2Psp17M2BJgpavUNYh2iFmcnd5xOOPIm+4gEfwIqu
tbaU5s06l4Lrs3BvkDYFm4eYH8kjieVe6DGHx5xkru5yjr4hx6/73+3yuHk5v0Be
8doPYZazUOcXkIORI9LRvm/BP89jnKukFEszP2TzT4zdqqxKAmNE7Bp4wTovuajW
x1JKILgykPK9UUVDqhADYJ5ZlDz26n26uWQ12q6zGOohFyp/+6uLVqU/yD9DXnve
S0fFc/ivLQoGg52Y2zPUez8nK6Xpl+i0hBTAssD+iW3N639UwI7d7aMG/4iPQh5n
78e365o7vOOPGKry7c/U/v+cCtQa6C2TloUq0TK4uq3kaHtlM8OQIKLEvOFwwzEI
ukN92CWuSlmvCDwdafC0RVkU2kMUlue7ptzLUxXCedCfHKwekl2FjZKK0XiOkzv2
JV9YEl1UdZZPelZy6cjhPeaABl99FbxV7PbzXMzpzHNI7utMLbEUjg0QlL2hXWge
KT13VlaE2o0jhTJDh/TD/FRAIjL35Kn8O4Ku0CzKjdZsyE3hw1G0yGOzK2n+eJjO
DPXTPPnTWQJs+ZecOFukzRFBvr9CAUzr84nUuC/fi15bGi5n3eDB85Jc8P8VxS9g
x8oUA4wgOsw+zo7i6FUw6OY8grnV/1rIoC8Ca4RBnL9u4CnHMhlNfAFNJtB09MpV
kI1l6+Bg1XKhJb0k1VSTfPajmTMO1MB9Tj2yktIeEbQJ5UyeLYCO9s8VwoQo5SRq
5jZJ3hRlSenMIzoQXBW+1mSNKfUfeFCfOLMtKoLs3DWr5psSd1s4+2xB2VScGl5w
P+boCbhgIHe6URkYbm19K6ZeZ23sNj5rzJDhN/+yIIh98CunWivKwzZmgfZEU6D+
dq6OlqgjY9M80XiC++rFAwj2AepSbCDFVsi97FTQVshidGFHht1Nr9UnUVT2m0zg
jfZmYKlPTb5KuumnRVKZ7Rm25yUeR2VoBlRanRh85yoPdRojfF5sC4T7iXX/HSJg
eU5yZ/PT7CGVN4zBdp3M5+PaFuFkgVCV3TQ85N/g8fjBYZrfB6Y/HqIP09JXBOqx
2Po7IvX00C8S8aQTrCe8GyxYYF4j2OghcT7i5nxy8Sy01U5BZdss8Q7w49zaJ3av
dHgA7wWP3cctWDlqoB40KA==
`protect END_PROTECTED
