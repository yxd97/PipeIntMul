`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Voygx7b8+SA3oaHgp3IZ88JLfn3sUtj2+T7PqrQ/PYgsBBlAKs7pZMXkmaVZ23PQ
NW6mdPo1/285jgO87kRfmqoZwV6Hnhm2Ax/DJ2fcQMHT+fC+6nRQU7nkpcf+YgMl
glNiQ3DrZS25uHtRa7HzPMZ+k9Ae74M7KT1eXhhcyDKt9MGcO98pM5bYCeDsejGE
lrxMu1rRyVYBjhMWCnSR9bf7N6pMV+Erovj2uz1p3sX3KVnXoVOlC+ZrmkNkebza
lJ9B/S03hznhEOFewChuFsPIE2741yFvk5yErHUEReP64GvDoX+mUTJAotedTGaI
WKuqPPU8P0tY9HEg185pUSPqUFNh9gYOVg8O5ng0RHNrnLrqPItZkjn9S/8abou3
Jr7aU3JOYHR8VKxoP5IbiYDtjPX2bfAaG8zGo5X0tB+3A/r5O4c15zpLb+gOAgg+
Ao6L7Nwi0mqi1xFBD1pMrZ8C3jdhhZfSkJ6qPjo/dha+Tfe46zxSRSvns5PWNfj0
n9jwWVV3UA9EtpI8BzcpAOI8yeNg5qAxVPLySV5eON0Ym89Te4qYNqQ5fx2KzZ4X
1qymTPj+QjG19aRMdcOjmjiDHBNVebLC9ZbG8StwOO97enGboNUnGgmWikiSCOoO
t10aAiTixww1bFd1C2xU/tbTwpIa0KxIXWSOrUT2d81i8HqmeRTsqvLKxpRpJeBY
jB9aGq4n4IzZ+xZh4cXq2+625aFgg0V98yX1LtvkTyJNxq+yAaz1ZJisM4rcL+Oz
hfU8hrVt9pDKVwptCitAUvLAH7KOGxjRKl8MQZwPm3nBv0hXUzsQ1sdHbmn2+ZQJ
dxfgTiJ5WoC/1ju/JXJ6PleVSgFO8oYovRp5oGDeNyPMNJpK1uWi+Hlblx3kWILB
GmK5/MTjra00yY0xCiqs7LdP9QjGV+93d9WaAejLGYV37zp3eh9moBA0xmZvVuhl
dPhxfeUpI8PGnvFPW1hoJA2SsmJ3ZgruWqbud5V934MFybMsRD/wIlXf/PYmow1K
ueLR0idpHsITkhYOR7rlZSPu81ZpASnuJhyrTsgCJz7zGlDyDTeuPCBE3UoYCV2u
GQR/HImE1+D4OIu7KOfF/1KcMYNnqnlArPRXLHmJUjzUhDsTFmoON1xur+gfUSaY
2sjBD3h+hp5u6VZIfrBEoDvRdkNIvrzDAxltrYOKKuyZaXlnBh3eCZw0WEdZfTEV
uGtTHNTw65SVVnMyG0ywk01hrqePmpJH67Visqj3Fr7UzXYWvlch+KNpZA9yW8kT
luGeoTfgqyFxzvIvCeC167/47e4chubpXFHNCX5hGeiyKyXqqAVsnqOuphsDx/Du
4zRAYKpsbI6tLos+rqIdKbMCwHVOc9R0MCfmqPP1tNrgBN5YI99nFALSjkCo1ytp
DYOnbKIEq782jjfLyDZV2SroxqEorLw6jGQoyNTT+yZClNsNfyn57AtELzsY1Hu4
v8GHe3oDyYJ5xjttadPoubqgTe09C1maJDN9akIP7NxKk+k8JFykdjdvS+H2xF7X
GYBjNGvO+O/VvIunK9IEwp5vC82tLy2tqJtgp13sR9VyqsEseO+S6qAVP152cq26
f/YdV+/OcfuNlJEaUpSsGbt6aCe3D5LcflctEflAaQjIJNH11I2UYJ02zWJit8X2
5X2iT9PSmdPbzElQOo5ZJPOnNSVQv5NL8QW6TsY/1YY=
`protect END_PROTECTED
