`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NUi88eDg8bp2H8fO/J+iaizBaAULiqNzucaaoYFLEgePjacIsylU+Ys07aJxBYwS
HAWIYW7TuPiJt95BaD3yTqNr8LXu/vrr8sCfcJQHvU1Wga6Jkt+Utmi9QxShpoFD
85yWJ1koV32nimOV5bI4hzQYG4y/79weXJFoeAE7khFtnoe3q4DmFLVIEBApY3zu
HlnColO3oOZY1R84gJLYzy5ZfqxX/y6D74EAKmf+LZ2BOwVLzQiIViueKAvyau1G
VQBUx9ELQC9KdCgXDe+YMFgRM4Sif4wCZENnJLH62W4fj24gflhVX1SgMAvFFwC0
ravgj0/gnAn5k4DX66dp/DbkiHXs6zan9vxFM7bdUYcTuqPTNfWF0D/DG6luweAp
eA5e68HaW1x2wmMepJtbD4XSSBZ58hfYd5YOlSNmg3AheBSgFug/AjKwMXO5t8gl
yD0oUNKs7M3buX3ASgMIVe8mA20bz9gpdjJ53xDDAqoKYO0Py3FqlE1rWFurkbCX
ELYQWZdDec0XqIyqAomNbPplfoy+XL1bGcYYRjXQAhxunqvggXtGupkaa5qWmlXT
zMCr9CE3AQOaaDiUGhd0Tr33Vlwj4cKgtQbGe0jDbiTM11NHBnRwSYhFHRxgk+gW
raz6vWuV4PBkKy+k8LqeA9PcjagkqqkcyK64pmK1ySnABnnhlR9NxAikzfEqdWsw
H2kllD+9GbeuWgbAWjtiRt3tDO2dsDJ/8+dS1ZIRsmIslX5mFle8Dqem5Q3TfwR+
GLXyhnYUkRpkvYtJ8hhfsauDo+Av4gL5O2iH2m8n8inUAj9qPEsdKKgAGc4FngRK
i9aiAeyroCtTUn/sRTLKVfXa4q3kjZvBn+0ZKnNrz//NLQSI0oyy1+kGierd4hRc
xWBIOgtz08SBx6RVjjThrmijaweInf5MKYoLte2rL/LNkrmmju4GEtM9/K3icmur
BYS3JQSaBjhbXDHnastPj/zJQEVTCg8uXJOUi+x2hLyo2E6hcAppw69EBOipJ9W5
k8JVzA7EN9j42W5FCmsuRG4VUORh6X1bpTDkBxSgx2rbwLDMbVCyafyyvzrSLeja
uFmIaVaqhACP+ZgFov2d9DqPDfK/ugtHNXNqrZZyKTb4aMt90zMHpdFeUuCaGtxY
cWuZ/2SMAKrRw6ABBIZb3l9Awyu6JzyLUZtETCFe98nxFT/xyAg9fgWouCwro/qq
U00aJDFBVOx6hTw2oNh6rj626jBgWajzxPMdNXish7lCZJT+6K7hIoLuItNWk+gy
wwJjCB5c15wxbgzXrq1+XzYOxAQNFsIyV8TEkJvIhfGoBvVe/dBGQ6R2rkGrM1Pn
BlVf8El/oaZhrZKq2b2ALtM1MullKuIGMz5apbXuojnb0RmV45F9xU9DY+a7NNdN
9uUKuacTJs3yXCP+cINm8SaOtkpkF7ZfkwJOZA5jTOYrwVAknjpKKfR5OrTEsdD0
Jy0fZs6f4YSYmnu6CXIlMRtdEgvOzgqY09UVNrNOfimRmZoGjsqNe+zWr7W4p8OG
68AVUhGw58nISt3NuG6df7JtcnX1Q+bnMo3sdowrURNpX5bXmhnctVH2eoWPQ00O
H/U4fHflrJG6NUO5DoPeZDDb1wzzHejAJ22Wr2xVW6P7bdGrd/N26agJNtw959CG
tB2mHQodCys2IGTTTC1WDl33KWZ+LEP27iSHWlqbk5gKeDG1uZL5OI8XLfZwIMpr
SNMjTEKn4ftcQc5N6wTNp8zbWue2miJBl+Vq3DlEFqJXbHIfmgTZuUEPcyGJeYG5
NeNXOgk6+b6/fB422nSl073Zu1FlEGZdwmjXqsGdua71L4MrY/j/GBgw2AS0ZTjB
S9IrKHwSWyz83hwub/KBNSrod5vn103mt3k5NystDV3j8v/QbxNGms6MNL7LmpcF
SEIMW1YMxmrVFab8wODWSEHVuba1XFdAajctmfJ4sw+k6dhZKyqASFxSsSEmVzCU
a/EhkVbOHRIRqNU/KdxjHKSoDwl5YnCVQE6PcR9CiJ4lggq0yeoFtDpH8IlCrGZp
`protect END_PROTECTED
