`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m4+j8J33dBbope+Pg2B1WUyprzng6035wLMT6YG1WB0QvhBuBIzkPtxaxq5asNak
b0Ay1uBg46q5q2ThRja3pQwvkWQWnAsDUa1fZL1gmcWTDlQ6OCWO/nnDKOgKBQ6i
NKtIYkm0RMiPYdIEYuNcyO8PUyiWjTkkcEPJDM/VQBxq7gOIeP1kvNFOW9vqRHKe
eMYyvy5jG2pBoO6nQvJlElwsjpouc3S+A/IpUQUyD6lzkhlAUNw3lieMjnDvpbCD
euStxZI0IEXGyn36Or2O1ABNbcGg60nhys5mgJaW2hWM2P4zMy1dMITWnuKcKMNC
n2PiaHGYN6KiyX3i8/i7+SXBq7iSf6otb9Emt4cSgfhvtJFP1UjMygyqvsZUnYDJ
XoMa78b4sOsdd9J/UzYFh85gsQ55TsuZ7PV1vIOsM4/r/n8PKaEdjgWrfCZN+LXt
44KbQvlVos7j98ILICKiFNAnKo1SotRY71icbVZMW1B2JTaiVvBRNXvALu5edc4q
IlhnEq4Fpzh9fdaDanKPIAqHZ8kzUBLLYJUXKbns9xSGQjTm3jvvc+vnYWx7updg
OxOuzuRgbyBNwIRWmIhp0iv2Y4aDkmNt/lSiFg2bJIyB/3GUClIej9UQ5tXgQL5v
F3v4K0YNL79HTKZPRpmPNl6FsNuB5WxC93QBKM7czKUBCV4lwuOsMK65XFOjoIhi
xYqIye/aoY4zy/zczoWAW4hfOCqFuL47Kn7d1O9FvgI=
`protect END_PROTECTED
