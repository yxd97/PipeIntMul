`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uuqs3msv7fKo+KEeDpHrPipHP7t1cvLGY315TI3Q05IKqdLQlyw8dH4GUVdDuPs9
AqD2EJLRWMcW7o3qLcotwrPg2qm99HgKB9RRgqEUMfl1MY7AAUrVL9n1MVVGNM/O
Z2aH9tqacKqpE6wNFTUfgxlJ+bGn4cDdBZiz4vYlylaMmQKkzyR8s2YiGb2hr+5/
g+zNUmGAX+I5uJruKIOraoQKVh0NkqMtxWM9xTSSxNKtqKWVve6COpC/KSr/7N+Y
KQFMtcmYHJHxzHNpzYULiVHfiAMcFQl2QirPXN8TIcq/G9lyzC5aAiOCqtypA3RT
O2iH4ge8p1dgm5bKoVh7Fw1qVSPIecRTh0uvlNMaS+t7/D5LYbVIXmEFfsZXS0zf
ZlOQU2PDydLsxvBHHxZREINYsaYW6yz8yjWujNaUPBjByI2MVcvAI+PTlrcZ7ZyD
ta7Y26TYBgVa7v66o+EOtbXEz5zadtM/mazZ1qHQyy13dVH+7A3D+5biNdxNIqbu
3ep8m0DQOTlGTGCFhAVwDc4qQW/yO7vJ4KrDZyvn05cLcqWlp2SSPjbjKB0Z8cEu
QlOmv7Io7dTbM3cnA8qYgdefOBRy/jAf9St/DCEFw9RVI8gSBRtBAtfcnvVtE3m6
doZNRTaajgEUl0azbSbOkbGdaBnmdrSdHwLip3vn4Kqcam3UDilw3vi9tIIwGvLq
r+qdY9lUcHcHNP1bJgHpkrGbA1T2NM5g0j5yyrTNeRRNOvP1ORd9hju1JvSCDGtX
4Sh/RQ1QHGS87LSsnod6uGCIJa3LNYUwKvr4v10UBfY=
`protect END_PROTECTED
