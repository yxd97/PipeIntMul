`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yi2x3kbPATWmtn1yNpHQZLIi314o4HOgMg3oNJaYrUwr1zG/aOMlpmWrd1yq1kZL
B9iBumQ+G6SMI5hT/lLIjSuB0AKAkJEbMydRr1j5Cpqq5oIMvgNbmfycWCuVP0K7
jSt0pUcaRqmuct0B4d067F7ZYbXQKlFvIk/odubvERVQ9DOQHVyzPZj0165wIrW5
Mk2yUIuPEbpYbGsmAFS6dr1Wz8on3QfyExYdMiwD0mIzAqIrMdyHzM3/a7UmAsi3
DlGqlAH5PnXcCECNdRJH6ftP8d/grAXq7YITROybyolKZPrFQbVrWFvwZUPRYUhD
V3t6Gox7lgASXTq5PWIlAqDuAm0i3z32SfkS9ZmWExu3cp6gfCjN9F3s04PUdwHv
AmaPVjmMYvaLpOcAFgrw+Meu4ioQ323MC3FaG0Fapc9FlZkUvscsMbBHao4W7jFB
mgqQLgBaJ997ploQ6m3nRkAGo6CuoTK4klnhlsBnCGGBadYueP8wos8v2ODpMRq6
lD/kj/vi9mfL5rkV945eGrfYBb2aPFu7QY9zJSWObtf7TL1V52cpKldwj10UbFwx
PGFTa69Yg6aNDU0GI+Tml6FMXp8vEf7xfrq7/WT9gB/yvfNndltD0/NX8YQLFR68
7UzgXYZBuZilaJCFd55gknPe+tVs2B7NiPpUa30KY5f4hXH3jgJF31c0xRQzvktI
njtzZwlPKroM7+40m2KN3xFArS0RIJCisocz6XHDkMnp9rB7NL6552rDFnSQp/If
x2hgB2OjticrrW3Y9qMwizhdRQTROUIPxVjo33FvmqRBQX9MvTHS06MtXAddaGhI
KJnVQtVzb+5rn1IGnE1aiMucQLjlIPbByv4KkgzhoAA=
`protect END_PROTECTED
