`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+nTf2y+QrnPENMxkX0RDsz9C1Kxw+ikgGGeiLBZL3Q9q9LAce/+vXhpXtzNACYl
LUgF0pHeIfWilaSrnA/rn8er0XTGD7G7g8aVx5kf/Q3ok1dfPXwIRl4UiJAqXSqv
s1F2VBcjh1zV1IXq7BZ0dL7Wz7KZWNV6mOQxcQqNOYvYCNf+RrdaULzKkIEVPdtD
9ZhsOp8GFVHtNCdC8kelXssVnNt+QteAip00VEfoYfM2zSkmvOjuHr4lkwOlWUBd
x99KPZ0Od4+FZk3siOoAE3Oo1LbOisXX3oS3Fd/KnVXKjGcT6TZgomdWkmiicyM2
dtJd6bwJphkOWK94/evpwGejYYxQ/EJR0jufsu6x+zp1CPkUkicRboe3/DOEpN6u
xJONd7nJtVAmF1H+gHK4PCj8wrE/id5x03WSpCZ9ISvrPzc7YSavvD5pAxE6cgBA
D+WEwj4EYyaLGs/T00KrtIW8XEbz3kQoUoYNBBFQMRhfhjMwsOptfx1nplNgf7Cl
pwKC1vT37rUV5G1g3FRu4mDayqSZIqfQt6ZWvjBiDJk692wSAujiGgODl/CCH15D
VKTwq795A7zhhQ4zWD521Lljl+pIUMcf2SQ7d86g03IA4rdvGkXMwcsz2YyC/vsi
VZ1itO/8+tohhOGYMkEReAmGAFxYvSyBWvf/8iIenKKJPwOBRT9oOr75NDCEslHb
FxxphZ+9D3gAnrYBSLkldjH9ckbKBjP+obJ8E6hFt3X0dM70mRukpKdZfzDhu1RQ
Qzy2FS8F/KAoqWfXq2bYHrGyH0cE4EW4o1XhHlxDpiDzc6OAKAOPziU+nhMkUYUi
Iyl68MFmXPqLt8DGv8HpFH7W3Zw5wJmQ+eKAyFPNH7nl/XqLO2UfUi1ive2kSYEn
r4en8HH1qvHCblD9+/ARxQ+gsj/qdn6MKCOgwwIOKYh4svj+quGCuMdNtrSnN3LK
gOtpBPaWInalXvU8szB28io+JQr+9U6rwEYVaaEbAN4Af3EtA8v5IUNWgMSr5Gvq
pHHuZU4z8mydXMZiUYJCgN+4ST1zKoLsS6H7C/4n3MEADZuk0cFUUKYIVxYuGnRb
uVAHERxIY8Kj90PyLmZQfwUrGqTTZvX9jaIT/1JNLKsXVD4icGaDqfCFxawzQfwV
hK6vFuiWhxrVK77dH+KJQLMg78YXhhTNqIotZtrY8qR++WOQUUtCpt3kxp7nNigL
8DITMPYhd36Rvn748yc9oMslrzkXrAVCELXIWyFoWZ/UqBZ02MhNC3J1EkIY7vGR
88TGSETEMcWBlpCfkBHVvc4qkyadmn9RkI0KVVvH4ehL/7nl+cpN5GydixJnKk7n
8jRaPTad9s5veN3fKznRRKlcHuppySmdBJPneeVDgXFKtHd1Tuhcfhsm7bD6dieM
QtkO9sc59kuZfhCB+VV83NlCUsjTW3a0jHrewDkNYfKx0QX6RLXyr9wmMPQhWf/9
3PoFT9ThwNKM9eU0QOh360Q11sPlsJKftBfA2Q3QAeojgccR8YGJNMzjA5nF5hcD
ZWjhwiKQs0KTgkEpABMPafzqAbJJj8WHMFUQRSbTPzNBo17foEuok+tOpdBP1EzR
piiad0EddGUQKdNzZR32MLmC7JKaKh/kBEvVXykuG5Aqq0vvSzsenq074STt5VUZ
islsBv371MfbKJtQWhJ0+B3enkkhn3C90LZOBNJSZ5psynNQfvNEPSpb5cqIJi32
d4VjYgbWkkD4L1hxKKJjrwg2D83xeDjOjelGTeRCkbYZDoKbbrU9n2HfTuCMdUai
1R7Tp4EsvLbCPR4jRmxnT0PtlN3CblAvyeQRCZtzY7NPbt9W3tWbBPj9mc+uPJGV
vl2TdZtSJbegnT0Mb5pY6TGRq7s0E2CICK8bmU55VADE50CnSptMZ6KFj0hP6zNE
bGeCbh+PuwIdXSu0O5dvyGRtSL8w8lwYGIEg+YDAvGbNZgsEbnT4lq1BKSI/7WjZ
MRgjzUCPHBl9BlD0T+1L54tG8QnX16Vud6JkO9hjHRgd1umhEm2YnZ0L3qah00P6
f/lhD3T8VyaTT/z3LnNB7o4GatU/fLVnVzA5rcXQlqnNA43YUXJW0h7sXpUmCaHe
F1iQt9pvbOIhI06QQ9QKfbqeyR4myEeaLYF4rt0AA2CcdyRLpFHLmZQXN6RyHktd
nzvv9b+s9spU+hRy0jRsjQf0TAaje77r7a5CLpA+LnwEc+UEMMgrA285IHoisyD/
Yl11YC5JI+hQSIR+RIYKvAbCLboGEM8xjSpd3B/ebTbKaAoXBCxTEHd2qZ9BVa3e
HjqwLfRTDb3DhwW5xiLcWpjhBbea9sbZYXPMed6XXreBETZ6SfzKWiqJjpbc5iet
8gpNoTGjyrudW7sq6r6bs4iC9dvbhNi5c6pFp+tNNLJPv/YP7jDAvLtuJpfwRwZN
9/hbHocbhNv5u0a/F6atidnx5jKPJPjNNZ8DXanXu6fEDshlCswvEfXI+CYmDxOo
RZugQfcXY8Py4GfU9JmMhE1faH6J0TjRCXkTptM6unyqR2Z81yWEPoGD4U/reiGA
tNAlv5PLKdRr6m3gh+QnnM4NQ+Gz8MK8ELJNOQzLZFFCmAAktJdkYqpwjhQ35oA8
QQFb6W9lnrj1Sg7BXNOLPQNaHlRDXVzHjrD7c41czOZe+XclvNtEdJjHOn5ZPf4f
SkBkpyMZs0ldS9RcOaTHBsLICxMGOJwzUQyNZYuEPgr/SXDS/pUocTBh4yfPFPeS
k7AS5cy2bQJjCdS8hopqrJ9G1daXih9yqViE8XcXSdl0q13rWrmGMG+ZuWEvR5Lu
oFeCHlUQQ1iaVvilK/Vj6WLHcz5Is66PEG/jSAywAxsErXgLcPTrgIla2XIjiwNB
smIobCh8/8vS7LBed5ydzM6JN9KfKOgTNCfd8nVnQfLv3FcXhkPPaUxjKQ9YOZsH
XZO+pOa6gqqf5ScpgaEgEcrmngEA5Q3aIhQOwAbMUfReRf8w4ueNAEM5HPF35bEx
Trkm0g3ADquNoyYRZQ/nA/T7xYKSrS6KRsZHA/hBSwfup1llpT4eDZ95RZJQcvei
vLBrwThtj+5ByXIcRjHp/7bq0nDYEhKhQwkCujtEp3L5+9bwTugC9Omz/g8H8h5e
JI74VcZrGct24hIlyP4l+CSFV+eNaOuRrRz/Y5VDSeeoCeZGOHZxoPO8HqYVHRJ3
JI0rCNkHxqwebp6xs7bokpOStqPRFQy4xAHAmFUDMxRjuA4FT26JvorOeJtgNzba
yKIqF4cj53rhCKrWPTCQinYX3MZvvZ5/Axq87WFxzZVABBnlcL1f0wVCCqFSgWar
Jg3agvn2VozIqDLaAGEN8QNnnGamSRUK4mUVv+02ii/xP+O4Ww6natiicBeI7jrQ
QaizMSTpnBDEh7roMK+oHehK54FSV7Z2q1qRhFzA71vkfGvODfhhcxewXvCmoC3+
s96DeGeIQ86yBPeMA8HXmUNt3qQkzN8MT9+CwNvofPQv2b6prjjuOXJbu7rw4wXU
5zMD0BVbU+1XmfJ40FyBICob7gQSJfMjineNd0+M8Xbfa7dqFSHP8KGISU0nojbC
B8m8ZGsR/qmz35zT+jA4nQeiHSopyIOl5BvxTpLj68OBYTOmbX7JKmE6vB6UcmDI
NvsX6Vsgwqu99k/iRKTPVd7xX8jqVghRENV6//h+jaE6dm3R6mL2q36QpGRevA6W
fFC96SFqP7/7Sebjbi1pkPkOc/dksskUwntwAs9gohoJARw269UL5rYWBub6hm5u
F6vz0rnPgZJpilC78+RPojmkzO/Adq+l+9XoGipSd4BD+KCfd+a1ew1ZhDmTcg2B
byo6pfcLij3iVKLOf64lw/WOJGOaZgjx94xq1f8+p1/vs+2IjymCiCVacOYPiA38
ewQvmib00tVAWeRTDnsr2Yi4FfO6cdN3kkz8bMloL+Dvww+GE/CAHU1eBmT+whbw
cvQJpJ930fl8kvYparqXoSAOwZVJvvq9/8WOsi6xEnmEynScalVlEaOWkDCubRA6
ejQ/X8dbJfcYhpI6hTa2ohbkbIS/HXoif2kU+MHXCP2eHB5nuwF6o3ZeIThFi7+H
50J9riDlzzwXZGXGO9VYCxL5d8Nx8PGGyChRH86YtuMbWstXWnRNS/fFAjjoBSuS
xALY2Cv4HxiVB2r4F5ESvL2LdEG/x0OGlTJhCT5dR+1WR8HWLHkbdXdDL5BTufHL
Mfpfd/dHfYQ4k6RD8v+Yl43S3/RSSeDZiKF/VjyjDSvvDxK0QEC5o40rXdTVkydI
dPWXHY9s6OkRBm4TlbKCD7f7psRvAYJopaFCDQwgCpSQAwxED1IBjZZdImK7LqBl
x5O5142ZyUrcy+7T/xYotGXzpm0ubwddCYULMF1nqosFXdbDfZpWYbRjCF6mBoo7
lrqIfPGmYzaxmmJme/P0odWL0PJkNoQIg6Bym8ycwY6atEUd0AsdiIgBbRn72mRV
EeqJCAGUhrCsjzeRggYGZz7Rmj05d+FGBcLYbg6irQ0wuYwEwai7IBz6jT/bwLkR
Zf6WgPTwBQ+M3vQCPACO1vnge1En/1/uNfBTYU1seJzbSa2fqfFjorGDVYEJA7ub
S1E7BG9Mmv1QFpy/p1r3cUejsW3HCxrnOwOpP5sUxaJJpXad5lHFag/HKAIFHkG1
05cXSvrvSnlTS2n2Tk5IRzxq1xZ/VWmSGn67As61n7onPzYfh/kYCbJzyJeAmKpB
0bbk7m2e5qqGbYhhMqKw/7GlatXNmQ2IRXPb+OwfZf0bUs90/CETh/GeiceQzOT7
pp3roUskqCkOaBoWgZWUsr9qBTBM0MguA3BEdy58VAnlFezqQuo2Q5f6j3ACPQtL
MTH8A0Lz/b0KKsImO3g/KmVM/7VrqTB40z6rFdMhVQj8WSQujQe0d7PaBiBuIYag
7+ZMopEgr86TJls1AumwwNwXBpbE5dsNYFHqaZuxq8EzvzKGPnTUSvdlSlCRsjRe
zk+O4007CyN1lzZbAsjg1O+46DOarPjOWFYvvwikRBct8dmu0xyVGwmzan9Oyfw8
pCrDkqIHS6R7rFBZRWHZRDccMxr+fFlCo7uIHKuVh1/jP3NLONJ335OrbuAyBBu7
ZbicDzHsJqfpGlv5temrVMMsMUjQWYBXMLq/uEH69tbpHBZLeMt3LaTUchXsUcuo
aHXLXAY9wHcgdWcIYROXmNC8zcrHmH2lD/eleLjqtOymIj/m929QpcrRSBzzAYmz
p0uxkQK57EoUCYkXgZZmMGT/d13so+NfC/7wgkLEnr/D9xfFbAfA0FZJys+rjzkh
V39lFbJ95eWO9LzwLVw/+f6pQTDhOa6/025ncYBHr6qfdc197XmybRihUWq9X4b+
pmdqCoDhjGd/IClATbxWNOfSf18MB+ZpXs6hhC0R2aVrZeD8OQTFC+OE1jQdmlsS
zf0KHKYKWpqiYY4SdQ/M269HHP6jZ5RDen+qASdWp2rn2pvZsUOvzog87X1/3aUC
3YNEPuaWBCVS6X0TOFwmI9FF/HBkcSPxtECg8SC+otIXzIBGGqaetwytP986PrUN
MIJlF61rWugT9SJ9RMz3XovwCcchIJ9AzU+9C0/4kXx9HV1iwD63MBsOPETlUWh+
H1x5WHGL4WlAKOFOlPkkUT80MEPnO0RMaPpMozZpX6mrUWiO9MtPEi2sFMiWnH+j
GNjiULlnD/71zutjQUJm6Wa1Qh5NEFNf4KbmdUFMqZsMqw0IV1tGZPKI2ms3Xyjh
inVrIDvAwwcw4SxwI/4jc6P8ayYblRg4zX3l0IhNfhkwMGDAu1QUU5jT/qb+myNg
ayHre6ldlBoqGG6Jv7f3rr3MQ//FSgEDrIzGK7m2BhpJWUD0roqLnqs0qecRQ5dH
AFq4cneqYI23QkDdUXPvc0yXrjK8rPP/b63CF7f2RFs+ZrYd5gVQeIRLJLF/uRrs
gNAdhdCA1N+nUv47gKL/V266gik1nlmJIlGKfLWZUM05bQDmZDjypUbG+S2kpJm5
IL51mY8ZAFjKVWMIDiWAktayM0HddhLzj+Zp3TOZB2yyH0DwUZmieCqsCkranO2P
iLIJEEc6mT8gvdmCPhd4r+o9R1WXjHQQpRIIiU62ppl8zYf1B/uN8y9VHdy0KeFH
3n310GQj1qqCjZmlcOsiZY8kt5G4bU9OuhvrZi8bS3FobF/ttvXRos/DLQ5lUH6z
x+ht+niAw2TlnEryEgDmR7mlU/2cwuM4TQxyd18VmuR9msNLo11LeDwfZCe5giWO
moxOWAfNJ6L050SlUFrIa+kB+uCWQT05VMHfLcTzihCS51o1Gzq5Z4p73CeEHVRA
Kueo+ZAQavhEzCrEwXPvNAQLfywykdSvEisrp0lLv4T3lIj5QXKYuzhRrPbGpWPe
/yfh9i/gNOaxyttLlIZzcdIZydhHFygo0LbaOGmVCFLgVMBHMaP3rRPfII0e0d3g
AvyjcNb2pqXQoyQtS+FnXkwLtOC8FUC63QHUBfAgYISYcXRGAW9OtKUHTJ8jgvAz
f2fOlTYm3u9R+T9q1Wsxg19TaFduspMg9pWW3MKt7sU187Zt1OuMopC8EPtY7/tg
jWfPQ2zrEitHE0r9oR+7tIHlKm7U8qrUTgMC5kIjcVuDqqfIelfo4AgabQ3XK5ee
Xpbq/5mBNw4G0WmtzZIxUz9giA9hTjj7M82zE+g8L1xGSgl/lizr+TSF2vjjmB88
8FEsiv0VSnqiyOZDXNf/UISVm8zEZuhgbd7LRqwJD9aFBfYuZL6RFvPWSLvl9G86
bPxUl3Iyok1hDz1xis08x7nR6EVf481pMksr0mabvZji+qeNgIWkgMFFwfu27yT1
HnB/zVlpn3rgapAuQveqa+rlD8xq/sRMixmnSXGIIp7oLN/414pZ7cmMZJOsTrKB
STSOIUHd61hx/+mYAi8SqXMr24Z7tTWP98Ze1wLTbLgJtwPApIvwZ3C5f1JWwWhi
Dbur5IFOo1OJWwIblvqWlnf2271nCsiD/DgVC4E8jeUfns+g99nlhitzssshk4Jk
SGkTWCxDo4PNoVQzxpRiHQ0NLEtOTQTGjpQJd+GypTT6Yp4fKkZCfjCRAKXgaHX0
Mo3daEa9PSCyWUOLMqTuTEzhm5oFoIG3l1Tr2HXyVsO5A4Lq1917wCY8PGvyJXWx
K4Krv1FOl28tB9MFn8l0XjE5uJcxTMK5r6rX6sRXonD3IEW8+dC0tTLcvcVgQ7ia
mq5rVhtgj6mz4OdzgQQIT9CsYTdEnpl0q7K1gBUDD8uFBU43aYfg2B/4l09eBiI0
vWjfTKRsrki4AjT7LlAJJzvhUWZ5NOnuY3jO156WMwGY29Mb9WnYaNU8H5SK+tUz
ITyssZecYiprU+/FPSfsqeqitJXvQUXmHatAVinMCVl+ZvoO02gcvdmtWchTGPIx
gLHDxeijyIzU2wpjTJUN++n4QaXeV/9tK1ko/2+xlesRxTY1JHJvZuAxX7BABLM9
fvoo1E4jb3m5EM5mLNXco5qUcySILc8e/ZwnZdYLmYmdplnE0e1noaO5VAfnRo/K
oKsmUCTU8lZFsn5WCdSETfNJOPr54PYCEc2CNMiyj7/AnGithXT5oaiA3ase3uJx
R9I69F8tNRVuyBmTCT9Jl2TD8T5iRsOd0Nrbm9X8K3feGfKFD7xILxRN2nHQ2Wpy
wYM5doMRCrh8utIR3T/34x4E9w3T3Jo0ZBjO+vHF+Y7rwM9OqxnP57AF23rEhZhG
luF06aadjGhmRX2+0bhIRp+NKPqq8kWoPs5DrPPxUC2mNmRdNCvl1xI2JlmjbzfG
ZoeHWR21HRY4ikAsfEDq6IkdfOiWzGUB3Ch2TeIXcQNY/VNqxvktjfycZHTNCwMC
Shzjw+UNCqMCLl9Y+Jo+112N9/oE0RxNmyBXUFNCS7x7P7EV7gnZyoaqDQEpgKZO
91h+0p12GTmqdNcb26zwEV48EtzbknvTGz2YCA3/MYGuvfVQG5b2JPA7Cjv3CyaT
xmt2xp6x2V5rR8dfOCnJT2h992Hya/rF2jmDPqe8NvmScnXGKuHBMbFjmwtIxEmK
ETWXRE2adPVyQmUE5eCTjhRuFanmshJYdtCSKFglp2HCWdQkrMk674iQlbajTbx0
0S/oOQ/58+SOUjGM6p2fNpf5GpxfC3NMGuRRf5uuBiVcFvRMw81kIpicQyyH5sMG
StxXpYcKsdpY3aSvTMlXjVIINYcz1d0+qnC3Yx+oag3gA9LGTovMmKsbeywoT7gQ
U5xKsU5U0aRFBr7SRicxqLXUB2T+OHJCXaaN/oIo5nfw7bapSrPP4q3CXqk/chBn
1R4gYu6iL3WECfmAFdg+hYZ11Zpt0FVAtkwIoGhuVY/rRa+5BFo+ERXj8qKc/G5h
AlV4DMeIu1VBEfyl3pnr/1Z85r5BQuN18hIem9NNRsL+huviRDIcDGYPqkBV+5Xw
6PaJoWHBwp1nW2NkusAn9ua3tFhxVbOk5Jnf05Ej6hi2NK2HFdSOn/CAdJC5uUCO
9OamIDJO0k02Nj/E7JVMjGDjTShZFUQV//VyguQgTCDwLokRTBKy27SrtWZap0v5
dGvTvIBtCPT/E3Kvubb84Tl7heN0VaaNIuwJwvId91UOCF8QdN+vG7J8DC4WlNXz
mvMHrz/YG7sEGfLYveZOM4vQ+kVF28sasUIYz841xuy7Iq889r0ioN0zPMDzog7l
PJrmrxH2wEOWxiRmA3/t63EXFE4xGnaQ7zSC31NxAa7nCOqEhtnGWBkDZSJUNT4B
5hXUYf8Q3fYEswzqOkrvIi0AhB5R8lRCYRvdV2F6EPCVWHIXvaGvDhjJ6baM+xq8
63ZfMwvSseYWIGbuIc5GaItugkCBLX9vOIRfxvBD/9Ai8UNE8AYT1Dnjj4ZnZLXw
aBqZ22rSuaKwDZuFUEtwBephxO7h+Ki2wOcJjIxgNpBswsYkqKfJM9LxCJSCyIWn
h5VFICEjBj6sh651To5lyIBHW02MFkn/SzrS4S6zAkLhFTYluYLEg6qe//TXNQo7
h5rWHvfVi3w7LleA0JOriunpN95as5dT2hedsz00pEx/Rcu/R7JsYE7fVAjA9oy4
1XubfeC6tNXw5dg3cUZyQQKrUvoSL14EahD7i2GhKIWW9+elmGWH8P2vBM41t/pH
8AT3Um69x5nhJMHQzIYQpMUO/cqvY2PP3UUn+nvHYg3jSVR1+rQeHiBQn9BWMK+f
Bb88zyUUG1jnU7suHIW+3ct3Tqy1BGcMf47ebG5Lh3lMlanrs3z098e2fsJFo2o4
d4YwoIkkJuwAEvvRCBDpTalEnP3zlvycmLMzjM9i+SLUl3UCXRB8FE6DcsbwWma/
uqxS2eAMJmQuxfzn/lp3EwtExDhXLAekzdXN5o4gDtMjbFMyMGOmeor41G0fJFt0
0RmIbgM7u3sdtn5kGEe4qp8rUNi2ArKB68K00qDa1dXaO6R8GDnEXKfidngSzclD
UcHhmHMDXEqjGJ1BWdXl0T3FPpZpkfDTipEPlFj0SlicKQWltRzN8EB7ZDpcnkNF
XuG+6h9hN1XABU+S7ORSC4z+UxcCD7iw5+6C35Ppu9c5plDWjPZW18/VlXwbQggq
Tmgnyyl4Bz6GVK0Pn0zr3pnWfoUZfKE0PeknnjnJH12cSK1Dgw1S2pptZkvIF/49
rleokv2YqY5G0uBR+2q+s2lLLDpbiWjMCRlFxmhO95uUVOrvfx2S43pznDO1pgy/
cfmxDsmIhYWlD93BsaqavItwLyCirlyP6DmFWa5wXTZZhWmWGEDDFDDUQmIfG21G
g6FqVGz8uR4Zw4/hPgEWNsJkpbnpyZyadNZQCQQEwZLjZWwXnzYDd2bAhXaT7t14
bJjA5CZY+WYj3Y7CXyfWQP3uTn0+av0qe5OMqyhpJvtUB+AuIKLgQTMHxQavSEHY
ND6bEPZMVHET5QQm6G6GzUn/PeMD5vmkF320U2m+XJ8r43uHPczJDmXL+KePfAQR
Uytrq94gj0KhKjvNgp7FP9nYivL/KtUpWHBQWHHRKlt+BVhRjj98DSt9dtZmft4G
o2quw2bFfbixJQEAdGcYtOmEAzH1uVoAagQUhJuVHEqrOHMu++//EamNmGaJ+7CK
FNwedCUF9uaJhQLq2aTf0l49Cl9ECC7c6kC5937oAeCnpxC5zlX/MrSlvZjVA7Mj
Wz8M5Nsxp8dmNFc8UlC4IibaVFbbeVlCLwq8Iz60Iiebs3Cb7vZ8EPaEB5xzki9W
BR0tYNnRy+dP8AkayRVzLE3iyRJ1y3E5eHq3nXpwVrEibygr3mpNV8voIjHsTob9
O3pAegyjvUzhfaWKaeinelteb8np/cB++AHen7ZKM2zvv8P8tp7F0kuu/Nv9WQlm
xBBsQnKd0kMrr3fnBlzkUgsNTAoI/yNhv8kf/BXchDAcF7v4pxXACHYtpSLT9Dde
whjfzWOw667TeNNDxnINCaFqGpherLOHk2lyT7lqBlPOL5GCI8qiaiNY9WEbkN4K
UOqlAatVmMDNs0+CWyagdrr9qt6rEgk75MeTOLYkUrZrOR6/M1qQvDBplr4OO1Yc
Wk4gz9pJpsX11zP808jUJNChxB17ETErMHhUcXr+KPuUn8XSIZ/wAD5C0QHONFYi
zz0cE47EGhBuUyWbO8tjCeE1uaGgfdK67+bIiEc2b4+A4va4hBN9UaU/IscA400f
66/CEJ5DkwI91dJLq/esFU/5379KdSYW8RENLKyOekgql93rexHRcPgEynrLclSh
kX2Esw8lQ4LqcFUpCZ+C3amaxXaQizS56MzTubnN4vVbWp5a1s3EVpQXP7I1vzss
UP/cJrdXOtuwM1FVeUCWN/wGSt0/5PaXUeY17LkRdZGk7udHGEMFvLZ+4cCELqtv
zyn+jCiWVnTICeR/I00A8En9I0gBbKQlZrWV+p2fr0kYJwgZ3zl0InrjEpXqxyaG
OC0dGI8jCG+iU9exn8qPXHEQcmt1/TFA91jap/UrVn5q4piSiKsNwzZfSzsbNjhH
/1N0RPfEAF8Q1D/w9o88bmPziZ3bYFuCD3m/29kbux6pYSiwolULSHmsASCHftXT
NPe3z9ELgZFSxPoshTjYPrkhOvse+vaTpu3c8yDUFAM0jEHQzw4jHKww54n00QBj
Hqq0btunhNtzXvo5IemDRuHWov1oegLfKvlfNXAhd2tHnSaNTN7Oca8tBnSViYvK
Alx0o6Ifao/bANYve6jgTfsoecnyGq/e7emeXUWrz6qwt7nOeuRos3dV9DTsiQJ3
`protect END_PROTECTED
