`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZNKVfN+xP11nbI00d5kZsMz9CcBevcEuZ9u2uAcLtlM8Av03Lrz/sXFaN6ZWk4m
YtDjGAfD+xxgYDD2/ip9IkmlqKJFfI5W7rpPu/9Vqc83cwSlMucqXftJj6VYRcHX
T9BFZEi27UgQmhf8zwdniggi5Qn1kcci7e3AXpgNlxj9yQ8fLe/+INZEiUo44Ug7
tLrmhaYOLsyWVgP4iIzPaJnA+rFq4uWamSx6v1f8cePfYpl55JnORHG2jRv/Ol6w
nBGyW1kFtyZbSmiT8xggLxC4paLMcZMZGPc8c0dyYWj9RlVntMZxMX4J52mcPFtg
sf94SrFvcQEtWSo+QfiMjhhEuTT2OxH3Ay8HOQDrDtHvMfYraNOgexRG4VuUgMYl
us35xlLHh+MyloDe2yvcsOa6DogCGIH5xF/OLilZAYtS4c0NVDZQTDx5Rs65+dVZ
0FA5Jc4Rxv7VlOLQSTH1wTHbzZAW0o7VYeM+e5NjusIfxw9xjChI5UyZaWD0fjNw
XX1/5rzqGHy9rhvfRprb8bDUPXzdsNjk8p1DLizR5m7U7VMurrvlrG8rAbbRMAZK
FqATBIeZI5PJD0pAns3e2lWsLf+1gKJausUPhksXxcdfNwWwr9tHHVH+WYE2Ev5p
wOx8aYwsPqYpuf7heOtLeA==
`protect END_PROTECTED
