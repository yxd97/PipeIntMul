`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vENrHYN/1cj8KEISf4WT0QFw3hjy0GpPNLAJuD1VXtgx7kdHakKb4TMWlK1ISq8H
r05Z3ue5qweEbJugi5YQ+sFDp9xinOIyIred+XJaKPKBkDsbyJrfGTP/8YN9Ds+s
32nJ9IpomYBbNYJRa4IgKG+HF4zK9It8Gwyekw7B1pGgeWRLwIad/qYLAjTQVXvo
d/yU2eFkKCff4+6bJScllofKj5cFDyY+6tffImNcz/MGCg7CI+wu5cS3exmAdgoO
zOkjEwsPeKFIJ0Sxfu1zwtx3YFZviDwGWANJAAkZEVbgkMMv2TntYWTBPn4kCnHG
vIBup7xPC2MspuPCPxQs341OyhsOd0a3EnjzAjcWS+Q4fSWB9tsfhTFk47t9aYiO
5kLl0gOEr5hKi5eH4qEzERhV9hde0nTeg0lBcBM1xJazZ7kCHPWX9UcQoSjVz2BD
FY+qs1Eq4x7qyauOZGVaSQ==
`protect END_PROTECTED
