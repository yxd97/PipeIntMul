`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N7FNKtqRmMLsnUmXwtAMJpro3cqrtazMX9W5VCt1t3QE06AlWh8G6Phx7m2E6UC8
OxBTZtdMYTjVy3hqmC8IXLStqQydu8nYAimMJzK/qyyF+CibqtnvG9MS9D3OyqZz
g9jQRdiXAjrsgYsU8XJYxZidTqAvX1x1/J8/QYV0HYLFZZaAwrfJjC0Zi3KADHdk
u6n1b1IDEUf5Bhp0cN4Km0XGPkygsT5IxtsW74kSGZFh/0C0wnOB9aKjskmoBuxz
iWj1Xaa/sae64kzy8c4mL01SYsFjrvvcbjteZVQ3BI8=
`protect END_PROTECTED
