`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXdPA5zeWtZyrD1J4u5wcKlikY2zyfChQJnbiXzJOCObEr9wFDRQi1NneWgQtRp3
HRMNWfwvqt0P/1Lb7BTA75UL+uz+FkezZIUaBTyEiFHSYyH9mrsD6GQ9zzCzQlzS
/0s5ED91UPi0A41hRQHQgAN6QsbEjBrhONxr86PTPBNSkoStjvLK6JEmpRlwHaA9
CIyaGI6d+cB+Vl32iaJ5oEr9uNN6r775UMrianLozg85xSUH7hJN9BwKAPIXXTgA
BTjfmRUnmelDDICrL4IQd0XCj7/gkn9Pbm6FSAw13WhWga1Nv4Dhkiuxqst5FsxF
P6X5cNEB/3Iayfc0I2VS74m5WmuwdFV4IdZxXc+ytBeFS4F3VLcveCrgiO8FUD+w
`protect END_PROTECTED
