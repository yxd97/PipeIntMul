`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3kwQ9Utx62vibMLAUpVpGV2rubydGd52DcfLgUBjp496WYBFiYRGmCsq2BCh3zB
aPP8HRlz3gRcHQhHX084Vzk3b8MAE0sbQFMXr1CDgmNM45lAR5HexKxJqNs+gJH7
SRVzoDgl/fOKFxZ8CjE2jy8S+nzZwbDiEZ2QIRgDfGaGUC9Ru8gC+Jr7LlObeWvi
nS52js7b9wDCdh/4ywOAcGDygP7uDINd/HS7MZk9CziBv/xbTG5nCwlDUTAFLb/D
AuIb/I1KsyqBUoL5UogodmukVAdOHrzvHUjmKL0B4n4QWd61qzfY7Y2kR/UmNkme
EuCSQZwO5091XFVL1wAiq3oeTQsOhi8Zm12w+IemvD12BpkFQrUGL4Jvhebzww8M
XyiRrjyjp7T1AmJgFaee8mr1O5VU//8hxQsz/Oqorc0PYWtALIzbR1GLGORWK0Lt
4DbPdW4ww89qbid87Z/M7uxVF+xnsVRm0tJ5yGvX/gY4yUl9MmmdbbguLeMte4YR
tkSILtfyKtR3cWF0VGuVfBKVZSaoi2Nd8qL6KvCcFa9oDsjk7xOoJlxtCMcJNT/B
WJLyejRcNqDcAYHbGP3G09skEtioTuGOazohf50qo8IAWuJfLaXrfEo/bxqAjJVD
4BQP4dOnhEKrzOplzpqB/eXoH2MJWKVC31iP56cu/ta93cYbK2JQI5X2ORTQ5a5Z
LR4AAdKD35RFi9Icw643tA==
`protect END_PROTECTED
