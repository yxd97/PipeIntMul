`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQBP9JbxkfSmuIP8p8fsf/t7pJFexXKU1XtiLuGIvUUG5I7kCjwbPN90V5iwkjdE
EfMhRu1OFqTrPRW6HQvmy9vTYzvn2/UF6L+G4WjJDy2JHcAksBQ7C98qW+TQoafX
hd4WivPLSPhz+mkZ7RvMe5KMkXPFYIj3LCRlWjolyyxaBSPX08YHwbVwV9zO/gxz
PQoTJsRYUWSFwmaID00xC3swf6yWdSKkNs8AGmKyYdJQwGlh1Xvld3l8wWDVlmvl
6NBI7EZh3hsLRPnqIoZvLqQgpCxPHNUajrXgDz1+7gWU7jyt8hKshj/6XVImO7CC
btjqx9zHmUw/FJusjG/mvx8rGDDVOlbOrKYhrYGoxBrQv2WTArlUtDO5r1soMtUN
Rpon4OHbN6zfZ9D0iC42XTNO+DQWxrra9pr44FcDg7HL9vlrBpcg7Tx4BZpz4vcW
9gCKsbe7AhOcuSbJtI2emKhdF4eBGrW0D8mrADnnBlagR8CDBm7+VxsunSTncMv6
tFCkIX85BcmwR6PhvXJomXoG8LnpH+Ad1xx0fj1Y7e7Nkb65D36Bcs7eVYEoqxep
Oyg6KYGjFV38XHOOH157zfy256+vLc9j5wEwTime43ucKIo5YtuF51FGwvPQV9ZH
teGyVmFkUKh/nqMqYCu2UQFQJ/8KBJTpeqBUfZluA9sN97YeE4CHhql9F3y868JF
CZ+kYHxKI+nxxdUyEeVdoA==
`protect END_PROTECTED
