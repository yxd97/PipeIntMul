`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uE1JH2dKC6l8Y8zXVWtTgJxkC7W5yEPJxnO/gcOjoexBIwfG9yGa/JVa9a8HOjn1
b4GJvbZNnzzUskoa2RfSqziy7qtw2XLrWaAf2EWIyFg79wBfeLjqbTXJdFkjh5Jy
rtp3S8YpTyrNGohy9i8tOZ4WkPejiODvPZ7vWYHUemLJBLolSj16jbGioVgNAuzx
59nojsdAnmHgVO5KNixeStjGnzPDgUQDb1F4bDTdyczNQG0EcHJj/H0B6OHdP3TC
+Sjxsv9Nyw70OEna2yGCOwXM8pUYX0dc4jeZChYM8rkMbrJ3cezjZveSydCHLWFR
Np3jwhoBlMO/ARvUgsfJt+faWYvpZVtlqiMdaZFCKFKGvqCg38SsmNg1j0czRtiD
fDZijpOeflfpKL1jMrV0vCAf0teW/NOyJMOAeRrPw3N+OSC9QaOzLAvzlX3pvFNe
vvfMAUAgN4Lp3dsVLX5qv7XsskYiOfNxWq4SOKX3sJFIR5kZrA93CdhCZjXz5jRt
`protect END_PROTECTED
