`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hV10kqphISTKVTomBNuDzDthh5/pzzCw6T8FvcwoYA2z0LKhhBzzjH8b2Bzsq+yU
xQlwVm14cLNr/vc31QvXfwSeuoy/JAZ3dg1qKgnqCmBc+jyjLGC6eKLtfVtMXKFI
wcR1sYMpESdm7dsJC2zV1yaNiOlm0uACEBfZM/2pAghm6Zph16Ch3ib5Lc1UuGfK
s0LWFu2FMLBmshZmILXQ5vKbjozO4/0e1OsnGc/B4omsOGV/XXAwOORqwLoTd0J6
AU76n45BQNrmLU6pmK++MYQqL55YQI87k0+0N1Eybwzio0u3SIA9O9MR/MYPJtiZ
U8OMRsgU/QqKJyfJs/mFwk+9Slv1MNDoDYYJiDbSOK1g/hRtIIxwglpEGN1d0kzq
Tnvu9n3YocipGPLPb2Y/G0B/a1RTrheozocyFWdJTdbo3IbPBA8I1+q+sBRZdLCI
Q1nrrCtsWx7dALkkSeEm8UJUa8zumI3nVU690yyucOQ=
`protect END_PROTECTED
