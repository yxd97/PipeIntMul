`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vCxC2PorzQgDJ1N12P8pisOqllVw8ymbl0VcYV/Q7zJxOKEDSp1PcHWJL8p6jEQP
bCVRjgW+nljeXzjxmMtfvQdXm+npuZGhfiO6wxSL6dJ61DprpGDqCrsOlFPp6yzj
UwHejLgUlR3q8fjBZNTfWgqqW9lhsse7gDr1u/pokVeaWcrR8V+CRqnQ51Hw/5D9
T7sCr8atxGGJxXbsvb9z92o8zMVSFkXrV5gJowP092sMvlLDrF/KeZaOiFoEUnK9
ZfpFv/bKbivgOs6MRBuXZ6P7LXvgIyHLaiYcS1wf1dkolcrVvo/hFqiF1ABI/qcN
HB1yZmwCHj2sQnQTGXLPcKmRJNwBTsDXNQED7PnSP322l+mhat1XgOMYTHJuIOol
jh5Bf3JrF5LIUhVFt20vp9kUIrvAreG3/8UGfocdwhqpO8aEgYzXse55PrWmFBq/
ZQb/z6quyjFboN3l8IM6mnQDibsZGY/KD2tiVq2SRSWmr1CpP3L6FGIjl/7tAgNY
La3byG4GXOA1OuPkTID0MbrjkYguwRif2gYQN5qPCzxXvNT0wePaarMjINl4/Ll7
Z/2USm5VV8Bk7WBe3bC42owzaCie1RVxDlUGY/i1dA02hRNztWLeBCh5gFRaz0Rn
ysRdz/ee0mds66OP3jqGaA==
`protect END_PROTECTED
