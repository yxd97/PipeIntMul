`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Om2Uq0/+Dg3CvI1UFWtzJ76XsuET8x8o5bktXydaKsll/I9sRSJCcUATe3K7B+FB
jnN3iBcvKMBveq6FcaVDRMrIbE3whp15cxO+fiCYUyuLjyXqBfWA5jle1fKiZUMt
ksewG0QOlUW2wdgnIRWt8Z1oMIfTwZ5yIlqXuixOxhINO46FBx/5eBFkmImUgl13
OLtsy1tWHPizvtMEkc4eeFaJ5uwMoRyjPTawOF5OQE0ku0igMZ8FKlYtfzIyln2J
hvHPfRoJNmL6v2va+U5eDst8IqBtQHWcrrEXIQ8O9pIjCvOZ4ApCMnPKWh+/sLjK
C4JoqqWy2OoVR2Uy9XckMqdiYDBpSfr0r8oOzpFQPXLYwidvsusWFlG64I5zDp1r
`protect END_PROTECTED
