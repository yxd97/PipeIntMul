`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3ur9QE/ZcExATttCrEZzivUjVHvUfgBXBhICYfR6af1TAjauHESNO6kHjFP4AMZ
VZL5+I6FmqKeV1dij513SesLGd3qKp3Xz8NnBsSnxt1IEx9GDn36qzdGXDYRDxrg
lfIMg6OAKu8N6dkYeoGorN08Glgp5e55Mg3uHxC0Up1umJG/bLb7W4oPEna9H6hH
3hvKTyQetkBiFZkvM8S+WLzGCwMjbPffzC/sAKCg9TDrqHRLoXwDlPKetc9qnShP
h1w1xD769Pdc5auG3V6qpR73WwFryDZ0atbe9C3EMQa9x5N4AwnkoJPjYDLdg+Lr
E4mtHUBQD6EdtbR/DJ7JY+BwtX0PWvIDqvGuLfi/H+Y9aemukDTApOekYg0HRpnB
FebvI61013TlFYaN9l501Il9Eg/M3r0RzsVinqrNLwUDGF/qO6mds4d4iimZId4m
CVDD1p66RZM7Qd6wIFSYSOc4yhQ/qcequ13IDvHIijGF3dCEkAqJYDo4HwqQV1Ga
IgtXaflnvgZub4pt1tkzomgA1z2DoMEjVD5k2B8BWX+dqtN9o8cVpWtRlYrVhvtm
+JsrDpVCt6t1lgzveoZWAKEB4TJvDI9MbAJ7Pie5wJURxCotPmsNFyYBHchWXfQb
FqiwhbxnrmlrmRqoBI7Q2HLnnVIHqtdS3YKLRi8y/UB9LvVIRTcvXkdogJ4toUWB
gGCUDPd9+7IwXWY+DXDED2Jxn7DTEqQgHiyWNZpbG0HEBIUtAzhAfMVNWdW1FhXe
kHxTnFInoYQyGYdw3tUSMldKTq7IKegi62F3Q7+6n+EU3516D24fqcdlKU55Pe8/
QhV14cYE2vDYsndc22xVJkvEoJHaDX34t/jfNuo2KI8TQQqf2AH535mST2oXPVnv
HQuUYnhOSZ/sqiWOqKreV9xVMTryNVR/oaChdP4CoK/FMLy95dvdQs0LpsZU+FJy
JF8u3DSo6z9TgkLh+cm/gWgy6bs+tr2QCu3eemKyuEKXzK9fNo+G5oqQm/o1o4vy
eLhDN9Z+Z9SqJgdk5sAKORjKmuKh203x9mOIJytPQKurDIG2T0sVJMv9bN9iZp4o
PBX8eR/hrMTnCBVltzMZOatA3z8U4MZRaSpottR17BeKUwMWoZvpyzXTNsoN5zfd
75JGkXZvbYIr0AbTnAN/bg3noW3nv6uTGqnu0qZ6Rj3cAjHMZAoO5CnFY1CIKeoQ
r7fcbXfIiWKb0snX9v7RQsoPeNw33HpS6agObKMOTvKDBlNA6hZJ7nbJDpbq//3d
94p51uElRqycffj2t+yoN8t03kKoRKMT174v+8y2OquhajET2ibIx0UfRM0dn5Px
nXXqGscqNTbgK/XQp26Pn8edJlE3ioOpR/eJBoNxjy3OLtwb4po1KAKqzVZ+uJ5Q
AP7VZHrR0xRbywd2OuUNIyt+XUH/z/Nq8ucVU7CHD3YbukO4Km4tSYS+4sxfV0HG
dru+T09nu7gZHHtqXVZgtD74F9/UrqoRZbszWCRyJP8Pk9AEcGFPBU9aO1apkK3D
Xl0QfiqNDaeZNEfu1DVG5mo/a/flpel7qtIvD5/RBAsJnIBXvGbz7WcHoO+XkUj7
RZbS3GEw8TAb4cJypktVoWVLqP0Pv6WJ2vPf4Yc6rU0d50lICzaWptlE7e+SjpEe
TrQfGAh94oZ2N5WcgFtDt4BoXJ5mL8Ht3ysomWVvuGVCS64nybk0A5TAXZ8+SHaO
u/AxqnCHOyELb/+t3y4D9/IrukD+sqgcY/gE2ZjPgSGSB9kjLQkvyLrfH6HWQuOe
Kp3nM/juGFXj0DJSin34LjxFNm9o8qPHmKMDptLnvgJQFys2LlaLX7DIt1prbcyZ
oZFcqDr0wxAdbNdD3ZUYMJm72KsgCHiiIMVr6rfZaiD4yN9qfwqiXd1EhM6lvlhk
VBvjd/tTEfTIAtbRT2WDyd/WiU3DhVAhrqzyHoFl17KecqKr98bj74EKZfN2F8i0
kBjjRB7iHMD+gJljkSIe8y3/MOMOj/sxLffk50+NT/eyS2H5f2lNgozQqG1YUN8V
Wy6st8F8T13ZEnsxl59g+xPupSExgCHIV8vd5h3Z5d5PNBR3uFWkRbU9TlsIWE38
uLqAodIwjiiaSL5vKwxeJwFhbJNdGtTO4J77Foghnyp7kksqBZrQWLQRq1PeBAdc
4rADz33fqTJ7rG+I+6YkqkUQxFPxTiGsXjjQoQNdqhT4BKehTesHFQ438JjwHOXc
5tPpNQcT7itwWA4A0AbOTdTwSsvBqSNIlT7jZELoYckGV2tL5zJinkBHESJE3InM
72tTVircGHl1iaXMz26tQdSnWY/Or0we9XES1qnkphBGbddVlh+CitMH0icbCSfO
rSiY2w7Rx6gFbsilgXrJfoYLWgseLYV2S93oVXhkfHifGBjndjXaG0Jerbiz019j
CwsF443xtu4K7VtFSjJYv7hKbzkp4bpw3TFYFJWfCevRGBDJ1+qzN0bcD/d8AbHx
zgkZX6TF5c5z/l6VhMW3gRtnCY8xyxEHwqEAjWbU7jRrffAsAHLDgm/0Nq2u5KdB
TUk417KL2PeOsHIkw9zsBwij3Cm/fWFKmkjBX0sv+oRc1Y7ZvKDC8Ea1AOm4/1CI
lGxcz1rxecGAz5itC2ls3058xV1cAk0vIAzcU4Ckzbag3nmUmlTqmgQx+PX5n1FQ
s7D4b/+mWFTQKw2+dna1s3d8qRySCnNdj6c/9yhlMsz/VCID8xMHjpJOhitHap3e
aH2NtCl8/K7HyfGOYyCginapVoIPwAcNPU0w+agDcf5bmb23E3Bv+o2YyN//IM/u
k8uIAHIwOmWUy8cW0Cd+xRYuw8hB6eXhn6nOkdkXWnjxu+c9fhRfJUdxh4Vysr6s
ujHrTdfFETxdeBefzSHlWypjw4CAH+PNahynUg1mPkLCstHQj8sw7Dtk1Qa9SV/J
cwccklwIHNJrWitPkmprGXMu4bQo9HDLN1Rlfc4yfrgprtrRnUggH7Lzw83TI+Zl
GScTMRgdUHt1tYRlWipbrMCO8RD7hcLy+W7edEmTfDcBTwkEUHOW1re+hLwI6IJg
X6OLV3HB7F8/CAG1rciSRQJy1Z7aFtimvilO7RiK1czmbqT2NlMVzaKg933lmYZJ
VK8k3rK1EVPhp1SG8orEfN9JvCNE4D/d5HnXJuLFF8LTxCWvVSE1wjkAptT3thps
DMWfQCWHxlMHfYyUURaQCFcqfloiX4PkuV1u5gdJxv1tpJ+MCey5M7jEf2BSJOe9
chptEsPSPHacAvUDT2t4SIyFzE1zKMdqatLwwYxbwpSxB6CM98dhbt986wZfdUHS
jIqtAcx3De5uPWQLoo2JbQDjddQFR+orjZDf8J3llQe85EjJ7rN0w5u301P/vPuV
2q4Xe/icMHTpSLv68ufrC2PWcgRehA1jha+Qa+zAbcG9ZIcc2ba8ZLBDRASoxB45
rV+kngMcWLFqnH4VEJm57ScltdlodklWet1v89zMshh0iMwczUa2Hadi0ArmLNlJ
2YnSRkH1+LXEcTg+luy6whPSx3tbvr3jJGigOxlx7M+fLf+Dbx54KfsoD3VeNqXN
RyXRiHv6lv+fUwbs1gcg0lMbOEggUxBNabi1jxzFywW1mG8yZu9ItbwwIlfYWT+/
SYfkGij6TGYH636IAGQWRUxBURHo1yFxva9P6TFFg6U9ilprlaUnpFHmqICn9/Jf
czzB60MuXYu9Sb6Ma3RxyNS08wmQ+LqG4hSI22jF0nAOh7NTT1nyy4HQXzdwzKnT
3B3HtvSD+kuwa5opu/EtAVSElxTCghR+fxa3bdZOOAot/ZhS31XxtBHAPXrBcen2
rFR8UHhlMN+3Kv66Iw+HbvjgVhcXXQXrVXZLsi7FeGOjhlPzm13wDPP80NAm+LWh
p1Grs1p09tQ4ovGtG5mh2OgfjLQZKpQplf7CEBwOBkoRdZsktUnpunnSDYkWemzH
iW2QSkrQv01BxoA5RmcOaGOwNy2hqFsHxIR6VJL2+T8QD65/XCf/yg841N+EIQuY
VUmJaKTNlQ4qfOgTaHLz5b2j2hbIVseyWN9VCR3GazP2lZGUFv7EH4j2luTF6lV2
bgU081WDrPYojed+JwEPPBxyW1c7sszfl/9w0l0HT4ORzT0Qfvfqo4VjlJ9WSpPl
azNSvJCzczHQw+ZlRlDpOZ+RFF8br/PAIz/0JFpRgX5pNtEnVKVqKIKOATPucoOH
3jMVpOdBHRjTrkZY0WYZLvT0yXis3VUxk/deyvUSjhPhAVsnT18Xot7wgWqPa8Li
w8kjLRBR9RfmGP1wPOwNUHWccAKCEqHsGkxKbm4ocwknX0kHDq16in7X9+LQ0OoM
IjJIZSW7kJlYQslURztVfHoxuBgdR4hI3DthyMU6zBDRT2BijIFtVvZJ0Xv570LP
HB2SUwzaaw/fFK828ic9wS7pjJYv+iIyHCxRdeS5vVkUs56E5NQvctpGiQtYI63G
tUT7oSgIJtvzvmRbmiurh0jaJnZ0EhK0zocCeNS7PqtmsyfQl9EYUeTzWjV0+om3
NnQp6KL/Ab5R0/b5lmeZZQhtmqOQiQsfK/YXTeYNW8GUnQI5BGTCnZKePozG5PlH
utowz5SzE1USWmC0mARNS2eCzTQg7fcIAAm5CwcDsLLu1kZ9FI2XuhVnjf1qiGEt
O+dKnIS73F23IPTg5A0E2S31EU5oDKDECnayP42sLtmW6DzaVGK5UAAD5G9NInQp
lP6qWhiqMGCqPX8XVX1rxd537+FWI4fMrF+sRyV/rQlpPplL7IrbERJwpsrMxAsl
pCRm7Kl+rVf1+tvTbhCB6IVNhq8NWbWP3PhwuszxDuExDUVu89A44Ipy9b4uvRqp
ocT3uOmpsOaPpKR3zVTph9tUbm9RhaoPveBzFfQikwjF8IGM6CqEPcyPTQaZApZF
oNcdjOw0xqY/+/ZX+WAUZiKcBYdJcE4XkTUAfpf6x4T5QXgA+R0mGEBwqs5g6MTU
ha8mm/U2CCIaQgFyOLya6YnpLZd/Bl813y127Y2zemrR72fkTKpwq9coIzCKcMSK
AC8p0q5Fd0B3rXtwKxlSoBiVBGXFYl67/XKcY/KS9UlS4TJ33lbWvYO8nodnTKG9
8+0e2Hbfp6zGxg9xbfrb8yFrQAixk3YpidX/OpSjfUY2ew1+5uo4B2BLfx3BZ3SB
Ok7XiPrrM6hZBSVihtj97E1A23Nxi3e2AacZA3hEK1scA61cwJcXRDI5cw3QRVCl
2srB3Y+dlyEUH+qe6H+r0QGadBSP8m45gwOSrHPnMVcY3Xy8erAkIl9VJ1suPEnc
4vGd4/07opR+6XocvByv7ifAZocRH4jNyd/2N00Mn3m80iCq5EjIqOdm4iwUzAQx
c+v0vBpiHhJ12KAKezzZFlrzakWGhC+oYkm2UOxohGfjH3vLBG0AoTO1tTBnKyU5
TL7C5mrvR0AHxrmFGo8UlZxRTDT1WPY03L/8fO4e5nLxkxcoBMyrZlIX1B0W5vMq
to8w+WH2zg6rr/LHgC5RoO1IiFNS2IoYGde6Dyb4ZVCtUHJmbU5JPnxr5XpmL9QD
LH0Y9oufGkj3v4ja8DOilvO8a9KenteISHBjmSEzUc6EB4+vZpv4nzMYQTWUPnl/
m3561Pwd6e5aWpizepG6PLGHkLeaoiNjb0EBwfUMviaOdhvPBux6m8oJYwxLUUOH
1ERXRpKcqd4nn6eyBUv1r5qAfS74r7gVzdkEEqCgEK2HnoLYL6i6cNcC4HAI3Ra5
YaO2dIdQkfct73XVnNYJGCOC+wkn8GmWXMZdiBFMnnyRFysEAISmKRpNvIUYZCqf
OEd8V7ruSk5/S5ekbG3qrRKy0QyKNrEH8fwjdXlZv+lbdEccItEItA3Maxkjm2tk
/aAfXP4ocmizqxj1ELs973h6en7t43XafIOwaIJiipLk20Bi8sf+KJYWXdPVdk3y
ByCG1U4/Z2c3Nu3PvvBdk+tqt3hMkzgdN2Ajd2ImVa8WAOcmVzG/4S8/gBjOyZdm
LGcvEAXLlEMpGeQuCq+hzEMKqP/xJe957xfJRZ5Y6Aaqap5QHMl3l0wbfc6U2E/5
NNneH+OveLa4fIevGyOclzn/iwgjan2joL3TvXrBzfWFqqGObyaV+vzwF9erP3fv
K+dVWNdosC3TSfcwzMTpLEu2PizZkw8/sHVAk4MeeVF3wheKdRamWR/ZA1Rfw/7W
hLZLzmyc0QERrb9OvBu4WAe+DL2RHsKe0sLPsHRBejk7DQkTtHzSF7l6LqhUj0jX
SnBtSj7wP+TI5zHm09+e/65BHw8YclqMwQrxFEkKJ55Suv6YXsH89SxmdMmD4499
qyZcxPXcs1pieo66iK301R4xTAZ/7vjYl2OvUSoTF6MkHrkWf23sRJN7A5CA16yW
f55pGf/V2/eYXIG8ThOXVofCUz5n9u8iiS1JbG2/ePrmTrb8Q/rlR0YxX2PyUAjn
MHwL/XfYlZiJ7IBePhnNH4MWwFaDwNBmMMRG7kLBzSPNGCww7zm7FjSmiXbuKn2a
XuLr0DWy//KHhUMR1KItWg76cW4sLo8UzuYTMOqQYbptla58cewmceKjr7/O6Lmq
0mHjT5um6dS7FcMkjNg515nDzaA2SQ2AviTYbdVy/ci6LigKtNulul05LfqB+ymw
OPo8J6bPh4Ey5wZ8wVMwyb+R0fVSAz4nMNoltDg9sVcftF2aQyUym5azAsmXEUpB
MnA6Km9vzQCqXJSY5Cj60fuIxWIxjds1lWjHX7ctKQ0Ioy5Lj+R596HmVgtpLO+A
WmBqCKtFO8MgCSMiNc+OMbEun4+TIhCkMTnzwyZxdcKP/Pk2TsyRZdUamxFhxl5X
0DNgS3gbZjBeNd8U24duyKzUxmVwsRaPqik6ACUYWL4sE8gKEu7pZG2ClUKMui0/
pSl3V7IImQ5Mk/NenUEVQ8/CuNDmLA6OyYzsC1SlWZpKUr85MCRHJaP65qZbE64y
r0BRN2HhUKCiAQ/+U+fm7mq5T3nRmBisHCTqETFHzw10M14QehMGHGUL37JaglrA
SLfXmaTFbBQhX6h3POkyJ/EzrlS5CaSC+xeJkEgqf4LprVi24DkMqWZ9YWgH1uRo
yUdPkmbVun3CRktwLUtBfhLlCmzwgzJYUH3thOEmNbfIoyo/vpXlDNocOM2I4ZkQ
vooN8D/4/nmZOOAL5pnehH4ak+dEI0O9QyE1pDd5OeHWhuJFthSGnFeug33vzpSV
HBdSf7BrHXwxl/Wh14q18khoUDRUOx1ZHGbz+45bebjIkIHkFNMp2s97DrxCHAGP
k0CwV+3uTfqHvR8YRo6ftvIf7IG9zhM0q96qEu6Jr/xsb3j+fMkT/KDDXU6+JcxY
ScmBpFSyL9VjTw39P48RMGgxr8ByHcYEe6VPVRA42use1m0SfG5a2WNJYH7qdLO2
7oDhWKpGh9DHsv4qG+Ip0zAFmARl9RI6EIn8QlFy2YWbYddut0XNI1nKOXbPWufC
/12xRALNBDMrB4/9WKZHJ4rotZlxdyVh39ZVXv0VkafWQ9RLMkroLDuj8p3/80uB
PF+qIeFym3Fx4a+vRjAYpAVr1kvgey+KaPULhbJn6xlRVdA/K2zGA+o6zmB+y7Tk
OyAEeZBj5X6ndPxgdB3MoVT0+dSz2de13p3Gj8CgIZQXBoGGvBU8uw6+MFEm5lcX
X7yVuGjUYmqLt37q2g1iUhn7k5LXN3Vv1nyCGRmPLi+i8NZ8tv47I0yUYFjVG5Eo
YNhrJB1a3fEPwIN+0KA7qhswz8WfQCLVd3tju7U08w+5zG01bhTMsBtyXdM85Fr3
2iYhF45/4QMKFViI0F58J9tDcyqZNPBL22LnIfosnyw9ypcP31mDx57UobteUpm4
8/KiANxyKM1LJp/Jh8nf9OZ3dtW/Ut/jrwh0ly6ywESfLdJjr2gZcpS2zq+LSneP
0LD2zHrOLjnV0nXgbd1F+qmaXRxVfSKplGSfosEmjiCY56kOMiciA/wgQyWjBG/S
+/CxarbPkF6WXqboqYEt7WF1VYBNqGElVClbfZj7RAA5GcKLER6iFsk+gm7p2hDk
OApwS/sm9dNpfaa6SiArJuWUqJ+clLaGedbw48o828KOK/rpbkErNC3dYpMgK4Ns
8Ggzf7L3QNWlwXqvNMfWoWRXwkVzgzPegj3C7DKvlRldDy/stu18/icy9ZHbLfeQ
fD5J554c4Z9q8kboRjqBBIIMSxc+Y/Ihnsfn40/bo5Kltf/BNJzAhl4ks1+sPsy3
wBoFalAr/adRZ0rLQHgQcKxNl/trsTSyhyHjMpOOZKb0Qi7111sbT6M2yr4sBHLh
qVch6/cM09ZgFMOlaRPEoc00y/oEwmtQtuej1jJFn5qY80OjJvvSjRe0+fJBg1H9
bWYufwFkYX3FNPT8hI6gGmSOYjxF1h7iUSJ/dT+kwCq+NEcAbQaehmfXMdTncE2d
/MYaapV6GqDYde7WehladP5I98aPFfmCekhkpmNJVKALs+75IlaQoTHF9mrULLgO
S/XPwSnl5LBDE8Eo38WNtSlRBm/lvYPSIjxxcA6H14UpvV0q3Jm5S7p2jRvnJEuJ
tXQT6xlQ/nqrvN+t0+0NhYBxptK8pKKWiv8iSxWNpTWed7waAqFmNE+XctKZ8kNM
MIGi7D/27wbyJhf7M2+2JH7JMPbHVio+De8tPWHIA6Y7mEoo0EWUlzGxALcLkjtB
UzfNFaUQM/8GtactKBDQdlU6OQy3GrG2XwgtHmZbno38pGO7OHsI6i5v/LKivYXe
Sv17ZsFvAHnRmNTH8HMetuHvy6sLg6+bdmiaXgRseREd2h/mvcu40rdaaY7XJOI2
DAt8DtKdL8GbP5O2EwK1S9nS7af3M5sCNf/kIwQ1JWonIpmCeCm99IxA7agjZppF
xn8pwOxvQM4hqLPHOr2k0jA0qXKCdAEZNOiWuF4APXO1v57CMe58t6oeoz/w04YD
D8iqv1CgDRL8YI5tF3oqEMTeOM/4hocQr4rhlOt06DrTEtoOOtlw/AIQoMrq02p+
2Z8V+7izEJz0u5O4F4RQmPTLbl/BEr/RK6uplNC1wwSCAKkw/i16xeT3Jg0PyNNk
G6PRyKD4E7s8jH6h9ApBtUAyy5i0Wh+Klt9R35AFn65whwGKXqrwN8Lo81txA//R
DJRZvmX1bv3L280tgbx+JScKQxSKwD0o3KvtZ5IyxCPmU39sbfJlFX/hEy0FAhO/
NCxoZyIq9/qTtzcXMuDoMQmx/xyP9oZ/DGuDyfX3EOOCDTn8MDBjwman2m/fduAG
9bi2qYEA2H6w7vF2mNsZt2yWc02o2NYot4Ew3Nl2K33YJsaN6ObDDwX0r2jrcuq2
5lUbDlv/UTLweoM20NiwMhqrxX/q0fI/FxM+q+MlDPhNw2/rZNuLOod2oTtIBWsd
JjEdxoAf31575JtisGdSSV9nIeYtpENzoSM+2adxEZv/MyQ6Wmml3RNmz4W1ScW3
3gj5ndD5TJlU8MpCV1w6+VM4NZQjHxlaazTtVOSU2FKRCzx1byMZpiEqJEMUlWZz
mw+Ok1xvP39zgBXSa+5pWTmOiFPqofiZCt8ai/9Fv2M+eyDzz18+3LR8CChAtzuW
/cmnbxYwQrpWRBPlIZM7q7xQuCoa2aYHIMCHp/D+/h/Rfi1ajMNlTOZiiHZ2o95r
5mdisOQY2e8vjA0l79eEDq3BZc9I0EzbA18h56IvR2w+kVgiLhSdGgBjjw7GxP8Z
fjfyc0ql5a5KYm5VmnrwDzyw3+5f7W8/FJAzT265cYlheT+/2ZqENan5rpFNqh07
Z8JqGvMRIEoCg/4UqH9oY12Yvpqa1xF45c6PadixQphkwavpW3ureVIukT+7ylqj
Yl2ruC3+sLHD0RqxBZoQd8lXCnKfqUxpVDgVWfuQw8KjnJ4MDgltu33pivHGU/gm
CVOoBKGnhRap3hpkNv66IMfBiMmeVePnEid2uMov/e6K3ljgmNfEIuLd4wPP0eaQ
8AM/WBGlWdkQK2iiJ3EEtGoxIe3HFdQxWvmPZA5LzupcLuomPyZSGlXQ91SnFYvn
rqruH6ISC/oWUklvN73mQ+E/dQwpuOgbgFhF7HvR7eu0aOxc/nEVjtUaBXOKX2z/
LgxFxiIcyAbDFLkK5U2k+owMKedHYLpVjbzggY33sQeJqetO6lWiDI/s1IT2Pqz3
xbxUrasEA+fLTwdFpK40maFVhEdm/CVcf/QoltnRxNcKOvmu1D5vXEGE0p3O2jr3
f62+jUOr/zox1S2N3eKbsZ/58IPdFhLxtr+2eKnRX0P6eXJBJr/R+TaSJQDWSfNY
ztFzhGoSLoKqylpHzdOGRyNsJ+bB8tXES1G9sk+kVfDoJxwUPx729q1Q8aS771LA
t8mIWw7trT6x151qJzPVt13wJYMXyyuqH1JBG7ZJPNuGvjGA/H7UtUuGT2ZKIGAo
sy0VdRNJ62pVmTaOfj5y7qlBj2UvpameMePzfT820uciDDm37aRttoSavfZFBkxu
4bK/0WDeYH8Ns6AQfinEnnBxMXbCdnQTfQffoRPqPSPC0pi7dNAf2VF1C+aUMB50
sWzK1W/xkaHwdqcBCdI9aNmnQ171QFveUSHpflaShQFPHGQlNPNsx/q4KDdnAnGV
hMG/zYwxdTdoH5FdAUPrIQbUB1brEXEmrKJJdNCYrILfvY6hp0aW6zHu8tYdkKGY
GCncUxsCaCFhCGbPqK4DF5tf4kNW9WXtObgyuh3BoomUvfpKwHTdxG3BR9berYBh
xYBdosyJKA7rfNYm3xZvLx9KUPQMZPpAsEu75+kvSSukpz1cVXGVrfwVTm3f1UB+
NuaRzvJXwVtHbZzRhu9/N2pL9AoKC4E9TJhmqT3EPdQpq3XYiqD8J/H6K36mOMg/
oWNfkyFUzZZMOmYn77VJfTXFvmBfUChGnqQmPnrLiZv0r9mrteBAq9gYz0Sfdewj
9zQ4CMxYPOpjoHnUo+4qYn4gpT+XDrxwU3qw0iDQSorzmre5/2bzSnAey1NBVntb
yNXDb2nw1I8y/41MoBE/xSMEnSjDXKM3smjC23nmIn03sRHJl3DJ0+R/pHLpNPpv
K/oz0JlBraNlg5WurVMKIucWfuKmWuph7vYi4R5zGV5fcIy65f2VisBZgvRySuQx
wyeDSW9uep/Kn1Ig2KXeP9+c9s1J3tDaLmbZKK0WgPqDE0bIsYMAJaxPn4t9PRkv
PlrUSVPH19Lqknlvtv2uNbpNgHfirVm8bfo++nCEfkngSIYy4yZyI0rgTGMCMfXB
L7GyWdUaoU68hyoXFAkVApopRQ8wxveeaeElI65RPwpgFc4pRkomgFDM4WWfcPy8
epvoiLB1WYq/8wyOatwnGZu2OQlEyiwFqriMNhHnwLDty4pXkk+NDmaG8G2XngtE
zD+WSZzU1gDtGwDy7e9qZGOEDGd+EpX6W2C7KIC0QBSio/HTs198hGjHsgQfPd8R
lphpQWFw6HiikOCc6QAZhG3lz7C5ONzQaSmniFSb51YNhmdFZ31aVnAJ8AX3nOOF
kOcv3nlnubx9uGUADO8yeHKYcYvFiqVI5Q9F6OWpn+bjlLN2n3+KAlSWx6Q6mv7j
/Btp9qaZ1aUPGcbMalC1LVGz23XtMu0LM+W7t9T/cxdyWxirOeKrP7p7fskJ/gkH
ObCVDMHPp5pePSppm/uxET5RPldxQx2Xv8EQ+ENJeqYsV2xOaCmn82eP/NVTFRbk
c1wB6jEkFZubp5DiiSUHMQ01omra24ZtgAf0lsN2DlidJT/fhQBszy34N/U/jzwb
GZ6lho6QzKXOJe56+Yoasf4ZQg555bMCS2gLOUFVF7Qv+eTUi/SuJworJr8UWX7S
GBw3iG753p9+HaOQFM5Er566y13GlB4n71od1xQQtSWkYTSq74VqBPKZ86z4LwlR
StaOdQpiVeZEixEyTj54OeUyrZG/v3ZMtwrLSLsTdvCkvia2Mc3F4nOGj5vQuUxb
qWT0Y33uDeQS4zZabmop0qvJbYXTlIEGXBFAAKUJMNbsJS3wErWIzl7fLg9t3lhM
Gcros0fTrRYMfLDfl842GdopzNsQiSH5MH10oVJz5ex72pAvlZTKnCz+4zce7UCm
mJ21RxiwfOUwiwxzGxSdedZC9whHZdJxIccL2dV/wN9LQVd1B6tX9nyw6+U/LyNi
8f6mt4SG9ysIoqt3sb8KDbVZDtRyvTKM8Yzs3xJMATNdhYR5IRbXvMXi3i1E/OT2
81KUq7jf7pA//veojL4hNPhUxKpR5ROHH3g5nrO73dn3r79I60GDcXAvfOP7ZdCz
Axx8aNGW2Gg6+wB5FnipSm5m+bzOhkxNOR00V0+KIu0Td9VS23RQEj7tROD4v7Jb
CWBsgi60o5qHLH+wt78KpQFT9dyi5PN4E7KtjlHOX11mvPdDBR+Lvv16st7Be/6+
d2bjhR/xtoV7bpdecOfB/iELCoq57YZcpo39g16D/8LMr3N9+IHlBLMqpJmqDPNb
1ayXTwCx3/wLN1slLbUie6903nfwFA04M28Q3J5vNirkeDAcSQ8R4yo5picAHIHR
Uyna/dYeXSSvX7ksFr/u23HpHU1ulvWPYzJjR+WQtIHQRa+lPuYsdX9x75g/LSlM
uOZ2wuNcf/hY7F5+Gdh11N3oBy216hn4uvMHCbOPKeOBlrtdDNjm83p7FjRjmHFV
ReL+q5Bwy/9P3TcY//Ws/rObw+T8aN5ufjeUDD6jXwP4ZRsGTcPnbMqbEZRrAFsG
Ji/Kv5V9xIJ/H0i7tUJK43H5kDPbZcPnaL1LekPyoicNBbfoD1pIs2pJJhlpNn3b
7HYsiIC+TF5Z6D1+9LxeE0QKizjVY6H3ru3hyBsAjhsOwRwDYehVlJraE2F4E3G5
BzSsb1pB+HHMmHLVOVgemLNaruRmWl4RvQKMGeIUeRqs/eMJMAZvNZEmQvBKPRpg
APe0S1p8jjH8TGsD+J+uEe/2Wiej1i+ZWeIYPWwNS4KuN1Xq0FuP+IcUwYKM1n3k
Nh4JB+pxEpiXLSyw0DgVTld+FyVcEGFR2KWwZYZqvm/OUWpaNIXFFdv/356fSHGZ
TCzIY2h9n6kggj0JxaQbu2LQcfaFNDl7I34PPOftv6p5rC/x8g7qc8UMaLybfbQz
uc4EvuxkEQIAj5UC/KJvdOGQlA+DQe7UZ7vdVgkPG/pC4/aXo1xyDw8dHureFDns
LZplw8Of0zP4sJUFkGLUrBinHiDPz2mrGhySk4VZWEYRWBkAYzcL2GJo1we5j9LX
Mm9JqpgtYwYRwah7r/48EhZKU/m0QfEVRF0uxtFCXOxcamCM9j6//qdPAGrARp7T
qG7vIH/cPWIdMaW5y0tB0RAo7G89pEi2J5sbgPoIGAqU9KPpWtC3oG8bvmIIExHF
Fq/ABgGy+p6iONkeeLvLlCSdrWOZA13ip87eW9eoVOeFXaIHFc6kwKTH5cIADMYs
EnKXEqOxzV8FfCYa4GiSb03+unzvlZspKZkrEIr9KwZbfB5Fv9vj+5+Y56QWJYhi
nb0XUjv2H2JaJkV25S3h9RF3LzMuOeO7C0IflsyhT2oWbk3/omDnDWYmOJzR64Mw
tNDqwARKUvcAk5I9qexQeeAsvwxF+1O/U1AqhesYjoVXe9fk1lo2qzWzrDjKPWi+
8nfDD1OiZLw2Zp8xjqLVuVCQh+i5klYlWFcPeHKLn/Gy+dFCJAvgEfy/9hbQqjwy
4EARP5BRUYYOJ9kS4mw3jWnMsVEoY6usJTYDfY8ewjBMGbXgoegdQxGxEvbundHI
7u36A1n1Tqm0OhdT+2O3wMIQTHyy0UFQ+NTds4NkZrY8tbN4R8gZ3b55TT0F0op2
dGru/lPkbZd9fRYU7msp45U/qFSth3XJOO0oNg7YLFfbdhe1RyLzXgOqnNWGmkGY
MtQZgV9kSIpHr+/1ETbF5SkMkkSwSikwn8rQZQUD3I0VWkK0M8xUFUHOWOtLg90Q
sIZVGpkcww8FM3oZDP6/NXY9oBJWG3LeSU5ecOOLc5wQBG5GJIQrea5fIThGtdep
HZwF9a3B+uGNpOFJID1ziinz7HerG040ZUSKngsWzrhySkS2rxyxqMIXeboPnNbD
bXjlFKsjYPYa9MW97Twlu+JVljBZHb4Udc5M2jcoHjlwzAmVi79G1JpSM+AHQbGR
ZVB5+p+8roKXKsfJS85HkrdTvQvrOzG0lvgkq7GhP02lG7YwsSm2a0VIVCYwFui0
fVdwA+FgTiD5FuAG4zjwpzR5FXCDWdXD0xjZVRsYj5SfxAo9Js5oLb8uR+viMVW2
KPxSJjvBL1QPQd2/sfBIf2jtGZd3183tuLv/1Pw2PMPq3ZzQmofXQVJd12dHrXDQ
Uj7uRr0xPpd000JProL1OzZvPzE4LfTvJ+ONCKRKRPbntl6mecK8YVN4gZtI6oyx
C526hv7fCcmkm+xXREjJ77cPaT7kSg9mAZuGuSWUqtoW3kUPfQL852K3XIY3robK
3RZPH24V9XEmzlW2ORyc7SHEwCqDfApM6y3DNprrLUM8JuCRda50tkbwlH4jeumb
Fl33nT0SrLmrrScHAxHh4nQiH+/BXxZdQw8uEwqNdTNnDPJUqxSljiUeT0ddwh+Z
fD8LJ8gGCKzaHncLsKrT/IYWuaP7YQIqrQJkttfuLI6fJnYJYV0YnZql8fQLXev1
m0iqDQ2WHh00oTWn2cpd0JuBOuF0m+jcoYZIOtL8U1sspZU2sVSWpPBlzRGfEPjG
X4jpXt6dvAtPOBiNa7woQ4RP0Bi2o0yqTjrnRnqHfFY2VWP2Iq3stk04SryGnEgA
Id5TLEQYhk3SOSmxDIP5gFcxOYlRpEcI6arLAqGrnkHz2LgzT1CpJVaPikofUup5
MABM52E9u+0+eaPsyTwJHCoAPFbUcQO+PtJnvug7WYbl+Hh9FHbKxUrfn8qUWMWX
B0oVxY8yB0PCis/VUoWbkjujjqqxqA/Ioa/EzC+vamQuLCl+gzQqBDgF/nOOPKPE
xvm+SmcGoxNhMbZYBWHHI48rXw6ohL0UeaS03+lQiL8bTJKh46H1fmLbddOrZwZ5
LkPdPWIPPDeNl+FzsqduHFpkXuaMC0j67bx+TpEk2g78Hic7jg4qvg9yqNbszFY+
dEv48N6WRHJrINuwPI8B6c5EcnNRgyTjHbnlHVWSBbpR+/R34FggJmXOgX3wnAY6
7ZppL4+t/SIb0FO4aPwGc/u+nOCQxzyLpEVV57snjifxv25QYgZjyPoZHfHT52Xb
3LKtrAZB11agzA8ahjuAOqFXRwcK71TXEeC3ngSRhaEd3jAZbQ+E9TeUZl8GdTJy
DYPrrhV4vTquS26RFO6IdQEDRlgQymANoUAAqceKFqy63f0KhnY+8RI9GBLjoA0x
lBNnWJju1zkY/jwHpMibe7zocaRPsocKX7SOMkzZsKwm6CkzekQlDnjR0JWuhHnP
CtROWwSva/PeLS0ADCg1WJANuXKRur2wHO+R+uefMHJOEL2E8nW46H8tdwAvRo9D
gBqCp3mH1MUZpu2iccRJbinlCkSt+SdGZjpwUnyV09f70vntHU/7eqZ4o4DtEXuY
vn/R+Fk9rM8ICX3FIIsZ9ngmfJRcWxCEFpvx+7XlnQOr37le9j8N2GjOwk08k7de
2P4iM4dvc89IegttB83wOtY+U/ITwmhb/MepsjGvihAJQ9y6vveP2AnAlcJcwN80
7tpBJHxMvdwasbnP9TLLRi/FzO5rzRT7MZfZSj7Tt004ecsvpYzJSbjkf1riVbhH
MrPuIHO2hvEiMjMl7AfQ9vAOhyk5x6agRB+COsqiDQmnf8bqO/Uol56iwIJXLo8O
H4hbhBSdMhKnFmY36y5pqLBBjVBg4Qb6WtW3rYii0ozZuQtXOZN9E+RslGiWQto/
kgGlWh+od+HpkoATZRyAZlgCyaj9tGKuQv+z8JdHDyMcNTRkfV63O9W7COb1JTrX
Afy5LlzoIQVyxn5gfl/5rvvXi1Brd7BA2jSKZdz5Rs+NGwJUUOlbpZAyidEbZ2KL
F07jfey3ZrDXE2Y/NrccZCpnhBnGgJ1pans/TJyMqSEL0ukuUqb1PBE98Fd2J6/Y
7OeODFx1ActxxSsTmZmRLauf58WzzLZ1dnf0D1F7W3NgCHbL/3WNoxMzbOQ2863O
kkfHEXZmr8MA4B2KecjKKMGgNjJHn629IRXBcOlpWgTF6T/4Pl5MQ97Xlcv7YFrh
6Tlv1TwAFGEwGZquaFwFC1sp/EyrCD2zGPBneY63X7u8sz3GLUJDCgOg4YpNnavG
YUoXPYSrszFkGfDc1LMWWkAbEMHqNtyYFMYQBTUFFKR7wSrYJrP/pdRGsiMKDsQ0
GxZcSN64BGWPbPf3YR7AOLoJxIUOs4OX/lFDoWNXNmxaX8KEA1bSY7moyzuM9UR8
PL5mSCRdHwRhYv1RQssLCvzkw0wzsbESIEFTsleH8BElcRLKnoFPK6EwKsWWyXXB
Uu1b56CVgkq4g0RJFOlr6rHC84YP2w4VZy9ICJcqHxynDltoP8bxu420nDvca6dp
AdI+Kqi58h3hp9N4VMyK+9X8h3PM2vKdCEpbGUdM0mCnyaNN/2fEIMljWWEYLydd
aVB7O29nvLuMXLpyXZIE+d8OSbIXvWEErfc+IJouFXdUVsTVtay6WZ9N1NbA80YX
XgoTMb+9G2tIEdD50Yu8S7vgE2j3exuXG7JfVBxlpDV8xDqwDDKQBObPuy3DOuEY
2tWmaXJx0ueAgmad2DSJl3hbKPtjV+q5yfcaK7nurkplH+LdMC5fMyhDIj80JtgV
Cilokc7P9HHsLNbjUzSeNmy0j5uQ8BwNsp7sBHT+EjYunzJCCG5x4ZPJwPelk/C7
CnbKwJzxjn2ec2idBPjAv+rrhvQaCJgW2VYL7RJn/rJf/ynN+BwfBi+LN+3PJP+W
dGYhE4aqu6vtDwT/Xcij681Ru7Dbjs/J0+s1fSgFgyjbIZOztmi7FvsadVuWx7lL
KQ5jvaJfICl3eQ9TsLBzBrPqLGWerQAI/YTBoRTCFJIrkWrB7p83CJcb2damMIJc
IdlgXjWbUR4S0zRVxdvbkKBnFEBOWM4n9iFDNnE/xveX11Q4RXJAV24pgBOO9tIF
Fg5UwuPRswW8rSfpAOXfDhiaVKBXhNrBSrfeBCajCTJAziHP0Lw01BWaBVbQfk4c
UPY+BHOmXJfmrvosEUYNlMiDG+O6qDDwnrHhP14T1C/Q4RHZDDY2nEprBUUtLs8i
QrnNIugA8G36rzlsZvrF6Auoj+WAPMJWRIZYeLapXNTkheFAY1DOpkzclMH5mgDY
H+mFjQpeM/rYvlYWI/KdlTDValRhwH6oYUi8iTYeJAMgvgKY5yLsY9zjzd1aoTZa
FgImEqFHKquvDbdKyQfj7tXKR7C7tyMnwqvnuBK4uy4PglM77yWFkS5sy18ehI1T
6faPkv+Um4d5oFVWZJHbx7kSoptKRsl7incFNDIvh7GSIIQN6YHr9W4kY6RIS5ni
CoAU+hYrM6NUHd1UerthfC6fVyr36UHSxjAMBWgpPz/g5WpSR8Gg5IoJa0/xGrxs
fe9bH+HiEyyqPGCxQnRfAMI+O3qoSZZbCkOqDxgFuATJnnC2bNlmK2mlgPKB5WiH
wqFdXyBOSuZtS1DWJoiirtt58OWYUkPkRHwg5IGUm32e2CL8k+5xdSR4Z/fN2rM1
aJVpAyEqHay578rXVy8HA8Kep64AUolodTwnJXjEyT5Tq24JN/+/mti+G7P5fMKx
QNZadRZ0vvU8X+oZ8/yIE5LzuNXylAdDqqIsREBIh7ANCpWWih+F6LGf9liiPGLE
8Vwyy7X9qcVDFCBj12b6ytG99iLjd7L5CCHeuE/YEylUyLr8Acc+XTJy3Rh1O7We
Qx3OzCNIefPwUi51xQc1BAwz0pM2xhM+OXGaUC72dV9Y0yilOPJwnCwhrZYlugey
cn1CZvrXJLPKvzsA9TeCp6XcViencmwZDAbaPhyHA3Qnw7iyJYVWDCvdsASd8Fyf
lLKrEHQDlepVpsD5qdWYTILI3rOwEVHO+h05TXXTQ9OPEYHeVbkp+LrXyRjH8TtG
N08xTd050ylggmToAIXpceo3aSttlmPfDjfmytZHm16rw6a1OmTC+sTB0olfHm92
O7/VE4jKpjmhNMV5bjUbCjCjvjIkpye+lpmRKWzv5WGQjdzIf0JHD+apBTX8HCqz
tSvvIeKvJk8lRnIub37ZuJQAvFN0V9jmB4/Ti7SBhTAkKL7djDBAyxNy0z4wajqR
h2Al0BTeOwxGJJi4WCCTTNiHnTNzMSHeEvDqoY3vxPlVG20tX4qxOy2TMG0NlLWp
9OXQoAnebDYcFgXGkBCKEniD5ttTdNz7Er1LHQrq6kiNleQR4sYtsdybIuEjUxLG
q5xu1IRVl8ARzpCKNlJLkm4wwg1Mz4SYP6bG40n/Asng8Lvk7s1PNWb3dX6u/Nt/
niY/IN5p/Z3GnwsPe1mD9MwEQkILmi3MBDpGI2OwcocZV549WLhCNv4QwWp2xMrg
xHQ01CxjJIGsSgNVNVdtjQFkUoALzKg1x7iz9g1Bfjsef8/Z++w2bwrGt1HnEyBs
/MOZu7MlCBy2+3//Uee70DmQYPSQXLTwDCp0f7GMA5Qb31VMbRKtvfP83oMMBr15
MCMNsHmfw3ZOfzYpIAYcXUAwAOI6rx16mDZSWR/hrvxvEsC40Cli9JA4uukbWUdx
q6osO38E/Als7Q4t6b7dc6dYP20CaXEMYJi4T0MohU0MxEaS8LQlp1GCQ0QCueo7
ZTyEj5PmTFLjlgGbXmNtykCBoSkGJiS9uOqlhfPLpA/umhxS0tIW7UqLB8d6Yt3i
w8lQQ0RuZDOeEIwZkF6MaI/lVvkZe7DKLrPSypHH4+CKXjfno55Xfct2OM76rAaS
eueWdOcLL0HhMDpCVZhykRweNPxOcQVPlRr5HrFLvIiM6tn8izK44l3oo/Vl967a
/O7t4nvaNsXTStLxe6bxhxUpYEY60HYrirOFfJXZ32jrDFdPzYaiFanmv77vIiok
WVa/Is5pE5RX8rV727Fa+2tsXd4OmalCqHDrEWZhKdrGxbMo/oXFP5EX982npk0t
0ONzhrMgxTF8vy0iYZ03cBN4Z8PRpC/lIIRjDuCa49to3hC+4VzsYUHqRmSgB6DR
NJjrxqRJCnom4w0ctet6Q5agnHEyqDG+QDphEu/R6sN52LnIo/AVQbN7oWGtjH40
vfJrPLh5SG9YnSL6m9UaTTOCjW7WFpyA8I8sK+5my0rMAuAlHxBgDd+EjckFkAXi
vhvljpvwHZIticMrFv+n05vP2Qs15SizDHqBEV/YwGGKhAdFfOkxUrWy70uDXvnH
BCU/E1RFDhMYwduxZG9y0lHmphXHuV4sdVhB0HIFkhxPcyCZArJf4byQEjzBq0oo
MUtgAAQR1uN1dqR8sJgChPFkmc/Dky6mY5yuopGoglA7Ey49LBWWhhxpFCGc5vI3
uQFQv1M+IieCWoLmfyH2KjbNMjSXeMU9ttwYoGspoD4kERAQ0T3XNIKd81U39JBS
o+QBAUf9RyUJpknyXG/05D8VlvaPH1T7bIBdjp64NcC54tEkY6IovDbNKu6V9B4+
YY+9VvHS+7vjHDdAK6luW4aSlVQqJjbNnHKYQJYK+uk5fm9ueYbDXRqu4TopzZF9
Yx1wt1xAKGSAaq9sHkZ3uJ+uzXNsaryXhquclKuQXW32AnBhlltZRZdemyNxZMhP
eJZzFJ1e85a4m5Fl0Zr1UaZGYyaAHmF98RbXoTXiuwdtBl0lLVTD+XrMVifIKZ1W
XTwGOJLbal9XV/w7lCAep223p65pBtz4ipOXa5Gi6sI+gUSUSbV7BlNP2idLf8xO
VkH2LtJlhP7DLR0jGNdT32z8MfBRkVCtiti036t8+JQiRd2w/7/I/3SUlWC+R6DH
xydyn9XlvMFailwhN24CbZjlOiuqK5JulWEzDz9xEm+WP1j6WvY5fII88gVDSJ1/
bvfn0fwUoUsTqtq/sJzTQyKrAw5HW2s2w8YF6m21PfJF1sIz8Imo2yQVn8nw/cYX
zJ4+rsD2kYiI9ehqgEjNzF07zt5mOAIhx1ivhObhE0PBTPI5E7zwGFquj8lA6JO1
Cv697Cfzpe13XwWGVs9EakPT0N0ouTMaljGF31WatyztJ3MVfQzA2Vlw6+F62Cb/
RHNf02PnPiewLj09Z1kKS0K5cQrJmmPUZ8aXYJxqBwuhbL/oN1WCE7PunifzsBQd
8fx3rOUf2MiX6qTI9sidhhvb1aIGu3HZvakWQ71cp1jE0NTTITTtZW0PGObxcwm1
IFGOOAtgQvoLimNZkz0pEjeAswfGFPSAagm3iBFWFyT91FdFSSFknM3jRIYP8tPW
Q08BK6qulUlFq/+LQZER174tzuPKNGd+AhkVHcIOQIgQ+7V3GtEtiQjE+WXc7yGh
48qvD527oU1eg1jM7N4VKztDJ+hDae5/eWz1gzLr+fNUB5ITnP07shaKAi5VBoFD
6NC+NBR0FpXc1t2kbODBLnWr4Otcj0QD8mU8a0c+xtR19NsxizHt8EsdZUV0nMyz
uTNASc0D3r9545/7iAPPVSk8a5jx4Vn84Th3GFBnXfnt/x/1oegvHDvGmO0wnTHg
aYEjQt3qNkKCuXFYrIOasswLMlGWcougsHPEumVcMYa8AKf7yDR01X03uP0E8AVv
Fftu/FRSH7Ndvh6+NKiI+wXY1WWJzvGkprtZvBlCUCz81A4HrhPV3geEBZ2s8MJv
HUp5pLcUhZb/CkNesgvJWT/f9FEa2u7SX4guA/pTK4X7kQKHd8D8lCaF6QlA3ncz
2MNccEPjq96fhaHl/0pEW/p96ZPkzlEMqJD4IfAgHcKQxGC5E7GoXujd14eP6EPD
PT7PiH5KMb6ld17kueZNTeW4rCj4+KS4msg3jOxewru0Vg8PVllhYPVtZlBPTMcS
DvadPjFLOsZtXz5X68diqbc07TGfydMtEYcU0GYWnahEqVOk2aBeTsAAOtE/LvsQ
woepjPdjibuQ6DS6S90X5Khc2N1hSwIRhJQcXNZPKtExsjBrSdwdP9Y00keu6wtW
yE4csmC+uMAGqnpxhKiZ0M4vKIGf6YLXRJ7+0OmMb2i0udky61I/jpTDpf4FXkOu
zgumaQoLLPnROeyGvf6jKCia79DCd48/rVq1hFcLbAYwm85H/yCdbp/rhh11qznT
/XQ7mpTsBkZ4SttcbYoAgWJ7IIY28gM+hFNlyBMZ1Wcr0ENEbBbjALRbsVTA8MlW
LDhGnBsRW8UOiVxC+JlPD5zNiFfi9KxyJ1ae+DZq40Ygw6cbGLzej+UlrcFuC/+5
KzDQ/8A7jji3h95gFJUEX+JPY2Z9kWcDeUQ1T4ITogksJTWAS5BXeaAn/iLUQjmE
FebmfMh0DuGCCdpJEfrWJC//lZoLbxgXJKjdrA/k9hiSUrTVYb+aLLG1rqB3sZoi
IYiK3iZJuGpXlRk4hZtKPcWyhwQf9cGjjiG+lMq6u75CYKYBiDpc7twxCXkKWfBa
Z21jrQgJS5LH5WPhWZSn5fKf+W+W87m20ztJiLuy2Do4JY3I7h6oxrdw8ICsJdp4
cFifGsHGOD9zgbD14Ecpj3QiDtPFD4DFcZtLTAACHddU0kqgLZPG3P6psycIsRdO
pQWBy/RZc2AlMmic+pbYV/QyimU+dfMZA82anVOgxnDNwLABrRhIHNWk0Iv9RnbF
tJe6HdElR4T8u5Hf6H2KpeX9ujzZ928PoI3whoCePc8Jd3fVSyKs749l/pWiHvzW
9LFxZyyBOPJJObBBuril69qO78EZjBeF+1FhQWfCUgds6gstgnTNi4Rsfk0Cwk3y
yBPV4O7/fn0GN42NPiYnWXKyBvORD2peK9HBPzOWBAxDYG5AZS9Fxh3JNipw6Z/O
XW7HHbT50ttK/c9oD8SOMEluFm+oIc3HQINhS22XhJdHwD+OjvVeEMYsegjsVYu5
jCthzhVLjKL6nE9HKMeVtDPC/SjGbC5J+3BDSFx/AP5zdamPd7n5gDfOuJ6ZMPyz
nmoxaDE7uEBaD+bSOJl4LrUcPRevLEsH7DRwSM53ze0Q29Yn87NJ47UbPpOVyafT
jX2V33Z87iDjFwtXQbM3cGJOQ4PuztkwgO8u1C0XR8QUDYV2GNPph99BFIF9jzES
D4Si6Rb2S+OOQljonPXEofzw9u9VyKHh1rtfkWZc/X4GDRjBYBWlXYKTcuuvL42H
Wd6d7B5Vppms1j22Ri9Tl4kh+IOpLh5JnePZ25Rip1ZJ3I3xRC5aofszNE+rGPTi
Kc+GsZI7VgeTJdl3LC0302qs9MZkJwPM6Si+Q/zAyCh53LsWQiCcxS9Poc5nSdtL
VBA0Nc0JDO8g79UwWtm8AgwKlpt4A15wz9BmakNbQcSw0jSOrZ5G+aMlRMqGILeF
du+Tg90dQxQnyBzahVATTa4j6RU9Y4KO4TGpOrRdVdhkHYJ77Sxp0Ycep/KjtkZc
1/e5lxGK4FCqxrusCw/uA0j9kTHIG1rp75Dam6RRY1UKAudSVXYobFsIeu43NBX5
L2mnW2ikaVLMKKdhyGvKONqzDk897VOwpyyzGzsK/E3UiD+JfKiSFlaKGyXzZkeM
kEUyULEDMfapdRJGV6Pp4UcCjAkJzvG7mnF/P4l7U2dxY4l4QFQQ20r3oZIHL1SK
opBJBCp3CfI/34dGco32K7tSQe7WxD0h5rPshbLuNEm8p5g+jmWXpAKpXlgx8m7o
1E4ibxG64lcjtD4e8wi4U7qnhZQLg7FLVfwkq42HX+U7ITYl32xw/7OA1yXYhLQi
NdU9CLFhNz7HTTYF9ZwUbZxqVQ2Si82crW+DY8btAACr41x400uU8AORq4ua6KkB
5LlvGWZdClCzM5veDpg3Ea4NRDCvVW2rC/uV2WxAg6dJSTtGuuFbO0dZkLYzRhzk
n3R2bJEz/11lMVyoi2F2aqjq9Tk2RI8BFUKq5PWRUWlmfueMhNLL+aBUcAfVYV+Q
OPC0+QAn13tFSHHIqpsdZXlzigLfEtw1ZwuxcWMLXT02W4SUDP4OAhtyT+QPOu5Y
DZJwtg3pSHV/uJ3iBVskV13vWopEUqUGOk/XV94VzchA5KHbaC647mIjZ3NF6NiH
E5i7yyBis5eHZqzBZeo5H2G6Py50gB4SOqg7dwCugcYr+6tBSRBWoVO8NAhtFDOd
0owJSPllYtW6whxWmgTbrim4DwApvW4wycUGF+xo47Bp/FtVsmoMhTeOSX8bOmo+
jZwA7ri8edCxQluWCYxnwDXPmPv2pgjHX/vII9aOBcVRGDAfpSxMjZq0UuxoWGcu
D6StYTIL56P9Yez7EsrvvnH0x+ji8FOI1/JF9EDdHZDfaZOxDWOPuUj92kDbgy/+
R3eZ4KNU04aO+AxpOwpecNPRfxIAG//IpbqOEdQ1aDuiACiF94zxPbSGo7rB569z
uPbx5ghVqiYviUKUI4YouWgYmFBrvILBgTAr6lEftyheU2ZCBtTpltfqgYdh+Cxh
7dvbiLYa+ToNlgeSfHQMi0JuaGL+bxLmxbZAump1GCOtsuq4TZTPll0txppVNcDl
lb72gN/wREegVzWswswrYmL9gZM7Ma4oHohUo6GMKMpNoJaut6FCBut7nN+0blJd
oD12PDnFJ8XOHrl915aYbEqTfqHlpKizrr55KFAbKsb64E3cDoCPOICIwh/ey5YM
3U86HXh66PWDyVc1K7oxcN4Lv/Lw5m7eWFj2RfZCQ08j9Erms9nHwDFhdBfeGZAM
2O4GCZHlzXdHvxI4zq4ryYWWWQQMorAXulG6vArL4XT8yxyFOcMWLNzkYObfeRUu
0rQBA4N3tDjttVbQCEhbes+8qbuAPZL9LCR+uIvcTGjl0laJDWrSaaEVROuNXcyr
+RqkamVFLfQz1jnTscKONxg5SGStp85URFg20oJTS0AAHxkvOlhpSAKO7A52KrNs
iPGR4by1gXkzwga61WVDCx4upVAIuW6CkL735S8D93kgSX0GUCM10lq2ZrStHvCp
4+PXNSaCOU9fnN8taCnCLPRIO3Ry0+JT83FXYwGUM0fhrGKQi6JufrAcC0uQfN99
N51APxURXcFMaA0fyT0wxlndVkVdQ69sluSpqeGpNz9z4RVhmIQ365/kribA597z
QMQRNl45GWvE+q+AQ8SttB4DrgzMLRocKaesqMuje2n5C4+vTKVFkrsN8JFwv++d
XYzg/yqMqppTDwO1qKpSCGF2sejVD4DAiIKdxPvVVpguLoLNrjJzMUApvPEzo6TZ
VZkZe3rVMI8EbVf3GisczhFY8yB+cP20TsHg7Gh51cqAHhZdNBkekViDw+KnEQlD
xSwCkpo6Chqw75V+BWZdE6FVmyhvs1j9I67xl+L8FGKtKCAPgt2oroksxqDflhIT
2c6q/kw6kQ6+NlR8+0v8uL3hQBnM9UF7U3msSnHm0UFCfBLLhlZpXR/Ne5pnoI43
C72fPbtrELC/S3G/FyS3I9sq8Va24PChWvE4/doLwE0wsqG9PlT8oQ/eDemRDNVk
Zystmncl5DiDU31cccq8deFb6nLMqA2BNv0lBpAgtKlyUj07/yYLg/XwWrKFBiGp
KU+/o45vnFCkZsdZQ3YcKojyltviYEEPdj+sQOBlXQgNpWx99TghjPvdglprmqeb
Q91t6BFrgVju/TcCZv3bd2KSvTc2IMsS3TAE+9PmogG296aun0ruW1ZRqjm7oRvB
t1P4szBrOCDP85NltlG/Mg4Bd37r1kOUF24ExK7v+5b/UB85r7hJU+7Q99L3o2Hj
7OR4nGnulBcHMzlueQJazscloYWcPidnwWQPh+FPkKrNLjokyUDNBbe9yZxnrOJk
yoLrQoemKZvPhFjcpM4mCR/O1zV/DVuhUPdGhgsQjsUDrtzMw/GP1Uc3wq3pOao0
qkn+Ow/cfKxdeGiPIXz9B7/cZWWrEf4sWzUVMig1zc0Lg7LLXhQZnA19zoKcVnMI
ufwugz2Hx5UnnqVRf3TIdvoqwuyBWpV83bTtfqiJU69DRLGbF7ViCvvao0JNlnxa
7b/bYhTz34NOJe0Uv+bkIU1hm6/LuylQRTBHm9/DSYsDgegCHQ0Y3OOOQpBi8Vdp
2Q2Ob7zdIXDU3Dfh1FxS2CPtzu7Dd6mSPfeflCeY3oQdNlMgkTIqSoSvhtP8PqON
Yb/z+xRxbqvn3sMTgtItT4kIQwGekMDyjYNxJsOwrK4WNRKS+furSXNqXHRv783H
kmWdjfYlRmfU9h1PhOXBSYkeKJduRy/+SgAZSf9Lokqf183owOjMy30q7m7HI7q0
TM3LSnr7YlKs73miqBoLuwTSITVkEG2f3PJxQNaRwC8snw7LOoq04t4JqVfPmVSO
GoUuv9V2mWpr5UPGHWY19RlluJPXz6SlyEDNVdfZ9cvJM5Ig0/HhwWwcYCAk+6ML
W10tr5TZTVwvaRBIh4O/qlA9TuQfi8PfdcVGYivXm6fW19XixtCcXg90dQ2Hkqe5
2dYg1EV/raJwDIAz65IUeGFmP56fhFUeSTms+f5u+p0LPYERy/kvH6E8ZHyEQNHG
ywTJ+9yU4N5dChbDvTKApCJ7COCZAVTxIWgcxTLymzEfXhNxuHU/lGIh/LV9Q7Ve
nnq03AqZkvc/9v0HzHm6f1O4OiQg7OmkZDKsY0Q2f4XSzuiTLFq76PwS1x/49pxY
edyAU7gED9D7dpO5JZfOTJ6k8eNacdYbvR5oC9FB4NmBBZHl0vJhjdSjpGR2wgrG
KtAfLeUcwFa43srqgdReS0tLWF4EGAPGfhunpTWevu5pLUB8RomTVmYcQITCPyxl
tMVMRNL5m6xsw5jlovSNjlHNZm80KYzSwmrwy+MsStsM9PtzRd48Wna5sMofxxnV
zmbrFVpOgpSO5zUos2PwjpPtWX9tdR5JB9sEnYS6sRdGGk/9F4wfQMamNI38A3Ed
DGHY9sUy+g9H004F001PUu/DRuKd0aX053wGMCqBzThZj83YRxbfW4nmmZhKD6Qj
FP5eh3s+MeHXlskDmQ9tx1v6NXSWr3J6FcJ0rKVe3A6QFE6pzP/BacywaM5KcMJQ
ZXfHcBr3UV/ugLF3Pl8i0ukomwt11z7GHFSHuk8eTfCGvBbijQkgC0HYySIS0/BI
VCwMkHOp+8NFAzfmZGT9PyJGCSlQtctC7Uvv/8doineOOtyvSKkCL48zMjutzyAb
aePRW6yMeEC8lca7N9sjRBWDWswsF5DwDeyp8Lq9MhGGu+jBsW0AS5I31LycWr2x
Fo6jDZsioafGGleAUGB7qlh1VpCJPfFgEKr50DuwsDm5IYp379YC4V5T8KhNB8Hy
f5dDsQUlrSoDzdqNnIqVSKNT53u3dWlMCLIo8hyFAP4DJCLTVIexbs6TTOBJoQNT
T+m9n6RUmRPxznxYUWGuBjwgcyTjcthmNsyYlN+wEPjQMEQNS/FYDJ17mSc36VDk
N7DrJm3UUpGU7xeLUfnfILwqaGKQasExDAfY+11eczwYX0UqWpEUCIp0k0Tz1QQl
f/vZXuM57/lpZbHNdkFm20Oxl6crTeXOQWKqbWX+nveklVTa1EUoV1GXnXMxC77a
LO+dKUswHNXZwd3wOrDkyrPR2PQy5t4xPeb5IuIG23ntl23npEAQM2lbAhpH5GaK
x5LtJ7w+u2tKhysmr326rHAtDtpW3pJbchXutF9QaOKzARuWKN4MYIFYGAStfb5s
MlEyk+dFbCre7kKEM9gx6Ezhx47feDFrV6EeGob0v9/u/fTGulrcFA3Z08SNaVPJ
0Cqiq0dKj1REDjki7jQeFKiiDd+fJA7eJDiKCpSIBQZf9BRwmV7GvJWwOGI3FpCo
N8SXINUFzDvNj3jLUudnc3/lIWyB6MP06se3IN2uFg6XUJGEOe7JzufaCveUjvdy
c1V22i1XIGI8b+5ULJ8E7Yt2BOXlEPl5uEjSUz9urDEUuPL8RBxAA0K59iB30CF2
P5WLIuHZJ90z3C5xd4D2SnfeFcOvW6B8mKmIIRVlzv7eiDV8DyV8aZMgkJZuO+Qs
Hx27r/+QqmVxUUAqHGOKk8qBX0mvJ4DFsxPZf8MeSKqTB7sazM4LnFdMHv/DfhZM
myy3Rv9ALfniNwQQoz9IM1OiPQzPvQAwhirqEYDlTYtv9/WwAXCRbzc5eiV8AeD5
ye23gTvPbXHYYrF/bNCFX+6cpb2sNudt01HG04wVvsjGMB62j9r6kPTa7vWnf6ll
XX0r67/M9dEwNu7WSw3hXCc4yHlHqsaGf2ZF6Eh6cz+NIlx2TPbtLo7cnkYasSE1
iCmX9NQPyFIMKeCVXdegz8yi3z7wA8AtftkJt9K67naU4o4pXTvx7rfMD4auyUXs
8AgUu1HBIiytyuGDvXDbYhRsZ+rZxRXt8yDpmLzO1Q5ycBPGD0Mx5Hq6i5yYBDJI
sdV+DADH0xk3C1ZhqGwfqdjjpN1ZslPTp3BkOIOgyHeauOYHuW3mI1woaL0TUES1
BprxhDqZ91OLSzM4vwcmUOJQfj122XJ2Ldhicbhtq26nvhuRnblXzwTJAub4bBzR
544TuQe1NiKSlTnXa4cjSjP45bL5FOpxJsVDRIOJS0dehh8Gh3C+C5BNZF/X5R3C
IZv2CiHTSvNcw0VevpLZKRW08Qgr1BZIs9b2V7lxHjlX2/o/TKpdi/+jpipxuHqW
FcAHrB5A2c5wC6gVePoGGicavZGDcMbAtcmBfaqd3O4wdmQm+NsFJepE/aFVkEuc
+Wc8Ksj6FU4dnuNXZasF56CD7MEBpx1hbo+DLt18h2f1Nd5HLjwvYAsHCHy7TA1s
c3RT8uRhvw3rdWTDHx1q3BYfeJ99FN7zNIEfIgPXsg/TQOWM+paE3jCeQXiAbUVb
L6tutzzyoRiGQhD9rgFCaRwTEhW5logV31MdjjCINuUsUzXohEOpdhvzMl6JxYmg
pYbR91b8+Xwd00YuIgvELIJ3oQOW/Oads7eRB3bd5TZSH2qgziv4ZEA48lNjv1aP
QwweFwLLuh8Xp90HyA6CuJXAndu/GKx+RGhjyuq0/ByS/CCoHVvJDNuh6ik4IOT7
R0Acp7TdbGmh6aYsR+0ElSOqVfFGTcYQJboDfud/9ScqCCndZPilBSyYYd8yx9Iy
rFgGnCM5DFOTh0eoEhgmMx9iqhvXHPRg5g9cM8Zgsywdiarwe8M9IkCeuoshR3KW
CHcGP8F4ANeJfSg+QYZ4RImWTiZlOo8obbpHco2cxAFZWaQu3U6+HnGAugjrZ9oR
Vw4xHQxLHI7F/YAWwtXu+zpVHnwr91NT2+akYf1kkY7gDjHKuG+BTOznUZCzy/lw
z7yvBm85DYWcZEqrgVjkrOhLeP57sLXerlgVuTXpefOTpazElnnI4Zt+Ys/vgoOX
pCe78Iqf0u5/8c3erZ52VBIwcOpA5QcqMbqYMMBv/qJtpcZF9R58RUPDciQHC0ts
SdeUN9LimiRM5w9WcAl6TN9S8TnFk7CxgsPEBh3V5lszL0VtXxv00hsRhJFhcOvZ
aFegmkT8E54kWkZma76JHWeZ8ITDhKI1Hr0fVrwO84G6D4Ec4o9+OlwtSCuLMAev
Z3lhweSqhU2m4GH6j091adgSJVu2XnkkdmCEA4YZYH9y4ru5/x6yVzH0OfAr8sXf
uZpkGADZMWBD3tSavBC0QEzdVyDyNGEseuNbKk80Am2w3A83SahnfHYKfmNLkG7J
AplUTdvMBHeDr0gLfOQCvl33saDO034o2gaXDJT3HxMPoGmWCsFWL7UdTanObj7c
wXqmr9QjpZAflvPRfeRNvtZsj3yKX1bZSfklNY5aRFbbCIRA7H2DDFqAeolVqOxP
ZIvrLWioz5l55Phrtj0ApbDxTUjCpFPelA1R7zOhJY1l/uoCQ+z/mbd1COq6mgJk
plhnbIky77gEKCnc3IXnv4p49fIG5OUUjTXOCVks++6zkKRkJHEXgBW3v+mpl6LC
XE7IYWHxOw1WK3YpjuPQCrBHrUUKiuvd/f6oXX3nWpEzyrKJ72Mpp8w+YQC9CBCr
6xkJaZVx2zqr9OOo3yHizzhN4iT1XlE9V5UcCxmwqxuBr6sn65hIWjYT4NUSwGRT
d4zrKDavr7g7Up+mNdkA+aMCFq3opxkU2DlxDMm48j1m2ds5JaCSLT8blnoAzxKU
NbH0EijZm0uFamjD9q0EJkY5nCbdbg1+SpQ3wTX63Q7bMb4jld7fEghDw3OXMc6I
k9FiEIChAnuIm47UnB6HACtiZaDq2SdbYAsbcZ/W2u0bX3MuTZHghf08/DeWJO3E
YEs+j5xFMYlSUz/1ZGcZ2lHisL634QYTLPEtSZgqA0KjpYjPxBkK7VsC/yQ0/1PM
STpBfTNgKGdFcwQg3AERIJwC6AZFfrqiiEUyQnYS7yLoZt4r6TbghYl+iZXTVkUY
VyJIPgPeajcsGDG2SIiJ6fsehrXjHEV+tsE7gKqJvTKoORoLLXeINNX/eKzVkYGU
FLNj7O/9NtPxoxfmIHXwiqewWuSKB6+1D1jDGrMcDEtNZf+Gb1KO2+K595XuxNSh
LjdTmR+cHiEABQQqwyok1PcjR+UOEBjU/vixIrEsfTqYgQuw53w57zdjThYIvnDR
sjDdYR4hun8kXSTFyPwQNeeANujGI/YJUCOLYx3Szeo7cgt0Y0BBg9zReJH2zDsw
JPjPsEg4PD2LCnVB7l+VVC7w98OIxEUHrYNAPxhlA3KDNaI7J5XCWOPTkii/vjKK
kI8H2FHMDPM6sly8CvXsrYLrx9ofR0siqz/WL9akjvHGCD9XNYTxv+4fDeUwgsQf
iZylMcdrtaCUANvwGOmwtvjMaVWnt3MzcIrjdCGZtsvkkH/KV523Lcb35Stdx9ya
8H6Tu3k6+jEkDgLW+XJaiLuX3igcK+sLsDB4UCtlPlPDKIA0Pfdyz1UMxZsVPhyT
pd2kMWs2F+9rx6lwiOwBwlaUGcy0KyCsVWizrdJJ+q9njyBwIoozMl+vHmGLDUIx
3En0OF+8rJO2tM93b6m0wTqe5ip/vLzWs6ebt39TSobOAlOJC/otdAlnPsTRiIQx
MKcmwfrmADXzyNKHDJN5RCCgPJuC7XXaYzUXtybhcewtlxWc+uJr+ik71ogRtLmW
jIW4+PWS84OVKVHr3pTBNIADwHR4pIso3dqDlK8QjbK1dbiRL8B+iHG+f108unZq
GOO5+fZM+H9M/hBovQzXa/WuvscAeWgDfHusZ7zForFHx6oCGPHbsSzyvLM6Fi9t
/LRfTVVRPQRcRztR/NAM3CemXp917Q4GUhwq9mM4xJZg82vZl3p62rhHWejNcnt4
a0rQjBjK0YQhHhFHOCVWGKsKEsvodAwBiL+F11OVxW7XprOcrJXjEywgXNNXx+OY
XPYyWa/B4uHawbJKli7qpKDiigm/3Z6KDzLk2dezlxxQbs5ynEC8fHFePTGT44VC
WSkrT/Pt6U+o5HhXP6Q+L5uzO+jnHlJQye5/Guz1VBBdUdv4YvotXQyu+mPIslsf
XNwQxx2P8IDJLlAgGAMIRPOuAkiWc/6yIEY98V03vfaj0e9pp5rcNd5xQv/SE9xj
rOrbhTuEty5lNcbyPLIPJ9h+J0lgBRgNpBUbAbEfwfXinXAf2cB9rZGYrORK/dbw
25t8AHxGJCH8twVreVh0K3Pm8IVhrSvryEz/iaOWCtRP7zG8hA/NF39W3TP1x3Nw
a8SvBOB3vJTLPtDvp+5xt77R9Eezh/bgdDwTxnLs5jZiIEac9B3QD8vWhdIJGZcw
CCJj4xt9OTZSYp66BpXpuaBnAkjJDf7VFXD3JL7Ap8QqsaEaWm68nrwYqjWMEY0a
LLVCbk8RRvKhdyHqdP/lKuz4+61j5obbisf0Fpscbqt0NXYuiy5ehnFuoDrDubbM
Y/MaDFoK2/atIC449RD/lWkjzwsMYVMFgFYm0hTfbQ0JmD9YvzOyx0qUN4dA4cbz
pV0uWy55Ga1ahZdMIXd5oczRfvhywOmTnhRRHiFlmpHRcb2lfGrlSmR3ZCMgWvU9
elx3S2dZ+QZ0oC6uwpV3B5sZVMyQBId8r+IIJR9ZyQOfP51Qkr/UnXqPgvDB7hnX
KJvYE9R8fNkbhCTuAH/XOTT3+7Dx32bSfovZmRQAYUjtDk3OnvthxzUh1Bx7NGTO
sN/h4UWehD9Cm2B9zKWVmJO9IhDO7QgTdKXQmlfr/ZYeN+SHpKUTK2hcF8kny/V0
TkS3Ng7wiZCIGDAizrBhLCLHyFXCMnObqNuZSpvioeWEunEBfAVbgfLTxIOmT+oN
SlQKq1Ad8a7dFrRBIDR0sGpNAIMB+h6F7pbWbHsGxgPjUlNyo7dyQ3lOjpdvg5eU
drWfSExsKrBZGQbnv/vv9MQp64R0NNmpDVrPxEXJ8gcEAmFjgTc8i7JlEsjx2mLr
QE1QcCya18JgGvgV3tiufCIIdqFBN8llha+JqCh2cpTYq9A4brU4sK3YRWYd3KzS
t7IUFxz7GY9cse+iWHr3PtDNEzPYdp+vqbpy9IWlsUbKEJHtoH+NFL9oqgByVDxJ
mnrPg8u8KT17SQwFpPiUrhWgySIOq+xn8jCyPCS7+2l71mHCt8VVoqkYKkxQIErd
NbVThiaec/pimrlGSKNyDnehSa3X0+Wh4GzdGPTWyCGRbExgTDrchpxAQC3Tsmnj
A7PWUlPGKCBdlwbL30muqdRZ8qqr7/HCWPpEWb5m6jSIgD+O8UaLYsstuXtbA6iv
VKVHVo7Hx6q5NgQDU5HuLOre0z31A+eqPEd8o2T+ChG2+PeJ1xy/PzOvcUgkvnE1
0ygX63oRKdD7C3sRAWAQmH2ob0CWTgj6f+eIj+DhcrsHxyl3ZCf5WDc4jGK/xCjd
deFHx9wYTF+J72lOvZOdkrIe9rokU81ytqyOuQbLggP5YMtvWLZRNMLNzM2n5na0
VsR9VMvv1R3UWrtENMNbHkkUpNHMOksHeqDjR2iNem79i8xyHzy7ycwkC4kY+0Ov
PCKNo210Hf8Idqtr71jnSsLrRtddJ7dGYfky/qpVZq29MTN/LldXjubNZGoljg5K
9qELLx7MFYraQ6Hewm/PoIJoNl5n/7+DN4WdXUrmdCfySDsXITupCfOgWV7t6Vq1
EEgU04oFHMz4T6TnTgBovyszJyGKAULR4Su8VHbVSKs6L7SX9kwgOneEfqXsgRml
Lm9LGZng0wqZVY8V/gjl5+n0F+RpFX+60sgnQVo6rkQb9GLZHAv+UVYs54LiP1jJ
WWvrKsltbsGAk/X2XAWhiuqcBwRn0Y4I+cN4F6Dk0KvUtbm/25dLocPE+Q0/yk/F
xY7qZGDUqsDpUjLUwknWAn3JWfvlKIszllweRln74W7aZQn4vCNe+wXvThG/Hkj7
3QYEcjnWthbekE2ZhXMLq2TAJEwGcTDa5Z09qZlJu9ds8zx8gTyLk3BIqLg8eQPz
bfAaJ1wUxByS0EcFoSosk//H6E3I2N9yj4KxN4PjqZ/hz7xp8DsMmR8qRnh9HG1e
ypSSHyvaglIFKMtUhAJdsel55WmenSQCZTItT6LIBYbJaZD/kpbKlAguxkZT2BSK
xQnQ0rRspd0DAKuhQdBrnr59TdGykZjL7G6EQqbopM+s2ByQ7AJAoB3hl+lq8txX
3pWzobAaqvbIg5O0EtWv7V4BfjuVCtbFvT1k9m1PRRG44OAoOPi5ssEnnbTB8nLW
BKEQz7UKboAGQihUGARj2JhwEJ4lzt/iMZsomzM9f6DVKrSxJLCpdmPQp/QsPgvP
TtovFy3Bp1TRlYQJ6F/DsniJZE8tpXcxPMtL0KuXmvcqLbC3WihE/BHQilr9d6EH
GCxr2tkwncjNPoovvjWyvTVv0/uXhmqmmkW3+j6ZiFZaOE/SWJp5dduA9erB8306
4Eh6Oto8Mmo/u81wGBCwA7yxn3oIg54CgbH73lzRuqY+5WXen7FXo1w5iJHE0Aqh
L7rM8FkzjdF9XaH3gDn8WvXoK63a+u0zfZ85HtLfGhSGtq7fO4Kvr5D0N49oPbFI
anruEpC3IY0NZgwz0Ubp03mgSnNil9wNnifSEscZgRhmdCWp121061IVShtlXpRd
CFg1n09E80Jdy9/TT0JAVk5JItxeU450lCMaZ7WynTxvcZiDYXKhC1cgQwnNaBLY
pK+qTs6rqGrWWuSLAzuND1ktuSH27qpSk4DiDspbw+R36p9Z65Pjc1XgxTmGyB0p
LSiW+6oJRXDjplrq+k/S7QYqsA9hAjXM8c3C4yreJ2KLI78hnjER6O+Hw11B2u5s
vbrF55WSKaBKXAzXljn/ksQ0c3LJeBsqp7yoAz1rC5PpcYhNeABwWFuXNAYpX8GS
oV5RpZ/etZOeGowT9JxPHVTbsgVOTrXxxusW9H4bEGNYxugPpJurdxqOXeJBKtan
u/OT2CTXieDu4faRrEoy57YTDlSSsXQVbY5ZXg1jMS+z3SGzqDC5yEzcyO68fFiG
8og3lsN2GKb7GmQAyCuDG3YWPjqjsTsba5SInr/CdXsw8pJjdJTIVs5be5prES8J
C4ApcMe6sPzkma94Q4kLV7J34kVcRMjMyAxhMncPFQoFZpDz8MDBg529H7AGiwoa
RjOFEXKquNRKD2IHm8EU+8Bldml+Ai76s4dN3rRChropD/qdQ3y2hQq7ZO/E5YBt
yFkSbVWTEiMTCqfmmIXz+awNIsJvJvAxPxEnIVwNQ2chpg342z34DFfrRuhmW6p/
/e/CeS8WsqO08na7inLk0IUZI6Bubh4lfOSKpteOL1tuX4valKn3RR++qR1WGlKX
D3yq0dyqOSVETlcKxDgiRjblsDKiTwaoQyUcYfkgpZBUih3mx7AMdTaGiVex9Hy+
nn/KWP6bY+DYxaHZXyp9I9QhOhxC0MNNIQyV6skd2iwulmf8dKboi/2GmnzgrZAO
x++sTucvMqNQfxMejLLn8/Y7M02DFsLIvjK4jpUruyOSeCKh9dM63oIs42Ijk5j3
haXxkg4b5Bf9qP1Zxos6qJg8ye6PX1t2dd076Ar+gZCB79JtsV1BmqNPUFV4Y6Us
Wa+C1RlB2pOAde2PH55lfAaCL94fIye6ZQlLBwuN8jFSdMNCz7AyFBnDF2OGsEU1
x7Gaer2wlh3h0bmzbgG7M6ub4NLC7Wh4qQ8YZ3K5mHbyOT4kefuqYlF36EHC6dDm
k/ltiAoEwCP353p5yOswZznoQOgPwv+NrylRu3h+KVuzPl9okAjXEi5Tk273HdkV
qwB9V4TjhRRsYAHVQVRER/DVAazR/53H+kohNhbQ78Q+PAf7MA0+bcQVqBlvoEJL
pSls6VX0q3Bu1agAaO73gJxgnRrYGflLQfRniNTkkfr0lA8kMpaUTYgKJ8AN34oZ
yxWBnz7oW0sRTWhhWD6FEOsdoZHcw5m/k0vDQ6it8yCIPePjl+IQOgHCthtOkNVI
YwPRJp/3C+ff+VlU6M45HBh3qBe4xkK6K9p0ec1GakXp6mC07k6HMYLFj+9OCLeo
as0zd7Z4bMS5mr4Y84n3IggtAd1QEEj+CC3wSpYqTdhP46k4R53RVX6ZW5+04rX6
bcOTfHRac/ARLHBgm530Xe7BMyfQyf1Cmeplmo7MCAt9ZVdnuxQCkWztGLrQiJK0
LhKzoa8UMbfp8tjo99ksJP3036JDssHPtnHKu5SB2BtJnaS5dNgVNz58jsW+Fnut
k7SDvba/sDSDv0ICUHh0dNALkiCHAzNt7baZC7ngoJAHEN8vwQw6maAr9ZDQapho
z+eVRNDJ3boQZCLh/5sZHhfI1w32CIVFwt2YsPccq2La9dTCkQTTHF9wptKcSeKW
MMVI7hpzni2Qq+UD/Utf3aH1Ln0ogqlSOPsvR7+4bjXuYGJNj4uV94dVuNyNSXmY
GhZ5WMW7UaEdPJAmaZqX9AUS4k/XNYE12dOtsPNIO8Q08eDYQSW4D6FuO8UZieZM
w0KVEtC6DBmK1T5qpHgH48hZeYSBuXBvlZwViQc6kfnuymaDLDHDIqbtudXcYdqJ
rPkBv8kEB05YCfyr7KBhn3H4E6WdOBsjZAc62JtRlDUE/cwmSokkhWbMWIM62jf0
tV2kcS+V2SimDoruxoPtgVOrbTR6BZdhcULm/dDJNIN2Rcnh7IqQnIm2EAg9EH93
SdfNjOaDwyMQZ4IIApxr/iJcGACQNymIJNdRTqoNCDjVIEIebzXmOeiNm2QgvSYe
6m1eqv2eCXPm5SZ6J2bCSWIWVbmNsbWh70YjFLLYwAPF8/uXgV31TSOyo9MiLZMn
Cv8Tq0Z9ulGyjqO238X6fJvGfhAIOWIPKN+ePMor/NliRgYF/YuCukewIk6naqMS
Fmv1IYZD635H1NL0KKmZLdkg1NOn6jxnT3uZ5r6swyhoq0jnU7I5oOsgKBg1b5RD
PjUIyJdVyllrhE43DkOYFtIHpUZ6Yy6W7Lcdq2eY/zpa6gxNeA5/JII40nMiVARN
cPx8xkcDHrK2CTb0KHOqRcFU129fMI51HtighrRcB6WkQHJlEbG1/PDxgc/Kzs3J
gfYjDYXGXnS5a07Bg2RrZ7521EiZphNdBjm8P+Z7yiKI7/ctJzTzJXZ2Aan5l3RO
rQJqY7/mnbl6J+sOXH6SIG2kwQp5ray3wJLLak2GjYTGlAOvRFppRay5P6QtGu3O
j/4H3a04vtsJhHTiHgeERJX1n7gTpdzXbdm3bLAwSwOpTfC39gpKuTtNld1b/b2j
JSniIz7mYWuRhs/4aBtu6Z0tLu8Ljrokm6etZIqElpxUFEAVQ5BdM7axB5ZcvH+o
2qoFGjKW6SYlyeRakmfQgCM7nsKE644LjVPMW0fIAnaGGOFS31Jcvhws9thrPOyS
mxcapqg3mFEIo5IW1Dh/kbCs+ZK22m0Lq2dJjnFCg6YF0gO2YKDnaLoYzyr0XHZj
+ScmJukgmpcDk9C7OiySkd0xSN0dE6x2NdjVhQfTLvuKOQ+ta+rxuNcYfHl5sg/e
hJYI646Cnbj5kZKMK2Fj4/hHHagE4T+qn/Hr6nbt2t5VG/tD1zcI5PcccfOrjlKz
kfhJ0yfQnVNzeyqxA/S2dZTSSKX5iKpygUc/2z8lM7VPR4GGFNtebpCt/1wxoUTi
uacXPHQFTKXUGU1HRjATyRz4Tq6ymQJQlwX+V9Uf7EZZ/bF0o2IOiaX7IBwd3W+R
nA7ehFPsjiTCYyvv7LZB/kPEXKAzg6i+0tFoSktJWx9jkBH67Sc3QJdLwFAhgakD
t1sPb9UvxQ2XyFkU1VDUSS2jQUOIpnm2v3cbtWQ7AZJ3zE3K9wdwLdYDNcKfwanR
3w29Pg9XdnJnetuqovIN2aRSz1FogN+R3L8JNRu+4x08BoF32tk0BL4ALUe4rMyU
okQzr6jSkVNqKrDaTK/j77KBhrfAB5BsLN2uuQKk+1L0GbOHXyb6tRGo0nc7xwVs
XPgjn50aFkbk7YRxKX2wqCwJeQ4sPHp1+qOyv4/wNuMjUtSIswdQ5gGVxtZjUqLl
VrZ1LFBDKHtOa3NY6o7/cKfna5BexMNDJry2yOhZvkiiX8zZxy/+9WfbpFMsqpeB
1YrW4yJlGYHlpah/3otdBmKSZeudAEyxTUXI5WmujZJpssvMf+gqM3TEzQnIaFlK
9EfK/+cHi1IhrH/4xNkCt7AqAyFCfe1AdiSmsrfnjs/V4li/xC0/m6wXRXKTe8qx
Wisnu5DrE+7POvCL+OIBOVWxBFElWclvVAiPuqeFQXTJ9Y6KYXbgk9SfInYYUgj9
6khTME89TFjka5KK23FQvc2+qPKjQxp320WU4oXGNvjef2UI71fJSs1OeOg024uZ
iojHDjUAmGruOBNp0iGqb5brRtWBs6Zqd/ChZwUAeuF9+3hAMqMSpYRPssCrP2wJ
nZraRyvw7CWmVugEr5vq2ID8R7e0Bu8i52CZuFx1bMNuHOmLb7v/yjsaAlmMplEZ
9BnQwue4HjpixX2g54ii4k8rUpsVTOrJ17oPO2lrhtucxpAOgY9G4+lBzNsZ5qBb
Bp4b1d2IfC8xK8ZmBUICwBGen6ol9dS56LC92MaJCXew8iffvnfzl4IMFCJO2TJR
Wttj3y4Q0csUL/5sGl/bEQu5FP2y55E5hEfTos1KoUZAUTgW5cgDyiAhmIrVwwO4
sfrmCwTUuJKPOCBm4m3DbdAYzCzmPSfnR//nPlvdxzEE4xkV+iPOTGoBSDuhmTVc
tCbuKZjKDgc373ieOdeco+vXJA2FnZQ16MHXpvkfCY+GNzAaXmjqu/eh56OZ13uM
22XzRKtnevEYvUxMLqsMSs2ObsMzuZ7nav0sbqBOAn43XEocLoBehLF/ZMaWtmh+
yuPjijmjbIP2D2pdjJrTmtYx3pz5ZZBE3xFk+cTJf8iRDIto2M/9lDkCUkDv1+8s
ZH0O2MofTBWMUGbON3uhk1DapIuDW10Mm054faodMIRNqAT/+FBlHKkQRAw4jzK9
LHpsFvJEhOVIxVVb1x/kuboM8tUBYz+1j6+71j+mkSYs+26lqzx7PIXiWjK8LBkS
9hXfj+z6Og2n8WixzGwswqm1b0PhBFEeHF1ddHqlz0nUsFnrogaQiOl/kfDWkOjI
4EPqVo2hyVJ3q7kKA/hhlKnbVDlHi1Wy+wqqZu4Z8cQxWic9sebKoVYuC1gsb3BG
0+kyYVVGShEuaRDRgdqrdbdrfW7lEGfDloul+I3sDdJJUE7RS0USxnYSkrNlwX2z
+xBhcKmyBdE999dS6HHE6r1BNLRv2SUquP5rjv3SK2dCiWdkaRhI0JMC2oO+JR1L
aLUwUUshHkFBIQAsTjkMsn4PMuRByXhHPNIhhmLGHZC/+lG/fP7VC14mK40TMPtA
2XBCl0WgAsqjkQCSxDSLrxgUySNMcUY6uuyTNR2CzveL2ddT96FKNXtF6ON01/As
Jheivcvnx/6/JTNgUpw6A+zhUiAOXAcREPbLeaHn0nbbYRcGa5Q8l4ErrvtQEX6A
fThmsDuCGDNLNhxT/LyADJFVltPRFh0GGwGIj9lLMCp2wZcpyfeLNccMlCX3xFSD
JLJ+8xA1I7EssL2iRjZtKLn68KYpO0Ms1/7rsXFIvVzUMXNWZcdQNLWIR2eWfIeN
SuqLi3DHkVTmhEffXKzXzShvRmEkMDvnGRU1fftInTFj841EM2hGuS1CvK0Bh09I
7sEdUZG7BR1yFrI8nq7vg61bERf3eI9F5FOVEvRNRPkwQENSSpFi+oFWubRSY1U4
naCnCgAhaYcqfZivoxGMx6rUmyVS/lijqFN2HuuXXQ71GZ+zUytjLInsFdrjFD0v
97WyyBPJ9B9BqTISAMFvzf/C2caRNwps/R/dwWTEObFrxByN6JWIKCGgkO1ZK0im
0Ylg6ah3bEE1VzNC38TVr97KxK/CyYQqJwtjuIqbEVebwASueGR74zork3ehwOtY
NFe2maxXkyKwEsHg6QF8ug63wCxH9nC34HfAmTscdG9f5txuvzDPqROom/4K59F5
1Q9E3F8S8Fe2jIY+RYTx/yEHR4Rrf+ynSitfSupqv+t9vEq2W9KQGsDsy0jUImyE
hws1FQdyUyn0LaORWSFcf87iDyFRnuYSMX/vXeka+pk5VEwjdDaFaIDP66Q+VzVX
iyw3maLhPjoOzzvPJV+OHMQK8OS7dglkaNYIc1ycuRj0WMinxvr3qn3CjwQc7KwW
5/C7GN1KsaTz5ILl0MereONio4YS0K6z02MAbZPP0zbY+U3G+EpCL1U7d33CtsPX
Jw29MBM74v0bk4dmBiomf6r1QVJnRua4XtDsJkCsRb0vpuUP9QjH6sAc4czo1OR0
eFyqV5DX5vyMl9LwKOOwj5eTyZM0bPC4d7zCwsvdFm1YfUCcy28xGCUqly5ZQrNe
ENvi5S3ChNgwBqptlL1UNgqmPJ2Uo5Ldrh1dFu+8MUJTDS4YWmG1UXdnI8jmLfWZ
ZnFi+aWVL5W68Buz9Kfe26HG4nvcl63cfg0rzL3ecO32hLvwLLA9y1exb/9gDREc
FZCW5vL//xLTZMq6tf5wlm9duwwm5r0BN6TAYhSkV320d6HaYTke/M78IhVwnvWD
hu5KtyjvoTiEG2OxIeH3CQV+EHxRw97dYq8k25T2OKClaXoM/GzjNWxH56cR0ySd
yjcPNrghWqyO+U0j3yINhqatIwUvSOON1+6aemUvITli3gnh/gGKGL4puqInng4x
1X34yhrAqDnZVwWyrKILeANxNjWwwt9yW+PlpJ5FsTt9cuIzG8fiqkHAjtSaJZmF
2vrPhBf3uH8+jM2GiuMgG7RVQ4Wj4eMp7cciWP/CLwfrOWV/xJbiBpTAwEPnwM/i
fnCClJcDGeAXa2+dOwgmSesCytWv+NitCCUh7g3T3LZ0IB9XLJAhKYNh4pksw2DV
TIE023SzpoDDHl2E0vV2UFSt4g5Uj5a+lSCjkHYI/XRgYh6gLCr/74Lj9R+b+/Oe
Rcnn10R4VNvfaN71Qo5lJs07Br4lDe0RQfvh9z249gj3OfN8Emqks0yQw+Q7v8Zx
Y5ixgsitcsgfyVc7+2pWZRSlhL5Jf6PtsyoitUHt18nR/kLwG2YWnod+LEzCLeGW
Y8bhjXW4jlbuCHwBJIYM8CVOrdcqP4wxkyOH7CW4Sy7NCikybICyj1d330ZVRk9o
jY7jsp6tXggcge+yeMNsr3oK9TfevdqDOLj1rD+BUeg/MV/jH7xKV1sDPS52ENRI
frVNOKL6n8XHwslyBw/KNcCoV8Bsf2/tofUpG+nmYMHyrEc9JtHKZP7znFda0iCc
epbkhhNOSDRlsDHTcgsmY71xsjfMCLlNs+HKSIEga4KZjESPE+5tbFQOmVHWLn6I
HW/TuRsXAPqssDDfEB0SWN9n+mqAOeKBE18Qm6cpKJXbxvAcNCuEW8naB6I5j6hq
zEdgNIaELqBIph2F0SmfG6pGE+CbnQdIiP+tZSkSUfSbNuhhpj+N4Am82AoEnAfW
HrGKSxI3YYcm8EG05UCbB9vBZQZ+gji+sR5fNgfiDcOzstY8YVnBG9uMcw4q32Re
aRxthhOYKY/pbzMxJYRYkxz7dcWxxOuvCBjHZ6v1+1B8ew8s7h2U0gj+ijHRKofi
maqrGtYStzG6fGwMXdoL8iZ4otfirmAGILlCPbKms7KKU2l4PcBopVyzgC7n/W1O
CbtZ8/k4sqSeBQAWsqtzKSRn6PNbW64QaVm5AJTmSFp7PVFjHchLhHU/KGfp3lCE
tplFdB9fr0mKI+qn5hCNaFcTTYk8lOOxkzQnOJNjF23h0OhFpcgy580BdlFTryuq
SAGkVA58/EoLUc7jwtKxVuiRRksdjkURbUVxr0RElwGPqA4tNYT3XEwG2YnLPkBY
ofhh+i2oap53QT/7wcHvQ+jwxgIl4tyzwgA9dR2X+uWCYcP3UHbToV1R/qYpIXwr
1Sf7lL8SpbZYtg7YmNue8S02cHy60Bb3c1HYx2uvPS5Ce1q1JksXHRG9NpDOhI/O
xI8s0ZiUypvGgo5wyIrPLPI5ri/DqN6ocxAb2yR/BjkmrgDfrJ1lMiMVdHiYiwdJ
3yBOMZHDmSHQmjKBJg0HnsFmkhf+ceJ9tuMSAfoacKqJI88RzbioEH05yoWPqSEq
CsMEQMWg5u2yYIPnnBqTb6GEYsu1d8n7JYONRd7n7XZS7yseUAF+Tkbo9Ddjxdwb
X4l93EpP9oYY0YaOryHRORdaI+yJl5hT7LkJHOvvNut4D7J+3gTWOgAwaAlzX+wQ
ZquhubPTckaBuFVeB6aR86tNiMSzb+P3RxQce35y+tdzNjOvuoxLWJv1UJBFJ9/I
fX7sHj0czCSqwSZxtwDLgw52NT/4oe55sUYv2Y8nz5fVVhQyH+45DAzcTgFORtuB
j1emrGusDrPMFEh3g4cebXK2ip9bWKZaiymq6JX3qA3SPThnYn43NTN9Hy23kZ3k
SqOFSvsb/W2AB9arMwgsM2fL+Q8y/frWq91jjs5IDdThglYLvJOgHzhXa0dOtwHA
Rq/tSgSRYJ38B8SrwfLOq5/7z8vc8JuTThDx25NNvADfn+O2mCPCLEKcsMTjC0RL
+shrdGe1hyPJl/pA0F653vPUIiATH3dJuBomwTEBzn/0Fu1+F4GtCQeENXf/HtiK
T+ZDrNVQJzMI1Mmj7rRUI1xB0QMOBtKa6X0NW/yIGnhEyNTa4FzSc52mO1hSkjgP
eXUI79Yryx9R9Vbj75HdYKEtdS51aSIf+JTsRcMDIhUPRs5XGLlGmT8zfMLuVrWc
lgaQ5LRhDPARZKulvdT2k3Y6ul3NB3AAoLSPBOOOsCw3OX4xszVqICXpt3NJxFyW
odpKiK42ZYSYsba7jL8Smdz2CeQ0LxGgBeb8pV7Vawwxq3yKYTbp/7kXNqU7nJvH
n7OmdUKz5NcizIpdhMFheLDBhvf37w/tJ3p25QQ9vzeDkoCskUed+L1nUdcC2VXE
qoSOtOHEdxm1cE40q5DwyLTPXGTLppeII8Wz8+qg0Jrl2qJ39ndM3MRcE1m08t5Z
mnlLucny5o0g5o3UMfwsE8VTJGkK7BZ0CDL542yLSIRMWI+i6pzov0TmDeIRDL22
zROFF5Oilxt9GNZLZ24ezywWiXiKJ+EgShQjog5vhvErpwayST4P8E4lN8A5bWIg
bbmYa75cxIYiUdrwrQwGvvCZpj69Nu+hNTpbpBNhuKnSG7yONNbF3rfweDRs3/9A
xEl+6ug3pcYSltWjMzq9EodUzD13zIL7oVi69zyBNk0Hq8DAWY1cqDF4rIom6lXM
PbzTWziItKYLVIWtsaqu76wdtP8w/tt1oYCJIONrKAVNH4K2BuXx495oAat4k311
lELxtfOqxEs2WKXSFGCFAh3fnxs6HjDq4ygbibwxJt69JH2As3D8Sp5+wpX+uYvu
snd2GQi44TVAsuj1daqeJGlMoKLFjpyGqod2w1XUrGmKTo9Yc07G6fioQtTKQNEv
Sy5MbdWZOCkJk3/eG3DLSGLLG0Gowz2s7gEe3HQEcFXamdnnRILUVedeQL0QA7l7
6t4z3UGkIB5bRvQk5MLH0n7VQVktDQ1vSA+XsZcXXVAp8PoI4KtUn2uitYUo1iA0
Z7fIuRbPVIYrT8AE0pp6rlccu3GMq1fXJTMOPJF2B4/arICAx6IvSLOlwYY3qZvn
U3JyR/XWQ8sZNxEXGD9xHXRyLVhmr1nQ8+7rBsRzP7gWQ7kk1cjKwW+au3eoBX0+
IzsYgn02iJWVd3tdCtoDqk2+PJmB6sxl3wr3IN2nOgA3YS1r8SffGimViKla9ED2
yLbH31acpSP4zuoDF//3BQDf0t0lOsVi2oRp2n+x4WspIpSk1V2QQH7l649efbxM
Ao7QzuLstVP5e60EB3Q2WB4apSFRChLEZup0qrW6oD7K/dcodSwoMA6gqV6lhpu0
9KsJGuaH4BCeZPr2aG/w2xbxnVXYcRB6z2GWBLu6yb1jv2HARiyPjXhN5Ybtg8YT
eZfAahO8kCm1G1SL7kATcxsfSNAQReCag8mhRTkZwMR+w55V001ZurwS90Wjl9co
/yeMT7njY/MIXcdDIl26WXWfJPA/jwgDWYIeWcwHKaE2k1b+Iu4rt6QcBEavAQga
L4dOqE9M1bEED9mlMUnCx220TCWHgDfJVMLL3T1R4NlJzmz9TicHfNzvOFNr4jIx
syFe5dWC5CWNDhegqh2TsUamevvZcBlgg6QuXi9iEZ6YlXAXTh+TUuSopFHaS+vf
06ueWAqIMqyZKwI5bknVMWfkO7o95SWVKt/aNe5sEP9Htllfg73HR7395ajmiSGd
zdlwJr9F5kBtK7rLIrFCrCyP0+1/lo7G/xoC9Y8ewFmW+0yQaTw0gdjV72yLPUvC
Z5FG1jzBHKrS11ZSTMLrIuWA6XoSvrYyPgU4R0LR9BAqIk98Nf6R88aIncBDvJHC
bmQpLKyK2vF5PGtoaB9oObfDMSkZrCfQkpIIoYzbkZvm5OkoD842V0BOAj91uG/R
jOOOhnUQS8hLIn//eQoCuaPOHV0RZuxpxlAbPZPyWxNoMEJAtLWEzMwlcCMGWxd8
fuX+OrWk1iCXQUub17kuE3mel4ucSRMKCYYdXDRswg1w0gpQ887oNKmNh9Vykfng
AxKeq46rhFjCW0Zhw1yJYHYqPIZAa1m5Jaq90ILWbQ8g94Fg0YsZdnzOkumCt8C/
MZMH1MOVadPY3GJQHImFAcaJ5cT0vmolErkG0jRXh6CNWhJwpyKQ/gJhpMv1L6uQ
/PU85cInszBZcJZhfL7q2RJO12B7XwsjZR2vb2fSyNGEUFpU1tbWK9AtOYk/2yEo
YZoy/Bvr6eZogMDWAae+R05vM9u4JDLc1wajP1q3pLNpfC9TZZ6eUC5y6t2EloyW
afnLVonverpgyEKpmBaW2oCI0jeC533kLEh8P5HrsSPjWAcomxYFwb7tAz3MtSUt
LTcO/y7J7ODXZeXSbvc/lUp1MQpgGxlA1w2ITbKGhNXpBSRuJLyrxQ+s/TB/NVZE
XpLTaWYHdHxg+Pskt2BU0k0FaAAtg5Pi7GTL2SXYgw4CIkdZZUNA/dqlFKHS3Ziv
mcgGRYbEIINHCpSFmmIOuFrgXci5DR4Z3LzoD9vK3pgxYKtaxPY/oeRrfxFrtPMe
G9FHYuOVxQHP5DFQQc78en5Bg8uto1Svt/qzB6je3l1kMgb+suhcMAp3IQcIm/cu
UhF3tN5u2f/EGS4xZhxwnvtD3k/6pc4FIi+7dV4u2i4nHYhWWFDhC5YVQ+Q/WGn7
q+TK7ZbcDTzmvoCYBoil/hf4o3XgfrmpcKlyTsQzedWsgrMl94VomRQLqOJ2sfNb
KlGZTeJgtwj8MOwdqgmTsiYFZ+onAUu7l/BOG1T8NcGrpS64haxGDIJ8w3aMBT9g
i/dUzD8wu8KRyzYfAe5qy+6elFqEce9wKgxCjYltQ7+sBjKytok7swZlGv5F5nZB
kZ/NYrYe1ph+stvZ3vlIQF/k30DWtGMFgQGOIfvk+TXtH71JY/6oxa+fx8bBNjr3
aZxilCwr6HLmbfnv40tIYyCZGEujQ8V3erRV6/rSYYK+gh1ZCaLVRBjWKUs6XUhK
2BEFJxXeYTRXqZgoQlxNBOGSFm+cwUOr/xm6HKUMAEIz2zG3cICFC4Tp85RPilJi
dNEE5rvLHxdJnMV/m2oziOTVO1KKQ5nNttAqC9h16ZRqVPo3GVK2JEqw1wd+G1IE
Es/DlyH5gg/5yB6CZm2jpB21YkvJRhxH1IkRbwnFtieZsfsIEaShQGQlV/7+tufn
VokKttudBNh9GXYlFWennaSMfetDH01eqo5AkTXyCQUs/DRmuoizQmTSQ6JEnQs5
FcXc4L7lRfeyz1dXDcicBT0r8W+W3lZi/TmfC9Khckdosa6gMCunDYPw5VXtwWpc
HYpYuTuAi7XZ3IHYMzIVhSPRv8JY6PWg8Vjvnt/h54kJfxr1RdpUDmzqiaw+onid
A2lermLXUFZlrSB+dkN61Jp+96TQcc/qiNJJz5OlGKcN5zPdaXHP+JqCeVX5AnxY
z6YCTsBw0Qi2q+rDXWEtXGI4BYTBIldupTzhZYjp2wcSG2rG1tGtku5SkMFO2jVv
d3qnbH4X8MEWZljNqeu7h6Zz9OSKazojyrdsMLZznaozSKMukcwAz7VLygzQYQR3
Q347KH3OS3ZeWlPovO+fQOtegN+ci4fHUQM6nlp8Q40pJv3C53YgSUzzG0fT3NTF
1BFu2HHiuvWToObv93Kic3quZDGemdZyQBJk/voYku1b3BFK5xDyinhSnt5RQG+1
x5Ko4Wz87rzyts4tpjRmfMDOt1CDl8NkUxCcD5IxI7ecHwHZNePifCZSN7jhU8Lh
3bCLrVnrU5h7Ib1l/a4Ug2xHAf3QOPKqlRnK8zzdJcp9sryezWPBaX+cGzVF3BbP
kvS4rGOCchjR9vLQCNGldjNScoIwC1hDx72CPabVEHRIDxzlYH/skNRm2/SeLir0
7GHWQaQbl95SbMMoVI6afe/CPdJLw6/00oqlbzJenKTYAipdTx4RAv9sGIALFsIb
gN1bve2u9lkU59ABMTjSlLwBy3sWHbIdvzJFz0n3vfYbHRaiFEvhKnP7qBlXPUKS
7nHqacn9tc9GJDb8oFYqfVtQeDdK8FREbJbt7iS3BR0ZC1/Kbb2K0Ei9GEQ1DG0S
4b0HHdQnRKDZteqvN+Hy0ZQq82+3IwqmTwiBfjraOZR+/P4Q8yj+NJiQumpRV+60
xY+BSEaX9PTWJ0P/9KY6nR6dQIkJDnwpknzL9nzFin0tkxWeqZ9OEHe8ohp6GKGO
LMkOcVfwliYiR/aMKvdMJ3p5cGtDyV8doXrrSPdLQOUWVTOQj9a0Vs+tZm+swmuD
zN9tCLyUBhb1GEt7XgVp1mSSZwLp/zPxz5u/EvbWHa2EvSiLG89o4HPymXu3lypZ
OGe6MQsEoQaBegTBzqJjlBuG1VutpUVHIJjnvZy++zt5JYEOY/59WTu3aHRROuFZ
yQTYzt7YjZg50R33+LEwIcy75rVRrmZY53R690Zvh5MiSUC03OGtJB7RT/j4Dbv2
c94VhTZNJBnvpti952tydXds20YmkrPxUIE4U0dPYrI82npDGE3P8wdc+535cSVj
mlxJefnM0sldFFLkXFNtO9ePhsq30c1TBVOcGkmPZ4bW71gZ+qMk4UanZ7HqZAdw
dGM59EYSmotDXo+Co4UiDqD6FpykziOPnNATB52JrpXo5CMRrsfLqaxuuojyNX0X
Dh0fhbNh0mGV6B2sjTGNR3gaJsRPFQyo5A7BllHuN+kTzpD3lnGW5Ra/v+ofCzRv
w1Z++T5gn17nUFk9CC7vQ3kh0p7+WyWQeo4ZXnX+eNaw4TMdjusi4agsJa09ctHU
Dk92821LzBoqr8cQnA6ez+a3AmuTritSLK7nMJO/OJO5ZPkz9X8z8Pvcp6VqIZCz
ruIp4lXNkj+iKC5tUrZ6pSvC88UqZ1H+ej6gkFpjkEUfFbR36MAeATQ15W+g+zpv
N7Wm7iMy04APAPGUhsKRzcCZiNwhLq0BwIkpiaM+ME7YPL7sWAGl/wx27Fk8PvHG
y9NGOFfUMiPZvrvp6ozY1jNI6Hgen2P5u+98vv6z81VGrg3QwyykYFa/WT2/KqQo
CleGHHJPNeirLTf2IsSLsns+DeQ0W3OoYyqQAFR3S6XQU2KdST1eYxx9b4H129rL
OqHD/2raDiuV7RatN767YuXPxbeUJMQ0jH5p0ZwqiA31GqOaT9uts/ERDy0PUy32
mykjc+2mDz62cQx7pXol9GaYFExROHcPUMsLsANhPgb/xQX2L7F7gl3SH9XRlq0g
K8+VXC0qWYTRw8PI+fapnxdoL7UAB9V1Wy9m87ex4A1w3W1BIL25uSj2NpdOk5h/
MDYO56m1Nu+UhXHCFkWn4sJpUhkOTRZAKWEohJZNc7rxOHHG9VpH6di0naUZJ4r3
/2mLSJ2fi8RALQC0yJzGTDJ4SxKLp8PmSS/aVQxRsBCKEfa4jplUdV9Sq4WYLCHK
NilCIH+f2J59tczRVVd2X9gYy0A8uEDb5SkzfDet3nPmWOccofLP121FYuer5him
kw8nK2/1qmFLPblbgHTC24hQ6DKLYSfeyGii5IEU03OVHHftyz7ZyyVekEKG8jNu
UhJhj9P7Huzb63nInwSvvPYQeaO/a7tcZymQfiV1KFEv2m1TtLi9f+A2BvvZz4H4
vwlM0dOfzvB882r8Ly2aSmlI1CnzsPfBngNbAAi3JLF2k+9g5uw2RZa4OkdkLBcS
RifLtU5U0ibZAbZNI+OxHS7Be0e364zMTzaEeLpsPBdl8Cg6O/ugWvj72W15ZBdd
HvMcj3bp1qLdp4QYBrJlJNxihTaH7SGyL3/TYlUDayEUg+zXDpQOWkfuxIUUCa5D
g9aHbclWueJYEAIcCfdM6GAmgNvHxQ2plgbEq2Khb2FnRr2Z+9jHIek+Ld6v5p5w
gPYr7Vz9WgC209skeHgGjhCAIsSkG4kTq2tjvxw7tO4c4jkX4ZvBVYWUFE5qzHFj
66tocU5MK9ymbI95CvUGEyDAjj7M1hyYvhHjvJF7JUJzNq/DEzYUjIV5BgDnEsnB
TvZQ2/vpuUucnBuyROdT/H1FOJHXDcYj4dywVCvbXSiXThSL6bg06EyWIuloMD4C
6WwRTIJh7Vm3GWNdgUyKO25J7xHGF26pN7NKNBNa1wY91q77ryqWj8iVdbpft+nF
+vsZzBKbzuX4zE1rz69oY4huH5IBQdk1pjM4QKCDqj8Nu6XsdncKkjPZ0VQDIYif
ZYSaai3s4bKjDbWdbyMb7Jci4S+GJTI5TeVYsoi7IXkGE4ejtecqpr4tMf1MsN+B
Rs5pFV9zbDiSStOOYD6YPHMEW5a8btuZDpmEu2C/9EGiMVxZbkeS89DmiSD0nKxz
vAPTkiapZ88zXYYRD/+MeX8V8hKVY0mP0Xpdbb1W0LaHrXGrdCgheNmBryYx/cFD
GN28lgBBbclQBobtjdYzw5rCTfKGZL3Ztj34I3kzHw4KNo4/uicUmoOA+dmHJC7V
a4i52FjJwNYjJZyB/Xn3we4QXviEGMQsJPzV+jHl1m12+lFEvs4oAQFwBFIOBfXr
9uX3NXl4sPGin1WPJbEbxygecUJWxjKdtx+GqZ07bDq3qnB+m0lQfp3l6plOgyKa
DN7hrxICosXFQbZxfR2oEeq22TN7dx6XrmW7oYBVkY5n5a1J7caUGyM5tSb2+jj8
1utxWhP1Tad90Sf5aI+XGBa4nIcxccqNNzDixmvMX1O6TIqHDF4WSVy83hqIqf3Y
1W6zIQSterM7+xri9SJyiGhI94h0VOYwIXsxVg0XqqWAQxYtbNflWJdDI9koZFU6
qVJT/UuIApc2JW5cXZntzoKhVdhMI9P8W6my2tSnG978x0YaRAKrLoCcckcExu7k
DIZzfpN9fiCF5V4mOvAiumKHDgxI0A34crg6c8Ez+aHOnKeVd3mn85/5kGYu7Ukx
btxpSiMwFkzxM1MRpbjU5wyvkrTGnj+VE4ZG7DW21I0duegzo40imV4RO+NlzP2F
0iBLdRjGFEeh+z06WZgZlWzv6ufPgv1+CRrwvjBW7+flAs2igEUFrESBzl908aEf
H4wj85M17Z2xFLQwTu+dNCb11WkizKf7e/g7jVR8fqggRz9FRhoQ2zCRI7ELL8ap
babnJ7w0U1pSFWaYYJXbpjACjHhchIaMRLXTsWIKwpKfMK5aqQSN5cAug6Lm1WbQ
0IrgW0ZqqB9kNfCfJdAklBKeTaNi/3vj92yyLzIzX/a9qJC7+zblG6ldPOCUWLf1
57KvgrA3f6nLklCcwsGkrd/5PYjwHi+tTjYdclUjg4jMYu452iNEH8wj0IrHZbtc
WWjcIKX8gnH/MqALLPBEO/LLMNdlaldS5K8FPNl19NYa+u7xLwZFsccCZgRZWCun
I98EOFrodDqUYRUKIude43+LOIQlpOCSo/1Ybw3Nz9fsVGVQROTNSBnOCYLEAsNx
8UdtOBFGL4r34DJ36WtEy26wEx2abOY4OGxFj4r6YGZ4wxuGDcot4r7vsfR3wdKa
XpBLJNiZ0d2HzqY5z9knXWnJui3Pt7CyZU1TZ4Zr96Y03Jn4riPNzzKVXSgAcR6X
BWSCH0U+5BV3hxb2EGaLWqxOeorChPvx29JN5hTQovMcfoGaT2bg+6xXjAnI3vPy
mhvv6+qyqouGC1Pn+i4lg8KMoA1q+vzJJBedC+IkDeGR/qJS9v8qL75DrWGtum/b
FV9KQZ2UoKjmKhTnXewCn4LJE/I3V7dv7nhQUdTxxwoc5rmTsQM/ht61yfKR1gjE
HHlOiUTWx159JSs4wBfQ92qNmJOtROftYn+Iv56sNFJHPoMdl+rSuhZZOYLX/qp+
sDx1JZT8OLC9eGFHGjUoUQ9/sGbaThxdOv4v91NLKfbP+Xu08PaFTOu7sRmA20XB
oDxkhQme80NruzdXhGnUM6iZMXlh5hsEh13iL7+iWRFP5zJ5scULLyB6rxnRftIy
GUcZZzuMYRZD3V2v7y9LcposFbRUVkn0W5ZZvi6cJOAixjYLhpknBcYNwXryaXPI
xDhiJpiZvvNdV6v7gB15GA1OTUuqeNkZHQDTrI6spOGVJhlo2jksnkur1V6XVEd8
upXMzifT0OF1VeSJUiilK/yyvksuaOxw1klJCxCQ0ierP0vF7rL8gsd3a3BCFeo5
2l7rtIqH2LYhHfTHNemBHf+eJSnFW/rAM8tlOiBijeAMuG8iYIQ4qVbCyb18cjWT
MIC2R538dsAmfDq2FPzA2r3CHujSxGUPGA5LFR4VoQAHzrnYFJ1jZG3l5lIEYj7g
iWJZYerW4eGkSQbGIst/BW3b1R1mqR92A6CMiqW60jUBIltlg8ODZMsHmXwF+CzY
vOjAIQNJGBRTIE9AvvIM4Tw3zhptV40hr7FNS+q+Zwh1nKjlaQbMSiO1SOZdJzAU
7qb/aHPKkFd5LBHeuTr5XnTxDySM1fU66AEGKWfpB2YaXFDYL1i/IkwlIgTnH40P
myUzZ1Bca82HSyeLYL5MkZ2BdkT+sYT4IOdyuIcOilbmspwTi8Xs9trUfKryrosb
Aiw8TVOGOgGymFL9hMUrItqaDBkZG4+fV+WwDcVBqtM4n3i2v/aMS5AHde7WfRai
nH0r++vsrtH+H28DAA4//KAf1aza6w7nZSkfF9tdUJyu1u+zEtkJCY2ByYz575RS
iDBDYfcEyoALVpbmcAAAR0Z6OnemYCygsucZdSnhEu0gLrm1fgJcvqNsGDXNlwNb
xuiDerm/dILAGs7qdRl1E7bihN9NVvWn4P5mK4sjNnYeJbIK93VJyphY4x5bjves
UKhoMPR8t5M4EYNPPpCuaJO6/jNtPNBsI0oFxXVG5d00JHrgoVH24sTBBdaqSqOU
1gq8k70gbI0vbQh47Mj9j8Q21KUG1v1t1kAgU9gThof/0bCXxJi+LNhB67XuyPwE
hbSBKf+8c1YmD1AwmIGcMiP5jF88HI1eN21FVq3jRNBL6iepizbJ+VYII6GgHfLw
tviJ/yehagBXJIGhfxOUvyCBauvE8NEilx+naZQVsUhJU/aVzGJIC/iVZregqA0f
u56jue9mpMspJvkorSp6VeYlK0I+fMFnR0/GkVlTo7i6nAiHmscv4p3jfSWCamTj
gX/OJXuYgv59vmzMseOhtR6FGR3N9Em/xBiTLFmdObV9w+SXo1GnkQN2NkNpeRSu
7ovg22N1IXm2izqGzigBGO4Sy90JH/40okcik1lJOaoL2hvYlDUASmWN+g+m85i1
6a0E1LVHzvYI9MNj1wX5D4MzhKACcaP0i4WrNT7KQMMqO8Eq8DcNeXehPiaYY5TL
1eqQua88NckjN4PMXdLoL2unHhXXhikW9v2Zzr9Jn0Cb683CyOvod8wgZWVZOKcz
u3VC2tkvdsmJqXoLIteB2ygTrGEBoee1jofYtPiTglaDORRdwEz9N8Y8MgWIScD0
AXBL4U6MQrvKf5At5Mirm1EgcdWIE3A8JdxUCwVkyxtFvxenIkTi5GP0p7Jh3foz
DbUlS+LEw76mUQR8Q+m9GQoB7D/E0Cu+e9JmD8jErZGrUKGDmd35d5QNui3oIc4g
ZyZcQPN20XixRAwyFhzAEk7qWhW0E8vs+tlrgEL4gaRFsT9vns8sHJYUp4gwow/W
/Ygc2WXrH+syW+gF3BdzLoRlcAol+Ss5J471n36XDzpMQKt8Plw7bQHUfiavig5z
8JqS0kLpxfyPHKEwRYQLgJMtiytVXEYNL5ROYLQ+QfLBBPf3qdHSZ0hM37oz60Z1
ER7HYmPjlM0nvO+MnaijVl+AASFUO/Mrms36XXtWLuQRXFDVHdzCcJuuKUgzKyY7
AwXCpyKGlxQQbP+r2GgLzIA2lGbJ023goQRM9uATZbCoMxJs15Epm6tpHyuFSko+
LzIfZ1I/RbR0fPbUCPrrOqq4pgFyijRAF4ECCVfjftUZVc6I3o8W2QTlA/IXNViW
yxIUAcoj9aeSYxqmxil8ADv6baEHGuM0neDbDRcpYzCgKmU5Jnirz1ubNRnDWR1D
s5XCbxd9fFn4bZZHDP72LnLhLfJlcJf8ajy4tO8IRzEi/vvlO53sWZn0ui3E3DUs
qklcNDB41TZf3ykRO+I0/2mFP6CTSsO1wVo8OJqjD5YssJ4S9EjI+G9xC9XOMnYe
piOpJYr1FjFqHATZh8r8aFTPNMBjyKDSFuGZkbBSISXUucC6EzPMlPaYFuZrR6xL
l1sTF2hv0BT5LBZlOBZAROqXMytN1X3250uhrWa/cicgAJkjxwzZc3K0hVQhb9A+
3y4ZRjrvk5bZ2NQ2SLUuG6XbCSDa1IxNuYSDFHwMLRlzaAL5ytNAnvw2QTjZhslz
b9QI21AkBvKHdUl+PVaztboxHtUmNSJeVn7p9FDO465jdD5iZ5eud2ha+DWjQsTQ
GP0k8QEZUZUx4cNsdpXiCwq1mlcJ/Sa/GUtg32gbTc3MIHcX8iUfR+w5+iEk9Y25
AE7cJxVZxG8z/vmRZjVmabgZGGFfcnPpZrpIqa9Nkq6rGpK7pDPUXIm0dpeCIUOG
fqd4bF0HYu3lQDF7YE7OLFWJbr7d39ve0ZB76EQbKC1QiskWFxAxKveNjYV4ulll
U+hGJn43JhaNh8rAc1qXnY0SkfoUOo9uwwWCZHVXWHbjpTySDYy2VHsik5QK+1hH
zgHd212ZjLEN31yNRp85GInvtR4Sxp/TlRdNajZIClzAQOEObFEl6pCIRFxrG/z8
IHyS+8sqcAOr/tgGb5+MckgWaz31yM6B8/8r0vgCUQGPiGcO+YM1xLXm8D8tsxsl
JatkFqmOa0P09Zr6cjyraxeEak5TbsbV/tQa9pm0UyVci/FWUdr4jYkFlnURUmA8
OXgoWT1nKZEOwX6NDGqiGIr3WjxAlfy6w4JC4Gd+iwp9/uz7u3re2v/mZMH4TK0O
HXxFDLrJ24DM44i4zQFNt4VbDosg/RnfBJmOsG1Nc6tXn/n2dK3dPwfRaG23LVW8
WX5bWBD7PgcH6M4A3R7PlBpNNi6mYIrro7rUQ7FVsuoP/sHaet+yjOlrYoIZR7+A
yALm2X9zN8AmUbc7crBLvSFDJxyIOapJ/KWEfIkeMOtKveKKjuLLzF1GccoKQBT3
F5/4XH+xRa/h7I0Sf2/UgxX+AurAJx9BU7zMppq54m+o2CSV/eQWrxVF6XHzl/SQ
Pyw21ep0ih5DdFPo0R0kH+RH00MoJD/0GuClstDPsvGR+oQOOIu76blSkkb9bMwc
fM7syrrBTC6DRFQUYGhrb2zbXwVS0klZSGvEJIuG/y0CJUcJU/Iu2LYYu6eWPf5k
Vy9bYnootrheBBTn/2qK3EaLKAtlFgZkVLPO265MjEokMxFNs+Ko8zAWhJUVCNyP
HnrABJ+XltlRzmVN3z951LCulUqd1NMouJqQZNNv63FwOjKpLAQKrengNqS7W0GF
URF84kqlxLuTotsHCuN4zwGMm+1W0M2z365QM4AD6mZ65sV/rcPSwl9eJSIu6oK0
DVIsXpheOJDfn2E0Vr4anAWtQT2h4TOtIdLNO/BCU8OgDVRH1pdMbTaPUYkoAn1E
Ghgn/St3BmkBtofzkrmd3yhS/aU+30bAJK3LKoGYb8ckqhp07/gubBUqfaBCf2Ys
Qhi24V4SKoI6G/PgtWhrcOuA1M+dHM7aBEsRhNHsUrL+eLtzxLLc4gmMjLL0P8Qc
fY3zAiRLnn7JuQLIGOTt+b6mOxKx9ZtccB7IFuAgAVwE3mGQUJGkf+CF5HTu4dV5
L4ok8K8604XxMb6mvFn0Vy8Lfh45ZeGOq1rvhhsoAWhiL8Mf0p8SM0tBkEdbPSAb
lCepmu5MSGjh3Iwbd2sy1oPl/yw17A/KKvzx3EwWZ5sxRQ8hwJlHmaAJ00kBEj/Y
zsISG/1MdUlCD3Hwp3f1ACie65GOQZ6cQvSyWjGnnk0YIavwBHo9uDRbmphwMHun
pqpYb3OZr4ZC2G6z7Fjv+xeeki+jvbDtoaAb+/VSL6PMvt5tD0xVrCLSaDt/whWz
tfVjl9rxaBturpD9rcHJc+evglu53yXvcu/LDWG1BmNNO1fj5Q7hkDdpc8FzTgT4
jJ8Cu8eJ/KEN64HAG9XUKE9HElAmv+spF0X+PsO44Rk2MX871YhoeJZWfL4CnYI0
tNuhCAyNxZZ26YX/h/JO49HKy4Gr6nwscN04qwXKGSoHfxPr9wXNbE+ZYwZOnS0C
pXNKhe7cbELXBFsalUdCnRhwn/OltPLMBlpQLJoRXz0kp0ezeLgtO3KCtL98emGH
A376aFAcXAPxOovukZnU8Qrp81I58Ss8CrkcCrGOyQmPxdPEIaUCnCm4SgXe9m/5
BpVO85v0MC14LWE8a7cwZuOZXWt7mjL/xrZlpGhRLjN2jMwM0KTTu+F04kWzbbMe
dhLVS0rxHoOQe63AaXh0oY7naKFPm7m2ZdxWKd/VRyuxh3ReD/SEAV980csLq83A
ZxDHZPMF57Q1IsANfuE0nDShAhZGeXbNeyQDzQUuOIGGOkuT8svfAlRaRchc0AHj
7rpTU/jAc4GO8PlPr/Hbete2EcQgQIKJ8Jc4RWeKyO0GqR9kkLUSO2QrkIKSR8IY
YF5BO2NQ/fQmg0SXjm4p/OYJWF9H/jDHMW473FxX7aS5pXSV9JzqL00J4UzvQHul
Nx1WZcUnjWXxfQQ7rGAjxzOvu/wjJ9DEU3/3d/XnPs9woLRMUbz3GXXj77WY1Vqk
kz4EYKt2q/5vMOqU2Cd1Yi8RWq//7r9a0SX1ORaLOtc5Uy3AO8NLqOZvq+/O12jc
iBZ4Dg/ladTBSsHmfUBr8fD9VM5ANb7uhaQ05WqFNe5ABC+scekeI01XyLsztyHR
Z3scJcnXKVrNx0NoOJRnX6o7Fz7RNE6VdWCw2bVuWLyONCsfMb6EJiIIN2yUknos
sX0G61KAwZRAd+obh0p5cvIgAjT14AUF6DOvcF0chtAIHlUndO4BWaTv6qpadLom
mrUr7mH8JeYj3/VfCkioswEsGsdJdyoIN4sqO3TY6pIookEDgQLqElM0l9y8YTMC
x0rhByum/qrdqUjNVwufuDgftjdVcH6eG/TLU54iBgwMBfIfv/Ei+cY5E+QEN9J5
88UnBsxqxuvVLzMTHR3xg5Ydwmg/3ffk65pDRMvQ3sA1WbI8R/IrGdNa+s9I9z7L
8D28miCO8YrabaIFC8On8c28ByT6muIEJAtlX+pPpOP+KZnppU6r4oziWtbh1lle
opAfEqfkmFhSDh558/nug/pyO8TdfUTff4ow5XyyVtBjcq5mJ7ER0rFbRZrXs45o
YuXSwPRYkMZbDOzJ4BA6g5tvN8dPql3doAHSzs7VbYGosCGmswRjqQBTj9Idgc47
oFbgRBwOBSZ1qeFMhVXpam5zpP2qUCRPorVN6BMk53nBB7YkUnUgZRBLfnO2FzxS
ucRtwEUaij5WFG/YY5Wqw3ko7JeYrVBNt2YXizex5cdYDtjw4HDfywD1O768uIFy
2bNCqMIHpIn3BNzhzKLKOXXrtKHqVmPTpGhaAHndTUBs7rwygR+LOFKeXY0bGvMp
Sd6YjwFjoPK0RAOWxOZczPEzug99c3qmUdusbOxcTXRY++G7TvKGjRKhQ2LBbf6Y
8vV0f3mj6zRWKYVHUIn4QlyYebgsojzZ1OQ43wiLmtSo7Tbj5n2epJMffgUH637b
VCx10PPaNrVZ0rBRGc08buIXz4oG21YLtgSbbIzlCmSzLyakmF+MBhsBgxx1ooay
wJcCck6eK8cHiEuxTKo9IcDfDw59Ih5HcHB1FjFRoAOJ/WZ2khbJSrEGCJIcr0Pu
Y1ONCWpzHD0VoInZ3ncmCOOpC+5FZ/BJ6rTL9Cm1WyBgVnOdTmHTzDXzWf8uc3Bi
r7kOUyGfMklknK3PM9AbmfHx/Fx2ElpXYmEFsM1tTgIQUnZSomWJAT4NIfGn0ZKL
ipL5oisBfMng5cet0VUvDaCO6kR7+du2w39lQDzRbbZUp0FEgz1fEJdex3tepVWZ
ohruRSpTxfFzQGRIS8yi0eru+SARLpT7cMXryE29EzkYumDl683R4jBcwCAXohqR
Al7pblA429QdyvPt0qN+IAab3OdW/iufslLweLcAgsltZ4uoB4C9zVYD7gYyS+w6
0wjIGzLpRCr/p1QaN6DyKOvzUIoStZXEqbbRdTnBJ0E5MuTt/ENq/GA5+fXxFAvx
IiaxNt/+h0DmN5GfZtRw0l6FQg0UFbZispGBFDOcJM179nAPArTU60DsvgT0fxL0
IizwTT+KAAQvdKOR/d6Q3itCZ+NDDIyFaOQE38i1eleBcXlJi9narcGuCEQbV7JI
PHxcpMavGgrr4AhNnio9dELCHcwt43AAbMs8p1Bovv0qRMvG4Thj78BGZmqeJMBj
m0aniUyIZsL3tAJ5Eik9CRfxs7CDNkLb5ja7Pd2+ZrDNKWygwNS2Tr2RaCVgHymG
aBAEILbDio0Qh18IMccQKuXRdW3tB2Q3HYOC9MsiDU4gLMm7Ck4ZAz58HWGOYD2M
8bQsswCrMX7ixlvW3xTBJWNbhJlG6q+KFWpMCO8OWBCGdHGMak36FJs2hA0kbcvJ
GFbqdzehI21bDRIeW9ABskJmwCSNDTGzDyNkJrHnEU+Ro+vN4pPG69+cMEhTRqsR
cZLFfrTDOslErhSS8WUSZPKpId7xsgDjTg9c4Zw2jNsDDQo4AlmLeT5oE2Tc4NoS
rb1yxG/cRx81gdIvw/pz4Enf07H3fD25lakgSm/ETQScoDv+WVG7EYHWF8rUG4GA
E1v73YSmzLkJDOkf6z9yVNQ23vjx0oeSiQtlIYI91FP7+xyjShsTvYMuiBptgMoP
aJ06dLiRLy9atr1zYngMD/yadKsKRso+ReBJzZRSMm1qmRDJAuoW7aH8o/5kQwYI
yDxz0/KzD/rdqBmrkfCkLMw5kkQQt1ARJgwRtjzRx0gJjjnOMLAyBMYG5etJbgNO
8MOYQFFrOQpdA1t8CvBtxKs/+c02pu6ylg9MuafznObFjp93AzRZcnUKybF8o3du
+JnF/TPFSTkcwFauQvAmbrl+G24VCRV3hQBJWQSc6df67728N5XSUfEDcLKEDUw7
8hpTNzEpUPpFgz3w4TSEhDcCGYN7ZBeGrL3pYLXD6hmzZNX42s37dOTXdKnb1zzX
CtYEkmNVxeL5f+tXPFt3RZAAvqUq0zgxxWLHQqKQGw6KTl+L9gLdfCH5BTcQ/GbD
x7GA4w86BEkqRDaPVKtHAaJuZyuVkzNXdLnWJLgMg3SqhGhuU3kD3UM6fW3Kjub0
NDwUqU+GZQStSnyk2Bg3PcJRiyFTJjUE7ncoIJe7oa6yDVCXS/xxpupO7gGKdQwq
WwWxmpENHgzBVpKVGdOsV1BksJJ58ljPSXA5FU6l9ahRUW8R8VJDKurosMhckdpg
sPC5Ni0wkkNRxBOGUhyQ4M4aNlu5KfE+WwsZdXUcuBSqL83EwVVhMuJAGNvnLmnb
t/PW8Yuo6IBFiEs9qz9F6hB2uKENUJqWon6Qwi0ozesuU+VhbA0X2Mlt9DDniHVV
9hk6B/ScVlc2uGv2b/2Kqh8+8Z21YLNa3OBeFz8hRdsobnik15yq9JrHsH6qBpMG
7pocdptgl6neTZQ6WeWCdK/Zog2A0+YHDOjR4SGnMy2PTyu4QUoe356pKcX/gHf8
hMKotf3PajrZATD0ogEhfW1r5PU8gDix3b3cnn6aWwR963wEviS+UelOaslIq7/R
m4O3yOVujuaSPUWodiv+5z8qWExP7jXwQxGkSq++wFfvXN//tuTXPFYXoHhpYJGb
5bBs9OQK89cVkO5/Fc8/yExS+/WgpMp9ppvjC5ceHjjORlC+7HWI47TXehYE5ziw
fkIxDcwvb8XsYkUsB4HkTOydrADpLaVGdt0z47pkDYkd2smyCqAeSc6Krl8k0W6u
yLCOwSHcOguRNIA237l2a6BDq+YT9KhS1v3al35N2Z9KxRamoKCEut8eeASbBwWU
0E4RCeRHCfCVGlOGJcbz1jICqcOoYMNWOelaojPyLertsCLwSCcm9Oh9qG3Qtnkf
sVh58vwBxD7uE/Ygu6NCy8N31Magnwlrt9H7shQiHu+yxZFkZfuvaptqHWrm6wix
l4Oth/uJOQnVd2i7n5A4+WUJ9GatfLGywTkpLH8/FYOblXZkar6DU5J9vKH9JWoU
lFn98qkYOevaIz7/A9jFLrhhojV51NJGZj02XXf7O6yxftIWnG6usGh96hcwZAK4
b8bNk2IZKq3KhZ7Xy4FX7FOilKc/mWLNiciMRFbjalXd41B1GMTwuzEVVAMm4qqe
3kmVzdJQJffTXw92hRmTJYfwlI7BA+N+eZpdCeCPmQLH0ysxMC3OR6gLwVU01VBk
mLuPe6fLrqMSTU5tPnks31PqVZI31bVsQEUE7/Wzt9cF5RfNRcTjc6msIEJ6WpR6
c8mM+AI1lXqS31zojUVQclrwVdmQG6qse8IUiKOSsognXUQh8TfKcmNcJsYP2lkA
zxtVtXs4koHmoMIdQWIhQJNWQUpkqlLwfue99h/FCIBFfMkDpRfHINBsWfH/THVJ
rIwuTAxJgxf3WFCfCu3y/5gcCVHdVCD0xxa5bWJpJPXH7ekbv32B70yG+g3L8RSS
L4VtYMMznM5DiqTtqmlEr05MzdEsYeWmM4JVeonZfFLhzeW2jxBQuq7QHIEVk5VL
EMvOAC7zkw+0qkerUStne7cFiAKFrkHXaJ0CueBHgCD0Dmjv1+ypvhXJD7/CSzFT
D199+iY7blJNdRgYB5cyxm2kW8J9FpBOhYaARshAWmlN2NuSQ8nHt4GIuiY0RRXQ
lmumVrONIFyStWW3mWnSxqH3OmAjANEAkAdt2OweWlNf3REqrZZ2SKIV1LfMeM3J
CyjJHC9ccwm8hnou3Fp+lx01lVTRoV9ti6iphonT25h8djx5SDRNT2hi2njidnZC
ImAjbw4svBongjJvUbvt+d/uoZIqv2vDvFEDL0ZMEf7Zh87RDUpX/T9JjimaQ2ce
KiyE7jRfyFafDfBY6iW39JdbiA7dC4meU9C2mfk1GnEdrVQObcRMMsn2dpMkXagM
WsO+kXV8uOTgRhQHj1ffDr2IQR9KnOMubkr4V8edb6JNd7EtIQKPE3KiYKXx0Hbm
1Fjsmcl5gWf/lSpAA+UB6eMetzCO0gQhSi7lGunDa289yzfcWdMrTzmyiUrmiuuD
D6RU4dW2gqMN1SCvtq4F/KcLUufxfRtv2uWMeoS4hkck4lcvr/aCzpofeS0qfsI9
1JOAQ8qQz6f2gq/h05shKds/HdnhgP5mlmIYXcY3dEZ9iLFe5NCdZhkPbXrxtoFu
HJqFcDeKOicZI7c2LSVnkH/pJas2i/h5KssGzlrqv7MSgwxbZjHPsosqVSIwFxTX
qk+ITvltE+gENXc0ojFqvhcasUzwGkf+wb6f2WMwHa8iKt2nk/OTd0LiqoyYF1Os
Vd7GMF798BSDWV6SrTJqEkRI5BFvl188Ai6b+pmgCUURSoSJjkFVWDZPrnH8SG+e
i/ZFJe3X4iguw4D7NS0gPijRRyMQiThkXUr/1QJ1eI5nnsj9DxP9tahmsYZ51dAm
oX4eL1/YCj8JtBnjt5RU2wBS0esoS+/+SH3Oh9HOiwP+aWruB0nug5jax8hUZO6i
0HEPHz6u8TYbgY+Xh/z5o+pbAV2r4LbYUVeBkHH1/XF/IXWQiSo6XzT1Ua2g2sq3
wt7kx+sWWFr2Er/2CoNrdKGDsKwBuxAo7YcqUZHEoi+XaasjNp0+20x6BJmgi7ZS
xI3Tvm+447WJqsa0H1xrBqGwGRSeqZCJ/WqIeWQjTCCFFHrUpEsbwhaTnTxuR2PK
kHFKnFjG/xVzIyOGP1FlLjjSldV5VOUCTfdicZ7kdEOQoWxGVWeyGfD/7vMeCC6T
AeyvGMKJ7httke30ecMWpDku2N7gIKevD78GPwMlKjQB06m4r0oLTXYuE6oQc7+5
BNIBvDihX9YmhIRxgf2Hl8bC+mC39QMDKV/V0Nky1KLeDxXAnTJqlU5dMj591BTI
YBWV3Gk88BXbP0i+W3pPSSsy5K5K5EAAORwc8G//LRI0vZTyJoic3cEq1jp1xvTK
bFbbsD+hNPrXBAUT82aKLwVJnRC3QjOHzn3Mp9keOzkz7CPU61FPEgI46yJKxtRM
C74Pw3gkrdlacvKcr3Qizcm9NzVDVwwNdaJujXkj41uKklRuJV223d1EemMZ6E5g
nxhA5bFZ4tBW1UBSIGQrnUgUaCCGc0EFaGHL8ng4qM9wTVmJ46KhXztg9ZssNmT8
hbfCXMlknOtWacxRIfogcOWqBWiS678oQ1yJ81eNSyhhsX4XgZjFlfAyBodvtRCQ
Xfjo/bgJ4ZwR0DfkWWrH1bz7I5tAUUMQegxDpxRiZ9MEzjIhXRKapvmfSFr80ilC
Wtrbh87T+hjRk3d0wlYontVqPj3YEOAOc5+c791C1uoWHgPPsrF0mkYxSgnECvUs
tmD3MwnvPDdAhb26wXZ73v3McsIEVB8ppHfYfrU9CUEv1e+vGvYiVK+ttOCONET2
jOSFBcMZ0ScS8FapLIcjaIcYCPy1iszaFu6s2462nDQNa9Gs1CrErfXslM7bI+Nf
Gkf9L2cbskrgKyC7jvtFWYWFzdaVaj8oHWRgrGekdPDlrzaXy1ZA7RN/5tWvuf3N
4SkE0qCZPbo5fAZ0CMZmNTPw8ziIWRTNi1lY6XGOkxSaKJAqdWKVDSHIGr8uBqEU
nbIB1gacE4OYauZJLEF8pAN+iLl6dF/1ds5AhYQnyoGPdzTXM/IxnW2CrQ+ri6XP
erIiru/+PjDI5xRmDzmfH7sKk9jgdncggd7mtFGeRLj3PFPWqjLpuFFb5wGEjMrh
DX7PXw49wLE2LJ4EBygNkD5uAlkac7o/TjMT7WootNotvAAjqRqFCQ5ODjBijAWd
BUGcxtwPMoMl78iwP7fu66O92N+XFQvGskGiRjl5o+OPR03/cSHEwfxOkDZWGVF5
IaSCbzWLKgVvgoEB4dIQj+oDL2g83ho5rKERaT+zBh5zBsXloe91BD/yZatqKWfY
nPBSb7n7qXN2J+7RyzXZ/evtCPHZKaEIxgfbvgAZ3UdDIRsj2FeVoi9tgdVDIsHG
qKOVJGirRgp+BC7+puyTB7yO5BTuXIqtkf5r5ojcYS8ie5aJJ6RymEUK1Ka3N3Yu
5UhBq5tGNvqgI4vxAsSyGF9qcuAcgfVxl3sSUf9O1uZbekIoTLqVoqg3PtLOmh3q
b8CWC5HxBndnJMjxRPFJOUvZtaxmvY+CcfJruuYA1ihs3liGaYwavPq6Hyaq98Z1
aZesI187MTVEa33x/NStqteDjjM9gXCQAhN/z24VCQTNaYR01dlkPaXwtwXLnU5Q
gGOzb77rvkPWWHdoQUTEJThUVEDzHrvQjQZ3pYE2Pa8GT1p/YbXEqDktHKuoRPEq
dyIkFrUjSj+8X+1W8THi5cXPnrxM4XNpUXaDYKuyNltjIrCFZjI8JB1//TnfXjyb
+55q61EOX+d1WXwywqSD90z5wPBjZfl23oF61HlnY6+J/Zz9w1qj88/LvCU9/lK5
WFq8KZr+7cnhcfx39h2gK2aRiaLLZCqZNXEO4TRvHuQ9G9II3YbPz+Pyr5rfpslU
l9oeYUNYDsJ9hImm9+cKBAiyeiE8Hzg6+D5O3G04aGvwpkhsvvcZDAe2hKUtGep/
XTxi/vNHRjfb1MNRLlCoiTEETyjl0GBKMCwKoqYablFmOiUWXrL1LOKYB9UJtfNk
4GHzwG0YbU2WfIXRPpeJu9e/tPwIDmdAHQ9ooYuyrzYzgQoLkFkyybRhFKIYSb7j
sdk9GoshLRVzIAdPExsuN+Pt2M7po4B6Go3oTeqeRI9G8iDqlyBGgzAo9WMFWWiJ
1aAqO6sQ01zqmHkL2q67uUAuhlHe2oEZJE9jqUjo1FJEiSVc6Ljw4um4IKqwRqXA
QadGXmC9aQDtlJgln4L/onXI0SoCtz5JZLI1uH9VnC5Ip9vVKkvY2qAtJF3zn5KK
jXKge1i1zYTg6By853Cb6vLWjb3+sZ/xQkWVnEe9cuE2dBrU3gVKme558NN2XRQg
tchvH52H4s8PhVkVGHLKpqMQzewcMtSeabfADgs/0tZGJ72dOncT5rl/tnsVe0DD
CjaOX+lHPRDEHik46bkK5rsIuOy/Je2YElqpJnFZUPi10AfU4vzd7tTLwgHY4xZ7
Sc7wQn07nBKndKHfcdZJ8wI/KHoD7dKh8BUi4ezSuRvAU/9/uhyDYLOjpYV8R8SB
2A0xoPVa65jPuDfWqTVBsbSHRhxnK5LT+q1Lc4s6xnNtkUonSvHhqABf0NfINfqi
vkouWUK/qv8aKs3YOWXxpOdbcrAbjE5TcZgU5I6b0GtVxtBJgZiU3KvIIsn7PekV
my6zj1o9zX0gkXlPM2zgmnzk9xNBoH/ku0lyN6iJUx7PIenVys3WPzEE/+kWEJy3
aapfggz7w+ub8ZU1Eto6KL9pjeY88dXlcSyoqRINx8dWXdU1iUDfwV70vvoxzmFZ
In2P/aQN7TQGm+Tan6ta87tiOA4jzJHgosdfC13GGkrTo/Ui4su7s5FEK2ptfOYX
OWYrU7Wq7Be51ci9jGit5ex5jpplMhi61OoA3e+4lpZZYIyaXidCtSXBi5BDPMog
fMjaTHfaqp0lOwO9M/Izo8eSzebFZK/dC8P9XgP0JfIFRuvl0KG61he9EZpcYScs
e2M2vyhMZ0hWhz3uFqXSVJcPPpXWTFWptdGI4oQfH2hor+j6CYdCEelaryGhsxak
zWO6VkoZ/rPiYmwam1wB5l21C4sNcndLtlufnLin9wCCEBARtYKUsH8+OW0z8yUh
y5jiwbchnr7VqA8oxftW/veCnXEsbRsgUNGRgqp8r12yPVnnq6H69yBgUsQfCA7R
OxEzt3fMPC+85GKym3EfuY4SsgDeYVhf0Xg8qSu1emJYQxS6nasQgKWqQUTfUY7f
7pzDdotaxYkUcAuqmoyQoMk1G61b5iTbwA2Wx8+Gi0z/Y+3VlU+FXsPs0ujYrmhk
SmgBT0sy0LRJqckzDSwxvRO9e+tDQVld47gUseSMZVF7SyBIX8LHMK154/8dK39w
cYFGdL1uvlEm84JObWMwTE8ycxuy+Um/pMvkECHuSNBxd4dX6JsLWUx3ehEP3CI/
tunfS0dfNJu9pBKRI/aO/Jv3Va+O0bR1zr3EkYknN5oBjhqKPmEakkwsmcXc1aaX
mjtxMC7oOgqZ1CqEu+DVfOnOikFobvDdmelToHnhke7aYNgMq97UtyBAh7eh9Vxu
EM/Zw/n03SfjsNOidZEOazqOLKfZ7mPLxqlmCaCcTDhuc6NKaphGUS4R2Yhiyna0
u6HAHkDselbYZ7nPpMdwXNoUVPRscUEkxPTcKMOD5ulFq7SamFYiS3KVoRGF6uJE
8ztDDPxPnEfxitj5YhTEgDcdYzwgcYFaaKKotlOYOLK6+3al4cbqes83O7s2TIbT
MZdto6pQpUPP4ZvG9v9px3s3kVAOG32HKC2zu6NC3iJOhdIJ7Zaq9YzzpthHUlTG
j8ef2AABZWVoZrAW+yHWK3ichhDoxOnxBX7Pb0N8mehOwzPgLrm7lyvKZFKjBlCJ
praMl358uLOUtXEQyN7vKrrDwOahqPadE1Qhyw4CJAz62TBuwY8UO2dDSSIRw8uL
KDY3GTqEhozrrCjFLwS5mwpV87fRJb6kntbi3xAvC5lzH+YALy8zATu7JvdG8ydr
dY6ZGqIfyrJQrXX23ELgUSFrMufCzYqbi7ZdyRZ4K4iLeTj9MGKU9F/ham3t3ng5
jBriKJsyyTAiJb0CpIemXMU/YoQ5iNdc+hGl5OrvVzhHmQUls5/qH6JihQeM4ED3
75z1Ar64+FMGOr1gXmpuKw8LfbhY5yHxe9egGzUoem7XQq4FUkBcExvdREbl0MoX
scJzvPaZrqpyb5r1eBd8L+qCbyJGnkukmRAdxEYKR5AzC7K1NjsqaFLKtrOHAjWQ
+oY6W0NlSiv/wclRhmuhHx0hVV9A07F6xhcXwLoyyR6poyvQ/VNGD1mCc6HNxaIS
j/E9f3a5MUJiYoD1aRgKwErrXvIDgEj7bvA4W6vf1x05QXRGyLybMcIS89I65ow3
M9ZH5Wm6LN6om7igW4wil9aDqtlXT531LStf6GWgaI0GjDpgFHHVrlk60cSF1Yw1
PI9oeRdcE9SdmkCpfxRRJbyU6uf9XVI7lX2ILP4JWEdzm694vXBWfwJF84VWaHhR
3oYumeydWEE8AiOlYA1lDt/CxKy0ZHgDIWsXi38RSyU4oe6iUhEZwAKsvpA73hZr
kTauTDYqVxJ8Eeef7lTHlF47BGTlBL4xqxO/N5hHn5Da8vrxJIUH+hEd5/LBY7ip
kpS+Ye1ajaDuKsRTURqY5b3wkV4UU79M+wv8ro9Nkv15nGZCXYjsnUZt8m4M0dYd
Qtl+PhGp6AKHc13MIf11fBdNbnbjb54h9O2TmjojgQaN/ldSBjj7roIK3QySt67C
uSEKc9/pqbQJMxp4LyLifA+W8PkLT2uhdYQsDyuOBvXCmZMkS9vYh8zkYA7gxXlJ
wYkHX60jCQWSulTLljMKeWD0PnGxO65vJcIdYU08MjmGdfrAlNFGdfCEfMuiHF56
zx3Oyc2Q6XTMIzD3Z1fwGG7/37Ooy2hl8erQ/O182W5JF6yizkxElLaen2eFff0K
U9Ybvgcck9Ts66EFxquSj2WJofAtXepgC7tbpAatDPl2oxyMzE51Qux8nYEe2hQm
Cayj3JxZgYXyR5qyycGMjtPxGmbt+L3EylGmhJHvET2iLtxki92m4GepA4AnOSt6
TKx/vtz3ek004wjMFnVAj9/ASe4iQMYqKU09dlGNSiw9Ryf6aLQjlFnjk5hX0qey
w2uzeIQr7Z9zsqjSy+99XGHtwp0MSPqmaRcxi3GhtXKDA/yev25TxA5XFJ+ZY7bz
tc/WGI8BPEDHcuEQHbJHrXfCgRLk4CLeytH28eFUk0n4NAY+a3oG9atx5PBe3gcS
uQXijbNqbtopPP6vo/PupzoCYTdtxrAmi//R3L0ytDHpaJ4WusD9Gw92fRXDL6Tb
rwmOukUJYRirRHsMOV+N2hmTuNvZs66zvazXLTp+0gWGf0exPxmHo7BHeV7tjgIR
cugc3tde2mRS1N0FT0eR+mYbJYEQjRyC/IA9EbusJkzNMT8/rSwT6fZl8hq6QR9E
IfgyhqH5zKyBuB5JWt55nirfj9yGdwC6e2beMMYpXg2wWHy9QyI77XNDWsqnacqe
wo6dZDV9TjyNM2q4oSzQRilZkC3ugN/ZKbrsFlU8xYp1Ngge//b3LByFjAj1fXPk
QCw7pJAMMsgugC/lBirLlDjkoAcLHHkFMDrkSRWodt8LFXrYSvAKyHTqcpfjVaME
rRxz+vbBiT3O1xk9gzB3yQeOf5HW9pdRlZEXUzbw8GMtazA2lC796vCB42ViilOo
mIry3l1AH8kd0PKA5WhsTSgkaXDYlZRdGhS+Mo1R0ZIaSqagAbo7JY7W4xjuN2bf
ebba08FNgPy/3dBcPEP/tXC1N4tS4RQMTwPYwVc+jYwF3uBnd3WYIOjVfpZq5aUQ
ghS1rLj9JUtK1XRy7U1KH1Y/ZjEUcuDmhqkglvyHbYhTKUADTNL36gjUbcRh709s
o901bIcvC7HdHJgKV9wAWglKvIVCTQCKMHw1v3IKvChuS1NOqEEhT8NOGk7xzPQ1
uZKmz9L/RErfyTMOGQIogdcqTe/nLvZDOpzW/2xkc35uXIqPx0ahe/ncWmT+H90a
TVGD9fqoa4kSvDzjov4FA2/x0YtgT4UzH2/tRXi1UuXevDE0nlBUa3w/ZGdOQN5v
vYJJYjVe7mPQbXI5COU/UrWAsfVLFpJDwCEU3KmyjrhbmMbCj5oYwZrTkCzyhyXb
8UUjCW8gXh2AzvGIGuKd9cTvNiIfYjjI+yg1C0FSxPSWmJ5OYZ0zJoNI2KDS0b65
+S4i+lJJIlTLknigeo1QPZChrMqzBAm001jCgKfmy2HUD2UanxTKdH4NzQeFr3w/
+4KA7nEM4VA1+DLJfT6oboHk6HrimjH8MQKvHJSTPXTC2J6PP7Zsn/ybDK7XkjgZ
EoXh668BuUNElzWEMffMddAVo06D5FeDKf/rwYWPdA2eCd9DRujb+/w/xICVyzhA
q5kDuneS582qWMmFTghROIF1WlSdynkjBoH5lEBvr9O6RjQ13dDmn6disEd0dvyb
SC07vfsxul1n3h10+oQ+3RBGC81rJRMSo51AoB2Wq+r1BC/OPwGQks38ZjBquB2O
uynqzqwiBy7PwFKHg5tPWKd0l2bd6C8eLjSI86Jrl4u/RogUyyd+EkE2OfqGLT0c
SF9zSF9WI0t9FjGzjEEOWH6p402v8ax9s9ryZu+sLdQahCmG2glrTSVEE8l8oHsc
Cz0GG2oq+pRStxWUeL0ssqeNur051tBSZy/7q6xBjACi47EXKnZC7oZopM4utP5+
w0C7JyQiq/e123CdrLixGOqkdRvnVpRoxx2VpxQmAGH0VkJ+GV8XRuyMfJS4aBLK
da9nJm5DT6uDy4n6mIRGpa7YYCALhNIuBWDsTKPBTe4tAfOLNzwru+4H33zwjxIH
gmKA/2vfeRnJELvYX5edveU8nxkmx3x8DK/rUmUbm3fscqsfNcod4p8zVStrVWlV
ZV3dS5rOycEEaNmgDqmD6zXv5eX58385w/gitxVaOAhCsWSRk8x3mbspws3OlU6o
V0a8I2VMf0RRn/oTvA9EJkZrIOCoz1U38hulSnY8J5k+PEmgRUGwPID3ySDskbgV
mORvprbOnGDEIibOmqCQoyBMyYTvh0gSp5vbFfcUVRLl6WSA2bcM5zCSgqbZea+f
zlkLGJJV840UAlOGJZc1BekBhUjznWcQivVClWhPgTJKJxBAU3Rfwbvn7DkltFZz
V63fnUBJUUcmtQkZR7SSHj19pl7RnvCr0RTSi1z4JC4eSzXe6NfErkyVbTrHTTGV
fAjMUeZ8lhBfZN5qQTmIqXNwq6GYXLPubcwG+ehmG2B7ldJ6GqO8ilYvk/8Qs4FA
DSsifpZAltIrhPU1l2HMw0Kt0v6DLT5C0+Pk10rqjVyX0UYmrGQ3nPNqM9IwsPez
hz7b5zinVh21CR/muRva2LZxngCxZ1yZw+4c6HMesNE+WtixvvcOzgvjzEfNOt4D
i3MTIsWkHyS5ocmt4uoybqZ1egmXk1gyqyZOzzpqdIbkOIzlmJQA65QWmPqfs8fq
A6jyqZt4LURV3pnz90OrzhmlwrrOb3BrSKSdTRji5303imaBSchcKUQIwy7RI8Qy
ZgPLetMjqVd6tYtheTB0z2lgrIxAdpDpmKeMD+/WpjB+OCJeYiRKQh5J7teAJyCR
96TIk6NCm1WRjEuBWv/HyZC9xICBrGLP0ioU2/6SSdLJC4SPr8MGmAdzzwY5izdA
CtZv0HYTH1OD0COM6fIgaNGRmtv8X4IR8Zn7Ac0gvEFj6C8caNvWd++gwh2cF/eG
wU94i1Wh3TQkmzYhrIQao7T52M/ChL++oGlPKrF6w/A0bihahn1B9hZ7+rZg9WWS
Z3/PTL+XL1I7hfO5QJHcQfEAbNuaIHo1DmR5fI4xyNma1dlwmOn/MpSb+bkHs+W1
xKXe5BWggBHwNuEApcc3tJoJ6BMrV24vuujEHGNyUEKV52EbJj2KZ1JaW6L3QFSZ
ZOZsWDUzrcf9O50tTr9BtekRr7mi75oSt6lxvXGa5MxjGgCIWWJRqmTBopLnhvlJ
eur0+gtGxPeTnaVPzo1qFUMs9GMQed/uktGphmVMys36wq1YF7PntsX84JDbFDRV
8tXsqNDdSQePR75w66a7UFil9dKJ8ATG/n77Vk3RuWBBnxxlieSn0Eb95xAZWDmV
MwPVPMGIqDBA42vR+BKS17VedY05SvvEwgD/BTpB/j6/ncvUwqbB0JGFSM4e1n9d
BpwGWL0ihSP4bHrEld35q9KTi0W12qgWF/29oDd9R1TGFa0MKcY16ke4aqh2osiR
QA7xH+uhzPQAJciS8HL8NR3H6ab+NaBxQ3VUb2NbW/Jh+KZj3vRSVo5YO4UWaXAc
g+qDU9Bwr2j/XrazJdsJnWyUnfZ4MqwPgkFwcgtiukZWh+BlTRpRcfsAaKMBO3qz
2FLS20jL4CNRnCffzjHp1fKsbMjp4jQJ9tHIPYrqNbSQwq0mr8hBlJoRaxuepMCn
EzD6awRMQ68Wn4RLI+u4lhs9eEI80L5csP1qd/nr2hBuEocAviu6ZW+A3v8JZ1JP
KwZ8xwYMiKHYyXei0f10GWz59hx+HnCVfOfEGa+n1b3giMXcEXysNtrOc895X0w1
DxSXTtIwF3AnQHLjA6wSjwtzrnoB+vxPZJ8oZua56iPux3ChWLNFYcbDJqtudhsE
EPp99hqm8Qr7Gzp99+i7csh3ZxxskmYTx8yRvFJYadgx/o+WcgaISeDd1v7eqJW4
IyXg5dmBKCVQ3x0mQyQTQrhbHdFb/MRwY1fVGiqLKkH4zQSmlFROsMzsgq0ihxr8
SOK2+Bt/ikljeOcdXu262Gb7xUlDBWD680dd8Jt9oZ0GLrLPeiA3+zQXL4RYM8lf
NxNuqPCNzOdj6c0nRTOw9k3kYdEO5fEbx1gMet13Ba/Ey8y9uIldsqJyP0qyMmil
GXesu0AIr+UGokKSaUmTgl6qLa8LFBvD/V6+0GeP5/rwmXC/G4WIA6I0QOWpHfvy
3nSfMGs1s/7YGy5xgnLprz8kp+7wWZEezz8DoOnOjp4VKu3byzk9T7kDpB6WZXc6
GS13UYlWednc0uFGFVijFjEouwxfX8po/p9NSZ1Ep/IHJ5jGTQHoK5JhIAISk4vY
5J0pbK9vasxntm6/ws+1To9jfkQq4n+lh9lgEPMpmwc8N9m/r1VklwqXKZpVIoxL
wm0/7vnwU6PDV+4N83XuIoD2NVc/FXE4VYEonD5I2EKOJw2qSHPyAPstC61FvGwS
fJwtY9fd4uAmRDLmgsboCTpTj5oWBMJBH73lKU9cQ3be0K5UhjBWXR8c6GS1M0uk
jj7pP/mVE2tp5UnAsFmS9XEfrVESfQ52XAHx5zJhfz2343dLfro/p/pG1xTXicgb
6dztX/m/0qUV/tDs/vH61YJoJtAFrZFEVI7AU/4svfsr+8sWpuJ/MSrAxIcNJEnd
kq6chXsy88zkmAD2naeP74eR2RtaUy2fqI3p0Wl1QtjIpUQSK3joxCcv4RkNueoG
5CupJ4Q8hyDp4HFCEjxiZKGUThdwb1m73L3FYhKzs3zXXhvlFwbl298EyYbLytG1
G78Rn37Gw1/8YzhcU+NXcOekYW3XLaLIBmyWOEP8RNarvZ8uR8mitKU1HivRGq0m
BHaDuGoDv5Z1LSDDzd4mPkgkTdk1LtZT5c4o6jXJneKRVeIRU1i7a/PObxix4kAg
dMgG43wv3DmqVkUpeeP9ZPKWFOES0EwEajHl7Pe7NH1uzAq+jZEoJC8QtXv/kQkz
Drb31RxwyVkOEbyOq56jjRSLAjn04OmcQSzaWMhiAjPoFTAuhjxOT7bK/CBtMrHM
je4Tyhxs76YccuUoPurve+bos6/ZsJCqg14RkAtUWUG7M6kJssJe+gHSQ09QYEVF
KHjQBcgZfUuW0Lq97i46gjFr6GKnuc+R4j/q4yZwTLHyBFjo/2Sb9fUGcsSHiZUF
xNejGnSY23vdb3EyO4SOJr2AA5xA0MaqdgPi6r6Pv0++6IFqsWwp8uz4QmkLGri8
kSGQfVmwu4Vd6LYGhxrujz7x+OqbUx2v68YNErZpH/6jB0eejPXYu4t0S8cgWWYM
doxioW7N/2uzUjwSsNAKm/BjggLF4rn/M7zSleUZxJEA3IwY0poTzDvF4Soe704c
DKe9zYKz1t8bql9K44ku7LkjMBhz4NkZaV3wg9hkEMPXhNXJsqBQ/zW9YvGpzsWz
Tz/jZzZFxEVNw7rEBcqCBwfVVon4BT0kb2oNfC8DSFJf9OKoieg/5e274dvfTXr7
l2mBP37uDKcdP9HR3E4/pIUTbVdQz9P2aSc3RUFE0FFyoYuLXsQerAL29Z71AWnz
bTW72gUQ6/NVf+Go2b6/WX4Kc2ZLQNqrHNdDAPEULbw/kaU5IsxzdLo/F1RsZt/K
GgETG5TXqZKXvAqq2ks1wPF60pwe7vZXNWp7Lf8jiWaTXAdOI5CEs4clItdsAbdn
X/iG6cuQbE9xxLpE1RnkW6ckXIFHxgRkqhxKAVjF3v0txJI73XwJpc3Ys+kvAFAx
cKgbaiSoLw9JTZoWvE1bUerpYiWDDizrjtOR5au4UbLiq7TdfCgM8T93VxawaHYk
XFfCadkAq1rLR417hCwogQtZ+4ulPNHpkqYqOZxF6X9yNxxRZAIOx2yJcKvUYw+G
3IrUAOIb9LQTBIuBAV6BVET0BSwg58vtfoajiAGJi72rlO0LTKyBFQP8V9xIdK0V
KFg9dLKYydxug//3J0630CXUfY4t0Yeye1tekCNUem8Afv3B02moJ8iw8Vh67pQw
cfIKWlNIQDbTx2dtwlua1XG+UaRMU2JVWHTOi5HQk50ZR1YmLB5RFBaDyA5BAVok
AJC8QXNl8fHAiqfPeVugehh5jR2Ckph0uWIWSL6usDtcU+mt8xq8wPQa+eXbOeQe
zss2OTK6OZaHtJ97uopbKAHbW3cgd9RK6aTUXiOBS5yzl2hNGQ/kKUry9lvn6Pmd
60E7150ZxgUofvbtg1YKQ7gmLqqFGaSbsEsKdsATt1wmS15joINxZ3+FVUjOiQUd
7trgKhyhcap2/WDgylHAy6Z5KNVaKxLadLOUlgXyn1ZJKAxBvE2tsEZ4DASjKDMd
jno2aP/usVPios4R26j8ZiKFkeLl0wwA+yTlh4UY3mZNH7yuVvWfOCgJpgdvNqjO
4eVF6MJYcS5h+A9AmayNSmpvwspwhREm2vVjhPdfG5bfiPIoNPQehlxmuw+PCvuu
63Oe79MS5xyOJrwKas/rZSMDCZ3agcPx2AuOXgOQv1SRIysZEWzoHpfkcpPEqPAR
9KOevuWNWrP5y8Yar/jA+6fX0DfwFCZ0pRIlQ0YTlIXGOnAgTMpysytnfGlo1OjQ
98B4HrqyZIA6El5cb0T4CAiI4F/rM1EzCEXCE9ehGbtG+oW26CerUV5+Jya0PULX
jnxTt+3HDzpmePTpWMihDxc8eQLwHkuebBeDJCT7TzZsYM757BTkIzNPPJZ7iQM1
2YywFqFLma9E4K+/EejOV4hfJH0mHyxoOZkJw+oopNuUS0oLV9aIh2OMDMxjyzej
Sf9vKiYa3YIsyOQ7BBnjAb5WKq+Uu+l9Zmsz1Jl7K/juDPMkIHP9lb7jydQbu5IU
jim4H0pDcPkZx+ii86krtbs7vsHhYrhApEE+t3GfNRHxT2CzWCEaZupjmDGehjbA
AqUh/KfGAeKsxVjM8YBRW2coBrc3DEIkC8LUOqT1q7byVG11M3xCv6hoo5Ji/Rk5
DkXp1YlLT7Pm/6X4ZxdCszMkRrykbCy6KWA2WBMVDU+bg1uSLuqFYYEK2B8gP23G
oFTOT1wD3eaoeAGcffo1H39knT7kU2ZiPUWH3wwbp6cjuVGoLArSKhk4GQ77DrUc
akE6r8b1AVM3OZ1amjibHE6wKSuWnEfoeIW7zapEsu5j/LGpwe5hzr04FuTT7kYb
vK12+AaQGP2/nXiGS8jT4j80yWGZ7JviKE3Z4OZruxkCplRTVsv1plEt2g9EoT1j
6u6Q7FiHbh2Q3Ukkr1DEkDXV2oW9ZyLIWVOrc4Vi6k2Eewv2zsOouyq9nH74r8Sz
uJmN9t0fFe/AIJdBOsI3xUReKdRHGEymH/YD71C2aBJzwv2i7a/gW+j2V72FteVm
q/TOhmrgEyNV3ljb9SvodBGrWp3co4Rmhg8ESgXCzjXLZo2tvpb4EzwBuGmiLcRR
9qP7ZiYWmHKxao3cuL7/XHbu9Kzfgv/tYQrzG6kzArkeS8xNgf+1zsLEY2aPg+ip
VBPrRMmz1nxqFCg6NJs3LZtvhq0OmF/B74U/ICd3lVZf0crCLOON9WBvy/n1nsL6
kW+Ua6c6nwLvd/6FvZZrkYcvpak3DTAiPO8CZ0bp1WdygwOvtcJIzpIXIJHZPXAt
yHpIbDsHiQoHcC6DAWG0oO8q7UzSf/czp2iaHV6C2BdVRyZHz5e++wtFLz0+jLq0
dc/Ou8BuJXiXdDpWbXuutlczUEr55VuqeWMD1sELjcTyygueWJ5b0mGIu2BzWC4v
65cJGnjWM36WrH0+WdLyOGCOaAfiIYkEToKaTkngiIVtu/4l6UEpriMQ07IG3ZXM
pbkovWTbrqBPLYIld4pS/kTVtvlp0MkllP6M58J8wiQ8KQiinmf67SktuiDRW7z6
hmpmEAKbiWPT1kwcmSiYoWYpBWamR5b8kX3Pkg/RNERslKqNAzBoh7LdvEKdKQqf
n+1LMsx1ci3TKgkUDmNJ2yLVWohuPxQXpzvvfl7q7vv25h48dFM+ktYQxYr6r0Fx
HwAfk7niYCMkaIBuDK3YhigtR5uqXiNsd03W8+mdEveuQyu6cnXIlF5EHtURpq2y
S4sThrMWw7271vD/LVDsPfG9UkSIxfs70qJCyf/4X73NmFWimEHKw9USPSjfAj1i
SM1/t5Hoe+drAjUpoP79JzvLnzNUcXUWSok+PeQ/UhkAhrn2P2qcNG+DOPdcmnaf
CwLg0+vks/Lr6hpKi+5G+MoyIok2yD938SVFayc+JKG4cLPMJDQI1U6iyDHADnUB
T990GVSoueQDMqTlcek0uge/G/eSNz3V3ExHAHep4KjOs2fHFEmiQP842bPU/gtw
J44CKrrcOgdpg5gtAbeSy7PvOe0VFyuLCU1x4cZU9gGJxFDodh8rM1JDfChtawQu
+tYM3UkxixQPkYWmgavVDybkqfIIeLXG0ug7h44RUMz/ZVHylR/7s8QI65zji5PZ
jLMxXmjzw8epJ9QthTcxtd1uKGGKeQcnoq4NQ3Ri+63z1WlgCLt1DMEerRx+14P1
bDQwLxYL6uKgVUcWoWjsTwKWGWCnLPSQkoxs5a5wvDGDHdxzcSb+5TN/7TZ7c1be
wPet37OCQKKq0dyfpjaBienuKuvI1gp7v8zyLfKeE6/DExkp8214YyHjdLnaIMf+
iqLW10zj2EKeWl4N0mF4FzGuQLKUNhFERTlfG2icP4gMF0iQsMr+w63Clx6dVAzy
sXm2ntDs1QXcv8qgDAAlgd9SH5gMryyK+BQHtjaAyWnB9loO0HROapeLIeDbGWhd
Fdj+lwljdEeyMszmRaLsGl6/ZypCpUkcpYeDzcLa9KfkgWttPYegYuZuf9NZVIx5
fvYUJymM2LwTLX6Rs9DAwd8VbXXiTpTDXrZoOhSUWdgJ33CzQW3Y/twxszES/xU3
4R3PCfCe0dSGsGZgYOBRPCM9PN4q4NP84ArNDLPMxAvcvDfM2zcqk4gGGRNV5d+/
Agy5BmkbnQck5HlzqxoEHZ3PJQq7AtsdvxTITT3Uo1Inhw3yJ/vZfMCBqVe1n4PB
dn9AeYR9eJ9ho1W7UkZ0CxXFhxd0fZEUaenAW9tsmn0hsbCDOwCScl47rGFrjCEe
fAezjmdnbhLKBY9qe3T9yUjO91/4fMNhFalaB+QGIsNjRqauvzaN7zjIgXgRqetS
X4hj+XoMHU83cDd7tOqydi64vFtFzq1dK4uFgOXh/+ZqqX9mZr/FJA07rDuXj32p
4TJhjDtduL72UdU5mB16QG5ZF7KaOMQkq/W1eyKM9LIU0aWNicagZNvXJcPTANeo
OmlTEymcFTYHAZFDnr/3fI5zOTwbUkNpMqrgNcsMdDC8DmqMBXCUjz3RBDjnUsud
sCBYiL4t3pfz1YLBzw2WLhd261kXs//wcmnKFcweVEkkHwZQfutgJ/rQx1x0EfyL
GjyEW1eOv+O3iKh19MjjKHKcIAjR8+pPaBQkxp972Lqa5owRzAqVst7foprXxX1y
dEFzWzzriXyGOpo4UEAMxPlDw6ZeW9ANrAL9GwP2HCPeGwpglX8YhTA+ZEwrCA+r
lq9muDSurXLwKB4Pewe7B7fd8UHxgXzhxkTzUUQ/NOhXM7ygKBYSSyONMxy8LkZH
9c9HbtFDH8NdaDspl000DUvjQvr3Ln5SfPBaZ6Tvw9FMXmh2OM5AXyqZzFSCfCr/
NVgnQhyPnjilQmxfLr9har6kJormBdPfNzTniOEhlnZBOIOyxXCB7TcXQBn2AL9k
SkDbr1kXY7Wic58w12T3xZcyPD83AZKravHGQSHE1PvM1dtZ67AjWT26HZkxx7ki
02HeQogerNH3l2dTWmuTo7kQwjdC4bOJc+pXylCt86famqdhRXBLFNF03eXepLeA
zN97BJ1/JotsOacC/B1zX8nz+vg6x11sWRiymh8fYrol1Y9FZrSMRnTNlgAFdnvE
HxycIpQnxfcZjHB3+T15Tv60c4Rqk80KPaetlVHJ/bdH0Ys4SrDZPFAjQDILJm+3
K0zSKep7lDXhSxWetJGMkeYJI9BGSjfP+xR3klZyeC8YJL8rr2Q6XcATA8KiruY0
o1WZHr9A7FklawQJsBV2jd1sfql9dcTIOFSI/+RPtbefEH0wcrkCQbHDrUMp7IDd
SR7/czq9+ZAUQGqzEEK78nB5sLhwXkJMD3jrHav9XmYr9/Klfk3GxzL79cYq1lRR
a1swR9aL+xluZ83KVlqRb/xda03yZjV8CEGvuBnGVIf/ajk4UmtPaOudLJhZn5U7
Aq0/zA6Vk0xjP15p9hKyRpz0+2uJnub4Ss9JepJBKfqdH6OgcE/kUDUhCvyzImHd
PgiWmPn7NjdtABBRT4kOuFtOV3tAyInXyG/GfX0o0y+zoZeBp2ejscHGjspcnrL9
imrmdemMFUKFweKZnuZJNckNjj4ZmMUrO8Cs1IVGsF2s3qNMZ7MAoCojWNwITLNw
CtVhMhP190ySziD8EjBNxJRiY14OQuw/DRzYKpa25p8yLI9ORr/YohAZ7GMgaD5y
uTgFpIoabyTi27SVrFJmorsWnlZdJMUeQAkV/4qlTIRDkLdsiF/S290HBzcqhibS
1efZtf8lEcB0ahzgaQOUa0hgxIdi74fmQVyl1VKRvUrBtHbjh473zd9oFdep+uFr
VDp9rV4xpUAtGp+EEOuNcSXG+3G8iKMdAZMEFdLFaqq9L58GaUbSfPp77USQ+umD
eHDJp/Eldz1z71fUfNyzib60sS+rg9Ok9HgBUub9B/JaF++h+o1KlkHUOifQ9BZY
6zNUrD3ySV6EbzU+18PFSgfW+XAS4GwPq9Xd8tq9A902ac7rwDA/LY8C6cxIhvy8
5pXk5FKTO4SvSA734ctNCIPZ+Wz9cYWZXI38HQYcmY9Vs7/v3ILTPjNnqouY4m2G
iqkc9vBNqjgoLVJlNb9ytK6BW+KtEKCgwYMIt87cd31lCrX6lks5ymjeJJgJimLE
15166R99MMUqr1C++DhFyEqGNFrotEtihsFliyqqkzItdy2XYHbdrZo1972bIjFr
mgFlji7uVBTetJhqIoed9W6UXh/WjiRlcsvcH4Z2OkuAgfQbGNJFl2C4C3qXIIny
eW1Pg5N/fikC+U2nlfaWHak856sXjk9WmdObe3cegwmVkvBzc6plMEJlkxL5RjTj
Y10hzQmV46rp2PEoHYeuWZEO2/Oy0RqDDL3JL0hBcaWzHpqisDQjwG6wmPSjD9DI
pVREy0TYDrcSCz0bIPUotmZocEsqITsfESJ3jUpazexA8qmsCfx0ydNYMjsiMRy4
qw0lDJ6nM7scn5vWmg6kRRjXBWwN8oam/+kRGAyeOpQHhd2tid8brCgzTd4I+oMO
GekO8RGZ1Okjym0L5bsbuY0Q1xynk7Nmdy/OB1g+CAsc3q2R8JV2c+z73XesYWos
Mw7ePl25R/c0UR0Q8Dlsu4NJgXRiaatDFDj034jfodMuy//gil1sHRE24WBdZ4e2
NPyPOonSyp+MMmr04Rdf4UEyWyvBhLRIUGMe3bQBjLselwjq2b7E7YNOthhW0xOW
16ZX//g1E+hsyOFjgWgRiJ3d/UyAzVP8/8CJDrFJUADwZezNoU1q6sz8QCatFTXL
pqmw/TWCJ6vYU5KNMfnSM8/4j/SWPDrOaEEa3krChWamc8ItZBnB9xYMWfSzSYcu
eEb7ufSAZ6CVKa1j7bI0vCV3xVPqf5zR79JngeiYDuWWC8vfPB1kzbCEO1on9ss+
Sn5WnhJiUvWQgePn2BkkgRStIyptz6B3E6jH0XylzZRxlSDmueP0kx0i6V/a/m71
4UecqBbXDeFWSRSvPBbOcT+rCkXwDfAEfM9fgPIeY9mJp4cmS1geUqq9YLk2sDj+
edHfe8URxbXBkCBBVaPkGbow6w3C6AdyhI2RagYY0ZV8PFPCACuhJLKOwgejRd01
BsQHocOxgd4r3njCnyLiRqcb//3ah61w7SK9hon/bssSCSP/6O1lIdnyNkwW40zC
2afdnDguMERYEk6V4FkYhy7PuJwicubPMQDyf09SU6FtLx7iPkmfQNGK6r5ueHNZ
mCqr0tKnbrlXvE1rHq/E6rK91l1HbgfHU9WVRlUQAABpQOyl/w4yARj2HRb1Xazk
m7tCeNU8+nNfMwFI3tiyn+bnT7bxRJnwIk8GvTkaaGd9/QZ2mLzXS+IYHBURApzI
FWQCRFq4liGwbN2TjsVJVPcYPI5AI8B8fUGfTQxAdxgsK/A3fGlp3SJsvCxMxAaY
Cvd97KKwqMeza2AUTpUJ5FUXdksMGAboOLSUS8ZRXtnCpx1ENZCJH0KQo03gB/C6
hjETh6Ald/YOw/BXQQqYe2WNzqNUIj+988HcDjDbb2rD0O4FRZ4ibLlMIVCkscNq
uI8tEG6rfBiAzt5D0umjt1Zt/KH5wy5Vzyq+SOd49FrvhVWy2mae9tgZ3IpFFwdP
8RG7T8VkyisblyoB0LWYt8NN3fgJySoXM7T4AJqQRldahuPdGnurMiSO/DuxpUR2
OZdbOyndwLnjsEjlAR6bue1nLfuspdbQkeEDcO56tjQgfaUlIP2QBq3UJox2NSV5
BbviLqnuxeFza4aKIXeDafI0/FbBwlf7NBm6tpQIFIh7gP8zlZEb1wGTfGvhJFD1
D/P8woiXwX3RjgY4jVpLZHtK7Gy3ZEYA9rvjMsiUmqUoOwxCXpY7msbOImFYrrzF
OvfxEUNTtpeE/l/FZtapJYgsO1ioaUFT/xHug8BrufPi6p1UTwhzWFwdn6T3FK4A
DaLSoFK5/4c/ZdcYK65ifoywjrDKeFVmLgH5kyn5kJP5fXO/YHDhK1ROIyXUwHZb
22ZZDV+G2d5P+qvLc7PVXKJoeWfh8+f0rfWuRUakSLIfXgrDfKlfm8KUnDYxd7/T
YerojDhCmrO7S1xAL49uI2YURcDPpRDf/BBTvbDgbnYqU2Aqoc4VJJlCEyrugftF
2HdVEea4w7SkQAhxEsQ3y6EY/ZM7qKPCHu7gYlO2xRXmnsOWsBFtbDFf7VsppC/S
lXGIrEav86ttkY00fPQd7qkAyz6sKlgOCDodF8YpfxnsOL/Xv4a0r/pO8NSOLc+b
gXTG6/RfX98RB9Kvitvi/AGNl6wCxusjWGgeuVWBSZm4fzmrnPxUYywWJM67GaQp
vvRSPRPYkOhzER08Q8wGu1Kl8bXG29nn3fdV2VgNcMsPNiZAZE0ZwxMGTqGoubEs
yKOef70XVhWJzseupvM/JEncJ9spKRb+XqG5J9tXLLDHFuGMWdqWm9Z6wcsUHUkP
ce8rJ7VaKVwzjuLtyQssAsXVVYtec+MM6TevSh3uKiN/f+d+7fuy7UgKAQj5/HJo
Nlu1WWVGXX7cwcRXtDneNdlIM2HVCw6iX6iY3N8vaSB5lY8uNbO/ZPVlb2eyKrU0
W6g3Op8Ju1fwwjhFuszhGQb9UTml7/JwCdigBak+T37clA+0RPNJngk88eFEHTix
K9iFpeh4iFMkTx9kz96tlgFVZFiyhSjaAnOTolqExtnraK/j4Ys9AK+wdrOeZz4r
rXsA/CNGrSO04VwYLDBnaEzBXp+55kw60vvJgIp8RQKcyU5gPq+lhZaPPhCXa2NT
QcGxMJOYbt4Wb3H8LVEkLrTbJygtvdAM3zIFzrOccP+xLxqeBlQvz2neM0RDSziy
L7wFkUCDIs0EK1vHv/phP6sX9+Je4z1o2alstRhPQiiW+6+8RDz47HSCJzhYA0Ik
NLKkDIoDvb+le/26sHnwZ59JVy58akiCEZiZ043koP9utm19RRzqL2DTnte+MsAF
3cabnyoUbNHti210O4kCdZqb3smNUChfgb2gcffweUnlfZYBgDz7u8hoBBzTh1Zr
aKxxpyG6kI33pk9PvqDmGffgfoyOFRIl2zTpFqRfxvIEcHxSD1XMjdE4LqIUGWmg
/AkbGjBgc+1Z+J6REBmXyRjqYGRb4hTOJ8/pCzFa9J+oxSRAKPVXcDW5AhO/1hxv
MN3PyuboJTzz0UvMbROaaoFfEmVxKEWQPto2qqn7XvAR1CWWGetWIjhLn0uH8fD6
c2tHb8fIQXDi91xFnmo0J6ZlQkjtQZEdVnOt6LYyCkG4+yNtj1Ky+Bq0NWM8PZCt
rYjK55iTiOGbvz5/xOjRc5SUbJLMXqiivefiPSnrb01ZWaE5nvnHuP59KsMgPAKQ
9RZQe18AjERny4hSkmlk+7Nbxa2tjaq3jXnMCbH7LcuJcjTCM8YKQNmtYu/3wC+A
r0JtFtdeATxffVRWJMG+iBgO6iqwe5WqTaR8L3/hRMORgDk8rc0hClLt7YEytILM
HKfA3Me6Yk2Uwg63Fkm3zh/+zzy9bgchKMu5+f1jwZSyZ7b2ZwkmCWB0Ud+kopZq
KwWj4Q8MXDeP3XZKCIWX8t2hHgYpUEjyoNg3NjKA5hdcBX61AbyAJZZgmeezme6I
P6tjvw1IcJRXbKqCK9UWHRVdOvnSMmRbwLE6QTJX7QVgYl8uL4sgDr51uQE7C/Sj
39h8GHxYpZ8BJGqm8ikGxCbPjF6rIZ/h6yUqvw5p9sXDxGEnlCR2aZ8uVio8V8F4
BeW0HNx1iktOsSZ8xxG6L+EKmbV/hPgiuhdAw9+4DqKEB1rdU5V+sfg4SKbvNaVv
kY1V/V2RUz3NtzHs9F1yVhZ7FURgcwz+zq9YRicNkYLayBFxyUtcdzkqaGgWdEG1
vzF+TuLOD1IC0uWONMfDOzg9LY78M1YuEovkVmEQGpYGHzntqLi6MWUKcmZbnQnq
/CggX1SGc6KRD0wxde/03Fp9bl9A24C2aOReKRDAq50nc7CioiapHxQ8BCBiAVrF
Yrnb90XdHyhd9xzeEWWzX5w9nD+QCa3eicGKBfTNkhFXI1wZwW8oSmEpET/C5scb
WfJgd/tpqq6Gl+pkkMBs7kA9nElYVwWit46SLd/2P4tn+y+QewVdFcSSqG45FtBK
ugENtKoHXaNc+Lisbf0OW8u/z78h5zhDGfdKOLqOucHvAJYDO1+TlZkzbuygf4st
IdJ+LMkjk8czir15nYmwBxRbbV7uOTJj/WdixaRD4Bc88RxgFJj0L56MsJrGg+0m
7I5z5qfnj0wkOsjSGtewy7W3rH8KYxqNar4lV8tsq9uyyQj6IM0T8xIAeGtk6hNE
fSbrpZK0l5PnvO5uCTH6gFlYCuJUUHx0/81cy0AgKl60GeodLIZpqjIWTvP7Mn4b
66pDlHVyjs7iOaDE9ZHsbwvGGUv/iBlp/bxcjcirdgpYoxZS+r+lrksLHexYrTV6
iLPueNA6uaBe4x3qJ4b32tXBh+K9et3hrpV5b+/Llwdd7/de0OU0i6IozSbATPDc
C4g/EZ7hKZg/bOHHtGshMT2UVK7Qovle0AhyQXE82/aqUrIAADIp2VScPOUIWHbW
9uOv0kElnPMcJY8NSP7TGJ4dfDVcAGHBzL7U7x+ayJHNi/noYaIR693mAidGGyU0
oLrHgfLyToFk90DdLCjd1ItaLTwOildc4AIU7jveIGa+8/qe27x9Z4cA/yM8qxIE
UrQc9X2dWnzxDTjx12Srd3q8z0Pj4+b60qa4dBvH0D04U/9FBF7OUuAw2J7ZBqmM
c4ch5wvgTwLVIYrLqV5oQSi2GbvEED6QGN1YL+7+sS+MvjpaZdyChM2l8pPLP54h
v13HpmYlfimtxonP5fXEqXzci6kOMYl0/sWc/HvYJ2Ox/qBp0WUvjJpnX38TSW2N
QvRLwItrCxeTgtlhjgTQzBjDn0zKsHci2o16VUegRf5bMSnBKZgOc4FAycX74CjF
CzR18kicpf9uo1wZvgutrMhg9FxwUGAA2557Bq8BNL52WxQiyLi0gUYSeztexGOm
Y/WPWC0Ijk5sQGaiCZSfVRUM17rMEOliPtb0wST5vNnxO8apxNmgAu5aHLowGiBT
uXlmxEVSqCDvJXcfQgBzY7Fzm95SKUtKQgIhRhWTcyVukcmxXbX6i+omAAxbUuzl
UNB4bkcksARjNtOXb6ivBlYuok9EQClPkWKnlpQhy9TCc4EnQu831sFaCLMfkxBJ
EhhwQItdXVvPa05+vE8ifbd2L01tFOdw0ETXJnUs2SbwN0O3VRHwgXRnWfRucNAZ
3M642pbw5oBZ7k0l7giZAo6zLMg+0/nkRDMgtfcIKaB6dT8KjXWRf2C+pX/VB638
T3cMjLV9SFXdZwav7p0JgNfDefTtu/u2lY0ZA0qXhKuBkPSOYOBqnP0tlIXZSPBj
mu4Ekta5UTi8RskpwPoHXe7v9QdekewRjtEjHMNsSg/dMa7VH4wc+SLdtyNuTnW9
SYS7WLZKjMkIWRLsMewYzBBDWLa8bOxwFCW0UhI2ikB1mIa7opaxNSr8VTtqyeAS
M7wzhnQBpMpVCyTY1dYQmMvU5NIE8QTmpuFgd961TWUnWrX84PgRfTnLApYukquD
9DHm6+uNcD8PT2A3hzNdUXfmGp1DMnDukx+aVQ4INH1jMVtboxx1dYyzIIJbIKeQ
mWy95Tu9d/rd4NFuDrLGqDHvWEMKRHDsvFtA+BY4k0iM6NTlyotB5BWG/l6cBbX4
uMa31+hZrWEHH87hrcLtAZGp9yb8aUjlMsDAujNlDtvOB1hUtJIGSr2jjyL7oPAQ
jOiolgw5f6ePh/W/tJr/9lEdBkn9caXtLfVKVrl742y22xpcaPSDnr9cVZU8V1Ti
dF2zvHo7ZfbJvMMjPuW7sa3o0x54DixMCJP3dybMc8AtwHdzz+AR7iPKHFVypcMi
vvt/qSl+VFqAI5r9uMrbMI19avFb+IufABcCJhSa7KLD6978sjELkROK2JjOoqge
k8Px2BFb+5cBfUurYhvEzgjdbKcMEs8i/YEtqmyRs0RUtke1WjRNkA/tLd57fZW4
gSIYwuznNuCrNWiTUMBqXH3kCf7G7m4PU8a7tCvy0D1UyOiD/jFpAsu1KGoPF4wg
G7HyIXhruuVKB4vTr3Jz6dAePL+i7bTghuRDDfxxxA+rkw3l/fdkz3+s3ks1sw5N
v8vXu+yf0dCwFwixxc81VAXkZK8cvh8wz+fZySC7vkCWbc20kMfW6Ao+YB+uAWJM
dnqnOzQJpFaxxNtcdJxRlHGwFvosiG8oIsKhDJSJd3F0t3UPar56LWIeew20iY6I
fF0aa4rxVUHOJV669sFeBSojGay83/kQ8aRUgM02cOu7/Ll4F8i6TSyJbHCmDI+H
YR4U1QOMc47z2eU2RNrriM3EhXeyu2AMdqEa7P4YfE8ZtzSUqJuUv5x3Pcy/3IS4
TM0dZJHIxQFObwPdeyhfhLlTwUQuOt7ditqRHYQlN8IX2kXXmAa5JR/wLX7BhM/K
hlPRuhrWiKz7gnX0VtGrW3r9qRVCKpZKuo8uCv0wXVMr2EJ+ntzYNpMiyyVwOhY2
JohGfV928XZuDV2EYDAEbTD/6jl6kDAyNzexgVGbZ3b77sPluXDlg8PPmUgTt/nC
oOMVjlpSuE0LOEBo2uPiBntGe9VZjQZqiKcg/mNUNeULH3kAA7kNPpMQ8h6L9j2P
3oBPwzO7Pr5LFA4MNIRie5dJFgckkyLxZ7aSToYNawx/Gnkl2oOGJMFLZr+mD6hM
vxoHGe0c02ti92ttve3NtuNc3s/R4PjgqS0PS3oJRAN30y7NCCdVROlpzKdeT4Ig
u0k6aXa2gKYt96f7tvJhvX51fj33xwSIXxlbX3Gx9rind979/UIebSESjtQQaEZp
Mrnh5UEjY+oJ4Cx1QjvsYE6Mm2A1usItB6c3OBMitvh6EbE4jr0P6Fbi+FOHu+tm
JsGsDBfzNqOHcpGghQydWJtmRs4QLEz9XyKdlkBD0WroN8H/ZwqcIWmEh3rJiY1x
zUHM2f4EsTVgiGtz88IsIlsgux8xkxrjGoNmjGA7qTpY0ADnRIr3+8i1ga8Mmf79
EgtB7Y8+yV+Z47aArfP3bEMuooq3byxJybEdrs91Unr83TX/49nB7kK72TtjgGWl
+DkEXneZUF8qzvIMHNrtDmb8mP0QfwRg1VqGVyID8p2whlN2oPIZbrrIb/BjVwo8
mqPkeVRMXpOUX3jP0y1nC+LkvQlo9o0fA1u0MFzA9lUkLgdA8lvbaGgR1oiRZo25
iUgwJ/c6evmHBZv/pmm4zJs/Zk5EuZGNOqRyFYf9Mt/sr8HdKy4nbgAyE5W/w0Ir
hbZQHrFNhvc974mtIhyXlq3U1wUP2EdpCJaLTlpe+wIYm92LCPKIlEY3yUJz10Cr
VSrTJV4XUXBYRPKezCQi4l3fBGakAUdeC+kdcFU3KSnD23+irO4B0UqGw1TKEU05
DWugocM0C5+ma/IsV7emHN4lnjF2+Ae7SYQV00qBqoGeCImI4RRwkI+w/HO08Ytr
FUDVGK9+Unhvj2uXkHx2k9eS3nRw53nlq9noDPF/ZHQHbjRUpXCZECPMlEAN6y4r
HSc/EdxSAU1Ps1q5Vaq8SZSWnm7thNoKJ8BrbyVxdRviY3YLs91agaqtrVvMxTDl
w1OdzcNLcflVoOdvNZqaF7sEHF8bkFcSaeYc3LMp5xZmXfV2qjzClzl/mjOKkvQa
DlI6mUhvBVUDEW0gFQNVXaA2Pk22KvtsChFFm62HA/57EJo4tXg0RKJ6ProYf35/
lnGu8M8NTbvkp/em6dUtyJm9lxu5qlLUfguiOPdAsnJN/vVsYnNcV01hlONYxvYA
SKte42O5F21aHkZ8PCdCbPpw6ND5HX14ApPZoDhbSRma22TUgAfasT6vztpm2cpG
V5jgZUGCtoz07WDobkRq3c6DKith2qZrhksugbk8UMPzjWjLOS4sQOQ2srO3NygN
0YracBc9MOODZsl1/Wg9/Q57ZZvifwfBbZkNegqDq8fQTlAmcpxUKwYaIn9dAIiK
9QdnlLucLBxaI/YetuxVIYOvFjQLrBi+FKz2UUyd5lhsZOCNGVhr8sPuuob+eDd+
CzU1bGLOPZzTWnI3Ao6RAdY6P4KLSLoVOF+GLL3n4Ia0D0/Yoj9FiMSPsmRK7KmP
S1Yuqq7CL/V1qgQJYniNuULREDbXIOtPSBgcF1rkjHYzdwMXbnc+qvLWdQp8+CxI
1iFEzjffKa7BNWsly7/LBdzPoWH5g+nckypQ7qzCVnCTTXz0udmAtwiigHI9umoJ
ji2/sU5zvVIUnSKQomMfec7GXtp7TSPQTpFUur76wMjm+TMta5g3utIn7Ypv3RzQ
dubgezI+oED1Eoz67MUWiozRmKunn1XJxn5b9XHZzdEQ/WGLOMrzq4yRLGNgiVc/
eC02WzDOHNK0mrr37HO0RCDBzszDQ67Uz6IohNBsPY04xc+5kCogn9Wcc7NKmf/5
DAKo/d+ep+RK79scsKd1H3lI3rfyMYCqoaN+rALTYYCP0NOFU1MdGoARRj9eRiCf
k2aa5fLFqi7D9nCissYYD8hVwhT3bfBV/NAXmIx+LJUxWucD65iSS4rH1HlXI59I
ev8gABf9KeD1Ia2jQOoQcQTkmDn295v2R1lIuiMlIFBdP469AWKR19BCAIrer53H
aXUMotxX7ooK/hwO18Qj4PKrVZSGFKkzNOXs2okgOQD38OJlSvy5C61BXyey+Zq8
Sf8sihraU5VsiJb7SZ+stgPTktZfjowkutwJVcxVqB5WMQFUjQ6zKAY2IIKQ7IgH
ZGHR5r3ptooOOfxQkYAQ7Wg2bdH/yryhVLA0CV0+Egd1d1b90jinMUyELrAwbPjD
Nu0QIKZ5ktM05Hw3jZXHRmqJdmrSwm6/mk4kfotTSfYaCqGciHr53mEmktJDjxCW
8n+wFcShocCdyvAPCOIFJEXwLIThGaC/eCfyiCVrYxdXhpg+Ma2hycoEGnqK2gsS
BIJkUrD+nwtPnZ769+/TEPh4unao0ygIHSwGjBbpbHvU+Fjn6bpXawhflFrklCCD
H3w95/ANNZ3mt15rh38orMaVpVf8jiCnz/473W4bNE/aZ+oARRrAAR4bQTQmeAth
Zl8DdI19FOC3GTvKaHZ6Ezs2DKJlxsR7m3MbDlZviSUuH5pyrZuenqbGd+HazzeE
CQSngTIT7kTYE6hZxTKACCxdaT+QxUPrZ5sbgFfL6L8/eyPGgF+8MTZBIJxKnF1b
Vl+dyZzRYj7Fk/8M13TE6pikMHRGv6jp6M3wJyxpGqZsrJnznye6gxB/HM82KWtB
1Jcr/3+vA9JJJ3OFNmxZaX92sjjiWT5vp6b6we6n/79xcE7Y1R9OI0WiwYzZJHqS
nMAtyAsrmkjbUYf1sPOK0sUkNTOdmYIGOPncsLWotImW/2GR5jL/HOV486sqs/2A
udmwFCcZcu+5RyGH1Ge2qQWoaMp/8PxvMmxk110bZBswQ5rMY+zrfjGvGNjc4WQk
TwBMEksQaPcrCoCk0hUaV+9+Y87MirvEy8VUkaLwjW+8U+XsLhSLhlPcoPPuo0qa
JK42CHuVIb9kKYOMpN2rqHpXC2Ar/fwY5cNFwj/9pOpzf/dnxVJlGt0FzEtGgEF0
NN4CWRX1uestbp6o4Sl+qqgGHkWNJG6039ALC4Y4zaMw05gii5ckNw1GSNagtYuS
vlvTO1dSy6mtFwQ4EjmxAjB/IvY5Pxge+HyhxuW24HPlSFLFi1xEwCjd4rPVMGtJ
ZrN+YlXoAEXXG1wozjCKartI1mCR1Cx1OYYgnG6Y7b8LNdGntmIwnBSpH59LBr7B
Nran8LRq58RxebIFruaXMK4AzhnpDa1MK3F7ycnc4LJcpje9cZR/exddAElasQaR
0F70vjORoKer/AZ80pbxWZu/A3yfDTtEM6iIyY4NdKsnZ3eO34K6zw5QGUL7hCWT
BGrtppAO26oSJx+qvz3YiUy4i49itnoRfThkCh/jo1QzVu9HOdbRkeWrt+RzhlZH
9UJlKGk1RtxREMStYcmo7q6q92kFG2hrmLliM9JZA8Qbeqg31YU6cKgA7NqtUWYJ
N3EOx5gK3relKQ410w6wPX7nwlC9cvm6cRDnqcWEyBfa+BGZE48zvS3H5LnDHTIp
JgGIx1OmOto4FHa3KJcVxCrhm3dZnXXCmpNSc+83rXU0bdd18BSV6ubnmXlmFDdZ
fuJCtaKYHx9nqFBdVl5r7Ho76VoStoU2WYDojKcOhMe3ThmUj+CBFBMbtoI1Ju3d
FKWqBbJ2Oz/S9UJakeAgUhmxm16vdVbakE8hbrZzT+ti2RznYjkg8yI7U1C3cOL5
MmHmzRHmpUYFmrNPnNMaFrnNPYgcQrQXbOuD79PKyt2yqu/C7amayQunbo+qZBqC
63nYWH+3Vsc/ROMx50rSd9qt4uFkwlaybo4btyOAX0rU896blk6zfDqPT8Y0y2Tn
gPqziBrwp/36XXhOS+zH+dy5Vrs14nhgcEsOUityyJLNlEano4lmuq+8UGucx4Dw
pLo4j2h0H/Zyu3bmtajYqDvcT1se+FitQvZuP99e+N0+8dNvHxUQwhYrsxg3fB3b
YZa9v8zFa6ezJhhJXH3ziso8IiAW6lZAhJAHptNIl+w2rp6PTOShgy8rcWXHkmFr
terDUStoWn1wOI6JvzuNzRcy1MahjFW2mICGnVGvZjowhD4qSSHfRb3Gml2iRAZw
SNwMRz/F9hJO/yqM2i2o2zTpB5zR8smSoSyZtTa4uNbHKUiidPOZ0W186d5cVtha
j6+t6SrtTHB0rEgQA+nPearFwZTe9Z/46KLiBfsH1zxRep2zIyR+2Fl0Qr7JmVGF
nA7ZkqbnRO72f7DDqOAhsZn5hT4Y/TPAWYVg9FJh6I2VEyl/VP6vs+v+R31pCE5G
/R9hPv/xrqQ3jQ4ZpGr1HIBR/G/QBmpvxKW5hjeHFpWJ612UaXxR15Xsr02NOisK
zOriyKkzLLxwkvl3DClVjIKDAhrWMsyLS7fB6WmvQm4XTZzdCkZ+Fy3AcBP3TdYU
Ok1wYBI+oHfwSbJ2xp8hvqayPznBgIp5w1fwiwS0e5mkGRZIVtIGVFYnCbbZEF4z
hvitGz3hKLVcXk9NmFUV6ZVtg6ZymrRGzXAImrHohuVf+Z64iZQOxPUrO77AMEiG
HxFjt18cojNMtZg9qGGTtaEIqsVUEh695yQSlW7AAqEr0AOhzCWG6qMNcREL2HOk
F/i9J0d5Z/05+mFHziFLVffXeYtnVecWQpl9a1dvxcl0NHa5Gd3VE1BbPzfWkvqz
pc/6sCejPOENbSoxEOjWTB+/5nhid7x9anRn9Jr6bfaM7jL8ooTlxR41WkIWAXcp
xdRpUtsMxV9vdnLNL3MERWCaBIgTFK99m+oE3ePzo7VJ65sIvkbiVnTCUTUyHmx2
p5boMcd5nQ3yghDzeKMeJdzkY4cHNoxeKYqP9OkKZT6wNi77hmPgrqzXeSwqOmfF
mrVWywS9ASmZwYAwv8TbY+VWjlS43hmtAdpSFEF9zjWvq99fVZjFL7wJb5YyOmjT
Bgrrp9cCEoVXnF/iFVQ6k0JvY58Caxdct7SppgftWzCSebBDBjnHTFpx9/Td5dyB
4JfPjon1jC56B8XPF/d2czJKev79Ounht7mkGkOzIBttL5ApgNt86+/wE8AbZZna
x//mCSivOu7Fo0EaZLU9Znv5K8vZYmpeEPr7gVXyhrGCbPz1wnDmlHoGroiPinm3
GWqeY0w0p8BnGTc/z5IVuqEcJ4OwYtixgph5SSicu1/rytpw6aW7Q6HU2a1XjEeJ
ahiIlnaJffDVPfC4+9pW2Me+U2Tb4GbCn2tEauWkDphLHy+ANcJBkcjmSXnTFyPj
5h7RAoCua5Lch5riohS8K3+O3X8Q0MwwFlOGtkuMLVzHoZ5UBgJrnKwuwVEawaER
MU9p/Ov0e9eeDaLTJiVJ405+/b4Svz8xSVflX5dkwFhtY//lxJYT2ulyAwiGizMo
mlOP6YA/27YRBV8xmH9zzGHuzMacpNH4qLF3bAUIK6is6H4BCaVApMXLbkT7n2Vk
7k19/w68mX086END/qnqjRDox+6WV8XQihYKUYd5G1ZoOeCGwL++wPGYjKycFTjH
aT9XR8gq70jTZ0YeIPmkeM2RJ2/TailLl1zRz8mpAb0PnNQMTcch9Orvsid6cG7q
10wZIQ/1CRmOuhGYzV+sWpuqEEUq4DiiPnclr1G6ZR8wvrsZ6RNDXQ0GbEZctPb9
VVWZf8xwxVa3PPO3JE1y+CRmwIGqV6YuHc0pg/qC7bScdj503/PUzrukAvTLkQaS
Wsr1eIE+0t9otH5uokX7mpilUYLf0wHz1FQQIZDs+pcMXACuZatQ3xed0iPOeas+
IIbtKJkT8XN4h+kmfdnQMbuoQBy6WpwgUFioDEKSjdAjtl03qmViuTc23R5FtURX
rxBui8KAbpHX8AKXKlr4AkJO4oNv8BorrGBq/7dKNWMBa6iVPpuOBDCq8hjmd8gi
MunuT0UMbDMn6ThECLTMTiawcv4wUdl7Gv473q6PJUQDYd2a3Vp/oj9K3l7Iew6B
2fBokFy8uP3FCfGIIbO/G+CrZfsSU3FWtG2poNqPfyIEVdeFT7cbo0kHVXF/ZEjQ
Z1lyD2CK9JM5YyxiFv20wJ5fo1RGaXnNjV4Fh/b0uy/czYH8eFWkni8CdT8sKlCD
Og8tbdMCsEjLLvBXf5mSjkkJn4xc2++LK1FajfxpIyQvfyo0wM0lpcCmdx8lzW4C
UncdJOL9Zqm5/20Hf2jPbZkrsbVQuBr8BvpBBbF06zwJxe3NJnZgcFrja3Jsj2v0
YQZH9A/RbKIINxUEASLrxDPqjTXRtCYmd6iOIw7c0S4Z85dWs9khnmoVL8gW1wDy
w/MURPpydKzj6CAj7oy31D0BXmaR/Sfag9u0IW/2VPysB7z2DKcBMjooDUvCdqBW
neganmNDejRTeTihIMPDiQXHoni4U/ONqubSZI/G9bKEmOFR1KMAMT5MER151u6H
Harix92abRtHEexZIPGhdoWfC0tTPKqbwK30Z0nDwBcZwsTXXecE7doTum9zZRtH
0ZR4cLCDmmCHDcwuo6jrxmzWSDYEiwXy6cWeDOPPIvn0T/h+4f32Pxx6AwBzfEie
pp6LW4mRC9ONhPECNPl6BX0NywVS5KZHYL1NEhZmswo3AJTAHEYuT4CQaQTJVyha
LyrulPrq219LUlsLpIdEqkjLoVlnPCqwUmTxNk7xhczzrqTFFLelXJ0EjLBKSRUy
Wwvm5oPdHVJdhSu8LhPA92lmJkDoLGiBZ4I5Psb+U0RqRYpkmWO3FI1AXAlEblCG
C+wftcFurgJJ0UYY8YPiu1ITTAiVjtnLzIgIRGEn/OfhdYnJegBlGQMZxy1+2rYe
d7y7xADzdA5lhX7UC7pBkp87ZO9uUrsY5wY/wmcV9KZPv0KkRk5WMqAwJmMqX3Ba
pft8rkG8wvUzzErJzh1rA9TILQBoiTRuU6BmkrN5QAOWdKtisStipCRHqcYB7XSD
tOfkHH5VZ6I4B06KcmOIZow97yVqQQCp+QWyH1jXsvCZW3kQFsgdyrCe1scPviH4
ONDjrLZ6oGOcfNF+WcML5fvM3HaWAilWCj5WfGJvk0xzDMu58sfZmF0iq/aowK5k
9nTd6tr/+oAfBxPwUwMNwyKNasmomfYboG5bA+hZXIiTgjdNUPlOd9RPORAr4SbR
DHr5fGzgxoQ9xX1b/LT03LmVuMk6q8Uzz5rQrfCGnHfsYgM1KAVVztS1fhYvZ1KU
EvftPVXf7KDFgBiI2rE/xFQMdbL4Yp4CcSDrZdTT6+a/ADtFTeNLUUJwLAupL3jK
jMEU2TKKIcjtNqGK+btj0++3ahoImoJ+OoHtdS/da4/bFVNUsFeF6pi6msMxEPVI
9J2kKcSiMLMlh+ZRHEI67O01JEKir3zMsNHiZI96uizF1hQFnPXNJq5eK71kuRlz
ROLs8336MB//vjKeswBjYOAAClb23QAm0PoBv7PYQVfG0cj4XoNgY8aDhQE8ynO6
CBok3DAhqkjD6tOi7jgjOskkuCASgi+DPYsMF2U/bnKOYPlM02BHfXKdISukc/lz
KMw5EZIyPfMb0Q+4iw9YXdG0QFM16jy/ugFthZnJZQiB+VVvrVF28iznNS5xsQAK
jKkGUjBD9/Uphnl9QMrnP1vGlDKzI8tNgqgvlKLcDZNgE9/GTrex+Nirlrt9UvG4
nEovVFy1W1iDxb9aiTCBfQbNoVvUXVy3v8QyDeSZh3AT6WiFyeREuPocHXyj01lt
4ICcQpeBFBcZmyhlrS4MZvGd/lJ/J9OKyqJ+LsMUyMjETCqYatrznqLld6CFqrdh
8Z2lFtv6GGGkjI53ZhberFBt4cB7ULsOcxvvMLPbUWynhNFx/5+jSOUWlavNbvX5
nCS7MtLdNaZqR7VRmtAeu4/myZ9WcbXs9YwgXSL5L3oqpFZq3uW/BIMxAix5mlF3
oXquaXdN3QthoON+y6C8T3UKukIIO4wHCD8sVDbUFWn8/JeC2tVwJRFTnUO40xJb
Q+Wx4p894IncZa2kRtBy6bQDAozD9F1nFbQJOh4MnkNoDMHCm5AmGQ05a3aHaijy
PdLslr8kzH8oQAoBe+w6Xo44bXWBjQvg4FQ7zV9VGXL4SFHktYTPdnBjLobE8Yp2
S0QMfPc043nl4TfzoAWMCGISMPmmOAA1DjYX5MD0Ie+v+bt+v0Oxdrxwv5JLziGE
9bo8lV2xRulJn/6cb7NpVyANCR5Gv+pGwHFejUeMwcTk7gLT7JQkFAqaNI+m+Dfj
vD3IYx12UPuh3txG/gp8sJ7IGD3RQRGfHbZyPIUN92R5enmc2GUGhZK9EcEc1pQk
z7DqPVYLin6mj6txQgQWbFDRUh2k+ZS2/EM++aJ4AIigJO/rGSTnrMgXigDPb+1Q
flby3wsFlin7BVSmgJzuLU6jQnayy+XPVZPviof9CSs+GeL8bo/V1do2YXiVM0tU
suVKdN8vgKyDXm7h2Ne+3tw9TpG2hokVNzSF2UuvwfnpCDT4YKuHug2fCu0f+CZ3
5Si4CPl6fpgR3M3FJONh8ufFiYHpAPlW2HhDQrSc5HdgHkAaEDV4Y0YdGUXVvzeI
pqMuSJSGoRsmvBGgXuhg6b9khEMoK7Bl/4l3uWsLIeqraBi2pAS607/JIypxshnc
xLtBWFcF6QhNkM25fKOoQBJ42+J77oTFa92c9JIT6VVkhp3MlD5chtTNc7ubGgzl
8UNwO/ojf9Yex658I3ksLQxfNCza2tiBg78vlK/HQT6on85ZNj2Gap5YcwlEr5PN
cB7zcpNlJ5Fkhrm/JJx0kpUflluzZgCKgvn377otAvg5oNwnyaYNagKwYElYIKK8
6AohW4qWCrDE/jDg5JfT1ELftFKqsRpN04wkkApTKRGBfAUfnSMWxuq5kRFiP3yP
HBrf6kFBKErClNMuXSmSFJaMPCkV90CZlYu4NMCGNWyFZsiJYuN5bQM2F7/plPD2
bjyXVwyw2YkJwUaOu9coLCPmLRO7SCzDaAa5zbPhrATXrg1A72DPGHYkbKs7/3Hs
fH14lQWYubUn/o1f3GvHJwSaxhSGwDiPnOQOE+eQH9OGrkerJc85335j2bzTxriD
cqoIduV+HGZq9k+jdwE1VaII6VIdxqvq6kyBywF88tkVQ92VN23wvTPMXnWZIlE6
ccg2NVPuv3sniC0kw7OuKzUy7aSMmeqXOYGq47qCRcvZTXB8FJqhiSpDeyhSYMA+
IrXOKBCPBYuo/OiP9DMtvNdwyamX2OH+z15kysCqswZJE1JtYFHxUOg5a3mEJNT7
S2CvXvwVZiepgjcLfV+f2H78u6I+hP57EoFnnzVVK0b+KQHsVNI1Ahb1s4/r8cMO
sRGhfD9d3GJPHxrpN2J14mGYRd8esKaGOcQ7FeLfTlrqgM4drnciHwJyCafypcWR
J5YqPsNhCOL//xCrgFHcmstFRa4qqiZ1CXRaqc1tRE1CBn5Sdh5vC3HfjboBZnCU
c5jJOS615rizn/Y2j3yoB3sARsWDAoa2VB4YfpecabQ5t2Z2VXBCQY+OdFCLmqq5
EylHW25KfP7d4dajh9bZGGueDW/esjF06HHsmxH5zHC3ty85/K94fJuCBOfTRvLD
obxgqCyuU2ObblPGh3kzvrj+0tA1/MdTdr5IdDwttXf4yxBz57fHo24XkZ1JCjYY
uUjhwnHr2IyDRHbs5LjOWP636qG2cOpXyAmK4DNVxRJotwBSHgGj6zmOtFIoCBtc
/sEyqo8d+eG1LvpPwejkK1FsEwZza2zs42TFf18rk06ur37oR69C5vBmwWYQFZL8
Au16IXd+kZQNAAktAeremTKZKObZhdGxy6zS4/6RfmlzQUsLEIE14WAP4Q5psUkJ
BAg6Kbkv6NW+WuTK5GvGAKuVU7DUxga1bsgxNG9Ef9NnZMm5vfVxKFGzmOeUg2ck
82qA1iJdSxq3j97ar0eQ71MOsOYVQFMdD/IPI41hLoh5f/wrMP3cJ5JcCzO1qdKh
MoogAy6iNrIilcKYwolv/t7jti3lV2RIRZOpx9S567/SGYY3iDhb8lPeye1v4KC+
PWVr6a1j5RU3shjLR85YwZS6m2C6seo4wAiAJvzHAvQKC2kd+OoKTdb9tDPVB3Sg
CG7ZhrbXJ6+iOjGcmNswYOu9pcorkSodl7KCGRfRn+9r5C7KnvQQl+YRRCRpdHvP
BRcfJsZFfr7jtrpF/3Etzq4qH/HtE3QME7uTz2Z4FCotHbby6vj8UpB6lkaU1U65
6JF4me1GCBGO0PgiN/Sjr1Y1SuVmrsgYVBODjX1AhjWEvicUNK1GJKkZMxkSgtge
LTggjZixOqgJIstMV/rTf3w13Gn1Ltc+wvVyCeuFoI3xoAqJkXj9d6J1iOYbruB+
UTPj1yfps0CtfFLGsgUtlLwY7FXJEnweKZmw4Nrg/ibylOe+rlswSV0vvbe4PKDj
xMVQNg330BOE/7qs4sPzAfqDuBiZ1yvOEF/39DSCpA/F9xVyuYNZBGU4bLgntTN7
uqxQHANXmmXJu15iyQqOqY7FG63pipNth9QV2my+9WXx9aBKJMmdQRzFY0ihZ+ct
2eeI4MV05iRZoL8AiUNaZOIdvspyGLJIx3jf0pj7AMLU4gn+R10TkOfyL611mIDr
L0G7fYACNNnQ+F6WVSzLfBAPc9i4gHmzCBDYttT4+KHHJB+hwEdfGJjtQgw+j6yi
rzqvoFpLXdo+p0ZtLE/l4NyemUuLULQo0uAnZxV4/JRsJW0fHnkTvnKBVSU3w9YB
/LJh4OuLtyfp55WHzZD8s/d/HEp1//0haTTscoLfXm10HgaquZCCyHDnczCytfYy
yiNUWuU1PF/LYQ3aZiN8ZgvWOvEi014XlqG6W9qCuyxoLI2UzH0H331pqFih7wYR
D+ZcUE9AWkQg9g7/sp+GiQJBoDeKRA+Xpl1aBW7AAke8VvX5waqEQ3iu5LN0ZUU2
IvhFAL+skSNkZgEdGHMk9qemRGsPwUrWE81yeqN0k4K5p3J4yTSyGWx4XbENYnlO
ysEd1rrGrNzzh1pY4A/R02xLhFtCBZ9NeILJ/T+dkVS+vLJHzRxllxRH25Bz8Isw
M3SZhMpRuCoUwqy/BfQI1T6UBH2Kef/H/J5kWj4r1UJTKandD/Z/1+dfdvciS8fI
5fJ2pow22+mnFBXsYLBvYEqmmKCJAZF6Ht2BI6IVhZEzPQjHs8+Ezc4LivHERoBs
RSY5QFtk1de073zcB8n9p4QB0GprIBpRaB/7FldfND2ORuyN9kXIW/ylNZTFUzGk
dmevXDSL4Nux/5WPOXi0f3I4jc0m4AaE3vFgD/X8iZVteNx1TMatwv+nZrtnLyJE
YWL4sCRgXzqZ2QL+1fFpDWA6d4EF12tg3xBNE448XD2+cV/jSVPQhhCeReX+zlDu
rc+JVm6n0DHNiz3KUaTeDMY6aC5sbygJECn2lb6WnD57Hd3r78HsSu7eaj/qtV+B
nJtLMpZzbRGsSz5+DVt+9jYPMcqQFvHxPEnnFzYpLrfUoZ05+SznSDDwV2z9x6VL
9t6zk80mAa8mxUG5KvmYJhta9qYR7JSf1jXAlSkv+02H9VwKDSIy5cxgPAMYpxHq
ijelnoHxFRTNmh/Q5CqX7RcPLgH4QF/He86SPRjpKr1ZzIbjds5DS9SvdbbzUIsj
RmZ2L4+BChNSbfp+drx73ZvctUgmWF/Jzd5gMxGNdSfklHErl72+3WtmYcVv0RBx
6CdJlJ25BRS5EU9VF+kMlwphjdMuNTQUk4WVR0APt61lEEahlCIrFj3RdlGbUabL
n0cavEmx1dBDn5GB2N3NhKX5fiaTewvmtC/4cVEnacFXxHTYX72diuwe8X2OhA40
mUotLvSvYOqhdKGTuSXikYKxnUexYciw71W5Pm4h1t+249Gj74vLj6wsvXxDEZD/
O2NOxciLR1j8e/FORO/NSTB8vy52Qf39GdJ/uu6YuYsRuO6fG3XTj3Gyr0GltkaQ
deiRroIL2POzJ8tB7QMs1w9RvmkqaHRfdgn9klQN8XzcaDzDkF5FRHdGnklpCPSQ
62kxN99fjD0XbQYT1W9W3zpbepsMV7Rj/jPp4yW/nISb+LVHGuK9x7gAUMWv5Pgb
4NG9gtifEPHr4iLq81mTWCcVXpMFgrf19P0qDGIDa75JNdxuawTyDcCxAiesmeQ1
ExTeMX+DBqObX6rgcjlsjd02zSrolHGpGWEn0DG5UzJ5c6DfYBbQfZtN1Q3JxWR0
xKEE1VlxmhVO35rSgTTYvL2nZWwKRGugk+LebB0XZicVqrcHC7xF8L2RS3ZusDTI
TV+PWY9+35TEaWqgoEY8BsB7fWXvulAezWTSplBDwIuYDVv6dBbZSuNg86PQpa5Q
SjPQfjGhLeJ/BTuqnwLnRjZ6pqdASMJIioPvgwfkjuKWwpSF83vpm0WVbBeLRtXx
U49WfbyoyHZfhoUW4QDdBsd4l1TmMA0XYN1kENHCJEtjMOK5w0WhtxmypYBjjgTu
ompwAuxqt3GHeyozDlnf9k7LsHA2rkMvHSPTxPpXLEP8yk8sgLdtHhW5tSRequH9
nLZCUJ93R+nGfl1bVfPBsGAGfnLO2xvWOvFDxR95H/RiBESSh26FCbM9OHGEEIQY
L9V1YZbAjmdUxFtbUKNtdd3yN8aWx5hSRehXl9bcO92sfnE/EHq1tPZstIBVZkMf
vNAHGu3zt5+2491BpMx79VYvEcgl6EMNx6d86ye1UubcMHZ8PUZVxJX/Nx9KHVRx
tiSt6p+BOE+NkgCsbTEtQCKzVhKg9REG9ViucXrPtwnZGXblqoJ78r59VNv0Lsn0
DyZL1vsXUAaGQ2ttrV12otENQKXG5lNR8h1aRTL2i95I3GqPpWXhtRb9Lw4hu8BY
kOyyOn3DTRJC+OhIwaUKF4L2V0ijfcgr8jMQrEbI6gXs6zbr3Sxs6ajJqsAKvAeO
moe8WjEq1Wo3nTHpGx95u7VhfpM7ZUn+Ik3CxPiOt7/i3atUhPL34+LwzoVAdbg5
ijGyi3M9h+6Ajb3OFSVb6Y7ctiwNmq7UR8LbnyoQWbdq2IoePb2AQUZ66ANbgm5U
fJuXYWvOXydvt5tJdyjT/uKkQ1fawGkr/cv/nqedyvkLTkzYNtI9hxsE91su3F/Z
RhG1tn54p7ZfxKdyYnQD2I4DWHJhYtocwNaQhbpWtRSXahnnciNYQVJ4SYm/CbQj
AydKDXIrgtAby6cvCVrMT0i7zdRi1CYb+1IfadaYQ7ybma9UG1mfs9mtcfzVWdIZ
VxPvIHNnOA3IjiOADxL63TVqutnoi4v4Cz+h4rIpZTQ3p4jHInQe/rl04nUTs9DM
qvAAsfiqbmS5sLsqpYaKVFExMTvsFMPWCUELv1pzm9DhnxEdJEb9zN/vW5i3pkg8
ps8iMFbstSUd8cnhQzDS3rboTP7XwnxS5TANDqEbTSSK44Pu9fD6l/vKTOQy+4AQ
ceWI2+j/AcupTiauvtr3ZJZ7rZ47EN0yddjpsKgec9fBI2CJ1VzE864EFwdo4CV0
3bCbtJIo5un2XWUo43xeFEfW20+JkJqiZuyMzQZxgKrYLYNPyMvrGwQ2n9FDzOI2
+5lNyuWoCdbi2wWnvV/a9QbfSsqoDTY2LWWdV1jxNj1QLunQhZdMS+55UAeagqox
28DdxnK0MUGqBkQgOHRxAT1DDtXrBrU5vnH45f7gH6QljDKycZa6GTeLDbe6bj+k
Tk1JpA+c38yKvAjwKdW0FHdimKL0K2LlGfqjwgvuiuGP+A+3zT3r+161+IjWoL3h
hctPyz/dQi99nhMiMKx1Sg==
`protect END_PROTECTED
