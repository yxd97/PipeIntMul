`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEtdgqrOEmGoFJ9X8HubXq0mBmDYR9X+IOxzMYwI+ZvBhXc95+kbDBovGe4ZUmi/
8CxgaVK0uoC67ezpesCc9nwCboNrS20kqITk0gycqifB0zzhj1YcrZ13xQH0r6V5
u+rJA4imt4zPX9XKYwK8prNoyfGrYfrkjX4LrB74Uhj5OzmeDx1UaUch2wJPPUbC
yriEEWp3U14P7/DohiLvawytD34gKpOKhNQojHZ8sPwmlf/X7QXD335UlzUMsU72
CorrR1rv3dX1wp37xWN7YQf94avlZAQriWDEDh9o86JwlFzcTPG2lfybr6Ydx2Ht
et1Dm9B06KkBmoD5Z6j02xdl/LR78STcJ5CSSaIkzz3oTAnhm89IJUdlzJDXgq0Q
ldCxt0BdYFzRvADvMJXARRcKSa2QqTBtseFPngZUxANDUMnHAnm0YeXXIjDiRQWN
6gJGklE0GbJ0Qh45e8TD9py/5jotOClQ2FXoqh5BKcEtDDvzJEGU0R5LSJZOLq8S
PGLK73zMuZSDGUMHWExvhDMK8L+mj2GHME60QDa/6M4mYAastrnib4rKbo00b954
Lc4DdmS7XNYSl08FsSQBN7rVc1exe01awrSYOamxxy7NpFrdvmm8Ss3XrOCt9cfC
3GIP1BoCNMkqnzxJpofE5VqRPNAzAA8aB/olTUJbR1oW3qNlATV58hNYaY7x1k5Y
f6iS6GN3lZv0xtltSy/GLFEk1XWzbYiMZRI09LIEB3Jnu7z5plGBW3vS7+8dlUwO
0QUH/c+JvE+psLJY9tnHgzRsKN08WEUEEdw7kn6sCW47wcq0RLzEzC+EmiR+VxLn
LcNe8S3p4V29Yd4lSzbiArEE5caDoWD5vIvMHbE3/6n6X1x7TPlZ7dyNDbymopye
wZv+6dJzXWb1byFtN4t16lnnplKTQG3jUtpYlHzIpO2sUegjlTIuncpZU8GxW+YU
yObenv+QKAXqByCFVk0H2PvYREfuucZxPFXjFNrlcF3e9B7H5VM656Zces6p7ky2
`protect END_PROTECTED
