`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DawT9wx8a9YuWe4whFQFZw4UluKeZe8A1SBI6fqeHh1ElPe+acXd8qGT7Pf9qE9n
iqZb3f4m+w6rs40v6T8tmPxwJDePZUZsHWZVOPSjo3lzoswQM+RI7J/UBBU1P124
xlXYshYdgpgi+wYDkbaNrHbVQsOfC/OD1tDUKtWsn10zkmB1uKzdWh5zMh+9JDWf
lFarQXNEAb0mpIaCImrkGa40ULozM10HSMfnwf975uunNkHU8YLcbLj+VJyfSKaZ
2iyXuwRQeGiXLRP8xU9sKYlUTS6ACCBbdpvGnQge2G7K12xtP62ViIPLjtH2Av5k
GhKpdmfWVDJ35y0SqJw9GR5FpEfZhv5ltdrcvd1H7eIS8p2S2Qy0x3rRiTf+9EMQ
5Q5Ru4Yw1Q0XLz+Vs07KHKN/U24GCQqWC256/i2Um5oS76qrbK/whmBq70vYqaNW
tdUjvx+uZvgu7M0mL32lCgLgMbdnqB5tILsDXBHzMXKaumf5NX0SJ3w5LIZx6r4x
USkSJV8poF8lI1Ls9mHoCB+z195VNQllyvoyftRFD14yxaAmVZ1Vosxt8vmYse+Y
fepmIsMdRWeX22n+Rq0a8yZblSxvvIsJwGsUnrX7253WhuER2R0IG3AMHzU8uuwG
kveg3QZhE71T6+1CioZJyppVdYVG+zsaQj/y+kTWuxVueX2SobRKue7Z5sW9op/n
j1hB6jhMt4k6HGE3tEZK/VnEeYsnLNcMDgw0lR2Mq2r6eq5W/3nBHs8F2vFWVzX1
SKEAbSGjFrYIjb26kiES0g==
`protect END_PROTECTED
