`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+MjM8K0eLLKXJBUOq3OCB9BvP/4aelrjr6psvB1Po2V6wsS95CLmjMP4NyKgBy2+
6cFL6qofOjQtboweskdLN0FRrg/uAwn2rSzmZBjcM94pXSsPmco3qePjF3xHgpeN
IPfmLUT8cBS+y3NaYG3PaXWi89hmXWPeRXW6N6GhWIHPxvCmNveN4aICG/pYp4vS
RAd11T2aFYZlMUXacmuQwgVDOv9NhwbbaCy/B2Ch9h5vjtnwTaX6ykNsESQ7v7d6
tp2IfO/enATzlmWYd4CQRUWzM0MKzTPaD4qGV9M4V1AbByopcWIotWPfvhdhY1Y+
sST+L8eTqsyLXRv7WcP+aw==
`protect END_PROTECTED
