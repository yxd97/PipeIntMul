`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Akqt4GJnUbMXxgr0/UnHk/jHf0B4iuMXoo71TbLjxVJEeOEvhdwwk6gCI+n06mRu
B8Yost7ciOz34ixSwKn5rx742wtnfxlGx4BlfV8lqirUso1+KoR1Gzg7+55HVUhJ
ao06IqBJgxgw3Am5oJSwWxGwp/doX3nn0Z7ndE267zTlRLm1tNdPwBbRxdUOwQCx
sSBoGHZzXCbvWK+dgHlTqo0f+ZNjTvKCN3TsAzq+DUDJ5fuLs3oxJ9frMncKJ8gU
jFE40wAUeFuXIqipb98JD3X1DvEoM+zTrpd29vMqZ9K9kOCMo9e4ZFBN0MDtQyj2
FhGvpwfTXjTHodJr1oWl558dfEwCUzVqpRHjYWvezgLTqM0gfA9O4RVIE2cieHlV
RRdDPQKdfWwhgMtvxG1E9QHfFIcE6sFTwwos1cEdeqi0GWyRq/rq6xxU1izUT2xL
nScM9rtGBRZ+eMuEwzWiM4EhGYg7htQuxTeBFLRfmxmrGXTSXmLq2+SH/bSEqUE5
cj+KUtMd/7YbpkUbCDnnCLoEPa04vfQSHfOUINIX1lQs8FC7cRQiDRJPehXroCpC
cJ7xpeEAe059d/zWD44+mmQweL7F4KsUj8OsQg/OWw1OBKfVkp7XCqx/7wFZERyY
dCHGhb5qa4OiqteHMyLbrr4KSbTnYxgAQtFYfwsl+CE=
`protect END_PROTECTED
