`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjgOoZGflvQ89SLLWdV9VHCVk00x1HoozM6aqhoCHamPqCHVCqRoTLzXvrMOVTr0
mckVLy1uUVD+TFz4+uv97YlOOPdh7FcnjU5NAfYj9WZ3sVwLb44vKJWuTGajmITq
oILcxirKNudUnVfoU+yuC8bFnsHLvy68Mp+N44pbeCEX+eWAMkXVqMN25ZAmNocQ
J/TrgCh65JjUbdpw9mwJMS6CyhyFWMjdVk6XSg9KUFa4/2tJptPnTsrkBdah0LfR
aLM6rtDsR9IPziSuhFQV5DSj54jZsTJeQ4Ui5O2NIlymsOB/E4PcGRGdzm3+6mau
/B3zRMMRluiFN5/saCJnZHofSGPekncv2p1BWU3JgWxY58hhPgaZUvs2L7pRbf+F
jiWbBDSD5bfMTBQbrEfS61RjrH28bpbs1CA+zpM/nqc=
`protect END_PROTECTED
