`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBatyhwKG+VTA7jebRPniZY0FTkpR5Akb02pwjJGKfiCgK/lQWvoLet0yadD4xfh
DH6hcO++bTeIKLgRYzHD852hU2yzGbdDKTZfKE1luJJfW3t9IxOapnSHCd1d8jcc
1Ab8UhXyXf9Yn38TsotsHt5JsVPQWYJcFSD/5ZjvRH0Hrk+KDxTgcFGvQ2H92/U4
0CWlCFLKNxwBL0vj6Ol87BVxtu5RUWTF0rY3/AQB+Ks9fdAgcCMJ5lPYRczlGERa
7YY81FAx9K9/P0yc+37dn+FSUbyVOVXyyzMJy8APQy1CsIDjW6PXsqJyUlbgSqsY
y99JuSmi8SaXZzu5dqKLI79nokjAX6z8gF9fRKwqffsR1A1ka+nfeRrrnEtGNy/7
FaG+yV8gd+ds1/cKPShSKQ==
`protect END_PROTECTED
