`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBeAGkb+3NI4NEZnX/z7jhzTyW0jm6ANojWqlftrJB5qIWVH5HAb3udIjIVAimCU
S0XoAv9ura+OdmbZfroKvMNagw14c4c6F1ULloxcqUCQC4QH2Ub5jgyVql8q8dD+
cgALkPXQFFRkguEgZsRw6aRR5X0bD7ABPaCKptL5y+qaILOI4I9MrweJhKf4Mzid
Nt85TFNX/pKJGL4ZpK1PrDUNS60S35X2aKKUYG/wvx29omuCsLYbsD+pgh/77EDp
/tX0qTLiAMHDzlOUAMudVtoDABYniKLLg7MYwEFDdonJbmRohk6nfJkv51mRW/ny
`protect END_PROTECTED
