`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Vl4xm1JG/iGIUqHdn5Zhwn1L6K6KPal5VPAt5Ywh5xBN1o8Lrvz9J2BkyxDc7WG
eKh74iFXIQJYC4f8GaZ29nCbvmTLyTNt6IXSgS9glhGr1V4oJDpDvvHBANsPct6K
9HSLQmk740JHrLR3TbZee7d0AvBvG66PbCtLD3r2Ga1wAj+VE35s1UVkJObHICx0
9iuBPwwLWDKr+QcFVACr10Tk3Oqx+Se9VIRVm5oTyEgu5ZHG/35xxFTQ6WzzAGDZ
wA66t7tkXEuU/8amkv+zKIqcPxMB9njbEmzhGgor0UwhN9kaWJuHgNs0PyIAXvee
7CSJG+P8qc8kFgmqtPcE5xyE23TZzgGZF17B17723RwrD1oVOOtPE93uGPm5EBXV
Cyx9xo2PNURf/xV45VMbXmgDkyMsg0a1K1HVBl1NN+w=
`protect END_PROTECTED
