`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rWHUJaueqdOa7+YXACLDMx3Qn931unj1H4hmJW0YBGWoDsJWHMO/kKzJMHfDRuja
R7bbAvBEcnNrZ7coqwEXMxb0Kn5NMDzlllUYb2nTkKsstdKnFX+tBtI3EgMgtcfa
sNiFa3+sATUs7s2er0xZPjrXnMb/yalvGxLnX5qfu9GB4Q2e97FMioOCUt0Fu+gx
45ljHkGc8KU4EYDEVztGu206yUPpSS2C0Zy2LGo4EzHqPbbSVw1xAVcdBN+kJuBm
F/Z/kSIQlAc8tvmD9GZNXrVkqy/Uv0rq8zzmGiolJJePtsZLdHHSPFr9GDPXqqvx
jnNOUt23nHmo5ylZrqCcMeKmPGXmTjsZw9JiAZUQNdk=
`protect END_PROTECTED
