`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EoXebL27K6oAPN9adDN7JC2ynf042IomJAH4A0Te/ZLNFXnf+CJXsyma+GVcIzKY
pskjZIHcRdrjbSzZKYGWULNswP4Vs3OMco6SFllvputCPyGTTFci0ANigRd3ba9P
laEAKpTyn0U6V/zo2iqOakPYzWICW+L9BcZYl1E5WYLqd2xvvqFCAkt8QMQTk0Zu
ks3JVnU9KXhHpweMxDAa90txlXEjdCKYfxjnSNh29htINtq7DWR2HhY2zMTyeROc
8u1ht9xiQ3PENRNjYYgj0tuFj18LGcZeOug+V0eotdtvn4yMt18RL+K1js1ZQHln
sU7lDw5DofJBNnDwudV0oY2r/T6O9tCJFUw3HTgtZl0=
`protect END_PROTECTED
