`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a7dV2Gx0XjcSEHeH8VA11bfYxQqbRkD0xBgI0hH1vQ6YzTViFl1U+ioVLV+zL85W
f6rR14P23OHQXW1x3qRHJ3ey+nb6KVuH5haHva8Xg6nvXzzcTxsmD1PLHiOUQgOd
6QnJxVhCWcuvWaFm+AsXVsqDAN9w8FyaavWbczr2Ca08U7XUS44aQ+qJ386p2WsE
MLQIstUv3b+Kzc0vVC3ozTQgBtTys2jOcaqruePkPGd5Ogy8S4KBoviRSw61AI3D
+zaHWpBfQ4FQGP4tTl+UD700l78EBwCkjgBMBDM/LXR1cy3Leu2XQd9IAAUxSzDI
V0jY+VIJlUfblkuZjUQB2g==
`protect END_PROTECTED
