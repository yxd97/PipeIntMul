`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jOhKkoJ4TlDwE+89DA3yQwIzcRX+iAo5xU9N15wGF0PAZ2sDCxK+6BzqDW4TnyI2
Yxnk/awYTPm5ilXuDsGKU540Z92TfLVEWZJ1liFxmoYpy46xhqaAs/EmzJZQnVip
Q+5+2NFr/Edb0nx8wktRtbwqF3KTBy0puPr8+Pf6G0HmqMvtcA3Hx9BhmWfULWTa
Ap4kM1BgEmHdaYUUfsNyI1f9srtAd0oDBKjlsn9fzClji7PJ1GOV7kkBjza08n4M
/l6qUvH5z2CEwM2b+oJbKJb3wvYcJlinqhrniAp1lAK2lQsWb0w+uYrDNq3P8cUo
GUdNbRwzdSMCax1vXswn66/e7Y2l6jcGtS9g5PFLrdHEfM8r5zjNf2OykuerpAOV
bGelyNGSLDUp3hz79FHfhYqqRHDhUySIHHuOltvnOVG5euGWi7GxEGrOqbPVM0GE
ezWt6drKofAvzPapOznphiaQKQA4DeS1AvimpbjifBs0jRKT67GDPDfaAJ9FJz5y
/pvi1/8jpZUMkCvQUbsbR5fe4IdC6sIhMke1J4WhLSnNhn+WOCgO8mKKj94nlwGI
o+w+wHvSAv3LwSzciL6B0UdE/d5DARlZpBJbW+XMRWT//ECoDv7G3fa3n/i0hYao
36BndFB2Z49u7kucAf56M7WOUHd3NDX2GOH7oswiY61CEuCNeXCjTyU+OyHASJdY
zf4ioRV1RX/J8QsWdrWFrNltHRMCCohnl0DOXVPJ9wv9pgp3/UQ0Us7NpXMBaSyI
GaUc97omx9+8L0NdHPUL37pkzu/GZcFq67Ts6JqZv9amIm4qb239B/s9a7StBt0g
3JFuY4Rb0ADc3KfMNbCoJw==
`protect END_PROTECTED
