`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zb/3Equgvxfgq4m7Rt6dACFSjupHA4bBiZYsrZqdJUXhOiU49g0W5+C18qAMqZX+
j1RQVi336ynMc1OQp1Dl3ARJXF+TPK/KC31W+rKYfpxrQKH/M+LIKgVJKZhHQ4ob
UpC04HH4zrPuG5WIvV7F6lX2iY3nNr5xz6sIHtc4KaNcIcnKBlBi+dmfYj/1mdsx
GY/CchPb+epF7LEzbtSrZSqrNPers3qP/uZsTUO/QWYeJ6hJouXTQ9qAI5OWtnAZ
Wygl0iPDz6t8d//7XT541nAapefGm/5NDhmFQUrmjYZRFGquIF/XG6HuEKDHMYTI
qUaQKOvbiqqtIWJHLS14kpB0pCGQa6uKj+8IySpa+VSvsS85zDhfXwHpZ7/lN28n
Gw1cM6q4Jni9LEnDWjug7a//B8sZX1iPRmx283D+1fpFIKCaeBMVRNonpdXIqNLB
kw6S3H86i0xRBjwASc5DWpA/EYCNridvEdsncX2Gu8oYyPr4TcGymo2K4oBgsrBl
RD/EDVIEPFlKs2lUcZ3K1GvHuTShf5kiQgZPkns6MN/6eyST6xVu5QOcctPV17NS
RcPxPOxrij/sylQ8Wq0osSRbVWgFHBEDP5lzlOJRWQnmrN2GYFJbYuka0IOl2RxX
od/T0fVeE9zL0C+DwAOEHjI4/fbosa96bW6DFKcibcx6/DzvFJ+doceIxMDGHTCE
HsRmSabS/Pu/XyCDl0QeOrtiLLA83wtsky5K21PD/w5UjlxCGNax4+QDAweqvR0d
XQXgGHMZMNrUnHokpicmTTCHh+h07TwddZKka9L+I6FCXIFDgs2sKVC8wC3aK1uF
vSEIiccFP3THDe0dIebj+Xq9t/0vK/ganB3dVjMsoYAOGuVZ35h8RDAmDCUB5H9t
CQFJ8YhG82X1D3LTeenYH0P7Qfxg2UdRALiwA2C0vVLh/dbOytomaZoWdSUzoqhj
0Jq5j6hIRv+9x3yKgDxOvUwGidDwRfqZAZao0iX3tUV1XgUYp+/bSXSINCBaLJqc
lwhttuYdqKXR5bupdqkuf7KtxBE8+8C4g/EDcUll6iHuqaabMTkBIKC9D+l2emk5
dolQYwk9uWiKHikGqpz3EuYaVLpq3P3trBbs2nZBWRSZvSpFy3Zs6p/SdXaU9JTn
nxlJttoQOpxJGME095RdvfDsv6Mp3c2jINjAodyJ7FR3lHN2LZs8oAC6KiM6fiTt
/Em3Ccg6FRlmZY50CRT+xxPj1JqcPVs9KQ+6mwNCKw3In7oshmgo0yJuA1USnUmq
8vSGBWmrvYLQXlwCbGSCTuza6B29RuYFVdyvB0Zn1yj+HZhUq4W45QX//69ZWAdJ
TehEYITlKW5mK1+QlUSrqccCbu94+K890TpgLOHD1DwC2qWFvWQuFHuuyBtcEZAf
BOuWR8tRTb1CGmjR0hD2bspXP3D4Ys8CH9/Ob/rXtx6k7ukAm+EB73szyC9jQPFS
9qgCRTv6qoyrTUMJcaLW7kk+VuFQ2dhp2efwJ/nFQhHc0r73yMMhpvncDSvRLlR1
GrWXqMKbIJE4F8rFmgGmKtPH3f+M6Whw+Ulqt4hEicZ6XwoJb2VTuwZNZ/DmC0qO
X8RecyRHcX+bIGTNPKMj8iJNYhoA9ehchhsQMJyhXJr/ALTZx7L7Mq8V/sabeyko
ySGy0pHakylxqY0flGXWuyMCnuAbLPZdOqCvx0pmklKkaXaNHvKRvmyVmGfRoCmd
1Th1eLlYh+kH/BTCVmqSgL/Td433vFC9zb6DMgT6v6LQjDv0J2InrgSYU609/l97
v92FOZXI3CkuFE8/45anUJ9FPD7E2bWUrVCjSp620dh0yXX9TEmj12CcYRsfQ7yB
Swz8b7g1QJuSplaBxw2kXyda2fRRMs7tp0vQQKqxSJxOvbz4SNKam+Hd5nnbEJw0
oi9L/qFDPbuiG1DYrGscZ8s0Ns9Rad33Zar6MVHvviEmiyWn7Ly3U2bvRzrvruLa
hFkDChM8dEt9tQ21td/zdzZYjVmDzOPOHiTTsK0slwy+ht8cnEI+fCNjtkxMlNu7
CqPGtg51K/B6fx04X8PDKCJ1FmM5KllCcLwgV7P0UvshxNAbhf7gpR2CAYfvEDCp
DBLNQTHRr3/xhRYrSh9fc/ErxSnchb3ta+uvrx3YUd7H41vi4IbebhuyrITfYlCf
IGH2WHzdQD1klp9OFC0LqxJ5o2yzLh1DOxxKEsq8PKl9Du9MWE2ClR8E294JyA36
iXJlrm8UXG9I5ThB7JJFhmxsm0yz9RfakwmdD5FTy0ikOxTuW3/fovwWQRSl+8ki
MGpSz06cxUi4IKz/9HHzcsfKWn9sHEDB/zSuQUx2Sd1opcsOiJuTVH93fxGqRShh
pU1OCOEA6/3Pgi6SKgoE2Ixt78wRYxY7AVZ5Th31LtMgfVVDbBhJ9V0D5sEQM9h4
VHnc7BksNJ8+m9t/6E2e1B/hQUBMEjbg1hGFKc8kANxlSTrzrC/cPtC2EiqC9RTI
mb7LB8O14KMqg3NjH7vWIRuoWPvpTpexChAj3oy6DF5wdMFrQA8YJBmeU/RsNkMl
riMGhREyU0JlY+GjZCZG4x+MG203D+vZmtYXRU8BD3ph65p7vecq6ATU8ycH/rKK
Vpr5Gh0E47GWoT6MFem5gLGRN46zScVRDQ/VbWmkfHMDMZRObxUbGYRXRs3houm5
BcpXQuS8pHwm8FI7WLepTfYFL3C6W+YYraTp4IQngZzkAy+gb8Qm0KKqdn8lJHyr
E9O1g2e2dgg6rXHTFv3G4RgGAG6dM8cN34igtc6krLt8h0aqVZ+zjDTDYuovAlD1
EnyWC7AQV4HYRBur3fIG8BxfN/F+uC6VXH7amObJt3/Fg0xl2ie21Z3rXmyDkPkT
IfHfhoYrvBSmrmvnsohSUU/I8SSifaJnKzm5IcqY+3Vboifmd9wpFedyhTIAsgkk
ckYdRQgAWTPKA9cRTNKtjr8RPpbbPAWr0WHwq5x6hT2ODYaeTbthWGDGt1WJiBIY
x3sL06xAK/1eEy4VUiW528PYbBzak5a/6otLRTHGWzT1e1lJFlov4O5jsd1Y6y2h
v2ne3VMAN0VHvPmUb2h4FV551fzAGTAOGdp/9Zi0PO0I/moCFGgpArhAXSMOgW+Q
59N4u+Zl9l0XoAhzO5B1/TbtWXr6j9Faqq/E00o47rgKMkgYewJMrrwDOlUX09bT
GQEWP/IID4wMM2L06ZdEO63MPVwqJuz3lstanZSw/7GhwI/a34g7B82G/csp1oDN
UzkRIlQUswCPIfpskfDmFhHVrTpGLQLPezrnKGRhyHHlCtHy3Mt8pAYUwACsYVYF
kL4OQDwkkh9K/kdbj+2IBGCNvfNwII3WAQfDKzb2JeNueTClSGN6veymgcIOWMBa
WEygTtKnsIpCMkXX3NL2o9FkJgl5zcneQWfQZCkNWqrtaRVy2/+WYhL8u4XLWczT
fUxYz+etJks3ylBvWmrBYh/8q2jPya67O/gm1o8dXO9uGp2wxdUVUGbjMbyrZEPx
rJa16Qj2zH4ksLQvyDdkFgAQOqW1tciK7/9orBElKIz1GCIiXhAz9PQIuMCA6e6b
tkqOzkrfFI8/+fYCyoVUhrYaRrt9uwIyhuHJ7BgpUFM3WKGhmg3FEMRpXaJ+1Mgg
3f4BgWMDaibYUv39GGTp/msXE4bMVZS7xiXMmhAL5o+FVKUwOTNWpmti+Xwr8KX8
0YCXoQR33G9Ty6cB32bz+1zIeUOzY3U6WwYU8gQonXgez2UCf1H81LKmV+QI1vrc
maEUa0FLvQHC55IN8XWY81wBaCZsZ9mA9XG3kEW8IfNOLBsDnpi62aLcyBdAzZHb
IiQZYxpvv5d1x+NK2Hb0KvQ/HBJ9DXqmcSkptWdfEPAT7iC50YnonSoE8x2iuYZF
63OWR033cpm0SlHhy4sBYETSqmrG3HQsUwMhHhBRc7ByMJl4kh8ya3u13kHzbnfW
lfCP57OrrT1F8KITId5StCgCVYNdHgHelQJOT0QXhj5z94WLCyfR2ja7h41YkxcU
gLwwnXNj9iAgYewhbNPI4P5GDWnFs6sB6W/zvB1BmKYMEJqllHSGff3NoPO/z0ZM
K+E7XYclwzTRKWNIFU3eJNesslq0Hl29KFq2OrsprdI+MiCQ5J6R9vRMOpbjS+ye
i9vP4QdbpQziFHuOsDsSqCVxFH+qbqZEmpvnNbabWbu/VG469ntoJDVCVAkf1Kwo
Jrq0lsQrqGUwYyeoS2OwV3Oloniq7ZBtyPn8+wXmnEEvJtRToY46yc/1KvcVKv28
XTJcBlm5K0ljAHd4olMhALFBosGeSUNnw6jZPPs6GDmPTrV7aVXNz8L03WMkjrxY
ouEdMZMacHA3B3Do3EN4E0OWasA2LDHkSyce292U6jSlH5sBBfz736GCebfzexwK
g+fdK6X7ev1x/bAvzOg83/Q08+fi6fv3/c1NdfZgArEo1KtwpqjLaeMIRF1Car8t
xc3sRLMSNJKB7ArDA+cgg7EMnusDRKU0ospA+F+vzQRxMa5mA1eMSor3/NcaajV5
dD5VfKg4ckJeHxcy2WyrgM8p8opKeMoQi6mEdyX4D27sTT28NcAfHHoSQ5196L70
GJc/PcRIB9kRWgVUfQahUj9eIPBZrFQ+ZxOE3tViwQ34N6epEEmixZYeVlZFCgDL
hYP1BZApnX5Fo2erC4nz42nJyAZvmR6o8OzqTEYH5YoIlu2op3XXbCoMpmLkLc7Y
kiF37EXk3vHnBBL6ztwScaqLt7X9mS9u+uQNYvgSRyeHkggwy1q3mi0NhxLe7NF4
xF2uKa1s1vE800r7mxnb6sCm/PB6GSCu1t9RCklU/IR654niD0g1/sANdlhE1k4C
zTeg41mrDzHNexsE9svGSWTGXv9eOUUYuaIVvJd2VzPryyKH8zuecZmU0h7pRKza
7QZs9gu74iDNHoez4o+jCcdU0VEijy7rnhrR6Z94N2AxfnFSzb/9DAH70VmZ4Gqi
1ohfFkefRrItTP11VoP0rOeAJg6Pu30D9pQ80yOirbPhH3Q0mvmo0l2xBT/g/Nlx
DVj9r8D8ZZJ8uUH5NIh7s5Z68uRycvSjOUPWPYS/FddJ0PD2d93Yhjaix2ck6J6U
D3bPJv3cbCJze1YjiApLRAAyTf8z5uCdRcrCHsvw9ZdxdwtzD71nzyjeoXbfxkbU
KotKTa4IYUAosBXEhV9gVFBchjqzz9PxZX/o1APPthvQo2aJ4T3jAPOdtN7JvdjL
R8rfJUpH1PynPINYW0aqvwVXwNTohuTVAW75BYo0s4aOUlModsk4wtKiPfE2wC3a
hOrnXtKquUtiqb70WwK1a75TQrSSf859BCTnaaDf4ecTw+Rj8cS4SMSHO2jMWAol
EFXt+a45Ns6nwzNthVUVKb8P0Td9VoYTdjNOtltodjTNU3os7jPZnkW0Ms8z7DRU
hOURX27FDHusR4R83rqsxlV2KaJNdw7lBnH9LOvdZ8aaRuZuy9e9vRss3V65Ridc
8HqGxF5t7AaRj23mmv950VAZEs6xvKUBh+doPhFl8gh0DV+nOnR6KsCBL+xQ3RMk
gTs1WT4UqEx9khjFICclRSpI3w/pkwvb5qPMSeRPFTc89++RfLeQ5EThvhNU81y3
B7pnwjz0thbHxA9FnxpMIWAgME9KLso5WjXNov4yKU12QUpLL1wRm7EUoB1sBVmp
xcz5r0W+om9HrueloYlEQWcDfeO4NiciSRKAzJsiE3YGP6rZHiL75P1jNGjsgM5b
LqWjaM2tHnsl0nwQ7ICiDV7AWewp0iUoD3sDXdxNifLT7piIjY4FzYC5zqWkS7j3
t0kB2ZIPHcecTO2vUR7u2rKbucPvkdPX6IDeYqXDqRLyy+Ro7LN98gLFmE8EQq2p
mVIgnojNSCVxA0ncc0+phKIGc7Gl1XBmJv6PnHkpj+dSrWFVapFH+Epevqo0KeIT
KqJUOwwiv1ZQpcD70VcsPsswgefLgaMBSaQEYdv1nXGTmLHkcAW6dLkLqS8oWTG1
KVNzvxSwXL3kb5wznxXfVgw1UiLmuDZO05vvbxhc/4AMCHCMRBS2DL8uY/0n8p+E
56jQ6f9KBUNiUubUxpKgEPBvv3M8izPCWvuWL0MTIjb/t4lVQ/M0GhoY0Y41/TQA
Ay2hQMrv3efdBmTF5dSHUWZWa97UiLZOptKC4NLxRXXg1IWYmrP9Pg57wXJqy8qb
h85b3F3UKxGq6hw4Ues91A588AS68GWRspkt+KZqlbS2BwYPodX8bfk575MTn0k7
8M8M17bvGr++ElpHROzA/Dq3aDAAIuNj5HBevWxd+qUmGqW3tCQ0qB/bW3YUTVCF
E8BjZF0smwUSu3/oKZvfjGFzS3RF4oQnayNjp7UjOGW5YmHGXU54ZoBiGj9mKpdq
qp4ek7hfnixhRYRrJl3L3RyWsKGN4kI6wDk5y3JNezlwjnJwfu5KwalaEX0hB0Lf
HMXaElciGa87JNm9c1vQVHgTuTCL/2ns+Gml+hQCz2ovgqhVpbmp5Qp1VaHpSgF0
jMdunH7UgOtdQ1mgJVKpTnpvuXYmZJmcYyW1Z7PG8KQpItGGRYoQKQ41q2+MngtM
YrJ7GjJmzdj52U4+p8VMAQwktR8MzsIAOD70C1otpCok/ZANbs9yVnZgCkb0bC4r
nh1CUdCrcArDNZ2rO23zWEojUcf6cdIrVjU9PO3NFqlBe84czj/txOki3q04fei5
iGx7CP7n617ODSIq0hH903815mhMc+TWVVwIYh5cO6LpmdHzn6QQzsDTWyS+C8Vu
v0bR4jWocbLyuymf+/XV6Hb4L2kZ1FBMOHE+U1tBcDMiWrTuvTg6lG4eiXfbqccY
damCg/YOvfw3ioVwxKbJ4iYO1wWj/bL60zuT4EdLcx6EV/M3MLiY1dylMB+uLiWw
aFnnGx5wBiM97SoXecoUZLi/ZXvw6dkjDgVspk0QLJjuA78whMXjrXB5rxKUzeTN
cv3/oxjq505e31/FJMZyhRe6C5+CTWA887a5MNm1SZlxG5qLwaKu42iY5ssoWoiU
DguGcvIpRstmCpNt4N2u2Poa0p/j0m8YHudRcJOcQ0eZl27op1y647h3DO5pDukE
bETuSD3bK+Rh80v6Y6B9Z3PX8JPLCCHYrcFr3KSWbCZpaOyhIJ8rHEqfoeHkfbR1
6DKndD3ejVwhuG7xBwGgZdnjHPbYEvhUJK0rcOYPmu1wA7G5TavlPwLwMfIUqfNL
1uxMsoYhL55kv/Hfruc7gFy5O9+aG2WhNryOsA9+n0EZiqNwHwg+cKpgAlh5GEMx
feh2bXyVPZAFPGK9rERUHRzCm12AbnbLesKf8P7TsPGf48Eka9BRvnqZXXcpL9ev
aiWb1brYQ7pMxtPj/8Y5XRdgr9Esp9yQUsncNBpJzoAxbHW2T2U8dYPM0jHlk80l
krkLuROZrCtNq/J7SEN9pBvkwyrZW7xMZPoheh2aT2vfJFRdTKkzpl5aQI8KuTZc
CkEXvSH/ijBVRBn/BGYN11GUhX1YKaPrgLaBarfKj8NR75oTCBpMqNni1YU19Mxa
Iopm6gghN6gt8i96OGhaxa+wLq5YkqnOAj5pQkGhaz/5/f77qdmlSDF2hlzuQuMW
OqthhAKVqhUKDkCx2MeNQKjLtWPwIa69eoVpjGuDvcGJ7JZlwJynkiiWdQCfi6Fb
oYl9Q02tKZ+eB7xTZ6P21ozRbYOObBf+GpxffxPkXrSFBYSwG0qF8PXyrXTXbpbO
lwKFhy/Z+PWMws0Q7CeZRme63bpZKxv2JV/b3LQbLXYVB4OoJ1j7F3iZWPWQD7vI
8CTfM6AVLJoV0nfXAFy0KzNtQt0X9Pc+0VR0vpIQaO6kd8OkqdGNMebhM8t9Tc+z
Pn4IwRsxFi895CxNiRqm56nfPqlWRpZyfFrx/SBl61V0dV11r9OE1FCZ/9biWEsq
yZvvaHX8dG8/TQjcJhLorF+fNZQtqCnXa1W6wSO/COsQa9wmLS0JACJBuC4eJTKH
Q+tH0TAX0HfCNZimx5ao7yMWXLhhl8bUg0X4Sg6pNAUVr6HCWeqBw+ONaPw74nBe
poRxjXOWvsmF+b2+g0m4DdALZDzOWNizaeYqcUVtje1ZeD5Q0yZ8guCmo+aK7OEU
yvcxqQmDAqBttFWW0ZtSQfmMW5gEykmdy/mSP1ooYuJN00PrCeNPryh6/hu2J/GT
WgTmASi4e4NCOCiPoVZixJaokEb4Qotv8SCwkapwh72seIVbzSOyx1WVisxZUvVs
yZOASi9ngwXacdGhelsc2Fj750sSfs4Z5DHBqSZrJkDxKs+pGF1NHrbDl1GwSrcS
dzpTMdaGvzLPLXBTcyahwHvrdtxQ2BIRX9UkkDNdQL/kicvAYQSkwednK3nQn7Xq
GfRAgnsgUem6LENK2nlviuEjBGGzoRE5DEttfWAzdD6kvGvSDt9jYfHYJCpygpOb
hr6Ptb3WphXTrwYEKnxxKahNb1B/8YnaInDhvpRQB77+UDLwJixQsf6BQPuEqgJf
vNDVUU0D4mPVyip9BS+d/jVVXtphAmznoUQl8cbXEhliRQlEHX5X6cfU3coWD2Rj
XBAc4LNLA/ni4UD+wzRafs+zxlcJFJye5PQN0eJl9q5d5Ea0tZSxbKr7Z7H0W5jy
ZPU1r/bZ7GIKv6xhQyQv98gOPB/OWCRY/NTXQoF4eoq9/evZEpFoqz9bwsPaIu6U
g8YXxYprw7K/mh6M83SeqLTujacdfkm3KIaPaF4Me4pxZaDGRe2YVnhUxYujfTet
XFjVhmu+nlaPumD6mjflY3IvHDh9C1ol0XRPgCC4bcdbEl36EhGs2TVE/qBLqBsO
LZ4ibTxJRvkgM/XNqVlMXbmvJh+/wwUediTgfs6ZIEiOdmxOex895LIg2cgq1q9d
tLM3o0yMK5SKRsNpuSxEcYlgIx7vvnCn6jP5c4Wl1Lx+cd8FRf0gnC1M8gXxlnCl
/isTJO0jK0fdfiKZPYaQ+Nc39OoSaVRaFE40zDEaWDCIRKUd6qvmop40Zl3LrMmf
kzNSeemqm5sqiYQ0YS7vrlru/AZyKn3YWbau47RcD7duf7h4ok44W5jRILocpPcl
+Pa2swoCQNcS6aRYjfABWjSyDovxV9Hu88hd4xugs2IMyojuWYyn7PgInmRyFzs9
vEjviGqLQf+VkFaKuEL1KVrxatEIQtYwHdphzddREg/RW0+CoMUdw6VwhBLusOza
V8J9uG6uJ55OLt8uIA5vduZaqRMooXBgLOrf1DOL+ShZ5bkvcqSqbnCkZU4CurP9
7ZIwMBh4z1W641lbS45jjoZSefnujZWLjNOVnBkN7p6SvlbyiE38qflSDjiVghsF
vIfWWvj9UsclLIfbrUluVLJymtxi96WRbBvGuii7imJHHKngla16rRgesQazt+9e
jPKixNCEVuwgI+Njm+3GugezN9+LQU2UjsxBA0gVfFyvceeXaEexJJIhFk/rO3JW
nZBBlCeuv+o6nBlY9MX/3+bn4tCR6MohUS1tClZ30mSATiIc2eiboQ3C6pKU9vLs
N0OXTuH3j0s8/3WBp7A01G0SdurMAt9Ijl7l08HjqI7elYZLr5Tqvkak5dHnq8wc
J4mleHnbfseAN+7IrlcaSRkaMfkVi/JoMP/n71bXcn01ZHsCeQ5Dosjpr4Ti06ZJ
zdos46u2xdiF9/1axAak9XRwyUSJ5oCW2UTSAHfBXNMEvBusJr2HCtg+rUe2Xvv3
HU6vLe4CAyPw7Gd39medSE7u9hriphNq3Qsnw4kxvMOF9ZaZL8u26MCryV/K+AA5
QxKqJxImjr2CdQ9teHARNrT7JPRApREFS5ROKrNglHoURRPIRP02iscs2oLx1Amo
7ZHLM1VCM2iR9EQfQQz2GSWGWhX7p1HZ8NuGYpCzPe5eHsM8CGAIS3OEGKQMHuJz
R+xvRzwVet9vJuf0/j5puVH6Yjyo2lqCib+oKzbo3oDeU9UooojnM5RrqTG+1T/9
zllRvQ5B4FVnt/NCdlmpAeklNOMt7rrJDMB4KaGSgW/pl8el2iNlt8H0rtWYY5kF
yTRRTZ9phZOrhN04lrx7R5qHCwhpLkdrFu2oOIex4xyuvhkk0WrdlnZA7PbPshAb
gLaGYpDz73TOZFt2z0BGuJApjsydZcEPCjS+5+iG/cddjlH/MHMiaxDk8sUEYZWs
lA3482Fy2tD4b6ZmLLiuQWoH2xZP6K1hu+OuzpaIgj7g7672MMkhYPvBJQyZLI5Q
bB0wrUjzWrKWZ2TOHKgFRvX/gpbHvnGiE380IFmdI6kbxRmUST6IRO9f7SU7nV3o
TiJZuZoMD/lWkkAvZQGedcxTMXb4g7zBWwIf5NQjPHPviTQWk4jw2j/WeoYTi793
0DCdbuEA8XJYWtdRXdUCyzKibIoTGWe5Nokz7qXZ0aRCVWcwGufxNv6zpe1bADOB
wT9drX7Ffrg8/mwaENuRiIPr4D/tbUm5nHsL7aLmYwRa30CcR90wDshtGBJUVx9G
4SlRM/j4LiUzUSmHfuL5xbhisTySG0IO7hBXXTZ62Y1dzCInwH6ezvLG/Bl62f6s
s0nWlCq1YTjN7sV3TNAMScbj1Ru7JUEPewdbk8xYvIdn+0m2PoQfeN08r3UqQv7b
Wwl4u3aehntEHSr1ePlkWhKxrFdmLxg2lTxP9ye+r8LhxKv9pCDAC3kE63ijBOPu
APDaql5HPgAJdasYm1t7YO3VEdwIdBSOJYBG1HFatjwk5clEEaQ754C+R+M8gIV+
jLQIaKKAXTEt7ZBVXquVUh3tzVjt0HKsD3URguofYUqWJgvu7V+2ea/7L2Tun/6V
r10PvV1+DWhMJiM2xZED9VCve7/RPplywj5v4V6Uc3Dr16scO7paYAZNnblGn9FJ
5aNXnd7DczgMvGsla20TKHmH4O3dkVQn6DjjPdxGNU5npIyoD7DfuwerWen9oP0p
22Nw8uy/d+OVbpQrPZQ3h+kQcGFCRiqgV8DNC9psZdDzMUlohjeXhsljhg7o4//6
O5vwu2EeROlv3ACumk9FKL2tRt6CtypJjCSmQePjMxsd2Q5oyi6QnOB144hSgSsE
gFSzA4ePtc72lavF4nrhHhS1XhziBCQu3PPhX/0IGUj9GYOYptSZp7AyM6NA60lb
8GBZ2qoUBkqcIsuvLssLUxz+zxc82ZmY6ifkZq9a97oWzA7CkNNa1YrwaXhyzuVr
29MeKGFWhxu70fYyaDkr9OFiwKX6SxXq2juhKRhQLN5fqOqf2MAfBtcTTDh9s8Dw
mATfOAYhWB/wcdY1TSeK02e090kpnoVUM1wthWlyWvxx7OldnD75DepRom7WymmL
B9NEaOjXKUVOCNqrjsQQrtfE/6BmAxuoaTGfpyf9inefgMxdSV9zymMgLRPYzCI0
pRZQatb8ZVUe6vwbxotM8zZjmm5PFh0SWxrfog7QQj3zpd4ndg9kXPmCxk31qxe9
v1srRxgh6mUV5ZrU96jAm0OOtAKY9Q9B+RsQJZHU/8GMIFqjTo3YxRVY2MMeb0vz
TdQ1KbOHBTG0eNNcqdi6nceFRgyOVlZZ00MmPMR5rCpI7pgUFKrE2RZWeJLhlTl/
z4l//A4y4gZvc6mpK/wEyNmYxL7J16D9yOdVT/E2QtxA0r3dXqtQDuhb70igyNVL
unb4xG3yJnNa5BdeMmsPEDj9Zv/uUrHBuq0IL8I7A/+PNS0/otqR7nqhHhPJ2lPb
qik9Lk0N/hzSRBBNRrnvWbRXryj7QrDgIG4IMtuFBxNPC3/UYyR+9TJbQXW4OApT
BgHI2RVu5wnpAIUpMGBnYOe43S/ffASF/fuILyVrjGA1GB+qYZc8c9zk6Gj0c9do
bF/9mASzq49JT06wX7Ze+pkLC89B9Xt92XGKrdqlVhgTToj5qi5iwRG/d8ozPg07
G+2Z3yqWEYpPDzWFQ3JQBPbPU2RrxvOq5lW7vM/BxEVOaNsHdmJrijnDnBPkjfOq
5JvliZcZBXxkCqt5EQyWJdyoyN08Vv4NY9buBP0zp0J2GWpG6/V8dcomPq5ZRCC1
9cp8KEffZOaFbcS3mv5LD6B4n89L9UKJFijY5MnkJgKd3E/CztvMyIfzglI9iCY5
JYUijDqCZjsyR5hl9fq+zaS7avCgW8BQXnKD1BuO/3VH7C6Cvqn/yP7khZ9/2k+r
MpnAInBf5w0/PRGWtZSYpyFE/L5pbgqGFHOwHNh/nYCUHPlmaC/lPfEy5m1FVj/Z
rP79rcyOQd0qVKsigmVSSDQfrdrmZH5PjtoJqpSezJfo7uUhBepfyYwH+sKLiZkw
Dx4qJSIZ1D6sSstaho7k9kQWMKEgGDk/KhAtvw1gUBvUsdjxIbPjiJWeUZwiNUHJ
YfMkxH1eb2R7mLkyIVQsK09/J1pjtt2mH7sHKdEK3eRX+70xAmAziwUuW8COJjss
dZi2jlyvAE9UpXpG2nYh9aQHMFTUegeiTynXMUMBHgPv4GlhLH0ilvKDMitpPWo/
CARCztqmSk0rb0XGf/UV5xzVdaqrU7qu9kR75kucBzs6L5cgeHp1/cfp6E/GWyma
2nDB14m/JB6sc15Cs8SbORZmr+KPh/nTvWyxgQacS2FFZLtAm8NGUl1uXPioLCyo
d5xP2MUhgtTD0WloFHiuPsFFAatdgHXgCsWK/UQp0z2AeNktTKSULRL9tBOWlF06
QKJADavjdIV3P16VsHLUe1kmeYDOQMCAEE8eN2fOZMRJ+9KqIq4WOAHXny0w9tMQ
Dm1gMEKHCChzVeB3+kpMCEFE7Y8c/rd3A/8PgxulocUxIFhYBMUYsI8mmPRovt1a
faEPOiUx8Ock9ZYK4dSHvlPl5WmzDcr/LEQq/C2qs+VPNCqWOXZtuCkxlbL179Sv
f++gKpT+QzOIpa9E+pGNU6PVsC0zh0waPhZX5DQJI6fARlJeNRejqZNya5yuXNEL
AVYbWmO/pR7vxUW+VOyZoB7B0OpsJwdOH3tmU+2VoQS5PwgkJHQDeRlEx0oT4sTB
Ybs1lieyKPdyt2bNLHR/BHCPkCTRr7D/yItKeDKZBQemjyRIiczD5dPBoNqC/pfp
k/6+D3VfQ8ZSD7ROlYjeuJXtmA7n6hmUVcaOUIl8Sna855GFvdR+FnybRleDLkUM
G4WAsWVrGiYmijc4dBMbjlXZtlyGs+pvH3B5PXxAwh0c99aejWDBl9TopLkKqChQ
wi0ygXYmyPSOaqBDBopz6x6tHcHBvFo/RoI4yQ2WPuDdgPxgc+MH/GPwVwiYJxo0
SdyGl2x8heShPBQlT/9+C7j9ov0bymx6lqKUyWFm33GYtIutfn3mhqA8m1ZMIBM9
9H7w+QJOKsOKupZpAyNVsZCLuHtkEuOoghVl75iCbXGEVJWpK2f2CEojC5pkILfl
SYnakffc0UcXC6QSBCrvVstmb6GlbwLJvyCTQUN2YXrptrel7QRsgZYhX/aTvR7a
xk+Drqxq32Vduq1345iZMuFOfBlYZ3PbYsPJpsYuQamvpW/7OGI9nUQEIXT+Kg9C
89EFDIkIqFMGKRGWn1HENfjDSPmSPdR6OVPMBxJLlqOHIOjXhrWuvQ0Rr2x66aQd
xZmYyzdndX5tZgUU2296VrjmajHyNDrH6smA1m2AnhNRNV1dMwu1jlXcaOYoSwYz
qi7bh7IHMB0og6Lx42Ox9L5MKYTVmcHgguJXG5ihePswAL9r4LHpY7GcjuKOIRbt
fCknC1t+4KKWKNzM6Kut6LIXbjwQwtpBReofDPHo8jRpWIh06IgVKCU6Mdwh3Bi8
9XSgBrcL63xexkK1PuIjj4pwbnEvr6sgDzrN/Sdk6hpOItJR1VMDVDbbUGQM7hBn
9hZm7M/iOxY1YCdQgnfPkJT6uejV4Ln5yEMr7Z4OR6D+GpOkqN+cS42nsSaeoM5L
5/XdBL/6sXgC9Sc1Eo0BGdc4xN9hI/iiVZZc8I/B/+0vqp1WBui7AewGuh3K6gGH
+JCudittJp5jBqGVsS9SDm0Bm30uXmpNe0jGDXKg/ZS7EyOxr3LapfgovutNFfop
hHbh3/OKDEbhP+oUv+h8LBBL1DqYl+LFO+insqg7dHlvjcFO4tp74QiDHTnXyB1U
CYxnwrJoXjpzNeWc2BmGyYhHxFAKAQGFR8ph6v1JVCbTOdywNus8RzxOM1mpksNc
yBqVkAY9Zi1WrpYD5jy4jpjeuQvd8axJUUb/ispxPhTuQvX4ECSezjvuzKIede/+
jSE912efV+3Joa90IkZLgbhe3yPo5Yp2wkGv4xcD4N8cabO0omSoa8erJziQ5fdH
OVxSCGfU9+WIlfizs6rotYS6cr0mVFA/JNp4ySHSBdv92brt/OP9SPueBdkd47dT
vy9q2dXETgsKqCPjzo4M277aaW9rCSEJJYkfs+Jo3es=
`protect END_PROTECTED
