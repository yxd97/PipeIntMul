`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
12AbRbVekhbd4G6wd9HhJqfg+VR2jb1TgzYtOUdG7q4x91GpP2CKSsYUAUanR5WF
OAWSgIOC1qt0nqA7cQehZSF8jfzvk56veQ6xcH82PptMqoEoT1ji9LBBsoX3dUYw
apgwSLU2VNhvZnFoPdniKY5oRyrrR2aDvlij6+/66uv8zdz3p+MozrQHXkTBclln
0hTQObGixAXFFV+fk1hXNmsmOEuwHUhjdxfPnIR9ERViu62nh04aSQMSUQK/1Fh+
NxPIarXRZzJ+x8mqTaxUMu1VhiBoepPYWzLP7B3vAGhjH1+14LAAZrIz0cUeNQgV
Idy2IzSIFvDix4aoxC7PXjfGqvRxVtdEyN/woqnReQkmgDG1Y+2gB58YHwRP2Puq
XOkk6Wq5Rf3J+2kQT2G3NPw4ded0gD5tv/j/0t7i3KMA7jOuUN7cYkvEMHJi6/J/
MQ1uVxLZcD3dWySR9kRE8jRtJMm8HbcqyUR6SNBPed570YD6DaBQB6eFO+0zbLxK
agVA9Xr+Kuye4XAroMkv9Hr7QxoccJ4VxCLBoCKMwGqn81dPGFeYoBj2k1eSod8P
Dw+98WoM1diGzu8ZUMtb7XuRFcKoas7IF3E164YIJVCZEKX80cJ+EluVVn0YSgPy
8grAn9fIDi2HbHTxLhhdWRTnVwTLCMIv1XUJMQ2ibx1SI4yb7zFXcu8qQ27+cfLu
CHo+3WlcJoaIId5HN4t3Nw==
`protect END_PROTECTED
