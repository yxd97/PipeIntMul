`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpCbjsVP6+6CtwEEhq4ZkDGFV9jR3Pj8N4W2N+BD5zd+3KciBO6t4pV0/oYdez30
RsMwfzXUPoWbQvLRy76oTxWI1UNExWkEwAzsEppMsYMKM0dY/50+ds0g+hwCTOJo
y6o5H0cgGQrbhNg26w1Lhp5ELnPzU1hfA1UzWRGyu6O1X65pampBxE6Uo5BRDwKi
Hr6xgxmKk9WsUqSvqKuckk2uz588NdAFvmzNn87m/i2IzjeGXSi/N5dbLqMPTCBu
WwR4195Sj9TG5JYq0y4cAmxTNjsELaS6hAVnisc9kj+qrzof1fpUd06vQL7C3MRh
JSJW3CCzydIE9LvAHShkSIk2zqP2YhMSWWO46Gd7xij+kDp8raHb3Ai2kd5EW7qH
VizevRF3Dq5P6S1BhbKBTBqh/F+YHkVtuvSPMc9uynivgSWFtQBQ4AbL8mOmYtiU
c6dVbHMAFlAIxmQpkzhO52hBm1IDWGSr42rn3kSTKUzmtNYbyZFK84UTr/2p1KW3
`protect END_PROTECTED
