`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xe4dE8/DlH/IQWSfL66oFYO59EAaDcdQo12MWceH3b/DAeWjP4RWDZDT+Rvjy+w6
LtYseIb2gO8KgIYkIGZSo7W6g/jA99d2QUokZ6ef0CHWN0pgrLkvKnrkxUsIaVah
qFvrQTNMMddUdH9RIsZPXnLtoS395PdBYjGs4Zzv6YNKutvLp5Z6E6gtkTPbetiW
2NVpqDTLYxhvFT10RcPHAT3giz1I1XZx3/iafDuxAwMNY22yWSNqmjm+Cqwot5bV
qWp0bV7B31DLt7gLjPi1nMbpeNMQ4wm37ZKPOwIpzYvra9uU4U06TXBg25H/8aH+
NbX4Xxaw/qaBZlurK45LKH9hFLH7oEYNBHemfzCxQ+aU4MKuKIpVoLCqFLRsui3+
LmNydpFVfH2tZmzJWQAXAlSeG5ZTAbG/KNdsAI8AL6aA0inH79DkfnFVRFpYJ2ml
iNwdkyVZ/IH7V2nX0WljdPkp5OkP4rZTQyK6xXHIjJpC+PPc6vyY5vs73M0ufwL0
+e7i5na1QPWI7++8baBGykudLKxaqRY6jmGf4lpM+COeX+xPD9uS3QQMCfVxLL93
2VpaODdmBRrN9bIaaUZhGXxJ/1BdYBWe9PwnK5Sh65t1gHz6wpMHJNIFlYsWxQZj
LRZA3TnvNn0bVVlNJPU7frsoMpo5FggeaaGLYVqoHKePZSBmsa0HoBed1PK156cq
3J7XZKAsEiVrj6/F6f1b7KsxJ27qflwguHTliSTNkkSlasw3H9QnMTvDnwD9rhim
ZcxR/VNaaPbIhAaU3Wr/tcv3sXdbpc7CNASZNgt2tkK9Y5kKNsg50ffBMI3MqxYu
gD+DuXDkIYEuIN9opc7blPE9uwncgnLqS1RiliVVOOHHPX8y0qIQUWI/PGJegB0W
AKjS/VorM171tWNASVMHO+TdLNdqGrkvYwQlsPyDC9pyB/6J9z1tqsRciGDDmBv2
BbCEIbRfgNPqICSSgZy5ycT1qHuLD82BwBw/At5wDte9eX/Brdb29U6+PfyzJEQY
y0kbQH7WYHPAdz8bEAr/gcqnAdJJGOZYEKxAD6PMkEc=
`protect END_PROTECTED
