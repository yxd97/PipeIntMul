`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yP3ArAFmi7MVL1d5/yyZNExgkRyQbfmUvhvb0de3FjlS8RlaomTIpzxDjz8Uh11r
pwz8HrKpvY/xwyVW6HffULPTD/QBGegFP4denPmi8tYU4RpHCeYOUeCb30otElPH
QcNmmYM2ufn7SewwlTy5AEHAvaQDSG+pCNXoSzG4/TRvqyzcQ5BjUnOxTDZ4w3YH
Hfe6lBp7Ss+dSshaN1WVjBWsIELeHkNF2cETe5REMxKA2rAkVCJhNksHvxwVbnek
sseO95hQ2d7uln6fTzZISVy50gaRUEislTyunawf3FGUxeuP2m1LcfzbmXV4TeQj
0iPL04hrL9pErI/4Sxl6z7h6RPMp9OD9RdvSKbmv36VJg/NdUl2Q0Knp9cR8CM/F
30iDReuBInC1K3PtOzFzWoVsNFrFD2Xxdx5ZcZe/CSzHUVpG26VwV7JZHf9vUx6z
bK/pEHMYY7hklPtyMTrZRmZin5oTMM1oPOcXYTvTcINQxVKF2VQGGhR790Xf4oDb
os7tHnM55Mzglql53g6zrXAxAGsrU2L3Fa0i96GYTd0+W/RFk9S4nDGMEnMg3wAO
Sej1p2bGKRxjPedPdUtPTPXmZHFHuG0beB9le27y7CwYyaqZLRr+u5AHCreB0NEN
JmHtPdII89luKndFF24EYuZbcRU35MeraySAO/fDwKk4/PeSae4rl7fhhLYCN6uy
9HBZy54GpLChwsR1Rwi4dTVFl2p2WI8d5pbYCHqTYYg5Y4YEM84y6poYfYMxDDag
DO0WRCtvnB8Wtsgi3VmCbpDhsOicTjuIiJucNvPYHLy1Z2Pto6sRELOkJFqXEOJ3
sWw9jjCAUS0m/uYo80jWtAyOAll0nILT3uWBd99AkA5pe72cmfB5FiuMeOKxcjlt
ohJMBy7+oJ6pfpzmwFMI+YBUZNWrPmvVETjt5xpaey8DwJeLaRKrSpV+bsSdvEfu
`protect END_PROTECTED
