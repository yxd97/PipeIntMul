`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nHAIrpVayewg+Wwdb83ZUKc8BQhLScomiEI8AhMnDpl7Vyy4QPE+3RYMm/MmPzF2
CbS8llpWRGI7XTQI6XrhnfVSrrM96QYGPumB/06J+sq9eZZTc0UGeXd894ETtRiJ
afbQZSUlebt6PHXueYmD/SU97E7P9PLwoTiXSmot022lW9y3NQ4n3GcBx+yMgTZ8
B4c1TwUBhlDYQBI3QD0K/EIFM4/cyBobAE5R4hN7RFmuIAxLiDdYxm5nrsOES2bp
XZU83HKok0Sy6AWZ9LC8iU6WRiq5p3NkAzFpQBsmUX7n9DDSdJQsVewJNsX9KktO
fsho8dKL3rUmVTYW67XE4CqFzHqJTFxCrBsdvfAO4mwOpTnpMwO1pAlk+5I6O14j
wtdqmAl9lHG7eArquGpDyrhuCy8xP2S9G2ue3zV3SRBeUs7SN04ZkfSDwVUYL6jO
3M4DT3rn3Vn2xcIa93tUI6dHRhUM7PLnz72LYz8ikrwECOTV/deHqCzDHCmgbBX2
/irR0iq+w5SqBpJhwRZvspcHVadSWNAgz9V4aqUL3KGxy1/uJg5Y+87rwT/yY5/U
w8k3tpGEzD+lMxaD7JjQLYRGHV6Wxv4twyDUshLAL1HHkTFMzPtUh4jwWBuKgPlX
cgG410miQdRHCFnAWLa0k2oRx5OCM71YSxg1XhbHp5iE93WAk4ZrV5fXyNaXFSjj
tnLkgLWSdv95Ux3VqHH2n+wR8Mw9W/6dqpj60NA9hrwfdgxVSxWku77CL7jnBA7v
Y1AUW+sQ+49es+LAMMRz6kX9AVSoMTZ108f3Nb3gGgoat6v4Rry5ZmOiNNY6WWuZ
8bhhNBsILF8fVl8fKL7MQOfFqNbIVE9B+lb3AZ70RdAUsq3ABpFIpq7sCwPFKbF4
EFVfK95QeDvDWLT1cJKv6eoFsZPSK4jLVD9AjLh4gHmOPfGENrexkO2BbOlp7fvx
yefISnrra1wcX0tGawfoPROv87x02j/bhuK5ZaotqCkSF/IcXTzkGmJDMhudmg1p
znJ6BqsYgS+72dlIDPiEXhxs9pLDBospvHpgBNL2OoC3H8dWWRWHBWSDs9js+NY0
dZEiKGZ/0MCxww49hdtFGfZj7CEVaw4m//KAj56lPfTfy7VPE8VIWWp5XJz5VMUP
QajBxNGpNoxujTk9/yJijNgKlaYy2HqlF3d9DnYISad5jgqtNwuMkOfvQUofURna
PRkmiJjKd68uV8k8000nt4OMY03WTUKYPtMLUYQGlnehj11E+w3aqMBUeuS1Rd++
`protect END_PROTECTED
