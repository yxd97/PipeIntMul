`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GoB5UHy7uitOTOA30iBkqvmjyrc2G4SjWfFtiG2oTq3SHCciyVaVdFgJqGzA1cxi
D/3AP6aQi/huuD6xehfBccGhFJuzahpjVKXEJasObXBPACwMiPyIHo7C634o5LSc
uKKy26+tYT84cBmJxeZtmUSLDSC/HHxu0sCJCS2u79SKnZZEmhhgC63IjXgE1DsE
ae+j5RXMGQK+xbwCOqrybIN4whn8r7WPCA9476f3JxR3cmg0RfTN9ldyKQRwfakc
OTiddvMJmiwW4romXzBXQUNkhs231JlBFHet9DNK/oa+6yvQVBQQTKVW5dtvxkOl
Y+xzBhxwXdthFwObRez+cgkLVenpRO+L4Dka45ZqmY7UKE80dDG5U51YIO1N08V8
mRuLAkhNDms5Ix745NENdauho0//zH5XD1fjG+WqKkG+NACJ/EgV7CQ0/Z+3bhtp
tJ/deQDZI+wXI2g4bmXVUqZc3Sh8vjzpz/cEpZsYDFF+w/U+nojusUYYNk561LA6
`protect END_PROTECTED
