`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EC7SX9mFVfG8HHiEAeUQpe1hxoNphC9lp2n+HZ6GNbUXz0C38z4GLRy0e0BEij75
hdCRhFAZZvEw02B/rrniOo9WBGUppTtTey3KE6OqjffAraYAx9HZmqsjy+87ba3q
jRPdvpYqgsf5G35YGClzDvu4b9k9WzGuyZckJ0EKS9q79pgl0c0K+FfPseaEPUU2
kHEuAU3h68Fz4MK7WajrAnvZn+snggKl/qU+H1Wex1nP2Fyl+mc0Uh0d3JpvsPVX
vgd4tKcHcArKbDeVo5RD1iRvvyL7v79kg8qh0ZQM9qxKlBR7NJUhe1nBMgBUMw5F
lIuXIAUsbLXcZZ0FcxfY4NpTD51sPzpSRbH+YFF9A+8FOnjnQnvsgTIaSCLAHRxl
5O2acPLtSoy3N564hUFue/Oa532Y7nWqNxOyYgUwLtU6RBL59r7rr/ydYl+WOrTw
`protect END_PROTECTED
