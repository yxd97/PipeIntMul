`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uUuwmIQZNmJwzV7+btobKt2Z4Svz1qZehgHs7MpQSLC001n4/ujbbX3BZNmImo7L
VnIITTN10CT+rj0BfeC/yiFFGVcEsa5I/z+NZEROemJK7N6p2bynHqjZr9UPir1e
wJHww4b9cNz5PvYQWf1NbLzmHL/FvFhQCCr0+mz1GegzsZqw52PeZ6qmzybetf9D
DxfiScc/3RgRJ9aoAKlH5YRgFHvvZ2oONUNTi+udOCwyVvVaPgB7HWU3DLPGo7Xb
v08mh4uzl6PBi77EB/R2AtVmb0/wm4/uSrsjXBN0utxHd+1iwNLFbvOJoAf7kzvm
qUZql0QVD678fk+MXvrkyjRNsHqC8AyWyMk43tgx+kZPD0g7pCVJ+2PxmXW/6Xah
TkIp/rHc7no5TsZFOJdJyA==
`protect END_PROTECTED
