`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrxATEbaXJiq2Xchz/1tmPMYf0Hek51M+tMkFQ8AmveCt9hCYGEFQbaQifrK5Skk
JEhTThF6FvbhkpnBzMfS99b1/NYi1Fn7OG7sNGrstG9iJwU7yRGxepK7KWQHtfyt
Kxltr6cUGusiffH0Jhll6xcbaoiGLILOvVIRPDhAArrU45d1qeHpeF7ph7TsVPRH
UIHbBUdzC65VgCuiMxfu08j4auWMzPhSc41NFeJfGceahsb77sNiutlkpUXs0tnm
ZgG3ywm4iA2ADW0rtziRSMq+yZmW5Nu6QD6UzZxWq4jbo98fyyQOCb/ZcGXa/2Qt
Fwe1OwwY9UdqOD7GovlQ+CunFsc3/gk8+FzDz/bZq+fomkpu2LhyFyIqPnJvdTGf
/UaK1a8roqk5P+LQhRtcD6In4re0yL8xh/8cHjNvJQ8AuAk+IAY2aogybLqOJyBL
TXZE1bkPZ4T1REkaqxbat+NpesGsuCgatyZ6XOuzALYURTF/bARaZ+15d/GDMKJh
IY+oewNFw6DkhzcR10W4Fba2sn7h1hyB97QMgxoMFTV5U1kKPUrPrvCZAqRSSp7W
zsnsl/vkcWJiGnrZjRT9q5Aa7CgWfR+B/5e20YwFKtIK6jzAGmOJvc+KpViu/uV4
+re6YcppAYlDM5hk3RY7ITzssYJ6tGdhl65V0qIX1+Z8DIjZseXWmRk8za8LVjsg
br6kBmhxKVh9RcafGfet2TzvV8XgFqVbp0tfCZI9gXYOItCpZtAQxchE00/FugpI
5lDh6cl0I3Q1DVuGpOrk8fuhlxS7SEiUj4udcWxsh/nkGiCh6o+CyM9k3bhT2u9X
TtzT+m00y9GkUYs7BVGioq8Jk5uqRju6Rc4ktW6WG7ADMKfTy4YNE9pneNPt3aqw
N44h5KXasQ4Hre8s7OQ8bCOf5SQs9YfsMfqLMBWNkdXi3LxgPyP7JQWR+tKGYsTq
BdG4N0hAZWRD2QDXT0wpJrwsuxO8cSmDyV3oA2NnSuEJawjRClnrzl+edWzYyjne
fEQJb2Cls2gTDAQ703DKjWfbVgER3a97SQfBeuMngTBtrRr2WWYtrbUoOW5QId4z
sU5xScfHAiBj7z69wT8GKg5LNNhDw15QmJ7AYy1gJ5GZbdi0FASXLqBRrPJpJwMI
ObUKB6Urtx9X40HAxT7YSe1JPVNbH8X1soOZAtWbdL9KjP/sXj0R9Q3H4ejfnP5m
1z4hcWFPszcVjfdkA25Ve7ugRrfCjOFSZgB22BU/rxX0P6cW5yhKw0whgiGY0jD5
SvXRfclA80o6QjeDXQR6WQfHvfjh7r/wOBqIyQEuu9c=
`protect END_PROTECTED
