`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hI/T0x9O9SZBiQ7XfV3DKfGE1xQJ5VeUohNGoDH/TinWlR3mx06vS56N2d0Y669N
fQEfJmFG9cAHsfnD3dKMLiKqipvalNBP0IMCqAAQTXBgUBTzmQFayDIyuc9pS4ij
3KF5nNRyT3U4SFRY+umYWXZVOpR8mjT0xE8yCKAhFfgWr8+7wRtDQvY7wu4YDuVa
y91J0kfCcaPh7acrddKYskmdJI2E04zMg7noAIuwgdN/zfMioUF5UaxajAIiShmL
30cYEJg4a2W/EiN+C1RZSq+nublEHqHgymQQ834SxAmX2YswAy7XvnTkRhU6IHLg
necjmpcS+XPRfCVC1zKKiIqJrKav2RtAwcmfIvH0OkkptVy+8cxQk/QQW/+WRv2W
WEsz1kEi4YgBabV/mcdZOVOVPh71pHxPGLIp7pNWL6hZk+1YymN/agsM4eyyBVb5
ScQ4lN40mWreZayasAssMF5fYrvedMSOopGEW7Xhqf1oayH+jP5U5C394wA6hh/a
TBfq0JH9CoWVZV3Iys9hWEwRQtOyCezRlXK2gxTZkm8ThmvpG77v8dq9GOlPUyZO
UL9+g6sd8hoMd2Fu3GQ2jj9Zlpza/PHC+TcRZ+xcdeBYAgB68E8MnFGH4S4KCmEO
2oNluK/SSHGqK8I6lyPO+2bV6UQNxXZEalDVUGmdqQywSf8W56FU0kzsm5eEgwbH
`protect END_PROTECTED
