`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0BY5Q0HOCxup6B1nAh4FfDle2HbDvwjUM85dTVyDqlYnk2mu/mtPi5W9IQTRT4F
lfxZtL7z7dNbzwY25VEimoOkBXSH5EtXj9N1GyLyY/YyTuVI3dNJzRPa/xDVmvYm
GREfnZKjy6XIFL9dDxCF8eAuTk41a4+seinFSmZx/SAosTDXaTca2hI6/v7l4qBE
l3brVMhuPhhq4pRqUypaFbFUsiLq/ZfBt4sbmSHGLgJg4FxQ2oLFGR2UNzuEQMF4
dFoCgEI2cIyf2qtqP7R3c8ndjatx8uc8YQqo8VyiwAhWKj7Gu7VytcuwSuthC4AP
r/zvjkK+EFWKc94ZAOCdpQKuQWxg7oJ8avzipnZXzGJcKY/WDiVxX/tu2gE+UWHQ
9qbqsj8qVIwRLxjod6YTb1VfQ9fE9gJGyzL3SSu7xXbviVXQ9oYPx6ZQy4hDk+Y6
p/HOKvYwXbtWMC8WdkQDwelnDNXK/XiWoO+tQjKJM/TADc/inygwIbbwMlghQhlN
GT60Tqa4tEIbl8F6roU4WVqhIvBARMIixo+c6IdXXu/Ui9a5gZkWuV48FP/iT4L2
+LEi2Hor8mZju73B7YQPCG5/ZgpeCTaxarsFxcl13FWZ86OSpXJjMcDxnX9G4VaR
dDPEbRtGx0nX9rOOcZFYt9c2rMQ4ZFA5D2WNHvQzD163wAY9+KKMplr1UFcnSjy/
PXJ26l1fmiwPlbi7pEGJi2d0Q6nke9u5N4Pyi5EU69TuQBe7xzmGOXXuVMKWDLTN
zxrFUVKKCLACqvVpXIGYPqtpLLhWF1gq7lGlMNq9h8jSU5wdcXBp67FpX4m4nzzt
V6NLWMg8NmUeiJdMOjtbxCfE4/j0unA0C6XuyzpgVbLH0VZ4br3bkA8ve8bAP037
02kaLfKKjkg0IR8GYP4kb9RTAceKzPA3sJRCS4qKcUCdBiGjmCYyXYBAElSUS14t
hxnmHn1T5pGgTLOGeaxQo1nYN6OFWPaGKSVvjYPAdqXeJpP6hlmyx9b3mvoCnnE7
x1DwkZOWTF/pmaNP1uOIIBAbgpdagdkDUhAkyC86oDkxVAesY7n6hpnG/0GDO+rt
pdfbykrstYqf1gis843IiTEO5vwEIi+3rQVYC2cj64YZfegva7fWrggq5wP4HxKr
JnjOpZxYwQlPDIiflSwIEDP7Q6g+B9aL4byMXYTyVTI0mp9yPVfhez6ZhtTeZEy5
HtsX+spWb6sdk9ZpruiL1edSCjWQpTkq901WPoFN1z9F5P89nOSx9QqPQ6ZlITUk
rxLJVBXc+Sg2EIHo1lhk8RLcASuOcABUWpEd0p5KLnCk+viY0cRh4xdU6l7ka9fB
1dqXlgMjpuT18nVeyacPLxV+zyrIke2v/lz34GJj9E5sm/sgOtSETc/6eDRzTpOV
6Lejd1FbAfhyQMBugh0tWA9sCiyiJkeOQiIiwJ0AwNttncjrcKfbUuEtlgdOYVor
1GT1yfnhX+peVk/b6ZwbNLkcG0FNIeZhZsuthudVtAhaQeLsR8bbziyouCrwil9n
SvNtsywXy4m9DzEr46Bt0POsdYzSa5WlDNdtivzukL6p1YeQX2GA+ku9PRP/bxqD
WU+oBAU7tz0y4Fgxecn85o6TW+oUiN7xpyt6dk4LSc2JUJWGoSXixqmUWxS5epgx
w1Ovk7U3ab2S1fsa71x3LANeZ8nk4NuyPP5U80u1a/O9gPp3xst2MewlPEraOOsT
rxW8F5FeuQ7ssp43hQEBRq3n7Gr2IUUKOBCmgDsCpT0JCSA9HIGtmjJNVDgq+XYo
3bojsD/9BEJyguZwhVn7n7mbK3MErXz2zlF4w6o27+CIm/B1Mx8Wo8p5nzZhGso4
hvzrx+L19dXjsYpsd/Tjh+uBoejs5oBXBu1mkHqP/CI3+9rykpxhVF8glrnLYEGN
xkyomuK8wryM/nl4V4y0B1CJEIJ2M6GLt4Feny55/DJQjZuTcdG2r+a/JyZpC3Kf
e7fVJM5hyXgyajew5HLAObu9fFKhbTMwjNE7nBcS0CmXz7om5IyQEptTmj6MrjMq
lm2Q1fTVAx0mU5fry6cUuLKF4DiJCyV/9Xp7VGWJAVdKcB0Fy+/D/YpMaV5kdLAW
gd6nsekCaGSP+f6PXqydKIDRidZrBPRix5DR3ozrdacjehVfCvVtGrvziYNpRPJP
id4nVCMacU41zheVcYuB50VwTYDkkusnTz8XrdtMNrWYRdeQlHTDCnxDoxJTvzY/
rZhN2VQsem6rI+HF48lVqUEIQY48VgjxL3GrB/5sBIsThbK5XcE7Cc11nxZSAMQ5
zxqP1ZLMm6Kj/HBD5wzuuzLibcr4TskomnGNhYXaX4LCBv5vuK6xke3kFT6vCr46
QtIotFLCZlREQ4cWnFdH2bq7Hn6KvsS8p6IN2MqFRLgwiXml61rDCvI7lMUdmlsw
lB2//5POsfLbv/pWIeSsxhG3uYEwofccAP/Cy27iAIGVDmASwFogmgyu9e2em7xk
ClJGH820nUG0ak8Tomc5hCb/lAGw1EGb3uUAyzxbtYAmfRGf6Wft6zPTgIhx9sv4
uSvS//DAf1I/jZPCVFRptEuvJ7UUD6K40pPiyFRApEdR8PMbCe240V32qIdkvVvq
zCp1EtAV5U99GdpNm3Abilu3Xysq3HFG/dNNX5gGrBTaF9cZDacyBXos1Kj4mRIN
sP0KJOPuguYaReEnFIZ8ANloLn5tJCz9O9qk6RLna+6p0gYjNzxXJ0WKb3rUZntG
4zt9QCto3F6eueSN9Z3jCH9EOA7uHSwi32wVFanaqOC7dxv2WaM/bYpGaTUWf7Iw
18zF2Gx7pJw3w67xJpbZ1deqr+VhhqrF2IOtqoWVZfB6UZpe40IAwt5KkJcbMfgU
Q63p7U1pd1+1FRlJ0My+rO2N271Sv2r+LILKXSBj9VrkETE7RUG9A932gSAxma3a
SJYoYnVtOlOCfQAgBNcc3vGH1T8gVqXS8AYWM4jkz1xiIv/1XwyylY7CD1A4SZ1o
Eu6bg1JtN0fYXRHve2oTDDsIGHPfIeviuEMPsQktQDXJBy/uc0SnMyLueaf0HjkW
4CQ5Q6IEVBug+hAPp0vKl2ysQQxIQzL/Mmx2KLtVvoTvaa644395/WAxhCLRTMMI
D7Nr1ZTm0hY5D0+G/bIIVdlDn9b4c3tFc/W5eI7Iz5YUV22r69l3oLeAD+RZdBKD
YyYGw50c8k3fu7OZ0e53H//P2dfH9HS8L4e+P3AvBUIwS6h6M9CTkTBjd0kgrcyl
TGk5USkNIzA5+qTR/UrJ9w==
`protect END_PROTECTED
