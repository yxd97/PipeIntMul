`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bI73blTFIKi6OfcjHQJfrZtAZSfqk0+ZvNfgPNuuwHmXbo+5KOfU+K4U3p5TvyQc
fxIhl0d/8OvRVNDKvx5rCp+A7oKGDFrM7fXdnEl6bXc31qW63lfvQjnjtg9iH8PX
+l02XplZl74FncoKrxNK9XU4nEQKg1YyX/W544VIRFOWJNY8+hoXK/3+EtzzzFy2
a0jdYk63KORaZsAS6NO9dR5pi5vLitW0vs0ZdEQl9W8ftiEn1c3mjwKVSlxEE7P7
eS1CvfF+rzflCSBVE9CbqWUWY43yFkD7hw4RLyZanVQqqYO6RlGYZx+jxo3Lhrmb
83xiYze6QqdCbKi9mM5jJPIVF/FRxKBfh+GjE+xaPTh6+llGMTKtnQu93GRdL/Ne
oXzdI5f4iWqDl9npXhiBVwtcA2a3NEHvryVVY2zqInpsS8Z514OB9Tx7A4NHjwMz
SCboy4+a4YbqY/UYFUUSPpU95hKjLjwdEbHkgVkl7fw=
`protect END_PROTECTED
