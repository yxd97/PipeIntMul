`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGiI76QHGLqE/iiUaManMVnqn3trX0q3rXQ/2wg7uGO1fVEz1JFdKUjaD0VsCe8C
iGQRyieF1FsW04u4AyTHD38akywrfUPXt9xgVSILvG3RIRUlXgmqe3kUtJozT4Zt
aL6B4DAjnSPP60ZGPTmqx+wgWbfk+ggSFw1h40WOC5ysNx7fh3nTxfF75mQginaS
4ATRe0Sy0bh5p06hTebBH0g9DWCwVZBfoMTehPpKqE4vZkxJA5qrMATunNG3pwZ9
700g9LCdYfGMhsDBYU+3oSoZJzEU1D1p7+31N8HMVzvaTYiT9N4s7ui9y5mUGKX+
5uakTFiM/IuIs/p4LcCpGYsXjIu+4ew6c5iJPMkWkFhbkvxChi/r3qpRvJMRMLKP
8yIs+JPZf6Z27MA/wMBgBb6V66SJo5FQI5WrgytTmlmPeHx6tazpORkXIzuoJbXd
YKZcYGVd4zJwC6Lq+hoL1h5CSkfEsoQaLvkldf/vWgDj9YeyRcF9rexU5xwprIeO
JAotxlcstE7LqRIvD62mHqlBVZO1dZSeEqq64IkHD0CD2E91/2gIVaWTDGnjrFT2
tiIuR4uPIc1xTovS8h4OlA==
`protect END_PROTECTED
