`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcQg2LC+kfHfJZY7/WMpizkJYemPEekZD/kCCfxOIdgYj8k6udC+ceGwZeXcDK97
iHSi8ycbPZRi1SyiWnlv529Y39rM1525ITddtt7i68MEGopgo0/ZCkYIoHM6KHrS
UYHbxVr2nZzrGbQewOkgkT7poP/KrpvCEmVNGAUiRW6UBQVwZ1Q5lHwgdRebOeBn
aidjH8Z+GqmHcZ5zLnL3KhtfXVbsrUiKxkq7oXvriwvTN/HGSsODLIcvYqucD8lD
utSag633zoY7h7bkQwIqtzWlPVlhx3i8G0YCqlMtmvepHEtPmN6R0bSS/nDMNXeq
yQNaFEtlneYLjsMUGIbW2fst2fb65t/KSMQG6oX95vO3ikDGOj8Cn3XCS4sy+2BW
DeAExuPncI0NNMi0arxKLmIrdFeGksDcBUV/BN7QQksSkGiqj1wMznBLba/sxaJr
`protect END_PROTECTED
