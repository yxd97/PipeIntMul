`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7r6bY7VXvBp2544Jp8GF95rnXURo+pfQlLVOv9vBv4dsKABkhZMfURb542PY0rL
Pi06LDVetd6+ufckQR1oFDHB1Lgis0iLBFB3mAXomG1hU5Ve/dJFQuRwysDqQHus
lNFzDNrfwPmKnsbRKYIE+Witsm98jvAYwcRTijN4HXI+HibLjrElQkpqTAXybPc/
/H8XZOVNWcT18yGMP5t6ZjY3Gphce6Y619GbT5foWpilJ8WCR4J4jKR15Ausgmru
TATiSDtCZyvCWfKCDaA4/BcCBIbcjEu86or8Ft9LQ4XfExgxK15SrPlfQcMYaK8m
7ku6UOTGhiM3qQXZkV9VrOoW0OAdc20fuHDWS5pzXIq84T3F+S5CoyuFZ0AuofX+
`protect END_PROTECTED
