`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uyOtzWk3Uxq4ocjkmmsDGd2dN6noBzDOGezocvd74oteOmrtHx5kEOA+LRWvzrBx
uyWEndoYorDtxwiYLqo7mFo4FbpNftw+cJGsSCBGG1MLuFbDOiBk5F8fiAEmy7c7
2ttU6yZ3KAheVZOeErHNDxSc10FbY15Nkd9l6eSVkE4L4HXHTaqWB4OQ64vRig3F
YiDI3NvJitLMEb4LosNUj1AcBoVyzW8Wn7rNXy08w4TcMN8tEu31Otqvu0Ov8gkY
Puthyb9dLLy4maavoc9OVRG4ouVIThOCkAorprie0AIWjVkqS1CV4L0nffOtZLkx
C9QqN6xe/Kmr37imoGNfxvDRYUIS3T05/vZ0Nb//gFjEwYNoZm2/EYXG07H6h6Xq
kJd7pV2725RbV5Y+hcnY0SLihlYXC1E3ybx+U8j4W6vtDIqKmSq285pzr+c5DHbQ
yAcv5bTUy9RhEGz5NUwePGA6g3KVXJ4kCo5s9h+77K/ETi98S/+lx0Mj/2tkGBA9
W+TRpGMlPA+sGMrNOFYPuEIE6lOkD12pG7P0Um5lX8R8VjeyPhEiULDRpvavnlah
kie58UbdInrZOfvTyBWdkdieHxRlTmebYAkEJ3BqMmjP9mCM/cJsGZ9tJ0Fqajmj
v47x2LUkrSNwoYOWJxArRhG2wMNfsvTqcGwhjevLij5rgM4Klchs+PRKkpKlk1fo
h1U5EqAJAnLULH8LfgLivggPySxWpbsj7sq/cb/ktlUG2OU5ggqdIAj71KYYJrjV
7IPHU4aZAgsrQO3LoXJZtzD+mcO65hITXi1kMmgzvbEIpvrwsl1qj4pjjKVb7m5d
CQ34/7Z4GjQn+rYhSTraO5y8Dj8TNwi6XPCcC51qCmNGfIQ8qnIl1CtYIip9rXPV
45lpt7Mlh4mho8TDnV4a+m9lXjnPaQVeA/7LMGUl1O1Tz3C8JKsKR2ikYUoxeGbi
CoRIHuMtbz98q0gmxxJ5JTin/aSLBu8v1Fsp8oVpQnh2jQF70a1mfexv6F9gXmGn
USEQBJ+wcoAaW00dOCOpfMwBD1AfsBJJtwjc+sNip+yonQ6YPwGo7skp9K4Cw7wl
/jugJh3q+nOvybKrn6oa3JAM9IRHvqmASvIHpBjTZWZqkdWoNDKPzwqdObVskfKH
hjNXLkArA7TdrTaPfayllsW427wNsoNnp9N/ReyNLBjXz/q4qE7mozN9gdfxJSLB
4Z/BibmYlKJHg79LtZ4r0zP3Fo+PKk+aZ0czhtVhgbksW54DVjnkXrSnaAlVl0I9
Kx45xVANdIEqQ76vtm2BSn399lg9iZR9yfkVbS1SAqfv6DFir7Thoo+57vU8Tr4A
hlEZdPWFD57FMbWqIYAw77QTsoTp1ePE/7LPrW9y2Zd8Jx7+PG/UGoCTc1Ei0bO/
g2Y/9DHNJsXh/SQUGI0bK8YXTtNNE7Os1SOESNrXWZHfkEIbVlEfH8XjVKgkYU3s
NtKiFWmNltCCHyhqZiSx2dtFTjE6Mi0vaYq7yTBMFZ2xpLogJroQolRgrUXhuxXK
uYF6OAzIyngAdFWblV60wGgKZ5nQ0Zziw7IX6BPz8qTD42oQqK0VZYHHeGqz92nC
cU0H92m+k4yg3qNntPbUTn5x/LozEGU3jgLNurRS8RYziCuH4ZE56MX3iQLHuaFh
TlYKa3wh4Dmj3HuZ+Q3WdPDphtyac6p/7h2jt+9tnOTX3TXC5cNhgk0IpZj2rFWr
aTWme+r0GLkKlGUUozJGSqRNuBFUTuDV62LyJBULuDtXbmQIHKZpaywHRyuBGYeN
jMIRqEYEvUJtv4nGyGouXLtbS5TYW8ER04XvprMr9w4kBF/USChA2Wj3pWpdYALE
BHQNzKFLQsH0pUAWQ5AJ4wZw8q61FVS7qqDu7E3jNYzzYcMqRwZ6oLhU2bHfZ95n
wYoLPX62j1SaG1u8JNreNrD/U2ybYbR3+5bdZSghXGrcOC15x3oxnwZPXEMLhhKj
GqOCHajhHQegeYG2R484phMoBWGAfnP4V1hsjiWcEg3duUljOqdG9CPB7ldWDy8s
qLXvcW0P70ForY8B7Hgt/OcobbY0S5k6+E9mC4KOdV7WSEofQE+SnRFc3UlWFqQF
DAGYpx2QJ9lmb94j6ZPg3+IHsyeZ1jmMPpCicceUdPKGiUrjCwdbGcGb9Bb519p+
02GS1VtsJj4dfnhK1zDjF8gfrzLioC7ywtrqTgHztsKeF+RMzUhtRpCiAW6GTTP+
TRGWQAC/BdW8s9xzRcgrAWo8TUS3y3lKA7e/KLC9D2MFnjuLysUuenYPoEHQd9fg
GhlXwZadjcWU+3GJqmQx6nnB2/OwhWDMS4VrkJr+F0qUmMMpR9uembaDr3hwZVEL
oL77h7trnPdl2Y+pNMjOSQwSeHoko6C2wINdHopVVEIH0i3z9J5lONMzQ6AVPrZ8
NXs4A5zQDhu4ScuX3S+YHIs7nLxDW8FTfhUUX/uUqVlxilpPvl80KKP0eY/q3Wp2
4sX3fMnIPOAaEuS7H/DcQgyAJlVwo6AKVnCb8LQ4prunIYOaDisM+qHYNRLcE7EK
RyxT0/omfTCsMl//lOJieSVKPzBr7GraUvMC1VJpAuqr9OvkWRipWGTqKe+B2snk
BNF3LS/4knzcKlNtMGY4D3wzFwk5u/OHxenOuG03y5kvJ49u92SfREmcJDMeCnCl
LBYYfozETv8WS0xhzjMvGio3erJ6BiOyu0H37y21gPxgXtGivGkApPtPP5XqWNlK
VtDpOeZcONNNqhWBsJzEaEQV/y6dW5yuha2DXrJkadCTPYRjh4QnEKOYmcA4spWy
Vg7dY1QC0EluOiz+vh6fSR1yLC5VejFzKtW2w7D13N8qfBvksH+CWbvUol64JCL1
n8dqRQTD8v7SW47Zk7cQyB2kSytFDR0X1MS3wcmkZL+8HsuJLapSzJzfU5U3YAgD
ing8mAzR+pfTjgj/6xoeq1ldv5lkmpp3bBVW4DRfzHUP1SVmhUnEX1yMt1g9ZM/n
JrLB2fZ8S/h6mHuuBiBriXhu7Wf7rISatp9viWrZTE+frcuVtsuG7YBtBJRB1jMe
Xo6n2VsG11X95DwymtOW5ej/DkhmjfMauIEDUyxCj/CDmCAl2qBB4uekSd7XB4O0
OmE9Hs5oUIOd3hzide6LIDqXWTKyufLptdFzAeHlTP6wFiA4BJREyn7fR4JM3hXc
UtwKBM67OeaWbyqkUyM0K+/a5V3gDEiE8uQSalXQlL0x1m7mlKJ+Yb2povEvYvH6
TWI59snqB1+mS03H5Rz2Z6KM3FcYwRWmDmzSoG9OYJAkbkX6ZIGaB8FSFgjoxLUO
pwN/z++z1mZYFD0zh1lq70FffZHqAJy80XRq6mLJQ7uitH94Gu1P75c06XgKnscK
4oqr61m5kqIBQmgJGiDV2U609a5GEIRtt92YsUl1Y5JifxFf2BDp8Q9ItjFPrJjw
eNoJypHmufSmaYG5ZyVAJBeSidxLAF8tF8tsFTWUvqLrgb6v9Dwyb+64hjgVWyy0
ZXtPHD4NrDMrpo7oCu6NwfSj6mdZncPXx0zr3tMf8/fuFpM9y2puB8nk2uvKeqtU
htFckTwrRqZYYQeyPPmn0kpvS9TEL5MTFZeaLthKJ73qo8ilN/bT7cAewNVKVnYH
n/AtDUtzU39ugf3+7HBZEgWLFAk8vPWAvicOH25n5tgYd8KeHuiT5HRDGrJ/omsJ
/Ll0Iv4MA1B5pqJlQDqrizTqAmEN9iblb303CRhr/5B+RSnGkMG9g2Ew0sHbOQPh
duvrOOppHXBrAlcpA0qUZTIIPQWeMg48iqKd0kQlXrayhoOw/6aHIWO+JmxMRFms
RX0++IVVGTk9QKHsFyT47em24Kl6U/3gD/0QhP7zLjaAWZiqQnPnqBNjHDYn6zvb
bF/CtryM3eL0686xtb4wG9fcjK08mswxGex53hXU8TBxovqaBEkQ93TLPBrZMsEj
Xtsy2+GRknlqaW0lD5Pa0/WE6OrYQW+GV5zvjwOg6mVq1QEB4fIYQyaLDUxBTunR
VsE0tJKvdFiR2iOq7AzQpEINgV/GAVeLC8rTCA/2wMMWIBO6BTp2aZz9M8y2R684
y+8k8Tr/AXWf0+PTTct3WE/sI8Qyvy1T+6/UM1vYmGKMCNMNV6CUF31M9bSjUMC3
H7kwbIvkwzcf1vxDAaMiBCPTC7mtIL5TVZzaJp30M+v70IzJ4mPXgpGY3xYyKtjz
DtUvsLlFjNypWfqs8WENIEtBNtSNU9IN4+3tdWgI2FpuMhj++E86hBRYppUn24nu
MSvVQNNQFmI6kGFiX45UquN5h9KKsVSdMp0Yuc0/40EEenTOOEyO674dBkEBTQkH
MkodZdu2cYE0euaPVnAhp9O3oBev7VakVfe5RvGTNxNvLWbahjNsYuHvACEEufzH
G2ZP2+TyvVNKInDAV84KDppezi0lqaDNWuXSqbEld9Dmj6morvg7iEtdrdfTTa9S
HRcluD+wFnnyqg6tw6cl91akdslXBLmx0hdp6CoqmTM=
`protect END_PROTECTED
