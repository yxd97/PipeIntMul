`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJIf6vrDelVdvKwoTdy77DfISxbr9gkVL6C+KoHnH0Ml4J+dWbmwH4IlBkbdPnnx
Y0mgNEmX7mHWpYxgKK2UBxp0SXjWQS8uEO7sl/TZ8j5yINdVoskg0ZEYVOnSlbAu
NhfNkO5BbaGSA9awjcHyFI6KGvaKJS0IE0bdCNbEDGMJ+MQDr3/eP+FUACWO3wgE
SF+K1kAmwqUOT4mDVLkOrG1uf30aH6lRKOwf11+avWRg9bNtBVzzsMTcQ2XmiuVD
AALrAXGvD0q2Oha0ErGnH9J33pTJCkbrkoB10pJ3bd04IHQrq2lSezDafUtMGp1s
ra1BMTsdtyHx8+gpLHT9q7OIiBgH1gJiHzflMEunvq4kGa1LBEKCsmW42lOs5stD
U97BTjXI2cbcRrBTuipRBVxTpIcYvGc+sUrRcTOdtCSJrjJKeBRJnWi6dN9xrt4A
`protect END_PROTECTED
