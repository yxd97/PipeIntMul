`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pI3hT1eLye5H3pRoxM1lQz5QFgl0cEBh39LzDyDcqaRawdgSuA7eEDGmDqYmsctS
aoCqE6Opgn0u5sOgH+9QJ/95J8yZGwGPMc/z6rOVkX5gJXPW2oocN3Us7g5AbGRr
f3If3xUs6gu+eymP2DAmK1HeKFaNZORv/zZX5pDJ2mowv4krfUmQ9TN4t/bHPk6x
9Ge4odv7aIxH+p0Y54jDYb+ODEpnPKZwxj23pwP6ANlqXwowqWY9JkymD+ML3UnD
Cz4Y5UhImGBEBoWsg8uSF3gsOy4gscKM3zZ0dbykKo6CuhC02tI7RcadxdiJPqPJ
ZkdXbDhRQwnasN5rat0LWZWl30o1W3x33QeuBvVGU798S1BVIPXcxzNRx1hkYKni
tM12G69Ko6DlKZH7map4rD8YdItTh7j6Xz8tSAVVT7kB/v8vLCefQ/1WjhJcFjHz
OnjNm+IyPwLhq/rPW1j2xna0zx+70L5VTvnZNCQ2QMFhobmdKipNWN30pkn9P86b
XwCcxjwfxzsOgSxg3cuZ9kS5R+eZ2d44Zpr7ad3MnTOzBjq73G868EiZnY6I5Lux
+JWFFprqnrVhFkiQhOkmC5h5PnsQA31J8r5DPZYveBK9DPhj/siz66dD0UfFp2gf
DVLiYMMhpAdKKMBHoTZCbq2ghB5qo0b7apPs/CSj/ka8DOe+OWxEGIvEcUqwvhYc
QL4X7fXzNoRfn4E4B0FtY+AP6BhGAvQ/Djo1tH+FSUvbjfKVMKA32gKG7MWJ9VlC
K7SUOcL2I4NHUNP/QrVxtpQrL2vczXaHcAlUecANHG4YRkNSnD7bz830y9BYDBFE
SxbYVctVzFf/iSN0Y0h7HxlhXM775y5n1nBi1aUiKWWZrPXBkC//83/hrOVxRVx+
v7vPT+qbbletKI/mmzTK/MrKejd0OTBLrcZe5z5EgU9Goddzf8srYmNCBGb96Fza
yuGu2TiX1d0UWyMK9YKseq1yAwDebMd9BGiwuVp0xaH6FyAxXCXkq4yWlNNu9bcq
OoAJyeyc8+UAXeNpZO1AJYGzuyWQsUTkpdbU2SghebifkjY6cGL/CyjET5uy+Q0m
shgleylbsJdImupkIBy5QqRxEBhn/57pE6m3+Xqi+2PyuwrUkH4QtQyTXdrWXs39
Q/dgONQEBFVlL8/gBG0kOMR/iKqakPoKYToTEpQ98Y04MFwZ0chEbEFpzMq4Bsow
nUMy0wS69OlbeM7MLkfC2Ylaneo8Kfm/H3Z2CnUuJ3XwCAKqcmhfq4Jm7j5WnHvT
w6Y9wtv6GTimIY98WbRXZwSxXHI1QGShalGXbICmjVIJq2sgbcGeQR18zFTDtQRd
TLlg/uChCLMjhmj3CCAlPYDz4AVtlomfpgu7Xk76a1XX1NEXQGoqNRIZ8Bw/tOtL
6zQoiMaesMP2emKTMo5AAw==
`protect END_PROTECTED
