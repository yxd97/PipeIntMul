`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3zwLmK7pW+lfj4ukd52sPzRQQZu0m8Ggi+cCazXdyT6OYRKEE2Pr5rL8XkDhq/g
FdecgALLE73Walbjop0KIghPc32d9y2JuC9AQD8omOstoB2jc80cAmgyDjI2jkya
J0k+VeUs8mYe5eWEpNxQ2tXnE9ZkjM3xnbUnJCqelLt9R+h/ZiwSD+0yAb1vaXYl
M7D4R4yP2LFRGDsATxQeTVsSJZLsudrVB8kjDotM7/Dwtf0E+AG6gVAr7Upa+TM/
GwPj7ozA2UhWekhQrIryvCvOFdI7SvRU73OwOqf54wv/WoBpaXSTTDgVdHSFsXSN
bcN6s/wc/05CvtQW+FL6CA==
`protect END_PROTECTED
