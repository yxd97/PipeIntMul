`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oXvEwz/9jMOgZoJ/hKY5CMBmLDVz1kZqk3SZkBOBJdYUWFqvsTgECz4IY58LqEql
xRNvtU7Q3DJLvXgbL2cl3msbZUIXnl3dBu74Q3mSeP8xFa3+7W7raRG8+Aqgp0/K
oajxkSp4JBbY6Wh0p5zMJvXbwJI3RUmqw6gE2sznAyW5E3yGeHW2wnePQ31tVQqP
bc4FQGwQETLlZc9FH5PIfw0KH2deBOFfxgbS5DePDA71UxQWZDKjQmyQKRwmeRGK
3dCkd/Pm8Pa7XuHftOl1Cg==
`protect END_PROTECTED
