`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qh+qkn7LV0swu70zwAVnoIuQJEMPj8cLxodjrIuJiWbVmdHb4R9vWjhoyEEpesLg
LZjwpQN7X5a7JsJjc7xkrcAv4chBGkGO+HbY+Rwy+vvoMbmfOsZc33CdkOaqGczW
JMRM/ryQpH4W5xt8huL0Dpp1YjQyYPGjHEugxU2ZZFhwWXTc5Crf9s/OKgMYc7ll
U72SK/D5bp6DvfbEs3Gn+y9Snp92prhnqWbSWvEmwMtwM++Ml0FDHFUFAxmA3RE0
Pc/cfSBKL5pbkEzZ/DMvlYePXQfUG6StCeTVO9ZNRASMxrrkPLTDRMuHVMVJ+lh0
fJsF0M6raocOpaxuJmSnRIQ+nby4EDOHzlSGDpUNdX+1N9Jp89FTz9yLBBWPSeAs
1eixjU4hv9uaR58f0o5a4g==
`protect END_PROTECTED
