`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NocBkTfhBt8E4FmZSNcFKaqAyTx5+6Utzsra1o5c2fcHYjPly2thDROPXhNL2xNn
TpoQzKtgk6l8dNE764n3mJryLvdZExxVrQNZmOCTklmT/OO5lCgv07sEV49i76QN
//tJclZhvlN4nlajpgxn6H8Bg7cn3irHNW4akmcwGlbZNQuIuCBmRwDNLU5agvPD
7i+FS1dHjPWs2BxHff967/X3JYdBd3KPvAC1TxZUIeGYICkAmeCLXwsUfcenQSS4
f8rhbU84qf0kuoKQ34Z/EBzhdU8Iia4R8osDB5VI0wqIODbp7rA2d1XZC6fG0Mxa
9PemcpVYWSvypAkPhOfJu4o/UQgA88//pIVfQvYWLkF9f5+YlW/PeK8M9+mLX7Xo
O2OcnqNOQefzqFNpx0qwpeP4aIwpKBKWr7DJuZ9e6WQVDldbZDOkz++ub/+1tBM2
65WQK579PEAQwyakQopCoyMmQ3VAMU+603aPfrO6LA0X57y8UamLA0FdX0+4XaPs
8gSLzweiZFECAFhK4DB7f8CIYRtAzrQWmbwn6RyHM5v2f5ohvQbNowhCkic/FFvU
9hvCaR2TXUJ8Vt/dmkrw/bKfvhGjYrSTAMw4dh5WvMw2S6sFG2Kdz5vwk+i3UNk9
1Q1owfZ8Pe73NB+wO7n3fI+FvZP+YLAg4Y7U3OJlFE554mGGDHfkQ1vC23W42AXu
hNanYR/ASZnQpr4/9OnWBv/i2DaMk0ElkzeeaGARUMjGllzSfvemb7i6mTMIpG7i
TcfbNsffoBOUbn1KgsIs6w2Z/1OqAw42BHJ5oLMFywkUzpJl+yoKgZKhH8V3rH+8
ChLQ9/QI4B0M1qDxKhdQB7wjSb4hDGl0GLLwvdGAHt3pSx7Wgok1QGZRFiqkJ9lx
kdBDUsVIxNSiv6uxG1FJJT293sXp7yi6dxuYMcbf61/I1TdZfAGj4zQsZsj0c/p+
dCvnTZBZHm7W6IJuOjC7y5pu0fDFbYY0MVjVc48EFIqbPhheUoPKPH4SVLo1aMRt
C4NQ/0hAoQTi0rm+5w9JIbINW6LICwv6CNUMP4pzI1pJ/l6dJnVvaDPJGTylCI5w
ieU7nJa1i8aMYvpzBUcYnaeUWBsurwgyRFSSCC5tbO1pTVw5M71ndHPjKYzlAbeT
0WS1bptOyXpOxSQcLoYanmsoMGWJX7qcHpecOFHF/p+emjNJBBwyEUULuqgXVAuk
3VNS416E3oRbkyxACrFaxbQOw+hYR2z7bPUf26BthyNapHiYn4KyFQDPBCbdMiOY
mQKgiGegDwAxVKZvto3VzJ1SyfoXa4TRdGXFk+wDjLWUfKWbz+n8srcOV4GRsZqo
JgY0Y+CDUQfzoICoAo/lz4q5O+kK2RlJgGdA2GOwEHLFI/xcggVMdsxZpHpo0JEW
LpYuGpE6O56cE9PGfw4sqklGAlcQKKFBkv5kSlS7EF69mOpkBfcf2Wx7WFIg+OLw
zTJA86gBXaFfvjTcuRiK3SdBXwJs5C9ACccELbnJNerGcYSYvpHxAPPXGp/Sg3z+
Jr20qHXBCMyZ8sEbgG3FVudR7sBptUG9nNPGZcbfo/Gy6OXTCtjORwR4SpgA2Qk1
RvaaSgMdX6IJdhYNMO08CoFFjo4o/1HjWji1KKgBdFEqEI2Tv2N781dqv4Bq66er
R6Su3t1szNHEG7G/bCkvnOHYEiyOaYWIeHogmDNvivaIcQ44v3ktaEsZZT5HprKp
su/yhcx2TbR7P3TAw0plF6j6dXtBatedh9El5UNcmzWHNfc3uSfFvRz09lrxFHAl
fgcKn9tXocebKcdIKiMqWF2msQv8O/qQ2Jfsy64nGKT321APVfihZForDB00Tpce
Tg4A+r5XxCt1kAuPNd4ChUTxRfhsuzUWGiDKFQvGVmEjhdAUgqax4J2XMJpffhF4
8EX2QRS7FFrEViW0JYu6RxxtzySP/A+acjzUST0W0p8VA7vn4okAs4p3054XyVue
I7LoEmR60NXpBKejp7eclbfYDub5b6B/RdKNqVG+LUG6shJ3QwhqcqhSsfc1pJ2d
UszSQMMMzjdgzoNEBD9Q8K7YjfBWrxoqQ48/e+NX0ZGTh+nKEtPQEE+Wgt9m/ge/
BEE4oVKw8E3e+wea67riNlMYhTEc2CN+wuZIB/ipgMxgWGYR35h5s2BkUt/QJlZK
qbrPqb8xPwu8wwE95SWTQZfhJw5VP7L1aSqkeIVTAjtNW7dHksP/ttlDaFmLlGKf
Vet+acHnLlEhbbKW1HvXkTDFF2g83WWP+3tcsOMi/1D2AmbJ1YIknN+4kjq//PXM
Qm16vjg1at2aI2IkT7V/CNw6RSC47kCzaaaQ+PMmn+COHermJErTT+afzoKISCal
H+86aCxBqU8Nxnn2pM97Wmif4MeVm1WKIyRhAn7sukEY6qg9x8cpG4cKBBm3+siS
N7uavhTGjOJpYCp/q5yEkSbd3pq1W+6yf1XXSBsXUCCKqrEckOcqe5iG4bh1FI/G
mHRnAxU7vqWsgge6lH8S1PCVrNZlQa34MnBV2BHnJJvhLVGfIMcMwFebS8fVoAMP
LtJaqKRlh3LBJZex8L4y/Xaf/+AhN0oSdbvF83/MDahWJHh2ftUJBhsTzgIhUr0K
mlOJ1/hKHZ/4Jo6i7q4mtHVToSfgdbR43Xxvm2s/si3tD1jyPOBeFwRbr4hutX6Y
OR87FY2pZgoniu+ZFJ+kT1hQdtpVIMwkUf4DeoNOtg9OZQoHWBvaPmeL5Pdctwfi
hdQfKoTRZnVkyNcw7xjLcRzlur7RlTwQtIp+nkXscgTy0dmmKzNtzFWyWGWangf2
tS1Jk/hrDZaIL8M4jLITxSIjlmyk2ZwnqgRAK4lRI/5OYDbKD8j+0eExwU1IMeJm
7KzK2sCAqeG89I+i1h8nyqLyMMjaX8umOZsfsJ56vexD6ZrftWvnxhyupPl96FVn
xOSmtqHfXAo1HEd5IsZRKfT+0pL7Ou31iWVMOl+S3LahaA3FsBmBAbmsJozclRET
VfNYHffctikGdLsf35h+n0vwLTA8cToaq2fE7sv7jm18/JsRJuwOh7boHZtFX9UX
+suzCyQUt0UXNdYjjydtzDM5mVpYVVWAlb8ux9gUhG5+Mqg97Hhm0rzmSOe3r5NL
OL1DDCMAV3jLE/TvwDjzIuN+owp9BD5ESqS/bWjvVuM1VX6DNL+y8uSriiZDJrCE
nCanOGmp15TJoyPCTlK33TYuWceVPk3svC0C3Pi2JblzbjT9GzSam4sBt36Zi3jk
MZVIddeNCb/Mpq+F+quIli4OP/wAFpZb0RHkffiCsSyDeSOQye0YF0jHhwCwms5h
fXJ/Qgc2H4vcR55iZrPjGt5w0AuC1vL07s8EVKszaLgMBa5hGlAx/RTk/gNblhmf
XcyNBf8UQwBc35mWoLuAGDF84vpmlaSSRBesZ2Nup+nKfbEHtwxQfWR398J/5tOu
vrolIbtoWYXC5JE38IOVQ2CM7LPvrBSQAkH3uiK87iVEDzPA0mB7IcwlVPHGApQ1
soi5AYjpWLpjmg1v/PwnunaK5HaBavh43TUPBFBtgxWeO/PwKolgMHxIRXm8OUjL
NwOOEPeGp3UzU0axTVL6sTGY637A4PZa6acw1ZN3RAxhqZ4L3j75Sdy7Rcfou4da
cXS+MWj/5RAtWPLZHDVG7YG8g63d73pOoIyOc+YrJNpmD25xmrRlfc60JJINdobE
PXKKJnz9Zco5ZHu/Ux9WnWBbxV35bbQNlzyS+m28mKdKOCSL1EBfKJBwPM0OYnOL
EeqXUUMvi92mKAnl8OyVrCUSY0BIYlmREl6Wek9XlhCvFqUpmFkbciNh1kTXFgE7
RlCDdd6xNguwB8R+b9yfII9PO7ldGYVUK5MvDc/gMsqzQwYg3UmBqX9u09CFZP3L
TPpq5f+borwNoQJRWNV2Wkj/kcxbBzcVJPIxvQixEp5vlJOa21saLuoG7evvijEx
Fc642Sao5z2/vkFaHJ97PjgjctmyH4OYSnj5cGKDk+ByU61PtlyB3sxwnCbBBnaO
QEp5ppLMiRYwhZAr5Nkq3ZhoqXOFLVHqQIRupO4/mTRTgXZuw0n8m/CmK77tLM1L
Vz5U0WYLSVObsAIzM/fuGS0TWU61bViljq6GekMNyWlB68zVsLtGAE5uL1XCdaC8
SD6tuA16BzHzLqoOPPd9DSHCdXAe9xSzXklL1vtTAEv0xjrX4C14gQynYESCiI9I
UxeKWcMCSmiSD+i5+eAMnthvfH2PfCXYrwffuLAt2VJ0bIfmSyqBf9CdiYbDvGmO
qIJ87A7jPKSgnsn5ZJFbfdTkxxZ20eWy5d2TBcZHj2LYhMjbKvVHGDkkngnQ86S8
t85QA7FOvvLwoR2V2e0I8eBGszp14eaX7us9jhqvpSLlwfd3RjDcTaZiA4IpawzM
BM7W32M4jlqCFoIv08lJUmJ4d1JrAImTPX/p0zpl9WTT4r0aJ/oLPW0ihwBMmD+U
rho5ZkS1Cfrvqas0HzOZ3oNVyuuZQONX5L67sA4LsZV+Nm+RTykK3eN49qApgB33
KVUtL56M1ceIwg44jPrTDWk5jbhwrGFO44Ye9v06wZk7REOwmxjxunVyB/gECh4P
JT0omNIaMBT+ES081s6LMFO6RQ50IvRZM67gsFHz4LD5FD6T4utViLzzm5vKOWEj
OSGe7Pd4zbK/3WVrt0sizVZ2+gIKXDxxWZju9iDE1AQ71vYYwArPQU9tnEcFBAyg
BdiAJLcMWrHz4sijDtiGMGbVByBM1bSWi1nHDqfWChmnERnYvJnSQR1yctUsTDIr
pE05d6/8pIk10YULc7DzyC+TBn9VBWjRJ6YQi1QV9wJ7Qq7AToJnZJJ4Fcwz9AjR
LwT+dFBrnDPZwTHLmqInx9IIBhYI1oIfvWA/ZOsdK4agalSN6wWhHrK4mPJYCL1V
s1FTSosHW9h/Que6ZKZPQfXELub2iNyw/HERpatsJzcvtoYk3/Jv+aa3xueMzaJM
LllX+hb28eQzS4F/SZr+sEoqPRrSR7y6eEynk9ciIECs8IFnq8C9M7NMVNqyqDZ6
Xj3PnI4Un/upZ44hfSVdj07FOi3t02OAzEo31bpQwv8ErqTzJ+LqFv7iACsNZfKN
ZakVA9II+6ALNJAw8jN96on64ZD8sVu1cBh3VSBOgdiOob7kZJsnLr6q/3lYOjGT
EH+oxWw7pQ5TtbP97UStuQw1haeEVAwxDm17c6zTj/vUY/PVInqxwxVGMFMXD1Tt
tbZ33eq0HYZBy9i+Qf9S6ipl2fwdTnEyntwlNiYH5C2ed+dYBQrhFvx+GHJnITPd
BW0lQ0umPva7W6+oKqp2uqItdBkr7Nx2V0BlxvWgDZL36XP72F3cTg6CndIcuOjs
qCDU/5QhOWYrGxWE8NjQUX4wq43c9S0731vePCI/6B6NY0/3sD/VXYaOVZp5D+l4
2TPins+7qtL74vN+3g0afX3hqCTkjiKBsNVqI1O8X+WndFBB49PpQbDz5DgtgNNt
Sj008FmFWBAqH6Ckehu1EmKlkd7Iy+AOJiB97CzKDOUajpjPuNyjg6MLityX33Jk
6oHVq0bzHYcCq9+hTRWfBRaFv2EOQpRDyAy0Vf8AuCcjlWGTJK98bhweBupHPPjO
/p5wRYnIBIhP4I0HrheVgCaUYjSnsZuOU6P4U7pM91e0RFekgo2ZiK/tNr1fOGAE
ie7Bod0oLk7XxodnKJz6PysV9sxjAMDb2MWBkuNh/aF5t9kUMxp1SdbakLktVByb
IAX33BjB6oNtQbZuhkuPrYEYGEoJlK2rRiT03XpsxgqkrtBBh5hd2Xz60fXW07/W
U648r/SVdbnkmJSxyjZYJuhcFe4EB7yoryU/SXuB4uHsEp26jjOl2ZvLpxQb3+iW
uOtQapQg5e/67baoQaqtKOZtcHN5RTgd1l5qSeYpK+n0KdM9WkOg6pJ0Vo/64qzn
vfiWiDymyjBk1tIdJlbiFj2aObxiAB/gpYIOlTkDwjAEn0R8UqCXJs/Pl69P8VTC
Tc1DkYhylOAOjMM3QeSUET1A+6DIGshLY6oz7zI/8dF4MH5CP6difFuTuTuycft/
wsCxXImW9XN1E0nMc8DbSoO3xgWYq+8IFYeajRBY+Zs/ew00WMGzvK3VDwVHTPnh
chfyccvQY+yVsgYU8J9v/ogU0bcTmSyJKLgo4hvG677pGHsNS7FHSoA6y5eRRLQp
sfOq/Fhst1qToZcVD+K5bwTU0b+M2snzl6p8XeqLqpWSUzCu1nYenu172Fl1SHoE
siGL89nrKhTUudsNd+e8JxJAthWA/9wZip0U6Bll5Oxn+JAOXnXQ8hu1DfVM3wLn
5RtUYoUuPv3sYix5U+TV1BW4sx2nq3aDgzhWrTmdh5R675LK9DJmvXHoeT/crCj7
+fa9UY/Mp3O+0NlG7V1JfNnPlaRWpxOyGz0piof8g8PmS7jQZY3OJtXkymheecdH
MKin1ZLKUf0PuIj131gpC+4Rc40vHf0PsPZDT5xtqfZWSgboEwWz0ZDK428qiymL
HLKebtYKrhuvyXvrQGnBHGFvKIWsWYzu3qb+V4ZEniizUlAOc8WVknm/FjUvVrol
6RpXbBS026/vnPQ5/az+Gj4I3lqSfwdm5oLKX6v/kuWMU5L3gKNL1nFRklU03OUJ
e8FeQpYaDdLa7Vi/Wd+PY6yJOmpY73WWLTo13SEekdaZ38Ylnp0OJAES/vIVsxTj
WUCC+QglOeAVC3KZtwFAxvi17f/cEh3KQ9MX7V49gmm15O+fu5o238sG4gxps24q
j7D98NTa73kiSs/TMRte1xgo+TrHFvd0XqJqu2N0Gd6mW5j/vkf7Z8Eg20oRYIyu
HNxV4T1a9QIh4kpkoQIX2hm6cCNIyFyRodi4rLdmnhUYWCqUnFK6e2x2o1seRPIa
pPM6wTRMcCLilwjIoEItCOtrubUdSzaIekXRR9GoxFN+Mj2Qqk6NtoO+IMUeiro4
CrXRqT2kqKQlML4dkmhIazEiaWqWQCpuNVc9A5y92mbaOSdMSCMwK0Z5M1s/CyQe
8W0r5h+Mhd0mix6+lyW3/utREP+Fqv0wiHVPApYLIpT0+E6DwW2rMMAKpoFhbi6d
vBM3WBUm14EpQzlcRwv8Yrj0InL1GzLYYkybiqZUB/T0DKjkyogxdGroRTFjA7Q2
0mbxkayEJu+7SDp6JL+mYa5SETXXH4BwrvRnD6hZ4H8URP1nZTjhDbMba8dREkOC
/xIjb3gNRBCBpt861tFOco7lZqHRVwBjkZXWngie5ehbeuqnnuvFehGfRrqn9FUB
wcgj9l334wVuWXWpIB5JmDzZVAVVinkGuJL1OXvbM5eFEDwAJ4pAKhKNlTarolZF
zwb2sXuWvCRNJ4B0yltGqxmhhGDWafiCiQOiosUFrbzSK0P0gn/yLPqKJYXjKfHD
ZUUO8OEK50TldGQTO51vM+4nPVe1CST5v4fCVfgofQD4rqfXVPzfn6U0iPfkpR27
oouVoEnYJi+qV1hencBxmiW9AeGMgHQpNXbOtZM1l3UqTxVw6t08gufQwCFD8seS
lCHEYVxAYKfYoWq5N+ptIAS0gAuy0uC3oKoi69z3xXMhgmAe+EV2iso13lYLe6hj
7JIo7fNAA6XT3uFFtjWPVOZG1dU19yjs1hkv0WdUbNY/elG9apl2Y3QsJ7Xj25Cq
eSyJy9HF845HfKs9OWW34EWYTtJcehMekMsh/2RQEAdG3uf3FI5L8eG1azJDAqaT
arl+nbWTV6tmyS310eIhf9rlw436Bb2GTIrXHueuFYL0s7Opgixyt4IIgBCmBaTz
m/NItAIJOzBal8XIh0ija/WizOQ3Cn3B0M/mle/MFHxC8RruVPIBpwVBEC8VJqK7
gtpYSfIfw3eK5y4pSPD6p+knd8nXTne22Ll8VZrHLwBUVQQ+rXwHq2hIIGEG4ttH
Rk7yF3s5BfTAydEAdniMBHeB6dCDmaLPLysh7ruiTM0xE7ksEpZ8LvUtYdtqxOxG
bURbSZQcWQ0/po290NKkv/hus8pULs9MfSDaQCu7gbFfzyxyakp/1+DTLFCskG0x
rhSbd1CfbpSZG8p97Ew4Y+IVTplSEFa1JARhgJea4vySFT5UfC08vyYRaASnQ5P5
5UarmW+N932EW2orBlk3Wmb335O9mF+Hi+83VapqPHNxQ0v80lOfk/efYGdGrWRf
KHia7sKsDbwUt8CnFpwawqMA3BBeT9NN9+tAcivim2HkZrRbWvEhvYMz7irtJ+mw
I+lz6pgtuxf0CVT0w/MKx69MWglcxAfU8ymFJYLJZ8N+XUxXba12HutCBtybb+wg
keMzLgeX0v7M19//jRFBT4QsoEXrO3dn8NKyzlSxm7Fa2vd5Vo5eOwWex/o7BLWM
2P5F2PI1y0evPFg6qM2pgpvMXe+8LezvtlSB/Wd2TrxTXMDbJToPSp+awqiHy6cw
t4X11KHzgd1EIKE+RWgA+vYIonaQSZilDHRSEMtqVeMWe7N6TTg+HxCLu/vQ9qNw
FmLYTm26Uh16GMk8NSXj67pKSXbmBmBOARdXJXRFiUwtuReDdvXdneFp4VzO9Q1A
qu7JlLpkUEDB5xLMpMRUK6gl1gTuu8hiK9hihq2PLs87vh8yPXyFEJtiHBzN2nAP
dVB97AZuZRpGTvBLhLk51e2FnlvljByIui9jb7ooOt0TPof3R8w7yfQhpITxqcZo
rh1EDLyqRF3OlZ05R33Y2/B8MZ5SEesxvlpDUOuGPUjyfCId7Ew7eap3M4Nuy2uP
xDoZLfjAMjhHJHvLqn7wjsGujK4NX10vxHp0Azyi63+NefPQ0GqDfBoSnP+evtp3
QyH9hiVkFmj4qtWvCQRiw77oHUDzFW6h5Cx9nz2NmJnzm6gdn79i6shiH7/HL/8W
rldlUz4nNaMcvboXQh2oIDgMDci8zwrPqHJrHto+ScfScHbtoZx30kDHKsQWKDVK
HdyTjA+CoIdKWyHOvb4tNU5DJFVHmSdok58yJ/rb7vPe+S0R4HdleH0W9DZ6r/33
doCtyie4fLLMjt48gJLWOzj5QHpN1udrPzADLA43zXnC9je4w+ivCJK7b/+Wpivx
U6Gpny5axeeEqfcZyUPST4KW4IQHHH+q1lc/LmtPbpM+SS4f+oX9Jg8fN/ZTrf8F
z70QQOzSQZrQe0cheaAtbQYR7QvsO9yTEp1UiJ4kxZvNPb2bGYPxN9dudd//p6dm
1mL159IApRu9QTJxfxXhOB1IYuhq6h9165g91+lpXTf+NyVZ/eD38yvF0dyYkf2Z
rL/5S1xZ6lTdDYIYKTwJSDFmHB8pk1VS4xiWPeg/vFpVnwHCxlA2QZCdlENk2+jF
MBjj1Bqr1u0MI6075NfGDNfG0dqWGMMufk55BUO3pkk1SZePtsQhBn/EaHYRfQH7
9kS914zfqYhbpmRZMPnUUEPlBBguVaTJBFJtPeLKZOqw76VouckMxJAtf5HtcTTq
94of4NkkQ0N9DCkCo8BBjGaBWaken13qnCKCaPz+v3TQatwmWhgjrVBkPT60vnR6
enu/JklIA95RRv0F2Eh6om3bCijdFQmkoS5S6WXNRjUC4SfCWRL8SUCIRA+W1zAI
d+o/G0cYhx/ATZeta1q1wSpHT3AgExSrgdCVk17XEhVKcpyajGmQ7KEi0Fquc9pD
XK5I9AGMcvzA5+GwbgefHItOGqHtPyM34nyFNZBlLlwy1GpfP+0APxaZ2G17XPeJ
orAHc4SgPVOR08xuCZPxQZG6UdkSqRB1RfFjgpYNwD1u2T/ih7DqyPo2n74aCBwf
qjQI2C1hZEKhCDFJMTJ3aMzB1A4Sv4/qaZ3EtAq+n7NoL13H6mTDegFdN28IRRwG
J6mAAv5grLOrI240zYkSsCp1ID5JryvT7zca6Nt5fKMgXterA9QfrP9ITkCK/uUj
oDFCee4Cfoj9gFlN8RRh9v+iUWx3GILYECf0Xgpu7yfsdT3JnXFC5mYuPP06SOl7
iYwZ8NOUHltI9I2NbSYkFWiQkuRysEPdJGIDib6wU929+CbyB8Y1KzNhflTpFJ72
4IlnALu3F/xPePMWPYkMZ97aF2qfgfw6wuw8Lps2BHB2KzBXzF2coJ7lg7GOqaPi
BxynPslmGiyyArqds9KnY7Q6Nn3rWIr0qQWMyQl9CNgWoPDk6x1b4KGT/7u51VVc
ngFpizaO1YKUeAxd3YQ+vlR+BuOTHEwrzBFxsevaFIvuuVIh5zmwlTaGM3J8RKKG
2U8O+XneBTcUsFX/zomiNpxxLtFQpikrac7Tp4A/bSuYSwm4yXAQQsZ4f/YO1UJ5
HSedHbR46jzH0UsH+5L8uCZvWRB/G/I0EcRzsswMxBcLBgEI4rcbvrY6HZMCXrtG
J+zhldznX42VCUmSKG6BtYRsGhKmxtAl10qTY9buGQ6r462M1p2wKbyKrZeMFLYo
jpgZGwyb3ylVokxbZZC+HKADVYWr/uW18DT1k5Ix+q1RFhZT3VVSS4YxAWdq3PoI
An2S8kUZ5OpOO3n+dO0jl3wB+CfrxS+yJaPajdR14zGXT4fFxvJnLWuID1kHItzr
loC5hdbTGozIL5UKyXgqNhjyldoCDqzGw5Ilr9uL9LT4NAn9xl8P3PPFLNC93kAL
5QFXaQ5+gJxvIEKlkIv0hkd+kI7ADl9bLzd3wb4Gzl7d24R2743W72LKTa+73pnq
Psc1wDhO9HqZaLxhE0V+GZ+23dnxg31ZYFEF8e7jrz27A7VlT8VJ6BrqW/sUvIQ/
A1YSNHIptAAj7rM9uQCSAm3GmNnEs77J3Y8dAs6bmBLLf/WOw1ZCmLmCquQAIbrw
i+IW3Ze/7rogQw9l7+0qObMM4k9D4PRoZOUR7H6W6AmmItiq7KwgNhJjBBexwIxc
TNOpX0rmQ6SUGNn6NPVBwUxbubrQBWXNCC1+ItPresAU8TyzXfrBI2MBdSbjWiwN
wnvk2c3ukRH1lpZ8sA20Yw906EoUxD5n1p8dwvpC58DgzhP7QRDgwIsg4DYWuapf
2csDX16hsOc8bbJWNL0xajOxwwsXRXfErHw01jek/BV5CzuSTePNy0+W3fi9tkIg
ya87fg2HU1h9h3ohW9N4GD9Ka5Di8xN+1BvFrUi/nkDjRJqt8z2Esd2qK/VGyJme
rf4wwUX2tMpCLFPiH8vjT4IhB/L+qcHloSTTtSSAhE++bc3Q0m2xK2W1v+FSM974
6rBtruz6ZxPhdookrWft0Nq3o6MsHA0AF3o/Lx5XpJsGd1nW9PyyRs3ocknKIn2U
aVUldhDQzwyFNKahdb8FNCpmZnflvj7lBnq8lagVWWNRN6zt6FMapmBPFji7nLvA
zurFMKs93cyA0HI5QVGDhqF1vS/oGyVTcGpo+aPnifl7pRVaFJ3bT5VBlHwRhJ4I
pVRneZKCp3Nz6mrjeIbPcDQdK6gN7QYaoI9p2ADxmTm9l+tEhqSTDqM3KKEsiHS1
DRTLdQtCpEaUqIPoLCeGQS1rOczFMwpdEIKPhF1V9EMGsV4jSOcgpiMM00a/zPF9
PheUdh/yHBBkdmEfS7jOyv4oCTopbPe90RcbU7CARNgQRaEfSZeWgIoBx+vJ1QBS
TS4CpgMAEt/el/7vAy8pNYyGa4EPoEWd5V6wuh8SfMLhFjtqsL+9+5CMoy5zI4uX
VYtYi4vZojGa8yPyjnNG3sx1yK4N+G7fz8u99MTm+K32yqrWxSdC+rK8z2ctASVs
ciW77endY1su5QOyxDl18M6otC3rIrcdHHo/nS9jXwC6jEkDn3Jomc+wB72vIMFp
VJlGgjdTbviaS/Rgp5Lfbn8eksQSutSUEjRlfGI2fIauQ8HCPeRaxaqJd+FU4g0o
7dxOcmjps7bVyhNtUlhxoviY4DO7t4RaZHGCKE8XopQh4eHG0vPrPHqzeAFJ1NXA
zu3TR4yOo3zOCmylLD82jznWrWZdJn1lfFdaHrZ4TBmrD4JJObM8WcSVJ3vLerw2
9uHZC17MGrb6jAs5VGJ98m9N9tvN8fClmPX/DDrMA8dnx2oyQ+yNGQPEJTali5RO
iE3IsYIbLzBrghUBaNnssuNa6R17UA+hPf62A99NNMiMvixZiRXddIhRqiO+7FVO
Q1S3I9mD0Q7G61bpOocOXUW6jB4fb/gEK13islL7eNdd4QPnqthgI0fZmLLpgwQA
Tew6aIszB4oy+nPxzrUYoMLOjfIQJD7wy9UlAJCjHZMbzzq3L/X5IZQkGnKcryz+
6AdBzYyCdCm8zuBHIgDt/QzgpDGJdiRtoJ9mL2QoGRG6PnGq3zCh5rlwtN8bnXCB
BCe1VMEGrCfnfRuAO64IgfObyqEsa/gTTxqiyP2vI5dEbHRoNHIiqG0t6g9pzhyt
GMcxiemOscEhnk5O/W7kyTIGwqe65/V+UAY3SQkp+5+5iDSjhuIhhORyhU0a0Men
UeHYyNIHyXerTPPANAJi7EyaMKFsxWtcJgKbFSu6dhv8ns7dWZG68U1v5WKGSVV/
kx0SfO77kSlZhMMqy1KRR/T9M0fyRRQm6/HeY+dqssRi3jIlO75NmUBxdqlvVHzX
ddu7aWtffkTXPvnfCYQV2kLI3uTZi3l7HmtSn5+tAuPMPfBX7WvwaeWVoIJzE9e4
/rBBWxnGzoob23pvdS2qAn9NbKFw6OLnm9DHspOjU3X9hxdkYCiwXsgtfLHd+yYk
ocqN1O0S6PjSSHSKMIs/1wgvCDZ4ylCgbmyW1HbpUhlVJY5kNG2fU0OOBhTP3G8R
X9+nkMWWfZPXCVpU9PtlzVWQkqnM6s20T1rwPrJGfKhVAnScCxsfjiI87jC/6gS4
HNzFItuxLaAB5jZN6iHvgtvPBSHDtSA1GedAncFUik76Maf592EUeF0DSsgJLTwn
NAF291K3o6WzXkwTVM1EulEgPVXvh1dC8/j9EX9Y40/FCYpeOOgRNnfqJI/d6fod
sagOmHNpADstHZrqxv9n/6ZhzHhvNghRD9I2Ype12PXsLgKKNQNEsVYDQPkIxclB
AXQMF8aTGUGwmsMjlrcI2ZocdgnHjxRx2H7o9FMsX0Q2eyAkvH8x5CNc53imCsZ7
whwXgtOt4ZJ2aqpVy5LgCvSloAzLmXRdfDgf5AbZmmvdqGeUFJKfBapG1lTsargF
RovEvv74oRvIK/7ICQ9YRukWVvORz03dJj6dbd/u2LetZ58ACP+lzpzVDX3wWl2t
Ye2B4Rrd41oVBMWbEFQlQ+BaqjvQMH8vk/zZJdhgRZHlYvm9S5vtUv9OjEVxgrnk
GoEJaIEk0ZAg/zv187M7Q/KeVjj0q4WuXAWzz8M9gB1JMioCz+zm3kkeBWYxbIMV
Y3CVE7prJom0POTq3VGJCN8nbyukQ3ISzzLWYVDmrgPLEqk93VvLAqafFQZW6YxT
Pkbh0Lc40kJSx22LZXOpiDMok27N2irsvRLdfUq+iw1RY1JUhWBG5+rSGV495l6u
B/pFJhNq3bo07P5RQp1vapqsHQ3KbQyVU9y84aUZxCiexH5xlkrC9mLKw6tgrHxE
dEJt0RJPlEk0LHVNhrhBgDv9Nn17y8tCX+Bg7N8wr9Bdfzv6wN5ZJrKzjrAAN9wg
b+XoKOzgJ0Q6hM5TejJoNF7ny0xXFyjvAz2zZ6EC+qlJEgAt7hycWApQEswFPj0o
AeVtO4z7/gpTTtNBmQLTWYk78cRaKC3OyqxX9I8UqocSgso7p4Iu1hYAVtAbdWkq
ei1gjmUGRb220W30r6YVxtDF7R3dK6AA4ECT/2eEdzK1cdAFY0f97DseAKqDqfwe
cV/uJzlRj6Ix5u+PuWuLBb/9fQSYHkKGJDSQdHXEUH1J7b54MT500sEUsoRbkVCc
c/taf9dinQOhOjL5dn7XU2/oRMrIlm6TA3/xgn71cB51qZaC8zjYnMxM7yWR1l1v
S8q+5W6A3zu6dNOGSvR4PwjIypMnsrMxaPhm9p0DRu8LcHMB/rkXcxPGkvmGDJ1T
Xg67EWx+wjhIfBh49/u4Hp+mwBiUpVyul2qqolVdIRbKeQ197v+t/DD6OwRqF7CS
ywWFapj01vH/2sZyR9yRuFqhrFk+D3c9qHx9fMnVS8vicXSjqiqWQzDbrhhHVNNf
h+aTc2lb7f54CJmeKjS/o/dDXKwxDANjLkLLoGzktcW7J/NXWG0WFeyT0z8f2M7S
7GDWaQUTinkzxPXzHVf8ooFgwc2dGFag0Zk2GWsPujLCqjNz3qZqUzSVBu6/92iP
TsfK/YsV6CLi5LgJVqWLIIuzZdMMseJULUq4GIXXDHgSY5qic2weigOjUhppynEv
kfCQKu2Elmo0VvZ3r1CbAoDRBo3hdNrHTs41d/JyfP27d++9XxNThqREv+N3NF/R
xKhqEoV8j/VcNkAsFB/VyLFfarC3AGxHeIh0pOitiEJyqc+gIaU0tdqRYdhHLICE
5pkk3iwxyqlt5ucit+B4I9e/rcBaSamdAy8iHk72NOoZWx0frE/eTYAThi2/LUPN
p+qtndFYwFyyeSz4Gsw6XYkCobAQczAnKgbZmIxkOUwtKm4xXB1tfh2ictMrDsU0
q7qfZg+CTtdqGtGhv5a49zxplNZZXj08XCUDJeXaZcG8AqS7Xgn5ZEt2G0yz9gaZ
ep3M0g9/cI/zzEPfzExOoH4qqvbQDSfilbwhUj7FDfqHDs6hNFUhJ3e8Cgd8im/H
Rja7VPNY57NDbWOUcgw8DDyNwkC4cRzFamUIrGtRZ+PJYInjAhQ1tjmBfNshWysT
jrF4O8+82uDbyK0hMRMUzld+K+VUZ3oZXn+0lp+E0+k6Anr7Ut/A27w68At4GTOr
IWMYpWy1RILNObPx3GighSf15faTjiOTw+S6vkJaeW722ul98y9m0A1i1tH804dX
3ykdc6HHozQNdhIG4rYG9k+pixIB4i5/aB8ngWBbVH1DuCc4Ym90xhTJLhFzSb96
dZCquJzFUtlWiX+hYSeEoJvjE9mZCOnRbUVTzo6RYcwQULa2K9iFKx1yNZf1Mfgy
oafjLOZgujioWSNngsaLR+LNpePriCOLVC+3X+cNZ6ilShGIMQ2or3lMbcMQnIbo
NBdgfHM0FcmKMdEUWesAUaAjT2M24qpkGXDE7cZZTakWY7C28oK+3p4swW+LysLA
wn7NCnMGJfgnwIx+cveHTZ8wiVOR63VuwCnIPn9cpzrHptMDGCipFhmGqw66M7LU
QvkJvCxaoaw6asNz3PXKDI/35cY6VmMT/sgdS20mgOfzOIhhzWM8PRl5N8QvUHFi
6BNbCHGIlmNGwuMaExE7lqnI6GnyQzRUx79uVBjen0Ffa1dVjhPG5i13yWGMYof9
CzJ/lwS8MXNPL0hUT07xDJM91pDdHvW+5Ylu1ZT+x9iog69946t8BVk7R0KUs9A7
dM7Lo0ZNnMaUP/M2RhjI0vOOaD1pBlNwMoxdAmseodsNP36cpi0xWFvZ9P8CaGeh
1/26ULkubAJ2vPZxJNmTxASeXA2ELjuo4Vfs6N1tZNAh3HdfVZ1//6MqxRWUuH4r
lgnAPrzEFXSWzF1xSLePOySkQvRKiE/WJZV2PmSeK28neQPTl0KeyyfJ3cCfEiOI
nFy+g615Rurdmdotf2a7yFJCx97RyX+xjwqht2L7/1lMc5lfiy9yDv/AJZzAIkQY
6olGSA6KFVKWW8JyWMP4VGIUh1GduM2T0Xq/Qy2eLEFvKYupYB+3JDO422wCyT4T
oTNRHF5kgFE0hkm6TTOJScPJoCPqMAWH6Wc8rLyX28pqsvMruLdJYmqO9WTYDJm7
M4Ynsf2g+suUBttjUPbzQ8nRNnIdVD/fROn+CO4J6hQa/JQ6hFid5jBexUob2mML
xJG097Y9Xaf20Hwh2I7+JkGVQk2dtQKQyPN0FKyw+v4yF8a15cGZ4Ne0aquTAMT1
wssPSYOzByqx1KTsYVoHw4RBIr70JmDmIEKQBsi3eOYY4KNOJXNw9tK8WSWb2jAp
YBToehSmmpn93G+/NJbZjFlMSc70ekCgRPzYbfjKY3KyK6uJe/WhDxucPnZpMqBo
6hjJ8pQswg6jhILKxPSPEaHA8GrrjI45jEAXFYr800vjPOS6xmp2qmXYyIiI/c1T
5xJJPwVal2zz3JYCX4XaGKWjHacqo9pS9rF9ZBEnF2BsRpcgfIUjkJWM/igZN3F0
XASy6zGlywGyFUCkF9hCdVTGTcoPEUKll/Tdc6eGxHPmxdrpADfQub36/JuqB+VV
H3alSAjao3wZvhYo/JXemllwFBWgddAl7bqKc0ZPt3zb67r5jC0+y40XrNiOw7os
bpprBCZrfgPupV8v9dah19vCjU4ijjbT2MTUs3jIVyMfn2WBDTK04Pj71vumjZJO
dIShRAohCjauO01qk/BfoXE2AvbAPxjd96hxjYlhNx0h72CLDSdNPn1EIEbcUq0m
lN37ZgT1i6Cdz3kNHXOZBZhXNrqKFMrirlFjUzk89w/1N0UYXBxgIxgxglEGayMH
y+GYXahExwRrMYhgUq7KR0sCtpExsSX1vq8B0STv7VzajmgQ8d7XQX3od3HGAgst
JMBjMNugGhOD4k/P4+byVPU9MZLwk1/uYggtHtE6AtczakTv595dWXx1yxQkym4U
UNwv09qiomxJRggOAD38uy85zEYY4Ly2cgajgC5lO6B/saFUbKbfGll80PeY3lia
b8pxutV9p8y9cpsi0R7GbUmNwfNHaXOQkBHzJKBgBeXX2vaKKjLPT2bYDLbZltox
1YYnlP96BbimKv1H/IAMhG8rYr31Qx6MGLtkW/hN7b1X+Q64u3DgDEqeYXf9uElP
QE10Tp2t4jiijcnVBOd8QY5ilV2X9RzALuV6DpFHsIBafuI1s66Pc++2c1sa4J6y
xszZjaIDwG3lZQrkT8x61jgjetYgA4UyHMxuYTKeLK+8+0l9qpGyaSSObgJIpENa
7gsEZg7mWNxqiyPb8a9VIrPAn7A/QRKScm65++nRpPl86HCIZ6iNdGgeFTlqIPIh
wmdDeFL+QsHQb4+eXWuuhx70NCo+r7mJoCrADgExfTq1W/LCgQ5QdWsJHtDGyiyA
WuQ3W18cn/TOlcz0T0I9TyFBEeCj4ZzPDbNR5wfb2pBaRYYZdcL/s9jRFPI/CSJ9
ZJCwJnpkiu3bOPExr/muKTdN+DzdjUqXAKHX/oQMgfmidgWDIQYk9R4S1VFUdJCg
F3we1JZSRQoSVohfxh9xVYKOlIV6Lhiua9gCFviWrPU8sLc6REddnfnzIZgJWWdP
C8PDrt4OVXDFZfNxNMJioFrrsKHqMGR+CTwiOKZyPA7YCvH7qXHl7JQ7lL+Rlwi4
alRWQMR3FXctBXgnJN3twLZt8+PjMfcq/7cOzWdiWeMQN79hTC5qL0hwy+k2tXYQ
Jwb8O+3VfS/QgmDpQpLqyKkMO0vlnYel9hNYjwcikc0H5g22TzbaeecuNgvsZ6Yg
Ry6+DRZrTDYqZZZx54tKpP80Xp9p8rLnJLrBOTNytkgreYPKgLWjg0KXCBQeXXjh
NrIuc31gWANYY6S6uxjaA4LWJ9GEMXqDFfTvBAFS+rgGu9oLERjHQoNlgBnxS8K+
00KrfPt/En25XdDpj5hPaAvrcRO3g+mKLaS1G6vqP8l+R+xIpDheyDuVBZ0IFJFl
21HLEeUb3/BDY+xUri0qTSJn6sfVp2d0IR3QAK40iDRslBi6YLT/3X4Bvfl3Y5Cp
0phBhJXhBVJJb9/IX+f5I3Eui9mZYDW+NEYS6YX2lIMMSqkAT5Gbo1K4r4BJjzJe
7SfH/lXyNTgNq+Q6+jM8zaKTe6PivAx2iaFMwewJYbFkIRgpAi9xp9YJYKC2pGH8
T+kKC9k43856T+zvn+uHeSNHQtcUKqFZlt37oB4HShboUVFezCdh6SWpHauITtCA
Blk9gzwPf6tW1oCGnhgOlfCxAmEbOM5xbCAWju/21eM2TzhMXcrIUtOXowH4zFWC
X01Q3SnySoWLJwtwoWutol5BMHGD4A08foh8afHQneqBilgXMJXUvFILC5fpH7Md
A1luUcTYHPYD0yPlWx9Kd/BsyOOfGzlcF4TATcKIAV1tIo3vlLR/Co5023hTIzfN
oAAXVX8gHOkcLeeJiZNxt14LkM/jUvlvk5q1FnfY81BDyDhNvSLf+NTsZYJjg+th
aGKeoMNML5Pb9qsduUWjsl94F5VTKCOtmvFCg90KHJPcKUFslne2T4/p34eUdbQt
0Q6p5lT68H933WIhpUXG/CwJVGrKFjfQ7xBFsbZrKS73s8HHWlWTtVrUvnnNyt3S
ki1dptLqBWnK6/JuVxBU/XFv+uoHV6XxYFIOAUBpAug0y/djQHfNHq8ztmk+ayB+
U655FqO3sPpt/zVD6/jg5r7l+X5mXloYe5Zsbqd/bVTum6c13Znju8n7ol9g4lRW
+BHC5Ykp8oJYpBEahe/2zsqPHKMSGDN9AWG6O922EDzuZQWkyHLqzL7jLdwb7bGE
NfFqRQjPcye0EA5l77d4dR3RyyxDYC+A8RCd0OU6CpxoV/uYx9obRmIv5VAcnQIh
DXkmnr3RxZAUp5Kj3QSq0jx4EEYaQRxY98rLXZHwZ3gWL/WO0V1fKDRy4bm7naiw
kaSnTb5+kvkWAiNafWkkFNQ9lf5i3e2XDznxFD3Fvf7nNUVKfUw03ZtHgyw8QgaJ
EcPXd1p3ct7LfJf4a2IDbg0rQ0q/qR8BdbeaQG55weRC50aNVb35sQ1ZkUgoiDt0
8WscvMomy3HpDFFjnd9kyi3/gsHChq4FlUwcPvudoDLjNLhp6qwiAHJhjHKXrPrx
gp/S/fE+E5nrDAvcL+r1ImnIV4luEx4zswuw4ezHGikepIIYJpXDVN/FLyx8EfZv
I/RCz4JQ6gb1mH6vn2PVk2I0zhcd9r+MXb6sxYldMGzIiRrruPc1rMTFitP3xFgt
KsUKR7lIuTJ1rHjUnAsmVN1TQfl8IRRl7U07n4aHh2GVX8ekM6/tWs1NWRmYz3ts
GSkyG2cZx0p2QQJEIRPUc2Q24eCBGvULnIbTmUkqz7wpvozla7JKQrXmTdijcM39
bWmnwk4CDdCaDihb7rGVY6qCISS3x7w7VA20jwKAODvh6I37N0r+3ki2N50KC6+h
wE+NMxhIbSy9+L6zrmBCZfGsr565SenOOIUdYPuOQA+T+CDkZAjBDXDLyix1OItb
YcYqbsr2yA7ojLKwTN70ZuUtloGpdB/3RU3XpKTkTNrhfkHgtQkai4awtFRIY04S
bKK+A1uaZ7oYOVFT0si+9nkoySYojqrGSGDxpquaQ41yA0V57KM1B9e1ql9C+N74
NJRaIgzO9u8Rn3a25Wd8cBHLr4WuzrTLSfZPvuJSeu2fUjBdvHiFBYByUBBqv98c
ve1bhGVj4yQ8CMtH/wspFLGK7j1uZ9d2UUflcgYFMDG5gLKCRAGGWLCsIFPt6/ES
WOj3lTegVzB4F7cEg7xEAlDtcmadMP6ICyFOMp6bIaJ6V/OneXdoJepM2rROYUOz
ViJmqsVCQzC718CS33PrvkDxj83udY2IFyx2yq0S9yzRRkMo6J8STP9R6Jp5ZEha
SLU+tLRCYs3XQMJr1LE6LJocwGtsnsLQGzhh+ENWTThtbAatj3T9/H6KgFBSauRQ
XbHnR+5O4TSaWxw2MCS1fRlcQ5Hqa3VFChf7dLA59z4OJdVW0N5OHUglbFvaLdh/
rnog0v1JhW1Qq1ziXFxgQXp75UeNTyrVlUeudy/8sTgkIDdpRAADXZTqM/zFf5wv
p5+w7e1EEfw5zO6Wb3Tm1tbTMns0Ka5tj66WdHEGWyZIUIAZ0fLNXVfaMiS0JMG2
OsyQtpB/THudbnb2DjgbUgBZcnAnnX+VDpESDPtTuJTCbX8fVJs56Zsxes4fti5C
PWjK2yB5ZUsNlmx9IhpOJnz4WMz63Fsg1JbcY/sPJj5F51UmHO7+UrXxEZ4Lfu1K
GjUXXNCW74HEWkIAmpmyY1fEIQI/nHtRTy/NbzbnvmQppx88InUqLtZZEhpO0+xB
MCcTKWY2xhWMH8kTR361o8BSyJm+ZsdkZxhAOR7Hs261FGVkAKwCswlzZ/a+EjOK
LiPZTqJZtHgI2uskEFr3PvCpTy1h2FbEw2xhI58StjUprOPx9ScT+M7H9D30DVVZ
o623tr9/Y4MWZwHqYM89izf3FneRLMYGDtI9V8snEvplNhDc8wEbQpiljMBBynJZ
qpcMywj1K76/BkpImmQxca7JTF4+mJuHjj2bjf2SdneS0DDKTnDAxeqjpiKPztzq
uNNWz68WyJcGHW0h1QD17yf/Gr9dk5uQDKmlP0jUI5qyAzFqYZCQZlirj/DBv+MR
K+bl2xemnSdYpVHR6lumY91EOprOoQj2RoPhsQQWxzXA3PPyJHlA65tZTOVSs+Tn
YjJL6TjGdMIVfuAk3ToaM+2uNi73WF9vJty9H9ZKfSyqoAiOZgvU/r/SsGo/c9E/
e9Y34c2ico08JCpzuhIWti/KYCV0ssvD+sFF3wrw/zlM+1MYtBLYvxNHnIhnntq+
LR+Ac+MHFgsz9BHQHNScgp54jL7Z1rzY9lVnUZc+IpjR3P4TSO2YOxshxy64zG4O
8FiXJzRsoeVAbqeZ5Zu+OBRM+N8jn4TFTXF6U88sAsKnqqxxEZj5cD2//AnfWiwr
7QyE01GmhUaOj5hfd4WuWtgU+PC2F0iNZWZQEmNL6IMH8RWTlGXngPt43pDqS17F
9m/gHdwkbFvzGnPzY42GUjVp9i1c7vKVMk1nBRabTYAuHvRSzmaoxRBHrH1qT/yP
up1MdlXKh+wGIuC2PFHyvHJH2R6/u2L21Zg/nBDMLlTnp0/c2KE3G2yX2iAcxa74
0Thb/jIgcP8jFOUKiBB/g4M2GcXBNs1oJ20mHn/mo5ytAtdn7tAenMxDMG23k49m
xj72DHAETUCJwPakttlHdZNvEHo63y9OQUl3ZPK0oVGYrek7HMCCSZ1xEQyHg9S6
ggH+rPlx3hgoJiY9BEbv2Nq5cgcWncfOgh/QvncW+x7B7/u6mflO7/3ZJ2nskinZ
Yy+DdVkax6GEMIICjvNgolWmLSVUg+aGPFt7cQNcmCgyBlXSmv6e/L+L6INcwVUv
sHQJdGX4Xxjp4qut1aggp5VbN+cftwNzbFxbBafoPOKO5c3rHO0k0yp0ffv3X980
zNP5Y0eihj7+UR9JutREnaofuh8K/Y4MkczZvSBSgq0kvAD8uREeS5ucKEkC9brf
JNyESHuErkIf0sLVtRe6C9NnvN3afQw0ahTEXIUltXySjaAVO+1hPlKjwhLsSKfq
Sm/Jb5MgnCsIbfMOuThRpTMnGTUOsIrSoTRWs0VVQ9GX0RVelHeJX2/rTwzBD2Gd
mS5JvxA/ngOSjVXx0wO36YYJPrbly1y/0l8RU5Iu4Df2ke4Xd+vt+kBWYIs7FrXy
d4DYQ25DwUaNdVNxtYfq3gT6ko+h8lEzAowh1rVtm/13Izvy9hs3DbmBjNzx6E0B
ZP0GvGgmp/O3Bx3rjquw54rP/Fle8gYAlQDyGngDstfyP0AO4ZN6izgUyQKq0w6n
Ce1LGCCo5EmfoJ/etXANSZcOWSMdbsLd8Ki0EuC//trYstBzlB1F1S/6aqsTqnQj
qLJq7Rhi0ALWDcI6Vf3QuvKp8zRRIvm22PFkI/w6EfcFcFlq7anxAeJxjI5gfEw6
JrAJZrAw5RUsfbgP8Zq9q13nmbn5awG46INax6n3vJ/xfWiUws6nOIdk9NUZ+F1M
6X2NOcxU8dgpCuUxx1HEslT4D5hTU77PT62slxRYzKNevPCiEvk65OQyO21mEPA1
M84sSGYqCjU50wLNaKt6bn7tia9yuXzJ9Ue42RHRcearNBX7CAVEtL1VVInG65ui
9BHfbbgsGls6LRHCutohWNwu6zr9auHJFCwOylhqpD1uAs9rmrO58JUAux4i9G5b
cHgdzkW3EYfkFHMoZMXH3Hfpm4mBJf0pKyQQ8emxEWA7EZJi95pm4JKhq+kQfXdH
pqxp+xsvqocIvqWD9KI+K1naEtVGmhA85BO5wPOv87YmgBuNfghTCMMyseG8jWZo
rlMbBUJlDCjNpX7LvrULfCjs8cGeSgwF6OMdjPlqIKtqOLa9EWO0bxz0nAG/ohvL
5L3FKo5plITCcE1VwHveGnIjkqsE1tAJP4f8RWlaUmB/75xPVAO71SGWxVspH+Hw
BANFxOEfYrs68oat9rtFCDeQA3k56Hb2f+/5+oVysEIRNEu7tkQOArEBsjacQnHC
kr3kqjlDtxmAJ61P9qUpNsBqgIoYENcszMiY6hPvZvxD0WargCmVgb6FJVgM3zvv
R8QEYLYrYMT+j/JQMrMsgaoGiu7t8qk2qjBha5a/z+2IeB+QIBnewdNxjSpT3bjO
IN5B5HaISv8AewTi45OAiOt5irewMYeQUJm5DdmMYNIE1f1QfqbvbZXEAETJ5kWR
F8g9d5t2ZtFqqxTBTuwo//aiRiEClLJEubjcD1bgiV79lN0e4pvvL01PYsnTBPVS
WX5QDX2rKA0sTXFgQN3i+OGfowd/NmU/0sPhYygGi23uZ1nEVjqbCHKub49vJhCE
LFcMUFWO6Eg5NZ/qU1CW+e4MjKjGQcNjNscXtRoZPEO1C0RdB7Ktel0HUNEdBiI9
Z0tL2eLn3FWkWGdo3riYRLp+1OGDNe2FPLiQj1D/IgJfoJCCpkibHrjdmJwGumZk
mCXQrO7mOeY8xwbpd7wungKpUvOA6GDXVf2BtrW9yhyby1+LRNLRmP1muRzynPSm
KltUXoGIwGEYE+aii8jSUPK/5fGLRhDjfsQa/WquDmeOnUw1o3g4hCckGR3OH4bQ
anfh7G0tf16dfwpQRx7DvalUDHSKHI9Rv9dD873/oJlNMKA3tt93FB7l6bIxHIYQ
xlzGRXuDV+xxaQKtw/bOzWZQ/Rykdm36/PbS2r0eSO0UysYo5YCvqh3aL92bXhxW
/bszQxTL67DisTZtQKF4B0Q0YioaDHrlwjNdu7qM5kERhAmhO9ryOXVdTbOBWMYf
cuBpwhk7EQeQ6urnvA479IiCG+IA669kIgAhFVYweJJeNhakv9PzKCsKmC6ZoNls
ooeu5Lra4KJiTmCJRJKYqNa/b4u6h6rxpsOyWZJ2UuyT/kfsXL+wgq9wqI971caO
trkdqWkCPq8+XuPDD0mi6LjG99Bc0yiAGC+Cs80F/PCI2Hv3g53aR1QcjY4VVLXQ
8+t18s5HjvSzxDAtBe7wGowJyDdQT87n5vYRCQd7videlZLZJ7xCL55MbIXDeCwt
Snvv+GTfD3DJ+6lTUqnpi74jrcRHIBJUbFxKxXf9yujhhHLHr935Rc4SKm6e2ZyH
rxWPuk5Ys8wFpRIMynwbxYcAFP3+Zdf7D5vShe33lYycfqN9h/TPg5tXQGNCT7qw
C/8qy+ZhD4pqCb4Xu3QcOV3CRaX0D3Z0gNMTgInIA8tbQfWUYvt9a1HjWfozdQvG
1sj65QSBGSzn/Jjkq4dP9rnbFJy17e8EiIjIc5v8l8sLiClWewN1mi4vCi7rB9rL
QTfKDitkh0eSzU3jnbVqznvhZXu3pnkR9G1KTkM2sZHyRenyIAWF9LAJpjVRhadp
N3GW4bNgcN6mk5zUir4ao+sTLN+kMpIO6Z6nBUp7fy0xIFk/MlGa6KAWAB/dH64K
cDxXV63ORjQyiGHubTYKDz2yOYjaX8MQ2wVF6ZaWMpl4LhXRCR3sXPcpR2FDZYed
LfTDHEN8iqOMi9ZFhEztTUm808Y8rWDfSs5f4IAzU3OMXmFY80115phE0qmrBADQ
VhuNbVYh0WOA9NhEG4QPfvBiioh1HlYNFX+LZQX+4Py+wx2REHILtJ4ZtGruDi1x
+Vk4b8xd4XDdo14yo11EdYQqdy140I0PFQSE7B2YmiES0gCDqg+ptCaYoCYx/wMw
mWbmWWOIkFC66PZK4/ir96W9SO/tdqn1RzrwHuL5MkTiSJYsWle+tQAr1Frwv4La
p7YCyab8/NjN0V+6SQF33UUIPMJQ8a4h/2OqcRNBfciXhH0PifWAHxMBqNiBMRUe
D7RG1gWqUkClCZ/P2N701MsobwEJSwS6rGZn1WWiE2Jw0IjoB9bJKlNEiwWVPJws
5PGkl2YjQWwtJjfM7n8iw391DLdOZfU8AyyGPaUK8ZucO1Rb0FFZZzNi6u476cws
uiBD1veMN30sayt3YTr4Ae5EmO8Q5NQVYhHqDg4XO0ZdgdIVhLNPofxvm1zV7s+A
2XIEJtryMORYI776hEYTweC0fEuJhWg+eDd0Ekm80rJ1dexmSv4EDe+r3ud8drY5
/HXQs2UMyd1otCtQTYiL6eHIZ2S3PxBqIxvS4NKHCC77KcU526ECeCjgNG7aIIj1
FyGT5c17ZCnayYfC9+UxU4tBQHRH+lY3C9Vwo82l9zZwdlpeg8a1M5Ktc33kNjG8
jF5oboBw9iE8IaLJLR+pocxlXrtlYSlB2BmNAkSiocOIodtKK3sSQRXwuWIkWKhE
EXQ99hQqc8JqdCGIWAE+q/MItnlFZYep+PdqAMIy/xlR0iJUz6pUyA4oRFklyjpc
wMxRp256Z5GBk2pUcuAyWZCoFis1mc1Cnc8T3OyaMYK9ycMQs6P7eFvgvdjwXpgD
6atH3dr+NUHL7w0bDhO0VX2kPgi0EBMA2NjaMnLLC60n31ZxmFBMmz6sI9Ot+4qD
CKMg+fWK/Z/C8ko3dgVtjuFOP1HM2xew822mPu45fZvbOIEMEUWj0DQydq/0AnRx
bDOdNnzpL4/x0vLfPej8WDtfIYE70i6tWauF/pBWVHuaDmpj7WchfDHStMttu9MM
PEJ25BCCQ4x2h45EAymvDz81/Zld/wwO126ebv4ckfaWGJXERnw7iAZOhzXCleoB
rihsL2oZeBtHrhmeP2nTw0JCvb8MVjwAA+PCOA8bHGkQQ007uST6Faosj3LJC24u
Q7iXqGzqk9Xo7mN6ofVGFUAgazcWu5dXWhxlKFUNKz2R6LqMgIvoXCj1C81b88kV
9mnvCDVZ7kQyuV82hsi2cqfPCsSYEk4mUuZaitZUPXc3XsErpSGZ38Itz5zUcfVw
Gp97su7rjo9hAtqT9wOGwYoxA0JDEOXaQvdY84aNAQTPjlL8qY4JnXTiWT5oXj4X
3l5zET10/cO3TmoUm9BrHjFSgCSucY5kBWYmHb+JFey+KjAt3ngnjzTtQAkpTk4R
q0FinFO1GYvETZPU4gqcve2ePOHG54GmgorEvb1CNHEJiBV8BLrp+XScHqGhX0Lm
HzeXXB4+AsVzLrDwesChtN83BfLxBT9fb1uUCTyAuspT0tqUA8nRUYDtIGsRNnPQ
zO20DRkBGvIqSmwDD+kP7iM4nrlW8PK9x79FD6RYIXM/S0DXs7ofFlNxlUHuvO7k
xtOkeCc3gq0+1OvhdFFtHow2pn29FyQTkdg4CaS0p8GLynAPCvpelTsPlT/+i7J0
U0GKEXFXGXmL18bzUCkOe0y9zVoxRYGCCTaMowKklsOsT2/ejNe2Z/W333LMzyQ2
SWWnoGEs+5uuRizYVAJlOjHdQ1fQ5yY6qDTrJ6OvaFc7cLKBuAwfMf8Mce+mtQlX
ecycZ9PgKMkoOEOKL3jNI4jbgJRVxdNxWxdXwTktss2L4OSDNG3U5DOn6t+7glfI
jUz3PD40Ae1BEB5nOUUCuKwZqiSFZDvMm7upmefzixZcd5OqGN0ZOkP2DOdY3KBf
V7JRCgEbz5jBsArpSU0dxmmNgv9PzCTz4oZWulqwg9eQMFfY4AY84kxDrSljRlt2
JFu5RS6qNPXGKqpY38zxe9rrTTQchFLR5TD4/91OLNL//zSKwatnvkz6BDjqbRoI
0vg/IVe9IX1ZWwqMrdmOKhIY5BtUKJopWH1puwg1Ph5nV2n3qH0Ym1W/mKkFogLu
E7ENDadABe6RWvkIGu+410deVHw9ZkRANx2NdqRiiB34Svr3rMS+EcSnoWppXkvU
2NS+MzUaom9JMqlppMmjMiIBECpofULqkvI//gsyZNKgoYJY2qRmO3k1cWzRVMNa
0y02TkEiEZvuJRHlwKitbRb0rr5oWtcUe+2cRCGHyBv56CemzweIwqMUkC6BZ9LN
8+kg/eqP96e37eyzVL7F+E+kGo53fWu4NbyKOzKt4z8BM7wBwOS7pjd6SUW8t3k7
tb4gSBXZWK3k5z55R/lfIj68izuflN3kPRRyerTrHPFAx5h22hHRQE2MbF7NZDd8
c+DSJVe2tTCPRSkgP8lMGgDZS/g30ZZJaGLPU2rlEp2cC+WV+JqTvZynzmN9sqNy
E5yFz24412+yCp4pJZoClqZrKVE7v+aQc9HM//okAJgubyG4kHQQ/K9R4c/m9X2X
EbxZgYtxsHfD0V/+wWK9xACiDJQ9IEUDfDHzM/VmYja+F6FienQtNv1SytXDBxiQ
eY4yES5hjI+1enSxXaL2D8nQ4d9alkPgKvaiCnJls6ABF7Pfcc0a29JXWK2aaWrv
gUgiV4FtotCqpDfBk4pg7RQHgQ9G9YDYJCgJVbnNqIzKdifLXr+ikwPsc++Qiwbg
jfUvbNqrimkLy5mOF4vmGYoTOwsk2v0RNYjHFqATMwmSOdEQ0/EGJHrpu+mNNfy4
zQIVaBQDVOfYDf8qCpvkv8I2Pg953m7gVEerV7RDnjeSvrpZP3ulfV97aEIPHsS6
LZVNiLYm0myt08BumlujeZ6YQ8AL3FNFd8ucRvDFnbLm3bMqevgP7+zl8t/NsUAD
ntwWdtT23rku7dGxT/L+cNt4kvjMtICToVfTC0QS9ujj1NRaVsaf3yRfeKTZOMVS
OGdP7787Kj/qZeuC42d89137yHHbQDzEkqakYpUDbd0ThtNuztNKpwjTtaIzTGbn
aTqwTeiuQDgGjZh3iO+3dPKfj8VP85n80fpfFmCAJXOsQxttouapLhcpwOQPtBIk
9l0FOMTIi7pC99bJAhs1sbn4X7dBADKvl6OJFBmgPq9Crg91InsqXrMbb1c4udCc
8nadt1k7olCs0jCSTtPTPHqnBTpxVh4ZqV3dDpqqsQ1l1pjw720qsfWZncWNBdY8
fPG6a2S8cuo3sCd7J6E2xGRr+Adr5BrIUfI1ndqR85tGx7LtAAaLBYnv6itjH7VD
LPoW/oAd7Zz+VR5877kvjNoHM7mGrajpCbNoSylDzS3UrcVwHJqSwF9aWoJ4mmZV
YJajt3RcflCcps9pJIlYwm7aQ9ta1Jkwm/+GRAT/7Sbk3Zih8RYgSni6qVfsHBpR
yP9vhbomvVr/AGlGc/xr4KcislkDg9Z8rjpQkbZFm7hjq33PFOEHc851USYrV+me
668J4C/nOJYau8tQA9GawF4ns3Wn4AKIq90Plvw5X99rrsS0CFVXWOdo8ZcyJL5q
zHgbIPX93nmXyUs9MX8YEu0R9roLn6ju3fxzAFbY+BGioEaEiZNWoy/ATz7LK0mk
6UC784+Gduem8NcxYX9Hpj1NA18rhejfZ04nWewa6opvC0zRxrZxImyBa3sH19/D
XEWQKfzYeB5DZb2lgN1LNu5u8lItL6gN1hn4S/40KUrIItW6kITxYS8oUUFk6VyP
9mKc+ytKzA8lqtVqah9ZHCmxfFh8i8ibCsRnUkndBCF3q+VCF2G4/ma6ESqHz67Z
2/Qgu40bPnUwYKuylHi7TRheCVbGD6DXxjR0ierAUJDAV0FPTrTRRGfwZ0ryJyjZ
Mzr/5NrgvbJHYF/CCbeiA5tw81gZEzpDi5OzAfpV7OuR884seSzGbvuKbk0Vto35
G7jaB7MMEpu9OAELx9qVX5Tz/qIjs+YcHCJPnMZAZa0T2M9nJ4ClQYk4rVb6rg06
g8/1NlM2q/EPLpSBHlU7nQAZbbUr5S2dUNpYmJF1MwEJcd3g7zE39EvdZulXWSz5
eQrAnL2mUKKIVO44p7P/SOH8HpCoZvEjfW0UKkM8oKKz9RMa28vwdB/r7b4aEPHv
STYWHo4Sb1AH19wxTryfZR1hpkfD27FEA4gCCR/b4+h4t2+jbV8LpKXGtsmkDj/k
xKWZoJSI5qW3MXwWMcVuidOctVlIy/tEWY+ogU4ThHuNStwS2uSFUItbORjDqK2X
NoTSOC4FdGHPmXS/rxgqlHtm2Luk1aM6A2pYPs3xETNEUPRns9PQBn/gmNOn0mLg
/yEsRfT0Fcx48iGKaVRFJgHEfLYisRzqb+0Khay5BoceyId144+ahwnDKl1oxlvF
9S3WmkzZ5xNO05tyhG7P5jn/Qyt9/5X8Ekbmzn4wgzrck3NY8C48Rm0k0PbGxgj7
al92lUXBUuS8G/d0B8Xyht91IeqXcNCb7OLNYf+IGGCplPv7Cx8XNELJYmHfM/EM
3GMObLryxavDxt8UgVNlhmJH2aopVsZAxXfgC6nVc7/4lyu/3x7h27sf1tzsP9+v
b3fY3azTRFWtziZtDh5Ep08kpYOB88v5SOxcl1kWz+XdEqv0UI4KmM1nx3REErt8
vY8nmuizXBwPeFHhw38bGb8sOm24QSK9+5AUPwUKGET84uWRPcvZmzZTmKTl++rE
LpeJryt0OTPzJQTHTNBKrIMEZHcuDkzevn9wMaYWDljFnJLnv6yQeXKmOECmzLDD
TsurqA/MlYAYtCSEDHhfTfNOT4ZwvEvXokNNzMNUF0/txMEo8ZEBU/6DF7jQ4JXh
9I2B6QwNrycVjGgbfIZR6ADCU6Nm1RzzxkfiTAhuA9336lkGdSK8QUp9RqMm2Wfk
BULtihHmlgdgeJ4g5ruScw8jY3s3t9/9vCwtxEbb9d5NN6+gV7ZL0wUtX6FQd5ix
Y+3kGEv92qmmkyYym5/BvKCYGUQrwdPX+AHxODdlDfP7MBzZM7T1eyooB2KTCnM7
Wca3aJKKgc75S10fJ+UKZDvXt0aP1ecNomFiSp6OCTbiG87WpnxTMZYFXbgRl2hm
t1A4ZCxKeQ5qozJ69WkGFGzR+ZdG66Z8gX6s4xxUXho+juwDiUK4xlsTv1fYILXW
WCKujGVqlJDXnhVi4MlzH5jh0kwGf3gX22JEYp/8ZP/Rot6XzyvtDmuOY6Lh/f2A
gauzhUUwiAks85iKWVlTIuNpyvfFY0vukUTnkyyCHBS4Lb3XnH5hY1sVTB7ak+uy
UqRo/af3rb5+HNrGXsyigw2VsVD0DbsKnYPvTaYriBGIEv2rHyBh/2uY9ErQfoc7
Zb+k/LCzk4SlJ+kPfpvctjS9a3pPCrlV/Ww36ojnPxdRHFJfx2hoStKoIAK+XUSn
Jiq4tCaJ6DEKIMNgdkc+z3oBp3d4q1hFTSVd0gxT94JRm7MEI5cebk4xLgx9mLE2
KKmuamDcwA10BpBQNFME+Tx4TyYqMLN69EEZ1YDdrI2799e5ntneDVmjX5b4ySk+
DJRVQY/MSz4cy0f0Sr9nzgxSlSktGi46QopOXbA+NsTxZjB4Lq+JcMIHHT00xkni
vGG9Q7BFlpApNavmPHFxAPQPkpSXkQHLy01GTXqlpAknjk+P7kxF4YImV4PT3T4g
ew4Tqs0cyO9HQoC9hE6v8M7zU78F514e7XcYrwVODW3hSlaD/D8X8eIG5Uh/vHEh
6iGyaHbqpcgNMCYP+tiP7ftTdueVOQDtCfZhmIL3YMn2OqeBDizWDBs3sJGlIgj1
ACBeTsBgElzEXYWXYmoNdUgpo2RwJBU26aYqyByWfV/bZIdn9sKoZg9K9u02wMvK
cyriS53UT26LKkRNQCyL0haols0iFFa1hgz+jDHZlmSTkS4/73NzDyrzUAs87sfW
/T4qwpK9P+P3JOBrVJEVzmSwxKT2jpRlXRtvAd2aukSVu0xOO50cc+aE/yElcCTT
By9X7CRrDxJ3uZHe6D0bdNYf/v/7PJOI8uj4ygIRGiGoNwPI5EJQG4p/Mc5GVG3q
Q1u/Z6OVX17FuceeinEQ5uWrRrqgDQ9d/2KGyzqL1KhuGbztEVyk6Asz52radOtQ
aLnsM/a/C0a8LaEo46KGgvU/E54dWYgAi9kIyIg1XQymmLLzVdyeuFvVbb714gxa
c0tSGRePrJMGzLx1df9P+YC35zgXbBPwAHU1wo7gI1yaOfTl+qXpLqYZAQ11EVTD
jrCoj848FIgLU1oDe0GuNWMh6EgtJeKecs7PPpUlttA9n5WqpW85t1TSTrxyB3ks
nFsKMIl3/by7GDmN8UAaNLI8FuYqTnhvBTBDNo5P2AN5oTyaq5MDJJBSQEEIhX8f
2UWknbSpg0LK5PyXRVBnnX5HhlnB1bZc/qweDNY5fFqYrieyCVKqZm6bThi07OfT
ZrjM0KRXPanZQ+fSGPL1zG9HJo6cDdijo9SyiYAvfm9To615RMLxGZLn5EQJz9vL
1u9rFncccPaRR9tNnqQJLzA7mcLg/0AJ7Fsh6HndLZ4O0NtYu8pHZaCYo64IOsNr
b6/3e220iJK4TnFux9H0LjVlYcyfhd5aUE8j/98NaO3GtXI2qnd2sVjCZisFcH8h
+bx46NvbB8xfsgEyxk8yUse379T8jdBAckFOC0ggYeelTjhfZZGET0SiuJaDgXHQ
oDXG8VWxLQnnshfBmKWr5wQaB2djtOwleL5c4LQ/fyt/dNajZK2hyHb1+IAXAjAk
n4HFFsvrBkfuvY9lb5/gsQwha1H5L5Mr4H/yoCv8gVCSmH3in8cb6ndix4XpffjB
a/R8hox+M4/4LXc0QRdQ3tS+eNflhsDi+z/E5mkY+HS+7pw/XzfA2sZfF6iG/dEC
7xmvfZ7969vHt0h7HPf6kefkWcTNUYEMWeNRFIU4hJmxj70fAJensvTxCkIBvJDy
rIh1dOGmV9W9WlvsYdD+5wpjFBef8Z5A7Pj5ToXYQpmyihuyeYwMftk24z2PM/MQ
H+BM9Se2hbC24U7Uu476ycA4DXxAiZE+gwxePAkjN7nmqiNR1j5GWxIoyLt6TBWk
LVyIVAsJZMSNGhlwDniRG1L9RmQTRYJW9bj7bx6CK4P+s/iPVhSfIKXi/OlzUcTN
sBkdUXTGddE2XajLLHAY96b2k7cGyCFXMO6f+ZJ41D73u2FvS3epx87evVU6e7la
hpu9UIVPc6AiC/ffHyNHgxSSLr8ZDnSJ3r7G5/mnNr5tVx+aRE1FRMnl4z0te1Vh
4kG0ERIOLBpzcenueHVJ63lPPGJmAj20JzRNZNLJIHANzUhJwzc4q1xMk66Q9lfN
y4PgrX/KfApGMES7/EP9p2VqJ+Q3g6mVKOOB+FwB2a6qPXFlLAwXEHrLdbgdbIVL
Stt9Om+IuQdFt6DbqumXEy9nfz3qrNayL5KdiLE7qWITr472PbPUIt3z7OBYZMMS
aEu2gFEF6brUTS8501ByCOVYAwdM3gkdyCw2T2Tb5HpVgdZaiI8DF7qNd0EhrqEF
cUa50KoEWDUF7kzCpo8hhpCHR8jZSDuiemSDVj7sN7nZqiUM7hfLsHBh0RCnpyA0
LHX4aNsy5inZdbOXjK0R/BvLVs3Ls4YWrmgWRzBkBu4tu8d4Dtr9ltFvZyds1uAA
etZk9OxWXYOsAWQ9v6wqLwVQrTQItlQ1TkOzQJQApeqTkmBysMTwQ1Pp0KKqEumG
UMUvRPuVlY0hDNhQc/o5syBUd5UZZ1+gxFeaez6KgQqst/g4XFeVddBBao/u3JBv
gpuJcudZIUlR+zW30nbzP3PFF66yhxowmSunQ+/mrj9nSupINVK6nGQu2+Q4iUiX
2vv7gkMwY4H2u9kyePEu0lMFM1jSVBs46BP0y6mluH9EqMTE0lT4d1w7bSw3wjh0
Xnhu3N8nqJ0PSFai1to9TTF9FQJdjpWJgeLXkfGsZ9g66DneLVp0lOQKH5i6eQL4
blnH7t0mna2YbYteXJnwniq8xTgJTHhR+US5u349owU14riDVz2IUqdeizdMtaqM
4RAU4bbJewfw1QEq9N2Ma6HlC3GIFZ//PeUY/w/ucBp9o6bseN4PNt2XkyfZiOJS
9uaCkaKR3ZtP2bxs6k8noo7T+gpwW6ap5flfv087dqR3EzEtllpQLzn/GxBjPXhw
rov17gYZ9Dne74mVG9FPBERwOA4Or6MVrOpsL1pFnme8Tw6CoH6Meu57kAmBwdSo
pMbpJA97Bm7RtRT2CoBshUOcdOXnnpBx6EAoCAXDHvkP1jLi95kc1h2c40eYIHrE
wRkP/QUQ/TkPKi742NgxpyGd6Zh6CEadC2p741cySXBpoZDNdk0KHPxMz08NSr76
Rz4+SsIaFcCi9zRvOShLS447GeS/FF7H27SlbcxNPBKc37Mkz33iK3qLWxsTXNew
ykl9Q6EG3HzN8Xr2dMCJvy1GAuvWTJzstUSwGFy46xKUf0BJ3003w2rGG9aOwfZn
C//SK2G0dutlfaY8BZJZxCucsQkUu0VXbAvpsJMZsOvwjpr+b77NKTVAC5lqVf7f
vP6s3DXGS/V4xEUIIem7RWUKH9gaNAHCwnW8Vd0VX/fMNrkjs+uhzQEqk913dHzT
vJaasuXU0ElWcq3zIh/qOThpR5bY9ZlV6DqrVwm6Jdb0MDKdbq+DnBaM5jRas6tr
sNQd5rsaiV10x8dQ6faRB+wmwHtRsvNnODzM6RRyB0HhHGChfM66cT1PAoxgFHqo
UxqXXkPw5ZKfgg+0DwxEXFxyaZvoF1ESpfC7Bz4EC2S/tolPuchuz0u7+iOfiPyq
1p7WuXmKZjYAwFO4ADFgFHwH4OQptLW2+27ANlN7vlPGjStIJ+7zTuwrkDFRUn79
kY2yDsC5SzgmR6u/1X3XOXbu0HVT4x5yGy4I0DM7EmS3Ret4zanysOlRptyjml21
hfM3NNejGnLmCOOos6wZf22Y0SHElpFWKNKL0guvhLQPuLeW92jGhx2pKS01rp9k
m/7FhzDyEsntnNjrpSRlkcllGG32S0J3+WEmiEkLI6A=
`protect END_PROTECTED
