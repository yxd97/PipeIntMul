`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LNDM33WwtC6S1jBD49X5vz/lF7R39p06BVPPnf7wTbz0A+sd8WyZ3E52/8xuiDoC
Fyd26rkjPMYA3CsiWZQjr2IVZMg6S0O+P85QmC0api79iYLSaW46IDqaNYlqW6j1
f4bH0VHGLoO0n6oFyr1jB3++9sSmTSESZEIsnzPXDDeYrrdlJcfx51oHOCvmsjJM
VVg51grwApeBGZ6w0NT7X3VhYGhnQwHBAl/SQ/G0P82ySqR2jLuP2zGv1ealDtoE
/h26xvv+W3c6dQtLgvCCvfdKI8HKTbzKdvq1qroO6hd/NQR4Al0O6lXMeZSP+/Dc
3nZ4hdypN/A2q4+aYOvBtQ/IftVz/xJWluHczF2A7gticGqvEwecKXVjKGWg+hQj
OyEeGfedB9VRGnJB1cZqdnQPjzibBrsbUu0ph28eOjpMx36NHhofEN3T/8xa/mTy
uSSLRFmJBwkjkkowO+gD6i2ocWMFFzz55pqaCtsCidDVc6i1vqlIioLk/pbQO6US
V5Ig+hAqn7Ppon5jLP+4hWVTcm4cML7mB1ZDvA3MGm5Val/lMf0uxMatCHVQOkSJ
wEu96IDlOoe8JbrYuJUPkKehsPJar3UCN4gVpFaKgmWDLzjlzDW5vmmDe1CusfIy
BhXOnal28ZawXf297A6nyatNQx6lw2ObOkxhGkgzyD/30UkBu+k5sau+gYW5rnUk
mQd/sWPtSHvWF2Hd05PGvGfT5jRb3PYIMIaZ6F4aE74g0QoZsPwFEhdkUyDiLhCZ
vlaXGXB32Z8yLRV6e9oHpNWdi3BnTqODABkZvZ33X03dSxoJUIGUQjNdmDa9HV2N
fS1h4p6gsexgRmnO56MciBc9t3OZOQ8ldBjVQ357xPjjhQIeA+0NybuYlaeqTQyh
kguhU8VW7oCvm10MoCv+LDLBnoHKfmxruTgOHYiIbyGmG+qd4wxYOPaEUr+0EWCo
VsFGR2YcS0RDVn9n9epy6lb4+A/9D/O1fyR+DHfQwdRc7wzXwEWt45X0V+xR0w6B
FYHau6ARPekG1EnBFIWYf1z6HyUm8UWiZ5uyPyLIANw215EzGrc+I7AJSmH2ZCGo
OT74RYUmQnBzq0ZPTjPXY77cFJKN6zF4anGeapW58MeqhwVz+ug8uF5yOhoquyaQ
afL4jS2fDfXO4s4t77vN0uvCtdKThZMvEPlMKFBejZXwQjFJ/wsugjrOd405ZHIV
zSTZFTIEtmNI/FQwA9GUgVkNBfh8gcibz0Bw81iVzA4YKiKHPXmbEo7z4KM1bfzH
xIHSlkj3/3SS5jFL8ZT5nbROXMdfzjHnDk68kjwhv29ehmjaJ++OyaaeyRHztj90
i13DnyRpny7xN9jDptg7rJz0dDesYX0El0raLu1sj9O1fmHHPzfQIbfGgWBoVdoV
ZluPQ+YeeCv5fSuLVrcjC6FSKWqOHbVvkq9Gc+YyxfFV1u+KCQAZBezLQ5j94bnF
JIR+47lPeZXrsQNfl//sNPzcEebFqGqPyYSW6EX/HFZLL0xQUdXgMF9pMXzJwaMc
PDfzYMdWCq+04y62STe+RbTfRTaMJnWZX1lrZ6MjbL7c0YpxW+eStLL+NomYXniQ
WUiVAB2QiUDN0Q6Fa0UlJ7JAtK5jrxz0KInxAxlWghgRGAlHEuwDkPxXy5gmCz8O
aWcoSx6OQb/lQJTWkP/4pQULpN6hKvOMs6xvybi6Q9i0c0Qbq1yVpcyEEphmHQfa
XyPc1yAooBJ6FZx/8cy9OBUFEbHtDcCVauzXPquK+IOKQ1z4YtB5gJskf1i96sij
KGmr4LaR0nxuJ5CNUgCK//F+ldRHIpgEGVnim8KCz3I2ZBwTjr53s8m9hoYmr6le
4kY4/e327RxiwVxZwV3qVjMVB8EpRgqv4JzuREjJ/8YtQRl4z2sQ6KS99cGjjZMO
rkv4/UQMvkpARl2haueTneJO0mF+kFIB2cxn8ee5ajx+sYa3l7z6+wf6YQ0Y3sQw
BZHJhdAK43j3fPCTuEaL2apGnM96g4xo9ICGB8cuMrWlG+jblWiLLDjhrSEL+Wcu
HgGnheUSMhtkdMM/IvoxYlvFjfV5HxXG5IU451Vn9d6sLlx8J8zWDAxWJ3F10n2B
vQls40F52mwfTU+bvRMmyiia+wnWDcu0N7/H345t1k3U29820yrCeqf5VCCwmRpk
Fj4DxbXDb0+y5q/gBXf3K+Rix0dzO8Xp/olr5EZbCEw7QGm+UI5N9Re6oOmMQf+9
nmazmXaO0BBHnVGXrubbM/EwKLzLtyFXkPVr1pX2dRqDLQKmzaUzKH896shVV+qr
19pPWdzDQKe9e+Fm3eoJNnHyNTmZoMiiuj3FVOXfyd4txptE5WSdzNixjO6LI97G
B04TKwXEiptXftaxo9LlSIODnEwg7BtT0J6pu3XwtZRsnNKMuH91NsmM/JRu+8/e
lZS3vMhZ2E0sfOdYNSSgqalTvTvcCbldcD2EbWlxI8ownpZl+OqghNoDpWriQMJo
cMatXQdKwvS/q8zbb/FMBNeAEavtLXVpsfxUsSEyHosrsLku6T+kWlgF73qKt+Gn
/KGo7M3T/yMycMYymnM8UATtVQ6PuNmpOSiiSwc07RVAzhBEDFpXMWfMTYwNFd33
btc2gKfusIj0SaJmEAZVro0lbUxb+tDGFT82UTnjHJ661KX9q3R0Vkxf3/8JLLAf
ausUmjEBwH8Qi19pAcfCUGUxJHwe34mm67eNNdd/2Iw=
`protect END_PROTECTED
