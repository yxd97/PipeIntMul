`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
grcgzI6GAksmmJUty0rM7EUywliwHVnDV7709ybKUqCsNGROf40nPXw8ljBD31ey
4o9155TuUEwujwxbCNeIMVKVPmcuHxHvree+CJUtMJTBIsu072Tb91PnF0UrZsfa
MY6xMoNvnhZSKRtm7xakhwaEGztrBnUs06smJ50BMtlSxSZAGEg5rAR9Ub3sUlbw
a+TPsXTPrcCfmiF/KV+xZq9ujRvkpKaxb0xLfgpmfdYwC5zbEYyXfaGfjbUNHy1L
P3N0c9w+I8aNng1HjvqarXdUKqGHcvE8CAuQ3zTxKMqpemg8pZ8SOvrjIy3q86sA
51tIUNEg0NpbVPDY/Rf0MCEmFxpdEhwKlrmn61E0RHT8/kw7VX1IQhbbvi1My+Qe
7A7KWYzioWXpf8p8uxXkCmfpzXdaoLFOHR2W21rhd4qLLhCjFTB1S49vcRK9P/4z
31oxTa1d5ccBFaLXBWhh8VQi4gsFLUda+LUH2CLqQ/1jxfZnaAfBOAUVPnDkj1K0
UlzhXvee+kN2RKLKJAT1tXhzrG+WsoypfFRIE+5wcnegmP2Gt5VF9fw9O2rIWLGY
5W2L/hTXhxFrw/FZb68bGQbowoFU04AqqXJ1Je5Rw5N5I9lJr6t4q2KiFRBDXgbw
eHIhpC0AMiJB8DBnqpJR/uC+OeXdfrNbAIDo37q7wTNgGr6otA5lCojBbAUolu86
tG8KgHqS4W6IgxpGkIE2f7OTXLDw9OolwyK9iQvqJF/Q447m3ioWvCnVMG28dqO3
LBXDZmC0Xb5z9feOHhqMFtGJkO4crYs5chkstsFxLkrAe8kQ6X4Z7ZU01IQDKYr8
iyLZGLiLb1cqTLUwkN05bg==
`protect END_PROTECTED
