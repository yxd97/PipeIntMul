`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ok51fVN16esVdyEWj4EZdQCLXjf0dbtwEJ52LIF32Bwsl1857VRYHh6/3QIFfe1X
KjncLphOVNxy9b4+Onr/LXtv58ioNjtSLFPknC2oN9jflgdCZIp1oH0bFrsm+tT9
y54yn/J9FYEwyILnVhlGjx8DJym9jGOJaz2J/yeVNTl0/3jgOOlwOZaW5gyzQgm/
93SXePR3Q1eqZmArPqFEVhR8OojCRLIfQgMgHPhl2UN+vfIB5edSUrwOgzxxKdy1
OUL4IkaiNNkJ3ZEj+jFgx3/ndp9qG5DN3lN6f4+SCSSXm/1V7cJadEodDaRMLemD
1qR0YXZcBKmaEp6+X4TKVRRDVFZUPk+TKTjLuOffNhP1MUxTqpKVTCcAYdIxA7A4
4nnVmbaH2mcT2wMNDW7w4ESRfVdcauUo04i2vWgaDgc=
`protect END_PROTECTED
