`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5AJBI6LSfABTa0v/FeqwRNJ9vDyiVzuhZ1eWFSPoDaulZyhWq2oruSbwFgWn5/h/
qTmpTNeNRaJHp/gZ18P02V251bumxjhURuEpQKsGXMuK3OUSiyA2JvmO6rpF6Lxt
Z9TAk0ui6oDbJt92bGpJapSGYmtCpGjFOF3YlE5R+EyjNyETUiUyrnIA00oLFiA8
Mjwloh/F2lMdRBIid78LxjSgCAIHmONsHhWAwFMlvdBgMII46oFmMeIZJhp2eUtF
RMSCcsJ9OXiPc/KjUYPQuDWIM1uZP0Ufpz9E6j4s5zugRjYCfzp+DoJcjZwNMD4j
UeEW5Nq6JOcAyPFNC2GlaOf227q5YqRGisFcibHt0AhlLBGeYhNQQ2enWdIxR46Z
yFOdR0Z6B97t3+bh9kSbLY+AMe5wJLeCyooEqDW5C3vP79yDPJ6g8/HARHzO2ER4
mnBby1rGy+DBnphbqab7iIfPdq7sqGEgRVFob33xGII=
`protect END_PROTECTED
