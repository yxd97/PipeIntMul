`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNZb89XmXnUeaOAh+AbFSQU0Tdsw40lHtdI79iaakFli7SB2JUB+v+p6f99dUao+
AM++98rBIGKL2dWhFu0moxih0PCYcy3rM7xPjuBjTtLCiJ1i0Svn6wDsudPjmOAs
sJv1Yo2uNazVaXKTxKrtyETGY/ebiN+VaBmAWc6bBmv8kfpTHLD+ug1XOc9/ikEW
Rb3F6p6wG/QK/qF23JkSRePWu0fEAjs44ViMT4Ko9VmmX3j7lSKsnpIz87r6ZJMu
c8ZRuWSEW97HHYMg0KIrnDk778boUaYOOR6ab3ZQXU/7jI1oqsdbHP3WbceWp4Xt
m/Gd0iiQNJqELUVurTK/Oe79/hAtcZcDpiI/l3yCUxoeRRENp4c8wfldl0oe2sTl
`protect END_PROTECTED
