`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXhcUTuxmqZnHG/wEbvtuF6z7Gzm68rs3LOA1sio2PFJbVhGYWkLfzlo/qzW7W/I
NJebjbb4Knj8DidSHU9ZYsT1bMHlABUYcEMy1QzLikeT1Qv/EEM8ME/Zy/iznwJd
i2ZigdW6bMynu+7ptFsRrGnbnMQkIQ7NGzja8L5WB5gB3H/ujyozuFDmmUGxhKnF
FShA5Dn7xB0/8BKjZqbVOBDgNJtUCjF71/K6/HGakLjeefNpnJHX2qQ+g96e2YOb
alt00EpwS3tdZI80+MRv9S/pAIb+Gn81urOy1XZ/WVPEYIErF+VXnu19HC+1yDGf
rpqs1qTaxMuRSHatF6krgzKK1pUIYayd9jamOpmIQ/MGluLp0txHPbGpRrHpTbEy
6ENYOqeIjDJ17f0lPU/0WX+upwghISYWqE2198JgfnPFx6Fjn9HZ51gXDk//0jxO
EL3G/2zR+rMzMlrJeu3Yc5JFPPDVBMLw5t/yp2SMY58kmxGaqDTbpa5uqQ+5sBq7
o/DlafERbtrLAEPa57OiiyKoOpooJ/0iKBRRkufRJ8WLwLKrhMay3kRBjH2vuD1y
sNghr+pOyib0mBtgrwCRQpdulBmeb5DHfNZJ8J33Wn/q8EBTIK54qBMRdOvlI72a
w930ddpZT4o4YD7cqfncvwQfWmJwV6MCwv1g0hq4edW6FMrzOOdvkqCpWHPl38J5
lwnUtbLQUVC4rT3niLbTCQ==
`protect END_PROTECTED
