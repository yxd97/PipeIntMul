`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZ9ttUCnjp+qys3oCv5BR+KeWSskKBIQ9NEPSm5vmLzf8iVexuvi0TZGWEfTy8Ku
sS+tbNP8jxtEro/2Ab4fLzd0xYfe42H9FC/Fl3juCxdHB7GDHVkaSud88mRhosUf
c0yHWQlqSGyJwPXOopOXTzcIipV50veL5tiLBEllgFc6fyl181afq6uzlT7PHDWT
bMPFk8WDXVG/9VNLv1bVZjIL9UUX19iXr2sWoCaWNdhJAkIdHJ/w4vifWnTAE5dh
CETSf5NRKDFfJhtBzqIWBAKBq/MIV57Q4RVI6T/4jFdKQoscPQwY5PRI4FfKOAF3
VA5962R0tEVcQm485Hhxh2vcMEeUlwJhrVBxTMnAnMCy5iBBwmxpINd9Hu9I3rz+
2diiDigjtHGqEkz5981GYhvA4m+OOVMt9vOWzz6p/rk7cdT0nqyMmEDk2s065KHS
6IhO2Y4APJqsH8yFi/g9yoZdME45m2R/VNh+Hyg4v60sZnpEYgPUzbrKriNmbsCX
nj0DnEs8jZBcxi2RiTbDIVgiGSbgoTU/sgaHBUFfDJxJTiqTpT6ZFwoSWs3wy1wX
mytjMxReDhNAtyU9z/3NVLdfeRXDCdmXPKgccloTbF2+RdO2eH9Pp5KFulwqnJtE
KrtjcMJ6RTdUwEgVhNObdAsz7aP10LncqWYf+ajD+3idKZ0BjuBDi7nDcB2aaYdY
vTEidoz+1YnlLI1IWgiUArbs/NXlqKfvJjzmhzpZhnlhzZtYDU92zrkYw2B5aqQr
cQWn6IsTdexAuFxFsm5qJj0tDkv8cYvDIf5FlyOGPKIFfq0HSE3P3w+8CkL/TxnF
`protect END_PROTECTED
