`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMckEMx0bUxPRgSzSRBRJTYQe8pII3pRA6YIeME0FIsfZuV4a4JJZ3gmwTJ8kECn
/+f0IAhUW0IQY7dnlsO4kmWQcqb0M4QFIqZFQxFL66zQo0TzQQJyqQzh8gzCqEmd
M4Wt7RID6Lj82kyfqQdORUJKZ+T0J8D9SHWNfLHZneUL/wNTZrMFxwcjiEvppZvr
GADT5OueZbubgKnAegs8ekpy6t6p9ZzTRfVbhWqUfnqizQTIoTMvEQhD+AmBiOos
KzJgW8HJpeWEq0a2yA7RhbnmbwGkKrw/Zf/vIYw69+vncli3lF29Scr5WHnJ2Cw5
3sAuu3sJ+BQHhVfK/EaFHRjgKSHnFFcd4iujv8mbtwwCwlUNj5ReWAmbr/uwmtD9
lBZx8W2aR5dTN4Tm9nMz5m5L/r//Qnx2k/0HdPiAhK+tLtrFXPLHEaPN9wyeekj6
8goPwT61pEi4INWHjyCD4OMhY9yU/yWpryYsI4/4mzzHElLFGNNSns5owRy5aoIW
UHnjGWAn2CfjeTlw6AOexuE6tPWI7xv0X77Tdr9qZM8IZB+J3VzeZSNOLcfxxdXP
uTQxzveM7u3BqJVoZ01yOUvuVlbDWXn+cig+hPfv3jnTxCLZEmScyfp8yCz7xLo+
V6cdEUFhrkSGP2hjtOVUEOM3wVw89jRoFVUBKrheaZY=
`protect END_PROTECTED
