`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+q1Si1wMh55Zah0203kCOpjKab2XLWLQBt0IIjTVnIR7zdc9AtMVgfoLtm+b3/q
uyhT73zTvaiXdD9A0xPWLTL1I7WCZbmpPCDvc2TzTLrXvjdnW7LofL/CDb5K7ZFI
+rz9fBGz3haXxLoeZ7MmRr0q81UQUrsO++OCrJDXkVQcb/s63u2x9AknJXFI2H1f
WOyx7W8K2xFyzCarxIVoohjMs+EummPSUUpvN6GJv1Mgv4a447UQfR/8M3R1MVeV
YQrWVP0JcDC5qrBTHLiYTLeAUVXpTHrXsJoyUrbyc9k83hTibMn2VMYQxZpm8/O/
Umra+6vXrxqpvEyBcq1sEAoqV4NGc63nyDOzSNNVMIpevSgN2Ja2CHaj3P+2YdAp
170LFo6P1LIJ2cRB+6b/XhNi9pWEkyjEIlnycRt8lRydr4U3ser0GpuwX+HJCOZd
KLo9OqoK4GvG08igJUtOwrsMOvpPofufKYZBaxfZDB4x8CrooGKj2cQ/LijedGLF
+I8E/KobD7UrFbT7NcQTN7naJ9wMZNuUHLB9pWiF5EsOv1N7XdJ8Wax4debUlByM
tG70OAAa+foqGPQYOdeT/Al1oFrYXNDXVwW4e4w0X+eKIsGh6k1slinXWvegtb98
YAKXQcYOT2Dcy6Mpol6AnGgNYfV3EtZ5hwMlFLRXnPkRClEOnU4IDgOlLpBS+mlw
eSqnObHjFU0zD7iYNXTA+WXolamFuZMQe5gaFGCi747MzGdIFWCKHIcDf0SM3VJh
Th4mo2wwSnKpKQ3/jdFj31RVRoZ/Cw4f/eTHNzjzHlstUBtfA25vApGSOcxVX+3O
NJRoGAwAfhp49EN7jEb49Sm/kv2lRnxCv1c6rnHdsEQc6uikv5wsH7dTGBlqXEb4
z0e0OCV2dqQFLRjzS3nJGCUojiJwcn1sdmlPs+YMmJdpyBOj6Hd141zkRK3jq3PK
xlg31WZM6zYBGpTxMsZ718qaCc3HaO9akB0hswhGw3AQ4c/lEq7ouNoRuHriQTvP
6wA6zpoR4/ViHKeYG79Jdju/p8U7D762U+yr+VxZx0AVRCJyuDIuCqoAyTU2oenO
/1MzLdOmvmTQkYRpJtkKPk2nmrExdBBtUECFXRPwvjNLbpAYAOyvPqyycwe7ryoi
NmDaXMRsb1rJbfrXH1eYIXunQV9xBZ3XVay2+VHxap4xVgKyGXZneGblOydEMVxI
6lxBFpsNhx4J+AuxpQtaP9b1i12IATDxWwiX2KSUduA=
`protect END_PROTECTED
