`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9U8L0Vx7trGWyLUtGIZhCb/CYpdqfSfSGMJRUb1OwOnNIsRPALvhexW2FXF+zt03
px6Ba3yo9jqMDX6c63w9/U+y7qvv5b1b3KFb1Q1C5YGyFFbmwU9lxft2pRrV/8vr
+IZo2dMMvfnpBrbo3Z+BBy2BL2x57AQ5Sv/tJzi3ZbZmVdHbr7w9YL9CVHnzNuPm
/m9DPnDCx53AtLz2wA1a3ACekO826hjITx30Sm08eEtE4+RaF26Bdiqm0EGHhcXB
WmVnOkM6cVKBET5hlW+Zn5+VsvRxLSXkESvAj8dvaem9xWxte5ytsVmQJLLCN92p
gYbOBkUGpkTf/5EII1odijzRhflVbJiJUGX4z35nMMt7m4HlinQimJmwK0k1CYo2
xbEg/bDjwFDVASoblW0oBA+O8TNV+TIohULPsAfIeWeELU6QVTS2cG8UQt3VJT5s
U1De7BfWT7yHupQSTze0a7ZeHJeyGVPdxCiFplxIZn4J0bf4VW+gtMkvBIeJqYd8
MZSj66v8DqPNaLcN4BDoZKiPa+MUNtZKJIdHZOdfLHuBf+a/RznN3qPaHCmlkpsG
Y4XPZ5EN8wALRFlYBfkDkXSUrhMlDPszrZIIfOqwyMjtVDQUqLvNFviyJ3oQZDXk
mXbyuzOSbFzhMiL4qBVbtf+g1Zekq6XXMsCpGean29G5Qp+LGIrjKEDP3H/x+d2b
frFQCJSgpIWsuXHH2E2AWZgCO08sV1jJHc1N5VGsG/a1Kg/cbHMgsdvA7CW4ZC3E
8NSXx/MMlEF+HsdY1/UjskuuESQJJnRTsLpqXphlT0oMrYZNsmK8U5VPor8gOWqQ
78HCDlPGCON2QdERJx97xdDNqxcNj7aOzlqvvCLWPeRc/U05Al/C1IPZ1/cGOH+7
vHN19rRIa4L495rWZzLpTYZ2rpcLC1sA5o761/lCePe3GHGSNnaHxlFZ5+JBlqpx
jRxpQ1Y4mzSt8zZnKbWXU007voTSmvi7OM1HRo/RMC/jbgoTP+Ui3rcWxFeSshaL
ugcaWPa9eh/c/uGHqFm2ToJKveONAJfy3arZB1lkfRr/uKzaajDRyiezpwGYIbpE
TTJLfclH8MNpZSdVYwhm3BVal0qRLbYrbcJ1Ba/qy70utbSweCWHPwKUaQ2+URUQ
XPCqDqn2sE72EFjXeAMY3fdVdx4qt0M6kdjFcCJGaNOhkGkpAQU/ibB6k4R3gHF2
lPJCxnf8c88hOFhDUPoFYttSWWjUq8JlKmPhVFmHYsWp1Gemf++rwIjZOXaEmN45
mhGrNYo0E7ikrdHKLp8oHhOOE0mPUvz7AH/mhH7F/iMYJJBczWoOnGoUtyKV0ZJz
ZjbfsPRYfbHuRFl5EwSGcHfXxpgthMJxOcZL02xM++YHGV0kvllvxWm9CDN7wdaO
Q9gTFf5VAhbZ5QpaytW0hqjhkQMgk3B/l1Rgcnou/NoFMXce88gRD581xKslPyC5
o1u5zyB8cGzo/zxscNrMZEo2twV2wJwz/kbilAT6aeQ1GYQh+zwdj2QAQXjC/kpf
7lWYhmzD6UpLh2P26dmaZvMRtK2b4t4V+g8vdjtNyCUxQQQUaypwERppcr7xlol1
rJs2SqgZUhv9JVZn+GBaZUkb9brXN3nHtWWX6nPy34tn+/e/yOo+UYbUQebC92ve
Md2iZS29aebviqLJ2CEWpoVK0wUaAMflzw6tRt8yOx6ppFAOGQmsVEATpk+0o/cQ
RWWgr0MjNqGwR2de6i0boB40ynI5HjkQINtQivYBmWgN0spvNDIg/y/zMVtPuHHS
MfxlrMt0lXSh0UKN7wTydFoFfZcZRvUrms/gDokRX/rAFfCl4MaprdBk9KYge8Jw
uHTTUQEKcxJtFwbIyzackiLcYfSpAitRm4jnmOdh7R9rH2Tlk8Z9E0wKhrwoA1Ue
P3dC8PVXmSAoMlqWXt89UxID+4Ri5/we9sWykminGB2y8FcWAZ+i1PM7Q4HAFJwe
`protect END_PROTECTED
