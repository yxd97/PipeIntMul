`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDTP1/1L+pLJEqNUjEvJ8jfZNFlu3q8zdIn1siD16yLDMz9ur4GkRiz6fxQbnkFt
E41W/lUSK4KQ7r0HzEbYClssSxFq2GgpP1tAOoNZhMEuXKw5aAM+NnjuS6ck4V+t
T5Pw2CG87cxjjojgfhcCr0L+sQK1V1uYMndTW7H4HDuZ/Dl6l5oUNtVhnSycClDz
H/FAKQRKNqaqKcOhWUIheFvk02VGzEUd+scXwzoY39Yg7kfKi6cDOYEQo/CTO8Kf
Hy/v1OqJRETawjra4mg+QfRK5wQFDt8YXtJizrPu37QwftcQ0lYajqpxox3WxHo1
8XFqFVbJ0nHQVbUwR8pm6S1uLTNHyVHxjnPaM1dA8PX2eriPLB5reO5voua0JyB8
+kQN2Vo3sXB+njNZLxtknNngEJDjQIJRlAOPvi7QmnDj8POpt8HWv05i0ULADK5F
1xKMgMTFxRnVAoJaHMQn4T/YQgPm3jfOVNmPvDKKuErQ1T2ZRNCroiU19HX55mxZ
Bm//C6hZevL37YpoSBDvcRUNtcGYJAXfpsEeMvKcpCuLtxduUCLcmUIdx+DSPUQ6
pMgoZRJB89qwNHCubcopa31lPLnEaeVKPBYkJhKukcQHmrURMOB8Z5fLKT4OgELm
iru1EupxHBFfCFj7yR8YKavcysaj2uDoput5BstraMymAhX+2tfSEEmS/jpgK4bQ
6xJrttecOcW4P8Cmi0eXAW0ynnlCFubx/X1jpX6zHmXqGSF7IOtNJ78bf8fnp039
oTwjTqY3jZI0T00+Gy7KPH/bbTbrJj8HXhUGGBI2XGyMu9pRAzyGZaB1PsUbeU9I
yZdcoPAXIxhCGe4+UL/kRNNYdiOuABpo3ECbSTyDZNzwC7epVRszwCESVNdC+aIa
Bag03zVQu5Ca97PxUiEhKDsFKI5epsu6+BaWdm5CvcOPcEwVFi8pR1hWKblVXsKQ
cj2Z0yLI3+OKuuZNYTMiyOEEAkTuUf252ATyMf+yPFuHl6IIV9Xqhjwt2pYV5R2F
pqjXfKWSvEjiqemDFYDjxdylIpJClhwHqJdGtuIHmrRwTB8eUvPQMXJv/KvHr8z0
ZsR0PZgcUe3ZpqV+HkDfsGpMyXo+BgrrUz1Nkz06uNjvq1bQoBqSVYgbrzy17kCs
ysl0NjCRumVwUucbXPV2BovGqWfbflSEkMHj/kOseSyc4tguLeHfxCmMXjn7VSfl
sgZhfz0NdDQB8RhHizC6k4P/8s3nXTyGpmHh4ofv0wNTZYbwUn+ORulBLitRXZ2o
s0TDF/4kQhDBoCB4SxDDfF0p6TFIbCiS8RIEBFYsDP8N1uJ45lxZTsSLH46lRdI/
rafG7/shJAtemUqs7yCF/XdF+hxnzp1AR9CUNiwMvcY0uMyo2UG93Js3tuCtTDxg
jlVjIXtwVmpGBiueG++RwqRuqMtjI6F/FFbbGH6cTBgqzNbN8PcfNrKsQKr7D1KV
O9Ayz3+KZ18qrU0EQS//svisdsE5G39jCTP4aBo04hdqj5nTEZd1wMY8nfzJ10cD
PmgD3SCcVPXO/nNTEqxhXHbxiUlVAy3VibPBdZrGkOfGog4T0jjO9lFUDksFJZPa
l5VVuXGfl/iitcvbDGOnHe2FntcOK6TyTnlwcQr/OgwfGHEcMarjZXUwZMRqa/Er
kUr/BbmQ2e1IuxSBGg+xceeV7W7RZynYuWignKvpLj80kwXsNQ/+K+I3nmDY0I3e
Ze3DXlxf04M2DM5dpA/r340j/44Z8MD2jMyKt99/NvWyXic7lc0Lv4BWGefayT4u
T4nR4wUFMkfFgijs8hA0gXsNPHo16pZXT/a4lgPpxlnn52FL1Xss7nqAc1VfZZC8
JwUoGI73IPKgUMgby2snwqLWo2AGsiaWg0gs3iHuQTp8+C0o3omDWc4c8BcU3aqn
zMePrmi/PzC1TLCjB52U+G5F4M96HbJIGiDdMQsJ4fzPchkoCrbR1pO6sD2pEMWH
oTiMLlo0g1s0Ffg0nW0wxFncgaRJHKv+h+90msPro9Enop5bqPSvWxDZTTmTkp1o
Kt307gK25A4x/lbX47XnITh6jOgXM4ZZeuDKSjH81qgazPmr3ugmccXR99RFViaG
RIrKfoqQZJefnpBtkG5A74TI3kzYenCJRtOtn1b2a6M=
`protect END_PROTECTED
