`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
co0nBHIEuNlaIFxoVC/5TRamTudE4CUHZdSpmU0DvdegTMLVT2bSwY9bEG8/bdwi
qSShubYIEYYsuzXx0Q72uAW20mPLr9SZxkl/VpnyB9ee2wllDmYOChom/rOfw9aJ
R66mKMaZ0oQRSFXC/wwe5bKZ6BxMhOgwYJxT4bZ7ojVTT/lL36exrE3qyCrB4sqC
q/G5RwmwfNou7ADEqsHu3uIHiA21CYUmu9SlAPXwCx5bTcGQfZ0a7KaY60mFZqle
RC4m3yQljJ4WyJxnaxTTWlKqDqIEXAXsUFQ07sYeG06pCVggyhYQKfFZbWKyB9Li
/eD4R7SVQ9iB9r6FCQyYnjUiAwRLpzdoGD/7WuXpiFXsKbZIZSohNIovtaHeyyBD
N0MfG01qBo+oClupTQhAtxDEmMmaHKOfW2x1T+0Vkuiza/vYWuVFiBVouY9CloOM
YKMKsw0av1bKUeKv40tpPzf2fMCrjjhNcqHAoI0ReiVK6Ya0XWGAqQLdGXC0TTXg
mqQztWFeTgxKc0IzrWyaxpohVRGzEMNlknmYoj3rZO+s16rx+OiyyqvurR1k0t3s
CRMdvqgMroVnJ1D8lJYb2EPBDyipsTHHO7wxrHGZ+fLvjibv4nparaDysqT79tGd
pbTJ6P6K11HTP4ydK7mlYoTV23my7I2CNXkeZxSeHjKg5cGml4fiojccrYFU5nSP
Z7q9RIAvVVkgGJzU5iaXsxXCGSL8qskDk2oNRpi+hCek07gFEK9Qlmv8xN2BpFSJ
Ub0hQuvyx9vB/JXZMLuNLL3qT7Gh4A7fPN0D0o5BKgoyRprcbr/dN0MWIkqYLBtU
HwG9uyPWq6MZXScSX0ea12oFZC2NjJsb4l1KoNWqKzUDKY0/18E+EVSdT0nbEe+W
r/h4gwjjQ67TkWaywzcT0OFPxjASzAB7cAgf6pa01DxPF+kajsG56+p1RYEZZgnR
`protect END_PROTECTED
