`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gdHjCEkl5FUGjfe9FANfHjAsmGBmxW5Z82zfn8OiOTC6E21YXyV1rGM8Fjxq4DLi
Mf2Czo44zIsmZHeLbJHR4EpEC260VyTd47LeOAoMOS1gHUA9t+HSLRBmRd6TkHuX
2pFt/Oiwubj2N22rLMcZ4aV4OnO/mqPTIvU48lcgL+eP4hYAk7vLOW5JR9lxN/bl
qAo8SHo/iGfdNQazC2afa2FNW6JFJQSMkMkvjoBHtJmFgDh37rUiDR+hZL3iPvdh
UXKhVUf0Qb0HnT4RMKXEA0NT/J3cWdI+blr3sWSbqDu6bKpQ+ioF5FckeH5+dft0
s/fpJVc7iux+wkgDbJ4h/4rL18BvzVsfv/zdVmD+m3rjZOMdh/a1kcdj/cMVpBud
eF6/Zf9D+sN2Owvz99BHuw==
`protect END_PROTECTED
