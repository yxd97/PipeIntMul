`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cik9aDU5te/zhA1UVvn6S4e20pGPgGlSBhHrjtlSSZjP3yvl6ssYamUcvlvzQaNO
BdxZLxasai8xJAmpGnFRM6djTniW5QTd51sdYhbSbMRRteK1CZU87IM8rC9IM3PQ
S+ahTYM6sD8Yf/ydDztaWZstSzYAUtSlzbpRkUhkjgiAm5LaxwuOXc+fJm2lC1do
tC6LmbLi6eyhow4K8qgXGB6wgGVTTmK8VsiHgMAD4ZfjhWYZ/wxuSz8Hn4SZ+fUI
Se9USj/jXrjIHNS3xg2zivUF3MQmlOTHcEDyij7fV8VKl67D28yW2pUyXD/veKuu
/6H8RgEPmPyaBZQP7jwOdLAbqZRTPI6/fe0079B2sEmmDF8znYBvwEppDSVe08EA
XRnlI9BkBrOO8+AE/LiWkt4A6mnN+jS3Gk8v3PFFVDXq/WB/lnycFJLevhyDkkPw
rFOg/j2FhsH4Ir7cLZKm7iomgFqbQtaQjGfjLTUvVMo=
`protect END_PROTECTED
