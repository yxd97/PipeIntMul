`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmUqvJD+h+gt+6anbNxlH3aSqC3qLwJQunJ1+C8hXOMbTE/ADINUs1R+VUjrqvFY
fdLjWnIhB7/97oSAzvOzLhfFJVj+TpUJ8TOdqFYoAcrM5jk5zKIfwM0luuW6oH3y
029JuFF0KlDJutZEhvWG4koQzecX/jcrrFs5TXj28OYIAUw08kjYlRCxqrQkf1jN
1v4011lhGFv+IK3LFJXCMYYysMog5w8tc2SKXObWdVupMqQUxAcYbVkRS2k1smpl
wm4fmEJPCX6YMtBzNJW7eA==
`protect END_PROTECTED
