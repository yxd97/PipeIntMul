`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yIb78z16fK4GU0tVPLWNcSRyG5UBUlMGFBPr36rnCoW13OQ/sQIQHLNJUnYYmDHg
sBoK8xAVYlect5jwI+5dkpokz+zG8fWUB9DjVZ5fmp3/v1z/lYLkSDCsj5CCprLm
8KaXuCjCwBWXshX8A17gJFUWF7sbPzZ1bEtecvPq4diiwlK04Q1poPLyI/alv4Z+
qbby7a61ZV5ISEHBmVaeb65F5AY/kgsCXE2MhP7ogPvZOtYcRgE68QFV8ww/Viiq
mZN2qSbuDWmpX/y7LUbyoZm+E0FP5tva5YRO7Qcp4BM+dQVzTzPEHygTOfeS8l6p
2/tHyXPlCJVli/CGHjHMgRK/KDLDFCSbeW6ArM3AH4na1149yY3nIZDRKvPLzsCT
moRAliqIG0TYlKHOqJsA/InUGCFnL/0Kr1RYhltMzEE=
`protect END_PROTECTED
