`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8e9ucdgT+72W0li/qC4/pDJUXpCx14XQu8xgd+omRE2BnEPn/ZZgT93yYzuiBvR
eAJX/h+j8Sbnb7U6Iylb50Kx9F846k9nKkHxE5TN7TuuVEcGggKdN42wFaJMQaEI
InVVpfn5kxVzq4NGVjUGl6okaP4lP6Q9P1KgOKwGyhkxuMF38gVfeFgkN0XfTo9J
IOjNM3JJhKYYwA5krHRdBlfwvsSQTLeUbg0bRlj9JJkb6bKhId66i5JjpwrzFesT
jhz2VWRf0iUt6VhXPp7TT1J3Z5vpS6r4oZ1BH2HV9bKUvHQZwFFxxXKXTCGXS8Fz
tdxnp4sIATLt8bmBqNTTvcnDSI0cTXpYc6InPB1pIbo0hWhBwj7q6hSNQxq05pkq
DoIX/hbVqvPhljCRTGqlSLHbjVwXoGfk6w3sYpWH81s=
`protect END_PROTECTED
