library verilog;
use verilog.vl_types.all;
entity PPC405_ADV is
    port(
        APUFCMDECODED   : out    vl_logic;
        APUFCMDECUDI    : out    vl_logic_vector(0 to 2);
        APUFCMDECUDIVALID: out    vl_logic;
        APUFCMENDIAN    : out    vl_logic;
        APUFCMFLUSH     : out    vl_logic;
        APUFCMINSTRUCTION: out    vl_logic_vector(0 to 31);
        APUFCMINSTRVALID: out    vl_logic;
        APUFCMLOADBYTEEN: out    vl_logic_vector(0 to 3);
        APUFCMLOADDATA  : out    vl_logic_vector(0 to 31);
        APUFCMLOADDVALID: out    vl_logic;
        APUFCMOPERANDVALID: out    vl_logic;
        APUFCMRADATA    : out    vl_logic_vector(0 to 31);
        APUFCMRBDATA    : out    vl_logic_vector(0 to 31);
        APUFCMWRITEBACKOK: out    vl_logic;
        APUFCMXERCA     : out    vl_logic;
        C405CPMCORESLEEPREQ: out    vl_logic;
        C405CPMMSRCE    : out    vl_logic;
        C405CPMMSREE    : out    vl_logic;
        C405CPMTIMERIRQ : out    vl_logic;
        C405CPMTIMERRESETREQ: out    vl_logic;
        C405DBGLOADDATAONAPUDBUS: out    vl_logic;
        C405DBGMSRWE    : out    vl_logic;
        C405DBGSTOPACK  : out    vl_logic;
        C405DBGWBCOMPLETE: out    vl_logic;
        C405DBGWBFULL   : out    vl_logic;
        C405DBGWBIAR    : out    vl_logic_vector(0 to 29);
        C405JTGCAPTUREDR: out    vl_logic;
        C405JTGEXTEST   : out    vl_logic;
        C405JTGPGMOUT   : out    vl_logic;
        C405JTGSHIFTDR  : out    vl_logic;
        C405JTGTDO      : out    vl_logic;
        C405JTGTDOEN    : out    vl_logic;
        C405JTGUPDATEDR : out    vl_logic;
        C405PLBDCUABORT : out    vl_logic;
        C405PLBDCUABUS  : out    vl_logic_vector(0 to 31);
        C405PLBDCUBE    : out    vl_logic_vector(0 to 7);
        C405PLBDCUCACHEABLE: out    vl_logic;
        C405PLBDCUGUARDED: out    vl_logic;
        C405PLBDCUPRIORITY: out    vl_logic_vector(0 to 1);
        C405PLBDCUREQUEST: out    vl_logic;
        C405PLBDCURNW   : out    vl_logic;
        C405PLBDCUSIZE2 : out    vl_logic;
        C405PLBDCUU0ATTR: out    vl_logic;
        C405PLBDCUWRDBUS: out    vl_logic_vector(0 to 63);
        C405PLBDCUWRITETHRU: out    vl_logic;
        C405PLBICUABORT : out    vl_logic;
        C405PLBICUABUS  : out    vl_logic_vector(0 to 29);
        C405PLBICUCACHEABLE: out    vl_logic;
        C405PLBICUPRIORITY: out    vl_logic_vector(0 to 1);
        C405PLBICUREQUEST: out    vl_logic;
        C405PLBICUSIZE  : out    vl_logic_vector(2 to 3);
        C405PLBICUU0ATTR: out    vl_logic;
        C405RSTCHIPRESETREQ: out    vl_logic;
        C405RSTCORERESETREQ: out    vl_logic;
        C405RSTSYSRESETREQ: out    vl_logic;
        C405TRCCYCLE    : out    vl_logic;
        C405TRCEVENEXECUTIONSTATUS: out    vl_logic_vector(0 to 1);
        C405TRCODDEXECUTIONSTATUS: out    vl_logic_vector(0 to 1);
        C405TRCTRACESTATUS: out    vl_logic_vector(0 to 3);
        C405TRCTRIGGEREVENTOUT: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE: out    vl_logic_vector(0 to 10);
        C405XXXMACHINECHECK: out    vl_logic;
        DCREMACABUS     : out    vl_logic_vector(8 to 9);
        DCREMACCLK      : out    vl_logic;
        DCREMACDBUS     : out    vl_logic_vector(0 to 31);
        DCREMACENABLER  : out    vl_logic;
        DCREMACREAD     : out    vl_logic;
        DCREMACWRITE    : out    vl_logic;
        DSOCMBRAMABUS   : out    vl_logic_vector(8 to 29);
        DSOCMBRAMBYTEWRITE: out    vl_logic_vector(0 to 3);
        DSOCMBRAMEN     : out    vl_logic;
        DSOCMBRAMWRDBUS : out    vl_logic_vector(0 to 31);
        DSOCMBUSY       : out    vl_logic;
        DSOCMRDADDRVALID: out    vl_logic;
        DSOCMWRADDRVALID: out    vl_logic;
        EXTDCRABUS      : out    vl_logic_vector(0 to 9);
        EXTDCRDBUSOUT   : out    vl_logic_vector(0 to 31);
        EXTDCRREAD      : out    vl_logic;
        EXTDCRWRITE     : out    vl_logic;
        ISOCMBRAMEN     : out    vl_logic;
        ISOCMBRAMEVENWRITEEN: out    vl_logic;
        ISOCMBRAMODDWRITEEN: out    vl_logic;
        ISOCMBRAMRDABUS : out    vl_logic_vector(8 to 28);
        ISOCMBRAMWRABUS : out    vl_logic_vector(8 to 28);
        ISOCMBRAMWRDBUS : out    vl_logic_vector(0 to 31);
        ISOCMDCRBRAMEVENEN: out    vl_logic;
        ISOCMDCRBRAMODDEN: out    vl_logic;
        ISOCMDCRBRAMRDSELECT: out    vl_logic;
        BRAMDSOCMCLK    : in     vl_logic;
        BRAMDSOCMRDDBUS : in     vl_logic_vector(0 to 31);
        BRAMISOCMCLK    : in     vl_logic;
        BRAMISOCMDCRRDDBUS: in     vl_logic_vector(0 to 31);
        BRAMISOCMRDDBUS : in     vl_logic_vector(0 to 63);
        CPMC405CLOCK    : in     vl_logic;
        CPMC405CORECLKINACTIVE: in     vl_logic;
        CPMC405CPUCLKEN : in     vl_logic;
        CPMC405JTAGCLKEN: in     vl_logic;
        CPMC405SYNCBYPASS: in     vl_logic;
        CPMC405TIMERCLKEN: in     vl_logic;
        CPMC405TIMERTICK: in     vl_logic;
        CPMDCRCLK       : in     vl_logic;
        CPMFCMCLK       : in     vl_logic;
        DBGC405DEBUGHALT: in     vl_logic;
        DBGC405EXTBUSHOLDACK: in     vl_logic;
        DBGC405UNCONDDEBUGEVENT: in     vl_logic;
        DSARCVALUE      : in     vl_logic_vector(0 to 7);
        DSCNTLVALUE     : in     vl_logic_vector(0 to 7);
        DSOCMRWCOMPLETE : in     vl_logic;
        EICC405CRITINPUTIRQ: in     vl_logic;
        EICC405EXTINPUTIRQ: in     vl_logic;
        EMACDCRACK      : in     vl_logic;
        EMACDCRDBUS     : in     vl_logic_vector(0 to 31);
        EXTDCRACK       : in     vl_logic;
        EXTDCRDBUSIN    : in     vl_logic_vector(0 to 31);
        FCMAPUCR        : in     vl_logic_vector(0 to 3);
        FCMAPUDCDCREN   : in     vl_logic;
        FCMAPUDCDFORCEALIGN: in     vl_logic;
        FCMAPUDCDFORCEBESTEERING: in     vl_logic;
        FCMAPUDCDFPUOP  : in     vl_logic;
        FCMAPUDCDGPRWRITE: in     vl_logic;
        FCMAPUDCDLDSTBYTE: in     vl_logic;
        FCMAPUDCDLDSTDW : in     vl_logic;
        FCMAPUDCDLDSTHW : in     vl_logic;
        FCMAPUDCDLDSTQW : in     vl_logic;
        FCMAPUDCDLDSTWD : in     vl_logic;
        FCMAPUDCDLOAD   : in     vl_logic;
        FCMAPUDCDPRIVOP : in     vl_logic;
        FCMAPUDCDRAEN   : in     vl_logic;
        FCMAPUDCDRBEN   : in     vl_logic;
        FCMAPUDCDSTORE  : in     vl_logic;
        FCMAPUDCDTRAPBE : in     vl_logic;
        FCMAPUDCDTRAPLE : in     vl_logic;
        FCMAPUDCDUPDATE : in     vl_logic;
        FCMAPUDCDXERCAEN: in     vl_logic;
        FCMAPUDCDXEROVEN: in     vl_logic;
        FCMAPUDECODEBUSY: in     vl_logic;
        FCMAPUDONE      : in     vl_logic;
        FCMAPUEXCEPTION : in     vl_logic;
        FCMAPUEXEBLOCKINGMCO: in     vl_logic;
        FCMAPUEXECRFIELD: in     vl_logic_vector(0 to 2);
        FCMAPUEXENONBLOCKINGMCO: in     vl_logic;
        FCMAPUINSTRACK  : in     vl_logic;
        FCMAPULOADWAIT  : in     vl_logic;
        FCMAPURESULT    : in     vl_logic_vector(0 to 31);
        FCMAPURESULTVALID: in     vl_logic;
        FCMAPUSLEEPNOTREADY: in     vl_logic;
        FCMAPUXERCA     : in     vl_logic;
        FCMAPUXEROV     : in     vl_logic;
        ISARCVALUE      : in     vl_logic_vector(0 to 7);
        ISCNTLVALUE     : in     vl_logic_vector(0 to 7);
        JTGC405BNDSCANTDO: in     vl_logic;
        JTGC405TCK      : in     vl_logic;
        JTGC405TDI      : in     vl_logic;
        JTGC405TMS      : in     vl_logic;
        JTGC405TRSTNEG  : in     vl_logic;
        MCBCPUCLKEN     : in     vl_logic;
        MCBJTAGEN       : in     vl_logic;
        MCBTIMEREN      : in     vl_logic;
        MCPPCRST        : in     vl_logic;
        PLBC405DCUADDRACK: in     vl_logic;
        PLBC405DCUBUSY  : in     vl_logic;
        PLBC405DCUERR   : in     vl_logic;
        PLBC405DCURDDACK: in     vl_logic;
        PLBC405DCURDDBUS: in     vl_logic_vector(0 to 63);
        PLBC405DCURDWDADDR: in     vl_logic_vector(1 to 3);
        PLBC405DCUSSIZE1: in     vl_logic;
        PLBC405DCUWRDACK: in     vl_logic;
        PLBC405ICUADDRACK: in     vl_logic;
        PLBC405ICUBUSY  : in     vl_logic;
        PLBC405ICUERR   : in     vl_logic;
        PLBC405ICURDDACK: in     vl_logic;
        PLBC405ICURDDBUS: in     vl_logic_vector(0 to 63);
        PLBC405ICURDWDADDR: in     vl_logic_vector(1 to 3);
        PLBC405ICUSSIZE1: in     vl_logic;
        PLBCLK          : in     vl_logic;
        RSTC405RESETCHIP: in     vl_logic;
        RSTC405RESETCORE: in     vl_logic;
        RSTC405RESETSYS : in     vl_logic;
        TIEAPUCONTROL   : in     vl_logic_vector(0 to 15);
        TIEAPUUDI1      : in     vl_logic_vector(0 to 23);
        TIEAPUUDI2      : in     vl_logic_vector(0 to 23);
        TIEAPUUDI3      : in     vl_logic_vector(0 to 23);
        TIEAPUUDI4      : in     vl_logic_vector(0 to 23);
        TIEAPUUDI5      : in     vl_logic_vector(0 to 23);
        TIEAPUUDI6      : in     vl_logic_vector(0 to 23);
        TIEAPUUDI7      : in     vl_logic_vector(0 to 23);
        TIEAPUUDI8      : in     vl_logic_vector(0 to 23);
        TIEC405DETERMINISTICMULT: in     vl_logic;
        TIEC405DISOPERANDFWD: in     vl_logic;
        TIEC405MMUEN    : in     vl_logic;
        TIEDCRADDR      : in     vl_logic_vector(0 to 5);
        TIEPVRBIT10     : in     vl_logic;
        TIEPVRBIT11     : in     vl_logic;
        TIEPVRBIT28     : in     vl_logic;
        TIEPVRBIT29     : in     vl_logic;
        TIEPVRBIT30     : in     vl_logic;
        TIEPVRBIT31     : in     vl_logic;
        TIEPVRBIT8      : in     vl_logic;
        TIEPVRBIT9      : in     vl_logic;
        TRCC405TRACEDISABLE: in     vl_logic;
        TRCC405TRIGGEREVENTIN: in     vl_logic
    );
end PPC405_ADV;
