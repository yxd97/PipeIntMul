`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L2o7XvE7EutOdWuWTuqTg02CEbxdgnj1G9865gVSTdpq6jSPBWx4+SUkuZYy3Tg3
qIrf5G4/VrovELXtUvKYzeK8q9fyPsBdtJx1i1uq8Vx5UZEZ/nQlaBAFkUhjx5d4
PLotpneNAhTF2/t1WDWWE6ZonzQ+DzmRJuiz7BkssXqt58zFLrYIY1PuaH/eD1fK
4iynzfcb0DEzrxTg79dqoI9QjQNUxXTnTCx+Xh19o/ZZqw904G4i3H60SnMKUaDd
u+Ez/tQn/FCDkYk6wnpAvt3LmkXhBDosXl2OwbHCmA09GMgAEzlugverW7W5/Fik
PgcmfEmqeODhHJyPI4p5aflvPBspToPjv1exRY4R/ZM10fs/O4PLorjZ8yT8ENJL
Ea3StKvvdpjWY7eF1ARJ4TLJPEsQeOYExy5SZ6+xZvOIJvMmMduG4e6Zv2a+0wX1
HqVgyNjy8wx8LdRhMtYvyt9XJK/EPY70MnLZiCcy5tCISmrOhndczVusK3Ff/gWD
DJRx8sjlaCIRZA2JCIa1Cjtu3uNpHN/wedofa6iWkWRdqmjnfn+zbwIztM/O9GNj
8xHArjWbn7k5qk7RpNSxlFwJRVbR6/sEpKtyE8kGCCc=
`protect END_PROTECTED
