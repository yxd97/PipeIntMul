`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+xL6bEBu0CkJsjzrmrePCNEpUPq+vzpKBKha83vxrBYTjtJNKqTqisW2NkOQkgj
BM4VW99pVEVA7zwup4cHLS3OyNB1XbU79IHtWTQ7IH50XjE8ID9wUSrDQXLngbKt
1XA6OdiWuwnWCj1x1J9g6vDyhJpYoGtvihkI1eFnTmMWIy+tGH4kGc2gFjlZIFkB
H07X4UHdeh5PRsnvUsoocsm890l1SAs33FEFRFn6565etcSe0+lRcf+wx8SMAm6S
h8nE1uowjmKJoIm+fnNkA0RGD2aZ7mbqVN+dWGCfbN1ZhJGKwdVhYXpQJMVqEGDR
2YVKXTmQUGCxHlR5pI+1J+WYDab2LlHQnWcSJm2gQ+EfEwyrB6JQnEmj3msjXj3k
v77eTmKbztIUOd8o9eFRuNcoUAngn8+NboXRwNnN1hh7AIKDVd41VFfPsA4LaeJ/
VsVmovQ3VXtC446RlUH3wpG+KcXOyQc+T6AzVcV7/cz+mH0DURjOhBXQMAEaXraD
Wn2z872EPYpMtHDdq+koyg==
`protect END_PROTECTED
