`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ruxlcVFoDfnsVINyLgr6e3VEbwXcmVmTLs5cH2oodfZJgVkL2TSzBY/+KyWHN17
AqYZPE4K0wmqsZk7hg/EydBmrIalNdoujFUU6EgywU7GXg4V7dRxDI4b77ZizlxL
+dHzp6em/pQyphKsTqARiapJtAMnuU2M3Z7C1AikVNgTvhqA+8vgAu5p3AoVvrvX
cxmDaemn2hgI74PxchaBnHFBGXRKPQmM7GREoyX6FGZMM5vgOlKWbjJx+tcV/X5+
qGLBJQJ7upYkNexG+3X5ltqJULq6E0rJvyR3VTzMtLR/mT64O62fZfKIU8xMAPgo
`protect END_PROTECTED
