`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8aYrV75sj3pubVWAuBO0guCnUGyvOePKkSGKsvtn5qw/j+hIc3Rz0Yshd0xFd/KO
KnJd7jcUM93Iu0i0C/dYtrMysVqWtsisQn0as7fH2t/786coh4l/rUjMJFWKlY81
9k/cW9VwKIsHD4XIpg0g501My3Z8dEh44kyhpUuaW5SKxx61ZhZSSe7Vf+1fKBad
h8S/YZ0kOwDh3nsVYAVHqd7WC+ph0+LGqslQgTg5mDN6jVv7jPJXoxHTg1Tw3ugo
fuYfHHJD3awfMWV6g20tnE7jmUZayBTjO+mAYZdffuz+AoBANW6zfxWpAxx/Pc/2
BVUhPd83rxVmxuljQ8vhmtamzoTRMtOa9BRlI/itFO/YDf43g7DqE/GlUJjPrFXI
vOBqcZRaUISc9uy+Vo7jzg==
`protect END_PROTECTED
