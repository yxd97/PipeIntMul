`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EXR9+w4Hu9O+snJdUUgeiVg8F5sBGa3kHXW+tSezRshngavzW2OlKGitCO6qPWKv
C4uRpZ2w44LP3SxEMonoFwwO4bBnLku+zcQjXkRQM6+S4kYWw2q9hmYDRhJdaowc
ZkMQCbA9iBdCWuXkn9vDqlyTJoods1FmJA8KvbCbqPq14GLWGt7s6DF9oWnQWQG9
PNMrdW8pscy3YxKhZPKt8QlPf84KJj5NSAJ6g/Wo1hHtDqWJE6uzrtlAM8OWVMYC
cqmITkNg1hTZ1gcHBLJffGJjA1Or5hzJj03+z9PA2qdaCKDXNcrLZ4zND1PLgokj
xVkuC0fvjfHjvIaSLyeVL1snrIfiTt7noNoCJjybiMpnMSWkDv9lVsp3XOcLO7oA
`protect END_PROTECTED
