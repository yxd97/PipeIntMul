`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1cJ2tETrrNSLdGFnw4AVXHRwncVe7RsKn1wDPI3CivdXS1dESRirniU8JrLtok/b
v6DnOW3jCMLMY+nxsYfXh/q6T4dK41akS3qRk6HaY813KJIWGUtpEzSmx4YH6ClO
I0noaKptmiNbgu0hz6Y4l8yDJprS6z8lI/Ua7uyjwOaEB5mAnKV4TGTnKVGAL50Y
sTST//S1d1uWxryZIe4AW+mmljSfa0M+FuSbNA1ko3b1Hs/4bSHQDegKbkgHnduO
vQMSjBjfp+mkSrkEdZILzc9fgkX3c97FfdL/EtbL670gYwN9QMmFh6Ch6Wz+1MDn
`protect END_PROTECTED
