`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oc2gaIstmu9jyKG6oXePUG3Rhy/o9xaSt6Z4R/IVLmMMHjjkFvtrQzMKjrSzNjcU
r0z1WWy+YJeoBaUhLl/0Jffc4au1Cal0hkwS7jMhr0doE/CMF8SU/zr9zpjVzYil
ux8YZiV9wWjwQx1yfbbRxqTbWnWUXXnwi1Mjn/tKw1T9foTDd3rfULmyBhVdGady
O6dGo7sozfhlZbEOyUFhhsDNgrQ7DHC54T/jE8CtOEm9ZhRY7LuXjRUX/T+b3KvV
2VghEERyiLOT+x0gozDnwmzuVTAQ6HbKcSzsAOLh7FjiykEE5ifgIRDymX1m7RLf
4mfmWp4ZbaShWvav/Hu3nWZ31h4HoVwM3Q7oMxJ8lopAJYXvw1PDkUSohesB2Nsh
9KRbLeQXgpQlMZYLymhB6pAVRUrLCK23sAkXUA6KuJ9RVTESVzr4qiXJLHQWfqET
EsRDVIxmzz70AM4VsVdMrJgjmQ/vw+opUICFxe7Mn+9wqVTO9Y5XAh9G/TnejaYr
Uoj2Gpgwu/OVMzc9sxp6IS1Jn8gqce+l4KIuISqTZfL4RseYNivfIs1lw3kMXxZW
E63mA+ZavHAh4l31eqG44Q==
`protect END_PROTECTED
