`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MUgecGobaX7cKcSQIWGgKnb89C609jS4yLooCFj071q3Pap6LCaVKAjkFN9ju28
bFB36jMcdFjb++zWSIz3wtKVrPsFyWAcNEXoQ7j9jriA1X/BbU28lO6vBHMrDwCl
iCNOIlRSXRzttiW8eplPatEDdtOp038u+7UfNohGm8bEhWNHw3EBvQ2hCaDWDQ/F
tQdSsnoEgJ6dMgCkRX55ggRslhHMMBZf/WMK1yRutk0zeP5QebcWQQSrpyBxf3Vp
ByvskbvNP0V3HwG7a6uitQ==
`protect END_PROTECTED
