`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0nymZJVqGGpGwYJTgKRmMimfeO/FMSdYVtgZ2La1P82D9lNr7taNqB2ED1RarEu
9wKF1c90ZWqLaM1K0yj4QJIysTqz7ULFV+nI/U0a5Uzikzyf79bFBDPhxbvCJI1n
BV4E52q84qDoQZT/3ogYqJgi/88ZaH0h6eA0dEHW+QxiszGy5JYzteuafThKcof0
aJ7tLgW/Iy8yuqZEdrWzy5oJasRcZTiqd4PjV8ovSbELypY/HyTUau6cDYqfH+mX
kLZgPm+c50NcKWnXV0xkV15VvrpMHzjUSXBl0v5UOeoIy6M0jfgEmJxvyoWsnA5e
owqvePdaenk0JUQw/XlbYGs72vYezGQykTyCNRmQQQvn1DjoknprrKWUKFus8Rft
isX7+WG/TjrMu7KiQQScdceRJce7ZsEGSIZzjrB9cNSpuNu3yInphw9zzOLpRyaX
r9Gyppyf8adOJFtP8t/KWvR+PUWXfVsWsyQGvPg+ysGPh9P9dHIMoGIJar4YVzXQ
01h4vISMXj/Z4saDjVQNXN8+kF+IHOHj6QDG44Yt/1Rc+aNcnVzCu19Z7kZVfl91
cuzAfFI9Kv7Yj2IoSwa8f0d/wAf7DQE8wnOIzrl2MBiClER3nPNKrwDgVELXsoIS
mrd9laiauS5vtZ+hc2710FaE57BhQHFTYJk+hcc1Pvetk532LsyBES4DtRpYA5SJ
5+hAeKg9OQZl5eR2WaRMYQ==
`protect END_PROTECTED
