`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ztx61jVNpGrNvzkLj5Ziqian1H91KcbGi5wDtzkfLULjrIiDZ9o4bV3ke6rTcNuC
Ig6yFE64Xy20LCdY7TBNuFCVP7LtISCNyMYZ3om8s94RDmfRn4GtAtKNSyhjS1jG
v4tTP3Kbu2rLVNEU88OBYahIffUOx1tiXsNCWjn4VrpkAK+Sso1s0gcxZxK3uw86
NSzdHwEfRYnMTYPc6mFiJCCiZYk5+o727fcXJEn7ZfeGer5JoMpkEGlu3+aPm1b6
Txdrk7l5W3/1cO/I+9fj1lyagAnMxTgBN2DvWkaZSpriWOIePNnEhQIUY4aOvRcy
ftFPLlHhZTyvIXhsu3GZGdGFWJKs5W0zRlAqrI184Kh9PNPcTm7Eezh2qTMg0pEx
0p+HYZDS0M0ckof70/tHuvRAFQchWhNJb5rA6GjsMvBE3qInBVzUdlnLQ2SI56St
A26+AyXRHQg7Wmx19VAF1FhfC+0qD7OrAeSajntN40DA+dQ/9PJd7RNU/hSrb+aF
Vl3luESLL2MDVelaAUx69DHZtRlG5IDVDktsQCmLyCljtdXpiDXPpGmUhpUuI5Fl
y+ex0jB5YQrICMwEqiYtnX3hzi9lNfvDnzG1+p9TEltaJFwl104Ds4f1qmYT67pR
OXUjcwmrYvDNoofUOjrOuYBPvavDgRXPAZSecYq7NfJlj/020mIVoOZUb0e7g7pC
NO5EDoi9Nue1Jq+5For0HYFEcc7HONnN0lzVLi6StNa7GB2hgPNG5F+V5vkm0iGp
xfaBWHhMKkzZD19RVTdxVbtOBFXU8GC61QczlUalOn2Vj2+pFUpnsCsNiy8OKM8t
UxISn3TKRuMBYFEEj4MFHmZqAugPMmMVFoxXl7W6jq1oudye6wwC9aKp5vEyGvd/
apyrhb0L9CGd3OOU6mMzxA==
`protect END_PROTECTED
