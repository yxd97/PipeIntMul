`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dz8rIqUvxD1CXcaltsRCVbpl4yng6659GzqywTiiS8hxL8WDOV4VxM1prEbgCbNO
u6CAYXn7Q9r361w4clI7Nth9jYZIw5OwuS+/vgSx7jIsYub1MWbwmNzceFK4uioj
qcNMoJJI4vFB9oMYG9aGutSA5JZg5oiI0Qb8PXKHSiFCx1hpjS9aZaAp+ERiPdgz
6JwGWiEmklvkLT915FT3CuNXImosk3IUNkovRZzmkEb/qEvTR62iODJdF8Fhje90
yLbGCV0z4xt7AITeJGQjeOYPQdvGCJnD4luW3UEzZICmWr2aB61pjdQKOmPo21G9
zSlR2x/thiqzaV3+GCeb6w==
`protect END_PROTECTED
