`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zCknoONLZgo2vLIANS1zS3zqYyyuOfs0KD8UETMd9FpHELUHtyo7ha1vGP770/1m
rTiC3kcmotuFqA4454m5XsuRVyiLDO2EDtS1r4SFDSI4zy6/qtLcPiKrg4AogLFQ
cxwSgLSxfqsJNqgTrRB1wxLdBOjN8m/uqBQ00gg8AhBN+XPlM/aoBRtp8wFW+VXJ
TXhpUB8/fKlEhJmr+Wa6rrFnPhreaoYFTsNtGU2ZuXvK4CaAkG+j68W12LeeRcEO
AQSlo+X5oIEQFoqeFqwJ2Jd3kM/770Y8WNP7nlioTrugA15F7d3E0Etcn7//ivGx
nS44TtFjkkYKX9vIgbtWBg==
`protect END_PROTECTED
