`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lx9RtF0W8+Vjbt20mV5U80ncYN3B5bWDXg6lF21YYVZW1X/hOR4NJ52100G5pyY5
RuhDfKh0rtBVgtiq5A9O0zxpnAap9mp+GAATkTlsSgnHC+Zaznor4trMnVBVy+3y
qqAF/hR+zvgcJone3EVi71FuEWrRIpD/gJ5PETd8IQSe0ZBwWnCqUCt6OD0bS6gI
vgHFWPRuRhaYPdL0Lzh1IRsBIm7xJQnQdb8Ut2+c5aMmvb5kD1wwDTVXTsHNL2jl
cDcp8ZJm+cj2qvR/VMh+COLd0CDePDM3Rfre78W/w+FopDkIExRalgjdCF7DAowR
si243BAhQr+vULHUmtQsTL/HX1fe9S/AjiC2nf7EK3VYwq0a3zPgNvKzQ8GGVimf
98bgQTJ22xLvTpq5IkvS9iEKKCcVrJFBDCewyuNsHCAGEqf+l4ZOkfhpo5rCt/tj
AOHzK47LEDYkJVwX9Q5W6DHVCDMq41BaPr25Ln/MfYc=
`protect END_PROTECTED
