`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vo0wGyeZLDPrSNNUqmqy5/pS3nkhGZM8S1pGdLCp1HNTENanNY0u7VBRdDgQjJ9V
ULsbCedycdDJWFUigQ9JBh0J3ltp4fUFMhYaQ+f0s8BCokw8hQH++ytCiqSjVexF
scOCk8EdVOmh03GuTHNHxbikfTCDYTcWjnuvs5yjJ+oDCXXya0qz1Un//y8t5GuB
d2tI7KlRvwhpyt45myeDy9u2mcumlaMA+heKfScbMg9CT/uWwSA/n5v1ee5W9R/u
wHQRAaY8r6FxKy0Fna27vCiX3Swv/X4fnjwyu75IrQvmULJ5Krad/SKOO5VDX2CC
IWqsRsPQiFKPuVlb00z/EBbgNZ5bllSTbEMSMw+pGkUfPrJjiqiyote7aOrxNwkU
uKCKkTA42glokwjymvj6rDjo60NRkJ0QnAs4DbPopCfXz9MBc5LW4UB5x/e0XUGT
6GEZI4h/mDrCQDgChvLIPJd30DlLpiI+YvC8IAdODH7j5UCUdMSRwfc/rZpF2MI3
ZUlGHFvU1ufPsjTcYMDfeozCPSErRoAjvCtPtqFXukHKBh/39Hj5jPvCQ55SKMk5
u36gw/U6YAkLeOCY60lDVTnywosUq1YpKAeyOx/g53K1HEObd9Z2y9pk/ufZMjXw
eXqchj3VaCTsPyH45SfGzYRxCBihFxpGnHufHuJ6UP7ZGcLmgu9uMHEKVsM7v36s
wSpRPkwv6JY74IA60k8/MDr6XmbrcUni7oL+4PO/evgGBmZOcSo2KSGpntQbg27v
nozr/kPYOG/ViNGG6s7rHNspRUpDuyIPT+Y7ENFCjHSH2FwWoVpfQyUrTdJ7lbLT
T6z0tEdtcy4EK/Fc5S3D3Rw8L2gUPBllPYSoSPySm6MGuoThMkqxVOLd5AfF85BW
Njs16qiSMWCMF6kJztFuk4BI3QeZ06BDgE6TH1S7nmM=
`protect END_PROTECTED
