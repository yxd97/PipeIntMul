`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMMiZBn9YzYDYkgbFRzjNKWCkkFs0PN+O3OiunURviojeWSlIc4ls8nVcfy6V4Cd
lkMBRDTY3Ahsc0Vm4cxDJVLRCjP7eZcTlOCZcG68sOD38iW7/ID4sZ/jI3cNxF2I
STpHvxURKlf6oT6YO56cVFXhBk7x0QNUHC0SBFAwZ5smr80pYcijvy7rI3+4T0W8
2DEcnMM3QgdLGiT6NyFVQqm0tg7Kl1W1Mldb8HDae3wl2ub7Z/Ga+Lsyez9D4Mlv
gf6s90RH2dUoXHIBOuAQNo4z+/gdHuHlT+mU/QxaUJd9NPi9GDJT23dfcyC/nORv
`protect END_PROTECTED
