`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
72mKcd0/9zHEh8rnkdi/8Np+Lja3Qo6vGOU4ikyUrce5oplBmIWI7GnvrmShRws5
yPRAurF9yUBHwvwY/cNSdrP/nIonIKVF07w3ydRxJUu2zTPf9ATR6JdGNRm4gr3n
iAINWvBNI26ZhDUkwbu6+p1s0wf6AV783azl+vRB8zdHc64T5PuOQIacERRJts+k
6lNLjJss76SpsA/2LNtCakD4Z8Wqb9/+09X/IgBxcjC1uQtuk4ZFWsmhMNbBFhxw
JDEH/ltmfolHSdjLVKdbTX+2BVB3UkxXBai8aJ0DEGYeosREDF+21ZkPDEBgiP4c
7dFnr0p40ncv/9SETZIbiol9I3Mw50CrqCQEHWtuK2hcVyC+ty+yJjJprHGTyJPm
3a1ArX0ZX840+OV9QbJXw6cG9z9XzD1Q6C38kaw5vUeV2PaIF5skqQ5sS/qyJHOl
JvySSZXAanOvlL+W1CwWiK1mtTrpTWRAdmRO86ZSoc/HaAOWyMYZeMsQ8ADrWITj
XKtdo1MtTgjYOtG+jRv9gvvdwkMPFNo1bKFZRNvUiOeCu63xs+0JNjLxf18k0v91
`protect END_PROTECTED
