`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vr23wJYoJCnpeVYzf2mpeaE8loEQjpnJ82ABG5dXBPfjQ7X3/vQb/Wg8WWHIBOtO
b9z32JiXVHEjrA7uSG0a/ACE31hGBpPuerkYvA+74tZ76xcXdrdPkj1w55sGSaqS
fBRRmM251YlsPvtr7YeEU57Kmc6zwTGAtO+EeCilopEUPR7YvehllEZL+myJxyuy
4X+/I2nro0aFxwRQ+LlEQAP0qn6WteKk7RSr4x9EJ9D+QPpHsGzJUQwK2NvbdJLe
QrP+qeUwOUUm+ISD/oToPKq/x4rNQgD0dU9O4yNCGRRGnjxFM02S1jE+bbXGOsiT
MBUKiQ0H6wkR4zkPFV+OinSI3EFY/mHML2bTEFrR11UAJ6hGHN+i1JmHXcPfV1CQ
bI/QqmPg/2su9rKpsuNWATVeS45Do7AXwjJEVgZ2MZUzofrj76iviLdK53a4PgnQ
oFia2rWul3Vejo5jUS+m8GKQwQcSJTiJf5LKDtHFBzh7Ue0L9iVwSt7tvb2D6klZ
FIA/03m8ubGp1uh9qpZkzct5J/+JcqFp491lO4ofyLG/48nxslNsmeY2APqqZYDW
JaujkISk+1um9oULye/cDA==
`protect END_PROTECTED
