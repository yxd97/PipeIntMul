`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+46o2XoIuotVZkgsGVKyzbGGNA77UnrrbqeStnes3vTeCcwCBHM4LcRakfC4VIXq
CHduLUXqahDdOXz4OP3B9cZFVUGQRn7y3HiFra/HNaSjon5TwNAbjtQUZ3fA0yB5
eHze9blVyDi6ll2rAH54ap0NKRElQp16Nb/A8iNIYbjcta/vlp7d6cJZTwv0sx6a
p/3FLVm19QCS7h25I5fLw0QU8XWN0nXFL1Dx86GJ38YN8bdpl2GI6ayzwPLbUjmm
cm9nJAUfJR6SJYMa3wJg38mKDfsZIY/qGLhVNg9L5lAqD9HMYbQ+uad3Uc6Io4Pu
4I6bk1tJaUcxh/f98HQhIdenANNduWuygv4OYqubyAT1CgJCtYVYnlmzojskoK50
+1VkekOiZ7MhA5mZCxKp03oeAP4HLBJzT92S0R0dzt92x8b1mO/ZmKn2RWkwvtlP
TEdE96ywzMjQF71RE2pGkgiHPr0WvJxr5DyooCvNBQK3emrKpvpd9NtQNPvOCXPb
axvxGgGpdcZEpAxHE3aiEAuSTiENcaF9JA+KGUG7G9ZJtKkLZMLcqnXW9uI7d4Nu
XBSXM5gjB8OfN2wCGh4THkd9ura3InWmjsET8fLda5hpeawQrc1qtWqILuwvq0xz
wVMNpso7QLYmjGRQbpkvgLUXva1rws6szl5xDTs4FRYsfS2SAgttGgoeZ18tedUQ
2rgzGgEtGCM2sQjpddoDNFkwMR7XCk952ZyJjllXkg3ww4SJbfd9JFRigr+rYEj3
AFoPSxJ9F2Bv2mAEntr2DEz8l4KyqyahrgnjO50fNH2iduwCe3XDUht/MC+C+CcY
bC8dg7SJNFOwjVbLtypAC5RkrdqjrYp3PXs3UDn29JIeADpurKrUEHZ0dSuX/f7O
ZIZI6ItOhuiXkkAwvngZ/HYDGQ3p8flZJ3ru/EfwnCDmjFEDP4/ls1mlbfYwrkG/
3tYm8QTbQJT5SSw0imPJNwnOsukKyZ0iwAuEDEpN8R8FlLe9VlsPHPrFlxu2fdzP
J1nH34IgejZwQXrBaz4BGEUnSVMpbIeGwMIbLG12qQZp8yIT+EYbduCyh93HQ/EP
b20Qwv1tlN+sa5nfafqXDfm69jlreE45fUzMQ4wKqJ6Mc9+3RANHLSeBV0llGv0O
rfRLsjO/GJyIZQcqLbKeM7OA3VoBfDOvUC5q/AB4jLyDcearIUGLGoBOT5bGI39K
c9AcQ6AicAFCrOK7QJ4E5FPWnVB0V9uGihwIrfC8fWAwxe8A8sdj+MSHZ9U4flyB
SR/R1bkbNs/8vPDN1iIL9zfa8ZD2+2CmKHGO557tEpr2FQcYrP34jcnXFGclso5n
LKd5ZnrSuG/V0ZeuUbyNeAMBgnrY6fRHts0g4V7Im2SPLr0s/HB7TscQv457Cp6w
Qhv7LHeJ1O9TN1Cln5q8eY3qdSIA8OPVJi8kXr8xUsoORVgRXeQrQ6DvNiUfxDhJ
/9UnOnE+ftoACuTHjPTkI2xGZ4W6SpZ2kOL9/XYau3H6yUREtr7b2JQIgvHbKHz7
d+KiWNm/zSwJN60WrwffuELzyaRhEcOz8DNN7i3zIMXtyS/IEnyQb7mE/CNILM10
HplVT3m+h9F9VcZAZ29GFB3ymswbWUiigPtPt+rU631rp2CUnxbG7UuSU7UjvnM3
mGIcKCwfK7j20SHIFte7YFeINZgvDqtGWXuNx1XUWbwnQRTq2iEt1HYhyJG7bMjm
32HJ8u4i8MY0PLLvivvJVuX7IW9OYR8zpJFXabPEaGIThs8hWgY81g7Yz/t/wE0H
1kIeX7cuJbISo1T1Bf/VWT9Bx98M7YP+C1cv7mNlZo+IEjnBI5KD13T1SWS5FRQ1
XSdBrck7pp2TLXfvc/pIcc/I6M3a3XrJE3bca5nB/x3yWLpzRJdJmM/wIV7yZ1dk
H+iboW+8l+Sbc/JScK0XuTDO78tRQVMbTz87R7Z3YN3IVZ+GgFGjOi3WOdyRO2Wt
V+CapeW4ziodKZ66jF0eBJfU41z/xx6ZHlBi6fLHxrUaJKKl9y+feSRJy99CNzKP
1gEGb6aRJWb+cM2KMllpGT/LB2W+jjlskyUQ+7/RhXIlKGaz9LcUV/AAwswjqOX3
txmNhTNf85WSUU0Sf3JcQ+Zw3YgETLFq4miDBQrDuVxuA9q/leEDHdd/BB711Uez
XTs7M1eOwPbadYIzNAJa99jcUMHRAcqUzgyUyPU6mvr8GTeLFhyK7K6/sjr/fYMy
F+inP52NdMptVmTkk7B7jPN+DxhEqYJDC55/th3QAxpNpZFy1HzIbnPGiQQs1dqC
wvyQPMzJqKD9u+wmwJlIrIpU4b4BsAFAtuJUgmWfkKoURx3jzvHX8bVNpnC9NLG/
Zq4R6yIKh4ThtH9mhwqSBjDiZf7pSOP6Ef5vwY8GEEzvJZWcezETsXkWFJHZvdzW
7hIw4x9rHNdRRxhdVg/XGJN+rP23QyjUnFaFlItI2Iy0op1xA+ao43GOkct6egfm
yduZe04a9SMtbLX+dX5oJr8D12YWttCMIkPcD1oJhVAjEu8iCapdBgW+VqDQWRRf
YZrhVEc8Fo15aBPch75mNusPCSK1p8UotqiBQQr0Vy7pXP/Y6XxPSxR/epJNBTIT
0m6aJxUlKZFUCBy5aCE+0UBUL9NcqjgwVV8WM+Uf0gRGFFWM7wHe/Insln+nvIJt
eZfaS6DA3FkYLjrzsA/9/PZS0A3Ow4XuS1JL0yObLxDymHjGunKy7jIaGjR1xZe/
o5IsGZ6f+7dGqJOx8asY+SCbNRXlW2DvgmAI8AIS4YCbIV3PPBKFYEMxZJ6AB0cy
SbUfaxtPvbeR7OH4nmwuTrlCiqrq/Hh3I4ZJHuWwTME0RTpm52z93qGIAFl7hj9Z
b0yaPlWqK0sdVEYoHJlaqoQo/gZkktSiBNbULXHT90sUO603hljz2k+tmI46syMx
XUq4vK8fC8iOhgaMpnkxKJr7dXPb4gBzqsVLW1O1e+AWhBaIqFx4tl1K+24kDJo4
oUR9+hiM5q+V1Uz0bSLOCDvnW5AeoFMX003pwAMFxo44ypM3/OE+BimUwvU054K/
7XgcobtQLH/tBi6fxMwxpgU/1OeHfGQopc44Q6+6xBLbyDlFmVw4/zD6ArFPCxsa
JQpMa2LiDKtewd6+qMOIfmujtrJy2zUblNWwjYkbAGWKSh1uP8gnHLLV3WRFeMpD
8G1qI1Mdgzae8alq2KoqTfNzz5cJltl40VNi4t7oAdyxzjwgSqz3FrMicXnmouYv
PUNs1JIWDPWRg8YYB4+AMXYB2i3jU0BjcD7uhSLVEbP+RLyD3WDUUB678QUR+bKg
96WUVBIxXyIOyhehy9sH/lcxq2Az3mcQezPrUntmvGSGKYAkeoQBh49edDGI9sLX
555dinQQKcXPp1u2R5RCAZrisX9+mdPWgHNS4CU9IEcJAWbyReVvTauFh4RFbgw1
KdNx+fj68bzxy83s1KgHn9bVeqmlXcHvRnnOW5k8dx4oiNOEF73Khe/0W7Zh8631
M5PEhZx0sLUo6m+EVJ188DD1So2CQmJByKf7KyXh5LIswbpSdJgQ+M5hRKsEwnzp
HIORnQShddPJeoV6XOjD0YY0/rJJNHhcuYWw0hidQkd8adtL8H+RCS+/KA60Mucw
zEu4p0HRPaNm1Zo3O0l5d2R1REPhzB2cM3zcKIEnOkMcM6qM2V0I8LHNUmJOFn0Y
dWOpD0fFcF9KLRmmGo8zo6TlGm9Is6K8cVzWCh41+qbcOUPySvoIP5QXzy/DUO4H
5QOjNzDaivZplMK/fpy3NllAY3imIJlNrV7x8qRZN8E7aERlBcf3AIxTPaiV6i50
Pnkjyu1LWxjl5hpzgRwaU7D7CBN7wqXluoD7vxvh0U4/ALJI/VemF69WvzXEgt9s
evJ+l5eVFdxRVFb0C5wUb2FUmiPAlCoLLIRGHHq9mnYXiXqYWBUHSBosgeTfuy9H
+GTY5hOTr/uMO0U45ZGc+dnG1PtkF6Puf8c0sL+nsICh/s5euP0BVmP4qaisywZU
FmdbtXr1wBsEkinWu2AP1uVxN3KRZ2tAur9whD4lP1H4N9fKmkS14SdScgpvV4dg
bMaaK35nGnzQhjV9t4XTNUZWU0157n27K3ynN0VNtKst9nBqaOlPebVlvw+gKi+B
yUs7J+/UQaeC6aMhT5VaXY0BwYGd3x8liUFwabnNp1YtWlnVw8rVd7HJq7tAjs4d
wPSkoGWeqUwIaXd43CcEfry8xfyF3IWP1ic/9vBQjnxqCTIPE2wJdKgiDPpcalUO
okgv+qCm5bbVVNNCLvg7Tz04sNdTLz+EczBkD5+PJ8SVJdQIoNWlRWiJL7ZBVRew
KFuY2B3d1ymiTWkwMh4pjOkALgfORB9bQMKH0hBe2f9XZgQCbDzwLzDAVBHDc2Ft
yI3xATGbbVy0aBltdLsmHe2TY9fqVPxH2tYcGLCfRTyWjvfB+7K6Y3EnQ4IfaYz7
7iKwhcRwQKiPwZZcf+oWJTOyElh9zap8jfO68iKHsI2HAnrpXhuTs2hEZxuQJunj
kkWS3fUSiKOuxbZaOMFEyP5f6SA6MMGubBP/W5+3L0T9t/msn8K772e4eh4EsxaL
zGReQg/VW/RkNleSE9kyNqTMurpA/u/mK6AxQGV1PkqhalTmjAH8TrMpwg3ud8Yu
24xcK+e9lvsd1HrZ5GCvNYadNp1va+K/dKcNrJJu4mPWHkVabPwpndHiT1XEZaj5
DBxs7cjYC8XxRVXsDOwXoIP+f3oSkOcOa/Q04Nw4Ti8CNsN9i4UBU83EI/286C1m
8NVHZFGkLSuY6etKfCKkxDvlvePNZdV4/Ga/tTRwCPhTQuce7a0/lfslV86Reb/I
agLUphEGRTNmtP8ovO1OZ1Eltke5sSKc2wiOX0kIzxqOgzvJdV0y9gIhzQNXnolY
S8NKMUir84kmI9WtRaTz/HYRdbSVtz7ABnJ7FDpzZi5j7nrhSO1V39NJGUgUP9MC
7e3qdWGYrTnUQVtGULKvacHpY4DJO6YEq2ebHvLs8j2DW2mT5FMaLEqqe4n00Joa
7qw+wjGkeGrAC9T/D4gFv09EdRTu+brjSWM6PCbvca62vlNs3kYXhaqcQW0QftSi
1xfvNAcjM2karbnD9qoCT8GM+EWHaIDUSh2uQfoRKj4TDrhiB0xyYD8CrzC2e/g9
cS3/VJ5IC9NthHe60wr1WY5sWeEqGjwzQxC4QeDyuwAO4pTfQx/VL5urZQW/HYaE
OQQ41XJ5rQzfMAtNTSA2MqjhfpwgRzbDrr4IQHpqe01xCGgzOK31kQDWehqvA3Ol
4paky2PLfXOA2rouX14OiHwyRoEhKIBc6vn+dKpCQ70WZp4qHm7pkVOltBTaNFNO
b+rfNQpQiF2y2HqSCnsVdsqzH8b7MiUX+HNG5wl2AsPFmL7VZlePQEC4Guy1hlRs
FkGlJtOlJbUfeBHLgqNaEtWj0psMMXZjcKQfhYWoBucwC/weiii8QVZGa/M89PRY
xzgvdpKGcvmvb4r6CjZI63WPo/E5INwgPP0bDCviusM1889Kvkqoehqi1RYIlTBS
r2uo741b2AGWoqri7I7EfTRPVLk9/a7x3YcOi7fOpolxEsyZM+2SMRsNaU4v5UcX
CCK4LpSuTzmGYghzHGaxbn7dBXhPn0jQa7IbMO0NKFIjyDPOs/5Z1f6rPWF+QOpL
QFmz/0Yi1jdFMRnus37X59aJ82gZVeImrqrnwwf/UAfQfNTIh+0kDBjxYl9XKlDe
wJd7ua0GzvKqv2AE1yaw7Ktl6k8l6XW0OnGMeo2FnGlQoxWbmOwbBFuUffIXX7Fl
XTCI8Ftxb2oFryPteQOUxHWfIYqI1lUdIHsPJ1xsryOIPYnLpfZDeeaZ2HQum4CO
sZPmypfMsQ4TrkpJ712L8ZOU2rvGuda/aCkyxNPJR9xcjmWtiak3YFrehiprrawj
Ze9w4sMu4TdwGLfSbvwzcAAVZGZGrsp94PuOSYLSLi6ZkqdAOu03xRfr7j6asUBJ
+EIcgkSY+0Kt7VQDMIOzipLaolDAlar5xmQZXe7KtTALooh4SF4VgrobaaVYtd1I
ZFhaKt5qvr7907WNui2io0ZloP7Vxok+bq3ALlUaJTdhzyXwFHP5fB6Yn0lBjBy+
48g2doNX5rcxN5OSWMm81A9iL1Dkq5P3/4osyWuE9JLU0o+tKyLQF3/owFfLTaVe
RZXRQz4Q7Ajngj3yozwmc6ZMCFKNDHT7lf6r36O6ekn8cqWLuW4/5RNhNIuuowVD
pBCAiMgTNmU7scamCdNB7qEb10VV+H2JePpsO8zQb5Xn1lF5IgWx/ie9fZBIVZKQ
c7Ri45BkSLfd+TA2yivCUQbqNCWD5KElvhz0UkewZLDdrKm5af2dt7mpLkN7EhuC
D+v4gZRXcW05D3GSClv/D2jXvEW+dq8p8iM66niI8e39Y2iP9gfNXB5ql4iFQx21
r7pGBWOepRG78g5D3pg9rqdbs0T6ITidQHfuvt88HEeHzecjnUqwSkUputOs8aku
lCQCtnx12mywgzvMypIvR/SUaal3t79/W2TfHgPHNTyhTxHNYuUHRnZxmS0kIa4K
Shms1WlfHRLpDth3ZNbvQ7kZkdbKudTG9qo5LWiH+0uv2oA0Z4lYVXz6eidb7Cf8
gMBoEO6dNFKfscgZaLy/8k1rIOhUngsYHcX3/SzDaXMff/gUgld9tvZorbVqZp2D
U2yXOcXShgY75U9wDzOwPlkiPwDt6Ll8gsCp2ZVTdIWhw+DP34ziAXYg7Kbk9h5h
BK+Z8BmOjbhqujLjh3YdVEHtwknkqceeQOw1FErp8aj8xpVzcTGQO4aemHaGBfHp
yuzl/6JTdn6PTSlfxb24z8Z0bFXClpwN9gZVQ0BFUfGuDwts69/LARzNgxAiyqc/
Y5QZOwI///Imb8kZ1pf3e/gJe3KmJInYf+LUgFxX9sOjocoVMIIJHA6zjk14Xymx
mcjzSnNXX234HhKIhbjVeRPRmrgkaWi+vdq+4s9W/gDQKzwHAGVWFgtP4Etnp4Sy
xKEZ998sZWTC34U5ryjWauYoolt+zm7lxVD7S3/TP8506aWaylSfZaA0qS1eqJM4
//ZdmI9RTyI5neELfUiqGfpLEB7gENqBkBzG0IIDqRLk7jRAv17pH4n6GE7JahiN
xNc7e/A36pZD780/IUiJ/yJk+NXrg4n+oenxQ1KSLtfpMTYzef8PRhnn2Kn4iRGG
3Hb+77basLRJP11bDjVMtISspEdCnVCpdq3n/NdVJcNZJ62NzB+r6DfLR5j1ULCe
Vh5VDjQQb6xtp4TUaxVocWtv3dCUM+2xOrCSJ33i7ba7LqfzKtm70iZ4Z47MwjDo
rjNeMMngH6G1YOCfhOhtMbCdXcEHhTJZyhjyCUv3FGqYBL2kbMXTUoza5xxsw3DX
d5o8LrZO7WmkdlXvKfk5Salgx3mX3PJCXhoOjPSykJapdDBhoxNm96V7ejBRnC9L
E/ssSoIewu+FiBqqwmPJJkyqMfftslBpqhqedqUzYAmdFtTUQ65XCx7c1c/IQgS+
qpNFELBPDOtnGZ4H4Jjfq4upNmH501JoS6tQ8ZbN00ZauxusoetI9DlPsalqoOqC
T4RtOIfuCaZLz8NKqj4GW8fLs6LKa6b2jo0d8QgPj501Mah6WGOfcCfkrmf56EBO
bAPJWWok/tiPQZGmlM8EOIq4jzCK1UWf4ohGC+GJvktszT3UygdFkf5nGVBOEkia
ZUKPYy4EtycXTQ8QVC+pdCkfb4iRIWSkmuYuftAjT0fLOLcSsG2bNQCtTD4vmCzR
CZcCQCxz1z5qGdPDOYUV1i5LU2cPrfwoP6mNY8aAn3mkpCyJmQbmx7uHC0GpZgEV
MVylhiltyJ5Ae9SpWjKw5qfHf5AbWKBsPW3MZ3oK37ZDbkmmNLPIm+EZUTck60f+
vdPa3xYr5DAvslf3qJCxkRxbaXvGAJqSmKjZdnmqlfaIf26i4dotC+RcQ0yNLdKl
EFj22lTyobcmMMqxXSVga9hHKnvAkN1zKiJ9Y7V1HxyjdoI5JgVTHLg9kuHj7JfR
+XilbLpBVCdt0KK7KNbTQnF4BttRFi7/yjlHc8Gyh222q34o6mSifrHApUK/xgzn
TzIFrX2QSRyf0v5eCHPbHKwihBvf1EX8o8Fsk8haxgz39u8zaZ2rrXrK/rVFk12I
wKiiNx81yKUP3jiD6HJpDxwa6R3G9/CDmesxTKIv6xtZ+ibdkjrh3C8oBjR0OK/R
FNDqabY9/lwKA0JacLij6S/XezhBjvh/sq+h6AAg6LqS8u2MUmEwd0KUbFYSvSl2
TgbaB2pHXiijkT5ak9+mEMwyzyDJxKx2GrdbC+TSi6r+J5T51dpv9ub8nPMUxN2A
xeiOZW+jsg19Ry+x5QXC2SD7VrSCtJ38pu1sJivp2WPbBMcmnSEyrYkJ1uEK5YRW
xR1tR8pgtRoL37c5/QqJtl7gWagnQ72prpBBDh4Yx+joTmRm+88VOGaagUDMczvA
GFYmaZryT+jJh7JZaTC7w01r04AoJITOZmwRFk2crEodaC5IT8nbrZvoED2VMpmy
zcDjhWHvzlH1znHIBYrfaQkVezXgRFmQpyYcTF+o1H8oFxotiyYp+sxlZ8O1KHDX
K3/js7hBPucj3Tr+DSUmNzaIO6RNoNLywFZ5HBXcsCwNTLk5lBuKFPlvWLoe4eR2
S9GAhU/D+sCn3mWPnp9VI06j+bXW6PUrax6lNvbrIqwGjNRdyfIjBtHyVh0BSCnW
hegX/WY/qqbc68EeBkVxOd5Ny2pYqbNhYZLYVK/77EIbqdP0LDOjfCql2On6IJO0
Fyqoj95ZfknDE1eyyYmjv6lFzKaKgpDYy4fadJSpPn0n4MNznaaXpky/iCNQbHRT
iAM590wf4TmhSm2inENtcrPTBcVVdqKyl77ONMPYj8KVrt8uM7sxFelc9EVTt2h+
TNG3VaG4uzu/MMVTNdgZ/cJKPPk1FdKjbMGJIYvrrw2oNc23gryF/vkzcJDzxTHy
3TTEz3PdLFGgYZqYdLhKfJtN6qCDZuvWbjCcw8keLlGrg78i4RCB28YmiTAk++i7
4R4ARlYrl1Ucr0RSmYu7gMLiJdzQTUwJYBK2ctOzzFjwuF7e1Ppy/qkMmkpwH6hx
yHmzflWWC4XofXNKou5De4D9EsJ5XiWF3DPwyOvE8DXPb5zLQfVtO2PPeqTDUlrI
cgVC/m9+4+FpkSd4D9OGC9HlapzJqWJ9KSl0QCSTBRzp0BNIWY3S7PsOTZuoaVFk
9FpBiJRF9EAdheoGtwNYMax5A5ovZvULrKx4DveGYB1BPE68zgV8L/GPOEDD99eT
erWTpKRDqyBgetFRw5WceunfizQx7uzR+Fi9YZCOY+jAmwYTOOT596RR3GQy9/Iu
sUda0rglikXKV65bsJRzstRaa9xrEo8EnKbp9q5iptOx6CDiInIy8Td7wOIQwbEs
n2sDAzpEjbm7pCk5paitBdoZWDXqFOOqvG4RwfDFErQqQe4AeTVReyf2VqHqJwyh
c1RWUuZFnempIAdbsNgIqem1LpX9mF1IQMJ//7GfiidjX8CO5EzmHhRR3R5iFizS
RW581Fu77mLsWm6iMacWqaolYjWljFnnYtX0XNaTn0p2bw0LF2XSm83At35nWB27
`protect END_PROTECTED
