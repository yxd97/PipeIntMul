`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCqYiUx5hnOhhgS9QgtK2hy4XRCIFf4zoDjEEJvbv6KzfvZDdX5WITbafpUeMco7
r2roggIFP5RnXNqxEfhc8zhU8DVQNbCYwBROwbM+sRty+fhfg7rivqhynzxfAM5/
FC6Oho4cyotmC7qJovrLLKm9dtV0MQpjX7NrVYXXwH6xGSP+17zh4R/832t25yX4
zc5RiNG6YXkvRT5/wPXvwcrCtyOovdp+D9SoKQOxJtzGl6aSaXJJgHIBn42b8Rsi
ZhlcUbJF4q0CCsfL1PHA1bwHVAWtzKvOu7z49XELd1v0goKrQrqA80E8tUOv41eq
UYkWtENMRBicH2x7c8uH4wV4qWlzgnX1AVmZDilWC7gfcBY59V79d1ikbbVxiIap
wgH8g2uvJQ67GPAWiWVKyRVyExNCAk1psxykRECH088HNicZvhMYE8PuYbhLpIG5
e0BwW/X96bWQI6yaCdYfe0baYKV8Dy6yUSNQdGG02GDxmCf1EdwqiL5znOlc2N/o
MTszsOk7AjryR2dM24zJtrxULLNYRPVzB3ZeheJkuiX8/674BXTU/uZf9/ltI0N1
FDLaxtWmmeeMUfcS8cTRrcJWgsL7ATry25lnuaVluDo=
`protect END_PROTECTED
