`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ng78qMbcWGqwNioa7GXTye9AbGZaXUu8j/uRfbhRjHe2dWH223xNISvFyQulmAQx
kj/mA+5izVawlnV4IF4DaI7FOS//qn5v24muZOSQocOwfSAbCm5WC/T1aoAu59Bg
N82tJFRGMjK8fBSu4B6NL/nOCyuwCdN+MvbOCux6Nv2+OAV+KtAZD8Aw9sIOYSFG
Us5qXnWb03gz839RR0C237AWWxuU0OGRSEYwUSt7Yj90DHzPRxdnlszP2fh74txq
UYnScOZtEsCwZNWm60b90IE/tds3kNXh0jhv0kx43r4o+I7hXPdkzjf8qt6SXcvc
/QUsfLelRkqXahIOBgbsJTddw70yesqSq4Y+ARGiE6nFaRTkoeq/LbQ+1ieOmY/M
XiwWGgdYfpxsRFqFJcu8fznYeqFqN+vGZ06sHzjmxM2xOpKpTJ03ayxTVLuLRK1U
BYgL7m+UOyS3VlBwmXKXjIwTug/jfYmiJaJnooaaU96aE4doAuJ1DKTo87ZZIFd0
BiUkhhaO4VKSSDThlcRYRbMRa7bCZC8MdkxvgqXU7O7qEfUZdz4QzxgyJdAy9lk/
kO8smPavcaUz1Y2WTi11P/ogK42soAzLpr3YR1pgBGlEHQxERUebvGA1OlBJfleN
MCZR4UcHB8lKEDdp9YIoAiAZsg/BAX8bjR5OWZiv1o4lUkYIHdBxTRKdf7qH7aMR
bG8ZOxMzsLqH4BrUQ5J0/SECGsbe0RTu2dnm46L7bzcRyF1V7XawRF3369IlcoEx
L2oI21OJDqpTFiQ2sRh3J06J62IfSHFzJEJFbo4a4lOCzRlqKwTF2DUGhtvezmaT
3i7G52R5kRQkErsh78W9A4o6AaFy69VReGx0Bvi9QBpIKlcCLt6ldrX06KeTPKce
p4btiLS9K6V1YHK3j8n/+poNBisMa2tGXCpGa5ivfQqFpSVpANMsNp3jwTNMhhv1
SkXFb/U4JK1JICNpw6oDvGIVjW0jeycEPeOTPzvtjKhSecYwaFx1Ofo6vMmvLO62
1Yv+FIZO/Jo8WB5/x8jb3t6ncIQw2fCPFvycRtFGWR6PZ2LSi/X8ZrJK16IiTzl0
LjnHgpvb+7OPmyCePSV/CACyEquEkcIsR+e0I56cMMxyvYiePeXOkQwESuwUFgx3
iGCxsth5/40MrPqoeHS1E/hYLiJc39Ute5EWjUMzJhgnwz8lgJRnYNVDAtjCFbye
sI7VPiwEsl2g6Ly0ebKjtOmbmMka3Dp4XY7BwuG1MHJzoSD+jmocw3dCAXboM3oX
Lle5wYpNVGIG4xCEoprRLxEdeHr6q+ljya4WWiCP9TwzI/9a7+OWOP8GeSLdxUBC
iKtWUsEMLr2V6vBtjbs0eFL4dzpI/5h/PoWdo5G+SlNZPMUSYJKPUNo3xSDVd5In
ZOilZfjxORerXuY95LsNcvVKx34erokAr06cross8WPvqN8X5hi7WWCSjJ5wCs5A
+k/K6k/EBLNa+iZiK0HI+k1BeLSIODMS4S5lJumMbeA4FC3GdraqBlD8WqpTMMHm
mtHw2EDgUwU1s0nUfWWMqwbKQcVgFwthB3Ek3OHBNqt02j4+lP+cH/KGl60kMFcu
fZRgmGSOX2/oPI4/SSaS80M93BaQDau4SnfkZmngu737T8DCzJ3jDhB9V/2/cyWn
tXnDmNYOtWXOAOUjY2IiUibgC+/uIxP1bSxcmnoQKLEMipdGE6SXzfHcotN1V/et
lLP7gFL8BIUzmWHUcXZbUbopvCy6rjXjVbCC5K88C4EtfimgLa+6MySc+N1mOEIh
kfPexFHf5amzJJd4GMWfC55HOrzOOrkxAhjdg6T3xcNiWBXi+b/w5rgdqNiok2D6
lTKPHZ9twhSFG8hJMGxlIe+aIflcolK84VYJP66TQCBP2hXfts9MZ7DaHHnU6NT4
G7SWNaQSy1Zfqq6WKzAfeSbsVtbIfbFhaSCPw0M/Wkw2tfV1KapfO9qan7PQz15n
VLjDsiykS2MTTS5XM/vfjn+s6nuRfz6L6tH3/cfLXR1DoKgNXFagLtwomZBan0QS
pKHeZJoWmfA93CoyuUp0pHQs2nNzl+zB7YVkz0vfDe4uLUuPBilvqRxOyj1XH9ky
pBQYYc7+VIONumsSAtr0+387w6O7yZIfQ/5fbEumHee+2grHj12Lkce+1x8V0FUe
URhP+5TYP9EZm8gkFG8xmpbVjDpqfH4TpkBXHG9qb3E8ohZp/Q4RG9v7ZvB69h9S
`protect END_PROTECTED
