`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xvxEu55Y7/B6vkyXrSzcQtexx1+tq+6X9GetE0xvkzWAKSF+EAIZRSxrR1i3O4OF
jSfzje+C0tEPu4tqKgaY2HjWRc4HOVP30nCAzLa2A1QGa4i3jd2VES3yvLn2yMef
B0QXNV2ESJ4OwIZGTrRClrOqhrs6PkT4BBALqF2iej/+cQQPwq3JgMxGlVaAbnAw
g+h+KzMskjniAL0Q/4gjKrNnvxmv/fCxAtJljZ+ERunUZVmE4OwepJmxSTan6ryH
VgL5DHX5pXUrqZPzZ7rszISiYZrJ7Qzg+fP0nYSEyP8ZDaspvHd4oIw7rm9I1ypq
5/Js3ClCySXa2PAd1Hq9Jvvv9l3Yt4aL3cDx76kS1FAQqFAXV+hqD+RBALUOSwrA
ccLeSROFRaWPq9bz0WL6T9zm5i/aNb9BVVv66sBPFxOn4WmgMGtcad56a16CBZBg
KvmvGzffdZU1aMRuiSXv6URg0MSMcm8FMEORqrEN+9RcpzIqXZeNR2euS/HJQ9BK
6jsxYqVWe4NgMRZ1BaL0DlwGJHYZXYJt4sOVG6fvpSI=
`protect END_PROTECTED
