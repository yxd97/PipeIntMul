`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hcsiWS5szMAkntPY6vkSQ16RtRT7SSoGhdc4WxIy77fEi1S0qeZ9J49yZkgb19Mm
faQ6QIgVV+9vHmn+iBlFyxwJbj6yzCtFWYx5pwgyTdwU0vAuZ1czHfeFLeRh39IV
gEnoFOxgjDeKVs3MRZPsi+2jmKrHYHPIXKkCFO0xt9PDQUBzB0/Ez3c3K1Z4j0Z7
4QY8oe6uXUwHx0PqQESq569ePSP/MRL0aMU1Q7+hnt6si1TehjiW5vIa2Iq7NiAL
/27I/iCkQANeCQ2LKsgFac33xBsmMrj2y0mU2FprGlhriFaNDwg8M+wfDe1j1FB2
O07FLk575EW985s0AvaiwQL6v076fVM+o0AizKZxiFYbueqwYgKY8E2lkMMZBfDf
z9FUMFLGLI+NfkM16bphoV30pfYJOBravUrF2f/lTrBhmdnxJq8eBs2uJfzteWio
1yplqJSaGMRIxX1mLMSH/zaJrDqMEmRJcPbnx5txd+MqDDanczVrxr84cB5IfGZq
I8TnyWmMUSMMJ7K/4BmdCR7h9FNPpIX9q8kJwOyfaoJdD+JNK75ZSAS5wyxdo8UT
g0XC1pwDH0o7hATvsdxBoJyhVNgzZWGheDGUQaXcGqMF8be3eP3HybVg/nhIogn+
y9e21tGrjAFtamNmEoP1YwFrJn4L0YDUy2AB5jSIalqJsOyO1k4/Vr99N80riNol
2Flf/xsq4pSs6w9UxuWxCboEA0IFp24GbDE5pwjuwLTquw2b8Km9eZQTqEWiL3vk
HiuD+cCqtWa3HkmYxnnt+B9zosPGpv6gBiK/IErqDiGF0Y9bLTOLGCP6Tk8IfupO
re0RCVfk+IJmMpaTrCk9dp4kIyLkuTnOxMoCIeHqVd4pV4QZB1Eh2oeDg6PvFZ/J
4sYNSFA37o/MSOaE1hjb4JgBxBmm68xTQGw2H3KuLT3+lRElvN+klSRszDPfbsGN
v4Fs2Z3Eomkm/8mlxuDrj9UfVEvRZLZknsv/sOUkBnp4Go32wSF8lQlXYildyt3g
EVVkQ6nVPWWiPIxVCtIPWe38mV0dBRHIQDL54qfMTCsRcqXU2Xuz9nj0dICKOVAD
`protect END_PROTECTED
