`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zckNrJH7gjysw2qyKqOEzZQexXTKshtoQw52kQc7Q+6dKXTWpjK0896IQzV2F4vr
WpV0EYJqxUF9QBagMBfyi0PIy73PSULDZ5LksCm4/jKFpG7gIwatfpp7+Bkt7wo+
pK7cRER1ew+FFRb6XQ5n+H1QaLHf9TaPhnoaOl7mJIInZx4D02UpG1jVBmE/pLRi
yc+0d5Y7D9fiDLSVGhz3gelGTiqaADANtGZNOuYg3MpS7jLQMlYauEOZHyRDUtvw
vQmf1XSEhak+xGkgjWMvqBFGuVTMZ6bTv8ff/UJvmpn7yzea5C4pMQmYF8ppeUbp
/YYwsOqlNUCDKKiJIVQoyGlewGPO7UeI2j8HJr8AcLC3DNEfZi6Qp0o79foNJ8MC
MrdLE7+u8RYs9v91xmsPPCrVF0ibN7ysXTz/4e7WlsYXprMJLLOj8hEG+He0dSZ3
oQhIpca5OIzRIMWzJlfWJj0bpmX5NFaV4Pv+JkPxGEXYSV+dJkgGhQ7bOQ/M8tLI
EGnvX7ksA/vg9e/XMNo8yaO8ZlE5nW2s9T00uv5pw2+cU2VR0MFStrvItHzOHLjl
JiMVMUCm/6Nd7LP7tPBdi5noI1HhlqVRzAH88lfDb45nfWatPeUJol5FAqvPTUwT
`protect END_PROTECTED
