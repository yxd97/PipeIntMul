`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLzjx1KC5sMMjtPzc/ZDrz/jX88s274KCf4Wq2hyGZr60UCS5MxoOe/8BOHBnejT
yhHs2lpEJJ/kPOe+JieXgZz7/a8kkV5RtwdWkG6Sz7ZRdBb5aE7fDyA/lUwsQelj
/sktakKZodkScnHwGhS5zBXqz5Q+ImALv1+mJ0RIS/LNLLa2MNXOHx5DT05fUEF2
57aKf3R9nhu6N5dv6sP3YYCm6cqVuCPXcgen4KNKCIJlqMCuPv2v9KCL3e458BKQ
kWs2uFSX+3GVSwvlPEh0J/ruNCcdlPH8hex13RErxYk81s4KAsMke7lv1m8rNV3+
nT+ZihPRo96x8XixiismeXEFKC5fBuEsCVuSDtlkHdlQ3tvXeTdUjirCd75hXe0E
DU42RXVq6xa7+fuXRNOybX/vuBEoFtPYXbQxC/OGm4l+VWrKZv8sY57Ql56k3YRF
TY/t4VcOiDQJWHRNMYmnwk9iCw/A1QUYTuuYtTBfmWV1j/gjtdoHK5Czn74c7zoS
vLKs9qxbkoPQzMKk5epmWR+kjZWK0o+MLMnAiQLJtEUlcKIwp9lNb1lZ/uJ2cCrJ
gfKDgdzea5rq/GTBcjcDFxEEC0inLp/cKktTjb2dKviCk5xYbxkBEROgr1ZW2cxz
NDXYu78x70sc3NZM4OH7vayKERAx5wYfpxcP9LW74e8M6I41PaGW5x5s9oiye0KA
`protect END_PROTECTED
