`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuU1UziU9gtfhd9NLymuTngQ28Xtm3YKgW3A9kyTr3M2EWNK5wP/pVwX46XMSgwe
ka4T5e1i/QzUjNykRgbFalDeuWSYliCga0kOQEbVruGvmGDel1iLsFnhcpV+4Fja
oW8o+VG5yKPkrhFdouO86bkOUQlYAaXDowpZr/XL+xOTXnWKdE34auLUpQsBU+u0
yQEwbvgf5K7YJrXEpX4xRzVP+1Z1crSYX6HhaylRW+M1C7VOrJkANg1fgB0wieCl
ELkX29p9AcwltPjwsSy7kLRzqwk20+bYYywwsJS4xct+N98uX8Mku3806LfeU/ip
owu918THYZRH7OPFvjBmKw==
`protect END_PROTECTED
