`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMq5G6+lnMnBQ+KU89iIjI5x4/L0IzoROtXtcVKTv7EpGqOgN6vL7nYoG9eJ5bSZ
Y+Ol+KQz1HVDfN4VvaR7IHq77bzOXLfoQdgHEB2jzBqM7GzfjJbHFbmSGU86g0Do
o1HRnhWSs9R0dWntr6TP0ot0GEOWTswXwBbZzKNZxf4tKs329sUb1OR6I/kitmzD
wt3vEny1p8c7pQK3GYBf1ymdF3emieLP79Qmz6blCK3FtnGxdcFxjVmlLNc64hk/
E+0bqtzx3hG/meP+odMZtfO5zD0s0VBvbatIhZCsoshxXmhxSDr75wU3Di/LDLW1
AVyPcUFFbPRWZY64KNr500OREvymXGexvkDJXt8Z8o3qDsd67vWIlkPYOkwnUhKL
`protect END_PROTECTED
