`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fl6tp9ZuLIT15pe1sqCaJmtuIgPn6efHSbWmDjr06W/wzWus6dSBnriClquVEIpQ
POBCl/FXpASLswXHhppMd1GfnrLxvujSkcWhT4riEXal7Vh6zUhtMwnM4K7HhM01
AKIetBAF/9Yiwh/YKX/RRa3/uOYIC/PApM8A/cYHii1YOQ4ATh4VRLtjCvpAIqhT
z2/O6vTjZdBGyC38qZXdPMFO0uHfksMGAZZ+YzheWRkSfkx3Qr5gHtkiHqXOYemQ
LuLT8Uv63ubLz4hHLJHE+zSxEhdpnLSV0xmwOZ8qANJTf6z7YN8/hqy8OngvwGBF
j2XAAuRnu4teqb6LlFHqKXkZZKItbbaX0XxFnQ6C6yS4Eap69rVJxDfcLQJ6st97
xTMmIp8rs1AmWCw2MUul8d4HdavZqenfCGYXu2xaSwH5U3wZMRP8J2lcrUsNhdQ9
f1/W31egC4l1b6dVII70FXWgvsR0NXifh3zOKbL3cuA5kiGWzGHYc0pYX0bwwiJL
9ZM2JH9Jml43S3OtpZ3N9enrLLQL2ZGLfVRbp6Rs18Q6cYwuA0awyXZDP4R6jT0J
hHjn9RwZBWlft2JpK/ZX/B50Y8zBR50/TwsMWksszk9yDLKmh2NeOP68NY/MgkTU
FHCEoplKAasqcZDLh4V2LVa0bVPH2lndT27VH+zrb4KNs4f4CT4MHXZv4lp41L+P
7+8FCSrnksbJ1ZFh1gBMC4hOTWmxvw7la8Se44RwH7kKdWe0j8PGGdkyYhs2EJ6e
e4qMU0Vgz7VVkArnMDro3fXi2uN83uoS6ydwh5jUsGOYrvENj+ZUNcBHV/xAa3ex
ZWD/FlU/Gu4iAweiK2ZVJOBldrFhwHILm61GDuqRy4bS+wP7lsA55j5EwS+SVdA9
ZDKxPAXXXt+tTbROenNZ+Q==
`protect END_PROTECTED
