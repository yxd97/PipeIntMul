`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FnMWUSzTA8SM/sf4WTAW4Sux7kri8+Tcbw7cKlFipZTxKq7fcRuZJnUZMdUrfPre
YHA2HZFJSJ8gBjr29zDownxWEExDLCK41chHT5MfZi5d/yg/vM1HTRbl1PBFp5kC
lPd4pQoYXn0sPwuNbiRJB/y2snjR3uFdJa8etS07tozYf+ZtG7KdGToWngFSXuiJ
zEdiVFpQrIDTzlEHktx4Mhp5eV1rkHi9vfB3bTlryzm/5+IUljlLLnPFkWw80zhw
vFT7ZqGgQaYCmc8Btk6H5I/QLBOmn7OQcEqCR0DDHlDQ3EW7VDhMdOPkyA93dLcm
SF7ORfR/gA3CrSKFqcC/3i+JlIaHVBWljIsotj+J0ExgQP5DKl3nM8lFEgzTHNGV
T/1di4ZNMQdSZnZMPaYsCRCPkYEV0xZBNle1iIj831p5WyXprv4i2RpCLApUNCtS
`protect END_PROTECTED
