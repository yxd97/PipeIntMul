`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BkUtJ3YJ/ESr2vx70Bs+xUjCO40GyTEKKHOkvH+vdiS/0xzORnExtRDOMXQjDlfJ
wfDq1ZiEfteE0Pvt3STwlCiv9VqZJ8IFtDTBLFJyQgy6AbADx89aLPFW9OIx/e17
HR47spARaB6Dc5+pPkal3lkmDz7X4De6tlEPuBzmfx4v4k6YERa1bcJKVuCryOBV
obUuR0sltR4MFzzRfFvIJ4lOIfNmPbFVFmasDlLQqD7x8cEpNdnsyZo0o1E6GrIB
kIeQiro1t6+RHSD0A16D/9mcURzrMhurLwEPjwczzZZZfAgvjjQbGo6OhpcGaCxb
5qgU7x1w+7xtgAw/NGj3Th3GiYQQnrN+Dkz4CfcFw7XuIeWIm5pMHXwhnSIDKPZi
WoAajHxf771SIaQ++ytPZw==
`protect END_PROTECTED
