`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
400evKyglO/PTV4Ie7sjFK0w+yWwiqOjzy8SgG1QNFRy1kFnOf6x6lGv612aCsA+
+moitNQdyLQ6lHVCnwtfdZHY8T/fX1sdYnxGKzSggMxZiL3iTACCJZwNJf8kGVy0
vA7d7UDhDa+53H/mbQenWKE99RvKw+SQC691jmdE6nYtcAu9Pd3O3WyIM+ar6ngx
X030i5k3xYh9XQuvfGGPs61ua1l/NtuwU6CO4ZUjos/fC+HoIkLg76eFYsFlN6gE
8RgMbLcuRdwqTzk/OmeVjhkVERa3BCjTrTxUY2lODkz+vESxjGsutLgFdA2KNfER
q4AHh5j1NJK67+WeoDtFIq6JHDVEeRuuZ8RCm5pxPwRo0dA7FsYCvrv3UsLjt9vi
JwAlqPtem5xFnXLH3NT9lBdznM8YeUaHU1+lF5UiUOsPgw7I3lHU9VVJ6geUQYnL
SMr3uRjH6pL1PZAWqbNGjU7uM7T38/48x690N0gzCGk=
`protect END_PROTECTED
