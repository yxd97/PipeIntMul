`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
li1bbnm4iEmnhVoMWu4FOHOIs2ueX+vI/j5UTc5BA2XN50LW7kVJ7ZM+RKVjNR5A
UTa1XlF2bKW+BuaprkUAFZ10CSGIkp+NmE2hwp/SZP7V2c4ArNci384yS6KgtCvV
hKgXIEKpW+XtxQNrm8w58Idp5F5AZmxHOj35ePd7JmsIL09rz7DWdpeMBcSQKl7x
DLV+xxV815B85jKIiFsoHRbTf2PiGvu1KHAbz8x/YrN7L9KWnznjHBUMjEfJh/Hh
uJ43fo5ANJaH212P7psiaw==
`protect END_PROTECTED
