`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knpHJNAKU4WXDBlVBwIXMorwvEVNsj1xBYQy9Go6AzIY/Yc6iFtKKcQe6sXSlh30
sWkjYDl+SfhwH3CidyS1iDmvFHjbCvjgf1mEJ3zUZc06w/ApSI3h2aBT5bv2f0Lw
xUhj0h5xl58zZ9aR76/8GBRuEEDnbdLu5iMdQ5lCpOiNPCECivGXfgQeA+UQrAht
nEXWA2bySaB3ZE8tkJiHO9XgdTgi334Gpo5id38UFI8Jc843KHgRcZd79tdiLYd6
RK1eklLV3+qWr2DPcJQFR0q8Ki02HfPuMRFA9aOXI9Sj6XuTrGzA69MzUMHoWgV6
Np8sGzGQv8l1wr7uGuNTsJ9bJpUEDfe5kjAQAtpNztGCFXTrm2aq4bGYRDVvRk/t
c7t65mLq/uh16fG6VLFPRF69crmlRoid6HSTViIwgvsP7bz3Qd3R28nrW/hGJ/Ts
l3gzWKROLegSC3fUd+7ih8hwXXKC3ULh3vYhf6dmqtZ7Ub6CwuQSu4h2cUkCgT+2
yT8CvEATmKVih+zglhg0wc+ngdbVMZtWjVbow+Za1890J4/HebO9UcfR+bFLcR4a
jcPxfso3lioV4y1KIE8xNvSKePcDcb/nZq45/4GzdYvtfdeiLAoiuNWR4TLkXmCs
tXn9nj8vcKUPWxbr7OFHU3Zv2bjF4Vm1Ubjwan2aVQr9T6yxS40BFMir1RFfIufV
syabUYRRr07x3/f/mdlB2NWt9X6V7FrWV23bo/RKjb9syKUZMIxuePvkKYRSak/h
Ycr5VeNaeNBY0lEHl+Ir7/QWJ/DJTt0obEe2fWnb3pvgrcB9KnRcLdCJNI6eDmvH
sT86R9JPxUEKU5WEPMahP2YKSX3E3M3jZCxY7hqV6AZAdOA4CyznaI+AYP5q3uVh
o2Ja+Pl8biGHHI+s+TJdJsPUSJQHePtOJ8j7RSwE1DRAsHkp49gYrzTn+RE2t6QG
sT2ST9yZP7cyAReXjRQZyzzwN4t2/I0ZXPwRmZWrwIYlXvv4j8J5ghg0Nn/FtGug
SkU++5jK+KAf3Ds3sofMzL4gZ0k/KNcoO6Auf+1s0LQNvsyETZgAef6CY4Y/8qD/
bGSW2Yf0nhLR9QUS5Q0aekpmGLA81hLhY8xlYmEQtn2mrCjimsLryDLjyPU4jYT3
dB3kegHd7pG94CpnmqGeEQ==
`protect END_PROTECTED
