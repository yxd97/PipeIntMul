`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TV13J0QaXVt82oBePfY/mpHbZC8NKYl7G17GgP/mWm14m5Tin7gZkwkDMeUgS5Zg
rpbYzKrMmjQztGnEkncYzuzOfE5HVdjpjGYcK5MN9JFOtMfhgAkbNwUcvuoZjirx
mWlzLzePtfPzMvIvJCSP5/pLfD5gmCUgztLNPfH2oO/EPPOgEIFbSPxdgR/7ALts
A8r5RexRs+Pd/tNs8iYe8ehahjNE85iffR+VE+ejuYtESLO4wfbnb0tNye5Gb4I/
gkZ+95pzO3e+4wg4VTsPiVjI4eBsWKDcoMwpZFw5QYNxwpixi752FVOftm5cXfEz
jPIYdklERMFuxcP8CVTjmJipf3Zqj1VFFXoeW/GypQ5SHD1Icx9/686SYGleQus6
8iiF1S1cXdBuDkmhHK93bOFAbN1S/A5VbO/vHUvDVwwOJoWbpTpbUF1SeUnh9Y6D
bmbIJ/FK73JimAeSi9TBgBjx6Q3w6eSq46EsdNKTGRhYHuLd7VoAcq6DZiR7DfUj
`protect END_PROTECTED
