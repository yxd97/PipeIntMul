`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NfqnWN86wqhpGJtjktJUVaQU+x82CfYXRPCdKCViBonw0vCIenOvfD+lXDI6AoV3
JglKhaU3jhCa4WxpllnChQFRwv152FgO+tGnlwfYJJ3OBdFnLqwyGZigKrLGDXYO
qm2r4UmXWguPlucdzJjTCFLAtVBskP+FhCYqRJw5DqBThOejfbRaFkwhpTXXByMs
j3D6T+bMOWwzDUCEz2b3tglkQC7q7U3Du4p0VSizAnpTrDDTYRY6ten+RusDGE7w
mJkrr+pKWnNlKWnv7RdqP7q2QTFTZX4sAADX3JhK+Gm/LQPrcByg45J8U47amS4G
oruRwc0AGr0wLfjIGCxV2zDhezTo9E0DHm8Cw+dokdUnAxvjSEyqV5FrBQ2zAKhX
YbLvV2We55pWPT7jKM2Zscs8/Erl24F0L74+bAIQ++6wFDmGgTCm+G5OtSnWc2La
BS9E+LFAIDrg02JWRITH4wjSf8WQDIZdMf+hOBy22l0u/adjd2oI19c0gN0fM9rE
qFNRjFesi+l1G/2uw9HFib0+enDmedOV4sLq0wiVFaOQPfBi5S0yj/HVwhNowgVR
vzYYHgm4SsLRIN6bOUGrcrKkxxWIC0+TWUVnZUptp4DYi90cE5DdtuKYR706tlus
ERFRd9+TWyuNxNngPQcYMhcAB5xwXH2FMFJWCzLywPavgAELSn+MdovacwK8nKZW
l+AINv74NtSOPvpO2dvwAQ==
`protect END_PROTECTED
