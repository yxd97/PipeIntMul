`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7UL+nVr0Vd+9BK9DTmBUiWRqytwi6DhhOuBTbIfxkAvcFyMwdLwePmfkQy17s1+y
dW8CK6R2dmbzfUo5lnBWl4IL37tT3uz3F+Le73tRGWm7q8wbH6dbi9V7Iw/bCNi1
eA2U95F9wxYsbX6Bfw9XkIGjT4vsaFbOTo6sHW8ZmGWWPSwK6wVE5MOyd7I0iaqb
yG1Oa5YZzfr1Gx2QjXTvbwbDkguiughz8FUMY+vs+Gsi2EmYoUS3cQXoN6OpI+Ei
4KrP57ELG/DF6qHSelckmItsCxNADQB+SmT88VtmbcfASjmshgNOuNi7i4WSRInp
qHPDWiDAwKaYFEbZejZPrL0DVKDgARxucj3+JcpfUhvaKNJHxxkNJJvgkEWrDxvy
`protect END_PROTECTED
