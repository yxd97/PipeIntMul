`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJ+SqrVd3GCQSrFOJ0tiuVOpwLA/3LeN5CJN2+tEwAb1KmLaPDrZvEqjBsCKILDT
sx5zPXTGhyKbg5ffKGaQ1EnKMP8mOjmKezudm4O80VUpgCJSyje6v6T7p/Ukc667
vx88m+DCXE3ar6AMccI3yibPrPx+2Z6LSmlhQKOYNBiv9klCa7j5LoYJuADJAFyF
A4v6MeV7ynvw0tXuM2/qeUgMKiL4ER+sXKk9o5Kc8o2GENaQ8XBo2+IPiQToW1rV
RCv+GURpFiY8xKqXYSsx0YsRtDFhZ8x8LvyJ/70ahT0ygxqI6AsDP2hyi+2E9HRk
qmODr1693SUePmOAr7mJLRN75movuneJZI8YxNkA8wNc1hXqTr8N0dYEO15aUikT
8XlBIigpa9gJAux1MymOU5JNfNzappaG5YSuGZw1N43mxdDhZcW7Pxt821PJJkQk
pM6eEQYPbUCUG0YAMgU06+K5AtzfOpXj0SZjIjZ+3RxjBxb91ZsmQguU1pHymr2s
1yclsDQpkP7hJ5x18sHo/JH0Wb9QFATbpOzoFtyW8dI6oiPKauJuqfI9ma3Iq1Y6
uy4G9PU6Xv3upU8rrU42ocL5wODyKZak1AqV87xtN2SmZnkS0/C3T2sW+BCUUhAk
j2HX3gs3TBLFGsP3a8P2vU4/aQswwYpOZOx9lklHpgkoSLdPffUagI5Sw/YRnrJv
EyuTCTqTHm6Gwq820g5G8w==
`protect END_PROTECTED
