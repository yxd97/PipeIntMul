`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
USxJVvqCgUq7C19PBvv6yx7/NPQSrpSbxyMpw9tEA7XwF2uvOyQ4uospJdQVKBmQ
SjYP13BgqKfzejWSdnemZV9EQqPCZIPkcuInOqJhdLL34kq9h3nngDG6+iX1aVO7
nm4RyRHPLJQN05E3Wcj7jNcP1KbWW0WxtV7K71rOWwkWyvrovywzVI+hVXxZcqBw
6BiTnfd+W8sAPD0NxV7VqBkSMmqGGNKQdbxkjK3w+gz/f6AViGo7GdEKpV7imYWm
+tRcBHDlOyFqt1pZy0SB/966VaZPK33D4dNYB1WPZNXmRNF/AlwSe/WWI+NlDkz2
sMXFiF11kBFUmMGrx1DoW+Kkz6mPVYnB098eOV0dAMxaxONG9izRoiaBxgrFeg4y
0BpUQk3Xz7PKLHj6UZwkUJ4O36jQ7XDWh4Fw1WbBP3Er/yILdbRip3DsFPV3JUy2
NOk55gLp18PT/eENHieJRhodUYfQihdH46+AYUrPzAcjsOlmTFjdt+GobYpjLUXl
Lkl6LodUJptGH3BCeHxgd7vnKkEMz+ED48FuOEIJxVHpHn95Q77d6BhEQFTqV5ZA
M3ITYwX3Jyt9dnUZMTEBHviLrCwdFvFN0M8cJCsGR8BeT9bvnAqZj2y1iAiRqjpG
C/FWp6/RaQ/LEqihymWJpUMyMLzVpQpufj7O9ue6EAQvohuLVUTtD8fPIv2+GSPf
b3MKWFH4br8WW2tTjbQWsnLcZyNc7cOIfjIVh6bi911sT6NQhnA39qsJUFshx677
bbFkFcM35xfZwrwbcuxLQIEmTe1rXDfkdDY3ORZmMy7K9VNf7vZZXIKZWjpCDOtP
H6sFI3X4Ts7Yuq8MbDEYPw==
`protect END_PROTECTED
