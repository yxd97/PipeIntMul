`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VKBjk2W5in84Pq0ABcFfKaLGKwtSRAlgGxSgRZrxQ+RjB/Dvz1dfXFFY5twZaGsj
Wpu6EgPRZsGhuPOfdHaKToM4y56xBvKb0x+sEC8anyLft54fImWedihZHLvp+WMi
VPUaaB1CYx0WHiXlwsxvTeotYr39hQrWUwpSvTPFvfJ2XdgFCgFM1edDrrrM5p7e
DUFe/MmJRDkI61K1/6AgsZ7f2Cyt6uyjcJwdkCHfflR2zMx/S8xtGZYJDrzqsUPb
GnP3kzeAwkGxuJ7rxZh+aKwHRfR2jMYHQH6TOxHpjcaISvue0SXivwJ/p4Z1x+U2
J6jX1kq3hfviWPtbMw58zx4+kEAeXogTvGU55Ab/xafIkd8QyAIpVow6MrOqhbw4
rwzL8OuUa6y/OMom4zkT5TL8rwvUJkkXH1VErOiPN+PuCeIPdgMzR0/VGbAZ93Sc
LzZ0SmFAlsdULsmI2LpYYHF5x6xyqUe2e357dyMkpt9Ij+P6KNwbylm69UiOqyxK
yxar5RprcdQbysp9Vs2fFZZ+zmuQ3awNCr3E0yxaZgTjyAKDry7+Q1pkFMxodYq3
NwC5QyVEPrgABFd1Jipn+Ns7FOsMKzBWXJkuPcovRsMCkDKqe96dmf+0NRTHo1ZO
qbkGXhJ+Mss6po/NkXzcyVWwT/V0a2FZsR8ZKs3aPzVojP9UczaOFG7jXzJXjWBB
ZOPeGVxlGy46X7VSZVzbG9Gy/1SqA1oXPHJ/wtFjHtHBFcGX4a4OjF1lJO1fHCda
bmEAoBkWZxbobgDl/bfdDg==
`protect END_PROTECTED
