`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeHqiYrOF2U+QG042bNFaNWDZxLvSQX8nc9x68ID3b6ZLAmyw1JWooZ/DjUYpk6x
YwtIwRNSVxkk6EIYe8dzuzOryeZuGIljHTwap9YN+5sSrmzc68rIQmdb+hdckiSP
W9Z1J8yzYKemRGIQjOqnpbO/IqmYYtZt7oJp1tSlPsiFkzN87dKzoyH+JN8Vak51
4EWCByumFH+Dgt8MRK93KDAujzkcpeRhKbFNCZhfGdzNCfYBpaHkpGNzItdYh1Un
t/LVf1zzlfqVX5FK4zaafdKzVCL+rATaqbZ0E3JuQkoe7nmj+XB91T/EW+/MzHEs
j9Z7ArHRGypbapiWolc/elCDcV9O/4SuH9ESdeEy3Qc=
`protect END_PROTECTED
