`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVXXEyzHDK6bCuFFUDFZ9maR1sunqXolAOQm5xgQsdRsDouY6qrxMJKPo1l2xgY4
8KNl7t9Gu7AQwufwkQRgWYcM88aNwmqITw43lQPSqqRWfFqEGYxigLBMJqw/Qsk1
DLKuVRTXnDK+0McsgKvXcVDMSCfJcNQ2I3COQeyBcwhLL99tVF607FdePBZOkhVl
ERP7+lKOzyTZTvdAIs/bxRNK4lVVasS+q0W1CyyHhs7aKYt6H4n34z3/JblTUDGh
dylBTRgQgZvW6l9qK3SUH+hUjP3XpZHS07e2LSeYNetvOBCU3RR8479Tcyjdw9Am
VDw8LwGKgaEWk1LRD7sKowe8NQv0Kc2o2NEPDNIWaos=
`protect END_PROTECTED
