`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wYspZF6QKEKIf+6fXlFk5nXaQsW4DM+6w6GPYdqtHM88OlosnKmEqvgrzl5hwZU0
mSKRwfLY8c8cTu/ZOyYIulcOX2WPalVtaoC1yLmAJKN7qfouqZcyru5WwEAcU2Z7
uY0vFhghaXjIj6IJOP8mHTNSvORiPilN9PcPVmVcNyVC4AwRupmD+GAQgEYQZTb3
OehUQIexnodYui1gWB+lXwC7wnBq9+qudYQvrC4fBi39+vX4xPneOr5Rsem5ZU5i
WZO/CpXU+YVh5EEHM0H/05rs60a9097zmk19fuwMOcjlBrVgLZJDS7F+pWD8VP7e
QfWOrzMAQANZ8CyDuA7Ymd0ON8464Z3jXforSjurF88m8RFa4vx2JK0m2+Bpx2OD
tuqH1CLbLyDSzAM2/CgepJaGi3J63uDjFY0wIrORrb3fSLV2X+Z7LdrzGYB5iUtA
cE+uSK5GpA2fQ7IgS1XRvzLh5aAox2yUrbnMzTa8PthwwScGAfzG2CEnVtcXPftR
r8MRquVWLsU7oeepc+Yv/w77qyWKqvxDsdDxnEOL+s6FXpcFNR0v7Ao4/VsPUYTD
YSUFsh8o4b7QctplOBtrdeV0xXO3I+D6CLNW8xGuiA05K4vqrnO5y19b6zcoCwGu
GR8apx+WQ1wW9Nl6OY0ddUUf/BNp4+3AWtNx5LSGmRdNh1QP2eT2MR9vLu+gfv8m
yHdZR0oEQO3oikBY7UQKHCnaT8oLsJlLxp20qFRz7i0=
`protect END_PROTECTED
