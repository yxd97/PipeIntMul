`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8T30MxtodN5DpFIJoPMWi4xktpvqxGiLXZK9HMjafeP4o7USdrh3fnolNkRXNibF
9e+vqtJ8DRKH+jrend0Iory11xbmoO6yQ83GgZJGFw06Kdrdqa0aEyZ3B9TvcPsF
skcNy662iLaWhOEfd0dkfQ3h4mBuSP/ovth836knCKx8yREmiPeI6/hcjIgUaocp
tYW0yVLgy0AJmd2gqC8puIURhLGf5/TcsQHtu6hzzwkeC7WMB/cpp+GmWgyFsC4i
dcW3lYdk8TWI7NUb373ghY9DcL+lI/LurfjoGTrWBzTh2utgoDeSeWEz1q0Q0XBS
cDICrp/TrbY0+8mBAwx3MfpfH8yRb4PRN/RsEc0zEUTgkxvlwC+qg0FRtwoUnyBp
3hle07ROoyJp79gIRcPY05uXTfXeO8XeKhyxbNbY85jDEy4AuS1PLhIpjSB06PVu
WlaymqzQ0Jz558JMFOHSmlAMjSUvh+3KlpRXWVsrJUk+UkvQuvJRU4An+G24LdIA
0uknqSGLG6ggtTh+KL+9bhuw/OjjJ5SHbJc8TPQW4bv4lP+1ZuVjTuvfteU096Aq
EYdIJuJBXSMfaC8HRsavS/q0NPcfL2YjalhqteYbOfHN+EJyfkW1ZU3MMcJaSOmF
wIyHVUjsWQOD0i3MZitV6SPsw2LjpV94JErhBhLUcooU5G+GWzAA+wyPERi0u26P
HjrHIXbaTq9/JecJx2PWd230CFke3xxiejPIlAng5kNelmZWiLDCaLZTIcPzW9I2
AttC7SYZ6ENOj9YSpFipQjz5W9QdImQl/NfwH2JOdUvcJlNWILPqGedGIi0csvII
LVwYIzYEn25TsM7DqUsLsTC3JFLwgDh1IfIqGqyEgMr+4N3qvxIhF8iaj27lUT2u
zHAQlFtgjddfDigig/e50hWndNhNmBRqDICsRsq/9rSrbC0th0eEbDAxYrsvpMmc
oPvXhTHOHAhBeUaoHa0eUaJGEIAuRLxqVUeHBKDGtXdpdFKA93MD0W506Nfvq2Tq
U8VpqepcGmxOpdaSXbtkW5ytirkAVq0GRUqNcJNTdJozgQM/5X13YDKmJ1+E/v1b
VhcBEu7A83ZsfRqGwqUxGhvhTbVb4zbILTKlGZ4vgo6VhEF2q3izsCsZ7JG/P6mx
56IqI8IpkBuNdWuoWTvOD16e310jexOmHCGEHR1qhC0M8RashPUPV3o2Lk8/9Wa/
9K7F0rKPUdnV3RsRGpsFuizrLW+eyFFbdSYLjFKP8aF1/2pfxtVtaPcYdcOpFSMl
fHMFwvlOU8WE2WvKVefhr7pSwEa6CCvui+uqbUrtDpSywgo8as7F43vuEGggA1y0
/6Xpy1P+ILSnkOb1iBdErdx8dQHpt7AjNwTfQ6GJJPMGTO0mzaNYAWlRV1lV0eeN
y4WgqtPfGCr6zWQmMXx0JhbTGeHmh2a2OnA4hkLrDQt81s3H2PsZMWo82p1IyKcF
uFqK5e01MysDrrTil/dQoG7E7OEGvFK5A8eB17Ds3OdYPYIta02Ive6HiAsedFio
cLiCHIG8oQ8/wHNqN77NFcE/gJ98EDr1Q7n4K4hyf9pRNwEihijyjufIdLyTZCYV
fgilF9FHgEDXWg4JH1pSUxnoM7kWdlljWPJdI2vH68yLoHhQBhlRTxVkNsloLvPN
9jQ1rx656/epFzxA6WFaaSu8/obe/Ba0A3FmIXMeo4kETEAeA6USaU7mSz39ZYXr
Fxda7xX/Cz2K/IIlUSg5SEHnd5WQExnxrHCbLyeo236lWKFik7359A0lemzZJQll
kNy/hwdYsRycL2kejMks5GMxHksVNGnSQ8nKE9oszmfMcbBX0BQzakrkG6P4B3O2
NswxyYuuO/Ua0YXiXVarJLwUXKspoTRmx5IO6dF44tUaaRPepLjnxPK6SydTwF0o
EZV2X3/wlbKosGbqzkGi9mzLBCH9wx7fPEeq5TsG2oe9D8B8+aTH/J90b52UR4rl
uvHb4U9oWUKwuIgBmq3F5fc4mHvb3A0AtN0zBjul598jPah8LzZu3EVLQWL+a/yh
/b3NECvgrx67NcsfR+0Mtu4xDBLKtapmwIl/6YFVj82ImxP6eRivtvKJOprYK328
RG5o0SqSY8nu+fHjkxfIvCxuZ9zFiL6Q6jAVKheY56vFZ36iaH6XWrVslJQ8hMCG
ySrq4PvN0Ibxntb9nt3PY2mFIQ4HE2b0Nnm7WfkSVb1q07vtJB1Jtabq8dZMR1GY
5jgvlJtKdT9fgxF7hrPuIxBuOpsZlf6U9KvwiS8KlMyZdofVOKoxSOb8REe4tSRy
TM033dc6r7fM/+6HFPFogM4s+a4yJ6erL5FtkhAFdD/aoRWHAWLK7eFGu45fvPEg
JP8aGX6hYh7FnvO3Md5F3Gv5/mZVhqwtL2tg5noYvkeyUuSwBz17QylloDYxUrUq
o3Ovldjb1fIC1p/zVCursMtJ3qNhec1bk8gecfZjCr7oLcaNX9+ahe2YTAxCwvT1
pAhLx3IKnza6N55k1jxs8jVk9MHxpmDGnS9tycybS4Y5SV88EeCcXoQR5ZNoqUiI
GsXOiKhrZeEFUjwCYQq3PmjWvjh9qEp5o1Qzgh0/G1jeYSidQoSVr83nD9tgIabZ
MwM1JqxzvqaH3S53UOKCN091EZ8KOaGIBlrHj9+2vUT98Bsjatb4yVikdHPcHUEm
7KmdZLjKqYpNJWb0JQHwTc8iNrwuiPyTno+PKOerf16XccdyOy1QxsiDxkTjnFq0
520PfeGLxIH2/2fy86lquzejmTqlzqVEaA/WUn89xoN1o3oVNeuVeIRNqBI92YCG
R+1VFHuARUgcZs/GcCpvKoYh7513ju9jeLqi2509s9LuZe32FKyXGq4sagUf5Oy0
Hi+NjsvCEvX/lbIrdOXFH6j1+iZx89v55T/Jfmu45IENhjACUtHS6724Vb4hZHnP
6seFPFHuAOxJrQIhkB7wNYAB4c/+zKtONdw/9/cPDnqV+bcFNadWad9seERpY0w8
ODdf8yj2rjHBHuOaRJkNqu16L3xyv1bq1v7oB/ViDGsaP2tQ2RmeijtRRHObh4Xd
yXGJ4AnzOmGKIPDmGqj0G8ugkViPHsm0QLmpE3Nna+cbC9/Dnn46rCysqbtippoR
gBWJW+/bmqsPIvt6R4bL7K/h+opIndqGJMXRhqOhKdThaoBn2+syRnUVu85PZxBr
LEh1ByDGgS/GpaJvWElGUnUu5ebnCPzGUPCShHR14dd9IC7IB1SRROhmiKBFU34y
Fe9NrxTMSjjebZoDxZ0hOzDTKI/DJNDt/byOk3P16wRndRoWE+1kX+vCH68ZYDhz
j0MkJYSLgMlVRHixfsuWk6YBPzNAi0JfpYNFdhTbSk1nEke1AicseXR6MhtGHWcJ
viQlQDsNyqrmRYwVfs7d1ULXr+z7wUA+nIE8Pbl49TrCmE2QxaeNXvH4bVfEpMrK
z2xqiFZYV0zREKIRRt+JSUu3vRfrgLeZb+mvZiBjNDYQkQt9Fx+SnfNoVpXoHywq
7N21wU3FfyNW3Qcnmar+VaXz1y9ohlNMaghoI8wehPlDZJsFV1rmCrPcdEsrdBKQ
yLRbKFRyJMcibW17/lQBcmbyFI6jGrPUME0P9d4iY35ITeY9kCwsuXr0xYSkLfdM
CFBlUADsqlljb3R36gJFFiW/n6Aoa5fCVfP6L9PaLNnCAcs4fPyDS74CuZnWwGi2
lKBYkw7b4+YzTa+dZ+3zbwfCTYUlPUKh/QqHHYhUNMesJL6WrJj9nvHkkrK6ogpJ
n1sf6wuAnY04GpxNjiWtmwFuyu1WaPs3WOMxLTYIUW0uTyDA/1Pcp7XZlcsuN8T1
ODMUbC3DAxS8KWFqbl+xtibDWyA7jbxhxSThPehoWijqdhNirzvSBABF8+dipDRk
Pz3Din1BxaN0lItDCkrx4FhaYgSy1Vd87LOEzE15LWSJa+36jQdmta+LqMP4tEBP
4Kac6S42pm0HHM6KLOOyLYgiERkAjV9R3FEnGmWPmevdUPFdOAT/UQfyIYSQ5OJO
tsotpyy7B95CGhg9nMZyDEuFsDHwqgzC7lhguPXj9m4p7yocuYYudrMt1XiLqMqw
ipgizvTUaCrRjHoPoKpFP7YNXRmmlWmXjRMwMBtWGZa2Aoe/ZP9BFRmovpw2K9qN
SlGpoPPFPoqFoHQVbK2ulq8ga+XsRGUDIsErRghFtoicZygu/+K4KCePukCwKpbf
tes8t6rMfSNNW9Gv8z9RRnXyPH/lpvifQdC1ixKAI5nz/1I1mBofLLKGoVWVPZwk
cEKsFg6nLCPINPa/OP39ceXYblzwokTgjb+OZWzrY6C/+GQn7NwI/H7XeDMC+NLm
Sj6L/enyHqELZNAKuYcNwOjrzq3KQpoozS4CR7IeMttR1mcc7kmUN6MxmoeIbsb7
ld29QxHR8Eme3Q6pFYH1ZGJ8jebZGHihuX+ZyoyxJVGmCIiALn0rTyB+GunZX1aL
eLfrhRWeS/BXnsZFMah1LC7C/eVUd/cOByDooN4GWbvejzC1zPOcihtnP+ikvgfz
t4bA2sE5ZKpaqRSuOJ8J5WB48FsfGAf7PaOyI7VWP1pvVgw5vCmq7AdFKLg5yivE
MRn/WGK2slMGJHamMiek8u4Q6SyRaz8TbUWtcQZJz/QhOhOlnfrMP1RmWex0ri97
5IoWRPvoK8PpHcXnCNrUKkpIoRe0t6mK8eK2Jo+YP+CyvN9Q7gulNaUCC24XzpxD
Jw9BS9Xk/CHR1crBcvkF0q2Scxu/ui7tQZGQJ6FHcyeWcyeAFZTJG8XCCg0yuPWv
XSIjK6rPMi2eajo16iCG78W91XYic7YB/lf9UVpUCKrRlA3jmDMjwfeQRdWE0GiV
Mo2Dt2Q1nEYWANtSTFmkJphyvj8Etx+QlsxHEtECIR0MCqUeEA27bIay1OS7ds+c
5fITqPBYK6y+f6OFybG1ZbBd9oUqX8Q/H00KmxzGVDTedHxBm1iSjjsIabd0Md+T
DKLfqqUQT92iWxlkrDVm573xUiKgMMdUmNCfdB3/R2DLpACEBTe2NUgMwST+K4e5
UZ0FzSBeHadvasglnqJrAFWMMfNFT6EAiyVFtz4BS72mpEGYVO+h8qZH2Np82TSY
5a7xWCNkj0sXFFE58ZaTzZ1xxwsVaFIbKv+vQM0kQeb3VgeZNnY3jLBMUb2eaa9n
KxV1mvJl6KPofQ1z1t1GU3vbN9X4P5QwD1Nvicp3yGma+qkpL72pfL03wAikcVRd
bqk/cqAUTIA0fyx592mYt1JKqamOUiK/nwZ9Gb2ooW1ymSpAPd+4QgshhirxURmT
9VP5ES2vEP0u9ElCDOoFJonXgGcB9i5BDxCcsnS3I4vWrNPpezJ3THzbxqtaEaQJ
V4c3vR84UOxSyC494VuZTs6wfjJ/GyhdBLICCO/tPdngFRGWQOsdyhxuB4/qrgBA
QFr0pVzdSpq1F0BhHokllzDSZp5GIRKBT/7kkho8ETKRmdGNllIqwzKfARjMeYih
CMpyfdQPdqmBV+CdedMrBZjMClVBGcwXGkPyBpMcu/VdrieY2ayCfKUb47jXbo2t
L50PQHEUA1pUbdSzhQN3LuXmMyyAQQqNeTQVvrWrK8R0SmaTJbXD/WhV0oCXzO8x
nh45wlifVbW9zuPAdf8uB7S8IU/nO42SqzucvTHHHYFoQX+MuOml9zZGLXXbL/PV
lDtW4thU4KDHXgAq9jtrJ+SYD2zDyVg7nDNz5l3nj8Qu5YJtbF+saHw3zDllgtD2
ELd2NBtcXyl1swf2hGuY+VUFqUF44FddL6+DD/jCaL/vS8kJdj+mqdAmkMvI6+Hz
IGv+ha1L9bvbBCHziFiBPfp48SPgeUfWFMDcjxf7eBqUds739bslj2EYPX1VTbi/
8LgAdwX9mlt290oLIJZmdu6UY3VM5DrlK++S34FKWzf1wutw1ZSdXxamKQ5Mfy0w
UwhOks7hVBSF9lUHvRW+DTONaCH4nVrBLzJ5llV1LE0KZNEebY8VsE7hMheN+YuC
WaZGj/1sr6URQXe1ysRwv8Xpl0+bo7QyxcsX857K2+rW9RMXuRwmWNhkLL742GZF
ZyUJFUxc6B4P2earRJZ0Lq1loLqs10Z2J0e0dnB6SxePS5t0CIKr/opJNrw818iR
QmLbQjh8LElRMB8iliE0pQI8LyaZtgQ+M+AjfbN7CQ/JxzPQH41BsrOrHLdMoiFR
mdYsRwnHXUTGh4CsP3LJnQM6TPUAPqXBa9oF7fPVJPZLGnDV+PunDOwlYLJzEgwT
fCDC9kub539Snesu+meP6IubszA/BnuIrb/RrJ2bp2sZ6CKbExEX4Kjqt+IFHT96
wEEkolznVBtCBiP/aQX1RCBBteQEm62YZG5ElfAtm32W8dvvzEfzPVNcePvaqomR
Te9oYRLgslJkG51mvv2WpczeoNYA2UT/Wiojs5bt3udU8lsFEEPw/OfoUXxdHVBb
x1P8x9a3yWUKI1WpAAbzDxerOTIpRWZgjKKMbPWccGT7WqKibhF+O5uPQtk+fynr
7h184mlfDAVibogru0c/WUfwVL+dERTQmomv/yjXRr8kn0mk65EPw6tnPSD47P9/
KMLtkILubfEg5Dz3TZo8J1YPxrNikjQEx8yrLN/9qx+9GivQTbJMC06ZacB9mecq
B8Y0UFdWPN8dZQky/0+aWFf/Hq2ohNaksKhIkcVLkqwHn0EJ6pQXZklRP+5SieLD
d34AWMOhARPtcF2K3BK6fz1Vn8tSiqqm3jKpTruHIGSByKxn2MrhDhoQYCWYojNl
/0P13vtMSA8taLjX/Fvg2jJMQv3tAblFNsG/aXgePFTRLkDZZ3jgNcFaUXpao9f+
X4BM8BjamG/RH+CLuDMQJkLTJJWLA8CgPuyozINkEQ++dhSCSGBrfsnw6ElVMHZV
k/W02N71UwifyNuc1j5GGr8pg3ciryoSDEcetD+pVM3fL+4l8lTdebnO6JA9fyBN
C/J4swS9SFGKbi9KyKGk8E22FQxvvF2Z9ATCxT7zkc1db62sCjjaWtlqmAjINb2i
JqKdkvmFpz3palFimoZCAnGih25X+kJPUvpJxYnPeXiVrGR2qDzDZxiui5ctiPtA
ZdmqB8Fo3XNbzysaw0M8KaW7ia2wf0q0oT5rNXciDd6wAjyP/3FuvTgYmMdhy+MT
87WQ1cOkn/Us9BVEwGIWUf3c5Pr6ZyQKLAc/0o7+gbosuSdpY0WdnVQo53hSa+ka
WXMvfclbPSZCSSqi2VEIa0svLYwao41v35W7SUQcxJq450/DEKgzdhPFxZmqwOXW
KxfdOnMc4HnmsDqO+FhZDJL6yngXRkqdYH/bTOd3kgFca3CdPFQ4I6tBPPoSG/Au
Ymko7RLap2ZCsV8eOnbAdYkU3bGmK2zXPYYeT9/FVK7n9rX3611Oda+fpoy+uTjy
2Cnnt5ttM8Jr1YVwH1W18OeAzt9b72OPQQU1MOdyff7xZ4VFkAtW9q65R6g7V5F0
vbEkevYQb7ciWeFZkTeq2xiIAAc6p9Zoufw/rfTyHX+lniOjMWg1O6XQLV6TUwIa
Q2QWyvbE2+wUxyIvU3DoJhrcq9MLEyF1dD6ZUithDkgVWbK0Wyy5wbpoB+8mOdj7
Es22ZA/ssNJZC8lh3PQDKqH8ZsSRWh+JBTqM+eaGk3tPhRWadong/HgFrVJ4ZonR
Jk3SBCq83SMBUW9dPYP/JjaGrNdA3G00K3CdpJlvdy+satWJuFJeayW1LhpB1bZG
GrTWcXGLAhPmyT8wYaXlwR8pIh998BTzhMqHIp6qiA4PXgW9d8tDNBZAkt3VaMgJ
ZBv1/f4HlDW0ITdcmejuI7fE+GPrHnmU+fN16yqC1oumWgFLOo9RXoq4oBz2EhTU
OLKGA8RAwq/tBN78hbQsFieP+TQNWbE2oe+dDr7deVCE61hJANDgrbKS3FaWMnie
qskqQuSjKuTy7xN1KPbby67opYkTBsYa5l0U4RTCR4uIAX3YnDjYnEUQgyF30B2I
Dt36iWgWf9d3xU4eZfo8vRPJenX8SgXfMB4aosfL4qs+Dk5iEDwRNuYb+/wkX9to
w9aqA1+pG0P1IoPXc8wHSlFMl58mt0T/qmstwzy+WcuGzAV0ZnUbbxI+LhISmaXp
vvFpDmpchMpIe4nrsF7RsVQFV6RAiMEf9XTQcgXA4tmp3Sz05Lfof/0BHDitv0d3
p5T8CFJKZa6+JO6r5iHm9S3dwG998hsBocK4wgOmMEHQeh/AO79/ST5xg46QNCpk
PtZk1XUBhQC8POo/WYB15ejy/KPRcNHTdO7KWpMAUGk511CEMMNoXRFpq5YFpXEi
emBHiS4gW0s1BOyNNn0iDs2Hf0omJ7bPb087XZGl3KIhDxNvPUUskC+68KZxcSX9
MjTs8bG+ciR+tfQj1SCI2zf5GHTGkrCRooKKjlzEt9iZyHw81slisMdnZnb9cskI
Ve6pZI1+7fX4uL5sZcQtSVR6DiToaucNPY9HOZL2ChoImbOSJYbNA5kW24Tg3WVS
`protect END_PROTECTED
