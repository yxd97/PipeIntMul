`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0/sqon3efwLpwdnxNEB+lSYvJraJ8uXoMDMcGfpot+dP8gwxf5B6i6y2gG/N93hI
cyrY+M90KbTmEL9SQpG8v0zY2qrcJwn3bB/ElC8zi3csxHHR7VCqtVRAwLyKNAye
w/gD0iIUN+1NOkIwMb6+j48npu4JcbFgMqHSQ3vqNo354J81VDuhoIm0pfCvT/1v
ntnc6/eLZsSDbQ6addN9LWNfdda4lBaFciuJo/XvDgn/IEGBNRcUAHKH3MKvkCqF
B/Ns21MmUcXNIXrRni30oGQ+Xc5wwL0PGEsJBlKAseDKcp4ttViluqdu6F6CtNnv
Iks6IC7GLnEhaYqEBp3bpqLbqZILFKQQbuQcaXdrJOIimaYrGJtksa0Fv1537Tq6
+upqmaIaMS/xasfrBOmLPhSba3Hw7b2Xo2QwBEE5asc+Ty8qBnmgGcxCYi6ypDlL
lc49eXGKMfWEU2fm4Pno11YNMtXAyZqnzoMxBxdwhRLIs4WLzOzZWTMNAENRriAL
rn3m8vWbaEe5hbthKCiGKIo/ebKJ0qJoKk5rINFoo9n7AbRr/QbrxIWUbpJtPSNz
qmWwPMpJIUoz1LPsFTLqJIAvL40ltpSKOM1ENkUKWQQQnTXzhEVpFSpy5Jj0v6PG
ljh+Pe2KIGYxBSBW4j0GRxWVqtdkxCCbwVIfgZDX7BJVFFUREnVCa+IZKdE3CxSi
s4ah15i30j90CXYL747wrlS+QhJC+oRL9Fatbji5KQT3Qr+VhflwracmUeFWTVod
BotvrRir4fyV7yfErNpKsL2txuXZJSd03gb6FK/u16AIgsa7HT8Yz7aWFdVWuu1e
eWr7JPigJcE31BzIh4U2zdUpR3RF/smCF1bybhcH7f0uboANxTmLqGsOy0YiAHIW
SBORO4zUs3PMIS1yFPitzsNCPYP0ZFBmF/1ossNs0iRDwxIxCmTmIgqqrPn5jcAg
5Frp6wqH841OWDLO8V4OgA==
`protect END_PROTECTED
