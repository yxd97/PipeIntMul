`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+fSJsY/lwsfqopFUyCqsVKGGDNrWDIffGpOv1hX70n/qK0FHkSYKE039upa2/+Q
f62Gh9HaRDSePPKFfj7knjcud9lVTX8IjQv1CTpEVVQevPrD70PBJqb0bJEXW+Vr
D21b+FT5kJTQFGe6rufIpWWWHe/w3/AcFFZ7wjha2aiFqtfz8wtEWmGQm7v8yqkg
C85bzha2zmfinZzSMOgHrlnmetZGwL7fSHvyRHvt72My1v2x67SAIZk8F5ON3aSr
cKcjGVKP0Y9YoUEFwcM7DoLYn3olFEYN3e8h0NyKzTfG6zBgEWsE4a4mhOb1d/if
FS5c/hzOWBuGOeVfydA4sJefYmjFn9BoEszLFJlTuvXAWA4fTyjrbhPSgTG1KFYa
PG7Tqg/my80wPTxvI9OdYw==
`protect END_PROTECTED
