`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KdLhOj1EpoNMhrv/XWK4a5Qq5jpUCkS2RKnX8np2eJBebl30aERfoCOWzkDMYdSE
Hm2v2JKbaxGOrewl4NWL2zNpR67v8JDamKEqAKpqOQMtirOjrpGnMdOuUA8GPe5J
Ffo99tLV6xXmhYk01qeuuG8qtNqp5qa5o22D0dD0AZYZH61J0G3UCixVqlcipZuU
Uy8P6W/89OAwXqZxfYDGyXJerFZoWPtL1xX/U/x2wsrDw9rdz5Rbq/YgcF7U2cO6
tOAh7aN8TL65ynou+IUIs7XI2AEB1JaiEIKLRP2VMCeJQDU0H+2XoKO7zsUWbfwh
67+KaGnbYVDyLJHmWAiLhPrTfaNXJSxEui+hY9vje1amY8cE8MSMm9iJN3/q5q7x
HdXamAsmCqxF6ymVtjr2RZieEml2qEJsBSpTy5ZtXQZPKrG1LiEpIxHagEjBK7fL
Ubj0EvS8lUw+33ahP7cwdCNHyniqQ3hm4LnAEX1aAjynJiDqv13luaxvSXNrZaJ9
PsMAa8uSckR2Nn1DsUdYh6pcbWzcKyvGQLZyylxUCcLoJFEiqaL97s6yBsj23u0C
ExH+w+RUpg/yrxNF4sYSN/ISekjLGA7Ok2Op/RFoRhUPFGZY6FltW9TyWrPYhmYJ
uUvyxMcJtv6LTxgF4nBH+Q==
`protect END_PROTECTED
