`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIafNPB8Qe6Bx2kOdmkcxXW5RIEQalhxPtn7VLEzgFpoSdmkWEmLnGreBZqGluJj
sx3CHTvpjfQvBgc/D2w5LO+Pg+XerDoDHgxQK5x33MqFi14EUL/a5w20IfkwHcKR
M5EwPo23+j31eoCw7VscKKPBwFxhQHs6zqwvuv1zJJSfVg2rVzLyGT0Ywi3xT654
Rwusy47xf5VpBh7VC33pBz4H49GwHdXdLtO0Op5Hxx3EjZNh6SN4cDI84FBgAFsu
LlBS/dZd72Bcq2YkcdiiD1CkxysGPHpC5yR50WoXsF6Q6PlsOMYXskeB72IoNHr4
oRuM4WYefRwQdjRLwJx2wzH/TdlnkgSrhustehYtNVIzYX//KdOi1u4QNSLOfTpK
G0lIHX6oONrCpSYmu8KUn/m3XQHStYylqGcuJuUpz6zgvpuKsF/CONhC9njAgMFt
Eazooi1qIpPs0t85la7PZpDwVGaDCy1U61xc14wvRedt5uRyfiNawrvZSlBm4fvN
E9iifSXFu9miwWa6T0ZqtOubxZZqmj4RcWpm9/kUKCFsIUSLvlxKWMdIBVUAHJXF
a78c33vKR2GEYJwh2JgKO/VuwBT2INge6VQ4IASmDX/iHJuTiK8XNUXGAAbkRT9Z
RqVn/ngRf0Wlwr8VdK9rp0WsetOSE2rITMVt/x/JhEPoyimyaZWsSIfjLH2QUblo
4Sy1ecTs2KnyDBXQvmMcuVCHrD/BZlCbzBQDih0bFDWbW6LAsA/Lgw0ujLhtejRF
oPuh4hKeLuRa313gVQGkScbJkQNTA9dzWYyJEfo8wkwpBFsLzoHQs4dezjrqFn/5
8Na/FLaAj0Gu7dMaJdMScapN/GlefAPlSJUjmi5vpQBmK+JHSS8yRLaiwGehrXCQ
mvLMvhhxLrjC6CcUQRt4kkcBOe9/dTPwcHp5Kh8M5Hh9fPFoNbBOc5why+5e7JZk
zx3PR0weYa6QulJXsp6txI+u7C9IHLbgfrQfNPAON/9UeQ0QJIgmC1F8qIB4ae9q
Z0JZuTYoQvAPsJ3/pxTrgQWrOwkvoKkJ0sTjLBEy/00cf3Mfp4Dm1t0VxfZFiGYP
UyTlNb4WFmwD0drW2q1nP8HAqWZDnMyLREfUxtLrprOMyDnzqfBhx2ENZtDNx/f9
2eP+8W59Dd/ULa1O0aQ5Ty8wOrIjl4+ghPfCqj7GlxJnFOO6Z/iNfLOkI1rME1oa
SpviIAq7+ljL6WYbmysT+oNycRYxDj21gNm7tK1Cbq9xuwA7I/oO5XCghIytGNta
vus8vaEeZX8cmRJANDmgTVyX/3GQNObZJBBG0BTcYKR2YRKL5Aw6XLo6TOcpkAE0
vKuxzn2JxmbHOBNqC8U96Lc5oe7u/LB4otFiBzw7YTle+wxBXhmu8O/dpqO/+mcj
bX5XR5MZ5UK+1YEBRphO27z1IbUJ7rkxITrwfsRW9P41Tw2jxbzj0d19e6RQRrgV
AdQL+xfes3mUjJ0VR/NEK2Xfk6u8/J3dBoOMP5xtpgm3U5uVs+E8K8PK9CpmqsR2
QTWcjETzafBwIr8ooRJ9SUm2+ZbFHDkKh+831bOKHMR2zIfP6i+yTtQwwWTizXuE
MCJYUnuXAPX/ldsOxij+nbezTDEvydBuK5n5WWxMo/aa7ihgiHh/ftPMkM3gSair
sHTyLm512awynqkaokpFzl0CiIWZB74gK5PIX2pzZRdONsB9iZpnOsW1ZtSRB0ws
o7UQ03EzAF6LxkjUyQwAsswx017uPWT9WrXjn1lusMBgL2DDvczdqalkhPOdVEvG
oCBMmW0hksVOy2h8EM7T4o4dFFVCqxxGBia1V+WgU6EKuYaHNveHs9Llnni+iJp9
Z/K8XCK3DKSvccjkpUfoL7L213U0V1CRJV+X0khNY3dz9hgNJo6e+pgil8fdTIa9
5Qy+wVdkeDyflHdsoGVawC2bYu+5hfcYgDJxTXbQPd7CjoBG7QBTPDkhcUtv+7s0
5o/EdBXrbJHMkEo65YiARAwQaKXaXSPZOMsGP+zzaOFKh7hsIwrgIQJtGJIeWNIk
7rguUM4M42Mt690WE0nso5DVXEes1aKOSYGsnflHq2Mn+Wgyz3iFwoJSJ/aL6FKN
Eao7loc16t+uTMMxKBH+G8J7kwaJ2YfDlgYv2vAb5R5imzYH+1ijchs23wgcgaod
HzkY+knegapI3/dlmXlYj/IfyT/Cdy8/1scSbr3KVWcuzb0FVfbGR7XXBL0+cCZz
rBrYicLiGSUAa7PRN9XP+/T5mzURjEI7zXGL+XQ3P9Q6JsVMtEEMbmmSZuN6JNaV
Pvqz8w7/4Zgj9L81VmIEU07M+pidy0YTn0BbDiyjDkse5Z1JQ5+GtUGJ8uZm4cOW
NI0EtN4tjR7iP6zYpvImmmX2g7h4NctXedjSLwoEns/AaDY0DDUGHl8J7rSJyR2L
9QIxh8getZO4oGHn8NC6u5ZQ53k/aiaxLW5RjfRMTwguw7kFWTITqIsSRE8qA5kv
`protect END_PROTECTED
