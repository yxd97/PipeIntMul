`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hx+M5Ml6nLJ9E0ZXGub2Cj6/iB22teLRUyIcW2OLYVQvYDJeAI0s6iff8pWg1ANi
i1Ctpek4IUsqSKcZJPkDt8ZIw9IaWUe/3uPch91HzZojziZtGotuJRObYABnkhoN
+ZRdVOQfwBQpdEQbq0IQz7/DfqPBYArwS2mMKps19IoUO/oETMcZtGfMcwW+GeZ9
BPqWgWq8zufgBUjqXqPd5+Y+/oBD7K9jMi9/QgSdjswtuSW1eqqIvjkjg7NTMWen
VOrbCk06sPtSSTzobR8QKuOWmn6fXS7L8YciwVWLX6B0yAiw32snLjx9V/gSJe+b
Sa7c6OcN1QAVid11oJXOvGb2Cuc0ZlZ4tylkG511B3CKBo9cR7QFNj90Es2crDi5
vL2anq+dWiSa0UQSrwO+NMgF8sHRpxmwE+rlSmosXdyZh4Sh7OPUnsKlSlwAHZFL
ubJk7jSkoflhYqN87/DB79A/xt+HzI2+rFd3+86PDuVwSclmqGQ/PQ7pT5mx8jLg
JoqqQxDm312uAYQfdinH6v50pwMiBQUsHP0UM+rV7fU+1ZJ6rTys3JFfT7N6MpVc
kL7+nsvtX/kQzlUCC8peiHkByq/C1dlfLPXXlXBwWCsQpxzirbPMhZ5u8D+a/fKn
C6saIbjHBn+QzOv3XZb/hE4xtAGyXMJNouD4Yjn0i73fFdiIF0BMnaT3Ba1UHNOT
heBDUtjNj1ZygrLdSgVjcv/4r4tUoFotAnMoPdWtrpWP8Xbraiw23GZdZI5qHbHu
+VI8Ez5xsOhvXCaqwcDf/XKIr4UjiRpp/88cP3hHFfNimSvcvgVsCtTXjBPx4cia
WRzq2y8EnZjZg6cEWh0A13SyVjnySn/1dWPOG4Z3icsihpkYHQ6jXIH+scMlADVY
h300ZMgZi4+uqvsqwarQkswvh83WQCC3cwhuQZGlvUgqbHypi7utaczXdreeOCOF
pC2tyxAamTFS6j5Lj0MvFCBrKvhR9wfANbStRgMEKpmrALe23KbasUgRP5ZCC7Zs
JOcRy1Ee4am7CLilTy9dKNPbElUl2mMSdtBg3+MhHfMNELdw3KB4sc9lhfoGPVCv
QMrbYs6hR2bB34TScJI3y5HJEbq+PEht6g0YmQMVyWPa3JYSMAWDw+8OSGxsg5jj
A0GPKNFuhBHhY4g2D1iegXnHDOhvSlsTZfuWWeafAl7v+7yD435BhKBBZyIY7Du3
GwRJ/oLNxojl3Al+Rklv/RZy4MgoYIy9B1T1qYQ6ryL4gan/j0pUS/jUdFvxXjBM
q2bM8FNCrRb61gZyVYZW4YVdXCHYLm6WpZq4DJuK9NW+o5jSwidbJR762wjDChJ9
uU6dSP+HO0Ko9pCB8lLA0PmFWKZG9FGpT8sMmJ6pPbRQ20Ws+c+41yZTVyjSQHQK
4YeLGlgt5nV6Z/7rU84gkFFpPXUYBVlU2QCvUmIU6RiF78gv6j61t3xLYjTZVcK7
6V4CzCMTb8H5dVLtIZH/WGmprjrjjDV5GMgLKFR5TJCQZ/pnD/QMCjb6isFoSDKa
9otrsVauxwlCs2/fV8KVCdb7WUzJztOMBeboMgST52Yvz5/w0Tso5Iqw2R1ue+DE
nZ9BAaVxw4OmM0Ni0g+ZhYFc57l8FbMeX6zxDm3Dz9JsWWfHeKi4/QG/wnMXDSZy
J97mfTZ5KAi6kVSMKv63EJa66lZ89QS7f6pGe4ASBkeaWIWzTITZ46dYaRFMmK7+
07tCpRzrD242w5AurYbJId5cI17AgJ2rfV3DQSmFE9LMSOCuqb4/4sSpOq69J/4c
pLUcU/naCdtPLD8flKuqWP0ojUIGbWgts48IYXIYGQbNkfeqlAQf6LHxuVbG1EY2
izXG1p7SSp/KtuY8ANMwxXg5+fEgNywLst6XDI2T1Depb4YQ7SqOBXJL+k/jz148
R8GULw/XxTD/wimECKnWl6ZQ6J6ohHf9sIeTk+juskUNbQ5w32GR9QFy3ysLhNyJ
jwnSKpaS8bG+bmiusp2qo1oeEZjwJEC96de/E+hcytetLI3uPoMxFHxNl6mhTkme
nB126XPPCMOBdIa8JV1UiTc2STZJ0AcLlmKU8SRA7dNgzeuU8HLag5beHAmR6uVW
INrsk8FSa+dqi5MAPPGoVnn+Ct8RgICSfha8zgUaHNr2VjRHkIYIBgZ/bywuPk+g
1W9YcBfA8e7O0XnbjZx4R+/iQmA8YzZofSVbYj1U0tjVqlzUPmrwYQJQ8HxiS+ch
QTmQ/1d5K4qTcVTBuuVVbhLO7+3K5JGt1Ecdb0cVIMTDeElztojAQWhrfUntE6wz
VsdsIgyex3piHb3A4VQo+ic3AsZiqyY3ny8Y4/B6iUdJ4XHS1AaxRyr9b+8hi3ha
wa+2UQdGz4rMi5/mTP87dO2jRXpdQITAHK9ITmlUylozcmk5FzadSxOfK1fanIwU
nqdVDz0FhkIeKPRg99X0QW6ebuhFXa2MtELgqWUlCEPH5M1y2v2eEcaTipxHYUm0
mV+CFGmhv9quwQnan2SUkaIXBK1oi8EAVObZ2KbwpVstIrkUJwO+oICpIEttRfZt
3xUUhtWoTSLmJJ8QcsGlciuQzbA/hpqialPvWjqUmgsLm59QuVYbAOvFxLtpjeds
BS3/h00MTHzBdO8SIej4OUgLQX6JWNUICBykU4TrtFQSEKq0kN1cxwVB5wgUUIeh
tJHujnFAtx5kwxYIKH9glmEXWgTph4WtdBiav9vyoHazr80vzhgvadmxYuUoTUj/
kYaUxG6rOjl02lxY9S3+Oj4BKw0RhofpINVQ7l47Zy4jLjdGddAnL8Rr/+Urn49y
PRxz/wfsS/04V27qdSyfKIDOvY4/90ujEeP9OQU3x8i7Lz6pO8PdUokYvH591o8g
uWjtsWKntFGS8VIvtMDXiH8qfndtT4dU1vRSzA7uegdiIjt+52gIC4T0z8wgTLOQ
WRre5oR5/JyyhIJb/Rr7wtKJeTkwM9KECq3PCezMNQ0j78l50PBt0SXvT/x+2opw
B3x7JE+ee1GOavM4Tt4Ik+Z+/9SgVe5Zb93N7XNFezEQog44jgl7AcNzP6KAFVnr
1f3jkj+CtALGi8IWd1EXal2GyEJTvHn9fyIEh3N2gHxV7NP/TmGlNw2rrCiDYzOg
wcFMUxvpIJumPg2ChG98Jjes1alZdGbobMswJJtMHJVRbthDY6xZQDLOnQTtCTQS
//b8DEJz1EqXMkWZXJu2lEDYxleeMBQ/QBbiM9yJ63QV1JAo/jjYKiyEikhMP4Fb
xiDIowviili46C4VrBsjewloHd7CFy9Q2EjxUP1uVGu/AS0NguY/qnLG58ZL2QMG
ShGXamiHX/u+EHfY3Su3CDFGlFGLbcrwLwbuVEsW2d5OQthlpsNGVwny9lK9YJZC
4XqcSmh2v6pZSMHf5OZF4ANm2X9m9j6htTpAZL9r8rzj8yjrW6FI3Mi3tf8R7o9G
`protect END_PROTECTED
