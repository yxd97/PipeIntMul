`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eRd4O5xqIRFoqedU9+gCGQ1DRfO1+JD7sH9D9LenRsObLiJEf4K7b+BvbY9DLcNR
XzOG1nIyyJn/lKAzY0sA5BwYhxEkXpxiqcdepjG25rnMnu+7hZfEzhLqzJrBayxg
xX1oJzUgNxU5Yc7hJUVtTFgU+RWCdRccnsIr8XM6wlUsEwPm14MnF2lzTS1AFTk3
AjgATNn201JeEj7QB5urhdpUkLYbE9oYJhFAzj8NhEnQYMOjfb0vaGQ0Q/4Ugbjk
5F8rxjigpTXLqZNzN/+rqK3843pYXQPINuAEIw/IDFLJxvJdGjZxhFAkNtJcmeBj
SB3EISgeiBR+rwNkGBkz2SgIFHzFnJVTE+vqkeFyRxfzuaZoGCAuJNLZVCnynmr7
IOZBDLG6Dpn/hxvKcdmUHdWHRU6BUFZXx141vfaoJPhZfc8W5vpCUZk3iapKA2VP
p1IjSmewXV/hQHhjmSrOl59pIeSS1EB12ccwJLGo8irzTsQadh01NgWcl/vN3E4L
/L4dJS0Wmf6K0b6+/Qrenhu7uPbQDAVr2EijVCACG87PXumFpTY3BPte+gebvEMO
8skdM8RYZm8LeRTnJbxIUMR3kREFam6rDLRKd6HwJ58HRVfkLrXh920Vb8gXsrnq
x9eIqYoyMeK9zKA+09vGeMgZTzeAt8h126CupzD3FlhbvlNJ/MbeHk2nTo9p7EFf
j/n/w8A+sXDxx8CBFLEbbwXUXEGiUi+ZWNSdU38PpMuVs+1tLDaQPS4L9TtSBqxZ
fDPqoizUpFJQ1xjJLc2gtxb+zns+I2/GpUoSPHshJeTD2jypWjF+ddF2fQH+OCvo
uJfs+bmyGaCdvzJB5P7QoMvltLDbAKWWN3JT+mfvwIfhH/ElhwZBQXQGAPPaFfe5
rstXwaaLgAEG69MR/PQm4xaFYvUkVOmBRIQjKsyrjiCXs1q5AS0nLYfA5S43zeT5
uQL6Fdocj7zWt+nBloFMmRAdWO+OEtWEG5bcV4Rek6GynHd8UvkiM74QeWUk3Nu1
PAbNjQ3g+YeA++wyomm+QVal3qG6AtgEeOe6l9sFQk5NSRxmbFDGrXZ6m5W6GAsI
FPiIqEQaUUV5s/zfa/6hfNv4jkPZ1gxGLjeNr+V0BD9IYQ606Y4gBr39tLCt20v9
p4wUmN2TydncZO/muZBE+35lISX/ChoC6Dup+8BGa3FpIYnQC7F14UzIhTaWB2uf
1gH5mBYbKoVDDwmp/qqGJqIhyJehkqXkFzJCOmJZIRZtCQCaRxPa/Gm6cWlkW9nJ
pnjei2igamq+VjwAT8bTgqfCF/qFfVQvGNZ0Z5SFB1VntZKJ3Cw4QZUxSV0CjV1W
Vn3HAFWgdKLd28E6nG142T/bgmm4nS5AVybwgrCOKIQpU6ZHEYylMxtu0Z06d7fD
UQmuIQX6Xqa6it11BRNk6BLOyf513KQHpby4GMRIV/p4VTb2RnBntksl0gOnFurQ
nrTs0FhLOgVfqRywKoktHWR4cHUc6RyQ+sKZ8dOuNgMLppIX1MW1FrRNrRHuWdQz
6Wb0+jzbIsHuW7b2TGtCJgi7HOjOVS9p2eRWKi2u62OoWEimgnBaHhv+jEN0g76u
PYbGHzlnR7FZHd4hTM8za9UkLn/jtZXEJGkt57JheGhiZyC9e3r5gI+tsmKoDn1D
vBO0xuIKl7oq0xS+ElE46nU8alZj8ppfquTSLDUJNcF8LJoUMlA4YqI5dDyG1Sa7
ZXht6eQZ4QnIMTH2QPPYodU51UGT61sl/QX1+lCs2bH3Yt0D5yPPLcvotNrrkhdZ
qje4axs8rTW49KLAKiin7K6XyfEq/qXcQZPlUJT08ZoQWc/KjaGtW1tt91diV13s
kn99DLd1pVU7pgOKM2INTz/jqZeilOl8W8VYE9LFN+RalxhDnlX+31H/+eC6rWnu
mBo/lGBPQAe2gW5hn0dDjarLm8poJFhWiXyDoizLc4uYUz6JbKQK8nCa+gklL34v
JsuvFdvCFH8aIM2hQEFsvop2LdzlN+8Sw/wIs+hXr7X/pz63mIuPdEQoJ6epRpE4
jtYap3zidrki8CNc7YWc8NcUPc0XWqO75B3KMuZZ8rEXON/skUMO7Z0p1S+lGrmq
fkK4dmVJGeX02o3LG41LS+EqL20sTSQjv9jtYFtF31DwhrdUjj8hS10qEp5CFuR0
`protect END_PROTECTED
