`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/u+mud2JQapd1AiFn0f72FpELc3iMkVo/Wap2b7tT+ZB86ix0sc2xCslFKswf5nQ
IA73pIUmffuXw363w5oG4P6z/gtMFzG66zm7noFF9h+F4qZHRngJ2OKNgxcb0clG
Bi0nxSaCnBUgC1H4X1EgdPMndKciYpNvFk2NSk59iJgHKPUiAGOowlnNw98+hz64
HezMYl+FSFSoYDrCkaGL/9yk6lUsc4T2V4bqemPcoKB5KWGi+obzIuzRqmyUCcmM
Gyl5klolFg6rjYCBuokDbZ9HkCTVohdWSWwGIw/lXhvZa2k7Eg8pwWCj56RxZBR9
rm6DlgzRmS/I3XNLFmyloPtg9/Zo6NYVd64TrYi5kiHVxHiHwXxG4tFRPXuW4chh
tZy+1gq6Zp7LnbOpdG4y7R9J6vpu1VeAw9+B4GvN3oVz7JhuGn5rDDT/KCpiWRGH
6p1wzv61ZFH1ZsRn66OTq6U3JJEuxMP0/8JtXFvUBzcTdxAd/cMVi7Y8gKNUzYK+
ro1C5h52k0zPVwIzDcmv6jCLO2X9b0InIAxgO5151wRAVrk0hHtUoZ7Elk6YQ4dF
vZJ6Flyl33tydeNS5yXrHUtzIIxbFkm0UJ43g4d8QkLLqHllumZZRk8D526lur4g
7miNaBdJSn84Dx8z//yW8dChct+KoRgYp27CgDY1pQ2SpMn55pF0UY99CZbkmVh6
2F0KYjIWYN69F7pF2P6wsYevqlqMpgQ+VYE/pJyqhtlBAxlSs+iuIOCQZe8JcFdK
EmO2ey4RUJGozzWDaSS/h+UOl875lOTDhWRmTdy2EqO+dtZUcNXszy76CxEw+Ehl
OClX98N0IpRFfdp7MeDcykPvvRNRvqNMT/h5Qo30bNwoxXWzK3xVTSUCnsHDQ1ZE
+fs1PLpEMXqkvRb7G3fCnLce1IaG8ze7NneSCQZmBluHPvvKZ5TVDf7fNhbUtDr1
Tq8nJj5kW/6+tTq6Aky96tFA5Obn/oDPSv6TOKC7XN56yxJDeWg8QY+k5be7swaF
h5+ntSySHFnoGGmKrb2XPgBKv0ybpOKu09E+iZ4UjEwOsfB3oHHP57o45ZHjoZd4
ZRn/yI0MP1gyBjAYXI0X2SarUPhl4Z7VOO0joc3cWsvSjkFKNzlZDKbgyqSL0TBT
9KKQl95EBt6HB4cxnLn+MmRJJRLDXpr5UgrkTK4z8lHwEkFA+JZqOLCiIwVyT+6T
PvmbzgTWlcN7ewbnF2JQmR5xowlxXrkDEAlQ3wwuDPE/dvKZWMahxW2H624kkZj2
muok4PoiKU7c2F2WusuEs98bU837hIdaOyL0JP1BERdFldDa5Zn30jMCZM1h8S2q
rSnfIUnnwV+DJONAlJuW1t+qYCVwxJSgw9vJl+bBezwKIS2hmUvVHidU3Ypmw5LA
2fb5KG4LRZw5tcQDmO+NTF3Q2i6ODhFi4dVlVtpOcpE89ZON7BethceAvZhHAHDe
wxXG3wSPqMLYLt4ModdFoiw+O9qjOqbFsfAYbt5IkVToCRBsatWtSgdQgXlmD64h
nuxi97yRJtREZ3hwfCt601nhnyAbfD4jAQcHBPljp2A/FXV5vGU6gKf5RFqWLnic
o5aQ2quJq7dEvNlz4bZUYWoxJ88efC9rhZsZnVBSQKa6i/OpGdzXxj7b0YN4tZKj
Pmc/buOXOdEN2qU0OjnoGukew/KY0Wi9WtHz+2fANiqM4ToLnTxtNS6cmlNYNPsh
tldNuC0xuHXbEgqj7iR21ooESkfklcEyEkC64XHKuSXY3H9XQIiO1EKwylqV0MRn
hUW3Qftvx21Zgwg0QvWoPEle5ASxhK0qpmsLoujYjkEgwdCGyur6t5lViTG7NCr9
yaLvAiDKKxjDOTteD9Md0huJdJAGvva3kdVvK2/GFS34Ubv295GtRsf1trX7h+1J
ikL4nssCdez6Ka/0weiLzz0H1RGCOnnctdJynnqqWYln76xbv2g1VaqCRf5XcHPm
Fn4eGgmlmzIfkZcGuK9aipF0PeBM6uyZztF6UHNJ3DDkyM9knKp2sMsLmGVxPWMK
si6Rof63Ub/GZVky7Q6c+uP+pw5a8sdvjZ3XwX+gpk5zzt5j1RbDbQqc7V3zDn0e
yfzZeBub57PW3ZW+Wl+QYo/46uOAtzZxJC/1mgts90A4BNkDNe8knuTq0SHEOj3W
hbZbWcaciyN3BYDk1T4VLgYqJ+B9qlKhceQa4OqC+2Et2LNgMTt3cbGa498NIKEL
`protect END_PROTECTED
