`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mnHZlZXcSwjnxln30eCIJdEHlYKFsjoMTpwL4kcPCFrwPF7aT3vkDPbeHw+v1+UV
2cobJ2FAzGLuudyFOQKkG5o22WYtvgIW5g22c1WFTVJDYNJf8Z4mfZV5C9e89kaZ
MRabAgcDY1aXhkeHNY3sP7kBJMcl9iX4BF/NKIGJiTCqXJDpdULXSiq/secvU3sz
mgBw/UosWJsrvHwkKju+p+Xbzr3PTpdZcZlb1+yfBq/Cl4t/Aa8jU5Fnh/3oRRn0
aa2E/xAmEqdHR+hbnw3gO8UIdAWZkMh3DoPmtWjvUxHrmfT5U71Sk1qiVNC3f4KB
lJeT6/x+J8S0XEyAYtwcum7CGfR4/q48pT1cuGU3xFgo5kp1ICMz/pdryaS2Zest
p6avdLUDmsW20PZs5mPq+M8e8mTMZo73js+wBG25GiWFklQKKnzKFd5u+Hi6fPt7
EBD9hwdazLv8/NM4ut3ktWDOfEnrq5OF3Fx0S05AuuuzQ3i/ssXicormGydpqCKa
jbaj1XhWJWY24Asf4gRbAHZ7XxLNKX8Y7LFNR/szYWb0kojsjyl15f+32Hx8S/mP
tq1ytPY+uMGuOxaY1oUrkfHgJmJhm5TU2ISmZd9Z3tt3mnVRYOAIjmiuVCxZH6mY
EmcQDxL/+6NUM6X6ZtC/H7TsB3Yh1/Sgvj1qUV8hA0MmJekl7126hI2DmpBPwQT9
8rw/uix9QFyFNjVMAjVAYSa3e81whCD8BSVl74xsBNvKJuQyR8yZDQw0QGpWYDH7
RJu8TPv+Dkd7438POAukMoV0/OK8ufJ+tpJ/C1Vx8aoH4wm2Mu75MEnt9JKyewY3
L8zZ8J7LJCPSs63oihO+fPs4E7+35NOlSd3w4dUZ4n33crAnU/Jele1Ur+TAIL7Q
q6kw4HKcSfzXCOxoEliTVB6MkTOb2K/AG+nFO1TC2d48VZ4PUzuWX/QLGn4pB55o
`protect END_PROTECTED
