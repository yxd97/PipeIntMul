`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OjLS9ABpBYAAU7k13LEKNC+YfOzbDGtHGiskzK7GzcZRU/l/x8JswtE4BPCqsp1
5wL6LEzKubeFMuJUpvs5Cdj6nMimCv4sdWXM8991yzfmBl2QIOTeoF7Hk/rhxo2F
bBYRVU6olQmSKvwFGw4nyGsk69pHgSRWyKuMEifq1LJd28gRBxyvAygqBtNoGJq9
n7iZXFdGmKDnNal22owHNTbNQODhjoCiHsFDoLOXq+SHiJaxabPUXfs6I/oevLNO
lnJgGYmAucohXdUFaA0TtA==
`protect END_PROTECTED
