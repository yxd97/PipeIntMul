`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
plq6Ndt7d65uEdDrd9lkmHq8cK6k4NF29M79jtJok+v6rZpB7ikGcvMTJCfCVkS9
8iHR2CEKHS1oDbIGHSI2mphhrd17IH/BZ08spgveCV2fHjHAByTBSDSTAmSw8DBM
vixf+9ZHs2j/DoyY2TyKTKSTGk6wUbNkZv6ovuV5Rd/FhUaCpWrpJc/u89DuEVDQ
GtGrQ78HsEAT3zBSwn8k/YHEPxetiUlE2BZ6qPkCIHXtC26qRjP6qjK2lDnakwrH
uoSA1SbT7Q+dC+9zT9o0Kg==
`protect END_PROTECTED
