`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4cdUEjx7K+8Ul94JzqFJ1F7TGSFgGuSuzHsy3dW6cVJMfx/iEG1HQjaDO/EnzI9j
pXUHPCBU5I7rBhzfoe6LwYdOukZdDZaulYtDOVDJUo1uCdSFQaFM8zpW0RDbMaLE
HW+UqNGvXJEd9tui4GlzQcVSMX+5v0hEiRcExG/YBSU7LbugC9K/sYHxalvA09jO
u1kKSLTrZS8O+UKEpNZKFRZJtIk9J2afdaFW73RtCOlW2LQJQmTmURSbb+O0LuMB
2tniqIvGupaXn/cmzsXvHo+CqMN+MrFgbUshTGXAHd+hUpLI2D/BEzbbwC6Qhqsb
+PiOHfyuVH7P+bvkjgJQjQ==
`protect END_PROTECTED
