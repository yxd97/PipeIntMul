`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SzERMfYJn6+OS6wZU7C8IgKU1aeSqql9U1Z0NADU/l1Kl+8vfCAx1ARQoCgHrhpH
HkgiK1EE9SFCJylGE5EjdVka7jQJR2ANt2IY1YgXe07FCKALcmEOCDTpE3cCvNSg
Mc6K7JNjKboC+G9WtpTop2pbBOUr3ZNEvBgvwe3LzCCOKU+vYvKtfOMY2E1o5dKL
cfcU1NDBriAzFRlszdPwn13kBJivG7aq4OHQ6YOWStSm/CmUIFqjcGpRht1CEh82
Y5nLbkViaY35tmWG4XPMlNjPCSPLnRhJka5kLmDvz556AmMp7vyCj4CL5poyVdW3
WM5Xyj9mtj3ws5ZkZ3SwgP1SgML7shvfJK0cevDBbcoXBGOF0pan38AiyIWumNOh
8hpL11cFIvrLCG8g9q0sh/tZ6wUf6yCjtyatIlkLRGyIWrLhE/GVWddtxxI/4Xwn
KZkL6Dc7NXyDyYJuLgmDG9yQk4g98oleQqC5hqsrV93uoIcdDfS5D3j86lFAgsmB
9TT0LUNLACXas1jfBZlFQ3OMG2pW4fcUhb/O9AjJrgh+FUPHEy4xfCqPsmlfm811
tQO/i5kUhi2A0u/TiToTVg==
`protect END_PROTECTED
