`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DpDoIHttfwCyB8kvylALRK7t5cjOsQ1yvzsTMsUwoRmlxVZ9Z86JZ4wNKha/m3mw
Nj3Pyz6CUrbdDYsaPovpmd95iA7j5nee47Gba4QDoHvTpJ49540nEARUfG5uGcST
JoNHp1PgcLYGU8pm0g0VXXcmMrZD2Vsba6Efc6TAzBwUSi20qmV03O86GpePQ5Er
xVu+cvWAQhU1u3SCs5CDG0AI9EnRUfu/MFuW3ogKSbeagDhcUWLdEjSovVU29aJ+
wCpqu2NX92v9yWwBMnHU7jJIQkqBeTVAFQy2LNU38H1nuYYOUPT31/U158ZwlN4r
dKn1hndkkdTh58+ccptdQ2FVhvZr95p+k1aTGozNaLUxm5bai1wohHj7N4l96fNl
iBarVxRGAlkB+B92VYmPmn1Ih5EW6YbjXmCWY4oPAaUL5zyoKHYkQh0jYFkWE48A
ZhP8lYlfa1sZ+HvjLvABZXvHw784PB+nU9dYFas33Xnp/gvluuB5MQ/bbSAXkZDW
qktZQN0phzSDw0XbkMkRVNQHVixKTNTNQvMMUQDYJRVuGctPL88n3vPNr4x+OVJZ
1MFw5iwCYfYa3Q8lwKq5UlUzx8zC6LZfnlfCONPprAzxr2YYw0GYzbZucWvG4rEV
doYov5wb9EC4uQt/roczBg==
`protect END_PROTECTED
