`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0cYGSoyk79v3bKWee7dG/BGOb0J7nK6GoKN52doT651VFHgQnQRJMYrysFlPjHZN
SgP7PZ/dh5qJKhcCQ6H4KNg23MUj//+/2GwoHqRNzEZgxm3NE+r8blZGYDpbF6sb
FyoGWGywABcpQ6goyyp29ebnUweAmvik7enGgvUO3lNRNP+T61Ccz9vizGe2BkHv
L7hNHgzYHmPJak3B1KviTzKcyRZe27bNgSmv1ESvVe9JdAkcCf0XhGX+grG4FwEL
+ToOgWYKfO9jmCOajOmqP1VfZ7xe8I1l9j3CyP2yRjmVCPbTY/JvOnBKpHMW/iFy
GvwTbgqKyss6t2rVs7bMDL1lNfncGHL7eFyyS8KWyl7IiQ8ZiSFnimQerRrVlD6A
hwBmATiGYinrL7N/HXbVT1BNgor8llDBB+B9t+ve3rht2S9HZyxplY2Pk95rZb25
xwZgLZuphIGhwjukGTJcz9TDDualnNMHQRGh6opx93o=
`protect END_PROTECTED
