`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1n6Oog1VJIvVQp/4ECgTbSq+9ghKto8q64iEBF80dbXUMo/PN1bKixYim7Dq0ViZ
7jmNSXqKEMHGQRZymKuxMRK6N+PNx9u8JJp3xMsh5DCb6wRJb+q73Fw/qMaO5KkL
aH902vCiPYSP/0TPJHk3TrOmuVX0qOVGpaq5SAkyVzvNhGAI3a0MdCx3U/PtU5Hp
yf1awWqGdqfeEDcUX2mvWmdhK7jGD+wWBKYoveohYecb8tqXTqxQm7ckeqjEzOx4
ANL0jvdXN0SNnLGyxDD3249R/WlMtgIvu0s+y+4Z4BqqeFPZ5+en4JRZP/0eLthj
IX5nX7xdSLPJpoy2bT717Bf75FcmRFb/YEhBJZrNMKL00c7IsJJCbO+91haAr0Oj
/kwKmSFrZ9w3QC5AJqXlJMdwIqkzVepXWErPYebtJ/m8oNRQhfYlJWdVTos3JUw8
wB/ddzl4RnL+a8D3dXDzlIlcOb9wzQUeYvmIYaK/GrbH1tCUhSjfkI/ETII4u1xZ
yYC8KysNYqp3OrMJqrJ25Dbe4uauqPDSLAMq5GZnke0=
`protect END_PROTECTED
