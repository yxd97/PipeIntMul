`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZL5+8lbmE7VfJ81c6zB0r/otyP4WghoffDNZdnkuwH6OTc5erJeo2xXMj5E1/7LG
y6qrOkMPKc34kSf9SmqgTf4DUFBhrZIs/zO2lFzZyG4sU3sA4TSw5fl/QYvI+HKK
RxjsAu/ilCCqj4wGfFXjpVsbeI5UtwuFelnS//NSLQ0JH3h7AGsI6XbXKOAV4WNz
zZ0vxpttSppzN1v4nxH+A0hs7NxGK276z3WRHREy3n1LEzz+oVjMhIfyKoO7lwow
OpFryfj4ajxeWhM6KiPkxQ==
`protect END_PROTECTED
