`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uns9iSA182awCMIfDys2bWGSp6cVGtfzHDGpju5tZHUYhuQLOcHB3QaWdolMmKHN
8g8qKbiAKtH+suSN/ouXh9mWla/2lyozj6Ua56XAyyA9cn49pGtqNqnh82y9JndG
oL77Qrb4TLn8ILhXMbK6L8AxwuK1gw6mhtSxYJQpN9ZqurbrM75LmsdLOeSuMIjC
q1Rte5k5ndOL9LV1ONQSznaYVXBbxymbQuhbTuyhmvcE67l8F4jDw5a7xLzRiLOW
cCBzHcEOUizELJabio6N6J17FhKi5zw2EZ7Lj5FjWl7tZhM9Gi3b/GGp+3YJIwwX
IRuuXdYX3yrX1PVK962FWz0eufzbTdEi2VB4F2kLS3UBktNXdpMHwtxR24iZQDnK
I3C5+EPzSLMJFEXpVJ5syJ7fy26L80x/hA+APsGGx0k70tPPanKI4LmEyD0p2iXv
/m1fbG6dSUS/oJYBc7UDFPpqgHzonsteh1cHxaLghhgWHe8TMyASh1Yt2wQBYyp+
f5eYiZ09usNG4htrENpwSfE4ppqxKzEsIoQhrzTFAGDNydAqv/bVZvhzo++md/IG
`protect END_PROTECTED
