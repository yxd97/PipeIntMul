`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7A7QNvnxr/i6kbgmwZZkQ6vWeyhj3c9eML/3CznTbIqWbuAzaIOUHk5qNmqXkcU/
o7hm8ygXk4XXnw+ePE2S7hhCfyuJq+Lcqn3ARZQCyrr3ov1RQ43d1muPU0uLIJTA
8pWlwwjzBfQjS023sFmAzjddNoVhatRKJ+4Aa5Qgh6CVl0Q6T9ANLUYm5ETLNYCG
3vD3XM45F+WjqZtETDkKMp6/5zfuUeajiYvHzpup+MlN3IBK56dzlwIPkGGInI2z
ww6qZk9QIuMu6Cb1hByjDVdVC6PeMbaDBm36RNpW+HtC/Rp7x6XHQH5srIukkKqs
3a4cLKUnSnVq6ZG74y1DpIglaygA6eA9t858fTg16xIN6I2ma8UvasW1MTCU95Um
KwImgvwCzldfqbT4lVAgazdst/xU9MA+vOXl3Qsq2W0ou1+s/e3q0yrqSWJ/Ihi1
yBc6fE4kMMQK09I3j8ld1OZfGs5nfw4uWH1ksesGUQLa8sKBT82mDjrdUKP5KR9l
0Z8hOTHgRQIFKBRAEfC3kIy8Cg8/2aRddBD94WffoDcrj88Frc19Ulg4WzsG63DT
chS6YzkszJm3yY4POlQztnnDhk3f1Z5Eaiza5yaMLfWAD9A4vlKIUZ0597d61WBd
`protect END_PROTECTED
