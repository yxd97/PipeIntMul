`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2txTy2ibyqMI9ZAUEP0bymjqH3j7WOPnHexXtRvSVx8HlDoxD+5VDRKBhtYHt+4B
u8kCtC4r4wAi0GFtONfMTvi3ShgjF8swy33OohGs7ffpWzqc4vr8qjnUPoh84pNS
uQNjkBdxGf5cpi2UaYXFOorIn0OJdqBCet0hBpWoYjgDounV8bhC4lAFIWqC1+0U
ZFN9kNgoSuMglQevLdTgk2tuovTVxONMAaI87owqOxnlmGZYi5mmVtvoELHRfmhQ
IOls/+GPdPaWBBok72iVAv5CkXr3YareX5AJsBdgIrD3ENsIPcu4Ocayqtx8nXwQ
44ZedHcTfv7XK7cD1Qn8M56AxaQm8D3V1w0yL/qbABffrnpeBbl4P6PkDSv5n8ev
ENlkHQbxiCOMn4GdqXnCOQ==
`protect END_PROTECTED
