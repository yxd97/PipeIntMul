`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y1qeqLH8EaYmyZcISoftZRBGL8nOuog0Zed5zgVJPAboKmerwnFrhQkVUK8QMsIV
wS5H18hT7UUxZSnyRcqweKWaF14jUix5EkrFPiHA/2GJFpGRw7q7A5NRR2O15kPw
8oXyhkdTxX/a998K11hXqqCvFFD2PmYmAoyV7Y+GyhJXSthxNY4aAy5niq3dPSZj
btEXyOPzBCSZn47MgzxejEfRYnrDr4Qm1mHwimLtYJat2kuwvsg8gChAskBIm+tB
bHa3X5RDwfjlhWJ+p22DbVUArX9XTqXIk+Qn3GBVNbeGSOD9iQTBCZaElQkQ8+pN
6gQTeiu4dqZZA6+wIUd+3w==
`protect END_PROTECTED
