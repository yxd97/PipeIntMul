`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZDOcm9hLejka31vbzZWMgLJdYAzKx2Evb7/P8X2l50Syk4bykFdewZW9SJ+H9SSu
8hZC9YROhUwllzzsKOZdoDvIVdsYBNRzuGroh1hKorbHCYvMFYXKZOH3h0Lg9OMC
Dol34N483SrhHWizGM4tzQ+guWRAQceNtfhIzUOkRkT2rkMYWTB0IoCg3u763+eh
crppHW/qV2wRpDm4VAXUVsa1VRbiFnMrs8eGJFnCpChZMrss0xJJtF75HEUHjNPP
oFOtcWr9n57v8Qu3ZN0vpe2gViLrshDbpl5laoo93dEnDwd62rk4iX3OgHHbvigv
zVQLmei7nJx/jLOcm8On7xFwPBLRj6eHKhUWZ/RvuBrxCe2/I8KbpbWDrz50+KGD
X6ESKYnOCqYeAKMoJVQzrA==
`protect END_PROTECTED
