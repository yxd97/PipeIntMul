`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBAI47ni28+DgeqsPcf0U9DuwXUdeIOfHXdKhnpxB2XWQeXRK+xJAyIaVz+BITd3
7B7jApYb8/Jxx9cyvh70U654/AHBF9p9NA8/xRHSl4llDkc0BBegvquzIix6wikg
3FQT4O81zgjqjG2xc351IRKvC7Qy/+xbtiXgngYOGqAKSExduMgAKEJHmDuBUXEg
RHJOozAXeAAZeExLDICXtyKuyIC+6IZGnN8xguuZSI8v7znTzoONYfDCaFv7Ykkf
CX4L3xgmnA2sbwNL6Gas5w81KAfqr/S3W0qGDHqXBiTZH1pj+UvhmhDIZGUtgcox
MEqnQGLr1ChdsMU22Qg1oP8v1MyhzpPQTrY/PhO8KGJe+GdYVKnTYZmzf/9g6BlJ
R04JKS3Zw3DtWkvmZqivFbZodnzJva05eCrGHxfShGQzGHf2f3jwFP8nsK9wItXU
CA6gAXNW6BlA97ztKUYVly4yrd1xnFT4y1smq0oUPPYVRsdyF6oykeGK+VprVVOj
Xs8iQpribK8564qCPp71CdImwZYkrlplif1RBRLKdfjUlubEX0r8P2ROhvu3iDiP
JGYnTS5xCYNGPxBdEFuCRKdeVMKC81jXeX8FvXHbMWqlFp2+ApjG252jSLib6JQE
pkYO2P850WtLWc+BFeGdMXciqSbUTDA0laF+I0Mh6UrVkohNrYVHjrHCGevcz+N1
JDYaDZQi2G3y+ypMiTE7VsozqRAWucoBljdDMN+T3zOoyeTOnEWNrDYhPhUHIITn
cZ+pWLWGMzn74heasA8nfw==
`protect END_PROTECTED
