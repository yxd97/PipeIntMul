`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yVpHU3lzEOSkTdhjeAaKHAnnG17G50YE1WxH1ccqXpbv5MKY74vjRxgnEH/p8tTJ
pMQNDQbvCSHf+vi0haFsmIKelp1JwYzOaPNOieNR8rKW/k2sKTG127tJlYttwGby
kI5ChdG2pc6r6C8XxClo5w2OPPB0vjFPe9SnM6hwmB4sQOBorAp37Lnf8Kug8LYy
qR7T8Uv4Ae9uKGgApovMXBGlCRN//XDFsnTGygfVm6R9ZOy5WydzGWNYjBvOBi2r
oy/z6z+6xqCnisrN3NJ3sOf5ITHysNMq8XibBccLhtAGRf5vUAkRKOUcEuTtYAjr
kDBEBgkcVgB1ZCD1AwRgxIDdY2P3hPbisjnCkck6iPKXVfJ582ua1q9u1Focek3y
halMKqOel+zw1Ct1HFkKlR9i11nai5aCR79JPQl88cp4Mgyl+owKM53COkaJJH7v
sTpzRdYfMzw+aeRn+AEah+Ja/iwdLu2Ec5anv+Xb3LU=
`protect END_PROTECTED
