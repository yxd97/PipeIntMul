`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mlV9fUdMDmO0a84sM5y9sSVsYBucytRRiRmaaPqAiXzm3PZpkNWewEYyTkEdcVIK
r7b/cyyAzjCJPcL10YZqUvTjONvu6JHl4rxVMRj5ODo3K8J7T5pnN3cxdH5kHp/x
mPk4AgYPeygDx3AnYUuQ2jpuxGibLCJadGdksynX8DGzcgbirEVMgu/vnU8fUMQd
krBV5Bmq1nHmkn9J9+I9E3ueLY2CvvjqhhIEZPnWXXgTnriuEO1OYCK7aOL+W6lO
`protect END_PROTECTED
