`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xt2o9jmEIkZnUmmc8GQGxugcBhXvpIKybKHm/0aHKEekk1Ih9TEm7fkOVw8hrLh
Ookd7+qIXBMKCwo9nbFXSXMSnT3/npftEzVANPx+eTYvyKwcs05/e8N8HSTeZ2xP
B5w3LMPVGxlQMg8gd6mN+56f4NSApyA2U+YlslH8mey23/mwn8VRfsf6fNhICGY1
KuP2KaxV3ZPyzbxB7W9h0EXKSvBMmOpL4YNHVSW98EyJv1IfeOOZDf67cGYZrMqZ
e6Y5uHUBIzdNONn0lk+zcEpwuih9lJv7ABAq43y5OxWVUyIDO2gMrP2lQA53xatP
eQ2Q1c5PPaiFVvrHm3OZ6119rSZPk/kVsxNJvvKh6Iwzxpq+Xogu75pKqmNROTD/
jM912DH/T17GjOH/REsAoQ==
`protect END_PROTECTED
