`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yVRUB3D8P868WcCZNGFifxZx4wPhtYugQLAOh3ZKk6oi4sCVh/w9eUpkP/dcIC8
5VK0dTMWhvy+6pRRU8sh76H2c8rNez3bRwmUlZPrVOJmV2T/rIj2Y6TynbP1VuV+
4krJWduSN5jS5Dnf0ClKzYoZHP6CHosiY+YVOtXeYzIIMGlSWT8HSnn5+khyjSbC
fAx1x4Wd8pexcpt0c5yT2fYNRKkkEmYFQ+7sbbJXYCbpOaJk/HFZlmZVDAy4+unB
0YXQRmpZUsind1+y/ZVeYPXx/t0rrnlB9rrzcnJ+DYKAC0SjPGWt83XJhSxgG3zg
iy34kCmlYv2D77q2krcA64E+c3eQLoj/+cPmFglSAEs29RekVOyGlNLDEvpJScml
ayfNvAwLByIVujlvcHMDD5TwWeYSizGFIu2UrKJMBy2WKakNS/mvKUmgWu11xd4f
zAxfTRBHA8lQnYt8nl9H4HVi22P3CBu3f52I4GU0r6pSWpG0Pj3fV1ES9Y5PkpZu
JiKVn6RxhWAbKlhDoWy9UNbrfFQRgy3DT8srh5Gxc2FyMXUPmydA4PGEjDLN/moi
rjaddAYN6Eal4tnM2RpTPKTs98WP+WhpdLQ+Nha5Z9CqB1UUJ52UUtl8wHWjFk5M
zwUtZtnxkCO1us5KlOnrRupaRaeA7LK4b5rKqCNlOiacpOm/zPP8MmBEiM76WLfA
`protect END_PROTECTED
