`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/w6eCgzKlIGoaxs8v6COqn64u4dkXUJ4jaJ++pTf6LwUIWflzrd2tSHn4D51C/W
utWQkWM63Qj3vuDujoWviwxzRM7TF0l5zNaAQdye4xm1BSgdbnL4eefnV0t/kMPI
DdIFgQtGF/IwNAUe59jWnmnyiX/ML+b09zARjYkPXLujP7w/qVWlFmaa9dbohc18
9GhdfmhGBTu3cVyK4MTzqDF1GceFIhg8ZWVVVU0fkN4KunhLvsvxWWVtO835JmUi
sWlPATMo/CwBP/jmmb/XDVx92LC/UqwrQ/1mxDJn9v2ONQTSFXASWfd1YVp539Nz
uC9cKz91AGEX/RZzItvJxM1WAUgwZR3ujM+tEm0IwuQm/1uvVCRZyLH2/oRnsWfS
KGKZ3MJVjQLRyFgL9JSxduW9oE0SPGRwfgDJflXDneySaXnphL03gZen2EW8fZbo
IQr9G5AK1iGkEOnyeYGM4J63kbUEhhwX13RYySlxNOpdfpj7CgFpKJxXgNxrihth
`protect END_PROTECTED
