`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3g6nFWPZouTJPYCS8NrsOaO6XRlIBugHZ1BDmpkAEF66yVQASHxSpWTV9ttlU3c/
gc/D1WMJRrAAoJLsWwN3UVnU/8rlj6CS3h3r/lin85tJ5ffwkubIRY2Xi+F+RtlY
Vdl9DsCeussbLiDm5MlR2MkSNmFNQo7xk99MUtnfsRR+CqM+U/4N+MT57rgYX7mq
jhDPjviMHZ+V1nulkArxy1yjfu8+nHVltHv+MPdCGO2ThR+UUEQgOWz4YmdtSvS1
GPloN1OxBH95HrvVDazE8UjRy67VcbActHzwrTKTFoAzwDaw5L7OwvWCjUSUKn2u
7vANHHSPKaJUuGfvrZrpcA==
`protect END_PROTECTED
