`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44W5AYvVatxCH87OWj+IWhMuMH0sD4ldlHO/TMD70URihlAKDXrzoAfD26Y7+7b+
pq5IeTx/YUbyPLxJRQ+FGaV+JkyeE5aN3r3r+I1xb/wQPmrPFnKUVyztcdjX7taU
OiZt1lwCVLC5ul119AzelXbqzGjQBkVxht1bdMDpaAFYQTkhywZAnQOU7nI3wOuY
2uJvwNOuEc7rObyJ5G9PwjgttZ/RqmKwI2+ZQRYJFVSVN9wngO0c3nZm+zVorGFT
qkXLqFxcdYAWNPcZGqv7CtXMGmJt6R7IC6zYzeqZRYWOt9I5IcXYN5Az6zZdKzEW
m/FcHNRiDh217z+pm19in1VKtvDc0AqpITY53cP0NVMmh5xcTSpwwT2MEi3b2cVc
/l3FggDsbMJCDpbxeEHbmvN1OyXgzShG4NBf27M30ZciQpQ+EP7EojB3pR4jQW0o
3lcVXIvGRTdS0+oRk3jE0Q==
`protect END_PROTECTED
