`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l6xwUbJG3nmaZZqNkM1yp6iRHbDU/K3vUd1FtfHdw4vwSvU+53CE95lvU3dxUAE5
7w5vJQqq9vYlLo/lbvC39IMB1ymIf1xlzvKj60fwqZoBLXLmWFyg4GJe9v7Em44o
2DXyM5kg0eXjfEudQO/FhnA6tAKuDaTfFBNa39OD/0Dc/27TOLSG4p0zxBeYaQIp
GzH8M4JWc3ULIP6cEsH8XugFFOeIW1/ZaAXB1AnMnJTSDITFXiyFweGCzjAhXzXa
jzNO2MtyTcoAsCe2Zy30c5ZVItZDQsm0potyS4CI+jPJ/J8Sch3PQuorQJNkKs5d
`protect END_PROTECTED
