`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJrb/w+i0UgXkE93aJN8PzQqHerB858i90zdmgLviAJaXEgorWPw/9+jKE8VoO0N
uTV+Kh9HQ5PGLkjxNPzI/W9sZ/olQTjOlREON+8qF3oSYWCxocSoTM0WSn/P+HHl
0xJPz+UjblOb7w7Kb6uiTPbEkxlvit8W54q6+5mOcsq7ZlpjjtTHMQMNVia4gzgJ
5TbALGaNGe1gkFVtZtaoHqPsM3suA52vTxWea1KNLlIX9jx1CuWwqnbHIcVnDZUd
iCdPVvInLcuAhn0e/DEPamXC7P04qhVbDNNCfS0h0d9pEy9x89o4B2zAYhn4A1pf
sZTiSf2BqT9km/xDBQFzMy3eC4WjaW8PtoC0mD8rv/Ic6sOQPPBaQnHG5gJhG8W7
A0By+g+6VLX66HWyVVsx7L/SKHTjlcl1B3Tv1MRRnWit1/eIfNjwOzuQSdSUodeL
/Omc8q6KUGI6Jvoe3TSddW7LN7YXimGhvtZ6X6O7ACRtOawcXQDBLIUSzm1skUba
HLq2b28cUpXDwr8UnVcLXzxRrGBnZF2apc2kkBW3fGkukmUQ2v8TevwGd01vapGV
yndWZHXISgSmtKxeSHWCt9J3hdgMnq6y8MgiyPwz0TxIHQACg8pPvDFr54Qpla2j
8RE644IuSq63CPymKhwKmgCIFReXVaEKw4LQarS0191lvlLgODCh7erKh3JG6LSo
zmuID8bFLyxSmZ8alXXtBmn1XNHNSmNIxVKzHILzPdd14ALpBojclfA5AVwip4gs
J/+478cZmYgeM96XMw3x2BHEEnTAPETnw1U4eG2pAOnC2Vnh+s8P+GgmVLj/9cKO
zL5kQS7OB8F68hyfHrmDZlYUHwTFStMkGD/O7/vs2AgICZTV2P5IfHu60HzpgrtJ
Yoxr6wpNzbYPVZUXkVM87C5kOpqUhnDITdN65R0U3+dx4+IqrnqgzgOXcBxV6/K5
Y8f9RhevjEYj/ssdh6BMog==
`protect END_PROTECTED
