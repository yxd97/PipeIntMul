`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lXoLdYfB98I48PC4YU7oPHpQCBoNXkFVxZVvJQFCRxc4mXiZWkKegN6VNcBuga8
RbwG41+TmMZNbqN/T+BS66HDajfjkk1XDXnLaFc7td4RDerfE7S6ZbTVFAM2oVpz
3O5teqPdyCY+YCuo8jZoRmNejyodANLblHbHheZboTGcxtY6PBrFs5I8CvTbP96B
o6JaC0x1AZcAb4oZvzzN19DXrPVOkQ4yN0jI8mdk38l6IrkFhESaoKNssvqdLQiu
8kM5EFBxtCyzfsadmWDq6zSWkBdiqQIfXW18+9Mv9WVbtD9Gfvz1v7Af72U+Di23
7mDTpkL1GRf/L4edtlPBStAThzfUTOr6uLs/wNEuKA1Ff6Yzn/upktqbzJjmKfPZ
Yh9Ia+JjpdlmlWxgw2nyKt7G6MiYdrtAzY/oS/zc2iA=
`protect END_PROTECTED
