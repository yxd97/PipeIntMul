`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s3tdmjZfwU9Yde+Kwb/efs+EyfOU3IKTCdelbqh03ZH49fNrglLRJpHYRDWJ7Mx8
8GpNo/8KovU7n24BajRHLOi3cnTmhGOlkXmR+hVOGSP0xh9L5LpRiQYdnoTKiPcI
MYPsSEskgDSYd8wZ4Qgrr0m86gLqHxGFE/KXKFUCMCDuXm26WqSwsmmcErqtJusL
5UXdUmou2dIeMl1HkH65g5DdT8iAY9nIiQf2aKEtdW6odSxGAwEzqHh3sD1ZmTRJ
0RClZiwDteIInARKVNZg6NDWRuUifcofMrn8vG0k7PbafX36y1VcP2BZTc8GhbSf
wt7ugZCcXi5OtOExQL5fziPCT0XzWfsn87+Zye67T0Yl7S2aTGdibUSJDzrZDel3
njB+oxzcWZYhdNUMWHxqtGqV93+O+ga2iM+todqwNjb+dp4BGZ2YmIdqEnGfoAjC
In0fjXn960D7D5+1gd9YOb9ztYKXILfNbZ9gHfy45kW6Ajatmbn+WlFJGktdjWnb
dye892mWWJGjRVf5475a6ot45MwWVDqeG1dklIdSd0EKkdnM+LgVLp8VPb01Mp7e
CKPv29xNRfo3UxlwqKPjiZthQzGs4u0tUfhvsfiBtg5GOYofUF0evxHCLeCWwAzo
oZX/gOAjJ1Y3njn8ZqdQ1d+ig/E7+gWa1Rn7e4xgGGL7iklyn50QzXwaB5Q3c4XK
UGpvEk9k7zJ0rqOmI4oCH95vNzz0aUkQWtwRfrGhNgSy3S6ALZoXLUrLMiOT06jY
pdS6Z+iHyg3Xltbk1Ty3KVskgdM/Y7KmCvR85KHc0V37PbIlZQTVw1av/vo5K5/l
tnUZmNi/1l5XrrQuxFvjzGaPF3deGwVmrobZfGq1qLuVZMkQNU8NAzFxGZRl6CZQ
gmGvEivwSiC3nRA5bZEaaBVavHcCzSy7ZCBMq3TrLGADu9EqfYr8j+LN4HYCTSuU
oipnE1F1vZqoBIw9/bDMNqnC6zIYAIM/KYGGJKX9D0rUUkqujbIb+zmbk8xbs4Xf
MZaMbQBIIW6ohqALV6glf6JMtzCZp+4Ht6/lWwe7Q8A87iUmvJkMIV0d6RVIG4u2
Nxnlg7OQsGkC5rRLyLWL53JqGQASqJ4Bx3KCK0SuTvcCrRtpVRm5o00+RovuCymB
38i+paYJ2RcDbb7yb2KStKslrDB0m2D6h1MjqWDEJNAXVIDAkfD4uw0B++F8hjpc
uIa65XRxHruhWpLLG6hBpu7yl0q/WSAawulMrG1zt5friLaXLC5RwwuWdptQ/Pdz
yB941HnFokC6q2/mXmaHdAmr7Q7vKC/k58Erj3Y8C0MwQv+W0cfCq/81R/y1ryel
Nd4qWYbJpixQ17OgFVDBuaM33QPrGUeEdryCzey9FuJgn5mgCKgIj0RER5403qi4
vZa617AoBKx7JiAMIYCEKltMLFAFSwhBcU9VtF2M/0Ktgvrg88TiCst09GhygtJZ
2DvYvYtB3yfKeM+quc8GzA6qmfqbvnKA67i4AvrqjuKW84CT7glrSysmb1eNun5h
X/BXhLXCT3XYm5q7QWF30K+YCwlQIXhykBq7IZHYqYdZTACGSZsImtMmHP85jog0
PUtUI2L4k0z2/wvywAfbtEsZbFEwjmFgArFB/ob05zQbrBz2s1/X5dTfT5DG+n4u
MEfwoDaPkUYYWGYaqPXKNC1kUXfdEojJlFb4Qj9X2G0BfWiwDIZkVWFAhdjWLGqy
PqI/8Uj2omDImizXnm3df0LtX1BXnfmkdDRxpxRIUF2AJyCTrrHFbgxJv3wEFo7p
DZqYGq+ncLebb5fWSB0QZ9mEYt6XEet0omOW0jRgI4+rO9eVLHk89BQ33avqBVwq
unUJ2T3jCS/kSYIQdd8r46ofYOx3zJ7sYcRGe2OhybJTSFOVbdN9smv3VyYH67yi
JXfxJzvVpR5/1qzo3CTYZKjVYev5aLeQrPlV1PNtFoJWe68BVa8dfXJ9iiFezmBc
Hs9a440bxeqhnuOsAOVOVjWxkGf97BS6T6fhO6EvauMRA8TadL9WcL58l4JK6Uv3
eY9EymWZAdbsdHTHINN+b89uPdkzTWmNSegE7cvHvXBxQs8RIg2IC9ukkmVyRcNu
U4+XwWBnXva3ysjxugnADrrzZt2K1Yuc/lSzECHfys9GiVXR5GBZ2ioioM2CIHxL
LmFy+AXDCDf9HRqTi0jKMMRcnBzXp6+lqnCl0BbD+gWXtvVTOgpE122Vlg1PtG/2
L7Om+bDZysc4qrQ0ZGo2r2dVI8UauYx1lIPFeydsb8a1vQ3g6z2kL70ijxl3ycJa
+sz1DpjkRy4DZyr9gJqdBa4gPNSnj6987yebOiYex6M=
`protect END_PROTECTED
