`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e7Q6sXiyZOH9RdQLOdkB9ThLRJYajBxPiNazEG5ON063EMRuCbHzeiddM2cOtsv/
TcKtWP3mg8wL6/EP41YiyiqbTl7ux3/jLj+IfaSlZatnUElLL3e4KNb7xuFnrfuw
sCzYfUyvEnZ0lUeK2QmS2mEeOYIvQkfy5JDH0UNiY+eby645wtG7QYpyQwAqNgAg
w5+V046Io2kzbq1eSkEi5pqqORE7xxvLOxGwhk2DLmU8SaUZ+WU023pmikwvwdam
m1mgEHZ8VcAz6fK7QHq7OxaKsknODrVC0hB5OGd+PmugWA8YXqt6mlm2M2YL0DAG
8RKViIHOfiXaniahVN5GkhzX5udg0fLh6TY5FyGy8xgQ5zrVcDwZsmC7J8wqytNC
N2L8TU5M7hZ8kSZB/IUmsg==
`protect END_PROTECTED
