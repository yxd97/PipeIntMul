`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29G9INDYhDl1iFeKH8Z3LoQG2m58YLN/eX43zGYRJbZM/Jwsb6ZrtLdeelwaCS4H
LeWVd36G5wRUpBo74xGKzaQ7OPRNPV+mZxZeKG8b7j9wKSf6pJbayfceEFKQClKx
lbTubT9SjuRRZENaguXJ7IyhgA2xxTi1cJExmlpWQQ15Z75fvmbi99uxu0TtMmZ2
sYpu5XHrno/F6lDiZiROZ2BmjMx4E1x6tbM/lEAUd9ouH/YxWPUWL785eUSIAUQa
FYs6CBK2bnQJztclv5OSung1DOS/BUJBgQ34aUeGnI16Du21cs4Yww+BiSvdQH4k
WdMkhZ9bpOuVMxomCfMzA+vo7LaNtjnD/WQ021jHDiHUfqT+xrLWz2a7F2t/jHcb
HrbZcn1J4Q0JVEHXZkYFPk84KOxWplMMq1mx0BTAHoVCZVtHShhKSqxG9Tmp/2Sd
kaEZiGeaR7hHRR5r41WQIy1+vF8nu/pFvFFEoqgN3G46IT12THhDteuqdzw1pTwB
gJwfYws3boh4M5yLgqpmAH4v+IcMYtjSSaPh4GfCEGULMe64ia8IttsXOUR8gIjZ
Rco5R3TJ8qMDsOeMDU4tYbpVA3MwpntVk4upMo2/B6OVU+i/805eeiOPaRknHEcV
XvWhf9LjILu1BQwxy8agVbmLrhLHmdZAynixQyv1M5BaNk1UohvRSj4STlYa6W9h
QxZGOzbWmH6ymjyswXjDNgMi4vLWXFDbiHIyZQMuqQfm2mIPZFzhaoHdoPIiIvas
O8KFYNcnnbOr2eFDtogfOjPP4b7VgcD7rKUkMHQ215z77FH/HUwvibwFCc3j0f22
jbosoBBg+mIr3mI4OufZy3jbv0n7p6+z++QdSJtnzb7CCx/3aqzwdIsEMCJGHICr
njzbh3UmMbN4dQg0/lQDev6EDzWhLCqI0VuIvRu8R2pP4Jb58Wc+vnriAsyFUXqF
uA/hNIrz+ioaUhKga+637nPeAToHtn3lyTS8FqStiGeYhRZ+zfGyQzf/RNqHob7L
g2BrNlSTxdakSLlBMwjhkdInH5m/2yHGHiF53hpjdvQ5vIQo522wzgixJxgfWAUZ
XmgUOonsBi25Rd11AhnhnwZXP5ctfDl0QrNTkUQYS/rvHmsp1AcswwuVyBG4SSs1
JvvfoRXiz3kZ7/DK8Co8d+FxBe9/tESK7ED6gIEJGODC6R2C+7S6i3UHrcOXA+Xh
ympgPmYE+0fnET9sZ+jxJ0+W2cGrz8keoTnJNlGztCgXngBw2scftGcctNoXLaZh
An796Q+NZVqTtfBAHNBe6xOs0Vd4ZJsP/keR3gj78TU=
`protect END_PROTECTED
