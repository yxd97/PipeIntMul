`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ct51hRI4WjqUvOnwxRO4mofq/5d/vi1oAKtkpAvq2V5wKY/YGT2/v/tb4OJ2rfNP
jBUZ6lYiFijCmuwjmY0u52ltDQfCmKMByqMLgTZDubzl34OLeijajBeRKWGTJpRm
1D849tjqiwnwDVUVZuoXM7L+W09XWkTKg9qeAhl8tP93ljVQC1UQKC36nrR8yxUb
epJeWDMMAmvbZsi872CpAQVnGV0IWb5VQcVXfoA9zeFnXnY9Wtpf5a8EGkbPeJKR
Wcus2jcuB5Bc23TmRtnx9WrX/r2Ypx0akk0wyYMCIDM=
`protect END_PROTECTED
