`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAS4On5KSCSTbuGIQSsUJrcBKQfCLF/nckV8wz3tWKN+svR+5T+JpZI2/glZAHZ8
TZkLF+iOHR3pFnkpir4fYKfyWMJoWd6LvrGTc2B5Z9iO9QxQphoIBSR6ml8uRVrH
egWNJXYNBpu32hArj430FvO38tQAESXpocdTvqubCGMPQnSJY2Bi3GD9O1tR2osD
JMqHt/Q3fxib2M3crIhDH10sCEdy5N8gVRZEJmha9HIL3KzsnD9EJ791o1Qek9Dk
5A2pgCoh20mu+YElLT8vCGDZHCcO5ZIkl/4VxBnGLRw889KJq02u+iC+TM1mBPqR
+rqJngdm/e8CdfKqSbZjimRZT2p+3Vw9nFE1jcNjCxMfUIE8HCquX4GnbkFFs9V1
Bg9onIgsaGgkssMfOJnXufdgoxnO9sbCcNG9qLFhA3i2ny6v2fa+BdJdfFTI/hN5
XHgut/t3qDrg1SoAKu1l39Fv6XXFtgrGUYzEeiT/EzSMmrVTzIVroQADxAgtWaQ1
IhZgiBfkuwJs/swT0uKtPtWS8JMIHRlrBpPKBjMr2+r6KC8g3Fe5psMyJ3HEFcb+
DRpL5PJ6I4Ud3K50A3/xzSU1IpR1JTLlpG1aaTG+7IBOeEk5qI3tHuxXx858Dv+s
x+dfqu0RAcNajACMHGn8MLPUwVpDRtlm1/qmdqxxkbBjL8xjVs5asJR7TZ/3rVvs
OfeS/+juQzkN/JzR184Lkls139t+GSQtS5V422+u9vzWNiK1MUX75L1dO2T3wsn1
`protect END_PROTECTED
