`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+SY4CZYn/Fq92K+sk/WzAjN/lb4Oe9b1KG3MjX3NwO1yxBwOPzhrkES56lhE7l+
wLFsCC+yPHM7uwbhzlkaOu0cposLziwH/NIPgd87oP9palPgdjmSLMHy+6mDv5Di
8LTUw4neRyqtRhv2Kuruh44wn580khSOsjiopTbPJ8oqi9pIll8RXyiEMgv3Iqf5
Mdd2xm5bHJVGiibN6dnvCMEwfm5CFjvRm/5WEd94IZjuCzIha+OOr0MWdcco5cMd
IeZcR3kLeWC5hfBlYsh7mA==
`protect END_PROTECTED
