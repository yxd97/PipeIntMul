`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6uV82k/mJMEAkBhMNKsdv7x1L8qHxvt4mFbdLsxqfZnN8zIo9UZ1aya0zK70Rcd
c2LLZDHlGrtI1FSw3t9EAphpnq7i4SRkmIhgnsIIr2EKPKEwV8S5SqOV1119FY7B
3+4eYogJrrr53eAAPlwN4d9El+5421Tj1aolG9jpGdO2jpIZIBSnDUmy7ZG1UxFu
EIlZoiV1yDM/NUnsKJuqw4uVo5uH6AVHcnS7IyGMUi9Dpz9B08X5+QCOGbAziwPo
TllWGLkP2+nLb29Zdg/tH49H4kRKNookq/nySFr7Dd5k2fu6CqHxCQyqUJCVyg7K
RUinn0TzpEETqv2NVdP89hY7QfOnGojaVm5DNlOsKsPldqF528KmmoWZs1Ig63DC
pLzc1rBPE79vTUjo0Jk+RA==
`protect END_PROTECTED
