`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P886/hyIcip3mqBz8l4vRX+cwYhs/ognlhLwZsiHElKdnXfbpD2sTbyeAAmEEjp+
/y10YnlYDMLA1YjwguyzLsrSfJlkjhXkXMKeKLu/p0vjn9GHNY9SkQ8jRyxq4G8j
9jBM2SP51UCHxySNAChC/s1HTXgxi3mqBTKLvsF5ro0ijL2RZyP6gRdLY3fCxGBI
sWSPvREN9ynGyx1wjZDpTUZ5CimAPFv1nZIGUkQIrDPw3gM8JccPF1cE3mBaSJkJ
o6dqV93JCE/RpAo1/QwsU9fXtM3JRUrcfIh5vn2rahy+mUcn+dM3KJryN++KWA3A
dqc2KDZQUUiyVATmwYwqRQyLLgFQp5J6qN70lbs4Q8i5gkSoW97DJkDQVSE1cT++
+x1VbGeEO3jZpxQqc69rrPTOYQIYOoVJbm3g6wu9kxViI47fHDk/K+8CvemE9YTl
E7gHCjdokH/oAa4O+qhk7Y+yki0FUWC4/WWOt15euWxnpNST6+jFx5LND0DSz31F
npJ49JErANK63+0LRbrxBdw9aIfqxGfeYoMZpfGS7IUseZvD5C7Ymr7Lpx8V69JX
e3E9CsFBztRsvS0PpO1aPPIQ7HAh79D8dROQ1DmMNs8CCdjASQWv401DNbfYmq2G
s+2RrLq2G3phuFto5UY7UOkcA1QIU6RKD2X6VHxGPAsWIJKkTaEy1FhHStIH8b8+
tpwxfGxbyXeeYXOv4E2z1xSB9pp79B8YXEASdKCokDIeyR2gLIzsQBCu2M8hjpiu
NrWcbtrDAnbGjeXKT6G77YVcuBW9Jlixapia1Eu/zSAVipokNBgsUDEL7LkEojZg
rDAe9H3aW/Sk7hksS/XwJihd56JjfE2Yxsyh8EaeEpxUuVA31GFYqJnck+tSkUBj
zXlgLVor5ryWzy+1l3iuwIEijyPKDalU20jjm5Q/fniZTypHrq9egzh8nKs6G1JN
g2TxyA6xwAbpAmRTjlJH9R7Uw04O0c8qDUHsJwMizz8j8ikqM8oFGvIQN2DhP/Zj
DA8DuvONkcxZU9LBdbIPJdmZ1YKsxbZur7w68VW5a6Y/sTixjcqHWyvnYtQuG9QE
VQrdDnH1bsBzU+ERtbpix0j/naehOIBuoXA39mvmdZx9BGqEx7NDvRntOuzLZ7Y9
QUjuDs35lQ7H3GGvOsF/4Js6FDlLxn2006EQi0ryml66OON++hTnAPq92s8dOPmq
rXUdtgTYmWbIKXddliR6i6QZDiMtKnvanPl7zV2jgki87C46x4Lu2fx4vw3n26QB
Ips1GjP1VxHnqWsWdZkCHvJWP6TozIkr53dgRUchigjHrc25fntOAg0fND7LlsdZ
zGt3YOVvlGnyPZ1OkWQGOMVb5tCgUN7/eOj+rYBSJ/dvbf+CNIiHrmHo8CgU/DyK
uJ3f6gw/+9I3AUdKp/EQ95meH4WaP/dXOqL4ySmj4UFOvgkSQgZvobmt9ZrNadVH
JQrWfSLiF9j3Kk+6JKvwHAc/EDX99YcVku252KABGxJQC2S7I+vU07Lir17UOJDt
NDXDcWj/uFQeTVQnVZFUNGo8215AXU98ObBsBiKxeOpQt8sHIPyFJm3jFOgjV8tz
vg/8FwFyMrhhQVMKzs36YcC17y+mxu9Z8701MKs6gQvKpObqdsoglq9oueTqbk/q
wcZDgyIOoJVLbTuK7IO/RptN9WmqpvbiTbB0NH9msuiM9kk/XaV64mDT+VovFYf3
y5/VrmkWm9JtLjeKA8VnwMFaxSR6mxPSRekq7PX34tg=
`protect END_PROTECTED
