`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
75MwfUXEN3barhreJXxrjVYjlQvcexsYAXk9FtWGnlwesQtLA/8a1YckNSQOMb3m
lrOlSPKOaFXaWtVz+2hjXiRbx4Ilfufx9N+3lW8Z25nQN0ks66lqgjzZ09OdQfDA
kx6yk4rYp4fnpacC5Niwh8TjpXR1bfc4miCWU2w5Ae3dRjEc6ttlXeoNnTAU7s3r
sbeVD2cVwbPrJLVEwCukvfJ3Ymulhg9fdlFzjbaJUi9YF/TqjzD+SZGomh9xpVwI
dTmNMnY9tmrmDBPY7fS6GuHQ8orzamZpJden35ytdRVb0BRRmOhbXUvYmDDQswL9
FqopIX4e/e17ygje/a44I8//rfIJ+leYrfub41OcCqsl1Rhm/NqhqPhPk3bleQr/
foRH4J0vdD7GGmMWJBPiAkh3pUDRZpo9NvAKkGz0DLVWPWFaoE9Zh1qY1Tek2lPd
Bqnjy3y42gWUEExdzi3RX1vPq53j6Wv4ldNp68lD1lg0fx6zBZzuV+YhGvJ6+fKr
nx9+zu9nWXJh1fp6sMfoFpq/Ox65jFdX4ThDGsm3e0FSbAEyf2wJItrmMPtwdXCn
vq4yJPo+14OQd5PDZk86czkpgeXqmSrv0ZdQmhCWEUepCSvWubMpcLqc4wZDZCOK
XRHomkS2xQSNC46nrlk4msx0wwJSUGUJWsM0GPJELHawo6X3oVRF7BvYLD/DBniG
7DJbsUEbTBX8qe7APyapf1UfaJamIxGmznRegJfacWM=
`protect END_PROTECTED
