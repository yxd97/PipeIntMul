`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3kWTlKqxoiy+vTPWewStmex7HByr6EQWwKR13Ufj9L4oozRnkr3Omgdy8l250O5
ooYWEza638JgzbBPi4xANbtKKzM0rbMg9A0VuwdLckMvNQaotDN5Vp8+lob1pcDo
VX4KVYvbUtvAW4Pvd+srYQ4XLWwNeZXHmt4qGA0ttSiWR5hdvVKR2Iu8dBa8bgBG
bMjvdQH0H8vCPe/X/6jlMvkkJh0ysFtaSF1PSWCI/BDOja6hZtYyXo9mHwqB9QxH
wsYpxgsZkINhkQDq52B+pRS/M4xPdIinfxGaAAjAPVf+pSM1gVwoBDcmISKKRXjZ
4V3Ri7YGUUvVGZqgbMI6OhA/tgdPMO12rBpYfGxZ4oDJthk0SGCHIR2j24gBKkMb
83GE+R7Xy3K26GLRZX0UJ4lIzJbw9Wm1vV3uahlv8LjHqVs88/zBmPTIGLckmAH7
TMqiMT91tY+uJNk+xmOGSmOOH32UaBgjA2Fwcer+P24=
`protect END_PROTECTED
