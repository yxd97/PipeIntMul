`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QtJ7d+am+SJR+YqX4R9VeF8yuRP09a6EgFKNb4FbO2vqGSPaLm17kld7S4BOZd/d
MPEBGKrHTM7FwIDXgEA/o3ulv2CT3/9SxdSWO07mGH+z2xeRtxl0VnTnYv7SqawI
lUIdMX/91Kpn6jAyertDKg3ZOoMoPVkMn5fYzx6JbJzpq3/5DGh1ymkJ0B1j7Bkh
mfqPthI6gjwjlDDPc2bg9FWg3VT2PfvvTudj+PKLX9xRxvhN2tkzYLF3gkdjCK7F
hi3JZwoxCCW2jXnK2xlkjPJBjWGCfgZ5wXXTS+3fRcyVHa43C790GGmOyQRsbjae
kkmAArGwce6g2xl5dYtZYDDH8URsHcDUQ+zCNarV+g3P9PUiLzx7mARYBKMAROxV
E07EvDPSn+4Gkux6VECb7SwpEGFz/W87fry4pnN0vF0TEjVdHhpVFGmoL1p0UhlL
7vYeIOCR7iNT854BkjsjxZtiksqQs5KVOOeudXEiBl2UzUDokmPEYeW48MTOghKK
hcqiVYcERbKcRkDlSeLqAf0V4+0e7geDQiPjoXaOsgn7+yZUHtispRJVDshYh2Aw
7tYRIeDez6oAJzXh7IiokwYhkcCoDOUYLtCBa+hvGQc=
`protect END_PROTECTED
