`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AX2pzbwAnNOq/ZUuquf3w0h75o7Ibe0rQS5mXyZ0j8mCTJ7FOviUrLurpPZPNbe1
ylldcF32A1xFQFXaoQgbnpDkKudyIjBQrSNEc1S//bFB+fB8egBnCp+H0Vs0w4OT
Poujh/5y2HsM2kCvOpNgkmyjIrZFE8+stNdFG8kCLqqHLsFPWDl0wr90pOS4CLZh
mVbGaMUkiZ7awyf95hi/i12aKCjGZ/bC8zadfjGrG/Qavn5z7gEZRd60z5IZQ2+j
hHNljoL3gRgvrWiwWT4B49ze9yT6mr3StXzHi0y/3oDA3iSggZe2N88ZOYXGaLgN
E2cxrZobkL6JIon0QPzwuIlMP0+nrjZDDvRdSn6OqorcdEfTEMG0CDaxZ55uqXqF
wp9+yLSzoBcxG3mixhVhWavZP1TtP+w2JMt9k8Kh2/jkq9d6Jes5zBVnoDEnEYpl
nXPTIn4cgmUZYDelFt9W6PhhpbQqpM6MvVr/YKu008KCaEfNFtMpqZzS2nnFcRPF
Zi7jzxSnODXmporSoaI+gCLJJJ8HhvERIM0EpS1QX/SvS5+7yEH/bMeIoIpvgKa3
AdOELhz1z1mTN6seonR8nrbt6K5tTF1p4rBXhpnE+pGrDUHj72dVhZ5D4b2Avrwc
VMEjqT4hb0eI693NIWhsNLWJ/0rnkYGGrFIZUG83Mhpnd0aI5ofd689/nX9WwGI/
PSIDjhVMh2YNcbAFGcIvZ6WuqCmsk41ugDOqrJPvRXB3fEvQWgyU1lZCWYrd9NUA
vh04BZ24vnx1nu8gsjDnC1Sr84SnKYvFXGnxOk5ngn8aj/HDKiV6coBme1RALFmd
WlXkbzAFypM/zAKp01LVdtYF5ngfJuWZf8pMepk2zB56SKq5VVGxsnMFArZtG02C
ndaKcgPGC3UAby8F8wNT1odOnXb+caj3HIdVNdyVG+vKtAqcItZ6eKBgIuqyy82M
7QV7TLehu96hV3eynoNyG8HR/eiXC6e9+5lbjRu4EcKWBtNL8jdtE8ICy3G5a84T
jQ+bVarfnhY5K6a8eLVtAOO1dh3t6JPclgYNrajnXzpV6rXxzP7H7GD3uHozOHL9
iVys6GaOp28k5IFKaqAmMCG+wr2vj0+yWWgu+ffItm2G0aTddAk0WJ+jW37uguST
FLHKpfRgmSqUpie+cQtInbr0DdZ+Ou/gaFPCtEChMzrlActto5mhOIX/I0ReUfHp
seOonPk+auoga35M0KB7rQWMrTi2TrJLClaL8LXVzj+ALMYr3BtP3TKGlndcsHz4
Ima9NhdfmjjVadPnZisbdp5e52wArLk742l5rmT4ziHP+lILHYXp9Nv3yb0xHXv3
kaP6Z2Htb+q/7Rdo238GjxVvoFLq/Lk2Ig2arS4WqRneIC33FkKaXyXNlnE5LiXh
dqNF/i7dNq4XoauuEPdp7Pmd4J60RV2jcSZVhQhmp2o1QPmLO6kyfzZJu3yGZ4ZF
25UXhoBf7Q92jPEHrSQnwIlXRTTDRuXfTcJX6JVpnxfWw7FObnu/P36D3CwO6bkA
CJwURYwp+URIhKSSgFKzZoZ2S/48Ibg43eZRCdxRxF5JMjPZZ/0TX9ktogjK9HB0
y8yJKVafF7cTykLUdbHGKgwYDmaCAv0yPfDkmrHcfrIvdQYM/mllM+FsUlQST1Dw
yYFuBhQgbAPVqaiebF/t2zLDAa51/KI32ZxXz8O2MtDDY9mONfcOZEeHGq4WBwSs
F1/kkRt1ruyUnmE+l04XVCeM1ORr6WMbAn7oAA59WN0DO2fiJrVDu/1GdfKzo/gs
HTJhnrHHWii2p4KP0ZeKQJckqt6wBvu9HIZbC1CgVLU=
`protect END_PROTECTED
