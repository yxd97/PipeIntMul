`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJ/4rPpebW0bBmOlBsy9VPUwOAnbaXOwiEN1gBpA4eEzPvAuwQGWAMlazCNb74LL
7ubXAVjTYFDT/Vc9fstEGPuKPd5hgHIGQM3DL/eEd96lQtAbYHqESP3K/7v9OoOK
FfL0Iz21GTb2t+F6r89iSfNZ5qmuAWYYGOc0FyKRt3cTYj1wsE5CqdlVA+L+9Hb6
krzn7+pgxV2m0CxZEYj3tMYk7Ism/lzVoKVYfkaxHY4Sr9b5ghz90COelSulibRL
nIKsdURtgiinQmL25VqUkIwhsmYCDsA6BrfoAvygTxHlnnBia4IXEYmskzmIuBZN
vrVlWOHaZqg55WB7x0LpthB7x4tdBn1tLUfqnPVRYsmyWvvlpybcaXhchsh7s6Qv
y8ZLtgjuvjQrp5eVi6UUQIUZ0K53MaRMdN/hYbzSDxpf03/9LZpA0yAkbkSPKuUG
2W112DMb1d88v6ecUBjmeVmxjnScZYJSmkeaSBW46QvPZrTtTxzFS6dnLxehNs0I
nDAhbvYiCFC73Fm02JjOprW9DDxU8x7NAsobDgvGWuB9L9dxX/vR50LrnIBfTVVb
rv+zCZtJmRwXGnhPi4O4IAmqs1fPVpXuVjmIcXtF5kU=
`protect END_PROTECTED
