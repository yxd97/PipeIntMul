`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjrDCbW4+8LMF3Evo/waduTuhLaNXM887vrNw4Gtart6eEDsSaL+TQE4bpMF7m9A
nHvvM1oVGWUoRpQUCYmO7Y7DrgQ89EFbvCDuqEEVFMJSKxpmTgNPYUPp9W8qyczN
iA+9XElCe47lDpbY30Xrb+N5WJye2gmk65Vxk7weO4vT0rqlAYWxgei/tSxICCTO
ng5fE7y9QxBb8xnfh9lPfbN5P4pX26hFz+udiQSzSRqTvC9DfcIRQ5Z4L/yNEX7A
OZMLIIWN2vbVZq1FsMMVsTLnS3jM4wvVsbeFCkaZewe8Vz4pi1w/jrfZM1VkxClj
MJQ0tvmwDSnKafaj0O0JUQaSVlEJmrx6fNSFSG6Wg5vIFtOdM/JBZomqmriSB2Sb
ZrA4IOinnTmOKeANxP0BIDNA7f/Iw8xh6K6DIgbITfyrUBOyjrEfYlG+v5Q52HE9
yt/uiP+dV/e+8ODcSTQyucd6GazbWXbf4TgswPjveVqR40rA2qgYxRUngspvvZgQ
NecaVAfBYdBWeBrcaofwuUo8e4bt7aTlpbiQvjn6Jg7uefVKCTvZ11ubt9DeEHpX
H+Bv3uEfF85ZnXwyjGziyYam2QMKfZD6HY/V5KyqNb+t96EwQNXdjOmMeBnlZZ7D
7T508l6kuxCTCojrsZrBGnrRxzXIclyeMAWXChJXrHo/Gv11dwdlo9yTTNXeYID2
5QuUvmmFrwP2DbZZyA+u3WIMhM21lQSZ17ziJG4yNewM2kiz5QCugIQsiBYVT7rJ
esed7+OQW2v0ZcYN6L+NeNYt4u6xwn/N4wOL2AXc1SnCPMFXiSYqva1Hmhitlaz5
c/5u854tgYO6o2Fhp7U8imy25arldXeAoRTpPgrLd74mCFMBbSx5l71AVAjj7qrD
hXqaVtRkco1ly1pYYia2m7NLozu4PS+4rGcq1t2QcTRBaVunKbzAesOAUpxdtLLa
AreBIQFAc+lbAKBgMovAYt8e+3mQ2bwqtfQmoFVqBQ/HAnMWB5wpDQGWXvlCa5YK
3cjD3VICcEAdlGPG7Jt0siuDx6XPwUrwgYkQdK7OaxYF0p3wlB/dE09I9PTdO+/G
nho7VUdhNmSboA20DYEozrVN8BQm8bTTdjfGlCT25p1+wy4yZmF9VRVC1/A/rnkx
4oiUdq+i884usN4nlS7yLYMhFY9MLZW0iHReXtJ8cnSYMJ06m7LYFhTnh5wXoUIX
7WuRCidhfj+1XAayu6/SsuoLqfuPcYGb3S5UZYgGGZ2RD14IIoqAIPFFSST+HraT
5Y7zqHbhJZvACqZq21AYxi+gq3xU+ivwMvuRDbY2bCXXAXQsplc4bsCugcjmwepl
Q+as7l3KdCRFx9t+aVRC9/fzx5RtLlR7BgzGHsOLV4OJflraMRYhzuIiZONNUowt
q29+gGuv1ujyODorjctk8Y5w6JPJ4U7UEpHoBw13VkSjv1e0ljQ8/wW1uKIslVQo
2QvPV3DKnwQgz4/1ceGtZS3aCrrYPPbfZnpLezF5xq+amx7LVWt1Ut0jW/gs21Zs
a5EGO24CXVLV89WDUjBls4FdC/42boqLNG/lz0eDI/37yVcIvtVnJlTExSDVVX+J
d0hQAhedX0XFJtZMe95c/ER1cPhX23ylhKBzP1o0MXqn2HjnEwxxA0tK3BeZZjzT
MvbP6E0AcCo79nJzJdKh5fiZWH8BeAqTiY+lnQhym212kdksGfPw4XhbmpEIAjIu
FBccYjrag6du0u/Yu+F1ym66YUanbOtnNZyLP4BoutYe9rmAfLp0t9ytSSuvFbQ8
NSJOM29d7B9EZWnTc2nH//HrDVyqDaQthHz3QsH5g3/SlEZHgNbB5TPfGhw8/qGW
dNmalFQPWHIpwXBbKVfgZr2o4kRrf6IvlVpByruYvhvVLO7qLXhP6tN/0OhO9BM6
nkch31lCIyGi7XZcZPy41QZm9NIT/IHU2W2PfbjgTZ6U4IBHJW0Av4zbYmsbzNGn
kPHENabHdIUGGV3900/V9yY0u27urND1pXZjASPUE3t5eFDMQ3ZB6ScthJTmrjZZ
L7I+xbZiSFX+fC+a9uRzQnNkCprlZE2be9BaPmSglE2e/K5IDjzA7zbrYopWiTz8
KSDLoGXMIoeJ4G+LbjlWoHIlPSh8Wo3kf2Xe+1UKD8qmg0Qv16NBtO5MUmIMR8dD
bKZYQgWrNaZV7H8ozgHMpgS+4wc672zz3I5wXS8fQTGqlhdt6mIqniF2thpT5hpX
9POreG+qBbbG5eEze1VQO1/6IMbyldVJzl87DEQKOEfZ0ojX1ICUjnZsC9MdhqSy
RI6ydPWoc2+ShZVgfabbafANrbjT2qy+8ck+/do0tp8N8PWrbEa/rh0DLLkX5qmQ
L44258qn52Imt4i5wQw0+5GB5IhXMt5f7a1J9H4BJiL+kU+lv4M5zEya3aaN+oFZ
8Dla9wUimouz5w/FoE4mqnX0CB0OsouV3snZGYGUgk53AF+ORZFvRZ+gt4VKGO0b
QixNbj22aBCY4YmERQum2ZkV+i6Y5JYQVjnIRgNiEXOcyLBQRJB87a7hV8RZ14IF
OilETyX8BA6VoiAIJeK3tYg1uxEagNj2AnRH0QslroeV72sitQ/rwPChjjhFabWV
Tzf76Q4Q7Bkw4SOBNJ9PLPeo493v2CnTYd3T2iRc86Nvtu32MdOLc4oDqeE0M4os
akIF3eZYvIZcntIGStiXruxhBfQkfinvlVyHP7h5jsNQTSrNKJOSuG0rICCjNb/Y
ywafuKve+PQ1UcSf0CkczfKXtswmeTDpiGvS81s7mPbn5zbjPh+/Wq7lTju06/qq
JDor/ZnMMu8+jqOd19SM/uV9ctiMDC8uqVpX6bRJRxUJKhHIVlckFZtFD82SeYnH
OHbzXxoJ3UZ9XShza+sOOwuidiws67Fhao4Lo23fCfydof0/F9PPoC2ikcD3lAJL
FwQwpes2c7djU+1FEHV+urrB7f8VrOTbALZd3d2ctzpIUEcixk7RymsOrE5sbdQu
kxaLLj2Yv8qEwt8rV1t9IhUS6MqHcpRjTtjy4S13ZiCuHg/UeW3oIfHxsT8o4MY2
K+LKmWrtd4oUrnYYJwgZLcYXOwC7zOHclXxzp1w6LlHWd2ZFDsLHHYIj/KgbLSiN
2CnEODafLxJZZx5AZK2vSUAuwNmTFvlSOULXheEPb8DadS652+6MeVKJIdcvECct
g6jQIo0pKOrpd19F2IrQljYvd4D+MNR3/ipHXAon8rnf6VXD2IT7La/UOIl2wd8H
yMjjeKHVcZRVXDUbZLeq38ATBBBb1vDb+OT5Z6TrSfasQhiiOajKM9Axek1Hh3NA
LH+o8eFTZZ3vcJ8PAqYK1GxVQdHvn50q/jTkRCGoVe2lFnolYYA48EQLDTRXR8Hw
dDnd8DOVElJl+TdCYTpajVEGZ5rzN4qCc6z7Jfiosr5A2m0xUAZE6bEt9l0Xfwr0
7ZNZ47Q/jju1RMzNkc3L0TT/OJ3eTWXMZn5syuEPOaVNwhYNf+z97tYqW+nhkMbY
c/ON35kE9rOc/tESKrSOIW/73zSHyHwOhltkrbsfQm0xfaeaD3+JI34BdmX5MwEx
YZGfNyU2O4SZd4VJa6f+0x0OGtTlMExKssyJ7Gghnn9m5z8zOerZiBhWdruwvzO9
jv7rpfgxbEAWJgJIkN77DVmVdKQFW6wS+qqNj/Oq5qinkTLI3sy8wME6G+SCilyG
giwjLDI2SAgLLmiRfi1DGbMjUyc1+Mxf96DEvqe1gucmhykkYvgskXNArda2cDN/
98/SWldQ4wa3t2XcbDc8DTebCcwzG62KQfyqerzTOiOy/dZiD3uVV0Iyr7Yh27Ai
mrE5KHE8j9wBIkbb9dfXNiPQRH1xCPtH0wKvVJqMsXLMTySxe1BqjBvJVJ+ni1N9
OatwFS86JEtHmgoXipvUqvgRB9/SWUUN5McQXHrpUmmtiDz3mUYOqRXEYR5K/nST
kRoXfC05ux4VEBQntRz8UPneOLwFlvFd/ZbWcdyNZguy9dRwUakIOqjvZQw3jrCo
gi4a9fYKVWMN8l6JBA3ysphSJ392qe63BuT4d46tvHOKJjPR93MoKA6NChERMcj0
U2tSc7YVHp8r+RVelHtLFvmMQwtSmbgFu1xtY4LtD084NPa0xbnS+5emCLuxgPLw
OGjMSMiYFShQNvIytDfZvzqLK+cYJn/mmepV3g2/HyaObcPMQNw/oAV0lYqD+3ON
Enz2yYm8UoP9XInTbzt5jdfDZrhOYGdKjtN5Y1h+zpbNv4TOvU8Q1jzRc36FisE4
mhhskDtBm7tD5XISiACTgmX40MvGfr+k2R/Tm0GjtL/T6Ccl9knLPARDLlXHhleo
sjizhq52cSfwEHu00qsNSiaDpOE+xZ7wzMl4Ndwzja3SrKUBIYnrT2NWDrO7WmGi
giod/XyAcnmKcfUBXmLt8u4vLyht9cJZ+YdWmnNAQAKraxFsgXOxB6H+z21lmmTn
gz59IjENenwJKrK2WMJ/j2tp1niKXA28E3oNepVf/5LfSGOvw4LqcRtSzv8ULRu6
zvHhGyr3yyi50lZCNe3Ws3UTSyf0wWAtDVcW5TekgxLVM8wDA90lBaae1oa18y3v
JjIZDSVXpUtW0EYEQv2D0sMnQ3WZK5hlL2k0CCyiIO5cqRnefpGcFgASSCdjkdkB
to1TRlSlrhmo0a/4dmv0ZdMB2h+CdKAklM+G5zZMT5Wjd/m1PjkNFAGAA/hBsgIt
iFkuTT0PSS5EZvBNaA6821Xf/1x5+IwYR3MVSLeBDSq+nIKH2Q+7QB+xZ/FlEhYw
hWfbQZPfQlAeZRXJjcsSgZ32tQjzTXt5e3bdM+aGbdb8XPjwGm3VnecLLbd0+ufv
9ihdqrvDhJQshMG5j/pbI3CtQxBugeuZCaeZJ6NNh1JEzaBHQge9aWTU8tpjDR9D
sBLCJ9cajDGjza516d/+2bSC90OGIdfwFrStJgIUsN3IWkOmrZ1MPjbonn96w6bq
0gEgQR49P7HrrYkez/0kTJJGyX7yvPteN+FEMJJ/lcfL3ih49iw7V7Mmu1Yvlt0L
qBVIadGqpqllPnToiArZl8QEhSWrpdOY92phrWpNwlTEeFfRQ424JfDqQU1k/PVR
ZxSPZgfhqq4/YnnyNkD573Oyn+M9/YZSVIy6QP/qqgNoOvrS/1lZEomDTsHcaVh6
YkO44u0XbXvrHSqJhBpof+IfTNLBY7KDyiXyGt/Qvcf/JPt4NYF/HTO7g84WxA9h
CIyBs2cLXtg3SmoTJxi0XaicYp22tRA1s1bEKApmyVs7FXIaKD4IxIPyvObENnd9
q3UooiFKdInsW5i1YURvanbBovku41BQ/cZWG4JQ+FdmqI2u8wZFhBhDktpx5BDg
NxYTJXC5pSlexBiFl1Xi0kp5k2IljDoK1FB3cf46qmhCmPwmeE7Lhj8rapSIk41M
/SpIWJFm6zZbdPv3Re/dmmTFJ9QnWm3gvK3i+u3grT+UoSt1j7o19Nqj1L0s1mEd
xFEYDokKKqiZcPcik6TemGCfK5DXeYK2EMACz76CNajREUDq2tobyBbnDPfpjZvj
TjL82RMW8ZGOTb+OedNohNvGmd7r6TbHoInNqbP8CNJxDB/Mvh5hb/e7wYw2i52/
90NsxZKXnqTDIDlnGiBnrcQ9a1eO5nPjJt3C+UVnSwRppYd/fDKM0/9fUg0q5dSf
9/XlND146s0Ru01KuFBsK6sVi8p5yrcUx3dWeH0uWrpP2Mgax5HtzMtyNMy0N9z5
d+hXxnR0Vs00QQjvZS45usVSz6CNTeJDbcR86t4PG3zh13IL6uC2q8eqtugLXZbX
5koZna4I47MYeTn2DnqYUv8C72tOS4Rr8CnnBSMSPbPKM8UjvAQgmobcpt0d0GF+
T5ZkkwwqgZhihNpy/90s452x0xGzn/5Pe2PFkLQKenZ/0/0R4wKmGVOYFlIgy3qP
R/Hd0ly/zZqRpvJVYcgdxJeyesALHp9gCO060JaIQa0WaW9yH3ksJSiSFPAdy65a
63j24wotlaHLHbsyLaQ3W1/VixDywywxEj44OYd0eyz7ZjpDVB416UKHHD02zOPA
QYCu3W9PwCc9L+sScQGPx4nOsdBYuGeUJkaFdI6bQkFEZF977lZo9HTXtx/nVW+y
wY8aQxwR6Mu0Shw2s3F77U5uuPH0AzE/AB/hbB7VmZAfZ8aMcunrZXw/oMcWrIEG
H6SjfeXuaT9/7JDylhSEcIzzScyEy0ouXEJaIWrIRST0MA4elsBOp7gpee92pMYT
fNWuJ/DB4IkKFaeHBg7QHb5FxZ49VnpgnFDrhw3bpX+w/hzRykgWIUZtxTZolZIX
eoyZkrDvIK3LAwQiqMVJDrzTN43DNSO5I3Cd2WAPC8ViLgo6Ed8GaYy5c0Rviww4
SbOSRTnusOmCi0MhB3CcX7Njwm2a6FSonS0KCobIYS7CKdTg/eUBmDeHkvny5kQN
YVNJXMI1tn88p8CDEuLifmaciRZU/3vNpuKP6HOpndVoybjxzHu5uh8GVNOWvjQj
gaNHkBEZssKbgptiFhHeUT5AdcjXG6E2z8UY2i4Xh6AmjJnGEuE/+7ROJBDGEQo8
dxtMtFQGR43J+kUjJ5PoWMp3IRWcFjDGAD0oTE6vH3VA911eHt9jec2P961R8nBd
txroQauw8Nuri+8qp9o5OdwnYcDiTBljxpqjNkVSRNTzFB0D1AkDCFtCW49GTJOR
2v6p56N5KMMCqmMIlTxaVJGexPoHT82OqkOfo7nV0i9uQU2gdOLNpvMLtZKnt7YZ
wMOtWhQgumPVA+wLcG1NgsY1QP3WRutpejX5Ai26gkmkSUosHuhXblwfHeKGQfIP
qTAQnA2o6ionNcKCko2fL8O8ZuNzBFGBnpkZZsZG6QQmkrvyxECNBpKrIL1Mq0Rx
CY0Y5HNYg7W+Idjpe16lpLsJAeAkNqZwwX5ZCkJwq+BremI0d0QbxpycQyWMKYqp
wAfmriGUCXWp5ZM1KdG5k11CxwBdTbtMrq2HWKNrx58M17yXgCvGk+hcdJlLnmdu
rOFB/wyK36n7LLqryxV8+7JuDhnKqiv45pCEZOqUVdRIPo+u1qVrZdvjRLfVzcG3
PYWRwh1xWzIP2Dz8HiYO2uw/uNgyOcYoQqg1BCrtv0c23PPMKuRoPsdzUSaIrSGe
DdXpUVLb2QLif5X5AZgvihp3y9rW9u41F7zQeOl5+ZUuHx0uXnVAwhJWZDJ6LBYv
MQ3cFHXA1j2oKTTX7rhLwBljhci75ohtyNsM/V0pJllC4qEtdIL6h+x2Qu0pqpwD
RDUpud95/aYrL6VXMQsupHabFlWItFFYC8Y6VBjbeMuq4IQxBp8KfkJoBs7hVfIC
M+pw7LG80nftREE54KemHRsx9PrSFWwWsYql2d0Hlmw=
`protect END_PROTECTED
