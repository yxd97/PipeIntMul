`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xpumbi2p71LuJkqBT2wdG9/3C9CbVy2J6RzvIe/R7EJhA1fg5XIHuDEmGA//n5dB
hJYLlxKNHiQhDTlcuXZ3Kkti7JBz5bb0oz/MSd/IiSSMr6mn/V+SHVZSEzcpvyRf
5135tZvLclKs5Ju1EFZGuCKpcAldHRUXHU0aAglw1DD7uB9ee2cIzeeWi6bWyVzV
7vg+HOtKOGY620QZjpO4WJwNAtFvbteWJlV8W+3qgNndtqTN/cYwv4kUYEQRlMY/
L7oWwVChwzHG1NRlXEmSqXtaUEoy83vZl2Z5/wlD9Q8=
`protect END_PROTECTED
