`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQds68qJGfZzmn3apInC5OjVsT7FhEKgkepoROYvKelEfCO0ilKCdArwFWZrET+h
2HITDCgF/bZ1JmUR/K4t8u2NtgDYws08qINNOVvoEgREViLkMtqXEtz4Qqm7CmpZ
uPXxM0DLXkVH0MVDTsUlaxx0ked9qOm4N8T8SRAobYmOYZMrcww8XdmTx8+K9ucV
0VRZHCz16PEBtk5ppdcyzCifQ5OO6xGe1qHNppOO4YgAPpfK0XvTnOcN6bp24pe7
ccsop1ZzplBNAJlEWNmB/Z7pHJPhlOgAMiH2melND407ACw0dvU2oCday7dKbj3u
lU8feA3DjyZnyQWKJbV6DA==
`protect END_PROTECTED
