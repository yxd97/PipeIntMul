`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ihl6vQTOhhUqV2Pv0Ra86qA3GDF6m/XBQlAxQIwjJVoNObn9icKmHjj/ZR4yUUZy
iAOqJ6qRx06BIhi1+4g5s1KXodTkqA+6AsiTSAVFk0+ACeahsa8HCQ5CkGRgRf+Y
TjX+em4V+oslNT1CUh82bbUqgVEEs9HBAQc6lZLiOQsfwzA8iMnCw/rqSp8BOFJ1
DtBNI0e0G/pYduvc+nUw2LPSQk8Gfoh4dHsQuJRAl8HqxwUcwR2CevabDRSMgxN9
CtzVudls+L+/F5oXFI+kWfSSa6eObHRPGvZhHVOWiVIeFbufAsBWA4ja37daYNcH
Irysc2WamaZMFCNVdSG7Xr61yD/UCd0sFAk81AiokxI3hGkVyXL45clB7KzVVpf8
ZPHU7/HeS/tKtvoTYisJFoLlNE8caWvZtCgzXl3RYPa97jVlMGPYBisBp7pyNnGT
`protect END_PROTECTED
