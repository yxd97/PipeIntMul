`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/+k4CnYYeVqHgyrKzhjsS+T5PaFrySuKdVGE+w78f/ICBcZH3SFSuRVw1AAq2HA
6zIgYNOrFbOi/foqLY9y4qmKtjKEG6Ima6q/ntZlhoJ6okStr2HcuXnUkdXl67DM
qFmuF8qR/+lKe1EavnQdu441fKUL7SowEKiYlCObWomapF4aKV95krovwbj4/LSt
mBB186qdT6eJSLSyX38c4663uEJYu7ELa1LBmuIEZG5MPp47+d+j3GV/6+me8eyB
cTQ5eaIXnoPj7Aqm6I/m73rkHn7o1Ac4O9cL3kSimXA=
`protect END_PROTECTED
