`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18HWzq3h/33/l1OtDiuUIkRt16TaCgpMxREvEyhW/fStU3i7j8tLXtv6MjSUX95g
huFHBn2ZBbXZ8iKfSoecLNWN6LJBliPLesoygJzFPPidloT7Fe2qEOR7NxOV9oIg
6v+e46qJnouK9IQlDONluMdBRsFqD9B1GgIndoFTWW9/H6fRaegbV6nfMcajl9DQ
w3vKxUChOe3w0TMwZqNFK+h3OVhoavaGJ0rcDJI8L9URnzwGA1fB18Kqqr+3tlOo
zzKzW8UIMPyUd7pkRrp8CPnI7HomhG3haVgSlSa52M9DiswBbMhxvAzoQ7bjLwHZ
/zevfmPppDJJr7qcr3jUtYwmDWWHPXF6zkjZrZ1qbgU8uKuG/pvcuRFwVW1Sm8cj
+PCYIlsKNuGDn0Dk+zdSPUzyrl5LgkfT0NXj9dXMa3E0rYjEa1mGimwnfzGa7YEL
0WxXoR2xGH6uQqNpICYz9VUEGFlx6LUlWPfDDJO829sLtqEV9N3pQheE0pWWfgFd
3U6HBWCRzZ3bcKWR9Xl+6MNnfZnd7ujJr5J+Qh1J7VKgaqPjMQS3KAe4a//z5TSb
HVSCs2jfyt/hlPE1UcY3kQ==
`protect END_PROTECTED
