`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dLixB7XVmmyayh4pi8Ss31MBn29pGh8lC5eXPvEpK6mp9n2Nxd01zWaRmu1nxF7U
+SGQwvbz5/GwhXj0pFbYM/zove+G0BRJ803vax3BmaCVFGjs4UVX7UMOWMMjkeUV
KJv9O+1tugvB7eMUZghaKG4egcMlADrBeM2kEjqEkSxS5NrPDTLjuYZG/8ZYMCr8
CjCbV0C1oYObLHYB/gcYtlLAgxH0OXWEBT0s8FI+Zeyk78Fe+g+/md8C2efsT5bB
VdeUPL3YqkZIcGs+6cM08XnXD/BiL8uqslJRGu4e71KZEqPWmbfwSGYh97Vdv6+4
SogUGqMy1XmzDtapNVOCvMbLecd8iwD8wJ9ZQi3qh7ezB3QX8FEh1DCUN4ED1j9H
0JDfCRup9ttvfcZ2PgvRwzwofFmNQxkGvurnMau1V7c6tulnVbMyZuHSZ8xTnv/4
gt3vtglCOrmEs5u1Ik5yXCZzi+8LqcwG4qp3UbbPBWRvKNWAs6nJOPg+B0U1QkBD
c9+MF31wcazK313BTRu+G1j5m4dSIrPywkPG5TbVNcR7sa/9hXssD4NoNF7And3/
DCwsWOlZ5ib9FRWPuV16OCFIazWOkjs+2AjVGOKTPzNJTx7CC8mbLRX8uyn9JV/M
GH0Fks+4HG0DauEM1qXzeAVi5hkflPgznrfF0JefMefeGBzs97JGl/YwKUEnyxDH
zxNXjFTiYS+UXoWYykMV6YLjUbIQxOMUjpogDf5CTIr+nh9UWoQ2tjdSU2AzpzHF
Sj4Z3RXabUJm0xti+2BQ+XWg2lKwmDjcsA4itUQtK3GoIpy/tn53yiUf0IMu2esJ
CXORVNi6gRYKhvtKtHV55WWaFJkzSzGtzphrDwxlt5CmostTKex8K+RdWKAHSiym
dTLB+51zvFaJY5uvpyC92V+QKNKJR7ACof2FlTvzpsFjjmBgJ4bzx2+riW8fD2xv
4FCeHSO3z8LR+6AUUnKjdYe1XoeSqsjg8ebeaqLWooD+VAwhu5zNWL/6cVCvIQl0
d6A2Nt+keEzJBlLLJrJbWXNieBkKYZH7frS9KxUp8EuUBBzE2eGhYK8ErMi64UH6
3rFzEOr1tfN2NSFnU1mmvgXGYmNiox2X6tRsUn0eBoanau3ww2mpDpn+tskErdDA
ZYRfmlZ/hy4Dvgsu2b2qIpKcZo4tvX2VuKVIjTbboql7nq0kMa2L7iePdX/a9+8Y
9jx7y7IrF1NmswLp5IOauuj8SJqU8vjjJ86w9MkjcvgMVJSpcusy/f1Jfl/jzIyw
U5FRJwhDdEUdoQdC8C8s1yfjilsPosVLnXYGOAvAXcvTiHCFc4w+52Hos0cihQhx
d2NuGW23HIGSirBKRxAj+0L5YRnVlcTS0wdggqfh/JnHqdiGWOd1tAC7Q8vddjRJ
VDWGDMR1LosXBg38EcPeAZV+7AdzZhOBweqwROmAtbnTC43+BPl46vTsbKhWkdFP
EUUI3HikPY+5MeZPR7UBTaX1WOFkXplI1vl+ke7LVrcjn8dOZVem1bsbd0fqyLxj
6clriQXgOyp0/1xoG+c57PpyAz7opth0H/XCjt2pnPkbF1lgYcV5p/BqVhtaAeLw
8TgOB4UMuzGp3b0B/4l5SlrDj2rO2iAVDvA9+XgutyW1I4zXVSgsD02sjEd5woqG
cXH8FzY3lhSMe4KL2yYXUt3Cucyqpv7VoPZ97mgwINZy7MhVCGQuKfpj7zULhbJz
sDVcb6KqBebnHWQ7UsXC351RnSodDZqvtUxd1sQr6Udg0Rk6UoJKqGV9YjqM3RAB
TzTfEtT8OAOMeL4W3eSe7Hnw1eKETYFa2Vt2JS6LPkZ24C7/aXOA73H87cm23huN
mgqsUAGO9U2GgEaCQI1g5OlIjWCMe2Bh4Cuf2O7We0uT8MfNcKS63ZeaiDAMVEMM
2/m6dYKHMd0E1j0OKP0BQ0V8JLajhpalNuo2ATY+Rl44gnNzUhvHU9eMnpZmnD8u
iKt85WQ7W1W6TxRM8iVtaVNpBJ3Pxdhm5GxkLHPeX1YIZxI+tEWYxrDfF8RMGnIm
Uay4VAIv2aLcj/49iYFWKut04IzfZluij33bVvmK0xFgaSOoOSSBrGDjjvSoEMzE
w2+cijUA/l8xSA/TE9bkQjc/sZt2Qyl6s+jiiZ2tRbpOOWetXmPJPROTH+xN1/gE
S4HRawUn47JJ84dZCScaleohmJvLou53SmJo98wkuEknMctnolDHZlyVdZGT1GHT
9Qed4ZmSKlmM4cA2R1eHQ4ZOh9r+CDUkOlPuXHiSayCzeHJ0lauTTWv9pbYTNaRN
uTNHc3+FqjH9TRKpxe+NVrOqq0fxcL6PQt08xzwhf/7LVzGSnIcTrtqScCQII99x
n8qIWi4paKsJBi1cTpj0GUCx9sbTmjWOjw0bSfwaBsUzq0Vrorv6bL2/Pi54elRI
ScfIFgGCPO7E6VExPTVPPvWdUuDGf3cpSZIFVmifz2Ws3r2sPWhYSZbc67N/nNn4
s6PU0S5HdAIxM2T97AwaPiljldFAHwlV4DTIa35JR+l8RSM5HQ3ySo4IbBztNc3C
fpfxM0NaQsKyvabGgBPxOHPaP8nguVsRxZSBKb2/DY9L9/blxUqySXvysxzLCx27
MJzf6G1SJ1PhbG4w5nXR/1e9nRdOPEaFFfEMEBjbq2OXkgmhR9T6aZMpJx/H0SGH
FDFkojz6KsqEaFaCR0O0Dbxrxy3JIJOidXmR/GYM2GLJEqC2NYVL+oukm6x2exot
UyexpUemY7ikiSZLKt+5/mr1YaMNCPgrs1PhAcBFYF1kqDDDxzIunk2cHFHeFKP1
L+QPcrpBzkNSCvqPcBwsI4nRMwUtUThpBy67uPmgonaCK+iUdJ7RZfuugdrVZRoG
P38WOy47e9+Kn5YilPob4WhcMWx348T9e9VCANyx36xOAigxZ3YI9ib7JNOQa0le
21yGx0TzLBbhYiE9RionRr6D5dRiqzlG4ngBTaiJt/x24qEobw2aRwiFtXGJr6R0
T4+8srGKdo+BEC82P8RPJmhbESAGfuSJgW2kB+EbbYg2sUTB2+dmNoEO8wD7MPKz
IjfGk30hkUzKtdYy8jqLIK2objSD1C/JKb2132JOWv8P5p2FNtSMh5v7iECRZJ/c
XPJOnNC2qLsuazqrROiABEIexsO+2F4vuBPZV9P5dsJEv5+hdGWHnoZvVhnt7UOp
h92ZVFkhzHqGl55Dp58ksk9wE3yztLEZhM4FyO+PJQYwZacfuOvT5+EHElBWqFm5
JvSRdt/w4kh8Ag6aopBH8suWNVTjm5C2Ja0O0O9voVcZkcpesYgMhcLPFGzLnvES
bqG9PJ9XZcF7jBAK0zlF8LIA9mymffHQk2esJzpj0jCHVusR/nHgv5RnOUXmbQRr
IO8gs2DnoBsOGbtnK5Du1AcidHCyIKZL8CSMn5nL/HmT/yDH5IIhy4/7bErVOF0s
Sd7LwrlUALBTRAoPuPstphAo7wos6G6gy++L4PgwvL/WsN0DxsOH4zenOs8bALBX
GVb9JxBZFaR4B/pb+5DD3KTMitLjk6SpC6rhh/skbJu5SmvMGvI25sti/BgxGpw4
ucoLvN85jlhnrW30CF/bFazFHMEHC7+m7H5THhRdbr0viFgcEPsi+wpYXRjrJCxa
tUa3BWnRs3sHTcyTiVSuhyeIroT0Z+VLL15YALGxnQgiN14gRKmxFgqpfxZX7kS1
YNZE6qwCqt0RPON3O00FPvdPMuUR3gMVlqIHvT0dz4+Wi61WB3ClMWeqGwb8vpGS
NH7VLUdjzrAYcmDW4NDjkMVJe1pbd+AicUWlxtvvM+4ehJHj4qjt2XfQw3JctJIb
JMua9NXqASmrlJTkVgXjyOyxDOyCSPh4FIdQo0zeDivlmOz+IVN0UWkbQM+echKl
bVffLGjlMtQOwGpj7FTNl+CvpWnDxDmvmlEDbKcHOS0GrUl+1lNd9u/b6EqozWh+
VPFJ6flPo/nHN32JK5tyjD5xUU7R/ENCkCRPN8yBIpKhyXIxNxtADxjRAJBV1xhS
4yRAJjqc9DNsv2WXZoItBRsfHucTGbgv/SothVce2hU=
`protect END_PROTECTED
