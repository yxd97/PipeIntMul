`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvl05MoGtlzY4fhg4S3P3IxzIDYI9ha6WWpj7yk0brpQb2vD+jRy6UyzrdxQsDaa
G+Pb2EviFHe5jsbJ6q83uiOxz/coUHfYmP6lrLR5d9L/Jv2DvMFpBV7QDpNZSOw2
y2YgaBn5+qojV8mlAfkZjZqZYW5IMu+T9Hj4z0LPAqNG8vcHLVTFYfK4c1coLirL
RM0P3wu26YK0iQntUNBUYB0zwUjVVV9NCZGSETEnQjsyt2LhUjgvf9Hv0fcCua8L
`protect END_PROTECTED
