`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
++IOTXsz8+TV2zvTxIBFSDVboycpc/EmF68+Lq+xadyTXIuNS3g5N9da7Ev4qXxI
I+dHXNpVH6MKbKeDfI6WsKYwoNgDW9eMr7a2VtptyrUPZIYvzjj/UMNEhWtG/Yyv
R0xzWAMqOsH/sAW9PhfSzE5JVzZI2izrH/SA7zDnaqnzPVE7yKX1VttyN+FuF0di
dPQPtC5zey/UHVq/0+HvbSbWWK2GEaEP679u7q4KmEZkcEqCZ+XJFpM2XXywRDZg
BEb2Wv7d8Dm5XpvzOhShH0+h5FsFNsNkpH/u+yBlo+CaqYWLS+P4axaZwalxjHyq
ZVxow8Z4oTR8ZkkQBcLbTh1WqPGlGj5Fl3hlVINfrBqAABG39vj9bOt5+GlaM55n
FiJP3HP/xkqHIZlb1vgGJ3Dl2TFQqLa85MUr3leMUjFDXrpBAEEzQzLEPiKl/7Fm
lFZKE5qqx66/x+cOZCpQOpiK2N9vF4NT/VoeAH8QRFPO/eupJR/hoXAV+pZq62rB
fSPxBkDgGTTE0w09Y3wLtisrV4DksZVuXBDOHjcwrAauFgYEYdhjWBQBAo5p2cnt
dbqIefqq5WHBxuYWgjDlDw==
`protect END_PROTECTED
