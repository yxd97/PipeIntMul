`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aiYLLAsiLo9hgIjqI1TG1nKJLoRJlAfgSZWxIc7h2SBmPKE+08d4M0Fr2w9GnVyl
jWkq4wgy9QZkICtDdVJG1oYUOYi70FVfT4z+FvQMxoGDfTfkqgYHAHjHhVqwkOgN
RSDf/YQwqWNcEELMh2lisaSwo7vi+yXv5Z9qb3wcV4OktG2yit5uUngnWrIx1B1w
TgEk9TabTsKC/84bBkLK1j+hGzCPRzTpj7EljMQJP896clpkiIlB1sgT+rWBkZzl
i7HTMiGOxxr+lZGQ6T/ivCd7z/0I08mBuOEkfPiV3k8Lqnzf8QzE+E5gx0BCVjYv
g3PhLB0zf6IsKi1fBamKiVUevYfC4z+X8Duh6lakecxg7Kax09SMBMR+KVWc4b3u
r2fkEVTpAiBLxbere7rgqwyeRwybSQCLgJNnEUaspXXTvjgZhXP0qoeGe1rnijaA
o4Pcb39Q2hTlSr1IImUCJLmIP4C4byJF8A/RFPCX1fZ+NRL8UucVzEP0fuKqUFOA
67QW0PbC040nzVhIznmKegGl106sMn9jTzV07w3fQqk2WEiwwlOWCRK1Y9pSL3np
QVLn04ANzQm3fKACQjZCsMscEV6A56bn/mpct0QORKXE1YWVpInF+bdWeB5Cvm9+
wa+Pfomlv3GoReNXFrTyAWfqZKmRkYZXCyj3ZCGD5h7tXvDEsQSUZaiZnNJRwFn8
Bpx4Bq7VVvz1VEttK+gRqvzSR6qJhHoxTeSoxIZHiTXnY7cbSzmnRT3ywA5W8Db0
Zw2uR9FNT9vOSJkyJGwOV9BdA3TumKYjUwz59yltk/y+HBH3zO+ALpkITQgNLZ+n
eWH+9eQ9xM+rlA9irPNSGic7viw2gbcYNDWWYZAUy/8PK6WmE+fiJrZ15i/ed4cq
7IjJIym8UcYIdu4qq42jbaZuAjF4uPpQJR5VsvKwDqSngko4FbyFnI03DTDFwDUc
7xm02PO2GoeQXjgrFQmfMt7RS0NscpxcmNvl0IgoLEnXCoY/oQdQgHptYQYV5ZLH
Gz2OESCL8dMI9V8z//4mhrYZd+Ww/RNpzAaVU7eCpytCFa4Rk1U0ZVa3ZLD/i04M
N4hdeTCz8I+hWUDYWb7zCOQDs0AtTSNSLyBcjO8Sx1HvkQBJqxPvYghAqAv4UJmL
12XYHN+xQtBbOPoYydwRXyYogTyLPAnyWST3uvfj66q8zFc5YL3swmdiJGHrKTAU
G4SllrqrYsevcAqWYHQ1iqez1KiP/1rElct1GNa24Sl40tmcLoZufJ3d/Il0jsif
UctPFOUca0y+qqdVRZFSYwo8VaZ4C3kS7TLT4oi0eMftosLCVkxuSRMlRbti+lKl
4MmMNcHdZa07ZHV3+mx2pJ+7IT46bBjyGQl2cukD7SnotYfSs2hP/lqxDm4ghCZV
OeYpBiwvgzzfDPH1eqWfZogQca+7l+Nuu0LTkmLiyzlVV9oJ1JRGkoyG580KQE1w
vQgeXnhaMmV63NA5AgIymTtejw/HGVDMKu8ky2aug05xYEsI6U2IhhMB0znfoHOP
TvKugcgcMa3e/4tB1ooO77R/9B6NXCoAJO+XJl35PGYRsnUNhxgDfQwfQe6Eu/Dc
X/4b1qPbH+fOR72YdWdlHkmPk4J17ClGxtGLE7ofsjLsEWiy/pskDQYql5t97K1D
j1cFABq7dN2utaHvqRLucIRqlksoClvwpL93XDNgr+3omHNMiQkcIzqw1Cf9BvNG
V54re4HgwJnWuf146W+ZG6UaugmYl33YQuKgltBn3uSYkHcvdI9+q8lB6sm/wU78
N0P7kcmYOdHlhjN0RX0AebUzJ7P9XqZGoA19f0PNdbGKj3+gfq8x/U3vszZepTvg
Iq5isMsjHhBtkRlnLr7IhKZ53MyWKWNQeF/Libq1pcIwsCKujXfmlK3T+MVSQf9g
PnmvRk2Tityg92ONUUM6JY3tEMcbF2S2RqhXr1ztc790TkQXXzguL3oRBotmpVDI
Al+1uNfHc+2TZfP9XGyWdYFeGd+MPHm7FMJ/3HXPMAp2A+b8tVZB5pb1JI3V5KU1
GrI2SFWVMq0/z86AmOP0H/PzWQH9udvqHaFpG0eDW0/Pob650gfqpKOaRIjY85wr
k3QKdLpAtPNSlwPDkpZoP0v1UY2X788GnLUo2vZTDQzlJWNOS6gJJZ/2/ehpmZmE
GhSBBqhDOCU34pSOX9mr93qzcYq+9HY1FukCa/aYkudkr5Uu1YUtutvRnQIzVzsT
ASW25ILOch/wC1EC5bethRx612aCo/PVgeIKMuMl7CABrssrVFc149HLy1TL/hnb
8wOBc7E96hhLPHxleE2u4Bvc8DCk/j/V70zVbm8sv3hefEYqWqoPZBrlJQhJmFob
QpZfC/+zlgO2lZtiwy0zVQ9LpcoDnWJN9TPexXTQ3dgestujCxYBneyKj2XSIwYt
lDs6iT6mCL9EAEzF3zA0JOvLW/pLBF9zUu4uJ6HC6DVtSbfdMAd5mWHFS5gH/Zqu
oMNJUBjIeYsqoW6hXNa8snlyuSHETn4+KIrurFXe4dMr2gE5wYPjp0uwZu+DeY58
JNZEa2gihMorOnN7DKuTk1vmVcrmFm2Zqrf870CeqT2T2HS4+oK6y1yuH9RKdeuu
CytQ8CgevfAXcDgR8WttZwN0I6KJBoAXXLBUjaa1DufH1sBr9Vn2JzMsUk0dqm7z
33wHzsnYYK4CS9KBm4MK69HyOb3egPO6Eio9P4wXmJZ94NLcZY1B7Q5+RzS3MFV4
H4gD0SMat+c6yzZikPFnKvGN53Cyg2O363PR7S0d65K3Y5Q+A0+2YkckQNxjYqqj
0ZTnTnzB8eeUxHQFczyx36A7nTj6eV8DjH6rMnkveGbPWDJb4O9FDWdaXSOBurQ8
XnPEDEFiI5ZLdP49gA49FDwGw32raS7rCjpqwUCDu2wqQgInbO3DPZx1fuWfs8iu
w+WO0BycfS3nskKuOqi7EBgLauLJdw+52umu/1zRV2ZvBcMGFDzeBIFx7yls9Lbz
A7U/CVAEKNXfnqzwdX54M2tR6zlSRKJYd8Dk2xhe2DjIenVklLfvOHSynMvIErV8
MAyrxHf10/aSPPcTIVghqiG3563vpNkmrYoZD2NtLk1j6EPQfE8p5Yz3RKnjbzZq
0ntb/5W8SpCpchEP+TlW3eECHN/kLMdBId4pjx04crATrYAGCvOBS2ompUNDx1AO
7/iN6YWfGuQo/oDIPCIvS6zAMp629R6lAbHsAy4PKvvSWKlp54QZdNesUuUlsVmO
rhvS+dlPoMOUPewGkiZdUJo206B2yBbLjvCQPcPa/f4FgYiLKVMO+/moA0DcdcF1
CAr5J2Nw+Zgwpnm8sGcMPfGm3IZw4nb0lC/CYpGoIM9kwfeTHOBaZ2CRzjr0zgpL
hInVRYcmql+IsyJ+/nHPVNcFKFZnvTmDNy6TSj8KPFQ77nlKJxS1YgiKhFFOhV74
1DXCF1JmlUTPYDu1zLQ+ohx/emrgcLD+YkdtuvQMn9OeXKiSGDTEl0Uqp3dJ7y66
rakwISaHgkgMmy7YB8lGb+OO8bHpuJF+vyPtsbmujWBRMfNDCUyty980EnQ+zPGE
/6bWxs3rcTPASdBoCodmAAaf/suJ0VDLxn9w22agde2WoABgxU/dy2YdyqfRHCbE
Cfffp44KCzQEsis5OCCYNqZyicDi7rhdaWDMLnd3Ga22rfpbUYD+dgfHFbDL6C1g
E7I2+M2nTLGSYfmAOHMGHK0hTMyeQXIkEHFGgOK5uNuGj9v9sLu/xjpZLl/l0ZT3
48wCK/Bk/MAn0DtYy6KDvW8R0NJWNO5M2OREe6azbNAZHTU8yvyzY71qlSiEAwA1
IEiNOCwnsLqK9YIzLgGxLLmnGFMQYpqkxv8EzEVOphfi8yLG9h5EjX4WvsD6EBzC
do1QPmSpV/3/1MZxGTrRKnWqGRlhDV1a0wWwObW+JECim7AtFcbwdVGDPkwn5np8
K0WelfpzYFGAMTKlQ//9L6tLWv5CwWsy8hBAHs27fy1SSnv26WWaRsWpBpkEaxTh
2KfkgPf/us+jtG95JoBf/sXh4ZZv7Lzjs+OcB4nnj6CIyQG37v77Y751RVvytlZi
3lnlct9f9SM5wUn+fyV4NWmOsdwVKarqx12jAUSmbLbKQb8NSOMZbuUZWxC3dyt7
ZfVAUzp4nNd56kkdViMlfIRU3zytx6ydPSU/ocQV5P+1LLNZepA+nshMZpGzzPcc
Bd7rBwIOU5lTwME35cSegpRe0qvj7H1L6ByJJzOm+s+OoM6hblbQbT8Q5+dd583h
vfNW1upYMq7877c9jkk91nVt4PcHrrkFaV0+ArAmuk0+Kh0JxtRJ3laMJi+p31rf
gxU+3g2FTKC6GXaR7lPwwCwQcUPpWpqC1uCfqCUjgEcSWpa+tNA5xHZ5m/uT4Re9
1BHA7Ydg48xkTZ22LIM9+WWM8ntxiQKzkLUoaemXd39ar5N5QZ7vnj9kQrnwTdL8
hs6ypnlSW5Dt8FtRnHnhRY7JkqyioqUxuQEn5N2q7l2CE/fs4r+ZqwsQQ/fhvcOs
NTxjx1dje4CB2mcEyFQd5JZNj0uPi6fzxtaXMU5xoI74NLHWcIrktDrEwbMglk/b
4otNmRbuoFn8V30+r6fPzs5pEZ7sULkMsRHgdkHRfx9fVMcQ9BPKCcwCVE5h2fWA
Cb+ygE9Ep8LU3ztiPhDWalPoft0EHbukenRodwP+My2eLG+pzHl7g8wvaJd22NAH
Z30Q2h9edlq3Q/hCxMPgI2Rk+ckIvc4OxPUlkhLoIuzrBSGKMgclK1FWP4zkOa4U
D7UOWWMqWI5sJp3Wgympfoj/JE/Z1RM99+akA270//dStizPTzTwzuse1fWpo5dl
AWB9rvrbyZhfxwn/q/ovmkiMo6Nb6ksTSRmYcMmhYA55YKQseM1irzQwrxkxskDx
kAnv3C4XmJFGCeGC0K9VRoOavSIDQxjub+mfuN3q0Yggehb84tSojSc51qIURJU5
+sAJsVfPjhhaQixMls4d5mFdM9hI9RVRpY3KVfT/fvWduNuI5bFasBZpIJCBOcmv
yf3V6SsRKgwW+9qodVLRoXWmqkw7SgM/ViTehlNeQc25HaJk1i+NjXuZNdBHBLRh
TTJKs8HdV6DqRPAM1Xrrmfyr9HwR63NpKCtkGwaM+c4pxcAjhGoR/VJl6wmlkBL6
2k79AruiPCkdl8chQnYg33SjKKDMRwofo/kO+4uOerlsWqVec4VA2xfAhsnRA7oj
9XV5ktg5jaburx9617hvQ9HKjS3NkI5h3sILioMB+CY9Ssjh1tGO3OHCi2Ai8QbR
rWjeOpHg15lgTvQMkRP+hQBJbIo/JQlrwoRtbnqpZC+r4OOULyvvEsD440Axj2uG
ILVBTF9T8yjCgYmfzJcuH5P5fqMWdjrPvCDeVScv6RNCP0xhYNJnKgokF6mtY5ht
zE14lXEkBm1TLQDhqnqSsZyJ9RdW6muR30QFE805FgDc4vQfqsbr2xm4QqlxozED
SBZakDUGJmaIPLLrWkSscgSdafIRHLfIzo/CMP+b3Eok5j3bpAhbN/oTQOKoV1/C
1YflefOCal1kbSTY8PnG5M1ScyL+6OwqDRYJYDmDjr0lUyeY0G1LMvuj5rHuposS
WEmOK0jg8aMxVAdWO5B7JNjPorhH5kYP4sm6sz9iWThzkj9oT/2g/ydUZkt8dbQ1
C+X4m5Qx444zSWwPCnho/YGU5WBULQBFuerXXDdeaz3TAlfFunQ2wvzfrIMWdwr6
vqYi+fw76swFW0HDFZf1YYLBqWSFAN9fitcXaLJEx7M/ooamJnN5DLwjtmJdiTWW
2cBus4PKMrE9DLu8tAlQ/P17Ma8Lx6ODVvtAhvx6Gw+J+Jam5xrgI8D2hAvKorvq
0Cl1kMOxDn6+C+UuTeJ2BXtdW9zSo2y4ZPumNfL85cjtCm1UiXA63HmVoYvhOjAo
zk1NIRVL2rWCpMWA0V5WYBHkGO0HvDfSKKC7ked7Nlvz7of0kYbUYws4JDGf4aci
G06y4P/gBon/mpctr0bRkyza4k/4OLn0vuoj82cKQuRK602hiFOZNuXBCMQSGIHI
gM4mSKz7o9+Xw/N9uwL4wI/GnaxiwEfi+0khUsLfihzEVAVn0bxaPzMFwURVr8jh
4PY9Tjq1mHuiijU5U0Ln3O6pKS7oZROTOlVhZpnsIEBRsO8rW0tg0mn68CgsJpsI
ZQvLIiW74q6oSZK6JGbpHHRaS/Ny5t+YZN4AsddUO2MAlDPD5B1SojnpEjOu7ron
I2pNnrZOnLnI3gfpmQICkUW/Ey/Sdi+NdanyxEuaEMxgIh1zRvwZpGNV7adw1K/F
dN56kkv3ImurHGf1RYmxqEuM+6LdpARkQgysdxgo+WXMuOT8zj/RgOZp5waV7yad
tN7nISR9oTNJnP2tbEjdCTzYWOW3iUlm+sFLO7tYwQAEP2A1pTBCLKy94BLT1bXk
S/veTuixaPTUdXk3TBH0/HKZUbvpAAtHULpHnfqGgT3cx0RtB6oVzRtK7UTHFJbX
IycOaDuajBxcsIRnz9YINsh86HAeA1iA5VHn0oVmI9bAE8WjrFLhXhB+avJo+bvR
FKudmH/6itvReljaX/kkBkCvyzK1vKaajf/bDs/A5QEBayzsTtCsDV8RTjUvS8n/
+VNkoeeJ8iir8BjW48klubiL59N2RIoonLwbVBbumyuDeOyv3jlPPDezAdYPcgnL
e+USlcpDRIlNCjckmlRNlSjAnEl1krA9oJCX4002H99huOxpNThmlLNF8drFBpd0
DoKqXhZsTpEwZ29exjpxHczXMz2BErkr19FrtobpEqGiPyGy3zP17/yE1eFkWUds
M0pxs1csPGHMf3zKHfYd5+n2YOs67+A9l2FAhS0yyG+7pztMjW7T1e2rc+npGBgH
1kN1M9i1/yW0P39hj12u38kj3ZOJvsjvYEy9sbryLDPDEXsfLSMvZTRBTW9GXWoI
EnQ3KTK0+1JjGGbKAjayLgK8U6B15k5HE65KrGQ83XPdGRAn1gn3QYA13lTCcsMX
NEMLRYxWUqteblhCzd1SM1w2cG6gm9LwQtgwlP3DzoZ3mDxHQPfgKOTjymsAfhas
s90qa64By+ft/JVvjEjknFcpEA9W08kDPZsEJfdX+azQdoZbz9DtFQPEAyT+YsAe
D53BvfXz5QO+uKqgSxrdGQ80mAJZAA+LkkedEZThrQjPfJhb9YUdU1ol2Do29wwv
mCLnAYhOAyJW9DCYtYnL19uxZ85wkxqcrG6nS7rl0780lIpHBeJ5vK8RoWDBFVrR
IjtjJBer5fkNosVcQpsMABCVaMckabjjUFjOz0lgFFswPkzMFHqQw2Amr5kI9u9Y
LNCKXXMwr43u06IBjnvGSnc5jXiXQ9R9/FIT2iugXwm8rgeIYyCEkD3P8kOF8oCk
850ASSCu2STAiuc1aPsVKg+ie+yOofWZpzUeKhpMlG2i1sIiJUfChq5z6D/eEjCb
lDOwOZAY5nrsKXg+d05LMku6Q9RD1FojzUM/rVWcFj6FjNvMl/SnSNbb4qE5EGZm
O8YNcRKHcvQufffEkCyMVjJngp1SIJyVv2MeWKv9VzXICpqqWxZnMyZ3RJvUDEYI
yRQnuR1B17m9WKapvYce3u4sixb2s+hUJ57PKLCAcVVL0n/gqALt/Zy2BRGH17W/
TgW8aRqIjR9FckgqD18mmmafb8bS16D6qidlYxynGhxJa0FtyrCpnMJ8MD6mjYcp
12uEEPPL52xYzUio1xVwjOpqKP1AuBwprLhow/RbeV/6s7F7RuheLFNWlwkNYWbf
MzPhdbNmSdsw8TRHz4zKOf9fCYETXqeU4TVC+P5qv5pX7aoYMhNm+RtBr1m5rNjM
Nvxz8NSrH0ptocj+Aa9K/VLAg3mqUzbf8wRkZwkdZeIG0oldPrHstiyYpPbriuHR
HAOEWvfX1A2sPt5sv6ajdZBTSqqyjH3lymmUB2DJB/ia/7hBm2fP9uik6AWHZ8go
+HyL1oqIJgd7eG+Yit5J7cHo56DKcIsbYS6CpujEbtHhmTD4CpLvtzhxhUfhOTPE
c+sXOpw4qm1hj5BpN6ze+Q/pUzMXf5jRyFKa6xVZyLssmx276oeHAc83b0rNJnbR
wwIdY1EfvanGTz423+x5hNpWjEri68ZHlkZmQYHyaywLNXJOebLuzsreLYBH/mNB
zHaF6RG2E/5Z+0Jv8dpYVOVC72HXQ2GJmj2Py9/T/upKnZ+jfcNHVrm54ru7w4DT
Frn/kpWwQi1RpFcTeWIJRRE0wA3HHz0P4+NdVkv4HkkzbbPMT0Mp0mjK7YMfqIuR
+PbAGvVJGmJTH2C2FyRpywyrPVYhyG7MyRgn4GRi2kT4BclxU4sSvsCixQ0GiCxk
Zwmy73tjHXssqzUNBxckcQN6OVW+MxrLygwi3iXm0q5aPj4aNAqibP9YWMIr/fU8
sSD8OKw0t+gAsfWB80A6akibwBwoHf354VLJ466hxULkPV9e4OucpTK3XNZqsXO9
Gp2mcOwMXEcSDH7PGalSD4hhHxlqYpy6swVzUVHjr55XvP252N3q4rHlC21qTCs6
jsgIweKjLvqIPkVLAtUfnAWj8nYJg9YoEECgp1MP2IUT+lg7cyvDFa2ic/Ekt0CL
zdgs5nsr6LPjrHAd/k0tGJQFLLPswYnL1gJsmjG+bwzMnN0FuZYUQpvfOLz5N74Q
kvULRKuNskH8d7aFlu5C0TJua+KIdx8zdkrPVlvv5cEB6xKrIdVk27mBwmvR71B3
Lof3UTrNy8VtZ9ay/vOaGXPbsOvBBWDwrhHXEUuJA0gSy0EbrmIExcA8ea2HME2s
MdBjJvEgrtddWU2VdVxGmOgV/GU0+4xV/PSAIEky4KjPVlml5DUoCxABcnclJTVX
4iGYd6CWvJM5UAQ5EuFp1xchfHtt+mJH4G7QjopCl47SxqIAYJaySf7q6w1AodYC
v2gNqnAbP4sblPDGazls33qWEDpkwnXpcllHlowpll0pwuQifNApvn+BJf0rdaRX
YSvk8YS4vmzoxc0ok/SjSVhAXUheTr41S2Bj/7bSOINmsH2Tzyawp1qMWU6YkXfK
fBRK3B0xU2L/OBx9GaNDg/GBBFmdWci/E3oo2YBsmhjJ2nAqboWOiZd7kABA5DEN
vwRj9mdXdQTKlQpqO7OBbX8RjjnG7QTtNsxgoWLzLL7NkaO6O6TSC/8KHZREcmGs
0wj0creFcKPs72wjZ1Ge+sePbGePCuoR2UfCfBaKjiwEKujKGfKCuw4QavHuEFDO
96asFMIBkueAsd1b66X6I6X7HEnherT4+USMAY6AeEqxx1/JhA82BOlhS0Q3b/tL
6vzqAoe3zZZf+/M/Ut1oh5bEvGzIniZd/nDZD/GLRUkiQE9FZWJY5CJ7EMYzaby8
dvzk8vmt2aLPpWBMkXrAEyme7kmIzssJ9Mbi/diZUT3Ph/sdbkFM8qmpoed1EC80
Y3zKRvvS6jHMOb/VVRuMdK0bYR287sP6e3n/Drvq+JFVrg/kVDsJkfjtAOKfvC4s
Hep0DXCt6iWAvKswRuaKx8F7RWCxlEN0vgQ+ULikzfvv4KDB408ZzxLBu0SwN2HT
NGbWLyIGWrYgSHD/wlJzkx45zYYAihLlm+M4mC932lz+9aXb730N3oANMJSY5QeW
VjnRG1BEu1Zea41BTD/skHbey7yMZaTG4NpYIquDC9RgU0+7fY7D8j26MI0s/y3T
7terKJ0ct10rBOnFuzWqbTRzcV0qInxjlv9vjGmtPvGKFWiuTtpUm+vS/u7T+vUD
KnQeWNQAyw6hzO8z7sCotTVh94yueg6bOvMwMoQYdcpAaqw64eOGpAmT2SOdZFiX
rNIbqtiSSf8micHcn/lnqB0CjiPGMKPnHKsq0/ccoyv7ayzZLsLm5kyXV1Hk5JvT
EGrYihPqe4u3YiqBXZUevPZygv72P8VJXUHs8faKU9O1gz/Dvcl2buTRFQ5NoMlw
GJ5Y6+NB93qb/9R6N53YlH+ehPNahqAACvoiiaGydhN+kZrFiJmvsf9rZEtIN2kh
62BNETOoBkMg6DS9nAcZ11qWrFRAsYXaXcviDxGYmwESvSeVpm436m8VjvYBhIxs
VPxQgza+3IH4cuE+u/roKsp+INvpdLLaRuAdt9LyRsztiNFDOsVelJ8WG6VQau3G
fZ78X06HDj6Yw2L2PlLF3SmC/guGwZbJenBLLwyIkPT64IlLol4Lk4aOUigdUs5b
Ogjfxt6xkDfa0sVbykvEF1sFOi66DWBxJOrGyn9XTHWTqC43PUwOMVxVsukApkVD
FdtkH9e4jJi+9Stj51wZKnFZuqC8BA74qDZSos8IZn2bCf1ygUUABbxxRkIBTOpl
aAVNN9zgsaRxn4Y4RhAbSmeTsU0WHaNWVepr2rhOT+1jlZ+0fOJ8EoOd5AqxKdRd
viUekkdtoWHvBBwKMC/IJycp6irVxpuQCNh3gd+BuErGmLUmmHzxPt1FQrO+EG+n
t+z9NLr0+Y0QFpGotL7TiyVEoGFIx3gwupxiGW8FKcqwmfkUEVVIk2feDTER+Frp
DDu0WnDtogKUGwQBEeMQPm/ldBPhUA4IWEDE5sJF5hv2iW3+q+V0WAbmh1HHVnen
vSfnokus/GEMvSz/MBDjC9nXGWIpGZX2Naujse+K7MfhwOkuGOzJI/E3JnwrRPZu
I+5Ye2fTpbjZwqaE4zUmWgfrVYz2QDOLdB8TdjbHld6ofUgTE3WWry+34+nrFDKI
Qy4T0srAS8Qo5h+CxiJ+ck9Bw7HDCckAK6uisv1f5a+ry37C4D1pbSfrmAHtrMc1
4fn/7Ou/M5zDRjIHgLIu24m0TduZ01JAoxJa6BRMIH/4P5FOC/Mvt5UzVZo3y5/a
XiqbchUiJU6FDDXeHbl58Bl/JFiW77vkpy1wb+VkuvH6XQ3LBTZk7m/c93qrGj4H
dml1+Zm/GTuUO6Z6JeainaieV5LFTmY0YjBmD+23+UIUIqQNxCyzXBhC+gjoVmeM
+1n2f+W0Sfs8DgXNg4fMumxBhViVZOvhZbONlxsk1Z8bUpMBYH1C+0TzszZ8K+4j
V3GnqpRAXMYddpRmO4PIOcxD7Iu+1avobSKbIEJcUq0z+JdiJy5xXmx0QUtBaDkf
JQ8RYW8/1LspYxNFzQgqXa967xq5eKui6GFczigXEVIfpRcXXCg/cSYKgwGQ+TGh
V0FQA6gcf5MxsiN+V/JjYrq85v1hMW6upKSmyWNCGZ+GSWqJiixZDtoUbWYj0l6C
Ca4eLIZuPmDu/IM0UM1i4NsWnHqaVFRjqVc/77wK3XJuXa507PCILVf99XJjIOyM
yQ0BxKboDJga5L+Zjn7PGVItlOEdE0+PsI65ZvllwC99GgZetanF9NwTdhRb3Ilj
JMCLd7lvrBzbaR3IyBnsKtygEnWfERErRLFKCwtfDMiXxlplFdzcpY/CbBBU4rfi
UD2HPyiRl3MM6Gjm16Pc2MiGNNwa3756FvHbaJkXhym/gmw1rAzExxCFZPVIMT82
X2fXEOWriSGu5D9AM5sxtAkY+ikAmcreMIh6fn9WkagUEgGznyX2/8whAM1lxZB+
lGYbQQJJ9oHHHKN2xUuH4NHd/vaqkXZExKWZMcxyAIww+1keZYQ/WjPz+BJ9C4t8
ErX2Vd/cEM85sf77lmExxRR8TSe9nhQRs2i1KZdbMEaaobLt5fxS/k69fGvFOt3L
CqsnwSRklMYBbiT/M/xfGzDhZaG3Jf4keogs587C9W/976DaKnWT/9WVr99qR5gK
G/2zA3GoeMooB1ANjsufUiurklJOVy3hx3BCk+yM7mKZdMqLiCtZJX6tJuAzdZ/n
+V7RviNC92eI5pNqAT7iX68jGAW3sW1qsPDs43E2Xd2IJtSAetHHvM9liC6ufw/C
XdjCAU7NUonjPvAmL6ruJSKX8OytbQoCgo63Hzfe2Y+bFXIqfpHiie40H5qXcnm1
Sdqq6uv52Na97hhqZVAMgojCoNjx6Fvok3qk+E44du4b0qNgSVRNE3w7Lo5bbp38
IhF87VMZqcVo+lMEaeyDNhc2jrV0BnrjlvAK3bGfVJikrfZgzrxdDlKN2DBhdPtc
HsQPyhiYTbTfUDRgNOcfiVv4hed+v3tzOihuFZiUopFZ/DlERv19hqGPZZM+E+RW
uDa/GMBkldBbl1GoRnciwoPIDM0PGL2I4y83trYWgtPxRVgmkuaKMkSz1ZumAjrS
4t5I7W5E0pvRtJj9htMmfiNVCVMMKb0QrJyfEufjvmDgMkdcv7F2fLhKOAXHEyxs
r9+g13P3ZDBqC9MRvWMvrvrJsSiS4ukuVVy8dfXIYAr+YdfCQsD5eEI4FOmAab91
66nady6vtBLH9Oc9j0wzQDRiZZZzd/t5T+QENQDoQUCvrQr5MkdUoZruiEbMXP6P
5UNumIsFJ/hFdHwXISM/SI64eFC2v+TAckewwDbAcuM2MrLRf3wHMjeYuqzky3py
detp8FOicG70ZIPm02os43wayBvdbRgXKu0wqr98JMping1EJO02d5aieoA+l+FT
h+EMEbBP6bE4u+nyhBoMw4GfEVOBGiMQloai21+2SihF/4ysUwnRRW2x7hpwrq9+
vtaLYEAIZ/kNHSyZY5mvwBu9BI24pQK2a49YgIrbU8iowErZNIJRBPL6ORuPJDes
v5Z12G3QYH+BxDHIgxKNFYPueTW5GqI1RlfP5dfakYQGnDcFDuoj5YD/U4Tj2LUq
bl+Jw3dV0SmZp8PJLAuURe8Zn7GL5sDoWEfy7yRUL4RrNt1Sglb9fO0wefVxo6ig
oRPPMfGErKgpWXoovGZIRJ7E66XaHTgyTOIqham3YwAOxrHpP0gRN9wJdasMZ2Dv
B+ktolzizUxdbvlYIxS8yKrYwki10WAm1XrrDnmlHWD5sq1X4lMkHpDbfjtv9139
mSnxHQyLS9HFqv6cGzfqdpEGXZRjYztc+Lk9JPp54x/EwgCvi12uSUG9lRSTcvHC
EC6PPlaSnx29pSQhr2uC+W3++SCdE2VN7cjG93h2w/9tCYn0Rr6XgYMXYMS8jZ5V
YLVAk4GYOQMRXeQIjPuLHzu8BAqpu7lLR1F2z9mOiYOF71gWA6+Ktx98kShZQNN7
NdJLJGt8j6PKAU9m66UJcJoI9xbvHhEFVAtE7NShoY0e/mjRR+O1zJbrqt4504G6
O9F7z5zx7U0pbD/ZnMO/Wgw+6A5ZxhD79NZyISSz+LrgxebAg/wMubsFs9af6NaF
kNAWsbcG2X8GFVrdHPntKMCyHS3B4j+wmdwkDA/4B5m1Lt2G369cwF/fDZ4FoD2D
w3LdDJtgEkekSLNIEJfuPXNI/B6upm+7ZYPsmkbHL6Rie2ukxMB1eQOH0KbLH6+X
0CuqnzNBHvNpsenYiOXIE+2/HkGrBAQq8wHaIk+CWoYOXdGR/WqF6WCZPbxA1KU8
cGBjYh2XWuAfQB3Nsc5hwbxhUBkXFc4dQTFPRZFcNKXc8O24n2aJj81mlSndSD7r
qP599if1Xy7Zhjz8Y52NUCL2UsauFQa/sFTcfJCthpnaH8e2+TRU7qfhdPqFrZ52
pDC6FRKkL6fRNR4zIn6Qklul9NpAqnYTHqaZWZtVQzNtVOsUTu3Sy/ov3s1FgiQc
RQB621n9cG0Lz6KAnbJfdOwuq5dTcMPDCTX26HB6wgaxGDkfm3HCUVFeRBrfFOMs
UyZgybN1PTqkwORP5sNIcJrhyBhv4xvdI1voVqAvRELdLVDyFJpCdH3gNc7piQMi
mBWtUNN5BU9tDLiD+EReiLmCTTg7Pz4QchXx1s+qlbDGVRjZzg+eZh5VCondYb0j
KsQLbGeBQJrus7ktCrNqeOXd34RDud5yIbcJEaHT3sZwJW3zPZktC7yMxWQb+mFT
Arc09zi5TvRDoOMKHDmuwD6MsdniN114pl42CsKPlvXATp+PxT4DVqGRgDL6UVQM
ss8F8flD1LBDb0TOUEeTsK/hAFd0HTqYycn/qeVZok72zAnu5jbOkR2RK7TB0u9T
/e8/JB8F/NK5WSEYwgMavJpsgQUHWmfKnkmaHQR+ZPA1eoM3kO//OFiB4Y1tCJnW
78BhL+a8W2kc9XxlApuunQQXUW9vUceDVwHM+QBSlo2kLFcZkPgDZd7LKyKJWPZa
uIrOoODqgjvACtbT5pyj6NEXtHucsFPfjyRfPxn5NypUX56tVfxbvg5Xo+tr6nBr
hMRdTT9DkRgF+E7ilVywaja0ClDLj6Lm+2fbzAW3u+GoD/pt86o2WMrOllcq5kcf
QuCHujbn0WW5uOjppITGkvy8CnQLKaW16gWx8BD66gE5gwsxN4i6lxAayRBLpOgk
0A9xquEdJDFtfE4zZbOM1Vl3CZ8ZQCftTaDOPd0EMTbI0LmSAUHS/HK/qDoodc8H
QkohXOX52dpbXadY7auWnVWlxDGPxOYwdjaRIEvJt3uI+VqwWpHyQ2vHOR4V954b
BucY69IJKDVAn60CLBaLeJpDmM/q3wOAe21orUq3DU5uQUL5UoBW/ucn2hdO69Ci
fjEpNRrrjn2K/AisjWCNYvLmbsLfEooscJmLDNC5Qlv5weIougDR9tx8nMlcBDfQ
PGtupGYj3uX+uG1ySo6dy/7Oqv2jY7Df6ZzT2o/xGVerhMEO1+3Nk1Hxjz1lwKmt
k1lQQCcZ+T9XXz8PQb/ZSpEFpUa6xF/PyRIHSMAwQiA+zVb1TPQhc+zYEVhVQ6i5
qO/Vl/6TaKtgppYmrMxyJ5PUyyGiwEaLD3NRd72kzZf5Z068R0eSKntSha1bxgrD
igqe/GukUdczs8O6yl/fOHuaEh4f9NJ4eJ5zNRD/LsbzLLg3234pWJhAxD6xBAXv
kf/vlq7qkq/I0xCREzYNcAdfEk2QbY9a0w/prcZt2/AFyS4JI55zrpOuKQNPLSG0
AlJm2Yb7iCNRvvqXP5r7D0+WouY60t5mHmIXoh6BTwWDVfTdGulSbbCZCcrbcAxj
d+elzbEgVPxamtJeZK8E7xTPoSFs7KarWcyeDLCzJA9wEeHEOfEJVOW6exHK7tK7
5XPWTOKqATG4DdnLu/2JJzptmuRouwzInPk2BHxJS2O+cqwbRvY8Zkc+nkeKAL05
VyC33EuNxbfmlkpc8fkqWqZ43D/OZeJIo2lZ5paxhzuotV3LXygOOVQfnIirYp8f
6+jwPNqHX8iROo0SnDCSuWBhdKpNHn6YJPhrsKNS2kJQkt3cbD7jD/1Rlqxf7q2I
TpqOivxqU+O86KOt3OPAcZcFn48FoAuDRyj3oe6N5WuUvOLvKvjvzK1Cqw+pd3Wg
ZW1bOvNJudR2qFGsm2m4ib1S4GWvQtxN6puYb5ABSljpj9h3hDwarp5wqHV2CLbW
Z1E6O8twrbt/4WUBxOavRZu0vVnNT3r80VTVvuvuvc0h+EZpW8WD9+i/EEuQ77LZ
wsyJpKq2giFDAA/ofsaJnbDFYV8AzBEjMBv5SsTXwcmjRC1mU1QOwJ3rAp1ZdV7/
ywBH6N1POCNUUo6eM4Vtk4MrtCs1zh5D5IabXdyPG7C3ONmVVojs6tb5GZytYCrF
OqlHA+M0rfa1oTxkB93WpRQ1e/4chsQ7/3xTKiA4ftRFEj2MiLiUn/XH1dFqNApl
mxqjCoNqahYEGlt1wH/hO699+uX9Ox+d7bOBHod1bikgYyzFP2jUn5MibVpeHhNC
40fXmubjOWKhrVuq3DFiIByjbeAKsLlciMkXCvT9RNPWdRl9ei8zldHMBTXiueTf
A/UO6yoxroW0Upl74q5969nXUO1o/XSOodlNdfnokjTmEOlRO+wbyBDI6RWXzef8
9JUYid0Ui2zQa2wpg0tlh7YbrCyn9SajjPtSOqqUJKLWYKPDM9AFmszO0aAAoQdC
zi8lM/e+R4M9z5nqOnYndG3T90/zsgOjGBhIvuaoEdpDQp7GDAckIPOZxKOs/7DD
7PdV9owb+0uy8USOKSBfNNCc3tPVsDg7E9nwGL2GSrcZLkN1faOkE10sL0hW7G9h
qbneFAn4c5B1VgFYoQcauWvIflR3MoX3ZfWPujIAoweYE4ZAvyb5gner9xBkIXvC
xxbosvceN7Qsr2PozQJKrUCDP5+lWAF7OAx3cgSf9pIxSdx1XP6RYY98iYDq+CKq
xMt4bBqU4GoPI7E8ZXAtvCWZvclwSwK/wlesKoEIDYWg96RkOwRZ/rq0yNBcb551
bvu/jq1mfCqUaXsg/3F8Dyxnp+uvydJIWa8JlpEjPNvzF4jXxu2pG+5qWAR+/Ba2
Jq8gz5WJw+EvPaobBgSELa2/QnROQqWlMrb0x+JvL2x//EOa/EHHMRWP9RzwRErw
4vluDz/imt67KI44oleVrkyu/FUAB+iVVDZA0AF+8jvh2ealEZP2vAiCFNfFl970
PVF91qQcCZ2pdcZJN69Ts/zbYY9j1s1jdBNmyawPMjKDEPo5aHGG5F6L58kwClNv
CSOaI5fIbvj3+3HxGjbyfRBk9sCm372/iQwlOWbmDus7b7gJaGcZ6PNZaI3gLCXL
y+1V/7ClehYTzsHiKjXt56++FB42hT4ac4GPYT8YYuEALH3VlUckTdrfyjOCiiIq
gDmW9pE4HWEZ0vFY1jy0kxTesB32W6t9kouvOKSDESwkITvPdgQZx6ZEBjRHRD0C
ilZcyODXahZLePSrhmpTP486KBNKQzOSS+fDT4bHD5fJ9JefokYHq7a5zksBfDeX
XjSuky6SS4IqlTsE5XW8uKxhN+HdXxuuc/l/euf9oKQkQYf3tesq/C8hB6VrUiWH
JVEr9EHQe0HAuiehS4tchYF4godlHuvcLQy2FH/YYnVE4hc4Io6G/9M/58DF/rBh
NMRS3DfVDn5s3MTAEw8FOV3uRQR/8XYs42F1dPavY93f6vQeggy+72egbd8x4CHV
Q3ttGH9KkdWX3Gj6H6AafDZ4vFANeHuoqvIW82R4DB1LVonitFliKkfiQMmxMqa5
0lp50jDsTBVxwWLT7fbH41/xDZoY3FqByySPiA56Xa2ux3/ghk0qR+vSVZgNFVI5
oD/TFHpqb1AmUme86uKOzrIi5M2jlYvEnVVkq+/E81iMKisZADI3IV1/WsZqtlGt
HkRMNjE9hdtBQ5Eshun08fp5WReCjBT4iiLRdH1kihiil/dPYvghGjTvCIBcc9EQ
cgNo7+/qFOHUWrqMuRMMv0JjBxDi6kXS7ZOx1j1O/YGPymWBVnhZ2E6Mh3o8AckT
TShm4Imz/fXyRVR7DqiPLQjsi+38JtYfOstOJoJk0qgAe67HUFQk00fSg9801ziY
LEdjr9rAn3X2NL6LQcIMqwZBqNgv3CYiHDyHZ8QSUAiQ8+tiaD+k1XOmq04J05TR
Y8hITGbiGbqcTZ3EkVxI86HzaAQgyJOVjvT40KFnlqVGHkVQ2L0x3fn5mLxn/x6H
LqGjuP/2zyNntwB4LaUZJxMUZqaIZNR5CUP5p0OvKi7Wj2Pv3RfmcGeAj/RjEaUJ
SYPjAxuGa5L57UqGTs14poCbY5uATcPpvJpEe7h1emIajSPcNtAE3amkRTOTrll7
xC0GbSPXeW10xBtdhOGsWB6cQA1Ej09BFN3Au0ExGHAmsidMWsuMtvdkWal4ZpUf
TlfEjsPfu+r97TmLl7Z0oc4HGtXkU1b35w2kGKRXvJRFplvvfFF9Q9+2unk/UJdL
1ouxnPjH7fonTW9x5Hiz6OGwPMyCYub82PNsun0xgBABPxm7vLCrvzIH8xtO7i8A
LSUL5Y/F7wWm28fc5YOBCRN9p3hV9VmPFrYtlHh3dZaafPuEEdFiV193jXT/uL+y
17zIKxelQgTlKSOgeMrtZC0TWMh1SQZYUfgbter2iR4TDPmPWnGh/jHyPokobGjc
epAL+eU9yZ+LCGhBshHKNz28syZJeT/FRg6Xaa/DJKn5IuEqx7Hw9gIfNIZ48+br
HgmvhwlQ/LSornqDchdXN71ilvhGfDzok2QIEoxkOauk7L6OYbtKLQu266w/AA0A
zU3HwvZMbxdPN4u0V+2S1dVR5TIfIcyLTRNgs0blFIDL75fzrodhWWKdgB7Ul+Y/
/Oq00dYrp15j1qF7scEvnAsyKHnHzGDsllWWjAi73UzG5fBRcq72x+IU3cpWkNXy
GP2JvYzaJBIRt9s2bxiDhj33mE3yx6TAjsJEUsSFQDavmkDhkoKtKeb34/jlUlqP
iVUy9Cj0g5uaybQuHTp0IhpC8mkWyr8MjoUM47IhLUuLiyK+OppY79RBap39I6P9
9BPQW+dX06ARjVW8hoHUkMyY0tkspSFHyr7W0eFL6EUvXv1T3noqS6yUdmSkwnCV
BsyZaqfAdJt7C6DQmZw2Q14K3+tCz/Ay7jVH3Kvp/eyKuZosidV1zoWxQTkiqM3u
FuhkKsI9L7x3pA8pvcQ66h6ePgA6QLkmYEC6yguB1SJROsKbNlv+6vXmLLAYmyF/
LMI02iDt1VvVYT7sE4EVf4nHvAVWwuV9Dq64IX75vmUMUTulrB4lpO58kg0YZZu9
w4Krx9kbTA1lrI0qCjGXDH/BYLB2crylR9xkSFQZJP3RUcbYzDb4bxkJhCpAnSWI
yKVby+bxc5sFfW8mugDYm01H8bfaiWHGCM0JONpCxvSp+y5WHwFZuscJ4yZ/ARj2
z6nSA+C7ChXRDknY2krEIRl8CAwg6DhYaqdAuAcsIYy8+5qC6TPkzK1S0WJgi3tR
dpCoR0Dg+fgcoB6NnlhlYGizJZ5qyEbeEDCdsN40JMrjxOVoi3VKANu5vMsBfX24
Uee6Q4zjLXmKfXEeaSpExz9yqIvt+ikMnUzSAsbaxIW/9TKFLwbsfoWM3yRJILK4
Mzls/5ngrUiTvFEEyq13fuECHlJyYVqp/2FIb9XR8RxpUmbSKyABS6tHNkQXGxzX
LLEtOgRvqDihsux1Hew82Zqp/4JGInyNfJl0tRDr3p6S4DPjBj/dPk75etTVEELy
gHecHEj+0WqIUFb7utRER2YztJQni8P5lKfALHMSJOit9U3Oc0nVY14godF3e1RV
KWBHwFmPai/FDvdmVL2o0UsqkvLATczlYPmZ+75cvO86gjUr1YvnSEmfI927jdaU
GcleLG5xvwbHtlbQ8+bhAVMEOWbiby9fC9AYyH66MV0AAYHz3sKt6HKHUM+UF1jL
e2wjwIJjSe7G6SVEgjxCnIrqf6C3V/nTNjuUjDJmwhydJFsacBIAhooRKzxu71Qc
MnUopu0JWhtccVMEfM1oDzbKc8H/vBvUbxO9c8YSVGImcQmfw5/tZx46Jsgqvv07
xICP6FmNF0plIpCGMdlYeszqXB6b2nBTggma8LLpUJp74ARN1exR1iZu/CeX31WX
YEGBbdH6Gmk+FBYjFBAcUmL/OTg4zKiFSO9LAKjO/s09XTCa7JGkEoeemhMok0FR
czX2WlroaR0pC5gpn+GZogXroSShCKpQfddojo6qFYTw4JXHaBaIh9K2iAZ+nbY/
BR2H+dgvGcCkFfOwPcNNIE/lHrUq2esPnetbCgrcz0q6hOz7j96DP0LKDZ6rlCXF
VGZ8rHZgQ6TuSGhzNt91xk2+AYN+RXqnCa6L/FOpD8Zrpy9ZGbfvYjgy2e2MjSea
s+afJ9Hl4aE5n0yjGfcnrmhK+oXyzd/+ADxJRY4Apisiz2DrGlA5lYyzsugEpYK0
UHf0U/M3oIPiAySMZ1K4Q/kBQjUVpvlJGLMcVVmyyiQGX/wqbHecZhyBkGRNKXP2
YE0PNJecuoPXKADe5G4xqMF+Xt1veePFO/OUXtj/bQ6nHk2EOidQrBdpX8hIpSPH
m60bSFiZt5AEz45bsQtBG0S/kNCETZyvIHJ2lkeklIPQoEuKxO+Vt36jDkU3eVmA
+wruak0139DtpCaB1wshsR/6bFXX/VAVp1zemWlS4YqeU894iOufGc+VnxxMXezA
czkATcKmu/gHJZUwlsSccBbMXG3bjKQf9h14fuvYcNIQ7eZi3vuaCloNSnJJYxVl
RhZUSxf+q9/BEtDVpJq0uJuWmP5o+bY5++l36kGwddfXukFMokek6gIZsK4h9eNr
ty7eGbbYiXOjwsKbUhqh9EL/S8C5T3+Ga1Ldz1vXnec300Q5WS/4Z/63H6zmJigY
1uY0Ob2KZKTsoMP+f/KIUkNL2PvkdBbZg2UsNAflpMwx92iuDkeC/tHt1HAEB7LO
4myrWuGj1Bp2WqfqvHl3RXfO5Fm4TDRiXQi+Gfhv5XOSlhzqsTJ1jTjtJZlMBfhC
2Kvlwdi4axZtgXrQahI6rihBhgRWcKQn1PF1jaS0rf9V6C4wlaIv7XuTdLguOEDK
zI61XI+eBCidcE+ucGBAv0aVoORn8K5wlRnzjShBE3YYk+AYJCFqjJiYf+ReGqTp
Or5qSDlNKJCz+RqodFw/nGBjJhm3CouwPPIQs3hHfhWl3zjx0szT3VYWxMFapqhQ
gSWQAA2aKES48bN4iOeFOzkaMED35m5T/vwBvOSBEB0eQiZjZWpRmjwZ+Qnd1K96
yPMkmYwMpiKdGRopmRC5w29wHBed0paTgb2e3RlAkxRltxb5eCKoaEiXnjJqIFYE
GRxdub0XSOpKKZX5rVREli8XnTxt4y44JSJ2zgbdT91+Op7scrHZ5GWsf/qPeJHl
bFwipO/o4JuDGvqBn5BXdPlFMTryWLrxxkEGUNkSBNU5PlRx19HqnHQY9R2r1aW0
A2r4auNiVigsBeS1wMtzrKPMW5eXQCKnqHB3/eZfa+MERio7NB6qF1rjdbhvHjoD
m5kpdgrV3piQTr5kLpD0B9B27+6gaPkem6mZKnukrYLW+ReqqlJlzsgFACziTmwm
pUSTGLc/rpK/surH3g3yEjpeVSv+9+8BqnhDyWymTXpXEz+4C2rdAKJSq+4CoBAt
UZuJWf+1DIn9rh+YowYZ/t4/7du5UReoaLVnf6VrjxRO2HA+UXM8j/55PwyANBL4
RgMEOX8pl6imGnwn85vQPYn11c4MJov/4zwr8+q9Mw6HQ6W48tO1DUIyotwwDgDG
nRs75PzuXYMoObwLbbKVEFhndKIcNvcB/rdA265scKoCh955oHspgxWZkczl8sy2
ZO6rRYsiSx9kOOGaZaeIIzLSau9KGmHFDQLlLbHJmwHqDaI54vcZEDHhpfeH3k0w
SrDb/XiXykx5sA5NyTgKsch5cjXLcuocQo2cr3DZgexoCfv+EjC1meWd7fUkRwu8
EGSCot6M2wF1mzpbEMPMH4OgZfJlnwn9HHJAz3vg3AAvVKCMZC6gKyqoleGwkSUq
xdU55QH/fIit/J3g/NLivrVQVJQMJ1S41ctlkaS0kDB5W0OPgGeVdigi8vdbniw6
hF5UQ0Ir+9NNK4YCuRMCvjATZ069oiMOmMOmPs5ClKlXRw3S9HYmqpzLMnql0UVm
FfvE+IA3cRaRIldkfh+JUhJKtwBfGSCC0R3y4K/SWZXK1V+J8jqPGxwG++FZSn4d
CwdJvXpF9hxpRh+x+8eGB7Ozxj+u7RDkXeV3OBeuJKJCifEW6e1782W5+l42Nop4
ZOac3DMbbYuVWSAWpfdTHCZYI7zEWFtbLYLugFMErND25Vml2ZE11Dn3/Hla33Ts
vs+uGG5euGY+zZx1lYyV3ZypBR27YLtE0biOQ+PsW2sdXHGhkmcs6prP3OzFZKn4
xoAOb/S09QjtkTZiTwTsDnaRMb4TTDwDwvFznAWLwUumHhj2c3ipUOOX8jP4owZD
zDPEYhvEkDDyXYKcQ2UqujCvHR6yHFS2wxd4UfdWUapiFLRW8+uk7AFlhru9Sh/U
ZWbhWSht3MMOuiLh6AIxDyrLPig2pt/0UjmDJXQ8URcFohaeJ9SaXHTvPxsbi87I
uAzYXih7C6FqskrvOimb99HoL9WGYJWHVDpPmWuAQ9tyR6YbmS5KhF89wWs/y9Qq
BA+1lnwpsTCFWZLH8DxDODnY4VNmLVX1JhJ54Wgk3a81xX0bXwNH7O8sReEKgrUJ
fR3iJiz4w7Gs2Qfd1RLMrWXpO8WSz05dX6jEQoarn7CCSU6FlxDdSBHyofULk7ee
xnwRLAwwpUXSB0vlhalpQ9Hs4feKculsFRH8UowRSxYpk63SSdiMwMfaWLodv7U1
DMWNQu4wqhKQQdxIsQt8/8q/7sRniCUfVBZSMPOtTey7HgNF8pC6w/vHhS78bFTJ
dd0EQbgQ6HxWgcFmn8ciLS2AADAPk0fNtijTK+SIrrp5Ior7l3LU2XQIVobu+BtE
O9SbuxDqUMXLoCrSrsyUm4IcsMZYxlfIO9uvAvxdekO5M9u7HPHoMnz3nfinW6/o
nw6EIeySRdT2/S4tw3jtVTeNwFKFt5mY6tphPRtKpJVv+3znV4OMboEuxsZW7fPY
rcjYvM/QMpWZ4xFHPRo86dZSlt7hhFjDvf/37Cw76PKx8kxOv08ZwyebhlHNjehS
qAkrxJ4BfWVgMdl7AvYW/SfmxW04VRlDLDetL5dY8xDZA6kB+IQjnTZ5TErY3G9R
9lTQYdkX+/2tpjhKsLZo0eiNjfnXp3usC+zDEl4iTKgUrjcisLdSZoru4ZtdaGOF
zR2ojRMqv+3uXxvo+cjSyneWTbuw8myzTvrFFdEB4Y5WvMoOH4HBp0jz0r+1DKcJ
YcWtG3kbfR6naELHc+gebCrwCjVMFHSGvXrxBCb3N7GZqH1mXBx2QPaNVrUzkl7k
Z8K4jtNKjOrhhc65sPbKKrAfEUxwoTHQTXzmsgXWlAixVuANOFljw4WJKhQQv1UK
YiYye0Sc3AhOaShencRkThYO3twe/BDnJkwsf6WxakuLOO54Tk9QHNFHlM+BTgAr
4Fta1YQ39IHh+tC+q1TJf57ob4zBs35cOEfhkzVli5sBlCBNut4ozrYf/S3VBmOl
Xgs2mM3fhOQNGC9oDePjSfAfF6kRN9ktVg8sNP3zoi2Pd0GsWySyD7+OhMI/uP84
UCZYXR6s+otvzHugfnPAhaPFfoginDfmyW59lv9XPpBZtQDBEj97BOdzOpHGlTlK
Vs8pHwvq53yqAa0/larRDxNdpPY6mp2Nip8qMm7ED+L8jk0HagWjESFivg0nRZmg
7vBi3CO9IrwAgRcueZWnErArj/1d76aGhEbZinieHRwzHFvEhoOjGpfLCiBJh/dc
EVnLg0SIprPLRFHuLzqiE6wksyN8b/yYW+/RjPAvr82DmJ0Octy/d+iUGHUkwr51
ksnDs/u3iehYKP7Uy99RCiScdsDKFY7w3/ZmFh7H2mISrlKn9xeKvjhKHNcNEIFc
DKi75apu2kxbjAy6/I0IXp1Ps3q4rRRqcMf1qsRlPhOC7O5ThnwIHR96l5u8crnb
abwt6G70nQpfmIa4/eEE6JUZiwO/z5V48/Mcv4XkvddAXphxXRe8mwJWRE5jwbb5
b+hwfsHtI7ZBQunCkOs075H14oe+KZF+smN0EiL4HrVV0ztVkd7pijLr0v/6cXGk
rDebUxU8tEJEwgOZgjLPzrOzO0g3NMPfMcromU5k9XfdV4gyBtbxzHCXIL2YfdEW
Ae7YHU71ICP7N/bSw3q3LDjSPfeqpo6Yh2Sd1bY9NMHSpa8HLPBTaXlxXAgX0VpA
gmVOsm5HqHrl6pVDiDaFyz80/va3ES198CGIGI8eJ/TadccG5M7HBUdy2YUzkmM9
fA4HXkTXKjWJPXMOZWyJ4LXCPagvipzqDOrMNlUHnSFwtl22PbjctWaeo3BdTofA
9A27ETsLM6i8kj3kCaqkzWy7D0I7+uHW5m/OlBS/D1UEuaYFQXvHqCUGXDmaH86+
sr8BIwr+vws90bRH4xeURUNVXM7FQeDPP9G3ljcYy8vVpLFLpt7/Ew95pDsJN2VZ
YBpI1wT57uACe2DNBEyQTVJqzXcU9y6P+ADfvOqyBYVi/9V4770ooayCl2bxtY/y
OibsvPiKgCa+y4WWhRoWONOMz3DpJ7VNEw/PeWUzXzhssyT2w5P4wPWILgNIPTBI
gnBneNj4TOQ0+bDsfW2jUkgwtaB7ZFEdIj1zEZ8th2U6LaUedAI4pK0rBdgxsSVb
NicvBHyB+Yi1bda3NMiCOiIUuZfW76tQ9qj7RQag/GBZLXu6c+xlcEtDYyUU/X4a
/SZ8CXrWosCdSkqta7qWhw0AMJWpEarPPUR86qj+gk2ZmmarhL5jsnLJYBFsYdJW
o+/PbWENpCa0zZz+pDiQWqzE+IueLH/V65g2pL/PQACeDJELEJOmq1xAtBlCyrv8
esUKHAOT6zWxvB3FMNKNGxuxI/9ENyTXeOsz2FJvoxdSbBMSR1IK5j2pSb8IB68A
e8h+bWqxiOfvBGD3PBQ/5Pn/8zs9hR84UOhQnghKrPTFJEkjzW8Je0/HC1oxZhY4
nNXwJ/paiHK7dWak/kUsynCA5TKAgYWC/QuvELq2yI0DUbQXSeuYBI4Oxbos0CDY
CqSYWv4a5fnXuLCP2T+pIzoBtKCvmm1Vs4gey2WPEed2lhjrPVyJCgqT6Ob1rPF8
jFGH47/Q1lZcSQLiXpFiILORVIsCUHrDBAuOBJxXOy5IqHO/8kvltDO1eG/Xg7lH
XCoNwYJcEPveB0DSEy+361bCZYsOrC89pZssFkx/akA3yMKxlCUL5LNKhA4KWpdR
YmdJU1WOKX1PWTlR1kn6U4F9Ngc9skk49YLklMtPVMy0/Wx5jxxcAZWXUfmfhIpE
ZOBAXXIh97B+45C6FG6G5WGudLhoApaPSYwoqLENZJv9MT6JX1LI0GgFiyBIHm5C
dZZryzO1BCpFllQlW1rgpeUsa1vlLKUbntrP3fu2uo8n65t2XA/gjS572YlZDZE4
2dzJdoG2EYPu1/jbJX9OP/gBCSA7QuFCh2w+IfUBtkDhyfGwJL4anHD4Ta269D6N
fKMCKMIlfVbnQREJxi14RrirfmYpiXd1OjcCdgTMqVsoPZasdz6O5vtq7TY0vAvz
TKwK0l+dd6SJp18Gu++oDfA7ALVowslJKKZOnt1xU582mZnVNgiduxYwPqi+bqmT
iLTKpzHCVWNkzoeKFXu7RMTFaBznslcyDOpvWLOWwVzQYzYIFwKVy7pEaEo63qQW
WL5jn1tmGpN6nlJteuqiQvQ8yK/uWIbgTPDSNQfXqZeEWjUEk+C1QTOtA+IvPrOW
prWoOiEaYcCQfEZjrWAoMiUy/2IMDBMDOGBW5iJXFh+pTWi0JQ8C5JMU7EyRjH3g
B2m+FAa1bvZj351ssTpYx5EtkklDwb9ln6JotLm/jf88SwKI3mEq+3nLUUfad2H0
1q8F5FzxBdBazRyry6aCRhKTrFNO123mMF5AxLYjLCK0cdh8h/fMZp+KJR19HSeg
oUMjFqePLktsMRxUM1wQhv/hSBNRymeE4FzwZCJ9hmL2q3jaJeqIYX/kQDRqkAA7
icHozFEPLu7R9zs8Tc1VqgjKoUQSyfh/gPrNY8B+pigA6QZwuY8xUmSAXV8bTozN
vcWwuqqcOGH6BlUcw4SOvG8K7GUvHo3iozIJ0YNfUF+NaP2IUmtsxPOvShc/FPHc
y9KT2KkmpxKtt3nqM7C5nkPFKx4N+9USHw1CO8ih4e3E+TZR6FhkHW64kpJpb9BR
XXZGFp4QrsXaiFqHGIhC5Roagl+Ztgglk2ZxTevO2M3wJLcgfcQqx1KfXekuhWiT
mmxK2F1iTlrJhgQDCcN5e5Poe9elvz2ixNCIJKJbhcAnueIdea3xcirO8QW9MFzz
A3BWbC1/UYjdGkzhulzi77nuEx15ydKf/a/PQQN+Yr4B7aBEygQUWXXvOksAtx9Z
7JRMw8b6CZaSONVa/C4dW+nLdU9HeFJnMpXzVj8MYZ/891yniZtGCmBxUPjtTlkT
xirmAN5WVtw/oJgNjpSzOtyWha77C8KwsrHb8cccNEH5YSZvYZqeXms/Wior7ESG
l9zH1NpASsC26fDUFilYatkMpldL7Nkx2unjE/i1kzwnclU8nbR0rMNS7IV2Zw4w
/uTTsAqmWBlsXiNSvZ6wMqRX+8XiZCG46PXFr0WhNmNFoWE/ZVEiphOpmPqc+WOi
bb3it/zRvSbzL0iLKyIPJp5WJYfKMS0e7n2TMyrcrJDYFhE8hM1ZaOtZ8+/v94/g
qpVHNKxgkLyeULtGaEaGPmSwp1+gLTwVMjOPM6GsruplTONHSPr9bjXyYXdOwQmQ
+LR5kwt2+teCqCpL1i+LOeVsmP9IUiPB26FdqsuNUt6+CY7x59ZfbcE13OIMglYx
2VKdQq/RZ0owlyNIFKyxRTXtpXey4YwxtbeaHrTxVU7zkFgNrXdxWbXSF72yxp0O
ZQ/csGud2x72ztY4mPV46V+RtFF3VLgMvJb0+kgi0//34zWdrUsp7G5ZiVRBARgD
cARzTQAiv8JRSA4s146zQSPyM7iythOK5Tc5x87ymx58qcrCQ7jR3tzUoy4QdCUq
MqGaM/6taVfoT04Lp2xzeTfj1pTpIZxxxRday4KKaQtFNPEiwsiGBRELO2pSCYvx
sCmlH0UN4ascSgcYgDOwb5WjVyFvn0n5v4q/DVa95FzggrUSDj9k8mdZ64Rxpd16
I+n/u44PdSzzSFldhGYR8WTJs76t7DEg+Yb5nEikiXI21KnwJ/mVp9xJENl3BuiH
6gMTQgltNnIZGaUUs4oBnXQvVPipGy2Ffq8CVuvTFEUBsMS48Z051unscPCFKxpz
+x//4Hw6wqXsUB1Kt0ey3KRMbQPREFOMcceWBh1G/0zAbvU8S5HWW4RfKpoduAnR
bA9PglWDFbm6pqYkt8NWKm/52vouSuqEUbZCIpCTFgf8W7JEz9ZHQXGOIO1FGGek
`protect END_PROTECTED
