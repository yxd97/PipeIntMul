`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uc1YFfFWsxebCabCcqSCp+UvnODhXLeLnZLIx1HnQKbTLEsjuO3xqK53fRZBqnT+
iZjdezrOjtbs7GLWPa4FLE/nrWA7HmFlMyyOwkzAm6ex9uEBFz4zgREL1z8x+FGS
PzcDWWa/hb0UpGqUZ1mtLfECK9Co1T58kP2kjgZOCXcmYFjWGBDI0AJJ/Noayo3V
IBMB4L3pF4WnlnGtebLBQpXRw9em2grvXk9/VecfnzNpWnTU5GV4l4Z/IhIFxtDN
+DE4U489XmaCiJB1gHB+WLfU3BuVuHHhtAjyp1R2CMRsXcTc87wk2tg80H2F+Tvu
H7roAERN1UlfBrrjB9l0zexvvPe8XACNFe0VhPktPne6r6QzaRTvqRw+sQFOkQ2D
0Ea5W5hiFB2Cg3zGLD6FwSjmyWuj3evaYRFBU4IWSOptLENIUwLn81AaV+cmW71i
B5CU73+1OsC5BfiblYaFqi2m/qd9hGBPPz3WDjJWZLkS5wV4Z1BpZZz5rZj7/XMZ
BX36J7QO/VhlVWd+Hf6VwX93/pbKtj48TXYtzyb7PZs2S23K4rO1WPaRglfw3S9F
YuAflaXjj4CkrGHUpVPGkM8eAEjjwqr7Yp1yQOQ74Rv+NaxboB8tWTxFPIEVV6aE
`protect END_PROTECTED
