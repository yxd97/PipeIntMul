`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6IvpekIiucLA4XhnBZDVZm36WJNO5Oihb/klagtfGxEE3pVb06K/vuFezJO3gFf
YRNA+EDHI2p5w9lhly3Ksz7Lgc2eqagOv/Yrhk3Ri3rM5eD8jnctRpb+FWxTiMYF
LQD1tEVb3eDlHwWMMQcPpur5JcJjR8dPeW4KQ9HZ0iA24q5wrcoGLifa/dtpY9/S
YSQKS8HiifNflEQYS9uGugg/1YyM8iKFKGanr2oX+Z/qRHPIacscpLMzcLecumfp
ThsQVId9mIf1F5p+wXuaZymmWZYYUCdLGxyJzV4uO99f6HHBWxKaVCtQVpqiyJ83
SnqglnTXNwrENWDeOpnTPHKr64aNj4hst6p02GDfdH++7Uxgfbu2Xw7CJ4NrcLrA
lJBnMwTVPnFVdqBwKWC72nCHmMm/aE15qsxXi2l9Hu0TdirQgjBKPbRPvdAem/8e
xtvEOD6r80PCf42oDZ55Qmrst4O6NNoKvt8qSJKWHxKjpVuN24dohFfrggStCO3x
mz6/1tohloOLyISVj0XiU6H95i8luRqmDYZfSOLjNVd0QmfC59hocMKGabd+N5Sn
QdyA1YVbHRpZf2SX2XVXQM9j643x6M3SgBK1HjtUKwbwAupxyDlzJNhdSSQsIkUp
avte5rcL3npIqOfYw3P9cIvUarG0GpGZrPyudRdcdAmMdKmKVUz3eNucyM3MJfAf
mhv/u74RwRSfndAyf7KFKktmxrFpX5f8MUgcuQqQdRcW7Ux0Y6ygBwW0k22FciDz
`protect END_PROTECTED
