`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CtFXY5SibYFuHJgnUJ98EOzNquqy41WU11HO577oSSLqLs037ItIhtjkIduQ/7fG
oLIHv88+t0WLd+W2FhoDXiythBglgCHOxawf+VDfKkHgWWjmFNnrajILYZwy9TVB
MDFevCRVSQ8NMnAb4gDJRD1zaocGZYkFk6t0ywKU11zh64P3J8lvjoXyazoCtALr
8ajhaYsij87iAkDyg7m+Y6CgAsr/uvg9Na1oaO+6bx/EWMC5XFJHPDFF9YkGNLmP
RKxhsQK4GAmLrRW8iKkn/qoqIPnfcArLXQUY4FybYD5BtIAEe5WBsdNRWQw/+CiT
Vv/bfdBwRTtQCc6fBxoHckIva55Ss0GkAi5cAPpcWFdyVtgPjyhBxQ4YKzh7e4wS
IPbytbwUazf9eKi4BPYG6NoZGWIjTsojB8Tlvdb9jJ4Rr+2HcYhYl8QynuCVkpM4
qCzknEWdmCFayQxe/zyME4+1GALqx31pWaEjyByQBqW3R1+Ax+Qap0YUP8mCJy2x
crTrflHhVQZ+yHIUay++PnJZ9XB2RtxbLD/fGIpAoem208oO5XLNHQ7NiH1bbSr3
KyylCD0Z/fHDFma0lD+ziKULvQHnIzw+wsOiB0FSmUXpnJXHlo81AcX54Ph3auuV
0MoVvl0ZFYWgqPs/B/V5Qi/RiqZr3nBoP0zawU7UpCOG6oWJl0ObKfyVB5DDzPMX
mJ0ChCmriPVdIrPweQoS682vDYa0RYv7r+3NNsHAKvCjoXg2MjJbfq67riB0GgYp
SGWOGGRkY9IQgjX++vDHY0sgQwrFjb+LWgpt3Rv4wsiJ6JdQAQdab6cdgooupGIT
7aU2Melw7Z7isjQ9FszVDD3IizwsGts+S97w6rxLTHHZekPt+JQnsBe+DwoaI3eM
6Kj0ines8LrMLBm4kOz0lLVlCC9nH1Rr05PKmOP61VtLqljylfG8wl0bRtQyDPDF
lIreGxWFUePVx0F/9Br9oetGivx7zDnZrcJPgcm2JtD8dDA1odWUTggeEfdUvMcr
WmXF9sYQgclF4Xj+6i6FKzdfmCMcmTkVNqak0yC4OwP2nIMyPdNnojNajs0WQsv1
YXYdelVuMq3PArXQ4Tu8yTemf67VzL3cGqtLKRlfZqf6mnuwC2xgj+Lpi2cQ36tI
JH78yTV0kscO+fQZTAJSf5nwcFejjQgH6P+hFePf5ksZUPX/nM/sTErQZ4tNCaY0
S9oHjyi9D/YqHUmp12jMUsnG5Yxi/UOYuy+moMLBsNK8pO45hAFxXts8w1OEZZf/
JNp0DaDhVFuPbM4XEivczVaB0Zt/P1I5pFz1/zGIEUvhTr00Snath04b8b52m7vU
6gmpina69DMKe7FiZSaB9LD9bKTo4R8BHl8IFakjMC/Mkq2VwO6r1y4MvIcAaC4n
towny6vECq99z1/v/EMWGhUdvV07wNvippPY0TdfDuEeY+l1SyLAP5l/DKdIJD66
HSuvl96bGkbWjV8rnkTcRfAQ+negNrkG+YVdulOOdHMsutgLEha9RmYdK/8YojCD
f0keo9RlmLoP9hdj/UiTu/hi45dGFN9Cp9r1/v85QMNGM7eyySDo3yB6CibeKuvW
YXjNmlHirhAJkTxo3DuooJWPZsRyZnbvZFB2D1yFm+U5hUSZGvfMmRnZSpLA7VWx
NG0HydW1H1gmrZfphE4SvZz3/K4guvcFWqO9I2dzkS8OI8NIM3q+H/A3lz+9DT9z
9V3PINIrj9YSSdfqyD3M2g95lMsqf2jlVY3TNSMM5cSCZz+Z+9T54BqeixXWhaL9
7Fc2zrEzIejeqNhQseovyhI7Urlsq45ZYqnp3/3/BgaCopn1U/675fvdOauMReXv
W7kcWcmOEWJRPdI7bGW/nHnIw70eCLj3ookySkaRB+g=
`protect END_PROTECTED
