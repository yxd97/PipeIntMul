`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XNhUDb818ECkP4EqHPDAxTCIWfCQgNExsXbr/eA2wKvyHTh/z9Qe8nyuhS1nENoq
FpH468pAr+rRZl8CH4UR1CFI8PN8mYKeID3lS9nsCXP1ReE1H/e6OlnxxmYcRZje
DcxY+5IH47c8Bq4xxS0/g13SW3NsZa48Viuxtqajmt9d3I2q50xcExdUjthYNBsy
SOWkDnXFU5QlZzzq0Y2thkTyeQbuF438RSkJxJJ6UUvKBeBzD0ZsGa1qTXEeXQ60
DyujbKEF2mQqr6WWSrsBGnzi794wbSc4mJtEb/qJ2rKuIU2GpMEU1+OY+EtOKtOA
VCVZkzHjiAVpkbWiZRb0Hc1vjFKyKvdcn+sYap+xIXPT5MH9oB6ZIa+FWgFX7FdH
+FzpLzndhLX1j+SZG3jybF5EQE8x3g9NMsD2ODAvnDnBfp0PuGUqpOd2ZyBtlOe6
Y3l/aeZnOrQ4LlKeGGGZfoM5Z1p3pGUcjf6nYgOTPI/W7/K6ONA4XrpFKSNjTH4j
muP3xlogt0zfyzfitB/9CmBDoBMq7LM94MLmZl0nydzvqAlCd+YyOWDqk3pB+8Qx
hYDWqitMODKj0EKzx34ln7kylbxywuBcWapjTKbpfVoL2xrBfz2pa+5oO2htXPEZ
dosQq8C7AshLLe/+CBO6NgHNGM13ApPU5xLa4mZ1qTuUB2jbVM9QF6gHPU98tbCz
rRF4790cWumJJXXumiMi6UmWBSfd/ZttaYJYQa/b0HVD8iO2JTCPzIVRtVIESV2S
1MUs/UEvyT00Ak55VJyn6kX8UXcr8/cjnjoZ2KOqLIHemgP8zlSKxFd0ov0KPYMR
VeRXhwX0wjmUdAlmNXrkbcY9eIQeC3qY0lWfVLHiSqTT5Nmow8wHYBSUTmXD3sNn
2xEXYCp6N4sv75VVgtnTfZeB/KLaarigbOWRHqAbgME8z9hM7Fo2wDapoNyfM78i
PRo6+G8c1PW4CBYX5T08F8qvGDGjiL9b0+zHvvdkAyPy4WphmKlcD0T1mZYuPeIZ
uRUD+ZNYpxGRHYPDls+rgw==
`protect END_PROTECTED
