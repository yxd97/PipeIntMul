`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pgbHd+xXy940Rxz7vEKgjb8YqKRhhfYdIbwSgiqECjDVj62+wNgKQeJqNWMvmzDW
Ve+nlGfYzCl6rWZzXj2iv3Hlfur55/p9WDyI7UVgZJ65/K7Xg768NCvsYsHWYEU2
OdBL6o3fLlCG/INAW2z4Cw9D4VayiywcnKdJ+mG7HoxzT1NW56Lg39O8QPG0QtOH
fWs6wye81W9/pWMK9yaD5HpXarki1OvpJxVmmSbf+l3NWHIZOXqSJfzdBUH+0/pf
JKR9XoJ1xo0L/bpoq+Jiuq0c1/8qX3McPlJfiVzJh4CbSpOhQard5to0akk9zzQo
JSu0JYLPcLBRxDBqPRVBaJek9/mXVWe6pL98u5Y3ZAoQFXyrr0pR77L6rZnOmt+s
23kOTHvZ1LGVd9uyCZNXyE2GtgjQEc1L9mSbRyVEbnyXxWgWjv/GOeHBu0srTd97
h5mcN2LkVjMASSmHPwahZhl+Q3AyNgT6izVCOdV4t6p+BocHhHKrqRVR8bkRhpvk
E0pCNYjGoKJLSgT3biwKMlS9v1DXaT+2fhjpVCffNbB9MHddlK6EjcK5PwHI64VC
xrft+0VQHQzGPNiEx4yVENG9yOvS0WUtXW+YqUpOtx/WZ3cfZtn+sIWEGAVLhQdJ
e/c5tL0x+1tPVONLralm+IM+CxWKtt/HdO/vDzZB5gFWZjqcRhXqR6F3TovSd+LZ
/MhsMk92XNAwXUjpWB5bykIieDqhY3siQNWlpNlutTQlkL9qgySmbPLOz2s4e74R
OGAc6ZK8qeMMW+MT8jPEf2JMOSYFL4jHZ8ms6EjhjJJDbe7mKI4uyTvp3xhEZOfT
Ovuf0u50wuQegobtBQ1i4VXD+P13c+hxcBztz6dSJ2VjF7ZmciJLUbjrRuAO8FtK
hkTEQAvoF9TxJkoGUUK98ih42VUZf1YRrP/Nq8l+A2hhoxUx3tmtojQLaSOJqOCl
eeuABkEQpezFB/d3erNsG0jt7PWmud0wQNRgCa/ll6dyJY3kJdbdGO84/q6WkD8J
6nUPTO4zuZlB2N4scOyrVgfT3UaItTVhvYnctvDcY0t1uYpl+hlizUvBCw1bImVl
wpqpx7BmSUjQt0Mh/l9+XpzQHvFtPL8n1LqV4bRQQBKvwhHx9yZDKl29ApaTGG0+
VWJAywqc1HY562EbYhZjAiKAJJ5/Z9U1RXcQpA8bByjyzHf9UsFsxFGO9SmZ87sd
tCLEyRxShLmXvID0nItiBpdxC2waFU4B03exaEufEkA=
`protect END_PROTECTED
