`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tB2MQCjYmOMkCFCi3Qasgc1EbJUVu1XOAuX0pG2Jz7LEAXGd7IfK2Fk1aOxXmL4v
wveLQZio2LUOopVD8Bzya7eofRmMx6aAYGgFyZRyyC5yzKwgIWyIlPOBj1JmijC3
ekOFq9AAv6pmhIO2g/pWdreyN6RUNj3a8IBdihxnNrtKwmEDAZ/PR6didj2aL4+d
RXuR1Oc9SdEJjuWTw2IBf2OewfrO73NZpAcdfT7l8l4g6gZaGFKbSnpCDETrCMvv
Io9n+BzMMfxTHjKfLWs9WVvdqBlVVgpwtTLxKUgkR3iJ5KVztWmu/pGCG/yfI1EY
ADf5esBEe3U8/DAXilRM5zmJqGn4HGIIMgPzvvxF6Jcq1sRlGBOpjfepPe8M5elm
`protect END_PROTECTED
