`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXdIVRfjSMMyq/SNhbro/6N8zo2TijbQKAvPPvi+e85DaPArKVW5oGVtuw4kUldu
RR6axrDVsqwXNcAVw4t7ZhLL/lwDDLdMPUdDlvCh0qJXFq+UUWcPjZIj/S3u/ZxJ
7l9RMWTGyoFDIuRz1oUsXqMZq1fZRRCAP1hbA+utmu91hNNREsrDMX1Q0IOFW2Nk
3JVoZ/TgmJY/5Vx3aBstUqwL2DF3C7i5nstkNHuqNkJSKQXVg0aHNOBXbobkkdFj
5El8EzmdgpAnL7sUNUPhsZVfClMfA69lkOobnjnKyr4PmK7FaoGT28Ro8sqrVNou
x2vIVdO9z6kXIP01q/GK7gAH6OGbbK3+nzPu7ZU+hZjn43js9K1Hywsahs3yOuda
Xp1s2xYGTUL2ChcQqCnzAzLbo4f1V5DjgDqTA1CP1vzVVYVEzOFSDHxENhp/q8jH
qMBOHrAM7QWrVfeSWI31rUpuT6IoeVKAZgMJdAkxXkjhj5m6CMdS2EnwkFsyRbLm
fWNeWxGwF6wC9bHsmjT8gJ1AOGFEhpGPlqtPQZZy14FXLfZ1oeYEz7+Y4gQehhOY
IahGMx00kqwtkhctmCPa5kAAfcJIubfPneEYaOTENqPHi4MZHj2pyf2HlUAkW/vw
DwnFF+oDhF3XOWiNcK5rGj9ppN2r34z2ZTTYI4y7weRnfg7Y2bHGRSpREmqErXYm
+ksTX7iXco+c4LzJGIiNC8QSbwCo/PQAL8a+coksmawM0MSv9RrfjrxMn7HO3JXS
DksEDPuMRF0/HCy8GB7cSlvCzM0skn/7urYxYppo5E1A3uXmC+XE4oa/Habu+1jZ
RweNk2bkD8dcZeoRYUqG92akdMh88MV+p/SZIbUj9ON4rvpkAd/VXwX5wlk7MgFx
0BY7kN6o+QGD41Q2tT28Cg5XSSUoUVrU4AgxWPOj9Z5owu4Akr6itqrBbqG6ms+o
Rx3YkSCGeih6EV9ecPdvOchCIzWb0ZcCefSkE+REUP955+bZrKjAwnkqx4ik0aDf
LKMHKClq47MGphMDxC8KY8liuj3MMc1hZfQn63zovrasP2TzKr7LAIAO/7OD9Aa+
ECR7IAGDItecuqEhx0oNyxfve2qDwFzkT92fxiXTaV2V2TBN63P3mnvJEquB7uNK
/0Jy/P9pog+XP1Ws7t/ZutQ5oGYodlybzebsJ1GKyblgsDrLXVsn37379r94JM+Y
NSR5QfVgs8oSrHI0XW1BYH2B4ey1ISzY1CbNMkDfyPbezVHVhT3cWuVP2FR4FgdU
nVu5XSb6AuRSy1YihljkzU6iAtXe0l47S2IW7IOYzR2qLKOmhr2hS5pPFCa3TBwz
+ujE39QvEIdy8uYrGEMkgDpZjbzO7DOXiqTQK6p4aEGl7NycXHz3dHQBOCA85zz8
DZdnm0hqqMkkrX5ixh4n7n4uH2QaDvD8/gSb0DYpGrSYTnM5x3LU4n+CgCsUdeFv
NTmnv7fj1k1gL/JyHZAUe306Ujs7cU9e+s6+yhPoqlTdzygFX1GdE8dDZOmaSign
CF+i+tTgEtWsm0VKGELp3m+OWx9c9pgHfleBYMkWAgSX5V0RxU60thceYKj/Q00+
yM9v2HRFyLWxOoce67wo+M+1zg/6fFM7PjIidaMrKMpgVl3OgDuj7YlsNiMICt9X
CpKk6w0XOle6ePKaLhLurvADdmMpoAYvMCVldbuUHDfgwy8GvMJjpe7HWQ7OBROI
dMsNP/g3vy94KcvekKyAK+/dMKNQI9ijSbKA3NsMWgTitcn+R7auk0DcRSluNrzZ
O/uNB5dtOYXCa0HcmuB7isXxm/C5Q+/CPP67gEkDKAL6gTPUCnG0oG0EGiBRhElH
w5GDz7A2m4srRLHn7jwfk8BHPewJFwwfkxeyD/sj5nXw3GMCD2UP2ScG+OtICawi
lbvYR05yZdKSV9R93RmSdq113K5krpnN4VG7C3+JZcFcKEuTwQ1aT44DFR1oFwVn
MwA0poDZmYiiviaexSgAWOUTgy05OPgKoLtHXzD9DWx0/o5zFM8+EdstoHn4G/AX
p6epz/K1davDsq6Z0SFV9zHfayqbvvFZmJpCM+1UGp+QDW61B4n4XaT55UFjOF1q
WDH7Xm+26ploJLukNsg4+YtL2IxlO+VG5OZjT2opaYLTl0O19sMCZ3FsnF2WbW4L
qxn3hUsxWN7sRWwMKpvBvdnQSt5SpWU64NjK085phTSu2eYJNFegcrIFSIHKZMgG
TNb9KSEHyTnCfjzIsAtoF5S7hyAi96UJsJnTPgBQsSJE5cq1xrtwLVafy1BQSPTF
NvsGx17f3dGVYo7IMm0wHhUvXvevVXpGDeUnZNjk5HupmKimi7AX0PAhOHdNRAN2
w6Py+qYFOo1it8QddKhB3Cx+uLOcWVejLXWEyT3x2c10/HgiA7TLNzpjvx8tKIcM
srMjfe6Yan8D71scxiUXYsMIJWlCP0qvbRVbMuxl4BOcjzryoxdF9fSBC3DtPJGt
5ElVSvBocY4uNqw6A8inqvvlULS3kJbkpl5pAPFHZB7kk2RnZdgCiIK8OI8aBlTU
aRrY31W7/wMgJ9N62LWtEp0x6SYlx/96VjKN3p1WWsyNA63+Zehq5lPszxovBxxs
+IoWglTxVdeHm/+GjCPD6NabA0+XD2wqWg8ehxLOugie5MW7oyohR5m5s+XT/6QT
kAp+jIcOY07FVDLBzyRzgM7xldscX5O9wbm0Nrfn7wO/FWbY89o1plaVVn/FVvu2
4LRkFzmti0n/ukO6P1RV/EtTEvMmwFN0oTSHp05bRO9DqR9dE7OiH6LLD93cMmwC
SHzyC1++Yc1mIhkCYNghmnzHTMaCRkOwOum2lg8+12cXCXcER6Pk+3UdA9B8WNqT
WrziuxYzn5wMheuPQb2jThYZqWTsdtXrxGdK4uevvcgTlbSP9biOhmA3E4f+6r9r
Zt3YKKNoBqNUU3TL95YAT0ikEaXa0/S5LZD9nWspBWiiN9oSV/Q93mFgI30ltjry
4t0jdQwA1VyO18fxmwA5vCGk7xF5yoAoZMjcQ+rYrPbkPqI9aIEOhHl+EXkbyIWr
ICHB6U1PrMcl5te9bRVxdBxWywxBqDpklgB5xRZrjAgoqv+LYN/+n8ZpG4XaqSg9
m9mcRFLCIR8UGeceEZScpUQGQAdkiOYMCKvo7J4XUTZ0W4exIy9coVbc5odpgv2R
gwLW5Ix+ESYG+tE0T/Nt5RuTXUKPqr8TPi0RDUIS3uQGus6bTHZpkwr7icmS/K43
GM7qk279wdHvBxLVpIWglNzcGdTQtOqu3Ts0XNFWNhfx7apHqC6NWN2tw4uSKmi+
znHgWM8v6Mneh9Du/u+oih1s7/LNKX89RrdknpQbHwqXUfBOUHgL2zxsEM/OGLNL
8QEtQuhHbRERH+wOOD5MhXybVDDGlv6sEA3ucyWJUh8vyMBBjSHhIXFR/wP2SX3p
o0j7J9ZP1fxs6H+RZ/wlMK8ZY3+JB/vi1g5qPG4ubk8eCVYZbxU1LngQz/N8ck8e
arUu0IVg4DH3+BJGJ+J7cscyFBljq97Lh1wyjn1pA+Or3MqSwr/26glu2+EJ0+B5
ncUURuiKB/Xkzrof3U5/lKvAx4oPc9xeYhbROeYwufQJ3J9uLyrHUzRNw50dYEum
RstPJN4723Co48f16/l0fnq7+AxjJ4svoURAEMPILgvX70j/EcoDCB1rYL8+6DCC
JbT2nkwyILFLpXiaXxeA+omaArxmaoQlM10/rrHsvD/5BIoHjQPFwdibANs4Rpnp
c5URz9EvdTkPpsDsE7aDBynvSzXFkngWFN0rFUa9mGEvDUhPu+lcd6D7n4DMdCfK
BTiFx5ZKj1cQFFJsf9SE3IFcxUVvay8IMr9IKZ6trzxDO/Fx9std6e9DUqTkxxtj
2zMtrGe1x9BZ2h3GNEs8oi033CS1DXqYvV/S+7dnJd9upy2koePQvPQ68T5EOPl1
vvYkKIOfNiXHMf7PB1DLuYClSt1h8sTABDDg+YC+GOElqk5I8t56GBGHtoqN9nOg
HCP48XXRW44oPh6UExXJD4jqtxhnQ0wcQmBfrggFJ2IxhUC7dAxb+kg5Jy1QWc1P
4K5A37eX9TiY37itHkJ9ky793fE+PyAio5L5IcdRIFl6wYmOlFGyFg+op9BIg3qs
eeuAh6zozm9PHqBfDxEtMOSzemz50yBG10EQSzdjuunEoyTktvI3iOIUY1gBWtWm
DxSbj7TL03/40c5Tcqn7ar+c6Dd0xMyt6eVH3cth2BVLapYLr0/XvB6UtAbKdLmJ
SI9K4cTO71Hgy8A9LTZ68J26UGjGj1mT+HpEqbM4t1Ta4oCvSrtDLNMb4n3lRbIe
z/4kTqGWHfarOyoFIb6dMKlY+jtSWtRzyuDIyP8/Wae4ltY5wGZKehNdOkybjaKP
lsMVTwthmfYFiM10eMTWs1E+GtBu2b347CNxrH0EIQS5rrCxQoYwpFJgTW8i6p5y
tgOpd8MSt0j80ZZ57Szw+CPXF9wqZ4vo2OIhh3uX7BTiS+pdnROLUVfKR0cifKWp
cyu36zaj5Fi0xuqpHFekx6Brfu809bPHGVmRUg6DamTOGZPxStmyrVO2nq7U0Drm
ZZ+66PpoSwD2BBhOGrf/hB+C0VyakQTcLFWUAY4fLH0N7Q62nUHXL8+KCrgaC8Px
z3Zyi4yDY/J665ZGa+rjfzAl+DHswBe61NIuAJtpcx//R5hhD10Deg/AyoRmkb0u
2bqUBymEglsVnmS0ZHqvYCMdgEv8E/hlZeBN4RVLEOsKWx3TjDF8NL20Qq3JGI6N
/c/NJWKfmrMCv3CXz8WedC+YbWSeGMJRDZ563+v6cjVgY/9UbaPuvKvEqf5uvP9T
tJxpBB9cIkaYC0OwphViN9IktZO7xy3WBewRJGwQEuhvAG5VeMJ9xjvvssf3KIbp
btSxxeSgwpQIwKM16udGW2kh4jjj/Kce6PDGLmIoifPtlrUiF/AuW7+SEiuT7bF/
0FSauktbsDJgduGetU0setZuba290ljolwjTaxgDPvtHnOuona0b8Z37uKS7sLFR
vkiq/KhqfOceY0lcEvsgeOc+cFCFA+wMDjQktpkZ+xK8g1Y1BgxFm2FrPO2lqHA8
rL6m/jCEEewb5t9HUNRmug/mqdpAr37wpv8xHLrHq9ewVfMpMm1hSX6F4r1hHszP
jK2ezmKWVz34FfK0oeHzPNKtRrEYqr7huugqNzlRAWp4VW7KgrNm7mcnc4H43mKp
FvPQoY5sERh/HZ4qq0TvS3HCgjcFA/AAryu9/46oQeTG8vFzg/GO8LKJhL+5l9fn
A8oeYUwwnYNyEU2/ibktf9fVeAXBRAO6FVlcomRr8meE2HT9vCNgbAh5S31cfZSF
sGRM7Ieve6GHsyHtEjyIbOyoFY0TL9b0fOuu0JsAB+eWt21mRzylagfp0Hx02iEH
Ce7E39GrWo5lLWDLI7rlquOcmb6vOTBSNz5R1Ycacbw/tncMGi1Up2extBKDvQnl
fmgDMWZ6n5q8KMoN2mHg4cGsSOc67ZiqFK5zJ7Afac+gnhOF5OIveG8b1R0TiXcB
tP7QHNPepG1Eif8uuiVAbSwSFrO7mQIckxv2bRgp9yuEK6OlwSlhaBotpBB6EAJQ
zsLmnn3mUeO/RDctYaddUDItLf3VWFy8YTJUL9e6dddJZpPRHlui+wF0163LRyKY
eSLixPZTUogi5JGdsRnEAjWcZPsFARH5e5XiXJKZl+TVk3RPKws6BMhIKOeUCksj
rl8FsfGOE0Gf+plNuhB/AgGWUYBGdlHHazGKHv1Ms7cOHokvEsvCwPD41n/Ymh0p
kSzzGJhx4h2T+xg9zmtEzNwZ6leQD+I7Yg3p1ScLf7pIgxhEF0kOguIlBoN3mf8Y
RqahGcUb18E/h1KSDdqtyeYoePbsulXSJAcJ640KQpaAfksq1Yxv+waZ7sXhA2D/
vlVq0/zrf5ewzZ3ODj4H0m2up5k7HniUs4ET+YAEKpw7n7+t3m+WlbZirpy4smpN
C/o4Xf/BQPueJyIBnS7IHpKw//8Fxxmivml3WwrRGzLvDhQ8lu/TCViNxJV/s5xV
B0mEFt57lRxZk4J9hBMoAq+QeUKGFEX7B09HW93qt1GvVkj333RaBJYDlB6nYw8w
HE3G0jT1OWjTfAAwrjC1MktkLM23brCjGWaNdz2Ym9lzxPSqSCTwWcdDnyLZpSE+
QDhmycfD9794pJfTAnu3JDJGh6TkGeQ1m2FwNmtPZeihV3iPvpNbv0g0oI7WM2FN
p1QoLeMEZAkNf0e8eBuxaNvSRJe0rv+Qd9nZxIhHtww3mmIzkwJYnTDhzDnloYck
t0m+V2vUFKCQ6ej58tbVqRy17FlrifZTp7ViU5nx0Clsoof90YSex4TvXT51MUP9
ZDoRc+aGWeHFJ62s9jLOqaPUFEMOUoXDE/bGhiTzDuraeYro3gT8pqilCuswHB+t
LmEz1N29RTLEJ9+hdJTJFpt1U6KWID4k8JmXXJxMrLAb2YtcViL2jt/Oq7lX71RN
TeCofAoXfQK1MnjStFpLitIvGtryW+mytbOkAArxQfFvSnOtFHkNwNn05N94BqsR
028kKoJWnX2N0G33kq8Qzz2focro1fyRiRiYKKQUpa+4dLGmRJt0Y5yWkUBcdv3U
WSSU4xPsKRbR0TFHNtfGY/l8O14zT1LoLYpoYcYXOoFotGPMkRGJ/PWqr5LaBjDN
jk/6kMmp9Jn4S//aa3B/fCi7DMqcqedt458VazcklJ1YLNrQuZlVxrf0SlnugYen
X9V+I3wkPc1QPcZaIH8kZhb8x7spSlu3rD/vOhTsCd+1QicRVvCqh7qk5qKdQ4/J
5mglvNjDQab7WjZga6TYS1jfNcET+1VTVFoIpNMhDEAOZ2uMkqzFJgyOOivHJDkv
OF0prnulo7mzhakrvDDT4U8zBitL8IfUr69lZiialOw=
`protect END_PROTECTED
