`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PuueeLP726h9Dvjad2RkCtn9e2OC7br4rcsAKHsyR3hQP6iP6+sGN/X+CHkP3sUS
MI19THg04q5Ta1g9ZxzqC/OMA/BERztSPl528wlWMRWP1n4bStyFivq8vG+LuzyU
5FAettVQc7TjwjaAoxgzaqPXrwKjORVOBX1QJXB9RtuY6wbux4vf4zOntbTAbnnK
MoJ9zhV6KBRAv41pkMAW54VUoQUjIOXcV/qWDeiMEodkpxpqzZEF315eVCoZ4BDP
mx4tv0XkkPuLVL4GQajnH2bUOLVoXzc+cxTm0bE2Yd64ck/5pliwBJnaXJjoRWr0
vea4p2O82xTxfIBhnGbrf7yAcYJxAhYQxFsCnYsRRQ/3/8ljF4HoZAXtEbBjtWzr
GgogCofNcL+1gm6cDVOXTiQPe+r/I9iuO55zQMcEQ4c=
`protect END_PROTECTED
