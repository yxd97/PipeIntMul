`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l58a6ZMIw6TQUQEtCNwsUcnn4HmqaLR94xUbbJHuWYqfhKZcAv3sbiS36LhYWesW
zasCC7OX0fdjA65qdibwinoajsIB6ViVyS4m4UHFH2AFQna3MSoLh608Jkw97Elb
zlOHsnhKNva51OxR0DzOUUF/ChZs+JloEhc0gMxCjKu8dYX3VVX4JFvxzpxrZgkq
dU1tk5/UXLzr/KWxFiR/fMKvCDPuprFwlAfrBiVA51IakTfRp8/lJ6sMgP0DEUod
1umOeM/9SnNi8naYxJmWLcaaMwWzLI5RE4+pRoDeADZtS7eRtOwt9I8u+I9CsVs+
9uVSn66uWPiTH374dqcGN6gr57GeIODKKMESoA+JuuqcgVHXlvsYP3EB6xZw+1fp
3LX1DHESz+UcXpLEqns9BA==
`protect END_PROTECTED
