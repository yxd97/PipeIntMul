`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yn3u4J2M69pv3RbKtl2yUH1YXkp6wov0VTRaef8qvZdwv9/s+4Qf4+uDZEgex+x/
jqIS/vmUxAD3xg4D6HHg3OVy3oiy8Fm7eZulvgeQrsLpAuxIXdK4HnnBQ5cqeZuM
/EzUPQzZqmjfhm7YhKRseZ6aV6sq2d2u4iOxEvWbq10TiVmlcRrFPKDP2kquMK0o
RR8xYvZc2ibyR8LDk5N8In7uGIre663HS4M8gaEXR2hs6jxnlBeCsK0ZCUt7ZlGb
+4dunp4zPl3QYla8RxhLYJ6SJNeIt7WLPz2RY7ymtAXLuYIfy3VOORTUSdlTUajt
NregfXyF5fP30DVObvTVxg==
`protect END_PROTECTED
