`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7smWEbTLQn9RweSCysaWtnPthqcxr7Hmox8/7+Beh0/grnRtDi1+i7jbNGBfoPl1
QsvvLvkeaPcwHS3ow8T/lMq1DdKj2cVnwwcQOIiTFstC9RIfXG8Z1Fj3wyDqFU6b
maghdWSJAQVNrIvvBTlcexUYgLIyONwgAwAKRNso+LTpyuPnvQFYErevVE1urshd
pAoA0dVRk+CroNq1PrhwdWXyApevhiuPZlPHYFD9B8ao+sRcytUKl/7xXDYn7PwY
r7OIEplVz01GKJd+xKOZS0hxkI8ZrxUgJCk2xngN6989Lk3S7OlMg8zfruOhZsyZ
dH6vR6QBG2A+O+hNPxe4Qy8laYXplE7h0dW+B8GLZFDuoA6o0z4NHRnPIl8KZctA
bmMbIGfARXlfSPEbvG+0EruCizg6yKxmxyzyDddyk7VUgXYF4a89t5dP9dUFvygi
dHzpAA2i0UyQVcTlc4yR3DODoZBl4XVT1XCyoWPSR1dCA6yOjQ3IWe7j25MotTe4
QvdgsooG9sCs3186hU/MQEWPZIdqvcFd3VNxU1jW8JN4EdMqRHhPItfWjKdOER0y
GmczK6SlpAc4iKwWB6c7nNM8bZjhvne+GMN3wfntRHqFRH7WBOkLvnQjImsnpFHS
bX5vJXkTBVQvCh+EG4DV/QFH/AjTHJEN6swRTkbYIr3VmO2MtysJ3uGD/FX2Kw5l
OA5fabw5MdJV7tEWwytRR1DzDtoZdirKuWp+97if6fQLgYP24Kxb45vJtPnlnTCN
TZ3Gix/41zGHutyDO5un2fBDxKDbRW1xCacubERE+woGRp8he+ZohFoD8UqsBoHd
Fzp70c/eW8Um16HC+20g/Q==
`protect END_PROTECTED
