`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AAyjwML4wJYAV2oiPw6c6Gk3aqOBy0nf1cXPfklF8XVql8xWLxJs+WrOQ0JKtz7/
EmOULdGFWZJ1KBSJjNsUSV0e41zeZqxOnurTUmK94jb4fA+NoLH4tgNmtawQBAih
itCdEwJph/osC02MAUv1J15+8jhKbaQY8TlF2PZJOCV/PWONGxfU86EwB42wPtiA
xX5ANXzcmwYvg/oLxHSXNQT7ObXouH+EFV4jvLvyCyYzfdKiuhLTta5+P9oRUlDJ
QTaT8EhhqKs3/roAcdDvhQ==
`protect END_PROTECTED
