`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RHNEUMFJ7LDdYbuonDM+k7VSWdOXI0nmk5+753cTaUlDlEbolHWkx8jwyK1B1wTM
mCDpjNW8U9HAXLDMP0UWa2z69RsKXLfN+MdcM2Nuv2Y/vF7AwOF841CK1dToq22e
MZtTjAWollSJlgMspQWewoiD92v7P1ggBcfDW3FNElkY1mwGq3AYbs/AzgWzU/CX
CYK+bQlWE2pAp9no7YvgA8rGxDmJXSc5lGe4kvvPoCnFEXW9KoTnNjH72KYuZ4fs
QP1gqHTwvRglnBzFd6rVG7uiwAxcAdXVUhKFkKCFRPUz5JhuSdAkiMPOVZqlDQP5
iJ1hqiLgUyjBTBBRL0pc3bu468ALMcHjuZIRP0A2Aq5IdlA2V2EZEQYTZr0VcNrL
e96PHiQOZMr2IRvTPkkJ1NwEpPuXYwGyBHo2B7Zeufm9hbCB4EO9Dsqb4ziZ3RWi
`protect END_PROTECTED
