`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uHctzJzDtVnUPHKM1VjfgA3s0Y5jNdSJTNZsEW/0qLDtvVJWMJzH7K9526vFphBP
sYTNPFARQLIXo04jMf2DI2OOJQVCrUpZDaTcDsgfyPVwRc9nx8Eo3+7mC3X5cZtM
++AtggK4wyaPLhLiEj32Z0p7vM3XEljjCbjrTPic7o2KU9OfikvXfBjPU47+osxj
3eF12PgbTKWjgK3hiZgdM5VLTFfYKrjwOpKjoTvtxkV8s6YmeaLUPSXcPG/FkOCl
`protect END_PROTECTED
