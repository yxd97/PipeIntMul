`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z4LpvKtADV6lHvNeyxkUGoFea860WMLLN1fgqCWcbQptsEvh4NJxyTw2rpSuWn5g
LdsFQKG6jmC1QvzSVPzjlSa2qgYMEPAP/gKIUQJa+c5UizzwsQUEsK4xWJ0fSdQ/
WvmR1ZQWwOiqlVngU+mVWNHvDYumeOrThDSHJNPmT15NX/tO6+mHnN5oRMTyM20E
tiVB0pbAuddeygJhtBRNmocF1rnkTWRkuQi1xhbeiE+Ugt/1YC6uyLwgR+3VbqYn
OAnYe56lPbYH+FZ3oLl273I7BqJ0hkHDMg1USnE5YHHlL1XG3DZfBm6bREtBFZH0
rhfrLzkqE0ZEcwtcamsnwYuATerb8fYWXh5d7i7rltQkvzCtknL7QL+v4WfdhDY6
/ikeXGKKnVYDlS+Elp3L8mF5io5dJ//G5Z0yn8HB/Wu67yn1Bexw0FRMH906b4wM
ni/ow88XVwt0NrK/XqD5H8jshkCswckd+Whoy/BKkaNUMdYLRaZ3ca7PM/ILTb6D
5S9EL0PCXWRnLdD5lw/W/Mr6Uy27JAtQ7K6VmGBLEJ/cHv05HlHVWF78yIno9CDV
Ad6M7dilHHgZKdYO3WWVPG7AjH2EE3jqx7jCW9N7m51XV8lP8KtQZMnmCfyHvJ2j
E2OhU/tQSB4nxmzB0dvcuRscFTbW1nCHK4XjI+eD4ydNF18aWevW6+C2Iiy+FhdX
Fg+zGSCnCN/cBUOojCuNC/Psecrbh5o0wwdflqjXWhA/P2dsM7yX/vlhbBgC4fpr
IfvM5h123Ma66LmxDKCESxl/xa4fEaA7DnQEbs3dfJSpPwpCxyIzoMgyxsoFatZW
idBXWkBUrK6y+L5JAdZDmQ1fWAcrtdZQ4JfRr1c9e+z8UyGwhtSh9STMxpNfOzDu
TEJUC13FabxEIj/Xw3WEMktQpugnU3bYNbK7hIDvfew=
`protect END_PROTECTED
