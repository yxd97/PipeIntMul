`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pduh7s3/O6Nmrk4O+lyj7WsG5EI6ISZPwMRegip4r0Jht2nutFbyYd+S9KgYR0+L
EVzLpAODyqeqSIWniNqYw8SIN24Sjds/0eWg2bN/18K8GZK55mht87C/2BoVNaEk
3wcI9YQ87bnHzZhaTpmWqdXCenuEwV5c5taz9vwQkLx6U7Qy4kZHOBBdp913AMWa
HkYOUFtj8PLPxoZm1eMU+PeEkgkT2QYdrEpkAnIs82nFyU476q5dF/QcTtKXubna
RkW6UCdPyiJM8mTKb+kjOcvWMbi/M+bCDAPqvYiR3iNry6fkN/nVTu8hY8UIpXLw
KiywJ2UiYfemu0CR3bgxyMbLWzXvxKwRTpT6i89PryQH9o6BUDXpvCclVDMJHoSm
VczYcmWz3RscPBZIGxvTnsCPWEo/by0Yaa7wXWTk3STd5ynKnLtbn5WDZvHq+Paq
I3IxSvw2EcYiaAAt/fdtwy7WBrqPlbrO2MKVg4bndRuUOPnUC3TBdws79WSPYwLe
3zE76pWeIzFEaXwkphQFrdJOsIQ+e/EznJc/lIIt25rk62JNLmhsBcm0IrBHIZlm
OzIHZDgJxJUTzu+chpJhszSteWlDMLuW88uacLKPD2X6/K3mRFhHg2qvZmITTjCJ
EGMnFD8bYYd3ynXczARDSwkYJIe2bh1EzO5Bejd3cCbxFiY0biFIDGzfm2MmKlof
3vz060/wPl2Lcd+pgyoB+MXJbKxbtKCgT+ZRpq4xkDnEmndXd04aPE+RmYDmdeba
buI1q+IpWupE43XcDkf0J14mwSoKW1gkU/JVmRsv6Q5DYoHIMzIOAmFH5SPutFkF
IqRfqzqyMXjJWuzOuMV/uYIwlhxG1OU8NYQKmp6TSDg2+oL1o4RizIAJQqWauUxX
1pql+Ex7VboHdqsnKR0ckxO+IoAZvoH0dZEy/5dk6Yc4B+hCUSFUAIG4YZyiHHB5
Uw6GBXGBLRKba4bVrcguZHEj6wHHMbjriCx+qrOJwYIELSXzBwtdEX+PfYW1jPsq
K9PuD8nR+4CDwfPJaFxawZauPksyOfx5mEqo7kgYmz7DlrgduEU7n3BU42abH5QN
AAzHM57FFi1FyvHZ5RII/xC2dI3ejtsEpUzfmCfSC8U3PgamDbq78DvbeRXmxmjM
dwBGTXLmYYhA9fkTZG4IFG9b0GH/zBXQT8a689ocU3EFoUlhAWgiQ1ZW84z0xPci
9hu16ZWzsLuvySVPNcMYf5hiH3MWi8q0beRjl3L5iYkdEeopmSWqf0XEOD9UA8rh
rnMtGlSYcuzrlXbWwpXmqsBatVpRsvf4O/l/OtVGBDPK1NIP6dSgoPs1dvx/MD/u
6dvEXe2HtdyFVSdF21q62HzRQS3s745L1+euVPl1A7XQL/OaH2yhictNsTGB/4NX
vGKG0s47N+OhY6thFqfBqMvEOMDChgzDjZZQGP5QyzcNjSkLCAL4FK54LOAbNyIl
Mmbd90RoakEgmRQI7q9cydeatl/RF4EvaBfKadXZ92+ShhD9Seb25BK4y+yM8ft+
Y5nJkgj1KV+t6b9t/Ls8FrmW9MQ5kaX9pYqk9bIRYVVaMttHudA+4M8z0sZP26iQ
Co7uWe/l7k2SobP3vV7pZF1SGAp2rdRyNYERyq5orUw5bMJYwt8O68QOZnQfqpdY
hg5aa+UlnL+J+3WgB+JLjmVZQjZazoO4gvP5M4SevpTVn0Vvc29G9OMJdXVBc6rJ
BPFM/I2f7WsVcYLOKBlYB+lQ5cdmtpT3y/pwbihIwhq8xMlU+fBCLKj/uFeIsBmi
ZBq2qPRl9QWCwoVAJblSP8A67TuH/GV+jD8XGPZhecJxVEkjEicj1jZj/KyISO2u
0x+p2bDuvGpx0ftmmN3x5z/5mzeQMYBmYsMxq3t8w/N0zudd8cmRHkN8jRO+IkA6
tW6xsaCJ5i6goMSfRWPxiuC65TDcu6uO+h2ZRkELatRdcdKowxTWFYeVZSlWQEHc
SZS/gpn1pc5WHv68TmU1W97RJhzYeYcceXpJMUj+/nCwVGUJ+jJ0NLr2rrYwsN0M
vKel1ahfhkoaCKG3mr4qd6NKJPhv8XRIEiC9OtU9x3kYXWZbdKQ+eQAMbHQIrURX
tH+KmRKuGU/8piiMnWSbTrJKAZ+9vtSoQFzrSbvvwAvdOD2z30/6nhN3AZ6YCeSM
M+Bh3B6EPjBYgWM3NoIOBfwXSW2rwFlETCoVN4BZrZhibVF6EtSqlkLUTgJyQqQE
gktPB0S6ZSFwNHQqlyjIJPdOUkKuGyfq8dwO3nyg86nEa8gBc5tQOhw5h3KsSOhz
NY1gmY9KS2lSe6oUISvQmzjrCP/rtYe4cKuSni0grt8ME6ySsT+UE/10Ug15oEY+
z/+D93xA1lWpLKONdJrVARwPSvzgIeYWGBBdzHdvAvEkbK62xcwYAcSfnziQ1eei
Mdei8/l3XIwdvvx7X4IXDeZoIKzUaMDWK4bX4KUsmzonuWrTdNj7FJ5/MkGJng8S
pislu4wOpOnG3LYeWOJH3C5i2rnT8xnKXuXA8uNAbt+42m8tbeiLFHxE8pUdXeoO
jIh1XfHewxgmfWr7KwTSH/DZyAHmEb7aoP7kj6CUaY7PyZX/ZwRLYq7A2LkoKS1W
XuBHt9c11+sHSuEszZSmK1S8f5tsqpb8Jsyuwf0lxJ7fYySmCRVgKsRqmOEtodx5
i+t9A+MtuKYnLNpLEYx9qGdV/8Ave+vVEWpqpp5i6wua0j3nC2KydxUUeUZ0hpAS
6w9WLjIQkgkYNvs4+ENsExt16zMExpDDhMnS8ubAF3VR42DLK7Hg/4D7d3NAcC5H
9B8qgoKKLeADWnxtUBgZ/MOHuC/PdJBtECsnzzCGY3kywH/qO5SH0Xa5BbsxBSQL
elEKYU/pQsKX0IRH4khaLXgL4j4gX8pCdWIqRN7+elwyNKZhwg0cEgW3jiyO48D4
gJfGrBBUxK2JkzRmwNiq/8CdM57I5Tjax77OceoB5b//5qhxfIFM1qvUWqscNINt
jqx5ThkdTbZuF4MHU9ZLlsvRUdxmh4t0S1SJVyqRteOcfS+SmxMitEZCuL8lUgkV
+31PEFiOOIFhXEeIzbY6ocSdatrpFgwsRjJq0culosXGQli69KmKsVWRrbUIEzSs
yVBKzVqhsfCFofipuNX5TN4hIv+BV+WLAVIqVlQ+5X4=
`protect END_PROTECTED
