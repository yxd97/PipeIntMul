`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/Jrk56ZzZXsGxEsjkRUK0MZnsvy8SKOGtzy29aAExj43P+956lRTh/eNgUROsQI
XhDgRb5oW9jwGrhMipiqCQmVCz3EAH4Zat+QbkuGvC2QEwM1d3hcgRp2QupLg716
I+Ejv0eWOvxIBmqqxEsVGMD1k87rfW8iIaO2dEzX14iD9EYDHiVxRGzFpEN9vz50
xfKa4iM1PFn4lSlFN6LcofVwNNxGo8JGRK7fYcqHXR/YAE+KxxP7jVDny4epkH/G
z00HWIQzpKRABqWwyZYVWmTDRparev3A/99oF00izWklEHMsO+W//J84lfjvVFkc
9LO7M+XN3j1YxZsvDhu86la9fBo9Y1RkhCOLkTsWY1+zrQqSsJvBGXwNi+cSpXRR
N4xfeTkD3njhWFqC8oQ5OH9LfeDepBaLbmLz8UH7Y87mTt2IWazt98V6zuZS/8pI
rlPk+K+XjY1jg9s8VJWcGYULm/ssV9faZyvWW76urD9ua4lQn0ufcJSQwmWpeA3X
`protect END_PROTECTED
