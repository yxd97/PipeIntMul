`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOhZ8TBdBjOMY0T5Lvl+oMbVAT+2o3tWdoptgKTwsw9hiVJyxRqDDFc216RG7mz/
rM09WaNBK+7ZSGNHxGDr+a+GlBdMqkQ3zcTQ+ar8b5V8DQmXXF3Zsw0ErStYnc4q
SXv2br008GhvW4jrE37Z4A9L8E62ChBAHsjTPqfB1yvl08c1plfSDUPooYgVhzwI
G++LA3Y6wp3Sqssv2czj3GydVK88/CWSArm9V3oP69LK22txIL3p9TnbgYLh0f2p
8tqS0NDEl6yGuFvDUDOoMnE3zSipnEaashHvOReWCMXaOLG4gH7chulr2Kv6Bq+p
+E1kg4kH8BOILCY2SUigRF1qvlJvS0pO0iERKe5xDv4qVJah38RFM0+pFi9WVlRG
GZ1mjMh2ZJNFe2sc5O2opEfOgZBggGfCfVwVGwljikmBaPVN6qB/RTt0pKrG0RdV
Ws9lTrZsUprEAaJFS1C4kT8oVBfsWRUTxpXVHJ+Z7TvZ7/HKA80GQvDBlx4Mef37
7eSse4/7TsKWpvmBPB3NdIqUaQzmBzc3r6Z1Ho/sfvv1DtYusK8aIBe7TfdCkqQW
JtzCuke5bWAJ71aLN4iJYpKVuHmoQqWnWfyx4JDuwT0diDwo1TEK8I4yujW6zTup
Dxm9TCplGNi1mQtK1iOjMS9/jPMHksOEvXDDIlAFYfIzkYu7pKp6Tx8SBfJy1D3G
bp7bctYtHqwLVeem1iZj0I7G27YK9IGvP4a82lE2DEpowciKWW5v0St6GMnQezaM
IvMEYHEiTz8tPIhxZIf+bJJvG6j4w/Zoo/6x4533zMC/V3IzNMLml3+O6DPuytd2
1DVXAAN1LThLc5VvOR0Sji4EhW4dhNzsfk9dKKFeP953AKFHcT0b0vWOzCaiYDB5
AEb2WxISbCBxcWwC6biflIsdC0HmDVwN/dwsnfl+xi1csumt5/Kl9vn0/mCUTN4D
bDFcECi83faWuYlHFFJwDslAjB52B8i4DuJ/JptwYNrOQzh0xsZXNPd5tVhrPrFC
tuIT9gmo2Ut6UhuX+2IxL5QpSjz6CmztwCnt0sTPjDyvCsYrgv1nPSuV/YXtaExv
Gs2qIxwFc9ymY+IoajQoP4HIJwElzF3DYIxL+681xqnCCouMXToewDz8gNsvHP+h
DC47tvVCCjcdxFJwuOa4IHVR6p7XKljsX2LkKlBz23yAFXrNdBKw8kdPFkqre+XD
pMEjGNSifPYWXN+VnEP30dGe+kq2Leiuss6TkxsAgW3+OQNknpOeKvZH1GEv4zrO
2Alqn6rCxKkxoDG31qs39pQO9thuNAe26WIhwYzwbr5ZybTNyau4zBFQ5dikLjb+
zBkkW45Ht7kmGOH0V4cQzahrF8+p+ybbWd+z7RHjqJxp0yy3ydaAdhmfrMHZHDpG
szlsERFBWRA7ssrAUSs1UIG17xZSHGScFijtKsuhRY1tRYmwKUDqNmrE3RSsNxVy
LgH703B4eib6JfEiw+a/3F6qurfdsGMP0jHuHvs+7jKSOIProgWwfi6xbGDfvMtx
CyqynsPTnWRw64yxdXfc0mAB6pSZ1/UyvjIAPwC3SWmL/IlLHD1dQE86XOmPLlaY
LSHLtoLMGTNyql8w3R8KusyoN1yRYI5qcDnIzt0FClDBdzsCwp7RK8nrn8ngsq2J
aal/YwFU7WnDA3SDEZyNnFk7C7Tl2xwH4c/ARU+3MwmkdBtVe6SCwIVFWhtEI18G
spKKw0uErLcpYg1ePr3jLBkm9V6CR3sgEm1HXGziDGHk525aQGl0jT1DWhYWEB/+
l+v1e0+bXj6aNQm7jL0xoJDIPE4/HK71iBVW8z4oPQxxtamozD757w7JzUKZ5Yxd
lyPj5FaWim8htE3sB4BfHwwv3RHjcwiGtRhVejc+GCcO87IQ6QCZqyTg/9XWG98N
ogOKldc/MX1reMFYV9lx6wawR0fJ8eJsVXLicUjOEtDieasS8ojMaubKxXMBJ4Zm
cQzO/rMAfPiRAIPck9eoVCpEM6rR9sahzIu3PoqpuP2Dy9WMLP6ct+8Xg8KMIGSl
05K+KSSfNQcLk+ooTVPRn/5/9+sBPYuxJYhIuyPrpjveiWD8+2c3XVPhZcuEQnKN
jZUtCdlesKJZvkHNwk6zEam95R2tZwhdZJ5DzE/lpr8tCYhatAb9g+3pAowKJOuz
7qalCHM9Z56p/DJZKacjY6jRRAHfyauxrLgW58Hl5iRhJuSJYONcypqXjX6q+o10
FzBjw9xTo/xptu6fYj5butMJopLQsPT22EGJyjcniczbmIHSGsuVvHr1BsH4jvJ5
NEjfW0kHlmJKm76ckFxbrXOpZ85SLf6s610xZvQzsJb+9hsjL4TITUrMhgzsOrrc
EmK/zaoCv5ckMOBy9NF4aMgl4swx2gscmIfNGa3xIr1QM9qsEcpcvM2ftaJPjUzh
h+dakYKDFIb+LNo8L1him5H6uLzXtjQYbUa1AJ1M2go2QEcn7SASuMvmwxFm8Nwb
cseQlnJH1h4x4CfCuwmk83t3ND1rae6ftIjqBqQ+FKM05QM8vHoTatfvIizA+4sQ
vGbYjBH6O7FuDxlYSlhq6QTvxmaBl4IZqPGqFIwpkj5ArA98wZnl0vnxL1xJZG0k
Hlg7Tz48EFkpe5EIoMud3YO+tB0fVmq1bLyxc/X1+R+m4Ug77c7LGByXZ0AXpQzQ
3LMQfv3uKi7xlC4n6rAhVHVT91ZFwdNGdyqmYJbMO0sURNqCGKTa3xw0tBY1PGJj
7hfseFgEcni1iu2Tm7LDY2KSQEz4GyNaOtvOF59IGkQax2QxS/0DdxcBK5ED+WLa
diCr5nbFmo37JcGp76/Co1SP6qgrhRDBtXLoBousI8CDaGQco0OS7IF/V93LEb49
DsUVM8AbMeS0+JCqJoeXXt62hNT5m+wpTr/H9HG0UB0BWbKTX3IuIKhdF4E+W1sv
cd2bhwSp5r4y8zgHsHIyBWAT3qvRcJi1pS1HnMAWl9Lv/PfeMIrP4jXZEjGdblXr
RyDCd4YVkSFfsqBXMHcVgjjbX60uWYw8eOsCuaOU3MUlmP8J6iluEOUVyKwBG1gD
JIqHXglRaOX4PLOplvm9/HsDxgkIuYMo6GmKbLblCIY2mF8h+yn+I86RmRhGYyRN
ef/dTugkrlLq0pPjJ0EUgD7XLq6tkcSHwKNHLO33rmkyZCTCDgGwqda3P3Wy27+4
T26V18GFuTcm27qRUZb9joS/VNv3zlmSUieW+0FNw5u7WtZdqThP7Y77VXodpOZW
Inoah2NADC5PoirC7Wnwt43LyJkT6ChdcxulXdiwLi6ZQO0Dis8Z5WV86r3lMtqp
GWFfDRMnoehIV6FDvZ5UyKpn9MWvv/hO/1ZNyzYROcdGefTP1eUW/5ORdEbyOsRj
0a6CNGCPu1qQriRkW/wh9z9uzlXjBN+7t4aD/RnulQ2a8DqqMhPmGEgounvKQ6mU
yPg8vd6QoiZKL4B9tUIJmb01oE0VMDepBwNo1sjR3pTrIYMg7X/I1ZZJNprM9CTq
La2wuCNxsfkERm6sJ9TzkVrGzDTvv++P08q8UaGgvyFiCSlwLZGLX7osJohqQN+G
+jA5i9bBWZ18Z6AaMpHTYnGigZ1SAxjR5neYoYb6jHdYX0GSmbKOCftkXuNQT57g
KULvY2Wl8K5NwfXaB5iyCA/VT3H2XcHmqeIi2KGM3/ADIbsNogrxb0rBImhxW43z
zKs0Lnte/DvuMX0WcQrSe4tgdMfd6RBoSq4ESAhAIir1YLTbC3XLCkB/ssMy7kAE
CGAJwlsc5ymxevSYc4WVXnU5iBlHO6pZauCB0145SgqIej31Om0Ki5nOwIs0NOvE
CfTyc7Kxz3FMyFxizey2oSnn0jpq25O89wV3sj0/O9hPQLOPEqZcisJSucscexUZ
2yK8Rg0XCigdZrnSSqPtiiNFj+pkl0Zdwy+G+J2ttc5G83BsYRVAsSoaALfpws0b
TArBU8L/myOXLYkXEgsolgOvXQpoF3mFUYdxQgb69dGicYdnZdFnbSeM3NazjZ5u
ArkhULqnzdnMRW4JsjmathgtfZES4UERPICEzec+UuK4ylj41/WVVBLvWaBrtEqI
I48fLlONZPtcsDgzeQrPoXCp+kknbGvUlTVW3gybiry/EfV8mRLj74mG5PdwhDLr
nAjjN0xUmzzvVRwFV/Gk/V8Gdn8ENj7jwIZeFSqCHHBAvBLTN78AGsdk967VBiYG
o6tIGsTVDEoRsEyznQucyFW3oJHx6aeY6Ekl7IN1UbCoFJn8TNKcQiRjvViBROfq
1G5ed3gCexJtoxVaO8T4+AUfPPxffXuWfUXY4sPtslApeLZESuvKdiCVPNpgGqNo
frZBeAm32eZK09/g+4Ce70SoKz4bWR8CF0/xc+9wndLSSFtL6nhS28ddYU1VXyEx
C4TZBv71xKu2+Cknqimnov9Un9x4LHGuIMYcJ6D0DQzO501fDv/pKWYKkl8HzxR6
2jcE1QMCbSmxBKHCaiDKj+hSj1ZE+IWjiTCYZuKnI93K8WZA2PHDPQqroSxmBNte
PS4nJzGyuHcbdBI73Mq2dJ1C3rHsVwSHVPja0M/5B6eBy/34CXqHVuTckgIRb2l9
uX6/OQpgMTLA4uoQNtenCAt27+LCXG2IelDoRtk9+r8jnUcuL/Bswm5eXUvp4dvl
my6E+38xRiP9dJu2+fvSDq3POzF05WAGcbNu0EwNYM1RsmWMOgT8v3hjv74Fp2Ig
xnQEFIZeJ/BSf3q6NR7R+/OzGbgIgfkjrrqzCzy4/EAHHgMANrtt1sB1tO+tH/1e
MnUZVlUR79VWKOiifXIFQ7g84Amk1dPQdYB1nx16M4CXsYL/WlLBfILDXVSK+Go2
sA+c0qP8muDlZ1cU8E1qg+p2iIA92PpyhQXx2ccebLynQi84ol54mMNCoj6FK1Mr
U6UCxq7+l/S5J/gsD2QAcIZVTGQ1BT1oXD91gbuUL3C0GLZPseeJBCUbyG0CCs/J
0tTGmBBAGqUQKfTTDbpryDnfJAgrezIeFtGhC1hmTQm9uxFyJGjZ+4kkVspCvtvL
e57c4jXP3++EcU6ZaNMbH30wG1b/HOpUT4Aih8e3EXMc8oQZNpvSTl5CaKUMLFng
GG7uwNy2FCDoF+yvAyUkazoKw6IClfERxsXw6zeekTN5R+XiGC79QRrUAhkXy9md
5V/xuiYrHZOV6pBclfWgIdjyK+RyKLo2MMNyLn7s+ty4rCKhxPpNLMwPEQUgY9DA
RT6YDEp8ojlDeiIrleJcGLbXW+RPeNI1d+ZIbqOctdZEbnRoXNxi2fLYM0k49fvF
JNj5waUNeVBcBWXoEv3ZcXELNeOBVzzFQJg6TPcK52O17bg+X6X0kNR0uHdPW068
mzQ2jyawTS4y3WovcpSFVIhSRgoccqP1IpdFoCaBWL5Wm+FWLzLdvmiuaHsS66sD
3x2zkJqONJavpenxAuBCBxi2zulV/282pFhFcyV3E8TXSuytMd52Hk1umlpDrjM2
fiRbFUBHhbh3LPIj5r7oQpl/w7uSbQfD/rDJDGXygm8ie4Nq0CJR9SD4R+mNWKit
uzjYHcNcKNXp8quKzpzqotmJpoe3nChtqkNoXXdyLf5aVHSbRkd368LUlMUJW1Ka
hUbBTx3iQcKAP2Xf+fV/3GGQk0l/D5wpAC3+50MI+nlGYtP45lqQiXDBex7x8NrV
u1abf1uWFOmY6yjo1iOt5VdB80aXzneETJ8R/7lzD8FQNVjwLJuUzrt9wP/ghZwG
2EFXinkMsa64/L161NEj8FweRdvN0BhuozjAf9YZGzTlw1JZbjTQ53AYdvvA+LV2
uc2otrvwXwGzWslqaFZnT3sC8296RkGsz5z9Iv9ta9wFaQz51JFxTfHvW77HDqwx
0oK1HehaA1NAYn5UIRoZZ8LhSR/5w/dRG/TX7KsiRTjeiS7A97ec0uIED2bdOqr5
5ixrfTjFslYz3s9T+I7O4Hb6E6ZYpJ31z1FyrIFUPSIYwR44P2KdhToJpwdXo6if
t8D9KU1KSpB8fHeR0Y1Dc0mmrh5iJSxM3ZqvJ9QSijxP5lOSQ+f3EGr15CvkHHil
eAm6hmHvgiJV5ta/SSS1CAgDJEzxdCt7JqxtTVX3D45QOlBOxN4ANcxrmwNAou0Z
huHOwj88T8Jfx3Uj5fRjDHQ3LwOUiqq8nkIygJG/xxzQILAECisPYh8ozBrbFL0+
V2znQC4XzMZcvWogj1h9nUrJQxriMLUM+JWVAWveQff0/J6B471pAA9DBiXo3QQB
Kb/SFxxuUyR7i51tJLDlEQgDgxGTMfpgjhgARvA/K7p7QYFsXM2zjMmjyE857BAB
5SRqdV27YALuYpQAoNGtU4PVhoesqJQf3N9833wF2XIC9Qv13Jtyrk8J2l9VvUEz
x3xTR2mJgt/8/dR4m4DUmATMPG7Lu66PL7s/Gn0GU6aKUsH54EFaHAAZHL+dXtiA
VX0jQE28d/r3p8X9Qa3QgrArfjmhTNXQOolUELx9Jr9rz5JZgeDJIDnbagnWZO4K
nb0HHPSvlfRDliI+sPhyopiq2beDa9qG4AYiCm7uJCLhzs6VxgH/froAfyTOvN1X
qDU0u4JeWcqz9gvA04METwo72hA9IBsgCszh7lmzBcO1GDYmRuydLlF52J375Mzr
GszQ2rMmBMElgxScUOd07pLmwqMbFAEBGdlzgykFnqBtQdrkdyYviCRhJlgqzGKe
UBPCZwzUDt5kfNeJ5dRQdfqh3hgqbFlBNx0YzTtjmiJl623toOSqLFAzxpeSb69w
ldza1/5Cq99ZDUeEj0ORJmSdv9AENt6ZSJFy72WERQuYyRpvZzWGP030l177Nn2n
yJTBojLJYy4pZyLXzU2kciBe9/pHZyUWgFpiHarIk782NqTnkDlSf7uDEIoyu/YU
QuS5UVb4INsTheVJDoUHDRI2lPorJeHkZzIHOEiTaK5FsXLJVpP8cgdIg2LkoY2+
Ffh6VrRZVOtZqxEvv2TEy0KnyhDKeCZlecngM2nykWixLavb5+wuzmgFPmHGHr10
Ggp98U8S6e/wSt7mTs/HP2OsrQFFPRgXW5T+lQx377Yu0Ksy103MuyoKkwLd2vIW
X7G92RL/jDQw6DKAGF6ODChP2T2F7xbVdFBOWc3HesL0qZsNQ7akA2eqO2WnpzcS
kT+XdvnabIMctlL06bHWimHu+D0NrSycrbW1hydVX+mlXyngvCEVrvv8PtqJ7V4e
6VlPeCjvD1zws9IRkcC7KsGEbU2Whbet6Euctmomlj5MXNzBOGAhcATH+w0srfsQ
Lc6bqEmogrhWYW7UEm/fNZQfdlOCDMd1mdN9KoV8OQjo1cdP79Sz3F3utLQITe+u
YGlctRZ+Yyx7auIxWfv+8sHFMs7DcaSl6IEGwxV++qAoRfgjTYPUwDoNh9l+8dZB
7x2f8cORqVdVD7p4tCqAwSciqOdBvdQrsRWQlszY390V+oo0+ZlIG2+EbknFfK84
ozKPdZoQUTteWJYp4GsEhLucuKHZ6JH7Ft6SxjXpjAZ4sxGB3mF3t842qFTy1R3p
87p64WDJdk8IDDzC6QMiRpHtRUDPm3ABKT96PG9KFJIDoPDvf6NC6MWbkmTW2hoe
zu5Q3dAgGfs8n2bdj2vyfhST6UreQ8+1+3V0cXxFSdO8PSzjTLwx/HlfdbvcBL5F
RBDNLgSl3Qs8zmlZPI+cn3GZ2QQ8zelFAvxmaIT6GMZVmZo2OQAJ1v6RXYFT8sxz
OGFkMYNksdNmf5r4cCckuzLb1IAeRW8I4FDdLdFrRFgh4wfntMag6/ulvAC/ZNFA
YwjTl6JqXo05ZC00yJMypxPh5OMYSBlyZ3WOTO62AO9KUKaldiTsIKG5fgmEY2HD
bMRX4qkM4XDLLeRhHLhLrXeYyjy8c76zEZmtH3b7izWeO0clES9f6vAdDO2IVZkH
HtEiC7HTEIE2Ve+R+dxWYzhwb0bM4PPcnG9oLcp5IU/Jjq3GBva5Gorjo4Hv0D6Q
is69fw9b+sHOmAY6whmP8DFbsR813lx4ED8ljyqg53Fpbs7pDuR8Amf46RDaxBX5
Y68/p3QuuRoBab/CkC8ynZARIaYOqGk3b9m4387AMsBevX4/GFu1L4SGmHMbNkrD
rdqWCQYv/ZWFel56bZjUyQmdF9NoF6OZBi+b/W3ElwYimXWReLtfp1PzFYgEgB5i
yGcUNR64JbQCwf2idQDHEqPSfsg2/4mxBTsjAsJvX707AC4yV4xHXSdpiicUeo39
MSrOR9+wSROfXqFsrDzhSzH9Zg9i3la/w99M95/txXAD352+hm1cBHHStlpjn/qj
LRQN9xdzOGyX/UamkEooZvyd/JOQQwSgpwCxg6SIgynqiVWXx9HhywYNcBizLsEK
xbo4LYjWGsrYw2Ay8yoRZ8w8XZ5CFlzeXjv/VWebPwg0vboaHPJq6erEllhZQFMe
0UNlnfrYN0tQRYxLpss0oLGzYq1WkdonKY+wkQ/gvarO7fmkmG6fcctLKXsPM21y
lCc7RBlLLo/w4UVt2JnFZNIV3r1moRmnOzOHVbAIFvBhxXiNnBbOLtYOXLB6QfRH
7EKCeb6A56DW/LlDlT81TXBIwC4DPq5GDeWnctxvVQsP1f219CuO/Sj7vFEaZDGT
VcYjGoCWtxvubgcHVAznfG1VIi+JQDMimBULkq5D5UOZTwdlb/75zeBjxB5OBDV3
ki1J71ZA7V9H9wmJufvBSibzJj5Bcz7eP0I6dka5sxR71/nLPkZxr2+Qid+qwSms
KShm87D1QbbTm/famwv8zsQ/sdpEzw0cua4dcLWjy+M7/r4eT7g0C3ewgDtkDcIX
YyIlUu2hThljY3LkGEJfl1pOmFL7CJi448EPNHxntCggrZKM8V0yOY0f8Rz23azY
EB9O9HqeM+GO9D+t+dl3LqJCsA199qvUiQJ5GiFmlEaFdo450ztHMS/7IgmY+FBm
EAP/KzWzG36tIOaOmVG8y0iotcTWTRqoP4ZXb4gd+jFjA5L2EpMKlOlwqIwJew/b
cABbLDhJwbiGkw8spsqVSTOxc0phXlh3tdlbu4QQVN0eJCNNOLHRJKbrarx6V9JK
TsFs4RHCCt7vh9VwxX0P0jK2cOYsOhkY6H1vCU295/q6b7Ns1NlaEHou0m8DouI+
MnvvNpUvcy29ceDz/36grUuwfScKFLC1kyy56c6SB9sHpo651/guYT8VzFkmFwfk
2XL0n/mzbshvQZbryAeqRtmFem9WYmq74ce9FPHqzDMDWP3VuZ/eeplsISVrBfmw
G9PoUfF4mVt7bbHZ3uIJiFvA3q3BO+rXCVkfctDezNhemG/YTPpbXeT8+KocPBAl
fv2voywhSQAaLHjUwbfl5px93K7NcMTaobWfbczN4TkEzWF2Ue5zurIUH08P/RpC
6ShIAM9X9lC7JasLEH5p8rYupsYSBq6W8ItptOO5H1X5tOJGg5WNG1zSWyhocVZH
nVTnObWrLmLezyGLBtJXzR3Uo58NVZp7/+BVw/KhxoiLpVPwqXugqMv53DaeNr5G
fL4sVOi0fTIboePiOU/2BZOJtqU3nxiQTfDY37HoWQGqYj5gmn1XKB7dsNCrMqlm
+jFHmcNVS2+amD+lK9RnqERh36fezQOAsO3OmzMbeN191rFUs+11kIytnAazpUCM
y+yqQWrIJhq7K9mUxTlTeeaxvkZ9w4qLaU3+1eK8xMXjlZGC7nRymXY8DMZlYw3l
xHox1XSGWcESsDzbL2Sl/0mA0RcX8kD22wVEHzyXEJe+11vxEIC2qHTKNmcPjXqI
EQAh0VIXZa14+MKU6YlWlyYQoNjSHfojbD3roPFSh5NPQP9rz7ESS/V3mYdai4EC
hnv4aV+vOwEMubOHV8XwvBQFxydm6pPEtH97i7p/Wn5VFqFm+B7rPtI+7gVyqe2g
1DfdLyQv4gtB6SvsH4moyWGp6hmhL4NKJejBjRzUwpqP4TsfJCDLc45oYH4gc6uc
QikrOyI9mADHjO8HcO5fPF1lhcn76k6QppOrhufDHVN/1Jch5XqVISHpAyIdn/6e
cLfrzcmXS0F8CiPV8jwo3hGRbmYWCgXJQ/jKAcS7G2WvMXmO66cPAtB7wCWYo7RA
EZmVCbFt2nd465+xwyCUTNnPHDf8iJE07Uu8S9/jRh7kTBIB8Ie4E2dcuNhKzZQ9
AwFDYq2STZPsiCqmbl90jKYvnk4mg8PlwGj0kCx7ohsFHhF1tI1zgkg+BB52bUek
jHteVOauNTfPevmFSKTR4KD2B7jCMUzu1/MNqRmmjkvWBWtKumKE+amCXb/XafvZ
jl+psJ73LcOQ/Qwpy20OkEyIQeGbptGDTbLqd8Yv/E2Yl4wuP0+3zZataADWibsT
Vb1TT4gB+v3R37XWjTrNGxMamHG9Pq7wWeI2OcKe5IdW0qGUw7ATGPbtjev8XTxB
FEmUTzqltfDRNA+UYDxlpoRV6jYN22g+pdcjWQtD7CSLqBN6p1sN37iN3FRKXAkv
v4J7zkhnfVRQN7LzCupes1a2DyTzKu7CZJ9nuFr6fQ5xClJP6a2L3qJMcrVbLi+q
jBGWymaKo4D+zd9BwSCEr4makbB0MxxTGRPb+6cTBGY1RQJYF54HVm/LzSMlUCiM
ONJUwhhFMgnazd9kJwiBF7VbpGDbyPZDm0lf2Ysll2Ik1g62JGefnl2Ny5Owd+Up
Q9o+GgGx+MKUoLKVXAjCFUN8MM2hjqst81YJNttmPTouIl/GwwbIUkqIKRjrVMI9
zIYc+tb5zBuYibOO87PZfPN1K1FLF6uvP9M8S9mUMf2OZuo1DyUGLHcqQEndxNM9
NWKjlIPVnCwZZu5miBGGdWsmhUCtPxIusCZukRP/rqwXG8mFYEa+SBtXW8JZcGHC
tMvzgwscC9/incPYKq73AbW4yZ4PHld8HOlD7lvApwr4BqaHnZ3JUz1j8NV8yLL0
FFjUrg2l2d/VxoZcvP+vvGBCPtDB7TwPXMDkGrTzKJu491DtDUmahlKyaL5XLGzW
swArhU5zo/2bhnoUTK5DnykpOj6QlbXb2e5+7DQdOKOQ8sd51AG3vO7TaR0rCSe7
`protect END_PROTECTED
