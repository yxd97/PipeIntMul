`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AZ4kkFFV1x6Nkl9H6TN/Vs9PoEnx1QvbMR4m1wRKZ9OzO8zAEywn7PXVIMeGgE1C
PqA8uaKi7ujWnsu+xZXmAcsB5ud91AaHtRACH/UyUt/n1u+rqVzB9McL6FHXaM51
TioRrYbOKr8tmiBN4IS7gM/H1GnRu3g4Pw74JPoDjLRUSa58ubow8/v4IxbuiWSB
m+mqIjAEa3mON020JlPYd2ndj4eV13MVIeLjbQY1WLHpJxz1truQ7YY3tIrbFEZV
881cVzSwbGC4+2+tUSh79sSbodqBZzRNKd/KsTsFmt6stYd3MBbth9ujS8vortLE
G8wWLXTFM6F3xKNHS6Z7XXWz7iMj73gGG9KaflCeemdPTx9DAlfrr61stK5CDwXA
aZTsKZXM7oF5eMpHMsx4Z+thGYw6stPTGlJBa02E50BSayO+5ijNaLDqoEwXjSuE
EoUW6YqqXyMb/1sMFHsi8IJI6iBwAtMmB8aIHUrGzmq5ky47sBJKUZD3XBzuUmmh
Of+z4RrQMkHsx6dSGzn0mM4K77+q5KmpUDhxozh3BrGB2RurVKO1Ktxm0P+kpVlM
bhh1VKF5ysQv4LwCPuOYm12r/ac56PjWWwXRu3o9Qe0MMlKCHuD9pb8XPZMiphfO
ygqyLL3c3nMrc+AsPSoZZ6hDKl4kfIF/614E6pfCPoyjmmiAVJdeLC95knucOp/3
OJwkAphuE5DPQY0gZ+boKGd0xVSb3cb+ZHEtOii0O2xsWQ2gO8TJ0MqiCE94sYZd
X6EWQTw8qVLwC30TzZ6Db3WvhNXbtoOBMEdE9o9Q83wARIr95A1MI/gDkvQ486ZH
t0rjzRaTCJb2Di+yl00WVozxfaiirx0WJpG4U+5iUWy9pjty8Ifo+E5bpmrELRQ1
6OaZHfdoaQF8fl/v7MFzHSLPRvSK7NBNrWU5a+9hsHf+2mLszWJkv7RCwLHvtV7L
Y7xpQegHCpoCv63eb9zZmayvJpoZNp43piQLUZUACIf7dZJdgsA395G5sZxhwxBP
E6NhLL6MrGseAY6ZeRRoy9bLGH6oHn6jPZArQ7OLPYA5qwh7q3arRrVj8+16Pyme
NpvS+UXvEBQVdY+4ArUgxFJIw5QsG3nwHOmAe5oHDtd4ui4T6QIidAwMY6wrlgIy
v+2N/dGrac1LoiPfZBtuG4C22NpGPJJ/cshUjIc3VWFhT7LcH0NFCGEk4pBqZjDa
fFLcDd38tXjaWB8+KHS0EpiZvzmoWnhHFGJselSCY/r3+5bm0LTWy+4UPjTPuHhQ
dUsjG1oJVADnSCsK977gVj3WmZokWU7ubtdClL0Zs8NtE8fX7ShTT45KKpweQsC8
FQJ2OmoiDstZXZOXx0qiTuccLX5qyOA19gw9kLPzrPE6Lo6BPUdUMgCSzG7SoaQ6
TVdh4WFBScLVaMjcx/pstWO4TKD2CL0O59hc7gMioOwDvLU6aw7gq9UpAjZD9x3S
bbELX1YFziWI0ZfgvdAo7vJ/tt9lpjZn3wvojnJ7S4hcqhRH2z29RvL//RjoEeJB
cCoaVK5Wu1ySUJsrA7KimvdzAUv3BCDMvxCaWKqIGkjbLs3uN83qYiBVR80N1I3E
6Fo1fomHE/TdpttEuiUul0ZAPwNLU+lIx3y/gbwMreTyeV3IWWxDbYwwqCaY/stF
DhnJSxv3zHP0J2OuYnpek/PslFZAtRSW5De1e86Fit5Vi2Q81qNjPR7Cs6AgeF/6
v7ZgmHPsGE2FwUknK8hm8j/KotDGZ7qZftvR+5TzsTXhlzlrrOV9hu+gyL4Z5a+g
IqlFljyVrsO/PbPOuVqLkDasLfw+a/V30Y4ogU179Lw3yOwzCD+/DeR/lIocriwK
6w1LHsmIqPO+blw0jPlfm8X6Wcx4Hf9Wh2nRHFfzplZKVmpLCoouwP7jYNj3lAag
pQkF88+oLY09inIc+0+l0FOf7+PAPRTQxZcKrTBas2rJF1XxnrAlMigavP+oLHCR
9NeCXIbq/IxgiwFqklFjFl0rdNzusQU5rAIA0XP52H3XYb/IW/EjOBZ2BGX7S4LS
SvtAO5MtgltT7PfNDNc5TMQlrKtxnZN0CTY1lFberJGwCefcV9egueRweFg92CEa
fwp0DMB8QYQgSoVAB+cMS3L2StRu+lbHomX5OollHwWpl5m+AgaWmjPaKym8XYtG
+P2jTR6OQEf6XJzR3urCS6ro3GQrVC+uifUiIRpugmjvWlMyrhfNfV9lOkkTppr4
p1nvWyvp4KBIl68SxplHYyc/y6BKvgR+BX7HzGntsEyml+nEXhcnmxOSDVM8FO5W
b/FqIz3TNdiXK4xSQnkYuoTxXvGvpqvNOpdlUIXPAqMhp/+U9129fg0+vldHJL1x
Hp5GuibkwD6lVYD1zM4R0VtDjNn8MHLR3U1EUwrMdUjoIwSfGlVi9vnRQ9cto1Vw
CfSaz4uMwqk+AFbiORgXwerkgYT1yvzgeEeyBrlTRnwLQtUXcgCtxQu0xxz8JOo2
ANJYmLpUyKiidvucJuSuYv2UyV41gVOZJHrJe6y7Z4Wb70CO7vXx90WowH8F7nTC
zu3z9t+LzJVo7phNpMTbeSbP6sjpaIyB5cnhdFh+hIWCp7LMQISkgdg0OXaxoxZn
U/kqSgzR6ovEgPQcPM1yXxTImu0lb0zmkaAZL29SyJeOmnkzKqixMeKE84OV+lMd
8A0BqOjb8eAYjFFLbBrRzJH5w0rYN73RemkQ5DbQdUnSwoCiecEwHLtY/kHbnLEt
YF7TriOIvsSdL1XAca1bYzNVxZG8o82vkJdgFAV+VabphgR8uqUoi8tAaNLpSEK4
/iJHZhXzRZl3YTqkWqx5XByvoPejLBfirkda+KEFnZgpvi30CMilaIbX060H5EDK
884DQuUha+dDO3xufM5zya6k+DNAMVbPODrv+5F5+pvwUeNdxUSUtfpjca6phaWx
Ux49E9aQ9aH8162Ua03v52BGyjiZmsPM1ZbJtNKBx/aM9d0q+0+3QuTzSyDWiY/Q
KcO5gb1/Wq1LB5AxUrWAaP3vawjN3JG4ZMhpfFboCvIb2ZVIufNu67myryMgLytt
UV5C33VTyIFpADE75sWsdzvy2kk02M9Y1ftR3Rf9pjWpXG4HCZajAagU7E53TYvO
3/LZ34RSzRigig7QNyxGRHPiDs66S8CDyqj3f2UWjiCaK6onzexIB2CmdclO8EuN
/fnr0m6WtPD1Wk+jluHHpOCOYxW07HamsD7yzErM8qmngVM8DWIJCwSo8gpDEEpf
7eTQ/1dyTrDNqvZN9DUNSN8QYQXFzTcTdwfa/8dhGb/tHGFWsgeSGCDwqnidtWHJ
5GaP14y4rFEwgLNCJ6jhpXnWiPA3Y4NEkdxwOPANQ3zV3wpwv+WD5BuvLwiq/FDc
6DUXv2Bcnp3Jr6ZMLTsJLjJjfR9jLZpG2Lp/uCwzXu94YOFJs2kgy84tgD536WnH
6bMmmlpRiEdXgI6Om4dp6yagmx6VPMiNRoQ/j3UXdakzU6t5TZCduoq2CxdkLops
5r8RivwVPPkKC20sahkoEhGx5qW2t6b5MD/fE73UPr6e9TlVRpDnrhBrJcHzWsqz
Hifa2gpyPPU4Me/kIixrNEweWCwdegN9fpEpXI9l8r4JXSuX4jyUt4dWIzv2inXq
z1rF/JDqJkVr2YA8YMKs8tvE5CoMzqqRsf2L2g2YP4c5pdBbZsMOGFfQeurvPbsN
AhPWFmBQu+V9Yj/frrtA+cYaRQMOtz/xyIRPLvAD5NsotmOOeKWfk7arkQPeaC1w
i84X+4Jssu+TAfLtBWjHgnvN8G7gqK8iVv9onOcwsCs=
`protect END_PROTECTED
