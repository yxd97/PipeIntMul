`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SjCyrrVCIcJQ4F/DF5CMaKev+HF5Tc1aGrk+0Boz84MMd+ydVrIO52trlE9mvpEX
VzBJiWBRTvrvtTIgFd+4fiiKuIcwjL3mi5kqdKnPCrRYa7svyPpbgnE0skh77bp5
/Pz4ulIcMKoHAjMMap34bQ0+fqDrUkSUbcxx80XFiik2A38kbxay4ie04V+fjXxJ
SN6JHCVlWvlKQEzH2sCFD6HMPnQlm2jDsxUAT29cb/6MlQ7FwCbmBxanSJdGvR1K
KD5HEt9MDOODeA0M8dG/UvKsa7szs5b9Q6Hod8D766c=
`protect END_PROTECTED
