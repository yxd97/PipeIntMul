`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2wP+NoKwN1QeZXfSy7ejWkNlsy8eTZ6t6efiqSRH02Pw1OovPgDYnwHzU8q2uhY
BWcgV3RmNuF5x2dJanLMqE/mbi0ofd6ma3iMMfmehj18U9nNd8x6mq1eEBeDNvQ0
jwsIsIiswk52pQovcTACJcMMkfgop0xGTFbekIbF2Qc7lhc0oqjjZFxCPrsil57P
h2CAry00nQX8K47cbv6LIB+PxJxTrM3KmoQMfpdYfnJzueskOi5ljLdkSwGcntWy
SyqDrExo4EIv90k2RQ1mztiK+w7GtALP2Jks0HqzMAeNOxLjemrxBwc0hQy2LRk0
u6ERyZFWs4NFxILVWCPYrPP0H0jBtOPJOlpOIdAlibsC5PmkJyqZZpXPXqs0hBWl
JWl6S+272Lqnd+tGllhY7T23VNUBkfY8SDcQeApJTHWV/grh3s9oQaBH+uqsnvUc
Ah1CIMhevQ7ZlScztm93Eksb0+moQ9yudYZcOkTqIhOgWhMiIzHULMVGaJLcaaS9
YzDu+yokWriFunL4T8rgh2c/Fr5Oo+vsinl1wBHqkw+6bOdai9o4Jls37a66me8e
C1jjYocWn6V2V4LhgXbXqAD76op8TwuhWymz0XB8yX/YWK6zkW2pj3qRvSkU9Gd8
C1grUQyR7SXs5OxIl1tZAGwmPAv+QdpnkSyIgDl6008w41IoANpU9C7QALnsced8
jbrjAMaB/mOZXFnrrJeXhS6GGYxgENyGvxImM2VJ8R+Hl0CouVn9NZFrAWbPn/yo
ptZbSs9EPDf78VOY2ydaj4MYUNtwds4XFymJusbYIbfieCgoB3iDPp3g4KxgIhNL
JWMISxFKqth4PLpBrCWmbIAxPt6KZ5QTA/HeajD9ayigIt03DeYNch7Gy/+0RpO/
QKTfJR9gk3p/fJ57jMsXn3lLT//0ayCFDNgGPRig9JuLmzDDuf5htmjikSBFSjgG
gnixNhtcXbMp4BQ8jSxAuT7i2ewDjC4XSlhDDWf4wVXBya1h3cDDMpYpiMEn0uIW
Pqc1ntjmgrWDVISVt4zBx1Nq1iQjQ/P2M4N2RgIPyqfEyBi1p73fgHzqcNFy6WB5
7vSWeL7yA1vnJpLTS4IUrkppwWq3WSTJY/E18HgGCPNJsSnfbLl7CctHzPfbYZNM
wiT6ccpC2SxKJz+NbHxQOL1tBG2ujCaET3N7l6zcEKoy69bUWAsQltdcRBRsjmdY
+JDz334Lj3tcFc4bS+NPIz+kiK0q/jZlbBOT9LI1Rj4fVxGU6Z5cN8AwoTL47qRB
6BPG2zc8QziAGy71ZJcHBHzbLTn5Uxtf+Lazgl6DAG5f6OCfXytbAJjX0Y6lE1rn
tjnEOphIP6YbXorZU+3fwv4WR4bE3jTzkhEdiW7ftkDAV3vzX7Q9VEqPDHDjiGAe
Xpu2e5chNwtnRSp4e7UHIA==
`protect END_PROTECTED
