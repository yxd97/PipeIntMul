`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RTedAdgo3BDN3UOJJfjlmIVacTMbB74zpts2RiKokxxRDtnWRYRn+b8Q/hrmMIf8
IW0XFKZZyKE2phPjB4pfsVHZ506IlQ8o8U0zuUKLE5pTS6DiXtifqwEsNxOPmXxE
XHleZ/IjbOLGjzAG7VvWQ54/wlakGFM1yDdgz5e1HWKD88U5KUtB8+dv5vFlsfQi
3wSDPoBMXi+5tfkvri5NMaiJQdP0aoM700m7emy0By/Sm4dQGm4FkSlsj1PA0z2P
//aLIY1vE/a1Mtsk6Az1GWKQlJ3xP7gMznd3vMT/rI1JslFlxPwZptnYDGXVD+VD
kZPAXmXpx7Sk3jpvMts6JfHfLcKOVDoyvNkzNRFiEs6Z0XqqnY8/n7EtGflHhCwe
pzv5HxVOERiOnwgWoBo0qCfWTmYnpc5J8sHDBVcQcb+FX9wxzvnIoFThYPfv0Y0M
gejlQOYGownXWcuHQPaSNF8ubuGGzyv64HH28OkrnwhtZsAXd0W0eOvf3Y3PRqYo
HVXfFPxlu8v3k4n+yaj3ELa1J+9o+XUnaUD/UG1oxzXgFlrmIJ2kil9Hbe+wxiHO
wcEHPGhPkp9tBpI0UTKvCbL8T4E1vy/1yXExpimye/T39iEkKEhlOftFxamLzM7p
EsB4vF38A8v1rcZQdbb1NTQyanM7WiJ4huFJry92AcpF4rlRLc85qyiRNPYm/ZtL
D+4FsmmiF+L0jVa5OXDcObQVmMoRueuiVm1tMP7XPpBIX/R+omr6kT1f0/oen3c6
NUu5tWBVtG/H0KDlacunZjlOrEeAV0u9zSssUlsllm4MWRBBtk/bIAw3W5v+XA+P
W2BXHrT//hlNb5LjIzCuni8awaou3GFV0Mgi/a+e5BJgNHBohyltQJswj/VbKlS7
U0tBoJVd54jiQE2JZLKtCgNdVJJX4faMBZ1xo6potsc=
`protect END_PROTECTED
