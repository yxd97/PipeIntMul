`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Uau0bghr4BgHYuWsj4c3mXhnp1wABL5yHxVNoplWaA7G2GkiyOhSGBQ+xWSwlQx
SwxHyRNgVxGk/j0h5Ayllwgxlr+E066Sh56+YqOXAUwGkxxrLPnwwqWDZACfu7Zc
mYtoM2xQUsrhm5ZURLYVlz6A2RPOdLQMw0zMboxFuNNyMB4snWCgcbJBnJewV1n8
zdAPnBjvXBxjPMGhJAZn14IWJ7rlZbEoAemGghJHEncfWHx87S31DcbZA8mu7/WB
qPamkbJglv9M0EG6kcRCTB6Hvpb81yiBTE1FkLd8fFq1pWor02xvu7yhhO1g24rK
r0/vx5yBoyoOUrbfqxx7NuMLxHaDN++K0LCmR+bTyEGoGWkTj2jw9CvqQOhJGCbF
g5PwmQS9m3D9o0bl21O0ZIDx8HAGKqYfNTSvT7SYflOF6rXM4tMFuWOp1nRbuWMd
oqYMou2zq/NvrbyECh+aFPPI3tOg/LZFBfYdJxXVQqDf1lE8ht8rpcgZt+5SBZJ4
C4QqKCFpz3N+zs4mkFTNHoYQw8W6dQmloOqv7W16BMkzobSNM4/O2LCZ2rDZv76K
sLB7DEAAl8vi3PxuLvfujq48r/rpRnwjZvPzgzsy5hU86eVDNAkw2XsOKORjOZEE
iWbh5pR6wxrIu7FYq3cD7EwkV5dDteuuajig8o7+sajaDlBISaZaIJWAc+b/QwYZ
2uyGghwerTFCSwHJE3/lVa7FY7dDcVP4VGGx8jr1w0xtowgOVKi/1tvBfh0MYNGM
S/Ftq2XVro0Pv+TNqwK+x+2O1ekTkYxwFMPb71m1BlmculLC8ZaGFqljtinnG5+e
B8ZtB1AvKeV/vjumjP9lw6VTZGRzFwY6jMdZpGgTEYnRU7n2K++Ep7lwoOtCXXAG
DTXLA1JddG4MXHWgKozH1zUVBQFrwE/hBR4cCmAKtj5M7qBthBiqilWWrtjroXjo
xztlCZm6xgWIAQAu8uYChb3Dl2SqZkIr0E/2Wh5rIg4TtogmslviQsto1rvu62xP
YRf9Ew6ITVc9oWLy0F1UtehCOmzqAYTBrXkWaVLN3truOXm06aHEk8JvzlwHPE0U
x5mxJNz1H5TEmU7GnJ/icBR9Gi50nhfDVY2QQjzukEedptQSKiugcwwjm7yYcmxA
rDNowr4Xy63V8RY9prTySv9DQKOq71IObMiQDBWl4r4mTcQCVRjqwdZVPQkVQuAp
V0Rfhy49d/UbMoww5DvsBXh0/loUOhkCJDHgVI9YIffXxyFiRmKMzweemiWyGhCz
9LO6AUNhtxoYfvnxRTiy8pJEzpu8MXDZ7wRdoLB0Arnyq5sg/qQEIWRmApRUvpko
pkRb4qhHwYU9uoNuOFMwdOFiRhs7aWoGiSUYzSK+0pniR4aMxcp/l8lsS+dB4k7R
ZZt5scc648cqWo42v4uBWqatYg0l8TIKG9t86MR1VEav1RcEaJtifXaq/uOKzBgC
A+heTI9ABCck358mveXuQ4B5bnaKTzkqoogrmWfWJy9DM3/HPMZ1N+NftUCVyBgE
Y7Sttpu934ZFvvN7581oNNkyuexOjTN8mRdtk/geOKfmBKsbvyHm3OtqUk4qiyLO
vzDgSY3iE8tlZdBsEqXCfYTUre/DDrQ/S26koKMFDWM0yNuS008H91068UjuzsJb
YA7Sk2+AVrX8WJpgo4xofUPg3DP+UJncxkXE6l14rulBH573mmU0zSGdP8Xy5MJu
Hq5oZhccW1+d/39vQZMn+sTR0wNLkT852FyeedIgYP8RbFZjxjzI2QxDIw4gbkbs
DQNYESIigtADLe5DkXKb4CO62Q2c+CJe0vtE613reLkmPVekCYWB0E2gdFYIleBC
P223TFKZK2nPYR3h01qyERfKVNqgj02l0NV7HaidHDa9I6Kb81MTDj1uTeREY1BK
dqIysOHowAWcpdOcZSOHS+/beWN3Hv3j8l8DCKp63nE/WM+SHosMxxqEOzqi+0+C
1bMNQaF+VNS66Pq3YrvREyJJJWPFueTpTtlcVfNfPQco6uex7tYTWMTCFIBSjY0Q
qsJ404jpMOvqnJWp/2qYxlFhJk5H0RtV9ZLg0ubUjN7sQ64BBx51KNqBEmYTS14N
zGsvt1rvyfRkS1ms1jFO/EtPBGBEI/zfIYoIQWFSZ4QoDej7CTnKCCMPhoj4AtIb
FOVwOy/afIGI07zM7xpHQwViNVWqiiM51mUAHVcC5r8C+vKH9nifsxCz4bd0HWUb
dOqe3zHGq9fn5uvEIpXUG4sSMfVOGUWIwjkLuOANpOs71Q22PlCYAAqcalku4UMw
0h0Qxe5YkmON3cj4lsKVIRondxbhy9GDVz79TL1SmXPjZtrIi7+9f24IcEVNqHcG
7H82+GLF13h1flcsrQUqGgSSL8khM+bIceSeP3lvKLFNA8c/IbN5CWHjN4bBAUss
wQzKwI1JJFBr3BQK/QBn/fC4y3ifRj2LaT6+W3x10B18kUAqZ0RX7v284wFiFuVZ
A4pfcQzeo75Vmwu+R/lPRfEGuxIcwx3fsuXYwut+4xqVuFHVRBI7VbgEc6v0+3qu
7ysOSMpIpwunoFHreRw6vpibdXHarfSxwAGRdi4FQtatqAYT/8FP4nFMslPnJ8Yk
IBMJHat/lGhrFkZVao6SmKMBmpGVqlJz2W74T0WAVmIMmm6/3Y3ADI9ymdaL40+o
3dz1EhKZ5PmJONHR6L78qbhEdhlqnSPlcJKtwh4O7SzxDrmMLr+tt8JcqOh7RwCM
fPLfkrJymhft37mdTeVi3WRa7eiG0wTb2NGmNecRyukge6CzopAz7OUX5LkXKbyP
/lVuaDh1cO1GveiNbL3fD8d+SPlzotdjkTqGQoikx1bLm9sDJFr3HHU1ygW6XbdV
FrWTAW7yArhqAdE+vy5PoyB85oc2+YMt1M03BsyeA2sE4QxcjaX0txF4M/RWln++
r5c8jvMxVUSK39TS+80n5+Ai2smiNhc0O7qo46UTB+Oo6Pbotj08N3wWG0r5rdv0
JYJD539XC1LnhwfJVecC4eLZg4UBXckxtMVQRUleJVMj7EUalmhdcV9+5kfBY7+z
0SvGeB2JFHu7WFmipNWGlVv6f9PrPq/QUHLMd7Hh9D/R46Mvv0l+yumwTJt8uLkB
d+Zi8+LqyWvt1wFHI23bXJZL0WWRt7sYlCW+rqeeCngsqB353p6dAxMXQwxcuDX8
peH10p3fqiFbLawa4iJ/wCvLbkoyT7H9tvZ9juiQWtZ858jm74uDTVRMuaHab0Ik
t8T4LnBW8U6jlA//F3qNEeLM1hpw60SX6qvdUW4Ztr29lCl47lw44pfY4AptvRAp
/5kcFozOdbTWZuzvIxasR7h2QEXNCU1QG6JzLVjrl7b+nbRI+3bCHVsuuRn9DWBe
Fhy5de/ndpJKczvMEGwyaliQoMdZzr9nN/kZ23R0FDE=
`protect END_PROTECTED
