`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qP32OmoyRPr3KbfT9uoqKVl91X18UZDv9Jc6h21h8lJHtH+JSMEQEvOn5E7evPE
/AHau90BZsRtaE006n70GGuFjpQhcpHuxXAzbS4EjWnhkiisKevLZbwdDCiY/hTQ
BX19+zYob6WqKNnY3fQvwZlYKOLKKOG8TcfcQHNHWUbIhG8HhOz+BYcil5JD+2Ms
H2Wlqsf5X1BFs71jvIO6yTjlJeIPGBic7bCx9wpPEh2CMQE89JiQf5/rsl34zL48
TgTsqcusAA8MIx3/P8dfqg==
`protect END_PROTECTED
