`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogVtCy/kXCPfjFtTDyAsqLl1J4HoZ0oubWF1u5QFNXyJxKwiMQ6hkQq9RyVfB0IW
AbvVAXC1sxRkLks8bmIfIJVOcHoKr4ivByDfjO01Ds7pOKlu1KOi1niS0fxfh78R
J4ZLtIio6AV/0WMmau6IE1q1oh4vFV8qwlfiJbhwmujd01XJs+4aemTuj0On61Gt
6dshlv16BD5f3IeKHhABDe+qfLyEFc8gqvtNtUhJiQRMGuFeF7IPZn9yy3pvnjY3
U5iytf3WzVaU3qVcPiJqtdr8KWu3FwMkFXZ4Y2BS1RDyM0PGdjnjzeFiW87VyzTg
Ld7mKzaSoMnUfNrtcQPfDA==
`protect END_PROTECTED
