`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BuNMaWXAW0ZVNmxBqB9x0bg34gr3+hli17fUFUdiSCvoKPGGaifMS7c1nPbu0erx
JDEpswb+2iJs0qZDQTN/KYXuxTNt0N0XMVP1fEn09HedtnDCDjQ9mjY6mRw2cp/k
zo6iXYTal2WDsu4qtBBhlzIWAeFKqXrJXgftl/3toYoX/ZATNeHYyTXR4p1eOYvt
KjoeLfGhGINTW4/OwM3pzrjPWdRgXAuvVYioz+QobasfQIZsFq67Fku59c/eqRbu
fK060sQH10C4RsyToRoI31Hfb50Id9TfvB/OIGZbd2amYR4CWDgZdePBTyzp9P1L
Fz2WHx/PEU21E9LI6cE+sLxbpwcb4vi9OfQVZLQrEUTnIRDicG+xuDfRgDGS6pvr
riB5qg3PYuTkC9Fg694FoQI/8YT83TnZVDYDhbKV6PyfOdR8ErIBrIFwSaQlk0Ta
x5ZM+NM3nIP26xRp9IDp8nXLtv7gxnboORDKTnTZqLM7cjHi5GVFV2NnZZWlAtQc
tYtWNBAH5X1HuOrFKhUpWp7sgXVteAcptNIZdBKem9BLOkSEaEU2fcs4gP+oDwj2
SCSflr4j9nDoggPfmnmjdA==
`protect END_PROTECTED
