`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVznC5BAyAlgoLrsIn6gRufA9dzGoO7FMS4EtN4a7TnMggzyOyfKCKc4McExYWwf
BQlXy7facvF8K75paVbLaJVwrzKr5NEP18DjKgLIySOSP2wTJt8tJFiAALuTeNh3
/RzhOwjYYmrDZurIAmtZVYzZCd09ePH9UIRnY2FiiHZHx9kxp8vU+lCAtpXNl6K/
79kKONHNJLK1GeCxdAE4EEONfZrIMvR8GSaELinN6jVWV2MGEquEzMjgQlKvF6ur
sFV+/KZA/J745lrUjHM9t5l0CvnkaMM56Glt74l3c+m8L+r5D8STq2b64k/gbIPM
RTVNfGWT8kYtyyuZfaPIU0rZZREjU8rMiTEqTkXpUYDbbrNIpuIbB2aSoTE4anAc
AnK0yscqdswdz2P6st2k7Uvk8IfhhGW93wBR5bJ2osTqJpBgql4DKMde4NpKQfPH
imtCyYukToN/OQL2BuFUlOCxNekqs3dtt3HzVKnDvRf9LQTA48xKn1HDF3LoHnZQ
NswqfJCpng2fIgvk5+aLsfnIREQCuKYauWFaWMaTkgg/a+WHOXv/1tqZkAzArsqE
swxoalAgbnKMfZohDW4pLeYqKTzJePGT0I6r8kfsBa0=
`protect END_PROTECTED
