`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Xx9+hQdEF16u4YuMHa2qv5ROvLTsTtk7togFwNqHuoZWGeqnRC39zo/azdbceWu
AfrBYBl1NYF5sdER803K40HOGLcjaU6XqSz+BERxKbYVhpFab72qlD+97Mib+IVs
WS+Bgd9Kryx+EXV9+ORD59izJ6Ui3XGoL86+ONwFt/vLCUbo9fegHZSekkqL0NO2
X1GZe4bZoGsHAHim6f5jKfNmUQk9F5PS2BytwFbr0rtLV63w26z8dSoSUkffloYo
kb1B0HOyL4Ov0MAqiijxpv0JhEwatlKRM07JvgVQUemsfR767mwVqB0S5uicPwHJ
N4Aeb0rWON7UsE2/tvSj0sVYD768A3eu1MEePfVAUfYNAOHYiOXx28LM6oqYhRbh
uQsNiqOQsxDy/JnmzYR3qO6yk5lqesngDG27fc/f0wd2kApAOOFrf8y/M55BDzUv
949Fhl2h1gLJczcs2K2/7M1Yf1wgoxnb+ECaq1+y0U8s3HLbuSK4u/d5YMBj7gwa
Lx+ps7RelM7EO3TmzH0dk9RHaE4Kt9PTOwWSvbeWKRlPAUFQoA849j/1FfpntF36
HcUP+5+mpNdL/kwnkzcrVQ==
`protect END_PROTECTED
