`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdLvLPheiuRSA4V0nHH5oVcF6QwlGPpaMWENy1ox3jN91b2obA5yfB5F65L+1kMN
uJE1szWBJQHTgRsfrVmbnQGDKo6NKkT24FOF3lNHRrUl/xZJMoWOxsa1InVV7ho/
XjxDKago3kNS51ttYQQyabxjuRYTY0Qw375HXTj7mOigFRp4oBSBRio9E+EWDGR+
xYHD4IEUh7Cx3k/LflUKZ1DLlKSneFko0dD+4aCaeEhy+xUZN2GJ+Ex8yaq9cV14
000SnVxJG78NFxIUgqiDlJQqMPbnJ0S5ZSQJz7TeYlim15EjROjv4FHBuBdj37xL
YkUleWHfyTE5OjgzUXSHT/OkWYQw84cwcyrHR5qYkc9O9rx7POc0Vy4K6FptvDql
wt0D5eqM+wU4KJvvI2h6ZK8H43pU7XX1Sw9V02fJbgBV/jQT0ZSKc5pddHqdf+7O
6lrRNO2IcEpsDlLxNfoGSB4efUArKulwb+cfBw93QptL3aQjfZUHG/R1mIIX7C0M
2nuKySF0GLV8KU2c5S+s57McAbCmNHq6JeEfRc44AO68FH7/MhganfHS6dv3mHSu
lBwEbzqK0JVgeYWQIgqc+q9KTBbHy5L0UE9ZEinmvZt7sonxeMkOjOWj2WWg1Re/
yjFpteg5iyhU7uA+jsJ1zm9OkyJ0xKOk+4pSiJzbIa9y9EafO3o/pXzDd3cMTgZC
Wh/V22RDTkpnv55odQ21D/rX2O6fS94viQRjOnhQkOI=
`protect END_PROTECTED
