`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gfxlUHCwnGRkJM1fpz5LUtxKgxntjLlvthtaJjyppI1Qrxm+yQQvPo+345gX4pIB
P8AWvTFu5C0nq9/lB4S2a1ZV5AJBDm+qwzn/1E+Ye2LGaNqdDp/tPV4HF6P3ec+d
wBlq6hGUnD7kRCyL2XBac7G4koH7q23nQ04gUHqf4x6pq3Jg+QtIh81MJWO2+BAc
iRZqrLAl0d19oz9E/L1rdT6KNma3B7wBoQD09/9+EX+1iMUVue1K45zSWC49pV90
xFyShthHYbeJ5XAGKhyYvA==
`protect END_PROTECTED
