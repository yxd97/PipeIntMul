`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oVPwekjJmyd333smpkL9wMbNY79reTp3S354uPEoD7cPgiE1+BVAa0OXapiTzXEd
4tJEoJHcb/cKiY8RJNmmu5owgOMatrCsYXqoHSWySjb/hI6v8tb8CRh+8TFSiFTo
4NWITwanmDluNBFjVKrCIaP4J4TK+WmIwBp2iF1obAaSLJauyxLZxQZ2d/+68AQe
cH9MyYWA5RZU5uVAzpop7+mEk+5++Tm3RAYrug0DhOPFzkSIF9CuXpw1BlyDqNHC
3SxHLvq5kanUfsj/JLfvwvEhBc/LHjJY9JyAXsH9GexFW5Wre92u24kG0aMRYMzL
29/88c1giWb7NRi2UNoSs0yj2u1a96eGTO3J5YW1FOGS1e6jC0mmRa2Stt1WO4RX
22dVdIrpuZoE67AX/hJtsB3tu1rRbw6ZLm/IqbtNpdJVNMXbH1x7kZ8Ra3wAMMs7
IXvnulfAEf31ClL5OncYVlXsykz8yA7T6Eo0qX3F+KgBPUpzQlbpd0690OlwxfJP
ojhyfMGuROAvlBq3W130mootDj6a+IoN6gJrN/257cWpR5lQQWdIkd/bV4An8P/0
gsgNHrcrCyXUxmXL92FtMWVc5JCnxckuY4iQA6Iz+R0pp9N5hC5bWwi6m00g3pL4
JKupoxbwRqBVUpm98zxvP72CwpUuMmo191MjNWa6KSYb4T/yijqXDNUCiQvs8L0o
6dWil2L0AYw4PU7SU8xkvdemXNaEfAGDdGClxjblj5i4xTHHrBd0KsKU+NxeH2m7
HQwTA4x6MSsTWuRZH8cqMd7J/Eg03p7SAaYmkDFWc04ruOFBJS6z3MisjjMtUhd1
4Nqb+P6OZlHh7qiL0RM+c9L4urZmWNZilCohsRcqz20fIkKFnDsEJhunncReAsWv
l6iGhilUVg0hLH61b4n6DoOsuX6Jf/Xf7C1UzhybjChgGcupTIpuzTEsSXT6nhwS
`protect END_PROTECTED
