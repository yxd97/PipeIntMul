`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aA7XfNkeZgYfTNBTnjX16GmQMj2XFQiZF9GQVOJOiSMzz/rOJ0evI8ay3hx4Ywq9
omYF0hZEHXzgHPfoSM9x8vCFf5/G4sj5ITcaGJOXjL5CJiUkoBU+d4IBnlV0E3DF
b8nNj84ChD8K7kpmisUPfEodLJYneNjbF/TWycz6j0Zt4Mr35mrGwsLzOc6OeN+Z
wCPQFp5Z8OqiG+pSmNc/rHEE5yOKEvhGndCRIOPkAIzyWszpUjq/6Rkj36Ea0xsK
37hklKB8Hz03XGVAeA4XHY4yGQgPSIgbD+nDtmtwfTRqiUVTU81BZML13/jwkN0f
7qhpq1aaAGKfe2s+53as2PrpDE7f2mQ9xAxVn8w00lVa2QOklZ/pCa8ROWlohYGS
shAUcc57zFSF1YbZwCgphYWTX1gOEiWl+twJCV8yA9RH91jomT4MSH87TZjVRnHH
xCTPKlNIbfccQmrW9+ManeJziRLIw3aCE7a51ghmx681aHd5O8IVNQy9Xe5TY98s
gsntNcWn5ydvlfcW3tAXnXWV4iDLbylI75b9AE2GBMg2QR1gZqAkJjiwv66N3oTD
RnPICRCxqPUuCAmh4uVjzh70o/TulJLVPlk417B9lZSEEh61Paw1tF/syyb5pHwN
Y1XrL7uYVmC98BQ9yRTJBF+RBlASRKotG/vUJtEKOsjtEpGPhsjZAY18Kn98Jzi2
C/UbPitflvmONuCYxXDB5RRmTkI03mFENlT0bMKWP5hqRYXOfxvsBXwTq4L95HWc
KzpZ8Fjsj2xddKjLsz9tIvKiGRlI+pEjJC507bcacOP7tdQYlYdigFyp5y5lyVsq
lYlFaNP1Dtnjw/scLNijFzSU4ICng0ONnpC+qUAu9f7uH/YgMKkAxd+ia0+9HmsO
0PBoitqLvYw06G01RtN1JW9ljgRva30DXJsZNRqPIcn9PJ3/lQN2zHM0p1//waIX
t71xtQfl5Poymq33EO5ERVTTuckNAGIH2dtTucps4D4qsTjnW1AaDJF5S66SvcUM
lXOaolkw9sAZ/I1OMBwDJgZAxWjIKCqT+ZALOfNkocwivUieRKMeqgLcYeFl4tB6
/MjrbEXgtZTNknviY6HB4GdTDrJogWPD+nK9wR2i9pbG7OQKzDJ0rSm8scQs+8Rj
RfcHcT7m8ePj9W6RplMfMEyQQKUE8XaVjDOgg6P7xDuhzuxBC8FELfFmQSdG/j7T
HZ1GCbGtcqVJL8Bz92Qiee0ya2Sebn6P9o3zX/k7Ymvse3Jy2eF0uX9rzgq9WDSA
MQdoQ1cy2WAqBd7AG+lhih972Oo/k7+q7SAfOZFnIxiwUNGjWswZaHkVQX4RSozL
87s7jKLpoVR/phAPzQJGJgyZqfAPnuOd+YgKgt59DmOhfAz3S9J8rncTB43x2Civ
Go85P0fUn3O4GLvaqjOYmQ==
`protect END_PROTECTED
