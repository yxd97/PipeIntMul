`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJs98Dw6iEmvOQHZdAKCTSdKlX7ilRhkfuqLuBxqpu02hb06zOtCDcbTpMcmEvPW
ocCtZcFN+a5yyZz8o6axC0sJqYCdsmaM7SPNwtINMf/Rp53Qg6pZJkqz97/O8Iox
PB5leC+7J7IbnQcntLs1roEMQh05fVMAgqjHoVmxUlXcIwt5rvk/9MHahvRJgnYG
T8QPJwlvN9UdcQIbVh/N4BoKRafHh59iC5VZW/eMi1RHmRuTHXdXqEHg6JzDd+Ui
7xKVYfNaSlZ9m34stgD97n1eQN7Kw44L4oEJutgSbaDqsYQHAU3OG8yP1NjSdIlX
QJauQW0ujUuqziLS3q/+1LqsjfJeW4B0hj/C8SO7rXA=
`protect END_PROTECTED
