`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a86zEBDTD7BB8LlLKVP0clvO2Q5II5sO7GOuYArjkzfn3s0c0EWQzZOzkDWXikq4
GSgaCB9AIDBoCxrGe8OZM3IoSLExv/+Dt2JioFk5h+qruKAJ5kVJfQq+ZjPakVul
5aEXj7uZBvjFGTkrTHgiWyAMrtdpAEh2VYHHx3M582k+r4uW1TuRUqaiL5Z/vn9i
Txyi+vWatt97meKEmMoeAEk1iAVMf66zgJEomUs0aE/TJ+pI/DSR7/3AeaqIAOcM
+9oQ59jBE1HTly6dL49A2L2SMzFWNHXPL5xAAbKJf0/h/6VXpUjW/+qqTYGb568v
`protect END_PROTECTED
