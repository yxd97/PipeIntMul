`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rK2kVcKQiwQ9jtfkWeseQ3aALwo6prYm950Q3YD74LfzWruO3L5uhQpJ6EGjr+AT
68SvTGKrm2JOVTQ05VJc2gDJksNxgMfcWsizTw8+XT7l+CoKbG57mRgk95S/CpS4
Kn9kWwlxq0EiYDbwfeiVdKKIOI0PeDioTSpT/fyfFL5V4ehEKYieTJo2bVoCG19S
XxDrXp7bbRhM5nCblEHW4csib12wEDFY8JGfZyJua2nNEBHG5PlLLAH/8Ph0czpq
lIl1t/i05kJFc+fb8F5c6QHtlgYUOOGtLPSfW0xfdGbFNnJf4/NfN5fsD0E0usT5
ya95MHYV05+qu9FhxmUi1YsqvkEPXyJkNhXNQUhBI8w19BR/zRxOgyCJ1m4bjPBa
+lPISuRjINw4T1BcU4zToP26UUlOiZWVKqwXyixbEOw7JvRbgSXyt+oijsdioXks
L0ud/OVKnmwRCsQb6XyxTROdT1t52GwJU2Gq7ynHM2BywkbKhsBddkP46hdCBZ1z
vLaQdcBftX46wCvZDKypcHwfyMhDFrrE97GaqTvj0jOrofDgS/zwHAraMrApuNhc
7NlEmLnatfh9bA41HyDc8/h/uJT1OnOS2uGkNyYs0ns8jNOjMg9KHnH2Kz50z3qn
Cxjtv+YWK+QdmW8Ob/0kdVpy5Dod4H76p2bw99P/Dxc9BliFCWSHnVzFVnt4RKEM
oi0ctoYNllCOcHqVMEtn/8g3ot2aM7A0tQMJ22Sj91lnku7Ii/JSKuvXJuiy1rTN
DTe1qC17wChn5lPKQLuy2VxpNvQz2CyUlIBBlNMowHHvrYtI09RGnaELoNNE4FZU
NVbcGRa+S8Vb/b/BD1n6wbqiHKoUb3z1ded2S/CnoclMVSQ6ol7RTHm3+MdP1n/Q
6VQxJXUW6ZQpr4TB8QmTfwyO6EG+7Vuldu8EmEWiRaSXlTiNCztPGA/19E7Imlvb
99nikeWsY6eDWLJ0azSMWibgcjlf95y1pvnNVaOeojytCY3kEjHu+xz9ezkLo64C
T6s9l/dMgGUnB7ee0WAKB+6Hay6qXoW7hCcdvfmwVA1JBlA5pZJ5mFInXUXPGrEw
VFQfI5a6lCHZKo6+3cJm8dTBbHpVqfq7f3NfrpenfY43A1gSq7EaM0m+lTFz+NsA
8yThZHmyIlxGPXO/ojsUa1HF9u977LUbdkvWie6GH1pHTwORlAaXvJ+aCsCekvIO
5Ud/VxxV8kq63yUjgHsF5s6ZajkTHAQsp79GRpVXnPbEtbjcx+BHg6RsuhAPYqlV
86kMnkpDrIA48A3Zbrni9LP9MLDYcUBA6gQH6WkC+W8P1KmjNrnl4/mYH6QxeZuM
8OM5oQ6MQ6z6S53vMF9QgvDDjW5+NthUW66BmIKPYMxia+3IJS5Ft+gc5dI3MNr4
R1vZkz10e1Fu55r4oTcWWnIRS6U345FQKokpyojLYir18l3RtBB0XWIeznVDmNdw
lQcaIEN9EQ0jbz5xMWspb/drd9X+025nyQTMH5IpzTFxXn6XdUHsylcOsykXA51X
xIaEyeov+viAG2sYWdvujZFML4QTp6w3UGq3drY2NQbeRnT3PZgJ/mgGZVenOPPT
g7xtOoPgoDPcn3Vq0d7DsbxgWu3Vjm/0qENRPIbBUEWn/vFOaF8ON/kwCe4xcLi0
aixSMohP6Uq3v2ukMhLOpht8BVFJrX+Gmmj22mRe8iDbBxSnCf+6wkfzjiYnE0RL
K95NUQCbwk7EO2kl2WhkIg2xNZCPSAJin3PrpOKSoDzmHp+usyD2VX63Ue+AZF/D
y0TvZjqPWDS8nKD59vT6GATCz4xsXnr0Sgx3QNmbdP8v05KHTOsqMdC4iKrRn6Vd
B1aIzSZ2uEcIEZIuL5X2mZIKkJCT7AIQ6p7sy+H91t29NTSxx0hgLCtnW/MQ+u3V
tzNSZnzBlTWByRGZbOfJm7rW/a2XRe3Nh6EHmjcCGHUogIpX6KEaWT4WQZbFykG4
Y5txJzg6tPhAbs2AYxdZlz6gLlORQobLnFPJ2KEcvd89qwRfFaXwiqnsJ0qJ/nkF
t08xtSvFLsACAEq9BF2Um8BM36dQK54RPjUqdthwZuzs5UpgsfDD4FEDmXojMZHR
8cZ6Fp/Ob0ANdixzEq3CIX9pHRlx/tKBYCQMLQOtmtVzkhKOYzjgnWWzgxeMZYAE
8KDduNr9rQu7nkFp6psZlg==
`protect END_PROTECTED
