`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEuRtkXzgY38Te8Qu9OS4lARH0NP+fjBP8m5UKtwgwIJ97bW6RRaiRiqi9No8o91
LBjlUnYjza4LQNKPvL+IbQksLxrQiqY57kChWCfPVhkF7odW7NnOu6e/alTzWyWV
Um+UpnJL9K/OoMXDXo6+5pUyP6vytoPhjLjveXRx5/n/BQzWswrmnNlGhgSR46kv
Ve7P/7J6v+IUwn4xrVunRAPVqdQH+XjmvWzUqeKAepw3bth9hwU1WZTTGqZCbHcj
juATgLmIUR4RTu2t0T5L/O/bmACL3mfUipe7tFxnk9TFgrygCqskBZbOPi2S+3W8
WQoWlRHsLIAaNX9+znK1Roe86x1uYT8NosmQyi9XZtKWMWwisOQE3sEEN6rh1Qr7
5mYAGsniA3kUdXA+uxHQdjujpypoxTZWxNvgA8zcr0Q=
`protect END_PROTECTED
