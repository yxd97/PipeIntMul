`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luJw3XmjOH+38iZdqSNiH4YhnKrSwKiQMigtw38hOGUoSdNYvdePGVFKDAy3g7if
wj0CU1OG6fv8JDP0l9dxB2s8x2zIhdzTFj5VXMze8BiatIUsLrGxeZU26FKMoWgD
5b9r4r7t4yaSoRt5pPZvf/UE0Zzgt5VNN/iTUlYAMH+illBnDDFL42nQjbusGssE
zQ0OMK+gXlhROGnDVWO0EhZitDriCDeTwMb6WUBEBNlkvAz3dwJMGXKWgRVyXqQD
FMNzIYYvgvw7uDd6KfQu4mDp07RVsZILiLgXFhYxf/yc9e4tripq84TIWtFznPo6
u+dZDbrE6eevQx7wEnigfg==
`protect END_PROTECTED
