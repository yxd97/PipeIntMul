`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CFz6wkUX1ggPxIqTReCb60rNH3Z9u3B5HAv1pP6pOjKhiIFFnqXhJG8dNKJYMNrp
pW4EYHX54ptZcdCzuveBmFnFbi1aJY1LywZiY7cp988J0kfw/0g4iirxrzRQSDqA
Sun6UBvlJMfhTaSIRW3gvlNy3hO4Tj3Q+Sk4xlj6JXs7PPASeoszvev9V675ERBV
W1GHoSPkSo6QtDfKJI5iE9nHXtHmt2uM0H25kg0AnKIo+GAKdfs6FlzunMvNB5wm
0GTH4mllD/Ls1XTKYwCuDLCo4GMvM72LeiZvIiBFj56XQN1htakDBPlghY0DDvPu
Tm3DJprJgt3Ni28fYknDbVkLAN6lWqUmU30pgiuQRXj43U6Yfe7ktR8QgFLJ5kGJ
8g3+pkjkgoHC/jHinALmJ4/kfV/Z5i/jvZULrqyKex0OyzFcfopTqPxeSwiEn1nN
QZih35FRnTkm47F4pzE0Trs60/qbBP89/o9Z/yHeUl045A99hE2L8lle6a6IaycD
mJUG65R+nUAgtuR+OUMmA0cT1GxOMCsa6wBhjmDZSGMLNH4zqRncAP0IdUuMjFm6
dg7/H+C03Q9TqxMDJnDiNzdORP0nqmvpW7KtU+dgL9WO5CHNwb9c5y4pxmHJvbzn
mWT8wgNmkrKHDkVE6P5V8VC9Rh6zRJIe5ntwBFtd2//55+9f2npxFR2N0p+EGVUU
vcY1cEKy1UpxeHckw7N01VH/PFGBNaBz12zf9WNeXb/yaOMWeVc1EPAGbr5GuGNI
wxTFq2u0w7mNlv+PGw2rI5LaqEiKlXN5fGQqRC8pFHA6p2hofWGQIVo6YMYpSrwz
mXe3v6b2BV9FyLYBAImoK3TOxuyEftfnJr/LxdzxNpU3K2259QWpbXChj4TuSjmq
9nFHbiyfNkEb+uKZJficd+DYk/FJ8vIJP/03AfcizzXjIe0kYreman7BNKTj2u9m
38TUyN8fuyekLcGoxBjecL5M/F9JKhsM7i7wwaQSoZw5JvaL+KUBBr+WPQwWnWdR
6NaZBy8pNsUNH3KSNW2+6k/lmhaMGtLesu+rmTJ7EHZFjuXKjNz5Vq3II26sPgFS
ERrislZXZBCPLlkn+G5W+vocI7YyvghogXRlKvTF/kVgkG66d0S5sbD6ySxqRNnu
RWYrfs13IVhaqbvlk1o1QpR0DjE3AM9qVARTZmV53F/t9WcSE+B71AQB+vy9mJFM
IWTkKy/ZQ0d4XAkeFxRWjrVcTje+JnUpfNZlB6khABNiCRcyyKktq/P0CjFxWX45
wUDyktTUaYdcvu7SER7tZMqtWd7pGQy9EUV3mvt462aSMowSw0XumVPoVZG4lyCP
HKqgcSYQrfFwLIKhcaelMh3pLZOM58tiYGEvcJTueKd9v9py83S2s+z1oP0iT5ew
0EwITrriv8XZo/BRjGjuFy2LYb4CdTKl/X7YJsWJb6tPZhbrx9GmwpqK8oUdIniI
xhaz3HxqZeCIBLU5xnWuBBkfbWWvU+GtYtGAx2a+gQbskGePAHac2/p8CEzA+SoD
rTVGN/E9DF59h4QU/jJYBwaKolkJABSRDzg/h9dJD7JpzEY2uAR3jUIWi9x6OqeH
15bF1FU3whvh97mVjIK7NF6EBwyoC1dcxb4ZM2HkiJtUcs65DeiHy42F/kZsar5X
sQMR4ees4CBR8n6khvzLtZ1qYb7MIg/sTQuHUPsmXTGorf9ifc5tJkalRkORidus
F7e4aaTON5ZMSlYfTqeALABd31EO9fNYNrZd1ALCG9oH/1tk1MJS2sFjQI23wHNP
XZgBJVyugGtf0+F0PluGd62WrkHqhnzXXjCmu57GBNRA1u1r5+yvScN8UJeLrO71
mvNANrs0GuV/7DaLyoW4KNlndzqTXUQzcVLlqJ96T1dWLLYQI/vKcNtT4CbM2jOJ
SgVtRTgeSegocEASNVW2zO3mUSyJBZFe/9qT3fUuCw+g6mACplVs6eeUQaHjlEol
3j7qNDz/kn/rcR4MBbMWvyuBDE2HY1yHVriPOENCncKxpUr/u6WEGFdZvksUgSZ1
d7D+X3tTS+YIytgcCeyzPk+s2946hqW5mUl6Z4wDoYls9mMoyKILBy/tmMM1u2KN
mGVqgAcJRlKg6wlObAXlo1yoAKYPI+PR673n4lQTqvsIsLypQC/OkGeJXN0WE+BS
d7puUI3nPal4RpXjhAf+2v1USpTbUuVLRZzpg94k+bbKe7mUd+c7ZK30AnpbyNUi
2MejsiBdgA31hZ5F+pFwo/AILwyK2Bb3Cbk1TeEV+vY+iaAZHIA41ZVgh6k4uql2
KJUBLzE3UaK1C7nytMv37y5XjedWEiUM/vwRFhGsuX/0A+hGv5WopN0o/dRvUMX8
FjvdeJ8bPEpEMLVIqLCS71LIXfEQ0O/2x7FwhC9Og3MfAA0zQ5AGAyRpvFtT+6LP
7cc+rI8Jsh9CVxUaSBr1xSJ6hoyvO7PD1M+1zklRLqEtfiLQQSkLSk7fjJ4K4hZq
1ca32MF0tMdQVRkVYi3Fq8GbLr1Pqupm5vE2MQAFwWP5/vQGSA8hOi8XdNU4ajNU
R/A06LbkTeCVK1bUXrSKD4hwIEmBF7FIqs1GxlL9bKwTvLQGPC8yWtQ7zMEJ4WZ0
7K1JdYgAkBgwtYvtODOmZyaGZ876zeH+uqjNfbNuxASQs1Y538kzXEF4wrDLy+FR
RuV2fOtYwr4h1ZaLvQrpW2bO4iNSV9aN69i3Rxy9XHzBPgQhZG7Ov6eHlrX80vZQ
29ONVERkWxSv7E65E9k83g==
`protect END_PROTECTED
