`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tEhSs+JShN7YjB5pyHbgtpvk7LnBYz/PAh5muEbLLZJGmAO4kO3yJOYulSq022l
irwuHJZ0VYnnGx0Gqa90OBWCNcXYRmRnL/OGtiaMrcfhC6KprR0pp/jMUej4jAto
h8dGQs8pgsDPk1nckddzDaE6jb/e0I+eDGUAZTU/m5KwJUCqnKqO6GMYVXt1go8c
MOOYBhFBa5oqUjyOK7z/+c3WB++24Gdf7fkRAplrEL99LfvnGBKzucWiy2sKHS7M
V065YKk/MQFE7oqV2c7BUJRCrl8/2QjYtCwPSPqFunEq8HDu+6QdJRFTnpfvmWz5
h/RYAataoMLYosB43HUj2kJNOqXkBWlZSCT+meyMoZTq9aWI33o/3txyf2jO8pe9
o/HXf4pXs+OPdmmg+p3dUUZF1JLxVGfwOECKDMlFIi+27FQD4202fOmlqdtNfJFo
WtqpIj4sNVeczy/Ow9QrjdEvKhrqORYaR006slTrTGztuLN1m2x4OUdwZozhh8B+
CFbB1zyKy+Nv3CdKOoiJYGY1GRatDFOM1c+IdgT8wy2zxUHy/jDXhDDaUE4sl3Be
8L5HP+V/+OV5KsgjdrGlYQ==
`protect END_PROTECTED
