`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1icSowB643CodmoiUIHLxLr+7bgpOSJtHi8SSl0jKay14CrdEhMHGFfwjTarWuW
gwtXQ6LseZybgiAZFRCShYcHQ0cHSWYwr5bL3MnECygH6pjzHrhwaZJNvfWHYxzL
vAwhea9pw6K7SlzPekTBWTHhZyAwP+zqGqPY4Dew889+LzfYUaYXlSjc+umCWRD5
wg1tT9G0P2kJcm6uotHDL9ztbwiEC/ub5qF08iu7GiIUyDhuKJv0mmQZ3GENqz/i
HqDFwI9ooKx/O23DzCPUHv4uf4hoKAEWydtb28LRTrJcMqIT5gN9b4KsFwnyJ2ly
TOsUy8YWabyEdgJPusS8O21J2qcza0/70DHcSbymsJ2KowIHyVGFDdAneRAoQC95
q0KBpZcMpv1OBtXvWQiBQt5P2qhoO8YeZ06X4H4PlJdUVHue4pw6rxsRhBKhMQqh
syKg/KNM8JSuLU50S4+4QQIrPy6VTXvGFegG+m3ytLCRucAJ9ZlpOwuKMKQgfgNd
wNc6YRA3gtUCCMTquZvguZn83I+ygFmIuMFcLg8ROfA6DD1zhahnPtfI7vT+Nico
nHPP8KRB3+xAsyLGV/b6dvlNxG2V3Bnt9BKT+Yxw9dsKpoovLs4szCPRlCcB1Lpe
Mdqtr78+O7HWnP3rvUO9Kh3VcloN1W7+F6hjWHN8mz1BVy55Ql0gmniuGNrOoTS0
73jD9iGZC0pqrIReVrNBWaHWsUSlT/vvI55/cM7EF4f+qFba/VPhawkxHBNe4BGG
CoC1FIgKHKBWsqTjKXhYrSWTRvR7DNGFwf85Xp5Mumy25jgSylhDWYZU9569fNv1
xhomwoXtm4PYP34mJAU+qbTDDZqZXmtwMj1e7JXFvCRKUqxLTku3MuW/SqWiLr4u
IHVUPiwStIPAEO4FKC+lhpAjy8aHDWeE/yIOrYlkv44DNC5vrrSUfDLtDzWeNpGz
8oY120VVCtie4ZyH9vVlkpRz31zQG8nbdLPk0cr3ChBciDZffEJ7+XevnX0wIY0m
dG8+mNLS6KBHzomZObIchBblwdV2KagJbZrZuAacgc0vyEEW2TAUTSdyaLurTrOO
1KyBiB0E/QnsaXtM60f037xEazEw7KIAfhzGyKhPr6rsapA+90xD3Puw0gMHPeab
EjTfvW5o+tZj0qRp9HGjtZEDfq0yh7bZVI7gHJj6jxzwmzc8EXjptWXXrAXcDcGD
VlieiRl5c8QEsGI4Hm6IETLEva/K8UZvgs1lmuhJInHGnJ5fWJvTwMQ6aeE4KDNn
wEB61z8EP4cchXYz8Q4EmwsfN6rOKmiL0mnMD81pK6fWjDVLdVdZRoZb/ViA4K5I
+0vCZE5cTbAlNpk0/MZWbRJREHLYFv6Nb4ryY+TumRVB8sqKLxXoLJqFCV0n90Fl
wdPh+C0v9NpHyVijbIZK4nq9XGZaA+2FT+GbBXdW4egcaTOc9RcV1qQQ6N3l1Fdz
d0F/lS8SGfo04eAa3fXs+KeovyllYlRwf+L6VZw5tHxztHJQcG6za9MvY8C+5ShN
SdI5sWQUR89842RcN4WvJEMhlFDUuK7H4VAPMm+arX8AhbACQjB8Qg1FQC0Ltbf0
8hohWibmfKSUX10RPQLrx3ZX90H0uItjwB/NQDH8egrAYVxrwQunIRFgjwihQDHF
tBDEBsRga8wFH/01qiJNnWuO4F5/u4ZnohXk085GVB89JV31uj6UwI0PBASLxlgj
U6tYZYcfFYavc5VQhAR4nZeQPVECn9R0G56Rbepm/FavNSIoQcIxOVzNKTZe7qLq
l1/JY64+JLz+ZddefGrKrd695CL5TS/eSKagCFwXOgjySmVbR7MwPXRJCldJDb1X
HjPhBiBaGUCfMaJW/Ta9AVn0xA6AB62ZxaFWkx+eEJ5508r/8nx4xuyRQopaahNM
RG72RZmfqjNM9zwb2juUeUcnOZR1EcD9PhB4BXydEheX1Sy3myDXNnHD731JxlGk
wqt30WmCOXK+ppZLyLNNgOHjeROzLHnbvhz6jTxfdzZJ3Q0XDdE26YPOxStWqzYC
6KNo66v5iLkKmlTGBYbh+CACnoY7UYmGtB83QBpD5ieHRGUv9FA4bHwxlGownBrb
YQ+Wt8388geUyyLPMWLOlCjhp1xyRZMCQ3LdboZma35GYEM4iDem2IKtBgPaZA3G
JBZ4MQaEKQ9KBdbjjOSdAnOCZait8xHYGrTZlqpo9TVSOdISWTVmyLoI6gyqay/n
duC7LAHcTjrSAxUBxwflfmYOWN3j/n8EpDbZqa/cTk8M4n871VvhyEVbmvqXkqJ0
Nee3HcZJj+v7uXVYVSkZNHFMq+30kiwvqmCQS81V8T+tSGWqczbn5yAo8hr7hZjf
HgNuYA3TyR1OcVYIiguiT6dImbhrNfSk/WwEn2y6y+L7EIZ3tvxKuXuAKnGvfRqV
/v2tJvNaBxF3BnO5WylB9+hctei1jEFLD9kHFKXDgEaJr/QACbdCqtaBb3UkGWyP
lm2yR+A1PDH8ecRtQ/pvaOwa1ebRpgS4FO8s0yk3D1qeOw6b8VBGwWpd7skpFIxL
hSv0hzl3je0h5cbxXb1c6pf9wyzCWh4SxuuwtKvhus3cwH6rrTjv35PUcHRqCMiG
XuLOgmvtrURQAnraT3qmyy7ONuYgfjDRE4tfmaTf7uTEBN3VE5Q0JvsCThyFxtYy
r8fdWHv0/LG7AZodL2ewJ27142K8ci7r4i/Ni/IlWVMxqdViw01MBCwMMSrV+qJ/
ZQrbWDuKKS7NhckeKl1YCZDJR11ZkVSy3znbKgCn73yofDhaXvivZfV2jsmt/4kv
Z4ol6iA5iPBCYZRsxua6LHknzFcFr9lMD3YaXPRKCXvwU1T85KeiCLGnB64PRU0N
nz02jNMGzNTu/Go+gu3b4UJESx4pm6za9Se01rnltVprDLfmhjSVNW1zUxi365E7
/5xwt5A3JdZuYqzm16+1RcBPZaqn2zcnJrTAKkaKNh39Buxf6/hPzKRJnUAIhEwr
VIgbyfzx2QyHKZM/pnjP8B2e1AiV3tyvGpjPuOuOVIrptxUtptLZa4pxuouF2CTh
gsOEbnRGnotAY4PmW5+lR/lgh8br3fQoWWGLUCyuSQvSV/R10zMT/nGNYe6kZ3Rw
nDynznqdCLeKp2FO20Hg3MdOEpwJP3nI87jbGWAISbZRmr+E2VvA/ebQqc2jkEyz
Lit8A2lQc/qbWSOE2t0EdrgykoupjSmO731p6t6ItMdKSYIA2Oo9mNKXGf8vrPzO
nuASSvRggxkgqOIiROnu7uzDxGGkdfRkReblPMpH7pFk8bzWRj1tyhjtG/3H+jke
03jAz5dYJzeqy1DO2cRA4GvqCprem2fcpMB6UlERyk2Z7TVTktXEAUT1V4qQJ9ie
GVw3/hl+mxbJ/E4pPcEQREbUsDcpAadxkPhi6YPtTCwUKCbXAJcKQiMSo5RlDbrG
b1AcejItnZ4aUjN3yOSs2oWgGRo/aIBZfziNNKK6dPE52ZseaY0WgMh5RFxuT4vB
AMFY1m5g1D9JPgV1TS/Fr6y48B72HZe6JxcauQCi8qpI+ylxjn3DFgePnjQ6GTPQ
Jy0YKNOrqFccAL0f2UYedhDDT72df/7uAVx/ly0Pc5w87nbS9cPVFYKMMRQCvLQz
m/lTpPXsBDic+98szAnNcj+AM3B/tIXL4zlcyDxa2WTRB7aaVNmNApDPlM0RBHUU
TzvG1ZAw/uflqHT7R7s4w36UUVxN2jjLplNzAHtvUX1F7eTcvIgc34vVIcvYj22M
DRg5oLzolGQmwi9ohGdgBRUwBatAsXSaVTI2waV3/zKhh6c6HxwdpNjL1hSRsu4G
rXBt4uw5VIwAY3LiWAcAoRUHD2ehu4FWy5QvtKB/8FCxIbrTCWdcRClNFjf0pPCM
VBQASdaflrXj0lZRUmrT93Uv67nW/mL1VL6n7YLB+AwX+bB5kscchhsnIkResIEC
UZ7YFfhvJAqLH9DIzxvLcm4q0XAvc7f5g8IA3fc/+rdzX+qZZ/d/EpAz9F7iwtAD
PMvji9znOep7xDzMCJw/p4Vt3Gno74Tow40jUlTf8cZ7/iRZd4wZHJaFhLJwwpIo
ZYrSIEF85OCEfgcO6041Rp48/oESH2bwzH4fMDF10hU5rR6YEw7yH4inMmxHGhcF
QEH29wwyiqEvglOeJbFY/6FkgjwiK0Drtxopd4vV6f3ERCr8pyIc1Ii3KX9fpUON
DeLijop5hX9taRigBbR4XKr+4W0l9JKse4U/siK9g/JNJSbzcdnt90ZYgsLSUAIN
Mc2AFDtQEwp13CblPQ/p32l3TkpIvoizjfYeDeXFwcwtRmM0NGi2ksHB3FJO4ahi
RbrEF1UfIKH/k3NLXEGpubw2ZOFQE/uABPewXMNge+N5/Q5f+L1e/MiGL+RvmF76
ZP+thjH99e4/iuCSMh3WncdC2gorf0wGLfuClNVaM5/zN8vy5J7x7aEfyUe16t3o
XUXXMqLMl86SYolbkQPDll6sNUMon3ea5I6558s2oJRhxRoembz5bHqX+PTYsiDp
jo04t5bkfu/sXRfKJBTTKK5LoUk7ONbT8iXhYEDbPlBvU2s1L0mQ3HJpMRApJBKk
tPl4rSOHPe3ZSIfRu1Bm9CFsLFt3r+FpHWZGvR/dg5QdjJC5VmYR8f2QOZAMB/Fc
AicZiD26XYPvvIYRrDYmI/jJAwCfEi8zeMfeVb7UHULkCEgXTBFLooHWbbC7cACH
XFS1DynCLREtgVsZGEnA8rUH8sHShtFAeCGxzncdW/AccbxMqyw1iQoFPGUBcUPi
2o29sRza97lMm0fRS1ainhv0ITxl6JGnCBG6X7nmjmc3CTjO9GlBi4XlYyzfdBTZ
Ch1okHOqIB3F1mIhzYG+J0BpwIrqBSG7mVHGqDpDbDpxPDN8te9zXns2gdh+RHQJ
Xb5OrmfNHElZXIZ3JSUM22qnltkb/RS1HWIaSy09FhlfXswK5IAAchRWOf3mRD6N
wXaTAYBQ3rfqq1mmYqVySYBXjfj7yRTkKxocevr6NT4a/VTW40hewJvAIW6+ju75
7QEizdJNHwpG5ItMMF5HjHCpASKQa2ICYiQ/E/vCUSSmpeCTu9C91mlSjurSvwnK
ZCT8Ig0dbCOWlaLdkd+ZkJtg7S3jI509dJNeZpKB+OC/Na3mu/fqT04+aQ8sVrAJ
l8lZaNktBOU0fvOuhz97garBXFgefh1E2UPS46bQSbKiE8+x525g0CH25Eo2VCgJ
FMl7dVXKCpoJAj+8HG3sJCzZxxt/xUBSKfws+zXB1DL3I9/uMPcC2/E+tq1Y/5aG
M4N8gboV2iOvKBIEdZAjo1/aM4m1m8FgLwtpBGrSnusble51kPeg0daYidSa2137
EqGnIY8HBXDNVT5FygWapf9dvxssweEk89xFQVHrSQgZLZkSVAOe0mm/bFZOcWTM
r4K62KCfQqmi+YHepw+a9A2whoThEYk9lYt3cg5bbcumxUvp/FuOPsaNO0opgl7c
Vf2YGA2iV+MIFqj6l8TXOf92gGniTTrdHev0kUROkQyT/ESc8fmW3n3t65qwX7B8
rQGyXv8DCZaeS81mfSTHzESu4ub0k3d4FS3Sn2cq2zvauBgq86mQyluv22apWbdq
fDdOywsP/IdVVpq/nHjCDA7lJHwNimw55Zl1/6lf/Cmw0ieGbrBZT6ExvSe5+oBR
JbD5i5BwN1loXrwpU9sPHt98uD5fKPQc+WZA2y8lPfw9fM/IY1sAeEX6xvSlobWC
Cbf832sxzZ3gH6JUUXa7acR6TPV/Y80utsHNbVxwgGHJ8KIbZa9BzIEp+EyGWqjP
0bX/nTFIIB4idtogjTdvX7iHcZ3+TsdmjrvfRyNeRyjv1lxik9rpsfIFw0/Hbkp/
y9NiRwiaxvVyaC2BD+5y8K5fUgAto1dlsA00wjLg/UwdWjoJ8UtiANVZ5fYyj/jC
X1X8FfMploy418E3n3Ifc0SQKwh514b6KtUvgE1OtFWQGmT5tPAAVNewSG7uahJJ
L8HThJ3J/0H3uqy5Lp/P4/TP7ii420geqwPR24nr3xhMe5OGIjXrHmbAUhkDjaws
CyiFbqBMfVrAv1VFofZyEcDHGv/nv1abnohvH38T3NqCjyFM/mgrX899TcXI3IeJ
eqc60CdZUqMHcepJFG1WcaIHaDxyyUzFWdVX4bpVRlQrCn0zXIkUq6Wt65mpG0dd
0qHBC2BkNOWMffv+TrtjFjaXD3nK6jmYY2/5P6GfUhoV6oN+wbqvbdFdURcjM8an
334I43X7jTxchCp78tJ6dLE3nbrg9aFKhxrTUSe758o3+4An0lDErJm4x/MCkPXM
WpywgMpmkuPn/2cKzaphNuCynEjS7cCLsTXCa/Jb/d+kpGRXJsWT0KrqjT5Lxf8/
4WcwIQrbG/9GCEsrAWFQlG+HmWFVmsRYmKDz4Qne2CqhOMDCoINrMgI1gQqGxiap
bEH4MDWkHv3O6DpD3GQcmaOi4N387eUlOt0pis5Tw7j2KqBiOFuhA5vIMCAAfb+E
37clKo9faDaLcUmhHnrC6Lt8/FiqVvfGKuDoYXfY25Pm32PIOx15eA7FVwi12lxx
di87mLteFDyO8AsQQm9AmlBK0WIgNTBeLqh4MVshIMRnYTaaH0ZySBPojULQxu+6
1Iy8IMBz7hBK7Xwoyf/Q185efNJBnNeIqU0QUJA0KrxQLZh3y9yVmghnvFdTKOab
unzXjFpjz+/G5xFIqf9niTLkVO/8E853N+zbVwpaN26s5eoBMHferB+2LZQjxnr8
ZN3QCslQeCLTOt/bgz5XCWcQbGXmyCS2ZeOB3ATWTS6qSeYjFM95fVg8gXKKgyVp
WocwysNDErOjQaOgU9YvmJEptO3xkqxMuRSEeIHFHxHSsHR8LPxsaJIKV/D3NjyP
GZytVqTsy1xIUiYYnpKsv2XMIDyTikKtgQjbuD3xvROMMIxDcJY9kixRb7D0zzoO
wMJkvlWq7ZhfkxlTqw3uxnuxosh+y1Zg1PPs3ZuFEFTU7nLHzxn2SO6p+iR/pDQT
uTXNhvxmZL3CoyOJhINXXV2d/jfezhim2QrRexEylSMMW9YgP56VgUVn1MYn5sVp
P1N0F+w16JECWlPCzi8pcUjU0jpEe7sFsk6Q09Qyzedh4m/YapyN1IUBGQBRldqk
WUTNfNyU7atIwbk6vGfBOua8VtG2X/AGXwsfgiJ1MoxbCFLwnmOzy807Jpr4VLAH
i3yuqO0IEIs4XVfctBKh/AVvlF6jkB1uNi/ELYAD8bUfvIhp3VVZ92Kytc3I6Sv6
oy05RxfLNNdagmuy+XJfLpjVIm0716GXfSaPtMkeUb+WktQq+TnHdFbuVM5omVkb
5KArbrOAUZQf2l0utnC3Bl4n1FKkHknWUEFoxiQL8LHL8ekyVUIpZndLUzyiD/2C
nZ3ENkOzt8SCs4VTCb88BHLEnPaydl3FN7RhVNhJLRWfW/BSQ51nFf7G7pEGJAln
X4RbLQi6CHotjTeG6PMGFlaLxtefLiAluJcTABdiXjYOsMlqKbPfHExdeVc3vDi+
B9786lRknG7in04GdShiZDe++ZTi2c4qAg9YsBYhUGWDl5NxMRnSSZrwiSx22cjn
9FK0Ew77SwEj2rckupTAcVfyJGcqN0svtEC+KOae1/UbXcn7ypwm0Q6TODz+PNDW
ou2LgDiKXDOLBzS7mgpCbAB1a8sAA4UvzQiAub8gCGoQNPwMRkgdRZqSVAf39Jqo
ZdC1jqqlTD+A8hV07ce07yvNTicN73vRgce1803Vfg37pjnTiWl2qt+H8d6Woo21
zwtlveqWa/H2O9UQHgrGuX1AT/tyZp/Pe+NZNuwieefW5kB1nWjT6cRiT+2dOyIr
pQ7HL83hB/4Y5qruK4UmUUeMVP0CGKt3Lgr8jBYdYnu/2Fk9VEPyMd9f2G0MOAhX
HbOXbqCk7Bxm4hm6EMNDTQ92h0CMbXOm8j5EJnpapKSSPAUA4kibvwI08OCUo61h
ebBqCKhT4Chqs/DzgCOSWhSmnXLZuI95mybiNjlreh+YZtzMy2DySJZYmpU9qe2W
nci0XHy7p/xFkscbJZhMjaWo1I3ItbyETv/T6iZau6Me4TJ2XOyrVo1ZbzmL4nr1
wyNcEwYdpVKE9d5vrZOSULQfwtJrVahlFMq/rmD9QnbF8xcEXYK44AWNIX8N5tV/
VzkkkcNMZ6ktKeKEHw5rlusU8osLq6J0xBaAv4kxXX9SF19jGCVPGcSh1ZBKav5i
mEoyLxeYyAh72boapn3fy4o1FQTk8QvUN+y7GsNsvmoB8SP+Ao9xebolaG7TMCON
QuHKAYmxjWIs7K2iNOYHtjcmVjf3AnpP5sIN07ti3IqU2W1qonIMAQsudiuzcl9g
83QUwnKmyw+buHgwl3pBAajoE7eiq5hwcqWD63tj+uhpdlcbPx3vN+FXHpqjB9EM
4Ul5bVuipS0Ld5tcx7SJ3p8b9nBBOkDNro4ty2hMSjbWYEDKjWJ+MDcri+jL2zay
gHrrHKF0XLmJ4FvZ80/U4yYeSbEg9KEU2195PFpEUBGDdFEZZsiIswJy04N3Bcmh
ump/H1MzpF/pyvU8Zjs1+0s7NJdiri+tN1t4+CZbJnF+t9BbBwNBca8nnLr2RY9X
g5Xqar9TNRp5FOhu24JfzxoHiZA2Jg46XD6PQjYKgiy8koUeqqvJNeDuNb3zOx2B
ocAv/RzFvlmT1J1OLc6kKMG7m7ON0lEAhH7MuSGgBdxm2aFk8RVBsbxQIS1bED0X
dvM6BdbREEcLvq2Ugzv46hXxwtMZtYg/RmO9D6KR5BZBU9WPpFaBVGVnf3Q6RTd5
vHpg/XAmsa1e8VXF+mVuzx3rf1T9o3jrbki5/h5aMkMiWh3OHaM0frKiCKZ3qtL+
3kdwrVRnhmAtoPcRO+LF4FVaAwYaSDyx+cL5cb/dznH1VsywJ4n+lf6hKOu8oW1q
GqhSdRS4J4KS5pt0VU3gv6klIMltjbHquPqPb9BW7htrR85sM0AkWNCsoMQWjIj8
B22vYGQpbPJzB+Hpki2x5jljdwDd4zp3An7eBD8gQq+wOpqdpAkJy+tov6AwkFd4
L3Hb1b7E23Yaru1ph0spcneqZkaPszHS8qhknPf6JapsCWEMtGoWEbbM5J7MmVPG
PsKWh+xUs52EEPLnRKux8jPE6Vczvl99rGuDEZckETFyww3VPKFWB5OLNrcDnX6g
27bBKG36KZl2kBT7LV5m/jDhTYeBzQRffUA4S4UWjtP3lA8HA+r+p7gF/nmlr/pA
liqk9uM/KgMHDbUP+4kQ7KtDjitTOK2Z04GRyn/vfCqdoAfRtzidOrUIbqInICaa
WqMin7lXxZlPIXRmXjMCrNv5rtEVEiY0PY8vIkR3vBVxKaIAREHaJewKQ6UZYces
31R5C4snkAI/DY920/JUm6/4asIQPvpOnkb2XnYBzgL/JwV6S/+GHRkWks6qqq7V
Xc3oUdQN2LBJ5lejHxt0YhZSoFB6HvzS9k2AeoEAszl9jDbxdcAEZQBqmCic8iYI
c3/6AD7i5tLSun9pglU7K73niQG3hFFlItTGkZRqw3QFwVTpthd8p3S+dZLjI1mf
HkeWzSlRSPuGEMyTugwofvM8P0/I/0HVHL6Enhk4FAEogBo4umdy/US8k/C3nQgn
q/MpdmvvRiMdZzPx8oR1x4KWVCI8EIFjc6RO5kQMwDm8ksbmDCrCCPW7i5mfrKS1
UbaHqMX4qz6BXNYp5spHOnjnBqEqBLfWp0mg9xFgpuMR+z8BwY/J1rZydjeyUWeo
cEV9LifJhUysUdFjZCl9l7iRg5Of1Ww1s8eseZ5/7Wp5gL5/vpUiHOG04aWicWME
7xJz/ZcBa2RE+B446MdhMIZop54KPksVK/pe9E8bF9fCUQ1DFsqkjhHxAmxs4nBK
NPKS2J68MwEMWlNmE4QLu67lsbed79paPvwdqMfJ59lAmwobGL724TC61mGkwEEN
OpztpvM2AWZ8vmD1agma112y6RusN2SHNRFFclD4kKYZTM5RN60YijxFcMX+tPGC
D2CdqNUNsxTz6pXOxvF3YjVVbYnh1a7OhODrQPjW83jfBjAIc22WXCO9ssrfMNMT
FiXHDq9VmkOrEsMEZ12DB1+bhVN+SSQn5QOOTSK63KGc5b0+LrPJLQk+dVw5AZwy
fQg6WABa/OYOrne0k9igSFoTh+Kg+v/1K/X2NtNvIj2ZolRI5TcY+VMDopvAkIqo
Y5SIeFmIfe+gNFpmS44hVFUbOk7MwAAzJnDd41ffVyN116KBmvQ8aJUNGBkKhY46
NAr2hcQ91N1h221acPn5NHAO4rYLdU6p02dn0rlxmI4mrXjRRDMp/xcxP0KiO8H8
AQqAuH6qL4U+J+HdihaXa28w5h8IhnPNVA8CV6q8o5M54axbflkPXWULx9yChil0
OgRnEl6oKrQKvFYzBkqCwGlSIikToIXbisdrXcCvszPzD0scBHG2yMM6RZA8mNdb
MeOaH2ahD1Q4ME9koT16xFx6Sv1WJci2WMo0dhNt+PEDRQNOsc0HlE1+Svpt/7H0
u3cwnlRpwzxgeD3K0tlQDYGzq3BRG5PhI+JGIflef5gaGdLQCKjYNirmSw3rSnJw
8aGhm/5Vskf89/CXSZQIABlNlHicPaRXuYHvrO328MTegoD3rRSX4gbH2aeCTaAy
Te1gDRZktQZbrzAVagGd0RpouGvGdrzwhiOHpADHgsCMa2v4gwhO8rceHwlT6k7Z
BzEShuzYs/8GDq/f3l3PuwcO1Xm3Q4Je8haXzX3vND+een+Az3141SqkgPi9iqks
99Yxc33EbnWofAcFWGnlNWd++GkjyoYQvFZUoatTrQC6r95DFd4bEXfbai+y+yd3
/3FUBXfIXFTPl8TBS4Eb14gjaj4ZC5/VK3C5+t/pIJ18JB0tW5IQSvccGWRqXjoo
eWwdUfOzKgbNV1IRlZSe76etHof2kjsOmb6vamtww8Z9il6oRRn1MIHxOQ+Vk0Pd
qRTj3EucIM3LcTAF6nq9XFNJ6r1+OXXGHdYJFWAUzY0GBv7C+JXA7ZrIe+95++In
FY0Lp9fKJkOaCYAoBeuq8U2yhCagl9LlFbtyPrtciLYEsQoLGyux7WRzeNL1wHpA
QuBXxJwtfhzpeCE1ccKXoJ+Mkqz6j9005LPHyTRoZuZ6WQzrS99eVRIrCXZJzmY8
9B8ufLXJIkya1gRsNydzwyHL8qS253o0CyvTnCq30PS4ZaoJ2bkcZihsEh2BTUW9
lbN+6BTZ4Q1ea1cDJFFV9s552R3rgUgFHi5wmQ5FfC+TqH/NxexuFMwzocmNJ36u
J2XJleQN8piWBIy5R5HbYYYBRzH4bQNLo9vko4YWzkx88qxBNxhfmxnPcmENNu14
sCxKL4eu6Q80Q0dI91EB9KNlgqzo7hBxXZKO3mj2uZGc+DfMH8+KXhVsdIJShTQ6
a7Wo4rafHhSExHYHMBshGGMLMYQdgdzpLMcDi8lrPCRIYhBXMHnam8MS5lgnK2PO
ZQlgjPJH1QOdSerZk0uiVHFqCh9NUgfCOJcWavFz7AwO9+HCks1mW9UhWnjkFifz
JzzXqQHK1FGDyUdBmeZb/jbCaRqSFTBObR3AzqFY9+HcGdsuDCLW1LpbWDr8A8iR
hXelXaVMyHtiRtxm1pk/jqeRWz5ypC1fXTu6+uHKQ480B6Wm3tlTIaSmUMhy0M3A
YP5fyg5vmqpWroX/8Sgv8LYShMmimX/LFAO630zq137ZQAbbIAsKxVTR4mZNv1l+
LOFyFxZSQBAwefCdTBOLzbjTkwEXZU/ReMaBIaJm8e5Bs1S34uHx9UZK0AE34Jg1
uI0zdU5NiYrRFXXQBUChAk3hU15d6isjxMTx4v4Vrg+VQo6DkqPNssiRhMtJrKO/
bFOQTS37PRyZ2UA0RMeJZ79dTYKUBbvSMOGm51Y79wWKxSz//vBujKGNxLCnpiDM
zg2Og/qFmaenKlsUOIH77AEaD0CJat1UTcmpLT/+QFVpBHCQ0PT3K9CCx+xLR+Lj
LHgEi1OKhCAtKDf7vmJFuNRP8uAPcFVRVBSSMHi7HdCrDHsUXPzmPuURZgPeoWsl
8zxE3ES6HLRfKKweHZRtEs2nSnoLxQ27e9+JCi3J+jr/r2mZCzvE4ResJJqm8uQN
Q00JDvX1hwToOgEw9U2Ah5gPrty5RZs4iupRXcSmCL2LzcCfld/GusIZSgLOVyiY
5pDVeVJEKyARTivdyd8LB1974YKHswa+2hLWVck7g6yQbSZnH6h/ZP0vH1QRIbCo
e82Wx5Fm5kJK78JgkmDVws0eXQM/rQvnX2Tsxwwo0vRIbkIUxJDOW7dblTJ56Q0Y
zYYMKj/FYq4vwC0ast1pQgo9lPIGxmCJfeTmTxC7yAM0MZFrdDYz0+uwoUvgMHAu
mfNx7JVKoQAzYA95fAzr3opIdffQd3chcqRj8XYdG/rq0ISoGUR8AvluCgqWz8rd
smTCqPeKDdMMuiJV8VYFPIqUnozvPAdYlC8q/WsSkb/5aWkP1so0+kD5Nm3jWCJJ
EsYdRaf+5YYXxvtFTUct4Qs0ltTE+ESM4zT9XqjpnKDhKw0PsYDVlA4FTa9mBoX1
AGR4S3aS8n5X53Pnkiq/+vUZKdtu0yesrgKkoGMYesK0anaMZs38jFX8iBDpwQc2
nT91PSHTgPa6qdnpxYWlAXPuyJrajj2NLHUMWjm8Mgx0YbeXy0SO1D9MOm2NpmRK
D5K0AsXuHMVuthwHBgEq/dGBspgQv0gz+olaKWPomRkANSbOxujNrU/ykc539G1Y
8lKjKQLw0673cjXvwYSZ8W0TNGl08U3JRrqe6jY+oSUI2kxlkUP2PF+3GZHHyNX0
ch37bJCrMM/xDo6MHqEoGg4ALVo+EFlbrVsEmrmj4aJ+bsw1ATjYZkpkVmfda9CA
P1w7hiKfmyKkfuPbbc4pE5+wO+ZkfXgOh1JBOwSl5ab2fA11jBbp/niGQQoej167
lchcqLZ1b798ROTnSbQLk5enS++Iu8lCMbmfOCgQsOMKCwXLv1EmgT4SSFi/QQ7t
3LGBtW1ywg91ADHJ+91+6ynDq1pazczWYR/iMkbWGo5htMKtwftGyoXdcjjJr4Rp
OsP2GQoshDw4FbwbVArfTl6HYZ+YKuQjSBETnWUd4NySvTEJMSICMvGYnj3cRYMo
ZOBR+ytR380fVbsjw41S9VCl8dzdGOVPQe7O90J33WEgY7XwKySEuvfnSXX1OmkZ
5ZosP7DlI0fsEcY9Hg1vJzwExIhO5HgXVlfcBgKOzSjDee27M/eFtHRh7/gBjfNf
5j8hcSTjgUKAdluFklAyF2Jmw6b5UfCCVjAJId980B/g64YuZU1l5FWeTiEQDAZK
XIE+Eeo43j7tPNectK1OVZUbMnvQUBhP7B9y5EOZiHhsyrNXdu681ht2SjiC/BmZ
rCN+1Yzjd3thtTFg/UGa39juWclsYOgqa0r71w9HCw3/Mhi3wEB6GTkCZWMxuLEy
4cdwIQcggMVEqIsgRDSJZI07u933LumN2Dc8Wa1m5Uudn6yAW15ZvEQx9rMTIcQo
XcqItiLxbaFxzTz4Gkb+IYvI0ps3R9AS+pFdCYJRiNkK4enRCrNCph/OOsbOQsN9
PoAB2suRYjxMvsiptE9X5m8WbZor6+aN47Wqedf2XhJBmSq2LAcHdldGHIY02T9x
sl9H4YPBrY9tub9DGUtii5+8mjsknvjFJtzqAWvnwcIqQvVfVs5c0JyluYD3iCam
eNAFvzPXy9ICTjuaaU0D/vyrky7YONQOTm3b+3t48RBUjT/xnRsaBRt3CLYzZxE6
CR+QJ298M/Kg0+Y7FsDSp/AS9yDOvgyG9tueuuuraa3nDm9OXmMFsfdi8+d8Bipb
xuiYm21kQeVNapgcakJhadYsZYBW3o0UXHIS8TXdBoeL5G/w8pG2FP29brCmMm9H
LCsm61qCTuazcUtKCvMkQDHe9pABZw9dsosdiaXDFBsqt8ckkytTZJde/Ig9/GN+
566CxIn5yqAdYwpltm8Cv7mIizIXFaNpoua4ZbJM6oOclVkYSG0SZXHgHkb+hm+q
pdUB7exFmGy6Liag7RwN+DiMjH4swb0zqqG2cwB7oa1imPYQ6ChMQIoA0dzm/F3T
BPmK4FHh1JcS/gAIhRpgEKbJOvryHd027A9E18hhizuuXbBAGMxXIfDd4+7sBG6x
tK5B0Ig0cI+mwDOI3smI1646jJ0S+5FYYqV+49pDL+JAPwzEDJn8TjtVqjHOBVN0
tSCmDe0dldkQoVMVuyLwFkSNlQ8yQEZdE+/sEPiiXybH04VZoTAe0rOtBYEH+vL2
THs9hs75BnuZXxXFRHbP2rsWiCOi90uv56+qgWd/WZEiCXqqeGJaCRy6crVYnfDv
bzRdfUwaxL63O1RNecIdkvENZ70pOl+N9kHgeQyKj6h9ksZ0Ql8oXVa3cpVHANlm
pmze1UQ2nbz0HcADxX2VglIrUEjbEfjbOhJ1S2ODTdD/Vwv5lr64YYzfPKflAxei
UC0osPiM9bPFH/ztZajwcYTvxClo8WRqF7JsXFzHo/G8odZySkh3P5kKe91/Uh8j
iEabPG+GMTPyT9WBnt4mhZDKGGTIY/rlmkvprN3mtLlgkEkU4PGp0/w/DHrGyEhq
JhD68Ku4VzZRXTyfu36NFfX+OuuyEpcm2sZElA6AA+oBHpxHWlypKb7Zj6fTNHDH
N3tBfWouqJr04FuisS5Z6ckylqFJ7bOhepD8Nm2AqJVhCjFoTd6Ir9At/LCJegAm
a4asionWj6vcuZVue3oOVeBKC7lKUHKEzM584RaQ4U5NkNb/mYLfubZ1f1U/JIlf
fbTGMN4w6NciX/go4GyR9qlAFvcRjeqKp33w43N/qyTAV5DzMkzVLYPEwDRDD6bW
FZa07MTK5s+PgnqD/4ZdC+gorwXln1H7LaoFBv3iHFxO8chWFBMsXt/X7fCAU804
iMdrou3FMQbaqXIUGEi5JaRxkNFBrDSZPKEjUP1jEmSYhrtOLhIIIaFoGIUsrTlk
VgStpRQF2nEPs9tO20z0iDalyYciXrLblSWuDpoEcIo47+AHUzDFT6+tMgmIMT4u
uqBRqDmLsRt1kZ9cQHZG8uiZhr9iSUhb/CV0z1dCArIPiwYYu2AevXrYbISMw8iZ
5h+wLi2+F7BxNa3CgDCoW8CxNe7bNFttjnu85IAHBy/dAJ7ZKEyihuNraXeeOrey
XZItws1INlWJG+Afmr5jYonpeVcwHrnKSa3283x6gihzbTlQ2alszqHGmkBuBXvk
oLXTKmj5QxD4l6p4CdqQUCSFGvdrk5XqhanARVvfmwc9HwfXx4ipXn0f7eDWBCaZ
Yx2kh41nVdTEWnf+b14gsMI1hYc3nD+Gej5wgDYsgcY8oE5DkVOdb6pJSOxi3gKx
28CBBM0ONpeKLOF4tYEipA54krrpoML+Rpwnu+bP+IkR2X06IyoEi5PePrtfiqhy
AfCgy2oVC6jKlmhgWB1l0EFe7wGU4g242GRVtz+XNOibQvG7gqemhsPz093kRB38
EwKz2odt+qTrSdswmwGB1sFyJQgnJDfd50+9g2uvU6uYuSZ7RHU5CgpDjEqOOvPc
u28/vTIf7tpHUjpx8YCS8W2llQhDXyimMykrzBFYBrcpls673c/fbG9OxX+IPkU+
2oNEN8lYEdw+2uN7xVEULYwVYCwTvssIzd6S/WVPWjcWdoPAk8/rcGK/mJIoMgpc
8Dn9iqGTblDoowYP4LMT2DDEDnTEoXvfXGz3lzijkmyxoXuIG8Vd025h+RQR4zKi
7XbueDOlpR2U4gzTm3p+lV4mNlbBiwIt11P3b9MUeIlmLlkPuIq/Uz2zobenUtzD
rvy2O56pskn003Nlf2vkxtUjjlq+pRVG75UFzMvzRzTZHHk/4i2X6Zd8B+AGc5C8
EnI/C2Irg/6FJr8SshnxdKZfD6MvGqVaUzyhk+6EM/3aUAJFfPkNHj0QwACvqMIc
lq5aw0W7DbNPp2vbngK1+h/dk6HGnLx8cUk9AQ2iYYoAi90Fosljg4FEdAi5lwYa
jhsA6DuJU39v65utSBUpOaQK2bTRdJCZxxqU/pMC5biW+9OO+zAeuW/PIj4eQcis
NL28rdzEQ+VHKjWiUGiwHEwA/rj0B422iXxp79oYrH6tCeRzMQ++fj/Sd5LyWduS
FpO4ogrTx2/BTcE/Paa+AxlRyeusyn5k/qo2HwdHGahjm93rXzMikcnQ3QVhlel+
vm7rHcfzW1rf8hGFmd4QbH5kWGF5mlg8DC/ahK4EccgvPQIYUNl/UDhJ8pcJ2vpX
ty+JfS5NkjVnSnsLXb/Xo20/dtKn2YBXlS8NfDHrQUc2y47tEGPnopD3ab8DiKE8
c5qECFr9VHKTh1MtT2+E0WGVv5yHQJy6fs8vtw02X8YojTk+hdbTPJLhN2SLaB/b
SzapFGcpArLxlZ3Fgj/1+VzN3+O/7jbg1PQ3gSjDKhL0SttJPjJCHJ+MCI09o8lW
64WjSTU+hskaIA55xxFzsxft8lH2ASllL6/7AbAo4sT7VjIJ9/IEyeICHg9RMyUh
OU8anrPpHjZIZc2jWatpUVwI1pkZscS45VOg5CQdaqANa+Lnz1rPr6wKV0hZ+pBP
iOFDbqDYp9wU4bnZG784qhV8345OPAgxKL1gJbaXaYkbEKMhj7knYUmf6zWL4+Fd
EyHY+xqv0bPHvF9ntYCRviv7LGerhMUB6cJmm8fIkjytuJQF7jN9J0ez2S3MuwK1
awAmD3suDsSVTO5qll/Qa0sfS5k/OgcBa4UqL/VkJH+IbapwZ5bc9Msu3eZ6t2Ui
BRgaQcV8cFCzVzl+ijSOHphMFMi3nX4o86r1poan+izVA+LSt0GPbp+vrtltIpkQ
4lV4TiJhKVU8bSfG7iag0feMyoTrw63ulzHmbVCE0CyIyBicQSRhZdlbwpU8gfm2
wWATacxo/UQ6rXzP4WvBWXV3i7WOFSBWaL+PmNHLdt5UUsWNg2/H74ZGe6TlnAyw
OtJ31AyHCfSQzGm8DL2L1xfphJOlK7K4lWCAVn76O/a7mOU+Q/qSeCvTPEV6083E
jPdRl/1Oh47rbbCzWs5/rY70z5pOVF6Ns5739ZcMhriaIIvp4FnyUZI5wpHJf5BK
GjSHnToCmk3P8M+fdVh/nRnM2ESGC/LO0qJiYGMh4TqkgiOOOvlLrqSFzSBzqD8Z
kYpEiMPfdMi3hwXCqyOJ1E8dxZWxX8MdjVbWpwsyYA8h6EFZ0pYeIz3VDEIr/xAl
qwmd7GPOaIt9y4LR3PSGxgdL7+XHZRWvOz1EtRFDVdkrwrSaZ+mv3dDCgnBOJRu3
ueOQ/EdfM4bBNP9UsVPYsConRRUJk8tG2BahWTxNNsXyR1c5/Nwg5duNhDsT6g0q
YE5026+gsEyM+Ya2v0yXQr+epY2VvaP9z6qgSkmnGn5SXM4+68y4xCafKo/CP5OA
aNWhhM0i0LbPCvgwTmhwvNV3LITcYsJsDRAxejlovdaX6x40mGP/+lCgRk3WnHJb
CnYiz9KBsMkBxKzAekZQhlrVr8PYUIVj/por7WfCvPqRSv9tKuNM5Z2TMobYbYX7
YSEgeEIMuCnfPjc2zb534yAqLpldF/0eJZcc0A+KO3e1ODzLnvnlsfJ7+fSKx1nV
+uVa02yyf81RfiaWDYQlo1C8WpTCVwfyyvmzfzz0qDkg9t4NQkVYU8QvUp2aKhID
AIh5QrqfT0mnk0AwkiQNxyI1irNoI6HZ1LVDxPMJOKN2BCH8VVtcU/B4hvvtii3D
Y+yL/JaGdhYAZSU/scHdn0XtSncjHj+bhFK+jPdJAAiobcaFNmRrmqDbvUYvhkUk
saFTdMf2Li+Th0BJPT2Nxc3dMC8Sj/vdNgXu66E7E82zCrQDu/dth54pLHxWBvnh
OFwmEjYldwIvKtKaUxuXHzAraalRONMXi2ofETtUxNsR6cFg9IDKF5Vto7r/kyDY
UdVD+k4GM5CUHlmDWf5mbj0YKaaBbTamt9kmjetXW4EJ184o07mA6D2lzEKTmOqh
5n8N+fr3f9eAnQkWTGeYPochB8CD16bTRyDbVEvDPeIj4vR/8tr39tmUtDPkCF0T
b4P7gql1mIYtGR5yDbkMs0yITY9OyqCAuuoh6izSY5IunsCPlhFPqtechEy9pcMf
JccHDoY5rS6AB1uOIfDb61OwqbGFMKfNotZn4RkC2TN7W0HTRYui0je9M2Zz05Sm
Scotg9COBEBOSvYU98YjD+Gs2Rs92YZjo9MOc3RvqVxhpfKeTxDO+ErwNeLEOxV4
NRWwForZ+m693RZdVefpIgd8kqh/sU1yXa/sV0LLm9Mn0OMn6ANtUzu2aSuZHuR9
oDzXiB2i37qj3LENmyChk3mixDaEg7bA4BCykC3wQf3T0WNl0PjtWdMn4nV7r4Sk
ClD7CprgryiRTPcHqpoMahyHH9ZtI8CCcNpd87fZ9rQx6H3kIYH3YuNM3f1YBHRk
Lp3erR3SsTrqCO/uiC57zfiGrOl67fb3JlH9++i/hUWeCoFAQsa00M0FiCN0OU/z
VpeVwNkwSY8tksVDEAZgQslc1SEVaZUN/10y3m2p+xd3vEwZXVgCdb1ocTTD7x/q
DDkBGGG5vAzCJixtXi1HhhcPsHLEV5xpqiwdS5l3nBy4wdj9mt1cTqXjUvq4Pkfs
UvDH+ZYzq1AxCCsD1oX6009Ga9s9T2EHp2HVZ1rfCPbDjFqY5coVbHrcwVhw+1BD
0XbEZ24j6LK1pFXeM4ryYHUQzaUDajb4FJsCIZCQ6UsvLcgRjeR1IznB8t7ArVf6
7KmfqOkbF1LrcYnvvqpb8j/arDTj8PJzrbkQPOAQetrW1wCRBGOOXIXIJ6etbWA4
VctEXC5axGd982FvnMvS+eIyPmhHYICDwaq+Vot/l8s8Yetmd/rNbbooBnQ+hypa
xI63jBKvBV63UQxdIVkTtoH8sH8I/o/EPBR8+MMjYUZrYS/g+InfwBqh9IfugF0M
2cDjN7M6kmVP0SuiP2oTWbI1k1YhY4iCoGr3uUWDXtKGo57Gp+ZR7GyyKygpKsN5
oGdYOmhS6OjEnoHtWvmZfV120aOVc6A2lhlZRkuSwP51jrl1hSwlSQWCWvKAxamT
uHANEINJkrX0u+SVk+HMn53/186Krajwr5gm3IuYNzHTZNbsL5queWjF2YfUlRog
Zvuudp/jmtZqDmSkmUcV+Ut9cNz6IKoF8jTZwlQ1QHFbc5k0cr0N57Z7uVti/J8T
49JX30h18lyFeQzyOXnhM/1EKB6SxRDoYujnezdS+GUYPxCu70dsbKuOiHaq4wa9
syVLmHUHlOzt2K+HJizl4pvFF5HJVx2xYHXMoAXlAvBsmExIgxlpgQBGKtchhwm0
zAUN14wnTc35Thrl1I0XHx6X/lt1iA+yjHUxLp+HxkraWKM8XvjDq9wj+DMja402
SA3FT9zSk9ZkwcSFwQlL7ddEanrd+UxNGlRTBMwTUk4OEDVSj6oUGaHzkwb82sn7
PpLDzYkXuZVK4NfFUWdlShMyt8VZDeLHseIWLYdFwVQNseB25fBSl6h7lQhKFaSl
U7RWiyg3Xtu0pQyndOa+mDPAO5jrWJ07Aw4/ZfGOvsYAYZhZByTiH7BIx9Jp3YLL
ck3y9iKew8ggGvpZNV7YsZD0ULm5ZUhcDBEGRuthM9c/qx7IpS2wr5gDZbRAL0sI
b4zK5KPxzwfOBw3ZlVcyoMKXkgdJafzLtfEILSPAZJbcxYMH7JR+UzeLl46QezOG
A/IbeAT28OAK3iUhK0w2tRe6dzNG8ksfAQP/qIF1NWFt7877QlQ8lHDhShdVzjYg
lzPTQzeb9MakVlqgK51ag70SXCavdsP/9OtiSy7y0YL/rRqQNiKjh/z7MtuX+D0i
cj5oPPprNLaKEpR+4Z5AWS1+Lb9UnRDqSFk0qRrxIg6SedKXk59LVAIOpbWkKT5o
JbIUppPemAuCCOBt30ej1yJXBqCXlCQRWIz9Z/JOB/KCn5s8NBj1D7teBCZvxhVq
WjFiUq9aXPpFgoi2adGD1FeUjkqzPyLu1+7zqJHkxP39ithTdUHRFe7Ip30EY9eV
HhxZZpJu0PdKxWnAh6qg1O02QTAvw88PncUhxf/XEU8M9hDT9r6LJ+TvovoSJW6p
uNGfv0xlo7IXxwQwWG1xTuU8XpRdcWJ9+CCOunKY5oPqWJQ9m/J9VKwZgV30BIGw
yZ8403e0cZdypdgUvngQaY90cyJoO1GN+fdvc+mtuUxhvnO52a+zCKfctcRRwvP7
+5uZQ5CL+Sg2avhfbZB0W1InQisKpyyDDWBBsk9p5uEDyoqAWnM4qRXjXMy/5/8R
mPvDhBu7U0/k1s+Beuxuxt1FgAdOTQFiLQO5kYCuAjQ/HLcbbpRmJz+6vB4QX6VV
8sE5H0ELtl4bRTZJgESiUw+QcZCwZswDp4qpS7rFYp0GWNYDjSWgPxPY57VQUF3S
HyK6rNqRQEEZuoIlD4L2PTqm8pPzkI5Al2Tqk9mE543SZYUtQsEXKfZbg0nDCWZs
p0glCSoeBo3d5kSazog5K5bWNHBXwPLZZhdRUkgDfb69Mf2K7VQ3nV9Bwqyw5/BH
NuparC2VCL3qM+RcRh4iJrkZSpUSCeZdrBsCEGq8/sKkg0H7lLuDDVJq1ah0EmkN
RTAC0+MQ5R4N6lXnyHtsY8C4rPfp+6dolb/BAmbq2Prb0knXiMNp3iSI1inG39p5
34gZx+sNX1C3ou7DRVfAijFG8roc8RPKoQUFFnYpz1khZBlXw8nC+jCK5dSEaftC
uX5dCCiU/03IddQADQG+y/QKLhoxV+ValIw5veppRFLQL05rGGPV/5gatYJ9Zxuy
Hmbq5jw2u9yR8jK4aZn+xu2AygDiLzMurEPpVgkgL6+++nEenqry5a+5PS/9P7a6
S1GF9+wgKoQeEwBsjxwunM/NKUhewtT7VjvroJcqa2NW2lFT7unaX2fB5zZ0aXuw
X/GoyMoX1U8vzfNDvsu83wq7AT1SYmnD8HVzuxUhcnBw5zlxn3SKHNujWs7tpFXN
+y10KKE4nyPKa4lyjTU/j9o6l5IZOZI2y5p5ramQm6yDNZL11tJspsagaKFIUcDG
39tSloPz+9zRFS8QOYBXoygMqb9U5LM9liMi/7eP7Vrj9NIuwcNAbSYXi6iIFpNe
VF9I/t+G4L4CXiGo6pP/p6gY5UAZyCMmVy3cB4GqAntqfH9fIPyo69RXPdQCSrDR
nOdpLTj6hkAJuUx9n9ev/1rt6hLPsNvV3Fu2S9Z979Fh3ZGpNDIYmMPs8RnOb88/
y278/000R5WJPNRl36pzInbDJrut9UfIVui5c7pO23Ws6X7eeelDY99uawehdhsl
t3DjmNSYTHmwBvhFBxiaLhb68cF+ODkT3sVMtVeBzkqWCsQf+infZZQuiqoJGkFU
d4jqibNTh+Z7/n3WgINp1elh/rYNNFFHJEaNdOGwtJtTqQXWaWDdQjSq3s54pQUG
gqBoi5Jc7Y1wwPBrH0EHV6ohAtRJ1eIgi/HzxbwaU9my1K8Z+CnQ5KZ8O1h/UgZE
+rj7G5bJRpP9jhTWjuSkvfQMMDRrAVAyZmaK+6PtY9JazxVOx/HhnbSeCov1aeBf
689vULt+Gy6+We8wtN06l0ZbrtlS+/ppjjdaASwRW7m7DnRfijJzFPAaAwXymL59
fhoRUCiEQeKGhqx4WsFlyan75CEyFaa9UTRcS3EDkJgFp/pFGGjmXCju7feoRSOi
wgA3d9XhMkkdbSPKBCMjlxWIdU7o8Yn4396WWlHxUhXX2H+7nvbbTgOdbP6jXIpv
DQ0iL5dIeMJG6lIAZtfSA0q83A64szwlM1hr0hd57JJYUiWNSvUDmRPWBb2+IPTX
ioLYX2exe3cWx3bZ9/D+pydREM/daQ7zUJN+gK0Y6w6N8ZnDb2t3KfA6VRVnrznD
hXwO2WCPCSZEXMzUxYCSCNRCmseQYLXtq1c+grhEiFEhpRsQYmG1nypSzUjDwHKV
0wtuvjHCOk5Ilw5MrtARRB2N+FKUbGqfODSvGbm22C4vBVPU1cZkyJmWRZxU5pQN
4xfr2P6UZFdMOy/PDS7IGKfHmHcU0Ux5IG58Cy5tKfnKo4/OtoTWKNw0WpF8OCoM
L+oPO39pO45So6peomCc688hRP4RwxPu8j3uh1oRtut3/rv/QWrPViwc9DNFISag
9RZApqmVp4G7jNsAzZAKcCD3SoKDmeJaztRUSWJg4ivIicFrvURPHayOJp7oky0Y
4mhN9v+9AXduNOY1vI8ypjrSDfSeGuTTrjCSPJ+YquxiCCr8SGSqoW1HKdzFqlMi
6TeuT06p8OA70EvwmYqTWhrHhUBdf1A5MzNJJ/r3i/AKqfh1cCDrHjd5f6Wyt3HI
3rCSHbkyu8TJTkABgAO6dQ7TrbL3ivA+ZuLRr33f2pQewofapyDy35i4hz4qJaRF
Lm97ZcTIr6QcZiHPrR3MrLNNyIchCYIdjhriPwBQTlbu0mdaRi5fuDkX0j1S7ZQI
uGVEW8pTTxOyEti6/bzsL9co0OemCVr+VEstK9E6bcJbGk8Dshw9P/0nQpstwRNo
TpaMpqWeaqfnQGUnxo0gwI7G/H9fuewtQUH8+3rbquaWCRGlo69UDqfWToo4e5Ud
zkQjXh6sG7IxMQ0Zbts+FsJycEAysJmlJqVmAyDa/KV/RWh1FER/Z6a4XPqfwv89
/RwN2B3hCC/7ZV20kE8+S2+kUXGDrJKGdhgms+kSVENnk8I2kXPT5Zze1WjyPlj/
V4gjib5zlEQtwdjsXfGpJRsjZ6IAGKACc10wL1s7Aet4tZx1kjuGKvl+kVYO1wME
WN0jAo2Z8CtzBTZg+UtzlX72HJqA1Y6zpTtcg6/jG+ALFpi3DGmsc8LLnGiu6v7G
2HGajqfHwEM6UKOW3GHsExHWIkraVmNW65oXr8zdvpQOycj1zZut2lQ6YAmyXA4R
KQlqHvlY9hhgBm0OwPaxIbhA2OjQP7FPy0T4Aft0WJw06UQMZbFoMBjJzpoqCVs1
T3ojtf28AhsngZ9rc5tq0MAhbNJp4yh2bLwxbe3pt9CaU7jQkaCViaXVPzcqx6Or
eWjifhtA5bB1f7ZY8fawXNy9aU746yAAgzil3jSEPeGH5/3FgquASlxoVlx+SANb
XIqDj0Hlz25hfMoNUreJ38xNUNu5a3qfyRAVlT/D4voHzQork28ASLMRq7Z60q33
9907N2yIiFErOR5Z1UoisH3ZcSeqUv+6pQZIoLcOC25Wexch2drJn04pl7Niktr1
mYOXHvkEgAKfuOMHJxZYYLpXIodDNxxVVJxo83zTNIELVNXCuFBtGDlq3FzJdRoo
Z1+uQ0EUhDpKqC3sDg0h7AYfNTLVLhHM6QfMzzp5dTnxH/TWx0OJRbkkixDCfy2I
SSODdeC51jMxlcbaSnybV3fR+eTib8FQpGyld2riSpWE2T6nl5CrmVzDD/IwsDUP
AgjlQkg5H770MrEbpsze/0cdgr3QNB/zjUPZ3X+I+pveZS+5E1u9evs5lVBVyO0K
/u8ogs8VV4ffJjVmBwuOJ8nLLj9b7I62KARqYwN8U3omJ0Nf5S5NOQymh8rt3q5E
4t3EUw/MH5VAxVYKCrCnywWoDBYrqyZQXBZ4G/hlftdaH/oUyBZM/03Lf7gd+cLB
MAJURZXwcGcYl1fWLihNuJ3+57e/uj29dd1pvQ5QkkwyW+2TgcGgrclASN9Oavyu
qHFES+zn1TyAgrKr039z7+xAwk9mMXRAB+URXwob661ZlwN5mzv+TC6B7XRb6f66
I+7zEPteidqB7JT8ZxK18AF1o6Gs4UHwve8291mXLZlLbgQPeEUq5A+rIcD0RfG4
h4JozxKmYYtauUszQKU9Rd6C0WXX2WcraZVfdFNDB0MlGTYkVLdpkMlbmnG32ca/
WWLv16p+FhJNvRPnvxEXilQeWE34bB1xQ1xE610hfmap11qNHKgTu6LD+MEUk+vj
Xi4Z7EUoBMzAC9tG3YG+4w679d2U9TMycOvEpqnUoc0p9S3+2k/EoAKyapxNDp41
KiM9XrP3SXiKjK4E3SZXjRCE0tO3cZah4JnJu4QxL6JM7K9oVyXbyqZZp4gmC+Dk
3jdsfY6WWtoHmj6EXX5ISwEUizxZg5a3vE8yhCBVK2rrSM1MiVtN4SaBiRyzU0z4
vQFVa9vnOvDE2Tx6H74O7LUCi165qBDArooe9e8eD3z6FDC83Qc/gxfOqhaP2/4F
E5bROTq0HUptqIIR1s+0Ts9C3sHDFyYw/HbcI86IqgcZJ/rzUkMw+f8I6877GNXi
3DVpKhBb9SMp1dcO7KYhlOnGruw1tM1Y4nE/pYWIttjXzm9peERn3EiEd7ZGn1oN
oBje1GhsDehPg21gUeW7GLgUHsUZ8bYZAefL6YD10D+sOmjno8pq8ubLSdkHoDmZ
z2RmLL5BwXn2Yot6QtmiR3C9jFtzuuiTUC85xz5CZgJPyLtRCGZAHtep3uCckUDI
t1Fqexd8zPmzuqOyD7CQEsKAA+wF3PIeoOIxHqbv7gAs9RcaWty2jyWlJXjJhKsh
txywlxbgggKsyJFdtg2Z5HpB2hkY2myZkIoHTkD3J1ldFpRbsIsW0sDE0TiaCkoa
KXPnJdBC//6s9t3l3HWcf2yHtxCzpmIV/x2NYy4lSfuQLdx0+f8k3zk1i1CM+yXo
hpd4ZQby6OxE0iXIaRHTvUsDLxl5v3FJXg01LFV8DR3Gdxg/GYhC1ykIUgFe/wYk
rsOu2YHU7hjfpJKTD4f9YHZbxoJxsdM+rJYLxytTIyAQVBsUjbGc9PeXoXRoOLa6
3srikecTWaKG7HKRP3yNmYXspRCGBnly4P7gFb3Z6Y8n/ZomymL3xhNJof/zEEbz
MScXxHcOu/ksPlY8olBLH4NmicoUYzothg/8tkk2dx/YzTMaU4N19qBFWaZ2Z0YX
v8GNLn5nvhYzoKWS7sv47BWaEkgdhXOT+7U1igQ/+8QYwrre6z4+/RJCZLP5zlbm
cxj68ungpimrjAVDVMZpHih3x2CTzfGohosX95+MVvwciO1VhfrQGkUPYoqC2NVq
EiP4pJg1WqBzBk1qK9ftl6kMGsuqpPEOV/Q8WZbcMuVtp+tZlzIBN4by7mWMwHzr
Ens4y+eXa2igT8GxUhDrBwUDlN4jrFuSBpXquPAv00WqgLyDtTsVqfv/0kzrbjzM
hElBYUKw5gVamwfjt2mTc5/TdQPOWWeDewWEkGAg2YXFM9N334Y8HJKicLAYFVxr
E94f3ljsJVTTwIA5XLNPUITJVARV7hR31n79h3bvGMySoKPLRYfVvVD9r+RNBh/w
1255ajPrLd/TmZdleG/bTxK2kN+1lxX1/ZBxGtlSUshq3Vh3VsX3IilRdzDgKZ5t
DyU6PQYzvw8GkmQVy+gQad/3fqTPmNnJTnP7xBZROUdNsYVGefTTOKX/h/uXDjz1
n/Ei3sIXel2J+BOpoejM/JXAsYlLm811lN/slYdHC5yFdO32LNjwpnOYWVzKz948
3IqFZqvg6VTpqQwiQZ56oP0FWkhQ2c43AtwntbVpWsFsZq/a+Q1CorrFdF2maQhu
rF0zwCg6yiTuHnO8l5qsJ3CpGoZU2Qgsl+FU5pS/QReKqxc4DXYJypwHMKcP9tnf
QqcR9ChjMddODglgLtOU+vcoljtaYjJmTQCQGX/52Lv3QwmFqCwBrzbWWEnn98jb
laWScH02iYrQrEKfAegIGgnt+vwx+8uD3rZ6u+kYnm1/L4zYOobI5KbWtA0GwRhq
YYPgqNzpLn38JLYhrmXSBb0gt2owBO0sijDzZdXx6g9dgY4v9jT7pDVDH44/oxOl
dHZ66brQhqz3Xau/tkvUTfAY5R6eLxgyIhFqs3lEQdWOcIDGWCCRZpLUgxNXeijO
omMZAYqsmjwsLiwzHMndmOxGi6S16EjbIxB3vJ8LoicscouL7ScVbjfFAZohyBfZ
BUmP2uqkBwM3bdnPeWfJal/JpOw40ZfL+K8hOII3VT9gcBwudkz21DcTanuZw4bI
ZyuiWnCx006wWuVBprOVXgagTdF0oSKaJRfSul1O7opBHb/1Am2nw5ybeH9RjJyh
AQcV1WztSoRxy+FxMvRW7N+y6+Od+JSIipCTxaRx7/lFvFUciZNYo1sfsK0jxRqv
BXP86toURlQHiwkHNvgB8zu51n9J7idlbClm6H12Unx8WY67+c7qpycT9SweGQS8
jA7HZlwdEQokxFAKQZ84Wdbq0u1+pZhw7LwINZw7q5pV2/rKsNWigw4Q8/F9kAKH
KrtPPxtvI7+M57uKA5cTnkdTS5Mjk1+nV+Q2ggYNTBGodtMPICx99ye7P3JqDJeg
U/gb16eQSh8K8X9/Y/edjdZo0i/xMpoBcKPBaPWH+3vbzYBxN7+LrgvUlNayBygS
fO3A2qDR2wjPeqWUx6otPZnvUyc24LiuzTGC2mhAQNi2shm4sD+N3uqyM8Zpe7qh
/Ig+zrWZOKWdYBgOAJjMmGYnoVRq50f8g02SGxps93e2CW7c0m9xAWYVQYKE78W3
PmPd7baE+zIdV0qsF2TtdvhgLVjp2o07C0/waU+rI9aKl05U9VImb3TxmfUGlj8n
lwubxJqfZtIrfMAgZbAXtF5AoVtGezV/9qtK2L65sKFpBjQiDTAlp/q6jFvGl0nR
I61dohkEzavrMlS2VqDFtaACCerlcC75F2BwPkPMpbd8xSbN87XXZaxOXVz4Dinf
Zay17X2AwtDiIpjmTZiGVjCELv7magquaN8D4kTKDRTioNqISlE12pfAkZTRE5I8
f5YoIkqpdLMAADMQA5WfIfhW0iVai23m1BOZOYQ2RISTC28uCKQzK/UMslV1DyII
t0Zze+iDyXVvr/aZ8Gt5c/2UlBk7VHk8cE2G1xLGfpe7Rlkzd6nUo/bR71v9fEAB
6EXiQSF62If38F9sgUT0/Dq3MAx5g7gx4PkHpxwltxIiSa4NJwCtnmYJrsPkqX/+
JbsoB1iHhyHYsu6IpO4VNvIrMM/JjKJCAjmC0ITcbL6f7ISuwhAAQOg9xHbpcok+
PbtCysOGVAtGKt9OBv4v6QCdjujIh3zTG6DI3cshHK3eAubDekV1cSiP978wszFu
hiHwbo6ne6DAsoLb6C/qZNJEoQszbY3/TWhpa5wOFt1OrTX7IC7hpr3YVVbVa7yP
syNO6eKJk5PXwHlK+Q64GBXs1BKNFq6Rf8SUq5QalRVxou9KDecnMUaYAsHxIbB7
8RBUoW4lmCiCvU7wvdoqIPHOc6Dhip+z49OHLQbwWB1B3VcdMBfThwhglPLpMvSz
VOu9WNOXjbhCwDjevVXxA1BQ59CMRGgyaWgEv8w/WfI9bvG3o4FOm517KEnLTQzf
Dct7Oq+UWUPp0U9i7ozA3pD8p9fH6ehu5Trp+DI7TncfExGEx6rtcsUZrr4oUfC9
6wjqaSlKgF8sRZBtfCCbdanmPXFLf+X5YtvS+odvaYI0NiWs4DSdE3pXv4A/RRIW
KtdlZtpOf2j6j0Lgx/SuDK0FtKjZUrLy67E19nekNJcgVlmHDtKSW40wjnwLSpTY
sByNEpc+2/8IVaIZftnEryRVIzHED0b12qShRTxbT9/wocbvw9ZBTYi/SCMeKRV1
g0eIBhWLSw+WgIVzpWCpDL5ROC84f3H17YjXa5Elh71uAktCj5L5BG5Vcqkza0aI
a/AGLhEy2398a4dW1L1jiO4Ii407XbEOspnh3GbB/QeJS1O251R6ugUncgHBZGyk
W33ZgA8PJSrGZ/DvNkyciyTGpaMcb/p3u2hlvH/0ntLzEDZ7F6nEsB8cMLOjcWF8
ug7P3H23PU2BJiYK84rSTr15gojslxcwIpXuy2PZA1N5yTi+pggU2wf57z2rBA64
Y7d4fBmlyjpRnat9S7MhVdcdKt9/CGJuLsp5I3nCHUYOmmC1V0yhLUmwFRis3rN5
PdY+bRJH7/Ind3CcJRN1FohRQpYHZgEvpZ8Rig5TtbSRgsIA/B+Zq2E6fxc92Zcm
R5INq/6Z0fUVpgRXrBpFRzn+JcJTmnCxNqFW+5IfNaMGzok24GxH60FO8cgJ0iqJ
g/lYltHVpPoJTQ8CxY5+4gR9EeY5hPGNbLgXZOIMjzZAlVaX5CHd2yHd0+PrMJdT
eQwnneN95Sfjs0t0auDayqgxgIZZIXHQZJ0XksRrRCwfHmERDega8I5J7amLRZJZ
MY3cxipEbNF5zR8Rwmwdt7tb/mZoU2Y6uxCoslK5Acio4g8v23Uc5tleh+FfvX5A
vxwSDjOxjfEfiI9BVIHWh2wQzu1Jhe8EuKJEjRswWwcri66xyvicm3gRtMlMAav4
EI3WNOHlHk0qY2XQzwtaFPld8QZHsCOhu68Te4MTf4zrxnbhm6brjsqtk5117JjP
VvxZyapqizfKRm33xbAsG1n8EM0hwXKevZ1gvJjQ4k3sOaz5x4DRRYfmdpwZPMBI
vMyTi9TLnYN19qVwi1C/VtTYwY6CvPvlpnCpUOyDoQESYwtYGj9Ws8UeJFPyhVfK
AwbetDyvqZ3w0taPQeqcorFn3gfeuqbhbJVtlI32FEoCdgpyOnNxtGWFllLl9FOs
2YOy4xa11yDxgIuqLb2rIAikmaZhYEv96G//AbLfwMfgo2YMtPuUOKrU3mpiAf73
+w00VW1cs4DFp3UJK1rNZ6bGXyQdv5e8nnpDxc+O9qrBkDGnny4p9JmdbyhXdkui
JYuUnVOvoqd2K1zecuqEBWzjHzJHgNSdbfIOB/jfRbELCAwfuYDVy+4xaMDTFNqr
l5fMBzo+s/Y/GugpCCuuXABWHlAYTivCLvmikF3DyC3L5Vy8C99MphGYDWjOsq5s
3JzGDhtMPZ62WhBSmtWGqaUWGjaL/EBENNA19+dftVAzZ95sep9bK/livpxKd4g+
iDeV2ReoLJvWnsseEasBkmsMfyPu6YG/Gls5AvPaT70J8CnBCkqSBZmqP/zhJc98
CUvs0H2be7/yZPv9jLf6j/B0FEz/YEOz1dkj0ECCkL+Y4qrGzovs89pd76W/GV42
7Xt8pKBVNQaaLPI04l3Ay6EpQwbhnv7nCwWraUswOWAjmtcJ6U76I1WbKJyDlyuE
hfrRMtVnMOQ7k6NBlR1XE4QaL9SGDayAa5xOep0cKZukQffQq1tN6Rp6o96kP07k
nerNbio1FQwoWKEAdCTF6ViA19N25MEWbR9zJm3vaVNJGds16W8nCRLSt8rB9wPD
CI06FoScHZ1HXhlA1ytsDJLAr7zwHOGkcUjGPZU+P9s5PNPDdlswbpPgkkU6F/Pl
+ZNFN0sO24Umxzz5waDYHIp0nqhSrYIMDw4/25rfULzw35ImqvF62O4AsCwiNUl5
/LupXabZ92yJPnMjH/DhC2u5ce8O/pEbcitF8uNBquDomQ4NuAq8HUGMfcmg1rT1
AYyLPgtYMb4FYWz08fC6kI+gNh0X2aZhVpEvrSBnhYWCcO2uunY+PhfKuGDXlKzy
UYkmzMLb1iF66XnG67YtgNopgk+n0yVgeW4pBdWxllu/9Zgq448OuezvI//8V+Xw
QqAyhwHj2ds93PojEdWSMl1xmQ1MomEx1SHn9RD98F7J+5h8SU0uYHYlykRlRhMl
p00nR2h+2tGXlxAaVFHlsTp8AMdK2ajP35SUnAULP+FWSb0k8u4DR3aXmP2w/VVT
2Kp1/5HHK00nYusC7DyqXC6Oxxv4zIu9AN/XuS8tr9+H5B0MLKSK3LokltZkm7aQ
heuaXwjnM/Rdxt5NBkJ+krMaWR4xnyVzesVCeSlXECGFezZqv2H0rC6DBLoGbZrQ
u2je9dJxH9GGbweqjfA6LOXG0V/GVh17mx5rFTOMm4IPjfhggR1IvT8tNwD5+cvX
DgK2Nabhj+za2tyxtXeO8PAa+PZHMkR+UQYpDvX2x0mO3+le/PQa21n7VU5BFgdG
tUZ2KTlxbC0U6wSJ8KpZRzMlQo4YCLs0+Wv9EzcWE9Y6nSbwlDmVcMQFWSCwVvf6
5KqRWLP9CPP6f9QxrKbtYSL6rF+08aIKFR+7gL5smfpGoMp/45zEGYzALLJLowjz
WGlPOnCRF8whq1FsJNbhbPh5dpQurVR78jTRF513FTc5Xyjd/kjOKWKrzRLaoe7r
RSxRNlQl5qlEY2THFt8phY2WGoGJIsDB6ENGUSH+hwjSkj8jV1rS/mLKq1UqeNgx
JL3PVVFCbJCZW70JmP5p8WbFiBBB8B0zHYOLGhTo/YM7677YJa8croD2rMrP+5lX
fIzVc/RFxCyki/swySVelTCNVAnpwxX2WeDx0UtYE89IWS/K/ZPLoycvBBZYuJGY
bDxeecf+wLoKToEyRjizeC6nrkb9q8mluux0kzuwo3Q2tYvQpGAxlf741R3x/8gT
TLZ7GRbieMWlHmk5u2p5nLtS1AVxkBfxZdAejd+SJeDlYHTGtM/u/hq4GD4No9/I
e9B4kFZMBoJy7+0uVwmd3ONvKQ93NOFNbWYmf5Bgoz27DZH6pmgOxnHcz/FjMRnj
0zOll2IeY5YHCdZTOXclnYE/jggl74HBdheJ/GrnWb/mLMvOWBhgbjPvcYJbhJJn
54+BCF7lb38HXcPH88GzFiTQJywRS+w9dJ++ai4xsKS1/S6CsUzhKDaav/kM0aj+
fH1yQWp2tujL54Mq+M6Tm1oBhq4moaQ/tf4Vky/X08rg6atSJBlYXQ4Ps01FYhOI
SWmbhnLSvVpzCdjm0ip80u+hoeV4VhA0R53j4VUK8C7qDgkDHfXsCY6uRPb1GgKF
4EBPag/XyFpZi2w1KL4Ux/c/q6k6k1fMcOxpvgxVe4g71LOg/uxfW12v+TDA+Ot5
rC0qSAWHwgUN39L9bHtGV4gAuqCuNCIWQuZGU/kZNTjQ3h5b3CqZu15Ys2ApIvv9
mCpPO/ZVLI867nzuvmi9EpTgGdhka/yavmYGRtU1xOuQ4L1vb0HyEy6dT7wu/FXE
ZRoznLMai5T9EiDXD8d1Y2p0iElztM6Ewx2+Fy4wBQsPjhFCg4S9XKky7ODxvPSk
ePSC5tF35dU5eS4dUdQuG62CNdvmf20QXJ2MruWqwgN0pTfH5uz8GWu811OjqCLI
wT+YNt77RApP265hDrDaSrkzyLL4YhsyzTLNBbFz/pqMh1D5dp2bDMJxHqFrZnQk
2za6eYzxK4KpXU9bEt6iVqHZZbUXk6H838SPwUqrnXru+ccFcKJf/VWn6YxIh772
hGG62l7CVCF6EkQdtmpHlxFu18Pnb4sSRX3JgNd/sBKQNewRdO3LWTLVFXIzmEQ/
YU4yeSuAJ9Wnq3EWtp78PFwsMg908OL3Dl3li6Z9d6UBy+/ObUnKdJD9KGg4/FHB
tp/ULzNErDpcY4hridXfRjNaof3FDrNdsNURaa2YT7aMLjpWgKIHl2gG3eI8oMtw
TNa+ka+Zx/4Gy2/Wx2xnPFVZa0hQFgIpfenCcKKHF9KQpm0FPG10cfiT7g1Ok9fn
rpjp1mIdtUtik0G9M2mIVOG3WUJ+tUsKiCN+IEabBDSXebc/jGSLiGTikzyfO69T
kNekPhr+kVAHkh7b/aphu30AZSfGHaHALla08qksPvXGNfnUT3615sroJrH6injD
W6qGh9mVIfDmAqG7IZ1Zy26wJ+ZERWhlNno7BokQtU+5lPRPqtyIf5L3jADq7GJT
2bHgIfbTu86A2z06mAEA+OwBQZKbYJ33yQyWAwSVW3PEc2tDnY0xZbrXVhyaCF6I
aL4BMZAUt2jzMTkPuW1Sy45R8GrVePUKLzIeGVYfqlcntd8VVMzbOijJojEAlK5Z
bdaBE/bBSiW/ZqkViMsUMA4OuCNqHx0NL+rWbAlKEhVJ/aKWl6LDh/jRFK46qnin
OrfKpu7QmH75JjLJsFn4pXiFXPApILfUYtGfSDdMBKFn9TVnYTgjwzJi8Uoa/7DR
crYE7r+i36k4uNlhF++I1dUG+owo8gWbmD6lnyxF98wvrNf5Ptadnlwm9hu/R/H/
z+M9hNIkI2VJNGtDDMGae9CMCvE/HumUKHAuEOcw1yK+wkEvPFQgrSXVND16qfE6
pG0RjDQpdr2KzCqFk1uBwj0KmK/Pbrs9LE9/0O31HU6Wux3TnJjXB3rUpncjDC4l
u5ZpDx+REA5ySpSCga1QEiV3ypqtPD2SXL67dpIhKC+QZVJ2hnxOUd1r0ekHZ8li
278rjis2bH3MLj+IArJLe2Nfxa88IZ862X1JU24WVex75JNGL9gcFuWZ+aDJ+hPB
J4RTCDIjt/pNNlUqSibPxzS0LZaU6h2sTgB4FXTjs+dmk8lXeaVnIEDgSIzQRJhs
X3UUYlFNj9I88SW4gh/HiEsrTofvq3Q+ZREPLQrry+UVOS8pvj7VdVEV+dUZg7NJ
16mMaJynPTQe37qKmpP7hCtvjfa80c1m0Z5wvjTWWewLM0QOq2s532bEPZMslQxT
L1QlfsTTkvGzxHsPNrlNZ814lUYCdVK9TbT19fLYdhdWSFr2+mBgA4Vh777tY5zE
wW6nfrjl7BoJanWAciXscdKjOJpXxRBGwPtRkMDAQywfwYB/qDuO7YFiTbweSyAx
aWEf9NlANcRHlm4l6N1//eM4FVSME26/5eKWYmDxC6eILMjC5W+kL4avpd6dN6Sw
/RuycvgMbRpQjMGu3SGN//DHgN/tMzFZUrdVMxcc5XEUHTkIjFOGeTPSBRrwfcTo
p+1FahM6KndItZjG1q4e7Oh6+48mYltNV+omI/rZTw0IOlFHHPhbsVakrWUWLZn7
t+dNUrsH8TgPj+xJFdBLVQXErvmb/Tw5eW1p0q3+aDRNC1pILMGZuRF/x9FCOp5H
8v7X3H4DeGW+9B0JGEN0Swi5Whig5LisyuypWP+lQ9VWAzuKV7nsC6afvdByP7Zf
B467/ORGlGdl2ai/2vJgxGRi2eRcVN92LnlvjAIWG5ceg7SA8H0tAFZ+uyll55rz
nXdL4qzmK0kJkVRa7z+J/1QcAW9alAinL/tZInLnrIhsmOONVIIDNfBaxaXUnLzl
A8vOMgUMs837y533M4E/s6Hz06aCrNj5G2LsE2GzX9NVoFRScgfOsxX+yiHmERRD
9+sy65jblpuNGnc907Cwe8WmR6wF/KwLxScpu/ch58PwO6+kYS/+3sFvyRMYQ8rh
ylKmMPEmMb7A7dTbwh23WnuI2h3nTMNd5+dhMCEaj0zB22U0zIQPM5wmJkQXPoC6
n4KlTC3EetpZ/PzB7f0YIXmB5VyPcOrvjSmqQe2tTBNmC+e6E/nFA0keycQOjV0p
lK/y3esLXqrjlH+DMuR585dDJBETOtZ3H+DaqQEeT8PmMN0nQKwh80FPg07NyhZP
kmvJTczQdOVfxDDyqtIHowl/NhzCtD8psuC4oN8J8y8+GmedpSfrmpHEw84kyVUL
TlkO2eZ6dnXxkLufL/XS5oyNhfEUF2yAcqx9pFPAb5/5W784oUL2KpKcNq+lfetc
DANLy2b2wv6/Hjand6U4C3FIj2EWn8Y8hB+5C2v06RUm9yRHQBQksOsL7QEuTaNL
ZmFDh+7lEx9KQZLddAxVZSUSXcCPnanhicaNwtt3INhJ4WOSyyBW+I2pw+KbWjB3
+XRtiSS4CCPiE+JIE3PjIkXKoE0EFoIcGEVIWknP2tsiH446Ad1nRmxIng01u4dd
ed5DM/pvviwRgi1gaC02Roz0pvKLyo0m1ZvdZnENWOXzdtX8Hgc2L4QDgVYIQORg
aJoIparm0BynzZC2ctDDPgA8teqJY9Lm3+2ff8Bl9BnryC14H165KrdEu/oefECG
d50R+kFAzA0+aGwHd7pI3KLSDWpp5j266Tmtcktkfnm4QPdwwHrh6EUYzWYuypyx
qsJTFp3vSnzmVkC3lsixp0MPJHAJYN65u9GEiKUochyj3oFehSlMMh0SLHl2qnDL
4a0cO5MQVzsjuadOJuR6WPgJ98yjdvxPYuKjF9YHpecTZPDyZFKSh2g7mDtyVcqn
RiekT4ypoOlha1YjlQHKnGjy/vG28uIHSlUBhMPk5QgpJrEQWHDSTBZYF1BFXy4t
HP/mfyB2gkrz+aixpAdCXai1wZcoXJJkznNbUM6FQ7YYawuQmBRP6KTkyjvZ4gv/
Oatus3p+bO9T+RPOJhAKmCGy/Gl0+uhRkExuA2pq54eV0KTOkb9UBkRxvdstIAMb
BocbMzj3jdlh8Bu4cURtOKfuMwGZNbJ+/yHoxaL4WIhyAZHC6FD2scqzjAOUq8R4
ljqWbaa6Sa4Z9rb+3tgih9BN3KoqRgk4K5Q0x1hi5h3+kuHSgxnKNPakx5A2jfb+
oHJI+utVzniyG82iXzAN65SNweI7w/DpQ4gsYO8hKCHW4Ce8avqfYhWZUXUR2mHf
PJvlgashgopOBy9zopqL1h1hpCfS3d9KUuwnrLPYrhGWx7Gul0b2jLGOo90YwT9S
hjekmpm+Q8lub/QL90fkydcyhDmKQK+cjqEcshwJnHxq7B8aOaERT1sFJRZrj0VL
UMW62CjueatnnWSxOb58oFBFillXnmgT+GXvC436XLzmeZEnLRkQ6mDKYE0NfezD
th//Atr54efH2S56Bf4AtV6tqgNzMIvMuj66IWCFa38lLPPuupZ2kSy7oRlFrzLX
iN/gCV7NV/Q8lx6EHivY4AnnoSZsH4bfiz0Oi185FuF3YjaUVAsUPT3MH8cp7Yyy
uhxYSnF14p2io2xYbMWskTX3NDMVdAyplNvzUnOa5PrBvjqGdiURP9DNlfdkpHMg
QjG1ApP1yOW81l+tD8KXBdjLD/q3Gh1BvjpGsjOn2aNcBatPuOvIUlpGwEoI6pEx
u3PXtOjaDyxML5a5HvEAQJCl+z4TsyfZYH+yE+/qEaJ4nSi8pIOOPIV/TQk8ntZV
vyE5RMhaXjEYY0l9Yww0rv+LeooPQxMwvlTCmgImYNq2qM2VV4s02AMKZsByC7hD
S/fh799Iw7unvwLpxpcXwkHA4m6+ACwgtYZe4NyZZj00Sookm5l60UbUyPaaoi8z
a6AdkXRw2cTu58Law6Wk8xFRMT2DpEuI4H4wIzsVQHplEbNLG32LUXhQb2GMBDiI
NgD7Aky3pN4zcX0UxMeYih37AXMNAxwT9C9ZqnMCsYLsaNnr4gNwl6IqldB/9xfJ
OdegwbXw7PvxXmrwtbE+roby0oWGwne8jM5PuD13dK/CWqrab8wc6U48h8aIkqED
pvEQzeVBKwfVXfFrl6aIjDdMGP/PmZn4p/t1RWfP6dHuFi5LVXNu+Asy9/8GHXKi
t09GG5f/m04TBEropki/K9pkiIMEDImCI1aT9+Etowh9h/U2DY/fcV3D2enYAOtN
U66Owk0Eu5410/leQuGq9zdIkqj7m9PrqxISK2uE98XFn3EzCtEZFlbY1242J09F
EWWXf5dv6K2c9rz9r2epGZNdikSPUiasnQcZ2AcXjZotXORKi2k+lVCYe5p5Uv83
pClirYX/h2RMbeobdshezh4A077+xTJlPvXCrC0s7/pBacoAvHt8gk3fKwVS86Lo
z0jEMJF1GBKKjNufyioMDeYolyFbYYkSjkjRaB6HrHkN5wGMkZ1IlXKQuvndVBwf
dvL3e/PjHSHqMDdsrjD1AEehlUNmw8+h2LlGJ0aBocIqefSJuqWcLEADb63y+Fue
3TxpbzQUCOGmU3l21mf/inYjfsNcia7P1GGALwkngo2OOuyaTzM4634E6waod6zO
kw53kiCgGR+2yfF60qvmtl8dF3MUq2xZOxIbYANPp5bUv+3K9UtrJGxZRgLaBjUl
e4vleMURAr66dxrJifjuTgleg0t5zx/7Eb+RraxZC7jevxNuSLGfqfVUqkLbu0eq
0N7ofZpbzhhh5o2VT8RzaRYjW7r6cuv/VcwH6Y3cPnb9J6BZzJI1ugekr6GQHH05
AkMGS2uMOG/WYVNJA+0pfYo1TXuPtdgbk3i+JRHnrncs9Qc5d0L0d9Swq97amLmN
24xXpdrsVZf7xZhw3QHkve/ygQ37X6f440Ir48hxGmTA7SGoBTIQs9vrZcPzFs+n
u7HneNn23SPGezrY8g0l9b6ChyaYvqdkTsmUODG7QOcdu2DT4abfNDfpghVNWptz
jziXgckscoEUJE7fkTbMjfBCkBUt/XG0ju6VjfpPfNAcHYijT9XXtX3reaJAQZxf
nLcCK5mq8fxrcOEc+83hzb25x3cBFq3q2DP3kQRsUaj2AqdA8ShVGjdMtxrKWNBp
r9SZdSqCV3QoDT3vdUqoCDzgPeRUQXjw7boK5cRCKvZ/vUw/tRLA+MtKBxbauDbd
P+Wb6i6PQGQPWLqtj3VrKCc9zSgkpz1NS/jBiE/uXB22tUvr7wE1RluUjfT/7er5
O1dUTOD5GYViWSvlIY75xDZZf6nNWrMKb7ERUy1o3afvFz78b647szbUj7DzOoox
BJ22TWl3JJafE/8NGX/v1NMWjLHUk/mHx7XVTKIwXkseJtgKFTuh3qnhePE8DI3h
6UcQxj6tieUbOT9KuHkL1Xp8RC6iszzeDMCDySMhKmAcIKuurn+12NI9NMMC2lXg
108gVkXjeIUF3w0+TJQ1rQHbHs+J4vgPu1QXczWSeKUbDTwAYomhgUn/KVbv6DZZ
jOVodGEWH5SZVkIieDy89rWwPIp3GCrpQ2/l4KGXJXOcWMM4+/wQqt3ZnI547smG
9DLcKct7MP+QX1/7MwbUd9rIqiVDT1u+e43kvtkdzvMMlleBnuHdLzsfQLZtdNPa
bJo8gHgOhDDCN81i4WYnHBn6nIxlvxatiOlXAcP32neKucvl27WUALAdPYSJHALW
SOrF/mDCiHyHufvJ9qMm5Uj1XVlZSbpq6huzJ0Ht86G9lyPZS4i4S4RZB57kWP32
7eFms/YhBQ4pJjYdBz/b1KMrL4kbB8Y1/giAfDdh4DsGvO8BgDwYzAuylbT5lr2Y
0Bkt/DNunasSC1UZvTSJL9V/7vuflZCP4GB57H3PdOCiko3UzE/l94K1c1GZU//U
4EKFUQJm1hCnO74zDA5ulRkrDyyGpGxJ9UvNbblBaiKBAhtqfx/tkJYKYSjO7Gwt
jNKOrn4JGFNNdn5sbLz8ysKeoY/TlGgIes3LefqQMq1YOEjoh3w+f2y9CC8dSPFi
A8WdgW8sqhdF6lQtOrXl/ig9d8zGWmx5DXP9eMahariP8Qu2Jc2TcwaGuShqCkTi
MBd+87GGgBeEVE4dnre+cpTjmAaGL0wZqv49RFqvmD6AbtHx2gHY751kto9j563q
+NOjmnN/EGG9Q7aZ+e9Z2VmRXV4KsRpFbX+wOdPLb57R3/O7FySR9LPcjrH1NOwH
541i4mLKsMaq5Tnm2C9bgJw9DDei3qfvlcCzrfXcWNRsaEpPJ2jm8YQOEUVcUKpk
R5kKQ+WKwWqQHSpxNuoh9KLZtdjt/YK69chXQNIDLcgIk5lzuhn5sP00TV3cTugs
4vYIi0siSD9rwGiM1GqEY9tu1YUtC4ZuQQc9TWHhkBq9r3DX9kRaCFm/SVJrYoCE
olHSB9A1hPCXCzAAkoQpVHppdpMcuTbGsjlryj29Ra4g830emK2CZ8snnNGbEhjb
rLCUWJKmGjA2oN+bkiYH7dy1ogfmi6s0Yh4Qc2W48hz2b4TzAnKi/nN4j0V7MLrZ
IZY00qApG8SgWiW3b/lRckp7VXcTLL0EYu8HQEOfuBbzKSE6fA+8YNx7bZyV77F0
6uhJgUFs0aeVTzwhq0ORIOAFPYtQCWhw5wn6K9ynz9n14gRZtLj8vWK5RmZSz6O+
3R446Xvx/N16/osuT1xwHKuQXG0xYdpwaIbUMu/s18C2EfpkI6trPyUeC10mSKIr
w+iMvYnorsQBsHORxOoBDDkEsDplGN79eOZBzWwrBwDpEh0TrOzR5TrUZoFxU07y
vHga6pdVHRfdgq+2D0GTzhWBA9khNo+vtfcDSt8nUKNaoCUz6PEZfBHQSKqeX+Pl
5AJzdGgFVYH4v47DfwcXFwIBlXRad0d5tb06B+zfXoDvQJnNrq/g06Cs48Cfp64O
I9iWe7oyqklcnflLNoO+hicWvhgQPXSdo2Wq30V5NvWFujmcg9gxz7sdrc6A7jbS
KhiW61q+iAlqFW52rIOyozy5rytPDdZW4FG/zQAawHviVoVesM/JPMo3o5Imu3a8
v8mp0D/5WHF52CcBWhm7WSDxvMOrb7jS2ZZVVienRfkypcM4T1z5gphELvCS2L+x
wtI6qz6uk9JQUT6wKYqa6IRFb3zWO9RmoHYrdlkylo5LBfM7w8yoZ3Kv2hCpTpjd
2+f3k/Cc6+QHMsQ48TCfeh4Kucu2g7eyp9BvEA+GBRmwzqY4TQ7J2W11CC0cne74
A60MrFe1ui1QgtNTiVG+Bma7pflzCI8ixZGIEFpscIl6Kx3rt2ZAhql46Rgsv63z
Ghep63/zG3njRSq40llY10bks5REwElYHghIH7Z9s0IIaNwxqoSTIyWsfmA4TcT5
6s4oeQjKeintM89yWZs1tThfsRDB3UQwr8pWio5oygl2tRl7PDeGaimXVlTCSlHK
g7uOqaSp2kYRpkB33pRJrZHJxHz21pTzoo9hP0P+RaZIZu3owZQFykebmwLBsH3a
k7Cd0piaQia+dJNJL5fDIwTqo0rrL3UVhxSfMTTfXLKxfzPtyWdseGaUnS3falHB
Sb1mnvCiUoPJr7JXyfSTU7O/JciFQDhrWP+rnUH6ZWECeiy6PERLR+nLlEztbb5x
PP2zuJ2XV6e7jbuZbxuDI6m7kIaaJjyp+aQwbitA10uiyev+XsBG36XZuhNv1gwW
JARixJsReULLW/y4JC0Led4spyU8bCmilucNYDgFcTF672pJqAwR0KyvJya0f8qQ
Nwjw2o4U9OoSM4MYT36VqeYFhZ5u2W+TN01XptNVaLbygRNqT2NkBCiSU2hR1sSk
Nz4yhLoMwVtn3qbFV6CAnpEwRSnerg/yIb/RVSNtKt76Izr6xrcdkIUVKDePY97u
h5K+L4mYPFejMuaGWXW8ArLv5KT1ysiYs/OI2prD1CoDTn76esmnrTzNLKa8vprz
Vy2kWLq0vFcQ8l30pn4r2L0xvDMThX7J4UxsJt75FhrcAOuiv1YVcUICAPZfT4SN
wDW6x5d7v3sErwCStjvop1QsExNtdrC+vEhgtz5AepMiIEaTXogezuny4TH5jXOr
iH3eUFgJxkdNNTDn3eC58n5MwSX90j3DfbmF8XdVZZzBMqUr7+3Qi8Qf5z4Z5qQq
gS3ZAjsFmp/vlVsMgDZJg3UaeTnrnm2D6aeNsGm3/DhdgkZp8w0dEc4DrAKUsAyu
9IRy6AfLqJCJeV6QucsavaO2TVCgVfT0ftkqRaNfi5wj0oQK0FesPOc6QzDe+7tX
wRF+5xxBUTj3jVztNjSQ+o19pmxPUJL9ptxPxgRK9r1wZ+6mGAu1/N+jWYuFys0j
UrTn1a/J5aTw8bMmOUs57Hau9oBX3QiJ+I9GkSgs+iLo+0s/x65QStO+4lDCb2Pa
rf5zjclnAvFTx9pb2yFNHmtWKpFf4UuZvL+QrF2CqAVs14CUg61EG+CzTeXDBLj5
mOHrl/RpWd7REL7MPONP+q8yLUKzvBnmZZgZKGY8YEsDA5xvdxaP2cXf++XmPHgi
dk64Gn0KJuinX1EBkW3K1BT+LwAxXxztismoPLFbbxiy13iynRVUIxvmssJOmFSm
3DaMwUGaKRqSKxUf/dV7BJejnymHEj4b4pZQcuCHX8yAcBGBQnOKkAvjnOjY6pRY
kzDAFNsEiSVJehKShS0XDbbP/UNBIrLYWUcDimtdOA3zNhCo/osqVuheY6UlwaN1
0wy2MiOPtg6qCHq7F48Mq6Xjwovfk001QKFFxFw3dBPjU92X7D3/EhMWoc+26Ms1
dSBD75F4r2jY3Q233UnwLtkvYp+0Ez4Lv7zbfCEQj6H/3L+IbQTRuCMmVhwlh4fb
J2jpDI+WmwG5M93wsEvxs7oPv6HA/KkN24wTa1ZOTqMNahNicEpqnf5etCbFH6KV
N1C0xtxDMj59jPxbD++61L6NaRqPZ40qihdHacv82eCBfGDHzS1HbAzrY1Hm4tRg
K8xjxhbat21nKuXYsi//rf6J7QGEji/uUmpaYL/FaIemEDR/0PicFPQdEKembIMv
K3hzhyZro7Am/uvafreG5j7+6bJTXEtshAifkJL8xFNPAHC3ROKcwSgnrh1EcLtA
yVW0K7SxQbeM0/+0+4ki+07If9AKEke+y8DHOzXLnC+bELsGZr+CJUnU7dRLqkfe
nLAhPgbfvBhb4D7KRntITozTrnIPu9R12lpk6+nCanTKItE3wUic8AUBvu7kQcsl
Ro0vi3LAvtA6vgeT6SOWUQGfcxmxsXiKt9vaSldpBTUOXdDsAoiJ2NbtiFNXN4i0
IsVizDSsrAvvxdAA4z7U43pOp0IynIvZJ6MOs2sQoJC4KYhE0ul9whxH3z9sO+63
4kWwGhQZbVDSELJACmRTsQOPO1JyIyKosUzoizmjgYXG9HcxB5+lY6EYEQHO6vni
7vbXp+ukCf+TIgT5OTk4Rf9emxqgi64Ago8lfMuvnmD3K3Ysmyp75vy+GFtcf7nf
ANR0wjoT3bcWh0TYg9GqJcDxHrWqSJjbMM83D56VmPXrxoMCT5AaArTomLAuknGT
s7gINbi92BF0TdB/6TrFe9T38K6tqKFuzgYPgqZIw3SHiKCi9omeTLz3qc77XKDm
5PXEDsi1K87YDq04BRAUaoxa7WvpgrcxnIdH2YJaQKZ+YF5hJCsUhYSzMNDE7zyT
4YaLrTqImMxYRWSP3kTX6Fqy7cu+jZ/piDK+wLcTXYuRB6R6QJH1hWRL0AbmTDnc
uM6vCEN2tbUU/r0KVIoqbi71p0JHu2VnPgx+Za5MTcCgvclcAKMn8bQ65K0bh6Zf
clRzy32ZNL1eKKQS3MWUwo+1An1SeixRi2RbZ7buHKg88iI4cgf1rhOQL62ILyBq
AZBtUH9LQGKdacnSHuR5e7Xokx4a2TMbysn9Afdh7hrgVi2RSJe8tUthvBLLA76x
DGaJuugWvVOeYtPpt4lx87/SomwkDxkKf+CBbS4sUfP5SoMNoU/k9ZagpueQ0jm5
WmiDoxuxJru4iz0gAJ4g0Rec9jLz+32c+3wcD6LuOwiPh/luIfwKp1yOKgmIE95F
bTneOkCggx/pFnMWBAiIffkieiGR4g5L6wJ698mXZgcZyWgmFqYSQY8tVR1aQNFI
3gHDq+VLfp8vx8sjUnXwANhrqbpcL588yK0V5Ynq86LlwpCfj04/GPPKqR34z516
bM16+Dv318kGky1IJ3RnmIRc+fjY7rAnzZFhNNJgS2q8/vfO+PSNutYJNnm0mPZc
PEForzAUOxxMIW034F7FOYeDQ8mYvAjGCztvFYUXSz5ZvWoCt/JWgOWtf3pHIYr5
FsqBbAqZCbe9tciicT94fpK9IHnuq5UJB6kFDh4Qx5hYZ0yJ5NkzF5vWOhCxbpCn
WsycFeFD+vGidiv/B2Wn9YEDjR8iW6qO/mLDJaA0hXqllpjoMf4xDA0+RES2qfsr
13WWf+VDoHRZezgg4FWT4UnHOmiHdSx7OqWLLu5OdQ2YceGM3bDCW9H/o4tf8Ins
ynrvBVCliRIXR5q7xuSXe0OQR+XU6dwtVzZN/DsqdpMyZg8WzAxui/GIDI7Swp4u
XFpzcGEc5BzGpxwhgAcsk/0Av9C1Me4pYqtNyn7lhmS/6PgMXhhKeRCT7QXQ9eUZ
IfUk6z8KoGSK4kZrH8+b3ewT7mNNC5hQ9KZB65+GiKav2fm6MEJDow86HygVyME0
kkPONfLiS9ZSXVdIoVMDqIhPMfDpAUWdqt/uNZmBnnBDHROjMByB5hYnF1JYj9Wd
wfpIaESSniYTpkjBHJnEQJ5pMZNWdQjJZ1S4EsJcfKclUEw5nMFsDPYY+wrCuMGh
VpHNc8b9kVTGcFq+d8mQKMH2aJVaRp5XOWbH6L4VAXU454jw2aAzy2ZHvdmLlYsE
iW+fO9NSG3hA9KF+LwMVGFMZ1oAXd5x1uDkYAEAgDN7myG5cGZ9icHk5MISAvJ45
vROr/WCX/NKwrPxuTiIsTIaqZQVeBXmv29Ttxz+rtkowX70SfQ91q7bw1ZG8Elpm
2HF582sfFCY/0pNfzQBN5grqVlOvnLVH6TUaE8HemOTiIu/NM4QH8P7IZBKuHolX
I9EpizFDt5r7RbyyAqhIZFYYtetl3SKVtlbS17P6uiRJtbQsGqoyOjMKX6MaCGq6
iL0j6cV9s01Bppk0XkgeNRLasY3jEGQDKsZfc29N80yJRWoqDOHRPOCPmxCI5kEK
ylD7HZRDqDOTfVI3QCs3egnm/7S73bHn9r3OzEWHAPILnDn9YovpA5g7aHJZETFu
8VUPbS3WlRJ0rxB1dGXKT6oRJBAT2jaYHnfSw7gA6pBlqETvDf3kCOvIwitJyM9s
bM4wSNsM9ZTAiYNSJW1MydweFScit3D0b0C4js9dvZx+5BYlL3GxkCnLfjAhbkNr
tyKfCVxI9CE1eQ4dYOg5Eh5bBN5ohYz4GnPr96Qr80h3Xi1eQYSnpYzl8F0CSvyK
9tq43aWJmkA6bSNaZxZtHmn8lQgVrqpSXD5/Zq7/JmBHlIhKvdL36QTdJVPO2O5H
dPXlJQr4y/B66Y7o0ldYvsiTavPWu9dmGF0qdmKknmq4IrhUW8yQGds847tuK/eS
p6tzVt8m74F3NGD76eJDIPF83TV+INQbNpN7CzH/vm7G55AzXMdmI7Acjf/wR3fy
gRjgT8V411LFkuud9sd50aeDnShf0JZubHv/tJAoF4Ol8T1SoafqoX0jbPODWT+B
HUQxKDyWupi2eMRqCg1SA2GFNDfFPQ9iXGYMbQncAKbjgWpmrheK5ALWsq//fN2s
zTSuuYMKBjB4EmPD0EmqenAgQM24cygtKRXWFuhwnMjmxzQIt/ohurS+ab85lmeH
iMIzJWhaIZ/KSK5sR1zK2bz1VCQ8vl6lV++5HAllMv1n3FhngedJzzy+f7ep/MVb
9c7gzBfV52SPbKVFbPsuQgPa8Yh6x4f/KNSKVBqLQgNr+zXBBGtIpXP7iGEt2Wog
aj3cq5oE1NzwsXAm0LDoucBJvwvC9rb+ENS0ZIWW4So3cUp1VRso9m5iTurg2ug0
Oa0hwixk3WubFCvlB4wZ3qak8q7uBo7H8eUA2NOFxK40XxOaU/I2j36KVMKT/GIx
TGjc2nv8/ICOLIpim/yE6VK5wOBmpscxTzrkAShNSlnNGdWuQASwveKYFRt8SrVs
xiHv/Gs4tjI5yj/G2px7TPFMm8c4AZwA7M0L6FBa4ryfSCzLX/XI/1POBhHx7IEG
eLK4pUquuMGbWF009AB9u3cCebW7PQVlP3Q+W7NbOQAX205sSKj1PUSO67wP81Qs
vDVnen2ftceaHIo2GRugaRMk+olvn5/N//lZKadW0BGK1091W6c9wqH4S3fwNjLU
PvkzbSa2GXDfWLtl3SYEZVSIhQI0J8CxCjG+VcMgvUx7oH0XoifRBrfyUgcXn2sq
fFKEWDdTo89BUscKBowywmRE2QXxbLFFxPY0tMSytopIIqe41xDGho8wO3TMGL1K
h2Aens4fAOmatQPjZEia4oZoWFxBtWemMTbbqy7R6h9uU2xVHsqMe27BX3szK7wi
09aA7FKAwOjBu4v/YZb6SL55XoOwYHZLI0aUXR3KqsQFIlljFc38y7Uu6vDVZEn7
JJrfOF0Vyr9a3p/7CSZTtkG4tSR77qJD5hCCFcoVdZTpbG7haXevWE0uJkm5mDm+
Sp0W0I/09CwBP8v6Y/QPsw4zpNFRiOQhvNgLxdjZJkTQh6at6UIeOzh91QGjhxj9
16kmtCvrDWsFfxLd0qkW4t/FtBD87271eBWE22hHGX2L00PdZqXohyTW//Tp4EZq
g/eXdWrXtDW5zctcx47GRbzmA2nqbESqERmOcomfMg9TotqYoG7mNdQ31Esru8Qc
kdkYoduHRBZ1kgDmV26fMA8uoPVMILK06vI2CTvarU6iPik7Zd6iJ61bq31JyYjP
aEofO9clodts4KZ2xWs8MsEHAfWw6oDjyT3Q0s8/U+7eeHiEhIGIjdgwNLhamJwj
nadUx0i2rZ+peOJDHoip02SivzQcaV76dDrC6KnRA6gaBLpjzkwuCuoMw/qEKCx+
1rxOu8eMhlwjQIA0cf13+BUoH2shl/ASSmIy6bbqCCP2vzlsaz89DsLNiQ9kIuj4
v1WrrpLjIofP8B01Sp2O01qXHvwy3gZ+aDfL7bJ+vb1eu2ZeQgGiAWBXMVCHRIk7
SRxBnCfGM4dQxj4A6xwy76JEPCBalwJ1Us6Vvvtfx2mJYRdOnXGVUNBT0LmmDSSO
lt7ntwXbZgAVCfUpkXC7zePGKZ2cYN4zJREZ2f4b8lFSdXVKaVFghiK0EY7fLlFA
QolDi6YNRzOnxorLpLf/irb3PDCbeIPO/6O6hUoxi2Uclx0ptaYShWpfJXptqrrn
wJBbK9wm7KZ+qLiwjqM9h4Uf3U7NXtX6hyF+EqyJvG/jWKhGP+FVwOrorVSWKAaO
IZS2EHDjqVIyANXDNk8f/dKUxDfZHs/kdmRZVBKxjs8EdBvJAIRLUhiDxBuTcQXF
Vkuf9+VdKE/c2QGbioPwJ0jMZKGuKDh+g0I6SO1rnNgeyfWf+K6rTQ++uKsNWPe0
GgIzEysMV2lx9Ba0kMxZoQ2jZC6rJFLN4VWTo2ZC15v5kp85mEOzhDZswVK0wLCM
`protect END_PROTECTED
