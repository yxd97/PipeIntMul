`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/lit382xentvEMs/n4VzX689B7gHsAA7Vvgj3Ck040QvU9nV5uHz7Z9nxGeAerV
C7QCD9CL0pNvRwoOeHkbdoJYzfvqjsVm+vq1kWTMwR4V9XpT0DHTeXRH0mR0EUjA
5W1AVuj8xSHTIvtPh/bgli6J/uxhba7f1t2F78VcE4sVuAJabRLsND1rL1moseRX
tnoThcbFQiZ/BAQqcwsaEQ7MwazVZc8qFPLFIbZf0QabKGQvfluZlTVqOXpjAr1O
S/z40Yfb8654ompAPYpd7HiXaEqEreVO4utjk2HufqfYrJwoHYOOGp6suT+VUFmI
CaPujwBKNUp+yrGvkAg2Sttxw+b9y1dTYbZcKTJ4iflqCReT0tNlIuJtDsl3ZSzp
SAomcotsB9Ys8EwQ8udn7sQ0GB28ZINFgVNYI2PB/c5hYxlBgSDbV68ktgqdLs10
`protect END_PROTECTED
