`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6u3vtbxL/ek6NgPM3YVQzT+e8gt/5SsCgz9ZPORF0PjIUbyYo4qoHK3ZLXjI8ZWa
ZDKfGq9O9iuYc154B+6hjZKUUA5UMODtqWz1q+ErRZAx2YPMJ9LrHzl+GiQomSwL
xlZ0v4Lsz/ApIgmArWpyfxBunE0Nr1aaTQctClI/uK0Jt8jWK1VKg9SyoQ3eZx3z
4eK9/R3rQfOPCMOlagU1FVXVJGTsjRjcCzUZPNHfM72Ccm/RKlSpeogf+Jyn/01p
XpFxHbhlbWaMn07NwTjy91SNBzJEhgf6zNi++5tA2VFV6GSYsDB9Yz3/gqlhsP1x
6SmVPVS30GriES661NWs57nVGpdrRPFsoFf1EKk+TboK1jVOMbc6wkDskntskQAf
HiHeGNEqMuUmrZZzk7LJIp47bp4APibKwnkKlMOG44NYGTot07xhgZvdVx8wErHq
QuKQxPOh1IZH7cY4iCr00b2sZRRUX6VWzGqeJnKW1wX8/llBDVG5zCY+LPcRA5sB
VgNUVQu8u5XZLOLrLUF1qhYt1PxaPLK+tWqHh2ITYko=
`protect END_PROTECTED
