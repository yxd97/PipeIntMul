`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Usz2je+c348ESuQuV/sAEo81VIdRs9LNWI/Vb4VtRPqTqlf7xowz7T+TFoUbaf94
kpAxgP9PRr3vAPTOQQBIqN94wJxDdCAbhiJnThM85klADPLX37jc750sVh3EWtfs
a2PMlbQiFC/mxhphxaPObHiSBfUmHZBsGX/L8oyVZxETsHY4OOKMIjl1Ei5Sz0yd
VHpDdY9hMQB0mwgJl0kt+KD/JlZ5O5bXF9gA9ju7QAtmdaUdQHdapb8nJ3pcG2c1
Dr64ErmBIX+f7kdiW90kqlDH7lqM96lYnzXQeDv/H8GP4EA65828Jjd5Z0CzOlwy
SSxMSMRxDGSNtK9hCkSs/k6IOBzC/m1Z3yyERkY78rU=
`protect END_PROTECTED
