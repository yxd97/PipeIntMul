`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AE3vpRkAEER8Pv2++3eVuWmnVDkYg5jbSzRKneUEW2VHl9fC67/pgSRmVSRhJ+EE
pVJaDqFDqfrzIxPbuIhZtge5F2AQOMorpC0UKmNinr617912Q7ZBqxJsJxw3XkU1
X9KIbaKwKq1iRsh7gwbbDVgYb8xImGwc876GUwhRezcHR6ySNS/f2dGuKJtYXowU
vhSxnnQvn6Pb+UOqjpi6MeMC5rvU8RiO/Sl+eGhgDKhG3wE8z/rvd82xFzrzgOhv
UZ1oLIGrP3oYzwZMeFmy/CXvejGaz7/P+PhzDOPuuIN+NSYgCttU3XlN6zjoUF/l
4zXsAJvbeBgxV6lh9VMQTNZbSg91rZkBup2oGKxQkJRKP8h+0SFtKtoc8hvEiyHt
9Jc0FmP+7HiFHkJo5BqauaWJDLsfoNVfqOoa0f570HmOEOuKukno3Ggz0xCtbguB
9KbQ3ftd+h64ze4AjqBrQExNAQX1AHNSNF5n4FRM4/DgQDyWwPS/mv7W/Zh7YPUE
4XZ61ExQojj3usWamZ06ImooBZGcbO0YJ/6DcH0oJ25a3E1zb4eIQ9ccvcjURXZH
mMPxy8/yqEmoeqJQ/7VIB8QHZS96j2geMG7o7lc6RGuldC5duNRsVa0+2GaKyyDX
+y+SGVvwttaqFMF9lEof7z+6M9E2bPA7kxcrXjUyLxz631nkQszfFDuOFVJLEQ/H
IqNU0CpOaIzE0E/0hmPrOdicoMbs6VbXhyaU/XSVXWWo4pJ91cNK6cTk7lhhGA7P
HkNjfquGU4ohDHxZZAOeUxVttVM9YHxEkIvhzkyjbF0/OzE4digW7HrjxH7r/39K
KLM8TU4q7ce1I/xYdepEoca+zhmL7pnTs4+hsm/Aoen6h9qAnCrnw3CNpXqC1w7p
hxcQt/cl9N5qufEQ/eAcC/h8U7HZxB6RVYN3toqbndsec3euM62405Q7FSSeNMdF
nYQtmT6F6eE/qpVV1M0uyf3RtS5EIB9yO3ER8Dco8WGMycGHGS5FaF7oGtoMUk8a
HVZJ3LKOgocHUxztbm2TA/P65M3g3KVM+FNhVDpyQqJI6SRena1ZaidAI/A8lzfu
7fJvFuJVUugeuHHERxb5NpGWLU8VOXKdWj0Yz5PTJO9lqz9j+Hi+mLqoS25kj5Oi
tAbCT6iYxYknokI4sFnT+UM1oR1tRS/98Vrj402+zyA6UVC5EH32XJQSXIO1UHHe
Ffb7y1EVRxu9GbxBCuYYyL04z1EiIPXFqDzy3BJOxn1PUFWsRorSsNAePyr/S5Nr
16Zznx4HXygzbA7XvJP6NQq/1Tn/XaR54tczULMt0ElJNn7kC2F4+05UT8GAz0FE
LjQhtkU6IF0n3fZ8m8FvauvNdhFF+Zdj6lw+bEV0cr9RTH+/MUM4NuXZS+ZmUsER
lr+89SdSs2PXiV6FzEkoMkuubUZkEnyEhb7Q6AJK6ym3vmIb8AYSEmKXUmDyaiBc
i4OMUv7CTb05ey+z5xWB539dFNFzzEoeFE7gxHN2mnaGiqgDW8aXAZVFz1YhjymM
zxtHYQ2nQiBDz2kOfSCBx84wq8bRsa2WKMn09TAvs1rxyV6u1z2WpTquRBjc3x6v
Als+1k0/vojjio2XY4NW9i26x56BsN2IXyxdlRjed+zAlLK/7v0CBeDRLKjZdJIV
tRTb9LSdEVvPJicbiqfDVTlPtrdOiyAUZa8KBnPwncQVG9EHxkzhQ/qDUrZEMO0J
xbpFx5xTu+smLx8Bp1BO27nlFnkPe+18CXX6cRwolNWVFBZ0qzhlLCpuLP2cxr0G
68ySMdwJeRhpjSzZ29Ekq45MxqRaVrNNEmfje2rRkMrl+HwWQNclvcXwLeW5ET4a
V3WXcPMnmbQ3CEYRjdhWmOpEVlLfl7MtioilHYQggISnTtvfZ5dvq6aP50wQR8GX
aDF4XB9RRk9G2dwExZbnqi6Kf0sOStb+LKxZsZzYrB9D1QXQMy6gNEBARjhqoHqa
Lv2fNWp1Z4dFCLeXo8tF2jr6XKe8DR2YYc+VVVAzAC5N99m3JmwSotUxMURvuHSZ
ClQbdR4howqZ4vGIn5YZbzXAHNIBtxY9FoHAh7aAnnlzZcffaHncTIN7VZPlTva/
vxnri7usuTrXSqVcTU0xT/XrY434GlR2+AMdywSz4iPnyB2N1X4+HGlPGYi9reU5
JFc1edqvpjddG9oS5ai8+cxyYvac2DBfKxGMCwsgfGhcCzlRVIYEwqn68wfCcfCp
5K9cXr4efCZs+Q3ikLWUwT89sdBgk9TrgJOLsJPQbQ9UNlTHG0vuiL1gAy5Sd8+F
Nb7qy5v99CHd5NKcJYrurs6PZOkwxsljK28wsSPlw56lZNvXiS0Qui+PcrGCQieN
wwXsm2/5p+B7DLX+UMdcemHksdoBWGIELv3mwKr0S/vDTttwNfdyO7YGmXoq8YPK
fp4QMuyan9Lamy8Rm/NivYK2BO/rVLrSv0wLegDxcdgKiApGCiMO30azoeOs6Ms/
OWY9jsxU48F6+CpRO4V5R+fqKdbYaS1KB/9bH1o3ul5JAGWoQZ4c/lob8OhrUJ/V
2LXrrEjXORAkbJwD+c9jrdqW/RDXA710zVBhonRZivQMCf4AAtaw0YO+i/8e4w+3
f9bEMI3p8WM5Cy4rFZJJi1B5jE/mkgzvZgiAy7q+3JtMOaDF3erk7mNwi86YWLWM
1GR7aHk0nkMjLumLwqy7/7LFQB52TUWmnIpGhEuQ1X+REnpke2MJHRhsXv/g3cfS
2Ri0rrACqmw9OS7qQTuT2CJ04mzmMjNIiMnrTYILpYHRr3AKnsOeIXy7INA2wP1q
JgGyDp0cMrGLo0d9IHGBtc7E4B5n2BID4ZTJXuTijmJyifGML19cX6fMk1Qsqomb
7op3sHxp/S3zP+cO9A50qwt/NhiE+NBztykLG4yhVhaH8/IxhYkkKncCPs9W7FKh
H61nWjS3Rzn+HPexOvdgSantjSa8gpvzextem4Noz226ajkRKPyRYi8FNRGFO0hr
aAGewbjtWDxJxbOk+ilcyn1NOmXWgjIdbDc0Nf2ibl9OXY3vHgdodGrzELHlMswJ
cCBD/VWYGyG93Ph0YslXG3Ru/Isi/g72174rlx2hjoH2NGlvFi7mfAx3KgLyzd8I
gNMg3aKYq7BppgF9QOGkcjmYwLhrppA6FnG5SY8vfmTAXG1bFZIoejBEcoC0FHF9
fw9EPOkJZgdYhFPpSTvGam6ra1/M8m6y+pWAXyfmCoHGq1agLk0XgaRhQR0Bou+c
bJ2M2WACfoFPZyzWxzq+w4OWGHkRytb1AWDU8MNi92jRJLl5L7aIEbzHdlasI3qf
YW1huaoqc/hFzBwozqr5CjbLCWcC6Fy2+QxhBZEGH75HgSfDId+TB3YaMni3Kq3S
gNjqno27uhdDdxFNABGXFh8scef2MrjIx7EGnxTDdoAoDd57JtkexjmfPbJ8R6Cb
ZreWY3FU6ksLMIUzWJHMiALaBWzKCPipjLf40/LdOS5/QDiwkmEr8nJedVIPWkcg
xy+SIomuAlsvjeHqKY04tGAidQ2lijwEU5WEKMri+6cEDTLa33uEdC2k6H/J7y+w
dRPw+LS65YyhCy8JBvkW/UXzQnP+BerrKh7iKHzpZ2NNhO3J8l7FmCS5XG/b/CuH
ipOuaOSbtZ7LTg6l+4LQOP6PR0byHaVItwq+A2aaAC6Nc63PK9GF/jqZKb2dNNbu
qGFEK3Uapx9xaPH09TEF1wdfk3yf+eJhXKr68WVVYH5mHHipsO+LMy0OXyc47c/W
3nJ+Aa9cbDH/+onYLrVz9k6J0b5a2mNa1q5ibtQfNCz+YEbSyzKmvJCudV8NdM7x
xzHZquZrelgviUKzFKm5xk96fUsKeQHVH1FiXTc9UYIQwyHbcnX6rjFpPzitMmTU
EQSEqhP36xc3+hEUFznsW4NwshTsG+9/rd2kj0WWR0fupPz+tu6zqrVLkHLh6KRi
JZOtbtd+V5HNlss7NnXm1Epa7vrZonP3GUZNPO6Hr3ab/dv/Ll30Y5hBWSnF7D4h
AnX1rKMxorW6NRvHCX55CZOA6knkPEU+eHOfaDI71EqdpDO2a9EvQkNEAszM2bl8
eupCNZoDqdo4yZCmepZAGSPlpnt2HSZ8pdnKIb1RaPjEHyggSgwulb4YuvQaivyl
2VwS2yco7n4F4pIPgfVmkH886VmkCdRjwgd2cjzK2ooyHoTo1y8IxpxIMDwgl0IO
8HPSX9FBEwMN1PMWZbQB2vMRaEFHqK/bLF8fUw5eF9bvzYYt+XDmwDBJNCPQLRdR
F9gCu+EO4lAMk3ab5wryrPmjSoeV0I65PzrcAtfyFbAflJbciFtdhSvwzfydlZ16
k7DsvVSzY1NI9eRy413YdGhHJuz6Rm7aY1cJZeAbfhn88DLXFJD/zkE3+YcE3maJ
Gm2XJRBfk/S54W4gRV9tHG9p5mc2szUQlhpTc0s9QU886x3gtytxwl6Wa9Vkf8if
fjKt1VonnmOzJ8MvZQdRWDA0L8mcBSumoV8qsykiwhLbCg6GOZUNf+seIlH7b0Sl
T2lf/26b7FM+CnfG52s57sK/8QBCLfPrDfcZbxT11C8PZnpz95j0EjuN7D47yu1I
DoLoEHn09Ehbznt2iAxwgMMkoNxIenivyWsU4IG2SYD+6wiCdNhLnx2WJuumlL4V
q9Zaiyrm9ZnNuXQe0ZBXYZDd60+RycLE6r6rTAiFpbdzS6h0hoyWf46saiMHcpdb
B9R7GBdPdp9f4n94EVQvXv55UOsVBv5DDnYAGlPmfHqyjastF9josALjkS8EecQa
fjP4/AiWNV4JeVsMqM0KnKmQw7pFzn3498vDXbEXRWgo7Us607pQ7yRVyAxZYlWc
eh/+AWXHoXQkaku6coBjDX+hDyF3Zwah0asYcYCFLda7SIG6d5OPZvbncR3ZbYIj
WzzkDI0LRs1wK0F4PjNO3oEWixBHiEtGIbrMtLQO5d3ayIp4td5Y2VYhbhCgGOyy
RS5cnUyv/t9zBxrT/Mb6uronmSVg+KEsrc0NiW/lEFybRfbmdomUkp+/sMTiKRbS
UQUUfE0Dk8m0tSj4pYRv4rJzaqXbg8FOoYR9AvB11hj5c+vkx7p67VrlgNywG2BV
yNqBGyjI/OCXIVNKE1iYlVkpmk5zMYaeBIp4R1YUpTZ9XRehyYIJ+y91tCreBJz0
PWRyNTFVjJSXNhCwfEUTEg==
`protect END_PROTECTED
