`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KfuCr4DB2z1Z2CSkdYq2IBlakkx3cA17j0l7kBxaqfwJDo9fmf9z/lzaLkm3Vi2o
DJxiqpWwCxLd12o3xu1vqPi8aRI0LfZbe4OG4nW7oNkBw89pTcpdYohi1YKCA3n6
wUhzl32Jk2+g68nBBTh+2N0UmorB8cA7gmwz5jgt5OzDZKBZU5sod/lFbkkFEop6
g3Wi6uhkyTAaq73nusKWRJ5hWaJkT1RQBMTNGGQguSLeNbKR3CvDg2Dq1lE+vEGO
tvQtGh9ihl7nAYYsB9FUJmBW3ZYTVzZPLep0hPDI1HWMANpL8H/Qm1BzIuvn47my
yTsOS8XKXS1w5cgpqIWTin/H//UZcCe9jbblKiqWzOl67iWbUg6FM3hVKtrF7Tx0
2aC3Fo8TVVss7bf3HhE/a1Tgupd4vrtVZbgUsfL7wcTbYpwPhM2vG6CpoNyqUj8r
`protect END_PROTECTED
