`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6tzwRVe6ND7vi3Q03zfW4WTelddZuJF6vJTmif2BvcTJxCNRv+NgHjNnRX94baw
vTaeFzlqEdIeC1GtNLpK2fvR3zIyjbrrlUNJEaxYUW0/fAAvuurHBFp1Ba1YscJq
MC3krl4fro+EVEsEx3q3j658b9uBVrhpoyQjQ38KhGDJCnxanohZWEcKT189Y2BM
dsHy7bXl5sJAGwetUh5jY5OcJZWycKoYxOwHghtLzODoxDigC+8Nc23DFs+PjKcO
TDaTRSAemUTSTLGSAIvidXu0LoChck6t5ltspSXkf1nIlPf4/KP8nU2UfmfJ950j
QoiECGNihWXl+QwTuQaEjZS8fIsXmv6EY6wo+6gucNznJ22+J4DiRX2b9YkxeRjD
VmW7zlf9/XlUORg83h+LysA80nILqCTsqTWqg51GhIg=
`protect END_PROTECTED
