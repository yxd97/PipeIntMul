`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUsW6/6YdLYbz/Gf691Z5Cw8ezozc3Xn6/6seF5eZyAwlZMigBFgCrA3b8yhBCZX
+1xnnG9VmtymH7sipYebVIh0FIJqRpf6qR67w4+Z+NYJKhaqqJ1xgLEseWESh7wy
7XrZUW/08C61WgsjmnStSyVpKH0RBmEnrE5hAC1Ra8wR0+U85kOyXdRQ9aPPX6mb
bQqPMt1t8CvXqhL181sKTs/QPEZUXSisSEyldgL4xmLOqp8OEnlH+AARg+Om6sQ8
Mm4EtgV1RsQa6P6EVE2CdVdCqN7XVzQTLwzhUXqL791CdOIVGlSxGTwsC5+rwwpg
TXgUSORTEgawvNWvl9zkQgFua6K/cFkUQe40j+vSrv0JkJUJivj5DM5g431U8Aj+
k9pnihVjZOVgLOsh3tyyzZppuhKxHdjl3f3LxNh2yW4Ln3o4Dg2gQAEooeuj6c6o
`protect END_PROTECTED
