`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i+p9Rgyd1S76bjoJcZ5dpT8zOAMp0DdrAJaIFhFeD3OFuXGjUCZ90lAYEXVzeoGJ
FmWNAzBmI+jDb72HxuspQSstnTxkYdwj2IGLwspK97ms/JOzKpu2rARjr6ViEEm4
i87Ceo+thT36q1ewbrkmUJ5pHW2lEFNqFRbZqrLfXbrEgMRbUJk15uq7bY419v3K
s8dnLQq/iGZ7a3kI0ty7pk/DzSp4lFKPZf2pgsCUGe8ldM6qirJIlz5AqomMlT1z
5TeGcML+cJ6jCxBAXlPKZSn5KQsAWTR+Dkpg5jB/AEL1cklqeqsW7fEozbR8ylJi
tjoSCb/nhIwmCqMKUF25zA==
`protect END_PROTECTED
