`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nBRYBAILNtoGjMqtb0lsloYuaCdElINC8N1ZbILOwWHgUC3UAv7K5rcnycTcBjYk
01Gtn/kGJHZt/IqjL5XcRXcgdajk7tdtKzsgGnNW6OWvmqTr5b5Nst/99upLnFkS
CyY6mTbIJ2ikAe4X55/wYGoBSxK/5wXFGjA8Wud8ChZQTevZngaUJNcQ4CNYgUx/
cTat5ha+Rpn/caDmRD7ZkV4PGmulfubDx9sDPSiaDWWLThxKioXOsMI5ZOvrdYj8
rWkZm3IQLZdN06ViH1aInHHGVxqnuIrqLlAa6iVZKvLcnA3xQacW2RtaSUcwCDh0
vODssfpnffk0OuaPkN+Q1QGtGHmUTomf4KPYZT30CYzfp34CQRXkj+EjE9+zQ9mj
C8a27JfcUEJ187FUfVZdbn0ucpoy56v/IEgFfSS3Ym/6hl+He2oHRgAGy+xnzA0T
+99EjkCkQiCXBUTS0tINmYx9/p0pHKJjb3EWzggxPeWdnWvggdexMcGB2qjNv9tn
oak5syGMI0eGV7NmtFVQkVzhcQtMpoTnqreNSOI81KjvP95pY9/3reRnikGLWnhL
`protect END_PROTECTED
