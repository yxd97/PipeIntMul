`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+j36rtvsPgSG2Z+wi/gL1KWX+5QXQDqlNdP7ANBTjFuGLwiw3ry/49ffCpc2IoE
wexnl5esXaK2LA6988vdLfBagc7aeKHGLBqkwBPIkbsuTXceRZ7laYS2ZPjzICel
4fW/vpk8pZuE2CxPculmd8+/IQump1jiQ7g8xHIqxPzyUBFzbAly9VlMxO2DXPbL
Fph8YMKxHKER9Xa/Smoj2wMOhHtKBhO3yt7I2UZyraX7zyaDOyWswSCjlQBuI7lO
cfAfObN6easijRRwxPlCASAy3fPbkqimCl8brOt6NQeHERk+NWwyAxhCxm9o6meB
sjE2hQPJaTZGGLiNe0+ToO2GYoaDgtZWAiLVGhutnCoPZII1Ku3rZgX8IiXs0OIL
dNL1cA38R7EggPkyZ01u3Q==
`protect END_PROTECTED
