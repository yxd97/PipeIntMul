`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HgezHEbuPbNzPU5DzXKfjC1vYbBSJL0BpCM5rdIeIgOLnsQr1OgRlpAlVuJ2hwG1
W93dZ1uJ7UMtFyhtBuGdw8aCrZbzIS9Jdm+z7HTxmdfnwh0jCknkA1N74FTj1K6D
0tT6Rt31KaXQkG7fdfP/lxj/FNTMp0Fxl7b6PtBpwfT0dCAqMkqA5ukpfR1OXTYq
7LNib8bfGvMYl5JRjvguG/lvPA7L+ZSMGXU+/cljrg16aK9Wx9PVx/hgAsPCbxNu
fXICpvgrZOI3wzxk3blARotPId8TEWYdyifSK9COjoBPfM5EDpqhvX3WWaKIaMsN
riMdBG/YFtF9NAuWgZpdYHzccuyDcajBzsmBzGMh5zx8D0vDJcIVKjFlX6ZHO9LD
QZoNNqOp/KoY8dLJq0JAdU5VTaF7AloZ4e0IuB12HKwx9TvTA2WEKXkPlAujL6HS
`protect END_PROTECTED
