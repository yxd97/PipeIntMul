`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D++v3yleQcD3YfzH6hJzQZd9Lu1XzspphEqwY3TPXIjz7/aX1zIpn3240jsYKWlD
LvY1HfB98xEfiqPpHG5ulsAXo0FBCJhVyMpXgvaxUaqCEa5xX1GMd4AK3UIgo65m
O3FkWTkP9wyX7ebZNdS0jyY6msEQPll9f/BrmnjBXi/Bfvuc7h/hxchvD7j7hVkg
fujsZA222nnP5eBZRMNcRrpsBiJOrOR6CIGVo8VGWhGhTyZRiEZQJDM/LQi6P5WF
TIIO89CeTpSsH4BXdl56rg127yT2wMqD8xzgEU8LQ7tt2A83IgLEKqF/wlUhIWJG
90lnHn4LNSguG7mcQ9umeSmbHWwhdLq4W33D7bHmfZs=
`protect END_PROTECTED
