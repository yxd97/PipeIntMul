`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PEF1x5evcVOXbQQSzpnq09ag7RRdCXWmjiXx7dPfIQoXc2/ylJwxfm2lCrxWK67j
dBo0SibBp5TMShQDqbcJ6hRsHFL5sKBx2PePx4RlLJxoS8jh/I/8PellgHOn75Hg
JLFUoNjjcYSkJEpDVVLIr1I4rO23pxu9nqBRoktimec16gf47grMNAWdA+H+GeQl
YCfZ+7+rWwsBbcmvBh5RSaDak13qeQUs0qUqWpkGKO00FemW3jQb7ROxaTusrZyE
FclYxlpXaj5R2tkOrnguxhu3qRFSKCgeJLtZLvNal/jsmV4Gy1ZJv4uLTnFduR7V
YBgBjPyclAt6kDoybRnN/bT+H+G/PGwnrTrq9WutRqAkkXKdu73iDZ1Z19MpoqWB
/YChVHcO7gX45usqLTKu9Q==
`protect END_PROTECTED
