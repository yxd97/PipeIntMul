`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i6RipNJmQjIjDEHS7ic29+hth4WiEUN4d/ji+HUdqw1g8UjNihkdKRTdwKcmZ8Js
PAK/4ORm9pk+hqAHOdEm+PrInvFhZqzLQRb7Cr7x7h8mImnSKQE1CG+DfoPj6j3Q
Bl9dyTm5vipiCaX7/s8CZ8+/ugZR5I1BjvgHSYuOfrc/PGxaKrh12GZaU2e3hrx/
GmalrOh/WEYjhgsx6umJiqNE05fVG8uHAkJ/z3WTlhdB2Zp2BBxD6UHvOf2TrWzX
mdJfkXrgZ0vgOKJKfa3F7oll4iwEpWc1yArw4ZmcNj9o4dEmME00HXizK23yFdjh
OIGwEN4b2QVEDgBFRqEFVhulATQ7sRC8UHG1f7miYM3pbMFIQyG06wm8ZR0+cJHc
tUE0i05RlAwQdTLdQyTvn6RAIGNI2u5Pn9i3LywPZ7o6XC4ZU3BEzlHrOPmze/QV
PrIWxA7SRJ5qYjNJ6IhRR490Nz9rL1RsE9yVsq2+84KtlrWnZSOhNJLx4d4wPr6u
gJtV+L0lzUpERg0MBSWwnj4fy735tmmLqXuBo5HwIDpGwjXxfvLJBWibXyS89MO/
N2odLqRy6JIxXhs8EVHkU3Sbt+FnNnMqtWlett7lZwPxnVmUmPP/Ky2jYRzLdZ94
9mHJC52epu4fHAlRRStRMZjV5MiGOK3cMZ1zTSeJpCYKoz6O+nRJ3jTgm6lEnScA
pyMciP3Of1Wm5jVwMZMOx2UIZqRE6WWd9i5W08+JSEImNBIv/FL02ATu8zmHWhIo
PjiihRimRYgr6c+EuiDdySrFCYDAvq0aPCVGg7hslamF4iW8nLmsCB8jEmstBTMD
9n3TvRzfuzIkaXB0/N1o/QA2MNNA/9EGCq0Hrez1pIkJC3dK97umEUMqz3mF8fNT
`protect END_PROTECTED
