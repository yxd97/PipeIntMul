`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s2odMyIUXdSR9qlctbEx8TwDI7FSBhvbkMhrcZGZNVGzBiExGXdvUEIV2qHucx5e
wLglJ9clKd1BfhNqoMwGZ+eugxAPG+HZSvfWtT2CosO/8poredrL0tmboJEnf9We
ucJnryk4sjrWwusQMxUlers1HIU+LC4X/CX2UKsokU4PZnlCNOyKSkKqu0O2YnZ0
nog/JMdHYiTTUgWBMC2fjVItL2n71Gx8ZZBl8q3WMwx3BY9HqcQMp3ybz1XpDMox
sFevIYLxmRCR8i3xIjJa2b0Vkb5+xxKWENfgU8zCGrIuQDF96yfpX3AAHfHVPmCU
5GzpG9AMPE6+tdIa+oXSye88ySC8WXVUeYWAQCVTbRXql8U+0EaYIyrN/I61vHmU
0894tp61TCRDq0dRv/Rnc8O+rjWGzmG/6ZhW4vTRNQnsT6A8BsyjR/gkVoy00LDa
e1D+Htfyg78unjhug4yzjtT6pyhxKjG/RfLLXiG3g3dKNm8er8gZW1A4UanfO3LF
7rIaGtpmPOWrNx9TR0b8bQIKF1nO3jordg0XUkR7Guujcoc5UhSFQVHxq41sFJsg
0ji8rxYcocpnS7/77W13bMqFN57bLu/Brlho1R1YJabqk/rKhgageSELWjH3iHxa
VAk8n3TW7bZeRSGgvX7V/VaUX8YFba7LWMrf9XxicMiWWK1lbH51hiSkKL3zIxVH
bWF9YI0t9+/jBK8PlI4PonfHlsFyD4mZYHEkhtx9cnYAR3+BrkjBXNWlYWlTr6jR
LS9UeBGrRgHtevWBleuunh5Ubez8JYodGxYQ+43onNdqMSymtTPrIdALgKHjCIOm
hql9yEE9BtdyaPCW8tXapEnjypt35nXYwsjECUXDR3faFJtzr5zHABLroBLft2SF
QWsiMjdtQzqFZexQUHB00+uIjOS1S8U4xzIFrMGxK/o7lsrIMhERgCJiffCAx4hj
`protect END_PROTECTED
