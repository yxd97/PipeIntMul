`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqW673yGvR4HER6jNzcVGFulhvziRONqAcLLAaYzHRO4uUHuCN1t4d0WGDiFJu+y
0n7FXr8UyxtKjxk62bf3tBtitJ2ku6LXzXA4N1tujFNJrx0kVS3rxMKXaTQMD4jh
BJaSjz9zTckmmu5+AiycvNk6gtS1ZYZRYTCwcRCZoKeaSmKJE3rHZjTHfCpv1R7s
DFyUcEUEVPHDqxGIQITjqtYWpbijvgwxtmbPBSuB7VdezftDEYSinHR8CxAPziX3
7AjrSz+QTaHUVGJLvA2fdOBlid4gBqPdz5goE6QokBPnPGcRcBHtg6gopFTNVPRS
cqO9hWOKzez9LC12hAzCA8BmZUStHCWzi1OHr5ZUVateuOEynTh3UNqjJVAbq4C+
g5tNOQnw+7i5G001QJrU4YMM/Icsz2dbeKgvakaw0lyELfwFmGL6Fi38US1o5ToY
ifh6DgiOz0CmiR8vUlXfuqqtzwG+39gyb8g7nZoAhWf+GM+BDeudMoZkvuv29mcc
D5Em2eCX1W6se4XiYNEsqlVj5RJ2mB4SMP9m2EaSPNcTNShGr/qASpqRa1ejJjtc
9L2m3/fECNKo+5Ky1uiHcf5X2IS2IgoYvuGCa5qySiUCV4E1ikfzGIy8trdQJE/I
mI6GCPOzRYQaGBevWM66CgxI475MDCN2Wy20iSI45Ai/j5fQHO8u7xT1Uc/p+ueJ
FLMpoX/vOFwW6nKJTNkcZdE5YzuBdswwA885/6Jh5LHOUk3n0CG8mbJRniSYP1hy
n8qTRRBP4UBlEY/W5439mtwp6/w6GhgtTTR9nblrvhJU3GVIlYLpkwyNQtpRg7N6
3LbzJwZHYImFm06e1szy0Q==
`protect END_PROTECTED
