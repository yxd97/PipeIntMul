`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j52JFfYrVCyVjKa8+dM2xAt0gC5/tnlDyOyt5gAvtvdPWy54dAeez5cBgqXJDwzs
WGs5GKf3EnDL6NpN+p/Q1BkJcSzi2gbAXs9xQede5FjFss00xsTPp/ZnW9ld7kjm
J9duClbyNR14J/ZXPTLiE1iIuFN0Jt3xCagMGrA7l1UTIbKthQA59zb1kIa39GaH
kYwVMBziaFKu+p/0v3DVYITHdB9Z4qkBqEKDLJ9CzAoA2sJLUfzW6L4Sa0IsMu2Q
jvuel9mrZanu/sQCTXf/PCHsoxnljP3G6v5VV7Xs2DQdcp6y5t1FmEFm/8G0b7VY
UXGcp64Z2qskK/+eeVaaHA==
`protect END_PROTECTED
