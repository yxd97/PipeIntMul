`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gZmLn6PNC3kyTdN/7F9t+ZAr5h/qmQTEonUHiKtaa582sKfITX3vMjRVI6tqd9iy
L+5DSKHPbHEWhuN/Cx1frTZg/nKm9VxJTYLiItd4UlMmVn3hZrcGv5c2CxMi3ac7
yM9X46wcXsmyTMNZGBJyzsRNMEn97bAWrmSFNx0cvTBvJC/diIzqQyVxBqw1tPsa
HC95LYz+Vq10cmEiGYZi/kHaT6U0Qs66b2ATz6FTrwIVYaRbgmtqSkVEOQXfbhU+
daBJ8CXEZgpN+bHUxTXTGQ==
`protect END_PROTECTED
