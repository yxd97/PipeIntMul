`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vgPnbTFb9sHYfr4g2YVZ0aji//l5rxJ3ouH04LJ8wO8d/YG9+syVygXRF0qX7ekC
VaGxsxElf0hOUzcpkBQVupFR9jZwYZ+oAWENhAzZrHh6dQaULIJoUi55LjdOrXRN
ALG7xFCShKddmz4p36KziHtWs3GqMU1Y/Y+fb2UCF8FKMzwvQaRZ/MnlZ8vmzURr
fyYVG6Sudpi4cgYp5rJ4RV5GUmW9fQapWPsFxW0CtNRYec6KCtsiNBx8KdfWF4bc
wd+hYDDl6FOzP846a61bumy7T0Pv0oPMj5j7Rc9YjtwsMl3LV1h22OS4EjAMVKD0
5viE6WMf1Ho9xx86riZ4A/oSNf6iCoIO3sk3F4T8y6caiFy0IxpA61p/7OYlwIeE
XJ+5j7Io+2UMVZ2Y4VsG1eF65Z9YEmTt93EuEbMSOv1Xpxg/3NZ/zXe3DbIYuk3W
GiJv965HONHoiUJpfYMIKE6EU/L1yjTYw7A5hhI0cDBUtoLLDfT6dDCJRFzAyR3F
OjkPlgcfjje322u0awu/ioA+mXXiPFejm0ArnAmJCqI=
`protect END_PROTECTED
