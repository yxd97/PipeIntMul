`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukLsxBNzPbLoAXGkp8/2OjjC+EZJH6P6CWLwJSFBwLu2V3on792rC0T4TiqoA3lp
ge6J7KaF5lxlFFxMVKPP4AKkb6VN7I4ik+cjl+AZMvPDoDWcuvfGnk1Y1zy6W7cs
PuXMdTjobo8V9u66dSx6hMDdGl89eJ+niB5gk7vGeQhGbmyORSjqWAZJL5yVAUhz
wq4+6WvHqvF9xMcwq9EuLT0H5CtvkwBWOECujtJZ7V5aXtSjgBAYORpaUSSEahjU
rW+T87ksL24aWGGDOAua4EAhYKptmMlNA13dq21qGIakhmNpoanPillU6xW6j65O
d6yLXnNNNE6hNBYiYCW3aiyr0w8Qc5keLd/XWkYr4rwwqCQtlf2iNt+PcLE/GNUU
G36mHvBlmpd6mL9ADZwcYRjeFegrESTGY3EvxT+DbJnaMFow17SpglN7aqR8zboD
GO/05R5Uzo4xQEuhigoXNBBajp5695pibAt0NBaK8XeF2eMseuQ0rMt34fFIYwQc
t+kiBleAUgydDxt9U/lhVAE0HKl7gk5tnGfdcTAS6RRBjr0qe2U/HR8qU48sPNVe
R8K90XlQ1RuWnkOdDPQFvd0h1kh+Hd+ZKCdVis80+NqTjznUnmvAIXCHIkCBlnwx
d6KPTcZq67UrULmHsCumFWBPTknp50wimk9rf7xWrooVP1Zb3eCNzYujuMuZR9ko
DNHBoksxxz1EoKDVPez3nM5T3HD4CoVNDRWWEbgJb4TgYlH4/fixqcYy2VYkGkgT
iyrMs6bmrLr6w0Lg5C7CviEmNex/4s6AvUVKhBUQgW9+HP4B8DutKyxb/W/SPHCR
mBIbH1R0xFDYQp9K0RDcgerAkYZChx5JYM9Aju4FrvvJSb4F6fd1lmxKcVBRkpZm
EAOB2bU34p+iWf4KUFJ/xQ==
`protect END_PROTECTED
