`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2fjXXPzRPGF1FZ9q1U2vyFw20B0zeKlAjEVEKxEx4YFJ4BQ2HkwXUVrdYGS026Xy
hxOvkcsdmBGu2H+HAzw/IyqaZ69N1MeED+mrN+h8mxCN1/sKMf/4UYMZkafn4y6V
6B+kiBjgCwNHDEUMq5NMLq9l6Iu+CEFdx7Iy8GjeHgmvRBsylLnSVCny1xdiHglb
y1tmEwykk2eJrQBv5eiOYFtp6WnYYw19o8fgjE5RZ/0PghsScSSHKIF7qfrPXj+z
YP7Vg/gSo+HZ4IJdbBUMBhZM4iGQ+mHejDPp+ZpXoP0qqEUaqrG0jCHmNXAvPdqt
sI89O0WVb/yh46GHn+uRT1p+T+DVqBoFA4jrTlYtFJVuE4v7ORb9/OcdhBfY+Uzl
t42Oy6DFNtoRGWRCJbAzbPxwpHCjEYljvEDrPDhxVBUYkXYbRuf6ns6Tn+9iT9av
R/T881M/eCDuWX8wTvJ4UZ8BgTMAT8Cc0z3qWETpArs3rPeckNnQqewC9ZO4tPH1
iNKaZc6AiuS4UBluUqEDahsayzd5my7DVGQgoL7m+nd+Ox12w7LffYiMZZ94sq9B
6YahM0BlecdUL+ydqo826+jBsshdcQlwlGjzoY0Qw5U=
`protect END_PROTECTED
