`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
APat3VRzemvbGLl92ZpwXXwpJaE0W626y6tN7IoiKxI4M+KOqeVa1zBI38Q6ePTJ
LB1nYCRX9JUj+d3cJXu7zoNiUZWRdfhcXRo3q44/fYeCVBBAnrXqPFZra9aJc6wr
iHdDbexDXbnjY90vl1Yq9yBz8SLGiR6VOFwLAzS3b/9t6E5Knjb1xCUbXVKvvUGm
hnw1BE3Dnr+9oAufZiqH2oms3wsdGjUDHm+TuGFPbDendIfBWtE0agCtYhaWyjSW
uKbGrrWx/b8LXKgnIMdLrUcmrATpYot+eSlmWz3ILshsAkJmqPpaeAP6NCnfsTcM
fSp3DRzNIZHu3CJ/Wry7zrS8gzZStr3EaFFh/2jJ3GEblEK/La2mATWcS6+kO0mf
eKWp4hrtIWjVcgmBVlLbhq1ro+VKwrMCs4MleMjUSr/mFVx2gU1GISfgZDA3Y/Lx
PXERCciLW2JwSSLta38q3AUkilGImjlgmzi76v+RtDAahcZonESE6UeMqQ7pc4vb
fWCNqi6fBL8B91cR25CO/G82nb7/e34fnTzZ/Yki8+IlgxCKk2jo8t++BKVlKLjg
bJZfsUgKgrhllpRu3Fbb7ZwkYFjGcYGmWmRnTTk5amM08W8mnlM8dMrD/N6tIJXc
DZ7BpX5QbkX1iQ7U/8C3MnIMO27Cu6Ftstb5IUPWFWyYDAUDryJB92fqJbKWzz7v
FIHmDsXXJJ30gKB5gmixOht/+mbDAj1NGmJUdcS3geKuAv+NoMIzGws+lGdH0AK/
bs8yYm6J8NGr+CrC43iy5g==
`protect END_PROTECTED
