`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0oeuuRBnRBK/Xcc5SMucTxMd9+glEpxzl5/H4xBYhmE/hA4CJAplwEOt6TTgD0jZ
TcKxkWaH1ZSDtQJ88oYeVP2zl94nLwHlMvisQDYdACXc3iVlkc//+G1wUm7p8G/9
BNmI8ubtzShWfOKv4AXAkx9Uh4FSIv1aJS0G+DzVADl/Gpnep6ZJG+Wvuua7K7gX
7BTb8WhJP29bNpQ6Dl1G7N4Ioevyctsk7O4DPY3vk55rKrb83guf5nwo37E/Mfy4
QgbTX86k5WczIeu20hT2xmw/D+ZhlPv4s85Puu+lZu6lEl54iJgJReS2vxLWg3mk
kM8QKPceAWLzh3gmAClOoFY3uaiRN95wJBru/86Trtk520lO/My0iPIhkxc7TBdD
v6AOBRn5tBCGdqbgxKhjItlN5dXaoor4rna1J6HhgSpFlDG39VCLDgpxg3iwEvA4
FdByOlErxZhAjbo8r/dCMZjpLxxPVz/7ADAuMLoHTC9F1k9nI7VJZ9Kza2H8f8rV
5RWzWTj892sc4bNqe3BsJDQMwQK8DD+DHiQC/F7KKmU=
`protect END_PROTECTED
