`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zywv5f5cd5VICPlS+az8wms0rURhflV59xWs3DX8u+4luhfPGEy+eZgFUDhggQQ4
Wc1Pgh+T3GxJpyCl/zq2Um8dqymLXMsaEkhFcYi1uqBADrbXuFWJKoo/s9xwWu7D
CgSKLCPR3JFieX/BToYaMQHzQqUWcSNH3Q7I6HzIv3arsNRT3nzKM+v7jI4NCSqk
6HQ0/BMu9Sc+0yWCFnOm+9JVXp0FlDzjKn44foPvj12m4D/um69jC9MelWhBnIX6
SegYm712xKjhFCMyS6PYlMO2iVoERoW6DM5+0uvqwS0JJGbS7y0opHs0Y2kmA/rh
lIeG8Poo5nZrvKStgSUtME5XHGv+wqfuXbIb8siSRj0=
`protect END_PROTECTED
