`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A3b1wSg+7a/4BBTUi2XGd/rN9rqUxv2MkpyPxmY0y17ar/tGdx3I2r59UrixBt74
u0T4vlNs1pqnoMLAPcMaK5e5VTpQpNF5pETrWQckk+Lh430dK2tLOI9WrH+vHs7K
/2Y1NbuRIbVAM4TSvWqVIpCsiz20XXRUblV20l8Oar6EnYVJuoDQ9qdzS/5pAbxH
ZGv955jvWWOf+VbxroEmDSAE0vQS9TODuo4zqiKDjdqHKh1eANVlsDYErA3d1P92
rf3jtng98EkDs7sqdSXUUDFlXk5EoH4jdyw7ArpaApjaGWgh3guRPYSk4fbxVwr4
`protect END_PROTECTED
