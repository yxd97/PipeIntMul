`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
23JGOBAXbpzPtYtI0ENtsGR1hvEGeqCoGTZ5QjyikxyWdQY9fzhflbC0AGm2BOqC
xE4pPekCe8GXfsGejcLiACxJWZoqOzA36Wxdhq9/CoEE6qyE6AB9GLEQ5BR+8jR7
ziHBwZNuN7cW8X7UGJubmkp5YFKgu0zBLoRokV9kLSJBxx9Bqsb6lPuXUgChqjNn
WtRWhJYuac4FHzyXk51tXmE3QEeixi8pOm/T5/46Xt5GCVKRgbE+vfQFIhPPY88I
efK+XQD9Ghg34Mv84Fb5vUEGGb3/B6nhQgAi/GelZkEmxh0ARE/77kRAjWbfQvp3
KkRTNCZqK2O5fYNXNusUHf3RejBW34VjEleKDD4rQ23uBGUyDEu8Sbq7aICSQoKg
wenIOBJfuwsqwRNiVcYoldWBHn/Bpb/LI47kxyf/DagYZqbfmpJfypPEbKZd+3GH
Hi9JUsvDAg5trBh6GwsjIxNgtAszw+a/+Vbr0d4x7h9PEbaGr8w/zD3D4PUu6RCf
D13brIIvEBiUP5CYUib8nyKic/wM1SVijc/KCQGCtQGQ9NS7lfPziggz9leVD2Ou
8aYxvNlYmqUd2mIWgO5PjkYhpK75JdI+QsBmH5iAFy5mZdvrKnwyxjzNbBMZj8+/
7k52S271Ltzv/zbsRf4PisUIdBRbODMo2ktwBWraQgH9QWmwIyULBxTSRZEM9gVJ
YfpmtK/CbXEv4s4BISoY1g5vypw+Db234rUHfpV7RmVGh+qHQcojLnw+AtQ7MBMt
m28z+191K22tFrOcDjp5AA==
`protect END_PROTECTED
