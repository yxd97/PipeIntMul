`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7z6hwTk1WH/0wTZwIEvhNeglupPZg+JcMQha46otw5eXNNUsthsb/Gvhja88SRm9
JDZIAijypX1m936XfuRlx47bcSTYDlAebI8rJR2xFGBUlXpa0OFM8AZny0MkrJxC
xjsoEIlUuAKANWdfY1YjXnn1NQvu0+a3evJFnXC7ZQQylwweMjONEAwbJFU1NKK0
L6uX+kb8T+Jso2H9KIY8esCGNSYmP13kttH8Gr5kHHO0MHYVwVN60M/1XPLrUeVd
qw9yHf3oh663gfyR4bTmGXaeMnDF8ephoWL+8nQ4Q4Jsxu3DNZHRNmd6MlmrMyyw
X6z3G3o743Qf4/IQk4PKsfvDMgVtXcxk74k4P3TBPh1junsrd+y2iar7NlhpRgeh
IIH1aCpeuY4P5xHSFuaZKmZGkZLwJ03y+fcwREk6IDDh1WkXzSR0cuiV/cY1TSbH
zZKU7hh/f6KzD2hp2nA8CmAXmNgIaAM6Yms4qyOiztyEq2nDUPR2upIqgnjDNwZJ
h9zw0AzqVYZh2jL4HOKtnhcajceJE0MjDbyiFCjp11U=
`protect END_PROTECTED
