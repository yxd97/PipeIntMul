`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qR/gj6HrUIFTAsOgKInr6/4pNEqdmwQqPDU1X9Ztux6pZyuaehuN0oJm0TfuN+HB
vjsGhnkCKxnOJMk6psmjTK4qnCes4KLhXSbjFBdGE6Qlg8gqnmgkHRXbhii7u0KB
3DoOTNNOKVvR9cabx5C6ImL0UD3ai20JlwBH4OCiAYCt+CVViSuVdXt3Tig8+PgK
8PpJ4Y1GNbgbdbVjPQGK0Y9pT2DC6NUwOdb3g9Ea+a8u+tGPBI78gsO5hUc/cYwS
5BkR0tG2dt/al+B1Smjfmm3qEoATogHyXDzyR9/WITl1Rq25kpF1f36c6+p3gf6b
e8cFwsAy83YvqXnuSf7WmA82QJSt/2rYwCmZSyeLEOlROQ8YSfX1Rr/2y4bS3aLZ
vMmlKeAiK5ZRHUudHsvvof5yk7CWPcZcMMyxsUonptN7A7aa5YjYj9mNDrpiYAq0
apJ0uBtztJY/tqyulWoHN1DfhsM3tTXAxrW/3mOafpyaOEko397l8Wf3DuzINmKL
5C+Ddcl0FV+rBnwfvoRYUUhinvuNUNZJ7ZUaHwM2w80YPGqPijV8+Y+SCm2D8N5T
akval8m6jDcnjpqSll/EbvoihcDb1IgtpMqty0LKlNOO1poVE6HoVdeiidjOxKTj
P61v45tGAek2xEcYf3iLJw==
`protect END_PROTECTED
