`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U539HZs304x6yCM/UBSvPFruM0svzvc6p+EclTRGygvcMMtZpNd69SSS/KTbI8eX
PC4GWnGGLoqDTvfL9qSHdw/F0tjenxkvt59VTqGtGgX3cZQQY1+eOg38drc5XmyV
TSTMgxi7G8V8/U2TIOi1dFXXelqqeAB6bbTm+6xHE1YGOowJ9tjB9utexaxgvQYl
HV6nBiBOb8nP8aDlpu/6muPa8QVhwNZ6DQIKXOKUUoeklmH27nn5/ibGcuqqd/XY
lE8GkYrqUR663c7YejZGaGOsgwqJA3UodfiAPHnueCQ=
`protect END_PROTECTED
