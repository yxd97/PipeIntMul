`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FFGS4uK0UevsflVReqQjA9XAG9S2+mZgYTDyS9EZXK5pvKhLSxU2F4ZA61bPY5Sh
iXqQuwxorJHZ38cqJFUrS84Jb7bI+rJNOSKCczkUFUHCuUU1+cZ3sBEFV6tCnEU+
La6V5P43G/5138564TEv5z0syDNXmf/i91Ii0wYh9i2nJfhLhof1Fh9+CpAGo5mI
2KYQEiBVrxEXjwuRNi6KHW5y1ja+bIXFTW0fFA19W4vxsvAhSf7LGIEJF+ju0g+j
e8t9yE1BvQ+kEeU1yu/MELIdKZ7K/GikIuqr1v25z8e63YBpbcDcxtzeoOHz/hN3
7kbO8KzGFMzWvjZwf6Sp5GtHTLi01j6K88qBpoq+0e0=
`protect END_PROTECTED
