`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDDfDTEa2YVe9zOU2//WLDD0jVD3pYkyJsjCy0ouyivyEm0LvU9KlDKNHNzz+FbA
nPvQIpw+4jFANIEHMV5hIeEgW+FRFJxx/Nqmrc4BbxCNsy5i+yjHL+VDpmHHq7hL
6x9tFqFXI65PaBzcg0LKqIgCmVxusL/KWVB6zehvSzeHWmcZGsV6TBFEsnCUbMXg
rYIGYOD+k85L1jv1gGV2hJGH56GxDmSI7Xe9W2E/ki5FA/d70mV6wAp3XMC7Burw
vCEHG6GNMBb7htdWTRcxczXh5r4iRO3ZvYopuKx9pqSYx/oEPdGsggTztMchKvH3
ldobYAaOjA93xDEoSp/2cpchYkckXJWJtJCODFiOQ2RemeqAB1MeOW/2fsn3dbzX
tfVXcZuL2NtARnUXEObReI0APhG0XpVfyIvvyOiHQdc0uMHaw0lppINUzpLK/iz5
Kym67TdNwPhDXhf1T3GJyktIW8zQapjhpAVxonueGUXq171k5ang4Nhylbkxdxie
JK0N3ZmBVAXGiVE/CxfQEtSeQ9AKSoLAI4nnIcYVEcVyz79fXsBjtXpgXMJnMDEU
XqUH8FxyKJufFp5HSb4E0Q==
`protect END_PROTECTED
