`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
enEVKcn0euZ9tepuaFs4pvsKVOUTCgdsaFEzo99aNpV/O82naDuRa5x47HO8a7Lp
1FX5+d6N1wILB/BEqKvrsdXRs0NblfRi+pK5Qi13q1ZJBzjYZkPsSaA1E2ckrt3l
EVltsI3ETPTC2pxDPA8L7doowi4jx/m6yEX9aDLZMytkt1KQGABsjycFTAXQevI8
8Q6nlv6qapDJKR4+79p2u6fWwPBsh2YgyDHnEnBKzS45gipD7JCCfuukFDfo4dad
CD65qqZVLLHTN+KRxgEYZhyUutnmtB7CnAXxdgLFNHpY1ZvvBhiISM+mcQlYSuhN
YOCVakZA7lOG9Bid6KOPQuZdeW9u07CFKN/+1md0iOdjTHWQPlSE6yvP+5gBZXrX
b3UYjyFY0YZdoIwAVAMHL5G0Wsn/pyNLN0mzCod9qIrmEn9TVXqKrQ8kxQXbaIL0
6fyp0ASlFu0MIut3RS8I1tH6gJpljO83yjkzfozuvnLHEVbgtsCxFEY9gbNoZD8K
hVvhmuvDLbdQMql9hzk1SXL//07yH8GLZznaJasnUFcww1BQk8uqFLtInkYaZYMj
jCKoZMw1m9g/U8fmqbMmIITphbJTihA2BkaLP0oFDdZZjReZnoD5apOTN0RAJhzj
tK8/ed9/v+vL/AwVKg2vboSm390Im5CjXzbwlME8qQUal4T8NPfTW4zSZPkOWZjB
X5S57GMcv5eFcIN0Xid/zpgxhYJxcMlw/BDAYeJQZLI3s8mjvpH/HAcsNtrHp8qY
fX13//s66mkPgqZuw/S2xupCtWGCOz8bd9scXJ0WA8goL+HVSF5ExzldfjtmSVs0
1p/XK0Xuq+cX6fOe9BqguYhWLzbTbon9S6zsFCh3DUCWThkkrjv1aj/k7GZTxQU5
/hC1xpjrir/QMJLyXFkW8gmiC4HKScT4/tL5fTwct9Lm2F1p+nNHGy8QMn4bWPnO
5v1JT1kfM20xw72Xx82PtIAHJ55DOwrhvi42/n7bFooVOn2YCmRg/Opz3zrPWaO1
d4n1eR07Jmy64IBp5Dl0/4oxuby/+F3S9AorGJIa1Ux5bqOuBRya8jxf6jGRxns0
Ei9x45R71L+cSvRRKZBm0aGYQ3Peg2/as1iBqH+8h3v2AWxy2omUwog9Rff+/kdA
4OxB51BpjdMIi48K1s0NZfxpuM3+21l/elSBanYNoRhGfMdSlg8F4sJPKe4IDVNL
R0NvTgnceptCIIRxCycbGo6y9TSBuX/DtiA9699YXETFqv4qQMV/Laexmp/Ps7ey
d+Ps7Er/Yt3FuAIhewDKPfEvv7kmMb2/GRZUtOYYEpm8lDpM61Tt2Ve5NqZmm3ws
i7WiWb3KCgSeW72c92PVU2VCgULTTRaO1KAkwj6ZJx4SAhiH43ntiHyQxyvYYIwb
OJrPPgwnZOsNi/hWx5l/PXyVrdn80WlfOqY9uTV53aUp67aMEl+v05X/2PKH1OMI
R/Lt6+IMVISncOZUZ9MTQ5fIDr44FGz5ZkD2oBwuqOXRr7RVGC6MKQPHUnPpHsDY
Qj0Rft1prMyQ7TDmPjcL73FcYe8njDYE60oYa4SlgqNJmm/Rhq6hVnQWU/2WetFO
jOw1q7QOocRDGrbYFDRxjT32m/yO8UZE+2owon3eOlqcVC3GmhCG8r224Muwv7V4
gUYi4ycBiw7Wetqzeu/iJSXynzrWSP4mo/O5abiFPKZnqBg3QlyoH1/gQJfzBgJe
+kMiEjyJsPX1j/f+7yG61rvoyGtq4MzAHCr8UKNXz6KuxInf7L9It23lw/3pWSWm
hcZEF2/kZQ9ny29jW3x8FTcVdl88xBlmJFmSEL9D97vQq6qKvKx2nOIx6KVMzLs1
cMhLdALGc58zzlFJ5QcghCjJxKVCziR69fssju+k9i2JxBGKoizjywWmqvkRjgmf
`protect END_PROTECTED
