`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqv3A9ivIPEloH4GZPcKv5AmYCmXDk+UkBwmLDM5ykfwX3oC5NlxtrLW4Jp6JdeR
B1HDA1qvszkiH/M8/ov9szniHVoN3spui2/PXK45URi4WcDtfHo3Fxn6O1yDAS+r
a7r4E1bGXhfzYmKz2y2H2X0wogIe9IhOh8vn14UIkANoSpmSnEQxvhhd1o60PFEH
vt1bpkUWkJJ+kvZyut7wVRes5ZFaDAUQS8Ghr/q3TR2uWaEN7Smzar2PpRdltTLq
yq4GpnDWXBJxRgAEi56u37wblKajTWcOsAg/ssyh+kiMTK/h1VZ6MPUv/DrU7GKN
GmRVjeof4l1AmSLDP7+LAtIcdXIYgkgotST5iDvkKZmcqRfMj7tAM7F/HglJRHou
suLWUhK9satQykd8YfbmSg==
`protect END_PROTECTED
