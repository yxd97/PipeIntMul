`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OgXSwygcskbZyXZYahL8DgFVBB+4junORzSr03OqbrE5c45e1UtfWisEYp8v4JYn
Zx35QSPJuDb9LyhVpV/KG6rMOt6PzAmGUw57dpIrSAlG15hfkQd06RsTPrCipybT
/GZjWxc6v4dK9VUX3Tq29cPp7JS7PsOeDGy6T9hxtgqRfkFupUEb3Xv8d6Xr/XP1
2L+3vFs8H5nGFny99ZioVfGqxTZENEXLh+SwEeQnEcNL+E9RCopqwJUcNTaOAwGJ
wvsfZ5sWo/+dxrOegZk+4BxRE4CSQd806p6zQJicYB4hQQicYLt9DqcQbOJwfKUW
S82wc7Exxx9SVaeGF+FxJ5xWOjzNtxsnYd1lbCQSBBny5WOxwkd7pItI92ugFcad
o+GNJr+4bdQ9neXo7acsTAkUBiXnf9xcWHqmoIm2NE4sFYfD5+DGmNYVRxQKUc5G
SrDjH8F4/0/yXhoRm66T4S2FpFbYBKcSqIJi5l/HiCN7uJIpm+B5Xs3xXYoCg3FW
wnGEAWzvRW6d4Zv2FW+utEs5QsTVKo/ipGHzVAwDU2hHiuuQaPPWJyRTrjoAMK6K
18fXdUHLG1povqKlkgOP9eKmvPnIunv/NkHrKl8I5adm6EXlvPKgaS9JpJ5sMnZw
Ityip1lErYGujVW9NarqiQBp0pTwnufi022/mLA+i2b6UY8+nJWVYKwj2o/o3a7j
tU5MZNlvyGOhnlxqDHOWr2QCVZ9p9V7En7pH78rDI2+mLN9WY13shFW+ktsxjdAk
OdDIl7ol2roNyXGM+NyhpF4f/muyU+jndo8iOKGiXwSRacxxlHfy+OXtCRbdHCRU
aXQk4lR2QJaG2bi0VxxvwiSEdkDwkSArYXo5tWp9i2jJDlQIwYmi9TuncI8/oYYP
O9bRWswkQyOQ9CDIVdCU1g==
`protect END_PROTECTED
