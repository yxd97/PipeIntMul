`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zv3QWBJ9J7InOx5kgR3PZCCg4nZfLUSoLsFpEmkJwB+Yt7amQTWrbhC7nRNEzi2
z/XklwcmTKwEERCchBFmof2KLEmJdEE6kTnotaIyov7trY1xtBWfL7/P8RiNEy7J
927Stgd682zyIfpHjS4D2jQF6bLig3AoePyTAP73juY0j9jYoputlXiy1JqrrwHi
ETyPzZbx93hXY5aaVqAn7E+sl6WZWUuFCNjVRT10mf+VFidB4k3KQ+DIRZrukqmz
w+IQnhbowy+sJQ3snz+WDk2ic6iqvdY5Ut6ISD84yUX5Bmh90Ii/urAIYCvH8tFw
BMzMABlzfhQuqY2rl5BhqWqudvHUGIg2LV+5GWl4iCovvSXM+oTFkaoTkytO7dQE
HlahUyvXXySAQPyxdGRkiT1mOw9WNld8jFnHKahJ9NGT1CTN9vMMnGobtRUH75iA
`protect END_PROTECTED
