`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCB2Tl37e4xphWpNPZT5Jf9bKND8bETDoFIC8SQ8Rkb2rEnhaqn4/AmMMWXntcIy
NsZ0URsmEsC2VzRLV5ynx60RFxJjnzArXmoZ9sXk01w+hG96d6NJw3QClQVIFV2l
NpDp27HsfWmrmHwMp4QZ9fx/2NjBfkE0Wly/ssNeLdMaNuVll2ZU4/s8y5PNjzv3
bmE6K+wreO/kZ7y0eWKRDbYak1frf9SdMH+kAsWcn+lQR0DaxN7DunIHAJbnlvWN
Q/pLpF58icPNjmlLzqY1M0YT/8s64KeyGNlcyCpBElfOQEijet/vYBv25V6Qv7XD
U/q4I6tL5tmOUpK2xIo6JmFwqyFr2C6ddlZuJG43UirltmyDN42IghX+tMWVvKQM
fmlqfEp4Zpd6Bp6wVCpEzYcUVypA0EExScevYIKZAIDrszmRQ+j/T6YT5g/eKtOe
+ZUotQWhfful7OacdOdLdLTr6tt7pumLamO60bock/E=
`protect END_PROTECTED
