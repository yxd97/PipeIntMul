`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c90nA5zOTEwTKhx77gAmZrmG9zFq4DOpUQZFcp9fBj2A0Yr6nzZ6aenB+cy4007H
o+edFcUALvKY9PmiRjrnIsys/MbB+PWyRxqYacgHb+iE9q0NuVvyaezOZcby13mq
GngjFclZYC/4YRqr6kYX0gp6I3rur7olSoOYvpuQofbJ9sDCbOT4UwnIyALJSrqz
9ySbzRJXyrx0voOBF7MepR8WLoZMYZhSvYQJEqF0bJ6GhBTe1aMop4jI+Kg3DlTs
ZSU0uSVMFGVyL9qJ4+ty1TDd1RzicP834sNVs5WCE9JRl4JeWeWlG5Ok4kOcWdwK
EZ6mmD59NYs0HpabX9qbqmjLbcp/xAgDeZwkpmNhWNFOCvTu69qx7+jbzWzbaG3r
F3xtux09pPTqu72KG51LVgaqgviu7xtlOfOCAe2DrLUsRP+D9X9oo/Yf+Mwkvz3u
SPFTxHbjuhbDxbV/ib9tBvLPyG0MVRxBlRPJF8pqYX8NFVgIzr3JVhIR4PmU8L3x
sE7WDjiTig/VfL6iSM6EagcFuW4Cg/T7TCb20WHnqiNBt5qeGz618EZiZLU+Z6kP
nZrr9uDp0ZBO/xyTAYGL+AI110OJjZA0U91u1rIT6gt+VFrUSJmsQJO95clYzYQh
PUHS0lIxfi1bHj1mwwj+tDKtuOLD2drZ9hILdTwlbgNpFmLVkm0d/nVRVgbaX8Ph
MQElhCdEpfyi9vsAFJwxFLrYdCbbTSILE/xUSJHB7WiodUbQz2YxZVXrONM26m3A
88b9oqYBRNPc98tJG1pb5A+PivJaSzoKItKGmG2htnk=
`protect END_PROTECTED
