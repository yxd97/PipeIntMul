`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WP83tuuV3q2QCXzIv02P6FCUQKfaOkNhpI3rtuBNoq5Lp4/KMWoFULS7d5RDvA5M
WvW8luOlT2+e6sBT0KyxcNcOogrXBCsgrtwQx9Gs8EE3kEBC7pHIigVOz4nL36/5
StTKYq8EupAma+Ryibijw1Me0SUfSmDiygdYSAjGr5rQZPE6dzEhKa7C7320Wk0Y
avyw9UfyxaBWwP6qu5C041jCAa8DHxKZUU/KfTrzohw30DR9wNFdrSSmsdn4TWGM
ifjWbc2QzT/ytcycfrxRjNwCLgAOycUyzUprMAESjIvINb/oHUrX+KmcZIv2SIeA
UoTSTTTEUaTMD3AQqoGcRRuzMgw3Vpmm1G+Sikbr6v22ndlgMi66hDH4K3G9nniG
PqdQoU0JDz5ooxpgcjd9i6sIjq9qjdq2PBZHOve7yJjC4SIZ1BYZZx9JTLHULj0r
TLjX3iZp0cu/TzSEQ6vyhpM9Sl/Ust0tpltwE4Xm0jw=
`protect END_PROTECTED
