`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SOub3bP4OHiXoEEjcMjBWB/2bruGIOjbptEn0yiMeIRn4QEz0YfF5hWy7tRpSiq3
Ldfvq5rzI330dlAg18NWdVbWRc7ZqtVcZJQ+dUGNAc34FbP77S7jwkI7DudJBgwS
qIZyveIi2f16Tvqw3vjqxldTwuC6mrWj2853I9A7v9xakkOEHarcp08OtuLo9wTa
lsCbAQrrSVdBcbmR8Q9/sDor1+Llonpju1QrMmiteu9YJyfZkmNdTytHFWWH8mPE
oKkFC7hD9GxnrcdA3LbmEQO9tx59jY1e2f5w8hN22q5ZB8T828HMFK85CP+wcNJe
zUsdVj3mZCPwWcSOwb8obAfEKdkWKhlhP0S+uXc/eC6LrJ2xidW+bhri+rT8w8Py
TcpirGFxVjOeAc9fIC5hk/LJM2RmZiqIAjQLIx7JwG8ifxkLr2079al8uR0cdmXh
Rwm55jONOIQtmV/w8Ds5vyRLkydWVWEWoS8ooZNId8bSz05os+H82plbz9OFQdwf
`protect END_PROTECTED
