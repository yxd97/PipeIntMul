`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KEPBcLrRiejoW12arrt6sMLziWcm7mpO+fSriLabiSL13IaAkQtfQygj8P6TZvI3
BWtpn8/r6kC8ogSvZQMxCOViThTkef0GAFd+lzXor/AbJ97ZuYjBqA5fIgOpKWwh
oB6Hx3lsren9rTD6HCbogoqmkfZkE3qMZdLy/15pEw44O5h1B2UNzRZKA86DZtII
3bOHFsRaBvNkwChjNXED9vaJfOVCVFa5n7u+GGTEl1jugpZaCSOTvAfABpVvOgMV
xkl1nDdVB8ZfQshPnCggXlPmXWxJHoAIRMwihA7v5l8eclq5GhujC7YynOr6Cchv
9OGWnGfPA6fDCs9ZT/S2tEKbya8KiIrUOaazU6nPnNTAl2UaNwXisKTu3uWU+bIl
snDLzNUnaw3WgptXPchD2T1k2t4KVLdPEdBzXIs3gavmWFpa0KGOeZgvi0Sh4hcX
dXTsfq9CLjq2dD1TyOta796bnMtXI1z3rR5rWgvja/CVEX/GMX1CcxMzZbIOzegJ
sm41c0cu2fUsW+qpk8ksIr81Y33ze4k8zu8rlNMx16ePwkCd2XMiINzOMX//mJ/y
Q/HuhwBi5HWm+myYfV1IcEGhARTsYFlnlZXe//IM861P5QlAwuUm6MFswW5IiHPt
WmAKLk7/EwnH7cvTkl8BWLsebAq6y/nOOTgdDv1sgxvWdXxu4yQ0ywlHHmd8yA56
jeGFYmehDdQwuqMu6mhg9aTy3slmCkUuNA33oXJ5jqxbDADIMxjrYTv1/fa7rzAD
ANnfu6YhW4NOwAY7UsG/nQU+nVVkJZB1Gxsp63/KNQW1ymkRHb2SFJAJ3De3fMRt
DEBDIE/IDwu+tmABNUABfV61qnM7CeoNUZTsVrs05ida8IASYCorn7756LDkfzOP
f89r7QYeRZhmhtKzQZWTuiaZZhsNxk8qd+iQtymfEx5zH75zTmEo3kf6Wc020WtX
VeZT1B5+Bes+B4ZbaVe9dsWp+fB4lJVhukUhTe5fzzVi13szkRGv4dSAdhZkuGBH
fRfjzd1lYm+KlCIDrY9D6yL1IhPWnaRcRWgq5kUvkcjVTzRLCQ+zpdHc/pQTy+5f
hL+OlPd9xEhB6ChccueT+maIHYQysSqR/PTxJXtT1OA5kYWs2dzI2UxfqOtsbc2C
9kGNJBAyaMTwXG6D8IqjqBYphv6jE4/EBKpmNpd+3gqNHqs7yHFPYEt7Yt/zLEfs
oSGzOTFvlvAR3jADBY7KPJTrEy8suFyUCYvs3SVsF+7lk/J20k8cZ+xmS9DIvWSd
VfYTkHoUVqwi1OHTTY3C1/MqQR41GwSCoND42OvDRUPPm9XlJg041t3CAeXRws+H
+pm65Z3JaWLzusCAsv1X6pt/5OHCojPv5DhVWZXFQe6xnMcfSe9XBWnzWaR22Txv
66fwZoU99keDoyLfOB6pEcDL8vodb8yEmtIU+RqlLIVKCXta9M8aqQ2hhEr/NloB
M/99D7OmdhpsRx6pjTZZW0OD/+Bde+eHnGzs/6uFPFlsok0VV3bWR75fZ5O5qn91
VBKHwMJDR09RLHiZto4QJePfL8nq053TPShuPaXKNWQ3K/zFPuxoBkgFBMiG88+Q
LpyFmkU0EEIWbsS34PPM1R28NxIeRuHwgwe6akyQPn212H65lXD8SpGp+oOTrYT4
XxQjaGubqmukwbcJN+e2hYcceAK5hhEUSlPmllRXg3AJlmXJ0QHGJ0d/D7PYyjfz
lKmNaSK4d6GACZ1rdMgqM4Jwzart4QvTpuowmFAgv5/KiiZDLDIb/Z4OcipekOM+
fIrIWFtGirZM+ciAYcPQHdtUHjGE+pDTcfy1qADuwxIbZDfQQRLOp161Yf9jTbA5
YxyM2sGmTAbGrWzOWwhA5pVnqnSfAeVFTTiLrpOi1yRZ+26GjgQ7Sj1jG0Nn9mJD
ZyIJKFcm8JKyGNimGxBwoqIJl49b2ZrAEq588iPgdCA73K3lYGm9KuTgkP5kizjL
sWiqW3uoq06Gp2vBXd7uzkX28BCAnZH+RIfSUbU1uZBxfJsPq3yW4BZrfUrVHE4v
XJl7v0+3+MNNmwd8eBTK7Evum2EauGdeQ4SsoGZIr7L2t7pfaiXX4kUBI8oNDNSp
M8QPp/53mgNiVdsO6rXbQYIbCGKOm55IyFQI+S76iFrEpiJUdVoaqLbvS4cwgCmj
1pJ/L2Xwt03TlLvmK6e/kMIqKtmRsYCJH1XbIdm31K6d6Jfimux2Gm63DdIrUL76
uqflIfY9wdJk/v+QFfJ/nKqHoJELB4F7W45raZTi+xLS0dvPJFgxyMdWkSeBEg5f
cLNzmBMpSq/rE1ek0ImR1M1X5r6OFs6L0T+E9vk6heyNCDyCLCy+WfeNAxGnODOn
vbHGsMgQr9bBpN9F4VdptB179Pi8mdI+pBAzH5pr0OL25oiS0NNOnImdqiaU0wxE
btu2WNfzck80gNuqnfmxK9LlG6I9rufu+fsqfpyiCkEqRUvtTG/tbFxXHRYpKv5z
Vfqis9YA+PnfuBdo9JHdaLoI5j3lUCMKr90u/Mlqz2Q6HUqOjYPfpgTDDXBtrjiM
hN9GMTC3s6WupE4bdmfhcCKx7diADYj8v9JN3sE2+S7WNiXY55FqFuhBxy36CLAE
aj5PZzGWtDQDtRdGklAYXQhS2hF74iiBG8uLXo/j3jhnoap0iBRx7Qwab8RKIuHB
vCpo6PTpmqFfcDNYwDYNphutllDDcdB/D8cHns1lheS6jpSRnfbqRV6uyDzJ8PcX
LndJ/DZLnm0dnoXQv9J3Xki1ZsX+1ANJv0epQPXQLWW45rMgZiedDn9ZV4T4Q8uq
X7AVKylvLkYOgALLulGKiTzfjA6CRX0laOSckIrotK/vlxa5QN7ebFvglfAy9Yn1
mIW1cdOLGYaIPcJjl3J9bgBT2xuW2kJqrgAeWe9R8LTohESiKA9ZTEhvHC1xxVJ2
US5tA+T0GrQX6yiwNmIsjTtiRXQ09oYdjcir2GOVE0yLt4oJgjE9iMDMqO319g2V
6tcODlSjaG0txY3c8pDaco8VdQpqFiyIfRMLHVgRNqz4wpq1M2asaZRvscx9iggq
4PxBkMw0aOlgqGyLxA578usvn0fRh0vxuSqMNnuucQk58CQZ3XzXbGVdwUWltMOS
nlTrtd8ndedcOKgfwAnTh61oKD7KmyVjZUx0PvVaMBCrzqyFucSVisNScfFncNcw
/F3ubx5REX6rfl052S42RfP2hnGE7dC7BfLxN3z1UzOYlHWlRke9mic6TiMtROx1
IWFScy2/MOcO/X4JRQK3Id55Nxqb+VFmS9/MFswhsul44jjhOccee78CfqdvI0Sm
++/UB3VrLWLv9+zzh3yiYvgikY+wZXfLO7WXuwVsIRaQ6TKx4PXhYpjXDJf5IUp5
TSREuFXVbBLve6At3cWEi5V3Xh8ztECw77L6zKNF8rCxPyq/K2wkMLSdHyy3Dw8e
6smgU/NpIoepx6mMhlx5szbSbuyatXCno5bk33/w8CIbfLfDIb0Xp2Je9hI0chIQ
3rbyC+dNWnjtpLnfzJos51c8bTFtZnUsBK0picC6JvIPJc1+4f+KFRlBv1mxedPo
S+aAJqoUQxnroAKukygNy/1jvvc7xpjVsW92gw1umyFlIWCZe25ZZiZKTBakez7A
C3txk4bro+Q0x2Ftmjexnue3ebT+Gf0RLNfKB2QiAt98lLhw4hczhfYHnYgFZL0s
lT5Bje2WL27KfhR7nSs+mLYIe4uV/p/sD7KZAe1Ono66Apd5RNUo4+3zhSe27W/A
c9gQNy/Ao+FlEC6NhYhQBjUqlEpBH0rRSUW20qyhYE5w8/CUl6EenZ1iCIefQoTb
CaxrktM0zbfFgrGO5j/O2CgtgW+gAHuhkjxtVhab8DZi4ZC+sAtbiBthnvnr2xi5
3IswoWvphOQLru/MeKEo1Olfnee1Kj+UJ76Cs4hEPiIFO5pRDFBdlebx0olNghiC
9T0bmpEHPJxxoCepMbGvoAZXKn0BSHgXffFRfWlVlRvRt64Pb44K4R7c4qcHxgbc
0YDWTeJYzY4Q5kTy4MEuUHYnydwsjeyUH2t1P52qFpdjjrIEYc0mMxXjDb2LPKbN
yPY7qT3Ivr9wMHUVI5f4cGWdHx19YThH01IO14uwpK33+kTdbQvFb5/S0z2byWNw
2YjZRBI/LYSo8Urww2qBk94BSug4PdGL+xDnCrcldlO3EBDkNSGfe5epCQ2N3ov/
ErrFFW5rkFW97X5I+mDiQ8Bo/cArFpI2VoTz+PlUGVUo8A4m5QNLZCLf8mPTuGj4
4iP1n9oAHRv0xk2IhLZRXYrAfCjVjLaf0NJHT0IrHvyd8VZ7OogmyKT4lf/HELcV
ZcqulPDcZ64EWJ4uNwVGLRGqoX7mE0eZCetXVF5bslQp3J4UzRnRAVkY+uhYo+9j
8QKYeXyMLPzEACWs5vCGhDZAsgWkK2pvI1T7DvxlOaSdQ551saJ/rdPvCQoltPH9
zAIznUmDhELi+xNgEyl3gK0K7X3JLviCCL4SOEpzm7AKutq0e7BleGPXS25Fvwqh
Nt19peDoIcqANTalBTEcBq8zW73mbEfDQqGoL6mtxY3J8pb6Utm/hsIPL1LgNZZ1
1kmFqnt5BkhNMQdhfiFJJeLzLkwyyjddIMHkOLLUJMv+jkdXIs2Kw0geujAkC1ia
kh/3dhKBP6itNHU7w1vYNccDF8QuhTEHZ1vcHXUD8sRAu4iMjZCzTeP8W/6olBD/
owrR9+8qSiZeW5yjnmkDJBOOIxufPydOscamxjJPxaLMw0vSyCFvEI+bO4eULmSD
55WrV4rYfDqm8Gy4V7KKQKb2NgfJMlwJo4q87hVyFgsipGpQdmZd6SJAWhP+yvy7
O4MqisN7nDPH/jOW2GLs9lcxhcPrvKdSuK9g5UVjjlS5NPqBeDxuu7JZWkAHLsUC
PQsYQYrXFLOqGL4SD90G0qaXFxruhMuMbzhI2/JKRRdHa+o/lq9hchfXl3J3pkOZ
`protect END_PROTECTED
