`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9oPOJmTf/ZG40nwBfSSJa69RaIdwTt+QKnLfwg08no9JOZJPvm3rUlSi+Wh9CGG
4Q49Bo7X4VOl4mqjogYNUgN7PfOpElubqZa1FS7NJvy+2VRytwjefhF/qctDf3PG
eHwbO/lpJK69KqkGqXv7KdwzUiDTTIVnm+f/nSPrrLBExC9bAcfBOY9jH8/9X7s4
60ni0IJWkANOuF2pns5KHO71/mM+sxqBJccyeRF73mTnZxIiZ5gOdLPkaNvnjL3R
wM3DNmWRA9yHuwriJVZGUWo+hlN181utcoUX7Msnao/vuDXpGSrKBQMtUzKJvFPS
xMOtnUXqn6vvLUBBdOrVqdum42UgWYIkNcH7YW+T87BVLSN1IO3sG8zTLNGvIzQW
lBAfWA6m114Mjk2ylVQvjjSvfqNtklYWyLqlXxp2QkjrDm4g5Me4kTIwhu0EeIMn
AWT5VahJ6u1UE3GjYAw834q27ChDpAYgrgSn6bA1562Pm5TtHS7bAwayM6Tp5Jd7
JkiPG74hT1vQM39DIArOnosAMvuho/bKBSE8UqVvtnbGiBSmPZhbcitY6DOFWeMY
U2YBaFOnETNxefsRSucKSuGXcP23+EJov5v/QxxQhtfMKw20vlkfAIooQ0nLYiHr
iRpIDBtqcuyGTle7XtL3kOdPVLEOnj3eFkcZ9uezhuVIFTsxfo0nOVwfB/aRFb+9
BXd+8cI9B1RrhVA0ErDU4wmpQVJLXJuo7mM3SMov+VK+7r4EmpUv0sxdHYzxbS3J
q5XZlq7SImG/O+Me8S3wIJzV1qsPC6y8Z4E/xoqiJD4WhQ6f3kpW4cjzrXFJSHds
gxQ9WFa1SJvs+cVq7uCgUMwh1uOxO4CBIicIZcCEczaQv7O9Rg1SZNwVAfv4jVtJ
gemIYkxQaXRVj6HugRwdLTcRKOAOA08URlnG8KILSdi8Fpm/7VQG23OHj8ol5k9Z
bDfi8INw26VTvFoXaW+i0xpIr+GDIrxD6g8Vz9oCl8oCvPETRKDpSq43UnaGndyV
Ytf7QOgYbBtdKzAvCM6+Hw==
`protect END_PROTECTED
