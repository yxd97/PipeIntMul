`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ghS0CHGxDLoO0fsG6TZCYtdAFWCGnKzf2zpe7eO85UIS9DPp9+b1+5WvReJBdvq0
7HA/uJ6ywpePTthNY7Wu5heIjvmJow30pxphiJIRZ/AnGxAWpDypWiBwtkXMIl2J
IC5emCs3RhtI3NaAzYmwrC13EKntjRfohXrIq3yr4bfGlbq3/UU8acue5dVEtJu5
/j2X+5+eNvQ1lN6A2Ghw76I2CoEmw3fZUjladtOK4NsS/85opOlOLLuqEa7xxyKb
6Q9LpNZMnLiVZRHbkuo9pZYQbq/VKpzsvpbPQtmW5N5V4kUeMu84b28dh8njxWpr
QgAU84P1rlABvqz17mq2cgLPnxH0uaScEVSZjzLD7jLSRwNZi7E4minAG/xj3NuL
az2L308akNmDHBvKmIk4r5SA+G8IcKBo/YwZfaF4E+V6m5Z9/uz78Mu+ClJ9t1ni
ViDWZIdyQwc6lneTbbN6bw==
`protect END_PROTECTED
