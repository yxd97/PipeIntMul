`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Ju5MS759f6DDJh1YIlVJnpW2K54D5TgiIofWvZbm4hT2Kdap/9aPVXuUmN/6iY7
/7ewOCwwUttxDuiHtiKjV1gce8qWnfsNz6ZgQY5EARv6eKOWewGUKgTKbaG4PDYT
KARfUUlqWsiH9Jz8nC/rpIQHX29XglNnePD0T829fbEncNkKdPp4bdVyb8ukJDRU
GepfwlHCXndpBMpzU3bPosBA30jlt7iu3Og78cPEdW//DyI5HTxNB0WtVN8BHLh6
uXP6g4WNJiXuRr7SkWpX60L4k0L5hiO2EIaDQThEeyQ=
`protect END_PROTECTED
