`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5v2dX7E1tWXtY7VYRuSqaW1bb5nGf2r//9hombvnuJ099BQzb4l6DZfuCHptCDZB
3p57gFLnpCVAmpCcLNs88flZPMY+sT8sgYYYq2Xc5CzmDW+we5Vmm6cAWi+8hH5e
kwIi8XX0kbWtG41/loOHGyrQ3TqCU3Bk1B5FHObG9BFQK+ZqU0roRRpHAS12vB1X
dHpkK3guef7KBLaD+tU42oUjjZv/HBhUVyD52jXE5AVmafeNrIKoLY5ZjJQGHZ7x
dICw0EylES7oR+GC5z4+whKQBDtK8+HlNXv2DkNMuAe1yq/YIxXTixs4uq5eybyL
Mk2lPnb6OBM1YAbUPw/Y47zCXlpaxyz9ev5AFjkv9yvqY7RTKUsfbdECrELriWJI
DlRLow87HMrpEpIaaojmIptE5t553NsJFn9XapTfJkSS7V7QTBDb516fdWIWsbba
gciTZuKTWCTPyPK/Z95K267mP63DXqkcKfgyrBPHsZaehCc2ABo5uEgB/JKM4hrR
BaPDZpOa/R8miNtbLvILs6+PDlKGIu6KXvnHHekzF0TE1EABKhtIMz2biK9KG+l5
r8+OYZ9Mk2Ne637Djr0nhCkATVINWoB0H90lafqhJltIlVHttvd31eXqxcUyeCII
3yYZpv+GbEPWIl7yPW1nNJY/kpfMQIRB5OItoFhKxHEMmZWJTSy9qC6+f6tmEBSz
HhlqKX4+xmBign2nTyZMJtbmtnhF/JCiKJesJlVqIf+lO8H2eexPy4XBVXOfYAq1
UMfI6/n6Mb+s1ULPQzJRlNpiz5U08iosevoYyuAduKWIxg2Vzwejt0njDdAKOVSt
Vl3ouCMNuBtwL5TYVPWVc/aJ1ni2hi1D0KK72zqDl2ttw87UX0wN18Qt2OfEIpgI
4jskrRm6RRBGw/IKeg5Elt+KlBtV7ic1puGEeHylj6fq5rhi7TZNteIMMYbuSApU
jhWVoShhnWNo0r9+0JruUSpoiOPfNRvN8/W5ETPV8iQ=
`protect END_PROTECTED
