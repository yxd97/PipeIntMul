`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHb9kD9XL8UUzcekZjLlEkALmxpS1uP3j3jw7wPJinwtxpV05oORCDVMcV6mjtm3
dEtVTlmhP8fsL/chDP3OZQokQ3E0AnjpdkRTtVLI4Ddl5DMOB34dWxrpsRogUGww
HBSAqUFFLX07nqjdpghm4rR54tLEjBKC/gfXU5DxPxRaQyfLPdoJN08WlAVYOF9E
ygj99yIiX/DE1E3KmRK59mmE5wtMXNeSaejaKMm6aRAYrWRW9WRnKQpIuF7PeM5r
7tGeC1RpJkJK7i/1jGMgL7paqN1zpgri7QmRcs4qqt+k7xTgIEceDEFb21UPXxMB
StbHeH4cOFi4i+YUR5XG1JZiZVCTK/EssWRYQ6/wj6Z+lH2nefqqh8U2vGAm/OCL
F0YyxAdnhHpCEWbkQvxxggVdv/BGSAc+pSdH2TjxEbhu+K04AEzFe2cdpdRR9v2z
G+Pk3F18URaW/TtqfRbMbAIZ9zKwDlqdln+gQay3xB7A8qIQSMqMWx/aPLo1U5Ym
/Y3x7LcOLQC8Q9AtacG2XncPqx9rO8d1i4OaFsIwXuBRQffEMij9wS3XMJOKYbbx
GDUno7K252uN+87bwBOtSp57fwMXOUMbq9HJ7mnfK0akkFHSWhP/8FArHTnPbwg0
WxhKfSwL6VGUA7LLPlQEakQOx0KVvhihd7exKesm2Qv7xDNpbVHEUPSr/QuEjPwG
iafck898fPjGX3KM1HO5bRW7196gVdaHwVSQ/vA3gkunN3v+dgqn8XJ7f1XERTWO
WR3Uk5dolDcuo1quvxIwD6lKTi6FOCdnpzrjCCjCOSQ4lFBr3KvUvDe1Fns9hxV3
XS+xKiplYilky5i6Sm9AEItjBXvK6j6esrfq+2Ue5wvI+7BLKOAFkdA6iitszwb8
8UX3vLisDYhpc+qTX5XyyZBQLckfkK8u8frJvx5Qp2QANndlaV6PZbZt3/SMwmOM
NesuPk7iqqNELhny7yDN07j3X2YsI3fpQ1387UawzeSrC2QuHDEk4L02KlgNmfps
AvmgS84kL9xgLpR86ncN/D1IZb0oke64IJnUv/3a0YRvFC4JQV5rKoX9zvOdwRg9
3VaWcGWSe/BdHQ4tB/r6YGWWcqMxwX/mfiAH8UHc5u6RSsVrPK5dOuENqtD9kO0o
wSsOCchEbsKNtcqOGq/7vTFm7OpfvPCNDV1FetTPe3So3KeKqx2pv8YGalqZqI1H
JQdluNW4StosV4LF5yV9e/ZA0Dn31D6Zh+YZ5jWTDDRfCp7Oqt/k+hlRktJV879X
WOQ0G4MVit1uG8Fy4J+vfdB9ANZa9oUaV2zs9LecQB+jLLsY5H0t48NxTAakaPP3
fEOUWrotz1J74DoEC9ouFz78EUrMYlseIyh3x6S8Zo5gjdqH0xY5Za98sH4Csg9c
CRAOrv5TzNidWIbK9SAC1AwODtF0hYHbPhC5lhXVRdypibIp2RlwgHv8an6PRira
nESuvTKx0A9RF1sGPlQTGTGeLOx6vggmnVsJhT0gjg1aI8rUo/SevEsfRshmZpaw
qP5n8tmJyuoLfa/8NNG/IvNoxBwZsbCY87XFWa3UQlDm1nRQf48pffCKMRIroxrE
iuquayb9Hvkfir99dVvn8R3yS7oGoaTBwiSo6DxkHIwtOlVUR7zJb2z7PhFMgGVA
LNsgE46yARe5+AU8pNk95CSAXghnUCgjkO2MpcypUDB3OtQgsct5HYMZvnOde505
RAcceOgMPIAiDzDesgCOBQaKla18411Uy94XzV27IYRxCtQBrnFo5ukpOIWzDqnf
XZXljWKPe07+JL/Y2tmXPo+OgdOyVUWVG+D+g7pA+AocagCyymjK2ZqFK2n8gSzH
XeuL0BjZ+I3+pbR4HdY7bz3PABHf3EA0JxRfFwdG6PdMQTUOHbZkTu69cmr/AJbG
/29gEmxCZLaMU0YQh7+hViy4d7FGU8izc66mXSqcq+BeliZLr6TKCaA4uxlGUO/S
0VDDmBijvPjnzwDxIZNuycBVg0UPs/Fn2qjx/7dBJgKqDxLQMVFyvfKgMDkfNEvp
T435UB8PnubIsFMyHr83b/92kBXKe9s7HpwswwOsbpoFTKf4islODWKyyYv7CZdU
4+S/R8GNLLAYTOq63aj5PsZahV8zfbtiGEiSm1c9eMd5Ifu5RsNnECQGL/gosg2Z
M9vQqt81Vlcu8LweBxFBuegtULNKSGAHyzliAz/6Omelsq2Ik/jjR9SAQvJpaS5M
5Kb1s3RqLcd8SX7mvojgiA==
`protect END_PROTECTED
