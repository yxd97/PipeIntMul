`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+FNQndeb4yHDqfCgiHfacrfKJbzI25fnXQoPcdCOFC0iV8TSynqmHFwfYQn6/EV
TV4G2YAjFB/qLRA6uGU7D6mL8i1+qFKgMCMEs7HrqZBGoMZcQ7SKeqKXFqeBgSSR
2y9JCQk0Vat1NPdhcSiPbqu1EiTK0n4Ye3KspOYQrqvs3U3YkXoHMbH4XsoIHAwN
5vXhJaSkNSoSCrm+5NZPjq2uge6alhdxu1PhGl7QKQkogHeJMiwM8WZQBKgjV8Fb
ZqzvpRJ1TFBLZlvEzbn3spXKyc2Nj0jm/6lGrpWe82sgM9VC4HSpx/ZhLG9De2of
pLVu8rEssOk5jNlAZvDuy6HJT8gK/gvoURLXDpZIiQXmabODkieIXswXV4+iV/qD
hFT+4iCBsUMHEgxi3VbWgHnhfmNsiyUwUJ4uDgobOReoYyWNodvVqyDKQqgFHvD/
nMKAF25io4ehR/DqKEEgsbaXPBhVHgbiaA8qjFgjTVs=
`protect END_PROTECTED
