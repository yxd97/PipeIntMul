`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKZ4tUNXIWjTIxbKv8xRscYofYBUIO6APjJYs7VE2yzH4yl3qjv6RFAcnp4XGqzN
Plxmt94BGAqkb7vLpkdUk+VtLEWJrCuarVHWloNSUCDc+OReF4ID+uXxXUAK6m8r
8f3N9WvzlyxsUMrnZzxc271/hL5swUOq5c2rxhwh/pPj4l+InyUBbSsSCTkigcWc
D/Q9RL+U/7nbl5m7n45Ojsd4SLUAUdp84Ux65v2/EuOr6NOQK0+07uvBUNCCiOU4
tiYrJvLLC9hURT+bYQhXRF8S/6tio3L23AtmwjmB7tMpg6lzm//jzmvQEPotQKNk
kaumI16xOa95f8GBNRCQHnsPwfsvwMnkxhiPNjQ9+toSk0SiccKwGiPnEKzWZWUT
088da7DBOjHrw7ZrjEjUgfxQs96qAUBBAdNbH9kx/9UiGJRTGQSEmPCzqfdqcz6y
hDJvao37XDPhM+YpuOS9xC8UocZ4fFiPwwDnn46ng3BGUvJWEoNy6HitDbZgL7p5
flJalfz93XJC+lruL4y/3wi/vmWuB63IZ2tVnaDsAEYVsRVQbDrCeOe+Qav1HZe7
tFTwiQ323UOEtgL9rSjpUVcFnEMddLy5o4dMTDv5jhEZTP5vBMkSNz8ITpeXYcgE
vxhTi2R6h5rai1+mBjCS9IiL/4nCz+bNDvWKhjEwce6YjyThof+C50Zzany7UVcj
vNLcPbfgQVjRQPugAA+e2I/GnJ2GARl8+GA38CFF73OEuLWn1kEXrL9fR6JjF1xe
Mp1E87OdPZWQvn/pm/kamXgQ3mNSa57KD7a4YvqaWrjJq0jEnlutRM/vbEtGi1tS
SOyUqtsZB80FyQ/TtXCuXoALu0+IPsy1to5wgCxGKJsF+jqDyX9H8pvTzV0UL/gS
nbS9W25O83vybOpc1yKVvkOtzoWZ+UJmABvNm6oIPdxzbEnQJPIki/Pst/bnzrWA
Yyou7zJvkdHRFO8QZ/63UL4pAoM2tIu/ldvBd1Ao5jf3M67kW/w7oNFcthYCJF+a
L9JPdpCRTfQsE0BXs9NnBA0YwC6WYI/1vOG1nshyFGkxtkw9Qb2tcwAZ9t2BJvlQ
lBD9TDWeBLSZhFMCgNdZVkGCuGO0KEQPxMtP5nyoSEImSIkUfp2b4J4pA46e6swZ
elG/5MgEgUnfBrUMx/p492pEO+xBFAXziMWUY4SuuyJb4G3YLUA2CwOvKuX0ZS3F
7LhrtutXrElhrsGG+mwusmS2qWFud0yoDgjcPWMORLdTbUbWqWy9obGky59gqrwj
rsR6Y7Xi0t2XLbyhEYGqMijktEe7ga/fe4HlbjUIiZQhqVulAaBMRXuJxuGy2UeB
rmXS/GfGo3hq6ytcdg932Eo+XQt3IQH1cyxTgUTqhUQdYuLNlqLIwwuMBskBNuRN
i4bp4vFkXqWLTkfazdhntcDJf3v5hW018HVrD4nqNQjpVm65tFqmQKs2ikbaCnA+
ZZ30bx1jXDin85BRuihsX1rvdaFNzd8uamxiJgENmn995+swpXsSzam5xZIUMpb4
k5wJHJZvQGae4yNjwX8GE+nbSBvcvt4of9EipCYUZdiFS3AaZCsKedR14FHY4G7t
lHeduk5A5gF7cvUKReayU9rNItW9KuvRqsVkzTfCPD1qGTKXecCZtRXqd2ca6CxE
tZFTjIkOXiN+vp1e8cz8/RQ/j2T+fUuEQH53drCwuEkbGKqm+K8TgQ86gErhPeJ1
J/w7TbrbrWJaGa1yrggvTHRrTcLXQAcQpXaWGiEQzVMm4zWnwUke5YSATZ1qsFeu
T9YbDAXAau3Mjue9CwE1atGWWjU+cKvNn004BGh4bEkctwLYQ0XS9+45X3L12EEf
z4+Z0N0Rpxz/6AXcwF5B5Kmmw05MRm99chU5QL7Z9qm3o0J7v2LRA2ztuLFwykkP
1vc0/INYmhjNp3RjlX3a2UIIRi2Lp6543WoS6d6W9RcxU2wGNfcU0a2kqTd2CE3n
BVXZcXihBskFaGoeCjgCGxQg/QrztU/e/nOrU2Ha4IYHYEcwXfyZAzbZGOghZGex
3WeN3Mc50yTAtWvWbvzo+al52FkZl2wV6gMU11UWHtzkjeX7iXWI8hQZsAJoXHFS
rf3V1C4YwmKyY1zy5dRmZtVDVBYYLpiM7QRDClUpNp42/6MLhyabJrluSyqr1GxU
ws5A8c0hX0aNR1SV6OrIzNCPGT1tVdr+xr/teqb9OelihniHDvhJzyaXXn1BABl6
r/dZg1WJQC7g2Jd8eKAF+SwwkyCkmdKfwN9hAFzOe/Jj/eJGsCapctVU0hIc6IX0
Gq9/3NXyuWhcGfkAGW7R3J3KzLrAgyDetHKIwwKXDEaHJt3HPkc8Fn6Cbb2d48nT
qEHd1QC2pwk4JznRAcrGALYJvKwyqTgDtWeM55XRxVrFmxqJ1ahPnnYIR4HfR6Ql
D93R9sRFjrLdWat4coi71Jjaw6qZnbHGHsoFXo2u1R+Xhymn0XSDUbQpOe66j/2S
EXSBE15Cevi/9iAGPidqK3GWzF9PPAKfQyEpGjhFyzALMv+402NU82uQeruPtwJv
b9W+FlO+7J17rLNTIRHfCBzFus4q4Tt+MDeaigZz0IsnmaC3pKFt7BhnWbP8vxfr
ytvVNV4XgmyCbkUZb80cDj570k+9Ut/3bS6CwrAbM9o/Er5G+k9VZcFsWehNdWif
G6iImyiMRx8E2t/bp5oCfXkSZZwoOmeCVbZy/GV8Lg8x082km6XrME+0AGDNMu3q
Fcqy7T+bHFO2s6tfEiM1RDnDCGKRnU1KH3cY+ILss8QpVDt4T0YMD8zf9MVT2Z8r
/9rtA9377VQHcwTR/68c4uJXFYsL+bC9ziGOrgRDTHZNzpa8zaU9Au/GJj7fjhZo
RhheiDfZ1bNGjfbzjlWtZFmmviWERKZ33mtlEmF5hI5WYKKbz9Xqz2NYNDH9bmmR
d/dFDFMKhGaFkk1AoOOwTVpbfMojd1iRAMdrLE+1lC56+ftdludgIYjh34hiWzs0
68YM7bM+abAyi1VyDj6cDnWtFUmi24A7nrBKs6LomjA8doiTMY3FdoP7aI53E2pZ
uKO+/fETJOx2+/S05cq9nTf3EohqBYUVY8a2EaQcKg7JeuPoj9eMIsvqKuer4bjA
T5ZItzkuRTCZ1AdEd0cwkTzyY8dSJugHvvb9P17vpyiRvj6qM40Pvv8EbHhvmtYT
OF589ouQNgy48EHVe8zn8Ah6MKCwQb1Xu5GGJ/KaEBt/vnYopDdxKDQowZn/WHBf
Ic7IBiS2Tnrj0bhNQmRUH/p0n4YzIJcWK6a378NPYg+t49CkDTQimg0BJDZbHcmM
9D8h9Iml7olGeA2cEoyREBRCb/1udxNQfF0KwbpE/qFYGn1aP7aqBOXVykBgaqKc
VAAMnmiOIyi6xqlIih4jsR6tdyb1YmDBenN9FfriBn5LLMMw8Fd/x4sUTS7V2LFe
sisKscFg8zIhT7AUg7YucZuN3h25AafobBCPZA+mO9z1BFyuqQSzivRWbp/Kk2nU
Dvxw5hZAHjKMRdQq0Ec7USEuamSTpdGIl0GX8kObF9e5GsjAVaB8QvsoQ8wZwLv6
WCgI2UGoUVtIpsWTBDSis90anXswnOmSPrn1xzROnTnpYg1CxvzY7ZUWf7wlNfLj
P7JY/8lKdBFpgTM146pn7ii+2ayDUmOu2miSFa2gh4bYc69dINmKdJ3ubvx7VySg
LHpC5T6IJDpEx6p03/wBOKm1wDyn6TfwnxyVqHKA2rndSWKXB1CDzsC/0S2ALffK
ncAbNDCnTOPv6ZnnNhcG3HsBEYHWXHcYZMl5+KSGgUcVEB/79dHIiKur4OJlajUb
gAn4w8vDOGqkaR9KkYoZIdNHEMsSSBU0Rt5PqIl0bhqFGR1xR6ffhuiiKDlfPvQS
E+RLTVYXZy/xRoAb0gNVBEiaEVjjt84Akivf0fUhxw7M5via5pw7N42/1wD+KqBK
H+JUvmD5aeuZX0bAbM2Pasg9drwTkvmt4SPAgaEJS8OBKmoWvavDlxj433A4hW3N
nMLzNNcppnemQfXYXMJWoitziYtgPlRYDS+f2NfUAZ1GTyfD1IVFUPYCKucLoevc
30GxlTmKKgJtZh8IUs7ZG8YH5iCthfHrk8o9fmXHWguIVzSPejn3ZnJQl/X5QiHa
jiEwQin0T5DLEJSEzAYdN2nIbLmfZG5YGN7+5jhmB9KR4HqQsrLjIB2Sl2lLFoUW
DXunLE0P74dkMAbV5uJmspaaOa8d8FqCEg8E4kCgVp7UzJxT0Eu5zQCg/HMFdG81
4qziovwkjpjYxhJYJKdVGPMm7AwYFsCsO9kmqh0M4wTjljjdFHANK07KE9p/enw5
GwqrA8GIv5ETk1+VSC5yDhn+hCFwOAFePROr1h9vJON+zFg70dRyPzLRpYPCIJ8/
99RDv+Tb4jm+wELkt3l4zjUzeRsH3A0ZejiUm52Q59rg8reYLB4BaVWvTuqtDC4i
+d5hLt3OovqfprSgV2Fcz1qYMOqiyoCwPtpn58bgPs2TkQEtthJZIF5KSJaTUuCG
4OuWtGIDGSoiiMtJfpMqMG7n6Xc++AWHv2xeb9JdzrNbmJ3Fy+RLldABilQILG0p
ZcB3Oc+epFkM8F//vesZ0OMmzy6lbXYEjMJdxzdRFBpSolygNuB2BQTINCwwAoXV
k1ft4/03ghAD1KIatAb7YJflHdibb9tZFLPRa5aXPTh1Y5dAZoGA5X/WizgKlIoE
UQIytYyua6i0zIftQQoQUQdfz10aIZAgzc6JzTtyelGmTSIFnWWM+GbODqAK1TPh
uSS0av9GrIaOKekDioHBxQR4w0tWSPAyunLDJFXuUMD3tXpHloU4PfxURrtvl/Rt
qQbQwgQtxlMBfPN3T/4+Jbm4GnDMCJtQEtqiBkeIUprHzXglr7Gl1m6moCBT8QfL
AxkrERp7zcuWf51Y/xyXuNkMJPz/s+dVop0fiCcx8sFyF3AktCbqpC31QUU8AaRJ
DqcWKah6P5HXxaiMOaqyJDHPLLHH37IuCknDdBk5MLAVuJ/xQapjH6t9h0zCGwaE
7eONKVvWTBDQqN/yi5AuxE8LhU+vwHseHRF3Oht/sW5vx6rKiRI2w8sVzm/AyITq
JCxqvcOi1CPutom/oQwrAC5Sxrp4EjxH1TLFWOlReHA+FAIl0u0LCNgezii/4a7J
AsUXUSlJ8APvoITRaaSpVoMKeGHGGbtkyChjjPXfuxPO9DnoAB745U1IriAEIAS+
+xrBTY19Pc1hvB+DxMKS6lxzEJeyFIMQnUA939Nu80XaXrzPC3Pm/pTLm+shgD7k
kOBW1jbwj70iLxx4W8Xsr82up91TYrsVYhIqQ97UmSzntBanIFirjtI0hfW704HY
Huho6HkyOB/xMwm3Lz5sboLW+z52CP5BGf9zhC/91rgNlRkZOw9Y8cftPcF2lRow
pvPZgjyyXo6fCKNqfasDIKjyOT1eXHWqQ8cpGn/v+Shl5WQkhtGiVdwg5EB/tCuC
RAO6ucPhfa5V2MAYGBTA/GyBuf1lpxHBnrbCwzVshX5Zw59v+6YYlrj5hAV99ibe
4aM+XrK+qVgqqetRmjARFbclC3S1QTT2+z0m78XDqtFMcfBPQWohaxaZ1GSb3mBL
ApPdmeRaIwjVD5bxakcVx6MUxWOfWzPiU5Gx0N5azDlBKrntdeH1gn0OeC/ugw2i
/5rSlzpfNZSzZRgX6C6qlZJ595IxETfLH7YMn6UiJLxhaSVzlAVZz8iM10AGUZoM
d3s3rhrFqOJInG4Qj2JmaRsVcK2vmcfJuJTAAffErZOC1w1yUsm1Z+OKQScx8aHE
wqGpgkDMw+r3ubb8acWruzwvnpBgr2aOPptnrGpupZnsK2y8WEOLFLHUEOyvDUU2
fl2RdE6SkjridUGAKVaf/iExomX7+KgcX7cwg+HGxZaNkV5sc7qM7HmcYMNjuuYM
Z1LXuNGkPDlzFExJrBlFRN8LWbAKQchYxr8qQWArYPNH0OosPYGfQmjFID027Ti0
KWsH++TcHoSDha8UELRyFzyMDp/TaEgQQO5X4RYQFndgPkB2/pys4pdZ1ahQ4JIy
xoKg/4Smir/D4m7+cquGKavq4x6ulndpl9sAgi64XRdBIudrA2Jjh2FMFPU9uhxy
/hrWt+9Fq3R4AMEyCoRbWjFM271XKScrbHNuKBPqdpRsH5DGI8CuJrInfQAyFmJu
XuEvtR5bSIVaqKSZJjm43lR7ZKfzK73CNepBWAtVVh+GrN0seLl0sJo6NtrkfGMr
7VAex+ja78i3ZTR6u/HaZX28ulf+6TOgo9vpGQxrcN+R6r/lhX/t3IqXmYl1118g
Kt3n/BiE0ZnsyeYov/oqOW3oCBvtL3ffG8qxv28P6nuGNzWPihwxBXmmO1h59Jg6
L/Cl9cUElcQBYBTTYZpo4oRcesslqGCYmhTODnhp9c65dD0wAw6RNZx2ft25ja38
DMcPlmWMTpvemkiE1QM+sqF9ErxH+pPcDRQ4erAfOyxwvaO3IprQuqHjCrwxWvOP
mD0/GRJwE8gpGzFb8i3u687HE1/PkqtukvNmg67vcWkmLJuSSpU1KOZ5NJluk1eX
Xz4mwKIRXguDqtZlt9y624ZjjdjeSMm6KOi/85cjIolGTQjKi81WbW0qw+aU2RCn
aOHDHVTK35WDr5GJMny0UmdjSZrLP7KHhS1j8QvpoDr6hXTeIoYWEkqy3wiFYvzV
aUpfkUc6bq+b2sSmYx9VQMg5l53auGVzsXvNyYFMdBw9F0D93sE9RCtU/PIVMOsm
MTbmzc8bdp8MjnsmoVYq8d+PzHayfKcTwlFNZ4AR8XdfaieXACMeiSvb4InK145m
np+OpyxjZ6nXxF8w4CioY8MyW+ksjQ/N4FIeszT7LUKD3nZB1C8Lds/y2fi+ow9/
A8+vHVIwWIyH7N+NmG0X+4BgOaPR2BhbAMHJXkqePCaE7nGvCLs3Wtm3jAyixJ8a
O1bcC1SSMsyvZ4ZOH3M3+BrLqbP+QOkWXpkms9LMIV+GwkxCISEgZgh3Ty5ulxsJ
Nhgiv2Z8Bu2tgNJ6NMrHX6Tv3RBEjBFcN2XGWXqb6vdNkpQgno3MNyhL3IEp5t7v
lyIIep6hG/cpKVf80t1qpLboR9kjQPmcVP4dUd4VBDc1MlH05ODQIzHc3gv7buvI
SyFoCC7KS4YIkiUlGTK8GsdXyuHZL/jGq4bLshYuylFMX5IqTK9AAjCIcM6RKUhg
E/DlL2sIDFyzPlk98xlKQLi/lLvh4QucMeTl95YRQvnqMbjnL9a+lWP2913TFZOI
jlcXS867YDI1+cmmUBtNwqTEhElV05Z/1ed7YPFZP9vunfBuS1rkwqgCf6sxxIfw
wN8z6/2C+GAfiSvI2/CGcoa1J4YsiAdIPPbWGemCfQkRL5IwuoTDLnppkhT90TDG
EQVBsg5WDr/Um0RcHGUomujNuNBeBFpKwmgEjeTkRRi5xXhs4Q/RWLYjJjg0gWID
BkbeqcLo2I5NcT2NeCBV7F8z3DpOVn8k1TFgqwOU6dBzP61gHO3udgJlikT/iyfT
ZOTSSF5ywHIXEyP3tmDBGpLCC2gXRpL/UMGYQ0uQCpodUDNk4qbR9AZcbNO5UJMU
TftXWIEYsk7MIKxSBxm3n/0AYo9nsU68BbBBiscXrlKLv+LcJTKWmp9XKf3VZJq1
HgKm6Y8RR2i3DQAhB0DHnC5qPadeZMZqQIsQPkpksFTBnJLq96+rHbamzi7tvV+d
wX44m9W2vJ6q7YX+3fRXFS6LUOxAueseehi9vTofhR5BD8gUheP0a5w3CFGO3cdx
uGhcqGKOXfx+vvaBhmV5RaxR0xXfJmuvJbeij/ORWetP7ECcEfI4VAfBpCM9RaGI
Wc1EaqH70+rw0sabMcfbPDDolsUw244GFfctBBOlIgPadl/WqyjlXMMgkk4y9OOO
weX61cd5EL+feK7w+f8tOGKz8jr1TCospnY8NLk0aIQknDfAmoKgXTx9BtndrAxY
d/CVowqkKX8FFtaxO1EU8dkEY/y1y0XqjH+Lt97jxlGVLxJSRQdOgi5ZbY7pulOh
gz8NUASrC2ktIVTVHbbEYilvmPFU6N7S7+ZyXn4zCgSFVS7qwNPWy+sWihT8LW/d
nej0tpulsUylPCh1X7B8FV+1Nh2G+c10RC5cGgq83hyWFLn5khEC5AkQ4UepLNj1
98Z8kKvmQyZUF5UTq4ZxWFd73HCnlCWy3SECR0Esm+GKp5sCEkcHK57dwDnGyyyw
o8S/q8Kx0CPq3NTZWpZGni+s15/YX4cOlKHCREHl6hrxI3jSYfQ+to/pduMHzU9W
Ml8JfmNq5Tw6IGvUX7Z0GZU83H/Aq8PyffwcHujc/hneAFQem2ZL6+eyf5ZLVe9c
UbPvrZ0rUbpQ5pb6t5od8mZ8IBjPIQqEmFvoPCUiOi8fmb/v5rf3NsawjdwIPSAO
zt2BStKkLgdGF1q12OoSi9dcwrAuzYjD655daDLi2aJUtc97M81/hvZxcGluguDL
DZC+vKFlLvo58l9uDmaKNcYtU5K71xzHnzz8TvyDDHF6arL4cb0Wsrtaj9xXZXzT
v3Y3+ErffpArL5j93QHc/xZLuqAeLUu7R0LwWbIFgMOA03qpita7VhjS8812WtT/
IsEzDKQXp2gVN50ZRbMm7uI1UmP4xGsqSTQFhUUzHDqwirSr7zNt7dx31vwfpTOb
jxqN+jeJkniLR69SZ7MXLuaSwBdMxXpqBDwnNwAnSB6szvYaV9b4bsAbhzv8pMK7
0gaHXyUv+u7XUUO3tK95EQRWr5eeeXQ5BTbxd90DETJxmj8uXvbPJRgdLgy5qIeP
jdWID4LogJ6JPoF2IyB+5i7Uhm9S4JlIDp+umMKqZ9zZUYG0fRR8lcsyF/9J3Y7F
mSY1fXPaL9ppOuxYexEQdxGovmiOiEKk3IBs4e9uH3YfgmZCdYbk+aLNglDEXsvo
jzaaRbTH/3DzGG9l0WSSyUaOL5PecUmH6+jZz3QS7Jl0hbhWZIcfq/zqE2D9yKo5
wO8/3wr9HGKp67qmkUeu6/3/bGa9A1PgbKQxCkdmYuwAUa6cLBWBh/gLws8/aCaA
2Hks+rpo9SpOunbkehYJ2A6LzH7eKXoF38lSk0w94Z7z7PvVE/2AnYGTexXjpjqG
dn+2y4CNd8eTyGaWvdRzqWpj7tobBPASk8Vb1mL8mts/BuhaobhwFs8RCKjIqr0B
HuOU7orhVX92AIuXGgvCivDWDJJbXZKVp4j9qwrI1/pnfC97z6AL/86vZkReZH4p
c8BNE1JBjV6SC3KHZjfRi6vjrzDgl7bw1Dhpe08vqzlWCfbxiUvVyrk6fdZ3L115
PUxOsaiHZkq6S81HBC/JuWDWrg3OmZrtgzUlLykqVtf/841WNFdMBi+08BcMchVQ
mfCV6VhY1i9jeRdTLkC+5v/okufMarb0WkPuhg6Z7+orhFHaqeOk/WIq9CP4q3ka
MFZgNNBQ+slwbw2EUIEQi9uJJdzGullnhrWaOJ+gvACnQvlK++JD8UbgbQkInMjb
hWQK0GkFdylYBDl6D94Coh/FRib95vlLChOBz91ikO48sWkhduHEvYn3zAa2qJbR
zGvWrNrLGaDgYgGmlfzVdY3Bwn7vOz7FnXlvDEYKNkHD5eYoobUq5IGO3zaHmYii
02aYstxFYgajuKap+vBn8CYCkTu8YSeJWFA0P6eON3ygVfZZkFymK1qvHHI3GNs5
Wo3RmYSHb3A6iJ++KksljdSoLCSitGzU8iQM3HEXO53ToCE/Cxr9zgs6mN7EDZ7V
6bKZgp2Iu2wfOWPs6fDUidANXxV6EsSUsu1P/avRhxCnLlpu1IhF7dLMiM804t9r
1MZD3MEQjlPkpL0bsTkvqZ9gpct73WsUiRQulbizNVSG9UnqGX5mDfE0bEJ+uM5t
BflaNdYezuVQFSCW/Rg1mEEcUSfGuhwJXXkEc1h9aWz3+OzBZrtjOqfLyv0Et4EU
fJbRFJCCytYARkkUPtrMRRPlFIjvbcup7dNZxZWPET83wD5KYw1LIYE31ZqkgfdF
IMkqa691XJEVZIHO+UuVRaS9tqO9j33V6p7TyfuZrZD8rKUKQte1MNut6bnJGWhh
yxDcs6I1gkVQYSaGGmnUZrFuyVyMi92egoQjVr0RM92yaOdeXkM/CFYr1bHsDiy5
S8vSK3iUsKJN0uhVkqWujXhOYfTdTzsf9XRxr5VBy7gUBHVWcwAyLTsWuJSmnb2R
dv/y1aJ20S6bSGQWx39hnUrZX87SavjbIRqjQCw5ke8v+MrP9kWGIwZKpx6bVQ4v
dSTmlq6wylVymplryMflztpBX276/KenD3+jAe/x8yqoOdAMFoibVu4c+zp1b0OK
1gGcijJ50UDnSPVf/8/dI5PaWZDR+3b5sJre/Uo/uVkj5JKq7FQw6kYL9HoY5rc1
IMbl3m4e2drfvmzCq6Z/Qxtt4XazgBCg4V79Ux/IIH31IA4ufiVm/P/cuX0vlK2l
HUAEmysCJDSln9V0tc5wSDXicQtBjnnR5Ms2MtN6U1+CIwFopyM86BxeW05V9xuK
rFfOVr2EBlx/UWNTyig8YeEp5F8Y3SKFXFZTfr581V2k4uwIPzr5CmTBWhfNVi36
ZUlCc+X/45H6MCHcl7ETJUqGLmbd9IbP/93LvdlLFSBPzoaBkePw25owu/bL5F3Q
YjF8OK8s+mZ3N30el+JMZMljE9COll1E8zrI6oP55MUvq2iGbD/GnuigsLf+Yd3U
zTUNQhtx3kayZs+SijxmMezEMgMMYSo/nhf/RfwwxXvVWnybEQj1M6OQkrbZMrpP
maL2nYec0Ay7b/KyyRLAgeYkL+puFZ03nCC1FPOfrecx5M3KQZ8vG2T4NqL+M1kY
VKKwP6Dkna6ea7Ly4gDIQqbW/KxPZXZ4aakGtM1S8qsES/hmjEjz5l9d05wkOnFL
nCPzn2f9L4fIgZrMFKkM+80RIrlwORgUgZawySCeavq+qnnKfSNKGLbzKqT2G+lO
o9tagX+nwzTroDVA2fxY4516Ev1HJcduq8cR1Gnu5BRjmkbyrZat4OvA5qFWY2t8
Tz/tj+DeqGNHpxv63RA2IzreLxl8YRdGh4xnPUgjVs0h7SMByBrJBcYWVHNlX7BU
LTt8ek/F0GF9+wd5revtLaeO+Re6iTgTLw5LUI304iASZVqzqC6v6rkgm4EbrKAH
713P9QUw874JwTE4CDhnMyKSNWFDY+XjlvTKEvbxEArR4TqECjShr+aHBfZODkm8
gFBvZXuAseNP0S30bV2sGOoiyCHRRg41yFt3GZdZdZB3LTC4XC2E00xqrJhtRWuy
B+o1kqbAJBR1iEVdTlCB+rEip509q6/ye8Md6PlWecCvyMTlKDmAPFCB0rs+RnB1
DfYhzojr1f2aC9JbiYa25M2redqM9QnLFGLuRtw3nfa4LeusABtBtnT9+KUbAwna
29BPGs0YM4MfJ5aJeTK97rSoWAWXUyvX+Oixu1RAujeEWJOHCC7SZoBDY94nDQAS
rWbOPw5BgrMGDVw0hVARh4tE0YWK0uVxFEgl0l10rupoaHKoMrv9/ujvrCRV6fqz
GvSQn7dv1yU1yRgj/UufWWwZvyoqDTmCnKjPK62MupbYeXiGNbeC4lHKVddcPBU6
NHY+epnaSQfT+Iimyp0PGIgHL1JdgNZhJszm4NAg5SRdpT12gXLUMrdv5p128tGS
NGnOaoqCfXF4IMkICun8nIzc0eiF2IlEDvE7ciQBKCkCrfvSfpgh32oKAflw9vUX
UvPOefodYbR/WQ6WKWqyy9Hv3g3SkelJhNwctWBrga/ZQGXhpAuB06KNdi46rW5p
XpCfLbP/7aBTxW40urYhEeENS7Ib/CJg1id3ts8RFJmG7wvAF/X7g04tJJz6AfPL
+bboNi29ObfpnwsZkmzVH1ZfxGIDR2T1fpARStvW3b+n9PDre2ImyHXuxMBY4nrI
34PIBBmtHKKL/d6oOX8MFw5vLA8/YtpqniYUzfziioxnsW6kLXQsDQB+Lo0piMbG
86DPuSBr053hUtMp86vNk79oC9RQ3Csh0/jwXDqufAzLCNWbZ8eRsneY43E3PTrY
w+nKDxGAfVEX1zQxy2QkVYSnk1YPcWRS5L3dWsp2QAPDok4ZXnSBErCT7wR8QrI7
TgbtpdDGkrWbCDrMkNV2xUccismJExzlbz+7TR5D9uiMy/Kwsm+Zf2PV+NECixMI
8dPVvfXBksz9quKToRyMh3QA+4NuyV7YX9TcLIjTLK/FFEy3cKIzOp7wMdIKZj+c
q3HhMVPfd0cwffDZJuS13ouXvqybxmWA5j3qo5KVwUKZdY/vE+UVYQ4y7QcpD/zF
K40GmaqjDOjeYb1Yt9mZcrLIDh9Keo4c9DcHYP4HDCK2QMCyA6AomNjFVXFOfHP/
GEkh+gDmpzclC17+RwnhXFVUg8xNBdntYdoFq4xsh4w+g+FSkw5gjWgsqLI1kNCC
GlXCH72MY3tIbhRcLBtTdRM5eu+uDu0dmWe6AUi5hAgSawZ/fTZxFwAi6JKS3KAZ
qqYky+yYi5daifZL+ScnPadDc3U6+ObBHNeDJJbOtDidrE9MZ8h73yUr38v/tInf
TSI1Hc/mGSsEosbFLYQM3Jq4ZSDkWrtl+/Tsw9Ha/Iv1fOxStkVY20yRuhEvjj1M
QdKaDBr9a6rSEMj0tJMzUevtNTHNp7OB6qB0NrgqKsMSO7FeF/Vziz+w5T3NHKzP
nUsyJxnQR3HSODvi9Yv6xqzGAP9PI7U8sBRVZZ/5ObcGNo9w9y/3SyIKLjqPlRzd
MxhlHrSVYdpJgNtktb5bx1XGnGnUwPsREFfeeEjUhhFODkS69f++eXCtSEisHDEw
xLSjZmSzn6//nBVb2NeOXHLehVivvCwaY9wrhAU9ST9DDbYeosBueX6EhEIF/XHd
vGVYbC3nKBqwBpqEA9B2YKvU3YJ4ulLDaYTydl9pmF9UT5lUXctHux9EDah3DciS
HlNkNE9aX4J2S0cV38U6SUTIatwb/f3wjd8NBJqBcDt7mNovO1NS5tANqU9b4KGN
cYarK1++rDzfoVdMCeAd4fXacre5zMH9hIqqqEoaixRSv9khzVIfi7Z52os1S8mR
q/IOkFKg7zV2ahVA4BIHDzEoK9OZ8/XgvIafqFmmszyccQlTm10CiUu9HOfDpYQS
+9WirfCTUrA2Jw3T9paD2jSzTziDYM11KpnAxL8WXkFdNrbXQeQIP8TdyG+X2l2t
pxAcaNsdL3lEEhW5TQMktHQX3QRkjHWCSsIKiQ5Mx6wPunAjA3QIxyLPgYNnDRUX
sYZdfCL2AQd08npXA7QCZacWnoJXWH6z1VcCIQKQLMGaGxMquV8sv4LCdm45Px4v
JNGhaqmEv2y1DhGKvahLwd3JAIVlRiuBVgmo8pXGvtYsDdHESJAt4JkaGT+Q51pi
c884T6qD4UwxzprCjRkmRoRvUieqsRVg343tyYGfPu/G6dczhiLce/V7UVITwFGP
kxhxYduY4AkiLHmjEMqANSG3PcJtIuExGJanUqWLyqiThtpEloXh9rm5JmltmRTg
o9aEqhRqMXnTqMeaNzPnyDRteBARM/Sgwfr+s6zfLjwzLjiy8gCiOpMOdeP/CBjy
DXp9AfUnav5WK1pVeEPn6nSw5iitMrR8F2Z6vSkHl8Cwwe6bhA8FGddNb1skehUM
9EUaNS8DG0TWbWV6q85qmGjhwj8uTy8bTc4WF9yZ8xRQ3yVTqRVfld17aNX8OXCS
3YGALa0EQXG6FEVptxodM7uOTbO5dg+uka5JqRhedkmJEL+St8ckGDFl4T92XSu+
KaSeleG+crrkyXTyUrzlwwxhV/TqxOPqUqJu9YudxkLNUoSo5+F75B7iv70IObGt
e0ADjS+AyDWkUeKfm1YesNWfWthePW0smEdSP9W8DsJql6Zu0zBSWis0LPoQy0dC
IXUQuXuTikF8RNAs5a7qUxJL+Es2/rVjAHZZYHVn6NglzRUuGopfMB5q5cwcP3kT
qM9LbCIwIFcoAJ/W2OdRunr5ZkjPA+k6hmnmvePIV48lzpBND5ldQ8nqqAQ7KinA
g69rE+zlCngcQBbwpgz7qOREeJDSIhJAyKKA1Msphbb0A+v5ud30chx534fOwY2P
xS5ppxz4tae1rAk2fg9PXNVudOJCf7rPlojpiMjdpPN5LDNoksmWDKIGb3ut4kGf
f4jC7hsqhSx75DDmvQLwY1h1hU78IpjahhQnh7p8eeGOnTyBbTGzxzSVDtVNTwmE
0wwc6zbijXBKfGS/sk7GkBYckpdsI6pJaCzmMlDrAIdedDw+GfgWCi9XTrwJ+bon
wZFUqgPUOT5rBB4hEFIU4NYVJzI9YvJQdPaLWh75wpeEgj/Accr5OfETDLMpfcY9
gPtnw4/WeTr7vhZHOs3S1JxLzjiMhQjtyzJuFTJ4jLLnayUXdOpJHyGf51co14+f
pDJxebVU2/219/XFyM4smOsCAemATg8puIlmpCYeAZpZth7Ss+F0mQGXichobxA/
/Kk4IblmH+J8PA3KFl1XhpJH/3i7pBhHcXUmlAQz79xggJc9PQJj2bR4NzaqfQN/
Nn2ZDbUavmDtomxYFZ28KRfLxUZPRL01sP2Un8I64t69JXYYXn2WEhk7B/HvnUMD
Llc6CwSBHqPcCeptgsK5EoUPoQ7hXOIH50lo555r/W49GKVjzongR+/d2oVUerAI
6vu86oUpyXUy50nAfUKqHCfiENgBR8wWqN6JF/hdUR8vrZWrqGLI8xpoTwQ7nPsW
fJsWZtaW/0g3gWpuYL/q5GKCD70SpycwsiA2BLwJLUbRMfDReooMaEcfMOdiM4NC
wTfmMXunIpCKPwoVOWiHIVkG2ZvOR2gcgeX+Va+HVRbR3DyYiXpOG5exRJMrJZDe
eXpzjJktaBxaMO3WIA6hPEEoUv0HY9PKumn0fl2QxeOwgt3m1Vq+pSEkHP1hN9Vp
lL/y0QbxjKMv7cdYMS/E8KuTnyCcJKOyxq5gqrOHvJfH/fb5bD7kt0cLIMx/5kGX
1A0M1g9lbFiLElq1P2+BSq77cqCaus31FcsFeGsdkE+1FVDQUr8IhX8x9aQfuo4t
sMabfcUn6Ib+6KvVO+Z0XllVYWYmNlPY6ULGsQjYTZXF1w3DExJyu4KytST0hGAD
RokU+wReTTIiuwsKxjV6EpJ+GY/4UvdtLrkmg/QkQZF4Ncr+MkvXVRLXKyFtVJNx
BW0CgJs6EFTuhlK45yoCZNxQIJHPpR4UKKzUCcXwfPwhDifhWDi0jVkQP55dj2Jl
6j/+IkcXpOsH5ZSrSt46cAZcj6IG4mfRmULYYtjSNrtWFsM2prPqMbQkkG8hk6fh
oytlUJAKwB0ySfN0mK+eC2RqB89x7VVkNvRqhoKWyCzk+YMxByIuo39aXxLb3Zb1
HHzJltJIe5yUqQz7ydNxbG+5qh9j/lb+SBrjZmjA9QV8IC3Vo7vMOydf4gTv25V0
O+mpgHkHDPAA4wlBog3BBhmQoXOs5Jpi3BIKoNqaGJd1Vxx1ZJJEFSWJn62GAS40
bPBrshFzkTiLcnWVLcHU+Bu+rerJJ7LRRJr8f53+3bXV1RiqMW3pYzmkQa8a1f5K
LramHogR4kqiaTBVfo8BS63UdR2RobKTWp/u87tscnztoq/C7i1BqnpCB3b4ULDy
6aHGOpHs79/4W4SoQ6UyG4nviiWG688SJpAftvWryv6yRBqyoHhjt3DRlYqRP5Hs
kHyZLAWK256lxYzIXTX4eDuKVceLQFN1R4+j3Lsz0RXWxb4eGcfbEMdym017QZKv
m2YH03ExzeMt/L/lrw0V6DqtB7UgUhJNRNDFuDGw2k0amZYY0Ur16yDe43AWPeAA
gH6/Tq5Rxg8hx8fpUpcGaCmBtzCyVcarynC4YsjHzNtfFcD8Wi7s7OqvC88yAurI
JHK1q89H0c5rUeHfbPUlLrKxO2BwSbWjca4aBKLkbzN+alxCyuOWz5q5SFFtNIuo
conVIL/IBPOp3igBvruWNe+wyFal9UzrKbZZrsKHLK/U4zy4Y4KqUVQ6zncn2HZ4
NhIbJovCxnzUyHOrwf6SLBi+WRtXe7bLWMgPvY8eOmvd62jkKgtkLHEpmGHDuG3M
md6j1xthJsJcyz72Wbo7GuTbJyLvehkt9RGF9R/WxT2OEDh5PYXVh2h3oOyYft6b
cqDhHH5j7SgAuyabjX9qSSyQy1BPqFoQ5xnTKF2iNdawDij8tkftT0Nd46m8/sZ2
uD3HD4mCAvAWrKSdjzG1R2zftRMfS+psbUtsUKF9psuLey+49DrtntchxVt26/af
A3/5Jr6Cq+SxUQw18VaBrSR/0xVcC9d4GT+PCk4N5C3QBo6LyreIad3OqdovZUhR
cY1+C68mC3llx7eJvGCiiZHR8Z7vHIRyPjYVXyphD9Qx2yeXZfi3ELmbN7qwZJ+h
TlBFZ3rZujw2DmJ+C8bs6WneP/BixHhXWVbGm8URfj5uWBiPYoU/ryX5AOEmALBb
zifncsbbAfUlbCAdPPkwCCHSq482wxolP2utB8hcLpN2Lvg4qx+FzZKTXs6sds1X
R4R+8gR/ZWxgNa0ffeCbLweYEiNyzzLgpAqZzDajQ5/Wr1SF1QzOCDtpq/Zx9Y0d
Oii7XuD/eL49EgL6HmCH+htyf+fDLYV9O5PUidtAYD2ig8hlE3EGzjk438MXs1y/
7TxSnM+FyKvG9o49YcfCD9/wDpMWgaQvzPulvBDfHVa3kajB1vD2Jepb5+MCI13h
ESgpCw6nO/IryWz2AEyTnLqk4GdPooHcQXJC12vU4cllaKWMcTTeTodIavEDNnoV
7oICV+K4/dH1pEE2s7Ad9G5D1k2fNfc3PgavO+nvTq9gjAknXUEyxBKN2crItm1W
vqmGEBWK1zsYS3USth9VsojwbphzRIlXNIMxDC1MpxawnXnL8QoM6nQoq4zEiXaQ
Gqyp4BWmh3j3X5E2xulYMLX4huGDsFlxpSRhA8pstcVyarEVq3cwVFF/leox4k4j
e4mrvEDchfdnIHmERpD+tEDCEi/eNV0UmYDpRuV4wKA7mKWRgASI13I94QqZlISm
g9WrlaokWavOs1MS1mKwzZfaO4JHtomUzZl0JblLK3NvezAK5x+lh0UKtRa/Pogf
xyzJbcxR1CQK4PRwmVjJ9J1ewmQQKma6zY3Y8YaByEs9Gnw+0vVMn6+JTfMaAllQ
bMKuCW8ifR0ULTK80S8aXZsXdgOusK+5FsdkOTyb2KC+W57nems2fglDTA+geGAw
zRd/sy2632jAoUCLv2hbgClfiJI1lB3fik7374KsREXbpuAziEE2qx1m4z+uiM9g
4vRdY1A6SzpjQ5jyGqh/Sbff3rJKQZt2uSoVIlARx4yvxKzELg0okzgcB7HWVbgM
g2BLsBhcYNwGXX3pPYz4DhHQLKCSuP/5ClFhmtSMThKVsA3do+meDvSp/AQhXdPL
1gOg4NYzBU62EC+/Z+9CesW3T6Chz2Del1fD+wZcWPjO/WkRW68D0/abtqIJFnM4
F64Ekf7YuFHKxTQbnCkcdP54ySb1In4HDFfMll/Lo/rWZCT2EjRHL2oUEicM3j2I
4H8alESfBWToUvNHsXOE4ctUBVHWkGcZvct7TC+s7PG1Ff8dRIcweClHeF+tTWhM
WDUEmIRrtSs/Vx4ryLYxzPLvLH0cJBGb7N2fGMmBoF9bsftbbZfi27t4GwAJa6Eu
3hkF7QplZSqNNctd6z8Du9bjbdBj5odBzIL3GEps5Rgzvvrvs6hqBQX4+D4a2ahZ
mNjjkutPQZPoWFU75KYqpcggstkoTquikNW0YAT61cgcjzKvV3o4asA/AVWjWarf
qAkMJgNNUhQsT1ggtW1D3oRdavS4EzyDRMcx92FtN3iqVceuAGZaaz3tNUmilytO
Gpxxf89rq3PAa2gN1CWKkb/oLCCOg4YozUq6cd4sEaUJYoFLSXcskt7lMlnz/TqR
ztK4pI72hmEoXqGMZUKUOiJdCIaPaEDoPJJeiVqEBtGfDQRWKRtOvyEYSpL8375f
yYaFnbKF6LTgLpFkotbWXzmPZCIvVzYNtPXX1kSlsEDAGPc4EsbDKNC/ErcsXJ3/
SBPwQrmOmzP+9mR5jiv0Gy2yVtsCb5BPJZmmN8uDM6JvcS91eHZa9drGIHwqe5SX
485z8aLUv765/adnDZU+WWeDPdJxLSHyHz7whdfe3L0EOSNWWOc3niaDBB8xIMsU
qbWzPuOo4xly/W71fHBSwchKoV1NwgSLxLUvx7Ldz4+lyp3ZcMv6scDdYvcYv0E7
2snad5h1d4zfZxqmabH3YcArmiiAWcG0NS05ZEDQ96os6g82TQhvZwvjmqrR5wae
MN1kQGXrQimFR9cfvO3X8JcOWab8+HiwTf3TQ7JXxJLIZjWwLcQMBhVia4ybJ9Ew
7+dZtgMW/2KVvZv1BQNEQrcbo6kZbmDBinGmfyTZpqYEDfQIkbc2pLaPlC/tImV5
XOJ/WV5Qe++mQA5bund4mw901Ee0+pjhcIxOt4hwQo57D4Wm1azjcBPcm9niFQAB
9coGm5Vbeo+GwhnYA5WcU4hxgUieoW+rbpI7BTrGFUoB3oEv00/b478BASUfD6ts
Rsf3v63VB+LjidaN2oaFVhxzeYcSMuKDhrLZURJCmuVZ8ZcLrY9s7Ty9op0r0l51
wFNW23oaW4j7ZLp1LEKrbUBqOyj1ZHkPXnBmtSI3/92sJSs78R7OLCE00sU3W2i9
hR0k487ME7WVJyMy0QBghTtHAfLdzV8p5jPMCzyu/KD/834VevUertKWpq3oz/CD
wZF6n5kTIXlbzCnpkUibISzadmEhkDjC15GEq+n4JForg0hCLXlji6jnw5cmXhd/
MPdh344tlDo4/CscAhxwR0eKwyM+iFT3iYQtT1bLa/ZW4fo6gUrgDO4rTz1HD4GI
4ePsh4FG8Lpakg7O2oCw46Jqzqc1vaJ4XYOaIu6SCj2gS/cOh7+1fLL2hJxLXBKk
0LZnaWoa4+ehO2A9GDK7nMiYsc5IvemB1qPvOUQHrWCljjZCxWpv08WNBusbdzDM
oSYqbs0MssatjhJeCaXK2/nVbhZm/rNpWNVIx3b0XzfTHVYToevzQVEZ7isrqJol
Jb742Zb2C+If+X5fM4CwFgRWrw1IGCC41hnL7cZRGp/43abo8QY2c3QYrf7hxeL8
u0E5Oz+s+pKoqnvlpR7rphN5gKAG9J0QA/UDi+30sGEka7cIwx4ScWkyO2XNT1Fu
g7GDe7Drw7qjkIPdZRnfFIqDAv4AUuFOFaSBKbob70baCxV7Z/XxhlBmwkNMiEJM
SGFLugacqO0ooasik8LBaBln1O3HZ4y91PcSmk7cpMq+03iGnbv2tmmU0qI9CrtU
qDfnlOUM7X9hYLC8egvpKuRecCCprr5fkUDyx44xyKdD/tMRIOUAJIU4bAEqq2hr
lBoZHUcuYWVPK1ta9WE9SfhOAIgFdEKVey1c+cc5syRBbtBghkZLf23uWuhfb9PU
WYPt7XGmr/V0mqAhx981K1jTulVM4nFLiuy5N8iv6lo3u3aaou282aQkf2xebTV5
Fe9DBPNMd5ApvrnTGThIJid2h6S014mOivDkqbtw5sljmdofB1XMNMUsfuFNe4TN
lQfUotVP6C8JzYv2blwjW3lnB3188m1RUGcyfBnCPtJ2DIH9p6vBSa6hgEy6xkG2
yn9755fjnqogGxqsxtOR/ombQyHdJw4W3RdUslvC2Z5U6g9zWRV8epvbTTDNsu2s
JAcngrdQG9bi3aohFzdNF/Eld+X+lSvd2REGY45pAyN0yyoEWolg/krhBpuSpbK+
kh9YiIrx+qJv1uk/mUv88LUzfs+tix8Lu9gZioV77DZ4uR9S2oiMMOmxFbfdgROD
XEQf9xIEYfijSE6v39EkCKi5MpIrQEgPWXw0vJPTTiYVwxW9k97ISeBVDLFpgmN0
7H/59ELHDxS6W4A9uzV+lf6Q6HieiSTwBBs94RBJCwi7oyaJOH7VkjlcyM5RQ91O
SZxBADLHsZJ89v04jQgk55IVBLrSi7uHikGv+sam2XB+7RHC7mzg4u5pSemavQ9+
NeE2fGiZMImD42ZfcQ1jM77WkPm9WRGwNo87KPub0FB++sTP3Btt6eyrQiLp7vo5
inwXX+JjEkdUUaNHlzovNB8R2oqwbVGrZqMTUoZAk6N3IaWkmnpgcEOWxJcq9+2G
heG9+ZbY+cPZpXMfUnhHWISKGf6szWgyUukSHNRckNKOo2WDgzt55HntEnvmOZJi
xhitfgfLH0dF9O7BAeW6uAsZ3uvQTzS8VX0SUjoUtRoOSf9gptOGW7vEryqtMSPo
gdVvVKP+JsAMJ6Nf2znM9IYO13ztD6XN8rJHk8otpZ+iyrbReFJUn9Lwdyqf2oAT
YsmhAWqQP73/Geu0gc1ArGqHCpShuTCXgPk8g9p3ZU3JvWUjbnDo0D98cW2+Snwc
/1BGBEbLIeiBSVJy9xaTOdcX/3dd5GGLnSLOheQ+w6FEKhFOvfvtIwuL+QcuHTCT
38tciB4DnKwrwdFQW+vZj5hshauJNjS+gHY4HKjopIICfbohSJyH3xPvTS0oauEu
cyHUoWZSEFm80UNmFSLKOK7sKwwTP5SHZ0qibwVIf/vCtsciTwcqp5JuVS9uYgYW
noDKnxeu+LSb9zM63XnKKLefXlJQUXMdPLCIJo+jHCWRz+Fqd/SHDjP4qenqkC+n
YDAqhEi5Uiptpyi0w0IQfiBGuvqwncKUTjjc2HhSlEH+tkY9Ey/0ZckcLsKo9Rtg
YqPDpEOMv0zeYgoKWSeS+p7AavNMZMbcAPR1EI+glspZY3MU5XGnblylAG6ekMv6
0iSlZ5ybsjun/t3RXMVhAOUdv2z5YzoLJBsHyDl5mzW5UKuOGgGHH+HS1mELc//z
3dIvXjZ7DhiTYVo1Q8MIijFMjfMkRRD9A8VZDplX03uEB7hVBbD0UMo9t5yC49Ch
ZhFSM5sXIVl9kvjsDlOwNj/GfLvO2gq36bGMyZJMHbI2x0AD9+IoVsJkW5t3YFoi
H+KgGwNqKr49T721H5TlSnX+dtxvlvFbtRW5By/gVhft9dpftuK46WyyuLGA+QbZ
nF3JtYRRBjcRtVlH23cHr5V3wVUwDVJgxp92mUHVkREYftf6apHVHjSkmlJ3muxJ
BTxXO4cu8pPkCci1IFBK/7h/Qac3SCGydJ/gM6JNlmtuYXC2Ppf289JVLy+J7MWz
PnJPXXd9r1Y0t1+uLgtujyZAQcFBdJjEirSLlZYrkKofMMC6R86Aw1PoUXFzBkVw
DQQwHoy/x1ZSWLlfcsk3UAo8sQYy+2AB3YtaMUzlyHFj9HFlJdbiUTYVGqQ3shH7
v2tcu1UQH8jurfSN5kjiuTJLpU4G0fnUmlYOFJOEaWdlyVFq8Qxq19akj2cbQXR1
jijojovaxEZn82N/85q+TBfcnrjD14nKK5s6Vnx7F5ouwZeQkZvAJhDT/GRG7PL2
51I4/GxHb8YjcgQ6FVBFeXvsu6rU7WTAVE1MNDRZrm974OpqUebmULBotUw3IulK
HoTrFOiXf/B+5OiPRdzsUFkerorNKWkV+4XBnGuBA4JB9ZYHi5J/b4AyVjevq0xr
L8X6gd+krhiFUTokS0mNTqb6O9wYJOJRzCuER6NOK583/hysjs2/3br4toFnRzdI
WM+UYGMMxK2W70D7iU6uZKJVuDLv6hPsZFjWWCau2+DB9kz275vmeIZhfla4EkJj
Cs9pWDOZY89rPFYq3CsJHgqOjYt+gb/66/vmlVuR/G7dk5FbpKe4dDSV7WGbMx7Q
iGR1ROZb8OF1pqkPysymoDZp+CK9QCf1wjrXgKEw2GFi09SXj5BDDG+QpeQ93pHr
b4lMXlXuvD4UXxdZdo5Qk6XUetua94nprOLotllmie5ScxX44WWtAeaQgcq4BZme
5Z2NyFjy8I4aTijIr2oNAsguEtd4VkOtVaVLYv/fDZtDD40CxX/zXdtFzhH3vgyI
uRcUTUhJDM3t4LW0U/psb3meVBWxemTiS+m7nY105XBGIiKBzLRj2DlZTVDaSZR+
3azV+o6rNC3sUC2DoORVcKwFhq4LoIlXlkXSok248j7cpFKnQuh5tZcMdIMk941z
4N9ar1g7sTNIsPlYuY3BO1SbbbQMxz47CnDNhYqYC1AnANU0OgC6tOjv1j2l1Q5W
f/us2wF4V+O8YTy42N+aiklaV50knXIK4sD0E8fCCwMZ+Pwwmxwuj8IHDUnzsJ/o
5irogDdwxZF/Kb9mF9Oinl57AbSwOSjnJSPOTp/Tm+ab7U4rieccENxks4QOlZip
alxwdvwkVODpjTkq9WXoNk9P9PEcYt1P6PHlC2LSOxw2R8BKwMnw3g1kDW/sbASQ
n8mzgqR0kAWMMYcg8GpMUnxxUfZ/p11OQFQmKFUzQMzRYhic+h3koTnjan8D7qOK
RC41N0jCQmFrwy4Uuxqf7PFXs0h7nzC4oLm3KJOPUAes/6bd2hNYTv2EpN2YZp9o
4RtwuwXNm6K02wFN3yDTk+nWWhrAUyrzzfJC4T3MRsIxIZBs593obTU5MVATALP/
JyIkMhVPbWpK9gKthHBCHoGIK1rT44GkbOqqr+t0iVRE/EC5hbMPh6zGeThesP5J
zAT4jWYIZlWXMnDtY/p/SdihN1LdoSBFDftIJHU/smNUamz42plXSVpO0TRcYf4Z
9dmdah8fUHtJDxHMbTvsPgAUiYsHxgefYMv9Q5a9nj/KfSxrFuPdpSrLjErDxgyj
iAdQRVL+su0Vi2xkVh5+H+4nuBtHXRr5Cxq52orfaqI71CwOUxTUDcs5/3vqVSKz
vRimlNmquawtUWxVx8VY+dOvjlU//QhVzO9xaEhoB+lIlhTHoWtJkyFQ44ThGn6x
2wSQlyZatY6fKo202ICAMyPSqshpePF9xeL1Sky1ldbyPZ9h9qtBsKpS24SXVEAm
EGiysd/A+tAK/yL05ngzryvVCH9elFrjNTE3W89oG6NSgD4NNMCsDwEbetClyRhF
Yjl2Yyc2tH8557VuBj6fhC69Io1aCJkhcEfjfJoDKmU8rST+bNs1SADjXXfhrmJH
RO8N6OXCkxaaVh4VX50Wsqr+y+IguUd+luvsjd05OX9mGt4SSBvObHXo1K+VOaov
U06WayWxQYkzz+YFJfNL3UdZCVaa3kvEKq5TeZacmAN0IrxnPT1JfKY5qMOLu/YV
Mo25uMopRP0FqE3UUMQ7MQta42WhwkyqYaM0J9R3ug0evOt4lyKpwqMjcr56fRRG
ixDxzninlad0nxNA3TjdSF4M2EHaX9gnX1CqsCAo/kOV7j75+qlLYFIpagf94sz9
g3X2pJAPbnKiu6IMlN60F1uR+TgFmNVEGvQXzfleJLhEB9VhXJ0OJB+ilVAM+JUW
WlINwSF3NSyPGfse4xHP1TI4yDNUklY68ezboK8SSDC52xC76J+Gn93EawqQfEe1
gGhIRsh7uZ7y7h8fxeofEK8Lns7yH+v/1ps5WYm/utBPTHb/CW0PkzHDY4pl0fm9
bH9f6Qoqkhidtnpl1wR1+Wttg2tWwJqsQFibNiH4YoEvaSa86bsbmRiSgBFEsR6t
ODoCTjsPqYe3yWSKC3sNq2UFtazmcIGoKVmuuUiQm9t3dZTaLdfsB30pMf/ZOf7y
uAv9vlAek8VIaWb/Km4NUHYhZSa9rm9RS8C6SCTHhf3rCYTOmDEWEO6SurGtszbd
eMKglJQHfzcLpvP0Lcj+RWh2juZycSsEhYrWnhgqPHb1SGUeoddoLG7t0a/PQXuH
fzFuS4B4UcL6pmtV/Vun2cGP+n9o9po1wQC5t6WfPtvvILZMQlmTGVEzbFm6lhWz
30m7r6Bz3GRfe/+5/zMEfVDO6T4F/blm9Elsj+WW5H2Z0ya6LjgM9pXKJ+Et/5aP
yv9jZeuTU7TlSxAq/DA5j/a9pC98IjwF0aEopnd5vFF/clbNZnuBL9TLhVzn7xRH
kCSb+T4dWlPx9eC7+2oOjkiRkg+5VKK6vnYenrh71xq+aUY5e1ACZhtoa4ID4GdM
+T2jT0iU5MJ9fIrRwj0Ep/dLhlHcAufhHHtwmEOCxK1kIjlQYMbt+qHYXYghlO3R
4bqikFzTMiNUhG2F6PC6d3iBvUeyM5QLoAmTLrJUZ+yydW+UhBpvqJ9JIt1RgHys
jalHq3upwKNM+yXhMK4U8GykZlLQMd8avrZaxV/SzaYPfs0wYUUr0MpScpwODOFa
j9Vu+PMbq2UGwEy+byIn7Ml8bL0j/sZeZUPXCDBzNPYrQPY2yiVsBSO2xRdoPjyy
pWB/Bc16rpABg0UXY1LKDF4nk4/V1pt6TIZJN7/H/4DKCdLYNhtt1e9caCFimBXw
o33uNgH7T2+BcL4cztHu7dxL9uRewnITCNkaOIh/KpOJAe4hl8rbwWy/NtVfvCR6
yA3fYRQIz1HLxySBfnWXNuhZw5jnD+yWLXQ7/blPWW1NhTdPlUHGEbQcvpMXN5IZ
J78Eavoi9+tLZfcb+0zS3YhR4HzIswbd3P5qW0JBc52r0qRuTCfSOxfNWQb04VlY
fac/mDFcJACHFETfn/JPJgHkqDiYBc+dvgOevTkwN2m+pqU/MWeIzFcBg3fgikyW
7mZAvEDASE+eCQCrk2ChjgDWNQso3ZAWqbmt8Fd5Foqo2jmIoEU7M5Pg2EyiARqM
K/hVPktA/g5ac5fPv+SND8VyzN6DYEI8N/0kE0wtNrdzrbSzVoP/E/47JF0u4qiv
7HFYH4/4qsrFIuuDo+/lSTBMjH1gcUpLaWLgSMTyal3zgOEQXGK22Qo2MHW2IaLH
fPLf8SQugS5BIulCSQ6yGCupzxFWH+caCBQkfrDXuC6GS/FcJcWwbKECmhv5ULml
ggCszIqvhUMJcNNFMZ+TWquA/x8zlYfGREviNh12Kw4uYT2tS1WKPLnNV4NEc2aI
9XNKm+8JKvx6L2H6hWbje27a2wBXotc8wk4gJYSAbwhzEGxnG1pcmG8YtxnecjnD
MePlzWeHbqYKgtIqDd2mhOvY58xEx6OagZTjjpJ0csMDKcBI5hZlm0MGbT06Okgo
RW/wzLpMS38KhE5gQCsHQCvdYCXgmbLO/r1mKaOVBGCT9nkIqNpA7qJq2l6EqwZD
cAKCmVRO0o9TEyO//quR1PJ16ffiPskikFTPpT/mBBchCmbyjyfuksD10rvjJyvT
qvfPeikasiNAHO+ru3Ln3UjsBJNm6JXqbT/Vq0wq/4bcO7XDTE4Eu2QnUddxBB6/
FRYyGCp+npQ0IOx979amxNek/115yvhkTjHLNOhls6WkdCX0dCuQT8OHQWPj+KeP
bYNY+dP79MFFotP3OjzIeD1fVyC8B2QBH7HkO5IbOIXfi0gfxrbV0N4z/+qOWVY3
Jr9UTYv5NdNLd691iYlhMRfL+a8vaf2WUAl59t7AfRrsMNLhDoiO9sGTz8n0TfMZ
MXVoEF1Qkpdq6L3Xu3y+LFVrGw13rOFOW2Eh+6v/YNENYfN59/ZiPnC7zYy5CjvW
pqHJKAI/SUFNoLV8NUY/+zcwaYsOvelyUfyRJNr12LUEineJOmmJhcdFDqnsJIg4
w6MHuM/+7KJ+WsEKK/mz7nwv5z4II5hH2fQ0A5tiyy+4PvPP/6pxMOrrX8Bk8ZbW
56+VIKh3aUjxXkR/TJu9I9rcFBDpAK3KRDIQ3ErSysuScg9i1f8dNL9DyzmL+nJS
hilGW2N0eIedCzxAB4I2oF4OE1avTjbtsuDB/yr3cQ1o39E4HKtSqtGTErCKXS9E
wqKyDokfYdKl9oxaxNYxlyAaiSYBqf+vvec/vF/8zDUu5WADLYbX4tPSKG+lqpBY
cJCCbCgYYqcrs47CeR02XF98WUX548l0ij9wU5kHDqYJ6wfvR4y2bsfItbWr8vDp
hIxy8Bd1evLw3uPKxk7ORt+p6Bi9geP3xvDv3uvyX7n9Ge88JszWBoQ5+bxJ87IV
C2vnVu6NCkWMtAFX9HM03Ux7gcuBeFA/3zi2P7BUGydVkfkh+2Q3c/bn+xlHsYgD
HMUTb7sg6jR8eVmg46KCtTqPW/5oYf/N7FWPTGrPRAYmcp6NeqTm/jY+hw/3VFUy
hOgSkSluWzKh9R38RD2tc2c7gjDW3DcLbx0rNEDzR4V6NGl+EVeZFjorCOfgQMsE
Q5Ps4sG6dBK7c7LZM3bhlbx5z7ToiXFgHS+2qiHfD2GtWDiFTzdtHqriYXsCemhj
hp1UWcjXbCkw+KVOqBYbYdr1NDknkBAYosvcBHg+M89XcVBo2ROpZOC5DJIqIP/b
RW2Fs+DfMezNqqTunqFQRVaEJLl0j9l45RrReLI5mnsb5lbr00rEwn+qCF3nHasA
1s0jP/dwqCNXilifpGqjWkNZpYZyUA0fuk63jQieTP6RVcqLrUU9pfgb+ha3DZCu
ViCr89oa0uUZPLt8j8BhfW6YuIi5CBHJra0AkuaKQ4J+fk3tzCGGnwE2kvFqbNaB
GigTMnFOj0yLpRhsxtNP90sLG1GMyamxEMxyzyED11z9wZyepfD+cXOJ5yg1MFqd
ulENQnkvGXiKmfihinaZBlvBKnwlYpLf3ikYUgH1//5jmBF1oDSfB3ddvhL2byxt
lva9TjE675gDQKPAW2PBPJSXlRUOCBqLdFtx/NWEXcABK/kcOo/2fIlqJsp2xEe2
PfObxxQkcASpSiOoLJTSLr1o6wax+2aS1UI/hjwLSvGwznCQy67RYxkxnDhzOwxg
f43Z+p0KDPmL5HEfWb3+Q0if3ENXWOaDoecFQCTCCIYJdT57FfNe3j9TSlWJ5R4E
qGv2XT5hPU9nGoKOnl7JORXkxGcHB/dlOjdNTqJrUQPYR8zEoHQCjPYTsnD7zzqF
rvJMTmvnAljAuGJ2n4uQKBWxxMURQ7xmb6eQ42picrvVz3tkwyBW1rdR1nVrfF0C
hNFZH53EVEIV3+V05cSmu2FWL0AkThcVJa+U5/yvIHJkuj641BtWQmqhOIOcZpAn
WhWZ76guLz9ch2SwP/OPNuBGL72QAvR3EYo2wZx4DD5BJHffANl5UsKSA7l4Iei+
Ub8dtT3lLgs0/X6lHFF3VAOAyYiwDjDz8p47RPV0dZnQIJz9R23SySYF3earhbGN
I/rOKEuMJumUXDdGja/I8q+6n8ADxZeF6LSpPsYMce0lcys5BHryl7sTDRvY42/v
tURYAkLLMh1lEvxK7g99MeaM91DgDoVpKpdLFRpsi62MQs9dIftuLoC7s1MdEjsL
kM0yNVp0HF+LrGXlP1mex+EBwU7Efj1lJBD+ypon7tFSGIdCT8kG1Ufg0ih3DiZ4
6ZsTzulJIRNYMWZVx4lqeU2SpEii3YrZtPCBs5l5oebsMMUlTsTqc0Ke/pNSX00k
+6LONo2g5mTyDaBpER3mfbdeK3+vqXGG3a9k3AZGWqfJtZu0rh+kqsdmSIOz+CSG
dpwRf4t5nYdwP3u6ZnxbWLGiCNFBRzDBFPI2RSxkBUoe9Vtpmlz7EbhTsaVUnxrf
KE2zqRFJPcixSR2cX9I6MU2Gtdxyx+nJt/6sVgHtebul7vBscXmNLTnrE2uE89o1
IB5VBPT7VztC7SpC3Mu+Mg==
`protect END_PROTECTED
