`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KuLlpkBSS1MQwPA9gbz2NRrSSm3zEVWHSwfPPTvTSozZCfmotw9Y5nIlAOAWmWjt
NeEzHljkkCwXauZ6SbUrH2LUIXgYts6QLX7K1npr9aWLWkiQ3cNvcaWsz52etyqv
Y70vqe+NxEcWl1TTl78vyPEiWJDDjSwW/rPw9gB29f6Jq5DJWiI+WUvTGfKYf520
hIwmyo4wKCNcaW0z/3cYQKkvoohYShRJMWU2dE+XCh3Fthgl7zslsDNbhhWlUZZh
bfySx2+/iRBcdTgLEbahhcBENPAwNXJ/rbu+5xLsMGLeayjPoQwuST5l3ebAupqU
6QJoC45bm+WRQPr8SpvvQnu2/PojvSFZOR6ZruA3radX4FpzWuLmbcsn8zE5kS1v
T+R2vH2huHvssepz7w+DUzAQxa37zFFCi3lTNxwmCkhYTPrCjfk0sNw/Eg/aty4s
`protect END_PROTECTED
