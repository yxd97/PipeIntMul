`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VCTrDHPRJfnu2Adkqj46s97/HuS96RVqamB22y8DprbZk2uhYLF7ZD7K5xC3lE8a
mGN/KvEbnG3H4fzSIIhxYGWvCvDEIOkYNNg3bHNRU7lAjlomUBs4mQf23y9hEYpq
gxpRe1TbGgAbez7BlLNd/Vnm0DJdd0TVM1mOZ7n0U7+obX07x4dWDU4Sv82o+8Da
FUrpQYm3wSyf0HVz510Wdrot3zDehTNdI91fltwLhy2tgqNPR/NGKp2zWwBkbyQU
tbMu/HXg8VqmOtwegfDO9uynSYqdLlkyYN2iF17TYgok9KQ34WnW7m85XuoxFLUa
mzsxfEr4ifDdDt4Cgd/r0BY+BHG8gcZ/4b821wYd4podz0YCSLvkMX9SpU0f9q8C
TfAZHMjCFgIZAmixKJ4CfjUYu0L3L+uUOu2QMSXk19xbfMJIt2nogZi+sJwLStR1
nTCm/pDjc8bLfwfHZtpjJoWWzy84K4M1lCNFIpMReQsBUeoX2QoYaUvHuIJm/dxp
URgVqEvz4kjrbgMS7C48B8VVhT7TAs1cyBjo4wQou9gIisRaAgPa0NdyM/4OkAyG
`protect END_PROTECTED
