`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZpCAJHNbE+k2prHEr/F60vhtv25L6DVc6chGxjYPYYZuZ8LRpLrZU21PSZWqicz6
dsSct8V+LJVvkzaiH3/oxD5MjBGtB4c4Mq2cRoFOHzowqCBlCBNkIbe5O8dfA9xX
XY+sS5DFkJ2L86IcgKx9oXYG8L2hfyP2qga2Y7T9+r0zQpGpXOL6nrYUtm36we15
lk6IS61qLTDSuEO3cStIJZq0hTaFrMgzi4dFEw6H549Aq33azHqv1wE0u6YR0i/e
MCY9uk4mwoFEx+mU/pt+j+kRtP0hBORej2p5uz7bCIQxA9rxyi0OenJKlKe2ALm6
2ZqHaaGn1TV1AbYeyuRIQ5SYjyNLY2w2gSCfvU0GrndPCriPJBa9xTBZjC25UOX7
YE8KYcMEnZHA0MDcbcqb3iMx2wnjrm9MMxBjv9zxR1XauoQk1ZRwBeNz92954yqK
hWvS8IjAlpNDCu9/TUkzYX8W8grHO+ciS1CU8MbgqRrpDYHHiRU4DK3MjDdVYWqi
6XURfQKKROHEnB+8ju+iVwM6U3VWR1tAYWXpYeNnrtNoXYzdSEPUb9W3pk2uH5Js
ngg8xSMl7vJy/pvvl1IIzuUaU9mRNqj+V7jo+mvCbWteteZHSOaLm41z4KG8kO8+
nkKb6plLbgkngA6wPTyOk1bKIsw+E6RHvG2dh1FF1PwnY/U11mKeoQvkcWdVM8L6
Pu7kZTz8QE9uNtZ+Xh3tux+159Hbzp6tDIQ0lEu7edKiteY6+lpClXKiOyV8bDiG
ipEkjv/n74QDSMx4cjlnyRrP4/lSFcQBmz94s33qkhNOWZHo42a86ufRbyaEDNsK
7vC+PoGJ0c7Q1u0GnVuY8uxWqAvE0Cyabk/gbrmW6+Nuu+GGe8dwjJGmHbl/lHVl
423uW+CwPrniw2GrVErS8KdjZ14xT2tcksgjk57huF4I7SM4tSlPa3oa84qmYQsX
mqQPSks+MvFnlvjlcPa5XazjP4woPafxf/GNTG+nphczyJ1cp/M3Iz7Km6/0v0vL
M1qQLCAnN6VhEeBLfrv0Id3i0e8wXvBhTet2YrucGv6xtWJO+OgsE1eomnn39ksa
PIadgbzPvtz9/YRIrQtVnKRrxr8dl8LdlBb8hkXnjIxLeLu2JFG1K0qERagdxyu3
boWgrMezBFF2eqaEPiZaPPiCe77w/+h4fU5sB+GGf+xJGGGN+Y8aA4j2H9ivU1OI
Kg6ptDQObLKJIaUhYnGOwaaa0eUDifLQZoT4urS99CfRNxFJ+B6o7CdHUjVVr5n2
C+1cxh3utBJJJiGVjvzN/eGiKMGF3uxzuwZTY3ykGbJhAFBH17pET+O65EEiEAaG
fh9A7MSnlSTDJ0nn2KYKGK9xZN5TbAEGjUz8nzogbimBL+qrE79kLHavxp3wcAzL
z829EfyYfAUXbXlEk9rGwBnM8tFkDdlzazoGnp9UzgTkKPhfK6na1SVFLhpeSqXf
PR23IgLf/UJoKHAsm6zdvOH9OFggwSxyvJTLi3xj1y7EkJhUR3JQgiV4yUpEwNws
D8tbuhbuY4FZhRVLKW5doq/OFxKhZ0W3NzhWe8INQ1pu2oZkOix5ZlOnzL64+rK0
RXzAlt2SevSRceIzeltr33Jom4p5cD2I77HqEQt3uPf+EYhTmiZJlZ01Mwdemutd
RM3lqWVNuJDckb0GHkKzv189laEMABDsWN0E/f3+SYwPpKXMznsxY8eVP2sWWN0v
vs7cMNuOQlMEdXKGmbiB6cHABLBqtEcFjELP9YckIs5UXPu+JMjftGcOFrio7K3/
9q1w6I1rog7DpSB+HyCjA37I1VyHbGequZ5oniBlIGnVBWA2JXo/u7XeFWya5VzF
y6cVbIxpg3GFTkI1Wja1Z7YZ02Bb0u9xIBKDgx9baHNeiK3oNivjPWwRYenl3hUQ
ELXeAP+Pjzh9pt4Mwm1VZ33FPghL/vg44azH0H2deUk3BiA5dIpY7GwCgSFwCCvn
2sRy+GMRjsXzkVxsuQFW4lt9e3NlfZFnhazm6U/y10DKDLVLjMuLqIw+wjwAUMDC
HJQhvyRpUwnsE/PLjsE9g+yv/iuHml7d4aBys0Mvf37lsk8WNX4GcZRNc7vY24kH
oEQT/52FUimi8q8yEVVSZNSsZVM9noQHV+xnAEZ1emXTZIXdg8KhLkbkZQe7vR5R
A+4VU0NBLjr88IvG3u3321csRurhFfpdK6Ox+wQXdVLhJyyL757nlc61wfwlcnLr
pxzJcojw2cgOcyjppvi00rO3G85JGbmjOlk3yhrlbNLdpRr0Fd2rRZk6HR/5/gmr
B4/NNde/MEdXRqcm9ks10It/FBI0nFQcjWJcoCWLs/gE8gzoheYwe12brGMzl/Ko
`protect END_PROTECTED
