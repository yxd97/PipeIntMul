`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Vxnl7IU3O1QuAjaTIVmZ1auZGkRQrpss5ANGG6mCbV/56sTunSu+Ntfev6OEbsL
M6bmW3qiiNyZUm5R4JDSTRPdVI6Wl7DB9c8+Pu+CYDUITnEvhPDEjs+N/dgRrQAn
RSlIbavx8ZfFoXr9E7VvYnViaurPV1rhnXB/ugdv9fJTKTkapQmKlJmIeAS4GxEu
ZJ6jLyUiHJgJBA0zWdE8PVAKeGMnOl+DfKiMF3hxHDiBZpCLwkzvs0I2dyD7U4Uh
ScYx+s8eZ4gsLxTnOWAEdzH+mP0j5xJ5hzjIEWtFdck2p3FIvCJ5HmGXVsuHk0Qx
8I12XoDlVsJv/Q3Baa+Cej/+SXRP0sXXSW2Dk/v313IR1IehVguGw3eO/0u76pn+
XE382sB6DM8TWr01Vo2x4o/7OcesiwbM//BKrydKMrFytIQ0kjBBQ/BjexQNZA2D
Wp16Ai0ylqk9BwxCbYQsZRSolCjn/kb/Ds1cwhf0DWcQHCjJwV5AmfoCrvfuVkaa
pA3/by4gYgeihI4DXgm93NqXr+PsusRpzIOPtPg5ajP+M4En0X/jlwX2QiXc6cMZ
gwbZeGDCrodW2J2DNIkCFMwz8jNJnpyHzgAsvUDwyLcARyMsArFFGfGfbRe6zYm9
kfh5INNGuMeW3LjG7IKdfeFLdi5yooG5XRHjrxTOPQMj1T2YTszdrPWzq5CS7Tc+
7a42Fwp/R2vu6cEDOcB6zKvahqIXUON7IUGf9UuOXtIfbg6hCZgIeWn3E/g9PvgJ
vwa3+A8zQOvJGMvyyuTh8vuUrqX6awVZNgVp6n+D2iPVX0uOWeJ65IBFMRjX+Rid
kAFSxo31vf5ICzB97DEcVn+EJshaV2RheyLlocJ+tSP9GJe5mUwp/HQY8FtiBdIg
XUuzWJCXYZuF1jagnUNtLGjUDNXsjMT9GKFgFZ9/2jWIPRnE7PLKtmIrIqXtxJTi
`protect END_PROTECTED
