`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VI3jRPnz0+fHaYBrRY93BxED4R2CPFlw12UfB8v7WEK/76tm+7uEkfAD/cKo4OF2
lqTw2IeZrSH870xzA/EgmALawSIOhmBJQjt879jQNVc99+Wz7gocPcstuTMRKDie
YT4mIz80Nep4UBGlsazJa7OujvMViNHEXEaM0T2CwRZ+VrnM2DttzK1fF7dd4gMV
mLMFFuEmhftfJaD0alXJXNoTPyUYg6SU+uvAkp+ywaLE0ZClvDStVLWR5zVdj/Al
tnn4qv19ooZBXZT22u0x3Mz+C8zmfgrWYaENpjJ9e93TQb5fKSSPERA816H9ppSs
j+SusBQUv/z71E47tIMnSTyrynwzf7bXFWqyZnkP5c6C+hxaxBk9zotdG3X9m7uU
g6jS5FZYqdaAmiUmPANWEcpesKuepwqyi8KXbfoog8OzpSXyKM2RpRNhu8Bi2LFg
`protect END_PROTECTED
