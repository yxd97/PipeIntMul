`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e1dPcA+daY8VMX8QhbdhWLwgszMxaQHNt1KVdg1AQ7cMjJibRHKG8n1sZkKIFkFq
mO9ByQ0UzSOsQfSi9d+Forf840hyVldJumMPG/zGMlUTGQpz1i4A1H0drwOCxw73
HgvLDx5tPd4MMoSTEowhBhywr8EWOPRwMMzq7NlIoaHg/kfS8ZZwPwq07Bw4qCPH
bXIeSmxpMrT9pf8aZB5qH2ohgQD5TFNfLxtpYj91IH/iUyoS1VFV+FZmxQaFwtJE
eGX1miHe8sDseyVIKTosXQfxF2XvIFRpwJ6jQ4DNqUaCmgaux91fLbCs7m9RNfmI
nR5bgWVWHlHxVTsq46t1uNHyjPOHR9orzPB/Rp/DT4Si4MAAPO/r3q5rOHayF7YW
qyCovhT6WsHnqABMvB/7PMYreWo9eOV5A5XbcaDxuAwu3HlXcUMu5or2E17WxErV
Nwvc0xmcR9/QTT/ITyJouuJKmw25vTBdWWevWsv11tG6ra7iQd5ut4/cHHKEDiI7
`protect END_PROTECTED
