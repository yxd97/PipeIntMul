`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CRkmcS2S1a56Z2hFOwiwxhvh4SMH1HvFGk5l+ZbNQLxEcGy5IVffKyqisVT5oecM
ULC8WoL8XQlKOAegLtOpNL0WpSw4ATTRiL11dI5yDhCbIfk5mJBGXJ/ZU1bF/QdL
VUOBB6gVoUaajicFEisYruhH5qIOXM9ngCmEA5hDihUKIX6poY62ovwPKK63UwCy
BIOQZokWcSE4YNLx6223jR1Ue06n3Xedj86tJaQqpR276T9Lxr/kG0oSHHAZbC3x
X8Y7c9CvjsxbJcJeikQY0Hoi9gnpVyGeilvefzjq+RjRKi5QrhpzMWpAeb04b7dg
e2S0qV+fgdl6b90wEP72cS4P6uakv49qgNVAdBcZW9QNn9XvptYO7/gA3uNichYB
QLDt2ej6LHDG3ul8+pWEBlxlYHUQiz5JGdnbBmlkC2f220fW59DJW0dZqSdPi1CI
cTMjRXSZKImuPyPHsz8UfLuOvLsrTkErmhKJLBL5+MCf+tyzYOz2u0mITWo01p7f
gNvO6JYv0scBD8STgnzD6Ft+Hvqh5B1TOkZJ0QKOA4Ob8drtRg8pE4OhXb62yRpQ
1F+entmJUKgq9WJNclMQ66yv5LnoBUDfWq/bp3H/WMv1ZcPxrnViUjGP9VUdQ40q
Ah+5ved+1GfU4NjCM6VmWCuRyAT1U/WLOLH1CjmuFpc=
`protect END_PROTECTED
