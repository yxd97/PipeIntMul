`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9seLPc32Ba10/kk8XofEAJGy2l+FTN1a4xAtT6N62xgLp0pDzVLE/ofPj+1FTmU
ZI7r29w9LcfwA/bcQs3TMhhJz8+sec6NpQAELpPeAAa2PQM4kvf3pPYRQKYyplVH
SpJk1gdAqyUgJL8jzDuBEfQLOEcH1LWIUIx+NL3FGfx3FHRrTYUodeGnMBJOj+jo
OlYj0fnfC3NDvTce7d60c0wuvF5gVqanMTsDecIb61JQxRm571W7sJKQqc+fF6bK
sJS7OznrvgYxNWnQMK9EIGYrCIFNM2XmTIRC7PJn8lkAw/aS/rhYhCRYbWOhKxYS
EyxZu3iQYliZvFYC3UJabKv3hlquKTp5UVSE4/M3mtcw3/+ydRDP9YBBprPHdVgI
CYfjXEJ2AoRbpEkEBC3ozbM0Bmv+NECC/fDHkmEoJhw=
`protect END_PROTECTED
