`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ir+vr2I2Y9pyfDU/OpRlzRx45MPydYVFKq7QKDPn12ua1JEFZ7nptED0Dh9J8Ww
rky+O7+ENHL1j2GOieySSCgEodAkfLCGRAk679AmD9jlFMlIgICOFBgxJB2zp5+p
ze9nNbaLCA6ADg4ulCVjV1uk9amCPI9JNBiF9QK5hSrEEJnwQBjg3XKnMQnrXYZL
qNVzQiLAcDimT/9o4QBjQERZoUP6zTNtVQOJHPo7gnum99p57jPfEGC3o9sO8WKS
jOmoU2DQ576eztDos9eFYwaPq2HqiClLTiyU7VYlWS4FV+x0fhQ47h8zTsHcCIVZ
42mcFGN5Ly+9UDDKIoD4xX+ji+arMiT+Ask224k/XItLROEuLADvAEJlnm7gGCXr
/8K6r0Et7+bkyRm0XlH1cOEJU86hxOAyVHx+BmO9iY+/AHya0o8kFa1naIrKyHRa
CPQFFl0uU0m+kAKxF1qvqqees2idSVOyVG/O/TntGVeHq/zFhHpAFm8se5DjPELX
R3llBViMqpKZ5kJ8Azta1KlTq8ZM8fsJOLlBJZs4vy/Kj/OT6ItAY2tNBlXR020Z
D+otDj0mgmlKJROiFfsR4kFLw19DDJgyi4jtmDVnu+i2cFIxzbQaFcWLCxkWuZ/l
DCjOmIAo3Mjhs2rJfdTJWWFhIVpLAIfAPT4ndeD+JH59/tqS3uFDaFR8YKe7TpfH
sJPQ9fH0ZsNJ+1trAKMoDxdw2XoyJzTAamExD1ewibM1D2zNJ9yGD71IB+MJv0+E
8DBcJt1wnS+rIvRVQOWoo1ZF5dt27yz9/hVaC8+yzUOH6WWOzaOum7VWL0v/PgQp
HKg5Q9IaicT5oc2FzPOpIDbIqPvQi+9dfAx3ymyTGgzNsGKgxrZhM70e5BcGKjfV
MBcBh7fCBYehzzStrC1pN9Hl5PJiMxIUj+2O/OQ3QZvkAjJOjvqEYni0XHFRFmmK
UbfSqrbHrSKmEJAHjVv5VD8nxywXKEqdCWp6hM9TrCE8PS2p2OSSLaRaRZfpdN4e
HqxG7ymI4pfGOGEl/C1vWuFBBcnwoH+CKuBEp0rCcXHAJ8wphQwlftytxsSh/Hci
ES/dbZ4oJb9yCchoU4+upOq/4cV43PDMuZ7MYkosSahBx+eZbtpMTqOa2L5GRPLV
17cinCmTQH78xQGleuEMcg==
`protect END_PROTECTED
