`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AE4F1fQIP5WOFCVHpTxNQzVhqxQbWmVjDJ5Yiuga6pJsyOrlYGYL9P9Em1PBOtno
4nOL8N9e0f8bpqugqkNX7sE/b723yEONTj6OPaiX3eNyaZF4jXSzZDhtrWUWfglu
InVBkwqXQoChRrd4OMs/DaMtlV+CI5PkF5gTWbD6c7NjK5J+R4HTOYqJce9y/EI6
x0VjbGV2cainsiugKrig882kCEbq6ah7DELQ9uJGIbj44ZAwGMFQKJ4abT017COP
mRvXkPMfUvl/pMAv7zs884LpJPTC/0sfs/hd9kUur4eKHd1Zl2+Mj6Hd9vPhyyRx
RtnkaMKS75B7LYUGr2Jjq8+8Tqnxy1hgnfYPW1l8k5g=
`protect END_PROTECTED
