`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ChqdoyY9EGDVmbZQQaZs2Amty+KZEisBNDHnV3JFf3u3qnm8xAPDew41qRTI0Agt
8lBIs7osGCaiLn1BAcXA0ndVFY9MKMF5Dk3/ZGjF03J7HFK8Mu5riAz0GfhFD81z
MFBGHUcLTBxM7/1Q3XPjx1Y5nt2aQcdK0aPumgachJH+CmVws+RWaIyi2stFpTRx
DMMbzqzPSKMPQlSlFZS/k5t7LnwMojG7CweZTp7eieExS1Dd13t6cHKfRalfWxvo
9Wt5hiwoJmx0DEnYKkoVU2NXTBEEtOiVEb/YjuR9Of6lJwQVlBcZV8mU/xZyxK9R
6HuCN18hgbLHKGI16Cc6uJAT3x6PmufuATEsxDPofjx0it7j7Bv/5i6UbhYgb/s1
tvlDDjSk1mcRpt3Ha3BJae7fpxmRcWQs3lxoNKilWug3qX69geggGc6OmGpL6BW1
Xd9fjF+T8oKD+3FYIVVLLmmaBn3egM2bgv8lVGVbgJz7PcGTDi84HPj2abeJ1Gqv
`protect END_PROTECTED
