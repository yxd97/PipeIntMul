`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cuuGX6r3fuj0OM4d40jDM0Ikp6MER6Z80xmkYFxQa9XW1V1N3VlRmdlx6yB3dVyw
NGstN8SFW3KY+K25o2e4/P9squQ6a6FHbcJTepCxALMUIMNpmnapB108TwhS+W3A
cczufRKHpVPjQZWTUj+e6qLln2sdUgmFIF5qNQy8rAkxhEf2Ca6jRzdGJtO3IBty
yIBNN2fsMCOWfjXTzL+jpLPwAWmc336gZJ18NdTiBnR3fbXsnWoatu7jurngA1t+
s4OgVUSREw0n4M3357smG9dvFQIonxf9ad2A9LnymOX8xzq4ewAjB5FNkDafKhPh
F70TIZ6IJMT/TPawc8wZJlb65/z5mq6/5MCovvnnkI5Y8JROuyMN5zeE6DeTZvVE
5AhcS9ViJrfGF+MQsCLehS/YJxkCQZ3Uw8M2dq8/dZi5QePO+6R0NSwxdDZgsZRC
qiz6ROa150pVwglRGZROemnp40iEXoUUhVsgrw/BZTNqKkohwTko0UALKtfTkucN
lFNDLvjD0mjGTE6bv8bPbfHoVcg90p5Bem9Uu0Rb0s+JsG0QJ4d9pTSfDURVAYsQ
lDrI/VHgnfmpCN7YRRyrTgqoPIktCoBcDB2UISIeor91U5IM/OlO6AQTveP/Z1Rr
YEF9tvieBcbUV4ZDH6nLw+pmh393LzTer8RDhfv3E9GyMIGX71zyZ0xydb1l83Ek
sP4y5B7QpMRJFpf8HydcmXDqtBdusziGndVLz1C6GqW2INOB5yGL+fASvnNyKrkd
NEUOCw5anF+KhO8uFHS6eHci/3JLitOueVHP0R6Xzw/jl0ZDXFnNYIKfxnA2ik01
59FwTvbJor7cY03LyVQjnHWRYBj0hrfm+DPfeoZkvxDfSFS8DVwt5yEfHXBFW3wI
TaRO4trCfUxsu8tu23/GMCg8YtEc3jmlbTtfxJqk2pWa6YF0GGG4rmXl+rMNu0Sg
a25bRRLEApfiJ544Y1GpKlDYo+hy/1EOJ5qxuOtKsO/ie0ljy24CAIbZ6Q/bk4mr
tzFEEzVGbynX+TVHTkxhclLvJSBbaHV9Rkt3lalgL8zWYyb3IuN6ME9K0V+RGgc8
LdjCWTXkaU3aqGu5TQEPG5HlTyZ5ZUvQInfmUh1mRs6hU8yuaT/uUfq0xjQbS/2t
u3+oidkx28ZX9j6BLWbuHkHt2a7+8I3LjJ6cjRNiEDePIx/OqZv1l++DH3V6h2ma
ctZQDTQxcpDWsZWO0f/8HurHqmo8Vgf8yt76+DDedMriHSWkJE4GXiX+SfXb06DB
0ACnABT/y7zeaeKzBI5N7NYCLf5t+BtnOZViuM3BfJHEFSDGggAZ9Y2JucmCZNin
hiqohteh/RcqwUm+ey1Nr3EDFRuXsIzTjbIVh+ThiN+8ZEvTBMiDi0Ay1gV5akzy
Qv5jelq7lmuBjsOoCgumBBsOBt1DjuKPQgrBG5kjmhemXLZhHE2FJ0ss42+/i3Hw
wUMA01cvl9xkTVRw4KycP7hMF3OGucAxiAySx5FK5o5s1wb41P9ubD02md1o9vAB
jrnS52SiNRL3hPd0aZNqQ6Mh12PcwxVB6Zecjz6LaSPIYWHhzRBs32CiDcwn0DEf
SLj1M1WxrF9NunOtdnOTTupwtvkL17FnfgZb1z1D+qFjdpY9e1PNwW6lb9UQdetd
sBNqJp7kBm3AK3BvVknfZMgudBe283Cm9JLHOYV1SEjfaDa+Q+ZrUn65rU/XxZvJ
X5ihOlbLs7TQUYMEj/+3eRX4d/UOZ6L2VlXNtpC7WJ32lT06mpCsf3kDf5TM9ice
tnoB+G6zxQfDnVvrnL9kIbqnqw8MC8ZcbtufakV7A6dRglSMy3SldJ0OR5kubp4V
zQdfeYLcbJgYV1dOw9zle2EAF8Nd3e7YvhAvAiWHJ/blwgrbcnQ1qWQZ2wRa2wyO
cgHjk6Vt+b+Tke6kKHaHoW8FoaQUbluv6Ti2qAtxq4xvzxiKARnDXMa/nOK1rks4
bNIK6KJsAUxT8v3VlZ7KGfrRhvAfAOtkIdcUHK7aM5LRaf/HwhbL64w1HYa6On61
Q//7GFP02egIVaJE6C4jJS4lwFjfHrp4beWxIdBBLt50Xmpv+6jHUtzeu0LqEYqe
tdq9UCApYbE+2iYmzfi41gSkPtwEVheqy04ujk0l7hAybPn3sUCpLlAuO1YooEaR
yJNeA5od7oFD+T+7v+EzJQyeS/o3AGUvOGWXiaz5cR290DDNf5X3jGqO1oHSHzO+
ZFgW2nUj6BUHh4Mh8JKPoO0Mr1vp44AV0UrCjF/j7Cm8I9EREeoi9Z7TGww2lIeq
jK7Ptta449KQrxRNf/tpBw==
`protect END_PROTECTED
