`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+onspeXD7z8fSTV8hevmKuI9FZcRJcNRp/8Et1WbMfGqsmsl/i6DhN0w/mops7i
aBFnWdd4elPCSMIsZjLp16keRLzalDAfgzQl/qgMjoOGJp/MWYVZMHXTr6QHIXpe
mgRy4+X3krDVoll6Mo78Wbc2L33Z0J/Fph0mNT0K88YbRcfh5hgYDfvPLsLpgIVq
HEGBSLzYLItfPkl5YlE8Y4RMrb17l+XTK0LJWh/ogAzJiBBz//mX+EeDaBjaDaig
`protect END_PROTECTED
