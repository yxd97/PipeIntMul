`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xL5xNHTlKKV87mU6bHS3t4LB0SmrNSK/ozZSeI+OnXQ5EH/qtrGeV8quRM3Mpvcf
qc9a/VOS+pmUIFjx1Mu798HaNqNAcnzY2EQWV4EmKI7yM0XCKVBFEKBy6JacjSj3
wK/cYZuWsU+5bU/ybV0+soV4XV8ikDn3au9JcpFekosp2iGBjkmZC3RjaqCfsZyY
pqqL6HmgtWtk8Ds4henYzt0mKqWV8oKpPf1ooE+uzISBGI3zrh3Y/Yfn1HBWqkjF
/CoXlnPxN2V5GyOSvmH7SE+HGA5Ymsm4wWuzisp53PIf+SGleYaKGf5/Zu5/YqRB
aB2KsErOmIvD6NGPHh5K4JBo1TCOGUn3BgKgjPllWt1P3ViseaADhVmrOCbfiUdR
lqNkxKdNJRdQt9BDNtNZjLZG6FeLSJclyE6++hf0tlT3GdMisz2EDxf6po/wAG3T
bPg/ZwrzSi4Hboy+SHgcUcaaJNwVU7yJxvuiKwDZLsA=
`protect END_PROTECTED
