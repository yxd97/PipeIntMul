`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6WzEtryLuE5Z7nssGNQYVmyZjoYFjgrZITZJUAuOwZlHSdH9HdGUKFgUkx+gYO+6
uF7o5zyvOGnCIRujsnu8AwQWgh8Mvzpr+zXHUh2msfMUGlm+8l8ZpOXDtL+Pub0/
LF/E/aV7ui9y1SWX/ai+5fvmAOqdURKEt9rrYHXCI38naCF1RLOAVKLHQr3qP5h8
ojV/w6y6ya3m6Z1Zxmdd4yfjUn47BvSuHGxnmoJVNy4lGBH6du3pTR9CDuG/+S9X
8ymG27Al2s2g4+++DX0m2AjNaBx/F0VIH6HsAuKl2St4CGMGFMXxKLIRKkqiOH4k
dhSVefcO6Or/oYYUpXaQpFUaqCK3mkoEc0YbB6Xy4yU7HAVy3JsL3ew2tHpbzr1Z
`protect END_PROTECTED
