`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZeWHG60SFVBGAh/nzpn1NDuEfe1H2b/XNypibjqFBpRqAsMl319xinOlSykn9zs
o9c1n38ia8EaCMZKuAJJJMW8cPqSQnqbMDGNUktzV1lZ0H38izdPAcOVtHfPZ0hC
0EyGGHFM7fzHbn5K7ddVr6nju70tjAzDuy0Cdb1OFDWBee7XtGZy6TKWnJHnUoKk
3yunlDIlXE8/8UrN/PK8rh6DP/1b/PqSRaWGHaGkEP3j7YQs8IzZrUWhbNzSQczq
pvSA4JhawRcgwj+JwxC0qG5sShyoQ9A63qIQ+7+l6uuBwwwv5p9t3s/bvsG+yKN0
SPr3HwPQ1AaPubYYYd5NBLKiuTqdIiMADTQj2S+5mEejx25so1N2UMLtI8jjAlZc
ifm+uRXmfo0GtnOy4zyjl9519xV3SEX1QK5wqBvnWFWouFzXqQBrkV8ngpEg8Bml
ilc2qcvajUItnyrD6zM1z/qMzG1zMqGFZ6Ho6uughAUEYCjUq6rPhyFHihD3hALv
v9e9SDmv7WYmKo0cYyRAJMogIi468eFaPTYO8/TjpAo=
`protect END_PROTECTED
