`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+beLJHxAZ7vW/b1E2xlj63zFElDf8cAxEK6Yh/jkHGGGWrbI/MKPT9mkIiphSzUF
XYKnT7CwCD50HUK/G1P0SjogJgWu2YNUEmX6FuAAEXXvEWtEyk2zYUNumMabQG7b
sG2BX9ev9cG9M1scgDu4M0hOaKTFecJe5qThH/lsTA+JSFw+BoXezi200NPcQp10
zis6QiZ6hrgCbzW6eOk1/P9vaEcV4z4Cpo9ez9x/chcIDZEDoiQNgUj/lc+saB2y
ej4cMiNd1MphI7VN9htEB97PSbq4JlkTVDaH7ESJUdcfd6P6tiejAVwd09VDFKyA
1Kh4nvVBhRb+II2w0QwrkEetRbCBLBlFF6bHEKYs9x2xoflLxmOPunB7HEpd+ghG
H/Jh2etveQ0Wpzb2SuDcrg==
`protect END_PROTECTED
