`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A+dMD/NgcEO3ss6TWctu5hHQX1BBYDXuFufCCUOYzRqFvvioBFtBFwCacFCUPUp7
1cssQlKMQr1MfqUa3pv7Zfc/ZoMHEpO+iN2m9QCbO0K07tndYc9q1GlcJ6T4rf4M
G6gMs0oBKoRZ3nlDX/7mhuhFnsBsUI1g75k94ndiWbvbv67SNFMQ19HTu2K3a9uA
gLYvmpKoLxcrlmLwERywF7W1+25BRCXS2weYFWmIY6teZV2Dodkiw3bNuDjh1HSs
kpHkat262t1BxoFWIwnt6rSo61bSjPAAxlyYAtJnoK+ZCorq0EBbBa2EbxaplYyh
xrzqoNyaW8dYB9qpkiqR4i4Hnv9/j2Zs7a2rbPnHSvd/c2JujTnAYOGeVCIqrTg4
IPBv/sLvXTgjTCaKO9He+cXCaWSrUQkMjScfibKp0HXKZap3SmFAuGXZcbUYy0ed
8QF7L5RxaUeGq9y8Qqs+Gp42eM3IvFsgM2FeBtfWefxNgm4GAhtyW+tTrbBy65y1
OZrbU5PfewRDdmfGVXxI70QR5uN2PJ75p7Ye3+coOZXiFT8/o4uykMfNcQPM2Dzt
/ykkknH1rCG/ElKLukkavoH63foa1qkHfKAbI4oqnpKtqFOhliIiEhOhPCCplNWj
6ZiC85L3KKZpmaFl+KgE0fHf8ZXWjd0QGeC4bHd8zynWxnWx+7CTFXvN67Y+Pfj5
2ebZ0XMGYRZDDuOrX0qfrzJEnfYG1zPFCpZW2CE0eJ0AdYfrzpBPOyGKZZoSryqQ
rUvox1/n5J4bTffi3hrsGCF6KXN26qtg5yem97IhFCyhRG1NYvCjY3Y1oTwKXmhN
bLjbR80vpM2PQUzGf2UBxez+cRE8EPcsgVax7Gmk+j8qsVcM+MzOjUhLfQPph9xa
+8DgLgn8f/8HUUm7M5KPMaryyX6J7xQZ7wh0M1cX+xQAMkQ3aqmjMso/IGr1KSgS
lu3txB/1nWHXZVNx8rKsZWfjdR96olzwOGe9LZ3O1k2dj41o2JC0cd4Y/Vp/kOWW
/d86VJ3SBSEP6hp9IDrF2H7GXytlTbWm5gj+t3veUJQfeOt5CuSoAJvLHRJxLNof
hnqscke5xKYjtaoHzjpcKq20aQ7TXGDjMTgY6voriQk+Wi3Ux7gfRRbH49KTx05A
ZlwD50LOaxxwZKO0osjN8lLlhMt08HwGmYp6cEuO/J4MEqx2Y4QBT1ROZGEOrQns
t+EhVUqDHTvXllkAdtQcKCNQOEkVCK08dqU1Hs/Tqbu1Pxy4clxH2dz6dA3olxJQ
rDAqYZ0TZvydwFdvSYtLQmE6AGAdg0JnpPlL/mvHfGx0NrGOaA9ndUm9q4cDGtp+
LuHJFlgfxQ/fRwK+brnl/AdXSNFtIij6dHKJ75o5tmogOmt/1GTJc4ljulCo3dZ0
PtZ0pbMWK/vMmd4FPkkXuogVt/VvZ/TMEWHTaRXnpMNL1zGwfh6dmiQ4Q6oYbJsg
6y6S2JS0Qc801p+ux2eZDX88+2IZgj5RV9M/+p9oCRbXkS3+ZyleaVICHhX62vMV
0k2KasiuilA2WcoT4DdzFK0i3ziJooFjNu827+PrjUgQ9JuJYbRlp9cyQWoEjR0x
2tlysXCR+ySdVBZpGhpWULw2/ekdz1/qMjc9B3svhN0DpwfspEko8RdCmCTZzHnV
ZHX7PlHghyC6DGj40FAUHChLSRUPyO4GXkyoM8Ikz8YqEnzI9fYbYgM/VyvPaoe1
y1l97pR3/bqHeAW6TwvU/0Azam3/K+ytg7A/vwZ2HsjXjg7jcPOs/GOX03o0uT/5
KarVv6FJWeI8+xGp49KfPaTx+/PwN5RID1hg0Texj/HYUC4wkpeXTl4gcO+qEJ3/
bmam7ASdoUer+rIibXu8kj3dJC9TczGgBpERsMdXAqBJDhwgsj779qZg8SFGIt2W
pMHPpaE1ZJO5sGzh/OEUsS+BkSVZ9gZCUJgsBinZQnwMhs4gtHpEBd9cOzSEeVnv
egfQxq1gYSI28bemES/S47LngmLWQ4+sn096OcfzDQwoew2b0zneJ5oNddcNRXoP
jWR5BCP6v4T2r8t7rNVO/4OHz4Ilv9FuUefYsdBxjMeIkTFEhjD9tz8jezVV8LAN
3Ws4ET1yZse9jOlFhjJQEUHJvCAap/y0NeUgKydohIjg0HrJOcvtjBtm+aUOrJ65
V7rbJOGedqPMc4Mv0Tvtn5/O73P1gSlG6vMfUvku3pgr9ocGxHhz7N65fXD7B92X
8vRuJJV0nkHkpr9q5P/FoHpkFEmR+bcRUFoDrKzLuFvApMDd0EpeP1lYcj4I3Fys
y8ZxTBlpfRIVenzrpsPziq84ei/CFsgMN931B9XScVjFgPFVap2V2RqIgB0jlAy/
hlhhCD21U1VwFzcoRIAeDhqL7FmgWB5kLWY4KjL/zX678YS+d84bOzzkO1yEPq5W
m+3oGQr28zBCSBv1gyYryyvdt+o5PBWhNK46/RbSdNGsjhy4BrGNocltmlf7LV4l
G9qKu/bmv2FkEZYJvMusWCie59GcstrTbteChL3sADuBV8/Y9zK87S3f19s075Wn
1jvD/RbyB6ZGzPOXEUp8x+qV4MK4XmbXDA8s2naSBHZ+BGPSdJKqRsgr8VHgAaGj
LPC/unLbHkd2X7mcWBZtpgSKSYu5WfIE8+ZcDkAVPd15/Ui5y5xbEGXj+Ca/MIM+
1LuqRb5XSj9zzJCu/tNgm3N5tywEEYhHZL3CyMBD/+WxPullIFZlIzPWDvEuKHex
nfBI6n5OAM6pHIt/geeraKkF4mCCg9Ok29JJVumxgUlcSUHlG4NIamXUb3h7PhVk
EW9eW4+vP3EBfLchT8lox9rZ7C3VFvDXfVqeGnFAkqJX2TT9swcqNM15sLlY85x3
RFdsxTJID/tuEmYqVhIwVjW7SSaZcchfL03Qfg05lFijrZ0IjHB21QCxXSYBe3Pi
EZY00yN5gUoMfYe/SaVxIg7b6pnapwEq4nnCqNuJvnAbtenv5RTIZwohsMYU0bPQ
S+2oXUE0D+lK8LlxQ83jHa6vOMtHPsWSMR4QCtbt4h3LXuyxx6PeWAQ7dyEIVwer
IcVZlpdmiZvU172fFTr4lhY37OCQGxFhJfAHBAgyqQE4Xds63d8mrfc9Z+znM3Pl
Cx2x+v/XLDVX/SGOe/gRn5C5omqMMH4w/3p0hYslLVqxuFcalGEgGbKgX+Y4ul40
5NRywh2aqC4MijInkPQNIs2RORvmDQ8/uuMnDL6HAiXWhHKsuSTfkmu8AMs/a2C1
Op32/RMQagYaDB8wGCW4+FeNcJzu0q0rbiv2oR7iznh6gatL2aqcV2jdh63s2Eda
hcyzU3omUF+DhehdCDe9JTnCfxtX1i+Luos+hSaImf3u6yTRIiB35r5Z/LCZhRMb
2CmbEkkMgNiDJW4WiAbEjVygP7zh+x96G/KuARkA+qjOu+ssgO4toX4VbogypX2M
l+AkElGFdfAwi4fX3+bP+cOFbZurUn09KPw1cHHU/XJQmWE8vUdqCljVFbfbw7Z4
aiEbFbwftL8paLqU931g9PqzBqY4sOzyh+fILmCgm62L/eyGFSsep1t7Jd4Yzd80
8Ouy/KVyDqkHHXlacl1s+SS4yoBP8eXb+S22/Xsy5zR0g3DhUmWJqov8SxStXcga
qu9v0dNN76YQ47eV8vH4Nq1GRnkvS37SHfEpYGoqlGQ8hWo5cCIAvOqkGkUz+KbE
VSkj/5kSHE6KeBbifMZT/BGDeTkl1UQszBn52m6Qm0Eo/OTKkYW0xMjBqJX/GIQE
QFSd1aDc1q+IJNhG16a/XEH7X+e36KlXmKzDQUpEOzUnspBkLhfaMPsLN9WCDGqE
nyuSJId/ZhltUXo8likNXCv3FLqhkp5yvwOz9uJf5QQZuNQLcyUj4Mqm+CeBwLwb
1dskx4a3Ju5CE0o2Iizr9tlElzLh5xUAouDP+VMxLmNclChQfaARltZ6NxQCxswp
kXspCcVMKCWBIGgZUb89UpjkJgRm3YBPgkhxrHZQOUVgWQxb0rUW1FCoulWdOPG3
D9QqqxC695IjYsm4pxx6Ax/eMbhY1utZG8K6vvizrqE0H/IRsJ9CEtlVMNeim9Xm
qWQOiGFn15pxDw0eMH5LwcOYshHmuOSdz/8g1otTK3FLloDn3+wYTl1rtTFOUefO
SCRDJsnSusIpcj7A6NOfoyN7Nz6BmZ769NpghD4I3EHGwzLtRyxPj1X1GUFtEPVG
4k6bV1ZnZ48q9LQgnrD7X9kg+smccRKDaGkFz+GnTrJ+tzMpwyjZMX1RoAnKpIdC
z4FWVuKwTUEOQzEZPWsh92a6yWhjycyIIyAMepqUHKVGVToJDArhQyzM9yQYz6V+
40C2loagnGtb6LiB1efZQNXMZ7jhrySTuc3YMsioLuw8c3NNar0D1rqpjeD2Stby
3qf3F0U1/EK1mzyPj4aCX+iAxesxffg9vnkZUPum1h13QcFSQyDmIdANbf3VpyNH
e0z9JR3nbeswUtwRRxUjw+kMqkkXCKkE5j8KxGSAp206ANEZ5/bXj58cKnsLa9/C
hDd6BGNUNucMBzvmCgP6nl0imWoBOmwZAHqw/nZilDodNbu2oeJwvr5HXuOXIj28
OflJzzWPtHz6eb3+NkHS7gmpXXnGDr7ZlVCesXKGQ6leA7yOBYuEeWSp+UflcR0/
acRyytusC+0C90wyF0H5eI8DwSpr/JyRuvuTjh30BWxtakFaCM9DLlZX+Ts0vejO
+odS0wWm88NeVQg4V4gIwPcX40L3jGs4LOerw2AcHPaE5blWQX/9jO4nPaEdblmF
3CSF/yNF8tO6xihMSih3Be76C4cWJ3yAUdrm+TgrgIhc+Th//BFT8ghi999mMOJN
KKSptQ44ApcQLnT0HRIld/rUzxYsSTHZe4+Myb/082r5hBf6K751gWXiQppTocTl
loYgFw6POMEUF1NuKR8zBQIEalZRB45jaosEUqAg9n4dfQ0WrFx8+BGMigZWfVX8
zF8StBsVXHu0CfHVhKcFclwywtbazd/96vhXSJNTq4NZYuMqdoLy7uzlZA1L1MPU
W3B56hyjGhVxm92RrVRoQq1J2FMoecxS2jOj9dtpIgox4LTCpcssPE7fl9Q2orFV
3pW8+Rfy9Vy/edO3GOfLiDfHN+FXs25t9JcFfD2vw1E6HoGPzCdjsjDCfEI5Slwt
u//CLyU7dFU01PkHdwz0+p2b1tLYhvGYpytHQjvleh2HJXIthf39nj5rJNiuTSbp
hXvHliwROlbWcnI2LJHEeLZ5O07lLAT9r4SntwJZ3AQpE9I3DnCp45tOAyUlaKF2
tgB2eNl8wjQwL6a1S2FfWMgUFGiY9j/Iw/bm6f+ppMb4/hG+G0qmkfSXP115HxUt
wRu8xg0dgQ6rQT/eZhDcFEFsJElbG47Jj1cfeg1ERgHQX9z9yGBz2GUMnZRwtUZY
Cn53m0FJGNZ+wb2MTnE1QXyE0u/JJeDqmfKFg7t3b3bP7Zn47QnlDvWk+ZbLaLk3
Lf6d/OCE4hAvaWHEh0L9qiOBvpwwU4pGZ2lQLr5NMgYAsyMAohvDw+4SiN/sXlTf
BXHDw4xvODrHvDkS7aQJAqaHBdgFdlwWFDGIHB8Wid3eMDISweg8vU71Hncc1e0c
1ImJjSvYpuTd/8qzHXfS2/fKLsYW6Bbye2vvFMzqjBon3w8PPLMHIkAOgW3iWt99
3brczYNwRFX5FvYI/0b1VpaBPFqL4N+wkSjgD7inJHdQIilbXY90I6qYebyhIdYt
Y6iYVD5/Yzy+i0Tq+Y+A4UZjRs5Cjmy6+9c1j7HobpPfZvU/NFZWEjuK8ek1eA+D
ZpxWyeTR3IRSRnAuPTG2CDmf+ha2Wt3wZ86HZ9aHo+TaYtvVp7zft1zZjU6nJeUt
C4z+8L8YAOIlCj2G4xSM7HD425bhZ0ITu49C99VPpyM9N6dTFIhIiTaCYB7ybjf6
AzGNhlcHilWGQVmFvYK/ccUKa9OA24IxgJ3ycVUDl0jyFKNU/wrl/j7Rpq+fMXxF
WGduLxmO2326J1SR1e+DN2f5C4QRQ+xieUScGKvpZyZFsHNWutzcm95ZtICB0FJh
4UyS4hG3EihDOD3aZ/ijA8QInzTiArqAygaIKi/IQYeWzJJDThaoY5uNHRhs9b+7
66DsUI9ZXY1vmaXPi/Ld5sG3gzQdRkxrUBw9D1ppvCxApN/wrVzpSlFLPQkHQDoU
XOxY/S9vsDMvNua9OYV9mz9zSyRFDwyQtFpDAuQ/kygjxTcBgiWaBf4xa44plQNU
nQ066C1/EVxUBlYuFt3/NQzGaTpOnVIH5sauqtC1bT7WVIhB21slajgIGDsqP67y
RAVBGvLq5IRwwMX30Uf7Mb0P/WeHC6peAC/1FoUsS0W8CkGiM5AYl/2awkPdT+Mv
dzfghVwTkA9B8T53aWWuk0FqOWlF/xasvhjwUntYqSRKZmGne+xLkKzJpQHIW/4N
tBuQgkQBKQ3evFfH/sOWI63055BltsXONreDaypP6RUvZRn8UI/GeUc64/Wujixp
ossCdG6opJCFRBNm9/Sx+/rjohTdDl7lyJOwGRPsaJsv5gnm4kR8DfNS5KotiuJo
iFwX6w13DHSgUpx3gzEdK1c7NIzprx3BlFVovgfLCPo9i2jlbANp2qjd5V/MZpAL
maoPBq3T5kgKCFFRCWJQvgaLQOFVFHK3SSr8HKOQwWvCjMS3YL4pCQCeEjYpGhIz
pFJ/B47JEEOaD9Ph/xVL3Sk4lDvNtcN8UbzRStEKpVGc2/c6hkNicW0r+VfrE04o
sD+jnqGHAyEDkuhSfxgBU+J0B+bz7FmTdXZ4OPSu3o19QXlrZnRSlpRSA//NQWBe
f9hk5tmLRyNYJgxmZf9mHOKJbQoVVXQqBXI5ciIuj0I8dd6clZr2i56oOr4zjv9Q
McglHhkhu8wcv4UCoZg+6b7jTcrZvTqh2YRDsLomeEADIhLXIfjRLlv2k99ZcdC5
wNNwhNy1WlylZ/C01mbuDKBACsXUM9wM1PDwGVbOo8TK698YMruvuOr7pdDvuPAc
vnUCu+BqJ8eIr4H9voLIiyfZNVYsEdGkRFan2Nk/toC4x+UnRXSHmg+oV0y/K310
Wa0HYfY7GkvBRcAXXUjFoBCAmX93ryRKf+ixYKgN4V8QsPKiY1I6wmkcgTmmtyOh
fyy+tPDAvRSqkAoFgnnTcbGBePqE5akyw0hIxpuqySHtWsxmwXqAc3QHWO1k8n4P
bC8DhByj7iVDbayiBNpz977skZKGvkSpa+5dD4VzIowRZz+U7bs7qpiWp9zZdvSD
4z7jhK0oFV59mkGh+h131Lsk2jv38rvNe+FOahCfUn1W6/ORF+I8JOuF2quqjPbK
gdJxWU9vmfQXFsJrq2bj3zfExTfQN/xwgJGb6wP0t8CiIkaO1B3cE8VP73PDTRHx
qEEc6KHoHZ5vA29t7BBTBESNPeSqRhEmViRxdgNG7ubBHrihCiOmAwcNTw1uEQN9
zs0o0qRunZw2XT33ttwy/AZGT2iP6hAaP2aSp0/QugiFMAKQsCgDFxgWrZhndrAa
xEGVCuEOHBALbyjVPAzmJRHBBPN41QpL+4FtSfWSbTPCjY0SsLIj50gRxD7blMsZ
xbPYNqm91vWqHv05nGwqjTKpJpVmXCakEi6hy8JIAegh2mUhsi5ogXXaSKCz8bs+
osDvpwezX1oVlSbcYG19857fvxtuzHP8NMEGbE3tCiCHsec3KUDc4h4wdEl4A2tT
L0bl0F/J2PkUmtWUMWWelP+liMaw9Mp0yj/yNHPQtLa4Yfbu1WLQVvQsJPGeFdHF
B9r0EEZEqfaV4LmfzPIevoev4k4iNkFNd5Y2VoVMCbjYgPP+/ve43AhEizo2rJ34
+pL9N2hYQHwXsrtigdKP8rZfP7oc3MRoLdddAFYRFLLFniiIt90I+slQy0QLHGCV
l6aIunvsSC7YCVhjpi1J4Xm1HXNwf5Hx5SKZAkRik57ok3vcSuhd+AIikvSeObqM
+CZ9ZUasD04aD6TcUtUwo9vpiHIipbb/+0YZsABDC9zS0BeRftz40YvYLsbpc06r
MLU0wqUlem4tQ3Y9F1ngGeZA8087Eo0ZOfMBEIQpeDrY8vka6QJFOqLqoKRRfJB5
vZ1PM2yZg4oJ3d/dtkhos3N6qM6frF7SbzgdNesvmMH/6ekqc8vxoQM3XzL0v2a0
vxyq24LmQSruwofZd0z2NM1oKBcqu4eTaL6zjO3xNKh/0SL6jmj7lNazoQaU9FC9
MOBDyjdFC8kF4ux7foKGlZPpck34oWbSUq0Pce29U+d8/NcOiCefJCfAlxQgDKkm
t1EssRnMGGQsB6BtxGf5pbL5sfG9ATRdgZwH8X4st4m7nvXPtQYfXNXNh7xroavt
RNtGZ0oANguYBH719l2D6wyD8jyINtA6xTYPWM2X4dBlHZhkA0qVu+5Zwu9jQiR8
hJDANdctt625W4XK4bXAUQa6coK9PnOGwx2HqWtODUdPVGo4EDzwW4iScpOKbauv
7BhhxrzprewcjjKrqx5F7g5xx5CRo7s0PSriFGzbolO3nN4BStMLzWY0V3Bicqpm
evO42X6C1/JXdPXnpF3nRgTa40Xa1xGjNSRMAO3JMDxVtIPwz2gnz4Tm3hcVT80+
jCRNtWGL9csvhmhDAlAsdbyVfI2V1mlmVN48kJRMa7ocXBfYoWTGkWCHNWIkuwsl
AStzOVK3CiIMcZE/8PfuIr0cjEM4c2zVNfJMsihsINpJcnLbcs4So3neHVj3Fyq7
F5rMF1RvZx+msMEgx9V7D/xAU+y7uvP+od/heHmnMGTeMbM/KxdojkCYrz34NVif
2cpxCFnp7ZOjikrmC9SEx6I4JyyKdWHO8Dx+qewu9jpAhzM7zC0yAEvf8F8RYeC0
LwACfD7D4mjDhNAk9veD4bFFDTmvOYbKewALoqrIGqqZuZiINnvsu30uaRmXMDAs
70Z48jfKGbhk4Pai3CoQk5wXisoFcIzEX66vGgHHIf+Q9wI6nkJl93GjRQ1ARO2R
TSLHtajJv+Vuwh1WczzyNC9RlQp+d46YSvQTrKAN5E/p14cVMLU5o+r7P5n3AUom
GdB9rLErkKU87psJHdy5HxYGBZDFOXPHngA80NeObYvpxxEmYYk9nEhhftGfMmHf
eRVqMugTzDVLBXAFAUbGT03HKXB8/Lxph5M5VOWcvx1/Rn4NsS6GRpxTznEqMwBK
R95GXctgQlDOVx8Q7MqyFOszPqiW75pGfn6XvytlJ4AKjwcjhLZJCW4KDx8y1J3F
d6zuToe46+N2tGFUwIZ7aQ0hbrdnhA3s4UBwhIyu0BiPZ/ijaUAuAKo3B9HLzbXe
giQfrbPBhgz1+curQt4q0MNAHFyz/dVBSHgJFLQDJYcY9I6cAbv+G7avAjO4Mjkj
A5CDCPh6yr8HG6EEFcdmGbvfzkT/UNTGq1FmQKEfcMUpT41UnUdczjb3UvQD3NkR
g4Sxwnv4TDMQZ0pGhdCyM3iq49U5qPtHaTrK3JwIDNfG7lJ+3BsYq+Sok9hUI7tQ
RAhmDXlO+1WWK976ewWFuozm2B+nSdzvh/W/PNI0goAI46uRQk2J4E1cZJ/ApUN2
MHdNc9GI2cCPeol88jZifI6mB7/BQ8pa4j6OVbf9ExcneMmPfjGwSLgcYaME+33n
3feudrv346Z4hRBieTfs4Ki7VOgp4DRzjNInKnEyuCHL9j9lUObY5uuK1deV/rW3
kwjzvd0lQ/LfaET3zomeXouDRmQ/ZEwFgOomkNgaeof6UABpx2THH+/em+X6TPag
W1BxDxliU7VyoO8Wp0KPXvb01dZxJhTOduzu2lFgwkwHpPdpQX5AtBZcoywYuFac
kAgNRnsAbIHUWQProk3fmVU6Q5YJmDO+RaXzo5a+kpw0CB8/xwSK9SbxwKlffaw0
zrYtgXgyWHQ8puUczW2+TSg0c6avhXnI/RxDM/ig4DC7iIesZHSfpHbNQtH6XgMu
MDQvq2O8ax+onnIcquvqwn2NZMy0nJafwGdNsSGFyODNO6jyRIoPmOYmL/w8p5Ea
qkgK5jPXISaT8B3hmuCig1KInymCyykfYUUsqT4RXfz8mfggkeiORgzHf4MpDELY
gdVnlXfjIgqcNbgIyrBVawrvpXQ5pE5kFpiuBru4JkrdYklhuOhV7NDjkatGEpPr
pcNNq4ThGnT4f0qpOP7tjNCpUmpu06gdry1Ce7b0UA0xkL6gcNqrjk8tPt/9yiTM
EOPuJx7UVEly/jBR1r6jp2kkNVsmjWomfurtcJj0fqs8tCaGoY06Y3qdwYWUV2bT
gtfUpLzlfmvD9LC4UQ4DlilrJW8wm/oc/HKEheeDuQyqEI9pJXECC/YKCZeHR3qk
rf04zgQIZYRbGpHLBXJ2GoPjZbgBL+M+sQ5KUtPhDQmyxk0tUCALoQearyOMLfUM
IxtMPJJh7CYdcnHSB0302g0aJTf05GlrIt/EJwtFZA96igGl11QYLaOrTFvCWvVS
C/zDLJU57m9mh5TImbLuoplNe3X6YbYDs6sqhHXr68RDt69sHMNiP88LuhjhL/NV
I/pg+H/iHEYZLrDN5idL53fNxzDq843hzW4iaUD/bTDV8m2FKbf4CRb4qMJ88i6A
EVV/nV5XGcdudmILZwLburze3mSE4s+LAA6v38H10TTh91mqtUSc8kFBPULhRMw8
2Louc3d8yyOyvLpaYJcYFjlIjT3BvBnxunknrsJXj9phE5zuIxTOhTfxpuTxhxiY
NvLvtvn2RcyNpZ32pBq8sWq+ntEGVVNH6mjM/dcb8yTpS/JgeCxD3JGthvq95Qoq
TXa+eVK9oXq3+8huDABcpMUweZpdGTo1t8/PTibzd5An34r/T+qeQow+wjijJfcE
reEhAvjWadDkhZZGzz0hM2LVqFenacFmFHVFPSyBndpK5YXNQIy7wNqa3RTy2GDi
+wESCPv4X25PGlXe9a9QHgu81edho7PLqSFSBtDsrBZwKlyOyk8cQ7xnB/dMxNfS
NCVTTpN9Cv1+KmBib6WkdLzdqHe39qU62Uc6RgP8Rp/j6VJv62s5xDAEfEaDVlOE
ZSQMmoqXabSdmMYrqDU80PM1OoRArEcYbDn/g3M9oN2BKAo4z64AiSplpxiThlfc
GEA9RDV6ceL6qOLVF7rG3ZFLKk5+gG/GVctzL5fmcYV5HVnq1dSKNjieCBVWDhMq
WvprazYq8mkRiZ64zENbpnratoLZroSPyBHVAdydE9C8Z8C5yQlhcbkgJMcFFd4r
QYvCA+myQGOHywDu8cYMluRigPlsAUMz0+oYhPdsAWdbGfZS1NGTUykdgsKimQIA
C/Y0E6m0qsGsdXkcCckGkjkUYRTU2sCqgt+P1zZ01qoF898cpayjLoDq49zVPfcj
T5tQLNNtaNCtWhO23G1Qnaj/YNldoN+B3x1EQ+DNi4oAujX+ik6Biom+OooZsvu1
DK1sKr7kJYgEZkYJY77lAuJMfWM7DU0o2+g3eYz20WFxkXr9/0tFQYjN48RxPxe9
v2jmpCR914tQN1gGHIo3x84Yfaonb58yCxUDWvTT4cFCtOw0dIzMbA6BOTuTcfVS
y4Vod0pqcgi6sSjzgz9k4L47wvqgRaQrOgGEP8wVJ45UP3N8qS17KVZUfviZTl7i
A5uJOAjIBt17Pzhuj1Z9vjwCfrqq2L47ekVSOgCO81zWK3j1Oi4AEA4FvAaPYwKq
qaQ9hS8fi4sf+KHqY8kDI1J0pT7uQisSR5fqQtAC471ATR8AlH2Ua6au28H/65he
TkedHsCExtQzmIG+XqIhOSo69xXiwhXPiGCxG5s1rwYJIS0FOPMxLhyg1TK2pPXU
YdBKlvBCFVThClEeXTYz1VpS4j4/UUMBv99/sQxB4GC7pTRurghJZKDUQ8MQz3aD
QDYWixDUYhrv4Ph+Ap6ZVWOf9kj46D55WzscpFy6f2lqObaCMCkN1vosVXqlMiim
g0JZZ37oX5IdgTy5LO8epYO9H+vVV1ujHXxa7N9JC9PHSbX1ohN6B+js5Z8UbsYD
Au35pJxyRoy9t/oUNFlGgtIt+R9NYzWcLgNaopjS3l/EfAAUhvNc34+9hSimZ56i
OtE5Svv3He+1t7ocvxXWcVCX8fbTHMzf1wiRuZ4njex/iiOK42oLKn11bT1WTelB
kjH9X9U5ybkkL0tcVaZsFTpEPerHgGGbhJ4sF8OS8gjOz+/VhcOabVG0ZrdvoEo1
6H4QfQq/qAgTzK9twZKotnEbG19YdQeF/ZAcqqCkraMLqghVR0SLnPUxMKPYgoV0
m3VnJHa1qQWCjXp/Vaj8gd2ool+XWRBXk8cg3Z6dOHyuTLOnNoWuLExOSGs3FZcD
/g18AiWr2+Ld/N1SU65f07QNUIEEQDRQ9p4ohQWIGVAARoJxSeJT3Iu6I0zG8QUq
Q+fMWhSF4xf1bLcejnpAIywVMc2eTWrhG6roliU/12Eby9HteylNW++MM4g5f9QU
zf8EQsWX4janZXKAmVLXGNWxvGpHNwj0Fcg4Zjsfd/jf7SPl7ZAhullODoTssv9n
dfWSjEEjFk1kAt1dtKEncnToycnnFL2vjETljsa3yHqf+Q/IvmYRd5ujwuHalJDV
jGzL6ETNtyc978I+x3DTAIkdBc6a8V7HiFMC9PZnem2bzgft2ijCAX4T+odTBwgE
XFOFYorhRJNmTW6fIjf63DGc7/af//Ph60dOFP7RwveXi20JZdJIPG/cUzTjwdjo
c3wmFSWPOBH4k2LpNI2lsETHcDQhv7Y03qZLJXb4evV2+gigVjbbhwuEN+0GafDy
biVvfw7iXRugcHgL3ttei5rREmPRdRE7GS8+fKZ27zhdI4R/Y1TbI8sqYQ08wc89
zh0HDeCb8q0lnX+ozW920lEi5QSJ+sLKcap6cM8DZv7bmKBMGZf9CyeaOknRGEDW
zIPoeD3+0DWMIyljFpc3mpOr+iwr+tY4l6DaQwixnCAmvzYTV1dLeOFJ+XT8wXsI
3hqAmrWacw3YVDdQkF4JPxzAb2O9RIZTs/WGcMT/4ca2rbMgwdSBI3RhpWMRfjHW
TBdnBJPI1apjWVHyy8emysB40qU9kT/ddjrdMFe1OaKRBzAp3h/pKMCIMyEFjWHS
Sk+FFwuXa0vN/Umut2WKp/h5zvzDcvhac87Hv+Y94HzU6z/GdHUKvxEdVC9yWJk6
csqfxRF1x/qCYDS9QxILCN5O7oFobt3WbNuXpEWsnY0Kl2vE0kwjSPG3UJxBqDTo
f0PbplvQDxrfwYIANfRuTxECiAdSTmWkyd3LaFNpngEJkUxkWMbkNgFoeUGlkIZk
yrg6KRjKPX1yWOuOJ1B+LIv/sYjY3VcjYvMcfKP7wtM658tHrZCK7HA1RArhp6i7
IRIaqbeiie2IDyTGH0o9QK4P9NZnm8n4B7AzXCLX0b2q0z0qpbXINQwcS66mgCsL
Y467HhlCS7yArFT5b7elTc2t5fukiWTuQ5VqS7YLB2oBf2nY9oQ7bJX+H4hBWQ1g
aigNig6sPv6B1AkgNholV6zatVvrxmBMTufu7fWIKTd5f4ozBK5P31L7XVcfaxsa
O1yuk3CUskBzourDHxizh6bINhxGVA442+FxokyQt+KE3l+e0ujbO0BfRmwQwCEk
5X+ZCnwkv/2lAyUMW6Q1rgLtiU+CTbAVfzUIWBvXNs/Bkokt9QhrC99szWohR+BM
8L2Yd4wbRRxoZljgH+IBggdU5ldQGBsP9zlBcF5RAgeylqAhDr5I/szRikZbA1pk
dbh+xkOU6Hqly34q1NmWOSsug5bkeE5xdYTQGwqOpIlxFyqhVUxRuP9+vxMJyE3E
bCidQxajerXROALTJ6WVM8C9nX04ytnroRGNbHFGVem7Kshhfy8RS1523sjJcsQk
qQiPYf8W+KFT9Q60oWaRDAVXamGyM0V10vGMXxKqZqkmUPwyRndwxZxrpaABscTJ
6qX3dnmINeHo2U6Q5bMybfvY38i3L8kR0/dGNtYiUIAN1JwlONn9gy+f4NHHeoVf
PFmpldlYXpZbn+ya5KIjTpFQI8t3tITh9WnnBVpO8YNU7Hma7tdQQmVxEjpCIiHl
0BimU773lkdmGu1t0f6MZK+hczVZ1zNdc7AQkqKEzmruGfJ9k/pDKIZLd3Oavma1
aT7FGynio6wgx0lyZ/31tcONi3D3h+B0ABU+UAk/HdL8rXDs0mq1n7mhCFUkDu8u
zWPa0DJtLczoiubfDomeuSFtPuklWd9ktO+0Wg3Vnb6afK87fBAfuuN+vWVhJwdt
IXFn9ZrI3TXuVKDr1bQKY8APzulGc+Msh3i2/Abf7AgpOthLx3MXYEJEtU0og3hU
HoQT6ZPvxoUu1WdFgiiNyGuwzKOxxsWDNmtHXNdqzFroPaDvvxqrBLo1gm7BA7g4
pN4EIctdWcudg1ZyAJWzeiAVwKJCuhy5vjp2qubGV8xph3/0L7zKHSvvwQNZqAjp
mC+hodQfPrePa5r9yMal97w4rAyMIskzZ5Usp6CEyLVlN1oely2MaUwO46d4pfsn
zKiH/pA8XHWDMvTj2qB7O7kdG45SaDmDCCjXmQ7m1oDdmaHm/MHzfOhWI3/pYN0R
o/hNFZipw8RIxoiRwSr/JTrVqzLkK5NoJ8lb38aYHOyY5jml+V2yMvB2tm90mheq
81cC/iRluqKJ/pX4aWVECexeKtlULkmdrNwhLCyENYn2vwBU4ltv5vYmK+/hBnUb
bpoV+PxPJQ2Vap2t6/EH8F8+hTXn3nzSdFSFGiDaYvHocKakpISefMsSgf6Z61Ki
t6XAJzb1r8WpA6PAykXZfqN3get8/fvmX3/U4E3ba3VDVrr+oxPp4XVw36cydZOQ
Th3wBPRZDCFyI1EeQQz68yl/18FtjRgsnza7Z8iOkOljQ105YhTUKsSvuIb3OjX8
2cZFyz60ndYDwjA+Ml1i7W+a7ak+aFex69DuQ0Yf+n9Cz14JLivtybNYLKxAFV+b
pnojGtwimVHsjp1SuwjOavfXWu7KPNrB94cdw1WhuAgjhupMVJzvi0sw/f2IwvqK
Nhjq8uCt2Y2iC3mZRdwv0WjuA3kvrkhHx3KYue2E0g3yYU4ynmvcFam8D8MIzqBH
crFYEFRiSE38AOJxxU83NOem9pliGRTA+64u9odGAeE=
`protect END_PROTECTED
