`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k4+agU2r+Nvg/OqdzSd8OmR3c9vS+jNqRO2367MZ7Da/Jk6cNp2HhixmwGdnjQ+o
l+GsneGQea9tqbY0YQ+nBd5YjNgIzj4U5MKkddC/E0qtSZD6pEuXCkLeRvQ2n+s/
aOorZYZu8Dzofib0NisVSmmGOcCBUHNjQW+l4NaSd77cCkZLbB4snJOFmxJpvnOr
f38wfj9WQ/mDFcsM5ONqYU6w+5vxdGGedBd/jApjCbYZAvZ+guLUUU3+bGGyaMU5
p0XKIYuh8Wd5HppPl1tbvw==
`protect END_PROTECTED
