`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7zVqgEB2CDmSTYZprg4oJX0QNIgUAM6j0ekNYkeWaNCnS/lzj9c7xbOOTOwJrHZE
4rM4QqCRwy7y9aXE2cMLWp2wpcu0jpxGX7z6a8Jn0TgWSP41IqUjzrlesY+g4Jkq
M4qLWsFCEMk3lM8k30ImvpTZLHa/1OGJFvBv4e7PyoLVvok4ojlahsiGJC1LdkQf
A3Gr+iVeQOmpJh/eQRUIPvTh8SC1QZ5YTloQ39anNRxUjJI3psXTi1F2ZORp/fY2
uZHgCYGdX/t35fE1JzIhQX0cf3PHVPbjCAxiU/fivRnRY16gTVCXlJQJxrDhZqh/
xMHkJjtTziD8vHi/8TY1Kw==
`protect END_PROTECTED
