`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S1OcBIIp7huVcUJquVA/Z8Din0tmm9asfye669hV9mwswSVQA0tn0JcKaMuNBirQ
f+kh7lAnIcm7LUgrcykh26OQS8QKy2mD0FUPQT20tafp2gxAws5dc14u/LDykg3k
dizly/TR88FJPzMhv2yjRfTOU6I2iwCcf4btl/fuFRJSX0Nd76EleUAUS8h9zrE9
CgN0dDntYR9IDZ2MH9EHJrTQ9Oh7r8EHpDm2VB+ieenqq9QQ/bB4f1i9QvxdTFKc
N3tXK9P3bkPNJ0Fpq/WwQa6T2/z1Q8YsCLbC3o+0kdLhRYxZI/Mz3xsEu8TEbsJd
cYvKAlNEJtTA4Jvp/Qq4zeL7Lms1Jr2RhXw+PNeBJnLN7F3sJlJ7XSta6E26wdXC
MAqfBPLYGpB0JZL3o/U0JX4rWJF6wbDOTDI6TDVamPMzNqD19fmnKsOUs00PxSUH
ST1N9DCTKNw0Jvw36AyNHysSv9/t3jrn8UWKFYd1wYJHIaQyWAH+XYg4CNz8yKiG
JqBoGtZ76jqBG/QdQOui2WU0V2oUWL2nR4pMvo3f2xAyo9ZS/FCHDYI0jnhO+/dw
En8098zjmpBXDFmYMu83WWCT5H2ZcUIcn2ZRZFCpEN6cuHPRtQvY3ehcUSrtx80B
nc/uuUVXI7pQkVm6Dh1UUe1yBrEQ9BYyI1B9eQtFW5VOQvy2yAkiZ1DHys6Pg8GQ
TPTt7ipqPDFBb/9IZvoMjtuA0gXA2G+DkMpUA+wgTixpZyU1y9HHbqqbdyVEhRJP
mmLDtE3FJaF6K94c3krN6U0M3oT+zOLU1EC51+spp4cNHK81+W2Ih8NQgj/QbWWj
+eIMXjgkXwhX8fHnS1vmcDuwwvUlZmv8FIWi+cXHQFh/g841Ao1LZdVPyXYD7p8H
2TkAULLLiPS+5PuPEhORIJ10an9GQMevPW6YTcDszxAgawwIr9JmximzJR6yLcXZ
aaNyHbwWNe/3D31kZjc75gHawddfbDF379ZZyPQbsrPPRvCCRIIDrkYXTkblt/Is
Wt9VZZgDRPX7dYOxX2IZDER7WHvwEsUKd4sL4bakil1TU+r+1qQvEsE7PAMWRsZL
B8A6xm25Y0IXdVsvtzatVlO5ey3Ss6e0+DqvtlY9r7D4PFtB9vF1i0l11YVWUto2
zXQzgeTL8/EPuk8M7Z/RbCFrGrK8RO4aImOwkonq4y8DL1MF2Xt66/Fh1aDfibEH
9rc32zfjasyfseAVnepWn1mCO4ZH1jLb1JQmUAfaMBc=
`protect END_PROTECTED
