`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lvu2uhI7SPJ9LvVW9SL/HK22q6P4CenpKRNGwWp9uHCaNWomW2KUPLZCXawzsh96
OL9L5PscJ8P+4JfcKiWg0fwF3xfx12xNZas2992SVQFQi9TXzxMiEon/1U392Lnl
RvpZEzwohNhEcOfEtymzW6MCbyDzsPrukW/va+8ZahQZStyu14sjkmeETxpv8UIO
3VMmZuWLowiLMo2TrWokF8Xod3H87IIvVJ3osHbhlfLWa6BlHuiWJTYKfTgUHVch
YrmkevOsrPSTfEsA+ezClC64W6ZhIs+/h3yIdI3IFgl+gZXEFJaoTJATOqzUcBJ6
9U1WNfw5dK64I6udLwC/WIzCt6a4WLQLvzxER9CI/biSoEH9VE9L7tvOlLNdl73P
N//Zs0J/Z+bLM8TZAHkDH2AJkFFiAEbcBQFgDky9Yx8ejpw04WoKvA+vnzibFR0d
9YNWaQ4gyK9aE0f3l5mKzqdmr96vIk5euxEky5lMqeKB3lUKUZmwiTigy3scDj7C
NEF2Vyu3T0+klrvQK0Zpj0JreRPPneLd5VyuwZoaVmKIHVg5hnsaG2t7Aps1derE
ticotP/vRm3cW3xaYXjLN3bZcGYNyUJqXp+h+MR2+aI=
`protect END_PROTECTED
