`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1z9n2LzfSYIskTarP0WASs2nfxJ0QNDINgD1d8Vkly/0aOgxAE64VfvDgP4joXam
OlKhMRYd1hHDZg9sp/ZPQmIqJ1AzqcWGtXIsh8ptIM7CQSrv0Fda17fDdQjVofGs
eLlZ976SNQS8z7sdGPM+XyH98cE/UMpHSB6R8kJf6llN0DBZJyek9vYYJJDGux2C
fsLbJhP4SGUB2feFuuf+9YiX3BNqRhvg5ivyCGLBIcQaoZ2EfToELa6zW+jRIyV8
zhVjMPRn3gEzGiUeoIvPJBQnRoaXQDEc2yPuBYLhN4VJ3duXmy6SAgLwwkQJgjeU
VvyTE0M0JaruOppIS6UUaupjonx2ewKXhLnsj77HqQSDTFcR7AWT7MM2d6xLnETV
fUBYlTWe6BbBnDKtrxiOft7kLh1tD7VkkPmnTon4vCs=
`protect END_PROTECTED
