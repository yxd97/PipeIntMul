`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nMj+GrI0dY57pYM4NTdQLpSnUE+V54YT5VToevhkTGBrmKjy6lJPyQXIDcrIEk7v
VsOe8OU8wQHtbhYkdQNqJqujp3UiTiuTbSV/B5A0RDbWcSolTTyB9q2KRLYE6t+8
YqTfzNkgabOBLOgmT+tkMvyvuW+gJ4G5RaHXC2yK/TN7ZasK9X/Ub53Nuf9OaXRd
qpO4zb/1lUTrxJKGv+ZQ3nIhe68rPcdUh+GDpXX2bPshU76l4O6msKW9Je6Vv/TN
c5WuxePeZxu1jZ9ODLaKnIN+cGfmuQeDOsevPKRuytKrKsPrW3tH/OxMfg2huHYC
pmQD5xSteVnUzjtJ4oEwCd06IuNYOmAWk0lO0OJXkH8OjVZwKkCB3cqTi+EQ52l3
qvnZYu4beRURIJhycB6/F/9gOE0+folGfyFqC2BqtcpLxAQwpPVBKbfJ2QRQ8hR7
rJ3XENFS+bly175nY+YqBxhQNhx01vcrfjiYQ+YudAj+bYkUDiMrz/oyN+M2Z7ga
PUQ8XIbU5IzLrmy56E9xrA==
`protect END_PROTECTED
