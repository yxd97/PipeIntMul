`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rztU3xrQ1gArJqdoQX2P7td8FFnrIZhv5QhHxB+/i+zCSsddZowpvN1f3rPXbiYc
5/MXIUfdSbeFAbzfAtKOfh6vcL9dO8WclsCClCX0i77IHjx8XYwqm4J1AIiozzr3
brY3UrsA+q6gTyp50b14+YGQLJoAaf5PCm4pExLcTAg1JBVBhyyNbs4S56YnZWh0
zwDfSWyo2WW4iOk+Ok7SgAj7aEPkzS6PvaWYWLwirSA6w6ikclZfd/r9nEtVjUJ9
hcJtTeb/LX+ZK2ZXA/W4tA==
`protect END_PROTECTED
