`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fcd9eZ8R+0QsBcUABCS+HnI+AA5c8BaxggkZ0XZPesPYoTiZ1p2q90a0JJ83wtem
mqeDp0EQ1YvT1HK/y5oLy/qeIixFUUiLGn4J+e6Z+JMcqHxNhJFy3ok8hCS+0Ohu
mmfpJkj76wmpE1zykpRV16K4gV1MHLCHOaHX2EKi7Wv14YSwn2AEg+0Of1HRM9Xj
8LOO3n5TQH3ZPtPO2JVIttKo1BjTAL2BbQHKM/DK4OZNKCeQOWBC199QvbgkmrCW
GBuKVM3Cl7qVFHxdYRiIY4YqKeDFWAMiXzdiFy2FsqH8sQCpChxwwDjb7vBcOWbN
+OMp+VVEuRDE9k0koUC+mppRjO3XhLnmaVCqelh/TQmPv+eSgFv+JJWyWCIascPJ
jCDavrSD8aFaBBg304tT/0eJvajZvC4EJMfIctU6fSdR0S6fC7S2TKnf48wn25tD
AG426DoenwuxKQyQQUB/xtxTwdy1ErLB/e4uIhF52AWmdWg8OqzysFf06gNO2hT4
IrcnkUTE4op3noR+3H3gL34/gq+BK/tfX7CnZQSTMubxU4XkK+kjfpehmOOJV+fr
dm7COaQsIs7//GfmKAm8brQrREl+kb3vPWSBi0J1rarjny3H93cPfK4E7ngqBFwM
K+rsTw3MOt5U+2QR7Yqt8hH+g5HWPfoVTOuU7zHx50y0znon1OQHd+d52tyd/IgF
964KQWAo/evT+xjHp0NR0DmJS8ZXVfy1hv/rA5kBaNhUCVWa2pOjWUPppOQBU/ms
zqmhuo7vzy7Fjw1+xJbiXkKnbUHXv9pUnj5fCXVuBuDtbmFX1UYR/kVJDytWhdjb
SzVJNjyAdi+vk6oz0Il4+OudHzCVVgR5E8vQB0iLpex4u6VAT3jUeQgQKdOM5lZw
au0BdbzuevHPuOH6e4pHFYqGp9K7pRgovz5+JrGUw9CiF+nHNcIwzDVeEbS2lzG8
X2mftwrFoMMLZUilCAApNr4A8lgkUPkULywc4r5lr39WFM5DIqU6Xggbwv4njL+C
NlqyAjMreUvpWK6Gul+P2S5zc3mDiU2MaIGLLriomowTML8s0Z5KZXvQ5edvgI9A
HB6OY0Qz+P9HFRRr0djQ7N2hHugdxPxu8+KLoeP7UXLpsQK8KSkHI7S5pKSO3JHz
wsfPIq0iJJOaMoASsZJeqmT1Hu4d+qWU6MAvGew0dWslCdMQBc0ufQtg2eTeWB8h
B46KP/ZcJH7r33kjmGSPYOmlOkWPyYEBbK92fCoaks2X89fQFGOhI028oqRaMaDA
RmfnYRJVwxqlKvYX3SEwjoCCk5/dzw7h1WDyH9M/zuVD7BpoSJbZa/MR7T82yBbT
8pOhBxi/9oP7B5XMl/S19bYMPdrGguZJ+GATbKkUHTPh+RSNbYV73AUV/B/WplTM
UeVz0qmCAIyQEw0ClZ557sZjRGRxpKt9ufFwudbYkSmFnxGae8do84HvEp12bNRW
XgilCLayJY/AwYvvE1EOCDQ4eWKOjWgGJRtPgU4TsezeANJPyQ470Xjx/ZrOUdMA
NCRPevFRW6JYTUw7RXJiA9BivDbCz5FpkSvozPv06TTW5yNKDBs4nrBLE8/CA9R/
FlojJmk/mrNgonPOqUZ5VVE11CF+OItA+Ng4t1rjj9eo5L6Tj/zxh9Pmqw4L+TwU
WOkCesqRn1pRqq+aL6L4RiLys6jk0oSCqFGLjRHJNoAF5KQAKqrXQU1XHIwZ1WkR
sVWwaBPwFLhWLyUpXZyjlnYkOevyz6zg+kuT444mPHNFmHorJZ+4EdSgzTJkzy4G
ghpaHqqETDoLZwY2KTZlm/pD3ZrYP6aPNA5oXqDtT24qAD9XXFF44hZ2z63e26V2
D7bnxeTcLkOAKGBeGt1hSTTckBj3doqOTYJfp3SZDbHuoQqIkJ/MIlK5DN8oCqaE
FiEKH0qCaC8cgG9Yl4tR72ItFKfFCNrtshDy0XAUsY8RcfFlfmvrG1a74KhwcGGv
3ueEo0aB5GaSU1c4Iv5cuDDqtX/ySfXl28PFOiL8ru+f/T5tCX7Y0WvfblJO/RD6
tKE7b0EoJmnxcJkKy8d0xb6p2BU5/QFeSsw6CIKEjjckt0U4zt4vQ/E5wYfOfFTn
Yb0VLLAmg5M8XI0xLC+0IMGZqlgKevKhXTudaft2rGRvQAzAewTB9DfYhhx5UFt4
qyHbnTYYBGmY2Xe0A0QjY50SJQifB5kVXJ5msFqGlrjjg76SRUK0SdK+hb+TjEFB
PReJZTt6qLVhpezF5cSnW1WArAVdujnFdbV/2SKGp1tM8rjQe4/aOAB04a+PMQ3S
H27H0Hwql+54CpebSOM/1whc6z45LW4Q3A8iIiPWHlddpkfmJaBfuEzzOcxnDzPk
La4hnKu+O8SzgI5A/kP0TOFdS5b4NVJ25+EsGMfvyaMGqiVr9Tcy+VMiIHlgVwRP
Q0ZGxfSDPIl1LZ9OTYzXfE/BndrsUVMC2h9RrUTCkVCuH/IUdfKwzzgX+jhPSko6
qN4qMI/4RVIyEHMRM+7P+Eq4tdTP/guWPD9ak5V4pAFJ8KYNYU9ZiYKfIOCgQBQ7
1OgDrfDgF7lLpS5WxIL1z3OZLx3uQ9iZHyHCEoEXLVM3d3IcLvSfeDbSxpk6CXFt
9X2pH0U221X1hOkgAwEEuIHxuffzjA1FvdTVRxscYytt2BPDs6F2/RD4XLD2di6j
ZFBbR0ZAMVMZjqUC8ja3a1Bd9d2BalfhcEw1pOTkDAyA7fNKzO5zOB6PHEdmi6Ks
rZxqnEYR9zUA9ijBmoNDep7zxylxBR1ghRzCMRJxyfio+dW02FP7sTOt0p3TcjmE
I6QahDUZitbv5mqwMn6RHuyS9Z7m9krLWmCs7JXAJnQ6/lWQKcEoCdrtnn4vA/0m
G3yQY3AVexMb4IndovHyoGRqdSdhjKtgMO39eBR7k2jUt1b+wlzyzcehy8MjI6sb
hz3NaTQC+k/DecOiImh6GutUPPDPi+w+B0R8gGYmipaGflzGmrTSOCvnrYVWX2YV
5ESkB7mUwBo+YO8mDv7X0g==
`protect END_PROTECTED
