`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VsxExFnpwHAPiThw1QxMg8tY3haQva3aOpFp4Jb2rSGyCrG60kQ7EAiY021NSyRL
zN1fGPJcUHW8hqMvapmWKr08vaTbFfT81e7soST2sPV0sZLDHIxia7jZXgZj7ymc
3yZ//i/Mz+BVhFiaO+TvmwJRmrBDFOK0Q2h9rqK1v+e+t4BtN3cl7/xyO/JQ4juu
LYkho61uWuvXlLhbv/Iry+yNZEoJsRbtAuyG0MvzRzzIAz62iUQjKq6T3g88WC+R
51TLwVJ30X0NcZtMbXu+DhCpoiPSjk+r4MEavyzX1WVtNUbWX1UjozHegH6E+nwo
0Q46m/B36t3vzLKEjIORew==
`protect END_PROTECTED
