`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0jYZwfeOIUIeqvz2jQnhqR7tpCSK89FnNmIeyFx0NOjKxDs+CY24Zjmn2N87M1KX
tnd7Asct+1X2lo4tT5AzE8pfCPMCz6iOXMOrDkYR+vghpEZ0CUPd5vPFpFHZRmpr
gEhP7So5+ObEAXjgDnsmEDlNWloD0XByGc8g0hnf2wpWWArL6jMjfFkfEIbPjglV
Jbn+htMDqjQViNMCdBRvTyKFnJG/9sQrBgQ2Cx/8Emtsd/8wOGJl0gYrifPRz49u
2zg9Ff+1sfU4XnsTdAJyYvrhuJsTi0jtayT4/O+aPXLOnkk6pxeB4rZJgW4JRCLn
8OJWNfZet/eEZDCiPXo9xdsNfn7HNRfCQUA1vLQL/n8oTwYH0lFRBw17QMmBR5fG
`protect END_PROTECTED
