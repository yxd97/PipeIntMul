`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afLLKzQ2zuFy3cWZDb3klOuD5w3wSEKC61ZA2Cfao/LwlKeSuLiY3Lab2VPAsVqL
CI+yG5LGcxvoKsn7NgpkjGdsWVOLpN3pt61jaT/D6v3zylv4F410mPQo/N6Qhdn+
4Sa6ksvl2Jc5gnIfJckEWShoSzxlg/IgyqGPumfPQwBm2XBGAGSgMrPUVyFrrtkj
P1ZR0uIw8S0clcVP42rjRWXOp7rPZgVxPihTEfdEWmbrML3DHMwLnk+ZB4+tNxB6
gBcDb32cS9RB6MlO+k0ZpzKiWp0AsdUHzvvA1sdP+G2sUW+LU4eEmZsz9bfc9YLu
rdw4wO5bsNMO4B+A6jR3RJnlPVgeid3ekMvs3OMWUVn8cgRpNWnef6br/TwvAuy8
7Xa/lqH8+fLsJSgvfr6N2BNvKlvWEluPgstq7Ptndwwolo+BPoy9szf3uq12N6DQ
dCQD23ah+i6llrShVoa+fettOf9HcEUCn5NBjjY2bUs3kEQNYdme6etf2XjZkpMo
JI7U3vPP6+G9v9S3yX8SJNKWNGXeN4XHUdkrqSOcUWUMH+3CaSPkbAeHSEDYlDA9
7Y97XUcMGVULc4dqOzzcZOZjJdC8S9SAK+DVJ3MglLR5jtFqhjQgBGf3eHTx8IMd
3gLapiPZ+C/8b2TxthVBh3TKfOW40W7LWGi8yBDyYfhsEXJj2Z3wf8O0ldlxDSxy
apfWVRQu+ZG6I6kSiSbsu7Cwn8UnUg7IsB/IWUvq6H+BDvRa0JXKhhmYDDtOCw7N
sr10Ly0yAtX9GDaAIXheyL6yOLx3tVHSJ3PtNEaFXOeQff32J6uLDsuaUFFVJsh8
4BXL2B1lSwmsGcgBFO6ISG6rlOuZBEXz+v/B9N3ijoAEp/67iuPBeYUmveE3o1Iy
yZA29GtZA67ozqnwEhQ5xO6u9wfpdV4Us0+3OXQZNuGXNd4t8DCsquxmai065Yrq
ZFzhg3/SSFIgChTj2ZmsQftUfencE0ElycvGiT8BpfgLAdkwUR+aFYTLLEWc5Dlb
+PXqjXPidH8FxDqGrHRsTUUTkgnV8iw81U17yrihclMnazELVr27YxOMkahk5qHh
XCUjfaPyxV/tFyXQZtofZaG5WhA21h+FH0SOzdGMDYox7w4IwlMuLT/UKDFocsE3
WA9nhDW8UTA1dI8dE8aWi+MmoX+E7Dzfl/QvHuScrf81P9bbbIIWOrJgNRkEIDTH
TTvbYJ3ktopl8Bg1x8aF8HBIvAPFdSqTPC3G2VYPsE/d6aFKvB8mefkSD5AWAZkT
0k6I5VIU9qqKGMpM0SOEREIlcrgU0FwqrG8/Sk/wfdA1l9b0IS9M8/Ua/GbURqG4
1g9gQx1WEobzzB/MJ8k97gHy1QcZRwnIBhK9+zlSp7h2nr+mDoh4fOeas51CqLaY
uRLadvHxuCTadeQjJidverp/i39b5SFAAG3su/ntUvaV5VxjzDKL0x/ZzGdqhFZ2
JoG9p07/hnvd2TO0QJyzyQ==
`protect END_PROTECTED
