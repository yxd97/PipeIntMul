`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XS3zW6f5HcxOO5n2p6YgKZKBrjlnVNX+SbskuUavbQBZ08tKdK3WfO7/CqsUtEG5
MR9H5+FWqvyQlV72Qo3NGxsxRkj358UYStmTKt3+PRWmsObWJUVViZ3xzRI/78uE
54w1qXTr2sQblSPcBvtfQFtftXNJTKxF9BPhB5bYr8NcG5KLf9Kve1Jc5XfmqOQa
gfeCC/TQzSXXnlA48E/YnHt/E58WRsYZbdtOJT7FLqXh8ZTAOKjqUbY0A+7hPNzq
6bbFKCqY4eWecxxJaACF21i8prdcNJ1NHB94phVvDohaq8+rtPhv/LYLif7jQIy6
DZlUZexRrduPyQq99caSSN0Trq9rRuT4d1+YUcUx0DJwUeFWJ5KqiYjm83OeY2aM
vZwZiqIHRGsBvXeKO1uStIgSD789KW3mxQgY2OMBHCsXYAJkt0LKtQeo08Auz5g4
r39YDADg521azf5nabTNI9IQ3DBFRR6GOLc/+3CtaNj42vU0fv3mjnSuAGOdGRCi
ye3XhZNJLJdUu5f2OuG6+cuuGOruhsKBNkVyYHVmeOm4s50KRZTt8rs1z93hHup7
8reRGEQUVmksxa552dsYAqjfpx5Kbvv/+DfneP6LAyGjNCG+eqRw8FKuq6sSOn2k
UExUMc0C3QrCY9ZMRfB01iCO+PdHOx4X5Du1rUDJMgX/8Dqh8zqTPqbYLKuH0DPm
0LE2td5BKzRz90d99Hj6nKJnljjlYf27C/KCFz4ECEjGi/NF7elWSRaMaGs0iYpZ
7tZtjykLL7IM+/CO6tsaBswTGvC1SykV2VppYyAEGSdndPDt08vHtcF9FI2aLMUK
Jwo6TMJm82lQuPfYkW8AwUagzDRbrchwNZ5NYbGI59sDU0y2097BW9KCNunnAGUp
yPvQ9f6T6bQPWl25HAVN48DPYndL3ESIEhRtS2m66WVMvhXrcHVkQqunIFyT90A+
UYD8uOCPC1ClioV3Y+D4hmU9Vf2EFW95Z2uyDJQOkPqRCXzdp6SB/Tp6e1Enaaav
sm/Hx03mURB2knolV5UScF+dBOF+Ka52e+UtHxv3mNikff8+L3xbaJKMuyk2vUyY
1LGGtiF3e1yr5WkSg1OLiXrUUpZAmPA2+h4ydBxTqXdgsnjfUjbyWZYjjXSlRtJw
bJU7zr9zUnDu/xVPdDxaJvp6yqIDXlJfBz4ebCSOtgrKs+W/+Ny1Ub6jn9y1mUWK
Zx5ONrKhnSixtHl8sYk2+XP9DVTwTMTRGq30D8K+4imOLOi8F3XzTvBXI1ZxgvlF
LP8K1TkT+saECR1pkGOhY2iTjB0ehu6fpesuU0v3ahlZ1yAyRerOCvLvVfioQy9Z
yCvFjlhoG5ZA6xnLTDbC4fKts2fWmt9vrQUdNB6+6oDt3GeAHNwMzQTGRTwYyUkl
Cuy3l5brcKeodGqFY0hhTA==
`protect END_PROTECTED
