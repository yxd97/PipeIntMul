`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWfwOFMCz1DGoljlxaDE5mC4wwoNQMZIpexgtItCbjxMMCJZYVoD3Z1K13qxvq+9
oGt++wqJphu6AnaVafesggHZ024mm1nJoB/sIBLdmV4fy7PJuMsweORU25CwgMo5
vA8AGEcDkFYUtIoofstdsSnEw6M8X4ljOqiFIghHtoUVqZW6ZAADWqx0xJhuFXLv
9DtrdCIV12tQtqMphTcszeCa/bOt8QipLSvtQf/eoY7FZNdH1BmIbIFnkIOeG4DX
FOqlGOM9WQKXQYwAULzuSvDsoLFcY2lhdqzOhLgOmDHqGNf+aToGQ1uDfKm24Eom
LWGfnUjJhM5BfIE5kBM+uA==
`protect END_PROTECTED
