`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z+8O4HFByvnKdf3wLS85Tu1m3lUrMhBtLbLokpQCPVq9EfcP6MUdDXvctH8KFlCa
pkmxW5s5w8VDoEkzZ6jBWc57TUdTFKsTt+XAFvmmKDLDTayikEvyihu+WS40Sb5J
aR/YLMff/40jZHKEmYDiqk4slCS/aShTvwYdBlSZFt0tIOOACLXUg4IQhwUKdA27
b8OW2eKEyGyCAXQnPkzBytovJIz45dG8ymYkAF9n6VfiAlYejnXwYFmiN+jsiHY+
`protect END_PROTECTED
