`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WAh+vH6oBcxVDHOWopy/0KV02ZpP17AcaLT5vByENHXJcxc+ytMNnSQhq4SHu1cv
vv9gRYEGJ8WRX9iKepWtsQm27nbmS2Idck/o5WvvnYeu0VVK/7mw25d3hV6ytZRj
H+E8ywg21fFhgPCtgfPiRw7Q5+xnUw5rOwu6Y5Uq8UcZ2xrpVe8KqCzkNbxjtmIh
YZBpA6rpgxlKCnLlRnS9A4XZHkuMbd37i/385eI2QYSTEAt2SbvTKoIdngeb8Fot
NdC3bpGmILCvJddSfdLufEny+UZ1ICtDcgQbi/rjiGXZsUry3slhKna9lWg3L6fe
tTBxoaB3Uks/4GqLHGeWO2nSBU89rXini08xWSR9DL/Ufu4/LbNZsLBmp9SCMc4F
MunQcRmtAiSo8RTC90VZLdYAQoYnFk5ypFt7myWX8cyE78gozbWmbUxcDnDJwNMY
ZsWeb/+jvnsbullvLYhjSITXtJHf8Xa7h5WHs4nBLOStHrABOgQaVc62HYiGUklX
Bf5eri4evMJfqS10QFFtNJ3E5x80NdNNH+QILNQp0VoABEs4TEUUmpPik+pLyBui
0n2En7RpI90JeVFdGSJ3+WVzeY7plk9f8t8waqgUac0CYTcFcJoelYBzcRaNMfG5
+8Id60sl6LakiAhc/WGXlup2GRvfcZIraVkGDtucu/VaOt4YqiqFVNvtwYsNoCTZ
OyoAkIGWz51xwlwgbF69Ai8QkvI9Rd+RR1m/iGYewvk936k4f3szpc35sqACamJg
mYvkhsn3/1Kz+V0mNfU5mZvdlT0hXqBpcz5GExrwZV9lmFH0QcEX2SdIz9QobuKt
sfOgptGq1IAYgjFhZHbkSVjClNr7BlbWOBz6Df3RC3klt0kzyZ0I41PQripasXmL
3MFsCi3OimaMCGD639D17n7i/0He6mj9SWd3f7c4NE+l/6fqDh+fKsBO1vnI8MfZ
Gh3xSsbSvP5HnHOWyR56iV9efTFuVvatAcBFa3VUE3ZsXzH3GKH6xzHBOyCHI8GU
TQF/oRxZY+8Y+aTlILV9GJ+T+mCMb07OfMHYJ/sARe17I1O8cNzXmJbs1BcGD216
o8qShXFtRQeRMOC0jEU0CPb/eclBBJUklglz2GB4hTmzQmO4i4TuPbW49aHN9lyc
Uf1/4y1HfOzWf6ZTF6UPmoOStzDIP9j8sJzD4PNTwvEp07cQfApa0F//dOiaNWUY
`protect END_PROTECTED
