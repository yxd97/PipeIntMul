`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W34yUbQjXhGbZSva0MunEU4iDDRR4i1TEIFpzMcUMl8mUYqLHxR6omiNEfMJo+Qw
5FPup7qgsnObumuo9woRF62CO0H5mEJY245px1gUBgjksgXbLyL5o3f3dcfsJV90
yEZEgABf7aHZI2Kh/gVRjAVz9vbFnu+mp0dBxvd6WxNsUa9uOLpbb447sAcNJWpv
xhcIMbyDSlG+j5L/d4vhteTdrXcbyNt9e6ld2enAg00LAaFBJGlx3C/z+hSl0F01
G7NSUhJWlfYrUXcCrcgRKsWS8WAx7JUj3MbTazwqRGD1rYtIFd4etQgwgGgvBf/2
JOcq+Fegc5ojrjSiIgBLfw==
`protect END_PROTECTED
