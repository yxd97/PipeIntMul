`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EyihujHMUdtzJ3+Te9EYL4gireeOtZScKiV23iruxZPkz5kPC0KZKHqqIXWd0eSR
HEkNloZyXZYrlguKgTPqAL3oqkk412ZV4e28WbmdAZIHtcWYg4Rvsrg6fApSoQkz
7zBW3IXBD4m5zMW5a1M9odtgwCh19HxzuRJFzRU/BGeUPC1ZO4dLO0zWkCZRWnNZ
VQgVWwiEVgut6cHD1YEk24A+PJfI8iykG0R+WJZYevN0msCAv0XBSQKrTXfg609T
lrW3Ajl9hCYoLdG/OVOxQKCeERLzLgJsWImxRAJ4yA34mlvc8yyCrjLxmIHCvpQq
IGk+oJwssrPCIGG4ZyaEcibI1FNY2n5B/iAWN5ODutUljUUlJSXnqHbQoR03IZ0/
79vULxjNxmukMaxo2yJ3/REnociHEPTmplDhy3t1ju0pDwvVzAKc9q0VcRb38Aqh
`protect END_PROTECTED
