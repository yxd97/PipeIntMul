`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ODryG95fpESdwTTzFISTs9s1D0hDnXu0DDHTNicx86ifQnvW7oXFotDY0nMzi9E
1uyrYyLAKPmppIYWYqGaG2tbCCKPHM5O8nDfMGkEjhoDJRflDiFfhHf3/dNQY8tY
piL4Y1Ita+afLzvLJRBzTf7BYX/5iHyQTsz2BjpNy7SYiENCPx62d4FFmnbyDE0l
Hwj+xtFe8D7JR1B3TB3u0aqMZVcbz8Km08iS5fM2hk9r9HSWhD7pwTV0OLUG6xk1
kr/nkqm2ngp+rnMozio5QkfveTUIj0+xaQLrdI9gNVucwwgNYE8FnQzTgVeQ1m6e
xevCOMBoBGpU8JEWhrao1K/nj7EhCg+HqckacZoBR9t6nhX8S0QHF7BVPs56l1th
e3XMlLrbxHmv00+/bpS6sHPK7h5j66EAqka9Znb7ElG0kHjHtQ9qJTVneyRlVQk1
Hz3vgB5djfgnzPivjYKrMnCkfrRX0z7q7TN2eeKliVszxWbRufsbn70FXjig/3p1
8bF8VOBhwV6KPczazs8TKQYnrt/8DGXBLLXVVqLRyGwY+9AuCVhdDsEZAQ903IXr
2KbtXxvZl9bXu4IIoOQ9O4wTBQTrBnKQGXT2TAASNupjw6TPOkmiChcnTWRyVUVr
XVhRaY0U193omFlocKiiKIZWtZKzrjLs8rlCUIgav54UkP1L2Z4n/vBilxrWRpkZ
tFiyVaunsKsxwhtnfdDvIvwslk8fo57LLm6WONHoDsIy1VMBDsbhhK5J7pkG38+k
`protect END_PROTECTED
