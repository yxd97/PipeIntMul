`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yXjcF+Ep5TIA31wq7Nwo95lT2DPaxpN69hvzBTurTCl9D9lr3mTwRqXGNdnI1Zs1
zQutoq8uPSah5V2yC2QXaap7mjsJzn0h7x8DaArPD6y29zzeaI9fQ+ghcxO6GV9r
eRnsL90IEJpZN++iHy16N9yxaVagy5Oe0cV+sSchaTirB4nHte+h+EpZfT/iGqm5
kAB9c3FtfNcwg0SS8Bwv304GL0KvQmCRDVJmpleQhbPRumPteO4uNHaeaSUkeI96
xUJw5hh00jClGBgMJPFNSK4d5nVYAq5O3vPrHRnSoFYD4z9SPZ9u+o+DlTo2DkW3
MXaKwv5F22BXp1SPSbmiwciEQME1OoKp9ZshClr8VFCLCo8vOjNMDflrIcgH9CmA
QRrXpgLCvUFV4PQrkjnxakjmuq9lTz4Y1vuT3BvLG046LKYSS80GkjiI/QIcQ0xW
TLzIzX6IhFis5++9KP2ktD9vQnjY8FqAnhV+AfvWd76dBbXZP9ZQx3HiGtsFU/xW
`protect END_PROTECTED
