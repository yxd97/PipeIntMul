`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOpZCyEDQMpkmLRM/+etDfrNqWTNX1FwcweRf5KDXgoYvWZokn0qKZvAlB6LRq54
SCFV+o7Sa0wSUYKPCRNJe33MuGOt0orj6E531TSm76QERSkXKpdayzOckp34Cwes
DLxbwdjBTYNEcaR6vfxhYl7OCdAO4WVDmRLDNiBpnEChc+iS0AAzxCrM9k4J9r/l
tdIuWZW82bbMCSTvaYmVrh7H+AhqNuUvEJucPGhaXbiwvIG0qgIBjYJdIGrBjIhv
+fqagmmIn0H8pzDNhs0uyatV/2DCxbM1Aj44oFVnHZq5oDGWnjfYqun8vo0c3Q8K
cGBsQ08jpg1oRVEbLh5fLiR8Vmj5vf4fdznBhU+H8RdE4TVseGZhKf0txkQG9OBM
8h0QtlPVpYO1c572yM791V77Tbev50WYor6CcI0yeuEisOZ+2UhdVp5B3I2+WF2m
P2rnwGg3T3kUljOkjGsLRqqTWFSh+K10exJtLMrwERrIBdRy2yRhIJvB/G4we2lE
0iUCXUlqSs/tW0T+SaKsZHaEOsSy4DXSd4B9SnxbxfYOJV4NXXE2Jan7Mahvt9f8
`protect END_PROTECTED
