`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0A/AKIOqwwgQQJ6RNzBiO9Aw6qxG7OwV7giP5SMVSz4sdH4CGJxY3UI7uTQlvxWd
Ntv8DEtuUuQw40fiJqTMGvGFlSqkl5W5tdQUmvG+OmfkK7QC7MsrtrgfMbQtRFsH
S94DIZbt55bTfj6qWYtlqniyNmOw+IQoteGZMvgbwTfthS/vOI2XifSpDXJBTcvY
ooPG50CNqvWVpSE2DoISE/m3TlgSAkU3i5NKuLhnf6EhBysACj8/g7v2pqcd8wAW
hRVwAqbP0J/qgHp5MnIJ/GLf/SRGb2utSJ3ZI8N1xRDPVue/nan7hsj+mWnXjElE
c+sPGbz8PcARv47eZFk0tg==
`protect END_PROTECTED
