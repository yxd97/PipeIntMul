`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3S+Zr7w2/CosOluJx8PkcNF+2sQ36aHxWx1MhPQfED7Va32xrHkis6SG64cFLfXU
gendX2yXxhswdYxqLt6XrHKoxMPwZ4YWvdBWhe7Bi+TBUHSKxLQtAhTwsR9q5vm7
59wH4GicQbA8prIUPcfnwoC1eJ76Dl6LSbs5CKXOHrNfeIn2ZcHGgIsLhMACfzgi
CehE5x3ifOUE3HpUzXqqgNdeVEyQi1FNfCD6wfZoIToNtH9oO8I9VG6nFrIkYyCY
eYrQui0UG/R4kxj8ZEsiyDS+KpIfsZpWWMaTdjFANsmtCIRq2SWRxRMN6qbXh8Gn
T7tOUC5kufu7ODlA6GUnjOjnzTa97kjwsSC33EAPBmA8PS72in06pIvYH9NavKBy
nXzkCkfWIPYO2Rp7jRf+86VJCLD55YyTQhziURgAXFaXmR6BUVwPtKSP+eHO0lDz
z/gJZL0wVK/ekpm2DpKQPw==
`protect END_PROTECTED
