`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KvZC9y8y9E1Atpt4shy1XASdrO6Iv1f4Dl27IHu1/1HXEcpWlxt5DyLVhYTv8tKK
3ENj150AzeFFrmE9HZtmtYzBFuvyrSnHq/ZzNXRqZ74YLXB+brtP0ozK97z1ybAk
IW+X9qP4bxCWyudAVPIGczSNPqWRGR4pdijHTwZ2MOtoYG3vbK0Ua2bRFGHNckeh
c7PmPvlogwbTdoaa6UOaeVJe19ofbjgYM6ueGCm/TMRJbc04hd8t8/oHP4XdxoiD
hNLO3ijhREmt2EkKdCKGzeUEl1UyCCMV0V2VMlwwwyDDC074rITIFAD79zgBBWlD
`protect END_PROTECTED
