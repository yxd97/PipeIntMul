`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLHaJoujvWse9rj8yGYPGPbx2vDEdQYuoFMhkyYu4XFqJan3wrqaEFU+ycN2JrC9
MLUu6X+Co8gcZsZ0zRLMH7aUYB8La6fAdKt8cDX11TAaDWhC5dVQhYy2/DxKsBUV
YjQ+fUZgzBYV5wqz0aAVIIpDaOHMuZfyxqJd+aN6CTksa1Lq0YpC+lB4PLcklyqV
OFC144hXfsE9x+tSJJ5wgJrHi5USl/Wt5eGw9o9vFrXVgDGrkqdj7qVexp8Tzudv
V7mcPu4pYcoLmmrDg1myzmBvsAnnJcrz6xhy19vDz5HYlkfQ8XdpObHsFwyNCS/7
rx/ncjTQv3/+/gekUBYh3BiHfV6cO1wlwUgXYtkrBG/xRuPhDlDRh+A4kCxaFSW0
tPMp/DUaDgchpE8kNzEcXQ==
`protect END_PROTECTED
