`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W0Fy1a5FTq5Gpxd/F6CV9GHXJjcxVpFPcX0bADQPyd9RIGh3D527p+4VGaZwgu+a
jhDSIvzEp+udKo8JqAr2uiHAgMAFi8rdhGjFULYHTh+pnKkqMJfgRj+eygM+5uDq
91J/YwEgI7aGjnk662lOuAQ532sPzw4vNue6QnXOEJoBiyyBQe689EAikHefanut
1ag0Bij+pHqAZ+A38vohG8A3DLdxH1PBkgISFozZx+Km9AtFceSqAHzZIppX10nX
uM1sra2P4L5ZngIXlt210VtpFHmRcFEBwnsewwViAu2Y2qi9GZddAGZrKuqznZG+
umaNdLmNo344lIeD80vA6daRuUkPkka9QASB9jTnk5rwTStdXuYZm/iGftWMwfHW
`protect END_PROTECTED
