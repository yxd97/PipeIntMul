`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dNgGcIhunahp3dSHbAcU+z6W9IPt+Iuntt49PapsDmHL+Hz5plI8OVyrTjO9gc06
aWTbSGvIqL/vSFKhrHwmLTTZ+XK1BHDgY97pkIqDM+N4jRemurvjacg29PbsAwES
9/S4K3uRWksP8d4hlzM9gieF3b/5SS0hFsFFjzJBL9ITcohkx51wx62F9u6D5PPv
yuXj2OhNiJPfGKBLdExqRZLb4nJRFArusQeLRTDVVO9sNToj+N4QV8WR9APZBn5G
E7p9linX6+HXLZL92CyhV4HfyO4Phnff4Sz5wH2cMh5dxNDJy9HRGAvi7r25Pywk
JFTkEaJdCaPnxq6MV67rQTXEmKXE5Ff6iW8Gef7nxxMp9L3idzqL0NOQ8Rji9c1g
jZABdblchbsSneNSfiIHX/j0zd+7YrujmdjFhLjImhhJ8qNNMRbndta78OhaHarR
`protect END_PROTECTED
