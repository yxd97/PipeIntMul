`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AmgVHnJXX+V/v9zG3RInzNyG53s0vayf3Iy/Z7i9xVN0L/1DOLBA6Yrv/2+RnAGX
s+78fnqSQFbAbvvZCY2W3NT7jaQqrYlxoKxhAjZ9BoCIZEIr2FVqNsPS7tOJXONv
+64M1/Oy6uScANjJr08d5OoCZhThZTZMNjzW6cS9zeBfPwaWotKIuen/PV1otGMz
twOEeEdJ34tVJRKBMn2xVUt8rlQToFFYAFyjNrX1s5Dp0oYmJe4H5as/aJXNUDw9
VWcjFKP6ml+PYuARrITfTGsI23xcMyZVb9IRlx5BVlOjc9lH0njHyO6Do0l1Rnen
mrByvJgQFJpnDZ/9jhDnZRG1i6msyr2XZ/891oTi+gA5IJchWAlxAIw1VObHM4He
c+guSJC5UFdBQxcrjqT76g==
`protect END_PROTECTED
