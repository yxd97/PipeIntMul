`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/CcTgKWH22xY6/ehnNbBtK5CjX+efg35M7ZlRfbOuXEn9VFhodAldvir8+KvBos
rjL0ULuWXbYs0+trex0vBp/Hn+JWLeIrZ2JJzUCwAGmE4Q73RYBFPljk+6JqmLuO
8CTxI9shDqudyASO3AIbsp9BcSalfXvUO9ZRURIKoT3IBzPIrcC7cE0myqVRf4Jf
I83nINpDMbX3clyBJZVpifzkjQd9zDiQGjXT3YzZDNhOm39AAmaPcr7dm6HaPHl6
O+8PoSAkEQvIZpZRAqD8kzXzMUrJcrYouQUqIjClJns=
`protect END_PROTECTED
