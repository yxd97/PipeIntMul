`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6By/2ot+yJNBZHDUTuarjHMLcyGibeycIem/UU9foszmU7CJsoZW79gWRsfUGRkC
gpxCTBZg/sZdAnH6NO2m7zZsvw6euDJ/gzHrAQWr9FKmAqZQAV0H5HuUBTarND2A
oEx+hbGgHJPQkveOrn0fBijVWqC/12hOf4mNSW3RkY6QZwcZtex0yuZ+utqWdyRe
cEEttCEJd7GxkciRb+V4fVl4Fn5qIFiy9fZIWjHMiE7mlJAJZkakBxJxfKTnSV4F
pcx+mxwsmIkRPt5gq6k94h070W9Mdp5sklYdi1+VBuqQ5UuZoSGLQ3vDiX4nSgI7
1FVAvdJLtY/F41oFL0I3tw76WnwAyFLh1q0xzJ6MeDnJSNcpFy6daU+mI+l5wez2
JvNW0HT71ijrKYkT3rkdhPU1mY2f0IbDkIM+SQ4sKlrWLIZsuSHUldsdTfkFeBXx
8cqNykFzX/kvIP71sJL7453cExWALqxdtPrxEKEqLxzkiYQ6VuNXvxUpPmYeZpkl
D+A8/qSTOMaxyefhN8U72VpizaNJby8iRj+gc2F7jBhl4Jv56hUzd/81WtFEE3Ti
CGAipQrAN1GebR0aM3OrKcSUH0/PH9Up5IJan/QwHHnY5tRd3YtAOuGldcdsTq29
TVVxBNpwSlXdHBnyovAXhH3Y/pXSstv/df9WZoRTldBQxlJdm0yQtmJvFEHf0br4
icL60kiG3WQWEx8CmPGLJVibEANe7HAiT96IvEs+8a7FQdxccxPVJV3fRORjPl1J
/e9HnPtZmJpF5VvB15UaY8DjRWOTjp4Xve4k2rfAxhTDdmx1uWxjw2m4TtxTIpjD
M48NVPOfLxYNCjLWVe3Tdq4qsxe1tymIwx+GyM7deK97Z6itNeiNtQKbNGupaLTT
ZWmfGPM3O8e/coREN9XgW8h/OUb8yztM7bYyDfk9Djl/ZsUHffzATIUvG51mNYku
oHK49l9Rh8iR5XmyiuEReDkkZybr9QxTf9Ez8AgaxqhncnNvgE4YLMzaxEwyanuf
ftoh9oiEd6BuR3CpD2pVZfYqym+52sT3zhUXOeJdud/OsYDLtmyykw6kWd3ylEWt
TYYb+McKzObkg+2DeplyM5shmr7aXN5dJAOnF1+oP9PIE9hk3cLz+g+e5/JUvvc1
15iSOIs17eXKHs4uM+6vaKzxjbNGkZJOPYjGc9Yf4llylydEPqt/zbW9iuUwtdFl
DfoVesin+kZQ9kvSLQfi+hxmrY9i3kyuKColEUGhHrBZvPcgvwV31xl4Ru3bZASh
jQWzOmsJCdHS9YWQRaJ7zmzFWwyzkMqDOMsMCMMeAbqR5s2hQlF2hNpV8Ep36Crq
IvMGMl6MHae1QDTbrdTJyg==
`protect END_PROTECTED
