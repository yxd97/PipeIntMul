`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i0IzkZQ5Dx7uDpk8p06VpFXR0yLgxE5OSeYFnNz1dJEuY2qIhqyZCfZxpQ5+8Rtp
OH0Zm4EeAc5iGOWJ8pWl7u4TZpkOXwcFwezgm/pfLuSK51tOHJNe2aJEW32prBP6
pv8ZxvBhw2bQsAgtzh7Z/yyQ8YLqbtwIS6+CbAHQ2wfQipa1z1cVvBjqCXxH6W89
zL9eyfF7dcVU5Msiu5t61bTzjie5UL2x8qpmQ0BpWt4Dufx5ek2jihVHcLxWuOoa
IiuZtJpS/5Nj4hhVMWxkGoc3ct5TSeZE8hdShYMZ/uBvhbQoD0IlBvyl6RiEixD9
unl6aU9SKeaS+3OENJ2V+goldoctkGVWsIBFqYLQm6NA/K5f2JDWKbih6nOGczNv
ME3nQn3HGLJHua4G+48WTHRyz5ks2381973br5ZMWwm3M9gbbFLhnV5d89V3qLns
r+Jdc4CFZwNIZXvuBOtM9zwzD8ZF1yqpJZTquNBJ8x65/yWSf34iv4K7nLrJeIlb
N8ICMCrnixOwj346kIe6/UjpjOrm3gEiJ6nSn4M4nkF9FBFfv6cAjTXWw/46qMdM
B3UTP5PrzXdSDjRp++ee9MPQDRu2eROjaS62D4I3B1brupFUHh4r0PZ3cousTkgD
iXLQP31BC1TbnWa9chgKdTaleE1Vat83+Ep9pc3j/L+Ov7tBC1LybkOcAtNDotyc
xKRbsGcWEca0AJXiNcgRTybF42QmSjZy7o0FCDynf/YR9Ojpk/W8McmNRpQXA/ib
Psn76SYqN+Ucfx6jLC5FizU6sVUGxF1mZ9KX1vI/CtPaDzR6G9tk93uyvJR6J2bU
VZHg2nCJh17bvEn2snrYrBlGKFfbPMjsNvj8sJRgzSe2Zdo0/T5/mkfLY3GIGXHo
lfou4kllIw6DnrJFi5qpgQI3q99qZZp1G5MnEERJPpzfQw+O1meUun9UU89z7QCc
KuXprOOOpBLXqmLbPgSkfyCqExJhnYxvtQrOrUe37wbzW3NEvo7Pen7ubGIkMeMC
bufMMDy1SfInsd6RnYV0eFYOZn68eu9f6UEvhoeNNiA=
`protect END_PROTECTED
