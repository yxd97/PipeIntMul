`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CFk1Vvf2VYbi8FamgM1jiYCJ+GHOExauJjeHR8xdfiQQOwlERu2aVgWy27q33jwW
9W8VMMtCBZHiRCpGO0OkW8Ee+dH6a/2dAbrxA2M6JGquSsoyh5MBlNxcZ90BN2TP
tmu1tx1OYR2aDm3I73KM+FRKPWCYDrKzhFDbMEw8v7xzN93eXATSzfhYS9yhf75G
wyYFRxUKS7cTX7lDBr0VLwZEE4G/jUPs5ow4qKkulH/458gxxOPL0ytANL3WVm51
ReB998r3VI4NrZReDo0L69h4xXKj/TQRu5/hTew9TIcqwbmt2Jn/IO1TRrIEDKtN
P1sUcH2fL/dUVs7dY4Oyj6oiKTrG9Bq/N6/ZbyRxf9D7xuKzLfGLtZLId58FAxK7
QNOHwWpLPEvNFiZu+8I7w6i4L+BXR64V4EU9+Mn2cesSL0fO8na1KxqYLOMijLkV
7N9Qv+2YrKXFbBFWTT3ENijboNGLKySIc91cXnbe33qkDi0mxGcnqbKnjLkjBlCa
8y1v0Ul3PuY/f/QmJCogN72wXj5kQDlhXJsF2tG5WjY2mkU6e9ON1rDOv6f+qFea
5JSCSTT0oEWfAz7Z4H12ytz6LfGA/xKpIjgVcoakGBcwpINjusan6Y0UWoQtppTR
qno7h8KEABmCLLagWmk6A6KpLnEsD8ihRouisz/rDeeYjZAAqNpHNIctyit7xss1
9ZUgJ426Yc1gNQ7dxm8MU7vojRunl/5EcuvPTGb8hstcVgRJ5OcZ/IIpIp16eEzI
yc0NVHzCvgxlT+ZOx6oGCX8i0cRclGKCnzrwXxe/az3RABqY2hFkFBMKMgO+u5l6
5aW8lhPYWXGbaZjXWqN9CvD0sahNTCcZoVWZ1sCuwf3aW6RX4JRGGdCwiLWbW1/g
uCjbcXpRWSDwRuivqogjBMbMk/hJ83+uCSt6ECyk1ysROenSEXzCwJBun7/iKd/1
QWV25097yvhZTyaNI6FLNaAbHQIuy4wWYnNfxOxAZV7btyPvR7oVn9ABNEwdrFH6
ux7P84IliaA1NalfbM4spAwWh4pspdgh21tXxqWmWJ512NLQQwuSOlPHc3ZPmVpJ
DxRagIorAGY5k6Zwi7XsN4d9FwI0YhJxH9I0B7cg7drldXnfP9x3Cw48fosGXZ20
TGzXHEa6iSxVfvsKufVyj5/5VOBesKHgJZUaFiiIkrdm4+USbFOog2nwu5/e72jZ
`protect END_PROTECTED
