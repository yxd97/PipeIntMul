`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uxqwPcB0ivH591SWPkOfpEd/5232a8emCB9jfa39EHQjxCWyYg4KaosZ6Uckk8KB
ulHgIvUdXhyf8t8sId9+SevDATw4DSKeF18TuVwnbh3nDHLEJ2BgQ5ax/rmj4Yq1
0jOkeBqeh7ZtabjYRCW9DVxdGQvPaOsnJ+tU0QICoag0J/tne0wg3wpo5WrOoviM
KMgFwSGhzY+M3bOwXyfoEHXJoBMoNNLUIkgzprDyeXL79WWMDu6y68C6OHfRRoqd
j/zSYu8SeWjvd6nEFSXr5c6TyZz8dy3lgbJ4xrTFeOX5VX3dCMXWg/Kson//PQHe
Ev8SM4Za0ge1786M3lkJMj+P8kUrQxkTrCUqu28CET7sj5rcA9qK6Gw8t319OySc
uxp+YaGvbl3FEJHy1SJDTX8LJcYBF8GF+b/1nqqiwHeK28ELFQxTxOJ+M/fJN33T
jw+CMDBTwNSAFT62ugQY+RHI7ZbhMk/dxwypccToXydh0ETeBJKYEuLrm+jdAneU
qbItt4+cJ7+IKn3yMogdSh8IIzc8tmnEScf6CN2mmmGJIi7oapyOlRZJ3pCz+s8m
lfzVPyQ/ntyeTKqNH9d+l8vBLZSJw6quKE991bRBBy1W5OJEFi3/licue8D6XYFP
sf6o2NX8WPMqwEISBPnvZ7Tdiu3KDoQfcWq7wSmZbO34GWhIVTF9iDfZHksRMs3F
Atz0SWzZOh2KulToUpYiWFvfEukh/5IpXzrVFvxfaMswjhiABiHLxI/Hc6v832ke
FraQmVwv919KmpWCjNXd8fb6oPcC9tajPa9le5M9MCw6F7T1gBL18BCI5bTANftM
Sl4OnWkZKLziFOFFZDNySA==
`protect END_PROTECTED
