`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jcAPJm8vcVsTsASnyRW5aH9SHUWmEAXRJ/tDQAatN1VZh74a9U44kyGxxYRLp6/a
CqpnFtaR4UylsNw9S21oi6dn+ynrktsbMvnL358PDPO11kq/hhC9DsBHwraapzcu
svYDioAPgMfS9PMuwtwJs7DNKMED7sucroCx4laXiGw+UV3j5az0lpPyzvmerrla
RzPfo5XirhAmtzuXQkMqC0Dm+i1foSJB4nfACp+gdkbeaXglZdrs527Xg2vFLbTG
rM5bcEb72OhCETt3xdONfwTRpmG94EfMIQtZYJ2FcmNNqclTgmsu1ZH52F24+/+N
k3WBU8vQlntj8QFBMKP7dA+YX370tlijYV1I21Ank9GAGDWE5LmlnEz7VUS3aHwQ
ByAOVc+MW7DRC3hn1VaYxfYZ2lXuUNoCYjQIkM37A6krKrsyXfvEhANf0ebCme6L
UHRbbsp9G33pBwxuBaAgz+i0X2preZBrwRJUT/G7mqD8mH9jz/mCfMN4BjQWWVQx
oTeYT/LSGOcoXEeDtE/w9FstMKut5YIVkgx5Jml94J6NlEOofJOscGqo/4ZMkDGK
n7JaZS7d97t9YOjySN55tgf6Ok8IGgxwLi7m8+GBIQpdRuXNpbohcP9HsGt7Mgf2
BW9gO9hEQgj0zeMiNxEOnEyAQBIOZTouDuEWq6TNaksK0FGrZkNZT+cbVjLc7nEm
j6anwyLd1zzacf2SxRh8Hw==
`protect END_PROTECTED
