`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rDT1b9MeZ29zGiakYFDEEpl7WmkwLSNh7GhqGYG5Eurjb7cKIKm0Stsq6pWa8Jtm
oqDo6YoBynYf5G2oGYqSBr9e3JAdi2/nbCKXzN8jyVOu1iJPUkotL+um+BlOlLEo
BC4ZY2/7l0B/BKbfzYhWV7aqEqBEQJHqzQUAmQTC3IVKXUjhha0LBlOB2Nfi40Af
k696YTcbN2IUqh0nY8p2cmsKif5s32nAwf1UAxICsRfuBqmEcZz5Xt4eY806N83p
AheQ09CHmdNI4GSoFAHrCen2v7DgykgDvdbe1hsT18ZHFrWnyBqYZSwmT7UeoGIM
0bYXMw4OC2m5oykCMyRerA==
`protect END_PROTECTED
