`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VqBzRc3YdOrz2nl9WluLffzh2QO2Pk7sqaQ1KkQCDZTR3Ospphpz2oGx5AbrNf6I
OGbeajLrmb0c0GeL73E5L6Z3EkfajyN+7SN1UgU/p6P0umrK/59xhx3hA1PrqreL
juYqdRxilosFHyy+3uue87u9wtLUa0rUJWA5F56IL0ZCN95XLTbB7A5T6ZgtyXhh
8V+myy0zoZKca3vY8l67/aHWru0OsX48j9q7GHiiRWfJMxAmL9FdTdcIwUObbFMF
XTSzCvAaZKwOASbXWbWjyLzvmozKeO+RjV+3veyoBLwBFEgEz0hQ2VNWwZn3xzXj
Lxqw8kwETN8KLhX6kpp+PEFGVU7uJGs1wMuUvPlwYlbBkULFIbqx9wlMNjl35blc
sU/8jGRxCJkLkSIM9vYARPWHa2H6t/TEhQOAKh83KY4I4ejY5JKblDuBXbOhBkBb
HWt1jEvk3mA0+fb9K2rOWGeVDsEXwA7eo+oz2q0hXvVcke/Pn3ZPvs4ibeVpDD4/
uYUTTStKF25v0PYAWJdZ4/q1pvgak+h7pvB7lDLfrOAHbFYQ6atvXz/c7otXRATf
iuKcLX2eXu3xkANzZrTe76Ox6pdQI9xY7KBsniVLLn2EGuqrKiujZ2/Hp4Si5p1q
`protect END_PROTECTED
