`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iNJG5tWZvFLjDpVAiMre3mnYb2rQBlPEwVVxt3mKsLQkK12dFzgG/3kLii+gv5Sc
/DF3MbpDMs2KtP9mnDV44wxWghyts9pkWtyNU6Cn3UbfjNho47TPUjsCy6fKqFoV
sVaxJPvLHqhOVHopsJGcFj9NvozbdUIw471lwwTXwkvrNijv6kpSp5XjtJg8Rj8R
B4iShCmbSlC3i+J3Y5hOrUR6FFZj8+eqm7tZaoUtbBhMnBsOdI/wu4tpUKYXDV3J
OKit+F3efNmdnsCgE7SbQRgfSJLfzSvZAXDGyBuFooV2qZHPM5ztF/yhH8isTnjh
J1TnswONXIsREmZj2eM9f3kM/5ZQBtuubKw1ARb2Z38hvbuW4ThJsgwOjIN6adq2
`protect END_PROTECTED
