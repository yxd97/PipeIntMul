`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L91REqfKUJ5C8riZcDMnMFXZugyGE0eWQOquyED+PVKWP1eBoC0t/5O1Ysw+9K7O
NwAg8YK/aluBSxv5CTrhN2blQIiCh9AjBEVWJcnzg8k/pt8A5l30hr7RRsXMB8Id
55MZBz5Uhe3DCOrphAntNUTOkpFEWSZl/aNm/wA3PKHUkhIyPRqQJQM+QP6kf5sy
NCxC6xJFC+I5eJw2NEFqFe5x/9gY241RBY3q/eZ/A7ggzB9wKzdqk8fCIv2t+Oz9
MQuGe+IUBY9Oa9gFBlRolEK2TjTy1uKlqcGZ5KVSd32qai1gnjyjApSJeLOVrUb3
IdKVZuqTKLiy46wxb000EEsyimd50nsTf0DTRCw+nzX47MXVMYc5wmmBui2YdMbK
aUyFW2oBirjdK34jn6KXzykoVtdjsomvwN3kt8dzhzpm1Eq16M8SJ4PicX2Z2GBE
+zO2MD2Faag3U2Wj7HYT9vYQWOydmIapZBpMV8MliABYH1iU+id/bq2/tlVbo8h7
Bx/Qtdb2iX1nmQpkhm+JbAJ9b1LDSpdJsvJe29mNXRbvzPREBgYdf0LtJZI8JD6h
14IKHh3E+ZB1I5cufL+KqwoyIX0K/MiO9GP0ImtMPBbsXBsRiYlmzPyZ+6CUPxjb
i5qQFN0M7hoAbIFJYMHw5nNUwtKJBRYTx4NlvpQRTf6IYliTIIFaTEB3WEDwFxze
M/0l5eZUZ3TTfYoqGCRPPfrZmAMcjs/mnf7SzP+v3D7gVFp173AwEShIpi3fk5oq
PMGYNANbJkGAtnxMBRtlfGbgFP4AReocqCpyHf3Kc5PRF5geJ4BEAwvi+xwO7U5o
PKBQY2awkFYImKO4hnXJjjCJJ7lTxg4vzOsu6BPblOTVEpVGY2vyxe3V08tTD3YI
V/ue282QS2K0vG4UvUpouwfRiMfwMz4/nWnKxjqPiARoZSVDPhcqB2m0LfftnAQ+
`protect END_PROTECTED
