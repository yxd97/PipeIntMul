`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DdTPxqqu8Hy219It8Jb6tQ+ETu66cIgRFhkEH828ckwpxINkUf/Lbmt9Mk9Gutku
V956tNvGY2gM1PbJmj4uVqsTqdPrZGUlWC+gK94wYo4dHKzltUThojy5D3XUQX4z
FIe764Z5r8G3g/FyLAUkfJz9/cB9JW8VNPCvW18/N+qvxGJZrf4HsthZN4Q7vEG2
yjAJQxTWIxgBOjvPJcPbRz/LebY3MWMLTq5AYEjURNDC4vOgQm1ewCw7htMIGUNi
YFGF163fLX07qk3eX+O8hKJNPc9BJWUWcC0dFNx6VFM=
`protect END_PROTECTED
