`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fIeku7DEN1rgIER+o7owt9Kra5Kup8Hg2tCcC+ndfT9XieVlBPl5jeG5cfEpsmk8
bVQh+ebxIX9e2tw4W9NlX5ps1jFOQXBTt6OX8MkacD1G7ZrbtWJ6hcfTt9JQahAs
o9vf0a10e6M2jTqsWwlWgIA5hylOjA52q4HLsR2VcH83GZfIHKDd+pNaUUV1e7v6
f1cxjIfxVaVOaVJYaroLrbMAjYdFW2MK+HJjCc+BZa1kfVzej4uEBEWWdlR8BMKx
PBQsxAjzsKoZ0ifuieHCpKRpcG+5eOM03M99bkp/xtANNZ+RsSG1VgEGNBic0mmA
1oUOLqe2/P7lhufshwFX/tAkTOOwVLPcaQ3l+ty9blI12BHU/mZPH6UMCTzs/qmS
JJFMAwu+Dm7+DJdGX2QeFA==
`protect END_PROTECTED
