`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qno/25/obRGfHdw6BHqRj0+dMXEu26hATh3L+kJC6qw0WSctkGGF5L/JWVcE82bo
OQjvsAZfa5hqOhzxsEju2P63nc0tk6HvEmuk4ZmnXVSutsnPObkDRlqN7fJxSMGI
8NQDiEtG9BA7+dgPI+aiDTWWmjY3o8sTB4U8cyIf8LQOHbO7tsbDRzpB5eNoDvUW
jBKz9318gvG0FvW344YykKEZls3gyPop6JfNcuSyEl9aZIi2gydTtj3Lx4j9UKk/
pfaRJMuwc40lNemH2g+EXt5fPam9oDsVqTtdXW05kjtf+T8vZufRjApnQe/nONuv
F7qHjnWF23BmAlClbvNLNNypJAmFb5Rc2X0JiMWatXXPiQjcUzUPYFMnBpHEwqvl
B2Me8hkmw8r05xmsj4rX4/pZjm01h7WF5Xpwy/3pWRW9uhlFVRqmSlxWSAw0B2s+
+HA3TpLLplileRijoiytP0bAT+RCYCSY/gzQQ4CggnfUwytmQV20CtxMN5cQWkmX
Kk316GBU+Cyuebz8Qp3vOhQ/rhaUBYirq4COJWUmcjD1/QiSQbtgd05/ioiTE/cc
2xwST4qrye65ctnMOhILOU55a9DijQ37vzMYIrblCHy0wrTT/UK+gxT/aNW3DOzD
s7QNXYHrskeoNdW7+WSUpuADaGgaj+m+KoJsVw4yz9HSLYeafZNIRelC8SEuTOu9
U/k5lbRtjDpS7lkYXquK29w5WXrCdAb7bDraX8/JuVX+P74SaU65qpuY5i54ClQw
OiKQFwcOO1uCfJU34wS1Fe446Cqm+1WhEWIV8j84bjOmodNH8YULO6ZyT/dr03Lr
UF9mLKOajYBGdrShwwTiJXsp3syx/rlcLEz5hCFahj1nLsmW3GfTfSzUGOUYOd1f
qoJsBfTNmTO/yeQfo5mNSKfTsHop9KJgKLdcBeVBDPr299fUiRfmmxsu5IWqrkxJ
vyEkjw35bQfl3lEO3UzT33mbqCDl1XeD/gz9VPH66zNZIR5yDiDY7B8dErSwKijX
R6BZh8n6p07n/5ZWr6t8BXOjmJD67K4dYKLxeGv4AEG7FzcTGvfFTN+xX0NWbpmT
vKgf1K/SRYNYNWvnq7a7UG21eQ0oHyZPxzx8xCV9vyfcKbTL8VpLHnxEgjmsKULx
G7vZ6+uEIQpVIRMy3BNuNlvpwCpsbohgYKvKFOlXLJ5l+i6QjboH+NcVOWE7ghBX
4fasnFddPFspDDPVdvwRk/YjC+NnJLOpa2ans9nYix2zJx29m6YMGMLLK82qU0dC
v5UFwm0b0MV2xeEpkQKNkWYchNKkXI6Ecveltwuijf7PUXKRDnuIQE7mcPvkrwbE
WSAFlz9tjAis/xKHfhYs0MDSO+PBNgdel3OnHcoHgAp0egwOR2fiT9qtxebcLOss
CRoIPp3yR0iQcTVAhhFW3KHwOSE7fnjebdM2uZOs1AWgjKrzI/8JZD54rvmBdgEU
ocShe14yYOAqw2L8I8JxYWnvWy1hyAl6Jseh8+qOwsRLTIm44raIiq6Rtqk+Ctbo
R5zCXmazRK43RlD2W9C1qzxbYOAfNG7XMha0rIIaIqdxpYXDMF7CV7RjG3AYEuFK
TptNVSRsGy/YPbC/UhAZXIcRBx8nUOL1EGZAKDdJBQEpbg4Fe8o9spKVwQY5Ebb/
VR+uYmEdD/awBszP29NpX9S4xqbCQgddoW/rZ5rA1Bnu1pnLFZ9V2VIIr0BTr2v0
xQlDx0Il2vcoLq4eNodbF9GM3EAEyZ5NXAM45ciCiu+XWMmKXsHVmvWZLFfsP2Yo
/NMQxwALMoa68SkVnue3yh6DzyJ4+BjtO5DCg+m7aDR3x9M4zqMp4V0U1xzxUR2O
Y9TFbW8ErI2Lq1kVi86BUw==
`protect END_PROTECTED
