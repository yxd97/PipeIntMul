`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gr6qQd+8BvUCmepzvZJ0oNLI/l+1sr+5t6/ZkMe6xGBmSiuAzkks4TiOpcfDsqjP
F+CPJc4fCrVXGy6uTJFF9N5JkMu2mxvIG2wuds3AH+tugNzILnzc2ymuO0or5wS3
GLutp01UhKV1axehN+rVKn3cClJlRF0s2MOFhpcoO9l3VQAiK0fzWON36ClHhT3I
tjlvEQPk4W+keHc4QoavNBKzCpWJDCQ3BX46wzrW8v6X2dTq/jES5/hSmXMulw14
XrNlACkqTGfI/10damKu8H75kJFYwrbR54bRwIiJE+TAWXJG46AtGb2myXvWDrfg
Y/3iKzUlBMSDRAOahndvT6T18RC8fzUEXX/ytU24n3Sk3tu4SzMcqmkDMHcOUayN
D5HTdgsBSc7vpuuEbcQPfz0VU801PuVFepsbpSdo8f8fnd+aU5gR3zEEtOJNcKsi
QD7jf2GR7eT/KaYVD81y7KzZzzyMaJNeF2cuK/AjWkkyv6xUpHX19hyECHJ0YjYk
Okzw5YWAH170gvvz71IfZWlZpHsARyVFWLBf1Vj+30oVM+Kg8/4ogR5sXBxjNLJ1
LNcuVhSBiyIsR/qz3l+N7Ao2GXSh2Nn3U93U+uREEuApPh/1ikvcpNuCbNIngN4Z
0ZMMxEuCbGVfc3yZm5JdD80IHNucZs1CvKV1o3RfvEbIzT+Olqx0gWvuz44iI2BF
DASCYtk4o8ioiN/quujg7zDwZ1TVqRAXxZOgSVslsxAtYNsj2RcFBPs+gTV6G9jN
eBbBmbldxYqQYf628RdxUa3wDu+/Iye/weJyUtu5/WtpimeQYqHVQXobF+UiK3sr
PMTSQKz/r07epJg4BGeT/FXOFNTo4cAjYWwB6NKOgaD9GW3mdjXpx9c+rtMQ/MTu
/MINKqrMUw+ex2atDU1AcjAuPLTaQh4hNBNjurNFc6sWSo8T9sdBT8G8lZQD2YM+
55J88J7OSm39T9JrjAtWITslguKRX1ldZs2Ibvr5rHcY3r0AOuG5LKDjBH6DEO/Z
wqnouyv7jxMbPrVS0dAR81VB5+KJnCF8Hd6Tdl8SQe6acL4CucjiY00br1WEetwF
8dZp97HXybdJzY8hT8mYKcs7OrEy/zz0HMcMu7mvcpP3eY8tXl1jZI28jP1FKdnN
nIKXhI/GcLDNEQaCIw4r1l2W7Tbu6cR4MlJzhRgQHDJwHVeVVGMAuIGsTfLoRJGU
AhWPeQo85kTssNKRST7BjBQUAxdjTuJTe1gqVNHU8KtsGffXQavcSlxDxHDTjttF
hz4Uj9B7wc1irR3zDHkKnWcREaEo0tMih+UFbabREnnM2l1xi82ZptORU3jsn5Fy
rPu42m+II4MkD8/Qfvf2pNy6bOBtawE7ojJLKSwPSHlYmiH3SVRvO7AL/IJN5Mrl
ieZgZmXAHZx+oV3IeiEGijzluySEoAl+3BF++2cA14iCsCBc57DpvD+XsQgyhjmK
rfafHo+wKu+901zcObwR32ClDA5B/wziLyDhUYaDH53k/4mGP7hNdY3Sp4SdoyLE
8QK5rqa5GWBdZw7Yk6qvlQENeJXDmSHWxNQ0RbwtA0LqYXP6vWeQmkuCefzeDWmv
VcF67pn6FOh+IAT2z4JF7b7zrtvI62+wIOiNuIzs3WPEljKZpTo0TqHPJsWEMASA
2+n3Y0j/RfY7LbZt6wE6EFEYyMCujQNYGonb7uN8YQ396ysUsNgKZ3z5e1QAjNsn
/2oYsugES5GTVcTyrVE6SELGYoBC+WbD7HyL8IrWMY9VOaKLTaKrNzdkQMLuzT0u
CEe5gLL+BjZVrxJsY0mtJFpOi0lvWmLY50q4wb9H7rblD444I/Tw8l7170BeaNN5
cTWRIyo40q7r/F+1xk2a3iPnUHcf4w884zDAVaCZ8JAPdeIDk6c66GzNPPIpTn/3
OUQawtj7F3hHdf8bCnTfUQ==
`protect END_PROTECTED
