`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VT8pIYYeMvhd43hWPQBviUZcN8sN5UTo7ld9iqmm6lCYnGDgIp4H46wZTEDGSSbC
fn7sLmOkuS2Emss/u6v5aGe1RlqO54ylh4u31QUWuAh43cmlmXU4TUtije9k2L3m
4SCJ2Y+QXnCFmRO7N4gj9g7dtB1xl/Ons/KGMlFTEpYeENtAJJaMSXueLn5Fp/ws
u48pdfgqMTZO3sG63E/bw+BDtd4PCmR0BZ7p8QGUMUtl/VFPDTkH+UfHNcLoyFOw
FrXCAHatMnr8326Nf/bPQMhp0rTOTSKub9rWumZ0AWwY+T4pdhaxCifX3wcQwFd1
YsJ56/onHLqs6PZRG3Xh7j5y9DkMcPsvi713k9Vk89ieYQJcfCTFC7ChR3FDeKw6
xwkEMCnl8ZMKeQa3jUGrqLeNsqmj/yvImqAgjxbJ9lBV8agm0rBsNU7TxydOHIZR
3jpitUcv2fHYVOaHUBPtM0CYLtmNU+UWUre1uA+yLswkLzR+8NNXC0kxGeiWhpZC
A6AjarmXWsH13qmk8dX8AHoYlk5dlj0y9IiDdzd147o9OPeW6hWxSHus8emF0any
A1qEtRBKH6WLFYwxclqwYj+wajDYTr2EZrE3p+WIKEt9Dw6eg6fe2AetzaTkY4p8
LUs9T0DX2Gln47DF1cgUDG/iuWdDrX7eF1S78dUeNzxuXPCymiRqwHy+e2WIc68O
/1P/hPmS9FP9O1O5rks5jHuo5TrOte3RLnK45TakxqlC87Wrq+RibecvqKy0bOiK
4FfZJgoQ1MishL2KzeiVjlpSVa/sfBxgN72/94rufkF581qmCrUHyyk/uF3t6eFT
QqT/CUT/QDCNpGmqXRlexZOHeWnnqhNzrxxxmXrbxi8=
`protect END_PROTECTED
