`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogdn1pJIO9uFy1EXgGB2kXGAJMl8V7GvOFG7v749aT5m5tb9eCzWbfk6P05O0a6z
jGqZsI3oIOF2gUpepyadbjaKTP1dECYm26y9UT425y9bMbwv4qSAYSNGLPQltap9
Li5eIR2jp+M3c0m7fNUrd3ya03UlBOxmh5oSLSF4hKN+l6f+/d7fwzUBhjWtMUKe
3vW/dSyKpg9yQN9JtY8erKlszL25Yt+XBqJyc5sjpDcThLqXAL6JCoJ5XYKjSRNS
5h1jQuVe+UVC4uMwCd6ja+MIZBTSxt+SIb2+OJ4Zbguh2CnvTA3PEVOda/Ipma+1
/ZY1TRqGj/MrC3nP0LedGmXId+h01zjzkSSFMMCZAQcousyJpfZvy1nXbzCEXT03
XdO2Z8ypTaPYwCjEmtT+TAv0QVFM6wbaj9rYZDDdTD3sECdVwUO5d6rsZ1US1M5S
jcPBEnAxRmzu09/T8CzgpOXiKAWNCQfJML1Cmubbvy8=
`protect END_PROTECTED
