`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZU8umOgZTC178vjBSF2FUswrPN84y6uIJjUZT0bxWJhssUnU2mNLhceQTbDs5VQD
M0Gi9s5M9SNkmjcrxPcLZ/3aWv0L4H16RyVabHlyW1RSmEi5BnhtR1jOsKGkv4o3
okR/j1MQ0GBvQgq5zFQ4qYg+mnT329gm8b+VGB+9FhIiv5rC59twzm1tE3lUfGMz
kpgBjVlmwl+3s/Ub6mCSiIylKPGbdevFaBaKEje5sqMxuyW+L/Vux6GLQ+WDIV0Z
KopwqHeCLDoNCkPqfP4cemUYtlp1XdzeQlyqBAL1Kp8z46mim3gdhp35cGyi9qCY
+An4Vy39y8kAJPaI6eanGUqzXzSng7DI7hQuACYSN3WfDC5C7wnU6xaoHusJk7TA
QrrZfdb20NtAMdUJ6y2BMLqVNj2sEElrUxAcr+W7QZq888iOh8GU6HSkvtgF8in8
3U7VHkebOtsZHzQ9jABACIMnMwauZZeuUz4vJPe7leY4QNMr/TNSMNSHD+YqVq3V
u44Gx9FA+LGYsH9KnogPhP/fR1fecA2VjiKwlONDT53qNkNuMckK1/fvVzQWaVNJ
Gr0ZBGM6QNeXydF9tWfxh97NRXxq0fCdySQb1PPYyXG7C1IsxmY4qgxlnwrz2xlz
2i4NiMjtfbfIvH5boFQbBUN56ZTpH/sj/hlX58GSAeOUfDNxUnkM+NhvLMbaYxGR
TSs6P7F2ujZupE7BOsyLcCelZICa5QyXMozYrEfpCHohlCSv8mO+oIiUWRau7cXd
vLNaKLUd15r8ezgyXDGYWAVYycUZnuy997AKwUTpE1e2ZaqpTqiywJvHfCRULcmT
vkD7VdnAaxlYkTl1RRsl7E28FqS5YKfnxDGFQnVzW1II0chhn8Ek1ECEwQpYAWBy
4ZdxUBfga8MNtik3LWaUAV1kzeFW7xtL0tzs7YW2w3ff6aDoZEg4WcnACtowK9LQ
`protect END_PROTECTED
