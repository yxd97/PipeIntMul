`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OGhOPE1nXguxTW+LPCmmFr5qMWH97RowiULpcFF5XYa6yS3jhsWhi9sdgbdQjKRQ
8MinkMRiGebuLB8omGojUh4aR0j8roz9lMO2DCRjH+ugQkqPgKLWM0/j4qe4UNVU
4XUJ7lFdBg0ttedn929LDGro07Rm0+kWlRU5WozvlWz7qhslz+IqjK5Vuj5kbCn9
prJQZ7SKXKZCAq4eo5mxC6GZy+3TzEjpiM/f/3uwEkMtOu84ZLcmdvxyovvwISPQ
RKmiULh4tMq7uDheHxf6zVkm18wWaybNKZDQcjY+A6o97pkCOFJ3qLlMiVa8dNIW
QikLuOChs+1CUHB9OHOB+eKnldI2SFtdmJ1lIn30l+fqYcS36/PTxju8Nd9b0Jyd
+0qsNZrjd2GE69zJUxCjHuc/jHL3R07CcPUyqm+Q44Fh0CEPtF75Ou8JMElOjUCF
/s10WB0FELulb0/HF78L+yMyAHsqQyjMJeyBeH1kLhG1EYYfnZcfcdeg2eCUgRxd
BXfu2hwHsp+S5GbVpab36/Rgujvt8fr0CoyDzqkB0fhmZpblRBGfmYTsiuT2Qau5
ZnFP7Ks7ZaD/O9Qif/efQa4h92IjWjjofF9kKlDPOOVpf+4KhsB+LOBMhj2A/vrW
k58P8KJkdxCs6e3oILatxN6ID0awEHIyicjqOre0bacERjVuiaVye2MJk5QR8XA9
rnF+9EHYrn4HM0m5zjrnihnbDmNFDD+kCbIoBd9Nq9f+GY1gMMsgg6O31J6wdjdW
BLatogGMU1WOW/u75vXnWDG7E26Kb52Pbmn+Yj8+TQ+2gxdILbXfvbt1McI/CECu
rr5n0mPGaUFh0PsC9jj3HySGaNVI7EZ8T0HHi8rthMi9SIm3GU1uXqhSmqqENL10
jDnAB+QPAmSDM1d6h5VuKir8Iy2Mo21Cod0p8hw2rw8sQytK1GsNvYrDOCIGYaKo
vuqSIumv7lHleneBARdziN9xVt7RRsNjbOnB8IwQAFk9Py4cSyXVaLeYw0C7Ajin
us38JVpdK0LAKZjoZavGYJj86MwxvEGTq7e/1UOomOau1Pj0Im/93wOqTKEuoi+y
SPtfC3VgOn9eUEv5/VlLeFL5tjpLEgr8nkT3k+Pe88UOdCpc4PFEdknhCYxWMmhg
XFz9pU5K6KWty8zVMs+d83VHzEV/v3MHTCWxZfPgwPDL/8LNp93Of7kRPlhF+SED
xGMFw3jgA/8mNqB9E6it5CZiJTWyxj+mJjdxAj58iz2RSvujrIDJJd7F+mKkaihk
IKaBDWhNbEPSwhLs1XfJM2omekys81e3GXwob1hPCt5JfVmx0sjHPV2cvOq+0V5H
dZkUgAvlIOuh9ZlREFKWJGxj00dlwenSnN5+FOpFQvLy94Mpi/iBIE3lSQ/lmo4n
9deAMCh6JadQvBLTk6degPPX+SdztFWKgJOtLOaQAHTHH/yAdHoZ4P0FAyucNYKD
iuzaw624epgQcOpJ3kiqOZyhPsLavwepfTmGdQ069bUx9mmtufP6bowmqbMTkiKh
tovjbMe97G1U6N0fDU1SLDDzaBTHIpPDQNfzYGIVhZeVdpjuzhkMuR5Qpo1Uv2g4
VremfYCq5rL+3wtHJ1AzSLtBpgPT9hyCTOsSlWhsNXN2GNILpOq1nPzp3L2v/cWs
l02rWDyldL/pDsiCYFE9XawkmwJE6zhrIEvsVNZex+CKDXTRWkpZxg+vvAGbhkiD
cvO3zDc0WJSuPDH4e86Ya2fimCn+P80i1wLcxhUiEb3YksW6JZ7DEPOTcclYXtmr
YVIg5wRA+XdotNVA2L1MJQwZFPM6YYfJfrr2ZvMA1zm/6Sa8AwpLPjtahxRfSGA7
ssASLsZIYbQDTHQ9hfUwPA==
`protect END_PROTECTED
