`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POJe4V2VCBGS7bBv1EnD8UDn8ulWNyltEYxUSg6F3gCFKiywndl0Gbsw/YCTxbF3
sMkRUb8Cwy28KtqZJk6Nb23KTMICHq3L82LalBtsz2mFBNVv4yXAjWRJx4Q5klfM
x48inbdazKmfSWjizvU+6nZmGsun1HfscuXMG+hju26PfRMAEubrZ8zt3rAl3as+
LxicHsDdh8+s7nZQw71s0/SGdIZfJydyEPFXmUqcIBvvYK/oTxPCbWMoGXOPpUog
VVkLHnzEvbA4KzjZS1aqGxAfKKm4DzQKbMQsDnCjNYRZXW9e7YlJcmE8H0jp1U4E
Nxzy8bejpyjJD4jaIBPFJ7BYIzQm1mX8i2R9SXToJWSE2aol37um8ifDCNbXKf/3
OT0PKG7tebk+DoPZcZdqUcOSHQhiXzptcaaVcqlt7YbQQwbOeFoEeotx0RfqF2di
cvE4+B3f57hkO22IGY7/dLwVRwfDzuIkNmpL47uSxdGr1nxZArssQ1/SDMZ6MHjj
0Jw4GCDSNgIR65DazB2CkwAGzwHMc0xSqNsK72rR8S51aZ5KWOUuetSE0WEul4ZV
icuz++EHMex5E29w74c8L4LdJVHVPfj7MP11F40yaKDghs8zQnjJKhoaS5u+dizv
AgCShBfqy22XP60UdcwXs7SVR6XBL3snerdtdB3qK+60lVJQ/B/yUOMiU/K+bdIb
q5HM8rOFZp6DwtfMa4gcoI8OswZdNcZnFXMCB2brorwYUpHq4iW01KNbAq/aECuV
CTYRU4+ErURzdTSOhkj8t+GSTE98LKkDJ18pHFwwCtCPsxVSEwxz/PqwyVbP1LzH
RLH5L3XwpDLBkI0TlDCzFlT3hQUiwyAgvyOd9y3e+X2moXRXDZt8l7zSRuLeSbsH
fIXiy8mx+488dV4g5L2QukAB/RRtQozdhbfucrw8E+vEurzUeK1O3g2l6e7Ij+mP
PQOTgOVrK7AQhGowIhtdXL2N2je2P1omAUgb7DdPgnrHOhWmqcaaYJq5hBIcgL9p
rQU/hlC0Wr+/aDTvZAkwoHggacEKjtk9nsdVYelVP1GP8VfL8vXfQ05ijASwDZcF
+GxuiIZt8xQJUP4sMEv2UN/YAbkS+IcxlNYckPzvN63wbrcLb4gdUwXr+kFS5KzG
HnDJhLvJ+SiNX2UxYPgcoC1pTK0hxfTlkRWHUVt2XThU6jq2OyQnIRd0AOcUBodC
krfn1tFuRw4xg4hcx6Fqe6zwdZ+iuE/mtmbxo9Q/An9/35AJ8wGftLlPp0fvscXt
f+xTVFZbxLt8E7KZeHn2u7CIa+SHtFWQo7mqNwGenWJvToPVKPmMD/PeRfR9bPfk
6Ex+/8zc4vVIkjNPq7wbOltYcgu0buU72+T7fsQ7xLGUDhy+PEj9QuTrpv5VVacY
vtnvVgLD/rzkkT1U+qA78zsAVPmSpeZsWvXs3g7gVPevIvYBvzRdhPrzqADNsn0s
4yrNvsO6jWxIP4MVjvctEOktv2UqhiFHTHjkjao9dXmfAXpWiMoA/D58G4ugF3VV
Ygq9iOVD6iR/eI+cO5En9xJJpMmVbmf0lVqXg+Lw3XfzmzcJ5YrttR5rzQ8BUq0g
H/EF0JG41hIaxks3JXZgjfE0i36+MC4mCOAtpE/LCbpklaSKmnM8PjtSUzywsGLg
vBlG3Nu+iO/wHN/N4pAALuxfQ6AiekQRQJ+beMQByMhX9yXuzz7eI0wSFWVJkBeb
kXUuYUyhbe0dBgQ/40y4NSY4LFyqXXn0bAZ7uUaR7LYDHoOshKV3vExihFDk7CkV
xUKC7n/KnxIZWwO6ye8Wj7r/BoQqDh12/J7v/b2bbjIBMGcbCkBG165sD72AZXg2
U48K8JVRzMPZgxYXb1srAdTPIVvzDkGq5qQEMf0ed1GLFPry7chG4SzNEQEalyvK
b7lFCaMXfpWVboanUWk1GSupQYDE9oCN6bLsvsewEIQg9p1XoiTCM8sXFzumjjmE
kYF6L7NsNg6+oIuWAohSdrPchwXoUBiwN5OVTi2XqVoCFISpGtRKpCBQpBc/6X52
4DgB9GJvHGM3JhtiVYYeLOtjUYLYd2gnfAKn8eJutW3bTzcGt8/1GEJCgZGGAXZP
d7Syr0GY2eZFZzADtFm/89pZujuQQamOLgVWccxypgYjjSznxf8LkbGBtDlFhEYj
JjR6Tlip+mj7/fihq6qoKz1WNJBE3BiDNsXAmOucG9/D3jXdFTifQshm06+A/YMs
0viJaZ6JPHvb989RnfB9scc0VGYpUi+7lh4U9/uv+uvlbON6xZkVEnORka1sYXKt
sM4RrdPxKeS4hWF4y4IiGQRFSHd641JzXpAEM++9YBCd5bSOOXIhAGdnTZzqPhvd
Kq8Z1jO9bVfFOktCGrENTFlmM9zmPx25dZSq+ReY9G+UrQaAcPgYU05xXOmCnKn5
GTVOwjHovMFGpMRo4mqSyG4wPLtUFhPCxiwsMTlbTKKszQsozCSapqTesu+98L75
jdGZy1TBQP85B3yJuKkWyTtlkmH+Sv6PKvcrxVH2HNX3WE1xfbSAnYvN3hkGP5nr
5nlZnQmHAGS/v6oqViw35HktT0HmJMzLo3hbsFi0/JHSyTD+1/Qj8shpMRpUZi43
75+ipIkrW2h2E/5zj7V2HTsUjgaA4CpF6BMUYILrNu8OnMsnOTqAytOEACP9Tetd
LKWR9kWi/1D00HDMGX0NJWxdgQ36V3abfd7FRgnpPs2orzGTPytY+EFJ+J/zEKHH
tlsCBPIUX2rWRfubwPNGG3A/Z4tFWvkV3DlUUQMXiDrlhiXoagefqQcIrfEjdvSV
`protect END_PROTECTED
