`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGBCLSKZu6E5JkjVs/l/ZCYhKQIBfFOqNz4To3yMcRx6o7qd5OxWTzaFiqq/o7fz
5A9TJg54AIGZQnwfrqnRYtCsQs++Qr8gLfMpi6FR3daq9ODw/8rcufq9a2dqYSK1
KD8oaqy66WRnFuyy/p6o6/LQ4+S6pVdiwv07zAVuIG1oqJtvcWQrvW/ztpOfFlZB
z++dy9tJwiyrHNb5E3TwrA3ISow3wRCIhWZ/usfTOWzIMbFTm5ettbQVaNuNMYhG
sNHmqIQqYhi5RLqUXBsb7nGer5VDW4AoNDsJSOy8BZ4IspMZbEylbXegeWMsUbUp
BfuF0i4YXMGMulvKfytsLGiDDFMWyWMz8B2r5Y+db4E6nexyMQNXiRd4867Wrdvr
OoHrrsfpeRHNDXKH2AEfGWngsnIhMZ/HLcLKnyA1vjfervnPNU4rXcZ4n8gJqh3h
G4+lIS0L5tQXDsaxLWYIZn5VyUKUaQWLUxK9BMvHje9A75p7ErBVDzIcNpOZKvWX
D7nfZ/J8y5H//yxLwdw5ZNO44vivUTIPJ2nFM7R2wnh25fGe+yXBaCdB26VOsGRu
ksWzUcTfzA96lxBivT7a3FCPd77edN6f1gcrFZfvU8c7tZN4L6ROovvqbUtpKMXH
T5RPULIEDTGNSv8U3ToIOcK/3hKrgzKxS7H2JXT9CNiEvhCRzTbcXGVWAb0Algfl
FvcZWpiww26CiFCub7CaFPDBgoTWY7XXCoQTTWPoXrjXKIUpoBJAzQ0hjE2Bn5q9
/yfJ3V4VZ85TDfM8rpOR5LVK96G5NcAfdPoegOOI2L/WVGDa2eKLaDVUr/H1Xz/s
FN+tFVBiZwMYWGrdDCKUjd2TMRT3+l55Zzwng+FRo+CgFgTOeSv669rGi6iYC9tg
gjTyB2V+NSnq7hZDXrjv4cYDXtUQs2CWhvdRLla55OYTypGevrfhh1C6mEbdcQuX
awWRaWc9UiYiNLtsq9fze9ZIRB8nm0prn4BNbqGVqPD+3ltPwUcPSLzghZ6F/L2m
PM62zddJR21uTQVH1RqBnPO/53xABc2p8P2n+iA6bvW5AVHwh8XlP29QnTQXpxXv
xm+9WI8sMBB9Ia0Lo2/m7KNC7VLXCAsbSnN5MChZ4awiVe/bUm3c91Ur3cyh6fQ+
N02uGO6ahexx1JTrGVtGWBNXGbREVFt9s/7KqqWDJSDcyVZycOTnuA5h4zEZ79sC
X5p98HErnH49eU6Wh+awCYLRXmyDkSHYs/fOOvubFpFPSG72CNjugfMCNMXlQye5
MyVm8dBooqOYhL3FB8HefOWYK9d9ORHN6cVym5NsAF/Fdr+Pq5N0hoOd2ep1qdDy
Shjy4ZiVwgEk4zXMANAM5aNYRdHdVkFS0KsW1SQtUkVbcqwSW6k9tUs3vZL8ahE9
V6FWc0aJCiFQ/F8tGJeSWYfzAtcPCW2woq957wX1jKg96yq53S9xTWAaTvIgOGbL
kYHK80zrB729CHv1vdPCkH+4/hEus0CVu0PPXCxB2y+h7l2UitsW9/atOB4IRj5w
f/PGbVhlcIg0bC/zDzAP2eohIU3Jpvc60TdFPUt76nbALFaTYKDemn4yx7xHOq4z
iivp2vSXesW61gLR1CdiAb5GnOipIxCkDicYX/8Dgt3P7L5ACRnsh16eNiaLpOTW
sxLHNUMwewRZ3jIyKc9VSVmZ7dQiqfWhRxf+V2dtkCJToR35jfGjqEKTU8BYQbks
5C6q5eiPyOur08SM4Nf/OfwfrpDG6u0CxzMhqeISsL4=
`protect END_PROTECTED
