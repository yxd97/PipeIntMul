`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IfjUo7WcJxbZZ7pkTog/J64hm+nY0hrl01lKLw1y4NZEX2kwVRElW4Vt4SpvNLor
H3/2EQfd6KEM+bKqPedtMphztcpPLhPjnVsUw2tOkprsWKi+ejR2pBqPYcG1uTLS
tqluUCvAM3jMambWdF3LHA==
`protect END_PROTECTED
