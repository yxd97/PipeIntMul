`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z1JsR4wvs+99jTKyk1LROE7Bd31FUhTjzF0YZh08hnOeI8jQIJbH/AUGlx++Cb3a
exCJ3hbPuIvD81Ov8S/IlWxY4wh/QPLgCNNqSbIuSGw5hOu2B71jHuEx0yCEfp3U
gvUPgqmo7geofb1wRuVJRRgCihps581eVyj7TBWsTP5oZQ0oANEnQ1z83sfcXKi0
3tp3wPq9D6jpzL25c9AjKTwii5xYR23shPOf08msw6fMytmkIUPF5pUEy3q5TtTy
d1IAIE1LSa4zocq0KAZH5JA4y+JipS+YR2iBcluh26WYbBz3MHqN1Z4D2JDu0bSZ
FMQXG98CoKHbDHlM3Vt4NhEU37Dx7S97ccJZHT7TtR0H4CghEagTDVgQuzpV076X
FIu7dsuQCeukXNyWXSaA81ZQ988+gApF5BAySYJ6dtsTrVBEopSgslE+ZbSJwsKA
LSecbMA3goZjhmZ+0HcbLOMmYhJZrsJShPu+dPNllglCXxnrFY7Urt5mR1j7metj
Fm6YGMTEfLXZ9M4t+L1C4EGUufJbAtkBYYBKw1EsX/CJoxf8hlrKNICkp4rQ59vO
`protect END_PROTECTED
