`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jnk7iQlvaN/yhvQbcYXEmf5dzQOOz5BRybyT3mVp6hULqGI7viKEWAxB/w1yuNKW
3H2J9D1pGfL6wJSbNIABtIdPFoarneRiwoerxczp44xXJCFNXIdix63Bdx5LxKso
rMdTP86bVguNIzbKApYM3dAkJSwzPmulO2isEJCVNmeIwkgli/KJmbVwc82BxIuS
S0az8Ic+hd3N7m2cC7Wa9P1GAuh75NuHwZardYzwiTpskDP+U31+U+S3CiLYf+Xo
YD2zTvJTLrtrVPaAtND9qI0FBgrnrAP64TjBLyG7brs=
`protect END_PROTECTED
