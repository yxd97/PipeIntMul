`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gsC6H2wNKqIqLIWdSBuQStHp6z7vYaH7NvDDedziWPM6gVf2BfHENSQSLJmUp28q
xW2dDu1Qix4EAny/RC6tLjHlDNbxcBGflAorwElfkVfgEr36kwwuSk14KBWAkxMy
mLi26RIR5MrBnzO68tLF84XslQ44FrwKtEi1996NVlbCyUJu3CxKBzUJEiyROe/2
ocCqGBcs8XYQWuRvQjk1TDnGhadYtQhSMbYZJETf7pheoO1kaV5UcAbdoDdfrx1H
AWvbLdfoUMV38khm8ripTy1JmFsBfeQH6oJDmWmeMPyEVlTQLrcK5DoEWjpbtLm1
TDJXmojmPvItkIPRmImhYV0OAZQ83fQ60YlnokGiIX6j8U2uwl5Q4ZqDk1aCHAEr
dPO65/8UhQJdshk9Lfilki9/3WwMnhQxVTwZ3yZ5n0/gCYpUNUehyUXr+h+X9T3i
9FBkt16Yv7YhFoCWVxU4+CDhLdI0thjJca2aQ32qx9tbCqePt2n5cJEQlB5bZIBf
Ft3RoshEnXNXiWndkSukrrYjLTjnEn1NrNv6KJFHOiScLGW+EtloVdi511WCQoSK
f634elW82gILjiA1oimqMAjoKBU+tu3HtMUbj9irbE1Ar9iykJp/kMNEwyOOnIcJ
IlpVb8crXVBsnDF3Wmbusw==
`protect END_PROTECTED
