`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nWjn593ty8qU8EpH+R7KQTOQzVDCAj5vx+9lr9qZNJgk2tP8WNNRVa8OehuvLIw9
NM3FGMBB2lBPiCW8LkNMfyd7pN947ayr+uRV+1WtzSnnakUXpSH1rLWK1r6HF3Ig
l3M03upN0o14wig5RhVYl51iown3UlBOmfjQm2pizwbEd/jVG/CgHf7HGodV1X1g
mgweUx8Y8m6x+mS+Hfu7P92GFhvE4dR+N3Ac4Ngbu1LaYA5gX9PVoNMRkz85Y/Eu
pU8C1r+EELr/2gpB2On7TajbbJhvBunENXYUNh549jMrjmN/7oCyHXkGFArYZIBG
xz/ct7XBwbNttBZcQzJswgJGG3M+fbKJ/N/WhASlqOeFAVE4R9+R83g5qOrm9EtW
bguGhu25UnxY6icZlJM9ZFPqc4aczr9DcHkeqe107utUXB+2DS9j3JD4VQussTy+
jpf5yKCXGdZMnhWk//cn99iWmGeAKoXInsACvUmU6O8=
`protect END_PROTECTED
