`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aCJn/VRLgFMQTd1n+fW47K67kfAewms7Omdoo5Xz6ihiu1wcr2FkLwjEyg0xf0Mv
1rLMIpvlSBj4vH3UorOqKdBPTETJXaUIM5LK/ujcd37Wa8OeCkXsr7uKqcRN36yH
9J0F5LsbBXt/1e/4i0lxLQ==
`protect END_PROTECTED
