`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jAs7HSGo5Ql3mhMOquiELPC9SFXipSDMY6eIuqmIr4qlaChkMQ4YdTPePSb+/uFQ
1E422f1lpM0ebzipJQ6DgOqwz8qrgq4olpr22Jn1bqTL3lfDFE5479x04DCeYJVo
AvDUAqP8EVKshIhHqGfMZs2fDrWonR0yzNDfE7vDmlFeg6tOkZ8gUynwaVj1Uk+2
9XKMuBm860LGXvOkodUCVxIBEFAX8DEmZV7f8bprUdx7LEHOLlMkm7YldTaHBpUb
2AkNMcEfObg3Q9PL2D6L+9kjzDfd81/2YpXsx6NCIWsyFf/M3iqDRfYREPfhxuhQ
UFJtEYiwMM/984utRv2KpxjGHJHz/5nuBYrsIday6974AjIHPJhIvnC4/3wFKDIi
FcRuiecjDhmYZ3z0OVFrmaGY5pA0Z7dBVSoUPfaFwI2z1Fuqgpth8oBnnPSycZVU
yy8mVVlIg7EPBf8MLYRqW4krT6RmjFgOFKy5/WnO5oO5kM6lGR0FhA5JdQ8jZ9P0
m9PgUSfX7NRyF1U9qp9iNJh7X1lhRl8cVAPuEfnXAX0vQqUJ1P1/zNWT2tRcC9pb
0TIGjC63JaHTrgMdEaohmA==
`protect END_PROTECTED
