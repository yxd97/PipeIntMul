`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNv61X7j9llQ8LbTerBAdu+6OFdBYQZXPJ48pmJhkoxWkcvbHioY0N6Aeb/+RnI4
aVnxbTo6asU/2UiWmJOg0ZZoCCvOmekrQE1CPyUEy63NpVfUTgtu7p0QKqTE54rz
LpX3UEBG7GoX1TZ05yYW5vp59tHeQ8F2hbc3DvIcJGXlf06wku+yOUSQrE4d6coT
Y+R9RTLmZv5y31/2Yvrs/qaUIRkwwyPq74R1HR5DCNLuERDVSgo+BpbCstNjJaLx
x0XVICkrxyVtConZzLqs+w4guIzsaf9XJVth8tbnM9s=
`protect END_PROTECTED
