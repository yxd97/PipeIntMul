`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Ku3vKbrQgKvEny71IeS118NskMFqYEbkvxyT6TvkSDYMgDkqId1ggH+hv5pBWA2
CpBDv13abh7gWtijvK8nXsnEoQ7kS/Cy5LMvyRaKLmZgk4eIIiyYlttxAUlfLAQM
WKubzTFhDNqqzbTK2dkxs31BXZp6S/f/lzAlw/4597ooA3eJxyt4wf1y+jNgQh8x
GmJpbEjC/gkRm3KRKssZ8cAJE9sWpT7IfJbeJ2DgpMwRgr6YFZyeqc4a49Ei17OR
qdvQ5Jr5TBFFpnelX3FPbtFkl3k3UNGfOhjJhSjRTnmh4kEAiamkBPzacP8vG76C
`protect END_PROTECTED
