`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pTqufhoFxBkD56SGQ1X+tzWlxq1AHBLEbymwXm7biC9LIyIQdJiab+CxuBqXJlgQ
ugQ0UEXGvK6rwyQWl1SNE0pXnG+LcrGo/IDor0IMZa19oS76q1dC3iWUE8DCP0mj
+TuV+4B6WOiCbS0UDTTJuc0/wuV5AvwwlAgnC7r3mN/puxBsqnNeGJwW08auRNqO
vO3bjvNJzRdzSRbr3Eokg/w3/mP5lMU3J+Lvc9sb4tChUHRjue+Ju6XhBzo0flrp
fau+hjuTTI4iMnS4ViGGyd3LGC9uQ6dKlA+0yXgFj4PB2v5lfPtPPHmfPIoGm4WL
KSWBLslpV0RyKmgmRpMGImcesrKuSkmv2oPudW93UGoUthlOc9vuANsczcDAdSHI
LzbdorDkhKDjgvDcAmVTC6ugzyREodam8s/EsmoMqs7In+kwWERDkIOxGgBCIlnl
mb16a3r8FqDzypMyjejixyvMk7MAtp9hkx0ZLFLpoCYWtqPFqf7XaCvA6Spmr7oq
sEIxudHsz4pXZCI26f2J4AilndlH1OcUrVOEVNqIeE/j5vWzEFiEoDWMiEPjmp5G
J5GIRGqt+fHbPSgwvrx16gABUgqp44AAfWX2OnJ2u/6j91nkP9OMKVz4qc7J3bF2
UPOLhhOm+xQceCl1+lvxWbctdO/XNcLFeTFwZlp/MgT7oMq5FYK7sUXh4t6GtB48
q5QwL2Of8UmangwNvn4YJTHSrDEr3mYAjFvH/7jw7mJ38ZVnt23Q9ze+L95zrbEO
jetoOCpiBqARAS6lOlZaUw9DlXqWdEBPIAbPvjArCndsGaAqUVUXtX5XXjfh4AP4
wDWnszkEglETZIGu6tDyCqkmUvOYrvuO5wfHnDxv/WSDmoSUPFzY403mlMLpjMtg
q3VI2tnivKltLxqGRc/0koAO6/oxNKT694kakJp/xVt8q/r+RVww+n0pAF722Ufv
`protect END_PROTECTED
