`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSapiTS4v6QzDNoiwHkB5iKvrn7TigeT8dH8lQXyLnTT4yP9ujyRzubEgSYbbD2V
aT05tXBEL05nwfWs8Us5JDYAvo0kQqcshgrjD5ePoyDmmmay3a91s2uZJpfXg0bE
kFpTq+50n71iXQ4+nUXhX6g5WrYFd+bsvWam2ffrePN9aapn5Fdw90ZxU/G4hlRW
VNoYYRqJQhkIs52+br9TKrP7iflHnii4DtisMpRINTtPdFhcm7yCB6WfRzOk0FGL
dz636vIrTujTgen9XuX2B5OSBUmA1X/GDeaOd+WuEThtFivHC/exCtC+fHIQhfma
6y5HXCUR2b48AVBkXVKA8gcWQz5JM3eJWyJALaCNafz6k8LhMmI46kc0QfSHycSH
cT5GgLPq9A1LFnH4xr1scw5RTWJZbYYM9vwprFMe0Z2OJHcg6nE1WlchNCdJT6BB
ohxW7WjEeoy+tbITYhJ66G/VgR4uord6CcUTSFV5ZiDQrx/bLxBgGjbkxs9xo7NM
ekJrGbyI+UoDpwdywdAGBUobt9apo63ppqF0on4gn7nwCKjpckH9YDMice8oWBSK
mXzwj/4PAEShbB5MgmAYMGo230l+YVEYdAsRXt0NlJPGz3w2voZc6R4vodXRZAyz
4I3TT2YJxtTOPnltdDHAuGe4mvewLguSsC9HInpDiowhvwVT3whD9lQSoZduZRJQ
sPHZrqwxUzfrAHcFokytcYrlCLYbue/Jq7jFZeXMWA4=
`protect END_PROTECTED
