`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zIbRKvXwPAB3BZNr7T2Ro33we6MUagcYP4EuQRwV+Uz01n9WqjH5Ddk9Vl7GwTdr
5r9SmyeqZMerosEcQwtwr4KNnlTn/enNh1Nr9LiU+Z8T0CluL/xoAo/GVMUG0wIf
UFRuNMHcUIhbqJdNiKvu+u1Iy6Ya12XC8XV8k/wRnBXmx1DhTmo3j/zNCYnHEsvV
wrWKdNZS/Moz+PT8GimW2cVX8uM01eTo64ISZZzKG1c8lyJBbPvaAMNm66gJVus8
ulUzgACHAcU//Wk0KKyVzvtXu/SJXsxyC25d6+KbH+B8qChdPVNhLZHkoZ7SLEsU
lhnbq/Im56MnK/t9GzrfnvL8buWw+ciwN/jOfHI1mntmJlMsv7QAdDrSLEXk3Ka8
9m0unZlKgov/YeJjAnNBF47wWr2PQeRux2RxTxKPOISMqcqkwmdnIYTetXkAncO9
vYTh/2YlpoGi7542BC1FRP5fBFFt9KkvxEGDrSi6yUCxaa6eeXYeY+YWANxyVoqG
T/LCo+QRXy3RKoOwkqbSDE/1MeZA6h+wH2/1w2+fuahabGWyX9R9S16PX7rTrL1x
LqZ0t9gIW2SqX/NOIqFpvgKyHp24PBhjMi+qUgn8vqUdhviuzCB9YW/MFr0nhLuu
lmCl9wVCxuDQXcGDO8hDp89A+GvMIr1pEruE0qXeZ7YiqHgm6ZDIIDn4QMmDu25V
rR5RDzS6Lwa1hq9m4EKl4syI5xMmTK8DXWbBLmMny3IOFQ4RBWbCdYoi5AScxc6a
l70ZgFj8hAI0VaWmH7W9UicKKEMK1ZOJvPtP2BquogQxceFwq1ZvUad1B6S1Ff2r
dm5De4OfuU4lFUZq79Tzy76dPwM003ZhfyziyJYcq+g3W/rhS3Ft6zqCYF7jFz+Z
u/zyUyJwxWKY3s1HGzOrS6wOeLwec3bh1zqWsgCwLSYaYva+qpLulHDqLUQq2Kki
qt/WJaG/Z5fMZJbqiY1mhdzINmxKqHHN2lO/3t7K1FjVdKpdAu9VfdovZE3Y+v0m
yd5fqf7huU3xQEarY1XstOT+Mr2wcc2ImHP2DHqzDp64O5Vsz4qOIBxfUUnLzqUv
awOxeZo77ocZDB+aMHJ062cm/fFybqbW6Kw7uleS/omwNVzD7zJSESDCqS4zlRP1
iCTLRHon1D+tzJpBjH6bkc9SXB1Sq5GXR0Ih65WXva7EeJJoivaRXIDhPMOt06II
4Neq2qJ3bOFNF+VZwxDDjJoMpOJ/s7VId/V5z/arEbBLF9aXOpw5juKsCiJaoU2h
ZTFHFAb4KYhPFAtg8m0K4L2UlzZL56EhNXImeBFj8iEuS2SBHu0Q1p/6ZaVn5NAK
i1SfNE+nWz/TCc2Bo8PsOIX9otmplmolfdX82L6zKPfnsskAmR08swXBejD4JRAq
y7mPWpRqtMee5XO4c/D5iMSMmQNXHR2MjQPns1Jyx0nnpeoCZpnk22sb7qYB0gbO
JY4k4m6GPWxsHm21TUySa0IVQIzyrriKkDjfatS8Ql9BZjbkO9P37fvxIrIvdHuV
su/vz0E3y5NxR3M7L1Fdi3PguO7EZOu+Sv2lQzgTfV4OhaeptwIgWprXLJUUM+kl
evc7zXG6WCW0at1Zvgvt+YgzuWLa5SY2/mN1X9XClA01BhC/D1a5yQV0dfWyvk/c
DHKUgeQgeGV+6B3mAWWA9HbstDfC7KijI2JaUJZPDn/4H6Cy87jafElzeMv3KInQ
WAiFxmQWiRNZzJ66/dkMs1iDkQngnagI8+mRP321/68=
`protect END_PROTECTED
