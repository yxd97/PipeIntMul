`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBgdK00jTYG4TpXYNud69SkIEA/jEwj4NWMT6gVBXRW1ZGLeFw1xCRQB5zc1PMS8
Jk05vAYozknsbxuP3/oo8VeP+TutkkPrOhG2YUNd7F31niNuZ5vTPsCfK24BWvB3
xMzQ5Dro015vSTsShyJeqy1G0+huqkERCRgZb2hUTKl5H2WMV+YfPuzLkEEUP+qJ
OfCFsAhKYLsq7Sc4fNPOr/dxrPruM7fEbbZGADq9eCclOXBMG2d3bmgxthQ86knM
39REkREoPCeBVYYw6EJGunbJXR9zImqw7nuQTvGgURdFgfxlg1eHqzK9YWlorQmm
ROU0oV7B1iINhN6/aGrA4+ikxvufGW9dCjubg9U6oqfdbPVOBQo6uMIu+m2/MSn/
0VQD+CWi0ICKPh3uB52vehgCZWxzsdcy5hDga9GaOuusixuSc6z/y1ORDsBcpa9i
JELgfgUjZ6px2XdJiej5rQ==
`protect END_PROTECTED
