`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ij0rnnN+rP4QeHjMpVq1f2oOkChBCiqRsVvC9CAqZaFoFflJl0Or+7wwUzqwo3N7
cBqA7fX5tNIEWzwhCkVEHF0RgIOA6cxoTzJdQC9R43Va8EX7lW4wFGHr6Y5/QV3I
B2YaBSu/QJLsT8+X6RXwlmPtkCxhUfJnvQ4bsGANrbExpautbUV+vd3QppIJU0/W
9ohtpy45s9su6057hn9O1p24SoINDRTrlJ89Bmx3iACJr6rwlkJdFCNUF9hTO8VV
iOW9EKrtbU2CuDwMyDKeNfF6bogpXFFB0yVAKMQbGmWJdcwo3c4qDRe4hSuPEyjH
94yaJVre0NQLXo8EAQKpIsD0R0qMdPj7R7FpNITPfRH4OthNqDb96KL0EZfA5vUB
QRlJ8ceSE29d8SGznuh6FV5HsCSAH6E7rGtHw0JXcWTVQVbLoaUR7JxfE60DOmEs
uhfyQ07GpNxV/qMdfrHlxgFJg4pK+FRrHXQQyBfIjD/ygdYSE8n3lkQiPv50T/0L
TN+XZWeHJuS9x3Q4dRsS6TJGoI693O8vRBDO08OKP2X086tmHDwMo0/ADL7gGOPw
079pP0GAKGlGGaajgnJ7Kj6aM+3jh3D6iblBeEZmOcjSEjNvCB5Jq+1UdSyEdNiW
jnNVX8crNkGZxAIfEfRmGYl5YiRTTTqFBPYgWOkQYegl0RH+E0kpe7NZ0D6Awbr9
sVRsDf79NTHMHNeYJv8yE2P7Zt9m+cj/ZSjomi0aX4BNcVDjLYRVvJt9SWlDPYDE
64+qmzgrOAb8wUpTDuxHlmENvPtdUUK5iijijlrEE/BW/mPdAs8hbuFP9bh+aNRk
AFWCiidsiEWM2wlxuGxhPHBjxB347+Ld8ugCQvYLPJEZtA8BhVIv1L9gLe3XAVCy
iUxi6rRZdvDCZzAqOBPI63xEMQpVgupjqGpS8b9WjUb9boF2zbtHg3YpbeWoyROk
1uSo3K1CniwxK5LT0MSpgQ==
`protect END_PROTECTED
