`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKOnPCaLbEUNpdeaNhl2tSCPKW2a/pEzW3gq0kwr9Z2iaDPYP4rHN/fLyYgFodVL
ws1LKhgXOWHYTPbw5ea/tYajLjhvl5fzpUVDr4BBeK97y5scF0Y9lzUiQEqOv2U6
8CKcd9c+RudqKat5izc/HFah4HxEaHBeMBXIKaMpM+0N5NlT3hHYIrI1vS3FUeuT
eRdkxaBAb2eqBSR+yLg6xPBpC9Ql1Tj2852Lbjq9wBfsu8ek2heG7FFFQy4Z2vld
kvyMips3QY0VZhABkrfLW0k91WlKi8uARiDmfcll2IabjCk9TKEBuLLXWIfrtis7
B6aig5nHPnItvHG8a77TLlsECXwWfkTfYQdhT8lYacI=
`protect END_PROTECTED
