`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zge7nInm7d4qXP2MmtfHZ7zboc+9nhNQiAZSR4LjAU4o8+W43wKGQs3MPDt148Q5
FTAztVfuahAGVVqKsVxHuhd63qXRSfu+VefHxRu3z52KhKbGLbGdVySOLlSVQ8Bl
2PsHgPzUkkhUe2BWkEqs2jPVZFapJcebgRc8vVRfcAlzwcT7fwHSg1AI1C3kOjI4
TmN957om6Rm7TU2NYYpTLT+6Slxcu/BZCcRafZJicLvvskxPUDaxDRfoTUULskff
HVZoyYSPGT27cWnrJ0SjE3XUfFFp8LnTa4cvr8ZPRrhk8mdvK2h1/Le5RXNq98ZX
IJpYL7GokeL//ErFXYVMPZw88tnosva51CR+X3yYmcLHbwe0RnV/0AjpAMQYnPEU
S+2hc1JmkH/El7aDMackT2hQluYLXbNATK7W3hjhsqdPHvvTow5QKDoBgVjJTYku
5C2voerARqSAAptNkxyezShVmBVDiO9itVDi2K7Pg0dE/UHunPfiPcXtVLeLOqTS
85f85DNVCkzeylI3bTPqd2Yi4PLo/oapwB8MD3a4eZCWdZKY+pIGd0Edp5PZlQhY
zK7iJF09KQUFDXFT5kFg0kOZpvujRPhk8r4JOHzMlHfw43gkTRkQYjzzkyuDuPGB
uCIpknloCZXpeLHT3aIuA/wqv2YU4Y0d30KCeqbvfPff59geE9Zo73OPl6Q4kxNB
4cTmWeqDXpoPXUOcg4u03zeVmvlzgV7PJ2zz9Qtb9GpYTxPKdBulvRETIop6Q8Bb
z4iYe0k57jKW+2MgaONpJKRpvOTlc7MD1x0i6O/1oAlVMl4DHKX8eLDO9s5jBuBb
anta+Rl15YUyHiER10/k5qp0OZzyHWbQ/XF1gAJWfMncIb8DPMi4FUqo4CCj/cWx
Q/m/T5FP6LSLwxtBi0/Y+w==
`protect END_PROTECTED
