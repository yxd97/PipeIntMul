`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J5r4+BCqvifEXTfNVh8I8wVbD6DTQ0lla/oS6tAfgPBRRZj/83LSeV3eGKQK3rsv
P09CvUZ+O8p4+9I66icZEsk1wLqabMDVkHDtHWWfDnp3ewKf8Qnu2DGo8oPxJbg8
UQUx4xOaoyOFHSany8Qi2CjJXbHvKNdEt1ZNTZbWJQ77AqHMuCSmKUkp8F0cZ8HE
7p7LiJC8SRZaMoCsQZSYat8uGTMMcDScjLjlDKTPgh5ylCKvypER0bic3jNH+bJr
WS0PsEAe+QSuyLmA/Ae8jrOmy8OcspJoIof0bPMNE7Rq0b+HtzKSxWq4vu0dMV23
3dOe3P4sLv5ybw5rd5zfp925hp4oMIEClnuVJLj2uh7U+JJaSMPpXa8bBeYFsKnM
2rM38MPhhdYQ2RUjJDyqKp9thDnJzRuwuOUovEtz31irej/25/vFPs7UYEeTv69H
hqHCmnAgVKBWWsx8idgcHBFJTpotBvgqeD4jhHEZ7WL7na3TD96dNcld7FlXBxTZ
bIEsZaY4GbRY9LiViIOH0J/x5xP9MUSvuZXdeAHj0yrQ5UDjKJFVBS3WzXMeeHrC
HQy1C/vw9G1JkgGrCTKMbsqvpg7Qg8CinRvlWpATRlN7Jh5QKiTfLyilf0ulbMbu
FL4NaQjEsN/0z9AVXCEdyjgPW2rX+oeDiNHrxf0q4gyZZKrKIp5aycvsjgnPAXCr
5icSfCGuDi4nH9KjYemlGohZ8k3PvTAc+KxeUs26MPNDD0FeZaU1J1GibnOIhOw1
Eu/PGmcVWrFaiAzYMgOruRV6+m4qj44lLfuY3kMi99Ieu2YKaeCj3/tUSBQI0W3J
537AUd07BIJcadmqeU+sOliuARd8iHQxbzC0pR0tP1xxcUmDdOH5YdoXcqaHV91e
oZiLmwWVVUtihSt4QqPx5g==
`protect END_PROTECTED
