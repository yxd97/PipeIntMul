`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/KDEdSik8hN9LsclaEADHks0Njf4BCWMGxyK04nO3R6zSxY//yEfLrY+ZUdq6um
m1iSW8lWz2CHYveu03BEbsw7FrQ2xSyc4FuxaPxw+6hnOR7RYZZ03FhAqLBnkVhA
4p1EN8B+mn6bWMnzKT1j7HTToGWqDSnTUJ9LIUzYLVN4Ss1W9pBi2L6DeW6gMVr1
Eib2fCmilRNhUCD66xtscKhpCtAkotheLC4BZozXeZS/obrvSu5b0H96mv0MeOLb
t32Ma1HRiB76UCZ81Mu3PO3G4ZtcBEAsLsUemZtOK+O93BFrX5vjdVFEbZC4Zc2E
vxrVt+kp7ejyqi9cTW9H/1RGE7+Ge4EZmVpeg2rQx7Lrz0KVnnjfQZ1VAqyU/Zxp
HZg1BUUHrGyozDGO/50MWQ==
`protect END_PROTECTED
