`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
net5BaW58AT5RDWx+Arr9MRRCu7xHxnm2nKvAskVteV1YIHQLRxFHhg6ppIJHyfV
o9X7PnsK+hPjqCJX+wPboAjYySiNWe19se6Kc4sUKVfvGotDXEbimxvSnUlbANkB
yOs1pWEg9gLBhH2YJycCfoZnMIbeyP1OULErchD8fNEx7rWI4giinLsEIojA7xFs
j6nXYxaD6MsEJqY39l2cB63WGEI4tqS0rFnoQX/MjkWjvW1tOB5ymsU0u8DpEHAn
TuW1ZgtidH/Mi84um2H0TKdqE0y7axUzk7sEStna5O311bqQuR49BFepELT1rKID
S84zElH/7tJMYPI6jYHEaYdmSBjqNVdxKS7cEM83KyctI6ZcfDpPvdNQcOR46xTu
XRkGYut2FezUuxJIEaQohw896+dZ10R1muPBC2ea5/ISVgLkCr7yf3mOIuHsRt01
`protect END_PROTECTED
