`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEUGHL+/TL9nnxQ0HqvV1kIvOblNApH0W2GVfIUscr55+9eo1KQPojt5T1NtWM5C
4wau2hOkBlYnovSJ/l5noZ05yJ8+D7f/iJS2PfQe+8OobdpJtnVW/RKboxG4ef/H
2FCrkJBvyx1DXblpY/YSe95eq4B61/HLDkW/G2KnO/oJBRF4IJcp7dTfhdLzjgQr
ZVawgZZbTqrohlorEzH/hO4IEFwqTIIma7Nc8fz1MHY8aXqEfXnAl5gs03XyfjdY
jf3wVc9opZv4FYG2xT/+5/9aiUum3yv6eFYHsxX6Wurp3337ZYdinMSm8M3aTTDg
yuK6cDRixViI1PnBt9/2DAhtCueWj07HXE851tT8b2jDAeYnZMfnWrtpWvDD/nu+
v7X3seFV+wt+bgQdQkgLFjKgHPLArHFtao5+WD5CUGOBzv16S8EWy9Ef9KwNPg3W
WpFu6D1PsTI6cJ0RU/oRGZAMZ+G+GbwKVrxeZFU6fLPudh53+7DfqpfeRuHtNstH
MtzTRkxeVKBhCE0x4T0Z3kPoRQCOS7m3563HL6Hnr8G7yZn6bcvFgg870eNHXaV2
`protect END_PROTECTED
