`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HUW1pp5IFUsVhncxOUbGF61AwwqWbxsvWc7bvyGUp1qeJdVHk9b2Y3AnFRtPfaqX
e1Seuv5+1jc2Ao+xIf/bSAV7cxporeZ1ts148WTN1D4UTha60n7n6sv3ykmCkARv
LiLX7Fiwk+B99HTSA6P4Wbtnbnx8YG8hcRT1OXzVoTHmYGgSPomBSod6I7LXBuGX
bciyBHl/eMui8VeTDv7NmMiW+1YnR3b7WixiJCIqszMowd62vWJLR+xBJYaz4POY
iAXhB8runEG5WfOSnh5O+aT/+kMf6fcF7pE8N5z73YVFKne9GDFqyoj6LF6T72Ap
VjkoQv2GWEDhNVm9rwh6//bdH25T5Qm1ZVlZnSFMIzLgAkMa1k8lpl06tMdDK6pN
xdRR664yz4fcRZo1QPI48CZDw5kZwi4RpC/AZ/NH84gr8wDJr7K5LPUJJhMd3kqK
Hdt+UizQ+UZscxcs9vyHH1iXVbfxF8lUPEyGdBGF16y3RP42MlbjQUvAYxaOcXb5
bmnulrcTMsp+eBFap5wzk8y0MBrPnUMxc53POEuf00c/V0G+l+2ojjD0M1/Orvdx
`protect END_PROTECTED
