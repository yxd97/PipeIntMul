`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69+W61bJiZvXZ4nF33WTT5B10EWDQXob8qSvw9fn5hzYt8Zpzqn9uC1qQ1rNY0Pk
AwXSy/XbCQDmoFY1GnDnYwGqWRP5VYqDxvQ/dMJAOBIBb0oKW4egI1sVCd5ZIkcF
AheTSwj6bgMFItPrP5br+IIcO5KrZS3mkBgOsKC0u4TluWd2p7xIn3anh93eDCpd
kcbOk5j38lUoP95rLewmD/1LjvxuZV3ZTo4mcDVpZDrbbZhUkRN0LJ4+rZ20Ri4v
8jrWq8WcsnEZtv5sSC9luV22CsOXybxEaVnPmPZQsFBb+D0tOQ8Nx/CWh9qkthRy
6Lo4Cj7tHLkB7UjC0ydwjYvp2y3Tnc9IRljIUo2tyCfFaLWYI96TA/Lx9DTUge3f
9QLDyHdsYs7ovegU6qFLx+zPYJqOHK/CxjDhtEa0uPSdFLSODYpwq+cXQOqMafSO
q511dnhh59W/6dX9IQbmWAa7zB7qWN/NAV50mD8h+LoK7esPd6gC1jFfOKNnBnIV
CfO+ddEcoixssimoAn7AynV0cybsmvcSFpRaGPawrEDbQSwXWOpaTwqpY5j6NW6N
fqBvWhgPVmt0z2jmQAphc0d2BDoqEa6ev1kgk+O9L8jKQ9rh4eTNSfg8ySFO9a9/
YkEu4eSWyKEEOW2mPLT09qc+FaaP5KHm8Fd8JybEHHn32A0/TlA3SWEbHaD/1AUK
NzcpziL89sUN46IAZjncx3ju8M9LDQxGYJ63cEFCtCurwy1PqPtKCfa7AIity+aM
pSLDSDGMsMWSXnCbCTsfb32iOl4ZCF2M64ZzgP63B+fR+wiBEBNJVybC0APV2wrW
k84Q/kIGU8AqboZZEZQS4S0ra+eKnswQk8UPGooUzEHANzAYmftPB0ApdNY5q7zW
mAdEkcA312P/16n2QXNu9f3HqB6crVcsz79ux3BdWwRHCB7kny9QtaMdaLgVt+0U
e3vO654p/98MKnDZY+cfxsYzlf9lCMEURwzpYTo9HijQciyKsz+SeX/z8sskn4Pe
wXmR+DDQwvSdbHGKYXCIk2EtfGdIybryIhk0i5VT1fkYRAASmr5IHKtu5nlQNcDJ
uMCaOhysBC8G4zrDsh4vUHdfZ5T9LGFk1R4tkiSnoyBgDQn0H79XgV0LdOzpLfJr
z2Om1t0+Fm5QsmCDiyGCwxWdeZ9u/3R+Ea3qdbhiz1gFvABbnkAqD9Qn3PyfhaRb
N04dRoLr7LABJocABH1lHPaF8YhaNBsiFtZb0bBhgKgw8JZZpJvsBXU+zVuH7e2c
P7yUFLOsWezQH0b7fL+/dhR4f3WeFUj9uzxYGfOLulIqXXbkuQ7FSVv64Lo4iuDY
7HEA2QTM/7IXmJZK5kU8YiVHHGI4xydzEiGDNmpOgLU=
`protect END_PROTECTED
