`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xMGSOd47bevVx9SPyJdFuCmTbih35abhPNo30okomjWMASC/Jv8dLDZWCMHIJ2wF
7X6O8SKiOc9ygtfLhT9r3sE+4wULtz/8SiL2OG6rFZdSBc97mmXzI61V1s2fS+Km
Z979MS+LHUhXgXsIrV3l3ZSwMM0ckaZKAmKxDCiw9NKRBriLeInaoeH5qrmfLNPf
X8CU8TIe9s+iwDtbDX8KRzI6+2LhINBZq67KmAI7c3kORiX11L3kmJZ/zjAXcYr0
eALrzcnJHc2Wq5MOPxyZhqexmtCiym6IM9GKAJCyVDPl/KYpPFiBHdiXa4woXVGl
0yIIFKdff91MDGAyvELAXQ==
`protect END_PROTECTED
