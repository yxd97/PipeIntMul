`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rW6N2N0HxaNXUYit2L5E4sjNt2z2OkKrHJJOhGdbxQnCOm60yt1LU1BanaskBU4O
hIYuAl4LYQJP3SrhrC5+2StEAuQDAE2N5ez425laLGe88OjLValuO+w9d4bDkUl/
Q2FGkc0eQ1ormG9gPcETyi0L613SnmqYgRbo/ahtcA5J1n7p22zdohT8kXGrwPN4
mwyUP7J2ZaNxRagkjif7YHVvL0YMjUenQKqQpBQoMlta51KrQfTU3HUEfSavzOFq
wzJgcrViPvbWcJB+G5m/vv1a1thKFUxPBBOguqdkxsj13aw1vW/zVxlgBjhkCM2c
CsiSLTHEZjq/ztJXzk1mYzjm8OYgDxhEw/H57WZxgLr4jOrKaWe4RPPM+ZB1M96D
Gg/5UnRaEuc6GsacYfL4DwPzbN8DQzUIWXlvpNZG9quHgwrkb+hLnd63IcTKemm3
MhUGhIheVuxPK8m9Oz09j8V1k4cXMf+WPSnEGymsHSKHDkGo+rrMgTMrqsPBFdyV
qyA6ql3nB0lDlfg4R6wB+md5KmvDcretdBpj2yRIf0s=
`protect END_PROTECTED
