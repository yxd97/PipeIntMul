`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VaHmiq3FESM7ywDlMqMwWHZjDZnrdzuCYv3c9Qdl+8/6/4udMaX5JJW3icufvnV
gvf4gGm4OxmW9Mkzmhww85RvTlBlVdmsd3wi4Y5zmKp38NmYLY+k+GMR4S9slUUI
YJIrWJ4xzvCL+3gd/SiehMe/O+HUaq3x6nXW8NUisIdOmPQyzo7iq+jnrSK0Xx7r
Wzs8QDabv7SsnxN1lM8NfiYZ4DCwJGzhcGbTinBipUgTtBQonfm998A8iZXbwd1T
FbYTPQHnSwv6Ea9qI/l8RaNU2rQR9FX/gwFb2SK+sWDlsILkIvUNVltbBa9cla/V
lbiy1kGpO7AUIdhlZpvO7Uyj8uoJMP23x62DOJe5XD2DtnEOEZ01FVq7n2b7ZBFi
fNr6vWtglc2TVQ7DFloALJOlv24ymqfR0wuc6OHcggzhRWZ5wRvCjNi0Gq3n1wTB
LTVOHFgQ8t/TGDEZqZeIaZMZoyz+v7bjFM2ky8FqGIPr3p5EPKmq6s4MAVAMgi2Y
hNP8JEYQa17tFxzq4aCsC7HQireRgHn8bGwiKe1UzmwjBclFW3w1Skg/ecrpX6CA
foinitPJH6Gk9Ps84/7/lvpNmO+IRyHUXLiDeAZKyEZiRSrcP4ZaMYo9cTJuMOxa
/zuG2rfcjrIr4e/7kwqds6Llrx4440ikHfOx20d5lzFZLdZPMj63RaCN3cZvv/UD
6T3h6p0Y8BCX9eV/pDB7TDMLVBoM9HxpW8ZUsunpwlkYAds8S2257uvmOnA91Qm4
7wBpjAH2SRlI9V/pZ2CvT2Jy4EgaqgpxiW90wqxK2KqE83QsOhrOeFhZCeSR10va
X3eB1nwHc69ZvU4H/Gum1Mqbox8NqQ5ytvNAtmRUODQEanYDHp1fDioc6SA0c8N3
nlyLpWUfQuc6bpWgPJ8r8iOQwqrKTqWtxABG/y3DvpdACgKcNyLbznf8NCUVyWqr
T2fJNow2zwfwwcHl5S5DYb/pCw0mB1MlEbYewIWlG/ItnuYyDJOc1Ow4GjJm29Ca
lMIpQ7dNtln2cYgg4e2Bg6kGc5Df+03sGdK9bZVNGuVhRbUKb03KMiaf5u+m2txg
80CnmUs/QVJFA5khADUkmuNLLMRqZuvj5zbzBb9mHn1LSQUN3VSwgNd7aiim9DN6
8l2BZ1GmeqWZueZ5gSJIf427SX3oeREbGnglX9b4k05Bw+jWaVKIzux1DP+YNEQd
Gp8DSb+wPukKaqhVAsOBk++HNI8rh6mOVQr4miofSdEPuHAyeyz6KnA4fKFbhWkf
A2barJfL0OCxNUS8LUFYMA0DkbGVGOeigt+kkj2W0v2kjKA5/lMOmt6pW/HxMWI3
zbLbueYue0LwTYLq6AThTk5TCuaV2T7tJHAbVULG4K0NdvAYv3ttnwFLTNEJOD5t
40MJxK5hpr/SVmnhxa+ftH3L1m6QMsdseWkWAkf0FBf6kY/hQ62wl7jqc1flDvmg
7kZlPZhCskKmGNABs6SpmM9Up1ZGqgzDUf5YZdK+vkZjlEY3wgEKYSTXE4PscIHA
3STJiRVk6mwp3XBDIkAQRqlD1/KxHElpftOzTsl98PlcCZdLmSCy9AOPIpu0DPqQ
lBCOT9PucwNtoSLyRF3lKG9x7y3sE5PnC8fgP5OK03I2pvG/jqQYSnEoYVh4xweg
Y975L2C6f4ZRKXZvyrEOMG3E8bD3lpr/X6kMU8a1IXDkM5381glKuRDKD5iXGdfR
oKFcn1qDWy89+OG0w0Tx86dNlB9hxI97QKz/an+JcHNRBDz2hnii2pEUHl1ixKej
ah0nbeCejn4WWvCYi3smxPXB+TDtADqzNqlIb9+Kdw3sy02RA9K8wQivhuzoKlmY
87aoUJY1nao3pICTzTDpn7HNhxtplAlFzdSfmUUK+rUI2oSeSWequchdUdXUofhE
Un3HTrB/s6TjCSUyd5r43DmmXTf7KuNjbYp4FI6qfI9WNzt0obF/ikRcS425Js7R
ym0U2YDnwG6A77Oea1HG3ezi+b3y3RMvsK3mHpqFdj9DsO1Aylz/rPWkLuOgilAG
KM3kNzE4a8sJQUZheEgjZ3LU3jqRSYk3Wa3YcdRCrLx01EPAshjCGWtbIKOZFDoa
MKODnLjkv5qCVADlTethgsCA34l90bazElpLxIj670gzShEW44oyhtyqc8ADXiAo
HNhXCVzK9vAAy1gy3Q1FYeFrdzUtTRFzKe6FXCd2FpiA0Gk84UaIi26LCUfQDVjH
tyRAl+ku5kejfM69eyqt+KkE19PpXj2zBdeWh4MY2RFfPIiZh3Tp3fkuvPaB2WDq
q4KeLcRAVX4kKcLFCO5jU8xf1yMiTtjBoRnVbx+Ppo6L9W6Ta0h6KmxEeWtVbMkf
xYB5vbWit6CNCFQi/uXN0c6YLTzyTJ043+U/rjMABI2FJLr2YvYpSu2SFdeqpwC7
qoJS3Bt94qssVQf/oOH2SJbQ/kI8ab1lBBlIdGv43P8W71uhsOVWgEdeP/o8gy7H
z/pkRsCNBoaQNVRsLPXEwdesjEtjmKObLhGVuNOc6WGf7vIo68couR5UbMe53Gn2
Q2nY+16XoMMmtFdygnVogs4J/vVA7glxNMCEkJnW63FOoSpTvIE6YXqtZh/x6omI
F4w0vXyMNt9qMzkMT4972IE4iFj9YL6Y3N7Y6E2K/fF5WX62hG64xzbMs/YfWJcv
gPo0l2MMrbI2IIvJGnyGqY/Y5TvNV0T0uTt4rfJJy7l1aj/z1p48YoN3HRotD/Wy
94p1Hc/c4ZLt9nicct78kWIqvq1MvkE6n/X/Sy/cKtvm8tMH7/ftEaleqTgW9Jr4
ovvD++VLoiZH1O9Z71j3D4ja4d6bvgfX5LV4rzxkD7k1bPhnd/zp/kcedWSIsz3J
v55jGrQD5PidGfHpur92L32m47yKd0f6ju+SfqCaVdK/yCPAm97mAukx7Kz9pTjO
ZMMHjinJAwUFVs4fh3XGpF1Guh/WkxND1RZv5s+vTjG/3vvMxy5ltEiVh+09Vx5c
RaV4mXjr98se/pVGER0xqUld3SDIJdRJPF+7XypZt9yOLrfQdOyUSavX+i8yxUEl
B2MrWH9tc9CVlZoaV6mebgcvGLhrWtATl4tni6x8wxQ/sGeyxFNM0j0sndp71Y19
wdzTAGynX6K0+mLNoLAuEdBTJyYrVFShCU8XndQy1rbGBHEd8V098Evv1GdhIHWD
ckUdrvRKWASyFybjFiBizcOtBwfgo4a/R+MRYokE14kQPkXtiZfPT5uIhl2qMxVj
Vyi+0GZn+cSKSkyChAoghyhsaCSAzJbK1buFMnH/OCZ1AF6VaHBLDLmhDin/G4+Z
IrLQcdksRGR1db17O0fdaFm8axwlx2bJY1XCa4MS0/QrcmcidRo+CIo6cbT1i2dF
nc+GKkSCo9EUeZiMG9aNNZPwdKHDTNwbEqdB71b5IIE3IXdOEcuKsUbPeVHnD/hk
iT7SRaeOz2lHbD06C+eA8TKBGsxWUkj0JQFoUlfCfR8MVNe/kC7H2nGq6zndhx8h
IL0Fo0EbEzV1ABkI3mdnuBqtVRfSst/CKDWjbaQOUpGr++JR1dcaqaHKW4i1vMr8
jrrYKvdaQymNnVgkOELLQXfez6O4WATJLqolLzDTqALVLKkIqoGbz2v8TdN6rAqA
EwkZVdoCMA9cgpIFC7RcvNeaJavrUIDOmst7IHkCPdKTX/TXLgFvK3BHKmKgZNg/
0ByBsDphCIdLZVXdgu6+SyORrHoQQ/cCA3ZAeIDxTPq8e0d1lddim8XbuHhRrduh
NZn+Ya1fDQorw021IhZpK7VMGDmtskj/Huahmr5hfRwXJQ8/bSH6T90aNhyv3FdV
ZjoASm2uM4PW9BeteNHgJmA8j4yLXdIcrI/pFbxwfRym7tcd6pXgqC+FWXQHjLVf
AKbcPec5yZ0zQ5YHnax/D5aLJIo1gpByoH15DlYy3Ilv3SYGnGGg1nImyQfJb24o
VoEgj78N+5jvo7uoqYuRkfHb1+go3ehCtiwwzkxpSyFeVAXaXTcjgxwgzbDOe/Z8
oZYDxhyl24yC8/hh+dh9E0tKCWT89n5zDhsg7aubronHiP7lIhFzWYNGIWiEVFe7
AEFExatkOZRhTNqkCxnq+SFmMujIxyDbSadVebDlf1j9kL73VR4m1re7Hi6BySMc
5M44HcOFk8v/C0kEzUBJUYhTO5ynrS4VAhszpBp7Kj4Y91/a0pUAmbqGcjLT28wa
uYaGv1ltmdLQum8nKAVHYaVXD2G6mOIuAH+MDgbLBB5pDPTuCYXW+Ed4OrZ9VHuS
FyuKaaLTIQ3fWICmPSVK+ifxNopyO3U8cdWg7OfDNwwoe3oiowTEUMqiH3iKsiCh
VinquCiAfq9D1w3rMJ9LlaeIF9Rve1IOm+0CtaYNWL3mDUV3AmGRLQ1QdRWplT95
Xa0VGGmhAC/PmXgruuOLJ+1ok3DPFONwK1RCrCwt2Hy54wI4cVhGArt1rr6EzOJT
57+vd+9YC7EPT9EqEjOc2sIJG7mO0Kqe/RzrFZATMhOwNBDUNCpQclf3QpecL7he
Qy96CNKHO45mQkIIOBVGppKg7Ci58w1e5pY67vZBGIJ0knYgVu1paTKemZpMQh0e
+IyLE0cuIJTjb9cDEKar2WIMMg3qwMmwb52juReGoHIOhGxJ45pQJDPJpN1P2aNU
DH9lmDea4Q5NHWS5jMj6K0uPbGD0JJFESvzg6MVagMSwJbJ73QCeMAuwsJaVhTy1
jK0UVoGLknypKORhVl+H+901Ur+yqISpr6rGdom23YfRbHIj62iQO62SOp3gsZMx
VBMxv0pbEUKhlEaNx22c8Wo9lQSrfocx5oWKAUFo/aFnjWbJgnmjxeZM5dXcCpP2
r80Z2UObSdo5NEF0zSN8jHomDxyli/TVcoULLx0kAQdnMF63y/DPZvtIcR9C4ymP
a+GVhwCq1FhxhbqqqSqzJcce963OeRUa65YFZQ0BoMhWvjNB/zTSYHpIA80yMUxW
ObHr/QrynfOBSug4AXL31mMzYIkqegoDXj0PhsHDKtFE7e3xo5ww8+1Zk3c2soZS
ppjHVuuBjqfttPY+Syi3FPlnWjOEqqaG/R/ZxZfiDvIJbqB/c7T6/hzNBbOPWJ4r
Ri/mN9J+Jyyme6AAuGa7ptuSPxAqwq0P1KMfrHBphFT6CWEoG6yf4i3kpx0y83yJ
+DpZXxv3SZjMbaw02Rf1D7f0MidtQrbVusQ+2+Q/qcURdW+fFE6PoTBHDvTztzH1
wlBm7+mls1lcnJOhxnMdKqhvKRGEi7nPQYPxwpt4ZVVZOkPCMf2sESWKaXuR+9DO
/bXNd0jTJ9L3Re2O62t1TCrSViACU5VBAK83LFwr6BoRw0okOPtSZU3AuwZcgwux
+C9dM5ZcV1F5++mZp6LHSe7NdhfX4Gw3iI7SUa+o6Wo6D5X4G7iRAKwyU+BM5F+e
y6jcL+3MXuVuzgwQV1yeDNlNcaPnqUwuXVszDHM1uDJL1PTj6+6uI2EyKIDBwLaP
OiBjV7qlZQPkL5wC3DYhh8riFAdpYv4/J0/twqDMjrEshgpboplfKrnmtMT91j45
vD4dPDD11+11aov9EzVh0ykJGgMZFOB7ReQBSFbiyxl+eQ9IriDPw6nZPbj0/2gH
sKYvC2NFZX1XiNwp/CYtdmuUrkO/ac+UeqQRqmp1+rxJ3Z+ZG50SzrP6mVKbi43H
i4kWG35FfxS1MRPdDOT5ct+uRlFYx4VreShd/d4JtFDDEmxYUt0QevmibAIwHT2x
4yCeQOD0/iUwvt99bvhe/lGraPykM6YTIsFmHGsjlGdxTb62lo7o/bvdfGsrJf3z
RszCmAbSspONeixpj6ZQUwNAPeCVbVGR4sQnnMnMYMK2toPzoJCwJALmKbB8oOLB
gR1J3myq5z7aagFIGcaAsyEL3lFCbj1v44x/vj5B2GEY2WyhvNdlMY718oty7aOO
uDHmGifwjJmdXg3Lc5ioNq4B898hpxrmkZ0xzNRKk0wC5TjM7odI0nAgNjFuMYZs
eQAWf8q2/7CRNQJBH3yibVIlGEUB/37xPUVpiIzBwK3zuVvXUzETeeJEkiC4/Bqu
EHXgcl5DPo+kA9p/yh85HNyzanvG6nMquezmXYGCvOUhShEbML9Cv5JNSsANZ8El
m10PrSUYpjRaQK2K6YFNJT+cjnfKKztXDT/71NbMvE+AjQuiVenVQLzR+IFVzred
k4jELG2TbQf3xCf/8Tyu77Q6grwoKZv+timF18POw0ZPripeN1ZLV7MQiEKmp/Qr
TCsUeuQxZurfvebqtJV9jHUwkitDNL/QLbLDQv+VSfjIoKtkA64hWJHP64TTbHgY
+dU7s3Cyuy+ydWLeSoJ81axFvUqu0ZenZsm8goOP6nDp04U4jwaVhzkjIk2/oqNK
7bsKBQi9811A23Z4t9ixIYJpGEIYTy092N1HfeLpTABBt+z9gR7Zxj7XRte0D4x4
lxfIGUrl6mJRIKCFNbWb3Zv/V1PVTUZLD0bpMvJtH17ZjaSjeZ4YO3NacG3UsI0H
6a97kduEoTxHU3+4jFIF0ymmqQsi4dN/OG+X+jbaNKXijMqpphQfkmhG1EeaYJ1Q
xkBdDtzw0Qhxs5UFpWkybrnYjBzyQWpYkoLtAY7snDo5Src86ss5/u5GZK48NKDD
yRtczhYrt3oRIiBpX++4nMlEkd5K4tDFfrjP7rNs9tjuaL163Z0Er2IJc3JBBHlD
1U3jHlejIarmleyYrPWUpJXK5/7KpGX/GpKajiMK2CNBs+vWJht+M7PlYUU0/7SV
ZrSmLRyO0GfojB2dbJn5uiceNCALzr5JFoBYKvlnp5BIgpPqTANNNr+ohR/HML5n
o075q+coryWVX/M8Vy4lTpTWc3Wa0e5oMyLuYrgupLRH4axBFnq0+kcrOqo+NSiZ
CFr4iWRrBFJGUzbBXHXujRdfNn2LPJcHK/QKQwfloS+1nybDrVJPOlqvJ1MGkG7i
dXLgtXZK3jBKGvX3as7CRcX0FYJOVTXHbqSu4ebgVaWGfbtScY1C//2oPlCZqfkQ
5hh/03n44Ssvp4z/eGvYUNs4BnL10672ZMThbk1mTCouO4geEhrXkWZEdUiOOVzA
i17jyk2u5knsClMW33fsH1TMmP4N0m38uurCF6RzyvDlZCUXUG4UrEVemhEjB2L8
1S5s8Tn3nSlLNaHVMxwgZqgZNYtDsOBeUzdiM20esecjN+OUYw7M8l5dfDzGm1Tp
ofB870G//n7pJnfUL0ch8URL8JUZVmpMjalxY8kWyzb1uuQVIXR43EV8rCUIaAlB
BkFRvs7doVFfMxiykc4Ad5F11MW1NDU3dLNKDgmg0sv06ut6ko243+9ROIaX7NHC
Yzy6RPfWqhaW1dbAOgWrIR2ghn1oqF61CWZV7nvhskzxdfwL92mI/CdauAJPvJrq
zgJ/OTHkh3lmdtrsHsynL9G0F4k7DLAqZWQfSkdgk9irp1XXHkOi4FA7/N+M3XeT
UFAh6kvCcy74XN7OZ1zt91ogF0v6h7vhQ0vSFsk+ckQO/VLemtbanQy2dp8d113I
l8a2bKCLculEMq+DChhddjr478MdpFPi+OnI9/2w2FGa+eceovyU9bayOFSIHRiW
4eEfFWl+Ur2iQnAKS/OaHUb+yDbBPqGZWJU5M+IYXP82l0JFdAHOvlECGjIFYtsX
tEk+K+06TMMZpg4PnhcrdX3dGc0vm3mXohI9kKSPO6VCFLA3l4CqmffGWhOKQRgG
PsHhgo/8kcqqk0Oaub5kAiQiNDscYmkMw7dV7Scs2WXe1Fmb44i0poAjwcTALG1L
oFzq8IbGCDvL4C4HHI0aqhwhHYmyeb4hmG79vklZ7ZLsLK10WYrL3cuN8uLaaNmW
ZKEIRL6BzMYku1seSncKfLnN4DULMzqzlSaHs+5VDMKw5ZNN5KUK1ngqrlWwwDpY
YDa+BRRcJ+V4DG4EJvVWIN/PDrKMvbMzSeK65mvQqK18629nz6VF0/N5geIUPvax
7X6Zh658cd9qihB5b6Z3W2fK81TAaffhD6un99HRy98jr3e8KdHVLux07eHRbjAV
gygBEPX456zrahht3y6ZS4XM9cLao7DhWHXNSyl7sUxK+R0+dNnV+Ie9z2R9kQKW
q4UQGFOAy2sPk9S21kqlNFe2bGEJkEtMA3EWnFFQPRB7IX5FDCFpQnLTweOGbbB9
xMSEsnoPz8QqzVSU8FYynbmM09Ff+Ew5bhVlhRJ1xFBKdjrwgCP4GMOVt+c14/Lt
EFAbyM8bLwVTziyyq/rqGr9y/IdCCrhUNZCb+xgET4NjJxHePAqK4+FoVlSUl94+
4bCjY+q2XRHV4lEMPpZFBraem36JFjjLt2+xjKG80i6mlBy3AQu2qLzaqdpo7Upz
pWT8UB8zaD6vbt9nR3luLvYwIBgwKrG01l3ScfYdrzK+/qLVneBgOwCGTcKHAGon
pa5UVIKq0F+tCEpIo/z2+PSU0adlY3QcPluFcMzjDgB+fOkvea9/XsTBgjwrcqqA
`protect END_PROTECTED
