`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYsaBLQ2GzUygUM+MkzAv6XuJuJ9kqmQzspp8w7mJtJUIoxUcTFtW1wLJ2N7SUJ3
CrLCK0wI7nNb16H6WJWrKLtuzBrd5PHopu+pOkHCBknAWPxZB2fFDLkEARe5K/hF
jNdtOjlKDvZTzfhl770w08EepDCBva1VmxE+2nqwQV3k1fZU7C98tcHJvphQ1Wgw
SFJGrc2Cmu8UBOpK5ShgO7zBEABPB5M7WSz6fNJIbWP8383WPJSK6X3ARvMP9vHe
rnGNoXTAPw+6UNDpwCr9m8s7pDsgFVJd5b3HvYJHdYY//waQ83N+yjVttJfENaL1
Um8P9xnZtXX6T2ZV6OVUq6XiZjbKsRiGNgf0jdV/vK7lCxmqB0PDMKyv43cAgERV
b6OceQ6QxYxhhrG+IaSJzIoRdk1izdyLyr3/mzga+2sc2GgDTdB+xFzUXqt7LHQL
FJYeq6VyIflBguXVoiWVPg==
`protect END_PROTECTED
