`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwuPX9XS4Hv+ooAcvt6jeE3AhB4UPNMDSbB4slQc49ASrMZ/bRm4anhcG8yfeQF/
Yi4tZJMna0/qwjO0aW/kAVIDWKjKV+gLX7bJ3F6DRokyrOb7zuiN0G6EMKvgeUUF
sd8h/ca0l5+Lm9kgpB+7egOWTvr9ux2rgLu2ggISbrlrOtpVtVTpQ+JNkwPvotL0
96QmKqxIaa2HOGR8LrRQPr+gtSyN0hgSOqFSIbJktM/bsrK4O9kKRwoJZ7hZwCkK
jolBXfDxZB30JZMMoiKcC6GoUshp53BEG5aowDx7hHOynK5vPer4L2GeM16v8a59
uUzUtCHzjORz9ZBQXMi4IpG6eAnLh5CqiClKVYAHH1pkb/HUA07oFFBUijhMlACP
gcQRR/YyweoRO357swT830tRZBzItVa9a+E7T1GW5V5LSe5uRZNqcciFDmBImtf2
lWzHf+odzsxkQM5X6fRN+YXn47QeOo/NQi1OpJc9lVHeTKu9LJwmbCc7MluFH34F
olKjkN1BotZ/Fg9uKXOugAPHbTC5tvoYPqq0S4V5GgG5vGXygL6VhMdtw2hvQID/
l/9PDpTa1v3pbpe+X2Ac685pDeSzXLfpMw3vB3/IKZBBAcP4bTNRdGzdrZeNadCg
tF5onZTyZ5DS3FSQR0eNBcDwa/0z+wkPb9ylKNo/qb4MeD7jOAkPKBR11Wr2vixE
rSSP2heeubqnl24+LeYeP1j3xd7t/e0/x3BVCEf0upJphqdUrW6Uf2TBrwCZpkos
YhJ0NlZ+1wW4sqYDofUPoYsOdT4MSnRhoAoeBdGU5yvsF3gmlnflC1XUIrD2IFXA
MOh1U7EHhP3/4xsqiT5DytgeVqTyBpJONB/blEHt88ByPzSpmJTAtWr6jE/8PH9J
cHXVGlpJ6whVse2k2TM9ie7OLWmuBpLReWWxaPUgszmayzqvkf2tg/WF/HX5AIMX
CjKAKJPn4dIQfr0ryLXutV0BnQuHRL4+CNMsGlLQNZVB7xf6GvzFw+puIPYiovYM
ctQNSq/98nh8UyzWu7rlGgvtZxAnu7ImN/L2HQQxpMSTXd4EH5zalVvcnD75EPhy
hLWrKJSqcbd0qlrTjh+JDL2FeJH31PUjA7y4vbR5uZ4AVXBcMPoInBjoho5UtSnF
c5I7pIxk1b06PylF5eBSBenV17zmS4oQXKQPC3fbGw39xZu6gQiIdc5km0MYP8uv
nIBB4nQh3Hix94ELD6YViOhtWBX+xrJruOVR2nhn/HVUnukWYYufflWUnmK2bzU9
ABNNwYz1DYPzfmJVljS6bEffZ5HQFiSn7IGmWPKELfH487YF2Sf6rFwudBcPvQHF
mCyIxKmReV1P2bvWlsH6uO4iAzelvUmmvWjnB4wcdGg=
`protect END_PROTECTED
