`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X31oDYNByiEi30rnkyCPNpjrHXjI+G18d5C91693p02Bv3GgcfD+FDSXx0QJupXc
AM/pcP9VNbG424mwyCsiPLnDJ+mWSKczKJyfatESmy8In+s5VxlPgNM8HHZtKoBo
6qI6dQHm4ovheTxd6udZCXy6DJiLrqe9uTI1/L7/qSs6S8g98sYD5ajU/VO4w4ia
4AuNi/m1xw5SwZ6yZex2xwaKf28z5dYTVG97AhST2/dmEDUcYNKzYmcGF1X939OW
+URFTmRkwZI/SffPS/hGr40qG9FCBCpAIb3MfwFJ3zHsEh7K3tR2fW5Qh7+EJon7
OqGddUttiXf1OTlJ8Wp4z1qeU0FX2xb1E5yGKfNCe6Vi5+v8axG912/k+hFgtSCM
HWO6/lxiEXnMsb+nLNJHnkGSGFqo7jpPC3iOo+Tx0iGahmYihhFGa7hX158eC6zc
Acf9j7ShO50NtHwUnfE47QtwZ003zFg81UH9cMDWEWPl8YzM5jFrRolbFb5zixU0
fFq10jDeFXYBiV2J0DPc0qGZQDvBxJTWTFpNGrisDWEM/SKKi/JyO/7chutVHyZG
OHXEbzS4xBEGPWuVipbEV6LV8iq5kB/hJtvAD8P4zUUOZ26YqXsbuFx+jrfOBmAa
oawpUfPVPlf1mIlIm3r2iMGnqsXphyrCLu9mrWhq7R0OY9Oacs28qJqZvsZ0rPrM
+8wd0Xge8foULbFWUfATnBuWiRkHtW/4M7w9dwM6/US/Sg70GiRvd8yjSRvJ2oil
XI1crGEPQobagFANYDwX9GgfRxKF9wqKbnpDhadZOMepjuY9XHL20EktusPLO/sL
m7SFmPOjJx3SSKhJugcYV66RgamgMWHALxXVY/uCyVN9RxlenHNXJ1z0tJk0h6tV
0rfP/sgMnodgfOYgWi/1qwZH5IGdS6Rp6W8h5UcE/dum7zjgiN+QTMZ7dL+wJhn6
xF+NQ9GpWMUGBQNZau4/m0bs8G2EMuu92SIm9NTdiaelrxToDgqLEBOPBdTEgOt/
zVxe/Kur3QGS9ZRUY30dzh8z4MmEPYWIfnHgXizWpmTfOp1HOWd2AI7Nd00r+9Jx
ANM0Rax1fo6PDvGxsS/Ry9ia5dgAL4NU6qqGgfKRW3rktIYqPHcCFDVpOP9TnWif
kAv6V6a23ZT+v52Mv/LEI/RNSmT5P6K0N7ZZ9BQbin8ihuAK/VilFk1/6/LE8wda
DLS1JT+6gr9iIwXwOcWyVsAFdD9V9lesCIZ9tPbuwUP1DeV7GTwp4N+uLtGKt4W4
jKuAq6Aj7Nkjk7pGDRyDtG02pwfTaqRzMHFQ8CdEiHKHfzHNYuj3ulLaf26hcfC6
/GcX89JVKab5bLxgv12paO1PTT8H5S8y+o/J6hmwnDXPvE4yFzqrY22lsQbppybt
eCfqwHxqoE3kULRQiAB/sE1vNB2UlV7ar0ZT6l/DiGYEiwBQqabGweMYXqbcWz7i
Utc/tPRU+1V8EUFkwcjFn1e5HJGJpLd9DCa4hGBYz+50vQYfpnymLO3m0SMwKaBz
t5An6nzcNNnY0b57PuD/aijE3hALktWNI8WX+yg+6dHzhZfAAGUO3aep/ySngUzJ
afsstd+12ifDzl0OnBCjaLcAG0W7NJW6VWGiSKPZwfudZpgKtaAtDFCKf9gmXRa1
kybht+3AKlXkk2y/lG687Nhkf8deqXSV6Di2K5qx04E0yXnC+LlugBz7MRq/2Fh7
w5tlDBpWMQBBTqXqk2SkYe7HhHPaMgbHTJfHjwEg7tgXgdpMC8A59damFQtlZJ24
TNi26j5OkQXRFj6oUbeCbYPUi/aGGGC9ItDDODUxS+zf1LKL2ed6yoA6i2SXTYWT
2P7BmZcbWRCaPlAONJlcAP3cNcYnnqYQvXqneHgFrWDvuDsMKjST5syOpp1fSC3N
VjfNTMU9brUVQ3+9Ep4xMCeHcgWwrWPAiK4RXTQNIhkWNLk+GLX9xXRgCo8sQ0Y+
y/EfHOWGL00xg2aq9e0swqUWKolvUk/4v0+LWQtRi6u+9iQP86zg9MgaRW1kGCmi
chGnDfDDGTWOKYPItEmy/dVccapttk+svyc2WFLiS3vZVi75J+7ISCudd4mqZnBw
V+3t+JBJsyknWG1dxhS+CtJNLLcMMubI3cSTCRBETUm2ouCbg8GZAkmRC8cDhltL
e6iOSjyT7HVJSIlv6jXjefWy4V+oG+aJ60mywB0U63sDTuHnd6dOdCIHK8OOIjwK
cO5qQg7nNd6mJfuDhw62Ji41kXChr1sHk0De0fabUww3kyPCaIdfcGtpOlWgsSbf
iFO85mvpxA0mDZeR+NWuDlOv7xC3sXZ7fxc5qWC6YfgyprKSOzD5a0spnIzEoGUi
YLHWtVlYTpP+iBqWZsU5ZEQDLXXfHAVJsagC5nNvqfEvPHiCvhJmNvMvZHWi2RKw
6XFYZlH7fTiZi33mzLt6x4yVqnD3sP10V5vhkxBVGZDFAyIoEXQRFUZAHfXdEkmg
hrks3iIVwXAZxvcpEo3UhRoP+a/gXQev5ri1a/JlVse/fQBMhCuTQjfweLk0DacG
VFoaVGA2ihQSFRTqfrpzBrV2YPRIxDO/Mb4SmIaO+JxX1njErFrHsnqsileYoX/Y
EacQcsyovVmr107CvSd/30gEiz2/nIiZRzo611rEpTKCkAy3AgaSqWJfhwaWDc61
vSv6iiQ2SLfNu1hairv3GQprD5SZLkJWFkv7HztoglomjtJ3jmuJIfKBslDRyaXA
XYjErjx1hcSEKW1oJHJof0oE1nLxFxqHHm4AslvNSyTlbnRTTjVFzcMyKEdjwufE
dmUFuK//UQNsbGeRvzjfOdF8peAKQMEJJr2is0oaKenUP1tpAWIEw4CygT+B5smy
4p0N1lh6XSnB9gBR0+RYRFIdC0oPkFGu8YcAUBasHrNwp1Pmsq+b2WONpP+FR7IS
f/5Z+iVQwLfXk5tZelJqxE59IboJVZLylOIL1NnouSdx/qIdvBXbEuFDo7khm5/E
zrmSIBzgpReoAHAR7+njRdSCdBt9QWTQRo98K8wKTYuTv1HeO7JC+WyqWUgMVGFK
x2MWz4B60yoTy8EaNdQdHySzzDro9rk28rcz2jmCD6JtZOgzIX1YJ54CayFmJUfp
KyXWwpdZAhx1EjvLAMxmzHsxiuJqN+UHYAyzasmC2B+LV5GvUiEjMo0WKZ62pccp
lHxVQGp593bB0irqXI+LXL/V1Ml8DzJi/nNWNEIjPrxAH/RM43X1vKeeAiWyJR8+
z6r9ltMDXnRJ1S/XazK9rrGJi85CVs/jVoAqScPMLYvjBA72a4xzo7cQhaWvXcDK
1u4lFxBg4sdAdwirH8baSzl0BRgYZC/WQXtjRORrKHpeEVgG46jvk0om0CbP73PE
yqtZBtI0mfhYjw/DYKixyuyEtSpafeN6IwzPs8FanpDlGRK2eSqblCSXIr0oZs7G
u8sBjzkHPQTk16/HyNdx49EardlYOGbKz9ln1DelZ18aC2eqBUpm/Gpx++XHoxTL
9iJyB6OoGeytLfHHq+s1R4gFl0JoyKVffa8DA5QH/ntkLSou7e7YBQwwHVIDDLU9
x7ICmNJgStj/1zVGx8U9EXbSr1fgA7ldkrvSAfjx9yXT97333rmC5y6/GiOlx8Ej
O7iJ5sAn3JVaAOfPtDoVT+aGCh+EuTgNpvqcInnWdrbvJD8+FAvNPRGtQT8tFPTk
AibbprTXJb36f4IoakuD9fwnH7Bi424i+cvdw3T70j24k+1J1FIYZPI4QqogoczN
Ym+yGprn4rL5AN2wAR4/VA==
`protect END_PROTECTED
