`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nwttGNCOB5XbgL9hhaLmE5suuXvkSI1crl/aUPI7sUxbFUAKVsbVFlNm2xOZ2aOm
1K+HcvdPT39Hf6dCCqYat6uyVbjeWj7i7zWSI/XRrDAETC7Go5gB1l0IrEc6DpK9
L8CkER80Zdm8b+xy1sW83zbGZJtODZafK+fwCI0sX3x9RKkqXrJ8siWdCJOkWnhf
JLrURKXp7Q59944BzJM32bIXluz33KKWCuCV7hOvDO1hKmh7txVDXFmjflZqbwT0
7TNmOX7x5xihYRsN4HoWixlQMRiRMk9KMsrJ+qhZkg6mLeDmq9RdVXLvUX7+GaKW
JUb5/JpzyENgmHOQ496i00jOaeQAHaFLu4iqp+l5vU4okscUxqDarYvzQSMC8kl5
BmExw96/q3MdRKRSxVAEj9eeg0dqQfJHnG187mLZZheK+igNHSS+tcxt55C8YGng
q0Uv35/MGegexf70wUM+fbdSwalM7UAVw762qoVkaHw=
`protect END_PROTECTED
