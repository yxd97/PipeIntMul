`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twahJUO6FffXbiruX3oUki+Truhbp3u4OhEsSmwkAt7nfGluLLLUROayE3HNfzQ/
MFOg5Frk0hhtjRZG6AtUoyB9gJTm4xTwdLvIM5syQ6T8u7Lo8KQ8rpn/+Co2KFjp
ZRYu1fGCvce56+w5pDPvMa2NG7dl1tdD8fsQhlDS+HMT+cL63IBtiIQvzXn/jbAZ
rb4sBDfmoGYri6Lawl3zufh536+yUdT/T8FBoP5KUBttTKPwWJksdfoJM3KyH9xh
1EC2jviLriCb4/NBLIZoQlZ+HoWwfsqFwJiGREGDnOMpccKVkZyOjMT7D1N1cRLs
Nw20JOLH19xVWEeTOxggpcl2+/78hKNP4YI5KgjL4TnOdaVbBxlbHJxWCUHBPnOT
fJvTabI1pZoU9Qhsa1ZlMkDTGIlukbqDhzFAI8tFTyc2fdcc4ZblbCjYUxKlxReJ
h7oQ/qJLrph8eix70JuCftIx7p4oARIA2khTxRUU1Pz/ht+y8MbBJTnDNmKYSa/R
SqDO0YhwpVOl8zU9yUU+rNl+Rv7uccw/B/TD0M+ThE9FoojqPLCGq4Vrc613fGtm
AWblNMrzenAMTdXVlSOXAYvV4nfyxd0ROS0NOWC+/4FJlbjdPjZ/ttO7Tw9TtW0V
Lcg1akPvLXi8l+czkIFklIvYtmAadWaNaJJNw7IvgHNjseXe60RZKFSYk13qSwkl
JJ+hlfSs8HTZbO7ZFVsTL0a4QQSBR4bbmfmfosk88Odhw/dnqF8f/+nbIXy62ubp
2MZ0OLJN8rjyODNz0lASf6J5Jx66al8rkh0vSSEFubrZnENLsBhWOpVIifZN6TWf
q92mHisFjE1Hi4Lh6JujUJ6Hf/m3iYTNl+m5FjNem/d4GE7xrCITFieVzcqyzrWN
b0TnzR90eJHJrju+D4JsdTh93xETiQCf2aDey9OeHqzJoZVfdEhJQjLT0I68SRJR
LHTMdnBdwy1GS506f9+3CQ==
`protect END_PROTECTED
