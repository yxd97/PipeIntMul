`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vvfoFG/rOK1Q6F/NReWNrvZSvYorOUEEszXUoWH6njy38bn/3/uaaEd1qRzYjnjm
GjeWP6eEQxTudQS8wVM7CWECUAA4xnE6FaSEProAODyCXozaeQtyFImcmbMiFbfd
MPSVTGiuicJDMJI5dZPatCz9qrkTtgWnspEwKTgXAjN55eKinuNPiYUkDRZJtRby
23GN4S61cZXkJ6/++xsl85Rqba8QrVVRSghp3Jq3ULCFDtIIvFfF/yNdZH5YTlX+
+1VRE6qGTXb65DCvY8/K9fnamOVFe/i3WMkfjfOdPET9+mtkq/UBiCRd4xHJ7gNS
`protect END_PROTECTED
