`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEM8CFCxbtQJwEjFeICFzaQILZziNzInpPPJXUPYdMj8vr7GNvOLPiB8KY+k9LCO
Uvj9wiCyFdc1RLHW4cZXuvPOnWasWJUWPKkyuM4fjjENymDgeUT8uq5kufzmYXCn
6RhIWAY0sAZ9KMag+Y4VHBIgKjmLP3hwQlDBgTPTMOPMI+MHjdWtbPf7WblvLOaO
9fQCu+colxqI18+kyZ7A7Mf4Pwgo4SEUysrUGl1oXl1H9AZ+xsnzSu2DwUtUPtL+
RfKLX8E7vWzFLkEM6CD1CMZwelVAeqegNx4t2Q681jY2k3sOR6gUkMaBmrskRTRl
DEXcaJyfsYKu8j7sXaDvpbV4pGnTYNoy+OuiYSIUVq4nvk74VTuRaFWSmnYse8Uq
ENG0vYY+R4u9oR7vroTPwtEFaGbMqZ4cNtZqddUVAIq0f9/vQBnaxQVcXu5hQmUh
z9eBeRe1MuDG0SwzTDINa3ZKZoovE6egmzJ+ogXx22ki+iu5Cig51rHfgB2P4FSk
fsrezmBQlEnfLJyK76HhzmGlY9oAriuiXzz+HLuJtlHzfFNY7qZdEiX6PbUuRAeZ
/98hTfupcay+fjYU+a/ek+6pafxKlY72ghLGs4K59B6xdvrlTFU+RTcFREEZTr/S
rbxTxKH8VQ8Xe2AO+Gr321RfeR3MemMv9iAaTFsqFzdLmAlWf8XlVU2dswRRcido
jq68vXfOiWXhQBsGeJnprlt9rayj5AbPrxht4xT+MRIxG+j26jviZNZPsSf8DpMG
a3jO1gGOs9o+/BwXLPCrmkt2ysEGIniG3a+AxU0mIWTc/NtLZ6KbQcs06vaVs0mL
G+h74WzckeMLzpnga81+DBNDlUa0JTP9/+o+D2INpAYU0OmS+U1yyvgA/+WfzfZ9
Gp9OICyBd5oDCQ1J8Gz9ujcUG3WSohj5TC553bmDluzUbM5XuLpnbaXY5dnaG7fu
v/jEgOulBK8bYUCNtLJ2HBvGXF0Dia7L8jHL2wmpcYR1kKirKGW5M8qySVfelwq5
v5ZuXLxAJb4Rwz9D95MnXYLmcuymTYY/SgoP5NK5ldhZWieOdmgHmZOkh0WBmldH
EOJIcqFxbU6Z9L1PMHvWITAuEL8M8SYVWJ59kOtwzYaKWjwLhMA5CKPkWpdTUaK2
hKRGrfhTk3lWx9pbdqEjqJC+JZ+WmkoKp7wxX0zgNp6arMHHAtZeJcr68c3Lrjl+
OlvJEtkhmummw8PXirlwPWK3OYacVkYctlGPzERSusJ6k38ohNC4FgSY0i9t1ABU
/tQjB7bLt+Tdbgf5OjB3vo2A00RWynDgOTI+7TDQngPjb6OvDo0qhgNkJ0bsTunv
1UWHHU1g+r8PdK7nks9aOCAKX+0pi8i7ATSbYYJuHsX0uGvu30vIHfMwR+Fqd7nJ
AqDgOUeaFgZt1p6x6xyr0DqwEtkyqIWiERW2N/w+g8ylhgP4VwUtEI4ePUv3FVOf
iCwmTv9WOALpz5PSijYumWOmaKtd+oq4VRzyK0F+JTqcKxgrWlktcan+exhScE9L
MGxWmyms26VBpnTm+TIimyJyScgWxwNUrRD55fjw1nqsw6h5Vg9EUGCEsQXmka1X
91lxIfMLaxb+gPOPfsg6WqmYn9GErUE/KuDMB4qGw3iNG6BxIjTqPxtPfGjI2inp
iB96vGxiikXOZBACyTxQSK1XVuUGC3DIToPIRinJeuo4BRzLI46kGA+pYVAUkoAY
QZylAU9Ppx/9+WvoKX5BxvZN1E379w/xzlGzNWz6Zxl6xkCLYP5MJSCwMBw61CVF
aCt3qtRx/2pP2FruJZoGSDPNNE3rYg8ZbOu2EX4mc0uNZRtPYZQF7Ct+9P1GZm+X
ZXepvdP5a9MVQa+hxcXc1OWXZJqYckp1S8X6SpyLR7N3Flc0swy+Xdc9pOdlC8lM
tlQBGffuolzt9Fn91tfVgr6dq+hR1YEoezR4LytHdAIPHbBaemwRUE0KhOXdG9Vj
rOFNhxx9u8HtRhefHESTykG9kvy9LR0ybg9kOI2M5rBVgzNNcP8hvNU3Sd8Tn6J9
sPnoUm72bZVsukKHJVjMjJSF/pSPTezv5+5xwODcwueG3n0x5fLKQlykfeZXg2dE
h/xP9FFtYpKVsGJK6Frk6yms4zW/O0UjfgkqRpTR138sLRiNkfByNPPD2CyQKauT
vYaS1eMwjCSGhppf0dpPXLBxdKQvmgZ9pyCt7l2PS+kgtKJ1kruoZFSYNLlKiWVP
ZIMX7Fw1ux2giQWXSU3fg+FvjWsTjb6k5F/7NlyLuLEyMjEJvzyXk0p/aOcmVVcD
v7mjUsD+0ZPRCEbAO24qvCF6iP2CIg/LzBj3ou+l0ExZivqGfidtDQ2kOTcagnE7
P2JKzNDvKnzxwG2aEP48NR4yQGDSXo2oz/JxT3YMXeNRXJWj+6UHw3VaF2T6vnlp
dMXp+ByfqsJU97QYHCbJu2KjSHbFyj5viMqTUrB4nw5gnT0zfAJiOvBTkvmtaO1u
917ob9n3lJT+zZ9tT4wPCBjaWwZ2ibpvLBaT64Pa1tVRFM373ezbtDFVrAvitpf8
8NMQYVVYF1lnHeOjh92Nccj0jKShC622GkajQ/yUL8rQ8Jby/okrMxnjdmSQfNXy
Z6ZqK/QxsKNtnY2tdx/1zTTO32GcBHn28mj/YEcIRoYvHo7wFZV2CAx7qNGFquol
wSDssQEaAsK6jIIFmzX78TYv/efuSlX6QZFNmiCi82552/SDCf0W1bwdMlM/mbZY
uDrgzLTovzdugJGelPPVDGLIHOcPVI7J06oyOAoGuu541ijjfDW6clxkxcM30yHo
FwmYupiFxYk8Ldl7f8eKjKsVTRnTFTwcgWnT5clTjcy3r385j/g1oN4S6XcHTv/Y
39K8ilzwf2VDkw2SaJeVSSqiQoYB3FWhKr0KC8+N/t8DwyJ4YivLOvDE9dlx4snW
/jjmdk12LG8HNMsDCSCOFydDY8TVH8YRzQifGQowGa4ZdUQ/8qbWMZkPBikZx2UF
UgzZmA0FZjOhGrxphcUKgjT7/k+gzcz979w+5A29TPAiw002TtI15qlC2ORY7b8E
0adb+tk6kv760cuEwEePHXsNLXssn/lyIvRYzIkkG9J9PFWgTH3A9NEF1rSKc6Uc
ibzDlLnbseG19ndYhTOu5OU57tsqjVLIMC2GSg1VEvpBNPS49hXoDeIDCygKi5tt
Z3ecig4yShKqTwWvm8vVHWShbqT9dPjyiE9+45Dk6sI+QI7hUIvmi770oxpVBc8B
jHkvPpvHwiK0x/cWtIsxmj+voT5ByFF6rbsVIRcxPUgmowwAMraqfwUBXS2QaLjQ
2F9AJjhciasv6EjAHRHgsw0JH7QZ0w+3PXeAdvHY5GP0h1Ms004Nwk2NKKqabDFJ
dRKURPiuyAR06kevTQtQMDpoE9AlzXiAgP4iBiJjM+ZpUfKHfjW93KnzoAG6lu6h
PUeiZv8KI74nGW9xSe0FNvOeuqQC04+uA+eJNtriPZCriPymeGPqVw2wsTMGsniP
C8hlVZyivn8L3WxyclA/lDLB44/qWad5VUHhwt50hCyo3tbNiJFsJaoNS8a0Jzn5
AsRnYN3CaAMZt/9cS4rt6lHOPoSldgINZRKSG5KbKHxFtcmcVeczkR0BkasxNDr4
kGGM7GR89z+MAVWGvqWnr1qBaTcjfWIiWgyu1gzZTTmw4FvA8bchemMa5cqL0bSv
9dORLmRyBbrHVoaUzVqlpgdiBhUw+sYqWwIuhLaAPr7Bi/8lcKrnQYuulcWfdwrP
iQdZnbro5n2ZXwwKQ9GSyQ5gMs2Nac/vwwi1+4VzQxPvwFOuqQd9bvIMu70HClrp
LqBv8xqzqZ1KnZIRkFTOt7OVM96X0Rt6PkR6bINwLwqe+cJq20oXdcsUd6pZcxra
h6qB7xhe7YUUC0nojCHOwBMQi/0fpnzs05XKl0r9GUZzO7kKulZTTVp5gW/67nf8
+SwA1NsZYNyVPkt/qh1Xk8X2lCkB5ksLB7Ug6CBHJQU=
`protect END_PROTECTED
