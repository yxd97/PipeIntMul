`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
13Jzz/lGM2ForSYq+iUasptV2+F+2bFkfDZ5ExRy8DAyHAMAJWx7qV66LZ8QSDak
y2D3MQd/PxNIISF3zcFj/0Zm1xIj8bSpbw7QHwmvUQ6yCfazIvb2RP8zBsS4+3Ts
7LnF/JXePYCelaajCyju7Qqh7va4KbQLSWMhpU8SL2d8b3ilu5M3MfzWcHmI/gdi
xkw5xUTWFU/WDVDp/DN4oIu84ixw3yfqMjjE2nC1sJYP+VpQvI8jgle3DgcGlqOH
dgqs/gPpUs+5jOpYyxtez1hbiUTeWeA8eUxOVZMdPbdPcBSV9NWVygWol5gzlxYX
zEwIoP2KZ5rHaFodAOCEm2mRSSxHZuEIL43mK8lON0MeaIW1vn4qBIHyqSan3iCH
fUmubwhIbTia6CMS5Zl+qhKFIf0hdpyc+zQLA1XrwtQ=
`protect END_PROTECTED
