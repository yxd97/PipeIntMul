`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
677Of91mAGrZUisX6T2JNajAdG+TLdcogJ3uGOzDtbav1Dacz6NjRpWsZvYWDi3F
pRIYwllaml2vmtq/m/s2Fw7sBQXcBp27q1T8L/7N2qonIkgkOUpzrS9XWNx5fRtA
sImp4a1vYJV+zB09JJfKw34KqPXLetxMsSQ5uS3SVffQoHYS75G7Oj0UhigleS+Q
v2+0OVbZxIpssIJOE50uWP0L9hW4IoCiGG6/Cw1gvi8HQTuR2q2XeP9gC5dxLjHs
ywDi5iqMVKy3DkYooGerBfzwOhBD2lF4zYbbWCDYBSQRzncTIX99gFAtH3m1pg88
NyPEJ44/XfL8V5nUQKg9sW1GksESzqGFr0yBbrPUDy6hQSpUnWZK38JYci09wAsW
BkDsxUJW3TPuddeKuhttp6+cwmyxShDbU1QyL1D0s+k=
`protect END_PROTECTED
