`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUX1RTSr2D3nzlwgf0+jqmTG+jYJPM0Sp6xGYkze7nl3xwcA03fgznAvNxO2AOMc
PWNq2nTekP6cemSSABwK78sN1gEEqImoeK8oSKzm9R9XxBEblM1UBLznmKGbzLKf
ZQNAy4Yebh51umrRngHgccLkXsoWA3VrWHB4GldDo25CvtMraX1P7P0oG71OJr3v
KlTB//naZcdwQZ0UKmK2x5ERXusJNMA1zxtWO+rIMZKIE3sB/0tpoMrc65yo+PI8
v17F18GZ25GR8/oR0R1bomTcPOcmSgPa14+1eszRusj9/mSDJiVAuGzZf2qzCGt0
sWOQglW+2GmljHnFNMluNYiN+DN7kLekyrtLmIU5mtcInlE26MzActSIq6kU0hTK
kEep/lqNXQbhZuG5SxV/gi3w03HnU04KigGGjyjbA1jYxYeEPHw2xLq6lL6yvnPm
1HUEPwykaOUjwjzTEhxvI+mDJKZmfYugWsp2pT3x2Fh8pm9f3rcv8FTSQ5mJFAee
8bEa4IAYwBoliwtd4/MEL4eZMbFb0YEBdWc+F2X67TLg9BCopynbtegjFOD12Y92
l/h4uLK6DukF38MeJcaUPUUAVRdVYZSIJPvEDhcd1QTB+gxpS1qyq+wzO37FEc8s
lRf21Z7nMtzMtVvCrwWnD+RACPPzezbHJ+GmnW/a+fLegUeFoTrktpL7IeURqzU2
zV2PgdHjzTd0aD61dRzGMLGskKc5E3TaozpbZppxXkCN+5EHGH53TJxosj6l5psq
lDATgpZI5zLYjyhnwjJh2Cce1BTFyna4NQOXftU8IZbD3i3j8tBhgzua6A7VJcvk
kITJk9fOAnFVrLX6vP9h6h/HPyhtZ/B5KB/M6tH5VfrARj50C5JRFoK06FnjQNPS
SCoHtlZTT4QBtcwn0iJapCLx9ZNWhVBmD8ut5+ASwkPJ1bKIFpJwbNvmvFQpN+Ye
8ZuBF2/MnvkTyTzbPAsdjcH/AuDbQxIedUYcCdKKzVAfa/fYbcoTOgRlai2Jj06W
EK4b9oAJ3MNsXDap3A8G4Jdi5fD1T1OMqav8AOBjSvuavPQePFp8Rm3YiJIYGIoN
c9Pn7+xE+TwVbdMjsHz356r+ZE//NPhi2ApdjYh2On3b3yNg+Lb+uwXvQL7ZJO5d
VJ5yBDyNP7VKXjMUCbDCZSdxnwbInEb7xlkuLwwsXMwEDJhIwkX77tVDw6vnxWhx
g6uKbtCcCtB3ezJ21pVYAgB7PBk7k+RTobbC91jvaoJmMvZd8bJtFDbaYNde4DBo
kLko/sPLLFNQbJwf6zq/AjsxlXGa66+H2mZwYc5n75MywmpqZjaC5KhpztsTJykj
uMtPwOQw77M/DXJlcudBbe8fEX8M2iimtbFU6dFgKn23aDeexYh5al5H8JPpXXgp
mJbDBjhvyArQ+qgHXuTmh5qqbP1bXicuZt7nIC6TQNBv7qvu45jJbT/+zdopeNzS
i9G/19RuaRT0UM8rQoXDzSlTWmDbf96tdMpjjvubPMnH0x0ysEDVo+y217XjnVZH
qV7WmGBqoWNlqKKfZrGTpFxpMFeYKvedc/P0QvnzGN5FjIG0pweXffZSPh/GExhT
iRwV8ObkLKXNvH+Qbd9vfLa05kQNY7KjWz4U10HkGVrl9qwfEyIVRF/dpZvVFHoo
TCbePRNg6JHLAUYPMpouDwyZQOLEslpuTJnldw3LpiTVm566E7ccfjphovw9xvP1
XRGNuol6bsCANBg4X0JvlDyQoN6KGKKTHC/qCw8CW+xwHCL5wkCW4PDwHUDi4tiA
4gUv2Ln1KeEhJCR+h2Ptyc5BwGLSYIGGU0LwGxZaJS+2G/1SoFNP0bUJS3iCMGbU
JLojXWH7OVanMasN6igE8U2Txx0kQesBE4rzhXpDyhcVo2s4KmC6T4plcThhpoxw
JtGFxCRO0c4JsX0RiXg5rbuNgaM3VR+27YBmZ0DXuEygGLBBSRlfR7g0Ulg0pOZl
vG7CoQ4MllyS/y2wJX6V0vtf6KBimjAuy1GUS/WL22mI2zuOB5GZR7Ut9ylBCj8D
nARlJ/QDBXmpUP4ItFoqxZ873iZP4lHLJ4Q3/a6RdJ9l+YHRd8LulCYwMYLrBL+I
tdZyr4/5VtQ5LPfOwBmh9eFujFEwaUi6IEQ/SZxsCCh9EhLUMLu3mfBbdFLuXnQj
1ZSOF9ngc0I1kluVKht1RUfUMxMKn2pg7p4yuiCttA4rEoiImMGp2eJ8u0b3sD93
G7gx67z3VDFeI3ExmohEaJ+JXJNJE4xADICWkCBRTZCfs6dMws3lDLkAw/0aNUKu
sumL7S2FQcOR9ilfj3y8LSX7jTcfXPM/73P5nKgl7FKsQT656+jFn5QZMQ8BD4s7
lx0OA4OdjJxvw9vgQnbjBr2WPgJsaUQ2oSJqGnurqPepMpavpiHrYCXvFgbENG9w
NUakpOf/pbFLQcq6aoK0Jv2PgW3fTZxSSiqm78KIvJo1DGxCpUxaNgbo3I90zXLh
2aqEoMwoIVFB8q1YVhajiYxI2ZbXU3Sv6Q7aPTeLlzQbKRSNioEKqaR0AAy6anL/
PZkVybMsc0DpOIuVx0lRACdkclK1pMbrRwRXgGblQ0espvvLJz0K4VBT3IqkLa3o
78zJx+amEKrQUduwHmBSaR4KMiU8oj/ZEtYH/DJF2MghdKS/QfxpPPEAl7ZnqfnT
SROw/HVQ5vC/bH3uU5TTF+NFcloSx7n1ugY5+KoCqs0snB2DiHTO+j4Spk/7Q3U5
tbcI1uj5+g0v+6XJPXb/Y5mx/ZPwUOSmyZsWWIaMGB98vG329NKgA5n0iTMqkLH5
QuULNWIP3k0WrUymAHSIwmTeqIrQSG1x87lSnjQ5i3d0QN1wLaMRR7JAc32kT6S8
yNg4/1L4LNibmAAz6rDZzMRr9n+KRnBVbhmEsapuoUu7ka4eDhHoQu2WeCAGkVZ2
dV/b/syC1lsmgbiqWIR0+eqp3cQrCNnAGqcsTp1qoxfynLEUDBofE6rYNYKFMT00
tVe44DyKg0uLdM1x4pING7GzcvidSjAgi4cGKTeGWUcZCwyVRUHE+8e/D2xLbdhH
0gByAuovJ4TAVtWOSjNf+E9AojjBDCn7eBoBcRPPcRmi4b+rCRnux6KkovYYR/T/
ZTIlKhhC+8uRvcsipmSYG9S0NREiDbZRJaLYtP686oflo+KO+oiwYtkgJxY4U0QB
Wzi7SmZD3+dz4T4tS1VSyr8YX8D+212EFJ9P9YSXtNzo/mNaPGMlWuUEGeOd9oT5
YxE9Tg1Y6SWu0xDL0mhJleFIZTUXByd3RUMJfrlWmM+u1ENzJ55qqSPWpdS9lO2e
AkG9oD+E769Xlfu4edr5N8yjUepOVrkgfdrkv9JzxrVSovfvgHwu9a4rTJXVbhR6
LlMXep3SVbcMEk1/ghMT0AiIeT9rW3ZZUY/5EpPHSowCpt4ZA6HJjJpW3M++5xGL
jvxAcHpq70ROGP7wWEks3DC+deqv3xxDqxHpOgFDR9RG5qqs3HMkhBgAltM/9AEP
ep3KJ7YyYPleZNoj2og+JhvmCEGXMv0CMCYS34Q2EniSYdQgbe+bcDDgfdlXTFI3
uWAk4sPTAB+WvuSUek03KN60AbO6FMRB9HhSN9RQmGbBcwLOVA1PaOkWh+3KUr19
g7mTPkDd04vAbHdYI/b9fX2B50f4r+iBDpqabunDi6ZVxpP0+lFUHkrqtHKnmpHG
fVyhGRhcVpDpvTfV2KU7eeEwiVW6EHt+jzsTUT1GS5EIQMpQM7ctLSrF4Qnu6qMM
7eYEVcKrsoSIKL6ensO6tSs+gCAZhwTI2f2aAPDy7s+xS1IoSV75/31wNMdJKlAM
BP6gEPISJunYzBHk6tE/Nv4Ri7pIMTjmoo7Q1xliEizBF3BnTfE7ljgSBEuBce5J
lX5d0h8zNZ2PRC3pXiGWuxJoUl1GBcIGroKU/5eih0JwBPrm5bni329qfIbBW415
dZNXnG+6uqRaYDl8pa5ztIwsmXw5xI3g1Q10OJSGjHfCGOk1c9b+6u8C8KFbuvK5
G65ogYHBLMxQoKiLpR7fq0zlaD4pPJXFTQPI485EYhWq6DgMMoXJxK578XGAWSd0
UykcWmT8qekxRdMLojJokSAjbwZep5iiefRdVslp7zY=
`protect END_PROTECTED
