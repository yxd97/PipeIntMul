`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ppa1uyVCUZQY2bXsl+KU7OwJhZe7aZYOzcuY5WzUS7yzvmvweFLATgAH8UdT+Sc
+rTwwADIhmZbk+UpYS0nwWx42eqMKJY1Jk991VeoPvR6Jh10YliLVDgVBJc7vyw0
mK04jWp0KL86qSBeTbirLJB79s+rXLsv5uozi/sLIcIhZfeMa36Vducm5ZR+TZWV
bo/CwszY+0sx3tW/LxS25ejHN7JY9WkSunsHXt74MZHVsN7eykhJ9UstMdAytr85
j5VQ21zsdQYh6exic3ogtBUHStUhgB3owpWS9O1m2QCLssxPVMCE7iKI2wdJSxib
1xc3FiTCAHAK33UDNVP0Zq63VvvQ+7+FZ5P1UE7JpDnlvC5C4W+94I6p6v6HPhcd
qhdvn8BbHluHs9yUNtkrAEBboPzVWXPhncfB0ktheNOIK7hhcK/Ng3R9Cz+g+spA
iRZ1ugGEvVFUDFSOMG0vy7V3Q7KqhLNhoBIyH0OamHborqs68QDpm2+ANl7PeHSy
ypw5e9IQl8DysDv+HSk7gxX+6i+b8pe42f3cMVGyeDGZyTSIk/NniH+8dSPdRTRG
9oWrjxmuCCLTrfiUAlwgJl67F98F3lzsKFZGjRLH+ZuQTp6C0ATPW1/4pukn230X
mJnya6l0EHio7IAidweaxsVq/iqWuPY5KrKIVCTeX9XD1azX+JsgnbgeUNUdxT8C
fgjejg7jRWUdN5vOi7SSDUotns9lGeJN1g7cUWis0ybEsTqGXceJgXTovzh/wDe+
tj8PSkNkxtL2fc5aOiIGkg==
`protect END_PROTECTED
