`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c2RwLTlZG5Cc1kWf5uX4USRNHQlatT3cbTU6p5DKBJBs0iGSaZfVU3PVaC/Yp0BG
2fCfziYzPePf4SLu083KpKuX0scCLg5YifgJwUU5pNlXQ1tq2sRYoxDjjGtwe8o1
H+Jf3E0N5wIMFPBmY6FiJ2fLqxzsBJiTn6ZstLr+YtD4BywvLcL1Wr+CWHP0pw0O
gKde7t1y9TbK4OlfDztR/ZoIw0rH+ZjzdmEbDYRe8zknZHaBwjllc0JrL74vbya5
iP0JI+/K6FcT5rs1pz13rH1xM3ZLy+wM20inK8urUzYpXBiVff6o7koiz7Dwjnk9
RIdYnLeeIeqSzHOjy9htXsIiXePwsdMEfBVB11dTzVuagmZKrUQfoqr5MIj4jK05
8/8K99s+phTsolwtBxUOyA==
`protect END_PROTECTED
