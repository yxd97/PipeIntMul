`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rPIpgM/f0dqjlKpGEXC/L0iiStf8irt1ZaVzBCgJr7mhDmkyZozE0lszgyZcIsXd
BGlteXctro6HYBEuPckBkI0X9oRFYLUz4zoz7DBJTSDc0W5cKzFl1Cebnzc4aIQa
b/63dsSRe/6PuuJrbllMHBPUKYz0r+rx80xxn9FxW18vn8K6efSGO8l+JeFEJoBl
T4DLN2WyIJt73wzFvcHe2ViCw7Yj4UnEygvuj7X4qxELGsdnmnNLdK4C2q03xYHE
XJglM6cc8UpAT3vQYCCof2gar/fna5Q0WjI/zk1XFSVr4cWmXSkhaHsV3z6nz7R4
8GE6nj+sjKwzS56m8fCjo5UKaf2jJMwYIRXo85psL7zvO7a1weHmshPhoyI9NbxO
FoUloirQxFHLWPpp90TY/kG46wtaBLzOYPybN5w/xgEN88voF7LXDuCeKlwkE69s
MJKBHoHWBVYS1vS+rh3EN2gjXGi/Ihqzl7Coq0pdPwRuzpwzd4JM5psnhkigd6pA
+BkmIyu5Alqkz7D21hkIWU3SA/q/kk5VRdEoYFH/6a9mL78QJMl0vfJvopXuwhuy
nnxaIY93Oa+ZWpP0YH5cL3xOmjolCenG5SDnYfA5HBox31S7rVwZHNS6gZrvC70y
ZDGtTWjdjZXolEnzPopFbri0V5N6pCRqllLEXhMCn4qlmdvKRqzdeNe16SgSDz0i
c9qqV0D8lqCS4hUfy4kkqQlQv5A2XSrLnYepJ/W7xNk=
`protect END_PROTECTED
