`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+jehUsVeCJHFERavUVUp6UDLdtECh+P3c0/88QJIq0kiauWE1XpzRPQiwcN4pmvP
Oam+DsMrqMTaCfNXvtHHJ/IapsOxnTyfvSPrzJYu6L8/tShTnOyYL6oG1ZqkNfLw
wdPTYsFxNVzPF6yComowneBOeW7FpRef1AHKGdFnHDB+v5/LRGdggHiD7d0Uhq5x
XCfBm8k5vQG4XLfV+DcjO9GPDnwLztnsKXZiH5J5bi9ATyP5A3NSprwebk32xek/
43aur2C1WqD6Xu3+xD72nmTymWn9+aI/bJGDNKVEoikQiQitqJ5rQ4ChA3IS5G+s
gXCUEwqV38492X7LlVqJGmBIVMgJq/tRJz7jP+SM8kuGoI+6xzxv0srFqtr5Sl0P
hDGq4wBClNfKriP4vpprdjHrk6YFwxl9l8GV4wQDMcGA6uwAmQnxCHox7sbqHnyU
+wQMgcesAHmRxk6bG7o39k8vVkuUtFYaffe/c2aKuzIGr+fAB5AXuU7ImXZC/F+X
`protect END_PROTECTED
