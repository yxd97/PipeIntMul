`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNhXR/VRGeGLdyHg+l0V0DoDCt4XfUCbfJFKNZBddKeCDTn5rrZ9GiOm/HzCRZfC
Jiu6+Jjj+tonTnFEv5i963zF8A5YA7Vd/DWca21PjmONcjmw0oAjav2C9+F5ZQzM
5yYiP2XimnzJx1D4wFpQNxW//byiWp41ffgXaDJ+meM1+NuEfVjcwh5c5vPWWRqx
yNH6Rjje3oBCEkawNNaU9ILux/94NDDnl1MIr+/qhgc/IwUbP2L4LqY8krnzblip
XaUFvUJnrESTCy+8MrGWUg==
`protect END_PROTECTED
