`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNV+PBItAPmHzsC8Xur0osRSRo7wzv/CToj4RSFULTR75Hh6sqLGigkecrrNH2sH
QAoW63kTlxtPAEjfbGlidtawG4BBMtK/ES9MXXxnulZRoD0NOdxT4zVVR7hp0e1O
FAxsyB6BuN5W40OfbUeFkKklyvmnJZ/JJbf2XCNW0zJLFwxukN6OoAb7T00QMcSg
ewkrM7+KxEUYBVHV1S9iLcOBJg8bTDSUXhNnHSQwQUDbN1xro7HXzT8XLM+0mh1o
t4kO3Yf3Wh12y2iouAvP+w==
`protect END_PROTECTED
