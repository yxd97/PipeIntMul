`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0eINqpC4kAaUAlxGIGP6EqyV4DFxvWGxtSO1eNmmx843xlarPbogEB2a7TEBXNhd
qLwxwFdVsSguyYhB9FIYWS6KNC/EnsAvOEPSS1OcrklhsPzNEYtJuV2iH4dSLalC
/MwZa3YQi1Z7894mT7sNxvidcK3u8pyM3dob7+cwBvTVswUnpaXkEgh0aAvdPVwo
Nfb5ixptpG3+4FeysHtPfMpXu/7BCYmLUYC5J16p3ycHYJa9Dnphp/TxmuRf0eTI
1c11CLEWdUjCzv5RAoV+VH6jxLpfUDcGh+V9o4r/t722+I9mSHdYFGFYSqLlnZPM
8x5p6jU2W5+R5/zEzJpfXL3W5ixi+VmXLjmJkvCoVSemymSFVc/9HUuFhm6Mw3/S
8z0GJBb5/G0HTVmpES0nlf7uUP7vOiHDRR7j2eRhgdRfKBJlXgxLrXV6cL0YWMUT
TWNhW1YKYq8jqZINY19XohxRomdSKKLiXzVXlQFLdYxh9L5Ae8duAcQMCQ5e4ur0
wH3KXHwB5WXpkmszjisJODJ11AnJJ9eXZCKBX2n33x2kbUWKzTU/iDNXDNFaj9Fc
q5JDRaZ9VEIPP78q/GPmBw/Z/937VC3UNTX0Jfe4fKdwTt/+01g9GRsW5V/9f2Z+
6US4FH8+04mYg5cS2BjeHjF200ylW418MSovIJ8Nv+6tM2dEzVmoSyPUCrERO2LT
YdaMYe27jGR+emmRxoO6WlTkxeTU3GfS3zZY2bUB+dUUVbSziufCrvs6TpAe2GfW
7UZq7QeiWPvAa+6lVusRN4+qldeLhqogkpnOm+VlUFWNbpx1utqFOXAklNPYEqqN
LahMx966NqEHYy42O2myeez9warLcA7GPGW7YOzeSPgz3v+J+uMorJr8uIuZ3CuC
XdLM7qmy7KmDSZoyf2/dX1CyqptiN5ZGk+5k/6gvcw5lSSEDnBQIqtaIoe+7bPXQ
LHe5BWrk/b+mr+/nniu81N32tsCRmqO+GFOwOmklF1Gyzmflq4G3f6TawZu8ecdW
pGWO0qCv+qWdx8vOZEczBcRgraOjaUcbwpNsFG5JBX0WnCk+7N5UqC2ORUjLfE0Q
u7wwyoLv2mQcRTaEik/xdg2oan/AUxe28HfrmnFrIE8U5k782crvVt72oBqycuC+
7ibOcSVXafoYPXIHToE86VhNPqVtxb+fyG5WwUmbRn6Oq2knWSyxEBlLm2HEBYRe
vlpHeGRqYq5uSJHuvMECJ9Xd/8o+OXhFfD+cGCPOzZdHQiy3ChlFVk8+lZWxP+6c
H89BMjoiNDj+v9mdBb7uyza8yx/BZGXVhTfXS+cApBo5P2GwozRxF3CKIJX18Il0
7vsquxxGaYe5tlb965oElbxITlIm1COXVUKndsblvJ00MaCAW5hcE9PiuHQGElHm
QHGiqXup8yzdulu1xF3U15wviQuCYa+tbX0mxFaW9a+lotGf5DOuZ8Fud4kqv7w9
YhP6plut4gXqK6j1F3Gu/Zsu+TYtqjCvN6I2hJOA47c6e/CmqIW8prGrvsgwDcDe
MMn+MCaqitgoHjSksXZKqUhGYyH+6nEXEqQSkYvha97iocfKT6VGD5Mc8YEodrQi
bVFpzCJXOVtUQgPsIfz67wK0ZUfKWqyJ3mY+Wn6VUFJAOCsCT5HQT9ja9Id6Ex4h
nI04HTqww4KKhyBLKrwnokG5o27/rv/cnk0UFQ8ixBnyY5fHr9NrZ1sjf3lpD9sk
ZY3j75+hImClUgSTt5jJT80BHiTzEcCgQyLLUluy1nXdjVgHkY/akGQljzvCYoA1
0wcTUGT2MBbgxI0s8UmNQbJPtHYmd7FERY3aMxe+OcrromdRkNR6LSEJVB8QtFVF
zJriGhHdJ8oSqjLjGYIGJ+9fqqfT5yt3l5iiRDj9SbDpXAxgbFNwh9yefqRLkLAU
3oWqJ769qqjLIxh4sgHaIsHz04OE6T9nz+LCiXO+QuAnAlE1r0J+clVpw+M1gFSt
gzV2wX4pAJHFYJhoaHC5jRKErtXvJo9pPyISUL17paQBn+2OGRoJC6dIeD4L5lj+
VxjV5ektXCOoV8eM6pYQZaPjMwymZ0T2kiM/NSsYezxAqBmPyqIV8vnKb9HtL7vs
mr6dj8vhVd8AecjwN1DfMeWNmQOxmepD37ScZ4RUkIVGewTNXTJZS1U+CMFOr9fy
PY0MxCEUmeCszVj0O5kU0NxE4zc+fzSEUOsxLmjUgSKZYf0qT6PEYHuQuD3JrWKE
Bdkv3NlkL/DhRogkAoiR50P9KuktmBsYlsRYns2yRCdm6qNjckSREJD8HfVVxnw5
Gu3ZkdDGwIWS3p15ach8hmQu6EHKwXbSOVPSzgbjGLocYDHz/ArdKYWCpi4ZrnhE
gOWnflct7p2jpSjp2+IKAXR/ailjHRjbxceH1aq9AVcCOhcpcqAhyFuiqaCOKQvT
jC8ithG2QKzVpzCpXMl/J3E9w0Qkdh8UwrNau59o7Ttv0D0G3vAq168vanrKNJ5v
h+9F1ts+INeXD7WFkV8UE4JRDiNoFUrVqkDmhb46ydA6aCwIqL3lNXvqozG84LqZ
ma0pDHsT2eOUlNChtmQgeedzLCzmJx6W3jmppPXOzCbrG7np6/8o4Y9IesVunjak
X9QBTvhdJVn84EtpHq5+HtNdO9Ikdp8phtNdjOcm7bxqK3IzbXOSslwQiz5pTfQ/
U+doUZl2mmCvuK9p8/TXCxvzHXivj39nTENFk2sxBh1drRxuF8iTuKn3mruFlUs5
Z+oZIQbLqcYBLs92/bDy/Mw1kF4/IamuhDJwmg86hP5D+iXzxlEwCMshXpLi1IYf
4P2eAKrvvC+MiVg+tJRoZLQnxMfhMVZ2oQU8tg0E0PLDzSnoNJtIp3Q1mGLiMp1R
hjFeA/7JRf/DQPYuffpSPf2W6ttxQQkcprV1Hk0AFVcwv3Y8BRGMixH8P95hb6xH
c+kQTQBbAikhJy6w8doXsPaI9sF5MON0f7t9o9znu3Dp/SgDQxIx/smxVHO+XFhJ
aVzAz8uwaZYIvRHASvY4ndNU0sbaEBqTvEourLsS7Ub6Z9ZeVlUkw4K084S7V0M3
oGecAeM5saLe+/+BZKiaoSrJmRr/EZI4ki0KMhDqlbZ5X2bmAxnR/qlUWDUozLIR
C1769oSHmmlCnYDr5ruZ+P9MJEWZOmjobfM6UZlWRavCITk33MGaq/Vyel7T+Va5
Ij/2u+yM5RladSkSvuqhqKLy9L62gNYrMXqYGONEERZakSpyHLAn6nTv+N5ye26A
C2ZH6u+a1zd2YqSnTNJ4B61J2SpyV0KFHsgg9Yt5IQCpsmwrAjAsORgZM6qaEbmO
K9CWsHCzaBbuuKH70FEJP6WOObHOFWTjmN5Ioud7NTzbaEn3Hl3RHKqc9h+DnFai
xuC3K0NvTdU3MDke3KJzotGpPKAK+iaYaoBRbI81sp/xcGEeZfReOr13pKfxZhQY
DWzzzb7M96jbU1Amg2Fz0osxnJLBdFACQYR0Q13XMCV5AnkQR5qA8TvzNWgLRrRp
4RxJB4RrPQ03L3FxnsStIyYOaaBrrf8muQQ2nIa/WiXdqCj/11ToO5N4G5Og0IZV
BfzbH4iEjbZp+XLyJYmMSvOtu1jxV+7v4of6YOmIdsXb8nx9zn7l8qmYnWgR4rVN
qPm5ABz22CkL8NFqtQWdaduKeiOEuc8IqhZRFui13iMOXR2rnv54EeoQcwiVNGh9
7fR5hNmnOsZoRL3NSC3nbhZ3ghCLDJncMeoEIL+6U9+p5VhLNCyKt+wga3UL3jcO
dNuQnPcO/NUHSiutt5NlppRKiv5fPFp5pVsGQ38jCLQKydI/RN9Ads0i7PyU1rCq
5IVN6f4ZKJi3bqCn7/WfpVgn6vsj6NLjc/T0Gu2/mY16qEVsxGQGo9tHgq0FF++p
CE0fFMUbIPqr8n3HHDADr5DBL4cW5SPYtJVn4LHIVn6J0KO7M4EvUZADzo1Yezpc
f5gDvxoZGPdxexILrBqa84PxIXFWdTtoQIhmOLn/CkpKWMEI9Q+RTbTEPsMo3Ftc
7YEKL3gktgLBPHUurJkzyvY2BZHFAEE7xN31UfMCfh2UfMPtZYBmF/jw9o+9OAnz
6z/lOZ9GCHC4sSA8PK5EXR6RpuU9TGdPu2C6oWNyEvde3cJ8JSgJCshiHUUYlLwa
DGCDH/GW2IxkMGqNWyvTmeo0EmV+7x0ZXGfYybFNIWct00fe/KfElS5UGDF9CsJs
7W3caWxMTWEatqY9UfVPMC0SHSuFzv+JiTo3BO3T+MJ66+1z8FnGtRKzneanmgOM
Ynv1zu7Rukx4TQC+Cbq3YJ9OfK4oWilmHL4Dh21FQCbWpSUlApHRWPBqDXtL/uP5
R+sWWP5JvLzZhFg0UWyh8daGayZUifOzAB4yuZ09tbZfXPCEA/A8RFqN0vkdqjR6
+1VYFIdMTfMvxCWUXlOXCSO9cdLwDBswLbYXcSDagFtM4FIaPzA5XfYQiNcl45WJ
xkq1bVgo6RNE1IB9LBRKri3bNyEdXX3aVsCpr+Omeb6tc7A+b6BVQ8q9wkVcpaS+
O781JVKi8dCWQWmpac5Cw6N1SbpRtbsZ4ND8yZfnLthtx6rXmucrvYnfcoLcYLq/
afY+Azlkuw37XmWWWJol9Sn+ebx1zooyAIw6LhcyoDZH9N/NXkGAJAlHYd8/OEz+
2r+EMNd3sMVECLAGIFed5/nMJFZ1ru8rrdUVAhZ0ksI5fxagyP9TWM7cdos9P5wl
Iexj84hQs6cByv9O9bBIQyIBca5H6xVg8fE/Y+QCP2HkQKD3IEkvw5qTdVtyD9xG
PWGlOTLizfgNUCCabinGMvaL+AxPFvI9qtzx0Q5BSAtTObw4KzXokpvBOcRidcY+
MPkfI+sS3VwkHSplBhwUJiPz/cLKmPMUvPyrn+8+MBFFTbFZgAQ7dSU9j/FKyxi3
QdPueITPfMyreZTpnUzyA278IRp0r4x1OJCL/tRde55WMz6BA91KaScDVFpgjmx9
O3kklCRDEgD7EQqgj3wJGS6P2j4o9iTvgD2CaRACpVFqqkw2JGHnKPyLAm/iEAlL
A97K1h/ojk0Vm6jWIRXQmp773tD1rvBN9MgaoUwoDAbJFSu/1IQNOx+WvCX9JkkU
47dUtaoEgfrUzLT1wcm+qU4Q20XiFXg6NrM2MxQZVmXXXJeo8ScZMstYHzXyHftF
sms030qONxFPFJ2TR7s9VLR6QHr2zPEmlHd/HXCktPVzY8LH53b2+Ii/wPOyGw4L
ocRlxFGCIT7emBKq4775nOJsVXlFFZN3AVvqeMnteSJ9qgyTSyFsnpEA3oJwBjkw
EisdFYv47eCBwSQBxlBNu3vH0ZWp/veuQAprfkPaKs8fkZd5V06fOQJ7jY54DRus
9+sM2nriq/AbY9kz/5Y1mFOKS+iiJo+Z+cNXmJL89RegX9WYrKTqbmwxc3NeWEnr
MZJDPZR+v2GEgUTwpqBqBijKGeI5y8BT6g77nusSD+7WPaKyMe8gS37NRx0q3YD3
QPKfWr2B8Yxw0T81kxQGvzJn5S2flfE+ZKKwRJDrqkZ+go0XEokOGIYVEx07Jugf
OhyvWIOGb5CCDQupMtRA1O1PoqgtRKyp3nriHK7BWjn4So5Zh0caH1kugvAArXWo
JzHPtUZmODSGdXKEMqKN2zzUyMDLGi2eaMJbj0qrCstm1s4ZC7AuIoKqtSohFlVi
v4q9qhAdmdAUcawb6NeiDNk/t/GZm7PKADsM8rKEsDyY664xYVpNpu49q6iHHl3W
GkbDxw0hpjQ9LlmRb4buafctRQ4PtN5q6DNoM13QkDdwNu5zols8mR/iHK7IzFI8
gn+vGz0PrNww1AzFioZzzhNLbnrTSka5xz3oa8XKsJLwNV0UzTVipkCzvY2mM2fY
nmN4RmikvavCo7DW+dFEHdsz+YeG+GZ8iazOaZzPKFbBT5hOIs1dBAF+a0eonkWg
3vGaXVhQiqXVVjH9soZ8WGbZH/SBFuYpuQYgsocND8ZKrfUWo+VrvHiebGWSINbU
BZQboLRC6jhZyiZeCdbIURVNVwVIny/M5MHTsS0WI9xkpr9FdjB/CkL7gB8OY7mP
RcQx0jZ6vznz8cIRf2yry+GynFuNoDFGVx/i9F5u0EGP1XI6oKCQtU56x3HO7PHv
le9yFn3Zr2b/tWSPeLhYTerVl3k9mAumJOOjRIF7A1lgl/DpUwNeB73Y8alE3Wdx
AgZipVWgkfsV5H0dEgsA+GF1r69zeKsjqCaWybZK6FUj6GGWpNmLLU4nB++cVZ48
suUJ4eyeGndNhau2FI3uoeMknIZl9wKS2a7gn769GzP1UCJ2BXr8t0ytCTL+8IH3
uvGb+FDU9ZncZtjbImKdsVaWmSfSSFnO+3Dnui8Qq0s8baa/xp7d4bOnywAifDAU
5CypxhImFJbLx6rOEjS0m3fwWKqLnIMEpJfzcvRmkA46vFDbnVlKmvXpEpWhRNNK
K4mGzA/OUUl/aKoAU0uJtzSJFE3cSf3klBfmIUbFgsR1cci+ilI+JPluATHbtRQ3
akdvoDsj9dMKD7PM5Bgh3Q1cdY6P2xw6gr8iwsm1lUCxwaZCx4O5noWxIkQS94ad
arcRfd3OtmNwrQBcdQ9S49Qg+Yq50DAfDaBjj/DWHeDk/AVcK7uF7id6GohuvMA8
SbA472+oVBWFHrRnArL0W0ExA8yjRubCOEaPL1LPXJyZ3IwAaMASjZT/dNJNUjm+
YIyR0g+dR9YbtgKouJm0j4Wz14aOF5t6C/SbhTgy0dLRwTF6t8fYos/Xwm+CstlW
giXqSBQZpTNN1ATKBs9vXIHeuGGcEH953El9pzgowuuPmn1nYw/q/crCgAnzWI36
H70uGcLlzo/zUYIiJW22W242NlP3MnKNAQh2NUnFe0ejcoTh1f2QfZd6fA0QeZzP
incFYdYfotF08lRi+TiVLLKZX28fG+vgJDwcMyKIk+ydrlf2iMFhP6+/K5dDFIDI
49sKiclR3vST44geogazhgPzjKvM4OXOYSOzWeCbe90vErXLtnSJDKBG1sldaQ9q
zriavnOG43ZutKieVjnue6ixmv+YHz/CNSwk2t8pO4lLCM3jtFjh88unXE7C4Ta1
Ta/9I8bMNmqvKzxa93XxFMbUcL4VjWYPnlh+pN1vudb42Fl7KxSbwahBoM79M5Om
rI81LRxSe1Qn1+Hngp4JjD/ZBOrtAJo44o0f+I32C9VR9zy3ifXbivdDiDu+849/
4qpseX7SkohPYxA7rxLKCJlp6gfPqweodjrtJhLXOIBUsGeV8oYs4O9zkX7RAA9U
oIvfTEqhNYPge4tNfMDYZt2L4V4MiHvTKM7zEg28GLcVvl+dJrrvtTCVYKfMqq9a
LSKa2aS2rOT7Z/hykyInps+gdlGrVxNn2m4OMVbgmqambBbBZ2kxMsfh2aAKoFZ7
n0n63beRXU02/CIFn0S6kyfoGD2GQNauGAD4qowJO/KJVlHV86+5iOIvHLc5ARjy
vHi4sUbqGQjrrKr+Yx9GoEcfDCZEXNgwY1MFmToaJDoaW/G4r/5W7pjXFbrE5vBH
3eFDSij7GiYkLxKmjEoOdcDTq3lGPhx67rhg02tl2gIDwkqf8wqVneUbYYG7VOMr
4M9x6kw2ObHBV2TOFoAN4dXhg1zAGnrh1/3l4qeQiiaPLAhg4M+YQ1RLLYRWlEP6
uNI0rBbTX/Rwi64/7CcAaHUp3QRgyZfx/Gf3SFWHD7R4aCWRLanb8O4JLVcybiEZ
mF9ocW9T4TyB19usZ3ztrdj6PngwPkg/S9Ez4KMZVWpw728iq3rfMNK5Gmr8mg06
wvDE8wzscsZ+IKLfNhLuae7NHsv5pnlQrP1GFaujdClBBOcCXUmngWZzjb+PFG/j
5po3yB69tn091CyIoMOFIFJTtL9LhInzzdbqTAuF2imDjVNy/jm28UmE55309h3n
G+/zMnyR6t1VcN+9WiPKi9XfG4xS73VTQwwq29FlQZqSU1+PkP9bcWSRTFt2+Gnd
thmJg2mP9gVo/osmdcGccG8roikJ3w/tdg0PJtxo4/BE4A2KEMnNNEYfYYxwIMi+
45Xd17i58pIQnD/3qZwBX4vJIZ871JFbRrqZtK85IuwhLla16igcxTGzsePTvs1C
oko1HPPtejwkeTqZ8/S/lb2BvBOiQtSYtuHFEwN42y/AnrpQB6oftRfx/kpV4b5+
rYLETlETItCttEWAWYCP8hNoP+7qnQCxHTGv3SSlEBRRfpn1wvJ12ih0SGjAkjAh
1EIowZ7YcJ7ltnTCGi4NOFOAdl/pJnwqVay3wvVXmeDa0SkYZ2oft8ei6G2foq83
MambpXOwxhPV/EV7BZmtTHTTGDopzmbmUgNj0xMeFt9X4p7KQ1nmSCTRrhLelPiw
P/jY5sdgi+iP2xEQ6ytXU8bMLwgqCmja7qs0D4E2+Kui4oxJYjhcOuu2Jnsw41H1
1o19WvaBrjt351XShttM+8V+T55srHcoDVUinDlCJ7s/7gdQr6beR0WcVxZNgiLf
K0xflZSb9ysD1XTml4AL3vnum770Hdk+yLVtxeR4Jqu8xBeqTkDjiHH1vPo70hn0
S4xCSObw/+YqIMkLXpVMu92ib2xgoBb0v2lOCcIfKdPxZ8T/htgBzi3ukMtqJX2Q
KrvNlnpBsyEMamB4Q5NnU8wK3Zv0bRQfjwJDkw9/gTGGYx9FZnIwYVGVMGMuxGyW
Ss+XoK6nNLgsc+l9/IoFO5TIUlBRSz+U8xI+k/2aYQTQwwjnq4Ca4CN+siFKKXIf
U3rNIqHpPHehThs71dTRG9zyvvzSRv/Y1kusF/Hh9SEQ3zvv8UEQUW8BKtURyIMt
FkSKgxoGG1rTFZhRRiaIHaoDoxOAa4dUH3tnzVMJ0pki755QhvRww/aCjnz8BK2n
sS0NUtEJ8511gREFKZjWUG8jgXRDNUsZntfF8JZFT6PAyBxUOVkLdNcmFFrvKQZh
A7ZSj+yuB+Y7Pva6XPpuaNgyCwpFIhiYWZPMFarV9Tea1CuODGkGlcqFyOLdj8e7
AQ89b45IckTtNm4Q8PX3j73FHVXYfou0YQfYybZm8A/k76CvocMs3E+f4/rQQXWc
QRvpC0+8ihlbxORK5EzJXu3tdOwinqAyaNzv2pocZOoC/kE3ShzmNHanCwHksLfl
lZy8QscaM9MjIdXGu31qwLiM+Tr4tIuVFLZlBXeMgztldW6bstZ9iSiDJM7IGx/C
mS9n9JTKePUswvhULnS6vEftvbB94SSNmey7+/qn3XNUp2NW1y0i+mitExzmF3k3
VYJBaMhjpFEim3J8vVWf2KMq/pu4LE8xgAloF2epIZmKQ+Vl5pUJirkZg5RUQP+M
FeEuvPfRTCBr5ZoC3zaCUBzMtwplGRl6ohY5xB1FORFIY0Ak5M94I9LQQ1lIY/ch
8LIB49fV8PJGFkwKofkm317ZJ9DzrH6nVmpVsL/D+4smcv5VUsNKjYk67raa8alT
VulWuzT6iG+cOfjiXwNutY4GED3pwBQ7h61cuAHmIavXRwmxU2nj/ot3NZB+GORb
surEAGDgbTXJQUmUhwiX+w++P7RYhdhC/AnF0AlaZ+hzp0/pmP5AuAMEpVw31V4M
GyIsKGUH6g0KC1cUwc7Yr/P1QFBV+1F8EKBQDOvy7GkWTSYRUScusBu5G86m7/im
5pGvc2tXSIv/YL2WPqFGIAPoMn/bBdpNGJKvQceGSP2Wp4cvOlcsiana/4/QDjrR
x4b7cQhozNtR8TdniCQURBmS7d1W5iqhwh0YPcLAqtgDmBnM+FC6t7STeOmaIj7g
DS4reffWH8cM8bUjpl00Xd1eZkjw47m4lZcGDy9Udw6wyxxbK3hlmgPd+izofwLo
eF85lPMZsxDasJPy77EB2w7Sby1ZC7pi2BODkPwDAK5vdatvVUtzY8KG9hk8ZLOL
kJp//GdOWrIjo28euFWJHSq26CiEfnU8Gf62wk8MVbFfOv4DEWjLMjUVeHV8nAbq
4GzkdM7a31m3OckhML2ToFWmdaCkGQyfMjHM9wc2u+czSEm8eRPlr7sQl1ZpEfkN
v6oTnV7LB7SOD30dRDExoQxPUbeLcHew1UM9jzo1Lv6eSXImBjkJ9ar/pMrUeIGq
QEg3zqm2xRcO0Qq7Qm6eX3IMZAAJQ3/hFFpobfHgv6gJfX0le36lWTlCpOs84SV8
ePlLPdD92f6Gii9zxT5l4jnvq4lC9de0xfEEAkOQ1taBtMO2d0x+rNmt3QOxC6Wp
gKk+Y341Y9L2qyY5E1zOe7LE3i8HGpZYxiPsaaXXgsAAh353fMRNKzM1KcYZqJsz
zmjr5VURhYIcPtsoHUZimk99c1RxF1o7c16jrUi/2uomZwpq2mCBUHXM4/n5vZlL
Dkm2JsOTAaD+EHSOAXWKd4vF3xhK7BirdFLsOcEWuUU+dwlZrSzAMbIuUcE1tClQ
Kwp6JTjWe/JsYqeEC8h6c+/jhrnBx3MWOgXqPCscorhp9g6D3MBFzNUln32SLqc6
PauOwy66r6pLeksd+HPl2kbzCeQIITRy74UAxyKrWIm4MNMQ0w2hq21cro1Sdfbi
g8KBttg0I1EQZApw2ZLP+prsksKiVR0PPV8YY7Q2wQnO26bkzEH6dl4lFsRqYb99
SVucswEkUuMmsazGYZ3a/8QOD7h2hbS7SPmezNen05Sds44ywTvGweYtJ921tLsw
Cr1IzIj76VQgaOApfWHr1U3ZDxKReEdWZslLL7utp5ATQi8qTPRHqYG5aX6CvOGR
mdD7fwigIc/rBCQNchsSi+e9672X7G6pTZtBvnDDguImqyexEGzunEH/lEa8nQ/t
Odj2/wWLoQNPAWlj46CRrTmxd7Mt6Eaq291uMxaouaZWWqZh8Yc186wTTeQDqxj0
j9PYWOxX+ZRwOGlFTDHtXaH1WYLCzjxqMKv/kOErC5pOhh1VJEjQjqpWdJIp/KPU
OaKaVSoLE5QOATrSOM8b0PzmDzpRZW0yyIAHyHt5r934TEofoxFMSaIFfPZjwfVk
od7Fq/cDtoQWUvh5nvrT4IwScnsCn980w/CYF98pc3Fd/NaIx56NxjR2d55ssHJk
ZA7QgPcGi04AJWEiG/xLO99BA2QddrxKZsLN+G3/7nGtNI+QR6G8jDhOrKnU4VOm
fGi6qFHAD9AsjzCCXYREbRbAAu4ppjqzI/JBwRrcWNr2m0DxyDF++45r9R5Ao0GQ
09FJqJAXWNnes9yvSMy+aQrTB9mDyaeNTbthjmNJqAKaF8jOibjpUxF0GYJnv/i9
Ol4CtBwMaiykwyjvsTklhzWp6frKaACF/M3xbXjyyrZ9boAAH/p4Hw8bjP0yZtTP
BrcHxOCw9nF+sFc6pUmXo4+8G4+P96cWXMQ4ry0zdMT9AS2GKSVZm6iy4bHt+Yqi
+UrVqNoQWzlTIMI6nKZCw45cWoCj1tG6LZ4xyE3DzCHxLD5I2HE7BkfKMY4o/iC1
0J64S2de6V9EzFrsquq9NoOGm5p0RsOF6r8PMMKoHcxwh6VmZMVU8eixTQcGqhBZ
hF2u3XuxilQFpmc18G93XEV+Ji6J4PWibvO0K5L850hijl4yWpWbCaJRro9mQ/x+
zuOhwSy/KhQXI3rIOEKJBZaYtfy6hSJRo8P+PyFhX2iZi5FiSvRfIyjG/IvarcND
i4U+n74O7EEQjqINERt1KmKDM5NZmlgLj8v877G6QjCbE3ZSXoSpjfNfi6LjyZRt
nl3rfVJhNs7IOLuWqmO5TLy6XCOoKfBzFk30uXGXoFbix5XGM9HwN+8JgdgN4HD6
fILHJNuuzpIOsO8a5vUz5tobVXE/AHtafcLaszRW2KdEqHzaixEks0FPs2U5/dI4
8313E6HNm5V7l+rtRbS/FdxIQXIDYVl++G0KTzjtgKLwMAVTz4CXsNfTbcYebGQG
+T/Uho0wQOaz3NVhI1ymH3m8EDI2LnDaDwv/m9Oucijec5AwokktnIEXLkXQfPCg
9+IcE9YH6hsbF43E7IfVJ44MGKezuRZLxG+m7osDGbf49G/Xnbr4ZBiAcSQ8/EHi
WOP8xYDJIFHZ5gKnPNWW9VhP1GRzZMbK9J2WahkgaG0D3WDLlQEsYB+D3oGIotqh
CFya6UtzDlqy6K+DtIKNz0AQu4+J1bbTGWyehjBO0l62noW7nu2qfmO8LpHcvpry
PWplh9W8pAsGfwDFvHJWuU3n0sg65nicUAa22HUS/DlGQ24FZcrlL+QPx15u+Jvh
0bsHCcrPdQhz3TsPm2AZo/HHfcxwh+rITiddhRzdFsF9tJqYhL5RIMcLKoIxOe8D
Omk76TlxIIAjGfXeBbpNESy66OXbuprMxg8gCJE/KptDYzfxu5rn2izId4sVlrkX
W7wAKQmt0SFlD+u1bvpn88W2A86ok82qoqq28cBsXGjvPGf1yoyeJUgT5/HAZsHC
Ui95BBRQMHt8QKRna9AsgNgfOlCgrnFSGCdgjg5M2wQq8OyFwZQtok6ufqw5HUbH
vXzHJH7C/AzLdIR/wtuQN5GJsPvTWstExe77W8Jv3zDipI4Drx8as1kOEZLW1XCC
bQ1J0Psz4Dmi2fJnr2xqcoz4K6FMBoioBnxEJiJdfc7/oPnsU527CZxjkG+9wyb0
8isnrRG8SqDdWxWwhQ0yUH9k/3F0QgPIPl3N3+n1SaQgmAzM03nz4o6ymlUv/SAe
QjM5f3lwX+LiVhxZMN8zu1sXY2oOjAOx3fbEqgbqCg/nm69MBYNntTeZGdcpVwKp
E01v2NNV6Osi5UrmoyqHkMhV7OvHahZY9dfmkU2QpjcFf80SV3GLAPKkdpoD+YJ4
XzYs3kTYAFog/kF21GxX1uBwarssGuVLgqdT6NTYtzjaYby5PgMC5+xloG7mJ7jx
gM7U5jwC+iNr5DcQaqu2ik9TzQ7xZBhnOgc0uGx76rrxS7hmUGGQdfLENsM/pl3c
fHpaOJZUTO7f1KmNrBMvQ4uCxwJ6ZgvHbsz4lyrUpH3w5IHIMVtJYBSJvLxy470J
1NVUEqSvsH+2nkQsXnH2XXa07e5XnfsYi0YXKvDLNE8ykBACgMdjGFk95npextuf
oF2F/w3BSkT2LApDaj0UEbwfIctXhDDWLpVGai5qw5EmRZKN7Ui1Onpwa/0XG8r+
ipgOCyLkciRFpJEQNMxEpcJxUVp2dcys60A05bpjEpSzGHaeb8RXlMtSj0fLpFpe
LTLVWhNraL3Jln+ptfz9HTYlx0D2KmwsTaSkxpM3PVZNxv/iybuw763m69vpXUNT
iounNYXu+MkTwlXsW3qV9lLlDZmumvSH3cikJ105k0IbH+wl33U1qPB3e7Q4EBEN
wfc+8Rc/HFB5nMJTwrKaww==
`protect END_PROTECTED
