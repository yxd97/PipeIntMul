`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zLof1Ik8qfSANY68FHMJRUIQC1pThtQTGjM0Ph6j9lJXqxuG/DXMNUCfau5KRRL
qe5ygGPs1SVQu4rWEi78jPHLsI/cIxppECkZnepu37d8AVE65dJoe20VY44HwOO0
EqWXpqaXMVggX12AFWUcYZSafyyII3XPHr3/pAQTyRiZI1KI70NsOyEVA9DEIbbw
tjsTsYNwPfenUukkjt3eOvSH9reRaVWtkHrl9F7yzlEDHqdlSglXditkpYGNwSO0
SIFyld1AbDhj6PZHmsDEKZKJs3AtQm2Grysq7G/xqDGLO2zvJ6thcfKAoZhk4GOD
/VXY//PKhR4XRYiFVC8LBi8rAouP5CYRi8wektmckGEE2R1spEp6uSiYTi0BWG/P
KoI7JV66Hjacqf0pymCb+cIbt/kSqnUFAmnVWBUCoRlm+utlQ3WOpXP8PcXXnmNk
LT0K07DhL7osmOJk2o9jR8LUxL6CoJQZ/JYGyAGnIoGIfF9xBNg0X/+jNATG9AKn
4FBPbvJtFWJjSYHvRTB1Uz3klpqKJtRqdX92SeYEz75qKmzajOL9fy3088aqqzxm
kI/wiE64NA2V24w8tAmUrzpNWzb9mKorgHYFBdBW5MthK/1yg+0VOo4wQRYocGng
TumZvrGaZdF9Us84SNVAizEzlZxgG5NlSRkdnGeiFO2hkDw4iSiU3FhHRTSSpOU6
+XP8ibC8OPIc37Jkla7CLs479PJGKwWSCyrGXSOky8eKzG5d8Z1/E3xZlhvcoLZJ
OsKqBj6lCyY0fylJzRcnCgQ3DfEgWaiKWCLNmnh1xeDXP62wl2pUehBFR2sWwU9x
1tkY3vM94t2qZSftVkexIFCDbe1DMDEI9zlwbFiw+0CZ1zO77eilV4a2y2rpVBL+
9OgOg06Qn4iHywRm/T/Un96L+eue6zvHcrBoKqAjCYlAUl4cMf3AxrRfhhBokDhg
yX+oXlUzWEt4jaJO94412ynSyO5fYEiffqnf4LXaX4LJYWvzKKrhKlDEnxbCdV8t
FFLCztMChLufemYCxbmkaggs+z/PoPlR1ScLcthTp4hxuB+MZ7tnbZ1JBl+67QJm
WlrRA+1miqf+M7y6Ex+RQECR1xtvA0GgOysKOuk8Q7qHlr34JMFZCZGpfC8D7Nft
nrDGr0nSAtibAVKT3QwbpzjnuUnZvYdqJhmUQ0ZiUhtwGfTu3cE17tnSRIk3P6h9
5WXycRa9pMdJeA8y7ygH4RWDIg8qJ0FrYUL0jSdEBFCmhJBRunCfStXCNhfnE1gF
VTJdTni9dUCdHT2iwYBwDwVPkUAQYIdNO1nUF86++rJw7CmcrD5Yjaln4GJpR9fO
idvgNWF2J7c6aYRXnthVYT8tZxA3oywJIW2XTlQ5SxUDB1fnZI4ubhvVSyVSL0yL
0KpIow0bKorAr01aoNU0pp/oM8nkYo5aNiIJNrGR7pg=
`protect END_PROTECTED
