`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O6eIFmPEUfk8PNW0H2XAY7dcGo+yR+5eTkOfmBduD1/7EioorW573/SPCiAivvTn
dvvhVjbQZsuZpWv2xTw2w4ZUIYgs+jajozyVVq1UmOCwS+Ly1SxySQ5mGhYOXE6B
vFd3fYPFTOsj2seo8nxZQXXmUYv0vBnTDHJiObV5EtNhpzRFI+xj73RS5j3eZ3CS
UpEKaOGTZtU8eiUHHmBS3t0j9LZXVPr4j+u6fcBKz0VTNLwGIlQ/xitzGvYqWRxW
t+fDd415jQOc6kGp55DaHi43UeNoYd6UnIfbGIwikiwkWkkd+He78iyA49r1M9wp
ulQFxqtr3GK7cqcuXCLafo4gFdKphIs0G+Ip6oyceusm2YltWE5R+9rHWaHSwwV1
sdz7SYdBmR1xczCLaRaQ0vKoATxY3HBRUT1MEq0rq4l4ZE5gp/yRVn304wDt/CM8
`protect END_PROTECTED
