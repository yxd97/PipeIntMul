`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yu08a+StLTScsk1BYdDph+DRLOX2Fr/qElsfaoMiPRkmhW6BAdxATxbwWujUpsKX
ifXxAAoFOa9mV0776LvC9bHHJfuqFVqtckDLXw6SzMxdQ+Y5PWEPla2ATp93OTId
GrALSx5BWeL4luz7ZQ9rcOti2lMyd1trck32X2Zi5SLXWSHsTOhTH6Ym+7+8bmh9
C2KLnl/njLaAmuGq5Ym5SUeFNfyk2OlaLCTdl5Q70O3ELnZNNU4/x6KfIR4IHcIz
PRi2p5ylrA/oxWufxJFx1tgTtJiuJvyzmW0bSsQrmpKoWEJ57pllx4/i60mMOIO/
H9TWPzpnONnJXx1rxbQS/+Kviu9zmKiXobt4uOIqYQYkTktip5bvbOd/1Ig2NChS
A60G852GFmXSuGnShAC6GaMjNJnvzT5fi147YEi93wa+UJ8+UtH8GzvUYVtGcW6O
RHsD0U9mcIYXSaMDx8NU4fvPsLm+JpaAH0fTY0KpDRg+ULzYsRryXeVtT6PKk1NY
vQ5reOOFjgUFMAyZRYyepKAFh3yWSe6PJU/uvpSnHZVd4+lKR/+4ASoV27TMl/ph
095UqEUloyVAT65aqV8zVSQZ6tOcSHBP+V/T2UFcZ6be5LuTLo3+3L7FJOwsjB1v
rYDrYPbFlt5D+/rYGCStsdxwKFHJKF3wEhWB+vIw9dXHIX8dwXwNItkIxcXvNWV7
9DEP3sVhVUMMz6UhvQeyU64Z3pqKjRp4JQtK58D7lMf3KkK4aXSfY7s4vDrnIGuL
6qnQEqtmdTMDyPBsrsB1lEfLoKGAjYAoK3qvdTJzyM/WJM474R+X2faGF+9HoHjw
0jHIFrnGorYPZvOi9kIjp1ToHMbinDDwHmGePEVTla8gTq2AU7vcU7m0CB0rpqBD
OZGmpXFhFyn9TolxsZtt8Y6J82Fm6j+Ljx9No1YRg8h8I47wlxU/0j2qhyFyhGg2
oFqmMdAPzYIyMQkYgDvFfhWiUP4EjuG5Q1bnFpuhrRtAyc6//2vjLbloEedV05G/
+YK22K3BL4yxB6lAuPg9s854NdYBbLF2zGyqDZwahSG/oqQ2rOKXHNdIyw8EZWQr
F27tTisAijZzji9O48JGs8hC7s0kDoTkg16LTm/XxHPNvXWXx1PGhmz8HCP12h/Q
Gaqkm1CHaTuZRJDNvw3ZByOTaATrlEGu+PfdQpwyVoqxFvif/uG/N7OwiOZ5OikE
VHssBWJtm/IrTY2b3Hr/izhHWoKl4333xn4sH25v9d4I2ppj2gpQM5ifTOfsmQnU
12JmIdxSZorsFGocj0+44yA++vgnXN+tlpSfHeFuCoypXhg5W7cPUNeUI+nknDxn
YSy2xj3DJXrX7BqbFMXxRoLtfkxykQXurjRb5EDFArzDwyRkG7sEKgkE8sfjX2sZ
bVog2j3wWv7OooDmLvb2vi+HI9twI337FYDYqBOGKSB7VIvpqVOrlLaR41dLVzi8
/7eyTKKnrQrkvjnChFPeTgqz2KfKCxuHnGpmreCdp2i+KA0BTNBD8FIU3cdG5Rv2
fF3kF+DOM2De4KWgcYKR+1iNDm/mL0+OLo5AzCNJ9sHPk3gG7mSpJecj9uL5HDuk
cQ5EmWz0+x9Kixyfx0psJgQEBXWJvEHPH8n32JChKRCvKNoNbKCe/ooX0IqRRs61
PNsoj2L6VWRpUOy4ia6kh35Zaav5QsW2v6HvcFTMp/2AL39b1w4rlV8+iSfGrQFs
jEj9nXc3rUVQi9TEbSNV4WY+UyMlH90t+cALLOI2+L2lXWLp8zdu4z8x/+vn4Kk7
PCnI7ZEJRfehcCYMjjB7drde8Xg2O6oSUuznoXIki1wnY2r77NAi1Qcar504FjtI
Kz3UP1S+sUnX/bpp4Hryfphpji/5yhCCxZ7j+gGpFLBPsa1EBByeavrvPMGi/+rQ
G3NHxya0Rv3BoPH5oIo9DuQXkDUnihfiWMynjlKqr1NBFVVEVgVm7NNQ3xXvB+YP
YYZwofD/FQObrmqTeI9iZA==
`protect END_PROTECTED
