`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FtGxgO58dDaGgmZ71z/bPTUD47GhITWycsbc9o2TYfPPkPPkz/2SP9DruFWPEC5
2GMilElqIu78w+JOLuNwON3DtIKrAdE2EBF/+v9GsmkwxBJ9MPSvzRDx1uRE3SIe
lWeglHjObp5006hMwPBE453UT2+htT8ua59E102ldIYSaRMnxYHpNlUuq16c7opy
ujoOc/PKLsn3QzBh0LpOLjU+R0FsQO8VVw64LCDgYVO5TMEdeTfVsFJwYV5zJeTh
dAQOwmgZIblKBRtxNUoxhOFJZlFKK/Ft4jdncCOzoS4pkKpjZu3PwSsGF7DtJfd+
o//1vW1OCsbnKxlBlInTubivCTo4Mpo27jQntdXo8YQ3pA7sElJJDVZmTePuerKX
3gcqZrlQ9EGuRnVlpm9NN8SSD8uKxFZpmZ6LfuGYGA4lnkkUPoMfJ0PnHRnoehp/
akr2DujaDW/jcz7d+LdrlgYrpP2U+gBKWhc1JYH9sBXHA8s4bptqtelrc4WhPGMW
RPxKTLppLuzYp4fqwprZi/+9IJlZDeD1iKNWBCHN5EAk5CuH4/2YJJ5jLrJfO87t
w9iF65ZS8RGrrfQ+fGMKqn0sNNUsigCMhk9/+sN08pOa4q2CnNUsswNj3UN87txV
qk1GNACcfLjKHULMITUEadBJu82ry+6GDTbcx/n8B11lRFwucZO9jQvJifNk1JRN
oGCMpJwotgEROzYnZfz7zXCVaFaGfX2tQlmFL6jvJQAkcVNI0pF1/c2oOXccOV9u
2yf+2tVb4s00ZmuiyWWHJWVjq3CKRMnT0jl+0p/UpQx8xbLcbeuM/5uRjkCjAOfw
CyZQlJk3itEU3qyYI9OJXb+x+RBP07PAkMzdTlW3tUNADqT+ZSJRGKosOW4IH+iH
SscpkWlytrZ3/1ZFKHf8loGgzextDEa4UK6btAHMmVApdrTw6bCWig3Xy7uAtnfJ
IsYxpkNaKBmk3xX3boLVHNuLBclzpK+cKT+lnoozQS7eL0YFIg7C/b4bOzZWSYMz
l8Ns0VSnsAnOIY6+aTU0DWmh+bNeH1WfLcKpHPlRVXVDkUyr7fwNIto1CqfuHWu9
eWyaDwFv6XyqNdrcCLPEUcNjzs1skp5v5xTGxDJlNkMO5DKBzPTx2Fifgo/wlCrH
8wAtT4QTbzY3BFPcKcrfm2qNPYIunkRFHUQ/1sBW2pM9T5TMjHApVCrBKVvbBsXB
9mB++W56cOTWLhsEX9wKjUW+/jdBQdnNIljwhNk5rxXSsFc5T1TlpxQxRClil7qF
sWmpqeh+CW8dHq8iqJgCqF12OndsPitqicEGACDDsFY=
`protect END_PROTECTED
