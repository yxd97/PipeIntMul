library verilog;
use verilog.vl_types.all;
entity X_OSERDESE1 is
    generic(
        DATA_RATE_OQ    : string  := "DDR";
        DATA_RATE_TQ    : string  := "DDR";
        DATA_WIDTH      : integer := 4;
        DDR3_DATA       : integer := 1;
        INIT_OQ         : vl_logic := Hi0;
        INIT_TQ         : vl_logic := Hi0;
        INTERFACE_TYPE  : string  := "DEFAULT";
        ODELAY_USED     : integer := 0;
        SERDES_MODE     : string  := "MASTER";
        SRVAL_OQ        : vl_logic := Hi0;
        SRVAL_TQ        : vl_logic := Hi0;
        TRISTATE_WIDTH  : integer := 4;
        LOC             : string  := "UNPLACED"
    );
    port(
        OCBEXTEND       : out    vl_logic;
        OFB             : out    vl_logic;
        OQ              : out    vl_logic;
        SHIFTOUT1       : out    vl_logic;
        SHIFTOUT2       : out    vl_logic;
        TFB             : out    vl_logic;
        TQ              : out    vl_logic;
        CLK             : in     vl_logic;
        CLKDIV          : in     vl_logic;
        CLKPERF         : in     vl_logic;
        CLKPERFDELAY    : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        D4              : in     vl_logic;
        D5              : in     vl_logic;
        D6              : in     vl_logic;
        OCE             : in     vl_logic;
        ODV             : in     vl_logic;
        RST             : in     vl_logic;
        SHIFTIN1        : in     vl_logic;
        SHIFTIN2        : in     vl_logic;
        T1              : in     vl_logic;
        T2              : in     vl_logic;
        T3              : in     vl_logic;
        T4              : in     vl_logic;
        TCE             : in     vl_logic;
        WC              : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DATA_RATE_OQ : constant is 1;
    attribute mti_svvh_generic_type of DATA_RATE_TQ : constant is 1;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of DDR3_DATA : constant is 2;
    attribute mti_svvh_generic_type of INIT_OQ : constant is 1;
    attribute mti_svvh_generic_type of INIT_TQ : constant is 1;
    attribute mti_svvh_generic_type of INTERFACE_TYPE : constant is 1;
    attribute mti_svvh_generic_type of ODELAY_USED : constant is 2;
    attribute mti_svvh_generic_type of SERDES_MODE : constant is 1;
    attribute mti_svvh_generic_type of SRVAL_OQ : constant is 1;
    attribute mti_svvh_generic_type of SRVAL_TQ : constant is 1;
    attribute mti_svvh_generic_type of TRISTATE_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of LOC : constant is 1;
end X_OSERDESE1;
