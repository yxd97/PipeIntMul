`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+DcLJ5xLLcG27b8kMOf0iwF8XFP4eO6uhghGMR4TJkgaDNCqsfavZ5XRgXbXodB
ItmtoLOzMLAKxVrz/Xvg909dazZmaHO83LOQIDz2cQrlA+J407KAzwEl1gMvXy5L
Q919HdIrXfUNTtUK3+HwRVKyPOyW10R4MRJbHdnQ1NiYXo3RooedyAk0Dq34EBY7
4GFCqbPBwtFG9sJXHrVjGpQe954WnN6dKq8HlNcI+7qm73+ygad0UvJnd8GOOmc1
hERzZhuBTxpWH7fTfBOm6TaywiMmVdnJ1/MOvLVywtlk+m88wEIFLCJ0yp7F9g1m
ZFSAHx99zTX/QoOvCaTSV4UgbLJA1OROK27wpDkcO7rUuGCDQp8/twJybsQizAjJ
hM4qw3uifh1MJj+H3sDdYE3QpVyC2pRr2p1MdYerzafyvR+3d74h/3RnmgujKdCj
`protect END_PROTECTED
