`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DeNU0qFXteCN4tDmHZsc0FoRG3xMqgMYtOXBpYIQJ48n04bUoBIslZHgrKL7rZ5
uNRV2GqFK15tM3fWAC6YbZ0Q/fgedeWOcjltes6+/YB6hFQkWnZ48ExDi/+PWv2e
b/zA8H2EMquPRXxR/AuxrvuPIG8f7hggJbZqIEtG1HPsFC7rSbWFthPP0iECE0V/
Mlyx4lVv/AXiIVm09TgpWbMSiN4UtldYyCc44mDV3Han3wkAW91o0+px/dClOR7a
4K4uJdtO28rIR1iWNkiOJtKlRqJ6Tm74zZpasDa6KlS5apmfsHElM/0TqSQ568cq
ulW8/84Tfk6/mmWCTzFjWtubRvhiB3aAY77wFQIRMAeyB3zK/6BvqgvuwSiYBnpc
YH9ijiJ2nv/zKgt16Cj70KXSLBBrz//jaqr2ytV1tZ4NNbYQtkx0HIR4y/c9ZF1d
lHb6W0thD+tlCMzzaBX73R2Q/nvMxt+bHyfx+wGEd7te/EO6fcYJsohzh3h2jton
6JkJ7R0GoSdI4SyqAVAL9kd34oDsWW98SrNF6L3nfvxRsLExJU0kbciTqutuDNhb
Mi+iCd9Dm+U7JR5E0jbj/VuMrITuIyiK10wHFySXrG+/iClN4haaoVKI6A62GQdP
kC+HI4Zvs+eqmQ5iRif++A==
`protect END_PROTECTED
