`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
02vTVjlg35sjIE+pnIrKDHoKCoSdZDYZm5GefSRX7jY+RjJzhRWwa0tdoAI3O9Uy
FLx1dgcA63/PRP0av12ZR4zNfsGaDYJ6ZpKJgwk6qm6ek68D8i/NBrnBndAlmT5e
QAnP2yqeEJ44tXOa2VZm7btFawYWIN2MjDbG1+DrCHCnQTxDAazQKr7o+1Ntlzcf
EH7xMw/WCrggfCI6B5+FwVwiPuoijUu7OTfv5gdGzvcwzBmmaOGWXRVYLs8l+8x+
AxhGLmZQLFXh1JVyaR126A==
`protect END_PROTECTED
