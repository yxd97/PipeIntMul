`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1ayrKvPgNLgql/R+vkkLerezoV6O+EHnTTDYjcfUlhMRBMo8PPzhUywhLSkOgdm
l52NVGPj9lIHjXDOrmi7UFkTPTRlvvS9f/d7Bakv6TStGN61LcpcjE+/H7Q383CW
+fGVuVx5qMT26YVVJ32WjdHLbJRYh5Z7Ti8vnO2FdRk2kBdcmOuEBxMGYvBqUNGe
GeKnuYvcAJea/Q+wqZU021mOq0k07cLE1+CJdTmxgXoNg/61OJwLtTXScSdHoMum
YZynGvaYAp4wP4bO/ThIEiWMDVhCmvBa1z2yTvNf5IIYo/FbalrZSmPawgMAgvSo
QwvtnA7c1thn27g6LLMOUA==
`protect END_PROTECTED
