`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ju5DdD8ytXZCDdrU+2B5q5Q27g8CD3qFO6j3IqQt8B7ZZjZGSZcJjSnjEl0xU0MK
y8SlILheLy4DdPx6Yi9cJhi3S2MzMKBqaL99NicMb71Wvu1VOCb9d+22knJ9u1/d
hvY/ZB8dCQxVDCWXExKxWyCwplc+ykmF/C+oIYF9QMLZlujCe6A4kh2aPjIl41ab
S5ugOkwSQ0MWqZYecLthrlAEZemCtUtyI/mSPbL9XR4zBNhS0HXC7eiT02C4IWm4
VrRYTm3CX0KLuv6l5kYHhjcaE04y96ZS6ju85iCuj3zwr70t1ZAdLehVQFaNHp2A
z/3mLVJs65BxPpZWAQO6K9RpMJ0uqYOlWLseiP7NsRybUgrbXwVo6/6g+1OlsLTH
Bgfuq6XeyElBHUkE+8oHmUIGu0biOxcJpHWFuILfcMgACbEzyG66DB8+bkbpB02J
omTbLZeX2yiwLXEXzP6PZEnWrsA6XsV9Er/quyLg3Wqu4/DIQGRMVf0cYmPtgPkN
`protect END_PROTECTED
