`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3UKnNKOf9acps+iBrGnTP2nFsB0sM16rBmhFA9mY1BmUhtGgPpUhlNkHzP0snJhD
Zz53sssDZDA6/aOQfPMA73Hzgj61PC6rxd+zBORdWsE/x7uc1YqdCzs8qg+Va/aq
WVEWinuHF+GlkqJAemuMbal2gR8TgdMY2gHjOI9Cgq/ukdllwTjfVNEjjcwzZyxX
FlfypwLqBMoKHFINMGTDuIoUCY3ri8tCWDWbHlni3wZZzuHRo756fJ1tYLeP70u+
oPNnqoNqWYJtkoTGf0bNw6q3PmvhbanKFeLTsK3ywlZNjwUcgUR662SVPOwPPlWs
uXqWxIrdpBmb+H3nYX6GU0jsRnaqEX8gGiTNPzBPP6R88zlNbEEZPE47HY9XNfim
2dqkaiefRwOyguiXnIdRpjpAF+SDrG0vnjbn6J2mlIlnSgf2IYnDOOljEYho/KAb
pB5tRyV4+nVbqHE9lGs5QjqRyj/n1qOOQSf6eU7D27dMHFkmNICnM3MPmhbqLWKn
P42Hw5e/17EC+s6ae1w/gqO3dH07Q8fmcDGwl8yWR9+SuNxH48ivVLXxpurlp7RI
tkW6an48DxopkDvu4BNbzrcgTg/AoD23rIh8+vmu2qVooAHE6/3MDwHba6SpQu3F
zbrXdG1gDSn+Bkc40x5Ljlef1PBui7fTSm/vXfH6gzs=
`protect END_PROTECTED
