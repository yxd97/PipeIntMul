`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPsX+/9uF3ycO3oFjuj1lLud8QnZvym4VJyl9qjY6ljgxSFopRx2ivmx4ylqpgUF
9OECKZbOZcUwRW/Iv8+352wQbm3kix68Wr+W0ZMyw3f8HYALKi9Sf7Upfb+I7E2Y
cfCyIX5Skd4c97A8eY7z5TsnR8DGsRRofxlO2V/jLAmlsCnMt6E4tAWTnPl8Idsm
orGkvF0iuB/EX/nahdJAYkqIpfLfMu/jbqVV+Wh2QfspD7hMlEnK22T3I9zxBjFT
sw1vm7B4Ec0/OLiEdJ7OqZmgxK37x45AmiGXGdLvzfW4Mrd5gaffIvoQIgNyJEqn
tWIL+ZMkRs6QCOHGqTqj6DxO7zma2+BKuAKxkGdnJOC5Wp89TDJKHTmhQ3SYfvS5
uNA+m5CpMryYydl4/SJ6PPMX5g579uzp3ifJSVFrdCY=
`protect END_PROTECTED
