`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eY1eQVrB4MwWU48u05B9dfZEvATd/QXPBYVBIVdHCRIQPGdCzXooYAyXfkTc4IOI
44D4gf8dZ/+c26nkhQhqe4w8+dJENUb/l4zS5F5BvBE4wnxEj42bp04WHGm8cis8
uOprEucu/oggxVaGaaKntX6MlEiGLk0LJGzXccoAAe7QJlROrsl0zulYqnRNxXVk
xY/y45/OCtR9/pnAryh68mxGxU23niSLmIHZu08PtUC8w0IicBlK/mlh/zO09t4l
Qr6a9o2i1Aj6ob1yrQMiTE7EbhJdLKuPsM0xDUsNDyF2j2wUSaxRg7P/S0PcbCdm
Ggan87t2d9Uuu0qS1RxcVtvPKwa17dnxUgXg6c6A7l3SYvhBOex5yJpE3ZVUghm/
YccbG3j4RSkfGRN02FTfaSvt7KzoZ/onZX3NKm+Esbn9z85JP8dWAHCsJekH/sue
BsVOT6VZR7VyKp4zU7I9fzoNJDeDHfpOJguqU1Jow5ccO3ryZ7Qup98HNWUlsGwJ
2cKCtxHLP8pFnQnK9f72X/3mWdhcozs3oY1cZI6TLCoEuULx1OfN4fm460YFc6YB
lgbMSADnR7xByv5gurP+AF5mveXPBzNS9XTHJr+jqRLLCiQmuMdAn7dwQ0/I6aAB
+OIsK3rn350RD6DpgOVzPUeQ+JP/Wd0Xf5yrWTVc+sJxWb179eF9hdLfdHJZ5XAm
1XfYUAlehPCBBFVLaFczjpt08LDHdvU1tq4QW3sPnNsd7Dv0rakQbmVnHmofRSqX
N/OQ+5zo59svqYRnDIiSmLJ3PvEJuEj7TGot8OkJrhnnJUDSUe4QreP8D27J9q71
0JGAdXFMy2uPnyaaNNOvr3VX6Q39Ax/6BhwREcRTyCHddHdAQxV9fNCmSDsKdeqz
PTqmxlwasI2yig+XQgJaxgUrxXGN6Qu5rzgvSSoNfpmfOzgXKhK81a1c7QgPXDpT
RS3dxo8FIxihKOMpSnBPFGsqnI+HgrPAytSjS1nniSvpCN4OMHsjRn7WSFHfwENM
+rRIjBKGP1YxqIrXFPfAd3Ly3UsSnzq6XvNGWY2ahoXczq1HIpDdAZb3QUroc9o0
/ggelUNwqkA/twl3EHfJ9DH+cVMO1HSJIe/LpoR0Iqv4VXyVFHq39QD0P6z+rDXG
/9J/K0YsZ4IjJ5MBBeShYz5xJghlPXPD4YpmaNLMYnW330DEAJZW9nXXISWPJvpV
SMh9d5RkNFkM69xLlobjamO7sai/iEEqbpE2WbT2h+6ACf1ObvE/kNM4CVvGVX4U
iulGPqHS2tMyNs3QP6Y7x1ASa2XGQbwNzrx/vr8LZFqehilIh8oCbaycCke0VmIk
2MO/JHUCLp1ui7SKlWeEwuNZBfwkrAIUFDpnskOGs6L065Adbzzj9vtWkJ+2gGk5
YKHEjRc5TI4cV5O4Ab7r6LQoNEMjpSm4CiUPsjp8mMjMGpnZnTj1Mve9c7ZS5W9y
V1DmBfcdeXkwHwpP13wjQurC/5U6deXWspl/QKXx8tWA/Ko/RVVSJ9e3snl8f+YE
GibTGW39pytiY4Vt7iy5bkdFdIp8y756SiNzDsxSWuvUpSyI+w8vH26M+vNRZVOJ
dXFDQgn77eXtTKtjpg6FO7eX/khEJslEAZTuPT4ibTI5A4Le3l89YNM2MI3ALx5W
zBgsmWu2PjVu2FLnKcbQbTCGCdgMhvEIov9MG75rzfU3DhtjuRPInkNoY5AhU6IO
SW/gf8SX8IkuudhsFoTLRCE0c7ThelVuI9OKLnOjiCSodawXRK1IDqQCN5SPLsy9
uvkoYDnpcz9rw4gKxaihRzQrTeR41w8K/oDFUICU8ZH72IFNUgSaqnUbd70gbDia
1D6sEZUaqPG/OmkukoATFyzjStAp26Y9oepG1vQE0sXDoN5RgsZAFKNWqG7NrtKc
I3tPiWdkVBMwn3pGkLmLWhuIfW87RO6zi1hLFN5AbaY/lrQRCME/gWRYTmwspNmn
hVCBD6Icen6865V0nMGTj7ENDSl/9hkat6LZVCA5rRkewiTREIyOn26KDyOLJ+f3
CuRGwbKeX4fICeeHCI1sXKL1/u1xVgtO0CvjZNDSHGDBBQYTgsNHdf42Csyxbc/o
lQ0JX08NQc145PvaDAxRkljL7ENl9rFydthKo8hqUlNXvWrFAz8/W5u5OAdtW8o/
y9DyvGmN4JtdpQYDFvttZfflasjspOmR0uHpyX0giBZwgq3d7oDhbx6elxWP8e4H
bA+ziNy4DC0269UkU37NfS/KMecQDedPh2SGyl6wyQtrRm7uUohSzbdQWrY6lycz
OiS3trRKp5M3ExmuurdjjTgfxNrpw1vZg+kMcROKVW9Ey/HmPhxIcHys0OgugQ2I
T/D1QyhL9843s+q75Tsfv+Z7SQimZZIKwAyZUmh4ukLeoRrnhmU6291H/oeVN6lI
/owT9HjHxzd2R2ffBczxrUJt1gmne0fbARZkjaUDmuYhxW+HbWU2Q1qKwMdI9xc1
pxAumyfEyq3qPU4Ep3cTROcDUcVhoM5+FSWuc4tjMwSVJHZBXR4PFbsI/JGtNBH9
5avIhZGEpbIo3hFfiP1XX4J3JqaiM8nnVWhFYgG2ZU25DkpB2y82aUUODoyEuWHh
XoROFAL30dlXPHuxjsxUFg0tWgPdzib7BcesNvYsrrdxjr0/bivLstO3AMfuBoFL
SFFhHqfXKXkxcX5sKcedpvz90gEkjYimo9hfPAhkR6f4s0IJUZBsyl0mjLp3hYH2
fOZQnGAYlfICQDCndbB/sVLYB0/gYH7hHcK60wLbuhDS9Hx/2mt0LTCOZHn7/dyi
h2Kk9tN4QisjciYc9oiWQN7lITrbtwa8XC2tX/FgGvQXXUCbSeKlrPaZmO838tFZ
h+6yErnp3ukC0yd0uIxFcb8RTXXV6I/88czQZe1oaNM9EGRD931CuuVQBiUHqshp
GaiszKQ1j1LyJ948TBxX5s/2kpxt/bCttrXbMLjOZqHlAT4KJeJmqThuEjBe/ibU
AJfceuWUEaoRdyHMNpT/7ujRyxQr+O+ii6BeZL37TvXnEAsz3Bshn6O3p+GjLnC3
nHLEgoWqD0NqtBFc7S3U2vmQAIUpV6IUDt/rWfq6FrpKig9IiDx5UtX0u++BBPTp
Dzk+cefhRstQfpuX3an9pNGvCOiXEl2stfzQvrn4W0RdIyajcfrJJ+/YNeFajqZf
iG/1wFGV9I8U+l3Bt7GXXB2ZVdSg6uVPQ570JJUJOIxK4OrLGZWoU9NW+NhcAKVC
+2J6ztpbI2eT2AM/Dsr6wipyIkcIJ0JpFb0WkewJlmEmnm5/uRaNf3MLXYFwx2s6
ZeGUN4x20gkwOD8SCJ9wxvios8BrWlzFEKt5P+8eDR+dSdFz22cDEKdicCuwGWRH
UOfDXPw+pmJ6Lz+pgY9qh4VCgg6yAfxNtREHybfiq2IXxblf8OhzY4UeYoNW3cBK
F1INCmjYE9xmGdlKmbCCgHU/l8rZsSAla7VQMZuYuKE=
`protect END_PROTECTED
