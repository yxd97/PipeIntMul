`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
icMM7+ux1WbOqh6/5wOUcoq+TfTqDySlmgsTBIXAxU+xPfyQe34vISR/gv4hJ5Oj
vLT3swexXaH/5WUTaWhwtVCm6cxayuRC05jigE6Jz4Msk0pGo/7JC75DTD3V2+29
uOMN4M6QxWowyjU212cCSsCeD6JGh1bLCHAlOr30lGd8IL0UPpmuv9jGUJ5leTMj
4J9rqaic6r51COTb1/blR6qU4eQOpXu6WVPhl04vIkWUk8rhOQ+Mf23xif2LxN0I
OSTbEeZ4he86YDIg8lSfs9rz/zhe3ICBe+5pINVJttugtCAhS4cz13r0LJTiyd8l
l61+/bIuT18tIYCP8wv6PhzONpILlT2cp37z1qFRHa0AkVSkE3/CoKlKkKNW8KtW
7Dr2JcUHmngImxHMSi2Ib35i6p58X+KLigOOEEcPBjnU14CtRGnRNkOzniB1u90g
XDTXX1g5isW2dbbcHGNiuO4GP9F29thhxXZk5kD9MSr/GXjzB9/2LsfekNIgk1Mx
BSBFyTqeBrf3vhjlDntSifDaF0pgi8FOjOgKjAuYSCQn4G9Dv1zVMF4USt+bNkY3
pRmXgUAZzdmug39EDPUamftohwroQfq28y4RYiJ1U54oOxSxfnkTiJE3cHPpkpdg
1tmb4R4EVdbgQEscv6KdSWA3v3qAZzzfQHbnYyUw6RU=
`protect END_PROTECTED
