`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2h4NL23QG0wdczbfTia6jk+7y+lkrDsENPqg8SnlfaATYHJEfjG2pcAZ/nIjv+XZ
53bfQFk+E0FPHDv73mR471EWqnHjGIy1Fq8+W3onwmj1hRXvAC44D7tqhOiWwRlu
bzKNQzIblPQrtaIrxEbQyCmCFkeHVtrq30ZA6Eih/p56gYEctnZ+ANVIYaDx0H6G
FUtiqox0FT+wpen88pE7oyEuLo3nPjyrrFQjUfG2LJTrmIaEpoEb773ce9QsWRHt
JBYM84/kfKGzKpXqGnNY6EKAJPYJoyBKxhoxUSDDry1iYMKrR3M86saLakdXWCiS
dR2UgCUN1Lee0rT6gUb3FxBN8qWyhWICzHFWjn4AKyoQLAcCUcUBJRrZb2Ivna+v
LmyC0fzyMZQ0wLlVcEyLApL+6QnVQ4yUrzvw0pB6mDs9P1HMTsMKX/Y8YuQONtza
F/uBxeKA3V4tk/bPyC1J9Oyr6PqHldDfsOGAn8adqOY9FxWkii4iBoVnM2VzTNee
crJR9ukUesxEiZt7KJdnlmNkiqZ17Bjp2335XIb57rLIlE2H1qzZ0YPPLJ2xnSmf
8K9d8AVxP2rgPQ9nXYoNTRouggux6PEyuzReSVl+CXcSppp/kEp/BNcIunqjJOCT
e5P8ZZRmxFe0jjzclGpO5toPfVAKxyeU1Wp1XNPhO70DjoCMCTIHyYmgqajqKO9z
CSg4jOMBQMOpUhtgNnHgCYrHd0nUKTkSl6dcPul05KUu8NiDCtJK8LPN5my0OA5R
1n3wcF6i7Xy0l9cWlA/eTUbmCv2wWKEbWA2Lw5v6bdqqUQtQUYhuH5dAJDPkYVai
CetGx2oUGrxu7HqZqlS/5H73S9b6XZRTiRr6Z8jp7AnMxTj95szOXi0KHYp49TXo
sSv1N4vPNY0AOOVxSjGaqZWARYZh8KeLb1fCgB5ATEekSM1DI3TYUiNVRO8Sgiv6
3Ff4k/LLmmhhRqQzXsVo/yK0znRkfXn4kAk0yQK/BbKdelZmbNFxrOm4wnkGwPmn
xOPD98j3aNBCfYINNk8UXR3Tukp8cSxmIZYielsryqYd7Cwtvb8sEhpVufGjHkyg
vmP5zDbQH6F5Cv+jHnrhTXtCkwN78/gBiDKphb3xtv0cqCYPcv0VQm/vHSULO8Ts
4wywd1ke24PRuEkoWxTRfTjtmTGauKoc3qLIiGPZLIKdJBqWK4ZIZkweRnfZlWJi
4QfEndYwFsM92Zu95M4IxMoBnH3XEOIxnf9nT7M8W5q3ZZYsaUqgfKXm9pTdrO6u
/nxVpJca+HLfKVpUCk4+Ktvsm1oQEBnpaqNB9i7/Vn0hrnSAdXs5tlSi+KbjDj/B
MXNBqohpgKLxLWQdAh9tfLXe46oiiWxr8EPe0N3ZB6JE81zJA9VtydE9bflC8gvH
+E7rVbxUkUpK81tzz/xPo2PkN//Y0O2qe0q48HyEwkNUq2jJcz21WeZYwvLVvmMI
a0wwDxojFv9bJM+DONsvcAn4EhiwDrqaomxFgOSlfAzMA6EGzz+W25ijmVC3oacq
+7756HVk6KAbwoKuETr1PgJSji8h9QlBJnE5iHf5UTTjFEX/3whV1DerKBj0krFm
aeA1vL46puO+2IjX+R4p5FrSGfATAzIAHvYk0UGav/BQkuy+8pRDxHKnXe9A2KBs
T+p+sJ00nJv+otpTNbRD0xqlLvMCfeLpHy41JbhD0vkPObAe8eBZebzZ0EVf0yu8
qm9jmTCtPRu0FQxcEgTu6Fylhw/aBA+5q36E/6UO4L9+d0YQBXJ+akOPjSwwSjx5
SI7QiXF/xSMrMeTn2M45eDF9431zizYvhk7y6Lemr4R5YCbeSBzd81JC4PnIg7BQ
FkVjN7U96kpUm+z/OPYvL7ruV8QsxuoRIv8myErEYUaELMcg9LF8uUyMnX0Q1CAz
GgRJ78K01jAGs8uR91e0LBrhUamxmBSnGYoRoXklkR1efRFtQc0p+WuXPh6zFtB0
GuX1d7KBgixWLDUVHx96ujQB9bRQ3qNx1hROvxV5WxOA246a+cUnBWKGJHXx/GG6
sVvsIqR9YKdpSTAXzIhFSPid/KfvOLMJfI3BCbxDNUdiFB0zx9Kxe+UuycVFeXP7
F+7aMo9XA0CiY/Te5apl5ouOIhb1cCLS55Iwbey7lYJ3QU3EYqvjyDHv2LJb+Ssx
EHUCtSkk7nSCTNV3AD4St0OJPy7/NA10CXiPgVMDRiSX4penkL3HYc6KVYTpYVdL
ENDW5YwsA+h7CcmDRz0tCxukxQX4k5dGybNAHn3RhFl2rAEflAevgQpQ6SFwfZys
/9fE9g3K51mKp4hFi7qWXaJZMlvtfUbVHyhpCejcWm3396lHX5p8ecUnZT5cgW/+
gTZ6y7OrMdAz+cAPYX320a3Q3bLpr+Pxtj12KgnfWjz6/72pLF+mKNSGG309UU/T
56KyYYnKLEuhU+aQjCYgqjWdTmlUWmrN808Jp9qHNNGjKccBrsHi8seEcQAYnBXB
BAI7aL9HEHGGl+n0oFfFHgGgaVB0VuNc1VyC+GlrkLWpmxqVY0695lYg/4M9RUji
+M9cBj4px4JTIHWicukIE+eT8bORR1B1UgjOBzj15lxivLkEnyvD5GmJoLjHwj1I
xFSqVVa9qDy72HHy7d17gcS01KewbR3ARsENigtfIzg9zj/7NGcqVgnLoIEjl2Xz
9ro+x+skaPBQ5XT4nrT9Vw==
`protect END_PROTECTED
