`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c6vf4lHUALKOoHwoWJiFyLiQNZJYzNSpk4PZSTZ7j3FdIn3VYd4TUa/yr4ggmLSe
pvnBiaPJKnrKu+IRW8AIdejBQ73VNH/yh6ugK9rWKWkTsdxTFVs9anNe42kBQnKi
jgSpmx2jbFuldWa9awJ7EtdfUxX3Wva17ZGOBnj9XNfA7N7HVsNyCuTmcIOHewL8
TpHfhZw+TFN1WuVFECyBDZHzhz6GwCPY3F9d49x6VqSL6y24CiXQzWpo7eJPG0P7
tM7Ti+I1+vn5qbc62uMhFiPH6n07jYvCf5qgDKGtqXieMpvA/qzCQchmqSAofM6J
Ach4c6e8gUcRDW7hfS0rjWUDjCaXFI4Ch6C6KzjSLUMN9z92MBrhNC7WqM5/V2uU
TrDvnk7WeERwP86xMKdawMWrLSKY9Gwuk0DCOZ1A3pib0nZKBm0PXO0/PN+OGlc/
DKVXWHY3I3kMx5q2nx5Z4w==
`protect END_PROTECTED
