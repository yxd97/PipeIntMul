`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kq+UXNGNPOTJp61wqjkrueww6j7yMjDXul3LCR345YJ5Ry3IJ8jB0WhpOPTcsp2p
fdVKQSMzOsK5F97JbU3h/tu2alrliyQqUMcI4RfbrXuCH/BWuImEUKMYLIN75lOk
i8f/OXEnV8F4lSX7w0k0hk5zU1DfraukN/GeEAgOoISR++kYf2ojeMEJ/gJHlqKJ
M4MKrximGxel0Z3ldjbxFu3Yn0VOWj6BGXbY879wEWavId33qtIxGSAPay2Iesuq
7BZV9xlJpio9yofySbYeJCg3HCRunL3hcfH6+njh5awnAnBdMePRLtQBX41LrtD8
gqio37DidZjYmVsI92vhkcugtH7SaavAWDqqbl7YvO9gC1Am9DZDn65+p5kJKJ6I
k0wWDMcDC+SCEZLT043ItaAlWHzYPr2vYj1eJOLHnzWIbEjvdfdBXc3W2k31kM1k
d9UCyGir0wd4sbsfieiIjvBB34hpucbKc1RnVdPcdL96bpMB+mFvvKrMLRSvroZX
p+CRQUy21DyKcf8hJM+ZOfbzjzJGLk2WZUhQ6LpupTObeG9U6xIFagwRKPnf865t
sseOwyq87cPX+6Eq/z/VPs5vTKJTaRZcRNdXrDiKzCirY7UCeG7RnZChBsist5Js
JisY+9oS422OKEOw2bAv+PGZ4czpFTTCaXucQMhwbcb8d6Gnnhb0cvXwzHvRqIyM
XaeyjKkgxu6BHweT2Jp3+Ri8Px05XDTs1BZ8TbOOvLPf/CEaPHNYD3UsBCIEAVE0
PC+NCjeIVTlOzqE8TiDa+CU6NwXdkain3m/XZcau7+3xcER0Pg08UfX9o9tUQfvF
6xxPwOD8F+TjhH4i/WSeMLtuZoX9W/5UyT2ik4r/jpSTaCTHnzISrBqk4Onx1gvg
a/fAGXdGmdd57xFcQeboOkYx1PnSMXH5h8U4mKkHPR9Vq+hMwUvj45jzx9X6rggN
AagBZ5A9Jpo+UTtkAbm+hlUx684xK7kd2XYxKRDO/fffGNBq2HvB7EBFn2G3xJ+Q
tayVSz35vcITwQjUwgdVhZn0l/I8q9bPfshMOmBB48gnAmyFOBCVKgyo2XaLZ7Pr
KJUABj2NwXObhJLpYMI/eLlanERnj8XkXjA+TRDOyk3bi+SWf+BSDXEZKiq4nYAe
sp+yNGLC0E33jbPMYDmYw67LSXAZ4Emi9ZmMV4Z7xut4wNlGGQDOcHNYzMUjkINL
GOoJlzoXj6Su9wyCs+BHYtrPXqDLG5Ob5G0HM2R4cxrZbLMubNDNzpFGYxJwo5PR
n+iBzRIPoQBc+cm6UezBMG7F76JJi+/T4V16y6cDCvVL1MmxJBGFlktSIXpe5TKc
LmxlaV/AgvSl1U5wIHxRuZKnrsr/iGLkTExS2fXtQWCqraRnU7S8M9UfroKBNgQw
UB7H04vNLTdccOxUKSFX8yeCHQPL986ngQQBLLk2S/CvelTY8Mg7XWwj+l8Lt0ZJ
w0qH4a0lwCBelTeQAMVjdIrhnQR7MqNRTgl1mnyYH+zUZtFOIaaSeCx1WHLSFBsl
4jlOpiql8BxeXsoeaAAxGAeCVY2EX1od+ecREzWRG2RBJ48lDXfDDawI9CyJ9Eyr
vJCIMGXZt6ZIYEWhZPXlsE48s2mTPxImZDvS0HaVYDE/xN8t/kjjmOGFuz3oUTZ1
oGQNIT3QtB3JU31Rk/Mg/fcrKt6wDD+AEs0x24NBtcFY1L7FSSmeht5Ls62PP9Oe
Qp8IjvrB5VbWmkCpjwGH+IMhLgmco/mWjwITTY0mwMOZQRtGFTg6gGduO6jqdghJ
BZd7ogQU/ri/NPWJaEutlw2a8dFPifdBXHuCgQu2CN1RWPsVXl7I52dG0RqV7ZnZ
155YE09KOmFqV0W6isYHfQXo/w7KKtColXpy6NeB454dVDhb9R0RK7E9BV7mJkJV
WgVxCyrMvwdxUw/F7szL5ga460JHz1a3pHYNVUas7pQMGTprm1ZjncTCaP6jyNsX
k8Qr0gbJQz/PQbV53r5R0Szo9MAn+0KoGQnASnVHUk7MJh92PKQP5l4qFGbu7/Yq
AdKPFHXIRIrFVRNzpJnDZlWA/AlI3N5y/JMr3jL+xZ2Rj/Jndp3BOJBKn4ICmvvx
JqNxCoeLH//C7S2pbR3wyhPq4PgHjrqy9mRVfkip8ULu5DwzAesOUeVgPtoCFqao
P+gknJiHIgY2/G9oSSODw9hbhWmP/+LkzxeqOw5NvU/cDlK3lXiNJpKBU5CQKsQY
ovtbtgBUPTPI8qPv6SHKKwc2ESIA8ImO10nsRuouNkohnAmXuDfdRY/w8ydxPYTl
aoy3y8C/g7ODAnjXrrYpTo+q2627NXxpO72C8B5bw8Em83xeAhMFYW7ZJjSU/ou6
7dncSBOMHBm8t6RwKC5+faI8S/SHxtRGQs6gkzyH0OQDvr1Wahgsyoh65znRG5K4
28z7/VY1K1K0AWZtqvMVMELeLD1ZWjEvNvM2dV+nJAwVrk5VQbZvExgQf9miY6x5
ZqZBUrIhPbkv0PLz/NSlxvZ82nsOzwVoP2sxKlL8qKULU2Qh/gzjGoIlhdks6FcA
8qXPuDt/c0R+xXCWKNlkxuiCm3jE33e+EnTGCBF+pztLz5u2kG78XLowaNYAilrf
Ci8ORcSw/H1ceyv9HBT/ePqpEZ2YtBM1+6QsoDZ3wy6romKWAXkTgzalB8n3gJkI
XMWnhCpZFnSBcwbarraP1g3DpEZDlyYQncgwCfnqrs02TP2p4sOCBh6e7UDSdhi4
xoc49AsqtI3p3IKLaRo/WFtjosUdD90L+NX3mNY83V1pBGWw2JNCobwwVX2YufE2
DRZRq3248dtK8SWTQAE0Jn0ZyruCeMlTYk5FfiZ95XOFVVDRoTqxdADbiwq1rHYS
2vCHP9JLzQMgz/as8bWaSBYaCk7q60Uv7yqKUVjS7RUh3K41fOi5pXBDu2p1d8OF
MTqN1ZAkr1HPoFc7lSzd9AgymuCmSm2FPMM5Uhbrz060eB4EoNCTtH6JkcE5ESKc
ZxdhiDOhS1yI+O2GgrK0uwtCWHf8El3f4qcjx4DDC6fF9IZKXeMF5ur+LNpHOp6y
LvfDrsI9ng/sGv8ACAey0BGyWE10mbPqX6ocklKTOhv4v3za5ChdXWWNj42y66Xh
SwN+te8oP+1GsiTFOXz6NU6XGWwA7KUF5owft3HAxq+vl8GlMj4CK2Hc5bIa3maQ
o0Gi7+d5vNlPjV8zfzMDecCJlDuKCQm9CIVPzqP8qjE5rBXxIGaPI06vhHqngeV1
83e2ZZzt5t2bEdY+knXa/VjeH02s0iZk6MHTC8zHPLGovIWOryjgcO8DDU9jfBty
C5nu+PZbw2ONsgaa7ZH0lYqICJn51Ri6UEetinCdTVcmur6YIIyi/yvQUJgx9a54
1TjJ4QVoiXHDp6ZqKXWeiNtc7SfICPg3fjgnnyYI/AQOjUOr6CC896lDROxC1onB
4cSAzitUzfY3QV5niKaCBsnA/veJE+ovAttgbvd9DPDRagpuHhVfRc424Lj3bPHb
/pCXxMgl2NCqywFAE6kcCckioriWZ8PZKR2FWJP4YymP4IjMx6VGUgsV8SzAM0Nw
AkzRJAMxz4y+hd7w6RT3bCCeLryi06jPd3Q01ZYuwBK2GTOj3AfvQacW41MEv1PG
t5o/NYX24wDIl8W8PxvNq/kFUqrH8mZAP8Jg5BbTphs7TQhjii3bMT4Y0twasQxz
iQfy7WY0YukCsRlwg9EFz05QT8k1z9EA9B4CI5BmZx1tnAe09w4SKKRrquzDnNWL
EnfP0FOYaiCLqGMTdpI23C9CDm3Dx/dE9m1jq4DtxRktZ80rfOs1VOOb3aA4JBME
Q3d5BCl+Iwp0PM5O5CciQ5HQloWuzaYUUx9YqpLhG/e1mcznXGfDbl2DuGBCFepS
79vPT58ynxLpQq8YvZh2KRO13/HLACuL5TFL7KmrGkmTCvcg4uxeOu05dezadJZY
RB0Mm9jv8DJEYUV3JIx9LWT+Emn08IxNI6tIIoLXFPYgXcR9mb0eC3yNFxydhKQ8
gJg2rAlZXpYZ0rmkCy650YMSga8Avfr6pLyJYarinDr2Binz2+ctiLJaVY3Fbn/j
CiUjNQvv2sst7Wd5ePzSd/YJFlo11usCD01nSZuk1NKIgpuMhiCOMPs6YQq7miq2
1Kb03HwXqr3inJ0Aaq08/vaLMTkS+/ZnYTK08X+X1Opn+WivXrVTQu8HvgGINvvo
0bLish6LDWy8pdzTdDUOkJTrmGIGrXkKNlIl8Mf8ZdImE6n/DoBmjmvbU++ON30d
s/NtW6W3Oxw86ZoVQeyAdfZ3mO3p+85PatZ82Df5HaIxL1nG//9Hbl54rEjJ5bDs
Ywp5ZTiUFx1jkwDgYZ7oFcPS0l4u65MRL+ejBGVJE2ttQTBXZPoXb9uDKM1Xg6xu
jlKlpJr541fLdbD/W5S1LWvSUyRanU5y+qqCZX4Y6dzfqFNdh46FCmkJ6ZOLZug3
CR2PHmRu+FXTVRN3gdws7mmUGg5xPll1ApjjBcTNmJDzgBBv8em3qpKOXbTLX2k7
JtkUiI7PWONWGHn9MUej1GhMsxhXSF5vangl6muCkP3eVCBmELcq4Om+NYdL4/i3
Y/MzweySTrIptHlwXvbc95LySsSCcrQgG+i6wOJjyzwIBhakpnvJEWuA7IcCHJAk
mNR+WwA5pxTMjX4Ad5T3/oGBNffc9EEhQwES9dLPdpQQvUR2cacQNjaI8tjenj1F
R90Womjfb0PH6nnJus4bRvszOW+YCO7j3N04kwf/1OjOeQR2l3rKB9xooe/nPzbU
fqBgUcibjwqBXh2SnEIcjy54Jzkm0ARlQ0IaNH27qRf7MML0mwquJ4mqL1EgbZWq
1gn5k/3hDpFxkxcwvmPB6fdEIVMZFVCH4cB2eoXMOj5x2jNc4nUuXg+rH3ZqPnDz
iUtoBzIZYIRYzZD9Mj/lu5pteMzxNgp5w7sWvx5wQs56JcTueUxePK8xWaTubnSX
9PE/hXmoBYlbCD9tVNWoDRG9RxU2+XIPf1PhgTjTLE/jYKRlFDYzzATobiwhozKx
Q3CSr2LuYbRHwDa2CSQmA1GkjljPQNjf3OmnFHf9f4VOnBYto7o2nHlZM3eiwx2O
gkTJnnCwpRmKwEN2swgP6euZ9bcHhY9xE0eQdC2Wq+f0UPwFixCS6yBuKa+pH/Nc
uA6sjnV/or1JIRlGK24MEn5GEb7AEX41rDjTOGJzujSnEzhIIddAW0Yzykw0qgjm
SVeULTsK2hA+KhqaY8uvJ59sdw7TKESMOSgfJ59oBvjwEE2tKjybi955VVvG/YyS
xMeCMBwWvxcnIt03wG9Cr60/zXVKc4kR7BjN8FdqdStTxXBFCWcpkDOMOA2yX1wD
isRwnS0IqMqt/8xxRUzUFez1nkqelTxhIX9kIu+3oYnnqKKxsHToJmtokpti7Qz7
LARpi2SFzYaX3Hgj4BzGVHo27Q/jL5fBAlBQXRl23urD4LKUeg29/+RU0lxdYyux
Et8KyoWf7Ycb3DjiOXXKdEtqnZZwtXTg2G5LMy1BEizgm2OhWwhT1wKKn1q2jt2d
NL6VR+2Rh+d946+cJeHiIYkAAYyVN3+jS8hEp6ERhUJOLvr6t4NkWgWhrk3kbwd7
38n5kXV8+m6bGSxUaKYzLtO+v0vcJTH+h0+aK6qJtNgx93E8vgQwzX5gVQ5h2bzs
tVOwg//rafDNzr7D6BcZOnReqwmW9nEA3SXKvCrbGMmUTvUMZHW0pBono5uJrEXt
IAZu64d7woqb1xyRuqJ6KAjo9DqvW0JaY/Vq9CML5kzEXsOImHA2nYbM/p/QCBbv
6a8GpvH6mr+Nz+HNKPosFs+LkyUN2hxZQFa3AHSF64G6s4pcowoXxCVYQ55+4ZWd
jmxKwjAt/7DHuSq5S7WE3/6SPVSgPQpLkM20srLiTHQzx0sdSnVZFqJYo0jpaAuA
pgYqBYnHoKJlu6Fmjn0SQueNmlNfkcA5OsmWbTMxP4fdpsYGyLBy98PwtPue3vqG
ZVEE+0y7j0TZtj+lcRCuxbsiqwdEg/VDKQ5oBoKWo2wCYYrCIGLbhW0z1YgPgFyC
IIlnf/ZUvxT4BpBAsfT4g98g9aohMcThyy++zYm6oa198UV/hQX+DPJYjsZjgdjk
k3k+T/3zNjcUblgYORUMonwpK3PALY+owvsy8jxiDECyxZ+lBPDTGgCn9Uv/149m
6R9PQPw+c3Um4naoOEt8psjyI2Y9h++UxKcoIpgQ1bhU8ORpNAU7wO4uXtKNFxTu
6d5KAa6AkX1jDzA1msdF+JTwv19wVXinfHwgQ9is2061rQlxLr7vN1oUyYcKuCFS
vtJ+M5QkYPmD60StfSCL6hingfnN/kKgJT53F6nP7kwxAObQyHAaE2W5GVptePhe
lnId28e87FqMQv5g4CXAgCayDxQmlL/PW+Z4qExuOulzGZvFAZbxLn1fOUKmRR8Q
cxsl5ucIMqQNJVhVNzyS0CPdTt6RT/Qarj4Y+TlorzCMItkKs69/QdWZTDuT+O+V
dQU0o/fufW8kpTXpEx89u6Vj8TqGVTYJOV1/A1kS6lL4K/r4uw8z09k4hLRqLdHy
LLsijh5EVKESHDKhx3XwYPUJUnfG70r1IUtKS1Je8Z4E33wmAm+clQUq7iNm8ldp
+bIyvo1yU+ckyx6bJqAmNS6n2tUL5gGqpy7ZvA/0MdxXMKRcJGFqv7NggWYgwJ0V
sC5M2S30gk3xuRqGG41f5hfrdW0kFxAmT9kaJjrcG9VNyQ8U7HVx7zSVQhByGSLU
L0E+WnYH4SUa9vybEpq9Vh+vp7h/4TbmDHJhxguP7UdYQLcZ4u93VEqLYKRpgP1W
SECSXIqHyKigec63+uidpyMS7YMrC3a4+rJAycvbYN4lJd0Rf+AVvWWUH0TuWI6z
jwZ2ah84ezTVrlot4vNsil9lf3UsEjT+xZhwzHzzqcfTzv14WHZUaZbCnhYo1xl7
JGmIlqKv+Wkv+o5yaIUFvqR5m21wZnPlBSNC4fVQFGcy7E2D6VygRQEK6Og9ji9/
5uBi8rmffa12C9rNp9lPqXW9HL+sjq1fuEtDFBPiv0b6CjQA/xlf273oU/izkxzs
NFK4p8h/bVnDMA+WUxAfPc+2zIXDf3Drx1v7Sni64D53hhU1QrpmOBn3agXG82g5
B+vgal6vXr1B6Ld7XM7m+wECaQGK8w5BOc72pvtc7R/5nSJ+zC73TA4hV/SggJQI
QqWdQXtdvakY0kFm7p8YA/LBW67E92vMhjlUI5wv2KcgacCLUmOlVb8nVtlG3lAH
uiSkUHbxr2FHHW367VIZePTDLBMDzdVmGw2EHZODiWTpFYNTNyaSljgyyZ3ip5v9
QesV9V3QpVh7LYlFojT6dwAfaeo/c0HglvdNEcHCL5+yvjo3aOaz7kaaTNwkUVuV
A0AfUeEmKa8zpD5Aisp4e/BZjfuJg+NHiT+byUjO2qEwQW42OWcBVp7J4iSUVTlX
2OxBCimuT/l5hogOYF+t+1jRsbsQ5WXTLXMAs719fsIGo0HyhZz/2Y6RfW9AZCLS
yizahAOEFo1SznQ5Xu8qw39EuVvYVmaNGzuIs3/4m4Tp8i72ryWgI2DWh5Z4WqQw
YNlWKYw896g+SwYrh2Z4Z5dw8VbfjXsc8Oy6/qZzb8EWlocDgYqcpBjXw9h9mZxZ
epnw8lNQ+Ej7yibBi7XAsHIoe/03DYWki1/kF5s6HK6TLPTHO4CH6LLf4GsI+IIe
plY2U/9hjrAbiVp04KZVqq4fBUBUrcywszPF23209jS2E73nQwFdv3lGLpQ9TpJx
MOiFemd4oWCZyD1xe4iHKFWalyZYxr1o6sC7CPC0UVSivKLlydosSuGT/IqtSLzz
OFjjDUIftaUiahLmJhAD7WcZ101xuIVzmVcvKGaCe243ZIqEnhnnTxRQylBwO4/P
o0lQOW9JaiZzq1heQDww7i3m3l5yVqfRRipb0WRZwwzC6Mb55ttdelnvN8Sx6i+K
Dyz4txQc9GlJZN/obkyaJ/OQ391FurJTaU/PxvzXnh171KQMADicqLWALQ3JUXiH
H9tBTYrlZHcc5ATKP9bGgRoHIWn7Kzv/HfhjLUu/2Wtvr4AJ1HmZ5rjln2OTZGtT
3TI9AjJ+d+2OP1ThRpgiscHzrUEyCtZKtvs8URSHJib+D7TSJPfIylCYmXj7U36H
5O/wM7d2aTBcrSdETwjGyGGhm2cacakQ+y4PW1E194dH8geJjnm374/jnFzbGJu1
qZWbOxbJgQu6/7EnyGLVHeDi2Qnwa9b+x1G9jAkb1ZMND52RFdTUaXL/FYBGpJSd
Jws1dg2+imooXqwjPeL1rhUYo2ZeQv08wYpiYMid9ho=
`protect END_PROTECTED
