`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zLU8Hi7jg65eqe4qmlpp8GeztafE8IjerEPSKl+GSNz+EMISQCnxiicfDms1MBc7
eWVgGt6RJn8z1G67yAvrTy5SqGOw0JG/eTCSwTBdVbYgOGPD5VF540ZmXTjh+D91
fPbwl/KhSonWD9ucT+Mp5LyFrea3pLT4tbwT5QdiRQ3l+vCy5VuyMQ9ilntwBZaD
BcolGKmaBv7vjhs18I5SapeGJwISINwlttup0DArINa3KRG8pL/NcN9R5BO2+lxc
+T/VYb8vbAuwHZq46RHgxH2HGRGX90HTTW0ANXw9a1jS4M2bQ0l9SGfKMa9W6TPO
HJhRNJdwVHsyjap4oFPNcQ==
`protect END_PROTECTED
