`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ESTyWs96uQzaHGfV+K8Ea29+F2f6AnMhTFOigXyvIDDdiL1cWnBJRDmfKBdUfm3Z
+GEB4w/hFOiGO35q8jxkfk/aPbZzSFJzIieVbr5cw2lxAV3pI9KIoLiGKZD4A+2Z
BvGwpKGDXW53kfQ7g1VL+E7pjEjn/UWXqDHUU7nZo6wrEF3eNBqvgfwNq7i6ftY7
bqIEuZmKtaZTXCpCaHTmN/AsJOJ644Uf+8PcCReX5ZOfnXfcN8Xi38VzafiEaewC
yMys1jzHCIneBHazG/qC5f+41ORj+XgCS6M+AoeeYF+/J7JVYQ0yh58NQ7SaP258
mCkblpTrfNdzf+DgdZuVwUcCvPICiEktZZvLRWUdxVjiw8ZF8wK2I2Kwid2I6/hL
FTSVa88pvVym2jiq4TGOWcxjhaFrcAG+NVxj0vOoMGdGN+C45Fp/1zBsIrF0MUmH
Fzj3su2nxROm3PLYHE8M9gV0Y1JWvetudoc+XdTLf80/qmOHABVKRNYOrLZasddF
oCI6Beba+x4p01irqBt6RcbYbpQzIiQ6M+/wB0uTpIY=
`protect END_PROTECTED
