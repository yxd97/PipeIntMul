`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aHVt5ZIqF8ymbBYAeTaAV1wDlIU1j55wFI63gUO4TaKTM0ABW7Ec+JDuZsJyVdbQ
FIabAsMaNKRAhi4g+TnM+qkwNEnnjPpOqF7cTW39ol/Y/OKkNTxS893d447xodrW
Zdok3+vp5HDjcEJ8dOdpcophzb/WPtzd1bmbs4EEGpb7bA1BuvgMhcEe/YK+ydTS
2wQE7aEy7MY5IQSTh7roWJ4gtfuXiahrCiwjqK5kVtSY0UPUuRxAwixr5SmoA+VU
GyCl0oKfMfcFQYJXP4ccLCZ0u4RCpWSRJQCY94/lXcK7Qd8WGqgdfncbXHOAx4Vl
0jIYSU2VnWo8595PPjVQiabgLIxuaDGz8txgxy2mFiuqqdc5WGm0WR9OAQZalSA2
DzqlJ8SkAycwWDVKC3xMAQ9wY5RruxkYUQGh1c+jbeJWCA9p+zRzasJKoKPDUx4A
/RyqlZKKXyxgrYZ+4BMtGTZd/fTMhH+LePrGBHgATGmZ1I6IrRsyerFP0zaimo9T
qKrSon8fyP1Fy6NbhJS8LQmAc3kW8JDq9wknEQQ0B1ke1XDq1BklGr3Kxx7oG+Pv
GGl6sp6HGQIUmo6Cn8es5gROwm2LbmARraQcWlffQbyG3bz409E3tUioSgZiTDoq
S1+bKjl6c8I36ZULh4q/jAT9HqCDEtuHxhAlX1vz94oMSnrsGgd4TtOYVCWpXWH7
vW1g9X+UyFr1d/4CCFx+fn/qr90EdD1ebbCCTcSyMoCiaXSO5I/kCFUAA2cINS/F
fY9ePB74EW1Q9AH0j4D4Fxfp0WQAXxdmL5Baehcj8Q5iJtJxYEyiPwj/G44QjDvb
J0hNqHUoQ8x+AQH9Xk931KpayYN1FXOXZHndiFRtEOBbQNtMGd3DnSqQtb7wkfAy
MjFs3KHW1jy8X7lp9eare6NPYTxCsnquljPFPEd5Yr6/6PxkTye92FHRb4NN2LSZ
`protect END_PROTECTED
