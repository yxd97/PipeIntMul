`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bxDd29QDF8oewonp1/Suyk5cnNnF+yIP0qVKGMSpcZ7bg3BLvSaFi4PAuEkDP+RX
6GHYFVu+8yQ7loxE1QmITd+3rlzvLD4AjxR4lDOcByDMhuptUI4Lr6kK5cRf2I+a
TSJq9MIyaIPH2QhHXCxQ02+txn/jnDKe63QGkrliUHQdFmpvY97LXm1Sf2CFXWZe
mndhaSGbXdlAPDLArmv0Nd9xKOv3/HPzHg1pEa7qfjWUxY4EDidH+6DbqkOpazWz
ojwcIDUStwYaF5J++w4BIE9A5aHn2G9CkRb0JYpJyXgm6EayadK0nRXxwoi0RGiD
IMxq7TzbtQK1CiEThFY3YoJ1SBYiKuLJ0HKW7DybqVPMzAe7/ZyjKn1iGwDYo0c8
Dzm8iBuZerFnkPlF2xKlw1XkAm69FjkoDkiiDBYA/dg=
`protect END_PROTECTED
