`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fGGINSHM30AHKpDj8kNnfzIQhpGzkxR7Zl6XebM+wyhcigZRTykU9gIH0lmeGQMT
LZuIrqPGN91p7oyNHYL+y4Cv2MXXusIYTxTjjezRp49lqAzhLZapLM9D74+atFUg
ANQOi5sLWHFTMLIKV0n8ydZ/9r5SOaHHCUO8SEe4Ue8vvlKIfh/8xa6zXGDsBPYL
IpcXYYzqwkMWjON6w1FqwjTtCvYhlmg4G+0q0jChggJpK/2MWZhfliez2mNnJfGC
FlQZLfn8x7BHScHnBhTcHDuskJ0sgtpQRviIy6y6bNcOA6fIiWHZYq+Q8/k1DmFp
c1I124b2jzAthZRaJdknHzxOlVE6BmjurjpvQ/3iQhlPUf15hVkFslXeMJ94FiXH
XuA+vxT2nkSQ3681r2N65w==
`protect END_PROTECTED
