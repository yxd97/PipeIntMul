`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0w2myrtG3ZytF/gejVupmhtMk5excD9wNTK2AOrIKZmfKdP9xMle4WGmaLF0egD/
U/M078tDBfbZSW1EcrlqmHPrqcW3FbFBhdjP3pQelB2BiBzLwitiJ6huCuEvxjIO
fZppc8d8+K8hkRsc3epTzxVJlgeRdgbdlJWG3pM1LLVp3PaI1tg4tDQv3QMoAR3x
eLcl0wwQtF4oKHWq64LMfzk5allfz3e3asS+JXZVpMqbSPeVmZ0MLCO2WCALB+iN
tra+7ROJsqvyXsiChY4KcsGkcwwxwOacsrAl0Xfv6L9pI5sFgxRiLPtQ7Jdka3IY
MlBPSe6n3WvkZZUQMP9CfPl6ya5sds/ne/61Psvjn6g4tiMo+J1QTw2N9CeTIUEb
8YOk0VHUveZkEMuJ7BOc1coksniW8+XimfLNgOlDiTFWNfX6zXsUsvFMisucXrwI
BeiEdeamDAVBKCkoyK8Bl70Txgmbvj3nZbMf8XsVmdJpIDYbxg9T+1l+1Tzps+5L
2f52N9IDlGlTegOJnK7mYpVz7IZM9h8XILDrZrqYCUkor1J6NWGIkBlMoj7FmbaL
YoMjs01RrhrgpEqZ1D1/FNyWwquQjeqEhU1G8excAcHk0Mz8UjEtbS7dCW+YXRYr
3SpO7Yon8Aq6oSW71XW99G2GQlkIg4WTTZCz48Duz51Wj12fCKCPt0JMxxMNVMlh
yWpmhOXqjxpyPvOJ2ojtOg6easRoWQ2UQWVwEbSUbim/Cl7Z0nyi51JDNLdJ50fA
lHEot4uIJgEf649JJb3R35z6XLch8DdncOLSeb+5eGpqsuc6DoZ4yB5+89dO93zJ
S2sXj5NbP428EGmYwToWXx9AOHoZhooKcgjus5QHkJ3ScOk2KMUL1B22kRh/Twu3
GgwG/qn8GKBMOdb7jx8yIQ==
`protect END_PROTECTED
