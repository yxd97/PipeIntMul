`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iafcmb2aavuCTLk1J5JXq5sKDMzhh3WMPE9y0xib0ypDHvvHPA+O5xXKH4eYbB3n
do7qTKo/QSsxx+U/eP/c2O4/yYt8D+Rbdts/XZt/58BSXAIvzyTvPrl8qAAkwjNI
9a8HW+6LfYYa5k2wxWxi39EvaBG1S9Qk8a2lHhK8TLUxXsfgVjOrTMd8InCFfyaS
Y9sdZm9LRsxQ3TpEJaGwdF7AjmFwzKRjVLBu7khUs3NaHa52s1KorxCFXqnfWymH
uA04XeRwIlfKTdcHuPANGEY16DClRnqvN6m6Tfo9QNkY0/RG83Xft4NCCWCiw5rU
s/Jpq6d+8py5E8jl9p/vZA==
`protect END_PROTECTED
