`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
irRXoBv9QmOJibfg400wTLuSkxtGVdchcnGD+vhGC4Ezj8g+sHQ2DxjSYTowz3QV
LthjI8YO6wAoKqkiopJG9JglNI6ylkVxIqMpEu4FuD6dU75s8pFJlcrh1LfhBa4z
Z/5VOUvqjsClx3CJwNxfj3mghLh6TlCXRg4uc2Y8LnSb/jhuL95/ei8mYoxIItGt
kYC2RejeEv557EalEw1L6pmShRjFvRaT4avEdv7eI3YWlVZSjSO9+1Wp4iGL76uM
G9e2fjmyJjCrWrLxOGLhz7jRTF1I+70k9AHfjvWUGE+xs8TSnbECuOLLKLz9tg1X
jfPDXqL76z5xBsyDzqsvCJr32TnUgQSM2bpGrMxMFwPiYPlM/ABGtp2YjD5FzGMQ
fXX2BSfizADviJ1eDctYeHEJpr8OemAo9IZS6rLjdQEgexABSXlbwCQGKdeKYKmN
IjpFmThYjO4pbDJKQriciE/lDfk+z2S3un+zto06rXEaQn0czMlsQggT20mtvd0W
K4OIRJOD8+4Uce+bSTBJ1sj6/4Vu2E/Ptm72wAg0AVOo73oJM4O2JS3P5NqHO/AG
FlRd7EjcUOn8Vyr2348n+6LpYuPs/S7cPEMDLgvqzdbDEJ+V4hh1TfifREoZYBD3
mW3DszefwUPJPSGvAZz4cjdmnaLsPEd5D2ayf7DuuDqgmxzssQDBI05llXcf7Nvz
LLBxSOSnmC3Qn5MPWxkGAV6C21oZx6S+NHpOJvnOwWOchOCVwCjU11n251Me2oLy
`protect END_PROTECTED
