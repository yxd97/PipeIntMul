`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KUrvMflzdMdhQ5zVklT4ebU+FLyf5jq/xvBLkg9+UaHxAK8vkz+wySdx7sy5kMZo
v2cSFW/XxoqOIAatqlQwGM0u9GZGpvNzBuszge/EWnVBcarEGrjyOYBOHv2IaCvn
vhqpVQnNBPMR4ZIZRnZwSZg3kD93Ud2Bf/qw6YJ8evRaq5Fw4vYifCed2Q2o1Ec5
7KLxbWbFN6tyds8usLtRlfdZWKzfenltzA/5FjTaK8cF90eP6pCmUh45I0njT3SO
5hMLcpmLosEmHprazvSlKQ==
`protect END_PROTECTED
