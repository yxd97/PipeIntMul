`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qWOMxsNLKvQ5et9jGQu/QbkHcYa9tVt1C+HNUj9ajlaHd3JLYmA+HnHdfVwdtDT3
iAXH2MeYXJ2rinyd7/XE7XE32MtUJWF7/Dzy1WEILg4mAw+af5+inhkNz9dhv4G/
ai1VyXUCl60dOKNXeavvEQfQTNv7KhjGc40EhewOZhsjr2BDWtrdJxrfYyDo0JrM
VXicNOuUL+QUGy/lYeuX1XEOPVUCZNCGF65rYvbmMXmz0yy/HnTHXzwlY08RD/wJ
KQpHAail032yMrR2GLYgzByvy32PhSHDzTziK7tP1nIOrcU9HL66WsQw32bRLaG9
7cytqb42q05mnvmrUJ/eSUMnzjAgONg90LDh+RM6hfQdhKDOOPgvTAHAY/I3uWod
TijFW1HkyDrW4ySchCoY/4jEhUNXMpdYBgn4CzLixZVLjVU2NFhsyIRRzajjbS8a
`protect END_PROTECTED
