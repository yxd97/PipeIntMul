`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvqLhsJZDQAfoGSZPFi/AGPd1qrAPE8/aQAP4Obsj4epUv9WnLHu8o1GE7zUiHKV
Acru035wSlg5S2cSitcuw2rr/8+2CjoLPR7V3bRwMcgSTHx7Y5ITg2q3+sQwJtj2
lQnNuwSI8XEfofahwj21wOIaj8v0Xt1gN+2kDVmWaSsj/zHxjwJdvjSaoYPLI9+/
k23wIYqjOMtr/SHjOqg/eIAgzNiOof9IRmxsB9S+KVuyh9+vkdhikLNx2llmDxdw
CiRA3F3ZXfgpKugTC3MBh58kGBXo9p93aQFBbE4kJfrLdUesRzV0l9lvF2M67E85
LQRgXCwRw02ELShsGFem9M7Mh/BKPkRdeDhEvhkb149G9POCxhNwidAFuf+Txmr/
67ByDHpEdpQs8WZGRkhVXk3IqXE6Byr+cKHN88XWR+8zY9/eE440J6TLcsBz7YwR
o8WTDNYswzWHFm9+EOApe/BP3tQm7p1M931xuX3eDDVjdlJuUARgiGAfR6wJDnGF
3XELxdNqgurT48qwK5T0XQGH3YOrmNcakeZLJX6Pw13r2lZ/pmUnA4MtKK2WI2Bl
EQIZtGg360+LhZG2VjqsVq+WfyAEAQ+uLnkIUHuOIuMlVmWaxtfbTW+52csFJIb+
T9aeAExAax5WXQdvEqD1z+wm7WUkdrdVBIwmvV1K9BAjYKGulUxHNMgqHqknO+L2
`protect END_PROTECTED
