`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UHlv6wmsahEbLgZT1ftFiV/lBlxTPzWkhJtOiKYfHe9ZALBLpkbKGC1UAUtqRJef
Ki6yKNCQQuz78+qulCSQ47U/gfe+kXv5JU1i4ZYRrwqv7gvnl9pWaKAYWgEgb94Q
Os32PCQvoLa1ymrJOhM8eQK3Z/nAL6rlnBScOh81+mY5855I4wIZzxLvGI6zdfk8
W7aqW/rlXnUYWpDdRRYLeat6jkBqWEnfmMXnOKh6A894M+f4cb/rzlyfSrgQ8vDz
g5Vq5mTvZC7XchiT41R6Oqr4Iz0tb4GBVB0Cw1BADv0V0IjZuk1QcIFtDRh9gBIZ
7xBhEedAjvrN0959NmoiQTZotIEfBqffdFChq9IUhUn/FH6sAY8SSrsoHhmOGTaW
36FZebz9qGUKmAKhynDvPbfoYjCMQdvG80rRu+eNZa/k5fVwly9sc4+IX1drNK2i
qyqYEC8ZTd630PYcWA03b4HQZy1jW6I2zC8A9CPnLnIoZsjJaAQoLk+zbfWWv8ba
`protect END_PROTECTED
