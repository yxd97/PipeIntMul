library verilog;
use verilog.vl_types.all;
entity BUF is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end BUF;
