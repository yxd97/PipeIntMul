`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cfN7/kfy66mnY4G32duuVPT1vPGpYwjJ+W5k1Jmx9MITXwD8sJ0CVVQWBpoiwBxI
PT6T5BVfevg1rHYSF58Z/j/St8ZqnsWZBwbaknDbaJqd+UOZfXAVBBQcxl4xUCFL
bsZkLCimGVz1erurjPs/36R2wqwxTphNlChe4yW9Vvm75zSYoVgy83RMqHsOCHkZ
W7yhzKPdBrh0pvWCKYxhUaSxMQ25mjl0DtS/3uku0WxoX3tR3nM06M5m4QltTz0Z
mc3vTxqoeyEhoBbg8dbBe4q+YX6Iig6gBZZGEfw1QxXz0Fe0rNvE3TWFRLq/nm/4
DIhlcIbFNKlGj+50J5Zf6xlqApTTpmqxXupz1z2IfWQ8Sjh9Y5hqOT+QsayA1Kn7
a1l5Nu+0Mku3Nzxz8NLbyk65EynD/+arzEQtYZEKk7Nu7pWDxkhPSyHAG+IAosca
5TU8Fzp7DV3qxDsetFqvawrAtmo4mGrCaI/9QGApPj5ZuwefoFwG4SVBjjeOGLRB
wX+HhQoRexkhdItBnw5AyuPzqJE1V2v/RxFMZtGunWymBPPLBQSP7AcF7itoSbzn
KNOrWjm9EbGRxTQBzpq1/Ww+yIHb1NLNnQxhsp9itjKXxRdT35FVJCDOjc5P8oLK
1Tt5WhyK8cuuM8ac0+OpsZVn6EzLlqmMRTEBsWCX0oLYyUjdza9onu7o+Jxeamlz
sgtiaOpIsjHHLeiIpJLY7xcMjU2iGF8RViKkuSWhZD7SH8H+ZnwVF2cwMcyT3lT5
SqvOEOCG1f0s4HJHZmfGKPQx9aBZEdIhyYtUjMXHq6kimX6fUWuzd7p6KYOozOtH
9MOzWQGZkkyik+EmTVvxSTesU95J+xzPW2SenJ6SNOOsj2W36XtdkUl+wEtMvyj5
Oz+gLEj306GD7/4F/vTzHOIR7P4/hWm49+6vgtj8MiD8CG0BGqgW8EBUSh4kRJUj
oB/Q6obxBCEPVw6Lz7rnKwqRfjCUxU2zCrc7hISe0Pg1ih7+DeEJn2Nxo5+Bgya0
eCPaGJW6E+9kXxBe2NGnLYe+u/W/HKbTy2j/m8Sy2H8rT1W1uqGv6NqMgU6Jqifr
kv1jSLJUviwNMP2TYxOhoVjqvhNKvuVL4qbUJF4URJikdOHBRfuII8HI0M6ILDxu
ln0A925RlZssJ7iInmrh3rbGnL4HsgsPH2FcNbkxf8PbaNYaQDyR6hFvRIUGodTr
Wmg+GCGtVQluTfLA+v0cwrHu7t0ugqJPPhrVOvFK94IzwoGH/OnuZL3QmYgAf1rv
/xFLtR8GhgHHOdQY2iHYpubuVyYCEQ70KFwfA0PZZ5jguCZXeceeru48FemmyELz
Ga3psBxAlGJIsWBQ/ax36WM6FBWy3cC8xl94pNDd3A9IAVMl6GZXVwvQs1ziEkLm
SvM/42Bt8D5PgjIOlPvS4PTrxGq3f6Xda+Pfgt9vsdFAdytBCUnDF/WVlOlN4ScI
9S8LoEAG53WxcRANuSv6hmHTsg+yq2URbs/szZYDkJXXUTbfiEX91rjNJYdz8sAU
2EdHNtYK4ZjOkOd+o6K2dODPMNk639wBeeh8AcmOPv8J0kgNVJE3qX8mVKq2m+Fl
yF+tRUQ7QlbdZxw/n9IaQzBZ9czDAqDSoysjUHs1hOqIK6v+9mV1Ev/3Oh/sNmsI
vQLpuO4IDBh//stg6bhiYrPnv0nD7mqMkXDUWjddAQemiDTJpk+ItsKP3q0Kydmt
PGopZNVU/hDXuqXCg8CQ2GBNqDZWsNlDLEv2qsChTGYsbstS8nDuQrwdIYDi/qlp
OxkHOVxH+EwoUt+ODHehKMh3L4pcXXuM96qCfPmgvT9NYY2+sZ04qpkJaRPb7RqB
2KCPTT1BxEGNyR45Pmrc/TUQvGCMH7gJc/ShlFbpjXSrnFF5UGCeWBly76JMwHJi
92tw2GABcaGT+k2Uwp5TSJ4RwBs1Sv/9ySd7/ywmxm4oXpN6IcgECKM7SyhbNbU6
9eTiZvDKAHLxonDZazMx9OElkGdfoG4aPLv4URTFXIfNKg5P14ombzA68ArGdst+
DI54Up7NtsJwI5dZv4lMJvdXN5j30ZNkXZP7OCRXm9ydAFvghZN5wS4wqOsmNMtF
s9uwJbU+bxyDTMyhCm7r+OnYy11xNfQtKYJ8HEAGJ8PHPVYdMqt9pnC0vtgW9/av
oTHw0e8zHNfui9WxHT8bZ3g+4+Zor3enqMasNQiY/rjsao1BvY54QK+hl376oODF
WUs5shL1d6X77BhT//qcE/wQEzY9HTjYyNMNCb/rK7ib1IFbdYFvne/IqdEejjkN
q36Xc2+eDu7OR6QYN3+8VnBoraU/jLNKVlqxfK8XzlWhK19MvXDdLLViKebDL+FS
GeIhBeQFQh0vLIqXIfn7QDKBqnN69/Ca9YLKgcizssExLEr+b65iimyLwu5zB00J
voAsgfT9uS3zs9JmpOiC4nUTZ7eYOQHH6L46C1nHuYiKA3hGh03q8vikktSPGbJh
JVgwmKxiQx2BqKhYdkw6JQ4F827MERaDNd0jCUW9yrkeyyfxTbO2sYUE07NW2QdX
PZmpJQzyQy9VSp2UgC1hFtkt1NBXoSPH0ZkcpRM9bW9jVmFXA2OtU4aDhLwimKl7
bllBpx3ILL8y8sPMjIS0sv4OkMm07m7nE9b8uj5bt9eDHb/Qb2Z7jIOYN9cx0rNs
3P7foCPykycxitMF7EsPyS9PboCW7ffw5w+VESk2oHZtBWHtlfbvX3CQDk2+QPae
92Q5Px9vJRlI7nXKK0gOKJDUj90jbUMkCw2/NcevExGR3NOROFgR80x3YrA/kyzc
o/rcKLpzv5O9ujdzOCyEo6fQ+qvUYsPmCUzvShb+1lzx8DvO5qQV60/Vg+I9Sfr9
5MCx897dxedpnVocxWvFxXiVPHdrnOc4KEGc3dcolMOxpBNbU5GB7ggv+U3Naq1o
+kA20sO+Tg8slxwwqUHASGVphoXbgVaTHT903hXXokEuZpZKk3Zrffh19WtgPk4H
sVwwk14P/ZyUqXC6zBVzRRz/VmEXvTlDLhB8MAysyqE85Z9C6PxUhvfkitj2BIU3
OZtQwuvs3xPdI3QZpkobnW2kqb9ZcluGJnfnoYbiicZwNPDzFvv30vGeehnxutoQ
4hYCN9QdgI96SO7JQe8VLVjP/OnM2Wqp8Fn60r8BwJmHdzyx6e2/dI1YZPdwkKGv
9wm9aDA64jy6XpC+NodigiHJDCcPU/gDgLHTJpcLlVaiWdU5jz+pbNbeG5aNSWLo
ziSPZEPskynxwlOIilotqoYjzMc8zx/7aCJuIh6cyr6ik6sR/rxsS+QI+q061nnp
nwmmzeh/YAi27q/2KVEtz6YEh8s0O+2XcSAvq+7S1BBOBEY1W53SpDN64S208zjn
3YCOvO5C/elpuJCLKyeW7drZ9rjBrppvUiuJu/On27XjJmzssQMV8k0GTAhryztD
sLrJjbMtb5/TxKqQKgCbW3bDBUhH6SeqtqAHEAseJGYnjyBTPYrG2tfmDPmd4nwg
mSUFC0NpCRPVTWHTfd/zenRqBnBO2VcDhpSv3cj8Ut085Jhk3QkSzSZ9THW/QjsB
/PkiRdAt0lII+GoI91suYw==
`protect END_PROTECTED
