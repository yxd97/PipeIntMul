`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+daIIqHJfL2BM+XVbCkTqbEDJiDOAv9YyvjrSJKRR/ztpzFGx8zZzkhEIx+a7/X
QAbUjj5PJuc9OvrFx372dT2cGKtCMqiNvoveROLa77JRbmWqX+yINJC/st9Wj2QZ
M3ThfjRop0q7sdZrNoSj/4hYifVwqIx3LVRnqf7FxMqIoN0cRDLUNwMsCgGPcep3
2XF+EaBKzyD8/m0Ov9VpSFB05cXw/kagCRDS7detv8WrytW6LpzToQ2sGdiRxaNd
r+0PaJxfJ7bHSOv57ZTorZUnImlwkFxvoCWc1WrtdfPVtaz8GEIm2KyZwQBBGYRo
Xu5wm6KuQN9nc3iYCmoasg==
`protect END_PROTECTED
