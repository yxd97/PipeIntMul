`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
54T/x3JiXmOyxcElCJdKEV+k7NljecCAtawVLKgn3iVLTFmJIQ3tuZWOplIG+sMP
LZKZrRdFjuydt/Je3J4uJduCCYArW+l5KSwur2kjEUBL6DpjdAJVmK172+8lqv4b
SYGqh0mA9z4W2gGK0uMWkXRXGGfPJriaGogqfAxGvnRoC4KX4SVBDBt+5sAWMOOq
oZAgUr/wGAlbOA0Fk9Dh0ioP59ksr/BUa0TlwGFaNzHlKhNawtey+lyCvOZyV5BS
Or8pe8li1j7F9NZeQGzT5E9TLyQMM80PYfPzNuIDo/grUoHbIaFCdMFJc3Zx74QH
GniZ6HldyY5nZKqMQAYGnhPy4gyFcTg8A99EVqQj4ZQG3pd9HOj+8imfLvnFLDgi
Itr/dGEjloo6IF15QUlMpNbk3lKDvw7H20RIaNBZUIpIVzDd8AsrRYO07iz6BX/j
vrYcganDY/1BcsXkl4Voq8D7Fp2bKsNzBznxx4op2k6bcu8E+eQD6J4pPiYf7t35
g8LAfBcFl6In8ra998EJ4UYDbtCqAvKID1UTI9V2W73IAiq9LaLwxGXnXLRw6uUh
ysg75IHyhIQTvbNZ8zgCtDkGXLwT5us4Cz6mnWNLxu2fPKLQi0mB8LckhZvcUbSQ
`protect END_PROTECTED
