`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WpbTDvd191nxcQWnyv9KQKDuD/hIKE9XsBkoupeNINjKkyJcCHCfsnwO7waCuxlI
3pUVFPlcL+g3cyDv4acxVdQY/EHOfNqdzrqt1taf0LWic4lHeyZz/6wfqm76LgNq
8HpguE+0DE4pkEIwoAMkFk4oS/2aG9g35p08fwscayRuAwACpEoZtOX7HVmvyIXj
kg7MFXoJC2t6aS0GgxFuCqcGrOLS8riN4zJtEC2FrvbunOZUza4TmtoZwXM0IYDo
PR+G6yMX8dTUWZclTsffF9eV0qkbTTyH+H6cdki89uKn7HeNE2f1Vxc9cirbnhcu
11i0Pg9P/e+LTwMe+VA6x+uESHYCNLn/z4fzTjpw4yMWBVNA9u9KmbCE32ER0Rox
p5881Gp77by5+uHYIl+RpdyI4InOt0MUyhp22YGqTSlUG/w+FaIOFU7uepnyMhV3
C0Ko3TvvDZ6U2IWk3+53FWqkDac+0A41oXjDnCfgU67A+sfiyz8R1pLZ7xnm4EXK
Hf0MusTxF/E56FTMYzTT1gloVnjO0KgI10P0b+vY76BhXuYxRMSLQJK19KvMd6Cw
Rvsckdev8OezpVm4SNM/Iw==
`protect END_PROTECTED
