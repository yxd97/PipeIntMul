`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gT2Jb7MmeTKYzMH+op1ba57gM6zquXOWPjc8cWtQMNkT0tmELRYwj0yHxCjG3hp
S8Z07jt10nsvSFt/dbmGiMAbIr7Qx4YS9OhWFe7f4nY3HBYD5FmztVok18ylmKpq
vE/GJZW/Dgl+czqwWdAgtQ8kXO8thgBzQL4fTmkOKYWTj/r6XfQySDInhTwKqxZG
+isAlDcta6m612aQXwC90J4CCtpo+RVwQxy8brkxfU2iUJPLounGX+HufyR30Yd2
xHbEgRTsH24NF2kmzJji+APe9XeQ+RLlG9G/Aa4qwE6Tfz5EzSJS3pmXPOkzrnHy
+Bo12GrcIp9YnzRl54tx6ZH9U48ud+Ket3IEvg8xtkLGbz5VvlZytgryYZVUpu0g
UpHWk2ZlW2rvkR5xrb8UTFpH3e+OxafWtYhIrpyFEwFtey8ADzw5Tme2BfDbHHEr
blSM/rVYzE0hCKKa6GgLLVe5dfOaDA/SLe6jNC/wPrc2dvR3w7yfe/G7HNcN6Vr9
fv/fv0yL9e3rFRFPSQ4B2M1gsaTcMi6fLCbXaLhSGQQkqbpZOtp0k48XfNus3o+c
wGgRr9ItHoUnpd2/6vXAgZclmFrwuB4F/qk1FDMJdhQ=
`protect END_PROTECTED
