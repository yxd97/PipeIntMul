`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6bqNebRJTuR1TXwXaRiuSor9Gm++5Xqg5EJMMn2pQByiCZ2YmKE9vnZhGGwbzx3D
RvJrYUeclAuGh2EGM9k4BUg0Zd7DvU/gWugUZQLIdQFZvXEwHPyoDnoIJ7qVO9Gq
7PdgPXXCNd7z8rzvJy7otkOmMMq22XiJ+wchiK+/EaneP6WtRnsErMlBN5NObkLe
LUJefDGtlYr9GuS6fW20yXbLI8DDvSumXvaDG51i89civUJKmHpegFwlfqINMoRU
vZ2wxqVGO0E9rdFBXg6VhCHhbRYEWHrP7hku/1lFhpceH9//GUKwWYlrAZl7XxYf
0Vpcf+cT88Mod2nB/Y+ArF6F16H2MaS8iBhr8xGtRrxEvOldNDVCJ3GCcW8WxSC2
SdIURXQVZDQETTkYpjAVImetY/XSFmWBPr9SktrbJpLh0q8cZEkMxYhWi349yAkz
PFsvdfi7y/PwBwMoObl/QBjwJHFSCXXk41+4era8zp+VHMU5+FAIvrbs6UOcVT4x
w9wfAMtPD0Ndp4aL2XJirMa6J6BgseqoPFm81iF79tPyr3ESiV2IgcBoDnEFKcf4
TUZYS3Ye1BiAjT/PByHqyJRzC9TQcpkff4MneBXRJTFKN1cE7dGiDiMsmR6qNuvl
p4R+URmHDgOp91vv0eDnT3W4EInglz2uVupGFl24DQ873Np1eysZgiQAnP5WOfLY
gMQkzBqELVwzxOchhqOKg1sdvF+cgpt6AXEUHxjqIEVwuaXtB/0KWVF5Wouej7T9
Yhp5r436tFizSLocGe8eDPfExlzxDFTugQP9c/wvgKbTGePXtAInFTLDvdwy/EcQ
hTJO+ifpVbP25w81ousMTg==
`protect END_PROTECTED
