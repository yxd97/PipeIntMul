library verilog;
use verilog.vl_types.all;
entity IBUF_AGP is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUF_AGP;
