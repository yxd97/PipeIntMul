`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zHiExg1QTmhI/yTOPNDz3RZQ3BBaSKJnBuBAfPzXHEgnMCxHfGJqRfL6Y0AzWmG
tlOIL0UxUFlMiAchDgizRux+uLDyq+J9Kmn7HAQw6ZFCvD3UvJNegCKw3rZ25P3I
cKb6jzHPr54hImj1u9MQLyBlwWUlF6KIPylWs5chx3ekEd3VY0SH+n3Lgkpeqb1l
Ge7Uq93xy88hKKtszlAwxy28x6fqBv8MBacLL/vxv4xkQx3oJwAzvmgDv0Hs3PXX
kWPhfEmM0ffYmjSblU0r+OvXVJXJaMNA/4rACzQ5Fn1EYPaQ8dJCKmCWcZEjRfrD
AdcXjGnRXGwH6aLNYBKrgHnIiTAofFZcdzEZ1dRG6GqviKOR1oYjJMWq0C3VyXZw
YZ2p+ZbiuW8whyKr/4BhT2nF9blYEtljMwaLX8MU/7HxtktO313P2EN4gexMnFXh
oiqGrDdDaZYhO4n0Y/d0FwDuKBrG/95h8Imp23qeP1hOn5GnzmlYQ2v7vxQ/rV0Q
LvjayoZiYAqeWmvZ0PdxssxeSRHbu4E7AdK+2hyq8RpYdOaH83bRys3/qYRhRJM8
3EolLEDKQLMDRTZigFwAs28XXC/45+N+/nKe3YIBaRLrkp2selHWD503URm2SsbT
ROBPcDP7gJhf37YiPlg4tv0z5QdfE8Red3mUATT/7wew2KjzaQyvtOuszT+Dn6Zk
PnDqUSElCtW3O3dnRRJexR/3SuFPXMB16VoORDlYXdbh5Fum+QlvFnNhIbFqXxEf
IAgJ2xK2wWMctYLVIfBOkTdf4SwDur53N6jgSmbVjDeCLRpD3i/UTYliJOZc6mD6
YhTGtJ3Jb22PCWJ3vXs+ZlxuNgOC9078g0c6swAyqRcSIFnycbhE3WMjIzycOKqT
5WknbfG36OzjHSqQtnSkUJApo4W6ue64Mj5MsM0f6XRvyqbb3RBVqX5CiLxVV2Jt
u5OA6qIl/p09QWJHcmG5KZNOMQ9nta1eGlGvDfz7R9Na3gPjXU7tZfB+Zr91PROo
P3A9d0ENaFU87COHxRXCR6kvV/7ftiMmAd9jb1x9bRq6Q7kf3vTIVfVHu6+kJin6
mZyL2SUFIC4sZ3Er9QgKO7oOmWJaI6dr5sTbuv/YOq1r7TwBdYeZtu3HxYY3qCzW
N7lt67D/T8L7JAfkxkbHbqImec07JpoxNLqbGVB7b50WHKnqyHCXRW/XBvVTaPFS
kVmqCmFOmA/z+hPPJHxo9ouLdJOxmkEb8HCkvRjL1yxyqz7IXE0CnCh9BuhxhzY+
aDv2BYMoMh1ThmRvBt8YKn7Q5KF4FPrOx1BkVI0U453P2uGHhu4nUr7ZazoykhfQ
RHWcAr2evCh05L+r6sJq9MI6x+CrzSrkG0ya2/CZWX1zaUg7Rec/mo5MEup8yWAs
E0FRq7LNO8V5jbmGEP+EP4TCRO5be3DGy/VixoAJQ/qMQUZwUdB4jWqo7erT3nPU
Hbg5TUhCQ8xfTqJnJDilY9xXq5FUjCTsg/QPW1+N5BZUZprBHuQpKS743qSwC0oE
9u5ehtZzD6jBqh1w63C1vvyo4BtjYPhOMJ5hol2j+/2Th3E6FEndCcYcPi0rTboo
+d/Evouqcx3pJ4uAYDaFEJjRFpyN655252CboR+uqD8ChdpkH+WBWXEsWsqwBXFh
u1LQikhZhoYRPWrZHZAj4yLgkQ7HtT3+vnnj4iv+uXEu0FSHO5U1Mr8NNm9C5M6s
8HuULmEt+UxwIpYMWh1jAz6e8UcKomOUOIskJCb2Vhonx+Iue5v3AOR7B+AO6RxN
YcaRSaXlB3FqIPcry1d0H0JnDIw/pKpsuPA9k2Zmq+B6Z3Mac8dSY/NsJAKZMC69
jAfD8TuZX2EyS0r+LCUyvx/zRfs9iarn235zfHv+dSxq0NcBOlj7TBLbZUuJmNPh
AatPOvAkLKXwnIA20W1uP97oQRtMfjAknMvYtfSmnKuNFGZXCpnJNM5BoQhNk0Ru
hlw7rkgmcnNpRjyWDxLpkzu4oZP49KrkW3R14iQ17uBNNDRPRIEcYG6NJN7PzHZK
mRfOSRtgSbZq8sZgRKLJtVx5z5W16U5QONCKsD5jX8WtyroUPsDWGXzzh2SUEJg4
r15Wzrxb7t9b+Dp3aAAvJA==
`protect END_PROTECTED
