`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I4gqTZGOimUr9SWkjw3yCPK8wmJjLCd6T1iR7LJCUxdGCPHVP8sLSjfuenqseIXg
B2eAeK28dTSCtPngGsTEs2pHNNYDUY+QTtvQcm0XYXp9feZZOfysUwPMVZB00o0H
k6xSXqzXRbco57UMPeLyW9GVpXmvreZCyEFO4OelgySOyB8Yy4U2pPkgcSJNorNw
XTCO69mHlAiabDRozrk792eYJswsG2LRrJGxnLCtDfGs+1ywHZHP1y5/r87/gxel
c8CpNw6MvEDw+xNmQsqCnVDvNd1pdUaBgBGE3N5HO4WzYKLym/RvoCY/V/Z/KITj
STz3oJq5uZ6ZbijpyRIcS/qLltlYr8qxVWaL2c/IvG/5JXUkijY0hTQlAnZJJAmg
srtDelYXXSgbpiatJkvHkiHJIIoHzw76D/eR+H3/8EWqKnEHb+h6fDQDv/ZEm87Y
Sodh+poLizdA86KBCGwGcCvmSVnzQIsSq7V8Y1g4IsxVpAC77xtO/3LFQP8JtseE
xCW3jXTm/FmaA86rFLsL5oXk2l1VVPr/5OcPiRT8yiIit5khkx5bg6bF3Fy+EFjD
ATo/SqcihZwX9EIx8xBXyz3SiNMsGE/WkjISgvBkYN2nz3xsFlYe+OTWLnUbCbZi
ccMvXX17tsqZT7TQNxz02g==
`protect END_PROTECTED
