`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iIujzzF9agcBYcANjTdzGJHIao/gDgVb3g0f3IwOGvcXqlNyMTgWv+1C4frLF6Jg
hAtmrg0STi6ksICjXfj9eWiXN/uV3ioECtZvgmwjs35qIfIMzMD8mNc7mjOadqaC
rAgil4s5qMSbizj+qOzDJvVaziqwUZyBBnRlVuNnOAgOMStgLqgEoDOwMu7vzk+8
bvcJb8EvBxwy+mSmyiIQR/rWt7JyEgfXkr6uUY5ec/wcbOWN7HEAlKZ5ow/q7Kt5
kB1dwDBlf59IF5m+L6fLeND3tmge05SjHdOS/T7s5Br9tKo/qsHPCqIYSQzrTMXu
vNu8IBGHjtyBvTRLbq8Bd37+SFFO0a/szIi4JtqhT/fRGG2rd2Z/L5ddY3tTp9Zc
8S5yxINUReU3rM6jk1H+iXsbEc66J8VdO0pnxYdYsXlMwKFKAzdeFyqBeUyObVK9
FKmfWeWNmwYpDTj5UqlIk/TXVhi2gYR4098MU/UX5WLjRvR0o1H4BVqh5bTwb0NU
TgHJEBoTKFuywAGwlThEHrMsv66xKN2MbnansFjuBCVIQlMYjFRmtjyCbolN1m4o
mwrlQuy+HWyZlxCdRzralODqPRH9lfFM20E6MYK2TwY/9MehK9EmZz/rHZJF55BU
ZyD2EjLmcxGmVLadb4tEEwRp8sY5mSkmJPFrDf5um/SS5hdrTlbOSXuLAU3whoyr
9MGB83p2U3qNgkV4BKngS+1NDpm1lK9RPqU1/BV4XTbJBNDlvyEmLVw/UXESOLWb
QEYqq9NKrzDbwWOWzuUh4SrjRCJmF4DwA5pLmfpwimI=
`protect END_PROTECTED
