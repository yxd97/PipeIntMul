`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jn1CQUhNFiqyT7te8wOkes24NhapJOaOqLimpTavGqgAATKncAGFKXx+r0AhlqkS
ifWczVzcDEHunn8dzSfggNszjZGIfekOYSuLRdNdGFAI5iVTTZWzW7UtXdyvQgge
2OJMkaPbY57LdVUiKAIea3DTHbjW2Pjx5Ja9QcIYNygdD+Y/zXvnjlgB/UjJBEne
GTvzaF+bU4rhnEOOdw0lSX0aCkQxrTEDn1amR8Ac1m1bFZgwraTxxFJQEUUxDgu5
7DSgzrKvufKN/iU3MhdvbpgUf2cljrJnERkoKR+JXrWrPPaABj1jbVVUyzeTzcS5
54NG8oLm0XQNKz9QZF7OROmqHThESm1LKPN0aza/mPtx41xkoXxE3O4eII2H9vb7
WYk6fVyO+LiUUHi1XxfkFW5qyf8xNetXVvfzKqrIIqZfVSn7S3M5H920sbSE50mp
YwS/JyycsjV3HWLWj18V5f4Ea6FPYNtJaPsPyDgh6XriIzyPQ79ff+5x9ZLUDTsb
BzA0kovHuns9rZFVwHcXtZpFPiOxERVTgpA1Fntp1zKuurlxolgY2biYipiI8f1f
I6CJSKhRWW4fPa40EEfKbDwi5ltRtA1/i6Bxu2jA0ZAxDQFDi2mys/7blRk5kYcz
qSffz6l3Fk9DYtLhMkOQKPIqBa7YWrKmj8WC9+lb00aSDrpn5vlWkTz0uctNRqgB
Dmh41Tlcs02oe00NZo9EEEV2hyo6JodcjBQ8bg+Un3TAOsKOLI4KIxvpmO1luFRx
SITjixurAM5v9YOWLCdXJPK2gf+3WRK89EGGCb29wKSRb8DG42mC0EAA0m7mHb+j
Y2ZRnITPeAgL8cjg6ZChl7hbobfExYgH79rL6ZKLR2NYCULfWYVxXZauSlII3cOb
vurehsVKcBVHu6pH1z/YEX1yV2dA94ELNpJUTyjRcHh7rDs0uvI3oXNBloM3qYpR
CaX24oxS545kkJ7D/WlRkCEM2wDVO7EbqZDJUQo77XOvL/4aJVB5V832E3Crkw+y
v8eO0ajIM5ExfYC7oxjcfXSBbvEL9j4PqHiimu/n0OO7RCcbPrGyqAs+y1PdlwQ6
7K56j5FkinDSldsY69oT1xQTIeN7ET8GxfdSUc/8Rd6fumtwD9FOVcnnS9UNMycR
5UkXulkU4lexlZkL8G7HHorkgFogHvahP9JXG56s0VciL2N9BZjVS85lHbVVElBS
dQyvEkyl1Dx7arYA9IOQBS3aPF3HNcOLNpbtadkaaqDHHQ39q+FsN5V/4stUrWGW
5uau/6pOGUvUsiflIfAqkYtlp5C3j6Uoihw7tv+awI7+OsbuGGLVb3i+mNnCXoBe
r4IxBn903rBQpBYdH6BKrKj0FrsI7PEt9veDAQHUs+0D4rvSAXDBj+mnQk5LxNQk
quzxyHmlnwQWQskfFyZDlvuAFv6acoBo/u5QAP2B56+JJWG1XRhA1lft6UXsqZe1
oW8VImX1zdEgdB8E4/5OcpzJpbS04aP4n7dDyuL3vgWq46J2f5ogHJlT8+pbVAtC
X2navsM49j/LFE+SLgl7XPBmtGnKGLJqDQCM7AAuXGryAbz1UivnSEd/thhnSTSN
66VCDrtmyWTlaPJn6uJ6j3yca7QV17L+PaJd47AYbeI1qXs4ZHhXi40uVrKFNMYa
8VnxBg8fiV8CSCwhv4x4vqaBKHSG96+oJGGBmnuUFS22ltIWcEqCZFfJPhi+pi+n
kc+nNANxQI+1N4XBJWYM34y7QzAHKoDEsLTsU8/LLLmo1WCotl4hJyZgKYkdLetI
sG7MGAxHz5QWeJsMtTIQQXQ3ckYV+yEhQulqMuOJ+SjKJdRuj9woZ9s3CfnPKdPZ
ltA5LRww26Oj+plADlTipU4tTi4T/Xp1nSwOnyGnz+awwHXKCVfitnBJi/i0WGcu
SBNZbZax5Zq1zjkiA7MmCvRaRdMtHysBWuvM3plKGNbhpqSwSGEOdFx5mDDhrzkw
x+mibsDeZqjd9x2ziGOiBmCiBMbNhg4sfRckFXNTYzvyhZO6IK5KhY866bJ2SQKm
K1o/C9wPem4NXz6cjLNcCdDsuYgdbkUFq1Nt8l21dVLNER9eVCx6ILb3vTltSn5g
V9tkLSdwvNORa8+9O3Gstz9lwi1xuETiz8M6rZXtCP4YTZAXsLi4p4IdSCr+I7GP
WuCd2V7YalSKPVfjaAnrugmdWt2nQw4wrKXIpsa5pbnfg7ngu9M/86nDDCReD3sw
nl/l9lS2moJlw9bNc7tGFaX8PX396WvxmdfhB8hOgyD6k3iajGgMB3UFD5qih6VB
/Z1s2DmZb+YAE0i2BsT39oBAtUiFo3OGgw+OkSgLtCq1TwChvn9uTch4j+8t8YWY
WJzz7x4kK+9Z3fEhA4nxJcqpNgZfvP2YYPXm0jjVrSzWmbA5uvJGSoH2pjvmrzFR
QyAVjdk203fUaEJp0y7LB2LqT2ZeZQl2e2K9hHGf7SrcOUzZJ8pQ6CIeKL/pz1Dn
In6YuF1B+Ba/SgDiqAXc2D4lyJZK10oXEKiNfsUJub6Xemy0kmR/8W3XH7FC6vB3
7bUh8dDsIXzI1MRS7AS1DIV7kT3/SRFDsxo7YbCpjBeB4ST5JFMAnCIZmlGnUsVS
z9fkqyEW3l9C4YD48mJRcAuUcaDqWlk5QxqSS0PSI9WwebdZO8+KVAaTCi61H5sP
pjkT1RQusBgONNy5MK+PvIhfJDd3xQxuym/qHRf5lwGIdtBtxQGdiukg/T7XFzIS
T8qbRW9itQ49vL5EYpFvPlr0wM4Qfk7RTOauEshStGQO7QiRrGxHlUGdntLo6GJ5
Aq4xwWxjmGipY4pLOfUvRjretM7yiHLJL1QPImfmCt2jnHxrLbDtcq5UNjQOZA7U
+CsmH4Vpf4KkF/PlWsgx9O2XJjMfO7bxWdkBkInbMTIZzBtcUurEgc0wQP447mDo
d1IBilMkBkyHzDvQ1LStdx3NVztSQ7uWWW/+JrRcSsX1OOnuvomYKK6JX0mfnpoE
EtNEjWe6nnVpqho1iQ+ettgrFJl7pc80QscW3kuX13FjwZ9ddKy1cDVpVWOWPa7c
gWQcjzF9RgkW9+K8an8fFnuBM78QnxOPTbVetB9FzCsPuAA5DBCink2euYWOKNSb
X7nDm6BBXUIqKguVRFxsvAN5MMpytQnR14pn3+2Dm9CdlAx5GXUJD+UxwUOVyjRT
RHlCoxBtBwHLks0yu/4QEHsefgOshN28quPuUCFlFx60ODhl/7wuUTa79S7GW7Lx
LQajiqiq0Fr1s2b/r5hov3AWjiBwoTO3zdV+ub9W+/l0o3N42qoXJ6M0q3IJC/ax
FMv6wKt+yCJUUkAwqpJkOcag3gL/24xuk2JYcVElK6VZAVE9obnJbtnVBPtcTLSw
PxzJEsA/u8QeDpSHpjkHW27pplvfIiOKTSLwYKfnc67XimKlC+gqYlBkhdt0Vk83
Rvnl4JkDJYdH60pwXuBDU/kR5/Z/FCil5uo0HQJWkUn1RnnYHgPBRVi+ypUkby1a
P24cqsPmRcv9hEk5hdTKssJ97E2c8dkVoK0iaI4m9EA2pRYoh86etqaBsDKr3nSS
ofGCwyEDkmKpr91FToRSmX26Z3KrJ3DBBVCGnxTdSrljwmL34cVY3/yQqLouv1GH
Y5y/XnX/WKb1fdlVz2+hW8n/04tlyRzgA93o5uA6BLo=
`protect END_PROTECTED
