`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gL9YWC8N9l0clS/xspPhnR6KBB1Yf8mCqvycNDw33rEPCryFx737R+ErgeZB+4Yk
+uofKgL6K5Aa4OwZXPHPdSaqNCLG1hM7LfbHi0t+GZFC0grxlkX2aupJukmjSTxP
WrBWk6C7fsxuzXxn6JOntNNF+gt3eNlxtDfBmoSEkjZ3mXrmEuJCEgE2PGy0JZzz
ONjb3+RXM33WNULRwm8Y4JjRVOj5Zhmc3h+Ua67yQqZtPIAlW69xTdW1GvFHCfAQ
t1zylElXvDzg7rJVbMMeIptQKptqdHDN5Y25PpNSnwERXjcTjrmX5PPmHGI3ckug
ZzR1S83NzAdiY9z77Qb+yQ==
`protect END_PROTECTED
