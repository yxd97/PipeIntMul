`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eqXak5wmXN4SeJwPMDi3SBetEaF+yrkj/iFy2r/nKUKIjVGlOxUzBX8TPDXDXKX5
bwXcMV3XVB5UD9MmPQYtOlxETFIVUMK4Qj79OdSt2MyJJeP+V6A2mxUbl6rEybIH
eEoIopGyMq7a3Xa9v4c0hDjs9HdivSTcKIsf9S4z0BHse5/FdRfMNxSfRy9beLaV
Wj7o62Lu/pfarHCGJ/G+dO+7HqYV5HqZRyfAqvtIIsGayKN0ToJhe/Sk88ik6KYv
Ytm1M6RyDbKVtcnaKnJ4PJEBI4KNhCPRLq+fsTEAX3DKxKCSYYLoUn2dORIesVyv
SouK4aaW1r04E65Ev+c6W5fnbbBG1zI7NuCIGMLnzsUMYkC9i4faDYVvZpxbABuH
iO7j2SplriLFMhEJrhudmwGcWNw+wdnlvQQV4zYDRd90CSz9waHJF1kMz/+SEHzW
lEFdEtwaoKuxD3p6Xi7qAssC4J2GdL51GNBaYnFzrLRWqxcVVrVN7MmoQarT3IO9
Qh954eS1y1NQU0KlYeHvUhic+DkBpL+mUQC5MYw70/HDhy8RAxJt4y3jCuFKP2ms
py7h/NnlgL50bEyPQ+j6Uje1y/KYSoYAmuYqhOGGWR4fIV8VmxZKRb41lcjZTRi0
DYAfB1ROMYfZdZ77rnkIpMG0UgAXY5UJ6avTrnnWsoMpa9jhWjIWmX1mPxJDGsT1
S/Cke4Y6wEUurmcK3VWUD1xwYfD8Wu8/wViupphcyXRe7Yte6mSPQ5hdB93peoP2
4PxBnKqq58iXnEvSdCUGqJKyxVwpvLQw5ZRUYAPdBvxcSRXac3VCbj8132+zTH/Y
TUhPntUbZyTklYvouBQOgKyjOu8724tPYbUlNYJNVHtIcp5oB6FPA7/QcDkMxtq4
UnUQGDJpEo1Yn4xmYegCWXo3ZetEny3lK7BDl2z3GphQBpwUmdN9/uW4d6N5puHr
gQeAopSYN53HWYU9toZnGqtv++BBr2CF/wmFdPcmxlXY97vgVI0nJiIjIscT4Oxx
H1zrYq/Sap0hKSNz29yDDi+BPruICJC5cY7Kz0ts+0eRCtMIMXZnH6ykHOaqtvw6
ZRe1Sv2m1/LfNxTwbdReTMlYMRfQRJRdqQkrF3c5BinZFwiQIOlmZyqoaoMecnpa
BlIAdCotLPHFjc7uDvBzwABFo8FzWecYPzkthPLQ/hQgzyaPgS5rkwrnHrXv2ix+
4QmWAY+L80Q97n2n7Y0WCTSR9/yCwgQZ4NjED9Uvt/5cWQc9uS8xB1Mvk7SWLJQT
iA6+59jWmijMRttfOfiAeufeHpr05jYSNMviW9JKUENlrAF7Qa3Xccfk0t7YvO/J
z6JWvQ3hJo8G8ot4aQQdrIiCcbvuK/I+8zkPySAr6Xa4N/W3AfmLTRNK4s8yAfOn
zTMz2xoN4fS+EcmtNJF/cjLUwOMIwDLcMo0anBkFEiH6GRFs/Vwb2FPbL86jznNT
HOkrM6ZhaRzDAiWiwezTxQGIuCAxB4vzEI1U+s6sJGn/F+cSPBWtI78RmuUpE72f
yvwL33lcA+4cAr2DcoEE6jf/0TIM/Txbp1sGhgNXui+bJ9bHEpEXgZprx255tT2r
N7jYomr3SyvBOsJLKPpDLI7z1rHDn6t6YFyymMVZ6dKzdqWjJwEk5K8g8UmePuSa
wDYWH7vu9XdmKVFvET6prE1bfTjYRxXotX5aiL1mrsc=
`protect END_PROTECTED
