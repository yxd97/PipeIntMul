`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7HczHaTXDQ3GJs1CrKA0dGUSEpi6KUj/Ves/kVuFoiSxRZz4PzjQ+SkOlOW6WvBH
UhBUW5t54jCJVXyvxMniciQLo8lqrL6I8rnMZZLHnely/eMA9aa5hlhxs9U0kEjA
GbnVpOzz/yGNZ9KA19LMB7hQ8ZykWPl6WcxsLzVp/b9AWxVi5GO3vdE0QlJDnjnG
TfynVUGl0DXwOncbnsH5cVTQh/23+xeIRkkhFLNixb2And+DIYVxhDPsqIF8Y68x
olF8y2LSfCkzvZReZUdV74GwOHlULBB1nkMwqBZh14LM1AHQlcHr8FOVCSHhix2D
FjGF+SkBZC7kZcMJiVpxq1j9qM/oxrxFV0aVXKT9c09bpl87t/jtBgZQiWA4TAvw
IqWNASJfPZGMiIX+FOas0/1jfwI86z2R9m3LPt/IoaLvU6W/QHo7FL5RzmjHXih8
Ea4iPVd6mizdQr74P9IahqsJ33pUmXpooOPYxesQMXn4dQLBZACKRcXkCeqJ1PIr
NwSz+VRZscUR6xiy+P5Ech0XDgOc4QMcRmPi4zhEjZb8YWx5XL9Fx/QTKDtnpUDp
kRceKjwjqH9a6kK76HzURQ==
`protect END_PROTECTED
