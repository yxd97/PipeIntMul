`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdVcUPLZ0GP3cCT1a14tzvcrF9UPXr0q7ynyX1S/PCgSu0l0OX4huRoVuCsrwhse
QlH+Kf5BPGSPzF/8yn8WQ+B19arSaZtQjlyVb1n/rdm49hY1YmOscmRGpAt4IGaA
/75AaIZzzkCKo/t6uql/MsFrdpw+BKe8ddQM7H6Z2kWlznWL2a2sic+nsOB8YPF8
gTswrhwnelurBHxE+F4q1Begp8r0UYR6KyrHXv+TaWT4B2CsWqDbXrBgy/dzbndl
E7dAgewzVTQW7WGTJ70ZFmThma4JVG6KawZc4lvoz/SSaoZQSsBqduXgWrNMd2rx
U256fonGsaI42RrhJU5nKjnGv8GzRn/It4ESNMJRDepFs0cIL0WPedUzFf7d2hMB
kINUFK5cE8+RAZ4e1uVsp/UTKqhD/ugtZTbvaYoDeH/ysG3cnBZ+o5/VeyStrrYK
KIS2UHWnMEO1uu6rejBXtwE6HRLH36kIjUNoRigmXnfR6Z5z5rOWybRp4/Z5kp9T
pHFphh1G/dv2LZFKgh3YKZQOZnpiJce6sYmq88GTo1UzsQOPm4DMQIl3yTZTidpG
iptFgjrbErrao2Xv7Se4q8baqtCygwLWtZ4fsgwUko6H7Ya7f8UjWEskLzSAAB5x
m25H1F6BDt2KRVoEoeNGTsRPP9rHL4llEVwWQZctDvedUe9FrjmOqMHaZTqWwG9z
9funqiigKbZ2yW4n+bUtjsoglxXEqSq9e4ffuH3ymp6jKyqEthRmOkwn1F2MofOo
CbOhvo35AmrTYDCW8TG6I2Hix7kmRptW75xWyVWzX6AeNggkTuFPFTur2CMrwjaS
tks5k+3l6CFWwTG+bjghcNsrYLIqhJyQ6Tua7fd1GOnYIaZJsxNJ5uhHLySOH5jF
wdpBP0x43xQy4WVDFYciQi30R0BPtXyEhlGuIcWD0GKTDAw29j+NR8wZN2kIUZEX
kjfEB32Jknp8CcrRlj8+jTVBgje9AllNf2O6cFoUrXoOw09DORFwY/V/tnvrwxe2
ZGl9cvfy0kMX/OzxanNBpkndigeFNvPeeBD4cc448wHxzGttzd2Wnrc+B9bOpHlo
Ush4odQ0LHp0wFOleuXtQlOHFy72X3P8mAp9j5Yuh+kFxjZPKVlY8viiC8mdwhA/
nUjFDo9Sp3dQvYns04PJgYrHp/cboeUEn3re/Q4uT9sBvZpCuuf9ATs8+Uvb1JlD
jNQpmh53Zg3TD2hIdxFRUDDZm8G8oovw9N1MyIArhz+5eFz21FSUKTJ9bSgPKcDJ
4jm9teM+hHTs30Y+YVaF7YSzEgrNI/5BY2f1p46COuFB6oKOPbioQM+SIRuGM1pQ
ADJXJEfBllClXgIpAgc8N3fjhwJ/u7MtMIuP0IuNSnPJZ5FvkWPva6h0paxpc73S
MDIhqPumAdmupJTxp+hZh5JYuChG0yncM9s8oz5gS5RIRL7ONCla/mWnvcamVm4n
V+p19+64XIo69sttOdtt5fUxclvpECb+0fw6cBHqRGZqcDKwWdJyyIbEsYwSG8BD
WY/7ej6EtIdgkYYJSuu0B1NxY1eKT8rqPNiusujYKnTFbScIWdiz+8ZKwXCYvnVQ
GAEmvnYIWlSgAhUgjiQVZBGwQpb/r+m4ZdYIP5XCY3zhUep4WFnyrAJnXi1AI7ZP
Qw4lrxGbWlYeaZD652YzJJPFgbESYfBIPW0dMBUEJighWxVN5E+A7DmFu6kbdR9K
gpH7ETuEQCQrNGc5a3o5Wj5EZ3+DfPGrL/Hdn0y/57g80cmQuFZp+Ful3zle8VHI
45/OTCV9f7Jur6sBL5IJonWU27kcJ4BcSh9fbSy4cY6mcsgh5rnpzF5aHzhvMBGn
UqFAH0FftxgY60NYlgKA0YvV7oCqPNAa6sfV8fRd1rFaCjA3MDCotToowuLB2xzC
1xaFtBYgsF4u9ZdIrDjeu2ZlJvKTZmS9ytKCGDXD+JsicHKJaOzDH8Ug+/QZ/KGV
D9DGTI5VUZzET3WHPOy4fPG/ja9SUwZQdekb0+JVKn5TQk7zDJscfOQu+jDkRepW
WUPhOmkESdrpeh9ENMLZ3glGQSQ00eHAytZ4JxRSkiDzw0ZIKVGyirim7ORPkRIM
RBF/rNNZK5ymVtbUj/iv4omi3YA/ZP+gZTVbqWjA1CwQ42orbSqsM+ZV3KYkpOP8
OeRrpY8HJgJ5c1lONpyz14aB+Ac6C1F04PbPd8SvT2wiA97OApcoj+RlkD/120Sj
pQMYpoXjMQWQ/+hiCzzhrUAhXTscu/OoLERg/W+w5qBEyMRWynTf1rjxg4D4sYiH
jUAIUcjV8uRL6yQ90K2aJL5VEICRv9z1UROEZ1TziKqG9GDwOgv/gEWeGlebBXnQ
40Y8LIBU+VILM0+PZLcxGkDzwX6wlalGpUJg9Vfxn+U=
`protect END_PROTECTED
