`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q4wHvUid6aGr7513XUGC397/O8zPBu0DM7e2IHprt1tjS1J2oC78XKJbqDXKTgu+
SXbz/6WnJMOYn53d65yMzPZHoQIzKr+kQb5fFBSSHicvoAa0KwnCMSbQaDjyb5n0
lwhlpNyHVQTLz2xp/F1s0cefRuaAJTtHeRFPjPL0FPoR+HlyV0X+bacfDPOyz9UO
OOicWzvertjMZuz/mRo/Hjy9uPnEDnTz52xmGMzzQC1ZBQFRvhjD17QFwKwJu8WT
8D14/CPOsg23GqQevwAp3XEVKI5XVNBMmTu7rDoiSjMiRocvP+7JE/360ek40+qF
uoudVSdBaSRa1fU5co7ckw==
`protect END_PROTECTED
