`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwHa/To+A/00GStZ8QZGDV318elaiYMeXS65GRUMWgfOzp0on1fSppNRoLkKVVcF
gH4X/ARRXsYzkj6KM3Oxr9N0+2kcZmK+maFdR6n0Tlsf03lMWK408oWmkDDDCwFI
EokrLgdf+XbJ5rGXN2tpGVatj0OQivDizL4yyDHkAu5sDoq6OfNTnYpV5JCoKDAU
MqCVebi0isxOL/Ee71rQew2ZFaEGaalkX25+N4I26MlyQwFYRbf7rG9esT6Gx8jc
MkvmsiMRPvBrCV0bIcvf7iGlXEDfQsZVyPy5DGXVnzfjxh6Le5GwrRjYGvuSTCli
NSJlUr4oVpR1kvl4e4E3kTNYoO6kDWMWwPfQ9nEAW35LcXYISRZlIjrYfVg8yncu
uj36K6h+ajFL/tZ38Pm7H8+Q5UcOd9nkpXCGWSEfS2zdM7Rv0kLnpH0dRgKNb8S4
nbmlnSXOn6t4+wE/OZMPomN69Td2LsVnKvOH5F6JkH2fI8Ah0obVK0s/quDxNby3
f/D5+SItOXZIfIjQqo9uuc2w9ssu2Iv7oJb3jW8YBfdpetBzMLcuUZH8dqWQ7lHV
P8kf/7NLoSyau5u/wVdYG7X5LBlU+44ltMgR1dtQXboT518KY/M4l/2eZ2TxxiQk
0fIxy0nT4/XNWCofPPJ/Z7IqVlo8NShAN8iNy8PcsLLbT8BHHxvyD6lcwhPHi/Qt
O0TuyZujG8jmu+HqhQKBYRshiHhnmhCOc5XUFoyLk2mug6GP5uwdmB0tuq/WR7wB
41wjxzmC9AjUpUzYW9TYoTWpYNC3CsPrQjVW+bC+4WJ3ovYYLUtjf/ykfYnF4yOP
KvWp0WZcEkG9nDbDq955Ek/+09LeDZkdWHZ1yO1aTElORuNE5Ncy1KhEiOx3Iq3w
rA5Rbxn3KUHIjVWAPVc+OVx3ieEQjX8jybYtCTraz6q6LMkLBdqrzjTsmEKbd/o4
VHjmEn4I5A6RPxHmf3xG1vwBNn4hDg0HLrDvvWivhBEgXMwDQdLf3ZHxsK7jvwpq
Lfau2ptdLCFX1D7ra+Yhuo5YuGahvDfYWPbTSF+y84UxjLxIS8QqbLvee6lEsXKR
pm7VISJgLbfMTe1RBOSpw0PjxutJJntjJdrUBo5rxY9mMHGx4ejNJhIfHHXAR81h
KRt+8oRL0wzpWRZLJ5VJbzPBkpmvhRS//RHMThZt+ISNL9PukMiVQyW352C1s148
sRS1wxqREim17jN7WrAZokMcvv4rDI9sy58UjVKo8OicUSTekNX84mQCOEqKgkbI
`protect END_PROTECTED
