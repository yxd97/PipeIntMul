`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/oHQPfQCTdXYrn8QGuAXTGhLM0HThZkXUzISIPUB9jFB2i2j28ImCqk0hYEw+4Me
UPoL44Lnc2us1EIFunRXFcWzHsrBqdFriTJf9F2Wm1fqc1HpEmqk4+GMcOfsUDV5
uH0xvTV0NiYXtXZL9Rztha7tu//MttxRwJooj9gfKa7eAYzaMUmEkX9eCa022Usj
cBbFPanwTtdrmAdkCNHWBtkWAhFf7ME187Y8ImAPpasZYE4EDK2WYZ8oNzqBjpfn
r+YzF/JlfZz0zQeGmYPGM3c9GCve1R6yOr1DzbYfCsdOzGiJHxSIb3VjOjUZ0HKs
1vL1h8N0mle1CfM+yIzqkdneoiGLuQo43TuFm1Zp05A+HsR2t0kjbe6z50vGzQaO
WvjyhmUdegVIR+4FF1ujV6qr+Lu/d3geidGy4cba53Kp0pUlJozRhZdVopYUF1/b
bSVjfX23IuolSGZD83yCJ+m/EMDR8U3c52xLvQhgqvY7MzczoH5pJ9UIrVGcrBTl
H8YXha9iL9/VfIHKoMs8dUREhQCdWuZOklZtLKxGp7sD3G0RkTo/s4qD9j815TmX
EbJoNTYoH/6jS26PfRPz/qnM06qbHEQOqicGD0Q2gUGZ8P6nxYq3gHlacio4Cc1C
HKlUzKN8OUlnOs06cwDk4S6/oa7Hk40VelQxRQSpKPDG4h6Zt+2popkuDzh/VgOw
FeoIYygZmjXlp2RP/Ajq0PmBLsywr4GZab3VnZhSGqs=
`protect END_PROTECTED
