`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJsG0miDFjcIHmYKojF9U9lOnTnzAGyLsJRAjA3/g9LJ8jzIpx+3oiOkC+EiN5GE
l5p6luru4uglhAQdBj9oScXLlxULAlAg1bE9xh+pdtrlIaLPwbT8nPprSJbzFocG
5+y6qPGX1o+hHJcCmTNsLn1tgHAZSqHYCYnHmMMo4m0qaxS2hzKVk2C4ymT2wv5c
8alGEFO30MX6aiRapW5qDAXjifavqk1EZCZFnIbMVCirLFihBj++BbsyIv8Q33wp
HrKsIwa0d5jHDL1oULaPwA==
`protect END_PROTECTED
