`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UhtEDfG3qo2SuF1feKOSOdfMSRIJJbuWdUJy1hMwdC7EbHpha96JAwKvE49b5I16
S0cIECO7fw6CpbRtFVIXHE96j22V0yAG7jvlHMkcL4HnmNM0hShNmp90JgcnUQDm
DD6r4TM1osE1EEiCDHtMHj2WPzaPHVVMEFukDslZ0WSrLz1jacMNZYI/J6L5cVXz
RIxoa8my0TK3Rc4vVdJMig4cn4R5jloKmKQAquSFMoa9ZkZb0WOAhtcaxUgudAJb
FmEoJUHFgiMMHPfIdbhfbUisqsJqZmRfx9s5P56pxn/h29/3B8lAf4V9ES1QXI8S
VpsCnJpGL/+1LYjssvZo6NAA8JIL0/McJ5sN67BwWt5IHl37xh8g7of0t+s8+tV7
+I0rRIF6iv5nhGpuqaoedDm+WY+sYaywquxYvjg+2QOw5DKT017ylmQfMW9n8L15
Bm48qB7ijU2gnuKnbA9ceiLJ5ARPzg1FRX93eiqLo4lvyD4c8t+FkPpSq/muHOW8
JbzM3V3pg07pn8mh9FtAabbKCluzMb2/qv67MmnKbFMCanQ9Mp8Y+CB1I3/Z4F2k
OdmQ48GAKpcOtvMLID7KnjGFL5/ETwj1o42/Ok5BbpGxQKDFrQQd1PsZJ0XAsDMk
m4slKw/XfpHuTrX3dVOzGg==
`protect END_PROTECTED
