`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gaJSQ91cnIlWbYKzMi29D0WmHJ2gHBSu1TRu4wGorcZMgktCkb6hShAzjqVCrnc
qlcE9DOkDIMYfYKVG8JXML4i/7hM3YcN5l+GoqNdxFpQinXcf7verFqFw5H3DyRU
zE5+dIdbNlKF0ufszMMCZsL/WAMfbpPtD8PE/2auRmiKXcD/k0xiJt9ZCtSq+SK+
WlyH5WrSWeVnQD5H3qPmDHilzeE/ktPx4jMP+NE5J15oMNtBaxnLANnJPHypmHzt
NHVcYb/KeTeDHq11waUTb4Jy+b7iEviC+aAj48HyjATZr4oXcnbA6q4CGFyo4gzO
XUkqL8XMFEcC9M4CtJIWooHb6O0NX8TzQ/XR+eumzApesCs4efoEQKlzD0ndNb5H
RtCKWMIVBDdNc7jT2DQG+60U4VKo0f7tgY+iKZtdrbk=
`protect END_PROTECTED
