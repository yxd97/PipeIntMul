`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z1aXio4yQMVvnaBL4DsEeFM7HeKIZjDeSyD6ixjiyfvSsTJUwqOKv7e05I7RatE9
Xpczh04hfTM9y68TkjjjQobGLnf2AWeDVHLFh3jpZpD/ZosBDSDV3O7Bqz2oHY90
gYw2z2/6XyDOd2jqIM9Y+BEE9y6TDUaYEhVfZom7bVy51llnrU7jlbfuPzV88FDU
YE3h1YxF1awclLyPKtHX3gHhrKa6nnb63JoisX8EvDsJp4a2Yn/dgQ/W48XL0a2L
+WhbSswku/I0nY0jRr/oAA==
`protect END_PROTECTED
