`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O4dhMGnUfXpn8Y/stKY6kdQxVqVz2dxHOSTHgiY25n7JBtUEbd0+nWBlGCJpD640
YO40UVdIGWCaMldzLX+eV0KdPEZxANn8OAC5R3u/bML+WCg0LjsPM9sfzesequMd
Dmi3KwJZ3n/fuNXxp8H7WafvDN4re/CdLdgn8lExEUJeMo3x7KKSPgBJXLE8t6pT
wPx4flNgG5PxDyKpmXCrE7dJ7X/zUeL2vxlUenVV20Wf7bPbdTHc9RvrK/VVa10+
Na9wken1zXx63Pa+udyA563tRNuRlKVcSfOgBShjRVQxJjmHRkjebPHe5dWY7A9m
q4lqSUiAHwiN91O6d75QGg2MqLwp90ktPa9EVzK2KWb19F9n9bX844gxuVm3rNFQ
ZQwyMgne2py/DxRFEcPCq6tlw7pfMRk5n/I/RpMDxVKc52ARbPoStkeTvA4XtABJ
NdX/OcNrFncmU0z8UslFqXB6QUqgby7857h2PX1hdT4IREy5o0lGrXjDjhEiug5y
Hlc1NTcjCxZL4AvkpVwmIihHdSqSKVBac+U45M4tPLi0SEAU7pt8eaDq45oz5M2t
ZdFzqBx9ee7Gc5xlX51PWM9KVECbqOCUf41cikrcRwh7sLaOLakUfp5ad41+J08K
y2sA9btSAF6+Oj7EeX3eECQYMyeqSjKPAUqmM+FhX5W24tadwD2BSfWKtl9IByCH
eBH6L/99Jij8IrcsqkzzHpLUrgco6GQf01yuhgqgAatIk7OpVb01Wky7Hadla5Rh
lfkz73RNmigEndRuI6gKLPYR3gt4EvvGZeFFKTEw011nX7cJLkC9BNRPxyPfFQcL
CNpsTGz4oFKdMalnBIVmuhtzUIuHe7aeEPTDPYhuENljyKONLqxoQ6M9/xG2vPdL
+Zlqh2+KV5pMuABquGTFio4UbWCOzNcLthG9of+QgVvrAvk1/q9vz8k1XzVwB7Qk
whWllrajWMg1mwHkCcCkuSZp1mo3mhyD8Tpt6yRpkhr1gAZOFvg+yKXKIUvSBR+J
jZxmLhUl1Mndg2YfREEq53jtOxxkl831sC7E2qzIIszAdwh2xRXUHNqOoPKnRP31
NV3dNl0sE5ca126iHnwSdvEHwC3F8R8Nqz4Daxi9j0lXuha3Y5Wwp+DaRz6YR7Ou
LvNKE12+ctwkN2/1Ox/6Dg==
`protect END_PROTECTED
