`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EBQEb3Nf7SSC6vZnEhyJKK5Faov16r6DPI1eM6aSVq32vhoHlhoQemkw3Y2EuCnh
Jx2i2dMCTTF+sBpEw85ZgiAEd2kfJ1s4cD7eFm5uRkcbUU5bEDNmmtHLE0l+sASU
RNWQjp4SJmjhPq+1bDAy8fV7rPeJQu1HM9bfIeTWhsSP225+Rcp58d9aRPshZMC0
thRCQ+iXGX1g6vJED0eg9qoEP2x1OA6FfjqObUFjFpI4fTV01yIlyzbYNQJUA4rC
ukA/w6OCXtEu+QJaHDisQNVXvRmxqveTf1GdFHp2+TP8eeLWHMGcEr8aA2bcErE8
4afJfPrvEVR3QQBmYWWex+PBWpRNuVxRQCxI86w4o60pOkmkgPJTTmD8ubh0Stzp
TzazhteDa67uqXzF6gkaqcccIVgBfl6fRT8iKpFvL2EmMsOzHub65Y8m7GX5T0pf
6HFsl8tUDHE8XtT00QJ6Z0uHT5HIyW4LQT9V72EZyBj5LEDzBYQ1P4XOzRvhY+Ch
gar6XwyI5lpwP/sG0ZU9lN+ZMs9OLWwPNkfRbrhQr/GlUDy+HoYQI2oDTfZcJqg5
b8NQg57sLF3Z7l5dz7nzpe4S9MS8LrjB+I/6P5rY1MtztytCvss9cwYoIzfZh2vB
3+1LipVZWTLdBgeeIlMzF5lg4wxH6og1s3te4D+AaqL+fjAaa/JdzbrSu2TW4eCL
bnQuZQlE6yH9iA2OwaBpfo1Gk9Q7I0yIvExVIOEIcMo=
`protect END_PROTECTED
