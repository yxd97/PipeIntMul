`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLiNGMzxCIWf3zPFjzjnUYFdghwM/MDC0NNhL4ow7XUdbZtHsO/gJQNA0HexFyxz
9kVWKv4KuNceTCktfhT4dwEsUoUxQ0dHQ+RdFVk8Y2Z5vo3+ek+gekuYNwbvf8RN
sv2AglJiO1vBSolXAlHcS5/gmlosISGcT8TldDG/OXkFP/BaWNgDnJg5FkfeZhgw
oZaPbTAV2fMW4Lfg/tLq8x+YjpSsNuEQTbMoTB87Iistu3fSNoK3qmWrPS3lE4mB
S0x/noM5KeAfhN3ZnvW+J7NV0KUgVJluCfYvFeF0U99ieLvXZnJzYxPJHq6/NsdF
aHLD/QUei/FBO0RV6uTHCmOGmIEMwquvgPx99zeQ8MPwVRIqfEbiLaOOXoBqQ4v6
Idv1qf55fEAYyPn9Rtigj6ydytMoGtUmaQHdoU4Xa9U5Jl2ul7DMJ73Xv1E3QsR5
7TofjtgXLyrA0u542b7cV2V14Ldyt1p9HisqaUo4P9sAp7WhpL3U5lk5/Xqaiqr0
pMAjyLBjgFQKfhzRRB/ZM3B6czXrMMHCzQvIKKkEItWRqfjrbAIuhe+I2d3Q9ECv
5mlCsYBoKRwsEPo8Vb28mpz3YKqolfBBJVBp8LUig2Wu9G2nYN6FiLsKSaP6Szxy
08FJ269VmMIwoAGDtkmZVinA63VA9R5Xl0nrToL/jsULHCflKwxYDNqzcMdYfQQn
XodnsyWnYBeYimA76F4td969uSflnzmFHbG+BuLEmm5vKR5uKtsoSFWa2zRG/T6x
8gdVkXtMCOvYHEqo7j+sx/+NbYr3/bujoh1WJRYzbjIEiQAFHfzSs7BwNRS5Qhsm
RtWD5p88bPaLVC2qSpQugz+vKz3pvt58YDnS/9L8SoBmmXekSmts1nczqz+2g92T
iiu96teald03aR03rM1ofv8fO6IBWxcEWrXL6XBfGBpfY79bl1it2WsF9Eeu9/UE
ipUqclJ9XE78KL21re4ei+VBRHQtSt/51up0x3Rp1G9yvIy0/DZZdXUvQwUYZUhs
EZC3rOnDQDKo8bRfJY6JAE9pwL4UtmfQEqFbD6F+QNMbiSa5ha8WqVDWrsDE2XAT
wkxetFS/k1NAzEeZWPwoC1OqKApa9h1TkfJqGQun4Um4y1Yo8PwVonOAM56Pw9cf
NSpRZA1vl5L4/gPCONeKnCpBJuQ+mYsQv75dEuzFdCOQ2BLH36bK2ZVJGAxab06d
qNnbxcfJN9twjIcLtydYGbDcQB20xpmRypxdhzECx1sPO+15l5GV2mGWxve5Ejaj
1gWoGmHv7w2lfpdE+mbRQDMPowefzdTkAlDniTVT44u236bgVakW/ZvfU3msYknT
vpJA5VXSFDL0kyiaCvAEeUNEcfV41lF6Eanw9EK0k2BpF3TcQSzs82aNjA/p28IB
EUULH+rW64lrvnlimvE6MnLgDom8spRRAF7oUWFgl2O7TW8K+iY6n+CVKBs8YNYx
JEeXjqsdU6TeAVS4+VQnwFq5AoYt1/4Jf4hIiEniZ9NzlHnrU6YLD/Me6P9gpUqQ
7PPx+sQpEP0t5QTzIVoEfNgdnHgF4Q92sxd7zJ0WeSk/ZO5Ma6ha67Vc/82LPzcX
BNasTubsTMijvVBabJpQvkgF+FIf+Q4GlS77Bru2DbUnqiHxLUFZRz1KSFU5734P
+0FLIIlcs/azH+KC/tS1TbrWyyjLOq1AWIEqUNfMcQ63q8Gs14gZpsB3WwI7dceS
js/yEg4z0d1gPP7oN5QvbrbT7atHScxksLdQM1hxXW7oB1dDjKOW4L3l5vkmO7Gc
76jYB7sMFFCMWJPgXUInsyUvXYENnqB3i26pRELy0tIUMrGFylnxGmmEstWvmUZT
PhXo9pROgSj5fZF8jJGLzSXfv+P3aMn/SFi4QW8CY3AIF+/tg1l1e2UuZySY/Vz3
PaRXb+9xnS/4RJr/i5JAbQ3mWtcsADQJ/l2swxgT4nx3Z1LLDBnYj1BTPxUBXcb1
lUMnMwGzlf+b8ZTWbRSw8Uj0K7fHdLRnNx7U2f936mUnLOH7ArCpH0cK2ZKuL4j6
DtI7Z0T+l2MKWhskA4wlf+FTTSvz3hblRT6KhsDOrkf0UEigolMY0qhatlYDrkKw
Q4XG2+qzFp1oAbsH1O6VrM+Z5EUjHGf8krG9zQgWruWOBMmnDGV/BhVsfvmb41SI
l81WjDvmTnYjCmFJ4xdibmPaAMVITJsZa60JHRXoFcJ/863jYMLJq2R/2qd9Dv0q
nLgGPoPWjQpDd99/fnTn6dVIL6iLD8WGfcqclcep4gJtV6YKBF1DDRCs3gmSFpdZ
5828H55P+UBbAEDWfYDJN0Gz+xw6Irm7WAwhO5uL/6w7OGICtm9t+4thP5sc9b6s
5OY43Z2VZqGZhD5QfRGE9cTny6Ca+sngXx1ysZqKc9YhfSotbiocuY0hgXTVy1kW
r7ktMbT6MbAaAPrkKSINIlw0eRyDRClxAb1UOzWDIYrDmjr/jQxf3G4vggM7ayho
Ms0yIuaRmNGhzHAWRVQe1qEs/78uhGPKn6uHQ0ejriNtJzqOWfQft2GoID6KdHKC
WUxtt842zb0k63gCnFhcYcIEAzZeXXrTEr2ZKBk8Uke1gyh2EXYeWdefZglvRzjn
Rd23gO7+UaLzBqExabRRNhAw+2lCQrf7Ib37swnhg+U2RjKuGsVc6oi6w6w/cR/+
FrQKKhQxAL61bhMEtX7wHGhGBjenws5cWUi6ygrAcbRYLPjlYX04sK727on1YhlR
caye+H8PvB5wjq8WKGWs/V0kgWCjJ5FM6fRYfrHzqLeIQkcx1PwxD3d7MaXVSmvi
f5icwtV25Lxek7+tdyNwJebmmW91PiuIVy3wS8VnxmQfM+0OrrWkTFAqgh+gPpge
GNRKHVd+UgKKd6ZVM/is2BV9kFrw2GbVUbs1HJ5/X5iOaD9anmtzPdIAeoAC80FM
iPXB8b6S0WfZ5iYdNVnqK63ce2QM/Y90hj4zgN59X4DIG7vgXk7Um3qzCwKs7WG/
drqEK/SoJUnGGaG+0+pDQvdHCmL1T9yTSzf9Rsbu3wzDs0HSDyxGWGD4c/gUMrzo
1rtxve8V8jAM9XXaG0SI28WRxtxC2nweKjt5eCA8eCSXn+Ungr1sy+F2YarMLVCz
ySQ+RrXGcWzmmQD+u9JwT3WtU6wbgSaDmciWxdATe1Tvj6WPNm0bNs5WpL307clD
l+iVC2LwEThR2tbjs39kLlFbyNOC2luCHhkK4W4pLFxvfQ+WZRcQfaiHSme3hxnR
YaCo1lOj7SWoSRTrrzhdkMXMM7MzFSiHck008yBSlfhHAD4R5n/0/nRICv6iPkJ8
rCJZ1gOylwGteBKHfLeemRAbxIyUoE5ZyHy0MeunReyiYRkvfk01vHVXeXK3OoYH
oXJPnzQjnkvFVHOFXPcq3wmOgARqLKNqhrIH09B7llVO0vjT9ZG3lOq/3aC+gSEt
uvFmuMCyjqtX+MYijBPQGbmIPi62rvvtuN7kzojvpd/cmJtT+ee69g5g/1ddZzh8
fCljrZAIrj8XBaN2RNFzD16Q3lxTNg/tGr3hzStKb1r7ME3hCvzKNSj0QiSf68cq
cj2jXjirg0IgZYBfpMWykAAbXdbMzHaK5XNJWirBNcbgzLsTJJtBp0yOWHmGey7+
+QiPMqUPcwmdqVK90WYo3y+Dbubfff3KMd1PNFCbgunkPsdcVI/xMqoJ+clJsL8O
c5LKIyty8pvrUVAISJ8ZZwp61ZvVNn5VPch08p2A32k14BRX2yyXw3Z4wuqHJYUl
c2vs+fr1xa1Pr1H56SYYbpy3Whfrv1cGGSRzlTXM6h4hFodQ9VzDg1n5K78F34dy
opeZft8ZTjJ3OM7mXl3YDSa798Qx49hLwC+67II/a+0I4qpj9ygSWNCWmY/Qg/pO
K3KXmJuC3qqTPRYBRkTXyizIjsEthAMpTeoWnqGNXVaAvX4z0UA75/NXlrgq2Ljw
bU8XZXlxOktrJgKq7E8ymFFaWn5s/vS95BzT8u7/FWgkcwHaor/s2OSXwGbAP1Yz
3fFJAqSlZbhmAImTV22Z8Xe4cy8ymeeh5zzAhmkqyCaQtTDB1/5Kxw/B1tpDzZ7v
BQ3Bp1Ar7kHJDsdbUcI9qZQto1IpiUvEbYbJQ6C55gwjj1RqdG1WiVmGdmKNj3Ps
8nKz+wlBtqfkRkA7HGZZvW5ssgyB33h/MMOBAW7p/JduufPnWKj1jnOr7rPwc/Mx
tOf7qivCKIdEdExymSGsncbD6nwK0u/Wj6ZOLJRP71gf3g6db9UvYtVxgE0ZNSkn
vN2QziJGo4vWWK6GOOYu0BgbX1MeJIW2HhmOXBD+HcvjIPT9G7y62O1tsMfGPZtk
R6xZetC87qsjKSYVpnQRZt+hRJGhibxDgp6dXe6kqUzUtLbS6CFQNxpW1Ua/mCFf
lR3eqUdBHfkxl4dd1drcKjobVv/vEaE/g5XQkp02RfxaQSaMv2xjeZqKTWJeGm+m
+NWbQ+ETNsdbfUsUCDygnOr+6AEfE/cSAM5Z9cLsw0w+kRFJEu6BedwXID5QWSQD
J9OEc9mgaOyCUYNhjceN1YuW8sdim+RLBar2uWgOVjsA2KAC9WlIUv42VEAD1SgP
p8jnc9o7tuJYo2cQOrz+7zBG2qsf7GsB6w1zJplITdZOguMorLSZPMa2kbeSglTy
ojyRs72ZMGkbogK+pPBYNp+xsCep6xQ86g5mX5Aj14gqAJggp/3XebHFMD1AIwEg
W+CUonzhp4cRGFgmfLAOVJ7ld7sVDxn9wk7dOmYRtm9WGonFhdHhmS0LFC63ogot
tyXfyn7cF3VXngH+YzRuXd8AvhcvepEtXvp1Dabpbkhn/5r1emrONQ4xLIwJccsO
7JZmRHQmEmDQd1BFTw0LS6NO16E5bna/gIDAqP0OdYtVpZqonu+1Q7/CftNN5E4g
y/sw/2kQwjOE0we6H4dS1Gli/hJNKGCp0FKd5zmDHfJ+izB3xVGt50Efmg1rfJhl
SF1FYSbCTpjYZwBsHyKAL7hXH2hcTc4HSSZVNkVPIMpl1Ce+/6QAyMCCfA5f3ve9
raQ1yja45RpK8kynzU7jDG16dpjWnZP7UCyaLzmLagApUHHER0WaZ2D90EhSkDmc
VyOkyar1Sn/rKRDD1ChJvxpNbCWP8ow+iCLNwGreQR+kVPg4G2xOPJbFbsLALDn/
8n/zyQKG1chvuJoOKhJrrBRw+UMvF8hcEMRt9to9+okrbTzAlZl8kICqe/s4SDSk
1RLxbKwHgwjIAN0gGWnkaYZqFn8an5TjaoojdLx/o/oMdhHp2q5r+TNc+bjJQuVZ
1yx60XWraH+Sewqf0hxM8hay50i3Bqz3jHmM3kz4BIlV/iLTAoWCG591dOg+vC7J
MaVmOiY/alLnktdhqvj4PLgT75KSziP2nc8TMnFv8IlaXYSdK/ac12dkoCkMpSRq
ucTPN+RayX78woN/D5axqP5pRV5pWGpLXjvlWX2u98GcCjO/TC9stySAoBFOhL5B
chI7pSSus5YHDo0oVEtqkTacRLIxO+2cAPZtbJYAgiIDNVHpVqUWn8xa1lUiHFzW
xMBrHEwokoRR0knKjqeRCJZK/GSIIPVo/CMANMmpoFlo+gbpGQbnKn+uq5AtlECE
ZcgKDZfJcDzGwmupmAiYlIOWXG0p+JvUkVFJVRAHFyiphxZyMvL2F0hLNbcytbX+
ZzAO/JyJoIU5uAZ1OAQzhbfTxW+1nykEihLBhID8/AcVR33T3ZG9b+804Gf+FY2U
R9vKF8bi2feBtctWjxHY42zMyzllg/VZqIr0gb6sX88WrSs3FxT2dOVEdBXEk8GH
Erlt3gfLYZEQqvppPIprRyxCSkmv1y6L9Iu6//LPQAJtnmatYUpwHD4pejeK0WVb
ZmslcJlHpcUSFz7XDO6oJN05+e+icGknZaCnYMTvhM35Z6S1Yzgv+q8JyTz1qUbS
O2Je0+LtzgyMWq6hclmFKFc8XXRrnl5OX2drboiQUEJ1tc7X7S0owX66CMoaw6t3
s1QMybjb+Q7nGKyKoDMgzGPTVTjAcQDndqtfDY08F6gsdXaNxNfuqyO5RbelS612
nsmZDTXOnq5yFizdG90hNrY3eOpRI/G0EI5W+Fst2W0GzTLm5q+ODQtR40dzYjc1
x4nehAfHuMUMFr3MH7+BPrJ43hOv7MY07g6u4vxMbVxFnF/j18BTViBn4zHfbxpy
zDYH2zE8vjb/4qHbYS+3kZW/7ecTGnmmh4uMNCtiKJb0n8McMUFqb656rOiRXEVw
psIKr1y2orfNCjDRL5YjQKKcaj3DKTcU8aulGsCme7xMkrcpXQIcOrvYr2SRhbCt
ITt1v6h+56gwT+n36XiEC/xRuKvkPqLbN23zfXzUlTl27Qh9HHfmpBCWfkDiET5X
Wea/VVQnHh59hTNKAMJXfluBJHYAa9UOaKGX9HNXx4DNxOLQ0WWX2Krm8qjC4e0c
+xYEWxrK0/Y2n3FQulMCi0hjkxulgSXsXymfyIvFIYI+WQajy1+GWQlM6KTqQweO
c4f7Ky1pDL8U+Mymav2qqp24dtVN0Cy+05DRBd94FU9UE3RrBvgnWDwYLb9k7eVo
KK1Xygrab5sN7B1F7XnrCeuyUUoA9ncv0YGOKphDC6av3IYlwwmrzJuIMGrXm9uw
/kot97cvIR3NJGsHf7O1YIUIBE5h+PKo5UKZkKtmW04dUB/d3JkbtSi0NHdJKIiy
ldxuoXU1Wjf0dzMTWMIbn1KwhuhVvqRHkR44xtB8jZ0b+pGHY8iz2xm4qiFKAVmP
E0RqL8gBJAAYNUbdpyKK1+/D+LE8PPgRG9Besw7TMO7utqQEkUvkttB/6tbh1t+2
bx/s4bL18SdJ0HV0dtmyWjbr584BZm6HV459+cY6XthlqgqjPc23CNvugFhxlwA4
66qgmSY2oAxryxMCKxF5aDqyVAcUZ/AjDX+W3ZNNFKZXdvENn0wZlH+PhUVMQhP8
CHvgG9F2Xy9vzsbnA6+oFFjER2JgX5JumiPxEg1GxDPwgIzKbgSEzO/kfI3HDBLn
onCFelCbXfIPHCq+LAQDuPvUxLiyUkb8crReDINejNUsA2ulwHihTDmkL+WumneV
`protect END_PROTECTED
