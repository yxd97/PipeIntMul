`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94IOpdg7rWYFZuTqG67hYoExbWpduTVqEABB3xooM0AbXojpB67Je+u5M0LqOAK7
6oHrO98B8VD0ug5OJdHmX1F8IQWHxtOxdc6/pBlbOrdb8/0V6CjxykrBdPdZHtfK
+4zkBRapslYunPjWveAOvXmkqwKQp3f+PsRwwNtKpNCTr4mVTcTWndA6419kTPnB
oiq3ejJiC0HspH+zfNsdVELALKXGtAexuEuQzpuBj0s+NbDz33Mc/Jd9a/4rAAbB
E9fMGiati3ctOaQx2Zcgrcctv8OGz6FupQVqOAYuTJUe2IsF3UwuJcJV8hx28WlI
Lyti7DqNJjpElwlYJWPPEtWVIm1B/3Prok60YTdLar5ErgWd7u8no7hyNRXv4R9G
uKVaiHDkQ8/oe/94CRV0Eq3GXqKruTCU+rkOS4qlixJ6KBNMB0b2CFCadz/xl7pv
Y+8C2U691dwIsRmtvGSnX3z39b4MwIUanBEufSp1D6fr4yWKb2SpaYKmPTCjt/He
7HyIUTheePa6cU9yJAk/ZQ==
`protect END_PROTECTED
