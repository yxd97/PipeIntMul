`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCzbooJxFNYVqHK+gFOEQH7Ul64EM4OFEXi+NQ1dkSiYWsJWZubs993QbQq4TuLV
U/y68LVrMtfh7DgN2UIEPykmrbc7AB7lC3IsEzo3u/Fzz1NhvaXEzw8Ipq9WIlH/
f4jD4L9DmnHopg9MI8Rt7Gz3amYpz5tF0K/GMVM2IxE3Cx5uZWGBbL5Bz98FxQyg
Z0Ti/VchLlRD3+N3agCE5YJZteWAuTsU0K0giW2RWf2dLKUmOlB7dzLv61CdwlMG
lI8l7txqK4cQ3ibqYLOKNARsVeqb4CwkO6cUHJrICmx+YKRdbJAGVVrlP5L84Frw
VVz2xiScaga/CAkbn704uebLX8awuSzvtGatKWGCr7A=
`protect END_PROTECTED
