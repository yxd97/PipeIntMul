`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dra/BEM+gIXs21mSTLDXZh6giRqdHNZqshlbfZMvxPje5FIKfHpGODBSKUk01/k+
s7YKBMlNFHkqTMNbfHwyDVn4rnnVKoL1/BMA7W9iT3995JP1KgFeYqTBy3Og1NIq
JzbZYzmlK0eKM9OqAkBjN/UG7LkEVqW9iEfSvUfRb7XX/BGG73ZjgSiR1FUONIVp
3djWwaC+vRVbtHsA/F5QIRWqHbR9Cl4A1qcMVKID8AARYG4Sa/p12QZRj/chAEh4
gnpFaufT0nHzEJJloMNRmbR8QGbuNsY8UmLedhT/293+osSFiUhLp6XBJxN+pWig
e1PrjRp0fnmfxDbp4uvjIiK07usAkeon4wBztD0De3No7y9BbDHRUbdYLdJoo6Ra
uoovkIyaXwOalUdmlzfeQqfuCMPxqEHKCXpFnK7+QAU=
`protect END_PROTECTED
