`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1vZsCbTJud6U3okvs5AlpTgkdvKJ6JDWYW8WSL7k7zGY7Jn8kMOog0YJBjOWnPz
SCx3gxOkdZzU+sd2pJ+kxnHGfI8Fh+j2UsxTKKVVBB2h8PPUrG/hTIvbIhFkQKVl
GXK2Fi1akMxztHb2Nn78S97tNLIXPuZ++sPBRC+bhfgN9hb98OUEn8YcfdMorwut
hi33ilJNc5LJy04XEQX5+HUf9APwX0ev19fLqRWff2f4g+Nq9DGz2llwuwUeLSza
6xxB/V/D/tqPPuO0J2JsuVzhHR+quN+ke3JCqn3ePi9j62ksg5BWuEjZ26PhKjTI
5YJC1ZLbujC0Q/cUaz83U4WcStyKGj+LDhMNr6VmQoNFmhYArJH37t9AWHA2HEXJ
2++8OwuatbvpO61qdSpCvvtJGvAfR5HL2ZjR7Jc32WaAYMZ87L4vWOFECpDJjhLr
cPExHxUrISUZUM1lm07j5ql/Q8Saao9viaiuEZKNRP8aczvsE2L1E36mJ/68PvEp
pbiLHP1Jg4dWqzlsYe6NqDxSSKFBufETRcTIVVQWgKcOzUlkAxsd4AD+08ejvnrw
yUdsoFCawL6sRB1r2d90H3S6JRAt4TjU5wanRWNspK6Un62q54hBrFODhVQWTxei
knE0h7BZOtmZ1xcaadPupzkV6rdeigUBauX1wKuIlhUeN5sTjWyrwtVbj7sicEbz
W6w/Ln03hKhC9GtqyxA+LJoCDk1b57zTxqouvBU2rv/aSkFhtuIVGW1N1WqByxh0
`protect END_PROTECTED
