`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6VzPutCtzSj5vEJ9NS9ISE6V9NFPgyayOcsasVV3j/X5mE8MeMBKyEzC/iDw2J4v
Tqiup++0HWpTE7ZhwHpfzcn9RPbZobmwqsnT7G4arQJchtxIKqklCnnJhC/ZXry7
gcmSmsxxySYKe+Q7XZbVODVNeMphtrdj4kxbtZiLoHsX6jZcdl91v63FHP48VL/j
EdrdDTOuark3PKluvBq6NC1rsh4dTNC+BNS1LeGxZSWf7YFl3j8wNr7cQEHiWB4x
CAw10w7CO9TqvmsQizrQzIfb83Z1YjXTAwQU7F3uAHm4xnPOoivTSw9V+QEsnZ15
Th3Qb2E8rl2OgU5RaxKR+NWJ8LkKFGgh+Tnxz++V+yVHNqXHaKW4gyzf2cnCzkRU
mQs8pIorolFJ92x4xPVNGCEZr1cXrbez9qZJLwaP7niyZ9nuo6PmnsOXFYh1JasB
MbzXuLwl6phbaxT3BDDhUhzKRtEFoSWeQ3BhYz0ypmAtLBOf77wAUvj8WsqUF7i+
rGEsqP8iRsATzlRmxOyodK8svXHNbGtK1Ip/+QVCYEgwGfBU7zQqRhrLJne3M76v
wxTkvTKWIEaI+1pY6ZVyQWdpAVb40+oVZG5o7xKsjEch7R1Ati557An6EI5jKo0i
NiK298Intv1lXZjfmPaN5+V8QLBeYJUslRa5HYlwh3CRnML6hJY/aXAuEO2Nq1uB
KRCdS9iG0TyHF6lxcn3qxAhjcamjCy++SZPcoSdhEB0LlqH3pmKO2feEByDu4CDO
JcdcjCuqP+ebaeJzz4lG2Rl3wUueD62ARMCcjEqBWgPLb/nxvZxMuyjWYjUxllj1
GLkcgFNdtoxx0QgO3nMRAidPu32HO3siacR48mqnHOknDWMrE1bYF1ZaSLIH1q26
iGTziI2eUcE/86pR1auQKQkhc9oboZQzl1ih1DdxOKu3Fj3jgDJWZFo94sAhQw+K
JbJoDBfPPESxnVKOx5RBnI+s6lJ4xKzNGdpebdXWApJSnWVvZK6gb7jhvpq8q9m/
pQtxcXrg0miQoeIQLVVpZzgoreAwwI93539xZQ2X+8T904yPS3HibNG5sw6HZJS1
ACNqt9KDZT8tzWyHf4ZNNQ5YZ+0tqpbcbl/ci2sDRssO/G5ruOi70CpuowRFvMP+
JeUP/mYfmU0xuFA11qa1A1UcOp0nMRZSVVQmFVy2T7wqY4sZsyZUhNHiN5G0sg3w
XxhxAf5z/QwcTDWuYFbFsxN1MCeaypLhxcpxls6qRiwl/dKhN7TxOc4KQxLRk2cB
3fqKmZDzqP8obOuoGWHUajuQygvydMsilH5C2PY9tUaENmNcLvWXTAkYVPPhQOI/
Mo407ygT2+AbmG55tuE0jOLOrh8ViOi5vX8tba0to3byiDNI5wqIQYtzs7ILHH+Z
IKJrBlyrLxOEERD3Z12f9xygjzK/BAZZ+IOv61HGvYpzXitl30egOMsGyUqEXY1U
1+ZEAzKElPS2wOdLK0NvOFP577C5YJjXNRNPiEOJzPbtUbv1SIUSGXi2neaFBYqV
86IwbgNKi6Ws69YUC3/BV4f/ZmF09EK/l7ddyGCA6WxbQEdaL9ucQkZduIgrOXHc
KkAurN2qYmG6B5475MMeZ1kgG3kvRk9wXHQA8XrW4vGR27BkP0Ktd2lk47XZM2vz
dbAuvbAcXOrLOLETql8mkUMxDkhL27xOQsgDw5HBEc5GNZEgsGXZ5Yc2G6iTGaKU
av46DqrTgoGpHEqZMAxYEZtDNsONFc6+r9g+0q7m2C+BEFkD3yoszo07l//2h+Od
8ReV91eyAs1VtBIM7PiqVaPf34Mf5AR4pVUC1fZIjrtu/uYgOGzHdNlx5dqr0Vcr
C3KueS08dMVxHGCgGLmZxd9CyqjPV5TbqRn9PpjiUG/Mm3FQAvVKV1X3uUO1lodW
KKJMA7JHT23co4wD9urfnLkvvX9sLaFbSE6NsGqdv92kgJcmAq88pE1nxoQXAnXh
1gSlW9pFRb/7UqR+91yQEZw22Kh/rcgLybXlEfTG5rNwcRU1RaOnR60HLHuiekBQ
BOpSG2+Kafd2M9tnaPYQyWssc69o2jz2WYcGSsoQCwq9O/2LdEFCYcxWWcX/KJGG
k8QUGDT5D5lYzPuVdXLEE0Fk9QifU72iilFOPWtUUL6I/y57uFOXukBv06huPbMC
iM8BF6obUvWnl1/nLRGyjZVeZQpB1VY2XcKznWcX2HLqYI39AcBOijCgyjo2O2yH
hxMPiTSYGgP54vrb76lnk/kFXzLKr4ED2GKl8mJ0HgVqB74i/Mg1z0ZXyZD+keGK
OIz3jIFiiL/2leiLGo1Q040G8ONlpJkooTM7iFX+sd8haa+MIX859pP/YbnHNojI
PPxfPplQfXbXSiqgA5nVehcJEN/igcMPuQFGD6Gk5vxi5LtgvwVe+YoqLEBGngqi
DZCzMEpqBL45x8+TLD22/tzP0s9jb+oc3b5I+qNMCT4DbD8JqzE+HhAIiRy5B6uW
NbgtkjEcGBgNXdlsCFdGzUdTc9X9WNvhJl76nFG3HWhlBhTisLn3XYltvCxJqw1V
kwB9oZ7SIoHhg5hzNgL5nduNvxkFzLUBdFZUS4ChLBqK2udYmCY7zWunhVGo1W/J
QUAHyGlC2fUGxG10hrPirluISmrJcRQuAjXOc8tptF4vC4gTYgWFmUntOhN6SxO8
hkVeugvulSclbgsDjhYA7EKC4d3hyXVpFNtNERbiMxE/sUslMll0F0jykEDnOu2u
8ydbFiPw1oHx/qA0vEmbAOtwo8Apa9EOk64idP1TIWYbzRl3Ik813Hrnauy1ZZKp
z71aN+QiQ5iGBJAxbWn2WUz5wKWb3UQUcrn682tomkAUonEREAbmmC5TMqprW2xK
hbVgqE9pAf5b2lsYTJC3eudby71dvw3csE0jqnQ3aqxPFtEAvAJXuQjwnFxD4+dY
wMB3oMSoIaOYN9EVW2seb26RsQSm8pJq/6nIVukno5+C2bVK80ukPH0GIK5iDMGp
w5R6PY1hzRG/mN6c217emfI/cppKL2McUZ/SBFva7i49NqRsX8NX2TPpoa3w1lna
32c63hEb5dO+A6N5Aytizfx0ALDv8DjzNoowQYzEbqGtT7MRgsCfUJHAR84fiBUA
uEBYmpE5eOkkLt8jioknzkWloEkRGSw1QkSkfp5HpOPPvaR5LUp0B9PWG00xxKS/
gJY2nmuVHbjFYgVl613rtbojJJuCESXfDDGrczJctGB216peYLGSPd9zJzs8i7Dp
O9nvCZrw5dDcrbZWDVHu9MJeRmTYMDBacOkv+/CHq/DzhrTuiYAuifbJd5S7o9Ng
y0i3y75cuCFij9hiC0n8FAuRDABXrL2eIZQc58ETcrHgHIrtZoOJgQ+qRhXTfwFL
3RDfOpX6SlFpe8Z6lCo1AT7cpDdqmDMMBnst2bntladd9mvEAbbWSWKCI9d/jdca
ozqBNZ/4jPCMMjGGRSOZGTQcA+sy5YN3jopIZX+4s1k7Y2oakiPAbNcsROws8Tq6
HuKJSixBX7luSyJrnIPGVwVLWoDLVCCcUiHKPuZR/HZUaKu1pKW4Kni+X22TLqMR
9U+vWc/WBHA80Rdc9KeK+KW7YbL+GB7cdi26zKg1Y0NWIVycKwcTDCQptunNWOCA
h1jYj5hWxhMAbKjm8EKQJpKXUwvGEuqU6Z6JPTSo0T1Rm3QjCQW+RnwseRIPaQcs
9IeNosIWsCGcLj9B0qnwUqibhrlnVT2LJOQg5tSiOYkorBdc3a7KMN/JybxHIsyT
1ImwontTHu8FipFRTsizdqfDRkdXYYyWmn5kdB410z2KAV/13MoNPoDPLMZ9WBS3
QzEi4So7z3DXKCCvXrO0iItyHQHNdrC4whRCbnhOqvmHUxmjlGhy9oRQ/Qm0KUrq
4WEbLBguwiepExFpdwYSxHn0PeYzDCtTCfuuGwTfLMbKVMhHquEG1QOHEJi3UBSx
DFFcn5L8fS1MYNoygbGFiFu58TKFRxygGZdsOjD1xywuBwz1wi9Au9c2DHBeuSZ/
5iWSjf4iDGMcx0CRzKMODeo6tbJEx2B9pYZD1EUiRZ78Qo54qI+apsUIm9Uyu+p+
u+gkxcK2CSSUNnJNhbWxJskEHImoh6C//CJQhlzFyWP4gSWtiQKJQhA/KWC5k8U1
Mu+y9LXnGzLMBs6qXj98hing5gjuBdmuF9nh3NkJiDRuwv7W0+MS+e//OdcYAUqV
qFHQmdd7GyeuQdXDBUS4uERejsWsJHN02liQMweNg3QdiqeVuCH4PFcnye1LO291
PLg/rFQZjWY+S6Q/DUGYnjBxknTWSaUrvpzz+FeUCtkMbNUODeNeLRvHVSYq7eN/
NJNyPw1Kh5RJkS3Dsh3myXSjE+xXCAuhk2rTd+Pw7HQw8w4QfN927wvwbosnUfIe
GisLY3Nt8Noxa6H6djHgiPp8hXcDG2zovPiANq1juZcPgYQIel6M4w4JFJIIc8nU
WSFlI9AUBrOOVOK3EW3Bjji8x3yPlytEoO3hLdObS0E1TZAnLU8ImJbRFoxssXYJ
MgwEb3yY9jztZSUsQA9kMA6by208dpuQnOASaVoVnEvdPlSA/O+yo8eMcak3YkmN
JB8D6qxV5YIAuutxbZ7h90fATKnkb4v0P95P2i8XCc1waW0dC9NUwBDTpuG8z4Df
fZRcLtIcLRCMBk4Tk4VgjrLNAIqtr/ytTTt2GctAfwyeQr5Vql29Xeg5DI11igt2
R3zVxoe05XqxbV/9pQRl381MXXEksm5LKBjWaBqclnybYpXzBrZ4UmPZxR6Kn89/
Vw4sWnSN82EMC68NsMo4tTAv+L9XOfSAB+OZgqItMRhHLKLcDYA8QzeF9mRqfHkP
P5uv8A7dQMN0Q4pkNcpitlcn1P2UzTKOzQGjdpZPJ/p9m9rDzySvxRIHZ1gqyG6Y
MPDGrNxi2fGAyWM97xqHQ8PBA0vnb8tQO3s0jy6/c+jHB0kVL93A2DQi+KPaQPDd
egJFlPS+fGpWvQC/6i4v/H4E+XtRvEPqzcv3OTByTxTRLevctAX9d4RwEpxXv2Rm
XuFvGl04t/CAAVFeOyhRQ6m/CKb/fQpz8Z0Zp/lsC2/xatgpuMI1Bd7XK4El1Otq
ptAwditvCY2N+x+wjgA4ttDusJ0QOpcn7K3EhCNilKGGaiKzDQGwabjZIL3RQo/z
zZ99T4WuC0TDuSshvhOZJevmiQJKvnEDwbDJYwgtml/nVH2nGxKYGK/MN/5ULr5l
QfWPvrhR5JhCjB8QahazAxL0D48r9hjxfhFm1t74LJ+SiuxCIrvZTMb+OUAtcbxR
nDOUvcHjd17mN3aR5iPGBZOPRXFTSdyz/QXkeD0qFMBgS/0hRctWbS3yXPiuwvKH
iFvn3n0HMSUvq4PgTewurxa0ReJSJysAdyUVcHgqq+RjU6SprRPLjdm/bgKxnc01
xPz6AUl1KZP5o2TdXCBKN2eI0cv/7ij9qiFvvnivfnCRoKjwFBCPI6UvCAkMUTL8
WkWj1T0ScG3x8EFUEQPyINPsIUA6oaqt0hPXKfVuqlibMpYhDHUAGDDksXQDe+4S
IxgwPe/N58wTXgmSc0sgFZhEfJWHuRGBt7bz/JCx+eQ0kOmf5zoUFC65A3ciXDiW
z+9Z12ts7xuMFsbGIoOCmzfAJrNPE9wdvy03iae1PQkIEOsVpzznvAbrRuasjoIu
22IG+ICatIwQ1rQlDuQlc3wDDFAWSXfNoOD/OHy53J50jjI0oA+0xAiUaw6Kh/jU
THVyMX/Qo740Wf76ckO7ViWP8530PFkgA+YDEAsFzkxGYXczKW7UA76ZL+HqPCjX
gCxO69GKlZEcm2ry9vIB/H1GH9Q6Cf1oZCcOQ1zBNVXYf+iK2TUFkdi9d7Q3Su+j
UuexzHhHKK1j1mjfz+YE0WADYXjXMk+geIW1uvnk8vxBKgFcDiiM7AZrJuSt3IPw
+UIrcD/ks5o6jy87p1HTxWHUj3RGMalGqehWhitFEufg+sfM93W2iVg8FGNn57CB
lnuf1PDtBsZ8I1I3QuwGazDykqjzChePk9z9Jo4bkK2n3G1ete68q4O9BtixJB5K
WGUcMjV/iHrlboKP9C7YJN+AMzTTIY5lDrqKIpwfLjwY/MrRAkr/v7bx1H0QXjcE
zdkYzIsk+8sIVE+6FWh3jyXP0U0QAJTuLy0vKfOEkzPsxUVOjPHATRcVIhRNKST5
hI84IfE0OOE5yxrcXDqT1bITanHYZt+BSzvO+FYULwCA0MXwMblUwaCQBkE6JCJq
Jzh79oeJS3jVaM4wpx2ld0q0hgTB9NoZi4nIxyayxnM8vZmMCJn8PTG3bbpPq0qa
7s7aL0wud004FvlEQVA1yfOT3NYNWDFz7zIJ/ztUHvLQgcaXOipwyibS9BKhVXoF
PLAU/2xCRqXlv4eeH7t70CLoHjRH+ONsryNPgDU3Yw6GsqGbSixCm/YJXhHotwZ3
Exo199oeklCIYaUfJPcOgdi22euaWMQx3n0aCtS5BBirqF+VzyAyvPBIkGtsHmz2
Z+dusE/r5q5OQdGjd5TDSMHx+c4N8YI55Wr6XDK2mdXA3w6/uulGRDOxzh0SxTPf
Z0teEI+TtR/pZK+0FzZ7sgvCezfSjTFNT38J1javXYuhHxJbZPw5JtOmXMn/Y+qF
ttE5T9LnNJol2u3uSLBBiXLVzKYs+YENFxwngKCrfjWEtnh/h38wIvjE3LH4TScC
cqY8OjU+FS8pKpECteRFEgQkLZ0Bdm9ybPK+X2PPBp/0cP/cerQzoNuon7o2HMhn
XfKCjZLMuaI2H4tybHyRkZuIWPCjPF9apY5gBiPmhLNSiZdGqk9wp/xKDEP6sGQX
QskFo+QQKNQIwPTmMU8frulB9q4K6SAg/FiM4PXlDBcVoWXkSEOwC4ReNdM5hNkE
bKToTncxeZq0QadXZGDxM9oXo3nOlHzHHOkWa3uPOyYR5IUkHWcIb3T6vHBV0IDI
GMUllm9MMinBHrt4EWats61Kp6U6of8yV1hQIHlyV1OBSCdgk3THOcmsuLaO/j+0
xx2yoeME4rXQmW3+27HtfDHfvLrkN+4tBDTkKu3D6EsChqgBzmAG5wSG3jx4sie8
HjRzouTN47PerxUBMni3+DGSOITmQsvxAj7OAOO1yEbngPqcCuBFwoTP1bAIFRcG
GWpSnwascJl+SY39473ayvgsNCUZX1jwqjVc9T3RVp14gjpg9yykFiHijKXIP83q
uUenOWAQ/LPhTe2kXXoUUWMQdsN/KNEYyuT/NG80P5mRVMppH7fVEBm9JOw/ZN6/
5a7HMsr9MZkTJkciehOmMriL4QLuXXMmAE7aG24dW5a0eofc1p63o0VDt0ExzoLX
QWVnHUhPyjl/wid9swJFg4ncTTHIIwS5M5VA7M/Xxgv7K/GI6/WlUvn1nYR42jcW
HlYU4HfQwk3WGr4GKhvsdUoNOKKi42cCAs4TImk2sDe8nMCG+m14KyD4Tp9vM1HZ
ngH97sINrt24e309EZl6FdvXrplQ2J6N3Ib0bNMCDOrQ03NLoL6dVuO6hEMOEtGN
sibkbOS+xwc/gqY0Gx9GKpxKoSwrm3zWB/mCyCcyDW3Wcd2tMj9dh1J9RWL+FVtJ
z+j6FZYqXIQ5/zJCBq46qrXX0HfLpggaWoNnecT4CXYSzdLun3lgYlsVTwAtO2y2
rqOKOeFDndd9Iqt/56NApwUQ2dpTUxs6PlS921jr6/o6AvHn/1FiTBlwTKtjFom6
1DilnpbDOm6ugazR/GyFOkWwpwcd9DDL2bomwxQqYy+QiyyLH2xiBaxBW236oK1v
LJ6IRlT+0BvrY43oeeoPV6QIq15TRKLPP3K2A7MeG5pbx297Oep+m9xkQ+V4NW5z
qBC5kpl9RImpJl1Au0btEQLEeLycnBbXY+Qs2S2O4oT1AgrVlv1RAY5BfjIZ7tmH
yy5XhmlkQGYE84s3Rl/YkJa1AUb7cPTc4i/uokjCOVfIvCvujwTbZugdZwgk8ZV6
wHwp5Vg4XV5248CSIOFf2smHIYtPixnGvpiwO9ubQFz2JGwJSZkI0s2lEzMEoKE6
ZKP1a/fE276uDsvpa2ceTb6oV5Y9RUHumFf/VHzCI/n1KRyeBTWqLWy7aSD4MJX5
KqKZeHphT+1pNg3a2bq9fAzU4noqOTFirK+0fDdjWSMdbc4F0xc+dIRW8lW3fdz6
S6gsflRfiz/oY+asf9ag8REA5Kg80zzmu4r2PIStN64AWaMoeDZUCcjEoMC9ddz2
NdL9S/F2b1mSluV5udJMF85ePlLDwRzgwAamYl6cgFzhMaM6c3RRGNoKNdzObweE
JoNaDAgzNsr47bKqAZIP0gDMQnnHgArx95KGj1eQXdCp6vKdrMrAJhqD4L7Riyp2
XwhL1+dwwTl/bgNbw8fe7bu/wVGBhNt/Y4ziMIL+U/9fmexW2E0BJ/qMVYngqmh8
BdVF5Tc04wka+sBGIYRQ4d1JeFBDFSlwvC5CaTNBcBQEl/oGsKkCkbh71ZyxIDxc
BMbxKKo2lu+HBPlLyN8sdnBrwOn4TJ6Wp0ntsRCeDtc1uit12QOaY2ssRj8o7tH7
27mDoDE2ctBAETPvDfRGmt3pCGhVkdsYZ/xSWvOVyYl2yiA/AXN/EZlPpGyHC2CI
0VhXS4zNJ4OA7RkWGCdUUemZyl6eJxGg7EDgnDrbEWv0zBnA8WldwcKa6CnL8cnC
4bMizyuRKlKBE8px8hqvj1Pf3hvZvZcviq4xJm2q0Q6wjLzFs2wZoQTInC/5BMHm
QsQ1mRSFce3vK7P9ijm0+iiNQyeN431o4AQl7MvdaEwVGDw8JoWVF7JbSq8XpY57
`protect END_PROTECTED
