`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WjjGlY9Aa61MEau8k9Eow5RhNeasOr0SWQvIm5koSMcmqKi66luJ837Ih+61yXMK
x774lLkU485GW1sZVCxJ3jP9J9z5XaRlyHue1zgmPWIMzKoELMxk3ktgXiOlhX2R
M8gNR9dCQjsQpPJPPRF5hozTZgDRYwDi0Rj11EZ8Xks2u2rv8A0/kB7WuaLKoVVm
Lune5nADUVJS1fmjuXSZQAF12h+rbcthoH6kjALDm7fWhrEpN2b6j2zoTjgtKu+x
mnIDz6QAbJYShiHJyBn3N+ptAMbITXKI8g410iCh3XHIQTh/ZZ1WphINN1HX+WBV
n89lldPZAsB/HBkA19T4kSCZdjAuypsG+fpoyQ37TfbUxxb8rTjg7hLa+blwEarY
FhwKYumM/P2DA+Tj0t7SIj5R2Xg9GesCIU2cL1EBXToySXrR78hswVv2K0GwgxDz
0QQI/zlkw1UbiMWwtwsvdEZVwZUoMLfq5X7dWxkIBbm2HSXpLwbKD9PGc4o1cAvC
GuhlRv36sHrmxN15/qaQ6sHtPHHf2dpULzLLatV5qu2wetrkhyFHZKekm5lVGarb
6mvCg5srBwcX1EJbD1iKyDD1Hu6x+M/zzv2niIcNg3m7sf5DKewRxWJipsVvoqtm
8pPFlt8EOtbVD4HShIhG1QpVxVVle1OYvvlDS2Njh0S0tsDtiYNttxjf8e3Ck4UC
kCzELB0TdnHa8VT+yLFrehSh1SfOPGaj9B/C/CPlwvjMaVGvHJS9SbM0YsRBYtci
`protect END_PROTECTED
