`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YsH5EII/yXQTcBHSqgeVTUoMaVo8tdGRr+eHPuLg28eDY+ItxPfCaWh5yedqxnaV
IjypHi4zJo7oFHrNVPtFilDJuwDjR/FQoGYSxPAl0LAt2XTarwahundIe1KicGIP
DImYfK7pH5B9c7HQetQln2sC5y4OG0zApWXRaPKqHSOiciQeYH7fTo5YKSMSTW12
U71w6ddopD9SUkQg9vVrnwOJyhwX75aEYi0QI23zikWj7iX4c5JeIGffyUSSg1xE
5RzjDYsl1rTMhr7MOByfybHUGwKJO1aarBCZAkLO/YZFFfy3YOTQF1qWqlSsZdAV
3D5yBUe8rbEPTYv3aTFzvHOPm9rzzl6DU2K+QRbA3MEnR90HV002MxJvIsAn14Sm
`protect END_PROTECTED
