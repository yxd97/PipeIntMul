`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Sx2HJuPG6QYtC5T9VZfnM7mmSgWeWINfFzkt7Z//VdTheKvuYU+k3TbV4ptXDfl
R80o9E4VbH2BUqDKL4p02YTygu+x5gML4B4ObvLyztQZu/8FVnvZMwKQfYC7uTcY
wlpqiJ1zwEREgY3pSDqHfde2U5qGaqnMcSSp2AvXxP693RCCUKfUtHslrzgK5C68
ZDEc70a2iMfEAULL9LFZDrUbNFZ4gW9m+vBSKUVAsi9YwVjfBwM6NKBSPZDzD0fK
0D3txBkPGfsBrELdgkQnte1Q75NrwtQwfr8Ov9sKSInOETtEs8KX5lu6lBQb8u3J
XBTQyb+YoQ0DFU5wL2JUQoemXUWIt1sKmxTDRxtgZOrtiyQyHzBrL3pDX8erylqJ
jH0ePYRfv6KtVL6SKjIuMcjbrY9h8Z2hDU2mNvuGe6alu0YEZkbxvCGks3rJ62lb
O2vu7rk+Gylwk4auciQE+ajVERJu5+VEfEF91M/2Qx8zBE9ricYiVLMTOI8cHgl6
hP5S7Y3cbpbF9D+tX4l8F5IIYAZKc0SP0EX/F7z2U+lZ1wCDuEwlwhsqwHtR0wzf
b+turyMpMyoZkCJhtCWg8cEZCzHGlrvvzB+ocZDUZDLrinbBGJZfBRmtDPR70LJC
IqVHArjVI9VYDkjyLdBwtlXxofkko2JvOneSF6JpNJAcET5zgIZ+K2cQdlwAkSw+
p8ueBhIowcPjE8d4AqMH+fPjiMK5ylNwHSnkX6KkWV5oJfN1KYAUBVZgSveXwR7b
ZIrHQ5xA9NeeA0fNL7OCVTPGnlTD73hA9e8BnNGAT4BZ/W7eWNwl+wBG+GyE2axS
LG7RUJDc1Q1pC73orRJ+OM3b4I/DVIwNPG1b/0BV3Lp1cbT3x2WpNGkhVatDdjyg
VS69duBB5rLlOJQ/FvDt3A==
`protect END_PROTECTED
