`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFkrxyfT5v/IwXxagX4rUt7ZmwQLweUaWQetwR8E4EveHo8lSWzzpmmh05MzDs1f
iL7lavZBuE36xIClHfG1yQgh2rcHfvh7xpAf71mFPnup6cSa0mS7x6HuDmc4Bef+
JsnWaqfCCesslwWIgOdzbeI/dvDaKiUb6tyHDkrXaNUFf7L5BSaRy0/PWiIcKIz8
IJYPV2bheVpQ5s2SNBlHqWGAKUF1fBO6+bvi4cgjaU9Rxm0SLqXf7ks4omaUK5nZ
BoLuIqvjCaeKoIl7buRtybtFg+vAEgqkduWx1wDcctayyfRWbohN8O/6VXXjhgy3
CbufLecUuH4fyJyUk5lgssMX00c4P0BNB0q8Ogmp3haLI2IW4q4hJlV3ufpQ7KWv
2cUzk0Il5irKKq1YfuhLnuskeNANHFFx+tqnIxFjozh8cg8N9rWIXFIFfLIEyrPj
QU4s5CpI81VG9fKkb4P0C/Pi6JwTnv31aer6n4pZKfB1tu+InZd+od9br2bCyz/w
jSh2+5+twP+F4V3Lk4krIXqQ+Rv867URGS5ViQxd7hf+VE+PCpHdOL2Jh38lxVLp
S047qo6mWCEvbt4e3fJqscAvCT7qjukzPXBjsc0vFxksXO9oIxq9dNM38+qxaG1D
cVfOEMBNCYw/v7HZFtqprSWOjIfrJ2pkMcdIj2IYMvTGbNrm5GXi0nwSSeMoNYIl
Vtic5TfUdBHvhcrLkICIP2KAh3v3aJTsY+bhL6O1s0lS1ECFngirejXnU2PbJgtT
n2oCPa1clyX0vKlafyDnqbRvxSswHJnnyTLMOSwK6Rym7Uv6Qhd4enAS7yI2ecLg
LwEH4ZXeL4d33gIXbHBnaOdnn3ZKbU1A9DPMxhsrgF6e+g11ulLxe5uWEiWGkzUd
FaftaTsA03KbOheHLw68ZQ5mjoR8cx0NNmymLUVNWkDXMVmtzFveGyUqIUuoYm8Q
fVStNUIWVapjuhNJcsB+gO37Th9hTFZ8LbXIwdJUlVMSKANvUjPJrGrYhXDxiBis
RbRSCKB+3NPL57Y4MoYd2x5sLjUQEcQtFe5s40dNBgB/vOFT0jbjwUqn5NbKKSDJ
tTfaJ/L+EXHALtWFGb3SuQmbYO7H7W5agdGeQTlNo+DX8Ffw8s4dhhIDOdu7VHq6
A5slG/WyocOsISEbYrxWWe9IciLqkon/SUcZVXVlvB0f+cDYKjVziIDdFsiVFKed
K9RURSoERBBj1MGeIPqtJtwnFfJx2LInKCipkZrgNs2YgK+bc9uPJuPtAmjlTuox
S8NrqC5tDjlgXysQUR1bYxZqx7/9jStqgruFPV45o+zoUFaPqGhZTzdz5Iz3jaQP
zo6bdk94PdvVcQGwjYTrjoledc7mR4swo4kKfuwF6Doo5Ez/2CBlroKcTRqPu/TE
gu+i2K4FVyAxIeT8+reOht1PZlVqUBUd6oTS9n9f1/oOb56DPJWb+OLYdL4bZOnL
wRSXz5v9TXsRd5/fRKkFVLgaK3/EpiKwv4U31wtYOfxV5Rm+cdVRtqiLx4nEVKi9
KXkmw40GBEzR7gboN97TPol26m6tOg7J50RXMfLrLQ/MmNKfSwc+8Wriq4Jx82Fc
+OnJBc9bdYbXY97IN6sXDwiCvC9mGfij/RVEMe4VhzMlvFRzdwcgXJgTgPIS9ZPU
q4n7M5LxRWzjE7NO9RgrVag8RaLig6kwnyvcA+tfKoA4t7Q2dNaMdlp2MhtVCWuy
xiu3yWxO/f6VS068GaL1xf5/cWgT0imLut049vN7WKNC40T2pN1uQD/mrmNOR0OS
zKTB/OPPA93fwu/N1zVyTdE3qjeqtG7fJR9t3BFwr8+0qWRo+JE+XoRQsCnfTk5j
YO/eqAjinR83fpweKdSWEm0aVEMVx5hTmQA9CLOXnlrmLEYt5RUUTBzWTiBZDpu3
j0VPIa0xEyPQBFHVU8d2cxFCu6FOBHKgTY9hVedvWbMnx9YmU/hECL+FZxGyiL5c
bbmvAbIfg8d4yy8aLatudqN+ynjC+QXolPKWPt74GtBHsgwHYLimPI2XwOWrvFFG
Ol7+tq/9/SIMOzX+5a3rTdLYBe3KtztGXYWaSJrZ6NkW2PEoNcQNlJR2Na/+pgHB
/DiX96Fbyrf215i/1LxaiBu2bpM7OL8XKe5RvGhaHp3Mcg4HRXCpCt+Xm4El544r
HSguT06W7megFLsSxcV08YSEzxfm4Ilnqy7SMQa0aK/AHkjHd8kv6ZSS0IKmf3Ot
P6Zt5z1F1O3rs8Ujo5bI8GF3/P0lv5AI4roFnIA+EvGcEMJ2T8AjkfEYs7UCVOQR
jbDBEKVpzmr34NCcXlTBDsjfwXG6BVw0JreEIsCPqRhbxuapHBp15NPbhJdg7ghh
viRRvxZ0ReEBGr2Cqn0dnlLu8VxqTOfcZrlXOjA8yKe4plzWcadgcwyMSHS5QVkJ
yClEdbZ2JA3/kx2L98huaFyV4hG0YijYGExrvY4X+LlmILb8tfs7UGVAeLZVA0Gx
vElCwkRgtwV0/h1GPFjNAjqwgmK+w7unFZO1s7NzYqS2mMk0m6NPz6zaoREoI+mv
3GPkJUKGOT4Zi3u4mzjIy3Z4L9/ZBSelgEQsmECYXOnerVm1EF5VixZK8olJOUcp
0YTiGlCPMqM4Y9xfFJyg39gGNMOcy8Xc4JMHuvMykbrMdv2GdEdoLP5fqtH3Sn6X
CufEzRii1u1/VT4Iyou+wMn6GOOmCm0PwCCTrArSMBP9AZ2MNbza8qRK2kFjy5vL
L8XMp/0aUdSRlnUzQvUFxy3G44WK3YfUlUg7PLWK80hdbzlTZngmc4ly8TXw5Ahe
GAW4HgmIjDxV9n6nXg3MS2P0gBe1btCDxa0UuSYdfjVcNT9WcPbA0GxbmIwzuG/G
HD1j8ozu6pvm3g27Xv3yU3qr4S1VVTtF4btyM8ZjDoHf2GL/0rmy14oJg6JzdqMw
jvhm6cQCxTNllIrNGilCngQvjAOpeIBoGI5Uuh6dgxPZUO2Vmnvd+6XZ9/Mj6cPh
yev2t6Uy9d4s7Op2KpJ07AESTodMSZELkh16ZTiU/aQde+0HVby9r/ifRlEiBAul
HXpSHe9mTJsxr6T6ePgpDA==
`protect END_PROTECTED
