library verilog;
use verilog.vl_types.all;
entity beh_vlog_muxf7_V7_2 is
    port(
        O               : out    vl_logic;
        I0              : in     vl_logic;
        I1              : in     vl_logic;
        S               : in     vl_logic
    );
end beh_vlog_muxf7_V7_2;
