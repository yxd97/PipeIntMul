`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lF9TzZeWeczwUTbTkcOVpBR5cm6KaIDUg1/BbS6k4cd85vvcbzPQThvNWh8moYWG
6gkoXvCo57wYYc1QuzD8ThhSYZMR/BuzGMxT//4YyPO/qBm6b5KT1QEoLCoWdKYc
kmVRALzWHD0MkPbmacnvReHbZ87zfcHaGBkUp6CtcUJmcMMzgbtxfheJ31/8WLDV
Hc10cvLdBXdC/zZD+toIFTR2qSl5s/1LM5q0zuJI+pC8jQbFBPzHCQDMy+RBW+Zz
xFHXLUlFPtYUiA6cWFOulBew45dd7+kUhklR5o01gdqpBCj5gLaES9nBUgO1hIJA
N0G+WzzOGFkwza9LoRUtqGhUDGgWnyYlr5QR4oMVgCCrIXo57OpD+qBSb/XdgrHQ
E+PvqWK1g7/4l3UafYVhXmMKjIpTeQp78ISbNbWGervTU5SZBpJD7hlmZHJU1PBF
0emNBVpsNpHIVCWprf7LOlVAB8+zd537RcXCgkXo3S35/uE3rrdk6cDwx8uW8MNZ
jK3UWYyI9F2/KTlYlML81nmclAQCec6plaH5iRt1mYVFkWAmw+Ns1Vn0RLP0EH6K
ZppD6ADNjtaAG1HzPAbVM4DytQHDRRmVKHnGq4I0jXvnFO2VWzBlkMwkdK7l69j2
LVCMsdfXkce1Qpctrlrdc9PmNiMTrbeBAYyVdr3y9HBOqwzqpfATUUSjitk6u74J
`protect END_PROTECTED
