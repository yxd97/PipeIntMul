`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4qpAPeCtaoFeLQRKMWyApyfJNhnieruxtUTGpzvo3WZzNl1MGUaRLEG/c4Sxr33
KSFjd4sepvVD3hKH3CWj0kcLxGilp6LmHocCKmYqW7YccjqezudCjKQvMb4u/CFh
Iu8rzOWzTuWubNvx6SPArkqgPZ/AUxc4WJnZTJkfb7T8cM7DsoqzcLVVGDMqeMXj
u+cGT3bTUyvFKkQ57ajBeB+eLINtmnAOrK0Us0cTO/7i0xs3pdK5o0VihaugEpV9
K+Ojo3yiIZ8XQ3saVV5vyV7H9bh7hbswdyHgSP/JvCWNzIwKnh2GwC2JDX5E1tzw
kIuEgBTFPNFzypCFYV8++RWsFR/8q16caUwz+movEM5vBz3cknq1shY07Smp6Fj7
GKuwEXo5+bO29PwFM3fLTDfA88vreZMcgi7KEsZJnm32dhLicD6Hp/DZJLoSisyl
FJX1zZzMTrTgjmCbWLXxuQcMvq+XCYpKOlM6x88nzfAO9U2/sCIIMUdCs7/iDxTQ
NIC3b0owO40sGyKgs4Kqm14GUbsfvpvN7sHip5gfU7ulP4o0ng7L4JBrbZ7G1JhX
`protect END_PROTECTED
