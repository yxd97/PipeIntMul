`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EEqXN2VOnsk01E4OSpRd2BrIMwgQMkJwuAd8rPmyGHg6hWqnyuIh3JM3figyqV9h
0qebnx3KYFANE0fZR4yiLsrIZb+oVEFTAAfObJpW2WivpWjiED6ywxACt68LANBs
FHSLPFyxGvT4RvejETwWMUR7+GFlRaaSqKl3+9q9d8d6kxX2w42qMGl4MCF6qE7A
3xIrTc6tWRB53jdx6EgzhBHdEGvRD+DS30HhsCUflACFYBZiQDdMnGa6RnWbKLhz
93cwixler3nRBXMj35fPb02Qymei0KJDRbfLN7vReQaQRgmolacx+s661zB74trS
OF6z7e5jz2UZ/tePd9lY87N4dIH1dt7ajC7ihbwLcvEryyov11qJ6vs4U+CSwWs4
yDdZzMCCIcrGJosJyWSvYTHhgQ+Tc+FpyZs6/6W9yAqj+Z207Yr4GGloic93fzUj
0W/PYkU9FGK8DptaFKhRfGBrS4gBswkYsHA5MFqrmJhB8b2KZHSlIgKWZexigtcj
lYB78Q0Knppu5+Y7DZQe6ePlPjNxVtz8DMUenKFTXnq915ugDhScvBFmaDDE2ztv
3PdKSXlMTIND9WM3tE5+DovQh3VnuKx3YValbNA1B/DUBXylTBsOR1afBDVHc/0k
Hw9c6B+qZilXnXvyQxQ2u6QUD51kWH0bRevclpxljial4ldK+jyGeHoa2QKz2rJh
t3X4lE4UovRZFelj5wr4AprJidnej0XEiKLq+CgHhJa0Ev8jP4ETHUFRQygD03Qo
90N63G9nD/J7m/ZZjwKEXZJ2wRu+bPq2cEu35RISUvsqSPgaJsffAxYLD78r3BkT
wbvUls7YGvndcRZlxtXeWX5X8RXT0efoVhN5XnYDC7ufjwpHS91XC6T2Ievwctz6
`protect END_PROTECTED
