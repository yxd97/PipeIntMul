`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3c4ta45AjUTkSIyaMVGBQZpsXrB/CCCSN1MSTAjOcm4/UFpMa0a7Fum6uwMrMCki
ucB8I2CDXocM1WXdamcsw/qOua/BYXyBe2TRbxEW8MMlxxHKqXz7jnpurjN2+bKK
oio6P6oX12fQkeXWar4LYn9Aimpg13MwkWfozyLXmshSQBEBYwbRqVx/bvua+IAd
i+kq98LLYZN7upWomsrZ49uPybsPy430M7YdRRkvdr+gh/RRcbaPd0DQYCUNrn6P
3C8geLUMsFZNEqsT0gYUH/OAtZgP47oLbiL2IpF1vwZgnLO1Jl9v7rOxfPfI99Af
q5I68ThdkCX2PxzATf+MWMsMXuX7+BXYnDtioguFyveGNcHL5FQPOUz2g/ySpiXb
5T4sVrvdbj6+WavStjUzVpf1ZBn+L/3iw/4WxQbqiS9YdnACj5KBwwXrma0PAlQu
jmTK5Dg9VlZ9KYf68qbWCFjUKY5lfkoeWBJrXRMalZk=
`protect END_PROTECTED
