`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tnQcKqY6JPA4CtO1EI8/uN390Psvg3XO2B1F1bB5UxX7tW6XQ+4Bqcng6avu3/fq
us1qy5oD0xaCd7hL/lmcqV1LzviHmivj73Xdaf+E6yljmOxX/gnH/+WjNxVbFhoB
9QaKQgsdbDnbPmBs5QAEMw6s4VbwsSKVuIHV+PqbQYjhD3SZ2Uy5aRTeP3bAFHn5
GqtEP/PKVSR2QLgFLbwiB3uY5bc7EOm8xaAzi1QpiQH51EgSnUQZuoJYVxyAN2HR
yGdeUOuCkooR+NL3tNm9c8X36QoduTbR16t6KaPkfFzw5SMXrMRNBlIeoCMiTlXw
FJlJ1+LeSEzou0bU9JyXMNSHneypYiflnlagGD5+uoKGP7u3bQrR64sS3OJxUQZw
xERfOwylgHGG4ZDx2JaHqg==
`protect END_PROTECTED
