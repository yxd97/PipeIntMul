`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5CmkY1BzEj+fByASW110zvTNY9Y7M7FAfBt8EWMVgjCGGVZOSDm5iTLV4ciaTPvC
GZKZJfqe7LrIlDhB7CxBgJxWaEee/NLS+rLE4edQPjkDgeuoQsUvKjYzhZaPIBUQ
rkCTeF6JiXRrUeG5dCVJBC33KR72suGpCg8e2WX3Rjc6m0vLiPhq/R+RXFGaOMpP
PhoYIHuoytuw4KRp9frlPg2MZsHZ00Fg3AUjQgD0+mbD2d1ZlHQa2BbDZEr25EkC
jG1nDkpf0xxtPWj2mP5hVWhLVx8+oeGHsEHa8hlbQsRmPfMMlAND9+b8potsBEj0
Q7qr5PMg6fZ73BLcTciWtqN3kvhJWaN1EXvktC3Xe5srLN0nwXswMrU5r3fxE33R
`protect END_PROTECTED
