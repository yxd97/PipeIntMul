`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/skKABmxt+KRsXtz62i27TTJkMm2uxzKy45XC/L4pGoscV5TGdzYkWA6FE8y7yX
RKpHPG341zZwyIqwz3xsQ8Dt0o9zwLLPfHT8UVh/cqbAOaTcsGxJiolgHLoQvJrX
6lgM+EGVZg8lRmoV7mZ95isvTAR6I32WcY+E8AuM8J5+eTZurJW0P7ubJ4A8xRgs
3f6L+w657vcOfVQoslJR2aEfSjlLJvbl+cVPAcawGtY/W89VFf85mUsM5Jwg7t36
IxPUmh3yltjuCQK3jWAjhQ==
`protect END_PROTECTED
