`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QLqAzkb1M0HEidQFovoU6fuivZRR7rXeZC1fHs/mtmaViRyzfO65eKwUDiGU4m9
QbbzspyJ2POJpKMJv8eUtZJ9hodNcQCFSC6TTkTp4J64LZ5vKpxz/aCVWmsXAPtK
TbOVyfVqY7k3UuILnzpaGiqUWRdv+Bq3SU6W3ParB9AE5lI0TUbodPmyAU2IEZ8u
wOMa+7blek2I0wIdLu6Q53aBjKM56NedB3Q6tTNNte8xw/8Qh+Gd3hQHXk6M5Jmn
+RdsxmPWxG7ovcflc49fu5eexyLnIWbVrnG4+U6JYaYsKuxhkNSx4NfO36sSt0RM
wCn1ETFfrMnKEpDjBkqZ/s235qTLYKfi5tV+eeO9RsW7vNlxeDPdXd5sM9g9Wnlt
bgpB6O1q+Z2E87EhS+mZHBjI2s37N6YdAXuUwQQb0bUBIZ3PlfJVg0eQA/O0N1ND
Qp491j7fUjUa/RUg98lb72Qex/iKHhVaDp0KiTPzRXEK6ye7/HhLGDEdtGOTCtg/
zHUjACkmQ3XHDuQqiZ7G4PAGab0tEsEor4GG3p5r3VLoNZkgKVOE5XZn49vX5sFX
a998lX4M7meL48pe5OrtlAwB3Vwxhy/Jl26arRL0B9Otl6kyWH++x8EtieQvi6Ks
xEYM1WkMZ14XkLcdPWRRkLoG/wKOf1/TcZ98OmAyc6q8htJvX2SVIjRyFP20W6xB
4d/FXlEWlpZJVj9dIEh4gR6h0xm9oWji3ZXl2WnWF+21ee7hBb/mMfy5Zq6IZy6R
rhPBeAAU+1Dpkqxj6P898qi/feIUyXELkTRabwdMMEFLXFW+7fCb69VYQL8nn4eI
uHnjUASAO0M47+E8H9tqVNwQ9LVkr+1t0mxzq0mrd5reiXN9CNloje6C2mwNhJai
oB3yFC96T1mVpB2YQugPpZCOKwSfSbxrCatdQ9Qv33nr1a21f3B13elxZ7qUjFTO
wp47/+tLMUmJpFu+rBGd+ynwh0NlOt6thGlUKFHXshYFyuqV9GQEk8R4JxDsbItt
BO8WE82teB8p5mvw3g+JIVTqJSPghb2nLP70w/wxLRzR5UtRQszgLO/enTRBhGDt
jGCf1nQ8hfcDuCNfqZoRQw==
`protect END_PROTECTED
