`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OyMQVzNPsaGm2wGVqs7TZzY0Ds/aP9X+RZJqX9NyKbf3UxXZpwFLQ/TAZDFy06et
fnnTkATL0CdyVKqunun8MGrh/xytomDcAqK8hAWucgSc46h65bfGfdMFKSLDxDN+
pExaPHu91AGmkvV9DdbmFuMC0sr5BQgcocpQUt+Mdbmf9mY3q7O05Ejx/BFkg4x1
GOgM/L1/0Kft1HgTgfLoQLBma8w2a/WdVYykiYWvLK3LQK0iDyH1/8mRZqtDiDjY
dBtP0EobgF2VXGNfBYOJKc8zIYrTPPsP3sy8h+kTc96ehGyJM/F1LTv4b4zjx+Ne
LmnK/d9YaYD+LXuvtbuUk04lPcKsGqzZT+3bCXTfGFQgM5JpnY4qv+cbC3XF4Qms
4lrqG9TjeWkDAEmjRkgOviTk80THwCEmh4/syK3DW9jMQULBVhseJe0Fli82zjob
7L/ondFZ/GnMPbe9BVNz15AYOGe7XWFRwWNENqFp3e4=
`protect END_PROTECTED
