`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IYc5aAxNL/ZNn5qEPHQS+J142kyBki1Cat66a8MwwDFB48aDNwFY060BLaxLlJku
IUHjBZc9qKPBMnWqsthUznpCs0Uq85AWHG1z3SRY5yyIGX5bW8zDudRf3Y33mKs9
pYDWrunJTNkucyP+T2Mgm7lP7QUg9EDYlkc+CXzuFui0Ta9hiciLf2nJl22nVpq2
LdN3yWy1tV1APGe/fgxhHXNUpQSieb/tjJvFWaCGxN5/p7V76317ES3ly6GLhiVF
X7BZsMEkBxkANAZUBVXrEnVBxFHwvcvkFutlRqWpubZFnXNpOCptUlaj/rhdxDuw
0FWYvYXYH3/mnuFVApbY2LxC8C3bje0wRUD8qqrtBtvLJW59vFrMXM4AWH2VLMWo
Kvm+OyQ6ulXz8nitbucOIj+S3c+oxHZJshk4QXsjaXwcXHDkeUVSMdNm/aOaiHpn
vSsN8rJhM5S/TjAuBhopa4i8EnA0to8hqtljgBp4ENhHb/II34Djnt2HRYswUyII
C7jXLVq5lsUHsA456/lTHtKjo6k2eTCehtNeoaK7eSP6mtlUCRvlv9au8Pf0hgwp
Dj40JMAhpFAQY7EcI1zaDx1+fjQ94h1VUWQ56h+JS4Qt/c8x+Twccc/btw82sM2A
x3WFR8KWDQ5LxFqwI29Yz8dcWmfuJS0GbaWoYTEATLIYbKuD+5nRAPdh+SIKRRUO
RQegOW144dv18RMYEAOkOXwO9DIqZC3rEfC8OKOv5CUV3gYlNvFm60Y1h5HqfpS+
UuIH3dLXdIj0Xt/hHDq6aEd6BNlWjf0qB3BT5GFokJ3u98YbFCoyaA+VRRMGz6mT
l41qe4MUg4uD0lwkQ7yLwFBJcjPti/Eu61aKq+Qg6xfouD4A5mGoaAAzXuYnsss8
wq/jmI/HJ2Whtrh+rmBMIatnYXdo4lUP4AxKYg0aOgWYkgTG/ErxdMqqBEelfoNm
74h57/dzBn7jZwoLCODUn0S5i5in5UDr93n0Wmp9x8kmlqkVaMp/Ruq1Bv/XuYjx
0zlEiC2Cpy0T5WTzxehqRMqlFuuBAKXpWtcJt+2kYfx3/+2GJPbbt6bnTJatEs46
THfdm4RInBJVZeYqQCfElw==
`protect END_PROTECTED
