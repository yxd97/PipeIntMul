`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QpNKtmE3k/M4hPhK7t/lDWXfrcopzYuNx8sPNCw/mXKVdCfN/0KCPbuatG8C5vFR
MXok/l/kLjeeoi3i2t+CQFCxTePr+Ma0KZMViAE5rPv6aMsZEwuDwSoigODSasNi
ir51+rab2TN3cTtR9ZAyN6Db0EnrWCgbi8fwJbc2tMksJ8+iW8ilv/2wpw8LtfJP
KejOYxFVMIcyP15QsXwKspCHMJ2rRNzUA2S3gkQA/RnvhL6/rVTKM5ZqWvIA8v1E
+rkCKQQp4xMPjN/1E/wNDvAP53qo2enfJ3txQh08ta0tLuXVH9ST3YtQqqGxL8Ok
2DvuWLiAth74ReFyY7xqXegGjJU4e8kxdBp8DhF7qr4ivFxU8Dwrnmli12SKVOsC
8nloT9Y0dovWiWyAc7Cv2CqA92t5ydkHnyHO4sNLbw5xZ1a7ApFwEUNbhidUav8g
vJmx+sFMWKUk7FVOoAYeeALbcecj2Q9Alr1MOZBxMsq9RGPogcp7bSVfC2boR7uZ
PZGG1Je8sMWzBhfpWXYdp+XM2Z5T0YgRJ1O9oRlzAMgNbjdYELxDTgnoemYxCuXu
LtzZRzufMHaNT43PjglAeojP0oj3GXnXCeWO9EahS8hmqtb+61zltFy2A6P6tVAy
6lzXht7G8jL+acstRblW7/WmyVYDOHhknyWsFy7K2kM6X9lm7tnTULLI/6NO6b+p
2EYenaEgspYMWoWTB4PD4rDnwW6XKpRvlzoYixpxS96V+tSGqXbe7qaEMiCOnGqb
W4KPthU0FfoQnqkwt3wNrblgCHWsbRFgsCKSOCjCAeZQT+MmJjbIePsKWfQYxFDs
yJKUOtCpcHi6vrhVikCxUjBbS1dPD2hM9deiqO0KNrojv2CzazhyhXt2+GRlOpUz
ZKZiVCrsHb1/cnu+V7hmZVSmkMtyd0f4uYJAPk9R2DGPf09UpkpHhwQsMQaYGQ02
QwhtngKQu6deczbwlvapZUydWy42tt4AxQ3fkAirvG0nTLkrcp42FffA1nZvBOhV
htplryiXCwTdPue0MSxpVXfRbL3Nxe5uHqnOzaYN6kmc9Q3ib7/7FS11MQhmN+iN
T0cQwcmXI/qkzHK1RmehrDoXIRjxIAfPU9/W/3iiqNN+KfrLoRbqXDqyb/9vb8ed
klxzXaEZ2o7YNHDUML8xPcwjeya4G2z0sa9UmkKwQxfK7qty9RrpSTQDHq8m7KZn
LOCubIyfyZzGYJi7cLAMMikXzBmpcDuTbk1SNK89HZbJ9dtu6YTcHLQqe61tDwjc
j4RpaHfhbyjsAlRDJMAfqbqupA0qfC1Kb4i6ZIsQa/QKrUtKDYT/mK+Uw+E+iMCG
EcLpnllwcf1QKg/e7q2oQWPNeTASr5igZ31UrCbkaRdmS25JAyJcHKxIrizNlkq6
e8p9tE5j0eA1Kmye27Y8fES6BelilK2nXdJMg3rAeQodwhFmQtwvUO6MUJFBATVI
D+wBon28pABPxYGaqs6k1pWH+T6kXI8cfdSP7P6QcprAswO6SuoSA/G2hPBXWGNn
beqvRfKYch/ARh5MOnxJBQ==
`protect END_PROTECTED
