`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuVk/4O4kTs/oeHsdSjRuac25fHQ5jdChFUpZTy6zyZId4qG22PseTqRV15NoODm
vtAY2yOuYkzfXDem6dl1/SwheUOnxbWEzjE6eAd5eoYpM15sKKDA+pQ20zXh0eb+
B+kVB61sdc61dET99YdC27kZnAqyUOC4B8ihcbrZSWyRuGatp97czSgGff0lcHOl
8oRXejmRS/p0qSdJbwaj2beMHqN5bZmrAgl253V7kso6cYYlBxpBnbJIgWm8Ekac
C1DwtOducZlFF1jusiE3ofwlp+Q8NS9TNX/B7cIggvz9IKHlwjMAWd51yq/fO2wV
Ulzx7WOwbwEHvHf4lvDLV+61AnVBU9flpQ2fCB7r/l7VWeJSaNJD9uaphYSHKmC0
XygOBG2HjCiex47tOL9fKsE146LRN/MOTTP2iu2Ytczz/gC+pPZlY4MRy6m3tdFh
xRbkCjrkUdfAirasK2hplg1IvxCwvY9ygJ6f2YJryOORQFww7Nbnu52OA1wCFv/T
DNtIo9RJFngFPgjJumSZ9ly2q7fF5UmK5Puw+tEIT4nliwX9Jx/fauNC1iOP+wNk
bWLiFr27z89nYbgUC/iKbAZ52bfciI41hLcYPLHJ3X+JgPrviV8pRvm0HToDjNCF
J+XSrHQafBJ+c7Llo7nVj4bvAspod+1IryY2XoNhgPzDW8vdfthxHfet6H++xVih
juM1/VgBI6zOtNgn19hBKQeVkoyXwkUSTaB2zt9AZ+BJx3Q5iH8P+caXbpiE9diu
1yd5vZCnP9mvy5dBVPUdIVxW7jDjctCr2C5Jvti+EvYkmVxqNLNqrJ1F+IH5ov4B
YKd4V9imdbnNBReauvLyUapcM/3EypwKpgb0+TSJSUszHtG0U8ZUDJy3bjcADkdv
yEf6o1Azingjl9rTF/wUfjP/h4DVsgta5fiK86l7Y4sKgts3u0W9unTaOg/ilBLI
AeM1LjzhonPsRMDtKveAVd/9a0g4orn5u2Fu5yGQ/1p18xDKvA3HAuwTRKOHz7RU
1U5DRGDeC56A5/UBNML7ZqBmMM7TkwTITkCBXRWGJopPAD9YiRUsk63ORxJSZYEv
/t1PNZlARcG/aE7kZuQyH1B/V9sJZnaLre41imEzl4NCID/ohfhTnPVYq6KxM7Nm
RHGCG8lkqmLm79dO6MFmD8MXlAgb1UtjhM7efQkVFg8DlW4NLjLr8r023gdiBGsz
jO452zvsFfH0fy/6B8YY7XJovZKKuKL0fS6pLVjNkgcJXO9Uh0OUayNoK5jglwcP
yRcuZ9l5NdW+wYSIxinjLW0vjdUFnGYqwE3fAABXRYhmhakVig7WEk53PHsAP/Sy
KhuVoO7O9hEmaA5TiZXIv1UWarRhj/pUTV6iG4xUOOppsoGh9KlvcdjO6RucWffR
Y19yXJQ2X+BI4UfKrdzhkqZExyngod0xLcx71T9dGO5sMKwLfrErxOfQxt1sr55g
rt2Mr0GqUUmgFlLXN212KLFWibnLb5ipWkgrxuL/B8XCzbpZjP/jy10UAJ0XQdJA
2KV2ipnrRS8KezygO+n9kpPMED8Dxm1+HpVXCq/qP/oDL3c1mDoLshcd74Vj81Qp
R9zK/jQoJTs8p9ugnAAfjXRPObA2pNWgiK3hhLdVq47qbyzL4lTloxGkPpoU9gww
YzbxuTRVfpN3DsbjcZfpfH/px8gSEgJxWiFWL5yjMYIWdYkFc4yswNQ6+Lmav4ig
dfCg54iaq+X3aiovVjLwpa/qh7GN8hbEGfhMLKv80NEbtehXnm6/WiWwLzA6VFwu
8BxOLFj5C/69kvO47f49gn192Nkqi5O7UeXyJdr4WWn7xmBXs30yZ0OqRloiaGjq
IXNIM0y46q0ETCu7SlhQZUGQFAivQRoivAynfavYLHINE2IWca9dgROFDolcWZPf
`protect END_PROTECTED
