`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQdigW+zYVXuJPYAzDMm57MDhZzbSZ+cjgqEkuD/adGUzARR+s3njYq7SnlKuIRm
95G9lfkODLDw+wPmmlhRKQl+6o7MiVn8Q7vJW6ANZB6XyMKu1Ik7h4dGuEtwQrRU
lzQK8W/wA6d/3S65VdB5P0O08+f5PuuozxXn7dXY4IoTkARWFF4U0dMuoVyeYr7S
WUVgpgk7dYAKN3UmIiLMdXWcLEsqnId5YB44+Bhmeu7gRsFamgqlkFPnGpqysJbm
g/wdwbaeXQ2xpHSJ+oYsXdt/osJG5V0wcuI/uBtfsWIX8ijlgwOx8GZ22zoIJ6CQ
rAm8KSZwj53WJybdOe8GUVtdljyHi1O75pr4Zwa72+XnHp+IUyHaJO0muBWwl2N/
KJlI919BRSWyxXTPKxxqH1QAgQi3OXa9rxKKY5ia1PVyvRExVo003aCokfNEAQbP
h1B/5ZLuQho7R8kzaEKnSHVWKroGM1qSxxp8wj6yYBrp2t14YSc0HCqDzDdLacfg
0oOn9LdIQVGNuHcTRi2ESenvtto9izETqy7e+yFYK1+rZkAUiRBLXoLPJ+73uarr
krxXHPX0/DkueygRDIUkAugWp3dGM/rMPLHB0d1waNombJ2uTJ2CUV/IbcZct4JR
TgugOSHtj199UmIzQCDahXZs2m23IPsv8WaT0x47e6w69fEjrSPNBjPBuPeSn+xs
5DWdv4MEAQrpzDjHvf0mKoXMIiNTJPQcAyme5O+3REmgkXuGQ1x2Lpg1HBd2l5/u
SvitVKJZ+IC4trwddhOPgpJOEP3yJx24YV6cAmguFCCjt5RLe0GU8Ci6S+zyO88w
x7/SnLbkoQmfgfucrqEL24BWC20wClQaPSh7vNfnh4wv/qYVC6JZqc2iJ9UvHfHS
+ItN+siFobyQIHlVX9ZFpGOqO59dfhvvu9YvHd1KtAs1/0u8D0neDmRuijD0nOgk
1hvMjQVZcRvL8TpJeS0YiAnKWy0PdvbTsjjSYWr0ZKWAqlio5vPZnI8EBIFuAe/M
QEPULYp2l2ZtRKA8rBQK4emLjvaRYhPZ82i6ya4qqKnXf9SwpM+bG1rJpxyFvZ5L
5fAIL83vBJNQrEne0gU0CKloGN7kRhePFMnnaEOVaWDRRGUB8gGQLidLkjFxzZ5t
M1vkIzohFLugKE4FwySOm+KL1A9ba400E69KqrJESknnbUVxVbnln1AKeKVZ9YvK
QCTTKEPjQV+ghtG7GZfT9WeaMsKQYPjZ+t26fkO+tBw3pBzriKZ8oAq9shodMebT
2zk8rQjeEXiti9QbNWy0T7uO7D9EGdd2uduIn6CjWEghaPYV0wUGhgDBLFf9L1gs
S1v5XvIQ6NAODemmMJmk+s6LplMOB7QzClD10RCk5OepJdgdKH+MmRahYkvecj4F
xiME5cv+zdCqFOjcAJB9VYmqERCVO1lY08VX+sl4bHKAinRe2dmtv7dMN3Xk04kz
8oAm9j5NcBIFNFDdO5fiaB4JVK5qxHcZMtDyal5YPCv+PHAX2sB7w4YcSNFQvuKW
PgoArlSwM9R2m12cNWeVoI/pG51r5emK4hQ11OL/UNXuRjSIuCtRAHlK2nvW++Yn
PGA02wBO8govYvTMwsCoUIOxbLP8LTZbwsjyPlUUxbk4UXYSf3VwhfFiTPTo/KX0
YEV8FaGVOlj8Lm1guC3n+tF1gho2wXsmzdpYkEe9zBYeCkGaTMquMN3OGy9ZHonh
kHNL95xa32BTMVSDpfiCY/tJR4jDVPlmfjvvshvj7ED7imzKTDN0WIaMkeoOvkKh
Sf7rPfbXuufdgr6KMD5KnzkBXI30i5AlJibV/Rc5jgrbsh08uaN9sSZUB4GaRqI0
cDNyfgpXejP6xQB8OKPMV9UZziGuTyc0WjvPb1bIwvpfKmgUjca/9FGrHxAQQbr6
ybAEY12aT/SMNqMlJlIqknpesujZCkD69Hx+b+Y5UDu8XZGF+DQoG6GhSPimkZut
QK3I6Rmuc9ckD6d50px9Z43Uw4wNY9lJbGBoJMgCfHwN4LMw3Cg2TgC+34PMuuIp
pOjswJa19y90RBlh5mh8JaZqdYNmmSG7KDvZ17wU6fDUFSdZcs/4J47/gpyr/B0C
0fGofFkK2Uck3RhtIAilHZVxO/7+swE9C2icicTEQs/AdqxmagS5Gl6QgpuOI4bd
SrXXQwHpY/ttrrl2+G+LNuSCGZXlVwK8cfwlZirDSEkGZGFbOakS5x2LGPPwl5Tt
kkt4RAOMQMqZpkGglUxV5kpr8HrmZKKDUzALUGAtcDaIGVvGSq0xJzO9kFqF/nvc
kDzEBO1ueIpejlfGW4JTlmm0oVFb0Yo472GcLm8amKypU6EBNSY+UGsFMPnsuHd4
qdnok4EdHvD4wzWnYu/pPn+pzAKLeACxgDaM6yF1NRMpGNO58Z/+7gk0kXRD4K8W
pLS1TuPzaJ6K3bHSl3PgJjPiIx52WZ2ZusW3NW+R6rPGN436DdA94/IPCkmqZeAr
P/QUr4Vu5JguzRHtwSgjMSVwkZ74MceHgpCEE9iNhHv6MPS5dMDA5cB6L7V/kk+3
2LEl5u3wV3R6D/a2xoSXi+mrC8/QGUxSZEqHvowncfZe2wfXtK+4rNEXQn/yQaqh
1896Wx5PS0wyudqSeH2mHZdEiUr4OwI6k2Ivxf3rhLHNRh1/tcwFWMGg52Yp4NFd
urS5gNCpr7a+IpLLScJ7hwIRWZiiJ4yvAVDZrPqKMX+Y5sHHYhAYDIJRXu+miWu+
b1UKW15hlXxbM/QBI/mPezhQdr/h8QQJ+1un6HOavXZ1+UBOb8LUQ3siw28D3OEl
GVOJYaSargQX/ewfy9yj3alSevKPg/myIz14ZmRtcnswyeVc+rI6yqHPohYvpmeH
HkLtH1nYYFAn5aQWeQ6U5HcxM3acHjF0qZvCZVl3tUNSNKtKPGXw2wUq8/3sHjDC
eEkT1GAIJec8+PtXqXPs4WppHcLmkKoaxIGnXtlyluKOPN31H83Q68mRHuGABsNR
f+Z1dFXrZdj5ntNS+UZCaWoIT4xoZIID0Cm/6pPvb8MXHUFF2eA4ytYtZoHzFZLY
dceAhHSlcJV2T1CKMppchn36LcW9ydtnmIh/cIr2vqBPaiVDL2taZg/9VDPwju4C
BfG0VJ8/g2ivPYDYNVCunFZm5YFEqCnXCA3gsZXCarl6Ee7yw5zqj4FeRA21vDgi
`protect END_PROTECTED
