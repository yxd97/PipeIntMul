`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IbLzPKsARHA1X4x0LEGTE1Gm3BQMwTgpdWKS6yEf73zhHURYXk5TYt3THXX0Sztb
Ig1WCODTzhC4TjTTctRHsvjkIyilyRcdYJeTbqjgrwURR9Hr7tX2CKO6rAkx0zvd
naAk0rx5YreMRdVQUHvNPw8ExVhi8ha/A/fWYSMcsLsmYXz47TcpfZuy9h9dGNqt
qHWKdifpJv8NX63NWyfgk7rWyjn2UfUD0E7q/s6KMU6JYInbYWZp8Guh9yGyUiQC
PeaOSCO9jKq83Xzk1lMs3jD9RR+rNAnn7HiShhJEp6VFrkgRapV1zaLcWpkHkkmF
uD5zoHMeJXMJSvS3u82iUw==
`protect END_PROTECTED
