`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/aXD3Pwm8qH8eFls89hjjHgF3HVOi8DePSQs3xQCQrz6esW0dmE7cQ+PB7dOL1p
rLPrYPWCOLOLAUJWOPXGNo/Ye8ncIiCQJKLHd4w6GU2IwuIrikO9o8h0K2WysnO0
WuLGk0qgxWWN/60oUuZtq/EQAM8lurVVe60bDq8z+g9NyznJ37Mve2SHqyY3aZK/
RWuYpYPbwBTy/nkeAEL2RD3fPyL+v39vNpjuFq33sjh4AxjZgi3SwPiqfRPhRuob
gdMh4KXahpjKVppb9s/WczkANAfGR6c+t2ALgXXQXmK/yvkNo43Lh0a0Rtm3GN0x
eXS3tPKkjFBLB5Vu9rUzjNrFNy9n6GsRkVchVf6iPV6t4k7IBPse/vUqQyUgRMB5
9LuDDFaY91PJzwHOGNTLyXKgGi6OivG5aXjnuStDQ5c=
`protect END_PROTECTED
