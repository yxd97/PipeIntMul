`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Si+aGrjNCqi1PZw98JF95rjBmENJFPy4XdR7YPuoZhNi0JUfTkPLKofeN8GRFQGT
XR/vitK7dJlBkIDDGuUE87ONP4n+ZlAH+mxhBqWHtSEA0IPOIsXzo8grkzKkBgbk
P4rzl1+EWKW28Rhv46A0y0QhDnaMtyhS09Bsq9vt43aDakNgNaRoH59gcf9nTVYw
FAWrOwr6cCRJrKF1Ry9tgu0UcI36gKbX+o4jTqjXqdQPv/xR0WY1aVurAuP/Va2U
WSRKdG8g7UBhEk6bGIAzc91X2rrRE3JDzX7nPgZ6rMygJZkXCf3CP1v0V7a9/eZQ
VrRi3z1r18H4MzvtedqPOAzi95q9+wIr6Yqg7S7nNlDuWH8u1ikpr3BmDDsnbQJq
RXlQmxHjSfYFoBi6TMk2dzABgy8T192tV5cG9wo8QKrRdM5TREDd0qHjIDd/V0v1
lV5/TD6zAroc3D/Cj/lrTO0zP5nSlPfzp7QOdjcYuh3CDSfv6MNU3DnJxVuU1Mjp
FwAaMPWTkWlcTJZGzf/YNeG2AltoE7KsQMbn17BCX5dX1sAELOQfVJrcykYsOz/k
N4PSBFYpzHLrI8z/ZEPGhMHfvCzuWyP1JZ6KJASAlALLCpMl3fiwtRY8aelW84wZ
r/z0ZHRHRACpqi/7TbPzCQ7FfsmVehPZUhTxgEbGUdTNk5P8L2O6BoWriIv1n81E
KVMw7FcvhmkjWMww6X4zEwSR/vSB65Gl4IqKR/ozHx3bjt+radKHi8lE08t7/+mW
OS0shfGFQmltsL9M5e1sd0aMHdV+r8Dw/zUoTIN5flfWdGx7mJ5SYPWOWVzCfPex
TffgSo89M9jiKBbvz1gUrg/oyUf4VxIHprUWbIbcefa/b3qDVADAxrZggppNF9pc
+carVmlQft87BQRtMUVhIYbMugS+CxAnvGYHfFpqfcHvuIaWk62y79DnBz0SyFK4
6O6EKw6RXBJxoG6oKchxlqGaZJpiBirRiDNsAw6sVAh75gAYA3Er10cvBff/O+w7
2lPQZ5YDX9nXNNZ9C3iCFCt1DPhZj9WQLk4IuhiOg57AIPhL+OQxW2TTOOqJqAsX
UEbh9ioQ2p3qZ+dsvvngZcc4uEXREXib85IF1Kv3fBtx8l5R473A/A8xNlqAbjPD
bqh6tbRNZlRv9AZVmB0EjpB9agVKQM2Ram8bUEq4F89ozeE3CKZNYkbZE40Gjd5q
7yMeIrW5Q7VaHQmi9vkY8DnR5NhNlRiZDQ4gtUtHZXhiGKUVv78TQr09k/R9XSPb
FDp0LDYEgi/zexMaO7PHUWbknk/M38qXSqxkiRr0HMRDnxkya99UqYtkpq06r7mn
HkaNg4x30okHl4G2V6e1HJ8wfbxmvWL1be1elRimJJsE8UB1N5NzQ0NEIet/7xY0
cQKAp/d8itJMxGXDwvKuSl8tjm61gSMo+ZdJTTxW9R1srLpqMaqqvr6HzACjPDIo
V346Zjuim8etnCJmKJbFwz9livCE5gJozBr83iF4np4=
`protect END_PROTECTED
