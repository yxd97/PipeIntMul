`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pD5sa4ZZK1D2uqCAkMCBOnADuhS2hxhcEgzyKfIa0t6dWO5pQA7Cj4MUljYkGzqb
BgOGqGFVood3P7IBtxTWb5ibbV907r+9Xm0RqAZxLgrizksm2q82Cc8fiqu+w6FS
0UrAzaMXT3xQv7sewp0DqTasXpBOm4LXy+CSFhRS5FaWbR3Av+4b7RoWOrvDu7Hv
K104THCEr+VtizbdS6lsclmDsxvShfJdtZ2EPq7RfC6GQDqVb2wBYhrB5/muktr3
ebDg6Hc7t2jMj5BdVYFtqBEsBnYJricx3bJbxAkeWYEg93jXPYxlSo6KXe8WPPGo
TBVNmTb698eVLPEZNpL59rh90+gVdQwpCMTBMb3Vo9yiXzcok4cV3sghqRa//Kwi
5OJJk6Ezg+ixKU9PeNk5dRQ5gL3w0zbgyolTq6RsX9xszwyCHb0D/cCMPbJCf3Vk
`protect END_PROTECTED
