`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sRD6O7k3V+8y+F6kCSb1qsZt8ocee5JZmCv9lgElbnQT5sISy407cVj0ogXxwnIS
tMNk8R17GNvYh/xHiJRgArfO+Yt8fcv68DUbJ/mG8C3E2am7B8wzahI6imz4FOJB
dYVjzpwLeDLt5MvcS1Qk3CdTaIAHh4GLx4h79r0qkq9c9aSj9ro3V4DwQEuxN7E9
c7kSuHTAcG2k/i7nARTBNIFse9IEpIoA6bHYhEB0TmyDJaGFYd2Lg9hj/Wt0e7kl
9IQKzulF4AHfkBvn2deK/HLIaMS7uKp9fXeioHsdHHQoXE00KDLdis8JoxNYn9FC
DQVeWnqqDxKnLXeFAmCPHQ==
`protect END_PROTECTED
