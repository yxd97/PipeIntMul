`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/UXzSAKLBeniKBee3WHufrKF5cwWOzkkB6P7Id9KnpjIxy56T7YDVmNZvb9MBzv
QUWkBpHGGqi1sDUbWaoOnLSDAY3xSNjxt380fNzGzQ57gdOhp8eYfXHe6K8CKaSF
2TU+rP147d6PiCmfQo3xMPpzTeq1Y852U5cXtRFilE9qerkWphVT0R2jdu/yZzX3
AWsLZhGs17zhCT65ju4R4Vvns7XkX9ejz8cbB9nPixiddUvFORc+gcHgB/cOOOxI
Qu63FiePyx5peKl3UnwCXQd4K/2PVYJ55fw9Ypnsin2kHI+cWbGkK5cwMfgbS//9
rqX60PcTn2lKb0iRyiD0RQwYCpokA4wfDDu+d/bLSQvxK/t4ny7grauU3XCTVxns
XuK+MMSsPJyHsMRGEgwiDSXntaxQljAdtsAFNty1w6C1xanR3G7/HnEl9zfZdzd2
yuEIWQBwQS8uoHZ/PFU8icu8xS7weJ7EF/dQ8cV72LzJtZBWiEY82TIm858ciGKY
d232fyWBAe3mEJ/LQBi6kaahPwLYCcsL1SEXjRopbVEOPK29bOQiGqn84eW9iaP6
wImNbLycDocpnRjSmecSxA==
`protect END_PROTECTED
