`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3WYttGQved1ltZVMRJCCuEnQJzQ6Tbcdz2nyBafzMex1xgrZpOFei6gbOi4wXPo
/SKETA5wH2Jb/yaDMPiRNi6bypHYB0EYo6UimIF7iM5ui11Kx5uCDjLItxMdU557
lRxKU4rWnBv6rOCAlkLWKIZ5jYOSwirm2sH6+fjUzbSdTbLyHV5iAT+7iLwzr7cA
diJxeGLkkaurUYj8r9P9890HtojMU411++CfzZJz1gVbL8T6tIBYLEXRK4Bpa49S
3EaWNecxAuykX4wNqFR9NMi71yR5srwomKVJjLEyz3B7p5YvH26t/H/AcmNLJAc5
znwDmNwpKSuxsUpmmcF38VuDOjWl/B8HeJ0mFYmYT7MXZY2+J8SnHdXaaZWCRmyN
j0U0n7yQc1bKsg1ovR+FfF9MKlmvX7jA0UMAonBRQXx5E0+/wYSyHQKefjZiuiEf
+nviTz+GY2vIsjaq2ejUFnS/5YwxN97f7zWwzcMKgaKMjyiPtgQffLDDXJPM/ckr
8NHGTwGXqc8/EDnuGOlSDtMl+A6figKJcHGzwAML5U2essseAVLjwxxwn9tB7a07
PnpBPq2tq4CoMyYv9EWn05ZDkC7f1Qhwbs7ZRTeZnRfhwixIJy6ceG0VHGY47wPH
ku/2eBhTLHxQFr8M/yB1RY5dG1xfl9T7Ymxv0MH9d89R5wlu9311B7kXuyzMwByZ
g/m6caRLQ3UqLlMT58qslGkC1lJBBnbx7niY0wbgJlhY8+e8noDtM6PZzPuO5baD
zXcbREm6YSm12eJZ+cbuXnL677lJTOQR/P6HYeXOA0P6w//98moZ54wwCqDKuhUu
Ws5jZGdFZ8Sv0HT5TzhWPBsCR1BcvcNNLAA+xJPi0Dg2JkMVBs3QuKuZuJLgfC/q
BoO3pk13tCBtY5MBRP9u0YS+BJThhlrhqkFJXbJDJxQ=
`protect END_PROTECTED
