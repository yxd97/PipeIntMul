`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BU7nanJ6xBfgAJgixyWD+6fukGejJY7Jmb5BaC/0wzTgNRBwxJHhXkZ0NWiA0mjx
OJ81liIVNV728nC3yieYeByVxftghG6rr0I60HC+f6yujWTfd37wwxFUY2x+YgQ+
XbchPRQ/m5f6VKezSqYKfDG0dqUJyal5eSlHGmzc+jUaAEw/ov6zlvkYJYExGw0t
i9RZkuD245zshmDXkmUi5MHvhIZyA+v0SZgKsiQM8zVYDtR6YTRLma+mlPjnadj0
13TTghWkEWK0EyoM5KVkdOqMQ/gfY3hbnKIyBicZZu08jCYvUwxFadPQmraxnwsk
7ddIdNDShrZnspSkGBUDa/Bh3sx/YxuRkXjlyW7OV7J2EP+7QtWByFN0EhnIo+NW
klQQxBKKMvutbjCpcU5FOqc/w5gKcqOxBOy7pgpxOZ4IWrpZs3T6HPcc8JZIHpSY
eKaNBuhqfQSqoIA3w0Le7OM3jPjGVDxWV6WN/eaBfB91Z2AegRCesChePZSClVrb
L1t5krZyKqWGO/LaCxH+mWZ0/bGwx5F6RuPHeEp5xXdodGSJJoNLizmAcvO4UUya
8HBoBSwcXUn3aUBBjvPVgO2zzyUF79JHiDudS3jLJkvVUzEA+bo8kFIbqcPHHaF3
aYOpKb+I5yJY2mYSgNyAfxTOcFNHB2kj9QEMHV9VfizAPeUrZ7995au00UPQOpMV
`protect END_PROTECTED
