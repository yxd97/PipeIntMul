`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bKcViZ33H409CvyAYYE9FxJn8OybkuZZLuVutNl8BWR0M8grspsXiIJeDIpfh0+v
QzzmEQ/LbhbAGUBz7KTZ0qo+TGdmfQs5dXP7CeU/F6ASUYAmuehkw2q3vKGuWRtB
po9wvAaNnYHRWZhRxUleNZD8yz5WvPl6lf7df12Pbl24XIYawNm+avIlkpP3YANi
KTTskkAK3OcgZtpyq+M378XBYfcX73gk2SP+qe38XDUb83ziyGwaBmkqns/KOaHy
FzBtU8JOE/YbEjxS+rU5jw==
`protect END_PROTECTED
