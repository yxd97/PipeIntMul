`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o7J7ZRMFvbIBFBinBEAeCMOhNVOu8ZK5eaaCAeg/dEKeePLAVLwkJbhvGUwLgRRe
uePpLTeLj+B6aPpweGnuGFlgfQODYXPwTH+4vRvO2RepBpr3oZvGQExgfoPqg60g
aeflnbziHEE809j6Qq1UhSHSyJ86c2eYTyCHI1m+pXgvURWCniW6+Kkdeic3u/r4
VXTNTRVdkXZ166D0+lxaB3zSA4VFwlJYaJNWv9eXoBahIvdt4IC8KisK3CHDGXMd
9X5axGOC9FfqZFakg1J/MkS9kHiSfFzT8JYNiuLVpK7FYzixTLdsm/surHKsM2lp
Pnphs4qkqGhK/i+TGr++9GSGfXb+qb9lVWI7RbQPrHA+JPWPkupngkONf8IRipm3
QCaDHtbEXJ2249J1/LDCuThm9M9KRixFqG4Zb/TTquckyLuZtYyS/lIhjFz3y9Ba
y4+4xVRhxpo1Wd/tA7WeHIif6/u+5D05fakPlWGn0fU=
`protect END_PROTECTED
