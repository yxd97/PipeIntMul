`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RnxJ8Gtk7AeCAr0Gz0ok2QQkVZYgvuHkcdQ54iRzKmoPHbl/kjJR8+Id2XAtwJ5g
y9Viu2vxfmdsdfXBd3HcZW90Y/dm6tox+PXYtdblD9Yl2VcZuucO5M2tdC8eXzqe
XJNpsbk0jH1FIQCVGAwMXgzNCw2bVrZlAYdQ/qLzwtkU7f79gB88Zg0QxLYzMQOK
69BO6zZah3TMRzKMzo68pNzbbJK2DjfuPpeiMR5lciyRrl3Ax6q/vZKkRru0Mdq2
jc6PfJNVaJg+IJH7QACSZcnbKl/g9kMbj5AAOCv0cNOpXcvLjBETZ8eVX5jECIP1
nyWivonkxcxs/y/xkiP0Cd+JNp3bxzmWz4M79pIOQs2mw3llkXYefWNgN79hn8q6
+Nf14Ats/4aKZkOcaS05p+BW37FijC76TmgZo0Hd83HJyj3Tu51kVtUcSzAUCEH3
/EZEIHDfW6+z8K8mx17cUoWh+etYuUUxJA88fKuM3zpNQhshmwp9O7vb1CTBVJxR
d0bkceDKAiMDHenpTCU7ASUDm8JwahpEC7MRPXQH50yXnK7FsJvgOJQmtZhZ6mOx
XXd2SZmcJxjFXPL+5C91RaJnYNDs92UtkIlnjFoNQgii3+FepOVmERNwxRLJqdZS
I/PtpMPglsBIQzCLU+MTUZFMkYha/IU0p6+OGvUDsJ3MxyzjOVZLA+70D0teY92c
pDtBzjFLD1snsgfhTcg+E4JrfZyD4upSuYI3eks7q28mgQO7ggI8/r4ERjGSkuUi
CE7XB8ODGoSF39Y4tfYzUPeiaTj4DZ4MvHH4fG46fwmky514wBoeRbeeYL97z4Dh
ibxljh/kHk85IpHs9bqDjyEimsRW7lErFa7LP5TlwWC4mB+zapjH376Z9ieCpIcx
bZVv3ojkiqSA/oGR7HAJoIyB00E8eaxRobqQChwSr35HxyjuGKfDFVq6btzgdek6
rPiiPekDOE8H97VWmAubeSeBep9zsaZcoqrVG+TAJmlfjW4UyMCPzhT9pcg1QQz/
2J4Qa9U6jHZR6p+JHXvVSkMj/u6V8siSTU+Ky7W25j9gh3XqLXZuW8iJ+7fjG0W0
JjsDf8SekkHLBTLsa6+txtdkbOmn4ZrCLKbu04HwldRQunDl0OQLZzrzgjD3XRhs
6Bqh3Vd2GRVGJTULFRol5dled9a8i4RfGu9LnX1oOVT/e7SWa1Zl83bmJMfCHlZn
QVYI4ym1HQji+OCrmqOmD3DVH1p7ODc5gtppYPRHCqPuBjZgeoqiK2aQdcHdxs0n
+DC2nyCNbC7DUF+OR2pjblsbmZEm1D8AHjhEbcL+10kXumiiFvjtxe02m67H6+n4
93eHh7SP6GMYkoORZftE7D8YCvVPIifMp7Xj9GZcgAOCiRUJF0l4NZuEn8ISkOlx
8ydjKt/tx4B0pwt7JtWTZjc4sBE+pPZpjoPyWQIEvuvkKNnTMvlHFZLwUjeLN66c
U7HXVwUMw7nH9XJtzDfWNvYPNjmRT4fb10YhU5xFYKy5nqORT9yyYyPWUsd9G23C
WuClSvGTTZksnzXb2He830fUsUQ3kagiV7dSYQum5K2uVbKZXely6DdlBTbMkkkV
p+felxGkrmytK0NOUzc8kgXZpR9XXRrL3pmFwlWxXgYYiqRGi4VrosxTV5HE1Pgr
LZpBWE5FYh4BKl/8/UmMB0K/txA7BQ6YfS6oxNxgKzj7JHdvmbjrE/b0VHBERrib
6BXLxCIr/G/qItZTOSi0H/OQWsUFrgGNgXyFUw0Ra5OrqGobprBwTg2RSpUAzBBe
g01Ya9aGiK9ZSVcEWHPZEFxGobIy/f2Gpz9RIQQM5VKTylnAEDIIlYjHo1KwyJVx
cJ5tUnB+r6O7PBxbp8Kxw9duaT1SN7/3QW5KZPq/cJIsFsNyB1QmqPnGUlczFwkV
pvcgN7us077Ff9l2YduNP0liUb6fSlsLLeWcxGzgzCJyo/WN3jD6Yhnv8kB8uvl+
cwB1SUMb1MLgFTTUEhJLxVLpg4IlmpXaEN1+jnx6FER+fldtGNLkzQRnXQyrsfKk
3HZTLGRAYRxne3lm/dh75pUgH4sucz7W5pQn1x6UMqs=
`protect END_PROTECTED
