`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtYJf8/H2/Gn4lEnT2QUK6pERwg1hAdQ57DRdEJhN24kD3VYT3h7nKWh3RUSIUJT
bsn9seWlHiRJO4aMb8GVq7gErQDm03siXULR4o50vdvHnhjcvrGNAk2ogLxw5pAj
GF6BMiXBcsfDj9TE2MBb0a2Iq6mFMT5AOYjLTNa2ITdPyFNUIqxoeRX+QL4PRKLf
qQx+a+pdWmVPTWGhchV5xPcxQxlz1TFplXRF9O6yGKKPxo01UIwcN3XY8DsiLOdb
iAtY84GyAvR0YNdWGVGk49aV49bgjGEitaUYlMTD+AMLKMr6PhjVF1ojd6DyCrre
idL943Mn7pFhwGqQwpchjRrN7POeAqCykWzWrkMACGeyE+3YranR0t5PxelWJmxx
RzG6UP/0EkIuOT9D1rH3jrV7U3yAYGnOLptUMHkcyoE=
`protect END_PROTECTED
