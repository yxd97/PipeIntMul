`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CPdk+EOW8vuuTbBEHjA+O5yZnx1/ir7RmZ12TD1LrNrLcb3FpILT0+/cNQhNgr/u
5HJ6zEfieH/KF6Si/2DB9pRtuDQHzV4GoPOOJAA+3wqF3/GvHuJBAASE9pMdgbW3
9VH4+sRlo1ta3dPL8O+O6b/B9JLzxpuktgbSL61U6+8iQtl4z7H0/vAXyZ5UC4IY
UJWvYs3TTVi6vx6D4ZfFYjplZINz9Xvt0dANqFI+N0Prr5ZoASWN8QW9PpXcIX02
oLKkm7mChOepVTvVe+RRGWy/khpUP6kOn2EMprS62E4lK6dDW/fqUdFCqptBW4H1
9WxByiYtSQLLY4X74ulYgUZYzZbOBzycOfcHuosW6xVpJXMwc1zCeMt2NPMTiGyj
4c9NlVoKRjTkvehs9XciaNyeBhZYPi0241kiFfMsJj2WHz1I0g37AsqtnnD36lud
EZrRh36C9Ua+ZlsGmATPh9AZDNoGEw0v92/ym+kaD2k=
`protect END_PROTECTED
