`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSvQDwOXfkPXgMpubNL638BT81J1iDOLMcHfcWH4JlhPTYQv8HN6lBbEczXNCO9U
IPnZsDaewXUXmqu+h9Qbf7SouJ4cB15ZsCL+NE+8jTnOpBb5QBCAekOczZk/n5aJ
DS6y8vk6tb4MgOZvEOshIVr04ITzG6lT9+ZQYHX6FgmTx/0wIL/gyB87MycpFi+k
1EPLt0fkKVGJzEZTdnBmaovybrGnwBv5zxD6lKS/rLui7LC/0ZJPLRIUArqQ7aCY
PSRVhCTMPvqmKZWD82+w1Q==
`protect END_PROTECTED
