`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+cLa4F9tbgH+y0jbU9ZJ2seKTps2PC/49FCwncVK6B5f3b8GwQivbWngbisqF8J
OLxg3p0fgyGEW+EsQ2c3tTumy6d5xXFvw2dkVy4gwyaCWWoKdZpapuUO8mVcIa8q
7M+R2guDChGBkcoBf6d4Bixw6vHpw6jK3Y3Xz5VRfA8VhHNqse8VRqdaf523YzTL
XBts2y6PjqX0BLm9N0rchB3oNETuJLVkCmMshKmCIvYSCVui+q/0+HbNptL5lOSI
5G7h8VrZBdKZAQMd45uNE7L0ekkw0jCo1D6lQtabkZuwEhrxB6SXm0rpSv6k5j/D
tz5ZLbEKYaMDIPRr7vwi2tswRNRo2ycI5ag8RuEK82bmZS3tn8/LbKb8wM/zTDTg
NdzEH4EeDP2AoRGhxEkHMD8xKGtL+kt7XrAeoTgKX6D3XCl44vd3GEgTziTLxXHI
5angO4CkO4HUK8TmmSf9VDXDNyHv0+XELsap4U/PiMIijwBOPup8gBThEkvVsQAX
L+bKVZprbE3wDsVRRpMxZteHDB5vTZrDtUydstBDbkdWhIzsG6nARl3/y7+jpR5h
kFdUUWaw/F3Tx1jHpYT5Vq9Fp1PDsRHl1AvZlTcOkODJ85pYnA+snB4sYsshmpmk
EzndkA/bbeBPkjEqsv/3ohaI+oWEGBmrE5nQ6dAn6uCa8SO6xwGKxJ+DGjuBKLCl
yn1rk4lnu9m6LhadNJhOFlbhwc3yv+rwA9srYMvur5MqTVuuBmnX6y1D2HQxaaAP
wgX+8rn8tPScqhYIzm7CqGRqGhqN5VIFcHUHjs4tbLXcUk8QoYSLrNUkzagWN8me
oaq0K6Qv2fVPFI/aRMZ6wCq4eQ9hY5cHj1mO66jhA2yIZZ/TEeCruZyXXDryhy6s
5cNTDvFdxoo8q4M/x2VaKmncd0i0BbXTso5YiyqbNzeuo4MznFEuDzhpqPVxjsgQ
qLEY7ZoC3YbeaAMhkt6dkb8bjJGU0tjGrxAEa2zw8diUu6n1+mlmOB/MLBpykBQo
2hPeMjbbUrdBC3pu95xjPzN/gtSx/l/80LH+LgL2A7wwYp7M8zIB3Xt3KLOhhIQv
nKNs0xFpXz1mA1Xn/SQ8CsMDDgdfxDreM5fDqSETY0OKr3PnG6GA0UBOYHQAXGWu
6I/2MD8P0wKofb4XgGtp1sbxyoCCrizlYICn7ZUaafiBQuukxIbRBMrPifNrEaAv
S3bY1pJXKbZCc8QwKrkhFBq0kC9y4sxudZiKkvk9EKLq6VnfJXcF/Vv4mR1E28mZ
svku7E0nghEc5JzqX0Ymj5o9fWeO8gDa02c9O2koX19aMQEh0Q5tH78QikNUG1oR
wJaksK5XkOckGkJO9r7+058bhAxsw4O65AFH0IPUUEv4HcIh9MqtAmzVHAnECC/D
zu6magxe8OklvvDY+pOEmZW1dvPm+wG+GopyyF/95p9Z6o2Uf+7cl9Ojzleeuyrr
CzFVa10vrEiQsPbdLTaQOF9TkU/b7m6B79KV9fwiNVa6D2TF5uFLCB50V3rtOt3c
CaRMgTh0SzZKdP57Cjc81rZNlRtxrMLblVxcgLvRg+gap788Pwt0U2XMhcbsQpO+
tdU4VPiV9V2TFB6tuDXY4BuPOtHzIBbQ5KPtQe3X4J+vIiI7z6oiQkpY7dbl+7+R
gk6JfSbauMsRos3XNSPIrT5zcqI1tTNcVGVkMKTIkeWrgky1qiN9x8vDHkXNNEcq
b20rTZNtiIiu4m9m8xIF/ubaNm29bKWTkYVVwNkb3RgerRQDnhYqE1XOGzpBiHA/
dmyVSNknJuDL6m07kuu5UTbsFO9Hmfbbtfom21TlDxCQYmqPSWQyTZkmG/TTdKND
HvPnnR/fCKQiVOzgTyfghNEqBFHBxiCCzHgle4dApSrv9tShFILOE8HTRrea67gJ
1/yL7newhm8xcoRGIU2OIZ6mrBX3Z1/IQ591GIFWlTWgxfIyBq5VxHrTh9pYjSA9
QYwYjJe3+lQoUuWlwOYAE/edh6jBa76y3Y2PUucK/Rft11ztldRvJwJFKJoZMfiq
OReUTL5dNSpexltzTxigAG0qtiJbJwCt3PvIzQ1j7a/0TlP1XM3REWDvTsemfIjR
Xojrfm/tigfEQb3cZhxo1NAqXWm+EUzTEQL7IMwoSibfAyVE7xC9Gp1e6FP1TEKi
`protect END_PROTECTED
