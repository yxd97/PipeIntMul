`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8Wwnoc6eiEZHnlM4h2VI0MbujNp4xHSDI+ZqjLPYwNNlpnF86C0LawZQxjiwMXp
sa6HMQFfFWgoh/koF+Syhom+mTw5M1AQvlyBpHBQ7FP41qQWJwFcvNB8jSCSR02h
FYKcN7qrGXb8V9D6cN98ZCZ4jVLnaqbii/u1Q8oFgq5D7pYxTJmd5aaGFNQR3Ybz
vmJwEuG4wCQf9Oba6CNW3cdhcpqGs40M00YKbXyZaS0aAb0Ra/LIWmJwdap7PVC1
/sBfYMDlS7D1nggq+8jXFKcQTzkVoFrwK6BDQmkS8QGrwosxCB40HrMP3InVTuBB
NIHKYRSBH2A1m+Veapzn12OBq13/gixrPF9rFs29iDfgTciHAKUo2K88JTlwMSjR
Y/5I/b/OCfFrQIvPWiNoSjuhvjs2BOpP8Ij2H1AvOXwobgoKUgqXUEFWiRVDvILZ
u1PkXwFIOWX3KA+SZb1M3GBtkxBLIma3BI53WGJlr8ZG3juMqWNLE/LANxUXO3NK
0aYoXsOUSp2S0CEo+UiM9+XCC6hkCyWmRO+cen1r43aA6GlYgbufWPvw5rm4FbLo
19Gt4SRr96o7HdzKmkAvdcR6qW/FcoBs2kTUMDnfaEcNRg30rV1W0V57IEeLR+w2
UxVM21y/zoAaLokLVVSmA9U3fwKPt0ovEWzpPaXZ2cHQlq/rzWNyQfoTGItDpm5l
9PdMxmLOzlllFWLViH7tqMayDZZiWNd582a66eSS0MeXuRn50PK9g6PU3KMwBGjX
G2w2JlI6WC0CvMqWUD3Tow4ksJY2fXLJDFZ4tGIPZASPTHsY6qubN/UCzopSEf8Q
2ePExWuKgbcnX7Ca9qK83gBSg4YqfmEeJNVm6Pdb5rAEciOYfI6j2XiFcB2gFH7l
f/acV+esSx8JmUIY+XGAkON1hrwPpb8hVllve9hFw8tSsNzWKgNTODIgSMJ9xud5
tcnGnTbx+Ttr43WydBFcPqhDPEDYYG9K4kT0HBe2DLTLC58NmSE8AM9Hs4rfE88y
ub3dDoooNXc0Tz44kdGTaCmYPAyFRJQVHvkxUcdtJXWNYJW3musOBbjHs8SjxdUl
bNuitMFSrwJjnXgDospHtKioGBwDrFbvkHsLT4hIEJkpO+lknOVEmwu/1hIF4bAX
Vznvale8EYoF22EpG+G105g1/ZVgYBnDOZkHPdKyFHOWLOmdNeLWtvGp9NNgJ+HJ
Mn9Ik3LMH59P91wHRkW9+QT4cAHIOjgwtTQRbmRYnsDAaxGfii5XVyC2ANZNZc6x
/TsG5e/0BSIutEs0CI8fV74jLFi8wR99zeMl4NAhPIkn9YIqQPHMvRFQBaWjiwNp
MkyDPyiddOdpyPFzeHTIxHZOOBFvy6rueSP0LpOKGa7HprbV3RojoXfN/VryOnq3
IrfEqrp8ZI1j8bedOjqj7gyvFudN+LQ/0WQ4FQhK+hBDgHS9hFtMj1lpIbAdUVaK
qnvp3JGEtO8DJdqAcq5OqPZlN68qkAPyV/OVf/Bjn3tpBaoK9nUPpaU2/R5gPDkO
SaXBEmj/T31fPaQ82ICsuzVQWo7aTSKQOH46FO0lZbfVsEdaxzMUrfGjXf1tov8X
GGLLWN7hdhAg9WoYcb9A6Fq7mp2IWBntcqe4cXf/CRSOokcuuZmHN0Er4YpW0xiJ
lJPen65D8mlS+/x+gpzsWJLdSkzQrnlTLvSXAvUml27oGG/pGbI138vZ0/U/BVdZ
HiERkxGEGG3ECFtyDBdlEQ==
`protect END_PROTECTED
