`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOZleEl4Foq7N0SYR4k4YS8IxWw5wY0piYAeVrPHGUrmNrWO575k3vBQig6U6kNu
5x7qUV9DgiKDT2ClofJE+suWA9WB1aI3eXINMbDi1C+MBpg9s9nOdTkl76e+jEJT
bwVwwAhaSfzg47BFPNd49ksrVPUPHt7UjU7Cx7+WLfLcIVwWl1fFgneBC9j7c/NG
1RF35SQD8G2yiOeUQftWyuwdwuM5CtRB5h8llVd1rNBp01gfFlmfiIk6yjBOReYw
1FPLM/8jZqjf20TFfMQk6FVZzd1SLgcvaiuD0t5vbmF3foZ2YYYmZcXlJo1pn8Fv
17DZLJvJzoQd1txKkifhcDgfTjnZqa4uWmDJvHD1BEMaHFIR5e8JBieAIyjOzhd3
e6+kBzS9wbd7U0LnhE1gVu8YjrsoTgT2UsLGpnKGaQwPoZNIVHdakin1xhSpmKDV
hPubWW2+cyhxY50Hl/lAR5uxHY0iG+FyU0o7PQWxviHaxurYgpfzXKTtxlgPU+Gw
FZMMxRbgKk7ij1wSWai4g0piO//VBLUW4Y1B+nOwLD4/qtdQs+f3vN5Xb0IcuUmn
H2mC2XOO+baUTtwbX1+CYgGBobbrDLzY8bieQySruWfIyFpx78Wxuq5QpYuGjg0G
iwM/JnS1BRsaCmaFw00Ggkz8iEJ99hKs4ZeMmM13gFPZyFrSBXxK+MxqN3RT6HB6
cg9tBA23QCZimeNjylpa8OdepGy+ssSGsEjhitU3NSnODlPlSWOlX5tkau5KXJid
V2dZjmFHWw8P6cwVQJ0XdwFP8PYdoJ1Lq5IgIHCHkPJpw4fXLPS7AHcNn3bXeS+3
mkAM/hg5ZpfWx6MsQBBGlyKvPjBHYec68OVhJfYxY615RJEkIhwl6UOKR989tnEH
epN5ujdGEm2L0VbRb6KOJjzI8J47h5DDcLU34B7qGE8atWTgK512hp4YZWy6lIYA
DgwyYBNZXMSd6zAkwrc611PNJEcPrvrtCgw0LpSdT9ASPOzUSKaC2JPZiHXdwJFo
JJP8ziRItN1r8W/sjzyYNINrPZw7I0HDq7omXuMGj5oHFMnIBrnkhLanJSbwfbB/
mmTngWPC55PocU1dT4VpRVrle+qRIY11fG5Dsx9fgonyf30eL+UZQlnggYBb8fNX
TL2w4TKTs05j7e/Wao+27MjeX4b86NcZtn3SiCcwt1ha/wX/YdFJ2vXRNMPKcgG4
Xj/BTelr1ljzwLcfJpGNMH7xUs+Quj7RtfJHbLXCBX6kSdLziZkDutF2x0vkEm37
sF5sy1CtrGSJ3k8sLmTe3R9SFoRAH2aY8dGf1wFGFFsYT2lppnRzeTuh2tGmRzlF
OVzoF+EIvRGDVkL13VVUb6xKbK5qnyWYFhZ2tJ471OkTCv/RFvb34FWoS+vLE/rZ
I5fKQv+Ul9HZOq0qH5q7/CQB/QgYonWZbd8ejOAvpQfi6vO/DnYb3VsQr6M4i1d7
JUO+32DtQEiEAhyR05WMMZmSPstskJKQX9xnNb4kBAAvFYcMrkSGdzaG/kJnEYpg
Sz5x8nkQZ7UpDpCMgNnC+HzVOEw+oR46uve3W6IgYZCoWQNW0QAXAui+0pJggYn5
W0tqfKHFftZlefqWQEXY1ZP8vJqv4gBwBz6RLb9iTA5eoEiq7GgP5Xh0xW0bvE2P
wuLEfdQ28dRb/AX1/mpQrlMV1xjc8s90L+9J3AXeMsMEIjPOP7KH2Jn0okytUzaX
8wSb7gSke15XGIt2ghCkGUSmtH7FEdzeekM93V62yioKysFqwLeadQevnneP91UL
XRbpSYu8gOY2+q2qiRDLuXp2IwimzHsk8sbjF8QT+eWEZnMZwGeqitctzTfWPqYu
TmjUbixgY2b9NWP0L+IYiyCgI8II7BWoiU2mnWdBJoveiUW2y5MiZ+UsJHsGGOOW
dW2ZE7VsGE0eS2SdWILKK8ckbK3e/71+7QE2CmDwge8RPIr8yB4MhxDnroGPz/cV
k8xiF26Nf2I3vxWySDWsE8XO2pRMdlFgEpG+I0zQM4yAJJ4hR1n5Jv1AH8ZnxWYV
ZBGIuMmaYC6p4lawKYpmV+MtJMZEmWsc0+jObh5jDvoUCFNK48dvikUus1m0XW11
BaBCraimFZo/ibUxscnOKcYSiZpLBUC1ggVk6fDhWfbm8Ng3YyvynEs3nD43ZR6Z
YDAZMQZxaEBTDMMYCnulXWdfu7wJbmpQbWCyXKyMK7AAkyYfEEDwxhEb0EKrYq/a
fNkNCcuYk9uANhUiYKgsvKaG5cmy0+Qiiw5Nl9Quep6UR6lu2L6SYaxMBX8nkO48
u94HnNVmEyAYLH/ODusuNIrMUVAnNwNqfraKFCc4kCH+aTRU3RuLYD8hG3blM/31
yxi22Yd1fSIHCysUnaNmy0Yj5FygI8TKiVFBQVO9rMlrSmasKmqd2PiRevYdTdY+
uzMpwNhgO/dm8OXUvJcjFk32wns8CBtYQNSqNJoYD6MiXTauGWgqKzooLH00rGOD
iDcvyjWJrUjq+kAHd8wgA/InUmsXzdQO4QLVBwqcEu2r+MZRqqMAqqkx4qzT2tXG
xalqkC2CbcFcAOLbXaIZmgPkgZ3WURoNnOKIJi84ib8ZjGqa22nQA0R6aoDh3htF
Bax0kJFIn8J2ous/NY0QzVFTTEeMN9CyjKKY3R/8D0uS88XL4z0I9cxX2EyU1E3w
A1VEGpGoDdxNzBTLXcAGLaqsVtnh/bwKPcLR9/tTJgPdWGDC4hhqDA0F47SlVC4q
D/UEzN8SBvHnL4XieOWRIp+3u6P0R9ANeLskcoK226+J4bHx1MuPO3F74RRbwnb4
PrOckOveZoGWd6srIb/SLXJOtGI7Bf5VBsgBuZKWM2EG+0yLd9LmdSBJaJRV+sv6
x8atR1lvgyg4/hH2IWctRZX7B/jL2ytBmhvomSawXwelgwxcig4zkvsitCtm8TEe
3sX0BrEKetDjjdEsIDzEeKRd/AWs0qtmyO6+KVEsLW/HWQrUi3MARxWFznNxqSb3
1URI8Zw+hM/gCzcWA+sP7epXrxdCFxDvtdUm3/OAkpGNDQCYFCVuIVS2q976BEJ5
Ln7lmZuOM+GLfJ4yjH4G+qy2bTKv2WAC03CoKzV1TSgaBk4DzytNEiimPzPYXuZu
97EXZVeHyQAZ3m56t2i43FTpwJhltBXVDkmtL/OrocDrkrLVnqbGqoxa/Q8IAPqs
3gjJp7FgAdg0191EZuQlQCMblarpgMmdQjrxzNJ9uRhePbD6oFXlD27nzeyEVIBy
g87qUYN5OXfWBTFwHgQobFR1Lv73y7+3sf0+MpBBwbpmya0UMfpe728hXdHKxJcN
XXoDZPlhzaCwXjYhH/5dJyS4DRfpTj0TKwt+KWYu3hZSFv8KOBgwq8b50Yb8UFRV
/ITH5/P14vJMjF0Mc5g9AwEko5XFz2aOVMmaboK/stkZ+Aq3Jqn07oIH1cK4RpT/
QIynYOQRKuXH6Hxwoh2GmFVOHOm4XGAb0Y8H24iTji4UhhqYaTKSrcHxulOAlobR
oZFgoPAoDTKXRtum9IDGBvfcaxONnNetWngONP2XxAWnRZieJtKN6c+rJi9Nxnpk
LBNiJPtlJrb+jAA04XsBmrxL+j8qcxFghcpYFrvzdzHHScyFX+HzLyR8K18bheI9
NNoM79316HKG9kPF5qIfenPFBdNzImzGVIc7ZNX4pJHV/z53ESEhlLi4qEZ7TIGx
/C/VmJaVR6njVgaDAuR5gLIWK8zMAJsduwxQiVf89Xm2uLMQS1V1zU6t7+GuLjjT
ykAk19NOghzHVRu1b92BNadUXU/8/MGT1jApJSrQo1zqSZMTTjnXJsqzfpZxMkhU
EH9pNnRmGEj0d/YsvIAo6Yg8nhMmXQsnPNPnmdBSu/xi/B2qvZgrSKzG3/3gVyjQ
T0bh/Z1CKsWP4q45uY4QXxH69hHubieRW/rKhmNxquMQr+35ODj9I8ztooLZ7pjS
2HKCSTbeRLSCU0Rsl28mx+mCER+ASHB+dZJpQoUyLZuZz5emp2LEZOIHVTUiG8zd
Bmpljd86DaMSu99RAM3IK0oQpL4FGEsLOTmX4yKz/cDvIMEorar7oI+un3CL595+
OPMQbgG7sA+sU5BKW2HDlfg7cmw/f/rWnxe4Kqa0gD4Do+9BJ1g7zuHLFJJO3MHD
hdkTJXYbcRhBIv3s/k+GbewYb8kOLu88ZqrHZpPNrO28qc053s1+vLv8/ECiktQy
2lNQTdRsTJS2UOVJMZ8Wr+tn/Fa3mlSaZNMLBopzEv+DlZ+q8VJjpaLFG62/tBi6
G1f7MyKp/kkrskYF0FAoeIGGuQQFQubV+djE2loQLPkaVvZLTP5j+UYRweSwDgex
sXV0AN6VLRBZgjpEqhBAVwKfG3A+TSWv+DmSh9zyJyBuXBNWGayOcLUs9ukWOuIp
`protect END_PROTECTED
