`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8pzLvuysB7sRjuTUePPWH3RIEZShMrFl9THiDy6BOqzeGOFgruelu0VhLZt9bxR6
DZ9mRq+o5eOCSqZSjnh3548kKm7UJaDpvwDE7KNLuyGb/keKRtrszWf55dOsoF2w
MPS9Y7RtLgnbWH/VE7m2wu9WhmJ8NLs6R+DgMnuhQo21WtvSGKud9lCNNbhDhJ/X
A21Rnymb6I4wiiV0nHTvZREV+N+f2B1r3qMadhBkVMueULt15j1mrEHXgV6cXYND
oBC2sNQC7Vr5B8kOQhxf6fccXB87LceCo+ZJzIVQj+/GbJOYGM3U0zmEDW96wq8/
tmuVDuGGs2aYTV4/XpViyQGieaGq6oIwdN8sbtQyF72hbE2Sjub8JcaCMCEfdJb8
PiKidXiYxf3idm5EYrx6kYxIu6MgV7BQFUnmmyBH1Koz6orGkk22EZoRLrk6xpMh
+n+6TuLODj4zhS8ts7mKKkRPRYrVItT3XHblm2yXVLw=
`protect END_PROTECTED
