`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OTL+XI4evmhOdl3D9Q+e/BTWepv2P6csWne+/7ZgicV4Wr46xDRTlFZ9z+XDR56y
9bqZTYBlCWAB4llmaMvZA3tCdC9bwe5GFi4Qsvi7P8zoHKN80dYD4/pVVZqThn56
emeonylL1ydwiLYR5zC2dWbQNz0Llmi3khYkmF4HSJ7TMdcb/Dy+xwVrUDGhl0z3
nTxrsmFbjcXWVQxtCPipXjN0qBX7PN7/8J625DkA5HMNIM3XJqlFMdRX1fOqX02Q
QqbKRU1KIrC0uStmYIKz0Tw9npNLpuESpk9bOstJHumcXNFsa1Ga5hP0YDmujFBq
ZYq/AnqGBHfLmxhxDro7FUxIe1FpJKAiOQRsF8/d49kRtkcE3webo4u10eobB2pi
7U5NFCkeB3Wjue2ZUA9ZeVH7crAGCyocuREPZRDt5ghi888VRIzlpeoKElzEaroS
S+DNIsk3Yr5WwDC0kanNvhgtmieZ8swDell+FM5aQNPe97bU+8xaHS46FVADI/i7
W+i1ZxFS1COoG3zRrc4h/h5ze6xWQZoq7dp4UHj3Mxnxx8VD2KFZU2LT975jieT3
Sm/SBRnpi1hcTV8069FlAg==
`protect END_PROTECTED
