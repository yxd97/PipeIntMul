`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63y3XGQO4Vx7AGp5rWIvsxr1WUzT/l0ibeKbgK19x83a4G6rQlDEE+Xs3a4MPE1I
sA7C2wa/PV7x9voHi6JTb1kBDyqBiXsojaEUpVlxNCria8fRNM6L39rizqtU5tiC
LVNZ2Ap0Vw1HxnGMB9E/PM9Dv7u+LAmJNMqyLw22J0IUodrzP8W3KTXhFN8pFk6p
Jd9WwxVfY56QUWeI7qDMVDHrT5+jEP37pxZDEqd4M1GVIL7eoc5UY+ozjnlBh39h
3fFteewmsPbmc9Qbi1PUbF2OQBYPY2LW4cl/0yMcZN/haSnxzLH439aEke8oWQ93
YyX0KWT04nrJKzGPTbsueS/Na+QhwxX04Bw3nhel/cyw5oSdsDLcTCSBpiwdYGg5
212Eg4T0UbPBAQ1ozrCIZOJxuB0tQlagzketToLAYZNtThYVcycW/D6Z1wi177jK
1ATYMqNXO+Tjw8Pe5JPh4RJFDkEBMJ1BxQmsEprGi+3jfSmFBQmpEWFhForh6+7V
mYjr+bUC65T0qnVozlGc0sXfsD/C0HqgaRQJvgGddtfHZMuWer+Hr6O86rG57A2z
Q3ukF89T5TsSbmOU7St+IbX1BBsjqntINNlm+XOVlGD02lYJAQAU7doFNdKg6AIU
UaT62TKYKNbCLXCrvAHvELbolvOQAKAMmSZWElyQTmxbeuvQhJAK6KpIBi57HVNN
dh3qUDnibkLpm838JRKSRLn8UX8RngSwJcOainzfufKZnzHi7Grd8cSHU8DaC2no
f4Hb8h6vnp0cK6qjc+mzkw==
`protect END_PROTECTED
