`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzdhUhvzs1QE1qLbK8Nyyg6w6v7qv3+4MzUE8ffto3ILorWOThPQoa1T6lFI8nL+
P33bKjtsXh2BtL701PxMUB6ODeARaBZOLeEdDjCkhHlEXJ29CwrBgMABvfvHULNE
C9BBB/kIKjpPCL5cAriXx0Ko27M7xN5xE32IwM5B7BKDV8mRfQyYvpoM3POjJXFq
LNQ7ONbyg7hw5GOBxZ/hkFoybBQI3OoInccgPFrEHfHQv52b5PDXIxRXiD5nzp9D
PhxhQr/QUiSN0BFGl5eJG8pXNgUF1p42OMEkhCU0txRDSW21BBfVUKxByoiY1qUH
9bi+eBrqcIK0g94dF2HbblRT3nAjV17q+oq2A/QuKTKGXlWzvxu7D+8ATeiaDzjS
edUn7OrL0bstQ/icbQuKooDSikS/xv3HI+BjE7fYErzHbP0mVDj5xg/awQwwCof0
QE8oeNRf4w0btP+AvxyiG11HoYhEF3hBfTkgDkW8D+qbKHvpbkispjnocen8sKcH
Yb5RcQaQtVP0xl7cut/tOwmaIhFDX9CxiMKwTwBuv3bFTe1XKoX2qbstBcU+YKQn
UMJ2CloUz6Ebrxm8RsuWYDgDkbJOBO6XFkTjub0iMCvyGSH303ojtmalSI2D5C+y
psXxpHNprusC5qOnBXRVKG3P20MJI9PkXXic95+8VCbRz7kAzDA/n+bEoheaaLlF
FJ5r7b/EzJzcIjPCuRfkKd+GINWQe8OPv2GWRnFd1JfQj3R27z0NWnjJlIGGStlC
dDgcSCC/QTXksu0juizAT0NxANqMyHXhN9drpErnsttp5T6nPwOxOlTXHBgWOXOX
eCNw6kZCsCTuBYq1xr2GB+6iqpjSxKt6DLLTZnlwgQjRtBvPGv1/CqBX0yAi/0mC
dK+VrnAtkR1+s0uNWVKiBA83dQmVF8JWNQayNQEYqrgS6w08spnvJfnOA6SVC4c4
GXIYqUmeeTApgHBJeGd9I1Ce1j2R6huIwuwp/CNpojoRfmtTaOCeMm37JUOHkPpo
PYSzreU0mBtdzC9L0RRoNt13RZ6ESf9IonuzPZUVjgLbel8III7NM2usMBHbP1th
/RzIYXhppj7IAJE9sct2T9I58CMLlplB+vBvU51WIqfiUztQlGKUoNQeKcZygYSv
RwQBeleSM+3tn4lhj1t3ZZn9H6Jg5niT33CK3ROvbYhkn+MBB0w1SLyXLC8pkXyQ
9Iv2j6l55FFDWUtiCow+AWatxbPoiFaQ3qKeTSi7EBgLScpv4jDVHvjivcKCAa2r
KZfmIoFgG/X0uzvXrp6L1WPMHvitAVkkuZBBgxr0POSGtpN9RNuXEKQDrv32CG2G
Q0abHkHdcS0/+mv0Hpc4fP1yI/p+V5JlU3K08w3XXPq5ijELxAA/f30ViLFVRYlw
Tebv1fas6Vikbe1prY3PA1YFxr640yhm0MTHdWq25u7RxT6lxy+f9W68lgAEE2Wt
c8K+RWIreR2kGynldV/Lq3c4r1jIDlW8VOUzwO9v3ZpKvDOKszP7UNM3i9RnGYCK
GrdgqXr7XkgslXke02sQwpLZkkr5Xa79UpYdgKXlpXnGYPU3mJn3m+zz5p3HcmAP
tPl8I6wptwbEDHRQFtEX+e0u7Z69w9bzJVVxUnPC/PxoBfsoMmrutjuFE9MTsfUh
j/ApnuCIyYmL1vII8QTbnKghnqu2szcnYh+59A58zaIrT/UPMnCOBQyvbXOynuJu
fvErFU/ucB1xPVaH6kOjAYZHsixe7ZrHh16/A4KuDEMHLDejk+cetjmEF3ZQEGYG
DvdXaomSsA+gwpMx1sNRBYsIVpBDxmhX8YLazI9l2ESDzRwqmxSO3ytRp+2zYp4D
`protect END_PROTECTED
