`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhuJtmA2dLt+RcoT+wwsu673NDlgEdIOu8ux/OH8UmkjeX/+xIx4jBh0xFcUswt/
lGxQHlYwov/PK4CSNDoXAAU3iV1dza6x4eIEp7mq7VsL9x9YWn1rF95OQ8Bhy9Ej
WJlb3gKhCXRt/77R8SRgBBNGqlB5AH/qNwPuxVjBOS16TbQvO35f9CevFtQqcmFF
h6LH6Bb9ySYMWdeIOyK5rJe7I1KjSle3WqtO1ObVnGg6KbyokkpA1LVDkwdCxzZ5
+81OS3rcpmpnE9jyCL00KEAimpKt7WeKnF7Pm0U79cU=
`protect END_PROTECTED
