`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wG5ToV7W6beSfUjSitvlmNCKSRL5fJkYwyAqS9rlsZ9COScvRB0ZGn+5kpmPuwB1
zKXc5VcPBxH3RbKSfXCgjYkmyVCrJIzGkt1oOmh90SWxAdg/p64OQrnxzjBv6N29
G4T8DyyZsOf99+m3N6fhMt58U2tSmBnffXiq5OzK2eaUq1K8a/6K9twFVtjHL0Gs
ozGF2kNNn8VcxIX0q3IWPo3RTA53pBUljiVygtEL2zGScyI3SFXsX+Kf4mluWJxG
y8wtRyWz0yyD7UrshEnAbj1JUOmaiL0Jk+m0mRZcnVu9QJfNRNYFhAR1Phg2OMwY
fbIATYdCYvU5zktfvSLpNUQux9hTsJY0S7AKyC31xpJaYeGPts1NXgnMruI1HKPC
DzOLRNdHZXfw9mJUWe5UTknbfwMtnV25fFyuujO9DH4Cx+Ibm9Um2hYo+Ll40Lkb
kdFMS2hCDAyBTIrtKOYctBTuduUl1x9dH9yS62jOPl8eQurujx/XOx+QUOv+nRCd
`protect END_PROTECTED
