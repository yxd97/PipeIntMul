`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QivXsKECl/JfRiA3Aun/8rWN+HcBZk/QawPrrvbP557+2CaqgMCDi5/0gWYIl5l4
bpHF4P/nqw8D6p60wtqStS+9Lh4ykRRlNAJ4dmyIW91UMnnRPg1Jaj5Ip13zezHQ
vsCxow60R1Q5YZreEQbWJ7b+VA5VJ5xA3csJ9QJyLBj6prhEmAZzr5Q4Tr0zV2AR
DqeRCz81Y72PYC22TiE9cX1MKoa0SQ4t9xU8U2B4zyJFmBrQNbpYfu0xM7na/9IV
8TZBowXGtUNvV3fygt+H0/tMpyd4d2wjxOIuruZpzSg=
`protect END_PROTECTED
