`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V7xDjGe43bLVBMN918qqgX/jNwGGZRNBJCxfQ2W3QxEuj3rO9sN+mM+9yw1uxysB
sDOlngS4U6lXcQCAUct2y1HrOsCYqNBB+Tl3hBAdpfU8egU1m6nKYdWdCY1aaWoi
1lLTmzSm5qNxEazOdKPKc4px1aUUYi1MHoJQlMj4dUNlyZnkScuigKKPQeWGMzOf
6+tjxtsIRInsDUOtMOhCAkB9iQXtKFpDKLmZWQTO9K5rK8eB39HKMyfkV4dHeMbu
fPRpFRlHq7dlOT7swA7WkrbRA3tyJPGZFa5MXOEGGzsITEVITQMKAdk0H+Wxg9XR
7yyVkkxBy8WeCsP9I+hMk7o89TgY3q5xgjAEI2KaQggch5/p1zEA+YTPI5qwj6kk
+O5+ezqXzvSuKbIH73jydyt2Kg1OInRjUihQE+NQX87Tn2nTGInrsYl5vdsIVOks
xDJPnsdSZlaDy2Oj/gNKTGDK4TL9vQlmSMSG++77delYyoAQQRWA7Y03OjM2Lgxq
`protect END_PROTECTED
