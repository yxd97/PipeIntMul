`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BB3KY9wmm/TvXBOXZJM7XMMQXO+aZfT1C/DvtXvXBuYax7U8NuWW5Jq37oeaE9Ea
eciHhX4uYNLWd/W/lBfMdZgEHPC4Yw5WwGKVGIKIXZeu1zaHcN4Ntr9TOyU15kmK
tC0KjeEqUBf1doYjEV7rMIfabh2nXOrGeGlibwhz1b4egaXCOORblKYkT1iVANzo
X9usdL8RnBGYgH95bHULThz0vHjw1OpaCyl/mvFcBGRPlQUrtt6cqecdkujr8/G0
zxceaLDRFCjC9VhFHD4nd4/RCniWiWf+xsO0bxYFiPoDxskgsFW3j+HPDHYAftgN
ElNGiWinXvTmtPqNMJe1hOA6Oov/8lQY4IybZvM8b/GR2U9msD69bbq9ZYImdMa4
m/Y/MDBFI8/s953CVja/XYPvoSwl6dXonZL6VWGzUGoG87uNwybeFaBo/Qi0TR0g
u4NOgOCtOImRnxqib3xfL/pliyFJq5l7/wklrKezJbmYeF2kB1he3fO+Wqu/ufDu
xsaLlRbs8tSjYvsclAqJjl6Fb6LQ/jjOKxU3dDm5cSpGTbXxtHFHibCjD8aYIIwg
QcSmcjzstaxscZQzcBQRLV1ilJyMcKWvBKRRYplHhmGJwGb1fiTEU5oyUEKkXHiU
SpNYfbaUHoZUeSbqi3GYyFHWVj8TZeHRiGRrFs79/KY=
`protect END_PROTECTED
