`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p5If6W/FySk51PAYKYAXj/DNeirGqUx0ao3NyuBRDr2G42RqVPKUitBbJq3gw95P
YrVK42Adf4rJ+qmG4zEnZnN0LiaFySjfk/i38r2J4r16LpjOfq81MayU5obNAYMk
gZRyhAgcowNm5kQ/XBcdJZ6pZTHMMnyvGuQUEz08XoLdOmETjBx64GohpMMwSCqt
u+FbWtqdWOOSTPPs7m32UUxVE9A4+kF78sWuhB6KM7HSiiFotp+JvJ7wuqr9cNka
YIkLjQXyW48czPrxpzuyLOWWQEdQXbLhQiXIuLjwA3AejPZw/XEWV85D0WT6O2li
+c6Mpz/DGNJ4syN9Dvh2VCKYlVYRGcWQz8+BBIFvSTyhKYcPqmv4F55QajduHvDY
sgBXRWPuaLrUndKBqRGJlqsTuSNuSWeqYreC78rZXvvw5Z80YFwXGXuCYYcJDglj
HHz3fU0KmVPwzdfzwfWnSQUaD362QyzRHxUnHfeWzbxCPwFP3vBfhFXeHpIDAIUe
OHNOuLxbqLSZGRWSQlnvwMxIItPpqIgCvl82LxoBND9YV8xH9/iAAaqCn/tNho+m
zVUtgB95fViw1+LO8lCPcKJFdfvyB8saLfEymWvFlANXpe/encQpTejeNDRMDbPi
3numYOH9kfYfNiUwHOM/Prq3/KzWL19gakrgFTyMe9qXFcx4J/WWst/ZatuD0CDO
lhgCXyHVL/HXZGr7SUZua+rfb7MRlGtrgoUb/3U8dbKAHmXtSM9bfGK7pAXkHmnG
0EyEJ4I3UprsJlySVorWxhW98erbwVbBwA7pajSkrQFtQLWXDaVgucuhsjaUy66S
UBc8bX0qPGtzWf5ssHcwi9L9zomr/Opp1ow8UZBm86oNaTIzpCnQ0TiqkPpmaCDf
GtEkw5ei4k6i764JrLbYhjXsVlgnSB5RgvDCxl3m4qwOoHwjJpTlS3m9FnfBmPjI
ZYbPRWC4uh4ihL5gKgnzp7rERyVb/Qh6DqP9AsFmjIqqyQHNa1lHy34YWGANSvff
4M8C9KYesgj9lkoVTIGLk+w8+wbbjKKheqVKnLhsyTat+XcEel/TM3xmBfLfE7G9
ia4F8e1b0hl4Lgxz2cn6yMfIqQpmPNfSK6qBN6issoH46dA/HzZUzTEnILEhOWA1
8GPoL11bPmUfqWuRlyY4uVYWuo4mOdvQ7q3AEI31hleATJPWdWOd61LOcu3OyC6c
Wzn4XTHLPCtZzkwtdNQuBEveMS4dwzcfUBq9PSfYdl+Xk/CpwkRLkk+j5ujHjEQg
vNQFLa9+6r1bH92n3FnU9AfRWCHhn4G0EbbddgpZwkQSEPbBq/tG1rPv51+EgN3C
rySXQW1FwVvycARZIfii7T/bi0pYjEvu2bLR/NAYf2vof1uNTxokhFhr2XSG+AFl
AJulalr0IZZ32D+JUhvsY1QY7wsczjTMvmyVef59o06ZhWYdk7TUX/CYh3Wltmhl
8tzD1WpPsZ7nj0akU9bOtTKaUl7G8KlEfpo1ubOx4pZpH+RA4ruy6nKTCk3jqsPS
kscZ3kKxU/JqYKhX5Rp7mnHYB12jvm2nwfTkThNWw1jQsNnQ16RqfmBNvadHtYtY
izuOoj7vbh+KYvN5by1WvVWId4Fsvleg51FSMJWfm81Hk2MmPCy/wLgV506j1/9D
7nHHuxr5fe6jSdVgJCxCTwMzGhg0ON9L4LVztfYcUP8vT/slmxA8mPclenBPu/dp
/TN2YcewMdZ94LtOrq9snDO07/a4/yDGV9LM1cWrcl7rrQ3sLmDK82pOU1WZr9zJ
G0tQylTCB0fzDVt7PbN2rFdmpGEGZ1P2l6t+6WKdYeypM4VqxFWo/pud369yJe3N
vKQJ+O6TdtoyyC8wyB8CmXEsE/jT89o2IiXVJuvzz0DavmNR+O2lfWHlXUg6XM4Q
chzIeCNfDTZsEG6cuyBtkyd+4D2bJ8HdSZUIe5GYeFKXgpbUoAu2GGnTs9jCIXLJ
lWDoER9gApGRApF9t4EEREoS7bvjiDyeuTeewrybr+FGMLJJcYrN9XM/zhexSepi
lJaOsuiZqht9n7GVroEbCudx/0SFuskho3Co9R4AK4Ra3ff2b9o+JV/jpR+IaBqL
0yw603qoJHjoEeUssQl3itOPfI2Gjl5dxfsk8quDxt8G/7yKwAN738BfOYaIZrPf
1sN8b8S9lrqHwZjhMWy1+csIq2sC+D1sUYXy0Qz3yyTNwiU0CDxToJ0nVk8NNx+c
l/o4V2eS2VURsEL5ifGyO5GCUBEaIlGsOCOBkGYbY1xveB8JxNV9d4HlriWvWPOQ
i6BT0uMr2LzzuGP8K5sN084Fm7yVeBFp/qo73EFRwsiPTpgrDM4AwciBqVpMGPeC
nGX6b1LRpBiZtsypELCII8lVBImsFNh4ggC9AI/DmUehoRAZzaAe5CUFW94uWZL0
jl5uY5aq8HM6LpgIlTd9k3yHhPZagrLkVBqSzma5N8Y4Ng3NAzm6c0DmIip24tvo
2eWSvtgQTdn4dymDuVld13d2is32tWpxLz6FioCnK83WyGTJj9WlPAunr55frHML
8vwYODTCkGUiQ+48uSZPc0relqRXgbhNjIh3geaptYmVg4ZZnpkjfo7Hdfq8qGtg
2IdZCwp8rBPHnISHJjXZTf5cJCWUlYNctT2xQGYwfXreDdQ5f2uobgfJOYze2fi1
utHvDFgsbnUxB3d+se/EYJI75TXbAG7cugZowB90TSsIDmqEtbHmCLmXpKabhDy8
YuQSFTdRJGp8pKOhKk7u4giIM1TVSmktzDbDs3BFPjmXRR19+Wx9lTMODiIsjUPG
gYdkqLpp97kX9kuxsFRm+veVeSRrAbEdPFxbG6AzTeZahP5iFPX8GKeAn5SteAMi
wTPrzLrqDpc90wcOcNDzhFIggf7tB1S8h3x1Qt2lEHKn98Qxjrx5BA1foYKr17Tw
1kk2MdfMYIqhL00HhjVHgOqazRNhskvTgK42gTJK6mSJLhS7a7AnpuXpWpkZ350e
FVAiTCEEPZ+mgRBtHpadHK7prvhCRomPaAQzUn2eew+x3hzIL4V9wXy9NbTdKjWr
i802ZrzD+B7480c9Mk/1KT4FUL+cRrwwLJhb/7tGGUpLWuX8uN8LhATOu5d/TNRh
bvZbNvI8mJDNiL5YM2CqbAnpxAGNrLJPl/VTD//7hzvdwKf9Ixf8FJ6KmaLjLtYN
UHAkNCR7yI4JJnzGuV7qI8+BHtdYxA9eGrpo+/uWiV1wQzFZDnJqJVLM7k9HvgZ6
DoTaPKw04pO1/IJue0RfTbIbjS8ETfz+3OqbzG0rfnjw2IFLgr1Cl5Y/A5U6ARqq
VlBkarCfEB4+pCJT+V+wLjngJzQlZpTGVWhrmRniIYX/32MGoCa0ekn4sdjG81j9
soC8PnItWurO/6m2kmmliUGBuQrnUNTxURA5hkoH9JWG9b/Hus23E2kCVVZW2kUx
fZ0aKMTtHvLt2eLO9oR43kNnoLaWn5vfFg9mMzgXPO59BmYveVDOi3uaxLhAYWrW
gU2gif3V5oMvD8KPBw6KRPcaKn+6ui2ipu2CRBCFKLB2wyJzxP0OXBKCm9JL/jCL
jKRVYLVVAs5v/SjG/ZF+lFDZhswvUVzAr/PsHW+py9+kQUbLPTMXDzAXlGaucbVO
wccebJg1oCCYp5tUZS2uqwXEH7ntQDh8IQKlEKk8sZhXXHTE6erRsrec5ix03VnN
xLjw3dHfRX4qO/6hZt1qas29fNwwYaCSvniyLBJ1bFt7opopaQ+UAnGZmwyOrWq3
m0s4bNyvsCeSdDSn0zz1sDNIY3rf1a8vpzh8UnXFliX4MP/MYveEopgygAIRNTeN
qeXwONy8N5CUWw0vBptld4b2aXdJyBCCEr6QJ7i5WtPF0jSET4Ozo9x0JoZ6F/W/
tfL/NndicrOBReKRZDGv6nWoVGbMekm9Ij3YOpcMRyUgU7YHt+GNe4WOO4oPGaK7
Kguzj+AXmI44he+Kauue7CZGj8mjX1MBU+jMDbCBfzuOjaqvwjYC9XM38Yh/gS0N
bF+AH/GjtjRpGefnMuHPc3R3evIiqXXmVtX81uiWh8hz/Cg1pK4afav1ivIstjs7
IynIm5TEW2MUKTjwF02zOwOZp33ZzaP2buoOu5aJppM93UgdOtLamHLCUEMgXuln
XEgavvCyv9z4DDK9TjQ9KzHZsYZZpGnf0N2TPMbCJdzxPDBV+COigwMGGkjEWzna
NMkScyFS9fA6MAyyne4DnyM5xofYHd0+z5nQR2RHN8cXoDJE3YACBeCrNVx4wmb+
QFAHEOG/pqQLNUsZ9mGw11pXccRGbX25/YR9kGrN5Ns7kMWoeOz8ZIs/Sk4TV88t
JP0JVc3YTEiVOo8m6cPtwYrGkw2BRHRz+256y8oFQ/SA3PvKCZnSZNmh796bMp96
WDHgsY/BtZNh3RcWEZ3sK5eNF2EmrPjWynYNfEY9PeKn0+HxvCebbZGcMK3RH90K
dYM84tBdaryyFjjlMjbyutRij5T/Dr0UPvFZ0geWTUorC8DgbLBe8J6S/CO3C6rT
6p8YqGYHcubxk1jLAtXFmHEH+/gHjCSAw5Tx+qkcKoVTWTx7ayIrGhlXbXSoLlP5
ARycjl7DlCKRemGDnVEWhaqrie4cZIXusUzBGYJCwAkhEV2POlMoiikBD1Fu+ORh
hHCjPmZIsO5R334Ua+PYW8UHQ9/Evhb7NJrD2YtxJbAghcah9P31ISGMkHkg1uZE
RcU4DAyTszzj+uuE9AWfPRZ8cu5CW+/2BOp6swSJmJQ6rp2cK9/YJP6sqe7fVpR+
zph62GOnWrwLaskWakliXYyRV7WMLwRrlHGLKt4yfIse1J82zXuk/HuTuicXxz/2
Rrjpqn45K+B/vuVDSVZmhhg5OMsQW9TLUI8USbWBTkuq/rnCskO+XFt0fMfCUmSw
IBnwbWc/UuEhvCbsJVfkcX/HN1E4Xp/DXTupCkPD8fIGmBWsfnllTFfuxoIY1aCs
DZTjXFjmGradlX7VNLLyUu6ReJ9c6t2lVUPjIeSBfKsyLOM0TZn8Qcjq/xL5BvbS
7JCpo5Uwi05bHhsG54TqRbJMwjj8EoZRIH+EHEOQ2eFKGxYyw7rszR62cEmEpYrz
Gnht++drP90+PYYqOLSF8GbWMyRXk3DiT5wDb0ZvDdHBlMaPkpe4eq7559WPQHwj
Q5otJmCmKJToaz8mWbYebrxNA6u41MWXJuRPhm1yKJeB74NSmk9uGAC3WspfapPK
z8IergQ28aWobCYbtgR6RlFVdvYVIKg5rdQyaqeeWkOdxF6dK1QfNfCZylQlwXwT
oTTls0FVpNRPyKrzifiHEumt56DKVlx4JPsw6cPb0Zrb2rw5hkRpTO09/tZ1vOgJ
FApFqwS5DXu6y+PbYz/Wqkdd0KEM9FWPCpn6JcR+A+9nmqw7LrUxufLIJ5sSE4Ja
nNR67N9pdUZQo4vnDegoqaTwJRLlqUdMB2wZ1MyFkNvWmbKcx8fGC5CDeK6BdsJS
spq365mUL2voxBOlWc9nVQb16c7+aHqPtl8j2etltPPE2Bw0HZl4i/g0qnfPc1Ta
Jysz/H0oJ7NcunSskIIGdTAqmBzfhCqPcr6Fjizsydu8yqzJaNFmn9Av6SnNHIg5
OB79CZTozTkL5MNy+xoRy0VctPEqoJtl++rZMdzF5lN1xZTxf88qyiQ8pi+Ycuq/
kVcQdFrjUufjl2bzUpHxC1XaxoqQY/Mzh7ANNiBjHR/IdfOTxoM0ZbAb+546M/R3
lHDrOGb0jx9GXDpZcjEYyxDnvJhLkiF8fW2kfWalhA/WzqgkLr9Wb5v9Rb1CG055
DpnyIoIuvqSYgLOumjsBGH3ClhzqMTCKU48k4hgZzgfscsAuW0RQPjREq/BivAff
gx/WhD6qTwQu6jCNeP8uLM+83Axw/1nQvPIlLhc3+elD95OpYRClkQjio6rJmsF4
gV6UzrF1PEmAwwpMcygQoWixlXyEgsbG+SuntdOa3ujEMUTax5MW7szV2DMl1Wql
927v9Xzzve/bXfjRKL/pxcvbNG2PCZvNCZEbYAZXoxxU8q5w85gTUje9bIl8eSf8
kZhuSE9TQLEiLtsHAUAWswBaSTaZgbY3SyDskNA1Iy/H6vQWF3ZEpyyJPzbUsb6L
xrNfAfjIqx3259JU87c1wZSqTLupbTbG3WkXpJq2TQolgOS+EHgE2n/UtVLkW+zL
deUWRbdwwuyLhe8Wjij5luSQuJ5euhDTJPZM0GLk+djvHp5tLpn9olOxbKD7NIlv
0SskMto9M4BQVGPlvMVdK+CG3sPAhGq+tu6V/DfbMfnHS3xeEOxItk7WIFgaDaIR
tmlHpLvdtskQuazspqwMB864uUD9bpfstQAD9Q9lr3sZRBdGbcnhAm4CYu+oFmVZ
wWsFjLfY2zkPVrgmPrW4Nw==
`protect END_PROTECTED
