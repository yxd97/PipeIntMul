`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6BMzDG0U6OdLOZnsjB1RCMFBDgjoKVTYUeAREP155zqztoICTN47oguG6YX3JqOs
1rAmeZjw5Fl2XaMveHv93uPv1C3ZTD8/G1Z2c0YyDDNhNQcWalpatbOFiFhO+UbF
AKx2qL1qQ+fyxo4YpuKi5lQpjzbKRVA1vSBmvsMVDbthusz5z8agX8GNetvBypiO
RB9IhSl2z0MRnC8GO5b5WTbJwZjF4wtZbmjV3XqnDXkV9JokPHkHrNoDP9oG+y64
fxUn7O6BphsIXR0fjsT4l3+h80msLMIMhyn2elV9i2HozqkChfjpv/H+QIHePHWe
3/eFU7Q71TKsJSp0uCMLSTAvY6j1DhXF6KA2uft5VmuJG9t7qJ3vjxjlAdThVU6C
hwq4d8ObbumpY5OJAjWi9EjUYV+wu6JWcFV/M1ylzUT/L29IRIDAgP3JIc35Mc7v
Ouxg5pQRZK/J0enKEwqDniahZp5Piy9veq9YrVacVDhml07JI7eRk60N1aC10AqW
`protect END_PROTECTED
