`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dk64oky+gtGfGBbgiB2O9u7gf2KI18HO2e4xZMvkdWIxx7Ex8z6dgVJomh1Lr5gb
okwdjKJp6a9f3/cWPpdIxxg6U0CMmZR+6jtolwhL/rb275SnT4UF72r44WYbHPhp
kXjbmYkj8SzcF2LJVbiwiKm2ZX0APfQ3SQD5Sv4RVqu8iPxdjvW1/l1P+CVvUuQo
78CCuCrV3b+byLXk28iR4B2Uf/l7uPmmJH48g391mN0JMuoAB0QXl8PTca1Qdacl
le0s6+W0ppt8eK/XoVWL68ICRnRNn1RkPLJ4v+zZlQoeFncRgA0GdbT1+F67sPE2
DJDLXApB8z5XrB9aQEU5ZLcZErMtws+4rbRyruYTR1Yu4IcJ/Tqf1SArAT/+Xapr
0bekbw273XeTg+DTSV4SWdPuYyJv3yIl/FRw99F9lGLa3GWqbP264KHafZte1PFf
1eSPLi01XO9aWUdz1vmqf6zpk8187C3XgF/mCsmNezy61wwFBZ9Wm575P+wzA+AX
uLpukD0D2lq+51o4TtApxDqZrDxbkzrJfpeaR+YeUxdYbvy5a0NCORm1jfY1hexe
8xpUTKdYBhvXpRgtPQgHifAmAJ7BT26jDQyibizyehRY5kv1LMUIdeuBwtssnlZT
RFIuQEc4NOuFANvjEpPMrOpscU9HVHYSiwgl7xbGEmUh05ijzPdNjzYBZFfkGLaG
HayK6CEZRWurmmtb/2Rk+TZwreOtMJxP/L5k3+rRNTa0wf+pvD4jp+sOFdANjG2N
uQrpt/XmWdx+ka/u+7BolA==
`protect END_PROTECTED
