`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EVjZHUqozHV8Wi3LJhLpABgCx6zr5RDNAwVNgh1qlwlnjnucN1S5olw8NQFE+GU1
ie5ORx8mjdTxYyMrdj+9r3hgiddaZnSl2yp8UGUWFZlad9K1xl4+p3djBlIc3Ck9
40kpkCf6naSjY5JyCmcIf25u2Rm2cqlfXlosuoJfBfmJ9DlLHqqM4UGmv4NAOATE
UI18tgOmZoloQJoJBq2bFeXgw56Vz2AcAllNZHLqJn/ZZN5ViXVEhB1MLEUN3o7z
sMNZzjkjtpdQd8Bxj3tKaCTmCNo6RpEuy8qYq7TuH9ly/MfgP61bRsFURSAd02kd
atfg37DYGoTwDt2xhFHhH/llv/Q312WBft+KwW9C3g76diUhAzPcxJBTDN70Oxfr
cTAuaTiLy2dto/Ty6XWLGrB6UFq0cGeQ30dduIqvwqQ=
`protect END_PROTECTED
