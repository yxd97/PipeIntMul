`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVz91QDsWCZxKxOYAYXh58QUqDvX0gkjY0wgYqXtpnlCYvnWnfVzlN0e8H4dyE3/
WLarUCi6F6wA3UaE0bVeCTb2PFL6u2LaAGYB7rD3eJmWWlr/Hn1b68lrhUGx3qSb
kciRLctZPqm862SwcLvp/YPrTViNp1JRiRGltkkwebcOTB7agwynN4nRfPuHyKLH
grJnrFcAsmC/bq9Zpq38M7v6HlTDk2XGPVLuBZN9wy3PARufuIqhZLHU+Ged9QVR
+aFYMTcS6R31U1Px3SOrK4JUX8GEOL8ObH+3VtzRslBiVLYxrhu7OnvR5hps0LZE
jBUA5q2+5XAxZRfgCQlFu574haKtiltCnvohB32ve+6h4tq1VZ/WJZM09UjGHRw+
mPExh1uOgf0eMz1UzSoManGHC6Mhgac2tzmyOyz+6XtVZ85b6YiFjqih1xvnaNNR
cP1Q04Xjt+NgxG/FsWGJqbkjgYK68UCW2g2BomPhnlU=
`protect END_PROTECTED
