`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T25HH/PrcWQvZIZlucLhjhPpUrYJxbWoMoUNGtd8ZG8+zqgTrIOBynQAXafpPjMf
GSTNpbQbJPVLWR0ZcOPpn0VPfI4b/TEb3XTOe0Co1AKxy0XbB50wGETyDuSV3iIY
Mcmwbk2Ax4q29hjrLYg7oD1zSPlGmHcir2EJZ/+LHiGo4tRkCC8vrP6NEJwD/9zL
7alesh8Pqc9/EHbUBqmaZHPefiWSl7D0mZWgbpuI75oy5W8oSydStXHQen3+jvzT
pjXgGLmQmhaB3MaMmTRzh9upMosZwy0pSMpHX0S46slovxk5bZYRuvzEnHyv5V5D
`protect END_PROTECTED
