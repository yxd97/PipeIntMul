`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/uFz32+gDjHVdYY/N8P8rCGs02u/++syPwaPY/a3XtWlnafG6wt7kfGDQjmuIOM
5SPM4uE9mABT9hN44tS+aKOGd6/+kLqePAHJ8DXNYjNdW4odMdEryEgOD9NfDZ1L
xWp+563Zvq/N+TiSXfMNfOWxGRTKIJUGRrJBdGpiwSwGFRIXFq3r2ze6mP36ShGA
hErBiEt/BvCgxiE7qV3wq+1YqNRdGcdL5JMOihgNQZzor1H8Vhl9gxMZgetitICm
zK7r+dFUUNzqD714ObNam/OS9M/cgJdLiYqGjMTegEweWGq48AP8wvAYASz3FFxj
4Lccq9YlqvLQIdyv63EeVD+ATnp+xY1+We4eyuAV0Cy+HxHKaXKyoNhsz1nUsjnw
owkqpHXhpTygHRVFeMoXuITduOAeeCw8W+HSFF9D6da9mxjFoqULGZ8q5KzF03Sx
dY70KqynM72CNvOYF8dzn4pBOiEKjqPyT8Ar4eQUFJmAX1sYNiHj1bVeUhC9u2Ub
RlsvGHD+33MC/HCRjqY8jbdT0R/+PL/v9MWRax2Kbd7pkPvVn90qlkMAal0srO09
lyywL00rYK9Ch/8j1rMRnBMYryE3pjM4t8dgNE9EvD6mPkogc57VmtTsp0tKa7SW
jPLZ/RAyGEas6REEl1QkIEyobmyDIjVMuQl9y/+5APyTm+fQ60E+RA6wQrr2q621
vdzSA1DCBZTYxCBh/bqtuP/vlGRhEydZdze74KhRjTAofjCm5CqqqkfcG1FroYak
wKcwEgcd+JN+J5MaCCv3+CYNr4dBVdUKtlVKn0mPd4Ux9vonsUTVmex/w8nSte8o
L/PiQsZZz2T5HX21PxOs4R8jNKSSsPg4mwHFLABJDOujvt4IDbJRWEkKgTwD7inA
Ay3jzls1x4crho6+M5DUn+W3pghMfHeUBW7S0hmrJGhhmdwmgC3Fqs/9dtbgIayB
7eoIcMUxSxzLg1K3nCWzWyvDJS4KCLRruEaHQOFUloXXhx+1Vk0MDXv0Ki96Xrmu
zNWESKjVPtUwqzT50sE++XB+0x/fl/ccaNFq3uYVa1DljeZXmv3TJ0sE5AyDr1tO
PP8vmdnPY5eoaFgD1mmO1ZaCterm9iAgxMr7zMy4O8oYRc8VZlQOYeO2qGXxEmSm
4Pr+sIsRPxF+aSp2ZK9LYKUfruat2V/E3SwOesP35CFQAlJrUxGUcXE1AAvFLlvp
wr6xzoSpGiKQLmnpmE/buR4kezTqCRFvtz/w1zeYkbDMdaOQK+V8eOsBugSWg6wV
TMsuW4HF10itME0Q+P5vv0Ei27gpq7qFYiRzqPMGE0W+AZWbMLWV1gDOKyqxuFbf
pQYBNvZStScv65RDSz8FGH95W6GBRzegFsh2eHg0OsH/JP+tfEE1v0mdJ+Sd5xgp
P28q2ECrW2L8BKp4aqb6KK9wNEs6BO+wa5DxBHlB+cykz5zoPAGugfWJgSPH9Kj2
9p26YxR0UFjMMjANg5SHMUtBtM8LxCA/hrIphvpxUWB/9SZNMJf0yfrNxdEKdKyP
GFeNmHt0X9re2DcZCdlY/A3fcPEr5QWevxink53N/1U=
`protect END_PROTECTED
