`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFfbKjJOzzQ6YAYdIh8K9gvlyj7D6RfErCN90oPSNXUTjyWNIHGgYOVuwmH0Ixvu
AdE7LcHZtoPOT1SdNDp3prLqtM8U3RrkXIeJCLNrO2nRDmgNsWLsbK8ebvpZp4s8
+P0fnijChmr+3hC1WqeOMkEgcILiok29jqF7fommdQuuN63vOv5sPe48v9NVIRcm
Ak6Urc22UdfKF2ZxrUAL7tDdWfj0RQkMtG7jF+4KNNiIIG6x9IjM26SCHZjjdSSS
rGlxJdN88kiD6EfAprUDt6a4XjQXv5QmfCFpiDTDXDeGwz/c8spZYcyY5JF83y9g
Ct8p5w78nS65fVMkOcFR6skMbTYDgZy6DRsYaoiLQ3sW+mdbTaaXtJdEV+oPzRdd
/DzZw5WiaZSPuIiljXjjopagy0hThgzfTSO3VwyZIZQzpqAvJDxPsXPUxkC6j9w2
cc6skxxKm4UMDGxyTGOMLF/nNupBAx6qfehQIZn2LEA=
`protect END_PROTECTED
