`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fn8LPVaaclCPXilsAYAAp7yOxkAnYNa8zpSaL7PGF6VMkxMxlNE1OPjZA6o3gvNt
oEQGvslcxmVYPNTDpdRzkrGuWiAEVxA9fihb3LkEkjs0ws5REol5GvDg60LA0kPF
8O1G1RmSGlpZfM5d4Q7+WvAUW5DIk34VQq8vbO9fMyqKk0ZTryX2oyn8z5OB2Iou
W+mHWa0cXSrKfdOGnMmE1PzAZqa253DupB7NOzw3JnDL16UI9nB+iQEIDlESaA0i
VqiqqNrXj6rlBBWlI2BsixMmAEywIESzd4QiyYEK0BTkzGG1dk24gZw+gO3biOlp
/okfJPAmjNBG1+Qa/rSIUXIbfdUck+6wxcrZMzqEQZcw1jSrOES+x3QUj5eG5vd8
FIRvGUXHbf+hpfZZsrFa4/971rLrZFZqVVrKPyCCz3YHNyrPXdSa6pN1DNj2gRAs
ZAA8ImmSIYu9rDDrTqWGhgYw4b1oqf3CrlFDwfkYOYvJp0X4rgGQCzecCstJeeDN
JLqppKXzKfegVBZZD4MBP/kvQO2tdBfiDcDiCUKEXumJvQ0SUodOLYmIltb1Q0gu
iTTJjaQwnHhz45T47icGLUegHhzO7FBRUYuvwQpW+yNBc4S4Lkm20v3y0n2b+vnm
bYlovMOXVYCTDnnxkNjvkQNp+74SXi4sir/PViuWL7TMGWjeEOqZnijN+4I2dOaH
DUl8fAWVsOJnz/uIwabT92sY8Kl+IJ/wbQ7xeePnxAx5qEISULb1O2+EEiNAgRt3
UEk1LCmtAhMnV1/KNLH5/gsNWxbcMcTVMS3djr3eYXFbSCTMjv++X088vYbhQHkS
xAGZRnmmvS8aHXUjDLtIJa7rYs/kElZE3rIqgnAR2Jm5JZ3lEYylPTHz8YdQF2gl
aY6KQkywAfrimqH4+pd/VvLSxCgVlpMhoEhR2HnKQ8Jiy68p+Gc/xx+K+MVJEHJ1
AfEUR94ox54yCCsfiDTl3LaBI5izpmXzY7KtsR4vgqmwW6eFhIRhYQ4AITtjMa3h
fj+pRrR2z/mzB85F7lsAH0K2KjxbREjvMQ61ddzX4TVSggFtdXHup7zmIgHBPnAd
eZFfMHiUX90ig9+D9D8gti0ZQbE7gnoAZCMqVKUZqhcFU/zzCEkBbrApyP75fu3t
iUQctqAkW2kQjvEb0nGBSTBSOXsIBxyvIzn+4ut4lXg38Hw42fvpe6ZwD4+IxWYR
edgWq/e4gLZgPqV0CK2z7gLEuZ16+BDCV8q53JAZXhnW5uDUl8e5Fmv9jhHaqc51
7mBYbOPbL9Hfj5BAAhglPx2b8El0mddrP5ZNdoMEllOm3xNFfKiRmwzd+uBXZoQh
bHi8BUvweQXU/qFZng7I5b6dSBSy4GmEYVzbku3IjyP9ftyecWE+Et+AAtPFLSaK
LYS1prz1KdCvtBZnB58Hydp36gWtbop626fZpWjkT4awqJ8P5XAAM8/8A9RRcKex
z4VRXFRF0d17vsaLhecWFDhQRI1dTUwMFeTt37nP3wV8U2eBrLnbi1x3pPcsCyLr
ujn5mHP4253zTK4ipJsdEszclLnFWwp272VKgMYw3HlKOpLtkU2G4wI/E0fEJHpf
lUmdO/VnGN4MG+3xMIYMTFqPliuBOkg1rfwM24sR4WWBHsjP1tGwjMpeUkFth339
WsoDeSbHHoi1PvLp/zQWuZF7V/avXXhX5GrTVKvMji2pZU9ioUfojpIsQBriM9jv
mBn6ArHHSDyOXX3EbxwYF8sP9ZcXem23kR404MSzYBwNU1tn9U3BtLsMB47kU62/
LLnvMUbedW/lSzv+lQEd/XEJZSVjNwHun8mR2PF++dPA/JlvOW60SIsRbcPPmyNj
ooaXLKInQYxy0+Gj95KqI6KclBJZhBp8XmApKnO7Ts0FA/XYltuj14b2zQ7epf7X
Jga8F6kQztke0L8tVDmvnuG33W2x1cX7oKgFEf8FFzFxO/zkJKtHshdGTSjh33bL
2iwvzw+QfaijyREMxRMov19cUa3tJvHLW3iOGJ4PFBEH8hCArT3YxOzMJb1um5oq
P/AFkWUX3f8LywpoP4afRCSFkQiAPqUnRzmK27HSoRVVvSqMwSs9FMPRI1+WetiO
DH4uZNxWE8gkoiZkXVQxD4xnkd5SgbLHiukSkz21eTxAhTBSIsf/TO1F9XQuizQC
0Lh5gxZzqKxdtBIbmV8OqhGo6/HhqUzDMRn8e2LXJakUtVswfre1lhZUrFdA3tWe
oqxQZQn1ZtqsUUHVm/PRuBz5+W6pIYiDgedbd+0qMAZvgPkVsCH7oS1BwFLtZ9Nb
yoyCs3mEC1CoFtrfyDFJ+a7gBVc7Npdw2uiDVFTUaTjad/a1m9z/MqnmfgEjKs/8
VSOd59YS6kwrbG9dJLQD0WvCtYSs9qORNb3pT9fvdoqD7G1V4ixaZaQfyDf+LRQ7
2dMSFy/qmP/Ar0QGYrKK8gQrfJMeEa+4OjbbyvAVEEvndgZ/mvlA4bqhIapGTvJw
Bx9m50Dfi7GW1NRm3XYN/z4USfBayX9NtINTccWbhbwxdm5s7Hk4Y4uT5gAK5NAT
gFNhcnCKJPHmIpHtCOAoLqHSlv40ej5447qpK2EvqfWIiBW23S1OMwteMkvJoJlU
ze/MvdEWkWwnAeqsyLLa813oCquAk48EVvIL6+w5N9py92mQdacNH3A+5eP6t8NT
Y2jWt7rKMsT6qZ64JSdpQAtuKCbgIIllzp2Trqnn3zuEZV4OkO4lWRYy/O4zC4nr
Mnvu9qBtuHg04Qt3zu8bLz5wqudRVtza3uCVdn0/8oGxi09d3Xg+74/rLBqQHKN6
RXH2PZknbU8Um07rAFpraU6Gj+K58CHUJHnC08j0Suu+JhMDRg8WgGNBXMqUKPSn
rIX7kRDddnPCPdf8s3f8khNEdg1QevLgp01YYISXlNUxLcSy7ucVs8ti/yBK3LHf
7QaOboITHS6YZPUeJ5sRN8tYDkV53MQX8HfP2gNsg9LXSgnxrveIha+aLZrlaHYR
kg4bJ/cgzYxSXNBsbJ+Qo7H7XmLCSMNGbuRsZwvlMfMpOABOflO5EAgRA125f/g2
d6Qv/PlCEx3IW3T/IL4zYtIpSRaXZ6FqrAZoMUIdNu9pYQkDMfCPlC/EyH1Bf07W
aIPOR9rOz/xxLBDriCLEBbe1X3yfKG4HgVRvjS6K4UgHmbBIViIsAe+xV/LGXbvO
SONjKdO+X3wfm5Yt3OBAPcpwW9oRtM9MLlecpbj7MlrmpPJVU7ruIrATLjlLTEjE
t0nxphyFi45yi6OkL1P/ZGtx2qh9FlGZ9QbNjZUC24DCMsCz18r3zFam7Px9lktz
a5G6VKpZVnvM7utY2l5WJ6YzZQ9woDZ44jN7h5eW4Zb2/qqKdQjbBewDhwsSQ5fN
6T4mk+EsP/DP4FyAx9EAUfpD41vke3DMXzBDdgeCB03w8OSAIGL8wPBgHKRVm5Oj
W4HxPdaw1Y4Jb3DfeF9i82T1+ER/ECDmoc7thyqtpoTLUPc9ghWIx83XsP/JtcCT
Ph+6kqCaYhRGt88zAOPo6MP5328x+ukRHCVmvu1GpMt/v1xsbi26eUKJn3JqUQm/
RF0B2NaLgtf4mhu03zf4ictS+wNsHqVeMjGT1xHe58DRXWohsVw/nY/TLqRruET/
Q2+jT9XeG9ra+hAKSqJ3HZ3+FGxj0hZzwBBgJaFHLTNdjgq2dHy4cX+tq2fmoGk1
JXQvzl+7RqYN5HmKnmHyrxJ06vi+5n3lm5e2rRMEosjGJDa1HJkerIpRsvk4Zo4B
7NB2/2QqPEG62iqL84/fVtbB3IhLfiCbS7TLnnE3o8oTi0qViJiiW4hzx6GdhuFG
JZHQFEzQHnKWtL5pgwQ+n7v2/Zl6YfHM9Q2Sn+LkPWBlF9r/JPNGB33m7U3dYduO
Da1tDTzmGqcTanVD87V9HiEcQmxFS/nZesXCNt9Us9W3tT/9Df0gLCLR5oA42IDy
PpkJy740SfsA/0qRsRL6hgjDP0PFVgAoCSybkQU4UJDKi0dmG3PbANz+kMnHcABD
rW0VSHFtkx2TV5II4qIgazcBGlZaiTQmi4851sU2O0d/ItvdMkST13wr7mk3zS1L
rXF/wfpHr3Sm9nPh3PSb4vsSa+OBuxoMDFqQ4hD+SrN8f0MdEMPiSFwrJnC3GsU7
8JUqX4C8OTzp8dgzp6/hFN1kDK8SMdzdODOSf9YSTysl25+VdaqDh27VbAJG+Me0
nCHP1In+s3uxb2fPUaZr9z3QPYJ+4de6VeDIhJ6tEzlZaEAuBREEcAbrOTvL+3UI
GEYUTPVQ8GLdDjuezPNU1x2lGEftHAmp3S/YrmUV2PqANPMIAY+vlufRyE94ZFXd
84khlPTcnxS2ek2Ky2w4CTOykK6AdfrpE2rOeHnvtflzQrshoIqbMnju7lRl9S+r
BbhhWnVnR4qtVb8yTqyMSuQjjZPR2s4howaQf7hdo3Y26XqLuwfwpVYwIN2DX/x6
VG9LoOwYOvnh7Ip6Ky+tETiazAZ0B1L8F+zPFK2rqwrlB9tWMHMUWQ+i5KrtNr+X
cnM8GxbP6Y0q/36j8LIjHih+9t8Z2UicxXSRAiv1JRmgu38wl1TTc6cEmtuxkqMb
lc0APNbIMc5NeLF1yeclGWoUOI45CFOZxDvZFTLE/v9dICcUEmIyInmWudmY/w1l
TdXL/5gwAOtNC+DzTH96s8sPbDE7liHIYgzMB/1kZSLDihmt2vX6qPgzRKJCWfDd
/diS0x9mVApDyjVFH/iRut39DY9fr+GiP/z+Hcy4TconL+6E5WXz5Aomf5tbNg5+
JKJbRWuXiVDROWyUmAXCWv7MYxHrTPOdtM2FblKIHaEWolyKTLTnCg83dbQFdGQC
LWponllaXKKIUoTrvh5Q2IuC6cd5MpdH66PFoCPCj72nn0i1f3k6jvebaxbKfYP3
i976T8SruwXW3uTa1thrBHrX3ra4vjQ1osvEbW2atzd2xnIp3LXFD4stUOQjZMiX
OUxN0LHdI0V/0it77OxSnGMJKUGN6oLpRbWsWqIyPhaDqpjzFFdIeSUqoRgq1ulY
e9ROsX69GikpxPxlMkFjpMcxIBrn4WI0FB2+iurMTcsGpkF8CL8mkx6R1TP5JHXc
et7+PRNXgJiraHaOp9Z75J4UlE5ZfPz9q3NZQ6OGeG0NkWlriO4LGHb4fZ5GSPsG
D6tPd4+A5PHUagjgavxXYsypRu1r6JDxe3ioSzcFTvcW5r1W8sXWAnncKD13CZkJ
YXn3wvgu6tRg3J35PTX3Wf+8BNDsNOaiT+s2vyi45lS5vAW81nGNkkHj1hkWeIf+
PP03bO0HgHsxuhXWzfktIHOYkJi1L3QB3eOhtS0iTCmrJGr1y0AE+bQivdnYnhrJ
S5REdqQDVIqxlIYF8MgMGoqUUJNXLzbkhfjhKgX/qvGnAg0hahBPjj7yieAgSzca
Oy0xFoXIRl0xljgZUPX+zcgEcydhFdhCrQw47cFfyfZsJUVmulwDGHnwsajwdkzV
jNqqMl6/wdh0qzrmBj0KPJqqQDqd18y8ba9uWW5ykZbH1Umqkt1Sf/eGuelZK6p8
MrmGLm350rhd74AW3BErN38XGl082p4BNBXlrzjBAYv47f1pzrC37fTi0RKX/2W/
kCQZDL+fiC5xOgnaRwbXPiC1oSHbC193lp4KO5RxwQHUgVxNOBRsqjABtRxXw+bh
MRAO2WAJqjIZTcbUBvJUV7TWCIzE0E5kL8t7Q63tBloSKxLVCn8BXv+P3hgGDIN+
TQsRN2z1DrFFeYS7RQUd6O2kdVF85lBdPX6YPPdUOUpb/6mexoCfkQV+S182AAgk
qt3TWI6QDS+8EGB4u3Z3j8cyU+r033SAOKMcZwQmQjuSbZW4tMbM/5kkSwmN4L7m
d3q9xhiP3TuFBCJQKfMAt+e0FypvzOsc+4v/8oyBAk9bZ5mqfT3q3VpaMVS8p4AQ
e44p51CwGInAq4N4QiK/a+YA9+jMZsTmh819SQJxwaf6IWagZOgqG2FqqfGA4VWn
zcIMUo1q/OB2mpgKmf3McdfS6hkMXHnvHrk3Gro7R1dOfmMg61WLbKXTAw4b5GB/
CiYJobQemp8VJeBpQx2vHTJ8SHlQWawKDblCAgoIXG01agPWdtV43o40h//WKKyx
SSObUyNjuAYcgyfV4NC2subGpvcNF1GCmEM4GkZAnDHlLQr4s2yZFWZelDeN47Un
Ww6rQf693vRzxaXkPEVnLImvWxYL+VlrTXEoIZh6/zNsiyRgqX4D6vDFRoUD/1D6
EFAW1F1r8lrTqThY2CR5oOtHmBnSOr4pjH87C5cmZVynm08Wb22Fgp0w4uRoYLGO
ESiu53Ngtna+SAsRpbKeGUGNbUFAOjR16Nc3h8OtOXN3anbK3Up00ntgjoJzoeff
31spb5TMuUEFzxShQmB4X1PzlHPGDIXMEneNjQVICNqnbkGE34qZ4opvkcypDywg
vBpz+Y1X0o6CrW4cjajOolQinaCvsfM5GRvSxfhhDvC4HRf/sgSTCjXzgINuaxZu
K8TiZtaE0HhDKhVAjOw0pA/whj4OYblTBZDI9Epjr/+VM9+TCdUsep3ERxGmraxw
gQt3ccS4XsScSUr9OfB7DmPOK+Rn31QUk7ZbvPwOGhZwOK2XW7ifXhQGsg9VJkd9
sVDXTSojuppZy6l5j/L5kewhu3/TNZa8g1TWrmSzA/qrdPiSm/4tOP/x9Unn/+Bn
0HHbQ0bu5j0XmTGxZNBEkqjXUXZTZW8mVwZuti+vgDH5ZwyA52qyPAGHu+QG8oLs
eH7PjjRERdUU2KY37EcfnXe/HPmLIMFx2V+HXymlHz0Ym5MJsM5TJ63g+v1Vmxqh
0QMUD244wcl53WXjSyw2fi0z+irXGp0m7i9wIJJSlnClZIDsQ1timQc0ba6ZSVUy
rbmrfccca+EdKpZdeGnE5KVKwly9bBitCamgf8NadUurn5Xvzv/znPn7e3fCIyWz
8Cyr9I3K6o9OlHPyAR8HD4j4e4GSBZKS7Xv+mP+jesbLEV/w9+lifRBdhZvPdUPo
T/pCwh4/9tzZLKhaMmL811a7uO/jrGwifjSYrjCC6ThRnXyMqAIT9ZI3W510T0Oe
mlCpa2f3SbqWQmMk1jo/MIzYR+L+C6B9R6wcPA6ACPLx7Ble3bW6ay63n6PaI3ki
3ksJzQPIphgDr7ziGBjlsS29J/Vc2d6aLlk5NIRPrJ4uva9KNotKomS8Ftcm8fUa
lD60umF6iy8+IKjzbkyJerRgE+CPO9mWi6fxcKePTPm8MFqlZR8P48QUOmRhyp9X
9vfsu+wk8PL2F4UYALo2JWCtx56jz8gNiLMWHc1DlTqJYYxRWvqf1BrqZUa/CDY+
kPTvJnAWKRWnTylffx0ZCahul+wHNlPn36PjKMpUNrvsrLg/UrVlBzRgOPcwB4lC
1h+lEzkOykoo2KdHenupZdbqSWJc7Md+6qDTRGDiM4YVZIYDKXmfd+YhXa6YiNzT
MUCKw8QOaan1ROOzdnQc1IBcN7oWPIlVf8imc/oi9joeLo4RSGP/YB3YTskHpfJE
5Za5vGpCHBBpJoeTATMoFn5bQfu/HEZFkUMWp7n3EQo7hguW7DmMv3JRaTN/yPrA
h0yf4WkuuKmhWdDJyzNq0nTVfax/iZSVJl1EpKR+pkrjc8yKnmXtRiV3K6E6q8gy
1nWqS8bx6da3tB/2T3MpRdW5L4vsXKI5e+WSiRI843TcymJbWj+mN5AJTrduuegi
1NREIVhOnAXnmHF7VehhJxEYSgZ0JEgWiovsq51spCg3oNG3ueuvFGbHAXR7HpQH
nsnaJqRqPkXrX8xBcMfRNPwhzpZZz7vhlDjQav3fJZGfeYJ0Gb9p76FKGsLpZu/F
DKQyYJgpLTDsnre+G0t7pymRVldrWB2DXesqJPj3YhkwrxxxK+NGQkPLhOlxA0LY
jXbFI/I/h8U2nu+uzBem+w==
`protect END_PROTECTED
