`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrTyhkPkE+R63BqdQZ2/42iD3YSy2L9GTgAtoyiwn1yMnS4iIMcstix5207sqBtt
1yO6x4zr86UsRX2Q786PO4LNijYYMZ8y7/8YGghZEkNnBIxbbKfNyXdbGeXdMQ3l
Gqbzi1OCrqFfYaUWxmEzJXPs5Xmv3zMLYSTkvkuGcOl5awHR25py5r+Zeyvsswyd
SiTbfp1tLUduKh9KHFUY0xChLG0k54AYuwMeZsyXAXsdkaeEa58UPmyp8/zaBrvn
vtEuDWZvOn2gBFbD3jjaFOI4goz/YInf8N2pKgQzZRvWt4j2s+av0Dfhx5gqg+Ng
yDJU7w6vs4vcg1yoyhfg630/Ccs5eNpk2MBVq2YyGmhd1cwIu/k2sQTBsWbbu13W
0w2ICuq3jRobi/c3UB8EJzY+6/9Dbw6D3HJPWZ7lP0mOmzaU4BvAWzzIHkPl4iJU
VzsRMhYMgfHDVzdZFOjQrvVMWVTqXfTenGLPk+6r22t8oQvqtfIdxFrlBmZ9ghWl
TtgCUMw6M9PrXgfEacDyviDZjnH8rtc3xeKBMtY1D/MTeN6CY6f+yGB/4dX9mKA6
AvzbGamL8TtodM+Saq16t78+xigShrDd0Xt8zOXORY6oujO2MEIFylUWOOQBuBgr
mQBdzrb5FuExyL26PydVRAuaGKefpttWwDBk/fVDCxOwBy/EYcEGGaSjCgjRBZOm
Zp437X3hRuZ1D7dUopprWtxqX0KGxhKSHndjmYvaAqyw781axgJvXPWI1n4nOQhQ
p3kekV8avtLsji1m+eD57H+Dhbt2T+J40nFLDCUCJQYxWmNJjyfXCEgvrzgCQHGx
O2PlU5y7Lja7eYLLEfMBE4SBHurCWnRk84HG5X8I44WfMx9/lWYA3HRpt0TTZoU5
KFxHbcsw3XEILVzUW3ko2x8osvvKOLxW7dmaOZqc3+1bcdojTUE6DfL0hsThcslk
6iG/ruHJMD3nQ7FnCCzuiPhsUtBGBnhIDPcpLdGiLNhoDdO3dqmkAKztKbVY3L+T
VvGtf88CEblJqywbl9zQgYzZPUl2/riiVPhpUt3u64lvImjpLH9imDhnULxlUPfw
E3zaMnxDLe+unlFQbgIxnq37IRrYOoXDj5/ERWAYOmmMTi7cLHLQrCaUv4gRBzDO
KcPjSyETg2D2nHLA26Dx8gSiCgwpdBKnql87dVJLM9Ko8gA3pt5wkujqdgcwVVW5
ybEDiFCI9girf1vVwytj4pSjgkPnfuzq6fRRvmJzTqUvJ18wX5YAf8P11AxQ95Je
+bqK7K9+Ssa0EC4ZIkYTzvrsl+Wr63bXg8Y7Z61JjosWmayHdS2PN4siSYIkgtF7
6dPItV0CfMV7ngsSNeR2tmlMOMCF6Cnh0JTxkqx8GEa5/nJGPThEcc5CKrsDrdx9
2x5veHW0aM9GQKvE7vPYKxtq9rnr8nSthVnFBmIFbXcNmQTii46Gu58B5Ts+q9HY
qimCovw9QRylZqGwjZ0WIb901mix34olaJw3YF7csL8HPELawPbiN7USCxvHnlXo
dWig5p9y+oOv8Ys5YkuuapRKvZTkis8Xd6YHqtlElDT91gVuwYUqkQPnSXbfrWUR
6ll1CqHlLUra2hITNcs6M/LD2JgAjoOLWOhC2yN+6nSLuZ16pQrtypkcoXuyhztO
vwSib8CTZkGTXNBgYI1ylMz+IdT07GA52l47VhXqDOF8VNB9VYmz5l3vAna7cSYT
O4X+3xmom4iFe6b49P6EpDjMo0U3Cf3Z6jWsOi5m0YkY5rfyMflRpGig8gBuPnRQ
W3ljGoFIpmukXI3QPxYXS9XU6fhVzlAeRMQYdsMmWMkWtaU8FYDv7td58A2FaRBx
q/N9FGzc7CnRdrs1queGJBS5kdj62fArEA85Li2nr+ZyJXRHmlT4+Am9fShBX6Dy
APdamJ5UtiaxAHBh9MSggVuZTzH90IUwUkIRdHIOb3yzaRXnpHQDtkGQ11fXvRxj
Vllp25fRhyx32i7S+YNwbgrb7+JmxJ5WOUZ+HAFVlUfCU4cMHEL+A782SBaBx38U
qeNU2cmnlUW0MgsE88tUfrvcITL3pIc2ryZoEwK6gAZFtQwKqH7zNyi2HaYRzPGa
PLR6aF48eWA/XBcYGKISvyoh3crAavnt13EZ5O1mlWHFx17CGUvym+diRZ1qUkJe
2R+kMGnQT96mSE2fAVxCSMGQ3apk9cDg7DlNK89ruh+aiwxNjT2b0Vs3km0ZJ64o
4D+O9OdxdsMfv66PgdrXx3VD6lC66Umz2e4SoxrxkMKgQJ+Y1+i+VfEd3bp0F8oy
md5DIcfL/nQA5up4kmhfs6ytXz0sp9xVrQZQptbNvzNbYawaiV5YzxKXEaj7SIxu
DsWsJcbRFJ7BZaR1xR2xIC8mwlau0Vuz9+gY4UX29bxa/kDZkTjBj0itl8S1EPJK
Mt9ircDWU/I/plLRZQK/JtV/Nod6Iybg7/TEreInJU7bdPKA+F1N6l0JlP+QGsO/
L7z/70c2NOek2BGJx6sNgJjewI/lrSovNc3GFZBH6GwaeAUCazS6GZLVNq/Uvfqp
GCRRFrTAkz7nVlmWkOrVc5OZF2fAkVkn2E41Yl25pUsvj0OWAosUCcf5V6KXty4R
hF9uMQVRe416vKctLLkeRljcvTQHklkRy5eB10VOshOoXnFMz1YXXblkXhvhKA3M
7b9EMZWRBY4eAhkg5kcAQXaGXAOPoh1dNFw8K9o7PpA1+Ga0vyVCI/vvq1WzTKar
ADi/5HjGv00AQTc0CjaO3JcPjsWl7wOLKOmo5KTqhwWqpwSG2lE6mc+/Z+6VMy8l
kS9tZ16SWKPgjRJMMMBWObQWvNRgwIq0ZKqY4sxbx4ZKK9ho6h18p3yO1FDIP9cz
UMClLuuUUVT+iaMxKxcBBqKw3DZ/sufQFbB1+xIR48mF+ragA/v3iwsQ3ZcbVfR8
Si8X+de/pQAULgroAxSMsdmOOE09MWahdlbXxlbsbYKNAsReHa+9SpKe5GeVJPgY
m/LWcqdmppvqrtiKLttUvw3jY/zZtGuU6wwvll+M6DUJvA8MQuz274F4vjFHjfVz
DrrKJSZSMAgHYmq2u/e6PSKMAC7KTONzVIPDVZbDLA96lGEe76zYPs6dCuqP5sc/
v06W1UvN/sANAOYESxsXAyhPiEHvZsWFEA78H87DT1i+dGHUmG0uafZ0Bl/GEgb4
Bv6KI8sv8oH07Y9xVVIl9T/LlR75hjctN1Qdq9PRlGUaY59K4UZ/1663H4ined+c
eY/oWXLp8hhoWewiI3omXmteyDu/DwsbdFAuOCCmoOg/NRRdp52XOjAGsOGalUN8
0oIWAJUKbLs0MXzZYRcRqzWpWMYy36XeelEGEd+314U9mNWF7g1Oqj4841rqMGYy
wLklAM6ZpVmwoCGDPQ2K0BiKmalYtAGKlVN3nAtlSoA=
`protect END_PROTECTED
