`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBrvBviBurF9BGkkki0mMD1Sa7oijHlTY5cUoOjt3IXEjGOyX9+B9+JinOuwp2NN
Ct5md84a1bZOIzYznQO3T7a+cyGQxG/ZPK1L3CzFJ/pf0h+ycc9p8AXUWufaKbyK
Rpzu2ustE2fhLmpCxjdlYcbmowMADSOaPIUYf79vmb9my80OzgfKpm7RiamVEgir
l7h7rmZ1c7a5GkPrr125im1wlNKIZr3/OfxcmBshXkqTJxMMON+Fk1tRvNmG1OC4
TeuqrvLId1p0c40OZ8MShgIIxw05xZx1qzRAFzg/c888nBZtC1tKxi24+B3zfvwU
AX/ZwoNi7VcCvUD7R9wt0ciS8s2uBZ59yH0Tds+xUmObkp3yjql830D8YEXr5u6D
it2NaOh4AcwfYVthjcXB/Q3Cgi+7T5BCxwEI4uvKe07/4beDQdxr2a0e+KsEBtxE
asvJwS1HNkSdJM3lL6G5CUbu3TQf0KpobWyxg1k7vm8=
`protect END_PROTECTED
