`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8uhp64AAXMwS7qtpm6tvihXcNpPyWzkfdiy0eZ7MUV9uTJAh1j7HutLITXDGynx0
eEWV0sg0HGi9OURJamdE9muWsNOulFmSeMTFhwq8KstzrmTkbBcI12af0lmOvvLS
fovSl68qijphA//ar+IhYm0CqYW6dsiH9DFK7NvDynxk7rmqYvI+rJvWf9uR3cq2
kdmDUBI8zV40wCY5YyautbbVbR7cLzNCI/FGwX0pV9zQdue26Bb+a/jKKkWcoBWI
s3/406StZd+D/lVkyfgovIye70KoPp2UwkEsLfYirQAI/YUScIQpxK0VLjhtkeLa
19O2SoKji2eWddB3vJLHJmKKrQrcp3cs7tOKIM/wIw+c+HozljpU/GGLzYUXtXBe
hRi3nCSysIhu/D270UVDMg==
`protect END_PROTECTED
