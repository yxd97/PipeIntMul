`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88iUPsEt5b6zUhaNtj7m/0Vt4W2SseV3Tvtmah1L0ng30ix10ffqjv7wQ4BAYp79
i7XRMOdHDqKNvgsCbifHsplq361TYaW+TOimsCPYSsectAwweECqXDM3Bsfoylxe
e8To/l15vnHf1fNMW7mvklV1GRjs91cIlECJ6QUknutka8o1fl+hvhcJoO/8hbpi
5MFhJpjpohDpsp3LEN3V8wWunX1VoGd1u4G6+j7lnexQejyJOWZnSbVXkJwemTF6
OyOdUiEBkO9CoN3NfEmihlFhDqqjD4nL4HryQvL9+aoBYt2G25dZb9IzVT/1nZdK
AtqqBBZuTM9KFEwNUNrX4GNxklKqHUa+R4FRvzvSfKUicb1gApflN5e719tD/rZr
LZ2uHd1M5jdYx8saVUcl8UiX+9M+3t0/z8q1zM8zcC5wSWeHqSLDZHF4zYE3wCIA
UqeO2ijObykhjIAL3v3UIp74HlUpypUBnpKgAp0MLCOx0TkPbjknd+iSk9syBNfZ
TdjMWpphpTVuS3zRLpwoYO2CXRDNkpCAX328euDKTuUeJi4CgBgG6LXCBGXxFyFL
go57K7atdDFGRYfqfZ3j7o5Ho+XuY/l+6KFUs3S5RNnZPUN3HL2wAdleinrIip0u
J7UbnNyE7ZWnxNb6tH3y4uVTYzj7+XFxD/6Tr2vaUWyWC047KtNkHzeR3tHKeTA0
KNqdoBnio+6qJh0g5O8EkaT92PeVeLNGQAKb32S3X0FuILcSUz1CRokfnuzo8uP1
0NAjO5859ur+vloaQagx2dSPk6aKsUASRGdH8MHPZMr7GzyDXLWq/CbfPRX2/Tem
6L3x39Dzqh0Pa5dlVwveFdyaECArekYE3CjqepqXsCFHb6JT7S4I0VUPdkzj5W3G
1Twp9A1eiKYfCVYwNekC2jBH3uhh8xSYECTG34Ubs5Lkoj4a/fSyRsUsUHdd+awJ
`protect END_PROTECTED
