`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Lb6cKulVRKUi33AKSkzkjn47x6aLTHpLMt6DrEgwRnPvJ2Ed4B0d5qwy4XWjuNy
5azOIc60nyMynItFiipdK+zbHVUlPBH3TgYhz4tCwNTlRYA7/hy1yKwtgugjwxEX
fxED5bfF1Gube29LFQ24B3WUnUBvDAwxdf5iIdLXMLEn9nhanxlcWoUrc8ltvOB4
jXPuhjrHmwcpI1lH1pHnleCqvPdlV7INXfeEOMy2XvgBpOj23Np35fbMGd8eYm4Z
q8SJF/LPYrOyhrdFMqBXMjBPRORLD7Jx3ObbKne4pKN3tYLSWVOmZvWDPUwtatIw
0tnG1yswEqkBIl46rYC6jSkBTcXba0LE9hShwSaeFq8nquzbdjikmXckMvBvMrLv
uu6zt4D4Aec74H+6ZWHwXZVIXRhurKhrpdC/3fkmgsHAtPNC9HCz1zmS/zfiTkpi
`protect END_PROTECTED
