`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s9vQdGmIT1oA7aa/C6njOqn3KU+gxQ4X9Hn+jMNfmNfdCYZswtzaOTkqoFg+eDZZ
s5JURrihRNiJvwg0y4ep6Yin6TTVa01nwlamZMC7m+Y+9XmgPCLA/d5aSBuumsqz
be5s4RkydYeYLod2xKBqm0pNFcGu/zHiycn6sfiNP0xn/WUvp+rbAioaP1rVhGb0
PxYUeMpRQ7q2pACjMFEWP2XTOiDMeVcfH5YJAIWuKM9WfVGUWE0w3W/8Mq4akIRU
WetU+2Y9bcP/Km/2v3VhKatq3tApd71zMjSvaz3yLN3Ryg7yeoeM0NVQvkUMOiyT
qBqU0V6h0Mo40uqRGmnVX22L69WP8zwkaDPuTgzA++95gYzgkFwwbOJfx2M5Ay5i
PS5XxGVgJ87uSVlhZyIilQ==
`protect END_PROTECTED
