`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YoJwgta0uJ4bjXH2tYDgGVTvbUq4ivdvhLDAffRTgTxwk7BMXk89xXqlW2YyWCDg
lh3PV4ntLM6DGfJllOTfwNgRSGrlhN81QnpB+ItFiRYYJIwyzQd4iEkFOFAg7faF
3bwSgbekJqnGfX/oxRlJI1d6BWcwtpXm0RzLAkZ/fGt51x67DyNa2PtmQZDR52FN
oWIJ72nUjkEuLea/mhFgTw36D5lJbd05aQyO1eFh5I4LlVZyqRaFxttfgm73YCRY
oMP4gx2mdZ4IntoSZS2brTQGWIqeSRMp6pdiMRseO2oDLdbJeYKDIaTCxyoiqdvm
OnrgUyBSJROMUWuqEEx9K7f83GW6sCbvhGBX4zChwhV02zBJHPrtYJQ+y2sCuKZP
uoa4jXndlepSWk2ysymFaw==
`protect END_PROTECTED
