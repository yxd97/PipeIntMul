`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXBV3Go/eqRa2Cs8OeYkHLT0FFyOz9D0NqjhKIyn26ywScbDkj9m5XlZJmpfZa/U
cAC6huvRciQ4iGupfbYC9HZPo5+vbjLd4i330ldkHc3mJOkMulSe1N8YAIeJC4Is
DHgguOQgIy5RoBl04UyVqziqeiqzRVZWX6tcWxBGpaML6ex/2A6MKJb90doAbGo8
5PLqsbpXgiyFwHfb6JYJ+CtwUa+hnaeQJHP+XMovJohavNssJgIP4S7nJ/eh18b4
xmRNdj4cbq13xk7Sfr8C+dolqSx5TVzp3NMjIlsLuVolOaip6l73+HtFJejOq71c
eJMaYalxdibIitU7jtCbfDLhDYR3LT+1qnUoO5d7pgjw1rJXxJIpspxvKhYZWvQp
WP1s/7wNFJ5NlF7qEW+DRuqGmpzCUUEl14ceIeldyUSE9ADkO99pgplPTtZdfRNY
voXYySuKNe+bGycilwCDWA45eeNLXkpU4U8YX8j8wFf5+4qwMkZfMJWnBCXxmgW5
Qg5Vy7MI4/XHf8jBleULZ/Q18NJg+xI/2m8EXH1N4qNB0bDSVhBkc9tAc0Bm47t3
/SJMNeBsYzdYMerHRSltXdkNLSwyuTXAzl0zZweLD/W5MkDEMJlzFWZKLPGqG+X5
tSqYzkOmsxbF3XWHyTNEz28lb+Zn2Oek4wKawy+LxrI=
`protect END_PROTECTED
