`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rfwbo4I6+1/bpuJrsQ1YDeYtJvMPW7EbZFzVVFbEono7GpOoc9Ph8tq3vvzNH5/Y
kAocVO768XGXufdx1f/NPb3KvWQljQDu2iAhAqqrp5yujkut4hAdjvn+B6D29Cu8
XFP63Xwhqcvdrh85rQwvxx28kH6Q3+qvAKyLIGCKZEIZTVg7txn+tCq1YsRlyy+5
bMCe+LCA0qEM/gkHzmX1gTf+80lLnb9is0ftuI5IC21T1kwKHr43pMG4MS8CUptx
uAOCTO5EIXB7wApigC/mbwn9iWQu6++BO9h/1GDSOfxTZuww0zDRdQO0jj5SvoW2
CMP9eBjsWHxsonxefbzciuqiNeSYYI+Whkeqok4Ws+EHbdQukWkJIRlhu/i39rUi
bwLl0G9A4snVLLGM9FZuaZJtr73nK+VNuufjPhLL3YEYeS9SiEUDsGvFUBVaBMyo
TopivExadomzIBF/ALKhOr1178xknUET+u2Iby1lFbiRzhi5+LHAnhxGIUeVF2H6
`protect END_PROTECTED
