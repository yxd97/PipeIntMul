`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3EDNchHFxqNk4jmApRsqDU9/6ZJP2XvsA+HKDMLjvswbvsQ4gq6gzAPIrp2Rq1a3
FpLfZ38QRJ5DZsmVMc71+AcV3mGmT9jKcu2nowq6kBR/vUj01LBXwargPhQk8ps5
bUb+I+I9bT6xZk5rZG06MezmKvlQjFJmMe41DVvKUJfdmeuzXRW1r0Ju30XlQDPa
xOmaE+3Fes2TWB+betuanvxzFg593VMuiWMyo+EXq9g4Zq2BB7zlvqAGefjuMfPT
ud7y1heAqSlLe9pUGEidrmnKfBHXcY7PjsE/ieLLSv83h/4K18fZl50XCkuYG6KY
qu9E53gIA8iCHDAftnsB6HF3/3RccXykw4EOY8teakOpednT0rxiJk76KJ7nrv8i
btgRuiVo/KeqhhMpvyUIVwrVt05wOyd9q8RHhixYamIhXr8GBTf+xAi/fHbE3Gqa
4CB7qGWbdsnpDoOb7plRVc8UD2UiHWdhbtu1qJJuTlZE38jexGv7/3eYBWKMoknG
ZoYw5u9WCVXhdIkMMnh173P2wcKyxyJGSV4w27BAPL3VIa9zOHNEqc3ywMlGyGGj
`protect END_PROTECTED
