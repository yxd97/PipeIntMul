`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
diLPubuVBurknAt2DcSIbKj/Rh8qoPC+snJ2cYLr5i7D9MCaBCyV4vlUVq19rQBi
Nu5PcDaIm6QpvFiP0FXyxS9ZReuuslKdPeVTJJLsPvBFVw65t/mIOevV6OepyrNR
/njJVncJH3E6dPY8spF2NGRrjjxb1n++iANdJSYLQ7kPxiLnJH+N+gr0B1TVWFpL
KbHFBPODK6AiqzjRYyaslw7Y0NZuYSurrlufyAH9bFDPN7n30lgDOyqBPcgL1qMK
r+oYp5KR289pRUMu0u3QbkB3NnV4isssK/hTuTULoHPuUAK+cJKAi+v+5irmeMI0
svYZGA3nDb56uQX+etzfrQ8YX/MdRkXj8hhNklATApYAXN4Ruq7Us64MUqDJCAJS
FnbaDUgzCYK/xaasiqTTUY6GIEYGgYRiZ2ON6SdF28z3cX1gj4mIwsELetZrHuDN
CZvv6HIv96K3YxvoXM9L+XAnz/V/ycPRZ3WN9TJkMvxva9lP+JRONQTC5CHgtEbE
rWzDwL1gnG7qFQLGxxgpkFR9f47dhEeLsBw8t2YWXAMgGy++L0tqv7+QCnKF0rQP
kmojdg5iqSr69r07U1+azTOq1DQK7wYlmkZ89U6x+caR2I5rZLNpqG2VeO7nld+7
dD85bEoV84ZrHS/d1+1D7Q==
`protect END_PROTECTED
