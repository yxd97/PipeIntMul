`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdtkPKgBAiYg4O4LGh1nOcZS4qEpu7MfSpYuMqlSkbWOIUTaeB4HwRLNwHyCdJCo
lzKVfTj+d8RoKUGnIaLZ6GcWKBvetqu0ad82MXsgk/stCRShDXyY9AF6VO50/PNq
ZG7txOHmk7rKQ5Wgrhglj3Yq+51ljbvLJNLRkxMrXMbZF3teltPAJXj2kg7wCYnA
FTzCBJHG39VQianPVLTVRmGByqCKAng1rca+Bk80fQGS06z5oRP0ErM7dM+CBW1A
6jsctl6Bxpq7rAw4DOugRozdMtlp2fyxRjZLk6HNLvjhp9xkPdU/zMDo5tggMS8n
q9lT2BOL3vF2LKAe8JfYIUMF0TiEfadEilEupAgFvute9tkQ1U/Pa8/MX2THRKsy
v0MOUcmhRak0aDyyLyAe9jqO+NO3wWxicGcIkFRewWDdVMShH3ihV655orWhO2v8
16y+kdoVuzNmF3GQFhbrkhu4Ds0Fsp4C/ZJ02Z0ceomESQEUAhHYFbYtowOigvT3
KeG5ehdhrUKjcTg56NsNBIzWStML9uRJQ5mMxcKGGZ8J74TQiGXzzBSgcxwJzvSu
HzeqmTqtKwwEF0ujNJGeANV1uCz/B5FOTCqbSeH51Xw=
`protect END_PROTECTED
