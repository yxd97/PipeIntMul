`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lesAHdZ5P+wGvobjPjvrZqUQIZwV0PFd3wdL6QBvhNWML8MR++dzaeXl5d4d/li
laESZ9xRdG69zFOqItDCSHKdLK9XQ6TaVnRmCOIAhyOKlilbzecoAal/GAEiLzX8
XnOLM4A9alE/prIFabZfEdjNzE7bvkgEwt+kMmVcLNnsFMJKElciA7l7KnCGmJDa
dLnTOYxP7qncVVJsLpRkzKDVv4mt4Qb6SJ15RO7j93vHYPFu5vU+gqmqyW2tw7to
/w0jeMpv/Q0yVJ610IFg65soX1UNtq6lFORCNcHgjg01rybJHY7O4v5KOJtuvv6W
TxwcrPdQ66+Gv2DFXjh3Dq2s9bQKElTk8ASXZ7hViaNoVhw4DXG+LKfzyZe1uzQO
f2i2hWVgQG1wpj01P9W53oT12JoHTcyKaQCrxrGxjNkCZ7AXZO5MW8cEA9kBNZwX
nryvrKvoR6a1+hJi9mb6LHIkZo9I2b7hvC81wTJPaz58wtCZrvOZJdhs9dzIDirR
EOzJyBYSyy98tT8NLiEAQhb4o0fTqh2uoHSrfC+Fk2G/iqAnqLRGfsMXK0mv0buu
NvmcxrIsvRI2k8BT1UKh6n6b5sBNsYXZ02wW8ElgFqfuekf0RZmwTaw+p6OMJl1D
picszgfKI6qOoz2haiTlkx/JQF6819Gf6UyWCGFeIh8cW1gD/KT5LE6OztZl9G0O
cPSzKi9LuQ8pcCKlDmlclgpg30HFQHLW9GKmUOSxQWtdoiawoNZauk9QZ9ROGtIH
GXCTBtrojFhgmmTAIJdz79CwO8UWrwq/dLmr/te8ntikrjKZNdLnvLUySXSzDXau
2rVWnAnkESe6/um1Lg7t8aQV4IzTVvYZ0l0SBWhSVCc4kTeEUvfJeQBbOp6ao55I
zggdooLfVVB1Tws/KIoSMwrlge+jnlN6jlE8xxjzpaF5gjYTKpUgZknl2zvC/HMi
6T9VOAHAcooUhPzmlDJv4MZFicI5dQiPOp5bQIze78yyJzHUjoSuj4l3Y+/6JzgN
UWHxBUikaIVbjKS+/uOxzhxuFW7A28Fe6AzbOheErXbgwzi8mHB1IgNPqYCdCEy5
w54cv0luDO3R2k8u2R7+h+KGDHEpkqEUXUnvzbJ7+xDINhzm5+km1Hft12bAyRnD
1hkyLSa3nmAW0sAeQaCcv5tVSbTqdKwaSTHp4DYZzFOGeZentDQEJhBUdnfHkShs
tYiv14RnMQ8podrLjOsz9mAq1FJw87fsZGr/I6s+3m93xx39llHDlPbtC8N1zdSU
uZjhJxkvdYdySurl2sTMMzbmkd51teWI3eZO6yb/6l+s2kahljkEtERVA8pXHYcE
bNrYxQ2lGJAs38k13ZT+BgJWZozuDqKnvIbQ7bWPzYXxRAaw+GaBQkXt9M2MKH0V
eSloyG0fzpph2sHhokzx/9smuoVk0j0YKKsgjYJK9TNnw7bs4v+0U0dOGVxVK76n
RqWlE4DtDobIhTuGzm1x2RLUgwgyOd2ByB77gOrIs28z1N8ZJrL8Tu5AYjPcCjtZ
Dn3EvkJmpyQ3JDif/esrKAtRYaS3EyOopmZpmvzY1RAysBPFzqvCGcZrMJ+Akp1i
r+a4jB5q+09d4ocrK7hVLFfZlUsZNI7p2/TQ28pkP7kysUSi51n+4bwBT8m1fHW+
5Pp28mr0R7nMNRdufHeJGiv5DcbWj7xngMZXpjDvB2ZvlSQ1Te4XeaxkUFrMBpeN
kbMH/g50dOMkOZ0zA+8dadFfJhVV7qjtvj5Walt+oPVVzgJJEZRbdPPPXPI8uI+w
ik6X2ITLjekY+lmxzrBpbf4Wm6m3q/CwXdF4sy2+A3Tcr8TCBtDuvtQY3z5zmkQ7
adszms5eEzmDTMnGeRMQ5QZtDwbrqr2r/Yp0EMtagbIvr27iGOdIQVExkAqCsE/k
prF9pDcgjarlMDeWYAvagROl60VVRV309J/4nqtxfcba9uVCzDYlc0KEJjJJVC2C
3ebDbQIyT/+PFclkUYEt4eJBOotc47FzSMr+G8l6yoavBZR20oNJ1bFbSGD0yPBE
+xebTplnW/9/AcSWkJM7hxdczFnLa5yIyFqeHDnIj14YWuoF2Lx2qmhc6/AmPcB1
HTQku2ueJVg86i1JkMHGaIPnO5CWVbL6/qkcTqq0BCJrwcGhTZlFQRfZGum3gsOK
ssJ+N+q+6nyaTrV64svSgHGKd4kUWROA7Y2StyNn/NlhMZkTT9QAghnBPQ4XXwxG
IHmtvl8JJc7NKe4KIHM+iYBJTljFXmUVPm6OMk57lmIFXA479gN26kXVVvHpAXO6
xkBBicdGJmKUmcvQvBWIfKW2lfjMbxZoksllbMfMT1T6br1/wkQ2x1RpMDOz1xWX
eCQUOnJEjb2OAcSnUNhmVMpo3VUpBpDt4njH2POFgoozVsm3mk6mnHXtbG5+wKhI
Gb2bgKc8AsdAAgyXvPC+ufYWnrIfJjW/grYZHOSGdaXc3DpdjgnfIv2Mm+YB9EjX
2B/JepNWD8UsrHjR7/Q3AnDv6qu9OjFK7Eq5F4ZGB/bBGXAJEcrSPmQ5eatdnPl8
uraJ44v4GPsRxBM39itjp5B4Vsp3FvcnmhsNrO7xZyHWzI5Dr+jy5+fbzvnU0KtG
Nh51ZXnLUQhLXsH5UTTG8YqqkLBF+0CCAs9GrAWRQAsNERnce4/BMNYHCSMfVov0
hnW8XPYJAz5l8kJpFKXsGsy8w+cjkofId55INJ2qb3QfD7DVXLHdZQpkXqsgTe0r
OyG6Qkk6KjJ/52O3C/a18t1VUjJNG7w2trSaP95LyEPN0h5SOkGEP+eD+NEDrLZj
gh94sST/WO5Pd0zfuE0N4dSiv4mySMfULZd0NuROkd9sWMVj8wv6h1SbduCj8Q+d
6cJlXQTvQyM7giJrLud0eDZrcF4p12ar71FU+/CpbO29ZloRkj1hj0E0SE1MgXMU
3JdsZP4GEkVBgVGcjFGLH5YhCBzWhmqVX7jgPLN5RLG4bqzw1eK1sCyLFdv1ArxY
X2RGhNzA8Xbez7B/PmDfLvVvqLSRe8r3bMTuRbb31ZFhzxOYMYNhksZHutH2ItSZ
tqYMAAk/Gdm43QIolM8SDugydLQDa1AZr+3zEGf5wSYgrHAGHI1Oe3NSG2oXiFMX
6tRrn+91k6D4Axzm1eBSbd6yOo9dSwra6M3SiALLMxhqCEWI3+ys69pX7GHHkvKB
1/NJxLuZbvccYPUUyBjllwI9TrD0m414OjCVIPvnpCwC4izflyhQL9Ywyu/1eHAT
+t3k2HDfvaNVSEkNxQ0rlgE+4Xw+tTRPqE9Kb5VjXG81/YnBcJnUxdcIrSFy8bQC
4VCa/f1VAFR3EKh0di2WUv+ZieAZWMgPeF086KBp29yiMf2Rly/jT6U48pKaQ/FH
5cVFlWhrrtNVAT92Zunyg/o7Pht1/rQXPMAG8SUo8Vd2qQW5M82Ud3P0E4sFxpai
DRc64+QrJpqN4+vrhcCWTgr+dBOHnuCGBCIrTVy4m0ETu/086TMR4kK5YYtHezG/
ZX04ry9Miy8GVzWCXKTG88ZhcBkqOm4suVYCjHNT4m9jcU8AKrMjnrULa4pYCpK4
Z27RnHqSBPJA84J5m8R/RZf4TSC5lZSkJgw+eAy71AeFo6KUsXnDOONbTJQE10S4
EBPytCM1Ga4fA58NwqhJ7DLHiQQdHCv2mY+LPlY4D3291g1P9a4vDB7WAeEMEtYd
ksk9C8hPb1jqXh+O/riy4EFEln6bOftmkp7fwUDWGZgaBFJkKYEEwkVDPKXaGHnN
DO8t0i4sBw45NBdNIHc2tkjPfGQ9qyK0iMoiCw7ofTfHst4n3M/gN6xuEXE7atLt
Bul9BijcQUZ33gCl9D0yJuMCLDkjT0lI/4DWJ089XCniqgB6++IyEpikGNRRFLLJ
8b4ID1tomrxgjfpkZ7BvK/tvMHg66fxBfRtvv+AtEjJuan5672JwDqIC6KHOymI9
1Q8K3rX987cikHj/gea2+wNzuyQ00+lTN8DYVT8JqnO3ZtV2juCX6P+8QmUtEpdg
KrZ++w1S3WQtnRL5TwZUIC/8BLlaMlIwLxAD37uZmG0pHQgmwd7iCVzWQKcwRV7G
XsLVmx7CprHR1bUREUhF2HJRijEJc93H8IMd6qOsLCqAsNQp0f4In2utEDW1WIzd
kMKMOn/66fkuFzJTVkwQWiTgns+ewF+gHFvCOQZP9ad5HXslihbXRrhMExgHdwBf
Xrv/atGgAJWg9AmTzZ8GMdcMf5zmBHlxXq55fqotsUJMHccTiEaJHpw3LNHqnLEU
zqiYlgQ20q+RGklz26VO1UWiBvr3C4SeV9+CPaBu+bOIB8UMVEISFtN5nt2+qMA3
rWOOkOLxt0Y78Fq1QmgY7JrPAh1DxfKVeSHwV9WPThh2v29sUDRbpHPqbmUWUzUi
diOCpYnEhViO0bm1VqtteVRZbTq3MbYAEdMr48H9380vMLBnzLRji4Ac0zUY3KzH
Vg3DV/BJpHqz0TSbYlf0csNce3yhgTjcyzfBn92IzjhUFnw2acWJ/vCJRQU3pzDE
UuWRdJ3HK2aMoCmWgpIjnS4AGoqcWXg3gAahaiMrpB0M9L0zbou/Xybcz0NNTX0y
V5D6Mh4ggVc4/H6EPbyrKpAlFlxem+snzgBpqjpWWs25FHj+uAO4bN0PfhP5Aisf
joK88M6PnTdoXednDFFcDQyd3MttGlLv1RCGfOcBhdw/1G91RgYuTUCiQKW88bfj
8krQdZOdjMxjd9EhnTG7qSDvcJ/Zg3qCy3t0/5SE9vc6WNNAG/5Rjpu8oQAcaQ2L
X2sLmupGmpLRvlDGEyVKBYJzuu4cwd3QqWrRRx2kEydcVcw6n39UnTv3wZw1zTLt
Gu/qhPHxoQVvaA2WIiZvLfgOzfItSgn3gApUWQzo1/c+w4TQTiICnMfZqLTG++2H
LNLpBvgzat3FBO9ADHw+NfXjhvinUuvRMiSCVhMw/0b1Wtlv0ytk7pKRhqstBXvT
AsMeMOm7O26HVKH3ZQa7ADRZJwBjIxBH045H7Yn4pJc+Qu94MjtRJfghteCMnlE7
S9lIIDtKwS679IAdDBa/tAC2uHQVJKV5fk60vWPIm8M0e09KvUxEeaHwOgMpF2E7
RWwGj8/tg4KYb5KwfwNNPMU1wTMBYeoYBHvVS1jKkDVpQaSW0btJk3ThgiyiigET
ZRQq0i/5zNFCwjEdenSUCgHGS/rllBTw5VIQTNu1yWv3rU4CjWsKFq2ayWTv/5FL
pwNQUimtHF/N/a11ScBFBfwFOxyqSKeRaV11c9jaBc0ybHRHqaumHSGBCq35g7X8
ltAJGc7WlvzsXkGkGts/z8S9PD7zMh3L+36vhjQ+zxWqLLdnsCPBmDPjRZHS4HBB
jsxG+UkdkAq+D2QuI4VrtWlVmLFceJf2nRi1ZsuURvtxXUrQNEfFA6+JQb4x2INd
fcUmFSefBz3Xcv2b5DFp4RYQHUHi4Xeeg9Guxa30RrGxElyquZrEnbcsqcswU4Ar
+MoBzHycz25TQLDK6iaPLl9DRu5IEsdp6i8p2nD4Yzpo6Hcb3Jj3R/PiFHDFNS2U
W2SfPzOoYWf+QCXD5ToCg5ig8Z7hVkjZyqJg4h9Qs8v+wPqdM2t+nrMu3Y9jHl08
Q3prNMMNmTkKv+tF9B5z7KN/xp00U3NgDcaaK7LVyCDEKUwEhr1NJ5A0wYaHjPAh
mUZk6GJP8RokJz0BvRHwkXfjKfNx48A/QeAnJx4KkW7nMnESeNUR7iNRLck7ZOrE
GWXS5Cz/BSbasA74lhuKgB0KMFfM6lkzZxBKcQCwaM+r7715MICaELUPWdfW8sMm
Lmh4NJW4EydVSm15pp+wV0ptWe2OKSkq9HdNX2MRhuMIY4D1Wt0s00DO7mewzxVz
H3ZjUfGrRgrFRzFSxg32BHJBLAT5uNmarRJFIMESZoo1s8/RevRZCczqd+WiohMD
y0rhHMbi76RmCoPql94E9mcy53PaAEn93q5cFwqSEvfrjX7AJi09IbUr2QQRIWBU
ffb0Uz/q9WTUPqeUEE009WCFJa1e8mgwOdud10DrN45kqUjbfgUswy/5sa6U7vwJ
IBXHot81F/oQXQ7xfIei7KTjVvayhyUe3ml1oISt+v4hyPmVQphB1gjwlm1EhEB2
vgoVVgCUltaLmvWbnDkBMTBYeQp6V6bSytdqLzcXDfOexcs0aMsHxA28ACZuUHVB
J3ie50zNHAHdWILTUhoN9Hxi2nyLpn6UhD4Xz20yBuH69oDuckRH5JrgW4Gw9n4K
lkgHqi0zFYN+oJPlwigoLdIft2rllyWm+TRDhCIBxRbbOamSYDx1Gtv5hnTba9YJ
ugKma9/Dty11mRocVsUJ6Vfm68ZFSHh/ykkSgQodcWSWWn+enW9H86PeCRzTKHvP
sYWV8etCHH6Z66YbjITfyNCLcFdYML+oeKMJMRb6cDcgnQWh/qNAlbUzX/SkoemX
IDDXTrX+XpFGGm5c2X90fKnfTyx3Jd9UwmAugX/WIAgybRU9NApGaLG/pyb/K7iQ
ktlYZL0DYbeLxv1hGyisfOY1AhhVW8sCaZPcZ4d1d7c14Wzpw8U4+YvGMwl5lZlg
tlBW1TGLRiRk4018mPJWtRtXtY/zeZDg8YEDUxGoTEMnqSIBHaKqSy5H7/wsd4TJ
9WXer26L7yys0G4ZEPCAPcp1t9sqBdrcqkddFVyLi0vJ2uHk9NGYaHMZ1T+4XT1M
QACyloId6mRbuSMnvnt5TARge2NDVfEroKfgFCByGDy8v6zFYbKJ+9rrgPqWnX7g
UXcbhXFlX2lt3Gdq9oNxAupKxot5nYB3akP1tzZMMr7irLKU/+EonBZbAyNJOVnT
+Rpn8IgfqqaUgu1ejgJmwRuTCZ7Rot/5qMujgEnvec5XvNjt1JnL/rRUHBpMSh93
8oubSnB7SrsleIKz9D4sYCGZ+yZ3hPjREpQYvWaToBWYzixWouAF1ljcQOgj9wiE
LgYki1xmQ4XLsIcia84OeJ0pQ3AW0n2SFUtqYPVH7Bwm3kfqdizIck+gfVPFiNhA
W8AXMgyX4tucecoDZegmMs7WhxkWzDpKwX6RAtAnE5ISzbpqRxxAd1SuHpv08qIU
OJBpQGtDg71zUmChkY4JZ+a8GgTpfcH4IIS8fnqCpWX+9Vja820nw6VZFAgppEBm
gI7j1Cvr3Wx8qWrQzKxeAZ+vivc7Co5RM38BT2GGb6H8Sro7E7bLWHDhvGwqhYtP
IaYtal9bQd7GJ7zokXcBLtlRDhhK0Ypa8EEMw/3+nzBs9vQzW5/SCHJi5LP+oLKO
QY45xSw2RPjFsFmigXWwkY6HZNi2ksLPPLm0p4AZ4l7eYiMPxJQMwZKeHnuXtslJ
1+Ki9PAItQs7PGKvIAQjvELI5kOfQlueNeVoX98ctZJ93THEOir2IxG02sYatLAS
U3MqZTh8LwzSb/eA4bSUrYa2JbLUyv+3OuLL7vO6XnBbU6g6BWVuovsOlHJRi4fL
zHjZ7ITaMK6Wj1zJAc4LPusOdoO09XrConGIb2O4u1ioHbcgMWKB4o/fDt1J7NDR
X6KwPYxySZTceTN2TOva2PCFncLLbZtp7IE2sBpojl7j77oJZy8hdXA1GZk6N4A8
cuBfNbTWz80B2AQj0QMcDJn8jxd4NAqrE+ocdYLnM3tarb5Op5bfH4Jfd81GY8N6
NOAgvw7f90vMFFyaTe992DdXgFTh1YCjWYFTIncxXtFor7PgAEhcoeBHj+dg65o2
IW5y1KISONwzkA83b+bWqSU7Rs0ZWYUwtO/yrgkk4JQhNid9pPDTRBhZYo8DqD/7
xapBLtGZcsfTSz0XYn7jjGCBiH6AGSLuNpThWKS3bu0+F5k/KYPFPmo9E3bx/N+S
f4Uz8hqIu3fIE9SHY3lO4ddCxL+ourOPPnJtYpA3/D8tVl5JXxqMD7mxkPKtKiax
4TLbI/PGLd3cnbDN/yjGIswtWS5r5H8NJGaB/Nifqp+f2SbNDziATUOcuO63KOzZ
Jh8OmdeTBf9bvqbSPiC72gNERNEeeNpg6jFDAN6nXRprslaT5jNKS4Aonz7A9lJ2
jXFW7UylA+aEOMtnp6kIp0ucNTIMcz9MBPVPUUq9OpRVy+5psPni5oxPE9qmqCeT
q8JgVx3s9U0a9S41QCY58LQTBck4x+xNdcwaKvEaBSq8VhX7IVacVh0atmROautT
EZLb+nmVD4rb4a2q1vih/9x6ttSLxxnqX1wzzJxnmRulmsuOYNxAWBEqeGH//Z/l
CA9LvbsMD1VLcJruObE1NPTXVjJxXqT2tF6JSluVY5H9I3ZBiY4Lu4X9m+W7MXNW
+S5DzldQ+dmsKdMA1jZb3aql/IPaS9GngaQC8UWS8Qgj+nZNyAvTpsz05mPedgG6
pURAvCaMO5MTuMOK5DQlG68ZhnfC11TauOLNX9zEKqxfNrvRCK336LU6iluwe28i
e2NX9VEQ7uxRbWy6Rb838lln5J6FcgL3vK0/KKgIoJEHDSsIoxRW3tTFxPrr3Rp3
EHbvJoP6Mo48GhbrBusZnJexTCwqb8lGvgyLWc4rntPwTTUqAH5JD7GQ1JuNexpm
gCq9KYBi5zRQPnd8ga+tK/ROwnAgszEXD4pDsTK7WvRsaTuXEq4iW1uJxeDg3tid
5uI7lMEJxC9kgEza5QMUffS4NHTAYtlvfAZafcv5ZGdrXl8sHGfl7Wxc5pucApi8
PE4eh3iSfBRFtTAA7nn9HUxvQ90+coHkkciWkUyHM645wRN1ilKD7qM/fkqFiGlj
IOy1pzzpnNtqyB3E5VfJvOoKnuluVBL8VOLkkpbe7bpPsUtwGGx0AyM5LjyQCic8
48omynPfKJyfNYrDY73edp4PdyoTTJ77Mx98TqmDKm8XT0QrqIchz6Tgkn2ddNO6
gikf9Tg3yoXYRfhCSNho6JYOuxmfGWmZbtj8dXSw2B8acZg6+9wkU79iCQcAr6cU
bnUmzHcU51VtJxqJ3mNgoMKOg3ojgISYtpqim5k8LX5hyB7ctanevepeDLGGo6Wk
1uMxkYhAVCmxuwy/ZpSYWBUZmEEPaRGgDJYjc1SKYUscbWpEDyLCqmh9s7yP2PH9
VvhcgUIwLwRxtFD9by1SzT+aMcoaWCf3U9qmj/kSMoS1mMo2rTkJpTEt590PV6GD
RE3hHTLxp9G3ABsngDGdsufq/w/SzeUddFGJCPGk9u9ElwUBj49CW/pkklx7rvWA
EU9okIQ3vsUmeAX9plOIwDq7SZs5aUBMj6u6Mw+1GGO0wl8O/7K9nJB81Xv8nCqk
9P1dnJ1RW20pXfwCCzF5CYm/D5biXciGVeh5EwiOCBp5tLKWHYPUxZqLDZTzEjQO
zw/VSj+GRh1BCyAcxUQ+7B7EoRN7q8Z+RqyzDEpBUhnGuTlnfyA8X0YgXub42X9b
fEHUWTDoyLMTXXD+cPztoBXZwaVxuwOvu7rNB6haW3iNKg5t49NL/anKDB4f308h
Un5TDgY6pRl/NHZg1RERk4ia1df3dYEZ28IfmCu7Y0btFL77Ay1lvWRx0xo+2l96
vvV9C0YsC0YA0TL3bMOEcuZtLrUFr7zFJVK+8v0b6s9bxCjcMAvY7wWMjpIsEnGt
9hwuyY1OKImft1PMCpbATy1DYfz6AuhblEtHXPhIPpmPVF9VIoJ+n8auPMoREaC6
zv3D8xsNlYNsfQX3vVlM1qHVrvIhJUxinnYEiOGxqwuZyOK7kYbAOjkDXd43YFAe
jWiWoD0Dv9VAkG8F3FQWaoXa+l2thp/k0ZtCvyb96WulnJ1qZhkMEaU00U9L8x+j
cAKEbNiLvucHSDjB++caOhUs+wwnprinSFggYNWxmFXWlIuGRPQUnKQrl+BEp7jc
pd6605VLo/8n6WG0M3F3Lqd6eRNePQ6cTppLFi+5wbhHVHEVQP+Kp3MxZqRaqgBU
DZiw4RqJwxSA9QxoBKLYxe6ZniDXD1d9Swohlh6G5qiGaZ6str7jPoazzGD+uX4F
7+SNy9aACMBU7W75VhbRcEBarschDmQyqN5Awvs5CPkpbmFqC73YMEqObTfaZm1f
`protect END_PROTECTED
