`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3LkylnNg1J74srDHIIK2HD9/bns1n75ZRHOy2Q5P4oDd+c40Nslf4ceAA2/K8/5
9U2RLdxigjnDjf9FqdtpIZqqFPRPN53W0hUEkJUzTSDouKtSJQMfLgh88hOjP+dW
Aym5Trjv8+ZItflX+tUSn4VYu1raHyClSosACZrq8iO6OPRPzRRk0JMSX82mmmw1
9YUIqEZOyPUS0aM/9cXZd9y+s2/y5BPlPBL8TTKpyjwd1PVYnwd7zwbsNT24LkcL
beX/NY5Ht6ifaGH8+NTZ/LzP/mhRjKbVm9izQnRtiyvxuIEuDjPHt0KVsgaDkzHA
v03DPDd7djYdJuekUo3pRkFU+iFTQMzxbkkWevgQWuw=
`protect END_PROTECTED
