`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oqTq6eHZ2LQUG/pwOi3oIT0ovFs/jklzmQ01Xm1IbZ5PBGRXz5ZB0sBSPDWZOziz
4QlYMaiwSSqZZAaee7XYGuf4s+flFSLws/u5lDmziRAxVxGN3MU8YIve1pDMxuFL
+q2kwtCgfzCbM9K3A8Nt1W5DVbyldtq3XViGFpHwPUvle5iMAdHCIDELuRK22NDu
qKnIHy3KS+GzVCLLadMDpBAUJXuJtYfEgciyaHma1UIx3eoxYbn+9wPO+EgRR9ir
cofQv6IhzRnSb+Y3KqTp0ytHz6ARxbi4M7Bq6iXZWZ1XncaOg+mH64D4bRZBMfHP
W6YP4pj78/hfcTllTgRmBVWiZd4jEBlgQVP3EDN/VW97ATZBF56O4TZSposYbO5A
BtFBzhLwcjVeMGEglLf4WxF/SvzxGPa1rYipjaWgKRc=
`protect END_PROTECTED
