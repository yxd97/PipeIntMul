`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZkUFzxypXf7iXKP5w+5Vj0jvMrFccuoWgd+AB3CS29RsWaiPdEhzoYP4KpaCZ8J
0qeOjPL6Xrl65Douv4GtqJgrxPSH9ZfuQIrfnH/nDUBdN5vDejVOJoiMt9Aw8x1T
Ih3qzMC3Zrv6/qRiR+FiHSghGR1hcav7YMvmHm57h3bf1A0PUCCdK60QDWO0xQPs
54LZF/DbLpAQDRZtb94q7hzVsvtN7Vf0DwchL+r6nGninksrU/POhgNaQdNwFJYC
QdmA2BKG9RS2mglMIfzVOYy/+47ndMeTSCrYfz9ZHWKA6BCp/LH3oCa11S3BrdkU
oJgH4xFhMqEWS98UMsIDT+ODY38PocOlGtMYf32lMBpFfMjZ/6XW5HajPpB3tvGR
n8wRvjO4GgM/S8vjqDE9PRzuLUU6pOkfMM7yxw7hHuCZEromWpcwGWAXKTPI45oA
LY8PUVk1921JSlzOK6sWGVtZoORFqKRnfcTVbbb2cJVGxWQq/LyqBENbxpTyrGbn
xmhRdFVYLQhayJ85GrEmlIlVtXIvhe+yJExjt78snae7E8e3nQM9txyQgqQxoTZk
Kc0J7mIZevC6ewjUG1qy2OSA44kifTCdTqqcs8wml6e9svPeyakrDSDKicKKzvzx
SiD6fNuAslsYQ9ZJZt1RRy52BYYj8J6HsUxa/jvYbIQEjvitGbF/V6XcKy/cy35/
c6Czvy7TbU1mBLRlgaeQg7MY/oP1sERr32gUVvK+JyLm9nkwDnhXtTpcjOCJBppc
1hbxWa03X5OzQiiEb3VyddF58/jBF9H5jcbQidQlv4Ttv2V9JpYiisA6a5hJm0yf
ps1Ve0gbzx5b21kgRoFiq5t4Q8FIQT2eZ45ZpAzDhGBOor/H82lVFJgVuckquShQ
+8N1KYI9YiwgxhMjjVfM6mjrInUtnK2QBBmUu+WMtK4K6V+QMB5AoBmXZHnApBac
VZIu8dbesgU1Ydq56IDLWE0iOFugm3TQdoOgOhCoKNpyZHB+QcK9zDXWBiSCSy9/
1b8cQAsL26PAwTX6UolWWWQpcUVqCmH5sOxTljvaAVgpHTqveMUv9+qHRXAnnOyb
KX5DL+zcZrG+Xd3qP3jXeQJeQP59cChQ1KHAQkJfAifs17aGeNrEVcKs1xJRp4Vv
4JHRLXLyervEzlBmxwJzIkfRILUmQLadhT+7ZsdtWds3FX8/XiHw7rX516yLQpey
JKSDCQYPsxdI4VNhMDhM1TCBNXTmqTyVdey406dKR18wIc+SkGiX/n2hGhVrD3N7
GyxuGfbwApWMiubYPqDvrBMzSEQxwtDF5JZHYdq+N3AVbpGcQY+q0cqVpTfSCT5D
bR8p7o79q1jNgcu/R/ahT7xqXpyv3/S3+5eIwhLGjbVLGXd5YD+vOvGbsdWhKzW3
QVFA3fbarzzxcgmqcMj+Jg1J0Pv22oqQ0hn/K+C9H8fc4BvXwFHa8uRciIA/rhrx
8KUWj51XpV180N02vARpsOXxJMtiJuiwU8MlaNFGI2QlLKpLodedQoF8SMpraqcQ
GBGzyCnTrFNYqziX/YdGunXknaz4oQnNm0MH0I65BmhliIKwMcCX8zMrFF5J54XS
8H2UD5PWkI4BzCUoOPamK3/nFnlyKHQpcYPpF5NWKxq+FBNDBDa8xNwtpErvljXe
gOweQmUz+9TsT5ezSmIzyVyCm5QDZJCynbsJhGxg4a1r2I52U1GZYULQPBzydPyE
BRZUbUY9i3gASFUoxHr4I5wVNMeAuuAHEZCfE7/gp/lNXyEaeyJKB3mZ3SMlz2/w
v/kyjk/OPYjSAwxcGBBpkifY6x2x2iYkN47keLSB6mD04jLBTlbZmdZHVGuAEEX8
kn0alRMKI3zkAWRtw3ia+MP7xbx/GiOGvJTnY4U/XVg946ZYSM3pP8Xj3mOyDcQP
I6WPbOxD6gCEavkRbS0PhqVEWSvMgVYzzD9j5g4pNGwuk7hObwPVtbUb6HN3puWl
6b95DOMTGV0/Em0SYPA/gESsvmDecVUUTa8J8AkUPOgh1H0dm9nQdfwShjKWRGOo
3jlRjyaEcr+VrgcX4crk0v3sawN8fYk9ExV/YzwkPuTUipoyLc87zd4Ji98Kl/fg
Zu8+kdSfp8WPE787BdyjL7yInSqXD4XtFHkKAs9AARcjpynbDsgHCE4MANNWqqn7
sXEs+dK5QSkumrDIq8d2lPc6+ZrWQXZsJk/bukLTe0Q/Ku/Jgqtgfaifom+lINwA
+b1PXtplxA2AjH8e8Uqi41vf4DzJuimSieLUB1ebfOhxhT8SIMSuE64naDRUDHav
VrF9Y9M86Jgc4+E18fnYxpjdTs0pwLnOMiSvYM4BDsWd6r/SPK6SDZvOvrPLPALi
IZjljWsTFdYHqMx/scOa7w==
`protect END_PROTECTED
