`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qkrSHushTGe0Xa628HueMmuamlce4X08dveLLXafxeVqIfW/kGXGtanq0n3zKtP/
hBYf20MhKR5gVE5Tg8of88rU7tnAtvamNKAOMD0Z7wHIRVeevN+wtqg1DL2D9DLb
SW5PHB/uVidAj46TxLGL+2Ne2P5Hud6hSmRkp/tvyachJmOR4kqEei96T9H5tDEH
x/7gl8vZxsK3ag3lz66zwVpUv6W0HUaOfeFAwomyBQEMi8idH+nwdeEJU9kGYhVq
KmCYVBcl3OAFSFs/znkc2//jj/RIInkeDZJ3asVjPNApqeb0fkQxnfqFrKvNmUV+
OYGIlpNbkxNa4JPVUurfXWSgJ59y7GX6Us+d0CW2UVy2jVvFh/FfTVcQUHDOjey6
WfXR5QUP+xQfyPzYfAJbfhcUubIz//sihHEuCvh7Mh72mvbdqELMYjEVf9lvfaSV
sggW/CCga1tYn7fNzuz+nUfJXeVwJoEP6vGWbn0E4cbmHDunQWQtUtq8vDBfYsfy
jXqh0R4CCf35a7zkDsJUdafYe4JgxW2CQl1nqiJlbvcu/eeu0ZxJxoESRRp9ZNfj
NgDoAUgj9vR+2y+KpU0GFLtFaJ/fW9czDq453F2x2+CJkznpnedBaC4HEp64VPqb
cf27+lj0KewjBVh5R0/RPKKR0fwr5lXVA4xnpab8cgoaDYFyZxDEhIRfdvv4TL8m
HhC59EwkFj0iS5zKAsNuOL+QUz7xPacOBobTOdHdHVr8BpPoXK1pX6xzr2MdxeFg
tFk8WejFPqvR6n6eK1OvzcHzsSaachIOnXeiczzBQvaGMNGojTuHtgizQESLP/gY
XIy3jDlTvbrG43ow5TL2ig8iuY5L3nzWL+LrG78orAo6G0yAY9hXQMYfjpBWcIp3
EnoAVKWESBTG9g2KwoWgbHSRNIZSzKUVe+rJv2KTB023FGvO7oQFe3MMIXGTF0gz
d7VsLoSFxMzWt9J76LC0LV2Lo3tWXt4aFg4R14f5ggQf1cbvlboCDMVubpHIy5US
NToXlSUQN8S9EIXQzXTLjjGtZO58VCq0qW30GuL5QyA9GkIukztk1aJoYvJphJSw
6tyb0hnOxqaMZ4OIkeFOkNBhctxfbfC2vmGB0LUam7jRKjKEPjBnQM8UPLZEJaMM
+AkStyXM8fG8azTHWZPO2KSds3NOApsPv+iOmaM5/aBYHGQfZtXy7nEj+s/NtsUi
AJi1NRjm0urTSYJq374vOx4oJD/RGJQ3O0X14LlHntdFnZWyjPYZ0hKfYq84s0aX
uLOjAXUkb6AOr6az8mEOo+I7RVhECVsONn3cxQ2t3dLcU6o09D+FY8vJSq7szdpa
ZlEld/ZuDlMpRvjOjyUs8GXhboukGhu0rjehverNNnmQV2EYYxpxd/yGVuMs7u7I
k4wnYd/68Ze29elNAdZLV+Jt072N7lGnAmtbQqnnmUIJ6bjcbU5z3/WCAwuMurax
V+LUjE4UBCpPK4UwsaY8AI4I8Sdhbts2N4FASBQjNnvseEh0GlLW7CCONgBjUP8I
CK5+STmTDjKkLxHuM5wmTntxdma1IFHnvgHGqLQyXxtpb/6KZJvZ6akLCMK7tKc8
KGIO4opS+6R34CiSO1hQaHnJ5wUBOvcm86roM+wtC+Tqp5hZPGnrVLXowM2tp8wX
WFKd83/4yuHHgG+zXMtapuYfqwAKHgiwtgk5GvOKYRy8MvtwXE9dVAkKuV+aH0w0
XvAYE9C3b18g+Y+j6KLOt9UCBzeygOROM81ZUpuuDMmTzH01XANcn7KmszBNu/rX
+cGCcD/QL5ZWzhLB+w3QWeAs0LsOI/oWp9wByi9dYPq+cF3BfDIyxfIdt6C0/uFu
pQWLKTEekASz+MBSYKidcN/iRWBudtLkzUo+oVnaTXdQc+WkzvMrHfAz0yeMMewc
60Ur1H7rbHiboF2cuPv5xvLt3s5/iPEOUiDxv/McrEyo1L3NMg1rYjyCm4y9qiKv
YoU48mTJ7ASSkwOEYQskD2xCfnygyRIB+H+FY+KNBNJo9QjCG7cr2a1wnRgqHbed
AbNZ+Hu2S/n8bowoZW+UtIOoXTDwkZvfQxofWzf0WtmbOelLJ7x3MlLUtfXT0Ls4
24e5YHKER2k0OOUKx+3xi5ggSeA5R4WsTZG9L9YK80uKUdGWDBQxta7PzIvI97Ci
opjQJ3NNtbtPMpjZwLqNkLSmNZ03Fta+3+qRtUswyWgTOHCT3fxOtHYO7ac00zYN
/nFGVVtnzoLsCZKOJMH/Cq5Rn50c9UY4dEZk0M+N6pFHn2+LaazuXeGaZIvgSxJg
LkSS/Yu0sKRSrBSMqkxw7rOCLLvnIrilZyhF+IyQrCgEQlxaoFS845Cc6UBSkGhK
OJRPLuehIt+cA0jzbwOmi7OiNoPTIOFC/b0SCr5b+EGhe2LIPa2SNtG6Upt3Plv9
p7TO37fwEMds2aeV9M+t8cMqLFDZaSy8k/zOQupGjBwi0mEXvLJojbUYL6oDfRky
uvSrg346dqIvVNOzE+3yRdf/zsp0++e9yR+JO1Wwgjg1WrX3C5hMHtWyUirf5/VG
srwFdbFhYuNqcrS+hfvv7pX7WIIiXLhs2FuEGyrn/kfDHx2wvmvXGgttdHREhBMu
eyyTG5XoIkwLYkzEAmNEUu6nNQCkwmM0KSMTigj/BaeVQUSc5sh0JxjrYRYPZleH
n4XE2/RNzqc8OBw/9Ao1ss9UTDHmxHMO1VVZxE1I+eMJx9ma0WUlOjaoz8URuHOr
MowuxK5NWNUB9fK/MpF16Hkp5dd+QdjOVI3yB9TdXdRSA/QJtjJa6waaNTiubKoe
jmyZzfJpbkHHaGANyU4qaxthEyMmRWzO+1uu1qWpsCVUuOiuTtZXGE5Dcrr4SaGo
Yh2AlBKw63UJu85noyylAsm0NlqqpFVEOilEvr5oEQX95TeBZyBPFwiPAgSHT4uv
cC5BlmfvxyeMqNu/aV5y4dC5WnS7+BIZAfGdlcPSG5ivbszjB1Deu0oh/3L8bKgg
sxi3RXokRexbCzcPhOVHmKF8FXLeDPdrv2VLCvvgMHskriy+gjS7oUwixBZ7/Kjp
b37wP5gZXfKmZjAq05vwe/q0f/IxbdzuR+s5xACg/YreV2TBbsaiLzwheBj2LzEh
FMKc9blbHbwyIg/iVAHBg9ooq02VxJ73WzuYdzgclLX2WqKy0Sf55b1trdHZ5vYQ
LGTufWR9kZ7drD+mjcR7eTq7cfJkUfWukm64wkplykzv0xMVekoi6uLKFrPHoQ92
AIY9PxeVcDDr4fUn7YZ5XuAEQli+u+rbBHPhfdnL8aM=
`protect END_PROTECTED
