`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKD67R7EHYdOGFoJA65rBxmJcc6Ajp1Q9jJPSFv7QP5CmIBVprW+qCb/0pkmnJAg
wvfBa6w+oZOMHNpNSU/LxocmCxlaE1/qQdJGubha6F/O/qOY7f6fJhk7Ytl0zBbB
gduKNfRM+ai5PivA5YMzzE9ecQHiCzSGCuznOXIVIrAytcdzionGVBtikcZIcpmR
JyaEm4KnZN3IRHyPfMA9uc/Wd17MqbnxduKExlX7p6XYpgKFYH35RqyzUXa4Dgvh
PUFR7q/eyXzkKZZpDpvUp6rHMsV1iAe4j1huKIag80zrergfBlI7Ma/m7X2z3cMc
cb+cWsiWhgxBGOw6j2AR4Jv41f8Rhq2Wu5H1zos/z55YGKY5ILSDsHfazF+KGbp1
pflSVweAZ2sJTFUIzyLREa75HcAt9Ds3GqmRKoknTZk=
`protect END_PROTECTED
