`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aAJpzCaA5ZoMaXbgiETDZWi0PJRBeie/8N40HYUg9AaPAO9NxdKkdznkOUXP7uwL
EUafzjLid4jTYBLhQGiM+xgZCH1W7giMbWaI8yzyjIkTeI1mDFfYJ4+LIJ1mWeB6
APL9Z+mbd2dRuvkOXie21gG+R5kArM1Jwz77KfdvkA1jF/gdBLude3MmRMEzE/e8
pD+J1bSENEZgGMTGvHQeQDl+EuCX3z4TxYN51fmZbIP226mafJWyVDF9wq0AqQ/p
T7GYUyhaiYLhJYHoJVHTWC+164b0eIrpsQTf/6i+52pEkjqvQQwEgdSDpRTm+z93
l1rzr93mmUmCYXh8a/CzUzX3yJNScRLNTHwYjCW0QZvBrqDPyMa6F4GxJC/pYneC
JpWhrDPgkVuAgyA8X98BmenwBmJMdGA8lnUcx52YW/jVk7z7depBiy2zKFHXgj7j
qGndw7a1U97HykWboShD0hoqHLOLTcAtHvBiyl9qOEixPCEepiXFJKlmuyrQ5ZD1
ddlrOntJ62GRyoD56Wd0wqAjoftH16TApDmu7w7m45H6QNftkreOkUI9o6qFwpim
gn4P8ZQGfAPUgdyXf9joBbp8DG1j3zvc2M1Bkb7jmIHiVq5NNhj4jtmomoTpfzr6
qtJTbmVxisa0YidPFLWE5GtffYWzPcqON4MCF6RQzG9ppKZh4oLELeC5dASwGcOj
EKdgD4OiSZxK0iWG+b3q6Bl1eFnnvskR+ly9ALzbG3F8wD3Xz6G4QBoJdBFaUOyQ
/7cNOQjvtV7U3vYBJUJvUCo1qPC0CA1ahYfcLMPaYJW/OKIiwt3TazgnhA/gzKKl
CEd7otSZ+niZRVXV7lbtDYCZtDhNM/WGotkdS/+OVs1mQOi4xJkDZvmigz9BusuG
YbbBcPYW8vEkyXUPuhWovDK6z9qv/cMCQkcKHlZ0Xm7oyyVhHaij8pNY2VTzorHM
KGhq6y+A9bw+0lRxnglBYRijfJGhrY4jptwL+KB1GVqUAyoLAVN9IpcaxRpNoVQ/
rK4BOrl2sQSQLQfyP+g3YYZgvQ06iJoGpfVkcuKnN+Gn2ME9TzNEK6g+hNwb8yAx
s/arOt8aOQAJWrKixhyFEpNTfOLAV40rV3CmyNuJFY7RjX8/SdoZ3yX1gm20gXEL
q0OsnjYWSbkYUdifsaYePulgZcEA0PujFzptJrSE0iMSXUNKkkWGMf/59y4AeG2P
KW9DiIBmZmvLSaOL/LiJl1aSbwzdvrgCQnkfZpDBuGP1bRgEPYpZTmrITo7NhXkg
Y9VQZKELFuDbcwz/wljWfmtsG8DA86QquvReJ0aA0T8eKEAnVPYxRrdGBSYJX0t/
zjy8dK0uAe+R6Rw9cjW8yjKBelEInQHMJc94XFDtb6Qcfb3YDng8v9R0+0e++M4E
Bh1rpLN48d9sMYT9P2ScjL/Fw6puTgzoxfQEejIsnqMJFMuiZal4VztkMnSxjiDf
AEQc01GZcrA4QS9LImxuLGRFasiBOxwuAAdU95u9MlnIy7/7gu6kX3CXL6OzFyuW
TvTWRCT/Q3fpdvie4OaYPQfrZI2qxe+gCj6feqPrlHS+Z5w0lIdlIvSmf5XTzb1Z
dEn9NUJOegHKxtkwuQOnf7pLwq+qPZeAYKv/Vfpi4x1yXC4w7jiGkC+gx6ssd9wy
13m9cfBAMPrBawjCTgcYrphRih1Ddhk4di1pEuJCYdXps8fAZoVJs45DjS/bh1W/
28dQgAev1f4fqjVmt1ycSsp6cYUyecdNMgtqRR+nm/HYVpFYJ0S+gJD0kkLeLtwT
tmQ8rvdfKMyPyScTC4+mFIvkcZNWr8kPsgRKh4fNlKMfnodIDEh44NmDLpnp202J
UW9QRwD4V3+6ralkgLZKPYJx2IVAfumY/ts8gaP2eWL04fSBG5DY5QnzpJBpFxNe
MWdm7D38xUkB/dLKIgQ233sf5U52gmnZE7MAI8MzGFPuqopKRdbMrCeHvEOsr6JK
C/o105HfsFaO0zl/C8oLXP+IRxMhpOpYkx1hmMiUHUmOEuGJe5U6GRW0gc1uDL/b
gQ8dmpDruN/Xormi37xhY6M6ifvTRM0AZ1gne4gDhsf4c4KoL0frjFarvM4Zb0Kh
vpAE0EFb4xTyHkrm7O+ezGdSpLr/N7t/JpIWvbbv8dbmThESLUmpjfKfXdwnnTa4
MBvW3rmsdDlrugURNCB6XRHu6PPyNHDVy99g+1PYw48ix3jOEsp7dfWHXi5vUv9R
MAgePPoDGKiXUTkUpp57M6AQIxxNJJkmS54l/JDc3i7FbS27Nx4rkhhH9tSbBaYJ
5uLJVYDAIgxYMjbG3OCv0BhK2LZRqNNfZWo6fFgGPB6q1dEsaoNOSqV6HUtdlH1s
I9cunsWBGneLC8Qn+gLVzc05Fa4Qy8woX6IbL19QCJv1mbKhniZB6HBOJPP0/O5N
HCozokoNz31PoTins6MMQCl8deOiBNyoql8Sdbs68UZ+xVdhZC8DgwM80uLdd+nc
DOT1yRvg+PnT8OnSg/ZoHXxd6D/J7E6ML0XpR6SYeDIluVInpo7j/Vtk3xKEA0tM
iPXwU9Fe/36GIeXlKEoPhe/mP55rJjqkNuq2G+crj4hUQXG8MLmI5pDqy42JtMN7
u2gKUU4XsCNwXaV3OGV7vpt5N0+lGBKD1YkMLf35tXNG59cH8U0EvgyPr+yBgeUV
tj3Si9vtvY7qKQfwKIG6WUIEHdFiHV/ZGBulnd0vrU6WDuNfAPNw1pHtEIi0QDs8
NO+cEuE3UsrZWtJKzc/05OkqhaxkG4ci0lvwBJQQmSZ8/cKxfYK8M80ExIJCVO2U
gllY/KESK6gZhfQGIv92OoFZ3uPMZvGGqELTcoAhrR+pmHjmkB/MoK8RObDP2d3/
4euaCsSGhnwQhFkcRXnv6/nJIGMCJpCaFybcX1NhS3a7B5J0VvV0CjgFM6tLyXVI
QWuOnoFkyodrDosB9T8pZi57/0IHQ4fLBDdcUW9/oRRgvr2lHYxNu1Jg7GvRaHqT
odSU1pmSvckhYJAexgBM4MvP1FYg0s7j4ARFafJtA+rWwYgZg/BlPXzYmNnZoz4c
MRz2GrGZ2m9w7ocl1pL89jCUg4X5Mg+iKfP0JnmhZiIlwbypGpAfp+hvUjmeRlzC
oTYa7N7FAiVP5vBVQ43Z8vGRrggb9Pxvc0i5abbwQVBufpJKmWyBxNkKj3TGNNVy
OjXEdcWMiHUqyaVphAnNLgLAJqxE9BG/RM2dEtLxk3zAboWcJspz9ieKj+L26xaX
eqa90F1pzCYGZn8SUgvgBxVy9gg8LBbi/kC8CDWf0nQlJwtBPLS08D3aDeG4XXSq
dGnGQa5hlk5nyy3y0AJl7o9x53nyUvVfFi+4m2a+wPz1PKa1sI0zbt4Td7YHtfiX
O8DMazWrJtj/7a/aRcD2nawjAtKoa+tiAHMawywcqCerMBtBsDeefnw9YA0Fv1TI
AP3ONxHmFc0FsOlN8dNWpMzEqfLrwm0aNw9Axxznu1SmK7u3IJLQwNURxTo90Xrw
6/YpRTLpOPoZkbuHXldbomFnRv2drJnOX6wx5vtW9QeU0FrsIyWeDyEma2iQt5Y+
TEi5eIzs9uRXyQNCvD8P5Vn3Ghur5u6H6vJVy8p/qCUyNbdzPmnoFmzY+uE5N3Zq
GEfgy3404ELeMGid85AdSQWalCfSTmhHTCLUA2TzyjCmlFlojDRI0CCPw2rpcEB6
ENtjdz5y7JQdl2f5pN0355fMZnYX74jJBXJapD+YrjIDAKvbEzwc+vtGX3iFxrVu
QxsBb4DpikwlCMeDRsRc8Vy7H7uB4aPM5Eotpq7BQlTvGb7e1xN5GPJAR3V8OxPI
iNbLeBUl/wXJHGqgIL+vl+w2lbGYVmft4BYe5vHv2mCvU7wbo0vkjSS6bgbB/P4z
FGQEfRyr6tZIRK4lkcAdbvj9cYmQ2b3OBZAts/ms4RIrPbhya5N139KwAu/eyYDK
eTeC95k1imkjKary1ntqe9sYNnpNHOy/vlzX8dymV0SJZ7HUQbjbq0o/KXUxDOoD
pcSjkGjsEa05X08UogGDAbG7cBmwqqvo8/OZBWKpsTbx3+7R3jSlx5Kp6s5m9klg
1BkkV4NDhR1C04+CtPlFsv34Zar8zO6DfjBTz/oNFvlOyUbs6Uefruhv8e3eQr5j
FPBQPLcSj2CnXNHQNH2IPMHgyPTUW6kHYGyYpI66Lr+CC2dy4kQQWPdX1AF5Zl30
tGh0y/kPwe/ad6tetA+57Is95euhFzia3iuSOXqvG48XSeYGlPHIflw2vTO//nMx
7C8jol7vl/cZTX3kkMS/iionVdjIdPrDbt6y0rwX5IIlfAKCYnx9zmCANK825D3T
BzEexod7/8HixV1s+pbUMzdog6b0ZQHGH08wwTzLiNSSs2rp2+k7yGZ0YMVXW5Hj
D6QdvWf0XlI46liWzjxcwdnYEOm9qOxWLNJduneZystiGYEmCoWsTF9+dKlMaFvD
v60IeltkNixUwTkr3h5nf+etlKhH8iHuIZj311sCBLd7wAa72BWiNNn20CJbzant
FtoazghqyhqH+Ra5o4rSshG2JvJulbVixALZH3sqwnIyNKXCh83FqyIOMbJxkfgL
xcr+q65CsIUxxC3iYLvJ8rmm9zgZ6NtBkkbdfuJwlhejcqh6PPondl4Ofh//YRFi
ngiRy+VW3iCVVzaMWnQtdxAydBdaGp1LRRNr9Z9beUQ+3NC0Bpr4+5rgQsYsl3OR
T3fQaDaT6ognLIdrPs6tB1izUmB4tYM+fgOauP7nrb1KPrdLMp4vjJo+F341444K
qEeSLD0pSg909C97LwtJlU8CDo3zNEwsletNG6jBT3VMfbALsG96FD5bnPmsXyOa
OZxXL/i8S2o7+wb17RfgAX693xWATyvjNToiFE3vZD4uuqa4B0uvYnJ7PyfolaG4
igAK7dWy/4ftDmEUYx6g0qRpRPlUHvzuxhzaO8PV68Zt7Ym43re4gBGzzHXwwQd1
deyq5VktcaBBayy+Q5PTITr9+uZ2pVOn55BZQ02CFZJlV3zn21ZU03PgfLm1Ujl0
xdJ5gzcOpTMyNAn7GRZ4RXk3rB6YPA3Id1hapKO79Sfbs5hZkhTVzN020HIfeiET
FlyCpx7Qela7RNtvc8GmFPQ/UjqilVdW4/vZMGiKt5cjqTwz1Xm29Ie2fXq8QLj+
P6NTOut/S/k/FyFQCB3kaxvCxyOGugDLqF35uDA9ch5nagaUbUQCe71y4WG1vzs8
VFxmYTgma/UpqDf2HGehn1SuUiW73t8h333cXuzskxTdpbspwjQqaTiPSUuMLLa4
T1AYrGa4AVAbx4NK+ijyD4GwFJeXbWTch3VoVDC/pJ1kuugg6oIyIOHuf+vvrxIE
FzC7BgbUu3dqqNrPco1mIGFdTf/TRsEn+1IeSFrtRY4ijaRo0z20i/nIXE25SV+t
`protect END_PROTECTED
