`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
owWkEgoqHA8JZc0z3Rb13RuQRSzNCPe/CqaSNSlDj8/KCL9n26dY+21aQ+ePUCG0
FaXwupuWCHzJdN3m2M31hW1+enuL6OaUx419dQECkGPzEHffWFprYC9rd7tpJTgA
Ux/OGDxlWeHk3ryTQtaVRSsML1jrhFkjgA2bitCMuZOKIzuSQaXLCMWc/ngWB4a0
/oVcbj77qrh4Or1jSe3VTTPv6xYbvZSe+XoJVfFkhFi8VCIqLLOVV3DTY4L3ig5h
xiqbZDhV6BtDVtHYzf9NVAIB1JTJAGlHdbIjNQulQLxg47SwB1y309o1zJxEmQLo
Rw1ul5g+/qerI8nHIg3bczvnd9nCsQk6+I3zRH4mNf+LvcUJNU5kftJySZ6y9jjy
sgHC8miaalGTtHoyKpQIURXAGXcvnq7w7JAyJ07gG9FEa8oBMlhhlwnECDiVxXeP
AGrwpF9MyHDvx24EWwemsaz0gUlER7Nf71nF2EwEQoU=
`protect END_PROTECTED
