`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kyURtOemC/9s9zorNZBRgZsm7TtGWFUHV/H5dwoKevdkPDNZYhTgGQlWOxM/xWL1
331s1gPw9zX9P00C27lgFSKysP0z5APuaLD73o/NDZU6UYHJtBGOf8sxyWsPXUo3
oN9KvgBCsKrOcHB63gmzT6H6whgicMfyvobKQfJmFvVkIar3d41pkiYpxmQxJWaE
vYE9YsINRn6sYDNFRfZc46RO+hEog/eu4h07RTJUxuvzJQjWFNLVHUkpuI6VyTTb
mDeVNq8Z/ElM2fZ07xgNjNBR9o4sA/uHAB6lIsM7wNP6D5RV12iCnBxYGVl+0tYA
+0dFNbJu35WTKRZo/N25XNPaZofkSSluIVD230wTTPaax8ziiSVUwcKk+Xy2l+t3
EHWrOtXMezu5VdHKBWZ+fjUxZ5/gDC7N7P7QgzK1RhmVAIxkNArM2cIWZ00W+9Rj
lOEpNAUgpD4t4SXWbTaYP6TLY8xlf/Dsbur2RrYJz+0YontF4k7Z9rhqXTfgz4t3
auXwxKwiNKhw4EToWHz+dVhqojCuoUXvYRSVd+DzFiJ2vRxm1X1V2BDCwEFeCcer
y78NG9NQ/c81wvfO0Urdtdghc/FPRK+tOC4/7Jj4hTMk3V6fxHADm16yzmjNX2Hi
yscn1n0xxP3MREkJJnqH5m1WlNwXvKk8Kle1RV/TPIGk4MyfnQxWhaTK0FbhAnzc
951k0tOxJVczT3CHLP/5PHX8Gz803tzDw8bHu+hGvimJp2wGQhMWrb3tgmGrZSGl
Sikraa3IIDWyh6fdhNofcNd0p8ELOGMOiHeA/Ja8LayTG6FWL+74g9dkCLWAJ9Qq
mUFCjhsR7Npr2Ns84nH6obRkCxSEgh4TLCpVrz3pzpv95yadRm2vbfJRKQs3J5yv
XCy+OidiEYywXkkNMhbuR2fTiYPB1RlBd/Q5nISlcrVKdZQIEIZVn/PHsjDDLSFE
t1hm/k3IC0EqFdTl9XX2zeZAjr7P8R3vndz3AiT5it4f+xigE23X6/AK17OV7S4Q
KjtB7lH8RzKG0j0hX/eIj2cKu256Z4GStOmMHalz9BKX+yd0x72WmIhtzsTc81a5
qcEOIONbD7buPQoTPfAPI4mXR5j37Gw1mlAZpaaenNM4WXKVKNawt0zjKUDuBu5d
LcGsstDqptkZMyqn8qMM69KFV+RjJu+I+LJfYAzbapbGkGtlcfI5cl3TtpcZE/I6
RffwgFrJnuzp9X+NY/gGkIfrQe4ZPrb0kRbB9EsigvcItINLoxYkSZn/nDV/RDLV
8B5qDeuX4pSkr04tcY4NGEg9/H8quFFIRHNd6CjI6of5cyarpi8c5eyFXnyU5LtG
jJGbMpbLimdBs+08grvbg77Cb75KC5TFEEFMz5UvivM+9MTnZ4yem8ctUS//OdjE
rCjXgHnZ+q5VONvdniA3JHSvBnA++sFLbC0Gkri3M+XVdm6asnUo9DX9UaftwnX0
8fSgqI74aRXNfAASar0zoWb2oLU7+eKPtiVC38rDFg8WLsrAM8h1HARZKvsMWBst
WGhvdGuA+ukN2AS+v5jLcUHM53juQAHLK664YPW8b5nDRFBprdMmG834sOy2QCvQ
qb1BYGrFpgmlj/mS8+OBGWFZVd4jZvucUEheFVEGbCzflqP/nEUcCvksBFg57hhv
Op9V0TAICVHpmCycPtwlJXhDFYd6Mym7IDfwLuLdM63zEltvfXbo/NHbezvTtuNl
qibqAIoeBy3vOKVT1P8+hIY0WIT0mzUZNCtVtpE6euzo5/Mvw5AIkF4ppXtkGPbf
7HBQUpVAvgT17uH5AjL7VagYQwLwzH1NaxYI06Lm8VdGbzsh1Ni7GVx8ignUbTny
wGZZ27fluHp2L6Ax7n9VSTWpix8Z+nT70NvSGBkTRVT/THs5N3NPFjGJQ5barmrq
9Brg0Bqppvkm96oqDwVE9/CKz6sL0DSX6fnUcvOyucljWZjdVOeOBlQaHp1jhS9A
uEsW7l/U6bMeP0lddYf67CLKUtMFYsjIfJaLE25i7zpCHpJgiNBqf086jrbs66CP
CvkI45MVz4FUe4NbWNoy58v9kUd2gNQ5sWa/IAyyJGa3DcektHNCWVMnS61rPFxH
gFxUvsqc5JB1F1oAJpYXmUShT+jTET8Hrh2TDi8AnxBI0h5mS/i68TLxxCdGBSCH
Vo4dDXYICFlsmQqNFLV9Vku/9icZoycCdDqbKUrF9I9gBmFmPIakBzBnRrfuquMr
xGVGP9vjn5T4hiXYBy9XanZvYgwzaTxae9LxKXeBf2Hmxl6QUW02dEAvgm5a46yi
hCQj4SN4I1yEmSwX1E6JgP++cl+vkWQPIVdjdyxgH03b0MHBdRY8/HJuiMwd0b1b
6fnP7BWp75w5dVX99CwafYEEuAnyCQZz2eiRTHfmkdP5wRCuYA0nvGYdAURpqmD8
1hZT5Rt4TdVJgAYGjA5ZmvVLPU9U0vzneByf/gLvLTF1QjaF4Xxk/j9OhwwC1eGK
+TE/8KwOiLGkaV2JMSY3t+mVhACls7RiOWyXUiBujc3Lt5VaD65xo3qH0QOu500x
HqRUaD733PfJGrsgnBBP0duUFJB7IiKI6lp54uPsiM/ji7ipfsPuyEjWeYlRimUz
iQtZkZGr+vJXMISo9CEvo6r5vrSWUy+HX40xL/isweiorFaaQVqBPPuSDUwch4aM
Msxl3JBNrzxmuzLFweWW/BXCI0Zjh5FkOvwf67YFH88RN2sp0UYPE88pfwzr0yMN
FXylVHEh1DOtYobg3tmtAMnYpnXjS1YNFGMdWzt3pfNtCv3itSklrOQfCIUCe+Ll
tZNmbDjKYzPX5o8GzZjMW8cT+aFguofOsE0bRSzBn81dCmtCySYiUaM5VEEm5tjY
YTE7mOUGMyle9a8A3lSbjpjor0PDb343hW3OJQVstmCXXr323TSZ995DwLcH7UcD
sKhIlpPukYkGixzCfaesVXEfWDQ/wC2DlpIaeaScvcm6ReTN8MI95k7Xra9kyDll
V4VAAWNF01S4y+obl4Wh4XwDkXCOPq6IiP8q6GGWHlMWIiIP/Y+1hNSMbaOSRMmD
v9trj7Jv96VCamYx/o7EaBO/yJXAohZAWuaJjMsIYg5ap0/hEIHM8vOYzlGkTrGd
euQ6LmlD54ogGl4uX1Bc+HPi87K7cU2xjqFqzEnzn+wXPclfc17kjha6vxMvxjgI
TrbFPuKrmlkSepF1/lf7gUaZOMg2/hmxY6luI24f+thlwmaHluhF+CyjHgUFJd9G
+2Mssna+EPEWW3e+5mJ/hRXAH8f5W3CGvHmXEyFF5RO+CnuRinZIEiDNTZYRKM9K
p21elw0krwkvv5Gj+oBBiqUGu5xK4d569cLQAbKSdQVHDFvbb7NEZSCA8Kt5IDrw
u171V9F5VDUZLjWSWUZOSKHxd1eEvfvVx/8kpi38GakCxekZbp5Qs4o2nnJmAQxF
5jpEiAa0Ygznp2TToDeys25W0I+2knoZYXgmzqb2VZbjOBWCFOdk3cqEha7OMm2s
8VRK5FG416AoAUDyMPFM5G7gnSX8qJJfnfGX+giF1DarTHjV1LZEDLi6gq93IT4V
fiGDQ2M35nbH2JZ9yjtTURACBjorSLcMDmvfwJ0zJShqv6nGeeKMerKh9qhO1p8J
f70OUncfPWuJDuIFhFYgwrodrqm6WTbXI+LVgva9jg/02aNSt/t05Jz92ATfIdGp
PcebfGU+CaL9ZAtywIl/hyY5EDW42bZ6Dh4X7UlBCrIv4XT+9C3bWyunlB6r8GgQ
UosW+gWOBmXUsZ/dF4mtrlJ5U2smv1FgIcELDI6X8PhHi800xksuyw6/J5XF/1mX
gSLcB0cYxvu7zNgjZLKheqtuJCci/VcPupP9iI0/txuEkv7brtD6q5StMGGlgI3X
HvQM8eSEEmmXuBIiQ9gHlhwf4qdc1sJhAZtrPlijvdQP40nWLZYogz4bc2G9r8n9
ClQL06wlu7BtiiJRsGekxvvo9heMs5kTvDh+xjwP00RiWwH3s470cWjefiuZ7VL4
SLPSV0gG+Kt/iqYogY7QyAdXC5nn4aG0Ug1VmnAuxVKGk1tMzYoVuLIWVxVbrHVb
8pKQGgqpgb8lyAWd5ZGjSS+CdTyicItH9Z3olab+iqJvAqmoCL3rQpKppQLt/vKc
dLiNdHDDgZxdWoVyFX7KObrTMjXN4yKZUVlixQn6QqiiGqvdoO43WcElC3vQjZE1
kvUFck0sdyzQAemGKQ1cgwb98NBnxbSEcY7B4kDIeQlfXWk/IwqR5hH1KdqDp5Ik
IqBpCp7p8AZ6V/D4AfPQmLzoImA5gAdWDByd0ZxiwP8NKegXjauGPLdAuYsV38ra
A5tKpw6SkNaSjivV5ntDHwHAUv5/7Nw1rFq6PE51KnqwCVkxpfTF+QFGxoXull8L
tDlF2oyYL5DBj4gyK0oErGNNrDxqBRPNr2mNWemOg+vW28hoaPH+R2VxFq1D/JSN
7z8zwhk4Ck7hVF+whZA9RagbJmB8/g8e2fkPYteu1R4vH6X808dBYczgyxVEc/Uo
s0IbDcns2Y2rR4+IhhimthctSeH52SiaPME0fMcMuLveZKs8buWFb4V4PUuiei7v
+bCV8Vr+SHqohiUv9GD8yJWN2ryfjPmoayAP6ePU6q6Y9NvxHnxAOJPSNkXARmV/
UwNW8e+aAosw/ApX7dQG/Imusj9GnrlSHnbqhyCMzFokvBiTyRU/A8pqdEzzhbuc
QGL9VHiI4geIl2VWc5LXjfGnc933XnpaUAhI1r+yO4X15ANW4SXM7dCGoj4FTSDq
mDF2UCxo/opKe4PZoE4ch3NR/ZzkmW8GEUo5gmf2lDLTDrgREZGqYGZ7jmXe3P6l
cjM4aFzlsR6DtSR9SyOC7MqXKW42R0OTgbU+vyohk75/YAnozocpCkHGdr7mWSli
sikcI2m4JmFO5zIK5KZbs3y3zjCMxC6ayiDPPxZ9HA1T3GkT/Xo1Znyc+irNZLeq
RxH7s/3b+oI5sv5FFBhGh940T9C6Sy13kJXOtfuw5cdBwA1j2B3HgxaTd4etL7B1
mciglOJn29Kl/IoBsoSKOYz1pLsxODjuL0vd81rCvircMgqj1jzZOf6edLmwLeT9
gYoPLz2fDrX9BjWT5AhvZoXOuwUe1yIYj+tN6Yja/ex/78ia6kDfHJR//7xvUeZA
Z/F1PC9SWDxqyjSjr5irFs+hZqHo/kWav8sJ6zt//ukBKxInXkfvaz5Kx32PCvey
ChJtlgJRvGUs0bIloI5Kq0mPu2E2xPGECG1Db8y463OjxE5HFIi7JWRvr8ikhkJz
/mUFa6EI/OricHAsYdi1Rx3nVUJ2vsbL1g2GAkjJZopopVUbU0Ro1oR8/jXDbIfR
XTiEhtQWrOXuUFgR54+C58bsNaIh8WMEbSgkBl8ynwwzQ4Itr16QQEVX63b+9s6p
chP8V3FMNMJJdIrbV228R8KPom1JHQMyk3Gy693kPE1ufzxGJZc1k9tw7sih9Jhz
kcCzQfNGJtcSMh1cGXHymyW3bC1sZ4h2l9WOlhBIzgDq91csUIQaP18t4V33eg8+
7XuLBgmjJz94MuBbZaLTTy3B+FxaNNgrHO+pkoGQ6yyhnjz/eyKwsSu+nmPjykgK
/p621ZtbPYmpriEZxaJfvSAv0KAQ5Y4YR0m4QHsTNSWniixATmQJ/7ebrzz37WmE
B2voLwIt+hUcX0EemLK0CY8pAXDOAnf0CVlD3viqBLnnl0RDhx1hTC6l1ZvpMhST
WkYJ9P6dMphVKoxEV8IyQJ1KWUnycSNNiZNvvDaE0upBY2a5HOa7MOe6R2/5YxTN
jL5YMXVJZTgnyAubz9ZlHq3KpG58FfBs03c0+dq/SrQOaavt1HzWu4r4tqCIchK4
wRo0JnRPgZ1EzF1bJPtR8b6SkLOO8u7hGYf6UJ/QSJOfkH+GcfaN75PQWeTMrP8H
IvcPv8Z1gQ8SrqTBJKpMO+DnhE1mCEdoA2XM6J6hg8ALEhqmqclzOU1ggvFeYeNP
wgoEDiV+hMQJnzQQa0iWw61rBe0Az4fle/cavg+QkuoKp9y3o94bgs9C01g0rAAz
1FwkMsr6An1R8K/FYQrtpsW8gZHer5yPKvLKD8xXIVZmOWRuywfI8dlFLP1FlQgg
qgt3V16Ubr6PTkFZW0KRLxVxYnx5QdoitehlMQqA9Ji9ThrkKpdwbLXsS2+gbBfE
vwgBtllsV5oCUgkAb9eVyCToXml/7nT406Cm3n0tqjBu5lQfQIoI0/60kYbhbNVu
ftQCQKWAxuJN13ERxj+ZPXQ44+9D0kiriqFKaHtOVhH89g2Nsg26XD/nv470Er6w
GI2DhheKh4wVjJ0yVX7BbmEk5zzkm27mVIueh39+10k1PeKxr1Dyi+8g/MWvUyBa
ACtSDRGsB4DFs58+4RoBKzZAAkRZGr29gAS5w/1D5edTFmzi+fnO1A0Oq5kgbTld
5bGo0ZBbw78Fh6O25KiZpcWKalLZ3QB8HhEWt/d83n2SKpv2g8NsA5cX+P/zRbNE
M6fJtlg+6fIgU+wKgbKSsLdeZrdxmO9PFzX97v5Alp13uAiNmjUGe56nvDBrHLw/
vsNzfXWcTNbI5alhc30iEn4fjOxpb7b62DJYLct9TmxmqSeEkM5FGA/vQW2GwVaJ
3P69yPeyJFBPIJrtgjGel5uq+j8bIL6WWTRuVBIiMReskgRridPZlwoUzBta4oOG
/kmZglTJZjHFvitQyVCkNV1+TXxtFuhHWdzs4ReHhkszQddLuTMrp1cc5B3wrBHy
odfQMyNBGhzi0BgByALTym+FZ5uGCxTBXEu9C5DCWG5V4XXaXZxOwM8kIJ0ji2WK
CMDKYsxBBq+Jbdofq3sVogeqf8pYFGE0c5a+BUKcYSZiP+VXWMQ4icLvrbolbbSa
u9T4QTVDVKokeaqRZYwRi581Dk04q5YC0fp+w2I52TsonM3tUwTwd9cNbpcf2f96
dn7jq+YsX0GpDOFcpH42j/AunTAVg2R8I+PKHjIMcGqA6lDGpTw1dyl4+RD7+/yI
r6xe5NNz10pRX7KQP5jzXfDBfD4qeFURSo2Og2dWyE2/4OTobSeAEmAb/Y7Y5Tgg
CGGjQl+c64M3cZjKu4dfTWOHglN5DPC6ppfA/ESpB9FgfgpFXsseIRQkEObi7MFP
gVzUf0szOKsl4TSfhgefs6uXJhp9W8y83GVLkSjOm1Y3gp6dR3sZKniEp7suhL7U
YkyJHcgFRZDzHAa300KBSk2SFAPfFc7F5x751Oppt1ldWhWXTO/mOuZX+tqxaBtu
+OYJ+183u2fQWmys3Asv0P7/h7YlvIqZyEboF+P19W5o9CVd8352LYELXhK/UG5b
4gXtONeuN70RP5AhN3S4pShhrHCvWqpGjfV3yfDeUQXOMzft3fsJALH6Ozy8z2Fe
oEtWpoPp5e0m9UKjolnP7SYw3985LFxg6BSHWiAQEaLuplr8bTSKex5aDDepf10J
UrU59BOfewK1OYimBFGofQWcduLxWWAnXzFNHLEXi25elN4CF8nHvp1L0X4HPfy9
6YA/R5Y3p28hclH60dYij9vrL06fHP0Npt3ZgB3bqZe9k0M1KrtHtCXwUpfUq6u7
wrXC8rfH27ciotx9Xv/9JDE1QxOi9cwMOWjpZ6krdG+mdsUWVJ7gfPcrBax2ZG7v
3GiY1D0Yw96xl7Bqzgac2vNDPnK7nnD1C3hWqm5Ak5uROJEReVh0xNRAPu2WEV7K
TCqAjOgNCeCMpGLiUHX9y4sAwODjDbPn8UnC6aAQ3v/3PFsEdM5erB/ZLiAz1F03
JU1mhRD5bUzrZUlGma1iXk8vztXFD671v6jIzNSQ9r8cy4pQ/WrR0B0PyrIEJnuG
tsxXSafF1hiN+w0wN4VBILny2ESpXFpEEY2ckfOcY8WozBoO4zem+pyOvlfNkV4v
xbkljRm4z/dJ0k8ee7aK0cR/HJpc68rd0u5ZxisUOzHSRo8SjsNJHIkKD3GoRQ9k
rpfYnE3VoL2tbIxrdTgEgyF5rmaLGkuXyAYBtzG0DrYKn5ntK3MJXpJtpgTHPggm
32J41akSC1PE1BMw1eC6iYO/dkxoVlhvQHdlrJ5zloXmjdmiAnq0Rc2lwCxBh74H
cP5Pf5UqfCSOqDv+9a2X16O6W2Zbbn3p0UW0vCg46winHz1Mom4kUj3ClD9wJLAa
oosxWlQUojPYCXD6rPgCrt6MAe+WOESd3XHerfUiMgpt2ZjkZV9YlMBKjeaF5yg1
z5vhCfNpLqPAyefe6muyrO62zJv3RIUo5m3e5qAKjjl8lx+j/QPLJ5hItSWLQFVt
qf31xMwQ7cAkRfJQBr0Oszjs2Ah9Rpt4bGBVDz7qZQ+x1G/eBsK98sn1+sd0M42W
uIHDHk9BT9B520hckfqV8Mkv0oxE8rO8X8SYsv14cm+Z6RYJkNAwHqVN4wkZEi6j
zJ+bAanrGKCwg37dnRYhUqzQ+M6S8M0NPrgCzYeXa/nkdrfwbD8PsZpxApZWcd3l
iDKGX5D4vNdbmcYbANhLp/RnbPXCPJ05uv0IHOW32TTqmIBzJZ/dwSLg85ud8mLX
3sTOzSFzNfK3KAQSrMnWPseRseasRamvVvazMuTWpvXH82/E3voAxgJGVqWImEl/
UzwsXUpPHGrAQV+8A8XgDCiExZ0RO+M8jqkKMXsiKuB+UsFXI6/Nend+jn6MRaH4
lCFSNygBWLF2ydymqFAcRIoqjgnMWNQ3dUJlVU5dMNjYoO2iN+l/oeItmdge3pMl
/7AAFyZAqxSSRQ+oPUx3UpC3k1c5eZiqmhgqSuDUaVGLtW80kg8kY0sNREw4GOi1
4jiwaB8cLhybdd6IoxcpyZ8LzDVzn1HQeuc1KOjXRYqIGMirnqojLLekYbW+aqF7
0BHQPBPy9Au7QUjDwf/iUl9yI9E1Sp1SEgO5+hjjnDtHLpGWWdNwaPujuTi7Wy9K
3Yv5s64FQdiOW0W2yKvl+DgBbEYGJG0a8gHMj7SckiBIMCbx1bTdaH8lXvcYBpOv
Va6fX7E0TCuk9xJZt9rBoJ5JWHqWF5mngSQ/DnEI9e850mgPWg5OKwAV9uUo3qRz
E2i4RWOEItGBby1GozZrKkPB9CjDr8sBLcKJxWTzmdafm0Vpv8Z/yRLnquYr3PGJ
fMohPeUwU5SIupM5TVxczT3lVuhU72a2WKDsxvLyi1eYgRGerPUJshgQPWysCrZ4
SHCgCebNKAPhrmUfDI9421HB1xKXAfqvXWKKCZrQu9gXR9tJVtrZL8WV+rSk3kzH
HXc754ZgSuRnZHg+ZOnCrloAxGxcpoE3PqwrTEXQNhvX7s9NFP6QablTvbqjDIDc
nKmdkmVdPA5nSDnZavd+54cnMElVUVVGB/9r/GtaFxZUNLghO5+qa5bvJWZObQOf
/7xFliu+GlujDH096sqONv187D7rfsRFl6Xo77HKC+R8Dh32a7SQgzEKnSAnAwgU
iVWU6hMzZbhzKyoJD/bJ5BuSZYrHRrIEU+4YjTNQ5CLqgNHIbwv3fML/oAzekqh9
Ca6C3fhsihXNIfPHAYqunq17nj+/lY7cZRV9Q1o0KPdSrhBRuNAsOuJ2544Ie0EQ
JjBVh4d1M62KG72vydR4sdRtM2885aDrq133mo/WDErh8+P2wL98k5iMJeTNy15p
ROc8k+nykQ7RfSU6LYs6jXaSXgsHtoaqdp1uwGFYv4rFLpuE/pi/JzzaMoP5ssrD
ed0uVwYGcO/IF27LM/d7D/UXG474XNb4KBJ01gx4HKlOHq+7ntVDx4wnt7paOrqV
NQdO0JsxrneyUpBT5NrNHZSKTrg4JveOtWxtvigDjx1hu0oT37xahgJJokuxw97I
1jJmtQpl5P/WiL37+G4EYZRa7O3/FTwEuiGpXYSlSI1OqeXrV/t+h0MsfBxA243+
5GI+UtWyhE30HwOTlJFOwlkND6hFiumgLJCRUSVFB8ptgwqM3TGjo2f8eKUzBrOB
T4ePd6HxglAvGejBfQ/X4HgUfjsCr/9S203xUkZbLDKU39WpbHrHe+Ag5CDLtvVC
H09zfW3S7E58zWkM2s706EsbbpMvx/9WZR1AKHoHZFXg0yITYqx3CDjEZs7+OnAY
h7kAYc9lJtypj1ANZ2aCwkWUDA2xDAtD4X/vs/5ZvX9LZn7QqDLtzboSVwi2+K+B
5EnVCfA6QcRUEfgaw52W556g2XDhhGgPntrbwcMt6qLPBx2xpjlegmBeuJJ6rZv5
XYSAs0scO/Upm0RN/9iVT6HU11KVhQTF75AtB8JYpkIaT/eR4mvUMCwyGaG8g2td
14Si9KcDvTxtq4l3FUq1nLTi7DeAEX/4UGtQQbroxWQ33RkCDFrWpSDsaA9yrCHI
AgV50aP46q1MGJ/iF9YTWg==
`protect END_PROTECTED
