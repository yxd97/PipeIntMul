`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+w7rmpjWvuEszGjKKDlAS75Fcwc/3ykWrZqytX7wmFCrGI2JDk5fd9Z8Ai9mPL3U
ykU0w+zI10XtsQA7guA8EdX5yh/YpYQSrkiaNUXxI6QTVAVKTbz5PB5RP/j9SLAM
t/lsZ+8D+eKoBuYHZzWZ38df8h/8VVNBnyiV9fqCiVEL6+Y5CSfkyZj+VnQW1Maz
qkUw068aZ7xEgInFgKoHKA0FlaTADA8l+Bg4QHyoURvrTJs18kodqo7eITaHZgur
IfkjmTsq22QOr+/LBpUQ5SpQYfqsdWWB4pNydmOFXpsgSGqHozGJbKpbPRLc582J
xTTxjJ+9Iz1wAw8pj4e6Q+FGdQyudO7C3GEtSZKcVy7YQvTVqhIhL+UZDxQ2KoJ5
1/Gd0Gou6MPGJqkUKzrwwtz6er/FEGrWvMjmhAl4G5fiOfmbOYGr51xf5W0aFpbK
N4UpVE/nqNoAzeiPVLZ25wU2DWmalOWRu8NV3jR2hPAaxjXn0Q0H8Q4SnmEChqzx
/6DemQzylz53jB8jAKGvRg==
`protect END_PROTECTED
