`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LAOmR1i9tcSATOqLXoz48yL+TPMzLUYsh8vJBXRhnTnNrc2nnIWmDMpPja8Q/d88
Jx6RxGK16mPllRh/9yiv3I7qd5/HITKR72z+Csxj9dWOjIRALblT3eIJ901iN+XG
o9KdBpjeixnK6616fUaWkDou5yFf/cHYt94z3RCInvkz4uYkkdWaGUpkYL/IhiOj
VhHllATm/UDlGXZtzzatHUbNsCxa8ecq/aRRQ+lWKPHPtuM+5FT2N3Q1Fh4f4Rk6
935k+BXmiPYaKIXS8SlMXP9oZdAe0L3XYzimtMx4xYV9Mv3k/ifyfZ8Pghi0aLtm
kMZ8HdSEBz+ItGOJZDYQAkDptVuAfHr56FI5xjllpXHztJ1CVLgYXFna3aAlKpwT
X23orwzyTy6tWjyPzRsTnZgGmUl0vhjFNcI7gyMz+pDSHrDskRDswP7EPTiWUs7z
O4e8yt+rjmiDu/2Q/gmaNdWXga6DA25Q7QMsSMHfnSmH6OoQP2QyxwKArr1ztTxf
w4+mX7ZjAcfvgAKp9vQ3Jb6lWe6DtBfn38o/COv+0w5IQOjx/4301rAz5o1/wAsj
14h4ZSyiZRhMqKPM3QX0Jw==
`protect END_PROTECTED
