`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CiyQBTJIM15P+kVJsd00UW+Hc/dm1rKI4p9m6LmV/FW8Qs4uUsKN3el7rzImeaj
tn9ncsNO5ZqwfujIBOYLJ0aPAM/hStQUGeLLDbxRYOC0tgRKj390RhW5epwiB7Qs
sHk1Ia6mvFhw3JIl1DO7zxIysu1NSMwqXykFLJLw+TQzKuLZzSJ2kS+vf8pSTCkh
fmQ24KOMgxirtd2Uok08hPyvMS/fg4PIq9d01dLWW8/jCjckWlCZ0Nm+CMTQni9r
erwwCMLKTXnj3E9gHyy/jm6YjrNGDCmeVLH2lFyrzPfwvQHwC4WwLG3cUfMCd88Y
yWVGK9WwzfrMXyQU04aHig2JD11VnKC7jaUjN7tL6tFXjWBAOcWt1LFH2ViW7GWn
1HN59Tf/rPQgpFiIJ+LscI32l8EBjQPvwipSItcswkX3XkACUqF8Ufo/DF4jzLH5
gkdhRBpIVaP3RQX1lzqhI66Qq89MBmrna3Ng+q8LQUBJkeygjNL+Abe7JKvWrGk5
zddkIe+1hb0CScGcVIQ6jidBAyLijI41pbGgOGjJ4Z4bWkcYDRL1K0XUyKEFt+pU
S7vX5x2I8uOHblUCsOMlU0iVME9QI2pkM/9gTWkqsGnn+dtyMmtKqAZ5tBRJ2sS5
kTuUTUhUCguWMCbWbED0vWRDIV/wXuKTO3gpnNoeCHNDY+H3XctCyAfmq1yEvHP0
Olv+Fy7/LLmEnwB7aYzmmZzX5OVOeNf4tz7w8gO58rvfB/EmIfzGzl5Ogz27C2Sk
00EMYE9vtf1l04tv7+lCtg==
`protect END_PROTECTED
