`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mfp+NUrwr9NyMM38J7fxDtaFPVwz/F/shgrIly5XpSDjLw/HYnAuKOnpa6bTXYvz
1RFaA7GsKwsCHPW4dnoN17g7XwToUghYtu2jJ3UyOOa8uKUtEBTWJKZOyDpfUW52
RdEX1k+hrwk7sr8I0OQrEJt7tkgHwyoJQnxWhit+citDeff3cBlBxgsqac7UfdJ7
z6IEz+qyyj55By2DMiCYNQqmeOQqhpOR6ntJsXDinwLT/yMQCIh1olhMagnfjNkr
ko/7UQ+TPLTQQrdjOA3XXt8DVf2PQJ4oC1e1bIh3VO9RheOd7TK2+AKNKQQechZQ
BGGCQjEjNTNyb6X7chQFqQ==
`protect END_PROTECTED
