`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IW2B87DCmnlxvtbOvvV7T4DRWFnxGy6xomcy4gbkDZMkoVSumJnmw2UJy0Nygqj/
a/ZmRdEUNlH4ddkr4a1tOS0UpcXwjFkFIjIwfBhBCH/b9aRQJLJEwKTizc0dx1bq
Pmy0OMKdl/rPMdRPWEtH+oH7fGK8nTctAGAUFAPiYnNIsMgpa43xk/9EDLMTvQnk
9Emck33DcQ4PfCG9Obbb2ci7RYK31zOva9PF/NhkA3n43a69fbWpSBxNmMDaQbIY
EP4Vj+kESyyx9zG+WCYyFAkuCj/vOjY46ZzH/jOoWSpJnKB1hPDxscSuy9kOo91Z
AtZV/rP+cveXHbQwcDGmxxsqt1tRlLrAiKkXoU64Z4Y8BgDO/8y/+C/ySkn9bZoC
GCOvRT/H9JvMvONid8a0aynoTj6tLm1PCvvrV49kuNHlk4zL0t1ZBeGb+pwwOd5/
Nf5tED4TW+EfUlom9U1hzhKR8HvxBLBl+vE2FXaSwDEGgpiPsmjeBhQ+iZTnGh6u
NgD09cFRGBuvPUIZ9scnr2xxL61/iEDOPZVa08ZCtTcp/V2lVIM60iN7WX2l1AMI
LlmnqOueEWa07Ib8GDOo7DadaJzlUUPWszrJw+XkT8kEKIaM/c6Lg2/m4l9qSFeO
5dOGQhITGzR+pmw7eGxm319EghKNqWQ2PNqzPzN1cas+SGnOSo5Vfok3sUHZUuqW
8Z0L9eANqxUcHYc2t927MCxslauciQ95eprgpChLKK8HCOagSXe50Ma9ctM6AAp3
l+JCXORapC+JgaaSqecwnN6LGK2Fmu2LoKFjnrgYBcGxXowMPfrdeOIK1xQLVld8
FeurUHYJhREBTXluyQ1kBbMUdGhArCCO5b7tuOwNGNbt6k4IwB4U/x7fJdcPxH4v
Z5PGs+oXlHW4i1CJ8DjI/OProU5BgYjoCgyLuM3EGlDw7NgK0er51zFTdajAKdIO
WUgubuFjU04d2qK8LCLkIaCXbQoDon1EGyeJCQ6sHLkx4KyITMd6LUBgVB6LxxWt
QNrMoQPVyaKj97lXecRcryEsjqFvz3xUaPPoYP9Cb0fsPXIOzRYTzkN5FHmxMhL1
ktvv5XLeCjA1J3dVNgr/wdBI5kjDLxV3sbxTvkH1hrqeailzVaTavHpXNoqQNwwM
bNvX43RTHLhfNYL59ytg7KIeXmm5Yz3FeeBLEIw7i71XJj8lf/Xl3DXa8Z3qI6b6
Kk8D9Ude4K6ILFD2DghcK997F4xOLsGKEaW2aYRsPO/NTrQJunEnof1o1aXiFuii
E5lX7Ha012ImEt6faDsnaQrbh1/XK56rvpfqrsLCeKhJ9J4DtwoYsoBdX904xTfl
W2LPsAp1gAth2MuC97t5Sg66aFF883J/xP38vkfC/fP6qEFPvWNI2LfKIbMFmrYb
eY71VBkbH6gClNmOkRfCfkVZBq2ZGhotY1CpK+ebN8hsUXH+He6YbUgJISnkep1c
mepANE18crHsoAXqfW+fX+nri4cFcs3h9/W7q0UJN0uToRihm7cTYDbqQoOGOWMX
/J44c2185+MByjb6xn7qc3Za7VkiSWuOwb01WuNC93sFS6s/a1upfbDn7TMjlY9D
ca07fJ7vG8+1HhxORiT1loAk6RQ9j7FU2TcEtmvCT5xsx7FpZD38q3rDFNvKTpl0
M43DSrprE1sV8oGg+9+kWD3xMVsmC9RSu/XYRSv/grfUnYXuMUal0Xq+yx8h3QNi
oY5P5RPDZGsp2DbKTcMylCAKoSyj13jGcecKhs/+dnKSJPS+uJg3+C5dqKQuvWb4
mUOip9mHSnnrnnPtK4/twfG9SIsNUAD5/FLMA3l3BzfWgD93X/2MgRfJdGs6nIU7
fWRlUujufZaOzPPMLhIqbpOpTnWrWPtka35dKSLKDrWScOYKGCcWqUliOkpad4Z5
n3xRIPZ7o98OR5OwckvLudKTCLJJux0IG59b1plKCSbgcQGAuDnGUBGs+gwgNaIs
IudfAPlHvciJSiYJoOOiFbCR6Mk2RfkyYT53lZ6yZpxdllZTQgZJu/aP2gzAU2G0
gIcd7vK5IO0Pdriu+LYIY1l9VEBwyRCwp0MUllJ7pzYUOCYHedyDTwv0Ka+S/VNp
VNjlBp5BiH43E/19EHX7IpL5vEi40JsmpTMVfh8Y03GQvg/81vL1anumAnikGGFq
/wsgkiNOm+VXUY9wGzxyU7rpPSYSWZtn1nTD/N1KfLo5wpPNY2n9PIrAPi+QBGZ6
OMnAy3D9nsjWB1m3+CbJ/evppgHg1GsWClXQ139/GO5JNUqmCw0odP/tO/7mYHbH
oahqSH+5WhXBkoteOmg5oHAQ+1ibdUl+0f71Dj2dfxek25AkPmztkGmhYYsm1qZr
mQk3B5tkU4shIf540H6GrmStGh6krHyhhGbxpSHVjFkqnXxiHM9RcaynZxy+1vt2
3a/FInLU+jcrpqpDeesy4f33clE/U/XToVZep6bXxm4atiOhPXdeiOAGHGfiFNDS
v7OBQc8H39b0JP0tHHDp14x+BXdG91HMtsryLqeVOhDcZc7uGu7YnZkO8zD6zDp0
wXmupVzW8SloQhv7flZpxgopV+xdqa+9mCTnEgcUpRfF8EQjO9gc2Aplxf2lvC4r
4SMs4Bt/37bSYKrkCtSOPY404FHTtpPKYyjmuQA4bzI/uV/p7FDjVL0yG7VXk7Zw
Da60Hd2CkttOoPfk30A39WEF0UD7xEgzKZAY2pw+0+ov7q7/kme5oicaBF/i7ycx
TTOup02cRYtF67r2PAxRDEB+6TqgwRKH5IXtfe0WV4EV+BUNjCyiY79YVA7XBKKQ
XWwUlt3nQYNVsESxh73MJtReIbGBz4Gd10XpqQPgtLShrs+T5fuufJZCkdr5Tp7J
RiKiHbdU6HaBiAMxtJAs9ZJDab2YWUR3dqB0GkVLcg3s/2HJRQZDVJ4ceccGHthc
reGf5ME779QxB/yqtm/XujOVH2rBk36Ml4G90Nx9mw7P88gSb/nk3N6fLnVuEoY3
hAQa9nRUs+8yIGYdZKUmmGXT7jB+GB6ddjzaqp5MmjKuMw3k955/iK9RlBBZmEC8
E08mXue4FsFh3Wmkl65tCHCKPqIq+WwFC9E1vjsoWI1Gz1pJKQFEZHgEEIBoWQob
gcmjoghF/2xd0sjNDgymdEDmRdry5gm7Ng+xR4Dmo8kIG0xiP4x/L9cqEo9IdmIY
G23u9wgqLtKMmpLUM0Lu6yvwzmk7CmPkWx+bcQh4zvc=
`protect END_PROTECTED
