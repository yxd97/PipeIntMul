`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oS3Uh6TceRd0FcICQyW32rI8SlD3/V6gfcvJ1Yw7M3Lat2BApNBaXEkdsyu889oJ
f5WSNNCrkAl0z7Kn/9BrOoTRO4oE+3Z0e1jHd770w6//RDTCuFrMC4obLHspDRvR
MnyFDfJBmWQlw7nLljba89f2dN5gMjKEQnA1r3YbsJSwNcYisYb2lHs/JFOaXv/x
zQ0L5bexS6q1Ch+OzqisngdcPsiDsbXYXIekPKDRhdXkgdJYNNqc5BbFg9VDXKx7
38hIJMnQ/DBBqAYxohc9Kye7IYkdzDWtkbG25FP02MZtndmjPUNZyZ8X9IyxsA7z
oFw9m1DH4VrENi6+0VLaw8s33b9Zgt8uqR+3z8KH9mtv0DvpXQAufCnVVqdX/BG7
/YzMq4RU0giguVqhFXxe1Mn2361hm0vZbe7/UqR9vyzrYAJ8Huq53f9Xmtlzy62V
`protect END_PROTECTED
