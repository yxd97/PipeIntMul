`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2qn22w2MHlMbme3AHODqd8g06/P9AMf1n6z4TSACeTjdiL7QzN/Bk7zM4Oj7lu+
uJJe3gAkDnQ66NoMWwTZAPg8uhAloyBkUzvP2KUaEY0ejIHpXlWc5tmOIHIhvl0m
7WUKUGPLJpk7OMqj5ujaaZSdLl7fA4wLOlxzJWA4Pk5t1y9GaY7aHpo8DRr3Bo8I
13w2Iu687aeYicuGX1gbIpfRNDtNtfop7Vzp3SKkuE61MGiIXFREGeDTGFK9qOfk
XT2RBKHtZein3QV9c6cHeZUiFKfMonuAFmoY7i14PxT3YG3DmGkLSbauks5vsJn4
LWn6zgEtywjlfoABDkktunP5AwvNC9C0MWeqOrDXuamoG3XlmBpmFAdpDhfNxILh
ryBDcESoHBFyGk85TsVO5yRPMr2j5GwPpAB3qRkIx53En2cckmk6J453EPhU7MPX
TyXyJiw0hp+Whbj+cwPURXBucIEDhdbpn6myXFnS4yDgr66A1IDjaiTR6jrCT7w0
nRe6505r0IZ55zl8Qb01N4x8qUS48H6r5Irl9Kup3ry0lTmE4+HHCrDAjyOQWzLR
cUNXXfycFUwvMzjJA01uyF/Lfsr9HQU32QlLfu+iGsw4Ph78uheNOB4OpP83ue3F
uyZ3MSDQffYbL/n1V3BorBvW8MVGFQunyB1mV5eiuZ2czcWaGvb375qwDFIq+ZPK
nk2k2MZrfXwiHDlqoxEId8Nr5j6tewHN4Qxd9EX68GxFyFcJeTiGQpdaX1pcTAyh
JbLgKV9P6OkYf7SfH37PJJ5FhFhDzra/APedonRWLir5lPRfU9ICJQSY8TWFDmSX
QuPv//frM61eALHMs+ZKqjzk9QmSBYpKIAgT6gvC6ITtg8tzni4Ys2ozBOvAZszW
QkuHOZiEhbSsizfy3MYAv23b9+7USLKnMvbKy7wx5vLlCNQyd1GdbHuqGBW36Zja
VTJkMUEQY8MfWWcaIUi0hQfAUbMcFQE6Z1GiEgMwXC/vd1Ntax+3xtaEVMpdNlOI
fRcisfEAqhOnHqh01BmS4wqbB11Eil23GYCUoFcMaT44AfYvp1JUBaLV3NNczaRQ
JiSn+sdcf1CRXY8rfghbSS9G4Gpp92HSV/ollrqgH/J0/1p04nAsd0DRVqSd49pc
CcpSBT/sTVFqM6z+mYyR5/+tXj8op4OVUW5kiCSHkKmc4NgODXu/qYxepCnMZwIB
H310KQIc+m629fGgRIqI4B00XM7iYoDrApgKPI32RN2/gG6gKE48LXveK/onO52c
`protect END_PROTECTED
