`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
leRWKu3FC8sqzM4rulaQH6ABXzp15H0rrdEFENeIefarXr335dq1ngR6k3kbp3sf
YO5dj+/qco7gxhhlTEIAIZeDTLn1xGccswiyEQTJKKleh+wN4DCPGS2sXGw1uBSC
n8Qdf57ic9/PkdSwJZQ42TdwisP8y+UyMKUJwkpwtdeDy7IKA/NfE59/ponIFQWk
8GaaEczJKqAjAcljNI1otVA0giIAKiaQlgMJDs7Zoo5dRWXcJQ59XsZ2QMAWgVeg
sAPdfJHcaZpL/xYIt2/KecB8bLq75OXYxelqlnNuLCZpa6/EyC512xFsXMfjlgyG
Jr+SHYhA+0/75PvqsXw/eqIYrrFV0Pfj6zeWXBPr+ye/PaOYX/h4ELL+yZcD1idI
vLfpGi5MdMQ8Fso8LkCBj05EQBhjAkLfWBoaFjf0pLgDChG3h8knoQ8QoFXfhN4M
SqMQNqppAARRjZ//PM1qRK6olwmrHF+T1L0jPWOoChGCQJGzUfd4vWD7R+lsuoSt
`protect END_PROTECTED
