`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lpH1AHbCybX2gUprvcvtiBLYilDCqhRHpgb/+SCh9Cj0+ZQNwgbdPhHz95cz1flq
ivm4PMdbeNJXi0wTpNvL4NytKGdh7YnWa8Q0BFKvN/L2SZRHrtWFT8zwhwlYBAIR
y6THAOxHqAJaU26aXv5XyzFTDfoX71FfRhHDoMPGMWa1WeAHnKzt4gG+ZXn8DWqX
HhtD76BMFvhCpsXGA0x3GymX4HXnCpJxW9EW4Atp7YTckQnjoya/FcHcOk6uUp7f
gx0+EiyC8a/C0Npo8qUnXZCDcxwKnTwF9aitGWekyYCl125fwKQcErQ2uaLAyIgO
dNNdDkEnjeMtMCHi/nCALAbtutnYzddcl4NYi8pS3YpulJOhHyXxA7kXajUAf50B
rhqdW62xBsOcljFJKrXu+oNQoEK/okn8/L55mcAHNTlI6ergfbAIDu40qlzUOwha
YK9LjsONIMpM4CtTA2FVRMl0zfgJQv4X9bmQI3fi10njQ8S+aPHI8PxDQLZbWgGD
ez32qo6bamSD/YNxcw8eYtLN2iGdC/jhVgBNapWMYLwU5UoytHYooUykpCJ87APA
uTPYLgFy559/fRHJXpxbEawrb0b+yp0I4Y2CIoedEYm/bmal/B27hkp/w3j7c6Zt
g383kNCVcnVGsOKfuqTkqDG/wAhN3YlaaWriUvhqInng0Nnrt/jFPXXks2JXHgP3
971UnpzvBvehEysRXOxCYo5zJE/Vog6iFfmX7QJcNZ+zxZ/jkOIXE/Q0+vG0LCqG
fpYgLOaqEIyB0ylV3n/P3jsbwtGy3FF+uYUN8oMrAdtif1y7qlMy4KqZrYiXv1Kl
XN2gGaNw2y1FSweAHUJSDKiiurQ8p6FKNzYSU0XGf/QBA3Azgyqln3bxnG3MxSKF
RJmlKOrZTsHyy0xJFSc3JBBFQ/f80C1xHNN7gODM0537Leh+efHpblpcYZx2zzMx
HbmNqH1AWXneX7IGKheDEnOcfRIB1MRtjjPShHFaOoTTU/1iWk8oCV/5WUuMc61u
lPT6tGJZ580X90g5S1WV9HNYX91IZ4UeU5mzu/YUtmtuHEorRBd0kO+i5Y7HAexo
ZYl7Y+6cIJ14n62vDPCGAHCDZ5lng//Yo6/hFX6RCGCJWLWdejRJOJssnHW2BXjQ
8CzPkeVjNcLrVB7Y+PwuD2aSl5QnsfVyvSZnMZWTZkusEcmPADVAN16Yar2RQIHk
hyHVbjvU324BmsQvyb55NhTNdz0LSHki6KrXi+oWQUwNsz1228PeDcJTdOL6D8LG
mbyfp2o9aIHKfxZnQ8rJdiP7SVeN7EIR3QSEg+V+oKsuebYdKsonxn1bJ7WKuZQg
YrY/y0xmGG2UMztUOXCka+Stxc6cmLFp7p3n7LKZoGgWaAUh8qt7wHoxamZqvWgW
q3dQeI0HqL/+gLXYxbNKdzUJ/Zr7mTxaSNe7xtJMQ20oRuxfQjU8HdyUwtfaY68A
6wXBQa3cC9lb159w8idCKkIzjUeitJTMuiyH/Q+lhSvB4lDdf+gjx3KkBL7k4Jye
QtiAixGoIszsfFpTd4I35EdD7jVF3DKpnqVLDHUDNo0TZ1yVx/vgjgOnio6KA83N
aVqAQcJkRdBrEemktLCGMSwz77JFg6L1RaA8RXu+JdIjGWWcQZ0iKlRevr8JUG8c
PEO27Bi+6EbJoa6u31PZRQTZGcoWVgIa+/QyMWXvkfDLb8MjEcyigGXoSO1NSy2z
lEr4OxJD6jPWijE/+L858j/ry87czPVYLTQrr4PLGOi+ucvFu60KIprHcwSHlkQZ
Po75Ay66z8+j8haFCXkJzXw/vWswtTXDzlyuJI9C1IcqSc/qZuYtCDp/J08erc7H
Lo0riipzz9Y7Et/cr6OxL4DET9Fw8UqtyaCUyVX3YhGL3KZQY6YwvJv45cf2RV9y
4k5REOhcHK5aDprAkpf8Nw10UEg3LpvmDikfSwLaNCm8QlyjcAvfOgoFDW7zjib1
uTw840Gj51h96XPraZRBl/EqeEfw1c31bAztoSET3UKb5TON6F7dIMF5mxt0R5ip
Y5ekC2FC34chRIA+4M9QRE3TqltRwdBu+RTafaNfVoMqjdSEgBt8NJTupb45I08H
Tc1xbat4TuvhkB0lV1koP2U5rtpocWhS5qibGseeKrZTRLvR8rS1JzUVh3/GAAnS
ztESN+iItPtA3tg/RNXuxGoIBmWWqC+dDymWBDADyl8852MELXWkOzVv7qgX9p4v
Mt1/sWFoBgFKqRgDsVw7HPrK4utkYUf0scgnjKII1we242ysYofnpMLaIFdLlrGd
nP9Feo0LUvSqOB6Z1j1cRSpRH78rG3Ob5bCuxhJXFdTlsPSxz+CVADDApd6ak7ol
m7RGwBg82SjY2uho2HdyOt2Qr6JaIKcxkaKlz7ghWQ8E2sGblj6wQGzWKVWct8t+
bB1Vq0c9aDesfioWQxoKgwpw8hPmWqkdlp+ZTXcu0j6GTBvZcPtKeav8+LrMzXHK
RniTGHuyAaFbdPabGPtvNwfy/ymVnqJR1G/Yw9cCsT5AzTd3xZaiX4Lg7m8FiRwc
5mK/xY+zM3Roc5ecYDxKmv+zX9ybOBDPHxO5Xc1HMzZQVo9TeR3/Q8cUyXY0uh6S
sP2p3NrFHE0mUWsyKwsEvVnW5HuDzJ6odbftF8RpDyJ8B82oRXgG4M92MzoKhWq6
F9zZYCenkCnhv4958wn9ytTL9XkGUiT1RY4hkBlp5HsMcnLYHDGTHw6y8fUgNUq3
kKnOImgRP0nksj/mDROpbgYPweGl5t040CWJyfp1CK48pysSs5BdSkoucgIkAdj3
ZzzQ5P6qpp+uUa0+5hDo/iFxT9sLcsWBPt0s5/pDw6agESd8sogRJzK+HDUe7ciI
1WTJ9SwHVQuTszu8Gjm2eUueU5Hps/u5LZ6jFNVNCi2k8veqBenAg7g6DQc1Df6c
X2NaUO5dk2KJIQfwt+Ha0leSyOBVGm+k8Ml5elLuKGEUovaYF2MHHqDyr7FjByfU
ToIMM+Nn8QLTa7vJoo+DKcqm9S9QMO7pfhb6G/EyECCBZgFmEdK5Qif5FHskeYf0
067nmUgpmi0zsipzWFLtb034feabziGV+wbv8Q9MEiI0ZofYgTDIV1RGCBzOGt4k
MRr2bJ3trdB8ypR64I9qEw==
`protect END_PROTECTED
