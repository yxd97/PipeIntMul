`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ex5KdmRMO6RzN42wlwASacsVYL9FxnHWXdouaJ9HPgzFlXbt47gI9R4TlpONZEgg
Eztd+2iuTpSmcibQSrOAjVi95I7yXduM5krN8qQfr36OpEWZBq4GoZ+q1H30JIwH
sOYMHkVyUWcUKteWIQFkgn5krL8rh6mPSuR3PDiKR/jyDZcyD+/Qx6d9SbST6U1P
bzLYLu4BtSguoCnqT8JaaYV09nsGfnFTxEDhwYzOUPILW5ydJuUl2xdp2BK2KtrE
4wP5wUwPC1jYORly3NEs1O6q6ZM50bOIsqWd6IpUqhRy9C5ekSWSHmCvNK1rSq70
Q89heeujv4Cq9gY5Q0K69gES1MTUxDeKeMXnwpb0ZECV/EaN6T/sHjj9V/ewhvbJ
CQAZ8Pf/I4HHzwMkvvB3dQ==
`protect END_PROTECTED
