`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGGY21ff7zJ/BMQTZpgeyk5IA1RK/mij3X4C5yofRYy+zlHgVlG5sx81Qrw0QtiK
D28Qaons0mAg0vUM2vik4/6+04U37Wsstj6q4bucZ1J/xFCBLtiuSlbBeST6iy5Q
ZR7aF0FGtiidduqjUNXlzedC21R7HSwSRPb04Mz/02feVt2w5/ADGBkqNVpFRuNc
P68Mc2TXP5zIYKYPA0rvs6YbLFk6/0xgmWwR9wpUx8Bd+tgP7Y73MVauxVkYK0YB
NKmmMd6ft/x8mvMldjY9q6Gwj4Y2QnhclJ0kGb/HiFVVgLyUo6no5Oji0PpKn9Su
iI3IUgVu2fzPIZFtCWjEXJRFCN0Rgilo0+Gg6L+Y2rL2AQPtZTZRqjZkgwKi94+N
6cjOhtctuddWKbVvep6lZQ==
`protect END_PROTECTED
