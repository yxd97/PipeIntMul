`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+/JrAF47ZbOyI0w7QEF/OltGZROXnsZrSqXDGYPLgQHuJzfa8bbXF3jmy4ppW0An
hC9YGrPosN5sgb+6y4IDv3OndyDOvpNVv2eBjh+CO9PNbj+qw1J/8Yz4qlpcwA9L
TOpf8LolAKaaT3sBn/CJ6aQwKzEYFHnwUEbWRLWlRagGUdlUm6o2rKHIS1x8/WKs
ZbbYzvT5E0PJDoN9Q95tr0mKQPySr3W/SIzQtI6H3PCfvjDr/9pXpRs1a4c7L1iy
PJQ9+tkrQc91ENE6wL9ZdeCG77jSo1DwaD3Xsc7TJZl17POO61Zm8HYh2QZUFvDM
t3iQmPq7Bd+SURiTs9UNUaLAjthwwOkkRK6h1pu8YlwcESpF4JzbGByxygfhP0j/
tS/Go01B4ImFSCTiDJzZuB+fxI8P3e/pogb5fNnaBR0iTnNdFFnhMSJl3PZ6t8jt
ElBKEAjoZFLPXJRdXDa/wLFFE2UoKByE9JQQxtU3brRps5WRRPmNNy2fdAOBjFqF
3VFSrQEb9d9R+YRutIq5BIp/lDZoKblmROAQtAyDMyHs7N+qyHEGTmqljHsvtNOx
fitoJKKOujDWc+1ElVRw+vsxxzB0bXWlyGWU+gFm+l8yCe8DeMAQEuyk3VlpZGUb
YyeQx76K25c4NX1fnfA54uguHsee9EhpGux7M0147Fg2xo4wZnQwGbGt3OlhLLZ2
cs0ezIamKyLIiV8rE4EaU96Un3fBRnOIH66SvIN2eDX1Jeh2b0QIX7WDau64RJHP
+iOIIqlGjTgbkOwfBfOt0MKtNj7rM78DAvl2tN2Y8LFhC5l0SQTcseORMIsV6v5Y
Oegs9+mFcbpwGoJEIoqrioEfiXiIxJknX2e4q0Vu7b1a7VLLr8auKxHmsu6EQeum
E/o509K9Wy7w6d1zSFFjo8FB+H751c1ZCRgbHS/OEKpu7Sv65LsPKZEoZU2NbsAd
1GfjCXscVZ0wtXoz66cAEoiA9T5vyN+GsOv25GZT59eDRVG6lJQ0I7gfgdyW0GKB
ITysehnTq5FLu13+i+gECaeoYyoVhyhqlOntHbesktj22tYMK6lXvG6+zXAW0Iaw
pEi65eSSdE8a4T2RsEYIb0HDB57SwMI5ryOvxoQ597DBvdrb08BYisN5pTQETqmY
PnXUq/FoyJjq+s4lDGijbxX+RFi9vS1EwUUFcEPqCkSSfqoIHqOIa1P5MVV+ghva
Tp+GhBeo/9UDboOimaj9FGiy3jtrzvpIHwk0OuUWa5w=
`protect END_PROTECTED
