`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiUbC/n3dDIanJ2VHspGs+GLNGirAuEjHZM4gM2+IGLiTVBwOqZqKSv3eUgHnXZP
6EZBPgIbYyZwyaIuEyHrPFlLRMUdP9hCG0MRzEIMOHLo5Dljw65tQ24c2znAVkIr
b+qlz7f8iilKXEn0Q2Lwn9QreQnmmr+HZGXw7UF1HzDp6xaQ/pbLQy+JB8ZCq8ex
RSzD3X0gnU726ahAHHlxEsecyQXdtdqapFTf/tZpkFYGGKj4L2pQOlmXWsK4mNWk
BEFykLPMwNk1cnAMZTxgUWZsKooVTPHDEDVGo4kTuGuLo9eBXfRsV6+ZeoKvLc9/
6ZdmZD2LMOPHuoaykbTFaUIpqsQARiBvHj2hWfj8AC/+3ONZmlO1k6TW6FJQ61Tn
YOmDyM6Ls0RHxJ/E2/kYApCbgHmgSJrZ6cbKkelPCBt5jQMvvljSLfk7Qk+GoHKp
pAnEfoBWJhKad6wK7VlOJ2QWP1/NK9CBTErfbO4aMQl3k/ft7GOOiUMBzyIaUqUs
FRZp7+oxMzzX5gcE/YoaIMrT02YmOhqO7QJBuo97/JTqCgxigRtXCWvA+KOqfUfd
/OkIe2GRcIGPrmSuzfS4yzp4YeTYZ30PjI8RXxEWfwBCLxxFSdFacyA/lhlFIctw
KggyQHMLjyi7L3stwKwXe+EaqapKDZYVye3MCKoUZLnHkus3IyqPxtInsIk7oOWj
DnRPTUZs67yJt2dIxzymcpsqosGENLDo0fa4aZ8A68tt+9XqMdF6pAVgp8TO8ZTl
j3SKZ2jCjGLBTuu832TirwHEfhBXBvBSNpW0Coe0Iczuz9kl+sGOnyukssFGfry0
IgJeFxA57FmiewqYcvt0+p1TVQZXRUD7JLp41xYPl7Y66/fj6Xe/uHZMTs2otebd
3NLSf+xajDS+6gRSdwSsCWwaczb3DXNwe7kD47x8fmmbQVrzRWiiCELpyYDUHBY0
UQOegGtJGxCAC8j5PFWfveNmKz/Uf2WaoX8hTIR/jOzL5voGkX5BHNu2JcKYbnnr
4lfJWTGCKZAeNv1YNPzSIxGMOpYTRffFpBJjCd5hlBj0j+N6SkVZFbKsBJQ7UN+B
Wnoiz3aicb8TrKJFE8GWCCmyTSHefDs5uSgonWREmFD5GxDZajoiHCBzeCkHptL0
4CfQZOaboEcpU3jP6WV6o8fpJVnu3sqH2xsG0Z5oOu6HqIdNgLNgHi1qfLfvSVVJ
ZtZfR9d9qYBsL5fCwToG5+5Q2H3Vdqn2AmBCdmRsPJb6lL8wi3gKnyLH8Y4EViiv
P+SAHjFtLFeLOelubmHFUUTfIQNvnJf1rItNwYUew2Ki+EO5zr320dWEH1Qhvb/2
BawbRKV51ksYwjikGap92lZhPlb9TxrT/7rbvR/T2Dl6uWwoEKcvdXi4SJVEen7X
fJ6Mrq1Nr6aaHKfPCJEnSzbi929UHCyRMgTOGsxsUtDf6NHUX3D5QzRImqzDcnfr
rpuZaDEES+u+KkuVINk0GTUzL3OD7rtrs2yEhXmIeW6D9JCK1Q0EwrP+LnfWraAm
Et8K/xvCa6A1Vjuvukwshf2glDlhmf3tsFPay0hYf262jTqSVvS/C88Jwv9yfdmI
3r9WgQ1glpOm567z7I6WUd470DzVBiLVGutK+3pWiuK5A/YvTcmv1gB+N9aDhw8M
tDJhxHaFB7OymsuDNvka28507r6OTSbkk5aPFVl0eawyGIa/JHw8jjfly9gl2pzO
LrXwXloq9E2txMgXDH8hqG6n+yR0xzC8OJLynik4cwdHhTP+6IgTDTpbkfLOXUUu
4NHKpx/lPbNIl4lomWj6Qfz8P5HssmOq0R7/JY/JkDeBauLaKfSTkRIuxIzcQ9V4
iQY2kZR/lOTLat8oE3djcru0JrKbuqSfzt38gLNUKC/TG8L61Almy4wfyjP4Yo/S
1nNwc50vof1imc48O64+bLAEZJTvi5j3jkhYkoMCPMuWRCIdY3nWzrQ83XWV1nB9
e8Jipw6BVslM1OF5OiA2PW0CliLL0uObFJwUby8KwLs0/1OyGkHjcjOYB1SKA3oW
r8xP2OXt7BPKXpKNdaL6UOu2bigE/u9VkESvbWDAyRU4w+VYrxyujDJecpLckTEr
lWKbAwTsQZYFhmph5pstbUqji+wjh+pKPz89sLOuWz4C2SFnIqBXvlXBUPfYn9ja
Pb/zqQUtosE5H12NlGU4w2jkJWy6D36zmdN8Zty2+BJasXGsb7qyGxUMp5M0R8fr
jaZyYBwDAjLmDd5sfjEtLzZnP/0VeN17N1nMiyWPJmp30c42Erwj+GrQUNrhhDdx
vfHqv/VC/y+Mcu/SpfiGYTlN9RotKMSPsl0LDAckiQGgkzMccF4719m5IQj+V+LH
v0PCLa71El5pITE7HhpHlR+4nlkqbx1LQvzj53annbtJOIFDNtYk24v7aQ0byfAj
bVX3kMzELoB8BoORTE4QtiFJWmUkeQ4JE0fneyEOM6wJRF7MaTvlKeWbFpakFkKJ
9WuK8eDMO0kxYLHlN4tozMDyCzmz9IUNiqJXDcdWcV3PvB7MzCKZDfgwQOkN1qUK
19vYMswL6ur7+ZWC8rdbpLTVmgUuNuAKDtD6T+PpVVDH7x5XaM2NsVabfmpFJtah
sG7VIx655iHSKazDohMKTPvdRujI810CnggneGwP+Z1wcYriiR9gFC/SHW5s48JR
pY9butxr70yzXHgEI31qlGmlmDS5hOJNTKwY7CB80SYt6Fse2sJvW6YtydEJyAIw
RV3BhSNBg9yT5CQ7CcDNdLlOjcR8B/5jDDyHmuW1emzgdFlLFzJiCsqqzcti4LrO
KllMc4NL2AdxsE4HUdjRqt28V0fhHypDKTBiH5xxehuKl6OHA7OTWA6ZrDYfWT8f
6Qr13j0SCsURlET0DIQVEOLsaBc05JaPjIyH5qlJvV4JCuNUG9GUIvgZnnR/I4qv
QxEtz5mxDVFax4rtRxylo8kbcwmmIGftoI2eV+TclShBoexwpgZIkOCF8SqjQirS
qSgdyLto0Y2UXurf+bHUTtStFuYlKGjxQuYnk2Xioa7JPZzH12jYdbw7IzbrW20X
UBfv+/+r7zgzAr5rxgQcyedwnBc62++BKgQ99Hr20vIcIrDTMvor9PquiG84CyjD
DCh6SpzbKJ49LYkyQ58kIMxiQg4KYKHyTSjKKwc2uBdtIh+Ug/OIozmBCpXO2ZSD
ictkMbKq6A8HbfM1XEi5xid4C/cmpjMCq2jnmQXW9r8MENAKEDmmmKXVTvL7BYNL
78h9GMxnc6v5X+L5B2j8mKKSCYKI7nnMdLYNupxxkXXDmfYnTSAHlONqnc2WL7va
9cP5T3QopGXtYEkcwZvT9A==
`protect END_PROTECTED
