`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xC6Ry0AWW6l2+7FjW1r87ihxZlczCkjavN3R74SnTVWQoIBjXo3FKbtp2iZ/7PPH
c7bHbRIafl/YsTHpLpcgC8Mzwli9QWP9xDNHcR1cGjM/TBMmvNwuexajhH03y1zs
LWvyoRh0V0MTlurginqfJs7RBDwL37VWBrARhs0qGB5SaevMU50OQlQckklbvXgM
dA6K2419VZYOTL8RgybkDV3ZIy9yiBIhtx5IwpLfRnvvpJ725kyKEGWqD0aHta/K
h29ax2uoMK93uJaThSXq+Ndgj1Tcpkp92e+cPzg46+v3CMzsMDM6F59sWk8FyWna
go1ni3X+QOWQE3b4ZwQgDp8OPv0/qhqfAWEhaG81NYG8B07QqF2HNtPuP/dlDP1S
EPkc23KWF5agnJ3X6fDhFlaX2CyDh/YW0h8INEOcw3yElgFVEkVsiey6AJAUZOJj
`protect END_PROTECTED
