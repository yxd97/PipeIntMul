`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QeJNkQykzjPspY+KGq4QpTMls4yaZTU5VRUmjKu3avOWCPazTU4LxFtJjR0ZT3u/
acGqOxNSzqDxGU0vaRcp2qc7Sj7ECZ5WBERayFJ8k0jeR7h2mUvydAlGCqFlw6cU
BGOdfgQJZPj+z4TJdqKaf6yeP8XB5OfSeje+HZlGL7Wt2Uof64oBVseKrnPTHRyP
xjaX3NRtcR0TsXqlYQ54rsKrBkJoy7uneTaXLZJ/+iUQgUpaCRyeM7nbqvcKoZ6s
yCcJoOq6+H0U9hsCYHey9Nvp/ShrMEmmnYsiy3m8HNvkXDxhILfgmXUIaxak53nC
0v/JHeVDJnwyEs4ZHBDklVN7OMmRZdTNPg3pl0NDCCjVaVBUMhHTalIZZijUy1VJ
0qq+jB1vv3rEEJLruAzVmAFqZPpaR1YMoCuQy3fPbzBrmdYNttufznEUVk4bRKSb
6ABz8k399RCOcOz9yuTCuDaXms+OYL4E43M9QI3i2jQU1Tyjx5YXb0Cg7XABn4vE
YVTIQxFJ2vBb7W983TVAVGApCk7YNXBBDA5fS8g8k07qTKBt9xgQAcUfx7hRoTgk
BGO47ZG6WAvHo44zOEdL2dvmoR/V3fgx9MwALJ5JvdCY2MFO7CmPo7rOTOpaJDiW
/bXYE8Wy1iCPxOJ7PshFlUW2i9unLKJXlvzapNWaZV46xcUsY4SyNQPHtahFK48Z
i5Xdl5J394MlHbe3RPBODCKcngbIi9gToFTWvEV5hEb4RmvVL4hBKMdtrGF7mL08
YEQssQR8xW5mPiysUcqpWVnS+4FPQQ8N2tT6IvEtK4MnBstN4fM7bQreVCg59DYZ
m/S5CduDfcyK8xmE0TxkYKjcGADsx0q1IsM+vcX8TOuxiJ77rOqBpNTR1ZS+Diw4
3lgnHDfLuo1gD8In3Vy5sElyznZc4M899pjEBTSVi7udsSwkKcdx9TlXo1qaUKFz
BM/5FhU+b6HL93OgIA7C6WYm5qhPi8VuYtlbXYLfuiAoQmIEwN0L6O+mBzQO6n03
uEWw4Pn8o8CaxVOozVdCQDRoV1VcPZLP/7vwhviebx4d8ljIDiM1kqxedsxXdxcO
ziq9YMzsGGWR1FjL3pONp0u1a3p0BOHBC+imZ3JZPtZZA2lccCwzBOZao3awFIpO
dKCNJYfaO8hL4QphjgR8dABA8KTKEROPEvJh6p0lbg9d+jSM3BgUTbAQYHfT5S8m
BiJpSViXJXQm96J1NEpeYMQE+CHOl20nzgeaoQo796cUdTjl/RrBbAvfwDvi7UAJ
JKgLAeq+0DHEU1mjfAjfxRMvtdjr3jbK0S/5GNSQXMmSKGM3CHeSAJpToHRaKDtf
6aPJIPYXZomx6Xwu8B0xd0V02ZJJvR8NgYy7Fx7YlW/BN7z/GCB5N1C+n1YDLWei
qJP7PjtSR4nf66n85ex3rrsoWI/aHcBbpNWC6reFmtFFPuSUv0d2SV7nsuVpEkVT
iv3q6UXWjZ+LKSQMIHE8DDRba+mlFnS8cqkYAl2vEvbk2qS4qXA3WVSVsbPMtTHu
51q4OdyeO20N4/FVFSnwN850d+x8s/fqE1nXGlDjGTNeFxR+q7efsdTp9Aw8aqwJ
/In8sOs6LEamGZKgJ+d0tF7ZCWxTOpv0j01d1cZhceRxUPgz32FzZOtyucopRGt4
KSdWTBQD/pASiQMr76Lx/E08sCVOLXT9LFfVtVyci7MiO8XZLh9LKnTQPe3xe33o
2jXhZsRCD3N+/IanbjMPj8SBUk1sLKBGj96OoqxlUtH2rOywOvKlVF8htgodIbtT
6Sq1vHMJa4vUhqhhlPUa0n6AYqB4eHGTPkBogzZU19aa91VGFah6EIOUpkm5Y4PV
31UxqOpQktIw3SsGc3sI8Shs14SMf77M5Wnr4Kq4ljML2DP9/C7puf303MP3bCBy
NAuQee5mCjHgwEMJvsPcAYjlrepbRVPv2DmZf81BcIjVDJJP317k5P9dpZbFHG/M
fzIHGPfJv3O229F+7gChfOzL9vAPHFPC7sdIYG8pdSw+IxcWC6Mns3NwGUWpgjJR
kr4eC6Y2k/9F3AFNlc7MfdI0GPP3jGnQEmmpW16uYMkMjHgEdfUW2wLSiQ+Jcs7z
CssHMHPXteEXqF5xxjkIHrl/xherDo/9Q1RrHcaZc1b4Qf0wTZ2hb2oA7hyTevTd
`protect END_PROTECTED
