`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/EPhEF2OSy3IAevFScmbUrFqrOS9FwYBKz8X2rNCQEOHRorfJkQtuL0J8c8oST3Z
5RcdRVZpbD130wQmd7chsJ6YYHG7JFC6FpJD7y/IAHTEsahomOf6uMa6ADIa1mRS
yL3mjJE2nPVPTU2R9TcmYTR22kyRpMmmPJjqRQyx7oG5gqxRRjDNYfXbxRVkdAi/
XYHP5858gMp5JOQifT1ybpu326rxoPcDjz2lP7jvVwW+L7D9EazeiAANT3iSFKvD
qgZ1lSR9R4i5YX+o2cKa9kqpQC5l4Tn5LC5JFmALrzLAc2PRFHIlpLo+JkkQwXdo
sM+OvEhaJX/bzc/cDQaE1gNs5V+b6dBcThXaikfF/AsWEW+lvwXmwqDb2/P442yy
791ukLzRTCzV3i9Kbg7kMlIdxIP8P+9pnCzhHWYNavA=
`protect END_PROTECTED
