`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lupATwg07rQ/sXQH29tSmgehF6ZKDs7CKCq+h84jABLgzTcVq//AJpfX/05UQIki
/lXRuaSljLktVRN1KvwHeF7JLDt+/Il9qgaPZbMKpjhc2soW2y9qkzxax/N7j9p6
zzOt2kRTNdErQy8n7YMLGs5v3cjixI3FKF791fMwRqogkuX8EjeAt4H81aE3GnH9
ZxpqDTaYUkvRPMT7Rd0STUKvYQtNdsjOv4xiWDldhUEIMFgLYZ2lzjx8KaKcXMrJ
FEswAe2x0JAX0qOaxFLGTnhp1/DepkwtJ6YeXEyXtpOAS1Ig4jshlJfWu8V7zJLv
iupj/tL2eTDSp9Lp5XxKLkj6iS34Ciy97/L6aE9BuRnfMcjJpi0TTPCl7OFQ8hiC
RMn9UGHRbfXV+GvOOOgZwA/ic8ZxXKsmegruXjxJUlzOZW5kMIJwdKZ5UUe3zqgK
KACEJATuKU5L/fkouPLfhYLadfNh5ANtT7UPkzFGi1etWtDt0o14d9Ljukoy7xkU
5OzJpKJEnd9PYwCjmy/5pzyEZjpQQvYL4rswu+H2uOX9CgDQvxw9+jtYDxIOk4YT
mM4u8hdgKOdMBje4oD/kZCBv77/gACPqdbrxRR54+CrhxC0+cdMD1xJ/Hu5gkShY
WoFdfJBdeBYLriKOdXY3py2L0SuNCvloRgvRhrUOvZDtyA07Z0hhGHkCUs8odm/Y
Gs9OEVSChi95pElaO9V+ijKqAg85FxLgySCjvcoE4SDGdk9JdsKuqRVz4gDIub7f
HZQyjh7TihDg4yokN1iZKKlv/X65PsZSBkbuekoR4qEaEFhuW5VU0Gz/ngqswx99
/G8nDFlQcjYVqgjLvc6UVvClwrIqYzl1Yakwf5SF+c/cbxrgJW6MmB/v6eDzl3Dz
WvJerTzAp/Z88XY7Z2nZ4zDs4rhRa8SZPvXbC7QCNgI64Ba2ZHo7/eVf/SGyyt/a
DSz4MzBgZ02D+J1wRrs5kKYdcnH6s9rdxuzJNj2BDaGEOvhpkv04uIetqKL0Ish/
MxRdCAaDwv4uLIMhqwyuirEo+Xk4Ak1g8FX3vIGH+qACCewXCFXFzpdbfSttG/mU
/NPIap3g/xH2EGNr45fRRe0JcCMhZVMOVNsQ9EBCEL0SE2vPC4UwXiexxrnVkQRj
pYp3/6CXel5I2CIE053xnl4KgkR1NHzsJotiLXZNhek/brqWEzm34FZNSS8gKbef
bUdcogoIr2DdP0LrivbYr4KDcjvBYHSSBzmyfw8UXKAtFYxBfxhbRIxM9gl8b2sc
wGmJHOZ5cWmj/rXfLQb/i4p8xoKDAjXcN2sF2EewIvSwdB8gVQHWlISIauaB84KZ
97ijad+QsMHWvc03wwxe0mRGC902nI2zFH05mFMSLqI2avokJUvvlfWNfioUpaO4
eFU7f168tK+fTxeaOrV/ZSmVSBxDhmh5r4EliAgXw90x805ZxiIQQpMMfm3PjxpM
Slfvlde0rEk6DXH0K2KA1rqiT/VYgo31gVxQLDV+8pwD+LXsHRDbf4CAP9NiuMBD
Zco/zE3Hz8OpUvHTOu9OKpRLo5aKsh4cAlOl03S9iJIW2SEQfulGnTPodLjyF7gV
UyPYRSzOu0/OAKVHQtIRFs4v1nZxTbakj9yMZveqfhlOVa8RM6X7tdEwW3zSrA32
nyB9Y/LQAASk2TBjce5+eJr2amFwFZ4uYFQiKpYpmYn//wB4veVKvOvZG18TTKyf
/K+WsjXK6/aBGMKiyGuvSAeV7aWanxtz1wQC2X4bXirS1VJTNOktfhiWhV8Yb6PR
MPA1d4XM2o+h9+wNz0jo6jZ0O6tepbuLU/H5EWf18JXSWlBj5qFRRvIxMy8ybAkX
ekptfQFHXKF63HhIQM8TOSZc4HNf8IksgEX7fJPoymEtwEosMk/7I0Dx218r3RdU
QnMzskxz+pp9h4r2nN0m46u7PfCw8d9V4rn5S+bf3L4MIn0JVIppyJmUWfBMyu3G
MMcL10/M11RrFsRphbYvSu07/QtCRn/uA7S1MkPcl8P6oaGEvqAyok6CmXvFyFaM
cZD6fBFqPZLHDz1UG8C7x5SyCY2VUuxJ7ucdsBPqKdZExk7aPaHVd9LCGl7SAy/s
Cfje7lvc93BUZhkdgOsus7KKBRjgUCeatm9uMydJzyU3BxcG83BIzl92Y3eAlxb8
xscIpPz1+QlIJK/dNgdwjmbvDFvYavyldR5wMXD36JzJcbgrVhsj+9zZuxXdKb2C
DwljLzgpIGS1D0MSZdifycNOynL4vgOxsnvfDmxuI4M0b7XdlxLrQtVEEwtuoy5I
3lXgHaLRZsRN5tAGg8e/mAsrK+ZoWSt8VgE5LJC7qr0BewvgjRDSRPtuGXACFCzI
KjQr/2205hF1G+ZJFk10F4KgbDUPWOPB87ZAwWaJWJpZVZ24R/mGxUkX1lwvnYNv
ly2qaDRnqT+k5Ylz92cQtKHbx+5dPfo+BZ1p2DYmplDxARNEQ2tS+eIIJ6y0FGQM
WHCJ88moSKFq6jN/IziPFu6Wwji8U+8StkAUDGPZLMcFlDQc8suxcr05YTpqwIit
relBQrD2ydQfaobp6zVyZZT8j2KfbV+GQ5fkVYqlTPxo42m815BrTLdnfKddBgHA
fSkZemfceG7l2cILFVa5CkaO+FB4DvXERLj63lb47JMQmxESznfJKWHcjgZkbp8p
HP4r7l6dpOMQvHrOY83KEfYHLnB6ao8pJoJKg2N76tZoKyh+VUL7IGG2EUn++eX9
tXP9a5F/nsXAe5nK95GzPO5Z642hGqyzwBmT0vBUtwSCGLet3WtZsq6oE+iynsKI
02TFy5b6IKm79CISBNaPjrd5gHkEK7KaKqQx+qSCsyHMbat2Lde4oVW8fp2rHJAN
CGnIrI9itfsT7WKTGl4LEn54JfGj94o3LpK1FPm1EOaGHCAXWxVLeTr56V3D7euG
FAGXwdy4G6V8mIi0EvJAXl7kUEhtlB8Nfw/nBZ2YTelfsRfXYJGHuurTsj+Er3vb
gTHk35O9dtwdsPOAJsDv95TzEn/0DbwpnBFH+tVYs3adoBCKEOwr2m+nTVADcEzO
u6rnATcS2HHd7dXzu6MEgoliB6EdjD1egLYjP5vXVXpFExyvApa7+W5qjzSNn0TC
0Pu/hQQQ7aQjUtMrm3EJxIVv9dETS9WalSGqNGksqPw9kN2oIKs/uKA4CO+yygFC
YZ7+Uy4jaP6w/5TkavAlEtDTvVTRSwDE9RvA5VC7vLosTUxKcJu59U9LzZfV18MW
EELrw6AouUWKyEVsHMXhzkQ0b4yf4TxestHqVNWIVSnhR+I1MrSibjaQQFq5pgBo
nkuB+Rmt4MHR5TXOiWbzzfAtDctQ1x3rn2YrhdeVmGMimRA0T14XYM1BnoRfEtGe
n5Om+4HZi63Hs28Km2d++1DS7NYQMmxsHgDS2K2fIfu/4dXLCgYVnSSMvYVnBpET
xgvqTx9QDQG1MKhoyT29fj3iGJu1rZQ92XM1p2aiExoP9RR8R9SZQIYaenItTXLm
Tldl7nHlQxIbR5rAh47zSQdgjAAmzU7Qrlte9LYQML8jm2A9cKwoLmFKSPw3QwSE
P5KHvYLB4Nd/wGY9is69LGyd/AKZ/rEbH5MzmajN++IMBM3vhmfZzsLNA3EaiQbM
GVjG/38rkwi7nnxh2IqDWSVTfZ0SJzQ7ncty3XHyn1EjjNuo0tk58Bye9xEDsq1N
jCI0OpxzUq9qdaQKSay6IEFC07CKfQGNIcegn8nm/HKhH7KAfzAw+AmbOao2QfOq
50+OQAode6kcf0f+MwwVuvgYQYYhVGc0shLRyTUj5282tp0EoDc25bkRYjzVP9Zc
dVrUgBRJSHtkclFeX8qwKC4f1sQlovJaUsU6j6lAx+aPoOyIIPauXun+HhUHxl9a
qFWXEZLVXg2MenWz6Ky5BG2LH9oL6yEceoel/oCmQNduwPDUK2lNJ/blTVjd7aoi
ADFUfcq2QU+YuDgGYD7zzLtSCqMQDC2Z0e4S/7zMZSFg2k/u+XFN4+G6Q8LYrm7s
W/0iWiBJBEHvGc+gIxMryZcrB/3vVLNCFTQnx7so88hrrb35hT2VJmx9dHXrHgu2
UO9dkU/rTCP3qf8VSRxkyDeiTLYFgBeN8ZDrjmT7uAqC0lpNZ+oBdD+Ndsb1UEqR
O9SHpjyVJnxG9n/dTrdo+hXkFLdguQYQMHzbxYdAAZHvt9dxUI0Zj56TiWqPAZTV
8F3LqMAsc3KarQUZQH9fGMjjAVo4CprQ0gTjoUo6v4x2U7rJEHHRdCJ/tTAqRCVv
x6k21qKLpVjlqotabixCqZVdPEqFOVodgcwdtdxdBn/RKS5/lZAZSZgp48AfaTZc
IqJPL8Sj4dVMmDDeeJ/RoealYT5GsHuYjIpv+GdQ9YU=
`protect END_PROTECTED
