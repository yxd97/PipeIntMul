`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQgpocDtls0gHUNPrskO+T63RYBJCTuSf7dwgdf+2xOLyY/gMTs6F2LuMDTZSN6l
QgAcPANHRvlqGXGFBiP5jVjcm09CHdGF54EMMu8HgXIDt1QBkK2xVvxzEFlEGAav
8kHhJJKyCMuscpHZI33vUP3Pjr7JRLOwCzLWB3z2wz+R736ReFd1NHZzQiS2PS0n
dbp00lmL9x1+19h3wq4wAJFkq2H1+fWkP7VM8KfnSiS8YnYXBAyG2Rt1xf4X+A+2
TIcRrUABwHXfoDx0FeCqDJSfLNVXbslIcq47L/QXMwTz8wzDOSqxDLIYsCu6fN0L
5XN4sYarLyiu8zPNA29WyCQAV6lEZNWlgJJnA5ooXoZZE6p7A5K23LkIMBX3ihLL
lpPIxBSdT2rlB9PGuoTttHyWHxFYBZiFiwojaQmDWGpDriCKDQ8Akxi74/3o8afz
OIDhutq65KNqDMU0hCSMFIYkpTK1AHtOTf3zOlB0jRvjkPCPtZmSTb/A6wg72FPX
o0Jr+itcw2GTlL5ON/EnyapZzdavr0suCIudpD2Zh/ZbpwO0+xymEtc9LZZdTzow
/g5z1Rj5ndZ0HlzNIdz8G89embwO4UoHm8NP3cKQrxNVkGdc8l3KTzEtYjtm2t4i
CQUy4SGfRom4tKPZJVRnQjtmycVOMeDTIckfgqeZ4Qvm1jCZTu53UBz5nrXRomHv
0W4ReArcwLLqx7DJpNIPrAaNaqCrZyHmEdTxqFIbF7RSDkGG4eiJTM7oz3apC/6D
bU7lcE6hya/6HNVQM0erOlshfrZi9Gt7FgYAS0YS3QRzepQ/AhXFp1NIrWQeGeXu
pzeSe6rAGAu9elnxMsUDDd83QF8rvpQ9+sVYDLRCVuHWy2jtRBU5O/bnyHk1Kpup
Y7E5qARgpJjNtT+zoNHb6M1le8bH9dkZrGTj5tplM6f3RBYMBpyoY+QgdAyVkUU4
woQvdb9wz+TudiQZECVTReWdTxDZDekQnjUTRfIyyd+tzY/sPwpDgy2SupSfXkcR
THR8xoAP+SGTKIjVwJY55q21zuPWgcm0VP3e9WtJLiEgXf5DUC3bPK8gMUoVZ5UK
b2gOzYASpbkGXopFfI1OtK7790KWFuKO7tCYIRdC0mxilQT6Fp/eP1QMZI2viejQ
e+afS9dXjBUXFVicNh/pVVOeYsu4khWg9U1fFVOOZgQJG903ry4qiZVZ1X54Q9P2
x3Ry0MNIZAoPDqV72nnNgSVkMZzbKWqVtQPkP8cP9n/uQvFrXTRBHjG/ej+wd8NR
pfqZ/UVDSaBPM0SgjAUQAb6xH3XVb3RgvvJJ0pq0EDomwIJMqHjlLE0Cjkf1dHfs
WMNeKpJPtjQuua/UcTpXGg5HkaH4RnrW1asac126focUGXucTMW+DTFHOdPWjwiy
U5X+90edlKrOxEiywdIiOhtIA1XCeourvRGnSg6cu9/fbfG5n15Qcm1Lw0Zbn+SS
ZOPDALKsjobiONDwM+SfnDKH77ETzWraYfayp0UG1NSxq/wBqWf4BcTaS0D1SbEC
3P/XAv8Bqmfr4rDT+zQh4qPdn7ZVdJZW1RecUcSqMLms1TAILUhUE5VddQroP0Ry
8AA+ikJhIUCAsPVkI74THvEsoH6dsoEm4gpggfG5K0YarbC1+jL9rBLiSmv47gUN
8xutU3NaB1YPFBIeSygWCw2h/FCgn0IBfKgskD/FqC280x42QWYfVZUA1H/iVuSi
vCEj+WeyEQmPhQBBln8ZIaNm1q/8aXqf3iyH1ZnzO7Z1BlrI5EiSU6PQB7PPqYU3
rShp1cCHiMmRbv3SW2e11FAHgLJtg3TpbbDfmN9DnmH4lZ27nf5rdzs6b9gLAStl
LzooWOZI5afRrIWD8nLD752XeOZAZp7tMGRdmfvrdPM=
`protect END_PROTECTED
