`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UXF3Nt6VoRF4qrdnXqRjhr1waAhmezdQz8HAIBahqu9PAMFdQ4FzvTri7qk41LKO
y4pMq1NIIFOJEAMhNtKThfr6RtQL9zf6cmhIPDVzA7TGt9sZ+zUtqf/81KygE7XP
CI9rjQM337cOdlkCN822iNK/NMmt+Ua5Yub97mDluvic+/18I1bFLUImH0B5qsXg
cKPYa+3X/b7FoBtdMEtzsabPY6S51YQx4Z4wil+zuZX7cblo7YYW2bJ43FjkMX6K
M4pXm8O8kQw5HxtWh5Bx2+qTnu+OAHd2BEfLgwE6mH4sbEQNhtExXRWuz5nJtle/
8WCoac5aP2eIR4dQerZ/djTLZG+RQtZMuXimtj0HoKCpc967PBcY6XjMqeWUiKkb
PHr5nGd5eQ+pZ2U+YAhXhHfJJP6xT8mM709V63u/sIw=
`protect END_PROTECTED
