`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IyNxcZDngYGGGg1ZqdXZ3Mj4bkY66A0wkOLwQTxeXMeEl4oxjo6+VMRJMGBUj6au
quTQGIk/rHZgkDDcEqSxT5r2fWqigd/8F932oNTBxRLHWr9sWkWI6eFuqS1HbEnz
OwhpRMefj/+3TxaBb7muYXxr+BW9utonfQnrmHfVIVLvS2fEiqPR7YpbcU+Ibg+Z
9T2aG4BeCOJvwd3MJ4ZSc5lu5rF0HVFXQ/EqgtoKdirv2YNDe8lczKq1gAjE7k4V
q3kpbCt8wgMI4YhMIHTz2Pc7Lp5JH7+Cj0q6tuxnEKfNTGpItkpeDIU7+lWB3cCX
nl6rfLXknDxqCFx4w8FvrQFEv6Q9F3qGcerukevEU9BAF/lSpfku9uzarF2aSQ8J
x0UPucqoAiMWDrLugHn/PK1Bk7O318lqlTRVg/G31mGTs9Gc7aZO/YokQVQiHGtt
mhI/QEhVCD7ajsG3ziKqdFa9+J+UtuCmDcvESxQS9pfvjEB3VowiCoesx/mnlLgX
sU7AjbkzpCGvB64ELZBhMLz/l/bXQ2WC1zlo6LzB1ytjIQ671HM7psohUdEbhQ1n
hM2dJG1ENh0qsmwN1dw9lW0lyWWmDlM/+J/OrU4h+GjwDG/ytJTILbgwL2LxUL4j
T8ay0/SCoFAmV6ln8GlaCQ==
`protect END_PROTECTED
