`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B5KD7AsMNMw7r/OdKV2N7vtzWAjnRcSlHoC4EN027Qx+QXcuCH6/4FchDHZet/dG
BVR1ITNOOzrGTlk21BL3quk06WhOMc2IXjQiiJxAg+MpVQIVFvDKp5KxxUplaPei
zzcBcfSONF9ben/yXOsdty+zxAK+zPd2grsEZ1kyD0vtsYuun4vTJOupMpSumrED
3vY6qvilN3Q01Q6Zinnn+zKWMDOf9XgED2vkstGuUHCXTySpKLr+1eCjYFCtWef+
FEQwMmI882R9NkfLCvTVeXinp/+WByNtZw0As3q1jf7oqJURgFmssZvFzHT7caI3
ZHC43Hh4PHWRccN0TeGIrRBG+AzF5zFp1LNPwUdQLSdm2MR6YhKmIv/kCS8BRo98
XGwEmPdxBWp1ik5QYcvTTd0bWwGFpXl5Obl53M0mr40ch+WXiDSgPJcl4TShoBce
CP9Fc9v99D4LwkNSZx5BOZuxa+PJ9hQJ8Fphm5qi+9I4RoEC1sralSRbC87H/eOG
HDm+vCnmGpuzTf5gEOMn40xft0O/sW+KgZGpzqAD/+37+i/0aFp11+7xmTKEmCfd
0+PcuzrwanWuQzmadBswPX8PflCVMuMVm+yFJsZRGm6O07QuF7G+c2d+yzR66/vI
23xhvgybfp9fq/SiMQzEHsZLkwJI7dSQ9s+1vNZ7xxAZP2WjiAH/t75QRIzX4vXt
bS5jhFvicRG+xzXS4dV3hdrJ+ClHmR5ALm8DsAdy8y1faj1xhRkhp0DJazbSk/Ni
MrOJ+1LiBT11N9U2HttrRoXvVNnNxDbJGRmFPT19m9oZJ5t02KQDbFPPOOPmtCBA
FXPQyfqx1fGfLBskRQihHleJlgeRV71apaLwdsYahfyaMNU6dHUZUV6qYBrcTHRL
/erx2vXqXTLnPmkgmLQV+cuOTpSxXBStVdS2frFbLIS8x6V4ZRBt6W9mVKXYo/Dx
z1qClVhN5hh8rJWEaFyx7keMAKxFNI5x5t8CtpvZ6pwEIgF/caDd6ZS8ajFmpPii
yc7qQOWv8/dNJR8wNjK7fjbCrsvGXtrRfT/35hMIp1cvnMwBtxHvBjzpzD99xG5E
l8yrBZeR87Jf3i3Z4H6iUeQRx62+xZjKqCZ8SJ9s8JhPJOoCQm7pgpGUOsOeJMs0
m2EfRlvjiUwFaA+fnQSLApNei1YGUZ42YG7tIe0SOp53/CBWPNt/Ak3e/lNCSMfe
sg1J4NzXhfzPwDg5ucBvVL1mLoVxe3W0+/kHKO5fZRSsIWQKfWH662UUoNkH4W2J
aCTSCxlcjHFBo0Af4FA0f8U2OyXRzoRJsPU+a+PggX3QLrYNi8dTAAiYZioM4PQM
UEsO7tDZon/wowF1kh/t1WBkUeTWcV6L1ut6ZK5+sf4pq/xDYHPHDdd11h901DI+
0L0SUmUkckXg4YCrC75DKAAc/X/CnONpkmiGNXe9nq0OG5BklfqvnYU5jZgrISIR
Brrk3aEAvDJsJaSR9GXfA0VxMKx2AQzoEPfdakSe4dwllx/bYSeQQWKhfTV2a7lg
FW3MIFy152H7LJaYJkvDsBg1Vw4S+Q70M1guaozUgiahhYyU7fhAPzCQTLUH4IA/
AuB5PBW34GnnJnKxYXzIr/nU8FuZp+Jypx10PkKV4osvcv6Q+i5CxvVFNyjkyA6C
bMAngoR5Wu1A73lew55eveRKBv6XJULg/mrMq+u5gKnLhxGMGIk1/OMd1RWlVBWZ
9C+gY90uhw7lhtJ3DcQKluR1MIQ+mWQr+hQ4qnNTnmclHZG0mPJHXylLUKI5ExMv
pRWxBPbiKdvSaOKnt/s31keRkhhJLhmqKOW4RitEPsR32Ka4rJ6d1/Il1rt5BQCI
JrvFzJcsvhKFMrLSeeRbN9Xa+rsVeyXAndwaTln31WLm0VcXSIdMZmEXX0ZeAqmI
HmboLMtaw2L+pMGQFl4uQGp1FCCIjpy52GYdVA58UiBCgrKX21mh+iPwT+r4rKJn
m+lSt+C1EI8yjS+NGeKrZOnm7QUSp2ccsY7EDeDWPIvF7+4DAA98bSFF+Oin88s+
JfbdtnVQgeaiSyMNsLT5vMHufUBaN1b4dX7Hau4s/jNeasYLDoYAQ9XzKL3w/eYr
P/e6dp95r+2QghL2CotFnUs21PfimSwYLoWdBL23pFr2t/aINQTru2QuTCiwnYHR
p0PHtu3jRsgAz73qzbw9ikIM7sZBBm+FQyohr1dGf/CzzPtZccRPPuuu2m03rLvt
jrwKSXkHsKxAqI8kZC6Kt37Qs5/95FHFWtlMNEKEIGI89/U2SJCXyeVEYFI6r5T8
aVsOwUC17MkZn9DxJvrlcFZ5/9ianm5CouSaDnAhiToF1ExynEI9UbdObtoCMx3Q
61fRlHmN9J/+r3Bb8xvxuEku1GHBF9BjB6l6VTMej17WvITt5xi6v8TCnScpRwJp
2r98xdRg2gkKvZa8YuX0d4KIJagygB4hApR/auoIIwJa6p8GSS9ph9DYuGeuxuGo
7ckYYAnowIYIKhGGNErwsqa6bZq4oULEQIDrFfOZo625RQPxgCo88IMKg/pewKyd
/gMq5FtXJL+XvtAvEuuH/TGALtfS6bL/Z4Mla1QtQW3/5MkqTwIFhe2imPNutTzx
ApOshlgr9Sm0vr1rgAUYK/lx5hE/dAwMueUnVj5AFYzgfChuPGvNTA2Nk1uXGNV6
47ITDmod+Du//oAyh+Xf8qGIHj8lpT8FWmFQfa/TSPNrwn0eLhWefYi8eqCe8kdD
ydzMcDfp8ZhCE8Fcb9F3uXHvRmZucu0En5KjAxHnZeSf7X7BEha4gTkUk4UD5/wl
58vEAJLy/GSc72Q6wVdF8FX1IBgan232v2+9gKnB5nB18jVwGRAhrSKghZt1n+XM
izM0lw4j4OO2lrQEiBg+xPjhKlJX13HzKR1Ps4FOTZsCNzlyWhjFAY9xTBgVrjQj
ZmI5WRLuxJf5+pTN6oNtFQLSVPxIdYhYnEYbh0Dzt80FHR9w2U2FsFsVA92xgVQH
CJZL/RnU/0TGTsaFslU3GcuYo7oK7AKFP+zOLOyYk4OMlUg2Gzzu2voCGA2TVbEK
zNyXlsjuMxTge/ekLLSGZhq+bWkpQgK8/mUECU5phuavrud+/EDlZDZgngD+kOoc
BiVCNbj8VM2Lb4ZE0oRoO0xKrxa7keATYKCdEIur4ael1PHIXWOivMTDn76YiPa2
pF34vBansrb7O902VnphMxrB+8UCpfiVUyCyYrf4Zldchtv0lQIi8RXrK6w3uyga
e1l12ZTRwGZ9b2I5597tqTCmc4i8RkY3mKTgxV2tLCiod84ndqtpdz1boRkeY1YM
XHpasOpQADWtfPJncwi4HVtuDLpbphvvwBGbIu0Yf1x75ITZRBmWGtoNaoAL6mmF
JxVX8oDtFAsswC4NFVXd4p/Ik5DZLWab2nPW99JuwYKWXYD09ZohLToIpe5lpFj4
QGZFAFLMGiS7mnlQ062Z5QPhrwDtnVcp0D5uj1gApFLhgThvm+jdVbWa91vVl6hd
yDbnFq/XaeRkpLwwV7Txa3gdxh4sCRREMQmqu6WWFB0yZhilL/l7mwkwfv1EpgOd
N/2HxoLPHYYz26+jbKARZ7ajNgnwN4ulf3IvYS1aZQy2o6J8Fev6cKkrJdK8p9fI
VhziIIhTR6NK82dqiQSb4RZWF2Bt86Db+6dJh3AX6qeNbz9LY+iylleEySRbJGdz
mI8vsNWltyQAOV8brH6pMX4VsTLr0Okvh3BSEq4NKuIWP9B80yTfQ6S4zdFE7wPZ
Kr/3lp1amz/sT002b5EToZv7+pLG0NfDx9ZHlm5va0rCaCRtTbmfdYDpF0htgE8F
+AtywGLD/Mi7AhVHGLdqFJBJFnjCLD/3nPh8v9Krgga6xxt89KGsPQ6goBLvMult
21eT5AyyReUiytDOUunC+CqJ6YchNT+Hnk8GG9Lbl2TO2qdoz7xHLQkCPMrkS8SE
BpbSE3xaM6IMH/8OzPLEm2aeaKL6UylS6CI4cyNW7YiOVGwOk6JLnJiyJvtDs0Q4
ceDdhTjiyHfFU0YMO5QvZU7uCKF8Kou+cEIEw0Ya1aTQEC4/OtVb+zs0e1qqkrc4
0LpsqzPf1bD9e+2yPfTbpoFX0ASTjKvP/WZZJDcFNoYgNTgvO0KafP439L4+u7Gy
GPfZfNRg5XT0uQSB/tNTDBIPXWX+l03nqcFnjIOgmiYhd+ZkDdI41ipGlxnz2DAh
/eI2fbhJ5vNdCsxO6J8/lTC39YvO8nNLIDoDrd5p7Z/8VuwARDgfA57nmZ5pS+Hs
+JyXAm1pBIBW2KogPtp9P9dZFxgah4qdnGJ25PlLAK5+HQGCBv2/6Oe1qSOvRmgv
MBXCBOvxjGTSyEcx5KBYY6vwrSlwtBuDXgIafTgBUT+Cm520N2+5Y0jSX34UXV6o
VhPCYN6QTCZ9GxxVAoGrkQkpVUeSVlVsJ5Q14CUMEaonJnfETY/9NBbsAPo1eg5K
PfYjYfcj0gS6lzhvumnJCuKH1EJEYOG+QCrmg60552jI9hWGEV1ILBxl6ZNpOJE9
/wZcEvoRJNXuAo0Y2stA1MdFDBV6S4vzzjfJ1dGz0r5/1f8yOcUYUcU233OTkWK7
Wu+oQDjrOrTyzx2o5efwOe6mfRV+qFNUy0C5lGdZ61eROJ+shgZlAj6s9e2f8fAU
2ye5NpsFh1kgCJlq10mPfPNEvXk59sHMmejm2w0Fo07543NBJ3H+YdiuYq1OCYow
j5lK8fGIZiILY2q/2C6DtM5TFjRyegNB4qaNWOGuu1esVpHtSQjNf9ycCdf8qoFP
rVKsYZnCQ3tacWcrXXI/xySObNid1Ftsjx+M/XJEWFwbStBHcNVD8J2qtchG0sPX
AE9kdYko7nwknJZM/nRadizC1nAc7aWzmwZ3sKLd+07vMW4NxlJHRWzfJ7EUGErY
TWyptsvK8rJci0l8bMnX3aFSODkOj2lcQSAx8BZlm80GnrFMu4LYTMxRw+ijatJT
tRvy6ugbjLn78hVHmuuZrIuE6M8euwpaS3FPhsTNGGgMe4ur812QC0u81CbcqkZP
DnjEbinL9OAk3QMc4h6Jhjy5Yy3mNWQurNKTdNdcKKvT5c1E7tagAHI/Vr2GOSG+
1lqqTsS2B+9rJfpL+n2sIdsAXEsukvnKbWdhnSNMFkU2DEBL5m9V8+spTSIL/b49
Q9mL7ZWxoNNSdcLciq8kV08AI+cHsD2k7/dNJdGsewBoqYfGPcmsSjkDq1FuZD4k
zyP9dHUnuNYBRs6ECdaXg+j8ca/J43rEklfdu4fKgxHw7W3DicLHYGTrzGNP+jUm
dou3nE65MCWOnxzaIQhhWFbqQI+XsnMDIe4Y96PeHC4qaipLgAttoI07I2Mb9pla
oSWRzU1YGl5ySW3riCAy5b4jcdYApxLxG6g3PQBN7Hgw4oFQxEop1j9Wpq06rSSo
Xxm1vfFR9CoatI9AdyvM5MUs2RMCwTpouwrZYVsbF7jUC87qLnJLP3GJE4OvTXbK
hU05KvBTc3jXRPST08SKZHiDu3qgHXmmVVj+XfXLgtKKLAK0l8pX/KfHhU8uVpkR
qZRNCIfOM5AQk4eOu9dREHEYcRahBx9p6R+QsGAC8x46Jt9cAybUppbIbPJ1oQ/Y
4S8VAEWvcuisIJICOtIiT+fnfHQ68o9YDJwipzKbvQmTanwuBjgInR0H3kecIjI3
m07I97RDxDKfoIh5j1Al5vsk0gumHm6vYJGIIXaWYDz+uUt91q9TjxfX86gZGVqt
RIfnIY3xPP8MnKThyGKPS8Ztc7V3pOjFmrmmM4/QpCSeYS1aeTP+w4B9a3jlAvfs
k29JhvMfFZe6u9lxhxRg+Rs6uvDd5enBoE9CG26a7iZa2Gol3z0TViO20PWrIQEt
FQvQIXNhlqwOpfyjfBF5FJPnGtmlA+CJcVNCi5uijfdiAKbQsRMbeqpdCcG/8YyQ
taXv55d0o+Dqhp8sbkP4yV8l3gQzZ0rfErXGnu0QaLf9EXJNw7jZ63H9WpzLOWLQ
8xEsOupR8WkeJDhxEmEkhJFjgPAkK50XKr4itlKT8aq3OlkFH7mdRRbfjR7c2a9H
DebCFE2SCBdzfaNLzLlVPlUn9qrM352AbVfG0sEiQlphJp5w2W9wl5bBPRSORoBX
43sDFJbv+2+KPzSCqYHQE5XfV2QGX68C1/RvGNb8csw91QpDjXaJiEizdh6jNMAQ
FvizXtD69ct++KL8ySri7jFDAeetO0cCOWye+FI/mcPvF2Yj4J4A0sSoUA7wVdUS
30khaDopzn+ZWpHdFxjUQmRIrsJmYoiWedENIb+sjL0VsBw9oD4qz3VCQuCqzKR4
X4bUgCA923nl5vSEoM7QsTeW/9qhQrQVCTTtr/jOVLE/BoSSNQszV5tkNJKOhmqT
wnOU+lyJ0MVxf54+G5shucce9LH1bnBwq0FtGa43G7ez2ihYSOUFYcLl6tDG72gT
9S6LRblRkVes5li6x/LdJZArnxuzelnI+fgM/ZIYjoC1r3SR1oFki1ijLoIAFFlU
yXQS2qwZo4fwN1tR58XOfTYRJYxgQARYZj6B/1oq5GVmc9Sx1KY5deJswEkDKsSy
5VPutx8HqeTHkxYA6FfugktQPUbMNcV6qdiAfypibOvwLNL0bQ5zAjoe2jwtuJul
eJZnY+/st8rBgjFo4LAJJIamaBqPdvdIIj79lINwo4WwHVVCMdkMc4xbwCB7hgdx
IWkC7lib7+AINqzOqZlwV+bK7yFSJhhKLnUvFSIHEOHb4wcwZo49wtzuQrLgltsJ
xMvbXammVYev1sd4LVU9kv1RMZ7JrcpWqZSQ+oMvSwDjCS5eMb5Rsceznxd/4O12
fbtV7O/qlwOp0bUI9+oNp7fFpIcC/QuypjzxrmTFOO5pRHccZRLR3bTQTIEwFfnR
6lOXuq6FkylyPedNblSLw3GpPMBstNwWxUDwOeUXJrP9SmKyMqD1pu68trCr8Tv9
tNKU0Ziv+mE83GnX0dfnbiF33pxhCKHfvhgeHeK4S3rTRfldL6KCVbEflwQfQ7yT
u6j7ESXAccTpZszHbaFSd8EIbfbc9UDDt+B7uXeI0Wci/dFdJtQYUZ63/ZMhY82g
wTexEJfdidyxn5tHg1/OC/auub/cIO8L8K2GZnElpXvVPZ//d8JbSgI9VFgteiFd
tUCpm+gwu8GyHyo6pJk1UvHpkiz7nHk3cefUt49yZ5cqDoHO9F7BxMjYFRFIKFN+
v9KYHRB8jAcfFwk1ALYOiOOQYB7NPkyzRnW4joDwjZdFniaBzitKua8bE1sZuiZl
95GwQUKzh/rceYfQQCQRd9rROl8VH8KyBGTbqwOyC650DUFli1ujQN5CgoSLXAqD
WnWFoDzouFy4qAqOw6evn9XILO2t9WPzBjuYZa6B0PH/qhGj/dPQW/VXRigvNDe2
xriPSQo4IfNeQoFwPNNF517r9pPULiJcdb19qGnGxuNuX94sntjuRw3FU8Vhew+5
+KoeQGIq/tz+ujfSQu3sPcA0JVpaplkYt/i8isQCT++cwG0ii3FAyO08qJ6wn1RX
JOycqvYNg+r8etighOU+nkZrKP+VC663S1nk3ksLCweav0W4/HPZ8TDTpdZS05xD
bp/Q5TpiljF8lR32p7x+3REA0Iy0Hfe4OVwCAum/c0rIeEOopxpTNjLDafS5rPgL
KWZ0DU3EGChqcEonpuBYA7IKGwD9QM/Z5AZw5eqC/AUb2gA22NtHFegW051hmxj/
pzjjfGpVnrZxh9qTZQWpjfxEPQskd3+RlkzvSeQkzMkDnia6+8EVHWR7yexNY7wX
JJcmk5OIt80Ej5hFXMLXr8Z4f36BK/t8F1pdy+2recZf1RGQynfY8vx4KwL3Tssd
iGGHxeQ1jgtQsfNnRCci1OmzZDtF0qflzi/KnrUuF3oyviV7rZxuumyFmWAhMAI/
up5tMfK35idhO0SqF7URsIO3yGlzEO0nDzCZK6D/csr67h7HaYqYwN0ko/nxmlb2
b+/sABynoH9F34QQ7wkxCix7VlLpnqwZ8ehyCnImo4+uwSmcHVSSz32OmV4bdH1B
SsbR7SxMx8SdbeCvb+XTUSVOPDLcVw5/aMgxYbqhQdNHF8Wf8Hxm/vMW/HuEYV+h
z+TuNe38d+3lA3Cd9L+6NflrRi0CAUCtBavcUv551Cpi1VfNqjt3Lqb8iasmxOlC
GPdb3umUv90VfkiSHfTCfB6W+pqy53BFL4vBxlYBVY+2YDLZM8OwMcUtydMBNF7m
Vwp7l6Ox3v3SFLGEVKV0NHKiSbQYjWpql+Co9ro+eJqBTpz3xfUOxBsgr9l2RQta
t2QxLr/gCfIu4bKV1ZAwMiWZQek2MmuJfjq/sZO4rMIYKWpak2mfhLx2RyUGAlVI
8SE1wY1rvo95nWLfse44c/ClAQtmlDbIA/O+GVjkC45rTaSZRaiTaUwSfO/TI8v3
s1LJPFj1JGJrmfTKy5U4SmNP8smWK3y0JWtswSUL26r/D0+MyjY34j41NxpSEgSl
Tx0ToyXCWVdeva2etw19qGKwN4z8e9De6r69Lf7OsTqz3t/zxIKZnFQGremWFKCa
Mn4q8LQWDnt+1ikMjRY7Yj8D6Inij01DV/eK6V3sm7KprTZ4YNa5UnRNppG+0HrI
x/t/XKB/ZSzgbAvwKVMM7IYkv1bZp54dR+m/iPR7RUIg5PZTH7zyQgxxsB8awRSf
sRA2p2KfjmGu10DlsX7IpJPIKasutmPWj8jVLfTcS3c/WGsj4vbzp2XRL+7csYH5
vsejFCqRVdWLsyGJ2U2szgll8d4B0uENd673dpFCNXJ5gC6HhhpKRZ/NL5/pNd/C
dut/mKs4gxsga+r2ZMZjmFoaahITR8bnWEQUTsljnBeANElAFpkFyga9a7EupMXE
LD18DH3oiRkVco1+RKPfe9G0K5s2W2HN50klqHOV0pVYfaZtkK+MHnjgRDp8fJ2Y
xaVw5NJuON77nZCBjntc6TKdxZqQ230sNIcd6vaPIL9orw8ojfZeEQAwLhNQdNkx
h7WLoEtRIdsp+od3nUW3knW54FyG+GuIDf9E10jRjT7/+1o1eAsl0aEuaCqc4Z/N
YrDo5WjBixuYcTs8mfwgVNXxdjOV/6JSEdBhcRk4TgvbP9vXkYExHqtBIwP5dbXR
IN6haLZvEhohB7xthkEuGyQl7JDZ6zgDZs7l5R4hFuE+WQeHSYQleg9IueVxc2pt
mo17GEC2mr5JCrm/BXSXc8JNYiAGeR5dn8Pg2X0bpM9+qp1CsvX8MsYcLTmmSiN4
aoGbWjSlJv5HCj8X2mhFBU4K4PS6a0VMkGfpYIm1wPcUg9FvDuEWATSVxq73STLD
mF5YJ7dJk9dOS3HSnNShjWX5T2gpLNoIWK0wred/rWy+hrTtfphlKZM0DQzRMNCt
JRBCKX9g09f9ATRjOUtQD4JQSkGMTPy8MzNQ1yskBy18X+vn/xFYJrS9C4WuspKv
C/dsoCmPyB5UPl5D2GG3Y3/0di/bEJsCrIHznLl6menIQXrRKhdz4y5311x9AUMz
9uYKtj/XV6OJY2kZG7u/xlvDpYoROynxUEXe2DHzd0XjeD8ZNuRlsaqQWswF2+hj
8acOMtwh+y+k7mEJdXyYpfZg4Ih6JmuiH/Cb5/3AW09D+/uLe/evs2ZO351wfBPf
XLxWnn3NbHU6aDY708vTnr+QOtA76blgnBGJ1/ZxpA1/Kc7E1wK4bmXQhsnaO4zn
BlA4hhb1gfYswvdcM+4qy38zJwimSrAIMSdPbYvJE22f6Qs2vio1F/2UauHXl1CK
q7xefNu4i4o2J0g6RGLvn/GRgn+lXpFr5+rJB94cc/LTBPheNh9q5WHAPFXFs9iu
73H3MzJ5eh3ZjMfqhHJrnMRyrZHo/FsHEwtFlxygJLbm3x6Y2uZZIibu0Tkt+POd
RJGTB4qVqirQc2i5ORiZeb377GutXyu8k2NxQdhp1oxZyt6VZyaI6JXgEbkdEOR6
QcNRpf0DKEs60UoE/6axP3oKNumheoDWIOxMup+lssns59NHfNrzWYtiJrBPj4y/
xhLT2PHvnqjwBmxMJ3jGEebl+AnQyg5R9CpLOotRlQjeRbzeuWQCFGm2NFKSVF3Q
thiKw45wJjuYDBkp2w0eBnxv8NU0REr4is7YK+sklftaLxdbyGNUidS+d0yLsDVV
i81QJq5YOR5Ilu6F1o/Hdp1EhOtkQsNV9ZhoWvNA/O4ua8Mrw+P0ATvzMTZ502hM
9qf3EQGLh6djYcUqlMhhhr0sT/4K3v9twFmVzfYBGg0EEkGmnQ9xQndoR1KzakZD
6Yl9VKI9MoUv3B/ihruGppEtpCj38FtbDCY8P/eaxAeXXr+DaQoAZcvu0KeBetmS
I2Adl8QXC6WoliHlSh7HMe96czwzKUqk7MH1hEEW5lKxsmdgLVmY4cm555HxS/V+
jxelfoNNBIi8/y0dP+P9oFYlJCOA+S5Ir/rkuk2R7cJS2k6jNNKszlGQt3zRD7WN
gT7uARZ+R0MaTcJlGdWEMEattmYgxjwdazA1qz7tvh2G4aKgUvIrMGJcW7JUykHt
rS6HPbK4EC+Y1f875qTEHOKHb01w2xkkH0X9QgG3/bWPEBx9nikHLTjjn8VnjYBo
SsR3f5d+iPtWVLHWUCz+nTOGSnjsR4UQGPOzi6xPpWVWPdVfXOjzbQaHZyPaWO5A
1ha69r3ZEEXnfKPBxe14yGMGgd4l1IcjZH9YoR3An5c4jMdgPBqkKvMBJmOkgO69
N1rCaIpF9uzF5TwQKkQhTsqKkuA13Id7OoKY/5eWm9cqGsFZAcMqMMJHwzyvKYYQ
B1u3/zaYsdpSCAbrkaPk/QSvvkZkekP0stEXjl1y0C0n61WoljWGHh2KH+FeiHYF
47D5AddL4oP14rA9KfptK3hUxKGTb0nvKtiAmTlfk/oz3smouJuwH7ylfTzAJxwf
sLfQ8MRFjQMWF5NTTKWqJtcEHrTKUTFrVyfhP0feKDjGeQuS+DvQZ7Z4NBGQNnnq
2c2oFh5mLf36g5HQqyJM0xJ+vkSIbWQQraKD+y4kBOVoegXWAv3a1vJviNEmK2rJ
1LQb1l5u+lmiTz95b9pXhLfj8sH3b/9B9JxlVqDWiccYAFHwYc8fNJDFmvMOgD6p
VvqYD5BWQLRr/gpju9blIRsOgh+FCn5yB/t3HXSUPy58e7IN6VPMPqx6uN0+o2cu
jymvxt3M1q+KmmSq+KU7JgoOFYDJ7dZzkxvu1v/pBCGwF8jbFdYK84IMlrQskdGQ
vUYi+dnfOgqtcr0uD721Pq+a97appf7fFx5HP0+J/Bbpt+ry/GTT5sQGcavqwuGO
w+hUyvY2KHH1cUyvvnZoGj2v3XB3fSMR6QFsUSJgh8E/IIwFe08bWRIA7QZF53aM
NroUYJorP7vmB0GyjsCASipSBxMZDnCPs9BIqV2+xBLt0ZiYtFGxg93Nng/GHekA
+bl8LExEBlLDOEXf3XUaTg0nbMb4/cILAhpNEW1wXGKucddaWP5e9bcWjyVY6FT1
HEr1kUuGU5LldUSi64oGiXvrW9Uvz2ZmuimJHKRy2bJbxSETJ9YldsJynSuck2Mc
cVwWsQy7eM4jIr+F52UH9D7YkRbC5DQwoSJVWnWn21/7f5kXuSe/B7ML1Ik6UDDH
NnkdQCYjw7CVXsa77jm71sMJjvcLD46jXvSpkt/sIW0gZJPWANwxmoZcdXsF4HMA
JmwUPd1c5VBwytMVWQmQXs/1R7CBJAc5whPBA1kQtNvM132sC/WvcXVRjsFuiuLQ
xBoALX/ibhB9CTu8/lX93ll2T+4gPlUhFnx2CoWYN1RURNzve0Z5tu8+FP8ZPdVJ
qYH+DRNWbxgTs6M3p05ALSBIERU59wbbYlK6zXqXbK5WeSEXkZ6et7yFfDYotMhL
jBNtYzNh0G9V3I8b2gRIhjiIZs59IT+hOt6zx9+12lBxbQeockr0LEPcL3fQizAa
YekpB2x22s+kpXttM+hKD6OdK85aaj2vyhbyARcmYBOdnEGjCnsg9RGepy8lhDnp
7tZVlcWIObreWbOrANNP4RLpBafYtqlPtv0hH8xEO7CiNUr62FmitcBNIcsn8Vkk
kOrwdyZADTpbqbi7jbAy3ephKq6PknfxXjS381lVU0ZOAoZ8PBJkePKz9j3dk1aN
9UgvdWjJw0YfpYPd4Mr3+YXkfUs4ZYam0d57vUZWvzKU2HeHL1oLxwVGeNdG+ri7
mVtFfZ7EbLZz8//9fWjXqosRfx5L4nHnwHjVFSfTDkHbxo8ruch29kK8+zH6SUwL
sgjc9dMVCsrFGk9Ni7YzdQumaiD6rGypBoTqLDad46yjEWGSqg5Hd+UnDjFrgstL
hLInswMLAj8jfbC6TZxm0I2Y5Pw+9KAcFSlLwr+UkdfiEVeMa8HavpWRzNQX5eJQ
6oDH2ICwH/RksAuRN9+ZiuxWEj7Kp6gjZ/tSmVRZEQ/gfMYEZXtwWtW8WcMuf/b4
9pb2Cg+uATtKgEDftvgCTB8tVAy0xi3VZ4Tea0tjRmkwvXS1QGfd3AB6Ed3ShBKt
p4fPf4Qc/HqkH2Ug6RgfjbDmNwZ3bmzeAhhUh4pnNq7zpVn44YoOcJvD70VtPtKy
1HtYZVlJqYAoUEYFHPANOVStSHq6W5P3tsNTVbSnIuvzjwWW2JwX++QEn99M2uH6
3pBbzo4c4/agH32bPn13wojcZnQ/YyF+VZ+9U8ofkKIi4gwi6MEuqcXH191riGWC
D26uFISJiNhElMv7ZtVZJmBorsHEvIyYFrcaaz04ZoYpfab+8KcQuXjry3pIP4yO
l/MkzkaXugvkare62i22hcOCD2zVZo3j921c1NXyn1Qp5eLBL8VPYYZqiUlFjFwS
xlbFxJoLxk71H09JCY7H72C9YO1mUqJEkubxaMhwQHJXAzzztdGirL/luglfKxPg
bHE5znVe3MialU1ubXaZKfySEyVikP+YFop3tCyaX7qrGXA1E+RW2eUYW0PI8jfY
FtiZWn6CNOfozdfXlOIVL3vdbGfGtDIIb1L4NJHrlxI/ebapxEI9TZfG75ejjCjY
kibst+qiKNyl8bB6aCEFKNrZWIV8Ge5/iKC+G9FODPAX+vI+8inamEot1NP3kTgV
EVZ69xWMZpsIrBxzUPo1jz3Syb9JSoi3taajhueobXNRx45ai9bpmXlpP7I8W2n0
IyP4Mheiml2RVpt4pj9HYr4L2kYyQURG5cqsbG21RtO3xM0ZohxOOBfTuHXYMr6/
1KwmSBVwK+K7/Yzdqbefsy9Mt/d0voJAO+biGOE0STq/DPc97oZqNk42hStAd18i
dwoqiVaE9LyF2Ai1LSoqDWRLapVC5azBoq2wFt3R2onLNYIYy7tH3tsT7sxMx9zH
r9yuicuDSXjDr6JfC3gKzAXkGDUYGHC/O2DtN8FV/BfiTekQnz0oWMIWzZ4k9/9d
fxNfT6mpC2GOSxUVFdqHKYAnGXbn4G5wcU3idPr46v5sswc6gAsolFt0raE+vasw
94sUNhq+IZV8NckHQ7Q6jL0HgRhcAlhsjpO9l+RoawyDe9jSRxuCd6ATxX+vbVvU
SbfYroIpuP1lbiO0a1t0rdSdcQuhCTM6lOv+EL+mjEPELnVijgsVsX/Z3pxJiIiB
OauAYBumW8rDxjMnhNd+iTfPDZbT5EWMHRJV5CKKjNlJ3zrIDx/3OVPq5+WOeATk
sjRpjJDlBDOrst7xOd4UzSCPW4tk05oVPsZDTbewNS3W/lj7QSZDwKlSwlHQ166x
f8TgwShkF47epuBUgkOzC1Ykx0P+e25zfgnv7+M8zF9nOU7zqAKcmSA7TjBwGPUv
jFzIC9RU0dk3wup+YT8ppN1DfkICoRMfCt18dppZys8rYXX9KEKjg5Da4gVLPpi2
lvV+dVJEabkYa67O0Yw/CXkiUVSz3iA2UtX/OoVYOcjyWfF/No6iEa8xKsDFZIOX
5fn2YyNfLjaA5TxjOQei4Yq7HvWebM7eJhC3jgTMi1p2iAxkt6A67XquYNOs19AV
o9ZSDK4kqfb7h58udUMjl+bFMaim4eEGqKgyPFoti6ZTKoEZtRHl94rnZXz1Spl2
PgkNigCr+7HEcyv7atbcA3uWVfnZwMNzCpLBSLevf/uV969BkHpqy9upvvR9iE8d
NTacMh8XIkAxuqA3LqeJguuWXRGxlBAdUJwjBUSeIY8V+70btb9oqIu5V5qruL8e
4SqzcPxWwp1NOWWLos98be0BpEnyt2JK+M/Bk7BHvgQZK5GmGU1wgwHLiJqS6yJP
I+wnqxZ19VhoNWjJZsN6qoaIj8YzJxSZqu7OA3a9ZGe6Ic2gXIip99eAbWnnnMRA
gt8UfhI1hGWO4iFPZm2F5nuy9xnUTiGYFomrP12eXf/GYA2XbKPkNomthzdv2fNI
MsWOjibfzMVyQ7KjEWwqWjSyMuQnf4nprgdrTRk1duLDUTL2LBAvu+TZGM+qA7Qr
N3lQNqIS/m13vRNRTraIP+hcilU+2kJZisLeWE7cJPkCsFNKKTJUEmlhQ4QR2RyF
1lx8qzBQ0E9WyJVbwRG37/30Xz8XkqzhutSPcNQlf+6Uxu/xFL8lBvzyri3gqjKL
1sAuvw5dF6a3mDXVDLdqZGDISyxHBbLBtaJaWkuT8EQ2SoP3QGP25vS9KGo3pktQ
4J8Ekqol4331CO6JxNOnxS4kiYmAlHCy+2J8e/7vAJubdkWKS9S1PSMHvozhL7LR
7uJBaYzVkbHJ6Zhpb4wgyWudJkhNoLBqzRDsqZbCNd59QAoPSBsGwKsg2neorlly
hsk1INskGoP1JJN+obP/xgAQ5Y9UlbB9Y7nyrIbqsDk1sGBRWVpKi+Ql00o4K7md
0If7OgibtVHQg7CZTwyr9fD7qbM3OzlPpKHXPoIWzD/lxmbI4uiwxH2NNgPG1nn4
XVs319DBnZ/NjkZMFJkgLKb9WbyEBeF6BX3Lnqa4a73ZlZYFonitc/2g+lYMtj5v
pWSMaoqLzvpTADYIKD+f+xrtybYkKMb4DwsXD5C4NXmGfz7sq2uuRmE+IPvHmK0m
mUktGCAgtEY4+t509xk789tEQuEqfA1L0TuXAJZ7Xajk3DUxWlNzsJvwfDwGsj6m
F0PxyK0SSeHJDOC/qGTVAFsI7BzDVLCgbO29XzWacxXN3tWDTdSwY8eAEOLC/CH5
/PlbyT1QZZ6eUGc0NfTewPMpGhB2oMj60dIpi8fwnazrwaV+F6/elvduTGa4j9xy
u0A5La50eO7TNGYMm+nQ+VXq3v13vjlR04ScVSy9uX0oh1wpP5XlGyPTVQyQb8iT
Gf5JMpoOIcfYAOxTVb/UJ297KJd7sKoIboNjSIsCJaOzRO5fFL7CKX+ftVP/+wrv
jvJaPOjokINUjUaCVKAirIUjoIOFZUrGUc+kYvZt/rnddiLkKXeM0LmEhk6RXazO
V5yh8eJDL83rOA2PkkRzaEurOLkZ3rAHOE+x5YyCF8YOKc76lxBlYafnEZWw47Dk
2bc+mqX0ZFPrl3MUnMa8ZgCGfkMETqY+tciQGUBhSNLDpvBSS3pO/zhMcRDbql7B
HqAlHrLDlw/Th80qRu9E3Yn5rMSlLcFT+8mPX21OiEku2mVQfJ8vrYTcMkn5JDFM
5aqU4ueDhIDDWE6NVfGqVIM+Ocux2Q/wyuI7te4ygV3Jyr/U6uV5O4HZ2wieP59H
ZTUYj/s9Ie4H0tvgRfI2UdHraMv+v5lMVvl2He1piqZfy/OrvFOWUus4Q6bY7Kd2
dLH2XX5q9VjYTSnzpLXXJr3QOGgzOEyqAt63oyWGZditOVvcmUEE//boefD0kgNr
0NtKiUcEBdWJA/hJs8k5wR80TBELVTXG6PUI81WD8D+dcYv8JJodRtJBmpvdnsYe
RSv+/vQn60lTr0toClktgROcJMlII/p6+nYlspicTPKvBiom9lmGCNFlTpRpLA0l
So4dhiNJVNjg61TAUIIyqOVjrGmuhjhF/4OHKxaQjvLiFwbKj2LNV2dD3vlxTx7S
iS0C1yciVpKikarVZ4gtwK7qquZGwJ2+gD5UewLdeQGjVNmipLN4RE0jfWI1MGBy
L2fjXwNJjhDVmRY148/BLo94eaRKAlWt5k1c7f7L+UIuzKo2CcfABlVWTkFTBTHc
TzUMZFFHbrVzmH5UnWilmJ29LuMAjufAjCkhOBYWPS593fX8w9DGIQ689fE4CrNx
qO4I50UYzCUQ2RmJzu4YaYF+6dwLP0N7BhtMH/Q/CmuLWRe2ExiEdL0Tj6iqTTK/
1Xonlwc7ng7Wu5Aay5TPUwgUUA2PxPb+FKYx+tm9SMEp/12N44YoTM9Z7FBusKoE
R+Qigdjcf5z/w7C9Ak+vuAF8WgAY8LRCc3OJ/Me7g1amTT1rxRKybiyNkB17qN3q
/Nc1sSj2SXj/XCFFy3+kt/cCP8INcgfOeJOfZ6gsyccOuFxyO0XDrPIYDiumgwAs
bkJz+CklRDgUKStEqqvNcD6LJl4vNx2T36bppbhLeEWh2StAz4XpE20MHLRvKmtB
amdufCEwWhqoHIk/VDTa3QvxtQyBUdwn5wjfJukL+524MpZJFjfYmZAvvjYTTlbh
M+M5Fhgv9LfYQbgkBdpHdTesrSHgS03vJ0JxJAhhISpk1aZjrDAaZeK1ZZCqYOFZ
bOC+8KnxLt/TpFp5mRui8UUlZM102ru1B2bnb+3iDzYd/Pg4iEu+lSCNgW1Afhhb
sqEeoHn6QRroILy++UhpXXaCGudacxqHqV6E510D4rEaHYvNZYZzYAwcEDvpqQA0
kUJ9c3VaV4d+H1tD46GTRlLelGJ7A4kvkkMDBciBBfUHujDRw9RS8b1vFNwg/ycr
Q1TLCghRnvEah+IGP32cxvfOsSYNyO6Ivu1nlAUZg/E=
`protect END_PROTECTED
