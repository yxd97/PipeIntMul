`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tUOurrowRW7Tho4zEJZQ5/56/D6k7KH/Peku0dyINdyYSwFnC8i81LK63qJ4nv4R
A/BmZErPIk3g4coB69kliljdde1LFzzvuNiVxSv2G9lPerdxVijac/98mn3RUjRw
mH/UcC87MdRHCSYpQdrPOL5nCRL3srJ1Zdt6+WA5NYGYJ/7s19H2bfrNsIOEP5ZD
FOI6bVUuu+gQRQhZmf4UkgdxDgGuI6bszcJ2unm7lJNIrPpIRr74fbkk0/o+atFs
WVIBdF31TrimLnJkoxl9fRBgnP3g7D1tr+54JagDpKOSrhL0folrRNwoRlzi83lJ
oS8XC+iHOiBdyIU6uaE3I5PSwe4aP8PnE6geXxBiknDgzO8jhXtOQ55bz/qrfU8Z
O+29vggndFWSofQF1qU/GNxyPLEn0BQdhECZqOtI+rtQapa4V9Mt2pwG730RumgB
VmoPciwRi4B7+PuDlgHtaixjxnDEN0TYAuu2lVvyH5BG0deVQ8cVkZT/zL7pI/DS
FsI9lDSD0gRDTlnN8vaACZ5VNP5ZiQPo+oLUDBPNR/lSoKoeh5bfRhxxbaeWFaWn
pJC50bvmE6ksX0e6J/mED0aWiiLMq6dinZJ4H2WdkDKj4IML3zvToqCstyb2f5OF
961gLNBnI9k+Q/Kuy5hqrLa/z3vTRf7kPltsx3pJ4TeZ/nZX+KP7BKF4pdI1bKO3
QOX6O1ZEBaTJgdJmrG7EF3GDdeUOIu5qdoJhJEdWQ/0+Ks0ku+rDJGAQTTGShG6D
85Sws3Jcok+RvChe4v/X8Ow+46JFVsgQg32LDwuFMuKJQL9/BUx8AxLlJsXxN/Uh
JVDIZcyAuzANlJRoSnUkucS3roqoHIXnHsRkDL7byhFOz6+vr66/o2uVt+Kj5MkS
ir5OlZy0UHAZYe+IM6MAhfUlm6Cp026dsByUncekK6hywlTyANP5kv8ucHP9wpEH
PPevAMzZoVwMK6OXD1sV0x97ntQPfq9lrF7rLHYHI5eMoFLl1yfDqoy4IalDkRAg
WRUMtO/N6rm2aZ4jkhFB0nC+kq3f3JQphHKky3j74ZFDlQq7yZrO2uxgLq4Q6oLZ
sk/7YY4YFuTon+DDcMex3FyPHRtQeBFJNZQxkAR+qwfn5PtKLHbyRg9wwNuZ4jdp
l1UTalJzlYcBywWHReqnaVZqjNOOJ4wC+gsRXGqUAPXSvL291kfoigCi1BiqBiF6
b2vUL6OoDS5eoKWdUTgNco6YmDcL0oMYinsXCR96wLItU8qXC2CzkOv1Saz2dW0N
kOi2o2YxSH4xmqeoFko43DmE6vfQLLwwFkjLiLH/jcWBPoMOO7S/PNd2AQHHIwOJ
rLj6zGuaVfv2ycG5Fud+Drfa+2GjS/mBKXkk0zbmI3vPSfb4QTxhHcELzpSZmXzi
66vtibn4DIqgAuZgdqeyGEW/nWz+IUwOlXHMtgLct70QaYGuzhZkPk8WOb6u8vh7
PmPagTLPQtdq8gpcHxFeiS/4IzEwj82d14qYP7Ff3grJNY+60Av1zODk0ibQ7giP
2ERC/fHpAtxAoPFM8R5RKZneJCngBPAE1Xh0xHwG5fIlm1tuVLkZOpqunxX3guzm
LQ85QSi7ptBoYzpQJbiue7g4fMPlOnYsHBNsteCNa467xmnu6HgcXGYSdtWhXFas
CiEcEkR8WLrvxppox8JVVLVzFotT4b4C6Us9Yc4ipEvHFCOM3nH+zuo8iAw8Y8/O
lNSj3q+Dj7InZMLB4W+jRLVXFERWHcZkN4qNR/8YUqv8elRm1T41/b88PjzmWDcj
ZczX0Vw5Ei1DxVJANviFCqMwKiEibAT81vPB5EB3Kc1vyAbxbiHd/Ky5+aXtFjRj
WSmiC+ba1oYlzWTbIiyUNYHvpdhT4V6vMbdyxrWs7X+RGcX5ONaP0vga4IJYt7jb
0L3Swu/Fr+b4RVLMGasiiETKRjksbb/TUace+iDQ122hOpc1xFfC0Anp/fq5+W30
loSkYkynTdwT8Jtb6JvEIDS65Sdk8gXcDxuhvtjDnVsWWFinZMhV6ONQ4WIWMD7r
HzgDPAdBnMR5BZLPcKvJ6b1DQbUdUNtn86SXdjwVK3ySFyguFcVZj3Jl/Ale6DuK
WW5XpYdx+Wa/Wzc8Y2I6GT3EgdSlAhrBvn8EZhnHVfeq/GYIwmMSo7G5SUfZhSvY
Z42rBI4MIcMGuA4fZ3l7fPQiZT1eyp/yqccxta90KNl9preQcD8XOMgB4CRZFDIa
pm81tYWy31ajEQzb4f/Qpx66532XmAKQUCuBhpGLM39HpC7WEUjItZMoAsoK/5Gw
SZe5gkwm8D0eGhoLF5k5UeBYyqr3umujylbmp5iF2vFczMc9T2cBieIqAoJeim4f
mspi/GzXgk7FqOxMCd9R1tCk7sGZ5gic8fB6DbcByA3XkDKW0GW/yHgOjEROhdX5
+i2WitCYlchg9mS9RfIGKKpMYo0SUT2M31Vej5xhQvk/gkc+oBGimUI+n7t/hotm
gF3VG10wecxY4sYeg+jaWMt3T1qvnUeVi0d2nEFe60O54UI43Q8TvurzArQi81RE
UBzmNKr/cQc8RI/0ajBkojaq4t4B8q9pDssK1LyRy+Z4QljMHNz94whyiYN0ryuF
zXLoF2+mQ0PuDnV6wZ1ljWYvE8sug4fKTE2ebDUvATs2kHfupRM+wQQvpcjCutRI
zLuip7osh6T8zyZA8MFBXrNxBGc5kDerk2RnmWIlXL/mqVSVyAhv+C44EDP696f3
wFR7OvppFyDajktj28/PGBZ/JR7YZ/3zLSxYZfLqh/ioueszGtdzWjs/eGYJB+NQ
S63Ysjz9UCVNGXL6oc+zkxcggUran5MXc9SuexvFUjr5oJYWCaBlPAxQooNDiU4I
z3pjIU4ezhioszOaOzbW4JuXcS0WIZLTk3a2att0lJik/XQRK5UJclOdVAkEeulL
KWq6nUHBTRnXis657LeaCYk1zpvZmkeiq0J1HMAggoMrLiZA3u8AFEyb9kKYQpbv
Ja5lBhekY675+HUb13j5MPZm8T74qT7AKrmGrlMnhPFOrDNCavjzW2WVwNx0+tUz
/mynjKyCESsyjd1o5ZCVBhJtPpjk4fsS1RmGmTNoyV8edhHnzmn+cYD3kQ36XKDc
YkW1buZ6HxGE9/mj+MCsOvrRcfwLjVbQmPFr+yqu/qh9rDNbsKSAkZ1LxQo8dKKk
TeAkjLty28KBZFR9zVgCshN/+BnVfdTZhurxvlCGT+Sc9KhNVMWrZm8jPa9Fp2v6
qx/yCPV00n/SHA6WnTYZCtF/cGwLm7MIxUt2he9+lT3pLRW/x3v+50zFHMouSM55
do+GfakUYD6qhT2rklRTa15Rbc6x49v7UQHqHIBOXnJfvd/Ox38NiVp8mYV8auYE
xIcpVoIRVjxc60aReLAlorwHCDWmRHYVP4ow2rGf18Y3KRbJNoD2Y36FI4TNsM0S
vSJpK4qWOY6WtW2mUOOtJmQUy7kTPyazgmqy07oGcwkQlfrgjJrHdDzgaoDciuWb
pLe3hgVcnOPAE5RYP8XD73uoO3v/tN7bvIL+RfuVnCedXsca3KnlY9Fl+X/sdPMa
B73qS77/fMYyu2ZQKzGMjxa4MDEH2Uxlyb2USlnNk3zETMCEHIyrYuk/iL0+h2dr
lKWCLjpJASW8M6CWDyzFMCTH8vsazhIPoIbik4Qkg93gqjhvhNrlLOrmATHfD+7z
q+1WvTwnTPrJhj9deXqlT5103vcAtsXNJL7R2T58+QAas8v4Xkaca65TaxdqpVT5
a0FdzQj4qOMXDvIGNikhp9EW27nlKWM8HA9jYxkEqPzzUjtVl7cD+CDE7nTp/2Dw
1QDHHYIBv48+4bI6puC/2CDJNVyp5KdGddDHrZaEefLgylbLUFMaveg39Qhpw/Do
9Ot5+IqxCiVGoTt/a1w+45bRfqyuolwKX12GTp/ORztvncthWX0Zq9UUZ7zE92/Z
Mm7JgooQBbe0dnpga14+nN8KIUfKVg1bIlUR4dbOMPR2ewfRHAk97NzwgGozYOD+
ClDiMKcLYP952uyFKXYEhr1Z+Cksd9MYuPWa1r3MVhI3F2xaNNtwENpW6qKdVxPl
VHoq5Qbb53bvlQ/CKS2mSgtkogdGEq6ACHq5Umhb5T+4sqoOGl7BipMTxHymFpkI
WGVdk/uvGHr/2wtq0a+NMZLkmHORMsOBVo/Y80dwr5HFXqfYgFaSl9Nb/v/PcSTt
qROjIWoz9fATk/zsbfpj9hD3upZCDAgrwVAtBEmB0AYnIh0fgRIaapI8nfEHWutq
APyZASaFYN18IWk3zMYIRn1ntE8VsAcCWinYAjra654OOnF4w0ONenlG3NdNAbd9
B7bHGsi228hZQ96N71GiB3l1vz0JgDlNEhyqh/PfsfcG6FFAZhXRdvNk9aDyIwaR
JkrohhS9DgaoyLFIISp45lwA2MCl3brp+GmkcjDErqO2wcoK0pVfKRrDHSfSCPSu
GdzJn4DzizsrnDHqFdNJ9rhTKxNn7498RfuZzHXaVSA2jGnBxQ7Cqlh+UXJPFQhy
kD9KQblF3w9d2piw+ZmXhkZGzafKEHVB8rBve+1Y7dYwI8yJ5FfmOcap9MPVg217
/VAEjt/sVSBMcybNDrEb+anvfKOpeFZTbKWkIieSZAl/AR5706WVkjJRafxT9Mhp
zfcxXtK8S4dhcOnIUNObeRVlW1vdB+DH156Oi10WPKtptFfHUUmkbk/G4inQLOcz
TdVE8HGBz0Tei58vOChfYJ/jn0CkM/0WDCtvLgy2POAG1kBz17SkQ5nXE4LFwOS9
uPiNBwmMfkAgQhieKvRRzs9yq9U+Hlz9d/e185dYEfErwGpzVgesbErAnvOm78WX
wP5Zfw5MCEO1OEM++ii33mQaKLGmPFBHf9uxt2HCFb3i61BmOSaxZ/zcyBX3EGgb
LfShvklrKT7xQj4xKHJsHNUx9oBB8rR9SpyrFdUEDt0VJal648EoFHe6/wzXS1Ic
o2CB7dKVwq4O0LOumckX4cvrw20OZOpB/7eccM7J8ce+/wprTIIrmK02T85S2hQX
njhfKcjb5xr7YLBzk+tROjSDVajZHm3cGYb2/U2aRJcg5fL5SDAcmX4BFtrCIRW2
mnB3GwXTfThjYeCwCBAQgmmZtvnu8hABOf7dQDTQtG8E94p6rHb0u6c1fuodE/IG
ZJ5w62Po4mYbjlyU7GB2XfrVfzidRnC8Tqv2PVdDBv2hFczJxWHHU68Zb3g2S0r2
inzOub+jAx1trBL6VeZyCe5V3QNgA/VkQyzE7a6EYEk5LHrox9IuzPIx8N32jsJY
b2CBKlaP53YPMnvFQZhlEAEntTo+J7lJOSKPyextdy4RkXljzH0EtQEFlzrVhVSi
q4adOdupNcJ3W/FwcF1CNA5RmYuNRjM2PZGqpO6Q/Ko+E0MR2rJp1oqdDU7xvg8A
waDtNjat7YJsGTAUfEjLfjV5kuN0hciBbiEjDql+Kq9GfeO8pJly6zJKMbDXMrDS
X6XAWfSQwUxVKbxbXKj4ebjEno5Zsgq02tp52Bg1S2m3/eNRbc4RTOpIQMX4iYvE
zakLyAyzB35E2f0YCG2Wab2uJw8ET7Sfyo3lRBY0UyW9mNJsDlMUIOremRSZTXsf
0dcB+yaD/1XGKz9lBmzawUCxdEGd6yscNcECT/kwP/NqNP5H/3ztk5SrQBjljTgC
/YBJBUKiDZAzke8gADVdwd7s9KcOOsTO6fv0zFyqAnjBHL0dowjULBNcIBkpLuDv
A8lGXjeyAS5Olh0xyVZweVhK+unFY5/fAHJuXh5VHA9QhMifP7kpaVb4B22zW6L5
B55aJ3WGidUL4zujdGfemnDBN+AzisG39mZa7KBdf3XDK1P1bpRRnpG6ve022KsQ
7gI8y6la6cdkCdyYTFd2ipnbvjtHseGFnLLJ3ejspZotvYy9lPi77XUsgs24u3XE
dItddveeyChQDMVVpJ3GihxZDK9vrkDQ5eSVGCLPEAQcXw+ZyB+pESn9KPAP3OG9
3igNlXM4G/B/MSESyIhQxnUOimws1Kl3Ek6Hhy9vwxj2MXw34kgEtpu++JXsbkjZ
/nQLVEB3SIIGQRANBBmRfR+8yNAASjT3Bi1PrOHX1X6mC1/AaaFo/5LxMuDSRHzA
2f+i9aBp94jn1Iw3HVELdp3H9x0y5Bjki5SqawANeXKTHwO8OuRZVNkPnKi6Dhw0
hz8eJfP2IcbC/tOb4miE9MrEY7yXCVXcrTEDwDHrgLUfeJA7WaGWyhW9fXbcKuxG
f31W1ux4VM3/moCy6KHY4oqgw1ve1y313yiciTq0ah2LuDaXqPeAFwfr18C881Tq
2Z3RON351maJ+JsvbyhwXW6BY9cbrjnxHidmvwfYFYq22+f4tdYl7kYJShHI8AkJ
SiNsrUxHhSayh7/169Zh0JR2uK5McU+kWwWwcl2iJtA=
`protect END_PROTECTED
