`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DC6ZdXfyFHPRDrJC0oIyuYlGi+chUQbPs4b23zqbMIdvwf6F5qGLC4pQWhP5gd0l
4PJAqhIUhTGRNmD26VGzKTcaP+6SNWJu4Rxi56lbIGnmU5UW+jfnZHsJ1e9yQh68
kWIA7TZVk+0gt1r2KTe2XPF8Sg63KowI/k11RoTmXXlGu0pt0Li4NB4nFcRSw9xX
UKGZV2XXGUafxyhhUuy1E27A3rQGq09gKBH9vlULpjDzYtSsXYL43VrGB7YyI+mm
UxviIsRw3OUwDtuH6lDFzOosUwhThRt0YY7f6+gWLlYDiKr24VjNENnsDBdjUk7r
S6NYsiwq6cG4VJHL0HssYjnPYuxuJTAbH88vGeP/97t86nTFXJqFNsejOWhEaUmk
47fWXuCfp/W4BOw8+PjHbgZmgohiDTvAGnZOxGxJebO3yaJv3dxJK6nhxg6HYCeP
Uzo2XVuMKl6qNiUwO/jUMhWQw0x0lU0M1OCeA6qtu/0ViXMpMBEa9PnbKrR515s7
Rn71SrmmA5MP7sOVOUcOBx6/AkMpgEW/5IA3V5j0cC4TGVltYPa1ycWTpMFQ4YGe
+SyAtr8TTgIZFzexQb1xuTD2NVALmDiiohj2IjHqqCqZ+QTTexlFvf6W19STqXqZ
TFRolRWyBGV5LmmQATh9IvFT5fQfYmU3sr3M+DvDg5G/1zqRWmqi0nDOF90wjsRR
D1FduGy4Df/MJGwfy41hMMIKibioqsC0cyC8emKs/ROLYSrEhyELNKx2Si+0mG95
aiAEjC9oPJMJsnTwUKREIKYO0pXIQp/K848CKEFxc4hNChmscCrjQH+jwd9L9rPI
SQmCjXKiyIVA+BBbu3nstGfi+zunLsFeqPx15L07L68=
`protect END_PROTECTED
