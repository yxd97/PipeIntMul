`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJ0UY8mvmr/ukvYIWAOz8xcuRgWsEVj/ukXijP+A1/IkPvdZ+aRdyGYOjC7qGafx
B0AqdbRgVm54djbjrLqgbrbNNeVfr6D1KH4vy4AiYmAl+nLT9u9/7mEZS0mIXjfE
kp4JMBlMCAlTmHYXU/q+J0Eel/uOSQjoGb+Kd1BoqSrkC9LcgrOrASzLRvf+R7sB
j2t/u6Fj3v20b10e7SBvgZr0Nws5ULvZvvJagG5qlba0/fmjN3ZQM3rydPVjsyOV
SS7/MLqqf8aUtwvqBYF8MtXxAG+2v0BJJIhPc/i0WnpwQsiksgViS8R4/ugHCzX9
Lxejr5sl6LMHo3nm4MNYMd8HgO99JBC86knhM2pB5t07JEU9TmDOtEdWG6piyHQk
06ys94ja2/Pw/tdtZwDM8PQsKJlyJIc+VTyFlygXOUEay4z1zzc8nJ+joGe7uVPG
D3U9FoCx6mAkqHfyQXRXpAH2AAXrPV3b6r4oipFocRQtcKWwZflwtyKCCGwjHH/G
H3qutu3E7gr1thJPEX9DmaXudSj9IY0tKBlzKthsjJa28/o0hokzL69FW+8iezUH
td13M0zXgTwx+mNDjeEZ/dIXJlMSQiD1Wg3FCczm2PaKXMcoS8Vcy18FUZT1nFpk
Ek6nyajJyE7UfCsU3RvfQ2mMQGDfAUv7sQ5kqvKN0DlTZHcBNt5ekw/3dyEyW2HP
mx/SmcyeotsU7maZ7zAxubk86oeD4c9ZYn0NleK77gcxpFiR6Cp550SJO95Dy60w
LY3AYElUwroGFXvhYf8GqXeCbO4Zx5f5yWrvPEpwYWz27A8Og10os75169osS3su
9wxhYXKdGVccTwW3CUXHlTIAN2IPRLdareiqE71mngiSPqMtH9iaxNSQucy1x4gx
W9ad49MRPbw3eFSVo4Vn0czUeuvjP7RPMah3dtDwFWR7tXg/FLAvyX8bu7a7Q43J
`protect END_PROTECTED
