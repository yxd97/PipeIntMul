`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxkIbpMCy6RgMz51AMn1hrTCR9+xFqkGUotGExvxbLU9CsR3MdK0oASgHKA/WeOT
LMSQ/y5d8MwsXchXjV7KkTM7283VhZ+OZtZwlQzHgzOPfaEvoWtqNLt+iKX5xuxJ
mtmA8BP3BorhqkNUTzPftNjdtJoKx0hLfV9qrYTp0xXN6p+NBA0hM/+CtTU7vU6L
rpa72Vr7EbjY90tRvo/ZcYRjZumi879hixGL1nmfgOvSBuU3hAXLN1Yvhx5m5Xpu
+l6x0OmvDQ835MIY5h6uoCbjefcsunplnUwlXugUkymQ8JGdqisrgvHijTqObTOh
qYa/Tjy5FkHehdxd6KpCbnFCbo34iNWu0p7QZjfD5How11m3GCjPFDAigrb+LEEp
A5Sv08X17t8T6eDRMGSsjTkGUnlZpItQ1bjE5Yys+2kbBPF/RzFYIWTk/KjFSiOc
InZlEuXnnzBjJLBmFVKrrOz7Vb9V2nQpsw2DhgROLl3a2LA08JRQu/oWt25y0TkE
I4KSAxxefKhRSwBe2VN3bH4NRKEDytDv04eQU9+/W2qKQoQtBDRgInn1X/25XprU
bQANLVupeN5rlxOe3qUYm6fVJ65g8pxKzMyH1iZ8y9+7dahvcLN82C2SkD7KPlGx
xqVhOL8s6yyN2EjEzFca/8HPoJOsLeslgc73aSuODvxGeuyqLA65dj744X31/bWj
DMe2BgQ7Ga5Ldjw1vqArERgQ9RQpG06ehnFcBPmO7VGS6k9tODRhd2857ctYB2SM
bJ9ekI+2A2sSy3Z/J4lzXIlfvDjPtgkBR/zu0TqvfItjlpgcMgni65qLSjO6R624
bHBWUlkeDHf1ETaX74ZYr5bAAeOW7Q1S6fUo1osrvzwA8T7H+KodYMNqRZfyultI
l7XCVCGRxvf2Iep5RCfkoRdmS5nj/GFL93z1L2rH4VcWZ/mqubzrj8M0+cvYvef9
RnK9NHjoQt178RLDR+WfPZ/uPFqo0a5LZ6muNspDB9bcXCpjK/rvBI1JuN2B6Vn9
WMMGiz9zQV2qojy3+z/HXsjvGCJ4amodp3Nfi33aIQBEm93P8wqj9Jax6H9vtwd5
fCJnS3LkKxvMvHB78N28SGeDz1eeiq7VbDz5VdPL5+9iONcFt8F4/Yn3sJMW5803
sZ0O6KGW45Su6UKLYyGzVkYO0jX8aQnDzerinsnV7qARSyu51t31EtcBoiI0pSMN
snNN6sCnCjEZAbmqhPDDOnqHKTjaoye5MzueDu9XbFas4eQLKwTZXtRlx3Ru9CtV
eDRHZLHMYudc2oKBEuyygXPshFiL8VHsnZ0nEOSecZXlTMxWde8J1KpRnR1pEasZ
c/WYDJIEyawGgKEYj9MhFLONjvQ2WERtmbPw7HN4MLNiVkIL2iYqqq6ACvrHnsaJ
s0R8sTRiSSV4g/HpuizlLd0Yl4z2VoEUQizrf4HgSfP54QtQjkXjnDtU4eV8moQn
t2LjHq9wQ68TfhyaoNJ2ykm9Tl9WAAG2QJwEEjHw4SltU0bisgVOxUzPAuDVbyDS
cM6NcWBzMEi0mfWo/pz7LJqvkx2IJM3ucCL+jOaJrmKpUiyVYjefLDG400cRfmPH
gyudqL4GfYbrsUE5m8+kC5vLq7kBhfv8bOyjg0GQ0Xg9dc7TGlV7gb9NUJtMrkrb
en10ycwEx//scuJLXxIuNRW1EQ3Thc4FRdqfZDh5iuH/0t6IuwPOQXm2aiwrtviw
LI5S8b9wYYemIV7YLORsxSrks5zqqUnSSZ++x0p6rwzgiM5ApNX/b0qPFy1ZnkYX
8dciEItByZIkBeu3nLr4BZg52u02raTukKOAa4ld0MR74pmvIdZG/1p8c+TvYXmd
zPSITAOMJSTZFHb1pruBuMefHZz2lF8VXxT8CnrczMGMvvcLrg2GnO7K49GPqAzW
lTyYy9fJjizYs2H+JYDgUwp/Hc56Nm6y4F/5WYNhAH4jJ/yo4Nte9AG2EXeVrQIa
YI5K/U2PhV7bous36gsz+0NksyWTwSuh4udfeCF6jHyv4qZTD2I3Bq3MD07xP9yd
6t9UtyKNq0eUhyuUvO+g3Zj9OTI0pPBQAng6wFbDiSO+YRJMqJ+5PKPYd8UJv8Q4
wa649bTUKCP0Sd2d75r/bCUXI8siy4MMk5VsPI0UMSlyUYYMBPSEYx3Uz8SShi3l
2KSuF6sjnpY2K0c/7wUBkcEL8xGVSrhL3EcEZuJiXjs3goKuKW4VY2GZU318f3MF
KJIg0PGfKRwO61lMKFcskvgK0eVr4FOjzS2rhgkLeokTgYNvxcnQZTjHLKlf98L0
jB+MY1MUa2B/nKGjjKk3v5Mt8XD94krmO6pIq3QDuZtDpygh5uni0xSLqmBAQFl6
NE5sJ1xCKR/IEwNDv/KTyMHBGqHSc8nInGsNu99SJgwl9Xi2C2JGs9KpJVn0aV7K
/uuVBvYhd3m+wdhS38vdEdV/JXXB6wv0a5B0oIa/aXgM8RIZnGiJ1P3ADyXWGQGV
eNlPZ3Jpx/lRKvK4z0BuRfSnEbn2DZILF8noxLFQlOKmD+atmFNaKHRy4akyL/pd
CsCiNnibmNlr4DjVLV6E2zXbuQ+fTBRXGnJ9woEbyf8qlyHCypNPUxZk0H3MYzOz
m174xaEvBYcT/a5zKh3/V297EtXTMH3wQr8tFBsy6yXM6bNJz0MAZRUXxa8KKpjn
xZTGrX/088v9lsF1En+55evjj6g7XwIUXl9H+j0BxNprQZUdOx6nSbTBAu0aRgym
IN5HlU7SBYXnLGe5pvMJAQlg/4TwqoCjSHcSGit9DrzbCJvpEkWva0W8nPo4Xyse
gSY+2YlWWghCNAUTKWE6zTw727uya5F9nKeRNOyO1C2qveCUT8zC6iPvgj3N1FJm
AKi8jh9S6imMCLBy8HfivcArDKT0wAd9kaJBoaIDFU9KdVc/QBy3pWyLjWbuyPCA
CK84vcsKGI4HjzHtaQy3MIxLywwxyG75fm7maS6gV1BE+iHbXlPyuXI4BDYI8zqc
m15QT1RiEC1QHoITmkBy0+IvlKSMFYBIoJSBrrO6jBi51PpQGt84RXBvQrXcl3Rp
/86IN586rQvFWMkUpV0xMdBSw8cti4ZN3UOcURFAVDZjxdIZjpdZW5/H276Ylr75
/qdH/d1NMOOIJoMcb+dtJSehefSallGbQeLk7YkucBD42LO/3+x406HbN84uzqhH
/KJA4xoiWGLy5fsdGrgBaFzrWpKHE4U7/YRzEBHuyomLzJW+Da09u/Sk4BYY1Uyl
atYptaIG9I7W/8gy8V6K9/v8ZXjFh+rdeFty7NROQdRulsXCFMz+tF2JEwyU6tyb
QJ8INQd6DlLTkXIv/35Mb7TACr4aRs2eiUt8vZlZKYJxlx8X+sSYre397tUH6enf
/vdQp81/CVILt//jI0uXIyOO/1uoTyBl3A9PW4AaIygTbiD35cLQ/DYKbYHDU+Qc
CVhB55exwX94Dx1qAQw/fDFauGmuc6Dg5Cucd6PAISDmngTQmb2NtL6wlY4Hzh/z
nYhXVmifMqSoYDHABMxw0LB6q8kKTOhKqzSrPkiYEaRo4xcqAvs9ERt2Dt+/+bW9
8PLWXPJbAzos7kK1aNgz3T5gWs+GvTLkkDigyuZSc1sN8aa/+pTBUgW4I908K9QR
0Z+YVpkXOftUNwQixJDzf7g4+f8kYH38lk9VkY0nBWqcVebZECG7rHRwIthxKBt4
BxIO5ErRA/yIf9yblEGNHlHzMpf6FgAewLK+bHICyuTgA5U5lym2WtsHUN97IWEJ
oo+k80E22q4BbTFJgBEtsSJgNHJmd/rjGr0mNXftBseDOYMgF0H6rudDF8C71RP6
5cqffaEIKg9zfxsNpQoA2Z5e+kDqYaG06zYc6NtK27zY0z/2XX4ri5ToyhS65kXV
1rVpqxCE1Gmt4kjuuU200xeKCYoEoKZj3dghQ5AK+7jHQLGmmAe9nsyUrVO4i+oz
yVvNp53RmsLnjQIsoxJN1QSARLd7MNlIXh+RbFos8CuP712o0ws31HTSJVA9pW8f
5UPdbcVgz1q5l9zmD3WFtz4hE0vttHy6jrbSHS/21IXJSv8NorQwljt7VEJ1PIZ6
oRb4tlqL8RPCwPQxj+YjTRGZTVjP7254rIxXIJl18mQMU2YaOaZZA7wDGxnrehwU
xH0mtqrYU4I4e709IOVJuE3BZvqBI8N+moW6RX4RjkTRxzgvO+t/5nCP3S/zGLgv
/K4qvEZ9pqo9jeRb/KOx71iikY1uEzypZwg/xCEpVJ0S98kHWHDskOW6TKZKJEw8
08tCmKYDDdWjt/bxuYj0CBPnnB5CF6x1AVFsXHOtKhXh/5dRvZLBezP8ij1iUDwr
6p4n0TsA2YOYB6sEiHQsPh+rJe39BEF4cQaTWKFTYMun0cxnoyNooo++wYF1riYe
29G9qJVUDMQH/DcMwQYY6nA/S9hNyaf5HpvJxSz8BhFOtyVmLTlajZ0YZXwebklR
YZQ7HfHKmYKbJ3MAOXuo0xqIaEjl7fWzfZYHvWFO7QjhCjKck5d3DZ86uzsFiHIH
Pe+Td0fZJkvFpvKPMBaMBK6PyzMIuVhcv/ckG5NJV/tUMhoXZ77YqOQ+tLmZPAd/
WKlimkgwYG6UcdlZgzxWHIWbG9bVrJUEEz2SUhN572hESTkt/fGGW0rNEERsqTA5
j87SAQoB8YLinq2foR28eyqgqyb6AVBAGvD/XOzo+9mrsSiLVhNht/r1fcVCZa8i
gafkMIjtbaUmaJSi+fZIh1KL015pTxrJNi7CMnjyzDM/AlXZABV926n7+KPvPqMP
aeF4AYi8G6upvLkAbNbJDgStAtL9OuJ9FBce8e3Cl7najc78L9pLGivcCWiLV2hW
Wp2B+ktLDvDc2fpcy29fsCyMnpTbp8u0p8njSwz1AVGetEYmh0vrVYlPxfT/f8Dx
IkE90q6pwRZH1t1wUECQfR3Ef+LUObyZ/tQ3UR1F2eJnLByaCAH4ppAwT16fXJ72
IVQYj0gLmCBkrE/s2y4TvAdCoaHMAkWZrW/zaSwPN4qQajAmUlMP3EgZhISi+3D+
s06buvotHuXvtXF4YD+AOusTpNJwqllpgkwxdg84Yce6owoGuDi3d1TsL/Do4Bmn
iaX5ykE4WBsfcKBGdSR8OotAoX0DOLr83HIFA57qxZUh/5ki72Yt5RA9BXvgY+AA
a3Un7AGzMxg7kDvHTCz2GoLs1NSeOGLREcxXOjgsP/O/5RBzoPMdRacuXNWLOpKv
isB1d9ZLh03h5P/nri/E+LYd15oa107VLrJ3q1H3RwbaSyreqFRCf4r207QIRj+c
kfh3elposh+fCvHIRRgv+Z40b7dIyz8L75JgZIdpLKGDXs1sgMHiCqh8lRdzd3Cs
3u+qGe+REdUrdF1QPzgRrN2aL4ht36A6bTgXKrdrIxbzkTq/AhiRfiyR0N6BONVq
H7ibOzyHIvi30O6cqGjIBbEweddYwl6w4Q1pOQstGSu5I3cmsbWGu0NgVYp5vZEK
prnmvrGFY5YvjmoGDRKZ4MBzryyCZjw9QFA8zy69MSL0Cry+W+P951YHOHwZEzc+
Yutb3zC6G3v0m7D+4bbu+nPAWFL28Uv3QMumA6fgM0ev8N+C+vl+2BMuzzX/X9P2
wJkzK8uyIsdu1neTR6H3STfI97I3M6LCTCtXPZqxuGfOI21zva3ZjxQ7KPGCe5lE
epMcvmcrfaBTRuX+hqSQOiY6AlepSFHZy8DHObcuVnLXSj/714J8cJsDJ+NNzrNX
gX8KQH9mt2MGsSkGf2AnC1f3gVRTBDqvG6+WaiN43lnY10Zo5Md92pJPDQDOTLfR
1A/Lw0IcFheJYwKgD2NWBQvyPqT333BcG5IzaBCOVDzJiCc9F0PQGNDvZbsiI04R
iXd1JZZHP+WlnGDtiyM7TMJj3nc4fjHWO3nJ08HkhlOnTF9zy8nw+/HSZ4ahIUJG
gT5QnPUuYoaBQJnit0llSWMEiWn0w4EGM+V3S7INcLSzM64MtForRimG8xt/OBKC
ATk8uVZiFUjn8xeobfxhGtP6d/6DaBOOV1qQ192wiGL0teLOskOZbR7BsHFzAWYe
6GxiBqTu0LiQ3xtKKdQ7HbkRvPQR8M1vbODleRg+Wfmq0TFTL/PBY2otkEwt3Y3Z
qmbpB82uVg7Qu4vvFsE/SOLpJRwlWajvaHA8bgmcdnQRRDbITUijdkffYNH5ZRSu
IJSQ/62Y8YNyWEObXLBGEckZGpAOcElAwZLxp2z10r7OHt2JeQNwyHQOaZKkBNif
50GjU+NE84n7nRY4dTDyFYxVVlBRaQJwJ/8pMobVIBHtHOe2gna5k+XVMe5zDH/Y
cBVi9yKux4qP7s9D2TtlqkY5+bNsleVwU1dw6H4vxSyHb9YsxCfbfbLWGlSjHtik
7eWTjNGJYSduLBuTb4Y52RigEzaSnqbMBJPay2G6l3dQdE782P6x71GWJDKRYAj0
pr9tA777uf4OQphAbSRis9AOMJNk40SqD4xX0gHZSNmgKHOBod/1w8g3cns9z0IY
0UqA1/K9PXsyj+3Tgh7GuD8kDssfuemYyAJyMLrbSMVHAVJCPR3jcUT/LVYVmIe8
b+qYWlWZk9894ahUnTvbwBkHdylCFFY1+46fzuwUCrI0mXqwDBDPfVAilRReRIfJ
a0l6yMEBsooraUvv+7LgJ3ZMK3Jjk4/JXDtOpXfZa9SJAbukk1mYaZ3O2FIu1mH1
Qig8+LaI6vfM2CZ3DKXtPtWznJiMATVmFUgOJubXYmtoreNgAwaoEMSwk34ukVVV
V2bknFCgqvbYx2YOwVf1l/IMI9uXEYB0NsyzTHlAAWt6u+1m+1Z5oUlRZgkPIr1H
1ms2+x8wwotvjDckN90MunbkVtQWJbHFYk11FwW7F56kPEmhDJKvHN5ud0n1z28o
9QGCvFOGYiHGX/jKgbZ/oZsZxiN5jwRgcBrPVXJZbxUwOOSONqnkuTC2IWtnn/7B
m1K8tM57upghpaY3qZ3L/koW1bB91m0IHYOPSgRlgf90J7W8A6EuqjRUwKJEE3Ad
7MxcVkUwG/hPE5Jfp3foEKSkyS6VAvgpvbe8Z3Q0WeF3mNltenMXGZJaV3SRW1Lr
xl9Ymj1GGV9xjKw0mn0W/1MaEcVECpzoxiUekcNA9L+sLHdkDiW9IXqTR4ywcov+
zzif7E8PwWjIvXZ/QB030RpRP/rBsgr7Ba8ngpoWUQDcJwBI1dPPB0tvTcPw64dx
ppjdUmgnvP8irnwYG7jwjRz/vGtBk4ZX0qN1bfaOcw+7xXdjQld3dCNLMan6sJaL
pGVkC8kU0pGLNmsqlVgxFoAf4YK7UuVY5q+TBmnrhb+8XcP719754zPQiXfX9T8R
Na6GzELEficMbTBHz4ykMdB+MXTHIIJYxwEP9VzhkWkbeSCrz+OKO5OHqnfUO0ws
gDuEycOwGtAuuL7QUKdO3kH0YSnLQa+6iO2Uf0vKlz8LjdmUg1nsC0NAJCySikDq
EIGHwWSA9Oxi7+Q+MBLQJBtg6R5srleoHsQh1SPJhgF0ihnGodlPrCq+hgAiDIXz
gSYth291ZHHU6biE/AZefKavbqBAh+i/PKpdhrfS+Iimi3P9qziaNjZsseugP9YW
xCPLg2UWl3yEQj7ukB0vJ0ir1rLxk7qqJWN86iUBdDGugiHTqz1vPfwR7Ev36j2J
iNIDEKEx7Nq+Sv079ZRBW4OqQLIdkvW+ZCHy0/xSw3mC7Y1O0qCMemg/o7q2EYic
/c5fIhiWQlORhDNDUFsjuyKXRaMUkqeiTXwarKlLFd7LcdGTnl8IEODeTBZfZk6O
2AyPqzQbLSGyD2EJqUJyZhQwoAzj1+BABwws3gX6sW5mmCpRopD17hU7v+c36zMm
9jWByWfK1x9LrPfJLX3kBNTlCed4VVu9713pkJKmIv4odi5h55KbW0PbcUMYt4M7
X4gPmmEKD775ih6IZqy2T58KhOJGkojDDGbOHIiJJo1CL/SUPAKhMJ4LCzcsezMu
7A/Q01JiHKMXtRdP56ReCVyXOKSv9wUsud5UvDEFIz2qWtFQLLl6p+h+5hQE8hK1
hfuvet7mddYiYhBd6JrXyaNVJ8KlZ7AevNXNV4ohpKNrE3yqJ/AqNFefMn1j0ADo
OiN5HIKjnMmuxj+g3MeO35kxHsgVO9UzYdUkqNnQAvaQEaPJYmc+8THXahJSv6AS
qbx2wI2qLBBRUxt2sHv2SUw8vcl/qeoaIgTeo/RXKAdd8LvIkj3l++bdKW8/QS+l
fcICHo7hYwVxR3ydqDzrwfySeiYu6s/bAaLNfzvBEQaiZZYsyrS7BvlKoqRz7aQJ
Hr60umZfqHPbztMZ1DmtKTUUzfU1vgPgOYZxQ31Sa1vQ4YQ9Y/eOsbVbrJ8cdM1h
FvVnM6AOMfoqTvfHmSrzq9IJ5O2qs9yrFVcLXZQKuLAPRwJQ/YDK2rAkBcMDhGCM
UXMIUlZHmARNznXsxzLvhTujW1HON8X6QmEUQwLG9r9nCL22G3dLAeZOC+Cv7tgI
ctRtc8osLIqhryekCmaN95Do9HmJY8GUpzTaApCPCoNS0E8Dalm3KjAS6fM9l134
zBILOpamgNX1kE9Zjcdh5HKU2a8cYbWQFDHsf0HbDANF1cqsB/CdZAepUtYII/hE
43rjRqgPBIrbXUauwBmww6rOSO4hL/arWseBOK6jMq8Nm3b8qitLdr0O+jEv2ioR
CDG7wN0v+Zy+OJHiI/sP7Ccxzf/NQe4SqnpyoxAsbMcRSpcpblVHOEVSK7yQKRZy
UkJV5k2kkn0DxffzG8Z2ScQOfjsi7dI0vCWM48FpzamBBNPPHju1MBiwlbY9Y0V/
gEsrLQkXwCWb3MHIprL7SbfxrgEkUHaLuLXVHAZgVdUMYeBWPNytNahxslSCd7Ft
WW7gogzJwNSN/v3oI5fHjFYwYiKuTUXjThd1ZDkbR/dLfxwzErDSmqnHbWUvipJP
eEd3C5mERb+0aC0E0lPc32jg2UE9mBSNNVKudbYce4Zq03a6BuFxj+qVO+ngvn9z
Aiaf5llIacMDZ641ZmDvNhHSwgr3+4fF7Q46sJFj4RycQdwYRurT7bH3fYCgT0gH
9cJBLR3tp16rLXJlWuUCFMp3Og8MaB0tuVKgPzTAugbdFDl60QkGyYEVKSgqo0R0
MU3MyIcLI97QF6vS91Ol6HDnK3c3q/XUEh4R5gfgZneqDA/dQADR/w8EG2byYJ/f
54/8tWnIIfq2cyd7KQ2mg8UWWrdeAuQqYvL6iFRenbxlBvxuPMzb0Lkr/B/NBi7F
FzmR65jdENsWzmKUXhfiW3dLZ+qQa5ST/j9WmMyksi+0GfuJR0hUWEe1ZON5mQJK
6Cx0UHH5PCALNYS/smm+e2ZKzbeor0gbUnYWZmuxFYWiUw60dhNt5napAg1C+dF5
1UT38AGwfnIVXP6nl2rLsADSb8+5naeTVldKm+6+x/rpzKrf6URWzoqxKqgDKKCK
CKVLF6lg/pTlUG+F/wI/O8DDHoS/FBtq6YlQCyX/nqYsmsN/bqpO9stHnmwGYSl5
EqPDCx6emt3U6kQWdVGrklD82UtxQoX1EFYZHdMLi1/iQ+/lOzMFvOeGiWqPfiDC
eS8OKW0ZB+p2skFyaZeDYisq1NO9Fov0pYYomuBvXocdwav82jPghMY4QwAYGd/2
/5a50r8t6WWSJ6ZhPir161d50Y8J7gul+otTm86PoCKTpn+CXs4gWak3XyGY9H0Z
5TCy5xUSFeWjAAowxVi6R4liQ0DdyyV6hydrU4AJNAnb9P+badBXILwpChJBYgU9
3lrC0OyvZ+4qOymNGPapV9xKqFbkdAGmSoJZx4t5Wzb71SuHZs1SYUmfmJGb+9QM
mmDCw7B2rg02Y3v7i5WhEBWXAAMsPSWVLo1CltzyZ4eT2h1SiBeNtBzmtIZV6xKT
LtmIH2yoO55m1I/UrqjUcLqTPGv9BnYDMwN18lusrLIzKTkomdvqhQTwVHJVCskJ
0sWY2O1ymMroY+DbqPhP1iCei2va6LWNL3w/uJHRRLnq1lNpPGOW6+9gAsT3Yrfq
mNYTVmdvDW/25rGTeJ+VeqkS8AlV70dKixAB/SuhIGx2hSIXJW9nq6e/oWlb3EhO
byFMYxg1nV++dytrFueejLt2SHQa1EieNMx8gNDXlaF64JSQLOkI7JS8t1CloaVv
DPvE5zUWZmbZL9nvqJCpJ9M0ecqX91zTAHtk+LE0kEq8TnlqXdgojkgU/mZHN1BU
cx+QJ759UDMfqS9y+H9LgY+Pe2SPBcPBnbAOYAsZ7Oxb5ItpyxwF+TjrO2iUK9S9
qpZh1m3WrIFS9SiLJURk5E+hh7MfUhoMtqamZc9EiPg8pNIXa6xOqECZhUmnuRxI
Ce1rfHSDZK8+0ThiM6zMfTRuBmUEhoBKSzPMfX6VjFJdzDsQ0mOqM7/KH+4vHjp3
EQll4FAuWw14+yZYoRNh/Ee9usLjP09Z+XQ77pjQcq2BwGLP0MdQKkgpUlApWrHu
rhiCQqFSavdvcc0UdAhlb2BzPcHtI3OsrMAnCJilyGhfn1ZcfeyhPKx2NMTv0l9e
iqT9wxWh6YPLR3y4jK9EEGuEAD26HvDJ+pMGa8EhTuFpYNthNn5KFzJQ65Wptzl4
bZQeNcS1yqqX8OnBoWckaS3F7tYsgM+2A+YGEbb5uflC97PhZX4UrXOZ8HofMzNJ
CZoa9Pk+a6W/Dn3h4ifD+i47vOx1afintMuzoC+ApH7VUxZwFKd7vaqdamgzbwoo
R8+n2LWzErxJHlQJzXAk5qhAp54UtLTKnEI1vJCoQehSQWxz7u3f8ZxpWdUSCctO
n5aa5kb7gD22KSb+DLQI/cy5dXvz8Cv1ZuZHIY7iVgvW9kA+peuOPEBKO3VUJ53o
3ukdZpnvp2DuYui/0mogaikKukBCMkGK0ETrhxW2cG/0XsdygjzBrozWJHRtyyCk
lJ/waeCRB3baS/ptTOvhXA8QLmpwG1560tJbRoOdTSevtEbvPcCULDk2exouqszi
r3XODPCpTaA9GiKYpYu2vFUSdtwaXBUCb/nBqst2vUTAT7CMvp4lVEQXoJcu//r4
zneOhPVMEQ43dDzR3sIkcdhAwyE6SZ4I5arX/ByySMFm2knr4hP3l2Myqxny1WF/
L07Qkp7c6vr3eJC+nvb1hkjQwi2GBDnmDiCIexpUWYrzO6CNeCoM1nFjkc0E/hob
DePbMtRcaTH8yZVljA2kyPkFukyU5nQGTDLJt3KKmFef7NoYoGKL6wZbWwU5dWVp
na7ATLYJIkECL2BFEBmOm1yQc2AX7+FCUTOiSoqKCbwATtCzBYUNm8+R7ay/mlvO
TD+tKaG3o+UPTnSsiatmh/RWPhH9Rwu/PsQa+YncXsnWphjTzrxIfm8Ur0DIBYgC
4mMayBtxVcz6TZs3rL1OdZ0wNBo0GaWQLBhLfemZnsay+vhLfnWC5cVcjmmISrT/
Vd8Fp5ZC4lpXB293NlJoVWAmbxye5ogTQ9rED4OxkwQVZm9OJLJdxQErgVhrBppn
e4gR9pnzKSyFqG5PuPiWwVinPyV3vmDQ0g2pmDwQEJq3Scfm53L8BnZXlJaiKxn3
Wa7AhPwdylAxA6lqEcaL/gGIb11q+3tsihQES0boKGrlB0/0D0i2kPmnSQpVu7eB
mgsPhTtoNPy/f/kgDn21oX3h0q4kvzGC6B43agN3NPLug8jBp2HUi3wc3mkzlynf
LInm/qwplM9LLEy+3+/LDtRSp3r/5yHmcdUAhJhXa/O8aaodM0oaAb+37/m6lQhk
OzIk6u2h4aFOsDi6wBal+8DBAlp1UXPlnW6GMT1aBhHfj6CQ79pme/JqhwdjtfSD
aPCaCbfTkYoOQOy6XdMMmqgONmW9th8lkp6vazXId1tipijFAcN7liUTePDSLlue
P2Ux1ui6n0QXmOd2T5zOlme1aaJhU4+ksaU2RbzHWPl/AQ2N0AOqxAlZS3jTmeCD
pX57Hc9AZCKEIX7RHUdo9yDnqN98toxfM1aislbNDRcMgGcBj4ZuviM3Pl/6nTC/
VqwSMO/3hmRBGlKuKl0bQHYmZLiqLyPOP1xGrtTPdOYtnCfIkRP5C0OVRtuiUXgw
RnIeNg2w3H2bOcYi7L4ZrpNLTJ8CAzIzoAM4wiW2Baslmemyqaq87AlY2uFkfMEq
gky2LH7qxt/7dk5ieg4wPCjtsrBerdOq7grBj7hBVxSJoAURpga3hDWDoru6LMTP
IbBwO3W9hrmsAjY4VERu4lXAQAwAZZRbEYRa3OnCGfOHORe9CTwtGOhCKfSLDqoF
yKI/+/pjlXBAojJ9eREQI1LIin0Nz9aRRliwKN1bX5j77X+MdXhFb76x1OTWljUQ
PKqP5H0AMnOO5RyzppNpRs2zv9zXqjnTMlx1Z8XOlfJT2/h7A+mzmVOEgj+5/C1/
ONdx8GbyBD/w8j4XxpVOc7yVO/mCRIdGE1cvielwrYtltqKYXVA5NenKdduoBNSN
k89uCVKVoojO2mcuVILCEJae48g28uffYVlNU04uzg3yFSzM0iy6Xo9Iy3uN9PS0
nkjnPc/mxmSRjjNTbYtH6JlVUpwNDmdaW4SUruTxqToN4aUEse0ublFfuNjr/B/O
pzMtuncCoVQJzVnP+cHsCYSnbuVzbgep9jhtq6qlVudGBfclQMlKczj8UD5gzVen
VulnP8pwXYVgPKRR4nBir3wnxrHr7ba1Wsyh8XZ/ccuvAdj3yaoCvhiNAZgGk+lW
E9F7nmXN0qHiEfIz02GLF88e77GNJFTntyGiwiydLz9Iv0oqJrVleQ4tSm6yO4vg
ni1d4ODbaUjYjVN3IVLCuwukmB4GZ0DC/KNwI0GWGePG2/yWdpOORRXJvxZ2hm9T
SUR4cSKBRWAV2/scjPRJWYP3cKEkQ4MV2XtEyAvQOD7d67c+b0o8VOIZY9kK+t4c
57xctXgkWXGXYHmUHm+ZieBsk5wSWAh7N03JMHRb5m2CCcXlCUEHTQVZFObjX/nz
GApWgXvWlSUDrhveiKCO024yAPJq41+CORqLFIgpJ4Uxyhccfi2O/xTrWcGRpVB3
4hQqrbxyjHd67lTy/fj/fh0RJEO67he6+j3e30H1ostUEO26/PfJN+RVcuZuUTl2
h27AL8KjvblChp89YOaa8TPVZQtlMt34Zv8iXTTqK4edPucRR36Z6RzxES+le7dg
Txqa4ciQH0WU+Tp/yqK8wRTPGxeQup6mhWsqD3QA98vocyqPtX6l62WATY04Ec7c
JLhL4+zi8aIXhSuKerLyoL4tob1fvBqntQjANSFHLj/gz6XaYFYESyVfW0u+nynM
XRkHwJl/a+DYoS1kJcLr8qA8iIyx1A0J74SWS5u/78iRQvKbwGGh5LNV9vgaRiHH
AQJX8PwvLl0J6sgvuzr93kW44NXQPRbllFZUvwYtZftVA0n3IxtrmbPWYMecJ0YO
/hL3cvqK9MD00fML1QolUatkryPRFm4rJc1t0R5oLrh6XjKJ3/mUmnsgNqrrH6lr
/iilmTvygeRGWTqoefxW9YWkrNXzNt5tIM8+AMVIBkwf+RiZ6c9a8o7up87j/ZnJ
FZ6mSKJYtOPGgQmba09BEQfPU3PLi5oWa6JqvPigvoxJLQ5Vr7pRUzjQDG1F8rIo
fM5ry5FTqX345OzI2Tw9ispuglbxmV6FRdnIZOZWFXqGy79In/OhLj3G0gxexq93
I2H2b0+ISzcDGhL/CySAeZRxnyUpx/ErQlHe3HowTwA44GXLKBisgV5uMeR5al2x
jxpO+flUFfHZPNs4rgEs2H/qph2biazeuqtGc3sR/gru8wiYNb0E8p3dl/T50YfG
YR1F4fX5t/oCggWRZnFJO5tY8ahNYyL1sF5ErLlkoc/n6q5/CHjbt/ZHWd1A39oc
oiRLKLbbKbnpw7j4u8j2a3wCFaGCt0WwlKJMVUWQSE9hq3xzE3FbZaYfVE6TlY2F
EUFeutuuEb8Zsz3ehn6cbCZ2hpiSeZlqDtFOrdRqxwLPACWLDo44jWQY13rWZlFl
+rWl8Ro8dOO4Kb0pBkVgC/Ok330c4syQ2VD5CvwKa8PAcbF6SqdTcaJhMyOR+SX8
h366rWnfiPzHWngCKzEHaURguLuJ4EpOZbDXu5u11A8ZD2aaqudq77hSP7yRrSGB
wufTKVYeFxj3DVEJA8jEMGPnYoEb6biM3QIMy5c13wuOflH0EuSNGCCv7PJnraBi
ynBXeRs4MbsTYmVQMXkDpXW0XimpV/3mZj0f7xraSZmI5ztm4f/Lhe1oSQRY/IV1
XLEGV5wLy47bLf8p1oCWf8o+JPdN51tIC6OiTjMQlzAofofC9d/4xosupvMTNuK2
LHZn9g/Nzkg9nheiU5tuAt1G/cVEBbygzp1GdcAIO0ATK6t9Fh0a3sEYkxr9t9XR
P1d1qsrPeb/Xz8UlDMkd8NVGASbCF6thiCPZ7XqbBXOgJJhlPA0QPQp4sjQQdxbz
hRR4YYSgAxytXltuCgbo5sEUzngZ65EqM6zwdxhRLjgoIIlmthbc3PUM3c5nfAOf
Wvo8tTFgHj60nznqIAk9qUrTHuRYhXvADRuj83p6+CW8h6Xrokfp7TAO2CWkVmEn
DV8JhdnV5cVkEZKiS6J2VAH5Bcr+3eVrtN3Mykkp8+3BZHZec+nqgpL1LVUCzQZl
ULy/CFhAaZdeXoYLwn98AxsTi5aCRm3f75VaEeAh5pP4V5AMYKxvnkR6esTm7vx6
i3rhIPlxTmk6UQbIebnApHn52tN6XdlgtpCJUeIQmvPakeLPIEIqszCI83pm789u
UVmvODeHKnlJO+sjTJ8TkgddpY9jP3CIwo9p+C4UAyMCZ9sJLm6YTi8PX1FHqHtL
/bNWWJXrFhMk4wwWtwde3ObP0PwOpLO/qfSJ+x1pYkYqVeBKmWGj20cWYn4MBlC9
yutkrR9Tn89YEfBONhAt75XG5HP2tyW/FuDPXsRfyZSipctpO4MZg5f/KoEYhdFd
6CzupPLiuAfFe3W68mpBHVnmQS8jSNnZ3D2wTkBCCFzPsAhbdHbqU70M79mpFrNG
cW6ROZu7EMhTbSO8DDPAXsmXHN6rABwyrL0oEr47tuE5McYZdN1OoCUCV6GiJAGH
pYglS9yS7+uPKZZ7AfptxhwbuzvTE9QwZ0UxGLBJG/qXFo80Ex0TcphSxFdaDdxj
oBn5YeXAFxnVDQryey4AXzJm0P3s8iILJ74dhyrBPoqdYN+9XvaR1Qvi21m0Ibxo
7u404wRWqYrRmkAmFX5GI9LYbJrsZfIzIPGxalQaaFIRPa+aYf9bC4ZiOT8CkNiQ
az+Ox7TJIuPEK56o0Pi9KtEZ7SR4ot25bpZXqYRkxxQ7ysJ+gc4dMIKbDIAEpbCU
IeG3aAGA2BTMrpYFKO7eUQ90RttM/ET2wBfmDLxQCJj5ggd+wHSvQq9EDcobc0Qz
LW1CqWiVMRi8qudU9rP6T8b5y1BvSNM882Lkf+65rG1bnHIqXrhbr2/Du2lyEZjD
yMpAGGUX4TIXpnE0GTlZvPO+tnZt9s6WUGpyFXe/uGd7Q2SVzTOMnn+qeNu0sSPG
5eppzTJZwptWlzqSoaZPwZyr3y75ezBHYHBKnok7C2uFVQut5As+nStFIPKPYr71
sg6F/4gzK6x7YigFExAMlRYsrGwupy01udLgPakeXEKfH/pMF5TbGz32SR3S5gHM
D8ig711e2EfZm+ekA40Cn71c2DIkm9obNhZHHAW8uVWW14FyKGExNFqecIQhWnxF
4gmSdAyISwPgAqgyDEe5U+MMwVjUe5nV44OamzxniZH3rAyQQPT8U4TtZ8kC/0OU
xQL1yy4F0sfpLHtYDhHDdTthWaslLNdIb3/BJssW/JAZKMrCFaNjyjl5s71gN5EB
sUWTcwmR+5njNE8WAlJatRbqe6bNe+TURhzo7llZ+2dEFzt4yDtxTYMdE73bawVj
yWER7t8W/C/8hPhxhqB0+ajDHvVsm6jIkl+xl15jxAc3H51rN6W8JA+KHaHIBUSU
JHvTX/Mf74D1DDKo8ksAmOVYJHs+LZ8U5J8MkbIEImYN0O4NvZdJwgZFNPDFJpo1
vXvthRQ+RSADU2sdMO1e5xI6Cc+slzlLRm15Ja/8Omrk9Xd90nqGDocCd0v8Ucaq
HtsQAnv7bDzB5Nbq6Dn3JA4v2W7f0nf47IHgTTM2ibFsA01lcLc15FC6iVLkQ0gY
S/XmqdE+agrqblfbKzaWv0fVnRmuwwo+FD3YVnAfzVll8VfflpcqdW797/xLL8WN
PgUkXMSjjcxIBg4F0LBEOk5i5I0hkaPhwrc1S8qKXN4ibAFVK6f/psZBvLC4dQZ8
Nw3gYkP53ZeWvh55ssm7yq4PzVN6qge7QZBY8veybbqoKYPAb/lkzRnefkG8BvHX
JATfUmMHtoWB0Y/NTlSlbGmQfZr8rHq+eTEzEgaWxiexgkpl5c6mbzRRaoLDKjf2
xXnyccCaPqJWKtbrpssY9IhmNeOwykzGLTZxSCZmGZ1clrN7M0Rq9HnmxzJGITzY
ynuuyQ4YSaktMbGsXlULqH8f/CJAxgvibOh+EcNn+0tX3KGt67UkwreceJW/UD3A
8ZlYAAUa4wVJaS6Xu4a9HWXdX9B0Z6ticVtI4c02k7NdWTAyz88ryw0OzWIpyBxm
4quejr6L6FY4V9bZML9oY20yhrV8KHy3G/XhdUMoytAhtdPJeNqAvwbeFfE6ypI6
GbakbS/T5nfPJYqArVH8QJfvH8m+k77FSf7Zyx18rxkIWSpdyhvohTG9ggMODqp2
Hy33MfU+O7JzsNz4ymedOYKqM7KV64GNv8XVjUUccnK+n+PKi+Rtx1tVfCGOhs5E
nrRrHjtcSqsW7a5rzci8JPtwk9Qd/LG+DnGri1ICeQizdpp9zp4yjGyDBjZsO/NL
L4LcEW/PmLX5qB/yXW8boqcbsxqeXMFQMEGzMaLM8hhG/agUWD0Z74zZeKL/cTia
SXvtvqak2e6h7E69BwhMDH16+pA5/5pjPg836SfayHvTIlnwRz0GsQzqX+8ihDb5
SCZuMLPWAlzUcMspirUTqlCerBDzQcX/Ck8+eMKA8dfPiuyapedh+2YER9S0h1t6
iPQyrb+gfjTDsa8kpGhrk5yyTAKDqymJlJknz3iOc5XsYHWQzTLRS1yKIDg3FwYu
c7PBQXv3a0Q4tNkWzx3cRD798lPsst7DuAT0u0MaIGORr3NAkYJ1/EsKCBQLQOqJ
zAVQr2W6x7ZsgikdeABUi73ctLek+LsLUsLukctcMfqRaGca8uxcjpUdJHYCI4YO
w0G30Mv7bM0I0tmvonC1JA/pwLswC3F+Bxd1Im4eylSlC2iW0g9NFBOlnQeDgU3x
MByvlTQ89JgjUbz1MzzzUpzPA3MkVurZ94PTuH7lZ+UtTmj2KPJwjyuXsEJbVc/r
AjFW4QF+/pARQ7zPfG5ZMuz4ioAtftA5LbXKnl6tFQTKCAgmCzYwYW9/FUcO3XiO
DRSRGk68bxQSOK26rphKLve3Rrmws4mwcXIm6MrZDAtKZ9uoZsFPSwbJucvfVocZ
X/l+MzkySmmXgjoYmvJKrlpfEVhur+jCHPYBTfE5srznUBCbJjdJZbJIWameAnAs
WJdLKKwGXN5CKYJZqgd5bC9iUzKEkzhwM8FelHnE2wiRCYO1AtHjwscvptv+Iy+m
rCXFVm4caB0K7lDlVZ+zasPZ8p3NDaE+o5ItkzRCAWAMReUzfBTGqZBUFskIpwIm
Kt17xoiJLjvNt8LkKpR2qIRn+r6lTBbfL+0EgHyOYeQei2C5Jt1r6wfxdJ+erom3
J2at6AO28DF5w0/UNs8LUq4+utZ1SVWeX7gFptHcJuzRAS2TtZN3942R80mIqH/2
GQvle5zeooL+Kg/yiwMB/U9FvHYWIW6iilGqXax90r8OnSyydrfD3pguEmFuim5D
X1YhOWTD+At0ifYMOlAGCfcITBRWvBxPMuvlNbu1NeU=
`protect END_PROTECTED
