`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sBtidsiy9Gxnb3JqklkcKWZXTD4H4cg78Vyno+Vzf/KCOdZO8EPzFgqyuXBacakb
sfZl7dbLaNQ2iPR02ZT4eLmqcOMTChDwtMEd0Y0rfcT0kxICshtHgsloZnbctPAs
0ANGodvU6mc4vAmRAud4bZsxuhznFlt5Hbxaykd0ZOy46oMtbjGDnwu/rUi1+yYo
jIBjfN/Buz2T+qtntgb83FOvjCvygfiBvYnW2LSTOex1VlqaG4Palx6ytqFRtppO
2fE46XaHtZf1Zj+xZfTUB+oHNcmEIH2Ct+dDlxWSW4n5WXSZz6/QNhW+GXbox/qE
g5uFVLFj8pCsc42EJkyONZ7K2Vke5dohqG14enJZ6rnwwkkzy3McLbaCcdbASSyD
m0jXoRfvcsXTANA9E7WqrGVcNbpGKc9Msp2nB1H5Iu6UU/GC3IP7sFZwhQxXuAKb
iUsIkr8KcRLiFnRKzvK/rzU80D4CtG/lY2PEKeWFIrtwMeLZQLjR1n2UmjqlJIw0
jOeRVay1tl5BMXu+p1uk95LFzlmNcypmCSIAXfTspulj9OuayC891zLr4t+l0Po8
yJ07w6SD8LEdtzvbYZqIuAUDyJD3iUzXCumNnNVxZnP5HAjhDsMSGL+FniD6X4Js
DUOg/YRPoWCGGQ8T3lceh92uXG7/mW7wnMTyyyCOHyxlzx0xatR4vfSXLAXQTrHN
ZDHDqJrSPuDLGZ+pr63mT1NvL6MwpHP6t8Xp+zJu7GwMR4o6m8hgtv/2pRD0s19p
vukeJVnrkcK3szk2064Bxg5CXP8VwR+QZp896IzFEF+zyumTblFi8dzMileGaA0n
h/d9k24ldWV087yH5ACUPihGAVwnEOMvd3nFeVjHh9GPFvvlqt3OG6nUBi4kfar5
K78U0aU737lOm+ieu+H58xdUrYrQYBIOTpc+8tWd4eMzWgeR7r9EHDKVR5ZQlD+t
g3omPu9m3tVU+DyV7jE7na5VIlrIRjuY5qMnl/e+jTbQGer9nqnubcF0XaLActhd
PDrhkw+QPXHtR8/uUJ/+DwTRzjTJUOy6Z9arTxZqrNOrb4rjk13umzWMdqBcE9WV
68jPh7XZ47wjpcUyGDDHV6PBzStPsqm6MxK4fuScIp63HNz7GFr2LI27dJcxsB5W
vKe1CjyucUTQPex+ZbHULCchVzbfK02ULPVP96O7jVqJiJNSdvbCIO0NJH/RX0/o
psBIaqguHAXUtci4acX1UhfI8430BlckP117OrRoiGu4zXwU1niPwIWhDnVUfnth
WQ71xdmCQHP8id6Ua2SfeS7+pPRXqIRyOIQACrT0dhMKCA2tx9hWzoCWagF+0jqD
uA4FwZM8dHFVKc71Slz/ZlqRcgkDqZfNS2311qNjfrMcezzX/etAPFttHxq6ibuB
Z0kDDUImGIp+YIWaV3zpQmYi6ReyTTsXMjMlWSTcdJOYsAtNikURI/9UxhQKSXlJ
YUQYUHl6qvmHmbUoQannbH83M9VZw//VnWfEeTE1wHTsEkT+jQ4zjRXhXDd8c1uw
mbMDNF7wsuPJgM0UwcmArdxMwFPe6f+qhRwhCtf5bXJklmUoK0POLvKy6SQbhBWM
HMnLHE2fGBK9QNy+Pe9KMPYLTDiIqGKN7V88te9R4j052hx6Pyz47ziFywa41yt+
E9WWtO3zquDv/Nnpn13Sp3UbVsremN/s46TJnNmG6ZJRSCqwT8rjelB6YB7PmiGj
IwjLmKfI0N8kOkKnn5kfgPLAHIMwiViagV2Ik59th17LKdkH0W7qcNbShlCksMLd
rJLgLit2j/BQTLZTJGoAQ+O3ayOQQ6awFsPiPrL6/bIbuAityIWjXj70Du1r+JoL
geprhqHmAMqxsKgoQ/WWKaM2ZoiYJl9glDM5m8kxsRnTcTkVXPIqmGu7Pba5Tl2R
+40ALjgd5Z9Z3t569z3+cPdwOdEwxLcoAgW6qVeR7RwUcJuV5OWnoCZyPuG2vP49
nZ+EZHCHG62EIsybCibc8M0ApPy/VZCpqPzWWphIAG9Vso6jFRQsLmMilARK66mW
7qRRMnHPyslCqeVQ573KQSyjyl/J2iil22PEiVHNFTc6+cmEYtEw1NBCkmouXv2g
vOfh5V7+BopnCJiy9mzxSvDLqsFbQOJfGHhWz+y344Ztsq4r27FpPARBK7szZeos
Ffh8WR8a5uuBFO14wWaK66+1MQVkyPwHqUS5zwEoNsPZvnvVZge7jVURKqnx2MUL
3og1gQjggukqbCmEh5eVZeF/Q51pWQmL5YjoNQo0nQv9FZVjGpUZbc5/k7x1t32D
xXuHGVwXV1vWGj69BhoRLKKBdNpW2jFnAgjtpQ7xoXWxERamZD8hXpNyiOjAUoTD
Po2hSSx92nyMI7Vjrri9Z8fAUhZFd8iG3AYF6k6+FKRhtWAO/GmWigpdprvc3/0j
I9JWOd3u7ATAm6bv7DtBKDjVPUFkDqW9T9SMXO1w3Qb2aOLgssxfdREmn+iSxnQt
3BHPwUP8w1nlWd1JoFtPLA==
`protect END_PROTECTED
