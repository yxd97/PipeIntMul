`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B/c1cAxo5SY7kBwbuQDn8JnRyfkxoSSAxXLK+3ZeUYwFEG7FSBGooU9QIqisz/yK
e3D0Ha6MkJnYpQdS0TtcVjn0dzb5I3yscCxTVrtT3AV7eGFbMiWkwFSXV3fi1kQF
yT7WLlw88ZH9EfXlxxYyPS13O8ROTSoIY9HDQSI3Xnigy1obL66vBr6sRQPB4t2t
jHQ4ze1kp7OVjpF1bHh/d/g7DcnOYL+Ovgtq0RriVfdNA5gySzQr93aIChuVwuN1
ALSzAm4vYI93DZzQANroYooF6hWVyoV7ctNZmmd1WGo/WvYyUhpT+HxNt7uA8gP0
zvpdh17Z55Ockw5vpRMXbq5KnKDMfujx/sEX4N8VnAEk0bNBe41jbKKmdiNwSTSn
gez5XKnLBu11RcJzpTgsiEcwILlrhRBkHYhGLAlEa078IG7pCLYhtXG5nMOxjaGE
gaBktMZs8FsAv7Qm767ap7Hznwk471EvHe++Pll9F5mWdOX0RuY8DmeNUKQ5n7Ss
JiicnEnlYstj7Y+xv4dr9TzFEYPy05WFyj5DEc4/waKuMiq+TvUu4iMoxuznpz44
axFY/lxEA1zR6686uXVyjdU5oVmQUaP2kFMRHoh7iz3eBewuM9eXFFVE4tIxEK3b
DWkWKpMOJkFTMVADDtcLd5fh/UcHUE3F/57bIU5XzgeaUCZM7Bwj+dDch6x0Iz09
0FiP4y9wGz8rrMncvJd2Z51ZIX9csWvYQSn6JnueQ2OwIxygYqhAUqkf9+eOppMT
vvCvdnS8/ptXJVx+4FiwuyZTVpJZ7rqX4XWY3OM5K90qqY88CIU/ymoBkxUBEXmn
s5KBzFzbtII0uWT3Viig/yuWIp2rDEdjYwRiBcAVyyY1WL9k0yMyzo2XIiZDpxBA
`protect END_PROTECTED
