`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbbRqBHzkrAYJizNuCuuAY+Jux5YoE3SsDIplPcQMMwjoeKrVmwrfrJEf+CNM9Sp
9IHYb7ApY5PspV5YkkP2dKH2puNyhSRt5ZLHxmFn0GynrCL0dnSKmJHHB+uYM6+x
YK9WGQ9MCtcz8oILUf9aedqx7QE1oyM2y/vQVZoSSzcQpGhh9jGOHZAB/FYzoMqJ
qegO0qV+Ikzp5qx/SNUm04Q1+h/dKVraEmJZr3tA2FfoRBtDwciNE43v5Dgc4b64
4VikFBBt7JzN2bj2/19XunDMejVuXEjJTnOb0/42CvDjOBdWCNqbw6x60MwBZM+M
dVXLg12Jv8+MAdaBoxzDemPCCMCRLAJIiMTCNqGV+nn0aJRM8vXQVsh+D6vk5jLg
`protect END_PROTECTED
