`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1AW/4oD2jjcDlp2M9Lva3pHwvWBlRh0bWsvOgsn7zMi68fu7Z3cGxPEnf6APDpCq
vKJUH7oJx+YbANZzbgg8r2wO+TIyPnsUJNqLC2Ttgs4MFVN4/+0AuQWFbNpBVYu3
vOhGPuL04pKiOTxtnrAkrXaihhEJcfwxZzeKkHvTVVB20mELb8oNS8xBgX8Ug+dk
6wgVZprQIQOewVcKE7uAV/P1M01KN2LvYvOBPNRHCtMRplIaxXAIk6LO3xaGB1SE
+hfY7/Irru7cukWR/1DGGmRLGAov27PLsdKTWaEWq8w+EdM5vNZmI+yDoBgjJfCN
RfDFQH8SmffWvW9qNnPV4ltHXR6JSoENTaNBgi3gcWM8yPich/JtREuSdN/KICy1
rbe41gIiB06C4KB5DHWnQN4hhonNTrZN1cjQYWyNDFVvk9GFbRt5mAHmGtUHqpwR
WnFaJgFKcn12nwcOu2fPqFFYHg6eDkKqt4WRqX5FdWUiwGQLRNEyolAbX+fpX0Nl
L5KiXKCqKBNAXjDxb2Fj6QvVolcw/DjpurogWs11PSrr+2/08Jbxoc9ALVBpqers
/ZrSavL6MdWdfuTL04uTDrBbTh3lwrfDrCW4pM4JOkb2zUwZmDqMz+7nUFJuu4+O
0GEuhv0BRLkJ0thVet/0zb6mRvMxTRv16K23DqtqOiQt8kcRk0Fxh0a0VCLOIOJm
yroZtYKKAXgaZ6l+DynT3V+4MSVbYwFMoNPwJjzmHc/welUWP4zZGh0I1xyeZKPP
ArK4UwSJrz98c5ZhqN1xxcAZHfcT7bSh4HmgDJzsbdeOQI82EojVPNjQNayrfjCP
2ol+V6nGbGHbDQohMhpOsObj4o9veXhDOdx4e0qFxhzm+BT1nd7sJFZfsX2JdBMX
iIQqK/4jsnNA3cB1E2NoU8HotSjyyu1zBkEGw8FLh+Npjoap1Xu38evbaCTIg7J3
sr5bhV2ExEL/W79s3fpeqf4P3t5DG0OsmVzJtizXjthA78L9EutY2MC/nLIJoYza
3p/74dC83JsulW4p/rCzNs57dy+6N0y6xooVNpOI2vDWvQt00NM8f9wGjK2yiotD
Nv6Oi19qxDfIxKSSDlXdRw==
`protect END_PROTECTED
