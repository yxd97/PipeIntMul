`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pv7gHBwjSMlU8YEfQPTEGuYEFaIFHJ+s9KQDPYm2oM07RSF7QRkpFZybe72pE2dn
2YV6/1Sil3wCMMV842KuG9J08uyO3qz5zPus2OUGqb6NYj8jCGjInyp9LiJKLCVK
n+cUTEtCJH4NN0lcybX5esuz4pFjAQyeHu3g3xxJYW5cEBxDMpBy6CM63ipmJyHt
ILXpOwC7EbcMYG9PYZ+iBJKZMmNnifBR5+BfftgplbReutt43ow2yNvQzZ/zvlDE
iZuyJ0CnSQICCvTfU6QCfK7K52XTYZk2xqNoyl9tJmIcvjCEKCH2yamMS+UkI6EC
lBV3B2MGeJXlABFmNdhCxL49c6kIC9baAz0a5vc/OJRwr6DSxPO8g84/QR92MllB
yMOoqNhgkrq8n1EMPWJmLmS4yUvOu4uZB50IpijTe600M/mo0ofVstUYuquadXmX
s+3D1EB6RaM7A7ntz2cdwxcVzzcnO2RdSsPTaD/KBK8ySp00dQbwRWOamkMQXSwp
RJy6CqIXZFXXgjGhH5y+DVvz+la7H9aku9upZAJZTobMz9XBiVXI/g+3L2RVSXks
oyetMPt7UtKJprlCzkrqjY24GshZzJJKkXchz2+bsvfw0DxaPpJGIFwg2cLCI2cY
hjy2QJhHZRr/qMvHiZjRLdfREwa9ZMkINIHuwnFzUzPftYCc5AnX4GRcpptv2Y57
Mdq0t6Gd/zQ/qPHZXwuGy1P8PLcODdXGUm4WwQS8xM2TZO3OHWd1EcqT8m/mzNtw
5wGxTsRxYO2qNptTHaA95FYd0Q/8ZYxFRkEXOp3BJfp2pnrDp838fa5GwSozFEOg
LTNIhnBflf26E6RXfZOvQigbUF7Gy66Qk1KD3xQ6ElId9gyi6Aeph01zwy6+GfQq
072THnrMnF/bNp6eoiiIehvVwH7mp6e1y0qO7FOPJnoGcD6gee4tf8VcsQNbnKvK
vGCODSC/3Yz+LSYv+nB+w6NLXnhjddAFih2EVdHbvO/wdtIp+D0EkIT6qsrZqYzi
tMKFI/GO83PtbDvLp/fpUkway/uYA3pZpaWk2UN69aML4hEKaT71lhpRmygNuHkM
ou3KpbR6fnfAU3S8cgNQk+EArkI0iaU6+6RkSZS8xREmfM2Xm6VFLwbypt+kV47v
XYAhONFmA1aZdJbl7SEuZJeD0JuchnE9+q9pllBk/bGuACa31or859weJOAkXN6j
U/8r/sQl2LnuZPOPCSSC2g==
`protect END_PROTECTED
