`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4AeF/t33hoU6qg9SYEiYwvJieb0+JPUasQxRVzxF0V4pcbbQbNJGXlUGwwqbOyVA
36v33NUr+gumVC/NC/Be4KRcH95aOPXvTBtiAb32oT+TtegPP7B5b1CfwPCC9ETV
PsM/DNmAOO0sV7byqxMXMxKncvX0/aAykSW2HdnBmplLY1CTZziu24INsWzMMZ63
5g34sO1dRdNMYnN5RZu+JyzJ6VtSnaSivkYX44s6B9cAeKguKCLAJ0jPeWWOln/A
KICWfcYJwktkGo3a+cPpgiZuxD9wYRU7E9B0tUhWPfdYtnSTunwaPCX8EBjs8ltG
m6LK8/aE9azCuDCHu8xQv/cn074n8y6KE1SQFxqrZmWMHjvMphfOYXkb/8WPZmXK
+GLmq/kwX3E5qhC4/YjWnZc9RUqvsZq60IJQVDyDHSMIs2yoTmfVSAaazSW45NM4
izMCtRLmrJn/piTUHSMq5Z59T/hHyHDEVXfAziK9sMzNI+RbaaBU/9q5ZUpBG4XT
FB3CmPgUo9NWh759/sxFvAWNjieOLs7KpKWOUiOFimWbEi2I8wQyWFXE+VJy/Nif
m7HU1JylK9Ms+RICz3v41eQegHCXIwRxdLmSQzt7FQmyrZBlLiOi9kz4EpECQHpn
DTQ5+WbgAkidZlAdIyEemjIeZzsEn6yhCjEmXYR30pn1IUlhkB16shTw9X+aYZfN
E7sQ4m17RfaZyq0TXG1Fh3iaR3hJfAIkhzpaAsc12lsfNZOf4yvSj2tCcd7r3513
OyCpOHQS8Z9AKUoSFZI29Nj2JTa4He5dUM1fIYioSoTZ8yacLaFO8iy5+uQM/y3K
lp5Re6/nQPeBKRPXzOvm+3vWQMGwWpUWj49rA8fjwwZia+ncY2nmHpMHTw9+MGjN
oxs5F7ZU6XcNpDgaOn4Wzqbe6fA0nmcCqUO4jsPtOnJcBRHO4tYAvD9uSPB8EmUk
lN0xbVSY6gQl73UlTL52MXikiY2yWQW65yiTUKzZ4F0LV2uKNQLxgeHr2ZqeYxaF
45RNBrvB66UVmnmOqpTmXMdX9enHIFA2Q3c7v0W4LOBIlU8HJJltVH8M//RV/zu+
HLxwsHv5UnoAF7YbjW6WMcswc3PxWcJ3tH4KrQ6qjB1m5qfUik4JiZB60A5/9pUQ
`protect END_PROTECTED
