`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A1GDaAZXct+8wkGSuAxxOHHRdedxfkUPcrEW0NOb6xrSyiTUkE0byiuksweB4HXR
V4zPH0olhlopZToLdgKZTRa6dj+3AlYmG0JsStG2h9rY00q+3NvXCp1vv4kxkIKS
IsZLuCqW4H3WBmMHeqn6FIjP0retVOtnGXuGp0SXV3qhMpyUZqxTZ2E1jdNWi8ou
79D/Mi6w+gTG3Kep1gDHFtb+zmBbaZrDeA6vLCFyegyFg8uZl20gMxUomXqCUtqi
lI6kdikIUkMdEIQPs5kRLCF1qd9pt2Wj0JmzNXU9zau9Li9cp+c6pJJyJBvKvqNT
Z7iZjG5Imcq+Ph3r8lGQ4aycgTSfNokLOn1OQ3aB8SB9Qe1BlWU6tAMZMP3+07x7
V8fd3sKiTPmQ1e4p8rBDZLuMit7t4s+eKlEaiDXcqCgRvepqbt3L4en/2MlTvUoW
ewRz5K6phsEGentLM2Xnv9+mFBqU53VmXc98R+GpwmPQ7dD6zr1kHknsmkCpa64C
j3B2tapR+jcCjW+wBRZtR/KtAcki51Gcv/jk2IQWbyHENwsFqrabA5TMpahciGEh
cz/NM+6bnqyg5jkW9rbagiVW7NEfz73+7/M9nWTVgD/k9Zftofvf1IIm5vU91HkX
a4zgo8nioz3nlNQGYosV+d99SSZoJ2hAzTkqb2A1CAU8ewKd/pprSaQ1rsuL88hD
8v9MarsyJuml8DAffITiL13hls17EEtbkGmNOBha/GddyokDnD5aCzpxA877jsvw
oO0FJxE1fRyUIoyD2RIhu0ZDXxsnRRTRLd8QNBYh0nW+JXEqsqXQkzPjPm6uhguX
UoqVSezboTFWKbwJ7q4/QkDA+UegQBqslZu+rbe40uQ46qNavqhr5pcMnmdCxaQA
LT9/CvMgxyVVCyQs10ZTBSMyOGrVhvrq/5M+NR26B8ViKu3LNVtxY9kZPZoIXJfb
I2brwZvoE3wePq+3REdOqkF7vaWMzXBGT8IIWPk+CCXIUWGCbG4+wT5dTsXhJEpX
tkqmDylZ8qdegSUHSQIJbEfA47dOkEzZGX7eBaX2mCKO8Y18/5hrqQn1VBMgxBWy
pBRIgfMTwALI9/Svcikr+HFMG2Yhm9Ks60gw7o1ftkP5C3WsnD5sVFvJjM0RfxE3
n0FnGG+KnlB99DENCSpi/k3F+l/8dM9nAQgWkRGwwhLdpiPSBXCF43YJVHx9iQIB
Z3JcTJKKEAE8R5Z9OclToPYhQCZ83PYqnTCOvPUfeUg=
`protect END_PROTECTED
