`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
onLCI0NlyCbpiR2I5laAmni7+GaMqtImk/tePrPoDNhvd+vsljZqqzErSFFlUZZY
zoDSkEYEb5UQy39nZCY0sFdv6trSOY1CY2UIFz0AP6/7jMXu0gAzcXnWywJdoK2B
YoL2kI3Bj2aGbFb603UU/CwD9e7OI0nBMS79ayR7v3lGh1z9i/XpEH+XQ83W9elH
+mxV0RV3A3Y1jMq9htYVnXZXlMmyATq37+Xi1/t5ZwiughevwsuBTVWtqKj8L+w1
g8lFc+QXEUN3DTBrOl3cciuBwo2KEGEfX5fdquc8hlgQIlfxg4jLgRCqjrc8N3yz
IybduHsJF6VKIoqctRsRC+fBaaY29KGDEXib8s0VuACTmAS2Svojkv/cDgvxB3ww
Q8Vhtu3yG4oli/kR+p6bbRsSTxPXo+Hye/RYMVIVhlvg4zeBYzldYAKJU9XF94Om
T2YhtI+6+4dIZjGC7SgKNGbCT8FuYyBEgLQ8m7R8wLdsgvGhYqDMSZCMv8zDbDjc
YIJwhnQC1ZPgQDRVZoXAQiBV2q6+zgEy4onG/xL07KExAZQ2upOq6xUi5LuzzvV9
`protect END_PROTECTED
