`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtRQ4je+QY22+o6S+NQrd7lR69pvY2R/PujOPyHQw/KRdlxwIhQlth+C++QVo1Gw
S9uIuHgXbuSVhC6+/54AXx9tpV0oS7QiIOVjjvCnrr9P++5xd8PJtW30xygMw5IW
W2k4ArPC+Zzf8PZn6VOclv44ZGGJfFNIe2B+1I+VJ92HbbwKnygMrp1SAwcwiKtD
TYox909VhegNIPhUMjQcuTE1wHVyHX6hlU3ATPuNEEfsU/lRLfgWDYuHs4DytLCz
7bQJB839IzXfh3vaEv6V+m3gUADx+juPYqfVY5hf7Nz7TCZH8eahtRZOumG2WwDJ
qyaw01fg/3h7yDTqFJHfmhozmnWjnYmXTtJ3jTPUpjrrzUwc6Ek8K3FxVOTEBF2x
e1lVZBx6vniq+jZ6a0w4gg==
`protect END_PROTECTED
