`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OuxnoT+0M7dlOoVhLm5RiY2mB6zslkNn802zn11K/T0rBXQXgcUIIJbjikEWEIIt
6cY9kt0SShD5gl9HVb3WLkxkBh/Or0veIzOqKuiPqRbtKlUcdFQPO5fnGY3nNFwl
u1lcX52h/KaJN7g4lTRxlqngdiMwZdELnxcM+LQ+5iAUgNmbuZaSqoNnEGHRnZMp
iA/s1jGPLMoq4g/suY9HNv2XgUEbN54eNThNE/w+btAKR6l5AguS64gmMLoBKzk4
YvqFnLHOOBNsEe4XGvCe7UVqXtzHm49muM1tV7NKTlUnPx6aAuA9jnNFIzBaF6xz
MX6h6vKYqreAgZKyjsV17SuOGrGopJxrYcoAYqXZsdGQmBDe4QuXC0/c9MEBRl8F
j4JkHqFTcDqyx9eG1FKCWXHACMJMwL6K8GCtrAjR32SlIrb5PfZ9KYAdJFWgsMb9
mWOXQlLj181NLij4+Ynzsf47oHRRGQW8DdhjblRJKUqQ50q2MtuYHquxbmjWqXtL
EASKVRXm55qjwK2ApoePbYg7KIWIsx3dJhoHmkpFmdyfrR5y4IBgFu0U5zm+VNlf
5Sqgh/1A01jkkpYWiFJgon2OApqcpzUza6rM4889Kf9JfNsb6DumEyejuKe2YfCp
ma96PoWMa8NTFrd9VzIF4u0Z8mgS/Auo4/v3t8K24X9WnmfkmrpfP5AX8YUUR4eA
7cQcqhLL2a+5nHf0kDSEvS8g4hN4R13aic8cNAuVdV4zz4ZwP+9DblJKMzC7oE14
cRRkk50IRaO36EE5A6EtLkNAnVcXzj4SuMxa46aSV/mc9UCYT2C6zwueanAX66TN
tvkHfaBVPbf067RlXQvoqRnMtCdkVyWIm6GooFh1gw6uiFZaNafNq8976+KT80D9
0sv173iUE3vzWgogsHeHWWyyNHDHRP2kJJzs9pZn826njiD5jR75MnPMxaexfbu4
kxLNuWTGYw0vd0FLS2AsR+bXQJyIzf0Xr5HyZjJdDx2qFUjz/ea3NUc6chybm7aU
+NlsAbKxgmu/8lFxzx0aOK9cI3goxW23KxwUfBikcqhPzJjiGXFeOVFAxvuee5bT
xgJ+a5wr0yVNdtHziVKVQuHzq4YIOeS062RCW1HV1Y6VpVK4Lyrn6qr9R/L0tQSr
C8v5hoiiWwYeOPSLgf3Ul+t1hg6v9P4mcOcA34FJIAW2tHXgOXtpEIzwlVcX8TFv
Hpq/iKvJGghfexKTi2zMCjH0e9w5tFnDbvy146mbxry/btBwgvQwTHBF26GjP5tp
oXUb8cXs3B2CdLVOdWH/exg3owt6rfNPinDGCY2lMqATasMzaV9rp490esfIMDYR
N+J1+9pp/5ks50PtnIOXPutbf3dp4t0xvLLEB2jOt3tSXhZm3K/XfEzTIuNsT4pC
`protect END_PROTECTED
