`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5x+ef9bidvo4EFWdUKWqIYrHf8HwD49arLHt0hWTomOtlmbmHfkIs5fy8SJXOX4g
sq5O76ygNosm1Dd9ruHdVKuHeAsfr+EJe2fh4pKg1x4Mc4iZcQDOYRAsm9SGZ27u
i+8xeKKHpzgszhChlq9wX7phKf7OJuEeXcNyW2xYchKhK9+ue/Rc2UqAsaGQVzMY
G1AU0O2KJKXqVjYsfgd0LPovsLPjRLWNfCMDPPfyfQrh6tmpi2wi1xRLWfNNZIS1
YWm9oNp6F5QOiQ6nID1ETtsUvQlykaaUQ+I4iqrp9B2iuaoBqboyGlYqt22/2r8h
l3cy/naIs+mCwVdw7M5ObyYshM9jzVbKz2HREd5PoZodKptVBY1jq43Fbv87F6ih
yYft37nUInGdHiwGsBeJSFrfUkwnrhET9b+tHlp7TpQ=
`protect END_PROTECTED
