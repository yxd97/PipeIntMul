`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbelQc7Jfbk0gQqWMG/5xQNKj58mEgtYY3m6xUZgHJALxDMfE/jWmxKhIbxzket+
3wqJACgvEJbfVe6gncs4fdCQbj+utKXt/KCgYq14TOZt4gPpd219tIEa5QfW2rMe
yp5El9uAkfdrpBT6/fL0qfIqGZdFB1vN5rY/1nuUKihms3/zK3aex5HmfWsweaRU
IJvd0kxvDFMpnexFPMQpkkns730ymmkRCZM8TbCFxlpiJPyjU9JMpmd4pBbGzR+w
ZdPSqb+oqzSKxWP10KJT2gM8tTz1qB9LJHeD8PQa9dlGAf2XJxpfQT6tEZy7bhpv
F6A2K2RbsZeSJp9L8DkOGA==
`protect END_PROTECTED
