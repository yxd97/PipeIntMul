`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ms4b5cxX2D4JGu0ONGJpGvfggihaoZglH9TIC0BLbfwgnKctNsTPBLd4bnFXNwnv
vbKZIIEQbnmjWotlSNb1Emi26pddusmGKkEdYZSLQWvjosvye1MhKZYYyBA54Ysp
s+WWgVLPtT58yPTtbMss6XfvFFDybqJqnJg+qM7qiDI/uOvk4cKgcHKj+/n308ss
p0URMJrtBZo84Yh9xYfoqth0QD+1wYcPduhWSWPNVcCfshPWKk06QaFeKFkgPzwL
e1zOj++pGG72pDRiOVoud3+myNnFy7OyY/egmSBUnkuedQItuWW5OeiD5M9y8BqA
SHvgT40WUXE9xX1h8DPmGVizgrpivYqTvqqEGtgsr4V5wt8WniUgdIZgnmznyWkY
8NsMuVZ1u/WOsZOs0aALWF+MCRNBJ/S9mhDzmaW2yXKvQUke2TuZl1i7CdtYihwI
NQwRgh1LMa1lKk/B/N1IkRdrAk9tc7jEX2+9OARc7SVB+jHrs9rqQbCleKSprrf7
h3E9qfVg/aV4PRoIPLC4GJzBpYVEniu+14k+y121UNROkZZdnQPw15qML7UqMhSD
uqMbTS0zFvkg4YHwONN56HaUzQbPOEyVgY3U8RJfdk2sg4q7DSB9Q4qiGrkDnDmm
nzbyPF8URdk1rad93qgKjv3xVg0KpezukTHanNpzKvRPdKj8MYsJKOJDjN62yVS7
JfY3P2uJP8VqB84m+eqQazujg/wJxnpmdTBeD/bdiE5ae4WIDE2+fo0/lgvh/wDC
AMQZ3JcPr7YOzYQFcLH8Qk1g+AX117Rc+41Wu9HlQRSaXkJBxxwdKwwEaQwQOcXX
S++VY2aR1Kxs+g9bpkLM27pHVU/PhaP5e9iuJkBs13CG3kf8aR3YuH7ZxJRkUXsN
9ZGntTAbMPAMJvAN6o+iw6JWAU5yFfLQnJxPUxEmrOVrE01xTeHrFfeU9MnyOipj
f/NDrrvqJO84GSUk28xqXGQ5q1pT12LTEuMH0r24CF7UCulkBGFdrrIQUmxYS3Xd
5NTeL1R+BMchnNIAF4DCWFAhj6c+P472/fP+dScp20eG/iEDCEGc4zq3j7jrB1sK
idMlAH0edossGZc4Xc7anFmE+PSzZ0Z1Vx7j68wpYBJxXbOTeu2+eiR41X7TwUZF
95/RYcBZSDzkFaAFlh4H6YLN5w3WsgJKSVc7rG4qVC04f2utGb056a2g4vhXDW1K
t+Bp+ytqIEfSSNMYQiNFeh0hkRw+NOYcpdzTAG9DaFsnXMitVQLHQZ4KsPpieO3W
5hDlgi4sL4RChph5AVoeBedCnXtmUVaFH+eerUHZBWtvolq4Q14a1WP0DC1RwVJM
zg55+xprBc1RJ307NmaFuwxaA7aOW6NJHiwkwIbCB4MoqQQFQ8+uerJKxw4kdFph
7/XjDFKtFZZu/QUpVYCZcXOlzQq/2HZWpjbsn7q9QhYn9IJYvWjDWc9Ck0DlJMiW
AdqknoWI/P6oqCCEUEgNCK+CnD2fenSO0dYDIi0EBvQW3GTEr8PVxN8J78tnRUog
+BpgO0oMJ3EQxPC57MmNjipsvH9s3uFsm/NQuK9kMkwHPodnx5gOQSyEvbPX3SmM
RZ1Q854EbaIW+Tmsc5HNX2LCgnYYVKfLIjaKAcqFtuYXKNbxla3wmL8At8Jq0cmd
RdCLt5TnrVU/GpJMNPDzJwGLOrDtf9wazfWt1Mg5HB2oKKemEHvH0oPWdwr5Gg2t
eTfvnEv0+fZRXGxdL04i23P78aVSlh+kQxRGV0xxtSIGlt3kCIFd6V0gD/BGQhAX
mgQJ5KErLdH5K8nMyu+PkFHR5VwB7cTfnquuDnbgbQQ8z3AVPKNr/Gw7iM6bWW+l
RqP7Vfcqk5CJRq14n5MkdE627cErkeV/1HHY86l+kvmzQ/o8M7OZCVLFaeoqtl5l
rkiHOlBScU95ujgJZ0udD15I78w3jh/APnclkDry1Cd00B15e1Bu+ba8qR3uPzww
hbhhGMqyilgjzGV91HKGEuiiO2Zk6tTPnocnRfEW0MjCmEAmn2pDqG1x8kvJuJd+
AyVRqZGAl6IirqBWTiQ/hIY6h0uqOnrYwFNeNzlMNF8J3M47Vy+h+5GTRv+7gKfL
hk72pJXpf1P/KgUrKkCu3r83nA5CERfPDj70/KhshkEWJF499wBmZwRHHp3kSw7u
5l7j01CQNZigY0Ceo4Vp7wOsVK7kX6leDlmasDV8TYY0m+0c+ce9zCS3caM3HUQ8
v0Kb3PRgu5+hx8e8C2Xq5TWPGMSBtVhlkFA5FCK0Jp0cgwf9e7aN9nY6CEH2zlo0
AZI60L/uXA42VQAETqt8GdizLlPjk+tAlwyR7NzEX+7rZrACt7B8nIrNXHD5gSIA
HNwqYnnFg313mKRvhYLY0bpap+EHQHPzXZA6+TtTZqxxV2K37EYSYgiJiJX3zFbG
rhO3+zgHtJQ1udhGJvY+V/aiZOIurnMGkz/X6CVwkYwxU2OuunH7KtsgCy0jneAZ
2KJV8rpiBh0DLTYLavqYEyhc8Iwo1/LFqhb8NmgeSNtZRAijstrnKiWHsf2wKK9l
9y3qwDUiIrofO8O9DiK5ztkezAEQnLoQlXzTAtBC7wLURsWQ9b02w9UDwZruSqOq
TjDPoc/HDfjgChBWxoGXuNvBHBXgccybMgrW+Vt643Taz7VgeQY8Zxx5uRjpugD5
+Jo+S8f20mXSGzl66hq5T5wRPF6gfGzPNAUQPEHxnPXHNSIoyne3TT4veeeQNuV1
pKTaYp1NWFip9DD4gXIDNl4O0WVaWYIkOLN/Ed/tMq6A5G6ltGGSTuShO1Sd4+5m
M2MxCwhJwnXOygrAi50/0GikNT38DdUUHT77z6A0dAqL7U/GLaOl3x6lgxw4yAYi
lJZpT35DXpojbhyexljoukRXzKrZ0nC69/fMPNfgaNjK3Y70u3ouKsydDdKpfUFe
iinBV72O7dxMRP8mEFIPSK2p/0NwFZBFXoljWac1Vum5pFR5OnnhkNTvoboPOlbB
1PfzSxWbm4e74CSCr6NgyhBVVaRrpEsFCaRU4C/cSredKu0oyVaNLhtVLxKWpE5P
YykAYXs1v8KYq1XASJk4Zps7ZiADB4ykPvlXGxUEGYGMVdVxahwSR94371VIlwtQ
rl7/OuVWbQxW/FLM9WlfxvMjfKhUYyBtnNCa8J/RXCZXFl2Jx2Wn79iNorr86swL
RflyAn92UZgv4+/AJMiVDxGBFhkdYEpQpXESyqXlbCiKpjzTecgwsyUHaGv0Trvz
chOfPSMsIx9xG4T9DKMRD2R12x4rPWAorZAKKKi5jPBmYYs156EdfsgQh72Z/oEO
yqQkimwaTH57DVaPWAjOqYOE/wuDQXvjdaq/49CAnWFS1YVgSDn5fmgyzbeegXg6
wp2QE7D1PnOSzpUDxlb22GvFnFoecQeTvsOT6mOEufv71FltW9glMAPPYAui2j6b
LJAnopQxpyedUh+GL0RjgK8U/FJUcBDNQOIDumRGqpY3/E8ynBpcbsWOqS/Cm65J
MfWSd4gkOV2RqZHnLIp4JEBGrKGdlj7jJRGDNqQhqfFGxa/LPKFU8g8uoWx/tLC3
5mGaiPUrD9v+07xAvU/SlNwy/2a1kydlHOTVK4MeI5rKNkVEN8asMQQHYoWrC76D
xCR6X/2s/iHfoDo07gH2M3+X1q4+VhQS5XCwW9DiEEOg/BULfo58OV1rTfMvSY76
dmgdGyt6X48KmzqrpSgWnNPFRlpLvw/kN2fv4sMvadM2m6kBTeZ+kkD7M7RVBfie
eF2UZ9XlJfIycwsW9QGhSgJe25VNvcYkvEhIGs+BBviqJJroEhCHIvrf5OUemoum
2K6tv6L42wgAv0/PB6b+aDx4fmLDnZlQSHgeVxSZYPttQbnTNaNXUKWn1GscHSCa
yEIn+UbG309oSNsJ1lA2xG2FhDTlvCGURDcDfZeLpGVv0xgP30nlnrJGGpr8cuat
KjlU1CoBpF7iqjGV+x57e31bdHyW84DiBGPo5F0JUr/IT9SESZUFJAgVMoXCu4GV
v/oXh5a3bMLWFBptu9nKPqsn3LHc5CHRJ44t07QVO8QiGGzKDH4C596lPnycLWiN
3O5+BcCmXYu9ZPa7zJxZ6qPILZXi5U2xpxQqu6MdrK4dlgiFQOedPfQT0iIbnq0w
fW5IlxWa43iUJQVsOhKSDf4iWgN7QF+NKjtw9RlYdpJmCTQtJPbXTZJl6xWV2IgP
DKFm/g6I6UjF6iNJed6wV0soLkSJUZhcUZ2x17OAgeiXMJA8v0hyrjSiwIL6bJOG
hkSr081tvqWqjZjdB2bFx2z/Qw7UhXmcnMRTIp2tnzwKZvwPbA7IXFWbW3bwkOKf
wXWJgJC9lN2MmBfs+V89mduTj4K4nDrYf55i1CG79Ec0HfDW1RphcsaX9f9LKdcI
nIfseF75W6n//kqbUcWpOh8fcSiMYYC21Ru6oPHUBeus0aYhvRNJyteWggA4x4Vb
SIha3VB8SfJzVrnU4CwIHWl125WGeuSwgmOYN95BVjvd3hFsmBtJ4fN4yw3OLtHo
WcuJ6si8Lnm7PtW8I0utAUJhemwytrm4Wcj9XRuQgsgCAVoFxHgi81pwWd//ZcOB
9mF9oxyIq5nJE9XOL6c25OT00yvGELHfodl2usVaKSJisH/PhRmJEZxyBLtbnsuO
2xQymyvA4f55uLKEGJNOrtWRaa0+QmXpiMeVvMjEzh02DGVi8E5+xdmudehMhMNk
kyPTrudbfFalNZEQSzvM+fmB13844fwukD9QiT2M2VUAFaCem0O7hXdLxcHusyLv
p5DgyZh+j7bEiYSC96jMi2oa6bCItwRjoze+j015u4eI8xmxQAO3AILXPntHMau8
pwv7u5KFdNYJEokVrFmOscrSicFFpEhqqhFvkAegHsWOR4oIqx6aL9Yl8lKaxa9C
EXCWgKpPAa+47i/EVRQkq5zulm7dJeHspOXtFotrLmV3utrn4GRgCx9iVV2hMi+3
Xmc3ciGcghXjUJwpyg8A+Tr5dhhl9swIdkoay8FwwOwBoZiAUfVm6e1+CkQXNpct
Jaif5JGrQRYbF1G8okI0I8FdgECaX8un3K8kDzQocdbzqq/IUIl/eo88Jij7b4XQ
9qhZexMvwd5etUWuaSbys4UMWiVvDrccHVY6blFlFP8/y/K82NHzFgicGwiPNGZc
aPlbx/uL5gzIUArfDa2x3sjaKi7CxmXw0mJO3P5erL1qt2/EwS/Dl5fwfyU34u9Y
gNU6vwZGMxEM4zxl53YllI2KQBV1RmPgJ9JUnQm+b+Hydp4AKWKy9WviZRElQ7Gy
MqL4jGm3IJmg6TBjlrKEGcmTrf0eKJswNRGFI1BauHmIl0ZQvrL/5P02fBVizFqu
3hwtZ/pptGJ0J0U29Xixqzs1HD6Nbb8fcBJ0WhitBe5Ny4olR2I/mFiW8Q7TCnTY
agXuwhyXt93Gz+BBf+DFbthKNSP/1XZ9GouAYJ983WBS/vUeLVIEmCb0Tdgm1xLY
FC/5Jkjvi2ABZm0lJiqxJsBfEJgkrzkdrKZsrr/CV6P0UysBmfhw4DIm4m6AgUIT
MlHR1lQZI0x1tjuGO+L6Xk69Deih7gD9Ne+ltfmTyVU=
`protect END_PROTECTED
