`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsBR8sAfMJyCkh9C/DYx3iOyS4dorfAGO+F6ZON0ybGXyK+6fwCauXJk6vJi15xY
hOqcR9rrl2v4CTlVRScx6yufyKCMLSIxsRwQl3JH20wNnA3TcBaxmGzfR+UPsn4u
9NGpVAP0GYDstX8ChwFwHRDgZLU98a6+k01C74BTFshhm4+sInEjmfnV2qsA2PxL
euNJ8SRLJ7p5LClxyFb9VkuD+I05p65jcrVoHIY9hhpo9aDxiazazXkTtJ8Lrx3a
WRPbilG+tLucFltsRFJOPyT4sg7Ztr/AFnz14ynC2HUu2hVv/LTVTB5rnSOwcpJc
jn59ugLq9/9m11Edlfontrq1p53DEEktLUHEMekCVqjpd6PM0glKqkijVubmKYG0
qMpOGBvwvtjQTLLc8+3L2clEz87M55oVFI8+1R4mFm7W17KU6iKydhUqEcUmO521
zyVwKP+CvbQbjOHnjPs8wJs/HFHAb+juNDBgLYQGQJE5OK6MKxHBdwz4of1HAacx
Bb0IkIPxVcDjHjeyGlnwB6owQY/4IfA4bsF1RPK2uxoG/o7y29UrUbHxvleUY8cf
8QNhw7RkfaP6KtVJwBMN+d/iL3NpNkHgbteHqoAz4El4KGQXQOx8nh9dPhUbQmWt
wzAuFlCqbOrkG/B7OmSOt/EOkbpsJlCPpLoRsuaCrhfRZeAgAiY5wQZwVoii6FbN
lVozRt4FcVY/QCyMy2w+rdhdVtnyj1uS3LjutQkKb9SRUZ8gS+G76XVuDOhBmXae
NislYURFBgTq0Ct5IrNL9Ut76rRDzTkpOenST8bA8/J3A+hlNFlSm0NJmDnLBmtM
I6b2s9nvBXmFzrhVNpXcyEDnVdu7cMbOvwWn8e7xe7J68THpLG+GCmRVoWxTd/4q
T5hEheF/F+OJSTffIjjfIaw7t89t0VB1rLRvxkESWMSaeEoB6wRlQySY9TR4av32
pdG67PdMfTcvO0JdEElZmVKNbJDeO76jBG0bmJuudnDifWa1Y4EcSMrhdzk5rWCH
VmxjUvCCzhF2dilqNKl+AhkKtzLHHGUJJGH7Qgb0xeWONvtn4aua7kfpp0GT5d/M
uoCACUXTTb6Ve/GLEMcGBtJUW1g6NtjKFO2KGlk2TUO/HtSCnGzaRQPAH1w76wex
Txmo8Pi7ZYiSGVRW2u55NCzYmlFBDW9FN2ctVwjdXT3fd4q92qcvK0u47Bg3J+VU
Eeoa/Hw72UgNSq9PzghRPtyjBkFO0CDnzAjn00CUVedtKjX6cvzUZfHNrT1i5oxh
kTYxk0iKemYsBj+vhsWHkBw2nVHsoVazCE8ld65d8A7FFk/rM6d+JpZbkPYGBe0J
TPXFBy/bxSLcPVbz0quD3yEMm7tZXnlV0CagUWuO2dyZHP6Df7SA+S3Sim1S/S78
Z7S1fg4CGHcP4M1BmAsWQJron2XR/r6a2qRTp1WBV0KLDkipw+ogoGI5FSHXDptm
UOvVLH44gbzNxzl0r+Aeu3/oBfV3bp+t8YFsM1g7RoljLREA4CCBrTL4Ct3eRW7O
`protect END_PROTECTED
