`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o12AYBczXI4+aWxbzpnwzuBcLkouj0fKgswotaZ9t7/hHqqmBCqqwe3IhkXtkbmx
lGXZCwI13IS6v3fcoVfsw74YBUt9h8I3abAESbLXZwKUye6L33ctlVsJAQ14vkLM
iLh6eKBi+hQE2/FQVjQ8YdengQJx1Lr/9nYDwtz0vh8ARMDUDfadxTtOj0KYhTJo
r0CmFoiFjzyooQn2ItjSTJeZOD6XSLxkTbLeDmPShcPOj2IAtq4bHVfispS+NdhI
Hajs9fXyWc9p3o7n8lr5gK8cHNVxswRS2Ix6vFj/7ojpHGLtWbjAsaHAaCuFzUW8
RJ9J2ox/YndL5X6SHrx8Wieb9k42xlyPo+kywWBfct5mrD6jT0ufsv8cI/eaUHqg
k/Y/wYLJDheQgFSolApetITf55pBwlWQn7pivi5i0aWbVsZad8hMOQP2PYQDvikN
moQ5+Mn+c2LWzwT6K+DrknA8UAO6DVzYFoaumfhePUAqIoXvNAE6prhlYmkhh7Ib
gksvxu242K8NtYyE0lXexSICqSGHII2/3bdjK04f48nHV/bmTWaicPi0RZo6YXMm
Pxj/Vc1sYvmatQW2H9GrOuWQk5khUi4MKZDV2MlfHNP2oV5keEt97L6oN/yH/Xqf
vHfUU9raW2QGjM0pboNQMkzGTzp4u/gOKAmQl8X7yTHkNuAaz90/G+8EvhSUIU6J
uGxmi9XzSUKOsMFV412eQ20Q5ZWh7M4GvSVALosBTIGWYeF0z/eoN4etNNCDXMmQ
XcjV9qo0sZGPFfXIK4WCnjKw8X4GV+mHHA0nYtG3mcYZlnpYf7niSsoJ5KuthALl
OSUIqbQrR+NQtaVr8stp56glGW0Ejpf6VlZHkW5xIPxZwXxCb+1szODjL1Hi19BA
hnFlMp6W6O4bUma28nozKlMpCU3EG1g79mAi8oEEdjTo3tGTRKd4b5S3/M+AK5dY
sK7R6k6VJub304t9xz39pfqL1GuoK8WC8BfcdcIDw5Nx0ms5SvI4TYW94/y37r9N
geMIdavJujrwr4Fm3Bbfc+LRnywUQwcvkVK4zMdsqUtSnlgKy1yYcFnuOIMVUdB2
h8x2/syc+LBA/JNVeJwz6ZiqumkDrXSfnLL5kVbPPy2QvrRkuPitS0mShTJNUniv
6OQ64IpVk97P+2a9QbeFzR1ZeonYSCUYY/PbVK7WtN+lHscP25aOjvp654WHi0NK
8iZTp+mKqbmk+TKDErAaK4taASFSefyob6PYvUcBMuy0VZZAe4DZ26ZZZshVo4ou
g4HWQSmbE/rCQsi6Y1syOzM6p2F2/CycOJu42xNPhs3I38IooyeZ8nXiPybf/sDw
ZcuFzsrEZpWi3bZYqYcI9Q==
`protect END_PROTECTED
