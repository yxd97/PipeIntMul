`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UjMx2rhaATSX9eDMSQDGYNF8ljflDPpRjjRJjMn31Pd8VhQTmc3QDVkRRDloD2tr
NnDnJbzhOZ5qgeIhWkgwt3t8ZV0/F8zmbPr+XNzRAYKTbOdpBdB2U/K9dB8jM27x
DXpsJNe5vJ7tR2KDga34AnAyD88vY1PbT19/l/sAzD3DFiCVsrruFaMpHOXRJsZA
lnHgid0W+fEV1yREtrUr6uKqWbcEROyZJLYQE3PN7xFjMtsPR1jBr4XKjsDE8IHA
DMiv/wGemfs4pDAk+g0log0D+WgoWdWF6UnNYS6RWRZayBuLJSJuiiQ/eMycNUjd
YqExazKCCPVI/nJLYaPvC56sSqM0JcerKoMQ92i9xyD+kEfcNU1q5MtXeqh4/2u0
OUPCk0EOyTibCVHNUxvg8xQ6eTt6JY2HJu3/J6Py+3IQubYNL7qxZFQOAB9v9GTE
1EjKAQIxcNqRfytx7yhHcFgvFoEyzexVcLp6l6fplM3IqTHPV5laCaNy4lvDaVqD
FGYqjzeNY+qOv1rTf/gbS3tz/3RdpubnVeVbPinDHLJZnILYs8uZDRkCSnL3F7Ep
vCEZePdCQ4KIlUnLmNhivgaIsayJI4n5ps+/PvTVfGjOJSR/niDHLNZxYnlHtkr4
47D1G0IKVuUOXX2LmK/ynA==
`protect END_PROTECTED
