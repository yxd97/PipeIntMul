`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O9cT/jNqXnAHNWexCJUTc6uLfCAfbnzOu5TCu1voPhXs59NE/BJ67l3IbZIKHxjt
foze3AOHjtjVTS2oa6Rr80O2OkHRBySowyYarZsYX2XRYp9HLz+CRh5l3SwY0LwL
St4ZjLn0I9BMvedsVLhXctA7QEppgjKYB3CJEN7g8uzN+txM09vSh6mplCXBeitX
Bd/P+Quy2fGV3ShClj7M0DOQc1d4mQ2s8KANbWut+3AYdzkRuLULpm92vU4gO3vd
oItwwnUvC+nKjWH4BzomiifANZIGGYtHchb+pRyYDpdurPj0tOrxiPfOuyYRX++j
uIFYR6wOVddKSvTaXq6LXhNXm9ajyeq0gsTDr6088rLQRcNgjxbK4CzGc1BSRTJJ
8woox2V6/jiwGcAqB/arxmqHf5OZ1wJlQ1o9eGCAsVCWNuBVUxfyMuzQ/awMPvgg
M03ZHZU7RrAurhHHDwFtLhNlUBQ0Vk7dIIJ4h1O6Y5cn3GnUoXEJuFTse+reUwoq
L0G20kvBfh+SK3eJK0akuOLzzUrR/hm0oJV8RhKuX6KQetpSDnicEs6uX1QAXjkv
kpI3z+8YHE/ZRdgvZQ7v7b5FHMlr7Wx7JcQWa0razlx+4rn7Wf/U4dURRTyMo519
DK44BvVIQ5TiP5mhL3Qcv0ldRFsErcuKwwONVvXaVoeB7cc6l/xzfW/hP61UaG2S
lqT98tjUZwahRDqkJw4uVwwtGoKVbLHZiLTy3wvuWf/KY6O0HsaYB68yS4DBigpc
pDm2+nvI44UoQjqJQId+m4GFNmggEZg52chl5EvCsBN9joB1OyV50Z+indBjbuKV
xbw16HS0+n2aN5oxZBtPWha8kxc2S6REFq38jvqw0Ch8icf1L0HH6u1RiqFz11b/
fD29uarKvjfum8lRCWQufR0cgeJOQzOiOvBn04suEblOEYaiSf31rGjx3vcJb0xH
tnwY3k6GC0CR4+P5ZRfdeXuEKxJszwbFRl/m46+VMo2twCiE+XxVMzY4hK63cPXs
WU6ND54/2ATB5U0YsOP7GeOIihffeuFjKGq7/9kY99vQ70OOVhrlLleO9leUkTfH
SOmkjSVhPneV9OO0STG8Rid84YDXmVB5y5QWibSGh9Vb4Ad4c7UwnAzOOsqHnbLb
Ef3jiCnpuhZVT3gNVTkeQLRKU1Oo/NmuY2QpGHgvUtCgzUldz5Bsj0XKSiOZb6ly
kCgsFlFbCegmC3VjpsY52CI0VgXhcLLPd4ioxRH1kfHovduBX5OBvniohF2IjOgU
n6CHYGcROC2LR4AOSFN4417m2dzlDQQZ6ADJomLEMmwpoRGSJRW1UFaHE07gLEic
nptaR1L6ruivJvS6G56qJYDp169E1olOacboRA7yOtUro4NDjCNktFafp7+4RNHN
OxfkESXllVQJEq7ZcmTilKqFtd1wmOp2IzAkRNMiHzza1k1ZOermcGZ48BhrRm35
6xIRCkP+/5u5ec0ElHykTFhMv2M1Djtr9QzTn2l6AGfsqQGtbp6/nII/B8XyK5IN
uDRizocvcmNnhJU6I9evtl2RGIhB60pRfneC1UAx/GM4EU9hIN70I94Gt1L2yIS2
LyikDf3iDkdW71CBi41BLeHsvW+TfzDgmBMbe7skz54XAMpe/bBHwcJdmvaXraKj
FSs8SAwbCK78C29vExxlAkjWbJY4z5jS+gKFS0FE4kB5J7fl9gFWoxZjq5ZOSrqS
pmjqeYs3fJ1qNMs7v5t2NKkzLpL4h28g294Zk7MkfWBjnjFLPImmmTivvqjZZiRO
q1BmP9FF8XkL1Q8SdsqdyRlJnwOV2QA5LxwNxkMcFDmae6QAYY6HJsEoUAFDxryU
T7IIdsCc1Ob7QKfHYjcvd1+v3WG/xFQOn75GA/136kBj4JxTZjnxa1j3fIsTOpGa
v/jxJ+45zJzwvUHTBuPf9kWuyN4RbloFqhpmhqlFFB9ySdu5djfACSKHOvJgk1PY
+heZTKL/cPiG/7MmV34LE6RIL5lgj4/jpVIF9oGuTo4+z+gDGqDSmxe69iZ8wiil
SUMCvIzJFMv1cSJjy5CTcZnaxi4qBCwz/yo3t+JxvYz85cNnjJzOx0xOhtI46Z6B
VYPBJE8nC9I7qSeFvam2YvwEdN74tnRsFo6rpennW/5rDFK30SCBqr+rIOHmNLN7
8niSLiIRS7WTazFxYPkYBOp2M6pC26gETeGRF9ORuL92zykChMf9izcg1guUlQKA
vvdkefwgfpawk+vf2tSMTQtfEHnN+1hVjuWuyYjIbTes0AgSW54FXNn9e8DctHiD
r3L9YScKXRz41sDgRpzqzlAlwF99R2N1ccdemLN6yPuZWD+8HMEvwoU1NJj5a4cC
KkDc7tUTqphIDeMu/38q5ZWqrUUbNoWExRkLpikaPHvSFjFRM8sWdps/LD4Kay04
rxgzVpueXegnZ7HUPC7rtZzy7LaNaVJIUNAwWrEamqkO6ojLm/940TeEvIicqKrT
3ivlo+XdZo7OZUbEO6n2d+wNHtgIY8RVrvb1nqb2lx0JeL3tvSeT1EQ8atUSRQkw
quVBq+N7DR5FeU7atPnO3nDeyutfE29sWqgYCmMmaDUyIDao6bqsaAReeDmUS880
UJgDFZB7JZOUejM1FplZTWemHFiizVa5SK9nY1j0KLTkEWd5G5o02+u+V64Nx57t
+oPc6jKfsPruejFL/Nl1MGtu0kU/4ynXp1CJaqNugXHmq6Ouu8chc0SFsC8GoYpg
cJE+1mMbNBhiOAZO+lWHgbg+kWGNglyQM3dybAzFOzQ5NjdSWJnnjf8g8LCFEyZp
QLF2LxWumPGOGl76dtlmUoR4OyxEVfnfaY+9j06QDa1k5kAB3VPE6MEaVbfv14nB
oxyWXTwGKcggKF5lh4gwOLHt4AOXePNumoW55ycmLVmjM8H33T3Ar5rV8rcptB3m
/l4lz2ijcuVJN+5auI5PgGs65ts+ntCn7paMchA4MagsEQThNXYYYDTzaSyf9U/D
YmK4hUgX9+OPxpIBI7+Pi4+comqS1MKbSaZto+PvQGbugW7kcNgmfH30sbTLNUNg
4Gt2VEZPpZAJlpVTFq7A/1rOOmYkT0TZYkecg7Zz2nRgTgrfG4b4yewvO8AHuunE
Z1Zhw2jncbrZG30I2TCZaw017cf3cCjGKvuciIId5VrAKCeVMJifCtjUmW5uQ2j6
+FMWYESNV7gQhdwFQEoYFfsb95z5CeFLA2a3xxGKqAZX5GL6MWbfE5NW0kVQKqyr
+ttuQ9OXdObt4anLz8f5yf2rKEn9Xpm9PpF/Els1Jk0Wk3gPoANwid8A1mnsQYUf
51yZOPqgQkcKz6JhYUp8XU8CYFppQuWJuJqyw6VP0g/+L52dtE9heVGAI7qi3zgl
FnrHLeP0DuQHL+MSIT5GoEIYr+VujUp0wlxswUWIhOpxFRjd389ZmQXYvsmE1IBC
TIzzT8jvuEMahqOneyq9+nA5gS6cH7BR00X1FlqLTr4F8VaEa/7II30HocJvNqVE
NYGH9cLGTdCsMjYcg0QQmashMHEl+0HRNABA6sl9Wqek8/Kw28aOXdYIAFFPdTEy
TBzwlCOODioIKZFJDN0hvmMonxy1qCDantI8oBNiDzZZF7JLN5SB3mRAn3iES02s
CR8GduXRmMWNr88TbJxE/KNvdKZ1qP6Akp9hi+gPg8FnxA54frw3pR5T/YquD+Ap
QnjPfwvWRmA7oEFHvFrhI3l2QVF/e9pBBlcudQRDZi1k5lpNYRXQl5eI0tkaIofP
7SkBupktKSzUkJKjG6vIXIEEhdH+u0bjNjx7EvpIBoHThwUkEiVM7tDU7FNni+mn
jtpyyd7Y0bGVXxKPXPnp35OU/mKo4H+0nEV+0i7g+v0yNjOuLBVPAIzztwm41KfP
XFS5gqm0YsDKMXS64fWXp9YmV9Bce7SPJxPLC5x2bfWfk+u4Y5PUgVlgH2q+q/S1
1BvG4Rh8PSRdofcRtyXReqTu3dTxBAMPd6VzLg8tMCRiWbIyDR4ehAgEx7s/GhQU
lIKqYc1x1XbXqgXw0wXiCVp3L/d66ni9cDPb9XPl5OPzel6T6KhZ6E4qNf9Ud/Uf
VFH7jvUQxBxLqIeJS8YErnpPINTfgqgWvF6dT8+kNmNL3aRDxJ08OrxmMvaBe+ri
xIzd13+jOvOG/KaUnfx6ZzaLXgEmTMQXiG17iRYa9JTEAblV91z82+XZjs4RvsjN
ZSFwheN00GvDe3VwuogsktXrrJWQA8nyi7a8xSwL9rtUveTYaRVCnGL07sneFfK7
qUIF+UlGYABLRmsMVdQ6vKnlYblMXEOrSZ613Fyu16U4Zcc4JNiI77wfNqzyW1FS
mKGQAhjegyqAdpt7MsIcUGyU1iOaLQwK5Wsgrr1EiXj2eqFtH0R9vMxkXvjQ5sP8
fUz2R628dWKqDneeceYz1MCUMm9d14dTmFIn+X86SPM/3K9Ezy+ZqD8U1RMVe/+W
vZ8T3NpJERqCHJf1hcVh86D8UHPQhQRGseVSqvZGnlp8LeZwWMNYD0spVc/a3Z3F
10n93K2WkIRgPdF7IVQ4CHQ5rc1wm5UE3IEbHhNE1gaRybiKKyz6ZGftyxgzD2cm
BN5jOJVLDtA+uLKQy0W7+mVF55eW1WwHPHJwvai9ZQiy0cGr8neFzxyDHfMEjh6h
5wqF7EwHKrcXBxJJkYABjskKDJcZ4BewPjFWDiYcJEXnt6rY+Wa+fnRjh+lIySb/
aCqitkgXrQT0XiF1s/sktJ8RwI6JTgjzo9RVPLIMpHlY7D7P36IYI6HcvJ/jALvl
Pkp3iurBAwHdVM5EJ/svq3mX/m95aT3i85uT9NjDazpMWevdAj5/rNnRRIUf66mg
juUQWRNiarDhmLpsCIlFrTZ1odjtagy5LSDU2npu2pWLzRFreHG843k4R5YZZwlY
sDwhKjhtMj8Es3S4XZa8KAMWHL+rR4uJ4SBEb90W23Wj+ksVmDpnYYjQIHSEH3bV
j3vmyhz+VJzPANf+6fxAa2Hy5+gR+5v/taUR+GSwdOZReybxlidRpsCkEhe3Cqp+
hAJjoq7H0k1e4OFhRUF6ZQlsT+uKNcelzPKv58OfwhXFcp+sGF0ClM7uGGQ8sNor
0hImuhcbAmvUdlzydzCfhiGAQHrQnbLiePs1Dw5FzLChLHyob7WfTlHubeEKumsZ
MhG6jP8fWMJj4Guj7fyLY24SA+tM0GdDtuYme0yk/MNDbpm0WkHudNIlp5v1Tfnn
HXLvO7VcE1LronUEuYtvWD39+44A3hWsajqfRMLBYrymJGZ7sUoqBLlu/v6m4dSH
4XuDg0ZXW4jM+PGBn3XX2Gk+GHa7kiYSNSchjc1zNqnxNbPjVY0/kCVT0+S/QCRg
Tq20ND5zRQeTETURWhABjRzh6bSPndCmFVjdfuvdbUAVIHk7lH/CCh4J60PIH1L3
W2lyJ0PPN5od5iyAF0dzSpD7N9PVsjtP032bDgsOXHR20WLApv6KdDRS62Gu1yvH
vNy7jjQ//dGf4IuWeBe5XjlhSOetnLGIC2hdyPylIjUAg/pEI0vFJhRrcF9HPuSR
02nolc0lXvGjz3fETtOiJdye6B9LTbs8s+mek3H6MDwiZQncZVCm1NujD+0sYnEp
AgbHCF+Hz+MiaQwfDeyzzB5HJbsIKJsb1awdlJD/0P2yWK+vqsva/FUtxZ0yXySD
yIYDQxJBGeOBXlTbdwyCdI+aQviRtrSbEku4eo0XZtOpHSEDckeoasqZf2+RvBZv
6gJ/Xpp0Kr1fNuC6xrKNB8JwVjDhS5wAaJ1ugmJG3ybyvhEGTt1dcBs6+DOlPr7O
ehNgxQ5oPyRXeW6JWkFmtD1yRwZSNjFCYTPQZsfajKHXnSpBhoJlknCc07JU928G
qla31kxeocr3r+9GjWOpUtKSTHZsuwaLQAASoMqk0jF1uAhzWE5RqTgXbxaU/9iE
2lNEJBbbmB0IR2iVYAcUEBFDow1BzXqjOkVyaHo079ntzyZrR3W3htwYual+/P7W
tNLw5DSJKbt/bwzPLPrD7U32KDJ3rEUi18VtFX2KFEVxx99RYmu+eIvCwvtJkIMW
25YLW0Nhb3mRKnUbhzqmxGq+nnmzpO8j5WrvTRp6P2wgrqjxuxEoPiFI3IY+L8kl
sbxS2p8uRxUHBDSqtBpd3rCGmtLcUKkAbUd5zhPA54qvBw7mKAF6lBb/7Vhd/Pfd
OwR1sZUoEHK/AzprTJEtlm4W3ZzvJsKk05jD9H9kqN7vXE0DnQkxM0K76xu7wyrx
qOtzfQYbvfpv9JLf/KTi6tk3kKO93Pkhb3Ptax3jRPUihPzgWV1jeWFYdZtzSe62
NkfyqQ2j0IMM19VrXQ93XoyCILlard0kmyrx9BSbrCYaZB6m7RLvN97rrEYiqtds
wRfHxfOFoSK0Hkp5vgTjUyrUsG1uffkCM/lsVfypjwmV2udnv6cXkjWSUSPyyAPr
TAsQd5fQYumxi1+Vc/kqG9TybhXYuMMIpSOVRE14D49hOVQBpUu1qiDszdsgcPuG
l+s2+ChEihI4v0mObY8ZeIfq8uRP3GTLWqDXf+Gnh5EdHPMrelWL8D2+7FJc3v6l
8pLMTi0YF/jJ51AUKs94TYK7xazJvx/VbJklYrdJPxexMUTprd0drOXv08MoJevl
n91HI3a75zKpSf/iCvuBIfXOay6dqSOD2R5aLu+tn6TBKRdimyCQH1liJ5muUXLl
b9JNkmNYwiCyX8C7hhQ3+VmauYkbNmWkQGU/a2qlh2sfggqFlaKbsjdroXljKQdD
erPAGWVfSIVXKb1U+YdbtMVCQTD8yYhibFifRjWLpBL05mcegNu/Exw5kZw7eiKO
zYBJFbQBcO+fxu3D4KIq5pau5UlyV9cT21w5Dov3v/v5CaFtgLV4d8uCNWNtjiNh
skM3QrktuP4kyoqZ4UiC/GNviFf5yfEU8gjgwv40LdG2wGHsSpJzHfn9sL8t/B0Z
DJ6Zk4JfEAEgiCtNDglIkaETxeantQ2VWOXlf/qqpsV5NltBKrvy4O6OgkqOlUEW
2IKHMrw2+FYKkXlB5Vnd0Vkd96hpDUo1jU7tFC5/81D+sbQFzwXRSJqTYaT6g1bo
sKu6QSKqiwXZcAvQ0OsuLw1kTYLPFW7x7Pq7gGrmtytvj2OdybaNzID/vGLNbThO
8SrDo/3GbQIzQtNRb9p+GG4f8jIfzeNj7y6nVOrJ2zoSQWBwlwywzEJRPqQN1Sbb
DhbSwjyUvVxDUPjk1wJpC5HIV6qfbynwj/bmzc4+DH6PWdlI/kBwTgrmrQPwRl7y
9bQl2dK4PoepuL9B0SCXdiSXwvues2upWalmSlIZwjO8jpKg5exHYHXPLZaVa10l
RfPY2brmEc0Km190H1NQ9HYuai/HeAmOWWPXvJtMuBvOKnSUwWlRqkFUhc+ZScWw
bcOc78PwZ7UY64jWh9JgVLihCwzv4ZPjeRgm+Ke2e34URjNfr+qiv2RwYrkGn+Ly
tuDTwwPFNUUryKcQpFWNodEa8I+PmDLGzA7PkqcE6pfiuczKvpoADnn3av90XwdI
wKo5eXFWWv2GQTYNE+cvzd2hwAIo7iVJcbwfoKaDjkyLa0C8GuaCe8l3uQpQRqar
lutrCXv+h2/DdyS50EITDie6E3YEdyL5Wg2Wmt/U3TZLN9gMNoAUuPFeGLi0u3Ta
5s1hXKy5UkvvbtWqFOxCRc1Acpvzftw5HDlLXh3GuIygoZrUkZLus/U5laeed7SN
wHpC7ZTkFo3tVxymSGlz2RJRGD1Imkt1Rs1Y9ptaEZV5ymSkQ8GfvRmRgEVAf3ET
Pj7hwkD/uOYfDtN/A2aJ4Pz4S348iRfouX7vVCS7HciDQnJSXgXvs0IiDUW2ulJL
hdYKOpI3t6yQYxtJ+clX1IPki9LSVn8UeIr9cGxs/MFWrROD2Rfj1e4s9yOdjPUb
WWlUVBQ9a/vu7SmEkS+SecjKLSfUJJLzYUA8YvwneBy5AmatI7QGv4jwuVkdhS3T
LnkPyPZ6P5f95go+kjFQfkep/qHiBVsGLFVXbZFprBMjnY6Y2krJiSX8n6pegvQM
OiJ8JSTzc/Gdku5H34eIvQ6rDSsfpuuzsMxDZldnC7/ldx/P7/5Q2b8XEoQn5a3c
8DHbm5A6MHZbHp/acyW28JM6y0LibIBmBdEIunRU/oYEyVpzN+B/klXcO7CB+kOr
lisJW+viyrQJ0nMwyOvzVLarVnzhpUkDYIio8/xOc4C0vLn2OC24SjRSOf/EJtDB
yRj81uYC8JvlIDZ63FAnIW5EOf172M92KkFD+UNrdgCJpWfZ+CVrqTFBdNPbbASU
g5vH4BuTzB1/TZTwoZHFKoblyR/OTzKBAab2+onrTzqKw7IQmYfLo6TPI4+qYiN2
zYfa22DN/Cu5XdVorCV3wcsJ1xvDNB+sP2M+C3WO/CgVdsyyWagsD42oJaNp5R7k
v6n1wssgc/TyvOjZQsuIWp4XLW07nns6JkyiFFiTs3WLoCzKyRWP0dgtjhphbts1
NpeZrsnONSfaLQdECM3TGoV2blwFrDbeacxgntnQ/Z8BJXNijU0CfRAR3JMGdRpg
zbyScQRuOUyvFXGugielI6BmL1hZMGfl322dtLT3C2WgUOLpSqclo8jsW3SWSdZT
4SGr3UHRwZFVRty9yttO0+9n0arc19faiGKPFKmB2H7n/0FZu4GbCLRhmZHpyrdI
vQWyErNbZQDfiLhNQh4ptZNJIptmaisLYZ9sm+KHKVer+xyeUAOgNzO/yz5+rYp+
ovK1fm1/JHq9v7GS7zuzBNgjOrI9ESe75lwrZPSTW1IGDnQe3I6sEgyspn3FG5Oy
ejI9ZmtnQMUbFy6zUEHJWpS0cUOz6ly8m2AFThIq50tXaJMVTJFbV2/sz+smyQDs
Xx1OHlTLX46GYgFqCgjflMmg9AJpf0wYpTEgl2eKwkXEPgZVDJn5nZL7hrL4IHgq
Gd3TEUEdfcuh8ey8c9Q1Fu3U37unqJEjKr6OD0H0L65WSXwLNu1lj9xwMSRojRfA
CBEhINMhKRrteDdYqLAJAOp8vNaXM+SpT6AxH2JLf0wjs4kPq9XT93j0P3Ei8TnW
E3bYcHcYEvF36YpUNqZGe4c9W7l4TA0fkMTMw6Dz7CU7q6FFhbeTJDxWDjvJ/UTu
KXEoglHws1iBAZOR2EgR3at2u95RqmRbzfFc6LXJ0acB5IdiCTs8DLQZU1WTlRN6
7eV/Kw3fw1A8yrEebXww9E/5rbrRaY8/lh8GosZIgBNlneer5LtXt/XDo62Hqr7U
JiAy15uVPhH4MMD4Iftj8gvvoFqUoHqLplFtKWzc4t8X6hTKgNOERMnR33EV7fA/
WG6XbS9ju1SLOAMscEd0fwMtH69OiInb78DKJZw9MmqziTCFLNsVEAlkAvtEnNAE
P4Aud5gS1LQGg8Z2cKgozyXwIH5/QEVS9A7GsAaUzcnbs2KdADNQ8MfqGSy1KnkW
caMNFoM7auXeFKcsMQZ6JJbpdzFTJ2DiS8FkfxOuLPxxr3AYYMcg8C6qmZy5C+K4
AOMtJDtD/Lee0wqd5BZ8UosDCTmxgwNvUmxY0qiaax7Zv6b7aWzgplXE9w+8U3Sd
1vILcV6ahpg0MSGZ9CTApQkH97IKmERP3eRLqUpUAk5586RAX1sZv5mk/3YfaLId
xF6nGXHho9BUZWMsMjB7+OwpdTbhHCIkdY4gjh0MIJCjXPc23V6m7IKoEQ1hKw91
5ZTD8WSLlIYYrTB72QN1CFOeMk7lmmqVwmjTxOZ7I/vXWu8gWBTyiEzxFoc40M0T
hUQE+LuUgCUGmr/PRQrwNv4h1I5aTQF2mRXD5fIjCUenJuAhlzGH0rsbxRH+z6WR
7+VP2kkzYtmqlQq6SfoM75mFlrzQEl2IHpokk9q7mviJyvFgUFONU8QP/jy7QVvE
qqVADn9h0EU7w9UyUgo7dbCBO4i4q4l5nAjzUCCA2aDGtvFEKkdKZ113U2Mg19xE
mff6SNmojVQyAUV5Xs5LSS+XefPZRbncaJ+nkv+QaLvhfMc+z4ao274swAXzQD75
LNbLOiIG2ouOGGK9NATx2za6Hm5qfJNyRg169xpLqERtyi2oZx3RrTdSOIMi7iMp
gaPSz4o1WJOG/PItfyzSPeZOaYB5Kb4rSznQPgTcqewuDsSWmzfNbUvwIHSC+cEP
HdoTd7qLOTKjPUpNRik4PA7l+p15tzmVHqpBYCA49AzGfAmZAipSkWkE8xK9flro
6s+JPS/YOp17I6eyACW71jyulVF4DpFbN27fGz/NG98HLO+t/sGye9M6kKb45l4D
VG9XBXYiri+kmVUkSBj5OytS3F+2Zm/bc2GWr0E4lrj8OJB6o+xoPbQei7EtC70g
hGGm7EpWtOInMfb6rAvWp7wa2xqS7VyGI/rGZlhTei4csFrc8qGh3VvTdWOYSLHa
BrMMYbCiY8766eAE9XlpnSqUPslWeQgd5dcdwjo00Q6/EpY1i0Etia5X47k3p4/4
VB5VIsmeVhluE8lTZYCBAi7Iqd0+EDlg96aH6YQ5ntQQSRbSuT0NJWtUFWcR4xWA
6x2c6+q5wXsHASiK0yRk6zvoO2ZC5O12uom7wmgnmMHaGamtAPcsOFnQx7xSUE3a
lFUPbK36kKDC/4y1/lRQBSYZreKNyHI4v/9AvBq/NiDa6kabB2GR4II0oEdYsxrn
AD8XxbsAYHxr1jqw2tLoyb2VqmgmCvS4DOW2WgvZ/YsyJJGL8TygxwwoDJOGMXuH
kdBA1kR/Cg/oWAX1R9gnHK4tVq5pcCIl6MjIhbty17AVIrTMweeEZC0v8RBuZz4g
ga1GmiVEhAoORnJcR88/W0WDlsgCyEYzWm8wpOKlVI6MzmRJ0R5D9+mchrM5qXCK
wO/gFv9fKLw6xh23bynEDLhkh2Q1lVg2ZaCsacuWlEwJzthsko0NCXf5QOIwZ8GH
3gQq0gLmd0XfZ+pI0+yx3Flm78KIs08w70JxAtSunDm98bGt2PkA7E6RBUcnhrHw
jIHi/0bxzFH7tbL4Xhy96F2Gw6X1OC9vVnARcuVT4Lji1g+2lWen/8pFmW0IpZ97
R0IL8P0+Wold4jqEiNs2ogmKZsu/HSkoS0tvusdtcoGrKf4BL9WiePQlS1fBPb/Q
WQiDjajCDIvn60Jid80FET6e0mqNgUGu4ZVQtNOdu9B8/2t+9j0AE8rcwYRwmhEK
DTJGSx6w7D4z273zr2n8yrV05Jxi16eLPLiQJsTeetcnlm6svRjscTabZsRAieXI
K4xHxoRmiJSP1Mgs2U5r1+oTa3PQDCgPJmARp08mMujfZjyVKjCZDREFXXsVysch
nIhgngc8gfBuR2Gs3UvHIRdzAw4I5jemVC3mNt1efC48mguA7JS1nNfgYBvVkMlL
GZKLHBbAg8X3Jdx94S7csHPiKKjS9FLB3Mh9rFrrDu0v4H8vVdninAJK6ONsjNM1
94fxxK/D8yakvNXXu+Fr36oXkvG+hH4S/NW2ocRacoZoAMEZQwyid3Dw/oTKTbpP
jSzZ7mvrXfWKY6HSdRi4ZKdfk6lveArhy6jXBn8KA8kyp0djs3xHv6nOQzR7k1AT
MH6IzB3ggboZKfx5L7bNOk6H+7e9r6Nni/f15pFra+hpnm4lmh2XW6SizN8Zvo6D
h3SNKTlVPdFx6g5VVY3RHXhZdSr2GXJg8TmCJKjv11ORHBo6KLt6hF0fPOPf6Q9u
Judytaz4+GBrHONdIE0KCGh4unoCRaJa1p/TSAMeg89WQxNwk5CcGv3E8Lz+l5xC
/GmMsGlThVJ8uW5Mah0ABCGRxNjDJ1F1RkdqNhrICq28Js2ycitV8HGPURE0TNs6
SlxFWICcq9F+ICboc1kQ5gN7+mZtUkIBXxKHESNIE3Wlb90Zg9F0l1ZBhso0KIJa
NJvVIuLOV6Z4X56RxEB5fDVs6frbPGtKFWSQKNNCnY3Q/ePjvmHlZ6Ukq+SwcaWU
Df8PJUfGjOk8/xQvR51FXlE7N4vfrXMv4cphXoKZ9BXVBUkRsCVK3Rw55OSDL2PU
T1XWfCprqpUy9Vq6H473EETnL0HbVj8yyJToVU2j3zvJKrBi2tAiz9+Bv+NDdAQM
weVvLFnE2aOpAHn1xQyHQ4CM649jFGkOCMaIqWUpos6qkIZsfRr0FSNzGeodo1ui
bcmRwJZknX6JZjyaV/wjdwyMv3nhtUVgi25LJ7wr6CUiSGpc5xIwAEI/1Wg/DEUp
cqT9dAnScf7xxUj8abSSf0inmaTHsrLChcCKteOMIVmVHBpNxotBkDHwhXOdEk+Z
9li4nVBdMmhP82BI2K5rH36+80Zuc6DweG0DHFq6ieiALrgqOK5sa0QzHwjihsU5
uO4HPLPgOC2K2vTf3tUSca3STnKH054Gz5OHiTPgyLHoLIaBcZw2TpXJqmixhBCC
EsuRrVxF9KiXNfLTuM5289E7RZOqPKQWGX6cLJT/4RdL1J9osejL34ho0EqaS/ew
0E+VrlpQ7Uzi9e8TNS5Di6hW5BJ1DD/CNkhwXcn7jvlqw9MfztpJAFx7eYjANaqW
/mrz72QcKSHKfxeKbnwXPOCPSE/K8wyCQizFWxHnjpi6ePAuIagUcW5cfffV3FAx
U1WH6+4qsxsxuSlXvHzRxsNsKQNboR4v+wF9iVEyDv4FeAxSwLJl7g9KYdvGnDOQ
EeCx3yJbnkRrOMmufsIF16sbEO08C270UOFTIlsbGC5Oon8ojnSmczLTUTeAQaAt
IyEWWXN6skvJnCD6JJqyfYYf2sYjU1+8oSOkcaTtTqGV/zp7VMaJOkbTZTj23ZUf
RjBvKhjhajI7NnD8XzteH5STwVNfaQx80tf+LgMY4ZNv9lgzvuZMG7k44XzV9cOB
ZdESb0OejSPvoqsYP4UQBH7+zmr6UYV/3TCWqnw+4jjZZEsS6s54LnWIBlpnLwoP
S4Gt9DDzIQ7SlzLBALyPXqBVaWUU4DNYz+lyDt87VvyoX6k7ZPrGZT2b+EU/guga
QHtwt5PoaJ4kJSuSY71L9GpWXbc1IEmE9I1jXQdCCjX1hW2iSXgLgMf24NmqV8tL
qMsW+/A5iz7iIYzBTbwWlvLtRn51Qin6Si4ywt5HqauX3KGBYC6RygSwrhl5/PIz
pGQcZG5bmvGm7nSDKB+RQcYERTsbFp3+Ib+wF1ovbwbqqsVwp3L7UfeXEXaY9IqX
03pLdfIH47438TZb8EgOakIEYX8mH5eE7SeBVxKgryrwdDtAlhoZmkbkzcN9wqvs
uMn6T/lMp0ZTH1xiijHegGw9atlMrBc+70NDGWRV5mqp5u5QIFSaUChdO65zNqee
PoPvDOdbZ9Ldl0uI5rj5kyoeaPtkVUXaEGK2e5L2VAzc4kVZQgoxROfEH/38+lbs
lDjRoJqny3ZCX1s1djKgeG2VadHekEWgL1Pv1IhL+uUy3Wg6cmKUWAJA801vtLgp
tEAme2P2cKTsE2258ER4yxjMn/KQ0gRNxy4lQtKRmYH7s3Y2UAhd6NvhkBAu35JA
H3hQtGFM2/QQQuSSphd97s71gwikovXZN4trbK3IiktetIklmnbOhfvXUARSXn86
yRGcMIvpTdSYZ08hPPr55cI6ZrtmTXdUlLL9dN/pBxNG0xciPIrr/Yi1BrwuKcL4
ItnTMaf0tzVi0bY71I1mMTk8WXLHcR6CeQvVyPy3f+de48VUQTG0iRfRnG1t2K/k
PtQHTiLbLP1HHgs1XA5Z3zwTaDnHPXwimN2KLPqw9KAFHWp3gFRx+3fOnp3Cp/eZ
MhvtkGJkPoVi9JpKgQabnSi6P8d5i3FHCeVspgqn0CcBy4lG/aejLQ0+KuqXlEzT
5iE4NcCkHxP3DXpxGzMPlnCaA3lXy5idzTpy2Zk614AhNq534ipK8ImTDCXwPT66
jltLUWESCF8JIR6uYNsA4eKYfDyCxkDBez1hAA/XfUuPnz8Rj0r5zL5+fxsbhH/m
dhVddOZK+M899O81E4T3S+NoxBBKf9eQ9f7Zjgq3+5aWzafaaUeoRbaXPYqG1PGd
YL/vbJ8ikubAqjsccAxMZbX66je6URtoQtJ3pIqt109qThiH1M2qHq2GhNKTp+4F
tLmq01uFmZ7pUb8pcSzSju8vnFi92VvxZh3cWN+NAeymhKNZlX+R7+JvkofM4vNk
hpJvdo3YquD3NgOLZJjp3Xj7w/xSSxKoL+iJImkj5wv3hPFFCploZZc5M9dXH4ws
Dt4bJeVuUR2fknziYg/glU2JI1/LtuY1wCLHCrwtvmzswIGxsIGgEzE/h1DFWP7c
VwpuGtHq60WB4bISmcPPHg1rpJrHyEXgWWqbo60j6VRsFcdooTGk4Y9/yBACoOEh
AI91DLlMmxrIMAgodZXVyDH/IYTm+XmK9I9v5+/FuqDJAXFzmGrHUht1xNE+Gw57
8FIvpqlySRflKTaEjgLvnnfN/WZCLLqm5I0GI9qqkJnxv1s7YRHA+qtYLe7vMfgp
9HHcya39khO1anBcghiLhXiFZ0tO2yWdhPEcrzoMrwgaH80SLNKkXeqKmxp0Z9uI
DGR2xSEqKNiDhD7379VAzWRAl86K6CnuCQc7uLNb02CyQ6xFkBR2XAWLJNN9aEmW
3ik48Y6tUmUa2EHDQwo3Sgut+aBxIAlfhlbtDLjiW0IPFHDxTvLD/aofCKBReUdy
LxEXEt7WBkX+MZXS+wt/22GksfNG1SeiEubvmANgT0gUYUTKV6ZTAzcr8gs26rVc
16RUPYmCoI+0xpX+W99sc9OIIl6qe1HK80HBvVaHd6Zlq/V1nweTVN0y3A/a0Xgj
7BeBy4UxLb2EYo9vhUJ3Z5aqMchq/eVVJbuNAiRA1qm+MYCirfgXZdCit8mJNnXW
AmMinfFwgQ25PoeDADvCtmROvC8ELAmxP1xIAd+BlbN4C2hjAHBp4oguGGmlFmqf
RkLyrkftc0zPOPozcvczYt/FbNv2L68EWkOs7DGiFwfq37pCZjOKmy2W4zrDNChQ
tIbU7pN+c9OX7FzRtbT/Xp0W0R9AOr8P5ng04GQH5EvsKPVnN6UXiQEYJWHl6w9Q
1XsIzbG5p+yG3bBCMvXHB9lHyfuADYgdke+XfcLDuESTzfFRxPazQnHTkGISc/tE
8DBZuwHOP7ujTMjWXiH7MNnVMaopzA9Z/Se7xPV3CYZ2m9FJupxuv9stesGtKMcU
pxpbHsxmrGOoVJzO0h2Gn/Kk6T7uH9pj0OuywuGQMSLd/m7dTdxkHQhCJNJoWj61
YHm1MhtfqFceLBaQ7BEMwuqkbv+TeFLhABcpil+Nwws/KniFZ610s7LphrrzTWrM
s61zKC/yd8OCe0J8jRJRwOTkLwwomli8l5PGK8dSJsyJgA5Usw96LBQHPTpl80rr
aSaWq6erPC6U7rfQRT6hj4eM8OIdf4rt8e4JYQDJ1sPTjd132uUCPGWKzqt6HNhj
Nc9eluL9Jw5u+2GHeHT+xXHsQwtSQhrqYONAcg/L94X7yuVY4iDL1vEelTVZgOJP
MEew98Jl/81CAX37J3L/mtsqtf40wwqCIeXxPIMuiNJXRFQXIYIksH699IIgnW0N
r2RhsdMvmOeKtzrE9zg058OOhCTuvfzGl9OGT2kMzv1UiBe2N1ofRPU6zthtBXiB
UN1dSKCpZ5Frr9Qez7bFF75Y7sr78qVwrzXAqo62kFcHoNWJiW4F/9NYpRzD90r0
ttICVnYijTi8Dc0DsHvqAf96ccx8owptC3IB1Ep9HEvYnCjlA5tGceau0VOrdgJu
J34fYBdYN8foAAf6mVsA8XOYia+R8gOY97bo2qKyikpi3I4AExFLLJlwDsORVDdS
66jcaogEowZXR6Y40UIgbjiReySryKW7H6N2AMT7sAl7LUgctGuw73Qo5lqCtdAL
lmx4KtQ2mQ+xKVe2wGNy/XC4dSPYUgjjoOFh0M7aLpGg0AfywRQzJeWFhYcuH1hH
W07zJSmVmQcNX4VBJUY/rZUmp9DncLNHnGV0sHSEViqpAphG/b42dPGGfE89nOrU
4uB6ISRajMjpLXLgBGZqcgqtzgzOH+sSNhXlaZISkGxt4YToJEUwRCM2ltnL7Lvd
Dq4ttumtselOa+1p0izbL4bIHpGJY3eGWfqUCxanGzvQnmyDfRKOIZP4e/lmt8Hi
SQtnm++742tGYL8gu/ZBeBqHdiQovFBiLsnAnvkLZil5jwqR2G5/yBIO765wcWGB
VwD9X19QkL9aQbKE9ZwPNZweWELVFtqO0RDJ0RES/ZXvWGmLujg7a8BBOo/pJ/7H
4P9wEgG6m1bzZE+rJ2CCe00JT8EgK7gntXdtDurGkiM1cW1XqHGKVgM8mUGaeCNo
ED077Y2egn1k/9/emO2t7SPIqg4mOx0KgPh9Gfkdl5mo/XE6HkA3WiuOBFSBm1v9
ytNn+vn/WF4loq3yRXrcPK6z9yNkZ7EEEcJ6YnSLQw6zYvMfYUGQBLshLhGiXKzY
3MQp9Ftr3I9w2jTBVhdm7qVDQFObqoxL0MN9zxOQJS9mtJBK9LV8LHe+YiRqDtAw
PTChq6AySVxy2muG9jNPJSSZ8esmmP0ugh7//BGnbLMjETD+KLmAkNfUjzlxh8tf
F0gu2kS5kl4i+HubDHiw/dz9IdQ/rADrVQ0pPyy8MADRbyXE54i3cUyvN4HVv/jz
PXKWnlY9VdyZkJuZI24wfTaPTe/DUw55cAqMGyGZN0OweRlD9sGcwLW4jtDoCJto
fQztof1RjW/Oe5dOeiO54ltUr8Vo/rbPxtaAIJFZR8MULGU7yHAUwNjE6xldvsLo
p94J0x+7KuUrmYjSSWGw+MfNtz9JF0cupHBG7XTwLrwsqcealOpo4n5riklcB2Xc
YD06cTzm6YHHmDq/YJ7D4dkv5pE8aZJxQMDOBCOFccvRsp6FlzxX7RsEN68U8rl+
86HjKjiTAhbq7zzhWqX+yozhYHATZ1ysEBW2W8EOmY/neYthby8CLAyE+gN5RalM
OeV+BBqABXecMisgPKOELBhkteMhqlQsbclmv2KTnN/E9pRPyv0DVmgvAqGdqUNk
EiQ84s4+3lEBg2iKb4p5+rvfG1o26/OCzRvll0qLXVzL3Ul4EqWap7jW6RIEMJQJ
VTKstL/X9IrRmxpWU3MmlksIGbrINOPEmXTk4eHpBby3fp/eRDuiFeDT2tQMoyTm
9KvVA6aMolAgiuyfOH/Yq1B3nuHJVQ5tLnmqHyUBCYjGgLJB3n9XrGbXo2sk7hit
xQ/pd1BQcAa+6mTHGKHom+5yeE+UJv0ANUvhlDawcv3s3s6KWKkTCqroyb+h6r/Q
6fVs12vRF1bqRNsfoXIYQdGNKyWfRYMy6PZv+NW996rMY1WuLT3PzAozpCWQasd5
nsBvSSrTJ9C2ZuX7D+pTm9gSel6yml4Oc2Hr5gHY8qdQPhfb48chPfzNYk0czJtr
bzs8x8m/DbxZBzx4iF1LLCAY7XxP+PSdncgkmFmhuELidLYrt5HR41exFQZyfpuN
LujDbl/Z/c332o6eRopGMNRYGzecexklDrkuMO63b28CpewlE21XnTKsEsy7h8NV
ciRzNB94SZzme5IaLvjYxsnvVSHWC+9si5pBDb2lxeVgs6717t6FtiKcoJJ/MwsV
kr5MAkyQpRqIkvx1x6Ayf1kqpyOTckaaScVu2foY/Q+zA4eKZSMlYrjl4JRTBTaW
Mps5w2FxR65SW2cVOIKFlh8RVq0btABMdRYUmj/cQpvOjnI/1zSw532Wlu/Sy6fz
vDGBB3QU+K7GmLmmaW0kbQCFfFYjQlpUOeD8ccsarC0oJBH3O1Kv+H5hJ15KyM5j
wrRPPcn3yPOoyOO/nybesEbM91rIoZJDFIqaHQN0JJrExbgOQY6GsQSCmFAek1i0
L8kqdXPjMVuCe4rrcq2wdbgyNJABMWWB2Az/nEDjpoH1soGdznOJdPu8JXjEkNZe
ZEJh10mtavUFxd2sS2K06OzoTVH/LqsFJpj97gDfz6zoRzJsIbJAfbawYtI29zoH
AEJoAlhRLIS93FdAiToFrg/acWPY8is/B60iDX3qC6uYZ6cmIg36XyRGBY18RT9Y
iawrvVL5HtNwGGGFj2xGx04a8W5Y9dpPkTxt3mr9xoR+jSpRG9AatLd2pramC0VW
sGbelYJfM6BoBAtnAOmDaFKOTBRbMhiGN2uEhssr8tMI/gj1KTCuhnT0v1T/wYOd
iEt29s4icRZik+ffdV6hw21qFLp/vM83oXwQ8EUGVEuxKcLavCszCDLErbCtXfFH
uMHgggSVvCl2FVousVb1NcA4B7YZ7OK5cs6xGB6Y34ALS9yXEOyJyHflAVu0TaKk
ZzrTpifpgz1Nt/kpe8ksBWhlzkytHxYUqU71u+AMbuSlq5jx4JmQvhgxzIb5j5Bo
szOYHOd3Fc8Xj6H+uVv4eNPLsoJHxLJ1KMg1ijhp33rrL9A75W85KujeWGwJUlOy
LLxxIBsJFOtznkUDKYCbp45QeCCuaaC2N35sUeAi2cudyzc8YYgwZoOonOLstKbg
9VI75UWRlt4MqvhRrdFviuHvmq/fxeYdjYH42sXiUc9mZEw40g7pIGB5rqrA0CDb
cQZciQJ4ekddBGgY/g4ZBONeIzYmienNTWI11FZL95Dz4U2PUuqCel1lv+bh0cws
x04mwayeOpsQxJ5ZDfBgHUTytGlkc4jGZ0eelPf+Ti0F5K3+45lmTjJ9A31aloYo
S/PmZquHA7e4qTiedPoNAUTx3yZkIrA3Gif5sH7RE8Ezj4eGfsrmxwdB9JfdKE3y
VSVn1ANya4kQxe+kkTQi3vpKMpZWYYw0RKwrUzWgBHGTl/Hp7qcmB4py0IxXLUn4
GAn940Bk5AT6ZW9rhXuOYQ+qEnW86fGnnGDS+jsjgpli+FQE1L8hi8u+EuNBkwuO
dQPnQT/eAffhLPgAqoJsHU6hWgHq986UN5PyWAIRT8hi4AlCa9p/dI/xzeaUWwyg
ioucwiFRuHpKx40TcI1ozBXHC5KTyCmAxuKOcG0wK/gUurKtf1jsBnsAyk2xe0QT
3bnwajTLy6WrJQC7vFw36SWM23GQXLMHA4BQExcwnDdqLIskjVLNX8QBOoyQhEVS
6tCg4Tg1qQ5GOzX9m9XPqZG3KZ/skgGiZZw8RBd2qGRmhjG1imUJD6WjACfkeA8j
6DbS12qywqB9oUpctH7lLo6SptMwPh7xsJzjsh3fPLJ9SDL+V/17BB+oa9ZZQVkt
81t9p+4TwGJ4+Fj1JuWwakLQ0k44rTVdKX+IFu1v6jh+camOEUAq98I4OhOUnrC6
OcLaJhM0t1hXuze7GZ/4qcgfJGg2+3UYRhDbWgOXQV3FLraMvgW2Pc1RERCJNO5i
aFtDTA5Vy2kw0HPxMKi/YtS1IWFA1aP4ucZUjiYwlHlYyTr0dSerBBDovYNy4Bmj
50KsX8xXcTWO7foa7CY52E6jIx5TY0fExOWTkeOMB4Z1pCpgXuJvsicdM7UaZEsM
DXTydk1hNyw13zYYeFRCUIhsZ1o8/p/TW+kDtVrthscys2lFFCpvHVPWZ6RxAIHn
Ib0JSDKIbJum3WarxXaR9EINEAyp08FOZbRoOpVkfZRjeEak5tZwC3ktqG/v1fWb
/Btwi0INA0kC1oB/mVWqPYZ3IWMze9U7M3E8zb5DIeo0SV+ZZ/xzmaZ9dNgBrWoW
EyJOs36a2VhMEd4r4q/53TQwhia1GpB3g2iB8ZQG8UyzuViT08uWWoXFFIybFX76
j6k71Iu0eDEMe+YtYy0jdTEX4mfVfwh/VW7Ijfg0Pq/nzIozhZeur+mk8+lRy8JK
aWYKDuyYmXLIija42c6Dap5LIhjfBVwF3s/DOTokyr29Qlu2sy0tQwlvACC4v9nv
mNkSeNZOi5c9xqfIklMXbc+WOVU0lHnMZNmT6EXKJUzz7PCIfll/MfxJH1hS1XIk
uz7aS+Crz9n6R5p615yPw0pZxAcd9GuTOqzjU00LHt5Z5PvFeJEMy6+RD20Uq7YT
y6Pdj2B5LDmy0bWZBXUEizeIH+Hp6UvsjHvZQZXqujJipq9oyRTEMRVz22WKkfDy
ZW6Y16YAqxJgrgzBoHrRezFNO6bpuAn7AMqV5KwBjV2V51o6oLsBZJfcGsFs05J0
278RPM5VZF06bJT0/JJKb/3IsGH9XRv5KfkPQacVdwezZS6sdpvdsSH8eXvuyiLU
fdJAnX9pezC3PCE2GqLZWBI0rZ8dvhn9WnTDWkq34mTMBZcgDqU66/oD4g8I4Mjw
8XvC/pSethCtNyagWarYFKEn1NS2/gYJLhxJfVOJyvleppdw0dBL5/U+O0ozH9Rd
QT0ErbYvIDnrkpFkwfm5IuP3sdk3scCwWHI2clqGYZJXA1bg25tl5ii2+NX2L0d6
Lw6l6eNWslyLudaiQ+MaWh5hkpHOWFcqrJTdWTOBL1yKr5JyX/AyK+8voAFPOtWu
Lk15jHVyzNcLOtF5B9xhEWKVjLz49qwCBwoplNGL+sAAImAtf6R2TiJrqaySXzXu
DqNZvhOD+SUcGCvLMCjoA9NYS9NqYgihZ+YAf5Y1mqEgUenui/TSO2+EUyJnj5Rz
5yJtKTeWZ0bncXQfzYWfQ+miWN0jmgAO1QuRO5lvJBMiqGbDHlTizz0NzSJe54j6
XBSSX0z420WvK7TiFzI1YZJZG0qj5kVA0BVqLhFBdHIT0PaiwXLObRnsVWU9mIRU
wfHbfY6guCMG/pnFt7TxzbKqKYXvssjbk8vgbQxCz0XD0DJ6OohiNjnpbyYZwv59
mZZP6SVqqMl7dK+jfmOQ4b4RHXNqiWxc7BVd/2h7nSRqk9X8J6GmvdUolJY/v27v
IKRKxyreCJ801Blpipuc2CVJs7wmZRCPDa7F+RSFLQuthwxCg6qdvat7OpxtRaNx
I1ek1maHdFyGUyfbAnNga0zmCvXiBV0LyKhsOEkn5gpsxHttclfrLwm3dM1OxKvB
27GZntGnfNaufMvpD+HN4iwtXtr1iSbwbHlzPO9cVQELPGklElKo5uDKxl9LPgbV
FOS4H3y7BLrBJ5WDexHffWQ0nlvdICD6eD5V+Y6iOLmrfsFSfIKV2nwda0daNVGT
YuLVTR+TIEbwGWSgE4pwOtp3zkvYri/KluoIJrFRFQ7KkKiVCJC7SCnG5uGwPv4J
XHiI5JAf+lKWpMWvBgjmSZcfxgB0AraQniGbjdnRbWyU4dWZ1cEsj51dAb2dDqIN
tEHNgCivLZw6++r/xDHMAnTh6ZJP7+Qnfp5ohACKDbdAV06hM78JMxRZmYVoj8be
U5XWVGT/PTMB9wtHB3a8tRE0rdDuLdWm2vuVbo+KuBBR0EYkb4E4cv4FRRKCGvoY
XfFkTQ6yeRbx2FblawZDT0pyWDONw9tfQ+Ws5EdydrqqnxeHeWXUtKIw2AVRFSna
NUdVV4TtysRVSJ8lceLBNr8m/G/C8DmeOjmmEFrI0dPJDvMY7fTz/F/lkOJH5UVO
q1ba4t6qpxgEG8W+ppcWBKEt/1UNP0FC27Lbbn3ALIrl5gb+aw+jA6frH4z+4AfS
VQhY2U9svOEibS6zcdedfYNnuqK+0hrU0apEVn6Z6rQt8t4S4O+y23ci+lDPutue
wJo2ypLPBKoOMZHGfdbbV3gOzBnvrcp4RLjMzAYMG1Oke718dc/bGe/Jj/aGBE9L
dKhcYMxJUQHD9NMnLiercv+VHIJ7sLVoBQI/GxxjCvxoJOcPdXC4CEt1oTjf8dpL
cYrlIW3qt9alRQtNDtTsBwc5nLBtypZaJId95MEVC/AMli24OU1GGVDMFmJm+qBq
ahrMJYD8e++ccJg1P3a97Vq5tM5J4fmsLDHUMargfJFaYo1YS9wOzyIuw1RYABxX
01G09pi1/gUBJ1OtiicwsnDP+3R4y+tg+I/GAJmRY/1exWdK+ny4EFvyXi9xI6bZ
VdRaj2wQNn1k13gQufpt1C/lIkyihzkLrWEHeNK0Y/s9i9SfOWTCA+5okOZc2LC+
XjIKAK/Qiwi1Chdkc38rd+WDMe75s5aTvLNBo4dlTQN10uVLnj2kEMZ2tn9kZn3x
oLbHYWtjPzTPbI8gO9BjzqrW7FmBcnfVeOswBzkBqDLUVwoJpGf41P9ika/z/H1u
Si2C5AyitiTLmrzo1WeYAPDch/O4l7Ndc4XLUlTICflqHB9u4mh6WU44W0o7AwOy
m4WbCgT1uFzVRHU4wwWyPjE8asRMdUAK/14InTuLf7Z77k6kgKkxliyfoa2+hHVH
GCFSdIHme/9d9CCDQ8aod3FMBGdI0zYf9AnmBJQ8S6flbT150HdOQdmW1oizxhB3
4Gi94+rwv9wH9nWl6O4lWKOrILoRKNltAafVULNzYrJzoMiiM7qWF8QYIK3SUCl1
k0Iu7rW7bevc40DN/Tw+zK6wrz0dLaojYVwtSM258zO3zAAPDf1hczAPrl+GZRa/
hCdxb+uLtJfk2Rlu5PwTtjKQ+tZ36ed8haaPZddG7cszK40xginpnGJmzWqV/U0y
VII+0/1gOXVsQvDqlb2cPQ==
`protect END_PROTECTED
