`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8igwLH92g4bh/1fjMSWKSfKCw63dklaTfQ4y6OOyF7tIOwS4QexSElt60XgqTSed
YniHn0x4D0DbJ39dzIXsvAiAp0bk6t/+ktCBFnnRDRywYF5eWJr4lyWR8uNW/CaY
AQUS433YrBmG/ZP2mZ9joKxd1MQO1hJM6PHIgsgulL8kYy13fwiybtwWrJ3JCDyE
OiBSKHPVMaIfQbV/ibKwSxfPOSxPix+dgPmuU8ylmiq9C2shZ9C2zyu2Fe5hdkG1
87qMePYWew4ohYOeqtpAa8CXEk8OFkCL59VftLV36ryvOmGTBtp2M+2aeNJyB/Of
KNR9UOFQb0/lr4/NH3EPeWY+JP/xPSmLIval+PB6wIEsWLLdNLlaITxfxWxPEucz
ofmAiGYVUTyh92p5rMVGuOC7R8iy/IezZsgAQwJEFDE0uHlShO4g/fMyg0rux9xJ
HjNpe5mVvrjLdnl53t4vVs1SzlkInbgCUVTfsHQ8fRht9g2lkDNdU+XaQqSpooAX
VVH1uJx6GB9g6DK6V9371NXnhs6E0GN+ULdyT64mWTyIcOW6xCEpZ5jtsDLLiizR
Ihfw+PI5B8pQeHTJYlHGpfniKu2inQ4PPMX3bZ2LBEvRdWUDKR8WdEiSAfuuZiCt
OujNtN5iV7hfzuGq8ONWBQcnK/4TJELkAwzz78LaxTDVa/dNU17lNyiq6+AjsAEj
XGWIhDnsA7DfSfiDkf4odktoknA5GC29GuS21juFrTUvxxUTrlSK8/uG9Z1WULrY
6wjRcnnO97OAFDxDg407mblAORkunENhZD8rd59OsCK9F1PdFtPo61Ol6hAU4wBi
8DY+5PSkkvUVeggTw9m0OHgjcYc11YEnRtjAsY6/7L8mLPGKHpzoJEaJBLzSSOdi
l4gUd7FLawvBFPgKey9YNTGgW7NPQNL2CxDmPnSUXjCtVXUMnmYheQ0ZYFZOOixp
l8krgJG07Bhuili4fMHckPU2jf4lkxaLOaGSh8y5elQLZ3Xx0Njy2TMRnp26p7fT
xzu0FSZqocHyNK5xz+/L3HLoYIbUD8DL3bqKNv3xSWpV60Zt/Va4fxz/xkgAM3Rs
5PGZJZIsQLEkBM+QgOjtTk4GplnAWFjI+FhbFWzB6kAifw1LQPT0YFVki+tkZs0l
JPIliVKgTSeL3AoAXH5UfSxgXkgI4ff4juu/DMgtIzrhFTMyFp4weUint8jVYpEH
oGXEH6wX9qEX5pMTRimyCUIo6NwNJLOqTyY/6XW6yzDL9DSGeRr1BJf8jYufACwY
D+BWQh1h8lW2M4ORZ9fCHozNqxNT56f/gDdd4mIdKBdB44XX6nv9p4sVsdKyBE0v
YRVunc9WVQw+UU6MhJiom/+58vJUT5Weaf/q97M56A0XrDwkGVin7CuMSS1+9Mka
rK6V06xycYoo0zY6LbM5dPhl0TIvQPOclN3GV1CFR+XLw7PK0/ynRbgLwAg5ROLJ
c8SlGBbbWB4uzJJ5O8rxQre3Hb5Z2rMX10aI0i3wJXnKumetmIJhB20Bm4V9cfmM
TXKZgOurIfBFcpozgnBl6pUWTkBNiAJ92W5MWQN9xdn+ekDo0qYR/qPP3wxLD0VD
qWaWHsz3KwWWvqXyNmpASjRT3pzysegwG0nOUFo4lNTVxoz9zdWUsD6NhLaCabnX
bAQuToDCrf6cJVUS4xZN2oa+aSNUqyL59ibT1hk3YG+ekjq+80Nx4wixMraU7lol
O0TONMJSb1KlgOLIEqYN0wGGmAMRlFh67C0vG6RSaLPWLvQ3Rtp01IRB19MiHqY6
ZNgm/7uC9LFFe1Db4+tshTXVd0rxrFytoBuH+JyRxd0/LQTJf0lb7JkxPspSrR1U
1+R+JIGKndsSuuMK6mhvII+COjsCfmBdUUNIxPFTlksb3SIUqnaRzSJR3S57gdVx
8JGgQjATExiDQHGQOya8hlGi1LC1SCAsy65S8Ru0S98Lr+YnkR37XTqrhYjFsZjt
ABD6uPpQi2DYK8aioHmEY11j07wxgvQCMmGnI9q3wLMLKcwbWMRf5/sSysYpVcW6
U8EksdBUyAXOnllObb+3VV0Hw32DKT79ak3H0BA+2Krxkul0UCs4zfpIveaAtQnp
RTYQXRyX/Khz4jGOvb1hCHlcRXmkos3rEzCNrrMjEOshpSVgnbYEV6De8ZqZj43R
nxLEBct3LO0lYb7rTMH5JzYQ9Dz+bhjqV6j6nLc6tsIXFu6GTkTPjq83urty/799
LHuGniOlPq4BOWXVJZwOFLGVYOuP7T2+1whjYr1Kk27uQdHWKyK0LnHG96RgUNKL
pP7nx4HQ8qjRJZ9wcoI3lWFPAoJIrY3USrKs/1Tkh2KlNM3GBJxIPIIARnepwGnK
KcuSuoysXWeEDvqSl1SotlRFQewmfUrSvlQe7N/WL5vr7ygNEm2ShMkDw7vp6tcx
ODNA4GtxoVwkD/6+7ASgBpJYb0bY1wqsIFMHEhM990sdowemZ20vr5BZ+At8ubea
FcZ6INi/kgkV4FGk8uzoeKRCo7SATZ9Ns/YbEY3a14XNi3YVhKPruT/YwELDwEVY
dTB2qe4fYhoPC8ZMWat8HtJMg1UQ1ftXQxoxibTaYHRKo01vqvhAEJhZZMAYbExq
jLSvvwLS1b11d1b0d8y0H1FTk6HssUbzncA0/OeyVt47suNRy7uAHl74w0rUnnHp
c5700ZtfhF3dJMInCM4Tub4E6+o9wRMd6QiaLh6CxYBo0sA3e40BJhu5mD1hIh8c
WiFIByIxSxjDKDqxMVJSJ6nmVu04J7giOG4yb0C+OJnLAWlH4WZ8RSpBSva6RfU+
mcgMzpPGmkAAFTv9PSBfCHKK1FvGvpCVqfoGMHOi8oViWxTHYLcQSnFXK7nzcWGe
ZRhIupRJ9iQxv2KlQmQofOej6+W3y20gvFnfmF34Sdtri/01R7zcw1Qd5cULXrkc
UYEGMoIecSEGDN3+6bnk7kLxp9VxOZYyFrrxxV67UXjVSMPvcXrh4jCam51gVfO3
6/QgFsFQh3N5k0IU5RqO6qw1Qx/i32gDczZ78+UZHZ9+If2lyOoL6KFKrPFXb2Gg
xJUSEWQ60u4YQ/NBvCxAoOpqf0QiLFtCpJMH3DCQeHMHdNyo5Cwlb4ewy10cjWQq
JP9qxZDweg0k21fXkFF0rePOrwlqkDZvXGbuyXxE7syBS1rcXARj1Vk6/T3jyXer
6loOxng+twL1ro8cnxJAHk+nC+ukh56MWzoSh/1N8/FIcpsgvpxaMfApWVLTRA59
YcBO6eFdXAsdcVaPuHGxwcPF+onC1XAbqSW/hIEYld5W1upbHYa8mtRTIbWD0n/d
TAWSbCOInj4HkQhQQn2Xpzrrf6h6was41VI+BhGAq16qdepZfaxUGN8U9MkzJA5p
9X8hlml9B+QjTICudbBpBgKUP+DTFLfkn0hT5vLIcOwceXEIOoLYGoKzJWqdombc
kYx07vvWRlCaH7wKmIKCItGE2cHXeGirLBrYf22JN4kJc/Lz3oYlfJBU0vm3ezSD
ORy7Ad53FLNMvY/LtOwnOBjgDBhjDcI5YEOaHTM1i3aqN+NxuD4QT4z8n2x7nsRY
zFBsWyCziVZoTXEaFf4GWYtjqlwUQin+PnVqNlUEPK3Cg1ele+oGNEhgjuVseDFM
tOEO8T2Vrj6+5zB1QtRqULy3dLmydoCwIi12KVGGcno54NFi9b6HKqE9TqMN3eL8
zDG1CykaOct6gz47L9hlwTLM4hih6UJUZDcCVlpfOSx6QmbJC5NcPWW1BMzOKv4C
eHZ0DmtMx0BXmW61f5kCkYIrML3zCdsd3M+6/xELk/K1GT0gfQM/zbe3WOkZjPr9
WT3aNATas+f+fGyGzRIVqc1lLZEhsyCq417IP0r9QksE9SShy9L9FFuCG4F1gPvQ
WboZWcSQw/ZwSO7r2wlTvsiAlMyCuGCQ5sp3tbLxEShnjSTljOtLf60pUQCw3PS7
dl3hjCvEv3+49ZCu2YT0EslSnYJNZO1cj7JAFQqkWxjpW1jZPSDTZjdf6nvJIATx
/qEmFUoTnUBRdI4ujwmv0xf5AhLSdvlneuStlnCH0mvtvcWRSwd5DsEo13dmu837
k9o4TBlIdxI8TRV0jezXB4ivrXN1GZfsr+3FA8I0i7fakTvVXMKP/pmcpC/hOFo7
+6v+hYtvgqa1eU2asRAkGAEry2O6C90/tKiiinyX6zKVeNUH01AUP1fCtkX0xaPQ
jzW3reoYG93giZacVNJ9jhmS7MQPd/eoX1RX2bDT2d8eh7BfNyzEfbIxFx67820e
UYDRS5fQ4/T2ou7LobAJxy5phL0FLX/zSKrdwYMgDWTRNQhynJ4aKnWdwh8to4oy
dlk3TbBv0JfscPNWDYRS4LDHyzVSdS1ImZ5EQKXFW1GzQXJjvIEVP/dfbim7PcxL
m9GwQWA6ffEn6mYH71lgfr8J4l/DIaStiXkoPbKzyR7IB/Ou0NjyD/XFNW0WmNRA
xtNNiE7Mq+0NDyaA0QwS/pMT6NwcxWR5L24DCpUaIJiQFrCahnUyUYI8cz+O+M/b
xM+kCxgZglag83TfNI61Tmvl4pNKIE3Q5v1BcR1xsCUXEZxvAdd/cYIXfQGgswBL
9yUkbvnbPPWir7JqhuBWct0sdy+509U0DTVsuQc9NabnXdTjQH+t/KHRPqG58Ud/
Lj+GEjHJjI6Bs+2c/a7XIKKGvT3h0Jsl3DMwRH5lwQB3PAAYYlb/Y6q2TMmoRDfr
9oogIUQps+cJ7K8CTJnz6Yonxz91M2qehdWz9v9j5ZN4l4hAFylIOVn4NLqtMJQw
oqBlHLoAPWaD6k42wBSvyN6K/1i278Pyb9IIvsgtqRnqM2CfG5t0d51F1oz/8kMa
5SWlHmrSq+6E/YqrAd/9xNBj63Ggn5b0ZXX1nuCk2SGaIt6w/9X1YnVdTIT+IBlO
VdFS7PG9NnD9ivvyfJvQsTGIAdxu7xrIolpnN1Ymk9fH3q5z2job54tSpNwDhMEv
8aPMvRLdON//W/KOWK0oF9ahr4GS9UJ+GafEVlAgcI0D48emsmqkaAieFeLoqdfk
J4O5fDj2SfL0wKv8k6jJ1AUKbLuUkO6EmVn8YhshvNMITrUSbG7baiJR4fXBbLnJ
08gPMr5p9kTuLRXVdFHPfb9R/oSJ+/ujRzcHPluwY8+rks/9BFFtfSK9zxwIOraz
R4K5EWm69SvlNTNTaVF75AmYQ9wa16MiAzYE+td3IMGyYiUVqiw07ShkMiE297F+
1bJrMHNc7ycf/MEPbACQVLr5dnWDJh0+5LmMZIDtt12/qehT39yiQly/Is3L34wN
KUFgk0t9/g+IuwqRWf9e6ZQzHbIbxkOuOe7YImg0VwiAEbTQfLo1ECQi233WQXzA
YtJMI9m3kuQ5bDDxLL/DVYv2IH+/42diZXAnBdz34ivyMDTbn+ewnmF5bg6mIpeU
t19RVSxPsYohQguDU1G5268Cm0XXUHEYQhMwkRsux4y8JYQ60Q3eViog9xkprcEN
XphdYxcVKuJ5UyOBzy2O/g1LxZPgmC0oyqVv/eau65ySt1ig2kLkYjHYshkHn8m9
PORx0MuyD+9JpNP/b4+jCkoJaEGKpC/RxWsrS9NzMVXpRB+mGxbrJoiOyOdHwPGr
mpzL/KNVE1hPBu/RrZssb1+/NqlMOlIH6tCfXMnYurmMHw9x8yHN4a034z0L07BZ
cpheqxSWehBRD0A/ipR6AI5cClF0hOQbRlFXtDQo9XyJs4/yl2MIgJ486/qzvwmK
DYRvF63h/4+9DF76FN4kAl+/FUQdocHXvYIznQTsBw1evnuv+R/iF7wYt4fhlCbQ
5MBzc5Ca7HG0RBREkzsGUQeAaSrEbDs5vD+ttTZdpPqwDBw6Y0FBkGkLbsvIDadR
K6RHpgrkXPLkGTpXc32WYjBYrCn5Iodv7YHFGlbm0CHF7q2qD/HNwfaKNCoQD+RG
oh40Jkmf3z6rMtm2QLSzcImmz9a2Cv0HIg8sQJN3daJQL6SsjT7VAWV8yiAKuQjg
1iiRIklm+VP4chaLU5LYE0ERIG/roH3IXEU586+QnLSfpAsGajCEfpfJi/NMl8kQ
KsNI2K/VX1f5wKcAUUdGEFrJg1YmkYYMP9cDd//5VXAg2bbdYj+ghwFN3qx6OMKw
EOrPBeNM0U1Hl7WngIfkcgupo6rJDjl+K3HEoI94FwZy+spYy3rzRdqKCDgy4rXh
8a4Iwrb3k8giIw0ZrWk+UXj1NKFTtzj+MEKbgVHkOPJkRHet4E1DsTViSg4rjIMg
xB4WeKqsCC4lrnCCzJMvHedRS/vFbrn8dO3crxZYgpxzMSv1CK2w3HvYZudBtaOA
Y4hNK82kboi9wKXhiIduYrZUQk3IIfcSZU1EHxBgJpyk5vy06IFFDOdDpzW5NTWM
qdh8/lngQ8FbMlCxo4uzc21Oh/31k+rM6a8/fNWw+xoUTN3Ey2fTOARFPDzi/X3h
Gmzpws+pjW5s7UfvIOKs1vg6oBd152mZLBy9gwnF1hFNV6izkpP+1VbUEIb4Cop9
8gDhgkclYFZvXkq6Ynh9ukF5zP8i7O0XiU5YmD7nogvHlXFX/clhtsWnMtZFpYDc
kUvFRdEnMJma0MidYrmDvcDNRpKHJiDJ98OA4Pk+WWx88zU+g8rTGAriotz6vMoi
enjCa4V9RA9JwtzLsSeFhM83mAB2BD/uQIOTzCiAJUw2Za1XoYYSw0ANiRAgUgn3
q4d7O52/vlug0nitmFNL0+rM7k3VN7Wdtd4p1x8FyBZ6OcLsvikortLGVEAxzVmt
J3/JzAzx7rKnwdY3kIRfHryYemcmFwN9OtxWHf1cc9bOiQrBY1gVNHG1XLE2gaWJ
nbO/EQRv4s9uTTsyYu4ffnEklM3OY8PwZKBV/nzzWD0PWZSUq9OYXysm1ZfErKql
eSiknKfrox+d8Pi9F2TQ+JuvDmxYIJTmDCm7NrGXfkW+48Umoi0cHaV5bK4pcvR9
azuWF8TBfQIJc0+26kDjN1FUtrBw53URVu5Ef3S8dWs/xTv4FBJAtxF/JLata5OX
ZSmSC1yfjzjMYPhid0iZx/hhouy8DTRVFgWhuN0wxKCni4+tprYTZJiXQHk2q/Ef
h4bSSLN0wsPJCAZJ0NZGDjaqasZokpiLl5PiwYf6Id457qoZir4jH/Blr05aQW8s
gJQcsbKeMqRddydUoc/VNYj6cBtgSo28VO39fhOEH29lLBHNFCM+WfvU9XdjYRSK
HAJv737wSU/w2pBXjjcxxnllLw/arRIEqYLbAbFBJErKFkb0JSwCJ5z2pjGXK/Ow
BklZPlgpDxBCpzYERn7o+nYmlDWj2La8GutmUrIVoUD+471jPJxwoAW4+GGITwUR
y3Mf3VhlWWbnG+8CZy82Pp4uKoOVD9avItqek2ZG8ZATJk8Vb85zYkG7DmLznpy9
UuVtOsVP6nXVaPwuq9oG8YwKUVugEEbX3Z1phXijVpg8uCREvwiDwbzeGkLfJSRw
rE0Kt0xZEs7hN1hv3/KEx9WN7ZxVLjEn7+bYlSrieuLlG5V7GPVpO0cnYOZlEK8T
8LKiX1OhBN7hGQbo+7UyBXDLlj9tMTF3eAfxf+Nb51Ko61Fbu4bX8IEt+9PxEN4Y
z228tAQEXObDR2zDvB8hWSyHH9GY8tS4WheLLFFPFxoLUGfwl8duqJJ268NIBx9u
VEvWNLW3QA+wSpwUYj9ocBlouoHIyKwBV6F0QICJclWfBi0OqZaYSLnnJW1Kzw/Z
6r+kFJKqjakQl9swVxIlvvyPvxwvfrodvmTR+837LHvOdZb9rcIXmBWSYJFgoMWI
D2+jOey26LHpybLtrl4DDo+5TkZgQp0zucTcwvCiLydqu9WN3ErIWo8RXcLqE4FZ
5DlZZGJJmLkYL8TI3RwPCLfgCioQk7qDSMw6k/Vcl/1Za9eZCWefgL3j367YC+5q
YndCWPCLu8YLFdu5ItjT+vPmVPbIRIxvABHAmG8ZbD2len2/xhfW0Q15wSh/R6Gb
AvWH4jtY5EacVI8FaSUO3xU8T+4Neq01ou1ZpcZJC0bBJXikUEbxtLOQVehcef8J
YyinY0tUfcwRcSQkBM7B9RlvK8+fKSrPTV7n4egKnFg50B7a9hpMLstf3m+KKmCe
G3QXXnyid+xOFGC/b7GvEXzvxZ5fiMXPHWP57dwcNw/pwFegnHzD8CgVNyfFilRA
M99CkYzepbm4H19XqpsxofiKNT7Ivo4Q1f68iuE/XbcEaxzkHyK2FeK/h87O9uYZ
nhziJhaRhBCrYJT+LYLxSREbrOzKTIK6tGOhsivS/7hkzZqnS8g15jtLfofiSTGk
x9s7iGVcFytlGuv3BnYYYfIoFpp+CPMrGdoDGBX+ZlFzIfhr49RVXJ1I+DKatEzm
9prY4DT0tMjWWbfJnfyhnGon4wYV3uCQDtw1iXKyN1TG0AGrsz5VdhTfubzBeIHE
Lm16ZExYdPhJout6diZ/3y4iJfeTfXkE9IX+wpE9fTNIklCdFTyKBJX+qxw37B0S
2Yj86wqzLwhNoVGn7cujETTpRGuRs3KBu0+UzuWW2NUMZMbxQmPZFBKROrf4hutc
uNyEvi5B/zWCH3ONaNwPo1FOgVLKh2qBnN3CevB4KT3j0ow6NEqMULuzLEGX2q2k
443lzSYE9h4kSvKRqZSW2BBj4boaxC9NtilFtGaDPAIiWCH/AHVX1fGsiqb+ZbP2
AVH6kRwOtEaz9tenCZIgkkz7qvu5Fv2r8nC5co8uDuOQ7XzzeXP3CdI+3A7vt8+k
CDXG4Bn85ko10iKQQ/siIzsDI3JAKqdCZanq7hEYRGhFmZmz3grju6m1/2d3NH+V
lL34lIYD0V7wSr9hfXBJOoLhhVfy/kAGa0R6mh/NlL+ytfHPw2V3we7xR2i0cv6l
NiSSRckF24ZGfwss/Ra0qo0Yok771V6bHW03IG8w49UraasmZl1QAzttNT+WzXxV
SZGF5UrJmytPifj3JtrSJvM4+w9gK5J1zBpF09LwWb1vZHx1kkTwElMfloLPGCza
wd9Ngu1uUGs0+7rJ5bencC16VeNZIuc+yMfaPgAyi5Psvj1UiNr5K83rRJOrvjQ9
sryDNv5flYpiLMLgSC5MYJOGo584nMnp/vwrzrUMRFV7xRYVetKUm7dHQJbnbxoG
sZ8grCwcvcqfE71fvXhfXtJOPacZIwMgOPWRgqOoA872HxjN0485duDcVXDyomBu
Xh61mnkj5xW7/KyHghtx9/uUp7rmHw/+zKBY/Iv7ZckeSM/BzmIat5xYcnk/nKTa
BtKtEO1cVcpxjYLp8aNpisJLDd4wRTR6k66LZ65yrvP+mPyM5HtFh6f51oztKhn/
fGxTova18s23jQY6vAVNnLxcvfTN8VGoZZrCvGMITgUolVFW7BK7SDGrHogu2gT1
tEO9KRl58Fk9SE2ts0qDN4wJ4AD8wNHJq7bSBmfFgDgNlGjnZb7mg5pc/E21kJ0H
w2KXPHQUrOEgziD57NCknXIH+D5wuJCTrdKIwbJJPc74IoloTCzK6q7eiqC/kWQV
ZP92TjflSL8gatclhowIkQNqevVuOvLRHhqGXrmhBLb9p/tRW8jVlMHUaq7P1luS
0IJqWfobs6rcR54JooZFBpQKi4ft9juX7LkGlFRdDgos9o82vetzhtwgHEKxdnsr
yh1Yobkm+dvOXxj9l/USv9SWUhdFXU2lvjJgPfbN8W/ruSJDcQRoAKWdCO62cqI3
vYWZL+c3FGR4qd8/CeZ6D56CtnZWVacbWxSvJZV0W/jYun1EYnQEUjM2swsEiPeS
TdGXpmry4sKU8WIPWKGsKS5W3l1Lc2bKTRkEyclv3PtLkpIqJgUh6trAdURstmv9
bFHirIDF5SORwNbZy8zBDjSUlzJYwqxF4SKBXSC1wyqZAHe8di6mTmJWsitDRvsr
Bl5k+B3ykDt7XuD8Y/Q5/e3Q+e7w0LLTKKBY8HdzW2W9aImxMWuSzK0DHh1t4Tef
dVMWeiusrSlutT+K0EV5qnLH8j9aZ8C8hKrfZu5APCYoF2YfZffVEJLSx+U1SrlD
WDA9/6jqEmDUxj//sVkL7MBS09AUwpNTAq2MAaGi0UCU3Y9KKU9sB/iIVzmmJ7sZ
x35cRAEi7c92Y3ITZcj2IjXR8cNZHnmAtFvBFWzNMF4xkeHym1e/4MfW5eKTASFD
9pVBevNubUBAZIb2IqDNx/F4wSnUzkgEjpUOBT6SDfe4PEhgYMMikgUZZXlTxvhd
Gir9x20vxPR2zHjAjHgo7HWpyyDaU9qlWTCXxJsdgkEujkOZ70jeuPdRqid7KJNl
SHY4SRjsW+P4V1h6drXWLRb9CYmm99UE8+uLfqPsxfMSkRJlUyKi0ITNRXpKXniX
NUjXBI98KLog+9nghJlHK1CGHMOntU2Vhi5zGRrmr3VU5w1pEgMVZ89pWk2Oj4aC
CJFe2YMfIeNCJQA9upttlEC2KBa+yBkKfPTdaKfF7S0JB0qxRRZOEvcjtJaHEJlH
3srJ6ozr+FPSxEJ2iS/Z28KKu2H++xP9Qze0+Q1toX4+paSeUSji8UXloFEUQLzw
FfbXkP94M8u3TdsQrYxO7cv/FoGuuOX8YtVp25iqYfrtMN7uFug0RwdcrkTA71Po
nkDKRJVyfz+Jqz2PNqqYF1FQsokFi2F7Z96XR2OfAq3zbzHvG4Wv25MKMAI0ZxB/
h4GyJPd2eeKO8jt+dq70w1H738qgMI6fL5H5CoXvukakwrcsNDR25HSCts9inOJN
O873rUAhVgJJWENVwf55rmlvmmdHb33mCI8Onc/iIq+iwyIWNnkGmRPfg7y8GmIr
5SxvDXVzodCZWVa/5Jak+sGInGQIS3Roz2QbmILEGsGXQRMkYkg8a+QV6jHvxD5v
hmgrZtRz4IGxhcSGD7s+57xJtH/76GPjvOoB4raz0ncwAbd3tg1ZKOxRbXFGzVbh
pQfVWAAZxLf/LBp7P3ju4dsF3tTCwPhTM2Fkx9jFqauYL4frznmzxmrsz0QQ6K0z
/hS1X7kar8ChHMUH1yN3B9lPqOJk6MBl3OrOBRr9Dx/+o3c6UdcHHuSSV4k68AVn
kU0ZtAu4TulyZCm1X7WZQIDxAd6UeCBG8MsHDv19olWB6oJ/4eWBDJeKfbCAsitL
UZPzvNK02D9FRTrw6GGl+kxJB0H7ut4SWdivI6bIZE3L8F4Mh4sEAqP+KF9FKrZJ
h4quHUvXJVjsub4XprUld/o4ZkeegPCCLhiVLG9QYwaYGAW0PBCHTFU/XTKucCDk
/mrCcuT8ZPcWDUjntJJPerZ5PWwRxeHPB/v0APgL45pKUdnRsgBvKD2WI/7ToJcN
QLAo70A0Vnrxs7m0aieKgwXC0fLiHzXyUyEq/iJypECGTmM1z9JTjzu1BnFOQn5K
04HfZsVPd4afVbWy9hrmWee44izf6GY/w4rfdfPq/xzHgAk1iyCBzRX9ohwVxHd9
fTSmLqLE3d1rirtMIdi3RbC7tyoKebnF2avDm9Hc2KwTInq/5VqobYEvQ/9WSpVF
OvctSCUNoj14O/KBRUeTebsS0B9FTUx0b1wb14ZEZq0UFnlwDsUM70PCyk0qn6q1
NIy1Wpe9t7/mKMrxB51FlnKUIwUYOeDmuaP1Jwcd9EL76HzhJdhJ7ce/+1xTNVcs
VnP+5Lc5R9+teobJORa+JyfT+vuSisbiWuSJLLdSGkb0G1YgUPzi2/lYL81P0SeV
7Crm5K3DiFzYSc0d8HtWAOlvUNCNU+LMSjWAU7DMYMOIg8Cdcii9nalbROhZMQcB
`protect END_PROTECTED
