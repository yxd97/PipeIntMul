`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1b7h1fwu6beo6NkdAFXnFbu0A680eG63AA44b5nhH0rGCMbpTQDpYQieLNok+Ch
CUWxGvT9LmSfIebwnphF7+Ji4PNuaOymuSHttyOq5B3af8l57GJ7fKo+cDqxOg8s
e3NuOSOWpWz086/uQUk5xpfGM3cHjObxd9NtPev4264zNcNDbRplfnXxP4TcREEC
uYFnm5RcmvSm36MgmGHroAeLfEtIsWKIqmrROdIp+fmbs04/zPZ4MV2TQfPWCYrR
buBs61X608s57ZLKC9j0pw==
`protect END_PROTECTED
