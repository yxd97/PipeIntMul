`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q5uufUohyWBbNgkqYTrdoxZQIY/ZEE/LTXQ8zsY2N0XW97wwdCZoJ23h9kOwOXFQ
bDsZmBlnBxB2Ou7tSmegFf926zY/N2M9+GD5ehuE+UEQyPQqrvO8gp0nzwEcpNlO
PusqPMBg3Pok3HY5/bMZYonESt78UQBgBCnHm1e8YW8//96BLUv9JigqtvwAbDlU
A9BThz4+VT0yxKDcvjIK1O9p6Fik8XjOV1PbGhgkHIgsE1f+DQxIM9BRl8yg13zT
qSrEibXqjRXN6/NZypehTaSNsT37L0HjR4XxU5tBGsmNwwS8CEkpdE+ldgFhOrq7
QNSFGqrbb+NSrmBxyRAEGFRB5phUAsxsFSHtiSMFBCuw4OCMbeyXxvbDmOsA3nwX
5ODmxzQtyFziSbHAdmLLQ3s0nNns0rvnjDVSHa/C5fWB8BxMxnT9/HNigyXBc7u9
fk1u6lMQBhpSvM4RxWGrCdY5tJ6f7CWQyAQNYuGc9zPww/w4+E6T5hZ8ldYy/GN2
3S4mv1tnIonzTAi92AI6999LAbokwC7A2CEW5QGAmRcqTSgknoPonLEB6m9yu9Mx
kKgKm+OBJkFcOozqFyTtlNQU97j8IeCt4iHRgwPAupc3gD1dbfeDf/YF2ZWcXDU/
MfCqLLw99O4+lGWYdUvvAQa156gBqYlyPX4RCd0xRWch4pHrVgfH87tgyKYHmsh+
A+pcgGL7z4v6c1F+RDUzpe/pNZNy89LJK+ZJzM9E5AU=
`protect END_PROTECTED
