`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xnOlOdPLFdoQliAAVdbGl92Qr2Fp0fDmTh2QLEc4gAA4ygnNB8oKHH6VYgKsTViT
Xdh7sO713rGuFOgG3VIM/Tjz7W6SLpkJ5Enczk4oAQ6xeno63yuZrql6RgS5d9s4
l1zQY2RJxYGfDK0x3wj+1lAcOI08BiqxgCosKMasgDMQkDomPU/0yxvRrlvoysNo
PRNVMnVFhODudJ8oEICH/IfHkxfrT6eA+FMmja896pJ4eMSPBn9OaVoQg4wC+Gbs
nX/RflDBNaEDmnghVMfKbTOvl13WTAPhCd85ISjwJStgj/mDQ/A4v8V9sZmyXmDd
V8KgOI4v73i7kkST9dgfn18gIecLu+XxWPTi1F8bRAc=
`protect END_PROTECTED
