`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c4Ad1JAw4pakbrWtnLu9nGekM8BziLucAxAXgnEbpP/NVRcGhDzvnsOUEk5/mwry
mkrXESKEJmyNRref9V+y6EYeCRu0Eh8i3GJKz+4RnRWeWCkbxK+fOrL35xJMsomt
zIIFwHnlnTavy7O/QMxSV607lFBsw3j7K4JIwIeli4p7lVUgp2K4QqOnafmB5fAa
XJqY+xb7OmBK/ixg7YT1z/KeZpO3+aA1gXw1J7Gi0xOXm+pBmMQV650y9aIEH6xm
AFxS1pVAUlr9FRGRZHdbqUtgOGcZGcdTUvs/HLx18+TvgtrcipTg6U6iHaDO3UI7
Y8NE0rvKNquyNRE/ICiFWKkhEonMb6V5NG+OkaJDhXeaXOr0aagXOvPp9E3e5xOU
KC8GJVr/zlZovYDrmbiUDigYYD2t0o9/gKcrsut8qoI8RUeooEbV76FXbZiC3FUn
aQVkX7zNz+bMKYABo3bVrglpEqAbZH0qvZ5ljfrzEJvl45hLoaO+FQcaSsX73AUq
whHEuPQMG8qbCzJbqhEvxLuMVTk3KZ1hmTTjZCCQgMHB8LyUDJywZxel9t0hntSp
2S53qI4b+Tf8OZ+gUtgSn00XH3YNkh5AZ1gWnCMyTqXxwDD7M9heMxp+3rCmIdna
SAck6zmeUOXwmxuI3gCZfrdVctnjkVD4FUyuuB7A/S6M4F9QcKrmAP6EgEBLM77K
TjhnWJ0ACieu7NdOMr1phMC5AtjGgM+GhpZQCSoCZ6/oRrMJ69NeR4b/RQlvy9/e
+KaTDaSj2ctmlOmQjGdu4e35OSchaJOAueVAIwg0nMilKPL3uFq2hqLQTaEpIVn+
ZnwJ5caM49+3w5xQNxUxc7ctZQEtcSTjKv3Y/f7ytf0I7EvRaC5unqEIkfXzs59T
c69x6fyAfmnaqDMynwyfXpstOMlwfOUDcdQwJQWFcC2mRiAMAzTIXt14ssL/V7nW
`protect END_PROTECTED
