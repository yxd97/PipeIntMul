`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PiVi2u+uLeIwCNkLHtsUCc7S1lWHJQ/83Wt7k7q8C/G8F+GZI7+x33SUZqNWlP/3
BlcO/3URz6+nIA6M3n2lRop7M9MJMUKC2W0PTUqD33duey/DYnv5t5nN7vQOYD78
YaifK+aj6BiZHqvSNnoz0SsjuLdOAfKOSlHRngpqDRLu3fGztMBXeMLQW3oDUclg
mJTILeQ1fgd0X2pcVzZr63o8ofgiYsmWbJTDJfusyaD4I/3dOTqRINcTPufdw2go
dh+3rrj33xcYAFqyt8ulAHJt85LFlUirNDQDYBC8k5PRTzWQlYgK/lHIYqQPiXBv
mfZm6PI/C+9mLsjoP7mCTJUVUVObZSuUuyyTgYHMNeXjQCBRwz2qGDrVPBIQ3Krm
fr3uzB37TseYxm/qem3Ufu65+93Vh5lRwW6CV8EjTXjx7r8koWVZOhiVeRlWIujm
fDUzja/X/e12xCQnwcnI7w==
`protect END_PROTECTED
