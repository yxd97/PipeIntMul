`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ps1af3hxJ8vIqYiQZ/eolGpFzyYuQUQMIhywfFf/KMtCebxJah0JDCYVrKF5Kxci
R89O9zOdWodAc5gCiIuPIFUea4oTRW7gvkm5PaeC+P22hXodcCr3JaMTLqtPsIIR
uLz6SZMPurq0MuSXhdXoeUQgCYh8UdzngrpYY2PohsDjsdtAX/Hsm+TNTgxZErmU
v6B9uARREhp56bx9zGeLqtaC873QkPTrQQ3LMga0rtz2vZ2RsQsCcxyA9SbMU4mt
md1Tg6LqQH4dPMo3jZou9uYRjSCNx/n1eZuJKxBjY3Pbr4zrJM7/I/oEmdnxbhJW
2J62bKJcrTBV+EoPr3guaskVmXyiszstWtxm61XNyA+KGpZUsCR89EzWvWW1JBgH
501r857MWBlQuKNac4rqtWhhWpWpnAzd3rcH1z4EtTcQPlOtODfnAFtgER3Iphdu
Elp4DeIWjoV0vpG0lxKR8EcGI5/M+UaUnf4zLID/WiXMkq1J8QHc0ArPRdgeptC+
LEXn/d40yjVdqhhGYP3PTrT6cEAZtq5krKvu9VQZuGPdBteOzexV8K8A6YWRpJSs
g8XrXufq7T+iYif9jPyhDHHQrQKxsCKauG97nRim24thLyptJ/+Pny6HTVS9AyAH
6n/ZOpS10U1AOZirTVEzWGC8O2VHSqfIq+Tadp4NSkUvR0QxhazRuZhWRIsXc5B9
AHXJ21ENgEGywFf5q04YXcW5EZ4dWqdv1bprw38GGP92IKX4RcXCbbOx50c8Vr69
ZRrhr2TyTUh0d3kKDTwkVUhrVZLza4h16CdYOD5B4ycI8fvekcuf9nr/VkTemejS
LfBRPkDxWnr9Eex8JeL+f4FjxsIJWHaUBtkdTiY44bMx6r0iK2Ogm9BwLEgMXzo1
YL0bGFnJkreIovp7olAnncdsEqFre5t4Ho1fxpKhRHw6Z6B/2FBcZ+5tOYhnqGo7
jcJYPxmibgEaFfCqAuMGzy/WvEGwi1XnCOCkxiz/PYPCboZFHVXPiOq7Clo6b/28
hS0d3FX56cNfppRY32cc5zvG/hrmvCjPIBHzFDxjMNCC/rLDciu05qvJOmBojFa+
ReAxbwVkeCPG3jm+taW7q58V0BYkey7u9/XwYrwW38/LNrTOnr3GWoIBlKxTK3u4
u6XCodsYE+RdRF0J655xL+mC3ibCa4kJ79NyccIgRxNgu4J+lu02cWfoMm8b23KT
VupknfxDdf/i5lnAH0lKh2YPP6YxDGEY4+KqlPwI7BFiUgETzQSjQIRul3SNZg+l
Kq3LmWALaYbXUVMYDAORdBK4AmW5JHrHc13eUBIHv+SbQv97DKTHzJwpQPS7+3M6
Ch9tl40LcPug9KW3gzmu8HSN6uB9MDoTq7qXkkuS7kLK3K2Yi8Selus5t5OvzWem
BBQLyVguz0Apdwfy8Q1fuf3Q6dIjHZb0DfA/xBPYBdnKeFIQrnWMDBAAsNE1ueVF
Znm5xf2/avVYd4gOna33XkXNGv5jpAn5FeZppIyGWchFJQ1PvVC8GFPR6z3G/F1y
+hl5+IRKxcWZJ+QI6WPbLGRXzOcLEowOpehkea+Ee4yCH7xn2ginSlG6FFmKk3PD
1jgueQcFcBc+85yO7BB7RsEgSB4cxsJhF/Kl9edkEYEr145CKNol8xnuK3whx0O5
64z/n5L4dDJmLhCFrLNPQ89rUuMSm4QsdvkSoGtgkWnvy5NMimkrAzxlDWUGuxlB
WlHUxcalEK8fEBApXHpBsuMGZD+Vqa5Vn+7TuiNVKzc0xytAGMM5T+mmThPr9MN8
dfu0auR1q3DjNQ/jdfuuKO7jSGkRtySCQlQqVQL6a+Fklt4TUxfnyikGbmLpV57N
OnROZXz1a8u1CE3zodpK+Q==
`protect END_PROTECTED
