`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzG5QIardb3Ael68KTwqDWcHyidTolD/YmTA7nwKtq+fBITX3uSFYAlAlylgssgO
QMnrIMys8wTOBXAU+n96g/CEhs3FyQyU64DwQpL37sazuuxSnEfy5YqatRSbtJcT
LT6KAc4xAaFLigFcK4kIKeopo3S3foHdXqyeDYTdqEVDiF00KorkM7L1aCYnTxRj
5aXX5X6H80eG6O8HPlrqjyw13RQk7Updo1MGxv8E4+gwxaWzHprUtwji9U0t6EEy
lB1vv3tbGIZPY/mjrJCf+VwfaFohGWfgqOWLg+DgOLvFQ5sZIP17iDicSkR7YswK
oAIFQ/kNBhop6SfZfCWQayP06npAELOKcna6KkbHTxQZUubvUd1SpfO7fgBhRWH7
gPVSztWVLoDaZm8535jHa7Q3E9+vKOA44gjw7/LFkYJ+H7PxmHYl+Y+Bif4soE8P
+t+3+zQC9tMRrac8N8ke651xT7Wqpyve5CKX4Zbo/pMAo7w8BW/CMZ8EzShQ3hMA
9wo71n/wZ7PCDhwMTi7M6ct4Mk8Sc5cVgTHAtCdDCnx2D3qDw9sDBvhJEyfdkN3o
DVZ8ZUiPVEBRGBA4L+9ZfegURsnJInzqNlbBXi/i6c63LfTsOKEF3p6TbOzik2yU
d3MaIqQEkRLP+/Za9EnCiw==
`protect END_PROTECTED
