`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xglxHmzmIl2zAr3q2Uk0s6t7baAQ7F4GVDjpO3MKjNFAEPSOQ1PR799ikcW2fSbF
6qRCgCyXMdBNwJSUPKvWa8gD1ujIWqiWQE7SXMvIRoN+eWN4+8lVc83W8Zwf4JT9
+b24Yr8ubojgvKTCX4I6V8HGhaCUZ6rFGxfeJQXBasT0M2kc38h5Fu9BCIZPyYsG
7SGON9kf3zC7fSjK5rvfvcBhe/3lderi3mM27/NXLbxe+oLyKAx+EMoVomv5nUED
lhuOiGMGQQnBUEjD4ysMMX7nQGH2rYEl35hKviaHjuNHmFqpbuvxrkqGKl1dqyF/
hJYCbykKIPTpsc4Zz2dqlc6cX6d64HWm3qa6E4a78Mzfu/dTmX0lRfnqI+UZgZN7
fVlW9cB13vpPNNQ4Bg7JtLgpsbz76zNm0X09YntzPA3NvFtYRE1O7CHekyhiBOA5
F6MsnK6FqCA95f8fGufZOG+f9WJXlwj3b1Vma+j8TgW3SZPw90nhe1/Mp4NhfItq
`protect END_PROTECTED
