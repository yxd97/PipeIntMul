`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8bJj0yoHdpMJkXcLUTCGXsNx7bqaTSRxogl3vFmFwgEAUXamlFMLUk3iYA6dOQXt
l6lPDDlbOe0pYn3h2QCflva4Hg1sbLKYKQ3lXHaOMaIyXjWYCnIhQDUghZCYtWea
PU8weUqmGyiJ6q8rhL/o8VKj8btcW5r5popi9TELqEAiVigZsr+372L5m76KSTA/
6OX24o/BB3ZezAduv50a+Oiuuy0YVPghL+/d1m8ZDB2hQHKl/CQ/MLx8ff1tHbH6
t/3Z02o3oIhmH2dSRsZGPA==
`protect END_PROTECTED
