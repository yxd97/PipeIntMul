`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fU4hM0I2KvPLFUHtOYWDVUuChH+6ErbazLBGhu5evC/S/HaESupxriY27nY3Y2ta
5Fj1BjmsoJgYPrs4j2kaaoq3uityRzymlPGegRkzU+w4+xJ8brD68g7swmSHLG6f
GCt0+RXKJQdhU8e2xVfaLyeFaO61CFBoZag461Rf/dBYmpmHwEe0XO5ShDrGSVPv
ldXBZN0YKCZSL+4SBcpU9nyEveqo26f+47wu7feqkAXpOX08Z7pZEi3I2JMrVmM8
qyoYM4uXJv+N8Anu1QFaumi/VNw1duHIH/r9OMBoGsLpL8zoQ6MWFAcJDKHGrWhw
rqUCIDD+pO0STdoRTMVIyQNjeqlrVACEgLWLYnmsZoVpEzw1N7r44zYa1tp73dNp
b93PNn19Xa0x4OXxyaWmJQSqb+SSP8oBorHW0/wNA9PwxKP5LMmGdOYFEeePRcWU
D0kNCQyORMDG2Xtg0+7cHmoBZguhv0mJwTmR4oyZujzeJSM5N9CDrUGKdP4ZP6mx
u3SkZBbl/L+7hJu/4AlFhA/jhtiMIDcK38XAG7UKdpBBEAA18lU9VGZztsLyTrnb
cCg8JGrcigf9XfhICcSTDOJxBR5fbTQPdwhuzwvXF1J95k2FeEqSvtN9ErUdQQqc
Jo2J7IU/rYDgs1eCYjqU+vHFbHAms8IC8uOwM89HaVeJ7AuuED0WZhG+tDV5bEUJ
Mx7q6S6jApPBBaSSBtHkIaMGVK2eTW+dVwzBVtwL2i08HT20FV2TnuA2cDOWowH0
OrnQnE405zMVbC04XT7CyRpv2/sq9im/jrR/cSRS9I0mwvgqDC8N300K8+McreVR
jtyCUaW3emNpO/vVyfgng/3jHZ1wsKM7B+REnyjrgmL0bNhiU9X5vspD0+T1JeH5
PLHpKghFLLG5UMxGo0SgedvD5MGv9d1m4UrWzt68bE9mvQ1gb01tPM4h6EBN6zSc
9q1fiFErvchRYSMnFPjP/hUf64S/55zAU+fMW74Mpy5ItPALkvYLRHGqT5wbkxa1
KEcpByDsJX7HtZA1XseCXM3Vcnn34nPeOzCLoNRFprG77mcVFRxVSnhHjlSsOOlk
vijagmetDeQFZ43MOfitHf6njoy13CsfreYn3YDBFD6z9QCa6I/9Vk6Q/TQ5Zy83
Yry1JsbuIfrcTo79F2+sZ5ea1vZu6JaRAGWaSrK6e3cMPp+y0V6I/NL91hOMjNPi
uNM3JxFqSfKMyWTYuADUIEcIAlm3LXd5mgu6pzY8jX6YQ79KRQYyale+6kT0ugxf
ZL7+i1qq2tDEpzeGuQks745bivT9g1heDcsualMxLrro70pxzIYWGUmns449TrMG
+ozxDsAuv9YNDN1vI4vR5E5Z3Vn7mWFsr9o8wxVbLCjqMzVOAoPe/E0/yyftFLcr
XP5rTcytOmUNescVcexFo2c8RnxSlQPOZY94r2ZpdV9bT9E78t4vLa1VUSiJQMkI
7ufVogogfv9leQpB6JUVJ3KObIZp7FD+HzcSl77uFHjafvrAfMycdviHDN9i/XGD
11UEl/+QgbeftggIeOTZk5wCfcQmD5G3PtdfQkuZjtG5/yeJHMkOZOUA/HxHIY2D
bD6B40AahvS0XAoPu159W83yKAswBuoc6L12puzP91pfMFYUxZjqB+ToaJOiVWXO
XpJHu9qstfY+rVv1WYaUWRbxAM09YINxBllbLSmkvYIL5VD8XMvd0qC0xigMPhzz
pHoI/7066AGIFwJY8pq7Fw/KQ9rmqE1c0ckRhOj777m6or94KQOEkC9NQsNygaA9
IB8RVrviLLengnG2nWBKCyQ4jJk2syybZrGQRq/0jjBMXQSzEXWMRXO+6gLlK8tV
SPhmdkyuXRguUAqz9gcMyqHv4wLaMzqGl6gFz+jjCxLRLMN022cwPkm5eFqWLttF
nVKs2MXeX+aIRirFKBKMFbyg71cJjzyX8OBjw3jtTruz7gVDBFTGJY630cAi9oDY
/bx1K7Ct/Xyyog3P74WwjL7leMBpesmNbzO4Ym6HeOqLlKsedaytY0LPMALqLuNj
uauXDzssMSNfxNVbOMmh24ZatL4c/BoKt0KhiF6cNbdOP8GL90OCPSHmijklu24j
jiWPyFnYCVi4ctOIAtAdFnMIsTdFadnCJCSMliThMp/2NHBXYKnNj5cLrHUEEABC
VwnH1AXMT0Q+tvB4ZdewrCB5WXZjZ6o/tOpjEJFttWkB0AQ6/lDs+q5R7iY/AEOT
ewd7lAEh+RlSXKX6P8yHrYmwCyWTpQNUAGrRjZ/hExSNT57vHRlw6qTxgY071N5b
g/9PHQDPsJcD6HldjB94JHh5pM3Fi7ycMBMe8CWdVMJO+8Gqifx4paiHit1Jx4k/
uP61whumrmv0DZ3zd6GQw2ag8i07sg5SywDt0gjyI5/rKsyujKnMpMTH4CMb+zwe
QQ4LW2h9qYUDC97uQiBCK+szH3uwKB1EcA/47+s87A1c+Q+HTANA+qf0JsjwJSGL
VTfIgrJGP+EA1nlFXMeJdmV5amOEImYLpomGXeOh68w5Vw87I590zptDUnBxjx45
eMkeR9rKksPeItKzBMQek/PiV1zrue++O1RWbkteC3nXvBwrsf5WDptzFXg2JdcZ
K3bs6dnSlpcgAwONNpxAw0SJ3hKvV9wLLJhTAmKquOMNTTd/GrCgTrwFk1Elwrc6
AXVHUlyxYEaCYrMg9bHLWgO1Nev3Cfz98Wk1Jd7+klrViGIuKhazXazgWfNPmPzA
HH4zl8J9v5xFb9l5uhs13EbtOlCreAGUIOlrv12+nfyx6Dyip0sU5lIu5TeSZ1MY
qdK53Gea5TLP4iOvDD/8RWUMaCTXkzg14nihRdmYVJA571Zj6hxp5NdHyRNs/0ww
OHM8I9nr9nKbDWZK9pX6yrdSfDmijMaezEfybBlD1FqohMtRmhaq6I7D+yBdywrD
yC9IFXDRuoKd2i1ZYDcNpyYMvTpNSpxs4xCUsGHPSlPIQ6lYofWm42w3qJOlE1Mg
mPiKvJvvlDBcxGCnmTGY9qrmZF2VA0kWbeE1dYxcudxNbejAuW8+GRQ5/sfxf+/7
Is3dkBXkPM0URgbOXG/4x1HOzq9xc1PvpFUdYD4akJCQpGpMQGl5qVnmf4+7iHwV
ljyfpfEWTLaLlZyvP/XrniBENcAj39TH4wLquYHAAMrYuC1NLlJnI4/Z/xWr05bC
Q3+ee7vhY60T04MY9khbuclYvXOttPCV+E2LnyAzor1pCzA+9WTeFRHQzs7YipRv
WLkyVn63VsOtI5IAUvFjUSOLHrYeiuosOH6d6BB1JpDjFT5/wbUsCb/qUCRAD5Lb
sEzowk0uIlL2DFDhMcpHI1GQumNmQOhtdnCT4APkICsdJLiAVoCpOTl3REz8I84f
SRZbj7X6wLt3DXJgG7fZJ7HYiaHwtynqKPkR/P2JngaMEKN/FKcWgBFjCfnY1gO5
6BgDUFHMYDgP4nOwtOMISp21S1vdK7dc7sQs4eLacMD9js6ovnD+o+IjO5gQauwX
7Na1c1hUPZhsumGW6YawfLVBuqa/RxH9TF6rD9NOstS0CwVbhS16cLDDUtDPV1Pm
e5fAANeS5vO/hUcB509aRcGNow1qZ/02AJT8XoENRWNmyNq11UbW9iLdyq2XH4uJ
XUzWmFFDt00zcjxAEtcf6BRrjm/qGKLG2YNjD5SiBXrJ92e5jHtzvpZID3VU93lK
eCCcwygtHzxGhNKFL4CyStkknmc9kuT7vGD4aK3RHG1SJc27AVS/HpcLw3SvYtWF
250UJgX59vJsyfd2BUkTH75MBvjImcUm1RlBVE2846yEWF7cek9sNDwzvLcwBJKL
+hDM8ZwOupjbg4KWpCkQV6gLSUePSFyK1YUj2UYVtqShRytQ4HEsdxjAakkvJ+rL
FDSkfSx3kS9lx8v/Xs9QDVGzGI5Cm6ZCtL+sM/oe2806JTlG5TH9J0giuJ2CZaEO
0Gyi0PlEsRIiw3nRkrk553p8NxNduq+IYWjFEJD4mZr6IhNVioUT1NyF6WCCUT3r
43QxZnJSCe5Z5P0vq5R+tJAXXDr4Gg209aEW98y6+yDpmWAqmg5wudtNfxFf+uT9
2rHtA0+5z39zwiJyo0j3oxYdUyFqZ6/pqqHksXMIOXxB+vrktmz7E+2sXYu66mPf
3l6J04crNn5aZxbPe972bciKWHhd9Ek8bEF+6Grqy0bF0iSXEa4xFIyFshot1TX+
vPTU8KpbWpTB/zE/yCLOkRym5ThGyWbzb1+VpnMlpumso1Q7KjK6n1Vfc3q3Aeco
bQEMdn+8nPwUiDL7rzbiFh7AVnzi4mha+IUbtzqqERmJgwYsJ8gTSDh1AHtuTSkg
3a24N7MgLvNjhH0m2vzR83Pj43vIJk6BgozMmoGWZBFyvLDEM/mXCLRE0IJYvxkZ
qVvQclOXUSukl1785b1jsjgrFWpMPmxd7gcuxd3Az8xZg0XU4HkhpTiZ7AYQV9m5
5XzOafJjYp2hIHRkHa9AO+bLLrV/M5h1gKzW/64pEJv3kZ9MYIl7oko7/GF+H2gx
V1qWqF/Yx//q4P1GZw53CJA7KFT4hQTSBfk8gtKM92rfghCHT/Qnc+ZwpYGb5fmk
91+qOSzTY8YGCtaIK1UcK/e6esxAWZs6+JBugf9NUZubsmNqVGHGkTx9kGATfQmO
Qzi+cNHjNWu7fumML20MlJX/O8zaUl1TUOji9bZ6bj5iL+Kg1IkCDIh/b5ClpmZG
X2q+WwDN83x9WbMn+kjj1M5hFef14NcblzCYeF1kBbd+ccHZZp7+I+onp/dziwqI
kdUzFpuhOnp8vAHLmUb3iiP7sSvLaTVim13gC07tufE4pGxLNL41I3ePpMBZs+6t
dw3ZejxsFJrxXaQxUboSjl+ZM7lWeVkaR4z0yRlkgjs0A8/hJJYyVNyFp06yrAy5
XTdHCMEz/7rfNsgJFxiF46j3g4HIIZJgHPMN+/R/DjtNEjTSV7cnV5JYGkQRpVBr
4vTCygB2VCRd8zk3Nz3zog==
`protect END_PROTECTED
