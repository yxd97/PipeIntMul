`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqC4FI28BnAUW5AKXsI74KQbwaqydAlDxwasb8agGPAWEvuhRsnYmmzGEAneKhRT
eAfzSSNajqgOf6EVtfhyKZy5hamVkRy+9b4wL0v+bSIbP7lFuwN+VgoN92iKbDDO
SZ/l16WFPyrU9ZajIadSmk1kTCmg2jEaSwJs73eUjS+Gh/U7DFc7Qn1WptO5txH5
sfXJjvPaFo88C0wW0hSEyvimZuEZJAcUxZKgMX5N1T9popUKGP2g/CEH5ELWJplJ
ZwTzTSnMAk80t35numzhLfQ4uDPsBs4wNVWSAnZ6drQTTnE1ZCb0SFDlC+oqyoXn
YmsANRJzUFr/G18cPDUTPIE66FhKlTig12Vu/8eOF0vbYNBUMSten5LWr+GEB+/T
CmnlQxRky5kBcleXsYkOlJ/tn5Hgd69jzuWSgfS6gJXwU+jiIc07p/rYxkQ800vg
RtG/HaIu9nr2B5GHU1l7oJ+xmdlp9oiX1nG8e3duxV4=
`protect END_PROTECTED
