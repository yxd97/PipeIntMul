`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XDlwyOfe+3wvpNzBDXb2xvQ3S2upsz+zMXpYcdfo0UmICoAGjRy2e2UArf/koN7v
XxRjE5Tp+uuyBNPcj3AFKqwgMzKfMv182JNgzeFazNTOfWLlQJ50mp1vByFlN0xW
TFN5HnMr9MfGCiBjZuqjHAOCSVCwHob02AIo0+K7rxDgmkTSL9M8lSW02ewINaaG
t+OlvKstEMmPyKp4E2u08dIBdSEe4N2/gwpvKuOun4a6p4IMVJFy03oSrrwDnf6w
u98rl1qnj6gGEFVcn0iFeIjX0sPakwTOZRU08hN0U+fL6plx2NUSwsgbW6rHtgo1
WXzDSTY9K095Cpi6WATLRgM3hngButhU23KfkQ0CgrvQZwgpFI+Y7AmdgQDJ2vHC
MqjzQEc7GjEh30o/UaC+bNe/E8unum3OWyNr32GavHeDXdUT/mVDVDdb1xBU811G
RKDB0cqqsUQhhjrwqjNpUW0KoOo+sJNjhJZiwcRIFgmyuzaJTTcmpOfitWlrEHSw
w2dTpqOKT5fjgMkBR71iBsDnbZdOkG7JxQFYuGLrTPi+80SAy2/KgXyw00hGaQR4
0Z3K5ieZCD9ATu/ZTDJuDYf8UBRZtZsvNAT/Vctyoq1M8qnRgPYH+hNUwgQz7GdP
o9k1qBLBzET+zkUbCjCo2nZlaIpdcPTr434f3OpoEidoDhFQzLOpk9enHMjaLM0x
`protect END_PROTECTED
