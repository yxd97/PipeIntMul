`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yh6LcIrLmhJWio8rlGQpb/3OmBVUL6dF8mXgOie8xUc0X4lqm3Q+x6nrnF3SDmhF
MxNism9b3xukrCZhI1X+Ml5elDwnS+AqBKZI/gg64USJYIf1UHkiMbrf/tz16jCM
2JwftksBwrA93gaL8lT0qbNWmsLzP5T7F4yYtkNpasNhc09TIRBS6JLO+nkMo+LB
zOyWPAOR6h1mFoMTMcEPOu4/+/8siA/eNqFHdRUuIzehcK06Nb7ZQnR8YsUIVWSi
Fiqbe/HbtUb1NBQmX+WATGqv4kMZ494lfF92U0EZUQ8=
`protect END_PROTECTED
