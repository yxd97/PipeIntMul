`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
93Z+K2ZQ80hAHQWNqO5yUQPua0eFijhVZQ6zW0vuv5iOyK2PYVHySD1DPWbV97QT
8raLVQsxqXiyEIlKcdr0ExCoHzvd5czLnA5ch6lz/e0nIcB/IxIYEnjNmYKz7EeR
g0bBfLLyKirwcqIESW84ATf5UL7zYk3yg1OU/2JfzClEMSITwEqzZv09APh86bPM
7RgihNFka5fETSBY2HJCiVCp6pqc+sk5Xd3iFL3F5qj0h0kt1ASFN9zZ2t8nsF5I
nLfyC4vL0g4ROswEjU3GGDUGedV2HW6jaC743j9taYusAI+65NyNBeywylaSD9+v
I55flyxtjwzO1HtK8cPfvW76w4yljZJvNNTF6ESSanqbr9N2dG/rY51hOWQMwBXG
bqwEOAgT+dGBrNGF25K8f44ybkkfu2ZIRKdpVMJSWBQlMi6Hnbk/gDG8k26SSct+
CPXg2SKUTI5TV+J7IW+am2NxbjxEF/JbMIgcUYM9r6zzfv9pbdF4v0NHLcuh7/ot
46iL0Xly3kV4XwmRvZdkNlTsmr+01KrOzu6NRYJhc4gBfszPcfkNkwG63vbN7Ajl
`protect END_PROTECTED
