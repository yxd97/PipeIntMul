`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AStHLHMWgFbNsi6PgKFKK5d/4vYCVEnw3bCHESEhf/WK718qJEVX35gHFOrDSne7
yIN1+0lq/50G6x5uLIwpDFZwo98/Yt+3nH88aOnw4B1H1lKUvZCt3PCtd7hTW15b
P33N0Z/Fs/wFiuSYTCAjfzFS5iRNt8ZWEwMHz1Q57DMP3birOH/0JOr2yLKs3XCy
xq6v7LPCAdvyGnmA0xres5yc985XCVfHGQI4qEYu/H14TJc7IstZ4mx8baSIHHf3
jhI/SovReuCYBrO8c7PbBecaXjetHAjLYgVqVs6AdfVL4EXGykmB129OWaKoC3ow
I6UP5nIFf54/tlmLE2o9JacgGOAzopTfcBHc1lanKKtnc5/yjyXpWnCrHrRZ8/co
yaL7wUFlJgWjSUM31Bc1Ckx1nibMx/Ub2DdadT3R49xTy+aLYccT43vu+HtdXavy
a94lZDWw33vGC6WbRTBg9huj0okiDXvzXaQywA5WEv4Zl6H6xRDtb37JLLyffNFJ
DBt8Au1qVOjJYK+sSnxhCy+LgTfajW5fufI0LodnaPbKL+/XOAdeFGOy7VrOkm3I
p5gvKtHWQEMFLtYTjjGi6lzu0pM2r7qG0tXpNkNcUtLw+GQc66OdPTB4ibD6Ctt5
W7vtbMlWGrTmmNoJSOSNmJakFl/fKNrGcpbp0a0XoiDtmL3om5WcUbFze2L1Eg08
b307wMu3Um0NlGm4l/c+vsUxpiXFkbW/4cRUwVx3YCHYAeX5dwbtE+0A8JkhUIUc
R5m5SYMSsqvqSNL2qNo3aQ==
`protect END_PROTECTED
