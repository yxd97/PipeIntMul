`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bj03b1LvdhZCuwggzvwNNLQhuoDbv2BVEtPrryQ4Xstpnpy4/GO/cCM958PRhNr+
4YAGNseH0vCnOiZt87DbG901xK+0bsFbNC3P34QKuXU69wBPeYSvAZNN0TE802sg
TqVEsAIwQQszu0reP+3upJG37kjLWwV3pnCo0NssWlRW3+1EiLxdIDYE0yVi9v1G
xnkKM5Ro8pnQm6U4tAmZpn8BYke2jaSqrOVKr/fmw1COPfJFee0gyI2Z2r2L86T3
VGtiys4NN4HcVmYSx0kRy2vEmVZYjyu0+ASOXO64GRAqFKpe4bxx+aUifGbnbMBB
Zk8jwJcf/i+fLLRL8poXEF+AjI9/aJyFvv2irg8WPsQhLEdhRwY+OSOUEN4Eq+8R
i2xySPR4mlhCoPBVvPlLNsoDA+plevFSx+RZyzSpQ55ttWxQOq1oj5wlNPN/KLBo
ErOTJvqXP7ie1RXVvpegSdqMLdnXYiFSGihKhOIejPzCejGfdhKMmapNqVUoX96q
982xEMJ63BdHBQfragTJwa3o1pX25MbD9iTAjD1JboR0kKFkJyaysc/tPjjIkJHW
mXJ76sg8iyiOMfhwpc459paetYQ5g7EwAtwMsEljx+GYKUvJYZeQTFa2/CuUpYk/
mujxPgvNCspLnUxWblc+7Kukl2GLPPXOr2T9kYWp4xRi3ySTVhCOykZLHaPp93L3
M46wRviVOvcjv14LA5oJJ5b4EnQdKdp2UGOVJI7BoZgGvv6XYAt3oPShbIbjfGCd
E5zVwu30QHB/TGv8B5AqoGnxkkBnGlOlD2+9HmQ5XhdzNrMlop5RKr2T2ipBbT36
sjamC5sPGRcV9pyufM8waFIHZlFL2szUDCjxneXxM7WZZ+rfcmyXChpt6sAuvgKl
zbqgMwK7MZb52uVHqaer66UoOrOdUVoreG5HqdQkxxVnK7W53jEsHIYESLKhssB5
gwliToUTPdJA8obMAWYOa9I/YP0RzUXFyHDEBmCi9Dcd6D6S3pWHfTJ1b2+7g7qX
ax8/kphO1AJxC+bIq0AQSkVNeESHgg6VF9jyT+g/wgKOkTDa4gIqeAn/tyRsDik9
Irj4mI6sLaMZxIxiuAzVeRJf0wzm3fZ1KTP7ukqYIoy2zGC1uirhhv6auHXSekF/
/4o7dNid/aE8GF7XpAQAMOf9Gw7shlwS6g84I8L4E3QQ8g15gfnTCRTXqfhNK8ko
bapKP4Q147PwLSUVYsNFB5DqBEQFk05TyuLbOQf1Gyf+TM2LmS3Pjj/DfUImIE/I
X0GmrDAzm9k3O0nq17q5x1sAPSkqsxIzDplH8gET4QhQlIZB/jhecwcT5MuV9OiA
3NO81UJTMRPi1z6tAWoxhUTTHAApe2jRM3HrN+jzuGsuWc7MtLMDYMsGCzwSQFNx
N7vhcqnjcclt279OEfKV9fUmNGFeuyGdwFm/4kqZoCxmq7zeig4QT/GePI6Rx3Q5
M8ul1fWJNegJmSwk+hMNU+pYekiaSix0inO8bBIFUwApoWmrz59rP2ytvnORkQ8Z
cdFtNmn09qet5K2pY4KPx4k0Tcl9Blhue3ugnJ2qr18+/Ez0dwPzSwf+iQUUKeUV
mNJls4Cv8bvX9GWfz8tu6x4Gb+7LgecMsRO1q0aKxNL8DJqM/PCgymxeddOl7TXe
Ecyye+d/Oa9HfaFFsdz9bGvhawQC5qFixgv2mT1kEFbcnguoxRIyfb1OX6NQk6A7
KEtVTCiUMC0+52kX60PDRa2Mw40MocVoqNTKBVqXrEJ0bTlve8s3+m0OrXluPyBu
v/RjoXdfSEXE+odOdKXSE/emkofo/rJbnOpt4r0qMJmIi1Mo5svd2eyj89kJ1d/K
tffcICrcEZqy1+6eps7gX9YPe4BuzG1+xzfIyDWuZxfNLYhY3HIw3vO8hAcrEGDZ
deEHUgn22cRQGQmP1/R63kQNkVtQypwM7HzugyuOq3yzrMAp18dV/uHMfGcuvdF/
YS70IJQW2RpDPIgIJ/e7Twn9BA1fUcxPnj70CnJHdqSYP3hcx9Hyx/nLlAd6zf6B
UqtM9bP+PMggdCKMcIRiX5cDhbGFTs+WWKHw/9UE0GjGDgIYIbzgvrgcDAui9Uib
lAOmgRB6TXRwPiZs6UyLyqm2PyJsECA6FgES3dwXKv10Lf7eAl5q99l9W9yW4mi/
TDrSyjs1sXGchKsG942SF4eNcn7tCcu0NNf5/BMGScioNPNTxalPmrEAJg+KUHa1
0vyvPqb/FMY7pLF+krBtcKKPiUDdPbx9M8Er0QIQ5NRxjP53Wdh+1fjoxO6qENaB
/TlgWdKjQ9/njSJejtXgeK/tOVWGnc43GlzC2MjhLThk/9/MHbFNh+JuJSwcrpP+
fGxWqcAZ44pF6l0/iQylQIPMgazcQGMNKwFSGNXplPcnmSjeRAhbXki2Zi0rV04n
i8M8bOz+v+oOPQ0KQYadl1YwugXZ+zWd7PMf/spULC0xV5as0yF9SzNG2Up/7zke
n51k+XP++LiXGv3a2l7u+NNNkR74YKJr6x2zXmQa9F0h/MLa7owxMkFlMPCmVHuT
PEt5IZJYCHdMdDAliTClI8Ewob5OO3Kq4I8+NgEu3plHGsKexnN2DZrkLNUfqXPo
Y6JIVNqym/0BNwphYb2b4k4D1/i8FfLM9Fk5xbrd1tMZ0Y7h4QiB7hYMxo9y+Wnl
hd1fyt3vgmLGVSTBZ+qvs8QLvPyrPwa5u1621/MCp4T8QOH02/EQCp25nsA0NipL
I/vWdYrPlQJ1baXaY3KDwT4o3Y2RVm/2BAeqrvYHmxCGCYCHxFJCaum5kMsMEDK8
2SSk55fJwB5FrCdP+NySqOyRHT2cr4se/wP7VWxJjuDGCvVCZxUnhKiQRLoiNRxA
5SUv/RAkKbxAguyZt6tJsgNaiD3T5M2WJw91in8t8NFqWPZOCBDu1x6LpFdwyXbt
FFojX1VLFGpB/M7eZaU9lSM9wvbnO1uDzYeQrRaPzULCMIzGX6G8QCWyavAOWG12
gBz5i8WS2Y0M4i/Gv3BSY372y43/t/4c1zaOaFUT8Y0FN1aoU110OrFGCtsK96b2
GhfDYvRdGExT2dmlMA94jr6qe9V+c18GPloAmpoueRYTEzh6fc7ULrvkbbdhW7NU
gPfWquT5wPTVKMcaQUzt6/EgKti+Bucqvcsp4mXqKcEyznl97cWvAkwfKhCPxV6S
E1/Uhr6HJ8N1rjXrxjgv8SBJbZ6ybzod4U3kpBtD3L5jb3vpCRvbiH7l95m9/7X4
qbGvGWSps+IRMzk2IebxNDee6ELIOLYswPMQx4cWcmeKh3chH9R1NKycZjUwi9yl
jP7nMtWofMxk3RVEyf/Yl7BlS4c1bXvyAKmO4T79zcHm6cFaUBBe3eB++H8vofhG
PdarxyEgxmMR1PeHmNdDPWU4a2QWIJ1QwY7z8sQ2uRj28uqGNXMMdYCh9u7jXjVc
LfJ4DSyh3sa3aML8CWyNy84r9NwhRb2PokhHIGoagBhH219DZOpsSrqZq8zgGrrw
AiQblt+uy+CQlsJJI8J5aqhmyoSl5lE/pXjXdkEnzM9cHwivlqooVjIgbfw35kp0
DUyjXoP/7PYQEb4UVJbvLo/IYgpuFTwN5SvVjUKsFAnZjvBPMHMvE4mSD4zG4zyF
e+I4a2OwnOaag2PNXFfHEJYZRwaZANIHPzahfqTMXpN1KJbKfIyhnc63WYdDitlC
KtMNbfrpeSkwuJ0xpDPXbA4XCZCZrcCrhH7rOItnwiFtxBCXc7nIF2Pkd2U6IR79
MtXMzBp7VWQkgW99TR5r+Fp/r94H7C7YHe73uVgB7I6EwXJ9jFtq41aZ+7IVhopS
dwL6CajQtoiqENIlQX9Eom1sSqDAmXev+jB86Z9gVYyRyy6LPh3o5UXVf4WdQwaq
2F4QNQ8ckJU4WuK4ZmEvR9vaTRMSH3UT/kPEwOZxA5pC0YCNqUti8YVXMpCu/l15
Udq2XyPchxrhgVs2RBWh7z9VNpDGkHTilMSQcTqWy+P8JS+OPITz/r7UjDskIgpl
3SnYPoCfVqNZooBxLGX2IHT7EJbnO/d/Al/N6/YYV2A0KLfiVIp4j0y16JpYiXIx
F1z0JpKNgm4yL9XcpusEPwncMehsxkU40OSQImSjz3KM8sBk67VJ96R7LgB6nFqJ
zhXpSTC5bZwDYSx6/zpBK82ekxzFzowZcLpe4cQ9QGRK63f1CipjYwmcgRrr092u
dM+AqoT+eEa8TYiC2kAhuoGTczpNHCg6Rc4QaRBBcmXZNeGUhjFunjilAoS4CtRB
GMbavZsJrx8iDwaD9XesxVt8qaKpVam4c2gucSMlss3NQr8ikTUCcP4Mg7qLG6qM
HW015gL94iVWv6jgHs8PtpUHcexVh8jP6+5NQPbW8c+jWlULB7wrVCXOZJAK+2Ul
7WNvc7x7yYsbmp0wIH1DfhXkQenxku99iZuImKWRbJccXqy2cOVBYZYNVBHlHHjY
mt1VwYuQmfmDUzoyNtifyWqiI88h1dncdUvAbyldIP5m1N98ceGgSerQlljamAlu
7Y+VEwAUyg6PhgXRbVWg8qMHDdb45G7o7Een/vp1wypM1TcQqp77FrzY078nO8rN
Ah/3Z3+jb05FsjSyXpM4WhynDg8eCjxcXNKK3WWTG5lCUpcp46bNE/mm6VcbOPDu
flvDgB8Jq8FQrON5bn0d6+id3bQPOJZT8xkDLInhq4XYs8AG5oi8UAr/kCUDjqSN
8YSRXsX4cZQWvTZcvpp5aanZFXzONSqCpE8v9k2coMI5uQHF8AdvDi41EmR+KP4X
ZxHsP3OfSO7PO7agY1mRqDUTfbf4Yf+CFsYD4GqdATNmK5Mpu7YtHFVDelIpkmU+
Q8lrFSNGc22ZtAetjGZiQgXyDUYWjozsNiwb9KzigasZcNzdUvIp/mN2ai4Zw8Dn
nl+quunBIvbvAgUhofiCZTchDuHAG5mkMDezsdM2pmVY0JzsUBusU4sT6UKRgqmQ
i71WHQxpKx5nq/Pj4CfcB+h/6oPAtNTDD6i6vT9Vps2lHGsiX68zb984ef4VpQaS
18bUIGuHW8a8QL0j9pkw8isPfQKtsmrfrwKh2FtDAp4Rwhp6/jkKR8Ir8Uru3m/3
4kMlw+8IL/N1BM8uBEPhPJPDi0jvXnrxFME3BGxyjcutUee+Xx8XZqIbP/wX3waM
iUOjTWvsAKEJH3g+5CVkvJVFNWiZ+MlcvWx7w4JPkXDxGBDA0zB013zo8gWMN0GE
0P+s27Dst1spZ1wVUZEF3Yw2Dv3fqK1PJRyPoUvr88dLiL5GhE+HwlGMrMdzwWkh
hLOhp+8F/k6zYF3b7I1ChCfo8VylO+YBLcbRooLI70s7yI6xJ5suJmvFAvy9ZRBg
eJgOcXon8D6lB8BCnzenEQ+tTp3o/20k4DKODIJJ7DnICQyL+BPi3jfstsnZVODd
Pw2+lZb/SHJMZF2tOnNw8b0rMfqu51n7q+uKf+tZC+B7eFZrjqgw4S9Eee3aJwgY
gImkecz/q5YWT5dwp8syP95kKvv6WjdKFWAMFh+Ktcfcxd9f7X7ILrqeKFBEK/Wi
iYyUGhc0iTQd2meIfJ1qwCi2L7hsahc5bs8UlPEeSTMgNw2gGd+NQBwtduSpO+PR
9FZxD6LzIDm7U16eix0LPwC7k2dscFeM42UXg6H1DDlv5z0f9WG5NRQDrUJEmozo
1/alfltF3pQjXsYGmjq6e31rOU9skAxVcwysfTubeXaWhSwbMmACfrP4itGv4Pfq
F9+qIHbGi5g9lLOTQ3FTnybSibkR94FQIRjFfd3SAFxNWMNBB7BJ4w/x7JzLVVnG
dZ0JDtoxTM3BG7uQvlHxN8UvAHG+jtx3w3iZblxhrUYdUGfoZSw9DFd2hB7T6iaI
1ZtgaZGQRfHcLUHGJyFRpqZdjf6ZNZdI2JJngyujk2Kge+HjG39bAOFmdWUfzO6R
BgZIGrwePuKlSdxI6sru+3VmgBqlNlKnImEG8RZg1ILqSKjNUdKSMN9xPt2k1Lcx
kq3gRJP4lg4N/SBhGbJbj5LkklyGQq5LPP6sLfP6iQEaXLkLjuM4Y5jpn7/Tsj8K
GgGNMsR+ZS7D6c6RBMagjf0RD3DGa0Rp99isxJq+zkz3Oj6o9yCc+azshu5nV6Cu
WHHNiR/HvXFCN1KazT18uA==
`protect END_PROTECTED
