`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bjCfyRwew3Z9WuGbHrx6ZEc8Yr3Q/tWoadkrhgA0qBere7db8PsIK4YKKhG8CFfx
UMeggG0Qd/jo1yJi/0RynjsVtbvAXqy9nS/YKvfAaonaUFP+sRWMhMy5ofTjsoYJ
QHru2dWSj92guedlgYx5fE94sR6mMMRr48Aid4QxbnUblNqcnvXv8XrE4MfWxslU
6qc6ErhfwHxfwGtLbCvZwe/wp16oT/gsBhnIwUC5mFsmjErEKLMPf8FwXxTgmfN9
OQ1uMJgGF6MRfgcpZ9nAps+2EhX+OraqNNDZK+Bq9KWTA8av/wfX6rBwL7KSWiQO
3MX+H6QnMARYNTOaHTLh3MhNQPrW7wkZEIgBVd1TiJ0QjM4vTW28X1NPuXR9NrW2
y3wf5m+a+9UrVXs0MQKAhLmphyxXgt39NYLkIQc5M4/ZxXUThs3mcc/Hp9EJo+KT
ucWANB0SmbDxYxkkk75HWsm0XdsFiVJVXO+ElBW+O58PYTB6NJhbycgPOdlkOWEf
0dIxk/UamFpRApUkvmN3AhyEdJktDuOrIHOdBdmQiUTeAsX456fznhbjAYAAz/v5
FnL6OlVyWd6CFo8CpKJm3BqK9UOMa07xarmoH9dhoI/P8vihS8QeQ6PN0kdGsh2P
PpKh8nE6Mee+bmiDIdetiX1iGEneOfEJkjcWxhE9Lut+ImRZvTcWU2TESBh80Fz6
cCdcvvgZdn6+oVqsEh986xEQLb13frt9sIC6GYCrQYKqGwjYV5YphwgKb+wL7wXs
gMFXsYCmLdrMUUk1j9ZOjFMkbSvTlPplCHnzdMhnkJADsysaDPYgmTFb7g1pCJn4
A0bNdr7VgnSjS4wdTY/WgJgAFljpsfTwmopVWNKaEgxcSmF0/CSHHjna9opmAtgF
MTmkxcHFJ/C087MxE7D/UQX/b38s6xu7DkbRBU7hkS28EkeiD9Y6wv4hx473LL65
T24mQwlrvsHlmvq1ME3kZBrwhtm6cGQG0bh1sKqyZsE1Imm7Jl8CDNvorqm74prr
PKLURPT/mxfze5sX1B4qCJf2ruZ5CIrF/SAJr+S5CYO9qtv0mwieWSRsSP6G151Q
+i3VOA/IhpGsK9h/BkFsuJBQAsDd6ysFvFFA9Ir2KN+WzJxOKgst4hoO0VZllJtC
04j8JpofwSN0oWIZcXG0k241eaXs02qOevXcMg6KAhEM9LdFTSAKVkA2FzLJ4exz
8jnar2NR1riS0BwCS62ZgtZHWgNwNPdzHSuK5+7tGMiQDuX4BtVz83vMA3THPsMn
`protect END_PROTECTED
