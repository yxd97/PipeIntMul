`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J9JVdN9c7deOW4R7yb6qbNTOqyMDQ/umj0thqaWFiEflS2Szez0EOAF/0MUu8N3b
+gWKOLxn/xJX3Tls0u3awr3D54RCnuBt5HD/GoCAuUr9azgsbLLLEGrNcydA8leA
17eITehY3KQ78G+44rC6bHlYHncfYHFegpYJwDPUq/ppBe6RmoU+pA2kbNtcnYcm
pZgRR36hPhHiNm7xU2Ic62sB8hAHmZovR5QRTaZFDVKvYDhvhv8IJXlz78FI3gNE
gc5Kq3WYpi54Uqh/bMHxGeqJKz2jcBS+jjaq5IVz53HL5fis9xKZOH5IMdAwsLc/
k1xiSo+ZAhRXN1MqGWHjHF6s0wfHLVNT4Fjmt0SrqtT1iZu//IML706991yANhLl
DU1C3FX0yhrD+zMpOKdIsy2ueHAvfGUZqC28L2+/UtmCnvYLnxoO4HZ9MGDS1OF+
7XNeXxDclQx7QDiQeeYqX3loieCaa9d0XdsXUDez1hYk98GsrSSTJt+0B7NQtJZ8
bnjHkQ1XvRCnFTZdsCZ7J6IEZ8ShwM9XSZY2g2D8vg7s9J55r4oaSQdilxC8Na9M
3ghR78UxMNYOT4To0ksDtEsX0R0++7Ilk81tZKWWwve2nQ12kztGvk74Lpe8Nru8
1w7Zg+yKHzWEVtfP3/8hGCCHQyPnB33tcD1RXkDVCCOlLQu7PBY9Gb0l4cOjcWpg
b7KruNAg5mun+OIg1c8o4Iz2fE3811uoRR+tq1K0AWjlzWgVLF7ZUri2m7OljDXq
0xJa4aK+dF3bneAjIYFZmbmcuKcHGvHr0Iprq4zEcL8/BHvICR/2sYilGzFINPcZ
ApBBxTlT6u9b12dcAcLt8e2JH6SxfUArmtPN7culncQQ4Uf90+dD1DkHJ7AcWBEh
70z8JB98qKZe0MP2BHRmYP8zc/vBHu2RoRVuocj9EROf+HK1gCXvN/SQQhNibq6o
C7gczZVaJ5od18uykwkVkIbPj3tgvIXFNgGa0hS6P+w=
`protect END_PROTECTED
