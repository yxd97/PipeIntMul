`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnCL7Tm8lyCQAD+kyW4GSmmCRPVzUtY0ApWFLoZM1P4HByUrLAnDRwO+gD6zNxKq
VEfAFTOMBnULiRS0NIcYL1GNL0IKQijRce0uPEHvssVSY5BjST/7nnweEGfq5xEr
rA5jFp2nGunY2k7dK53ZZSpyVLz+9EIYezkgbHH0ceZGjVkuEs7414VOgh02XGBD
sBMYRoiH281NGPwtV0ONVCLNOxEkiPt9f6cY7W2OrapLBGdBGXPDBrXc9AsuARyz
m1IWsPyZo1n/OwbTnPoF35CfAi9+nsFvTaArsjFMUN8B3HOa6jFtUm4TDDJ1TPxf
Jr8c439WRWgh0UJ4ak6bue33nQV+fyHOlLLQDahWOXyVQ2J4Bf7qVW2YqjnUkkoG
nSM/TcpwJtGqJRIcq5a5GlgecsNzWgt8WoGsAJWYQ/6eueLqCG/nrsYhDn64TXgT
PERoxeiDkagOZdLcJis7fQI2JOEG3Fmzk2XlHhO7CsOVQUcU04T2a/ZYxJZIt7Ox
59wjcOvGSTcSypone6cyDbbHy7JN6+x6G4IL67F/uaU87wY3lbdDNMeE1TMX41aI
`protect END_PROTECTED
