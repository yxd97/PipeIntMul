`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIbadyH46Spk29QUt8Rd2WgRoX5LT5cXSehcWkcynp/CstwiIA4VUottFY3ATGpP
Rs9WCRlVBST/1C4LrtNwnUxGURwFgcCgGcKzHPU8UOYnqIRh7tTrm9gQMa0dA0zJ
nmtAAwdBGhmEt1wTZbNcCBMxOeiNhKXLHTwDIO0jHsVJh4M9Kg1QkEyj1DGQ9MnY
t2gQMcWoWlHYsZWqVM9DEiN8W0y1vvB/TREoVgNP20urukBSiFzEpimx9M+TjIVV
FpHnMAdX+v4CvjA0TRRioj6Tt432Hmm6otQZnoJgEIwoBKXCWmUshAespewaYPew
FVB/3JlSevmnV7B0xOEMvf2p8mjEhqgsMOgFiIhwvU2nxaL3VFTvtWJQVgA3bmTw
3rbLHcIbyezNl1lkVaSqHM0v9qSavbhrv3SeD4adkXRh7ghcfUda17tBWoccjPYu
`protect END_PROTECTED
