`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9IHLU7TYZZ/KHqJ3YQOzNaaSs/0dsaTRM9KGxUHIK6itUIQs3YLslV4JTL2o2Zt
D1XAos0uyHxCLfJn2lAOPsKNCiJh82PSSALIimKwxHsCClqaKTiPQv/AR4Dq1hpl
L4S/Ue4WZCt5NGjWD0tGwVQnD2m68hM8xtwZOvAlHmoUqGW7vKV1387sO3GHyzRz
m+IzflkkUowuyBa/pPJ+vPW4IhAVyz8uvTKMoRkyBJi2rBiw5kt5IhocqogeYaVE
B0BHqQRWQNYfIwNQLQhfErBz0EbQW7TQdrqHDRZRtC/ai8gmjRb06ECF6+Q9CVpz
ePbqnM8vBtY4siwK/47XjLk8230NcxgB+zvmgwBokmw7ulV07IpT2Wv8+6BWlrqD
R9YTRwUfWmdx3fwJ0Sro6XSmGvW4stxThgFjap9xly1YeMlalanWSSv8SPRv7Zgi
hl9GgkJzSMy4eTda2hef2vrVoV2ktDZzfYW3yFv5CWaFvLWtl+FA3kCAtr+Vs5lR
sHVar7qQjsOHUCtRLC8ORlvVM6Jl/yofzJ44yoU9gUl6opM3SKr9ZsrFVND0i/5c
NwEui075TO2eJPkxXVlCZq/sfYolH5fghe2Er8QxFMqMCx7btIMUp5+DxNMq46LC
buql2UY0WdAzkX2o640LQrDBTibvv9CVzL/OYUVTUmcjF1MoVapOhStXab0jxWI0
9Iv0u7cRwasP/GOE5w+e3Gi4APW+EK2TqlhXdjEHYKDXlwZmspvh95s7kSGvGgsC
lOrMN/aQ6qzm8XAZeuUwInjleaoHMST4/i9kfE345Sl2ek4NTQjrt6yTLtFzV3YK
AGt20zLCAuRyQ3ZZRaWaZV8oeDTdYo4EGJYV31Q+f7yFZN/wJiHRdd2FWq6Hc3Z6
ayw6w+Mw12YBBh00LWkdAppZVimaDzpcyfUZUhYvMLCV1pUNFAaaezlU0niyTdaM
F7KFSU2492UwppjQfr9yKlK2eE9mAtyIldZzcYyAC5fqnY7pzDWdXEwQjVcz3e+B
6KuoKHLRXFAYESDC+cmkkA==
`protect END_PROTECTED
