`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JdnWa06ayOLMDj8xWpp7hXDOCm1ZJXN+VUt3foVpwZ+OycME/eRL64MEYjW8lC+l
6JzkCzdS8MVqfuOsWp90Nj2xzHfQtoAOaKpzu+cOEeGuT1r651ou9HyRXP1mbEl2
RHMOK7tTTU2ZLJiO9mZizYZnQUrxtxeIPdEe17mcv6yvp6Jl6XPZcsEYOKqn+sXT
0duOrqHBY5+Dt27UQS9C7fgnWfsfekUOl7UY8hKr8iqoBI2yt+okP7C83PINQqWo
990AXvvH9ABfYlJ89uEEqMeOfVhO37luuwah+aVxllCTza+oyImS1wrGc/vvnjc2
ctdqvXKg3I56J1oQP5Gr/Yog1QHI4PageScbOWUodvk0ad1KsSWyTX5pKhGsfLgH
dNsVP8g9TpZHxAWY4/5GfIH4Gg5OjF9s6W+U7+k34XCzRhfxDChCBPK0BihAe/8n
xoP/psrILh7xgUaXjPflhwWZZ14vit8tcTPhZJDauVtj7rM71yHAjVRpWxkGLnkZ
VLdOo+IhrzP6rSoNTsSgeycJYRsPCP+jJvr93Cn7uBoXvJYBVQpFrH5lxvOw4lIL
EAFHawFiqCpjIX19ukX6GmGrEKIWMvM8Tm6ZZ3diLA0+wCf2aSgdzRgBvoVCfBlR
IXJRO8R+jN9ySvnAah/NfFAroI1Kc5xZfnOZzk7IHFqk8WWoKlLCIAhw97GRwU/M
EeroXwKRtKetjkN35uzFNYZoBiZB1umhNdwanow777EeLoM5p9QbIUBRR10c1kOC
n0EnExCWFjbXSnuD87Bz5yAnM3pQNKCl6IxzwErADpIhxOLSNA/L/TAHm5MGsZ0a
AC/1uh6rRizKt0l6YGQ5kFdcX5PVf9b4ezCA419yQEn0w2QHqHWk7yjBbks5LfUs
Bg7KHr0YEejUtswypIytxAYmKTj+ioxVBLGybyV4vzViEJu7fuv/O2MtMySmxnCo
PRKbTpqsMDuPakKGFdXFKsQujlb0jbda8snOp5t0gxgu9S19WKY7NxOhXzpFTUmG
/lHH0zJ20hUM036Y6zo0CPysVftdnmO/Wd6FnfBxDMYIpWdZOoSxdTcYPvrCA80b
Q+t7LGQKt4449urzIfICdjUyKKvJqCYkGY6efofU8W88ZKXSI/k0J5/tJTvFaAsA
f+GtO+o3Zrq5rEYqfrgsYyOAqUD/JAJBGsxDCsVVLDt4IUKCj2kcGAQjwmkKussc
cBISrCetApEmVDkcVuPGxXPWgvWcpdZRHNRSFCxMQrLSu/6GdQd88dhCIRUrgBMS
NNhD/qCshZd7g03znyslIlUo0HkTidxksu+AO3olYYMLT8Zy0b6rrxYcXiRrMsQn
8dFzWU0/4C6VSvtBLnRjiRgnPoEXk+WY88g1vGlqHDzRjqXiUD3obDBzx5ywtqoU
VHdXxHTSfx6yjl0Nb9BjHXQZeMGYTAjuwYBcmYEcGlW9tQKau2ccboYsG5YZ214U
7pG5f1gKq8ddZIsgYLUipAdNlKW9+zN5oq0QaCZPqoQ=
`protect END_PROTECTED
