`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wkoreZiBhBAnVZriXN5Bz6UTKePDqo7FcCUIlKUYMPdFv07+43V0UY/gWDg+V9FP
C4VGXRb5AVZx+JJ7djgA0GVKmJWObO/aJhhX0M/R2dZu1TxGERrpShyAnLzoLhnI
59G1w+5Hj+O2spICPZVlz9Riv4UBaGXFVMMukimuAxR1feMSZ5vGimPcjaiDxXm9
1gUULtJ1zppKx4qpmQA8vPYArxk7lIJMZWpGAjjbF1gsB6zXnEg10P03GKEWRyxY
c1hzAbV846GAYm8BxXKJMA==
`protect END_PROTECTED
