`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jbEiQUs3ieWmiVRAbqEMM8/aMErQ17r1TnyyjoImab0rWLh0w4d8TZcNkmw8QEtv
bQ/RtVWY6ITzc2K83LGjzsYCcJoh/UVDebECyvDGXYKx6aJfAEOYpVbwWYujnc6M
0fJ8KMHlgYS4XDDqoD8BHdghJly5njgZkM4tKOcfoaUR1jraCxuEqjusUPb781sS
NXN1vJLAcScz4LgjgJfnlhvX9rDKOTWSEiioxZdVbWGFHQfcuzEtUKCbxEN+AVpz
cxglT4q1k0eA81WxOzBnbQm03bYhy75MaINnUuLJSn5Xa+aF8NTGgdHd+22AbDIU
BCd4/FgK5vESnwPNUS/aZkdreuOwCgpwCf9WWX8/tvZ/ZiTAVH7bxQ82XUvVqUrH
+lt1HFLSNeTxEvA1xgoa4mRTBxHNzwPYkSvImMxBvRI577aUkTZw/KXIkXp1PqS0
1TJfBsZADpifLViYyhuUpnArxxm0NDH3hlEuc7+NZQXROt9xmVHsUZVNNVAy/IzK
00HLJn5mf409Q+AzWvlSliPsbD2FB9XPYNMqlyTELeyGz4UqjiANkdnx5GJCQzHZ
88lR4PKn7FsPOc9LltXixD8l1UC3ydI27sncfRfAd3EWCEgaXIXyRpmwQ9G8Zy2D
J6YG9rzdwoL2ucoe+zZwqfkgl0+z7kh9D4mfKtR2GKwr9hXUKGw/PgEbkyhmSJdQ
S6cS31ReziY38Z3wMUVxyj6I3+bFkN4nAocbx42sThgcTPzoqXUMC0nR3wg8cob3
ppPpg3YSFUny+Cx9BAtwQHyQOcVkwdsnlQCLiMhlCjfoSa3OcRahRbTWrFe3ex1J
jtKbzQFPKb60uZjSPSJ6rkaGphskS4dkM+cpb3P/CNnfuR+jOt0DGoriWnFF3ZbC
5lOOHOm0DOz34eSiR+7qLIohUi9AwLuBQc7+XlAVbpnUdbWu94/KIvJ21cOPTb1k
ILfxGpPhwmRkkoh3lOfJW9ugVeBdzTbiB2DTxCz9N15Jy9BjY/EgwS1JYQBOkh4u
YFD5G/UFjZ0kBfZX/+6lTZgIloGfwu6gE8nthxGDeLv6Wb80U94uUr+AV7S8PuJp
CRIY9Li1LF/dC9s8+2/lEKKqMu7mClF9cLNRpO6+H6sFqJCxGpQnfmfmsDaJe4DL
uYklrZJGx17eGeVYF30VVb41Rx/MJg5qDO0G7u++O5tC3azyg7DarvRiKq+irGrh
f1bpfKvYtXZiExMk8vV99A==
`protect END_PROTECTED
