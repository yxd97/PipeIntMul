`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QetSNxJe4+cf9v1YrvGjH/680tLtKmb00eEjOuX8fj4d0LDz82wd7wQem8a8b0wf
Cx8ikLB2iNtsX5/Y7BN/KBaZTRKSt+ztMdppkUky4Renju88tF5tRZIKLRwdxf5l
lBo15Ed7o6C5omN9KCQMg+YNy9tSQ6MOMGHSSn34W+fDF3/AY15b5FklcDluGcwN
8tu2HhO0JrcAcWxEPu43XWjOa95yRdqTSYWj3B+xnCF2AYeFoXodU/otcC5uaTCB
Ov+UWbdPOKZJr7f10CrFHRbRhbLMj20DC+7Mr2Nz5QGl2DIPcOWLMfS/VcEdmDyK
fLznySfxnWiGlxW/ptbw+UviQkgCl6aF5BQPjq/PPWMb+AxeylK96I/8seeaTJj0
LbjLafbOZPTH6jWr7PGmQDsfiJb+JJEQi0RPQVguVP6eyvVdd5eZRqoa8A2ePBJi
EE86YXJqDfZD+HxMvXlrlkEj82CXij8OogAiRTB0HgxB55BTB4gEkR1zcmbNmcwB
EoyWw560LkiT2ksrsddE1QK+4mZwkfAclx114y87g+W27X5yt1EKmsLd97lf3nFy
zLBLtkRTFyelVRoBCcFfITvbfnH1DwAmcDYqbWQ+vhsXBYMMp5MnGZLiueRXxWl8
O5sKxtMOQem8ZESL5yiL9BdKWYLP5JmfcIi7Ew4VYAd8uHm4e4qVsG3nG/jwuJWs
hHg1gzHUCAvmkYsykiYRcbcx0183adMap4ZIVhoOtag8fDRRbG0nKDGmiCvSPXLj
jDMnfGKo1RHQmmEum/7EwLykvEr8PgCeW1l/x1LqQm18HxqXLacUpdY1wha8hwy8
KlMuwU0m0DxFpN7og80xaaECSjP9rHowIriJgR7QIvWsIyjPf/peQ+1gEnKwhYKO
5bQ5sSgy8Cxsh+ldhoMS50pNYFTW90c0qtNzI2peF5WdOt8/fqIFkUMfMBTqwPhQ
/VDmbGQNijdGPxIJojOQ3ao/C8E4CERY5fdTW7C7xZ9StVaOveODIP/VgvBn+Egs
fCl0Pbwt3yAlhBBav8mqW+HxUTlRkiPe+vrdGBBWtc/eAfMnRsxVgJk7rkxNoiak
1IonO8Hcn3ok6oVMnPEWBfbnTAWky5iveZkQSS1F7qz43dW0QzIJ/R8v+iGBVUy/
hMKcdaUjhds3cAdGRkf7fYGTqGkoRIZtALJyVsSk+tHWx5JA04PeABC5e0dmeZga
/RGFFqFCCJUsZX6LD3q9Dr+dCWgjr0RCENCNyiRoeucq8D2fIte2YthUsX3qCOFY
mij/z+/1aFgOXNIcH2KYHSVvfXVKSn2K/mQ7BbjNzkLJTHQ1ackH1J/5BxfubNK5
Ki38+Lqq8mfuSGpwlW0KcvDoWOWfxvbXEVvP/teFHonLhv3KcXvniEZ/bnTdB6LT
dP6ACLmmuLptFvUmkXM9JIXOaZ0aQnOkKlBsBb5ip6/Ppvv/ycDXqJ/p+3ZiZMBL
5Kr2Sgew1N9cvilrml2CLZATjgzsUEfXkMhkcYzjEShAPuzaSq0UqqvyIkLLkhGW
NBNvB0elas7YKCp01q81WsBxshqwuCc9lY4Id6TfdDBe6bdG2FRuO5DZ2/ylJ9v8
vLTO9I28Sy16T0fYoFti68lhYJxjL8uI+HcbeVdiJXekQJxVlAy2CAqphxfkCXO2
f148KO4zuiaNC1afCbJdLSbSTcIimAYgl1FrtlpPHV3YCL4Qaifg/p6hdc3Wxxpy
ML5yCcp9OvkrvFe3rPiyM946ASjpW/S3iS53ROZeUvI=
`protect END_PROTECTED
