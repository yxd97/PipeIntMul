`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NT8YoRNgIxqTw4DrkvvRJVwdrx5qxMAqXjJk/AwT7OszqALmeuEIr5nJ9tjjSV7i
ltgMVIuKPH477/FLpTWb4uSFjOl9Nb4rz4u9RVWZ+Y5BBY2yjST+lFDfVw6BzN2w
14Gz8sLNf7hIkS3HwUyLfarV20Pkf2hCowx+5a/Ty4zcVmrVQ44IHCrK0z3qu6Wt
xOwsYPq+yBHej3+36QPJfMdqk2AV333ZIMm+sZgbeGKtQAlbqbWHe7g2XJnJJdp0
Swg31f2IWYAXDw4pXEsn128iW1IGezBCVgTxt4ndGY1r95GqavHse8pNy9SC8U9W
13UyEClTyt1XRciwpMDc4Sb3hwoW4t+tF/O4jCg2fi1rR8K3pbgHje9uyG0kKCwA
lnqLXwCtsZEDTQYvqZkyx4XVXXH6OxXoiXRCTevX2NjYsRyHPu95iVBpj8wnmDvg
B1o950KJCqA/H/F3ebZZ88qvt6szfncWDyOzYIGdaIbN+p+i35DRMrN8S9acqMNI
`protect END_PROTECTED
