`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYtQ2ScAyuop4q9cz7ve+0FtPgNctTPGfh+Kf7cqo+vEy2kFK1JhBA+V0YPqCzDy
Q25EwhkaTypNPkyRcwsIRcKKenkXvJxx5JpadgCL78LbFqR4rBBBzPo0+lpjSu2i
t7/Q4KF0G2ceKSi8grdx+wVoCdsW5UqU22afZp9nHdS02TWQ8mzXQFACIXlw6JtY
bujh7pJRrTqZOwo7xTEuW/zwL/qtpNzLyfXsYJ+L72IOR56dcf2OwsromqGCM5xD
4DxY2wuifgu3WGLH+u78lZ4wx1vf5/JJFLAbKISc9Ccqz8yEhzu4a5jA9dixGOaY
Qoh3YsqsMx5RPoxNsXug7g==
`protect END_PROTECTED
