`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bvdn1T4pLu+dpvdZ5SYX5UsuXZQsmHP2Sw8w+T5+5m/s0AJc72EhvyXCaa89fg3K
ZLhBBObXO+8Id0rYM7uNbsyv9IPRuIei3GqjwJ7dgmSPXulgZvQ3cNRh9kneUPDW
zn5z0zn3+UfbDF2R4pGOQyMOfcJwyA24ymvtqL4djhjJyRBMXHTRkIaCFGoj/8HD
NEeua32ps4wR5He2SIOxNi+8kOPkG0mmziKK5XFgacQKsoW8B6tr1vduhpGb5tfE
n0VbN3DxTSemYDLEtVBpZaQRQLepp3BvajGKiuZbhmQ=
`protect END_PROTECTED
