`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tKOr6KiQLcxw19XibFbzFyBzqBOM2Gr7ERo+/gXieqF9Q1e6OkdM39oItssonEsL
ua/z+6jOKUSNT/gmKzfh+DE0zslNLnBP5RhLM/yguyJ0VhjEveFsmcKmgoao5bEq
2Kxfi4GunEcP6rB0Lsm2Iuk7iQz/NF00GkAch3Xux/Il8H2V3eBKtAB89hDOp7RD
7nzDXP65Xwh1YwtpqFUERTbPop4w70e+3vIItZ8YGTudPM13ifqnuKJ6tjJJqolh
CP2foDskT9RnsfTF+AypvKfKw5e9AJFY3WdWiRXtLc3fngv4X/kp6Jcx3bavYTDI
m0JtDYbg0kRhYOTv3c5VQUlZsfBr5+H+Xvd3Jn09Gi+5qLazglzbWXuXqaVn8DBS
4NeiEgOjfoksIKZcIJq09+pf6ppvF7C8fvOc9BX0OUznd3jlvpw/c8+bgn5uufw4
7xinY0xVy+vF4xJQJqvmEwpE7ffwXmasOg0AG1ikeRx8nauBKHDzQtjYKSAESZoa
b2mwa4vqWEpEAUM14UNG8IYs0xOsPhhb7plDrdVwydLO6qYfvoCqdEKdnls0drV2
UM89zIQ++gkxsdwmxQPBd0RPGMTKvGq7Z+nRibvEZl7ajwll1SwS4MmCASe037tJ
Cspyj6M6lKJL2KnimmyZGRQ+L4oPH+3X/wBr4xS4Q5+FVrZqrQPLmBAsPuLDDhH+
0Ue5CJqhjepwmsG2ttoyf2vSgdTtfVOJRfec5cB2cnNm3k6kA7kPHBb1j+v488g3
3XyesQX3ojLTHOha3oJFn/q1PE2aeL7wdPK+I1mhxVMVgMlfcnO+VlBD4++v+hOr
xTMsnW/rSdw2lNcnKHBAE5up/zUeoU8tPUZYixiXxcrOgcXf4bD+WlU5VJ8kvjAt
JGbQbgscqayKAOFd8HTv1hRVN3mz2jSpf5U4yrrRVcxti9o23DZYyHNFRz/JeYd9
31F4/8jPQCxwgNKEiFBLZRgLWTmHDESRoAmUVtSzvMqalsc+UqWN79stLkCCdmG1
LRmtDp/SCfwmmxhhYzkd3WnIRGClrkU01AkPSi6ETMoIJUN4Ex7YUZ+YppO8rd90
lS0vbGt1N1woUq7xpzd5VhqdZrgAfzCnhiJ1kHCrQVqquaS3EJoZxOr6MpFrj0Iy
+i5ZirlmMqQV3sKdnGoiiEHYXth0Eu31eHWd1obbOZHdVzE5OHXxf3F9qhsXfaNL
SCxSbveX2iQVjMWk960nNLG1bcwTUOjkFn/n0vvpdIu+wgEug5C2d4MBpKCJG4RJ
AgZXYwq3S9Ai0vh2rC5rJRqB+tjqmuMCeLEZ9/TyiQ9CSzc4giJZsL35CbrfNZc4
yCNhYL12RHI127sWoexeGxbR3uKv8u0rEwZXyMvrKLWg/Hg/CQdxzGyBdXbHSJpc
w0a9bRCVFRusD0yEr1b87cHPeHxNRUfJZXswNFq3CoD75tVB89se5wnJR0cWbs07
DD0bxDrJCs1RkNTQAXpB1OEnFus76E+SLuJsWOZbRrGf/FED7QqqGDfJCl25XgXj
9FhLJeg0t2PA8Q5A77iyijcUv2SdYMVDKVCp4fmX5yQl/muPAx372XoF5w2ERkYr
0T0YDqjXIkyVJ/1IOU04BTQEZm0qcoWKUHjr8m/CSDIfHgvx6V42PxwM3LiYtvo7
d2pUPQJQY+scuLhuiXZgDhICFCngCPuf1rsuSO7p7KNQKr3kfGvO1dNrE14zKApW
cwNj1YJDWlQFx4j6k/X9V7akIhuFYmFJqYixTqo2wFVqz1/1VLiYOoJm6Pzi1O5m
vAxAsEgCazhqUloluL4Srhz8XiHtb8MawqzjyH273yztm/lZCXszkIAfgC2o96zi
b6nLo1M8zl6hkAVpc4EM2ZenjslGNh09I2v6wAX4jWzhYJgM5Wi3ZCE+qDhuDNy+
FUx2NM0s2zckteNDLyngkJrYjbJefXNzJN/ayIQIv4p1KlNgDPpQ75DxWmvwbO5M
UFNXx+EclbRO8gZNQ1ZQqovjSgqmQp7cXv1mLe9d3AR6KXcKGMi0GZPqKo/XZUDY
nmoubNU/DfXQabzCZaB9fsIuYs4Ip6GgQMx4K2N+/KWu38Dz8khjqRVenFHwD981
jfccnLmFtEQicrGSYdCQ73VfvmTU2MY252ZNnHbzvA9+4YiesJnxspyr0QtncAZS
v/6iNvMCQ4yCaFeaNoRNkUeI5Md2okVs4ZXucy+K38Yhy/Pn5Q34ZEM+wrWPB3d7
emyJHblFI21PLWngB8gr2u69OmMQmHMfCoQfGMO9yQrdp+m/MFEs44bIFOsx+KWj
`protect END_PROTECTED
