`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9p2HHDaOmWmElsRi7a6R7QrdXA3D/J0wFOFMC+QS0o3mJP78nGVmcw97kIiyUtBu
UD32uoTmfRlyFi5QCgOFf/WBLbpmkABTPfROsAAry8j0fnkYCxVwxnXXX9IRXa7H
B3h/IbjZl8q+dfJPl6IyBfzLY1iHQ2OkN2/ABDaV8Zg9920YfrAv7bj7GSPu+67B
g94HJ5nQFpO0vDC3Hc46KBgcE8pWLT2hPWi/iZXrsfTxor+Mg49kMNh4d2sSyv5D
dw6e5mwXorsHTFEfr4TD0/LhC1c/f2RZy9fBtcxDLCHZ03ZEiUenOrG81MOr/Hzc
Pyi2BsecMpETLKIKoTWHWQpBtqRTnFqW0prSrE2obuaG114a62pU55az84rSKekl
CEGHZiHV2cZ8mx1TY/dso6c2r7F+PEqmDGf0CYRVNPV0bGZl/ql1aKjYgsO52G9r
UDEYWHQbbAWUlD9YYilIs6VhgmQIubI2t9q6/tJGhxNqKqWnquKUEmMl9gBXqXRM
z2hnpZ/GfMQjjWwbX30X/8Bm1RwyyZOGv4CBIDSFadVad2vIQdYZfyl5tFYCpmpQ
eX9LsH+W/Kw3jwY5I0iKCeFaS3BXStYluG3MG5VdUKU=
`protect END_PROTECTED
