`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5iF8WiTDKAZx+s9xT9p4SS4oMe53jZWEP+2eFkz2EfQ4sEo9og8MLlrS0WHvKqO1
l9g8sBRx4ZP4ImluIWQxB8egKRB7DoaZacHhn82TgCW79lgvG0Moh7FQLkJ4BOAN
GugrTMJs7iYKPj+i0LQOV2S37cvRbKCq3aR98mEkajWGCs33HE+jNLsgALmRiHKj
nBODEfRHeaGX2Sx8rPu0WGkl7fEX15FCuutRBPfvdy9rEKCs8l8oxiYUeEwH58qs
6p5G7roqe4gFiCJu9W5BZgb0BtKp7ZlmFAsepsS6GbJd2n+kBUSCz2W+GMEBR45B
rODqkLSWgQx+wIBDsTR+E/VnZpcNyAnWiyVhx0IS1s5e1+J60DRLPcCVGoXBuIu0
zEv+Sngt/0HDnA3k2w9ZOqaqBTD2ev8zo4Ll/5PS+2dPCHVDiJhfuSeKb8Zqp+rG
vA8T1Rb4wKpclTj0Az0cq9gOILtHajtrmUOrcwEeVXjQrHCIBAWVSqYWOruC1Qar
Bk30tWlcUFb85gsk0LXmxDis1NGMufde7Q5FMgs73n3SGjQAmaq1DN24v4tCue0b
w+hUdgu9DDzQuQ71NtFb0fMniHrwELv722GxVNcF1PuB41ZHr5hy/vcXaS3vDzPc
MnquJ56skyKtObm45B0QXWvEOlsKxZUumdWIepEaX7kvsFvciZmRISFVtHcwPnbq
sPnxAiX0EGROOBpv1i3aPBKzQQ1m1MWMzbf+tVfg/dBEGuLtIPt1pVwx+JwiiC72
cubpaBS/pWzMFU9TxrKiGhSdTj4U0MPXV2zyuFYkzy/pv2/4TBf3dcrJksSk9n9w
6Q19AwfXeo7f4qOsNuq+FUvELKlmODSWf2pdJ5mhNOLaLsyIjFO0HNXv1q64tYnf
YqxCEtYZYSInawVUWwch24zv+7r/bw17UJTv3XmE88VIhizTbcf8WVpKBAiPLXQO
r6b+3fVvDD5hgBKP9G9ti6GB3RFVFm2CPelUBjOj8uomRzpZs3TXLof5UyuEAgF5
/HmxNa9/Wb6KAXVZmVVuTT/lylCwM7hA6L3JxZNsW66OV9R9Wz3xun1JieKMny2N
RFT9Hb+ZYQtZgXfmPoNJyLcHEdKrfj3PaeW8u1jx45bJC6+ngvCwJmqfKxVZCbAq
WqmxkNQMsvOVmnXB13GPFbmrHaNkqXC1kP+wWO+47mnpbShwaX8ZewY4LhuPoWlb
BsCi90g/qb0NpyPNhbQsX5Ahw14hlxij4vEfRirJlg2DxJ6elt43/24ueo4fwl5A
vlI3l1NrfmU9Z+kMkmOZdJKCJav44FgIwFzRJk6+rVzfRWdFM182zQusNLdu4bEK
tKjMtr2/YbklcXz0SC8/mUQm62Yo0VHVlhHZctFmtbrJ4Eggp07srQL5Hc5CIICN
CUn/lsl3hqQuiNV9hts97koFvZ0EcH0mW0MzxKpPQCapIhFqf/lyiZzl9HbjgYcb
g0nbf6D9M9Qw36iDKftpsajtS1eBklwHcT3/J7labQx0WW/pcXTPHhNckd+cqVFX
+etotHBHdQUx6/xbJ422FMBUtzjx+oA6EB8lnXaKF98e1vMN+6F9o8UIBeXRg5qO
7WbNlYDB70+8nOluRN8tOjxytYuXYcjci9+14ZaxBdFm/2UuhUv0sQFceZHg8Egs
MlndL8Cj7BdsPyJTJd755UJ9dWbmQ/NgI5QHMjvmDdxuGj+/FkecsBaB3mtntIuE
QO4lOuXK1PBYA3SKiF6riXaD7QRNuA9RTHglapVO8TccyUe1r3zKhapHgEtGMsoE
eFfZj5BBR/X1k46KJ3BcUaaSghOT8Ned36RgmPeQK/E89R8hjycF2J9YcPc8RFSF
0zQ6MoJGgnAWj5PMa8M3tUk8eovLYmchR6Ve0pPzuV9DwN59VIWLX9d1RDW3v67Y
J2To815mAFkHxGuki14FaJwF5MiYmpQ5mo4WIN52+UwXshhf0RP0ARzfgyGYrlQy
HqpWSp/qFsR+e16lEPiGEEJTpJAmphKCkEykZlPGIYzpou/iw1lSlZ0mKVuLOOYe
km/i4aV4Dnn2q/ZRWvxW89Y+Q1upjkPtrnx9ef8rsYQ=
`protect END_PROTECTED
