`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y54RV6Pf/Ffmz3GF8WDM86ef6jQbk/g+Xt5aTw/cTQwIe7mYfRCRh9VHK+jnt404
AxaEMYsvg11Tkw4Dg50tYjVo1nUUsISMYnqIZ07ZZBbyruT/e+BWSBjQxGHQYtNx
9ASpm/GHK6//lHTSHiOls4GCEbP2GDZCbxw4Msl68/TO55XwobZ4rUmaJXU55uuP
p3HhbN7TzHjqavBb6rLIxFvp1JErDGu54wq9a4e7QF9nW7nBWRHab22LVcwjmy/E
nFe/2zuMi7/nwvUJpDx4lOfA3hgWFKsfjFJA3S66Et6l3HFoRF80mYSxAr3rMMam
zDp820BD6XJL03kl/7+2Cr92Dy+zFB2L/BwiWR98EfkXCjElS1xNjT8VMXWQLeAd
MepO83GNHLajMDfRHro4nuEmIFbKpcfAwR4JAHGFzNlxwL4/Xh5vFUtSfVdNdATF
3mGgkExAtoW+rn1Rv0H1sxcUgYPbaziDTC9+ITW2SYnnnemVrFCfIEY5sh2gEly0
/rHvAGaxQKHONoMP+4Rq9PIUU2/P0ITAZmruTI8t1nu3GYBOPCyBimiak+ckLjJP
INTaSbREAk9oyQaO3D+jBDzVociY4JX9wchk6B2ET6mAuay4kg5jA5e0IpMBhXxe
3DUKMel58/k8jcSjBKMznQ==
`protect END_PROTECTED
