`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
miljgeaNWoe+yP2lUEPEyK8HxCLKfqtRTlWPtY1dw5YrvZ0EWFBVjGt8KDCPWCv3
RRvFcVa1qE0LGObgjGKkzbEfLL9P1LzQZ1VFD0dFk/CtCmOjItUnmv9Iq8mEFaDb
FOk05E9qmiHvEijhWX4AXJ5Xmt4fP2+vscFr9nP7GWxSPwQ4sUuC6SC/V/7nuYZ/
e5yL+5o3OOYZiTg8VZLqZ9/ZjU8IDjEicRe/+rkwiAP147sP4u9kAa4axkEc1X4p
BPOH36FdtEsMu3Z88+tjdE4N4Dui7mdr1yrqe98h0uHtHb7kBj5VW+un95ob5PoK
S3v6ZMnnVgGIlF67R5I7wXfZGmfS2iUtt+uZx6f7fN9xlOl/iyC/Vny0tPI/CS8E
JnkXZzvhUMGzZYdVvco/4qezaKfHktZJGJnHro//ikt8zMg0j2BOJwTL1bUpJeGe
UnHZl5bCodX/UrfGC6fA+1eOTWjV4uxMdbuhFLPELPfBODdrCDgdLOOY3uq6OiLc
G69Y6RZKI2HgzLl8XEfFA6V0a9aed01uahFvqycCt9o=
`protect END_PROTECTED
