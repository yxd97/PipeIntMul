`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KdyaONnaNVS3MJC3bW5qT3j7WrcDWEntCm7wssnsqmnJ+uBAQf2Le2wf9xV0HiBQ
s/b1VcFgy8xzwh4KPMaFAhkdleHquYwlw4i9J8DbbaFtodO0/3xlqbD3ST4aKKei
RApvDkr4LjYZJJ6ecB1QRSSh4inGXur5XxGuj+29v9PxeDwFsFlwbCQyVJeE0aiu
uJcPLXTkcRzr2sfPsVLMyDBP/1GOrwdOsKBlMah/0YTdC5+yrrOGi1UaDTzTnOCK
mwCC46FK1xwsoi21t/on9BSw6+wI+iIp3eZ3nfpnm9vFtDtEyG0D4DdsZeOUS2pr
tB6ur4ZWYlthrCTTKhhfjP5MvAdteDTuQlCmzj2X4WJ6EIT/IWpR2HU1N4Ke2zjN
C1dzBERC0fiuf3+JTgXxRDoDUPgudm6N1lPYxc+fjtfkO8zb8vD2g00KAs8WgyZ0
4r1xUi83bE/eFDhtpzd3KjDYRS9rsHL/eWXXVS851+eQzFl5zj57exOpjLSvNl2P
ApRhIurX1l5BEUvIbFiyi9a/zmCynv5X29dCXHv+DKTkJKNr8RbNLhbfoirpp9NI
zPt4GGqGHpHliResIIeAr88TxJ/r0VsbMcbh+MNqfNp5a1w90ouooJqtVNP3eV6s
bShiHQMT6S8swfV2nctxrp7HIJbs86IaARUqc0ClSnIu6K307IKW4BsO+OKisS8b
M0n3swZlBZNdB7xMC8AlHiB7h4d3VQQcSlNV30MgoRIBlpKTLy4BPdVOicAzTtXA
XLsvuF8iVMY+hrMWQNsqmtClm02UJQ1TDSypur5FjeEHTiiktzj7jG+WBKf0lOoW
JNXDqiPZr8zOOVxQfLx91jsY3Sc2A2C07UDi2hdpwpQ3coEn8sUcc/r7bsvePnED
oViajYeCzhcW9txYuC/yU/CrExKPPEPO44/0toigMFMDgA3kiq1pVQNVBrUelEaC
p9SFlT/vYz5KwArAZRCUWQ==
`protect END_PROTECTED
