`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ntpQgzCKqBZmgur02a97RNaceYlLBHNCzrgnyruB6sX1Sv98hUQjOGNEXS0fcWF
13RJf5Zu5aJMPaZpopdVSHL8CmpL5ovfam0Xb7v7zaJg2KMtZMZ7uhbO3YnCxMy0
aTOqyFwrkiYiJDEUy3ppvg+fmkTX71mmmWPdlYTr5TzULGkwsKy4U4pHEsvLee9U
25RT8IufUBtqM/VRnd/LIByef1bB+2tR5LNwm3BciCNzevbTHjanAa8fwOowbpsJ
2ickdaw2P7ew6V8CgveMg1bwEhqvFucdEaQ7YpsDxdrGWYXE2GKDmDNS2R4P7iW0
tbB1w3biU+hRtAPYxcgMqTxeAiOkdNtxsKKIwRUFAckMM/gcs2/uG6QdJDsZu/fo
HIwoukb4hppDhMQHFqe7BWangQd6jQO6xDFZZK3xO/yJvdYhsQU9bGtPVFsavtfs
cRcwZuhBKGMzJc+kJag2QmetvPPdlVr6effgaxB8zTRS1ZVVLRrY8GsgbSRgKef+
q60WecBUk6GCsy6V3TMLxMM3Rzdvnkv/w2Uo0D9YIyxHut0iG4hxHLY8P/ALySX7
mSK8lmaY24kpkGsG9CXuf5z/M0y0dgStUVaJF5Vzig+JnR9mPdAvNf9RNgH0ieoL
46SJVu6w3EaTvEJAxqVD7siE9sJPqWvP2BfhbdKjtqjU1LclMzS4WoOWXJr+jpq0
pRLYtOF+tqvCT9qfpshGROSmejKbKbte6/j+2sDrDPM=
`protect END_PROTECTED
