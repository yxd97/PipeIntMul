`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzHU/gC7mG3IkYMKFn58yHvocH25KbXo3OhNyk+xXnwzBccLBpzUHpsc7+T7JDNP
RO2R+mIl+SQFXob8DBwB+0Ki4tU4/b21r+mIMcQ+Qjq/ea58WbxIKC0XQ3at4YE1
n/S+u1o/6Kuj6iMHZmcOdOvrWWJMOdUeTKTfRfKMEKsQW6NCL3ISQt7O74uwnxbA
OsB1OVsVUE/uxvqo3sGXKJT0X/FMqtrqwy+XAsybrEST1vzMC0HxeV/tIKuVdhPW
VbC3GHf13toqf8HzmgcJy+wM4t1BVMlORKH0ukTH6bkTF0jrZU4lvB02BLZ4W34V
9/fOhdanEe79+F1q8g4OlJq0t5tPQUI/x1ouBomoE0/Ot5QUdpR4ojB+LcPp5hh/
yAPKHESIJ0LGvqv4k5YF+Xe4kAOu9bK8WVvfKg4tRQwvgXAP6xuLPgmor4jKjyVf
CSZD9/uFjeeFokmVJPhDRhoKSu5plVtIroBj3Qz6AiZSvpe5q7zCPdO+JESrxIRP
g4TD+u3J74To2jy2yo4fI0qtrzq3Ci3n2mgYp3rNbN+xFUUb145PVHtdaWSUiNc7
dKxyKhvv3XQ2L7e5C52+DNDj2RvzFFw3ZF+YmT8dX1me+hzxd3FNUajZC46VxjQZ
`protect END_PROTECTED
