library verilog;
use verilog.vl_types.all;
entity IBUF_SSTL2_II is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUF_SSTL2_II;
