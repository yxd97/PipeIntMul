`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kx9wgHRHcMVp3NThp/KQ17RgFyu5hJnGs4ouE52JVyxd0hOu5Rzz9nZyYvhoRvnc
+6XfMoatPKuzzV1ojQXw2XWTUYu9qebOTUqOg6d/3vIy0KCkhzP63p3eaGEny0iX
kay2vizKJC+VUHD78MEYIc00Yp6JeLIICfIIo3OYb7/khFNRfUOnqqOCablwzUNZ
Z9idK2IYXfgbd35zQ4q1rSyrq4pU4HghmrIGeP8icAH+IBOlU0f+TpLWP0sAdDDF
LryXcAJ4Kz/iWsWvb9JRaEHQ+d1P5kYF/FX6HQiGbCQj3uS5DPfocfUowHw3V5y+
2SVIT5dvUxjkoRjBvV8M/xfBxkAIDF0Pijd3llQTUz4zRpNdcC7xSohRDvUC/Rbl
06bT9rEewNAUEgB1W0cUvey8sh5AdABumppXhOwv3ouGBkDOi5krCKs4qfZWfv3h
awcoND5JNE5mJk6iYepMcEY/SU5FgjtvVOeIpru+TqHH2mHTmtixZw71Gzq06U0k
6Yk+5p5sO6LC3sdKEtBvBT+bj0G1ly7lAhgk4nnY7l5eLsiEBKxaIGMQpq267ToQ
9UIfbeBpPQ5quqSPeiAd8zPRRikXBwpRFdtObn+3j1OgaZAKaLW61MhXWcdj7Fr9
EHgdz3S2VRlE8m1seS8aJg8RbsIc+qLAc2YVzc+pyI+18yUASrycslqw6/4hiJum
mKCZFUkxAh7zsEGyhrZ3tq2CbcaD4r8qO0q5awzEHApyc+6DFUTgyh1/46qI31/l
hkU7b2EzetOBYRRMArrt7p6EeM2CcspZreNUuTtc3Z+d2Pe6ajJVpli9sIGzq7FC
uVFH5GGT2ekceVp1ZQ74fKBp1d2ru/NWn/jMXW0ZTswFrcR+lYodQEIdVc/xZtb3
VHg/wV5OroiBUtZjqDD6etlUD5h6wfbo+Y9pWF7BkcjvysD9RzMXL7nZsoJVMzyW
tIyo9Nqx+Nl2aiBDguAyKvMbCBuMTDwyZvGH+6UNwQm6CmwjFawH/+S3DC3XK7Tn
Xq/OsBbnfDJYkgkiFqrWjY6LbQYkZVr6j01bI1YWKBVcrDL2zi3O0yjqlKXKTYOl
LJ5oao7rOWWvtv6sj4+nmubJuzrVKELCWKn8GkdV1z+WN/+x1TiDU2O+6P+zuxVe
dcyjENqR+8QVJNd8Fqp9A8s+1vqe8uM31e2Hlnsze1PIHGRUkc8fxjHaSDynLXht
+IwX4Q9HDYnvk5/ANQ2pKBSSBe/s5ZewqJeC/dcm1R6bMlzcCASczSfGvb8Zjc4J
mh8O9C1ST1ciFHp9/KTuzSDnTBFnEWY8J+DSmvQwxw2/F7YV9hh6eXuBH/qs9x/L
FXW6PIPfzzvdXuN6XBVi0FfqdDyi+vZZRXyElMeAIBvjC6y6onawYTmJ+Mt0A9/5
`protect END_PROTECTED
