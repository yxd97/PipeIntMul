`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4Rj9dSEWSutoNnVwf5T28c0PqMdLaMnEBQeXNq5NPm//4BxFJ0ls4kAoCuXZaZa
5ne3mKSel5/LDTRWPle+fynhb4cSFOJHEHcRbwfzOZvFSqXv7+NQmejyERp7KvPT
0569yFRPEK5KKi4V/+B92lj/3pSW58z+LkOm0I9ByqrNGchJjvFjz0Awyb9P1B2Y
q2/3rlrHAI5fkVQr3QIukmQ59khwrfxhNezMeybZM0fRrrBo9PPpbxiHoUJqDTsR
0Uibc+tu6h08C8NRX+XnVXNz8pqQtxipXVVbm5C+Ho5hmgWQc54bMOyaKYGIalUw
jqJyxLidtbEhaIlIJFRgwykK0xXTBcWkeTrqfmQTSQiwU1LiG87Kf6lx5jOuS3kq
nwBH3j9rG6pZAkLpbgnOAg==
`protect END_PROTECTED
