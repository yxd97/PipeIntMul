`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gz+Kb3fwZAgbd1cpqacBGqFIu+KlCyCO8bXNr9h6VHcT7JHPr8heD+r6nTQes75L
M4n1/eI7RrxmxqnHL8rDSc7il4rJz8MZTIjaeIx25Zt7k3TneJ2TlL7/L2I2MDFY
d0j8bWpqROSWBk6po4AhwU56OlHpH/ONEHzbQeR/8ZOEG5Y4YhVmGPFLJq39CSxn
9pMwgp+y7xl32b9O9qdFO58q0KsnMmlVKm1byJQhv3hJSFYaCGnb1G+yha77TKBF
qantLae3pyLlIHw2Dvkhgl+yyGagObyy9+q6kJEx+WMCex+VHa87MqyEJR2xa1op
3IOL5jZ4NlzHl+bhNIukr2baX+gdIV+aw8PsrcptNgOtiqjfQ3EOqrKylWIENzbz
aeOS48uB9Xz/09uVeZf1kgz6a6KdPtrMF9DVcvHh0ubBmhKqxscl+JX9Ni8CdvPK
it5um0OlAp9CfNI4JznC3KBmTNwthhLjKQ8zKQhLB8+NkEQQ/DvqExLEK6D6T3DR
cAHcDJ0vKFEdoxpafjT7ZcDSwQQJ/MivqiJbTEsaCFmBEvahYBxR0yb0b+2JgYvK
mKvmJT3AJlj26Tlps8cseryeYWG5r5a+SwfeTU5aV2F8QbSaAGV2zz8WYDNYZ9sG
fXHb0hzBioTlNRyZxBXYR9W6GVkbVV/2aLMU/Ab0EiJn7ogyuxWD4Ot97OlLK8op
RH6ISprrJmB7ajASOxBmPxdPvWPD0URP0bRkxf7f2Rg5XS/0gN2NajM6gu0uDXnO
OXh+8HtuVhmtheG3P6rgfH5K5wg8NGrsMsYuYpQnGJcE1XCqzif7Q0hVbA5e/4PX
w1Ah0pLBAm8B+UarTLfuOkKZsco5X34WVX/CNsF9iteQ7enAYA/AQe/bdJn+Y4OP
ZsRxyUX+ueemfZ/zXgQTp05AIJKDm+RVsYi7w8dARzRSYlXiTGNrdreLwrn9y/Nx
Fm6FnaNyuL4WKAP+G8YBlCOGk4FO4UaRmUQchQ2YKED/Pq8GjvdcRvfiPTa4CHBP
C8XE2DtTSizyPel5dsR5+qkrJxgz7hj5b4NKHEr+otCqZlTIyKbDzEvsRkID99kW
yxlJeqE+FYmSfr8MIoovv6efxYF0xRsACdB3XMEL5Yj8cpX736782gpwRWA41fVk
ag2ZFXUV6UeFqNFRkQv63KGUb1haw4E1uPe4PpZIL2X1qg+n+CR/AOyqd0LzhnV8
izzToNnnC++vRteIiETrV+xXjA4PbZfLsUIWbjdN3LwO+Dk/ITOtuYRgV0rmd48H
JIem96DWVABLknXpUOcXczy0aN2oS57tqg4hLMaWhPhL8sI1lylMCJkiqYv0eDVV
agkJvo+RiEPbFtu80UMfvgQY/vqgbg9S+Es24Xnef7ypmX7bomMqQZWPTUEHgJhB
xxW+MJJQWYqBz+0rTeRdVYIuxW0sxK0gJVp4CkW3NLlrCXYDou0rikrzc1dgpyxj
1mWOBzeRdZCaaxLCnYBKhDJRLgwTRfpuW5Jz/cHP7SILSHU2NCZpapSKA9YicOG2
1RKCMJFBSH8ayIWgxcSpb26bvpZsW04gxs+hjP6m+QkzpVHTNRTftS7u3swD2wfr
RjPzqYk2ZEiriV9PJ0RTPxt2G6EmIdtjfvsDctBhgiLsEXnMHFvr3FnwtfiGB6ks
lqZa4lRuKLWtz3mABpTeakM9T51oxTx44urrYHF7YIun5uw3Ux4X5FUtLE62ee3D
dDGMhZ3eOqbUvyg2kRa3ig/ACeJAL8iQAOLTvnAmKGsmCzfw7fFWhfRq5VzXiABA
3AcMhOwcajtqKJOy3TWxt7RUts1aCeGkhCNfLT15wqnxNA05NAxpd2ws6QG33CYW
ODvFAQhT5ISZFlSHehqKPaDsXLJkSYp2zMcQ6toNo3LgJwsykjiGg96y2dC0UpEo
kCdNgM5mMBDFUseb2ngFFeDccU+GgCDxuGjl5b3DGS4uvpGeLKcXGOtFsJsFH+PW
7xvoc0NGrBh1tE6+GbTHDCwnCZq3oaN6CurM1otXrOwKeMcIHB8GYGvoPNu7l3qP
e4kS+rNdtLhe/VxV1lTMnAccWNZk2+SDF1n2hbrDzD1GY3M5TXRkcF4KYW+vNANY
SdCfUERUOLCV59pgddnoPwYOPEJvVGpRCimLO1WZlxtsu088SRaounK9Av94cbcj
MA9OuhKpHmV5RL8/l18+yotHSGb1rwQlCa2WzC3S9JbI6MPnx9zRi8pk3tqA2hfg
aYoypIxVAjUvQoDfrhM3cQzT5uG6RMwYC4RQmSVyqbvdXcptIollAJcBAe+b5Z2Q
6GLcgGk8WNMcKT6AiO8QNHlB0ijkAHjtlT6HYE0Ttq2oYYyHLNjwm7+DRef4LTTr
GBn14pzvfffdKNyKb/2A8zh6f7mfivHvM3NwirFDGtb8f341DceDmfMSyk53LG27
w42RJ0v7q/UZF32PpBTb/8D0ce1lT8JZsKjP1SxizFgLO0FZ1PyQr7RF++OprP3/
BLLDkCNnaE4rNlj1JLn0wHB3eFboMTD9M1TuqhqZdDHbaFRV3vYhTaotxXsCDvrz
AwDTht4x+s26tGbNY/e1IcF+alPs+17TEz4mcbkCpEYFyIfGbH2QIYBXJCKzXnN3
HcGegsmHTa3I6Qw7GEj7smPcTkSyeehnAbhin5LmnDr/J9rqwkws/KUjPjZFwODQ
qb4U132kuxdfXpWr2Dh1EpRjKkrfxxPRxPwRpEa6y6R+YbaKOxvmc0JHdCvaaO7s
FVMbIlOWqf2n0KsoUFdlu3/UjCSmrKoVJAeMKZi2pdtlP9tIHP3j4SUASABVhQ7J
1wGU6HC8VbgBpQSauD8KgLfOTw1rhcF8WJ+GnUuGgOXS/qtJEaMr04bBP/XInV4S
zBXEow/vfa+behpKBsZKNl8qcSbdvcePjH3xPVqQtwm4iKYu8pehpmtN1diWTgOG
/2RnfRoqQJdMI4j5sL/thIaGH3aS3CIXXRewW6xTcf2E9VUVGe/C4BwRJK0eKJwg
yHIvF8UyX85OndAtszz7Vg00ijo6lH+2LEvk4ROw/srw2zD/Pj5v3j5D+em+jkED
0QK1/km1WVJCMHnDV6As6Z9r+YXhHBbIq0ItBGRU3g9eWk+RRM7oQ/Tv7nUJ0VDZ
rUW8WIUApaWUyfjJz76s1YAjEvxgHeqvTXiPI/f5ZRNOHlG4vYWGjgLWTv1hOsFj
e/57knvIFmWt9Uccc/gUgCAUbVZ45rqPimAnQ3iJ/XLrUpH1oxOcCyFresni/0Ux
YcVTBSI/Jkt7oDtOJ5WDV89Mu5fdlmXWLSDdvvk0d/6JSWg9etCAmusWH5pudL5f
O42M9ICyRGMlOPL7CCTrgt8Xc0vNO9gBtd3M+pJ+OguWB03UYekK2u/I9DmTV3Os
XRyzuw75o+JFj7CJvPfn8HwTGng217NCaCGBF2X9VUKDiCRBl5CwL5fp8gyVWNQb
D4YH+FtrQhSGpN2+qU3XSB6DKbtgWbIMMVryn9RPoGTrFkGS9Nfcg2u+FzcPYplo
y6Azlc0JGScK8Z/RuhITr45bwZwsZ70SpPcHRMNRz5+qg0JmbE3oDMtqEgr5v7La
eL6YEWIqMl+9RmsY2IO6FCTtkW9dexu0GfPfFfXm3Ygss5XZlMrpEEf2Kb9z9MTc
letsPXdWQ9iJnyuItpVoCnUcVS9jTkOwN3DIDRwkCRLhNilRGQn8TZ9/ul+LqG8k
SaEwHdWo9HawLhm3ZD7FJnJj2/0jW3KLRwVsKxvnWPqdZ5imPItx++7nRPYeMoHW
3UM9+TzXCSIHUlo2d+2T3DY98xzlGwPRDf/Zf7m4bU3PILB8J+K5Y3p9MPr8fq20
nZhPS5qkKU+aH6WNeK+a825fiGSbo5YvAj+N3CySFtxTsYr48D/XybTEd7jK6h21
ctKmmxcpT7QVN3/dKgWMiw02iQZ7uSE+yZI23uQn7L5zJkstV1HsCG4XjydRt0Ta
ryldz5SjFc7MIjDM8lmNwACzo50T/jVmXOcD0m2/vFhLQZKRO9RUiT2AD5/1AsQk
3NlFwqoOS2Ci+nX/eNmO2J2vTg66B8AYaoEjprxEjnBPEj+4vXJXglaLKb1tX+nh
+dMdV17xhNeNA+aCfr6Jjy5F0ajawzkJB3FFTFLkhJC9N8atdEwJgidzusrLQfpT
JU2atePJDZhK0gY0PVJJslhMx7UU5m9U3V7KmGO/g8umhGqPuEdz0sZEjLq9OGMo
nmhCbjIYbpO88vxICZJZ7qmze+XSfWlGfg3V8TQ29DvX6PaM7OyRBoUqf9Lf9Gab
Z3xN7Lxag0c/pDsdSImdHVOXp2rWrSRTYa5ZK0/UzI0nviF/IFdv7PT3AHeRwvuQ
UpaxI3XDkypBpb7keBdyL0HqGhf656ag4GGNvdKd8VtmxEyCEsVMIT6sxz7OSzrR
rZdFzcvvdY5Akhklf9ZW/Se4MBtVEdDqVD1m2QwUUL2NDdmtfpQHlHWpGiOxDYf6
2pP6EOCZjU55jOhPMWFPfIgxuN372xXNPzOv3T0P8qQbOq29aYg1WJhIHJ+OXR8G
VXaTj3UJ7d9yqkSLf+VkClOgF12RDwKkbn7mJhYS9rtir7HB+FHt6h0VlRVFU8IW
Ct3frYXCycDUkISnIv40Kvxt8R8ZnEkenxx301sr1lzvd3Ruw4APxX0ZC8p2vt73
97cp4rq4WMUnDCHkDCsdmQQaGziU1LwVmSxQlEZwwLqhw2icCph7HyYt49OliAGr
37XHgmU8BDxpKlPCxfdwX8+oy8Q+AnK9Ds0ECPiycOiybjnZjw7Q3wLtMPcqEFLh
dYVyLzopgrEyRiU/W+APGMrk7q39cKZawSSdKBwIl0IUkIl0GHW0Kem0E/9CFrqG
gGgG/ZmGAtKFXn5HYbyDvFsjuY5s2JkG+yIotRCKJN8ITSVQLsZWNxjEkSEdDiyA
IEGQynMYlFUXUB012omZ0y83zu23Ju/nrcFk3FkXm8jEpLS/rscJdHHsuUq6LG2o
wIwoq5oBnIL2LfD8cKof599OIYr8wZlfKdUdD6xoD0Y6gHTOe4yawmBXPRyj3YSa
x+JH3QQu5APpZFmDkuSpX0zpZp+2Yf3m2vGR2KOzdfdSb0VHW8UsfpNRpY3DGX+V
KcjyuvG8uD4bsswouXYZUDW7RWrypuT7GkIUSUHJbjGXdTtuulmzqTGMyitZpAzo
+zElic2ZSrQyehIr6t5QtsphcbFP0xK84S/bmMen7wdhQ5sHugRb/JpUm/7tJEi6
PJA5jA+cji5klqNFe/nq/cRFC5kKwNwjDQvAALNn9tMDA8R6Efb5sWTsVV+o9Ig8
c1XXoPsTr6S9ZqywAiKouN9i39YcIft7z74HK9q92BQFGZ/qgoq2JJXiupIOn7Jr
TP3qCxxh/76JEn5u0WisRA==
`protect END_PROTECTED
