`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5nQ2p1cWysicnBd3SMy2lNZHbaotvB2ApCfgr6xwiQtfP8qiA6W8Tbidd3Mx1WmN
aH4kqljiCn1xYRMjG1a6zpCcIlFBr5thifUHWZAOzZLJqpvpNMh2+MVsvQ9YudUK
o9mrh/S8HmNzfzkiPgRzlZywZzjp/r+4EdBT+u8BVsGbvyKKeFnawqdR121F4uYC
8967rc63dE2TSmTkYGcHzDhvBX2At9iw3kS358sXGsLmc4dHlEB6FrRiaYhCtdWo
eTv0FneJD9Ny65Ly1K9VE0ZGQHkRiuDZ5iWAoH0XZSKNS9iN3c9f60SURyooKqCu
c522osAMLkqhJEIiuGMnGlfTedR9k01JRB8lJKWM86FdGXQflaaKVrDHhFkrTlc/
soTqljjdJ+qugfrTe6lbGtRW2iFa8PGhTUJFAFrvH49xAJr/ornrw5lEPPkITJBu
MeIgdUkb96xg+kxXS4nueV+uMR7HnzTQYjojDXMrSsEj/V8I31rQZG6Ci8NM0Uib
AbBiieMDW9wM7b1608h6w8wwkbrslVpaNO0vkaG5w82pfcK+GJBMKSJcIvMHyiMj
nr9ESyNRfESHdG/H8rRSfNkEWm0muPRoWzE5zDpFGa2Yu87MHLfFIaeh+dRUnBZV
v43mbtj8kJivo9VavE9ywXrYxSENKoyjEJRMMfk/hUYioTrIqlJmaHFo2cksQ0Pd
`protect END_PROTECTED
