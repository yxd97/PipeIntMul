`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQ44SurCL51kgRhV2sLUt46WXkPbjz0dUuAj03eePxvZ/0ji70TGLukhDV4w0C7w
u+3xfU7pz8uU8lLMVQQM0+n9FD6dRTPQfrRAA6sONyvaW4JcpNU/P4NnYe3hFNIE
IYnVJpqAfVgUwhBTWmtPN0hxKUsnHcq6Z4qHVvT/NsvadVe5GzaK9Z8xeYeDcOqv
PT5kwllrl+ABX8iRFLBnsL56CXGU0DAUvOGrnaO99ACwhX+3CuZCSdN/Zdfom8vE
wUHPuVcUOjYJLvLD9qG20ogPcWzos0KFIoGruPlrRmXehRfCaIhwB/Mr63jBtknN
AIqBJjhpmD1ErlrEQ0pcHmKvQ+I9QtXUGFgPe4Fu7zV6DHYpuo8JXB+beeqCiG0S
oTzgRIaU6w0LgizUiVqsZUIRpfk3U3yx8ZAkrZcL2ZA=
`protect END_PROTECTED
