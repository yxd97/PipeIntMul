`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubdNrJZLSyyIXIUV4c5ktTXDJ4jLlwvOhZGqF5qcauSNix7bgAlHw2FH77ihscFg
y0yIWundbY4qOIXUUA/oe49BFM+pjcCqcqzJkrySTqlVwhp70lkodG76WI7rUDe7
AfAeznZ3dV2CVKei3NeHibvzSs9+sarN6JfZpsUo1dnCcd3JX7ZZtLjYP6PxjTOR
EAcvmv9P5YD99AM0cfDDN7fexy6+FtHcgxVQ3I2En2ky1E/xOxh2bs6TyhqetUSW
PGjZjXAmL3sjai+x8LmCGqwJ/pzkoCuoKWuhPeNc0L4IZdmJU+eQytMpeg8cGZkT
zdaFBJDBjRPWlLtjpQ5i9spx9Qa2Mczfef531mf+h/+kdTD12jQFIaAyOFPbLyKC
1RKfDkX0WoVve0AuQMjaxA==
`protect END_PROTECTED
