`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnswKlsHdUJXTjkCk4pNec/F9vwfNKHcZV27B1KMq+iqrE5A1U+0CcGtL8FZMuU7
6LHEPT9YNi8HaXkVXvsT4gA7lVRateR8tU6KxUQCxCnLzZw+tN6z6QIXxCNu6Ntj
tn5jsVF+IyglOtLGqwfc0D1OyC2ZgYzXr18dpIytv3YAS2zxvq2DLjdZSvL//unT
wDkXfznnGO+TNCUpsZHRMX3psH56BY453sdmHm8tiiDs2VxsXiTBR9pacmtNi5Ov
gMUWBgWe3B6t/9AsRMJhdadgUEbHX0QDdNYcePsUrVPpvmVA0CHOzzRNZ93FAYhf
DvvjJyadt0481qkiJoL8rSDQ4yEJDnhu2PrHuspL4FMXTGLo23SKyzG3Vs9r6MGo
ggxotSBtztU3Thue36+IVLlZ2a50xPF1iZlRGI5y1rcDr6FwFov5T5BFbkEuirsT
ivRn6o8cOmZ5/U4u8Gmk7F6SA00U8AqHtIK6rCGf0jr+o8+8tdAqJqzFdQtpgxdy
gxcp5Q1WyGUjNW1wdifI/gwu3wNisBv4uJnUcWvlVip3osHxdFOUkXCpu3Eyuf8k
0d+N7LVR75slouPO4MY64Kj/+MZ+h8DUboA8+eE5dzJUxBlxrQoWRiewZn8AC4Th
eLU97em8V30aAXWpztbT5EYAUe/XSR7/KNJpa/h752IslQDpvAzGV3y6mi+/7iVu
Q6A3S9wFoANEj8Do/6TTZ3r6HknTKgzHso7cXhDMsqIRmcKERGDw6RbS+RTcpaQH
4j9leSOvE9M/yNCXgulgOUhg+x71YHpiUYecT28aFuP2JSofSlg4fFfOr/m3dfJz
3Tr2tZds2ary2MFxM588ykuBVTAEs/fHyKulu4J4GKIW1DC9ass+qZ2PZyWBuhIf
5wjpiguE6VFf/Z/YLc5Ik1aFVmbYIzVR+FTNBG2fKs6TumxOffX3Eyef9JqEB9E2
hSApNELuGGBLGkby66dlpqqyg2wv+I6uhu9o+wNVg36IDFA7wLSLyrDnl7K54sPi
5PoOcYGIpNWFU2j3mzMgUc57RGjwTXmwR9Kbje9a57CEMNeXHxpg7M3yViGkiZ24
3/2i6toCEdo2Kf69KRTlQyiB2afLxaiGOkMSmbEpr1Cj1BJrIbOxkm1uzrW1A9Ef
BTi01oEuq9VSWWw92aASp52hAOQfqDgo1k/IvMQjd8Y6nK8LPIGdLfvbD4VVEymu
jNBDvir890XqPbuK+6GWp9jU4yGGBIL3HDG+tyW6Cq4QzHJwvlYMGraLTNfVkQEJ
4+y8NVDT6Dsbce8Vl38RuXqpMaVu09PA90a5e5/MGpp0teLFw8y46hbsTM+c4dLh
44a7Z0eeOGVtbyNH4v905jsg4Ck8zC1YSihNaB4BFGeJWoe/uLPOJVrC7hz/RKR9
BGN8saM87GXYJXE8lMFHZkVs6Jp1uZtTAPdJjCbjAX7XxjEQpKpsV333cSiuPS51
h9RuoLcFUFDe38Cq/xDnHww0OnVkWWTHQpljaP9dGTjnirKefwxRRlG3XfsSiroT
rz46lgf1pzlZLv1Q2F3IYt2/jWLVjVLxRLNo9toujtN4os2jUc9yPibtMjOLB9fs
8/1Qb2CJu7PadzZvjAp55OOECTofn5tPc3Mg59ueoSX9XMKIUnqkVOa72fHdEiAE
FXa0uN2i5ELi47UVwePr9SN7Hoka26fVrtMq80WAsXHtd0zEp16HQmAJJ5LGry9A
DqvMCnewWW+ZAzs5/7ZcTtATMqpXdGaqpCtyTasLzfLkgs2ga0qoMylc2ni0Ealt
OdoBPNtFaKhW5seP8+rzUYOntmvFb3f0+8olyM3imyQfugfpiyUhkCX2xYy/Ju4O
CBAdPiYk09gwvIylyhpw/JmrG9U+kNZQsm+IzdOjAwUf8jw2Qh6bfsBZ4U7Vh2LI
WiLhFqDsGQQWlKna7ovuYUMYBKtIvG3T3WvImSdbYDTllaA2ZZDIu/dTotAfecVX
Qd0f3BJDrriieEskhlqMxOb0SL8/RcXnL+2m0Gj9FKhFdLHzL4Ztsej+plBNlKk0
cX0U3jcw9bY2/fl6esftqZLZ/A/Sgw3u/czhzNWIuXI0R31aAljdEx0WUEcrbWJK
sIarWYUc26MOopuVXCjEh6v1xGlj+fAZiD19EhM4WjZzJg1D1FUx2WSfYomWrkYx
nWfwIumIDwG4iEBw697/yqGNgYqnjuEKTRGSdZ+HavD9kGoZac00IurUWGxz+GO4
rX0AD7RWzU4bT7Fj10hcAVlm7piKhJmdTM3o4mufa9Y2SCDZh5YVNZNHBGJKPryF
LMrsbyfpvNtvpTHEYSpCKPH9h87R+FWWzogxnK4TdDj8dzTsaSf/rRzAud0bqheh
dJbRxLIJuQSvLjnAC48/W/fIbP6u/VuAsLFu+gk6AuJPbhZOXk1aWxFMtXwxCPk2
JvEboxba4xyDqCR2bhxbwlkynFAddAPH9aL7BcfLUict+0KzIPX7uC2dJU6GowIn
j7nawveg1O3bwoI/Ks7ezB240Xq7Tko5vPwHy9lUI9jwfD9L7d3Uw4fMiAH0mOho
TWHQJoJ7V71ggC/JLX1IDNbIkWQI2m2K0nInd5Q9gOYenc8sDgjMIcoTUEdDN/EB
`protect END_PROTECTED
