`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mb2+nxqRQyvevBEEYwp5U0CR3ylbS1M46G2mrQZkD110a144FinYav/m3K0GisRh
H7nJitavZQiNR9yE+XiJVuDingEVfzphGusUMPvYCmYimkHhawc013Xrqtsuwoxh
SSw+NzJYjcJVIEEDJ3DA3PyB5zI4VD9pz2hYzHDj9rZhNA6d1dW3jb61ifI9LaPF
dfrOVDSn4xosdDxMBlaD54vjeGQG+a8v6XKH4ihEUP3bgKEJ5xo7/u55A0V9mfwu
YaZaDA/joZww0JhK6isC3+tgsmGyECvU0DuwHvkQE3NjFe5nGUDatMOz9iwGRtDX
CnN7jSZLTS2QzxBDVZ2prG8IM8BtXUBkPoJpECaWugfj1CjPk+3QamQrVxO45IE9
t7EL/yLo56OMbslwQ6EyMSgWxX0bIQN41h+3S/J5hP6hDtIalzT83+WJJ+ib/jIP
h+N1AUXzf3vnGUwEiwe6iIBjfiWsmE3zwe16UEtgfnUTKyJQXN3jggygCOqQxVtB
VJJ9v12rCLhzeHk6VuzOmEFMf9qPwUMGnUww+J+QN+hv0EGwuGM1MTgJpzEuhBG3
9JbDQCZmnfpVwhuO9FerRlmbXO74maWxVf9KwgiekBpXWRHKokiN2Wv17ia9Pc5W
mqC23dP1nBzmhV8i31au9GA/gzrq7FEEpLRSLmV1bteUPIBxiqvnI8VEHzgTo4Vu
6sx7CFUx/wGP0x1J8mcMaIzY0zINqM2ZepBdOLyUWRmXygAl2sC4sKQQvCPEQR/0
CXSF01OGVUCbC44s2Tnukm7PEnUZ8DjSdxNvfns8nsIzo2Y5m8cxbwV5zGrg/TLz
CxQ0mxio0gqKlK6gZg4Xo1sx/a5n2+rw4CvfHiDHe1ZRvC03tbKUiJimKfupk7Ho
1+F3WtQ+Cv7T8aiiLjK3pURLQb31JVo47x3unzdI7X/SWYfC53WlX1CymuC2EwL9
wpVIffjaGC/VRVSAkF7s8A37hOAT6orD01Lcn5Tlj5j1kGQ3cmEJ2oYtae3f8AdZ
`protect END_PROTECTED
