`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z59O6gaQAl0FbS+Rdv+S7+Qr4ujCF3UaCHGYvzQaDHHByRu/1N4XCqiPlfTH6arD
Xajv/Q27T1KBJnN9jRp5BYe9fHWTisWBaLuvYuxcZdq3rD/J2GMRNPrH0nbvCYqn
oRxvEeT+pKmOCQes/KiriCJgWZYE1hEn0x9ldoWLeMmE2Y253CxeCkipasRm0zAV
8dbqDJeq7JLB3MDyYYSeM9QRBByHFvj3jNOvzPRS2bl+0iFk8i6wQ2nRrxDBwyyY
eB8cERknyG75CHjQZShCjA==
`protect END_PROTECTED
