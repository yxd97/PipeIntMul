`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuVKMD6L7NE2lLpLptuQw1lNB0LSZGmHfFplKSCnFQh0Z+cGj69IDDAI3HDg6K6k
OJWH+BaK6+6lmt1HTYVgp0AzGkNzEs/F64mZ1n71X0OdrX39Fdhu62kgOSnH0YVu
CXAI9qzRkA8s15RDZlDheQzUYzZge7LX6ZMX0sxW8bAYRS6I8HJhdfR0tQj70yV5
qaLWcohBkskgeVN1czABoEQr6o9TxXa/LFaZRMQ9O6dfgrbMwMIle9zF1YJMmtgi
S3NP0Qsd4d7rGEsLjwgIaC2nArhjl6KK6qrHz9DXkUIXjBwJR5zVcs6cUqnW9IgB
YX5Fp/1109xCw6LAc0TXyg==
`protect END_PROTECTED
