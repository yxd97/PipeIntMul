`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9V7SkhCu36oS0MYB6SUcWvd7Bu4cW64SIs6tSq2fJ2+487CQ1QSOoqrz3OV1XYp
ClWHAO1zI0J1BxX0wc1DJxALxlidVI6xAOaRrClY2o+uzLbAqpxOrrEqzI/xM31t
i3EYtzjN11TgdZ4v4ZpRdWQmurCOnQYGn5+1vPtjDdyfcZsBVvnttnwe5pC9eB3i
7COiOAVFyabF9ymoAj87lrky7gKUKw5OpIg7nY2bA+mdRchmunP85ET7BxNqCufs
wCDYzk7tas/pOKxhnTaCd6WFa9PD5bIZUEgOcu9YFm2O4HXhHW/a4UJNR0Bf9g5V
e/krZ2kHpjkXKKUkAu17P/N+voV3X2TO9mGenRsUczqPvo4vHovuJys4DMdS4zz+
`protect END_PROTECTED
