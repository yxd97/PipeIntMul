`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lNx87sZ1gjHBHP+8YOhKhXhAeLl+0HM/sYiVcpmNXcfOIYLgAKdoQjc+425w4iyu
V1jr992aEsaKeRc163wbe9Kolwu0AUjds1XsIlewYU8PqAbJ4zuUftAE0Kfb3357
Hf1qQvekhTsThMBou9BKeADzY174gr/mq5lkgy5aNNs/uEFvww1Uy+F1YD58Vf/b
XaBJ+lEH7ZYvjYsVW+NhwwoKKz+ZhFho/+/WWPZJMzmNbwXOrUmgRxWSASYB5RfF
iabAPancKL8YXgFHVO+3nuE+p35rXpuIZWF51p2AmV/MxQtyMURUYG/iZvOhcWMY
aoR33Q4pJxs7kJ6sgw7X1cNU+DqVlpSfBqSfile5ivmy9v2LJDguN/q1xG5pbI7J
k/YwuZFeRrzCoPcbX/inS1ct36112U9uEL08/aFjR0/2/QkqfNtWUvhgk+lhc6LH
WSC+QhW5OUHh7Gnvsrk042G57qYWadFGOqx71LptUDq9anJ57P9QHdIbCa/wLNBO
8O1W/43gs40Rp+3pv9GThll+RpP38f9Icc5MOoFJHC0q7FS/660+4zpBijhwEI7y
ED3MA+dbCDcVJe1WIrT0pPJUXNGujc/eMJDTNiS45Ibsz6TVLt3fx2oB06HFzfF9
0l86sktisF/E3uz9JUOCv6pJwX4PppAAlaBEejOHQaXJnhGAiQ1lc8+RwJS9jd98
nQ4AzCcDmX1z70BfAqvpIJV5Cfx649u2g+qEazhWgafr+Weea7du9PA0hw8yf3I8
qMg37uXLmKEDeRMu7iPyLl8aNieu1n459joBdoMWmqU1cgqZJiTQcIZbLFxxs5hl
TbamvyJanYGWA58AMMc8q50gEaZ6TExTsw7rfPXkeIGRGXUPMN/zkCemc+aLuSvl
`protect END_PROTECTED
