`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vWLApsdwWVa+xt0uokI7aFm/NTVQXJUd1iJMudFOOhp5VWBetM/cTBbDl8qR7gVr
Xc++XtL/ieXQeizt+8em0+Ef6gNRVDD96FzTIJsKPJv34gyqvq/WA4zEiIzl1AZw
VWD8bB0KDTa6QPwToCQPm12j8DRMvf6LWQYHSZJMyU6mtXM66+kK3m9hn8eUP/id
QszYLKfD/wAnYLIjTLq9qnWsHMGDdhjsxxaawtIu7EkA4dM9AMaxxzfo8O8rIQJz
vH+QzL4oOstAhopwkM7S736eR00vsIUNQjFk8nLGbHoZvWW2A5Hhqm+u90mwc7IZ
zGUvroJcGraNLaprnfhFeOr/tn7oH5iUvORjAQnIRcmB2dJ3nYhABkVvmAc77n8f
Fkb6Olpoicy06m3eEi2CHUKVsqomJ9LsGIk25MeIHXqVt//hWF1w6ilj8/8/9rNI
aCK3ZpDRyow8Cnmyt8Q/GG/ZeVyh0cF/RhlrgNIfxsU6BgDoEHTWdBgHCXHz9GFe
aBqR/BIn3y5fDgROAgFq0kKGuZx/L07wENoXrCHn4SHEN64dbQVVlkYU0ODduOfd
5grvI91GlgnXdhKvZYnS0eaT1K71QbSC8ZvR6GUT7aJR6o2PXlytWj+dUjPN5KFN
AIEEN2vnCVN2ka+fC7AEViPZihnXxodk+8Q2ZGxFaZfcXBwpoZkXEatp6SO8Tm/j
oHidQQRBLAURbC5nDIw0ZvjT8z8kBPhGre/1u95UA2OAIMhiLdvh/iG8brUI6Zrg
O7gcm6x2RCgPT4f3IwzPOw==
`protect END_PROTECTED
