`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oyLnAg7k3NBkv9oKyoH0PCnMzUjBtFrZ24XuAe6RsDt2uQifSuGalllTS+FEaHIp
AFt4CuOAFZN3Gc7Qprii3staZZsoGvTzvxfwGRFousG/gxo+Eq7+WdkbYG99Kzaq
YTQhP8kO4z38GnBpe7/ZR7uv8Z7+aE5auWeeqmMZWZpNwFIu6pTSTQUfEL2TYzHF
88H2x/Deak5g9jQWsMDgpM5AsOFKBOIsm1y/0x+tUrHEQptjOueQ8nb9q+ZmjInR
vxMr7u9twQJLZv38CqEVvJPmN9Gpuz0cGLa5vl7iM+8GDSuM9IVfliFcTKY65eBO
uZZJAVFcAE3eqikpsLWMk3UgEcnspU1MjbBA/VcDXyXZlDJOe0xCZTqw9b3f9nnX
BUL6mfTZ5t3WzHrAVoItZOkkkLN0VJWq8wcjhadPYyDqdTJtqJ+ouY3IoIsvwTxb
OfAgtjOvXyk/4UDD8Z6f+A9xL7TCnh0x2GpAk24RcdA=
`protect END_PROTECTED
