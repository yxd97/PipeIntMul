`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VI+G47DObct9fPfTwynHj98Lj4FY1RXLxSQOV9Ht7ufm0DVYrsOKJP+a1ga1HogG
1RB12c0eeucroTlvb2jSwdamHcU4UmOLy34fz6Cw7QSDiPBMVOh+zve67Qw+KQY5
f7w9GxXefZGBiq5DG5vgCH0K64wCZD4RBmT5281MDyoRnr13+2Lt5nwc8kK0P3HJ
AkSW2ohfycV+By606tbe6oZ5GIMqQYqgONVUgJ8sH1YrOSB8kkHcUz8rDqTWIWjx
lUkBzI81+IkJlNh53obghK2rn6gaYylqilm/8IxjFGKJ92bh09cqh9r5aRNs7338
aT3Swr6F8FsziaGw+XBrNt7I4Yu9VtEBoCH3md/5Gqt6tMKMRkyrusRHEdY3qO14
7qjsLv78x3tRwWGhh88+ycYD/G9n1a9Bu2W/v81I7QSNUzNdhSLmPiURt58y0IGy
kwJFUKWYdyBz26HMfLRHpEa72/cPh/fjlueNNYV6y3pPKU/wgLOCVuarwPygNw5F
UaXFqSC3LcX+PvyYUqHPlbvK3csI5fWHRjlE5TnHOkaIucsxq/52Jk0cXKsxwpsc
/YEgIPXiCrLgRhocQ8Q/dK8rboijxjApGv8ALjK8y29/OKCeo/CKs9xuh21tOXCZ
oGhvBy8c0uBqWKcTiCzoOOqsdHUet9XTp4vJHCdu/dmglNJiWi/lMbJWUnQUIxjt
EQUPlB2w3J1RNt2245ruPUIPr5l6qhQkl3Ra52Ik2ep3k860rfim5wN9aUhg82kD
RyL6YEF20vov+51kP9sGzg1GCrcRLxMY01nZnJ0uijcIKrKMgVehyAQZsEDIX20n
1D8VOSdUKnqxQ6Lnz7JEG1wENr93XoqSM7xHWL7qHCE4W2u50fHutXzurDzCrzYW
7/Hc6yIPzeQbHeamYsVlIgfG8WuuD6XZTNDNgqNy3d6kQPvoZLQl7OuY4WBrfnyB
gGQUwaV8gHj0aZV/yLAfquQoCpnW2++TifEK7iqlVlHqaQBOzhNzxBrhdf4oCOOz
zZ+H2tZ758aUNQwlq42WF1WaWJvqdN0EYze4+sf3OTmzyrkeK3w8L34rVwqtaV8v
WcYY42WN3WCKqk/33TCPhKQ1Dtkf3123vS3BGwFW8kjem4vrde344VsRloXJA7SW
eIlHFskjvnq+Ma9ZWXgD9ify0zkz3DPKvLkcmRz0DQKmwKEgE2wsW3hrdaFVpNBp
12NCxDPYmGtAVUoqhFyb9lZofuCkf1bwNVZS8HrRv/QYfwi6YEixU/gHdrPq4o+B
`protect END_PROTECTED
