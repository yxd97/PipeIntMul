`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAMoWmw8J3YR/DpMVIiuQ9S2ZNWLEJxfv04rOKVrOZ4AyQ0gTGZG9P3o69OJxj0o
/tI/9ATdLnIT31nak0xUjjSxGirbd0ix8zTBewMn0z+VYBjoBjdVBvm9PerAftbs
uRU6dbKVENKDHBNtNaU74syfuR2BN/WJhzRKRMXPWBrqhpiVN87A4Zt21BzRipjO
yuxvrN7Pa+W/3gA1I19rJh/xnubpZpnp2Jm1THtEY2PQWOzH0vS+ESDjmtAlF19T
C6YLcq4CQV35X+xhiKnpu/zJlMH45aBwpB2/8fUK/WgHYRLbCRX9Ma/NL9e3hP9Y
Xb/BZYtZRBcr4DOBHwf7yQIPmeJgDfB/qm/zzQlUawbSDNUAFts+W8nT128Oaf7A
j3PsZmZyYWS1ot1L5Y5EA8e84W+hYvUF61bIDL2GSbFFp3/XVrqztmDC8QON8jEI
xTRaiIQFQPW1gpmqHsPtVw==
`protect END_PROTECTED
