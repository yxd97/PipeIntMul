`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mBBMR6maBfb+7lkpVREeaaf5Si48UbyQs+cCJxq7RbXY9HPLpd3mwedp6g2jszQz
Wi9GRSO4Y6Y/JLEIUcOvWnWBmoBz7KvOkUe8WCLKz/DFV7gPy/25LxpempplKj5w
hXoJq27j5MU3AI1OL4ch5JBlr+/MBy6FmNF9PKqaH8hX217GAfsXO/AcxNDTht3/
aQzLJOnfB5oCOJGPkDr5szScqOPO5drx16JW3fhD8K8xHkyRROqVDSaZXf7CmSGg
BcH3W3piD5Rwq16UJ6VwVnlqltq7j2wwCEPvz6N1AGx4AYm9uXXKASI/1+NiPqzn
HZueRgZ7gXjVbEMoDvPq/bx2dkFfmZF2QHrY2njSfNbVewSaImtQKrBAIzuWaeNL
9CO1yr4KH6wAwuzuW3n4sOBcCM51Ol0yY7UaT9lIFDAVwYphUNtUaa6DYbdCuGL9
061MdPFAUTxHWA+wYvn3ws0cM0M0d30rsKe/PsHR/hpgQu9DVgV0zG3vd9YNHR2A
ZyM4wFBIQG4ixucHsnaQvk/lLisXNa/s3V+F3yFWlt6zqGEEtYSYPygewnnqLsqf
Xo6Q1tM05lbvDWHxgSVilUOE/lEYR/lY2OwXYMj/1XIuKWdytqMUAXuD+qJlAGfb
7Whg3cndmZvoRY+VsxLXjzuB8f/1JIfz6yQLUTtu2UIaYP8kssAEac4tuOXcn1TY
lXbulR2VaSwODIG/mBeoLw==
`protect END_PROTECTED
