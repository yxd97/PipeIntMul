`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gA0HJEWJmSpnm1k/+I+0DgZo2rGa1fYwdWZz6MpRil2r/0W8OUJy69DxM4/890a5
i3j/FdvtgW+5zEYkTUxTZ8VoYhqoccRcUrwPikvvpXFf1oIGjdqetvS/AoUejamF
Gn7DG7gfaXHwhjxyyEP5wdGgr7mnJnqHPmLxFgx9EGhCF94XgCM8L2tHerK/aj16
lVBjEGZ4g5IcLFHytNCwUOcBMmYSfhL98v8e/ANKXbD1yXNMhuCsAOnPcH0vGVIO
1dCrWh4okcmxbjcmwNRXLUwlE8hjnTl9wOiZXHxT2wuAaaqzuFk6HeUxr+ROd8rY
gSaBmUN7idmg1iI2SJvSLsW/NgC7x/khsLjmMXoVVvuyDrOrP7mVHH4LgTDNlbh2
hbGhZ9j8SiHhifbDH+vPu+YtHv1v7RvNIXngu94UeaLpQuoZ5sDuXn+raeYMnA2D
WRfNbKEFg/RA7AFqs+K6Ztzf+M3Yy2sHdYGjpa5+lLLSCtpPMnnUYWAt/rOPjyRw
V2bBRWAKwqTkKjSBVt+H//HztvmOb75hEgq2saNsktDtkuXaCqvtYagwbLWkVWsQ
qXoA4mjQwhOjgoj3+suBktmSFvh0bv3xRhP47oyQO6k3YEtKu6TbnGYmxvHl67mp
OJeUdanS9OqKKi9OR9NGNsEMyLqCpow8x1PXvkhcisGp9iCR6amxVt485BYiB/7b
RI6IKQF+f+4In/XVQsEe4GjLl9ZNbOQc679VdCaj0+dpRbEmgwn99krnYjoDrTD1
0FFSxf9mWku5ORGuBFkHXjwIPOr7yrWsMrJM7YNAzfyqE/hzS81HyH5Yl+Wxc81y
TIntoAnCTigcxF4hs6CbVlNYtbzHssalPqwTKkHTqtxkS67aCZeFZSrjega0pPLa
l6UWEVyvcix089uZ8Ir6LA==
`protect END_PROTECTED
