`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I7RCWWIxCSWOTUfABld0CGnzECQHoQR52Rct5+hXSSk6MeTL3uJy9baIweErPt3J
p/WCnuzslXn4p994B2QYSIdAGiikDFWTXrTgWTeedCRzZvoVbzwNeWc81Vbsn0vj
jYK+6SGQMLtmJ/fML2m1VG1ysVLS5s+Cq1SF+JdoYkH3MdUX6IZiweuFCP407nlm
xBOPGQU15tqMccSWCRUp0NlNKQdPjAMA7s0QE6M+QMPZUT0Hb+GYcCXOstI6y0cq
xhRwK93c5zHjjjBtAvk8E0ke5zcw6daGLgrHGgeirT7I4/+87a9vBUkLyxnfNQii
4/IAiexWsisNCtpt5XL546VG7dW6e3CFTSPBKg0bfovcZ3ZR5UXQ/Lvx4jyH/YJi
bPyC//gzq6ec3skUWmDjvw==
`protect END_PROTECTED
