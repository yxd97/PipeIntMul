`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/Y/L293UmXVcK7hq0BAwDY3sFcOPX4Xc/xW7H7MGlmWo2ajPvI5QPDVwrxCqPMw
QfWGK70n5blPyn4R/aV8UK59zJeb98ba5iCOKw98zojwMaGklidvIpZ9NjVwkTqG
LdNZ1ulfP6Jj7aQeXhaEzDl+FtDxZPprfORIT3+TQxusI4x+Q0/J7Uak7SOIllIF
fN7t6i7ejwiQt8Pqh3jOrnwB7e3rHi+05Vtt+28q0vmw+38Bbtj9o/KUeudU5etz
6JGwwNYpImtY2W+Zhs3Z26LuOquznjrDOYP8ahCFRT0jNgT3EEDkYQ2Zllc91zmu
vOS0rXm1Fd2gSjvstWKB1BivP6eg2X8GucKkvk72DY2ybCndXFPds4vBcY/W6k14
wHZ8Ux5zsGzWwALdpTg+UBCYZYs9lXi8F7OveNiP5crkqIgF1JFDYmMs1iyLBNQ8
i1smTnKj8nQAKMTOFnNRYpSsmKyLmB3nImahP0IHk0xJWLLZfoNlssRRxGOEbIrl
`protect END_PROTECTED
