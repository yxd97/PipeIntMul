`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59O/nbRBtmk6aoAoK+Y2Ylu3iL6KOLuTUd5zRdoETKuXp7UEJSTawOyZAV46bWOs
cZBEa+7VdYg3I2Msi0aKtSg7PtXlQ31ne2fvl6ulwDtGMqSNEFNeNmEyA4KTnnEq
bXnZ2QeC6f/dVngOXgvEDrq9XfLwppLVyK+wLYEGjBH+fSqnnIQ/3h0vpOselRIS
4j+aCjn8K5e2MaOPRcQpJKToURL9KRUApzxRbhpGYHqYEqS74kX2BSksfcfF+mGx
hk8TeKVsbt7zKz2wTLH/90vz9AEXySugk2SkU+VfCPaQcoCPxQkAJ9hDZo6/B2uf
KnTghGPIh1/qKTOgC3K5VA==
`protect END_PROTECTED
