`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5fSfoskY683pZxaoDSZcDrKrBnyD7/ApVsqyAfqAQXS2d9QfJAU5y0gmczfzL3Au
yfx0zUFM0iyNV5UrRs0C8c2Ru0bO2bWGxE0RB0sBBRqWq1YLXVQEA8C3J8qwk9LR
PvLn+apvlFjuIboJNmWtumm8tiP7kkAcone+TX3E5iUVUKy5VS1MyabjK3ZaZfZS
Boe+RLcIsUhSl6f/v0hK0Erhruc8YJu5+6kVY02JEXBcK+ob6fc6k8G+d+is6MsM
yaDadQIkGcDI0hwFt0B3XYxojoQ0vctgjdNwgXEJmAsM8JLxox8sjmEwlYjnMYIL
L2evStWsCsUPH1PGUblMdRAyZBFiHWaErDVfEGEhoztD+A4eapL2HEc3faqPPya7
h75m289EBxHKSFaGumFJ8Q==
`protect END_PROTECTED
