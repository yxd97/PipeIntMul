`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yESjdaPDPdiGd4txL72Td0csrOuSQ6aQfhlSGNectfilHq1gI1GxkTry6AF4zz0U
wlK1eoxPZZHbBiLxxE/XfDmVp3eHJ+Tv/DIg+k10n76d2a2ZEvIMn9H98Cedyksc
NfbxEb0LqOXWGLMNI1MMGzFShck0zCDotpZ/T3IgkrgvVHvHOYzxE2nmEKZ0wqto
vZ3BedZRUHmMN5tHfdHHNLFcBYDbsDdQeWB7S7orDAb6Fk6QFJ4AIxzxJ8yoLfik
gtLNLwp6O3OUC8CB3j+0b3oA5kyfC8JxDYE5ZrF8vXkVY/o3UXNDINiWCEnlXTtB
Q+g2u0YbAIK4qadfOGYggbhNufveU1NKSatyIgHaoCQ=
`protect END_PROTECTED
