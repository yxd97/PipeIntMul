`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ladE8olZTsJNy2gq50hURWd/As3vL0fpdy7liBg7/JhgrszeqJW9tv6PCit16eiP
d8ssHTzVeD5+j9KLwtvV3NuBNT81nt25Au7qluR8JSAg5B98Lhd/9+lM9pJEH0wU
5MCRiVpMMSaCqmIYss+rLjDC/Ml342XpdQ48v5L/nA0d8qMRpqCLFEgY614ppqMG
hRDTcidNtZHkRqxy/lhuTmLBzz8fujBORqvYkF03IEKeFmiVq9/X2b3LZesBdnUu
8ANNhcANVl7RG3fz1yKIQpLBE+nn92ztefxLwglKbezKryyhxhNN3SfeoLFWSEjv
ZsAqffvSgfOQArEoaLXv30fLPpoFhBrF3dS03Wdc8TDjpl0o2dB32WNbAPvohMxE
dq/BME44b/zkgQH9W7oTsfeOpvQ/97B7yKm8ptXzf1h1IYDIpb+J6byhblklOwYm
nJGmmXiFQ9oho4LAgE+CKTMFvzFMy+Z0fpI8Ielvmc95ItKDSotWupVmJInowtnv
4nG0GtTnxz7XIV7dcES7S9H8Mc0+P6bgivOBncCeCrKH2Zxjs9pG74+/ov2PNzWo
6A/2G79Qii2oTvsMeh+KrMftL7vZtsUNBb4P+UOB/GbTgba9L8jh8z2rjVXTJzmr
AZcstpCYr1a8nWJiQHALBtx1+SjW0T/V1jViVLB8VXnppLsSd09T6c82UGmpghwb
Fj9lxOIOJWx+hSqgsMReAcd/vJvOo3k2HRerBfamwxNWF/JbK0lZ/9qdNaYL3R7D
CD+Bnl622MskaqYGCBq8ttkFPgDgMfuIPob8lR8rRULKhAMMz2RSe40fGHADEj4O
equW5PG6xgMzOVq4pJccBYa38pyrWEV/tcUjW/6obzeEyzvWNapKpYs/M1ATQUQ7
kGdSz7w0XMrh/qBzsCvMekybdMQNOIhYrEmaJ8KYTnKHh2ywVhjIMZ1eB82zKvEP
nGwRZdd68dPamxC5rM9+5uY+rbo7k7P3JZtcjxOaWTyrGfvxMdXdJY4tOzqQORNN
2cYoUibbfstWBRbcrzFY7jUZPh1N7zRVv9leyXTxs6TEUWZZVGkIeaSQfkfFVUUR
u7vdDPwad9YqKHqYZ4V6FIdwTZbNsGBb8erHbyS8L72vSRTHGUbDwcc+zBPtnVi6
kWq0jFRQFal23BqFW86+jZKa9fVNINXXlqp9YOgb5OTIhSOoyGijZgEPywNkliFF
h4adxmMZJywUfZzGGruhy3iDgC3GdJ8aTvqWXchWx3vCBhaDorz44nNUbpw8DO/l
te1yUjQkiME3VMojD64OQ3OINNHiV99/6LVGdHdCcs8TqnPmYmQtIH4PBpXhxiJ+
vEPin7GiH+BynLwpEIAnNhAJfLkHHAkcXATD4JJd8yAv2OhfoCcX7wL3ZgeU6fK8
CitXIoKSWIyUuJW+y/lrSsI0fealQQzU1xD1p5ew8vz/61LMV2pjJ7qoO8F2diZB
0gFXRTsySgbcFN9FKNEPKeBF/vkAzxSEPE63AdyEUSeWQdrt+7L98U0dXawI6Yjk
s+r5evgDVbsA2AHzmSoEcWXA0e1GxQGLCS1EDgusPEDkPhbpiw85ADPYiw18leCd
AN1pNLbM0a6/+LJzy7majcI4PEasa//SSWL2/ER1au5PcInPIBG8SknmBnlZ2LZC
z25cS9WZymxFb5P1kdbjSdoCLovhhIqOppOKAcTw2pZh+bvY2zwvNMstO6EZ+szk
J15LYv7KAberzHqJT6rdIg5674/LcQqM1lUFD+QI7TiBFV+9HPTdKIO/9k7CDlMe
2KJtYG8+VopjAkVqYdCtTsZXaux9Hm25+lcvaQtCwFq5GBfiiPy1YKndoN4KsCje
EX8JtcwwLxenifC0RCov2JGbx1v4OpA1NZQDcXigqI6Sft0Tud/DpiaWBtv96JMo
Gw52q+gq4UUIsA3sFL/lF+kjuSVGk+hJ5W7TgpjwQ28Q4Fz0N1VRveZ4l8xn36ff
TaBEFkPncc5vFa8G/xf2xNSsq9npOyyZaP61nHtvgmD6zCn+ls1ApqWKQ8lK1MxZ
c3g6BLE6RpA9EYXDrUnxw4jK7lBaK5TZMSKGONo0jFf3g2wIPx2VKB9HWqc5C5Tt
78AulHroZ8ljJMLTWbSYs5lcFpbKneZ/ImERnOpdL3YhStUFzfliUEAQRWRDhbIo
WLUJndFn8Z9z8GuEdqdPvEa9xrgmgAAoabO3ToBIzvugdMB8JpgtGaS1A99oRzhr
WMt8Yozryi8NBu8mODvTiBO7IMMnCguIaEhx6/8+zu+OHdY2RVgUPZx7G1xQLDB6
hvmkCyAzrcIwZkG8LJEPr21pgrfiwet3/3qi8AX4Xh0plOLvPuXKu3jMgUgpPh5F
pZfVDkj78ncVXlAar04pqbyKIH5By1r1zWrrL/rvqZcsqZSvgDZ2uhmX6CQa3pt7
7lAQAdxpm5YbM2/Igz6Ha7QARa1wy+INqm8+o1v1uc0kDppkg0QNllzj7BHhMTEn
I3gNxLzIhEBrsECR2wENdK5Pk2OPfocn+9f8edAyvXeInUknBrJfVhX0htrmfL7/
vRtOQKxabn597GeZSCQ2wNbchPC3KFXeYbR5gj1u3idkroAirqPcCZJBPJuJA6HB
rxwk7U9WsvQgvPbKGt56G4c1Fcdwsv8iuY7vWc1x14l/LDGAbCw9JCVtgLYrH37m
QNvUjt7cJDcK73mEMvfWBcZvouvlgLGHX/ooClCDTh5O8UeBzuqhI0hBH3T94LIP
oPmxVCplSoxyIoblld5o4iP2tcCgRIBIxxme0Playp9rU57jdFkyvL3ARtHG4JCs
4cBDnt7wme7AyIlgdVk/5g1QAPKxeopVCKhmsm7vqFU+9f9UpeKYZVuOVnEfL1MI
iAg5G0bgaxMC/wRy3SOKOf5tZBYKhUL/hxjei8j5/0GjoQAgfBb4uBc3LE4DfeK8
XPGpz2Md9o9DrUF4tiqxoLISzVIDioHB++7hyU2zFKr03aDItq44QF3TPFi/scng
ACqPSicHsTVE+CHHZLoGRhfHmP8T5k4psiEgSTasoO2ajJdg/z/zWfS5tQABmXAY
59nY7r0C9+UtDIXnRSjUVq/HkJ3OEpHbMYchaa9FDJ/jnE+txZBU7TwcCcBiGRUZ
0jOsG9feYgSnkTfQUvMT6SiQBDViI88uE1jobnuHRtsMKymzyyRGyw3aO4YL53Pc
EL13yfyqJtgvz9kWBxvIfIxo6RzL2YWH8aYJ6sePk9DcUgT8tpO797ZsipS+eq4L
KlJiQoWXYmGxjnTk9GSbMxfOB/FCJ01zENM03yg3wb4sVZc15AhQG2EuWri4OK8p
ncBacjydzLAiNv8zqbnj/qwM3cOxjW8IcyYCteXiW4t2wj3WYV0uFgO57lZYfNmV
NcxP3gNr2hrjDENVeWE/D0Z8SqbhbM1ChlP6fYzpQQh1XYomd31UJFdP9hofbpIQ
ZF8KkOXCVj4k4RTBYapRw07lsX218iWfINIvXhM28vqMnaRpf6xo5wVGEL0I2Ei+
G5UuxZ0vNPaLtEI2q9rhjMSWaA4yB0PwsO0rQf07MkoDuJgwqat5IGR0sbWERKtz
d+mCjjI8D0jPCV8bAHVZ+E1Lgt9Si/jr7RBBN2cDEURrx2UeVy2WX/74WSo2gp8n
+DgTuq40xQgXDYgu42PcQUpqBz9mF9sSBssF5qkNW/+UTB4Nfbwe0582Wk3lD40G
slWo9xBoQDB9aghQNlBgpJWQBf94LVHBfJZChOeyH4mxeq7K2d9kXoHSt8iAZvhX
sZ++NCGSv6ICG+MMO4Y5kkt3RHGc2Ef6qSGqTYqM1xKG5w9SjVU3RcH4Sv60S4Qz
Uu5SwjjfJrFge9IubBPvFuPrF7/G392XhsQrLdBZbggYd6354EZoTjhvhbVnr1gK
7uSWoFyfN2rhc/iFWeHxptnwPK49FuyVZaQpmp2hzHL/44WkD//QvylhhAVQg9tX
zMZpquSzkY0OM9M/sm2K12GoItoNow0qUQgsQIxmobwFfX4qZZM1SENQWdcYnV+o
omxD9h5prtn/DHOMV+dj7WH5rWnTR/Qn4rdr5uocv6zJ3+ZcJLJ7S4Q9sALTOlku
awQ4ayYbjrYn9oKRfV4QhLKFOdteA2ROFQ5NNaUXzU9TRXR4TFNlQ9Qn/3KZK47q
CisrmbHktVvTHuxdDoQyUOOq/xJ5mta8aDZRlc55wL8pSeLaUANv/GcXllLZSlPI
JC+ITOFMnZ5tQZy1ELLi2TCv8njrMi1jgAYkEmv3MJso8EXcvtNDOpXMplc4YT5F
vtay0STVXEA1tDGPmjOH+MkJgysILvELNs7tQ2pdx/rEQ/nfFWjIW49aJrMprkfU
prOQiX/8dZBX1sW76nShnDjO7H+sbrKGYMO+WkOHZi0E1RpUUlXuoYVNYSdUcUw0
GnU/8CYSdfOQb99KYLbwzea3TZ0CVHi/2oSJj/6/hgfzTnfqXVUwBOu6GQJphxCj
/0RPVrXSKyLnRH85u7oZg5TTZRaeHmIFqy524QGCbbFeop6+F7zXz7ZXI4M5r+fD
SKgjQTlXAp/AsqLHqJYt5EVGE/CrSEf2zFy969ZH0vUHgM9zVxn8UaDmQpQSpbdM
hssidk9ERnNP8+dl0F7IsOJ1xSaDJCVzXPohhaAgs42DCntoPwvgkKJxLOcCyrJ8
fBMfc36a6pn0vEekCseNZ0Ls3BbBYVxRtQsgXx3KPq/73WL+N6x98kGEO6ALsnkq
o6r0jPiJEpc/Fia+OSQO/0GKvIIGwe5mZG52NRhVcJfR8x9Bz/KtijFgap0yv4xU
yZB3KysH9gLZgAOiSLkMCxdbheLI6cnz/m1Y4MH716g0mBmwmKSiBwuClYbRCcLZ
T2p0S4sSI8uUydn+msvKWN8PWS+GhvnzvKlZ6vF0iiTuDqtjMIJQ2oiAN58zXGnG
ub6eQUd4rNmaGQwRM9vPbwClDuSYnSEemJMpR0DLDcxzmemvoNbBYF0lwmMzR3EM
5ZE897SGHuECBCs2/fiAJ5NljMUxbMIIZPM2bJJSE4gaOAszOui7TTxMLetfsHQA
J59snU71N8pk3yEBqLCbDPZBtYRrKtlY7CvN3R8XwdU+l6qT+c+cfl/kDhfaF1l5
YgHj5wOO7os9g2pHNOd5CuAOPIKvuZXkti6cePi9XQ/DKJwnsDXr8ePx7xLC9Pir
I6Y1GcKit80mBHDmrMjTimbrBGY8lEN4DlxDeeoPt48SoHeYD+5lxkGveR+k4T/e
9aubFKd15YBtcszsTkzaGfzgmGSn236rb/hiWbo0yVDvIBmccexHGdxW2hhPSDNj
z91JAtGRlHdAGQWpl7/uRqKxztIFK0O6oaUJWhFVt+y+/HkFvQTOAP42lydV4QRq
C1zFXP/rLj0A530KPkwK2pU8SlVw4hmgLtbj/r0IAwolxguP7m2Obeic2ok41qmu
UQWsy8kg0m9y9XeSFpzcpOnl1y9wWZ+wzVvXr2MGn5IuCc1/wtbzjEMvnBVin+EY
9nfjKwn83Hh4WwEjrTJLtT+Ew428RcjBYbatXhI5jJqHdl9sPOJbzHeaczKrZ1Cm
PVIVI9YWkLYMSyK1AwhqH24Perb0iuzglV8V4LJJDNW4ieMxt4y/K/FBJHfdn3Yn
wgqKGL4euhJk8uanO8cTS3QeBhzeEbN9VvGSOn1TWG9QKhFeLczcLI286YEH63f8
VzocEkdXQgU71P5mQ5bwOXrRgp11a0L20GmrSQQ7/GErCALBrY6jPs+Rg1685t6K
BXVrZg49SHtu6t1GvQKSEVfxl1VPrDcKQNHjks9O2Nyvtnz4WHvD3CoZwI3VEwAt
Pr/pIM0l6ZNEiP/0l0TP+jUMYm3tdvUnx2yimui2XqMftrUErwGkpYiEpz4Ftc69
vFhFUSEf5uEAX0E+CF95pR8KhCUqfh1da9QLL1FsUeFUzgq7SojUfEN5kisyKl3G
ZHlepzRFQrrj+V0DSxvWQKuSxXrK3Cm3slgxUDrqxgDY1/vmTsagXH5lUNq9DbhB
o/9LU3pea0zVLeUOyQzi8x3uSGXbhqeKpp6OYkkNctzwWVA7eccRzx+xTsxcBK/u
D7qgL9NbrbBW/58m6vEGZ/4mvJ8wtQVu/Ua52EfGWMy6LV+PF4DjYW7oEeAWIbZ7
u6J4rnsu03wlYv6YHq2/FOj2EiPWW4mYitVjDFDEduQAtM+qTEimMsjuiXzdiGE1
tLZ4pjnR23DV0E5xYfeEhJAvYSYjNqXddTjRMWzRPJOKQiKcIV6gWbXQMoRr7sg+
X3y6dvpcWCrtRebauBpS//+UsBIJJZH4lxfFyWkPATG60htQKeDRSKfdiyhfH0fN
tpAbxyRNKF8UiJfto4YvjvAc4vdaIJtIpmg2B+iNQTznYWydT1VOV/MHAC7ODw8c
uIeuho9L+DjY5bKy2zoKb/ddD3qwWwDTR8ZcxsbCf+xKRQFWyEMTVjhzmTfXOt83
o3CnReW68QeSRl29qlxietphDYJVRG9WICZ/7th2rSIQJESSuHPlEMIUX+Lf4Er3
MB+JanhqEiL4iAuhZRJOOFf8ziT/i0255embthxe1O9msQtaAC+k+g+k6koGoohR
yl3D5SN+Wi3YMxETT0969Hshzvu964DxF+5If/gKtCD7b+EDTFjmJ8EEV6QAMYzX
Z5BOvk3ODJfaHKeqoFU6etBLAKzlyiSUu56TvzyhsA9laAzxhU30hZODdlLkMeAJ
I+T8KRr1+oeg24Egr9zk0BLZW4HDfD7/3RP7w1UPsTtjTGC82bNGcROaFcGqw0gZ
Oeq+rX3RhFx/h+JxxTHDC1v70MGOhPUiphFPtzzadzvBA7qs38EWwLxtaMYGO2aq
k9Qtz1kr0yQAR13GeINKMI8+idGmeVYGMlV8jKdeDeuHt4sceTRJeOxlxkcPQATa
8vorTN5ckklpo1UHepB7THfkAOm3VsQivlaHMBW2/rFmQx+3E96t7vWQ6CWSNYOE
ibj/PC2UoYNfRPZWt43K2f73AxGc7jlDvXbjIQ7OW6+9jtp9k9U5QyXKyYy3KyoY
q7+/Mk0v052kszyTW+eivaD+E5r5EmdkqGQ9itRSEiGILbRSAjG4PUYwWnL8quYL
qqGl+7lD4WyXr8QKSwwZYN5T2OXDlfw808PVA19AH4RaMI1Nxi7wBd1Nh0N7PVwu
cpNdmknWdAQgTy9t7riEDhypbUABW5DlH6HgdCqL67DDAhxNigo1LPlx0l9JAbKd
jG3CVzu+y7bmqfiiPjLHqnexuTX8/GLMgV6UsMP8smIl76W1zaROQ42B7tNo03vu
2fwClQSCi7SuXa6s+uemm9kHHsJhm69+1DMq135qBSFIVFTePcPU4suyw4SObvJN
Amk5ofC5uWrV05s7sXrBZ7ffGwHXa5Vv6NX9L8pX7ZQ1Mb/b/8HBBe2VNV2T+DGx
sLaTg9PncxpM7Wf5OIeIBbORYGlhRv4ndN4mC344um3q2weCt1Xo5A49pbap+Bnz
vbTaJ8l3hmfyQYxSiVcY4BKVyCvwXWoWBv9Geh9fo7IVfjMXJkUZ2M5FRFHaRzpT
IcB2bIOHVDy+YO43mR0Rje01Y9vKvMXRrLIe8gXyVYAiwuZYJmfX3pf+VxMlJr7d
PmvBd+Z10VhEvQY+WqJ//rcU3EnGJ0gKSg11UHY/jnKI4UweNHhDaHvNs1LQ7vqU
jO2o3LQ0/A2ClD2l7iPMTilFVDdMiX1MPVvbW48qGrjya6ZtzDAk5siCdrc5w0ao
U1X0IoaX9pTiScHo7xOXxwBfUqYkjquX1oSaGN9ct2wwE260l9NNyjKiYLiV7+MN
HVNvPt5NSwoDrCo25pp81kEwSQ9b5hUm1WNqH6IVzk6855qk+2p3joQnYGdm/yfj
yGa84JaNDy3khUtQOT/T0lseWg69t1rWRgzuefiKaiUiqAQZOmeV3zUN/FgaPrzC
D3kpEz6rS29sAhK3H243nbCOiQ5QOFnsZIdC9ExbPsmB56BIgsFi7z1rNV6dP1rk
OST5CdLm7f4/C2WI84l8JWipnYHk4vL+uhaL0toKyNDFf3IRSaXUJXoYKQjGRUT5
65O/2yD6PHD+PE5UpsFPo21DkI6xA1pb6ZUSEwSc3Wnb/fvInV1eVnvD9u2MT4uu
44HHMK5W0rFR8B6u6ZRb7GCkD8JdXUjT3KVxNvGK62ppdRneVyxxnT8Fos57TOGR
SML352q6imoUWuXB8Qkg2skPuiIC7t+HvVkNQit3lboRuqPzhfdWAExny8wyj4//
yhNGkFHN4Pzt+jiUfaAXqr0sSRcdCXnTFKAulqw27ffBsZOombXqrSil5I1nFz1I
N9yQaE6fUeH08d7HD7JJZfFmtvjTqpjjxtLKKhcbDEx7rhcJqwefR8Vhjb47U+LB
VqWl+5C1fZ/ynaK5WU9zYvhDkpFda0+SOIjdcM6xMY8IX8shjt3WT7D3hyGf3oQF
tYMTdKTFGz47HnuMrSkOnx4ptIvzzfAvThhKeSIDEbEJLbcc+/bNAULczHlpr9kD
qO8DtC/FXvkKXBRIgjPrXmtWDFWTPQzOhFtDv12NPf71nUrNB2auyOn2hSRG3IN6
B0HRLEhgYoD/RQ4XUHrUysiNjHCeL0zF+lP1u9mX/sBwzTJN1nO2/fbVWZdrQr0y
OVoXbTjlGzmNYi0HXAotrcCgW1PWtLXKsXK4PKWq4Uhr+NOZiRJe55HgCZVSCZYA
7aBS0Pt1Hr3fDHzw42SXoWimnmuMSBiHOn8S4yqbzjEFBmH70SSUuvzCXqXf3Wlc
bVKe9Dxp52f67thXX0/GwQZS4Gz+GQlT3OY8BDkD9ryekjpQWa47pqH82Xo+9xpU
lTQGAsQziXDfDctoxW8CKSHn6Pgib3TK6ysxuJFLpu5BMsO3dtUFDLAPlgMC3W6v
d8Ui4qIcahFPISoAIC1Q9+Oq/PjFoKQhJvE3jwbHXJe3nr8vEuPyaUPYp5pjy6pG
uHVCiW3CgpSawYkvkfwcT92Jd2ttP9GOVEMQcwek/UihMzGgxDmBdtmtTvMD4/vR
3AbVcpTv/2ADTGvlUEanr37xc3mVXx2jon6EGM8SuJ2Q6hMw8+K3HLMJUrNnoi+Y
Eun8BeqkwbqUXdGRUU092dv0i0a9Pr1laiSLGo94P9tXl0FLzbRr662F4Y24naQZ
/R9+VwsUlZ2iDUSR1vf5ksvFIlug2jEH6L+l6g4NSBEkck3ghXRMCBUfgmmQnXhy
AuKKl/j0kQdd3Rb+FRZD9r69Nwt3L6gtba0/nkp6TYqcmB7ln5MLw0ByVhplPBWg
492q7pCmSJgBFGbMGTHcoNbGRX5B38f7XQ2/gwdxLXeFD/ulAknikDO0WiLK58lN
GanprVsv9UPuj45E0eiLZabOY948DY04TXV07/ptaa17cfcEij7dS69N9KrOWCFB
WVmRa2hGlh07b2nIwCKXe9owpD2SvfsBiKK7f6cB938UzTEallkrSuyG6c5gYhRq
VxeYPgWCESWSUeEJLlKrMQJlMHt9kbXCMQDcYdgxfe+itpdHi8GzCar3PcBFdzIB
6Dqn95ZDY5Zul5P6Wbdo0A==
`protect END_PROTECTED
