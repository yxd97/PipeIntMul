`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2ORQWng7HHgc5CXrNd37ZPOPzOMwW2yYuihGooypKRStsxOIqtSEMbh43R8J3Hr
JxU1xBECKLmlf9T4znlS9Pnqz3/4HfZlNj1JdtHdzxbRv95mVKmqy9MdXVf/TivE
LHOUAnqruT07xddeDu9qaDFA0UgOXwnr46PrYcF/EpR3gOF8S7/AKaaY5kYl2oFs
5b6dhC9bohSESDi/0d8KLk/Trd3EuvRdGYWKi2c7TJGKb98CkUB2YYWxOrf5SDyR
T5UgXW2q+pfQ8ehwpsBwrBu7ebUC3lV8aotxdzLLhjTylCdDRqCW4sYKF/IUQWPn
3HLblAwRTH4i2rcMRjL6Q1jU/qKwuV4Os47T+xQ4Houm2W1amF770LgIifuJqtqf
l9pWhLFiVWwPIRlZUf/tEfKwANObjnyxdv3QX4SyikS1Lj2Z9TSeYjhVYahIwLcu
dLDMajGp6vVo1v705yz2eHpAdWxiPELa0jIvF74d8cHqpfgd8UKbd9+DgOEop55a
`protect END_PROTECTED
