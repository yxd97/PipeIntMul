`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exFR7/Lv4jeGe7f70oDdx+UDPevLsMNtSxIYMz4HsDX8exjaCUf4DHwQLpZzo8f5
roOqQMmu0CYC1OE9wtjv2SAYA0I5o686OwshgUTleWln/x+uDefgGOhpTOsCPAwM
42d48NGY0OROjM9M4r0ZN5SOSapAM2Gljxf1u5GYoieSntV6inFy2PrCYxR96yb2
+Igh2DGjDp31EKUXmmtKEafJY3lBDEQgjTLXBT+eXyhO5Sd/TFbCTOrznIF9PdYD
RXkYwklfQfDsnRqiXjC47Bb55KKEnSTLhWzIcFuSavIfnFVYPq4qYxphN2IHlumM
N01aJ9XTdP9Q6YIJdrOXYW+XY+DpFMn8aoNuEXgdG148zufUKrOujO1Az1U2kPnK
v+6AfutP1pDLqKrP+MP2DasGYVDw5nGhqg8KPfNOujRiUGTBzLBMYpZe3wOvPH3U
nS8notSfZEV6Vu2HHqxXhwIV+hynyxKv8h/FiTnBL8kLwf0Pc5MXLKv+PCu5h6Ns
WUgZbh8EGEW8l9L0t+77VKTOgYxXmisgYncArppyzO9g6ZOHKHiTGgMWP+7Yfkpo
ZmkkFTEG20bFbpB1toU83/mJeb7M/QfyehcKB/h5/VjnZu+tThCwK+LEFy5sMo9r
+8iT031S29upAL/Wjt6/GQ==
`protect END_PROTECTED
