`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vlcd0r4Ysq17Pqm06v6g0MJW8+wdYxz0Gf7W5tZIKIyFFWqmb6lmewwpEU7Zm+y
vBFi6HFB2YZOwGgWRDSyE97eqXdchELoTXovHxadY/gatlRm8WXqOj3pk8xG06ZR
hveRB9rWjiVXxnsDgl69Z9gq4dGblInRmVKUqogktlvSVRQWJ3Yiqp7yLcdqxA4e
TKCDan5D1MbDoSgU2Od0mT8uMiuGl1cLXXjOp7xh1hc38NaN/sevnERW6jW5DWwt
kmfOZIyiporrI+aT+mfU6xiT0N3SZjwtfdq9+rDhA+wzuGqCpAw559JqjbshwnbF
ceMe/s/1PboLIciweS7Epnx7RaPA7+Na/UHkvxHKmei9AG8usbE078lm2aN04dow
F4qGcuGrqKUDb56OWgfOPOlOcdwRkXMNSjrJYhLur8M=
`protect END_PROTECTED
