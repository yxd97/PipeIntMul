`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQ8Wk9nfmmyh7C6eSPqq4E5P7gnwjVk01h16ATvCsWUGU0h94kz1QYZQnHbKru96
p+x0Vm41axoqiOFMWxHXPQeTAkONJBjUvdT16RlrzmbTo/a9DNkpr20AXc9vM6AF
xi49pbsVXJNB0g4G42RfBTelxYrN/7dIBtlOJ1WUGMZXQzCG+OeoFJ9AayBkLytX
wBp4jgxXhjLy4kIXgs8h0fnzYfufdGYHirjS0zhsazMdC34XKlUApNr3qYvr4f54
qF5h22J+j7SY6+Sa6bEhTmaJ8BVTkRsRKHtPX/jlyfFeqVSrCbQYJJc3e6lZh2dQ
8PeI/2MtD59cpGPPPrHM6zt9yuKbyXz7tUMaSYZxIWeAaMutXpD0QQpczLeWFXPO
i4q9awIe67RPurRLyPcZjQZsO89T8ogSCFUwoA0/cZyURS8TlaVPkFPudPvgxKN8
TChrPvPL0Og6daomYiEi60vfbF+AmYhGAmrXXmji4i7hJxKgVyu9EEEXrsj2+xrU
paL5Ai8JWzqtkBH9wMwheRxLLSac6ciqW9/PRWmiwdjBOZUqtPAMauM10M40Yn+h
dbet25zfiBrg3fh1GYeB6c8soam03WHO4wPGJPz8ZkvvAQB2cm1oiK8GluBSLbsc
/IBLLntULxEfNPIumvvaKTA2QxJClK9JAu3pBz7oPpzqgBiS/e4oWf42WVw+hoPh
MU73MhG1CRreApdH04a9OpX7Zku7s2wNTuiFxcTHDOnaZifvHBw9/mfP4vFVsLFi
WxW/8gqsU6bP1D+5UP/moCIE2PwZMQlsR7Zsl6q5FPdtUtuiu0tL5C48Ujm0IMe5
4a/G13bg6pAz2kOsq+keiL5/u4leSrKizWpCepTp6/8eI5Mz4RQ1SHmON8O/L8S2
uoOJn6cXoc/S7q77U3uIwLV1GhajUC3/6JwxExhpjgQjN90Vs3UDWqsFQwSZmmzP
NNM0XUvc4JvvLKyGdee5zGNVIyVhNtfDuVPcIlRVMtdyBBoVprE1FM2ekd+gMIKN
iN29JROnYwqSFPpecDZ7jH9G3Y+vI7zqPVzgbeCdYOhtg1G5y9JxN1OckalUmNeW
DTw5HheuQ/Dab/gHDhXSYaM2TD8xAWgQ1tO+RURPxv/H/sm+oDXK6HrDjOPrHQ3m
i0kNrZT0Y6i2AzjAQ+QvLa10oZj6tKwtcuNHnxzErAH+G0CUROagM9hwWdKUed2l
uRzdoPlHlbO/aYwRfxMKutZmkji6XG2TVC9XLA/+kaAplSO7FK/gxM4SuPywAyeP
`protect END_PROTECTED
