`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EKwltxHeEZk/2TLjNQ5KCpXisf0BCLm4zuFuqYVSji3xsxF7lL9hKZg+BtxkPQRC
uyh1zgVUSh75h1fsIfvzPJ6gMwAGgbtm5xZTFnXUaI7WULwyutRb2irl2yP681FF
KuLjsmmZ2BbS5BNp07W9HMFIUhC7PmivNZGYKJdHu+eF/9vr6KfptUFWMC3b5lhs
tMXJaduCFTQgWp8r/bAse2UHqPRl5yBXyEgcAtq0Pnkg14S8y7bpkL0S+uECWbhN
xza8amd4fUYScxoD/laFdVdFKBSkJ634zyccepkQlvUoJLHr+QR+2Z7D1QQknISC
dkLjGXMqOHv0rzH4CcL+Sf9yNWC4EpQ/XmqorWI/tLwg1LJ/v7l5qwXT/Bp5FJgx
A0ECDXuh//BpxyJO0+Wo1XIYV5lLNH3XBnQQ9nmbbu5jsH1ayQRSfkIEymf3W4yE
iuep6qU3E4HCTgOw+8q1dLaWhYruBCZxQwj+KboiK2BV4TIvgN5bJXV7ldZ9MA0T
hvdHHLTuaEOOBW8B5WiDW0Lkebw5CklYnJuZ31Y2UaiKM71FZEXvht4ho/VeCh9G
ig9MIPHmlO0LD6rHCcvUsb5t7F+mgo7a9DbFKvLlthqsHAm9PNa5SZKvmoarmwdI
mE9ivvaEAN22+auD7ZCVR9UsoHIQ8xENhxRGFHos3CX+PuPs3PL7SNHaSxnT/r+K
PJVp2bukE9/S9gPu55d5FYLlgjBI2zuzMFRcwvX6JejPXA4vq1ivEMhbTzlztRcH
Y3/4SiESW/n8NzNHCq7VNGjb1AKIOkjm/l2GGRwkzsKd6vqNI8mU5cscSDj/vTa/
iClOZPjp/dtznw8LPFhdfhrrYrPNUALjdjfrYeWtovSHk6aZI0ML4f7rZykBnkqp
0L8+04XlsBZIN+QN+6sNcD7bPJ4mbGSNM2iBANEn97QavswkDC0guZAHBOu1/4ld
`protect END_PROTECTED
