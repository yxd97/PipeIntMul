`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2xsii4Xi07uOZvW7UCSHm1APhSRqEhVjdNrr5M+FEkoIHF9vcNl5OYlNZzO1IEN5
R7pw9e8Kq6JuyBmUbp1aHWyd73SOirLIktcRIWR7D6GyVdcTF5DNGdqQKqjM+ljC
n/avBSCIqzpkmvTglq/BHgmMvcL1sPjQ1witDMqB/nkfNBif8ogwKTcTfgpTdkaG
BX6pJOy+9kjg2ZGUeUAwzTkEYVhXWW1tC4SbLugc4LCNtpI10yoMOIW9PJiWo8Fz
lXFfh1aMgGAyUKN6x2KGXSi21jJ4bZfK49iuW3yqtkqlw4Gb7+P7fyzXG5KxPZm4
llvAiW23aYUXaTvicfjYtwV7mU0p0aoCSuQnJc8BAXYPpMU3p2s3xYt681540s+8
oBaU2PXjzGSNseDXoAocY986nBvIF644OvCkmb3ZzlUsr+TyjpHhL/ALNDlY5Om9
/RGWnXtpoKq/OKwm2Nav9HyWYWFaSluDzQEyRq7bv5I=
`protect END_PROTECTED
