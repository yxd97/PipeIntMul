`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OuvaBEH6KhaeLtgHX9ZrpjU7HvtIZMvkkqxT9i+soECf2QDtbfCnhP5u8LCzNN6p
xUank1ZWri80kYz/vGcCLb0eiR7kaPUtHiQrEy7b6uAg2YuBWF5nFD9LztBbggGQ
TtoFyftmMbGQIWIlISurX/fYf1IUVaoftTbvI5EgW5O0UXJ3fxxgzTkarYbBliu5
qhf48fdPy02bwR8s4eoSwsorSQPDjG156yyyW9NLOj6QeqCDKh+pOI/me8gz8skd
plPC3S2qtrh5eBy/UFiVUC2QLbHNWdNxAA4DURo1aEte9nLOzLlga4YGUCosne9A
1kp8Agg7C0lWYujxlU3TWIhmePDYgk/zVbnkCboMx2Wh27ovR7Uiqq7LT8LnJrM7
r0PtIeABzThhPYZo7vIhF9dxQ6gyx/+BZPMTQTek+fJNooimJCoaYFxsr9f/mp61
R32iJ1TKt2mzIMjmvxnTtAWd/5ACsc7/wwWqbo6Zk6rpNpn/MKkL7pKQBNHUFke+
uBMlSiYwR5wQpxLmNLwQRkogT5QkS1RkH3xgQYvcXpp+rCVr5C3QehKg9ok6hjCB
U/FvESrnMP6786YZGFfLWea0lF8o1FXxMkExvpJLn2k0FsdseuucVflBB5tCeAOU
wGoybBP9gqE3QMjbTVSEfjflu0zP5H+7ooHJTKFg+e0hoFVIbIUIGOPhql5wOM30
NQkjzNiXqKaXrxwCJyHucEQlzElA/e4ihYQT/tImVoLoz9PLHVqXk8Y5oQPtBbF+
MGgLD6BTBr54Y+ru94dkz3CMsWKIGrKmLHIhpFa41v3UI1zqPJQTwP0NtMHdbuOd
A6svu3QcF8O2Qa4QofQPT6DrSO8ZYHAE7mv30OkljSDRujFd2eccjOHn1DIVP8KH
XeT8Zckis2SsZ3RXIkZc3Rrf4QROQBvLnfe+skMlLQpot371jnaks16OHUp7BTvy
aU1oABP2oCAHdicchytbIZzMKd360dNR5tgGSzX3u+wU35CvgZGlPCSUYcXJR0zo
`protect END_PROTECTED
