`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2FuHy9TOUIP3oq00aqi8OuWVhINLbrccxfD14ujOgCj4vh3HMourVNZMrXcmX3UB
Yllet4FFsD6UeKYl3QbHpqb74i+rJRwAeoitq/Zu2gkpOrFfVoV53c/PF2OKwVvO
ChJXCCGl16XVLdV9gs4U1ZV4Y1dfNUkDJcJ4ZJoOatZVqeKp7+I2gvmz0y99LFW7
WTTg2cbGyBrxXyUA7gWbdFwsilb0j1IclFoLAphXAZofSrcyDl3xXGcveBqaYjUa
Rz8AY/Yk0dpAxedKZbP1jMjikU9c6g5mcMDchRlNtJ7fs/1PjD2fyW/at0kt4bg3
OKUpGAJrgS9rpnJEtIdY33rnn3hmv0YhnuPyUdxr226/q+hBl4uZzQYGQ1dPCKKG
sKUjCsIWXZIry76PfNhzjyYm8Of72JAk6sIPNvkbBklv0pCecW0c1KMFV9MsG4a1
9KNw7YpLBKvmd3sodHvjrnCuMDNs+WlM1KdBNgPbwcX9c0011qSL7k9RdjTsr8mh
kLFeoZhhU0x/K26VmyQQjlu5bjr94TtoNTpCJlKRZwAxr3pB7ljwxx2rZzMPAL15
WBc/Qefii/SxxgUcnnsN/fOCt0EMAeRVXFX6sTCHc5Q=
`protect END_PROTECTED
