`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocDCmraPW/PE1+RH4Flvvd3YCfME5g7RrkGuFrx8zF3DYasKfl8j7/mcSMSBPP4H
aODoxl4bRXphXkFRQRBfwXYSFqPKIg8e1KRL5p+YP1r5VlLjlCzDYvkSTLCRjF66
8owqJdEQF8pxsK6alQoNLbqU+/c8tGuo2RCg8jHz0vgAUgVr27K8zw0bduBOTxIa
FxYRjPsxs5tGfJwUJo80QTcImhkSthd8I6bMXt/NFdA9BoRD6NV0taioDI/9nK3L
hoUL3LuYcPlKRCMJ4xRjg5D0lfap4c+kZ2IbOEDyjNYuU42IjIyM4bq2N17Dqsa6
na0q3WkdiqpRpYtJqBfXE7xDZVIHQN3SzxZ3jtl5USEhHdE1BYBbnEq/U7gQOLjI
iG+p86UvRQf2iSj3mgKfo5pX+MKewIORDKJH1JIejfqtKlpiAN9NgJI/QOv9zFvd
9DPlLshHyVZuik+NNk+GtqUaFraxHAoYDbK6QWiz3dKTMgpltY1JjtpnTuJzGedK
`protect END_PROTECTED
