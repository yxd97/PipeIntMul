`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZDGIFu877YL0Wy4v35pdEt2iWcuXId2lD6ULZ933kugsa3oEq+nwYigKY3o63Wj
4vE5QV/6ZmnWmPW8uv+ms4iEiQsFAmRikkC0EyrTSGjPadiLaTC0SNWwJM0MZDWy
fFHFnD53KGBzljp29kzZ426b7rzDAOndP/mpBathWfeFJ5fpymOWQBZV3Dr+uPGx
Nujj/OKrEl3neEBDlhfCSIB576O/7SwYKH93JGBm2JoKei3JlW6K10g0v7Sj+rJI
6I+E53+xJVOmINPprDtaXM0g5xdwI2VwFfMEcBXf6m6J/5p/Ev14u+qDxoitqScu
cOW8Ye5/9KERccraEkQbzaOvg+IPPXPS1Su3JFGH+7Oe7Xa+Uy08YDjXmD2HXICR
wjUvAgLQjVPNh/XaqzdcycVhip3obG/ydrFCwL1CBogYIkBB2yxz2XaVuTRhKJs/
B5VrxC30RufQNhfk+gzs7fjV7GE5D9EeMhVrvK+wFfaFqiqXvHCSgsR7aWDRS3SY
dLopNjB907Ufj2yPwr8aTFywJwrQObl7iZd+jocDbpu2llebGYCgMBX+i1PunsDh
w5pzlW89EWBwby+pfeOFZ4PGCHGXVWtvcq7qT69XLvhmdOBU6U61HkpU02W2O3Rg
1pADXGYmzV0ZiRsN0fV82A==
`protect END_PROTECTED
