`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLoWLCpIBqU/e237M/Da6YuyQw4XW4WANpYXnGjP89XWmLBQ07qA2em9L4RTzYuw
xYW7sN1i5lfj9ViTC+NmdTcisIUf1q0Wq6BLfpXEhuR3Ij3enKuJMAZL0oQt+h/v
vTTFAAWirGs4ybdoXjXCeD5gFEVBiMZ92t5VUuPC4kPMoCMW/791GTwqARJSmycS
+0eqjYloYmnQHbmURsIYtYwXxMY/EJfuR4KadOO4yWx0MOKNMXxELEvSYqfiPO3F
DByHDuwpBDYNcXvl57Nf+i246LncXQlAoylRadEp+g8H1ayicCyDxcbTgtkY9boN
i4ljSHjwujpjZbP1Gx5gyKeWw/NdjitWxf/kfwdv0vy/+2J4RjEHrBRcJs4DUZWm
mbfzzjRLqdabS03v2IqCTM1bM91uErRQHsmM7gn2OjBQpxulJwNEu6p0/zNQxcEN
Eepk9rnNPnQd24zJJfx54B/Ts0GSTjhmtxFL67G+xEfpJ7WID2TfQqwq7sf+kWCq
WgJsPCGTEvER76TxhAji0BJFZuoCkyVno4RKJbdqkyZZKMoz8JQaakxP09DxAjuY
mex6GSqvUJCjZmX6Sp6ZgwpnNGH+quiIgkChFwH4pHKs0FoI7Mm5B7VHHt/Xqwtf
6GW5HoDW1+g6oAm8HM4+Oum7AhDF9OqcMlnYmFWyg9gvq30nb9kUDgH3Nm1wDJSZ
302PzdE8eSHgOiUpz7EgDrLWBEDo/Bn7OfwLhcvZGwfrLXelJ9+xvdzW3qkQIcNc
46Gkwai0l8N/zcf8ECjaDVc0iGzDL5B+gtBROCv2fVgZTa9tdfbypoavcccchux7
ED3czAxkEKqdMjJL9+YRP8TOfKhmjDyJNdUEoTZVCz6CMu0+nyO6pccggZdaCAmG
sWRH72ZkB5sIIoj/Ls7enoTmntyJSt9hf6blW7EWm/wod+rt7/rA0F3JKtgDkG/K
`protect END_PROTECTED
