`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sVWvXOtlw+ycaIgJhT/izhkzKGT/MBDJxrLboo0ZdxTB37jgN7Xn0iuUo/SYzP3f
Svop1I0Vd7TxRNP5BSG51CUnywofpohXjbpyWLcFcphay+E+k/3vdIl9VhRLCM+h
OIz0uTUUOtpmUVuUoMao4KGwMlPPidrpkzWXyq7X9g5IvInmHlVhsrxTbfvS5ZQ8
eWw/9vQ1/VkhcmrSaf2njv6ng5YiqKezw8ejjFTFcDNCmATxuWJG1QSVgxddvBnS
IE37kJYt433CownIDUbOrS5S0znzHUmqS5Ws8XUaIupz+zBqy4ciFToFTwdfS5j0
cA1LAXlsH1F9qwQ8t5j80u+da7BQkVen/SncGxbz5YdKmJeROUU1I8pwtA0dtqof
jRYg9v+F1bvkU5dWBhcMlTc1nmN43hMUgbbcdzkb/vw23g4rcazbLUDf8PlNvvKC
WdpmXYGtFQ7zXKwqglPp3uYaoj5fReJUfJpNaMQmlNuH17hhshhtb+hXf4jnbR7I
dU1225i2SlPvkKzEMNs7XXRsydo9c+h/xPFxv671t1TPwhjyUuW1YdnnoYFvr3jF
0jajLuyNjv94M81njWJtFFHCOLF7LK+5C2HKX+z4P+Q=
`protect END_PROTECTED
