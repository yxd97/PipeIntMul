`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQ6eBrbMI30MMkXf4FkKiUBjTSUPVLpUXoXbrbUEvdboMvkfkA7vLEAwGjJu0UbK
FT01Rqeg2Bsg7ovpSEEVkNzIj7roW5oOUbee5xLxzXff4BZ2UjExAxq3LMlro7JH
3qiHsdXBSdD3+aDgYPtotNSRcw8H5q9OOMe9BlELwaQv3j0yn3f6PP3uSZfDxe24
+UNb9KnJG1/YxoRaelrgN4has9jJd85qswrGkCcb2iHk0e34AvoCc+ZYxZ4y69C+
SSHMxMbXU+SPhLWOLwASY3cavbsjDvCt0auYOvtfEEbtQlYxDEHOjz1KTsbMHRlk
i6OqxwCkM25oP6iNjDcTB+0xVGVizcpJbwAKq6RtTWlhpU3wzIPwx7NyKUtbjqCy
CnPckeDwGBEA1+WutosI9BUsOB+1/0lNc8NZ4nKiNEmGlCAI9XVCz/z8ellxU2+k
qMXKuHkALCvTODtZSaz6f8OsT+hQ2EiDNlJZ2S/ac2ppLA86HqBG1BPyf6BZViKJ
`protect END_PROTECTED
