`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPxP0DuU5mIt5UF4481R9Fzl2ydrQ3X9LVWxUJJN7pCTURRlvCaW+X94mcym9iVB
fRqc+0ksQKFxK7QN0+GBzIuVEV8i+xR6jsPSuW7mxPxVLfygSIAPiNh5Rc3hcDGN
unGotxaXWbmNwbv0eDAFUda4JfpUnJPiQy9/cG7LYPbfjqh4NhwGm0wrGCi+M4CH
J5yB21uEnAl1wsTTBl+wwNs9QgBt9nJKuUCH1G6egpS5mcEb8YZ0js01yW8zVeZl
msp38qf3LS8BJx7UWOqt2uP9INyyOtczNA1GNtig4+NBeWe+htuqDpkp/Hw6o5eO
u5chasKOJ7To1qzJq2nLQE2tMDWdJQOmq9AGqqdc0v+CtUUa4X+0faQK9YMFw1XR
35NyF2UT+H/WVsSqXdgxhvN0sHtuQU4CfBXeTDViv4IjVVFRliDtB79cIQ5jiGfO
9agAAwmekQQ8M2OBPCzKIN3nPHiVo+RNWf+Rk1d5xyPb4bkWkhpZmzPil6nzVAuJ
l848/zLskd8qP2B3XbnWJYkRUwKO1sXRBA5UN2NL18ccTzdYgmJ8mvPRe2VhB1+Q
HywFV9QgZowYgdx26XhrNA==
`protect END_PROTECTED
