`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+uqh/XqiUfo+OKhf3F5JVh+rEHStTPuHNJfMyz/naeekC44jEgFBNBbBXYVtc1+P
4je+nLhrF133ScIbPgJBPYEr90xXmUEKlt1Q3XjkdC4EAcxa2pqIHDJaek7anMgR
jfbZuYtWs1W2PAzdYSctWFg8Q1T2uBqsmDq8Npwltyh5PONIDYwINMGDfjjCvc/V
o1kXMUTegV4g4Rr3JQY0Y2QySIZxXo0N10d17qNMSTLDMjXqEVeFepCitmxsABH0
c+8tLkKV8ljQCcV7fQavi/ywHfgNC9rLKT4MZpoO7urodYLPQ2qodrQAWmx9Lac0
2aG7+9qbYtRmY3DuukMfZw==
`protect END_PROTECTED
