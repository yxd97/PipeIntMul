`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRUVEm8mtMO01powlIo6RtgyyeEzm2dRrCok7Uyzs9UppxLNYVw8PVaCU321D5b9
xSierEpv9sTHgFup0fIkD7Q1fiMWNP01ofgWD0yTRwvhLyr/9NkRJ38zTO8KE1S9
lgCmb0MF4sZelZ5vmTlhrMYzg4+9+z5J+0lSWfs1Cu5TPK7ForjD/ZQ9R8os4dvh
F54UaSqgGvU/Heprf4GztKUMVyafm+hVJe7NS2Mp9l8zQDjR8ml0J9IpN/0FRac0
ey+DzbAkuGhXKvzVoTja4SRbZJjgXO3+qXqPbbm3lxpcK5DR30PRFIjG7s1S7qlW
qOC4QQDBIihwYRyR/oaaFACKbA5vw/+EocyNp+QEuZQ1hw4HMfht4na76G1ljCuU
7BAIALgm1UqW6+5KI8kHgsyCIBLhcGZBXW13b3NKlIM=
`protect END_PROTECTED
