`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7D9oqveV5Uv9kDSpPFuo0UdUSfzqlHdIqoq7UilfVpieqqCPuk03gSzo74Ms2PIq
+WyGamevqLmzB+8Mp0VyN+67JJtunNLrZ7JhM7Twc/3BrYFYdZviIotFs0HBGjyu
TT3WcFyE4SXa7Aw1Rm8gMWvghgYQS9Xtqa+qbtj3I6ygxBVaCdiVxlXGTTgEpfEf
sSX1G4fs1wMKxsOEPwxcgscE4R60uNCLQm8fdpkFulnLIVZO3fJ3MRzizMHoCsTo
/vQVALwqFdoWMkGXA7SQ+LHHx9nH3P+oApCZ2pEzpqubW0cvmsRvDD7C327eTnOo
qXfCMpmK7P6N+PXncKRqJw==
`protect END_PROTECTED
