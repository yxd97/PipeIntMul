`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMgx8UtwtxGn4sYeFb9vaeAM6Ci9hNuGuIYnAyNMEmF+FRbEIccWPbBOnB8e6F6M
HevzpSfN6NQJlytZ5qgJemRHlIjXPjWIy7/SdJ7eVyoAuK7XCqZZtWS8kII5zA8u
m35SgolABTlFJepDEWBpTPIoFqH6tbKeBRLaw+okrih3ZgMJhBEj9ujiegOsphxH
WMl0V/6GkhmhM59x+w/0gmHNqbYsGtWAlT28A4ULlna9ii2N6b635hFPs2DvTTSK
5sVx97dOtWxQliNBPW88U1tPSwJnkz8KaFinouHUtHjWfubdzZdKmi9u1oD96QDI
TWD8MF9PeJ4xnCAvH5sQ1Q==
`protect END_PROTECTED
