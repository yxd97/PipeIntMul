`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XCqZgcKb2iRURnM2F5WT5j1vXz0M0kG+oMr9hkPIsTf0oE7kYqUFM/UJs322Uqjw
AyP794SQ5sD/B7u9HKkwSsIkHsaA3TzL2ZRe7OEGBH0q7G9yrUIdT80EPCLpYNM0
0EAOdj/eN5WMCFaQA/ZHk1G575AHjFRwv7tB69RnGEgTtHMu//cCzYllsedSUtqa
FCDdwvf5ABqZj4rehkWcQzu8OFk4GtHW/5hFnsknswzocZPWXwKmXw4VKNEM9Q2d
NnLw1oEnJssvMQqa7wfp9doSdzTPTvWUgN9AKiNkDCbqyrovk0/cSi5YPuTA0Yo8
+L/jTcL+TiNek3OkDSGcURpfn8LzbUFCoU7voTECds9u1HPrxArz361SGIfvIhR5
wsO50r9bOn9/aelQySYAge6CC+xm07o3cxfEYe+1zZ/WwetSbJ5gcHjDWxhF8HlW
UGhsutZw7ken1/SXksZKpZiOZhr21YtQHQujO+Jn3hG8mZNMciSm/4yzjd9Yo5R2
exbgMW/JIdKDXmlGNldJjiXBG7vsBFj30PR5o7Cozjq7okqdDLNwAtu9OT7LLvQf
pLnj8PX5Q+5r3z1y6svdOeddSlfiTW6/KnlwIsWuyG8zAlM+uVOmNE8kd8ISSZZT
P1dwCU1+JwFxxV9QnePwKzRjXnRFwX9iArZhLXkfZpSn1l03Q3h+6qAf4+5ZRypb
1/b565c7ROcoKnAIHP/8Lb9QHoz9BSYAsLlaHyx7s1oCM+VkUe7FDQG6sHqoFp5E
1fdyccmgrNCn2fdLqln5Y7UFBhSWbzBsEbblWybAGuJzFLmXq4vNbl2TQ0DGy2E7
T6M+7ldm91r7+CSUixUMwqcB/YGAaUPDvGNWOfrRCA0VbFb2hpT+YZKII5Ll3MNs
qkhWPwQH9WDbwwRmApj4xoipORi/dULKzSsFTBqRDICtj3dnhtE+qPdRcVJNWwVV
pP4wFCFu6iLoaQhhp+j9+ZxbHDDjDMmwGU7mxeSYqaBmznC6ZkTs9KP9ngfBzzPW
qUk+daBoXdb3wJ2z+CDYuZDRKYX9eomDNu9R5LWyE+wLu7LBmH2zo450m6B0XXnO
P1EovU6WVpjcTA/0fkm2Z4DApJzbZYfiSlYJzwzDGRkAa4I4ljCqPPfBK9wy9nM4
fWswzGv4jvcuEmXEPcZUB8uBMWGRnId1zIjLIEMilfxCs890okw7zfaHbXq39k4j
i2/hYPHlyt7Bl7ORzqwDtpKinjebJiKJsWU2uX8xQxUCXH793PxbjXYRcWe8Vccq
rkTF1kcoZVFK8KmCrNos+5ZVOlB2GXZ4OsZkavtyCmBQoZxzrzyGqdvSyAacss10
P9tXp7x7fzHdvySWbn5hjV1gIy5bCpGvqzhj4d00bVnYVkCssNZ7yof1ar0MLeSQ
l46kPfKy+yMByWHqmRv19X87bY1D8H+m88MFIVugtAPe4HXS6qPc433eDplhlNdx
X93hErFBF5k1IaPNwh6xTazfpDb9GV9dB8mHcGrrmIYKPK5xBcOR+Pk7ep+FaTuq
tbgE4ruS40kbPP07UBgiowZtPj1VWAayhIuHFG6LCqP8JzUUq9jJ4zV5WU9S6yfh
klxADm0Tb8YK0WMiK9KN2eM2z8i+mzp9IbYDUig8z4cu0lcbDJqA3ZMlnZSZuqqv
DSEiAiMttQpHKL9+ycS1ihiuq10GzaOx5hJrz5j500u3YiEQVIAHuiptKfzBnOjr
7RfGMl5454w9DMPxl3TBk/T6C3XH40JenXeCGgxqVIxFAkKkLKy+TgUtAhFUiIpY
o1smOxWB3AoVxT9Tv8+h8PLhy2G1NdC+UDtaWFSwaVz/SHwNNPU9Oanz9CeFADJh
dpkpmBpku0WF4gm2w5SM1rNVJzq2vF0NM7eenwt0h5UWZ3aca5gJ3tE3/61HQppL
zMGuWjrPUsOdpAviNsOmn9YbrroCv1lnUTvuwQXE2tsQgYD4hQKdePqK7fgAeVCn
wf0Na9BR6876tMwg8ThYqfLUjHL3uFk07OWLpCf3im5DW5dKFILwCet2aRHmyP65
PQP+Nf/Pv2mOqsDua3FbtplQfh1DImrZTEj7nYbVax2EeFz+iu9KMgyNauqmxE/v
oJf92A21LvDTxvtiKcLfXLAher5ci5Bl8JF3ImuhyNTZTo7t5j9ym9a/Cm4+wmaU
TaUyJ20Quv9BidV6pObtLO0hVqatNjPJrFk5MiKD3TbX5JN0AlTjOnV86K5Ns4FH
C46dHdrfBVkgnksFCY+IiWom4zTxDVTMcZz5hLV9C/WLO5KbOiJxQKSfvqxG50VE
8T2mHDqfy6jyTpM9md4OkLz9sLa5qwUfnl2AaT1UMQlW9q26nf+iQ0UkezKqfeR0
p1ZZoSTiLtyupTaH/E63G15Dh5LynDIYZs8n0RWA5fc0xARb5cOLJcxh9N/pRXSf
+PYUETYaOnFTFJ/LkaWQHews8kLYuJshj3OYafjvSOJwL7yFyhz+zk6FwPj0X+un
pMMjifuppwZLIP0+q6F1x52sZXoHFvijST4ff7zeeYoU0gglzswNJPzNRD4Xl1BO
RA3Ddpe2Zq0xWzbyTQ+iT+TWMWoyfQ8gqRG4mN244jiiNJPgaFVneWCqrqT/a24o
1OAUjUPEXsQmuBIm97HdcIeTRTP7zSEAquO5QPpYHXPc5P66lNokYdKdWJ6PC5gw
KQXVY0goAyJtMVlnXe/z4bBqwtEpliG3Hh59m5RpB1MRHxaYVwkUjfuSbuVsrzwD
Kd5Q+6kxrs2e1oj/h9DfN+pOfpzGYh9pHxvVEPQziLQm2jlZh+wzYbT1kCw+u8b1
vqmPZpZxGo/m1TvKwFzotUij0slg4uouUqHS8ISJW7jGVkZ4JeP/18y/8/8jWKj5
eulo8xH756o8BaNTKvPqPuA0Ax7JzbleNZokZ0d3mJ4xKiasZOl6U/Jg+JIBei11
D1W+R1aCNPorELGjLqox6C51TARMmZoQsMkATOvRshhsZGrU8etIj1/5cIioAG8E
rcJLc7Zuk03TPASAgH5KnwmuDLgWt5pS6qo6829/SdpjWTdBS2JYCFGvjPHSiNhN
EgqisD2SkAch1NZ1A4CzWSHLL7Br1i51CAqbC+KEck1YQHk2rSDeNoJyVEmeR2SW
WdGQyTv+R//Rp9WGDPHVBYfk30YbVPEjLFr0pcXPpkDfaBo8UD+QnFVxi/4e3PGa
UUlMBFPa89xyeWDUj3FcnQR1UyasBcXKBy4GrI3WbThk7GMUhiEWmq1zc5KkWZwx
z+ldbLVXxEuUSjjqAVP4l39UPDlBz01SOw0kjYMZQeepMdiaqNk+Cjt+ZADvGDJ/
2zshg8zRSUqTety4sup7OM+ktOtK/lb0xU954bUCwOA6C0U3kpkiEeUevLTo9n1e
JuHuQdZwAdu6jIEknb8tklFC/NeLib5kjNXT0VDAfOmROILN4xJHfrtlCAzykTNn
WlouV4tDPw65kgWSKyGTq54+OnyFqGGu6MQdpEMexj9kAeW0cNG/qR2A+1UinDsm
6deIfl9zbooNIAws8F2VopkgNl4f6LF9j8vASOCSji4+nCaeFxAT0QqsjBAjOPvn
2hd1ZDHgBzVAmbM6ENuNzVkq7Wbgl30gPSXIOUXmqv5DNNufr/ha/7GdqZIEBkaH
7lzoefTfgB4R5cFt2Ktbh96fv2YwxeCKvTKfpzjLuiX21xO52P5Jhv69SzIp45GD
7ilUXzMvXv5D4cNqD/cB+QXRSisX59y8wDuZwSl9A78dpAMa1GjuFskGonvOnYx2
tmRJ02afPGq6z8FwHSUf7CP8zZJJ1RybE5AeplvqtlR5DRTr+tJSa4MX8WISIgVT
finGjRDd3X206lFW59YZx1yNVuHjpP+0MH2lP9K7nctJaI0GA4s5isuWy9tQPGbg
ozbD53EtrACdM9jCRWtwYw7Gp3cQn5WeSHnQFjJwW4gJ0fy+c3d01SYv+adifvYm
QTNoYr88XKs3XF+njupOpgbZ+3G92WidNENmXhZDlmpoL99tJtgj6kUZCwrfs+K8
YTGeTMQOsRXEbHQTiO3hhwCPNQZ/Ee+YiF53qD6EZCJr/oBN2XbWl4zlUcVg3Ynf
BaP3BDO1P4zJklk6V1edzoc+3jKf/PYd0p4yN+ohzj8uhy2pVhahBvB7VvEnmnI6
Tn9WrwXNa9VhKB/YaE62K+uSLz73NGYYCjxiwk9fKMozcZpiOiccbBGAC7nfjVUA
M5i0QhXRRbuBs4tc9d/Gz66fpX8IxWSVegTg1LzAP3Am4ID/xGMSpFD0qo1vdkTu
o5nl6UJnuNBDSg8rIEqaRA==
`protect END_PROTECTED
