`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LygmobPRXODVFBT8cB4lZj90DewPDa/cf1ZKXHPmDgovqY2P0g2XJFNNb0h5KQQX
d1hXFnUynoThqTVyPrJfUWziK+I7q/mss2LAKI9qNSelm6xRmIIPDQuPdmbtkEUu
BHfU20OShXg3ev/5MO4yJgHHIakciMMP4PJBMI/eUrJhF8zIDSCvPvxbzkVC0OQw
xjZgRijcHacvbskq5zh/Btb+x54t9cPCHR252q+hvr89c1QStX5a7M73CZ8ZaSNr
z8NQgE/ty4TH/wy1N3qXmdRPIqyO9U+DbLn55uVHDE0tmdFiTFCyorIdNXZMJtpY
XVo5YCs7zVr82pQhjlnXBn1Tn9LmY/uohjmMzIew/Slo3aPTql98Q2gwAt65H1lU
1m5FG2SnxZ4hEGQF47iRmEF4b5Hatdnc7wRx2yCF67wq6cJg2Xc1M+bmrQzFH0Y2
nvyizrAhRiEj5a+ylHe4OUwFkBDr0V64R7WGdL6ByoX/rC6/klCDLH48ntLqALlV
rsSAdowHbBn3DZm/6oH4vmIWwopHAgHeQanbW5a93IvRzFFgkBWFFOO3gI2wRuEa
j5+wB70LCIAeNNQORsgtrXAKXipaafCGXDlJSKAzWvsCczlxcy538+uxWeJzqfML
WOLGS/rSsy41y+ZrHm2K/7m2CHFSVmL4BNTqGF1YpHfPZLt2ACdzRB0jtQkhzE/4
pybxCmDipPcUIDsaeQFxC+qp0R1Bilyr8x0RfidBZYomJJYUSDSvlaPqQ3yBSeB4
oudjYnksxi2bUgiWkytQbl+EVkOA4MoFg1OkjKTHdbpNaqAi87nlziNlM3fVbMJU
hgiz07pal4oQO128wTxWnHsmPz/V3aX5hJIQm+bog9PmLpPqyY8KU6D3DYd5Q31x
EyLPMqOsBKi2KmcLm65fWA/SR1wrLl/EP50G/RCwzIKyzjvKsjUGmdIHAXnOrtoI
FnrlbhLYZFahLLRgt32KL7aa/bZRtI/BYLDxRcnKKakgaT/o3toJIjmdVrp3hRJC
l8WYSvZRKPuCLV25i9WNx8eXGf6TRePDcnMmmawywK4j74vxLiyJk0vXrpsOUOBB
JbmMZ0P+5rIJAqfuDQOd4jql/PXw9dIDDomzll66DQpljkRz2JAyJFShf3mv5ZUS
BnFP7y7qnNokNuNM1zd8RILNLKNeIHsGY854/qqR9IMoHJymwpzKLc2ASXHGAlom
lZsEIdy+vnNQHR0+w0vo046YNUjNfifHtFOrL62jbzbNit+veQQjzrA3VLx4hmwS
MZedrc3seHxBRMC1tMMbHfegsUCAh8ivZUj/qvl4bVrVQTBPZOTPPVdLKoZODbkI
EMGJjw/nK044Z53uMu3LfP9rL7wzIyxh1LA4GlVNELVrxSqu60BIGEE0aKLd1usM
faBmZBshaZHZAizH7Vgc7Uh+FuGMrclPl/zTRTeJVQVJUrOqhpORT225WDu2pkln
a8Q/uq7iZIq6UBGvyVVsiUQPPnkztxW3EhR0bfWCei+JgOiCAEtnSUMu+hkRu0Fo
BBqZ+f62UtuHzRv2tG5VMzGQWw3JG3GtYUP9B7oLxqQpGSdMrp7D6eoXjmiSd6ej
/jJVGdB6RaLjU5ix6vorhOowhwa8MMa1VI1MkLzMIxpFnIbJF1cdsl+56eEs4sbd
WPOgEi7rwK3KUWADfk9DY/qT3NpBPnah87m29oQSJcQz/2i12REvmNLGZV0SRSfI
9fkwazFq+TckoGKQCu+bUOnOeBRkaGcJEP/Cd3hdpp9PPHbZlzthJibqXpteFSZG
6CxUvC5rSWUuUfjHG0OG9iGsaBQUBJa1Kyv1EYuNeH4GHs2Hy2bTUIGZw6vl1f7A
HeD/ej/paPsAxR7Es6ce9w6T9hGCrGL6Jea8JAjr27nnaCXT+UURAS6dwSbpzEHa
DdWevrNquouojZl7eF5J/tqJEU5Hk1PTXCiKImPjTWKkUqPChWuv6waEJhIrrxFE
GUPp02e0miXZ6PzWaxI7tIADNcJBabK90YcOnSu1MiTXc1VCk+TiwakRQSulcBfY
hWV/f8rxYdOCIyn6fiwVnlNw+vCrIOdLFx8EjgxHmS8Cm7hdPbFRc3ltomDrghYl
weJGDrLiFWymDV98LI4mcHKNnrfotmL/SXoiIFQZDWPUdKIoOmeHG/8mkHyqY3Xn
+v95hCrsm2OS8E/KPNHDMnhyfb3DC+Fblxg2ZXhuOTAhYTS+RK0hfYKYe/t2v+qm
+0CwvdFTc89sci+GvfxoOWgw3TTKgccZqMT7cwXfH0PDCBTr8LDfPMq/8qCjEPhQ
rb3sSQlJ9aBeoWhfiCtqkJKl2K0XlYyeWN3A7+wYG7vaWahgNsmUCEqu12vFLxgv
7/Pgpk3Kt7r/1S1tiQMHBwHKfV80xrm3MgpDW0YzlR3JomUdUADDdybmJy3nhH1C
bs5P3r6Xqs8JxJDyc0FinErjNnrbBQSIBZUDJF1S2Z1BqNUHMuNpuCvnNDouLCMN
Dcw7hFRM0X6ukJ1U+bY8fkT63z37g8n2I/X5VLlgcXwW4DXIah1DlReZRjuZsB94
sEui77vjDcgAVe+A/STNX55/RjkAFkYmSSnMY8kqoW1e3VGxF4X9437CodvQkRoE
TflVuRttTtMYJ/FBBCHYTLxqSJac4y8z3oreB4dAgvo=
`protect END_PROTECTED
