`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jgxNWzKODN3qupwGFxcwwG2i7BlFkpAjJRkrrWhzKWEv83NA6Qsm76Bo2/PY6Ve
lwUSfm2VwCyIRWfK//RRW5iTnjYz9RoDATyBoXVWWHKGt3pjoBv6pX6ZsVhvIfnG
qIUzNZeImvUU9IijaVV+W/AF0virCIY8z4SHPUee43RCji34fTUCqtUFvu0f3um1
SdjLT+isgehSeEdZji+Q7i/I+VhM6+5vFE9c9Ns69RUc3eqPhaK6syRTVBbMNmPY
NIh5iRpayy4cIwlG4kx8zuBhcVYD/U57Ml5qG5uRQGyUWJtktX5htCIbjuggBWEM
9Jp57AlTDmXKFAJnzh4+3gbZRQfrp1Qq0qWImlx9x7KDzx3iyzEfEHjXgFoefnG0
bIMkaEY+aiVJb6bnc3dtRQ==
`protect END_PROTECTED
