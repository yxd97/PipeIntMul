`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OpHYNWOa6klHBM8CVrLtQpuvK45DK3WOaCsWbI0fQMnX37lVJkh5VWVjj9fawulx
uZR+cso+cKoVk8qgxpTk5Ybu2MivYJiW2vfvyoqIzTJh/v8dvgasdHr520QKuBos
3nAqbLTV1WXfJtKqIuJrxuEPyyTq/SO5FNk2HVtkhr2J+uF0BjvOMEGGGLZvzYP4
CJ+uzg5zBZqQO07zV6UprqpLArltkZDZzkh+APtcbgO221Xlw13ca6X8rrNo0YXF
OJqWLMT3oPqv4WG+5OjdcvIoSsD/pWKU0jfEJt5/dbB/QgMhiqfSSJTDLSpQs7/T
RbqsDKavvjxVzVguIEKcr1Lr9xa38h9OTC3G+3n16VzuRgezUlRklH9w0xKraXZS
nbi1AlIxMYPJZg5RNq86vWXnE/bVKGJFl4sQrrcmlWLPOefvCsutIr6p7lYWO4cS
F1ySeoTu1c5gGjgJUseItcyN6WufGhRn+5uC8UjjW4okS96dLC5xI2Qiq1/3F0tB
WV5Vw3zmO1LHlQFy6qMcgv0PLp6hm1O6daYmu09iOVIOsdRnd7vtrYUSmBzFF+Sv
Vs1CFmbcfuHED269Rj6mfA==
`protect END_PROTECTED
