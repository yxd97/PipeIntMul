`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSXjopmPzQ7fAsecrzhXoAYfa7Y2+NvHkS83+LMCWlAL628C6qE38CCJYhHZBEPn
l7x6Z5sU9nEHttOC5czu0qb9CwC8GBhyz1qz7jObGG20th2+y5WG12gM9GYH+Dv7
nGDg37g4sgojnFy2vQH026rBDB3/mVbR3CukfiowjsgA8bRtqggTxgvchh7JiOOE
fRWntkmvn0XNXWJ+Z4m7N9VsJPj5om5GyQ+k4ZGT2HpqABnefGO8zlZRqoCwq+tz
kHpPO2569ut3rVWe4vPdxzY0gwR6VKZ4VYT3InhtqMmnvqOJ/btXGPMny3QemIjQ
1U4W9ucsiCNy7/gou3MHeFAa4IMkWhxd5UIx3BuiecSFVroq1jhEuROjQ7Kg42OB
mZKxNm14NDNVY6lUxoHEg4vqU5VkweGeJs2wNPD4vuhVpPk+a4nRHC3n8qFKsQ0o
gvEiRYGlZ4dtg7WKVIXW6iYyPfHp4IB2JcMWzxgMkxUsa2PrW06IQBO5vxYDQubp
qvOMW+hJLyYV3w3LE6jYZQPsWonIzkng8Mijj/Jr8TeYN7OeCBBSupSUZ5rdmgEP
YyXu0F6T4iXxiiN6j9enWOhz6u7FSGY4cotrKSmE2TcvARy/Htr2iyXZ0vbN7sE8
A9KMTaNP6sd0IqGx6S6aCA==
`protect END_PROTECTED
