`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZpFN0/FwILHPCRIXm/v6keU6CR+MrawSHzLn+WUuazAqxLgtnUxbygU1aa/9rkLa
okx+d4ha1t6fo8v9rVRcPOHTSQD9wax69btiIINzerOwqd4VNROZo3gHDBmr+Ke0
gX7l9AU9f40gockAi+BVpTrGrf1TVr4UifRpEmDX3QIH09dwOZzON4875cBzVA25
WuYT+Rgj+E02U+DVWWlDe+7qph7+vmbv06iyf0gkQQxuVFz2oLMQoYi9SmlztHYH
rGoIwy+Lm+KjPuG0YNMFSixix1hZ3dw36edaKfDSl9lNhErrrVJNIVdORQw92DIQ
960n+mNrDBfkcxK+VMikB2lF4hP1Meq7cr74Vj/Esll9Bq5NVAaufdguv8aS6+zo
rLMP42j+ByPqQapXqcBthw==
`protect END_PROTECTED
