`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNYc0fzyu4FIe+Cz+w34EAIdQaBm+aA3GjKxNH4IFxA2eLGwrktkaCe0AhELrABy
Yig9cCu1wvOorH3XYpCnRSW/Iggkwh3HsE9RhYZuJGDcP+KzxYMA5RuxkXaa166J
PtERnThuMnGZtRuRY5TUhxQ6IEqGEDUE9yM3F4wxfMD1fM6PGMw/x4O3xGo1oK/N
lnA61gbw5UUYEKtgCVo3pKxd+cSc0pA7jwpbSdfkjrYbt+x0n8dmymGEYGZrJ8s6
9ZP7EO2mkGZ9L+/E61dV8Q/YuxVKyd6xfapv9BC1Dj4ed0xM84iwtpoxlN+5wMKI
eSCtckgGyDsyUXEEg1FoUl0q5+nlMQ7llBVyvmfVLEIitAX5wKYsMK09prESVbuJ
v/JN/ofV42JLHTk8Yz0Da0aoozCjsWdpvYtM+4mHu9E=
`protect END_PROTECTED
