`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O00bJSJG18WjiGk4tmKYyl+nX2waAsF6X2ct2aJfxTJyLOiktqNIHuROq3DEo+z3
v/QuEHo08SPnToST1eHdrfhLNShxEfrpJ1QlMgqE0yinpUrKcDJn6uf3M/2GxSVV
OsR7BJU38YqO7k372QsSbCkz2TCBqKuEqEpKdyO/ljrV7egyQqugawxOoSMAmCjL
mzjV6qsKNEwArGhsaApCpPWOiqJzbKG0oPrmN+sMKwtvOAW/YSVE9YFmmHZb8NLA
y2DDNEw9NbkFuxVz00jD3Q==
`protect END_PROTECTED
