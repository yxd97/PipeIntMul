`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jNSCEWA05YlcmckPjKMWeroBz4F0U5fX3DNQ0xjayCyYNP+/xReGX0Q2P3AoHFR0
p1MBliXBwuWMaDRTvZMnYdpcKIaVml4fc2Knt7xYa0kCXw8CrTALQpvwLqTeZrib
caQ3k95rXi4H87XAPFazuquexkR7d5jR6pOdkGenICEPIJxo2AiCFmbTM0hEURfB
CbC2h1ddo3IW6+hAEzIupygTPle2+WzojlYHfnqa1bYqGOxAeA19IQiK7mi5dIIv
7hizPScBsp/4nYhvLYXK1Lb+54aPXs/RtKOvBGf4s3/rfqzWf/J9uwu8heRL2fin
fq75/OByt7bJy0oXC+6fLggwAYmnrmbwUujG+lEgRdhSAHGdUZ+Tr7eNphRhK0jg
qBU4qJF924BKNCYWS8aTMLFDsK5qLD2OQc+PijZmejSdxdxMEBb/8kjAVvHm7aQw
JPfjQcfVJ6ZQHwFptlKr0YmTlNb6PGlCTNFKE1HmghgMW/ux3jlipiHLjFqepIr8
cuzoRq7ddn4TfBRzLhyDVI6dx57hYDxq5Zeon65Y4y/BXa82PI9tvsyqhyI1kl8T
smXqSeQMzK3kPk4SaYSHzKhASbgJwg8I/fW/VQmzxYMOR7jTZpc937sc9CpVj8ao
FJGAgpg6mb/NL2uvICGGkWsnpGd5aZa4cJhsGAwbyHZX9uiXITn0Av+jH6HFTf12
psyxj5TTNv6KBGoxLCkzJGuF1Cji3CjqiBfDK0FxvMUeVgH91Mx4A21Jx1i7zbOt
nLT0OT4QOBnHRSYBo6+W7yClBnTEO5shY2n5MKdqfBx2wJJ8knEGwKIiKoIsjz50
y3M3RYwFJM5I1GuywW3CbggWuOWab16aVueUxvmz+EsX8K3/ZVV6BwnBurRRof5C
D1++/nwFySBEiiuvB7fdiZkLF1O2k3noSMYhwF370sB3EJzaGzQgAk9/M2TiZ4Gv
tDU4wO4j0HgnhHPCUFKq8xQfUEnmAWa8aUy+KumkU17NkUyJABPBJrIXR0SrN+EF
hI/0VEZlLDxCEv/rYhBkT5oPEuJMTm6H60PCif9Uar5qRmKX4azdR5SniUFLVU2K
Mtdy4F7KyM1FnBdYepvz9FNYwZMJOKfweC8q1YzLFQbyLDXsTE5x+n9Sdi6gP5KV
A2cpiHawLmF7sxkZx5hICgVvK7qnuxlf8zAMKb+gOPVEsEbFwmZpW1UCxPrR/i3T
yBf0rvIy5r8OzwBhI19IdLbGF0pU8m7NbIwRnowwrBQ837d9+3yc3GqJEDlz58kd
`protect END_PROTECTED
