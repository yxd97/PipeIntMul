`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uW5x3dWKUkdrpFAMo3dYdh2ucJKcJJviDytye7vcY18f9YyZyQYvQX8YGpu2j0Ui
cy/9xfA46sDmxBYC+9S4Vw79pw99KxcBtnxNBUSJDn/ehxujZ//50YorMAjvXErG
KLnGnBTv9v3ITKxZ/7mOmNUCZqD4VInm87JFoY/ad9nsD42uffyXhTSAaBAzVE6u
mCrwrzbkqpfskexiFnFFabBF3nKZvjAk95m59+sDof5BWcoVNGWeWfls+bDwpF+1
nulyz2ixP7WIcqcp0IXbz8X2lL2fohSuULqKoX31+Ws=
`protect END_PROTECTED
