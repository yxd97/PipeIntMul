`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAM4h4nZxWfFXTBvZ2Yas+ovL3zwDSELgxcK4TAjE5UVWWGsNEC/u0xaJQ+zISSC
mdKpQv/M2LppMjB7a1iF0pfM49s/FWusLMhlKwPuGcy1MDqmmlN6oxdzpVNrpMt0
2hrIDZMIjwoMwro+XIqXFRbVcnwbO4arkO24x+cYxFoN1Rg/QLTwbfDEzaNUdmRs
dszJqNonWSpbK824KIScYUj6r8awCcUujakBvnuVWLBNVqCSRtKkUidAVfSrs/Ea
Gg+V5aiA2oDvuLPWiQcAr3cCXOnxh8HIPySz7LLeCuLnbzjENy67fawPY27vnGp3
vyxjMbETXnclP0ZWwCo8oASZJAJiOf8OcEtRIEE38MjFXGRa8hLfGkze3cLMt4/E
Q3uUHgjHOEwm29A6vsPEuczm/ZauetOF/mF5EeVRIziaFSUkwoUP17YMT5pu+0i8
2d/ynY6K9pIj93gUHwgcBL4Za2h5r0/EkBgJ0e8E3pSvdWCWYAnZ+3z8blB072fL
bbarAegIbE13ABVRPcIfAk4oICLsBRccAzgMixxGxil63agvm1pWWv5iQRsjP/Bv
Db1VYJQxPqPCffZsJM3n9iZT5fSFDNTgE+mvb/K3jnacZ0vJQTS/Waj2jRAUzeFM
V079F0mDgdPdiwxO338Te9ZPyVYruJNQ01yZ5ScIUhDeAYOn45HEZPFytOPGgDWG
010htT2xjBgR96rHCx7D9tmOJCOczCjVYdC1PO6uAOARReQZ726v44TA2PDv9/uP
ydeHzP81pnyHIEBi3bkoP03rHRznYbxLJy1qNrdFPItORXRiWgS+huPMjq2vAH4d
UYOFR15ZqXJaqw84cG+uy0Rc9lCmsDv/+Ds++jm98w+e6UuKCjUahx3c30PVTZ75
h7Dn7jjipRz6GqmFbmSM+GOnjIlLdfqxL1oTBgmW26u42Xv5cHBsqYOIZ8avw+Qx
1YMtXdzlEuFcFLJFmMhkxOTx+dYEiUJUwomVbcLNup5dWKQCpmNuDfpEUhwcT5ca
bkZgNapTKn1aR3gA/ZN5c1SuGZSyhng0JEdJGr1zK57FpGEPUQIasjoDo4Z3D9gg
oZy1L1Fm1F4Oun4B0wNeRW5bg/qvjqPyH+NUZPYJfiQJq6dQEN6RFq6h7BRrEu9J
kzpf5fNCBWCIvnDaxp58s41ugjA6tlAu+qupNYpQj+/V7si04RdT0z1suI7JGvsu
Na6bUbaW50iMRVoMHw62jcT+KDpirfGjM41ev00f/NDPZ5/dGWNKCPxUxy0NY5Uo
MTgj9u57IC3OkdeWIjLFiFGVY0z5Ap1Qj5vqrpgllh/ASDYsiVxD5EouJHuDjb0F
HMENsEpZpcM0GaQkv9miyUA0Lgira70F0hAzEnRvh1BQ5SKpwby+zBVShMxzhkxG
OVKwbUSrLkVok/IDU2Fp9BjJhzrTnX5jxv9RvB2iczvR+Yef/PacRkQys44GQOAC
RAynWbZXoU7T2Lv6l9wl1FWAWYBl7hU0WrUzBgXMQGALZFINlfVEq5sCnHULqO7E
nFk9RKv8xepOvF/Juy8h8abOt7BYtut5UzeLHdnngzeJtBA4tWAMMzS3zzAkf3Ao
eK5e0vvEDSe9tC33JcT9H3DMtpiKaNqFa84vSCdTfYilJ0q/H64EueD+SuiELR5D
QcersUpfIAuneagZpdnYE/mpPf6tQa23iVkP/o6wlsEgPOEa9rAa8aSV6cdQdjPC
kB0132Ds4VT1C9GHyOJSkm0IjmEyfY58RZIC4lnhKX4odDTrqekRKGTM1cf0zUbv
29opM+zuyJgZFGTzUTH/G7l4LuTvHaKja8xyoNoXDTwns/F/6/x8ujIegXoYc/7D
LWNUoeHYhRQYzg/2HF2S/XD/ImTuOO7FA0mSSMn+Mvw+5oGlHwbtyC7xKsRKcDJO
SZxCycRgQG0DJ2Nf6va9UA==
`protect END_PROTECTED
