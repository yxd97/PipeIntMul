`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Id3D2L8DPOupCA3D39QotuoTVmIXR6VntGsGfpvGnwh+KZW3o3aOPziyC1rdWX+
dhSDoe0+t6FEj3smZ3fPvK27yaBsCcXDn3HLpSJar8q+L34B2vyA8zNj2uCXSxVd
BSLUkhMk15xkbFXyfTRdvExjDC1iU99M0ZCiXY8EP5Ln6oYKJgkV+dOr8qofa9WK
GBlEmzKLc1C810u6CGsFow0fwQTsNFKlaiHkHvWucLwJ8L/nsJ5t58zoerWvS+eW
ZXMGOKHGvm4WLh124Ic2yi480QLmVKEJF7c1WDYy9SI=
`protect END_PROTECTED
