`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrC2P0/xW8rEkTxstqNpsdfOZrYiGeLLYKnitxZ6daXWRWwT3e2MzIIp7XHdeaN+
cCJKHV5Biwvn4uVSlkZIVCsMuzm43qX1rFN3T+iRP1YLX2bablpwKIYaCsLLdI+1
G0hBY5YQwi4W03dCOYVSfHGEbu5ky/HSTAk6/yyiz9HAbR1o1LqhdEv+XFohbbl0
F7wz33yJj6ezCquMbwEcX27VpuQYyUvwYb+ONIil6AWGqVgGM2lHnI4nV6mIIwIk
a+lpx07EcjIb9aVTQV8iST5JTfzA9m3RA8Y/Sf3Qz4Wpd8Eqqr1Np8hGHWfuLBD7
q0Sc2hoeZRzcMB+LXzrD8TdzLESeLRk2HvH72vAy4GfPBiJUHJXxpJ5XQQi8oRTZ
s9iyd0V2cwwqsWmGFE/kpzD+mUWW+nr3tKOpdm22pBU=
`protect END_PROTECTED
