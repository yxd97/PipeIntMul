`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZeu+7WoJZDVucnImZmYTCT4WO88Ks1tQL8/JvoMLTgp5ezEv1ci9GzKbi7iBt7d
uonhybqQiLnHQiepEVsX4loMaoqHxlgPvcnOp12I/Kfn2Etf9WE+VEeBXqZnOExe
fudmOdN6Wy3wmr+MErf/aYAV7zextI9d85s9XDIsgEQGEASFnrDSZ7y1GYIdq7dI
F4ai52RN9zDX7YUxx+JC1ZitmCjODo2kCOFywnkTiPgeJNKwT8m8Xmljd/BnLDaq
uB2OGi2Ue0aFwst2ByBvR9ItB7pbJNM1Q9g6130GnTpTFM7di5rUkiKluMzSs2Uy
3feZl3w8V0to5mHsVPsSdzPFq9YQNKkrtPKFjBbOjNSi5qQ+cRaNDSTu/mbYIULJ
I2aiiB1XLXERhxvgTqq/EnRxjA3ZkhheAj6ocseOXPwRitvY/mxy7wRRlg27Y24y
+ZzvUOaD1zDinLYVBBDGEA==
`protect END_PROTECTED
