`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5JHKdkgJW5skGeZuCfACNJRMUcTjmG7PRVOsIvqu2ao4yFthefqtzgXqEk7+hF3
SEpDZ/8lHFeDHfoerOr61Gbd6xTO4dAq1oI2aVfunfVRWi+Gnf79u5pjdlWMbqQ8
iFDkGfW2JniG80yald1Io9QP63DGOdeENDmS6vVmdErCfELr8G2EbbQTQ68UcO8w
L6GQml8SRqsUGkmJbQRLxN4IyLCBAWssmkNOroFLVLPFtCxVKxlXNgDO9qKnrAio
qk763h0K71w0BLBsDxVc9Yp+hhQuq9REi55x5Y7Hn+adF85Usf/MFtR5Y5FXtufo
t5prCZPh6ghnGjgM91olHpy7duE7eTYFnxy8o0AtAVrh0Ztq8s7v8k12jgDUPdKR
54ecbAqCsLBQqXufAeHE5q1CsKCHcEPbvs74SM4wyz+MYt8JoydjK+KhHtNanWNW
m/1YG5arBJcp4YrQejhLyLMCtQUc8HRK0DtAyNYHxQoEz6pLB2+CeHiX9gxnhKvP
QSC8hMUSYzwDLSwKO+qlsNwg62M011VtJVu7c+9WusHFYKurNjNrGV+++kUyy5bB
9iGJmtCeux6URKx5zKerkVkTiatYsWuEmivA9jEyyY72KBtpTZCL5o+k7jbGUF4C
wnfMEdhytvDvemMrnhCv42ucZQhU6RRlxzWSz4ySun9Ml6ntFHjliIs011+Z3CAC
iWB5DRKqm5cJWpuhH+1Gkhn/TV3teHakndCljWd/Iion2OubUokgNQCeNH3zOBzB
d4Z0f+ZEIzKQSH+A/ZnvteFBdX7hLZXKqNuHdkUHbUnhvI55LP+MLmUxlQb4Hz0j
qh7LTYS6nidPzp8tAzMSkuRZz0RbNGIqe6zU8yuSbTXJVeTaIPY28j8FuaENH3yF
SfCd8J3sgMjtLj6dNaLXKGhmaWs3HnVoaEHWLtf3M6M=
`protect END_PROTECTED
