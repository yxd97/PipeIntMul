`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zE5zRJHa6hxnAf7w1TK6S8i9vhr5YFc+R9DTnq8PM3E10jn6oes5Xz/xEnfAi+Mb
cp9PjPiiBq0aGsTjT6+FH4YzkLOOSeXQqNdwCOgc8Z1ftT0G4DuvQYYgUe1dDDzZ
2FF+Ih7cMeqLIrNSoEjRPjv7MNUV68lNCzduFFzcxGv+cqcJBovBSLESBXhr2P5u
0bHJQ967rfnOme2zXkFgoZGMwHhIjsW2Ezje80TXCH185mnvDmGg3WRkiHxe8nn4
a53H7CxIAomsFYuwIdtZoJaDkwXZ6OI+RPTnsKBRXZSs8IZTdWKCO3SXiFxD4nwK
/NF/vPgM7KLaNPEyHr+7J4sx7aLeQMzTF+Q9+6X4ZMFLtnit+05JAWl0MRNj5DWc
CT1JnMeKb+sYXkaRPBCZ5acOAcJBwQ4AfyAcVh/NbmFSnKbMwgt23rNhf/m+qa2S
SPzIWJlL70zc1lhpMIDgwXl5qPDVnsanlQY7olTyNJTVFazCckLp8npuszc7XKlr
`protect END_PROTECTED
