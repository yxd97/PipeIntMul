`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJdQK05HTCbX5SJja9XmWPGwslH/AlsxusCPiTqHHrrEUJw/LpdK7/3O5XzO9wK7
Q4DjEdIrsTZwci/LlexGNdnpXgjMQYROrB0u2QJ/Nu/R/pybzIHoh/2NjIHJyEzn
dgAMKea2IgTjGdwyN3JKj//pUTDAIfsJYvfgC9TkX7jygV/CJXrFDqVxR8NkAqsj
Ho3cHZFXk44QAOTNmUuJonff7RqO5CTYZMSo6hjw6PfhQwnMaDClySrfk1buwqTN
He96w3BUB2OoS1yFLg6hlDpF72H6ivJwvVHJFfhipCcfrjBTmF01s4PHxKiPmekT
`protect END_PROTECTED
