`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EcgCtYh8OdW0ARQqpSlp98I+SIFwkaSCDOb7a1yr6CN31e/ad8OpynuWcVoncsL
zs7zzeARajx7q7PfCi7AAKj05O0ZjRoQNAu6c/uHjvMCOi+nmzzhOv3SxgZ8fV9Y
7lSAkbQ5inF95kj6q6GdYuGFFNgvxpHX/+dduq75g9bIl8PvwabxM/42+VrhxvnN
jxkTij7e9lMFlY0CANOU1C327gBYvjY9anPeoCQp8fuYLi5x+N5p6pllpIPU3YaP
xIbqoeoxgV1NXYXE35ALbaCL5quF+3ldmPmCmoWBLtupLTG77H8xT9NT+26qdztL
4dV7gQV2sBNQ9pmXnwPg3g==
`protect END_PROTECTED
