`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufsmoUBGXdqU14W69MMss91FiugDhkLHRWfRJMzqgPgecqmIlAQkeyQcFpJmjiq4
vJCarjvnBcAUKRIdMjh7pzRCBZzDd8/a1/DcTajt15gIHzDzVc/n58Qn0AJooIfb
cSXnNrlZhnajqYcDNVLiZLom1BaC+FU35IW0vGhDnAX+VPseC3K16Lwbe2hTfkAn
Ed12JFTVN5+08hn8MtgtHkVElZqMB4QHod/VfkXwaWrSJ3pRElb4HMrZi6dWfj+M
qAQEJCiioGUb2NCO5uIg4LqRhdmg5g02e1x89oPrUiS86g+rLP9Q03ndVHvpFBKQ
RSpxqaag8HJBQ2zTpZIArlDAadziezVkGcdKXW/p8krUZwLm3FOd9AvQkNz5pB3D
fWUNIsgiZWowhQyZ9Nm3AtY86OaIDIq0W3cq7lZ0nhlLcWSiwefRIsqnKKxpKIsn
y3PbOOt5pdRoJyw1VSO/Fk6pLHKVjdQTGzZ5ytgxEgnnLOKdy/wvZgSUWN5A1+To
rsP86c2ajy3VGd2E53aiXwF9g6CaSAAkwgdO0s/FppOLoFB43OFrZDeXue17Fplj
lxm6ADsMlRPAxABvqcWuTLYWaWgPDS1ZuPZRn10feLTCSVn9wpVklFE/IeWxgIGr
0tNRPtK51ClPk53j73a6V/yRrNzb7pNGpg3SDDYCLDPs3IxcQuWWcci9/paIPIc9
ikOa70EQwly0lkmHqt/OujrNEZm+NVQwKXD7BX1LIfawSGyV6wVpZJI0zXNj3zzc
0VDfsUmxDv/JRVwx9DkEaWI4qb5LNLtX3d7stkgjN53CFHbMwMAlQ6VouvSi/ge+
/vX8zx7X1WVnc1NetGA3C9HKy3Q9CKAnr5zUh1XV5VKu0CpiKc+RhpWtb8VnctjT
87PMauvo2/HRn2OIXid6CI8G8nTMhZ+pYn9ngoD9AKchUzO5T7VacD+Yv6MLjMGN
+xwNZzEpxE4AEZmHJk8y6Ci0jeQjw5bWwkobb0oefSv15Ht/K2fna81YIKYcmBvT
5rWRRzzGZgdqvcvzIn1/lMAPMhVKrIZOtLCe6V3n3T6k4pNAAYXbSp311N3zv9JD
JqvxvTt4MLL+YKzLVxWiIMl1/wnPL5HQj8JslUqjO9eDMFQckVTT0hkp2AW0ARAk
WbBmqGSVXmyqQqxmD/bIWFNBBZKrKm6jKiiImqKaeqRG3+D3hHJUbu7kZ9H/nX5Q
NGG2+sIOPBBCdZA362bKVrR9NkyztjwBjhLrC8/7vVSdCJ50Y5McLdW/WpdkJYuq
EngXmTfOPeUmu/s1GPp1/KUYKZg6f2FR4GylgEJsc1+D+Jj7k34oGiTyhfI72fUS
D42GNt1vcTBd024JsoFs9bgagZrOWo2fQGPGBIxw1izxCHI4DGErK0kwblVj4moa
vqO6XXOALRz62kgBSY9jVurJT/D0ZkJG1VWpao5SGFLYo7hL8zgWFTQL1qCEj/Gb
LBe59WtRxlUO5uHclz8R0hyg5EIX87B/Mr9YcIV39igLbe5vZUYxJ8ZK5OIRkGF0
TlqnIvQgIYqhpmHsoWHTUfuADBDPa0kfwpNym9Wc8ZcF7VWFAwMkH/qUBZH7m/Ko
+lR2HAQ7SRiMFC3JxeytHm6c59MDzio9GXw/oANWaLWyrSVWsTYrAnS9JClTjfOQ
01gQvQy4lvfVJCWgWfYlcY+WM5Fbej/iWSwiJ3NLN5J3uUEHiPK4kr6epaNzIOIU
`protect END_PROTECTED
