`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPDtY1YJ3U8yYPqnmWa77+oXA/6+lBW4GlowqaOHmyEqP9qIJUypeiXfDonZLyFI
2Vn0/ilfILKoMj1oUue1/NZZYPI6IiUDpHucgJnw56eBxAIyjVOq9XY2MbrXNxyh
ZywDwfkvtmu4wqZlpms0dx2aiqOH4A9TR4eUukGj9q4D7WQAkXZzzPAFv1SbNkpw
prVjfARIRolu+c/yL5H5og1v49jEuTO/cyjdQBCgUf4cq+0ivGWrKe3yHmO/PY3s
veAG2JM1sz22P0GeFxFQVZ2ELE9F8anvi42f65y22YHY7SMGdQ/xcRf9YQNqos2G
Gp276M6M7UEu5npUzzKZT8cU/CLsupWRJORQPwT2FOJYMXX/R5B1KIJdfZQa49PC
yqltsrtoVcI54wo52apKuioqaSAhGtigqzfbCCGzV18=
`protect END_PROTECTED
