`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ovzmmzbLJ/jerMh/ol8GTZW5v0zUUJqV/PnG0ksJU29ukLHvmMGGd618vlGoHer
759MG+xVcABCSQVNw9Yxqe/0wQgUfTrrbG5t2JfQC62qBsDX+amBqLlRpmB/mpe5
gMl0sEEm/sUS8+GXpPReHz/5k73r874XVb59nqqrI1hNiY4uzpTAbek1yZxc30uh
5pZFQE3sIMcLenb0V0pU0BSkoVfvTgojh+RZvcKnAzPQYvy3wzNSIXiZ48cIbIdl
`protect END_PROTECTED
