`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QNZZQzoXViPvLyROml+6DwkJ1ut8QGms1BS8vvKTif/Z6ZIDLlOg4Wr7pQHldbo+
pEEYMZeVfCYcYEozf6ax0pVtAW6wWeupOIXXJVwjKMIMRAJLt390ZG1E3K7+c+j4
HgDJinxO+AJ4NVJ1GYBCYLt5ExaKysKTm4jOvr9RNHFRMi+YFL+nNNng0rKxkRH6
TKNaTQSbOysDQkmA3eYdCYqPTO21Y/R9evFJFOUsgSSRkRVc6RNM0QbOkqtL6/AT
dOViGskGDHHNoGSNyOFoOA==
`protect END_PROTECTED
