`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
007tlUpsrBUMvD0hCzETo88SHD4w2E+IbOvs25ylmBFErB0/MpRxE2MXFN5uEzzi
niLo4GICdALzhZQQeNRjr3M5Btc/rJOqHmvH8eweBfH8sIWjoXtmvYi2TD7pcluX
a5sDnheccn1xiQMaCgRyudJo/OKuGHcehF0/ys4KnKl75R7PQp/amti9TYtggzUv
UhR53tYPoRcBOylP77vtIc+pDYbf6oF1+3TiYRu0AT/2FNrMBwawcqRG7avSZt01
5iGSevzsY1o+qrOd40Iz5tvFuRtZjfh61XV5k8MimRZXLGlWvThf65YoS2KVyyu+
w784RHcDaxLVPZuptzcv9lNZRjYkmrNChBBtlwoZLgE/0UuHqOuC8F3OSUteXiXf
5t0gHJn3/2rGRWHPx21VVlFkzds2D+GuICvCh9U2GQd9wwlA1BjCxQiGo/sOUAZ8
`protect END_PROTECTED
