`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/fZ+mKOL1eNWwk/+0e+YwS+VNof4CTuVKmpcTStglJZUvrjqGCQHcq4d8l+KQZa
nwl2LEqw6jqUhKW00dO+j93qn/M8OUksIpD4CyIoyeXWGXwbVvjpPuJtIeSRDzi1
83NjUdgTgRjVrLoHQe9czoUchdK5a28JigDsPv2d3u6c1Kly/YpfGvXwFeOEMRkj
WK9hPUpQrrnoOV96jcnP1aJoBfH/a8zATGqLOpPxHwlTLcXsbmiNj1dBKHeMsIXg
pMCQfUiK2tG35yQTfBhmoUA8iqFuHa5wNJpicYcPXgw8LvZFCnenN/SOEz5Rw12x
aFHLxQrjRcU8WN8NUj+/kPqHiGh7mh941HsQjzcX7qORxIosBtm4S/KgbLpThZ6l
uVXjC/4dPY6UJEXjHacAOxlsrE69TiPlTg6y4C0s17SeM2V3ygxXmk+n8OJwU/Rl
HsgfhLuwDGRGVDwnZoPnRA0EyN/mmZlqFA4DVjclj/s8UtBqlr8UBTRUS50HioMF
HpDZ8CVraW7MIAEW9JS+/Ebf9ZDR4bYk/A6X/UyY+dI=
`protect END_PROTECTED
