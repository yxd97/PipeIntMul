`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBWRIggllyc0aarEx9R+RiDtRvrlzC2FMDdDgZHfNi+asDDLV1ImlrdJ6NoDDadr
tYNc85VUgeF9XbUoUN9oVmlPfmXnx+N+7CbWIVFkaqdE7RtqUaMv0hOHYIxFKEZc
SM+f5Or6nqYTTFkbbWpHQ5FMPYsHSkOto05ILh6vNJQ4NM/FwKRqq2y83occg8Er
L08LL58gJMw6diQy9bLtdsPQBggcd92lwWsIkqAZ4LAMuePq8bngDMoaV/nlD72b
HqRvDrYP9xI3Xv+rVJqeD6645Q6D6BXBVWoqbl3eG+A9JxqQTg+84Vsf6FZPiU07
S+H9u4QNrhyj3NdeO38PKNtZZ4YNDU6SW4Fy59Fqz2J6IwF+v93MxSr9dCVkcJCq
kiUvNdPw511DBKbvnsIgi+IgHguS0mk91W/QXlkr8MVCeCpoBqYPVm0NV3NnZ80W
/8H9yvtZk/s0TpOpnZviQ0R1yj+x7ZEhS/0DyMHLj/SOMVDstDdPWsqK/UtNSXiU
1beFwjCzjJnUOoYuDLwMTpNWRrBcv4lLio2HlMDnuAIoG4xxPT+h4rYO6taznaLh
vY0AlWWuzGhLIvXctlYRQIwSHZFoOBB65q6eS0JvxIiOvl/A7u1X0fEzZj0EL1d4
ceyqt6g9TB2TQAPT7KkLi033Bq0dvZScR6prM3wskwkL/RCKJ022ftH9o0Ceg9nh
bO4rLkj0Spa98kZURmUGZyKc3MPyrSLv3KUhwDgGb56LyLKy6oLqA6v9dIJk05d9
`protect END_PROTECTED
