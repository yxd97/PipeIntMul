`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ze82lQAwOtyL9JLBf4eIWzjTuLkVv6t641ktvrvmLamla3Tk75mkzJA6d56foPdY
Ph3JM8ouskfJ345KSEH+JFdAJrDKaK0XwdFnBIftbnj2YtKEt7LrtHkkh+XeAVGY
t+GmISbEufxFbLwJtE1PmuFCk2UDpWuj+dcrtRiNP+ctXYlW1OL3SH/A0DDGHncB
Jqt8zGOfZOrQ4FZluNEljwV3QOffbHl5f2th0YdJczApnqXNvI12m4zuvNrV/tcX
QbLVlm0t8d9UlvKtHNJ7mbNPTrJf3NqSq2acb4xdj7/xWk8kuxHuXbTgabbglYoQ
XqdtxpnPncs3Lb5/CLzOuYIhk6oxGSMWjebQoLUXol0SSvY9Co+v2CkRXIhSyiBi
JIqbkbzxAGR0LAo1c2D74g==
`protect END_PROTECTED
