`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTcnHp/liuB7LSe1Y+gV69MFx9Gs7uJef3jbWM6URdSWUUeXO0WMcaFFJSoRNFmS
LRtwLwfuJ0nh3W+DXtYY6T4ofgMgiVDAlyd0zJVcv9RCd+CZOpBw5wUhBOYFKUaz
iCn+tZtt9ZBBKiCZ6nS1tW9zDq/UOj2nsyE7L0wpdTjred9mjwh9FRm0bgsMNORV
/bP37vSStHfzeH3RJjshJRcrwJ8hn0HQy8IwIEs9UUwUJiyo31mqkhKlMc6iEnMZ
n2R5o/5kDD0yyyKJI8AeS0wiCWP1/cXX9rcJLK9HS5tQFFx0fv9B+qZU4+1JJXjT
PmXMYgvnn2uEmn1bDFVcNUQLJI/MFDVHv22dUKII2dLRF+2NYtituRXBrAFdjeJU
wzw7pVWU1C1d3kljfzBpUsbTQrqOsPMyQpmIjR4obS/m3qyrHO9aAQ/ZaE9Fo1Az
iVJJm2vK2Ccw5cWG6XeBdzJNI73ccvmCl8HI2iG6vK7DC3xwGDUzyoYGSccBwJ9F
mhBbj3bK7urRAO05nDumlXzZ/ZxeF9F0QG/l+ryNNrk7OrWsh/OxuU7vAW32f1IL
n+sfU4K4kppi/QRgcfPBHhdVTprySvSBdF+mts3SduBuezKfvHkfDSscUixAPnpK
GOOR2SgCYS3OVmOvp3aEhU2fbjBjnkR+YQU12EoaXUyKl9UqBTpKk0segtpx5POd
w2DDfmXFyb06qyCXUFK0gAxR8gcAubFqCKs3orzpDYl2yZ0Zpw11KitNBf9W+iH2
n67tl7RoSC5HCeY+a3VdBYB1j/OoT1fE0syuVW+6bsKQu8r2I8g5RiFZboSBjGTb
2kb8i2tl9uhI4Wepl4E8qaYhhgzl4V1fVU0v21GWSGkKnY8JifhxMo0v+O6+x4nG
Ap7QqRQFCmZmCceI/p6F2tfiR6xuFgpDjlcehsSA66g=
`protect END_PROTECTED
