`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gfitt/LBQ5LkzZFQLpwNI3ixon592mGuqCdub4yLrXX2+66PA6i+QbPs7BmWEVUR
pBRO7QEfhNyIRqJ8Z+L6K+iQSR26yh01KyXaGKwxAFQGERUGXZnr3REFm2EQqOUO
Z31h8zXbzTRzVHqMBYLpuRWUoljpSUx7PKMANSPyzFZbZG57nRUcqCLH/MIbPcy6
3jU94gpZ2O7b9E9Fnhpt8xRmz15fTJNjstF3cd+OqroekDh/LD/wktNdTwFzlo1F
0Zec5nQzzuO8U1XamTvi8ILB6dsFHoOK3VDkMKHyqrW1sYxkDGXZC6HQ6IBemOtH
/sp8Bz6zu+U+j4c0+P94zUX35KUqV4FNim7zpfqBrWve1t9lazkjpK9F/V3EBDPC
RlqFm4Ri0AOvTftAHT2bQs085gWNJGks/Yh6r9PkMFCgcKSBxHxz4QLJVDrXccSB
HdBQBzJI989AWioT96T+ZEtAYyzjtXbmsbOYr18ePLZGnySsOLNuovMWhUCVF5HB
ItVNzXPyNjmiYXQMXRC3lWy+SuDvzpMDtK18B/dfDv0NppxKK2FLo9qT/MaD8BYp
CvcTYbXtflFnuhMGleprS9/J9hFAspHrrAaaPk8Lr4kSlhjZ+jig5z6jgGfPmsaE
4fSPN54+B5whLYW/IS9/ezdjMRRMiuKRbqOEnDxUZk4qUy0NV5lNIEi9wtKXF0hd
Bn9uQo3xEKqQz/MLc2zsCPivP5oq/lAvG9L+3iCgFkO62NEauLJr+fWAvzO5BSLy
s+Dk1VYDBtd2VtlaKGYMJ6lJfC5bNrqm63eeXXgbJbGCvbkljG/9F46kR0sNz3Zb
NSgqy2fcPe+J1l13GC5oUmTYn/f5oQ59p6NY0M1lZ92NANz1hZiZmLwTJqurwKo8
tOHIzzdp/mfW7RdMISuIaVaTEsVYWIuIKsKrBF6TmX4aQurPz9BJRh6l5rxg/s8Z
Z+hNBGW+oiA/0G4BC3cv6hhmicP2g6QwpSNHLcA+A1x8jMeWu14BSKvYdqL+SFPf
Il5ktr9ZVEhmhOmxn4MxtAI9xxPgOqUdRi6uRAjHujRn+yFzYUjYEVs6rGvFwKW+
c2+2tKLZeHPKB0OoiBkfBZFcbxvDkSzNV177x4xZp4cuumLa11+vBu19Z2xHBU0b
tSU33OffUew3MPFfAcVyofZJie+VDZmNMepAlgWKdOKTG5k6ZIfH8WW1HPqnRoLD
07mqB36eIR/NQgXqZVtiOTNjYIOpFXkZ0wXEtH90lJDK22M5n6INnDcepk85s40F
8rB2rYi12uH4QVd0iIBuqQ==
`protect END_PROTECTED
