`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3z58n6yMfDpYBidQhyCU8XnB2YeGnXdj2QMCmPuh3FTIfgWClVmZSxwaD+kHP6k4
LUKEDFiEww50udua5crONlI7EAuJhfCowwZqvD9+tXWN4/LEca5pN4xIRBSOiMdV
y1jYZ2HcOXq3fYz526PgoCB1Mz3xkOV2D3im5SxZWscPTQ6x5Ar1iF/dvisMnTeC
H3VHvXfWT+mjRAdl+V4H1FhbDaw3yXSnlcFq+KMD1UJxJ74NnXLLoXo3F2b3BcWu
L/KUPl1KgRuGaI5gxvDTMQt0d+6sBhTnD3vu+22r94724fR+sYYkf57vAgbFWfZw
TJjfu4f0U5dc+j4eMuJJesFB0mbUUaDLWzE6qmIEwR0=
`protect END_PROTECTED
