`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UdPmgjwnN0IgGUHtiJLuw5q6ppgrJyFGYtS3lcYciAaN+kMezkIPZRU3cqJoT7Mu
GGo3KfoIrWMYyBhKL3f8fZT8FqeLPNDiuqjn7x5fsfTevthpkEkG2pdLk/gWINbH
F7hDnUdXsxZYARdF5+0uyVNNbqAE4ogf8a5cUVi6n1njWtu6ZipMmunZ/3PXNsHs
mvA0vt2jeJGneN+04xXIw9m7aGPq45NNAtcj5boCyNtV0fuNJUFmuj8Y5xFIQqQT
dZI4y+H+ZVZMeKi2gH1dWb/FgJIliSNKI5g5XMJ/Raj1hkuhCM5pct383blZcPMl
3P4cknDMqY0lJQos+D/mvSM11fUuMQ1NRhu7f1LSet9rXknh8xkP62v7bPHw3KEe
ffDzvzfvgq4cwoV1tSIS3AxPPjDS6gZ/C4FRpcUJe4eBVR4rjxwPpyU6rBQwGj47
I94sg2JAb5NXok8Kcjhnb3W2FC3zs/VnIFg3luMyCKI6BLodUF4QRzk4R5FFGkdN
5tK5f4WnbiNQvRSsUEkhJEZKOn7QDRzQO9+eDH1lrNSRpPr4u8pSLmX71x7AhnpY
XUDUDkETpEH92uP/BVSTJ833FLstjUR8RX2x1NT6fdizVgHhh+x5DYfG/JmNsWAM
Aif+Y615jR9jQ1Z9gmdF818JxzesflaRecvF1XjWb6hMGT8cT7vRCN+KiVSoX3kp
1QSPIFPduepyW8ANifyyYikPsiScWsrXYawKBuuA5DV6/Pkg1/1uaYYdY9DrBfdH
zklgI2AJHcQryDVXbF1qDLQGFu1Ng1Zba5JrgqgRT0Z+mtWbtxkVN+yLL+PkYO4P
09ZQxdagcgZQ8AGg/GWRLPUhYe7GsPCyiG5ymfMg8XegilOeBGfaVL8aInRL6vlG
lOOAt7umMXgW3OjFN+bFSRryQoMZLzF83QiiPLDD3eoxdN7dC2I2YGh3nlzi7dMd
Pw8wviOGHeSfY+RJooPJqIfkI3POHG9aKnR9tuY8Kh6lsAy/5hT89KS5W0K4lMFk
BOs4Zw6J0wYad8j309Hekyj4B+DMgWGa2qJe/6CB5JC/aXUuo349P1jPo9kIFfPZ
4zXX0+JoHUSLBrImMnYoBjsBBjir48w4p9vmaw54dpLEUX+eSZw/rop2Kxd8Fmce
5i7eVzpJZA/EtJwDgq3AyjcUuZSpk4dI0TUVA5cOkMtGYb288IQ41zwng0kJThgN
lUSed+lVx0ZDaCXDXd6h97xWuALa3+x/ZMO8/BwwvOTcOl3pSnx9gwbMvwq2P7Hw
nXDwGkKrFWh3f22ZA7UD1OuyHmixEVFvOrmBOCNiE8TblGvs0OGjgbzY6jRh5F07
lY7BNRQPr71qTeBljTikhjiV2Uhcv3UiSk0hYoSW7xV2RZhc2+NS9lmM7HfS6JUt
NWYWLNSbS4dgvDLof6j/jqquw1g6UJbs9sKHXinBgR1GuOSexruClrmCoDoqAxxY
syYBP90pPcKfSq1858OXmrIBTY3niyeD5LLW3i2mCB1EMaFZRUHJv1vlodxo5ymB
pyMx1WfZTztYhEqqGCj+BQqvtpQPJ6ELNuYoMGozy7GsRo3diQx4flMkW3HaZs21
Wt08AF4unP6FXG96jUmzQIflkhqkCTAX2LZPE12vgXNeE7GgFDjXgIGvMNtZKS2D
F3d3Y6eDSHRCPQJwRg9de9GqazLIGVovYZOYSi7kOR0IMXs3egV0cg3dLJxfhaSA
3Nv+0FPXRAdvM2pZMd6DG0MyjplbV5O44apr2AfSP9cjIU9iSY+zI43d+828+8lc
WakuVz8SCarHH/IeLUhfjSNE7SCTb9+z0zHxqQ84aZjRD8B9Dqh+VQzcU3g/fJpS
kyUeOw3ID4GjqXrbjiEn2OC/kKO7wcIRxsSOdJIUtOS/rkHAo3x5dAP+lk5nvTDR
QIXQKbMl/rpQBFyYnJCwBcRX8moj1O8qZHmcKm/apwqGRy2zvx1VgtCevFHH5aeX
vhsfaHrD5RtQyaZMuRTllGVdOonOL111pXlNvzDvcZaVm9S/rv5H5EK4v1rPLLpy
u78F18kbKs1R044k9ltfrKkBaxneUbduoo1ia0wf4Iu2jsvD5enalTNUTKnNaeMj
ZEjqVdq6i6f0K54eFK5Vrf8+26FDCdlD9YF3ZU1+Q15x0ShobuQ6Ax06+X4lRDzj
tWSR1p/M1RYauK9xwoKIWrMh4e5Njqw5hTWpnPmHlqvSnGHgDRfXfDjEU+QmybdZ
Nbq6v0UwELaIL75iAWxXv6/N1zy/b7BwZwAP7Bc+o/DTUY2DyGfB6NczQogzx7vq
gZWNcvbw5bdGWH2XYyAnZotmA9By7GqQcMa5SsCWBaIQBp0CuHjImQg4u7JzmKso
sIYFMW9DLfW861g/Z3wgXxrMa6o8pA+5hx0mPNo4Wkjo7R7KuFb0J34ZsTLsDnxh
7VVhjvV8AjgQGuHo3TQfBV0fGcv04MpngtlLxvBb7Dc=
`protect END_PROTECTED
