`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwcEg+wk5PasoSnY957WDUdwAylMRchGc2SKst2XmI6kTOlUnG342VpF9ueenw+6
s2sOQIrrU6+2B976G5Ty6swwXHlcsvYfDvwyQsFRpg5hyF5j7UiahSSh6CRjHea5
dB1igN0XffNXEGGkA+ccGwVgL8sGV2SHT8J+NKM8jWugOWl7ZtFwl69mEIL49Vhl
UgPYHXUwVlKLAu22Ulfz42eNV5Jd6czK4mwGbdRDSXbCjgb18xuCQScOmbuRzF53
qmC+Ho+Q9JHUvDeh2esUPWGbaHu+WaH/kB0nAnz1ZktIhGuKtqJVyWRv3I8Or8hw
ceOov0yh2va1uBqC7wHLURArSixbybhWZ74wOrKwztnBzgcmfRPqITpdgIn2+A/D
FNhQOFe+CoaMbxcviKTRbnNOw4XCvifkgHmzuzGMb1zBC0WdIrscvexlf15lyVJZ
Va4uhbW8AmKt3KeYyQLkbJoTWp/uLu2PB1EdB56P5zPzFswMGsHVznQbk6TC+1Wi
jRv2rhJgtRJWFacJI+5dwQFNJFTT7BfC3/90J4nE5rQ/5aNiVOFM0Q6xReiH+Fgk
PeNfZmO0+nk+C7Y1CVaSmejIqvZMT1PGsYVtXh0N+ALyDinhfcngjgleaaTFtyN1
UE1u+PARcL8iCZf3/btxXfEiYAvnR0QQTB6f7GsfDF9Vl8+U8rtZtcnd2yfcLWPE
IpxAy5IegWp5WzIdkC4tVGpa5R5/L4I97BfCNxKzjtfh9d13unz5T0502qCklOR4
nWFnF7Myqd4dv5BvUh/88ZNQnjOdxkX50QqnXO87IqeqLbiPiuP72rprTKtD3Foe
6y8f7R6tDPmPGeDuEiBbAXwQiBWBhMg+zRQIFpjJf9bDXUuLHGIxpLoGpj5RYmMy
UkvxxBOERgscZ0LY438BGyGwGpZLVA2jCJ/1IJxxQMo5d8Pm1pb47iphdwXwKUjU
4bonUAQbZyZ12R9+cgwxPC33lwRhAq1TyS5r2PygmadfbsGoVWGdutpVWMgR6l93
uJArwKMfM3jCrf/T9u4+0um6BRKWl4Wvijkx4++GiKtUSaqw8wpIbY7n7F5++5i0
eo4L91SdER1V2T4jKfPMwTaRKpYF0ZMEf2jj+jur40TlaeCkRaWVNLJZyNh5dB1s
`protect END_PROTECTED
