`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X8AoB9aqQ1YdwKlqjTe/Q4eOqRVaqzuK9al3C/UWj3ZUDvNd6NDbCDafoLsfvoe7
pHbcQwcP+re/lTx7XXX6SJlR6ogCwd1AkUnJiQjLMf2lagek3er9cNlELtR7A6cF
h+UqByNfTh3WyRvOIXJxHgum4g7eCzaXQ+xAmR7x/7pp6Dsf/bURz3M8sqbovA9g
gEE16rpHtY2xteu7q8PvYxGHSYVk+wy8pHsvZsHtc5FPnKFcvg+PXuphVG4amCee
JLiJeFIlWfNQ2D6Vo39UKY9GtdTBCynR1Hk5hgOrdEnf74Q5v+maV0/v2mP2iElm
nDCml2BVkxxEBkDguVDmQQ2dVkihudUmwGnEmQloI2dE21D9acI0tqeB8ST9u6/P
eOVZIi7XBPa28jx800WT/LTNnL9Ex4mZMf5KVhZ89oTLZukOH1aDSy1Fa3GkHM1N
qTq5I7uIBqexo8pcsFi9Cww/cyLQZbLe/7VYZ0VfBhjcck/etDAsUMkA2Apa/Wre
bKHd8HuPYG8WBmDblfMKZQ/+cJJLzI94jWvrw6yM6x6zimOKvHy2oVc8CmLc/As4
`protect END_PROTECTED
