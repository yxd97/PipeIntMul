library verilog;
use verilog.vl_types.all;
entity X_GT11 is
    generic(
        LOC             : string  := "UNPLACED";
        BANDGAPSEL      : string  := "FALSE";
        BIASRESSEL      : string  := "FALSE";
        CCCB_ARBITRATOR_DISABLE: string  := "FALSE";
        CHAN_BOND_MODE  : string  := "NONE";
        CHAN_BOND_ONE_SHOT: string  := "FALSE";
        CHAN_BOND_SEQ_1_1: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_1_2: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_1_3: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_1_4: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_1_MASK: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        CHAN_BOND_SEQ_2_1: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_2_2: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_2_3: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_2_4: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_2_MASK: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        CHAN_BOND_SEQ_2_USE: string  := "FALSE";
        CLK_CORRECT_USE : string  := "FALSE";
        CLK_COR_8B10B_DE: string  := "FALSE";
        CLK_COR_SEQ_1_1 : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_1_2 : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_1_3 : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_1_4 : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_1_MASK: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        CLK_COR_SEQ_2_1 : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_2_2 : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_2_3 : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_2_4 : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_2_MASK: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        CLK_COR_SEQ_2_USE: string  := "FALSE";
        CLK_COR_SEQ_DROP: string  := "FALSE";
        COMMA32         : string  := "FALSE";
        COMMA_10B_MASK  : vl_logic_vector(0 to 9) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        CYCLE_LIMIT_SEL : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        DCDR_FILTER     : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        DEC_MCOMMA_DETECT: string  := "TRUE";
        DEC_PCOMMA_DETECT: string  := "TRUE";
        DEC_VALID_COMMA_ONLY: string  := "TRUE";
        DIGRX_FWDCLK    : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        DIGRX_SYNC_MODE : string  := "FALSE";
        ENABLE_DCDR     : string  := "FALSE";
        FDET_HYS_CAL    : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        FDET_HYS_SEL    : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        FDET_LCK_CAL    : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        FDET_LCK_SEL    : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        GT11_MODE       : string  := "DONT_CARE";
        IREFBIASMODE    : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        LOOPCAL_WAIT    : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        MCOMMA_32B_VALUE: integer := 0;
        MCOMMA_DETECT   : string  := "TRUE";
        OPPOSITE_SELECT : string  := "FALSE";
        PCOMMA_32B_VALUE: integer := 0;
        PCOMMA_DETECT   : string  := "TRUE";
        PCS_BIT_SLIP    : string  := "FALSE";
        PMACLKENABLE    : string  := "TRUE";
        PMACOREPWRENABLE: string  := "TRUE";
        PMAIREFTRIM     : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        PMAVBGCTRL      : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PMAVREFTRIM     : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        PMA_BIT_SLIP    : string  := "FALSE";
        POWER_ENABLE    : string  := "TRUE";
        REPEATER        : string  := "FALSE";
        RXACTST         : string  := "FALSE";
        RXAFEEQ         : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXAFEPD         : string  := "FALSE";
        RXAFETST        : string  := "FALSE";
        RXAPD           : string  := "FALSE";
        RXAREGCTRL      : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        RXASYNCDIVIDE   : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        RXBY_32         : string  := "FALSE";
        RXCDRLOS        : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXCLK0_FORCE_PMACLK: string  := "FALSE";
        RXCLKMODE       : vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        RXCLMODE        : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        RXCMADJ         : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        RXCPSEL         : string  := "TRUE";
        RXCPTST         : string  := "FALSE";
        RXCRCCLOCKDOUBLE: string  := "FALSE";
        RXCRCENABLE     : string  := "FALSE";
        RXCRCINITVAL    : integer := 0;
        RXCRCINVERTGEN  : string  := "FALSE";
        RXCRCSAMECLOCK  : string  := "FALSE";
        RXCTRL1         : vl_logic_vector(0 to 9) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXCYCLE_LIMIT_SEL: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        RXDATA_SEL      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        RXDCCOUPLE      : string  := "FALSE";
        RXDIGRESET      : string  := "FALSE";
        RXDIGRX         : string  := "FALSE";
        RXEQ            : vl_logic_vector(0 to 63) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXFDCAL_CLOCK_DIVIDE: string  := "NONE";
        RXFDET_HYS_CAL  : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        RXFDET_HYS_SEL  : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        RXFDET_LCK_CAL  : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        RXFDET_LCK_SEL  : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        RXFECONTROL1    : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        RXFECONTROL2    : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        RXFETUNE        : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        RXLB            : string  := "FALSE";
        RXLKADJ         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        RXLKAPD         : string  := "FALSE";
        RXLOOPCAL_WAIT  : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        RXLOOPFILT      : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        RXMODE          : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXPD            : string  := "FALSE";
        RXPDDTST        : string  := "TRUE";
        RXPMACLKSEL     : string  := "REFCLK1";
        RXRCPADJ        : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        RXRCPPD         : string  := "FALSE";
        RXRECCLK1_USE_SYNC: string  := "FALSE";
        RXRIBADJ        : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        RXRPDPD         : string  := "FALSE";
        RXRSDPD         : string  := "FALSE";
        RXSLOWDOWN_CAL  : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        RXTUNE          : vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXVCODAC_INIT   : vl_logic_vector(0 to 9) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXVCO_CTRL_ENABLE: string  := "FALSE";
        RX_BUFFER_USE   : string  := "TRUE";
        RX_CLOCK_DIVIDER: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        SAMPLE_8X       : string  := "FALSE";
        SLOWDOWN_CAL    : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        TXABPMACLKSEL   : string  := "REFCLK1";
        TXAPD           : string  := "FALSE";
        TXAREFBIASSEL   : string  := "TRUE";
        TXASYNCDIVIDE   : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        TXCLK0_FORCE_PMACLK: string  := "FALSE";
        TXCLKMODE       : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        TXCLMODE        : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        TXCPSEL         : string  := "TRUE";
        TXCRCCLOCKDOUBLE: string  := "FALSE";
        TXCRCENABLE     : string  := "FALSE";
        TXCRCINITVAL    : integer := 0;
        TXCRCINVERTGEN  : string  := "FALSE";
        TXCRCSAMECLOCK  : string  := "FALSE";
        TXCTRL1         : vl_logic_vector(0 to 9) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TXDATA_SEL      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        TXDAT_PRDRV_DAC : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        TXDAT_TAP_DAC   : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi0);
        TXDIGPD         : string  := "FALSE";
        TXFDCAL_CLOCK_DIVIDE: string  := "NONE";
        TXHIGHSIGNALEN  : string  := "TRUE";
        TXLOOPFILT      : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        TXLVLSHFTPD     : string  := "FALSE";
        TXOUTCLK1_USE_SYNC: string  := "FALSE";
        TXPD            : string  := "FALSE";
        TXPHASESEL      : string  := "FALSE";
        TXPOST_PRDRV_DAC: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        TXPOST_TAP_DAC  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi0);
        TXPOST_TAP_PD   : string  := "TRUE";
        TXPRE_PRDRV_DAC : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        TXPRE_TAP_DAC   : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        TXPRE_TAP_PD    : string  := "TRUE";
        TXSLEWRATE      : string  := "FALSE";
        TXTERMTRIM      : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        TXTUNE          : vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TX_BUFFER_USE   : string  := "TRUE";
        TX_CLOCK_DIVIDER: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        VCODAC_INIT     : vl_logic_vector(0 to 9) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VCO_CTRL_ENABLE : string  := "FALSE";
        VREFBIASMODE    : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        ALIGN_COMMA_WORD: integer := 4;
        CHAN_BOND_LIMIT : integer := 16;
        CHAN_BOND_SEQ_LEN: integer := 1;
        CLK_COR_MAX_LAT : integer := 48;
        CLK_COR_MIN_LAT : integer := 36;
        CLK_COR_SEQ_LEN : integer := 1;
        RXOUTDIV2SEL    : integer := 1;
        RXPLLNDIVSEL    : integer := 8;
        RXUSRDIVISOR    : integer := 1;
        SH_CNT_MAX      : integer := 64;
        SH_INVALID_CNT_MAX: integer := 16;
        TXOUTDIV2SEL    : integer := 1;
        TXPLLNDIVSEL    : integer := 8
    );
    port(
        CHBONDO         : out    vl_logic_vector(4 downto 0);
        COMBUSOUT       : out    vl_logic_vector(15 downto 0);
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        RXBUFERR        : out    vl_logic;
        RXCALFAIL       : out    vl_logic;
        RXCHARISCOMMA   : out    vl_logic_vector(7 downto 0);
        RXCHARISK       : out    vl_logic_vector(7 downto 0);
        RXCOMMADET      : out    vl_logic;
        RXCRCOUT        : out    vl_logic_vector(31 downto 0);
        RXCYCLELIMIT    : out    vl_logic;
        RXDATA          : out    vl_logic_vector(63 downto 0);
        RXDISPERR       : out    vl_logic_vector(7 downto 0);
        RXLOCK          : out    vl_logic;
        RXLOSSOFSYNC    : out    vl_logic_vector(1 downto 0);
        RXMCLK          : out    vl_logic;
        RXNOTINTABLE    : out    vl_logic_vector(7 downto 0);
        RXPCSHCLKOUT    : out    vl_logic;
        RXREALIGN       : out    vl_logic;
        RXRECCLK1       : out    vl_logic;
        RXRECCLK2       : out    vl_logic;
        RXRUNDISP       : out    vl_logic_vector(7 downto 0);
        RXSIGDET        : out    vl_logic;
        RXSTATUS        : out    vl_logic_vector(5 downto 0);
        TX1N            : out    vl_logic;
        TX1P            : out    vl_logic;
        TXBUFERR        : out    vl_logic;
        TXCALFAIL       : out    vl_logic;
        TXCRCOUT        : out    vl_logic_vector(31 downto 0);
        TXCYCLELIMIT    : out    vl_logic;
        TXKERR          : out    vl_logic_vector(7 downto 0);
        TXLOCK          : out    vl_logic;
        TXOUTCLK1       : out    vl_logic;
        TXOUTCLK2       : out    vl_logic;
        TXPCSHCLKOUT    : out    vl_logic;
        TXRUNDISP       : out    vl_logic_vector(7 downto 0);
        CHBONDI         : in     vl_logic_vector(4 downto 0);
        COMBUSIN        : in     vl_logic_vector(15 downto 0);
        DADDR           : in     vl_logic_vector(7 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        ENCHANSYNC      : in     vl_logic;
        ENMCOMMAALIGN   : in     vl_logic;
        ENPCOMMAALIGN   : in     vl_logic;
        GREFCLK         : in     vl_logic;
        LOOPBACK        : in     vl_logic_vector(1 downto 0);
        POWERDOWN       : in     vl_logic;
        REFCLK1         : in     vl_logic;
        REFCLK2         : in     vl_logic;
        RX1N            : in     vl_logic;
        RX1P            : in     vl_logic;
        RXBLOCKSYNC64B66BUSE: in     vl_logic;
        RXCLKSTABLE     : in     vl_logic;
        RXCOMMADETUSE   : in     vl_logic;
        RXCRCCLK        : in     vl_logic;
        RXCRCDATAVALID  : in     vl_logic;
        RXCRCDATAWIDTH  : in     vl_logic_vector(2 downto 0);
        RXCRCIN         : in     vl_logic_vector(63 downto 0);
        RXCRCINIT       : in     vl_logic;
        RXCRCINTCLK     : in     vl_logic;
        RXCRCPD         : in     vl_logic;
        RXCRCRESET      : in     vl_logic;
        RXDATAWIDTH     : in     vl_logic_vector(1 downto 0);
        RXDEC64B66BUSE  : in     vl_logic;
        RXDEC8B10BUSE   : in     vl_logic;
        RXDESCRAM64B66BUSE: in     vl_logic;
        RXIGNOREBTF     : in     vl_logic;
        RXINTDATAWIDTH  : in     vl_logic_vector(1 downto 0);
        RXPMARESET      : in     vl_logic;
        RXPOLARITY      : in     vl_logic;
        RXRESET         : in     vl_logic;
        RXSLIDE         : in     vl_logic;
        RXSYNC          : in     vl_logic;
        RXUSRCLK        : in     vl_logic;
        RXUSRCLK2       : in     vl_logic;
        TXBYPASS8B10B   : in     vl_logic_vector(7 downto 0);
        TXCHARDISPMODE  : in     vl_logic_vector(7 downto 0);
        TXCHARDISPVAL   : in     vl_logic_vector(7 downto 0);
        TXCHARISK       : in     vl_logic_vector(7 downto 0);
        TXCLKSTABLE     : in     vl_logic;
        TXCRCCLK        : in     vl_logic;
        TXCRCDATAVALID  : in     vl_logic;
        TXCRCDATAWIDTH  : in     vl_logic_vector(2 downto 0);
        TXCRCIN         : in     vl_logic_vector(63 downto 0);
        TXCRCINIT       : in     vl_logic;
        TXCRCINTCLK     : in     vl_logic;
        TXCRCPD         : in     vl_logic;
        TXCRCRESET      : in     vl_logic;
        TXDATA          : in     vl_logic_vector(63 downto 0);
        TXDATAWIDTH     : in     vl_logic_vector(1 downto 0);
        TXENC64B66BUSE  : in     vl_logic;
        TXENC8B10BUSE   : in     vl_logic;
        TXENOOB         : in     vl_logic;
        TXGEARBOX64B66BUSE: in     vl_logic;
        TXINHIBIT       : in     vl_logic;
        TXINTDATAWIDTH  : in     vl_logic_vector(1 downto 0);
        TXPMARESET      : in     vl_logic;
        TXPOLARITY      : in     vl_logic;
        TXRESET         : in     vl_logic;
        TXSCRAM64B66BUSE: in     vl_logic;
        TXSYNC          : in     vl_logic;
        TXUSRCLK        : in     vl_logic;
        TXUSRCLK2       : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOC : constant is 1;
    attribute mti_svvh_generic_type of BANDGAPSEL : constant is 1;
    attribute mti_svvh_generic_type of BIASRESSEL : constant is 1;
    attribute mti_svvh_generic_type of CCCB_ARBITRATOR_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_MODE : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_ONE_SHOT : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_1 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_2 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_3 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_4 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_MASK : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_1 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_2 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_3 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_4 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_MASK : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_USE : constant is 1;
    attribute mti_svvh_generic_type of CLK_CORRECT_USE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_8B10B_DE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_1 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_2 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_3 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_4 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_MASK : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_1 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_2 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_3 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_4 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_MASK : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_USE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_DROP : constant is 1;
    attribute mti_svvh_generic_type of COMMA32 : constant is 1;
    attribute mti_svvh_generic_type of COMMA_10B_MASK : constant is 1;
    attribute mti_svvh_generic_type of CYCLE_LIMIT_SEL : constant is 1;
    attribute mti_svvh_generic_type of DCDR_FILTER : constant is 1;
    attribute mti_svvh_generic_type of DEC_MCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of DEC_PCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of DEC_VALID_COMMA_ONLY : constant is 1;
    attribute mti_svvh_generic_type of DIGRX_FWDCLK : constant is 1;
    attribute mti_svvh_generic_type of DIGRX_SYNC_MODE : constant is 1;
    attribute mti_svvh_generic_type of ENABLE_DCDR : constant is 1;
    attribute mti_svvh_generic_type of FDET_HYS_CAL : constant is 1;
    attribute mti_svvh_generic_type of FDET_HYS_SEL : constant is 1;
    attribute mti_svvh_generic_type of FDET_LCK_CAL : constant is 1;
    attribute mti_svvh_generic_type of FDET_LCK_SEL : constant is 1;
    attribute mti_svvh_generic_type of GT11_MODE : constant is 1;
    attribute mti_svvh_generic_type of IREFBIASMODE : constant is 1;
    attribute mti_svvh_generic_type of LOOPCAL_WAIT : constant is 1;
    attribute mti_svvh_generic_type of MCOMMA_32B_VALUE : constant is 1;
    attribute mti_svvh_generic_type of MCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of OPPOSITE_SELECT : constant is 1;
    attribute mti_svvh_generic_type of PCOMMA_32B_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of PCS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PMACLKENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMACOREPWRENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMAIREFTRIM : constant is 1;
    attribute mti_svvh_generic_type of PMAVBGCTRL : constant is 1;
    attribute mti_svvh_generic_type of PMAVREFTRIM : constant is 1;
    attribute mti_svvh_generic_type of PMA_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of POWER_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of REPEATER : constant is 1;
    attribute mti_svvh_generic_type of RXACTST : constant is 1;
    attribute mti_svvh_generic_type of RXAFEEQ : constant is 1;
    attribute mti_svvh_generic_type of RXAFEPD : constant is 1;
    attribute mti_svvh_generic_type of RXAFETST : constant is 1;
    attribute mti_svvh_generic_type of RXAPD : constant is 1;
    attribute mti_svvh_generic_type of RXAREGCTRL : constant is 1;
    attribute mti_svvh_generic_type of RXASYNCDIVIDE : constant is 1;
    attribute mti_svvh_generic_type of RXBY_32 : constant is 1;
    attribute mti_svvh_generic_type of RXCDRLOS : constant is 1;
    attribute mti_svvh_generic_type of RXCLK0_FORCE_PMACLK : constant is 1;
    attribute mti_svvh_generic_type of RXCLKMODE : constant is 1;
    attribute mti_svvh_generic_type of RXCLMODE : constant is 1;
    attribute mti_svvh_generic_type of RXCMADJ : constant is 1;
    attribute mti_svvh_generic_type of RXCPSEL : constant is 1;
    attribute mti_svvh_generic_type of RXCPTST : constant is 1;
    attribute mti_svvh_generic_type of RXCRCCLOCKDOUBLE : constant is 1;
    attribute mti_svvh_generic_type of RXCRCENABLE : constant is 1;
    attribute mti_svvh_generic_type of RXCRCINITVAL : constant is 1;
    attribute mti_svvh_generic_type of RXCRCINVERTGEN : constant is 1;
    attribute mti_svvh_generic_type of RXCRCSAMECLOCK : constant is 1;
    attribute mti_svvh_generic_type of RXCTRL1 : constant is 1;
    attribute mti_svvh_generic_type of RXCYCLE_LIMIT_SEL : constant is 1;
    attribute mti_svvh_generic_type of RXDATA_SEL : constant is 1;
    attribute mti_svvh_generic_type of RXDCCOUPLE : constant is 1;
    attribute mti_svvh_generic_type of RXDIGRESET : constant is 1;
    attribute mti_svvh_generic_type of RXDIGRX : constant is 1;
    attribute mti_svvh_generic_type of RXEQ : constant is 1;
    attribute mti_svvh_generic_type of RXFDCAL_CLOCK_DIVIDE : constant is 1;
    attribute mti_svvh_generic_type of RXFDET_HYS_CAL : constant is 1;
    attribute mti_svvh_generic_type of RXFDET_HYS_SEL : constant is 1;
    attribute mti_svvh_generic_type of RXFDET_LCK_CAL : constant is 1;
    attribute mti_svvh_generic_type of RXFDET_LCK_SEL : constant is 1;
    attribute mti_svvh_generic_type of RXFECONTROL1 : constant is 1;
    attribute mti_svvh_generic_type of RXFECONTROL2 : constant is 1;
    attribute mti_svvh_generic_type of RXFETUNE : constant is 1;
    attribute mti_svvh_generic_type of RXLB : constant is 1;
    attribute mti_svvh_generic_type of RXLKADJ : constant is 1;
    attribute mti_svvh_generic_type of RXLKAPD : constant is 1;
    attribute mti_svvh_generic_type of RXLOOPCAL_WAIT : constant is 1;
    attribute mti_svvh_generic_type of RXLOOPFILT : constant is 1;
    attribute mti_svvh_generic_type of RXMODE : constant is 1;
    attribute mti_svvh_generic_type of RXPD : constant is 1;
    attribute mti_svvh_generic_type of RXPDDTST : constant is 1;
    attribute mti_svvh_generic_type of RXPMACLKSEL : constant is 1;
    attribute mti_svvh_generic_type of RXRCPADJ : constant is 1;
    attribute mti_svvh_generic_type of RXRCPPD : constant is 1;
    attribute mti_svvh_generic_type of RXRECCLK1_USE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of RXRIBADJ : constant is 1;
    attribute mti_svvh_generic_type of RXRPDPD : constant is 1;
    attribute mti_svvh_generic_type of RXRSDPD : constant is 1;
    attribute mti_svvh_generic_type of RXSLOWDOWN_CAL : constant is 1;
    attribute mti_svvh_generic_type of RXTUNE : constant is 1;
    attribute mti_svvh_generic_type of RXVCODAC_INIT : constant is 1;
    attribute mti_svvh_generic_type of RXVCO_CTRL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of RX_BUFFER_USE : constant is 1;
    attribute mti_svvh_generic_type of RX_CLOCK_DIVIDER : constant is 1;
    attribute mti_svvh_generic_type of SAMPLE_8X : constant is 1;
    attribute mti_svvh_generic_type of SLOWDOWN_CAL : constant is 1;
    attribute mti_svvh_generic_type of TXABPMACLKSEL : constant is 1;
    attribute mti_svvh_generic_type of TXAPD : constant is 1;
    attribute mti_svvh_generic_type of TXAREFBIASSEL : constant is 1;
    attribute mti_svvh_generic_type of TXASYNCDIVIDE : constant is 1;
    attribute mti_svvh_generic_type of TXCLK0_FORCE_PMACLK : constant is 1;
    attribute mti_svvh_generic_type of TXCLKMODE : constant is 1;
    attribute mti_svvh_generic_type of TXCLMODE : constant is 1;
    attribute mti_svvh_generic_type of TXCPSEL : constant is 1;
    attribute mti_svvh_generic_type of TXCRCCLOCKDOUBLE : constant is 1;
    attribute mti_svvh_generic_type of TXCRCENABLE : constant is 1;
    attribute mti_svvh_generic_type of TXCRCINITVAL : constant is 1;
    attribute mti_svvh_generic_type of TXCRCINVERTGEN : constant is 1;
    attribute mti_svvh_generic_type of TXCRCSAMECLOCK : constant is 1;
    attribute mti_svvh_generic_type of TXCTRL1 : constant is 1;
    attribute mti_svvh_generic_type of TXDATA_SEL : constant is 1;
    attribute mti_svvh_generic_type of TXDAT_PRDRV_DAC : constant is 1;
    attribute mti_svvh_generic_type of TXDAT_TAP_DAC : constant is 1;
    attribute mti_svvh_generic_type of TXDIGPD : constant is 1;
    attribute mti_svvh_generic_type of TXFDCAL_CLOCK_DIVIDE : constant is 1;
    attribute mti_svvh_generic_type of TXHIGHSIGNALEN : constant is 1;
    attribute mti_svvh_generic_type of TXLOOPFILT : constant is 1;
    attribute mti_svvh_generic_type of TXLVLSHFTPD : constant is 1;
    attribute mti_svvh_generic_type of TXOUTCLK1_USE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of TXPD : constant is 1;
    attribute mti_svvh_generic_type of TXPHASESEL : constant is 1;
    attribute mti_svvh_generic_type of TXPOST_PRDRV_DAC : constant is 1;
    attribute mti_svvh_generic_type of TXPOST_TAP_DAC : constant is 1;
    attribute mti_svvh_generic_type of TXPOST_TAP_PD : constant is 1;
    attribute mti_svvh_generic_type of TXPRE_PRDRV_DAC : constant is 1;
    attribute mti_svvh_generic_type of TXPRE_TAP_DAC : constant is 1;
    attribute mti_svvh_generic_type of TXPRE_TAP_PD : constant is 1;
    attribute mti_svvh_generic_type of TXSLEWRATE : constant is 1;
    attribute mti_svvh_generic_type of TXTERMTRIM : constant is 1;
    attribute mti_svvh_generic_type of TXTUNE : constant is 1;
    attribute mti_svvh_generic_type of TX_BUFFER_USE : constant is 1;
    attribute mti_svvh_generic_type of TX_CLOCK_DIVIDER : constant is 1;
    attribute mti_svvh_generic_type of VCODAC_INIT : constant is 1;
    attribute mti_svvh_generic_type of VCO_CTRL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of VREFBIASMODE : constant is 1;
    attribute mti_svvh_generic_type of ALIGN_COMMA_WORD : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_LIMIT : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_LEN : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_MAX_LAT : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_MIN_LAT : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_LEN : constant is 2;
    attribute mti_svvh_generic_type of RXOUTDIV2SEL : constant is 2;
    attribute mti_svvh_generic_type of RXPLLNDIVSEL : constant is 2;
    attribute mti_svvh_generic_type of RXUSRDIVISOR : constant is 2;
    attribute mti_svvh_generic_type of SH_CNT_MAX : constant is 2;
    attribute mti_svvh_generic_type of SH_INVALID_CNT_MAX : constant is 2;
    attribute mti_svvh_generic_type of TXOUTDIV2SEL : constant is 2;
    attribute mti_svvh_generic_type of TXPLLNDIVSEL : constant is 2;
end X_GT11;
