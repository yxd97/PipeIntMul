`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pjrmAO/jLAcxjIWTv8ABNTtSUMQ+mEAr2CMFeeypkNi3H4br5encqrgu4S6pXMzr
5IlPKn1erOQY9LHd3VzKZJCdi1bMThaYqGSTjBFq/l3L0MQV4NEVq/UQtaO2t+Lh
fpF/6aQwqXY7KsI2kPrW62dIBDuPKR6Nz5nrqX3W8iq0UlSDiCRLCYd2mKqNrUhn
uBr6IjHUyr7yOIqMPflLq/DjWnksaoh3ZTCUfsJuMaaE2A+wjAIGUXQ8BlXwMcO+
eAnCKdCLynJg8ydYdGy83CifkrZkOCWFCczyveBLYbyR/whyze+RRYs1PEeYskNI
NwfyCoQtCIi+8hXHcX4L8w2oZTiIKFHcZ3AoGbwnsbykNGf9rilHVRaQ+pXR7miG
MRtTPC59+7O6UQRA0g1cEp8RY6cVyrN8ByRWIvzMWsWQYUpsT1CZ1on3rXO+1rbq
CNdSJl6Xdk/n0SAT+6fbDMCErQBY75rEbCvr/IOUZsx56e47hlMlMd2xbthV8Xmo
`protect END_PROTECTED
