`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGOqagoR6TwYrK0puRoZOGXaBRzASs6jkVg2Himtk/GGjaYGkD7ddlkgPHK1Ada4
dhjkTPwTdq6MINUZ4w/qYjPFsGRU8OUJ8CcKXUKALQ+m4tCxZjS5e+cUUc8Z5K5j
Nes7T2PsnFc27+peR0+VJGkerN6xyN+iBwhK0yQf5Zvi838afoW2zZT86ShriCOu
IsE3pxhHTzCqEftki8A2y9b/wdNkGxyvMm2oD77+Jf/Nmtp3IqrcHSobluraNo7+
eouFGFWepJ2ZuOiQFwRILIHYEJ4YQP8o8/Rt68W1pYRxkGoTDWVN4edjBjCbwBSb
8eYWnuMk+XuMaUy/emagG03sNxRQ9pfGkY6X1UJ/U4LwXXXNafMc6Lb63YZxIpuF
`protect END_PROTECTED
