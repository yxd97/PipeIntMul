`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kvjALrxD7JU+3ZHFuwjHSPwwLryI/76Iu3EaGN6HMe1mW+ZLAlehPpBXG5xY3NhX
U52kE2hGz8m/WoKeaLhymGEuBVzYGNTxCM2+Q9+/mD28HYQ8doDBWN36T9eUmW5S
F1wNCza8aSgdfpqCSXl1MMrRzx4kbE7NjsJK4I8aZNIXBI7M5CaesFUEhXS81KZg
LQ876LLOnuNOwAlxGiAH/xdb2DVtRcuVYB0lub/CtfNXz28xxcBQjuTz/LnOZ67D
G3haNqhM+InlOIpIFLoD2KPN03UR1/IcmpK747asEL1RAg7C0w0xd4M5v8rSVhSJ
MKWgM6+Botaf0F2IK25YDn0KrRKzRyC1ew5+bPj01g16qr2RVx1AFMvyjW6jOAIo
5P1zpKC7WcmpByNevTdyKxLQTKcSsctgBAfeMjUbwSBF0iXuT3vAfR00NAweMZpX
PkyAd+kruXiGFiKUlsABfV5eDmj5sVsFb/dnUwh0FrfXs9wRFc4FaF6rkivUSBpS
DqHYJOc5tfLtAURrk0pnwud6jbteK7G8eUyM5oP+H1nOwVJ03xWx0ttU08mHjQpY
H3wLXO8aQH7v98E6hknQTg==
`protect END_PROTECTED
