`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pm7IMA2qza0XMfx+UfTPR8D0VPRCk8wQkveLk0UQHMPLiV4l77rilT/PpBnRYu6W
utMZ2iuzWSjLk6pGfxnqhcDmVIPO3XlZkQTyJemKZby/Rj/lG5y3alox6+/mbrtM
8Ih0zY1n+Zp9+vJOsUpd39lE92p86dak0tiH+e3zFyzr2eg9ZL4KSqFBfBMMmDKt
w04JeaKhT06UfCGHLYUr8Xn9rvSFvTWnSdbWWo1XLjwQ2pNVDjr8vgz7utLpdYTs
uoKPTL16V6Jphz972mSGR2gbqMn43Lgn7dz83IeJGz326DzQdjAxvggCsaQopNYJ
T7Q4BJd8L3isxMeFNexFkA==
`protect END_PROTECTED
