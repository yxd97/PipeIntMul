`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlJoL2ULP0qOasZ36z1JhlaQ/EEPpPpQYqh6XcRdSWGyW+1Feye7zmKXWCJOnrTH
OKPbKrE6tCalsPDpipvSdMcc/CnH5oZrGlAVXX8ee/aBaxVayWHHB6yBsiArKbkI
HI3njODDr7HFhVkSIHzpQbCBUQZiEJbUXoGK4pxUpEzLky6W0v1AhDtljB6GOqgp
SrV4wY7RgEhGaxhD9PGbT9fRzlh6hbgckqLtvcfuDL4HzpBtSZ6c9V/OIXA/MFES
aWm4mGascsCMT3oo/Pljdh/5jc5Jue2+j46pHMee7fxEeW1VAfk63GhvwoZABedo
EMzp6xaOsx0LEWI8WtMLxg==
`protect END_PROTECTED
