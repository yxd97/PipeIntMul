`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mc1SR+BoutRqZsTI7tHjk2X1vqWDq5rgHxq3Kpi5GZW4u/nCdq/VQK3o64IX4PX2
ooixGpQJBIaoVJkoPMk3lV387/QOioRlo5ZjhVeakJA/zBwvBfNpzYeMjxSQwz5a
ZNaM5XkUob78MP63uT3fMT1c9m37V1u2/UMxpUCgwdFMGK8EptUmJ7oyerj2pXp1
3rv32+DiH84VkJZjHQdfSlxDSFfmsu6l3SG9AhHMUgkIRmI+CjT/8xb/Z9rgqfEM
hlanrtBTEjautjxSBtnI38CmxfgolpNwk7TiOdPFVYOxUxGrJr5n7hMNDQxfQEI7
sKlbMa2+17xEBKsJ2v//H+v+LG0N9wrTJQX6XrPVzAR5Gf59AhnffolF1mVsMiAI
03THXgi3VZPaWclZUqtjZkq+NAnkT8Wzi1zrBprQx4S2GX9jMbmEuOc8UbNJYADO
OjUf3tQA2ZlDdU4KeYrkHy66gDNE3FmVxvQ8BqoKJOkHAH1w7gNWLjYOyPD9jv0V
upZ6q4cMox1Kpp/dh7SnRB6OMZxisUZ5BsofJYLmSWN/GUyr7LBqISu+1TmYEmnS
veBIchqy9RjD5vazoMjfV/R+N6RJfYhLx2feCEOLn2s7GZZvkMVtjEWP++QrvV7/
Kkq/4qrgXJhC5s905bOz2AFg63BUJOfz5OIl0SPl9uvankr+coYZHhl7C3y4qpcB
ib77Dp45yBxHw0INSwPfJBNAVrJBeUp4pc/i9wP1k+9jseq2tA4AvHuUG791UhRb
1VTwy2DHGRt+1Z6JRG+zY8sRzF3gbHNtrkNCIV1lBskWxgAVctseAo/40EUZpB5t
gKxcP/iyk5a6WiuCnU1+k60B4ZdN9l+WdRZowGXz3YWAnqmcNUS3U5qbgsl1ls9G
DHq4KlA9LI3ViGkrS/OTJu1QAliFkPncI5pVHaFuBwQQF7qGq7CfgimQbC7arLpU
aaZO52yO2drNnmy47ItRQXo8GbbXr2PuL60wDHOo2kaHyyVUb1OoM6610/cgxb1r
4bYv8EBfqSvzrpSeP1h5u1kRyjFot/bI5LWGI9aO2i4vHQzpizvyfIksOvQWB4mO
2f/Ex6XW9ezx8W8naXDaXf1WZd1oUmS3PkxcBDKWMRNwjbSG9QYK59TYxD5r1XFs
UZwdIRFRchGobCQ7rSohvjx6SI6EQSuZAPh7c84KOrx/O7ZYl31TLjPHmF92y6h/
ZApJOMI1r1uLansQLd/84jD8+K/uH+5XWkDALq+Wm6hNvLWrFex5AH16f9+QF6JX
w6LaNW2xe/JlTDBDorOgzSIEw/3f3pWm9ZdsXHM+nEFcaopvgfx33x+sq7vuJ935
w3fW2wswQmZouu97Qa6z6IyEDL+AKROBj3jmh65zxHtduDKZyer0kuccOm0b68rX
pXCbTbQK3g7C3RcD5graTI6B9OW9HQ+v0oCZEgL+Y0CxGgbYr56ynKElF7AHJ+5U
fraR1EiZewjmF/RF+8UUt/wwhpPetBRSpsIqMt49SjylYdSAr+4pc0E+vxCiAlQM
090RUzqSzEGUq52FRxygoYNYNT3VV0ecASRdr3uzi/02GlR+4MJn/S27pEpmln0u
Q2fow7boFtuwhdupwsmUfiWp05Z2+GnoBLmvIvmm2vm66OK8PDqtB18CIuB0AQ2s
C8CBweuC5wIK7H68FiMoQnQjHK4Rz3hz961XK3QSYH2Md+utLsnwGHaj/Ft6GXws
KXtPkCpZWyWE94Xv932E9dxYTPJ/nTj9mCD3is+DBOyQqiTnhv8Yt9lEOs7cbLDL
zHqOeIUVjCvR/Bf8iFT9YF4JKWa1/ipgv8NP6awlarTjgRQI7l8RT3XlB56T/12L
SM/Z+BPBrD2R22KVjo/QfZ8/+AdMSIkHRYuP+1DF129MrES39Zsahjl4i3iV2jYd
yTYYIGybhFEDG9WFI8QbnF13CS1KHttVACPpprtfXzpdgemJD+6xNpzVm2mS82CB
y+P/XH7g/9kv2EP6knHB2zU0nsxm9ibjnITlkfTJZwL6cmYrCR4cCiomvdR9uUM+
Zfi/IiZTK1P63XaGdgZFHe+3cebGm22WIgmv0VFvWrZ2oewRWXC0aylHv2iofOZR
wwSx6L+pYH3wPWKF/vgX4qiBWl8+vbNvGjKTYSTtlabT5RFjZCMbS6qPyT2ylw7K
V8kSmCFyBvncNz9o9+MprZt7oHKrs42z7vdC+je99+Rb93SE4KYqiJchnTmmtQwO
FGUnjHH7LX8mQA04pM4NiNWaV9ClndvxdsnwNWoKWAA7bwgW5IdH/fOlOJ2beVb1
PKq1nzukn2S6h0XkJAOeLMrJFfcDfXW7fJNQojydmDdEbloKWhnPdbvWoOXau7dn
5pvwNPpjELZiPWmFMmXbPt8yLzi55PSVdwaTPv9jJxLy2S2G8A9RyLuPh8vvMNIq
Gqq/zhOe60LuLchhbHp+aOQqrmqcMuLnvySH0pZMsUxPB4XiknAlOFRE1Gn0lxsE
crMX3PSfj/BirKEPxHE4uKdjKG8hpBwHmJ/g00JFEsqdiF4n3GxwnlZMvZnSdxqv
mxwF7UsIm0+oQzwieHYXLCo+OWl9by77t3dYQ0DygC1XJ6Nt5u7ZWWdGlRd+KfvB
u0+YYCQtfsbesNXthWL3S/B/+33NCXzwHvw0wi14M6wwkAglvmfmoURoeO6SZynk
MQKo35lWDhEl6q5x2rSf0RCLRc+XrvbhXXF0WvFA53/LtiFK/HoOHBgZWoC9kqOQ
h3mdojzraibobWrmGMzUS+SG9CulPgIpErgHhmqziEZ4pOm0UpXxG8zCjY3EJWuX
a6q0uEl0NFBlJu5QPYw9ijaW363e7WeVrHWCoeA5Ek8NqFjDjbYQu3viYvFW7RXk
YRVnAEuqNhKEwNT0t/7WK0e2vcZJcNyAXkGEioiikuWSlHg5HuBsAH8fCgi4tFjy
tNosZMMvU2bMdHna7NQSeO3UoMSiUJGB3iA/6Zs5ary44icbk/Zia4zGQVFf91D9
SAUgun4eLQGONjH7h88cjrfJ6npOdUOGrM+9pI0MwYfm7KA9Qqb4dDjQq3jpna0h
kTH/SaUfsuFma0S6QPvgwNn6Kx4R4JTn0ksWDlacdX/WlTww9c67oR/egw8mzUud
/ljArpGzKyWZKsIbYZ6wZ0E86TrbDRZABehbBwWTuCmTLnhiVH6/UAQnk0pj0gmz
7TnWS5PERgyT/9QSVbEYZ22g1gI/duj5Tu8qyMsdHPoa8YGgYkKJ60eaR+KN6DDS
XniC0VwfhnBRgQkP2dX2NqrdpP/l4xbb7jt6hKmOi6hmPQXJ1pQNABBpQTmGMnYn
ZD83ps8gcAXJtat4MpZ7UJHknJR+SPDYepdj6WHi3HK05XQS61WibOyeGMiqRjFu
EUeg+A/3QL5FeuL7WDtd6HUTtR9kzU7eBnYYJgRZ7NP22BTZsU/4fZI8L6oK5o4t
r9Cqodd+MH+3wCp/NvP+nAfyl13ozPQTGCObg194rml1SkWRUiKCdk59VTlRD38V
zFKJfh74N7/K0GpBH8qMHyZhIODR712uT8wB80J2sM6yAm8BqSgU3Z/DI/D1LJEX
UphBLFbVGw9LIuk8D14/x9AvZXtvwIR7oTvlYzQpNpAWBkZAGw+xDAKtwJ41HEns
MxmR3zaj2apmQ3TO12wbToKYxg+RRbST3Q/X8PWKKkTEyuKyi7LQob0PW9iNHEuC
bjPC6VLdWeaBMaxo73q0rDyPMfqFyMHSDASlzfmoC7tSNbrEU7kFIVY5XGrvZsyr
0weWLVeytFuzQc6oTHXfqSH/Sz2dwyQAFhy6AP2mN9zHkyhwm3Txi/ivo0do3inW
lCxFnOPy7H4uotCE/7/P8lK1yRoecPqb9DvWTW2SJ1VUyGx+pt7Jmp+iiPn8N8Zn
+Hc7OR10CErmR+/I5U8WJifVqEMwSvSqlTeVD6NsUkmZgxsqu9wCUuS1EfvBxJY/
c6P+6/QyIWlgg1gti/q67yjR/sEcowTUmrqhIitaVg+XboJYAz5Rd6GA+PgRdQwK
O127QBa0CELp+Vq19SuDgW/0bpOCJ9hUywv2vCNjWI43P4p8wNlhpYVwnaaC/wsL
D/ATg31EJs59y1jGHup/yjYOvAjsE4x2Rh3BWYZbMR6fp6WCqN4IXDDDKk2oKpKw
hzXY8SC2Gm6mVKyYVhyckt/TrzPsLwAQr9gQ6Cpnd0p+HJZ8H+vYhw21HWVcQgot
t67UtYsb3BPIQnT6AJ8nCsK7REozQV0QKYNohUHlXeiSplIQFl2/4/aln5V3e0TV
0s83v5JTUMg0xW1PBdxyZElplEWDgaBppc16EGpVuLHVcLmsuIxCt5srRdzNHbfl
UF1lbPIWe7ilJr6af94Io4Rhd7zDmR73c0gXP8N/GCPQPA7tVSg4RfXChQElyiyR
7RyPV/d8CIaIEPj+ysSDmslW3e4x/w8uLipgdejoCBaLUt8EEmb+j2eig8JK5uyF
0rcUZZA7v202+7tRHsk698u3HQIGwiOF9vzo0Ob6WLB6VyDGqz09GCDVGory+CXL
iobORMoU9mzjM4VPaLg8JV4EiX2OqVPYFpVJjIRPl1C4sGav5O1ylBGtlPaUwinA
k8z5/aq76oCg1zHTc9OyWwWLNjqpnGFJ9fgkt64PIExhqByTQIHyZ4QNoIF71Tbe
lUg+lMwcqeuYTm54gF/lQbtvEAS+djFeQRBkWjQj9GEELACktxzPr0MPrG5vh4sT
cg/f1cTGtqMlU7KbnCa9xpBhVY2kKZgWF6NrqumEoz2nlm17KzYDL5ViDIsqyL04
Bb247Pv+fmDycot2o1MMvCPM5OVWVEge/zdthLTpbyyyPauHxDBoEDqidOLzW23u
jqN23x0Fcjldmms7T94EGdg6qnr/gN90AbeUe1Kso6upX5Gcl0BQrHxh6mtOQMh4
FrFhxBLstotQXBDPSn8P/JBHSsGXUklnwdHDL054WaQCmx3qadikVgU+ala7nwhG
2CSAqABv+bvt0Qjl3fwossTGi2IyK+bLzt3QLMWDrG7tu0krtxtbOav9f1gSYzL8
OwD4BJ0Dsz0NW7+V5aOLDl1zz2EtQvgjytwODs/yY8g7e0wIgBi/dcYa0DLtvFeG
MxBIDTmpqCJKgQ68Znje0x6pqbnr2KcLUylFjghKlXNZkd6VfH1Gcn1Ojei5XEuy
5CvSUWuQm3A4djVvIsZbiwsJDXIgwtH1OklWsHWtnpZyaKW4v7U86TpFjxeyrG7t
NkmWgP7+bsu7L5aKNCmHyrrgpaDYwcTZkJiWEg3RvqBoOhcs4ryJq2rqPaxUyBx/
eDyRKaJ43VlG3cfsFg6ZgmITHsS9uUf94sdd9MRcGbp1hdyet81BfXCFw4JV+HOz
+i6sGhlo9KnNPlNenQYEQOsW1vcRgcsf65zuglNNJGGQ8bxi4/vRO94Urw1IjJru
7SBgrCbyFVlboC5Qq6y2cH22ol7sepJV2IEBvoCbRGChTpHIE1HzJ1HFMlBZsbJO
xqi4x2zprsNsMUWv6qgWBa0NC1KmA1WXKr+N1j8N7sQmtEwaVMVNMqN5d9FFyG5e
B5VqxCH2fgtw4T8Qzf/g0JAXMcOxiG9LHogPuE97O4108Lzp1kQWX8VvUKgD10pQ
eLJFRVdDS4eLJFZxDkJCfV9K4IbbjVPpConaF6WAYgUlW1h69eOOYsp7IhX1t30h
zHz5IkyGnq+B+KVJpqqtM0qvs1/gs2SnEppZuu4/CIjn4AqRXYKPL4ChITw+Z+Qr
vQ59VFgdCxZxhPdy0oxazQ9eY/3mdho0atpzmlF4Vaf1mn33HN1rUeAh6we6OBC0
yhnuvRqiY/2NYdldDB9Eyu3ye9PCesNVEn/otEMPh1l6TX/rNgkjI+K3XU8251PU
B7z4AVU/k1oZTZnj7TsRzvrsYY8eYY4sPJxXEuEbzmaR2Iblmh98ua/cAyMg8Fz7
vyRqcfPNNE9NsK5BeIOdL7iQD/x52hthJvZ8rIb9728vt+/+ilWoAzp5cebtcmqM
6T4H2mdF9PTDSQE1/Xv7h+I1+OoAavzpMiqcQxSy/9Sf7nZWVXjf9DfdoSQ4UYYR
dhDTQHpBbeIgalavAW9hRsDOlrZI8ZRgvG2UoZgfuCYSgJIbHm3XyFXfTW8a9wUL
t71TP+GP3no+oPpmuDEqW0aSetRj8kGR+F14LGtw1lNGb8egteKCFff5o8cPNh37
ZHiipaOqTd01gxEtsLkFHEa2TKXbC3k1ryyJPv8CrqUcRUT7v2EDZaiHf+Y23Zvn
k272zm1vwR79hJPeVLXz18FSnRgmcgETJhJgYsKGuF1WIt5y8rhlENcTw52veDvD
eqfEADgRxtYaT8r/4ht92Sf2TSNr0TXXvfdhmuFtbeHi+3CV4vHHv3zVFyeYNIsm
HH1JgZtMwye7iMszU78Ltg9z6C3tIcfhqwknYT9JrcdoszhHTe/XrhOhn+BbXQuC
v25/Xll9J+ohh3pDGLXRxUyiK2kkmylZRMl9iU/itFw6iGL97MoVnbvPl9xvZrkw
iMt646Ov9dAMwZ+Y7ZQD+OZKNb3cxiqKz9quwcJpqnpU1/HkHUtkMVF/gQmAu0AG
cnZiW1rdwOD0hM6hCAB/WkB2Dj5ayIS8m3BDdNKn0ypevohNB+tjuFvtXemgUDUw
gUcK//CwW8ipU2vJRWDKs/lkP9ZA393hXDr2OhVJ53dFoYxq2GCJqGgTFxqCtlIa
/IFhV51BrwVn4FPwaZrq3jxUU9lbMMnFe8YvP50xBiNQrj6m1xa/L0Psg3JWU379
alFWy4+6JpvwBchP25X6oBFUkAMBiSDf9aPeduzQzghDOHvjNMx+sy7qRZLr4A2r
AvN7juatQQRfRvBvwyR/dT7N680glmZeuBjmoQYSQ177f4WLVstiyrT/hH1Ke7oA
bX0D3iZ+DErfkBm4lSX1l6C4iUpr9i/Hob4PIINglvzVa/IDZjqob7Hkcz4PmeD8
0MWJ6mEMNrd237Gp0CoIv4nH86YegHydIYk9cJK8XagSMQ+mktNAmzt2y4SNFujt
85Wa/VfPoDhRE3/joxgHRkRaf1pGhKzErvaEiv4FywoKGIb78GYxwWRLjX5nWWMv
rDTFe0phKRHAvEwISZCYQLCfE+pGM7pCt9DfSem0MJndHdnOwn8fh/y1OlLgvzxA
jNKru+JMhBEjIkJAQjuu/lUHCq7OUxT3wX4RHSOqLib55OzKUTlUd7YZvTyB+DLW
/KhsiO4k0vhbrpM2RrNWkLUKUct/X4jYYZjO5WVuTsltVzDZWw/E2/75mfkCdQ1+
TWWGM57887zCykQz0G66PFLBl9A5tAfQBfXsesIqCviN2pcr+joPP7N/yqQL3m5y
qQJDkshP2TXNHPW6cCVuR75ZMKD/8Rw5fMVP8GK/NNV81GznxgAEoFjVNmo/K3dw
Nt6M6nDOlo1Lfz8pjo58fOaViO6DbACeTiH7f4oBOUo7ZgpAGNW566Z4zO/QGWLX
2MYHEjzZyj9pfdco/sQvnS/rSn61rKF2xbnecJbUu11w35+RTaNRd9is92THaxrq
YZcUFmiMKe5U2hZ1muzPkjysVena9dKFabTe+vVjqQGPQGOu6GnTM5SFRBgUD06f
UZbBo9ZtV/zoeoPWwGbSTYZp2scjLRfmVkknkAUChpMrqZ4AQRP3dBbpCKQGR/g8
x6RjFnrd32gxSyAwnhvsaWY6E/1VPWtpfEm0Qtg5BZvYXRj5Yt2uXfZjPNLvqQlt
0QkyYtdOmUlE2n7jblOK4zIKKdW52R15ooW5yN4BnOVmmprrNlS49Tqtf7x/mX6P
4P3Xoq1zo7bhvjX6w4j/tVqFgxviP1m1bwg7hyiJMjs48FfjPSlms8H/sgoZgqDT
hNCa5051wWmCFxi43AM9/Kw+QXzmeCbz6pEWYwDDmLs4IeSfTo2P1NPqbHja6jW2
4gWLPjc5WysTkgoezyA9wIDE1FgWYFpJHm8WYTMJNmfbAmvXjUPu/V8c7TQz94K1
Q6upWEgkvYMacO9ADzhbZdTKKYydqk2hCEsVdMYVmjBbJdj5b7jABRTws8IusEi/
S9lrc+78FRGrCn0IqTgmk6sf9KixfglRrehvpqTR5QzSj2N1MoqMkEZichRxePIX
y78NP6cNM1vGBvEw35/myH7IdSYjUyyuj9YX9YW7R3gd76hVm6QFrZnMVfhmWcPw
kwFR9qNmsuscPVTfAVrvqJQ+eVyfSiE27WIv1bGTO/8yDncPzo6youBCg5eYk4Ur
Tedc4rq7tXuvFO2tOFZj80ksjZAaK+P7t1TuQCUmWPB+aJFEf92cT4PhYaz+BOAK
9AR39WVXU7PqoVo/PzyKjsFXAOW8p5HjnYOM/cJxYUJ09xQgZXqO+Eyf5rioNssK
2vn4kYpxgWd8qV4hGkqcxlbYlw9uQqFB9V+9DxNFHdON5OHLK4mNH/Z0iHTBEr/X
yr47jzSQI+LZu6gpI4vJv8qhCzD68+o5Rwn0+oDvZ9YbM4Ry7L+K9i3+W+Cm4VQx
FpAWUbe9mJ+6JVQa7ErY8uWevt3F/om/q0rY3Q1gqHRRHv8A/MJkctGSLSf/3wNA
e5HXPiZXAuNiVp8sr6vTeo2Ntoe4sXpr1HRfze6l5AAJ6kdxBFwLvyf6j1qm7N+R
G6PZlQ9xTc4jH6l4Yvhblb4hHaDcHkrMJDS6h3Vd2gwRkyNpFuEF+36cXzr376ZO
b8nusC3mrBSktmHq5887OcvDWJln3JfwVduo1axh5nYWM2qOJVwe5lqOx/ga0Phd
qM73NE7C1cX6dCXVO/bphsKY64FVfRwFiaM1zfx5lvjdcCIx3jgm8W1IZrVCagRZ
0r1LuZJ/Teg1Phw5bOYMdI2nCPaeADx5QDPbqXVzsZBHOA3FjQOPva+lheLx1Ykr
4LQbTXR4WoUNd9jGIdXzl5M2LEURoVbcOKKXCYwy5Ua2ZQ0sxrABlSbrbnuqfMgX
uC7bHuyjvcQB3TfdrqPaQ6GvrdB/n1Xy7K0HWVFU02vSwlmfWxubgMDiOlqSUmkP
4EJkRYdQXCKsRR/v6AxuxV4Exiu0pUGfzuG0/ote2n8/Ry8EuDrbeT+xk2qtTCO9
tN50vSYdlGPiNVSOAochk5LKhR45r15uGUgdXi6nlHUfpF6jUvWwK1TLFKxivRFe
W0VT9vZjwC/JL2p6FmwwvZ8rL/g0ZKMBLKy7E+ynSnRa4CXyxDYhjQu9eGO3jmED
h2oAzfEveTXlYdCo+/j0r4jTi07EHZKkD/3lky3HKVQWsxhsmxCSyOc3eheHeIaR
ziLMsnKwlHBNT40xm4SPbHK1DgaqvStD/ABGYoswO9Wa1ek4hSRJekDZw5qth0PD
QAwZ/4wQGpEnIQTW1QzQyBQZTQT30PkEzErq69EtyIBJCM40P7TtuodC5s0hTfsP
GPWMKYojlSYmuN8pEVcF8gywrUK+CGbG3eP1RfhhzAcgfISyMd6HXIpXBEE7xHSZ
PFS94knfkzPQzPqGe1XUg/OmmiVGK3cC996BSQWAqOAD1e7bHxrwQ8fWoKNSWnCO
B4QgdZFFc7ONjb5oNRKEO98LwJzx59ZJ2FMN6g7OaZGueOtrURqGJJt9cET9tL25
ZbznEOdxSTp4ELDSNC0Y7uV2gCCzx7wwTS+0jblaRlblygAzHSINg8pnpI8E2Fy4
ENfjYHr7MPKsPP9CcxHtwtMuDwzqN5dDFtRzJxJRw8dZLBSmZdjKY3sSS+LdvLPw
2Pt3uyj8KbITf/N2LuNUOpNHlEPPiklMWYy82hnbq0rpzf9jPOPl63IyZVmwWDsh
wOndsteDhsRS/cK/EVJRWtUzjntXfdOculDhYWjIvXmCeL49PNKpTS1rNXG0tYp6
GD7A5hkGSKeUnViAO9ESr4hWQ7Io1E2wLchLgKHOryvyM8bp9sO98zR9dwDkYjKX
KCm+Rq4kP9NWOM2Mr/AKZlhjXmG4fdb6c/tX+A5rEIAnlukptuXLEeAIvItjZ05i
/7V5Zi4MKbeLrkkHp6sFBtYa956CSRRUWmUgORE/9kQc6X8UiZcdtJ2ZjNrWK1DB
lspRLoKzS7Eq49g9Ftf/R6LQCBnSeqr7pwkUkLcNZVCmtComexlIu0J+Um5wTXjW
0souJlbMxSIUAG0hdTxKmneeK4qfG4D9R8NBTlKSZdA1G03GYioD2NjRtd8jUojD
6PndSoPVRFZcHXHWT2LJ0p6lO8hmskKCxrDC5AyYLpz1uBnjstuXkY5ch3uRaAGT
TMHGtMBK/jKXfmHmhvTcyAzKlfgkGKD5u2ojPPeAldRoNdXQgsZMlgjONj54sE3L
KtCONZLAc7Lt417UZdQjwuPZzFum8JvIx+z9HTIifBqtIeuJKbIRjKjqdZCmaA2Q
Wpop23+Sk304JyTAeh1niCi59DM4i88bwpbQpJSyVsK8L0VCws/qLkBT+hGWptkN
79QKVobfz8JxNufKH+BtHpdDRUUTVD9hp3xVnc+Gy1+VXEyC2Wmj8My8Va0Y/SOR
RvYVFoQZP2iRzoc6akKS0uWfqlsJxSMWtJXuv7qTMOP2NBUqcGl/vxGqLDbbhzT6
qwl5l9gqhJ+12FgFwX6oaIFQISERmFguSnnDAiP1IFJuhYyW0G4HqcwhIoJYTmD7
X7Fdz5rHynv9bDgs9e6IXsKFaky49RvyoH4ThUQpZnWmQsVCKPEKoUcrSua6v3Ih
lJPnsjpuThM5U+gXf9uWKtfXE/tTnxEC2zevKt5YXAyLVTylOCe7c+0mqZIc9dFS
vKOMflrhM3Rl48CABIcWmyCkdZoCQCOCvsxfv83LZkOZtxFHXH0mwYu0NzBx1yzw
sUYnHwF4dg67BUZ+pzc0SQqj3JrPyplTNUU5GlAhR6Ck92X5bt+Ahm9D4HdeYsXC
iReD25ri7aMJwumZHwJ3CUNE2EfAMBt1invYEwL13bMJ8aHmmUGmy5fmNAGuvdPX
LwNbr6Xo5BOYeEHaS6vtfisSyOWJIenIXlvLiI9mcX6otUY1rLLukQO55zU5M4/0
dwczdyATW0Qpc/DuwV0+Sm8I6y1EJwFDslVzy1ajQ3SPJUOaNjB9u4lM8sYxFzmV
f35NIEvmGfK2rJFMFu8rUPGTlvFqL1TqvqbNofP10cxGGr4MotDQOHYRB+YeqRbe
KCai+lK4cbXNwEUrld5Dbwv4GtVlE2E0emWvDwmv5wFwR3u69wjNHcd5+4lKp5yp
JgflzqwH6bPYBz4ggK3Sdc5k6RmEP76IKAvW2eC5D+cxancuKpyRmo9cLSpa2vT3
ZdTT2yIwPaRK4SWuu5KJVMblVpf3/Qj3tdjcFXxrCqvLkeuB3rZyPmFzpQc+RQPc
aSpeSfsAaPXHpAF6M0LMzHNT2lEb+rqX8biaBgWY3pPJXCY7BowW5BwO0dw73Y5P
HyJm9GZOxXbsKzWypxEiLRYDisW7mI73rxrYTWKZ8UPHI1tGD4dEj+HqaoXDRwxW
+/0JPmOzCDylTYrd1j6bZmhbhKgaFThssj2I9m2pitbWBN8UmtI2RKmTsJUjpOKs
RSGUiAg0hz6Lb8ocCSxhtlmW0T4BJ8ygEUDWjIk2Nt8V7AF/tludqOUjG70MCJ3h
J0/6LAjRhdKHzA97NHDAUIAc7AzzVodKC6Bbh+SzQGJIoODAFgq03HezYAdTDOqK
OiaZ5rIXRBe3mFWZ0G1i0iUd5o7bAMTQBezrfBjdvg/DKgM8pDu/LHnOZMoOFFxn
kfbeVnLAYwo/PcpVdSYEWQjBBMFkpisCTaKu0CUln0ZlzsZxOyAYz3vI8hOylqCu
v0c2EzqOK6PRYA7aHnP264FNZnUGUxojYStyF+freCPnFMLdvVGbWUn3UrNKtL5C
4lSFcsdTfqSmpxSSJPQ5X6ougfDlLasM7AjGqR0CmQApedUa4XDH5cZaYpOtXIzU
5oDluJVI6hwRals0s7pFbZQg2DSvI6xjFKP3tbcNo9vRvUh4ODU8ObfAoBZ4APi2
n/EC+1WwZ1wyPPf90zF084L848oi2xlfRXbWIOsEor6bKxePjESnlBeMQB9SPckQ
LuD+RGcw8meCvQsalNI3wDsdfNk6e/4HUCpTyk+OGAm6oAK4dRGrtFrVRD2DyqOn
w/R+X8v0vdGIsOGHNh08sfru6U6jz2o/Inxoof2+54Fc7k8NIZQd/c0fMb4Q67lh
Bb9w+as3pRjtgwCnjuMbPpjFOb5znvdfb6PtKigIx39N8uoWElTTduSLS6pIF1yu
fRJFsv1WP/P+wm5rRV0bHePxXp0/xvqP0GgPx5XLnBUJ8vnGMaxdzXbdCcTcAEul
2oiueMIRvhTsI4H3I+oZtRBw5MBqrdxpwiR1dtYNMlNNaiqQGrKefysZI3SQhEC1
syPyb7yTRI3pg0omnU9vxXZ9gK6gkYGRMcxhxpQK1mvA0f/ldp5ezk4ua39tQhnW
nZ7KSDBNHhPHaBMujS3DD9U9v9Ci+XdrkSC5FTNAmL+ITMX9vYcBBulmoiSuNuRm
5VKndcj/FRGqigJCtw21+ZO7yj+4yV3AdcY4uEiLkEgABP8Hp184MnQs3eUnHn9F
taxeYmvWxwQvAmnxfdnGTt6T7LXhQHp0Eo3+GL6p4mN68adv9qTC+vpgBvBlub1N
pXc7djI5IfeKamStstom1+4f3Ll0XaXSAoXwiQKVEpA=
`protect END_PROTECTED
