`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCXw9WDjr8akYM6UsgUIJ+xaXppfZ23JA+wHZg5yTiXDHQDrItZXzFjNB83nT1QK
oJOb2zl7iwLnxX/pGMDb1jM31j330n1VBFLpykOL2vTvQJOg1psZ6bViDU973cjC
esFpDrSd3znUZbvmkSsmVCw32G7DBpUu2xEod82s5LBDHI7FV4szKHdrRukNuVJC
Pfe4hFzvZAhGibVjovQbUMDJgQLQryrHtrGvrp7oGIOeBK4bjOvilQ19M5yK5Ynf
KsiT6gHbz6LxeZ1tUfi8bXSPrQPCV8B9C0mkfo+VFciDhLlrgG8hWNcO+X4ZezR3
7gRtmQFxQULlFj+0zlx7q3V6YnBpXtC+EZ38a1fGUJ7CuoBOJvP9LhZ4kedRn4lV
ba7JguZN0ZlnkF5wrxXdtFCJGl3dZDYmpcrI/9DiBt4vc4McYNgz9OZkEQL41rqV
kz+FHfTrLsJcszlstpl5Bm69GEi6fkpkC2m10/tDd//vObtx2L+lcNbQEC8+6a+L
DsaveTWnd2EjSnpS4mqrHe3eBxlefs+jHcM3Q8yPUdJ01LGR2rYjBFa8ZVU0Qs3g
+9UbRQIZxu+bcU02ZKZOVRIHO68C2Rs1qUQe57sZc6Lw7k3J89OYNpUEqwaIMYlZ
LURjMTNWyXR+ZuyqW8jwvEq3To4zt6fGv+0/6KIPrTrBsCf8kAn+1FfJ0UWKq56Z
y5x/4Chhy01pb1GnAHCPPAa5pEufMSS3c+ay3KkOjeFKtP7eJ/EMscJJHdKNBkAP
FzanAZ/y+mvGVotboj+Do6uZvbxlDjHHbPYMIGJ1gdGEUvXPK8An3t0kzKjJRRGt
+SlhvFODAXfuwNJCgDdqecI5gUHCzwjNyBaGbPwqNHcMrJg0WoUJnIFfqfiKJqN7
cWQ6HFp0aUyBlDPSNotDPoPKCYfA9/CIFaN6Dupobij9QuV23PgTR6rGEw5k/+kI
ignAtg8v+TzhBLGLN18Z28XMHPKaMdPZJ+8uGNcHE3or19VPAfT1LpVMQZb9JP/l
axQTyH3TMZbBK+lchSgr7OfaEFkYG5DfJLK4e1liNdu1O/L4/g8I0w4FenY4n79V
geyB7DnAVi+InapTI9sxNSDFanMZEf6bAIltcqpx3tHpTgmVdUvTTWOO6Wm3gQHJ
FPzuO32XlD2yZW/WQZWFLaUATzQar1VEST8K8n4Hc0INt6IW3xMOnHuC2WHo1Cib
8s9uBdaCYRL53Xrb9pyA5gaQgsYCoh49N6SCRUVqzLyHG3Hk+1xQk/ZCQAWns06R
Dpxaq74mOiVB/HBqS8GzrkRSGQfkgbe+M/bAtUcCNv3DXpKQmhkkiJ9+bl5iS+4g
R8AFb/6MVxAbD1sW0pJhnwN6YxdyiSco5rDodqpLXocrk7wVRoToevgMY7j4slTf
loBZOPfSr3RVjvbyl3hc/ORzsD3MAIWfAZ60Hrkpp2+VUI2S4/kOcvJWU8lrfnNy
v+j/m7HqPBTjL3dXfm7n/C34odx0aXRm3994Zig5PYrOmxFznG/SixHI9J2NoYBQ
jR/PVqTwgsVjLPNjMUK0nnyCEmFOO3az7oI9l8VV7CZfB6HRueHw4xbJz9pSAW68
Yx6c8ER7fknjEpmcFWEpbotZ+yH3jThakrXMbWWUmbieWRb789U+13w3a9YY+jwx
6vS7zrSe9OwZOI+Yqq/tHnH5jiVDwWfPgvqkBXDWLNQEcvAbZy9Gm916Hiuv6r3o
XTXK/4O2GLz0P46jcGOoZggd27fqkrppy6pFd6Zrg8p+B5MB0uho/rgdu2FEEBKE
Q6lXGi2nSHoxpk2TTaFxr7kkeSJ74OmebFC9RycJm+D7+BJpFKKdDy3saFSPPBAj
Qu5i59ZFXImivTOi5Ua614Bb1SAq8z3L7DrSJd0rM5YUeAo9ahMQH6gcCafh+buc
AVQhYL1uTtk2m/DGw3D+ThuIyf6vEuMp0xToDh2OuJkhIzsss6UVxV9uBCHEbimC
8FsseztGtqBSE0iJKE/Bn0cRdCz9MshuTJxwzDMni1BZJMtm6GN0piK4jdJ9y6M7
FV7b+iZkCD/Ox5Z11507DXEEpfcTS7DaKCnpB6oztCJuvjfvPbg10ngX6uJE9RjX
u3Vs/uGtrxUWhlfAcyHkclqz0gCUqijZ7BWhnkqV8+gEYv3+8SoQ8zH/NoOofnqm
JQyUb6+JharbK75FBdMmx9f2WsEUdlR/ANMpZHA9T4n1v9OLAQSj6c+rn3tQU6bw
4P3uNbJeP9WwH3iTnrbWTjKnbLj61rahsVLMjdD8iD/LPiF9s62/JTu5xdJYvtmq
aiv8tA+9PLG5xo7xVbgYfOwpzjEOdwDWF/pbxebhbv1leKUJTcvPj+xY534LBwKZ
CqKAOzAlO9FM9h5qipF9yHegxvKRZquxdpL1tT7EsP3dS8nmAcxx7gu0Qsd1yaGR
mAxQahPNlLHxpL9CBzNbOC4+GxLFy8Yc5mQg0Jy/3CEd/fiIcqV9/yuDpZi6uDbM
asXv3uLuUQ3KJ1VlTEgit+tl4hDN+tOmEzyZnMDobejVxC8lzFOD3GX+1fjjqySR
y/Yap4azcbW1ywkpwixlKISuQzfGpF/LWGGV3vPeJLHzPL6nx832fP/JEHhssLIC
hE9b2sd8TCm/6LPgZk0s4KSjf2e2OZ+jU/M05aElQoruzeD3JHT0nlRJ0mXCru+j
GF7jvFxjvNTqI9at14C6pnKyyplqZvmc6QXZBJ+FuJXq8W8n9CTVeHjXuWqugq8C
clOr9LJfiSm0IU/Okl96lEBSwLyLIOInpm5S8RcuRyc=
`protect END_PROTECTED
