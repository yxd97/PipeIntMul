`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kBkJmn7/Q+V/yRXof9FngIbUECxwAV9VTgpxu65CgB+c33+MdjnE5GTaeRTjh+Y
3ICRW6bWTlJvvlhg0UkbBydusFTs/lFFCOME+f27+UPLqKC6Ba5Smrq1DTaB/55y
YzJbYtDHoXJRiuSPsgYddGmBFsG0mwonTxlGMgrh6/QQheWJirfjObtyn+l+TtYl
9fghhVWkAwYO4NFCYu4cV2yLSYbmPMl8IQQOcGL3n4mCzfCtV+s67RUVkHTNpvvL
P7qwnlPCHWgKO1MTM2sGZ1wqtWzlYJNCySfNpRoYKcJOR2lqf18/dseZAEWksQWm
VQZENO+ln05l6cwifw+e57eIR8uMcQc7YGT3ks4sGXbIgnGphYfHnk15bNv+uO2v
cdC/hkbftUXidrGnyQLtWSoY5ns6d1Vz9minT6Mnu2O5uA6NVd2Znf+0afY6LwSK
ZLdp43y4mKGPCwYatTjxDK2vbYUFpJC7vqFnUOiX0XuOYoQ6I22mLf69aCqKiIOF
jovP16zrdGaJLoerxwHWio94nsLMDCQPYSKcphQQsEBQKJWu98ppjTVtXBEkbETO
HdL3tLpa8iL9FK2lEwO8oYQcMzT+ObM06x10hz8kMcEB+uoY3MkMQul00T4xwSaB
MCXjfWFykEyOYmiq7YE83CPwcWww2P97GlySXS9pyjJmL23b4oYoNsX8WCFBKCK4
0fLLQvxa6bxXoTsXiB3+r/Q2sfboSsIy5C+Cz4ZaW/+1XqA32qYO6p6c+dUogN/u
/qsK0XjNtNqhUbL3LMouPsR/v4WnxodAmzKvRMTIFPlO7KE+rq9sOA59ZxBcuKmL
YZDwt5IoQW3jrPlwqLKdCliKwhQqS86mKniBzb6TmC9RxXuYLFEtuzLG+zDPkkKv
s2zppP2XPq4wti7pf22V4EuzMAWSRyFxaCAtxbEpIumVEywuSh8Xt3Noi6XKiHuV
IheLhASdfRR24F2GLrtkDrIOvE/tz0tH3kkZwJkczwbvA81PwaAef9EJsS7CoPO0
PRcT/FtjgFytcdTwYJ0++3XhMt6QsiPKihVF4K/1ESXOUDVzSU0b5KIOtWF1CB86
jUo3urEp1hZXMXqnExCrBLVszxylop5lXs/9sUQcrEK4zy5O4GQFxcfZGfkENDtp
4ytCOy0AsVBirpBfX6CA64auFmLLbJrrE7QVPgPc3JE5T2COHOmBhWPAgFIto0Zj
lgfIkdqbnPNSX3eo2geLBPRfpNxlgrbF6kN6BOdwmaGrue+gITnB2VFQ6qJDISsv
rQgxvAM233Ntve8QkH2tWYhtgDZL9+VZUDP3dxBgp04bvzYS95WZy+C9n3KI8PCp
2r3YfShBULrqvBPPp73eq8R5f5oiVpkGLPWJoOMzqvuAu74aPhU9rAGnVFTASdN6
5ZyK55s+QSgMkzDlU2iV4bmMBzD5lRd76lr56Me3lnFnTXglVkI8VBt59r1NjAL5
ZNEMTpzzlSsd8cBJODlDfaD5GNmEwHvt6Ix2BbnnJ5QRga9TZcCVRDTEzidefSJq
H02oQVKfhLQRVqezTQ8rzg/eMsr3lXK9Ujp5DIX/RbZx1//QJoz+8/9BRhFMvweZ
hUN4cfZk4vKw1cpGERN/YMOMPHEX2qpSiQ0B7c5n2tMqW0CeK5f73JPErCnbv/EX
xnXChcnZ3tMgDo/tsCw/5RgMiEodpOO/Sn4cGJPv1MRi1f0gN9eADE/Q4MWJ15/u
Wwwn//eue32tISLgf+TashPTnRK6Kf9iO53ZTkwu+FRji3jYcigp5FbBBuoNCtW/
GMjVXtXWY2fbyuJKASsYR+QZLdZ6OwKSB7hmO+5PPm8zAeIa4EbNBb/d9lLLd3yk
9jGyliPWlzSsY8Xx63Id2xBR0TOYSe5nu3Yspqg3HGkF7kvpciuCdQMEJXJ/lBtP
ZDd0DeRkoWKM+bo/piap/EjXIrtAra5hxd4TjV5YxmVResYU4QwlNfRmkBkblJKc
9DAjs/IsB04UWATWsPibV9MtEGndsJxb2h5OGvOeS8AbqWys6/fwG3giirdAqKya
Q2nifXe0wAAJPHxHTH1R7hYXlRZL24pEETCrGiltLjsrGbaTIc7nQ5QQZ12b4o9J
j2VhwIh5vAOVVYk6M2Krzf9BM2OnSd6Zg71FoZ6hhu1aE6vf8oOE1cmfNxg2Wfag
YjfMO2kfINv4mg7rSiZX0MvfECeo533LVe9iAiKoceSmGVjLCJNZoSSvgzRmoBKU
Fx1O3YRhazuHepWgKpYr9oWC2OXMXckGMVXDm+hzG/sm1ezofjxq4sI9M/UARs/f
pGGH9ReQ9Cy+pnFe7DQf6uzyO0Hm6jzqYI1yM2VAL74rttedcviZCajXirpSURJ1
PpwSAiLtMuK+VScdUwOA8gsSFAV0HVUfx/+UPAjviFSl+SOtd/pEMLe8fYOyFrOR
2fx0IgLCVMUZOzIVz+3L1kCJAJmhLkX6zkoLIULQkkLWP0lgub1ojaJCsSEJFLXG
m0pvX1wLfyHaG30aUvYi3nHW4NwkVMRJ0sTig9kR7v3ofI2EyadM6zHI5zI67p/t
2XZPyPUmPVU7AhtOduTU94RrsT6pZdjSQxJVdSex+cIBcvJkDmziKx0Doh2kRyAv
T8PX2A/lxlOX9k4aXMHBMFJKbchbDjuOEkI9gX7YUVtH9ADyPsZLdGOl9i7HiyAD
eA4JVpy7OVE+NDeHWI5KyJN7IFghInYFeIDPai0T5rjZMV/o6koBQW9E2BoVkGH8
xE099NRe6HK/MhiVXhUsbsShG8cBR+318yQj/TRJP7BQgkUcI8oRElZ5eI1UDDSr
Oe0f4ARGmAPLO2jD33P9FIdQYxUwu/7xluvkx9DMmvbG4/1ZBg6SbALbll2QQCi2
kuHS0peAYazY00NSkzCNudrZDieAyVuMxMc0t/nCVtnWwKsL7VPwC3DywuD/IGWO
IaCAe3qqS+FOOfH6JDDvxoq6lN3uDDWs5NyerOV76mGqvWr2RZVX6+wo+jIvXN1C
ZyOjrmAMCFYLTDZmn9NdihvOKR9Irh8UkARJ6/jLJRBUm0IxKhlSs6SOYeK2msFY
`protect END_PROTECTED
