`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MY4WF9jHaCpfS2bwA1fD7YfNGhHanA4RiHyAtu3jFyAxOWsgTRp4eeyTr51vnVCR
5nKgLdBswt9GnBJorayE4/8dkGNuclE5bIJYcjPl7zR4FIgdfLCBV8+jsueDZRqo
qJcZYC/44ATRJmnJ2Q1E2Nye73iSNtHDkxmlhHfxxToYMZAGmiY+zxPb9rFaKae+
Q4Lik0jfpz8efMcswIDGx5gLm4qXSj1dAE8AtOTsNRWvv/aCx3gLq8ylXkY102kg
T6DL6diGDKl309MDhFeIZNEgPMgaaG4EaZQMP2VEWjMls6knE6QwkACQzL69xqp5
mFcWeyJH62f+TrQ3ax4DIXpve5xD+tbtteRHMgUJY+Jpc3JeRcUf8G+mMaScw5HB
j5cGrXN4uAssIMxEiF+WAZLtZAQ24gw37NHpTEpjGpz1/ROcs1HW72ptaXGyw3KA
7BFYZbmABHwbuh0RJSiyqHGhBdPB82O7Qy0AD/Qq6QomivT3sqN3vA14nyiUl3P+
`protect END_PROTECTED
