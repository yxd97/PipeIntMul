`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4oHxHDyAwtT2BWWGQlfY8c7kFwCC2Da2E2LnM9u7usMEAvkD+kUNs383ityRjuf
E01Fr48GBfd6anLmzsSka/ly3F2mRgUX9ifK48mUmCSNdPWB0gXXq0FhB+abovRa
G7Pk0zAmeJdJ+8rkUxNaQ12tTpl+KcbGRmtE+VxktwdlMx+aUggh19Y8Djvtug8N
q5JtiN5HJFY+ut4HcFN0/tHuhmS4ALQJviDlXyLUq2ZUrVvXXC3BRmaonRI1v5Kn
i9eHYhrs6iWOAPgJmbL40A==
`protect END_PROTECTED
