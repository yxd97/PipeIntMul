`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+uS/wiLV8rXFYx0ACVD7+8bxpY4YwdZONqwFvFtLCwW6Qs8KMZlgMQKbKQjvCb/T
wTl7OM4GfgiivFKdcHq/FeDZto6gW4iYzItYLOYjGALeJ47sMhZAzfy0ZQrXTZg1
XcXOqe2mLTwTQspMGS7iqsAoGiH9dE85i0pvAYeR+48TUfaNt0aJ5c2oeEeFit1P
gcicZhKugBu8Q33zc/YfCJPIxQDg6Ue6eyiZg7bnNw64yJemqmdTXQ7SJdPVdI7f
CB0vmuOTjrJ+9Nc2r7j4DBD2x/Ustfn+cXnwJbDfqB+0EKFfQtht+efKzwy4bdkH
Cg+POCdtPxMXqY7LgklXWtpfG4iqBD1wmLJQ7S1l24EcPw9L7jtoWXvbqfgNQTP6
`protect END_PROTECTED
