`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PP4LeFqbCKvZASqgOxBz4y4a4f/To3ij0HaB9IeIax/D9QuwriD6TOUNoC88LbvZ
GVcr++dagEs/Uy96UjMaU9lSPRDZbQvmFwonsxNup/IaH7uC+7w90ZGIlDXlg6Zz
TMI0RiEH2lIoXAvSba2I3d+abRN2FfB1p+epskFt/oE7I3fwAJ8UnsveKi8/mF0K
pHT/COGaHb5TA/Y2HoNfRJPNhkkMWGYhi8h2YbPe9hQ6wd/GiRZ292AwV/AT6Nhp
r4fkRFwf5trXl57mySD9L8qvm3i2HeD7u6YO1iQikCpyuo4lxpj261VaO0Ch+aPj
R+ke9PphVIoTnbUKZH+WlT7bAJlizSv0yOJkOX/waUNZmkaIxhnhlaeZl7UhmTKY
EWjQ9hJwM/LRwMFAWUC04o5hquP01CJte0pfle0LhCTAm9rNoroypj+LLHwgmI1j
IPyA9EN5DVWQZQtfHceU2zMKlTVIgmKdqYgV4VXWTQE92N/a+tPhJpWR/v3KIKUK
7Xn4+1/jn6bL2p6NZMHlEBGnJ0R7EUdAWOykvbSowIeoi4/r0P8gbQui+LfJeh3c
x4wLHlTlZvrvmCS45gqacCzxmE6veGrbVh2AhcLt0cQUvlBNvJG/ecSjrG70QarG
ycj0+/o+2hYTfRQbkqTt+THfg9LpoK57VrBcWEJlikcKZk46Src2vhcfraKR/Mer
vv/yKWBkrwpdDKpjk7TjLw/wrqfrn1K2+nha8OVNPlU=
`protect END_PROTECTED
