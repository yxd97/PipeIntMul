`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJJirnlNpuEUvwAs8sln8KOQ1oQl89QLpH1IWks65pb/IsDylPgvDaGXGCswjTmS
mZ7LkKVrB7z32MWDT7GjnqyQv63cYMSg9UGY4vmNSxqDxFe8NVgDKxf6AQJAgGwV
M8PLO2ZhiFONJ5f0AKq/7k/wrlJsbLxQOXi7P0sCqMWSk4g2oU36IohbCM2bcAP2
xtm+5gX7vFAROgHdfeFyhz/fP0LvFjFEPTgbHzwHkb8FS5P12IH9OYlcOF3btK95
0BAmTjrsjEt0N6SpVe2t5XDq4F8kg7Ncrhz2tq5wvyk=
`protect END_PROTECTED
