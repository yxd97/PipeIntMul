`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dcpiec1HqNk5rUkFSM6VAizEdVKVyFlZFVzFn6Nec5TQc0BBI/wjPfzdsO4w917Y
dWg32Nsf9rFHar0aTgonWPBvYpXMryvTFLG9IndIGjOGIriBCbBh0Vvi5X1H/0k4
8EbcgtV5QlAT3uMGtqnaewsdP8SJBVh7LU0ROlzzAlCpGJGdxhJ8272/hPgyxbe1
dOTGxB4KqbfzEX31ZiXjI0mb/TyilWY4nLLJRkbqnJ5fWNqbyEv04vp88P3mVXL9
YLXT9wSqz7p6jorKe8/Xv6CbtSrSsjOa5uVLe8awXHM1JSt+F1s5bDpq2rIDwNl4
wc+WlC54UdeTQYXgHuSEpAbACiQSzQ11kTVAMGLKulsYW9qmjMsHIJoyZiLpAn69
UazdxXFIFrDr/RHJeZLDL6J2LLKREJJAgiZgnyT5qJeEwG5zsJksjH2zU3W3ejwz
/FjR12MFlU+gZ4k7KVcgb3y8/EV/SlHlmkSslrlC9PlMzFfS71XVgvNu1BYsPq/1
mipIkZtuUK2KEwCRRta9d+DvSIcV/ZBnEOnpbP/Tb/wOPvAHXUJ4tcE7hUJiLioR
8p+9enxiN7yAdjLRb2/bHlPu7Wa2Qs55cG2hoi6SLNLjIAVNtZJNjJwetU9wh5iy
Ca898xEVuKMMz4J9x4nmIaOrg7bnc5RQGEx4A8H9eDOdT107QJHOug6ztnclGItY
fn2OA27woQIFTO6qbhKHzwgvylKNwce70cty3Ac5ItDXup1UWyyT4pi49VuGyhRs
amH6IXzfn73QHaZqN9sMVqKEmRhttYPr0sgE2j6/k6K3f526LiQOsdKbMAGOv7hf
1coP1P3BX9Fy37MdDk1/IL/J7OGn3T6XznEY4I4VyGnMtSJMvu6XndR8e7gQb2HW
HzNOS2corbu8nS1eUdwsJZglyLy9HM1mjCwdUmrxj70g2VSFFkLTpkdSRLX3GMqO
gXcEJVNoaAREK3UcWPBGpVq6sCo9/6HpkMcSD+DpqPSAyLB65LOobCY0SThFWlLz
CDLSaV/ope2DAIrke0+u8u76PP+bXObqOetWW5DDzqqvp+jP0cdfU8WemZLCl1M9
Eje06z8l7rtojUzuFcBht1jjZh7EpO57mIXuGQC+4S9rjQ1PeD561xThY4knWkDG
2pIqX0HnoiGId3VJ1qVXcq4Sp9DVzCEKQGSITrfsoGD5hPiMSMJ2qbQNfihUFKBi
LdX1465mPfumk72EU2aoNSqM3fCR8RcPJaFlt+DQckNdusB3jTN6nvE10swwxwFT
UkPHUQ6jH9am6KtHLfbqe6c99XRNq9qmeYMvwX/itvMyumjGRxmHm+7OVCvpz/M+
CCKA9n4FTZwnt3Asd/segfZ5bTPwEJSu+AUgVZJi6f6FJPYWsZVAU94dVx0c5Zz4
ayuBkMstiMk0bSR0xnA6hcy//VDB8BEG4KZBKHXwWT1PXAfKYVyBemVpqBQHuQgH
6t2rjFwkUzb83y6d4WETTsCk/hnIb5CBKCYISBQynOWfeuRec9ztfNKORws2ywH9
a3d53ShaH1od6IHtfVRoYZ38Q8d6rivMMzBHRpmg1QKL/6m9gA+NaD593QhZmdD+
ZqisJCdMx9bmTVbdVnARhQwKWN1XBCS4OSOOnms/fpg5QSzd/18RqTZ3zVQxwF7f
BX0Ta3NZ5G8bPgJAMWHYA6j2Yl32S0NtpZCGDhAi1dKDcIAPKKUqeCFwT/jTnYWA
3Hp7I4wtr6VJBWi5+EVMhnqB0st1MMD4+PK8aGPGgZ3AUPVr2h1XDB5F+um8gPIY
BKC6HvAhuabOlgKhfWe7dbQpUUigVg/SK8RNCGWregaKvN+Qb5E9Gwqtf/xzhLdo
sHI7VytihlFpoTuZmE3TNtpakci519idiF8CO2Jxd0aqSp3k4UXPcWLCqMjP8al8
BvSHLbLdgtEHM+zVjAhH8nKWtEQqyHYhlMPD1Ax+P0My+WKU7lfb0XZDNhX5ihGz
UJw/rLaU6zjDXEBO4pyL8Z8b5wP9a9k8jlsPFpDhcAU4DoT0ADgzltojSArtwGoP
FyNaMJgPSysgLnSIZ+TVjEaIqu0rgAtCUZ5r7O2+oZo/rilHJ/5TFmh8bl1O0iz0
SPeRu66bJzFl1LxBNReuEcPCoamUDbOAMdLVvYD5Bvnu8hTKseUIQMB2cLsfx6WD
omjTEIaa0Fb3Cv913ZqWp5vOgh2osUYuQLbSi1y4Jn9uPLeE+T+jXTRycYJCsB7Y
nm3M9xs9hrcZEqzfBSxIqVTafywSkCO6FWUZ78H0pTOlt1IScmoY6ip/L+5/MoK4
+5WxxcbyeIgzPunUU0jMcLvz9GCZTKVdk6rHhTMXpefovm5TInK0sxopaoiah8Aa
M7csQm49DEbS4uQVj/zgnMwF7rUQ5VVv99yxaz0paGh8tWwD7kVqRlUVZuHvG3zk
ZtE2RXeRCH2oR+wc7aC5pll7mRNM6NDKaJRuG1O/ebZl8lkymodVFOHjUi4wrHcV
rxxv+CGW7ZMCD//2omxUuE9yq8kRHBVcoMnz+BPdmtOunN453GSHATGzLFKPr5WO
EKJksgLD5oKeUsA8JYTV3Z/BWMxTomRJk6W7gJJHZjtJpHEepqswpXbtcM3qeBhw
qeNKV/+oP131Ym85tId3s47GhH4PCDqRzKtHBMQjXfvxVIy4Y8jMS6EYF2VqZ1Vd
hoyJaOaYzJCScFplZv1OyMlT1jdCLtjeHxlNwvC6yfOCQKe/JVjBhksl23mn9w0X
/01wqp5JbTXBcaAeW7i9+k+NaIByn9nrV14MxcdxdSfp/6A1nHcpvvcB6Ypc7pTg
IKiOWL5NcPXqF3uFAjJT9/+RXxzpYjOQT4pHvb4YR+IH3RKIah5EDfRaqEy8EMi6
fjd9e56RCZW69opOwJTZBLqLUqrA2nA1mAYSpPYauII0oZnngt6Bz5vWTCAYoEse
mXWFH98deN8VYXJHdmZ8kWj/LFwJYsW70mV0CDepUhUgw9+Yd1pLh/i0eDNej5Cd
/RRXhoty3T5XcDL3ayo03/VXdriNygvfu73mBOUoxwYZ4aBYoEu+DPAm0yBpjK8+
a3/zcIvjSR2wmx5j+Br1XRvQhLQBNPiPuP6CSyBPnIsuitVRAZdKZAi7kVYjKIWA
2K2/zarK2Scmr7oy+4xKNQNr1ibHOBVAcnlSsFdngSpTDtAxzKSXwC7I1gGXVkfe
sgsaN3hXtUlmgMsaB5TmAhfwTvUl88zrc3mjLXzr0VIrBpnt6DamMI50amn9JigV
yT7vqI8tZKhjd6lEDYvWUiv8UB2deAqi8TreVPeof/S5SThKFxoy27+QQd/7ZRaX
AssCGFlNBlaXjNL9vPHcMsvgXDcZO3LBTPD1bZQcZm7lCOx6+syKe90AG06NAP1J
Kd+q855RidJvZHEsK3WDfawWIVvAef7F7N/RolG9s2fQ0d0Q3xi63M9/0fNsrXtJ
mBnwUjafUmKAgIQ1AtGtlFnVBg4T7exbK1xZjwOkoSb8ukL6rZoHgqSlE7ILoppJ
JiSzofOf7erVCT4HCsq8BL+yC5SQ9YOPntJ+rVqdb/sQKdCSxR85pgI2ZVecM3Ha
0OM4wcG1JB7/+pDHlFoI2xrnaJPjdp7lGBLpwdjH7Pn9VNPbWTlTwn7/bqsX354D
5FxHO2D76F/T/P6yb++neJbLEINEBhVOacFRz6CdhkWIeofYUC8mn0kCUYkE08y/
DknFccrgtTkgW0P24z/tI9tHEaQ2BeBySppuOKe4XSRi+Hl2NEc2HrNRLMLapJ58
CLYQf8QEog3mU9qxuHTVyWbO7JfouZDe5NcCxQOBG3gHtd2ssFo7UOo3F+NEvXTa
lvxycxaHV3yp4OFlpLnp2CQoLDqgVqwPY42FPto0y0mZMfJbeV97zRCpxyV0pa23
BGdpBAGX5EdFTFWqhe/SRCjv1LpCZlbArz2rx1MaPNu47lyuF9IGc3/2Th9VChV5
0XZQoEFKu/2jpIToMxLTyRmeP8Dbxsu98/htdRfJj/nHBNZ1Xqg3rgHjEO4j1Wuo
Q7NrX6gLPT3CKYQ9VzmJPqV9V3Tf49IOxu9kGEHfIgki1/0ULjZwbTdMKF8qXGSK
KLkZn/x9xv/ZpGG6byFhzUaOv4tvks34U6uEgOmG3SjKj7O2yLw+gUuQG/rK7jXl
icRZ8oNPHQYnDaGM4sMQXjvOmjO0oa8aYuIxYa3CsQQ6xTC6IHz6vCVB/QzTNStj
pXCWy6XnQHB5HGHKlyxmitwsQHdIo3f5ibceBIQrOR1S2ha4YbS03SgR2OE6t9i6
Sj84RqHAs/OUTTFVom869GTWqKHlULvJA1nOBMXX3ocjxF1i66W8skPWHsSsJ6Kg
wW1ojfx5o6FfoDkFwiR8sDcWYpAtGmVa20Euu79aIklkOBNNzfJR3NlqrJ1pS+T3
WrWWzF1Z1bP7bAIfKhmiEmFSmNDxgmvjeq5W1YkkSjjHkWmaNhLKBnhTQ9xR4at/
d2n5On/rAJ7IeoE+43PFR3QCWrEummm71EG6cMzoB+nSwFo+KYWuDdkA59mbri4H
/CyxsPIio2DSUR7o+MMT/W6LJYbIYnNIJsZqg5Cj8hUYYtTqBF528trsZRiwDEjI
JkbOaOwCAXgtNZEk9QLupSBSI1X/PNojUVxMY3KtxRYvCerTnFyh8Dk3bQbKGLyV
P1VTFP5R9Pee8HCIU8gtbvmfDEcQWthkUhcUTIx/48Q3YFWW9FAy1oNuoOAHTMjq
HCqR8wbOugGgxTtpQ9emmOFEciq9Cd2sktp9gDrXe87WuXuKgbiaUmgi5wnb5dvt
KnCuMWm0fwxoYhzYjnZicRM7JK4ttvNDZml0kEEeHqWIt41D8z59iQ2bUvb3K/KU
Tda2q1RDDDubWIAeGc4DYY3PPoOfmPQSgljymrP8Z95p+sWKT9YF7/qeuJzXvA+z
1KMHiJRpo795E+rKN5jpFDjvkHN+af3LyC2vysehk8TldVg8gjtl+ag97dsrLV+y
JVKm0jSXpgAPZaFbmMq1mijxxGU9WXEO8oEGPlaYLagTNGWoLP+SLyaj5cSR5aCe
xqJy25rP54DGEdBl2+jFTzFiA6NKDK9qYi9bvdY2j30zxrQVFRT4PoENcW1hBEfp
FLNSEFg9NzS8+cf0C+N7JAXJ2WUWTkzamuTZUtKEefLWOjn67n9FzuATk85PlNio
ari9wpvd6ynNn8Uv5s5Sd3d/jx1jVGyShVw36LMcvB5UOFfxK6MaAdKv5H3fYLkO
3c8vUesoxwuYGASOWDNB1+0ZT9BR5jp2DtDpdGa+4jMoP7ZuEMHLAP/IHNdCAFPU
2n6orT9PegzuaClUNNgU2A40NrdvIUt4T2C93FvNvhTb5kKj9xWbEOsicwaPh19i
YqngC1ULvFeRqcn4COuIhvCg7A9a1Kz/e5KGGY7pLeu8H44Cuat4j2e4C3PTL64r
wocONEiSPxJ9WWhJKWvmtKiRMDusiQ/XXEbimruuqPSyg5kSlL74F1vZ/9+RPy7x
qEn8FY8WXp40KPmiaHbFthrmd0uAeNjfD/0XWILjyELts33ZwiDJZG+nlrmRAuEF
j+Q2X3j62zJ6fSwfTJd89HeE/k+zwsVUXU8jPBRafl2GvarPGE7i7bpvYOiCNcA2
Nrn88CUBQp4CyKhYyTXHbhEIEomJgfaiwWIclQLtuWX6LybZhpGYonWc/pwqferA
i9MpTxXUg56z/SS53dpsnv3CX/AWOeSOZBOt6oZweoObXTgl9kP8UMSolDoxpk/l
TLL63t777wdjGcihDoek8p/7/TDYkcV/YCtFRliN/AsLAqZtstoNBlLIEZ08XoHu
Q3BG5yFm+QvCenLaGOBcjJlSxl7vpadDK562vFfHfeBARfTUhn1NHfimfkw4NAEk
rW1tGpreNpQhM0vu7MsxwKSBJ0gS9jE5y4oKMD9gcZTmZBRQIRvuTj45rd/e+0Gl
wYxZ0HlBJXWvXNa0ko+xfdPEav61LUiXM2QMICncgZcmr31D97r3X+fG4TFb+Z/e
iCicehd5YF2HVB05wG/tsud8lHQuhhjrvWua3iuR221UO/HW9chlcjFGsNqHOjaZ
5MiYrc++jqcKPlkv6ycRxlIn90latclf/AdqYH8cBhLG93/IjdvRxaBBntBWdMiV
Xt7+CIeloXjdRIjzHks6nc63JTom0Y/uJjryimLa02qkbJlrpKo78WhIfFkC3Abd
uaRd4RYe0C2FKBFQ3JZxSYDHBcOm80FZhZUqR14mkBfNp1MfUPc9dV9m2imFteGp
vWp9C1h29vrieNjbi0zlKxw4ZCx7MN5OLerULyGocAT6b26SSiy7EQC39zHrW8y/
PDrrxLzAHEtUP4zZeowwSMBaTd9inLkL49GZvoUZp00UFfWrC5+/TbvVd0RdzyJv
BrVzPWsuz/yuUD7sfV5uDP3fnt41yhpWCXr476nQ/zQvhc1tcfgnM9dJzHYPzy0A
k9tlc7WI8fMkJZpYhwtM3XCBkQr4z2dM07YS23jIbroDr9AcZ12M1XFA0u2lC2a5
Yfswv6rGH5M/Sk7b7xT8964RX1seJRJw6oD4z8GERyn9t0d+/hiKJHqvfRUldEA4
MICAzvH4P7hFSJTMJ4jXTM3CyQYZvI920XZfPQCqqwL2VG5ku1ZmqMLDgVe04HdN
79MbbOy6iw/KEDwfdeEKWgjdhzjlrNIUlRVwywKtMdjMX7NTshuI4gjK9dTGrViT
LLnxnlatbX/kJhQgBeugosk8uwaRjbq/URagqFr80YfkJaR0mBexX2AVa+hfoe55
b8cVKizYllLpYbza5LL/Bv99T3GzY09m5SBCevpRSSPbbLSaoUAerdZSYhguHlIP
XDvqWZ73ZH0P+DPHMhHO4UKqKm90pRi9Rcy6h35NfduJebHc+FxG/CF4j1JoWRMU
BdzlD/CJocimtU64QZl/xEyES8nLkBsYI/TCrizePJ6MMqPMH+5kf5tNod7/OAUe
6IY8/veSAVrJrc9RxejvzRe6VjRu5L9uKWeDDg/D65rJNItYaH8MNTCgzZix32u0
thdJxjpJDBEnb2s76jKQeZ5+M33+qHSCLr96TbHR+hGWkHZXJRMAiW6blv+sk8tD
4revmCpWS2s1NaBGTEs/C2gjW2UsuVA2uO0bB9AwztQRL/dYeBQf84I6zedLY0v8
dWeI6ci0qUIHr7QvMFiJ6UomZY2UfrbXVXgP7mXMe3iW7aeN2MzJ8coPRUYB7vVl
IykjTmdizEoJtxKIwi77eRekiMzUUN7wxl28iN/GnzFLqtT5B7QpCOO9Qi/WhkoD
oOnMkAie6IhkfQpk5NkhPGeyvuIrWnVxHoV36MgRQfjWCFMYI16hD3tSzQ7KV8Q7
a9hrQ+WQ61QP9P2BJ3s9Ijvm/aKi1pKJa6nzPytQe5t6KEalKlFaKjqXjzSX6BlG
1qEyOBi1eJXWjiSQiFoGerZn1N3/T4v2mIn54OiGz0Lgq6jBaW6PS1WOntl+PvP0
by7Sleo2D8MmCllZFvgzpomgnEwvjMuoebWH2sdL0CIzUncnVLn9XcUrx0J00CVu
eDo9ZGZpWwHSqo3d28b0b6AZCBLFDhn9BS0cdRSla5IbUj66a6Qlyq+OA8bVykfS
iTtsZ8rHl1PObH0qNKloFNNrYW4Mj6rQ/J3Ujf80fPRwgbhh9wcrNHMThptdUxkA
m1uwSJZIzdOO9IeYTXJBNHbBMt2+D6Zx/pdsVCruBuEQ5/quW8XLOXIZHN26Zroa
iYBmpDBu0jJHryrxtIbYVYIdGSfnr7TJqGhnMxlEedXg09L1CiOensX0GUS4N4m6
tZe3M/SVIYI/+KTTrbTAH2OerDXD8ustxBiejY98omHEbkLhU4JvA3rpH/Z8HW/9
hensO5i+UfQF7JQBPMA8UE6IlFUUPm6nsFZDe3ct0ZfEebXfKy9IuXqmdKAzbfMa
eTvgobFHUQV3lN9ZJGmAFfIKQd7rqvUzjCAfZep5/4Wfbrm/gqdGIsUWQnpYfyak
1kI1Eyeg4wDv8rPOqVemknA/p8wBtrAG95hGUGLWcZhfXPB+hnHP84/HHqTCcE3z
7OpjQKHSBaD8o1ma3SASPBkJTncSQv02WuqHTO/U+ShErWMLcGaeDU96BQrOEwaC
gs2h5CIhQVfWcAadHwPCLtohL2TUQiAgWze+rVYSkOnmQA072CvbBgApprzGzRqw
0ojAeOHLtOOJ+5o3jq1yq1zLF8K2msYKj75c9vZpzgGJJC5qaJz/knktZ+/RMfk5
yf3FBGBC79SDkOtVqg0Qt1MX6eW27tIHVNNGvmWLl1YZlAauz3IHoYWZKSa0TDlP
ztdUZrIkC6VYXORrZt+jXUp30ct9qNDa3jTgpMYhv+KFHBESNVMcVwN1t4+6m1QL
/xJ1nIjoyH9Ui5HTXpaH2jTxzyHhfcXLmVuiZu2hbahQYYMgMzIOy5HPHKY91oRJ
+cxpMYMq8sc7MabodGFf3iRyMaxs/P6TclvFpndQVUrUKF+LIDFI2HgP3CQ3dPKa
Atnk8oGq61vo/sBMyODWU1MrFK4kaz3vpEXUz50XxZ2Q8wSCzu0Ze7nkC6MjwIdH
Q5vN+b8ZaeBoF9izmj5MCZh2jPsnWuT2JG2eSur3G1IomDvI+U53K3k6U3K3/m0T
9vdnB7IsU0kRkFLu3VQEiTL3BxUz90HmPWG61HrAXSza2xg5atYNxVIc2HAU4zWx
lsj9YczL9xNo/mJTzegPC17aT4O4tZyTeGbI2yqDnLDVJIMArWnxE6aldH5Vb2YG
mqFHW4p8T0fPbKkWY95Ee0liJQnfPcfv7DYIucYDv2kZC4fkVDa3iek8hqUOKUWY
cPQmntou/ZpsiXGTI1zicAiXmaVYN59PIEKfEKoSQBClNUQ3Zyu2QsnIwJOmXSmE
/qNzyA7smAbbb4ndHUlP+AVjlLL4/fFF+7pAVdFepHEuLewWco6fN7QrKrzxqXtb
jelPvLu+UnzVJpLBMu1TvI6kZF6zhyxXk4/SG6/UpBWHVlou+BQNCu3pk6bYGOJg
PGQh+2wnv0APitLemhs+hgP22rnzFGX/R9p32Tq4R8n7ByHXK6z64x/tSDqZpAiv
mA1IpqEfAEEZn5Pwi9wQivvVPIKCDLBjhxRRr7pti0apk2TIyFlFLEBJ35Lb8B1Q
x6S9/9k+cBLD34PGtTx/M1uoysYc7cCzXlIZk6Y4oel6Ouijkslx9chtdUUSP5ve
pLmPW8dpagZqO8fqdNPl6MBHg1F2cppAycgjrK9JXy2FzqB8XNaiVAsn+CultK6X
AouDWBo3LbzcbzCn/lLdNIM21tmWwmAgO+q/rMGS37Hz/bX5a6lRz/M77SZ0ZYZ8
JrqvgCMe5la029ew9cu0niYcUcV1Z8/C4TxPuTlkYOaueRYIriPxBpsq0vCl+DiF
PJscOgIXSjOoCK9LiAEZxEpItac3CNHZSV1yz7uje+S8ezWrha3wty2TC79l2Cuc
0FuHUzdrIkBQcoDDEEIc58bo+8+A8roA8IX9F74xckweYICC2MCIzdAKb4kaGsPs
jovsiNSzP0Tz90KrQY9ZRJnXi+nHyQP54KQF4adLGXWgOke9cyFpkhn8v0wET+ir
4i5015MYZrOX/c48rHa0EqibY0Y3nT8CMmvjzPq0osDbQpBa0VxlO24zG0C+oNLD
FYXjtWxksprKUbxjrqjSnbsS/NrvB3Irj/laqIqLSk8dk5WLWP3mN8HlfhvC7+eD
v8nIV9bWOr6DRn1RmVtTkryckabcwhY48RTaXVCQorqx2Ty8GUK63DzbM+FnI/MH
mVb/gJ4CM/e30zp4tmLx6Mzlp+0l8fvy3YWn/HuQY9Vwm2M4AKQCNNgomK4TkCKt
gj44hHw2IHmQwZKGNEsGRohGW9v9WPNYgLFccmFOEVLNIrU4X11G+5QaBwRQ8SY5
WuoLV6dTaexB7oK94RQ29LoASAfskmO8901isFxj98znNAMka8YzzyfV4utUUZxT
Bx1e1m5M12h6e1gkC0kKvc/+lEH6a7+ywbbbG+7DLaQCKSOPYYFaMUZyO4HcFywr
QVAaz9SS5+JM5QaNyMdlsOHOYADeuWoDmO7a4D/4Z8JUsoGuAqLwczuM3os7IDcc
4ReJ2lnbVqmPyQS9WOy0OdC5hq6HjYk/+x2O346JxbnAGJ0b28OkPs2ls45J3K01
2dcV7oUKRqS3pbiLQedummF3EZjsBCAQILMHQcFgxOZ38beKfk1qoZ2sftNwd+6M
8SnoDh6R/nMfAnWZT+m1ACIhG8gaSX+XEYtzNfnHbv5O5A1Ed6jR14Jv6ccli3lB
UOGf1q/6hGTT1RMLDMmbMYBmpMA/uxqnSS0KW5+CP4kBiA1SsUsIaiQFAvRA2ZsQ
UK1ijYMVP/N+sZfzmSgKNY/8xrk8EdH9ofZ2BWGRNIJ7VJaaiUlYXNxvmFUHiSnb
T1C2VxC6xjscvu9WMZPrCdxf4F9Z7lp9htG/XVMHhr/vYCoK1+ZfXvHylbqSSxvZ
O/T8CSXrwbvxlXi+RGV/92acL2H0nhyOUHxHb9+0cqjEMNKTU6jm2D1uCS4rU+QR
KQ+C8JNHHnwCjpXsJpcQHSMcCM/gM9c+2CAuAPestm3wA8g/nJm7dqhYSXrXRUN4
7VGL4ve/hZgOzU6tK2W+Kubh21b4jECrc72Qs1y7M2BFDbUI0+pWh9ex+M18ol+z
lwWPY3gS2c79DElxohZbndLwsjloeXmPIm4k81LQDA4eoRCAUfgVes9qfZAy6LSx
8GcxMckP4GA8UeMOJqtJvgGdrUWuEgWD9mUA/WmoRRTT1fxrMB9HS3T1xZxnM+RV
tDHLJUre/G008rBoRwJry4UUtvVep2FTqEtpihrpUSq1SZggYLW/CNec+Hwl8Wnk
naFWDlviPRSX3ybf/EqZR1SBnh2mImV1qlq22Uyf6sJVw2Dxca047GPJ5daX0KcV
XbW/lZ4djc/mjcq5vMwNO3p/PSGOVhlwtFU6eixh9JvvrqnzKSekiwvBjsbospp+
s1aDURCOw6nowVdfuLkz09KRQhkofDPKCsaoDfxSemY2kc+23gGzF4ddz1Dx3olz
tsGFksD3RbVsJldiTQD2v0LhlMJ1RbbD6l5oJrR/BkmtqyPnPmBxFkvoMRMLyebq
LvBK6R3msQLl2wLZLqZq1q7c3LGY+JIr2JaXHd4cdEVLHbK9Cb5/qbzJq3/r3Qjv
OPDUTeX6X29YUdJsRreskmlfDeMj0Ydb09DuLmw+GD3Of2gU4mkUcNZrBP/WbDX1
UzldRXtgSMLEAOYjcW4NbBzBMm94j4v8eQUbNT4TMk9qib1wONALDyCUbh+X+nZ4
zRKJQRNybX0zyjeOxFtJBbHwfhLvz4c5+Usb8Rb2ND5nHsA/EpDbrJZCesY/n1Hz
PX3Biw109fGH7VSD4G1QAeKwUZGANo7gTPDTQokNE9QWBrs6IA+1Ruq9BdRIgUa8
SHA1qAV2d3s3IYbcg/nA+SeH5IX8zzeBMSaRl9cRV8nt4M3PW/sdSdVXrzXbAE7J
FPKhn8c4snaOKI9N849t7QDdOp0V+kTjUWb+5dLeOUJ3YmX7zF/cnqXpQXydkv1C
pV7jMfToWzC2QxPoWP6G1Og/X2xR9iisWxAQYb5KmFR8NcO6prqqXO2PTtcUiA/Q
22myPAxWL3/E3xS7K/R2tFJXXGoakWcAL5OnjAExjvDDZTvXNCaeVGVxxrXz+mgD
pe7VevsCbzcCkr4Y/pydxAqPGTyUPgPi5M8uqVHO1Veg+mmPnZRTFaA652pKFo11
fBUk2VOWvamT127+NbW65TBJzye+rTlL1lvfJxU5mGKfN4OvZAC1Adl9HHUyUquO
UBL8JAeAR686mDiBxYrWrp87qelPHJrFXm0Y5LRQWuyV5Dn9+2TIG7kfDNKmIS8k
dmJprHBccv3359z0OdLigb6HhC3PTAzuUqywACsd17BNp818GPEKpq2ED7avAlpt
8S7qKIC8rRf/XZ6tQqPrj/C0/noJcdd4pAZwB8EU5NfBQQ5C0xjD5EndwWt+oXO7
e1zZvcYKOzGdHb3ZFSvWsI0rNEQqnBvxh24EfGGglWmQEuaBD8AaIymgDkJCqU5V
Z161W6+QpQDHL1vDkQuc2MCWYWDoxNkXC94dviXT6GTCkOyTvpGFKRw+VhxnK5St
J3PJTNCeBcznhOqu9HJA4IYdaPihZQePIqlNTjgojYN2f/WQZYJZK7kNYNRhaFoY
130clDDFS+0KLDl4kR8fGl5kaLzyPzBH6M2EzsE/MBKVe0qIzzv94V0ZSmKamrN3
ux3DP2Vyk2YiZfcHGw00PYjTtF2BVg/ukc27B0RMnk/kySzBbATAP3FF3CZCq76z
Q3wZ6AGJHx/ZGCr3CfP2KjF+KU6zG1DM+/iXE2w+O+ylCcBLr64cpa459iGBF9gG
LvX7HP29Mpg+vSwqOjG2raP7Nws9h7BWxlhC12Old+G7+hTsxmZ/30TQTxqZIJf/
ghqIULbE6ma3FCvQtoJa+EhvqjsXVX1Ziq8W6/4AXWxD54DQuCgeeQhiyDt1rgDJ
+vV0GlDUZ3tBrhO5Hen2iUFEZbifNO7KQM6fRPR6lFSZdVbRdHFlsEsFQk8AO2QB
M/Db6PsJ6jcQO/1cqAEKi9pNG+IAs1uj9lVPGoovRe7apEQNmxhbqksBMX8Xj7/p
2u4JlxLmRjRxfsjn8qTtlt1qrNARsavVe/35jVLXgwN0/UXsT+6ayTHSey8NlO4P
ZFGcsf4eNbA/k7ZSlnb5KnBay2CU+4jNm/7Do4LSN1MPUfHOZAcR9iK3LeICg0fG
RAofNMdEgoJIiQOZeS4suUrZk67nNm2tYcwX//YO7ktCHwGDTTtDFmAXxa1v60Xe
zlJDZjZD215mbwYESr6aLABSTPmFROL8XTzTh9vjXnVhHeQeOwyGTIPKtHeh4kbw
YvJb3wCjN3r6lEHg4xbKGyt2e0dd1g62IOl6CX8uxAeUkZOX9yEjJeqKG1NPILFU
88YTiQTypy3ko+dBXhEABByx3OmIsNFvr5diy1wfxDCPOXjEKvU9D8s4gEqThY0z
hAlsdn77VQfAxKQC5JD8iX4j5GK5TT8Q6Zq0rLerZ87DucE0mDDr9DHHVkUOrKrp
TWvupYMg1fGRPMRcMon1rEUme2xS6Wf/WnDo3uiEo9OPmN5r6fZVAhPexByAPK02
DzAPlG/gNABHIIDDGlFIXNAN12IQrWOwLZuLgS3drDRzscXwsqrXNWgt/BKAxGvC
+clfedwjMPkooOw4MARoT3SjsEDbCHWdIKxFuIvxghebjS1+9hdltczYKCoOo9oH
sfSg7smkG2Vznp9M36upvHEjE5tp7bZjbJjKjIFBZi0QnPElyWMkJFUYBU0/sSEU
Gpk1BjkEFWHafTN4N49RG8Oi2GZdaRa8/qqxImDMQNjcvT25lEFjwXL0Iumlu94N
nd2O8jeh4sA5kiQ06rO3ODn13W0SSDDvY5/QuiMiIgyVeQyOSm5hj2LVQcH3ewxT
Mk6ucnt/MU2PnZh/IzuN11cySiDC8sGNdAXNozH3UDLq5zqQMRkiCqwPzRcALySK
HwZhjpe4gkwHkY7H4ttftHGs4Z1EVtLao/1BC+VzAEnZ1GlKrIpKlsnX162tkjp9
mN8ekfwLrUjKupKCZ+VPjY0U+zYor6ZYLeqpSuu7KTaerPg8eJqz9vG9v24TrNcM
c6hftr1DKI3Zl26Q324WTwlJWVvKJCl6Dcg8RVUWqnIl1J0CTs9IssI6BCr0A4jf
+tGNLV1PlXk20T8HdadWilqq/wjDP+xIuQ9ExRKjjMljijmDaq+3fatKje3f4SAo
9HB6SLDv+Vmedy+bSuCsPRr16/f1OJxFS8EddMgqbc0uDk9IKA50DaPeVTyCz0jJ
kcLZnoXftvpXXJNzqR/ESAsDhMbW6o+13Agzs8sptUVdrRn9sGsL54sQ7j8Yzbrz
gitjR1ObL5KOAThcPWxQwVxZVhRC4jvUum2iwoPocHWkdHXrEMQfIaJWchAQP9cL
ANBhXv5tgsg25qEO4Q3tqPH13XL38UwUL5s5B7Yv34S59jbVXmTOIY6yunzmdZA8
21w2BV7aafpsJXNqeV+5UvX18zLPI4YNChh+hVR33XIJizXVNz/AvVXKLHZiUUM0
u3kgMAk/9au/LO1HCUT/YyJ5xXdYl6+vaDgH/Iw0qYjkyiXuOEApyk1zNNxUN6bB
EpviVuvgg8FEFkB5pR21SuMh3wVpMnprIgYv2SyrHAj7glotiJA52kohkMwS3zG/
A5GJUCLyBzS4swpTT9aQb/mlkbNZWNmJLEbC9jx0PLigLeKoyw7ZS/OhzlZ97lyu
Upbk8pxOe9KZXHn6Dq5kF5xyYXTMZex8Qat9IJiTtZvkhT+eQ3T1+H7VyfFy6KJX
B6om3k9P12OrsrrwsZEuACv0SBPe46YTqxCRWukp/xac+INxMDPS8RKUKr140I2H
il8dsVuKLzBQcK3oEj0KP9y/Fq51rkFY6cBVUMa7VBYDiACN6/Sjf9QClH82gTbi
RTDbA6sFOph/pqScMhdFNY17/RZ/K/ol21MpW4LIh8rEHxtTH1g3fY/w8lFAk7ff
jq7bqPjZuEJ/GvVQvtugLNobx1yR0yVpc1p3RkmsXp6p4aXxf2T3z0NV2M9kikLb
lLcDVHp3lBZlFhBOp0CY94Xq7DMv1St33Vw8pjEiEhL519zl08Fu+02SsO9ah9Y/
nibrifOZ5xSxHGH2KQggI3P2bROPRvrbbEdTpowEKcmm5Aw0r2sx6bBlNyg5KVT8
i8pYLdW2oEYol+JPZOBW1d5HziVFxHFu1JGbSm6lIiokG498EEZQuIvnk8yXqV0c
zaOm6jmIis+ef5SeJXzJ0ixFuQg6MRw6yki0juGGthDh9idE+BtGMHvq0Omjs+lf
fHvhSFvkOXWbDErvNg7JvhUWB7Zynv1SmTf1A2bqrHYgSM5bfhHuzRjqnMLakfFu
SPxoZjNCsXtJFyTv7PTEGsTVO8y5uMoiVnAMCDT06fz9+jMJJQDIpbNhSplqkiOz
YTqBg18zLDmzmgdICam8UF9I6gmcvAI55cWNdAixxwgF1J0OORQ1VQq2/DiEwn14
I5Fh+//0u1l9DosE5+UKWWrefVqJ3/bk1QB4sqA7PSdRa2lrY/dC1xlNX2HGMoWt
6P40L0PEYuDcSQZQ/FVSmpsNouzQzTz1Vm6Tfb3i9JyvBmwzeWoW1tvFg5uiU/ci
lO0RzOH4nDWvHZ6XjTfC6PNFTb8pDFM40kRQlkS4kxu5J2v0bcBbQ02DBJcNbNhN
/CDD9auIP+xrdgcvPHjnjOg3dBf1DJdomQfxtdo7pcIn0+aXj/uX4azjp3WTyHia
kqvPGYBPjG3QHSdxP7++FInSkt/H3+JGcheYgTKocWP5/SxCHLqOOMKPIxmOET8Y
n9GvTxUPCvHJvc8Gdj+2+M8CYLTBidHUdc+UPi1pnNO8B9/q7a3cI+BlIDBt/4Fl
splPq4kNgVkXEh3ECOAAq8WSUQRrvegnaK4b22S8j+TH+YZKMx8tzf6ivJUP39sE
F1j0ABgEBirm9uFuadLHO9zJt9iGpPAm8fkquvELWUeWm/mXM1Jk8khl2RDeSMlF
Q4ouSK68zA82sQVfUdhwQIkLEeogyG1OuTDLdODRN2hpG4ZJikQldBeBNH2FKZ7b
xmx8Cf9R6Un0HRpN4QjsrsakvMahP25Ekn/Lk/x77fLq5VE5ObrBYzrd0agAirbQ
c/SQUdRAXXkN4UHweuPxjQf2lMTAkYnlBD1c+vntgMZATtHkETaUzhw3Umms798I
xVDdjdK5SOxgqRaF0TaOQTfFnwoVA0r7TrW1qFPI5Nyx6Mo1+jvC75ksA29x2Ljb
uV9CWC81E67en3lvzq7yt/v1/q9GpY0sxBkmYunWIvypyv5ZWbE5tS/+5UOD0yWw
+4sIXhHfCe8McKUykInqb3pUXvwdPp+Xd0V0HdSsB0uPyMKD8bO12djhDNMqPHpD
AJeRz34x8SWNHJ3HMwp7IFGcLX9vgK38jMngw3Ho3o7QUoIQ9Kwe3JKUHQmKTAxC
hf1ToMomeDdBzZaYBJhTlYzhlq+0Cbefvtwr5l6aYAnIljumObXOG06Q7xfhclkg
wz902IxU7S+9CxzYr3Ar2N0JbDsZwLaXV6myRPFXHE8TmzpExhaam6mR8YsFH7RM
YX4KB1cGX2H2XnxTcaT/pyY+GOgKe+hU7/q1q8JioNoTDXeTAYXsddXMnEi4USh7
YI0kXLbGnd7M4pKEb7VWwChcZcybj30bVvHVYxIwzFQIHmbub/jbaQ+GF7pYD2G8
vHMoZ3d2+u2fZGsLVCtd8HMVaSc8mnSCxMNHEfmTBmCP3uajFbjkc7t1ZTt4Q4s4
OOUKgWMIX5Eu2bfz9mWGMvtapJsknE3yimu38OsJfYQRy1I58nM1bE5ZorlXRIOi
QPrcvxim+FdImxU3zdECnEmqse0b5OFTfEopnJb0xujfV8bBguq82VQ5YKyWcJuH
L6LgJ3Y82gCdP1Imas48ifMo+TlaKgmEki+sEdG36wb8RRoE9TT+TjOhIOSkJwam
7PdwmYQJBbgUe4UnHrV4Ei8yJOBx3rBF9q8gmEmVi6MEIZDut2pKtiDb4fXE5gYN
5O51/dJYf4r5lanh9EI5dZwUiA4b9nX5VY83ZsZihCy/MWQvwy4xeUIhOywX+VlL
ftjgkIYzhaS2vKqkJ0gJJSz4+8HJZOhp6+Dh3T+WSbAEfgrbEyhgGOgVWm52Xxk8
gXVLkUfkAOt48SnGhBnIBJ+sl7EIsjlfQ8tIC6XCMAeFrIW1tYBzoTpEN4bkCaqc
y6m1B8vbRqG1uWUjy/jZ+iSiI/YDo2EOD/+TRwoweceZrK25fTvF+iicz1ogK8SX
nmhlqcCZ/0Dic1fzSB1bYPDsxA3H7INzwx2y33hSpsG6QzEbJ7pXOta1sNfpQgS8
nJuseZw5eUyALLB66HAuOeL6RA9h6kMeyxgRMhehcSbuDtaYVs4KQ6Nid1PG7r3n
TDO9sLdwpKRoRASmSjzgNHPE0GeEqsQq9znDT0Q7g1ol7x0IRFJgh93T5Ypbun4V
/LTh+7mYdEA53h+VtpmtWWJOS0v+gaPb8CLAnjNhPQpeAek4TvU6qWN1iuULTA4T
C27haO8LnevMZM/mabmzmL8PCmZHf9kSJ+frYMgsrOxPTwbMbODlXif9cSfQVjMc
x3Fz2xTuKZR0SBbueiTmMID24xpPGu7S/wFQDzzUP1dTHdFtNaIaO8uVJaBVrgMX
lKG5p154RWsCE7krTNVsnnt+v3iDow5F5YxsdtfVW6e+YRnaNqi7BJOOCs4/zehz
LEJYDNEgZH7aDf4mcW5DnuF4Eu+PBBx3FvfYuWkuneCrYDw9AJetVzUEyj5SZxjf
k7ggaZ3JEiO866BPcsa8tE/OqE6UXFS/Wv8iVtL6bqL/UaTHOQPTYv4CfGIt9mTf
QLecG1RBFTZCqGkC7K5e2z6ZO0vlnraGvYPNmy+YGIv25eBbI5m5tj/mSn7/aMi3
ya8WwoK/cFBdwry4r98VxI/WWCkUgc0weIkmwLUszvdMfhgOSK4EJxqYg++4PBEx
78x6Jvy2kcwMbKK0RyI9qhxJLHhyIVS7aOhE2ab6AJSu67FbGX8uLW70zFwuMUxF
vSXJ/u9l+m+WEzpVrgMYp4mZEkOLqZgbQDCfLBO0vTsnlBfYljvXOJ1XS7n5ct/3
BFfLD8APaeH8p4qLMEWf1qZdb1soM8ggZk+W2Jp9NT0tQ0Se6z3gXxqGz9UTO5QF
Q55daQ9IWk5IYKTb8hza1V8L+TTyEZXgyg0wN3fNNX98UyggEfTusPl806fY70br
Cr+nRg6tRYGM/wT8fqD1gVSAYNmiH5jZDch8rqyWUGFHA5TApDpHL4sHq4Igpqu7
tphoI2b3L3SQ/fRFH+gV8ll2rNT/QmzHHfUOvbLWvn1rTXAKANMOKDcagadhloZT
w9ACvg187qrBL0CW7Bt89jdLYah45Ff+sVrGYHNtFdq4dNleZMNif0LiQsg1xT7m
JVjiguZm+uG6gpQUP+fkjXxJZyY51IUjmPRaAzRYPlxfE/Dixsna1aGZomECsu+/
alsLxDxaoBqyasIELer0tz4WsQvoEcTaZoicNqsmn/MzECT83s/RDAXn7Mggvap7
MQjamboTisxo7LCeG1aQ96bbBbErozXYvYXyfnND/47qVz+PdHAqCm4AygQPjg3E
nQ7yZsQCQvqWUEklbJXQi6NWiojxo2+74tUQW3W68ANFI0OvUsrmHi2NUoZiWM+a
lblgEfRzvceRyjZyYDUBYppuBkS15CcqcCtmXr/GUiqIi07yX6f8ywTj4orLWXXk
WQGoov0dXEVzTrAVGTekldUNEW9oqY7DW962KyCUkksYrChw1/PYCjE1pnYXAl+9
nNj73Z2y5+k4fd6VTKx9NICkDxCZ9lM3esu65qznzkLIWt7GM9tkLnOXVS8aNiJX
vJVQQow77LS3uFr/3fp/05ofn4TEFgW2k4GAa4NQehTfSJpdHo9Ulq6WOCzC7Ata
Fk22X9mlLSTRnbeu8uTB3bPqysRFKeGhbonzJCwk2XnX7icrZAvLdyegcq/v4fyj
Y1qVKIUB/sqTg1r+flaNuUXLqDHo6sO6mCumBzPIpoMFM5PrmvpqggcWz/pTM2bY
q9mngJ5dUV49kehQYQG0xnp7vxYerdmwmGz49MYyp+LU/nCC3OX8VYp/bEx43LBH
PjTYG1REQP8VV8jhDiNqe8o2vymTx/f+H492/Zbghl//uttykftgfaMJQwW+MCLy
Gns90x++hME2Uu3u5JYuzPlB7kKeaeN8Tp2OhquBN24rSrEeYvpbYbDfp9r5nsnj
OEOFvfXrYzs1GcGXApKX2KcaglsTcpxT978IrPQaCtxklBBUoTsL3F+X9BqC23gG
ZoRmT5MiZg92OxDgP27awvOzTt1X2WgumyEvzErDAl0cmLwgtkwIw40hF74yCndg
O5Jhci2/YKya+vE0T6OqpT5bmHuw8JtG6ZXIjaGojtKekRNMyB40Dn2jjHQTDBRD
tz7x/zsbfumwAC3mu/6XCx7jVxe2mC3lqr8gG4dni+bjb7sv+DnjfmlT4qg749mb
cw1CegydyJWo2lCugxXxTIJjX6Pw8NxR1nKBE3HZ3NZEi/n+BeJTz9gnZbS1LfF+
lgFhot3L2eUQl9UR8Q9XXUMO4eW7EbM4xpvfIt2McwmYRaRv+ZwjdhqPoZil0jMu
tJ9UeLOF2kN0Cq8jc0fpLXWU8enAzdB1eYUAHTRVA2GG7EqjaPikC1x30Q9Zghmk
4RK8kLXz9a4v+qiPWC7HjIvqlDkBfXt90vV5kct8BSoTnwKz3xbDsTplMtUwau+I
SAFnuz9w9uD8aHexl4QznhBNN8XkEH5bjHn5NEUY1ysqcdP67Az6baM/q7eCzQv7
vWUS9LbHFoDmFiYc4UXcvgr5mKWqEogosadQto7D3BxteDu7ZAcbWbi/XS0TmeqR
jCLPJ5+qAzQSKKiUOgx27XdldYn+9fOTiZ58HlXCwLZX0RxEu3D3rqjWGqRf/6fF
FKT8qKrV7wgAW/xfC+ttxj1vGKKaNtAf+1DifRtREA81TJCBbHfKy/UkneSPs4AV
fBRFzElNZsL8wYCUxiB4AqsIV5xNQIhVPlrD36G7VUvqITXYaSSC2xgA1QX3Ba7i
LC9kuh99DqBie8zwc3W9CFC80ub5hvj20Txb4jjC81sfToM7oZiInXQ0LQfa/i+U
uUDBSVh50z75WD3Lw87DFvDsMgGr0Ey0lmVLOjTthpwDPRjlbaOnBlzATwSaX/dJ
c9ZA8hSX0VvdGswi3/RhkL0TIAm49B/K4aJV9CjN1gmwSaR/xKyUgYplFDSDTjjf
M1QBC094hGtZnKCKf1Ge9fBpU55R1Euu2sTkyUFfGvdK0qVHKsKbfrza5m7YYoYD
lBjmej4nqZZsUjYubYuqytoOeDkKULMF9vTGh6hj0VxyBEVNd05stG876urFMpFh
+HNgopTXwkLOb3ihN+pZmiwobbj2mq8N6cNAUNDwU4J9Ixf+eLOfxh2UlD6skgXH
d13LURCaElj1c/9D2X8MjyWPa/ABX8iNLSHPlXXnzdnkbXT4u19Nm1mzegAtoxpO
XU198Qfrtv+mK9Tjxwl7H7+b0GiXITsycV8qfNvubAJPi/sjX7H0wpmlyQ/gMpJH
0IDfANuCPF5jCI4mcSaPIRVjs94w5KkHEx5rjyZ/mha3UT0lveKXOMSRk1MjzcII
vMWOcoU6kt9Xq2dBQnyKS+KA3AzGzs/YUd2fUBaxMEDD1a/WvqwIu9cKolVwoXCO
FhLQP2R9b/xCD/oDg9eT1ZPguvdokOf7IRqxWYXHVxYEzEosJyNLVM7xcxUaUMV6
yvJmvHneZK8f50NmSbM4LIXp9Spnj3p9ywXDTCvLUxik1hXODxgvBy1ZuXIKfDs5
ZPh0H5vv4x+1+vqzXsrTGHmlFByke5IEB91bcu0gpxOwJmwBRzD8Usj1u/fAw0An
TJZihpbAzPpcqKmQFx/RPHWYliotLAc1FMrPgnayvS5kOweIr18bh7RaZiE4ZlZ2
vGyNWZ/r4FXrn+1hKZRzSnL2fpOZ4utNUjM91tvBHLRwGQ8EX8IFh85b0DLiG09m
gpPufTE6OT2PWg5lXVbGtYD1Rn5XbOJgYVK+V4a2gfnrl0UC1OnDbQEKJYCoeH9r
neEDdaVrsdVJm2LbKkY37GX6xFo7BdfdVG+ZEH05MJy6dezpNIH1mL2+ElQGdda8
i0x0jk8x818moEazN6FKIsgBGyDrZHac4QIoKDKhtBtMbLSHxDrwew83tlDlzphK
AbsR9ryBCNUWEHuRKuesk3gJbUyYovAURPdkjn2i6SCPrH6VPxta3k/RWhzNs5gS
SMObEMA4NF1Am24gKiY0FhtagNm5E1Lyl/kylKV5UGGiRrUYl0y5QwWWT4uFqCK4
DeNb5Gfl78lCYUXLe9cmqCp8nq8P0/h58ILrnK6ztXhH95guJTd5VNCzcpBc/705
60rsAuk2UId1TVQkdNMIG/58cVcjuPwdbtWrQrm5VrB0Rf7CS24+TIDEgF32awNv
IrINZCPt7SN+vZpcg93CqfUzSPZY9ff89Rn4nml/X3FJm6Hy8d0EK8HSYLW9DIVB
xA1G2sjkENyp0N4qUO6GkImNaUiV7uPzxjAekSj9pq7ToB7Qksw+Rj3DV7y9C2Mt
i+X912O6uUgtSRqpOUJ3KfS0WuLBR3Zh6EVxG7NDBDqAaGiQ+4frSqb8Upzv95vu
EjUVA72926y0zCdczyjgQF6r+0JqtsJCgVi6S+OC525Oq8UyrGpW6cBtXG4HK76m
mwcAYxLwQ2WaAEHCRxcf0SunfVp/ZxkS3akSzS6+VdC3NfXD4Vo3r1yJRlTNuGJ3
bVBPrMh0b+xZ9/SW6QrT7QG79cyzQZ11XbKH4PlntXjoywaXQW9iFbWJUEOnwn+3
+zPTCuczj+quMnpM+fswc4yW/cwd5QjNTXbtwzSaVecq8+YqUExKiINtNVbsth9e
cWUh2livfVFfdejxiW8BZ0CWOOku0K5/Npu4LJUB/lapWWnMS0g5v2auqZHkLz2L
+wF2ANP6RAvHox6EllKreys4S9+iVAABqbbri6bNDCFMY20T2VsvYtzCpD1/o6jc
x8pfNXoF8Yo/ilacuYlgON2WolGHjyX1Xhj3sIe50BQrkTSApR3Zhe1PiPOHk8AA
hQXZa4sbir3gCdMijY/X0+8UeKgZxo8/Q+1QJRacH4h8swycDlElBcWnjZSfj0r6
1okgMCPjLP8oYyVtRicBLrE10M46/5eHz7FKyJszRDaSOgSW6zG68Id6iEXAgaPK
nNPRZazJ66UJ/v4xK9rtj/KWn1tut7+ccapCYKROFX3eMd8HVAKZkTjLPFORxHa5
FUP0e6CDEa9FNJuAqCDZkxmjgVbyzfY5fAAwkPB5FIOCnnDZ6Z7vH5DtAvxLaGxY
Dt9wC5uLEuTv+8P49/QflgUAU/XpDMyLjtA9bZ/HzXtLbwuFkhhBgZVIBzobjK0Q
j6woV/epnwV8kHZkL5CZ2k4iUPbgN+oTKDkT9sHwGpxE2SNYuMlZSXFvfzMiMi4k
jau7N06gl3Rvq0wDHRKVtbLqXW9qJ44W6qaxk1rrBEQclr+er53ZuJnFe7DY32SU
7gWsepbH3nFk2cnxDkx8pWfuUCJrp0OkytqusaNIHn29Mqp6m7vnQXHWGdnKhTD2
ZKZgRLy0EaYj529DvR7vL9MMbz2Crqh8/JBFI3GzwrhrXC4TlljlzBq8om6gZZmf
0sYrglMKyN9f/TRHpBZRc9uthHtf7CSwzE3C6juj5Zo8WB4UguKeO+GXew0ZJcsv
64cVgVjcLyW+qpfZbgJGJXLJVvnrTuIPyNjDaFoOWMrfG3J16+KJR7eWivve4fQo
uAfl5dH4ffXuFn96ORhg8AtzL/HczPrPUA/ByHmc/oba0ykTEWUOSMljibG0AymO
RcDvNxkzyXhcguUcIqxszIuIoZRAw9XKfDjworESgccoyE20ELlQDvdJHNsPBF2T
OhHwQt83fjTpbWecEfmKOxBjwiju7clZRDW966JVNpq7xvhbOQs1mjPy6eH+7ZgC
0bfW4ohzI1idDFKVNd/vUdHA2wRhrrLSuVMpkZ8CPxxfsqZ3kxFhgi11sBOZP46D
gwcMj3TPkMvJ+oZsSaoae7AmzU1yN6X0RJSHtywHe1U0B2E5+Qx5d2YrYiaLAJbk
/EiozHwH6/w0/mH2JoiGc3pATEFX+XnjaVj7D4IXKhrMJSn7AnwSDhWAnE5Ri37z
KgT2hk/6072cvaETgVavDzcjl3WTgE+1RbKDKxZ1KCXp5++Y7CHHmezNs/d/7tg7
jQlvVNdukCkxemtSULGUsu5KFswWQAH5QzCuqPri4bUyWjhyQs2qJ4eLNrvVog64
STNcfOGw3niZG0RsSn/UqVpQnp9ayhfCwCos2OTapxukImuWGDqZ9NkPHewyiV0J
R3UB/LAWst8apGiLCl2pPPT2zKBYQj7fbsrQU34alCaYDiXGwTNLCPARTUwYpZmt
w4EtC00y1XYWVf85l0WhWipsetfHogIUqr0+z1ZX2vYfSPnAfLAwam3tyj1LEGoo
AvV/tHptTiFV6zG0/3p2oY6AKiyk7Oqtnec81/1Extcs4YLhwQauEwXBJMM664Mh
Ujwrx6jseFgnp3m9aD89zDZalNcn1MlmTP8Za/7D+1zGGRE/rOeNEMNcswvfaZQL
E3+oWo2g05TY/JPfUgGd3RSspoAyptSXVfwRxyM95WnQndTqa9AYf/VDxdP+l6VM
/vwdDNMLi7ETV96jaP8wtcLwokh3Z3CaHdFjzuZX7yZmHHhrdBMP9Q8NiJnMGCqT
XMLrWNneWv4G1wWZzebmqc9FNI/v2dxIUOEfAW6plSRI70wjX5lgXzaJyno39LSb
6pnaDFHPaZZSH5B5iUvL5QQioi2AcPZI1eGQQbCnst3YzBllifsTUipVbMO++SVM
uZi/4OnyUyAm11a8wdrerlMUNe06yDyViE0YNNK3CAtnrjebY9bF8af+89gi5Z2K
vvGCnNnBNZWSRNfAFojX+8XM/sy/DFh0iEMN1xo4jOK7XDlmFlCSOkAlcX/fYSsQ
SZU4iJLd/5GOYA4yy1bKJFSCMQc62oq/+7UmkuH/58N4JKJUuOJFsE6tyrjIIuzk
hPQ48Ri7wDqPxQodKamli+/IsW5zk8spa30q+AOgHR7B4acaLRyswEhhD36rOmb/
M0dNe5U7ssOxE3RmNTfcNIYfS8hDw2Se02RQD2SuxeUf7TgUn9U0Lem9Xghc0aBQ
S112STxMuOzQXcMrxqnu7AwaII1dRyZlHTnh2iEtC6BWwi6dcwaYcL6ioVbOkSNc
FR5rR8hR/TfwkPnYYAeEawW8TTDhQejsctlXbLa3is2/3ykXuPYLvxbaqMiOO8W8
gvgqm66gbvFmahg1aa/dtxTIGPGs7GHsB14DKcGr+cf6aPoVw8IBUV1V7d4nOXHN
pW1cpE/SKDVlpGENVRDJOhcwl6ClYY09CkNO0Q/3oJm5lOvFYCQlwhzg1iz85OjA
RgSzVcaCpGpUp9XdQTaqlWXNjhdxFY6tApQMn7D4ICy3BcY2yvyFVNaoRAvEgo4U
X/D/QdVcPKSxNoko9HP834Tp8/3pW94YFvqqBLwmQoF/9rMnyKS3yTKuDkql4fHv
6NVq+r6GbmsVh9Yw2Zy9NIlyK5u+WqSmeuv9fCVtP1Ox9pq7sar0u0v7VA/wzXTq
aiHAfC5uyDvN7bNMTa4KpcwwDknlCgx90U5I5jGJr+EKxXU9WY9uFofepCboRg4y
HSFBo404gUc+/P9o2mjrekV2CdWipVDe55eXwJDgrPbzk/2333F0xAsLiVhOnG9n
QBTr9offhW1ncVnvHOd/0wkV2kbKXYLHuoUhXuVCsZE6mGstAb/Y5xyJ5rLfp3du
63gzOlhV0952PqYq0gl0y9I/kjzNWEVY0GikU/Ba1yPQreV6eGVDfhwPSAqNvCfF
C4EnetvDWM2FETF21olsSpjPfUbMYBrI4o/RspE9xIGmT8CgaS4DTBt5nGOKJYt7
aGkmbChlwbUemYSSXMuSspJ3ZpfTotyu4Zj2G+SM4uU=
`protect END_PROTECTED
