`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5cNCZFmd0pTPzVL2xR1o2LHLDUedS7ypbGKKzRa/3i2P0t7XFq9Vv8CZEoG6oGCi
sX7v5U+wNOI6IRDewdEuWG5reOw6csgWih5ZG+qG1QbAf9P5rjz/AoO1uqopGGZV
ioB1pq8ZzLI8Wj6evtQjXCQpD5jUaAO+QgUkgx1s/CbrxUxpPDppALU46j8Omefm
vfIklXscxt8a7xOEkn6Cga0XWCGmJO/w04UJ3UNvAoZHxkz19YtLSCaSpCPaKcH1
ed+uU0ZyGwRiAs3xDWWtLUiPCqS1NyoG0bihIjyHX+s7jsHIAWuHIqQwegwRWM1A
TNmFRyLKncXwCXGDEbsqtwABknpW/HHE/cGOyo1AEjCTDT85mx1JzuyJARXZzJDU
PL48mUlUP+WZ0CfYWVphj5v1A13A9Cqzu7LKIew4vLDHJPnUOZvhnetvgeneujH7
prQ6BXBQwjZa2PCr3t96O07fAUfcC0vK2RnbOO2O02shCEfUPlWadGKHI/87RDEH
RWGBafANVIBXm1hU1LVCXe2zuU2mhR+p+EWqbKnxYu7/XTYjgq7GHmr0pQIgbarj
FhmCqf8E1p+9wq4dOLSLdQ==
`protect END_PROTECTED
