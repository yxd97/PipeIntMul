`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x31V/HfgmDqMafnvmvDa4PODUTPF9c7DUVSsshaD7tsPCxYJqa3gCACAZo8kpBvS
L4afOhNrR2wmgC3NRe4wfidHQ0X3vJhOp03jeBZeoLgaHoO4spaCRU4NQ7OuGnbo
h+VELhjezcj6YAsfY8OmbXaICArzC49yzFpw4xcki7oyKV+//Y3rhoNBuVZ/F4/h
qETDjMxvnrDzIK2QX2aAl/1GwfhchwkwWnhdQG6wcXr+iDFBYucwpe9P6gGlmLvx
LXxFPRmDBTrx/ldobA+e3wOH0uazbEWaZEOXbc5l8kNeUW86l0+chlhleTepjTZs
z6lGI5kbRNw0LvM06Sg+iw==
`protect END_PROTECTED
