`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oM8XPmr/4StKx/KTanfM6JEV+gsbTWd/OkJeBobY5Tk7tXATlKxQQMUtei7ffhNd
QaOebnK4LB2F7H4WtvfbwGIQGJqMiMXH7yJtv++eV3ynDnJSQIy6FHnw+a8UGN6X
4asMS+I7j3BJ0MiXcslOd1mqwT1AJfCNfxxgK8wvNxkHBIn/PCYhn+MaPz8asib6
tZezeJVr2c7vDnveW70Ms+nyzJaR4RN0781sTUwmsHRUpxVfFV9eJLAJ1KBjC+DS
XguFP26Y7Lcq9uA0vmIYQvj0VV8K7fU+2KI0tH/ppKPzGaO24PmoK1AMJaZIAQAS
IvDd167yN7EbwpLJ+7QY7WHKXlOJ19ERdbdQdY7mmRAuDlVkH6dHXmdRq5HuqyrE
fFM4ZAvu6ZzKQWh6FRy8bbziEn3HUtJclngpnF/k2urIly1noKKRXaVRxyEQwNZu
rOccEGl69KChDA+UrG6pLUAsAyPZDy9kwliGdVrm8cmBEWwC+ibCYyGKEtSnnLMO
8+9bZSrbpUa+vElW2oOsQUUGhKBfm5ccHPgmZPb2jBmkXXf7j2j8BQyxHaMkMbK0
f0CRXFbtKvbGxPTfMBLa7/zWYCAzO4SKAIRtFREh9+WzN3pqKL4NkhSKuSZvUnnH
7hEltS5JP02OnfG2cZUS6e8o8/fEHLKiqIpFsv+7MxzfHjn47hBnqdij2zLhg8xL
`protect END_PROTECTED
