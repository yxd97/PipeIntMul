`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sCBQ9CTnSmjtfmTO5SyrcqtZMy8LSTP1E+gggKDClxYw7LRChK4cyMtbQ0IW28F
gZU5EeYpNJ3GTt8JC1S5fIC4mL0D59ehXE1IFemPtUnQMXAA4WoklaPSReubU0cO
0NYIVRIC1+XYEmhdV1w6DyHwaNGYS7iTxFA1prO6f3g+FB7yLljCJmkD4qPn3LJw
1uP8qfJ4Uxxk1rI3XfsW3urrCoLOzlMp/6Fc6ids3O2YXr9Dnu7wJJ8g6AdKyQXM
/XPPC9jMfqCi87YokVr+KmkfAPHLXi/8Dxg3MAESkCJ1V5TKEf4QoEOMAEgDPB8t
B77a+XSkpXZMYQBGJG1WAC7HpcolMcvRzWh8lucKUqRyiw3ItfpiU15RGfM5eyWI
nWYfkW9X0aVsdEIZ65afu7RT9bhEysj3FbnBAxiuf0E=
`protect END_PROTECTED
