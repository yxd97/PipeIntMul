`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4Ongfj9UCUwOc+PteuNR1mYNIUw9vY2zqh1dYheGruv8oKxGNcOtsC04DgzUREg
KoC106utY+fSKryoZt2NvEvcZk7KDd4dbTc+nQfnDs27WvZL4xwMqVsiIEpQOcmr
4WCgG+sHAqg2bMiNrsekR2AhxPESB48vr5u5nmECx4jsIElfFKgfdnwCcFZThc9D
BZA+J813qfFgwMpRYWubzz/7C2U9JPG41qtXbxc1yNhiUTiaXRGnPyD+b+lmiKHv
xw7blzpeQymFKLm9Dd8zcG/yhWDq+AaQBeclJzCZEjztS12vCc4wanIbkSgKWzDF
ybqKuTWLw+Sjtl6x3HIm++1JE7XbJ9Bp/WJjivtqz8RhTrlmo2I1Y512O5FeInQ5
wFbiV/qk8ye0ALeiywRUtceO5aM2BgTcC9VcXolAhNf1e2x6p+AEHgqYr9cPy0i1
wqwtdWl2DhO8RT8jv6KG8cHQHjxEK8BRbbFzGUxpWbaAZgONYh+T9hTFuET7d1Ua
`protect END_PROTECTED
