`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RoJCN0WmLDjKY05yxtplbY/qW0pjRGgfNuY6e5kcl+PQ5meIIL7dHDL4DYoHr9Cp
89ssk5Wvv6uLmLguSUfkwSfXjiGon3fd0UtB2h6iSh4RKJDSM8VHOzcehCOrIHX7
EVMdeQWyieeH0BBG4ZdVuPAssAqMtPromC0T35ehJAgnKznUTBIpbzmABO2peBEQ
kJBKo5TBVfZogs5IaYoEJ9EnPFDTkrpsXxb45V4d5QQblkL814f3P7sdCz6sJfcV
UrH/krnR8U/p3OxJT24nGfDYTCz8ejgF1k9BYx+LMdI=
`protect END_PROTECTED
