`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5bVCUcIDMYgyQk2BD5grxLRm6LETNfRihi9gphvbXU9bj+THETFu0AxAkE0WZdWX
tfY2cMjDE/djnKqlcY8xexW6rlSMFgj+SpgscjklGvspVsZ+wzEqwBE3dF2xTN2I
zUi2Trf2nfedyeBJXISiYZOLINWuNjNypzLAQNbnNPH+VxpZwWfO9HIhMDXPCPrQ
odERCNqyva+uucqeuIHR9OXiKZVZ+1WabH65gHuOm28DKFQ+tBNrKON5LxD8/tGr
0HZUB92/1N/OSNCU5CO6qYpsPBzuS/5RqGfswy8+dkDcIMloWY6EFfD08HIZPMJY
NiCwLHO6VpE2PiWTxiihC3JTpeBbUdbI03DeageZoFp/k5L3w3YOas15JLkB9Qx+
lHzxOXTnSc7/W2Sm1xISIod7wfbamCzK9K0RTOTMRwfzKIJ70QV7IzdytjCsUAbT
e1rMt5luLR2jWpNAl4tebxE5e9W0Ud8FFpu+wyhA3SkJ54F6RKnbZCb8A80QO9FI
`protect END_PROTECTED
