`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s37SF9s7O5/9Gp8Ym2ZV696VlJsSlEQO+pyteW5eJsWYxUwnxvphs5Jp7lYLMnX8
PmGhGEEkokeHjGPbHfIQtxYVrE8qcxcN0JxxULFu/dpSGmfSJa+Nl9X4pDg+yPfy
znyFSDnhLWu4qxLqaGAlkJTNv4SROKUYjaI2S4a4Eau2vRX3A/LuUhgcrBNSFFRh
A0iV4yjBrqwshltFiPJ7sj7ynGvwAZ5pJcdq+lSB+Pr4+EnAmU7pDtUxsnUG1Uj0
85/Vh0RY5kg/+He9YaEnWdLL2S4q4PlYBT+MvyaDEXwO23l7ILLP+6ya/JT+z4kI
vqwsf2DGaC32t7kjhmOpZDsu6obtAL2uYQikV6vAkplZr8FcIsRUe3LJ+oYMEfUN
2ZrlQqwZS746p+Ksj6QwnRn86qHcOCiTD/QvIoTVg5yRDFRyjn/LXGzV/00RFkin
fboQjPNN7YJWnSXNVox0q8mRwgWE7rXBEu/T7/OADCdOvq+xcY+W2Mn8GQwQtMuK
ZO0BmScDAYYmnm8k7h4Nz/pIwsu+f4jUsmLylTMbKFsV83QPp8tsBnt8lWAdjM6K
glw1APp9xJrl9SzwehilSxkfyN9ZcOOepVOnt9RonUUhv7f9XZrn3BRT3m0zRdmc
UPfb1oYBCv/gGYarwbTGBYZyjcGLiG+eUG3v6Fnu6g2j7CSwfDyNCeFylVWBxIBO
E4ecuZQv8FjxFTjNJEwwqfqm+IUoGCQinGDWKlU9DzqXPuKXgsR4isu/wEWbPCp8
xJxBhDcRx6k3Zqjfzcf+RAnMmHCTjt4xEnZ5oeqzb/NaMSKfet5BjJajx3RiutPp
OPmeE6EusuaJivwGQb9cLoRtYESd/muy3bzhEdkiqPg=
`protect END_PROTECTED
