`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pj+oaIx3VMJr2crEOtt1oNB8Dbh+DGxp0/uKDHDwyJv/cxF+xUEZf/ATITqbxXq7
lOyVbEYDeAr1I2XtZxC6ay4DRV8UnO/Lw5ZdN8pNEZxQDrU1V1ccsCr0Fun8tj+Q
d/qjSAgi7kH7ui42nEeaK4Wf1+DTpdM0wUoxqgGshLdqZehF3lY5tPtMgdxN1QcV
RddgYPFyHFWJlIz5O0AT4/qvhyy+ISeyEsyU/LHxaeHn6IfMbN0BjthrKmxIPbcb
DjLOtAPJqzZKWB7plKa7r+Ln8v3+Gzk6BHMHAYWdIyzov78wH4LYqZuRW0SR19Hc
9jfTdnveCXp8BH5zFqh42s/7NryS/tOCWYxPaN47jlrJHCRq8JtzJmQxmN+PG0Wx
MfIdURBvlPPrh64pe23UQ/LZYOwvCkadIjTEaR9A+kfeVrzY3yyxz8So45bF6/ea
H9ltKvgwJnvZUYO/Tw3bxxszpqThnD4drMpYXnq7wnQaznJ2MTVSFdjXWnSswRbR
Hq0Ic4InDhIs9dlumCSjAyFwBXnNNg9MZ+O4B2JEDjZIt6I7Wl1tzaOc6Ex5AHr8
Jwl2Bhzyez3wQs0/sHwONGE34nxYsdiAhmDbQVSkt8MNwizGkHpapKNj/TnEd5Fo
x7vLuEpWWKEtwf/7TBAVDU/c5/R+CCI2wTKNC5EMaReRmZkcCVnv2GM7bj7sK5fU
CPXUOmatCwAu9znkTVX0m+rLVf0MJvBarwynrRnZcSxYNtAtj65BVOExo7ZIYxM0
735rLG6iqZ6JsDvmHuPWhlqbrxYDJWjLlPph3ArcQln9UHAc4b7+F4yRDUB4wG5w
dwDd9vPRcRNd/zRf/j97JYKEdkBT83R9XNjZ0cISKo5uFJ9fAFU1j3qMqwGEb5p9
95lRWkvMbOGTK0iJ47+QuYj+aZIQOM+b6F/Qu+OcDDc9qqcNjKJVie4vF7gNR6Lg
lWWsXwuEt9nRz6b9DT8tqt47KCsgCaJZFMjj+CLiJQjHhZ3gUsQKPLEFbg3FlNaF
E2xgD717K4hWHZK0Uw6Wo2TktBtCCT5Uk39+lr8VqoEoA/P48Tkl+yxevkJgpZQK
+pKgJ5do+Qn+qlpBRHcpuvyuRr4AS7y56Zdz3nnZeNfkS5RZMiFPQnbrcafz/kl+
1+ynBNCtinU/+1cqNuSUnILQujG3hP8uLbC27Xqosju/lIEcTiHj9HkHod8H+7NR
ywHJOHb9YEGxUJc0C8VZRBzkAn3vE6luu+E6vMUkSCAgdTXAsOPZonTdYJKFb/8e
Loh6nAF3nTNBmtXafd22fAz6dTdgHVMrN+E4LeJgZh+KLI9FrjrcfaDCxc3vgG/2
WmRo6VY0OMq1wHx+p7rwKRajPaATRdC9Nf3Fbn2W1tnCLsVfG+/AQPmfU7LBJgd+
Hq0wOd6tDegLjTAIyzCNkluBqo35PY1zTf/GvW4ZgDfQ4yPXrLv0qIsl4v9mf/Qi
6NE9rco+M+K0Yt5xmGt+h6Xzm4XaumJNuv3xrM8ZzUE=
`protect END_PROTECTED
