library verilog;
use verilog.vl_types.all;
entity X_ISERDES_NODELAY is
    generic(
        BITSLIP_ENABLE  : string  := "FALSE";
        DATA_RATE       : string  := "DDR";
        DATA_WIDTH      : integer := 4;
        INIT_Q1         : vl_logic := Hi0;
        INIT_Q2         : vl_logic := Hi0;
        INIT_Q3         : vl_logic := Hi0;
        INIT_Q4         : vl_logic := Hi0;
        INTERFACE_TYPE  : string  := "MEMORY";
        IOBDELAY        : string  := "NONE";
        LOC             : string  := "UNPLACED";
        NUM_CE          : integer := 2;
        OFB_USED        : string  := "FALSE";
        SERDES_MODE     : string  := "MASTER";
        ffinp           : integer := 300;
        mxinp1          : integer := 60;
        mxinp2          : integer := 120;
        ffice           : integer := 300;
        mxice           : integer := 60;
        ffbsc           : integer := 300;
        mxbsc           : integer := 60;
        mxinp1_my       : integer := 0
    );
    port(
        O               : out    vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic;
        Q3              : out    vl_logic;
        Q4              : out    vl_logic;
        Q5              : out    vl_logic;
        Q6              : out    vl_logic;
        SHIFTOUT1       : out    vl_logic;
        SHIFTOUT2       : out    vl_logic;
        BITSLIP         : in     vl_logic;
        CE1             : in     vl_logic;
        CE2             : in     vl_logic;
        CLK             : in     vl_logic;
        CLKB            : in     vl_logic;
        CLKDIV          : in     vl_logic;
        D               : in     vl_logic;
        DDLY            : in     vl_logic;
        OCLK            : in     vl_logic;
        OFB             : in     vl_logic;
        RST             : in     vl_logic;
        SHIFTIN1        : in     vl_logic;
        SHIFTIN2        : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BITSLIP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of DATA_RATE : constant is 1;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of INIT_Q1 : constant is 1;
    attribute mti_svvh_generic_type of INIT_Q2 : constant is 1;
    attribute mti_svvh_generic_type of INIT_Q3 : constant is 1;
    attribute mti_svvh_generic_type of INIT_Q4 : constant is 1;
    attribute mti_svvh_generic_type of INTERFACE_TYPE : constant is 1;
    attribute mti_svvh_generic_type of IOBDELAY : constant is 1;
    attribute mti_svvh_generic_type of LOC : constant is 1;
    attribute mti_svvh_generic_type of NUM_CE : constant is 2;
    attribute mti_svvh_generic_type of OFB_USED : constant is 1;
    attribute mti_svvh_generic_type of SERDES_MODE : constant is 1;
    attribute mti_svvh_generic_type of ffinp : constant is 1;
    attribute mti_svvh_generic_type of mxinp1 : constant is 1;
    attribute mti_svvh_generic_type of mxinp2 : constant is 1;
    attribute mti_svvh_generic_type of ffice : constant is 1;
    attribute mti_svvh_generic_type of mxice : constant is 1;
    attribute mti_svvh_generic_type of ffbsc : constant is 1;
    attribute mti_svvh_generic_type of mxbsc : constant is 1;
    attribute mti_svvh_generic_type of mxinp1_my : constant is 1;
end X_ISERDES_NODELAY;
