`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9DQOHpExHxqHYB98VgfNgSsj2sBSc7UIaM07b7qwTa0ikQ7HSG//AWtv3iFx0Tj
luH1N14TM1B9MvhcRbaSfcRkZjg5HCbcyxC2UZHWfnE6D2ILaxlLdJgSYEAFCuTX
yXOa6wAQ8qesUfOuIcsmZgHM2vQt2BTVFRmWBFJKhWsFYbFK/6GNlQ/g9wfFyswD
aSkrmBZhSg7B2WyO7lIMx4wjmNDJNo003dCoHX22oL0/18USq8ex9ONOirnjxNtD
O/FK1K7Vt3pG6xlliCg0toq92d24EpEZc7onopDzWEkMXToWJgAv6KaoAa9w2nrA
r2IP5eDiw5hdB3BjnC5ncuIE7Ecj4K+91DQpsuYpyglcKglylrKyzRUsX6okFDHm
HNZc+l0mFSCKYV6kVSecBp6rPzG6V0RjxFnlTC8fLe+o+azLI9lOKnFJjjVJHQXr
HzLOVQ6I1MpUi88JNs+f5mXPGec2er9lhDOhi3Ucan1wVfaSNlMd1jqViMs6QtLs
kPDWMumEu/n/whFOkQT9OECU8cfuk/tTCC3DMXH3vxVMdgesIHosyvpqBcmBuUvO
GsYdsoc0WsTLRQXXn/Isgb4UwO9GaL9z84xpTRY8Ajm+yJLcJkRKlnev49cOEeHd
Wh+r9mI/wmmm3npljn5Q6Kv8AR5asX1YxRtgO3w4Xgx/5GsZwuGeysbO8LScZCuu
1SikBb2hklcg+EyDZiFrssDEG1jNccgp/9D2KSeyULxW+kbutL/3NJoGZ2MQpX9g
1o4pQuKCbRpZMblL72YEGhgR8K8atlHoSnAJxF3R08h9DzSKuwChKLJV6h2LcvPT
MlHhDTf4NxgzQV76f/kWplhvCym7jdMSkR8ZFKCtjR9lPGyP+RAXPNp1OsozFjnv
mh6os4/WMR3p72Z03e/sBA2lLXKIO9oy1mOKueUUVj1sgDffKrmsUg4tVoCLeD2Z
3SaVgV4fJyPstiuQ+o7PJDoiOSON2fHrwooTgmFWhDaCJlICYT28SDFI2Y8MJ6a7
DRmF3Jhi0Ws0PxWbLEcKxdNJRIC6j08+GtbzoipROY1MJNCZOdNpvDrRjowX03tY
kEZmW46OJGX5ZVAHADGdil2331ZfFH4SFdytb7MicgBfPYddHUlqsf+NwMLOL32u
bk95WUu/Nstfgw/2/sw/ymdEySmJq7CmPZePQGGgia8o489ImidqmbeVMglI8Dut
iNnqW6uIbfvJWFbOalNziybSf1BX1WNvGY61Ie3R3e/fQbdKo+MzGDJoHMWCmdH9
gOPJFm0DS7kFEry9p59eQFnCiFdzFdCdQDuIMq8jYYSNoOqubMuc4Ycc7+dKTZW3
ENWgAS4HrEWeXEreDY2pZQwD9Y+h283fw27FrTd53CWQlKIIGrxkvZxFdCwGJGfi
cMklFtBz3x2WhYftwPnN5byTCgDXm5b9nKKboAkf5zS5+41tUZkoV2YN6M5HKL0M
vX3NlHKiZty++rOqwrp6zfByaJDjdh9CCV8ooqQicirkTq0+mCHRA9GBQIvXWHVf
Kp3XHQ7gh7UykFVQwKxDoW5eCTQt3AMmuANl+ZwEmDwD10gtpmncgaREdzpUtJ6A
nOvR9bNn2SYsuchFMNEg+5CZq0ws+aVnzSTs9n91py+q8W6Z89MHSpI80IWvKk/T
AUf6b9uEG8k8xrP6TePP+oeoh2kj9j5jL4NoUPSOjZKh5Xa+sTGvsnk7DFNyLB0I
sMUJVQW2yDuHe23jQUEFeouEHie8MF/9IhrrhVxWdPVV9mG6GZaUNNo3YLv59Kog
uoPMu4NBAWJC4N6K3X11kzz3BIWL3g6rt05hmsDvVY4Hi5dwdUjIKE3FshCxbC0U
3I46Esu3u2MWhFUK5NZn55E7ZmQPgzTH7eX+7iikVASAoR/jUzonGjXbhS9pIlDs
DGrBKV/lso4+u63XVXgDoB6Xkh8hl2AHjTfigP+geo5ZbXmDv6rtgoJispPE89x5
2Cl3j/O88TOfQihx26qguZy3TlOOy49bUYuoyEZQWhUa65RXzLSIzW9SidBEC2qq
nckLUvvQFCeLOXMRCotEOgFdRgc7o7MAxcU8aOn/7OXkar1Q2zCpkFUlCUPx6BdQ
ozYPbZRZ21G64sm03VF1tbMGZDZYoEI6ueL+T9HfaBSrNpHYpHsw2xuPNR46DT1e
MNc+4E5s6coDVhrowOF0P/6wWslGqnLJ/XBVsMoGuXZaZm+u1tCpgh/amFyFi/cl
nBpJQyF6qDmH6WDgGptFShyBNYnDfvux2IotQpjWmlEUlw93y4P0NnM6uCzQrUBe
C/lq4a03fsLLj4ndEJlSzNX7qqbtb+I6ZTZSbxGSWIVCdlQJIQ2C3//DTcHtmtvo
7n3m1gmP0vOxsPFuhKcpTC1Q8miFVREu1Hz1YJHsamxkSLedmDfPvI2FSka+j8zl
nFBdiUAjNPEZKVDaz9Vh5My9hvQC7w/6pP5mavhJfSm5Oi56k+0fYwkqFIsBlpNr
d6Hak6D/2PWziBqDs5d92/37Qk7hFaXRnI3KDRtdb75lhEHD7PYNGOw3S7OhsM79
SZaB+uonc0dxoR7M+dXTWVXbGc+gLufbcp1Y6mHzDknRwm2GnDHpylPeGEtY0CEF
o8wd7doREYMHBc4ZN0pAIBiGU1XTa8uzbD4VtKy5wbPOAdWbfh6sxZ5AmlmcCZMs
ePXHtXMN6wAVNOM8b5qQnYcO7Vtia6XwV2wXpBU3S8hZJ1ZPabuMDB1CDmeUxUd2
YqPahBJUZcWFudwYsVA2hsfMD1txNOTb2N7o5aLtJvgyg7oxtqA86rTLBGscRfDP
P05XS6iPydq05CtRXrb1G7TEVTVt6px7eOxUdAC5FVn6msyHt97YePLjXrYAzPkY
MMt5Td5sdYjUvMUQetHEADfhvCpJoYz4DCJKUPdqTNYnJUAYnBpUbpvzhZtiEbHu
Yh4iw+z+YQBqCrnuESeCk0JC1PRGNT2gOFvrRv3mVORxpd11AkL43yDy3FbZAtEq
lmdcqqi5AiTqdWJgI5gG0K3UoO5ALh8x7aflGOz4u7AxUa3X7lb2RuMT9xFdlIcH
H28gwE72QwpeYkJXMEkq3BulWoUx9iCPRRcDm6ApcuAkN97nCE+fSBXLSdETghSK
/VCD4034t8N2Gdli+K1BS4jVwgNNbECqXKQ2xwHb3OVdj5Mv7NyLUB7YTYhJoD8u
3IS806ZzSRMzVavP7DrKHou0LCtzO6vZC1GIO42J/wuhejqf980eJG1IWpX/Lehj
5SKcQS609QmengYNITFNcMxa+qFQDXEEbO6MQfaWvOyKJ0WZgUt4zkk3KKix/Gx0
zWVhnQbIP5bCetVmrzSo9ImKTeXqYknBpvhelTvMkaYx5CBip+eBiiOL3AvCuXil
YGmRcIq+bHu0QbozswT8AEENVo6/Owq/xpB8vIqZGLuEEKbIlf+PjKbKLPPY5irs
vLyf2Si9oPWvWmKcfFnbr62tv+/QYtn/R3K6BycLcIONNRYOwnqK77pzYoHyju2y
okdc8Kz5nQ7kzT83wxehyOCD3zwkzEm4MDlGSdGLEuAlUC9ogbaXWfAm47wCwNHr
a4p8Clf2z8fl8zSnOHGR1r6V1Hj18daFUMLZTREnHBx+kDx6WWMnsJ8d8lijLn1Q
IjfauMeqJX8r5KnPh29x+KzWPCTr+ALXi6l2H7xBIc8gYo6BG3Ay8DizYs7RApJr
MUij1sJLLn3OMNbx4RgIMEbuPstLUz3vMBpsek5Uduvhx9LFjxf4wl3w6wJMAAyA
8FpqSk72AZhCyeBTTZaUXn2P8lgbqQWYzwzHNfq8XqRFdmvcMBDr2hcL5bAHEGVK
bhqVPD90YddLx3+4eysErCplbhoGNLaJ4JrSHDZgHR9fo7XOAzDeL3mfVqKXSWoc
ywOvt7ooU05sakSCmcX5gM0by095536QPAPEoMkzuNC1SsVoXg5VZm27aItyeMpz
iwnwIaj7X3rDEHTbqudEvcLKUq6SjPUWcRnaMiqOTlI6goXAPZtGebdllPdsU+i5
8TG/CmntWPXHXnZMkdEse3vNLAAcVG/sZ4y5Rdx5HpLtDYqpaycaegUhxa7DxaP+
tv7TiV5Osp2VdnVAR+MeXfNaNnAsFaGids74QCWDhlvSoSZPLX4Uz/dQbeHoAlAd
g87Q8EoOcEOVgrOhAR8dS/fz8jKSR8PJYqF2F6ozTjvj1lWOmF0zSb024payKcnp
6OWWb3b994ttiPpu6DIWT6ZakFQZsgRASkYvpswmXbs0oQHCz68msVIKXDgHeMcg
vCPnL76w8WiwFVzvQhBj4udEJOZpJyBzq4Rna10ZLnsUa7iHdT8cT9B6ZciELwO0
eEZYTmt5gHg4UQW1gb71xc4PPSuiUhzVvIMXHUa+krCidOuoJc7N/R4viwBh+5HJ
bjLcQ5kpSJSFHe8ARbut2QojZZ/niVYjyjUDpAL6zvHZDgojSUppvqQG0+AKc8B2
bSEdfos791AZTeB2ggvEeixx51A698HZhav+XVN7pnVC2wyhNFalJo6cQ3XpcStx
8eW7iI0TAf8XmGHg/IIAolnuF+IjpCt6dmjhjyQsSnH25vb4hHwTTxliHS7+tgXR
XM+7YhUPUhj4tUVDNM+yCppn7Kgnng/uWebQNsl7Jtn+NoGO1RoJ8LXAUEIZ+ET/
qvLPYukgrHQ+i4LyFx8RhWeoHvHs/LihH8J3zzLuoDtUCqFcUZRZx6t5yD8bdWbW
mmGTTduDJ6YzPbOHa1U6pof+iVtw31cd4AMhb5cOYlVt3icK0CPYCVvW6yxKkrdE
u33tao01bdlOoN9Vkd/UyJQtyxlu1KZjhbHHNSNHTc8mdHlvn0oe5l0lqi/rVWpo
sMdjEyAsCuB9ZdwGf7MBWEIJF7vo2yIF7mtgYQ/7VFPKSr0/flR1jv+c17SVck2q
IMRH3U+NAOzCVUX4BHD9a0zdnaHzYQRTZdCAKa+uKFG+CLFUvxFuHsvbpAUu/JoG
Y9XUiiEIhnaOIiO5QK+gAsTN5KSj3K9+QLoHJtr1EqIaDdOgDqnDN6hY/kz91AP/
WpTwyDzga5SIhHFEhAiOJP6gfcWRI6woIJd92mCQc7lWmJDipk99dtqCNiTjEHKj
4Y//DIcL7jnb5pWformtKUadebuqejg/7sPlKXLBoqqTj1x5IeQn8HbA7zuzdQ7y
JR5EwY6NNJjXTaKLqgvbsds6WiWB8T4rACYRtoVJIvukvH8/eoJhY4h5wfJ0Vpx3
4oRNFxnj6DNkpS8+vzLZHdbifrevq7+VyUKDoknq3YzzeyXPI6d/7owBtJpw3gE+
XnwHOE7PjDbyUwpkPoPvFeOk80iEP52eMybslWogoTs+TkY3Y+MZvGFP816P3QmD
sQV4ktra8r8OisgUv6e4z9LJ1wEK3n0pElzaMez8xiaZcxhDhoRJ04nL44NeTpku
H2pwuPshFyLMQDWhHnL/oKBAPs3sbFcM6voBrCmZms9+Hwa3JzhZNJXelLqUHlZa
GvlBxFRZMCBoUw74dsoXff1ZKEfYsUue1tAX18irDU9EkEpM25m5srdvEyxbY2vk
K1E/VkOFydlrL8YFqfXKrbhQq+kq8/77FRiGCKvkAFeQ4DaT8htl3/1++Jnv3ekG
wi46/1T5gqoVE+9eQEMmSfkmZ318+N6DkAuCCX9tmNZzmnEghOQx3n+JI+UBM209
MogyTLugCZaEDfcfmpxodJwP7OpSEkO3mPQ5Pm484B+eICoAthGbYPR9P1u6Ic/b
Y9KPcFSXtZjZrWFmyrK0lYGin43akuZnCvcuZ1foyFXHw2CSM664YeojttE5Fv9L
EcqBQOH+pr+dA2pv1W6rn00HKsu9fWyTSlVgDFoY3uxiU1/uU8BKPPZE28I+D2Y3
cZRQ589g7XmwEtfWDnYmjyy2BlMqTlzxaq6gf+sggpsgeYzplRbM8X7V/hgUQC+7
ccwDlqFK/CzBbqOkfOXjR05Bfja5MBHHVkQojfxd+PecGnq2Vb546msxQxnVM7NJ
4ioidEBfcfx+9rXOA7dduIFxmOLr1QklNFlIipVtGO13njDhr5R3uvMYbVy97jOL
h3ngWb07QHHebwfxGX4TRLAMWXrXIVQuf0/dZ0Zxln9VBnLgEA2Td6uuQuk/sfdH
jmo4HD03G6Zh5J37k/dRG7mnFFoJkDapgrDxw0/pjWSrWi74rb6lkJ37+X1qN60/
h2idrtWBN+XPbHA2yPiHMEtv4HA3svuR/Yslc0MmnOr/sbuS7jad87QyrsEXv3W3
g5ewZQE2bP5JmW5jRUvSrRfgwQsJLxTpNY0Ltov70SVE7OI+raGyck1Ze5lZEHXl
H08FcRuOuieCDQs84pPatGzYy3KlUKzQ0LISKQM/x5ABzAyUT+gA3oUrAC8/Ag8v
DBI6Me4dd00woX6FIJDrAEXzAvfTu6NOEc1GAw6assN5bGyF2w16c1FoekF1Q094
kZHrscms4m46iexquzMo46dwk6HAHP3sRrhdahU3qQYa9WkHy2kPPyhbxk23Vbpx
kMmmzG6S5V/Z75PpWKvZ1h9cNJL4x/bvbmrDh3GbiwHQWmOef/ZSJv556xqRR2Bf
OfKe8ItDLteolVtzvagLEqRV9avM44CtBUk0u66Tx8IQdbX8CzByfkAo4Jj7Wu70
BoNNz8EEFp5M5dhNvSwTwViaPgMFLsdYJSamdruLWMZLkijHKtl6MDbbY2m4jmv5
n2idsGMrSEih2mP6shsd5nQ/WrDZrgSIbpEjdfAgMv8SRNT/H1V6XA8nvjEdE1u0
ga1inP/rWIkf0WpT0J2/i3ATwRMlg7yYPvNRvhqS7+kRdCrBqA6nyg5y1l566fzC
l3oFHAD3LKjHlQMog80Q+mChHP20yzrqX0xOQGyJTD1VtO6pB+xZM2Mr3ZfhoiWQ
X1Ie+FozVHWClqxZS1AM0u3yYA5mD0pGiCHdXb0Jd0Qq5ZRh7DuypSMPmZKxA0r4
dks95CMtafy+zP60S/GnpBGSafZf3BrHTw5abm3+8AXpt2smVlyXAwzQWrPuWd2U
n5+zzyKkFhg3HlUWcsEcwQAAeE+9qQ90tY3YDn/8edp5HQKg5LIRJnU1DJRhJU7f
ZPnpQx1Wk0qosmvTqpWvNeuQOfCW/UxnNaE7J//zy5s54gWBeygy/V6sMKCYOJ7f
DuMXzFnleXxqyyxbKMEkjuPJY7NsBoprYHz1dUlDBgqr7CHNmunQ3I7tXzdSEy9E
Dc2Yj3t8pkUyJz0URBBom+LANiuWApWd7izB4Tdfs+ace+Um+C4pil9pWNj2j8Du
7N8o7CHHXPRbnwNAVQfnCos94zRH1wZr+yNwHVrCEdWUh2fpoUC1/faBwuT4+Ri2
EmvVnHA/+9rWUSZTs3t2OdmTzqezqBoyTOxC6N18MBGjvhC6JeJcZn/ldYY/lStp
C8PaYEFDw+Pbjm/hTsFcsj76kLFaLax6Bll5GTFpo99AP6z3/NE6WyfkMnB2LrPc
2cW4hchnppLePiYAC6567MbU2/hZkHvDRSU/v9ttrU/3SXwwXEV1SZgyERkDhJlq
VcH1X0gsEvfMZvfXJh7qkihwy7QwtiWzdRWCo/zaKjQ+oPh7qgGt153v6ow4i00k
z+7HwyVW1ENBo1QYTrzdh1F+U+l3gDXoocyAc/JikLKWfFl3A3gLk5VM0C4cDAPm
tu0C3gw3zOYyH5hp2VPPyvU3RuF1TUh+HODj3WpKoaV6OMbiGHRbrzRCA385jkiw
ekY4EF47gagws6WruW4BEV68gltF+TavurBRo4zHlpzY3KIMim+8e/vsZ3IfyaiG
RQeA/s4W5Ca9e/TjvdsD3pu/5SCZajJbwG5kJJua/BeEEO5aqfUH61W/kkYwbGnO
C29yJ5A9YoYxhLKkevJJoUnHp04nrWuDtj3Mu20wDMpbUpbsKlpI9fTEqWMKYEg5
i8NGfqSaA9GjiIMnISfF00YhGpfb/GnEb9RmHeZ+ZbwqbIr4VmUrxGSt9ij9uk+b
tzYLoq7Jt2iKPK8+H8iGmaldh3Bhw2zdjwCPFZDPn1NMsPfJc888ZbNJfEWYgUr6
cVY31nsWnKT/HYgRuzXOfyVsPvk/VwvpPt/yRVSGUZBpYSPtrmJrRhEbvGTXgiW7
pMAVxUdV2kUTwzN2r8mikFcsROFQo3bZL06lSXdVksVVdvzIjePmwCxEGQlkypfa
9WB8zPVupV/eFNZ4gbWBR+jH5NNVNInDNdefU3+u0hSIKIA9MViQQVMaE6gBvqDW
FNUvG49ggTcrTA0+7d4S/vYOeQWqe/vmfCdm1300/zedByQ+X65hdLXrxQyteOaz
vzXLfNhE5SXLJtOV38Z8Eb1bZyf4tGEAEYKWHKSL52XC35C2V+FGr3RpucX11uvZ
x6JfPlpglFR49I7zrBVvUjFKTU885SZVQ5oT0PVpY3kzyWQARXEn65glX6hC0xjW
mY2r2u7TjRiMdeXYZGxYI15NXpNBkbVlru8M1aXXbjtRYcOAwjBi6G5H9BPriD4w
ca6s7W6rqm/v/RNHe7rKyori+zYoKLZGIuWS5aih0U/KmW9uNO6lHCtClTOH5teZ
bxSY8F8tCOogu3VRWqbcUnPte1W25d1QwJlGXH62eKl6bYIKDL57m0ka4sY4hOQy
gGPkqbCKY5VdXYY7WSkkI/g5rGIXtt0DW9lKSdmnCcU1P/x7QFNSmd0CbznDQmmY
6B7oJq8SgMHV6Q+1hYjXMJbqflooOOyVcpgot+4SepaYwefLnpK4nzPuwIBWzUuk
B+dRajPVqoU6EdxN8QnKjI5Cz60rXYGKEcssHfnsPFf4zb+nMrBUzobC77VOatnb
ul0CxvuDDtttTvYEAHSzAgwgbfBlki4dsmUQU+Yb4Fta6QE4H99K8V0lD1vcns/I
afSCqpfYgl1GyXdlk+xJr3zzWSFs43j+sDLgO/rL3XWARe8cQ/EjzlYcgISKFLGY
J9rR+3CY2T5vrOWv94JZIH90LwMdaoJafqGpv6ERh/bA4IQEX7QFHmO63K1THyy7
MsrcVGzAoIpRUZViBVRfUmrW5X8Pag4wTTsXb3PiBY9KWD3QSphxd0HC3EO1kVXz
AyPRqYTlCe+E7Bzxyj8aYaaQ523tfK5KHl4liG1FsIU+vushtAUyXYFt6gl7z3D7
gHH7jLnUdZ5Ii09/+hPQI0limJIvTLglk4GCOoplNt8DyGS7k1RTzTIpnXN+ovlQ
BJBkpvn3K4Q2d74vV5qXMLgP9pAE9KngNbrV+1JKS1W1lgMNcMfCx6x8cqFkZQsG
JdMi9j+u26OYTivRd+xF5sXb/+sxVyzgaGeK5enOM3IlFm2e3e97C0G2bje91c+l
3H/vdPm5iuAQLKck6Rc5BYxZaiFS+ltTaBlh1FBPwxVHkL92p1OXOnt3Vdt79FuJ
qnCdvuPFrArgU/sAZCu1In/Jgfnsm+d0n2kFncGSYU2ThurJAlOsk6Q/8IKCv+wm
I/cE9B89xvRuTjwgluIxh7FOBMjwM0IJVhWfUz8iXuF/fm7/eMqZSUsZXOBFkBkD
Ua6i0FI/SG79MyGzvdslaU7nYSbpWOHLDAFPeaW2jDRvGpjLyrfsogbsocNzCm6r
6N1xpjRFRcUwhhADhStqLGllTmg0k4HAy87B5Ktt/sJi/O8ZOo32aLtYtDhE6Ot7
sM9muT19t6ZQPuX0XdOJ3G+Q9vlPy5y4xC9tVpw5D2dxZOGXKNyHDR/WNdKZrpbS
aPFODoXKYFfciHVWAfWmLrQhvSMRUYsoQHyQplkicNU8TIBkXqvGUWqEK1KIwjNQ
qCnL5g6bV4SZE1HJz94CbxP6/2s9oRWABxu01/tIub+yeA5+dY/iu6gFVxpQqkwa
SrN8++Zqfh3BmnHG9pnno3Sv4lHXWGVp/w+uIHlA3oSeEVaxG1I3Pz5yXXUmnBDF
ooMT2IdtYyr3strqMrrkxFfiyjmYbILcAJr4SEEJI5bwY10fOzaXZrjYRPNe3rg+
lbhEDGk7xdxGHO0xA5ev6300DKKL51PJba46VXIzv/9mBoKlHxLrbmf3PzbSvP8e
aHPn/3450FqGXeCWzE5zUjtTMRi6OL5KPqWoKOsXxLvgfwvh0STnNSasAtfadkkZ
n96lrIvOzcOa/JbBhYA2/BwLTar63CbLjw4D6kxAdcrP1vqs6BxRlbC4T0+gJtex
HxbmZfNKEgIljFdOoNoN4Zd6O+lenpHUXp52yjzafr45BnbTrOCCm012CPRalVl+
`protect END_PROTECTED
