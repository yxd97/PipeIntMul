`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P++MpO5pAlxBM+O0k4DDbQ8o4Hlnbda8ojvAe1IQAMkYL3s3vjBA/+WrD9ywo0pw
tnc4bntPiaupMSGs3NotkQZz2Ob818cS4TRmH3jqlykE3qwPI5AA847Lcpz3xLmr
gQLJsu5sDm7mc7LzRgvExlmKj5P63ah6TGqIKSQl4Q4vTt6uBMFZkEPM1xJ6wA+7
4njbZT7nrrxFhl6w+C5ovHbdabkrZS46af89rYZ2w6W/JHPzkH43s35MC8AeWGv9
KGIy3I0EiHSe1N+V/rP2ymNzRRJFgdl5nQ4/B5PKnINK7cxcezHSonFS8/P6N2fu
LdAX5Jg8dvBiM2sehCKjGSprkFJ3FlRFf+MVVd986ZMInj0FtQuGO1VeN1Be62r4
Io1lQwW0qW1dL6HrAzMOqyDqF+sjumjLJtGK/TSmZ1Y=
`protect END_PROTECTED
