`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2ov6j8gSiF/jChWJSV/w9agYDo1lIaTaGgMiqAcTsWdLFxmWUMFrfKSQ2YVgdZM
pMYLmgceMtoM2urc7mBVoU6y5SeVjF7Q5kFS0aQAHsa1P8AiSNlbrDqz+GDTsE8a
Z+533jsRxGXpwws/HeB7H4+cg0OG7G6B1KO7b1TWNJMgZ+oRPwhzDNcnFErG8nBn
mx/3jss2ruXFzLp5vZCHET55k00ThpmxEfj+Oi36kUfo/3UTrsoTXskZzGMTCKFU
WSB3GlkN+i+OE+0RvLsGm3ldpDCBs2YmzYZCp5LhXH0WCU2QvRJ4u3NO+NHQDAKU
VKcfxOhxbHyyKhbjGD+RNUbvtKpRNa1KQZ4laEBF1QtFIaONjGb7AZk2dYI6xt8x
LJEEdHufehzb5UjYDifNGnaSUzKBN6zy2rAa0pPlRiYzXaXIj9ayJa+iD0wujmBv
+iYGr2HPX/Suw4UEunuNFlptJoQn3VTYb5CaxCqkfBTtxBwFGhyg5HckEIxPLpSG
`protect END_PROTECTED
