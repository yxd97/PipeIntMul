`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJXgQOCwYvpvpUBx7GBjo3stnvPmB/dZNctZFsIzqDYcHF2FaT6bfg2vYE37HhQo
H9hFUWsaI+fTblF45fZCX+BvrlzS1ObhEKmpaREwIaaRp1nNXejV1FevGwZ0OJ2/
4WV8nlKL4qLSbU7Lnsmt2UB+5yhWd5ehOrQt8Jm+Xbkha4+EsPqiT8+4XY0L2nbD
QPJbrYwKmVPXrf5+1ag0+ZC5whWKZbhOlSWKwlpj/OvO4E7WFVu47504HqS753Uy
x1lpunO1YphpNrhWB70r5CZaOcSkZJkVr78KGENNPEO2mJLul0c8JpLBVVTRGPXw
2MQ4o7l6qpmt/yUE8rRuWKDim06l79J1YSCk/eqn8YeXkToMBFepd6CwwbeON57A
X4Q/HfeFYnTDZB90tLKOK2MnkynSB6vSSz7OehaI2rU49gPaNh6xdPhBukQFAGjU
41JVU3A6bFmEPJ/YDbCl9PKALFE2RyHGtvgUNmoZzYlVbe5s6YW1D3FcTRr123ZC
ztETuM3/H22QOWcWQ5Nun1bl50U+lw33a7GRtgJpULSPqn93bFRDyMEEf4gMZoP+
k1wFlHAfDXPsB4PZK5BytP7YMx0vivzPBnF5AyuQcPHtpStdsNbXWEFyEEpXz+Qv
QdcU8NeE0N0R1FQ4nrKtwhOLCrLj1Rbc64a0PMFvppDuZaSzvq1Tobt0XdCA/fzG
5c9WqjBFEDWbAnatSSvHg4TJyBiqrFJiaGLhqiN+xSKvS1k/KPec+LNDp7D8L5cG
XrotUv+rfWECP++asOSyFfSefW0mAh88rX7A/QUBAsxdc6tosokkMaSRutm7eRGT
QLMKVKhxlGqCVNptV8NXRxoWD7QTDsCH/cnK/AUjxGudui5DpqTq7v31463w7FwY
DpEbUiCcgBnPXKr7rv+wJ2zTa2x8Zr6Grsp2EKTUoiIUfUTaVo4Flv0u9Jk4akdQ
AT3W6avhEB0attFBTokERgR+9/tSIAJxLuXFzVKxE8YNGGXIKkpyAVdxBstg3LGL
r+Q8F5fAPO2lnrbDCokw/AS22bZrcyeQVuDvymXwoxMcnri5BHHcSJkFDeTEmRWK
WgfJJ7WymTP7M/VIue7n8DbCjeZoyH/uHY8x9qAC2/jrlvmhibiWfw4j7wGOK19E
CX+6apB3wkaTorvSF/uNF1V04V5eHjHUcaAUnDrqLAZnmDQD/U6bLX7RstgIhgWg
UgCgCWGEn4AsSuZW0ab/YDb47/U+DjvC0R5V1Tuq013g1YqbOlCHZiHUctYhZqgw
a+gTj7iUw+MGBd+U0fiS1GfqzUfMx4/ioLSxw8SrNFFItboRCCuBAojTggP0icSU
r/qD+5eB7zfrUpjSqEzFRTx3FTxa7AzPu63fFIXQ98kkPXt6T+rRMv5D4YX5YQdC
8NBM6N7bRfOik2Yb84H4PyeKQGmQW9QchuSzWom3zBpKvCdVkD0XuFzXWkmg5Lw4
Re6KRr0uUSDfR5X9qRKeL0uRtUMV9hPNKjae1stGHtPjIYq50EUIan9iC9DxEqJ7
KKxNamZ8XEd5kF1u5OibP+omKwBM/SUJe7/SYmra2PxxlAqFkz7Z9tad1Q9XUzWY
fpp6NrJY0sgX6MGZP3OgY9cQ0ZEl91Gsovuy7OKTTEtojL4BWufVHk5Wti9ZkZxg
Z3rCZA0KhfvtJ/nZKrJh1qImsg3CSD0kKv+CvtDDODP32+mrWiJjb7ln1kKvRLRn
e0k1k6sA7WG9zuBi3zRPU+VkZvixT1tOa5MdEfCsNuA+49xkqGkUla18qGgLgqn6
Ig0MwLq01xnIW43iST2fEHDySCiHDZJrp94Lrzho7A4wAY5XN/BqX84nJ5H5jY7m
yGLSGbRC0B7SwM4BTQc60o0WYpeKrDPRRtNx37VSHp4aumvriPR/hAxhTdpAAgVM
oSH38bPOekKvDepl6FfjRYUgFUYR19cj16uP8Mx6EW18fsSVQPbUv9/RNTH6lLHC
+vU645hwT1GLcTmd4GUADTxj92ekR94wlh+JafqyBWyzNq5rULs8PwztWHYZszhE
ZeZsK5KRdfkld9t3SLR7ZcIExNrt0iNz8xxV1w5gAa71K4g61mOf0q8ZHeY49P4c
cufW4HVLhGI4P8QvZ1fSogS1UE7QhoSV7sQKbLBAsqVgAwnuBc3oJnd0Jfx25EaP
sN9rrAIJdkud9+1W0+ziN6lsUD+wE2HwH6Y3I9AtHzyeuAZS1QUYEriDktr3XX/o
C7YzR7ZQda32/S1H9T3/gc8osWq5ZJvOmNdBNivz/D8e3JeLk6xktj+Hfy246vhO
V4aBVKDhGhT6IOAq6orF+YdbfPbj9/i5Pkv4RA3hUI6exjd3cVd+KPIbYZd5C4Hn
oN8a7WtrSaNm+YG54mCP+wdRtP4NjnBI6q2BVzHM9sa5PKW7oaFFPUwjVumFj3f7
OIcgWmhfsu/Ka0v9lF/9LiY8qRGf4/l2Zk5ZUoTC0i9LQ6TP4+7Hl/EreGbWXU6c
OHEYkChRh+jKAvLjt12LO7G+nD5kkDJzDWLwjDPv0e9NEWUC7VNlKQXpn4pjAhIy
EiqMny2lCVh3yzRtR5AoHL+RyrWQdALwzyNCaTD4c/f75SciVNhMDV0iP5y8yvr8
MCM9g1BdqIRe+4G6EhnsPGQvakOue3xzqF4GQ0WU7fdBqbUIpXoqjDaC4ORkb7dZ
WQrk/NYnARYJ9DI1Ekw8ZL4UEQktbDRBW/CmmiwfwurxyrJk4y0lBkAE9jRYzv8G
3dbTrlwniZg5tNBh0o/OwmzDhmbSBhHAy0cuUwPs/MIj3xeJPBPX33R89+yHIq4Y
SCyhz39nIWQFODvHFgHvQzUa6/t2PR413ikv3FD/2QX078CIZKgUxtvZMooa9U4n
kb6pyyyuiHh5/spINj2L6b0Ewibfxusy+7cbbNMcIA3pUFk4np5PbxfDmag4T/Kb
WtCQPn9ZNQB9nMZSwCZSm9KCt+Suv0tvPmV321uxZ0GrASnUnBEqINXDqVAT6XKE
Tn5tKM/EzcHgT55xDCx0WbBJn3RjmisVCMwwAcr7SeEdMaxSNrysLLTK0eUFDeC1
6q//cJOemriI4vXOqF1hPGklV5NrwzDoFk+uOFZ+Mz8AVEBv2/zavjEF0aSjLrnB
1sc6z3kFvSXGpKBoFd/unVu83pZpntXPhYAHegSqqF3yO8FuhuME7HTISSrqCmbT
ZxB2hVmSq8DceBLV5sfMLLKl3anhhZUkWksnMB7PWEpUwkcAWTh2AAh2Azwn3oA8
6OwbGFgpv1rD7fC+jR8NEJGSELMZHRScAMHCJqnuYN+g+gSAimpYd7qNpn7tcMs+
8X7EP3u1rV0ONw6EVWpPfNYsTAgWDdvTX+aTX354R31IxHVVad9bUTQrkzOpm5yH
zCiBXJoP24bCeIDBjaO3wz8ArZVSMRj4fuE4JD8rxIK4N7sVzaVeL2psKvl3e3P1
8FU6a4O28bsodto4+Jp7WMEv1myylPFio/P0zlASfvuUkdsDQFln6TBMlpQ/9+S4
W1eSqhyItx8wKVbY6BggNH8qjVZPpliJA2GMwdeXA2ihabdSovDJnXLfvIeGSdBu
FJ3B6W8KJTsnJs1y0X10KyF4Lp5mZs7bA2L/7FRbc4TMLkBUsW/bubJJHYR3pqm4
+jNZET4Yc3AMsL7qsukq75HnC+imUolWn8HC08y66UBP4Z/sIAOTADb0CVD79eS9
/E5U4aAiPjX7E2jMUdUYY1qDmIlVE8ENbgoaAxskmpTGajGZMeBBxcBebJ9Ffqpu
GOmNEc3tPbCy5jLk4ow1JT6ID5wWxwjN8Kfzp5vl3v3wRp2sKsAflCP5sUedeohC
8hUv5mz8jqdTeB/MIzHVX4CnL7loRtWHTFA956xXRqol2HHgFWsPT74w6x978KGc
uzj9/lMiSGwYL3YR6SX/noHQzrVyEdJpAHJC6hOIC+9lvHtPjetBrcHez5Ii4ViH
J99Gz1Ymn4CVmpybMfaDAk6t9ybwTFPgOcLU3oIisjOioJCjZckxyM96OVpoaGBk
5j7uUyzk8MhuJtyv5rDSUhu82LPvd4/Xv27nB0yc0l2T638/UJ2PdvU2oIjsK5Gf
blDjwlVblW3/3iFfvm54yJEDG9wh/pRa6uHyQkRf2ZmCQsyNTwh/kg/D7ov+K+MT
7DQ6qhtefq93RwXLlpw/1ywrtbg7IagM1aPmw5YTDVzC1aAmyNCeZ3AePRYhcNSI
KiJg26HCuOtiv+MUCuRBOc4rTWyYnnSCxBBV2LJ3hW08yWoYqBKvF6+SC3z/KzZR
67a0yJNmLlUgB/zd9GlVKOlwYFlNaukMgs9/pxvG+oMaheXSN6gMNYgCv8PaYZxS
6mkZ2Q4YDli7NE4SOlXrATVqZgpxHy1uTTiJuuJV4Yw8y8bF1GIZPm6YGFV4316c
f44httVLGgcjyN2iDFS/0vqG738v1lXQIxfDy8ayN4lXPYDBKVMzshc/GfvgaYdn
SPTtDC3dq/DrFuQJ9x+QQU+SDOiVDS3+ndQYYQuSGxT+ehIYr4cEDJ6/KYEk7Ozv
nYHklTPNDxoF2H3n6N5GEw2s+7fRr+QKivYrjEOcG2ys4cUSMiY6Ns+PBNRXi+5T
fxQrptl8/2/iuO3G/BrX/14HnULDD+p4q3gnaJTOwYpPQh+3YgvG07ZwOghZ65rb
0jzcIDIWRJBd/GqjWct8AEHXUNzdzPhP3BclOI4KbYCxfTsPnHSdTxL25jvVMkvN
sD+aXaEmxyTSOCo0GaHF4goFPlHPhx27sPKwon8i61hiys489xY2HGBK2my2O3q3
xACd3r8LSXX/wb92e0pJmlhQMjsB3y+J7qiRPLLEvor4+1cc1QdR0ujMzGWyMmQs
I0qYMCot7zbfX+Aq/iYIGxtnUqbu796pNtBsBOQwKZWETvZ4e5BA9lt8XLFkFVcU
1r2+fcOUFUUrsfKISoayCwrTxf672H4SRlsdaV4BMUQQvCUaXd+APxBU6LECeg7H
6BR8Q2bSnR57rabUi/PseP7gK3g65pUUcnk2MfFruvxclVkJORD0bI+OW02+B9ux
L1IxaqVxtqFH2vg7FeTAXEVKU+nlEurR8WDXR7qgDD1P/ZNbiGpzbNh7+b5CzjcM
7Q5ka9E5WoI/JskmkrE0puT6ryg9k7+kdS2TslZWGkatzLNzBULZm4JghtaLf6uH
jNQ6/S1I/2GbvQFiPMvqmEAmTfT/X0UR2NeC6Qq4noAZ5rlFElvxOXP3u3OdOna6
UAxTym07Pj0opJZPf/WXKHGJ7lxro2UGRBqbb/Yzq0ropUZcNYqqffFiATXmygl7
gaixbwXu1c+1Im9YS0d6Vt2sWJLcI5BIGx/RKCBYAxKiVTHlaRIbeEz4fY0qq4lE
YSTYwxsF7t0NKfoj90yhfCg7q8t+PyhGTFLDraRkU5GYX8hWjWpwnO2Om8C09zBZ
0b03AhkZ0w8Lr7XLNttqp0fR57yqQy2Kj+LrXJ556sVdOnOgtScjkspfrWr5ETaU
iE59s8UWuyFFuO8JfDmBglMg4Ef1GL7q00hWJB3hnsk/n5CkkQ3iAFBq6LXObTwo
sSjMSnnJd5QpaaQULDHi19jrF45e2J6qkkNw+gPP/lxxnA4X3EdgBW492xAvi6A1
tnoRNMicFMfOtA1cHZSZUBdq1Mp2TX3hd48mT64EZ5Zulcu19JSlGEQn8u369EW/
CrllAxbI5z/GTzWCG3X4lm05mc00d+brRF73ZpVXiwHIMqYpJ7PcEh7GSjMquWT4
GK3735D0DzS1uJfS+vBAS8V9d2Pq1xGwFwhHjZQINjrABoCNP5TlgiLwOjnhGvuS
/2/JUMcEInZAFSa5WA1JE6sbP9owzFLowFsb+05KwKbOBy22ZOHWSGi5p0t6aREb
yGs+NPA+hkQOv/PmQEFTfGsaGAb1DE3vV0iuqj4tQLxpiaeuZsgb8xjmJULyR9AC
oIT3rext/cfROKWmTCG9fFhltNFJuLvbmZ7NKnueCkN1gyb8AlZtnDNBAl7F06A8
Z0miLdLcIhDOXFLDZnb24IZOrSa8108LZAFUpLKLy3AN08h1UuF63EfW0+MDavHe
aui4AmITwCChiFz3RK0vn//u8++bn/2208fV9OpPKdjQI/q+BX9Jq7Y1GhGpJoEJ
btyRTt82L671+EScWXmtEOnjoMX6o6iOD40QPwst+3Os5rxf5ue6USu9rT0vyNAB
UlNiA60o8STLbgpbbRMQ0nK33qA5f6opTIRR+pIQ5Clplb+DZ1BjSAlZEIxE5tJy
DP6NhiUtLfkAInebu7WDcgvfQlMUiN3Oy8NZudbwXFYJIlXWzvrSDd3w3ufL6dRi
ctu4htXU6KCi43r5aVvj5x4i+NoUSYG03T31ZNjBGUgOvrtm3XSOcoNSMsG0fpaq
8nK0cl+leIVq8PAbn0Yqsb+A3pc3kKO6py0wPBAqAP7qn20a1KyCuVuMGo/EoAE8
yZoqQLe1ejUr3C982+tyhrxMDnmN+vMkMEQ6toCVrVOJJgFRycLibrtIpk1PrQO6
xAa9BUOvcsobwQ5lYEfkq/XxWmuTb4J/N+GwoZHd5V0q6E+/b+y4B6eSu4gyqf/8
d54w3YYvPCt8OiIRdYixLaLylkoov2czvlIRsZWBonI7JFeX/qwzYyl+3efvZXJK
Si7yPDDLD42gtB8O+cdjOWJtLeRQB5q+QWHGaYNpwdkSvpUcmL+omIz5M/tJgJ9t
87a+Xm3ZmSslwyl0D5B6LRYBd64McmhFbU3YMG/W/MFWbQUD+7X8sR+b/uCvTHZX
S+gjf+NyHNB507NvRNfsm8uuLj9wYlT6sZ5UyQxa0jxJdLrci/YX03VRGnZpYQ1A
tZ/BmNQgKwaKRhWeXDBQ5ho6BgCopD6Q2a7XbxswamcPGo5Vs/5VBgORdYurxfvi
yArbSQtY6szONWex1QZOAjiKM+QepwnHG2pedBAGmfJ07AsmGPCoioNdsjah9bZ4
wG0y9eV0SPnMSAEp7OfWW6R1AdPKohWWWOwb8vvEg0SoI+wXWxHt7sWBMqEOeCwQ
Y6icz89+EKuaYQOWz7PvT+HRW3HeFPzdqx0vjyuYMWmMehdCfdJXbrM3gNdgMxXQ
fNIKY0AGrrs1+fSAvfdpCAsjiiQrJucDG2EdrC3n56hq3V4nTWMdfqGo7Ma1Fj+G
5khzk3VM6Ic1iuqoe2L5jmhxKbSfH+3XSqwuVPBF7lvnzyv/SPjz5jiM++y4gv7o
jozLir5ZB3JoDvTcpadGxqSOVcxZkeTPccq/z1u3x+1JxA1RYAZ3nIg7Qyit+AjH
SUgFMalkS0FVpUTUOc8BHNbxXEGTS0guRBkz4LPlZaHxQhx8gvWsU6nkD2wfuemD
`protect END_PROTECTED
