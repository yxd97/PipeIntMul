`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fu5aCGXM40CBjBBIwoHAJTSerqOFZwbjXUNHWRrS1xUjOgvO52fn1hJGlxR2eLeZ
gRHnC/1z74fX2EJfeFd8xvN+BbPAIkP6DSgLZFD8RWixrfYftwjPljhiG6ltZ34N
UU03qOhNPHSowX1rkJFa3mDO+cOWDmxibJ8LvqheIeYBaEFf+dKf+FT42Gj+M2/j
zeu2vb1mGpeXrrcwLhY3CU90V/hZ3LPElfa51fqFisGK7Ki6rCUqOKolkdUTNa5g
MofKk/Po2Vjb3I2pVzs0fjoz4nUHqUFJVAYsr0fNhI4PJxof+CpjHAT2/Fq6v44F
G9/zYHgPrxRcE4cMoNQR6aMqc3Q/B+9wxHVuu/Hxrbkf6p2PZCw3kJyhZia/883F
7HEZnqMWTrm6B+dcr42l0CuEurB6MWt5VDBchRlLFkDC3PPptmeumyoOpl6Sl/vV
QMpI2xtV84d1r7eXOdKRRgNprWEDkgIJ5oPwNMHEr3hytI/ZxFteZ4EObUK7oYtp
IQqQOTf3HUokG534nQIrnTInRsUqbGy/Sk5tv5CBPS/Ct0atpYUBgpqXucev5q1F
FmnNxMLVkTfwYbZHdTXLRJerN4+aWiSLCokaq+al5+PBZT9GYNFuIsVcQIHhMDDg
wiWc7F9R/1JgJGZ9hDGW2W5D9Dl6BVHCIeiN1Z+6YnL4MTNwFa4ThRZp34ei/eZf
gP8OFdm5v9VuT2oW2cn3HPgtr9CrVKaNisRWyZ5OFu5/lPFXU7vseyMPNpZab+H9
Ozv8Br2i2YyLolIXkxRNNp3g7rU+cVkqdLi7FAekdX/33o6MnydyHSWTX4mk3h/a
wQj8QmFusz5oTka9yqeogLhwosX8p21QdGUqnU6GDcnWYt4otjcm+aaRne4jgrdV
5n6JqYUzp0II02YZzFRBoxTO98RsfM2ooXqhrh6J/klowVYp3z2Eu1BWgVht6PIa
DnAy0gNSSKEwl6IEda4ye5UdhBTynfEdvsnex+6PQgsnkmwjFr1Vp5uGQaWvC4Ke
jz9oxKrg98FFdj9hIxG43ihItQRnvdQ91sKZvY/JaoiXuNZrrfuW+ccADQnZGzqZ
Xdo+mnVW351EPrTNFhSWJbmBOIW/7XvlQxr9i5LMokF9JE49XExrmG5Mn6yvZMLM
E4yYOseU0sgmy91HWwWQnpcDEu+CA2WS1FZpnMOyudsATXr3w4vQku27BJHz1/wI
CnGR+wsB1nizts/u1bRFUpgrkYwqY8M7bMdViPCwjmOY8c0SGWNW2IKR+pb2esLx
1utqCbRUC3HbliArtaZXyymtq03jdQC50p9Jf9tmPFBtxtKXv1dAPNC4ARdMcxHD
ej7C5Hst5wSFqNHkLvqUx96p0XJ5ujjMCLfiOYsev0djaUkvNNbpezw0pKLp/yBm
4BhrEOisDGkPH+XzfFa1Ljvulplh61KeI5sZQy/muXseDkwrVzLCld/mXCJTGfdg
SVYpwdtWUG7EKtxNnajsLIlY6q2XCeEbmLpZLngzwlQSVsq8VRgpEmgafb2NKXPe
NWs9yqw3Yx8zdDIkX6w6zGXcPHWJJ5lMIO6oUpM+ZkE8R0xhS9uaE50D2+Y4gr3Q
n89BKNRd/j0hzq1AkMEAW7/Vp2Q1ybitFezidNh2hpA4mbCHbxehCvGQt46nOk3P
rb2JCUUHiMJ6ZM874NHvwzcrp+DDyZzSWmWcwtFNJqfgI9VCfIfDUYTUJIn2iW8H
sRPp7Y86oeNQdd+5GOrJ7WTwtXdBSnZn4kv4VgkJxZwcCAxKKDnXeDkXz9AhSJaZ
TEhYwTHu2gaUjnaDfRg5CEUOuvjfswUSZqgqpCtiUidxbFfh2Q3lpsdcmcDmF2ZM
3Z3iv2+2zGe4MqrIcolvTMU2og5PRSCLCqzoNA48c5QmqFZ/uFlkvxzSnKQQnkRG
9dIcAMwRuS+VQPT3h2msSDnuHQOj70qjsltojoVJ3pOWUeWjam0tdVu/miyl/f3A
UKILmBVUq7ipU1AvAKqZpINbuff/MPBdy4yXKoCdO0mW4Z/Fxzv0CYvl8YknU5YG
9HR9TvHC7MYpgFVLqtcI7RjEwIw4DIl+qSYfGAgcPyODpIwA/8fiwPA61P/k+ZiB
UIm6LPPaSTKx9RZWOXozWuUbdJQ0Of2UYuI77nC7BH6k0KQfAzkZRYvFwmrsxNhF
AF47TjuoiOJv1l9MSv+MtLAXlrfTo0cgRfWEgnzU2wM3IZ+VQlft0ug/dFTR32wp
+6Eo5AYuJEKN9HGVetsRVDJmUwBMq03c5yilU0GhTnKe++Plwt9cBVfEjtZZBQbf
f2xx6STtuHq1KvqJ4i1vSHgL14gvrSO9+bFdegTbZ7cChb0x+oHIzJoUGV44da3u
lZ7nMvu+Q1R5Jg7vf2KKNONTOPJV2BnGAYF8uIPcikbPr78X1q7AICUPrU8YLNyR
qLackHaJ6F8KTO8D6r+a84UBSfwGlXqlPM3QG3D7N84MLCEVPzQQcA4l42VQWev0
wRmlr7O9ghNcUsDLNpkSny4jBNGHVC4sXLLhCCq7AUgzFIwjs7EQt0Dfzy0/EpKx
cs79qdfiaywhrM26bFVJXjtBelx5uGIr4OYKooimCjYkhW9Yb3PDuEcTLHVs6K1R
YtdA/bho6ZR1wHvOfBHDuq4ROCzTOgaGuFgtF+Rg22XAgcadNbq4+XdXeyS3HZao
XKUo5s5NSQpMrhbr61QyLbph+iNkIVnMJFAOnZ6uxK/QHmnB4bk1h1IyvQFmvf1S
vn37s1izowLpWchGJzIAzas1C5Se6LrKe37xqGhSHsj9Alwm5z93reHOswxIlQZL
C0lHbzS5lZv82KExUum78rEzeJU97dCbCVtPFudeLIPaPwPsxbpHs0MM0NHgxFsU
oVldcEf0MfmiAGZ7KhMZJ0yxX/Gek0+zcnDLedXXErtzJALQHcqjysAZp8/xT1pe
bPNEvvwCrxVcb9iDudvH7HX3+M0vPp60EUj0jQsduZt6jXmRsJ0grFx7vsa6oC78
uKnxvT+usWSY5gG7G6erz0sZ5npHTw1iKhXVpQWQcSsBQUmxCxBcan5A4vmkquBh
VdWaiOvEu/b3sTgMnDwPNuyd8UbynAElgjjTzqRVAMpGv/P7m5cLrxu2LBoGCOnT
hTxe8WnLQht7Hy8KO5Pw7T8zvzoDPGWbV0rKogNBcidrt5ZsLZkTVhi240yZJrSJ
w87FssuR+G+jdqSIo1ppGj/tTyobBLpYRYIyXBojpDYPVvhmLddQKAaDuYtaG63s
3MWL0z5NWnb5Ebq19aRctIyAPO31EqppHTRqV6jaC2VTotNIM/7pHihxXrbvof/b
7y17ZnM1vGYTHfes1i86aI+qER1y01JIFhUWY+j5oHXWer9Mfk8FdT0MSzFBtUMV
bDWwTHIKzCLO3r9KI4ggdeypKXqbp87okPfZoyt+zZrFhYSvoviMry2w/R3qTSjx
XwyXVb+9XMuHeImJGYs3fYCkETBxIqE6OEqCLmma4U2UnwiwHL6smlLVpEYbXQnB
jTQTpvxpcuz2PfwGtjw6nTLNqHK8vzocY1lckhQ+O2GPJij6HN2pOQoE1ETvEnQO
s6HwyKohl+sFiz573ZEQnr8DEcCX4i68TiNFkvWEuFuOUg0RF8lWT/TlHW6R8Onh
qQed3P20hBjly+Rfq6IgnX6FU5v8blKYdAnpUsUk5UmEp594/w2whVCmIRFozcgP
5eHboL/qU6yCFQ3pov0N1RcKqCiOhR+7xamWS1SnsmpXwqwEPGu/QAp8CXH2auDX
WwQoDDPOeW5upJ7WMSapZRnHdHtf6hg7n8Eel43iVgXkKi4zxGGb+FAre1jA0y9J
6Br4nfXZKQU+G6igd8gbmgaT54h2Yp0I/jBIw1NAuQFowlA9dZn68pGBV7Zqj10a
mGDGcPjCoZm8GtrmZWY3Js1DYZBgsGjzd0x4m3+ENSitvAn5z16kIjrpwZfQY4Mp
VQsbgcdG++yKC/NMHXvRp9TzZoMZ7zVZXMFX6XEnPdQfzKpYI95tAmqdK26Cwwqy
cBeALIAAS7Pk+YXIDpumO9ZXNPU6NNGCsabI5oatSu//0+25KrrWMOidS+5poGM2
0E+ARxjH4/FcAQ+6EyH+KRm92MtHy9iW/oZMQtTNNkKqBhVnsF02i2nlVzAVY/tV
ek6wma+eZv0MxMOWnG/1sbdqwI9TvWjFOCbvYv1qV/8iQVoMYMDpNx8cI6xBUSHT
8fVxC9Gu3pDzaaggrI7cVsamRdMfTyOr4V3sWvEmkvMWKhLjVid3tYiIJgRefIp6
bNx2x4KglwOnCsNIZmAuJ7bs9O/AUO8slp0uBdk2Oexc/c2av4AdTbThWfnyOpOn
/xFqc2nxFMB2ejRTxNrgXwlUqFTjG2e4DwJMkkVdt61MATOV+UXoihe7lpcycMRu
1PHQUGSq/hUoVHEzLb0kNmK3KdSxosBIWxJpF2MnLDmdSw1Lfu5HKkZa+mLrcNqB
OlTrZ3AJ+72X5H7bjGfNj73nj1d5S9StJ7jcEC2MjSqXYHBfy2QFHFDCbbhr9FMY
w076yQvbiLy4Jj+GAlKaORhSQtaZ+O/QHKH4edt5norn6xIvaxfwUoLzuI8LK8Pl
a1cyLq4pHRvTL+YM0Z9fWMY+I22AANCcuYMFxPG65IqhK2Rcje+TLeOLJi9GZoQ2
1kbZ8gAYDM5k+cIsWyZPVpwfx19fZKMQ2UB30Aj3VntLhV6LpBXgudbLKlzo2lZ0
ZFkDnQyH93KbY/hxoO2OPU/nnzZsKwz+muTJsSoPBbSH1TRFdwJ4WQMwI2YtupoE
ZpINCQmYUJDvCJCLDr3gngNq1nZhNutc65V7L8sD5VdJWVuIqvjB9U5SLyss/kv7
r2qz/5wEQ9QxyRC9j76PlxnxWO0ly7Sgjopy6CoOmAgzmYXShP23kn1K2JGa0+PU
H29jJA1eFi3qkkuNAtyzweKWcead8t0WdmlYlWlKs9mev5hCn83RvKB7sc5orWqf
1gMkszpxka4kDio6p3qcCg8S3YbggYSrkTdQs4jH2TvItFo9ATTzNAwZ7d7v3j0W
P1yGn0Frdi6rE1Ac5D4enR6OP8pqy+wzcwW+BSVfTAy8GtpxOITnVwiWRs3QbqAL
3b8ENIK17GvfTQyK4qeSkQO/pRvsdJm7z0W10XV1YcqoaZ8kxfTfoMlPzKPP4HvZ
vJ8qZrATLYYYWf4JfQf7dTloOelHbLW93VsKu1zgJzoOPfSGduGcKulU9W+LiFlf
EJSI5Yo1DbHPR+PoLb8R/Uas+FfxF0yj2OsZgwRoXcw5luDOMkrsXwF4swq0KFN+
+2rPqvVmD74mg9nuF62+gRkKG9lnotxreUz6s7DY3D+4N5ZqgJFuCsT5zNhFk+qD
RedBWJjgiomw8bTLrpePtqgQGEBPNesONu6b+4i9Ayg5H+R+E/JxOe2ZQw5g2sY7
VklcgvOgNyCYLcpjITiCfHiNsqM7rrr+Q7UL9DnTh55yt1RZ0iMhz3fZJOA5bz9G
6185ZUUhgT/r2a54fkksXADkWBisspdW4E2m5sf3MQzsEv+BisYkWGkiiWJ1+QqO
oQqLfVbjUkagKUQeub01huqjpbBcm0vAfV3zVN93E+vxv6AUz6g3daZhv+AB+/Nq
EzhpM9NWrDb21rn6d4g+kNeUD/Jwz3gvAuD7BPGkp2aLTrSHI3MSA4pttd8sUeyQ
q7sZ7UEaHWC2gfCzmVd78ST8Z9+4cmmFlWmIFuQj6c0NWfk/9+VkJnS8Tfb9wKaE
mmCgSjCliRLNztAGSR16bR3E6W8QQzUTCmgmyVqwvb4RMdsV8oM7+mp1PqVxBHU2
C+AJfiy+aps/roVMcoZjNgqtlJ6a9UWag4d/KsVLa29Tjwa2pgwrtjcHEml30p0q
ZZFZH52ob7wH7r/+krBfeeNx4MTgDalNLo/rYrnlvYRaYZxFPBMhDYK5cW7CyNTa
vJVk4j51wD3BMIPdgGuYQlny8O27+i3vHRXizEPpswcOU25Dzjo6qtZzElH1291k
tT9NaPU5s653O78qheBJT1qXj0RAlbw0K2WNxV48Xf2vyvvsM0ILxNVMUVq1fJF1
qsW+qFQf5yKBBeqr+ATQUe04+38hj/WiN6H8dR+Nav6jwvoaKI2jRVqxb0mpcU2N
qJOhBQ/iALKbAQRLOE3FCTK/Y28mJ0rapKZlO7dJNadBOZX2d+cICCWOhbaHFSq5
jn8VdaHuZTp9ovrn7DAyVZDRfGO9LgGtvxEEO25mDnzfW/YkxoFumrwOiuEqU9i2
8j+vxsqPn0hXf7UWxTtoYkAbcT/8QTLvBxU19Twdd9rn6AwQas4EDchxuaD47yXw
ljeTVi+oiZSokWeXyUUNArCDtImEiWuUYQlbMD/7emvSHBKz8a5XtNKTJTupjbmm
lQD0rmLa6TFMEpuwCBuoxtFtU6m3mszoxMEJI+6sZ1gFNrLoDuFBj+0IJqEmEgok
cvAlQ2TmqMdlmuiHM+KWJiLvUbJIvpJgRCGjfIF31nsxtVHOasUcoMfkhHseLYds
4UF4grCd25W5l2BDhYyKQSS5JYQBX37Kt/0i10Dxsu/1Jdzjre6yQu3KO/VlZ8Uk
JYzvpWMPKsudqZRQKHNm5eXonITFaVq4VekNgjo85fHSzqgo2sgnI+QCIgGVUbWU
BFCmvxuYaJEQ9pw4l5qeWXeccotgFswPB05ygGqOZw/MArGsxvteJKO5P2XlAf49
7OR4ru6vovUM+BoEHHdr5vd2t52nhz6kHGQWMJJeEEvRgoGlgeBSw/5A6VvQ1ow+
atMhbF+JwXT+s8sERhMCsqy6ADnoO9yNpFhv+JihKJzjFU6DYZp8VeMt3ygw6Qen
TrVfuAUSYa/nEQNzvxo0zJXaCjNzPBUfcKUa0S6ypknJPpAL8KCwg/z819EaM4uy
uiyqd0rclNi0yGcucd+kxCbIKFcx7c1YsLLtQLsFBSzHrEWg1tdi+UDGZh331zmU
zXwHpCWv5J+9aB/trElFWDzii/TKP5b9rcSnUbe6515p7SpfBptWts03okrTD98J
HTSOo3DsH0JT18il4cnHF9YK4lz4BiYZGR/c0vHXs6Z/02lQkHzxZNclkF8lgq6g
Xa/Y5PKimnmI41gIhnCZwYd1l5FCFCQM0wldGvkc8G13A1jWwJVMqzRHr6UyHaYY
ZnmDWCr19v1CM893kc+icQ==
`protect END_PROTECTED
