`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sP0QqpH9hA/eLcTccBXD/0jnZIVl/7VQYaGIUtMRmPbXAs9N3to/OJDbkQkUqeuD
//Vs9bytcLGu/28K7TkMPfEB37VQVgIzqs5BijgwznDmoqktZk/fEvpbA/8qN7m9
wbRva/rDS+gLuqthhoF08b+SF7KyXuPSI5Dgp/GFB/VkcZ7J9QN/BqZ1vQv2MrW5
nzZRT2f4JBeupltQ29KgwlD8w5gPf21YFCrNJKuvwBbDrN4wLaXNBLeBNa4ea9bh
RCZzOqFvvi+FT1T9YkoWJggvJehwhoeJGQ93zlPdC9uORvvhrZp2HuqIRhM4/fc+
bnb/Gqc3siZTsaNo9D0QzG2urrG+VEiS/YfuPRzWp6WNRP/TTYGUUVKdmyuImMq3
DCQIqhXWrxOWOeAm2kvB0HMc5cnZph8r0/LO6mYy4uXB/zWc4t7tzsgWX+H+hw4B
xebWXJP0KLRwHaLZWFAOOmtI7aUEbgSO+KUkcTqsokrUJHghx9N+nXALCASoeVX2
ReK2sfEboMBcfV4+Pbhx7aiYb826vQhmj8d6uFJVOKFMMR2cOqecifhYdLUNSlyS
3JiKpmzv1MWIv9MnMOl9zKcVCy8PWYiwLIvl/Rjg7czABgz81vKDlUXa6POLULZu
v6AqVmaZGMyRAzYgFghuUGp6fIqoDoalwEGw4OR/NKY7YhSOo/+cWxTDiM1eP2ph
u30A4OZT3m1UR+9U56D+MJXnbVsUECeJlQLW13HhVXDsynkzvi/pCZ7kOTr7Vfty
O3Boa6gS2yM1OUmWKZvXbw==
`protect END_PROTECTED
