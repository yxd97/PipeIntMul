`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Doy6Nub74wYIxrbnwYuDRL7jmH9i+/ENbPVrVwINBW/UIxk9OWUbzu/P72GazG9Z
4qmntq/ZZLvWJ7SCBOBIOV4GKGU8UAU20yJaC6eKeKaN4Ewb1Cm3Sem3La34GRdz
gLQu2JGkLCFalb1VnQ/Xlgx1yg/qI57p4KgIODkJN+SyO0hFcR041vPobVo9LiM5
mT3ieE9zGYhuxoEVYa7unYF3qzLJkDeiaraljXi+6xr1im/4LicC30AxTpfxQe8f
/5wehlNthGP1JhTD+FISUg==
`protect END_PROTECTED
