`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EqWPjDBcYuKlGeN3/HtLPVPrwv/1I6Hx892nZNLh/ubeRtu6sd4sdLxSKKK02IZE
/PGK3DukStpl6UDD6CBFaS+4vCcypg8B7kzjjnH0pi7F3ZAqmVrNx43fCfxseGGK
tAAQfXuBK92LhhfoXFPPvlWgtd8n72o2xbu9RWUf68uqU8cawNb60YyGw196qboD
7BR0ks8EQVRBFDHkI8iNkE0LAc1otLBmuq7+adxRa6Y1hkTR5JJLSfVT5/9KNgAx
yOCMOto8eJ52fjhM70Zw5TMOs2h4SQ4K8k1aoEFmtoGojqez/pB4uwz1RDsyCT0+
wyHDMZzKs2E4Wz0QwEsYrl3mkMPtFTQBMYKl9aLN4t9TmwE26396w0+Xc9goYJ8U
V23iJBz1MPDTl9d2HS3pqPAoAC98zhD640OLkAjmBpY=
`protect END_PROTECTED
