`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wofhu7LWA2vFsjK/csEHHUf1voo4nd7/O/KhSCIpyISFUeBv43y/hLRffszgBFMe
qNnl0maqb0mK8sLUHA2vNpGxYSsSWN/exqVvZjDGhovN+ja86JyYJccCQ0X0SWw9
bOwgOmPppDTxtkjmPadI1ABfKBwotaxEtvzYa6aXMjlUGAcnVq/MAhalw5v+cHSR
Y0JQLGOYFC6JstrZmr5G0YOUIakBGsBH38dRBP7sqnORWmJ3ZhVxIJQw217EWWpV
/I8NHe7hRbObQsDFsNhPnEu1pvd+mdaSkYpFefahrFZlYTSIZMlggEWGkEVBnBaI
vuCpPWBvKKmGLVlQ1MFp3Fw5cvhvwbVEiMzPbwwrZlrFou57ZBS4GVQdlo+MWLil
EMGqPgj7vjkKetD5Uy+Tvrugl700XNK6jhD6WSEOnph1o9b4d1Y1rGCX2AOjXk6q
IEWqc2MiIeHuQnOEHJjGNR60RLgtPKQtrbv/3/xdA6EAxXJq1g4T0ilwkI3vvt3u
clDa+ARYD9i06I2iV4TYysw9HVjoFS6T/rm3DAqmoM8CfAhIgekprWEafQUsWG1B
muyllUD/EdHSP3BY8NJsGSudVRO16EJMk1xU7TcnXCtzsnA+Ie5uyS8btw328sWU
WaEG/yTyb26Mh00ApIw54YWa9axiP2CDP2OmYPwfkogBTVKaKx3PvLQpaGAcFaPN
9rQHb4QeUZbG1AhKqkgCngNW+94RuENyDDQPRgZJu2A9JfcG2vQLPhY3ZJ4hqn43
XkzUH/a0Mp19CR1an13/LvqyEUaBGHJ2Es/PSr7cxvaij1jm1uPHVMraYSpyn4MQ
zMI3YtWGEpfjBk9NUYSj3JrchTt+N7tPIDJ/oCBxcfO0MDpeVQ0VqOqQte7WlFSY
49dRyxZu9Tjbaj91tnD6Ht533j8I5RiDIY9Tshj6itOnQBxehFlIjSCNBOUtTjcz
XNwS9y1Qfmmk8vdg1GSb5fH7lFjvFa99z2FAuXTdA9gwjZAYvP9QBf5wUFzTIdAv
BqWYeiPHVnSEsw9oIUd3NdwzVD/8dWwyh1slAQMVhv/mpMAypp1Q5yVI10dulGyq
bWgGK8wM09HUHd7txCqxKFerpeR8eFciMCc5cVyOlClH7U16+iLDE/VB8729BHdp
SKuzJ/66m/yaIKX1lNKa2jNq4ZrHF+1StcSwwKeqrWTIDzNEr9jeCUaL6PsaGKA5
i148jAsl927LuiCaJ9ESocePEc8Miqq+NJgIQJf3u/W41mzKAhz6RqZqYqQXgmCy
sYkSfBEaB3ySSeE4wwkj03I8HPiBHav4T6ESu36cIKGRWW/pJRabNRmtMEdRSipq
/FiLy8+qyEJjFxT5kHBzwryPvV4nL6KV1K/wrT+d5NQ6GNPk7x2+GQElGuINBd1F
DerJzuT4Pp2iLIdtXvXTg0axM1KVFRqXoqELd+RFWR5uFAerr2yAyXpI4CccW3Kt
hweixpdZzE1aLe3rxJSuDOa5J3lb9cHAM6JtigeNqDG3aLD1CCzT6eKaPIl+AiWC
FzzR8lhDZQkdq9/uLWNl8ZcaeUSCVwtAcuH4tvM86p8lT0KVxZ7vq0S5NpZOOHpb
+4pPzFdYk4WFTGz4y6u43MkdAX0v/7tFrAnFLZ7EEJtQ4cbf9oWV7QnXhHhfgalG
UOT3BEOOXoYfwnThzjKQNW8lvVZELepea9AfKxTe19/ftkBHpiQfZglg5EgwEGWG
vinz/zcERbeBsZOLH0Xho9FeL72ANA5D4Ci26Q4sRpN86wWJhTLBWVhUXkNjiHoN
fGbvIrXC6LQrXcFbMg/9N0CHCjVw5Z/nUUdYfUNVadktS2ZTkabkn/eKD4gIrIVm
dGHdJULr3xZfespYzrz71soBa//yVzMWnjIipPmHIHXFqN8bsd4oB1l/8htS4IWp
HNt7h7d6DVxFh2mUTSrwPHOwBBMMY4lyYViKKkawRuF+IqKDlMQ6xS8I7t/RTsHJ
pfiquu0KgsLNFjHiZv+QAF05q6lcO3X3NBLgkar/sezFqFKqdJdN71CGlliYgaEz
HvrvwptApZk8R1cJmAzrda4O4MHODSE/7gYy0ourxD8=
`protect END_PROTECTED
