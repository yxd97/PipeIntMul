`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+G6XcjZHaYrE1CTheejGeVJGv7z2Ycmiz5R5skwBOZVAxl28h2owjnfVeKSlxhN
oQ+b+Px6Zz6wEZeLCLeCJVvhj6OvvCeBjyJ2d7Ly1DbtsiGygmzb5c6Ck7U/YFIC
rLMmSxFrxSDlHqysq9uRDX/21qRIbiDotj6NgFdbRv8Q8jSVIps26XZlcRKycak7
dSMMRvw6VMmo2RFK2eMk1SAzit1pq/Xzn5FF/+ZlpXZChD/Shvyp4tB0jpnY1jiG
Tzs9/Cw7/RsNCGIKdSOHlOen6IpUFS8bHSIDyNc2uAkEyEiu1xvDCIT/NvEhN3gD
KbKTGM7Hi2xy0Jnq81kAaC0OlSzypjH7hfVxO8Yum4z1hfQN71aD5+TAPUSfpCNK
c3gejMcU612khm6Kn/RXKZdbiU0tpXnxlm/X+YE7lC4hGhrqz25B93zY/LXbvZ+z
KnVaH/nhfVmitFX9k4s64buKjsLlmw4VRfAqGAIRAaBWYg2wsQd9VfLrySfxPVy6
P0X6eM7L4V4kfdvZBm59GB95K3D6ihNPEnEU5wgC1jst32buhKfQsJoMSareFXpD
`protect END_PROTECTED
