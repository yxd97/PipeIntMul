`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0EVZsTVikkca9Hdjty3D78DUWGOFOfK2u/YAMSCIMZZVbDTlAXnr/+aHL4u2qyJR
eOxkeSj2vSdoznRUgs3vcRtrx+saeEwCntMzR+RxGKqYsfUf/qdx1KUHh1h+8zOM
N68sOdVpHeGA8pWUdstT7JEhuYK/OLFIjiN1+drcSBuh7OgpwnYAcl/zWSrm1WoK
NsNdNbtKw3APBubQInQpGPKvAievE4lYxRvH+3zME7l8ctDnXzZ6pHipx/JuUCEo
mkhKnrYZWnlnz4YK4K+iA/Fgbs1MyHYTlgD6t0pSSC2Jy63ZN8irD/JMNwaXAp2z
5DL4VBXS0S7LLkVJ12A2k+NTXIyY71p9TVyY1ftzv2g419xJfsK0CxsWVxKTMFiw
xJ6ds1LkCA02sGsrcHQPPcviZWaj4F1Xs1NrUGmZIdvo/NoMXTTCx5Ozj3lrjlXS
`protect END_PROTECTED
