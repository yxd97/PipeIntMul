`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uVe7wOt5QsFIPuzSsvwY6V4Mt9aglRBbgfQUBIK0rGFqcvmMnRIsKpx103rsq8ET
SS11GAVDtIiSp4F5njU67v75Jv/9EHvV+Pz2K50YDyzEulioURCaH49BX3T1i6Ry
I00mZIpRqrdrc76nGtwRDQ3h08ucTP5NH7NT8adDzcjXqbdAOrKo5p4qxcjwkLg1
eAAhIZApcgJC1y+8yvDXJzYOErC9RSghi940CN/utmTMesMp2TB4BXWRwPukCoLz
DTPBwEK5MFysa5ok113idDRXqPGzpLwXScck3t7dOWjrgyDY3SfKA4/DFCOG+AQq
wJe/p1FoAycJ67BDcSdD3A==
`protect END_PROTECTED
