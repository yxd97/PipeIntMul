`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eG0JKKgG/7ZO9M1EtxbLZxOIrsRxm0z8mORlciqsvFW+gW0FW0SmXSDWk6qsZahC
txawLfNiDYv2wWGl2DWdXOSKGS+a2mEeltrLyRRHNNvwcNof7JDyC/r4ScK1hio/
akPK7aVKKALDbiCNcUkSp5UdLqL48VDiNEhfH0EdWZpGhlvAA+sFriD+0fKWhw68
WBFVmoLe76PXti1vr/1cBz+j8lVhPKJyTli/qdimb4kKYBHY1mqYLiQmOSEFjo92
klEGrOkM8blLRx9mRY+Vp7YcWFRXH9+XBjSWJiceVOKVH9M22s2HCaGbtiXRI+Ot
mLPsedfbswu72IJ/VWvBdLVnDCtMbzfxa3a25XjC73rhtP+W7s1g4rwD9esR1FZk
z6sOmtUtBhljwu79Y+cL1Q==
`protect END_PROTECTED
