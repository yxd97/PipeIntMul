`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihY/BYRilV1+3uhd9MgeaFrGCoXBjD4+0FRvqvoPNj2Ag0n3QE6s6YMsQfS1dqvx
sa35ta2uLjCxr5Tl0a/XVLPlZkskSty7jegETwZ93IDhB0Kc+Lgurai59CT3QXH+
z2kHs1D+MHT0euf7zXRHwjCaKzJ70Qg9guJyUPQmfo0utlAik3FZgYogg/ZNVeiR
1xXncfidEspkZilL6itjKurXiPUp2KLnWEksBstSQmC1UffgaXhfM+DDJBMl03X5
S7TU/5jIbfWi3Vlr85y7WhW3OP85TcTcY/wtW+YKElOke/xWXu5uxvoaDNfVjvZ7
eFB65AjAhvk18bfXPNEkOdkbeNhyvpBZqAWJnfMoPJxazjHoNVOwAInMpkiEy7UR
FN/F00RF8E7wr3KKX9NpWgaaisBSj11ljn2gI6d/CMi/VuB/2ZpbKaY4vXJTbywK
`protect END_PROTECTED
