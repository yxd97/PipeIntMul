`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYc1G9U/5QGLptutlDWli29Yyg5ZP6gLPJH9pGbsqblGHdBshugJYVaKA6obF16m
ib2zRqHjjdvU6soncSElmk2IdKPq7Fr/PRWCw2mUZqAzHqfAr0ivp9La68FdquS9
CQ7753dRtdx02VOAguvT//0Wt/+mOLqd5QPIN5VO9wnIQMQ0VOaVWCS4cobMPEWg
GMaS0G9KYHkUz/RTXox6/Ya+79tVDmW2vqiNGaP1N9Vab/vvVkq07ENk0ghLX5AX
3S3wdC1bA3u1F6zA3YOaVuVhCk4PY6eZVrJPiMxy5vfw5F/37tG2DyLMIWPEqXf6
9ET4WDXufHMCJEsE61tNfQZt7+vFHb4ybIlOBUi6WxSQ40wXvHz4ryssjonwy5rK
UYk/ZRorUo7jOwBsnWYjmHgf8AW0haw7EqM06LYJLCrf0KrPA7M9dg7nXYQZLg2U
3Y00lx16UCp9Ru4UDZyjYTGBmfSK5xWFUNLpdhQE7b2q/m68EjoVQHOnq7JjIMVM
1YGRQNzZcPGXLtwrr030TaolzuUlcJssSUKwsDi5B1c8te9txMo4BF1EzWXeiu1f
JH83qf0H1CFqboGoET6kTy40MeIv8JthYee6UkkmiURTioDVo5jd9aRVp/7UCZ8B
z94Kh7iuxmsS+T3uDD9KB+j5hX3VxCJaXRJeJOYqNHc=
`protect END_PROTECTED
