`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjrB0qoetPAOO3k4NhlRj/4eWqhhGxbq07rFnMuh2zIpOXqMmD77EjEsdCjJC6Ua
MW3veLniqfx2OOP7iNtkxGxlK4Gz8/YpEwIJraI55Nc2AlXIKBmk/lOfCwcf8iHh
T1euoNlBIg0bFgcmnGTTf5E9jk016/cPnD/OkIPygMXd0VZO6lLmW6oGAmPItNp4
udtONVlB6mAHSn2JaAmGFITTk3POe/DcasoeoBuWI9kuw4nmNwZaayOHxkthWEQJ
tXHyNzv1Ked3SJnGofl5h11AtHykCAKRbT2Y1Z2HzMbvGQDv2TBfTCJeag4gBTbt
7JCV9ghA8sPV+ZpqQOmVKRoQraxvXxtKcehRVGArCHBGst5AHCAsbZJR6L6oi63Z
/Rejw1e72/8Bf+DQ4RSCJaEQklWQyefM+zKJTxGDAYwO6IY3JaDEYrlj3sxyhKyd
PbNBI7yBuANqj1Pz6VuM1ISchOgIjZiWJcr1ozat6zxDoRUEUt2XVOVwAqdQMSpo
`protect END_PROTECTED
