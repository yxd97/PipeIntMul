`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlIIB7o4P+pa0DbyHoMixzDiPC9t0wwlt265C6X5d8YOAlBumir9dXo9XiB7H/1G
nZkTX6I0/Tun6xToak2Vd2QkreBEXKtMLPhZe7EZy4O1dNw4lE5vjP7vBCEmpdbO
emt73rHGR1+OgGLXHtcH6oPg5bhKD9OkTF5yLaZUzD8V6s5xvr71hHYisKEYPqCt
eVyr+bWTj4KLTbhSok/2shys3o9CI3x6cVw2NYG7WmDbkeAUx2o1l9sVU0/nHqKs
HOtvtWCivDseHJ/ENBstmzrtNtHV145pKdCMS7fYRAgLtBSBrhEp9m6dtGvYkonD
K5xPdfVFrvlx9AqEZD6bI8jcF8RWrEoLeIDPDKbGuopZ3NZ8H3o7/qCgtIsg0sHH
J6aXxRv0CT6UPu1+EkduBoTJ+kLOnRx2gYez2V4s+MQ=
`protect END_PROTECTED
