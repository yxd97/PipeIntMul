`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rS/J3XtLQKO2Zxzh7CHop/t5rvJGaMckr/X3JitGBRyK9t5PZscXh2YBs/adJdKP
XqYnWqP2ALu8oeadsv/ADzsrAGp1XfSoRewt3Kvexr8BjIgQlg7P/nIiF2j5npp/
IgtrO1Q5Q+4KS403wdze3AmMw083DRPDRcAkHz5ih5w9001+qsmgyUM5DuJDISk9
sD0VELCoualaPhYM8gl8l+UjGX/QXWCskJwNrqkPYcrngD6hgZ6HpuO3uribJY2V
iekspjSwTtMwhZXzMRB3oPzWetOtpZhJSsXxJ46D75Q5Ftb515xwWSs+n2yfmB1/
jl2Q6CVXJ+Umw/D6VXOwRcQClVtTzERbSuH/mdxWYVhK8csBf11EF/08GM2jymJ4
b+LsLhd4s5WXcfv/7hFfLbUGpB+drL9z7JOBlXqtqn8nvtlwZA5Cr00QEAzPCmvb
BUyCah5+ctsbyBcjaedKF5LM/GfsANsj822d7p8BRUXUnIDOxZ/TRe8eIHzesqIw
cjXiIrLVxagvBINTt+CnWkKrtm0Dkl5MWFCBSbUZLAn0JVLnJ/7GaUJMEO+34Xqh
dqqT5mKKERKLvJMSckjXC+SofafUKQfwXPnXvdrVWLPZTthKIqneUd4ThlQsGEN/
wOSblb96F3Iqfal6pGXLqPB1cqg5GpMGUlZmD3hOJIOxiC1bekyM8IkiLQdSgvoV
N57nHHgARcgVk9EsuTjOJ5spykpi0bLe8kFui69fUsZPBSVQwCOLVVy9tcnT3vG4
DV0b5TKJ2LxfFrKdDuOpl+Sg8Re5NFn7MIorJVzqexOOH6B2dr9XXYsR50s+4wh8
Rx9rZBzoBQjXkM/dloBHjCUc/SplazQq4OXEm4WOnWl+wgHUoSF69UigMmS/19U8
jAgOwd9y5u6MH2dV7qcxIRvtqRt7zJpA67FrmD+/j8zT+9nkIc4AdQK2aK3gcrcx
mcrjTzXoFtrAJen2L6pXVdJntwvgmtMzsevtHl88uqjRkC2o+PZS+c9AAbfs9VLX
jf79o6GrFlTHeDrV/0mTHE/MjedxBOfyqnwLhazIyQOOIvsZOyOKdQsZzMOT4Sbk
/ho2mlH9ExRKZku6tEx2dgYvSBpQ3ffXxH7fcnwv8gxPWKTijCbsH9KC5ZNnDiAo
Quioh+C4i+wfyq/6atx99TYwaXX2khqI3B8H5LXO/5Vc5nAlHl7Kr3gho1Hin8Uk
NmQIjL23NqGX6jNVJ9jB5XRM+hMWcjExBwMNDPJqmaJD+yev4wIhWmRz7n35+qJM
YdE5p0NnGfsteI3ZahwYzICSHcrHVDJr/XdRItRL3/kHF6ibgcIVFD2fFsIZVIik
BP0R95nctZcQ/nJQ8JatIn7NGUT98GKpv0p26NsAkEyGY131Zc7sxUWEl/Pn7OdD
eMHxJuXNvDpMg58OE7xW9n7qy0jtynBHcQzK0Pz/GXy4UXEsPaXZQps6TO1T9Fv2
Zkgnk0GB20xEsXFav8zeSEfdm65/XXKK1eDRdncnHK8/WrMjgLHUie4TTkAdURxP
`protect END_PROTECTED
