`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rG14bJL9xIhK0HSvCNDU+rSZU+TKKNufMrbfbDL6sMh0gGfd3ktFCJ3rvv584em
rkq5jTRm3SX9VVBaQiTeY+dV+/dj2OISWZXRHZ2CLhY594/33AETi2rYvwSRbuG0
A3ywh17Fo1JEJJZGL+QlVWtYv/0OmLFc3RMsHnzT5f+T6vYtCJsrF/tFzNnghehH
i/QYb2v0TF0CnlG8DGIj/PirS7/i62SppM+NHjEvcU+RYBVetosouDTzubt6cxz6
AWD5fssi2yoydLm9AcxohJ5RIOf5CQRXX0aBP7ur5hohGcm3A8RHy/uRlpwyYrWQ
p4d48u8W3BlA8cfJ+g0jCUBc5z2WQ+7DxQev3CpMxdhK0HvIcFGLAvt5KcmlPyAB
AjmHxe5o6ZMIw8B80m17bOpsFQtSrImQE6imWI+oztc/8PnDvVa7nraHkJ3zH7qV
vsXgEN/7ZXknPRVxEEVbKp28Bn5IH/08d/XrbgeeOL/6kpzRoJmtiuVjZf+jogmQ
Wsf89XHRmG+s5DCxOU80yIeUMBEWjPqWmGmTq6lB0G+BzTqAZb65y9D2ogjVSKtb
PzsJqEJQ4SN53eoOCLMQFh9Y1oLY3v8emGijKU+vua+HewIKeT5BC+pHB3oLfDOi
kboxUV9E/7lvTKMDMgGESMN6IYOJLlnhNUVhCidZtxsoASLEA2eojwozCc7foPan
RGu6qoN09K8c/kc4ewVfMdYiHLmBOfcS+22FhFQ+BiWNuWU+UpiKcjZOeRg8NpXP
+xIx9lpOCBarj0RLJ3TmZcNsPdvBLvGkd2UHpW3PpjJTmOqCpTEqD2lYGWCpoMJb
Dt6UUwJ1Q9l1bqeyFIIJAV/anjwLrvrDB84bpH4Fd7ldYjiaJV+rk0peF+5J7WRi
3M/pivghnDbpeeRcA2GO1ClvtuLqg84o1mgvFkaogyr3B8uJnSgLtm5UvLzAdnpk
WQ4ogZ4/lHGmiZvKM8zjjuK6bPuXqQQ4X0yxK8dPxmQjfn4sOFQ3A9HSk2WPUTiz
kBoyooXO9UC8AQjiuz2LY5+SQn3QsleTwBva83Va6pGcCgKp55cbLqpwJ6LqGrKb
r2V+2kqRATBAUpNJ51Rw5QBXgZnAacVyX9TPLUkwpg7AlIniKXsTT6s80+Ns8Kpy
4Z2LZRNk25KdZY7YGjPLsNi7emneTsDD/s4F7MOxX65KqmBeHsRb2QE2RhicpOVP
EF+NTgaFJYdOzISnE+48ehJVIdmQ6eEx7PLf5Zm+dakX+gplaK1Lo0cBjY/XOFUp
X/aA9/gn47q9GZv3MTdnGctsVgzSuy2V4p/ygGSEpOMzmRcbIko7UvSXdGvVEAIV
v2msqErrFA5VdXFwEaHA+mveP6xqQSbU0pYFN2weIlAdAswQe86/6ePXEMoMpvPZ
osMNs4hGRhoedWae7D+WnV8EhphKdszmfXNytPjX8gPRRlJqj2KP6c9/kIkyAr+Q
DRzoFuPzGwa1RvuRWvDPSvpaibuF9BudNIrW7Y3CrzVScEI+1SQzU60FJZdSIvWu
Dn97e85SdUO9mJPbhGAb92uutJjd70QzadRnWmI3ed4Egou5oKo9obMp2VDapX0Z
LvuEYacOM32S/j/+xWOKI1ov6e1Jhjv6DYToZbYa0TUG5dssXRGRvBSjw/QV1Fj6
q4vfwwmVzvnxSIBIjhfTamZtVPQ0L7jozXesYaNwKBZWi9GN5yFLNLl3UZO3e1Uy
J/o6neKBayIeuG4pCMQfPrwzlL+pXVyfPcmUAc5VQhSvdYtLt3vcMuF43UshJ4aR
Xj65WBJfCwqqFPNJu3sXbl+ApWJ7H/zXdKRFMQ12Eas/zMy78Tdyhux8Q6JHQHET
SiXXuyLuFXo2MKdWm8nW9i6HdZ+U29lYUD+Ef9x1C6fnZDR8WmaK2jCiA/UvwkE1
n0QdaaLW6gw9H9PP0qB7awj/D7/JQYb56Ji5zwgt9sMtTWehMo7h954uKDrDuVUU
R/GxLreDRL6RUJP/vY21k09yKXle1dVFIJk7ERpbTMQVqcZvEAV1h9EdUdmQ5vyG
If7KgROgsYZhfKnbWV3ppt7lMbYGmbZD5PPiXCt2Wuse5zcB8XqJ5P6LFfACxUeq
QwnnT9E7n4d7zV3Xlrt+Doi4n9x62IjUfVU38O2fflxnBEluaagv3PiuPw8zSO+7
M1aLQkNBfPTBQn0Hc+no2D9ogqSmhXM3YiZu0TXvYruEGgE2mCEO8kZW3Ja23AKo
8BiHZYreTRcPlYjfXtv3UnlSt67aSJAs7572KXAkuUqRJeL+cF8DRdffNqVS46qt
OIwX9TKgMFw/TunoEJOyvDHIUFlKIEn0vJG+zpeJ6u/IRZ+62y2QPpu5yZKOwnTT
91XSWqcgDXT7pj0C0PWpVvZDtdtawHRYuAdPv2q694UlRHbN9SU0n5+hIgWrD1BZ
M55/q5A26uzUA14pEp8jjc/IqV65VyhcukzG281JJZBM7GBOAukI+OIJk7oP17FM
+4mcXnhG2OhtC7d0fTv6GAuZXsVPXNbNIF3mWZEVrbnGysSQvkDOFj12DJFqXgwU
E0C/lwFK5dJDdp650sOxi5wSYCDcuNUW+wEvSFMd0YMzZaNZBc7m89LwuIthCe4s
zNhvbvAYBmQPJlof1mNL+6LRxRSdym6p9OP3nDnQ5DmH96vNUkIo1VNFV9MjyI4j
bGJS5x51c6hGkUUGcCtwr/7NjCQPUrU+8A/p7G+pemqwvRqfbO40tNdu7MKeh0ti
IRkIRqisRvQTNfui3PYyUn0CwsbXXhRyWtzahzHV8muQCOGB4cdNaWL9GFzOxmEf
unfgBbs+LgjTphsdCjUCptGPNFfvg4ERIW8n9pfeTnBE6TOylJr0gPFmwJ5Ysrqq
Jhjby93+1y/Bgj96Igld5A==
`protect END_PROTECTED
