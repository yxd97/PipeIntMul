`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5PfQHQ+ZH7hQflVzVGmYhx6jJVZY9bvMgQtWqx63a7QjpQ1ozKgF8sHnPwTHs7ll
WldEuaSWeVRzeap39nDAyLRwg8LyhXNAK7rs44Berz6OdBejiOlU8KKtG0UX0mPw
sIYat9Y90usgyrPRXVYDAWn5l1qn0GobDPKqq9YiGK/nXpwmg2JJVzCljR4y+szP
ZolFpjpW6aofGGfpjia+L4VjUDCTmgkLifd1YMZ9R8vG2RP1SlgmJ3t6DeZtbN5t
Ex08APt++sdBKAdF3yw7teGYMubHh8+nwp1lxR+BqdEVCA1y7Gjx5eFOxlQZi6LE
/ko34otHw7bZkZFtIHyvLPfyUjlbBF4C17MgFHbh6txYa+Tu9Ok1Z5wDUfiomO8g
17s48RlyTsagn0tF86rmyPUtJ0iuKttwMV/pt9eG53UEtcHplwyZ5RkCQo1/MPGu
sQndPqZaFkbraraiudyaeWSGmtGrnKwHb2RJUj0vcvMcOibM9VoOBVVUysH6D2Ox
q3MfNxynumgF8vBkOGuj2XyoFYIONvQkxcpvnukPe7MTzCUyQp6trF9HergM2bPt
kDISE6BIFnYAMzdM47hqtGuzw1lVeFokLtpyMOKK0g6GzYHso0xSTsxLRDP3+2W9
4Lgd+rWnInOZNX61snBBM9pQ5NcxtuYgt0b/QZT0yfyvFbepnIS3Le+IHVuwVs7m
Wk3re1AGfumALFVJRdXe4eilGcowMw1FSG9M8YV55VyZyC4+JhTvsSyLQbqb5lLM
Xm2fbnRYbxRmapEczYcPUQ==
`protect END_PROTECTED
