`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2SfE04qxtukAnsZSsr8mlruvk/aKXdzcdtO/BH92JqUivV87X1WFwcIy2jXApl4z
Z83iORJ3rvY2MA2t67rZZseVlRlgEjC5A6AO/468bI/qz2MBTf0FvW/9R2DeG99c
zviTNJhp+3JFgWveukGK2Xkac8J9e2E02BY1rJDdzpEVsACMVftk3KrXuwxoEM+t
5Dzt9ynDNVFEVes/aHIm/916/CtgwifHEWqgDB65+nHEFYYADLKzhL30icWSv8uK
NNH6RkarUSSgwUhwlLcWrOfZ6eVnmGBMecrYkMw50mVwDHIe9H6Xd4+1QYVjQlAZ
acDrYqBqDPbBGlqnO3fUDuZ5R2vBfy8Eg1JzB7DY40dL0lexo1qnHS5xDZdP6v5d
DMpWXazGIL3iGAOWsx+sdaPJd6q/eD8h6Y45iL0gchfSpG5QHNU0X4sGeEX/tsf/
`protect END_PROTECTED
