`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VUPJRei6tEO4PohsgCCyy8F0i5/n23Nnp8BmCQugpqsj91RiDJVTOCoYqjfFpM3h
CpHfFopauf1woVvOiTc/iX1wAbRec9QgW8gvzo5j9nMCiIE39oF6FRw1Q2RVx9BN
+h6AeuDY90vJrTM/hveXLVkc4rMURSgViuSQJ4VPUsBmnw/8QbwaaC5KyfEVsw5e
LoKus3119W+WrWSfasUjdMDMPKtANGGk8VqC+ZHvIXgpLKscJrf/bBWPK6zB3OI1
dd3wUt3ZyhbBbYggGUl/Mbn6MIwIVs9kWdirRA1PyJyyb3YgaaXIULWNQqq1erC6
RCSgEUBn5IUx2mWc/UCGdZ/J6ST6owXWJNtMUufufMlyXBmjlDE502mnq7+iylN4
ZmGD3L2s3PJAXlQRKvNprUrK/7GPIKvfHZJAw5BJJ3oNwQUUU2Yei1GqT8pp8fB+
0zN/tLByo7Y4hNLdvLMd3sNO71lV5zuCahSAEM8UZVsu2QHXMZCxDIpyUdvSWd8y
SMcxCsekoosb/YNodenKzU/uA6JBOcJ2+LYvqnsvGAfHARg7EKR+aX1P6gOu89zk
BQYeVMkjnIOqwjfQjKo2HreiQme5i1ZdzXhrlHFCMgGh4AtiRfLbSvHCJBKMiL0E
+IyEA2rkZJCL2l7r4V2e5A==
`protect END_PROTECTED
