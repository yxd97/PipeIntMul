`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HN71dTPermHT5Icov7nry//V9BEyi9e5xPFj1KEr69pYQS6dh6TnPcnlahLfKHzs
CZ23qLFIEdfSEaEgUcZkZbuH6RxERHLgI3DZ2NiVrAg+3wwioPmPLXI27bDVSr1V
2uycE3V/qJuUJ9f0BCylbA8WnQPM5lDIKyukQzxnBvo1sfpWD4+jexxYDOG4GytT
Qcc3Q2ANWFAheC1xUNkT8e3V+Lsa/Dn33ljiT/8MdZm2BUPAdvmQWdc4ybiM6ByR
/EgfX7Ro4W0/L2sDOuWolU4OX2DIQnuus7hc3mSY3PQzASHFYTgI9D/vpA4KBCM2
G0+NnHn2NTBm/GZn8VIQcogUPnF/qQfs/HCCFSMQ6d0xnaEntCfuToUdjmMVBijg
f8Mh1yxylpQZEQ9FpMohgMqJkIWkZZMdNCN0NezHkMV132PhsBMRFnrKNFsNdpCA
RjvNe4C+uDf4aVf1A9t+c69fza48Rn+GY1nwuwO1HB9GVeArATdW2wJnLZfM8yiS
c0zppLtoSfN781enXwMEZRw9ULCacE44on0cam4HEp8QOK3myA+mDtaBX71leAsF
TR7t+7pi2K+LEOXUwACAxu0X0r8mzb6LlOCGssgVFcupzXJ+4YZKkJe/eHltOD9L
MzHmlT2s5g46CKzxMN31WDVV/VB40RC1qi3A/SWlzH3LaPJEyG3TFkee1zjh8WHr
vJ0JKukuZAen3Wm86bfNbRJoA6Px/dKBmNDQ/BBmhiKMWwredsTcS8TU+84BKSwG
VoGbeF6jhGYXvaSXLrbnmtvLuYi329yzAkphz52EwIQu6NEJUDBoKkKnFCp/PwfZ
9PtXxi7Py1yVECLOSk6Dy89bHSmSOiRwZU+beA+Gko8Mi58aXrY3nNFCyedFY4iL
SfjRS1Oe4xOuvytX4F/Pgm6e4F0YM0dbaupJYf9XFLIkvUI49gTolZ3emz9hmgjD
flJOA5rabyE19noTXHGPWOyyq5ycAMOHjnQq+WCyffEHy/Bbjhx8YTrJ+0SiLgeN
F9Fp7XM6pIrCl3o+xNYds8S/a3L/z9BfOi6znQ9u2raVcv3jAN7EOv2vsltG/KNK
a5dZ/2V7uvBtIC3BGyDE4K2aeysxr6snVYMy1dePYTVR70BVS0OXtj+UfKTMNyh1
7WjK24hjCFh4fNtisJD9Mc7a8oRpj67QTiJrVntVEmevwdAz0NEnbMtr/sRxO1pK
kH5oUh9OratOAxULNApwxGvpsXiLdPqDPhM/y0abSt+P+NINd6Evaorz5pd5DgPm
mFlK+Il1TRtEiqauGre6qxltply1XFCnaTX/sSlgBjXaN841CKUfh+IBEB7+d+OI
twNiEtJRJ2SNtrmJ1eY0nRPq1gfuu6X+ekvaWCLgxkld6FQYbFArRSornZg42aA4
CZHyeHWFCONvrLmiBr9E+G1r64IGzOEsqHYwaztWsKCqZV/LuswuzQlIwFUNUT70
j6U5DZAXnknjKiw1sEd+78VzXs8BG1UOZ1l3viHVOV9VDHDIgdBeCbEVnDvZ0WkZ
d0LVToSeZ6hw2r2KhsRG4cLHlHuOpDpuVoYJ1KyH/V3twFrw0R2MPAZaWgCHue0J
nBqFb/D42yJEJ0WG5cKMdhaHmil515iNk0GEFDsG9ESaKtXHLYBoUEpHA5nK9Cpj
F4QZDRlT6u33koLshfRjFtF0tVzEhXYaHpQkI5E8UlOF6RBiRfdc+GgfDQQBQ+sA
h9O8dTHMp9xeOjLXRizvyLzaitiic+cwaK2qugaBIkQAvl3nZbVSSpaYHJyuBIky
OgsY0Ie80/6B06d3eNGqvx5wjQo0Odx9Mq7vAc6fUKstG018RAvS4Rg3uhTie26u
DKAQO1YTEL6eYcOH8ncZPruF5jhtCUSxS7AJ2ePVr9cCLYPui9UCTIhyWT/GiQNk
oC0qwBGdRWy/FIyXVCZ1nzwsK20hGEiRBt/tnmtH06wVXghNo40JffK4vj5KP2OA
7rqswCdaUGGz0UuBHKSMIZapGk0t9E7mhswmC5z59nh/ZSrKKQc2Hpdlv1HXpWR8
qsYOV4VPAwjD9ZB9h4opUNKKR+xM8YJqL8zIx3kaYDg5oaOAXGOG6hbbpKxTCWM5
5SDmkfAD8180lzO3Tlnd4n8xY/ZAmZw7qGXI6QIaS8Nf2VD2wwLBj68HeuxTyVG+
0xwj+Gpaj5iXKvrdII9eV5KlhLKdd/f2PE5uL1P/p5uWI+N9mxNZ/e0uhJXmGyi7
sblysfUd4qSAEXo8VnoC+sQDu9XVqlP29ySMYv6/1biA0VqWEHuphEJ5wu4JOu2N
f4PdajFnh2Wif80Tzv2rP8hnM0fih0+scN3YaAfLiEkdqzleBHBgEFQjjF44GEs7
q0ag9GQCwaQIwGmN2+JNvylyStUTtJZugaonbfwciQH6lKTNuU4xYDFyw3FemA4a
QSD6Ce+Nsp/moib8KxMJT0NTipYUAodAzKZtAcjAJLW63W+AGckTsSQxPo6MRaZb
AkuNfSyEtaTXwsgZenkSdVRR24bU7kmTI2OyBeB0c+E7MryM4KCN8gpZSjcF2UuL
WtZtewdgFr5Ay0ji/vLerThLAiI3rlBYbO+PWJMLPb+kwo2dFidlTjMmNfH7b9Ic
ppJqeN+i5XK5SnCi+YRaQLBRpa0CNuSAxt5Z1S4mt+355yj70iWd3var7kE3qGjI
E5GkKt0TjoK+z/IydbDuESSAdYob2ff+X3dpZ35eMkv9F0bIWY0LzQg0m9Sz6D0m
GnnBmOh2GEqorf4h77GNYZOLuOrwrrPMqgBMUmtmfjsy2hIRfC1qJg/ADnIQ3Ecc
YAwe3MdA70Yp6MjMRZKHxIBmEfcasDacSwuBrMxNZtYO7xfVkq+6+BH0aUT04Nsw
apvj19ryIloVV6BZ9PuvFwJ9x8Ow8eSiVcNe1IqE7GVJYXzYxRBkS6YKoKH8VxgL
e49ZuYXoidT1OnVgsPzQjmDtjfzpGnZwRxe9iQ/6szAE48C5OpmKh2eZ5ENhwmuC
n8/jeheQvPlAZS0jLVqZNZgUx2IUnj6EyyHNXxPGg79kHUSC4HSE9d7rhk/PpvnD
oztpzteiwKDJvibtzNNjvOtRe4cQ+Xx37qf2HRs8kwQgnEDAtFqII5A+dZPDKiIC
rruPl6JRYTvkmuuwCK/RNitQX2BB2mroIjutsxMvERzhdpRROPAzzi/d7TFAFZxM
qrucV5pX+fTzyrURmv/qoX82hJ3HMbq43VJzMZM6dEUljBkMlsze5Om1xIme2pot
ZP5T6RmE9yncANd/8nWVAz78LW2Oi50vtqyjUkllR74cPOJwGAA5g2R4Q0jYHVb6
MYYfN2K/FEXug80q3K9FxzvonqLGqxtr/KIu+kft4t7WXeSWwMHDil+DX2OZHjKd
INDQY9rawCRRXCX+jGZUOPgVn8r6DzrNiP/+TV/e80cEidINZrphA6u5XfzQKxg4
Ms07jAXSIOdG7eyaFEYVxe2NSLfhjBA6UKmFxl99lRXulyDeKtQlcQvORYlTxoLf
7MizIHBDYEF4yQrjY4WUWGmQbVelIA/VRYZt1O8cnhh1XjFjOMGPLgCH2SQCHti4
+am/a8YA8bVzor5cfrrTqOexBqb+sxDP3w61k5uO71zhbHT2TE+WUgBp/KIHDGX3
eiHwD3IC5Iy3suJK5UTgZIamc/JUW0LJuSZfqdG/NBTJe5vZ3GfU/iEpcvKtFNho
OPNDNLCKcj+Uu3t9jDBJD9Zy0bHpU2xLep1OQIid9uz6TvfddZsZfXja9FrOKEJP
OmdZXdAVd6a0QxG26uiBFbyskWG/pt7YcUgn00/7dCx1lYTUFBvlXmCrwnsSf6ww
TgCUkkCNo8qVve5k8fK5CryPIJaSWbiLWi5pCrr8CgQ0Ae8ZXXZSKwJEDyCSWebx
4LV1BBEL7OqKFnK9zUxHgH+cA/QaNP/7GzZaHO5qRMYMGvlElqt8EwJ/lXQlOUOd
MXn2/CjtipsOz4bNvdbHf+fkdiHkkY2N3BEo1ucpJdNJ5EkjNQcNp0msY0ci/pXt
mkr89Oah1ICluxMsVzyYhZ5Xv+TXjhOuzvZDqBumRCl+E9UC4G+8MTGUlxFg0YRA
uOC6PKn32XJB1AgQ+8y3vtZe83mrAoN7N0KWarjE1Q38Az2+O6DKGW8uOHsiACy7
h0NWJmQwVM50jNUDTZRQbSxyfQo/Ps8WFSei1pWogB9IIf6D9mYyuzslMTF4rolZ
rDhJIUa2BSnvlnbkISPN5Wa4AQRjzgzuZ04GTdqMO64J568Mjmumb7Q08iNZlzr8
sOgwy5VvozKpsW6LIO3G0YnZT+xwp+Ltpw2cxpiPQrptaCxxeKW/TAQ3GCxKcxYB
H8GhuMb2VysGowsvMbnfzgFMDoCjEW+tX54J6NWVuB2ZPQfoCuWnryw8lHMSOy+z
Bc2Sf/LdIE/jiz1zr3WxpqNcOlRokFqa2v4asqOhfxcF6wI4n2pIpKbBo1BQL1Dj
9HTGhT9IcaTlDfWFrTuinL2DJGnjNSVhc156NbJUGeVaHK8VJHqWf8l9dopNPxVK
oGdP/XAxQNvC+GezrYB1nfcOfaYhuNLSBAubLpAslGdAIzyPL+vnjlVN/I5So/Ml
xkJ7gVzW2VyUgXwMXr00LTcLz/NGr2PXirAfOJ7Q38Q5AOt4254XdI9lsvuy8mEN
ec4JRzdXZxB4tgIMAmBepi76WuWQQ82dAJJhlhq5lQT+3LgU7ZPLsL9zKPIZ84EK
dNsFpFWX7lUC5MKzoKLAJigdTQvvfqTmmX7VPYc38MiB92SweLsD1gJzNyWP2PsW
5wppJaPviJAolLgv/vSOg7qxC+Ai8OTMD9nL7YvLchOZdEH0yyPHIPpYmAjM/cu8
gJz9528t6EQSaAnBAfEv1v4zXF4cerIchNad54ksp0PcMyZmtAlHCKPjcZsIz7AQ
NmUVlDIPVRkMMH7442WLVgSXO7V+g+AucRqP9XzL/IObude62st3n06+STPiQr8J
D81v++RfJZ3B1TfK1YlBT7mmEJ46BO1xyqh/Eh8Htv5Z8L9QmKYZ53xnA9i9Kx/B
Ey+0oglrj1XWeqOCihAbYeyW7P+satH/3U9O33n7/o4ORzmFPAVYt/+37VCIEdwO
FUNuRo/+dwOT1MTnMcYboWUF/mZ/ZCstHmY+LyDmV112HxVNYx2598blvE12V1Ss
tZ/uzrEN//qx6GlL4caEOyAtgz1ioMqSc+dtNm4BrS46YRTugREz6pxZ3XVXfuSk
ZscrjKUldCWKKnY5Zlz21vOEL/LjUXocIc8e1K+m0+p8ZcCKwUlFyFxZO8Zmgy1z
1L124Ho2/LqLhMWm9Ophwtx19v3R4JG+iXBFbbKZ3YkaSXnhTP9BZkz/mvDOgW5r
Cfj2q9UPwD6B88FhpK1TL/Fpn8OIXWTvj/NjaYfTRHSyGpemoW5Yv838d81aJ76M
hYDBiNtrXE1l60KA6dIIbaZ1qpjqArXutXCmvy29yw9SdyQ6V7zlhRH15KNs1fY0
9A2KTrVArUvYF4FiA+C2u7VtAMOwXRcsVOu6a5IcFzdvwkXdb7fbFaNn0R24bNi9
sFp7YnaxO7uWCBBmHJbqAJW4QSKZSfO/nGH+DauFWjFzulOc8rw2BIMH/Vt+ZJiK
HO7jncJ9lhmCkmKbrO44oxAzbOt3T0z9gHfdJvBjRnuHckif6DgIK1VqdDHVi4Uj
LWWJI8ukuAGHi7dsyFYnt39xDIKSuo+J37DfFE0LciQAUapuxe2VnWY6vcMyx8Ak
eIgIXXSjnSvSDux6s7zILQKTWLHWZ24p2wJvHi+ibi6NrvsOOyez3QdzKlbMUwoo
SycGo+TrT5oQ97qW/q7WTfd4u3V1FZnUqR5wwPk0697viOY55rUknSRAoQaPglaZ
+2Cnq05Zs7utu+dHmvNweH4ArwaO3nXkZzp3k0kr7y46iQtPmCM0tdUC0k2YaVbY
Uvq0SEmQehA7xSsl97EUumKo1t3mh7km8x2wt2fNScY/F1aSjsaS0D9O3Oorwejh
aUs+amZH6D8P7Y8RQIptWI0QhlE3r2te2yVwOKSL01eBbsWRNoNK0WTRw4f3es2w
B6w7N/oYb3a+fMyIyjhNzw8jZoZDFaYNbD1SAVYHWh47TjBTQ69QulNoLkgJ+zVH
BqlyhntfInr4kwQCjPc+Fo7vxl6fNSLvMqHHT0YH4BI8UZZnW1u9imNIRx9dIpDr
stMeb22lrMtuh5OrCXY3T4ZFeZm2MvhvueqxGay9Mst/ho6rqF82pzjODaN97beD
cH3N/1PFj9aTZyMPXHl+g+wS66YC+/I6X/dh6udXL+9B6YuFW/Dj2gqxcoKiwQyh
/c7oDQezRd8DvF6AQmw/LuehbjcYShZ25c3KJFMht/FF1pNBEY5TYBmZxXx+3zZZ
20Gx0EiVhpy6crf3ppYb769cj05IbFgV2o2q+eHZ5gcs6Mjz2HB5mhNCyQ7pt24p
YFZSK2pdgdMCqUJkUJXVoquAqz3NjFczy202oESZJL6qaALnhNjAso7QZhmGWcYE
tcEpXu3hG6lkgIl0F9OfyjH9scXbXEkh1BdgdvGeLa1gV76RrrxAI5+OS4I4EaUO
Pf6lHjLlJkPQH7P9j58joGRQUtQpbd//7S3JDjK+Cdp5062Mx+Rzrbk+V/AUSpkS
a0BxkUPvzzVWkAIUbNxJdycrs78w1RI69nedyvfL3X03hRYsovJx16o6xiMCbR/x
4bjy7WgwvFTQFOPUlrFzNVK7u+z8+6l6LiPu1SRsmGUhIqgF/7iAKeNqiLBSJ/aE
AR2GPiCcFVCiB7Ms21+KSZHN0RJOCiUzTaJVft8NqZ00SDlIb1ojJTxPvxBC/PW8
P5AUfkQzQPShdTY0IwepeF2nPj8AmjCgZAHwTHgBn3SV6wdPtlrf8ETJtz93JVE6
OoCgTcqNEJmmjUM9KoiNForTO0/DZU0AmXixLsKgzEGaozCEjJCir+TOVwCa3a6E
50kwkWcJO60+WB3L64+LraguKLbhMN6EwtTf2xSk6/xYPMCAIywVpwB3aKM9p2b/
6DA5Q1pRg+v4iJAcgljpM4Co5AJACe2zwQAM/5zJ725iKyNCwcR/0eO32XbHa87i
ie9YITwsur8cefPi7nyRdWI6WjZ87gSxpQoA2P5kIh2y0vrYxq1EkaA1Eoe5b9HO
LsZfysI4k03A5SjCVoYgZmhXYzqk4+AA/SGarMRXfy7BxZ6KuGfhmr2rD2BpAI6q
XAzwqfjZDhi6XbNUQILKEo+5WbcuAAXDgI4TVD0x1vNi9ue8Yh9XZgBtATbnkHxx
gT/MR7niHdT/fQZJbhWtG79ovNRBXP8VFaw4dy8I2BySFWLrWg6x0Z5tgpmdMuGZ
NYSCK06AqmQFxabVDetBarwjZ++/di/dY1jPrGjZRSugZW7GJfc878x4YHj4dQXS
40FX3JY+Ix6iG99+tkcdLh6FLn6F4/lDbVPEL6Rm4KgeyRdWOlsdGpcUFROhyrZd
DdQ1OttNIJYQsVJfAxGg/zhfOmv49EqUKbxPDRGqHDZxLyJxlrNMe8H4M+fqYiyP
0QdQOR5Haq0slTf60DNlU1N171G3GRmbE1ychsKb/J9u9/3fC1tfonzIaIfSVDh3
orYfebi/X9vAIpqXXJ6/WvSBGcaClA6dUEr/6luDEe8CoPQVKFvN73rrJ8kbuHE9
BwCXfQVS+J+HIs/IrKlIotrCZzMl9XAwB0FiSwf78Xcr0nof/GMx6Vg3M7yaIsIs
sa2FH6hqXUV0iPHODY56mYL/tNibYMNtolsow4OwpUuzx2XcS8lyTdmXQ2COKAxl
PiDXSfIGRl+ygBrVYBjS/HrLEJ70DiP3I5CF3UDxMWcGkeICz3356Tghldja9TsH
JPnGPffKRjI194rhRYSe0WvqWq3ics7iJ1hHu+5HHBmMhHAsQApsGbuqLa2HFvbh
Mjj8alMoQeksNdGATTw0eWRhpY4wp5lfMYHVnqhpq1lOW99Vy+ZoLRs2PXNTyJvF
bGqHnaL1YXiwW2+tF0qsxtqLknMwUrh4/1JT1WChedP+dmns+hig8o0rqUTkPskn
FydMIwNQ7Jm/SmBlOiFxZjD5qpw5ZpPnWvThXhguS/iwnuBhTHv0yk+FuxVxBe/W
6YsJMiPL0gaUqb1lNg9Qn/mv5JSMy/6uKi13Cs3zu/AJ18H7fAPWezuPNf0+DSNz
pTlh942ejZGJHuaO8TTXKaSw8c4ze0wP6fyChZxYRGFlfdlcNL29nAEjtCc5JAhU
HeLnTLpvdSPwO1bt/Z5DDYI8fiaWGn6VDQQhQDoegShTstLRSB2LM9ipqJFPI7Om
1uYRUMtmY+fPrL25tGed/+HzpWEPpkTRH34UQYLfyeVe4RT31Tr6SmvK4ENfcxtv
SesUU7+G8FNp1Wuhsno4JjHH/I0Uev9vT2lY2dS/z3KoPBYa9rOiQu1PTGZWYggQ
YfIuQuZfUJ0v+ZCUcbmAOkWNyfFEnWG/hdsNrzxB9vSVTq9RDx7r3eZ9aCEqXiH7
SGsqy8bS0ok8fUOdehRpM61ryJNBeGXy9iskCxpEeaDn8wmbWoBSAa4lb023SRxp
m3fv0qO/XMpgqyE8Fg5Gu1CRf11jmBBdDh6K3bq6uz8HGtilYpZY7MF0sLNMT1oW
VAhA55kfyEoBnZ8HlL2PnK+WRuCj4H33kSTwtVR53kbhmrJLymYxsh08H+g9dwCi
MIO49A93kqbrxcj2unJyNBau66wlAOPa0/QwPu/EQuMnunTnkB9g9LEbXKHl41uI
6SWhTc0e9++BllKVWZAlo8MfRbnrbHdnd4kZ8aFf3spULBqucI71nsSf289M51Da
TBBV686vqPp1oRf7Fef77IO1BQC1cSHHs3VDFtdlEJ2R3HExYJUUetVmtxr+4WhQ
lRrpLfL8SYO5EwTWdxv073erFObYKZEet65HKKFwvIqTmv5Fur+YIV6TMLK+30NX
elB3wbfN6hw91rP9a1aY2VJEtGgmQt8ByphS0ZysQiywk/MWcnnPRRO+JUOimw7s
4sfgPY9tOdIvLRbyah7mlmOrgPch/J5lb7Q9Cks4jPAH+iOFeQ7mq8tgm86c9j/Z
k7tn7PyrwCgCN6heMcjREUc3haQdCXtqvQuA6Ct4FeTUPIc/g1DCUcK71qF6sPbK
iBbvExNWVI0toOWet97E2vIbfbx4rQBn2yERKbPBdUXyBRNZ7OOTAfzCsSCHjch8
DF5ccV8tInTJLRZQVLfNMFS04Rlx05Jqohjj9kjNwHoxX6w5aRQc9fV4k/966xzL
SEqCiFfciBPVFoV9Pd2lNpdQYNT6mgBpeWc45Ex7KdNnIsLXVhwSB9hnyIFZ014W
7dZVDFP3rlZ3eaqrJhwsD6KEFRTQ/Q0KNDNvH1dxzzidDyYPyaYoExi5zyIcEqcB
X985NiEk3OzfBDBklkLkFRMXBABsf4onyZHbcOE7z4ntz8RKcTCr7doiJc2GiaJq
NEIr+z4Fkj2ZEm5SyO8H1x0isaTY9s5otGJiLXmEXmOThavgdVBtPdn4BAHgSw5F
bzJU57cRT8eL3yEZ0EzNtxcmaxtXyfloE1VUKxjmnb/MmoYQN9L2emuHvoM0r7ml
llVUgFpoBCZFiNH3jwF2FVMPdUyFKF1z5FMoZda0vSP9kmVn2ww6HXcn6L+Z/Qkf
qwHnn3qRtXlc2OOwjkqT2zmaBGePXPA3R9M3/OBEMqswV82oRI0sJzS6l4dyHAR/
lAga985Dv+00l3rfIDycyL4UotZSkhsf6RONH2/WKULcrFIl54W0FF347q7U33Od
5XLaKbwI7lf2/4L5lJOuVemR9d7Vtnqo2fPnN13YI9xcOUCS9u/nFcBkr0o4f2xx
I6kEP+YSsEyR8on5CC1vHnxPRAvr9bu7ifgjGsvgTJCD4s23ePFdIH0HgsZKh1VU
Q6uscAXpTto1lCZyybQeRYKOke/PPH6WIr0jJ8IL/Re7VoK4of4SLjwOnL8P6YMh
8mWULAg9qyoF/xb4YnSFB1sMhjeBGhnQ7jBFIDOs6ILMJxXQeRMBgVQWpW8bm60b
YB1hzaGivI/+F7ej3kYatGE93OqFK2gF0Y4+7CcHhQx0J2Ib4a61QfhNa4N+CUU/
UfyRWpMR6VIjtAmOAmmy3hRBsg93Z0k+Q55zX+XXKGpjMW0ZfOI0eOGspcQIIr/w
g/+LazZza+hXBs5ScxeIxR/mieZyvlrpzOMDoZaNVg56tsD2jgqpZy5KNlH4ERiI
2RB0jW2uLRDNFyy+edrf2Gp8ppNinks19uRuCl598EX+L0LpSBjqisYeCHCJBzyH
M/d7pFqc2FAJxfSMocXe+yZ4MbUa82ahugxkx+/lFvRubKFJ4kKWuYF7Ur/dVyVa
asaF7T7IkupBlO+eP7Kv55EVwQTZyEIvWenb0xl/3LVcCii8mrS7ic43NWkJ5POe
VTAaJu6Kv1dcTnwbux5q40zzXV2gEWDBu46UeGR0K6d/srv1oGjaQnG8VLYTW0dz
Lyrg0DBmLwo0CGTuy3nOPSJZNtb0FsWtm8sVi49be2l/1p/fPAj0Hfm8QqHz4UmV
7tAvXD+BArl/ExcJsirgXl85dB2+NImReBOX3EecWbAbMmgMxl3sJ5g4eByb7zxS
wo8OU1qOMPG6TIpRVX8cP6HTPGL0EvgGLtxDoZMLc/KnMLCXXFS1fZ2GJ9NufLbL
DOWr9isWV/G/hbX+Ivngt5vz1KAN2cONU4VMvBw4tGPJvLyKfPbj0N2TZJXbHwkN
5oVnm47vIUbrIfvFfZeHrkGzgL9Wr+TljyXd3o74ONeuPNe0Q8qvDQX/LdefRiY+
7FVjNvPcI2H2lzZlUzfF7xvN6bJFkjdzBdBjJAPxVrzkcXpGbT83bL4/XVchALIo
FPTjKvp6Sm08ab/kvcOFVOtxOxptaLgn4X+ZqvczzMLbLKJo8lrZ0B7owWGjQMd+
8FVOv85Jf1F3/9tsoSAsIs12FBatIGVVcxgQ/dJHrOVFmMLDfh6Dy8yL/1Zwh/LA
NnNl0vTRm2KxJrJjEAVRNS41NaEddYCdx4afhRyTB7fc0oRQqqG/ylzBpC84I069
Eo+QqQr+1rFyq2aj1LdYeZINPMDcPJV17OfwpsG5l0Gwgkw2t+vz8UkQNz3MvV1s
M+mSqhoUPDYB8pOVhET3gTuNBzFxeByf7ERpitDNWOyUzVD3gDGhT44BNJgXj15V
w7op116dEphL0D1IW6XdBfqMMrBualWJXiCChNg8mgH0k+agrlDP14e+gACnWxsj
niTN1AAJElIj+USDshIJcz4Fe18gXr849+VNPbjFLlqons+3K0TOzz4tAqhlOd4N
ZFClVI/ImIesOPhXhdRFFt+YXuPKayAzidEwnF+iMlusenKs8ygkbcZdV9lgObJz
r0XcMh/A15/hodEHRR3vavEwK/GtpMsTFsfTs5We68mcsWNKBKYunYLM1w76e3MN
uydGUMEp2AKbZ3Qd6vdN0F+tXPucb7hDg7I0hup2SkxaTij90ItS4WZky2ULkLRC
9Nkr7x0YiWWROUXTdekl9mN+phULUygNtIRjSYaQX0KBzrFsz+YTJJnZHg5TjF/Q
hMzL6MU6oZ3pqoga2D0lnLOmJnWlOJADOf9zdjld2JJYIdYBdrZPc9nylDXLyLKU
eavgcHULQXPJweM3dmUnRL1qkTjU4ei/Tx9Z/vayc0mocLbH9+oLC+Y/a2r1kYps
V46DQkrhc0o+NILpbCm/oJzZ+Obpw8NK9Coh3WhPlPjXRXFkb5IyPpGx85TX1Sop
xtQ5uPMfroEsh56zwub0/w3W2ReH15mkAI/S2Wr62dRjxcEElf3xRSQfH/gi8r0G
CB6rKZTHEcppAwPEM3W6HVm+GtWLt9rhksCf4AZEwBTEXMfibO+eXSobmkT9myuJ
D4QV97jUDE020pDcgimtryJemEGnFKoVge4ggaoURrCAHXSnsfJ72Y6H6MIAQrD+
5d0Gaakn0Z0g3SaOBMpDdMVHopaYo8wdlNf1dSR8HYBwADUiPFuP0LuIhFNPQFtt
Ahy+K7yMKWJmv2q1fcavsdYQ+CcU0t2tTuFIvu/VRCti23kWQMKP4QUSnpJ2rACn
LYlJ4HPlFFH4wOSh9CI/E4gPk1mkhNXUW/4cXfkVFPv0lOVaLTBZmiF8jBnyx2UN
9mPkcB5evGLR3l4LMkUWQCr8PcVPHkdQz8jpyyLIlFnvctALA7uSXXOHAkW1Bb53
s7nXtfPGnzfw3LLdbHiJg0FxXfT7h6Lhn9XigcodPD6QXRajI8P1txvke8NF671y
rwAh3NukSwGE9Cux8//JYc1ikefy3FIhlx7K2Lz823Hc3OGIeuiyrkIrKdJyTJwy
qNIwg+55cyQMOb+dd7I5cG3BH+eSw9SIVdY9OIjVWqYRxr+8HBwLYJqiW9OD802B
qH9eBJmRHUcSVMzR2sK3DLxBdxyI27GJY6YvC9hcUtLeb68YbZNdWKt2bDLc6Wn/
A6zfNNypB2p53Ighy5V/nSZEmsivf+vmNIrN6wWaUR0gtYiJvAGXi44jvY4K3g0E
4ZyUKlS0NDN4vP37I3bMUjcnDr5fPxouacrUoa54iiHxhJfU6QGO3YlUOEsnUcUG
j1m/ltSPZLpsbhgtGHR3RMoXpdcRzpnPXvrIWpDi8SIWrm0xSaEtiyIZ4CzcUilH
c+b7GCN2MKqgzelqmWitI+lqgO8FO9/Qas8GDQ8gEMqGOW7FgbLJA2ZLZgUMrD6n
EeOtBW556qNw+VP5EitFb4fZRIFcavSLAyZNZGxVOtsEbe+cQo9WDTna3pD7ggPJ
BcqSBWCAaNFWzrxjiPZknv8zKgwsgGWvCTS+iQOaoSCNUx4DDqnRNyrUn1uWWu0h
1w25nTWglBJ2UIfMTkHRray24e5771yp+Pyam9Mwk9IDKPF4krsbnPXlQu+4zPV6
mo4Wz8Zu/pguV8G695gBpihMVD56hl2Z+cemZdo2Cc4d2nnIcpJ/Os2IUbl6GgXF
/gCD4k1tfdiomKjse0m74Yemm6HbUuoaucj3BPUSMwWiJFZn1rtzvbiK6/q9Af0f
FuEwrXKM6osIut8Ih8oSh6wnRjB/vFnN6UxGAKcfFbb+K5xrd8yIdwUgiZxoPiMr
4kVoK2mdI5gPM8MHEUMcnCNDluVs2wICKlqW++OxIiyU0XgcUxF9VfbxQ8DcsDcN
44oCeGFQSOjiri2lEsYiHstOw55BqkLg1gAn7LOigqz+RGJT9eaj88t2yuS5mxhs
DyhT/+y4Mpszj7dewEJBFaSkknrGDoF3VzLaUTv15Ebf8yy1wPQUj7+NSZulaRVM
BNGFo3VFX+12lxHhN4MQ62BY+K+OVHQPJI5SodZDDvk9P+18y7qYv95MsZlptCAk
7ODZ0Gv3P/cJ6LdrH9b82S+RWuipBCHLmI1SD3m8qS6ZmVvfoYE2gXKEcPZGKg+/
506JPps3R/7lt6v+iSpV9cXxRtsXG5qpsBUBR8Eu7Tz55lFsCK8RoyAfG0DyyPna
iuD6CHrf0odpDzq0hSUsL81iovjEcJE0DVIGfSJDSnxRH/NmglGRVYHHkwMScI86
cjTEr6AjeK7X05QZ/FxeURMj7ItiPkIx+dc9Ixs+IkFwBqn5LqG2qg7DDuhMRDxB
lqOyKaRITH4vsAf63sYr0rzOnp3jwJdmPfhA6UJ4ZS7C3JUtHgk/FP32FI7JBNxb
2vkH8dzdFYMskiB09deZvS1p/0iKGtT/HDzOX48k/yo6HIZ/aMdSQZwpbLk0QQGY
V2qHAFFsMLLWZgH0u6/SRXBTJKaIQoKOIpL1gIGvidXF6o0OrvfqNfdF3nhiCTlx
1GmjUx2RifGAZlp3+pF0HtEvRkj2HNHTpTTcU/7spWo+hw88kKkPNlBkMJ71X999
rszv2algiTABzt0WHuUELCRRJeuZ0dAXboJdiWStJlQvRwwHW9wBkuztfiSs2mr3
6k3qn0tw1uYgpnGVxjtzGQaZXeqryWpZzIA7mzRqruFd0fSxccdVeWhRZpZhoafX
jNouS/MfzVB8CwXpgtJzNvfF8sDqu8uQupY9eJkvjUTyCZU1oxNQynChBT4BAcZf
g1lAWvIIjcoSGyyRhcZelrFgBPSe6PE4KUmKvaK8cQyeFI+aJ1Dc1bf7B4H7qTVe
jm8E5/9ZPPE59hO2gjRscfa7XiDArPqAEj5O6qvCo5tKVrUyHnj8Uaclh93WBJ1Y
ZP5MJEMM7NYwkC62cdI8PF42T2wTV3UnmKAR8onkixC8/re74cMAsM1VgDh+7j5T
+O83gC5Gce6vYO0LJnMvkrNf5yS0caChvSPJa/KihKyqh0HGXdCFbBAw9X6jIb+s
xgrkG0I8b/21stWZINzvNpq6QM/L9A46/RxjHWD7a4sa5NQeXNPuetCEbu0UYiTi
nRM5Qll0KCGBIs8KDc/GhikPNsWqrb049BhB8xMfHHbvCL84yeroEQynvczH6ign
YJ/aR00008CL/HUmv36MDhNLEnv1a02KucHfN5wC9503RcnSgDW15E71LW0ImmLR
KkcSsEQdnjLXYbBoi3H1bC4uaQphGgaS3nPKE9BvDxnk5z37949xghXBMKDBy4Yt
PhmZB3V99pKyC9bgLLG2nxDt9OkXyneZGAW/i2sqwRjWPu3tKubha6ViNn6gU07X
HKBhb8KQkFlcdVxWaf7A4RJdKP8uBrn3TBLTerbPM699vGE3PVYqOu3dTlLFm79X
hpCtvYgc+szLCprYwR6AgLoqxa/EFzrNY+o/clYkc0+9ecBx9u01EcKgi7Jg4T5B
h2oizC6GoY4+ybmzBfkCzK8cfRqU3XBV9OexKHq2Rchs5io7XeDvSUSP35PU4yNQ
4lD6rYvX39Bva3zl84O9EBRBcCiC4CDMK3omokhxgo8KvEJLJseOj/l6UH/zGrH6
X3OGBF9k26ELgr0iYiRBXFo/U+mAlFto+HZPQQs4I2QxeIOET8tpLHkUBw3PLRAM
bcYfUHOddOZC58+D+NZYcEw4t9crNHOWZBdOnM5fKZqYW+nw7gmW4ZQhvnCF/ajm
Sz+9uXSuaeo0tL4QvH4EhCZGdS/hIhjNYqmCSYTcppycIhLZHF+x2ThL16TqSjqw
Wj+7UNNGm8/91GT71Ab85MC28sClUMvAH40xwy6g/5I1xet6L9sr8zKPZITC0Nkv
PISabZnCnGldAWEWjBEOcm7Podpass2Wwngw2bbA66IuUJokEtw257BrfpJY1rLx
r4VrAEq+1GFPlWNZh5BXUcz+MLwA8f4hY/nT0zgW9o072i+XP4pTZT0EIm8klqst
0nVusi8Q/Fxi9BwgoWregKjhrF8D01LoFl9ih2KVThzRjCcqS7kZqpS2m0y3oTbG
`protect END_PROTECTED
