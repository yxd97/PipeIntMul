`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pF0QoGdlHjRAz48YaxNP9bMITsxUo5gLv9EX6HUxlveoiYps9oCFJBpl2mtXXljh
lCExzZYL06gy31awChYOYRiA4Ibqeeepqxe3kopIWtfNC3MuwkRx23yS4M8UPmr6
4vxA2Q5H3HMkEPUEH8FcZ6eleC03+ijoGHqDIFrNbEfH0bw9xqqZO4VRHlzcGQCR
MCykbMTc/GFK1FCwKLaqh1KnIEd3z/zTfPcnv8qDPmO95OPlJuhprgSLRi1YgGB2
q+0HZG8s2Wd4H4u0XBfOLdCo/QoFBGaN+vip48mdwf4s95l6IvzPyiHpMe1Z4Rbk
FD5/fQKUjUscyXOe7dXiGupPmRjvK9NGV34Yfv2YSH34lIbroyoa1qj4PECpBrcS
ojLP++Z86zAWLmP2ihcAT4kqQhvQu6yIl3+AN8C3EqF09TsnqwuXdTEJTjSeyPTW
gtHpC/WP9clQT3w8fFbz9PnQ4szmES3T7NILjlu56S4P2TCPgkk26bAnMiRhOP3u
fPN8ZQzjr7OQ8JIlYpsKPgh1aIDqzdilEK/5ctxpDNC0UEh1VDcnmLHBOjKdWY1Z
DaBu3XKtkuCHpL5FJGM0I9EJiw8jStVzAKZ582H1+aYvZkGEiPC+PHmeSLQBaOZw
C+ilc3u1+pxTTM5nSIr+ndnANB+WejxyE17h0lATBqxp2pmi8jMI7H9ofsyPyjlG
VEHDj2/6Og5pLcaNuiVWvVH7npxW/AFRFsEKEgLCMu47CAz8IBrT7Dj7dtiXgu31
PejY/HaGbW+83z6N9hQxoI6HWx2+gVhD/14s6bV1eKfvXWPJ1fynVHKvp5zTlWEK
H488ZgJbOso3uq8Sb6urbyXA06igIInxgMSO3k2ym7Yplpcow/Uj5HWPCQbS3uI/
rMxFC1oPA6ZDlTA1oC4U13XB53mJpIivzIEaf8dTe6WWmD+3Dsv5sA5ZmPkkXQTx
m75VMOKd/CHFv/X6rhYbojktVy33W/jw+FaY4CdDDUmFFlLbmryrsAECcQhwnkyZ
OuUiErpynTWnvCFgI1Y4rKz20bal0cmRHZGkVPynr1VlJtOK/rxlTMxjt+KA41ov
/bnrsfZ5EsFu7G6WafiGwIs2OKRe2Xy8+PHF2w/he21KWhENzhyylrAm7E3PhMjU
Y1ceIIUkhw5knqXs5jQQmQPqukx45P+fLIT9mJIFBUUPJOYOjk8NkGih5gs/ECIK
2iu4YzZ7EUHyMGrQziFN41hgvTlJDxrhJ0S0sTQs1iew1ZpLE7mlg+61oCfTesXq
69bOPq0ury4jv/SmwVdijHK0ZMQf5uwz59Oddvea923bu8IZpvmzwCKdNTQ0bEve
w/y+Sbqysw7N4dSwcBx+h6gnlkjz0yFU9PcyCFYbo6VhAIZS0jHBpMj88OcBfNCH
b/EGJoR8FCfoT1lFlFdUUPW4zGNG1/BLSG5BBHejzfHTnKyxd5QzvCL/4OyeVH5A
FADVFOUXufeCRpPdfEBa0UFjs0gZIbZU8URRcTF7iAIO04JK/xvJiph6o1mCwgBW
ihS9V8DbITgG3DTATojc890btPGihsVkNgsPCuKn9rwhVzgyM1R+XQspnCpXemQO
0BfGsyfAE1sfCgQO7jUKNljogsGFbBcyI6nYydvypjfEVBfagLFMgU8Fq1eTVh0Q
/Ln5zgKpfIFhHRwqwlHHqXTORh898O3kJePK9b2HZqZV7yAwE4YrtYVqi5SEh7Dd
SkqoxsUkpthOra59ucrviqYf0UZgMaOJtA/gfaUmUtjlOWdhhccwo/r6jl1WFkmM
7kB34oNSWCXUznJigL6P1v2p9zghmrCI0ezxahXoLXzeGPHsxNEMKubaMNcoCNtK
afIdeh8rzWN/u4lnPQcRP1mYf4DsMGrjCzWNKZL9sfJyOIIwoRKyUy11LAY+pbEj
JhVs+h1s9NFhRpbcJSNzgGLcvZprhkN4ekZbtQ+Ib82a8/FNqZX2ArTdpr8EQeXQ
iOaDP/lmjV6ULXITNemgZ65WVgGxagdo8lwcwgBGtmtB3VoYXASC4jO6d/l/sf5L
k4qD7eMjt1f+SAbsOauplGySw3q4KFSUlMIzxnPJEbqfvU+4eYPHed9/mCaEivbh
mJtbRTYV/R4Ub++qXdNsHKlc399/d/2OTu/fHDDyogmqxPaTXdkz7r6SH5/XaF5J
m2g837H7e14o16Ygfkf0zGUdEXzXpx/ZLet03aswzC/dDVIN4dLwCaO9lgrDC5+z
6vov7z/AAWK2O7bJGGUo87bLQ32xfA8Cv4ezAjH30YYOxrbSWDN11mtN0gL16sq1
EYssQlZdwa776nnycMB5sjiQfyljGSe4w7GvVEPHfgXPVFvwA/nJcNdHf7vo4j5i
JdNFpW+XvzPxkEr2SOjdAnt8v43zkOQWRkj4v+ny7W2u8mUH1wgF5HoqWiEDPKjS
+p9+osrIUJ0Yj6bXCnzsBz+d2XUIQCH+M04TguyiTvTSq1qwQ6cgjJIHmy0JsSg0
n/gIYUdO9wcSJLN9bhcuFDDtcEiepmiRIqh6BAHnIByd0Inu5uWmsKVEhchgoVW+
JOJY9bsZYCU5bO6UiN4Rl2hkn3dB1nv0RvDj54sFNNss5ZLX74dzzdKZStDH9ekU
1x49lCMz1knUBF+oH9Tj5o+oD0ZoUGa65ieO+IDlfC6Av93jVx79nRFdeXgqZ1lu
dbP8ZmtgHrpg4GGOwxhV++4gyazqstT7x14iog4GucrQvGT3G1nprX0g81rZ3pix
uE3/DN+KvbdhzEygTIq8rC5W8aUTB7v/4UFAFRzYT3vLmChCUAu5jmsnm555jnvi
cX1r0a4YmklbNenddQS3A8bGpyiERjpwmBYQddBhJ9IM3eAsNUdLrY5LEDqMM8Zo
fQMHvm2c4V7wCCdPB3IHBmysMLAPLXZFDi1AEMH+QIBUk78IVoZGLNO34lYecuSg
pn7eSAgwr+6Jh65grJWLw8fNPbRQCmPOOQO5FVBPxfpMRFNyM4eXvPrB4XHl1yX3
Ne39/wGBd6ci1hbjE3xreosFg6d+VWcd8Lmulf/2Bhrpy1JRecBYrSowvJLjgatp
5Kj9CaFzGNEEhISJ32ToM5/BxZTQlLd1nMRWvg3fk8xyH0HFRG+4EFxW/EKNnPHc
syQjBwybF01kcC4GFHP/LL2Ehosa10e27kDJWK/IdQioXdCpswkwSdTabmKMPllM
RVgiCyUFV5mCkBruk/h2Ql1eqnx1j5vGgIb1N3dScXyrsTAoQ/ZN5CDKhtTAtMu/
PQkiglNTpAQWu7dyZgTqeq/RgfF49lzDEf2AfciijPsJiHhe0i6TG1wWl5+RvcWn
54YlMJMEfr5fQN0Ol1FpRUsOhw3mEdKiqqItSfGMZVpc+5qFuuZ04fsE1aY8HWW1
LNIHFnt8ZFAR606P6jLOTojDkd6EAeURFekeuW5O7hM6DjGH0f8/4kct+O33xvXm
cN5V9qI/W3vAri9+r9X28dnCXlvWHY4DoqiJ2GHFXWmg6QGcDC0dvyc3P1Ji+SaW
aSZz2YqEozwOaRMapy0SuHS8bpcuvfoMtXcJcPiuKNS3mgjULZQt+PMKvX/ct/BP
nAU9lzjU8dDCA4Xg1IDiRjSLTY+hr2o/t+1/MhQXNYrRNWYdCOFvv3U1aXuXtcoy
/4FXuXuGpC3fFzY76eEom74xDCV3YGvO/wsaq0y2K+9XEOrZjCCOOtSldW67uSZ6
PCZdMvdXpaovKBzZg+rlsFZZP1vqrV+cKz8feYUZXR2kOoM0TGI7wC1ckbu6zW1a
/oH55m7fDNMiGQ3z4MSV6NErPTbgkT3zkvXiNKVYvdTXcIOHb9VSYNkaohv4xgfX
zhruP0LD8a7gEFSBo//YyCRWVGGbgttPE0YncK5A5O+wx91oI7YDKrIOgB62cYGP
cbSemxHoXM8Zh3+BSTQvUVUGT1/LxU2GEzj6z4MaXfGQWmYU3BmnJh1QckrtP+/0
0LRSU2maAUzpcIal1XQF4/JiNglMDmTrUVSFdcZWdibc0NN6Dfga9/ZS1xKnxbeV
IcyiFRHY19+AiYZsXZdY9/wGa1SiMuzfvkYm4KUQX3iqf5gJLyl5eFYRbjPcCuA8
cIqYPfp9gD1bMtMnOwlgOD0rxIwggGY4vuYYveWoTrbv/ubD6Nq6mMYWj8AiNT5x
3EJOwm8UoHJK35tUKsvmr4uGK+5EEYLYCVnSHX/qPGQtR6oQZFZuaBSioBqNeSKR
31qLyddivIz4xkIHyrmWRyIuADY5q0XYjhx4MXeiaEK/645t4rZ6QDQjf/qHvK47
yj9HZ4VLaFIz3292Ykv6T0Ipy4jf1aK5oD7TEd3FcLAgS+4zhzyAtfFFr1RmeWfQ
uI+Im7pdDjeRu5fUm1fovir1ihrEn12iLBzU9kWW3IblhEW6g7q7hh/uuV81YYFu
ktijW+xFY1mdBK5QkYIr0or/XdVQqPbHfQJ9Tv4gcn27Rb1ZGRKCvYCiyOR5kcmz
00UJD98nawIn5QVBfS+bEwT+M6EsvwKXwlPBH7GQEqprYU8SKbZUbP8eHTpINDG4
IZ/gfXCCoaDMBUKTlocxeacnIvAOZaNyRlNXfzrpKEC3nLPEzhjhkXeJLv7bTp9t
WQte6IcCPTe0PM5W3lsG4nQjRR5GhbbeI4XgBa/f9UfGK5Xgfu/qVh0axSzwDO2N
Otz2ytWtt1CVOVbtvcpLqMc7s776yYP2/IGTqI+cqZUyh6fwH/GnRY7I9pFdA8Ke
YJetBE8WfazdkiYEg+G9i81mNC7AHtJnxHKmS6NFG6Xase+Th/4TEvTfiKezuIwP
WXwl4ywdthZnHUMGLeGX7VbuPJHYV9m8lnGHjtZ86R0OLcfdSMNwXQ1XMuI+I1ym
eiVU6cFFZHNbo96tbjQNeU9f2OhaIWfTwQ6PYemS7xr4zzIhL7oL64j9OJ8Io0FL
epa4XcRkXkVtwXhI7aVg81VT6UGEj61D6FPubkDjDJWcQLsBrUb2ew5kENgwr7+U
xSwTVTj4UknrD/WZVfVqlYqZnguWlZedSMWepfoI3E3uF6Kk7DQ5kLIc67cURVRK
ccUWnUllAwbNHQnqfghSxEq2HpjjYjZ0ANKv2RspAtdN4PXxVgBilrKNgusZVVcT
+noH5O+ilm/efr7hfjuO3CDmGbIveWfdlW8uNcvjPBBj88Z9thhQVEABA9rOhgJu
ErFm5q7KU72JhhXXB2EJRa+uClGSh75lyzwGZ1jJdQ7vIe6sPME+EUBKHyFfHkiQ
5eFyt1mjC7VMlW+xdnpPjK+dCFLofWvpSgA9Qtb69aHi7nBEIg7ThFaJJLVkSbPP
yb9zTGHrtwwgc4TD4Te5kNKsDZbhgSyUREE9aCOKETmMmtKajpS5dHksryWNzaF3
RJGjVVyKQP2FtwB877HIjxuYLk9OrhawUBGq8k7gccD6IJ2d2nvlPbd6nHoYHBov
kkLyDQGjcoe6WH8k38rkJMMw3WsrHDMvLYq5aWLQxHN22p4TlrIXNUBA2ISEdWmi
McgZHK1QluvSJ4z0I/WWi19fHd4mP1x9HTzSN5Q4OMx5UqUzlY5+wuh+dZ69Y/Oz
LG/m99rZekCT2vL8VHiGZSzQg4N5KuVqEKE3YDaiEdkixplbGtVRzoZqGM4U2+qT
ohwWnbEWpMhRrZAfZIgDrfrDXnkhxvVbGLBOhTbcch8x+vWMPt9kzzH11I98ridm
EAx2a6VqC1vmHINvF+ChDB5S43dkepiYINQ0gUFHTwbCknkLtIrBtbCBbgFRP6wF
710MGQvhI+4o8V23NHKx/otCh1wcVTyab3t1CEWgzKH1x9eT8AIpQ9cpg0+o/RUl
8/iAzZlrxrD/0BwrlfoMQuWNSYIGMdm9+5kyzDMGvaAwNK3QJskEUZTyxGWZwSLK
U7uKFf6l19OyfCzsvXb6W2AHdjslJFLMAwND43NLRSN5esQ3jeOBvRrf/8N88VQk
yuAzpJmZ8Jvs3hEHw5WGhSLiQXy8vIQSlCg4gSdHY0xnssfRV/xo54+EQXUmnCF/
v4Rv3+/wwfPp66Lvv+OcFJBzTq75D8MhRJw5e8TKHie/DbQsFkFjxjoPpn6sB+Aj
d+rB5Jm14bFSvz4KYvxyzPW/IMTkTKRqcn1FiX8snuqtpdt8LiZEXjZGx3KAO69X
2AjVtA09QZeri9Om9zZ2NmAPtBFkuNlm2RRfNVuYiAaQY7oV2ju9efDHSCiasjsF
fwOY8e+VO8THJz6jbKzGM+A/O3YbxWhrFdfh3CXWjUDSfoU5qZcQ2w7sGJhMSyx+
t0g4KDwNBhaurGsoIHulEvCjQ4Q0JLNToALZNpRAuLSDLAjtRUc4xmEFJz7F6fed
R3jiTyTqtg1sV7WQZjg1ljE9+pj8UJ7glC/SW+2oEZgxrygH9SZrDShon5sfe5Iv
zAnwE/6WVDrdt/T4jXy0714Wop05DWegF69U22anXHrL3Lkoft/tRzXlH+jEvnnM
X4EekyczIO1PgpSoNQortGaDivhWJKACha2RYaCpOV6U35vR2xiXobq+N1Mb9Y1G
rOvwy4DNq8CksTAN2s41sN8+8XI6QfgehWN1Qpjj6IbR32W5DGvh8iXxKUaw/Mqj
9QppTfkUecsq5QSQ3WF/Drya2LzJDcSiW9jzRGGiWWKU6OJws+xaxEMcWzBzJSjR
gn8fXNzRDu0euQL8joF5857PRCx2AUHt9Z4DaR+V6NKE1X31e2J9Xb75gk+GiNTU
UMA9C3NGVy5Tnq6/1+S2rhMLwKRUM7AUVkEwhW+/3MHiMwbw1uErZA6f/rsFIBA6
YF+WTxn1XtFnxovF2nztjmrl87pdMoHILyQdPj6RBq4X9VqrHeaX97sboIBGqVDy
ODDMKgJWakfT2jkuJZAcKogrdc2PUTSPYsFfr99JZolIALD8fabfb9XRHoAwZCRD
9ca/HURQ3LJDobPtnvGQiqrHyRy+AIf6EvEl1p7F4C0cVkNEvOX0Hs8jaIYdSRkn
R2HjBdgnsQCze6unshTTEH+DMrgTDx7eGM7RXamKDluQYk6s/jkXjuXSh8mzWIvC
/rvP2O/+unWOGxFOZUNSA51i7Yq7TBJyffFiDS5dvpyrdaRyMr+4AU+tC3jdZmi1
oKtnJRwnSlWzDxp3lSBzb/cP9TbrMr8S9ltX7QVNYLNVw1ymD593HLmlnU6P39XQ
VkVznX5eiw9tB6fHHo0G4viLk5KX4X9gc46eZZ4Mzp0KwcSDX7AsPwW0kQH/AAmy
UYJpnSLUVXKwc8nimejBUVdsyKeJQcyp3srrXmuINtPtRExCWri3/oCMeRVOM7+s
SToO8wo14pVIBk4MXwPv+4706kLpMCwmQKGitqDm0+9mg4ooZBiciCIiA7ZNmIOz
tth9SylGxmr04nhJWQq/vJD8JwzHT43rva2ZOfHihj86H+vvCzpG6eluuNi9Q2KJ
Fu8oTQXFdmn/YRuPWlq08twTSe/sDSKWWYJWgM8nU0lhNktgHfw8MupFd1vkZBYh
EBaQW46cOP57rJmXyn1MOvd1T1F4dn05BwBx1uOa5yca1xRdM0KuLNcezIcoiKQq
JdKEmuiN0ePppELkVv8OXDY6ZuXgwUSNqr88b5TRpNUWHgdmIVR1S2/kREmTfadp
aEAbBcOr7sFtEmXEkSU5YNKcqCP5Lv35pcZWKUon+SdmgTrFPjyPV+mXxARB8lc5
UnBvDJedkwR+PhLRomDELurSCfrZE+nt4GLJL73VBsCiTCV6uxRVuGMRtvsf2jSZ
KfIzS4WnxNQFQOV27fWgwuakW44KAqiF7sPtJxzUEQ25qBnuwYxSkGBpaQcSQB2n
V7sUMPIjayS54folAgGRcDcnIhcASzxGcoOAK821KvqzrIVb3D3Mmmb8K3OT3B6a
fqOKEDk0e6Fz+swnbLR4HwIRmreQ3P4FFPeNhu44C3ihefhm+erxVjDutxuS1v5Y
YOgcAHn1DWqlT8WAP06Y673Qhw0rlNW7Ly8IlyUtwGWtTKFEOd/KI/Ov3U0jAYIk
8frvFXhShGgLMfeb1nFhQ1NIfTnC5w0qeOchEOjXrR8UhQBuxQOY3k+XiuHxAYWW
10dwHMM8Ys7iabcm53QAyXy93tH+mVAdQDPnmLzN2TEYVBL5Kj8l9XYQXKUBYXFJ
eCvn5qdaPIlH1bmI+ySlCSLUAitGiolaR7FSDjkYdmVstNznQ/macoo0TFcM1cQl
SYmr2DnnW07yMrwB14ax08N6Hq651wFKxWjb41Vo7z5Zs/UWclYPffmITGYFhk8Y
GhvcZ8h9RttLL5yYoZlMmq93aPhrClugUFFQwES/IHSyRhJT9KmhPCIdSaF/xj18
fYKqOzLwRxY2KthYWgsy0EdImA4tetAE8K16vcAXf/xez1vC4DdUMYLFf4dUq8c+
l+dBrPiOElZRgT5E15ShUjKjEVScrJw3lqqGbM+ZTJl8TlZ2+owiMhPRsV9EgD5u
lkQFVT24G/GDMIkak8JuOdMgbs2bXNZKHT8UKU+vwjcn0DmITGJKv+DYiLQDW6hT
CqM5qQrtdly0n8I5cP6nadhmRbNWAmXlLu/9gu2GpbUHCIURFpTt8zZDbwJZIqKW
JHWdTZrt9ikuxod9O+JE1JA8LKxt3u1t+H/9vR03kdD6I0BWOePqEQJ97U9Vu0L2
ucqd+TxaTlp+wmp9Xq/h/APzY/rzhMHencBioB985U55Ai0XgGSJEOu07WBuYH+C
vgCW+lbla+FGqeTXjMAH6Iw+zQIVAXSBaxFWP1nTrCnZf9Mbyb0WvIIZOmXz9Jte
RNzyiVLIqkCVQImeIEbC9cczmww6I+PnCrgkgqKizBoe7WCuG7NLpknAhJAZADvw
n3hW8hHIhDg0siiO0cghvLoNCA3Ft0uaiTUPC6cIRmzIK8thBZjTXs6l4fRvFU2y
eq2N4aOdtYJtnrD6uFrA1dQXBgmTB3bCjqKCKBlV4MMtfu4n07uKhYzelv4ar+6Z
4pKLKYz5BuSG9c9eHqOmscuMgbTkAoqNbZbJPkJDOGOq5CROyULX+8c3A1+KoHyD
JTWKuXeV+9hunlOnNbQOhiThBH9xLtHSjJPVyviz47DVFWQQ+Go7iHin1A1y615l
wsAwug4r8NzPBPFMT5Esdo6wLaXc+zeX8cfOa3PwNLS1IwditDf1QFtuvEua9e6K
8FEBMfPisReeUkfI62byrMZtJX6Sf9wV4P9yfyRJgm2BxLJPvf/Jtrxq0VjZBZxS
bhLKrbEkYbFO9aSRBN8KWCUQj8szdR05QJzTLnDjq72Dka9uZrQKQ75+lhgldMsK
arW6cgnKYV60PYecKz4C9N+0SxOVVdN3UO+0axrgRgGTAsPmRQvtV7guE76gZGaU
3Mr1WQWPpNza7Vjeoq79X/bdAoQaHpr7n51NwBqQTHL7MfQ3+6clabYLgIpwDjfU
gYMnW3psrqVR2tPiFVgD8Q9bwzP/Uovhq6VR477x3NaOyR/y2/8SSSEpVzP7u7jU
yZsA08nDL5iRE5YgjxdlC9hT9fFH/c+UTZE2EAJ2RsWeVHifLrsMyMMMRlA2o0i8
EApdQBqP+fAZODZ1mBoGTwnirGTg/dXVq6djv2lXxWuLLYw3Xa+eORhuwKueNKev
aFkSmNLtio+QclFcTNC33qSL/cHRewUxBFL1trKm4KhCVIWxRKatQOTAZdOvNDu3
mcq9IiYQHHCWHB3pmov7rbqfixjvexqdX8hymli+1p2f/uzg935/aW37zM/2HfQ8
gCgeCxTJmDxOTL9ngyMhzRfT6Kc9DteM56RfEGmFxQMmmuukuztTgv3RmXjmtLcp
RlP9Rwvlpa1pGeMk2kARHOeCjAAIQxMTqNYpoQf8v+4LLDF7yHNwvLtAZ+YKXfpa
K2RTyAAOXE7x/rmVoGPbopajsi4gIM79pFkZVtq0BO3aXL4a3SwFlApeGr38V8D6
//e87Aftwn53XoPV8ru0nIHPuw0RSMQuyI5xaA4jGZ0j5MS3b6+YQdxGhtpBn26r
XJTUjGIINfZr/icyiidDQYGafcrfeYc/jG6TOx2xF/KBy7vbbSOom+hWEKWp7b79
1ttm8GQkCrxiJC7CvNjpwCxUDZMdpnC1CkoHdRJqxUfyZbe5mepyzdFnYncjoDzA
7jMrV19rmdCscZCHljnzQAnjbKjxLBL3Rr3GUrSK8rqJEptZd8q7RGFu55LNgaMH
KGvtrHdmfdazCK+kuO8K41UcxCimCs9wS1CmbGqXkPndcw91IfVM+PeGynGU+8Td
Guzsv3Gnsoz2j8F++gjJDh0keZ9URjhea2KfKCrbY8p9XyZ+MJh9HlVDMKdoFDhh
gzrtQ4QI6LHheaXzMMhh97E2FMM3b0cBaXOu7NNICcAeF32dYOzhe1jYVqkBGCxo
DBWbB9hcPXe4r+VjNsWTmnl9ND49IfOS399QWGCaLWYzQnSVyxZzByhcfxIN2AFK
DIBvgNrVMWtGjUXkftDW27WC82oYL80nOT52cBJGx/jPodjHF4no+ujAWo9Dx475
Beshmrswj0iN0aKcfw4j1PH/mzgJpxrwIyPiYYTGvZNpsQJLTX722UQM26VIcVEY
3C7fORsfUQMiy60rxEeXujcZVrwwiHEmxBL2mlH7EznlcelXroFx4vLhsefwiWbO
kjvJRHmtueN43sGEkpr5Ic9N4KCnicM8YZ3GNUSbfB1ukQJ6qxSjixV6KOhxkMtF
YitHRAAnPAhyoxMN0c55DGztd3USWI5mgwP0FiQWH2lMZ/6GReFGtp+p25sv9KJu
7YqYB8hM4Ao0/jtw1pKUtHDpovvmZNdNKyoCUwTX9u2rkyK5cus4u39v08xjBGuS
YcLjuYV6rwq7IjK8hefMKAm65QYXZUHr/nxzg/U3+t8puX3KWRIod6oUGkMfwSo4
VBN79yYFO+Enxs0+cYKs70NSdPBxCzjP2sQvaywIp2boJB2adnrBneXgpSMpWmyh
AjXC2GmHqyxLGcUfTRq3rBsx0WzAGSyViTUwgTmtiVShxZzt2yxQ+a710/oqp28T
0UG35lpdctW6LtkQ4yhpX80ADK7DzoQjjycEKI1mi20jLRQkxUdirzIbHbNjzIwU
w5YQ95t2ljzbjeNP2ATiVN8aWflOT98Qj80gvsYx41UcODIYSRb/sv1h0LAIy37M
qxB9SNpVCx4kx3GmUzrRKB/wFfXhG6JLW7kwnCS1vGw8Fhb2xeStVd8En6hc/TLH
U0fhwyep+NHciXnR1TKXbzkzgr1Rno7h/8XLS3BWRll1iMWqAXy9n2xiJM+4/Z7h
ijWwT7v6z5xlQkpZ+jdQxonvdtAawiwXfjNpgcNRSKrWFiGykAs76pyT+bKFU/oV
TSp+QXk/8fb+FbkWh5q0b27yxqt/7sZb4HkFbFInirxT8MC7Pyf/+njie6FMdqpz
w0aROr/lITgp90LIJ4VAq5gcDdSDCKKEv2AO1d7cq3NH/og30KofEP/8gyoNRjcG
S/xSAfYZ7/DIIFAnRPL3w1L3B+y+Wik3grVsprYVNWSiG2yA9VcIOS+YhthgpN3/
msOoDTZ0NXA1XxiJsTMQ3IUDA05vKqCBtYf4LDJwHWo6hliIsHCA6v72jy5tLS1u
MAYfSRqOsHrgw5HcWRrPQdfq6BUc/x3bopwYPN/RAW4o41jyDUzn2oviTh386GPF
Ikp0CmRrfBgEkyN5dijj9V64Y1FlXVWGAqrnn9lV7hcwiDzKNAMs3LEaFEYTEirN
tnlB0h7WjDLgZ8QfuqzdiTFf6MqpEpocwk//KA3jpYMcgGx1eYWmL5ACmNykT5PH
/WrC/9HwQ8Py8rsJ7NqZgcfMwdLezeecTell5U7loAz16yhwt5QHKzkszitRIIKV
9mmgEZNeNyfMc77FtkxgG5rCknt0SXmENn+7ml8VI+Hy0z29j+J025e3LJHmiFxz
6i1IAOth2CKVqZPygxJD6/BniTGcA+ggn0GhKS7Gx/ZwV7uT3PlexPGeL7Eqgn7V
MBZQdrZFWIEeVqyKE1rW6cfdRu6RMsf1vvcafo3DNXA7vrgkTBGXd7BygIy+4Myc
XYQVQNJh3lVftG6I45uw3kz8I5t01Ywza4X4vX115VA4ak1N8qoh8ZzzSZhqa/QQ
BeRt2haDHNVTwDJHn8wmS59ZTR0nRRESuRTjdMAU1duh5XwoMb7v5wgWeaYEM+Bk
Yyv/sjW2pp3pOPneqwnbvdEaz+2B66lDWEJ3pSxAriWgnOJ+aKUKs5VTehgrYlxq
3JhE5dZYeWFSVeQU0tKfgqHKLfMPKBtB/abj3ZDtv3/SmUSHrhBmPiBudDVDBghl
opIGGeWDQAm/Uxg9cGlRfGUm87wMFo2kYaQ7FUc78dmXS+u4Rzhswp43M0hKYqGq
mYNcDWC77SxY9Q3ujYYDi27LFaT5o34xeOUEDNnYSi7yN/YfSoWTy5oSWxaPwwFF
WW2tBV+FT8b/27dkVZo/AAdwVX3aeTniZk3ac22KQatyI7/dtArA3SwItEelPvrM
LQ/X6c/c69+PMLcdbjXY5RKNrmLu0dfDWhSfiScQbq3bFGnsSIzkGEeLJ6v9MH6X
dQ92VaLigBxv/wyBMjwOmzA+7vnuaUuWjD4vzcl2krvdnkDhwnrgb46AYT/A7dl2
f1Rdx1m7vzrEQf29EejCtPUP31TxrIoaMBXhtnZPdnyzCxAgT7ZwjqK1RghDoqkO
MQoGIaLztflbtFme5nbvXm+ismGhoPhzBl6BMdot+1MhbOuSAkhSAymRJ8GhlDO9
8kFKWvHArDpN1ESlTn3mih7Z/jjpPKAok4GUKQ8ZIk4vzXNgYAiNYS9kKKrmxcZk
TCBhXdJ0AazpDb4rMUZKXojb6iarosw5TmHyeKa8bKGx0+i+awmWsghMs253yjxy
k5fsnCOEN0J0tIq2MzWy5yN0QWXM5eBhypT83gSZygOX/vbdRc3izudR5aF9is4p
BMOqae72EtIh57oZTSCTwztUXYdaIY3yPrcPvfu5GJulBGEJZZMEgITzeZ8SOMxx
b1fmfYQECLh0VDuhmiW9Hm23MTObU6wATzXenBS4D1UFCCV9wadZkGhmMmrNMRVk
zqg76Eflo2Nhme+FaHlH0zLSdWA7XJRiFRCxsOhFey4kDfujg9fUHq45VoACJf5x
bVfthRve9fE9fe6P3NZ0J7QraPu7QPxPq6IrCjnfc/fj5Ig+BDZKY0hrbzHfCQDf
gKc4xGRlsr1NyKM88xIk4ZnW8jSIYRjH9K0VP/JX+0YgvCw7SF3wKHr279aX/TNA
r6loW1MB47M47DflKKVNXEeNkvTsfrv7pL3ZMCq+MTkr/92G+gY34SnHm5C8+sFv
YlHhkJebGEpxmVhaAQmoRikYaY2JcB48fnZsyEDwupPYfo+WJxVhFoma18yOl58x
SUPuUKCexQBZa+RF5peESNUvzvvCYl+PWiYw/X96zUCTwOspmoR79sRpbz+PoGV9
unL+0J96IyywdrWw1qK99Ebfv13xjLFZMOQg3Of/FOSBiCvU7DFjOG5HoqyHigX0
GM7u7rjtViqOyV9lVfksiwra05b2OSUZ+t2WyWqzZfz6KQ1pfooxj3i7HArjE614
CBjdP1sbSzlZsoB1tuMu2wQzeH1g/1/VTqKWFFtmAe2GHAWHHIJ2pUMqiYybP5bR
8I7Tr+mAaUbZu0TmkTmLIc5mXtqtXGO7mdXNBgMB/6WFNCxD0xuI9dk+gRCm80/j
yrCuFh16eEj4MDidhacTwATaKIt+BZNIC33AlHEUSfd60weHtLeRUbygaZRTf5Xu
qcv+isOE4kRNU6EsqLp7Nemg1lam1mJbV7KLN/WW/h1Yv3CrUucJkI6u4T1IatlS
b5jYkxEn460VDSEB7okt6eRvyQUDMjwq0rr+gzsf1qjqOKfJ52SgL1WQ4fGNOIX2
ieIcrjut6+kJXL8Rg4ZDkdPxNv/Ypw++36YHLAoHCPZ6k+zSdJiqY/ec2LQJltt6
UvHcx3zCzK8SXpPij0wo1GaS2rHzNmxi5s9G2PP9ZZjaUpCWv7RGAYiKgnUl5AbQ
fjYJBEylKBIbYu9dSdz/yAw+CBN2xjXgId9zhF9TItHiTSFDEwQr9ozc4CKOX5n3
gPKfzy6jS5SV8A/XSX/7FCOPvmiH5tkayMEKnzOzH/zIhc1VRIX2xYjV4beAwqvz
cUo37uz/ZunrnzHlZRQQCt0UoSswNMF8EqhTUadKRugOr2WClDFZiNBVzs5tt0Ui
yy9CM6ISfIhRS+APJD2l+IholPsdXzapMzhVXoPH2ZHjKHRaeWwj3c6Eepa7ALca
SmaWeosBtxYCNij4Kz3Qi6ntET6YRKxMSbpTiF8M02F2k5BNBRxYgzk/MfzwbIUg
wePngy123Ihy2Zqeo1YLQ8bDByCvC4HSrM3oAVXd9AiATVJSeZrFZWevgOb0LLrQ
phwGxAUwoEfL/TwRGAAkdHmcgjBTtRU1xl7TPfoJoAw5CyQhpAb0bLPaouEvKmEm
Zp92ZrU7l+Cv7OmiZ/yGXyWvcLpMF402cHkFBgCAVUTnBRxowygODIW27OaoiX6n
ZJXvTJiVrV2FL4oJsJjslMP0/0I2FNK8zdq0Tl3U66IodGEPvOvmam+2WwdGJQlQ
b89LXd+dHh/mTKdrkSosy6g67nMmPEr+KWEV5j9pFhunJORC2dAZhpA5PgMfPgfy
OVo9hOjpcw42bNeG1Xp3C/PPSaBtms060gEmOGD5xS0aVkyVQRoMTP9cW57AwDKH
CXj5CRRx3hg+M3id+GEoWOMEzBMhsIpj5mHl9eDDahIogKgtxZN0lNbJYahWs4YW
kaehicMof9yXss71DY2M5M5+Xd0cPVaOpVOOGhyhQY+XX7233vM5/9jyH3wo69Lt
FWKIBYaFbkSRlDTBkC8niMQde+nEd89G7eKZFK1nuiKufyeH+PE0nDmd/gFKZ86R
3JTaXc8Jr/FAGAaISUcBOcOTJNAjRi1zrHue+E1nHLaqAFvOuwPlXGvV6wnHsVYB
P+61UTb04LezeGhBXadsswiPlS6nrgFHTmP4ZCiHdn23vrDWlsZzcMWl6OJOiroA
Vs49Vu1LO5NoDBYIW3PfUt10itEPpJlkX4Iaqxc8CW0MDgsLIB7vVl4eATllA/VR
5Iqt7UUpndz8OeTZKMpLSO25L9xoV9tDqrTZmE0jO746wlKySvfS9072ODq79/lG
OQGXNUEV4TiEpxNU5IRtB6pP4U+ernE0yG3i1zQH37bWnY7AidLTQ+8qovlcSUHg
B418QdMHbATDVPj5DYJbDRi6yS7P/gJTGOVMxfovvrHF5nbS1zyMVMf0tt7YyIm/
nO2NCad7KUGhRUiIA8aQChQ1pfmsU/2GpYiWzBcxdBlZTifO+5qoBiawxo6A7Qqo
ZgTWuTJyMKrGe5lWTOTbdmVVsaG2sTuvRCeuZfOL/L17iuNBy8+YlTvAiFQO0doV
XyTitu6dPuw14xl2hkFOF3ZiDBmaTSiOlGvm90AVcn5r+YPYjBVWAJT2n9yS6D9s
NIcVEWMlciqLhhnw4+6r6AR7vbl5E6dCYqS0XziPXUP8p6HGqH2xC+2KYn1tFFAF
SSSh/vMi7+VZMp3+1xMhHPTMFboTo8Uw5JrrZTyqxiYsZplZSEzCRWPiSRmnXV3A
mnynYTcCPrdg3tq0JFBcXgluG7uDcgNmDb3dh01vbDv/VigVOj48MAZttlSn+fOl
qwEai1qyRXmAWNXg8nqK7t1E+gNQROT/4CJ+k4m9zJDFgZ4BKlPXiwc9r21Ql1L0
s8Ewq4MzHkqg3f7fEv8ZFXCj2iVhUQfz7UyUtHqXDl+KU6Q0lSUfP73//cCQZIG0
vG3vUkWBRNuAngc3soxPR9ukQKUGRqcEeGFSiSYk3hYkEadOe1xSjHtIVhPUV5Y4
Y3o0luuDGK3fvx1oS8wZst72OE2ke4znJruCBke3m148OovIf3zRQc7LGJorpBUE
hb7HEefemPqEXZkbiFWdWdjDE+8UiFvkPGIb9AnRbpU4y7H4ZHYq4yM8XORuoR6I
EKAex3nEFj+oWneKEq/UtiTMgBzEY746b29H4No4DbkqGj2gFup02ac1t/uVqske
1GhBd0RYW6dNvycg6CI3GHeMrw23z9cVZfEXLvwvIEk/5+tELS/f+Du00elBBEb7
TDvN6uW6Qv5Ja25VNlXouVwbW3+odvbE6Pj8tn7VZKOIzKJ/CJFPViLS/tvazYPw
5R9k87nOVnnhJP60Xjjc0AvHXcoN05tLl3lBZThCb5q12cwKa2JRXwTWvGsHghWi
rWbRAmWpVuRABEXZ3tICIo/xHhZJ4qOfGphsc2ExsCmX17dKBsCsVbqOA39jhvH8
9QW01DhpNn1aavORXEHsnt9sEPLJx0wee0qjcC7XURrfB/sw5KDa7IcR7LukHYFf
URuI2QBGS/ivXYwy8hB9a+iGdy0Dx5qfueR7Kb4abs3kanUVR2BQ9Wr2CgYsHPnX
DmSkYoUJK5XlGmGCw/6S3/LLvs9xPj5f3PNGWwgLnBVWRdKG/YhvGMIQb9R3wCBY
i8bNZ/tYtS63daiqWLBfqv2/+C3lkUx3GbHs1vDvuyVJ1jc5nQGWcR5eGB/9qD5D
uVuhs3DUPa0IehoOBrfAEXFaaETFNxdEsiGpmoC33l5/Rc8g02UyOL3DvAp8Wl/5
QPPZY2acGbMN3+urcn3MkwbWdYEnKoTBwhre0wLnxEW9XiiJrryWAwvp4eutzSvT
IX3BR7Rm38s0XlzP3MRyHWxV719VLo6ptIVkFImWT3Q/zdNbgtX2kU+1tnYXLYy7
Uf7CIGdDjNZ8awwXVGLZl1ox6O9qopT11QvmhE8hW5iASwjnFIJqicU5Hpg7JHVg
l21zozfWh/ABdF/jarlDHYONisKE4aCQssbqJfFvoeJqODA0dya745Oxk3E+SH/d
FftXbMgJW8p4nXCDDa/l4ExcaNKAVsWUsB5HuVwikNaY5A3FX3SAmzCLxnyJlybE
8o8LSJPZ1bBXod0J2k8NkJGozrnqpLtax5AGoNPXkgKF/ETEovzFxBQtWfowiAUi
//OviGtOIB6kVGa/SMPrqHDyGMvZg5059mVa0rpWnXaCfx7ffAKytuv1TYZ+bCgt
A6KqUAWFuGNPahg2F9kAOlUUTAaxcZTvsBPdqeAbDD7koiJj6feWB6dS77M94CFq
KKTSoefZMy5KsumFdcWL7/cDNasC8e3BOgup0Tuvapwee0zKifQQfYHoDSt8mvwZ
a7Zbpap0NImifU0rOxZBpNEFVBa/HgnGl+3WAOZJwl7/dhCmiOWiQRWIa0Yyv3fz
p11dNxPJ+6GLdgZHRqhmFEfZTaat/Yr5zWECZ+uSR78lskb97DMSom+NzCH5zjI0
gdzCNvOzR8witZygb/8AXnFQUb5Tn31/nqclUXgWG21YdZDVSecMFD6TWTX4vaMf
2wWld27DCfOMebPb2ZkqxseLqZtV+Enmmi8r5/+MP3XHghoSz3ZpTmXdmUJwXBzZ
WOzWnNnfEUUCNPpaDhM5y3A3VL6ofw6/Y6iWpxc9ajv/7ficNAM2oO6BnyhjTIiy
9JinyWTz8pUUHUFEyof/wdp11holHMOjqPUx7riSqYj5Vy0fcp0cR3gh/590g1CM
StikuAKVCtbrBbOqn9BM3lOmV3U42Ms7xRh/e9gY1ubtKF4f9JxRwMUjz4s0SHja
5GlKnEmtlIOCMP8gynCZImN0Q1eR8aV+QJpMLRYoZ7YtwrsAAJbU9EfN25zJ64ou
3y2/Ao+8L3beut+y0XUDGZcwn5eS41uOGCB+vYUh1rhKbN0mGycDAGkimberWk2o
2zyXQj13wgGFZtW69O8Y47J6jqnbsdoh3siT9VX3Cv56ADypUxRLBV9/sa4cyECa
A86ah2mDqcV3Hu8r+toWRwWcDQhNxmR6m0t5xKhWOyFjpqFJLVWnv77osZycdpX5
hWZaVwXqY2cigIEMZ34cT9+s6uhBqJBLBe2HKyh6FsrvcKnMeZ6xV6difBDEn38A
gFBwy7/+YAZg7l1wD2SxIVhsIbvRQzmavkQ5qsGfaKIdMS2OmdGu/j0yi3DivEjZ
WB3v1trWyZRGQS5Sz0fYd72KaYfTcOeniLvS+bmHWSNaVnGqNODuE/hu4rcmsp5e
j2f2Y/2oAJvyZSiq0yKufv2T2G3LfnyyWHc3m1NPMXlIDn4iImo+uebZKXmLorNa
HtwEpsIIgoJE0QZH+aIPmuVD0JEr1ak/5nNnX+d6XXLK/9ONGTYE6Ksz0nQwvykV
oc7zkdgeK8c1mmCVD4OGlgwY0WW/tJko2jZ0OZOLELN0ML8vf10WzY8AsZ1H3Y1J
Z4oR6V9pqQGFeg0bDhiNqQuyLIqowObkSFEkfTZQzqX1GR951weSXVN8icmnFbvs
k9YpK+Asyz13HFwnLCjFUnYPagHq3cRss2ia7w4VMo4hX82yFYsvWUb83Adj43D6
fFoc9OrV0s/nIozQQlK0/DLqwjyQC/yL0eMz1vlUzPl3HbnjYa0pr+RDegPol0XP
fLRCCEhsjWxP9qkR2fQfe2MAcCKMlPaI/7kw6Hzg3FbINY/5Ta0fq9eRkW+PjvZ3
gaqL/VsgCDUJ4PvuOxgrxKdY735QGBt4KVLjtREzVEbI0f/dsyGEWd7lXLvaduAc
ypVpFOeh6QVAC43UhGZCgsS5HltQ+a1//I9DUYwNuDxYZAORs3Q9vbJIOKzCfANN
O0JfrcjOqlE60Abn+vLsuO3Wjg0Gm9XCfZpi2zJc3YS2zwnVjkddmd42FNJJOr5K
Q9XRdfG49W9E0KzU6Ss6jNr/ctOG9R1/859zA1XymR0d1OZ99gwHuFhgfQ0mwhKA
1yocc7XLaw/VlRuj8O6ZMf15ogPvXy2x0Uqj6ZAasOtWvrmgwppcbeEkv3hI6dsD
LZbK83YwJ3b0ozVgKk946bVlKbnAIaLvXlNqVa+dFNqB3azKRjt5vYNRw4iKDwxP
DbUe5ivcYrCwJ8KaRFUhrIagv2y/BWtF7mcUzWBvWcjGNQXNXA29QwReo0Rhz9fq
cuCG6ivI/SpsyjG9hQ1L6wdUgCk5t0DWJW9v8IpRgqRmVeou6G7GP7nOK4AMq0Kg
ix4twKKlxhzO8FKLleAg4rFPboo2f7JSQJLfPIkTcotxluEDBtiDH6giu1VVqIF2
wlNgtov1pZQZBxRNmBslAMaGNBZhyLoICbMlfg3opHGsvCcg/OOM0HEXxMwN3NdE
8lsRLI/a4m3z2F9njRY/GmnFY3AB73ikjkUj2Hvp86jDwdhb+CbR8LYUzF3hsUlb
kyt8hD3WBZ2ZUuLeTW7NpmpHOXuMyQIWFEDx7RrOBm4FLKdbn5tYfz0mxyGattAl
VSDL1/5rRt4t9kMmzYVF+fPt4HFiGLPbZuwRTJo/dabXjeq2ngmqjD1LTZ6o17ke
TOuOBURSwA+++8cwh48KTYHzof8a+ddWoORPUlwqk4bdPSz38aEm7A4HTHay733H
nIxy9lno6aH9KlSteC5AhEaJpv7sRgOvD16Vj7H08/L48ZRvght2bHhOrJmrhHR+
lQohCnsgsXZFbfmPyOQIfK42MTnh250RWR23FyoO8dEcMnWe75lBZrXvLNZRSAm9
u6qAKZ03IXzgG6HSrBrvkp2NILuCNabBsi/DAhm/5UIKCXJ+J8BxZSKoLhdwTnOf
CyAtZl0giPdOyq9qPpzeYbDXM3OV1LSWAYDaFBqXHxygye2/ShxPMhzVKFtOqLOs
UjDHdkaq5hTIw04BGizki59uVZk9+Gho0rWLT/0G1DPTS/x+V5hikG2WFbda/b+W
LE2EcdVKtW+e+zBXkawOq5Cgp8GBn88kwLPiZZ3/9WkdCb8k0HUqKaJpTCBm6e8q
yIlj+r/VZJXPfTwxH4Ourj2JKPlnywK7rOGh/nQfF1UdEm+gyBUnb1qpGM5LYeX/
ECs2+/OcWONQXraLlpR4S1JU//h5/BBdFYKCGgodnYMZOPZjHWXKwD452myLv5K2
HT8Vm++/YY+umU3eyL6JfSDJ27D/VQP3h+4IGoKgMlzZ5G4Kd0uQL2HTzLFLSode
+833Ok8mQmWHBrQ7ErEVQZICnTk5KVLVoF9OQZxL6VMjEONE2whAqZySqD6e0TMo
mu9rezpAbihfgBeXzuNTmRZsrZhOQA5u4Dlum7tsOvEFLo+3kPxGCuW1n/1WeLym
oM3DmIjislnj8n7cv/PB+DbKqJwykjhHdGbEnw/DEhRyPqkzBZYou7XgqrEIixwL
Qyuh/UCrJ3NkUbqzf/vk/RxbM6LPCraQe9Ua4QMUY532+xZgvJ5FDh3YwrUpxl31
JFCDDEvSZ2QWHxYDHEt/jyVNvKwPjH3EQIRT6gsrE1foZwwqPsvWXQd/woTUOIBY
m9t9KwpTe1SyQbdYtuuf7flouoXSONAr20qF3DGOu7gt0Fcgg7vuhh2GCblXBEzM
hvHKr2pJZuGfhZGt/ep7eqDzIRgaHuGXwdhV+RaihDOBJhRc/1aSpFU0u35ylOoo
zig1fpq+7SlkEuVErMbWEo8cCx8fFoGFuZ/fwvxwvRx6mjPwmiac3OICTgLKRSnb
ruQ3drAk1t38MsolrwI062U24wN5mwq+MQAKkMmDzTnmfm9p61J8rvTxkLwjogIs
0tLJTfa630TOMT9I/QekNcsvFZTunJAZafitB71rBexEPHlJd7L3s9seRnNwsePH
tJsjmerR4Or9ogLrJL+xpgHM1gYwxNYpJSZl8EqX2PHFCrl2spsoMszAkNlvJ5IN
HD+hvANq4R49qOscWcEpzxXCe2ZmkubsIYkrDsicBZrHB7DPahEfDC8UrMkpD5Jm
mjdjej8zRHwqmiYKN7Ub6SRUGMw1Ivt1RPEWAyIhAxBiByYqgb7yB4pheoRH4leM
lNXup/uMjKPSWoRe0tR6RdfmiObZ7N0SsZIKz7CVGroEHasTSWEvJJQhNKzVmrnQ
1fJfOrRbwkJJ2/h/7JlAi+8+MeZXSe7NPwD1eQOF8QyxLN6aLI/gyUtJag2vifUZ
QEGNFkUXC1Wj2SBIutJg7sIN2rvZ9XWpc+I1qbQFxEd+6QqWxPN4qgouRcx8CLvI
vrWF1aQdkdzNHFS0cuyhogYxluINWwWz7OpZMySBcJnhckok8jVy0iZomudU/aIg
B9ssmlxI0fWyj8HTxuGwDmuUishVNKWnqpBnXFT8KhPQmJ8kyU4+eqzYiBVSPM2i
Rf2ozNbvn4/PJVK3mfFkKLa3joo8sjcUasIOGJ/nDn6gpT8CLFA/Wy6GGxHDbbHK
p5svp4cnJLbQz6dAWMLMIzojwdxR+J22ZPOluYxg2/O99kVrdTvIjw0S++zp8PMN
wMEpgsUr89+NiBZpcPLvVB88fsiYfEDeaJHhjoKxaaml8nur8a7ChVVUQ/j0+MyP
ridVtAVLqEHQpEyJHzlTIpSMFaBLcdf5O825q+qSQG2om65wLzFHlnqSq+hXJAUS
wXhDHl7hBs5aVDHqPjuFBComNiRcRqxegPKk730+tslJt9gb/Q3kCStgNphmz9o7
g8O4pk4SJDrdqZ38N32NchMOWDBofyAv1ILMPh4KdlTN7Z/ITEm+/O7Y/qlu3Lun
mUdVAz4Vj54B9yZnwa29oKtluCANKq0AQJDfAJT28aEOE9dkcusOOs86s5fcm7JA
MvwK/Jg9rm9Xz98+xsb1i1bRb3/WCRDKlEmS5Rp13X/541gPeqdSpShUqkXXGuuo
I8yAyqKpqNjxygJkR7nNHSMbOUkUkZO3Hw/jbQvXBg4BGCRj5XvO/L0r8e/PcdB6
Vuzeh1bpcsbX45jhk321oTFxWw5mb0eLToSnt7RIujESyCjx/0fwnXPaIPQjydhQ
I3C4F2AdWKW/oQxyd0nXWwRC8UStGmNJhiVlr7GJfeJZL0aqnrtrFctqiTfKcsG+
sErXTbwNmnQAyLMQ5Au40SqOs1eFhfdZzb53oqebs2UgjPopwbq/Accrf0jUTOno
e5oQ2f5Kwy+5inKTWe8TS5BOcdN8iC1D7rruf2dcpr/6IK/bGzuFX+XLj/YLoIOB
Py7pjQ8+L0QV8jdGN5B4fprIZPhLW1THgg/Vj7x/yYUG0p8wE5Y1Z0ccLuHoESPS
sw46NYzb5wD6B3hUsjLDiy62JLtiKQa66sCxdNzLxU8zJAu15QZJcQZJWYCLUdyh
CwGGD/DX0KCzxqJTK7jAqGDnIpM5wBpps+RDS1P0DbkZQqOQAu5BNKHFpVXeGIG1
108CWmxxR2QhNRTyAEPTlMD8iKFH/czdnUGX2iIxAFbvgmLxOYCmXvPvYKCuLwWE
fImJXCQ6TxyR+rOHAcWmhsp+7esOHyz6T6GHegkJ3u5itgCtDoThP4oiZh/yuLZZ
ozoitrdmPthjc5bw9fhsecijonT5UWsR9nIZ9jw8M45sN4F3bT4RXl7TO4l1s2pz
Jf41YmH91jzzN8NZ4lYGo0B1y3VO/8UTni9PIwpxdJYHrVUA6+7KINYe8FG4AhzX
0B3HzURgZqJuDHMKndD/I4Cn+6SluJ7XZ49XNLC1ojhGjNvEsHfHu0zyYp1dJ4vs
lS14OpzUgQ0PNQH3Kb0xLpsDO8zBjqe3bNpZjtCPQhUGvWYORwfm813TzLgswf/Q
++yGace3mFBTiIiOTcQ5B5QW/lBSY+rT9GTbsQDOdaWxkGEkpwy+rOp5AgWvMC9Z
Sun+IO7cQc98TgkYKj+oHWz22Cqs0x+JYIBE9hQzDvAzj37tAdOPT8KxoOHPrlu9
YH6Nk8LRnFP+DG/GxIVPAt+dJrp4mFwgt7CHmPdqAGVO0/uOCSVziomHBjkce7E+
yT87AGCzZKuUVSwVzUzJPiDHDGMz9eD8c/L2ZkXDg9yFM6IYe91CUTBI2jYmBDKy
OUzDv5kZIemaKtYOmwZ7KZTaIkPBVBd/AtWvcqFDtSXCyrMhvQJH33GbVGujNSzv
pUeX9AfjSGxrSiTKjE5qqe1wEKsXKhBwt2+sCSVItKVJZ2u7J9PYdkystOOZMKUI
rSfCG9631XDpseqo2RED/Hbp9XISeFRBBaKIPU13BOaU7pX9eSDbLprQ+2XvaH/T
IFJ2OUvDjczb2K2B8z5yUFuapUpKhxwO4JNji1HUC872yh4Al9hGBTOGQHCoD4KL
ZH+v2Bur8VXOiTkxZjqRysoa8+pKgVyI9rxbyP7lqVvwyLeApci02VAJYTFg/fr2
LXlrukfcTl/CCCF8ljgYajRK5+UMOb2ClkSYqaXgkTGOtbUk8XZJqT10iJ/Z6w3p
EduOr8npHZ2xSX9I4TNRMa9O1iXLz4Ym9zTTHDV8HnYhfZ+HXjD6p4bqSZ48mxpn
lHEIl4TmMqQMzObyisZuFxKJ6UmglO75odkhPScA9nNvxlq+5KLgtMOlU5PFwTd4
9Pf6n1ibuWZb6Nfr1nEu+xgxbi1pZIPHkFtnWp1JetDd0VbmBMYaMiGOdMG6nWJ+
tsY+jZdOAPu4XYNlOJvL4lLGViVmoqMtHqvxmuaOsMN04jaedkeiYwDGFwkE5H1F
CJfnAitvyv8VVmyQng6DL7s6BsHNQZlRrJk2pClND5ssysUlRy8MXlYuJPutqhfl
939oiIHM5RNaesKUS2PoK8dyfF2iseBatPCA/P4QzjG4bPk0Jv4wTwFGGsX2Vb+s
7ANYJyBe21REOXvq8uuQl0l6vohOI60xowaa5CP7IKMEp6lnTktGMobz7gXzUVL7
rSTR+y2cmb24JmiDfg7TA2U0u2/zetOwMdz2H90PZbS6m4NWBw7JxtUJ0q4MsnHl
czklLQ4PKrk8+ka0o/1LRECUmasq5Gl/d2dHqZB/6c4+ZB6X2E2fMcIMDjNcxwt5
JtklnEGg/i+bLiRGDtWeD0zfcRaKstg7zcu2djjZ6H/s0adMerf9oyLtt3ovB7OK
9gJt1nUtmnoVzEzzq9DS8tPwFnTc2ji7y0lVv8ciMaQBepcKjFmCZSw2hBf9kBQY
5QuIzs1vqB1jFUalH6rWiYApht1ucCYmwlmpK4o8j3NdhpkeML6w3L6fRcuv9PQQ
sJY0G9ayEByuAzo/wvrV747Nhq59u0ge8FMP7nSLB8W1F3rullPKoPKtcTgWyjdq
MkeZH8TVEEmcx9OfJFR4RuXJRZFSBXSnAYQJyiaFGWkx1dxkNQKtPVf4B2vUMQ/G
BgzZP96056/bcXwv4zmkwIdCWzs4Vyd6bQSe5otc9PiRTlaKRpF3t0FSiRjsDaTe
ml7HAn2YuwYzKDG80BdHv+dUmhs0UOK6opCWuhl8hd8vHLsD+OBedPE9M3SweEv7
vH7a4WV3TVPLqqUsmvxh1baZ7tLVH+G2KkQsG6DS/Stq/Gth943cZcv6VYCVFk+0
rc7RbRBUUnR+jaqKfMbE5oph9WWktGXqUMjoSojKLlRukMf+5LgDqQGC9Y3JZBZg
F74RvjQp4xuQp1tSPr8v1cqf/n2yRenScU9OjmSw9g/Qgb6ZDWcA9NJr4RxW6TSV
L+mz/PDs4/HC/IFxUliVDbw2id7N0V/9tHsenBIRJDSLtafepDRqGF3nohaf8Zca
0ZtkPbnhfyj1cz3LHl78sdbY8IWT+MoFYOdKBY/6GWJSZW46wFhFrXPB431fbx+z
OZxj4vAXweShQEbXM1WszxvsYvT3EyVtUBij9m2LmOvTTYqnzvGwoKOx1p8RIhqy
4zR0ZyjPSkjIPfaXI25E0UfeVyRQEDdKh8vGKKv7XiHgK+v90mf1/QM64NXJ1SpC
sO4kJY/s+IQpaMfIZL8KaRQ6Oa4goCKH6iVcBI7BkYawqLFj/j+I5LvldDCs2jNX
q99Pu5Qc8V6y+A+eOGRsorMaUG3r0ndq2Tozt7XXqsG9g5DsUo1KoR1LGum3jX2R
kD0CUiNWAIkKEnLdpsNsDguHBqT+wnkPEQwA7S1iqBpNdT48MvVhAkEZfP26YOoL
LOgpeT+LAmjLFvNcUuiGR75YZymlvcpSZlNTogP0WolV3s+PGaFocpiyutQ79K5b
+3soC6XXo8oat1ZFataXvNDJrEfzYY1vrR/iRR9nxBD6NcffQc1sAf9TYIFVkp6V
PESF9pzassb5g25/hJiDKoynjRQYNXnKSa5AgvSJUb+gI5CH/Rr1soOoBCV+YiMs
oMImy25koGEgohwOmjRl83D6AMuW3mdZ7O/kmpEwIy+AvRjNNYGut+bpzxMHrntV
ESAhRIKLjvH93HseK6cw/R3dspTIXokBf+1TDfcCF7sIaVFDoLrb7vSIGPucGkFP
MZeH8IA/6AgjkdKdB+ayCKp3rAdXc1hHNLUgfVJc7/4v5BP+9SW6PCERWnsPDco2
ruxNMOk/zAsW9jKdeZHw+VLYXCSuL7hAb7nNH7C2f8XeqXHc/R3H9Byc/6GQ3f4P
aR3pXZTRRpY29+oFQGTWIhIVFzkiMS0Auj9LPbrqbYGLN4qepe1Ij5scW6FyqLwj
ZVKxEjoX43IYhNpxsnpk3p5tail7JtGpPJPGibCqzECrv8frIIay3TP5hkjl5K6/
LY+QHHaR+dA12fGBgsPcK2SBIGV7Xu9/seftve7ZMyhzsv/eCQg2q1TAtCUkopjF
uv6GjlQUfoVAO4+CJuYjRXqB9uiuSEdosZe/DYRfeLbTRNUqM6anJJafoTNLBMhp
K0zISqUtPkA4j8I77+UsUQiypDPiaBNbNV+K6MVCxvTON18EfOyT4zijp9UNWA/l
3LRJFuvKSvOM0EV3JjuK4u5h+MS4XAK/LRx77cw4r09HtF2apjxD08FJj5JZsNwo
dc7SRtCup3l4hiRJO90ot7pSzn766x4b/nAOI6FZpUBw9kHbyiYDE/CqFw+G2Z6H
8aDY1kzkQExvtss7ish5omwpeY2Vw4DLmZZiNa6GoiwpBcRAZCYM8TQapwsvMADt
D3OApZuWg4MFwzXMCIsIbSnLq83JlREREVc15Qqi56HlHBdmSEpGa0qAlMH74haE
d+l/4slcANYxYQ0IpOew9PEG5fAIYLzkNWCXSs0HEW7oB+tdVno7gC57hYMYkoff
RBsqyq9K/Hy3e8jqZ5zr/b+m2EekwzTJMqsaOxnLTvADpMA9KyRT25/XXho7hraL
e5gFpfa4XEvY/cFEgiNwYyrLSwDoPQYg+RHdqBhDiHGUk8O2Ff6pDI5sEve6gese
z3CcS6zIZMJt22x4mC4b6Qbpf3kxSxMtrIRBdU6U8x3gLNIUQPLfFzw3rAGT0XWH
cOzEbLXgNCO1YQJpMeOr+IQqbABxxQ9fg2G3Ab5RkvQs/MwChB0wsi2Av1jTYgLa
5VkoyyuXOOAZIVKNiT3bsppev369VIZ1IPUSWp80WDKLlEhBwwFH/9PAEAHfvZqG
1HhYbg8TMQHWZm4eCUodUQxTaBjH2g4TV0LaYZXwEZHRtBF579YZeo83XGdBVAPx
3rOUAf4WLbacNr5OGNmLoGyWs2qNV5sBZUvlJ9ciFBgl1T43DS0OdLLQaR2MK7Vm
S9LlZJUJAvnWmLa4/+F5dMacdlihyruRzfn5kgQ9p/DISTlqxtI7thyyes/9qcE/
rdyMknC48sDMnv0hiNQkrciAlVd6A6dG3q/8tIAzZUl54xjcEWbNbQPMxNHWaC5u
eirLLRcwIUAGwG3Fy53GUuJ2KBpwY2sd5zgiR6sXWZ7r2utsN13SQO39piG80Fi7
0Nnkc+EPcjY+hHtnEQu3slOyehjrQ38OWbyP2Q+mYMgywHusj7fZjUllt+7xWbs9
9t6dfw7xU7vB85QQl8EWPSJf80xHH2Ifs5kNCEl3BSdw5n7y2rzmoZ4jKBAmCmP4
KDqJJtqsQ5utkwJiiy5f8VjLx+6h0EjXYLngIlammKQeE5+Wj6qgvBQeIEqwG+97
fktBzc9/h1pVYmfEcnm0KcaMlx3TSV+hIwVh0aoohpbBGtE7oMU0ebYlm6HB3ufa
JKnXG00INQL0yi1ltnzXoGu65ALSltFJZ6GnIPJSoqU+PCNuIPaie7dWfQmMpIy1
v6vCR1nRFDD25MH/51/W/JNXdla8spgKTZntwD6K0DhcWKgHxbCpLJBzMPxJG4WG
F+SPGfGJDoIt1kPZVuI+NfEVxLJfgqUPrHlQ+dVAYMnNTf3OH1sd8rd0xVUXHHwJ
ru6UOrJrSUsr4J07YzbgzhT+D4DAry2VFELUAh8xrzz7hAtR4/fvxmvbzRknNOXD
S4WNbN+wm7AqENV9oJ5SH3/7Oa/SXRZG0lNcMciUSJvX9en0I6o9+vGlYjwM92BW
9aMwoNzVMsPK3iE/6MxHeUjS0hYJ2Chp9NQvSUEmnXkYG7p4/c+tlNH+TgoMrDOs
+VhFoOSkvHDmzcLn0CgXOlIqjlyCNSb0fbiOO0NUJESqzykGya55etzIuFt+6vD7
4V7SZ68y6nBybbsd+ybbXUwIbB22NW5L7jO8VXbrhq/tlzMVZs8cCqkxtkIcVE6o
NOksM+/qr+Om1RJl7dEi9KXkzRibGbUOttnpe0RRPYKTfpTkWG3poy93BYsz5Q15
OuEMYnwdmqtSNSXMF4CRDRMniCc5eFTPjBhA5ZTMpnKL1cGjbuN5p7dnSwODLUe6
y+SaeBpayb7//MvP5IqWOuKqQiNTnWtFiYIWsu/e3htsA9UWFmI6TeQS7vHeuGyi
UDXDc10UweYr/m05hLIhmD6SyLSFY79Vvceyix4tzhhHzSC0GS+ifmXzvHP2piWq
/EUwCoTicI7bXe0lmADNceon+eq6bzQz2vUVKRUG3yje49W6ltX7Vps2J0jQQXfr
Yu8jcLBtpKwI62HBqb2xo+hXYlZQ3XYeRH+ayGnhc5qJKjCuZ0PaTiFHEuIUfUXO
rcUmWTcabNcWov3NaRTs6W1DSNq2xo2NnpErrJ3Z8X51Ky2qV8SqF6j9Ap8MdrPa
78ZCp40jMhVd+V0uw7XffImEnbcLpntqdUELwO4jTbD5rDsGMZY2MPbKgg2vEweQ
5bR7Te8LbwAM1s52/DlB2/63kxN49TJv68nlT9Z47zO4rbwplNklPW+iQsB8vbHl
N2WUuNGW+hKAEsd3HxDJHEkiHkHcTJrwvfG5tjlrjPXbmoUnDa537MJwWIPxt4fn
1qCrIjHvjwcfGeKDe7nZhx+el91MxQHsKGawUMaTWMBicrxhgmsXhn5Hvjk2Ec6I
Gn5Jme2mDXgAoeeomzoclM0YemkaqDhqvFTv9UYYmsW37hXG1mBQw9VwxsuvJPO1
p2qFNUtGlv5+BiqT7PPsmjK6ZF+TWCndIszus8kCHJRg8BnXf7QOqXM+mB2NecGo
+0KSUIUcC8wiDHasnHKuTwYGy5kTi6iDP883Bnf1LNHMJULkmPNI907OB2Tyksyx
RM9wqNHaJnE1A2Af21iMdBo1I4fSZhox4xM5UVGWatXsrzlfs+nwe+uGr87+FChE
2RsvzL5KqOrorx0v5vZds9WAIp3hUAmyHrl56zn3eO8SPYugV8gGgN2nVg3gD1b7
EmDNExiHdTvzphZXm7mesOp9DreYvgCPXpiI7YJRJ/+S/YsBnUayMbwxsJ232Nkr
cWDoC+pplGBfE38tyK+Q3NLSlDK/+AfjxUh2srVxWKk+hvXXISjsD9PuAMUIC9zN
1auENXYKd2xyiVuY8atSkTTbcf6Y6ky1SjxP4v8iX0DcJKYztJdKkJCAaLYDdMKS
Xwp7cTK+FcEbI/DhQSlNoDEbrTba7Wb0XI/9NfKnpynylbh+I3K/GLD+AUWPVXM4
oNrReIvVDo1dwaLb/8aaEiex4haEwecJbWSYtJUpfVsOq74f3RfzQ4p5zdo3z1f5
BBugPnZl6P0zICw2kyJNFsgP6+YXUPHybSyc+ADqgHpQQ3tejQ6ktIXLQI9FywSo
sXjj8AkHNWfitAr37Mos0jw3B8+W4GfF9JGyQZbUcBRyogEkLbbKj0f4t3ftSEW8
kGOCo1zTIxZ1guj3cVO1IMhS8I/cjlVQ5w0Oc/oSNAfgcE17uv6HqEuOECH+hgsY
JIQeA6oJVMDIkEAb7K4atL1/B1+y13ksMDoW/OtkgqzL3w0uy5EmT0js60uaNHsP
fMgShyFt2VqRCiw8s1KwoSEeCofSR1LOX3iYxAEJPT9h8q4nUFYmq2/xSz/OdptG
uuomskqJQbiTV3kzYN6SW95UzyRUtumVzsO/NlrwIXLfgiQ6VsB5hn2EGrn5nHFU
FpcWWpHEdKbypTNpNldDnnaJpSKQ1O83PKj8H4UckptjSNT1AopMQpCeBxnWd9Cw
/tdHPqpD99o48UZmsE1rqyi9n+39fVIzi90pypbCqd1Vi71K9i6fdSbCUEbgLVZm
w6cEnDuyuJg56+ZSRsPNMJ2m8GyxoHIcz09pZBZwbt55OmAD563zr8zY7HlqOqI6
vzqmYAh0qXSETdoVo0l7XdZCOQr+aDMYkWxAIXGBkdmfPNG/mlcVRGvodc7e9N3W
URppBod1N73PfCO/lpd6fmBzqZxw9HPR20MVeZ3wCZy1qkqFtCjAyT0YDcVfKWAX
jWiyyz9nQz2hGRyC6GjKjhtPaEhRVeHArjQa6E4jx/rnssbx3X374zNc3aLOzH4T
WqzLASeBxddX1/HtKJSBV8mAHQAcx3tuUrQ+M8TAxmgesuZf5l/0aGSS2Tvgoy4T
cSEPj4U/QpQiwZ+zQSvRpB0LSXptvdo+xZozo7fc2MwX8RONMi45y0xZALT5avgy
Ul3MQieFo28JgLpKBrmbiUi3v5oOojEl2kAXtw1KoZdJPWKdbivRnNdDKMGp0Sdc
U6WQ5nB6DuMZ+7pvoHZ6S+tkle3G8iUf2mzPkuAwiwYZolDq5kbTcPx+Bo+YhYid
OrKJZ/2vG+hybUNnnWP2NgkPTlovkdXjtNEZ61D9dgXiWs6HWNaukEsjTT0Je+/J
SAERjE50M1qqWBrflDVFBN+XTyu4QwSBGyuFlP0D0KjeJrkOmyIa2hB3RsEpQBnC
UMlvcOP9WXNqpxlA9UxWjX5Ap3+QpNRQB8EAEQ7HfijUP0nRMGwYGwSxidmjp6Wv
syF3sEk3QM8SygPBKvLStKh7oB8Nc+kMhvX9d0zEaMc4qdk085QfxqUBtY5xUodx
pgYb5AB/ZiPWrX0oom7HDYWcJhgOsHY75L9y+9HgcrJXKDssyO2tZsQP2pkNBteK
LshaTCXI1rss12TGOY8tei5PiR0dOgjIsOkP9zIxmHB6PGx+i6Uy+bwvZxXO8qn0
cALO+nued3u7bpF5IbrYcNMYdTN8tag46L+qXSrlZQDKv0isKEzOLQ47Iq0rE93E
4HKfGFa4gSXglJQPPdijYA28eNpff51XmrtScU/gYKdRX7B72YMPv8cqPyTodYtd
OMVyjC1RYgSuihrRmGEB8ru+NqekPKByO0XY0bAf8FIIEu9gmDDc0GrgpNrp7C0q
7/hEAtBEVYnFgzFo4rqlwG7GcBeCaaR27cSVNIim1oUIpJifN1lxXoIBC7pCrGJ2
7E4Kuoe0PVXuN2SeNOhzo3YWNAqjkSFbjOZW0cp+nEINoJmlt8LIa6GzmtDkT7FE
Zn56b5ciqbBCLSN8qXYuP5k5ZKhcDKIolPGOwc9VfdunwkpskZpwmWsq2fzrq1Dz
zIxUuWUoRsqgxWB9zg4aw+S5K7zqEV9ZB3CraPTzaItWD+TbgoSkcwtvWWVeeIgp
fQYUOYEhV9WlGCoDvC+dTNA63IRp9QkzK+sxs9L9Luk4vKbeuB/ZVpgvW9v68dCh
mjQC3hORZDDLu5PI+iuLYn7Jtxo5MmmgSwGIgucVY9sAwN9dWrC7SMYAIZZpbNYl
cTYzfeTkWUY8Isaby361kJo5bjvnCT1fG+p29+Y/4kZT40u+3GYmGNFRl8Lzn4Fn
cYNmAF4k2XIH5kNvCG3pzWVjhyWATFMkkEF2jUJP52lIUvCoBX3/UcDvaoSjIVIt
JqPH25jm0PJwm1hKQSWATk62sgagw4uTdzVSXoxL8Ik4MK8/g2+9f9MlAxxNGupT
F5IE0zPF1GCcVFW2Es3iQTR828e0aHnR6OKhSqQxvUOmaTcpm05sL+/DkQUy4EUM
/q8QLFBZQfaXGB2YvrLX5DWmE2ZXAXqzgPEqAvCG+ilogKXv6wE5RUDo/PGZJtt1
jOk8cbZqazhGdWb6adeWOAdF6+nwEYi8A/nrmZWvfX62Ndlul+b0t50C5LldLPj/
YT1zOVNE20Fxh3IaHAcfyrm3R2FIzfpjApl7mHQhhZgy5y4FouLtS6vaCgRX46pj
rPL4lOdHhQBCS0WYjAjvCjd0XoDG9ff87iI3Usmqg/huPNsapg3/nc+XzWeZsX7X
vIkRbbJxkImWK4/xXyIm0Sl9zWvAW7LQc9tn+DrArYKVTv9FwfIUGynHMV/CZlEh
cknsAv2bS8Fsf8lRthciHHZw5YU0JUOa3mKgb1+vxDAUyujLOV1h/O0oymPRqSBC
YfH2+terlWT9q6UowK/q4gqTVZEwBAFIrV5rfEQdMLKM6to1nxkZ+9faBz/w4/eA
EVqXiv3xN4JH8QL8++eg6tENClrqgmHg0pGRxLmFC0jS6DpAjAYMHPgJ4fKo8tsN
+j/tgwxpZdav/CDEruBh72nw/Lxt4Jkv1QaK7UTL8iV3cyn+PCds+9NRO2dAQm1j
DLXuPgqZ+KGt57nGydgBc1cj4MDHCfkBwoqVxl6VWclix/IkO2zABDkqnU6h5qeW
TF5+C7YjXqAx4SJkoa3/mnXKw74gAKI2gmz+9jrhTy+cNmSSegwnQSVuGPxoD2Rp
DbCOKIqi/Bxm9aagOoAHuNSjnGM0OyVQCXrGksgyvVMZcUYTsrlxKAuh6Wg2ZTcY
nGOb+M5/WpyL/7y19+Ai0DwJQS+4oFpt718nQ2jG0eO7PbJFPZUL4Ttl/tgRFUrw
RY8jAcOFOaZNq57ILXCNdxD1sHA2dn/5f/OOsgUmU9/iczriI3uKdhb6lRPE4mC5
K07FTe7VQnMjXb4wEPaLc0NEyMRs7zvNj2YvrFT0vN7GFj/yrBUl3lU+yWX4qJdJ
H2JO78NS5oGnA8CqoyplabD2BAhwWYISwYpQE4Ic3W8q2D85qIqAJJapOVO8Fib8
ianbElFFQ5ZFmP5HiJvQXr43W3y9QdivTgbQQ84NJYcY+oT72csGUWWXtCeMvAKj
yN4/08glcIXQ2n1p9z5p0Q8OFfxOysBCAD1inYym4XEPUELsDAbRILwUmxgi8oR9
uwcD3XNgq0qwo0AFzHgzqtgd93T9+MVZ1yO7/5Bgut/glfxj2Y56I4GsjkxrE6hX
Jf6OMMcqLVvU7BdzElgyF/a1z/XsoyUgLLy7VPJOvJr5CeNbMl1ocIqicC8VWtuT
IpWQYl97QRq+NABoh270L1GkLm0zZGPl2iQNSaSNLn0ftRAfMpZ2FEd0AWM6da0+
n3TC6HBajxA4g7Pd4R8qELG6FxVhRaUaua3kIUJEQv5BSMTmaAEOo7jg8v+YRh7h
nIJ4iIHUA0MdcbmtibgNQ6m2SPKSOh7XQixcjh2iBveiKcJwPb88FWZJOtiqOMTB
wyhZMSuIx/U7fgDX6Lrzf6A0IiiXhZQA/xBavK5kAD/V5Teh8S3m9cpgoQZ7rhSn
Ya0RRmq6qtIBqiWvUesYhCIOz88GDxuoJek+7v/6F72KVGJdm02MIK94GKt1PRlI
hsH39bjKtHZePCqnWeMQsy6UgtAudNbUwiRqHZsCtYsdxkXvyoXzrdU5IzW59pF7
vnRnUOckX1NnpMXpjhE2aDqq/pvaiQsznfZOYgV4LkZksvbV9a81nmy6vYkG9YiV
wwg+WujYfkWULfwXcQvJclDHRk0OF8MubTyzDIHbU0uKxy7iO19XyivAaMlsi/RI
toq1hnS35wXNONyMReKrD7ylgWmW7rWNlnnyQv6ikcTlvX6iEDllnnwn/DUuuFpT
VEF7osKcH97eyY9oMji7JiX2/tnXx+wzPKyD5Mh7PpaI9j69SB6psr4vU2k9N92z
dlnikFBdm+gj5v+N796n369LYLnMXIz1jA3gx2a1f65FGFTGDpQzdjpGY22uK9TE
VmvyDVtBv2jC8SDEieoGUf/k8nYaXA+flr7EUmHj4s34qlp2wmXKzgbGlQVgDMW1
5xrDhunbpMsVdaSqHFRNDFd6tMdmoctVw0SLFy4oktb0Q0RMNgXayNbjXCl9MgXf
pJOMCPOROrjRvZcgKwyPqUp4/gcOLAnFIqHVW3KvSLf8yJKAa6Qy370TcdI7YnPJ
LfMEMK+imj+vuzSI38J2e92Alfw5in277SKcxo8RJu+73LDxeWhBzhwwbRCgolCU
Y74bqpMHmGzj3JOX7KLgoJaK+O4SNkp9r5sBnMsqbPCO/HMKx62SRs8PLDT/+UyI
Dzj2GjVE/MkERzq95heZWkEeW1xqWDjSSpmxOhuqq6y05GKLM3ACqQ4jR/RR/TD/
GEcdak8xCLiXrtTSNOlzCkaWH1L65qroE42wEcAWp7YEqTCRRD5d0Jrt3aGBF4ST
5HFOLvZB8HrEZTyDT8kAOW5FrjKGLhphxQGwchbpCiNaMBBqFoYYywQyNKLpphkz
gUm2RYfGTNX2m569hkLhLCGOUIDTq9mW2bTygeUYwwzgzB0xerwqBhS+mcTkccry
bdw/u5MXY9VtGpDWmzcjPVYxdsg4SCrbaGs5JwbW3LH210eTokI5r2oO5k3v+/L3
svI12EO6mxidHLP/3yRfMab9fTDyOwap+wngNMU/IfJp4xh0GinWM3xIRh0tuu6Q
c/CpKpOhC5ncN/RJPdFPBUiE8GQ+hZKvPvfbuBymKm2gEBkRIfNXAKVFSQnwuREA
b/sDqbz2LdYTqEhclLwfJaPTnE3kKmf7CPHgrudINuBAVAGoeZfAN7tkh4nbpP5F
aCTwKIjjv7nuV0PDu2wRGswgdIfo/Y5f/UA2x0VWXXJv5UzvnerZX/Rb6bXXN5A1
ue172yStgObhfj3rJwBqOJiwnNfAD8YjHYBoeFwMExJWTB7V3Bptlw+RGsECuw7m
i66D9M1BIi59KtHPvQJiSmBg49PirYqWUBltZtNe5tzVC4Awoop+Ic+jNVJCqpqh
Bul3Z2FU3jJhK0gsy5BFhKOmmzXOzr96iCn41use2JLtIUJ5TBhmDfBrSRN1D0U5
dnFKiuh25NI1Cxw01LHpzlTdT89VP0zc0W5my9FUm+pQ6yPywPuEiQdMKGpZnpVr
BPwjZJOf9FWyHPKaw94ML4o2WjRU6ISrs0dCX5XhzfrB4e8EJ9KYtHurpQJhzh2X
PUM+BcWhxYEimuP668ji/box+Gd8cggWvxiFpcNl59Blw1egjFgI0cXIiK5PFVCG
zpumVRD4bEuS8Alpmzwu4UiIEX14D5wyHJIDv6bRt/q+uzacu9xrBPhH7I5FITtw
4SOYdhXM5L2d6lCTaymldSx5MTXWy+H0XLpSPfQiwDsru1MktsMb144+XSB1d/uz
Ll2yEE1vw8AgOJFna0IdlxEJ7yd7G/skSGa96GXecXp7xhCeHz/JcoIjgJSSPWSf
nQYoCK/ur4MDDuzmYV6LwV45D+5mLg484OpdH7v81iTU1ue33MRpAXTsZq4m5o9z
QMnwtU+xWN8ukHWSkploS8XwkMosXhTtGCW+X35J9c4+/S5HjKOywKQ3Y//BmkPa
N7XLD5aEPlxC0Dc2l9x2Es0pCCPsc6GMtdSVDx0pvFkY4OyNsstO4mM9EUMChsvK
tp0JrYSk7hhjvSiDnXHn/ptB2nZr5VgNKm4SmcCgtumVKwAagzt02w3drPT7iwer
qqoE5bwbeNH1oZHU8NQ8caqzBPOXMpH2Ypu8COryLuEE5zG5uIGKwlLI04IXpTya
alJMePPkzlhxKkcv4aLi0mxpII6Vwxxh+W0N/WU845iE5JBqg8ONLoKVDswybbXw
OQLUp3TGXe8U+pxec9w6GrJnSioZsLUjknDFTqiA8JtX+S4q82YQQomXDKNPADyG
pAXUaYk8vfphzt5vgx7Kin3uV9+oO5B0XgSx8QzSrmFOBuBebUZpL0eCUzw48dd1
CI/XAYj0NFHRvJc3utHz7P1nBsFJ201XF5Fk0+jHT3oUiyUeIbsC+9HNIjz/g5KG
+855o7o/LnWehqPkE7m3F8VSyXPn2qGAX6To4IzqEGwmQIneadYwkcyMsTdZ5fnh
3FkHV7mCuqUxpqJnlfTUSLDMvSr2dX2MY6TeXcoVMAE3B6cR/OZTX1EP0JuYU27c
WOXkwAlbEzxZKpiytugiQNGhbkx7lM/YMg6Tf5ALWV2tKQVwj4ymfI3ZnsvAdp9a
qQh82kwDeIj6zjvk26kqJVvlk6Jjdhm5GDZbfw1pInWDFNTQ4xrTymS6VkFvhORH
2r9hP4Ljr9+W7GCQmtFdn/+XSE3mK1fKxsUy4n6fYZxB9Oa3lZKw2OvfHME+SpDt
pobw5EXkn+kcy/26xGCy2s5+bPkICKZqdIW8G7FHWjQlHEZYuKftzBQ0lRH1bHuM
YxFp/iOn07Ub+yf4hTino7NyeCFrSHKPVuJ6tZ3cetofFsG/On9EJGKraAVEQ/G+
lFua5j2JyWtJ90MvM6Tr0BgfDImKNyBnmO/J8jIhs19EFvYUE4Ww5TNeOi6Ao2zA
FiFc8ioB5AiwTtvr6DqYu3IntDLLL74hdKs58isQGqTuwVFhINGyun/Ifo5MfQwp
EgMzPAY/fDV6Z02wzmQ1ISdIVIqSLw6ga8SPsWgoitkUsNtrxZNTdQJfLYmqggHd
38nQAR22ZdX/fboKOAeepcYOnIgdGBUabTXQpGle85LfhbgLE71uNEbUfmfYk4t7
Pw9vMy8g4g/2ffOgHbDEmKyXNjmegRpkD6L0aBo18VkqaOyB0Ir4fRgZcgZZXMgE
tMwdLmdfhgY4N1oiR2XLmX0q6++tFq/rCPiLMRt18YfhMd9q+twYsYoHQwCuck84
1iHCksSqjk1/9w12L85kyWxCiWRXJYw3Hmn58ga+AmY3k1vxMznoC4juTSqwkFnZ
gj7/pb0udp/4yZ+WKA6XZu85nKoZK3DTh50oeCTztGZeqWV9AS28f9gapwsTa+k7
NJuwkM67VyGYNeSRuJtp5Y+EgKkFR2sLRNu0/wTRYSimQtWkMyVl6nYymgbFCbzo
29umj8+/vRMqqcJ4WXXwxwQrncYF6BISsXwWfYq8v/koIMfnN9e/wk/ZyrQql1xC
VowgXbWyA+zLUPjPjCzcbdwYo9Au3ptn8UM775xL6PXZQIGZt4gf56JdZHxDwbPG
mm/IIrCD70sxmn8PrRuloKvGNzs/8SLiHJ8fBx1TyZGkdsm5Vp1m6bSjnneJCOz1
QMY/4cTr/KP6gES2NZfy8vh1TXf33Ihmjc9ypl4JtlnmQdI1INLA+h0ou3qRrp4g
8oNHHNmOq8zlytVNtrSJVZWLu2DgE3ScIUT/BSrIXsaGH4w/GqTDdK0BdAqEBcGJ
gZrN0p7ABz4rthN3tGELe8uVvJuIFAW6UtSHfISvRwhFvqAAF+cmMTsra31sHcf3
1J0vf9lWZQ71XCu560KeVGcD6BVTYPJhKN+ahX/FwW8bKRqbkV384oIZeEFKnonY
wLO/Lvft0QySGuejw0EDpA3tH5hcmiO091YfcyGm6mel5mepqnsDQDqqa5ptLaPQ
zeCxUd6E0RAG8L647xHMwn8gEzPxqpQiSP9rGwiJ8ULfmKzbXNmXNbBDs8k+N+dz
C2NKKs2EiB2zC+qvy3tjpYxMAtZLNM0aj6IwC8ewRw7t/3SCROMfBsaovvQYAYkr
0S80everJnoJwkGdmj9KymGAHXYb4VGOeTyOYR8D2tFA0Ta8E33IPEcwC3IshEC4
TvU25cAXzjD/p9+OzSOLA/SAwvLaWK9Bgs9APvatMSWw27D5bSts8/NapsSYbgXf
jmYmxpInEY4cLiAKGMc5/42TWoCiiciBe2PC6JevESVeI7447NcsvouDiPZYu1vT
PzPm8/EttnEVSdEsA+tV+JD/mewis0a58TS03bVitp/Jeg8mFL7wxfMT3Q1z3Ufq
SQCqzXGWBpNwvBsjyNDI4gpGAVSKN26JHhLkKpNLzToCz4d16q1o085YKmgX1bc9
87rTvmGGKEAqgMsUo6jVfjHLCgFGe5GXEEEKM1a/Bg9iDuRY3JYyeQTQ5ytDh9SK
64lbvp9ajpMWWOWtDIveGWD4yJiAf6thCQHqy3NSotVpHd8DGzuRQ6MUXZ71x/w5
jNXMjpE9qLjGKAkGoOnRNxFJ/E4RlajGwyOrVQccm0MiO++IcDuK+qbOqdAd7kXA
k2XadCnmiXPyh+OScDVczEhy1r2gK6MCYA6Gwc+ulbGTLdyEo7Fo5VavBMUFTNuE
GkNEcFpgW08kZHHbwugq0bVMi+B/L0lmKZgNhQwbOkRju8kZvUrEu/UWC4J+hDfU
BVHEQomLGO3Ta0MJZu6uVB6kNW6d4VoeaLXJGFv3HpTk008HcLAJXHbO1ZrXohM2
RZQFfdF79GtfDHtO3X9T14mrGJAk5N7eWCzFA/I0dCsevLvvRs8//EVvoIqwhWkE
KAdhC+Qj6nqh8C9fTe0UUcC9TxIAuSnEK53jeVX+cw31mj/F8bqM01FQL59/6gZF
bNcioCqfaKH5y7Z/8IH8gr8N7Q6wDCPMg4RNR3+x9shoqIxwuu7IzMOAsWIHctEV
9qHLS7xK2fn8qhb9EY68nNgifc4Q9YWzGN4/dnMu2GoAapkUcm7awf0y3giNAQFn
Q43YXb0N0HCnmk7YW/M4BvHdgFTxa102gf4Oie4IZPiFEpOdiI4I+oidzbeUHNuw
Yi9ZFcX4MhYlHIN5pjDKFEEWS57coanjeDzZru81kCulOiRaJLkWP55/G0k9peHX
ajAjXiZkDCPX5b/ZYjrE2DgM7QPHpFwvFYpQPomIlmIE2nq3WzafACKdbntqxJnR
OAuJ+ZEskt+/MRdSysB9PLoF7S1Z5EZQl5/JLfDBOcTja9iKut77g0mxCX+0zsKT
aAgKYtBhKCXagsjL0XzcZAoPcenvar+lA/4uivEsf5gwh/6DXqJnyrK/SV/Qne5Z
72gEfYZhP5eArr70f1155Ik3Mc227GQ8QqEzUUHHx5X2cK5CghwamHYUe8Cu4iXs
Coa+EhGTHvgpGKfw0Zp4t+dswifUeilHkdwJU8edjKoJ+C6OmYZ55srFeQV1xnam
eHe5WUYUkMdnaWTwu0+jynmfqt9gyV30gNqaUTy2bxPaQUZBhoVScKa1y0iBGA2c
lJOEhm8blmd4EJdGvJ6LZFtbqwA2xGUfdNTPWc93oCDQhmEko+80nPVdmRm54TL0
b4V8/4l9W02FckYg/A8iONTx4ZiQZ8vPltr1gIj7qNG/5mZyrZu4CgThdbGplzk9
MR5oLBFmHrfqnQxfRgl78OERKG5lzdQc94R9lSWCq4vaX66Tv7VxmVnYrrvWx8QP
8LItmKBCXf5jbRw7kP6ScPazuW88+Jznv7Zo47ZmhCsYAyF0QEi4hu+OSDBc+V41
UUJk93ilxsHWRI1GadfCXyfug/lEqC01O1KV/VR4pYwgHLtvDEcZaRgucE+rWs4H
lKSwZSLG8xyAU59gB0bOsuUGAEfPZwxnNt2azF7OiE18Wfq7JfSyaTtJfjpFWjhT
ubxg0B9vIP30LIls3zf4J+V1Fxziurc4znxenDhhzVk7itmUr7lpkp1tRawPgKsw
2jofyB2VMbB6IlXqF8CxivZVGH9GSF5zSC8tABmM8Rv7Q1wJqzd2ZyV55jNMidOt
lhbsjilO0ZTZYHX7ZxFTtpdXF2mxjV5CsF7H7/hM0g0EvcULGhj/NNlBDMgkBH92
pYBHIfjC0j8QRAPRAV5Z9+fwntGGYqhArrbUlWwvrJ48wLmSokXHJ6aw8CQ84lsU
dZpDi5Jd4TNt+SwtZCJr/rZfuPkOknGcBQRw2BQ6YxBQFf+eXWpSPmwf6MQDoJg1
mjxoxlAy6p3a+ydyLYTXGa4kydQyw2V3PaG8N/FQ+/M4MadGsT+3DMfynecN5h7G
3SGmEuAENGoQ6FIDsSRDh3HK5SMNoON+fSk+t8OrRAKGfePTw+V5fQVX4h5Y69Qb
jYrD4x7cNCKsDSOUVU7tQBaTaCDTu5ixraZ2lEYgDjT4O+DRsUriRkxNUGjscjAV
NUPTgjQccz9aKuvppH75/p5nbzNYrRNtlpSJm78RECKn2XEgqibl4td/6elDdizT
rBT/8SnOL4IfnuyyotKmDZPD3fXtPXFIRVZsQiEAPsgdHzNLMHLb89fvwMkEZRfN
SUhSdalhhncRA2pwflmD1cth5PKcwONg1hyEPo7J1hsmXzPnByvL4HsHQnVaJf/x
X7J0TmThTYEGOXARCnAmr56gAqW0zvbwV2pqExM1JAaJkroO2IV5uzlgE2WxWpyV
B9s3nDHtGvPORdixUGWW73H5i9WG2+QYvgS57kBLasGrmQPO9S11eEdAjQ+xXpie
5BPicaiYWHA+z+RfjGOZVUVps2jLvwrmvFDjKOMVIBiwho4rJd/HDBbKWsbd+XW2
8YunD3fVBWzCn7/SdHLN+NGWDQD3oU4vIzOB5N8VjY08kle7SSnzyoD3jxo6ZYpg
b1jxJ5UKWpLJ3GJW2kJNqJWEdPCJ5jmr3CPCuGTll4Zx/lIv53HSWDhhYSTNQebg
shjC2OAOlQ5eQP4KRqW/wr6DhJMpYkeLMEBepSGMEAbx0NN+deTh8sJKPOZXBMdO
QI4A3j/yBe6XPRjtNtJHCoKxFZerKIeNKoCGmAujVhpbPdxbQGi80yNnoy3G6+y7
qS0GPJypEz6cHMxV7N43lqlgdWhxf4y/DDKPPU0pa5OnpqQhfzXVSayX6dgcX0uK
EGTJTAMfhXPzf1txH7cVGUq2z2PFOx5KRifOkvpR6ruF2e1DFSTxhl7/Cuefcdoz
e3RQ5A7xqN/tJ39mI5gORjktfQvgDeoiSwAwbyBddJXbSfrMjv+jE0o1LwTt6NCl
cTPSADlNMagpAMfCsR3uN6hddNGY8+eZkTJpQBsoSWULDC8gVyDdD5c5edL965ql
FpH3wdo77AB4UQzTIddsnmHH1M1agYxe3CHY3n1X7Yik73sS3zyFkBM96AACBwvx
vIUcQ6t4BtlBGjU/DdMs2607BKhYSUrDXDq3tqOC0qyRTfkMf/GZiqXL17pcxAg4
z3bu3jB7YITO5OWt7PB/YnVcA7h73G3NX4yaxvmLbCF6He5JkGLIi5zVtJA+lS0u
hEtSOsWwFwf8Rqtcqvse+MQSxckgLdKx28I/kbZQb2yeujdo0Et/yMIuae5rlPVJ
4nMkL0izLPUYX0l5JJ5+pmRj1cAB59iMC+XZqDuRXzM/n1RkPPbD0WXR7wOVLMqK
X0WHr/8f4Pn039S3oMUXKpdrN8giGdr7wh+Q1aHXtu04tWGDnONh76yrr6Mc3aom
TDG13PADq3jodSqpkEC/M0X7VAYSH0pmeq4PyrM02HwBjJZbeSrk9xkaC1Qm1o2F
8BqhSJAOQlTRxNu+dOgAlM4oHYJsSytuxRT81Ad2OBCfn0nKWiyj+EezonfePz8G
HDFdvviWlbfVxv5Bs8+1sHGikf6L9wDKRImOLhDacqZWPuVi1i9a+lSBtvrB7Uya
srJ5p7vezgMlKL+FXC7GsGQYjsheuREAmGI0jVOLXH2j8joNbNHpROBDF2d0Bs9K
gfoU3t6HhEXokQavyfOsfoPq+rR3xVbs4G0ViFcYPbHLYZ2rTdtN1Al8jG5CTF8a
KwMRlueVjTD28HTyk7XcjuA8L+WC0Kc+BeZW24TxSnFHjoO2cyPugh0SdhcEl9Ha
41CeuoxEeqV1xHUvf8aEXAHyzzHsqehxIM2d5TlbcCQGa3fQep/+Fe9XcPnwdvcn
Rpd4Hgmo18wDaAVBhpOQnbY2L78Aq5XowAVFgMmAplCyCxV4W/B90aXiChAtTz5D
o7e02bQhPhyG3rWRlVSqSmnM22PX+iEq5hdYznc1FQkThfLLiaq0l3+hTs6s6kbx
YISIs/MigoPPsUphBs/9x4pIITqhjhg/wfIEGht9FRUumsnU9hVTqaWpdhu7ZERK
b+uxla6zOu5E8OIJwedbaBOEEvUMHJM6dMIAUXo8T4EsCAvtAauTvbfdsPHfcQmU
Dy4GYTEI8njMdt5SvSy5YGZV0L0EDYPveQfS3C/Bg5EprVoT2eTqtdK2tDLdYRJn
YwIuV9Hk4iraaauMpjxI5qThceK/krGBP6kaKShZIopEU9omPNTo2N4iMzXN/Q6F
GNeD+r+vVrUscoFFNR9myuoH6zfem0tiat6lHPQjBehMR6uNe5DfNnSpREDHSHkK
5//zemmETmW2qNvvAv47eRiX7E4BPCu40cvMpaCIIdLZQR3PJtny5+9vu0Ytmf/A
vJFf6DLp7IcHZ3Yebvn/nPt2SlPv9dYKxLaD3Fkifi6D1Et5dA81ON+qAtNiFRQr
urlTwTUgQwRVIqnXObZs2/OGWYBR4EmuQJ1yCAMHFAMfCDeio6ycbcMFWLrA6FlG
QOolN3ivNBRG+CmXYYquS9UxFeKy1jZPoscWdsqIWTHkNeZMu3kR02vGkukORfQE
lu+WR4mvkDhtFD/SwQ58U7DQJYd1AiGbqw/UxgR7Tw3texdlZJ4NdLbJ6l68/QwG
/Mt405SJFhpHE23rDVI3Oo2YMo185gDTWkiwM1ylhy+gf+2nt/5CWk9qLqACcL/B
hMLZxcYKGTufO0oHY2t/q+JSB974CBKAhgG7o81U8zQIT4t+dTPkeNq7OX28O/5K
wu5lDHesE3zj3SxoqU0WrAQ25A7fb3SkVR+YqiOCMV5hH1WSIQI8KLvU0T+/W6Ee
1UA3GcBWC3r8CVzuCMz68dgZaCbR0JQZZYXf/7MXZBaiRyMC9s0kFpORwLF1aud1
47ijcXE5QV1FtBV7V57HzzYYmbVHbT2reIy3oe6lSVlpNbtB+x4flpFrcoc0joIj
BPlSyjjmpqdSZ4XpyRBYLdt/lGpvztXaDQFfqquKUtdqpMjsG60gCXXDBQGV+t04
PUwiAEaOs0UID7L4Iz3bCezDdnwiqR5joI+09Bejqw/a2a6qaZYDtO+9mBaAEESY
z0Nyv5nt4ExwTZvzJ8/6CnByuGORj0yDFZHWWPVEnAjsltSF+4QRZLyzkrr/Z2RI
iGu/l+ggaPRFTl6Rxoirf5FZOnUx0TwvvGQlX5Uv+z8XQ0OSAyTis16ZLKk1fPSF
IOo8iC9UgHu87STlAn8umdy5YVMNAh7e6cfHyrBhDg1fIwjhGw4sIdQpt2N39OXG
2wNK/CaI2KIswlvml1MCvZloADcVEE+kxtSkJZkPRJS+6Wpqahe5VJddMSLkhoLV
OV6IlnRIuBdpc9Jy50kljVdftIv0QMWBkG9z5fA9iYsZXCnEOLj/aE1zDok75iQC
aJE4uMOgo/sl0XLD1gmYR0Gkpq7UIf+hSxIeEhMsemyMyz708TSk0ZKaTWeiIfZ7
uOIXJKWOlQLjZNwj4tiKm1AxCjrUXHDrBXsZh5j/0LeP6BQWFF9d/hpb/zKeh66G
avTxZOkNxf3w8+omKwtdYNMsHK8mHWvex5OHOEo1RVYFFSqd90JaLY+/e6bOnbmS
HJoJ+AhOXjzZJp5x36HyqY4kztEUCSTVwI2FXCSxHb+iUQ2D4TezCDoI1e4AiDot
w9N8IJNZDx3nq/fv+xLmzloG8SKRFfwHyM5F8W9Y6Da7RX0G7nVZtEvQqpyb+PeT
A7EfviYCeDENK2BNar/PnGOJC7HNl2/9/kxQWa76udoaMyclolbm81q4R++3Dz6Q
cJDRoE7JJgYt8z19OxVWc7h3hr1Fm4mydzeJqyZ9Q5TomMs6kR2LuMNnk39Q95xg
rvIEH5h+ZFTs6a5UtMGOoDJELCyhAQWvDSogMiQ4F7/WQURe5d8fbwDdXAeopWs7
wffPb9yZwtPu+ghMOL4wopkcx9sy0S3FskcDudkY1EKk47nQKdqU+UQ2nI7w7Rm3
yncW4ApvaTxwi67xSeypjssmAT9xy1q2Wqt97lnlLM/5D4No1BvLw2XnxVvxqmzw
zI+HydwalowQFGsvlbGGVFq5w/slYz/5JCd/Ja9mPgy6Zj7glherjl4lfRgiJowT
2TLMEE/YOHqXCB2ITeKtsyiJXsv4qG1aDK3zbVkDln/C7uM5I23ID4jAWmsrJqhe
Ek6u0tVNNJ2EQHfS+E1pv5STKknGKk4HV6jktek74FpfbXecGyKLk221rsXWObLX
JSesr+f9Afq4tFyAZh2YgHXAJ+9ymgzmhujbmtez3Sri8HqMsoMmxXTQu14CU3dl
AfbVQVPLfV5OmVPKMNKw/IJOhITzC8PlgH/y0W14TfF4zLnB0eDXxLs0doL+gHFq
fL0zQVjoPhb3PT+z7zKtsLbyt42qMvVkeGsOy3xafKnarak4c0zyGnAQvCtd8pjB
7sta3fnSt0XFVZ//IfrrlnyY9STbcco0g5s+QPGQaaLyPGG1nwQ7XOYForNkh6iJ
RogZnyHT51rmH0unw1rOUMI0W4LRJxVvA06O6R+rlhys5F1H7Qp10ucbZNTO0mtW
mEi3RCN4I8fjT+EDfIeooJimiBK8yBjYBDCkwKD16zd2HTZwbpyeY4oX0SKzA7Lg
Z+9Y4sbmf9Q9c4YPUZEnQFSGzk+LYZ9oiSVCqcy9/Cy9yuujG7VoJcM/L81k5/CZ
7vaFDpsXfamfWmC2pumDlqQS+EYt7M1K/zn9OiiDac3Hoihs3Qpl+Xohz+w0FQc6
MYMZSxUpa9In29B/g0/SD/FTxubgfVu4gfPxFh5kEZtpwf5MoMS/DZkGJ44cHu3U
YsoryxQun0FQAPX2+5o08Hl+j1PuthhVMBGl+CvxEmRE+3YzE7LFhXauzuS9FwoC
v2Orhuwbwzqtim68XzVxcg1OwIiSShHXjEkypkqOTxNNyFDPaSTXuT7io1WDbTVO
7BUszt5xxpiuKDr3cxDsAkujfLncTzrlk7XDkTyoF5l90D1+0+xz8JPRabkYuB7B
KyD8h2E3fw8AAaOHJOGzvAQbEQFeqd58kgihbbTi2BppGW4SeGYWLCJFrIl1YTOO
kUu7qRtjDuitA+yMuPKbK0dtjMGX2eat82AMlBRo5cKJOjk41t97+kHge21GSzkq
+1Vrvv0n3btpMOLf3XJGBwjM9eFBskECW6ooPGGLr5IefK13JoogRhi5ggj5WJKD
sl75Pk7DhdnJQAqFvPD8QeV/DNcoojPztI12DRqFbqSu10LMa2CGn+Q2dWhklabH
K6JW1EHW52kqsCKyoqRIJSbzJ2kS6tcr1FZKjBD9+s7s1BGXK6HaXjbLzWO+ymYp
mOdP1TBBoTfGQDPgFsFJ8v/9o7Cz8KO5rOrHJV6mEhQELuBItkHe3qvtABdu7QSU
ILg0VuQSdoKHEmlxKs3egKInQQB9MwnWzpVLmv9U7eDC5HJsqgKVpihSCqmeYQhr
DxRW/O7k3H3JeghTnn0FKjyGw4GGFJUaEREkkJ3IjUE4TWMVfBv9wIllak0CkYHX
FBX9VzEgynF5uDQw0xEI593Yy8qP3bvjUGzIuJMbMTk+s3E+rc+C9haxU6bjnkUz
P2sXGOuIdvSKPFBtdg/owDJwCjDiCvK2d8iKeVaqQ3ezHF0o3dteuKxwAtJw0dMv
o4M3hPnV/CFryRVJO0v72zuPLTKekYEqLYnQTCBEQwyYW4C8aKXn+hyioD5urcqq
czx3FdBnOzZ+O1wo5zRfinBBPiSbCrOn67zzEMaPA2Gp6AtqP0YlKidQDgN4s7j/
45qxL9ru5i/4JRSHrQ534AEFohgIzjrL3/DUzlD7cJUEL7I0w5o1ijGDCf7KHFGK
fWDNszUBukUnAySIDh9BWPQCAlz/Yj/JoFlvRxcOpTTBVci4zlplCH+HmtFmYl2F
3FoHysmPcSymluB4FsY4MO5DwIYbD46lH8GvBWVecYaZU9E2d+mzaQKha+FTfi3I
AqWAw+wYLKCjnCrYVAzWt+WCE8Vbn2XOj3eERIgykjVvC9Zuo0sYr55El0Tu7Vyb
u8ZNpM2Ukh98GyDEuqftz/N7mTiU0oOYg5MJQmIZ5CTc9rJgaj8nOBfEUQE10wGx
qvoSOQ+Tibl2YoPaMyQd9IOfKm4lQHBHxIyQTJZRAVXb6N4Dyru2OUbU39bHdQAX
3WoGhBujoi6xRvbUX1VQVgInq9E2S8eXSv7As9zTGCLVL9OjHJB4PLPfAISNgk0L
5rvX2KyzmhF2B+foPK5GR4nPCdYMpHGSQ++SC6IAmaz3Oj27Z9VLbJ7NRznW5XkA
V/imtRIlVoDlMSqxoeko6ZnxCsyBuY/omW/qYmm0hvB7g43WaPO1pWTw6ZvbHz27
nVgR3348fn4RcegvZjhM4xaxYT/Bv4ncG4QIV7mHZe8j1TphVoB6qBP+2UZDyNy4
8GjHvwsn86XTeVzRiWL1Zluz/7xLcaUycO3tJ8SvnR7J1bgo85kp+607VLhieJPo
7RBsvdRt0PM4Fm0AEjBrepNyJ50z/MHqzcBb0pm5sh2yJrE3WldUGXBrdaia2NUH
naxcpocp7IcDYiEnS3YAMCWkAKgT+/5I39GvSh53mebaSlRLJgT5WQ+ZONEOCUTT
hz3eByjcIUKPhqrj2w+/mowtOejjQcUQVErC1/oCFYWrourT2zCd9MxCeB3GsTRl
W5KA30grNqCoMfcCcoiRAJEahi2omW1oZTDu097kTMTetLgn5+2JYG7KykCCPxHN
4McXZ0c+GITFq6A85xSyBOCv8a6+4k/PlDuvzN64OSrjLm/6dzvzSjDrFzv1jOT1
vOwf74BevaqvlTcnfzA1X/+H/HbueQpR1mmWanrG+VYtie10Lg6uUzFYRhH7TXf9
3sqkRUXO02wb4Ekzu2xqnqEMJzLpP6PDrlgqfHj/l2eb55crOyJMBkPUkM6N1MG6
9hft/uUY2Knl/JplpQYolwXciHSlQhi1ahCnlxNb6deSZYebHRLjCwSchFAPGJBT
x0vydARBXPoDZacFZ3nwz7ytT0a4JWqlL9w+x8iKJ7aeJ9PcS3biCT7dJOOocmJ8
2NQZLS40YVtTlp2XAooDBu//ChjUBsdRl3r6EPhZf214kqQ3Beean1aAiLwZLfy0
5PNafK9AjLCH4RfRsD7jaAWE7ORU8ZgUU8H+K645Q9728q43E8+YlXFW0rOo4spe
WfWD/o4iFa4iDQNr/s5YFcy62Ks2nCGU06gXWORSFyQ9ycQuOL9Yt53f7AJlRmHF
mL14NjKyPRdZl+S6/wSuQDwQ6N00q+ZqYINCmyA58Zv5Fabd4YP9kq1x1Q2W16KQ
pW2H57aWM+VdxtroTCMRAnQvbvm7E35vHYP03sP4YwLX6qAAzi/n265LQiLiEzxB
yMaHI91cExtNnhK0scJuOud83hW40aiQFXfDV85ZH72dYkJnldzZZpRYeUY1XSUi
RMJeNhR0OAPYSc+u08YrVrfdVW1dYAd85flMwSD92NZpHWMD3FZFNmZ9fBARdk6v
SRHZqL4u26l0rY93RghHqVu587ZrGQ831JrzWMkrK2SWOsOfOx20dp8aBy6u9XEx
atNhnxs2Ib2qyWY/ZOs0hz7EjKjvsDb2LbwDDjbIBw9kHQo1X3cgNEuB9PA0a6N9
Ohb+acqdsPFFPpZANAUjktO4oaBKTE/+QRbG4IbvDaP2HkjXTe2No2x1qugvAUwM
xHnw9A1sWK3XMYjCrtpa8uz3EKzxg1lsMVTjSlXhColS6wo+hW+aI999sNjH/vCS
PreXcj0SB/y6D88CYXKQsHVI4P4K5V1g6YPwemRiXBfd31eDt87xbFMMC+tsCy83
pTsWrWyogelr8nlvGwBXMJULlLydcwx+lFhcWKlBQwBRi4xPFvnWWlQHTCd9Wsau
93GcEUrnBh67JKX8YdYr7QrIPxjVN9VF09x3XXoceLa/AuJILghQIsdIlj9zbDI3
vNkujHn8tUQJLEYktU8iL4BcXG6chl6FSPIR73m2Iw5wEip7S0X5de2ff30GCB3I
QlgsedhXnnptinTw5VXrbaR9cFm+Bv0nrIzKqwm0y2dLEc66UeFQu7HMyC+Wm+S9
cY9eVxj1FD0BZd1dIafMoSYyj3J+CbKkpAfIPLyfEBwO4w7WPbjJ81wUM/JRj8Hd
Q2gdYFQykE6k5yi7rnZICIr6IXNtOc0ljhNSD67F6KKFpTgPrUozVDewwva+kP1E
yN5uY7pBALUPVnUSdKJJzsli/BgK/S1TA9+VZtKtDghv44Vcj5Uu/oXhO4jhsFvS
a6ZPf80waL1pYUsfAMChcxOLCnjdYS3YycsMxhj5oBn8TiRzdd6bgLe3waG8RLrM
j5xX934HTn9G2kMDSPunf6qRippzgKDI4EORnEKc02VBxV/HEKt9h4uo/St3JqFI
S5551ZkITLl0M04v/0nYZmEiadN9whsR+DrGcvnbWQuCxeNqlDZSMO97FO7PK6yi
OUsSYotQMgXVbDty6nKIrxMa0swei1jmGMJvE8lxqDG4MXTq0hixNK7zRK6dfOJZ
ioteaD0NF5erzbQ/ae/gIJAAHYeJpHG6iEJbMs21f1sqmqFomOGPdAX+ko6yokBN
lwfi+bm1iVgGR6CriAORU6SghqPgcvw1oZeZO+nqYte9JdGgq77rIb10iPYKeVhb
lsVDxx5dzcVQIpHsaAJbGvsut9/XSj8wNw0MifQfmj7R0cZ5S/UFOUVXSoMpzJWV
47BXvQFog1/i8YH7XYKgA6pYKJNK9W7fAKJEpfT0cv2sbBJ+I3x1A3VmO7SJJQPe
qa9FulJoGTj1PUeKeXWuXukH42UbPlt46p6edSqnFjFR7R3uRjetkWB5+uWbQiqa
i7OwD3R/ITHy+Fnque+f6g+/IU9kqwMQBNJU+BgEdNYyOrLctYKKdY/QXxMFygA9
RTrrlFQbCvxB5yWSaETkys2qijCuK4FTS7ErG8JgmAom4KG180qncm4VjWiFaUmy
TgHj1+mGyXfLBMKUXROMV1kKL7NjvfqNEZ4TQTPFeRy6Tu3lvUlWS3FgRAyyR1h6
ROFram2g1sjgAzbnfVsQn6BbghxxqqUtO6fgH6gXdiSeR0BOYzruLXajoU2DX7Ph
CRYPni7IDUfrVUXxR4Cg95ZW/uIQuNdCqHsXw8H3QE9IVe3xqrxirHqniO6IPauL
CSgQb59uwnKMycpyZDDxXz4LrfCA8Gr/Ev9j9+fIHO+c7tgJptD1unvcfO0WFwsX
sRN6L1tt/7BzwR5wSoQ5ds1tj3I7MvhpuEzGgqwSGgHpy6+qYyteCU9qONsgq+gE
Z0J6N2sgi/bzApkeE/h17igMqNm7I+ckyKvHpdkBXGiVea9iY0kdIzxeGp0MoBeN
EfZITOqhSONgtJHi1EEtvgUbKFac1nzTIF3OYcDaFQRg8gbeaFGL5/i99drDJAeq
qVCgbGjkNFKiuvQbZ6gN0yg+/VVqZIYaEcwNBNumG11cTK2Ybm1jyV1E0v00frQa
GoWOqDAPSIX9czG796vC9qItob4TENwiSbeV+aWaY7JCAg4Wnwz9KfscQ5dw2NRA
x994aH/4L2vKWSd/cXfSUbDIlpexJleLjUmXrkislNn4+3Gpi/c9VRJ9/cb7JIp6
gFIzzxTSIcYlUtjzF4AboL5b9Lp0dYrKzKooMFo+js3Ktjl+0HBsKMCEORyE8Uh7
CCdRQh6kpncSxfl1WVKhrCuW+FM+hQP7hvED8t6QRj4VnzFSJzUf/TvyH3xaLYcF
bLmsKO/mKXiFk7Ze2dCkh9UjRWW4obTOFBP7ex0NW5oROesemZZJ44Fpg4CU5dO2
yLL5sqgMT6pUxqUhbTyEZsWMlbaWn//W9kXAdLxRuwyeOvNHXyncdtQXCJ9M2JhB
fvjkEN8V3UAR/BfR5XoHdsCHIfnIXy0oYMsMDVagphjap+QmoqYV7//XDRMT7JsP
2gMcchFZ9ApBte8gNeeFisffd/moEfnaseauH7W85qdfvyucMJWjUbiOqOHblxnl
mW3oCwOsyIkyJzEHJ8CuL0Qy8880ebjOln6cnnMXvuLwf4TdRo8EBCVDUFNKcUqe
dik2S4AhfHgUbspO+KEgMlrhSUNBCJQeyGBefTwWnqMIrRgGvK1YqfVLJHcVL32Q
o6F5mYdg5VnyNqSOXRSKIytgAGpzYgRZrtIATA8Qu0hiL59mx4pON4Qy2herKziP
suyg752xRar+DJSdMCNZVzYE1kew0fK6dnN0VuVJR9A51xFi6/ERR55Cv8dGLiG/
ZA8x3xGEtZCHvjba2d4YSfV8JB2VfWJILMEo/P0JyB4aocnQmWTaG1ZpB1pAEZ0s
mvLoNYVTpNLnMC5Xhy4qz5/b/zWCdIhDLfRR5v+NNrMZC/4dJ/2mCONDNsd5YYkY
n38C9/Opzi56IcmZgKJuuai4XdJOUZMxRVl3w4sGtpH07CJ9kuCRnldgnaLQ3Yp4
F6h5LTtdBV5mRRGqy2mwUK3qjD0RPsxHUUf51DmoD3GoUYRg+JZtYY3+3H7Sdets
uOj6h2/f/ADivM+PMh74SpxMBLBLG99o+9dqgywZiQm2Q25quO0NMO2d5lvlOx1j
5UpvyZknQFDWuyHvZFOtS7RjUBEhg7H2wFZzhBPM1Tx2set/Y2fw4s2eafUbYIYN
zhxge4XpuDxKdTFHq5DYDA5U6S5B4zkTXYGf8eYyW+6ka3DCjzIEzoAqb9FwcUzV
ql0QuiwepAYpRjZKuJobJ8H/IddXIMjcA7dqI3UuEmseGzFxNuIuEkHP351Q3v4d
nGYDmATAiPWuBveNAjKHa+EKXr6TiLanY3NOSVqJtC4hAwQP4yJzd2MzESDJlNTf
G+cpCVSp3Xxq4J361KCp8XFeepdv68kLQffUnha7pZZUjyddTL6lQ1LiYHlksBUn
CdVwCC7oHE7EX4Q+Bb5tTphmDwuBY5b9WlMP+ZRQkyiDFBMc8sicMl1VjfMLJH3Q
qUzaH9iELDBBvwPiHyW8OIcU+KQAMRbdzoFET5NyxdhaIuLSyldskniV6oifnl/a
OAt3yK9OOKCByFMD4THaPWwnaMM0faY7KN7VzGbfYTM9DEyoM7PHVUwap4nEsk3x
49sO+CPosvFoiHv5qA3EjQrG0/cnFw+wZqAftKb8ynjWUxGZiXle5fkD61Ltu1Bq
3olwCzM558eZUKZ9WQC6cIx+vW+UeVKMZsd5oIGDJjlv5dHvsXD+NHFxbMfKgK9H
e1Rmv1btwFiG6QP7luz0HUgZYQ61mpoRttcVEDnv6rZQk/gaFJSw0sxo/b4LEWsC
yJci50+GbnFQ9UM96nCAKQ8j68kCOQhHaPQCEK/q+6aOoqXnh1NoIO1okdZ2RB1G
6cXCo+EjPo3Ow03KgtM4foSm7eQHjfVFNUdX4ikRXQaxqehwp9sctdbKgtSExso9
SvLQT6hVCXZ43XLgfF1bzbwr53rqZU1fcCrcUDuteDouGWyouFtNYhOkNX1s6bic
VW9DBKeu0PoSl9GkfRMX9HbJXQX5yoXf2FkC4Ozw83pl8xejTyZV1Ad1/lhpYg9p
+Jpo1XN5L6y9xZgyfiPRftY0r14qop8wsf/bcpz6VVqMpujtMwWp0WKRZMEtWHKl
anM41xGi2hRjGh+jSsUjfuNrH6FMwjXO2SLh/Fy4nJzEPRBHfHQjSM/EqO1LVKPV
IPI3E0arA5Lfz02rupEFW7MZwspUPgl+yPO1GFLkOqSmi88Hz/8u50Cavzcpygqg
UffQLYxlm6+EsrDBxU4XfQJXyYmnt/PvYi5r7OIN+zjSNXFNcMvkk+C8ec6I4t81
xV2q3gLf5pjmS50OxL/1ishfSgF/BEbDWMTJFHzMWwS+AMOOuPH7z+McVO+MykVm
CEML0Kok5C8v7r8nWUmI5z2wOu9m3WiHpmCIWMmNKkc7P0u+5fkqF4g6tjbpS6yb
VirFBOaT2udy4jwVMDuFJe+USafHzMkoyNk8PsnOQP+8nsfEgZrzfuglJ+rpwcuP
ZJWOQsv4umOASd4uGmrTcNDDIn3oMe37AfnYNQa3RNQwl948CTqqid6UIq3FVz2O
NPnDdlhe+olba9be57Kr9UDt81awEw69GNjvVJP66vqiuaoex9uQTP8CqdHny38Y
uHvAY0gqRu0NacSQgmm+kGNR0XzCuGUdcs2Lwp37m9Ydcc3NRsvScJjr56+WjUeg
yVzHmn8VLx50cTfkddOvaVsn9wmngIXRqNBD7RRr2Q6L+EasoCAS9C9ZI7Nxztqu
wfZF1fqxm4s3j1h0qDIo5UNGlK3R4M9XDgrEkPheShzg2J+0H/YfFAgpXFBwaQVm
eQdw7DwSx6Hus3m/QMRXlWJfXzBHRm4IjyDeNlBpT3xGP2k6ment8m4J5QKRWPod
OD+X+aHd76rDQyWGp+zxoFW8P+2sz6gjXpLf9G+zZTLX4cIg7pBJho4E4yhR8F+w
mRe/mZxU+0+ikr0nmYkxCTbOynLxT8gpFmm8u1SlJUT2g2QAryc1Rl9k7TFr6UNv
w11slYi8O7T/M5rIVOQ0ScN6i1rl/SeRSFTveqUKcFbCkXKVYVeU7MX9ci05Ei9r
8B2zVDwv+hax8+ZFE+EvnRURhdZ9Uwr8CSv9M1j95HJwcVOi/EPUgeSoq106pxH7
CKIP3uRw/cxmz7cBJNC3fKob4rX8wf9yIh5ykPh7bsNYpVi5lqGptkx6OKCiULlY
sAetk8+YK4JiCdNmXhD8QgU5zbaR5Io8lAqy5+WcKgI6vtt+hEMDU6b37z+aM3yq
WWvjSqYe2kBvep2Evn2aZgVbrpamF+lWWaWuHk9tj53CGNv6TzD8A9GqssqiTuJt
o8f+f/dB2ZSK40Acwn1Q03FywbR0I800tZNy1nDsooJdS0W88apGaCSPOEx3c1d5
Dz7s+XkGCQP7EIQHyeXK4kd4kE572nYuhl2EFkSN0QMC49w86Z+Rd/kybs9TLASX
1N2PhBldM5wPpCz1FC4fP0oATHW9n2FVTrj0zkIZ8QTd19j428OKoXFffgmRrl8D
9UOYxLbzHhtZ3Ooc1hzJTohOvMxhczrsAR+qM6+mTmPHbDWxhnAgwFYKKeHCh9Vo
gg7UmxpufEQRGGfkFt6a3TTUazsLamId16lMHVYUKWuAKuJZ0RCREXHYVFZ0jJ8o
5Gw4vFqK02PfnEswxFcZAua/aeAmRBsnR4DHr78fZn1eFww+ljfJeP3yfeU2PlaM
B47gHwe7LgpjXiDk2riiW3JBfWIKGDdzGEuermZ1aVVjKxteINS4mAypN2el31cX
Ow4Nrokkn3teRCcfG7CsN8Cj2F9qoq1LeBJjQjA9P8XLldYQ955BNWfICywYcxy2
B9XjG+Ocu1HU2GRQSQwyjn7zaDXr83hrtEuKDB+KJ8sRc6doIJSAitUSJj2jAyzr
fxmWnWbWOdVFyAlUiLbsfthp5Ce+NDJOqyQXDMN7JaN7nr11dr3dG5XNwusHddx8
B3fymO7eUhvh4VKKBrTmyyjbqVu/oxD8SqNY1jU771QTb6NqIsuX7ULo8tHr7N/3
tOISu1/sz1VXfqXUzlj5Ff3Eur+5gtRuWmuTosMvIL5V9K13Ssmq9j4Cax57eX+7
I+J5bITAcylkFkO5BAsUAImB/0mRTmMaTeQxk2DH73Lj6/AD9m8lFc5b1BqkB1S0
8/9ptUM5PLSjaCcRckasGAUDx8E7OWDj/5oVurhUV1mT/cf1zMeP4GiHN66FsRqG
auVM6Af7gDQFI7wt/DqTPDfibp4O5MIVH3bZsNap9hBFBb2wv5dmbi7neykEXQum
DjRTHiXdbLac9drnuUxYlNFwC3S4I64LkT49Hopz4CyVIovJYJVTJHo0cBUcP7iX
jUQUAkpYDgEGD4goN9tef6kS7OUJibEm9SsLR4R5B0zaRJcHQ1fe+7EvzRpSVjz3
Jhgp/AEnwFvyeqg3dPfhHkjhmnHobqTHf/yab96ID9CJNJdy6A2rfh5tRiNNUrw9
qHMXfAlSUv89+2SaJ32nRJymI+t2EUs1yqjuca548JEGeYfAqXu8uhvSec9nP2db
mIXKiacfGumLSFM8heFkgSBOP5rW9XQlujsMKHL/bwuuQN/wW5YpjElhBLTxdHf1
oQclfTW5dDkr8ghb0Q/hp07dFaTj/CSa/9rL8Z6/X6kxsMVYlK8f4N3/Yr8rL/Z8
5tScBzzSmtcZubGu7/F47vxOm3qOi8mj0or53hoyPHPt/722ZXCOsyosi2MXL0RQ
Vqzi3DunXsEQn4DkmdFnn+Zi0RiilIChuVkVpZZVAJBkby2uoYxGJ/7Szgo9e3Nz
kFnCK8dbSJxU9E/+8Gnd1eGlt3aGc544RgE4NqpRTgX/ivpFKiahz/UXT/3SWpuv
2UB0uPxGZYOj99MiG4Z1GGqQokwJEXgqRWgEP8V0dN3VRTd1jwbmmKNaL2Dv29YT
8ZCHqMDd3PzWJlT0KlCRqt9yzLmzRDC6nCZCEZsPVmY+XdE88Yg6WURstrimDv7T
citvUFyBt9agWnsnSn2vLwGUbwkMh8SEpTy8m0GMBTBIaXL2aIArk39ygSXZxn9O
F5Z/bElopAv2nn470MM8F46fuG0VbwOSb5oRrM2xXlFkPNvCiTBwblyzwFFq4Dbp
oIjMQjnwIOvT4UjbK0l5dzoxDMPmLLVncon+6PmlHv1leZhYrKfQ08eQdH994osM
HAiDz7Sl3QPme38gfKgCOXiouuqFsRvgZWDEXyyGYyKRCrKAXt8TuYlMQ6j6x8Ur
bSgKJBuata1S8VnDl3mOhkCRw6TnbDb+/nd4l6YweXjAh2tbhSgR96Cu/ujz3VSj
sAfcYayQ6d9eJIMGY4URm9a5sld+/iZn/kZmohoiqfVwvo1qYvhR/zInKuBV708D
w40f1arXuYrHU2mdXH2bXKwk8MXLX699So0h/KiwFcrTTijC0Q7RxybzOFOOa4it
H/ynA4oX9SUXEyoXLqF5Bcu+kockmLK+O2CF3MRzKqfjo4RqYHuJoeZ09iKroTaq
bL0hheb4z239mUinQpR+nDvc+mwDnkAeDkTc1ChGv8VF4ta+TWjtfgDeUGwmfWPu
/wy5q4C+M+qhFeBAQH5MJ8VertYZIehiyRGDYobbh4N8NJ5BMFNCSOngKYqSs7Mu
RHsvczeLOVPzhfsKDXBdEdQzuHC7ahdcGI0w8Tf2hhCJN3Ob+ZGchY+HZEVmCnUf
7utip8jXXN15RofoFcrBumNGKw6VifOlly+k1PsxeL4BcA4mCFB1EY5m1nWaGY8f
BQAWBaKOd73qMtjrgTRpBuoOHmhzaD/TgAr9fmp3IwxgzGeF40Ve5PMjrWflsFJI
XrUJOIfIpt8423+/LjMtV1Rn5GcBlfO7dzEFauB+AN7un2y1qO16lmguVA0nVsG/
LsiNocsZRUprE94a4QKaxMJw1nmL3xqgWpU8BXryGi5yVdL4bkk9yvz85ga6cp0m
1qYZOBxOicAelnyAa9/bnECXxsG7D5cwgcxovO6BxlJcNCf4rkYXK1RZaFBX/5zE
n98Im9B2HNpEivJuxXBzuQU6vXBCdPuTTvrdSU4zAgz26kGTJzmouTnuw4ajysxc
ufGJpQuYiMS6QaFFSo6GKCu4tDKmcLRIYj6YDYPUIa86IhSSk/syIEgdtsab5vE0
moZbLpXO5wyp7bW9CLy0gcJOeLI2h/aJ4N60I52Ua3+sbEdT/GlTeNehacaSm/WM
44wjMH6qQBpkBoS66h9QzCJx2fWj/9iWsv3YD0Ys3RV1ejQG2K5QcHHOA4rcysBi
y7ud5rNp+aJQSoP5fuVbQADfymcdG0R52E1TsPl9JaXvpGfQxwHSG3ED+zLAmmyj
vcx1ktxR4jINqPWZC+ugGZ4VHBtvDG5qFtk0+HgV5hOZV1wWdhBhdhC0PwbEE9e4
y4OnnGoUqjtlLr8B19rLj0TJ4ZRZRmAkBnIs7DRbVBYG287icN66ttFVnGsua1zO
BxfckNR+ITJUuUCkIuTHPv91DzFNRb8tYpeB/L5Xkdbqx21QlLSsmhnuT/A3e4oU
lzShDnyg7lPdcNDyZ7kp/YPiQl2QqgRuCfVRvn8CvDAxoKgkqQU4hV0RyxJR1qA0
rqqxliwD7lYHxJ2FxxxZXCffQDdTIsk0vk3/ZIAK7tI/e8QsWmwLPI9mnPlUfGqy
/O7QiJThY9ZqmlH+TTiwPtmeL1IuKozXAqDXtc+I65odhRA4TvaqUFGXKyCGg/8q
/jVjmRwVYRdfqmAtKC0cIkAG1iSH+5OSrdYEMrZOZCUYm3aacmu/2Hgi1z1Xcxqb
yzI+W06jJ+IktpstJWW07g6LfWuEA+f2rydligptlrJzxREvfJ7bYHudVhsnZeC7
`protect END_PROTECTED
