`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCUinqXFFraIruqXYM/6TBUQHtXHfE6SZTwppcPs1++4+cugHr1JAJxamlmYcjzV
0Oi0LEU3FOW4kwAKHnWyGfykUPDZe1OF8ewMIEsFm7UcPNdYmmkpYK5JlVkQrM+S
GeGL/qqX4JdJfi0BmN9Ve3JZnclM3nFyLGsj5ThYds5Q8vV0dYFYLEiuv3xAJmcU
kQDl//giyktnvuxcqxvI1PmhYVHn6O9bxD1pUgiBnLXLuy2S5ENW8yQ/5x96QE6Q
n/jS4LT630I/yyH+S9SCbvXKkALNRAezBq5gPweSFHWYmRV/BUwIjXVuI0yb7Ac7
lZgi6xYx7YtSoMJhD9SSv4FzrJyPG9SYpjZ6+0e4uzY1feZAu4MbJXwrGIPfZt5R
r8kfsBfyuCoYYNGVZLgOIHfJAduApmNtIZiwIfKoamc=
`protect END_PROTECTED
