`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HGsZIUkuFSDdjw7rhpyN+rej6TPPW/yXErrb+GpHodGApkY9SPLgokB+Fi/Ht1sY
TPY4M0zU70KhDcLHlgjdIGnXFeokDW8B+R2gq5WGyTaLqBIHJ/Z0vlpGYAvmLR+z
dL+vtooWrJ5HTRGTXDrF1ADLfPtKNJsZCTHmTK/j4oHnpF7HC8o32dhGhBzczqgf
0fDfoak978EkJwYDNj5hNT6a0zXBUAdNDi0izbEtCl67NfCiI55zVq4Cpbe1njAQ
MnLfseZRd11Su1l+F42DHeQGEoNqVnkVEgk4d5PmFQJ7dKrzu+krCswk1B7b7RMI
RXpNtHHVcGUHPgPHjazOKFebS/9ucKL/bRObf1xQhFMx9t6aKAJEJzpgeszlHMCj
ZkzCBiKLq1Gx/mocgvGpDw==
`protect END_PROTECTED
