`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
utMY7+BBLYl4ZVC4xL3UzJG/TPrKl6a4MwagwWXIk98dGM9AK8NPpGf1t8ZvEKuo
BV1+fy5j35cQgVgh16G1ctYwfiPuHPFRXY3xvbNv1KX5ZWM84ou2PRvUOibbCgCY
CKXF93OEsB4ACpDWfhgohLkHhZe8wM3/B0oNI01TzxvnG4BIyjeEvm/mEl/9A3SG
Pb+F+p1tyEP4FCe/Y7gda5ULoQ1KLuDyaTxMYmSBdXeWif3jKzpHtR394hYyj6qk
2pPPfEgt9+8iPuUFQLRqzCPnbSFNrsoQMbKOXB0ltZk21Cia79LRtvNfRM3xyEqy
myJdRA1er9fJR15sbaz48LaJnhKW+ZQHHkTaxRUBzPyE3hlczVQiP0M/51cMTLLJ
vGmnfmAIJFODIvWPEhE+xOmgKnEvvPazK44ZlAhp9EBEZSRV40RrrJDXBHY5glpQ
7t117K168nNMOKTHUtyWuhWWFtemBkV/4sU62oIopLqvoSuo4uGYRX+Yk0iwvkQA
nvIBngKKIS7f5vovHi31R1Bc9QYEfAal3Pe33nmaIABJ2J3zwhlNzG2jsVA6dxSo
MGfes0U2VtFoB3Day5g6hWwAJcPfRAvkVrSxXGzmqNw=
`protect END_PROTECTED
