`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bq+J2cRb5FxZGXbkoOZ0FPTGt9mASGDDNgjqPWHK9ZkCy1XmNi1AmbuTHbcbKHg6
ryaOYY0tQQ/snmDHbYEHiUp9diyUrROp613c8hO3ePC5O7/y/xqXMzrv69viqSRJ
KxMH9COPrCRFUNpRsQIHUcza+zT2rTxzKjCYkVBfk6XmXXasAair8GxHEspoCsv/
rSPcXQb7fzcqH5fNIKmuBcc0bNDKtRFA+dlQAkvzM57Bpp1rIOESlUKe6/ZwFqEo
+MhtEM5c8wIWwp5n9JSRK5XOgxq7jNSwEH1FR1CUL9JuLPFDnPzFRkUdhDRh0UwM
8MZe4JD+ZUBKCUo4/OajKczyP22lDzpzP7fpmCdJX4E1MNXLsfG/YYCVJERuN46J
bpJPKvC0gEcTctxlTmSZqv6DuRzxPP4YAyjmf9XqMDuvTlpUW6jLQDPpSZFMevAp
bzlKtxCXgUhDilWuDSDGnWQxvEq4lAzjJfZBsv55QIxtPJLw7fZXXhpPjHm7ZWyi
D6dbCuOoP2ZZ7YQfBLqGzARrAyoqZlY/MWsm+YY7dZoNojdIa/Dq5I/Y1Rw8RMvW
tMmpjzsrGEvclQGlsla+aagRxZeYBCV7WYfv8SOL9WVoBJSdYvORrguG7CenZu7y
eQu1M3vlRpD36jaelM4CzLFpZaW5NouU824kvWOcUZh4mACoB9CMrE7Ou0Bpmk/f
vyf/vkFzTM1vJ0ZezgB8ZSP/CKYOx9tTZ5Gi4ezBjS5vGxRM9YI6ZbZlN8tzAiWU
FDLAcFj5pJqV5KpFdNuYbWQiJQruTSIHjFoWKW5YP8nwuSNIKg/EMSQrlI+HafFK
KqnUvkWXBAptYWDDHQgGuJKyg0SnN1rz4PTCOVb72ZCH78pNy4mvvj4I6SZ6Pupy
uTjEetZoBn8LK/Y3dvHv4JtDb8UVt1y2/EKZ17Xs0pRE4d7hMtpGPcQHh8QZ6Lhl
GQKTjAQm5AS47YanePvY/HvdVUjfP4WyWMhDfkINV7c82ANf5Sh+xVWwoiaQP5lc
`protect END_PROTECTED
