`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tLhuMFMtt2Rhkh+sf1lFFHXrAf5Ez3j5EfILFJRrvfL9M0Gqhi0nYVjba4ZryEWN
Qz8NCSZC8DtmXdmVj/lw7fMhqmJ1KLOzfMQWvk0ABnkFkUJvLWL5ET433rqiFVMA
Py/VVlbSeQh5SXyfk43FTL75DnWN5IuHzjEDKhTDSDwgUyofapuGjiEDlmnugEsY
L9dppHmxvoYqr+k8uV4kZ4Ybrm9Jpna26TFbfp7i/NGZZsIL9f5bzMhmgcwIWqYR
6+iyQelfr0cDsVWmpYuTwauA6hInd4kwXK3lPnY+oIc=
`protect END_PROTECTED
