`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBTiotVeoNfE0OXVx7cB9GJZY1uIotf6hGK+p9Ijb/1HVbV727OG8Cjg7l5Ynuoa
hjWVY+8qnka6QnTGaGM/AS3BOmJSLJSUyb1SW30KKXmkJfBNOkoxy50ycuhjqfW6
IjplPvzvh9tZR+aRZ+OMOs6r9ayb6f0w4xXrnIe0NV1Bw3hpu6LcOT42p2u5kuVi
+lB2/RWFzD3ZNsEv5lNmk8MdfMq+knOBhAgPjJGXQyPYKesqQfY8De/AiGMxeY5P
u3qZMluwbG2MLRrYuYCYZeiDRhWuLkVuXegbRRVOI1x55mK24A/nqwSfZAoQClW0
SukNWX88IYRmN7fA+OnHT9Z4Jaaa2taOe/KfGzjWotAZYRP0YjaLsPBxYLR7PRWc
XCPCKIzbLNZcXs0E/x8YbziOz+wI4OwGPrSb9TlmeDw=
`protect END_PROTECTED
