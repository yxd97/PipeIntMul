`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N7wojQR5f/sKRi1UGHhq0KNHpBAIu9WgLWKMxVLoOOyj80mekm51fPVnvqx00Nuc
LiZUEcFPBJ2b/wixHO2c8mspheum0zwxWbO9PLmYdnDVR76WN4j52EhfKRwQNJhG
bJyQPIF+6sDKqBqIUm0wINAkWi6z0ruvnr7bIyQ3TCDqsaOHOjYPeDP/2wK7DRhb
fRr8NMNfcuBXDthfndmRZJleIxaFzONJ+7oZZhWW/7yXpJ/tMMb/ZQL8Kbk8v+kP
yjkagbCY96bUDXcs35hI7MRP+AUVkRTHP859xd8r7AdOUkigF5yyXWvOxK7cmyZ9
EWW//Mtq8r93v7aaBP1PVL8E1BpQgzQsY9RPyQJNkSDhU+2VTTItS1DWjVoYvv1X
BhiS7W8VOkshnEjpUyNZGWYCFRQZ+rdi+AybbFeDp9YNKLZ2AgXaqPAyvKgYxntw
`protect END_PROTECTED
