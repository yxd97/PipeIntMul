`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i78lSNafa8gIpCmQVYA7jOnSL2YEOuqv5nu0hcqCRw+0ntWa/dYDwghtcEje2/C5
dnuyLjRan0QY8bbNwjk/vH2Ijfyz4B2VuwKZ5AxUQ4MOcafdCzZbt7wMGFMozP+j
5UyY8xDELG4Yy6NlZIrwgRnAvnoNZ0ikcbkyP+bEMeGQi+txWvS1MFwkQIDgg2Py
F9qqFXxLFiZNP+KtjS+oqbW85cvHr5l+L1BLPt8F/2oJtm/rSS/zrUHHwML+PYxl
Iars3J/b4z4nl4QOHwmi0k+7dJQPsO0TF2zi+jTSCFU=
`protect END_PROTECTED
