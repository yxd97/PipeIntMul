`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NGPZ7JKu2/EzCZiX6ZiWg8nHgfnmWc/al0RuUWGKe408BNvicVZAgtesHSFyhbGW
zQQlknuMo81gtzO+FPUOzSUk0Ovu6wiEbiwyukYL/1jL9XYQJB3+nHxbaF+JgMC4
RpNARb5wU9MGsMx3q3ZiGQYPAdmbjXZepaF55zY6CLXF/qa4G0IksuYaiFdLkOKO
QDOBLPeQumWJL4Y1xyHDp9Q8HHGkfA2alYM69l1rbX4b8vcJRCKWIyOe4ISYhLV5
6A3aSBTgiL/qxn3E4X24BqdYRkOuHet7wUK2HCibGaWslwYAv49gcevAMbok/6VN
UYWzHevQlJ92uGmqxgXBi8RLQm71MOzxxYYNwWyULfFw96bEihGPDkuy4ivfhSx/
/q0C7vsn03krLprCfpaGa7M5Cda1au+44h2tRFwX9hxewdkPMaK1hr9AgJlMgpSS
h26eXJbcXcmEEIeUcup1016cI045P/WdxVydT5aoMR66cMZIr5mtcH4szMsX7OPE
nMoQ3cKg0xQtHtL8WHu+sp4rnOQcZBwXHWp5o0FBj8hxEDOEf+EmYIQzFr8Yic1w
hlSOizG7hx1FmzRDugvQ5mF6hE0sygYJZbgvwu8Ur7QxxWb6nn+5SOENiMKg/veR
PaCPOuFTktShb6ZJRN+tIxDlL5yOg1dAYcQcFcVQ4+jLZ4PHcsDswnmRlhSlbAL4
xF4lQVNRYs8FZbjSss8AOHZx1o8mteXYejmQyiqg6w76gVeJt04ekvPD5zzV5Evu
tb01m4bFNtThb6HKVkO1r5wb/XztYSgmCJQ/tdf4dVy1qmYDUGECIqGvrKRzv1yr
VDoZEhKlhnGVDctkQmzPJY3b5P9Ucn3FPCigRqBblMkySv78u4gYBFW9lYdQW7ak
9HxZ7tox+i4m3C4I1bvIM/WXDjLStnp57iOyDdlFn+f5YycuDz89t5+/EdmQbuu4
cq0BeHj6WsPLOtvHgNLxbua67rLp+rdQPJZ6GirzlB9A1a4L1q3NWx+gaOD5a2He
rsTZswK+f8WN4PfZSX9vZImFbiEu2MFbHQ7wc9AMm7F1KbFPjRX3+CfyUPZgAQhT
AFjLpt+cAQ3uohDOZHqTBMYHugAIiJ+GAA35pAzcF9lT4+XzwuI1MZtA2YJTI7mY
B2Uo+NDdMAZs3pNXBd+xDA==
`protect END_PROTECTED
