`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AG5HB42sJNomWdEj7/symmj4UQY8KBDk7nyTxmcKXGatW1meDlfosLuqAZ79dWZl
HLspQJLxpWQtmd3xrIjEwnyMHKXPKLbjkfrXw0nnzvYBjTfiBeScZFz3GxTPyR0j
LH+C9XYvM/yKlxjM9TpqUz8afNJdZPOcbZ8DoLfATYIxOc+udWOI06QNFyA/XLJY
+vvdrt9SqNG4w2mMtyFRwDYSkPZ2kf+31zfd7CLhVc6Ndllg4dFGtCNry4jIgD5G
KiWSOlLoRelb9YLo4ErR5LWh3cEIHZ81kBEXidhAzyEdeGt5SM3B9LGFnPemqsCf
nHjp7UEQqOnfdOJCaMaFoxRfVsmH6iBpCJ1PhVpG4Y/7IhHIYhchWqcTzGOtcW03
`protect END_PROTECTED
