`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wMtmmJmDRrxLo7bNaLjnWAplF7nXzo35X4ah/CRFghM0jMbDEvhbEalKfRelPmFz
DrjmZiJLU6sqcQG16ZjHd6jzdD79i4dCG1pVLgKeghyI77QL5lkWtFQD7sCdewYA
ZEm3u6qnStGiroEFr76n4mMrjS7/7KqcfjvabYnaYcu4ER/WzyA+fJ6iHR9Jqo/D
O+n4JmkKMU02j9OgCl8ktMyUE2andbVdoqpK/Yem/EfgcCEzgylgwk5Lk1R4bbIG
CGyv7flQaEv37v7EbOhthw==
`protect END_PROTECTED
