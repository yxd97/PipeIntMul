`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LA1Pjcg0i0pUdz+ouSSqQkLLY60jOAne0286a5MaIt+DXo7WLxmGgONx5XZQn8Ux
WX7M1q8HTO67WSObRpx1Zu9nV4Df0gXmnmb0QNx73e+DnfO2ToSHichCcaMA17aB
Hq+fcVopOmatcwO0fY/oZAZQlGNrWsUvAkIJUoEp+1Vesl7zZzLesMdjNESflhm/
gkTYWssafGcxflsaF7CJaurKIX9ejrmHvehmZOtjPs0XOoBu+J9+rQ8I2zKPWf4W
aJq7M4hG19zpuBndu6dUmgcjwaa6JmzBoBpdTuQL1dVKegxR9PKW46uBm5eG5lnL
7EgPz8aBsLfhQS4c4C8TZfCG6l6aoISBt6UDKb2/QnuHSxC3RKf02BM6HCy6t9j+
hAONpv3B2McFp00qotpL9kQU94JCSzCcJLjJJlyRtZ7kZaMl2vZ5hUOEfh6mXNaH
4H/y4dycZFlqICeWqOm+KJxaLnyQ28o0sd+PgXx/aRG4lIFVYxqBvGTYfQmin14W
AxLeRD1ms1mR6RsLypvi4Y+c7k0mheQKpzLxAUVqtx1KKJEeach2VOXoRm/abmZ3
bSjVR1W3ivxJiUUdK6E4ORRBPdbCp23Stbi4DCbi1nnKv3pN32KY758hPEl+I3w6
p6wxl/z+V7ir9wIGm/lvSO6xYmr+DJA0TLetLYIC7uqy1fv8vIY51iX2ZCvZ6t4Y
OfLbe2yxI9zauZYleM2ZnS16lAIXM9iAmlV+JzEPhjFlg3iPGKnD5Jy9CZscoCcE
X2XxVlmH6ylI+78+h0TRlAu1payC/YJkZxrG94tCgrKL0rMObeyT+U//ST3MpK0a
la5KFKNQ6Cbby21VGuPIStqXcGeB7ys3s1vt9psIJw1EHUmAaUtHM+5Ojmv5aVMe
lrDCWkOZslQw0QVmW+z/BSXhCmPeCrsEOxdJJWLfmsfJQ4/3ztvonRrujSgWvBt0
69zKCpKQX+QHly6346ToNWSATNjHIjs69Df0icXIil+nkKt+LLacv/lPdZO6cr71
`protect END_PROTECTED
