`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1mkQYRMHyjaUa8QPcOSPOVzi956HIDXSlnd0I7bTLNXugW7Yu0uUxob12kN5Ttx
jCVzqm+DbJSs5t4bz8Vv9kUdpaUw5MAMPfi9aNEAfd+A6wAXSEkPC/CKgzIjKU0n
gubtoCcnsvGRDrv/7eYYQzVQM3GfseQVlsNCO4J2nx9VOyNefsRFGfTgkwl4E8dT
xtWAQaMfZdPpp6u4UZwXfvLg42gT6r8PaSRuGQpn7y2nDIKkNxw3Qj4S7hFD+UiL
Ywx6W1/DIWECxmTNaELvqcC7ohOC+fM75vnQLAz5rljFausMNJyNSjTCV3G7d8Ph
mm4DtCYIdniT69rTETjI5OZpGVGeZnsSMbrskDESgF3oXPpGbImU7SLkQ5/37A4M
6Fkm8j/YytJ5gTlOQ86RHjKthu8MqopglWOcwqrMQzWlWc2uI54UOkGYO1OuUk9G
xEX9oLXjSefpQo4uCwmaqAmdhEC+KSl9hxabMyyNabo6ABkDShB2RHvRBNXORqn4
qP4xNKeeWUTl5RrvDgz7wk4pL/gKUCzUJ3HLgwQkbB2HfaJ8NhsRNkBzJonc9V9+
tMc3HwLFbtwuCmFT1yL7pYSTBG2A4NtaEzBf36MV4Vpg3xyhnzaAJWPyKx91a0Vz
zCT2amEa8FWmkNAPakdnq0rbW476fzDA056bAqDFUtbI21CUgnEc6Vl8leEPJL9T
bFxkLHS0SJPJPQpcBYs+Op49DmfgYdoUlQCGvKbJwgRxOMfHG/9MeZ2V312j+Ng+
OQ7QNI8bQDDi/PuUQTIyE3LqezypbGLEspQTtq3H2QwexR8ON3xzHgsCXCHEDjq5
niFh+PyuEhDl0CSIhjSvWKnh+dGKHikc7F1bw2JvHh1xPyK34R220yYy4i/JgkpW
2z53FvQQK7x9wOtxA6YBqTToQpBNFNgY0OLyzyHF3zvu7m0uw6hl8GBShgKiPCrw
RGfb6ddMAOTTGodEcZDcMZqJGNvidx3VU1aax/LhEfblEc/ulEL6V2ghBdTPHAFA
BcKQZeupaO5+i+1/rfPOtA==
`protect END_PROTECTED
