`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOPhcGy0dVdvPVilUXFxWFzTGImKBUzOWIT3AgUtqfeVM+BIh4P+il+hJFe0iPCE
E4yigMf+G7oLEBHPDF3+Ogvc7Wrjndl114crmXKtdQRKmfJ8xK4cMMlnRldrmPkv
Ev1O3s7tlciV/mmL/+QFTLXZGxelpGFqX2BOVqEZwP/hRbnmbkt8/AI1Ue+G55r+
xYWDZ9fvrhIybmwd4quofI/H1BRnBPMrS7QiXsZsP0sIXutYsRd34gWxdYtIOGVO
hTYE43XwhS1NVfVLtjBOkEVOcDQGgv0YwEGVJLr5l/6hyflAJnlSMD+hzgkYmk6I
OnsPDn7RIdGCZ/BgqgPlkGGOdC2tGoIwG0Vpm59tuY+itsTYyQs5By+39gfCw3Rv
f4ddKn3enFvafnL4qr+/y8BS6mWRDqxijCR3eoZ8aByvq4nXx7ATa6x6BwgNOawI
UIYZ428ZKfmuMvdh5YI5ZoV6EToy6R9dSEsgObxVUxnG3t++Tqrf4hGNvNR1FR4l
3S7Xcny/Jl3zvj+UgrPLvXG3bAOqWoJ5D62YNMsp3AeuM/wlgPmWdTzKyPPGk6SC
vq3FtngVfhd4Um7eyzgN1sZ/F/5/Hw1cRfQHnJQgMXW4P3Oq+glcAQ4fE2ZvNRaT
yYNAOrHnQJwOmz2n1E7OcBtIdvtB8JH2z/0Ly8iy8dttnyhp1T+5bHxNfzF8abxo
wXPNNSvsN1/IbR8v9tKEXSIBUQHZ84ONTD4W8vCLapoDFjx9DS/gvs2yqhK2CMGF
ZPefbW3rV8G8MsF4PwPoX4nCCWkqj7c790GLBOtxS3lq7GVoS6l0Hg8Tu7Sw/heF
7gvcYzj8wzmv3gD6eULU5d9NOiDPzrxvwz8U6+uylEdqganQF8w7kqoTO8c8Mo+B
LDcpWpl057nM5R5F2aM5HiW/75e5OupL8IIEg2hARFIXU/NsAL4hCojPq8FV67R5
hjrqKEf9MoDaNFcOG90v5ZmCF+5QIt5GChu8FeGgHyebyTMqEc5y3tU/ON3NOuf8
FP5F47v9Ui1Rd0XAXPTJDOZHglFWLSSPPZ6yCeiwH3lr34Jlhf3OH6VNm2mtd0la
1mnSV2NuSyxbWAP3+1c/zmfX0dG/+eUt+tv9et6LF//Ro3pc6WhgSqzVYL1cy48j
96juLcmLQR+c7UA/vY2uyKCh1saySwLTe27N6wHjDa0m+b2gp3b7LXndit7a0kmm
9HSX+DLqM38yl6+PyEKkYIlxap3iLYSR01hoy7GEluA442uo2VqprTy0V/Fu6NfL
GZqSeNuBPXHfiR6dZTs4agw1GvSxyLcZ70Q1HDgaxwBjHXmiGIXOULMgAHde+YMY
ROSAbuJ9Jp5givxw4lBFQMcpC2Mc5536pLeevY+7Tcmw/xAXXXyX2q97+Rg+lAsT
OVTsB5HVsHpEtfG9j8Q2k/b/O6ecPVUoY8v2mmNBqTa3pH/pS/tSax0+ZpOeyATb
Z32OHqz4HCKsOBdlPY6vZXk7Sv8GaATGWiGCm/uIN3XY6lBAKylI7AslAduzLetD
tVti37kI4hEL/YuJVSx0MT4Ao9qJCRlZba6kwqL0CghDBY3nSoLgVWE6RQhKrydV
526OjfeMivBTvedmqvLaXMWu+7f0eVidDF5hSR9shBE/EZ26265zz9Wffu7vKSuG
Tug2Uuqp3x0yzjMs2MbUfDMMd54cwC3l+i5EmRb6ut3kXPOmw13cyc7AwjGCchM6
3ZUA9zW4hmQP5Fq/ehwIKn2SGgnCLdEmweme1s23nPTRFOp1Opdaqv3+XQucZYR0
r1VI2dUUqiXzkfA3PAf0BzpUsiZeRzX7eBsj4R3VctQnU+UcRzPGLYKndW40MykO
qEZqcAS0mvBY2N6g5Kzj8Ipj46gozI765BTAHGuxRK64KCEFLKNe0T7ZCX4ZnYHO
GVpv56qhy6cyCx8Mz4dPX2YiLuXUK9srQ079X2v20RYTb0Tf1tbOuXQHyp/CgEnQ
0/KG/VN4p/H4alG1UNKEQHtvzxELyX1eX5UJ4n82fPGM4bylg/WfTUxVOJcauEVo
sIWHPDZredmbUQt05zW7GjgibiFK4broCOdhzPKYtXCbe9hmHvNXT8sVjNjwYgZo
RQT/UGoj/4hFr/xsc8+Cp1jZEqpdTtr4+b6r/cIgp+mT2hhmTue0+J3lUXkFfAkO
9qcX+l58Ke2sAt2ec9RAcj1JeX3ckLxCq6I2eWJHyMLlrPuQa2dl/rGkhNdsBA8l
PbnpTzfIIDa5RpLUI/GYwa5hwDO/t4ZAOhqBurmi4PVb2Rj0BqpI+9nt6VD7tdgV
4lykPxZ3OXJE4ds6kkpkQVLkOeLOvd7H9PKJxKQDbjzIXO1CDg8GXNhFEJYAu2eL
Em2ivVYfEr+LsxCoVI+5sofGCYpDp72Me9BkMoAoLfweKH6I7XHkATmvSiUnkl1E
41zt5q5whuUT+F7Ner8m8z/SN8e8S/x4+jALVUAirt1rjet0hWLBswYucfIR0Jer
6Pj/y/RPVSA9o3SYFGu+CF2RU7r6+KmEYPUEkoVqQq/R/XIXK22sX1SAROwmPQCo
2ow4I49qBM3F8jScw5wxDojYHGmAuQdjwBAYuyjmWw55o1VnNLrvbnd37e2HbF/+
AJJFZ1ff7AadBGM5iD5FczJzS+5HE+dmQVtzdtWCbEsWDB805HhBXibIWUI2xYdq
q3+KTN8XGXLLmcM17JODnhGr9oz4x4RrME8JfOisW7vV1u9ZmxgPEcfJuBpf4zJ1
Tumb1BYW7hk738qadAMBvpUBKtRALXZRysd2tEzH/HFV3rREp+MDsfs2O7yQ35+e
4Kl1B1Is/9EajF3t+SkqeSeNHDv/1Pv7UMmEfCdavuzntxQCJF3Cl5r+oMXUoSpX
n6Ghde0tmLR9up64cP9pZmqttVV612NjNrTRyL7URXCBN7m+Y0I+YEKRF3HZ5/ck
SLk/G6ZDruH4NM63g+3YJ5vmsCfWwt1s4CdL18N3NLXowuYphtSKAzAn3vIokmm2
4g5FRehH1ejm0SYeg/1HHwBumIpQbiiCPSFllkLscs94uwG4io8Hzc2NZPg2QHw+
ikJ5AP82eVLWlZOYiPT8pz0uCJHL3cYFWQXx3GKbnTwqQQ+mhQ5EgOG5ke/GqSie
Qfu+ZegkOk9+O5yJb9fuV1S5bIfZIePbkwnLSefZGGpgOq2Ty2K9JCyMMBqUHW9c
YkLpLxw89dnXsI4ugtUSiMlutjXL2ioWnThJAl4koqbH5mrE8UJfzptuj04nm0YS
9+3nxzSWeCIzp5/gXOZXVjcG4T5Bq9ok0gYhmnj/Cru8T8PPNUf8ek3svxehhMlR
sdruArQXuq8y87GFJp3CYGPJYrslbU8ag/sWcTiYVox2fe951Im0xDXidSGTc75h
B4N+zTS8lk8ZLMbN7wjwlknjtGfNs/BH21tPc7zoPH5Hzsb5L9CKsehVnhasXQns
gaUHjSkkSJjscZGRws4hr+viycPIu4DYj7ymK+YSdtgfcHgB1yFpVDVpLpxPnaRx
y/3nTdxtn162ZXrUAVo0Tu8Sy4zZVZBUfp2F0IWjVSwUT2wtIuSQLJhXnEfwlJ1l
qJcRjeK0GGj8vMIYymoQCVrOlNRBbAPfN7u8E8c76XJkW1C0S2EOXw6CUNF22juU
Hpg2nGzlbJIF666b6935y6KLshiKcFaSRTeihQ5BhTqq3D7JXaK9fKvGZpYc2UAV
Jt2qiWqeb2SYgCYyDIxPW+C+VcHSRCHPbqze/gtBWDrSL8w8zJ0t6FJWvgx3YzPD
ZxkUSgd0vuRl8fRFWpT7/vgV/zJ41elBrescAY4k6fCiZvYK59mM81afdvt2lzNK
XGUvfmYbCgXZNPbmJf0RPILHUoPHWiYEVGJ7gyWucsaBs97VfHjrg/vh9Tq8GOnK
610bHcqX2vuuRMYEkCBY14SvdLknIP6ZALfj0gXLehc+mIJ3mNbE4wLdfCowd+NO
JEjJ0kP9y8JzDtyB1DWMzc9fRQI+3aut0aYRsfS+R7KRQwXX3XjQNxb8GDTxRP3K
1mCLB/jCj/pq6T7UvLVGjyhDDC764XrviXTA0f9y8gVxJ0CjDyz+aWM4QCPWnf9p
29Cv+HodkAVwCw2gvAGfMNit4TH6/AcewqapJBIr8dO+amVcZbL9A5q3t6GIcVLJ
oS9+7X/ZYUru7xWIjg4wuUkoCy2Tltjp7f/2SOmVheN752QL+af89A8zdoogYoi3
ZDjZlzQT+3FaVTr7axrllgQF4wJPFQ3Q+QpIcABx5dyLe3lDc1Y5mGbP9KblcseE
tpXraDKdEKsJ4QTYaR5E/aWgXWko6fwwgwuWvGfBtL+/eCHABK7E+r1R5LEaxwgh
jteVsjzIfHhWpO350jgg7cPbk9Y24+0Z4W36UoaYcLyr34+07YtVGnGG2JM1f57Y
f7lmw42LIhehHumE1QBMFv7hfuJrAbfc7T4hYcSHomxAHQ8RCKOOJVcIShSNfpXf
iasdw/TLr2BbXIgLzDxmHdyV7/UUhBkNDJdffh8zoD2H1f/YCdxCamX50NyVWZHG
LriCdW0jXsT3dE1JIiFrSr8C3dv+dkygKss+/L2XR9fz1eyW+mqY+c6H5+iGomSu
oPNy1p08+Launjj/bN3oXI2xE9GCEXADBjOsk0YcaA9QPmwY2BWGYK0ePrGQb0tI
tGncQYXw3FOnoQGOkoefZQSvuHZPIS9BUlSA2VGbkWovgypPvWtJi1SfbYn5+XkK
gK3gZepL4B8ejAnOSIXlLWkbRLA0Q4qQcQLKpYeEzrYRtFwdIJhmxV7wQCD2Hpjx
pcp44DrIOvALE4lzJlWMpE2WgpVmjYhFjMerOZDLZy/MILDO8U+qg0LPXkwrpmTC
GUSC65LPbj32ORRmwMjztmOFieV3DDkh1wpyarKwGWleBdcAVh0vJb6B62FMh1iz
rHRrs9IEq3ocRJP9bnBebm0y15dlqP1eJacyhPCNIMKBI/jy7LWFWFYmHVDDVHsm
HewzQPjTG9DMtewotXl0ky/dbc7nGNlMmTIFwYdORS/ep4OJd3dZ/aajI1H41iqf
H2wvbUwuSWoHf52wINzdpqphUFGdCBWipAQUXEi2NzE2kednP1x9gknTW7BAHUnt
6sVr2y2GfDF63UPn+kd/eYzb2IaorMqHhOb2MiSIC5vqiQSdRGJUsM9qzpomzHin
YWYtfGDwVFr/Fv8HJAFXEpCZuoiM7t/SGEi7DB8R68k0o44dBFX0amDTffqGkLPe
V3FpVukbMp2lxawWdIYwf959G4ojPZBwbdA7RQJS2TvAVm7yyiQBuvxInWOH5x8m
FWqCfiWASVvC7bxOwFyJ99qLfvb/hCtkq1l47yiDA+OjjzW/q34m8/L0Fgzx8lKL
y45jVTK3WcEkMx3WvUb/ijBkxUZWRoAvNaKdWUJzzO4mTU7xWKMdxJtf1AQ14dso
Q1GCi0YF5BIg1kF566AKqZIBJkkOUKC1+5hXMqSmErqsTEVjErlsELed6uVDDvfY
LPaMpehvlHornY4QWlwOz0ywZ4Y0oD24Y4Gu/f9Y2F1bEMXUd3KXTF+RrCXU87te
iPu+SM+qXW4mon7QV+HGrKX82ny3w4HlPPKQXQMMsMXh/sf45KXRY8gF6+bRqvFr
aCcN8Ih5agoXh38YBWCU+2CXDMnfvv4Nfwc8mdWQKx7EgEagRhyBqyM87lO+Y8dv
fTqntQ7t7MjJbLfsr8VXp4uWc81jOviT6nSxp9m+RWqOA2Jes7dhu1EEyydWihda
zecdYkXFW5KI3arEgv2ptKwGop9bEKQcjuCnJhkTJTuUXn056hDCr8tOnOl4tc++
WfhWYgs5oPC/K5CcSG/YWvKXHpmKGjbZQaIAPEg2y3O8BEYKdN6cZOQ+ZsR0+d3U
z9RTIvUlx7jCAFrSUHbMeSNCVNjTlTXBuJsnCYI/pyuprCkS8rPwoXsIvDvOY7cK
ZacEjYSYgUj3omHOLyNYdXyv3YgyPHq5b2AU/6JM/FU5UKaTfbh3bKYBSxybTOvD
x+ze55Ncsd3Xm6D9nKCjsN2lshEYAHUkpUmRYyc2fSzWSTuLoyTVH+Fb4FrBZJEx
qzbO+UgPbXp43OkmPCOZYj1zMfVHtT5IIqOV5Ke8JIKGzlKNs0pp0e+kZpn78n1H
aZGsBzE3tshLw9dYWPputMXrW6d2nbbki+l+wpW75nr4Je/qKjS85WJTv3uFgVp5
uFK4xkmbxbhzQOOcbvz5eqLgdTAWoRmFG5ltwJqidPp43/FsyYwNyH7GmOrGPe6q
fiWBtnBwlQUsmNW0uN0CvVK7xvGh3Umjw7u10HpKxloHKuZh3LfwfDvoNMpCEBEc
zFqeCUlRn+1nusGg3WlOcbG1vlzLZh08KaqQtYu63C22nuwGmiRVqsMgsAzaJhhh
QdtDI45d8Dp676yiAp0ydG4WxLF/pLi7uOwr0DQVVOgPXCUO7ZaLGTdq6kieg56K
djmR86m1jJq0PjVSJrWxho+hOB1QdxRVJ+56gvv5YMLX42JgB5IQB5MWjDV048Ph
7fG6qvSLxnAlZXcpp6ctdrSl74orUz4ukTgzN+S6RBkAOC4tGVyzIbooXC2V1ImO
xBldhzxwE+wSR9P/cOiGX1XBCfh1oAWj1LITpusir1EBlle0yC83mtV+ajYgbJDK
WPKdc46QmSA05hbJHvxdBopvjHegiHMWBgMbZIGYyGQhvsN//AQsUOnBLx6zN3PB
x6O8BtiGR+WwiuXh/WfIpIRX1f9dI8SjGF6ZMh+B0tiChJmdjfJ66pEcl8QSuaa9
MxT58SO5tsH6s8uJ/o09/Rb1hR6RI5+KYDLilIVt5qpNTpjkj+fPzkOqm1gqC5oh
d5NZA20vVtTALfNsSW0KNkfPCqJkKWRGKSsGnLxmtBwYZ+cxXDkoz9V1w/hUrlf2
oIoyzRTzzrq22cpFfy4yatbIQsAzIV4hzwTj65NJZXKJE74zdtV2V+ycMmCvNAkV
xYrmvyr4nBD9rIoztDS7rNoJy069hV+3HdowhZDk0z8o/G2UKvJTY510FR4digEn
aRpc+gRzCthE2FtGxSppiDyLFSPzExJOXU4mbVjGGjfABjuVRSeCBcJ5+HL5Nqc8
GCiZ434jZkaVVlDIkcb9/F3uyivPv9PBr93b1bomjV76ujLBhSTG/rXpLtcK2qLp
b1ffoa7xb4vsAAJ1RQybHU7/w3O0yfSc3+p8EKpITa3fXrmJvOkkHsyC7xOK11d9
p8ktdGiotZPheYFFvpT6RFdDEcxbolG7D6HXWiFrFxiV3UWSni27XJOx0Iy6Ps3v
KOullDKu9GKORh4/d9SDLE/b/EVno+hq6kHc7OmN7+bcD6KRsrslX3+jcU/4G1+Z
+iowTZP8IfcYrx1hO8hG1Rvr80W/c0P01txRCUoLx4aexJvs2U0nt4I7ZUyBaDnq
Gopk5+LOXCe+hImHHaqMqQzx7P+A+JKScASDo3dKmVrcNSRXBQF2dJTuiv1QTQgf
ocoL4mHQGjEtCVsZ4qpOe79AIClXPiYkiXW2dx0fAiYDINZ7Vb1QkqvGL+oXlj4E
LSNH+0rEsyDu0p/OIJn37PKORuKuSVqrMnDncyGtziRh5hqiFKmjEzy4RsK5rNb4
SdZcc5sZNWSeT0HQ7r7CIvCE6V5BHQT8rS9yoIzu/r9ZV0+IJtsHWf4IKhlm7TK/
QQkwwjLE0JIkgRhFvKMa9SXQY7OEuQnNhpNIhr2e6pyHYin/rACgBc7810R7Aavj
2yo3bW+jrHrBte/rghMswGNwFPHoHmoQsoqR30uV+PApbGW/zQfid4WnkIeS5D6+
Cf911Z+qy8avLUEq+Uhab7loHZIbS6B+OHc4l8W8gT0l0lMzOjHMTTjobqOJljjr
yemSy0QQSlaXCMuFhRbb4JytERqmfqQtkIy4iJsKfGggb4tfu6HOET0oeFGyr7pO
vy63YGIbmeQaqCKRq8taEQJ5MUCQYVnIbCDCcpAuN1mB66/Hs0lkB7FNdiSm/Xr+
ZqjxN7G0GdETZzcajD7ioVPLrTHztkKNX1eI2Qzhypuaixk8kwVW2MNvIdIhY4Iy
BxDvwD4WZaEtVpmk0bW299MpN6ZPysphU03yf079XEis72FRjHcyo3DgQoWJeKPN
X0aE4l9SPtCz3YIHG2FplE2VTXgRZffXRosrYj66y5hc4ObIy4PPELkdOZ0E4Qv6
t81BNdcYVJGH2fCrGlc3Lv9v2JA/o2JDXIkbjyJqbfWEaFGKDOTnzkjDrizNq+IN
Dkh/rwutOpjjEfXwfVQ7cN3ZYntAtHrpPJfLSIE2/8Vrcj/uPI7CcOO0EuGGwUzL
uMt+A0QsdSIPX/wWOekQL6ec6UMcx5EuAzbyNeYPQZ5ChTNqxIXx2iOqc37HxpIc
MZChvEXmsURu6qcZ8uO9Zx+0ZWEQg+IgZbsGIPSRvIa4E9ZPY2+CZQOtRaVB2YR3
4vXhnfrufAywO5N13pbVZHiWUXIEQfmV2/34QILAfuEayjx8YAA/BCokj+oZKuBm
cMl7GAl10ejMhtf+R1Xws/94KiPQWrW0K7UAAVSgxo0cEueFFIznLxgovoh11juU
5LvLChA+ivAhD/2xVmRBQ2P6fvZLeY+i3hKYabn77pum9SnMQgsOvlGiDHA6lzuQ
2dyAOmtzNhZkQCLwsmoXnRjEYYNj27B0hMOtDLZbxbXMxKcBag0USxU3skIHzvoA
hbns/UCu+rE93HVIDlh3qFWD4VJS4lUOx2dO+DBs7E0enSGr3LTlQnR0Po2FIDeG
fyQHCn+dT4ASr4MfDDdJq0ypF7qeOCEsCNDwjugEdcuqZno7vHqj/4h+xLJi+QUx
KC5jRN+NCB68QUaQsk9BRsJuQHokwDlhFawzUjX7gcQ4Su1f5Y9nSlc/fcwUedoa
jzqDPtSuQCj8dFAADKvfwok8TSLeNSgqiPW1yeyollAOXyzPV8hWfGD5tOGnnP4I
3KKvbhSM4OtoPpIO5LOeCefk3QD8aVe30xO0HE35ZS7khgn2J3iwvwR1rX8QellY
GVBROMLt2YjxmhLQnh5uYGr3VWDGmgo41mV9xVntdi2Rq5GIlxupGOzUzGAUjgUS
Z3Nb7XXHhIZwSOY0goM+5GJ7mM/aahN5dvybCEZzZPzqyxTTLKCrJ00M+g3wGS/V
QkHgDFqQsVVt3PlV/6t6iLKrJHk4YPzC/qQonpuo9R4j8QzqCrs5KCM+JouJ5cau
due7mqo9mTGRi1s0YV5eXzPu0xygRwrL9ciTK0Mka75La7oayMeWrHimwPoNROAL
8YP3OG/lmCuvnE+nkHw7wNLjGKslyfDnjhlSRHPNJKeDeDHZfNvNol+FgfIV5OMa
zfMD9sNzMwU+o3kTuz7RDcY62EDs6dCXCjT0DbQ4e0tjUW6n7S+26qBV8f5fUs1v
sIFN/9Ln7PS8Os9x58zLXn0yx2kXQYYY+mLqO1+der3PofQE73iPnIHzYlas7SLA
x/NNAJL/pk3+KtJyk803YOiwVipuXPc60eod8O2JoGCdLNSAAkUiOs5qiduWDA9w
RgHJY5lkASsD1iHqz8DeHfillk1ye4vOGEA4h6shtwEqB8b0oydq9m0gRE2Uab1G
ryw/vovjTfd4Fx5pqro/u1EFqn7cBeb+iZkBSbXBJR87dorw236h1kxZdb9fk6iE
FZRzX3YfyMBPdoR8brigZRoILiBM2s2nhiSrsH/bOjLNl+T2Y84NNdMvIFtuCuac
Z7mqNOtLZ1L0ST3vEkN7MgWCGxNw4yDPHdYXTtNzbDf28OO4++NeXfe53ilR8IJI
4ES73+LkgkzA46/4QCA1tJmzDdpigzQvqnVd0O+rhfGYuh3pd9dVlDWat3UU5ceZ
60lvoJZn2l1LuWEgVAhsNLE4/YGQc+LZ5bBNfghZOOfgENL2LCBJ8i9pKAQNgGSQ
uSuZpkebplzT/bWCFBhVoDO/y8SNmh5K/rJM9/4G0IlbGiEg6CFATsECHLQjy1VZ
nZNmlg5VXltiv+FXnT5/EjNN+Yj31puZWxBKvKKf/d6GrHOhU1uCKXcq41Ebhyc7
VmkYXDuIvLwMuXYldbVp1l61wabhF6PT58mzxmrJD0H/VWWtvlQ2h++iAMZ8k8mJ
ppM33m+dET5W3qYcTI0rJYXMIOeVnftN6jmcjwXHXHN4gT0jh3c+/W9JhZGVphXF
kKl4B1PSfoKamOKAKuQp5VeXh1sGNaw1nwL34DxUuBBVHyEjG77YCrW/30rcZLLN
a1+dct1iL94x7F3CK+DhEuPazs5QfN6kaVWOnGY+ALC/yw4AtbBSILaibVot6Dxa
PtToBG7QNFpxPz5fqK1BXcEaezVoDyvzgcglEBPFBal+FpCjD1W+UbFAlWGrjtFF
L9LRXpGYbhh39+eWaLfRW5+9f3y0lvoMGKpjHx5jm3359f64NVZaMskkvAoXLml+
ffNmEvKAAOyN5bGWP6wJvWwRaSt7s2czJMkiAkSe2+z21bvO8rXgjf52KCIgto/2
UYhwHLqu7wxhmYshjXjxBl3wXNBtkZs7RdowRCOg3ruTlsi3GYeQbv7j2iCIHD8F
J9JrerHn6o3k2vpQhRRoi6ruAFWGPmVaTj674f7XuYyhqkGD/6+vciHvfJ5L5KGl
Kr47irTgH31sfPB9sQ+5GLQWxwtTm8+83R/SYHGOiXZUi+gaON5wD8JTfOoXLRkD
47AC5sSQeOKEv2gAeM2ofy4wcBNDG8Qscg3JNxk6GITK4mErt9H9L+7eUTjElcLy
XmXYlXf27Rg1dxtWxAqVmM3+oBw4QJDZS4yNg1pSiVNqpqu7WMHqkKLjuOe/FepZ
uwTOPQaH12rygwvseLjh1MySuR7D8DArcfRCd2aOE9CpvRlShhYsTnSAHsUAVu1X
MgbLypatqTjYd/7K4f3Jb1TzFIqj2bGkAecHGQxsEGMvjyn2Hw5kG5JlefSvy1Ub
0smjNWQqQc/svAmrZzOILbpLw5UV9Y7lwsXlFewDqrL1ehki/Rd4XxEHGCSHp+OH
aNc8RoANoYs4DKZpbyc6cc4MoYQ5THyXjLsivzU5nHgSgo1Fcaa3yFvYQcGWoEfg
GAVONMgocG+GV9wRZC03cFcfCdBztSeNzgpizB2BGxu4MspJ7k14X/rWqTlqZBkp
cUgQ2IoIEgKPxkQxdPWRBP4cTpNKLeN7a9C49DOk4wkKk9PG/H98D8YgqHN0GEo4
gj+MwsswY3WCt5FlSlQvMcaXlQ8xADivV9YIenMqwAiAHPBycV8LK8o4nhS8wwJk
Mi8dcN5A5zfv9vwTwJ7V9teHOFWbixRA7VELgdSFsMDfk8fNqMHST31GH1oKk7H+
fCX3wqLtftuPT4hY1Hf7EY19D0x2HijRZFiGVsVWbwim/22bxTzkKR7yE5H5D4T7
GPBM8oMdr0SIJJxoawZ4QtfUo5GUiNb/5dXPaJV7UmpgybYcHpiMe/SeP8vnrWC+
vKEnieJ8wno+cRePlVUnOP6zdnsXhzgj0h+lqhKPpJMAEZABsu+zN8KlD0cvchkH
u0Ha7hSmh4OLx1SR1zgJgW8K682uysXaIGExdlIt9NgG4hJiCY+IxvDsx5PAj7Wf
jB3S28TtmsByXa7Ox9KRjQiaKq07KIwUBdNnqvoX6nBsDSC3nBOADEwKVKoege6m
khcRsieSTTJfoaC4IY0VuJ6Zy2i3Q8eKJcmv8a1bTDZkh5x8Us3QfhtxDIenjhjK
KdEupabIO73cbJ8VTxxdAnWCmHOlS7gJzsUacFQIrzLidvpRbLmOoBFMbrltfIzo
Qjzny7NLoO9wkGH4ncOaw9qfHyclhLJKIF01lvNzOnqmXq9plGwFXvaHVZWiqlIt
Fvv0E8OGC4JziLf74CNOsCYjCPQh2BqxOuYWCCf9thMW2NsTgm8f2U871MMaVRuq
QwxPKJxc0Q1RUU/v/bUu7pBvjUcA91OXPQ2bKHEwQH40uwiWmEnynGkEIChT8EXB
7d0BZjSHS/xzzw+ZtouqLDb2QamWKlZ+Btv6eW899VCtRuENSBTt7YrmHlr6dZff
3YZIcFsphvfS14WM3nEriv43JYpaJ9tZQBk5EnVNFpJmhE3IVRE83v93E3zj8UPO
NZC5KhDh8/Oy+hwhTewBn49VpG45PCjpDAr8MBuB6f9zKmNqBP728P8ysWYuWFRZ
KGp8zFtrISGtTpR/wg6YbfBx8PhUmQcCP4k4Ab1E0t4xS5irhewKqQGjhmKIXiPm
lV+GVrQSU4Rb+miLXEeRuiRNu2Q4dEVTdaSIn0rCpMXKBQTsDDwqURIk8QsC5zBO
bBZYIHWlfqOeh73RACaK2DXTL/1i+hnbjJ9Oc+cFc309Sezmtn9+nmWU/XQ2hrfp
aSpTRTsZczel/U76GMQ3mtSvxjXaRakdRZ5dFZ4gZvYqzc8D8//SyXpL5Y+dbaSY
plxpvYBZyyVtZPYTGmjPO7q0ILvT9HhbKIGoAIdetgDXcxz5C9iBa+R0JdKLvM36
zt787zg6lAFPT1QrfAQlqMJaU23DWNnpQqonHz/tuG4vpU+Oqy1ipZNRiphlOBWk
nDTdwvRqKA4SElHtjHeiUxfg4pMdZ6vYE+wfXPrMw6JGZOHAERvODXIpPM6nMJfe
CRscZ8R2IIN/BTiuIc7pRN50AeSkjVfTeDvoGSCfEDIdTEV6rPLmii0LXDxdd2zl
bUQHSYK0BgELzhOSFrbBZH2I1YCG7ocbe7I3icOGWyEy3FRqpmUP8tOomPbK5IFr
cuC4GuanCJrKYwpBRPj4uv+B7/+JbIGDymFYDqtXgLy0HD7FLEeEiEf1swCmombf
FLcB385REzZoaCAjxwzIIp12uRrA3t07P3StAB/GSZVHH6CMJAFwscR9Ea5JSILV
RPS1w8k51Qp+2YMIQFQAKUZt3aKlO8WVtOXdn+9CpI7QtaqDn9uoWTPQv6qy6GCz
bnkY2CBhcppq9gRYxWEmYpsfFw26B5qUHNrzt6R4pcEahijvW8M2s/1KUKZeC4/4
9pQT0Rgd5+1BiNs/2jrSK6yCwDLcoNlGj0QSttuM3eKY508dfLOCfQB54BcLApKw
eSBR0sRqTgHWQ0CIrJ6hFxe38DsSQLDtWg/VY2BMHb8U4ZNaTnY/kyhN2gIfxH0u
wIi95B2ZcG6Q0fGHA9FFQ0zONl4uEdg0iOsX4hftEOOD3Wb/rJSTpYuL13pO1OyF
eWuo9ZZ3kNYCxuK5JHSklvh5/pTponWbyW9AgUzNZA8debxjJnCYontOlHF1vsN6
Zj7CEo5ykl4TPdapzzcL6uuIlNN91T5uXbW7Bk3hKr2S+0lS4YLZsaYUj1UNUW0u
lRA738Qv0qmvD7V7NEAdfFqLLsa06HoafQcnBQa9IycKqZybVCicVPG3VG8rrDY/
1dY74krRJ0Z6G/HXPuTr04NffHeRXrMaeNhMQSGfQvrlVSJt+ItIyj73Oh8hNbex
RpiBT7TKZ3ycjYQmK23GiM0eqOJsKHrnQD8+SWgz6tZTQfuWegnAYT9koNNYlSB8
Gt/4KucYwUq17//toqISGv6r0QVwz6IFT46VPGJHwzKDMcDkqBjf2LuXXEEMUDyx
sAtitNDKT2xh+PItS5K+yeo5BG81klV9p2ma+mZ7ESOFIdGqH+UV1RVxZtDok19Y
+hdCBIB0+MB1l6dh4GbVZw7tWYtITHnxFr8OGDfgZLNhYBLBqEvpHxlMWoH0RO8x
kRZ8bnE1bkgENgGfHUuk2GZRy4RiVukJF4VXMiykVe6rkYaMb0365q9LAbx13RxJ
rWjTS1DPAkGKammOVO394g5Pm7RpxRt3bA67zhd2TZ+Gi2T9Cy0/jW0EhlGohiTn
iB9rB5AbneOdZRMNeFHJBBpbEBMinz53Cx+YR9AnsUFCzoEJt3ZTG+pZoXCTf1eC
gstBSsX46199A3mjHxWF5bEQvBp/rbnd2LX762c58W/Qz66JOcE+jzmyMqXZlAvS
G//HMmylPOZPkCGOXw0z3Srwxvuxd0ztx2H6z7aQHrU0Lsj7Eo+wt/C1u/z3yM+b
s1Zh1XrzVsGQXlP4dZLBtRF4UuqpQFB8Ge+iQ9IDqDfsvzvLWgMWmV8Bhj6Pu5ms
O7hBNMtVxN3qZt9bLk1j++BBn7y77+4BDj/pJw8Of6r4qpP5EsCjZFuf55u/GfSB
EuWYSUgSqEUVI8nPDBxzdNl3MO+9HcWMaB++jT9MSrCWefCceCs5n/1Zvw13WfpU
8Xd7A0JECw/sdur/V2vjHuyMV1ekvo5zEXIdcyXVXCRwXHKEC5192L7n4OyetmW+
jdozBEli6wYXZRteHkRaRaryZpaUxPusQ34677I1lwTvX0Naaj5APgUVf8KXGKcv
93Ee5IwvbhmRnMxgglb5MSbRIg3ahgJNcvQk/uU3hPrGvLMmW1uJqHOCnNX5Yl+7
sHC+ArdZDRW4VRrwzvbv+SP8CkK2XEylpW5T5jL4aD6KAhJrPXoiYyLQJac/wR4p
IDxjxcBkp6aVCd0AkEAlUW1RcoSc76VAI7GDqf43lUl2ocqek44YcsV2ivzugTB3
PYU4f64/OwgGffc4bymkLv0ZkewW+mbnAM+WWUNjOw2UWz9AonngS3ku3OzshJjc
1mrfScSfcBeDBtk4cpWE2DQ663U5NHuQSsJiAQxckebNc6sjTPW7QioyBMC8Gw67
pm9C2eWeqefX/wCPRNzLf9CT11URUEUBNrhlRHwrYfoW51CiMjgEDBsLo19MSQfs
DB+bYyNazmVIL6uXh5ptBZNM3BCbFAZlYorQiOHyYDzKDdOp65B7w8upyeqRH4ob
g7Qm7u09fyAruW2BmoMipb6JP6A1iHi8TtIeg6XI3Ankvp44OZZ7Y7VoBe4bwfQS
WVs/bgFAPd9cvJmK8yDXc3i3LdgnN8Ri6BrYHbktj7DrGSpr+OBmDO05SLD/P0E6
qKfA68j6tHWd/9f1zjLzSqR5EMtlesFDsV5ORQKQpBZKNe9Z0fHJguprzy1UxLBF
QFJu1fCxc67CKiJ//Bpc3TMmJigl1FYsSDHi2I4ywgKQm4Be/BVImWJ3w0wYKDca
0f1CbsHw6TPglZQ4Xi3S5/ZmLvbfyDL2zgYe1lnN6MZDPUDuWaVZjyDnRHZairLH
6bCy/Eu6Ly+ea0g8ZyvSTgrquAXC/PrIJhE1Evg/QkT2MnI+dvhlQ4KtAN+zkTue
q8wk5bAQpSfdbYXzEQbWl+wSk1gDgmUbA+nSk17yltSs9XBJwfqPNpWbjlzp93rf
q4U8xOvj/Yi/d/haOLt6PqKfKgi8jGa0WMO2Twj6X1IuZlCDgBvrgBmgJNc5ojpF
GEG1AZLknIpT5lUO/8NdocnnV8lvqUxVLCoP8/snd7j4Tzk0eB7vhwcWYqRoBnyN
1t+xTgzB6MLjX6mryK05kPaeQEP3d0dRbllPjwbeZuq+3ewI8Pgfmf2szny2PHK2
FzIErj0iDFZf1IOsiHKek7+3wXTpdeozj9JWX+nTRXSgI5H4pZxK0GfilnBAiQoU
ISxI7yX9LqhUComqtmvBQfoEuNKvB5S1QM3jd/SCKdMKT1HYqKA25a3yxyUrn/F9
PuYPQOUQk0QIiLp29adQ5J8XCSFc7CYMDBk+zXOgeggP/Iasdyw5zGSg10ZvMpBV
MJheedC5coefXsdZeBv+ndG2PqSaTk/jkCqGRwpyFuRXf+ZQ5MTpHGYOb2SEh/xq
GIlq+DD0mWTmlDJs3FJIvffEjP9u52K7s2nMhJ4QVr9wsSveUvEneH8dgZ2NSnSl
ODz+VTT0TynEO9lJ8HV1HfmUZV9pRA4DRNAR6qZpjULOOTm8fJFSVDNPh8V9rGXk
U+ie6waWPVCMSEnxJelIWOMFZGi54hFJGWiPgxhdyZMKiztkSq3HAS3YZpc/rzPK
/tDwzcbw7KDzyLZa+/eJIRV7uM06QF0jeNEGn6uclhP7EBWPzIFonrRheGsSVOYa
YbScZj3ORypoL6h1OtcyJHaFWxVfuFgc3+TbNQ87dAm8YosEULat6MmaU9cXZLg4
HaLW9ts1NdSIL7RYte/lwXRDqB8n2PzGPdC0Z8UygiIZDovVIy3hCAufIVfYWwkg
APAf4wfVbfMpsLqwThf9BEJnpB5TC8GmZo7Tl197I8QqyLukbUU4u0xMVcW9nEyV
aZ/TvDG3Ha+mF7APSdlx1mAMsAhycP1I/+FHiPFdkI0+foPid4tFAzOYjZGjUcJx
faJMmdIXm6WUm1SdWIAOdvt5PAqmv/fgtuAbrWfsOOGIq7flG2rR5VN5A9UUzbrU
BrMBk0Sm+jvKiMoyKkn66RklxHGux721JIA6YDJgtvZYCD0Vs1+KM7e15/oywP9v
JdbDlvrpN5vB47VZeWDdhDjORiSVzbmGEUVhfz6poVe4++1bLi/mN7ac2X6J8mtS
6sCpu8uXIe+j47gegTBauz2INW+/pEyp/4yaMbZ62fuzJjVdeFmo8zhunQmThntv
FpMvKfXN9MVyp5Q+naaXIipj+tSWg+pbuQi6W+A+z53eTNvh7dA47w1z0np2RFv3
AsKcJgTjn25Uv+5cWi2Xleyzy3AQv0URovBP+KyvwXw2Ytfp2WY8mIaenvEAqFxY
h8TPHRZTPuBbrlWcdEZ55HDssVeeM2ENJhVwplazTKwVfiSna49zTivt4mkyj7Xh
o7fe5pOvn1kEDHTXeT05S/BxJJFw8U/Lbx0yi5AoeiHf58Dn0YNOiwvll4VrSDWC
26kSb/Giq5zkmwP2QyT5rpHvZf8y0DfgJgznhiuAYE5xr4rbHpESPGJeD1yO2XWQ
bp3/Qci+OLmouMRW5j3SS168+Anigfyhkg4TYvDAkc0JOk/FFPDePqr2SZ8ZL21T
iOQ1RA4h5EbmbP4j4YMvkeXlfQUn7gqsqKJf/JK3F5Bcou/Ndb3vAu6nNUfVFu+N
uvWo8VktuQ/jtXReJzUkCiqi+exZteW82fw3nX7XzVXaNIOQjl281InPn/OudPGb
eHEjlywdx8/RlvDuBwzQpN24ZbIFkzoUoR8I4ygG/h5HzIIecWLOQ7h5fIhS7RZ6
MRgbI2LPuoMRvGVR0J9FcqUaevRK0K6G4wrmosIGckXUBVm63cZktftJgzZqRoDL
CqtmwWsTZMWaQkW4sMo8LqK0SjEUA5M8V0pOF9XgqAAixtNcKrVVIFNKZoCFTtq6
7AcHHhBDqotVOjwFC0P4x6Iw3hvh+6bScFwXAo8//yXmXfQkiI5K3Fh4kCEcIh9q
8nB8TYlu0HEjtoCUPLIjmIQkBDbf35p8Ty2MpNtcJpAcLjrX/qfdG2O8jIn05bIU
66d7Pwtv8XU80UphapHUi6cuYiyWpOlnYvkgN55hoKRLuD4zgXkbat9hsXLo5rua
5EhYkTNWLK2R9pNvdb/QtoSevh5ASC4D2EuO3FPYRlG5Rs7Wu23yKwIy0l3Cl5yV
t4zEuCG57pDlaFY8Y+MxG4mB++k1jvkaqfpMIQpPe2B+12eClXzqneJOc/TbK0o8
nzcXNNfdokEWHmxHTKwQJMTRVL/WkpHIs7VpAqWpEQTyDbskWQKkc3HR7e+zJFYi
XI3BA/yFI1BAif8wkI66eDh3GF7r/41wB7PcHyW3dmPMD0GCWOV5a7OJzEfALCg+
StIZLwJzfEYpcwnfO6CoTYJVLkUEVBbv2HXHOuL5g81079OCes2pAZUSY/7DWrTJ
GrG2AfNEDARHiCogQewjLF5+hRhr3HZQHOfG+cypytVGAQJxFg4qYT/ZhoMhPgZ+
22hXG3RFHL8u4Ot7W6Tkitip92/o5sWXYJlplMB8fi4UvVvl8ISWABBXnHxEhCuT
UMxNh3GDuW63hin9A6b3bsp+J76f7rIk7vzN/cbMYWM+NwO5z3654YU0kekDV2VD
eaoixnpJ7kaoOqFDcoUm7ODR9Xij10zJMF6Wwkgget71mqEknXODD9C8B0NVNa7O
5uGUyUvuRBOWsd3iH6ePY7Aw6kgP91pbnQSb2APMQIR13KgZZaEerJ5dKLPP0F5b
UXVAKqIhjnJ+qRoua5CGiGjpd7SK3Ie8mHmjulvEoUW6Q8X7PdEUUoAKXIM7tvhf
K/dBEWSP6q+c3S5XQFB1vARJvr3LDLeMC4bREpcCLK+nrIuiOdiEk6Yuszv8HrER
j+Inr/MTBpKyLA5eoP4LTBDpaw2TVxGs2pFQSSkdWm32qvlyjLaFMkT4t0CBAXnT
Qhto66MIV9LDQVXrQQYdL+5GhblzvhMCYjdendPsut0qB9CqURt6dIM4i12w43Hp
njaFK7rd5PDDLRblB0XeG7pxeXRNp/Lyns7n7y/m7lQlOQRIExDM/Q4I9FwIQ2sx
63RGNdmp6HEBPnj5saLu07YbQK+rTJXkDDVci5DVH8BLr0/YdBzZMjrzZxNytLo+
N6v+sxStcqKun/KwodEhjWmZGgWk6AVIaA7j7r1JUQwBxc3wJaZfA9ArNrdnsW4Y
a0E53df5L9eNAWHVt36zA8W6a0m67NsomWZv+8O2dvg2Iua+xM6mb3BKvcdTygVc
9v3QyHOpQYhxx/crer+iYchlayJ5n9Ast0M+wQayeBhs9PRwzjTQE6b/qZ9u/v6n
AO52oSXCCGHa4YrY3FrjCxVpzi7f1bH5OKjDImD+1rB7j58zzm3onh2IkG09FssU
A+MbWobpLbxUK3SMSJsu3dpHbHuAqA17CWvI6jB4H+m140n7uP/j+6zA0TddUdzC
DoyCU5iiuV5qQOkZBnEd9kpFh/bhQZvqMvUN7mUekwMkpdFQlLZcY76sNlwQu2I8
yocddjGYE5j60kV7snBL1isjNEINT/2HSSd9BpAAL6mYq8tujNSzAwIry6CJwG+5
F4KYTl1pS0xmTJT+d2s0FzxWIYmS+1xmbASDRiB4gmuB4AUo25BrYQgXu94gI8Ml
g+XyMsUBwvqCIm7PjC49nTlHokFJjw4usNZ+Wv+Q+i28DJFNQj18zZ7DW2GgegVM
bS3auVFeJ2/KUTngLlu+UYnx4Ln0ykBKpxPjInWkl4LY7BUhrCaGUR3UbNEO6hA2
NNKkx3gnqVz9dCL5FvGdpmYIvSiVdKIOCnG6i+VJUtK++URCjd0fCTw4G3P2+SvJ
FIyFFly9gvXwYDAbP7Uj/LdbgsjVlMd1vUkxewP708yHg3ZfH8OuYGEAMzr7nYye
NVWxgKd3Q/IdtreCxs6VhqF3B3pRTgwPgJUy9J+lH4p1kJ3pmB0BCnyr84Fu6TrD
qeyHjZrLRaxzE9OABa+ksCgOB9x6YkZS6yhJo5Hza4+ucmCX0at3qGWcrR3vtUDt
C+wzv0yVIJV0bWQX+fO7tL2trVpU5hgir5bIvqg2gGD5j/LHET6szVvyHFenmVkU
Xt5N7tEiqACBA32U92RixXrNFiKgKLg2sBscMuEAf818Qk8uPjRhbES0/Y6whWK0
RtHX+ZhvfchaKq8gNoVVTFLXRx2lD7k73W48qQUEQo6D14GEVSNzxbaJuIPd6AkS
sRFz/ivIHk1KoZnSUnF/jNsiOBZb/SRB2gkv6RncxoY3p7xbYm8XpvfzKh/GTvuK
WAeJO44lYS9oQdVtj5j/v92JpIQBXIYKKmDbwzdMJGB+dbZEi9r3VNAiuux2a+dR
WWkeJa7Ea1SOsnkDG/e9zdShximiJI3MtkkZre74rbczXcb2li/23kYM2IbrNnDg
dQMNH3/q9S/tuZLFTTsT/a5YYMKWNtMt/coDwNsywfB3xl+ceVQlZID1uOIWq+Qc
8BWL8vKifcb6uGoN3jZmsYF1wSYPNhONFRMHlbOE265ozU9Me+4Vi+c7HBggwCrV
Jr5NSuqUVIu2idpGzWa+HCWnESAz1wW/H7mkMj6r29RHAYHWwBmtjxwREjYzvqhI
yfXnxbXVueRX3r7AZsy1fD5/sXn1drhrKiGgOle6jeNZaEGb2+8DG8hnQWbpIRCk
O+hs+zViJ8qlzvxkDwc2cC5uDi2FY+X4Fd5LhN0xzOxmW9WO/7dUtGmwzx2pZ2uB
nf9SGs5TnJjyIKCKv44VFG2a4LtbUdhwRVfpKwdeEK2je1MxKedU3TfuoKvPgioa
/sUQ/jNpBMYRmur/1W/dWcTsrqemsaFSH1xqAB2feP6o4ktFq9DStikQD29ksGpY
hS8NBofclK5w7CR9ZgjSzxNAzGlENPHyr9VH88IEF849p97p2J5W39PV14dp0q03
/Klk/jlDhMp30Pq98eAXBpAGFcB/5igsVz9FjCYZaptXEGAbKPgqeWfMHkCZTB7U
TIf16Q+LfcsfpVbGkFv9l3R0k6DvojzuGtp+HhkA4Lmz6muchuUFHIarmbsb+xWy
Pk5xfhOsTxCbTGIRjFpozR1mzgEocF97hJUIfQpmy4pP7bbe0UxtAU5s6G0Wj2RE
pT/OVawJG3Xannx5GvcBBoV3Hk5C6WQchlt04xCYmDYsTl6VTF1jRte1wL3P7ofi
xi2kX2vyhfl2YESROn2q6LWjTxOcYiW3rJIiENFY2Ue6dqbSqQJX8+BBaquMj8bA
V4hkTpGp4LAzBBr7VIBEUHvI9K/Xw+cDVkKBuIvKXYP7ZyI9f9Z+821ep1QjaTtZ
w0OkA1YbBcrxHA1JVeT90xepO9nBtQBC4W9F1kesmcESmJgLPXuCCwdfg3rb8hM9
CKs/qxWJylUlLb4d9hcupqWDHbhm9wqQcjiLlTL6To1npwvAp6Z9ABCPTTCClg+b
2HRDyQtSHrhHu3S2dl2VmMBttKwWTVs6OF2I7JUKsfZMLsPgwj3rmpaVr8Vcavu+
hmGV/2Cj12VRSvhNsiPGsO0uGURFQ7Y9f3zc7HLp13hnqUFIpTaMM/VNQDHIq0Ed
p5jplSQX8h22RgQQHATMB3+//IN9S01vmJ6gneWHE9rzswijq6iP171OejxYK7Bv
7hmxQsNFwA+mq/NuRISHzcgVzw3PHwBhiZ1UEZQqWDN1n2O+er+v1f7W9Z8CWT90
Ogfbn8N0/DTJV2FB2NO9bQMS96+qG3zoqs4UDb8hxGX8vAj5wgo0YlgQFlZ+rQo2
Z79aH7KnVT+3D8NZbmIQ0XDUB4orFcr+neqUv9Y76up8roGvksdJX3MVu/3EKqi1
gJZRT0h19a0uVJWE9guRUuzF0VXI6to/IuYbX0j03PODg3PJnG/AGLim//UEKCzg
LRyiJOGXmbVrFntN1OiriWhuS8ZrAZgq7TRF/21JRzS/k/Q1AD3Aeow+tWKb/izX
lEIjPuxNkXRe+a+r8NKfuOwArw2eN+mMdWeb8MD1tSNkDaMPDfAeauHq5sjCzmB2
jlfP+ciA+lf5EwBI4ibrtDA+F4t2BOQPtydITgmjyLQEMUIvjcDWaKYy39GKBVrg
QwNJSFQtbAHujneBZU/RTWnLnG9wNP/s4o6UnTS8WUYJFdvx0WRIlqKHSoSksPuE
rOtRWEi6gVNgwDCKD58erHky8fuL9xqlCykfcdmS8Qx8Sdf1rbdko7WyNxDfwh0q
KQUj2lcclzyUcRrJgYQMK1p6RUxAJhh7fwmlj4c8Myy6kVg3nVW1uajH/efb8Pil
cmsUFgJFYmxKiaFE9IkdAs+LtxPmP6cVh9hQaaheHhCCKfT71wbVPCIHw9DXHG2V
Pukg7/kFXh5AnOqAND9qicOBJ9/KI23AknrlygKHSkehSoW8XEgGljmYVBKErpKQ
G0rQfty/Bf0gQBfxFBhnPiLkKxypTCVufkEm+8vfgnZTDZaZv9xG110achfU4MTF
loN3D5CM+wZ64IXKjOQ5L3W2LjTaywlni523jvjtWU2O7JzPxYztGtoPJ2Ul0pTm
zayek5Tv4J1rtQ5zYnnvGB4ykVwo+JQhNc7/RoET0sYe0kTVtpC1K508Nfv8oIs9
LhD6iTN/SsksFPZIK+Rz2EDvzzGgemYWHjK0KT9XQPU6S2MXUNYF58xs11GYXg8U
njnHQeUMKQ75d5e6Vq98AdrUhN0cTLpZzp9lZeY7rz06E3uc573hdND/i/Ih/XU0
QHOsYa8BCEZZg/boxxe1t94oFlSJV7Z7TV697GX0ZOncIedD3ulI2632rLtxq+Y/
VtkuCRD9Jkm82RtYSgtVY2J3dQCkeOKVuWtKFjxJcsfJdBF2Pntea6BLywuymyNO
vWjCyXXZwwxZZnVnHb5Il1sJ2xJLdhvKzHehzSbMJ97TgpD/rx/0qhpfLYRZMMBq
8CZF25tiT6WsGszSjapg0ndtNeg2XaWxIKIF9PhOCeIGtiNEuuEkNGzMqxewST8U
gY3zViOSdQ+DsClEGvpxTv0OJPL4Eza9b6IhOn6Ypb2PF3JxPjvm47fLLnmwHipW
BMYPTgDGA+KN5YoA4Np0YJ98Fyzw0Io753d47bccaKfMlWpJcw0HODAuHBDMEIhE
YyJBPpr5g7Tsxlly3JeOYoWRngOaa/EELbw3OKhf6uIZ135AgtAQ7scUPaK6t5Yo
o5sLOEv4zpnDi+I55K3D0RJnbEDrsGXCxvJ9s6njY/+kTr7kP6D0NZ6hP3QIYfIo
p4R7gIdh6uFnqVtCiUZ4MPLUGF1QU1PliNffppbBRc8LNLAvUzbUJ7pTlKH/RM67
ArGQCNFCymOXomvDxmjNHxwXpCY31lOUNNj7rjX1zgaJ/Ed5ODUsywEftDrMxVuZ
+zbqZYMbH+OixMiDbUnsmYY07sS0Eg8tng8KphP0ypGPniqyi3ln+asmkkRZrcD/
WNbztjNm8ByFcIGrHnAQd23gMfbsYs1zHY1kOu9XdQaH7J8OBEomE2QOBTwJOvai
XIeY1CQL/heb+h5Mayh9MJ8QxN9ZQwqN6jDvvyXYHLp1wrtFLFjod4gzjrfiaEut
mlwDg/8Xy4S12KR1JCtVQ+DlK5O3JbcNgzToGoTFjpUCuAvf1bYkdE6YwlJw5bZ9
hRSVuSkKuMM3RjYVu9b1CUdHaPRh3CWWuEp6XCuSb1RPczoJcVk9bhAI6rBVsNHU
yXbEQajqSjYI5CCMtW5/Zx2EW/YoZdktI9z3E1qmMq/9j93P70VzS/e8TS7AG98X
XwJQStGBbZGcYMSbSbFhZ0iLUjG23arS0JaLP4R1Qs+jCdAAruNvmqMUx9KgWtcl
u4AMrcy9j0+kJcdG1YtEVovSbX1J1KhIg5DZLIPSQswiQChffZt7IJVR0afE4yyz
xfYGikf1eOEjV5hdhP/jS0x9+MHGS1/WxyMETkSx2Qs36lhfyNrXd/gdN8JTVvdE
Oq8ov6GBZ7SIcZZpEL4b586FeKK4TzlASV+4gwM868LYTJvKUsufuSQp+215nwJi
N/javXQgdiRmyGObB+7qPZ5nseX5K5YvdJxLmOsmaJZKTiBFlVMWev80/ysvQpp5
JvfUckw2youPRReN7r7YdfbRaypvxFqvHWy8vK6VObmTQvuRG/gGfQynrGRgEhhR
OKgtG6zCuyy5wnwfYx47xCRcryE3AhSWg8wJOQD9xvBZdwu3iDLbeakPnkhHNMCU
VtTW7zkMYmsrIhXt5qPxUfMMMhAYp2+3aPx+wk2iyQ350uVDbOeHEtIbhhRKd1y0
KC0Mom00GEDVroIL34r1u9QEa1jLxoNh/jYlfihhM0/wLIkUMWAIrQUwGJizRd0E
mWDuNr4nvhE/ldPVizqvw/riH15iB2y4gFV8SvZf3ekTsbZ/BsUt97GN5bKQ4qIS
vv0dOo1chSyHzgH/SgR2EmWuQrw1c8LBlSQ0QApknIoTt3kRS0gM2R3ievbIvaZw
xqBEQGxABZjvfuMsWvqHqTCFokxUDd/pEBmSMeAlKZP+IvthLjTPQWJ0GHOQ9l+x
oCuY/XLC59JbVrgODenkWfF63Or76yKxt4fPeOUaCHpMD26JP/YIKbJeOJ5U5EZq
uMlYvUyAG/DfZaXQnAg86H4chQiFEhprnQM3jN/Hen+83m1tsRrFVyNTbFkgJJru
qZBEvHjcfS89wJv8nBwm319IrIsTc5r7kyx8WwUlebmcDTDuMLDR6HJALIVusibe
VaDMoI0EThcaBZMA3PY1LbbKwUHHfNfvxVc2V4/A2kN+cRrOBIUzXD5mJGx1HGFX
YIdnZlirxrOKfhxgd5IoWGIYG2al3joNsIVIw3ET0zZ11MAMDWH6a6PbTZM2J/7k
bMTpRohKrVlMSAzvpxGvNJYkmID7DUFpvfOwxoQLFq6Wk337bDUd7vtx0xHwzIHx
4cjeA797Sdfw/UlMYfLUFXGJ4171BjCPZTXt7y+17ZhzeMZsatE5AYSN+H3hHfy7
+w/DGp/VfyczaBoTAAYrXy+q6MzLTYeF0/PTf+6KtplCFHT6VgDDfkMvEMd2xxqq
WRRE9/LluhTyAOwM1q2NhPU+RUyZwnrtn64rsPuu4tGYMWNfsPlpARbZrs1InAKE
H+V2XgEqhnUHY7vWFbrkkTC3Ll3EqorCgyBe7enhkBnZ2UJSCKHeqHD4erkaN+6R
ImEdDG7pQUs+AXGvih39P95Hocu4lPTRkfv1f3kYg/F+o4O2SQ0a0MjEgzUtZtD6
RC427HrJ/578y3FlIVArYbzsxaz4XHNG7wnLuzdqU0R1x7PQ74aRvMLD6CGomvKM
JMNmGsTS1dqM9KjY1hJZhCdQzYtRd3ryPCXlAd4mdx3XWst4JEOHD8XArgcUHpEt
IxAGRdk5YqDlrBz8Bwehk6djH1p6ub5sPKa+wTcVLWphhzVxnixKTvDM8ibYqH7f
8e77qA0djB8zDFM0Dyv4XijwhE097lQZ6yATS0FJ6ZaHc/J6u9iRIyUYU47rpd0i
77j2ukIQxZrcLX6/CcQcYgFmGfXn5sVP4LPz5PaHYMUe6yxt2KGse1JVeHhsnWx8
ywEYiA3scPbGuo1aVNlUGm9AITteFcclSRfS29MK1GmXW/ENIc9a41BtCQayxea0
bLHSXkQAPGqbaFkmaMKx7JWe3m+QGGZQzpdZQRFMMmy44n/3pttkUTfiEsS7qYoG
lkyjBeIeD7LF+nrrT0rgNNsFHttFduQPaqZ0n6YZePYxyJ1F3x3gfcvWsGaxrU4A
msio+jOYgmOGQQF4tKEnx4c5QfKsIFJ14W2T4GtIQgv5oqttppn+A2pJm9DyWr53
GrPAXm9HJxk7us51AVcTTZPKk9q/KGUiogtxUVjQnqWo0eFq1QmK6ermAn4Uvxiq
BieZryNY7lDNUTdN9LMz36isPOnjhqG60Rc5TydzfckA0RsJCPhv5J/dsrKylMh4
49udawW4EglAmJtoCmfktrgsNYudeB9NEo1tEbdavwy9T1Qldsmv75nr4NB+zLpC
ud4J87zv1kzF6RxFZAroLegJsXY2QNwFRqa48M2TWiD+NdWxMNFdFSY/hfcL2tqy
dxc6Pl5NQHrXdrC4/hdlHoPm0yqLraOshWiesBzudd9ncozMZadtTlzfcF8LMFjk
lokb55YHK7s3YKoIUz6VuiTjM0oepO62D5NUq+LeDccDxXOsG2WPAHEfAYEgqBGc
F2FrHJg1TG3pHrDDL1SoqEzoJxVgkNLZZ8ALgObNV61NHOGf4KckTvcv1h4H3LkC
ZjMc6vKI7TSzdE7IXgaHRcsfsQvCa1x1fjvbVybTvUOF5GkD3/FCv0A2OBqfKD3U
RYYF+oqKuZmJFjlVcOnWZyj0/mwT2B51Xhj9RSfvC90XYJsf2RqShyNk43EebABV
MRxUDL9ldQ8zhe3xAfpuX/8uoJ8/wovHXC3OvPfCbySIgCSlyjGs8OZ4z8ci9LUb
HWwd1hG2WUGEDkfYWTrWrIwq0p4Mf0zokrw9SWW7lSpwZD7ex7BGBDeOHbyYBuyJ
VL07Ns2Fpae4I5OpghehUdJb2AqSqNYPdrmyz2QCJZiBUoG9i2j8RtkSyAp440ub
4JON8a9aUD7dnjfDMzTT3y4vpmqbtSjGeOO7TeXgdVhhYpNQrMbbpwpFBb9+MNp5
iQELrif2fcxmlmOPjs1zoPigKidPc3cxm5uak1if7gYmy8Bv6DxaX037UmIYVoiT
qOgrrgsgePItjoan/Lf2EtCYNl+Lk/4PjaroO5UvV7GpFt/BE87XpUsFyMNtyeiL
074QirNzzcWI4oqI9TE2tycXcGbDO9yp7bFo+bXgfmop/y/4SbkL7nS9DBM4fOGY
QGbQ5XxGtKHRa2+jWXY0VuAorpiimCNecbjuaCDp1Kxq6dIMZEqoJVtyLpnvBqA2
6Nn+mztKmrc6xkFe6OmXvwRUsh8k9zF7SHXY5YwnE0q+wxKT5Bhflf9kNRjP2YPJ
+pAmEDlEc663jvaEud5AYPNLZU9ckO6dc0NeoBAbuGXE6R1n/Q9OM280iVMKUOr+
NTECHpLo1CB5fT/20dBkSQBikbHWFydli0qWtaJTS92zyWtslUisX7MnNzBM42oL
Y+iEfSJ8I6Ala0LPA+ytsSAuJDvP61zUkZD8D9EkbpIuJqQh9NucL87Q8pZeM3AD
lHEjSiJsxAQSGTeP5sVOSKIk/JFW1xT2OXyrvzkGAqE4uPHxBuGqzo9eg9Vi5VM7
wiBwhFD6aMcIWh8Rh5q1Uk6u4/pmq94hIycoadh/+32liE/EmxGho0DNnldz4MNO
YZKt1X2b/0ebDHp5r7NxygeUGDI9Bayqchg9tfBdoUWHoTFpAs//VHYcDTmXuD6S
ybviNGC1oIbJBykCumYdITyu83esIYKD9aKKTEaTeqS0YkZg72gWG3jet8sdGHos
ZOSYJl1G29ndzcPVev4ir7noCInhRbKo/BaWbGO3SnT8CYyVq6BPBOxjGpLXRQT4
MbCYjYzLmAYl24djwBO/qNlpHO2ZSgZ1V1M9zyejZ1JdnuoVgSrrMhRiKIO2GjV6
1R/azR7dJWO1dT7prDgKkJ+LdSOVdjOgjIkoCEvjWZZ2FcZpD1GjbrvSJAUXUE2Y
w+XINt3VCjqx1lNgr/a5tUT8nPq8vez6U65i6OlbgQwS8SHUWnEgNmMSnM9XfKBl
sUXTjgalV8k8Ze2bgEgie3wLA3RJCLQ3R96WT8EhUHK9u51zlPtyFFPP5Etu3juS
xdyPzVUtuaKfnFQ5OGjFXvlhO5M+z3rOQ5bOJFdtLR6gHrm90OBtkoyW78rJ4eN4
1biZfwW8rkuna1ZXJ9FuGZa9QRMrbgwHjIpxYVDoB/Ekl77fHwcPDM9scyEalIDw
gEWz7Km5+kUnhpIFG5Hft8oO8ZqOVIQxSiEt6/Cn1zAJJzfOeUCJyE7ZXf5sDt6N
1Er1H7fUA5jafxm+99VRLHFljb2ViVBV1GtXK3mzRtkk9z2FV1xKJjw69VllEIx7
4dmQIPBYhbGBzWs/r1Bw7Pm+R7j4iUmhLWQprilokMIQldMIZfgJ8SnXG4LYCv4z
CRo2ZSCDKyyiNfItV7FyvrmIVhGflodt+px2lCwY3554DrrA5052I1iyC9jv6myb
SqKGqiq1uiZ9d2Q7h2/FwEpF72K3Oo4YQty3DrRJJsWwrRG4WM6veDyG5h31u0Dl
k76s6tN2w2sPF0ZdMqjNF3NQwBQ0ljZAUKLZo72ZHw88EMqElMZIYtAUQajqgpl+
4wmDYafP2Hm5ICYhjytrQO1U7zvccjcVWNWH7duZGEXxdX9kvDL9rKLutk/L6aat
3lOeLxjPCpdZu2wJuO9oF/GpGvyJre0D3d/eIZYe6HUDUeHAA4o4WR8zwf+mAfHL
B9Tu/Lb6FjX/jTo6blbakgGrrwFdkWHHaC+PqvMfB5MNj+1X6FL/v/+EJ5P+eOKg
cHiHrfasj7NTKC5SQcTueh+jqLxwzAiO1GJ+bTP4k1YJS3aRf6COoj+l0nvZz3Tl
qO1zvaoqXmMcjcOIq5c86V7swtDmsh+a6gc8bAGrYP4H9rNWGV70XqncRHZhr3bV
sLpdwU2GGU7IBkKlKB1szyPu0QBqZ4bV7jrWMyXZQ881FT0xmN0+Y5WoFNloTje+
bc8LaKL5yJ1JPzLDQmspbFT+hFO6aWvYFPWEhTiQaDA9DIsSJ/wwpVZeR1BAd7/h
3OqSmvMIeSMT7SA1yFFHZrIW6QmbIHQiCpbTtfVRibqM3xERhEFOH2zwJaYhvhUE
EIFVQTWDmz32xGnXb8eMf3NYuqqQJgYERcdcse7AHfs3jFX8hhexhOFN7GMyG9w/
gmdPgkyCzluWxRsY6C1541vtpOuUKBJBKNKNCi4YNCEkSHhxjoMxtDtqhfSMi0QU
U0u9JtPXwPkpgpMtg9dN9mHt9WynBGXSQlDXdsa30Y4C2gx1ZwLAxY2/f5FeBlXl
4fJSXkSDMTYmU1Qf7JB6DI7QyGdYbdPXZrF7tE0tEb3WW7KAA1hT7oJmzeF3lsxD
RyjgASaNazN1TMplLDK7J++qxBSl8mAuvLeAp7UC6cqm5no0WZyqhb7tJiSgC3gY
44gIe1TXAeUyNBP7/Umm0t5KpqnMM8caoUBHDQPh7P8jeVfzUtpoTgKanddtfK6V
wTuyGtUDIYH0RQ9C+W7TLQnJ5KKRbrA52I/hT7jN9iFgCiXTEjNZceoF/IrySjct
btNAgo19KOOZm8pkF6vCT1gCRByig5KInQx+trpUcmuy3i63ponu30hq/smE88xb
QbsmnuSyLpuqvEZeRsWE3Cne27MimciJBVYaOX4vpCM5FVQROGdl2SkAHn/h40IL
s5S0C1fPCrW9qGqdcctnOlzP+cOc66kzAUCZaEVGsxBJ3ztY8SsZFXXMa0180xT3
z5HGJciUPXjB2BvlVjCaNB5rle1/+wH/z1IVRKP1ZdnneWwsxRXzMm/TgaSrVVCg
zY1x0ssldKk8zu8RZTqBSg5sMUxDUE/o3ZPAwJs01uJaRG9g70g7ek49V2sdtPQl
w88z2EGz6bPJsxLaBpqwSV39Q2OTi8tI+h2sl5FmyHfN3tVNx6UJC76xWuw2fvaI
kDKTfV/VKytHcEiCxeYVttF+/Apfhpl6eCg2tn6auaNr2ODjm9iGcF7nzCU1L+Ma
5rZPu0b9aro4LOQYzjBjLznqhU8a4rFip3pn0m4HXAbaAZstpaFEkiWefBVUNF4F
BXz2lX74X1M6Yvm0PunVioRbWr7pluEHp7PlqjYsJanis1Q1YPaVumJJP+IlW88O
9ythRr/oJyL0tyc7DWpSnpqlHpQ77mCJo/wkrDL+SR4T2Z0x+uIuhiG5JWHK0TtJ
YdR/THMVsRgPaxtGAe04y2JlDVUw+MxLmJJHCn78Qs+CvjVCpxtfsdyA94QuHa8O
bUxjTkGzANaUx2+yMZCpCtFRZTL5L4m4CVELDgjROFx6Y2IxmBN1jA5xmhE713Dr
6UEueGbp3vC9uZPnamN1lDrtrrmD79ubyghqvzrNCD/0SkDwhLSEwQvRGlpk5DFm
cH2TNNGAiIJsxWOaooRCLNGwwqGeNVSSN0zew4jTxeUcWVpmz7qY1lYt4dgfp5//
XTTJ3YbuShHhauNrNRNl5cFokzlYyNDki7FNKm2BwEV8xoKoYr0nHnRLeL9wNtud
chZoryWeSfB9cLkH0zNRDXlP7SI9LM6BjhS0mFlEB7U1o4rXRlbOfXsX9Lpqmsdx
5YaMp5C4L1MjwPnQZig8K/It2ksHyj0a3LwzGy05oS/a3/KTM8L9lgMp+AP2ccWy
8WoZOCv6d2NXdGiJ2CS0SuEdKRPKLyvk3gwDCxCdFGDzytL77pQKf1D+xSAtElTq
74SdlAQOSS3/+ddJTC6R+OzrFXQuoE/bEP4rdw3v+O2D/7aLSLIUXvguXIThhoJ1
JL0JTgJ748U1O2xP+vIO2yK0Lah2+gFZogxpkJWDWK7uH6IvANcQiWEzpjASrefy
lRq6/AXBEyBCpzFjnWr4X+JuH+/XICccF3wlRhnseG6hVZ6Yb2no2MTAhwvpmeQh
JnO/z0ijgaz4GyJucRralvLwHd/hv8peKtR14LsGdIYq8NQmV+Ycy5+FUGw4AO/q
m4tpRevDpmXpKZTEm17iQjDOarFsdcKpGPs804FTObn9Y5RU+Kc9BKXdbaKLL29S
p2r8O44RUYYcln6X24aKomUXi8hdqEvRgLoSrB8JUZhRU9zYRChWs7QAc9JilXSI
miHat/l90AIiDah2RWUfT0LEmxfj6L8mD+YDx8rP+CA6oAIodaOoZHqKpUzS3UIC
9RQKt7SxYgcoZjuDZRnJZlRT/ySRbQZA2Jp5r9zMVqB+6w4HXJCZ1s1kmw6HRPJG
ssRJFcXc2uQ04BLg0ySiKI7Xw15HzilNmHm/a1Y2uvqJOsnmh0UKcSpJzyI92s9m
8jjkS94ESMuZn8Ct7znZ2MnzCGJ3dEdpO2OyLLgbrGu8qWkCOoLe7B80vtVDQ16n
Q+fGnXs+tMaPYgRaaW4KofNO26HZhyXQl1lHnvo9sIoMA2ipD03Nb7ciovG9yYhn
5Hq2SUIbx2KwBkZ+7krrxZ+D8knsl3QhZ1NKG7WUlcBQR5QMcnr1kmo9fBieZxlx
FkVMIH4zK6QoA8ndx0dQTnGE+S5KqCop4w4wRDQyAV4Ksf+Di+Mba4fLqgKa4moh
IluHNfk83kh8otkw8p6S0MsjVyIEHa0KfUSNAerichnx5ZDxXQ5PFyJCwzypf22z
OWGHqcnXYhdR2jDqzGD8Aylx6VAJBWPMpnYaD6wdAOy5H81MSr4SSXdsh+wJq7Gk
SNpRrJi3j66QOIPP13NsEETawdO5eR6qrN8wmNs49vWgYARaEZ+i7T60wQ98dWao
pNbmeQH/DHjeKJk+hHcMKkOfFaxgTzopZ36mOmR55hVHzMPas3HkcxvAEDtBGiDn
InUpZiECXV94ntvInPNHL2Uu8B7qZmszMiMr9GGj/j5Yz3n3Ae86jMXHAGAKKNYu
+RJOgOT4bVK4GnKtGx5gCoGuCHxr5JQC7yVKfyL4CosrnIcpAtVrBhiMc7Pxx+hc
VwzNsCXBW3bJIepvUWsEnj/z3wuk0qBBGOysRxq2lA0nzGe0xzsllUUWRI+H+OI2
FYuOdJmwvM5T7aALmM+Cvr9cbxEshfYlPDklcbxuc7wDDQnp3SmBq7fIy8sV4Vvj
v/+5PKumHYxdIuu8HHrg2FOxuECQNX+rIsEF8LCw3dONJWxHzaw8MrqxdByytA3k
vJ7ey39b2TtKtWd9is7jAzlwcSkgNtDSYDr330SfHE8S2SV7Hvmzvy3Jvz4CbBj9
aaGMwmhWwdKMRA7lk2S6Tji7nXI0wrSbkuUp5StuJUBkVUavpS25Jp5otrSidZQn
qU1NFVY13Q/mNCrtX//YP0KKZVNJmyGMBCEqJrVXTetYvQucWMaf4UggZgh/jJVj
SmIY6vSNZrsFk1RY7MOE71sOYaxFlqdgaoDfaZHpAvs+hfOVjJqA7nLfTJy18HrA
Jd6X4+kac329tL3FaVQKNLebmqDYkIPxWi0FLwpZ69ERHeKjMXbAC96ekPfC2iYl
ow3yjZa7E+IKzUhgi7J6QEpWetgZYJ5NHmGjwQjhMlweTGkaREUgl/rBuU8Le42f
KUJD/j1IVlPzadb+7MG34LSW5OHmRCSsbQ8U8HvDCHHkoJtPRt6wbV5StC86PXsw
cy6L/NbPNdFBiRGzrUZZM83YkZOHwNEByPaWArJ3B0B1Dp6A/9NMTURJJoXRDEb0
VVR+pm0DwbjiXwuNA2Y5ou0s7IlyPsK7kM9u/LT41PgyVL+V9tyeSTb14Ja0HZQ1
qVZKVzVlMi/6Vl6Gn3Pw+U3fukHEatQOO6t6mH5Gb2wGfbYjPkdf14bYytaUpN+r
r62CRbMcL5T6124OmwyYNonr2qS+FPYsT9a+dByOyO0lIzDw5Ta6ziiKnasm1/z0
tYYn8jNmLsfQF7oICmfeKkVEWAlfxnacrB+NrvzOZiduIXBjxt1PYh+Ms1nifroJ
5rDI/wcqeDxTzAliKBZAOr2bxyJObsJ4OyMq0+ai0vL14qEASQKxgnHc21YNxoV3
WOoHRW0WLRJyYaYFWJ84aUi6TWzcoOS3n1BHUyO2q9ogVi+/2KFnl1VcVtTYLLgX
l4+TcR6zPDmDx6sthGiv1ipeoS6YQCthfVMnYe61pX78MnivPQx3R5PbMd/xbzsR
slbz6BCp70uFZOK/F1kohfs6oYMI01svOmk92mOwarFRQPoDNSudRlGkMomOjeUM
H/Ad6spwtIwWbVUKO9SFhZrutN2OmX3eXzy/NDAC+8p2DsBn2pdNXkRNmKc6rRLF
NayGnMcDyW+LucMoa9KiUABljl0HwvTA277WG5qmohgCUhEM/XYKm/xSaAZKhBn7
gxCaw5xuWa2BAFaFRDbvxO9+8LV12eG/KVaFhUpA4JnhNXAkU0jM9uOFA8NGXmms
Ue8iRly3PhEjcJxk9G5D+NsbD2Oj6KhCdnJUuSNpOioKcbwTH3qqTlJvfA8RmZgD
fxmdBOw/b2XHnAnArqx3yBP92j7b6Di1GRrb90m+ohrC6KVcZkUbgyqG3c06TgT0
tYKr2bSUrITlgE+7EXsWr/qKirUvwdjKBHr0hEwoQf3MqGLgVruQte+ONnTSqMLH
a9jwafC5A25EdFOW1vOF44YApYHxRySI8EpXX7h4RmaiiGwwr6fwGckDUl+cG9nn
g9Qkr0A0kLncl72JrI8B8wEGF3bCrRnzekDlOSz1rOkhoSXcfkey6kHCBUrtnOKQ
BQxXsAN2LgXTdB/dpIDoXVZpliV1ZzQrih5LLEYi35Z5AzcYc6EQljJ2GHVDEQuU
E4GkJdu5NrhkqvnTSSzL9Q/yea79GaEzqtMpzrgyfx9P3FCZWcD3kMBW1jSDZZbk
UtFgoA7WCWdqQB0hCLiQQzTkA7FpVmx4nnLdIBs5xyJfO7PKQkVG8W1doZs42B78
oVkLGBbg/uXSlvNiX/mJfxpCMTiB9Pz/MIvqgV+pancCs5u3h4BuxSvD10UwMKkx
CuqHsw5wipcYY6me74Annuwm1CYSd0Mks350JglkDZc1LpUOBCytpG94oAlU0R7P
wRImUuTV0cpXV4qHWKjaICU+Y2e2nEnkHHaoXOBMUSjUUYNz9+5A9qXFKYnvGJmo
YkxAPQTPWKIjBygDgsdlvCUBerN2fO6JR08HW0R0fLW/cgg6J6jgM/JtOoFMKlR5
58+hryF7hq+oO6uOGXm0KheA7q0rc4ZOno+qcVcWOPVlwm+pOdgn4mpHqE418PBj
sPLHJpolcIcbXLQ9wM6oYqlpCbN2r3PVIsogMSiuI/Z3D4oA/IuDEgROYwdo9eSL
vEZYhzN3LyESOgethPK55qb96tTIgb/DcYF6M0rfeNfI/UweXv/EeX93ZsYYXDI4
oAgPI4jD2qTm3KMJIgzsbfVyGbYzGSf+hR225OsfbjUx4mDGPcN6AqmW0FJwH1c/
n6p/v7s5uGnUzDTKuHyjh+S01+DQRsKxJPcigeD7e7ehOay9qKBKDPjMhDvDZXaD
H67RrIuRvk1INOkvM1Oht9hmSCYzxnypudwYtp6DejDJaDe1k7L1VIhgbh04jJuX
mj3AJ6aiyFvGncitME9BxfSg24L2/qh7AFqyOWs27JgAvnBbMgkuOSMQ4GEQxPNX
da0BiHvUXwvqWDrX95gHxsN7LvUEpSw9QmKYULtEg2JeTxkJ9uxxyM7mecsYnFKk
3As/xzSa6PUky+pQstnj97yS5QSIILvd/f93PKQX0zMW90xJ1l3fKhZ7TgJIDcyF
OWfKMLtwYkZk5iq81gMw6GRC7sxiI1Eu9JjdXZZiWzAnqdwUt19fmptjSmkrT5E9
dt/cydr+jUjAGfcazsl+zqxPCMgXaRp+ee7Q7s+jG7+PoY12wFJTkYxWhWUSDLCf
FA5qq87zvHsCxmsT+i33Fk3EnVNbIJP3YzGd1MyjOqQcZf6JKOSjdfVPiFtLvukv
YQOAWENPX/yX8O3O2Lj6LJEWg10HQJyZRzRBNxbx03cWS0QiExkRblQQb2N1ezo2
NCgCg3Jnhj38NxpqE11SHIPiCAOEgg3JmTpoA0ZhEgzzPdwXS7vJn326JbOv/SAV
VpStWn84uVh7iNiNmguxXxULi+n+jjk1oqeC+5j0QqxFBtU8JbrpoAAByUkFEUFS
Ona/DI93jI5ahkkdWkgR2DheFh/PT9orf+eZY5PZRPfp73lE8BXecNfwjwrdvqUV
qYcEZc0L7Kw1WF0oLPHKxDX2wCUm3WCb1bdRGWyRbMII/jXJLDk8q+COYv8XZhNg
9G5ITudoyw4Pc9ku9v8wnaKBRoj9RC/NK+HWoH7Bg4cOeV1zHnAKRLrAN+rzpJdv
P/3dTAGKSTgHNhYCIJm8BUzUXtCNRjPYzGHZk9LOR5Orjd8vWD437QKFMti7bEnT
FviSX1JGDmpBaPSGxLPH3HPRydKcxxmpPiOZ1x5OnzxEnsPU8pQD7Lawmol3YnW/
7E9H6lU0XhWxFZzbFADkqxmq04yFHFbcjHDpAf7oWKHQFrOpQl6s6xB1PlMLsarQ
NPSPf27hq6+NmPeffgY4sv6Iz8+0gm8SyUNNktNaqA2OugyPVh6uv9eZ9PKD5tUz
8bSqvCGpULIhTHyCcsYQZ8MZ05JVNN4Nf3ZEJ0yXXWMi7e1zhT8G/HfdOv2sbMsY
DcP/V2yWjKHkX/Bm5ulwMiByiZn3msjB4BQhmwoNskF7aWUmQkNlsUUPD+ik4Wiz
9xY1t3GZCfDHQrLt3e7quiZyqpiLSodKvhTi/T8vwwAYRE++HSH8ZZQBUsII3NfS
arTSidpQh047Rcep/jV57tz1hLzDfVx4Rt8eBCsy12iiwQWl2YxqbZEHmt37KMyN
hUP4hGuFEiW/BV3AuG2/XmZcjgqhVr7N5dd++mM8VEY06MLJ8plSq0/Ww+zKXvJr
dRXRLh4qyuEDBGJitu0X9RpfpR7xqeUZiE9pG3ech/LLhejSylDLYxIWw6yNh4ho
4AglmTgOe9Lb0c0zHape3wZhlnedfevV/KXlIvIKlyx+82FNdA6p+eVcexqWiZ6j
nSuILC2jzKhuJcF0SgZyX68bNIi63lG80tPFqjmvFNTwdd7j7V8ZhxvP6S251704
d49n31iAQ0jDmNMcU2hOd+7tKkdXryaTFsBjrQzraKVmxrxLqmXj2YDlROKGaVhm
HWf2xsrHi7aV18+U/pbCjF6BFkhZQt8iF1VyArDxKvGkALx+GpnWStpkU8Oli9Zl
6HdOuzPJ9obUuWTBRiYyYb3gVhmZDXupE78xwGxk5fxuAxroam6Zm2XAOlQRDUou
78BJpSX/Ff7nadnoRnXaqbJJBPkoVJY2B04wpnUIDyJpwguYWfsgTgda+kvf0dUJ
hqdr5xtTsLZ+NuNvVKnIpi35lLLBtZcnsPAMibgZ1mqv3lipIYseISrK74oebSi4
a8+Vs0KFi3bmS0vdTtrHTzjvkDMDDyotDaEhVVLNxnxAMjpfdLsR0ojlSUm9e+Cj
8dDEdUUJEHjStVGSXdSS63kDjS2IwcG1Lcns8k6mkTKQAmNGI+TxLCpk4ABckV9O
jobe/UjIdzYvvRzyHMpGCuOiYh8QCDmMxY/KfA4A2fqD/tOXJvUS0KwdeLjK+HXk
9Lt4r7yfcIqjQ0HCy9tLkLi4ukN75iCNODcn9d89N0kFF7YhAFa1ws5W1Z7lRxNh
f21FkkgShZpQyLTAdRULGcGVOM7qQlKu44fob91t6AU30TeiHm35NCCsv+olFk09
RrvtXDGfcGD63Ri96BJHva9POy4B2pZhzjKMHnvG0J8Iiu85oU2B5B1duskS+Npl
SZixYoJ1k1HvaA6DH5KV++ZxY0EDhrY8EzJmZ6XD1zbQZV0Gzvt6tFOsg3i4xSj0
6oniLXOGU+zoxFgoU6ycMGUMRFeo+yBnrdWNUxuTAvhf7vp9OAHBORG4DQachzsG
0+2W0rmtiQ7pNnrc8fvDNlQSAPfhsT8cSgHcAhmSMW0FADFA9xl2LG12Zq8n2OwH
lvSUGkiREDU40gn9l5m3SohyfdQ0DySLcnluyoXI2gRbVPnRgPArX2qarfHwDNyY
NjZITKGjs20kQjbRSYPQ/Yu9uK1S9pLxHJY5CWX6zLuXY/9ug3lFHlVSgpQDdP3P
SI+FeuHCbXTY8iApo52P37977ahcVduHyOh3Qz/L5BKq89kBCsV6So4AJ7bAfQux
cLBw3FSVNpv8qANoQUbWITcdaUSlDtYND+Iw2ITKs3uSN2Bl6XEWeIeQA806i3Ti
QPXwQmQAet7TBbGIQy3Xq8vcb8cKq+9BhwiQPL/S9ANVDoZ6D+gsa4bWSMcl7uQ5
oC+ZANBE9WUt3VyJmzRXA91t4XBKv31FwKusDcHbBx8NErrqoLbzU8V5FBfizsBS
EoQlfAc5cV3EYp921mdhPvNRjMyVBYeB4ILrMMPMFpdDP+/oNcMhgIfxx3uh1Nvc
gU9KevpeMkBj/8shW8wMNiWQ9ScCnf1FtT3h7WjScF2zoctLsSwt4PuTRjsaApH8
xu4AVJCOuXmXc6/5o6qbwkhQKtwr+QbNcs19l3HgCc9bHdFAmwSrT2100lh0jGu8
GrYbJcbz3hI6VbNcpym+KCAwLtNnEpZVhXKrOmIpyq+uvGWYU1jQsV0OKY4S5XxZ
JM6nRetENfBv1Pcl15WNMq5An8fMcGjl+WD92r71t1hfT8J7XTKa+Ts9lDHFoOcY
PaJYJ8+tgMyjBq7PD++1b0Jvrj2Vp/zcV8kGeC8yXThZxRhJvOKO0rNSmCjEMk+o
N2brGgM0bZk7qF6DA329/W1HqrC0coBqdFRv9ZzaONZIRLaeFYYadLEKfhcXafnk
mQkW+JEzEAf4dUq5VhH5oiNQmX/s8IiH1KIKjQo/ZYiiAyZ1qyebvU7Z2NzsScpF
Mlad+w9Q9VY3hUH9qTSxZa1Mo6zRs/qSCNy+JjlZ/KDaVtHGbxloERN5uU153tx7
rcrGkYwl7PHyZF/8pYQUdNKVWdSVT0xWSMXEyDJ4+Ora1Et52k4qzrpY9iBAtsOj
XkS0iCa2M1cm9lJuJqXz10cCMqyrkpD8vsxQKCJRuDOKw95TLPDsnOl0SAtoNEL6
YNtWQCnWiQzzQhZcWDgYq57VJDn5ATmTPAujOxfi8Wk3mUVR9/JKQ0YUdRxDPhbm
V0Ku6NKLocdX9yzQpL/NZRXKEvbthti90twVAWPJi8bYRoIIYW3FrbXJXvfr2Owt
BQJjbCSwWRtdrKSzzTUJboQflSFjQhj4fgCMWWoNds6/MoNdweImz54MpSOpQlC5
r6SUZF2NfSJDz9uMjOEe+8JdXdODOU8hQfz1gQXUwP+TRmCEejPJioFHFLW4rVhk
UGlf4iqH7kMLUQLIcXtEW+qDCGb8M488HreAUwZw9gbWFKYBm2kYvvWLuLF9XBbe
pO8BBEru+UCyT5UbVPb8ELBJeVG6A3GwHVwHdZu8DGvQ42UupDnlNAb/kX4upv9x
eEO0nfyGRq5GtoK1qAamGI0UX71um/mYkg2dOO34skjDT2S5xlQuxkni8HBU5qtV
3mYi7ZiS51KkYAar/mfAa8TImDh6XCj380TK4El8cDhql4XeNKnjzY/Kk4ifzj+a
kaZn8a6d2/DwnxCQuajxHkg8ePAckDR5VWirjAGvu8nHOghyuB0P0lMf3iYuWsQd
dtpICEPw9xKxyz2Xi2+MvjGi/VFL2u4zaX3oQB9x4t4K2VYspD/OMV29m8MI9HQb
NUIjN5Sq+G+R0KY3wI+v9DubNlRl2JMWECx5sPH06MRXmnNTwRhwyH6QqiY5DELJ
S61VAcVDa4Q4YW4LEV6zjOkaS6C41kJZ36xox1rzBSeEWA43XQFdYuKw9R9z51jP
Y0fTon56heLZsvanbkUIj8vyqPZ0+zYRWyU7m/Rj9i4nOpavrvAlH+lmZSTIRRdL
VCMiK5JyTGh8R4L1mtQo9oJOL5j/J7pDbv+F/wAvTlW7ureFOt/LZGdyMt8gmy7/
jM4xBckqchi5cRClnYZTne02lStDVI0fYXaAukK6wbYf8SBobe+TVLvg+AFNyD3Y
h76QZzsA6t12avxTOREPJ4Q05Zy/6EVudyeTXN/3UzHIAAYLb49ETmz7SXU/Ib//
skd2heZyDrm/OOvo5SGoSb7mF6Bf+44ZUlO4UqL/lo43cJheRnSNtK7iE7nGwP/e
RDTWOyp3yJEQEDz/0zSE0fvTg/ZYXWb3yPDMQi536ewtFV+ejgHINbAPlo6LoEnY
EOvhRhY2Ge9yWnmUTkQQSfyOXeYNSIAj6ULNW8Vdb2Dr+VGPsaWNQrYWGV9dENif
ybxAehMJh7YkDYwzhyZ7tiKvgYkiznxjAleMUvX9L6ErMcR3roh0JixFVTw6mBOR
H0WvhC0AIEpaJTTeX9myCuw85/hUV0kSV/0IPdufUh/Kr/AkW8E6IolnNCkGmBOM
EDOiROr4ARQ7GJsyNaE/jZqjeqtYGxh/8KKknWo+zqJIpl5/oEHx5MdU/dE13aD9
PxyD6JP7BWty6X4iZO/aOcCwyGeX//a9iJsxGDadvZ/8+P3d+BvdtZUuZVJLF9on
UyNs65X4n+Aj0X8qRxqnSRLse58unN1nrlBg4POyPZthcfG1przZjZNDQtrjJkYE
AF5jXanNdpEOM3avBl6rTt9qOv70nhoz3m7OfomZpw+GpfsNUm0N3bwfdBY+SoWy
yRjSA1Lk32VpQMgvSV4sAlkU2kRNYfvh6v6CieANu4l9AdMoNCJACFhgRWk8QyaR
CMArGVGUrTR5HXH4Q5YEhpR1wM2O4zcaomucAJKxwRsuMuNeT9xJn2Sjgh786pgI
uVu9wOhnF8ejUc1i0PKqpHcpAFOJelmH29hL5tieF6yA1bkFncKpQmJDzBbDq9fd
25s+Fc4veHfC0gd9HUfxJKa3i9m+RbNQoF0srGJypv0h+ebTlX0DlLZoCuVl63FX
AtSFBzvJUsFUkdT/v5IJLy3LXx+p60LJWnjDEnAKEMULJYlRDBVjfUanEYpNsopz
vPd41R798q99lVeoGCceRS1uFjikK3J/J1I4hR4jf6iSkroBhTsR2LjrJ4PSHiKg
Qr1TipMZt1ofjb0HyZw0Al8fWoYASj92T+1zj8itb1MPszwixKigeGQKJELjjdn4
dayhT+oXdfupcx8Vh06vNPYjle8bbwGxDeZkedYArzMbrJXxfkChTFdWG1+vw7MH
jLjzQOqLyg1+dE5SpMtJAQj/ZZ76qIflWlZDYga2EbOnh47I/Qc+ZuOkzxUbifeL
TKM4+eG652hJXZn1A7/QKP63H7b5wW9sTNA9W75SUVq1hcWY3NkdBVFmspNnJ/8J
fB3iNP8KOHcIP5jwDlETGhPHbMgob9Ffc+8kbaqUjdgdIhcIVkaOAjCdf02BfXe7
Ho6zX3QgttjddB3KaK08VFyhSVw0i/OSiRmOKDM8kOoVNDQzHgxQ7GhPH5ELUMYU
4VuKTpQloIBJoCQ0VI24jcoQO4w9b/CTk7MPESsH4EfvmX75MTjdrlRVbkod2Zr6
yBV74L+EHEC/2sk5VflnFgcebMXfrPVb7rqI8btUtfa2jQHDmqZq2ano37b6U3RF
JtrqSd6/ySTvblvRXZE0NGtH7kG7Rsvg8ejo7bnAMf0OcZsWqEW05Wx4gfPP7r1n
0zve/nTv6g7pqunKYu+RaLyKm+HIzLbloVYLjlWYcAH8M91Mlv2ro7CVEF/hJuDF
sXS1wUKXDJ6RcgXL1GrSrNJLnGesoQC2Yd1Caxf0sTdgOrizZedsQM3Czgi8aBJj
hS68YDzHZrTXLVMvi2rsSE+63DJPz/BVgxC/stTjkklCrMW/81lerAPFAhIyOwDK
i1yuZ87jCr7iB1bDCuvc83qtCks8yp52v0U4xNKRUfVfSx0xv+kbeKAooSuc1QEj
XVkqt62kQdltgNDR+MWTG0T89ZjQSAzw0PiAYXkXA3Aho754iwfHPrK/vLToUS/B
SAxZQAfOiQSJSN/wbfjcNYtb2We+ZhKDm+0sgJUluF0vz/sQwRgqn6Kj88Ji5Xsk
8n33GBuU/HqXYuWzykZA7IHl59QJiIzklmKMmsCu2Qtfyurl2NdoUjdxnleqUJor
QObJLcB/JDlDZwO1R1Zf4AY2bPiZ1rhDCp1whH6L7YIVGLEfFVnysKFOj9vu/m59
BN11qV2Lqml2KvQQ59d5Lfl66obv3WxhZGxpviI+iGK40Yd1AwXrribvxopBCFed
UV56hujEeY4Y6Kjsw9eFkXwmSz7aUqXsHPf5EZ/pYTHU5CriHmhslfScBqI+rlOH
B8p5xzooa4sZUjiCP3BXiC130Of0GpRLPmXtzQwD8sNhPtNRFKJi8go8O+wwx1Xg
r2sC5uUJdVa/N26eo8wWaI0OOolO6WHrEVNdJLft2IvaLiHiS24aiK4xq32GOh/a
FtH1zX3vf4yV1XSXJ6zqdfX6P/+3jLqcP5CeBnp0ofQM9RygPvfVAj/PK5GTU4gy
9VFLdFZHt7MX/PD5UeIWpbPrRdg6WzeM/GTV6W5h0RO7Ys7XcycG/SkQNHZ24klm
7rqKossxDkXYvlNb7jx4yqsaeuYuLQB5/8WGlj3hGaNTO+vqLkLQtPOl8FpkRnG6
dnQ+20tR4JW6m+qRGRhBR8cucypsUBzhPjGCQDZBGdvJdr0SnMfua1uuu43E8ERn
NM43aY/rdSamypwF66t5JDaN62v0HIW7PXV3Y44wVS/CZ/hm7z3vJtXR5PyOSl8Z
w2ylZXJUdzMPpb19SQTqz0DCpqiqPGwlBUe4CPwDr69WFl3bOVC+fpTcTjcro58R
EXqDVH3bJdVNjuqwP5jzZfCApMtcb0UAK1sPN2kIcvda2Sngp+8kPeASxNfp2rvM
Dw1s4+8CbXKgLq/xiGDmkZHPL2g0svZK0IT2SD3PROqCgeHPg3XnnFFv7KXP0ujW
UCT2LBpY22nX6UNJSOmQ/eAbfz6vfCfr6EcMyuTc44+/geh6n/EQuxLjeRNYrMtU
UziTk+ZwNNXi4QsVJqxJab0FdFyWiJ1JXsfMLnnzjf51EXnOw7qOXp4Wv4a8o0W5
0Z1cPsud6lzW/MZ86qBrWP6o/iNHP1e9SRoZ4CyChqUV3PXqJjjhyieoqyuQ0Neb
96HarPEZ9r41fGfKLrDt1vzIGZRAlONkkU8U31Ms33h4NMkQwNPZsu/iBx/rvv5B
dVHjtg132aO9Eo/pw/GRhA4UMyiwGwSvmJtJd2yOmjaXqF7Hv5lSiw7f4o/nhEW1
tRnAA4UIkOv/QwX9N/+V1aP2njWUGYMi+b5B3/ito1q6LsLH9isDAY29C6/daH1f
VrbNhBwG+4CjzdMo2wXFrfTVt+ms7R2Sbz5AqSdnpIW+pTq1Mti+pk1cHUkmQdqQ
uHC7OxAnrSdupNp9jDmesAprDaIrViiJhjmuTYsmniJmr3bYRqJYcs2L9/P9bOVB
igtpsAoD2mk/X9/0jcYqdSdWwmojV7xUnwOPwoP57CGZDNQTH60H/fKoU02GPets
Q5XkPdKZj64JMCq+vkgGeogewfASdHHl7831qcRLY7oQk08n1g+5dcoOKcA1C8eQ
M0bI+rPUhTww+hs4sEBrthas6dIy2dH6lV1lbWbK7X1GPA9J+Pm/nV0HWuUuWkVR
tjciNKZmu3Uy4LPZpqy06+g5vUnP563+h8u58E2iO3T4qiydIbYXg91YuDskn1rJ
r/VkmypDORrlY9c2cueP+vrq64am6TqSZf2c7xYOv4UUvaQfmDgMpuYNXyI4PXhR
ghXdfEyDBPAl9b0ZpHtoJ//S/Q840LZQ3qJNVAht84MY9ujiSOFmYhUv2A642MTT
i4Fqj/LphPNsvzzl2n4yKH/2TDKXTyOe0Hsn4ZXT2cDhPs6tw2BkLja1ljzVXBqM
ojBDcsmzeJWZvsuzz86CQgDBQ0ju2bGF8kseNJ2OUmm00CogGjtC3+1Rw2IFHoJa
KY2+y4ls7tKKgZbdo3Dq4HU7IgJXpph37CjgQnLkY+rdVsdLS8kQX5jIDcZ69DvA
zJlWAUmShiQaBRyPjVjuPKmxdU/8ndaQ5o28bAomskAT5FesGjocTAeuJjBRdmmU
4g1vfwJKiWd/wTkbQGycpHYdxIAuOkLqE0r3hD35E1EAuTuvcU/S5uyt9nhoprYC
75rBRawcnSPmSA2Y1iz7hy9m+yBa+Q3rzixY6vIvoRrsE3WHW1fp4FumyHjUJI1j
kdLbRa+AlD3QAZ2zi7MRPzN+pqpuyUUgzU9sAW7+WNGB6DosyW9fV/cfLW1xYk8i
4EsAztVHI285D38nueaQjfDcuo5BgBd15VmP+4ORLIw/we8021vLqcCfFn3Ww1Wi
ZoBNvPouGbNkyA/fuJ+jM4t2lSwtUC6zkjSAGcTrqh7gbrVVKAFQ/ixV4L5sGXy2
JwgbTRNevOvG3X1cp3aIJX5/Bs0esva1Z4gFSGsvjQcUXg6X8S2Rus/5FmvhI6Xc
a1sWhmJ8kbLjKveOqBeSvg8Ol2XD/IiZirOfD0s8JInmToXOkUlL+tpa4Rx68A5a
8h8BxeSODd6Hl4k9OilrcqNJoFKTd9lzTko8snm29C40MSLrOfuocgGysOM2wMyf
CF6mkmPTR57Mpnkcx9UIkVH2X2EHA709uZyqEowE8tBZsJ/zXNp4wIiU05ggQBCB
NKSDOslMCVbc5zCJSJ7hedlJk5j9YxulF+hNx2NxSU1K4cFoKAm2/nJSW11dWA84
DMODiaW05/eXNKi6D+O69/B7c1tD/e39u3a68u2mi1k+GKYGAiQj3u1IvSugkyX6
tltSj3WGw4lGlqRMGyjtaDz33sjEjJkiq03iZ/o7paJK7jaeALec7Ii7nw70hPfF
bNrfdA0def+gduk+lJ6b0dchmaWm36YqjZWEFmSPmeT/X2lzQ7rA3xp76D9txw7U
uhH8hsdC/njDvwB7+umekpzxRKhGYqGOI9xzcNSIGv3jINZkzc7Wg9X7FyPs0xD8
f3/lHltvXZ0dxlg8A62U4lHsk6BHGjPv73+jaoWazM/4hpGSlzcW4LtiaAbNvi3J
s34sgVOgIjBRjjI/TpXgCOpkloWCgObj/T/F2wbQ/ylTIgmtzA4FpdkjABj5tkfN
G25fpENTVgKgmbOmZV2X2NmX25K4xpcS14w1WXDfd9GV6SKQ40lXkN3tSuNns/sF
qZQhisMWnzZBOjOgIDbgu+/5ojsY9RfCUVu2aaCAfxRSEDaeE8INa5vvZibES9ZB
LrymURUdY/XuHAlbzN4+HyAByPUGu/Yr+UQgsOuPfUrwD0Au8zXbdN92nrPrsZKf
mdCHsVGZ61Dz6MUrNbo0X6mFZUjOD6d7f3mFNWwEv9I0irJd/WLouL3oxJffvRgC
BDQk8vKzUA680AG76CgWzyNXG4K8NNA9azSZrLo2vwhw2nX5Bo2y5QjkFV4mVgG4
D37RWlKZ935njjAHFZbZw6oqk0Zb0lvEvnX06ZD+Bm5FqgdQWNqSX2Uvrb9sLsU7
R+EVGW8+ZKRXx0VRiMNF6dsipN7kEbzxJE+trIBkQ7HRj4Pk4OAvL8LpLbI2N/dr
heo5A0A6fWtUUlHjq0phrjuuTqyXNAMmUefZNdn79CA4jKXivtG3gDk0WfgNG0eQ
Gucewb/6wHWbva17MpCDZc7pu6tO1mN7XOQbNDuAWqDr+uimvVA0QjwlETkRl8mS
lVyCb5+QL7Z5cmBC6XnTAj7xdnuS8z7rb+C78MW+0HYVO7y15m5SS8iXFfLVSNIq
Y3hnhfyhRQn8P0vh5/FefNwwF5Z+y3rf4W0uI/AFzmju0L/6W7Bpj+7wfrH9TNej
69OLysKXOdsW88FjwbbFgDhZUR+P0/tODQEb42Jx3tfGD2BH1drMsVeb6S4K/auN
8Q47c5i/2mPZt60/EGGuRP5D4DJR8beRevHSVuO1jhhTDyu74ntMiu5WMBTsFEQZ
ZOyHNzA/MWO2In7TyZV5qSXP7HU/sX8o4gDRcGATnMP/gguywM5Eb+oXPJAtaKsc
XCRTEAG81smQACzqfATS6IPpU+w7FQP75uB96GImt2zPHKmWfMdxHPf8DJMWkGBJ
fBtok7cSFTrNm6Oenw6uT11SNcAG2Q/exbeFyOdc7nHphCdHVwjhFaYei6sFwVGa
Lw1EgbJBuj1cdDcNvu+P2UiQl4dUR3gacrHota4nQ81B53OmsJVcAC03vlaSpFmo
K1sbhw56L/YMQnLGFBiGonBjh+B17pNdVN3x73NHDgkpvhYL3kp86NjIZA6cRjyf
qPayZiYzQGc1WxSQXZMvKW9FQxwGHe1cBR88F1XSSOyqoYfTXTZoS9Ro8fo+MNSi
IBReDlHTworDOnDtGJ6iHQ5r/mvaqRLNnEi0Th6L6YurquZAI05pDW6XAmNC+zW+
QNa2LkI7yEzbVlqYhUQ4B3p7hUuz8HDUV7IafsLLl7jDB1Cjcna1fCImWrlns5EA
EgdeUsq0NPHoHIJZ2cjqMvMD8oUvaJuPIwK5EMf3VxrOOzsQ7GTy+TEYIbJF+i3d
VjA9IdcTrC0/3EGiM5fHjDSnM+neJRyYGvSWgGH5Sv+qf/bl1EtnBa/VXQGjidKB
bnmg8per8itnchmg5pCZ3sS1/CLmaLjEMXrxohDzW5x/uwl8VQTk4rgb0inwhgl8
M4NoE4EhPllMEKhpb7+s2ezApaV57fFQy8QA3uL+Sgwc4TOfqKGYoP9i9ogHwkvd
dU6/DmxNK8meG0h1Fz5Bu2bizovYi/FmMgbicXhcABGXuLJ0AuZBBqO6C69N0gG2
v1OG+WfQqrMkZEoTq+Luo2vsb5OFsKC6EprEiIhR+qoRNWq0Sar0sbjZ9RZCbA1r
VhWTYQe8aMG3wCvuT7TBdD7H1mRk2IbpbrQcf9ELSArOUdgZPEKPsq5D9Mx2n20n
uqI72qs72krY++IcszeMCoqif4d9VEa7xbz7dMuEVutZXbLyrgfY8+k+pqOzbLC/
On+HvuWSWknafpa5VTp7AukCG0gImklLHSE7EGl77TmdTOkQyuQzCrE1YjLhCSg2
PSIm0M15iwgvig8TytR9RjbyA/alCTYNOut/abGXUr+4ajrps4h7ZX4IECpQOLsY
AEYuxsisB9vHCnC3JjXqSd/107lqkT+RNO49XW2hBXT9ly/O7pkj2FRLoSLx9g6B
SSxhGxstt4h4WCIqNt0ny/iYOyf46TM4o9tkqGpQa8gv03hfTSFymj+1CeHu+s1u
sh3KXJx4eoXwJ4/2C8n/4tsZfmV3GzR37mI+VBPxxbqxS5oK9yK0X8pcZgj+ONjI
AnQ0sorMUE91O7mtaoVBMNBodfHP3p5XduAp1QxnEvfc5XB8mCkrttAS0WeT0puh
fM87BBgFM0e6HRR0elWcEyl+2LXklivklLc79B8MVoMQnaRuk9/zRcdWDqqIEAtB
qYN7VR65k9+3IKEGq79zyKoA3oSr4dIGRgLfvAAyJtLe6bReb+Sw9cY7Ztr+Q060
7ITKCO6wja+1mjYxvyurWi9dkLs1BFml9TQoX9gToP52mjVXnhbO+Y7YDIZmECQo
G7qCD8oAz8CvNO7juDduQeofVEmP8n8Pdjyi7OOd34pKqvWS29HAIKP5iCuSzV4Q
I+fzAs7xQ3QxenyxXzA524JLf/cAN8Rcj2iuSCd/ImRlRsD6LCISRJYGYwtOqlYT
b8CXJKI5DFezbe50+IArmytyJlqJV7AXKQ2nB1G3rIjObXCeOcisZkVLUwQluAyl
vsundFVQkdzxRia0D5MP9mE6iZyuhcn2JeYMlgO4zMPcDnzUCe0YkRNcdE0xX8L3
RGutBVb4JMdiqZPBJtzxuLZLsIdTJrPGcGiUYyrCxBZ6v0lHJJlgKXavyUjHnYZy
Rdnkxb6L9mfCaj6unruBZJvF4/UIErduE9/c3o2Obgpxem56G42tDi/e7+6lfjja
AmidBY9UDVLqKdGn2ZtMkwJRWlzoTk5OZkDJwFVrDCjoQrz28dVyTh3b7YEAjmmm
9lL4Ql0XD6stHV3tPqNUnTkxbaNXcY4QfkaoABHZawt/0xXMPU2PIkdL7+AVn10g
qJ9BxTHyIt6zkz6tLdmF8R7SIGRw8USFdj405otneNCnKfcc7AjWv/A94rtswjNj
CfgE4I/m5y8XN8MtCCP67yiNp0fCV8AnHSmAZgKRvLCj7vQ27xWSpLyW9rWRkrvv
vJv92mEUlSZGL9usw9St7lZE/d6jI7j9Acdme06yh8WXEUA++aH9ZBUqMUiWgCIt
PgMTG+xcSskv40sYlIpGvKEFBEODE0M/eAav3C64YMR+AtNR5oCxLPx17LQZ8tC5
RFdnqxQQ84iAng/u8QSIfzjei5NQzH9Kd0JZSuPiRGMkmdKCvymYa7yax2V7Gaa7
mZiB0C5ZstPSrHsOWlaEyBR2X6lMFE1TxTiYrMmJZphNnvRY4JoCc0doSwQqpvu/
VPCYE/v+AVO6Xq4bIt/xDcZUGgQcqJ/jwSI957C0WkKOKPnpU9EDDo8bymzpnsTQ
/+jgOOUjy8iiYTYUe2oH4+EV+G9DC2hQi4l8Mhe4hktifvPmh+NbPjylxAN6V/Jv
KGn74lxfqWeqNcL0C1OTKVikDoXilFrfur9KuCowqXqZYCN42c/TuSLHCSPvmiPb
JMQSi4KPdEdk0Wi75CoTIxNDpJLJoNP0W9lOoNDfuVmkvsmXAFd/vF29TRQV9n0n
bmDN0CejEFWoGnzyZXzoPHQ79AY/ElZ4VO6eVRReAzkZSioR01qED/m17oqo1Yj5
YARvUcV0nFWwDpbbyxXkCr2Cxzh7kt6ss3iZpjIcjerhayyMVX4PNDbXPJiOQfNh
lRnrBcquE2ZI51bsiY66thSxyW9AiNJE+qRN4X6Ov7aYKns4itQsFN6965dcXFLl
viuCuZGT372DvQOgKbXmEr9mbZN8vCp+0vXrK4b4MT42ayRMNIcNes55Et2ccOkK
nUWBsF6pS/UTs6sZ0YaHDlZQDnjO2YhIoLIMNDbpT1SQH/YqxLhTgMj9BXl6hNA4
0DTo1uLdpmroq5qURwmH6tUOqGP0z8uCTN7CJD+rw4wGGhDsDG4QRZqi75y/icFT
WV4D3hv9isr1iA1aL3wdnzbLp6zboafymp9V5YZdF2lXeQvGMIx25r4EqGIbgOGB
3rTgQkQgvE5SrlyOS6xsd7WK1rHT94AYUzW/nKouSNgbjC1WLdTb8+IqF7pyGVgs
mU36j5MSGyCjR9arqRVDEX4qNZwmN9lIEhJSkwkRkAPjG49ly1GeQLpIBrCcM2sU
rxNLevvnhv7louF6rhdUPYHEqyjqBdksl4CTEWDXsjpYJMzG82tO+tlxaqqVBgA6
HMTwPQZmAEzHsabK2/x0JTuJQQJlbZgOQTcmvNk8WOCJWYFJc6pa2YlBikWBTzum
gqVvWQlBLiy/vFB7lyCsb9nLePfAzjTBWXjE/a0GTMbk/pVlyRNOgsLt2L3kpuT+
11m3VXai7m8JfFg5rkGu4qh4iYd31fN/eqZh/Ys7SNpQbLnqkvpj5AlCtGVW1TVi
tfnFK/Yds/cJfJYKVmlHlfjFoJv4HY9jeR4WGv98pnMlPUVEbJsar3NPN6VUNW6A
DfQcSGTvBFkQTx9u+aa3EGmKhkg5rg+qGx0GFttFeuvx9NGn1jIH2/T1mZguwsD2
gGa5UAVY7YJr9tY1unUD5Dxn/1natvL5uMfbnKaJSEr2IezDfxSqFD/I2jMjrwmD
5JLU3IIVQ5/gc2F53yR6lyZLF44w60Ffix3xLf4R9ykKS9+pBxuDSdfAOSYwhFD6
mUt3+u8ta7Aa39iQCVsyU9IYXdysIDTjGFK4ES2y2SMFsX7UH1YP3N7N4s1g2L2n
jz1rUeD5iEAE03FFCc9ZReJGgFhWzwe9O/xsHbZteHfEOxc+NcctHhMKCRq1QtEo
E/qRfHQPM4EeKEToN2TAyz/bFTQcVH/M0foJXUtnpGGguNWAfZKsXbpXMWwHfftx
2Ny7+WTxyZKljAdVxWv+ceY2pEQ8/uk+R3PbS1+dHMWxUFD9gr3EIqWljECVGyUC
fowRh/dpKSXskI9Kve+qV4gEHJBZ9n8NhBLcgXR8LZv6ITYZET2CU2/Q5CCZtrCV
Vly094oA2xHtF6FrOWdzd+vxqcoxQc3Ufma9zpdKgH2jml/OSCNuVrKkwRFfTJ4+
C1w7Om0p3tRDU4+/7PMT7g1L1dxA/wCb8ZNWHGD91eO4IBluMvCBXHF9CctY/o2e
3566WeF6lXIiz8QnBuNEbUIpfGJVWAtIK4gJY+b7Gip0ukPmUTmxK1pIztOWm+Mw
A9IYAY4s4/X8gBAaOGm/6GKwRjm4Tg/ls0p9hguHHRFQAmsOROJ36VaDA0/lXXWC
blYDDw8IxA1THnBZhTRlWcKui1I8de9ZEmaH7/aUEhx+zHR0GA7nQB/AyI1gRvTm
KxIWI6z012PqSolz3htFYqheKJRl06ctCTzTonExCpItm4Lt4YCf+yfEbTAI8aIf
IMfQLiF4AKAsASY1qOpMJbFfYwgpHqRqkiv4i8V2AgCho3zb646PX/OgGtSd8Jr8
yGF0EVSIGkABDP0zK9jwMp3A+WhYhsA421tyCnS0bkaeKuEBurRnPVQ67AjiCvAw
f4aZHN4HA24pH83t6Nfs+lyvY8jAie4uA4PltrN0dxB8ffgF+4lq2ecu4N19/qcT
OSGrlrQEuXsvhpKr2mwlEPzYxbgjDlOthqDunq7tYNZN8QK+Y5av4swnHuA9yioS
5Iya5YQPd5SEp/CYspDTOlDKojoAhFKvJEL1XzfXSxwkHbMYvKHA0q9tL0/6iQnU
lhM3r2ZRXjyBK+A7a9MsTkF/Z0NJDqvR6zMY5d8G6vuper6qnjqN8dyLVb0naarA
hl9Ly0DdYdnJMDuoUSwu4oxgnFvNHzltqURWtTN8B3gkdTkIqkbmI1JSFoLG/rYi
ZEg6Ukkpom3yqikht4PcXIataFIhy6tyCoAKDCdkxzNjoKY1qKEpM2AVUOT1t+Gb
kaJD3FVUbGx/7s2KnAOywvntmKNaIF7tEhoZljEcTa47TBsEbd+DBEiDWuewIZrQ
Z1lyoNm2Xhc1CdvGInGj6r1hqLcSN0aswQpBMsxhk3MlG85nPhAfuOgHh57RHFv1
99jEPXcLREPJVEbYARbeBIpnWx20VVLb/LGqDLIXcpQTz9nfNMWLHCq/uA5L9DyY
du7IfOmdJ0CLKHoungeKBrGS0+Pt9D3Dul2K/NcUracqGgN7zVB2dMElYEeWdFA3
yInWzllESd5CpPWJ4PqfW2JW761vQOg2fZXcZBfYDXXo5yvxiW1LeCfEgQgwE3DQ
5DOQ0RtLDWvk6S2lwk5oQOaEr6RxNat3Sr6RBWRE58yXeQzBXsBhKtNwONKpy0VN
AxSDz+RIMfKPUdoLd6SqPqHxb7vVi5gPACTAC6kRLVYEoq+C5LtYlSFCCukFnj54
cY9/bEF8vWIbqmfnOCU3XPdKpTlu4PDSkjLi9MODrv5X8/VGQZmU1pF63nl2ySwR
lG/3nPU2mno8TzOufWMFh19+dZstokJhcOW6r8SQ1/WijgywUSyyIbymMak50aU/
Sp8ycss6LdGaoEZB9fydYq1akcg3nusq1sNq0Bu/NZOg4pIk/RZg5y+cBu2wojGJ
EupyhuWPQ3TBy8jGT6/mKEACRg6yRdg+4hi7HBUVpjMNKYS2k0MSzSQ+Fh/Xqtfx
/KcbCJ9t23eKXnRLmmtFTN3lBwMqJMiKczHkhG/CjxYGthmNtVbabP82my+fqM8j
ltlrLdRrFSuCFo6gBQEdGvNwYUps6YmU+EygE7x1j8TbHBk9o09FBog82ArGqi8X
O9YuDTrIk2M3uXel1GeUgGzCBlHcyvkuTawiTjcFOT2EOcWWMn4UKn47sie5A9lv
/6tZRrTst1hNukGKfiHVSp7p2TyquYCMe/p9gxnSdp+Fbs1pMVqSskS4RblzwUKS
d/GkmzBZBf0itKMAIoVF4TKFMaRTXdAYxyhu4Xw21lLSmjk5jJOWtzzE5LacXy2A
dE9mitzi7447AcRy/x9bM0FmO4FYR+XkEmI2G6/VOs+wCsUA+RyQxMJIlK4T/i68
1DViVLO63/q0EOb0Pe1ou2CRqUuY2iFtdSjVkpc60cTzFNkeJWxnC0wJ8Ndj6O5d
iZFObFoC8ZD+/76Pycf8t52rOlRiyf1p9tC9vcSShxlPlW+mkNvZreNF4526U4E7
GoIt4nmlrFAu+71ZJT6FQ3fJpxJsD+Gdk+9eEu9lgeMc1aI6O0ffCQA4l1lOGYgz
BOGR325pZeS4rohZW8GtwTdRBWj0Uoo7Lpt+hDA3iTOToYkHifDTr82VMckoW71i
ziKx1Kn9t8CcqaC6oGcu2Cl9WA8hbfFcN6szR2NWID7Yvgwnqv1GkHhUK7xjLuiu
6z4TjlI5rTgZlNi4GtiJZP1QYxTX/Nqe0T/M0IpRRi55o70snKrOuRfMBOOvkQ7z
a9kDjLdV6+NLWWTwVAP1SN+StkRTD0nVa9X4TFVfRVlcLSJfNRKix8ULrMaPTEO9
vd/rKTJwZj1CvazsbBTwX7nxUjOhyYDysADRlvsCVgk+GW72wNEi1lXJwddBNF8A
ZxxfPe8z7aMckA7LZkOdbuyQv5+oc/XyPn5h4aRJBg0ZGX2hA7j0QtaJ7eVGpXX0
F7JkLQW05HK/KrqKjSsoR/QRakDNvOLQyTYKWfrqQkMmn+JjqLG3LKGPq1PTINbv
a28xoSUCHWahneSJte9PsZGGWcNdFYKY1vdVNhOE180fLfL12X+ruppRvta7c4EZ
enk7kAlCVEPrVUQQimWPXu7oVPDcoQb4GZuLoj+ARfGjmxwJly+CWBm6j1Lku9PH
P4LtgPkM30JKFeQdeK546+ltLIR/hyn9ytwp/Qigbq107MxyyR6rxE1GeFcvElyv
hsuMHV3l034YlSnurmlCMfyoaQ+cmAfxsFP4PgGXOSwD+UwOzZ41dV85ceHJ61dv
Qd1fiz3TOyG+H9c/CuMWnOs6ltTzFEl4+x2fwWt2TBp8rxifSM1deAH6kHjvdbg5
dGu/VcJUqNHjcY14fXzoxmBFL1CRXuCbSuknJEjGo1V/SveifkiCqt0w5LxTS77A
BhVQeKEImWXmUYEh4HlDd6USiqiWr9QgMxxhKxf6dM6eWTWOH6sZYr+883bwhU4u
jp3GPJCTEPMaYiXlf8LckbTiVVSW2ZLV27n+4oehNQl8TlrL7++EaLMG/EmkKW7Y
Ocrep+hvXv/c09Ta+2yjJ5XA7MDZxRWH6yXVSSXQN6Q3xTiEAOtpFpeeCP+SPUYb
uf8WTfSZBi3nbAYJl8xjrb73F5J1Y6jPcsB0CxOfpjy89x6BIS85ULaq31xjZcT5
U5ZEze1ihE/5LP1ktTrf27kLaLgZXyGDvA7NPOJjIZ9o4Z8IHiOAO1o0p0qb6XxL
hrG++wYruTe2in5FyE1uucB8XpM4MZqFO75alFnr7vQSuhLfwQRfv6DvdVajX9dx
lxs3v/nNJHIcmDqUN1kQMKsoNMvSVfyZs+9+4tfW2FMBpY8kxO6xyJacA3+f3Q9F
NjA/88WK6PN18VH72Onvq3wRu4vOODtR/LeGfefP/leftMdfmeWluL4uBqOSufih
qS7z45fYoFE8A0VMbHcjYDPRrKARxBL89t/OAVOr7BDXXpIZ4rksKJpGyNtvY7Jn
+EgGs4u8/KO7BwIFztCx0Q9TexGffV4G8p2mKIZVaGE+pgpKSVOjLNk5ktxYBk8N
VBVuPlGSnYsFf6837X+AduVd49e6XoRZGDP+wRbXcjbxbEsdXRNnnqRXxK0BSk/U
fv60yng8PoTCDBpWgcQ/6uP/5Gf0KxKq1nvkf9SCoR5Pk3DsgIaXCr3/F0mIkfQz
ZvbqgiBY2zoydCeDZmERHp/NSCIcYUxqV4U0jFUfsoff0eWKDarklybbSR3gH44a
By9KmhhlyYeY4Uwp6Ln8J7gK52lCTfSs8oZCB8XtOqE0NrEdWQIXODrmprJ513/T
uxJKnHhpuhgCWygrnQ5DeQ9jzRYz6FX/SMmluAcabhwZYPSU2PXTG7NGoe+Z4t0i
zWQCwLy7XYN1Ky7QdXTiOWb7zQOnZYNkoCkmA/Dh7tbOdr3GnimarFgJxjUNhfTU
/sxVr6eWg+ppo8VIvpvn6rtIX0tYxdrfsP4cOzsltMXUsUTX2lKFOYKNiW+ZL4TU
lkSEkLlpgVlGgLkPj/P1YGewkOT0HCwgwo8lGZqmMIpj+bC1NCZx/smNld/bYoDX
yUNtItAbfbEVSgIQ8vJup5KRFnszVo6f8hyRx2CLO0W6+8HF1L0hW5w9D26V1ILE
6uErkYD5boktMByMpfOmT/fDm+vDCfBCjy/BSurwAAENb7aKCEaRynsBhk6HEnx9
C9xyhWJ5swh7SOgWW3ZcvbeydORRMMrVSh7UiZ1Nn/k1fho07Ta5ookeLsUtUTD5
F93TUDG6wkMymfVqrNmxFjwT7jFo06RG9nhfwa+g7peoi3wcAkFOam9GjPu+MlUH
ufkXvFC/yWZyvwuPhJxlSw3pO5FsCuQ75NgNOQihKQHavSU4XqzdCD9mGdMwk7e8
awaRezkeaqdKpx57Z7xIpi5CE3gSN8GfHgsL9hTb61OoTElsQ84iaMnLxfhMq+Xh
12WlN33CT3dvGcnlnv1YuEDkpkb+b/LAy+oSxaW0ndbjIQAt79DvwKFGPCK3Uk4X
hMuj0ejQwaiXcX6I1a8MT18hiwybVLqNXxB60/lZjXvdPgHC7xOl5aChbm0wlv9b
KfubEbVtZJsExxkP0K9ogj++kVX8mlXFtmCKEH2WoA8TbxuUXo7kf06W1Rn3FN+W
Dl6HYfbE7E2SHvOtZxJqjtip8iM1J0pE0t1bh5jr+NM2FKtvvZdPuKdC538qb0xQ
xZMlNZI1kfAEoEiVigcqP59aZWqHqO1eygOV3Fag1ItKijqaZ44fykKVPFYTM0S5
80/axi3g8DVm9rFigByJg7TkWpGt2Arf8zwLwAPTEK4zURp6znvus96Ct2rhK8pp
ab4ZlEFq4JD1CTxUwDlB7jI8+9tHALczctyOjKHpG/V+T8X2G9CUbsjy67SbI25H
y0F3bmyuYYP3Oxq0jPJcgH2gpWCu57wN6FQjZfx6dW1uv6AUSQ0ztCJzapxynvJo
22A0hsuZTndPjlNPgBzF1VMKrdLwkGzmMMCUyBz2ebERZpl0SdiomK913v8Pe4c2
UJuQ8ApFHHVtfFkXCH2QZ/fd78w3KgtqUONEH5kN2ibhTb/VpnmGcXiWkkr5LuKC
O7vTlDIFErJssVwnVzTK5DoUgmEY0DYhQwNCgFHsotgAxvQqE70r6Hq3TPF0u9+l
rBSB3WHikdTE4WNUBtgh4l56OTJx4BhDawpR3FFEWF+QryEvDTSrS5oYKorGksZf
jkA+UWJ3OXfwvtv5JZ9NB8/Z8M+/AeVb7h5a1JC1+jUo0/zQJolCwqSCc04kibji
U2kCzzWzXEzivntDhIoJIePuPZtT0SrRG1MHpWLVq50BEFOJ3o1M0FaXe0P2QRVh
srEh/+SyXGf474mReRYofIGYH9AetTaymLWecmCMhm9CW98w/jD/NqKBI3TEnCQ6
9wVfKEZ0p+DrALXrMCekPsFjsYPLapP5SpZRSJov6mW8+xzSdE3mIo5BwjTsPHlP
Ue0s9kJwWH81Ab01fIixVtpeqxaKv4Tq1rQvVimUYeBkjRyMmndY7XoKK6Z4FoB2
qPT6SLmWPbLvbvDtJs27FZBsbEky3j2ovltjZzSau4u3K7OW9eedYRvfn9lMe5jE
KGLQCN4ApNvhcHrVC81xwGbEN18Nfm3CoUFfSaxEmnp/sas6DBNkmrARipz5rJoz
VuFtdOHp+WCGvOQ22GeUrYnpJgAnhiq7XuBAhZu2ohRuRmgK+xwyeR0DIcL2vvyQ
cJSOOP9jleGcLlvOgfe9Cx8sNrfWjuRVWZ4jHFj4P7uXwAul1mqwBJmKx8ViN0aQ
0m497ch6tyEMeaEAJBzGfd2BWrUvF6GrGef0KFLOz/6jjuUl+frW7xLMpp71aQ+e
Qn5RHThjzc+4x7VRT1G6ueQaWnYvTywdSW+uB7nCqPY4oRnNnkzVdsJaemXplxTT
cQop0iqeWitnq9W+5ckQgmUSIxsCixY8w/a3VahiVvMpgN/BHP/keaF9iwvkKoht
po2/PxQbHMobRtykw47gKpL6G7YSzaDLKdlRqu3EXmSHjYoHebS1A7brt/hx469G
ILFFAUS6JUHDiltFzpgigh4KSKKBOIbC/pCVoZ9Oe5f9bMt4NTeufHMzvs3fMv7o
nYgq6VWsh0LntZpvoVNBojMVnOI3mj9Ke+DbWHVoaTUIcpN39IufyouyWBcmjZkL
ho+4F0DMkLG2WKoK1URhYxkHFSqTMPDMQuIyhVgK+jJ4WBvhsjZ4bqVe63Q062eq
P8x5u6gOtGGY7bggCn6UTeVlBcttlnss+Nh8etPlnaDiCrKkOYOQC+POyym2geQj
f1LZmDiln8ZbGNd2L367eW9DUiO/3VjMQWeJ3/7w3m520kXy8HG5G4mvlbITWeU9
0ptTUkL8OGtkF0Tr6evqyr5TtMK6vDvPPxxxHp2bPP65GnqrL1nCkxNnM99EBSIf
7o8WCgEPVBY/Rw3UAscI1tTomXitz6HchQ+5iYTUl3SHW1aHefkyB4K639/9Sxpm
WOP44YXX9r6W/nAA0X5BDzhOkqqpt/Dy0x7AOhOUb/6Uw0waKVdwQGUN3kToHyz4
xno5sHYc98MHWx7Uc5Eznl+6U4f1QmGCOvIFYQqePdjIvIBzprzEEJoJd3XhCj6r
c/0UObAfI/NEPfIAFUoeZIZe7JZU7kRy12HHgKIDRaCmEE7rH21DjAckO/R4XmFD
CeR3Uwwak6YG00KgdYpdMe42yLP0gvxK+0UgcvrqbPRrD1AUOHJWpXHV5M4pjL8f
SHxP9qSuz/Fd5/k6e8wDtyBYvbMHJpIufryToBPG7s6hP4SQQ9gqJg/bdwSk0DCH
Y/9+LNclqe9SfE4tMTvxW+shHp0NA23f986cvs/N0wCX5tE5rnqFAslqWX+77Ze/
aeSTxNdnv1kzIJiqOAJjG0yvfAWuyQdLFJL19O0c2uqwYoIkWKzIZsevS8w+ljk+
rXJkDWTJRy2DR0962pRrfoYNoZdvTSvmLzcF6Xcsi13k7Fsa1NpEv6nI5Y8R/rko
Exfowe2gYOZggPO65xw6WCYBrsnJlw0DgzUXPLu8txHeDMJGFBOmmDdOOAzrP/2T
OKQdX0VBx0rMhCBI5RhPl9zNf0HqmZ6HdCHZBhUrBvPWX5XIIe389R8iK+UAxw3J
GNlHAq1r3i+9I+3rM0+0XjCjKxHWa2XR86155c9AaipFc/HFcbdtNO/oQSnRYbAp
xLbN0c8VfB8bmGR2EAnwage6baOpb7fsRPaHlO/jDrWglx2mAwuoVPaI7+ESJB9V
Wj0PS7Chp4jPLon25x2/H65hptS/JiJeip+nMSzcAT3fIFdgD4mxk7P0ltIDA4VV
bCf9tV/Vb0oEOe4QO6GZzvjNA4eitbXsfI09PaWWTrE2lWtCLlE3nE7M6gyQDYvY
UY6WuwnIXGlztPcIHIXLwinC3h3g+7ZGSYyOLgT4CppDlwVEufl+B/rwDrh7nAJM
x1ED8Me9tGTr1rm/4YLVsNJoLGnEMlKsPQbS58kCox1GVw7MBNpsGJpZdMxlJB4r
VY/9BCFsENQQcSM2KJ1O+cho5BYKvb3kT6DtPtwBy1cfJMqi12Jozch33H88tXCA
Gil7um9xYMv3x++02lYVxDk2BT4MZIQ2/WLFJhZ8orCeKpyuAq6Gd4lbdb0f08TK
GnnZpj7OBr5Mo5q7qmEv58rub8nhfWYUCp1uE/PrcaYpCKd4N+j+H39c9/+9P8A+
WKuNXbdQY3JlI0BuJ+SamOhGKOXlD87ZgpE3NsPsSb/yQZ6I9TWS6xTtrutJrpcJ
bV6lEk3Ms3kgjCE2Kf3s5dvBd6ZmkkkaYML1gOj+bfp8ehL4Ix4DFlVGv0gfDwT0
6eLLJX6q/RI5kYcy3ax/HQC0kKZzDokr1xgtymIgac+AEdtkfMf0nFOAPhhT/RYn
A4WHJz4lhzN6b3MRc4XRmrF0Www8VBRJQ+WPEDaqTs4gTr6A3+R8D0ZEcc0tkO60
FLyZaOwbaLv0XGh5ZLOVg3th2OX4s5l44hKFu7A8HBMSFsUevdtfbiwTHyE/g/z9
Pv2sj+orOKSiYjYeOomlGJoDNJ1AqR6wsUyYBr8uKKL0c15JepZNoO5fAp1Qk7wV
DwAr1S3XA5k59ZLJpAt0gnUaGYGr5rnYvlDc2pUgrjAi6iN+SmB/ENLHC9KaYW+Q
ru2V/QinsCBQyypFPhu8fi7gmoJK128WPcPnnWGH8XYHNe1sClcNp5c2thVrtxze
CcNkNNwElY7VvJgRGW7AmON36XCODA1F2EH+zlNm2J+C/l/7KVpFkYBGaRvDF+S9
8RnBLMM45U7Bd/6w0Sh5BafShzhTgswTaS6g46QuMVV2UyygKV3GlNfM0i1KgqPY
M59M9TgGSlfG9WcaLX5YdybfU8BvWUq6jpeBoahRrnxQnq3L1fKZiSfcxGhn5Rt1
yS8FacAhsLr6k6U8oQTR8Uk4Afzwxusx9cOutPxuk0eXMAmEBlPt/ljhW/Qaw2GG
kwd1puwIdJc8KpGNG0cAiuAd9hTIiCqZ6xYoWEhkled97qjFhOHAMO2WlnJfD2rh
Jt+s+eUixUqB4l4+XhlyCVN8vNHXMSePvFJWYpHmvIvY1UDQf4YHN/T5AgrzMzeV
QwZHiy+4440WgOzNdnKnqppRj0OAzUls5Vgtx8sK7/7KnEPB5OYIi2P2OqCGlqzn
V8JhDRPbLfw6gEvYZgYkmt4T/upG3++RHjXDKuGIRKv3z6GxN+BlvrRo7dw7hKDA
ofg59C+YaaulheuVusXnnimYeBqO/Rmbzz8YNqCxismhQV9oHgmkqmbAPaPhO3Nr
GgoEDNORgd6CHe7YYydKRjY/hhh7tsE7VdAmqXMu6pQ8YWF+VXDM5p3Upf0Xexk+
i8Rn77JeNSyvf2F7XoQSPIM9Y0g4f1o625WO8FlAkf6fr1NJ3/fmrhEvIL1phNS3
xx11++rudGv8u6MCChllX6e3NXYu9ewXj+6aQRIc2Gbe2bl9jDt0IWVcfMsviAoi
wkUMrw/lRCpMYW84OY7xhfoebnf8CNcV5rn1vfp0oV/GN090PYUNMpkiJ01act/R
OWH7qwalRbNilvy/VFzUn6Iyvs7sMZ/RBfCfb9Ni9ZG91P0g/HxRb2K6NXLJ517O
yxX2wzXJWk986jvRJVpc5h6B7YOJbw96kVekY5Y8vIJWtRWWrWmw+gxQ18FX7rvK
WJ2btZBsDSgHtBscoEzoSnDj1MjhPtEM3/PBQZufSokp5ecUVPeBYB2QyDA2gkU/
mInhkBtykxGilG2odQeRpw/DYGoDX+lp4eaz1BxVI1kD36/NuTS15Oc1p8ieMHCv
lgRyYoS1Sbv8v/CzONOL9v09lhrnbPDua43HPMVyZa4r5ISg/JLdQKCsIsJC0WvM
dCOB8cEiRUJ1D6FVSNkQkl7kfghUj2eNrDCJp/5xN5l9I/SYPeqQvLo8Ws2b297r
bjXa7hGX/mSEORDFJUBzwkjl4WKdArXmLOLPh/VRMjSp5s5JhYuUT8YGqF5sB5Zd
gCD4vJtFRrvupSDo+BGwRb6seyawBSCNN5RsEh2f3PGNgMekirGjBCdMi+8mVYyX
2Fg+7zebKRmiago7OEmtWPIkQctOFIarc312w1TXhoBpmmGrpDQM6RHhP+0NWtyB
Xe8xbS7su+YtBmjFPGiXeGJmhK52IRaEnrUDFqQYNjSkwzXe6N29JVKyiU7qGvKM
QcrrlQab+tFq+CWDqBdYFbWJHTUegSZI+/eThUqJ5+46BsC/GouKTJznK1J9c/CZ
dphvQIrlKMYPPw3Z2g8+uqqr7u/p3YmcSN99QOhWtOdOJ5ePXtylbkjnltc/XYm9
X/yLiw2emCrQdjj3Pcovw77lrcYzjUw2Kfm7QVpTlyrk9PMER9kVsORhFRz2V/zu
ytl0JpdiJEwKRFFS7CFtC+CjDgec5dHyj859xrbu6dcjM5fJBnakK08TKYj3zCES
xL2QGltG5ADw11JyvVnZ5s55ztHSFMgencEOuZYhodVA8pPBz+WX0GgLbVDTEBoz
/z5zOEFnv6iU6Db05QP43oir+p4D0O8A2W+WAj/oAp0V2HpKpc+LhgQh4O2U000K
egzrH2++6aLkfmhnIPjDvWku0pQdSfjTMq0OcrB2YF8gP0yp8zqEe31gz0ObNTSU
F/xBkah7TovU5LDBUomO3zL3eGijbNtTe9bZWK1iqXXbdHuzbo3WKmWuQnqdeUEn
XLj23XJuXd4rQbe4Brr4rHvFt3SUIc7ZVXSDClFtHC+NFLFFLizWWns3bIDgEJgD
q5qh/SXxlAdwSOgj/iEI0G0YUuAUzMqWZZD3yYRti3UaxrQujZdi3qaDMLXMymnY
mSGTei8JR3pdhxC1KhS3fnCWoRQegO8FYDKCXOzmNBDxN01UrhZy/RQxtLzy/WSZ
j66GzDuIK+M8yt7OMsVsZlLBwbY09ZVfpiAkxIuc6VjO8R/CNgMypeBXQfoBGyNf
+2vUv7cPCiCD7QHzNEReZjQT/uEuVnjQe+TC70u3gwVMF0U3YI0m/iJBTahEUlTu
5MTPjZXtsbzY0SSsfcQ6Jf4zKjRBlExeZBOYcjI7UEoCYQfjW+isW3qGu6/7+H8P
8gzBjZKTwyx71tYSI9weSMxfRS7LJtnWdp6yeSOIxHS5zrUZqyPOEPnvLurYlEgC
JObWVY3jLTsQY2iU6B0r84qbYY1c/QxEYKvx0V4LEcr7EVnsP+cQ8kqexXVi8pB7
cYbuq2A3gn7ZXs0vgOMLb6nZt4CTOD0f7s2vvgzieTUK4xK8sENuYQ2OqKmCtOoS
7Mn/pFLxT25X+xbJvGGAJTCqyKVMZ+3om1b3bBpy5TeCHoiZ6QA+HoRb+DOST6KB
gsoMV5IIEV+RiZ92nlNcBgaDWNbSTK0uSHyNkP688mmm2XCq+rqRHdNjTX+7yZ64
+km/tQSLmXg+tNc2hAmNYHeWvNoAESMR0lucLr07fqCRUeudoYhmeaz3JOsjjLPf
Xex9hIo1ZdQXzh8sM/JhIz8SJrBIyR4BaTz9stUsKr8+AMsjtZwA3wjldwsuvK/i
m6/NAZ2kOy0mKoll2aoL5xVaTzo5/cYIc6KfNuuQw2dh5vgTFA0Jnx4uARrMumao
P8fHkx9Hs6jd+Pt+xIH1i8PM+8nQAtCD25p338aVhqNlQI6SyiyXHF0i7Kn+0hNd
77oYjJ3J4ZDg2aOKEQikbmm0VtdtVNGmHu+DkQkuoXv5X/7Xr94vIg8qWtKEzXOT
leUX2AGfF07mr1NNVisdsQ/p/hPTD8zIWiOWLnEk2YtInetG//oiApq181/zweUM
NSBqgpnWRaztWKDQryvA0Hs+K/MCcHfa5+j6oWlsLJce+Tvck9y5pKrbP92wB7HU
dlLwg74tbW3oWkoIrPhKeMzYqLU4dl3jWX2PLInEmeEK5OELkguPqTmliCuI+gqw
Vw2LZ0o/3+3VH8Zwh59c28iaSSLLH/2DCDNE6G13lJMb7c64c1vJrYwGOfYntT+H
vcdF/ZFv2N1UAU+9V0czGMNbz7oKEIZH2hggW/NGqkq7giYEUkA/cATWIKzHV/iW
xpPuhK7e8MD5cWGQzHAI0sXHcj3HpgGFij+JvLxLrnFaig3IhB0cKXZ68YFex554
GU50wOvtzSUuPXC5hAE3G/Jum6TTrhdSEi/GDlyjyNoxvCnTE92rZu/LKxgICaPl
DeRYYf/7n58lVYdo/ybh1wW1RhMHf6Di4ff6jk8S0763X60NcicmUeGnv6ozGfX8
XyGYpQaD0gOirveBAxR/KNH81TQZNXm7zc5gCSG4CW2f+GS0nwRjF7SAPagXeeRp
J2Uw8mr1WfEpsfD1S99ibV3r/8futzM5WBmW5AcFapMnzFoUknurkKZJCAJZCNtW
EdGcl+M1kMLTOBzLQLAq+jB1lQCYlvkFIswHrx7YnlfA1tL5x8kqfmW3bbKTS32O
nqJakx6koTDcQtUWszkfA374kzGFBiRKko1hGojpmHQkdmFa9uDIIDhGsVCW3dtI
38eZ6/HbV5qBgUvdZohlVExKawBz0fxiKtdeoTPDdJD/rMZlBEPLUpnkVkiAIhoK
Oisuc/Yla28Bw5C1okc8rReCzPBcggT6h7breviQUvui7Ke+QwgLX3dk27zR1s+M
WinNen2E4zZFjD2JQUXhv2DaesChCOHH9BvDRAsxNpmyOt4YyrIKpoSyLUR60y0W
6MEJUl6LUfU2uNtoALVdamvzT+xNxkGe6E/hijW9oLF1RE0Fj3ISN9+5XFK6d+RA
4/vIx8vdNTkl42HYZEkGyuOcIDijyof1Of2l6QoUiFogYP7OQF1R38l+PnNgGwrs
cGaxoAgkOVr3Tt3bZJiNJGXuOFj27QJbLtsNPCM4WelhSwHkym+rzot5MGllS174
O88S3S9j45OqYV06uVHW0Gy9fGh4Otv2deYJxS6UWMy2TA+rCmYQl81cebOBPjVM
ffKpSUDhIP16f6MGQFcWAYsZxApvbqVV49C0euG70OfmEhg2pMOUV3OSAxRa+HD9
IPtx91tm2i9+b5v2IJM6kVKei+RU1zIAxpAnsxN9wY75Nvti165jzLHdNeokaRr0
bUNc7KX3JviTep7xkZitgUjmxpSoKpG/uaFhlOPQNT1qC3qD1JccpmZyzxy0DtuG
ZpkFB9qhwHwGnm/Wwb08wIEkuFp+3ksG72P4otBpJ7a1NWrJAuXuZFRpfTKVyx7W
6rZUhvlGnMekpkNu4bbKtAOKJF5LXxCLdoo4U8/rneIdqnwF1uYk4NZTL0aH/uP4
Y2dqEpIeihapOmEdf6lZDUjWJEAJFyrEZKRDgma17t6Ky3IoZI4hZXchZziMk8d4
3/tiEvhFD7i9EwPymzP0GC047+EJJGqMvYO1z0nZappswYAuuuL8B3ugJPN89EKK
2NfrDQRprjQhGqe7NgRkSWva3guzEFM3MI2lMKzJqijAMB4nl4aOEZIcigH/iZjE
0cJeIa9vexqESUwNHKG9nV8SisW7lekxcqhivehnEHTC77vvJY23BgfQWVjExnWN
CQqDImYj843AUBxxxfHvflAd/3OoGo7IS9/pA8OB2EPUe7EN2WdAMJRWo8gf9mmm
IxdOMyRaFP6jQTRuVtpwvwI2OymeC580R+3flJtFTwYjNAKQOoXPNS4TCymaC8SP
8taOhh3vp6BoOh+peEyuB7yiTQiFbJ36HvU/5rpS/2X8zOgdE0E+ExCs9fWjqCfT
jPCytdj9UXePt456QGvocT+hzW2pDUGjC96j8Luucut7fQAt3zW8jVmbnsA47hZO
d+ytdbWn6D9Mg4zejQx87b9JfClI8STJhFoq9+DXNDmCCtETm/fhdgkdajX4upai
YHqvcHv0CueDmVeerc+RqQ7NMw9BVznzJyWxsKAceMWazrxppPqlyeSMFzc2Ru6f
k0XFMIf+lbEsJCTaP6olbaQaGM6Jh6qaNQleJz+FKLY0pIzUG+XB0I0B5XoT5LvR
yr/0IWdYwRqN1JrY9jpP06TdeDy+9W5UbNW+ZfWJ/PCRK8LtUt5QlqYEAjY3pjny
BrfeYF+kJuEeHauq/uFdHpPVm5AfJEB6E2qCRZu/PBTwoU5nuZAVSuHiNG5VBqjA
W0YOLZBv7UIOucEq8B8rnxePKjgOtBShplMoM3YkSHOyRKyZ8+8nR87cmHQogA04
h6iAJfl+qDuq/Ad1OQbdUhLsTxR5CT8evFzgWH9lp0pT9gmeFpYtl5hFFjh+vMAm
o2aeA9hbEjDKcMUU8WN6K4hPSnNb8BybsUWCAMHSUcTFuxPYAxAwfifcwGErb6FP
FOymdiHR1Du4FYG3vJJb/qITQaQ6JsLPguG2JDBBhZb66qDCL14qilmp/3vUaPZl
ccYMqJ/gRqlNCa6djmIFdkGphDtyp3weFSLlsOolkI9fUO43PAU4QieEzaGmEwJF
HD2RMc/9K2GOdP+7D3/2qhEiADSwpSt1hQjMcoZBx0Zx5w/k7OrC4Cy4EvFM79Ca
4ChMmqSEusVG5ZKcDOMAXSvSVYiBzXLv6MF6sayuC5MFi9iA1tAYXREufKpop7aL
JeRZLp4iNfwMlYwLzukvla8jtrYMn5FPABpNYM7crOz0ggh5dMqtYavl7OjfcoyM
Y3IYwUx88j1XOzxAigZCejT/OUldQBHz1n/VlfhsCDNwobmkxO3SvrxrTV1xlNjk
ObhpZBJdV4mrmflLExgE3LFIQCDg7/Ghizv6w82PbTLjuHikfOxGBKf2/nppWQcf
8Xt+jS2OHnM7VvDoOOQBSqZVqI9dJ6tZ8PMpPlJYu+C/VHx2aKotl2e6bVNuoPLf
6tpDm1OrhZ+SVTGPYwcNqQLUcTtJkfQMOnM2zXkdqGtO6c84MfXaZFDsP8wrEaUO
QelKkA410GMAWxnhjJCDim7wjg4NxjSMu+CAFn5BuaIZu/hFBNvR+vO8AcG8W+Bx
3JTwHc7t8z5szszbSrXxFpDMf5lGQs+8U/P/sXrzBs+zg7Yr5DetpfmkpJ8Mp2GA
UqjT51Djsidsc+p+cQkVCD/GWq/pycCmqni/EPX5LJXwygdBPR/3/GfVvYJ8NZGe
wk5kTJaxNh/tPz0QD+EsgDAEIXzwYLAwg/WrOP9rwzZQKKt4vZlNYy/W94dh95Q6
5XWh6hvY/k6z4eYP5Zz3XFjBaiLIBbvUSwmyqoldEd1MahmUZkSfhgNXbJtOxdLE
oO3rZ2Jt98V6zV18Y1l4S3U183V9fjETBLXhXSM2v9FJtfLF/hADmgqoAB3ZV+l/
c9EzR0aXKo6CMfsV3UVJsK8Cyl6uvd072hUg+p7oLWgDT965bjVtNPfNFVyM4AaD
oEgAcg0/EIL+3xPbPwzKLBtlq4iQ61Be4pRht6jqTwNzoggiydlZzWqOEImxvMxx
oldqhbFeupc4AuZ0nVIbzcA4xbOrEUNuva7sCuNLcdPfxFVLyJawcrGHOahneA6S
HNXYLKDJvhYmCVdTpiknaTW0ojXz4m7KlazvJzrrWjMLqBjGalTKSTuJVU71eOxA
CMTyhh3WURP3IjcAz1k2+QivURVrK42JtQlAYBQB5cmoc2bijZb9lUhm4AkDHvCf
ykdttAwNWJl8QhgLzYr19MuiHi9WuN8JYF8vZNfJzWUmYNHsiS2TMU+iIHbK0aQb
wi8QUJaP2dhTcOFctzOHvsMsKmyPmMw7K1NxjSeVmY4aSzwYcE1tKTBxpIPzoBtj
4ijXMTSu7fgQgdODLf3q+9GV7RZu6Ae51yWuhpm/ksOWuZzaP+ZQO/pQjImTKhIX
JOJuX2TzE8IHJneCbEHupm4xiM27wG0E2JfqlnQqdPfWRYbob7oMZINNqtH6QvMU
XfJ5jT7IEcnTPA086ntbF3qEAONmkAttKJ3gkMihfC/Tn+coUWlRBNjxDrtLQ8gM
lpVY/BjOqZrICu3KzHCUq8pkjetz/rBESVLG8OOTdGxZDdJ7I+Z6nENkibCjaa/m
yFpxiJH7Yoy2ZCrDkXS9P2uQLNPAd4XRdAS3mQvHAheGJaREjBmxX4LFYnBeGtZY
LR0V8Q7SOJt7w3tLsbMgnVWvatb61B28jTrWJjqlK4M2dPjmXrOT7NCqm1RYD8ud
KYrUL3EH0L6mP/uZnfvxSFAYNxmrekTkDwtnZP2HAxU4mrGJnI+BBAnIkjf58phY
1CpYMNmkrN3joeYb9K3U7atn3+5Mkdx4O44QGZw/jToQIpfAHbDJHXj2He7TE1gU
wyS1hPs7vklT1ca6vH6e9W/DmeQ49tphYZvE1933VCo/TXJ8AA4DFfR4Sj8rqMn5
I2LmQcV+sm+D98smhSy16yNCT5xhKVK8G9U/AE/Lo+a+QnEA2D34WgqlbPh7oskY
vkLV3LxWY+GwwmAVhoFnBb7V0Hy9ArXqKYNesW8W8krjd38pJ7BO7dGs+k9SHZyl
IDMx20giVwEkzGSpN0ge4gzccDn8DyBdC6D29CjHcfhu5zWnBcm4+V7tAmZCX47M
zopxE/2JLh88joY1fy8KWzNepjZAWG7vHx1qDHks5Bo4NpoSIgK0TvLvHk/JMZDF
RSvg7EnXRefOhJuMwqGnlfEMUKm35HXmPTLGa52EvOMGDdkiFIz90ol4+zVBaa5I
MwHgblIMGJzDc+gjCpDFv06ehUvNFK2uEtTtyh01aectUHkBWnAJ3I6CKV9Wo7QJ
9XnRayWSpUqs1mSHfty9ieqdCqWj3MbDWyxlCiUnvIa5MpnnsBI+8hwpdYmkIPRb
laKbuyOvQYZdA7ae3gA+6iYRVtP9xPrZoKxKiXgHMAeIMSCvx6Ncy28P/taXEnbm
H0XR3Zf5PkcD9iW1p/GBIpSHHRNyLrIz0u3sMFQbyPTzgHR6AxEnmSgFDM3bMLQM
mrOvVBufcVTepOzzfsIUQmliNnasMeVegVoxdj6VfpGnq2vm562ylOnooyZchPk5
EcfE3HiqwD8PiNX906pMHXdH+72I2qM/s79oQbfhpBzTGORApDigSdqShn65C9Ga
24FY5UKTFsrE8sI2udW/J6n9pEscwR31w11soPdS9zEkfeP+sks7+ILh9BD1cpcV
OLON95tzbJ2nT7jO+y2FqVRbk7Q33WFy+gWw1TThNAu/TQk7Uh0OCgQ1xGuBC6UU
n+jDoXe5uN4wwgugrs68IfG1RbkreGaQtrcx5snLMl7KS6cTnqj2JjSRjbZ75ZFO
Xfv+WoWIhG+pLKcYZ1D/pdWF31CI1TubnfVWj9R1VFlZVdKvH0k6fYI1LliXm5wC
hOx2sYBkAOlP5CZLxmYJ6nHvrRQuDSOokSzCO+LbV6ASqxEohqUlgwoibyzj0KHr
bsXyuMlklkEpZDRDGqSx2sFsp9tLEidrRxj07OcJCylmzHrKlT3U+40+FhpVYANl
PepZNUc4gfs2AiEBFlxUA1v+aXPG1g7jfB1OtdBo2AXbEUD2XyqmrJwXLMY0X48z
vEea+TUtS7nzgoAyz+KLaulzVsHy/n/1tml/I5R1aim2PUDgvsuOhSs/rYeOu9xZ
hUrx/gj5FeMRCMtiL/MGeDXWeHNDpqehatYPzN4NvMc5+BtJyTNNGBz0G7flZNSV
zVd0MK4xdpNviddBL8Ci60EXg5Udz4JlVuEmgb6qHjeU7uUtztOTuTWDtAGYl287
/aTDwBbjB8ybmDe3KYUO5nh1rVjPeXOm9HmwEZASw1r4He0zufkk7ruwmjLxdNQK
7Y3p2mgp5YR6ENScw+gVkAGKqvqGHsShixQY053npNgQBR0USrRopqrCXN3jt3K2
PLYVgsRFw/V1EBqEnd6HtRav2NJNH0OD/VkhIdDlUx5AB/0+lNoQ7bHZxsJmQ9Lg
6k8hd0jTsKiSi4WVHflxJy1yWqWKXq9xnDFZ6i6ghpgpdLw7IANMM+narsy0V1oh
37u0PxdY91ut/yt4P6TdrITYuPfrcB/1hpWaZYKQJx+hx/bKt6VrbsUuxviwNUE/
bL0nVXDaJzhytjb7s653jHz0MR7Aym36mM1k8pd+Cq3SdCDjOd/2a55V0mp/DpZ0
1fvAE/5Rx5I6CkyUxS7Ng3t0T8osjqwGm/3kaEtuONozlM2EqQz37GVKsMjS7oPg
7PBhYoREi/Vwl8tThkcTJjyE2AyeDVprug4Ya9e6POl9fCLf8hbkleN0GYGfBjUS
ACixgwIVoa6tJkUTYLyfcQqEf0/gzbpWlEjSOrplj2FeHoyn4DtHXHWBnbqeVukn
Hfs9wxUFejkET7qKTdVeZQ6aaJNMR67JNGRJm4A2Wt8E3sIMF6gMRR4S3oT4CkCT
3eFcuq26yj/1ifPuTY2Rqp8wpGhFMgUAtX9QtnQjrHOIsRW2wTcRDh2Iqu0yc5aG
yLKANMCZBP+TZVXC5NsCZfGBvhn5R2A/ra3hvGglcDxkiqrNIaJ6A6hTlwk4hriR
Na1ReRFNLtGYjzGSHczpM6DPAa7r38HSE6aCOMcCYcus+1BPd5iDjaT5eGcZLxwX
B/bhNA5n9GCLO4iJe3CQ4MHFxjtwvpIwVNLrPLMavuUliTef3i0g4+Z3kyBJ0iHU
cIFrrq2nmnBERrsW+7pE2ctQLWoPdXaveNpPiE4FZsQU9SNzfaEc1AmX+Nk2aq9Y
PSLfivqpiDU8D+e/KiTkIiSTNbrYcRVkmr80dOXuvQ9qj/KtljpU/AXCY2Azk51B
1Bg/ckIZuxP6us6aoLrERuh4CDpsu12ROfYhvNmhg/4sQ0fTyeh/H+GaSIjOPGKF
chFRf18x1nmVxjuoNGObvc7qeWrxfnwXHFweEZ7fnYUuP5HWQsEJxmhzRt0aFH5o
7AUxhJBW9YG6XE/jhHVlG+rt8ke3aCbxyeX4Pwe4E638TVdy7QwQyoIchbxnytyx
tZvwirKy2Yd5giclPuHezRe0qRg5a7e9K2EAgSG95h1JzYtSeqBVNwZlJ++5JwuI
nswrta7vhExzsT85jPbvVN0K8NWpiJdZw7gkPzrnQkGmegqwdf5NTgvNQwVVx3Sc
ac1wQvLO1f0YG4qH6ZqYci83YLxfoo1RsWkFm2MFwcst3OBniJttShfD2ssDHNuK
xKmOR5SEzc0AExQ2AO41ZK6jOn0qxDRBEzJgUyJQM/Yv0PwF5SDJKGlO9BjWGXwi
LfcTSAJ0hHGABrAF3r3ZW0ROgYDkFFfxeJAR1OjwSiYOjTglSz3g+XbU5tVEJbC6
DLEGJmggEOSFQxSpqcdFrDx/bcb7mMe/E32H0d4d2rmHSiWyUvKu0UBAgGk0ybjO
D4r+1PiI/fgwlbbaiBktBes418RJytzHLYRN7US/jzsgBaC141Fg/cnmbshDD97m
X+XlQCp1ygsW8/GAJd2F5arIB+e4wahvplOXQj3kHRngTGh7wF262U8RbT15Bqb2
4Rke79TUYVZeH9Y0hdwnnDVgLqdqoL9k6oGmtIak/EKmZSNpwiLgaxx9PjVlffi4
l2wF9S6sulDJKM5aZWIezAIh2gqSdRXp2IdqQnvPPPgmWyatdFnZT/3PHRZ8W1Pf
A4Dxoh4wQitws7wXH8FRroHxxRY7S02XnPgMTKfRdXGeolHsjXBrx0uyKJdr833i
PSvzMf8X+uONRmotUi1ZT9xhPf8KndDA6oKu0XKtckRhgUF5IIXwPF4kYCA1slas
jgLbIPBTSyqeKFO/RYs3IT4JP0m0vB+evIsGQWng1ktu4p88w9K98riCgWtFBQv9
Y2JIb4tZbUvBd5Kb2pNy5kEJjAUkp/X4ROqi9011MtwfgYk7WyrVpTwZIN81DrZl
+s5G5LX2+isFYnLuuNnrTF/AmhlnxdIycyqcT97yfrNx2LL/25+qzjI7ph6Z8utI
A33dFOtRVwftDu/sLEwsWrXDmk5g1GFdXEgkD9WRzPepjKEJSgg1EBa7Wyw0HZLX
ZP2ovDcnDdweXGoovG/rpeEiqrSeHmXZd4Nsd08ISAlZiaP61BNQrtrSLYmM350j
KnQugB6t0VOEW2urYe0Uam9irVAKH/uUsPj/mCBs0fMBIq3nQKGFi8pKnFNuSUjt
ml9nipY+x6eXF+xjXAWRZd1TFYCFaMJ9lvcCzl2Fqc3xCKVxiZ32coLdcOgkPsjk
9j5mCtSGoFRUBKfXlGqcLWFi/0nA0F05+kKZoSqdUHFsGqTBhQkLRc9b3lFJElLL
+6ghOg7ToFmjgGwqLP8skxLiIb8LO4by8U/FEGsTvmd/yYBVZWDmAizG3FK86RNc
ShgyAFmq/pJILW5jNuOfGey2YVcKJ0Zt3b/X6vrSsM1GOqRuVbF5GcxLy92VtZwB
/GUDYH/PuHtpncbYHKgROfbS6YkoPDt+G7eW5cpECoR42BvURhUeVauL8swQrrLM
UYGNTKdGKOMhBYPHE3AKucRW3yDTvPWeuHZ/9p+Rqt1sS6f/+0y1YJO9Qno5n8Mq
EvFZkpDCI9gmPudOJGk2zxeSCdmsDuwJ+Nr2NiudkJQ6CylOqfnZV9nqvF+33LJW
QgcJnVU38aRTp4bqPlrvr70BoIfKRxmTgKSKEzzIUhwPwlik9GA1pQCduzEXrXOX
hPqJHycICTHbQgHnweQeQXbJIkGpqE8tP/0lJyLF3B3R7D4uQ5OUclJaAuY05LCR
NlmIZua1pJxliaswHkxcAGFqMSbdwZsL/dR2GlGwKwLjlW91C6LTkLpHiBe4jPsr
EGJyKVGry5gO2ymNL0IGU+7iQrBLOqFNL2aWZAc4u+a+pRNx7lNIaMWBK7yRZ2gq
Xwpw+YdRy1tZkn0UDefnyCJhSPZWU7yM2A9yKpkVcFXhvOSNrbDgi7Gb4jFn/BYW
ktZ7n+8/IqeC61Qu8FlovM8vbw5pwrLKWrYjh1EwDcFbhMSzXEgXp/JLLFDKawgJ
TDwpm4FPasIJ+KtjoF19K1+SYSNPpUwoFiiF0gwkVePTSwRjlb+BABFqeCJPRfVz
CXlHwz1UY0qH3VuY7Q//1lVSwg0BCAPGeGjreU9smGhjFp45k43Wc8g9BQWp65B/
O7veiknkEgr1h3LiqJEg51Nr/q2g1dicBttxq6aOBmh1mpHpvHihAUjrx4jsX8VQ
I5ephUmAWDcTHM63oe6mURXLwoP1nAzNGUWo/5F7Fgz1StOtcHIgB2Nu0EafCoJK
MjAttQ3RqYC/GkZheF0UO+eAgdxkss9SHhlWdWKx2GV8835J/vOfXRjcPea0+x4m
mkga+gUf5NXLUfQesTJZcAPcrafK2N9O9Z20PYqMnEDZVpAN83yDKRkneE4HpeE0
RoRS559DM6VIxwF/jiNkuqKqgvO3o0u2KlC/Gw0T+eYvuvBKPvlgXV0Dtol2FsHl
azW2Q5XdX+gmTesZdtngBRH5qQyHnx0FZyKCTmu3fdekBUofvAOeiR4b5ZPaJHv0
mlQP8+PqSWlLxTe4FvzBT7WdN+XWZ7CrgxTAS6hmsNaAA4NribXXs1B982ilrgL0
Z8MZ9s6ecdEtmN3hxEBUCFB0D+MxoPkIHmWlo+LEFakth5t4ISG6CiHA4+2r1Ly3
rXPvbLkVsQQ3JN9T1Frxe6/PhyOpRWMDN3+TrPgRPOdYXoXoukn/mzmOdWBupLhl
zalYY34m0LC1i0A+obVUjHuT/KfyH6Zu96qgXAls2xPlIOaHuQ7p3p0pte+EKfFF
eP2RBfNKQj9qJfr+mjlwJeRrp9dPyA1eOrtZ5QSYE4pfW+/Cbn1Dv+wU7wLlAV+0
M1sXADNPAJxPA2ErqJp1kan6Zt+EhzsgjRatXFnnK7lzG4p2lVs/aKvzhE+9nO2+
CnnZIXIyHP0DfnoUSX31TlASPMu0uG+08nJs/2kYRXUP2xDw1Wb7OeNzF8fWsRgw
odEJaboB42vfxa3a7OTWZGY+Y4d49+mLUZF0ehtTYX3/cvGZDf5AGqyvanajNr2V
beZMNJYfynUBNwHaGQqpGS/xXUSIRdbfxwodRI/ezqcpNWE+sLIxFulCdHMnveVD
SAegR5+TAK1qx8+KukSmEe0tnDpg8CG/CepyWGMOruIMi6KpAHV1MMSVi0kYPYrv
bWbS8nEaNcLUdqI6XEXDhkPANqGwJre/JPaw8VgxtEob8IG97nBNvumwLFc90FYL
GqShQ7lm3o5RvNxZNG8cCxP8/RWXKvo8UFBl0fn514q1GVj6lzI/Zr8WDO+CyVDo
0ZF6MFDEkhBON7W6a+vXY2SZpfI58A3kd+Sp1BOLabgdW+uKWi50on/CA52mexZM
jrb0NNStvitkKYFQ5yUz7Xp8L5RdFjzzFEXiCQYaTJKiCKqkDgW5ENsOZJ6ImTQi
7SJm+P/sHsNyUFnwtD+QkaLHteJtB+tdXY/ltqoJO8vuhw+7fFSVz8atZKGzg7NH
/iVWkTiUydlzzCloeCqttrwtPECxXM+A5Ch/2nOnAkGDLnAIiZXQPZyuVwZp7D2w
he72kCxANGynu9U+byCHm9JxH0I+SnwSSWv7PpSocEVKp4strV5TMOCPQ9j3Rrvf
PZflONgBBK/wL6uL6takyEWUB/A53pAZB0gq96BdhEiHlCo7F8iScWud92sfYgzX
44Vs6WWw+RUytRo+/cvOQ7x1gsaK0k2ujJnF+Ep9zoMNGqUM6CUAozFkOqLZUOgU
ZkqS85F2DQrMfs+JR11g5LenxuMhTww+J22X936ITF/n2A58+9esp7BtmH29MliA
u86RnI+2v0esCG1PWedj5utcWJrTiDnWM0LhWer/KlYSdsgs55aQUQPfDmsw9ve6
n/zf23n/0++dyAszBqa4MSjDdAxjASTZkbUemYjO70ket9JMx6IjERc2n4EyKXTx
ZndZT8SH6PwuBInoYV+MkV3D/QR79KQesiFRx9BVD1S6CBlY0xMgPsr5bCwvharm
6zXyili7IwyxJM48HtvqZjl+uUHHrV3xLNB1FLBtnXnwcQ/FYmRTbW2lVWGB1P4F
lsjLvaa1Ncedv5VFnADwWr7O+PNPaDS7adT1mlGwnlJ1HBB8ZnU83KCOtMGgIuxr
06Jp119T0zxilUWbhUx5ckW1O06QO7QBFeTdorImHqh8A4780s7WjNVehOEPh3h2
uu3LBqwrFAObZlWoeha+nkjmSXoE6enDbos7gQjnd8Ly8AGnR/sbMwoPBU8lQrh1
41HetoMJl9sqVHaPgnv6aF9EhuODMhy+3rW8VSIQcDk1QhjdZP4wqNdghVbyqCmv
LCnr3V4H3qEH6UPWNALo2d+4/o+QfJnoLwANh3cqTNmlF49TY215Ozd7DObrouk3
gAfjoAEzjStvyVCXn+zGKkOWLto/Bo+SLhGqfKWuCzMRMeJiWhH4PZCaARruL7EC
xA09CkQSobQYhRS5AlYDX2ZytVyAGiK9OleZIWXtA47xJz1PDIaMbRl061jCyGOE
NTjj5SZOWl4Lqzt5ERROWKD1T/0f3px9z2G7bqLJkuLktxDs1rJhufyquhJXtpj8
MD+ss8/xU9pbpteu2fylbPoQBgBDrZopB33F+vZoYoixC9fTsnhei2hkrlKq83WZ
p+enVc1jGtQQ5wAjEWaVsps8AjAYA0Xv1xtV6A3QKMV/WwDlyPJd0QYzP1tDI5y1
F7OEw0gqOkjxQUbYMmP32xDWGwftJV1DDU8mrcjDdxSHueKE/RZdmMPjbGAK3euN
n+aJkQDVGDTVcJ6d4y3GiMdMePDhDmedgZ+Jx+BaqVVuZDwefbR+cXOB34grUZPU
gXLGfesBs4pzRwPoaXUhbnQ0HkrMP1C2o+t7Sq5I38O2tj6o9pwbNzAojZcrFqMp
sQYKIlq3no7eP03YyclDrp9htzSgA5WMhMQP2RMo63oo8jucQsMRFMBl2hs+1UaW
2QaGwk0rjoiYhQfxqmGV7Xvll5ed4nFCWoCKExR1TZvOcXW0x+y4If9YJ/fTta2D
Rd/LJl+XyPAzvrrcoNV1yfizq1oGWjmmnzOOgLJ2qri5MYDkrC2yR8jppEMgDTA7
mWNlzthTQ+W7bIOZoO0RHmRZMvLxfngGV7UZyuMTHLEDo9jKhfBtiZQHXpCeUd0J
uHBF/k1x3Mjyl/ZYEah8e26ldda2R0HbyeNgY7a4o85psTMMh7eJtQvDAdQFEr/x
sjShzjDADZGAVxIJ66O86Tny4OrH8AgvDytcvZjEXUQnwFTdwwGiMpoXkwRmL5zX
mY5w/VfWIJJB0BypTawTazYGYYc9RephGRp2KP5HFNIM8SK9c02580zyfZvtr53S
KIgMtCqDGLsVJXgZK51UohChXgPZ1EBimVNW/CG9iSn9Wp/N8JFE8C0gmwjoZCuu
NlwAMYL0pIFr+2eoDwocs/bSBu1Gyqrq7MS0Qp0T5NfYfMkkzoWXRVvRS/Fr+9rP
Tio2UaXtvyr5rQC5ujv3KuKHRLaPXEDSvDE1B7BSgA1hAkTS+P4fJNUMuIxD1ifG
ub0YRplFHD/gTmSTY969LkTAZGDNkMLLLrNJ36afs+vd05J9nXwqdUIHrLEJPyNo
p/5DP5JbQQd81Q00gOTAJA7VSv5n7u0lIZFGwXLfhNOjW+4BukxDkoaO8WnQ4m+z
p8F8NCRwePPzx0u5ZZ1V5XCx0gjBiiMNYnCtnU6FLlJffDYAdayRJuhRU90bXr7E
Yxuz32B9t1hghlHO6oPRNxABWFwb08dAqRkA+3Tc0LW58X5kK5GE/aFBVA1Ybfet
pNSKajZ05z2+FOiEt4/+78PZq9nF7qfJ0NMxxPp9gNKSNK7TQFGee4JfuszOVRgh
D65CyhVq13XB2OPCe4pkGuLuD+mdxQqWJizd3vpNXp4SDZ3qFLOA5iuO3bei8dkI
U53cTKUt5qv6fl88zoJH5zQLjXlwjiimqlEp/+NIXkd7uMh4dWD68shtqxRGrZVh
tn9PAUFGP4vbN8hafHToQHlothzLkY4AS+xXjU7x4MtH5ZjQVT85PFZB7KuVwRlm
bWLQ9IfSPMbDpGmIo+N6ei0vQL3/gccv2S6XzFSyVCXEDhTTB+oT6DN7m4oPjqV0
nSZBnhn91KsAGqQ7OcCgneBLh8d4GSg88eOgdSjxgegFSXeAS/C8D4dRd2YPbggi
GHwrdNWFDgvIoQN4a8WRa6hZUfYC45iCJvhFcqhoPT+uefLf56oDbwwwrrO/ft7m
dEaCo4fW582+0B6wfl+gq8NQKNlL31TI1E+pYoNu5kJpYLR5w8pLAWiYqPuaQWw7
8jeR5ahGYHOY7dtzIbQ31E0Qvj3ZymeeWmdBCRrqvybUeXx09wp1YTMfumxB1AVB
aDTHAe43mRTuwxV57MWN+mX5uC0ZkFmmNpb2y+atacvbhywrm7ub00nYcQr/1kZd
Q5ZZpfBpYm99G6dhZjdDgtYqOUVGLPOndiiMXZqLhQN/a2E8rSCTWS58DtvjvSai
X1iJAEOqIM3qySZguJNg+OHA8KLGbP/CAkpGjvD8d14Hg9qbU5HiMzS4Q4PDdCOy
OvYChCT0H9gXpyn6NpIQTUZ1AQQsso6JCv/SNFb/RlRvFdZ8jcL1D01/Sfgj8YXY
4Z6RIYCdKC/QdQMKArzCA8NzRsE/LdiX2E4ZUrRhs2MrrdC854UXVpLd594hMk00
oQDzQy6f4GIC+kBufM8YZXQ03Oym9fYDgfzkJi77nSxqueIIpu14RIelWkuPpQKy
slygeim5aJqFdXUrNtUFMxqGwQM34/hUsd5J9XA3S9jigJDaw6PdodQYy4VVSW0E
QsAMhqS5+Goqo567g91T7PCtPg1ya4VO2zwRqES4GjUJCXRpjSMgBZOJIVTlTU3r
lYeZdux4+X42DbfsVamy1/dhxEsVID0vL+QyxHOqbU+G8nsnEjLbYQn8yPcz8RWq
X4PzIw0DcDJOfsyV+kS3pswEAUwL0y90bWdoW9NDVaC7HXrqr6lINRdC1QqBFf1y
J/HUzd/mDCm19dn2camlP/7jsWI25eCYvUm1XrpwZNPoQfjDSNlq+5wNyFpYpRbA
NMbUHrQYJPdpjQMfxMaJdCgbFhCv5yJaCJA+JMzPCVmrEhg+wWDSb+bleFYWUrlO
SZr5sKH9UB0gcevxh5f9xQIURYqm0ZTLJPzW0JpgoGF4EYnLWhfMQ4xGDNaiHFX1
v46bEVJY8KoyzPH4p+A1PBHKbu7eO7NFnqwXF6E9WB/WVn+vkmNlJHVT878Wr50g
nOOK049I6bLtI+vcb0FYbwx0wwMmIvx3nTINgMgb9Cs3KZRytJx+XdI68dn1aM/N
06uafTdoDBv2V+wrx223/TsLhsnOi3SK6qw4pFUhIXZ00eITjPIvql/62QdiJGRa
RVSB1rC82w38uwcISSeTVg6BUKsrPsz8a3V8AYlZsU+4RnGlGifTMhCcxB/kEg0Q
zSIpQMDT4tb83Z9ml/FfP5HvKQBmQ9rNmFec7/RIZvRFz91i5a4ASAhdSuaUEoSh
yTlgZ/nWcw55oJ1G3vwAhxeVLg358UCBB5aPAD+tt3a849igdyP9JoJU33F6+U6r
T82P6p4wXepWbbn0hLIrdkmnMf+AStzrUdnEKoqJ4vK6cCVCCXPWNxR7ELYZxteg
XSIU+6N8CwolXu0Oy4OXQeabYmoRlthYxOrIYcWb9VGTwdLqmkQXjWGDm/6EAPkT
siY3R4ZHpox6u2UpG9E3BZrTKYUiL0ufTeEXRDSFflCLGdF9wZueeYZnX8y1XNRo
PJDGifCuaOPfhc5Pfr/g5RazKzQEHH8+ihdfXaSbGjjxEu0HIXHbNrodC81dCgGu
LvsVieioh6zxhkzlvf+/OVLtsYtToOWQjOaF2beH2IlxGgZVBLC3TrZyOa70eGJt
Qu/VbNr1JANbtGYUKEqAobjQ8FT59j7zJDLBL3x7cGT6Z79+r+MuujlCMkbNBX5J
euf7Q2rM5hELCwLaRb5HPhfKEEUWQo5ZV0gmjsyM0lM5+YFb9MbkIvSqphZB1QZs
psDL1Jdc3ibC5jj8megSG0ZrXO/yq4OXD7kg800OH/3zpmOKOIST0041IKTQToTs
W1l6GEVhrRUIAoiPbVnQqWQUBHWx18Drit06TeQdJVkDXQOZXfAe/jiY3+1nRRYl
hAwTnfj5VAjj82MwqC/W4V2C3bix6Y1cRUmAGrd5P8wFz+Sd5uj9x/mwW1nY/IDw
mLgYoJekytD8pgvG425jfs+Oqq9NfhtE+cH+qeSrX+573Rky2S3oWWKgpLxWALmF
4HTIh8CnAD4tMjrjq+LbDuFJk5rpNbT6pFNlkm/Ke/MBKHcG/3zx3bohTilQ/l+f
I/x7XnhrQCUAm4J5ZHfCUbI3Voo8yABtVW1mSoB3YpRUHoticgQ/LDw6kHnzcGCh
6aOWrmCPtrLCAgQwhNIgddxviKNlqRKs55G6mo15dBN+2uz0Yu+AlovKmQgKEQtI
u/AkA180trWHGFS0lPVIpkFmlEglajr8Mo6F9mP9gcyC5U3xqWt3CX3H3FEz3LbE
n7yFH6cBfxb2m5Usv44kn0i7NzxD8CILTUa8BMrc/xyp4mYo9qKS+HxIHclkGxIB
CoGvH3DJYIMSmmkKKAxjAr52ymKnTde8FQt3BTqqcjIdgCrBQLd0zsvJjkaQrTJN
LlH8RIa5dDGcHq/5HgMaOEPfdsTMubNjWhJz17WNAE8lgkXj8B28sI+WjijmSIRn
2fgTEWg5nFTMUGPq+FykvAVsLidOBojSvrPq89abtkx8gRECA/AXASzEaINUEPCZ
PRiDzAXEX2KgeY/4zvCWIoQ59NpMGhiF5qdCv94B5Ym2oc+g426/BSGPniLzwgVo
wbbXKUa4Zc6RwHFRwFc93Udd5vj+sfvXBL8ZAwC9zmSJRQ4Oz84DzM5LpoesegRO
O5xmKqfQw6hpCfGkrSjN6AL32dUorDQoYZkb7VD8klpAeRlY0gd5vPswt7Ras5ld
eZFvcoHgfrcyPG7sPukVyGGbxuTwH0VXxt4iyghKakVLx9NPmZlKIirCMo47rURZ
McbHDAj67qp+OK4XOzgpzUmBqAvxGbFMxbs9cHBidtrl8TC7JdGFdtccchIuBA9S
eclxrZ1GJlM6B50Bj2RnZIOdRMKJWEGuQ4yPoLu63x3SPUzq+3eXCoNUOZm4x5aD
olTiZaZgcZ03a2wC0T8JhOTrMWH4GR0S/oABryvfIzdKw08TbFqhOpy/WMVjAnrs
XhgIL1duCgK1Ic6apLLwcuGWQs7i8MGX3EkkaXPp6zUq/vq/bWOkMefadF+nSql6
KFJxh8mNOSRwnVSGDmV/g1UwqxF8BUlYKzLsuxpp+ANHnqscsomCo15ZqBw2rB5F
q9xGNlhIWfmpdnBtHBOXwbEgNUZxMRjP89BHjx7g83H3Ydo5EjZzoiVtlmi//KwA
Jw0blt/s2kAzLLA9XfmWmI/8UEBMwJm9AUPSkbPdVMhYJo3lvJ1l1TjCjgYX1qE0
NoqS39o9/jMcrAZyh+Szkp8KAGVGd/Wv4HcjL4A6tvAgB7nM+4EeEaoLQEcIZFtu
HeWAB3pi0J8D3jIQKp7E87GRgBMP0N9MB8FmlWAf3vOscmDCRt9qro1Ey/r9FFfQ
T8EyeCDFIQ2mMBsJb7ozF6VG1Ov9KcM8YoU9SGG0SvR0swGpHiZPc+q1qCU4Pl2V
KZocJFMYppP2mfWlsZGyCYph2KB9IfPmqSc6bZX4OpfvJz8HBf5HJfLIHHAq7b5+
QJ06XFgaGlahQvt7iwDyt44PmwNCyDVXw+9mQJtTRvuRupA8YnUKwssDJV7zd82k
GLKxlM6xoaymEVz/IqP040XfOoVIF7AsaezJSM3+XbnWXuucd/V9Yx2AOTgUal3c
WUIqitqEO6tjENmaGE/k55eRJElF7WJGYZ77vHXuu+4qA5bx9Y58IxnMlSJBRbzH
4CVUaYdmxmVOa3MOVO7a0Je008AyVUid0bsyU9j19F9QyS7tOg7Jf/zu/K5B75qX
Ai3dK17LVdH3Grn8NlhftOiWNyPL71vm/c0X6SpNcWDSBMG22EBfoxItn3JwogI0
d1D8rzjyjpUgnqpkwGb2+cEzjEdNBOZjv4t3wYZBJSCu0X41wtkZzT0LRbG1ERoC
wlnU55AAh3l1x75TVTGR0rGSGwMA3brkCjADrEqWkDKHpcdwu0tvCQIl9Lkwbg6O
i8BwrT+nVssRGN0WWmcRN4aMMK+fAegHDM7q4zZaxmNWoYbN2cvJrwGTUd3fIdzu
FVSNN+PuS6ihzCwyTFxw0Jn0oonlXgcxG+WR0IcopAArbWr/rF+qoLTiHWwOTy2q
g0lOChQs1FjSIr4BxIA2hIu3ZV+ckDc1wvRmO4dMy8W51c6H+2+xkq2dfdYSOJuK
HJUocyG21DNbxkicRofUCOc4nz43L59syJ2VkzsTXIlJGCVC0zLbN1S2evWdv+I+
BzlRYsA4mF+E0wjYNWfOIh7zqlSDEPzCm/s0iscGnO2VI7wUR0TTktE6OgoiuVui
GautxBSidn3C/CHDwT5iT1bafkAKR4OrKxRHiVf4ZtOXHyvYVrnzPnA0gNpvCkjU
/zWxqBdWVpZtY71ZsNNZpij2xZA8fOaukoJ5SkC4i15KWFs9tN2SQf0+/3jQ8vwj
u4WfM4a2skIGVT2m8nnGZe7c5rlSxHD2kYJw0m68Dn69NhoYwq2ZDUmZNVi4EjaX
THNz3cxBj967xORyFxM1XAPmyqh+IdiRFRP+Q2SyRq7xDh7U0vNywabGhgXsxCWI
F8+mdyX9X4f9jZ5rcVu3k1awzjVP283xO/ouAwjL7L7g+PXaTdq0SjdWZD3+tGT8
FKb1YOBbctjVQuz5SECO5HIpQYK50tHEc3HwmChuDyOl1uqLU7Os3YFcpGZxz3DY
mfJj6j89cmukpx1Q/FEaGiuvV/G7FZkbOGQ//l45cVerHN2cnsuPWaCm3SlxN+Hy
VqIZvdcUdisynHTgq4xah3L5fQxmy8G7/pGXR87qNvNiKXv0UVdY1Wv4ekRXiSuW
3XxH9H/60qVyAVHpjqCap4hFNE93npP2SNUjqMpP0F7XE41aftNKBlbSEdf5wTLo
xHGMVEDP2oHFtzDo/6eKjgOF6683wN7BC4L7C7cbAFZI8V5SCA23zMWVE5Gxkli+
m1eDsckSLLcmA+vSpdIICFE21+3R/cK8siRLcZaUc7Q1nzDQUAFZQXBogLrwXE6i
jcT/qhtfaa4pbRj8RLF7s/eWa8GRR/aW8gDbc2FS9gjE/+8FTErVxwVeiVdsY8bV
2wCPpuLkDqBwwh7MFzEaPKZnf7rJpltRTirqns16r+xFdLjKb7KKRuSLA6YP5aLg
LgwFz/Vw4hubuXXiCSB5XYJm0DshyBZTxJgWlUjMjCFQLuMQvEuJGiaRxjA8QX15
1SEGTprNr+gS3mb29/vHSXa3Zk5CaTxVpek6TGyDUY87exSqRGUGCXHt3aFuHsRf
cOSw/+esyMX8x/IpgoO2ArdV/S1HFQRXPWCXBoWsViB01o5lfNEtD0T3oev3HmIL
TJNvk2hSqs9x8i991xl0ff/dDOeHWHC5SaARHLrF0zi05mnMkIoIGrJUAK+CrzGx
VuS18T3bRylemZP6FM/m2S+X7vHBPaWZRV/VN94ZeHt1Wi9Gvwvmr2QBO5umRlgk
sNGOFwLs/+1Fd2wOiQt8D3UNEz5l3g3BWR+5DXBmvUm/cJ/XWG4rX4N3rTcurbY/
0nO7FmHHTwiulroba13Kyy9w/ZT1623FmVT4T9K/FO2SJZMV1HzeneveVphkHFAd
gGgkuI++x0kY0Y/olK3ZchKoFY0tnV0R6wd6A5+bKKUpuSikV8djZVAzWpJAZGSA
7MbP08VqRd0lOJRDg6kTBtmSwcMrtAuaqVYXYPmdP+iP5IcOyENYdbUmQeiTBB0V
GVIpQ/v5JIs/ZhdAVnD/BobqsdyMNWnKzTn73iVEoY5/TdeBN0ELGNn2B238KrUf
N6Ux+yyl1fUaUX/SKOy9RngKnEFL1LwaGIv4gQzTqSmdbivw/nq5Lqdye0NCVX45
bCO7ItNrNehVm86d8AeJavwuAIABVLeE0jmNqeGIOPZUGyPnPYiZiPz4aH0dD6um
q4DD6YzbTumKnS/BQNko+5taCKa668xQqvrgJOU1b07RPZkFvYmdQbLZTLhbllJF
zWD0qXPfyOG/TO2biuOOl36gJjqevOuvwKhlQvxsFRHorUPTtE7nFyO8++FwnXGu
234KoyxEt76rQdlpUhnnyNT07UtFFM2Q84HpcWGZUYvLifubbBAvsEjhpR2VeFMd
JzqYZmEwzTMC7t24WkPWeVTcCylQ4kB/UthAX1HTqAg520CYbshWEUgZPlMJqTq5
ynP173h4YYk6FT72bScX03Zd3LfWcjTxjx0QUTgMNBOdn7xw4tRJKLe3Oqg2AWcV
1YrCAsDj0IU2H/LJRp9SmDU0XzxVr6xSgdJg0RJFS3hrQdw1tKKEJiN2R9+YY4Yq
O/7w9IirLaCHu5q3L8dZzOiE0gcbEBNytl9hajfvxckbucXCKOb0LPaklKr8c5tY
1Bmk9UovJ3Ptm+5n08M/Ys5HnVoDV28C40xUVvO2PCBxiOvpWqPiyjp7hU+zDY3A
KbLFCBNrN/9x4NMovmvrtRUGnE9Y87nki6Try/7CtRjBb6TN/yWQg/pWMqdS21JB
BGpoEAs2ud3+9xI+Tk/LcMCNlGUfGfyY4f6WTfSfJq6KZZ7kWOIIpMV+JC2BpyFV
u9paE/VnLEb/ungF3hDhVRyO00Wt+1dtx7LlVPXEgk2Gth3B1vL3+R2JspAWFtWx
ID3RDVcvb36eooiXmOy0vK43lGOrPj7XOGmCn/I/iATnckUGaOYcDliB01Ssw79c
VrPdIdiz8LnKNLA0QgUvhdb0pgBCPz0l52TpEqH67VJvfSj4VtVoNIWYmW993F7V
7faZHMMql96AA+kLoT2ZP/i9xhx5ZAIuvJssLg8B/+xIbbzPotR+V/wn9Pwl8PsH
pB2FwoUq/iMFqHjwAUZnmPyHsF9g6zbgRpnT/ufMwGcGSWigfE4UY6Yf7wkGFMc1
Bnwr+aEBEDenYsUMg+yCw2mZKJATrBc9BKeFitUetPha5T2pswogQ5WjsyNdfBUu
WcEFoEco6fmRO/iCtCkYryOCwCCuiKdwby1GR/Bz6dqnlUMUWvQgoAgbXkYffZyW
8k3jOnz/njH1clB/MEEwirPfnzVbBUbt85NGT9P48ESMKMXfdDbXOLjx2AXXVK3B
/1m/HHxRMecToyVs0kfI9qeNCzJBYXMrVvOF1auLNkNkR58+T5QN0brLZmEpDRZj
gA+zJOdvRdbLNM3DzKpZN51qUfO7dIvRzVcyh7PNWsR9F6ptqh8ZaimCHoTEKrQL
nljRCBCRlL7SM62SmsWtSM2J4gLkHfMAdQ4aYqoloGlyaJ9TKON04ZsmtCbGW9ea
7QF6axr88e9o3s0+9HfY/N9HiSRFL13QTSW9mZKUFNBVrEPbJ68JKvpzWi993gq2
b6U49Unvt93mYTpYt2M3kcccUhGNioXuKj8O/Qa5bTWz3zv/Mgt/aYsYZpFKQMbs
wZItYKY8mJvcTScNGQfN4QAL817jAwCXyymqKPv+81I03hYZ0HRYiGrfRLI3zCdi
xE8B5/vG1Px4mY9aR7zSCZQktqKcL3UTP/zuEnfktW8ZCpw1pPJ3dvyOlvqWxpux
NuFo/eyrHwLG2FVVM65320zES6ksBp/VidVBWKuT4uMyiq3lipXUIeS7NLNAO8cp
cGWzcHHhc2KLxhDIKMJ04rqplTq4tYvbjWw1bWVRsK5isS4nH509k/uHgXunxIvM
Qk2iL4yrTSCxwVunO4d0KBByni0+KGGnfw/wN+sOmNZnalJBi3OSe7NvPDNQ1BBB
OI0J5JBegJEM0ltXZE3/8n8d+7Cycg0H+II9DgXSWyRoq96nkVbfBFZ2RR8UgZ+V
funMJXGk8YXGrTnP1CZOQSZ54C01hN6XYBTQF1dIBwAc8hwnEo5Bib0aVCRop8Ha
086NZvZJ89LZQBkwnIJFo0Fi6UNlN3mms5XThcd22ZipfeNQm3lr9PB/QCXhkYUD
JLiDNNoO6287ImVgDpL/xrMZAGPqNOXDHYKNPe7ct+RA91H+FZtWCIyDM/7LfLJr
x8OhK0+eEXZ/ZkGjYi/hQuitI5TSG4XFhffE9RAXudXbZt22e7TnItZ02sHEpJLY
KKKf39SCNgOsUtnW+gWabckzJGngolzeJTfhSkQcb2PjNqwirIZm72DGivx1/YJT
p9+tXWAX5HHOiA5FW+vi6sRih3nvBjrXsWxXLN47WLHVwnUwINam+bX5Et5hYOSl
ZfCTdKEtf5T8ZVbDX4Z8ZNhwlGEr4ofc6HR0kT38ode8IbG0gWsCdw7z8LwGyZwN
HK7dYF0GxcP8rxmNPi2E/d2CElmM+7fe1Oi769aJXuc9r091YIiS3gkCCwSEIfmq
z/j4e+s7dX9ZX1I6Zzr6NuYD+pPbhO6kFIX5DQmHamclJnr5X3S9Yb2zagUr4PcF
HCfCgP2qL6cDe28gdBJVw4cSkbsNKeshvr2iLKC4cUGqHmY0wDjEydl6TQD/9ZOE
3l1IDP8yXyth9/mZGzCQPn0bCt9HWs1dX7+SQoiBF2jejXbERQB+x5yhb/K0WMON
qxGaWPUAFonaA1NIki59Ah9JujCyYMamWwVVvelj12xCgFK6ZK9NZ3QiWANJGq8Z
5Ya+6x/6NuL0djH+nct6ApxIYqK+OjLP648tQt8HT1liFUuDlfPWX3bZny9VISVA
QAkqQbRWCbJpGRLtCVlzU9FCfg98fcMMsgzCSa4xI83UlhiY7xXa9EcP4d800yKU
QtJLpA1GSnzMXkODRRXsVz6eFL2KoWJq2L/u+ZyVWZdhvKsPRzc5LM+KzQbk8+P5
sKo3z3qmQLijFT4txZBgHMJaDW257MUWfaBLOI7/YCxyqrPWpEKKvD9gTMkOjWhw
8Wz8leHgugrrIRYA6aM2exgARU7ahs4FrG2gQQ7wA93MgOSFa1ctx7PuxNfK3NhI
7KDl2SyDh/+ZO5ogw7kCBRt96nCWaQWXPAYlvZLXvB65u+spj30H2ba8Zd8+peiy
C6nyqg3EW2P+ikRHuvH0i45UqNmWXvMqouLHy6ydnoxrjOwX/Gk4OOk8xfCiGAaE
oSo9yR0nmvIideVv2IZlzP5ToQEuTA22Ggo6lJDHNmDDt7V7N+mhmrigXpFBxIfb
MQPWCvIWG6cSmpP7GKlsMEYMsgcVAfMqmmJeqWW4hT7CuSoV8CoPkQ3R4SnoYaHT
em1UxPe56z3QnPa6TJenwLmG5OEdiD5nweWTBzeaoLIwziwYf6I8x9IyRIGTKiHp
TXyXBG+/O2magl3R78P4UXT3p2VzroWaokBzAAa/J7vKvFbpZ5Hdn/AfTCbCCtng
FnRnFV6mATJbnxmJMjv2CMJz7g0+ovsYZiJ+NLwzrCVF7kxEoCVKou9dMGIL/gop
aP1H1q/1ZxRua90yqxmFb22spWagAdCsuwPaMbAUAPY3YTFEBRfLzLi20Gomcf9Z
Yrp+r+p8gfaTqZx2huXmFJDf9LVbQmcwSToet+Yn+QEiU3D63I96mdxQ8KNix+KX
MBAGUPf/gHMHX7/nHbnvyqVaGpMDmwVvl1h4sp+WrrBXN4bKSiVcBOL/W5KZI27z
8N1pgsdU+0Bs99u7dJvjQjF8V8zq2A/A5I4oJ5YgneVNsEEI/+3xTq0R4vs8uWXA
Xq7hU+zFmelm/GeBklvfjJSl7TXvX9mgcSXg/DC4M+UHFc4X1IotzH4bl+865jOT
U6/WJxfG68PGiXwSr3y0ombETl15LdDRN1kg7xchO7Uv0EIocPaTB/L30ZB4sr6W
MgJoueoXRhHP6S8r7hrp0O2xxd8ZMvIsHdoZ/NdLLnpGxH6l7BqXCdm2uY0rvN/E
FykyB2KedJZ1tAe4RLPqDF5IBsKDtmoN0rpQfb6gqRGXK8TxKYOGPAxVYCa0LrpM
gYDqlK9H9ZZd7RssKlfQ0oDKYo4YAKEJP3+HWz8jGU0xddIkZcHi4FlaTQOf555V
LAGHaOhPRkWgW6WOqTOjOSIRbDP30SyueiHZxdPzjJwCJ2R5Zgs6gpHYyWyyiSRa
zuDQdnPPoLu1UdAwqsQOvDRjWf1J5rRmJwpkBrg8MYa9b+YOfc2iCPSF3iuIP6sf
MZDfrIQc9ar23rMBl6v0Gj48lrryJ9VfhTY2TB50IshjIC0R4aiSVSytJxhcx664
ht3bslDfy2tma+0KOiiLXDBcJQz+fEgTAvCNPK1L7O83tEelft/MBjsg7/ZZiYpA
f4w1GL+qkya29RGlvTnRb9QQZgRXbx5lpThIyL9zVPYkX/PJMpIExrJajl/ZF1KY
fqL9HRH89VmbdC3s4eLJmkxtZlPsBEuAajfrbfnfr2pOOYgiCwNv3JSqgXVtsOwi
Sa1Oeqhcwxic7LPVO8+/hIAFJVcS4tSn3QDi2J0L1nDlGdNnOIFhtjYo21MHhlxC
r3rKPU0Vlgm4bnAtrf1ZHfht31VbEQbkHjgijCjEgEqefkME55NCxYjc9k6bDoUa
f8+Dh0PzIdwTT0kG6gH0RuUTKiLf7oJyJOCmKn1fNA2IQKKpyi+kyWTkagh+p5G3
QDaXMSYzQMHelGiGGCPbZZ4RVxnvjPcOyKQDbD1Loyx1eK7ymTAi6OjNRntx1g4K
vZna1lKVHDjm1JnXUfBwNQJ1cIU/wC7Q9RSbM8PAC1lLsgSnonwBKxZKMnc59GNE
AgaV4F5WpCAXyDA7Pop9DpxjHjr+IJaZJI+VEEyDwqm82+MnF0V6lPc05/rQ/Xc7
mcjjQ7Vmd2lBJG/4ZEE1RvM5IIV4E90dlH2xoTs5OV1d2uq1MR5rT+eMKU/pE9nN
le0BhFfseJ8ppEvWIHyE+YBw3g2I9RIbacHl34R/yLULb03P229y/3DQwLqpXcGw
zc3zaLtJ86KIurMQjwelZ+HAKY76MuUOtgng4Pccde/kudxU9ZlzPct/pLECVjhW
NYA6O/hWKI/UgDCXFRht13MCXl9/6XdORMJk8SyjtSX3eJGWkkamcJC6ua/V0bo6
AO5ZQYW5YzCuHdoQ272+tviRk4XwH+RAb2K0ahF/R9iG4pJuFRLuUcJlHvi4yB5O
J6la9yRO/j0pDxdSvfVaLtEGicYesFOm+zD0/82sMOBx3PU9IR1NwBtYsjmrya/p
z9GlsLJwbnqL5pBIdtH4qMn1AE44F32t6Ow/1LU/pWU7YupxtqoOZJgQdDXzl4Vg
6qqrOD9Hv7eubnPo442QpOngh5wfZn8vG8QferCZ+UZZxfhB9GNKfheHTbTqe4th
ZbbWv0N+K+uSGzh5ubSwqTGwnpOeaI4t7ytRsm16m/2+VU+7k9oZ5zf0bOLHKCLe
H4gpAJKdJK0A674iqs0I/iEsyX6eD9KhHMOfJ9GfIyKEFZAhroA8fY5hcG6MtUbX
muqvmiVF1c1B5h1FUROFkY6MYeQ7jNm/Owsyc4QBjjPTPxaUOl5g3gXI6e6NyKH7
rbDvqFebFVQPq0/+oER/AFt0MVi95pMT98OsXxd9CZEae1AwiFMlP3GdjdnwBv/P
v9xFudUPD1UPjZbKZ3yc2n9ZuiArQN7HItJiqX0NhG2/nrdw1h+UBVHNPNp2Il1w
DwG2n1FrRT4lmxUfLhjXzubgbZYQrnUxA3U97fgU2Rm7DP1tS3CruXnpPX97fa01
QCa/5b6k54UD3H0BDJNdk8U22fFtTLKHFp0tj+j6jDjHo9+44J/tcVBCPn0Gdbdu
Q9w69VeHXeT6doaLzBc0+L29IcZJpNx6b/gvzq++MGDE+ayaE4Qbnsm8XMZXJlc4
bP4TTxDk4DrMM16oyicMZwbp32G1TGZll+O3h6kJeTufd1664oW/bSi1x5897P+1
yQ4rsFmiCDUJeljEfc1yP27BoHL2iXoTCxsCRSy9iLTYLYR2ibXWkL0R0EvcC8S8
YR9G5qhLnA9ozQL3JQHfaZvqOWwJJaDS/6Xsx59Y7ATaAE6DbxVbpcLf0n37+Lr3
9m+HPK9T7z+BwoH6mSNYsjNrgoliLb/0zswBssZyCzpi/0VLMB2d/z7UjwtXaHNM
lD8xSHDCetk/zhugcOZQM8PSAG/bP2v4kaQVxqQMyzd0mENi7kbC2uLScZ+xoIJi
+akAw1lGBcKnRQBuTgjCQlbIFy0o/7wnbERXJIkbBkj0QI7H2wnj0zDUvluBP5j7
5B0E/denHNSxlwGEyLbRIEUX0hHFEe3RXcTCYGkHfDUYc2bxjj6F8lXJzfM2KM7O
lkEMJTvn0YV/6/kIH7mdFpqxd72gVCQ1Sjrvi16sYL3ytTg4oPs4Bde3M7ztzXwZ
8b2F4riBREEyr5oflayL0qFdUhAvSRsL8GyekpPN+pHclHiLKpXCalRD3yvBr9zj
RH4KSbb4a2AryDl3FSeirChUtYXk1nkOR73rZ9LWExgH2+e2dZLnYbfBfe6QAbQo
RdXwn7YFMrNAFc03b/1IDyYHeLT/DWWWdyn8aaI24opeb/8zPDqx8KR4Nle5oNoe
J6WWbgNpgh5szy4FgCcSDdh+OIz/OkFU37tFoP7wboqTu4T9NxbCxgGWAJqFAvpF
QzG5FCqPNJJvJLpOJPEdeOw67fiCIH6YHCE/XUTpOWgM59t+GoM9I3LPgAAx2sA7
pOQmxI0b84TGYGY9wpNyFtdPIGhD4CJYdHAtzo8ZHtS0c8QGGGzQL9YBCTAzf8sB
5R+1iY+HgTy5Pd1fp3kmCRZQ1LoLY2dm9XxxG1SaqYfOCFgXo/8at++3DTxg/eA4
/RbrzSdq3PkMB+v1S3ow/dF9Aw3vvjRz3YDqC/3C8D8HUIpfkYp9ifrQ6shmkIhX
CgtVvMuUAKDLNCAKGpVfdakyEahcSMHgoBsIMVuhkr2YG2MpdQH6vCQVmKwsSrHE
oWjzoprEQ9CYybyALS53JviUnHFryr0ZCnN8/jNWlTxcrHddYSq65IJiuBT34tvk
2gjTQ8ABfF28LcypAG4Wze8tPEjoFJfh5uiz4G3OYfCHKcH3RCrG8FI6VtgDrCZC
TL0+ZutRAGj4O3eckQ+qe/6VJZAea910TVn8Uenj8tOPdOmGGZXs+fxEy7JjovRZ
ziYVhIFD8SGerW9LpIyXPhEWEcTeoqt4iDxt1a8/nOy8LsAbwU+bYu0+Hqyh2N4C
W2vaF9Tk5iXlGdL5ySKN7thm2CvKYjLNf4OIXUuI/FXbVirSc4zTuhgClpgRx0Hz
Gee7wMZ9HTGJV68czZRztFhGogSJScOTcr7Ggq8GEhnwFjnmHqYcFOYxHDnwM2b5
2/hTrENDBG80MLN71HiIm8uekJAzCemqARI3T0MjyxVINOp+BTfwmteeQ5YRHVI+
C36BdqVY21CzUjezxnFr6pSbdKBcsWlM1uAta+kG6DaM5lbG9+K89inuHAq7b9tr
IOzVDB8MxGBz6e7eWFxYdjGss/dEl0jvQQIMROcjudcwcmxIa2m8DpgDaaC2o+6Y
Yyukj+e3zY1DM+q9cgcv8HuyDLOUQnzKfDquhOLO0h7CeZqiDWnlDrqcMBPt4Jzx
NYnAJEK/bimkZyOFwceXxsm3NfLe2C+4Kd10j2+8ojWPJ6aSkSnFYvgrG1vo76J0
X36y1DcPAsSw13/JCNBxxisydgdPsh1Lg/oS2DvsRCpskmcI6eewQNk3uQ5Y/vvr
wqhkyX02dGXxBL5gIg6vSoDYX2lMHUQKW7wiukQ4hsf8uR8z47zmMrdjvPBazrsS
ELG8UwsewagySddf0LHS6BUKcKT5uS7OyRzL/Rfae4a2I9lAwfNvS6RGPRRMkWQ2
sYXd2hkqN2xxJBQye1wSypQ3U0ROIxxloHJntoQeCJr69mE4x1P7P3ck+gMOZuJa
gTPNz0SmqevrkWCw8hv1skOot8snuy72BgLPxZLJjPf1U8s6CG8RTd3uQshX43OI
V0NdQf0CaZRIGTra8d6GKZV/DEIkDAsQpH3sIEdRdWLERsksU/OtQmwZ2Knd/JkH
vWUh7T7dTwz+xt7JO61X6vbT4fNMaTdPY/RaE7jGBECanaR7d/+/FYTWBL/2UXEF
efmtfLuWJL2Madyj1IzyJzeuIuOzp8wiDnVlUonGROnsj+HWx5QcvyaLBOt4XRx2
QCLeUxKgE1kQGHzVLefuhtS0koANEcCyr8/OY9YUmlDhMJz4vwgdpmqJyuwei9vw
jNM/vvUyXEsU0LStngRPvijc0T6NCfwhWWYhFgiLq1pSUAlTipWh+QdrlxV+AtTp
h5Ut1HhKLe/3rO/wFtx3CAO/fqzHKlCXXljsGOb8lWumQMT4TfE+RBRPGVwYbhZF
6znhcHyZObdqg5f63fNmRzQ2xXy2OhrWwcoouNKmkIO90t7/2gFutNpxz38pEJ3G
uE4YlBlrW/nKMTkZi7R8i5To1vNe5r6V3AnAQmdGgObPh/DVIuolOcu506zqPEkD
KoZGBmlirovwWo4ZR0D/zImkONwJIPxVOFQhlof0llD2peSnl6Wss9u1y+MFBmzm
JM/VZmSTvXerJFaS60Ryju7ctGfuk5chIu/SgFlcJwUISzDTgJbL1smHuxhkgVZX
59QrwiZBK+F+glaSm2/w2Ly6UpxdrN1q75DPWTtGJMdpPPs0C6djApdCoxuvovl3
SbUgGeQqJnQuosTLUIPTsbYecJjouyS//Igety1K95VErI9VTzRiUdCOcHZ8WJJG
XUnfs9ZofLX56dQKYHxwK6U8RfgZf07IMRyH9EN4npofDI1W83aKw+fL5MGEa4WB
5vj89doFlGhvS3K0kbTqrc+Kx1pZ1upp9G2ILdaH2nexgKY6s057Oky0sbuBPgxX
mKUUi9UPZYXTd4fgDtgPEiJ8mkSvQ/DPuOcC/FQS9LpdD3aWfgbzY754N9WRoH8i
62kE71NZEElvmlK3aHzs2cZG7ljL5+048W3doagK3x2DpG3NkAZpMcV9uClQ6cXy
jqEY7+df/0ZsvnrHcNIlhvqXfXN+kga/qegHVOOXB03D6cRXucxhl5ylv2zu1bAO
CshysN76mlQRLvrDATUcGS6bRPoYbE8j7LivGV2J8QljZVwxr1PRfnSaLHqOQ9UF
9ID3ydXSGs7FRpJG6KIDXqNR1040ZB81DB3i82CVXbpYqS8wXQsfnL0PN9WwgjLj
wZQ/c42pZbdpL/8RnwEtGdLV7bZM3WlhQX6cGkbthOGcfItlpwf589E01n4t+rv/
05cNXIO6wLryxMY8L0LpezJwFdZXwKVHMaf6m/VvyKu01bsSEO049/lbqOIawfxR
+Ggps0Ea0e9y7iVnLLnjRHB2Bo1ud7yq7r2wvIVzwxRhl3bDYnkIHwubsVuq/NnA
miLcJZ1YrUeZ2aSMR1vlpE5kIMKwEkQnyZui38Qs6tFx1KCGmD3Cw9QvYRY8sb3R
gFf5Kx6tOPFl1DfzdS1SS/bbcqlre2z8KnynggdH7NopEL+1MWdMDD9I5bL26l+p
hP1j+1mKM0PFapRBj70Ldzo6VARagvFw3wMIr0u1UAE1APlZ7kqGcrqKSR21ARHd
9DKd5BU1XAyGuGowso7gb+lKSCOxybZpdiwLsD3xk3tuA9pLA1P/HxzCuDJQIf+1
JAvHuDNWyT/JUWwyGCm5LjB2EEJZ1wlfL/s5xOe2+KEmNQhN13pnUOF/ltmit8nB
CmJfW/tOk/dw87BIhUvj8H/2glC9bs6Gg4XVZRqFluVQUnrbd1MrFP2A7lindwk6
d4WSxKnkDtSLmFMgq9xEo/DHrsj5QkQbOCcccrQDHbsdB3+858mxEUdJKgpeLdZE
RoN48IjCvb5tmfB5Ou563RKEH7mTKhPBDde/bJ7tq0dGviNfMmpbuSlaeKl/jE8R
DSKyNEz4xf3aKVdINuP6My/uyOLU+6Zwb1Q/ZHwn0QaB3qpcRps+3SJkQNqZ9++N
pjZikCHkeCfaPMErfn1CbKLR7UaoaEt8blOSMng1BpIiqxT6oC41+yE/ItvFspLE
JHOglW5T7hb+r5M7N/QcNHvpvCHw6BoBEEn3WRgM6w8xdOcTRfQNwpkXkVG+1zXF
NxP7qaV017q/3LbFRKyz8vWbB+bLX7GIlktiRFZ/3Y1uLEGFojakFtmsQZHbvGrx
5qTA7nQECWxYZIU3+KZmQRo2jReCaEDGV97CdjbwK/r2fjB9ak9KX9pn/CzvhPPR
2f3ZLAH3hoFsTfgyxO5+xvoHl0EsCOvUHXKMjlKj0TVmCn+C2fvIK8R3aGV9T7Io
Ls1c3HdHbR2TOOkhW4pLNi6ocaHSnIUaept0O4/YQOgBiL3tdbRGGedYpNv8LCMi
DEim4ydFEV9qJRHMQtZlVlKqNWirwxQPWmIopppIkiUgB6VoxKFsMv/pM5+PP5lw
TGDuWytEp4j2sd8E8fO7w/lE6Cp9heUMaAOQrYqQffi8juIRC4WmAILWbDQ6DPpf
Hr31eyqmywduP7h1JA08Ogrplyi07qDrC0UNn3kyE6ddyf5HhCNAEI4+JRRYQ/i/
3bb+Hzf0Vs0e01wLBkkfU1HTd1JDkFgt3p7/8zK/ZhMmjt34YDWxqIkcjqF9B4lI
ZCij/MjR64+5nZvQhCeP21Z+Wcv22oWmtq9qc9sNp8U2vH/uYGMUkB4YsRg6zqFf
IAdgsvD0r3F1YYsY3i0Izkxw8/j3Elux961ND1dIyoX9zt+b0Pij/EDdDgcUolNb
2McldimFt86Afim2cWnNNDhXt0Ex4JKSNh0u0X8I2SI+BT4+L4GpzUMFOu7jkd/g
I1GLJHnNzwBSUF5obb7zEWmRoJx865RWsZjodOY+d3C1xltWSsM1bDd5Vqc+chua
k5p/8iYro4bUakOZdnPwwA5IDeo4jRzg7P+/k8VSvQgic/Zk8gcPGtZT9Du0CsGF
VbwzwsGTkeejAeG61bWWPor33Eio68Bvtg9BY+jw3a0L4XAGPHKTAEFGwiRcPzXV
f8y+2xTUMFjwkNprh1vgZp3pzpeZoSeAAzawQsD6ER70NogFASHoeVIhv8lexq78
Rwbr2NO9Yfe7K3OBxbbm4O1SS9vAEWV9vvdvYRU3cBOBF7dF0S0k4W0CdfQPMM7A
OAm188GlRXZmVxCeGwz9a6gCZ1GY/rGxhqNjnCAMtI5DrlR6EOSQVXsHhH9EdJ2l
NYa++lsJiTxQvNgWS7AU67goudvcWJUpR5XuEdh6UToJQp8Rq3IjPIIjc1GP0cZs
/HuVfoA52V6tZiTr0AU4prE9I3Ord4x3XV8qGeIZlOK8IRFKPlBxgGs29vV41WYj
4zJP6IrpzSWegcw5aUYyA5KcPtiOp3ZnJYe8Kn7CVqs49hs1XHoxxJisfGQxS16S
yByHx1UuesctZ5XSLL8tIjEX2No1xPSxrxWxgYTEGHX83u5ggjBm9R/D/vB6HURI
LhVouwQuF7gSfY6XceO/6reI8+Ty4B5mklKxkw3NxhoAEu7SE3Nh0vG+KfRPBTe9
NxU+9Y8s+/X+tWo6tu6KM82zTwhW55Kyv6CGd2C2zjsJtKxE6LyQXor26gjT/KdK
gz5C6ENP9kuIUvc8DMvQcSJ+vOTEHnz070HcutDcyGuQIBELhzQNPZs6TOf/c1ya
X96BQx/TcfbH5GxS5Gv98bjJpcHrnwRg+A1uxkznSitKcRJ3sEKYCNJ9JQkUs93O
Geqc+cEeYIh5J/4GRI5CWFJedKH3Aa23vXVrLYtdinXjI9gFU/V6/k9jBFwFcE5S
yGjd3ZBB339cMH3CNxl8TzTkBOhzUcbE1HL0I1QvNJnhvn2EoeRkNcokak82FevM
Csw9ey2Hs3dLtCu3TfGKCIn76vpMQ9WL1KawrOmfRXdewTY4kDaALBLPGVoPQeFm
JdMd6qgvV6ekZG0eYGLBgFva7Js2Bw2FqbpRpu215oFJDXiK+1PryJlGKdIztUCA
mTaYfYPIRiE/kf3smTL0P7ZTmOgcfekPsKYC6wxF/hMTuln6SJUHeNV5fSKbSegv
NdXZgfDgNJ/1YazAhLT3FVIVP2ZobuJs42T71L29+cQKhkJye0upCq0ldNaCBwvN
aI7lWqrTJCZBp0/lQG3/a0B+z2ikVzoaqjezrr+3el3hcV6BfiXAcVo1YCfKX9LY
wW9zgPfm3J/935JoCGkgeZsXTB2iFZiKmK78nTBkMtnEWQwz0Ip8a2g/XVhpSRmq
GzBpHZi+knmXC3ahsoCuosvVmutEqdmTngd1uLnOAHHx1LtscNH4uLKJeHCSZlHY
xyKmmNyVZDzB749AcgPP3n5AjCzwB9tNfpJ3lySPJlTUpCt+DlWMesBpR2Djq7ng
0A9apr3w96YSWeyXlZN3g8xJB6a5uHsvclQoklqyABgQ3Hu7wjKPtPabUlozmnzz
0YL1zZmgqhOa3H5Atq6vTF9kDUEfQCqIZJ3bWxZ2w+itXYLG9+AnS6U1TtAmDeT9
7/dMu/okZO1mpjUPCxDnvIX1pVAmeHeRF/p5AKWVKDPrMzEJj5E5i4hbUXcczFsu
jF2gBS/lVPyctvKNlzW24DcoFxAvRDxIvaupopP5GsYl/QrM6YOyhgpB+4FkEnME
4k5FegBViAw5GbkCZJUKAUTRPFlTPy85wFMe7QLidy5q3qyYHJUqqDpVCr1rcPd6
G2pbJZkOq9yaMI1yJ6A1aP2z6J3SEp/77VLS8IEb8wXJvQs7gPncQBIVm/kzM3Mw
OIdGziNHv5739P7q6K3ZIrI9E2mCbUxleZKqlDziK7b0FA4KBAQTM/KPVCn8//J4
TYnVqGb4SHNrum/FYbFWgOsqPN3D5dHF1YuR4UUvVxfJ5jq4f7zEt8WrWWTMPkTe
xXh2aKoFWi2guPGF91AV8HyIlqTk5UY1I8m6B+V73lVAUw6Dgs6N9BinSnLKZQZV
2cbTKbOHoC2kjy5zQlASebuaqBX7/kyZp/4DITYGYnQjlGJ/w4Xxs57Ie8GLvXuC
S6p+o/Ajvv9NWBrAjLh7QYnNn3OK6yq53IlkM7vIAKAGHxnOQabNp+7rA3eoGoW5
QWmbGI+xsf8ryLQlZNk+KmUZfeenQo++Z/IoBNtp2r1S917w4bAE0Ja2YahsjmYT
58sLHW8FR+dwGSwOr1TefETCo5fxeYAgN/6DGc2vOD3+5cul1hCZj3QvWvx2BSqd
Ag9dz/NVZ137xoS+4yEY20mYHCcAtN4dH36YyIxiA0ow6ec3d9Krfb8l/srIoSX7
0jDIRH9mic6qJswIDGRr9YvxGP2sfKIvV3o5QkKvQKyPACb1Pp/QxQpwGMFoGe6N
FjnZCR9XZyV4pUEzhbVryo7UFzuWHrqVojL+4TQcsYQRU56nZxqAp1oI0Rp5D5xE
9a9vLatWsT++x99W2EI5ZV+XzUVqTPNGdJQ8J3YlN0UP43HeLc4wx4q55OWymwIX
melWJYjzvX7gnPqFGKmB9vG81SDkstbXHSdvEYUt3BXF5ZszxZIjFwFOtgK6WTjL
/6H4rXkmJHnAHf2IgspFN5VzSSwlCj6P2FnCQ1qmLcmIDnKERgDF7VH8S/yXfA8Y
MUiEHUC4aGWv5eBvwpTE46AypFBrezP+ieJU4s7UhOuBq+RMX7tn9NaYsZ62FTMz
GkJ5cu86X+31P1KwS6ncTEj/ycxgv3AJJ2fOkAkGVJdjQPriYHsD8yjmG34dSDX4
OfWJqZ0HT0upMvJ/DpheKs7UU6IGfBgEOF/+VeSvDDBxPPyuPoGREs4y71+isala
3AbYARDkVusmRBcc9ugPILQVE59PMJzjOd/pyukLwhgk/cz3dgtsdOIv6EklmxaV
/Xv4oS7oeyANxJB9MGwexn/CUdUCNSKH1Sc5JLPSwq0THJZcztqmkff36XbFpFOe
iK5HdiJppy39TFSnwl3pPjONhrz4vWjxpX7HMA2ndskrvkx/UIQhSii65NxjHekY
xRKYynK6JnPJ4j/EN3ShfEZ5K330Cht9npEz/yUBfsmlum7bZ59kcV3iB6GJB0vI
K2citKddqz0bWMJnZLY//jCKQh5e6CCBZwDnviG1432wj7/X78LHA70aNdYeMt6z
U/yUVUR58dhsrj9APa8z9wmFqfRsya5rUtMrUGGTv3JvEY0w7Fl6K/sR1CnJu6wQ
inUNUyMLL+KrRcbwjXpoO3ti3UN9P4AiYNyNakgZ5sl0gAd//k5n9K7yByYsdpTm
KhjkG9qC9OYSP/R+2gIjx14jmTRpFVFrw/D6EyPaGRqsHE90UQKtm01ZqRDU2Bj/
Xap1qnq8MVM88CeN7mc0bLfLmBimWxlwRTr32pE78ndD1YLMd/h7K8rQwgekjWfn
dAKpPlu3qEKoRbFSkRqyd+VRgA5Nmgj4NSZxU/l4Y4PfsmMjC1kHLBxKk6Xtts/6
xCNpbFxpPo797oA/3KZCOVZXA8E21nkeayrv0zOxkQj1kdnEOJEcIgHrPzikXgAO
PDwmPv8a8LkKngyWBz3TcPWEQFhRLSjo+LflE6tBwACEPzc+oF/ASxZUlXEdqDD8
aTx+aLxB5DDUrXqKNqvGG0iv4FCaRHTAeEoElu708lEFVLn3SG20k8xdjB44hvEd
ZorXNn1Om8NBrD8Q3Z1fnp24kX1sI9Q/c46X5vbDptUmNK98AoPyQET4Yrs/3oTR
kmLR4+NYikpv3c81UMP6nwFUfmj/GOwXojl92mVMjElSBPadTdqfv6TgkL+UT1nh
fP8vi0Cb4JDPLfqetnYohN7Myc/PHiuVkJCmoZD6WEnTy+ICkfIm09VTpgL6PDQR
lFAJfuivmx1w8/u+Pon0aiNK1tWTaGr813joCuPP2o8L+Z4lN/eMXYRO/WolLcNg
QJKglJ4LM+Qxf2JEEnLCB7/60B6joUpxTPhPw/uMJbagL8nXK8V3gYgtqImPiHUQ
UpRLZ/8y4FOxyvYNMUJ+Xk1lxs6qSV1psaD2zOlZ/qX8srnP+nEi+vlJWfgnsaxF
F3ItY4ukNghLlnO/uotjGIaOgpWm1QDtAn6ccJtBZiWP13/YGeshEjnWbGvyCHly
nyesinoCglCB+eqvMB+hr6aTaeZtImCB7ZZ7Xs/4vRC5FkdekGQQWfbWeGr3OOKN
0wRDCP2CRVhg8s2dZigutzgU+xuVgGygCFiiEbXXjpO73nPCb2Nt+9U/cEoQ9X3l
RkgryEEKojKKxmq6BMDKoeQCrNCAZQ//A8u+MRAvIqBrwQVWozvgvvMPMeCT8fGn
Nl9kiVgSTZskrgQhQKkuDOVlaPa51MNUA4qzfqn/hnqohHSxQfPZAViy2nGBtLu8
j4rlhYZxhqgiBnHPWaa7X1nraJ1SCtY407tlcuwb+k5PmbvivRWegUoIStNdi7Vx
tzRWCgGngSguMG/37kmlfTac2j/qVnjqIgsnVCDze9M2PJ+fY1b9rUBOjCsH/CRL
HC13lrssqq10h2gvBJLwunLZCSMl1P5dORM6gJGC/nwqwThhJD4Ze/ZJYDbi1vyv
P2eV7sIZpWmQJq71pTl0w8bxQZSO7tapVSt1a40HN0DEHK7LQOSFfaTW9MEim11w
IXBAd7e9FH3Zz/8yLwzRPL0nnYdD27br4ahqSSPmdOaqG+CeKK8RYVKPs/PGP0Wi
d28CB+lkuvr3TN11jxArDZCRj0dldDfDiM/jN1mB80Q4ofRmQ9pc35HCLi4phEtE
2YYS1tB8j/5Ry2QVbDK/hWiznmBQg/zTsmLogDsfIGKJhThelA6eZJbRg6X5YfLy
j0EupcvHzGrI9t2ejHLMDoQRKXkvWVfPijaCj0XX9gsaCTOJqCKFby+i1VenWVaD
GSLD5NzjrBZs45NGk2ney/2Hy/Qxu4q5pDCtK81qvRkiq35G6kZNsRKiFywSn54v
Bfjq7+cYnDFeq+Xmn3OKi3gzYzqcprm7M2/nwduFn3h3Ktq2P8xF6qGvKQVUiruj
Uqv6EOvJTwfkGnzaBKVqiP/WhUztyEnaaoVGnvT3BOpx1rnikQB2+DI1zK0e25nb
Bte48MsOeRuCa87ulCS5evl/z2GuHGagFscTocF/jxssIbOWzlBxafGdJQxARf4A
QP5837jfAYVYFf8ODHKiV/M6xVx6CiHzbuNAFUclXSdATigEvkuuAyurMMeCKInJ
ZApo1QjILccylVpDbfsOB0zdloNdN0A+slO7OqrLj8Ec2ULA3kUIFAhAn3isYZq9
lOkfW8xEDUYl4/zPiGLSJs3BZ+GnB3M/wX1PXAgypgYG+PIurrVWL8iIdbiHTkyS
2Z8GDA+xxYDfOng9XIe5/0KngSi2ad4cxldaVQxQ9FPv9Qd3QOzGCLxgcnvgeK6N
DjVMDo9eQiz0z9Ufv4CCUBPoXHHcPT+hXfpPzHD09edkC6Q9qISUsok9s5YPU2hT
o+VLwOfdDRXPaQzV26uxHJivmJaZLYGuomtA21CHoCesfqf4goGyNs9vH1OVKSYl
DbbUCgNRUX9t1z7kSqK7PDa/N3m4ix3eXI5p/PTnt6WjEN6r0CVG5eo7cD8AESKC
HJYL5ZEnm2rSx8CR1t1oDCpj0VaUY1zra5/AQgMd6vroJNByengVkPyzPgJ084Oo
pvIV/zDB0tICNtAN/MseoitnNkYV+u2NbQ/vU/Rm9XiVAcsrzaTXIXFXmpJB9Nr+
rhjX4qsuFQvsDRFYKnlAjK/dprSskvMuKdsuGBoTBVNMEgr+djwpZTgeKqZXjsP4
9nwQfF8kFjHiKRHHteKiq8U3nlslpMZ3Cyc1U0Am46VIANXIEoZQLh2Ge7QG8g2n
dEKkDve2omItiCB5TsvhiDCvWvviE8cmDEqpZaJQhipSZDpnSfXKt/TadUyx8tTK
udPCJ6/oqJDIbqZklC73RptwSFrRkd+6/E0abO5puQD4avX+FnPwy0o5C8Oz6LBK
jXJm54K1c8fG0uWCgknr7n54ibcP93R8WrbTt1s9JHPLMMzEmI3BeXTdhd3PaOec
QGp4D9hSclfA0HQJqZRybFd0Ta2kYzYjsThC293ZxXHbitMONf8eH80X9F/3PJsz
hCXfiV6HhMauW3Cme2mC1uYBIX+W7m/zDYCtxvoyn1hjr1GDOYPtrrtONiSfLlF3
K3XXamaBw4N4Oru2oJT++gSbJ1L/dDZXb+KUgE/qHgG+LxlxmgMCEM5VGXv5ytCR
z56dVXfGc+Fl8gZtVEnpkbfdEUL11pCAZsXgl9cwA645LkVVzlklKf0op4OxiFU3
eTklx3to+btRYYvaYI82FfcMj4wMxvkLhjbcjOFWWzUnfOca7QjISbIXSIj/I1sK
CaZluSBN6nti8rPNhHdziKg4uPhUX0jSG/WsYXyQNmFFnLorfCsgqzgaHtawpe2e
rQPj2EvBB6jFmgtfqvoSR/d/LnLcBGTss9JJR0JrQynFOTA+Nztk2Q6qEBqNPdnP
4wP8FJQmJHMdWfDUEK4O29HnNIwJPMowlR01wzwYvL8cPneaoUsLA1n9lVPGjhZh
oqFJ2xhiZzhBW4N1yDD56lMw6P2eMp8ukzZSF0mxrY/tmVycqlGFo3luR17DWy7W
Rhh6T0twdX5QamPrYBrd9RRXWyAuugxGZ6IPnDI6gz+jBHRmpUxiNEldsXRyWqzC
Tux1VylWclvOmw0OX9c/MKL7AXrikpG869hMgEPGVbysEo2uNIXcRli716YAvJv1
tvtDA9aytUgeu4nBNpUP4cO4e/NyLHfsY7iXEYSbEc+KrN9UFbgBt0RDURIhfDA2
LV9xEBIuz5geGfCcLhvssscprFlxRBs5Bof/FOG1gyfM2dyRR5L0A2jowwiTFH11
+jYWG5CrNXcWIIhw+wLDVO5GcfwczOTYbeZFGk6qO+wbuXn3xQ+/FSaSGwwZYEQj
Wow7IhzOMrgLqO6QdOBS8EXGOmtLrybV+stm+ZEmR4KJ9SOX3rTOX3+lUl2sB0JT
/i+BUudRQkTYUpPkqx5DnenKrMH34q765VjAZOEGYXMAdt+6KtsVuWE5lS/Jkpp/
pxand7esX/TVcWuftYfkx5zzRUZ3ZI9ssIz0vrvJv+p9gx72f94Dslhc9gJvdA3O
SaRCqL6TAe5c6oo3yUZzaU9XQzfTHjS7h6QsCo0Hv9LHdKWVPsGwlwCtSyTP+pkY
avTIshlpgquqcbR5a/Eavg1yspPHYBeu39XRSvm6z94JQT45H3T8nMr2hX5Z1Tv6
SErsHlhqB0Tbu7JoeH6BB5nbl0I2hMxTOrcmO5DlvEopYEktFCnmMV67ly4LQJ3f
z3B0HO2lenIv+EP6pB/1PcbsIfmMQihFNx4a/ZChdZoLnQ1TO9rNW/LYnsPn19Lq
EpVWQSL2yhiRhY+YUs2t7D4736ocpdk1eO+4BobL8/88/Ioly3dNuC9UapfL7PAv
CNtanyFz+5n8eIxY2lAX+maWRLgr6xq8UXwxgIvWPeeAn+rog5bK6tnSTV1NNcz7
FHTfbB91IJx6eE/v78+iAJoR8s5He9x93c6j2UsuCnbK8Ib+6QQxgu3lunf5lAyl
N2G3+PPGrEQWJ+nElWX52Q4VorA0NVtb8VoN6F4QTZtZhPNu4d3O2NBLIe0ruE/h
BeLSJDl7urEm76O89ZVO22ZPT8adgN93XY4EC7/U9HDCkAiyeZr6EHojbtb0QbgP
0n6hv7pL1h9biXZcjHvhJwtUpcN8bz3MwCezJ7FJKyw+Kcul2Iz7qiT+7WlWoO/i
qRXp4U/p6PV7WL1ynd7QmZKBWt381VvYc9VT+qkwbMY2o/yOk+Ve76VTONqg3MwG
RcyJyYbMAMjbYospBn0LBRyHnr7Of426275KFi58Fx5i41xH4TTLvJTgzw65MBxT
ZYMszeJ6XdmanNHGMbkho16LiOFJBXO5Hum7HNtb9wEP/joTqAGTAWy9ww8YF271
qRnjaK4t/x7giJeXL97Q+zitZqDt7gFxnioj5SiIUyATMeAu2zIkuhGX0XShXB3P
1Ce/l0I6ah6H4PYVQBwnuF7gV4ZU9QYQNurCH/YXPr9GzC1HhpR1rCvFr8x4IDeT
gs3OonmB8/xzTDF5cBM/lHCVRB1630fNZVMLZLX6fqs+9bv0TKD+wJr6k8Ibi/52
zYeRqkmIEXV0xEEsFEBHPGhvVLMRrNzYAvLmXvbd/Y7OFvzls00Uh2FuHlT6l8wD
nr4BzKlxL/D2zYgsk8xHUIDTE6vitvlISIKqGDHctPIxZLb6WzV4PMYhGLB4nTev
CIu89a0EuVGSsbpbL/XllWgMJRNl4iJEEPkkpp/u9UileJiVQ3bUtOkYvJ9uj06q
6d9xXhNSBtmed38AgikKjvqdkQmLAPnd9HMY9REeG6nvsyjLBIKN/txrhrtCn1ht
QsFH8TMqG7bBq/tsROQwuvgMATAFMownvjB7UrsV6CdTAUdqXuT6fMVT18u4iv99
4zyBuwXfY4Byy+0EUVZw1cCTxxpu0Bs12pG+QePTy1NYyXGlLXeOfZwX4/KvRM6m
q5Rqp3WZc+6gcATJU9g6aMhOHe8iKddGvG5ZKBuUItgV0/Cp123RtLFH3tZ8oYJT
LHSH8wI9v6KC7tGyojX+zZe3n7yDalAfjZpm1J6XHD3b79RvP2c7uVWU8m/ZQH38
kGHNMDFntD+KcIBk37vG4GWLr0uBPgVEaMj9eMNpYrkO8ZNg2dtiu/1HbRrZQL/0
4pX2rjoPFCzzpYUiHMhXVl+eXU1vmf0pGxXqqTk3oQPwLFovcm9FKbt6tiVkJvj7
6IpjmH2OWXcrwBIrtcayGhohSdcgKbc3t4VtSrFhDqOdgjgmLymfxUGCAF/dPebn
KB5ShXsuE1DLu79ms3GZAtZLabJNoPSoAStgwALMJXX9KqyWVMBzTngMWR9Ndbt+
f43ghaQiI9vTxsw3EKNx5KKxfdl/EYCN0TvXqRunhizOBmeYvLjrAIFOAHwvEayO
MUq+0qTrAEWy7jTvHvQflULn//vuCUVcl3gXn8I8M4eALZlfPtZLMjPZZmqbXYD7
vxFkfHgP6ubPe3l8PjnEzwJutu4o0y+hxi7MQd0S92K5J3mSNYs5l352k2wnsZAs
5npfp26jl/LRRchN5+88JouxA0B/Z/0VLfG9sp67SnFVJvgS8xuxal6r8+PnmTg8
a3H+rfwD6QJGE0/MgXNCA1DBQ+JBAe9TGZhp1CKbaHhfcDCgpd+tD9tgX+gSZkbk
0UC2KdHSt/VPSIO9UaM6N5iVILOPLudhtKK9B0VcIohuaL6SD/dHGVUJMHY9FeNa
vPrA/KdXagfHr4/C2FQtgJbgUPkTt3YPSnyHiprdYOwiDbcB/Z8FI2gKWFxjuwqU
bezfCXHN1LOLsanokrLv3M0bVmj2yiwBdQXw5/Gd2ukwlw5wt1ESbKzjIuaSmYBq
a/llxFlJhjig5xVWrlFOjGIxM/pbisDKxgYn/rM54a3gbGURRXhFZinuVz0U1RqR
XWDt7I/0dJWZM6RUAHVq5eo7RSrFADnitMWmoZRKooxxG34M5Jj8ger3PfKTfEMs
tQSXdjRKO+wzIKCBgfoH+bHLr4aow3lk6yyLBgn2wH0mayH36xi7NphUFgIPkA+g
J+9U4HDaLwow4REQpQb4kmrcPuXiA7XLdxb5Pw4wb0RLoKZNR3ISclizgRJPSqqR
Wzt/EMg55KCnA0cRa/NMrS1uk+7+CNcHd5KfHKZ22XBt4+Q1wC8DE2HSzX5aazJx
k/+lyK0eNTmAScEwcsGQ0CxXk2/dfHtPZz0zENSC7dYC215qelWo2uTW3cka+c0E
ePbO4NjO1tWpRD14OZA8rv8l96pkfp08KAHJrOVL/+KpQ1aeGe5CQonS/v/NeqIF
qXRiZtlJd5S/tIjSvX3pv4p2aN2P42agrA689vakF0GDEzw1ial42Syi0v9NjVfY
3tk5cxzT6w86SC6o8ZyrNn+tYmKjeI7p637Ehhb7jgctKPRq3bN7lCv+qphN7Wm6
aThdiN65/iDtx9jw1HSz+asveipzZjKKvggg3EyV8QlqbezxQK06FIYHd620AzPs
b5NCuQrEvZ2AYLFQGoidseveDG8u7hWQSHO8HsUqsVqf53n+4qQye9f2yCQkYUM8
cgx40aJhUtv76KolJ5waRnFTJeLMYHt9iU4b2MudRQSapV+266r0j0kIO8RAlE4n
FC5WHqvIL3CLpronbhmVoLocGKppMtY4DnCputEZnTe7ZJYeON4oAHtML0P2LJmX
7UcOBGGSfQKcv5zo8fuGwLqau9M5pjBeO1b/otNngHQWikKG3TP6JsbWGM2BFkxg
NTztMwUyRSbopgVsowgmi6uPP6Itp2h3EEU/OmfXQIszcEBhS7uZ/p/1eWE1f9Ci
Sm0i+Re+MkLClyb1kRdfftPwXwehOwluopJpZIhaPo7vZhSbaAcii9YG5rljpCw9
zrfjRG6SErUjvczkDMktQJVn/Eob6IzI7fb0lpZSineMoN5EJyQ1mbN2BH75flJO
n6AlzvsUAebNh3fnxIJ+qTNsuXi8UQogeaFhoMvBQg0IeQnZLnrGgOgxN7Tk8PKd
qkph/fiqBywQ88R7m53kDC95OB91NmWnFnaDq3DVCRv76IYu6lcANol6P41Cuj1H
oiRdqHtjxIdRqyAB1JR2QGNYWZ//tT7WdG099HvLfJ7P/LF4QImV4iM/Nq7au13A
5ilbiNC/XxcORMW1NY20ZDaepTxXvscK4Li8sfiOeYG42b32MH836Kx/cTPlAWPN
h7VQ2bmNTkA4oNR/vvuK4ZTB+JDNi/3pRWcorYWYW8Yd2k9F1EJH1kHDabc2BBAs
g3sDZYsQlN2OoYCbZk+Y5/cYtYeznJF0WTKkc+NrY/eoXbUCapOP1GA5CTNYV6e3
f0D2DayMLjzZhK6HsTO2mXtkzg1e5wAS8d1h4FXNLAcRmNfRJ6uiSXqA5xwzHkHL
pVUeo2f9yQomK3fArtiPlCKOqfgsEILGEVUdmfKuRrydJL0E7/vv/IAiVlJDfiB7
gN6oRhhBXl20xlbP8J9IWBFuQmL2arx9tjZZ5VhDPwB4+IVWlkiC7DVR9c9F/2vV
6N4rVb9OMCo46/ZyFw5AWkMimEX80RbGg91i69lQbDcBD1bQuT/oOJj7c3IDE/Vu
+TEUMGuM1Mzw+CofSn6jzWYzNlfQbZzUMCxsRTKng/r7uwDktkGbhiJ5GKczT6zN
Yn3BT2Lxd7eJxtQsf6pVZO/YBPuVCcuQ8pAH5eGFMegOawsVSDa2K+yTJrQ/MDBS
wnWAiTEO2xvNKoPzxwL8yoeNATl3GxaCDPw0l1ubw34yNHHF5keEd5gK+K2w5SxN
Z5eY+XkaTSSuFrfsXo5NzD4L352qCJ9sdDvh9VuUQ2kirRq3vWQh3zo63+khVVcr
3eI5MZeUeGOWIZmFPf5TqzlArRlcWmDFFMfg++wtYFolNxOqMXuFpTc83wQmHB90
cP0AtpdTK8Y0dVMkXW5gTpr5xaDPQ2g0NFxcUFfdVnFcEwewSjoWjbrr5uMxwf+3
bx05yc7/7D7Dq8pXADqe5dqG5jnCboxOa56shLKKpBmiQ27ZlWXk/7jEUd3Ocdj1
78/B04DspygfHQFqqRf7RPLmClWE0xtIzRnMBKhihVFck2Qat3WdDng29wxWC9L6
84MmsZRnzDXG/aQ1plw0h/+rL2IcR0F0TaBWfhguRINbFLUzuabOCZq55LqmnVCq
0TKog65QBDME8dARmw8A2tu9RRLG01YugpgZ5EiGRHB0vuNeDAt2ANqGw6+kXnYN
Q3sHKAaA4tj4ys63TuNKli9pr1l9Vqqxl6ifzMW/VcON4tTRP8QJCuB0oOFR7ZZK
gVIdKiEbkR7yH2M+8F0WaQwRNEGc+ALZkfUIscrJaeKoeT5iiomdlHG4J7W1TGPo
KvF1cQ6cDtVGpjuok6PfHuh1UEPo9ZSDHiCo2Oy8yjuw/4TbvVMk87FvwAhimQBa
Dg2Kjtrp5twswINurMMiqKxNWTobILdU9bg0kpmrk0xA/A8KdbzLY6rIRzfU4r00
Lra0L7xrvavoU+sGlV/iUOZXLY96TFZyrf9Bvo4Ra1EfrE+yA4PDkv/fbxqvC4Qh
piDH2cKM5lFCEnJY0XUlTE2UiT7BZd2wT/B2J+zdeSOEWedxN7AT/QB+dXG71mhH
xzFoZFEq2GMHxB4ZGZhZGPb6HzdazRTpcm7lAvzXlQThCynNIFJB7cCLblSgMw1e
958GiQ4lDKccM3EZ4dMMYObJ2ZDhlSks63JHZOOZvYiJFyF7xvhFmRJVk7p3V1Lo
s/DUsMa1z+h1rtb7JU+SFjytbB7NeBCvbVKyuMXAUx1WQ2OUI0GN/DTkolVnR6Pm
KuGsxonEvfjeg6H3C1ocNwutJWOQ9u2Abub1VHOTaXbxExTNcGpR3N4Jc36km+Ao
2G9dslaXLDm/A7DWeR+FXGpsFJ2sU8mErFjb4qgAdCp1cm7VCpRqqFqr464wVenF
x3sOZTtxYL3zNNOFYPh1CZk3bXvdMhgVJ91x7Nwn5nQRM0E9mxfFy1Sx/FiMPNzp
Uhjr+bBSfFRLu+jgbxadc5zmH9bcavy4ZEGrZZjvBWU0j1sBi7iFj3OXYYoigN67
UJDWxK4KKRjirczN82woZDeLdyBzgs4FqJF2TazD5ZKuPNaKGqxlVwnFdWG1BHGO
LXChqVNJyzEcq6zEj58qVFWrr+LWJNI1kh01gcrw7xZ0k/MfjA2I8E6trwpOIEmC
qSUS/TbUvD2CpjYDibamq5PuP/EmeAm1/KzJe5+9BsCN9AMzULyPqpgoSFvmo54Q
FY2kZeXLB0QS+995XzQtYAKbzo7FwCjR68pumdKQfD9S3ooX1E3G7EgIy07dI6+7
NPRAPmWuQFVzjK5oSeh2wYdLpAEhiu/kLwX5AhKRrWOBgVHAnjo9igqflwWUMi6z
FmJU56MRyMA5qh3hvaE4gtOXqwTnLYgFR6KgegEiKh/7R4Rxyzc/qWgkrM8hi9e0
+Mj0qRtP2h9Pew8HDNXOUxJ5K7MRTb3b7bj2yT8AQh6rFu/sJ8AwXzkxaEOCzz1H
P0PhQMwUzPVvTfnLWBXghRwHd+ucJzp9r3VoaQKZyXN664obXG6uPhHd51RmUXfm
2on9SB36vd887NxO5/5HDKflX0Ez8jEazXyM+YLD7idIuj1bqkz21gl7UBTDMUrw
Zk+AvGr6WbH4eceaAabnWdNVRcAxxc8FEQQhksQpRKRaLSjUohd3BU24J6yN+NJA
XR102f+vmlPK0AOwGM2GVRyy3aMgrbu4u4vpl0A9y4WSDLFW0Dorz9cplvFlK2qE
HZELw9Hx5qafoYkllEmoI/bSHjcq8HYWduAkkd5WBqnZ6HXbldSmNWfX67RnsYcH
wHYgjKGVVexiYGClfnxL7a2BSLr+NlLQBSNPfuGmd3cI5ZUUO3aZHXyrQ2A/OVAd
uv4iDQA2zQQPlFcCPSjOVbYCai0RbTP4k927kzIgvgDfYT4np72UAl7PqxiLu/6x
ZuOuq/RRi33p+JBMKpG3STxF3Y9TTaglkIBW9wE2En4BKVC6oijMS/iZsBktgHYd
23lGaxX4IDMgldXqdcUdYUbm34Y9QOkri0496VWToZk0KSX3pvmMVt/qKp9KU9Lg
RKDGFMEeqbxv93eRAPP00tv0sIZOqXu/PqX6DKHIjNBdlBeGr9HFiNyyh2s9QR3S
P1nNulrc2b8RatOGDRC4doe0RSl+/f6QrPseJe0JXs/lk4+EBGu6kI0VKeXJzJtM
Lw7q/nHWZO9mS0DEuXlK/dKjCNql5WUKan3JEnE4qBfeXIw36OZanfZwxKLYuGVF
OhkWzjBtav8lljpIfibDFQSBHkk0g6HrvQlhUvoxztO1e7cf+1j+nBmJ9gJyzqAb
9jaBtLx79hrY9KSlKRsnLTooBSOSzf7hldsr0fOpuuRFHoupAcamD9HvBBM1B+Hy
Rqjf4Au5XfVb0bo+LAZGQMVjT2QL1HH49CtBVE7TpYcNCVQseKQyaju9yNuniGJQ
h+Vsxe+gL84T1KeG9/lybvZfFOGOGlwTFmdc0H5V3l2+Da7rrzOhgg6wzmRpOt4I
OK6Sqyg0BgXSrdb5sr0AYoW69WnllQNkjhPtAxmhpdIMN6jwQgW+38ckZig61rN+
KDZ8dJFJt7iGLtCvbSOVwa6Z72ef2F+7tpNk0RVlBRnaQ9FUxSkcLWSuGnZz5sQc
tt2BpIKjqLU1wUBZoFu9bX4/Af06WMO/t1w7xwovDJUhfyQ9of7/rm22N/Tv94Tf
DXYj0Z8n/1kbznIU8Q/XZYfaYcwzinL9ySdo2uT4PWFr6m5WCXCXp0AfFvcJlMhL
6yOQTh54scxk7tjJDmFVVtMydswGxS7zPk13UqCDv8VjR+KYIjbXw3fYhhKiYezG
YXSOXLn8R9yywu1Y4wq2atpAKvJhcV37ntfscDoxbP0JLGma/8S7o7I5CitLSK2E
yFIEsakLk+1zONTiHhctbrmFVrzXKDneRWoxdG/GxhXTgt2QhFv0h18ltA3tOb8L
RWJkZDKEqoXL9/YY9SKm73LvyOgaP3sygxI2NG6onrOWyu0tGZaqCqor5I+0sYVF
11an4oXWMjfQmSzYPbC1NOB15wb+9VbFB3O3gVYM+LMZu5sVv8anyx34E39ARheJ
p0nK0azT+2J4uUmsFoHZTi/wmMRrBAMlkYoUrupkWcjSP2sdoygYKXtD4yLZ24Gz
LGeII2TfZ1yCNwL8W1nM+L94mJ6Y9XwilWmxUyh2Af5sdnvzeABiaIvIKP0bdc3B
NzzVNly3sefBMuY2wFBF5b4NXD8pEdRnXOLM1eYBjHxMQ0Qb7atLSDrd+5uYWUSb
A9k4wpCX0uU+S5iTHB699LB0uI7TRiQcWN3a1AFaUXY4WgWzXaoT8PjNlG4xqSxJ
0fgHevRUs1BHldvap/RmctzPb+jNdr2KXLuiuCdrs5uCTie8LcwFV6MZ1qXC+fMq
r2osn0ukxqq05uKI3CSfFqpmpBBzRBOc6gRXwhozMvTUiktsOdQvQiU74ORBy/4F
8uYChutXmjgp4rNF23tZqdYZNNEcmtVEgTBoDhG+e5Mrr/4nfsDLrCm4jyDSybOM
byr3vzEe7LX40mgA96NBFYO0zphkoxi4kXTpYJOIaOpiammWVj70TTUhKZxQ26up
1ztKBDnx4odYhj5ZPbgi65sZpsgAhCEsSApqEEC1XKlQX/F8aeaywSdxYFtHSJfK
O1cBBoKAqdD1J5OhXPEZu0Lofh3W3NZZRnRIlYraWqL/rHefYDBFJJaQcyOJYeor
JEy3uXLN5b+DHQfWX6wp/d+j76TCJUcygXagd4/uHfGdn2vFySpkrg356luUWArK
sKdhf++JDCDqZH7NdlG2OPvXDHVuzztySmTClZPk4kQ9/1dp9YBPbGtqT1M9MIP9
+t17lT3pwG7BjdZ+WZotPzjr9h7Eh6Y0ne8v/gKQRhITVHmJcm6UdnSdi7I0gxok
Jb02i4HFx2fodWa3sNFNu7+p5jgV8PvgSSizJm8voD4/Bu8aYTN/WnXEqkMjkrPW
Wc61Maldnmn+2ZeN+2m0qH/tAKA1UUBv2VnB8w/CvpfVU/bUcaS1UpYTxorK8A5P
a68OgxVm3MaAbnyPeWPeizHGLQuQ6kJdo8BeFn9Inre602iClXbalTWomFoJvQva
Twye/3OZDbDRybcbJmAMKjHR3P3oZX2jBdjg9TJkKN90kuEMKsyuqC9oaTWdtexj
8PkTQC9nmtwBdvtg/dwRdQr0xRNw/Qa8psTw5ZaA80aU4O6/Y5PK4N3ZgzZBMii8
X9d0V+qciJAH27kslpN+fQ+6C3w8w+QYDsKImR2Tahg5bdyN2KB0pCp4GVkW7BJX
K4cBiyKIW/zOc4h894czcotxDEDIwktSSKgW8TuQieLjsFZ6Kc3esLQ1qxea09qP
IumPl5Uh0LJ4wTXuBJNayowMeMCYEyV9OIAIpcqWCo2rWq8qD3eaHlin2tafPuon
7vwvAHwz7/P3g8gqqhDjf9OaycNjVHdqTLlriBZpVhOt2zhNQhJrAjoPhrDl8bnr
6q2uX9dNH/QjeDzP2Vq5/PA09UPKad3BaqmJJkiVSVnoGbzli4KjyZjKzq1ZDHrD
0tXP1Pz+N78+xoQQJqIM43/MgQYJerp29Xjx/y6P2jMXZWjsxJyyQD9Knk9q8OG2
OaW1VWKtnf/DEQCStLSj6pvWmcFz+fYyP6OP89FymWcKF8lnEeznALMoIiDJ91k9
YD87YNZGHRtdNrclHcB+avtarhVeeMoxF2ccztIEObN6iivxML+BOiHC5InPjYOe
tJFJYGmm17xqF7+CuFZa11oZVKVAJf6A+qigXl7G5+KdMHovBt0EVcZsyEBaOFIu
6WZBWyouU0Xfx7oeYjjhveVvFZ7dKTIB+94Ly5vVL18KbwqojMsWLGvHDLYar9tJ
kN0gqnNjWikRy9kUAmvVjEryrwaqw0IosZJxHsPezjn9qSaYTmjfkZGlZXuGkc9x
RxXoHm5KPYQLH3eRNwTrOdw7+te3CdjYuBpLFMp7vKW+cQrHsy1k5lkfwNUG3cpw
b0ksdaXANBBdLZh9zE+yx/JpCIXdTwl3nM8pI4aH32UGXo/KRMVeP067fxbqQDed
fR2+IC8G4mmqQi8kamCYmCbDV17qVzhw66zePHvX3AXwostrNqkog/wxgZQG2BgM
heQp1h3mcr3c0vXOdzQ8HpHKg90xz9m18928hwDe3rSNFPgxIdPEJXcehfor1cgZ
ktIRGfJgqO1PuDu6SUbybO3Fe6OFhzumchYLHqbhn163BDEQy5Vuxc0mnSVqev4T
T0rEHXIBvzl0i15zqqSc3h82t7v5q0AnDF+x2qtqo3oQ7wbQeJGV7y7cK8ItBpfy
HikSxhM+QmXSwlwRMxf4S+1U4yfP5tBnznMjoDRlHxh70zIki9fi/twUZs2yIxBT
4DasR6I6rwqbL9h8MPe7IZ6ls1DxqEs5IJ0kMrHwcFBzVvY4LCg71mf+cRzYkyPL
XXEb3YkYLBUdambXE9f/Is+eZQ86EWwKHW5W9nb8pOMY3DC6gMepwId5X27cIMI2
K7bW0JSMlNrymwGTmq+YtnyVVkYDW7f8lISzZzcFAh3hl7mt0AVhkEoVzkIod5pY
geNRqWot4lv2Hku8Fbv/I2/OSTMoummE/K7JkxNpOXOFeGNWdGYtVjV6MHv9+MdC
q2WFgS9TMdJ+nJUPcrfgMTMzBaoJEOU83opLmtsZdfiREfXdkzvBXalwYQcu3J+j
gCUL7Po2PRW6QnNjF4FSuBO/hVWxy+SrrNiScy82Xv5mh9AIWJB51sh582qClbZw
XaF/MVtn57UyzqzTrMG4JY6HdLa7VrFjxAYkgUelzFvmkCPUB2k4MwVWMRekAegC
cTBGe2hx8qj5o5a2C3zlA0NbpXDso2grWzrSJwF25QkQtPksQm22a/XGdtXu6teC
YEDdQS/wIcQQmJicb0vH+sFYGtxDW/E6IWhA6a5+NXOIS8Rl/HFnKMVmcwRElcOl
enfa2LGKfomMRQjLflxKKbP3J2LSsuxawnb/FIm9SXm4paWBXen5kEMRvrp8Y3kT
llZ1sYjQGOVx2/mSElnU9IRFhV6ZCGLBgOifOvzJda2UQJ3d9yh+YXcFASFt5PSm
+VvHlGtoK2iFxGS71M+FmFeYPGJPdzZmkAa6hadKLIpMNgLTYRa5GLQ3aSKvJVnX
cWFjfG84I11lqXzqFYFge+2RivNKIQI/NXPZ1KwihqbnhcrzOzQJYagrnEKhuvFU
Zmd8vbvbFhdncA6HdoEw9Q6z/qReGDHeQ7+lhlvw+r+k4QVuCqpdfsS+92/ix8Gq
aM8LXfDWPasZeLaSKdjkI9kC4iNwe9IPFURBRjuwv7MvTxY6WiCETaVvJmJN8+3p
gicBbrm21IAhKZiPKVRyqt020p8oLLoZvynPi5v/cC08eQ6hTJCWPdv7Y0Z8OhOZ
iItnEb8yUSJDhR/gWkKyqkRheiGdFV/xjTX4Lm+rYpLBqGNaRAILepu7EWFbTy6k
oWGFqQSSJF2QXEFJYcPaOqMBiM8XHysaYrBPZXnFxr8mfGpe1+iiWUH3VqRyqQCZ
l3qxhbfUVohOVH3yceJTi2K4KSsU1cSSC2GaOuy0Z93PrY1dvCPblyj2I2Xe+4Yn
oXZRwDEjjKZnraVr2PErNlPsbELJqR7gRZQ3asjXMne8CfrYYLKk17xXVSxnOb9P
Yr6OaNFRynlAr4yT40EgurVnobb2HkhsRvYBqasW+7IVhYU7boMbZdlOiqFxEVsE
FoPL0SZVcYi/udZyBzzn71vRGbfWCdvYGNIEBBG5xytU+IoKKpDlbcPg3UfA8/JI
7mB1qwrSKfIrgje7WRJFF8alC1lhbyIDSB8zRY9XvZmpjvaIcBG+zn/xbAUT4yKA
jWm2q5Zk1RA5RkATRTglQXcuxI+1lot1dp8eFhq0nCVnW0n3vFKtfp7oRt3On3uy
Hka1ktjTXay9lpVz0lzoRuww2vzV1LcdoDmCITAViKqDcA6B5vBuGT2PTcDUIhVH
FTAcYoCWB/XDz1EhIL3Bwd+g/hx6ShznUjPl5ZOSvF3XJuVrMgW+WUdiJM3NjBpG
hU0DqsrT1++yeaE95qK5j1ROB5BKrtG9YxS+LR4r3lGSJBtB2f5c2yw54lkZP+Ge
1DWOpGPhLhSD2NJBbRraYiOSbRL7/J4jfYO+v5s5PZDlngGn+BexENRAJ1/7FJhx
nfOZFmYDiOBdRrD7G9ZE1LTJl5amCW272HWhnyfyRi6ZUgqtiEefUDNBl150jpyv
q7Sdq4+/3/QP2lybrY8hAnVW9/l8bjLdT5BjhBROtx0ioAZh80D5u6tlpyrRRNfy
oP4HCXMzrD/601E28rglp6W3KP+sB9ui0o6w1Fq9xtksmo3bLL11R8TXeW/PF9i5
7gBwyiHMH7GjHmUSvBKs3smXPjSwQKwRVg+Bu7w923g3lxbtcQ2YzoehGw93x2np
DLl5k/KkspWqdvKnlEzDe+zA9+CvIJAm2JlTvO/mVqsfqZNzwEXPSuGtDNX52/up
QZCBgXSyE44QI+v7GAhuX35FcCylXOUFhAPtTRzAFDuedEwg81xMIey4SkENt5GT
KBaXMiXMwbAm2emS9iEi0jbF/wYuJ7VHE68n5RwoclYqYwrp4F64UZasinraeJrA
SWfer+1ROuUcIV/xM2Gu/ZvDR6zB+5lXIJpI38X6oyrNyHjBtK39nw3V2ofMg3G2
eRQ3tfx/1G5iyUjEfJ5wQAiVwcYO3lJFVbAhjo4t6c3ZLJCbd9UVijkbLqR9geOr
tBp7Udcq4NJcg3FltPpViur1lA1BcYgbmlbFamdRis7d8BDqQt2+tZUxjDKJMUzj
4oJ+QOaMR3MEd4OdAbAHtyFhRLfMRFuL+fUIpWxfNJgDNakiw3eN6GZ46xBZ1GwR
+tfxVRNrlRQxBdDn7bxz+mOu2QbkUMTDfeCKE3S99lCYGLookNClY3XDHaxroCGj
0pCoX0nZw1VXwbG4wv8lEYrMREYMO2OvUKVD870WaHZrqUYQ2dl79cthvl70jzmZ
7lFymw1mgDgcgaFAxsvCJwsdPDnf3VvD6UNv9jiwT2NBf+04Pz2C/lWSR2UBW5t2
XMygkLt4wu2M97M4QX1LXnw5lVdoueFg842Fs+dqa2ysakVoBJYqASabXbci1kbC
b0cyhD4pJLGp7q8Uyg/Y3+p3nNt4q1u1X52D3NvLeToM+qNc+yfXkZS9tLhNw6tS
sedp+RNVYutxKDFdI2ODA+rROJMHUrGUMZeS/cXLThiDzH+VceYLqeKbxNEdHowN
Qv6R9cvfqKT7OALrfoHvx9C8mXy1IfvD+UKMe99ywI7rCBZERwIBFGnznlcz3K2O
yoIznOvg6iwQ461dTiyVWO3Oz7Ao3xDYAEw8V+HDl7krdy7kX5fgoRh/dnnyVHPA
/nOtKz8ly4N+k23yQVKKza0Qmxi2cFDz27GvIoQj3IUEfzK1bJLzv6yPP9g9MT/s
7ByIvj4ALqheIOKwzl4HZXLCkj4tNX+h2pSHfthntLQCB7EUGUuc1kLurkY9Mi66
C4Nuv3IASWDNd6fDSC3+eTrdG1RUUTte1t4zNoTL8LM/VpP/nxes9r/OlISos8gg
a+FcLivgKcz9CPh9r54+2BKtzm+PlpQX6zXcct6dVbJhtz1SOZihbRnEIx6O82ki
t2BSeXh9VjVefuyIrgS6aahCi1m7d8Jm7pPaq9Tlj9p5gMY/MhHmuVQcVmCGKEYx
5F74003/O758gc/Dr9uPvqW6C8IPEC5nOZBHrbBtAkh41ARJePdr9rmd6TprYN/F
0K2GzGslDZiZCj99K/HxHbkQ7nVR3uy8zIWylJXagRQvti/Onqb6iM3EUs1Mbs5i
spU0Hzuu7fajwoSdJHhI9i0uKBjNO0Gv9V3ief+DjJvhoi9ZCO9GEX62tkN26W5c
E+B3/Iq4K1ATZVr82UkguSn5Rdv9xDqh7DVAZEUmwlnSn4a6xvWT45owuDtKpk4s
OzezsQCs2q16ZCakc+FRRfV0jMhh3BkNWY+awkcQtn5dlXRYDN50ULgAL8FBQf+b
jqC5OzZc9izb7cmMOTJok+sHJpnimFdND/CsZ/rhv6QCt4jsa+JyAdiFFnWLnhBE
51V6VSLbt35d8agxkahyX314hEuS6fbLZcFr2g2dpat4ibZbYPJPgT/EsIuD0dS5
Ss9Qt1hrtiLLgalN/4Gax8w70vdxK4NmQcohXYp6m3dhjSbpbnMe9+AWfxKvUdem
leRyhxV22Z/Ds+bXdK/ydDdVi5mK+PvRHvC/BHg5+vJCh0FZzXgza5xyez0AWHg+
SvFGl0AGAfJUIgdrG7mTSQ2qZLiJYyJFZeP/s39d81BtdnZ4unULFN0DXe/8EiOH
xlOcFITou0+Ug0pGxTb9Uyxyq0/rc2Ki1y8wftDgve2w9Y0p77IS+8nsPvJG0qiO
wJlxYRcVOB1TJX1ciOm1BfvhfmgoqUb55Ns4nqWWttCBuJDrRfS+my+RJjpQyZo1
L3GevkhDNcx8WWPLDfgRMBbtEbGFUupCk9wMjpjtwnK9ufGHnawdSNLiJNJEXiPA
rjHCav5gJW+yxXE5rLX22eE0uPujzN58c++s5cJkerEWCy0GhHplyiY+H6uWS2Oa
uNI0RiUm6S3bBoUAiWf3UwWTcS4Ul4hHqDjUcY9P/UdHHr3++B5iFy6/foDodC0G
SzKvYWMiFBBpFeSSwe26ES3dC5caWv0g4dDQIDoaijlUHz3yOkYWHKRZpdLhqH6q
Oiuc0Yv2ufPGjdiKJMGv18C0BtSHgYx/+pr0QLHBXX1S4ssy4ozMi4GBCWY24aab
gmL95M5UB8Zt8JvUbb1U4kJiPAVuMAnV9XbLaBJfInYTasapZEa0rYCSfPSVWDC2
DOH2d8QFzLohgJmXce/pPELJ/vxO5ivi0lh5804lESalRHBQigfzbcFlTRNxMHC8
ud7ptL4PAXwuLebfcsSslNYYbocVxOyE9lnMNnBIHTCLGzLbw3uq7alXDQ7EkVpr
lNvsrYOV/R6lVReXI6vUicJuXI28VArozMeCHsoW6VpCp5s3L9Hqhx2rwAZEIiPG
rHUByXvKs/n73JuuDLBXKx1ok0VULpUKxdXmyyDr9bfhOy+WN9mnZNyqEoAzZREk
YyKkD7pcCZoZqgqrhY7VTLz5A/c9hnO0vMaPzssGF0NIZCpP5pX5XYTgjyiqx7Zg
6iv51dBUO5FT/orLLa2cLEFp8ZNk7jXtyAXKKVaTZEu5ci1Sq3UoESKpETgs3veN
6CFVJoZj5pIOfAO2YwR+SrBIq/rqwZJMIPDgT1k3WvAw0/fZELJaQy6BJWWrtf5t
oyXHilbtjUrrhLRBd9TQV314fAv74SWh0v9yhDNqhiA0n5PkVFmDbdXiIQNBwaTt
BNZqFZ8nWmecbcezdXPtbA352KGgdkzL9dSMe6ULrbHoymJudZgF8u7o4pEU3zvX
bmgj7Dag1O+dntaBrs4aBN97C7nRplHgQhHWdjLrZvoA9b5RtZ0Z/e/WOkQjUEzc
JnZ+yWa0TFelOmMm0N3THcXqdaDxZtYu2t/EgpBWb4ehtlbO5tY+7WMiODRQwdca
+RTbL9BGtURRDJ17OO39BS1D9V2ZQTghFFa2QmnOTK82Jm4WAhRyJ5AxiJkFGqDH
RONfobdch6tEuZafFOkvSKz4FV2tJxWaIXq8nfNASTn8/W317SSiNy9HDor1i4W3
4PlMaAFH0QBwVCv/opW+LyS6uREAIfQc8sGnrOtMebvylsiH+nLCkY/Ujjqn51v7
O/6Q859eY5Dj42YvcPULRDAbY1YErJ4ZrIRp/unkium2lu2OUpweUpaKz11ELfoL
9DOfc+pZF/UTsC+IR5xEhHt3F4q39MAYDTpHjKz4GzYELEY4yLsI3W5OnoYlp6zb
MnHFtHh4E+19r4KH37E6UEWgtFEr/fGaMQpojVf68P/LrYxbCVU7xKyVY/0Ybiyk
Ts4/pztboU+tXm7AwyTCChQZ66RDJ9FliRh6NL+3KCOnblC1pQUdcBQmFLzB7VNV
CoUEKkIgFP/U7FDRoV0X9fAu9/ZScgIgYY9zPpP4I6MCX3Pa8bPfLlit6jfQRogO
CF5K5/P9wlgBJcarthnVGs3PJ9stUBqRePELsGCnrXsZC2YZ5osSEyhfD97IdG8f
UUrRTy/jgex9kxXswaTWmI5rYdhDHRJzW95dzkPlC1k5lmDzgyvLkAZfixO+bi0A
S85bLJvtqF143Av7Xips5iO/+KFocIq9Y+S/3O6pQ/Jl6phw3G82DNiNzUq1oa/Y
o6U3lfQVP0c0cLHd6l4zMkXipZSGNEBd9r+D1dYjUq8YLaQlL3ORyKE+zmoa+2WQ
u6WGiwweKdXRvoaI0O/EmKn2+h80oGTi31R5Xo/c809t8nRu8XOd/fCMCFAzyHcd
cV7iXDmSFFE2DgktH/XPLkwZw9OVchEFREjgFzBq/E3eVv+Bh+sOtcnTCNZA8kQ6
OxIpVQRBMo9TsQcUPIx6mPro4OikTVUnCjnoZlWQu9vG2DszQM5v4Gf2BXmvXoNz
paIfvOC6LWwQgkRWT+VsVaPX2RDaMzwRC1bGzEPf+jKwcqJAwZtGIde6EZ6eJAAA
w6oEYwIzuCaxjf5Sd2RtJTmhXyeObgWnNWtGPv3wGIpRVmv/mD7BYN3+P0eSpWd8
NyKaWaIDh9QLLQdEBzxlBvZfDJieKpMIVPQUWi4CRHbzG9NHX94Mjpztm4px1iRb
DbCjS97Hsnc6S9KlZuVgngxSpyTSQwX1w8bm52xeeusYD93hVJBCPjlBh4fVwxFZ
2+lIsKJvTsKZHCFqwfbmBZw0EpV5UmT8yR9dCwS32vbEBR4IVgs19YYztLrNV1QY
CPQVaDAljBLj5ArwsM78gsBBZIXNrgOCxZtq4huxg6LfAGnd+YgL58MfWix24BDr
mt6SY5hZUQhadrpqVCfnSmhbiCBAv5L31dPHgjfE156V9m3WCojqsn58yWXxOmyK
onYT0JTsHZ14TzC/zetfUoKEXgnuOtrFEfNb8zDLddiI+QOUBKoDt2XTgi2hz95X
KlKaYGB5+Cb9mD9LmUZjQ+F6c1aTMoWNFJ+y2x0R0JTmi7oF5bSbOA2hM1VqxSjD
sLR+3qX1+GA4NYT+fVjWK8GCiEiIiar8p+cLYL4uIXUavJ0Q7Uq+GTTTmCvASknO
aDr+oYmA84M/RPb5cssf8MYJa1IyeJGU0hWRXFCnnsYYfF0FR4J4MjR4TfHCv9eh
+K/a9fC13PlzdLTsam1CeGGE3hBXdxxDUIseBnTR2J6OAFbIy6QEEIE4E8jpCu8I
UFOjiqkohwWqky7D9ruIrkrY4qe8j9MCJ3DHvYFTjWt4ZY5xhOTs0j/GFXRYxAMd
AwIIdHT8Hic7LAvS5lL7P4s+9un23ImmjQwzwyp/0JZuuhpnz+psmtttq78aUADe
HzYx5IRrJbPcqoNuVdN0N9NHaggjA1vG+pDILaTmwICrnMInvVCRkGlDSj3SQQbe
u3d4QPgVy8PjHVVc0SMuvAhSw3PfaXUf27Bn48WVCtMOurrnzAiM/Deim9e0p4jb
WlOgkCP9KzNgGi0weogu+r+SWN8aHH6zH3ddi9Iw1fz36GnEIOFq61L3UTq96kNw
ZDOorsyCOGXZIoaWxiBjJbgPTvfI36MKevksDA4tg4uDkxfRV2Tl8AVuj3c2SU2W
X4GknIcfXNYE0Zb/b3SzyWr4CkVc0kiRqsPkPk35ca1Kp8VSZuWRmWknumlww5I1
v8+Fq0exOiHHhgPAfFGlR6XP4b5ETekdNNCUoA+UNSfYNPMa8HzgfQXiFnFIBk5P
W/c8pBajRfRUwM0PZystZZv59szb8PfdKpIu7hJsfz8fUjXKTZ+pTnBWURLVUhca
7LnJO0j8yNcgOOUO0QjXWJls2ln6J6UHJ7s53XYeXthOyYqZ3ny53e7e2xqfytDP
MqqetmQo3o1HMlQLGbk5eS9TXAQAZDR0O4CuUYRsc9wzEWFWKzajLFxc1FS26mCq
hIqgKHgpru9K/UOuRXRypOx3kgYVMMe7mPJUCwdG3ySYorX2xpOE634QzDPDICGi
VDXh9EMsGmQL8OJOAwuyuPnj69HUQF2WWirkN9PnGFEZHzhkSwymqAm7ml8FuNsd
Bm+MyO2R8/2keOUTPw4tdOCYGm1bUiTT8HxXgUFITLbezrzGp4gw26Zul27o507X
YC+MH1xLDkEQx12e5z2noj8aLAGiCrIV0wh2RZtTu/3+3t4qPZv32yt4HEdWyZ5m
rOdx9k3s1VFnRRnIsuIWGc1L5v7miqc3AzWVUWQg8Pl8G1W4lyTz4hrVIVXn9hxU
FDLt4b+FFsSINKUXBLlI5twSuNuhoNTAh3IyIx1YaqDGuqv7PNBeHHtgVbAlwtQt
zxro5uNbPpyq9DjDAKRXlCV7k+zRMB+5FJl0kHSwIcooT3m51jMdR3bNpHmNnTZN
TKGJcaDw4O9zZHu6NPNz5OkpJS6GsRtiNwxjthlQeqqnr5Z0GvSDsTE4wBsStNbs
q7dhMQaCchUlncSCzTe2hhffIEZTw+A+pTB5uu23NnINKR0oDst2kW8WucUXnH9b
S+aN/+RvVn2L4TECiqOqq4GEOsbmNqbKRL8n8Ot6bT+mce3oLiMZIz+nRAeGN8Gp
fKVTtAQbNlJvCAGJM9ioKBN3H715yM9J00Qp+5ziVhBi23GHmxBRmy5HSrQU2RY9
GdPll5Pad3CgtjAgND8vaYHJS44JoeOFpoAqsU8IQMNWXnjdrGwu+zpR9MGsJ+7V
vw/482riojoIu6QNDGheM+4RCYUonzl8imZb/DrWHRvRqP3vYPwzQM6yBRg+gXZ9
eSogWmqrCLJRyfBgvAIOx4repM3GyOL7Mu4fvIwxiQv8EW5cAfIoimonGCkShPi/
xWkN2qbl5HaFtTnU/h4+SdrWuxptVIGXszwJrFuyPoPbB6u5iwzdOBSZ1fzSgIAq
cw66HUU3nBldG838trtZbmDIWpq/FUY64fdiXTvqt8SksMuotkml1jHv/zYJULR/
meJfyNijfl5MAn1glS910c7kKkQLCF8TLBPUzl6xT71xkTNTEAAGYxMhcObEbeRM
AA99J7/UgLHsyK8ZtP2PtGX2T/qANv7zLscDjSY1He4qm0tuqOQIh+wOagABrVNL
S3Mt9t6qNCIbdRtsBfSlt05rmyJm9JKisUObRnsstVjHbAnRVFhnGVVwhla9/5+c
X1a/VAzLSdGB1ItO4GdzPHxQzf23bzCRx42+nX6bRBxte2nipkTkrC27HyAoVLch
iN5IOd8QN+0M7uSSbCOAj0zDsGyNRo8sR7PMn1xDc8M0ZpoxHHLbcmOmfduicn0j
bUSHVHlcm5oGj3oO3jvgHO5p86JVXWn6VoDyXYAkCsiXyiVjJk7ea0D/xYQhRKcB
2Nu7KqzGaZ2jtfO1bZljPfUstc/arg1Y5TAWWHnEfNoGU5fRvSh+NEysBSZKjGgU
z7lfZ+F090SQH/dRxlEnmxNsIYeo6ySPa8eHcEALMsU85Hcr51/F1M351pV75WjY
Egn7dSibhCexDhkllOnc3aaYVjXbzWVrm14MASAhEOk3JdTIashyjSZmGk6rhwco
+vZRpka+AX6A199GhGeZ7c8GH7D77ssXO4hUNjh1t710gcQujizCp/OEe63+H6s0
+IOWCJoROZ7ey1A1+kfYG0GFrqXC5389V2qEUAZ3VUasYv6DWo36zv6qFWWgky7t
QQYz9sg7GN81wf9hxY0CQdZC/Mg9CrKT/Z5cWzF/aFHh2wje1rAgDdxLAzGHvpDD
sjJINLZAGhkgce7HA6O/XqAzn76qqJBnqQMrUHLKHAIGqKXnhsyGDeKpWbcttGIM
oNYYtjm4ecZVF0hHNIEXXievTNgzODVDKb+xkA0nClq5RKOF+f4/67tePZ+TRM1S
mNodh/LI74TO9AJWjB9wpMadZPI/mTlAZZ757vcQm05rfGv+coQGzgZg83lLAEW1
h0EeE33NrjGnu/47u/BMvvB93Ugq+wgHyCiXgEK6xaRZDv8wpjCviMONhSXU5DJp
sPmsqlDuwlbZaxdtt2RNVSZgv9z0v9lFoyNwML23m4WGk820XTArp+L9dyJWaOQ3
lc19B5ZolayqUxUQcIvzKzJCtI2NKxXsE72PYntUevrM1Ajo1dPWymQMQcijospF
k9IN+rUDzeCJ8x6Gs0G6S1RSR5UVo+biv6nIlTOEKn5DumOIfEZS9cry4a2FnhsL
fTDGTAWhJ4ZL9dIuzb+ZF33LOffP//7005kFr/u2bM/5lbQVF2ZnWoTbpJC/W3M9
FOm8G60OmMcfNERFM8nF7jSD8Ymt1XFNlt8LbrC9B6brgDJDXjS7V+hGxRH1UhMS
OU7aPQiMMUtqTXoQ/Gf5B1jJUnzL0pERSpXKrjyMBo104fgCVkaTR2LkheW5Wp8/
tKVr6v3AIqzvYnKncfMpSkav2lOUdtZzUly2fIXlK8+njpwywVMVgSxp5B593gMt
+KYoLyAF+xOGylYiB2pifEfm9QxtRf03UUmL1vVEGQP3gbzd5kZzQO1OqDqDRo/h
EsRaPLKYKo6xPfP/KQlT2PoqlR02Vf1UGZ9xdCm56xcgE1eeXVEWmpRY1EZ9HSmG
QiFtvk246Tpw9ZG86+6avgHIRUCIhsQacL35saDy6fCTIfgLIFjwjw/LloNBaMUY
9cehxBXA5ryQ7rlg5H+JKmSuag9H054k3T3W4Rkqd1FYiQa4LSYGFb4t2wUHoKDP
L5ozXiZOsNl6yfb7XOPchzXJX2msNzTalIAw4fqkQBl2ii3bWX9L2g4IZxAjkBqb
jt06GhfrDa+ET3pjUZwk7Ph24fKUOTESkZS17XqoFSmG87TSFsO0WLlrkTGsdRSi
k1ygp++KuhnL48s0GQMyOIRu3/4yYaU9C9Wy+j7TmBm9EKSWlO+ubLoJ0zFu8qqb
veewlprkSrXHkXS4xZzfB+PxRDAddyHFgG5FD/deMsCbTSrz8r6COKc3oO1P4VMY
FaH+sv7IFB4H+8HywP/h3Cyw1jLEAR+UVOvAGqQX+3YnSr0WD/LyUhhXiyHgSWOj
sO6ffayrFSP6Cu8PIQksiSzN1n+9EBwpsrPT4YW7iY2aX/GKqog17fZ18eb8PHDp
f4Cp/FuPq5yV5FUU0YGv5juQzYyou2HWioxhgcMoSS9PuRZr8/00qXvLEQ4qOxby
fe+44NFa1tGbwsr8LFULFflWpHMHt980DRgtiKbPm5IFqB5niE7WKlwStuyiahfK
5nZ5zkMygXsdysZ3G55TRvSCTwRjsXKNW0A+0RsUOcd5xcpoJFL3Sv69DyZRTjtJ
JrBDdyKPeqH7dMepTK7BRa4LFfJxfjnTj8gBb4hTzq2Ya8dN6y4nKqMdGVrmCoN0
WBKTiv1GEQW2bFGq/jBE+mE9Cn++IeH/rVOBn6HGrZbAfskT9UMPaB9OgI/JcS+w
WBI5jNiuJUC6Y+yyYU/U9lH99gL/wj8DvAJElkEytpS9nJJaqcNGaaCl5VA9ws4P
fPuBRBjjuEr3BuNLYr2Uz1Z4PWeR0oJO7dPXThrR9JU9naKiXAC5aairUv+plS2f
25g2xnsXMLABRDGut3grNw95davM4nlGia0I03RBB/biJfHUr78nE1PRqCunZF6J
LLnPbn9wKNDQEPxQDKSC9XJKVWtNdlIN0XZgyRabpUNWhfwNXB/5WGYjGdwnF+Uz
ODUfFcARkRJ5qVvR7JVKEVg8+AD5Qzq62Cn4yki0m18k2NAwn54p70iDESLQxL0E
WTZRjWCpFSgzah5EaXVsKJ5Ng0LOPIZfzgcz9ohdjjRo+cJLu/fmwmavJkQUsqtZ
YpZsFs08F+mLYqSXXPkfsyZg/D2LS/7qKHuP4S4RhVwAbz8k5dsAPBdV7RCUPVKo
6YtmqFdC0Xa/dYgbz2HSXWFGa8dbPAKiWSaexxAj68C+gS/E5PhKAhC43wqw92LO
mdvfqnw0ePFvMX65y1NM2+ieBIyDLPQIXOnAZMBfkKqDSUndUAp5bkpVMDhMe1Mn
du4im+S1wIobtE4DVmhd20jnyp7HWIeC3XtD73loQmfN3bWf8G5QRxwBaSJMQDDj
cSLg50Xz7c83Rin8T7FvR0DLoMx5bRqiwWyz/TIp1YzNi44E+b4Y2Y/vXaL1rcbN
DL2OJvzo2tiI6HXI97H8VoZpljs3MsNtpLQV4ueqHaEpneH7GdkpiioUVHuFtqwM
BMhWYJzQPhe5Fj/QCvD90kyKHGDBbHHS4gKJDG/hLZ013gjYy2eNU85F58lPLhp+
eTdeVV552sxb0qC4kkeiCQ9eGWMis23awkU+2I/gnqR3qBuvAFkw6Mgn1ixyTkkO
MoPsT8Xv+VmLC8npJH5p1kSaFYsIysu0nOZu+vPrxqfX4MgJInZ0w91s3/sb5kOa
Um7+UlkVF/Z4nH0yS001fKN72okOTYjEgawRJHM7dIRlXYs8WQQeNwBvmAAQroXJ
krbe7KGYpqn+MphRrp+yupmA0lR14eaOfGYddIPirgDfH+7tm1LyyNv2wttCCztN
D+WaY6MOLFy/Q0Sw7f/LzKpgy2HQ+M+L9/C4JorjiB6J35XQW6IWKkhGl39JgJGl
ZOOGf750DEjYO+tq986X/gsMEBdgtempUxYrUlBDv0L3jRSJBN6omfz20qjOdK+p
rih6fACj2RX+C76QU4q6rJkWfZjAs5x1WL4Krwymz1UzuciiWlKllaErWy7jwAWo
+5aDyG5ff6FSwAXTju/B7bwkk1Wde4mp64FjmMJk1OtKYyxPp2IQeNRrOQftyMlv
UMtFln5oHi21J+jaGaCE9MuDyBUmk7GzyPBTUd98UjNIx4xWsmgZigoqNLrin06X
Sd5ubL0s4ZDwS1xizv2wheVfQl0Fq9N6076S22vQksvT6Nj/M5rIWaG5u1YdkwL8
rTJ7S3/CEO8PaZhs3gQZZATYP5fo22/FvFsPwLRYBpbCHFwQVr8pUKkXUDGjzHIZ
hDy0nOviOPaAhNtspkHumTqfl+ENGIPF7B0vt3VPXZlD2ZKIXRGcnD4zaPyob0M2
er2WATwoiBQeelGB6Dw2IdBE2WmBfhCWn+qQqCSGB0phqbqK5pgsAxwMOVY5HeNy
tOyfG/YzR4Pmeknfu2HM08GmFI984ciJgnAmr0XaLRuKiLPId06FVX356JPuHl9Z
1h6rNTKu3r2Hw/ztspbLxMGJia1pfcylOmrPoyNxARC4Sxf/5hTW6Ppxd5xtv8O4
vZVuQsherSw0pKkRXqi90yElDs7bd1bAXmMpeTadth+N0gEQzlKdFE4WNMtwVMVi
tsna4JR0Z80rzrvrOwQ9IT7gVByHWdJPAihKckhJYWcCORotWpc8YZ/0sZPuC6hO
reCFK+KeCx/NI9lIQCQ69obP7KV7Wwrb4B14Rz/w0ETyCpE8u1UkWs4hDCu3ca6W
rcZvw1fB/WJzbAZ2huvHfSXucNvhN3VeKDsUTRBWP3ZMgtQAv94yYGYrfuKTgS+S
q70vC3O1G8pHEzy8PScFONv+rwEY0unO9I3fx/AI+jIK0oZrSp4kpbz5tdJbzqGo
PdNLFDRqCsHisP3Zkh6Uzbmw6YCHfa/gk3oBjm8VoMV3+D7Y4zqmD0BrOujDTSu2
eZydvhNOUho1d8/aYOsOMcc/G5CjU5PmA0jc2FsrBrMuQr1rfEzM4fMjny4CetY3
FctiAyKO/ncBju4QLegzoyEs2CdJfuDG+x1viViJl1G/HRQ8kotXvIvq4gvhMM59
vW6+vXck0qH5I/pDnTGipI0NcU4xIoJXgK+LR4QG0vvuwxyEmReVUIEfqqSnlsvn
5tzPea3ff0o4DfCZmiC41X/HW/5+q036dxzxzXc34cNcXa4a/niywSXFFyKoQ54B
h969VhkVk5MSRHpklvUC+Wq2n6Lb+aADg4/OsbL1okpaD2etOnLEmvROL+og062/
xucF2wxeeKsZ9UYRJKMGsY/N+xmdmqAoMmVs3ySYBD9fWGg96NLH5m8Et9vh7AKY
RNgI2Rld6jXK453NUGx6j9MlxUOvuv7UhZXFwMTj1eD///SrCB8I1WRmqoIjHsvh
5GjOiUt2OoNDi37M4aU1qMu4qTXERB8I4eHxwrVHXKSuXPDD+tsVnMUCjf3I0z/c
8f43WuJ2arfc5KH2qv4jcYoFk/hYdOjsnyPcDE3A/ZIQSM9z9q/H10BACIxk6Oc6
3cGLKg1Z8DB3PyWKIw4GAONlg9VYfdyHGujZaYDrKgHmaR0WweKcq0mAe/Ckm4EV
/hDRjEd5uV9+lxRtwSkRYgXiB1uuVzQ9GYp23uptedQz81U85N3Mo0RCXwuoAzmJ
IWxtsXOvyM0WJpdiQap36zub+H2Hm0YMF0PGLan6zY36cjETiUlLHfcHi1tJvhlH
YfYb5V7MpU9n75Q8rw7PdQ38V86nrA+V4JpqGyC5cUEWtWajK8s8kwzeYz2gJ8D7
JFnTSsJgPguoIug+VgWCQ9/p5zZ5xMQZ/mioAEHM3SUwEFz+Oq8mkMBupRdzazsi
5JXSMJDeoDx1PZDuMcFjF2TP/GS8l4ifVY1wVVP/jswxmcWliVaubdj7R8o4wmIA
/j41mdbIzF9T6ghAQH6wMtynfqwVLc8JiDyLOos+VrmfC+X9p20ksIEGpuwA8ETU
v09IgzmakU7OafJQ4IuXAwGTUymd2cyPxL3cIPVGeXX03Ufg2N9aed0IQOLDomQw
sytghbk+54JEpnEvTocbs1b1Juv8zXeknc9TiXIuUqkeBj0YOmcv1k9p1Zjyk6PH
1PIun7GdIoGtxnMsxFTi8apyOYhPqODG712zTNIo/TwVfptTsePdWr/Z9nQZ3gQ/
trf14MIIWE/r1IyktPDsgwgIendEUBYMjh3lKO/m/rZzHswlhFEGUuZIS5XsDuzx
JPBw+bnLknv8XNxdsbTqkSVTUGYu2xAzwH4WbdZbbgKHzzSpYy904SmpMoPE1ew6
u8WKredW3hB9jFpfPOICQGKzsofGsr9EkV75cZAAlTHq9RI1E5x6ORJ6d+RaaX9B
fV/qTKVCu6mCxXXe99dyNzb04aQ3VTG5Nzbik+NATUh7pf7uzzMseSZyuhFq2QB/
yI8W1u3CPP19onOFvHC8IdjUEYnhKyxoJ83M4TnulTDf5chHlaHUw8H4kmTkh42k
NjtK8rOqD0LDOTIRgNewtmY9IRftmNjr68c2A6KLOlmHtrsMbJjyn4SYxMpMgayo
eWJpTMwV5IVvrWQN+jmugqRXNekmkIquZ5Xd1NWno+gT0ltz+mRK0o6uy1WzlMbk
2CdGZxaTAdNCPqxLjBLcTl52fZ8DKbMSJtPFUv36NLrNF7eJfW4wou/rLJULr3/M
UbZ6x+vD9RLT7jzrgd02tOtQFn4yL8otyOuPA0iPN7QQNGOIt1l8mB7H1grKvAfO
GpQUUMlEe8/NEjqZBNtkD9atfLoAakffhLv0USBURFdBGxGUL5aR8WUCNfppM2lH
ZaeOz2zRwCu/gZKyA0/h+nNx5glAETleQbc3H7uBvsW3HZuOuefScQ+yDpUthC4u
DevyXfo+hGNl+yNEsBSiKX0/y7ZW6atg6vrTAKubkhMsdpMsz/KYFSWiINfQ+lUK
zWZJHEf+WLx6GiV0xtHU52g14R167K09ZyZz5N+oTDcwOrj0Ea8gRZF3DhmwKf/a
E+y3r3sV1E8B4/DKjXQLE13bVSzsPkKXW4Yi+VyesN1AXOLBhdPpNOY/aQItpv7H
K8zk/ic1woEssqmLAamRWTOxMF6+ahY851/nAcIS3OLy1Z6O7Mjv6RqA5ZA+90Pg
5/sVfe+SLBcrbhqOv9k2u7plDI7p/STLzapnz1O+ehcHOE331Ud2KMQYxgOeDYzx
WSxuUy07Lsawasksti2sU44GmQPzRe5uYVaQhxL5DmayYm3pgBJdRNj94y5+3CpH
tf09NaYydiGoQwK25fwrrc40xSCee9npAQeDdi9lYVvMv6Zp4avVuQMutXrprm16
1sJRpilJCwwjL6KzjBnBtavRyEyhs71dQ6iH1IdWNsFKddZ6Z8AMO+LE9Y8ZcFTB
OCXV5erqtUweuHntYOJ6A3Y/XNfsjCezD5A+igLymh7p/meTmok8oDB6OAeQ4TOF
R6KZFfF3FQKzsskNLLyzMe9t1qdmTBHU7UsbEJVLV1kNiGiLNL9UGEllyIqjAo6F
2Wn++hC+FUFMDprOhb+j4OXYHJhk8JsrAJprMyRZ7pTPRa0ThF2hMYmDhcKtKQlV
luxDZ6Y2DxYt9OkRWQ9hEhKHKFt1s3V4S+xHKE37IK1QKn9cA3mBimfAIpZq54J7
slNiGK3BxmQFidW/93xQZHyEJbaVow2Mv59zqwvQKoLYwYwbkgc/ALjPNrvCk45I
hEnVjyZB4T/ixXug415shA+l4EQniroWz5wPoTO1KiHPhLlRk+nHq8LMetJFUgji
TXQK8+akYi8FFxGlhNSsl5uMgJTY5vHmD8XGMufndGH3x4EfJLn4H9Ixo4NMz7/A
IAi5taNZHR/Twm3jkXFVUUoRQ/WIHOgVEzmFqqsFo5vCqO+0GLnVR9DQjuhJJF27
p0iB05czsUDIqGWBv2GVR1RjX0CJJFsuiZ+sf5IuRKpgdlrhfrZ/BOzOlwpIuGYd
jCsnHzYVKlTREr5yWF4wSVfT4Zq6nH822P6sHwfYqMPf7YWeCQ9ANQa9E9cHfXLD
57ggSket8988hTK7bWr1Ukf8GSWko4XF8ElJ+nMWLEIoFg69lz9end0dhPhhrnwj
mOw6eVVVepVwjjCNpGPanuz/M4Wr5qpQj3ZzQWdR6/TW7gyOisuILsp2wZgnRwbt
BjG6xDAHKHeA4iYx4aGLglw10BafAlb8BKTEmD0UIU0qC3nVmEVM/Z0Tj0k00jx5
MHMue+3O26j8GdBuE/TAcnTUI7VfKL7EC4mnKkFpGzbZpUwW2/VXK5Ax14FQg43k
9i9EqkiSnvgBqcrgvs6xQuBCIcxPs7mhMEPSZ8ANWiR18hyWKeAmlBYsRZA/oqGh
XUipISDLMmtKdTfHme/eBlZlMB/QbWsF14y7h3s8FTPZ/5PorcTit6nHAQzy2heb
/cIHETTeKpUFhmqInynEygfjgVzEFlN8/acm4dBA1orSm8vkaxnsECrLEhl/QJ/d
+DY9JS9ny1k6sqS89SnGCywsmhvmolP28Ip9HR1DVS59E9CGvuVpyn3w1Q7Y1AGX
Hb/mJQgMu+gRD/Y/WBuk0FX+diPwhZlExP+4BhVoqvEcg2aXqmPFwPYngbAiR1aw
v+icknlxUWxvWVrhZaGklQaz5XW6IJMkuKgwzXlYAKlklYOpXSVLItbyRX9H1h1b
gK1wSlC0D9a0P1P4pJwDDqw72pZjHUMG1K7s/UBXaSdNfTwwbBnYRkVUpFiZ3ZnO
nd01ZASchRxf4ORcz15+uOsj6MSBSvBdqQxCpZD4609BiVB6KmNMMEg1TBoGW1lq
o6/AbLyeiTWRSx8OlDIDUC+LpWjwwHu0Qd4TKmG89+VV452OO3yIsV33RhK7X+wB
wMAm1t3XmxKCeqbtxd5KXheGYBufwkeUWlJEzNRPtdWUTELAdFbN2b4LgOnenSJ+
WSiCbCwgQ/W7tX+/NN4i8bXeos3kcQQea++8GqbO3Z/gYVouKDOUYVor204kmb+t
wuId5WjJ2mRlcn4qD4iTvsKZAkVLzuEnpmLH34w1ojBRmEbk8P1LMYmdJNiQhDXO
0VHP7J10nEHYTgXn4EvKvD0l0wnLFDWDm48Llqb4Qo2lXb5yQCfaTn/gMSS5LuGH
91Kka4Z1pwCen1wq+bmB7HrtXRqgJMPM7Kn4IR+RU0k/YlLocZ1tJxUmBp80D4Al
FkbuvHQgLHf3O3RrIK5bE/TxL+pVOjVWGRJBlLx95AyL43I2ty4frALQiWfZxXkl
W2h7ySzfbTi+nFZoMbH/WcsRsmQv4qcrh7ZeT/GIMomC9J2qwaiRKBMscqk8P6bq
7bhyb/hRWLAuBOuO5eIlOmMQshUKtz4FESqwpR7Meo1ZYZEUHTXou+MBj4vcpG3w
DAOyEzXwgmvrPS9OO3u4tP/k9VC/j7cuLzjLOMsq7h3dlvQs69sLX57v71obo8fD
xdR1L9IYpjy9FLx3cimql6LODhR5+RLsg3VBRfLlxLh/JNgZfTZ+rrzLLL+/1BdG
+5r/Z+c7f/CmuZQhpBfgkUH64NTp8wKH7Mlx2qmMWDuYGB0nmszLnTuicEwMyVLI
Wa300SRf0tyuTioqwxPp4PnlvLyiTLuMWtH4Qg9AYwIqWmsNl/UGg4hoAjXfXEH7
o6yxZ630nm3ORQomPQiT9Un0Clv+2Hf5PYLQIACWN5mxtQiieEkt9rykM3+L3LDY
MD2k3Lb+saHhPEga1ER6VuLoTrIbPSAHlNKwGGjdshY+Wu5R3aCSuX9DzQLL11Fx
SRl3p5dBG1UOSMME2fPQp08rFMAOiatGjEKv5eDnhT60YvdbdyOba9hApFV8HLG2
R/7GsnT/nVDVmnSEDVRFvar/G/gxpQV08shhLGiFoNK70CQzLhEzR6R+9E7KvoXN
DdQztPiABRbuS8Y8+Q7V612cXzsyxbgNItimSfDuFgyi/u56sH2GQLsv5HT1Choe
KLrwesh6cZ59/BrddoAkdumgBHtHRknvEUpZNgGIgNJpCE4BhWBheQhZUSDXrM5j
B9PpZb4689WTlZkaD25njtaoVeS21EllkqhW/b6m960IFvB3sgSn3Ons5eZ1QK8V
uNWgfy5HxmK7EZ/VWLPD8ugplAZAhGtqEq6BGJi3OTPfeN2S9eAiJDemrKtQYrmw
QAVdMX0CS1vHWwrEsnweTFlLpSkDrF2tQdBjHA6Zi4sJE+ifdZSfwjUap8JPpWbm
kWTSVt5h+fIEY/bIOuv3k1CnjM+n21XlAXaWu9atFNhorQ2iQGzWg68ERhc8CZbD
LiFp7LSMnad/WX7vaR6wERrBLd+4MoAoFBjue21tYJ3sPepTU1uctU23hSyYRY7h
1rlwtsFTtKeDfxz2JRd21Zi/E5Ba0pR1NWa0mDlGyeOH6H67ulUEflCR/poiABBi
TyqGny085UofxoIc9QEj/bCB60gd5+xR1GpkO2ySPbJifDMk/VDxubbCpGt53AJu
qLVbFdysTWSe0qFFGkD7N1v9sDMQGqnlyjwj229GLLQDZkoIplI82EVlT4w7crsW
OvCyqWbBSTMkJ9AuEkIEs/fBLgLqixEUSZQNMz8AGzDQdmSG9JOomKFerhr7P/l2
ZOWCRCLN06Ay8toQFwHqbK7m0H8U8F7EOkDtpYOMIyzE2iAt8TRrd/cK23OWIzCt
b6tpr2INbzwj/0qxbCukIrfWPU5VaMM0U2DHfjHrmiNO6g0fl4XjMyO5o3PreC7t
uWAlUnXX3iEyU3ZwWJ23W6f26CKEkTjTROd9iyeqWKSyioBew5Mazpu24Utb94RX
oPrsUwB/+517KFI5Bqjs6TRk43s4AFjjN/HPnCoMtjZb63rKLrY4RQt8n+jE3ml2
k4Ygd88M2wDzzmMZuGmMHpJ3mYPW0+I+dKW5lg98stqa+4AqIi8QAwGk8DZgUXnM
yDaQKugewhPJMou9tSd0dLH1PU61tHXHDMI6gYfppd2tGq9f6ITimGtIKyGaSJ86
5KCh4SOAxU0xhJPvuaUW0HZXtMRQAj5H2fuzwNyiPuJkLji6Fd8ovi6qTPXr992E
3rxicGQELnJ0U5QWI/wcbIsN6FBtXBrJh+hsBmEW/ilM5F7RjtR/o/npKm/CbDSC
YQbp6GMiWDLv6d5SNxbugBBuXokruxc/BqRNCGf25HAPyRcBCGumRCmrLB2qSbV5
+JudEVRxpLm1U+1ze/kv4ATCbVMEa/rxtxMlMygE2baV3meNgdOZ2EKTVuq6PvHl
GAKBHlzPwMZY+AYHYISqx3pMMXB9vyaM1LT9PDHQqnqgJg1LS5EBL3OYKML2LSfB
fsdWKcRqWR3L8waif3qxkfSPOK/EbiU5/BmcUWbnS+Y3+n8tfbWyi6zYJgDz6G7P
+57YJpZsVFVdmK8JFeaetj2K0QJJvS4FLrDRgBDGdJ7mp2181+2PntcMQWoIFgM+
ZbzgW6fHt3UZYC+pO2SFXk4GFuWeSHRFK3sv4wMZWyZbsvfKguRG4Z3kUQQFLHqh
Pk3RNI2Ar8cX5KvF7Qq5bckQmg0p47g8KgjNK5N7nutmfg+jjEth3jzFuEIsFfTQ
Z2fi1HfgDSTdV5mxe7pXYtA39qL7tKB9l9xYAm0GYYmTc3aNblXB3PwUWxwxmvAn
R6oO1VkqEQus+GzNqbJZaGFgBNHCpK0Cn6dVlH1iO0hJnuavM/dFKfJy3aH+TT9s
aGgbEti5nQj9kfAm9CVq7c7bR2CPriebenLkg5S/Prr43CV5QxArnIlYgxl3sLCI
2fgYEJZ8vzK63lmUHytElqaXTkGux0AhgdExmsmbyjGzvmIQxTomo57yhVj7aZjo
Dnd2T+dYCImH41QiuXzPDP3PetqXHIQsYYqfWHRVzqn5es0aj0q3wn0Ch4HU/jMv
oZnBhAs9nuwOy/ruNxWU+T8tAiPsEC37Gs3PPFLVjfI/QYlNQqM4wJH2Vdw+K7bD
0ywgHSKz+3GLR6zMrv5BxdDsIwBqlMABBTvfqwGd2op9sjpENNnPbK3wksBSWtWp
EbCGE5t7JjMSh3MBBqWO4kjDu5xQR3J7qFm+jBfP0wwMcVt5prtxT9CCHmefRHpn
FRstpx5/7vIDjmCIRkanQFfTnA2sr5uxxjb2gVapH2+VqYz5MdS0VHxPnxRxPYIK
D4RRzZVrzhwyN8b+rSMVyNz3US2qR9JOLzmSHz6kRyXvwnvlkOLtsYhNCD0j6YHt
cMA/wcIbPvvBTfS8qvZRU/ImEUbBT2WA0xoUPPtVxVejSSB/0m9b0esSM1f7tJd0
sUKd9d6MoIxNkCX85fv2oqf0yUc5KUB4gsHhUfkkCOEOKnRUG9BPdk9dC6ZxXRny
iEUwYrGNLfOYcGzjLGg3fvffR2MuXiN03n5yI886424Z3gwMiso6nycXHocGolV2
rWme5S9I8PyWVM91YhLaUq7WbMMviqZNyq3qjCsHrrgirsEH65QEiSERghmYvkiI
MesDz8hZRtmCcxAJaynDVh/hsYeoxqDVuFdRSaxmcYrRctyOk783RYmFluqg8Hp1
v+2t+aD5Oz3IO+3EEd9QfgHqjkYDNucUcKk2K05ntrE0Yin1AI5lm66hxuoLTgU9
UIbC93SljkYahY6XC24JUB7LNCnGdyPFub8m0R11Uv/7md9GmFTBI6JgVFz5i8qq
lmKBHFDuY3VNJjSzxStxb3M7j1n7ZZbjHEiqnRZtkM1iFMUC4o23iu0j0KabDlpe
inkchDD8ES3wi4e/f3PkKR+O+UsdAkf3ht18Jnp8YkvZndff8PrfmVvjFE6xbsW6
EgMW/zotd7Wmqf84w6XosRKtt3MftYP9IDR1IXdnlzkwCTMLQtqwHXadSHh922WP
7Qwdtl7tTFjzl8LSTSzEjA017P4wL5fHT0myMPvcJeTTuWFXfkhjna+M5MWHN1vn
UjIKmnld1foY+44lhF1B97+k25l2wCfnF5m0h0+7938VaB1Wid9bwOlhDjZO45S8
Bl0PLIyIpOUsZ8FLPyA5aPkl8SyM9f7Y+jx+szEOa6N9fKUqoqTeryo1aEvh8eMT
y9JpPlHgYtqrbB0SZ6UjYJJN4zP1y3p1LKig8MCtXtGKY1kmAzQRnaViaxhCvLdQ
kO2slHR9xTHY0jOCYPc2xHpaeNbr77YGfD0NUt0GOjqZQ94GV/Oakmh6lI6c2e4+
oDG6bhKHGBe4NjjQI/vK/s/uL3etO8P0Hg6kR6VxHUd6JXrErsaQUJoa+TjWofxh
CAgKFU1DZNGeIzUMBJfpN9wihPwrdwFNmEMInQUgn5/544ROqqvFZ05qs4K64R1f
x3bbieOUQN5rShLCrYSZEZakmtZZxCKSPBQUVbca1Ie+/Oos7XUKGG4D0lCEBAJ6
7SI1FTwvYDp3M3dL1hY02ZJjf4aX0FfMe1IKsD5HODHP+15HJvvJAjlqoTcUtsLj
F69MUAuXxdxY1xagS4KKw3RmAz1b8w58x6xdm52n3prWo0MhA4DrbNRyRXKAWw96
4xmvME+SFSNj6ACG5EjJ7teadC7JA+d14YYCChmjZ8WJx/wwHe/iH2uZhkI59vvJ
l8DwSd9yBLOYybYbXMrbogUCCNdgQYKQh9HFUxJ+E72hTHV763myETgVM0Lkwpg2
mmTUyt16FoRk++yWIFgZcFK6QucG8ffBVfmGVxRuZ6LPXfakBpZo7e+6ub6AUaNd
A0MSyIgHikXjGLjbSCxxo7rrQ2JrzntgrpmWgLj75DGTqgYVmGd/ERnVovgq+N/I
EZ84TLka1/RbvdTu213wdZCehUnQOdfPlqzXtXbJYvFVzXQ4AgXQ90bicuY3G50x
Uzq0NqsoA1eEyw4pGXKaq7Woy3wZT93g44rMQDHKgri+hoAXDExnS3KaahPOMGuU
9ZcPyUz4SPe+Mp+7SV3wyWCqPuPVAFHPGr579pYM+1TVkAckNoY/zoqr86rZqTEU
Otp9n15cO6scoNeMEEAaoX1Lo51gBZCegWNgprfqegK1PmVMAT1YXsZxGrjL0FGx
YzqMusfsnknylVlTI8z/1ygeNbMHSikx7Sq64KepCQH/SypxTRNcpjP5uOgS4HzL
7K2c+HxbGZ/2wP0/ROiU2ijJ6pcHPoqMAQbaYNfJP2bsXX2hxMDB4DSD5ViScnmA
rhB+HaaN7Q0gTmF6zmAAt00mgfRagwRyqFghv5iikyJLVp016ai+DWTBScoGOPbl
hbYqcS4crRGpjAWdIy4c6O4SziWtVVgLck6E5Kuc5b5x9kTLAGpiQ79Z5EFIm3zf
34nuDlZPn2bPFT3qumN8SK+KO0b76Tabx9Pq2dwKsh2zN/SXG0nUMZuNWdgs2paJ
OpOSKsXoyamUQdFu/TMLw/IYy+4gsYgXJ6FIlPgepxuhzJGnzfRVwWqAwAX0t8fF
5qdSEBs/fKMeF8Qb6RzSfUedgMij4pIaO8JDFb4pNebTwd3UKOwbndCEMnbkBYZv
Jv2HKTQnfUdMrc0XhqMIBVGQ5+W8rWZGsKYy59L9IZ+nc1wN9RrWLyX9VL5SD9Ib
m2pGemNMS8czOvdK7eKyWMS8osJUNgsiBrkOEXxLcLfqPtM7Tlij0DzPAXpAfdxh
g4eftU1+pkPPi6Xgq2jlMdqz9BnkDyTXmRTPOavSUCEwb0FJeWCdQq4MQCKzoSMK
AwHPJutY0cC46wH8jOhEz+RRDV7Ggt7MwHc3LqNNeRTsd8qSqPq5ROePnD4io5AZ
iTloTtczHB+Eg2CW9QrHiNPti7eB8dllov+4YiLte0r+BKfjT023vWHAFkBkgMJ3
HBBa2Acdy0j1GPiMNsEURVKDNnsFQG9kJU0Xmyn0DPHK98abDPfeK2btiQF4cK3u
YSjRiIj8S4HlMD+rVYimu6st0XP0hAK1ZvNI7SCGhyJoEO7uLTOIk6GjwDN7HQ2J
GzE10MnQXdLfdZ4368JwFSKLpbQkDc0IqXwLlwC8aI9SKpml05S+A/6SEQifrbEk
bOZrXAzlIuUzVmal7Y5yCT3clCFUsHNoaSAx0Wr6WVnvF5Zno4N/2iSQCR9EACeA
EXgG0hkix8siyOqxarOapJKkmc8/M1setAMwGzDt+k2kVQuC0055yvlVqwlAtJ2x
dooE/iTPrFr0Be7VKvG6XS4BACUms5FKQQ7vlrJzLeWWmKZG/+i5K9BEAqvMu8ZH
g7EYFO9ntrC1Jekdqkz60n+6zaeX4ajSmgvHCcal1SNslDp2irXkfT6cA4pKBvZT
w5lRfH1NcyZ1jLBXiO/iLKceWghw84YY00/ZCMz5bEEWR4UMNFfl3U18BPbcks7j
3aGwZ/bedYIMCDKvVitchc5YSbIUam4Mde7YdTdxjysCi9GCjLBB+iv64WMYDwh8
W+xuJhK/ZoUsiV56hh8VtHEhaCewrZGJL7F/oGGhz60sUpIPTwgrtfBSR+qRDh+2
vtYb0CZTiM7alVQaKX+RjLhKnXDQQz+AKrmvCDHMZZFVXyXHwTuu7hXoRpuN+L+t
Lzg4vWKymEVsxDEFuHi3+LeQtlUUnsTeldWZBYO7l4nreMuMIWaneNqXxhF/VFf/
NLaR4RCNAUrm/d3oGH1BbMPUF7YHo0RiebWSuilgJJvfzNpnqVgn3QuVMnMNXe4O
XsJ0RMpQF4nVI1QSWXUAKCBVfUukCivRW9nX51bys+/3JxgTmgEs+cIQy9tkiA98
qXPi5JnliGBcMOBJ22lyZQOBMRIiXbbgO4pN634feLjcJKxyVKcWYkhNtWUSXti1
k9mBc77Y24NSeEj3197Ra0JcI3G0hiphENM/+A5YnponsWBlZHd9USPluMZzlsjL
h3BEv35T/LS3X6T+pRThvmGQ3Fz4HsMxy7q+imIXteBrzczVXfu5HWjYhZ7LMCbx
aOdycnErPU+LxdoDnsTJ5xb4j6Tc59AMP0O+BTzNvWtsVB8fb/1ebTiDhf1gyFrl
D15HlhKOBLqBpyLdMydgXJ5smdvbmCcs/CUsas80MH926K2OROAbN+hjBHlF2OL5
WdHAjy9uP5I23tV8OCVDAM/f/D7JuQ3IgRDE2vcfEW4NG57ab7aTPtaPCHE5wt2/
Vap4RA5Jba+vnAtS6EODjO7jQSgcZ/6Yg8HxvoJGbVYN1+rkGxbg09SnCx46qEos
6nK2Q3/0e2cho3qgpLbx7Cek4fe7TLz8zL41Iw0wwQtGmjDwNEqpYn2pTeJ+jzjt
KbRINIKWCMmKn9PB+1gCNvcRuk9fZj0XlIbY6TvnY8v8itds9tS3O9t4udinH6za
d8IlXGy4fd44EIl6/llSIMKXBjkKBTajCtRuT7p+x7nWckJcZC+jSWiq9pPCRqUu
qF2SWu36io6wfQc/MD2CUQLk+oiyv5GIRUNtilh25Henfs2tFEFGFNn8SBGtZvyF
dfB8Ju/b7G9qT0e6/+4uyStrQCXMJyf5Qls5irfnA7bKhlUT8CDscgPwh5TgKkje
hKVR80eDFbGNI2AFtsUS2BGU3AiqFi303Bs8PHimxqcBDKeZ+0F2rjuyRdQs4+P7
HVoCP/bHRGVe77Pb8NFT7ceIsVo2I0SuPdVT94S1Qz/vJPq4UuFBbeqE13G14+ym
FkCpwt9hX5N4WYhkRWPArXaJsJuUyPSU9aclEcfWsKmjx54tFdE2gkAKJWVM5xQd
+Q0vpQFdSHXiIRy84i5D8b83TfA7tVNsi2z8O/mzhptcITXN13Wlp+K1qY0MbmBX
qKIDl3nxb7f7k0jqAu8u4rAHk633UKzBKyRWAA88LuVFDsllkwIKKKhraslYa4Ef
g/zsGm+zQKE1GRfwuYn0bUlYGy92XwLOpx7q107Ce4FVqToYDJF2k4eQYvd0bGAD
jsOszgGKOV2GEiOtYl1X3TA5w8Ouc7bz+SOKRrwAd/mAS+7XYHXpna+S3+hDcC3L
i3mamtUSipyCMrYwa1pi46XF1y6yjeya+3PQWyjlLE4MEWgoC+FhZbu4Esma8UDx
FA+AMYemWaj6e7oAgBtHZbjuUYBxwZ4l+uYjqkiGNePNjRzVDq6d0zEpV3nYGe7l
ReNKgvg20pFJGGQCFkjIm2lpm89xLIp+3KH2R50IidvLt78/cfvA4L8DktoCIyUp
zcIz385OeFvpmyi5OATCrfc9vM0qdg8bKYPC6wm4FJUPRVDVr3y4P35oV/uM1KXh
pH8iDcRLHAr5S534E6AUc3Wz0LOZW7zIAs+DwAVrIHqcpnWoBWO9SXm0AN3S3YaJ
x5L62OgoxCfhyJRaaJ207lvnJO9cV2i8y6c3bAjhBH0p3vbQaFWfiWz8GmAdRdO7
BY7Qt64NfzsOTthBlfyyvzHniA1HGXLFZ+g5iDc7Zkaxo/rMva8mcwSn+5QwxgNr
xzp6bWzqgp9j5kkHQr6QAbLIDW3dbEO69Af3YXf9e0PpmSB4duepvCH4zgM6JtVn
cPky1DPnCb5lvIIS6zTyoxO8xuuW48KB5nvzXiyEROd0QEzELBFVlIdwNPM87Ynh
YA7s1uDgshC+etYIOxs0QL1jHtlkirpG6wG9RlPgJTK3jNOsCRf+VPzOd8i5K4s/
r+QogJbypVn32eBNzqV7OsnT7dSS5LnC0gmDuKB9xq3mq84q7JnHDvKajABvyjn8
0V3HUYqjBa/bu9vAaxyKKQZAxdPh0ogBOBZy5kTrecBqSZbaX5Pm456tT+N5P5XS
DhpqM7jLlQIx32i3Vy7Q/d8axevrm+d41rOJGA5q7kJh6acba9aP4ZaXX6kkJsz7
mnSxIFb7xEh9OC3qxFyrqQ4EAmysg6Lt8fRe/8yuUaIB06VVal+3ZFjgbq7p2PxB
lTqIVtAxBSHE+Sdd5l/KfFXhQvPx94svxEj49n5btECX2xEazYYMyJ0s8I2IZ8+7
JKE98driaXtANcGfP0XS3JGG+JlQZoNrPWjIkXK30764r+CIfWZIC4jzqPUG1UTj
JVqhySCIscFkpVi73YgK9xnJi38k1KkoCGsrW/dPKoe3UPGZEgHliwjPDx8HykOT
91Y5L0b/biNpMQJ+aKkA7qBFZITba+zjGIXKP7qp/b8WKnWGLMKbpsYAO9jc5/mT
f1OIBSgT8WBpYCSK/abrACUZFeAbZtzF7VgF2ax+PagJwg+mByZY1kKNUYEVnDE7
zPZBEEalhhnGe9k7bORuDrFtGyM63ypoATXSNr+4MI0OZqmfUDfy/s3oDAIu/qgm
11fv3Uw0CsKE5g5WofkewzTJaK43IUcre9ZLMQIeK/HO+dWcfFZMVgu/0B/Y/jUW
qJYj1namgkGECWR3/UOlpzIPmm85itXKVuAuk203t4QvDX0LsG+lVnK/9VRBpBk0
YRdCZQZm64wcrkP8aVuwZQlq6j78Cg7jLME8QnLD7JXbmRxtCj2gBWZFXhX2d3Rz
CnIZcUf1cyorV1/bhko4ny9+4YSnyZdWF8ewhhrNNy1HqRoelAyATMPBIH6v0vv7
Nu6MILieKW30hIIMTUsxb8RajyL+mg7TPWfpsl4tBxOeNAQK7smXjLT6MTnrJBtH
Tm03Ek3C88YSyom//0yAFrrmKb/Ud0/Sb40pIEl437GgyF/JDQS9ef5luWZ+bNeY
Jp88An32HR62oimH6PvtwTUqFr/uYCYWmEKo48pe+znjYaZXvILJfBmdmgHMkGx+
qX1YAuucPkpcBORqGvZ1cw0JxFmTKFdkbIHSkquxEs71UVd9m46RI3pYbOGgl0BX
XbO6zmDw8rBJcdgfhlQmaFQriOvT7lXzU8y30cDb+ZC29P8NCWrfFmmJf5TIxMDr
mqrsMiUI4JaWOTXYOIRA1STjPbm7pcNzQiC4bADTn3tQgseXfH/RTggkMiYHsV4b
CSz8oJC7mdoo54RTOyIPN17bOkOthBPb6ttHJXUc73pndEgAt3SR8xdA9qXukKiD
NK951ZjGvAbO6BrUvCuq2+7lB1SiguhLfz+t5TyhtlgW/JEdu9y/hY4u5/CREuPu
lMoKXJEGmGxj0ZAAcjLscOc5xd3w5gQvw+Xs/whkwpDPGoTyVTMxHj+niodKVQNh
oI3Te/LXE5WNCyKsqaAuGYQsf6QlmI6HUEQaGssxfkBzGHySwHd4FGhIUffbwJex
I9Gx0/OHBY/56ndLx8IW/j5TQCj3w3yZkzl03fHHrRBqPnohxKAYjl+aVYpbTiS/
kTgoGUNKDwm3BHEnuUivNfGg8PC/aY8X2Zyv67YVZh5FFYUwfSN86QBDvPkSaCsI
GViNJeRMWricOuGbfOaO9YI38P9qqEjUJfI8wRU7V+6atWpUlnQ4bNm0bGkkO9hb
8ajmRORihTuE0bufO7WS2SCAhxm3rJrFVD3TrijHCNn+jGfTORZb4agGyTp6hnDS
7n9kCuPKpA1ntwqvmK0qhrjRNhXq5OMKOx/LEiJAK965HoKvVDDciJH0aMmlhz7B
vU6p+G6uHyiDFCPRHte0uwKStjMeC5PJ2nGAkO7jit14hCLjHYfN5zB/2htP1Ccy
8OKWfhATIPIPcynTtug/AHqfE90X7sXjm5hf4euChptc0xu2Fh5iv0WAFjgs0P4n
6IRMq/JOQ7Omf1GMzKeIlyWNq4ZrFEArnopZqWas/3FzunwFXBR02R1jqDGB34MK
bUzjJUgGH7ReKZqqLHcdglXbjBeSnD3QhIBnv5nXzcGwvwMEynTDoXo/JN2DM6VW
oNg1Mj/y6nX+9OAd69LUETroe/S9FJ1Nd3qM2vM7I7UxHHjYjlptBm0onXnUd8JV
oIAvQPV9Yg90xbq9+Oy3GN1ylwaI3jHnnfqTjFUEBkp9paNsFLSRwr+G+OqlNBLe
H80eJJH5xxUfjVU/vptehqpRDhAHrSO0sJRlsxaKwDymRghbrP7S8Eag/93zlAbW
dl9WqiaU89QW19+TJxbBLwtccE9Ebm1pWx+pK2H8jKTW/shS8pZfeazruSKSGBkR
GaPNHR0/v3O3ZxGpw8Yey/Neym/BgQSnOHuK0hOGo2Jx0yJxOWnIHyos5Axk/QAQ
nKMNwjBWzTkIEx/eOyl/uz7cd6Ttye/jCxlgrS4m3KZAV438PfWQNeUPvfpatJq7
uBGlrK/llc+NpDs3GTou9+KWKrmPKR1Rby1hqRP8rXlHDSrdhTu54/KuHEVaNlPQ
VDi+8sCvr4A9EOaAOIwzO01z0VJ811jtOCdceDHOHy+mMlWMyD7x14Xsj6LVhNGx
N7desvsGzGyYZcHWQujhZJKqPWRY0KxuQayHDr8SE/VYLMtWWOQGPL3ZVia2K/Ao
bD3Dc/ag5vDysgUw8tJ3lkAjmor0sYbgsE8tAqIvJGsdlCDojnSt+mCXXI6ylOTL
uzaM3QGIXPgUWNYnS8zZqlB8lncPc5ffNSe9bM0UVPYNXHOuR2JvHNPcyAABZxA9
nCpy6nOXpZlaDJn/5AzC6BstEuGZD9AagBv69Yzd9PdeOFfObbDe+tcNgNX3iTpD
Ajmg2yXFr6nPgVa5VhDEi9I4pGBequSQe6lB9VJSnlxDAV1icPF5K5yA0p/7rWJj
t9ZX926lPhjTqsNnNIhCpZvgq5O+PzJZhMz6AiiCqXUacat4vwmsY67S4AcpvbRg
L8oI+557JI7mYBwNrTp9UxuZthqmWchgGzYChdz1pdhYdB8PHqMYNOWBAZDECf8t
8YNPhX+31aOLGIHx3FTpoGXhVeYBzscFeapD6BQ7XuZE9mf2IwDepWMq0gm2i4T3
QwLNHS5bUe+HSF/fKqgnJ2ytYFxL8GEYw/VQnH75KYeKZQ5429i8Pr48Mu5u7Dm4
1M1We58WLzNCjfK2d+mmonIIB1f21QhQqN7iYPQ1zB3afRZPQ32o0QZ+Rw5yjVK8
RC94lvRKysiY9I5jQXt/AkdHSZFksF1g108KSZqt62cws/iwk070q6YRSSLPYYcf
tpGM36IUwBhVl2kWskCFfn779B2zdvg9A6i2ipTGVPzff3omVcRw/F5/hMcTbJP8
1Si/XCMvJ8AAn2OSZ4Z/kNz1bDNHaM+4NOFvPs33Dghn0HOU2OVqFYsJyHBtDUoF
szoeBsbxkz6idA2x3/uxYqY1nrTkfY3pwRux6K1dNLCsTZno2qaiTQhMkAXF1qcA
y4ZAHe5UX8ZZ2qN0JPWTCbu79zosQoZ9CEsJcyDz0bZreJuGDfm1ZZDfRTqKkJJE
lUAwBo1gZxymSmxHBn6idrKLI88P02FJpX8Sn11gD2cJMigUno3cYoao8PbkkdOr
z+U9aJqI/WkVAHbA5c9lZ0k0gQAGvjLZQoqR3GqHxZ5yO7OaHy6E+7+qXe6P/Jpx
n2AqKmdONdeqs6lVBmi2GZaqJ4aYzDW6/Fqspx15Sb4U1Zp509aOlK6XIvmxNHNi
tAZme5DEhJHXWEwPvus3hP34vpn4zUSUsiWW/2piWu9aTHLvol759zBTYj4qkawU
STRc38Oqoq25/U3jd5pVR4PWLu7iUk8H1ycfEq9Pg/IzFHy0LvUVNQNyfLwmteXK
1CSjsYo/+5dFSkv8yzQr65XQa/qHzxmvtaGKZe/4wDUVjcIpT+aekhN35la0O3+k
0vsGYWW+3BoGYlLcqJXwin5Rn/LNzJrSjFXxFswr7HrSjWnnzylYYYXdm8bpqgBT
0qm8RAMjVhxRR2BeMB4WxYcZD3gG+Evd/T748DfRM4kTvjt6lDp0yqq+JMg47V2H
PjNkXgtthZN8vr4Tm4GXQLnm0aUxZgskQJo9g0xze8XsQzoMnZCIgiRO/U0P5gjK
yQhNV9ADuwS/guWPQCDs6xLcOlF7suvsKuKr60HogW8KQfQ7L0/GUvA9Q8VRVPS1
/dHQvnUJXvqiqGIfQOETw19baxEW43fKr9DTaMMNaHvoqDKEOjwhsu34kvREEX6N
30YLXv9OdY+wjvswhLkMm9njH0JQy7ja6sW9/tna05EJHzg8uxVtWHrgM9+wZ6VZ
3fUSRdufQcNQ46QTy6IPekByKaonEYH2h287oJiOKkQYfAq1BBLciPjpVZe2FZQV
zVarDR8JhFzRA7ySILl3QooiZBLfCZhkdqqnp6/kmCuOurJXG4bp+x0o0urXZGbO
QFotde4n4GnLNqP0GCsUyTFIgGbBoot4tHPTiNbERCJD33TbGr+L4VCNEA1ta9CP
uwFLJdThXphj5sJLK6/AfZ6HuTEp9nwxUOaCN792XmXFVBKQIST8/zP0QndhUztb
tUJNjceUnIHg5VY/eSytBpkTLwb+s3Y8l0CWS/tLiiLv3l1wjc9u8RQsJcRhGS4W
jD67hFjzhd12SWYS5FKPzUS9XS3MSpxYwWRYbXct2I5zvSwh4j5M9rdSbt4LINXZ
vAh4X7KgiJNE3i3pzXVVPhZVMgbJRMZOkq+pqw3u8EdMUu/ACG2x8632o2QVXH+e
RyKj/1rh8Co+cNcDFnk/fptqgjJXyt6WL5CrrsoyNi0bXKwGvmvTZQtE68JnSyxR
U64Th0a4v2Bp5unG4pw8wdrGrQelrkC56RORVBCXyiV0P34rk+/dqHQs2Sl0LxhL
9AZKQlL75wV7ulMn4ByRYiJT9MUtB7unn9GzRa/Yf1RQzf3aLy6xvEmBh+CsERr2
8ynIgSrLujGk4JesoiLS1hDcnmZLcQz7e0FetfT9IkjLQ9zjzFUZ5z4k8uEmLiS3
CCo9gGkZaCxUs9WJuNAuVSgjco9AlRHuAFXKYV57b4xbVhFVqUdBt8ZVJr7A54Jj
1M/EJK2eMtldei945xXYeV2rU1tah7lpEQmXuhmFk1j2PrR3WfWPZZL55kw6SuMa
y87n3m/+Ok6EHR0fVaWlMSs8cIu7ZkguzgVnFzoBqXocKfMiJ8miMBarvZtHiJ24
8O7PMaY85iXw+FzQFpT5wUu/iXVu4GuZyOD4IzcvosYFpBTrB+nOWHS2ZvtfaK7q
c8tMfTzdSOrwOX5XdMVkuCTer/zJMXUuAZaZu9+dsSGqtoo2fBQXsqkCNx3gSTLg
/6s4UqDGOeQgkiYJ0ofFRK/k0sPw++c6gReDXSyXf+u3Pmlsenl5Z4flVfnYXzqM
8yZ4zkOvgomZZZLOQUKyUtDuMupmId0b08wKllgmFpVcJvTJkx8ZRAbDbKN7+Otn
Ur2nA4ymjpVD2DdXuQ/zV2sq29Gqm22rkNw36FK9IVf8+bFwvUBKrSBNhM9Vu0Q9
j5rsG1gESlGkV4X9mVE1862zUG5nctaBVThu1Rp0ALc+rdHL7GrTmsTSFQb81iDr
B2faZmVn44ZhAk8lDNycdBh3CgaEj7Rbq0im6wPqMMPpiMSiGF1RyMWG7NkljNUg
LVZAvE4e6qqigThHrsWJZrXxPnULp/WA4nGIBJRaVvBeBVEs6/nltwGKSzfBHrxa
EEdcZu4sxWlVoz4taBbWlf2pxMOd3cDqwH5TswcYK/uBfWUR7g1Slj/ZgPQ+guKD
Pu0YN+HLr6hL7iTw4I/jimrJMBRwPUPfelMiHu76fAf7oA5gGHnCzORijEUgQqKM
6Mq12AWz5pepXIGPGGPe/GEUOMga3ZIHExtDyzfY0MYoeVXX1UwQrBnEmjcDkJBa
nkdQhtMLWb3tpeS/5ypb/pFIQPTEmhEhs9yOXABthV3qkHZywcwlLvNMH1vGEn8A
B7Icqgiq6dB2G7nUuy61peIkW/vQmlassCq/OcBEBqQs+/GQKlZL3eq9OqwAUJhD
T2zVi87oFkE43I9IL/bW/icAaHi4NoRoK40yC9jiSrn6vq61PYquQwBi4HWLB/ez
sk25noVlEmPnCfbPr9z2CBtQAwIh2Ocr3aiDlkiGyLJXm4Szob5gd/uXABtO5d6K
RoXG4ZUenbQ9JK+mzI2aRZ5UfObjo26wprD3LcmS3UA/ebnb2IFJdGpVocvK+B6d
yR2FYWUactGDRQ4J5SlV4gQzwbv68yoZO6xW9jekEamJSF2yT2o2beIsx15uefxQ
BgUWMz70z4yxEjvfGkIZE8BJdBtm/IcIerAYltpe9SOTYtBOXWihEx+ZSYP/qRy+
N6wShIzY8bKjUqDxQbPdgG25T7oabV2/ibo9k4RPJdjUQIYPP1E4FmuriM2DYp3j
LhT7GgicZJlVNn/jARMSp8a34q7Cx7heDMCmoxkaixuap/6l/o0PsKqRHy/G1QyD
35LTrUQKrxV22U7Q0ytBTEcc9Gx+YJsD34Wm6yUDSeVcmAzCh8y6G8iAcuX1PreU
vgB0ox5SuIjGILTHF0XDoQ9qPEo9XuSag8ZVUte82Hx0llukpnL1EiHKGibVUfNi
Gbjp7YPhrXeW94HB/4c+FUb7yXFpjqS2W1+DGSlGx3aamvic/kuzx8vEtFHY+IxG
92ztXfZcP5qOty0rXREEET7VfOmT7YwdSNqS2PcHisg48r5wHawqc9h+AFWj8iJE
7iptG9SEyKbOW3ZnW8HdHhyOx7gi1Zn85IdERAHHQ9FhLEyW6OCaWveXJwbLaSfz
i/2HEYLF1YYYrQklvDtuq409iZRspLmmZuL/tc4AgI9tlSY1sfieOh3qefr/ATFx
F2pavMRaz6RlfJf7H24AUqozdnmjXflHDBf0Pmh5kSeHcnhEAaFGbUWQj1rpZZk/
M9fDIGBtr66Ohsom1W7CZZGAq+aASJSChBogdHuj89wG5wdqlbpaEqVKkMLlJ3mS
XePSyuCDn8mOr9r+0YLszTRVhxhuRgvE0iRn2Is5p5+cs+lcY+Dx38MnB4GTr7f0
b1die3gGeR8k0KYMFqYTMmdQOEL3fGgZdKp9kTazgfnNEQ71HPYMJls41oB/DMHP
9atzw8AwCrccbzynBooSLkJx0EZYry/oeqHIrInNCBPwosKmdFJLarjPmD1FJNzk
t+j/9CfqgiAY5Gq4bQ98yOyvYNRXC7mm424vqgOPiEYqqcuUF3QTScUr2g4jk1wd
8REtozI3Eo09zrVeCu9iTILkfIs1JDHW7uaiDq9/glg2oMJHlTQcAvy125PfKYEO
YMiZ8jqBw2fOQvmhUcr3z2dHX7CiTSgfFekz/3g5yDRaOSKq314qhxqMVxWzSpsA
jYtIy95Yh7jN/CyoNgIvyZ3B9hL4pE/w1yvoGfSC/xfgfaSshdFKqmLCk4om+FnX
23uBhj74OfvHQ2iV+ufXB7VFq/jHZbkVf/mU/pTuounPdoG7zZ9BB0UoAKUBF8X5
qAjZHH91dvB3eD8DIlI72p+LqUjmd18wgjEwBDO/VNtUyZpT/1ytGObDh0UQE5zi
R3GD817qXOPOJlZErdyfbmRfz0Ih2C79mSELxfzpgi/YTHONib8Djd38EAsiSyeB
gao54Y1y/BSsw+aDzsTqlvQtwYfWwddHQOCb49rIJ/QS/Q9G/L8f4c5dpcWPo51N
nMvVrRwsww/PXL2UawB3VV1LD0sOazIW/8c9ocDAHucny2P97mWCCqOya7ySsIY7
4Fn8YbnBrrvFA9GlyGj/MIutZsdq3SBY2JgC/XWQHrWGJi9cLKSq73nSdAUxFHKa
i7kmZe3cQiwx2zPRs0WygPtjff25od3jesrd55ljwExKjU80HUqljrsL1BCNZyKb
8KDT3PHSjlFu30khGmz8kNHMzI9ETdE5Mfe2N3fuP1C6uRfbK12bHRLOen+Jzm1L
8tpIhXEDlEtRNWTd+WWJtKcI6ZVPZ0duSTu6ZHNGmxOP3MznmfO8mVVD3YjXqK2R
02Kh3iKZuEMQPXuNR9AJiur1CLC6F5CVJIE6AMWScAShf7qBmTXnDH860eAS4jRO
Q3H8t0z2lVbvh06F0+oY2cpN8qCLEdXFzWwbP1zen6TOridw2uma9VPVthbslEc2
kUYtJkLZuw2IhotyATv7rmTCGguFzfbVsEnV2Ogx9MvXFTPw1APM5CLLsoCUPGAd
udU3E3GStkFt0wzf6PYLRfpwDz5p2pI8FXLaTR6IOe+5yAuwK1z4jL9wtTZQ2jS1
MKX2//lunR3VH6pMvHYzhl42NxRdvr7MLFzyl5XxQ2u2qxIgTp5m+ZY8jXHoOoEl
M+r/1rrnpxbSWrDrGmPo1HtiLYA/EJNmPpmOdkhZxyGHzBfDXDHtEN7kyaqbKKSJ
w0HoJGL9WmNGMbJcOG3e/W++Zc6XThELDEGTcyGbImbEZ4OX/IT5VtBJPKKs0xRD
ZE9boc310HQYF+RnB2cP2J9ukNDo+Fr5lDln/0/1F7cqJZNbYe1zyzOMxUxPVDdQ
TWeaPT2907qO40I517QO1LeoAowXFgk2DXEjsOzTAixPplMJpw+25EjJJVNf7fBs
l0wzK1ZReZWDcQJlF8FVD3Q4OYX9lw0axQwwQTQo6SZkrT5f78HVYal9Y+TfXpcd
bZhI1LteaKMljQj/BQ3iSxGgX5aFuJ5pjczJHSayQc9/TO/j47LfMnWN3pPLj8m3
ptX75Y3K3J/wAmlrELZ6mZB57EX0QHCAY2Ku9c++Lbf6WobumliyjMS9hinT86Dn
ZBObA3SFMi36iOBXCOH3mHQPvNTT0esglJW095WifLvWNftyy83rYGPuRdAupqsE
KspT20XeEAz9kjcQASyAYpYIGnwXif7sMTnJ8oEb6RzoNso82AVYGOSDvFhTwNy0
dqevc/9vMPRh2M4gjkbpq/7fybVB4tzaKEZ0zjAvnVnFrFIIkuNmgwjrXZHCs0xU
ejXK9VzjctXrnmsp7fy2vxkHPfdoqIQ+apefVHnPzBkQuQCK0F8hiMdvIkTrA3UL
aQPZu6DQTuSgQqBOkegY+CI8IFs+P4dsWr5awcJk7J3A69T/I8kfXyZtq5JPLHjl
/6WtKhZY+WF4VuUTJd3hdmZkHLwKgtAVhuBDLpusUSBQLl4G3RJJpzBWL+tJpZhk
VhwE9x5JlX63r14bHIRZAAlkPftDSwgK5+qRsflMEhpGcGLJNUUr2pNV3rLrblAt
Qv+X6qspsVpy8uA5v4yH2FEL7/U44MvvHZa+gQAE82iE8b7RkNdIv9JsN4IbZZHs
NZT77OnqBUN31L19vFyzf3zCPB6n5J9TSGNhu9glk2iMNgeyiPUOwD0vQvVdtJKr
8HVpEHqtjGGi3nDLqn/gbDESQEItOI7qhldNMDiw19zUM06p1CaQJfZpyheUBMe1
Jsv5WEPbYNkJPsWqMta/OsNthv/SlINGRwk8UHJjz2MsD8Qx1LleL7HCZiG7NLsp
j2duJhTMNbqjKvFIAZMzgSj/uyXC0sv3CssD1RG6dW5klfzapVhVZXTIM+ZL7Qjs
x8+jIm7ZpD6teKQw8TfONHqY08hAs6olRhY9smlDh3wcLfsBzdgBUeSUHcKHs7nL
UD7hxZYbr+9mVNgA0VCdcADkBCRD/o5a/s4X3EwFZc9jRLkOFZxunlXu/aKCt6SF
8c6hRsZhporVF5Frt+xYcD1qnjFax5Tsae2X9BNhwE1K3fddbKMkAaMdXnqslyVU
HDDNeNyOMCbBmiWZHXN9dxS6oLwh8D1BB9dHLlX5/uCNAz1P2wnIxaq6RgPGyJJV
vBBMonWZpuKOl3edDfTpYJqLRGL0oKJT4V9bzD0XYHN4QYBwxp8sGC7X2vbj7e0+
LZmFQOwjuFq8eVr2Dd3oueY+qXtFJq0bL4JhULZCoX6WXRAx27+e0BmPV0nxlR1Z
BdANzPb6/ZvpTdASVMylk2aluQlYlDBb5+fx2w7pBQqLI5TKDq8p8Kv59D+PNNri
RCDBuLC8orBeXXUdpiOhqKvNdnnh1YDlWtt3stimj9IPcdhacov3Q2emQt5Rnm3X
20mTbsr368zIi0zBl06HbK0xzMiAd2YKPI3dIkxu/Mgq3oin61j9TWGo3b7FuMrv
mjs07oHn/KkqbJCm0SZ99s8a/gf8Db3UpmQN0YDsgA6oilK0Z3OH/Yr2YU7K8oXQ
elWegFxow6h9vuqdVrkEIPfKFXHq2x3iKTHaeD4DoqiUaJkobBVwWJEhQcA4F5Ce
Xm6FuhDgNv4f+dMcgHb5r2ZRn5BVto/3Dg5aVeXfHEnUREcMsg+xYczFmvYZBP/O
QT6n+D7U3pdSN1NJnoaRKHvi7JrvziFBgxWSmoiAqqMJXnXD7H+i1cRNc7nsnhxl
q3+TAp+spWeoQBnV/LNzlZ7HlVkbHBZMfZvazw5JUMoS6PMOTzoHhfNxwWbyngZD
rCYEe4iYFfpCCrolzBR2D71NenWOjkIG2BwzoZaf3H3aveucgu0JUtbq4c9qRxjp
2opWtn+TDIu1eSYDCqx8AKjL3/WRFYKHSSc7X6527/9aNSR3S+6mH0tAl5RL1TN1
Vf0QTFFyRS5xgVsd85iw+3lNoYueDlclhgwOs3wjV+Q7aaY0qAXzrpqkq9VvCceV
vB5B2N35Api75e8LtuLIBuxmLoHyUAWfRNKiMbx+36VNOXLFuhUrcyVDgs2pSZW/
WKbvfFwyLvg9zWG6dXMX/YhViACKRJPxAmSNra9IaylUeNxS6Gu5lsnuZCCc43ol
/Q0ScQTh74vBPp6QsrDuxFuUjT4/CXhFbkcJf5ujU8lNAYMEkQQGn30NBa28pf5A
+6sKlAf746fbNtyZV41HsoBsPiZqONYGUcGKAiB0n/sN1xCEo9Ht/lynOuMP9t54
wLZ/wTQcRULcXJn3PFc6fDdWcjB+LYN6/Rjw5e54KE4z/OQ0mtlWVetZN20kNO3k
Rwh7b+w310WlT+rKVaB0LV1Oy+aXmyF/A12d/TFN9idaEScjTIwOT/v/UXrC1B1/
rOdJ+KCRYgm/sVZEJtQb4/CJRBMrq3AXZHV26tiT36yOWjSn7X76XOTrQHxC3aBW
b4JUjoOYsXv9thLlJAbIB5xW0ZQHY5tVILH3drraPZL0bywBN7aImw2ln+aAQCrv
UDd61eypaWGr2sc+3PJdCsKKQiBYcnOl/ecs95n7S+XhpgjmRWjHeHLMHqIjcK1F
m9B3sbl58lbtcEVDlwDJZu3Yg/TLza9Vo+d0PcMUn2DrDI5n7kOXEqKcMT4f0UYZ
iWVib6UaRk7ppep12o1h4MHwKI3Oh7haLDJtO1vUCTU8luKi5KN41Mvh8shfQIIe
rtAmPe7yM0yCXGx8v93tSOqTYJyXreRGJHeeYgbyOsJgTcmAMlFsL2tZc5Sh0kq3
uTgK24UBwjy28oXxCw4EwXHWvkLyud9ntZDtM8zIEeXFMozhCi1SlHVLpTzhLM6n
6cGQ2cVZD/kU3x8AmXz/9VExLkKzCzUO0peAs4geMdX0RhNBhtjqxJ9RClFENHfv
xYGf7DtDW7BxtEtM0LdjgH8Om67exLnEqMimrYpINCBwY2kMPWiL0LzfsEJ8gZkk
w+eCXn/PGm97oI1HXE9FT2Ll6X7Qq97ERBx156jVfzji+2iIaCXxAWiNlgjXk+jy
qUnA/FcruEaDWTSaMGWfrart6qodgbya2QtePNzYmXC9kF3YHNu21HnflGJINfu8
puvL6cDPKt5UsKPW3KtfbBSKNFuQFitTYygdsVTrXp8NTsgRSjEaA2okCJVq68Ci
EnDEbBHp9U6JW9oKtlKXlkJ0/LdWXu/wMV28GUYyw1m229Wm93hGZkZnJVAtzDTe
MVM1mNETG5p6RyRsdesHQh1OC4UJp3I48VO+JRLhdZNubQ6c0tKo1n8JZUQ3kRDR
/A0aovbqhJtjGzmFYlHQuFi/RpK0aSisgeHfZFhwe1jmA8FjQqccO5+Ut+xqIxPu
eCYhJVlPVq1wRRiZGajbTVOHXgKoJ0nArTK9D/Te0aj16YFz1TqHfCM87kplJAiW
t1zxJGJLDIkwhcYawbLPg4ub3yZ6hz4qzYuB3qNua9Od6iEwFJiTNyygk3nK6Dud
w94S5XpJLYfBNNOsOYlFDEPhpp6KADRsALREps/lBOR2g6qR4UvwpBW+hcJE3EU7
MA1F3nSHJVaQUAOoVX4MXhgqZ2hOhKjq1rqPneBDRqc4MQ8knK5Uo+c4tMJHVBwf
a4GXxSoz0S7s8ggldA5BRr5nsleK1zwBD/CAoQAxgHCY4zu+KqZpZXcjMSnXTtmN
2qHGRXIn08pIbkpZMNccbXJRE2MACxhn8cm5K/dI09707NEf/2OBNPYpw5lxPPkj
DvtWmFEGCCq6+i9sU47k3Xzqrx9Vr8iav6vvSoJYs83DLVTrNryrDHAroXJAFzGU
f+pIU2qakp13w5JzwVpXf5+txhvzqFqmzqQddkI5wwTuu/+fH/CXz8tmmFoDKnow
n5q8C/VqXiJyqeltm/Xi4aqUGjHTXHgJD262YmzrDOO+EjM6yv1qshhFYr0vapi2
GUEWTsgV2f+s7/okXGjepoRRtP7Qt0NqNIj1igrZUBhe64Yp/oDvQxmLGeyv2Zzd
c/o3FpAlwhCx4HLiZFOjszSosdusvQ/BUGhGEmkOFVOc2w78/ndWka1V1LINSUzv
CtJ/u8fTs6Rw1CEoEeDQfcd4+pDZsBC6cO7y7pN56tqd1ZTg2fEluOHCPB73sr1o
5WP8bqTm+HX7zaKZl2kupMTsD4z4ZOMzUc/p5Waw62X0Jb5HjV+oxCqd5ZCv9/aA
j96etKlOFO5OTTC3ADgjwTCwywYPHEPjigMlDTleUNTFDtf+UftUzEYRU5q1w8xT
Rjr7ORU55tvD3uhb2iSPAvA0CRRv6nzUmsVJivhtZod3o60MuMdxpNp1RHLSks9x
W4NZzscXc5qqsiq41XwkfhoFB7qzJFG0mRcfY38CXf3mc85g9XZWK84C02jZWd9D
TgaVgowRfLYFIPDifFUvow5rnXDPfFPM7alyv6lNCdqGNfQf9LuAKOU/2BaFny1y
tMjv2n2YxkFHl+7a8fq5n4i9ubgarniUB2mulU4Jz9n8beMZTVuMSWaoLLE6Ihbp
M4fgZJh/fiD9viJ5IjOwmNaB/yg9k0csVguNFbacnIU1mp8KYF7A3UbMV3gTGZKi
zexru8I9PvT5YNEX1z31r+DBqHfX02MQiJU3sk08+LWT0NAPFmdH45xCqSc87Qj/
GvXra0ClOi+lf9zVdl0OItrTzr+FjKbTiIHjs//HhypEeNza8d1DT/uIxo13Xfjm
+b/c9aTqCP0kQXC5zH4o4ShpR7deAl4+1ieFrRd+CeislbJK5QAjN5u9R1TerjhD
QKK35TbPbdu4wMfKIavH0uZsmiVeJMe1XdBCtludkXeetnT0+Kz78acQUfN7wZml
rILF7O/HYILE24TKmnkPogvMTt1DmHdF/RwC7KoF5KS7GVKstgU01K7IvxjcIpdV
kZ1fuUcnJw06DrnxKoD5/Bf6c2dLRIXZ8C85PkeIJySIhVGBgJwDgVQVCopjCU5I
eCBMORTpS3BQGoxYnXAPqezM4nA2LaBY1Z2q5X5qxWTj9fuoWXGT+180gDTCv2yJ
QHSGqZ84gfi6LOEvjLwPwO0Hy6TnGxFSQLEamE8RY7m1upHDWRIWTDJY7YP2Hfw8
Y1JS5ju9D47dWZj9rS80sBmjvQAeZTEGm1kUCv2qlOE3q41n6paWy+7XO6ldY/2G
r3N4tiWKSIgtSwHJg/V9550jNxpj5p4z+SzFYyFksFzXhbSfOMUm1jDmLHfgQb7x
WBaRpCk9f9EGh2rO7OZvWTukdEAGmcxsaLkVaPC2NYdoqvh16kcAi8Hj2OflFvFp
vO9HBlit01kjD8pzN++EEI3vN7fmyv/250U1XrGBUNdFV7X8lKO6Qw3u4qd0R6eZ
exxVl27Waujx+59h/SVmd8XQH8tuBIZK7jsW2Pfdws6ukLj0rV09B93wlcElgIYC
JdbUGXsi5WRhHVcJ5jlI2bMYtxqRZJbkmfLM5RBMlH9iIrZxCnoyt1OnZcPkAivc
qL6Nib1xlqf5jqSiM+YnbLUdwMmjGViZK9Rn3cYPejS4vg1AIEY367vTH7nstOo7
CJfR0SawmrWalytOQJduuFypEa3H4R5Amy+FZ2lvXqlblFXNFcdFMBdGcr4/s6ph
YldianJqe5CZ6b82qGH2FYgenAvn19lZB1fb/xB0+5GWAX5OPPJTcVhagmA1fYpP
HICPYr8qE2J8yFF/kyN8yB/zlUrd5uEI3oEKZbpSfb03bOkq6EmNjtLPo0ocvuSy
IwvPFEIRg5e80HWCzXXnG20XVeGvz0n+F2Vtc+dOok61Td4hv4vC5uNmYbPvxG+r
PeDtaaeDDsC+K3n0YToAq9fGUOCh8lxCI0BP8/V0qcoOHkNQ+6/4UdIKHuqtGAPX
mn36wljNfz5HjpOmSzW8gtaRMjn0qSt8AB6a/M7bfGLJrO/fiyLipHP9cxfQEEhW
qUFZXh2ekENcIwPhagmA0NlFU8zgzP+9GP4MzIalb7VMz1hRld0QJ30rKvL01eb1
9R5TTl3Nh6gcmGzSqZFzOgDsgnW2KDDR1NE2/Z51xySR8Dl7fNunHwIGCFIJzP+P
eBFVl4ZbpNx/spjOc2QXg7wi1OLliqQZgo5jbdmZzOKx347d25bzC2MAkZcNfdYl
mixUD2/bcfHJgBeqGtvgUY/lgCUDDRAPAPp970Pr1GlhvNilIxi+CzX9TESxu3Ru
BwC94t5xCMpfvnyVps78KmjiIBADjc0okV67UVb0xxOcj6cvSBySMrBnNOLAM3j1
Bch0g+OB1BzRJKnt1ucj0Pu4np/Cz+eciLN90SJezYZP9yKKw93FuFfbTHAVZ2D4
zJb1oIQwbnP5+FTrgYoVRbvFJzSjgI1tTT2lf01yOGrI0F+cT8Gol1ZJ2oNlHxBJ
MWltPy4dKXImPiKYPdGKNx0Y57n3yXWV1hoLP2RWVR3ZhQKrZAuNWwwut4tni5eX
cgGK+ilou8amNxHJrHtEk3plOAsQANPS5P+dHqxIiuSoutuIo01YykJWbpR0N39E
rWmEReaqBj16mHhXlabkW1nQkxBbzLl6MrJqqkgYQVNJWzAFI3Y0YZ75XTGgJ5Fy
8h441XT41eF5QN5XYHB3tB45H/lysUnxTN8+u7nnjd7E6wdmi5L8zK3C/N5XUNhV
KWmkmSFUE0j7JSouhW08IhNbWfolG2kpp1xFWoyki8bXf2RHoD+QmJlPb/RTR8ZU
bjxw3uHYmkuRtV7s4S/rsI5TAt8eS9WVPMwzwksBB3a7F2RDpGwU+zToq6dVfWdI
rX3f4BBwbwVH+Tf+1J0Q4z7JuXNRM+KARtnyZsjfWcJ57ujUpLw+ogbYGTT3A0uN
/iIjJtzG8Zqh3EpArpMNgIupBUe45yrVutreZ4Y20H5LL9NjGSa3L6hKnbPUClK1
7uNu6zdbSsdLzhGmdJuegKesmSdpKVlKR7zGbKjjOJ2qhfiDLxBuBQcuLFec6+rl
dbDsjJ9Fx6Ux0PsF0xg0zINZNc1q6qfukeF4u5v5juNt+BHBlhwu7OxfsQFJXlMr
Fdv4egMsO/eMvKAjqTqxONLnTsHLfQIsUkfg6UYu/nl6vHo+vMY3royvj8uwcCZd
x8NYbwuAQ2XW3rWQfwmc86SQgL2VXSPF2NFruEf3X767LknzBccDV3qSphvyFmu+
71vZtdt/EnwcR1gQaBhQyCceTNg92OAEdro29DDsQyO1SZKG3iuOSsJeHeFOub6Z
Yq1u6/+j7X8H5GuU1fRVJzbXWnuxtdm8riHlOOW4k8F6Nn69ePwDVpzBuhbsApS+
EJVZNu233YQwsDNxTJ67ZCN7Z51nkH8R16JOmX9StZcfc/PW6N4erLjGO9YtUvYe
40ZoAOLYPvJrGbm6MmqUgSXp0GVaZ5LWVwJfhcPCoB2zCzBWGTPQguQv39XKT/Sh
CkLzwKnYaFwaar40fL4oc0RvDoD0k/q/mXKURb/HltbHHwvjZoegSlw+vXAsRwUj
jix3n6KmiB1o5H4oJZufGAa4vAf62E1wmxPfZjFkGyCRQlzS3clhcTSUI8Q6zbf8
zfkO/8zwn6RGZgxFUyRsD6VeqL3/HLm9OVvJxjbq6rlu1jWzcrEIoVFbYwzpMGix
TpoLdN/6saspqaRh4araLBx4jz6a5mjAGmyovKefyWjWw88yTrGCOwxFWGbRkQOm
dPtdtpzEbWSAE+0xijOSiVDdnsQwJTy+OSm/If/wOmb6yUkYx5/dGnA4jSxptwcq
54FjvUg1buh++3aebTr7S944xDo+qilozICwfVxsb8Zk9YfmJE5pTsmLzBtsiDZg
WIh0EoYc6xwpLqg3op4EYSZmD09mmzExNcIKFz86Z7av0Ed6fx//EQL1K+g3P31K
ifZWeS771cfeRkZGJ7V2ePwA7tGAaujj+mc4SSQZAcPiAoXW2e2U1PeXjB5OdwRQ
VASu+/UVnLGCrk3R6bpaq7wEFPtMPKFMYNj9+j7aBGCYBaamj1Nn3odevWrPrZCf
q0mpPmUb64WVUktmoc0GiBCV3mLAnZspfV/uSIET74gLuXny2tQkgND2HzUb+ME4
RJeguoJEXmQToL2r7SiRmdbGQtGpt+6OWPjlE7lMwUrh77UPgG5PPcuZdH7x6vKJ
utawwcNP9CIU2jeS0Ok2/nVD17mD6fI58CibpIvMr4yvZZll1EtKlFgNzkEvSG2A
RHbi8BnSBOdNIr3iq8M/PxtIgxFdEFLlmy8DZ3+hBxLujir6pJIEDEJNzHJnD3BD
3VVrxHp9ZfQYASzGHUGQbVEWxPc0wkbS6Sv1x+iHiWL65B5Ccw/RI5UbX64f3yFe
T+Gn8VCdSPR4O0lwVhkeV3wll05n3OsBC1CSn1tLnR4qZtdEd08BaHEdm6ecPs8n
OpSKufHHi2vL8C29fne1qmYmFfTS5BbAiP+2MT9+4D1p5P6MZJwdJwqzoOgq3Bfw
jpngIIEnratqwV5bmxYMAfQVdURyl0shFXA0a3ruYgHSeakzZkUmCj4uSs36ekFS
xTQcSvx7LhZDDW+se6pRROllRvCudlNPyPC69OxVs/Hw71mF6OKVO6iuzxjMM3yZ
YFVG1iN/KsU77227UqbskLxM7BgO/bVBNEcTi8fHljv6pDAKzQLFBLh7Ckfay74S
MN7VsCoktxUjbMLoptMLPV+kcT8/4jcWbTj3Kc4RXbWQG6zGj67ACEo3ZX/zJ5ct
odmwC9j3m0vyw+mSQp29XgJEndwsaAxC0i+uOGK5jEiPmRs6bZOO0bDVJHuJQSx5
yHnY6vZwEps4wKRepq7wEb66gnrJz5fpEXYCTxPdyeZOjHpGqhIa4n2pMMJ91y1W
1cnN9hbH1EihWS0+EPXU26VClEbhF3B1LgC/4lS/2PxEmtiq93gTCW7FcpG2ncuj
/jwpeBoZdvDxGXPwyhaPX1+0GM/is/hpdAfomeXf+mtJ9uq2PINb8cvpFI2v5r3/
VmdEaaknvAuz5xa/+gmOVffTTeZKsWZ6P5PNjRr8JjTJEdufxBMq7mUFD49E0Okw
jF5bh45KUlAS+SrY7y0P2JipZF9FfXuoQIHUsBtHDdQ0COHZ35KI6O1YnhkxOeWJ
Pxqupy66jcw6/Ol3tUHMIw8FjOW8L7SRAOA6U/FbKndbG0KVMwJCeevKZs+4ze4z
SqCwqLJQxdDFV/pMxO/XGdItb1z1OvpMLObpjFmVfJY4en6TzidtFj8B7TdFFGtr
veJe3QMebl5jdMU7dLjE5jHYPcge08ge9cRA6uOczKaHLTPSvktAN/eGegwdWcAJ
9qb/J8o+m1HqZfCwxdOjsDTTpM64V+z60w0mGFsnZpj0LISkY06qDhJm5XdMr1fa
W1rLSQVKVt2fI5lUeeXoiC0KtsuskcvKwz4Z76X48iPhvsK8tUhJCrU2uVhBcAMV
hWP4IsBF6l3IHGS+CoTCmph2nkTwwOU6j+goZAiWQUJJmeGWqOrU+AYGA1mltClo
lOzbC+ffwz9mk6/3QRXCvTTIrxxFMZ5i9KoFBf5dC1UB81bMB/sOSMr5GY7WBHbM
LwuyVy4I1AULI4HEbzJctREPBVTGYopSrGqguEv6i+UsKG3xUP+xGXQhhMhSJ2+V
HB1ugmhqWjd+J2NgyAH7ZDQSpDzmI/ni9C7POc3QBriZZx14rYYN5mLgfIA1D7mY
AZeOX2r2bWzhhfMiM+Q8NbMPoxqNV6TEGgtihyPqx9SSmGQp0yniZ9/ctkaOgzxQ
ySMRLYeM3eYqaGXk199dZSM+SQDCKFxzpXPlSNnQF3VA8yyg64cVgcVf/cZqkl7K
OSPCuFqjqyB6b1crAljuZAm6VRsAbwX8tK/UaWeuQV5855gCAPqBuiqZrhrDvdRr
4TrgGJZsfIHbwyBjQeozDmCmGXc7JoxzOrzQ0UaNYm05i1GIDFLMWkSlfjd5nfTs
iDDg8pvXssV0Yp8Stxr/8bgsesYNDlK0XeZocVH/BBMW+Lm54CwcMDV4BiIe5MLM
D3Nq/h28GDlSaxT1r16Jst49S4BRMG1Bfe0YYBVgOQA3pbKP35Asb6r2ndsMyRMp
v0gDqaYDjEktZOtlIRTa0/b9TuSHqXql/oIckzZAx5xALiQabj9sUuP1FYPwck1A
Q3UgQnOKU1gexFfeC7OzzTIAIFL8am30Pcv8sudteAk7LmeyslkjOyRLJ2deG2iZ
tbfWqLEQqFRPQxpKhp4DYBWaD2jmudtl7FyeeS5GAP+NQeaGZxM3Syc62zjpBFVT
PqOt3So+SOGtzl+lhONgGyKL+paDzYf999nPho1rStJEN/HT+CnPGgCuVJb9GRwE
wZpqZk/fFrDKKevwEUxg5jmh36B6Qi9j3N+FWnpvfgRSw7yeGa90H9MyWp6x8jBs
yPZnTVYL/+Juuja6R6IPa5/Tryza0yPFajBpInPB4Bnkb61mwEq5Tl092Jc1ObYR
7F14GHFQdPv0zGX22EVx8DjkD6n33eukKolU2VUd1cuGKUZI0ury4z1YR23MNMLW
eu1IeLz8SaVRlV4vBvUVsxg9ceUrlXbIUF2uVhhlUcv04TQc7wda1yZDl7s1XYuI
LTVFpkTW6OOQQWrfTWhJZ3M47vxitQWTp3TepaJKoZPRKB2oZqeiV/YbCsAe/mbG
FX+HNKorDcS03BojZEOFGJ8fxfK9gR9Vpwxtm/qeP1l9oKOSmrPzGGzgL3xtFjhO
2UcFLn7wcagr7YCM01UxFH0eyUXb5+HCu6vLzm1MJRt00poqk+zMLQNM3p+JOun1
T1n8ChnO5uJ5ZOqdb+3ZUc8XB0I8sb7eES4ayAsY8IDJ824b40xXjUwiUzWaQEXc
0voe5Z7sysLxC08LOdHd8xNQhYTeJFayTzxZHHUqVcCicv2H1MmiQRE5BL4ykpCX
zYDt/8FdKaGxuegx8xCMXt279n4cFPHSYFQudTHXYxGxSoqOJoBN2OPgIWz6W0F/
Vse9g9TjsnlKyeBWAmXuATLH+HEVVrXFvWOcUWYyvmt/Z6GV3/P8Dl5qUyzCY4mC
sZX0pVthymkzeSpnmcUOw53u+sXN8jwikyql3F6Li6MtT0AtQD+NYPsP1gCGZ69V
Zz1V/mmlUjiJc+jCHq1DNu0dhUxSdb59W/O249pLa74rp6RvcnxjWbJMm63X+Tdc
ZEsDdtIqi+5TFLU8kRA3dI5lJBZO1E4JqR77QMiAPxjZx0icKag7/o8sGpE4jv9K
VSleI5uiC8B1ePW7EE3dhdCJVlIMMGwWOUD9tq1eQOomlnLaWV1UsNhgBWFzyxIs
KE0DW6MfHl3GtHQUy53wqR0tCI0rdmtG7TJA69YdbkpOpClLPjkxUXrdpdt0Gr3x
XsYPWZBnW8ZP6mG1/NHTf1MNE5meu8JZ/RJ3aXpLnsqaC4YlTCktQ4kN+nZHo9q0
oLxeslqk/zjlNWCnH6Ckt31kScuqRk1bQyN6az2G8XgbLwT092GWo93PSMJmBwXk
RtSn3DzZ3PpYDYkFQLOfvqFQZWNIdpNIXOyZpg9RdlwC6jPJPzT/YlSLwSV3+y+k
+87eNUQUBEkyYjfNWuyTHB1itmYdFirK2R1U/ZdFZWe01PqxYWCP5r69CXA+RmBz
0Z2zKQ7bNbSxE8stNnX7rbT8IHlld54//D3+tPNodr/i+TA2vN+INit/UfdyegDL
e5xHM1VpvyLeiAbAInm8hl3xo39MjNbkBj2rgIxI0aNvhWdJqpJFDahh0RolK2q5
BXmuhPAgICrVkky/Cwct7yyztAkvFoGNsq191w+qBz/xy4NlwVHgGFp6jxiOXmgO
2Frp65/CRbibU0/lL282X5txr4vzx5J7Q/ueS0Cw/aLenDCcr502MRB6QLA3ejXj
vBaWB8aIaqynZu1J/+rmjciGgjoQ3VcQBWF9dzYPJPJ8VmKzYonj7GJtt4oJ5FTk
Kc0aeZ2FkODPV/uOQPX3/WlxWQSRv8elrabrNkx4s+CHrCgXmCiJGMOuE/lcGUEN
ciMmOfFbLlBAZ0fcV2ynM9ld2ujMrJKv54Q9VqfLI+sGZVj5WIuIIDqGNYhIzqyY
Sb6cPTofaO3ysY7shs4+80/CEFh8VueNkszziSnfhllwn4YebbL6Y8lgyCVke8B6
sylzYhbxexnjvHLgMP/fnPzp3yNsqe76P1viarZzRdtwbSKHTuFM2bu4hlSQv1ZG
9HbGHZ2kDSe3XaTlCIWeC0zdJU8KUEPvMxFsM58J71IFE2VAfujs6zXpKTyra5bh
Ta0hKBB9LruseMCh4p2mLLg+MBKtD7pegVxc6jozBWeuTCcFL5wWwTWDF3RTfX1o
G0kIjdAzJG997rEc4/+OwWj4Bt4PowiUW50/6HfjO5d5KHmTeR6twnl8/VkHkcC9
xh+HzJQmmqSRoh9ovKZiXQ5RPUceE3eNc6XDM3RVz6libL4sn7x9k2Hm3GDfSkn5
PeGFjG3c3qo9R8FPp6Z1/58zGbEe50CJ6z6MwNTBDiy5OlJFh0T92YWf3sMNPoOX
bSY/+Cm4jVCM9NdbnWkhd3DLlgbktLt4KsXBDqrOKg7KSsXFgZ+h7w02t2tLcYA4
cXfvH7CNQGfJIRVqLRRIqKz/OqeMqq5Ux2U4iCby/+O1YsqPAdyLDVJ6ktMyiyBP
49LyvX2GRNIeXwgnimW3PWT6VaCRamPIL8g2cvCn/nOv7umaUw5OVrZOKmnyux0E
Mo7idzZFuk0/4CzQhchFrcdsutDTPKHlLcCxeHk06joT04nsaraN5pCkT2T9nenD
wPXJSiGjkvTFbJjRCXjPFuV4qGQxpIU19JuDGdBDxuH5U+WK86wNWhhFGnKhdpf0
LF9ZeCH7w3+T8W8LX4lNeueCiI9pQ86jxeAggLligjj0CdJUD7V+eoZkhE/bW2jq
E69Df6btRzAaPCC5LjL4hno/Jd6tjMcIUHgNRLnH4otc9mRkuXGhDKn1vmyIVQ61
q7jw3b39gHuWd73Ln18KcJr4mUtoB/Htq6b+VfEwY5Io2yt4SkinWTT1ENKYsigV
vKP2ANwTGc0T4kuFxqUm/wExjHfQTqkk6xsasNaj1oH1uhA8MGJ04dYfA2sGUz/a
mVHzKXdMtPJBJbielttMBSGA6K4IVtcbYirLcShqU2S7KiVzqiG8d3tvqGZuqWdV
bFN+SMEO/+nEhStDjziA5/aIANLoFQNBQg22CplTvdA20yNqHbUt1FRmA37u0ZE9
1A3m7NWyY+phVj+/g5g9YtxxHgRsiNvjEZw3t8tO3tNQ67NYFYeDGFVEDOnU1xw9
CI7uGMceHmTsD3R5qHG8v/SQ4qKsh+3+Q9OXCvjSBjvsbBSHbf0WUk9u52zVIqXm
j2PqaFuadhtVP8GonXLYBsLfjBEQqPCYNzp8Pq8jPza1rTTWX8z40d6j8Th6oss6
93Hm9jrzbeZmwNAgmJ9Y5Z4mLYTPARnbUSgkLOBhmKvlnyH+R5h6sRAE3CjseXkb
7FFiqcjaSFnCNEb17CgOIMYr85gbKBtHadkYSjDWCAcTq5zgMx6ehEy8KB3l2fO1
5esWo2oc5PawmL9OlttB1pKonpRfsLMTHfc4Nl47x7RBEK2isKxguHHMaIZgoHwp
E1zcpQgq6BD48zEg3kJkE+0ZfDsosoCBOS8tMn++L4WdPqsvfHBhHRbSArllZgQe
3SRJ6/2Umg2UYfHjaZZ3ORtDbX4COYYID1NDkMVpfUkDzzpp5f+OYTrzecdbRJKk
GvMTkoVAQVEJLjRawtlcQT29Q3OOHyK/uhsFDaPLFFNnKvTEZDTcJcHYXfVC+aCg
beSQisTP0hvQuih9z0M2kYP4UNXiws2LoF5qA4Dp7M4ZRlawC+CjZ2VqIiU9J12g
BqDl1Y6uXbrIINVqNUfLcD0DfMB5CZptd00OdzaqQeu7i6yPzNVQJcZMyclqd9NU
ek/2gQeYQQNXBBtJDaRV6ItgmVYtB72IdtU99dhxYf5MpBDP4fPTQflHGJwHE9MC
nFx/bIQlbt7BB0VevftQ1Isw9RhH96TPzwxezq8exQvrvEjxQFUofi8AAmwmbQzk
ilNzAWrlUqMOvqdpGwZ3jDvXVoI/3OzpNWgzMIyO5CyKfEZPeyKRtAg0GN7X9yOk
eVOiFi7u3l3T7FpSS5851ZbRS6KvNWPtaoY+KHUk5bp3W0gUpphJqYhQrDEB/c0J
RoZSFZfOoUUOWSEeOEup1T76JXjbocuhaIFCUc3bg5bQvbj3xY90sF4i/+Jz7hG8
Oy5cdf7jTjIAUXfBwMWQPZPVnyZINPPxwkjkyNCBN6g7dZ2Td1QWsykWC17r2Pek
WpzcdaGw3lKMBW4WaNkXY5WbFaXmcGgts72F1fPbhW0uv0QPhX4GRfHJ3ifcHHNP
fgRLE8ehUFUYuQV75WjAY6acAh1CxtblUlE0DbZKA8sbc6l2DKqljRCSnPBiTFGo
ymJtGQPEsEXKTS5XXHYXwunSIlUjg3yoL9NjQLQmV5E4aLkfdKkSGC4YCA2k0f3A
KcixpBxX81h0A724ntdrRYf4xLnFsbAD1Mw3ihQx/5OnTZ6ZPkcNXOtumDx7eMUZ
e2Eh5mk4T4he42fEeJQ9pEwD8+AFVLMsA0SUml03GE0lfxeKRvvdiLwOKuN3mUGG
MCFw5mEvSfoyHyig59l3eNJ2nB0+5jVjbsMUZo0vBTf1or7JsrJdBJ4TbfFUZRlH
NBgOXKbUuEkzGkqu8lhoyfpdYSb//D/HEFl6LKWgsk+1/TZYdR3wA5tpc0hCT6IT
Cxpn7JjOMX5sfVFaZzsJSvGfEQUBtUclZBEYVuF3xuXicOYXJgkA7cnkw6M0M93g
MTVDsA42L8L6gKwk3DpoO5soXp35TKuDJONFF+BUAyCfQjJbYoGVmhGOBlBYiNjv
/0VDV+EruvWXXfptW29DBuqNL1S/6+2RNLnGmcvjvny6mHa8IhcpAxu4mpJX3Cll
rNLzLcagpb5Tk1fOFiIpVZaqooyIej3pLALXC0ltq5JG/y8wwvnfJtEqD84aM8W3
DWGW9otafaOeAhMXAgtG4zVou0IHbVvGvHuK8L65XBQsdDLhIs8XYIsFzRbkBvaM
xKbuExKfS9eWftg137uQoLLiSKHFkX6xdrb2WPeuH4jzAEWPQ82Ec2qi7RMDH9lS
QwK4VfWgAV4Flr9iH75Ijv9R73FEw24n5hz+4zC6QP39VSUBWzKOY/J4NTT3CrTM
pN/XZIbASxghuDqaUQFfMcbzSUXrUNQ0JDWQ7BVWCLTnKLxxghV7JPgDt2iRuYDc
QJTI5Xnk01epLQfxInqrl3gjPCpyMSQNBF5i8wEIRrIoHeTAphAo1RTg5DyhX+UX
H7z4hleyVn/DaTTu7TrGEpAqH9R9tDzGRMpK50WqDWsdX0amcj0M3nRAcWDmzftQ
dMKfAF63wHCYwwMBgkZxSLrbbVvFi6BjsKvjhMQAVysidIfBnKb2Zx7pRFoxgdvU
A1nN6L1frXdCGHidJSuCQ7w3bbruCHvWTHFBX3NYZGnP2FUcNfGjrPfuYxdJCAhB
gsNiW3YkWGNwojhtZsD3vLhZVf3g4rq9c2jHaYL0Oac0aP9KRbVHZmL+c6VWDY15
HDnRCuYaHhXNFBc4rxrEDMuB8/mYQ/6AJK6kUPvWFYFpH2Cc8F6PM2ppZNvRlQid
QYaTG/68XqlagMDpXrF5iNG33m8vbF1kCFdS3TskenWz7Wx/FJpwVNjVnjwl/8/O
se+KkdZPH1oh0IU5AKl4J5U3qm2kSb3HS2kJAgRj2IWYOlzp1MlF9Cl+S+3jdJ5x
rG72P4YMSD3s7QA0OjaXucWnUzTZgvruC4NlZYCy7bYXcIpvrFxAFG7A7BNxzbaE
ecitn1hX8t3G/Qx6asb0n8/+3MTu0aT6qa5QwFFDv8kGfIAN2kKDuKKVVB+qDrj2
EJIVD/fYBtA1PSBCo1mJAWNAhZ+TMCa9mTeSrUX8HvJ7t7DjV/7mtKJJr7bZ8n0z
ptXeUqtG1G3HBzt6SrNwWH4UdoBb/5XgsZBDJ7f8wnh/sQ5zHEOhkYCJH2olF4cm
szUq8px5PXd0v9jQW5D2ft9NPS5VM7FyNj+ANt805eDc24Y9tokbWS6yCTembrtk
5uZ4wTgLLuSz/Iq+UEzumW6amOG49+ieiDPPHcSPDxZp+Cq1Pm4EwHOXvvDZg0CL
YRVC7K0penly/NWbGlvRkmfVL5HtRwCPIIeQOhMVfwEaduJuVQ0FNyjG0FT67WRN
OJlC2FKADVwkUGnlLito0oDgLyMam8+Jg4FDf0KAnweWtVCLYGFWU33/RZIUf9Fk
zm+8698fQJfnpj9wV28ujrczT1HwyO431IhIpCaD50YKyv12LjiyXuGPFhdUNExE
iLG+aoHAK2kxvzryTL0FhzVQYlfGW7jTXrw1AniWF23SLgbfHl+FpUlaXAzqnAoT
S0NqnwPK/uISfrEHksFOhjs8gKAQlEEIalQFAmj1ZPFMHD5VJDpe2DAcOO66WQQE
6GXv6AqANSYt0UDzyqSPoE7P92O/YK0tJVT9GubYJgWdGlxwztYLj5Z/mtjpQnIV
t1jw62L1udIQbLA1Sllm7Gg0LockDPijS3A4q+ip3bfb//dFhje2NOCFjBPFkTGm
HmXkOdF7jyfd+hophoQI3gAVwpQvJrN7wO7VWTgxsKRTB9jSs4J5nCfUoVLgbO/F
y/OnRIl3vr6/RiCfiYpRbfV5nJGBmXZ+uA/IzcsbrEfG5a0VyGmiYSpMhG2dRCmC
Kfs3ijTtcFoHLS6S1xMmbyXVEBWBTcUFYY1D/96nE6DNf24OwBLqRf0j0NTWnNM6
s23KeN/a0SCzJUjJnvZAFFgnwr192jK/k7+Brg87c4HaFEzrbKEKs02Dyxbe26cc
KyySIpsU9Y5n6L/P3jIwEkZiTFbFSUO6lRU2DOAwer+Md2gAilxrT2w9Q/YWwUE9
SMJqRCCXi9oycrshvxBzfYZb/NDbJo+lYeHBdOg3GhawBGrOn3MwU9fHjNzGM+4L
tXe47sFTs0IoFEnBoJncrer0rJCjpI4JBvgfVIvEbHtjmJeumNpw6rwGX0Gdb8d1
4Z+3RkOmBY+0nNluB+GSKAOglRS317Fa35GIEEAJuYwc0CtIkvoLdjquZnjx3ZTf
5d3mg2tmRUolHGOmucqoiplzKsxZ0EGs5oRiC9sDHLeyhKfea/nRseG0e0S+bgI7
3Zu9dpNJSwIDePAg8iL0Xw9qoudVAkNKPmDhyIA+e8ZJdtfzU5XBaNE62ssNNfp9
wWry+/bxVRWne3/D4/GmlxolF+1z57pgUwXxOYQhjbN+nyFirLuI82Mb7V6CTeoC
i5oLEdss0Tr9GbJRc5YNELA6jHWxUSipRNPJnWC/kRhpn+t1Q/e7VG5Ci2bgwlH9
YsPdlx96iV9sKz9AllhI+CO1q5kFFfrfguE58y3kxj+MeOITu+aSDgPLUzDWkRZl
q+SxAFhow9OUUzlJBFFBFPdz3lWucvcVdJLOao4JbfXuKkj3EFpWLPLdN5ONHTz8
5DdcwacXO29Gg/Zn6kFYkU8IdCQ10Dwoa3AwLZ8QjPvIzUlftB+tFSZAspzSkTMU
lswaKVM91F7NJxxPjT4au0CmVcm3kioJYDZsabxcdwpamctqNaudkK2GCh3YAja+
k3xItnjlLpr8kpWdTKmyhbgdt+Ki9r2Uq1edttOGJ+IkE0wHdE8Zk59JbgSuPHLq
Bd4x4jVgsJwzvW9Za521LGQTZFSMRCkMyZA13TwbiwRNS0kvCGW9B5ASriRm2Ete
TIsrSzm2QgDrNayEF6qVBLYCpu/IBqVIpnufa1WxkUD/vcmsH29oybz4fz1y0M7s
OdXSgyrRhZwa+5zmDhKQlWkACdp7BLGe/YSAQek49z7/6eW30gBlQh2ikOd0dT7P
mKTJ3UU+CiKLpB3qT7zOxW+I6jbH9lBgZErQYfzwx86x0lVs9sQtImZMueKMVVkD
vEex08lmKmG6GiILcmCUqSA9H3ezWAupWCsyphxT/vyVmDGC4NPHGNYqwawTFY2w
4hDNTh9ce11hpwWPQGmyehvcg39a14uxkcb9EzV1SSGPGcf+xjbg7DD5EXj8y2Xb
ySOIRmLmkBXj8vDrlYKWClFaxyYn3u4Ss1PhU/h+Hjhx60cjtCFcCEhr2Mv1VF7M
ghf+l+ZIy96Lh8wqIVhp4/G63nHzzNxbH+DocAL63IyuPXPKBqGje8l4IDI+kYBd
e9xU9panrc7ap+O4c6o2sZb7RqxXT4GEECQxwXFN7xd0pGsjNZHcD/iG309DO8T5
DEWP1EbeOQ0JIhHYwIGpm1R4gr4727TslPXxWUCC7XOYKm8BiYDaZDjUyrJ2tNA1
Wt/3w3HRaJSrvfXTngvmE9Eybh/D9Xba2xEBb+cFJCASvZruBE7i4spESPLAoh7M
iptxrTJg7C6Me92LWf3upBn5herq0eHbme8rwx6jXe1xHIfrNq9dTu6x7+ZXt8dH
CimcjM2XEET7YRy22fOgdW7da5Y/s60nIRetiI1zbXdpCKTykEPA4fqK9qYFvoqf
QCkPXPe8kli1QgOjMpr/90vgfkhaKK2AdcJOVQuCbh3HzAg80Wytp7k5kA6ktCRQ
dt2fmQd4zcVBhmoPnKfVGd1T3xxSm9d4ck3ncjjruNPmzXtAp+iyff7wFDHzajHC
ynd/C/S/71qQBJPFZPPgVvvzzCCTKDAV0wvjVw4c5cwcX6dzdFzPlPEmkkV51Nf3
0PTjGhzJecpCiIKEiTmB7DAp8oD844E1TY+BSapfkYDDLvSwauCCIJuyovkwnIk8
KhWS6Js6DGQ19xioiPiVCJAoyhU1hHFpAuFtgs6VoNhjhnQE9vGmxAx0/HNn1Nhq
IVs/P9N0NhvTiK6+cTqaZzDzwinm3uNN05gLM62BfFMpSVyE0sWZ2fxj0RHvC1JM
2ghCqkhzDmkkTYiKzRYgv6JXPe8cYJKrzFsn/bO8Mq1E3OtuzPM1LbxgHx5s886t
KRythhfH2SxobSSkG4LO8VYtS+ep6LJQ+NWvtYa3+atCWjpnR9WeOhOtENcFWEUc
wRXumdvR9uMWxyMiu9+GyCDS1m7vqVeL58xaIrE2w6kfM9VxBO7vu66578lEgB7C
MB/r15cErJV0aqyBVqd7f0M7Jbwf9kDoTZOWO+HUeOtJlgta2zNEv7tXfiULnh+Q
bdP//JFPTJyM+OTVgAbEQFpOpiJi1+HA+10iSujDfDoBDnQNgc1nuXfHtk/+qdcV
E5U+Ax63g9dF70Tt5gizsZTfxix0mhz1hi1qlyoadFynMEhn6D7Cco+pI/GYqBut
9QQ42159kxB2kBNFb84WLw+sDgX4vs7c/2X+PDPQi9WxN/dk4BbuBUx0r5QQ+Ik5
mFVVptkTM53hlBCLKrKx1sgeWCwH9ogctwMGf5P4yfDb0yja4yh8rDsoYu4dZiZz
N7xvQbcdd0/X6HYwASbIPZhqk3srpCMWqS4rpRlbskGJbHgF+KXkWD0nSMda5tX3
119/Dmmm6qsL65rGePBm/5hLQNVu2ryke7xoI6tUGyqqtX0gWV3YviljQh1OYuoY
EnSCvYOb4BUlWaJwOq4x379ye19my4eyxMquDPdGtGXN9+W/ZSdd+ZDmvYk4q0jB
aBuK+wiqFEhfIYRtMmakOYXxFaTv5/exgIoxnbkfFiDlEkCXgIzJIHXtXNKDhoiJ
7/Bw9hdCd5EJ9GdQztrTsKUZsaXLdbQ/52GYmIpCAFIKPByecshx48vcdnCsDjiC
Fk5BllSHXGVzwyt1ijT6ZgRtJPiBD1RzQD2acfsvhGb4R8JcxsKsFP+mKJWExL/A
o47wiwkAsPDtKmjQB7fbFb4weut5/iHVCkVssDawVoi4ghon9DHDvTioVHy6AvXB
/H91BoTVVBaUQ0bwA7EpZY5Eujq0WimGWJBzZtEsDsVZNF1cTMkBDQd9jfX8CjHJ
FvswHxcxbMbJs9K4iBX9FnIc6NKo5XIf39Z4vbwhxwe4hH5L7lFWoCSLaSggwL/U
8l/oFp1F5LNn/OJW+wYOpJ2+zOPLtdSXCOX421ElDbSfAL7zXBc5RqS/WuHygWNh
p+crLMtgYgC3wvykButglbjrpx43Nf9jhFxyHQTO9KKOI30MYjCsK8cu2maDsuiD
a2HIZYAwLDGUOfnpnNlMx1sOo7SB7dbLNWt7qs4Wqc1fdERylLjpDtodDPncfptQ
J8X281/3nGPBpwoEdBlKaKkGLauWfwuhX1G+s6Q+Mfze8nunySGxbiUJ8LJxEhlq
eKbyo3jaDPIKg6aADW/rdxBrdDdLixGZYfoZ5Yipt6RcfdYFDZtIoi6uHUI2LSwB
kvuolOUjfIGKCO7srABdaibe5low4p/MqP7Oyae5cckRSkAR31cZxAxCwZP4zY9O
jTesIb+i2Hi1wedGkRWHtLDitt+FhgszLSRmwKgOWEVnjcG5x1Y3ipMUzvQ4e8Fp
OmB8glTDxa807Mv5hL1zCO+P8veHeWtlrkpYNvwslrTO8MJOUQ67+F+h+voa/A3i
9155P1ygmHzrUBoGMWF/9CabDKfamWk+BggAGkq9C4SyND29Olg78q6tgAO7zO/4
heChtkpzbIOwPnUNvuTq1weaVBoMGFl+wtlPIyqlh8KKYG66LY09EiF3uVpWUBE4
zfeELWHjr94yN/NVwH2kRqLX43LueqounlDYw0ek7cWylVn0RvZm8fUpbhd+GY+g
GgOwrC+/Y42LtjhezCM3p5mZ5GUw5iv191+TibwQqNdMEsblZxnbGHB5W4nS1a6U
xUtK2N5LVta5XaSmxF/pxo9apIdWJJaja/kyBAeOm83EjH/fm44uZKpjaL/pWwX5
6DS/7G8HL6mqZWdxjOwhmjk+ysA/lyVWLyVF4cwoJ/eGd6iGhv16C3JiEK1N9Hqs
G+vcMuCkLqJ1ctuoxaAGzMXIrsxRv+bghyLNGTxiIrQk94oAr95X0GPkIciTmHBX
+sXuQPR9Oi3FC0+P/qMTCFblcVSQZZJ7JRfyfqs3zhPsGSLnwSLB8DRktwF1YFCl
+V8kzoOqo02V4KpVOXkVwVYfr4Z+r4ayQKBUoLb3S/qw7NuMfFIfHoDRN4nsvLPi
9StH8TzVrXS7536jAnwTlXesl+OM1HQhfSp0AOXz5wFhEIY0iod9TejXJyp4qFDi
w4PmyE0mr7A+brkDNglIWfrp0esQIcbJ/+3yY86c86Uxb1C84lNNSoRnsQZf89PO
UzQsJp3gBIVxO6vjCqRUlck+Il6GsqgL611fNbdkDp9mMZKvvOi9u5YtFApGorce
d+t9Zwr+Nr9/LklsicPJWbAcB3LaLmXj0H5AzRrfxiA0M0ygsHzFQukPkvXDUtCW
+HQFLh9681EYM8wjFs3TnV4H8O6O5JmRo9XSrCPU7OWveRC4SHoBy9Q3xWRxSShv
H0vke9hidjDDD99atMIOrWWmFzviGzykD1yKigqsHFKrGGWVheO6uBWygM0LX6m7
ynjkOGR56oBbBHBS2tCqfhlRBgvPrvlkppmG3+BF17PlHSLPEvH4KmXYYCVL3h61
qAaxBTGXAEkjSvWwi4EYK9G9n3fmh9YqB2EHF/wFnbPbI+uYcPA68kC63kCqwT/A
+UUKsyfuehANdLQbjwmXtDHRjvrILGGbcq4fdUqAX5X6vRRSSlGjeYeOsUH2YCtg
5xEl+cng3U5WiAyscxXU8IHRjHCD2YfaUKv5QuDBPea8gQOBodqfPy3kBAJX+bOP
yYZhpWTRIZhln8lgoL2VzBovH+ynhaQQIFANW+oK2xAJjO1nb14Oww0mwtkWMWO1
Uxfp2LKSK6DFTo1xe5FHAcRnnI8fjw5Nq3PxjeOr9CTFmbJt0M/Lw0yahs+aPsIP
XsQKQJm4vqTaQ0uhzrZGD9uqxvGJcBRXZv3DoEUlXHDIjF+OVqm0gvowf4XCM+fY
bd+c8Cay4ijBntdh3aX8uIxKlfwycgPPSOwRvYccCrf5tv3bseHlKmhrsVu3c7iV
E2blIsCgJMWygmnYRieCs1buWkjDHAOhnmr8TixjYaaQDq0WNlrGnktyEZ1tmb0b
YDhjBkAI43y7GG66DGRaGy8qOnQFmArKqWHOU/0ACZE9CE0eHvWeycGsI42SFMh3
OC4AiPWO+XzVTJZNtp1NgMjzfh/3YpygROVogLSrKATcHrzqyjO8lLCtSroW3l6m
8zfPSC9wIem6VKx+o2zD9tMF982TwFPJK3d0IXXPUwHo0ex07sdmBHz+bXOVJXWS
ZqyIo2OnwA01pH9SNOYSPK0wNUqglwvsk9wWq6Kf9qopzi+N8Rg6vzZPyknLEod0
GaSH+79dh71Lx/GBpGUk1QidT+bldQbdEQeg6TLUKeEhpNqWJq5aLllzyBt4TVp3
PEpyZwJieXuPeXehnGd5U9Vk73gBktB/G8LYLKDWEbBQ7R6RFmy5kxPM/Mv1eFJ1
evynTVgutvAvwyyxHLGlnrAq/B58XlR7SrdVoFNTV/SQ1/KZYhT42nXv5AqWDORH
SM99d9ayccwP/EmpKZc0QZZL/qGmQQmhnkYXfg3ysw+lkCg2tjSgCPqfXQ/hcS+R
nbipMRlTwKUuxuPR55bd23XDtpNv12TxnpqtAgzzCfmGaBV3W/v4RMAb6uzQ2dec
KUR6nsjEz4aDzL50LnEqk7On+AmgIyBymeb8fbBrPBQHShGhi6umh/xGYmZlQVk0
pDL4leWV/bF6AT1N5PXl15Jg2WG9Xha1lvnXfjFcMtl9uz+0JOT0Un65WKS0bCSu
tXkamTO9m5WiPA3HAG0ITXJnlUDClEUvCYECOsvOK6brk1zS2ZbzYqyIjJXR/Vn5
fdvB7ubtSICWn36kvbD7UclQqFQOKvLkmXTf1IwiepTuNDGh42ki0+s7hRJ+4TZ5
pxLaYBjW8XyPhtB1aYoD2f1n2VKV9jzazavdVrka8jTH8bobavt+CdrV38vDyPvz
f+aLuq3V/ifhRVA/efgQeW7h+oXkfN9kS2K8FtfgQQ6tZBTISmOy8L2r4roiZdUB
J0BlgQoQf8zVNe4nsnffBoWlMyMGAhQp2NVNy++wH+w2Kx7P8HkPoePPsevOJJka
H/R6EyfrH3nDCIh8tELNuwluRQ90DH4NwHyL/l/FKwelVMz3AvaiuQm+XI1PNJ8Z
onWiBTaYF83+QpO3Bl2TwKqJCBI3UblKqe8x0w9lQF/2Fze4peAqVBftnW7q+ZLD
OKXMZ2JVpJmeBh4IiG6LwNKrkfw9WRTCcxnPDSt+OrCMTquESuoPFfkxSxRk1Dru
FMY6yGpN3nfzpjuPzO2Zi97cc3/8ooUtvLz0uelddW3/puwE1M+up1WlXr/SVvhp
F581Fi5+Wu4MOIPf4XJw2JUjgJqkCFTGKfj1vobBSc3dqqSK2sSU8onDPyxahsdu
7Dw38W7P2BzYwHVcuKk7y1sJokoBrvF38Re6I8a3ZHDPXERuQDIyFSWhJnvQPbqY
ULoypNW1e4ZiEbOaNVtkGSL4YMTJMrEiGr8W9Wkq8Ff5c/wezbupX2egZU37x259
LIbTEP93GI68vWT0M49xwJp0OUGnMpZ5YQh9gU1m22XXd2ZQLTLeGenpLylh40mK
edDRDvaFggrmRT2L10QXjMddtvOIr/Z8jDpIAu0R++yZtfz1hD1F2x406KbgycSd
GtCH8LGlXM6w0x/FxRIOGEJoSr4vRz1xPQzIEv3dwlrZD37Suqty8Ztlpyir2Sbt
zdxU3Facuv9vvoKoMtVm+2MYxF6zUH3keMbECcABD0r3pSBxqZowjxWtZWXa1he7
jQTh1H12k0+41l1IUbiOygZU3SYEkjx4hf2jrhpN2ImNM1BdekqtTAyZQWAOUJH+
uRbITTBXJzSo/OTKf1/YZc8z9k6fZ9oC3Y3YY4JHITRv7gjzu6SIPKnRmD/mabr8
xTChPrW0rpOeQjE49Ibe6P3Daq+t+QKtfcCwuQkhO+oAeNv+L71kKoKJitgUEtu8
YGWqdJ518LFi5LvSrJt2QpX48AAwXHqpVsp1n4COc1ezuWP6GMQHHptlrtxdCWJa
b8btkVK5bIBJAMx4WcROt+YeWAvFhrQbiuAHi6Oyh/g6NUsXhrfkRxax9x3eq+9C
tDqr5yNurzL7XELxKXCAG642O7fcrL4b0cfadF1cF0St4usP2QBSvGbpDPpYZ45l
4Kk35HRj6Henrg/KdwCohV4jkcIRb+aEACD8mPaDsHr/vKJn2zeQSwcbBXk9S7AJ
4UJCY/fUHGemVGPHK9vA57IpFLe7812YyzGEUhjiUCxlUeJcoz5vvkhwEK5yjsgu
dIoe/8FG6BPBdx8bxdouSQagKNn7IPqcf1zP4SZuSym2lWCRwftb0kXeggdpyQm7
61DLRN3tDtj1GlOueuCYw/RHI2j5z4vjZS2A3oNk2BRe+1qWICRVMls3QB1+9Het
Q8AhyLAmjU2T960neCc+dXMRdVpCF4zAIQnImKMykFuYhDv0lz9t16hzo4QcPxiM
FPGAFfW7DxIs8wCteQVkkEN7StyJGEPm/Q7idmmZ5knondIj3RRU6w+iLr4jeNi6
WwNNfnXEdPgmRC3RsAYBoPhisE3sRXj8eFtLSSUqDm682jt7Y6wgeKc4BsMrzpdr
Grb3ZwB8GX/e6H6FsdyHe/hzyiLdSnk3uyZFXxIogipB9yftlZB9bm2tbjx2EwG+
lgDQ4CHuPaL1p9sU97lM/Y2KqiVU/SZDOZwib34YaIa+4agSnyYtNHR78nl/YAvy
vf0oJoL2IabsVWNVbBR2dXxcDddBOXBeT4vykAHZ+QJNUQRy8cFv8aL0A62i/vZN
tJzs5+iJMGoLfqDORQCPypBLVYK8K1Uu0QUxqDlx99wH02Lk+5UKBSGNlZVhKLMF
AMMpQXCs2RWh3LzxXlmFOSh7oBadccFpJwnqZUVC+7ZEXsC2gsdEpPYCveiaEtHM
e9l7F5n/OlJNrfu4Nhp8ycPAHfzU+xDTBC0QHzLMF3lzAFGOrgZPfgvn3NjA9Wju
8wbUHXemkz885H6RsLAsqnbR8WqgWWKKprJ6lkrAlMn8vdBm7/ymst0cVGy+oii9
BuuEKQ2CkmVkNJUCAVoWkyp4fd4u66nHPC+St50EWf7IzjsCcBpfYgrXUKx/f+uu
DkQMu9qK4NLHlYFBlMbJ7w8WenPO7JKQ9EUTb3qPm64kyGUa7j8VciUz073R7u54
UVvDV3ClpCFk9ouLZt93z/rdnDzKxyoJBI6Kcohl2P5TroejOwzSyOd7nzNZFgEB
YRkeLFZCRHw7V1nrcMOwqMvJ7sMRmjftFiXQxcLCx15TAYnRP+eePtcN6HLodZ80
dI4cHvbGqEipfiUM6wWjqz/O/uWd6k8fbmSa+InDkZsC2+HQqOUqfAlQwlGtWo6i
VAoxM5qYtRTVxGE4bf6rSqxbXsfSxbi8AaWSCWZLvCxQFkwk8e5fIUalUABwGro/
C6+33zqbbYVga+EQT4JbfGMbPyVNHXrmClHDBwKlYqvumTCoVPQtup6lQtjJqmOW
Jxvrqu6hrNE9wxDS+s6DV7Oy2E/nXE4CqSIBTD1/b1mRGDKViK3mlP/E8Ss52Qj3
cCvrr4oHVtvoHfLF0uJ0xXiyCch62IJaEQgJ2tGh4ktV71fXljnenF0AzoW6oeZK
IuJGmHDlBMwmCL8xWiq7PXK/e0w5RnWYY3C3tBwNXzl24IH0kA/xwNhr1FfGDAT/
qPkS7AUvhM+nSoHx5eF+/CtQEXa9aqnDkH/b9EIj6wVJHQ2eerM2n/I/tCj2t9wp
KXMdvfvR3o9ck1BN7r5BcxcwFAf7Fn5PUuGK4VlypaSJ83fbhWLcPWVza0CC2Ykc
cDyLoB/JM8wplfeumgSty1PnH83d8nk/E0U5aWzO2IBcWdT6iDDfTm7PctFO/K5y
/BnutHLVZZE4dj81N7HhdygktHXnfniO3X3N+3ZtJgEi0WWgGBBmN7s/7Tc0lSXH
lYY/8MSOhFa5FgigkWs0c8JyMh5W7SoJTOezEnluM5pmqGBRIaeBV9F8nXKy0jnv
3xjyhPhz0d3koI1TS0byLh0sVVB/ehg2+rTENtUMRV8Hv6/5gOSMTvN9yZtBIZDU
PoYdWLqWsJxErP3oQiAeijBIdEKfPfPnTWN7HnRV66UUCCX0OQkYCmakTEi+pKcJ
SDL6ByokR73sucBWLBfGF8HDrwDy1Naui78ZqdoBnIA8Svrxn0QMhPgGJro/P1Da
xilbWyXlyXQU+jjNbszNcXqbEQ7sGJIp//fnv7n46lGZRWAv+17ys1sdyw5MUZNU
X54my/9S/LYp3Xffb8LZVxQYJdQXvqggtHIgDej2hMu23O4rGayhC8jJupR52fwq
ACyxYJT/r6IYxbEF58/PitFDwMKQEv1D5eBk0uE+2ScCUMgcrT8nQahfwVe3n3YJ
ZxV0b1RBWg9/qRAv2ApcOvqC1B4DXV8nGsIjSHBbRZx2iVl9tl8V4NPLfyOxzP7G
vFsmuvzYeRmFvNItnwn/cj6e6YnTvA0QvSgv2YSIpyzaBAQ6HDwviIBXiF2r0Rdt
titswsZkE0r0c2nuMqG4DF1i+5Wwci8FTwVb5svrcS9ID5hJBIKCCg7ORWLDAeTf
pm1HtSdmCf24GmwfISnJevq8oCs8DVHQGJ4sRgKseKdzAVLd9GF/SXw95RgwjxZJ
lqW0hysKYOO0LIM/3r7lI3A5fE9bBdXhUaGSc6XPbFyGWsG9gK/ZMyY6StpGfK7u
fp6QE/EVdsZSdT+d3wD3hRxtCETbq6Or9ooxm8Wp5Vi9lMTOMzQp2lNAZyOHHozS
gVEopziclfbWVCHnGlBmp5w96OW+qMuAYv7JSbS2gg6LlZrdzg9PHlZ435+nEM3Y
Cd8szX1z9HCDCBiqyFcEMIuyY8aRVdLA2yAd4SsRo3xzAzUJUqDw8QaikUMmacxJ
2RNMEVgfX/SlsJyOk6PS//NtQsIGnZNC9xMVnGOdx4XscbLkN3Juprh+0IM1Doko
d1fLuObttf31QxaIRCGOLFy0gMYBQ9WlVH+Tlp/b9ykP2sG27l5/BdZ7qP/QMyTu
ghywB54jfGQF8UtUb/Kt5svNzixXQRv05p126DwCakobcSFYsObUTwhjHYyqmvU0
AfG1blS14C7PUfkjGopIVG+opJHONVBGBdVwdVcX/NQo3Y9eiwnAb8SUAY62IziX
jg8SQN7+Am5/B6Tqw94NRALHzc/rXaB6Wky7UtzSIlJD3Sd0SBMF/xsplyYTO+MU
BRPn39BMNbfg4iaLvA/RtabrZK/sWYzo9M4QE7wRd2t+gygpYqJEg++LXve7w3me
ufaH9tPUqDQDZUUsxS13Max8pTnzemEI0+LumowwQOEjqvqEUHu8EyTowSHpgYYY
CRCI7Rq8zfpdDpyTSqMpkkZQdhz92bzcv99DqesrTWruzkWhew7mGt4b+cDue3Z2
kyBtQ9OMj7y1MozzbdJR2UwRi5HySrigJQK47DjRQWOgtu2SXmWrMZrGjSZxqaGk
ROCiPq0j4m8yqg1t5RZGoPqewSDCvEPzTrbfNhtIeZaWBvnAgej3pXCdK+q3ggdJ
BB/Knfox1YkqAjghABKM++uYFoxO/8SbqH3a8KWFa/3PTnjcvrB9oV/vBE0RbFwy
8/UVL/ogxzM+M+GwX68o9bJr7SyHiTTU7q7JjG99+fmYBPsy082BBOIBT8ajk37e
Yg6M16sAiMoixH80kP2DCpp8fmT8Iyi+37WQbUBNPn5EXaVmnTpvWmUynXnKmmNU
E23bpx82V4AhY1l2DUTG5CdXGWXuQTqWgl9DDA1pTX781mkYo/+Fhn5nGwg23SbP
doQckYBL5YVkqFBH2uzJrOQi+ZQW7dl3qM+rmWKvHf6NtyMofUApNg+OY2sAcvrc
DwCey7a+RY3+99XRuqOtxbF8uncFTbYlDRQFw3NAzYwftYgg0Blfauf5HRxr3Opw
u+owadxCUG/mXYatg7xOdUsAPKTdxYhnM7+ia2MnwzeYN7NOsHtWXOMQrHFsqoko
sDz+kgqtt7hcZTNYUQwjBi1apucNmwvpvfGeAiSWgpW9L84RqjUKricZduQrjs+n
1JW1rVDKsWOZPrwLEBBmtIrxCfogcemQsR0LKi6htdRE2amrav7HwFyElK0HQJan
ryhgfyyRz37T3TzlagIO/RAON/QCPHhPbjgkMWf2q++vwtH8LbX1oMKS/84AJYAO
eLGFa8AD2QhqQuOY/aWiUZnq1GasRb6jdybTyxJu5XgAx3W421N3nW/4c0LG7G6V
dSAkFrSIXybOIRwB+d1bX7Ujw75phQ5sB1T6fZgMzLksIbb+eBXgZZqA/RJHhBlk
P80PAf6OcEyOmu/RQ0dkXo15Zz4kiGUipxaM7PrpIrzQz/34ImjU+ZzKS9OEuvjN
fx/Wqfl1t7a7N/k+v3FXCqKm0BeNX4B4q99Nh//dz+D6K9aCHF1QVCZ08KZQZNcG
x3hc4XIoStnPxfxWHpb10Jq6p1mojtP1Q/XSWXtVvTCOBU+VReScgENHUJMkxNBJ
3UFpPx7H+7/kYSQxthNTkxcKIQnvQJgXO2Irn2vmIknlSDSLHheAFm/DbSlxD9vI
vdwFKIm4CnoosAwl6Edp63Kzm2VSMsQlWpYYf83WBJMRVRR2fV8aeB/t/qqzXokN
86JJSbdJ/hubhB7ppL8cHlJuVCnXkyfmyf57RNHSDAnlXIRJhdSUE9mu+MiF1q0+
98wIEV3uxnMaiA5Wcqtf2lXa2f0ty3zqbAOkhqiKeafeTRAMSe7iB4wOXakqR4hg
vz8csmxIDet+9ix6PrtcV/Smi/AxA9fYo55Fje1kBqg0CvyYIkJm7vhozB+feR5T
d/a8qA79aDS0KJiwE3US4+65R5UmFZNyQDrMymGNbeb9B1LKy4QVxAIKCaScw30+
8I/xuoVr7XQl9FClmRRZ/Tz2m6cIHb1rXTY04Cq1T2poQuGTi4FQYn+l/psXOaXN
o0ufg4UNd86LdeUIJXwtLI9xhWqeCpLeQMpVuREGxP36a6gizyYTn6N7wHPkn7WI
vsJSE42Ao9bWCgxMOhRY1BMemqAIwvlbUDZ54XRm87733kobBQNO5VdnM6XWJlSe
eD7DeGJErbSFCvNGHVOvQU/edzhOk9zf4YtSFddQJEfjHN+garb+Px0A0WH6rpYA
+/fPYr1kD+Y/zxkRjg4NSWXQ/on/sFbiNi3EZwTjMqHKy522yX3z3nfAAmRWaH/e
1xsX0dpwDX9O0Z+vYesKEZhpqjkbaxQyefNjjtjLdMl8k6kM8eqB7wVMp2LptxPE
kpdScErrTktNpivF666n4EX2ighgC+h82FwzXW1KDm64HvzaQPXgwzA5AUry3dik
JrhbSDz2ZPOmG3vWBkdlj/4QHsarb+U6l87Kt6XYD6i7oEzeeEkkSbIEkQE67fdV
J25NIYH1JoO7OSr4rShk9xzzRGeKxRkQino9KgiMsjTpTsrGG7rQTXl1YkLWtQtx
vh0Xao0hHfiYG7bY09MyqWBVMPKX8ruSK5PVUXoANIEGOe5l/vT1Y3HJ4li8kT8o
qsG45KVckBut4ZvRutnt0R6Z+syxF0rTYRoZgQar1sEx6HfyoVrMMEwQbjCeCG88
2NuiAx4bCLiTattSQWhlQKsPcg7cQaczVSWgT+4ENYjCpj2uy9Bkf3WJHRyN7Nu2
VGXH2FXEwaVgS0mcNZvb6rRjQUg7xzrIN5qemJTSuHNgPGveyCT2lgjIORoMAQjo
Fn4pB8MORrxRju2kIB2kQ6rrvME1OsYM9xbaCfLr2bsEw9qBxHi2eAF7tfb9378s
LCmf1/sFjhL4Sm6cy2W22wgndWmabAxa1qnhQJuq/3ZnUfneHZ2l7Kv+zD7CI0u/
sbRr2aI+omv/r9mFKnbub+d9Gwfsh/YbuoHz0I1QMW1KKYpmoDfnZwLl65AOhKly
72Pa9Rwcw773DZnLl9Y6ck/V8P3mmHraRJW/3ayxIngtGpOwNlPzHcd6o7yBjdv3
+EGACLDbP/ojzt9gD6BuJ8GL2IzhoMvJNCZzAmyf4+hZfRriT5zv3Ayc9b4Wl5js
T9LN4FrBKemWmRVWTZwB+2zRUGwmc/1cutVITPS5J47UbgXdyNxcVTX2EJGzS+9T
otC/kxukmBTlaSZqD1EnrMDFT1bwI/fty9TNrGKJb6u7KM0vOrcUi16xFcpmyOPx
OPetngg2yC+WTJILsrEPG+8EpElPTnqt8O2NwupEqUBXEb6f6rvzKhZGicurdiex
lW36xUjfd+N00kYe6qqMx60M4Bve02XK0FuWmWTO6YldSyS0AY3Qw7j4orsll0r+
sGYeM48Wpam4mPoJnXXNFwXzEm63mLWc4nYbeiojh0o6l/izmDwsmAVvV61nwDL4
6PqLWgbpVU/1OGgfU+tyajaZpmi/ez7afSjpkReJXWz8meXHfGcMm1VoTUHHjpsx
PKysb9r6LVTrh1YVaIBF6YWzJRKb4IHMWLMR+Pb/opyBDDWjOGi0txRAa9dp4Zu+
U36HsJ/x5adl/HzAar7qRIK4J0MGTh/CEVIuoA5mkET5wPEt9g+DHwFzePD6YRT4
NABvFnS9nUc0QUrfp6kkDBF0cDj9aUpZU3+x2zAE18UrXsokRvsRBHqNXhiMrfHW
2d2YYyZVZ/jsv0jC1/VsXGL9RxfGLnoEjQhwNJ3I+k7+W1GNmpYT6Ner/E9pufYU
/WS5vLzouPS61V/ex/7Shzz6V77eZkBEMUvEAuA6jQaL8tAz8u55mF+qmTexo0sH
2nLklKPQWa1qx6zvbKxYPkeQZdXTZ0X4CDr0yWx0dcQvWPhJllGsqBB94xISMsYo
BlMGnPw0g0atO+o3MWsWC913H/NvuU0B3fjNXFTwOElEjvYbMj90LFr83zsv/L/U
metKLWUGHkIDO99RVOkVnef7DxRLSSJ1X/koVU9fv36PU2PQiZXevZEX/GkFE1Lb
Y4yyQsutKuPlSQJU+U2g/Rc14BigA9P5ORK0eKlXAXccQELP3bPqnVpgcEpuWtEB
6macMCsIxrD6KLF9+a++9YafCBm6hXCAqleXVC9iYPfS2DKT+DLDb2yNWPSGD22Y
sper3cTCO8RzYJjMvw0t5S+6Fq9708U/GJ9JMWNkiwj0KtUU48xP6mW7Rd2fIV+r
983mOfRkAtrGEhv+s1ZhAhutN/Me5JfhLgnZft2SCAdL3IBcTYJ7CRDTxsD5yg9R
yfTgjLtO2oWTFViktvFYIdvBNM+G7lNCioWxyrm5G0NrJwUON1BHRrKnk7uyUFG3
pjGFPsqeEOOJWt/NQpIb2PCO8csNCTu3rMquO5V0JhF3tnL4E4025jkvSCbf5V/F
1MRYmyfW5BbPSFDse7J5W1+lkFWipFclvsN7TCotxdRqakgtSFxzDIkrU/A5TMQR
n9QeAZFYRq73aYMqDwVgWOOH/NwYi34Mzbk/iQyW5QjFUVFngM0j/mL4s9/ZLRZ9
IFFQa3/+2XTvtVc2zf+VF6ZdAIp6nrNd1+vYLRfmQgSdIY13qmBWfdGqm++Ex6RV
sftoqk6B3N5oyUdubhGPrEzjoNXeYvNqukrRoh7c9wQG+HpwCcTHa5QaM7sX1SYH
Ka9M9PUpD54TIVjD6pRyOza5B0zNZAGUICwNXv8LAiLhMqcH0ME6VSQJvGMyAoE7
vyRolD7Uni7y/mvaBRS6BxMfigyKQ7yEZbC5a0mmn356HY4FcG+79/CS6OBxBy0d
mSid6gMtXH6lJgDrqWTMPCZn0xtt59gVo5kVvt922C0wf23tPSZ6E//CGFBEXM8T
etrOh0Dyx8yMAMb+mIsNcwZpfKoFpvkSRE70dDaEjgoidXX/EuQ3+wjtvVaWS/Wn
+M0Jqt0R7oHx3vTz7wDIJOb/a5Z1mri9DRKHtT4Slp+JFyDq4D0D4ja3MUQJzgSK
GA5I00CxIRnvqH/af7hUqAAqyjQfu9/MaBMcwW9E6G9Fl9SpnuTDd8bVtUhtdqbs
6TQzllGkO793VcFAtHDuyi7kMmmxPstRS0I/3VjcnqqtOnVTb3GMgTL9Ts9XjLEV
iPFhM7HjaIIyY5FH/6Vf5eJdMEtAXVUPEtFAI/O5hIsb7xQ2wO1hJmpSJuKExIEp
QSmevh/a37/WWHVfQKsYxa8sSHBax0kyycwnFmamqagYGPnBORLykJbRYlXjnNZC
WBoeqaD274D7Ba0VNigchJ0BwIgUF84VCanbIo0knNClglUXuhnN5Ng7NKAcAVIJ
0VC6Y1V7+8rLoQuAmoXsN/IOsKhxjX6c2XAFuW8P3kxxHNEtczfkeK3euFbas2zx
qKGYCzJjbmTVDPfrQFL77YKL6fafXoWR2tWv4iL0HTyBTDfPGeO3Dq1etorXTofA
MijL202be6ghydhepLQaZ9pEQHgKlBswXjWC5kjNrkIhIPPHz++LAcPf8MBPUeLM
c8GiZU7wDynnfASaKbUDrPdxJcA/7hyoFGtiiRVdEtBBH1nugqMNYOFgyzlw5Jdd
UjHP24FFC/WUsZSoZb5UmWuFF6JgdTUHkchFGufT6otM8QiYlApf9n2UreK/kqU2
BM4+800935zwES4nzLeop0/0LRJWdz7kcLZ2scWVSOYqPBFv1M9GNa6KGgTJIJ3V
TRiG6wWF0oMbVkoB9mgcOjUJ1niFMryNICwm1bc/fla39zJjNKWZTi8GQXyN0rSn
Ry4uxSrMgKbPTPKV7dAYXeCb03QQ17RI3EJntIHnsuL/D5xafSsbmJhTTDNtU2PB
AjzC0AVpL3dvmw37t3juxsdryGo9FZpeEE9mlSouniMKUj7jVdN9+oukRAG7X43J
0XriVxE3Bj0ItUFrTD9J++3usZE6BbeCLDt/SDI6+Ho8TQSvNbLFAmbOhXLNJ7ev
nZVbCBX//M9n9f4+vr2nTUV/AR0KlO3Ddpo0ck0Dn6WRHn1jRSi2kNQBPDzJW1nY
xNz9z1SEM9wOhUstjyQmKKsBsiHH44MyPW+z1SUornpwEUzFA55z0OdovraA/sQ5
A9I0OwuN/2fZJGJNaaHUgtjM20mIROFyio3Tz5em8n/bmuH7pA/+gnRJaQzFx88A
nvnz0Q5Btiy+/wGGTugKsmOW8xgnDPH9ApMD5eLcbjdvaAb0eOF4QLELa/VDKxIo
+oVQIdyiQlNAnvEojVtfsYJ+HQ8PhX4ZXvymEt8EGxARyrIG2Q17JJBjh8lm9wh4
M4BBis/9Hcvnk215WEFQ4dxLX57/9zLtBTyjVX3XTc/xZbzzEm83IF+VF+oz+ebY
1qLm1gWhS3Z5KBYRAr5GAwFtCjdOPMpH0FS09JHiZNZz6vTxchyz8k/yYXd73am0
W1SFE6+TYiCyDl8uLEXJ94R0/y9GcDbDqvWfWuwzrWqdXapdsOk97a1TY9cTmCRE
iZQTsXmgjhH0QdxLwhNVZ189xF3hlm9PIHCxfp5CoUnHBTrGcoIEWYGP6xe5xxgi
vgGhiCoEdDDfwIrgmoR333vVd2lSQrFT3CZlWibi/YfCpjBrKBzLd2HNwZN8Dy1f
0EI6IEiDWTaEcEtxgfPx7kmOhZIRxgFO9HZ35YTLLrPoYxuGTxAo/IxkxsRnRGHb
fgfPJwj+SQwyGGYHs6r7QXURfVXEFFHnfjCUu0G1huMZ3ngPCRFjqWadJwpALgN8
mitgywz6+WzPrp260HuAThJRRpCOTQ8Iccf5YDzEaZWJEHobEXrO2et8TufJcGTO
fHkg/l42a/Do6ku4g7c7gWe9bQm18REUbFSpoH4gh0KwPlbrh13CeI1HUosv4Rka
iYKjtZnMKOU575mELOl1pOokSDIzj0LKMBbtoLT7GwXRyst0HXol4TllNrLqbX/k
+ZZYLPEsIZxbZm3YHScjk64P5GMnGCx5qjmB8PcWpIZg445qcQPG5eV0WDWYd4tL
Uc6HGudmJxPoCMaIEJdEo6QseNt05BImgK5l7AZyVN4vo9uBGtBzTjdTIdrYxci6
27xcQOKrMR7uztNeWT/L9SnM6gIke0cS9orn7oAoSp+1RZu5lemTnzgA7ybKggCG
Wzx+cXUKpty6CxiQQ48NP90g6qqJN6L8p5kBvlHgrf7ZuI8l+/y7AYYpQE/NrObh
6O4Mst1C15FCqRyLjNc30D5Bwm8dDJLmuObhky58B7+FFBcgkVfZb/RRrROoGaj1
xiu7uLIW+lCZAi3+T+nCNe5G2ZVX6oI7CaogR1bXOrznHozJOHEccIVuvH89fQOU
imqopoahOfU/w8uBl0Ip8WdCMAJeDiM0wKLibgZRrExl3bqRj8eY2N3vFhPC5y/4
Kmkw8PuZSxnxwogKAGvwoVK9+yw8pJyAGCnejrhEAHLKm5jjT11dXPqff9LdjhGE
wNthADkzkBo1kHvZJzaxiEdfwVOJOTby1BLPOeSRQhMZEapkMDkl4xQLJsu/Yezb
PIcowa/tHPGFkMIRLy+zq/umhpHGUfm/IBJx4b1ge9s1R8WozZxEXY+FBuCSJSk6
ZC5T49ikiQPyWzQTTiE6GzcBfTnyB9K6almFN41SMbV2+cyIwUM2IC+zsH21lQGn
a0RkBm8AumCr7GdqNmf2GywT2fr7OUnS04aXvmWzhrbr/2K7+xytHOk4jvOQhNnS
U8hASaRb78uqkbXMM47XcdWK6XPRB7V0HyM0PdNRsa3Pv2Rl7OdTdP3+yVFsx0uI
qSZ6f1U/tdYLJ18hjTv45WjkHpyHjdUov35TknTX88E8SAIJKO6TIc84UYW7OdWz
p7CIVOWoVY1HRRRMT/xF2Eh3ve6s9XHN+KuPvMLLA0VtrGNnwzIVrgNcOzj31YCP
hnCSRESlBRc74pSsFmEwpnZ4uKPcyifG1f0UCHPluJeKQlZscPei0QGoLGwlbP68
6BvJ8gL9rxUGucRY/N7jHhLOgUXQXJH6YgaiR9tvm4JQfuWEdpWtmhQGuSdEE8FR
tD8Svb8sZx/NqZmOcER9bofPNsK/seW3MpjQ6xEzFW4k/upFrxKMj9ZdWng4fsRf
cWptjCwddTC8ccYLOuoAHR0ezCDfVbuff7G7p+k5B47u5fbYwWOvTUQBkrIvemGF
riGq16JDxYLSc1kQNAX0BRYjjf6KKWvWSoAHgLkyHus0EDdGCfbdZK8EmhScwDGa
7Fw7FYCTh2E9l9V+M9yXlGADJr/flM+mB2PycNFhkUUPn7YLB9OoeScyixYIKF7Y
F8H+8wl4KQ17GESPSXSn2UwR5OJK/U72JlAzpWsUQCILhxbVDNLJz4cLb/5xk4kz
P87xbuIE25Wd3MMTDlM/XU62hAjmxjuOUJWvZ2UeQSOMmOm5TtegaKLDNTUMfPbV
Zh6xncwva1RJXRFD13wQcqSMTvXTjfDcLj7fIShW/FHfWdl4BhD24+L8QqLyCKlD
OO6H+lNoAZdd82HFJbrvRtIgyPKD0c5glNvtJgf+KQ4WPTZWU8T7mkI2VmtObvsE
k4obnulrpb1NaWhFrV3QHGvl0M9q/n+4ZwK4MYC1snMkDvpgwzwIupDG8bhX3AhZ
7CqHPNA1ZctmJh2fO/0b5NyjEe+sGTbSm6tgQunoABJnZmVxwzfUSoLx7B9AROvA
1Hafra3M4LwoyPHLXhfJ//67IpIO+sQYKnt8VI4IR8Jn8DRmGnbpMUnaeDLERRF4
RHJfx8DiQUQh5uwH/+wO44B3Xx8QfX4JYwZJynBZANOX5mv9M1tYc4/ZZ9TMAu6G
FbMZO9V9f71POfLvxldwGcYFMKv90DZqJqQ/QcbRHPdztTC+N1zwoQuV0HA1nNZW
B1VwqkcyAcjA6nbxZj62HuB6HO9ar7k1ckLL1q7nvJkpruGP2XSKgiRK9ZSQaFui
Gh1S/Vah/9nhIPuIo2naXBcIkyNem3GVFQyhK1pn9btMi5fvH5zrt62X+hr0H0Wt
VWanVQvZKCynxLizUpzSZrjVTCXxQQvVuJUwn/UurE0BUB2uRdv7xXalRj1ifXYs
EcoaLqgJabWitfQ/qh+arpqz/Ptl7PY3czx23oFNcji2Ioj/O0doyyw8xk/vS8ZX
wWGRv28fn0W+CwzV82Hr4kYvoTS0bwrDrEVZTKYCW6aQBjfFfkyA1Y/IN6uDlUFx
+vhvo2n1ewjdCx9p2Cj5wvFA9gc2BYVCUz0tPMmaHsAQItXfs9h1UOx0La9TyPSI
H27ehVgmhcH3tI5qSyy4b8qepWKfZpu/gm3fEgYELSPHtyGKjERYpySkYYLg2dG5
4Pq1PM3Ch18R6Xak1ZAiqUVKmcJhEiuuDQoe0otTvEjsARA3L5ZMpbXyd53ti59I
Z40HOp2+T8vYodRNyIblLxGRWLelrXdpC9/TUfJ4elyLTfRtB2HjlrbXZE8NfDiw
b0bzvEXX6pz57PslWwSxbNFiMuPO20itdF5GlgR6E6gxw0uSqcgqkFflXYrJeZmA
6r9DJSedPZ+QoA/7soON26nhRaPbzoNqtOAv9516QqMTNihpxZc/oR4BBJh/vyok
6J6b8A7dBX/Sq7ImWDnl8OkaBqnl3WKusSWTgRHU0ezjopWAyDG74t3aGsSdR3Kp
aG0yMs+OOyolry2JourmsK4b2DPe2gu7VisxTSHT7/3/w5W8nUHzt7roPRXGyhqv
Ti0oMJjs0Z4sBvN8lugRbim+a7rwSZ2aJaCntVj5u/dBeiWf0bXSY6sEagec9t6b
bTn/eyZkHmeWt08wlEelRJxZ86qYy0t4UKj4s7BcHeVXv9Agl5PXp9rEN8a71vW0
Gi1q4I4+QBtzoA9DkXbaqhUhzo5a0hMHG0ME4rokzloaLCDABRkiB1A8yJfPgg19
gqpv1tE71NQrS/dzx38dceCOzC4B05XlSRN5GQqNVHxgdmIVLjQWbLmn8Ba63Lza
TAIQVlZfUr9UbqWbUw6M3yUK/Sk/3qbvs+RnnTIEdna2YYyqAeR6mkPdogB9l+Ae
OVPDUHrBu89UtdWRFpo8XfwsVK1Dwq7o4hjV4pahxbU247VlorfnqQLFTQTPumIE
KKXiihl+KljDcWjhMcU2BMIzksYo1Cta/AB10leWACsPD1jzpCJTLrEqr9cN1vIA
Z98vlxKyUiGhy1fy8WLSsNN4Xbgluqn+qo2NqWSlQCSICXjz6VerP2S4z97WHSzP
AcZYeSOf0Yf2+Hn8LyeCzEz67mdvnCIWB6SI8TXhu04yUWIwW2HGY7/QlU68+tSh
CoJCDFc8BMTnjUh4Rzw1B35HHRVbCErKnonE0o4OMYRTIX+aQuMMvkAHj+0JFqkf
FmlIc95oG4ik5IcuVWAAcIzRZ2QYnTV3J0apgw0PlXz4jff0xbrcGxv7BxVOICin
Sn53bOLAYXtsgFkkFLw6xh7dVpAKRB0ckeQu48h1fg13/0dCoKG342lF1k2I51G3
eiexAcq3IHtq9Hhy+nTrr84BvekaNj8SxkQmmJVJtgC+n56kOUCujcPnYksV/Wzj
0KfkZi+7wn0Vgspduc+Sm6ACbkaUpSzO5CStmCwL91RWO9T0lUrXAuxPGQypELrI
2aeewZ+RNBSZxGTd4r35w4h2JMtcomAjiDVHG9/g1Y1WVNMBI6g+LFLpQJTiYCf2
OOkTNgQ4IsQT/7bgvWeL/V5aDMC7BkUp6c8t1VEtbbES7IJeET5EBfEUfC6MnGA2
JIInfrD6XxgH3l/J+7Wg72BsDKksXD+HPFgelMs7d2ymFqYFiF6l5L9fJrsk5EsM
9T2V9/ghUefjQ5lsCkZcNvWgW9WwwnF6+ST1iWBaT1RiAKg6kfzTngujs07uu9lw
4h2V7wxhh+ZEge6GwnfzFJHJoET4Z6LVHWX9a6VSiy3GSHrWj2vKkktTU5D4G0sS
LXByLZDQu33T0izzvsPWpmS/Nev5bQScE7J5xsiFN0OmNpqLuHUn8w+xmSVD+RAA
fNC1Z8JnW3HjJ75jAlraVQz/OVJs/yfFTMjY4m07XAN5NJWzvW3lWdQiBhhwnNud
624iGIbjdycuH/o4GECDbabNGEuptDSwzhisSFYmTOV9vbhWVpJrw3HO1XXqrfHi
jaeZYXdlSn38lNT3h9P2GqsZeKWT+fwv3ylre2CdKzNY/mEiYMY5zdbM4hGsTdrf
8NnplzBQHk0TlxJZ9udD3fXXzYRLiXcIkn0zpffHDRALjGVP3o/EI9McAmP9K4sM
Az06rZKzl7KRg8weTwPWPWWx6FIUDZR+70xa5sOsYkMqZ33r9GJz86nteXONQ+eS
FdK/7bYb5oW/NXSy1FrwwXdgaqs8sqL1vskxO3cRdeiPDrczuvOw+2mz3I49jJhH
vQO8JxQTOAT2E/TRvVni9Y9QJoWKuPlrx/eoaIDRM9tHq9HQ/vSJY+sW3b+kuVbh
Rn2n1qsSTWKyOvLlu7jCKZ8rDtgfzKDte9O8RnDrCTugo/AxvZGCmrzlMZICc7n7
MM8k+0OMz49W51ZteGDcLbx0h1yRzaAJzbNsXE9ujiPaNASeOp68/qKu387Lsr7Z
DZe69eRuvUlfZwGJ9hpc1njfYqVMPQT9FMCRQiXvYkqW/rFOYHgcLjV3WrWSqKKQ
J0R20xzu/wauXa+4j2ibQwi41HJnRGbejokQ8oLdt1bkXyHIgIuN1y3Cq/LUDx1W
nScn+MtcPBzvsz6hIUmu2j5CwtDJ8TUPdXKsodYiENjNOO+C8SjtHGFFTwU3pSgL
N6o0/DvX0+tklM5GEeHsggGEHfj+v3PO1K2ZOMwK9Z76Up9dcIOX2X2ysi5FLBTK
/Kcx8V8kQm9Rlcrvj11/1gn9kvuUshgUkPw7zU7XG56QS/mp67NkbnnvAMlihXn3
KvjphT08dIc3rT5pNcFnAAammegLEyzcPpTGByhVN3h9nfQWS6pCAZ+hU1m7kGu/
P0m3yawoEXY9Ua4dQP9WGsIedc0fZ3j3tpYtyTU6GupCP/kMAhg0uiWYHDfVz/9C
p0BiixoruZif1k6bKmCivg5vHa7S4ESHO4ONnFhzpi8B0jvDNNrxlNJ6L7Io+TLe
+gKkPXIei7ec2vgw8oI+k+oMW2ZEGhyHn9nTzxiRiOj8JbzKCM9Z/v1jIYfGILSx
DaRWgp7j7bSM/3POxKEbTFFmgiD9GPYEi6SCRP6WijyPV9fd+Uvocb0j1PDj08pg
SJNiFYzMazRW0HYs65STkiMAqIdFdmyq5QrGwS0V/adX5h9HQ0ZKFF18L9ol9Ubz
XNHjIT38Ojk3Ihhgekkq8DjAmz8e0NLjgd5DPsH9027t8CUcDQI5lHMhooHxVgcM
sGXZH/ejwnYkghHtKimoSjy452PCAwlKlQlPJPDz9O53n9xBuuj4F/L982LvIgw2
GhqJXUDslWtDzMbNi/GDgwjguxL/yzlohnGxpZpydfVSEN+17IrO7g4w+IiiKItW
47awDxntGEfFardsYcP4pSmyKH2Uoe5Ci2IkSCyzZMATOsjS7MUDs+PBeuhWt8zv
M5Dpw5xyiEOOUv7cNLzeOF09Me+Q7dkh8KokZiFlHg8hIDWlkfYUaM9QQ3hqsC6d
kcR4/act6FEV2TR++110TBz8kjjCzYdI4/JRxBMDQSTdq0ZVdDZo8ux8MGmNFNfC
RmDDk2yziW0vzCP4PP5VMHNcDOVCK4+qA1IRtLCKU1dqrael3Tek74H2xd2+lb5E
MBJ0Eq1JFJxmeHeyxG2GTRnCJntd4waKJHntZrSfYrnv2i4OztW8SajCGISJI+Qe
N9GjKVOweKZhOndBckKRLUQ+a3+1QyMCRDxoddqpmSCnAvV0wDPA85efmsjZYvZ6
KXixlMlfDZloPyzfUUd86GPB3bheznv8Cf5pidiCmCOpRMTPHWbjL0YCmfRh4gDj
PKmrdggEmt5zvMliE52bHo+vSgf6qSPmhJ7J2wgTwrUzkwlj64Tz5uZceEPZpth4
sGmsnEcw0X+svUUWeSHsoH2XjB3cym+LYNZkUJ1Pem67Jr6+67VS21WKuZF53Wix
KVm7nw8OEb9DU6cS7VgxcqYG98HRKHwi1kX/yeZJkMdLOCnGH12ayAHU2jbgN2hy
f0RN2M2nSlWRB+pXafhIoMUcpBkN9wjBA3c5eKwpUnYuG+Yc1PS3H4V/yyVqTfsh
NDyN+w+jnrCH16R22VsaHH9iJB842VmXcpV0Fzjjm5FW6dtEOHxVLfoz8tg/7pXg
8Xs1GftyOD+VZxYZr/tkiUFh9XIUf+ph1cmy58tNoxI0TxvOSnZhwr0yCa75G0ut
qCSbf2HeM/UJDZCRoqZAZvDK0aQ2lfPCZi2zK5tju09DRNMAuKw3yAA4L56H1ifD
l0bV9E69wuN7YyUBmL6DkXCns3etVx8umfcibid0UNJNO8R7W+uL1XS8aDGAFx5p
brp5bjd/54XrUcUefzC90RB5C+HcfPIEG4QDfY0OyWND025PzdrVjMd3MfZmAvxZ
dJl6cXYBrJ33WVBfczjaG2/3rRiyux1zTZAWnhmcv0bUMC8KGntpkFKpG/FfkJ3N
zGg0BUduA8MYBWtfYPYP1uhUy7sUMm5auqdJYtWdDRi/qKcSu+X/8sbByH7GeYI9
o/6VAW5xiLbFBQgm4L+cx2OHlmOP177vSZ8dgYUjqGO6YtRoltIKezCZIoQLSv2A
gKxmgV7ZpGF5C/z43XA/3RKtrrBty/9Lu7ipyMAULu8/aV6WHKCZrvXIL0V5zB0c
WCsIr9YCJv8+LcXFvH9NGSU1c2p3QFKGEpwfx4gM/FLbawMtJGzRex4IbfA921mh
dsWgmF5gwozauFtXQrjxRtztW3NQvRZUjldWZ9HtG4MohVIpgnimuCNkvmZQ2NSf
OHpdzDXY+5RxMSH0tcgy+Bigskr0bTa03Zfr7eH0+23tyWmrS+Yg7HnPAKyJtmw1
Bb2DgBB6Ahr+I35n8glnVkvJrmCmwg+TC61rJgdNiQkHAo9L9KTsqa9Gv/gf4u+q
KJABjBbvuNn2AZjWpQ5jQu0Xc7SBZdo+XSYlWCBYWXk6BK/FENfH/selO4tJtRUu
fdqi+O1fDb2gVzhD1gzvYgm9ZoUBw2dbDiQ8xgZURsvSbYAJME1T2O0OBASKdw0h
OJZlScwJqAmAqoEgc+g0qnru4tF864ysqQt2Xnq8vIug5yRFvKGqNfPeUln+sH3V
jSH2P+9ypvBKT/++gQhNmbt60y3thvzDhdCb2/WP+s8JJhQcPZCKyQg54UfnnCcs
VgrP4309fJ1orv4z8J/L+p6SuwI7d79U+2mqpoNdeBCdMXjawfvjllPkp1jG5IZf
gau6pdokifTYaYGyXHAO6qKTO0meNMzTYwfFHHmUNkaA56RtRuUCqo1p9K1ecnhv
khJ8NJ0X1G3G+WAqsYwEVNqpt7T4JU+exndzPaJMO2Kg2vk8UskznCM8gRu6lU+x
VUyM3kiU9om5ntm1PXNHz5FhkAqeUhULBNyVLZONkDQXBz8AWSj94CASfCfRgX/L
O5qA5lkQJ5GEZezkeLgT6lvyGZfJo5HzTizGvnHg+F/PJ+Ss1aSUVZStb3zvKBnS
L5wTarI2yyQntppQGzuCl7nBdw0Kdn47k3OJQFlIVEvhoAnUiB/6AUQ2zFd/zOH+
28jWYYKg+9CL8NbHdYsl+TRhutM2FhRb7SLvmaYP2BEevdHqcz/QB5OUs16aruHA
+2KWRepWb9rMtydkI6Y8JE92MCtkdlWlAiFaNXon7Q3GlwGGfKDPYiZeupFEEH3r
068IpO0GGdIpxsyqIKlZCk1pwJT54WU6pDSott66BlgHeEu9aytbc49P8GJE30N6
4eTjawNxr2xEbQsiOrddc9FtlbKV2xw+qtoYS50/eF6PLk7gG3DWUTxJU2n5YpN6
r/Q90R9NYl3e/sd0O5dWGlnW2FkxZPcZoDC4XCoNYjI8T3dWYVPZSQKG1c9aEW9q
nL3lGIS2guxevQR+voP/BLy/Zw6K3oB+8UQaF8POmRCA7Jq6nL9m4rBiKb78pzzv
7skQRnA1UunNGrhu7Ll0JL/t5aoyLOBg/AMmvvX3xKvlHUDz4W431hdBQAZSLgx2
6VUTpQIbihwHqV8Ex7opXjknJ+JohOWGUjdSCDjXjnF4gXkduwG0feubr76Z0nvb
fXRrIX6v+gbGjtc4HF/MzXv4ZqHwll/XSdCfdKXalfvwQXbAq3kA+S+NRenP0kW3
bYGCXrZhXMRNuhmbyD+cufaVjjViJ6jzWbrA4xBHo/JlFpolC4VLNeQ4Vhrp/LRS
ZNLJxY8P0SUdohrvjBp1ZixQu3jgGgnInI3RGxU2cB4jpmCWvX+u5l6PklUMCg69
M3yErm1coHoRyB8IwYKWDN+NWbQhHpzRugUmK7/9+JAinBer7oS/+IxHNW0b/8J0
+KXBn+zL/x2ihB6GTD+PxOZHajuxzr7p9mucdh9C5ZGEGUIy7YiCZO4Z5AYe2Sui
LfTygXd4A8F+1VZw2gn+OHb+skkXUx5M6sVvEWn5oCijuqLOvI0K6xx361Enku5n
t7keYRFAfYo1JdPqv5NL54W5CofqBwevWtk+9+VVLUCWydYz4dd/8cisgdoPW2UL
KvrI6H8DpZS1E/TQDvvgv6wZdP00jRIm6GiBxCBUkYZeTXVTpBOg3LVOjcZh3lkR
y1SiLV5KFYYM50kY1IPSEvr616oME/I0i0nfNQh9U5kFk/WTmfeZwUW/b2zfzhAo
1cIahotxkwujg64a9r0xQ6rlYSy4gCkVFGH4CzO5inNZk059ZCDKfFl3UiIMBfdw
DGJfVCRJR1OHKVuyVXHGYowYhBMbNxT/ZaeGsiWqVdZYVyNsWhppQ+bo6dKDFb85
ybWxzl9IQ23chEpMd+Qk77EulHlXqyIhTV+U4SIR9otlFq6BKbJKZhPucaS7q5d/
A7RkabC8crR/yBwoo82ycou5Q/kJnZyrVfW2QCHEo7nHLQ5Ci8gd8TAD/yOwic23
18MNeqQFt0GZ/rt4ZV7hSbeSapqL/pZhC9dxgFvyJ+5ZsjFj2r88OSSN5rEwpfIW
XQelRRbMZ5OyhRsoHBqbdWAHpG4/cnyle+lbLZhrunWMzZR8bafpM85eeTmxPUsd
BFyxBjdWcJNqs/IcMn4mFbtcr2jvxrXA8A82x1fVGwm+1Y11l+9Rfh9+5TCHENaP
eqQT1mE3l6Qr4wc3Z3xlToiFkG3Hi15uucIONWDrQqzfEzGZpPtlWzZrr3yO9Idu
3M8Hzv3HiQoaGlNS6i9achv4GdcGsnDfVsgalePRHEeGu3ACQ0FW2lT6XHm8QERx
P9HZUTSMLNFGuog1Ej50x8c7UVstei6Jmd6z1QXMHqXrjQBKlVe2s7dga99tlXTi
QxI6RgEtAuDKDDsYPOpJubQSKq6zK5b3ScBwEAiV6oMIj8ZMjs62QPh3j2MojdBs
p8D3B0d8zR3mjAJBfZjqhwG3RQdrLlz9AMvaKK9r+lgsCDbtj2KRmUYW04XdSTCW
LikGC1Z/XyXkGv1cUXRzFnw3TKw3rVupm9su9V9keLyI0ff+FfOsnanhUKeZe9BD
vg0CbN7Z6VR+CLAYjpO57XS8jGa3V+9yaKMhXXNxQUHPhZJV4E6zZ//ThUj1bCdp
63dOcwLhm0rQ5ImZenHeZd8mel/rv9K2Nf4M7ptOJy3O+/3rAGjJBtEhjZ4nBUMm
u/1jRaom55Y9eR72q735U6nrvmd+/kXmkEAdEgf1LsA3US7l+LD6eeYvOB97oIE6
fsyAQOm94vjAt08R8hBSnhsO1z5z4qOoKoXBbhphGLX/TIL4jRvZV2CLHFwUsRQP
s/c+c5VPo+2IY5cgLTiz6Z0WZns+QO0F/z3edhZbvR6aL+C0rEMSgjW4Y+pTV+2u
9oGgEG9fCAVV6AFZcWYyRsZUWaNwAf60F2jD+clGOe76p2nG4MIJKsolVZ5IwOcK
QSfZIs7HrbrmVvkMTds+DjukpGrEDQpMvAQwk7rugYpg8AO2gUPSJCAeyQmyfj8n
fD9H9sDk3Vnq9Zc9CNRBr7mvtt/6cyc5L4xCE+YvHMeANgs44Tou0+5l3BkhSJDW
TTBNGJK1QK2WNer/3JzW+hhRH4yjmVvibq1FhXwOj2sK4/Gr0zTCnEuiUMcdP2VL
y1QtHoPzvZrR9L0RUL9C8Wi3jHTY18fj668Q7b7oKw6weO3c7Wx26jVR/8nYs6It
CDVso6pEf8NIvUng1hmt+ON1X0fk3p4QLCqB/wDZkUuj4hYAZYwbXQpoqrEpbY1o
vh/RzddXFDmIpkAPOsqaIJ1ThWtA7gKEFIKIiMG7Pam0AxTU88syVk970AuiTXMM
7inRyMNY04DDEvosUH84M6jNrUmBOyoHsmxVoaGs1upW9M55WTSY+JQvSaRTM9KT
KYe6TQ+/LvKE/l8hq5sP1P3pOYu1yGryjv+Jfc1vjQrJMkYi6jkcM8XM5ulIUtnu
ilMBdsM8ef353Yl3Ok9mzcOrE40El488ElyrBm8NU2TFmrnsibG0229WZrJk3JhI
c1l2gZsRlKbBPe87xvuqNsBrCixLEHwOmXZ9Sq9sawEgr7gFh0npIV5hLypPNfAU
UDi4OHWA3k7qIAbgTJqVLTGl7ToBX2Ra6iaXSjciO1tLhlJ8mLHp/xiAoldHgLvJ
gXKsVVlQ3gDFCa4WiduKtls2LT4NdtHQOjNig4ve2OyhUmKvuEvWXdTOIZWiUQ3W
WaieorU+jIdie+waj1+kHrSywTBk4etcRtfY6slWz3nx+WSfThF06sM+fTioFUK3
KMy7IXsOEoLogIkXAUHJ0OHQG02FTYH6U1DK+7AU7OVhgBhtITENG3I1h6qpLbd3
mM/l35Ar9++Stq4KGoeqYO14dX9yC9+NSm2IzopK8fKSvqhVD8Kl3BRvTTeWs4Gn
z97ND1XVTqAaP+nDxYp41hKMMu5jDKZBBic2QZWr5UinhYn0pZmuVVK750X0eqQC
KRo5d92J6QOXhirxgGizuiqwxT8QUOM3FFRZWBGmeCGPiVLI6i+r8rUYdk2tnBhz
o+liAbxw+5DEbFVEB61gmpRJwYpkZNde9RU3DYC2c6rUhEqvZnalSCqgMKTEpHNu
29qjGel7c180UFfYb4yri90jOjUxI2upd8HvMmOSRU6e4qX5k3xHA1lgOWyykEoq
EaObK/Ktt1qw8IFi7jJyIGyKVUc5psj4RTNhDiYRfnEHfpOY5VRO2vsg63oiHiyG
VOKG2/keIvWUa03nguzW9jmwDUGcsEX+emuWDV5yrQpkcAoM2yBNcysQBpsoUTfk
4Qwz3Xe07bcCZk407F/nhhngr74dgmmyn4LJ4ppporBTpu0eWAeztaLQ8UEI2EFt
Q/em12ttmCv0eCugS5hl+cfFmF/yBGsBWARpoORCScf4hF/P2qOd/7U9tqCLlP/F
t2ecYKT+pYe3CTvav3Yi6u10/p44riO/E5CeULhkf4YzZectGYm6JJdVnu6mtEDx
5K6nlKPDTtYj3XGwe80glb3n7wN6RcSURLmS+B2sC3brFxVEFZJDzs2UGK8eTcQ9
QYtqrMqlWh1VI0p3IEXhoewApkpc9voLffA2Nav/sh5NXa5snITbW7VT9PRoTepv
l0u89LFNobT0gB1lnGDgfB3UjeW9ZcFD0X5N6aDFBFAI14VPuSGZXoBhNayxzs8h
hW2gSLLhQzmXc86kTVKnifblDHmo5NyePJiDH+2Kd/dRzdFr2fHPWvB+voQ1szwY
CT29dsvkR5b0Ne/kRUuzTcsk5Xs0C79RaS9HTxV3y4Y7Gs883nawx/W3ggOnvvmL
sB3GxHhmtVG629obeu5B5HI9zRbFgaVBn/ru+BaTdOB6HawRNRC1QuELfU5bk7GH
DoH8j2HWp70ktP2dq0mlPkRUi5Kj0xxDuCGU7stUjlR3y90VBxDyigEo7LWS0/pR
9Ped7EkHjPLHjE+IJKfTf204VW2u1uApU4ALhjZL7R0oP+AufH+41ppWRVI7xC8g
HUyF6Qv6TeBZ5Cbpl9M1tNU9unKNNGeVFV7qmYdmV6IRdGQz8eqgQlEbA6lz4MVJ
jonAuKO8gX1Eg2M99F6BPojNyq+s8l11ltuWK1pjbDrtMpM0zg3XWQIBis4X+uHR
6SmCNq5UBvO0rGrP/YMUjvCFyMEWpLhnTuFBsAg0mA3OypvC88kpD9yM6o6I7+Kp
heNYLtPXkP5jBwjTwFLoBU7wY+Cbbx0Ho8QKSAy8l5Ck3l8x6TAMcHKQpGyun25w
a6H46kkn1xJYCT4SwImu8Sa5EO+WZnlIsRZdePwLX/cZTafqsjLYO/lioloKfPH4
iq2twlTAlG2jB8iP0ZJc8fOAyZnUXajJDPUIuOoRJvQ6M0JX/7UXZLtMfxaJxiVz
AmVy6puYLjyxLytiZ8UhGe1NB7t1/kALHdJSsCsvI4MPeTttYRN6ND7Oh2vDULNR
jSN4NpwX8OeSWNCz3Kv4b9DKKG1MA/TNvYqUilblfrvji7Ij8+zvb6rlvoAvJUUZ
/3v4s8iq49RLKgLwHPWDRTwPO1qrzVI1xr6cONnEW2FlN/gQX6+q8QHKqT80Pq9V
EbqKz36141EFS9aVe24WFL+5ZUkqeKK7LBBrh6Xz77OeLiPkMSwMyCGxAYw/QMQc
bHx2GDAuHuzlrs+Os2Etct6OJhbzUhT6z52lI/euERWH9XOVx8386rVHtgDRObEE
TDKg0xid5rmTsJIS7VgbJqgB4QW5QT2I3RSbg//92faKuF16sCoQBURwqqa+K6oe
P5CGBVGrndnCsj7+sQV0FJWVb3ArvNKCBRhaJSj9wr7+AUrkokMF8wnO0m/JPEzZ
L/1poM/ssFULFu4lCjZc8dW9gWsmwvYBBRbdrOZXKdgASyXrcUIqMEVN0kNwnOab
mxIkjJ/ug25Cehron9kt2j345tuBlbPmBBMTR99xxfFn1vabZmmDKUDOMQwmP44b
tKeVm4zZDsO60RD5fRS65QRc+uxu4QqPS67EsozBNGd46QYeG6jda8ipWAaQVhCk
iv23kQlS/6Za8Zn9CPJ3luvWHS9g/rmAkdQhQSbX02nqQGesEEmIbrZ0Ek/6tIdN
OC0tcMMxGwl1QpKKs+aEed+dh01CSUCRZMMb3H24nUGxS2U/jjbbgXjwXswJ5Nwn
Rq6R5dkBt5YL7ULHqe+yKldOhpWSstH16zkh6uGQbBhrq44FBGPEsjSHqFWedNmZ
8slnfflWtH2vHEj1uWEaDNAdFJpPYkZuzOEk8fJjDEdyePvMjiYHLZwKAMU8B3ts
UaflieRdcLn+sUaefw5A7HxGOyKfQGStDQp7HM9x1Fiv09o2jNITh81YFg+Sru3u
7n23MB9Itmx0gjuRGJ1ZQMxyl82B5D8GRsIwLk4IpXbz0wtYYkXQbJTwoOeda83f
qLxJa+Z4S/7nkx9asaPhB371mPU12F1Ipck0kqqehLzvy5ngNsafPK4Yku32kedH
nyZ8/g9LYGHIrJFoyThWnGwiwKplotaUANV1c6wJPhH7R/ijDcNsdEjkGsEDZE66
UEbhvgA1bHFuuQFjb+WID2bhYorDHoAQ6FbNMxfIj/bpHslDEzlq3G65xLgb4Z6k
GHWGkQRZHCA4d5yMg90RtcAtDVTHt+LEbyNQDd+Ryoi4Oap6ktUWTIy67vqT/nMR
S7ecqwuwl6b4XgEe6Bx/V5IP6r6DiwDv59JGYlPcIeNhQhQeiiqcIhOvQq2SRnc5
zUDI/PoGg8my/aMN9ALqnGLb1RoEu8ttlEwPjuoeYqPivSS1vLk1mQwz3oCOWG0U
ChCna7yPZ1KnbKUiKst4W+aFcrGlLaNrqtE/mH58B5LDDD6kzFyB6vsDAQuW0CWX
wDgLm3d2Cw0eije8BnBJtXuYz6/+3NgjpizwtkFO7ubKyYvFVZd+TsdBgV+kHOR5
QQOG9CLyaGaDk/r84dPKQ/RPuH1oPcuUurboe4+R75rIj7RiDh1pAHgXezG4eAK9
gq9Q1/hLoQQWusQHbp5QG+b3k3JB8PsdpPC5iclKgupx7RbUOnjCI/MydX+h8ESb
7gjxjHSvmPNYk/AoWuF1Ww+HFN6RyJHfrn5fBdtnlfqh9r5Hd2xf8sTroGrtzofb
7geT78RbCGHpuhnXKlYIURox9Yf+urQiaeVRvyNQ5r+QU0x1b8SmkOGi/JvVev1l
BpAH0k3sbBaI+AhQU0NKr8Nw+N51GvrAODu21SbecVLbukgmX5QKmGCwR/UA2xu7
N4MywRtYPH62ZMYGvwML+D5sbdP+9YotTcciCiTsLZ75YD9p4X/5kO+4zp9kEnfZ
TBGxBWab34QKKflQW88tZWWqveLQP4mlqXYW/nW5v5PiheJXjsm7v4egJJBc6qWm
KNwnoyxzbWRW/kKJACv/ZN3jo+g2insVZf+EsS6TyOCDM1MvWovMu61/qi+SsxYP
q1/QJUKAiU/1F8vtp3rSnLnYyJnvGOrhvB1H2AqxdM9lvqey68pU0qp05kptnMSX
tUfWJGov9pOiorcG54IToZsNQZKwfA7bpA/AoHoxHLCHfAMXciF2b+NcGOHBVd3O
1cWs3Syifpxk0458aVTFNk/yVD8W830QWIbRgXUaBNyPkK0QljTisd1AIZmIivep
N3ilvYKwTb/NokzyyyqkmfdyS3o9aEsKFNY92xkp2J++Jibkwlfgj0AKV0qLv1cj
Atlz5zvSGL0GDrjfWpBeN6hhoHCDX/04TRsccTPPCgk5v82gLdQ+ZobwkozEewfp
4F5m3Zspo/6Wh2NV7a06tYu4XgvDW9V3Pk4AyEFwATSlQT/KwXsyXFjcX3bF4SuA
f1DBlH3quMV7Gopc6V7TRp2bEZ9lWyQITE8oyxGAOtSfhDUoaunB6OKjfTUYqrCH
Htr8PdZrfiZ5wNJUhdLZpnpAM6HGDuizkQ+R1mbMy4n2fgDfyufdWPAW5Alhuz20
tvRPnj07X+6HmzaK6qVYQIP3CMtJ73NWtnWZaecypBq2NgaM59lU0j134kgS4O23
jksyVJiziscABfH0kh2qqXfp/2zgXso04E7MojTeL34vk3XYjT1NHh24UuriC56/
GLJRYViEBf08Co2BUWu1aKaEs2F6A8TS9vJ/6U98IDzQQl0I1O5LQn+jQkVXeXvk
ZrwgPlqj4bjSrTcpqMZHcaGmxdWpxCQ8IPzcA5QeCKSKmiWeasFokRdfvvyBXIhM
ZAgxleO3sIr+/n1rRw9kOy5HZdxtJUwpeJuASg6SayOJhm/nIOMSJxmMVePuTyPy
C5nRWEEVc1MzBrZmS9utgPjUIcGVCuag/YTnX2KfjXKZ0KS1QWbp9QCgTpit8b6O
7Do/t0WE3SMg5LYnrrwt6r1XBLCJguWeCUuHAbAzK9aA8owfkVKf4Pz84c1DYFdT
jv5+xGByxvEayPL3pn4GHVK6h7g0LlrY1pHZassvvpe5zWzzdlkcf15Wy80G/WN/
06++0WaZQfEQgbBJcGRZ7P8rt5PqSiGVx20emcwrgMofmnKQMJNSXO126T9Pwri6
yrlweSo34HdMK4t97l/Qlkqd4fwU9WjtVtCCxq2vmHsJTcFgtJwTk4Zwo+pyexru
kbiK59SIo48z/3jRaT6rBf3dIJ5rcUtrURpxM65CqohjSFbz6CZj+PtZ5LTbGK93
i3INTihLWPXg81ifK4J6S4vaLyytDfZWM2L2bEla3wOO1NjrhWW58nhI+DnbPlP4
HWZLXRwnlkfZSFADAqkxXPyNwCSNr4j39kQEr8D4MaHUaUdvKFTdtWbQVbI5aqSE
BwimtVSTZk6qmZ76YaMSH83i2zS0Z6wcQIDxSfI3rHzA1FuuxJFCDvLFTCEZYzFK
288Cd2gYEhhtv8KB/d9YnGSLYd/C/aWAaV0ikFRUhOJH0iCItORAfdP6xtoW2nDq
Dyd50iOyVnB/pY+lrO5Ap825/SWmCKICTUfYTlFBuqycoXY6c5ByYsMc2ixRQ6zv
TZnrMhRB+BtfC1Y84zVFSFoxat/FCyR2JzhW9nACiPdigWylGzx2GkM1ey5Vj+JJ
PYDGd4eC4/NszGjQGQ6wl/1jrl7RofUdseY5VBpEyYDoZcvcSwZBuLVrZOsQWeK2
bqvZY1qU+4iVKwyUA5byG7a6Sa6cUT2ZO+BXLJn4uqsOGnFoYbtH+8G1zi/MUigF
xnLq62+lzOKPrgjppp0ogn3jiHquprBnLYBczbqsK792VNK1AM6qXYzoWfvY2XRJ
vT9L2wGqFEXWZ6en0h6a9xxv5q9cY4OCiib8axiMjvAvEJ2YKuRYz9OoMjXSfFYa
y056bsG+2vtiEAL8ug+K4mFJ+WBqI4ZV4dRPu3R8jK70cROAl2b61WsFVq4iFnc+
Ip4hp7De/ioqfrJtOw9PhPF/wom7veHtmksz+uiDxOB581xPNaEZsTg5LJSvx/K9
F32R/09CEW9x1dP28f20K2Hy2YT7F4Tc8dz7dlf1n6MjQKRp2uN6Yen4ZZDJmLZQ
sorsEMkz2asKIcnGpi2QTXrqfU+uhHRMo2b+H5I8AcyHf5qhDSG9TGQGfiaHTHJR
aHseLaI0orKQ9xg1cvIpgjDB8lON8SErZQqmU9LZCBK5kTX78Cq0cLxDIPrCOgWR
ofF/P/g+THwFv9CbFjDir1rqXdb7W/f1Wq98SgkNR7kLbC7FOUUXH7RBGd/llaJK
k8ACGHqgMGZCeznzHUW2sD2nz7YY2zd+BO7M2Yo1quLpx+betrfMNHvD8xA5GPZz
3vj3voyp3djoEl+cN2ao4lkue/KWDIg3r8i8pfCza6GFgJ/LuQZe6UKygMkAIZgH
PSkGS6ER2cuJebGUgX7gzJHTtboP01ifwdTdJ4oajsVad3qZ4d+u48lKenh0Fk+V
gPa84XvPXsiuvzWT6yQJ1w6pY0OghZajxoA3w8ZFfuyh4EgpG+dzT18RFkD+1BLX
n9jbk3VlkK4vfqfzKAY2O9UDEFtf9ZMZI12b34Lxc3h9AtzuhhYgdxUUTz13Y6hS
MeRrfV9FtNCgOWBfyOzFgL6SFvxX2mt3A1yeT85BUSNesTM0RfhJGz+cgdz79bvS
eutCPPtGPgPpJAGCHCMamqT/op6yp8CAFuLQAU4b43EuiqAb36sQt3P0Ry0u0qdU
Rxt5L8sI5tZ2qnjPUPRylbEhbfx84K7Hk28LUP0nFr2wJhMst+/6LqZaTe3kc1hD
RD7xBoT+5a3RHdUsbjf8p6CE1FVqhtl3LkgTYKrLdnt6HsJdJULZPfmKO0fwJ4xW
ZjDN1HODtvZ5jTH12oXZLnW0+qQjnFUI9aKTWiBkChzf/kdlQD9B5z0lsqJMagtk
0/MymitnvOZ1LtnX09Gp3EsXtwfwlT+JhVJFIYuM5VrCwwBPxyjYfnqb6G6LZnQj
4PY5r1lpkTTVyLLJ3nuD0Kmcpuezde5ZyHusFFl401Tuk3uRpgPO6Aqbl9PC3Mj6
jDTi/qJcVCE1Yn2kncSwlh+xhXa7uzNAqcpBLz1lb5jH5vpR/5ryOchwFw3lIee5
nk44DZH3uk6BHYXpSYqpuph1P+Y1tjXK/u9q/zc0bJ+CVOdQu/j7SIhD2kZDL5M2
+r0tfC97vCPN5D4NVyUzdX4IQ/37D/dt91Z8FCvhLEJvmKVNxLBiu6M0Ryzj4CQn
XITTHTtWI7Aya2APar2tmXDxza0OEbsUYtVhrrk444xC1gDQ8KkMeWGZeOOBE7oZ
PAFo3rlZbsXQ3+KMNq5HrLG5T00uz8peb/GF7hXmNOPaHKU6AIoqsacTncOcfcCH
8ykbLDag/sLaChrNbBwdd3kymePqGwuURzHFxPu84jaf8u9uSKXLeVK9V4p2f1uP
/eEs+KyIIm1d+RktakdIlp4lYpr+PQaZlhXjZyPUKi78Ay3T4tw/cr35xPmAPj+7
Sz88BsP+pXC4DLLiN10dLReK5Ddi8gJ1NROVGO1cPD7oaRbaPndFrzIV80g9szA/
niHx3zbxt4bfH2Kq/ysN+u2aQUqVqX7VujPSPJ1zYgRROe9eLVNUpBT/iYpOLeb9
rPxqeuMwoSaFvR8n5s74ArYTMHrXXUoKlcvsOW0X3jHbNNu5NSU8YI9g6NCdia+W
Yum83SB8NpSOQ6ov5nONFfX9m5r9bEZDWjBJY09kpnzklRznT2MqNr9qxzzZiOy4
MklxosifwXnGxUUs4uhnd/ALlswX1Pl50Ya0hBcqLN6N8JmVWGGgnKNT4Gv/nSGa
MJkGj12US5v5ZjM76VJFvgA1ZIEBckcGExJRMtPeNQdaWbTVvnGWj+bVmvOB7X0E
U7S40qgJOXJNELQ7mcqNTde8xFml5oGdLURin7es9kNSfTHqhLWsUEmpr6TsDNmf
E9/aIrQDB2c/8RRG3yThVt0ZTDByluaUe46eaRJp5lhSzMxC2Ap2oCIbltN1VZmN
d10TndE8JuLYW1orl88jTIRG65WVgUAnh4vQcFXD+s1CvXuQmbC/rGDoMUzEhgn6
f2SQ3U7rrpwTfXwVMfWvmzJQC2OnNeW0trU1ICh60NuiIowRKQpIjMwlYg0A/cRa
qhQaGSiqI5Dx3W/kPF46Mvq9f0Lpd+c6kJguwaAOlHMyDbnogFxdarvR1WUEgPTe
DgNuFMPVCu2VOdAQNyunjyXg1NHp3jDAhEOlZGk9ihD69DLmA4A8Zdn0xDsnlcge
NI4uyqAGlITSEm7WpNU91yIjwUQKQ5qMUiViwAdQ7yeisV7Q++T7SHxlZUCygBVP
U9YK7VGYbrg01SgQ5EoUc3IADLZUl7VDdVYnxJ3qX7tJFA+XRYLGDEz0rnVGPMGq
ip0mWHK8m5p8D3o6+F+y8beEtqQk6zG1uBDUTqiAvNLhQRIvqe+B4crlNjnzjikP
S5gaDyKKlE5XzTirLX6JqtJeJOly3fBnNNWvCw6Il8Z8nElOoJ8qy/8egG4kn4T2
L49fNIBiLHyLpD4f4/xlobCa8+0yt9lSsRmZMpMPhy3kPMm6CGu/sF4pBJA1t30S
WVQ/ziljaQtuLZRBcPXQeb9L+i/M6vzIpy++EIrqaUndols4uCZcIjBwhP/ZOdum
tM+E64vnYLLNbBnulwCDw+tcuwiKmSg4gtXpbQlGPwCUepKLR+5zpOTugpTiKhEy
sgs3q4ZNquaYEKeov8kzSWywrrxlqJkHx4C0yn1VGYo83bPxv83PFC/sQKNzRg8g
ummUXsQmL4zvozwLUUzwZCu1IgSxYclnDcJQbFbE3K1EOA2OJ6aKwPCtooCGEybW
X5pbo+MKame7nR9TTrau91aI3I2rjXiN9P6Dxtd3ZBG0ZjR+q8cb5eRp/hG10vvn
vNvN9QvetsdLsuFVE2jyd27o4nWA81r1XTKTZRuSZLfBprSbPuY9G3CsegqSivLs
9r9ua0KIqiMyYi8rzfIg5iYXzKTVb2zdWcAjZZrxl5GqdimgqX8CTT72EuwWYd+D
0mjoBYk+Bi76YVFb7U4daGujtWT2hcC3H3CjrSekPfwpvtv3iCZ9fvJrlIEy/bS1
0O9evsKcjw4Zf3euNHBB01P0QL7jfxxWzdzHpTj31PvW4N1aXAT0CnYZoI8ynUKa
s8PaejilMVP/CD0czCMd1KaEH/R+VTM1r7a4reFXz3bkI/ZgNL/NCaUd/Fn8pjyH
0z9II6B23qiwiwPnfQDNTTESmaBZyGO7NUINEG/IcCBXLzPMiAyG5PZwOfUsEv3n
GkPQB3VaUaHIr1R4VHZqtF+mtoEhvj+nguUXOErgdmEHMgq0fY8fHs0dVdBYI/85
5+/FJU9m+Qim7XXaHg+I7Chb/XlGYKg+L6nNw1gOpGVsdVWNzpfer6aFowkSbcpt
maKMw/LgilYX3tWkVXecyLn19IC1mPKwn928pJafYCnWJJ/fhQjxs7h6LFULmt6X
B2ofQJ6FEXvo1K+S2f9UTqsn5XkHSbPAOXfFE7fXZ4IvE849vzrToCLo0pyhBVaN
EpwEGHUdpwv3rqywEkdyM8u7TOij26ukctL0gO25y5BBTrTwLTEDT7O6o6whp8PA
VkwNMWQzRuQ6Xm2u60j6UBVFPQ/HyAkVUd2RTsRpIwwWDorZ6vKV3GMO4u8fB9y1
ele1h4+RFNGKrmzMxyebiUupwb4J7s8XjReJ0i9POcMXpAPSA+4Fg8ZuCim0M4uC
us59j3wKhnM3r0B0Vx/9V3Iev1u1J9KBN7dFVWaDVeiL/II5mIIaDTrkDEA5U+dX
ZgT9NqZzNmhxX/kPZg/lOAJnszf/Ts/h6cphu3RXA8fOKPVTnDZi7eaBS8Oo4G4K
64KEXmzyNhMCO+uEAuYyNZTbaeN4yMzO2jdeswPX1hKCN8YyJuzAWKSmJtQznw+B
cRDO/rpzKmJsODf9e4G4/ROah2n5ij34SCQLLXPv4hFqYdJAUO4OMFh1Uaa0Sb6r
oD9T/T9+pc0BFPzyjmxIkgSeGmGjWE4wceTWZp1IYPsDTfB60juB45tUzv27NFly
icaAz3Zo8IXUVX/hf2qp2Bz5AeRpsa60f9rsnDxR1+S9Ind2ZHzpuVdC1L1pM8l/
W70oFXHoxccWjFLlftZOEO9U/bIRunFTpGXQjkL6LSv6juKfWvuce+SkHEbsZ2nU
RZ6H0nGY2qE9YV52lqfTrnd3yikgJBzv+XYoVj/Kw0EmnWI81O1JNvV2ZjN6OSQH
dPuQu4IMFyhVRYVmRg0uUWfUpz7VAoEqvC8jH/RamgoCmDO7YNT+aF4LN/62nwpK
R+rsJysodXsTsgXBd6Nw/Oqc1SMzfYlIWpGcb9o26BrYl36zAAxBYzbLKu14RYl6
Edf4voLPn+56QLpehdhYC4egJGcpYeK7jIekTkJWFgXhqGavGKi00oTI75EnViel
SufF/mCX2yju2ovHYaSJS4uxg2ZlO7FfyHDgsZ9F/JSMq/1dPog1TsRWU9yq+WRT
1dARqRDrKrflBYnMGTLA8Y5sGQxweeqkYsUzoIbtpAr3eCn2AVCjBJQjZ3PV/7O2
+KseK+wmBEY/cPh4mGTZMq2ChlGpnf4+xw+cryvfS+c3toX095bEnmhGVo18aQHR
iD72ha2V6kEGKHduZD8AYvFx6M/EFaHfhPCA140wr6m5nXh2ycBaJ4OmHrX9Dj4Y
OUmVFESnSIZ/8nwsL+mau/bixoEBJorum6vWeT4t/t82jySgAR0isXMqOtrf+lEA
gV80VhdGEqNv1oIt3k5C+/is7dGJVRikE15Fckgyv+pwlS1EwOsqeSbYDQgAnhVB
dG5D1pDAsvfQdDki1Kkgu7/qYwAVgRl2Ao/Nr9pDmejwrn7qDNOhoU4Yr2xqZgCF
3RTl2nzz0rNg+Sa4pOdxGEeWMlGuiYSh+kv27ybo60GiuMc6UC8nVKJV15bYNmnQ
xCiYPS/RC2U6tDreTshH4UuVGVN+4ePUpa/VUh28TKLuIfWaA/Xvj8DmXF82+J3z
J4nWQ0WfBpXsmU2mo7bZuKjr6f8xVMyOqFIWv1YlBxDxoV8nZc4bAIniZ8gt7Cd7
aU52Nz/qk9QcgDfqYVxdsVxXZ+7JC9+arShjF544xWiDX02QEsLGNJc6xN24w0Lv
UCYFJs07/hWBm9hB287V0ZEYLT9+oMKGwXbJ8WgNU4AtcxiFz97opcVCfBu/1Mmi
IfY++19TahbkRdFT598HbYjlHPzLHJXQlX8pca5XDI8lCqP+E+20eleyKPFFW2DQ
a9/wOOisyABBqjeAtt6l3HfriB9rLp/lOyvD2PYbJ9LTIJzKc+3i344d8y085VGp
jFrs9G/VV6nr0pGFxY4UdmzkIwnOn1flrLA7Dj1cNweJhnG6jz4F5HjJ95mf2rpT
ioVgnEtD5xHssKBm10r8+0Xb9TXb5lhFS+fvERUDw3LEQt3nkHt6IMzkL5TV7O/Y
7kgw3jqhgHXRpNZ85CXwGkvEPPJpjCfmHsEp4Nb2sg1qfBbGVcfbUnWD6QcTHOpM
oP+WwiSQwtRwdNvyNoU1wQf4sZE2DNVmd7V1VJv2Wm3HhOqTt0205YZDDDS94MQR
nHfgIuSschX0zoZpFrN66naDTWAkr39liB7Z+7EJRaae04O03tHLxLJundaLdM3j
kAdeNsV+9Zj+3CG+Fj46Jl//EcV7yp898fXOOmJbI3u+WR+vUi+EMn+F/c3Hku1i
oLVmwVVYOxd1cCz08+OxIn5jP6aB+bBvejTRsuYbCFaltGCqOFlhu/WLl+vg9kIS
o990lnPTbE37Y904gUkTSsXNEipRjP2QVD6AGSYeAqqpK+KQCBUegQ1UioKETnuM
Yy8QqXLWZdD5RRtWU442SGbPvmABADLgqp5XjEGpa+wcAvWB3hUU+Or2/M9EGih6
1yXR5adFptTeh0kmmjJGBkD3Kmnw4Lvk9Edxd6FUOxIlmh74//Kv8QAFzguTZt4p
HVGjYkjZXPv3eQ8PXkN90iNX58bB70m4wOl+DCNUez/CdiEGN6WWK9KTx7/V5/eo
vpAV4Rx4xND80Zz7wpdLeHwNO6Ye7b25RnmIyxF/QxL8VcTzVFVCS0Xmkw+EeKf6
hfHkdtv/P5wAqDdmYoEx2M8nCpCeOBAAnV5m9p5EpmKChtL3E6BEdxCrHu8zrd0w
s6SumMbxqw0lywgS+DJ9VkwyDgTgckSOhgAJbh4gx4HbEdnQIZEFS4uCJduteGZw
umxsNChfNA2G73I/y5UDe1G4C7h3VnO889Deiue67Q96oESgHUOvjZDFdA2uxmj0
balpm3a7BUvAP/aACjILWCY38neatCreZXhz7LDU+kceQR5W5Q+elUkZHbmFWTnq
aQTeDvGejg35HAcQ9htug1FG6ph31MwfC098S/JhyiVIM6BZp4xXOdI8yLKAugrB
OOMEQXvlt3qp7fLDYn+CdOH5dwGGXD829Ccy5QrQsf9AlbhIK6e7Q/n9a9n3wrZb
0hGtdI7jxi1HtcDd0RYUyri3ocCYEZ6ohYOHjguoKdqs11xcposwyZRQ/6f4wGx7
/15pJYIfVOd10Q5auQAAAL4c4FqpDjM8bL7Xpb/lxiaPSSjvhxByLKAKcONyyAPf
GmuGKNODctJ94FPnTm6fQSu3B1ILLySDAHUlCfMWXhOREd0gC2A9LAnfU6C5HFMn
nGjB07M6i6ByA5/214iFBxmBuVNlv4cJhu4Be4KRfeMv7VY6AIivz7bCoBX1Jc1W
BcakL3Prhnb80Xigg/wpapQUImnIToW4Z/G4p5+V8SIA21t5dArV9vrmWtwbm2Ba
YzWiPjQxfHc8jqIu5STi5O01MPmI3MhJ+8PdzmeMZ/7unNcV7qj7GZ5XHLRg1/Cd
h7v+sanl+jFjh4FtTlZ6XU3RPNrOicd/ooQ36BVtsxXgnr+2IiA9JpgCbWIGADXn
VvKs3iwmcm63aCfFyZL2stjQ7hZEYUBiQH+tclUK8KPmLrvhWx6QExENqie4THdV
iKfNuKCi8ik7hMzH5JN2zSv88RsrNGQwk3OAoeyZud/aMrCHytCIdyt4rLXaIKW1
LpqMIZAZkrTpEDidfh8U3j6+0oSXSOsJ54xN90YTQsiVsB9xQd1NsJ35LEHHgeWi
oHBZk5j+1SgvQdilXzP71rq3mA4AZSTOw9SXTlvLb9Mh17ljYyKSzCbtbH0EaEhG
klQ4zvyrfg92v9TSMbTBsx1EcumM3diSlzfPNW707H7tIhlhv4yvstgf2XpCZwAr
tXIQruGvCA7a2pyHSJ4OPEtwP09jJJcgRnbTTIT0IUxIyiselhMTYFa1V3TjgWYs
hsMmmAt5QM+YlUR/F4ZBgdgO06W3Nv0JmfzfFYF1O0Kl+zqJQQGyMNHpELBFHt52
GlbGjZr8vZNLK3ayrmd+B3Mp2N24BZjEB0TQN4oj/6U5ORwmk8H2ZFSvsVRS5UH3
mrXyWou0pN2ktALmxZW1dJgyYSX/INxpVNz4i9ZpnYDwf9i+a6cwPYjMLY1Hwruf
QJsJA0qfXGuSRSdFtKXQsDdVOx7BXIdUIH3m6btGev3iiSEl9dXc93VPQpLNZ6MQ
CrBi5iQ2mxzebcCqfRW3tpRpMsTInbq+Twp7lTCoqi09xpGDTLanegXcQ+5xU+70
XlMqubDHlWWF0Be1BLw4fgHyJmrfd3H9ePLwoGoEOCtIU1+SzvYnnmXk2awy+leU
ARl8PTi+bgVvwZiwymxvOc89IZw8iVcZT2CtTOIpYzX6T6tgXYocTbSUmBcPnj4b
xtk2NTjP1Xa+9c7++DmkWGHD3fFUxWVLZf+YqqGiKuxg66GvBrv/g+H1l5+h4o6x
aszamPMYT4VGjWQRwJGTsO8O4mdim6GVAjtaRfb0UYW1Ol9AmKpRG+7vfV1qHWKl
E9/gSeaQgKj/fKr7gK9BKHmKEYai6+WYzKCeS7hcry5aN/F6kl/xGMcY4g2CxQVY
JI1ny4RWZ8Xc0RLNVp+ur/RwJerFGVhIiO95vmt/4S5EuSe9GcMo04uYpbiNSahN
1Axqa1UkPZSv9joInaLzFrubVIQqh69NL+63XjNwF+CTqN5dRuS7CghgLqwgdrhs
/pNzQWPJC3nsgaftKp05jLFi44U6sbZ/yPRwJcKMIYYABsziGKyyYQ6CFRj3mHd5
JM7MF2N0SwBYWyZTaL0SzOFMG0v1r9clCK4I601kuR4fafS3xE9z9hhtKL1wg/gU
MScLHQWG/lGAspf4KtoVGSWrq1IcpQnURjTtBHTwN5BRAPL/WN7o1a55ENRSqzQZ
KAycyB1n+tCLHeb5nks2plTK5KDbbpcICC2LD4qoEXxH22zGHA2CA65L6ZMml4U4
blmiLHVzQ+EiMbR9LPTmtXyhlVlwVkX4K+iqybT/Hajf00N6HbrxC/VTr1hUoS4f
IZu60jPbC/D4iX9tBV3Mbl+J6YCOy/+U6FzwN3J9o1v8w9llzpdmSUeHY5HJFAzv
dCsTKPdFPWAz00apelSd+diTSyuevcCGDwNDQ/0ntxREODbYLwygM2HhxTPbh5q9
F1kHwdhEQ8xZGDOJh7ktQQGViZelctDvGhOseeSRusIpeVoZtixCJUuoR5aTBBuH
N7mxz4XAydn5C3NlPNpyg8nVdVAZOitw90SE7/evphPy9qfYX16cgl2T2pUoWLcS
3F5GdymaVOVWP6WkGJhRp1d3Grbzp5SDXWsZTfjP+/WQqDWyCQE+mvDv0Q8f4F/Z
VKERb7kZDJQ2mNNReH9Lk3IrX6p5qcS+iKlGX0Y42bkWpuZ98OhnK7RZMeS8aK44
UG0gWroKWhW6zIYimFPAgUoZ5fIoAdImGq6kkf4dPLVGrjubEyuRrowv5giki0o8
+xIa+Jt29mFpRyFM/VJFpAnLGzJzIml/W9oRPwxjMuTZNTtIWZpEBPaOCNTSIRwj
1P6oOruk6zwFzg8CwvVrNRtT+rF7BOgATRY/FdzFMAm5gSmj6vH/Lb3g8ytCN9Ht
0cF2BjYpGzwf3vD9PuSCfzItyzsBBiJbi7QrsOKkNyTmQ/1Yyyi85VL26n4nHgl9
k5H7JkLC3vtwPR/xrelpQqFfjsj0vi3VS/LMAnkxZfu4e41GnW7t9Y+hEQLMaMcK
E6nxTIZadgEOSn5AlsKw6QzFxkMhYUCLqiyBSZKLOFNAACzqbk7rBV93xwiLq0wA
rzZD1C66R1uT0+Ca50Z4AULleLgwSslB4oWxE32kdD2iDy8AB5YZkP2WtTeCpgUF
vIkCz8asYXXYzXD7b4nodJLQD7xCrCj5sx+1gLoWL3QKrqE4OI6c4ETJnbXKAxcj
TTdntbvg5mz5LWyxEoA45BD8vd9Dl5Owa5wY+4KUNkwhd/4AE23g4F1lAurvz9/z
n62AZmZ+ho4MdDS/8orq4dY6CQbUiUq+8WNYihiMHyltCzk5zvxTSpdKiDFrRJEP
DqHMMiGLxgqzQeBYl9AeRWkWcxB5h6KDW8dnB6kQPcqUBeD1E6MdEufNR+EKapA1
TEToezu2YymgpybuY95Og0iRMWtyBtc5GdoMpDJo3SVWYCr2JpxInrHn39BG2MNx
ixRNPFAgoMyxzFzpMcbyDAjqCFB54899m9WJoIlwP9vtPWwQT4KMCVpPNkXG1SZM
5Cn3Z6xYZDZSNH0JnksDXrfIgpmi42emZKPbL+YyLLs3yoKbWh9ELptboKBIhMS0
TQEvm2ycjcZbVfMNNMVBcjKUOD0tnecUEyL79MKw1Qs0XfdLq2N29ew/HKekUCSl
TttW1KJa+9VmUebOp4rFDjtj4HecJvBhStf3GmWxVLkf6tfJKgoOidOpsWvAth/D
mj6hxcD0KoHbJrhdoi9VefMhWXs1Gs5CQuZbf3TgU/ht5Ak5/YeLktT00v35XVNc
FmhjUWaGLdEPYlXH+/dXqY1k0ROhOR/80dS0citMlqK7/CZ96Ye6FMw3EiqYZLEJ
qsEZTiA7Yde16wwbuF82ixKhWmdLMGkwcfnpu2oL+dDjlQZeKOeoaVdx7ip1Jyfb
cziCRrN8o/Ls3uIrQVOJCWPNQL+Kw0pPBaCMPTkbGOmaH0kJXNE5KXYchi3DC0mb
2Y3yPoC9YW/P9Vq4SIXKriI7KjOSupvjKnARUBYqq1vrFEP58SX93DYbfQk0jO0+
U3YIG1WBWkba7Fel7jbnw7Tty5JKrKbBnuIK3Yz9qU1n29euxHjxCHCAIJd6fy0T
pRYNcIVozSGdwDHVMdFYKbk29U4m/lEQvaa+8qG5Ko8wzuMToNXLfPtDTvrU8f8W
80SPCu2ld6aWnLZIISCl+NrhdwScgyZPsI8qhm6qsMW3edj7PdbhBA/eV1qbfTo+
Foh4M6r3TTdHvL9T+jrfEalZDd0m/pVy0YIL1lcUTRJ1InqNSxGAggNPH60IwY0F
YGD4lR+fFqOf6HOESJyFdpe0ZkZe+b95ETZ4pgchGU0SUL1cOTiOMe6GN2cSmNFp
4XiBU7neSgaj3yOQHvZnFcX1c+W4GdGiamsQvaCkOSLArqh31dx/U8wQCuTanqVU
SNZlJiCsxc003oIV6oPadDcH5TKoBDOIdGkn3wsZvVErvv8U6/2cbqxTTY8zirvt
ytzSrvdEIi39v0VvkuabowBz/p6j5X1m1YdeFzJ6VRa69FQlu7mqA2IXg+toS08U
m1nS2xz9eAxuZXFXCj1dGvYFTk21HaD+0RPO3Hnw4RQzUPjXtmZbGMgKGbjtGWP8
guYMMKyD3H5slA5bSHyceATMcSnXz1s8pDX9jyF/qKpBfXDIE4UiYDF3zGUF9Wz/
UOfBIBNC4xedVfPnPmmuWC2OB63CG/MIKA4JbHdyIz1kAA8NquclmXRLp9dD2rMI
Cmesca0EkqZIigKYc7KHsJqbh1/afJ6DPU4HrDe3keY+EP9IKvn8/sFj5CUBs2f6
vhnuyExhExQkf+aA1roeKAac3g3LCRQqLX96xczFYvxc2i5YKgYy7Hu45/bAO0r4
SMB1HhPpEYoqbeYgPq8LNlraNSVvwit1GHubOLhLYHRPBCBJfpEp1sNnZKaIJwLM
/l3d0a9GjGEJTNquvxoKqwaz+CqjW9No7Wti6nUhZM2nZb9bUGRw7JgUHhechQT7
3BmnkWkWYJF2+imyKPHuyXbvlo5+A/+3UTl6R983dFIDWmaS3eQ6wCGiE2qx5eso
8mdzP+WJxu1rLgIM4IkKek6OuZxp/BvsvUy/XGhY+lpOPrczVtc5vUd7k2cOs6qD
Tq+lpbQCow/ewZaYzDizDlnUMHtx5L+DZorLaGpKf68oTooIRqAl95xdsCbNqBu1
m3poxcjuq185mvLyakfF09FQ5rDrfprDSM9NqtOPEjK/Py1iG8KVtDeNZZd5el+1
DiX11FOWW9M+XZE96tpNunC1l8iocjtGa/+8H+51MWnavNk1GGxVX1Fegm+RR6sx
HDje1eJiSYMJGv8sJ1BwTAQyvMW2aQYK0MvoekLjAFWtF3+/cMHI3sLgi8z17rsn
/Keg7OpNADWnjkHDl1rD9cKceOr1jPxOkPBZ6uhBo6eGTx1hMJlNSHGn6ZD4sY18
UCP1CpOVreoe9RbnBs6mwaaBMQlXxkDPIITczAC1nqM4KY2ia74y+QBaRMWxyr2G
7NnyU7ZblnoWiqdJPZGiQv37nM+KfpnDLtXbn5cZm1f2wcvaEuBgQNBdirAqDzCt
sVlxHiAzXz9ncP3/LHtfWGQrbQd5FX0a24X7FJpiduRsEcl7zYbM9P3NP097GHRm
YdXAYg8ATw3CPOIQsMCTk/G/cnEU7TvqCfXuJlDdkfVvHSTEAmW/RjPHP23ms0+R
yMW8rFYcP3YdXGI0jpAK7iI7RnYGXgjS9zfQnf0tHMnJWptj+dod2NE97dIrbXT3
97k21hUfCOZ+me+kO5gkHFSesP4p3xifOEFF8PPEbkHC/8YPlLxQQjVKwBLmX5PU
Wx9AId+iTN3qo1NV+A+zV08BNw6meGVee5ialoaDh+8YBW7p7nuKZHJiOMbAlhSO
A1ziBcIb4RKQqfz5vywgl7eRT0T1br6KHwgR4lryWcnMSwLuabgrJQzRBAQ1XGcq
6NuksBVYKtOc2x+ynGfZkWoFJYN4NPsow8QNsxd2wP08pAsYsCIzdQ4HWx/rNCKA
Gw6Lf+wI3JSLlv1ibPaMpe2RMq3hAuaIfnx7KvMgP1bmywhggsH1y3eImGr7ouBo
OUe6X4hV1PzMLUFSsCflzSEIrUCcjLie5cGXjgsaiE3ph6lLn2/kmgKBHrNHz9F2
1gMUoME/eIM18hFzHeSwVcFJYtMFnBbC2zEyZjotZepV8CFsKshZGtlvo9d61FFO
vbw04FSklTOLpIiMtzPCHNUUM6PEqOBbMMX7zIztH6rEolnZJAD40UOcvXhVHwpM
wWXe4H/iiKr+d7SXEYChClivIz4cVGzH/vqMKT/9UWj0Zut0M3lWLPIxrOvL+xg3
xG4ewCRwKo0MydcZTTMlwA+mEzSh7LCol0MqqGXQLyWaQAWnvMH4qNStbTXX4FSv
n8jKvfG9aRlQE1H70FAoQ1/wvtBJG5LPFbUA8L37REH5CnmhCRw7a6H8CK5Ccy1N
qD3WF/L6flUQuUgn0ijakYdLORsmbe7gbzgg/8/lOs3C+vo8/O56+Hd0mcUNhSF/
qHe5a1pcbpiJR9O0F/AphoSEHX3R3ecHjexvB7acjiBgAZuZrKsa3hnaQWgsPuH5
WKE2IEKoecyet9Gsrk4Zr3bkeDk+REJhZpUO+CtvuLwvyOQBdITIJiiisuSmLlg3
rSOtZqrd0PCQzgg1qihsyCY8WzxtUJtvheOiEwe92owLpi1FHWupFQ344HYWPdl+
Jc/W63aoTj24xbEdoSc4bDwMd7w46usMm0DxlggL7CQkXTeoYKxHttAoR6RZgiYq
pQVUWWW6IeSLqH3CI/jT++jX6TR079KMzy6+Z6y835/gi0kwi2FRLQu+XBLJ3FU7
YH+QQMEyPqMX6Wnsz+GZFVhHk3QB30vMlkgpnaOsSK3VZwt0JyId9ZTc2hlmRFMK
Y79WA0JlE/Jaikehfu2MkfXRLhri5x5Z0WCFOjjlJFcvmtFIgbsbafM/lsCIP/rC
WvxBRRpz7f7a9F/evYiemIK3arLu+WJo36E3prM0N0ciyxfnelQNxKWcf5L0ttO1
X2241F8LYCjl/lvThRfZS6NbH1+dmtNj4xVFIdO14vU9bP6uTJLe91gjGq8TXVQC
UYzeVsiKbulnpa6dLuViX8YZzt70TdCVExwG0HFiv7cdB1FFofEswdUgJGW1FcC7
0OjFC82BjupFe1xm793ssau1jGu4mu7wj3W5s6N3yrI9hQNht3BSR9zqyPfTV/r2
/w/kQxpo0XAF1IfNP48QwldIV2dtJ3o8jPFBp4hBHAgImC+YyYdRdFTAlmhca1lL
bTbISy1dkU6HQ1seFL8L+NnbI+yX4OWqpF+kHhOSh6AfJQ8nKhddP1yU0svN7fkO
PQlsIcDP14j4IOy21fmXUOUUUAlYVaHvkeVpWBazNrbGkE+AdrWAd9qlqrIb9gle
P1MgvYvQml4V/DcVfK2TS9WElfzirhFXNvAeBgLegB6Iqws+yHvTrT2VOs+fqTH9
yT+GLuUKBH8R6UoLMzJVRuWuQd5Khhf2x6JIQ4AG6+krXM6csXR5Zj8kl8Y/JDzh
bYKfuVU3wt/RaklWgOLL0e6rs1g0Qus/wWC9jYpggF9edKb8oEpttoxc0mtcffU2
NnDfuBjBuzq0FW6TBEcc7XhBZqTurJcB7i1/rBp6CpPkmg1IuSeM9cyD1ALI1eO3
ot2WY4iczqCxiEDIEJY4s+4MN5/f30eJ+IyAtO7H3JRTZk7hQoeMe+rhPJfWnNIQ
Erj79ou5lq6N2MWhl2VOuLEj0pD6lDyJ+5HxHeoN1LidhfSQyMEbbPrCitc2mKaE
m2h4YSqtxrDPjoOwA28ahvypTCgnYVaqKw9cVspoTWk5wXJllthXOKZHWh1FZbLy
ioqCJDFv55xgRnWSb05JbyUdhabA5iTg4z2YEXO7CTByIdrOatxXnqY+A5pbr0Oi
xXUfsG4h8AB012VTx6wWgJqMcREptcc/yd+8og1CbarEKtKSULoF0f+0yeNd+eOC
Ykql4miEzTL81UcJF9sjY0xNArZ25w77vHe+JrWldSaD0EIzs9vHbCzHJGjpPctX
Wn0qXb/NlPee0mlJLqDIimzcPN0d4KcJifeffE1bBKr1en8VPGvQXmWjubKK9hvk
nco2bQVQA1MwMyfpG4ww2NQ0AxDpUVletX5WxP5vzmfTTbfbJgNdGIVQ0myrmn5I
t29tZ9+ZiBThv/Ayd7Wnvd3HVqXHBAQCZ/dUBWVBrU2XtXK/ljLfzqVMoJswquRI
m4dtKZDHU533Qm2AEJ4o5Hva54DxAK2652yurbkLlgjmeCGxczYooGuAc2wfKNJP
APhdJVorWQ9pRHqQbHOrRBqgf5++jGfU/NedR+Ay9TWT1lXDV5C02Sl4wB/l3tK3
BPhZ5B4co7Rf5X8Qc6N56+dakMlfFwSnkiO0XHaLvuqQbpOMDaoTW9ueNJh76q8j
2UsMunFol5jvqY9HD0vP4HiNb0kivsLSQel0IAdHX3XUp5TogrYd5YTQlSVEt7En
ehmarV2Ig7P2SXAgPFiE0MquWkTaFmIJJNdQCG3acL43dFu8EPgC+TXIeDei1jjB
WJDr2U0dFwrFYp6jPOEP92YKzJzELpCQ2dCsFT2tO6u3FlwOQKfCOKyTTI7mleC/
bintMO8/3z7C+qhIEbfcr9HAnygoPzAbJWoOpTo0YVtgHKtx/GVRTs6WOqN+EbWV
RWetJ4Ia2Xrh9FrpP931KdJFy3ViX+OzE+i1pOJRPhd3XHNod/uRyesBwakPKst6
ygUdUBZgJev2Ve8lAuFo/vu6VorKs9x1SyAS/EJm5cs6ZG5t+B81UeEjWtA3DIlA
ttpvrZUoafvunaVFHFbznQo3xXtJka/oz0wDVFk5IvD0xQCIdJKmUlFf7uw172+r
9ANKfXMSeN22EF1t/NN66FrFCRKobEuEYNkRmKj+Xpi1ZbtBP3c6i0/JP9+dbgZa
098aIOYz6ms5IO+HgBIyDzBll9X1wGinCrWCVqts0bLu1dG8MHfcHdA/ORzPKz+h
RAGQMwcahbJTSY+f1BD2z+LnOgGxHqKK/WGewRc2KFrXB5gS81K4MFaUxhFfRUrv
IqV8r6yQAI4vh20vbuIHTLov3g1+liTbfFYA9kcpwW9RdgCfvN7eOMncmYvUsKqJ
RVVSO+EAshD4Bbtj02SjVc++oVxzRwH9r3pdYGOaC9eUET2WJ4auFwaVE47eEdGH
d6L/HxJsW9+f/MYIpLa3rKRRp7nq+yoXbTLifnd1WSL0DqmPRZAJ60Qu2Ymholgs
Y27r98yMfelfRVrm9/chK+fI7OtxO9dlieIq8Z7BizfYFaZG0i9uKAUClXbuReCO
L913dCgIPxzd/q3t3eP50CG3aLENjPKxVQ+z1qoi+xL6fh48MaFKGoVDi8IgJUcO
4DkGN0JYYg058H3tyBCOLuNFrPbgTKOSHWgVZkojGHwAweNHwFmM5yAXxKWAyb7J
9bS6HrCLOT9GASaLPJmKmHK+V6FC9SIHRbkeUvhwgjwY9EnoS4Tk3kUrGs4XoVKP
DFlNt5I5qPqX2jwDhLLzVv0L5ztjHkybsiO08pBLyjwwjBe7dV2oR5SLptcylxDA
D1hShKGkgZnw1wJhoQHVuvGZYYER40+WAO6qfq5avf+3p6yAXbxR75Wiq1t6OVwf
t04DsCCT37LiBl0YoFvp5ZVnONnHLY+NdkqT5QfWZKsQ02tm4QafeTwuHPibXe3L
CU0TNeBW33lDeZbX/AaSLI2QnlbaQTOQVrLS0iREOGE3EEnUzGhd3hOmlg1GbWfd
7Hf7qAoFrAVSqZrMgp1YGLX0u1vJ/bZt+x7pY9b6ySfUtWqTKki+hOxO+0m9R4pr
zq+Uh7kYLA0gPHhbPbLbvzcjJTWoHwcvay4wh5csPb18myQ/jet+9tyv5JDUNh8w
qVs8LC7HLpz7FdfemH2lUBIr+7fOkNnX3XsTJaXt0LUbKDdHZ4D/KfwuosIKMwMo
FLJh0UazW6umPEbdZMaNLNr4mlC65Limxp5CDAAL0o/Zh47pv1iGcHhT4Y6GZWe4
t5GQOlZWU001vANAQiUWKqGexLrJnzajnEioUqnr6W6WKoGKOBzFUUzzn1o2vLGt
h8c3aGueOr7hEvhMVA7mMRQCXwMQOwBsiSaiyvVM3RrF5KJASn2Q4DaX6rDFuneu
Wanj0XPh8dPgQ34QfEFb5nbQhAqcu1TRETqwuqTBAmTlOPJ/vtbYB19UhRhYsTl2
+Fqkhi38U+iptmuRi/QVIiQ4kdnY1Zg9aR0hS4IVXoOCVMP6uq+m8wPKpOyQKT7b
vDXSEtGIzmucRt8ut2kbCim3dh/MsYUZZ9tSC+uW9QrXhVaIsCsZae4U8baWHyZr
yATQjGUeK4EibqkyLmpU1MRLceTu4egDiNkMSsEaCqoq0f4k7ny1EKM9y1fazSKH
GoY3GXQfyDorcLDI2BO3tpgY5qKBF+A41MPkdFF25M0KjM25T1CR+YzNX5l/ULFj
JuEa4bBs93sKQb3he2a20gsqJS9cVyXRZ+DWSvNd4UcxOeBjVcX/X1UGOQQwOpwy
kFfEWi9t58FnhBceR4608HvPmvtC+BvHTYiuEGFRdL1Q4JlNN2ZGeQhz7LrQaI53
MC4PKNnyq/qp7IRCob1nsXgGRXVhix2ueXtuwmQu5UNaAn62e+A1Sc/ZKtWbb7YC
v2DBtGgoCM1KpPl9v6A0rNXVYHSgjjR4S7C0mUN6mTcai7+D8+lM08olr2Btp/Ra
N8psv3NdABkoCLdSf/MaI+JqPLNAnDqFK6G88TQUXA0H+wFxulbttLFPGIt0b61s
sl5vLVevni4AcKu89MTSC2hTbyR7NA3hrW+wxbAooGU7youK1nJ9cx8oGpQsijnU
Q5uimw3e6kdCLeFPFql4nXeLUsz91bYbf7mauLXnh317LhfiJFFgCAvsIeROKuZV
Wn1r9Sq1PbUxilUyhbi2td33c5zp00i8gP91mI+Tj1tmklanD0rofDhgV0+FO41n
spzpmkrAwYl0iDXctrU1umxXESoha7P+yZ9cxKPwiNDBJntNT/le3uWsloUr4prP
F4yz3PUDQ+xSQT49zisQKd4y2CRg3bSJZrPaABx0yx/zKX6HtnA+uQC7dWJoB8wk
OQ6zKlHiCQr+X8R/9MEMrpxf/PEXnnzCPdx/aVAlIeTXk/JDkzE8Q3Jl3AvFQB6c
NYYx329T+sCaUXl53myw8J1pNJ9GuFp2casyQF4JoZFc/55cAX/AGIJdMOwNhaRw
6y06xhZ7LgSKb3twkR1S63QQFsikSaWXObuxAP7+SCmek//sgQ6LWlaiz9FJ6rS8
IClZIez3MR8Rja+vRqwLrTbZgUFFigOlxy3mVDLSCpihupbUYM4I83+5bkk5/RLx
33atN0rBAnH1biTpP8cL7Etlo5Oi4HXdvTgOofcqVa7E0kPaOc9Pmc4kIu14hiLW
gdYiWGEL6jPIUp/p5PBDsyM0TFIvNI435+w4B8gfb3n3trFAXmr+bma5Qf+xpZWJ
czg1MYud37t1wQe+euEon30xVZ+6iQFZkBp+rglq/L1qrjxNKSYFbf0NmSGuODkn
MFzP+cen3/FTdXkZx6E9UtoK3JpuWEqQnqyxbIgmh3rjtsuOuJzGVMWs5EaJgrv4
otBppZB7JLDjsuA//vRcT63Ew83psNjaHhYcPe2pIXtQ3apl/b9J85DCpHqabmnf
L+OUW/gqHdcl+1G5vWykO+5yJnMBkAKvwCeO61rswBypaOuy/oanTF3V/iDAsFUL
r2KHGWQdQYqWdS/vykSp/DWmFHP7TDp0zIIoO34rP26re7s3xKvxNTeTnp7JzVlh
pEQBDQ79Dfc3dH+oYk1zd8m9grUzT/fkKu6Ie732Bhq3YLdp26OFk/VqjiNGpGib
vxxce0vQl7oIEU84cRIrdVMAh+WVOJQKN/fuQ31wr1tMD7IS4yZQUJAgIimO6GOu
zAtGiT8+hPIFrvA8pk3edii9dz36bwGJnNNaASBjPN0ZTMZNsKv6UQRwsmBHB+/A
BeltNBVPksIRSZkJnwSNNLpq4Asl+Y7VsYFLWWzNaWyZngvoRXfHxuXRmJDZX/pD
/JSw+z+X10K0D8kELQHaL87n6Q725WaARwFQccu4pVefcKFR4CesR3y3boAZQbfA
XddJoALbL2oFK96XhpZT0nodrJ5oE4XGUed+f9nFs61JwKgKXTeaFdHNmqV/mXbl
4T4Jt+plldzZDvMQFf140W1hMgnSOE1+h+/mOq+Q72X0L4bqQF8HCCUbHXEf/sug
GljG8NRDQ2fUuCT3ClDkkC0QyP+FuitbB71d5YMruGwRecytOf3bnd0W0vi4kPzp
+Gmh0DBY8Etdx9xvTMxUzl3t/OQBdZPNkBHowAJdAPDHHGvlokZtwNjRoBOC4/ep
VC46heGVhvyqapbE1/2ZpfVcvKJhUVJU5CMlLuaXOIQbP59wiQZ0xfQS2Q8WPvlc
XdhctmD/J1vYuxHbzrQU1UEhGyXdfDCcW3kC1t5ql0bAtZeFo98JDknNxf2RdF+Y
gGD/9k4DTv+Sapw+2U9vxk+s9Zak2TPGMddAqnf4qBQbUsfbcVkw+kqtKrJ50rzx
6a1CeLIe8VfiLxyfs0D1fpZDeuvy8FbXo4Zqo265K1+GjGtpCLBjy6XphZ1RUte0
mQhuM9qAM2r1H4Xzi4H2GIuC2nSbb5sh13P0lwW2CgTgNgZa79x2bW7YHtJF9cGN
MiZ6UiqXBYwvzDb4fBkoIk+jdJj6shhcFiqDj/GlbMKUIN3I6gYQmQTk0+AFEcdc
9QjfaXc/aHdSVcE4dMVeHOWuvkimm9R/9vesJy4jU0asYeEZdfVHKl9Pi3/KMuIa
B3CHS1Ri9SgMxXmhUZb4VyTj0Px2G98mrrs5fAK7JygftAJKL56DCCyP7gH8jpna
BbG5OkLt8xxN4rKOuc5Ck3bXXRilxSqaihyTLbEXrWrME9hefbryjv5o49STKs/1
cMminGUCfOLLdc9GUttBN4S2QDZBT23U86hCCh+41Da02lcsYgtsrJ+z1J0XhIHT
pv6eKJacRHJbwuVCzMndMAbgcnELAIS35hl1+jfE+ZYYNvBRZgvS4wJS5eQRO8Gr
APQZmMGWGNue3wtlg1fRoLtUdA0SsgP4CPBex7FYyQN/he+PHcyK3bmijqfn9AC7
UgfANcfEHqT/Z6mnDxjkasfIQqqzIlSiyGUPdgNijxXq4HjYeVvZBdBOTCJTOjfy
schycm5O9w+ZKxE1avnMItNt4AqFCMfokS62SNxHaG/F1ikA6IUOLgKuqSDrWQRE
yOZ6gzx5nMuRSKrbyAe5pUn47lu6AIWJ9wn/Soj9HIGCz0+DIjZPTh3c120gyXo/
nbTMRnCzVbeHx2wB1ypP6f/0KNPKapzYCUCaHt0DuMPEsRIHU8bOt7SpiMZujl2R
DqQUKt1SzWGs++5VoqcZz5lewvn3OkhT1atcV/2+05m6hWO9j+Y1oQijSUasVWQi
L41YsUXBeKbkqKaX1SoYJ/+CDL2Mp0J2FLWl9Vu+CqVS1MbIoZ+MQ0dWxKt5yM4u
RRe2K8W0oY4B5i/ZsoMhJRJVhX++ZXda6PxgrVquKBvIPBUsF2AQHpik3mthOjFm
QuoLsdYbcdZy83dmkKKXoKWxWJPnVcMBH9bV3XrJLNjQcc4XyCIa+NcaL4YV2lW1
7vJeKGCfl4VdN8uasyDyG/RiLcH3cUZzidoKwD/g06yHaHH1ISIOi0s7KCzvAjK/
WyyFmULm/EYVgexowXXWimeUcS/SQQmh7sPG+by/FKsN+EduaMgIu1oXkI2CBhp7
R1zW4LUWyJSs5+mxdbtPt7ohWcW/y+7aicUJ/WwE4GV5YiDz3+Fw5HidwXADdX8d
p4Sptq49lO4568Q0xiRZ7Ar99twBbN0eZWczKTCwCJQfiRYjJisIZ8TLiN2/KYe+
7ov0oJkG3DdmrC7LQ/fhFQWhwKk3d8PrL5r7S0Y1j//ljY52gSd4IiJmtVokWQin
LvBKztJaKhKRPZV3KsoCGyNpt+QLWH/GlB1izlP+jZqtoQPlccRFg4nOpxjjj29j
1T9J3xm2XxN1H+dx8aQwnWku56uEuSPGPs+KYKhmgOFK3toPBBmZLv44O6GxRW9E
ica1xD9ESZr1j5DefTWok/JhqjTiMzIGKiVKK2AC4ezHkeebuxyeYu/kTyrxRWfO
34EZaeqUzdDxJsQ7IPLqVtcsgWVf8JHK80NjluLLfAJqZuvvi4AvSUkbZTZhrSGX
Ho2wVW9eTFp8eJjXTyHdck2aRFB+918vxkFEVaAQiL2FFSUPq+f9rAsgJb5ypzzU
n1RE+twlZfJTClFQLeF2O18GryxYZAcg5lDhAwcytgqTZEF8X6xQLlMIsKdB3GL1
oVaDUod7ZsyrUN/LKvlLTS+fXfGkcTJg823cChyOgyqT1sG608rdMXoqrPqwqsJk
tzReWEPGUwEJ//Mhxg5xPZOTf5CemwQ7hxb1vXAO974qDMdKEStXiG2pmUdmaXyR
F24ibXu7NG1yHzTFQ7S0BphPIPMeGbah2T2saQ33QZ0q6xbR7fAOSwfV0kH2mZls
9la6gYoOds+4XuuFhE/gUn3mfBMtQrMbdlnxsgTMmxqGljQG4Nanyup9YzOPB2hC
r5wT6t2wHcVWrUx5TSSVB6btCbg++Rh58KDFEhc4YC7i7RzDK//Yyl/T9w6zVhHw
q75JNrjvx76LybnALhNKOkx31WCTP5WqA0xkqRZx/0IcoTp7sZX/EElr1jRBrDOh
MkSxRzbFTsY9gAJdkbmH3JQ0bVJCyewvXgKb1i9eMMrltJZyUlRzrKZCHtc3W/Tb
wQQjtksxF2aj9fzgeFpiacwLxEzZqM3a0XYFwxAE6i8iGZlFmRFw4OCkQzPlnaQP
jaWK1txoNMMCA+s9lLKvteAJJbIdRiDRXv98j1qOb+ifNj5HmKOl0VP0U+f2tE5d
edriVU7+Qz3TNGUeiXBAL6lbkCb0yuAe2XC4+mEsmpRruPuYfwRX44cneN8P7M1c
ZznWzdAMciN7NOT0cF4SCuEeuMLej67D0FyaUY5T7qVxanlQUjFLGugYtMEJeHCI
YXVyYgIMCqgpRfZDtCU1rvBll/gt5QQTCuJVsVuYVL4TQGo5yMxxwXx6tiwT5mC0
5IZ7oKHhr+x/5DFR9w0SkMkMgh6/GwdPeh4K5bJT5ZFd5NeFWpzFmSVkLfX94v1T
skp/wrAeYagaj9eHT8O8ezqEbFcNtn+pg6qx5Ozfx/cx+kA0/Yyw6dRnKd6bkA3P
ypNY5QoZkgw9z+isyIq+i9uiwIkQvJ+Ib9EjwOIW7Bu4qhTehejE0erOuPbe9uIN
ok0OKKZ3eDUCH3igKbRfAW0i6WLLOL/J3vKs+N+PjE3bF7Mwjyd8ds/JboxhMnja
vgbuc+xLFy05G4KP3Q5NUoGNyaDAN3BIFruiLqx/Q/cXby4a+7iMtQtzijeK8Jkg
uRRyB+CPFOjOot2PCX46F9953HzQMcNWKSLhaHQqj6i6ut0yyIVqybsXUk+RGOof
DYe+L0X+raKZAudle8HBXj5Q9D7EEll67BFmAEKAumUJ3qcfFcc6/G6Rc0bMxz4p
Sw5+sHV3RjXgc9hf0LbwceJ/MU8WisyFWy7T50Ka2YhC/QQX4ekjMf0wz8M5opaj
6rRKyf4C2C1nCYUqDNG3+NYksSWd0HR2V/HonjZnXZ3ozNQ/DUKXYDgf7WM1kIcs
1rjEOs8qZHoQ44d9C48v1vw10GHbqKK84hw/4Lh143AhG9BgLpD775+Wp+biEqOK
ddus/cZVXCUrommI3ya/X85woFI92hQkwmgfqCAHfenb9Ho3i+2SGYaT6CTM7r/u
+FFQ7z9X4mYX8wmPSlu7lPWpQkBZ8S0rHDiq1WRaGrOorceVJ5isxPR943WPfvsd
3qa5wqzWGjqh0NeHs8iFTg6JlygMaRuUYbjvmk0GRfTEo12tW8vSEK7hmSQwGS/m
88zRerG3tMoEMSzIX1cMihiNQeb0WtLTedxmR0crTWOTny5hVm/bL3SiasLVC1S4
bTMbl4Qmw1L3IUpBfdYUjxlA4qnTAEfKSaaj9mxjYjwJvPerBUCsT+F9LjcejgO1
JLKEksDYzK1172A5jBfbvYWi0hF//4uRjZv1TkUv8ftp/QeYbOfbRlvAmLbp+U6Q
s/RHATxFoUFPamqOL57Es+TSckHkh2406+gw0q4UJEyT5igMMi6Er1V9lcqBLNS+
VzTl+3Uw3EH0r14OYJkHqr+h6Xiw0yf131YihzGYFECb9C3IiN16tUjKUOKo2plD
jj86kRr58DbvkrYVR9aoHT8DeOE+Ct4HQFuhMYhBmzFNdjlsZr3iPZQrpVJ756RZ
HCuzgNpwp5JuAh39ViBd9KLiwGsydUFUzKya0xpJguJ6gcU4Cvc+hjxeHQD0rxdn
Im6LUqGopBY1LXwe1J3yky9CDgA+stuIi8C28LYrauoDD1tbR6LvKPVAIDHqjpwM
3F1N3OjsxieEJLRwLmbsZDh1IEpKG1uGkFzmARZzZwcAciNyCS6fUUom71JocOj1
ivJJkw2+pb6yyQjj9QgP5qFF+HGULXFhT2DlDUSA9IdHXJqWuzg5TyaNZ3KbDprU
7d7xh1etA8MKefi8vkgqY2HweOpix3HFP8QWzMUXPbS/WVelYXhvLa9nBjo1Xgn6
qoOvEVVbwWn1Px+0vnAR1jKHvMheKAA7BEDNqt19zm3az/BHZdYj58dw75m9bFuo
AcvE1p5/apzb8VYoXOqKueqL6WgV69Ar5g7ocRAacWBX84mJvcGbpysIJoo7k1Rw
LF7LfrgBKDEzuA7by4X2I58+2gxgqIV032hH44QRBq0p6IJ9qNscy0Mf6RKBk7xc
TLicR4Ri3urcRfWvOEZkjsALP5Q1ov7fTR4bSgVXKtqIzXWbyMPqBw/HfH6k5Vs4
FgvV7ZeXnFUjXbNU+dlt6O7OOeobvuYokdyNmFUvuzYxvkMzoCiU2j6j7YY62vZK
GTwkMTYnp2foWtidFLxFWpzRs6NkjPaaBTRLlmuFm4m382fg0dUL9tqhR6uJCun/
XxPxrkmRnDiO06Ixhiqt5c9xQM7i3++74tHEZVc315g2tGcnM6jKli60M2YtKPOh
hh0ZR+0cTwgH52WSacuAVdhPKg2Bo35r4sIJcZDjmbZbky8DsG5D8GCuxPe0/S2o
6NJj1l9CSrd98MCn7Yq+gYrxqxsVgl+6HSO/Y632OA7Akn+ZRZafSWoP14yKoADv
j3RhCfSGsSWr+tgrnyvMW0xxuXI5hNLhpThyB/nfObJcij9ftPb93GapDmdmnINU
ltnegKl1yo9+LgcLwmWaBdgnrPlJcyeMF+5OtU3SM3aQCbMLMSgBSMSoOyrG/btx
zDSzQjvXLnWYNWX/OZE+qcaX20ZYmS0bXik1Nus7O69VrYg3jSpr4s20UfvoJIMM
42CYbTVv9T1Q9TvjgwykAbbyj1cfPr7Nu7aOeG2C/zxksSeekArxlxqKLl0pDJAH
XlEp7T6RJLZjx6wyHiV+UOhRpiu7bmt37qgre2l5ABG4YIIc9oebsqzmPCFpoTyr
L1f/9CpeqiSpY03GaCaZCaTpOTXVFpEOcdJINRNZBNYHhXBZylJxlf/0U6Z/v06j
lDOqaM1JU5+UnbxqOML2Bj5HyHtMrh4jOT7huO8ejnCX4uTJ0dAUoMTUR7Rmth9d
/jxTu8+nPW4M6hh9gyg9rI26EryPrYMGo89nHGlWN98Q2ZfO0Gt2YjrXUZddbp+E
Cug/UXg0HFY1AFw9PjN496GPgXX68HISNqxyxIZqddrvw/hn20I7tEramq8ajiKN
mQYifHt2/SxHFCfLTSHVbduVtjdCyU/J0Sbz7A+63IJMEjsuKhf27AF2e7ED55MQ
U/FuYMMF0k3it1XhzNQry6hC/6ApnC4gBBB6DZc8w6N1vULQr1tPBGosDhEakmKQ
x6wcslF2A/B0I1qaKOrgJeESEPukGu9d4gYNEidIw2dHw9mMBsrz1ZqrrX3lLysA
aEusXBTKDvxYhDSP2uqzQuPJjsgvX/GKcBO5GADJgwN+yoEL3AFZZX07Nd0ikEr5
bZAUQuPgYJYFJ7uckvgj1lE+wZWU5webKhi6m+v2AHzCyNwvWgP1wzRnFo8WmSss
m2u5zd3vjjkI/8ecnKW0qvQVjlklREKS32Q87iRBG9OhnmS7hwhaLza6AhIrCQJf
ECk8ekihSpy6sb+AS/SYPUcp595rHZ0gSVtT33lcZhbPw3dulPJuoX6X0Kl0y2Ez
/T3mmubTP7IooEssM9rVlKdVgGQXOPMvn1WTxCJp6k9BODVI0fn8VzzHFKhQYpmS
ZQRNU0uJqJmvQJExQa64l3K/hC6yK776+8oYto7hye+UVYUXQuDPx3Qi35TWQ1aj
BJt6a/YpUZn8aGMYcXI6NgyefWqIXBmZBgscSnC278RsDfUSy2vFf+sJzenyCp4g
86TVc+wQpe73e/oe0qBkZyXXKk1/+NeFD7SsXt4M6KSl555gGKEPBX6NipRkIC2k
If64swbXt5Sc6RTlfu8wauH8lFxAuv29sGXJrnCka4m8bq3t/eqVaYCPXi1rIASO
4B6mGtpXa+ngsEx4j2gE/XFLIdz9dzWdH6lpI8+eAsBUidP3M6A3RVl7ZuPWF9XN
Uj2ONhW7Ek3yiKb9pVIqhwfKsGHSOUrsWCisEGI+GFDEf9dpCqc2oOjMzVizGwRI
RgxF+SC78z7GH/CqU4wGN5vKM2sXCSIiByDCjrBNxSYF5uvT3/Xi2jfWFE1rEtNB
MQZwrcxjRuPrB/vAOmnNl2sQcU/e0Ta7wruHw2wB77dmu/HMCbNmgYJghzZKSNwd
gxQKEptU/MDMGR7jKquWVOpKUB0Za3x7xL4nwuT5m+jCvtudjuLbwFwKGvS582RW
bnUhQ/uhWijLm8e8vwDpu5htiCVL1MhiUyAiasijahH3Sy+uyrAukjrTdiXemY3w
PTLT7mc+mTpR7TFTF1TRf+P26t+9vZg7CRrj989cZTrZlLJynKLfMHhDcV3hBXrB
HGKKZOIivtb4TuATtVWu531WFfiMKqyuIxzffEP7U+qKkyOghXru0Le8U+wJ3esI
lAfTMvDHuIjqdG5XHMOytdOAYHlvLADTMABY1/05ioINjMBcDdAXK6Slc6aMn1/T
VeIdpFYUUzKaG7vjxSyMxu9CqTw+d7wnsbHpT7rEykGEeVrfk/AFEGE2Mu33tkun
vUq7OtPmVkkxmJoyziSWBLMYY5ILStgscLHKYnF5A4UtQIfIqgqPnSp/iF62e58f
ls3BAWIW85PIrJBVvMHClyt0IWSKQOkGjqrMjKip1UcKyknFWGMcc27gY4RyCcNM
vjrMERB1b90YCxogKJkCHMjdLoiKFTE3vEZ2f4gWQEr9H6zucBGrDHrHz7Zw1A2A
RQCV5vD+tbKj2jz8AvVD3vJHe4UDtHQDH9Q1Wd5xg70ahY6lEIGip/RvEPOEY0C5
6re2oBWfDsb9y918KlLEY/yMLJzGVJ4b/Put1jw+c2Kwe0K2lncObxxNwQX9Q4mU
2zBdk/e9Pc9Q61x+T7OR/vkTidgSJGFO2A+gBQSkv+xgRJ6jTyLvE6ui2hE/81ue
vi2E7xM9xMkv11P4slQmqS34soJK+r3qDUqj2vExOng94s8PMVlK2jzZvHcPZrtg
hPhJiVty5ZVxYiZIMzqIz2BdGTIOXhvYmEjuy8Oo35UgHxhoWXf2yX+Ns8DxR7o/
mxmwNoIRyxPe21apNArMFszkHUMAU8VNzusVxaWNddOdrqfLi7VriP+Y4EJPdA4v
h7E/DtiIDDsRk8ZU8TpbxMy5aKDEHj74I7bzgIcnDwOkBEDtSSJ/lGnlEY473HNG
gAH9T3cNSPCW2Z7lK/ZZLlsMibufNZu9mbtiZxvUkrXskmvEDDR6HHbJYNB1RwdN
L78T4jgoMYmk49Xm7admczse8TnRaT2aPyQOqRXGjQjPvKvDgtMeuml/o1DJh3JQ
fSY+9clz88XkYp4ZBAS+DoKBdRRbXCC6SiAa3vJXFB4PJMun5czHunPnQTorXNmH
TNqz3aOecxwM6K9vl7xOJNmyJMVWpVdfkLAbxCmLfzouT6AdU8r8U0oofvQzLPr3
aiBJNouU+KfqPTwErgbQRHkypkkO2KgJl0PP4D4npiiF3Qj/BB7z1xm/m0D9qhKh
XAsB/i7mVf7W0wM9csBeFxleg9xTM3MQ/PTNjz/yUf6hjbspjd+gpB5A+XWFuEzK
h8+IR2X1AHO8YRB0yLQ6j+YFKW3D+91ma/A59StChUGuiVKGhDND5LoEiReV6ZFh
fGASBNS5hOTN5PZAvToqvgsZBeNruyrZjhlSh+MW9KZyeaJ9xlpY17KzB5vvRZ7/
ou4jL3USaO1Wwt3mirQJzR2b3elHYvP+tOQ8znKTbH6qVag0fNfVTZx4tdcVFI/r
nxkYOXe40E45tdm9Zem372JnsQu2FcmaqHkk1bWv5xWqe0RneFUO1SCt9CZ24fYI
d5q7QgWHNs9oxEGD7Hz1dbw/zfj7LWzJqAcq3iOV2uOff3UoZaEUzSUz6OuZ6BNy
VXpvrR0BMrSE+JTEvNcihB8xDJyifFwJ7HzuNhdlgKaKm8GGGqjoL+zQUvvM/CwT
eqBRuDOZkDahQej9fNivqb2FpEA6fk+2V8yQvG3t+yt9ZGhTJkJ0w6et5k2MVHe/
lWfFNmZmEblRpAofNdDHgd70juJ52qDi27AwGyYH9BrxLOXYQKAzq8oatOjZqU38
bahp1GgsrgD/cKKFqlitJk1VqkImDJmyyoQ0SuvAlPEckWsT4lsPkmPVxRj6zm78
RSBqpm267g+smaOCL7O1l7aOsoa4eiYS20ETVCJLGxH/PBDbcw092DcI/QeWEIwt
iJWAbizDafqr+NvbhzOtWmYRXygWd3i5yvaTG2tqwoQJ/3D3AAhjdA3HxW8zBdjR
fa5j9iIkJBHAjsUFEefO3i08GZ/EVexaT8nfucF1C6q2+lW8DPVl1tVHNrTwP+Mu
ZTKMYoZCIc2S16E3ErymRhXXsPZ4tN0IhPntrBdvNwLVTS/53+Zyd/0MWzms2ZCp
RTNgf6NcBUOfKMwgo+b73fgC0Qo10kKRFJThDKEkcO74B2WVQOegO3gVaec73WGd
InwQkif+k4brpXr9PZqCbaIhO4kEdQHXoNg6JgIKUPtIx/RXxLlumOD7O/LiACG/
/laUviEEGcpP+Kk5uPx4khombe7ccY7gP8zG5jcyXW8u65eO9hxpqxshLeMqk3Gp
Ccu1Hp7RqmCna9LaNWIakFaF1x3JlnT1XPatriZdk7oxUNyejgNs+m7joIwIO4U4
UdB+sV+qpEqH+1bwO9nGYSucYJLaPkuuY5im2LSUxdqhoaT3PSXIl4RA6ahZ2zbY
iHTQswf9Bg1V1OHDszU9uRTJKw94mLrV+edsmMdMocs8GO3zVndtYrpRUDLnu8SO
bb4F6GSx8ygMrkjQIjGGP5kuuJOKDH2h7ERiCfjgQkjLzu7NiUeUCSEVAvgoMsC/
Khkx+Eo+HaWtade8dxcQhqfVC6axAFLWeu8RX+iPwYOcItCw3BuhLNkLjH3NqIa1
nZi3IDH7JJ33nLvDf1LuLGeDHDBN5PQFnmU/2N3Wres0lg1cRArNNqcb078XkY6u
Qjn56z1SUy80SRoHu0+eVHBsmPeTULLBbLBBeYRQWX72y1OgjTJuqm8vMwTeZA0x
baVtSsrF0uHf3H8k/0jl9GIiUYpmZrF5+g7+1dPYdKNlrqa6aiOHU6xsxq4nJ0aN
1SaHhGSCFZ/6/TLblovppYg0mWV/Qm207hS3d8pHAWq6i+8p0ui3gx3Pg4JDKuYM
ptqsRTB1hSQlHiOIKbaxHZNm42/ns3Oj4C6UXF91iaQmOqZGUWeKqmV0H3M5l8ff
B9U73MyBvQimDe0mH22NTQHdniOtA3kETDVXK4Du/67VeUsE2sgpq5koY8OhjDUj
HUURDQ0sFsscLy43pOZO04zKP13frkyWAhzRjyujoDErLzYA3A+mtEtz9A/kfK/o
SuXCLPhYPB73MqPVv17Fpy6qiwVLmzT+3PPHRDlQKKOi+x0evge/dba8iCpQ9aar
pzAbu3avSPuAjuYLMhwoS98oij9JSrdjQ8Ht2TtbwmYjmxIrZaUn7eM8YdG+BgWP
1OdKiqVy2DdIYv71hev9Z656f62x8GgqY5SkgkI4ayU+jUGVwqraVf1Zyrw2Ekbj
Zu+f0CcYuk1JYykUNErSGn9Oaeoi7Tg8c4KH8ouktoXOcehiD8UwRDZLK4UULbZJ
o5fthlC6RebF2zrjk/MQkIyfD/7CcLOOx+Badly3ge3IkCmePJNXUVTuviUNvff7
mrHjVl37sW/MH5xkSH6LVe4vcxDQMB6jKKqTbi0OokozObtfBSvvC7ld5g/hcIFG
/EXaSO5DJsLFJYZ6MST0JRpm6lw/YvMDJTratx3hpfDf5JMz8Ev3Fm/gwdpJyJsP
W5KpXTPymToBagQGGd5fd8F75rT8nhEgY2RTAfTx+Hs8bFVvRjVe1FniDjgSC+FA
1ro3u3ipIez/i2Pp8Tn9N+ssxFx890c8Llm1w8tnMRTf6sdpAyV0NbqqoCp+cykw
vThekELyQkZlq0nV0YB+JkR3aqcW05RaI3R16hozP96cVWWs3KJaLdzcT0j4x2+V
CJazPkZ5WqLHQgH8Ldx0IOk2tJ10tF/vKPnPk3hXmsVVCqc9K2RRUtzgm06ZEhAZ
q6ijhNTHZkaG+kcCuIqohWfUfO8Wlv/iNp7DZlU9Q3gsebYMNI4z6QS2RzDS6W8D
2eR2WFehaM8Swv/qXR1tINd6U2EHjWu9goWe9wCF6RX/cSN8vk9rKxhRYyPG/tw9
gSh3Y7alpBU5RZ3tFLLs5Fzd/IzpE8txzHINmDn3fKuEZh74NxRilN7TvQwnu8P5
BvPyRtu1HYvn/l5p1+FcZ/EjXdYWkJmkYkqXGDmKb/i/ICANLUo8h+MdQ4RdluP1
rLC0X8PhHQDFGUqXFqsgSrhGqmzlaPtjAU/RG/jyNoBvvlX4c1KXs4Yjqf1Mo2q+
K3HZI7uqN3XUZ39Bd7YPNLcOPUvfFLIDs2+atX98SAN4rXqqBAfhIXMi/HD09rLB
QS06U4DbYhpLSJt3zslCV3HjXS8CVM5Uk4Ae7P6bHLCYY7flsOUJ0qp8/uH3z8xX
A4ehOEt6o8mQnDXUTkd63DJqsadMT76Jz8E+KinimLYqEfr/P/favCOr9ej/vHzQ
Y58lfayeCQZ9aPFEF1ID5ruH/EDiKCMsD5gDmJizU/ZH8lnV3t4VTgC7cFA82+O5
K3l4vIKsx8bjCKr6ZkO1Pq7PzbZ6rZoW8kUpeBO+RYCjSRPQpQYZnNeL/aMrOpDc
dOoIT+2a+pkOsDGmpKSKRtwdyXlBU36VIB46iwMTlKKSZ/5e4arQJGPFCoZIkVwY
Dp2yUws4fSLf6U17sx0KF1X+rpZgMG6R4YJ/XVQKzf3Qz1tOh46n/tpxaf1eKrmv
AAxUTqdGV3aqYLF8PU41UQutZgG+6565cs1HFAVMSn609ndaAGfctFSiRR33u/Kz
PlWzSniBnZ2oHzClI78Ewc/RUxVu7TA+4ogrdbKgduUpzy9hREnpTgAh+G4fJTCN
9d8MX71LZCbWK4IwFqOB7LDe9eWK+fLKTmQYnmmGhg8Ow1Zw1F5ByY1Kd9tEPepX
FISJQlKP6bWCu4Ine/6BzZC2al4U7ZYAq/yL9LCLUSQO88dmEpbQSL/SwZa4cCfl
MTQIwIXhsfsNc8gAGJKq6Qjjj2W2sRUj2lxC9eho9OJsP2h7ShohLkWpIDPfh8sw
yL6+20f26wpM1JGV2dwI8qwgqX8xhBHeP+KBN7afi9Cmc1mvTpxPuhmXQztceLna
B0mzd6tTU5ZZAaShSkfbKpK8xGCOfgjoXXlf3meNBsj+0G2dHl7Xea7xK44pbJs1
xFSD0RUSFZ0/UDm/2kb22V+ci0uIkIKQ/qC+3iKYLYV8u3vB3fVhDDIdTmR2XlfK
c+7coxG1PFK1WkqduQca453wnTVUhE+B7X9ru2OK/0z3V/SBAeI18igszj8E/LBb
LvOJl7bfHa8FKQNCnA6eZPLwZmPF+g7/vSHWXNX4m4LfB33hdzU/F7qJcqlO1upN
eI7mSywdLtC8EeRuPLbe0dz0/p/ZtmUz9BVEyl3SXw9Owzws190+npsOvftRMb1a
hYxKFCsI66SxAD6QFrMBsRs4AeGX+SPQaQjCL6WImLGK+ykdsI5jv3gg2L1luj6Z
kvX+E6d1TzDyXtrUBUvXj/yqKUA+oKaTN5HT9jwGxyMjNDUqufQ+4VbYLGA0oiks
zNTQ/db2VgTFl41i+57dGilC3N626QMSlinaKyyfzla1ekY5TeCU9opfaVJfeOHg
PEE5BCsBmQk5fcYuzWdNd0AqJlYFLqtxpVhr1VjXOFcoCJv71Ri/Xmhu5ubp5m/8
EISU89RyXmbG93ItmPWvg0cxO9bPZgKewK+lIr26XtgHaTLGv0AjBtZwvjJxWju3
Omt2mEdw/YVRQ/PXFYJs/xI8iXgBDWYDc+mbNF90bJL0OYMIC2qDznKdZQ8Jrk4Y
zsEvS8H2AkvrhqxQWiO1zswPEiDeNaaRQJK24oZg/XymgCAnVzCJlMoMdyJJz7yt
lhRsYjmNL3EXFT9lAeb6uMo0n9I06w/eI4kd/tV4JGV1j3p63LVYPjzOKq9roXdf
awMLGSwHZrN8lhg4MK5vUzxrMmZklaDW01o0IiysxHpLI/ZxRQ5lRlwoCxWN0D7q
htkJH9voK4avx6l0mxUgKcjWHhKreyNxddXn+P8YWzwCm8fozNvIWX7ZNGP4IBoJ
eaBkYj18NyZzxwJD//0rGhf16GYaGGxZLR8aEou5EsF56sgo4x4037CG7DuigsSB
txEZXskHdKcW2H5yDcb8Kz1XXcmnU5n6dRGR2F2nNBNX6on3XDO2ldOECqUPXeal
/0TjmrVXG3GCVZ8MciJRQSfU7+Hz+19u4MDLyZjDxUPDmwnx1Uu9l0J3e5ceiIaq
CWY5uqrZOiWl+6QqSmGppz4Bj9NCsTUM+6OJINjHSNl1dYGEM7mZHG3P1Oul0D5v
RhqQUpv7SyYuX1LDrVVzJOcdqIHlVmwBXjhTn+JxyrIHR3VUR6oxG0iRg1ImpgLs
s24C5s9zbH0pS4fow06vOabLGAv4ll/XawmZUsC0P+1vl5nIpd70YgvVYWsDSF8X
fYapsitUVN+on3Kjbbdo71IhLWM4R16hSRR+3i31fM+6uLZyfV/s1uvrfdfCeKgc
Q5v64yeYoDUhhl7MYA7gS3zsZWubgl/uWmjPoEDw2YA77CQIcPo5w4Js7FZJsn+b
/4LGmKGabyS0VlUcZOi7aXTlZWUKv6oJZ2z+4XhGJceLiqUpfo/24BdkeaFwqoP7
ZRrOjN3OpSKjf3UEE6O40mi2ECy3n6ehSE7RiU/VZBvFL6AAYM42krZQmuT9ickx
nq+t8PW/7fQi8Goh5uaLfcbPRKEMbVPSFtIo8wpnFk4O7Jp8jK4EbOTwew4I0p6M
JmOen6p7cyb69A4T+xTZNq9mva+qrtHhELJQq/j2CLIs1ayugFmGsvO/oJ72v41h
q4NuqRkVjQHlHuOPv7YLjw/aKdCKw1S0EvM5fazlQr6RM02f2k6l24U1LAB+lcKO
856PnmLZf7ASnYlvXl0c95Yaz8a8C6cEGhxJ9Ec9/QocI7J43RYPyfnKLEeajHEv
u2+Bcipb98zkBr4+tIat5K4MRYvY9/VbgvpPBcuYK/xSLA8jQGfSMlCpRxLaXukX
IELAalp0UKlnGQf1o9nqNliyG9vN4uz/RSqPCyfXT9sx3FTg151AkbswTcz/hyg7
+fSt7BoAdpCxjKIfhLhW+QyK/5w92qMw1YtM3ImO5kFOWwVqIRsP3V0YDStEbwxl
mAu8P9BmdfyUHNokbrYlS62BdUZDVP25viaS7GeOC/u7W3++TiVUODPkvKd+5KST
GeZnQdW+qWr038trj29GogLwrFxSwH3uEKgl+fpAi65+zGxnN5agZwYbTICRJ0cD
09dnFCzVRUwYl18lhlrcdPkEGCabL69hgzPEIqTS+1Nnxw4/Hhcug/gKcKnGQq89
Au9gGQWVJfs4Oi3cwCICU7HJKUnrDW3Ua17Hh+f/yf1y9ZLpaTiNRh0kTISiOgA+
CrTIgoaSzCe1aq2s99CExe8MKK2cVp6q+0j5JYTVvDV41A0iyJnzfHmbeAXNNv9e
QWPodaW2E+EMQfqteaNzMddkjvW/Zz2F+qRMftUCAgN2IAR4kjEFoTqSeeg7zLam
M03eaYDkQbr7ykm2HXjRCh6f35d629kSZAsTCdF8jmZHb6753ySsXLOVswSEMllU
JzeNVyVKg0MeRPS7GZUbndvlBa6ZFZ8ghiqJ3K8Ut+LiIjgfGOGZxcU1Pw7kG2zA
miLNrcHK2h+2CK6m/nemn9Au6BSZkUzqFCeZnJNMRi8X02UR/MqB9ZlDCBBZiYrD
866UoaSgeL6dlU0Ai6wVscdIAp46YfT3knQVLz3TXsdU2VaeNujMfThBKeeAvvVf
t89X+Iy47ivQMeIX0/91b1ifmGTxT6m2adNQEp9hzvwyFTtTHowNKhOfhdX1prOi
jywpJIkFhZPgQ9x2/CtU0tvSJ5J3p14HZyC6oW+1IJx4oTp3+G1UgUJk5xTGnUZS
VmrsIpMGN4yc3tmyQc+wLMMSoIWbBLRF0FnfNFaHZ0rY6lmOOJion1Wdt0AdrcjP
em25Jbqs28m/dceMWXXDXzotHIZTK2OG8wCSIz7y2cnzWQEqaBOp2Ku3axciQhk+
rJPiznN5mTU6w3glLKslDzljfjVID42eVlVdsx4/Kff/gO8v5bXtglE2j/KEIXQB
D6UGio3kFV5nfCs6250witQRbUHAJb4ZRMG/5PIPngKzIAD1x6/932Hrqtnbsv9e
vuHiZXZFv9O0gXjgMnAQu7VM07GbcELAldtUkN9XQXCVhNItzPKAq8zz7sBb9NaG
oBpllhkdXNv/U77ZPRG+V2cVorPkaBAN6yTQnwMl9mlRB8d6UZEXlO11PUG5VJvi
oHmzBDCgvCxyJB9PpkkXs3bIJbPbNGEWUHR5Q62IyAnNfeUH4EDx3b29Xem603py
iw6ed17rxuFo6j9dSLWOUfECwDnOV3QR0nqwjnR4PceDz1Bd99Qs2tKMlMktcUPQ
VSWejJPC5kYDAkT6wbm2RMI2BN8XgPYxKDdCxFSCwq+ZDCiEcc8zaIHnzm5fY7I2
O9sqxdbOvd3q4g8Y0N845E+GNGpg7DITDrwmQvq4vdCtDH8ZXVUG5mx8+QAzPebB
q4CMBXjW/fcUKkLxkhsrE4ghYOcc+AzuY8MX947cI+l7IvoICvwGRvtNpmRg3QTr
SnONgtqiEArv7tMXfe4R8hNBL1dbeYTd+taigrZ3LGA0Wf4eTVuPK73ruuJT1zIv
fvSWp8N0EjOGnn9oVJ4Grf2i1wxG+woZEarRq75RQL8CFtVYa+wz/VGecGmBC+R8
xisbFbRa122aAQabQMNQ20ypgxp+XfkmrrNtajj+VVctAqKFe5KhWgfVxHUwvSYD
SWoB3Tmak92JFT3UN5ECHC/vLJv/NZ9ryyAWclHYbEoe/JzmpY5wzsr7JisVPzj7
27FIP89G8/yAMgixluS2Ai0HK2c1XkKOoRrspumav+BJExheT1k16uH/29jF20wc
oFHoOFormCc8kFdlUM8/egnR3zYzzuVX1XnE8f/0YizMEWGop8J5x3EzlNH6S4Er
U3i6Qz4VmMW3iep+VytwH5SBKFSeFmpJm9lrHKjjkGufCE90Ti2PeLrKR7YlkOAd
MweKv6I68kx1YUmjCc9VokhVNfLQRIapuBT5Hwv1kGml7ke8nbhCPxlxScZuPJhe
xz9Lf9LN4D0OMT0GZx9RNlburBNWb9AYCrzFk343lxQ66QSdVWoWGMA7+O406aB/
f+TEjyVyuoITBtIvPHYG6CoFyxHjOhC+FZ1Nx5cpCMsy4lWus5NrV5UgAsMv4qgr
a6WCmqTZD7NmE80gUtNJc2nKbjkSmLcLd095bazkfFMJIQpzxPSmgI1OMpCzowKH
j50vdamVXEePzyZn1H16kDG/ZHK1+ilpoakbi4wLQLEEo5faWZaQfQP8DSpMLkxq
T41r4cgo4N4YkT5HlPyYkMN9sau6KYlt1ALtaSma299wUGwUaPA5NbiA9jgt8/gP
yP8lETYHy58vtkvk0Iue96PNWrR0Z42/vHaNHdhD55EQpdtcgKkKiwTc7CNuxPNm
XcmcKn0QRrMsUFGWvyAdvlNvb4moTdWufu07N8SaE04t4AWEgp8UcsyXsMbAkjBZ
p9sZVdSQALx/94nSE2G8OAM45K+wWWQgs1XiQAwH06DddMdLjTAo4/PlXonoAXyu
xaoHg9VaeOEOAiih6WRHGB7geD50yJjwyofqyq8L4smJ3mtucTtbjacSv8pUZOQz
xh7TFSy/J1cczVDLWMOktukfgYmxLw+Vuug/EjcHTLQ/gBLjKI9RjK5MTc3Y9eEC
JlV0dYGAcjgMy8OQM/SDeFeeH75MkJo7KFtlSgb5HjoguReli0nq0ImSbL2cqv7l
89+370eadXZOUKrrdvy9mQsfyhKYX8lqQ5rx3NfdEGc9vTng5Q8WcYqFpEjqafim
QZRruJf/AiJq2Hn93R4jj71hl2VuMUlHhFIvZAtBx1MS/+IdequzODTsosrxyOuj
CPfYIzpgBth8H02DL6JJ0O50BI6tHjYlRBrCgeP1m/lgdaT0vUzOAnYi548PV091
qpZwogl1G5fhNs11cby5TgAl9i76GkiMOEMJYoO+RZVXBkL9AhsRNFEO/NJH0nQ3
HA0QY7lsf2RScIthvwqQVq5oBaszZLOWUQi4c/n9dAW7t/14emMWTEQdJqOZaR7I
4iYan9HsXMvTAazyLJDZQCB0OPDzQI+cf88Rx97VB+Dq16+ZtMu31AcNGisR7RaM
5HfmkyPDrJbF6/f4CR6sC3zPcAE7PcaXzGDTnJ9u6UGkYvanX1gJZUyQ5m+UueFU
l5XfmOD/XD4VpJEJemOMADgADhu8bfC6UWxr1MgL3sx6lQpI6lNXVoX28+xQMUYT
p/LQ9hDZ+M/80M8GoIVmoVaVgBhYmKzcgKAsLQWhmOU3QagePE4Nxi0zpRtbhlDC
seiuArBtAFoMB+3abip9MGhB1+5SCpFuNyIZE/5cvcwmfXog2lMRo6rf/JyX6Xj1
ErjP1eJv6wEEZsoBIC7709DDlRJpVI7f4fjAib8nJQufp4e2kTnSc8x5dekybQqe
ndr6LCzTY/QxhoBNA+fawzfaYnsc0tgSWFCiSwhpjOiaRREYd4QBO0hw7x8HDAJT
SSxmM1M3y8p5DtpAeNfK7AEeZU9usuxkFBNOeoWis6mi/bhSh0u3a8E+hFK9Jkyn
WDlKG6CLP+gWlnZ3h+lHH7sXIMwjZ+cfO8TDrVw9xR+dQ04ImeX0Q7/l4uWJr589
v0xgr8gVTiY+zJtd11eGbAEA+GdnoW6UZDJTNAAmtdmHuR/cCCOjPAIDJt9qx0Ti
7MoDuydKfgSh6P+/iMREfOJw0Um9w0cHI3MHndb/p+FcOboMQscfrJPgQGoGqo7y
uHKMjU25LiG0KVKcvvkzUL46Q484BolMYjkxTE2Q5J9uz5E4/soFRTZPHORJrJLM
+wmf4xEPuLHg6ufmj6Slba/tpEXaApbG9i+5iOHNb/4aC6Yz8CwUXJMILYaZGMq8
UImKmOIRb2Cd4zkQjVw64wNonD5yOgqr4pazN8DDl65dn9r5GghevXDNf4Xpno7y
oYBobdnVE6UlFRKXExbT3I6O3NnGF06zNTsO4JoRXFngShekbY2URzhHFPCZ2DlM
7VC+roy0Q5wnn0hD+FRGEPhZuMIQDM50anpqqitVB8WRMNdENlrP0P1pgb8G8fSO
G6xHIF07pSJxcepTvsQuf5lQdfB2FjDlSPuMT8XlO5Vv5mzlSHqT8ParIb2oAbNz
xMORHUjfG5TngrHLgrZKiB/v7vA+FalZa9GSAgr/6Ysv6AwreVf3f9LTq2E0ZHGt
lijXuz/1XMnb5TflaYcc72EhkiwOp0MT4/TTz8TkDzZqOHb1TTfuWtuTkoig0Vui
1o5KqsQdLwkCpVcTmyLMoG4Q2Js+dCHBVp3vakm1VV00pkRJQLL/ALmaPLob1I3V
7LHMmAIlnEE1/Jw3UAHt6D8Js3lwuo7sxWGrWOwPcSc16tLK9IZN02CMCWCcrFhn
QPPez8r47OSkDVoRYYanj6ZgkpQ9T/8t/qif79xck+818+JuWpxGLOcaYoZKwdQq
/k2BSrIrpOd37KfgNY2isybzz1x5f9n8n5LSQBopuC9o63/U2qPyVm7QlwZUM1Ml
mnxq7eYJeNCI5Ol3nkc5Ropf4+gTmdxArMl6YDmUSXHeImURXUpwJ18FlS4Bacsv
Z4jvcY0/BoiBr6/mR/Gzq4uw2hcBP4SQpSlrj1h+H5c6HWipmswsDCIx/7uD0jZI
KUlKtjCBx3Cae4XfxROGAoj6v6y/JrKhOuhd3UzSzSyJUGrXzii8m+m7NsLKtOim
7s/DCecgBkgjjb9oOmRDDmyr5ZSfw/DSYzv/0uX+t6GPugLkFN7Q36duv/ZTyAjF
Z/Zei5cJB3dF2LIuGBqUL2uZCglgqGHMj84dOblnt7mIHJGXEBZwTkA5WI7G23A3
Gl4sEA+8jO0s6F59tv8G28JyziJTCK6+MyTaMoTL2o9MiAAkiVC4VtGcqlGDLLvg
Mz+nRcoY2SgH4DMZswlFEehFT7TLOyJQ8LOI09BpSpzZ4SoJHD6Sj/4PqQAKKw7s
DznWvQhTpNwS3yIPD0fdXhAiRkWUb+DDXP2gHOkWAMzhssQNXYGmaQrXRy9X2YvS
XY/v7WDOYm6ffo+m+F4VdhqYIB52eygct65VDSwxJdQPucjieqYrsEVCZmON7O1y
x44QUMzctImh2GFNvSnyh/aOMBnoM30nBtCMoJzbQf7c5NMrciSfwOR53sujiKEQ
S84kX/DUAx4DkKDVx+SffpwwI+NnfblwNx8QOixGojoPz00eG08KbAvnOQbVMoKd
uSEWK0H2b5lx4g76sgRhEFkCZXiF6yXRoFjxK8QRbJOchfujfSDXIM9NZ7Mdl8CG
Ihwy0U10cnOGUWTWl0M0bz+xRkBeCp8yeDSWjs9Zk0v55WHicrerA8F0IF3pZHzo
8FVfgFNneGvgG5ExIEOwmW/T4V83xZMgz09ujMPSrHJUCyU7oREHVSoDyRWuWWv+
AkvZMYPZeNKDLGErE3itA2sKIYtV/XVL4vIoYZcVOWdg9bezrpfyKffilpOFg6+7
5Ksue4l3J7uyhEDe2j+UHiaf9AVrwa/0M8tivmLAz/K2HWdqVQMppm4C4y7zQpw1
k/R49nhivJ7UZ2JFktsW8QxBUCpYPqXWrlWstXz8P28xyiuzUgOkyejIGX4xY24g
4yBA2r6gHE0TdSVBN9ehHbpCIHwW6ZRldRUSQKF/YqpaPp9QhnG5kZWXU4FHuvJu
Gsq9UQaojoaxFum+ErC+DWInZhCtZYvwQsivj+6cMidPOid+/ERYfpx9URCDPPoU
flGSo9xoGmTmLj7xml3czC4PThr/VspU2ss2kzi7TRbkQSYaAnvMOPQw4oxzVGqs
SKfNdyepd+W3UDAhAlQnLtqfQxuBZqK1tZtq0vA4WoSVnF4qT/wBaRjtTyVvwdp5
Ko9+rvtvMdxhTIS0sb71fmohPqdlTgPRo3y7YENLsPBpb1UDEiYJ7sOLI9Q0WPZK
RD7JfhVqfg+mwQFGlzgqvNkjLqI5zN4HdXFcKN5oQ1h417JxiROATzjPafQyU/yn
62w4lax2rr3biZOW/FpfCslPcjUo2p6KQkZ253M4lYEjWq1dPiqgeNcWavZNrTTv
i+sW6hAd/5tXinnadrzWfFje060FXhRA5BPj91poExjdI85EkV6NOO1YeXhPZfa7
M9Skd+0k5Q2paXhdT2Hv9veglkssHOASQcJsPAIAKW8vAidefd5jwCiNSLBvFaQh
QWMslz04e4Gfah+TqjJMlNDE379QAW0Ri7uHWWndExmHtOZ1Ju2OX2gKGdW1//SD
e0lCz0nXIYvwJzLJ45Y/9xi36eidOsBUxV4qtgwDqfm2nVAcemo+s+pijFW9jAjz
rI9tMDwcsTdtouX8TwNSDQV26TxrRxN5QgMB8/SGq+i/QXY2nXzFKtKw67rzKuUz
UZgTToBVf6qZZwMX68TrsSnVXLzNLWrpIwwAmCp3KveqarHtmLmSj9+AfmwVNeqM
gWYchYTql2hf4ze0CD0192uQ9iEamUOUUwJP6D7R8RLYomQ7egPy9WVPvNwjllX+
Mp+gnxreLQNv10ibx7tthmmsygi+fjnae7J0gpo9jKgsPGpot1PGlWgkjdnMqYlr
LeVK3/wYHOxZiX4II6vy3HCrolWodTs3AP2ZaR0IV8RcRwIlmehZ2+qJCKWNZMRv
xLtVEW9M+C8XK0cTmNaOJGAq+u6LcpZDJShTb1abGSX7/T51bO1nrWd18GU60ihr
mdM4ZA59XPx/ks+GQfpVOUMQ+02zT7QJDXS16+BaLnEnKGu5XK1oSwg9F5D2VSpv
MG3CalJHG+VIwTXgmWwGl9xkfzR0DX6KlZsBZVCCpntGE0ZlUsRa+vTdOPW0wL52
l0DabGt4+w0d3NdCpNZJVFDArdE5WCzJEfmIgU2Y3cwakLUm5hUTyeddXqZ+KUeQ
ZAp6Y83WrJAIMD32bvrllKPE4Mz/Uo9FwjliaVFLnAZVTlHsMjJu6O4QCB0TJD8n
FdeT5EyWOoihJBjrUq0ogBWkbQpdzwUuIxFg3lIPRb5P/BE/wjzBNlIMzCCak73Y
/G2CZifnIAhs/R+GySS/RshlmfW49ramnNz9FIcbqoBh6LYlUfqQphKuzXAtvIew
tB3DuEV2yWf2n78up4swXptNFoMLk6J0LQPu9iOwVFaC5+ZIartHZAdTYLdboISC
vuHHcxmglWxCqEuWlG92LinYOZy5P+v25550UZ8DNnb/vnOpoGG3SGiq8YqZ1OMn
q605fSzRCfrxC1OiD5RePVtyaw/5zPgWD9z6IMdUD66EGtK3OnSb+3T7lW2L4JLk
VVR1ZGLM6utgghazS6S64Yckxy1PivWx+lgvZAZ7z3nxsweS6PwkIJYoi1n5jJC0
/LH/TFetLt8VRrrTk1n23Nkhh3fJ29eWCGQLkldvI2/LNnW9V7VruH9Qf0Ol06g8
rOuCZnkcIU/dawC17lc7x2jQsRagaIobTvYZbeh+c+9F9qpud/VWxTDxhga55oVE
6D0OJQKT87jAcXh55cFUPU3f8u4uVPdHnU0v3L9jlh7VH9oHAn0EztKR9U12bPlF
V3YRddVbfXQDxHE5dDUKdU748/sC7UN3NrZeKtYkmY3WJbFk+kKa76ETng4GEsfC
25GYZGnv4lqquwGcZBe4mIrZ5pXoMGd3D/Vbb7EotRxt5fQqjIey21Uc9EjgdcBu
YJ+ULoqC53v+m7MqYpPwtHxJqgpQOHsTwyfs4GnPKOSsQTCNO0XUOmenWjwnF0t2
x2CVRggemAQl7CRVfvQh6bJtgmeGSrzxsqH80BzGKyMMTqwM2OgueRhobNW1yNzC
IAX/BkwLSnIiBf7OCvlrIHond2646csGnQHz4wA6tYdvO8wQT1MXF/GZL+XsWjl7
rMiH/fREqhIWzRE5rRsVWW2z8coIGYp0i4h8XZk4Mw8hPpwrTJ1UrZPgb2YPiNuI
z1C6Mhg2AS9GlOyPVSVgyd83UKhNwzbgPnatQqkW9sUWcmAFHZC4ePK6JzqS2b3S
cMkJNl6ZQ0UqPrq3bi0I3eDkrQy8YSMljUMGj5xf6vmuoPARbp+Y2y4x1esGXmDh
1OtCdH61fQkOcfYDLWds8P/QqYKG8P60HmK7SrjYUdcn8iRJurs10JGb3ebk71S1
Sz6lqyhsbBcW9UoYhHkl0bnrRIrEgXxyPi8yd7qo9Z0crnztQHSrixW5TV5twasp
r14ihDIKaL0Ytbh2PBazazMqPCxw+OK2Lk9g7LdSie2mn5EUfbvzrNbD8Zzi4UR4
KuVTKwU+3HgsWpCYuozoF1UKyaMazBmToT+GYDu2vmyHHxIiIGQ/NRbiRjJF4UQI
caaviKGhTiP+Fgm0aHcRLpi5LpOcrgp8i/ogO7heJRMM4UI4xwm+6lEH3vu2YKky
uLK8D3Xid3V/UFBlh5LoTV2CfXwcAbaOzy6eevVNrPd51SC0TchTu5QKOFdC944z
4NWS8sjCnXH/vqBtifMWCohQu6vQoKftS31E6FaLLTyXT5I4bwOSResHl17yWbQ6
47tOLn73zwbLkY92b9Ur5rdAhSg3yk31LKDXreAcmQnxYZvvOdinmuX/HJEUgD5K
T/RIzeriVOpaJ8qWStA65g4HYyNTQ9EzXMtyl7tKUkLKocqEenev0w9vPShcNMIO
GZdXWUkm0rrkbhJqe0kE269c4OwRufKMr0BEi/VbSmDwMXeJrZg1ylUMY+wLss4W
kEXScgvxaFStZYEmNG2ldkGIIDukont7NgH0cgQomWI6lR2s8638KRejGjL0MfnY
XKCqTzfvANKQkadkzhCxP2AIGS3vRzX9pQFHwNFebefcF/81dm/1vhIZoyjknIaC
zFWTCLEBgLQnoDNjlY2Gvek+XqY5Ga8dGaeM76loVVYrDUOloUJaVwSy+rKPorxP
YzCrcJZnYAShz2Ba+kZE3Kk9COXXp/eWdq1o8YVYnQa0bxii5OXxGs0nXEvSgbIl
R5yeeQ3BnqvwlYfjTWwmlYIwOWUbNYSPVMKDPMT4iCMmGsrBmEswq3NPR7oZ8MPJ
pivqHMBlPPSgr5Gyx07zD6co9ZkZtVbztzY0a8LWLjvnz5pzHUO/HoQ5I27EAYQt
/ay09kcEkpt5OP2NmuqyuVlFE41wIGNbhDlXBpvVLW8cANceERc6guHIQEoXmJZQ
4wlIdNSZi+I9Zd9MX/Ak8QgTWvQrsnWWOYrIg4tNFiA4UivC9Snd1JKYNpTqNbJK
iGviG3YMoCdlpn/6Yij8ZxhyR5PbOFLfVQavbAfnaj+rhB0aHcqEb8HMaFXZ2bXR
nIx443YHvrtVmuO1pX6OqfSVEBlyfIOS/HumRTpEHsKaM2C1zrYBavrpkg05fAX7
bsy4UtpVmqSXco6Dz23YrWLC3pBtNHD/cgEhytU+Hr3THkayALgM/dEPBA4b8dHQ
t9KS22+2TjF9jZbCTKfO731NWIJd6O9PpA03kIpKqiw3xwXmUg+fZj0Na0nZkCA+
eVPaYpdSHhmXI8ALB4wc5Kp2rmlu1RUi33qizpy41yJsFhq3zxn9/uIDmanTdo5X
mm29TcE9+iOPhGjyka6KKPLAxSTVuqoGuZKFRc9zeJNjf+q2lLzWSY3CI45lkNkQ
Homr+r+kThnLZcC/V70Th6v9S2z8U/pI06UQkrQuiOki7AMilZxKTDsrEv3NbJXq
9wIC4HruyjyJLqv4g64f3/ITRt+S4h3fPv6Anedk33H+BDtKapJ8W0hte73lY8HM
EiAClrPb9gbsS9iue8bBk0yci5oY3GZLxXhW4vZHE3e82QRoEXrv6TYIS5baeqHi
z2lmW3LYURWjCnp6gS1zF0PSYg28CnSnE1xzw4AFO75l5b1oF9/PIi47/NIV6Fec
iwxJgtOhjVmw/pYmM2PxCURQ1PsnG9s+VuOiuGc5a8hoM/LAzSnUGzO5NtO9BZBr
n77LNU7X1z2XcpnWFvnLTrn2UzqPiZPqQlxW7CkrZuEI9Tar1x4gSwPme9p+gP3I
F0oWQUACYTa9GsvIgC0Oho2mkL/vDEtgowp4WotBGoAZQWvg4wHmD4x9e8ck8UoE
TEXt0EuYL/d5h/TopoX+akR+d8J2viD721rSCo/JicTnl3n4SN18NS9yYHTIOHId
x06Rr+PFSoP+I6ig6PY1prH6Dr3IVVaUnRNeM3yfrwvRLsN3wZTS3Jgm72F53ZD6
HMsTklNAn9Tmx/CAO+mJYTgfdAcdFK5I4zhf++XCc5Z+lX+SiRMfGZE/2hwZ7VmO
I0UpWwM6l92V2DWxCrdeNrC1ztNXDp9Y/WSTgwJlQbOhvEd5yoLWAhZCUYdsRyHI
Ut9fZxPjQNCP4R91J5VN4/7WJhlDQ4cv/FrMNfFKwX73sKvuypXS3xHsPa9f9KAc
fFXes3s6WkmkLLN79p3OCPYs0hqRf3rJWfjX10TFbzbbYvJ8U1QA4A92TCauXe2U
LEO7XnD0nlOgwxcwwyFfqIUV5PMCE/XIHkfSXNy0KiGcmW6L+/xXuySV2hi9X8xE
RKlm1DXglngl+xIy7ATx5e3PldLXLTnN4h5lHsCrlbU932EtqhTyhZZmQzu3ODZ4
G8l22JUnDnAqBdPr17ozaHtme2mHT25AKRaz5BKBDkCrnSxRBSIsJHbZWUYFyraL
eBkMoSXpTo7OyaxxQaKtCBM0eZB5MV4eMFz+rlbnnmtvoSxx75Xgn3iRRWkZF5ZM
byvvAAxkRKrLYx++Cyyhf3WwWptoAAWh5mP/jtr7kma/8mfjSHq79aURR882hKGA
cFPgXcE39MSsd3thhj6I5X0O5h0HluBIMRjp2gEgX27Nq80N3W6Tsfi1iRxPwbhd
GNihE+qi7ZK1ElVHqdmmJUyIQD79EgOcnUcrZKSlrIalX86VZLSQbTWXaFSL2wCL
2OXuREx77ykq9dHOL5rD/CZdlBs43QsbrCyfwTEItLw2QUcdtSS1i/mHPHUmV7qf
Xcf8HqtRfEJCcOqUU5qk9KpHDC0CQQNdv6Qw71w98uqD6YQot44ees4CAbDmoxAK
7PizsYl40VjqEC3DdeD0EvTO7hV9qIR8Dz7ASg9TDTDbj5/shBSMwY8P/yTB7Gap
lvn+m5oHOOXw9mZzmrmDLgzm84O3rnD8AKeL9m6VLMmS8FGKuBGdLVOrds7sMdYa
J4T3H+J4zHTvCQ6ShMg3jj3xZqHBF1gdgQ0TdhjoJDmXNNZimmnzMZKFuqioZ7kj
ha4BBF6+MWdbdfcGy80cQrkjSLglAvZrmxu9g8uv6haujHkepHwSHMiHckNA6Y/J
jqSo2Z12pBhkvyen6V1dZIcsZdEFgTJ+N3JcUrq1bALq1OjqJXd9Ew9BYuIH6d3M
bx7rGRlem+15Elkcw7MPvS64JPtHbgFbFg8RVrOwjiobpDoTH6lsdFZT3OO2Fk9p
c3OoXDKjVSJeoMaO71XW6+alJ4mIYka5aIIljE4DGxfwrH54MiH5VvnwgNTnqdMp
iUzdujAu8GIMx/qB4iVzH7Xvst5J4H7mdjf8yajlkzjxtq0lSiEFcfk3iQ4XrnHm
ufNQY1zY5BYPGz0hBdavGVbiSm1AemMgpiN3UhEjswaP9fR8R94T5HG+AyOLX2sZ
4lrKM0d1DNrt8YT2u63zdEKYXxXD+3/n9xe780bPP302HmJFVg2k0gGkvIfRpqje
dsojxYNZD8cly3Xw1kqP9lJm7X3caFzdv0yjOiWWZt+dLcu81wbrIuaak5JXS6Cu
FMSHM3gZfAh8FJ7tpclqBZGQlt3rCpijhroQXuyAoM7DdFjfF2HUdI4KgnvqHh+Z
8LXOhj33SscQCbdwFAydxG7WYb53Mr3d6JMkXZJHmbep6AR0pVfkzGxrxDw+FRo0
4P69Wu7M2zqTIX91Vv2GEDH/OnJkaVqh2jdh3SB3vWSBuIRuIiaoCSD2HUtSDp9X
9/83idAzMYW4c2tt/MvmMlRiz22gbOoYwwYWvgTlYlxQIIuRaMuGLAJnEkfkQ2vE
dzdTD7z5+jlI30ZpTCQCyWEtgwb/uLTbnRyVt8xC15h0m9m5J7HlMo0dbwMLIghd
4D9N3rDA4/C0aqvtYEjarWYbZD+9CvUCKVEC7Jto2CIfpwTv1xG9FCjUxmE+O+JY
mwSX9bSi/Md4E3x3lS65TZbfFeMgnVJ/UQQ/8vtyBQ/lBbF9hKzkRdFkZk0NK/rX
LWhuJb34WzD2LgwYeK/RQUqLeNjmB9noUynMmPxZVjOkSx1pnNvODkBFsEOrmnhf
d24Em2dm2DAOVzYd011VpT8KNoS7fJLQXf46jA+a978DDXdnwTLiJx5JePalZ0iI
4Xc1MbGtGjWBt1uHKe5LUBgfNJmsH8YeN2AZ1qSGWurUFTspGbE/him46kBSbopA
snouu85pI4ICawoIiWDhXl7wY2XRqPb1t2Cbbaye/BbizGU6fuCrkzVDU/h0cCL4
sDhtaASs16bSti3c3oanITaCbdP6rFAOaAWuO+cQ2HkcuDNem/72Prfswk2a0zx0
/H709jfdCoFl6WAJAI2TooEm9vc/6J98UY0TckdGl6eTOycdc3HOtTG6obyi/tFO
lViF+B+w8fTE4iK1lYS7jr1l+dqrhTBICdzvJRky+2cxM2GrqKdjsVp3nKBX0x0i
IK9Vw/UHCv4EWeJ/uwqASpC7anw13XQjUfs6PRJjIH7P8dwzb2FszG8hEQtEYElb
WiCrrmNnUcvAommdXUHfbSikZl3XjS8ZpbqZ8FISc3attAVG9+CJ1qM75flU5c9/
MYA0U7Etnk2I/u2a7+ty2kqqYiUeYPff9OEQrFnpTt5h9XHoaYXpXbyGDn7ZiBNb
GJxwb0lNArZFlsNyZidI8Y+him8NA4070Mfp/Tt7wL1muQrPeulOh5bBkMCwdgMT
p+zdHSNtCxopy00Gf17w4CyY7xyT931qbvrWXc48LN5j9DMZHPFzh3uWNlJKZiNq
55D9DmxKl8HQbjQWucfYv3hIgEWAbYOYPGtogBbfuV4WMcvC9v10LzThrvqUDSoS
cS1kgL2yYimkc91oPVB8RkQuPoG0cdE753/FDjuJjxp6qlNoMkItDslmydReBDDY
anCfEJnbq+zXQ0r8A+FU40CyyFFWDKQNw5WoRMPHq6lZpOH16kUGaVjmScqSFKYS
Ht10JeqvCsjNCSpnNkFUxQYOq8KaczUYweJ5Vi/0XSLZdoYS2LcL2dEylBTsk4X5
pwQYIIG1f/3WoPLyRlcr85DjpHekLUyzlkcmgUPJm8E+yA1N2xYK2owGhaC11wxR
8ywOL4RUziZk4An6QX+lCeazpa6/knkHD6Fop3hB1uIqjwRRzRZ4Yy2Zys8Y/Wga
kW83kshh5RwP+Beo6jN+OExeG5bD3jIOQOsfE6eeSRjFbK1GRvuSzivAYYNV2gwH
d4swFg/MsU4CwzRavurU6el4BZ7ByyAtsQtacGyrJVxIOIZhm2P+QV62XLyKx3/S
cXryUgA1qR/sZqLCYw6jI6BX0ysfr7NlP+pkis7IJrW1LAGqT/aIvMY8r8JYGpYa
0dbM3HbP2IrWChZHK5z1a3tMAOh3lHrDEgl+xCCP7acmA+Nlbnp6aOZlx5UxT8gT
Wux3nyvAhD9XbKL5rAVvfkLaZnaOAsaC7Xzw/ZacEDCD6IBFgmD8O3wF0t5N078u
N/4LADgqiIXCtRwsu0aVlvIIc0sSkefOS2PC+a/FdW/9XusPZ00nXmz8miLgnAUP
J6vH95H/edk43Fs4bFrAo57QU1Kj48KzpHKQCsvWklyJ0k2M5Mlccc9ctcZOPbU8
J5dMPo3PomKaNYrTHC6Xmzy6f2VlzXzNdOL3dpFkDRF1pvFjFrHlcEhTXB3AqMqa
noP9Jdm95x8s2ysL4Xdr2/DNHTUNLsIIHueNDV1TQl91OKphGkQhfLL8ybGF0Voc
eJ4PqwUJ1YnGMvMkFU27VCj4cwrJSNt7wH2qZUTN7HH9CCv4SOm1lE4Zgg59tsFy
P5NTq1ojbP5RShbcfsfGBu66Dfim8yF+DpScfzY67nhbDhY9DyQcT+/FqvEZR7FO
Pi+Hut7dUyEf/9uc3x0yFwXsSQN+8zutm2V70Fzzfs+J1FJ99nE8L10Kz4Lgxz/7
qCCcOwJfCD6LNjcg2iLSrkdZPvTg1U6CioZaBirWzk42mfpXk/yhmmFzRTK9WITV
dHW2gt85b0+nEkrB6E6rm7LmE1PAywo52UqYRaJjo63xuWDSPc4+42zEG5o0DH+M
buEFuKh/2gG/XVXxxtZMM5jvPV5v0bTI6LwLyWrXQ/o297lhzTYrqqNTqr0xTtbb
sejOLCwNVXp08xJN0I1jt6+DmHYnZyFImoLCgxlC03tGjxB0p+/TYxRvPmjcNEdD
/WzKzziu1BKWlxJ2H5hRWL/F5BDyrQGbkqSYmvPLqVnCoRtH56XTr3XR7O9cU4s3
HPpqgVt0ww1RiHpcUo9paDxCTjItM+wDQUO+YGlu5XpfdeqEEHbHLLCxUgF12TDb
6vZuPxNj3O9HI7Eo4loEEbj4WiUIUJ9fUpreVijFS5yhehZfnASiNL6cjxM9Ws3i
YOGtqrt1Pz9WyfZRplvatHQlbjZeQPwbdT+2nPFSTko+708+hyAnGOv92UIiNimN
SK36nDnZm2cZihFgz9+v9hDuUHLotnsJORRg76ECg/hVX2qRiFOzWyKjETApNOtf
JYwuLTRJuogzyv0HGUncje/i+pwZV84Kw59W9bN4rdsJz7vRXNGI6rb20XxDfa9q
hCTj0LvXFv0Wgjxf5F4XF2hIYcp+YymOOl7ZnL4EJglvvXnuekeH5Osnoa8lscJy
/65HntS19WJ8F9nGmHahoB5m44OwuvZTPYbC6ogtrPvaHvnCnakWymk7CEheOT2f
yseI81avCEghk0OkYisuFiU6jElC8YtsfFrQXaJCD4eY25gVaxrx+UlI7ftYW4FW
zArM7/3Yox08pr83PXGcMrn78YBbfnmbvRYQzsloEUM2Y/Ef137istir36Vcw8gy
QxaCmtCb1wxUnRRQ8QUAP3VMCH7YvxHQ5E1te1ll2bDpkQ/u+6jQ+b13/IAhc+FB
rVE2SeD9bjm6DNB8pyryHtExHXMn3aFZbbOxRokL9FZ5m6GevbnNOBHZdfSYtXEP
I0IHKqzL7rcBADMFUtffefN0B04HnMWjgS+buDYwqOPQwpKmJPeUg9PEeNjDnJz8
Om/CukzBWdMy9SMdkwD2MoTD6lMa0mRHiMrj6TSp26udPMwC9q8GdHchvitQpz8w
7vO8FNMn6qPyt72pRKFarYSbe1Jq12weMOv2zrICQWufiPTyO7ObshwQx15drNyh
DdnHDE47BCL2FQEfbkybfblcWCMQFFXYq07PgbXzAk1I5BsuBxuIYX5LWs4zQVbI
O7YnRUOYgA2zc/HSyl4lrloxd5VqRLo3w/ZwddOp0zJYu4Ye4wniJZdu0D4Z62mf
s8bCKZmmBLgSOebGcVN/I2ICjC840h3ss6fa4KucZNnvt+N40I0pxoSlue3FwhC8
vwXDsLHPFgkkSIKOaghcGnJKsUj5Xe+Nc5r0+riYiUrGrbmY7fYR7rygEIPXLr/d
qdjfQNHTPFY4wF52qT1+kGmzXZVjm3zt+PXjfRMZ8eFon7Q8cJE7K8CpFjXn9QVQ
HhPhbPZ3c8SalPoNlYcxVYFwLsTsbvMjxuC9QzYNQeEVsgIXsp81L69LiQl1yfqp
4bmm788nuthsmiL5RH7dhMlWVh136NQpYjR/N1WLksWR7MzRgwMO9G2lvU6SHDip
90GVGPgIVwNbxeheOC7MgbJfgEK7XtDJs2JvA+eQnxFNVPtnFqpYkKWbBVFMjCZP
vwcBzpv1trBqUk5MilPSO7DW0o60wuotv56ubL4MacnLGuuuQk7qRa9utYZmr/b4
53544RByarcVZhAVM/ReH0ikB6a4J3J1yAZduGjGtveV6lx5h1HVISZNnGju8WtG
1IT7kdPHeGn/9CxPPiMVkg3pLH41xR/4bnX+RAska1rhX2mH3OIO1Y2oQAXvO/Eg
ZDStcyTZt3GDcXph0rHpcScGa251GaENrZqK8q7Z1Ga35Htq0YePouPr24anDi3N
VOb20a5lhnjFtAAYrGuSPB0xdHHhVpR2Xpu2B+368ZZNFo2YvGEuKW4M5ZuHz5qV
FdwFT3vCaUkviaia6oiYxZJ0d/CppTjH3Y4aCbPl3UEDMPG7SSSVjMd1UtFigEdy
WA/oCpwAwKLxZQhvV8Ctrkfh6DNw//xM2678qN2CkFDNzXTfJ67tjO67nbpBY8Zh
hvLv51Sarxj3V4lSGLZJnSx9v5+nKg8rURgOUEBf/ENCUpuac3n+sgsQ46UKOBVW
ArvE+Y8REwHGUVDdmId+2OQ3uhONidSRbdANeOIwnF/3zEmGVtTIjJPoYRECQh1i
yhTCdzOzxtw7fPgF1x7j+y9F5tBk7zRfuntpmSzVOAqsPNBLXCGtPTCKZ4dwPy7g
hEmARLGOIpfN3HOmxdeZUcDM1E0rVw2SzDbotlisr/KyeZ/Tumln7G3WChA2KPNR
IadgHg3+oaXvNg7SthInbQDXoOpCjngMOWsPUrk5O9Cj6NNV7wWSxr/Ht02y+ir4
aKENsJIUBgyK1tTpPGiiGeXTjXcKGVUpAd6JTmZJJs0rwfBUqKeP8aDmoQy/QNYj
iDV3BHUMTuYobE5Pbr2UvdiiHwThMhpvGYLrdMtC06ToOy0I7XMAd3iAOsz59JR2
Dg0f4cxqnWLH6VPj4z3UH71qEvbLxZOceaK+8es445fKpWhZA413CLQ30YY8XsnO
j6LDdO/W5LYf8uDu3g7uzqoh8DdbxBLJIUd2XgB15s0OjxiYz4jXA80wGuVmuEBi
B3yGPUeFcbs2DBa729SkYqfBKo/A5rcHvwwMzsMC9G4qDlCnvzmncFacugnewr/9
JoJb7zsMzcT53h7LvUn+VHiePny/7fOUXYHOYye4HdIu4BkUqW5xASa+t0Rxf+8v
nenKSmlc8OWwXrFvrMhFa/x8y0jfwxJufPUNt5KC8tk1lFTzEhkzE5Veeqt2tJqY
gF2+qmeH2EAm9Dc4qK8MXjX0wgk54qCHl22n2coiwTCjWUGrcAyb6vgq0f9glUzq
JKHI6bnVzrjvTRZPlgyoixbWdZUVAaYnSqnzeTi/NnssmPZ2jtaphGA9crcnHzvs
KEBuiDaY1SH4Caj/7W9eZyVNzGYMH937YePLZtskp1+xeGJfjNo2agHdWw0gwEmD
9009JGw6HBQIgc6z3OF67UYdR28pP/O7bhjM68Bg/uFn9zaxz5L2c2D9AgFtkwWj
2HQQbHocf0t/1m6dfKRkkoPLKiZ1gsAEIuYe+rjwFFDIR8xd29OId80+90pyHBbj
CRBoBXTGsbQWXO8ELjsKjjswSVerpLYkR06J2EMzUK4JN4a3roX9RP2/d/+D+Qql
1G41Ets5vExkKUPQ5d2CBeFtcvWjHOnJcZH7X2UMW+tcGR2fNqJ4UFSoj22pkVgg
dj0ER2hX6mmTaiJ7vDE0hAL2Fs7XrFmaEPqceby+rAqHURU8Dip+LVHux5j8SV0+
6HtUBE5k5e+1Kb3VjLcRB80bdX6E1Jws+mSIKAvVKL1IbKAS5WNEBZf4qsyYYZ1i
fPI9/07f9T5zMlOtfrBOGCYvgoAd7mPqKjmrReBOcftwbgWwbtx1ogYsKT8jZIda
tlzZoaD8IO2reeaM/HIys8rwv3dOMUn3K+MUaDJeLrKhs87AFK3rXSoD9VB7I0w9
Eq4toGay52X9Yr91X2cn832qsIj7DdzbLNFee0hYCyo7U4ZhzcteEb9gNB8T89bP
hmMsfvmSgW0ptM0FvSC/6m+0TIIJ5eZgpVEVFzXRG1YcD7q+6r8SoPSf5T7galJO
E48SU4dXpzWW9lClgvshtMQZsPBpXNj30Otzec7Tiu6gMAWh2aw6eb1J3pzfyB2Y
90RZHY4BE/f5IjAQBT74B2OWjLDj8oEA7PJj+CMXGWDAyzXT75pl2U7oewoqIxUe
coy2da69uwnAKQcshzYGWhVbh8fmq7fVzSeYyhmH7YtElbae3Fo/8Hg5UhDbz14p
YBYOe1sPQ1s0ThlFYmX3eTWPIH6DibjkirZz2crhuBJC/NVR58VJxdyFJDSCS919
ASwh6u5cCgdy+A7WgIXuEMeiIrbw39UpdQ6nFzsXQCMzy7uxG/QxHftL84i+/zrG
JD0wqB+UBWICB5LzyVpLGD+Y1cSdiWdBefgtQeQHK2DKkY0A2ZxNBC4SXVdhqNIO
AK5/gVrLjrcdoLKhzTcuGJA32eJaDI/bMVhsktptGGws52FxWg1RitCVNPT2DaH4
GRa6jppt321zKDmtmv3cfj3toHXsx4B8FJoF7Tuhy1JlJ+r2EJfH8IB8ZsOP0PFI
8N9n2XSZbp9CAFJBye5ubgitzTJOguBcMNah8aBYMQGIetd2KaYbcaiYHHDHWlt3
OTQu9JDU95ru/ChgT9WDpDherxcAPunLi6eLCCXBPcQonxAtn0/V5FeSNCSODR0e
6blhHrld0FO7OeRSPQrEOIA1WiXxXU21YrfItcqfd6MttDR4eowFUGi8bbSDwF2h
8tGM+bNaYsdjgWC9YMhfHnroJOxt76cze7OMAhnI3+oMfvpluBgEIeyAxkX4tUk6
f6U97QAJyp5jF9R3Qy3tJG5qx95ThKBJrpZdY2cvff9kAHI2mrChwkDUE0elpyY0
PHVdFqbJlEd0ISSwilEqrC8usmfdeAn9RHxZZpxD2T6DWRa8PqDT7tugDq+g+Aw0
R2RffZyiCiFKaoHxDrJXcqKhDqyPCDrTYyfkQITMskQsEDq/OG/xwMBkQuod8I41
P9qgM9apHq8zbyffQI+wM3fNHvlgptM9n+M8omgrWwW0thHGyTkjQW4/UtmSUG5A
wnnEghqS2pOF0Pd4YToqTfUuyCZcxeGIUy4nX9MVYSGYWPluX5OETMsi0NKM20cI
N3ZwhVU6GmO6hMcQ0ZBrHWCDmlwzhp7s+PXf5IpGj2xK/SOdME8zVoWT1pEnXqV2
PCxtcDJnW9ddecbdk9ZEH2+8bL3pVffOsu2hwUMd4IfLqMHKEzlacTDeepu38GhM
BIg4jVRAiH8dKmie5mv9+kto5mOvTRCzJoh9p9u9jd2sKPdyJNaaQF6+SfWB9UFn
7C8bfxSZ2uqQPs8tr8roELF/uQZ6V+SQ/UblAAzb0OwrqAia5oC4/gFeAznUqFr+
xH+ie+IHgmFaDp/A8EfBPr0L03UTC2yAr5Gj+tEs8T98PQNALXrXTyntK+rXhsiU
jfeZz/tImcOd9eo3wq3NfJXjG6IJjJWjAK1HMG7JneRv1E1YGzlFxo+wqMVW2J0N
fKmLpj81dLXCiVWqocIXnTFQ7B+vrAuAzqdna7QW+1r+0PpZrPCwvxKb0rQHdoyE
lf3TosiWHMt9CLBu50F6SZWjWgXJcJb2T1BhGulcIBIO81WXnsMoVM0mhYjb8iaa
C5IjbJuOjB8QHGZPvm5nzmn7B/n2VbmCOOsKips6phUYtnBAP9FQ8rMRUd77OutJ
yTnbH1Eik/sITT+kAAw+/RlmA188lT8yS8otyoXzhpV6/urdcdDK1Hd7+y6Ww5gh
1zZL9Fc7S+00b/+s7zJYLn+ZwV/e1mnEbSqaAqDrd6G6RV9j++0dS4F83UB/QQjp
3MKdgIw1AibHODrKDUrP5iOHQiIf9LzVGspN/9SSgfFOmlfb2fQ/26WPxMCNwBBo
a4VAJJXguIw+VY/4r41JZc0XIs+25xVXseFMfEt7z6lTtZ5QCQAWhHuKluEayKl/
3QqUdLCEJqwDd/pNPVu8Q2k4doyk7DhdFL+oEAKTuh66tOat+rM6z+BhQKGs8HnC
x+8TE6oVt8HEHwjaJCcrFk884GMT8d4jynWaC3DV/B/R2B4IcjB4Xy3jD7OuKbMp
+0NgMz2YZV8jnPeWWN9n+BSyy6bR8jhIa472hSf7Iu5ewpaLNaTqEu/bvG5+0MNT
BWnW6GV09rT1Xmc67gQOHtaciiqeYXrWzggXIclWXoYoIyp16F6n94yELDS2i/iD
83R0C0u2mmUllDfA/ci68nXFqjiv3Uj5vUL+c0638Akz9Y1yLmBzmPV3U1LWCE39
YafO56xqQ74/uhYZBP++bPm6IsuL8EcWy7ExBh8391iPYftVQ8yM5VNFX2VSI2X/
FRvcVhJTEdvwx2Sc3Y/4X1/QSKWMRo+9eRPJ3sIAUrqguUm99nqDa9RDLh4HuNve
hwYrSFEQYUElVZheSe/h5GAnK2P954EcygzykjLq2ZiXqHCUy0Dh0RZwqp2/xSHN
GIa4LlafTKCEVfhOz9BolErA+JXtaLxddv08YaIftg1vP9rtiYCSuKd8NeuSofDo
L3fZDf/P5EQYrCRwVcP4Neyxk50iedQ0nwC8qxabjVO40exkHluWwmq3CJnxbwfn
8FCHHqWEkms+rgqNAddAVLYNQROD2BDZ0BEEIJQZr6V7RbID31dvqT4h1bHCFMVC
Rf5GIegru2t3TpnWncPo6icoCm35gTgSgKMinr2HTyeHsN663K5+j9nP0/R+sh75
BgRVoEhhek/1/IXfs/sezF8i/2+09oc9FXJgxHpg1JVWNeTXEI1sgfRkBVlhtyoW
EK6MB/oNKlds8O2ykeHjlymrKn+OwDzkTrc/WUFNS6k22QAdT73BFXt3Mr9tPT4C
Hl9VCoF+43XR0cSM/C/qW6lXaA/I2iK4pMFel9QP06xI+ufBxc4TsNKJ5pq9bjMx
Tyuv1a0kzvnD6Q5So30zLUEA/e7pITi0GCn6dEJkO0sIYazifb97iAPpLf+M5kyD
PZUiaPD/E9z9BEw/UWFPdLeKmryzbhjEz65bxxVQIm2hQAso910rwbg/pEKlgYp6
uv/bUJFYsWLCHm/L/TvBqzQjRDCOmAnktS6J7VVSY6UWq6U+xwjGXH7meqcGUfPb
yWUaok34AB+LbqKH9BakLgSEQW7eiqKfZzUWBij8mu8rzwr4viizyPNY8HuPvKPi
Y5RFG8oCf6abe//eU9Htf0u0CRF/1vZxEGCQxaRwctRxHhR/TNnkmwA/ggYtOaNm
8ilHn2DD94tKLPNRdfO2Em8lAhCkadUzMJvI1n1oNtktckm6XZdZrOzIQ/HGfIP3
98yNHbwQhgRkm5bXIehGkQTOq/IM6PA1vGb/arU9ziT3zkHQhZiQQljJF00KTRfj
HrrO7tu6jwa53NH7dEeDDgrjOsP2VCWs2YVm8Dg27+VXtDQDoUyabHWzoJDUmeuS
wYRpwjIFahpC15nHuFEwicziGKGZlP9gY+zo3NgeoN/QOsIwbGbYnH345XIYYxvR
SBGnf40/pX/cXPjeW6zOYSSErweq29CcHRigWDvNUbS+E5DduUVSDUTydUGLGFqH
7KxuhMdThHFOVlgOcLMSd0GL9UlQotddSzIY1DljfVHh4JlzGF0fV6XRvoUjuj1M
XMZ3ql574M/hQN+0Z9Lu1PXlw9/RTuKnjjZnG7rpDUXhZxdPag1D6am6HZipBCbW
LJ5Ehcsd4T7Lr/wuwmY7Uea1lKOTjRhN7lakFv2u+pUoIVmJDu+7pYojsGcBpa41
bfwc4/0zJhISPKeuz0iJxdR0//tenEFwtgK69U+GR8xBDnCTIpbpae6+9ToSxUng
rUjfluYWty4grWWW7t32eT9cWk7eRpdymNSql6Yqlg4w9we9e1Lb9DfFn9+7biGf
1VDtoC5zvsUMmha7sRi9kRQ8CXPinKiAnCd/nhR1siTN+4RlLSs7yEz2z+SEHTCN
/2fKjfpsdtKFO0PgI2UxeccP8EiN2PcXI4lYr6zw9WHj0Fz+IGqVYSImzTNsUDjB
hl4MXBQ0xnkG7wZesj4rd0oX6nU4NxHiPQ28kXbSjYC5BFDlc+a2sG2yhHpn3Ke9
GVRd/GUrV0bvZhN3H/iBxplBd8/0fFWUISGFczGg3yuuvHTinNE1JzEK/4DNHScz
e2wogOMijuw6cof27v9q27U55OnSH+2zheHP/6aOnQX7b2XatvXDMnIvUxPXUlLg
66t67D+5VW552JEYhRfWp5TV357BNBV0H4iWw/tYg2k6nggwTQS/X91/Ch33LnOu
sH6aUa9gZhLv0+m2Uw68/WYLu3a0OFJ4JAGNhYUHo1RFGiAgN2+XjTUdViu1dUar
oRJCidGDHc94yvNvcOaiTCR+i/esZn7L3IhXF3w5I7aDatnCvlTpUZ7Left3awpe
M7FKGF2UMZYXuMBDHXd+JE12lT/ZSSM6ujH8tX0tl9W4umpU3irO/lpYMl1gqGb7
QytG+Uvdrrw4FNTzAz9FPQba04Dma1uww96jY63QqAeJzNSSUSs7GvwhIchl4L04
PTmXmkbB16wz7dJV3kcW+eLwhl3gnPjOMQTz8n2gj3LR9Fjh1FMQctfpU/vuONPM
0e6YJQzzsFxv8OAnIbdPunK3QJ2/FwS7q2633suFFO/s3TYFvpArTlNxRx5a39OX
2SHMPz7cl7Gghjr4S3WJHFacAcsNqH/jNzOaQTgaWIcxpD215FkICiPGiyJOn7DS
ZPCav8qEIkchpxDdWhtFt8LuzCEWiEmPcvPWYbeV+y2pCdeC4UR9BT91maKI7OKs
cdJrd3Jya/I2mBzh2pXN4Y5SxyjhoZpiODYkXuhi50wV4USQebTO0uh7pp1WTSS9
gkRvddd2s4s8UBCI4Je4K8Jiq3yoNzqHwh02SC46iZjfeaNeJmfW/TZMojIP4qEU
Ptlsq3VAhV3qhoLwNE7ulFigszWpkM0vvcyxI3qtrmt/+9ZyiuWvaSXsxrG7Fkpc
Hu/Ug5hQfiI+ulNoEaFnieY1cafQKc3D+1kXhi+a6MZiLP8C+fEOoZE5gdTFreA6
7nMEqh7dv81l6vBu3Lkbc9p/snWBtiZWqZZeEJC1noo5xgoHoO5g0xnwTTQbM6wR
c1XynBZX/ZkXHPqvMY2odFrxD2AW1z8uxKytrgchT6y/wZHMwT0oQ0nVcoJ+Blpa
wdmisgmfRn1iNnTERdXUFoUxS9tnzk43T9sxyPhcMIIuzegFECsju1Y1Jwgf8g3k
E9t/K5LhO15fyljw5glSP/9ZCW+PbsdovmX0z4DczONlZ3RG7/iS5Qk9yLLSxJSZ
+L8r4r7IgFK63tZKvJyiWvxNzeTb3ADPnuTEpbGfzMd1zQZMnE5bNEF1Py4ctI8R
YPHRTIlTPrgAYQ8KzDDBM1HZHCaLxcv13lii72VvxwSWLB2rdink4TYUBsW/Vrkf
epzrAPkBV8EbolChhP9f+i5+AHsLSQ3eUhSM8XhNwdIQ5QZG7r+jl0QIr3zmohly
HzEohtCQJxqzoHH8UbYIBSLcSiogvb0GWhcIZAWCc9D9g/F2Y1mWNIq+bfcK7IZs
EwWBum1Tb4qDcN+hNnV0zhTIuKnh11HQtCNhXDPTNcWfY3iUJe4ITcGfwVcju7bp
Y478AF0XTnso7Wk/tk9DpAgBJ6+9dRElPHSpxqqCUS+SHv7Qosfl14Lb9uQDVYXE
FZfCL9tefbsS3Tph5cinoW2Q327YPUkCOULG1d3dkdz8x1JI8vypqnnLMd4DIVWt
YFLWugcd5fO89AIpeJEAEeg0kJcP3AhmhD642MYbLtHmqMOMj4RBqIiIJ8QU6YjC
VrYUQVz78bz4y7ABeNlS/BrDv5J/93KXQaGe39eifzTc/6VlgDpw2Kda7AUmoZig
y/+nJEkbFyeVIdrZx/LAJHHluzB4pvjTDlqvtYHrw1YMsvfLS4vj6ZXBDA232oxh
8+Lt710nF8FTrsRNAZwdEWxk0bFUUNgyBnJfdJOaG23AxRxE/3c29egej/4eRwaX
QYBnQ5ZeUxv2v4XVemQ7OoVlU6BBwBOHomqHAhAol5QEsGyqIkQTeqhnXfAa/PT4
C8ee1GrMyogMO6SsnRxBQRR8qJ1C0vBcCbHmnzzhafuapmdbVVwnUAgJqqrDExKe
lh2dBrSJ2ifRF1YZOq5842zFMog6d5AIs2+OF34+S7FDHQLy3SMjgZwF9ALTmbmf
o+48I3enakEi9PdMe+aDEta923P+1hTpsxr6fWz+cq1htZtSPtS53wItnH2vUnGL
5y+QbBzCjsfjlxc9s5tFBM7EnZE4vo26kqY/G5jJFR+dLxWkQYgtNnVmkdVG8vI1
BTYgok5gWIy+vcW+BL76ABjIN2DP7v+vccuJaI0GdOl+B9586glxFnRLyyoeI23F
NKMTshOlwHxx8A9ueRJ80lsaXrggiozfPRD+j5xASj+r9bo1LXv9kF9FNfva5oDW
hQxPa7zBEH4BWdgO7wS1YzrNwRjOQzI2jgiZee2dFRiFxDNxv1XIKZae2pPC1A18
oqCxm7xdZWeIb9tELJWlm5uARBtFdEH0B7d3rQPW0nl3AsoDs5YYh7c0ou/Yf+au
uAEPC5MWT3ur67JU54pa1OKNPvp8ihcIa0K+ovbt2x4gZyIV2Q/IROovoIQfTu33
iSyKr9i781y8QH7qeOYJJRmw+qUdPmm+KPr9ooophbhmCaqRCRMDTZC5Eoi+fcQ3
dMbQjLUTWFp312gsANxR8Zbzqg05cOyVIRhtbr/LKkasdQ2rmesjTTvC5PZ8yMyA
Bxkh9V5Zwbk9sImE3K2q1pxZdom9i+qdvkZ+byau3mSdSLYo079sUaZhmP2TuTBR
cX1Uf44BlN4y/pu2cSuvB2fFMXYWAagrtB/dOQZIzxh8e6X5eHuBhOGD/AjzMXEr
mO1U/f+w8gi1wTNSGgkGF5CmvTETHUmosowP2G+ghR9TqoNxypqwaWftWmyxaCzA
Na+/7ACYFFU0xP8PWR4aP2w+Tr6/XfwKS6c3NjwBPPUsD+2SvMtUnV6rp9T/bJVt
OgYa7PPNw0g5cIWAiBsQAHjnsk725GnYwSWY+5iiRDtCdjV1yJfmJ3oYgaYdc/xO
5z2LFhFx21QFegmQ11BFpGdtTtboDJEkn9jVz+0hTbSagHgfciHpXlnsPqrOxVsL
CHT5JqnAub4K6ZyVQA0WbBIj8LP7kwmETayJUkFEPF1ogE+IBXIrSppmjmCobeyB
U9wspdYzox3fEU6Vi5pdSgBS5GFyDqkCTz+ICedRSYGGBBpSQAyLRL0Gb2y8wjKZ
chuRuaSKujF27bDpx77eYUi/wUAsdy22gZ1nYgaLTPekrbu729EdcayY7yvLVoKA
B++tHEn+M95FdAs01cyDjdERfNPEpMeIU4m/8LY5vjjahmtFDrRHRPzAPFEw2jiW
hcqEsOknzE9FFS9WXAt+BvhPIgO2CG4LKMYEM+Vjq5Y1d4bde+U4xTx67M+W3cjI
6b4A63XIqllx5USTUvm97EZxBesx5yvGzOcHLv4glpfdvYlOW1VayUXlqlTpjGx8
IVBHNQ6ui6QFyvKFT5doVreSq48K2Zepeq3kEAQVG2axMuPVnVcEOBmYI8cOTEvN
AFfz/JpPNtoqb0TcA9Q8cpfSo2rveKQWGE3195gztRv5LtMTN/bObCaTISwNoVPN
UBqzxeiC5/yv464r9sous2VxZ5bfXTkr8QTGOuv09NsHhvurhk3xowY8oP4ltOMP
/4JNtv9Zv3s1rsdQltFztk3rmbQwd3ozXD4A3ukf2onuAsA2gOXjOXugA0F2B2cS
S8NdAar7xEGnZnHZ3xvhVU10s4T2z/JO1O3PtymqPfO/7x5v0XrIEljHwcFbK01i
AV3L1J5VC+qMnA6vKMEBO8N5zSqut877ZhlQdByZqXQY7iaVsYbmCZh1+2hu4RLY
5HlFczVYaAcEdo1F6UsbCHYmpUhD4PdgwyGZT1EeeHOHO840ML9R4QgXcUIc7TF7
NdNT41og70taJvQsimhfWCzZqSAr2rjcD5/HaSa/fh4BgpGsW5MwXzicdIo//B1V
itwQmx3OKHbklIaoJO2YbHiDfvfLz1HVBAbUDHR38OP16xOkAd0ONdYExuHyVyAl
g9aYjM1TKEb0Qt08kvXIWBcT41GfIaWUrgDxIgV31LBw+lqMCsXHk1hhhOOcQ9X7
JptNDPxNh8VOlFkSV2h8apc4/tdRfloQVGzXTEvR46atGrYNf5bafXU48DqA/NQ1
qyw0FnYwRWUqc7OZ13hQTcAHUnCSu636sNJo+DpZyFSV+Gm2NOfiIXErhy96txKJ
zxiiTFs7uKjUVNwFfl6pplG1eeEGeOfH1cLYfiUBQQ6txvjLXGTXNpbpL4qGg/IE
w7fgNM+abcUUWc9N4KCIsvEvU6K9xqtcUeTNJ+YXMsXPJiGKRUt0wvIBYhmtOaln
IjthimZheIf4h383BSo/+h2Cwlc0mqe9KL0drwhWzZORYMRiPV9GWPr2K261iXAo
BTYBHNoWdF4WjzyZdUi/PTBMrKHURCJS30ProMGpev9YxO9YxKm2HR6JKZH3YsUE
UTHqLyNqAy1xh5h2PEA1xMr3DitbTOJeTpVGd8MBTHgS8VRib53ss3TUmlCO17i6
8+0fHxdZIxbqf630PiA6IkKeOnix9w14vkHt5WRTnJRkSb8QI+HtWL8dXVKRbKSb
xQNDB4yK3YHiLEQVD2n4e+PN1PLViqdRb9scYo2RKfO2zzlGK+6xb8jOkpkk5SPe
BaRqF5AJ+EdRXBlwI3RW6x6bpu6fqpzRNz2pjY6WrGqXa3B0Vi0iOu1FN72zTZ5u
mcN+Iq6uRw9ltVVSqvAW2lagxm82cUawaKf6HhgNtdKl2AAiMdtW+tyosDT/e776
qvO9lNlIaRVgHIWXoRNIdS0mxKGDdIxr+yuQ1P0HQizQLhSavectO6ZlpHaCQ0R4
L2gmOKUXlBsDgKVB+TN7+hXAJhW+EVzy7hm9swI7pEOXmWDMW6QyUVjEsB8toGpx
S8z9vEEkUVCHrEMxDYw8snt3jp++hdGix7xCqfGjqefKvP++neB6LgbBslL2fmnB
LUFFHeEnqs4m4OuLXjs3UpZRNUcRp5qA5B5GpJati8s/wAtxOqOEIBRYyoL0jPeX
+uN9c4M/p1kiX0HrIN9K1lU14GIs9T4M4ut/Ow4J5SIIXWBP1XslPgR6DY7GIZyR
qX+pCAGPs8iEh9Gre85Z0KQlbOsdDZPtlKNEXv5yZKHl/Y/WWW3G11/7ThCt2oGR
fGYlNYnXP0QiyzIU+f9JIhTQ/jiLJXu1TTb/dGIiyVY+/9e7Ijiy9F6A+XyC/IPG
1VEOq1uXLjbz5fqsFiekM/5W1FLz1PeUA5pEgfTbvWk1WE/IB4ELpexJearYRd5y
JaNwCz4FUVPdZfFsKi9N63N5AtWtfE9abTej+ED3m7HBtZg6TyxChHGIQf31tvcV
zTDHciuEbYQxIVnA8oPIxQzBbI98/H4PeG6/j/3HgF/1XorUUDlIO/VB0WSBTk8h
4ArlChnY53SUgKKy9/uDmOh2my8DVm0B/M5qUGMU/W1JSSv8ExqdmcjTAnosZvsk
CvHOXY09r6W7imXHcNSAFNaEjCfm2hzoRBZ7MQGBWNAfKRhClupfPvuJWahUmf1U
4xrSIX/lUX86AjSOcbTJtlgBS/lT6vDlcicfk6/4mgOs99hchTBwQJHqcGQu6VXP
KBkEg4uhbKRaEfwG79FZOLA9RynLq2K/zwTRR+f4RlITyzgkL/76JtKLRZWiS8Zy
MFptU2wf8bNG38b/iO3QtQRPNyWD0RiUvO1az7Wy7212XQ1WMM8CDOhIFqc++xHX
IDbwQotJm07w9mnvZ9nzJm7eC90cOXpG7AiTzImJ5XKHHkmbVCgRYT0x/CtCtGrZ
ugxe0BAQ3SY+HWVu2EK1ddM2c1bw9Bdd4xnsmz8fLaLsKc3UBhmaamdL+Eah9UTk
NiTeIFGhrZIWOmtUcPoM3pa9B8ttKxL8BOs57+BJ7kebWhZvC7kROtYykuXUwjlW
6soSRg3KVg+alT/WwYhCfNjQNtnA3FXk6U+LJybDXI0ZoLnqL/HGsqSbiXnczgsQ
y7uEGyCkNTp/xXOhhcUp4NkEc2ZhhYD/vObHeQRmfRe7qEP/6y/THXN41tjeXe0i
BIVRIaxCCqTEslMIrffxeoEtwjaL77N/Vx7LQeqqCSxo9ICOe6RYW7NVwYzg8rTI
oKJDzUKWogjp+wMFCgDm1rzo5Zk8BKCz7UbOrD2Wd8kAjX5amrvPh6OxdfjSCXxb
gFp6hK7hRgchDN0MzoyhuGSr36nRAt9qNI296t8Xf0REU3dwEni7b54qSbPRFrqX
Iob8mYajYq/6vnZ+aoTxdSeTaQQWEQzZIP1QokpxTpK+HG4Odj5dtx2apPnU6igF
FzSBVXOfUMO8Am5b/EPoXsFltG/2+Ueg1LwthLBbM+ZLkIPJ6nqYmsLPz6xa8HeY
mJePoZKwRBTmIqowbf5GeymiffyH+auyy3+gqsdjYqUNLkGh0C7//UEPtrPATdrC
adlNkwTo/cvW96OTan2xuNF3BoLOf7L9oHT7R8FGN4pErAqooGUih98+8DKy+9Ao
B92OQwOgKTIZrpqQB4mesEioLcgEIHjas4HxRI43BHNx+Pp7Ao8ftTHWxaptNGlc
IElF94H9PhNhfRpicEUIRp+k08R77fRtpBm3PAIdU2QBrdoslXEC9Ff4VsjdVgF9
5SU6Lf5CGRdXVRJySSnefQdlE6TDd4Y9r3nHquq3Jd2VR03VnluRutuuvKP/1FsW
MWuxcUpi9SezZPFhtQeiEyoz/9g99BdgQhCp8ShXaLGaJjPWJZtoYHP2tPo/Awsv
C+vQ1TYITTyozmNOTEE689DFzyPQ5jmpzoW+5W95RAJSE2g8J07hdhgoY/O1oKka
HYE6lKPBgFUjLKcBtpLXfqTLeIxY3LKp+b1lDynq81NOaVoenmnT5c+89eAfIg4M
UHQd7O9D0F35fReWTqmRt/jLADB+wYXsRroV1seYTXVgzGkB0pKfb4ZAq38zlFY8
3+BdUmNWAshW5c5pnv9opI2bjHLepM0mcycXEL1K5Q5mLtMRLEzJMG3j9DnBGRzn
yqGeKrkf4FVbcYLiE3A1GwBGuiYqIyM5U6FMSn0O0nSzqi3Fj6mJI5no6p3zco+T
RyCLbDkxR3v3KibAfpe53a4BwjuK9oh9W8FOAVV3fyj1SVekC/rDjBnYQ51deRAT
Qlj5ZDsRyxahnjDSgFPgRCbIFyv2H5gZO/2eYIUULautQmJ9OfVLD0v0wXmMX24G
iLno4XFBDRwR1tqQkwgeb+D0st/WqQ2EQO3a/P8BQBeHD4vahpS3eFf0kImFUlcc
nOCYgR71n4AXx1KnBHf9cKJdM+9qBP6GgLIoVwt+J0i6uOfiQauggaJcfogJNTKN
yoesPxoDGp39KRcVUpjER1wVjsOncnxej0VL+NL22KZlGhzb1AvfZXajVE8wQt3e
hIrxVltIEUEqdOdzEpiLy8cUQtzNfTH21NQEhYTNuECT3ViLpc2bvMVrgZ3+TkA2
PkU6Tvw14SXW1RJum7hG/hxhihsyBNcuSzGi07qmVTbr192iggNjM0GzeJytIslb
Roi5DHlaFUtOsyKZ2pLsqNZVM/7SAJQ6otY4dDjfF539Chgx7aKgmNEOIK++OII4
cPBolUyyoZReZGgcmVu6hgMY63EAvHe4OUxEQrxNZHFLWBI7f39zy6STVKDlvzL3
oErsToUuoqY1S7ixq7oMLL1zvQctmk+BZTFrShzobTr/P3rXgiOajwl9gq96vLzH
hJnryH4mv9a1onbJH18xbnBsLF4jYsCDtY4GTqTlB8ARcIhLoo1hn1c53GO0buML
wNCf3LpqkQzLUv/hDgurCE0wPh9B9+fw0OW7ywxjU9r7f2c8Xrw8fvxCuHMbqlg8
RaROw292dp7yOIJ8rgDpqKnpXFTH76LAHh4xIUvkwg8hMgSo6usax9QIwz6Q2lZz
QEIRQWLQMcxQBiKGdZ39Fu/O+Dt2MmrNsUs37Ojk/4sMq53fvgpi2QirIojSSzww
o+nrVIDKWiIAUdZAK2kPjlvXHiUT4gxSmRnXQNiSlMYeMhxNDceq2LMGPo9OPJmc
ptL80Mo070ifL9/q6jVWFABZbdoo2QIcDer+Z04R5Eegfx87krr0AlmUMNEd+/pI
h92L7Ly33tNv5ALPbEstKfzdThZbB7HlIZ5HSrV0KrHo5p5snqoiDc2EAh5TtzPi
AqsWUrGO2qyTqSpD9vldhRAfH9PDDL3G+1ToHEwMdWjLXtCtBIuBMCzWb8kQUZb0
s6rJxf+oFn9M5KpEnZQhixT4unb5m718YdCzRm0yp+banR4Nj4H301tFSENj2kVH
W6sqxuVHE7uoKzdTlz/kIj7Nc2KdR0X43H8qhPL4tMWqyxgXwXxjHjNLiysyWeF1
PF0NlyN0IVbZ6kMvwakXo9sjMvoEQ3p8I0dWYj8+LZ4suFHq0BxuBmGKuvnS2MR8
aefn0osSWYSNb/1DZU4Hclna3TITZiDjkuekK3ySvV7Csz5s+spjaGvSBmczV71r
oEF6fqNWCoj1kaSuzA6chBpcwS75DrRax6nD+f/iVfLKJGqdSmqNIsFJ6FBBPsSk
xGb3UdMH/bblyez3unj5tJLTOPJIYP6z8dL2ZMyRqO8qTkeevuKQ99A32H/ZqZUb
cbCHLCsun1qH9Eg+IjYMvrmS0CYIY6FHwKDG8GyyrGp/ZRH7zTgQM7uMInSirmOV
MeegwtMeArhiMdaMY+thjJMPRRXo6kGoK2ySHYSIFEcDk34AmmibvZU+WUolEtIa
LtVgwL4hAWHyqup46TrzcYhB8kdV8JDQfFfGvYoURoDXPRMOtBDWg3q+uStRNUiZ
SPOp6hx3Ds+oSdE+9g/K6wmi99z8oaFdF5GP3mqnDXaTl6xfYF/7CQQP6W6GRbE1
yrmZYlf1mxhJn2eNZzHtAvPQSD5z2v0wI4pq7UxfrvCtkkt5hC7L+cEZZPceJQZo
4+OJwkfPPucU276DoRRmgQHkom21svtcp2jsZ7RjH5GcIdnf+HrOVoL57XAMykW+
mtleLQWu53EcUzBsPJvkKccSVEq1BYZ+KjV8d0dW/QRR3rr1THs1LN4x6VPcYSib
0b6BjQs+tSBGLfVHKQb57MKEkN9NE2TBh/BAEQR35XkU5L9nWjP2Q2XyTAtV86JB
ukNgvhjeJSDrQgVhCvMFV8bT2t82iOXvI2Mc2if2VS9C4W2UjssKMCUTb6oKbj9J
FPAxeFzRBFhyCU6W6wP/8bx7o1qaE0SOV1WjSsGTAyASxuV5audExgsZb2L5b0oZ
ChN9GrJecgjfVofaCT55HvGEbhizGCnass2MbCsM3OmT1MzRZZM6xmfZhU2wLNhf
kOJU7kgNBxjre1r5KdwkAogyw2oK42Tpz3OFaCVyM91pzLi/tsZlFAb3+Ji6cIiX
YVqeYYfjtKdpzHuip60NccL6/PiNifbT1wY9YP0QodD0uACOEvFbWtYscxnral/A
SAgCyX81Q4IUXyi3fGHqtoV8FhRcA6jJWz/foycA+5Y3yOa5ZgaYnU+wMddsD4d3
20QP4eiwhhkAaogG1Jn7SGITJJOhhCshPV5EqNmL+ibuKcVQyzrVTqpql1ES/rIl
Xzm8LGHh+wK9rQGphF1Jms/ERNeM9v4IqqwD6LRL6b/9mwchnFZ+8tYbWmnBE/7o
yqWjmw06ZamWAhYU9F2wzUDnWBhreTWy/QpIl/D7HKwv0SARZPGbP1Q3roSRerjj
C5kfHdylTB6x0oCTi/LGtTU0dwjPidOTc8zXVSc1Sq/s5HHcL4+BK8ztr7ds3J3L
yNTT7Fb0vvQKx/IkIKZWb0QvkrHQRbwJjEJaZOiicD1t7NblpX0XzFqTZTzOY5Jj
jbw94d+Y7EFQjZqc2dDFkBA9WK3ybNKnEsqqTICMxMpLEKkjIzkAQDp6wMAwd48S
S/u403hJ6k7ygLxcRfc+fnfB39Fw1Dt0PuO2M3Mw7pMtnjYwMFUjeCjJQHEcmIVc
FBd55bUa+mQmgfB6WBfBN7ry1Zha0orlOnU3+EIJ4Jq/yEfHTSXyiUotLCyxLQ1w
ZJSg19Td0c+55W8rYd+3RhnSXcpz/5JIiseBTZquv8nbCC7IPvOHjfWSMTDTXIQ/
9ISdz/tnnghAcVVYv6l+emHxB/eZcSzXwBAMbazvz0Rw3+CNvKFNJzcdjgpbxRxY
EyuT+xX+9seXZxpYXWw9bwtiC2zZTArQfSGvG6hWKkYe94ruhcGet0+rB6GRSn8/
jlmBE5DWkxt6ohzpYjPYbhNl5gkdyLEo8GsMCbW9SYWUpjBhdB7AIjj+V5Xmw9M1
zK3h7uRPR4/L3Y9eN0DeTmtKhd7X/AUPB4mxqHl5RqJUPssqwh2hIGSz55HdUWu0
gdB1lwKpu3oPl6XQ7rAhz/jAxp5keRBHJYwLgXWSx7qla/5SBbspxXZ1K6vgDyx/
hKGCDzuNXAomT/67p1sZfJNI2XUBgCFkuvYZISKkUePP8uaFtShXZz5KbhRSeLfL
/6ac4da0iQy1m/uqpKzGXYJ35Twz2eMxU7S5m8ia/tSa9ev7uya5sUDKY8OXoCEC
BfozFl4ZILsF183AbXNWsXZRsfJUUOf7pXgprwIoYGCbxTPyVa7/rNncKrvL4bQt
gKYqrDKDn7jIF5mQmNenTlc084CPXxBXxgU0fmQjTQr8gO6qLiNQR/Z9Yh2KgOuE
IOqLHUskoEs1L0m4Phqj4TrBXd7LC0vcIhvaQuZvOIhWhnQYkaM10MHZiLZu1Irs
zNCjleEBKOFSK05FC36vpYP2E0+Um+6eFC7oZlIOEq0U2Aiikvm3n5kxjgPEgoqv
kG8baKcGP2rH8drQNOFsLGC9FagDOaj2+NZpjzeP1Zr999hJWRD+na6fFx7RxbRQ
ZxtBguUhReAte0dE2gqa6qBExgfppHcjGe6NAeMor6Zv0OYBr11EHPuqr780L4q4
WsI7MbPP3+VV4LJYeglIOjswFTjI8QvlBhUJfABQLumCevgH+D4lE5hGdxNoZ4+r
0xKwCoJu+5fAIVV0o1414SaFekjQJ9srtZn1+Ef523i4e/n6yVfPo9gTf0iVzT1Q
AlxNKM1G4eEi/9H04ABpXaScIoQh6r+bIY/zj4pi/dIlRahdI0+YD58L/Y7C51D8
piJ3pqeDkmj/tOZQdZOMXAOySnNTdiYKQ/TirmuA+3uj5mVHBA0y9DxevUsdD8eM
4l1FR7YU0AoM0abW1bIY6sxgS8WmtOyoVKggT22XG/kI51oGUR29kySlUgC55ZLo
YpZtUvhf5gVtzA3RQavHXWLtNRxlWSKHsrkTq45KNwFniDX3N7wUlyIZSaYFnzbh
JeoAim0/4kxwkq3F6FCp4v6WRq1ndv58UrKnVx0P2g6oAO1MQOfOtfhPondijckT
DYIw9iQX3NpyAl5J1siKKg9u7PMp39n7BnhsMTuUOdMb5n5X/kFW8ci0uirXyld3
OHgIVQkCYj+wTjdwzWJBuIYQsCa+ib4adAGLBpCH61kG/Vp9hY51SI0fjjfY3eZw
jhergIYDITOnR7+JONhb445DR/ipq//Xum/k2g7FaI2Q98f78GcsH7XVAZY0W8Vc
+5aNGvU3CBRhyZ2mDMOjuaGNjvZ55IUTEuVAkPdSsOPz+EmiROR+xXgYDpaDjW65
VE4eIT4tbHdE6SN8yj5Z0lyema3cYVTVFAqxsoDioyiAsG6HTgHDl3QlzjoX29RZ
VD5M382Jyd9CW1njw5SsLd1SxhJU6psAhzICKNQsKxc+dDYcFr72lJyx+5IyTi5d
7vzzdX/eiCJIPvZd8HzOkZt/E+Ll26qePRD18DAf3Mgp2c/w0x6SZDDJCnV5ndbC
bD1QiI6WM236+7j2yO8ZFOqMz3/RbOnQaHkcsNo3D1uWSMGK06OCCYY72kpbZ9cx
A1K3wNLKVxbsO2f/DqgHn56/5CpVLpL5ghVNZMbxybr698JwFLwB5IuPKrbZHAyk
m3jbY0Vw8wLe9Q3tix8VIYpn83x+cJjwpmH2J0bf/9W6m4rvbqk4+gpreQLDFJ6e
OPT5LObPS+nsEn3ZZeh5oQfnbzsuhit/n42cNLty0hV+lFse+ABEDKsONCJl9O6a
EFaIe8zOceB9SfxM2O96LIwjpx/1/YIsqXm62vjtvftcy1U/60d+PML7UNKf0U5k
kLqvKvbm74MKtm0uw7DN/2w+/XxWqU1tgX5yz4xBUsb1tt5m03ZBoLRf3XF95fNV
kWXmFQaTV+oEMj1kkalVXTwqWzYbHPEqs0JsN8yKDZt6rTM7bn8yz+0zIhImhFKv
tn0nPKd56PnATefDmIJJBEjCPLXgi3pHuGbezKtQL6sXHVDuYZoyNgk8JfbSubNA
Gf3zSxSuSIi3Cii0w19BtPwDhwc2cu+KwgI8ejGtFLdbxzNCyr9DpPTwsB0G9O1u
KqCb4QTQSvIcdq3vLhseE1Tk2FcwwZ2Ydmv17u5wX/GUkDYeShj72WeEJjTDqwaa
i/Dr+FTxdBJcSMt8E+kapbeA7l0EbTHw7DXoVSr9EBXyTraSwVwz8UYWPXbh0W8m
2mbGDAuwdqWCXFUQQiJ8xNnOxXK65A1ToSqb2c9sFNZAa+YNVSfO5+TvQnru4X+g
4cG+UwZpjQ75wcHtsul7WIITflcNVgQG47kRm3ne1+BWBaaFLTkdE9lH3wMuCTx+
ZH/Qk/nWgrEzZEvV+xpthZiUrZZT694zkUvtig6jYpJSHer6OQyX/4hfGhTi9RCl
YaGhAwWDkd/h/Pa7VCwa3BE02aaoWuoODj6pvzZS1va88FkPOL9qNCs3jniXkVJB
9tajVgTbZC8XmVIPz3QQpoqBedScLQKmXt/29grs5jp9NsMHCtCQlYjLMlE2eto6
DgF+JDzZ673aDYTtqCRYdzNr/qZunPZSMSe81iTWBkbpsaFljbGy2IizbMv2EbxR
n6f2tmCCup9jQ7wAVW0oKkck2FKPfO3b4183f8+QnTJ9tIHDBFxrHytnOfztom9O
KDFaT5fXjrNaSpwGKRQZsnzaNR/AbNuigsnhlpD18ulevv9zcTTSle3Vz+IyXrmC
GXUIKq/ytQZ8rWongQzW1Pflj08dmyWVY5ohBpBX8QYST9GD3bjGmy972EfGCZ4a
SD5c6HgZ1Vb9W1b8J+POKzToxeHo6NH9yE/tVzKa9JWPN6iip8vabFZa07B/yP/k
M8XYIl7zEND/LYYCxU4JL8AH9P4d/HOy8h2dSeaGR0yIarv6+7xHUIWe+5O6MJ1w
Pjod9QGq163wL8MZPlSXfF4MeHK3dHxtsJK/9JlMYn5BbPkg5LXIDtScUK5VlulM
L2SDZi73ASDpaWyyFJ/m6aI7KVn4WnQYZmybQXH1NYNesAEvozRv0/YuX1Jd2xXH
vY6if1BRljQqldmBAKNl7526E4CD1LpdYmKmJNbArz5ZfxGQx4VFD5hgPEiafesp
/won7ENCPvDYdEiKRP+BmESEBlOp/p82pFPFiKPjK92+eM6a0YaTLdj8y32LAYis
SFYy+mwN3RjcW8hGIIhbXiijGfcX1jU415KF1eBckZjbxQJ5iqTCRhaLOogX8eqD
lMFx3FTNNk3esbohOhJaUz4gIDkrROcv29osVKb1qVfEKdHR3px0yF6bxuxeWnAJ
Xwh6S4zKyI5ZppzLQAtPFC9l0wkUM4iteoepoADYJOC5l7QH4Y1iXXcpE+QYYs21
6bShOgzXCr/JCQ8nktjkYk+KXZE9PD8HkPYgbFlSG5LqYMgCkKrl3JsB2vQITYlS
FQBkwxI+bprRJ1FOQLuvtdv/cbCeKLUeRjU9/JHT/52pBUsCc9Pr6YiJoe8ujUAX
VNuyJSZ7yAupncpinwmNJ+k0ksjz8nvsQs3ahZbji62HPWd1ZhX7jEfnpUokslHb
e0/L+01yOzM5fERPH9MxkMFrPQP9pckzXSJSXea5S4hbiaG+mTsSwA0GYiKMXTCg
YaL7TUupOWq+cvz8IVpfBIb8S/qB0wUA1C4LxL7JzPMQAy4aekohsTih2ftOd2BG
WCu6Bd+ReMldgvjpqOXJxe6ZMMp73a+7js0hzZBMZJTjiK2x174QZ1s6bJvfhamV
CohHm0kpgBAVMroHLmtlSZPLAalJa5ikciKANax09/1yWEFj21BwwUONzLGwQ6G+
5YR2LVU4Jw/66OeRWXzkN79a2/eBCTLyQjiGlpkvjPEHmZCbHCm8n3vr9L0+K6r7
ksLzQUET20esCzrLgV8cf/7uScRXTsk2XxNqg72R2byk4xWGI5gJqxhaJrnyoPPb
UybMk+4sjclG6jdHLnDr/bAIbMPOhnBFhlnJ3a4MScZ55Y/1PkG6mDt0S6SUVIaN
Qcz8Xn1sDMRIdeT6m/NHWRC9J4gnawAxq1mZbr6SHCp9MMGWsFAVgfqLqcXPdEk/
Ial0rxveoTYD96jXXcs2p7sUGwo6SikCGPVbo/9wDQAvg8h3wh+C2TCq/t4We3Bv
RsnHk8jIPgjCJ4+4cl0pyuAQeqXLcZ9h+hcGdaG3GU0gPAiXXjTgX6VQoqAHh5Co
MvxhvcpJs4qntpRRE4k/ZDOyTZmcugR/xD6NdqPvxYdcC3Mo1Ysf/wHd/0kDys9m
KmyFp1oEee5dioFIhipYHnGKrXammYw1apgG8NBg04bmuqWeL3aGSPanMFKw5v1k
6zUjAXMMfGZgcMPVyRuozJN40Ib01RYWvxFmpy1vLV9QdZDMiylSP52Hmtihbb40
FN7MobR5M6ZUfg3UautLdnE7mMDA7E2BLialzJoSFjWnHc+FxxzmLdz+wOtTDkWK
c9wKtIRk3k/pzYds3svpFAWnWA35v7dgkEpqCVbk80dsgHePEH/7iSiR0ww2fq0N
Su+h5nRAXi28JzVNTp1uD9MeS4brQdX2yp7TxUIGOmZuoTKUufmQ3ZNoiYJ+GMtj
Ei/V9SnB3Tbya5JbjTfLYTNOPBMc27UDCLQCHyryhEl0v51rQpe4RnLnqbFeVRR/
gQ1s7SjNgBHFMT5mhFlhvL7mAAAg70p/u61qtpdECfQxb5krxjdBq2r1iPIhut4x
uEISzQt5iIRxcRObXuLdsR0O6qRds/w/DpWcNYjbKzd6CwwdsNl+xDxkzchpG7/w
HT2EXzhgrGxxfaN09YgrZKBxH4QARdWlUndedLXmrwTa8Q+Nky5c+oL0ELdl7o8G
gh83cOE71h+I6Ww20CKFSk+MvXDOLm3hl1Iv4y+EpJu95KP3Owk8Q4+A7zy3sXCG
9FbHFrVtSNDG0NOnzrpyFHffHcMPcGYISMGtsWVFObJX5llZeBM0JjaUG+nBw+zT
axz19bOHKR1/g9PPactoM+dRvLvwhbSZX9X9BPfYd20j8j50QDInlpiS2W1Fsjyw
DHXiT1vhrZfa08WqY7ZM1MvfOmCa+Nwf5PMyYtsh4TfSrE/ywEjliyW7OSn43r7j
OqUSAyXlNNp7lauMfkyUzf6T8cI12dTeh0sZt+opAE4SsMKD3t/PPLURIBSwSTWj
Qp7zUkof0FigwFQCggVYWo+Bos9WtCRxfDVCRfw52VkugqYGN8+/RpcXja5mc1es
URPgvdxwdOqjqBHLbmzuuul7uQ6Gbb69UrpKygeWimsCJ2Lme3bVVqpPxxV8w8UI
FYWPBfZCH7pcBPVDVC48H8wFJAbr69gZImWz2GcuFQx7vG11b/CnPzxzowemKVon
sQX/AQcTJJvO9eL2iFZTfRcImVtakSRLiw4V73LJnrm2mGtoyYW/WWPCz4XK84aO
upUVIRUc1kEf36BMF5YujzmwzKqs0Pe7QRgwAvnygU5ovonTp1cwpZ/U0deylPzO
TLdzxXfK36uiQ4RGyD915Ol6XkO7Zqc84/WRHhJVB2sp9Z9UpuRBvrbDQEdjGOVQ
ciy38C74C5wJPOr+TNRlozILPjr01dD7J0jeckhODPHLQ2TV0SI7DCsXd6f8YH/8
6HMVzk5tsaCzf9dk5q+stDbufsIZd7VZPJSergJv8I9fusHIg80+Q8VnSPbVGt9U
vhlIe7wZ0Qd93Hd5DqqaZmKDkpIyuAirSwINhr6Lube3/AySAoamfaU4wNKyTCrI
6HLPzqQvU6it/mQBTOir1lj3wMuR+19ECSFZjqg3ksboLZhLsTPBiBgIs1rnS5Ml
hNzRGmYpL37Dg8aZguOOr1YrjHNXCdTlsiqyTQJLIqxMa36I83nu3W2WvhZ3xOPZ
Z93fOBM/619S/pi5hmlZwIH3L9YaDBcgGOpVqiknbrP4PO3+xLXxQ0Xi10EyO4Ht
wFu3rpajVO7QtM60q0YJBwCWBV6vqVLZDajB1DGKrMI8GkOVoM04ZeD54+kYxkVQ
uGhckQlThGBfe5IqtH1Hi4WaeT50DorIbFxaIytEYESvrF5PyDSJ5PTgZ40hhtOo
Ld7hdu3TSo6Pdffypbj8873ZnH6T2oY7yFR2N1Qq5FUELawiWIPXBM5wBlZMV4Jz
ExFm1f9ZyHaQOeo35T5kry8upVtJGHgB5DKfHEIGjozc3vFYxAw6FhnJqp16ndXT
2g8BysBjNtZAJg4yPOfPVUfAJHorJz3Ly+Oc9ErRp5r9K0Pu1sPwt7VhtTHFr/1j
A42ZMeDxk9e+5kAQifcy9VwhvUMzqjhF4kj7lfQpqpEUgVTz9jeT1o2Tw+2/MRyx
QiR7zVQlycF/8XEdmw1LsePp2/AccvdD0IxWwnkCYq022HMuldZWi6pb9eq/NSxh
qqWSqkYsDMOn8O0LGDjhm0AG0RNcactllEIIgmZ7VKswIg6bXyWBx86djBNVKogt
Nu4WH6t/iDBbKgpijcUKKZyib9IKvbYCj1sa5FS35kJj72dLzDqi/uKQ38hWqK+W
a6x0GvWLCzHq8qt6ed9Vq5jqHl3re/Px/e6zS3aPyaf2k6H1Vl/LT/ojjk6x3GIa
FNJwNkbyaj+I8//91lexZUWjOFFk2IW2uIiz9pt7stCWFGXaUDTbhGxGdpaLqzG3
g5LVx5qTEBdFq9RPZi5632wKvXnFkH07CCX/cNCWtbOSYmOIqmLMyVtOy2BJE9oZ
gWSRgc7E97m5N5TfWsq3kJLmMsi7BaKaZXavxMFyGztDohnfd/LIJJhd478kmnK5
iyjP0lj183JsvXgI/k5zeQ+83dXaFd3408SsVWHbASePFFGcmqFpFDI6oCLjJd/7
9iFbmccDPZ+KN/5P3UhblPqairQnX6JuLfeRN6anoiRx9SLxuiHG+/PkEvmBrJ+h
tnjWJvjASJwP88JO30u9/BGbQUi16bc2cXAxduQ0VE55T3G0hB8tvlZRd+SrZAXu
g5a01LnCudNcKT2aeJZwoR3Z2Jhb/P8Q1KxqQ9lX8BTWldqsYCwb6D66WetyHw+7
P9kh2lZYxkaiKr6cSxAf9tnlj8e+kp60tUOrIcPKhCWIVsQpM9wKBcpEXeEPSEVW
qfh2a4w6DIFX/c3yXSkf6EG8nE8fqWIv+B7WVZEZVsFsFqXugc5aF8yLY3cIlfHF
oD6pzRRITfUO0bhKuCDJWoSjkYVUAmdR4BifgWUWUewD7EHN0Wapnp29v+f+2k6J
2G8ISfJp1/YYeWSoiE4NRQ5uL6sbpYgV9rLU2wX6TTFvf5lFhYe7hSt4PL197DqF
aLhTH503/7JL7OWlh1MiptSQsHaH0kBXoyXpC0H4TylkCR3njCQ7ZlgMhfUD7XO/
SfrHmL5paQvOV2cCSHej49ysWdO685bmz4yUgV8ge3c1gyg6DrdEWKBHrpkNCtg+
l0bXui54rdfuTMppBwuZhNDylKCsBilhpxN1cysvEmqT5j+BuT2CQSHL6pqgWRLp
AmzYR9NSeuQ+Q3wWTng6EN+PGxONrx+Ab5s4rnD6jfmvi7tpUyrlQ+fTB89eiGq2
SVLjKb3DymWLrxWLXa1UkHED8a9nRw9jHbefGDF4AUiFC0SUojwG8lPvEK56jK12
LgqGQklcJR4bkHDMc4+14KeqEIbis42UOl3VsUyEMABCeOWaO082TeOW2mCloXFU
ZC2uPrN9NJBHwb/mZGmqyD1HzfUauKl2ZqwBtnFr89ffBI84rFDjABPcvCJyS0s3
8DV26q5uW7EkPcWXU+DehaVWYcCd4vuyHELqz1+krezUnG3F7Qjh73gge+BMoI3R
iCcHt9c23Sr5w/2iLhocxWDs8wxkudeMS3w1jetkR7Zsk6AGfXkihhLo+ARKneZb
41uhSsAAZ+82lSfJqopJ97i28ia7sWBhMUMrLr4RYjJviZtVNzwWT9S5Ran1J5dl
EwJ+54bsXJ2Hp5X5eWtP51+IC/0hL4wimzjXskCysWhZ4SJtcOMNy8LO8Mi4egEq
UK7avL4XILNMITflwief0aRVid7w/V/nuVS3Z1bDjm9UtzG5BgKHrij8NObvEFFV
8kNe3LeOmf1sBMq7oHEmzdvS/KuqemGM5F+XCZgLWnT0r6p8dAVH00+4Wd4/kQYC
bVqbcyAAeczp/+YVRR/lFII2SbfY0PeGJaE+36YWJQ/XXnjtAri1n/RWOsZbEbwp
ncTCmRjDmboAfG6zjWC6GpQeQpDvWCzGBJ35lwZ3qzmBZ3fc564jJD2pivQJMLmf
DOg66fP/hDmFzEtO6/Lr7DREkFQJT1d9GtNPSFX77q9EWW6sLGhR6sSpGUPfrX/l
7dac19C4uiTZ052bajKq/Or1KBHkypq7T1IubiF3WI9/xhqE6AdOjcH0r2w/Hi9t
c/KFQdiAp4Znn2ja+GxDCcljplw93D5xZYS3N3LdkX2ONms8rgiM1BfL9QHcI68x
tFEzp+W31MUPGrq1tNRVQ8ckh78RQklVJFQeO0XaCLrwxvO198PW6YDshkKkBNcC
Dsdvb/THpc4FosSacTCQwir30p6EwtOO/CmCKL5I6IGWdmjJ1lMSRdoschzGbL4r
Ng8ZAwL3S+dKPnovK027Guynpm/xrc6MnZNXmyioOTuFdXIEILCo2/zdxPinInP/
ftQzGxkW9B1HbKuYUY7cHfh4N5eNOqV3AQe8zb+ufPoyJFeIOg1asGl6tkr6Vc9c
mklM3ieC5iikbTzukVCoRc3Sh83iSaH9b/BzHoI1+xR+vcAA+G5xAX/nq6zLaQkM
whOZwEq8B4yIwwKrb1hKoC3rXz76C4lcUHTFRdNsxlqShsDwpTN6ALtj1ekf0qou
TPO5cLAsnpTaL7b5gNiFs0jGXaieroM2Cu7kbMEjNlvl4VbmJYK0j7L2ZS0dlpnZ
+nSuN4v3WRCVB1sNJPVvUCLQx1IOGiZaX7hSb581+YexZ4dsozau8AmV+WpyiOr0
yrIlaL5Oqs8hsgBRHy349WeMbCB63DTSERNjK267L5RuHWS7RSfjaLuVwNCVM9iw
ZEC0lxnwDYOFpIXgpL/ZrOpogu372+drleJT736JRs/FaV5hUvR91426yFR+7WoQ
m+6v8soJHWDIXw4qlTEoiXLlMrhkIEIb1y2HaYJD4es8gndw3U3fGhiwKvqKwZn3
NMkRbvjDMnoh7q8TCAZlDWXUuWlQZC44+6aOEeyWdkfiDq/yiXpf41aeZw6VjphP
fuyS3Pjux2b58e/jBVjIFkLQmrM73tq1pc6NeDa2l66X3AYVEZFgWIfSypMagBG4
LXQ5xd3lXUkX8+L80NJP80aaa5wAyhL/TleCXKVpP3zbZsDeYCyngNoO8+7nkWQX
ePNhEFRxYfrdbsSwgwfEPTIRjQ4mmKwyJmn+syzNmPcdLkyX6iHfkGZnOKDxWRAc
iVKsFhaHONuLd5JUV+DrmJVBkzx811Y4ZSnlKb5oSkQbsoPDhhegiasJGOjIFFVw
OQnMtuT1TCLlrv0hq+mHWryBfS5C1w0kF7yEpKzFjgi6sHSTlq8oro/2pqPRPMtI
wZvuD1Xx63gu5ajkDuWv09r861mCaXxrC6grT5MAVYuPHeP1QmYDt2IHdIitqM7R
FKYet1yPwAp7hGHMToCLLjupQLK7QbXip+GmD4izI0a7Erl7IW/4c+mxgKfGJDhS
kg8JiDDZxvGNrWAxrh/DTWxWW6iN403YCiVTX80k+h3t92YMc4yMLTdZxoP+4u/z
DdcGd0S6jc8VSl6nXgPRspZa/SyeBLPpI7fu+B2a/PNdVB3ksNi5LrWzitU7akAS
sgmJY4QeU1uMWQ8fW4aGUf/eHVGuZ5cCmAVzQq+4yifsA7qOVIiXV6+MSh9K1mAA
IxDe9pMWKmaFEb6z3fRsPYtffHLiBWMNqp/FNmLF9+L1HCS1w9BJzeXgoFvypaGG
QWDO+nD5v6qu0Cqkbf1ZaBJLCuG2IUC3uHoW61B/LL6TPFXecyfBc3dLDPkS1jRr
kPQRLA7Impsyur9F+mlOFApryqxqJKm2uwqQINSXOiTRwDAgsdgXdiFp1SX5lqbx
LgagJtYH5UeArp4r51Fd/IolVdl87ZiHxHcjgknWme3Jcb6YWhXCRISLNSGgMV8i
1/btPIOUwru+gcU2NmV5rogvXwSAlVGhKmgFfoeaPW3/shJmcMnnxqQ1giKqbZKt
IB40kW1XXNop4ooi+iidqDIUXzBdeb6aEHOmGQO7/Xz1sCNboHO0tadb1Y1IfGuE
8lVnsSXxf64fjk6x/Kl4zn/bVFlIgc+69cUfKB63iL7NS5nos9lMSoFokpvrWiAJ
rxFMVLBpfeWBtYkvLT54pp7X7pgstjw0JXJyRkCR6yhrfQy9+iTO7SxuiM0kDUaN
60I8+xzHPk5t9dNuQCc+VmbY2FbDUc5IKJJ2PR584usMx1bF3bHbpMG7TES6qmF/
d8bFFZHpN/aGXKLGJ0BDhkynmrkN4HOBgPsc20S5PAuYfc9nZ+ea9vfPQyC1aMeX
nTD3jUtv290XII7PuYizGTo0UJFt+1YdJgZKirnH0R2tCPU/eZSA9A0UqX0p659B
lq+S143oiZMxKZyM56xx8Mu2MnkFcw4BEAdIZylzEZwaukOaYd2yF8J4uURv0NHT
ID2qT7U043dpDpckGQEnotpZdMIjjKrfRrntVkkedAL/6Lioh5vnXNLi37jguROW
BbJEnMrw+h/viZsaTnbBke1aa/ElPPp+uZdl6g/fEa9lss99mGGno3bHOHdrwVSJ
4CD2HvDfvGIavgR6CFiGRoIzkN8YyeV3fhvOcC+PKf/MOExIDuQEXmI/XhVOklys
lCHgoEKHrHhCg3WyvbDI5xRPvIJQhEj3B1coQt1Hj0wCagUkVHJSxAj04DVRV93C
WaBxXxuUOeJym1uTvu3pop3LAvJskvSBPeGgzCoRC4llbKt9MxE7tDGhe+GbbDv1
rZmzK89GKLUk7lyHiyrMnyqRkdZz3lxQ1a/1dAPjVyQ+khq7ApJw1QgnAUnNjEzi
ykqvpO6Px3QtiuIm1Rs/ZEPyqfZ5fOXlp5LTO+jyBMSR8ire9xQx0k9rwq0Leokf
2BzpsYGnYOBQIHtuJmc1UvZhAopNftRB2P+Pe824tTGvMWz9X6qHdQzxzTpBowzj
ANdpH8GIXQo5rysIP3XqiuNI5gZQRLEpsdYK9E9+lLQBlEIiE0Xv+zY6AqrXi7+m
2eVh7RImNF5SLvA6lybynQLRrzkFvvb7y/Kz25lRxhwiStlwZoN9jkDm+UELTJVD
WDwc664z65/ZjgpkcYnxw2c10/9462KCYVm9Ns4EmguMd8jhxeihHbG7vhYpnjtA
toBsggL7w9xf6HozOf+RNPgF+/YoEvffTfwam6pDaBIgQm7e8mgjZ1VZ2VveXtV2
i1j0dek8PujMecgEpxdiV34qrWlJyceqSdr8Or4oEowk1PXcui53l9w1h+D+dIRL
Rq3pXR4nxAYqPpM03eIezfnBYSAHuDG5IH4XvLQikBTLF08xMZROrW3CEut1leTC
XrlPXYRI54yM9MOAMvh7NagwKaq3p0W9OSFIfi6WvgfpoQOTs34wQekn+USK0jHf
cnRGfvxzi6mHpX0Wq7OWhiPO/XQlLZJRBqfg3VIDnbeVHsMpX0C51e9yB79ntppl
CptQ2dF85uG19wcowu7+rCurQH/vkaNlT1V/TBqXKVkXsOs0lRLGtwfVlsInWdBD
/3wNddlngyt8r1fuN70XBzQfc3xiwtHIATN9de0xD/lUecRjsaB82lra83e3umKj
+gOfbb/SUi2TNGojMiowN6dJ0mYRmIhoBtj2r9saRDg35AKNV3YTHZ3SUY5EG00p
Tw/U1jus3JX3NxNp80/tHIwt32J+Q1W+A/GhdDgQWckgO2wbsnkyWE7tMc/dnDSQ
/XrxFiXVVkwq1/f6W/l0h3UiAwWIVoKw4K3lAjLlK0vDCYzHGHq6aIgCCRdy8v13
MiYGZDXNZ8OtDLmnO1QsF1S7nUy9G2h9QjyjJc2fYAkRVfKMTCIKxKyrD99qUsbJ
8XuCmDfcgSaI8sVZgEmn5PKOOuHaQY7Q8T23LD3ARMy2SwNzJ6EgicxZ3QquZSA9
PalZHOqdi/qcjr7FfV9+SG30iDVDGletDrJ789dOG7SaTmy+lrTrlkfF+pA3/zxO
wQSH+86KAmeHngexTCOU1XX4trnDKlUB8mqDoTEsqjlNrr9CWsXQAhidCnCMxcXh
nKt+w8vBRm0LACeoRKQnQw34eqW73hyNx0hw8UVVaXT6zr3MOvW+AG3Valf8EMOV
cfmX8PGy8onmF4RkYORPXwNBUAgALVA5vLBn3u3KmpFqC3IG2DeHUfi5s1pNX1L0
QPu+/tPNN9YHS3Rp+KJ7mgtTqJPnsZ1dNwRVvIgajt7ycFPE7CB6qT9KBOzq5/Ic
w71AfXVa1WQegJKqByldMa8hHkxwkDw9E5XeeED7n5hHXOMAX3l0n9nkfiM8UAzd
g+xuCoCoZZJYbgzq1KRIURslxRtGYiTvOKKNg4VEN+M4BHYobXHQeKMfG/it1MoX
cbhAP37HxmHE0GxsdcrUpUR9ExAHfC6bOi6beDGJNxLTay2jKOzKluf9OPI/Es+A
sLQQ49NO+U0tIuTpZn0dWjfkGxKYoBFmIvDJC4MdUrUMfi1UCPVCheRjpAN1Su2o
5wVnVcw8UuaIbKJKMuVC+tbTbRIU2U79SclrXRRtCyeIY/lPMlcWbB0Ql1h+ZYgD
ZqIa8KXeP/UdGz7H58ou+5tQN7LRCLoW8bhhw5YCfJFtUkvShO4TcNNF8Ose+P7O
jT7JmwM+Kf9JaoHxMvpBWOwLg/+LbDdaqR74FP+etcA9jqkop5rj+hgS3NsqvshF
q7whNRDLj+S0g5wRua1PmQK8MVwMnQLkPPLMMSuyJww7EMPTpEc2vdKzDuwiNmkZ
VKRVMG0zbiYwyAPhLX34GD8q13JM9lFJDkmM5XPxbwzTQbdmQO2Z2Mf4Zj3ZzVYe
AY00sDR3SDUd2KTRy4eYUi1fjBza8sWmT3+WLVq+IDzsp5OjYZ8ixs+VH24k8FdK
VWxPLnTyOEPFSXi526gJr/Cg8UK+4Io0gms/BCOHvNdSnsPAqh4vUvnyuHBmPrYh
ZLlUdKPiaxVsrreRYo+FbFLndwCRu9Gs9tzYS9dkgxz0f57YbbfXrt6WPUdOKQAh
Pkej5UZyhf4uxxqSi0U7KWIqx6OnupI/AcNt6otjtJjlzVsQGEXaT4LFcQe/QARF
o4Ziclgs1h9acr4oUuDPPEuEUGVrntSZlFENdZYSBXcDuSPQCdO/lHVKFX/hzOXh
LTwLhVIO3SFn3LbKparHOQODLuxKhwXPxOG9W/F2Vv7m5hBEeqFNGRwRSi116k0I
oenI/Nm793SiT6bGFeIPjY0D+z9vPETfl84bE3ARdABq8snI+/lRjBQBeYBWZrAm
sw8B9x2MfBmjoJEhQAnBP305dvHNwAtkG9iQIO+NxEoNQcqYOPw5YHl5hLQ+g50C
okHSVkYLkEwbAezi36c7jSzoWmo1yNfZUoOf8DzzGyY8IUnLVZXTlHKQG0XiADkS
pNd8lbRQSBLEj8mJuyPflFelBH0LDRwy/aeGkD+26GQEXN1PcxaBK3z9atv6u4pv
+eufMkPwzsUqRXXhOdsGTtp47MN5hMOHWFnCkXDWzIvZ2w1y3t1PNnSe0jHIHeIJ
pB05CeZalrGIaYNJVMtcdjAlQhu8cYCMJqAZ2MUDwz8sGqyp0TvCyI+X/m8OleGd
U1m5mzmgJ9q5tkx+7EQOfrTp4Tzuj+SxMRo/7Rf2IQOYBs4vIXOZzdBW5E9dJa8e
cIOq1bf9KkT2Nq0eUiEXlngh0FrAGiaK54m4TFTp1Tl1+npZPswo1lbnwiyG90ta
mIUNJO8HWI5KuqkUDc2LrBIbreMKM+/jOS5iX8L201VxJsQutJ9lX89REKfLgR+Y
nMNn1fGnMLCApNS6k3hi3dh13BvtHqNIFVgAMw3HH1H6cgB/Z3ZPgcrpCQynEqNh
n1GGtVUW3+iRMyxs/KTyHEvBCAg9aummrhICaIG/zHEjjPYc2Ujdn+pjTFypQCrH
KzBHHMBuXQgXTUVVNvTuO12gNS0/+8lR+k/t01JKIY18lGTSmF449gMqkUyy4qfI
BMq032w/nMAITX2q0Bd3KoGqRDbxRaKa2WtgimJ72iP+G5+/s82bMJ1qxZ0rwYaU
ikSRzDfUcXvgFZ0udZoOtIhnj2tFh1q0diP/gSXohu7QYkzW0l6laNaN+KjyG0Br
gybnyuNpijfyzgQowVNRE71tGATSF6RG6MKz6GE6VyTpU2atpqukNGMpqezgWsoN
3URIkBC3jSDwmLzPo83fMLYV+K9hd/CGDDBNJZmkNUUpA/p9xhYnqHHZqDw4mI7d
EppyRb09/dkC9GO8FPcSI7mFLD1ow2oodIaI9SEUxPhnrYh+Dh+NFGZ7IMUDPQWr
MnAZZTHiqJmxb9bj+1a+PiwGhjUhgDHp/u4ftFcy6R3dMKsKrkEal4SkfUqxWKxH
Si7lvb9+MUMLJMd4C0MuMM4HhJ+QoopFxWk+JeEbcLFYxpjnDfIRMRSrrZUd2/J4
VZyoj2ut30TIk8sX18NCbs8fAmhw0V5Jhv6VSWH6VivIRYVDZhLFxOoDVyA7XtTo
HGRdZ6+VYwDWH/6qBiYbSG9EOrHStwEWibIfIkkXUKNSyfJv4X/rsTkRmoJFktjc
7RV+i1Sjo9s6YZYXzA3JsVHA3KY947kjiFwmdoCgJUgCMKEGoCy4C3G4Q+4/NQ/Z
JbHiLbVEBeJ2ESrYKMnPHsvwxhcPDU88yq1ZSZnm0pr1k+if5WPwZleQ3yqxsxoO
82QVsBR6TgrRls8YDO2z3FKEoMzXdYm81TulNDGdw4GOW/GN4Olp5io4/oKkRVxZ
wHzK+M+KC2Z9f3hAlGuBp1gBti0ml2PHNhzhJPJ9YZaZU9CO2wKF5h43mlNzAsdY
AcW00yaOSizkHL1H7XRqdtacZ9nE5SWGsPYdxckArmLJeQbnqQSF7B3Rcs/cXIpW
hQ3/bGxTNj8/3ZG2+yzCQzk+tYQNGe0Sr+Sw+ccs90gq8hKHiNZEv0GImuTDZqmq
hlFfIkSyeWj5/Nw+gWq/X7S96h1sk17a0+h7SQ39NUkXyWKnXEj7G5bki42kM9lU
hII+Q+pyzW6gxdByFCww7eInILjoLjpi+TqlVa/44rWBIrSTLhdrIXzZjLviIsY/
wXwP5prhpFQtdZqMB7OnU6IgoQUHKfS2RoamXTYH8hTgKXYyWRJBph1LERpByj/+
koiqUfIV/7iEjfUUN08Qq0c0bSIs9zPeX6go1Z9YdPdEqrk07o6l7pp4cThHM1Ty
6XYZreehY/7rIvMSuTxb/ynPhT93ZUhtds2579bt6traaxKA+UKudYCQcWpedqQq
r4QeBDAW/1DYrLkEepSrwPFlITPu71XqARassRizkPEnZ6djqX9AIurpqjIfLNYF
L6igvcgwp+mglme6ecFh2f3GU+67n7KlyqwCDm1NzpUJ7jpv1g9rx6oTYLGVvC/S
piy2rsjwU4aVLGZzrOpEizLYLlP+VA4Zawn2WsDZsHc49RZBnI63Hv04rUQQl2NS
H+2nAzhIEuHa5i9B8TWcy9MHQBhajjFDqmpXnmyjfLHPTFQoP37W7jOnfGo1z3W2
X73DddfaXAbbcP+7NDdPRheHEyshg6yF8CSzJ2R62iQI3C1rctottODswcgP35OV
JHOx97Eh3zipGpOSD1YzZC/LqAOcqe6N7rJsaaDKrKzMws14/kx2zdRwaXNi3ofJ
EBYHyn0rbtMeSC7cyU38CtRZr+DfHCxqYnwmy4aNlNVrrz2awRy081wADKdW/Ekj
2OB0SwGEwNPUmsazS4ljlm5DO5wEh+V3ONzRBtqbb0mTvhw61ti+ct/6Znm6GIu4
oeeECnAM9Bjcak30AiMs1Sp7wLsf8dC4oCWgy7gg+7ctB74vmvgaalV8Z18T8obV
baAQAbHqJ1WDIrtfDYBzP9liuYMQ0oAw7lAlJ/31EV4NB+kqh5qquIwFFq6mP8Q2
FlZahbCZTuNlbN8KjNAO/8GWaVd72Jv9UXc0rGnsZFpabI0sAioZA/R3YrQcEVYP
a2y0980JKEfGswt200nNvgItfpLewUYyuCvNHPAdtIf8eOKbw1raOsN3LgdZvmiX
H1leJoFHjdLOr/UA8PKscIXMOEjXihRHWBOhA7jBfPXgg2g/Dy0Oe74T+RevPEg2
TATZwK6wBD4XbADHQDH6dyuwnZAdCGCKpJwISZnpUcFBZV5bCJQj0kDj2AWzz/FM
x8gz88A5GgKqRhaTMsfktYjvVN7MmEN1zQFcjSocIaQOof/ZABlW5k1vVji0Bb+u
zfnxk1uDOVHyY2lVhiJuXn4lEQZaqI9ph5NUwE8IwqezmWinygty9tP5D+Ts6CFO
O1Aw88Xrc7n7OybsWWB8xGCSWML8FjyC1Ef/aIw55z6G6pkkn2Hg86WXn7DeuBMT
Kq9rbnkdZAaGDvLaIzylknckS7UHLhOlowT8cIQCl4L07G1umyGwsu9AeYk1H1m7
M3Zy7hOA0xipFrnfaXKblw82+vJqDzzhSXEe9W6P/18FBMfbigMcn56tc36FfN8C
K0ybC77Jme+HhNHp4bYGJVPgdyBF1lrcncKXhMGNrlhZtU9d9S8x+P/wvuJwHX5/
Vd7zadJ5QZE7JlziIU7FRbqzBL3Nw/BeygrjVbWZdf5sf3XnnAhKCj3cL/KwmL/w
aMKNhoOpbGCClCSGZoeRDz5NMLJ93lh5a8qgRDjEnDjCCr4Wdz4MgtXRiUW7p0Y5
GCHPKWAxClhmQhDS1DWWU1oqTonbWK2uffXWS20eujj1PIM0uaIGE7+fu7BCybMF
KdT8ImeSpEEvFwB28mPvZ9fyKq3B3M2mfLr7424VcV6u1IREkDE4eJSB48fgStQK
UojJDLnGOwqSTbMkPd4FwEZACV0VUxCPhXENfIjaCUKWSYuFktbsNCcBAm1ak2ig
o9ZI8Ow+jk1UmeP6p68w2GSrjR3mC5rjx5jbVzx3f4+FU7R10DbNhvvXnZISVY70
J1IooFU+sVUgqFN/Rqt6J82bLbA3g+QE4VAL16/RUx8+KPUa5Iszvj9W/E6tU4TU
l/ulkUFCuz45FFdkb17mWzK1DOoNjJiSVaXerrwRnKUfkgaHg6G8FH7S2b/9tBR+
RDB7O+UimPfMFJMtQw9v93IjrKu4P8gsKF7zrtPvkHLu1T45AAqF70sWZXD1aOlX
LagHnN9SBgoitgb8C65kgny7AmTW+GZhf5lk0xd3EhRBadsY2PA222/rNackXYp5
NsPp+FHAanAtOTc0rQBeNaFseVn/hJSBaZwzsff92ZerbUovQpr6twqof/mAP4lK
lpm/iGFexwFY9PWao+A8CNVBVNNnDJseN6HUBXURdduFyyUDrMLV1YIRx3bR3xld
drOwPldY/DCcxz9FLdXjI8M5ZFZy8QST7gcs2grQzFX4nwOmFHL5+pXsKEJm2Qq6
XEq6m0C+xJ90bPffiBstBtlxyzp79+VqKMk8fyUaGUGwD/8ZtSU+S/uk3iXM6bR9
q4VLm4uJj5VCJoJ2kna8Pek2r8tEcmQDdtkeHc0X23poPn/sCHF2W8akqWDqeUXG
RdX4ARHD2Ykk6SpxVls3YIrtPJA6xiKxmU+STMjZOvtzZT/B4luiO3GsWP41digG
ahmzVENXOuULXF1gveLC+gTr6qmieoNjRipa9YPUTtPvPCZP0nEpFnptidoazfgW
Dpsb7O2ynYVM06bvey6j1Hv0uEpaUqvOloJHXf+Kx915+C1cZUOIyrKT7zSCUaL2
dfKYtaRgp+YCDp0vozZVfbss9mS9oO2jhZ6qM2ryIZHjT9uCtrD6qrU7We6QUbQB
0LzlH82AYASCnT27QBP0k37SHpdOWUZAAjjDJuoeS0A4zAbc3y4zaAn4uHibhD0m
ZHVfs8Kq7exADjoGBhiZ8shzPhvnbg6knH4ZCxV1He2Zn32yzIVgICzogZZAJkq6
7ICglp0uBsyjGk0zWJAYlwCavMcvJ8H/qxOrohrhxgZnC4aKnYxfhGLFL5YNI+r0
b8b87imKHzjTh1HFy3Yqc0kVmHsAU5jzc8skKrBjsgDFqdsa1tkLA4tM7v01mwDq
CPM6jE4GjG4fBP7dCy/tYfHDuA3DC5oVgS4G6noY9epjY3JX6JyK03yrvuCvNBMP
uJGccP45wMBPbj04RmwwLos/s6scgE+Ez4v2wSJKgH6eJp9laLW8AiDbkMnH4cdP
MLEchRCFbDswEN5FU/OTQpby4A+0Dc5nl4UbFOFTm1E+4uy5jGOiT9Bb9RikPAzC
26Q3W6jqF7ECAQ42fcB6T6g0D6ea000iipvpCSZhqkXNLDeGDysCGCpmi1sIRNnA
MGfxG7+iUT4aTxBn3+2eZOqdNswaOVJhF256/X3eBQyORhKk6AxGtIaX8CchGagw
jLRhoKEu8TiUg/bcBNDgWpxyWSIImVIpnvBRLHgbRFqb+ksgKAOOkJuLZTBcld4g
/jSeayYiDuEC5EyUideIb884j7zpJXmQfpIU/ZvX0Y0W9JOK9lQf+rordyYRLdoO
aW7ojSANexi3R2oQASZq4R4xqxVnXAgMVAWi4OzwQPgOK0fHfuJziOTmyq4Hqi27
xcyqiJiB9dKY3R9tS23iDr3iYMR19vPwQJkBWCagTP8d+kHMnP1XzSKS9nnqbP3H
7YciWNvrBPvX8n3B3c5q6pRq7RcrlfbYVBGe6Lvv8anC+KD/oHRgfkchuRw/ja93
usmn0f3yYRL5h7XMysaB5zWVKXlCNiGs879fItW44xsYTUl4+d+WeW84y96XDEDH
YVSj1/J/oPzyjeRVqqT8YCX7l6Hz2ReVhyvIBdKY10ox/WReO8t0wzMPS8i7TE2q
qVmXyQCUq7u5wflSKfbEu1Mg53DHDx6j6sK79SfCn4aM32tfeMxPzNHyUr/TETQX
8V1XqYafEDcDvi0xgaG2nE6lIPR1hNKMb7WPlnuoMsbkxZvLgmLop/7Q0s0V5X6S
CwVju3kGw91L5Iv+piUfRXZHJmtUSHoi1Z1hE7wdt9/lPKhkdEh643ECJjxPY/e8
xnvnKPEKhz0i09iKyW64iJ5KD1E+I0Vcu36uahvuSwM4Qq5CcCv43RuyIqjj31Mm
a/oNT0Prq04w1iOUwPbKffOr0bNPvIvKLOA6R4vhLj1JvsrvmZLToYLTvd/ThF+V
s9LlQBj2tNk9AjtPgFLzibiUG6+L35JZ7JEDrJAgiExuT7+Dxulby5YcfiUF/vRY
K/QF9Eix1K4KDeXG87+OzJw513B0IN38GqMnLdLDrnfSrfQdWL9ux6yBHweUdMzF
jyV+P7KvK9S7bvrGlzDGtu6n/YdWCeEoWGEKi0acqx3eNZxl5mX/xvSzEMiodjqS
2bElAHtzyCOsHg+ntan8cH8v+BhWECw1RR84ZyJf+kvmW26ivgsSyUUC6yPaHftp
2EETWaeIuzpUCCrq54EsPdU9A/PgukfpmWFNq3QrHxtjPwL4cEc6OvlR8aW5uEt3
hhXhckc70yQbPHoIUICB+0F7sgJ6ZD8+0IbhunkBcz7p9ffXaS5CqxClPLgKs037
dvVr8zZ1IsD3TPM5KL0JHcIaQcbu/YZG2D0ltC5QSsi9yrlgLoDNzMVhMbJBSwyv
1Sv8j6XThXKXQsJKY72mmIxKyAEBhy5RFXnC5dw9I1NafKgG9KgYuHkDecDTVyUi
34bh1FN1F5AZ+c6sDbuL17n0eMjbndvF4rWubZ5rbtavZpSJ2/p3WOMNJ/yvcUda
gb0I4Jrhm6Ntgp974t2s6Ukfa7DUiJgTikObY+/XjP2YcXeTAvXy0CetQbkzyUkb
bc0i4QWTTQ09B/oaxQq8IHT77VnAyl7jiRP5z/z8b3FT5CIwoUCIc2OfiPmVwWgd
rH/mS8COFGXgS3GVoy7u6dxZb8L3aPKdJwFJCwJKavUcqsJel4qhia4KdgrJKkB4
uMjaYtJEEt+VjyVG6EvyTLFKMFPPjP0DZeOvxHNpxz24DhCYbHSm1z2+rjmj9H1/
X5CsDV0LWzizQas1rVbJ7pJgjsw8/QU+2uQzIRTqcTe/NM+tO7x+XGwDZNf05wBc
2qCCgZJtSezeTD0riTuRYzxpOp/zYw6n1QzZEAFjL+pypYtHfFNU9ilx+UkLnnR/
54hPznnkH7Aa7vrFUcsfheWUZ/qX14coJDfEb52ycaKG1F47GNv9vTX5JdfTA1EU
StLvCKt73/8t9kpdcUyHlXCRYXhM+diBnNSqyL7KydDNsHN64Kea/RjVJAcQGZ0f
28tB3ZaTvGrjysuS3mZz4gpPwDILzF3zrS88xdY17gyoK5IoSU94zGhgsVZ97qlR
ZKDmbeQVuLRQ03SHBA2LmtvZWqABr02K1n/DzqcbfMy+fWitmVU8ep75qAYApMuu
rZQTPy5oSrP0x4eR3equbE9OruSn8uyVu3/Idg4jHnIAW30ouSo0IXZ3lODvVU7W
iqpIuZ/EHugczV7x2ucFxkL6F4PFj+D42n2esFkr3n0mmnqfJRbjQXt+IggnrGAp
wEeNQ4Q7cBmqoJNH1KnXR2BazDnTqU7o/YJKZT1JumsKwD5p+Xtyen0jX8DIocZJ
22MbyB8+/WZVVU3e6KW4B7CGa2oEHyukKTP5PnVELQH1u5HR1qqa5FJvvGOlGDsP
3QwYabJBqrYZ+jVd1xaJiDkZlOM9xF+kqg/5DB6nfrMIoZo6RljQf1BLw48nv7Fm
pV+mK3GyOoqUGsZrbVC0wfJdHUlQFlOHE5hxXY5DZ3P2HLlUjAxcEeEWX25rbWGu
6pUOIZFG2hlI8gG8hkVd2Gf0Z+VhIB1wP2BTN4cla7yN6/XIrv6FVRjuzPtFcSFv
DSUCc0JZOuAaEzmjIOdeq2oSEfhp5g0MvaVAdhJ3LsgR62rSdJIHh9aI63IHE18q
g4mIbd7FPUVgfVBDcCYmUGqEB6Ef+Iav5Zmq+wwK3l+y2aBMlXSxVEuiyMDaEH1+
MBu9MbG4YnWGfUlAb77O2cFDBuHetGEEaPymJHLHKZwJILukkaASG5Tw9Usy+naf
3x8unoJ+3gzvXi5rexqAICvPj8trPebxI5YtFaSkU9PlNp2rbDr+CNujaK2Zeo8Q
mp0SXR+/46qbLwStgx/AbXr/1EXr+Rhb6nVIuqO+hzQpiTRQeohLdx/f6Gsj+rhx
U+xeea89c4lDgSg8+VuH9Ev/OBl8SMmgFpPKpOXRfffei7IegR8w8cDcb7x9nrzm
+CGAhJmtjTYvbenqVL81PKPKHmtmjLEvoGw48uDW2CLIaKVoLfhkPT+g78geG2Nu
eRxLNr+mDgL0BndMbd5l0g1d3SzP9qsRbzrPWV9t1Rv/l0KsDuDtwJLyWqEeDo1e
Enpv6FRFFfuB0IktZvLI7VOwHToVlyYIVJKy5EFi74gT0g4rCKm0Sk2lD2itCL0U
Oo1F2e4ZJKy8adGl+1v0RgJO90Xdtsz4fsSb2VPXwCJ9tHQbBLENizxhzOdMJWhX
9tPRaZa8HAUbIDcCQj2WUIW+MqXF8aY2rl/jWhClRu0zpk1kzSXQy8dD9olf/1jx
RDx1yp/c7UWS9/709dkfEc+snkP7aMdCaCnIYsXBR9YqWNBABHqduvyWmWcJskLo
EwaFiOY9NmTT1KEh/Nuh8iE4YglIsgvAFYCePb1fT3mrEew8BdIj8WFdqhuObmCF
3uxAQ6KYJDbKUlgYUvDNyPLd5cmBm1zbhlhdpUXTGaqHaSmM5cvbnvicTxZGrmx6
aex4AXsDnkrcC+jglxFkc6IrwsA7q5VzfcObiNSInbt7Kw3RPmt1yrpZekEMVmkS
Abd1XT0HD1A8yj/KLmWTRaH+OYYdB4KU5Q5c5Rs3l9lulPts0co2SH3+pNvyqXle
6C0EhkOMdNKry79FqHikA+2Ji0zB12yxv9ZBUZSA2HiVgVAnSId4Az24ceYZboi+
2j8VNUOFqQdw2JuF5p6O0MrRaPwmgfYPUbgneUgDpXWhZPOePmYIxb3Xh7OV9zvm
/SXqcyRqZbpZ9kge/V8iDobs3RxsTYw0BRnMkjgmpxoYCA0oP8tfBwIfK5A6UD60
2a2paimh+CA7V2AuYZuZm2A1RkGh4qMGC4zIInQNqwIXBPK0lQY6DiYBqLuIq4Qm
yb+qGOGiLlZBK5eCpS2YKYkon1XluKa6rGt7UHsMvPCV4mhqPZhDfbDDTBahwova
2auPQm04zXyIYsWPxXzO2Wj3Etq6M/30Tb90XvEi5i0U+1nTcmI1KAG+Yl1nnWVQ
fG3kiBffrpXq99ne+uSwGmWE0FqrIcRFEyM/DV8M3jAxMzJRZSHMPVYu5XZf39K9
n+bFos7Vep9mmsvPDyWH8KoaSzL3j5wQmFQ+sY4Mh/wC/6ozxcTvla/qcxWc7G1u
hGNPBuIndSuIFTrXS5ujg1I+M+mbgedooYXNX68YPkANr7tmCmTucEwrYMFvuYvM
OqnjBitCIfD+ixr/jA/gCFdYMsSSQ/VOT8JAV8u80v03YuX8v403npqKErqJjC9x
3fDhaLPQzqnYotAi/4SfGaPcgDycjkoK9T4tm95XyMWMDJiJ9AVhmu4/ucxrnJRE
ew+Y+NmNWlU57zFpuPfq296vYT6FMMYY4Gtj+N+VYm9MuqiHNv8f7gTEtj5XYd9R
oLnJGBhmKUcSnJZ4YcfriQlzTmG1DdPGssb2SS1IqOI61scP1HT/lR+KACVeHqmN
I5FRvNR1YjvTf0MNN8qA/FLRSyfdOUixjdc81F/OfklmCuOlSpeEuvNkVdVjsihP
iHksbfJPhVwN5tIsnFSOBC5C2e2pFExOhpvvARQS9N6OKPpNWKXbTBbFslShdkQl
1fEcBfFlWUEUFGrK/cDIkgIChwb0uZarU+JiwSekJcLVkP+5zCtEjpsGviNR2R3x
9y5iOMCgcntgfPtZU7hcKVRqnetVMeVKJ17XGdJYS9AjXW2YORQGwvfPytqok7tZ
xksZvYOCCAB6vx1BPhyQ9Kor73QN008ssHDzIIZqwEFDk0sKIIFYb3NoQtl9xbwQ
UvAD2aR9jw+pA+oWif1e4o5zOAm3n+/ACu2w6++Y0BZ0zyhjMJEQArT8jFpG1vt9
7JmLPz5zrbJi332lvwn+ycBa+eFBi49x2rX9TP2iDqUM4jlFaDShsV8Ma8/u16nj
bKdI0F2wUQaL4ZaFJlXWRz9RQurRU9zAo6bS6sOvWjGEg9MOhErs1n+Wu8QVLsUk
sVYNPaRN/qvvPy/lQPNmlpJEF9MlEsGNyPTdbKtB/foVIDi5dg8+GkSVdDNgrX/H
Rsh9mqx0hvXSq8royVnmZLkKOItOgU+uNO2F4tkPu1MPwLK7MW/W7FxmQsHgiDh/
fUv8MwlnYWZXbz7HmWxe9QtDAiswQjbgdJcZtRg7x8xb10/lNyJTBZcxxD+AvNCz
7LyOPlF+RTNCC8bziK+WPcer5b94CJK/uBS7ovdWZl0nmAf5Bk+TVOSM9VjXpRI5
OmS9cbPKdxD0rHU/l2eGVDkw55Cwq2NyvKQsiTUnz8kxYvGHbo42xwrF7znDJyaW
JfZPmDUoxydJe3IH/OdeQjmB+wcgaYBf+Z0czRJ3s4bUXqhumx8PaPKVYekPz1TT
Z0hzEtFcoYhZU6CT/oBU4BgRWM70xOUz3AGiMrdO5B2zWO5WOxGMd9KditQUG+UK
Ks5AIsvpYeB1Ku5Qr/4bw0wHukCg4QEs5jTqoYiPiu4npaEvCdWvJh/znCwqVk9N
83zudQnx5CtyFIH5SvqnYsXo3LGbXtbOKSN/NojRRkt9lFVxPhhjSvU83IC2SefX
73wG8cXJ0w31wd8g8UrHyCyzsFv5TUQzUP5z9+rknlRfBaMrZtjUx2U5ykLJyTAw
UDNGAu2OrH5LWF+uNWxs/GE2cmh0tM5bFpLMumGyQAs4UwAcJPCzbC86jH7y65vt
P2IrvjjVPU4qvkO+0z61bjWwn7qk21RRsD7b8axDusuAmsqZkHOxjw7TiA7nDZPQ
iThzKcKAXyadHEGrSbeX217SL4LKiCk7jSaNBUCd8RwxF5+/TwmAyXBRUha5TGED
2JH7+U6BjJw5tYn9l3AV1fFhW6rxY7JY8Fw6XtUN+M5x3vYQSnOyVUmW5zn7Vkhn
VjMNMAvUDtLQNbXkrDTCYv9pBliTak+GEmmwop9uq4DOEQbnYquhTVa1pnk2kDGO
VrM3xRs9Qg42CKUiuBsht4phso02hDxNkIxeHYbVNiaA/LG0928Jd99r4jMppUye
4c0tSkVlqi420Py+Dp0lrebMJ3h2VzxIXkG3tq3gYZIdE+pCJwjAZyiqcuRlQxnu
1+HyVORmrrYih8WZVYfjlwyM2hX6xP11tFcicabGWO1gx47HcFRGOTpBVGUvF3Dl
y6Zzs7OJIlFOB/xpGdngfu3O31j3RDR0KFwPfNiV/4AqmlKdmU8ioq5oOZWyAJZT
ehTRtYbMZRoxADak0pYTEL5aDJ2Pyh14v70tXPyVbtRbJPRC2lxm+mXQWxkOOJf+
oDjPK9/43ikcYcHX18GEkDcqXVSKCOWGGTJSgSNIJgcILIDVr/1lR2DlgDqLxamy
6bK9ahdvy0RvnSaZoBkzVaYe8tjzKP4TQjUZPieWXcoOejLLPOqyTDeWFoxvt+y0
CmpC9mgidT6dzH91SfhumtSpprUmsUUUxTzQKglpCxGCpXoPrd4+9HhBeGXiE/bJ
QyTIwXnAHaeemlC5t1nCr45MbKk09lLrorCGiJOSDlaEhXbs7n/AMB5xkQtv6B2n
Np+ngFiUBF6/8ATbZKfRYEnpIICQNg/zv2iiDywVMXAMm2wqMpJ6slXRcKnqDxUi
AGxHCW6XifmupU3h7QWPoN1cUF4gw5bZgKB+KplLlASsqHcBTWaIbWmZTw5eAE+m
xIXniXucQJfDYm7ptqaMVPDD3stbnQ1mTq9XbmCALhIcp4Hj9ZpNU6kf6/2dl2sl
MLm5RWffOSaZomm0hxYZbC7sxmngvHKkF5/dcNDxNZ4fdXmeQxXMcWELBCtq7Utl
Uzmzsv7bR3E7qMD5IRvzYxLQQ06GYB/5KGClNCQG3LmSq4xrttSHC3vgnVvacMKe
v2GtLULma4Dl7Yg0VihfW21zAnVT163twYKkdWWPaBeQUWm42ifLKJEObWHW4P8y
uGfO3ETuPOrxRFcmn/NMA/tYGkzR2YAtjKtkzuQGR+bDPGbPSjfAc9qkn/FlCOqx
uO77TgNrgyev5jIgh4SkiR/BUvviZBM3fubijxOm6vJX/Lx99fR1nr1/xYZvq68Z
9yqv5SL3J7lxuuccMSqvo05a21a+s+bCzu78r21/6b4yzrnsaXEooSbR7bZy+iMu
ZJ0/P/c6dOGRoenhiDyN5D6EzrrsWRwCDyD3NVUz4ETJ7VV17oXUJG99aiR222fI
fzFMv1V9It7JdKEbzBppPkb7R688XdFcMT3tjow6nxh4JBQ/ElVlX+mxpP5jsYm7
QZ2gd1DD23Hy4ssIjX2eeCTKxkemSnMsrDr7yrKSLQb1BsWAqXfwQZPrYQgt0sbi
ZJ4G4Z94gOE07vZ7UQ+6lNJka2N/U1xRBZh5DbcKpiU6IkS+PjyGgQIadYVicm8o
PK7c12lgpqdnkUfr7VebTyy8TB6oPGrPPdGgiFG5v17a29ZBipLNLS/hZKSqjlh3
yOcdMq8ySS05Yrx2XWpEi1wjYduVAlBbCowMPVOTgK7h3TzlttqtY61orZqGctt6
gEIRWxZGHitYCHMHi3eGjHG/I7+6tWV2JKbQUqY7UXdyNuLO93MNA5m0znFLqqa1
xlhAhrDq1XKaMztSoBt/m3xpqBnhkRkIS87IK3zYwIrqLL0WUrw0x+pi6gCltW66
P/a53TKCtrg3h2AYqnThFZYrfv9keCAkb+UU2rJ2Uh53U46wQLXCgSRDefjkXT69
PnPnp/J5K3oufb1mZiHjqn58s7sV8jwErSHmD8pMFSpP+JvTMpB+lDSIrtUTMuzK
v+2UaGWINrdSS+/7PN+G+ZWSDTb6TrooPvMXVixhcKf9zFFsqqs67fvlWxNuX5U1
mEhHbYip0nQVBT+5RHeDsTe7Nt6Zj7UJsMUwA6BrTI8net8m+5T1m9w1zr4Otgzt
kY0c9gYy9O1oEsI3eB2JlzCYrN1sdFs0b1Wb36x93kyN0u3P/ssFSv0OXaCDHJGW
UWMU501fJReejajbeWhN7O5Q20sRHtA2XJGxa/hMzVZZf76XiUFG9iNtGt3iSvEE
UgAiGH4MoMBFhFjJWgYh7clmBtTJA+Y/9olZEhvvf+Q307q+jiCc6WRXwlxa3EqI
KWaMumCNtlyjBIfc4GegUBEdflQdSQZOjgbP1O/f3RrOIWCBKbLMAelhtNgmttI/
hQxIXatn71gbYzYw6XCWgImTLJIAA2S3cF++u0/DbhcH3Ss4UWSRJLfbrFZEITUN
eAHrPi8SBOQH2reCWWsLUeCTquBG9i+S9lJjMlI7bziNVzgEfOC0ep9DH/sE0Dsd
bRnfH5w5Fh1AMFD5oOHaDcuPXdHoTGJHKWWZ36wYAJpZeCKZiRe1nsJmR6f9ZbE6
mdkZ5PYPIGltKHanVfPe8dxVXDEQ+ad25LEHOQ/yBRJKpMydhka0ujmSGwxWwuo4
EsBjvGsNcfYTsefwNbrGqrISAuRRTb4ETyQYJpaM6FC56nD7kVJSQm+IX/HmJMfx
+a+qvpajhc5wlKJJJJ/hrd2zxWEPZTtA+P+6kwEHRAw8LRL2Y+pAXfZQNNtf7Fd3
6zWtfrR1OlgEMVaMqsraKQuhgCZrMxR3GyRFqjDByjKHhV1zFrCi3k6rloxE8GfC
vNRA2cO7Fwx/ejiTe/s0wirSLmBpX1eIAQ2D4T5lBVHjc2++ENEzpE090296RtQO
mGvOt+xSzDQD6NsnBZ0LsxYaUGOFxMthFVIpbNO3RSmFE9T5POLerFMoayq5MmvT
dcFr2I6GK7b4YBYSfU2HMX2o/399T+KI3twNBIsi0XDgISQvAnYzXd9x+oIRAaVD
tDvZTs+xV/+MXk4Pmlp5vjqrg4ToGAyQw2jYdlgSJWzuOGc+IYNyTX9m4EDm5Pxz
rW94eKPlgWQy0yTgkQG2JLBgQtIoIu7RKcUP1Ngf5BiJy320v9TIwehVDR40ApwY
ZqeiKiMMCIvHGBlnPFM13sy7fT+msTcQNwqNIC4CAQLoFX6efFM3ZyVNtgCFTC66
zYFNvjNELxqgiz0LPTpiCbSEnUmkC1PqjWkg6H8DKWwyT2iVE4PHQVcE3qM/U+cc
jiUC186/9DF0cUINFqqsycvZDo0lRVfCeTM83UzdSR7yW996Y1J7HDe5KMcQEKya
/8nog+kRLOUST0lwY85Q2Gu8PCYBJPjNELa23SNPPNwZDE2+50YvFJ6nl5nsIzKG
8XYeOhRS+TICXdKRS/xdnHizV0clL+MVunqYfI4NEo5NjxB43sgvXKRJ51rfCA97
5A2jNFdu+vhSP20P1XabI/4Zd14tj6oyDIzYyMiL2li9nhqVYNtnqQ9AYoEtqEwA
Fo9KobBrbK79dx400Z8eTqMtYg5WvEHIncF91ClzdxZkkONmTg8fzu8e4UOSyZVV
L8C/dr7VOik42jiGEiQka2UUGVpzeRd5FKyoRi1xlraGDt+ml7o2lg/x2P0szYFL
cDDXi7GnAdlassM37Mn3WQ5bg/yaIWkdHszTr5kmraLC0piePl2hf9RIquvvIPs0
/icPYQsyb+Kqkd1BEqjOWX6fnuh0P+ZhdAb0lY8KrAIYovAm+zL7IDN+uSp15/fT
xlee1q4r+yVHAhQvbeWPwqkTER1z6hZJ5x9iYv6jto+SiKdpy2+xodfuAVBqkI4H
PmnArtHWP1sjnGXLQB00T6lGsZFEEq4jUZoy3y0JQ0TqYr7UsyR82UPNMf5fuDjD
nMoTTTtXMcfAIMayjioTGKBVT10KMXUxWKuT1VKaiZmZVqQRVl6Db18ayXH2kWy5
Iz9lsTUxw/DVYAtOrK1RtmofWtjQJkAOoZy8M7ukVyN0QEbgS/bA4wHiOtCmFzy2
iTE2zvunFolyBrQQcJRASSJI263iekHVrLHUtJs9bOcqpSRtiKMh+z7KypDkFwyK
TZmE8h0xsjm5mFS5d7cPrYUSKtfajkQ0jjBor3Xwto64k60mTVhiBePPi7+Wmav6
ucAxkI+0BbToFR1d3yqNdthA5LWaVEb6zrz4fueCMA0qw3onL+14vCympQdjPGfk
UhtW4Zm7USWrUi0ny2QMZZ5fy56Tiuyuiyt06xCqdIsSuLxtuYMglxdRIsw5o4wV
WPLxlUAUY0capglzKW9vDM4XoQLookSex+D1J+Lamy1MUgxiJUm9MQmOcL0nWrwp
2IAaOKg900BKkI+oaqVKeYA6o3WJwyEmppzHhLFwq4rZlPT9pPeUEP1gdUVpCzdL
Kxe5CeBl3XTxgLPbdCwmx6z4dRhy52r5YiJwe/7hIfHU57QUEix1/Hj2mO0iOMVk
nzfc4V+veFIBpaTSJGCcEd6POiXiHA9E9Kyvp59+/fjgvOzp4TXpHqSp/2K++QtK
LhQXdD2zGmDfLXIrJ6bNODP8Cn0kTIYW9W6mqUV/JXoJhNdmC7C8AIuDWK7azUYz
LlBYCo2osFbiYPtF4Z/Wnlue2ZKkRoSJFMTrDXGu0hbH3xHP/oRIcyWFhZb7GYKf
1qinzxGO3VgT0D1Lij1S+t48JEOqNX+mLuNrWGm9zFrmwOM1sLgUogQ4HaQmTthZ
pKSV0ffJhZ2mVo62EF5iEaOHEF5QfZFpoBzUXGvU8jGP78H6y4TUjIAMbmfMXaHJ
6pCtu7Xpaw7rG6dF2jmB2xFbE5i0jlt0GLmyYy8sD8Llz58lFmdOwoIS6s1UKPxT
rKLo4PZuCIleGqfyK0pPc/Pk4CaRZbfzNyTeyGr1+YhF5y/4tGAxtmvs5Xsp+rGV
5Ztfnh8Q5urNpv2u5tyJmnKGvLEF2fq5X3BsKxeJOYTO5AKkhSUMCp/ve6emo2DF
NKl+g1HCWH7g9v+DBmNiDKdy96ck6B+UGw7LYA4W8Z5aibTCgH0h0z70b6Dm/XEh
GsIEKyRw4yAKqXfU6Qjy/GVFEwyKdzEzYvznDjAFy9Bt8YEnc3g3pNO5eZeOl3i0
smRTDbO8Bw+4sxG0pJdx5RhYekdm76thHLa6KCVUwTBaaGqz7hP7bbQmwK/LBOIQ
hDa+AC5Gv3Ar5b5PE2GAdoKPCKlcphMR5ZCatUHdtpaPXq+dW/Yp3JCoRvXTodRf
QrFUb3DNXb0mIwSjF4+bfmeVogrkKlbNKSRUVzmFggRT5bx0fvOsLhxb7ocH1SHD
PvLyHnZ17sGjUp5+gBMKsPG6rou9T5wUZuez0Z2XZgIcT7NsHfKsCxnCevvLt4Ub
Q3mY7+DQ7zymlPFGI8nWuOipgFGjEHcemQjiCdAzgPGtYST6v53TgIg4VI/xZ4E2
8rUJIO6Et/A938riOff/c4hl1Gl+iqOLWXire21DjScQmx7nTBEzMeS6dvuobgUH
0hV35UMtygdohC+b+8qgmQcBl7lKip1t4iDe2LFuMw9BeHNivgCtbIA3civVNQI9
8Pn+RwowDvv8RjOxSMUl4EeRBzJPnENUHKg+sOG4nKobgiH9b2NKQGcsOSOwJf5g
OblikR3Um3iPyDGBXr6B10Qk/sOdDe1qBRIBTjQQIFaYDm7JxA3z2W5N77sq5AKv
o8KvvpJ2KFpVxz4pHVWD3L0FbdD0B2pQS/49k0+7Hff7BEsHqlx95S/+iIENO/2i
ByFSMVJebQpQt7UOEQ3MQNEQhaKMKoqKL+Gq7zktcD6nXDBpuAWCgJiFIBlVRSKH
gpsxcuG/JHie8wcqZTjS2DS5ojNfloDqy6DrRgIZepjtYi3W86qG3UiCxOS9KAre
zvazXv+G7eprCOIkJ6lsk8qkXOCrRVpXPelIe8gr2lCJW9SWAyY/yn1VK+IK78a2
6h0T5F6zq8g/lZarBDHt27lrlazL9GBQn6puP+JZCf6ZiTfaoWJ5g7BJxSg0ktLd
b2JQNo9ViADA+LG0sY2ShmtWABPt+yaRvv2qAf5swKKdgL7DVaAOJC4AnvELh/ej
GhRmlbTBNHhz41upuCGxWFx8PMAxk47Tgaopy5uu5OsHTSiKATRNM+CJBOKBLpOb
Gzg0AOUDZwOuN9WudgzyPpH4/jpqNKcsSbYXRpDDFwK8oN5Vbt7v6AzN3HTSxn+p
YCFifuGfaW6tcJCDvfy+nHzcKRXUq6J0N5d+zoHjYj7bJHe1TLHAJW8KaSF5N1+g
And+2NTR0/LQ1NaBH6F8TRn+ezmLOYQ/ZvbKywJF+Lz3DrNQF/Sno9msO966lX/W
d3fMPA3dsJNkVEUGlkcQuU29RLGjk+tTRaB9N7u71Hm79fgdWq7W1xZnjrHwgFlO
V+N0GHwPzRdoStPGehml0dOAcvEfpnsPYlrk88b0s0nH/jpxcLdABUq/lY/51+ns
9G/0GHOfkkx5l6y/Yd0SmHAqW0VRZqzBv+3SQshUa0JfDWBXH+nKqUpq40Tc0xfZ
7aewfiJDIe+eJYwmZqIxtIcSJRk7ytsPJE/MFR9GLpmumgCwA9AJ8HYdKFBJz3xy
ou+XpL/GzyIY/83eO1D/GpVDm1PJ/AZcwDBev+XsiRbuOG/J2kZ4UY0mmNJaKOdd
2ZvShEtYurpC69AnY8KcQHN0WyWGvwmrKqaNysx+0THlmqA45pKHAK68LTmbPSA+
EE/CcklIsoUDvcEgPBXfk/j00Hn/QeMW3uRaZmSilvCDBnks824t5xetpENsDpw1
RMSn6xbcsRSQXIuvpNKa201hIFtQRt53MyuXYwmUJw8GzY8cXLUky2YKoiRHXrso
CBXajOMNPQu/gd5S6h6dwM0JFHwzzP2d/vFOWUviDb4zdgAVABVXF8Xa18DSJkWf
8Dj69J9w7SV8Y9qEguBle/LmdUxh4G2AzLSQI469m1zasgaBlMahuVxcpFa4onim
eR+mOlE39Y4E35TnWIEGqpD55PTjRZOmIOZvjx4f2N4Q2iIYKte3xAZGXLdrwUWT
vWroCNsmdlVSlQTe5DoaFyjbJSwuOkj7bqzd6Ts1mllze4MPYgmsBViEMDmTKTEO
yvBRp4io2paFHKaUig8oC+JtzdyXcmtGuyhPR3vnlh9pQaa3X1jMzuxKoGBGx/HV
l6Ev/q/JxFpeXPu571TUk1VkUJPsA9rW6AXf/VWxWkvPn7N/lvZ18QTYI5ELyYT/
PQCBIfgSZv7WcGHUAWrJM1hdibJ1aqWL2pyiiqZRm4GkFqHTxJJeCLvWuP9zwMMS
bHy2ID/wFatZspFEYYHMbtGMHy9FQA/sBBGbGHsPU/JbiV5Fx9/RDtv/o2/CRejk
pWSscdEnmISBixCyEnHdQoFThkc7Xgtzunwucp38RBmlin/xQMZfo4aoXPlchG/x
VLEW82zFd5uiLEV0OTSkqMVFX7OR9lN3V++atUUf3Lit/LPh3GV+6R9MX/p8fGM0
4QXnVB87Guda/rqRoRigsDIm2MZ+ll7mUTZwSgdajC90vgGbj0UKkgvnQXqlBFgX
hhL4TT+67wzlpealrr9BwV8ujloGVlUxxSxKPYU+AiIXtymP6+UMR/YLkDMOswmt
fNGkFK0OGlridUNmddFTCUZQL9SOjji7oqe531dxXSq2y6kSmmdWQLH6RAhahPTV
kbjls47WBEUOotu+Ax/cl4a+nwIKNJnVcPoZ8VeVbhZugVt0tspP3/L1CudBTtwP
523T5Cf+rkvCFGfA/UhBHDpfAMRD70OGfF8vaZWqXua7ySvlrkuUOzPKPQPXdChk
41RS1Oelnv6H5/wXyiCKfFvAhAaDeb9yEMa2u68XXXmVLhAASDThQ8dxayUglBQy
grjRRZd7kF64JYWNrQyxIfLMtLvJkAri8c5sz7Ar+ORlfXwZk3qLyExM/Is3PB61
LJlzw0aiH85GZbfTODGs8iV9hJYD/bg4pTtJWlEziCSfRHkC90d1Afh+/bSnQBg3
vNo8oDoMwi1MZgfLxNlsRhhFx8gI4GImsU0G3BCAmhZxsOBKRol/Q0kLqPSRoC1Q
8tyPk5s3vHoBt8in9cs/EpEg5ULElRaWL4NDwKkSPxIwb4iYQyQbMClE39sFRv0f
vTYDW3N5LOdG/dy58YFZxIvg1KJW5iwK03fCYgcdMpDLMT3Gmn+/sR22CXab56fx
EA/ljxwkC+/1burDaar14sMhNMjCpHXjT5qsHaMbI2n3djxRo80335p2MTXKyffU
OgSeGW3HPgYW0qTIUGjh6aaoQWPyUf9yi0b1j8rU6NJft1upJUN+dlZURzlAt4ez
Fd3ahtNYzDd8WZTjsiyzU8rZCdSLDPXk6djP0uisxzyvao2KBjc/HUOewtUy3/iq
hl6bGtIthRS6V7UTRLH9LvPuZ9f8Kh8kf2g2wMc8ThtsHaUfieyJmGgZu13JxEJ7
A7VoD5qWrnQk/JKomcDVSNF7j6dQoqdGZtzciJqRF4h6NqIjhx8CzDdOirnWPxBs
G5ibT+MaGBK49qXaTkUuF6C+fnApZ/7NuxmWrFrDNfCAOiG4k8H3YbaBIwFK4Fmw
EoqdWAdbkdoysRJtuzDthMovfKvR/8zzeARXJKiPaLBEl3MLvkuBS5w8gEV2MuP+
X3Zsg3AqEOcN/k7Ri0mQFtwdYv1blu7HuvJPLoqACARHTrP1TK0xmtHFpBvMcbAg
BSY4Q94S9usUHGdDhyqeuAhEZK/9MvtDToem45vQat4irKEZOJRSNA9szVHZ5FBE
xdDz6NXqqw6f+mcOJT7LM+e4JVrzHbh8Bx+8cLiZyl7p4a8kDc2+iEwEuIGP0P/h
LARt2BsUlb8Mk0ACZ7JV9veGN2iohD6D3tCPsBN/IuqemlxAPObMUv3DcIizBk+s
AWEBXzHcCXC/MBUx4T96cxIRfc5t0dHnU7mtSPHR+pVNMFmX38abWlY1kff6KeFL
Ur9AMhNsMmWwosgBzNliW5V9oqodtZBhIpwJ8aSSuESiJPCCQ+/EG6uEj5svHoIR
cLShuv5tG2JPdMNI74I3Uwmn5dKYXzEe7VFry1HVERZlIcccC/7E9UH40hCMozFv
YnvJixW+PId3dzkAF6As+7HDJ11wE+2q18hvCVYC/vhDju7S3+bCZyDX8kTnIk9r
rPs1vT4Tyi3KGF+Xz3m0fuCoI/1kgxY7EaMO1iDVvEqvegZ9HjVnlp9Oa8Ox5KwJ
zQiIfNgeqHquEt5iNVSCoZPv5NFxONPaV9zP2y+gyrzuzmFjKxHQr7/FLdEItD1Z
xUluRsVGo/ZK/YwQbxIhwb2LZ2mtrsNVKFUS/vS688jLRGdkXJ+jGt0I5NN7ampS
mEubkYt3Nz/KLkPVczDvp9TZiPVQBSpllJKfHZbwLukgrlj8Qim5n4VLUf4iHvh4
Inxu5Ad+GFKSG/puHxtsXYa/uo1TOtibvxZjwwqanFXuPD74UaEA/hO1nFC3P0Wj
U7v2ErixUn+Y7nS1orZRx2R/rqBs7uC4OZa2G3XZjl1ZMLdoRBtLogrytaaYXSAP
T+wF0zUEO5I0Ctv2msQTF2jZTjQLrCdeIJJgV+6PD1yECpvnW3Hl8B0rR697OjpG
RZcceP2OgeyAXlq8dVyFZr/V4K1z2RhJEcgJ97sYvoipo46IfzlZOakQyAs4Prmb
dxQMOCtbmDjuaHiZn4XRoYXYJl3ifRb29pEMTaBzSalZCqTL/Vvdjmh/ivJwQ/TJ
9bYSTmZqhFxccqYEwBC+9kdQVZdW+GbEs9T2eVY4Cf/0mQSJrbxJoh1+WUSF/te3
ednsleOAOYS+TnCu/zArAQwDG2Ne+6R+d1UKhNGKJ+PzXgwsU4Y7epjLvCsGQ5Qy
aq/lDnhb9bx5y221S2bhB0OcmF+Q1qFB3gjhnHTsARpgJnGTgNeGSSEf+lTSA4tZ
MGr2bgFKX6vpkvP40XAn2jJbE+gVbnsNdELigehj3T4j+vFh3nt5XX9Id1okdNfL
ACL2v/CvkxrIm2vPj3mZ4sOXQcVynh9pYA0D9hYIiPpkapvfpjvXFbtPPEuvANlg
pyUMh1gkZ5GcA+hkf14mSRi6z+CUANBx3ccMRrlaJL6pqe3xcHlyIOBSkVGXYzsg
00VYAHgOs7xoLHG5ndU7FGyJ27huW3b+8yvHGCbH5HNPQOimSx9WMJ40nKljnoQb
OSknA23e4Cu12XetyibQ2pQNU7Pe1+atS5okxxqORALXadPVfNEwep/uSTXYEaNK
4jxnOoI5BC9OxBNApatXvTLQBXcfJUJ3Gh5xCqBRIEUdaWWtgJ6gWxeDmoPtjjKC
Pns2FSgjXkn05VLy1CrnXt/TXmrdSDvtNiGny6RZPuaJZtDoUhLx20h2rfPU5JtK
Szg7j7J0lDJCKdjfkh55legOc8BctTour5Nu2teSVha1oOtKRXFI/I38Xc2Nqatl
M38KlNqwvoJhMctUuYOGaaevYlMQqANh8TwJ34KbUn1MUii1HRsGKtjTcKpoV3uC
q926S8T2OA6DvFDh5T5ZGf0zB9g8OMD9kE3vbxpd17qa9zlPKAcn3qVfb1NyTFLR
wOAx/FKTFSt49i1TCTsNx1sGu04JgXR4RMzDYupTnAhczHo5blPZCsqV16/48WVC
qzI/gB9gsssKn/anAk1Ffb2P6ZCh0kVLERjk05egVdklb8hUKSOqeCtUUB8O0yOo
AM3qMXNxX6cwbqnKZlqW3P4nv8AWNHnBk0xjPR80OHIz3/yR++TRrPeEaVWFjy1I
31qcKLzK/aAJHc2bqJOIAXZGrKisPp7I89MANvO8vaoYcuoMHbwn6BIwpMjFyYlJ
/rRjzBL/5mgevgawLTjK+KVvzP+n6OX8df2DTJ0WfTwzRqBTtOCFit1Yn7nyy0x3
hMlmw9sMIqX5gqbPLYd6hM8+3Yc9M7yAwh/mIKunX1ZQdQIfoj/+h9EYlrPYMxHQ
OpiLl3A2tv2nYfnPEKBSrevOvkxRAIw7L+kaENNH1sL4TCQJkg1Wx7sQMy0Uf0hL
xXe6J62hHFOIRcARZYNmQ6uUkEFMoDVn842pT9eG+Z9P1mtLtlsep6QFpG6+0VbR
f4mz4nzde12rjWb6qrz5gJZIJfWDQZWGPZWFT9LcaiesRMu2HQ/7gGRgx9hu3OGo
/ri8hS1RhUS/4aAiOVNgZ9GY2ezcJTY+3rBaP41KAPhEmO2iycxvj14cnr9k6ARI
3Gk/g9hRPgzVLJukQXENUFf2p/xIzivyq8z2Zxs7/ekLWABrsQCbWg4kMTfwMnmH
06o894rw6JR3UVjjMbJbXjghJLxA++t0oTQjUAzwD+irPI5zvxUjxHNvfxlSB7Qz
wejCkUhiJ7PIjJD3jRgFtp7CPIDTqd1/XkbLnNwMJe5KkhMx5rd5r/5sdgsFqDY5
WI0475W6YPLzBuwgYIRTRsx4HydDMF1L/uDgMXHCVh1xs2xDBTESZdTmuIKnghpn
v6amnicX5fv4jzDcyWnjrkrLoh1N7eawmsRxlzKvGUNdI1YC+Y0aRV2HG3zYNUqO
ognJPO/Oaf8Y1fYVyxTAVOpp1x2ZMPQ1TJuI4FDi+XFQZAdCjyc38gQiNHBGKEuY
9Cd+YZpS+3SvN236qZAiI2lDN5GU4yZ6xQP9yJr7M8exSGJDrwdCEtCG39t/+t+6
Y1FdXUhFZLFoTvceHUiAS8+m2K8xHhMqvPN4q6fZadsXNgioY/LTPAtWsyTxZl+2
Lnn5t453JjLW8mK2z8q+oLMaZ5cRmQoh8YKYy+ue6mK8JPb1rEM5T+TkQNSzJ+Z7
/BzpQjgV3AbS30yy5+S8cYgU1kTE46srOhJOgYb5Oa8VKb+9obiC+dHOiH84O/wJ
nM9w1rVlqBzqwmujsNlKjSTEcrGrnH+XsQMvK2CwGND+yMBl2hAuPjTNypEFu6S8
rCX/JlgqY7PcGX/O5G9UW9Flpjd3I+mHcv7y9xucPvKgDO9CqttiwOU1nIU/hzf1
BlVhJLXYTjqxUm5JcEDIi5IBhorprQQ13k0ZTdMQS/dR2Jotemxi7+Q1+k3nw6Pv
48q2gDWXdze3+7LYHnvZrLlkSt0wBSso56IT8njCGozAp/rwggoxDT9Gahd9f2A7
aIDn7uMyw/b4TIRjgEEsBab+RJYmGdHqficbEZua22xV3u431DYU2SqA00Tf+42l
I6wQT2sYwFo9fYeElTMI6DOUZAepFoMIKdg/qZtX4M51uPrnkl2nah9mJjUQmy0L
pusXSSYckab7K3ddfDTdESEdwpRg31yJHSFmVwUdP/sG65fJOe92pUvfIdOz3oYH
BSSUgfOGQN1tcZqnylpgqbN03J+E3YUcw+4psi/+KU8wSxLmjXl/gO8IiDfyY0vY
+gmlZ2mDyQQNPpN7al29Yc8Ctj1AWMfnOi3APJNngfehEVmB6dtEVck22//IXhhb
qUkF1EnjRpRQYqQFDKWYaqhgjmxh8iFL6KpvvXMT+cqZ7GpP0IQeFzgc2X8fa3i+
VLSfvnRqPC19COuyTjqDhG6SlpVkOq1wWKVFHLQOw8Gw54WaplFdcikC2GbNnV2w
8hpmUX+RcZoo1HmIo7glLxSrdW83GslJJcfgLRZgxC+J6IdEYdv9b5mFVFzuCJPw
RD1fuadB3hzvB6R1R7ylgKf6uVmnuV1VN09pjwFHNhi60Y/S9bnPNwEMJvR7GQKT
zJMENK5QX4Ty4ALzolOPBNHORBR/aXr+hDNsfM3iSfLtI4M6YdMr41+oHakXhRjX
cjN7tjsxVbBBsMgqIv1dBQQbRVkpasHWfndf0WEKS+Tm6ggH2uDcpb7bLm0fSy+f
FahO6C7lE76bX1cKRtt8ex6dDBvD2c6zpU9bqnOI8nOrvjuMlHXtxVyPJf7aHb6p
KatfgSHHddzU8Z0yBsi6DQHOlJOqJ8otGA7tniqT8PvJoOyoeSShfnPUcvMz63r9
TXc9Xlu+i/VjHRgBoFsiSD3xlWjHfBQgT9k+8rwnVxPla9hdqtWggPgPEJbqVrdx
GVW+fl5pF1St0yX00CSBVGgHNH3Tg+Lwz+WbvF7lyQAFmPJ0XcK4Tz1Wp3Il2igE
j0x4QZaUK3tLPYDhEQhCc6GzHuNkH7osciPDLMeVsVLu9gydeNjXN32wnzuzb/de
p47Ba1OwWwy9JoezzzUXVvQ4uDmmBcYdZ75IInFUfhv+u40T1uGwMwF663zvnUVl
l1aqfYcfIQyW6c0lfHQJKSsTBi+TtQzgKBDw4fdhumREN9Al9jxihqi3AhpkwUj6
6gObaFXJyM9Jwejx088peABdaA0ysq7guUqwSsmh3c1o8kmZTIj6ymq/kWXCpPg/
RGJZfOtHJbN8HIkXJyEQph5UlFvKLNr8lCaFnIHL0mO1bKFT2C84Y6H9a0D7ebKF
uzcaL9Q+otFYjiUHXskv7LwtVBErQx+Q2Nk1c5hLDgPtukrKT2IUz9bunoR2MD5T
vA6C+wzFg23hPwnc7JJ0XP3L1aeePEoCWEosbpBAUNPfsG67yMdyIWj+NQjN2mcy
W3TyoDv+r4apKiYnlFV18J4roM7CLeTGi29U8tNmEcN3xfzJYXfEvEznsRGG5TQH
YLG+CvzBKNDtVZcxEIKddL69nGuMgLaCaglGwxd7H80aqeXgFSgbR5dQpybCdbHb
Ea12cJfb2BLs3XDhn4GGLAkpcO85EDuzp/nTSSxhEhnEyoO1lR4GitKVCeJ2yxPF
2z/igImK1+QPOBjbXH9xKDrsF36zf682e+mp2aoR5TPdJbNqoQsMweyAZLFMrFMJ
Agx8gxw6tqqmaty6/15YxuVn78r2QIihkipKDGjNYZlqJudp3MIpYYTVhA367XVN
XWj5Z3HGGvusf0Fz5U1y1jUSZAvzdXscFLBbEfg1atYGEFV8vtUdpD9YuGj7HaSp
o93/kL6+LiZewiorqjJ8OvNIBpLq0gWL0nnb/j3JrkA7NCJs98lufhvBKJVk8AI1
i0WoW3jWGTaDITNkHDKbRxqh9pfkZA7iFDX5E6VDMtESnrhT8zjDQ/njivPyIP6c
NQWrDmGWTODxdacijKoxom9zxSCPLRvhHYLBApYEo8/GequGdS5a8xVE3AF1DSqS
NidhFFO1tri+Est+T9aglEfxrIlUFnZHyPuFHGMKvuk3EaC8R6FAmUs19onQBNVH
zVrfelw09/BnrOqW9Px/hzj39mG57nGH73SG+VLN7n17Pm3P0o9WL9Fz4xa/0tM4
wnQmAUmJaLFGw2C6drWaJldre8xllALEimjC6xa2tAzndJPSSzBabgoWmHhAF+Nk
s6RtjdTJd70JWJWTfoOWWQS06/7tQNH+DIihJmBavqz+kewu5NqYCj2JlbrWJ+PW
NuEHMH2fUJTwo0w5bQFO+wYI7Ycd+eXRtdgiqbaw4kfB31F8hASDTbqFPwJyN7T0
6sAlbLrYgat4qTlnWqW4EgFfemEhmoD4JGFntYEE+w+ixuJab2cZEgTZp7CgUNop
8capgNfrC2lj9Ts5FePLfepkxI7QQjg1h5mfTl+2gDT7gIlH1V/kBWFEYnq/+Tx8
l93xe/QQ4d3AXnyPw0mTHpWdpgLpuXO2RhptYugOqDpaBF3xPytKUwqt9PXNd5T2
fG5ZXnsdWaeyr0N4H+hQUX1uRXrANT5jVqQ6z147B9hbF5M9yUHJcjJNLHKL4c27
FWdmtpVQupU9JvWKaRgKGGfcW0Rtf8FdvTa9uWA+Q3+Jro7Am0O/xPjb5lPp8QFJ
9PdWFdU+PlGjh6LpcjUmJwXZC0Psq6zUsF+KjSkRAyHp8MGqC/pUFABqux0zv+W+
Ys5l5mAvl5xwD4e14sAiipmzrshzJPnmhMfQir16jotJVqi/2PnJJlVG2o+8bk/P
ygg211ywUCafw2r8U+LGzY2dASOyVvSaRN4HM5GZYqZWjQgx36c15m7JRuZnjA2V
KFZk++coXHxlnPeV53S3o40pfSbVyX6h4yEFNBKe/vy8hgU4FULIrnFft5vdHM9i
PZNz+GqKqR8Mwm/Afkcnbya2pFxRCjhoGnX+GR05Yp6OBwSuxnVLM1kT4/gF27yW
cpBnVl+Uh6f75Zz9azer1eTOwHbA6wisHNJRstgW6zG4q6V2/k5T7AfHxLRWsQ2m
f99aQmA5CJKIMusG3+CccoivWtlfCqLUGx0hxYe4+HlqKeWpl+EdDKqgwjjprA2X
uozUHNFrbVl6k2J3Lubq8eYvoZnHOGL6JvJTa+YUnuh+1gD3SyE9+F7xnicCBL8k
LkSHO3ppXnAbypnDSWLd+nAsVkTp8cpqDw9+9zw9/2i0bAefDKK6nQDTTQbNoGsL
gWMCp/r+lYA8+jnjuLaRAzP6pF4RxyD7b1lje5xFBdd96I8wwwfeCUPmxaBZtYiO
0zMYIxS6QSg/F2TwhmmNBCvRN7LgC6oV3KK/t1YgK1EEkG2EluA8mpZ1fOksAgtl
Y4PYNOivGgbWlf415+v7hNNbmQSo6b9D3o7dstAF5b9UsBRbWv2gUK+ikrVRL1Ve
C54NOQTrmHf0uml3Bl3pS1Vj1UY8ix4Wi10DyjMEyro1qtRltZpZPvu4NrY3N1pd
z3+5VsRqdoywVrk+eFCCstSqaufJIHBBQKyfl6mSU1SKSU3PcTSPjjDZ5Pmn56HN
n4i8vmxWv9t/3O+3bHOiXVEfh1hJVYEAD6a2HRUDDEECR0x7T5VvTps53Y8Yi+XH
XxtfAjH78kEsU7HAmtxU9N6OJ8PFLT+j9D4EA9aOQSYBn+VZtz4XUtzf7dMoik0g
xLHOdB0DuJtf1M4oUH/xhd8+411ab/NbZplNuhT83b53kwrCNcKPnccZwzyYTxya
ti4P9vnFiT5H2+sm+UfSWKHZHsAhVo13wwPj90nAG/LA/+SkEYuSN6H92qZTlBru
qINeVwkVUJvSB6oEO0gudAD7H+vsXU/mo4GIjfTddl0vySrRtcDqL7RsRSl+z0Hd
NT/aIOCc0+VsBeIBAMC8RbC8w7hJ8Sw/2ZCRauBai5goNOHRm+J+bA/UClsEbVRO
XUzsInvp2idjPhPGmOfMTYBIwUHW9bvwriSa01Z9fhnMq3UODf4GkcaF8mDHK74g
/trzQhwrmKkWxTv+3uaMrhTvpalPtpgoDENibHrVGKzt0PSLY0a3uh+Ex5Q8kjM9
2Jhs2OoMeBEqDZw1PoixJSegug62gBvONabdyJzFe92reoSESC/IBGs8ijdXByLh
wjRaNipGPdvjei7i8+dDcds0Mk3s9HGy0MmqYVLYFDNPWagpypPj7gtMrghEiXba
Nw1RC2IUaWkEd4TadRj2Wfd9EaDhcF0KdbMTMNDxNUPNcwW6+i8nTGL9JVbBqQl7
KQAoPqSS+0XuEMlQE1C4bRzn31SB/tcCjjvUh7EfJHgJTv5cfzxD8VjeEFPwsHTQ
vCjjfIhBSi70/YVl7iKSsuTnI+WOWaNwrQs1VX6+LqqWu53Fw/UdpAmrPYOH9gwj
/pv0hx9pKw5+1plrDo8AkWrEvGDu+ksdL/fVi06u5EEmFn13NKZsXVpk00eUWT/q
LTzCVVnTJ0jh8CeJBFrUYyLvk3lBCc5Kn99BiLyrwnQp+eBdl1SZMB7SqpbDVHg5
o/DDMexZzBe3dUPdSGOSXmzV3S53zwckEXt5P6farOXZ2INfjSsiVUKAR8WKu0Bu
aiBRhn6MWEwHG+PmcM2DowB0P1o+uX9ToDSTIa6FTT6F8wZCwjRNjrFUefMog6SD
AmbqilGxhC6jQ0iCkfPlT1eiKtGADyMiXF+FNtF1gapKUWTp0IOORJrP7UwrCb7H
xRLB8WrHNAOa/0WJqBpD3ILlrFzwJtFHTnZzHwV99WnGsWf5tNG+Wny+B0acefx2
npYULtIs/qYyiqNU043M1MSbbZEDZokaa9Fs+zrxVtb81iE186clGIKU3CQ0vVEn
V63mVoND1dXHciBZM4oYDcjlFfq1V3BEt8tZGaG4VPVGl616M+lxlkVKLDX+ySSu
dgLOLyvI61RXrOoy311UiaiCLQRcQWppObzNKiy3CqId9p8Hkiv70WureakZwTkR
fRyYYSNEzOQwnoQbsq3KchmfMjWWZoUsSoYJvBd1ciDqLLJrvOeuV/mYLLO2wP9t
8C932FcjpQer/HkZYHwKhqiaKgKMU8s8rd68s7kdEFuII2A0aCQUQpIIbJrw6gWb
e5rmPKWs2plovOdrv4ltzLoETUcaGXuKVqzjK2SuAtMnhMk1/KCBzyeUqmDi5pN/
R7Au7Uhno2NbsiV6Q+Bll59BRD3gS8M9saxiD3Vo4eUm9fN0c5Pa5uWhd4Tj66p6
uXRzswgt3pEzx4RJpXJF77q9+R9qiZkQFz3RSEeOoGPf+kYjxJV8mvCca91C/V+I
kwjulC3IR7ERDo+nEhgeUlNUIoNn+I5XjfKSPrLR9OrJsLXMIPwiCPHz2ORtDVPR
lJouCwrU9cFwHBYBTtJWDBvYxiIw/cqXWaZJ7WWlZ2V+mWxx2dw5POWbteyNBwOg
xflQqU5iBj9/XUd0IuphCCcepLEUhoAMQc9S8djcxuCiTyGS/QuYk36DGa4JssWN
gvKHAkMPUx++vGvrCPsXaP1975VWEMzhRTmhSZOua0UIxmCgEnCY4APR0DmV+Y2k
KG6LucaAIbwZt2YP4O58f4REEVR06zQGx0RNndLD9qY4eFZk/b9V3Hx0Nd08UdMu
R9nwEA7dPuA0CA6PlSnQRwgNdmtLzF+AVOsPGBZpte30eVg2/QCrjF61fBvz/Lmr
QnqBuE+LPu2TU7m7Ka+qx+qOM5dVarDSmLnXM1GrQV3PhbH42tsE5Z0QM/FIleS2
pGIGvhu7XQt1gvFYdlAgjTjbU52MwbxM6VwueHVkjIHgMuaQ6XmXaVUkNTyfPjH0
Fk440gkO00fiYE8SX/CYD9cl22h6whWer6J7ICm3XUiskpyWyf+lgj74AFumnA8h
7oVtBF+BCjcKfN8DDjyv/8IsgGQ+oCp57Vo36+aqcey5ltX5fW8nfekW77mO+Ofy
G/gn9/aXxDkguIIYxsmTGGZe/0SHaIPNQramSe5CJQlofn26blmP8RhGYMeQvolA
7PZMzjiGhBLGLtl8klGdK2/sVJIPqR5qgQpLEC/Jb08Tcj01f0tylKuMOqncwPKg
1KNFfs+HuYUvC+ngVFIs6EvWtyqPG79vVRycTM3tkQRdIFGa2dTqCjmpfXSSIXla
HrePWwcBrvldhQlwTJKFEJH8Bq730yq6EvweoRDs3BB0oFRQv65m8sfL/QAjw3JB
LitqPEATm2tgFADMk31o0tgaGCnv+5fsURG/rop+6COVTF35pjKraNskfQ6HF1O4
CbyJy8DuzB0A+yDyInQImJdG+cal02RMlimlnRSPmqdqCc1fecHqo8b/vSwdpkhO
TSDBn1Itt1EyL152i//zUZje5k1QqGkt3IolyMROuEvfWHfcmNMN5u01TqY2ApIJ
GqouqCjX6hwNSf6jtTNaqhquR0wIPEz4TXab0+UL+nemI0blO4ipw2GkARWTsB4V
TYjHTo00DmsMAVQQurbjZwvbQgoQnkrOz5r1WEzjZsg8vVbw6ySGXHTHsmhxv3wp
RYWcJw0cSXKxVWtdtVX+pmPvIgrPMWSZwxbyY4rzZnodpLufllamkmsY+MFsPpag
5YOemJrHqjx/SP5o3+ZSSJJjiKBv+BR5rRYAKImo1THXZ6ITf8eeB75d5eqJ7+Hd
fralc6DxhkZX9LEYgx1l1k0AvWD3cH18yVITuehxPtWHb+IZvhNZpNRrBg7Xjpy+
QVfmQdl3OusvcIzoaua50iV4C0kv9QTpy9qNlqKkrg+HVEPMkmcc9GEsdRCbjR3k
EDuh+BKmrX28OE9X5pruwwu1nkRHTiGPeWFaga/FwfO6n0GYHU2rqSSuQnK+QW99
t6aBs4xDcM7npRwKrBdSlOM1Ty7oqGPDIChnWVGU7DxLvWxQCWdMrJ9nzI0RHEsf
+llCiwAbPkRzJ7dCBuSfN4mexQ1z6UyEgfjgm7v91oU/2vTRgwWMo6TGC3w/9rWA
+8x/tTvpyf0GQZ53ROsPhXj8vjRLoIZqMXW0wtuER4hRWQiDkTcq1xs+YcgY7Jiq
z/MCMtftOs+NalfRHbysMbe8KcFU5d5Z9JINcw2H7h62Ri8J28JTc+ZFIV8+UQFY
fYLU2eN4cXK5VlVrlwFMkkhlos6j+1qZBOmIJZ68yYNdDOWg4uxsiG+eDtenqEv5
1a9bomZCeEsVYATn9dh83/cHwysccfvRXuSBLIi1B2RmanNnrVAgnBEllmI8iRM1
Rgrhv1PpM7kqhh2bVaTiwcLgyQSA/8fDb+mBqMY5eu0j1s+61weVQmuYWYzs163D
K3p8AEfrhO+d8XYwoTQ0MFbZF5Rrt0A1x9wbwRjlbFXgqaN7wsS6gbmNm8wXmaFQ
D5cJKZdByhB7CzmuO5OKtksvnbU8p843rm6rLxRhdso4xB2bY5ZS1vw7nhz7GVuW
d+UPz1qvWWKzc6hwtwgj3sKb8O6WT2+1jZFeSvLMCnFmBAEbpES5igmu8rOUn4fr
No4e0IhBrbeL/GlCJqtc9zqD7HnM/szTI1XFDR4GAj2+HY8lh/Xe2k05/Bi1tUkg
4o5MwH+grGQ9aS3ahSh2C/yX5rZ3q1GRqknJGu+Ar3e5V61WN8HHiWNSPQkZ7HBI
K8EarGrktJQ7rtkvY3UWxYHS/3il7jH0oNvkxQUugBxP7eR5ZrheE5gllr8GRyt5
DO5C3/wGrcnY7V2BX/H0Q6PSskm4OKKViO2AImdPvWvs1KUCB5Zwp4CLMhMAoCAG
JJzwkZXJanZnge71o0r1ZauH4OxS9rhYkUjMZM1zAGkB2Kzyh+6kNcYpNB3gYEPb
auyx34Jk9BTWdawVIJY+n3ZjR/X8hECWBh4dqnCNNhbWnh672mGXSFi3rh+Kun/h
atTKsOa6HnW87fsaMplEuu46cB5djh3BOLhruUtwWEUrDc69gYd0w5XtZja2H3y9
Btazc4AONZczBLStLYxkTrd7NlXhGrIDmP4TWQMebFJwbZfjlDtEur3I+UohNEp8
IMNU3oeflbeQjt5MAciqi0lFIsOB9IYKChwN79MxHjQKSR3CXNO1Aix272mJY1o8
F9r7Gel52yOCTy5Z9y9v3h0x4gHab+DqwfLFul3rHdI1gEG6SPgfMEghaUa6HWR1
Q85OugNhoqLE8aGZvCe9cx0XhFLy+lm6ku2x6YiqK73Bri9bQkrey3PIUrfcdBaN
kixEOkrDQXGfRUQAf8RftKz2z3gVf0Zjo9vHxpmXFZUktci5XR9xfvzJ6l7C+6xX
WCflnJmK/P9WdtjnnrX6Ikojl4QiMI11Y+sum2JEKlGHTYRBvNGReJnpw7ks/KWX
rNVgR49Np6Gh/g/9hqGxnbYEtctMH/DunrSYxdjnaz68lO2Q4laXbN3dK5Z7TqoZ
QH85HhgqI71bmNzv1bqOsg28C6wVxvEe5XQOa6ZjYUnYEbEgAnYWU7vHmqJHAe0j
2J55MO+siltfpss84ngenh7UxTMcBEDIYwDm3h1vApFQ4W/tKP0H4EOByU7vbZ61
wmYBvy8vRvksInXgJJJQMuKLfEotcLBgBPLwh5pzjV+OYr9xYFDZxGk7dNZfKNJn
laZJRlDlp5XeKz6GY9fL8N9yqZKGQ4r3XQATBzR79zZ7agRkiPBAmS9Ho5NnRijG
UMVS8mbUkzZNDMeSe7xlhM21YQLY4OEfozaZDjZOVhdcav74eGLY86Z97DYlFOU3
2oNv298vFUG2yc89B8rAGx1qDhYqLh4gEoJWkDIyGJpv+tFH+PAfnncuc7iv9DIQ
vAP4k4C+lGAHO/0h314nMaDSCKZlY4o1VRtFf8oEycsNHTdut/UIMHrmu6lx/JcT
hP14cPzA2oCTSh38f00E9u1YZ3kT6cz3dBXUsGfByMXHF3doklwzZKVLGjiaDFoc
/qn48w01e5BNVd1BdY3XXwfOIPxji+5phU0oYYIYEXiLAsK/hBVKh/HdKgzQj1Ra
uMrZOk4SBjFWH5XUm8y2a2lO2r5UALzkNX53qqj/C2Ql9c0HgC37pljMGG+eZI/i
EqMhn8AHx62g3HZCJON2xPBkMgj9EJ3U697gABYbrabg5k3ssKIInbCYrFwja36j
TfwI4wc6xpP4JShfqPnKp7Novx/ZhXfbpQIr0sDdmsXtzCrYb7EPdBpdTcF0xnHD
rkxeRIxyGpNqbM9McvCxbi5bVBJ9yQnix9GUsb5TNmDqDUnlsqL4lDc+QfV+wfSy
AbvaM4uOqbCXtJSRtdZUZkkB+acx2Xx/w+wyjDsbfg/o1Yz7J9snD1yHIeXq8Y+d
ET++5ELnmrQYKiZgj1L8MhrMyyvO3TLItpJBhxIDSU1Hy0R8ccMIr9puHjvFSbbW
hSRBG7jnQDEg9jHRSW25sqK01hpV0k68iiCcm0d7STt91YCHW+Nd+/vMmiDFiZui
/4o24GmdSTBU5N/flYd0VkyIZg9svW30qDBB6TAjHUJwJjJqHlqllqUzM9fBKaGf
4/TZ+JXTGbyqo5XPbaaWW2WAM9kA0oIkIsEHboUFb9eYfLE9aJdMN5ZKVfL7bgMs
uOXbcuqY1t2KhihLBtSfeocJKJsr3ao15/tVFldfpJnnxO2MuXq+Gp7Vs0Kx+jAm
LVb+ALK9jZFyOWamr8Mne5HP2XspMXDGC5QHzL/NJbUwCKEnox/PA+WxWET0rMmH
v/Yp79uWr5pAVGRahMSXP7EfCbnZbbhSneXng5J+84rTMN6+KC89kIiW4NUWpLuh
DDNbKMHnuxppiFdgAau8qlsbe2H+eJILnJm33DB93ZRNVfp8pvegd+PmELKGNE1d
bkwmYCaODbgY75KVmh6QVG4EeXHJZ8Yn6+nxP6m2niIHZ8s2uCpqgfictk5eOQQ7
vhWaNCXTqYsuNl2mWRVBg/k7e4HArRpsiBMtWCOC0eh4Sd59Ytxkda2OB8TzH2Sh
Kzw/ve2qysQFuTyH4poTJoauLWW0JTKDKXVd36EWX0H/5CbeYsl+5C0JrGVrkU3K
z7f2GnLoNOyusCxeFRdkaNSKEe/bJ7idUEUzALfzCgCbxLXx5KoJWFHHGHIKuoMy
WylYU5+8LlKkVKoJ4wOK85L2KN7JsSecH3aD6xCa0lqLXHnIIt1mU2rPuKxVi/1e
cnkDKMG4I3r9b65HC/kk14KBUTMXvZc/+X/Dxyjzh0AQ7U6b/fWE4nQRDlwu+5P2
mtTDEOPyqYTJX/1bagGJTcbMfj4vuqUOf1ltNyBgjn9atcbRvs/or0vtaEnw5j03
n5Jk3JRs2OiYyr4a+3/qaWs6Dsq6nBO3mD7RT2PX+43RbfZInKHp0QnENClmiIBT
uHmd3Z/38rrcgcw8YBXnzlL+aKpGsZPDrf+Ud28bFH/PbEZfH+fRzNDzoXQLz46t
J6PQ3ObJmi1B5RzkLOid1+VyRCzzcmxenRARNILJn5hjA4xXnLwmEDiEb1r02bMj
x0cB8u6/kA+nRlCYiwGRcE8GI6GOcrAxx5aMt90ewD7niTLe0eXCJtve1G08U2pZ
lxdHRvvGN1kWG8fQhXAk9mt8CcRbf70HpU3l7RHSyJMrHr/UIzbrTLu1tTTMGCro
m72dRYwCV6gvu8hhkXp9OkY5yptcAQu4WqFGuzbB9l38YLWYD+E1K8k3FtDQl4Jr
M7hf6ctFl69uafo3AZLGP9O2L7f4guBL2voLT3bEjHVGpPYwbhVwnNFv2O0gqW6H
gosbUl33qpKETjJUKW+Fo8UfQboOrwHJp2E8Mu8bhP+kqiZBGkfAuXi8Jn+JsrAM
SYYh8l+1hTuX5l4d8iWo3xFVTZsuQ5gGj/3d1TTcpgvFWPjZqx/lSHcmStVqQ6XA
oaIsf6WYm1iGcWQW01rYK3Zqm9yXn0LDVXpq5jTJSXoa1eFwB6bmnaFj0LRop/AJ
LMVzU4Tnk1mrxY5j+HZzNovv3sgr62aHiGOMP52BQegodqLAvsHdB52pYMkkbczP
rypjlrkaA+YSvKTyc6mbI738SQFhcRu31JqvHNSCLVHmjHS+Cn7rKRayFzkWkb8X
o9AYsj3LnZIbeo1dO9SnbbFnjgNlqlruEbueoV7zQXsyr+eg6zX3WYj+zTnIL6c/
a7u/9Ph0w0gkrtPMM6YI3f0aumzEW3s29n1b+tDz0Xp3g+l6d/OJq2Gy8sZcZZP0
8BZO3h274L3TRff5XMLIfBvfxYlHCcrodTk1fjy8WgFcjYlFhCPEJoXAjhWMw9za
VTH4q7JQvx+0hx12llXHuek/e/dFskRIZESiDvmXlZ8SGciGW+YS4ZCADMkrzcqq
j1ZhPZFIeu/lKkDEWCT5P6okUmf39uRXQaKoNzx4DDzqkXI0uuMtynJQBC3ixbeu
RRZ0eEFyoVB3XvFlgx7FX9nkkBpHq77QxQET1Bwvvwj6zmXBVO0NL2rDXxgcRw9u
6r/G1x4ywTyCimtJrTB2v0UPxkSh2qQqZq5dx//IjJ8toBg5O9BISBlrU6rIC70d
Lzk1DHms5SkvDZYcnRVcC2hDXRmWGbulILQAG6l1UFXAV42GJt+sO/A13Xo26gBI
U4KfPB2YMu+N3j1die15D+scfJYG5FkY1KTE5N+1+Ds+q258f6inqm4a4q+T2mNB
8U4u6ZVQq19yOmjshSxL63mxfgbEjGKaLJt3cXNWcpDpaaoYVTmA1E6eQTKuY/gj
naSnhSiwSVlzkabQ4QmAEWK9Jhi6uboBaoggRPEgyjdnhCEmEyN/TtaFvHnGL74v
rl90ykkjGlxdeTzOgoI2PTptDAVv28jDwVJMnKqcP6ThUu9XRM9/u27/jAsEu6D0
hhvLkWUbVY1fdWvZ5+k/HrswbJX5oHv/nZV+t5D0ozfBs2Y5fcmzT6X9eaxfd+hy
NrwymLq4JfHy6TJf0ZhqpG+PVI6SzyNBcghOeCfHB3YWU8jFksnKyGZoKIB4plX+
l5DO6pHZGfujiIueVqXEvTGRrsmVNjF6puqt5fQZTlEk+haE3eKKO58OKs7/3/Kv
/wMZ1irPtmQOW9QUOvYSV81O8+VCh099BE3dsweMPHv7s39LOy1ifhqg33L6iIeJ
DC22zCsAPKo9bycKIIRmZJlSlvmB2csVDJWZNxZTOriKKvxrzToW6+N5Ll5v1ES8
pF91xgDhHTGpdo2TibW0tdXwk4bsue8vYJTZ61KPUKfHx+ClEQ92FmUl9HXhgE7d
THkjyzBIcU28egLJ6PSYiZQd78PQYizgVkCL8MlxZmYHuyhpGIUw+Pwuu1N0+vcJ
LaKwGWJoJaeqgqEN4ZD+dK6mmqKWlRlgKEiAg6QXWWFu0qOmHmBQhqsyAbLNvhHi
EJgCTTZhia6CCjGGbwW9R6AJKJ2+WTOzjR/9RIVd5bXtQAJxX3m2tA1kMB6eHpcB
lb65U/DgcGkzwh5bBPUB1iulUBJ3YaYU+SG8kuyhjk8J0p8uk/98MMFCZ1IR4q9Z
9fMd21Q4zvETo+RvP56eBv/U3JwnG9bN4rWmK1zdHS4M+Tn1JiIDeVE4YGFq736C
IQ8cVRaRk3oHY3mabKOeOgb4AResGJxpAoonSTg/FhxudXq7EGLPrVORbY/0sj3h
mDKb9wEjBSJlWjswLs6vh1q2Z8ccL7dUhNyEkcSnT3dyBxZ0P0wMK2aqLvubS+aG
kyef6925RekzyOQTTAoAPMBfj3d1YSv+GHBzz9J5pqTTmepot188jiItf0QFoCvK
1Tnn95IKvVsHoSKUFJDd3zXlJvGpT3OlWk/Pd2y9Qyj4jTHPE8hKVqzu6TDIOpiL
UF4FHWyRt4vX9N9mMmpT0mfwqq4RfnUf/RN4+WB6KyNIDU5Iws1MthTf1PGw7mUm
eqwq8fjDnviN0p975NODyTsdOvjjxPbxphkuegFKvS9i4dWrNP59l9jmYWTyAYKj
athtVWwXEdROUV9NBHZQNrPjQilzRWT6ypoxcr0Wf1LOFs4ARgAmhteGVMcU6o9c
IQgtIhgb7aQmA0maJXOt1fYaFTYKvBZ7KaSnZOT8FLqbdjBlYG/O20NJ9l/sYMWG
5sxp2oKvWaoAASG2G/FSErQ0yecVzd2Lb/7Lp890X95SsuSHcPb6tViEWivTg1mC
2OrSp2W+/0y0XXhaft7kU6Vp5M85f1SYTKH859EqFeME0OJzj6ahflAKrJ+FMSP9
U2NW5Or889v9IR192xfNH0NvV4CLRPH3HYBWt1gdv0kqhs3ZutJEThz5P/tatTEC
RlZCppHTty9XVJ2qb2LNApBLFeo5K4dKl3xAA8yzeXTujd8fO9Df689L8F9gVCkB
YXhW2Y07TPSMMpwRZP+Q1kdH747qbkc1PRgyp2HqWU3ZU6M6s4K6QfHMiolQVVjs
cJIQrySLagXUtNOBo6jye93099GaEBawDa0yNZS59BmdpzfA7m8WOOOSGr2Uidbz
c9ezJZqEbTHsIibj6jLSPMQNEjRUKUFcPAWfEaPZB8XtpAwK3RomABXdEsmclEj9
dBCbnYIllrmUIjkFhCkU3JCeybn935XrC92Vi92Y1QcU8bW3FJ/mTH3VTw9/IdO3
YvxLGxVI4BelQ2JXwqRdwrdQgp/i0G5jD0qOa8OA4XmPUGky/Lnf5LgCCmTxGt/q
8M7nu5tSQILATkvAhn3QWhrJDPbF86vIWWLSwNFCyOTX50/DOb3JtxH1+fSTI/Ck
Ahdf8Zzan8IqPBoZ7O3JgCQiLp5KXUwX4dc8A3PH9iJuwBjAI9gdK941wqQqZSTe
bfHMyr7kC2Nt9HI26nWFgaVT8ZgVaySaL6MVouC9dvYW+SE0YFSApTkdcCNd6iQe
9qU1n0vXvDs4zvgGnwWXwwQnE4YzV2KFNEBYzEMJtnTt0Sd4ZYA/aYT8ZuPVnAF/
9QAGxvyiF2ky1X+xZVK6WZAarzzx0iDM6X6DeBO0gFpc55kwe0I45Wbpj5/r3Zt/
NdViBTjzccYe2jCDirwgP/MeqUpdClfXJdBts26iRxRHGzWT/19FMSTnFHBHgoOy
puLkvwFAf62h4X7IKYnr9Vk2/f7nAIAWs3LVeS47uXqB7AoGcChqXrqJLyXaYdGS
YtQv+YORlkddtDv6LMXq6sJTBtb05GouwFl+v09fsZs6oMzslBd5D5MJFAFR3r+O
t4vW+ctRhZEa2hVMc6tqw8JbSE5y6jLa7aocGWGkkMlprErkgSJKspn6jlyHSVoi
EglsjGjd5+IfcWpWmy2zqw3o0PmTnddUtBe7nP8vaj6dnee8XldvyEE3uv4KiTqh
OcFFREuTj2ksAkjPRUMyZUkS4xRGwOI3sUHv3dvJO1mdhQL7bJn43o6PTkAVXTSR
ajeCJmonjg+dsAPQxt8o6x98PrZ5EIByT2NCm+LW/sv3nfJ8qLolqYcBCS6UVkH3
GqSz7qx96gSoWnk9riH8AQs3UZMFuqwVp+Xfob8cOEGiPoVFav21lbaec3kOQYGX
hgMyXCbIRwfTfLaeGliSrF8K2UY2udumoafCGgYZmFnwYF6/xfKI57uzJFclqFZF
E7eeynFwpsEahGUOdyTx2x56cH3DRSSI3TYptwiAIsxSnY2lQXSwpGZGQFuA0Hro
JQdpTp6L1X9iALJyTDtkVRYv//MbKnGosCn27+hryZxdfuZa8kbqKMi07tcPD3S5
mCGCPNZjtIi3+DKuroujbeYd4V7fLrnMRO8qw1qjdfDixj6z11pgfuBp7Xx6oq48
Tt+o77ylfm2loOxaVDoo893qjxVG1fg3ocM60G4AMfVOAYewauHYS21xz25Vg7Tx
OtPuhPBr5S4eKVKx6T7RWlb8AjVivoe3AdRuveSdQBZvGcJmvUbF9elcEhh5I6XP
62lTTLeOd+yNSQYOttng2oH6x8TZ1ZGQTfJrK1ZxmmTUEH7F0lX0+64BF5Xgc5A0
BPQoNKmiD8KDqk9JspVnBfhIeibCaenDEu21NUYBuIWa8DlF1sQd9VPNPXnOqze+
Jcy2wPcZovbm/yU1rvT8yb2v3zfLFIP04lq+Sv/Nuv2P5SttrxrIyoLfANK4HXsO
XsYD79RfpRUf4LzPx+CogwidZsejlMXZ37Unlr6zEBD3fPkgNnZivIa87pzDgCpR
1oCm3KzUrcdz24h2hcKAaLYby45WnTATraukortcekWg0y9bJWPgDInndFnYrIz0
D3/xKhLWSsf7Chm1dK0BIYs/1bOJ/SZOrVW2Lxki+RqLySyz9cioJ0p5cE3GBWEq
hC2KAP9mXP4hvud8NvE8/HHnM4W6srltE8uUGTp0xIPsh+5h6P9V0bM3Bjx1gsPB
4YzQayFICS7LBBk/fcOyjRJWIZpeW4TFH0Vd6P5+LwnZlc0Kt71DzTR8JO3wnL8A
oAl3hbkP7Cyke3UsQzBIcoDUuxpEDipfveDtfESE9Xt+l7NX0u4HIENQbulgn6FQ
f/HMuP4R++sLO4X1zsadvOBY+WHM94ZTLZdjl67mWX50wiKhG1yFjNmw1AJgPX7B
8Xec6qpR7UcR/Mneg71zJuCW3vnEbs7+UbCyiRIbjAc/IK0wu6L5l5jqZ9U7oQY6
Q3aHY/he/yoHoSookQ8MBNhDK0B2jEGBEuf46PFlR5AQxuRuRtipELOiBVX39oFt
8pFSC7ByvSM3uzXqbs8MprgAVp1GkZnBPOvgFQD6R1Mhi3AV4uTO5KhOs/ejJT+Q
T/wZtQ648bu4K7zIZu/XnmlIF0soJAmp4DWkNbQk5w3T9BBEwZvWYxhnFK261JH9
KTU12ZBxUbZAIfA3rzHi6QIM8WAfFEUCjZRTrLqFEViSVbGcG+WvNjXcB+3lxMeP
mLYYlSLTODsUjlJzwvqxbK8EayZdXgRRUODhsDU/wak716glO0G6ABGImCFM/IXE
cj/jHtKXtYdonJ/z/QRNzLXKKw1pysBntyjrzaCkLvpzZyX2URYaJsI5uL4ANWFJ
Dghj4l2hLF9x0iUn3/mZ/xfbqMC3xC0ORsSTjeM6sG9P4mRhLsQRnrUpiOIauB6Q
F+yFornv7yEl42RPtNOfKYoMYgd/XxDBQUtmVGUV03zjOpVaA1ZdFIUTcHReUelP
53ZR5mb0jmDcXPGPqiuekDJ6iRbGJaq6atAdFm36UtCXJjP4D/N1j7sCFrsFgT42
FSY/U58sK0UOSJHo+K4WQKQnPHkA4LXXwodNr/nQ7t4Vi4AeSM1WjmOPjLzoWe/C
5nELTHf5+NTv0vsCFrH/S5ffG/6couib8IvGsS1r7rD9mesWtJBdFcRDxWp39Fk+
jfxtXmuClGnH7Le+C0KCCYU9qnIe7qqQtp/Q/PTa3frd93CcgtRPdH/7LEIZvSXl
vZB2FDfO+zyG8WLne3Qvb9S3KdAOPTN95L24IXewYkY0M4VHGNsV8ABR06CDtvlr
H10dQ1HUEfFewnOLH56PXmrY5xyoskX73B96U4xcJzKShXIskkRfeBvtPUjxiGOx
AvSn19fFDhVPBEyoMZbTlKZlXiEMIeauoX9MBmdmehynCzyM+WClWFoBIIkvupA6
pGrpxvYrVpqJ7JpMVfGI7KvzeOqqz5HqhpuYPN/SO8BRhj8TphSsAnaXdZZbToVA
DohHMi6HAgaukJowYGGe4KNPhMhyjuE2S8fT1p2feJjaiBd7SAoGGGC1AD7CkhME
graPN8rCVJuLFSvrt7SyZSSVH7TxNLvgi/uSSElu6eqbc8UsCEL7CGeespOGLZeA
ahp8MOioHTtcLP0V+jiwyZkHRGTgVfTJdqyseRpTaNMin2ngRdU5AVZ/dQ7VwA00
BKgRwklqIfRhZ13t0vhy1YlGHvUbEi402L23Xm0mGQlCF8c5TQsL2SzLACIhEm/p
65C0GMDvrs03aaGpN+r5MBIxxQfsmo2CBqIQjfjseH0WimPyrDbX0hsFZrs/B21+
m4UV0wLbqKQID1zKoV/pCIxymxe9U0jo25S3nz6Ozdq4bo0lEr5S0Q2mo/7k3t9U
pE6XasRsZjkEeeduB7BxwbCs3MCD4/dq+uhwTIf8tVVMQa2ZI6BaE3//wslYjHng
+cWtNzcdLpnGxk0X07xTfLa+qpiIScXUVohqoa4eEnQTnHpEgnLgCYvkfjmSiPbH
aAmgQ5J7q7nzn9nq1RvEA+y7kt1G/8X8aOMxSfa8U9LuHl178S7eerqCw3/nU012
Igm32dcaqQSYQBtmgrfm0QVWyeOGb6ont9fX7LY4O06cmNRyqBepF27CFgYvtDm7
W6+Jea/8f+BAMDXvjdvECnmFp3wwpLWth84iz9nHidDb/ouonV00TQBs5PC/Zt+a
+cVuqQ7lCU3RmA/MIvPAJjkS+F2rmYHFMnKr9gVgP8sKsxPJZYWGjTsGdFlrYs3B
6liIqTPi1j2fVK1KBHrGICqq1Nw5h3JBb6uwYd+7cwQ7qP8hex57GLaypc9bPfDD
8CURlxj0bib+Y92RpIxWogOsaOLC8ATNZAI7YP/0wzNDpMk6FRbouo5jfq4+6snP
huXiO/eTF9nAp5DzV0haJCqdJIG3VOH6Rx+7KunbTv3Az1Dpa4kG9cLUUfq53p8D
aNZ8xtdgT3qKdxjh4mSS5c6nsZtsKFsVnvBtDE120mX2CAU6R8hCd6yo/bg8yDei
hWbbE3eQQlvqIIPvVgcribSb5eQnq0XFRkitfWk7LRkseHZVOcV1+ZA466DfdEx5
63uVWqwnP6JV+9Z6c/1W3TNhsCHdU5pjbhcCmbKxKMMc3aic8JbA/OSFi42LXf0U
fk5DdpHZpUBtB5RHCOo8zZskiuBdVevyoCpSjK6eY07+LzQ4aBCE0B1WNZ0olLiP
KHZNqTxDxLctEDAZC6LVXL7Vjn1VbAlNmzHMPfp9n7S7R3vvWowvutUK6bOC3UF+
3dLYofDfHm6OSi/KG8PIGqiBvGQ9fKUIcraS7ivjf39DzXxhWyYx3spOAudx82wl
BozMS1PDA0T4ErGoDXew78hYMRVDBw0trId03Hf/IyCwV7vzhEOB/yKzQY/3UCr2
csCCwqV6CgNYEVsBll8YBE92yT5JilmXoEftl2o5cOPgswtFKJJMT8ohCzqSGlDV
0wLV0tgh2iJGPu1Ijd/WhQVdFIqSZ9BXXxs4e6iPq6eD1+fJz9vXQECudXHVZZMG
En7hW4AXnVeI4a39BAep2JyDDYL/UrnbAyqpty6saxPqETpPkcuc7cfBGzu31fza
mPGhlQGUqzPgdCvQ3nR649OgRCLzJbESeblbKMjSs7AVWbU2tryNPzV/NV9SvSGs
fPkl+bkcSu5H4NW8VJuCNaFJgxgnNkuLPlukaKqNva3XKBaHR6wFPsTThjHEJfVo
FJAbifa69JFYbjU99wZn57fjBfaz8ctt4E8U03hT3nNSqAPFdVamzmMzTFUS16eL
oTMLGL9/V40dXSqLLSLxC7apUbnzOBN9rupK2pzWProTFyEu0MXL+E+CHNJ/VF7p
19hXCwvQDHQn8fQyrYjWlA7TOlEbB/xp4OaJaJhV5YnvVh1FWEo9rBhjVKZfr8pk
43B65tMlgWokgx9LYFTQonhbi/GH16bV84EbGXtj5WAw9DGfBfibJ96eJ5sWK2un
Qd6EMo+4AF8KaGMV1+6Q1D4CxF4GU5+4MwujWwHWtOrA+8HMoYspV2e8BclRR8un
x/BNJxs4cWu0vcWG0nnnioOmgJrkSFXK3bzq1oUlWs2jt1Uuu4KH2PeXzNq2kOTV
Kvh9CPyKVzUbg6rXiAhEbkHNIVplytpjoTTjjdYLg5RIG74XBxRVnAv9jHHAfFTZ
qvWVPEp36A2RiCR+xjrH7Isjm2iIYrwx2K8i/bumkMGPcEKkJ+OjkVWzHcQkS6Ij
21jXP3yiOiI+Q/atyyf4DtPkwrJy0FyF+zHj+7rQUnzhMqdpdtX9DxmXELPDBw2R
7+SJugDhjKpg5GQ61wpZogpj+uoR5PPz2mS7xf1dV7wABUnSrEID+XKFIGN1iZ2+
EtMjC7rOivGEQPH5xqwWHi2KR+/8zmwxhKSRlXHd0alL++l3uzde6oDLiaXRUJGS
JbJp5Mi20m8vFtUH3upLOnkflhzIcjnaGOK4qs7CulIrcwWLePknGDxEDQDP9aAF
C7r8FbAXmxO76Dn2omykA2rldMvA+BUozSWDT9KXV9rtxRKRAo96cZrdK14deVt2
MC5a78GfYnuSecOrjvAApbenqYb0OwvUhZ0zY4uJ/vCVnu4i4pzY1IO6uYrGd0U3
hLnsd8yBbIlVibHQzpOuefkTjFXdTsdLEZPiyLzp0KwFm+hThh0S4a6T9zrFcLE/
YAywYOWSOdYqaTfFHmPnJfEwqJnwp3WbngkDnnYMVC021nXvGrQgddDJByTkQpgg
0X6PzC5ieZCJAs5RbS++K2YtA7/3tXVj1nhUGLTzL5dWUGbOl/psutkG1LgzkinC
2RDEQeDeTyYQhH4kSgtBQxpmNC0fogUOH0QX9p81xBSLcvJU8Bp9pMYklZfNa9Yx
Dt68gEjro23fAjjHP5YBLL8l9uz6b3YFynu795+evMsO36eUteHCZdtnvcb0hPp0
rKJMb0aTbMlyvozFwieqaTa+bmI/CboY1AyzllD3XZSv5z6HiJLMHC8017190vA6
gLv4BB/GJS6+s10KhLmC//RHxblmEeKH9m7uXooU0pzQwlHta2Al7dgCPvyuKa0y
7nHp7sIqYTk4CJOj286xWSc95IhtnfL3nDpQ9ovyaWcJ6sqMYCGYhi24doQcOPLo
KVFt5UuZoD0h55jhCPqxPILxba7YBbQNxyByMcYRcGYRr7eZ12VzSStlPZLtYrbM
3ALXzfwleVtdhkK1xr8J1p238Cn5oddvWrQiSF6QwE+46scck4D9HPS2gagA8b6r
zjXeXdXzdyqI6VR0/qHNR4lvt+c8B9nlKzfRCCUv6/53Pjbzlc9G88PrhIWXcIuH
awDVfdtuZhl6P8aCwnm9nY0zp2PvrftW0AUfWUZFA3qsSxI7XtCt4o0N5h0CJHhP
t9gAE6Ci2lPJXaaEGKkXti4duMhKLk44x4BCvmfOqXQhRYPBjRrdSic/j90Ag0CT
CU0um98gapXZaPeWBtejzi1+TANiSDy/BGsznEaevaLs2Knoxdpj1dM6zSqRR7b/
ZLNwRAupuT7qGHqY9CPhTpYwYJ/J7IKxHVwjS6kZbOQZgNP+xr4Rsd7UdOub1PCF
p2rk77REFDXxHPIFoVlzJXGI9kabuhIYnhXdOba1Jr9sk/ochJf7QE7Zl6lI+8yt
lM0vJAuBwE5JvpoRDgraPlX/CsmlsSIKMMz5ULwkxQuK4tL9qxQW5EmUDA93f6dW
oAsNe06k0MFTF9qulwSDlbRyu0ARAefkNNBC1TekolXKB4Ys0y24wihxH0yD3rlc
0BfFcMHEsvOvjff5OJoZWIN+j8iw4rl+Nr06NcCu/CjMG5mQIxKsrwBKv7gkKUJR
RlBjx8YAD8lzNHooj/U/3gaqRynLg3vqBw09znDnJ16fo3WVQyDff//OcCPNXzKN
JSg9iDSslPUF5JJVPmSi/kXzpWura/qJcmwr4mslXfyPi/WtYuzrNlRRS+73sdpw
yroB638W/SA1HmyVwLlL7eO0CMHRX7FKjNiDsFg5PTSKcb2Nku/jMVpLYzZWWhMB
coPTXrGRet3hEaoNNOm4LAn9JL9CMuhQtzgw0WQLgdm9++A4h3X7HtQQU58qPF3A
OUQBCrkJjLMqqhKWfW2UdtB89U3ug4e1jTlnQVFyWtDDXW47sKjlK/dv1gXqMVbc
hhq/OcVF4EmCBYI2a7fQd0qurzWHLmIODt+geU0BFpqXYVAU/1VakGSyjUkEgioB
66EWhUN72zUkIaf7BQuvwPDfV6heL82j2x3Lxg6tG4Z5l09QzylUvVbJyOhqXL6R
WUpFGAEJcltPC7JCj5kbbiLxGj0D1PvW8GQ4uWJg2dtaSZZ4oKIE7LD0P5sIMsHi
5VdG2X0Q7ZKS8LSLhvGmMiVOewIU8Hb9kbOpg2rwCMu1rHSUndYERvIMVN/EQuFb
UIYoxmr94g/8T6qBhaGngrZgDOVkqwwOLC2TCfOS4IOAxI16+h72/Tw6X2iZ5QoD
gDpF6H6fIXalN9CL4MuuKFrGjdnF1QQp0aLdqBRd+FK7CbLTdFILpptqwwFT1Qk6
VWcSrfeZJl9h0HiotQeToPGemAl0YlMKMPCXSdcmkPKyzOtORQhZMsaiPPqAX4jc
96vYXg0RZMBd8EYK64m7jErPMA/symMvD7ySLA56HVJ8T8kdpahk1rXdQPP5V3/4
AapCO6MHRt2feG54KNJO8mqYyiUO1mHHiiLCA3RkIGFFnPUgORotjVjafwfkTv3s
m4fyeeJ69K/g/Y6GJg4bCSF0AJPsVMJhceZBN6NL8hdbcE9mLKGIZfp3zo8vPNWW
BiBDiyAU5GgdeVrPVcL/T4n8ZCaOfkBIbA1e86WN+1/yE7tg3GGJW1kQsglQ67eJ
oe+h2cglHx5eYAQHp12dON78t7sezsqHWKAj64tBfmSkktMayt/OM/IRWBTjdN1N
6Q8ufTHZbdVxoUzMikbXedcibTLwQDh4ZBdS4M8FkoWV56s36gpUKDLOM9dEDKwj
wOUWoTufvQywMEa/m4rbZHdBnxeGgI37sBCXHJfFNgMRQYPvnv3ADTXawONqp/2x
1ZfD1kCgfJ999u3DvPDp/tJjSF6Yb+u0PlLDoEX8fDvg/FwhV6PmE6XcCx02KgJ9
Y+cb4gB5VOnBJqxvWpVSfm/k9U+wowntVX4KrvScXTf/VsPTinFaytsRAeozlOok
1LGDVrwbdXqUea9sjVBMfEQvR+Q+y3TlpxDUeHZkW8ei0CI/qrs94VpCwLojrr2z
chsvMsFX0HGSDjRGKvDqIdFGgSjfnB7w1qjSfMS33l2tHRD8lubhvRNG9SB/+L2k
PD2w0llfRVC1dUUUQDNBxZXNIqwuHCyCy+WlO3ENSIUG+vdPmukXrEuZUvCPoFBu
3+3cnQJ917luYJlRoIXl/zRmLDhJj0evy5AEbbxfzGovtQYFuSO5DLlosjecCy/v
Di8sFGs+LqDOFLL/QF4RyG8JCMvMTbUWlHc7tmHA3rCY98V6EjjmO8TFRs1wvIWB
w4cFFITaJHW7Sj60CmplQtpNnxNSoPg45SJ0EFIytqJjp0216CfJPaKLsfjDBjrE
cvS0zFM9WBOrDGKJ+omRy0be6FQDuG8g7y3lazgJ9qdAMsqnQ5AzdvyFZOa67Xm2
WOVZs5ejA3drzyiGEyPAX3IOj9rPbYDnX0Vf+GiHQiG30OqCIubG+FB1aFogsFP+
y6ehFmZGj4UGDgTi9ah1i1+iv6eFhL06GAEoEMvHUir8weYxiu+OR4xSe1XTe/VT
E9vGO7qeTclhHrEtJbiYc746wixwpUSRePMTfcYY8ZzXPWC4hpf3bci1ms5DzFvv
ReHwOlrIBN9sVWy7GHsh2M5Kc5Q9QVddUGRz9sEevrU021Zob67ythhb0n+SvcjY
xAIQMunEj3eiCjHr4xD2OY3S3x5T0ol4BCaQsJhC94+xD6yLspl6bdPrAddgzdKF
Mo8O3H1nkNVt97eCVD8KYqvzQyUBAwOc+0ATJfbDltWH11+akTo5m4GNp4bgdyMM
6c5Pke+biPaNfGfwtQgS3QRQYeOodCVRuyAWabWh3wvpOhZWj9PCC1klatBapnqU
j4BIu62w9aGq4MxlPRy7o23cJ7Tmvxf2Ru6hUS+dei3xLuj7N4EZ7pOLeKbD2yET
Wz4HIgrEcKmzGDxPfUuAW1H3Z3amgaVXyWZ7YpGrsnvtnt+3RmDbMoVkdYDqPjmu
Cbl9ZBB+vyCJqx34nSyXmVht7p20EHtXip79ttd16h5IabBAVEn1lr/umWBFd4qB
Ycc9wHStRCxWGyxt9ij+Eu9vJjbRFs37x/NZ/MvHAilxv0+LjjmmT03S+5GOFOGX
HfVgqwIfPs3M1ocTurNyKqk5KdWheFhNXhFr6pQwCdX59GPXOV+Miq01+d7wAfPx
rQB3DrqhMJtvrYsDWknJXT98wly9wP8c7V+ha/KGLhP25HQIYMzgChGZDM8wplHt
tf2Pr/bEosP+eueuA32Gk2Vq/BwFlOTXZJ3eSOEw9kmtR6yHotbLvVomhF1dWf2I
6cTLr45LXxVw11nJ+5MM6IdEHJ6Z/4f3eLCuf5/RY8WG1O8OMCgEmJa5wiRIHJGC
vf1YTMk6s3YSNvLH0x/XVuCEarnwD2NsChq3BSUgvZrg6zJI9h7rXVvLf2mEESZQ
5cNVEFc5Rh0D4ysk4zbtJDpXZWKQEzozGv8Hanqi+lapC5eY4Ywy53zrxj99Xnet
mwvsmfxXQ3fqjJcFeDY1GV2Ad3Qc4v0xu3B7FYB0H65mysYeZohKiufbca0hjISn
6Wx33kuYAu0u5xNnBoUxPve1Vj9yNF7+z7tv2Kuj8zBPigs+TmaTFsrNqVG1X3tj
ppxW/N9jbYR7ySs9QHsHcJqdbc5LekEXoEPWMBDbndNZWoQqQtwIiFyem7gKpxk+
+pQSWBoUENUuX1zUJaYXxsj0fgcNhZkrpWtny7+L9B5UBlbYvD0B1/9p4rz6S6tO
sdBlr/OWxDyWyif4X1hY1ZAogocfk4Fe1Y+FD1nnHKxqEY7VSISsYAIoBoON0NVn
0IBfQQqywbqWgXCwGQyvQ3ABZvP6uEso2tDHjsFXOFdr7BZ47QLF3SYnIVpIMNoo
rBvXvW51t5wYGN4HOIojoudtlhQsxHsbHc6KiCRkMD9LIc91dP6DyZqWjbkXKI2v
8tYTrrhxK9Je13gT8deGW8Gs0tKFxx3deWexHoKHnZgRtvkVS+XMUWDL+UWzQVsH
AAnePdtdbdIaPSdnEFghvaS9xRca3IbTV9YK2HHWdiuPx928juTZfxO27AXyDbVT
Mo2+uUX9Fvpy47WHKBSuwrVzCziHR64Pv3zKJ8uufyVwdjKPXPK1kNqkrz7XDzLF
QsUK+kbp2NX1ly+sOfrK3CfjsPe1jRiLfX7Qj4MP0dwfjRRA6buX7ELwvpd9JgV9
/OtqtE1kLMfamCYq2AVpyzfUd5vkxhAkj3nitClFtLhVEebfdRy+HFxV6nK61xRg
Ajo7NaHYu9at9gAwSrJCFTyLt+xitofzZPkjesRY3LAFo7MxWDI+ARarvTAFg+Z/
SiJml98kzKDqQZ0Gs/xvMLvxE65d7EdNvdsfKGwKfP1UsZwABP7CLrqDB1SYuzhf
1f549xzu+1F7GnCmFmR4+0750ArgfEzur3iiaCSZiTQbpAv0xjJQzGIYD6wb8s/9
a4lz1na8Yv7DpGrvQKMhrnVDDVo7u7s6Pv+A7PlNA0FGMA39CpuTIJoPrMJ8WiwX
ttwJ4xzT8bCC6QOrdpzlbpivuhpJk9aSrz1HJzd57JuCNV2Kl6AaODpoPujjDXW+
Oz3Hp5kR/2vLdb9P05hutefEaeKGD+drR7ZuWvykqBwnuZRmcUVlaTVtIaR8DGFd
vKsm7q8Ax0NdG341xhW+rjZudBFPJsjOu6vKvsApVyD5EVF+4hlPZzVOl2nxhQ/r
CztJd1UlQZcUyOvCM574ilwEd2H+zG9Sj/ws0FQb4L2cWvJ0TuV3Ebrr1qKTtiXY
3Y7IlFIOEzJHNOMv5JSvM5aFiJLAkSdNmVOPP8P08hHD7twO99ce20b9fN0GgARL
JcBXkdLRdrFyyzOkkGXpThTdW09qKVxhTc7tlFlioNGTgTs9jXiGN+PuG3gKQZio
ecXKWdydnqJIPCtFn0pXDe4DvtCSyO++mHe0uispQc2fGSWGovqGheqqkWFPol3n
EQ9NyphiOaqU4RZ9omyvZ/qPKirqE3iEmD8UWzODwvkrtNceWIrvxhmdOGEq14vH
o4xnnwNTKL2uZ5b1svVUtxAmEFXQd8i+RgJcv/hcMb9H0J8Ff3EtEa/pPmjaoZAS
98BcL8wUwTQyibPQPxNcXBCeJ5Ly+b5D2jAIlKojvJKwovKRXV2+0peGEkISxm4H
NICVcpcRAosFw5rRb4oU1dxweaZdFQ8lTtAKpp70/ddaxd/02xgOtavoTixGHeeJ
lq6WKgCJdizdnZQGM8Jr1rlqZhdQoEaB6SMcMOlahp5MAV1hNA9r8Fa/72a4sU0h
S11eaOD42Ysg8sKU8LjR60h+lm6BpJWGeEnbvMDEohjmgFGo2tIdmtU7snJE3/ZI
PFG5xhXZJqbarjGtwl/NVwpnGmCb2y4TwtGDAKYQmGvvEYQSu+vVlRD/mmUgxSvB
875zSG8Q89XVckNnOOQL9exHDccpSs0QIUho7Att19PHHaagGNZy5Pf3Lnbfk5xR
xdjDg54Ml6Q4zwl1ncGtZ7tQ72+JL+B5QiRLhaqRCwCSRkRp9T9EuEgvrIQM0L/H
7kg67WUaMflnWuTQlYl5sHWH0EH8jFA0WfeoAOabTAOfHR5m7BfJYH7PBPhOwMH8
teSesKR/Kt1rMCNsUnXeC0cgzZov7oweVaD8S9F8OrxbDV5nVlaxyibkg6XQ0Qin
NYyj3dtZab25k5bVew+dDUg9vtXwCpZBE+Jl7QzhSM/iSErowLf57LKUZreg1NTQ
u8Xspsg2EWkhK+/s4xBtJuNp7XCD+mTMtRqEq1u5GUH/28KdjTsnZHEh3uWkvUg0
v3ROC2oj2J9q5I0Y4X9DQVD+qQlECFd5iYYcg02q/PiPJdG0ZrN240c+iyNW/CH+
PQhOd/KGW11rREyUDfcUKd4nKMDzELemUX3bajOnFDE4uA6SrR+CbAte0VQQUVIt
wMNI4Lhq/aPqrynrMb0e0uzaXVYhsNhxjV2mfYfT2W04r82LSsgQLIdABDIsjqtH
7Vrl1TZxfgzarhUWMzodXvkRBpmgQkuPmgzj3u5VKXqJHKc3Mzb92cGWeZy/lVgn
AnkvTgXnNwKLNlPEZNwKH1HY8UkPlGFwo9KztPzh94tlbrYpLgRYhpuUt5ptYB/t
U26D9EG4fhMbT9Bf4jkhHNTbMqy1ie/Z24pnpoyKvj/doyZAQVI/qWPPe8emqx/4
MUk8aLTszjghdm2NvsHWYOgLLcv0+jD7fUABnGvf0sDoWbsj40O1JYevYJ5TVUA9
PUKOWxREZ5Bc7/iIvb92bv9otV7mXvJMzwzLHhciYN95H+PQ/SZBiEPHdHmmZ+eB
Lm18YT71yNywyIj69qpCLf24Ylc9IT6fWdHxbsUCLEN9rVNRRiBVpnUgkzjk7h2v
J4cWkZJmcLHrohLNxLpRJiOi7D4FbtnWF110YgqnAXJ9rhn8kIu/SoDxngFf07MS
YfTdqL/NH4ta01/2XSrezUo8CTqO/91J/80uAXr0bjZuG5D88x2Sr0t7ROsCAkK2
N24X6g6KQ5d4o3iI5isrtSbY+6hMp3lZbhTxtE1pcUjfaCxokOSId32sytvPObvU
k1CIcBl1mkROygqxFBS+o7tZtLHze22mwdSYvTWfyA+cfopx2dGqj1WZjMzaIpL0
H8st2mkXOIpJlZF/W2apy1hbrH1oZ7S7E7+hEp9UhU7h9J+9Io89FJV491i3lC6f
KljctnxXc5kv07fX/5JOiynwZU2f8ypRGo1hT1A8mEjHrMS6S1DEEf4L4AUSN3Cu
0IT9b4J8029xx4SnMtYHtJM4D32b7X1f0PkuokGynbGuraF2/WwRNQbu0oZL40g7
qDUmnPjzPnNiPRy9P/Njk34RtZM6+fYSWSu0WFSGR60R8uS+fnLS7nQs7HFO7HR0
CvgtgWGcOVYCo/vBot3DhxxirkkIRLPXL8KYfih1V5kXmoSxbYIVbimrj9PoLorF
eGZepPEOrmMcZ5kZNB6I5KIK09RHV72GuXUCwQQVPw5u/dU2eI22A5UWFv+nEam4
Sq8Y474VaGCTQqNMI3zE6BmrN2fun42PZzhUAueK2Ql/Mzt+t4sL7+6KucaHaG3t
wa2sIMYQqcIlNZSMrpNdp5AmLyXSaRcAawMD/PMwbV3qrJDlZUWEraDeDkB3b/yS
bp1OVrFy8wXA0Je7LoRu5WKR5yI3Id6/Ge3WjraV+wtzYt4iBweDjo7jjvooYKoe
O6Q1D2Kio9L9XE4UmI5a1pGENNpfhN0ol/foGVTO1Q2oTGmpBpcSPhSQfQ0BbbyC
86uN5wxQcrqs48ps0ULiMDCnfssPr+lJk3wuCzWrT/iPeVKJAjAZVeS9VAyYL2Fl
hQGDUrhTuZg15aaPQgNvSxt2TdgQUJQLu9ShCtIbBa2K4wQk+zqB+kdGqChhwrM4
oblL1h0ufDdr+yQZXjky04I2Xt3jml/Uo2WI8IYq5GTXqTsDXm40x3msgtMxwOfx
K7AcSvO5vuSX0yi8NssMA1fq+nzSj8TbBfVtx9yw8Ggd6p+wkD4dIHcxHyN3TCh5
Y23osINJk1U/9zSliVcBh/gF+DHOCqz30/ZtZWAnwLItYr/U/nr4vaDqve719K+v
g1o3p6eyiW093WhmVaRGNROidNOH+yOoak8a2wzhQa8IZmaVxNtTw13VzGQy1AjO
iNcTCC35Fog1nsS/0HP6bjnyoKfLbBUQijgcK3uiezFZaBnbw1TbublDVfhJ91MN
foWddPYe6LmmjvxT1J+2cD3Co1txII2Kf+JnAMB44xROFHjOpsChVNTICm/yvQF6
cv1QRBPemayhIymgQHEBN4MKkVvuRE2uOrf01+IJg/4/cmFTFbeYsw2ZSdy0yhrq
J7fD+4875xaI5hQ+AQ9qFmFdI9C5PNleuNPCKLCj0tQ4zq5GcXzP/HNFwkr5f01q
BzMOWL5Wq8vvm6takmfjjzCLOjb+8/js/gRyuhRmXhnFo1oGxoTAAHS8Nm3Mqn4a
dXLygZ1zmMZT8IrUd/vYDxsYmHDYIwZhbBqwI70+x/q4a2Lobe7rkM7DHh5vbgVy
94Wo0WUVz3FI6/NJ+uL9gUDKP1KXBvKLn9EcApB0EQfafH2a6u/4R9DGGF5StDMy
Y4cYeRy+7zJnhTcWm3ECai7Y2eW0YQkVrgtqJskWKWsbBUYm8Syz6+PGOcJnZ+Dr
MpsioB2JBXwDIjh8C1jsufzvwFLGA8eYv+IELIFdzUTIcaNpENY1u0AT5Odbc2iz
SiUsAgXRv5nxpIv+hVe8SGcFU0lpGjHBKv1NkEFFZE5qkrQQLtrHswXGDfV5B1Hm
bj42HhuKygxNcQ8tfNq9L1Xzosh7nBnaZqnBmlayVVwb0BkB2qdT+PU1Iil3+IxW
VynUfhwpePAn6/WxrvJk5S3gy5W8M6IImGKNk0lLNmRvljXx6gRFHv1TyQJby/Er
mosNFSeI2zVlS5NMmr9Ley9xSszE3dX309bgPKZMTwpP4N0nsa+1PZ7UkZWYx6J3
xSY+R8D42tAVoor9ypaTtlMXlF469h63sMCvYA060oqK1Oz4TNCVkpVDP6Vw4sSQ
/7Ip+mrEpzDf46NVeaP3K+fe7LSXNTOtbHgD6+oJuomtHA/YdPxkT3MKNaVpGCZZ
F4SNOwjLfsd7u1U6cytRe68kPUBvg5ibB76I8Xxa2lqy6503p1m/nN2SeVqQmZ6U
UJRf4gXeG+Gx99GgVQ/AHImWimRkjj7S/0CCoIkIUgk9iJAZObiK/z6370G4+Wgt
CVv/zp/9ZTpwG7yc94jX9cnxns01RZO/+irWd6Bhx7Wg0RBJgv38YS+tjhsRpiqj
zRZAKmf/Plw7wqH16SjUwUxGx+XY5bijzaiy+Uy+NTdDOtGSIloxMY7xUct0MAJO
EIMYGfmUpj9pQD4Ix6ZUQ2FOzTGXzyjtIMazZCQzk3fNCaH1sSfRfSULQGDNhrg2
4MOs2O5MEiA0VDOQAFEdCj587ZC7FrFwOOX8kD4M2rLKm9iMmqG/TsRGL7jhsjnx
hoo7TgwuEpxF4jGU5V4BoVS74tyLFd5HrFh28DKc++LSa03DKXSXsuggD7QD+cXc
Xe5kffHfu+hNx3HavkrcnHGvHVrbEbtBSf8/gpaM2nwznuOTcYFJTJx8xFI/B3IV
AgDmzaE+cIxSBA1A2tvQyLcf/8RPN+Suc81IZA8gfQfQpJ+F0qV+jL5OVynS3TXb
LmOZIUfNcwBEpIQE/7dpET6ePPUAlyWg2LHUYSncvKamXFedRh13hFUfbjXm3ZHp
2ogn/Hjk8jqHNA1jSQKol48pG3TwXcQkAab6DFRoT8WvZK1tLe8jfqAx7IQ6yn+w
9YyJPX4UAHpvNFDECPG7XKPgDW1csLpi/iWkSh9ESTFG7p7uGeSCOWqIvMmv6oLf
bW1AxG27fpCSIc3T5SISwG2GLNNNrGAu4Lu6JIcFtqyES9dNKQLhN+PLaDzSFjBo
piV4v4ylJa7CUKO86Isxd1BMSjiweHkZo9l2KDTSd0ZRKN78SK3Wi5csfYZAMTJG
eI9zCvzQMe8E6DxUVOodGl9yQ+N9VC9fnxwUku46nYNvAhHkT/GBYTFBV90F1DSS
EARTXE3JyCPU7RZKZpfxzhoGKeuq6dgQ5dpJRRhoLnqr5NEX9jS34jdkyW6fbHVc
rwaJoikuePHFfPPkYJloVkijDG25JiIyR666Tkv5UJrbLa0Bi9rI84lQ0iqL3VZ8
QMYsM7TfJlaqBh24eAciW7SS1xxAADyGet+CMvX25+Q6+xeMyA5HhfNgVQXZslX4
ml0LzFL3HivAwutKjSW8eaQb5cQryRaVuYLpwbSuBDUEPprIkEut6Ciq2cONHp+7
AjE8X4h2ckn9HNMMJOub/aNdl4PcD6ZmA1uTX37oe2DrujCEGx1dKzz81JzdtNxv
XnbFsnfWiSrzlTq6uuC1+s8g5o0GHyjg7Q5ll+Y78inRcICKrXs3hX8QX0jddGsW
4ePV3dV0kQSz8slwnqCy7FHDkaMpDgvEa2OBiKBnu/1x5rnUKLpZYBEjUGr8C00R
Eepcz24Qf7v1hN6eOfqRc7WOxj5gIKyDbOwsJHJqPIFVSktVuNcRFmXTZCB62s6f
NJ7R4q2ISBy5Z6xzdrXIdwRAm5wo4rhVd3UNs/wX2dfQ7I8/nKhWle0sEODC/GBD
+IhyU9ib42xt4QGOWeJGtGIy+xo8hPcu2nPAtkA61Qe8OHBOW3+ISug3CQqhv/v/
7aYCopElOmHbObGIoG7WuBauzlIhomMKkYcIFE/+AXGHIaEQPtsC7Y8libPr69Ed
6Z+21HUayfj5wvRFBcqryHserLlY2kw95yFJHChHEAYFUfdfYZxRpItCyNd0y3ff
DcDtP9OehK45cduie12QHVmeUNhebTuGlX5+8NatRn2tROhPAgRT9geTRLrJibpA
9FJMIZlStW5xUUt3kxFnwkXxhhxIfeF0zzyDKvSU3N2F0yaXWIKkzDb9IhV0+L2E
lRwiXZ5sLLCOOOBDz1CC7TYeyt2qcZ3RRwOTxEZKEsZlEAqu4MYq78AFw4ocFy9c
rnLSviCuu80AHKHvMSWVg953YzbdFMmWNdEVbFsBgEOyugH9lJ/3oon6jyfImLMx
Xco2rc52OjEt+MzBnXk+Irp0yegizYs9mwlnnxyrh/O8Dnta1EvY6AX5k1sIZKAw
nFn7KdaHRvmglNtHSZJ/oPebiFaXJCJiUJcoPKdhdhv9nYC+VmreJnbZxZQsORj4
oWCc0xvDyAp4VmelfeKQbeHSaDnT2d7YNLQpUx3jQzFGxXrd9k0RRN5d1xk9DXIS
7f8LxNjowuUoto9dGjhtMWL7/L0hThFAlpSLtEHxpBLynidqWRo9KxfzJz4FWdf/
Vqd9Ot4mQy3dJVnGSGVstUm1rPUfGc4b4bXU6sLvcKbyz/HxNBsM42+hvziBbaae
ezLCgizEeO7nt+5utDwnpS4hThkzaT4RQJjFXg6vCN5cnTW37ybR4uf8OCcGi6uh
nxDCpS9lnj4qVixezBt73wERrDGMAyDafu2qLzLiKP6n5mqKgqBqvigOPvumoLQ1
3eOBKUYIYFSQvKEW1x5qIu0i/F1qHuAB+CsnuPv54Tl7fL/YAsaTJhFH4N4Pr0zm
PD249VOCZXnVcnG5WZbgkW4pITEmZ+y95lqGWMw2J7hX2scg2cTywSEUxAj5vtbN
jNjttpSRif4av8qRv6NfEjnCQ91+3hhU1DwI4W0OsY6oSdREqjsaUGiKqYkjOdRb
wF/enu/KNvwrFz3VeFcle1ZiLTLEsekMeLwc4ZPNBCEpAry8hoxS0oYyMGrldWC5
ofRjYKHnvBFFJpaSMcb/DB52GG993QcLFaOzjC1cMXjLdayszY0D94OeniaAQZhA
dhNvdYTbMU/0JsubF0UzI8GugeC0A69NsQxt9e03JC+gEms/64vKdvvoe475y5z5
0ntL+O6FTx1IZgHbftTIyG+6IEHGlSuP6eNomJnXJxSSw7X3oI4BRH3jA08jFMdc
vQpS8bMy4OxxK7qmyV9rePqe4fluFQk+xaOQXgvj0ckufhGrq2WSFm9cUWUOhYvG
CTv3GfD5p5ViUt/MT4xyxC3dBNcPlJqp4P3coqMjfk9eUiacnRa+O7yLW7wbCm2G
2CSYePuwBLvYiRIBRxO7SepnpyQKmJuRqjsfSfJIgXa2xa78pKCrYwkNoFw2UhMu
lP8BDbc3JkkWEGkVB5brLsXBWw3Q2uO9CdMOsy9LBR2QQf5R3ytMJeazuHfgWufT
wNSmQJWZA6RzdfMSZfkBPUUinl9AON+9UNND90QK8HmaC47f1Lg3V/o02MH1aCNw
8t+01lk5DIVz0yzKxHbpb6wjSDIntadLb6t/XsKeAh7nryCPsOP3TIBf10mc/P6p
/Cp+4b/B/S6HDs7bV7czYyoh7E1C3oz+pwcTrOJoRjUlcafCvMrnr0q1WzB1EoH1
ZW5WLMi0eWvWzQ34Z7SclHeJSg+l8AOk1zvzxykXluE/8hDVj1M3Q5b+L3Q6knPC
asSaPTdBdCNefMP7bEK3T3i52ovwi/4DuN66h3Yn/U/gXI7eCozjPmiJ36x+TCa6
TCbkx2NazcJNDwv1s+hGNSFmsMsSyIEx4h9ELwxqAea24tLSqE4oP3FLcchiJqmi
un0Lg3cDVfEGiEZSrFqtU3UKiUoc46XzJJnscNAh5ZYpJ/OKODVnkPFz8IoFO88o
G/fpNrGAr/M3VlYmsQqCChOms2lp2lJmOGcHZZiOx9YE5FpF5Exafc8QUpoHsQ5p
3OLB3o5jBdVqT2NHf1ozhvXmLiaUngq0hVFG9o7O885BK4+HH3dlFsm9zUQOM7ez
WhGZRhIylUnO/4Dt/LDscDEjTvCNW8UZ4HXOe7X5KJVbY+xh67NIMhi49QpfnV/N
wbhblkJ2wdxVqZagAWF0CtYWwjxXEi9GOgQpWlZ9C6daoTbjHe44z7chfNpuoJKd
7Wnh6FLyjan8JpTXLylGy0iR0cSdkw7ZKiqi69Ousiv6KlXM9KSWg6S752o8Kiwv
I3lovfpYJZl9alBnrX9+/N05acd/3BSc7PGaXsKehwmimXVoZvNJkPBpYAPrAFAm
z48SPbn84gsXbXsFp7v8KJdvp/H09J4+m7DP+F/dk/e0ZMDOarDSNCOe8pQefHJR
jY1E0UoqwUtib+1Rr7wS+x3J6zN/SEvYuWDcNCLFPQM7ecFVbL5MTRYJ72ei+vtW
sCD2CzJnGaKqHfDp3x0bC9JnEYr73j0Nnf+faq8kXJUQgD46p8UgpNcNaz1IK8xf
QAm78JTnJX0apn0J4Eto1WT6RN0dYzOxSQruAOiTQMz4/NUJjwtyMjBhywh7iy29
Nh0BFzfFuvNLMVcKWjeFsFy/Kp4Zc/LKWnUfGgZs3Ihsg5uiElg3PWg1oGadnyS2
uZ0ZZQinZTSzG4GSs3MdM52wO0iTITkA42A/HpHOjOdziVUgvE9ciU3Gld8uqSvx
woOkqWZmeqvc3nlHwE1EbMR2cRBrEOtxYTQBmsX7g1Q4zxB9M5w0X0CorcxdBBNn
7jZg9vt8SBFb74zHLs1umBi5zj2FE9xxfN+zW2OcZzrarJBlhIi6NSh53yKgigG7
uOBTinQdPj+UcLPE/Kw5Haij1EyVZqTh9fpPv7DFN5jODyd5k1VvwqqCJcPNzYVB
nSSSY2S73YI/upytes8WLM7o/pjBYIRK2G6WNYgw/JCgAJDKh/CDkFPoj7PR5pGH
NeZdZ6aU3mlvDRG3KzCKMH53OfrEl4BrQ3wKEu5lUI8x689MCJlZk6RRyc4tuBSb
AIdcZvWojuMFzKiG9stohlNbZtJku441BkJXtCKGvX255NjAg3rECwoxWfT2/RFz
ddjUTApzuzWcXBOFFOgFSbiALMQEn+Etr8NX7dIIEBuYl6Ov1lJGjs4xxRBZ4OEG
elyNBPOW0rl+nkoFl8OZh/Y+YPI3ew6/hEphLq0fJd6L79DaCsCpEsotQbFeZC/K
IHqNZ4d4ObazFUj/wrGp0Hkq9yz5T9EKjvImNAxXlRuZtZLI0oOQQjRt2U8BR0Ol
VcyyWOAYJ2RgidIAzYpdAPPRNze+OjxgYxMMvTqbPiEIhqchkb70uV+UTSMiaaFG
vYRj7SYMCtDZF+4GlE6aQtZZTexXSuPwjnWQnSCxO7etiVem7lwOWix8XV1B8Jry
P4p9CQQc4MLNaijlv2m8dPrcuu4sQ+16dfzDorZHCYD1Rc74kxiTBcbE5YgIyvxH
QV7cvnm0GxngJckMVZWdCF6bWV4/A4eNz233nx/VT5Ssvu26pXRybCy2RZGcQCRP
HjcTcjIn8NBsiGFT0Raes2M0HeUjUzgYOG0NgwDbMX118khzXuyBfOSDnLGrTFxs
82bogi152vsgpTe27GBdAoAHq+L+20vCar8xACKgeRZtj3tnA/vjsO00HTB2R2JI
u8P18QFyW88267qFowDjOKLSamDdJ4OzqPDwa5wYc3af2pwVF7re2IFCgcrPDo0S
mASiHzxcqCE9aPPsR9ghmJZycSYkM/wPce4v0dCbtcbNPeB7NJ+7xuY/NZV9kIxo
0OmV7RLWT5DxCIqP24Jz5SQXHzyb5gGUhLQ8dgkjjIkQBwbRSYwlgUdcDmyJkDBz
bJ+U17GPmwUMG3Yxz3OKXzvzZ+LQEUCDZKFfzs0oWKdHJnQHFMJX7rHdyZOiuSJa
2zqlM57s1xVGrx1Y7Rq6jYAd9ExE9F6NzFsz4GxfUaN3ZYbOezYdPT6lFTxSwi4c
1ONzToV6MrPyEZzHnaW+oDRteeUcevbwoTNUTxKcqkgZSSStjU6WQdog2Dji7uo1
QLzT2Gy8/QCNE85H5M8BPhhM8QuNLE3/IloAocO2yCg6pLGqY48Edypt4OajtDuT
X889UM7/M586g68JUQINBuUqEzeHM+jt/mP9PbMyyu95mkgTTDoXwbDswOVjH3ZL
dROR7VFsbC7hp9jsXgm59LN9UP5vKIPx6F/rCYLXzEPwetF/W3Kdh1vV3Ak/mEEb
ZCc9VhAfIVq5rJxDlYj8NLPjdKoIHfuIBvXRg9TIdVzqW0sLF8GSAOxo6ReER8TE
eJcZKPvHPs0+psw++OAaHPmxdatqIOnt0DRJxsocNeimLCkvcb28rAvZj7Yw5S9s
w1Wy41ADbOQh6zuD3IuBVRCl2d+w0gOEzuzWkkQUtiQYT0qok6/mHH6QWg0UOUD2
xHVg2bnJ+AimM5Mf+OGkh9SJSlRjz581ntrz90MMSwsbcT0EQ96iGlErE+NOoWcl
hpnL7Wg1ypEa6tmkWI89igNN2JralEceO0qlQ2F2z4bSn4DODsdELhkEQ0voHZcr
dwT010kMhF6tdLEfrgNEqq9eRsSzR19XVSOM633sjvAJd8DqGoBwHtYRxB41T8H7
d5lRQG9l2b+XQVTeWF+s+7YxWPa9YSATwBRtCrl+rpXGgR2odkzGauqXa+N0ksEx
LJ8CQlZvJa/R7HwceLrxf9RvdXKmB6MrgtyqC46OeHOJHSUobRbgWn2Id2osQ5vz
XZkarM+JR9IOsc57FduPX9g/Ps6WNpmr20oKXKUzpQvAgJvWxCn4nUFFO+j8kC55
veKuUpJx3dfkZaEf5UAUEHmI+MFrMe8n15KBxb1Yupo5ryPB9onTmZbHV3bJIC/h
yN616dsFkUuAUirMp3Czz1u1wZ0eIa1uUFzkzUKmWhCvP+SMXUHyHQMBrkNNKJg2
mPcioxamUpyTqYFR9ur5uFmdCR1jGc8aIrjVPFC2NW7SMebDCw5F0i9Y3wxg60qW
JI1Ep3Z8YEREnAXus34F9SPKb/IUoNL4o4JhL3SrC3Q7qQCdc4cTRZqLAPWQlkDU
4IKC1jkSyRx3VV9s2InhuhSpzTXnCLY42N+uqxVEe1eZZWOSMgcSE2gwoHLFv1Ys
+bca4URl2w7IijEuybBtc5b02WKOT5G8GAibW+ojh2clQJdIbEJJa9M53qsa1urJ
Loi4PTUGyozavMveAbl1zOyYGVcVLCr89GiZQOOMzCBOJqjj4vkmqaZ1XQ/D6Yiz
ZWoR0k5rPrXvZ0xB0p+ZAZy00gbgnkVo3RiLzDeZ+6azNIKGTt25r+ADmwh0y7qO
uVyvXrgrwpKa1CL9zDcd2l4P6B/coF2M9R/WTayXCo/Nl1ZBw2TXy70PIrvzkoV3
RSPtQMD/EbpEe/VTm7JIFOlVO9FkQVXXKwBo4g+vGjimvs3FDjbMhO0HQR+pMJdZ
PGgOkIhIQpOZETp64mTWikLm3Dz0FZc2e7ItUmiCEbSXLbSVi01c7TvshpEFKT/h
GCSHIz3y41O+eMQmT64XfbBjYC0LvdK6tcsOtUXhdkvFEAeCWfKhwdLZl9XQW7KZ
NGU1wYF7fqsj3ZUhi87E3btUvs2XQfpjb+DiQSfR+JfHyMwMPArFfYGB44v3odDj
Xw5agcJaZMNVX1hguaisAPI4wtAFPgsf+v23kYT9j13iD4M11Hs2CzRmb2fp84Zo
qhzY6QHHybHNUsvuAMOLpeoSo+FEiL2g51x9Lh6J8r/Ba31DfxiW+8/chKZf9Vcv
xfAkHSaWBHCOUPWLS7R7e0Fp7j2wFXxyHjjEeZTkN/yvPc2gVyLCLarJ2SyPX6+W
rupUPw9FZeulhbYfu1aQZjouiTpLkFSdVWdHW6iPQNy5+0J9LH7BiX4ehMDtAHnz
giolwCveNGruTgzQQTIrW1dpBsIYfk8UQ1YnECCMzsc8yC38ycvVvPirj6BCFB2N
JCJCiIEcE/RNsPCtK5AfaWNRgrELUq7IEb1ZLMP5qb6KU0QozkQfG/e+IQsoOPnJ
XUhl+LGOtbY0+USAreMvyhdUtHxDS7wHeyR6jTvv9O2dDxVlmNM9DZm3mcqoXYpl
P/loY7GfLxXcyGP2s8PD1G0gvA1tUPk6mYLSGVc5F4TBYJeWp5m9Tsmx95GLBT9l
h3y9xDkpq+2Q+D85YiFpW8Tnj01JHr+f+P1tF0tB5dn38yls54FMe18eTa00rGW3
OkZ6vTTI0Owsdjefv6DunLn8KcXEuIk6NRtdzy9Z+cy0Co8WaRgAO8gLx+Ie3sVI
DlFRvqW3tOylJvOoSNg6cPbiZgGvaBruRXZ8t0ppmxkfSOtpVJTW5cGMTWZx9QDb
cKOPOFjg/USYoMnfGtM8ouBsUmyZm/91Xim3PIAynp1uNRSgXaA2S8I/rpOz5n4L
TQe9qiEkmz9JXZk7eoXuME4d/+1FxcaLZGeKlK/5Z4BZ3/PWk9qj8/1BDiKGyZoj
BIpn0nLOREjAKd90be+glAGMnWoqvOHKlVeuMbD1SYjO7I32FBO9/gm3Tp0aPQZ0
hIB7TdKqsjL7weiceQRUEUuKZu809WxCOmlyJcoapqGRtEimrlPH2J0mepEuy0x8
SB/ENLFhvVkyOidlS63Wp5TZvPJrPnJN5MhxGeZ7bGZVtehDknVAhuDOmuvRY8A8
WCWP1wFmw5vXoePKDNzmEMBOv6UvxmyWTfOBE0jvnJQpS1zn7ee6xSBuSmGfkrs5
VgqpZAnAe/H9jBw5+yDAsIapXKXUQJ3nNmKKJkbxvvTTpjp9+Jm857fZHnAQYgA7
mFTGRct7jim/p7+Y+Z3XyaREhQ8iGWfXr+TNtDHHHwu77/tjTfVBM54B5DesTZYY
BCmiDhBnsPEcGV8mf/ymcPR43ZboAgNdccDrcQxUukVd+PttYBjRkUvVH3pT4KT4
FGLR2k0M7PKBfec+tznI1NPL0pshyhcPl48cevuP+RtLVSDFAM2GX56POTyx174X
kU+iRR6tDOVouIKxx5nlqqokfr66LEGvCKDPYAA537SxfDUl+e8PIuvicOq5R0nm
jzUVTNY7RmCZcIlMbuMhmnJtZvNM6tOjNQNSuEcSKMf61B4ySj1XxWcVxCSuzaaI
tRKCahN31u1iZVC8OWsLOEV9ybEhHUoAxp4c1oJpcMtRzu5mxWkxN6thHqajtOc4
fRxr5WXtMaRIvEv6LzCjEjMvHKmLEdksObIRpCvTb+xwGlNLYntJgFYueJPYAXKt
NZGlFCqeA2F1+hs6WO4aF5TI60g0JjHJAzbtWN5mTlEtxJ8dMrUbQI9MgdLHFNes
AAgZN9KB7On3znpU6GEXZj8bE3HD5OrNinpkbDcoYY3hJDs7tZQTOUw/KVAQ40Tj
tIU4dYziJO603KQyLskv6i2yo9Q6zs2DpeQwV3OYpl77xe7aDR2sDZsBCPorcb8l
KR/GDlX+/7u2+JRWXfpdlu6PFwMgxkP/GWWPoqWI9qjcvCKA83nIksmSwm4ejc6f
KZGTJVWtP85+1NrLZyt/0do9h4TeChxa1Bvepf/Cbmusolg7V1DW+W6/Rj3creZe
0990rtJHbJhT9F36uOUO0390TN2KzQgJUNEc0wXRi6imBwk1VhKlYvx3Vl+xRN+2
6boL9cVRAGbsWihybA7l0UQaFOhFT5GthqsrZtzFLMCWeAhqwLmdjXyV8teYfy31
7vtc9hqLSTMM9hnwpPGzeuNaLWRfUWmnFUKixF08xJ+Ad4skP255qM/4zGKjQkI8
C+Y7Mi+yfPu/iZjpDK9Ovh0Ng4EHHIC8XAodqdlapr5i1oLW54PbegFVwgEf8c3M
uiaaikIyHUXm1GEgWOUr2XDPhoW1de+OxR9zxhsMunYgmDnDPePIgx47FQJbXkbc
yXnCuFyrBo0fz6mlwfEdBUo8oEx+cAPfsRBQJf8+ZD/MIkfXZhd+9g0xx7Lh6T9+
qL0xuuh8pdwMKsq+Cl5Ze+f6SvmHLupzw3SeW2ALtFMlR6NS1fq/gbEzr4fHM4we
/0d5Sxbqh6tByNxFyYncCRjtKLQwSKBklVEy/RvG1lVtpZjAqGh5wp9duAeypu5I
XULJm4VrSH4rRjTz6M/xrbcl4E4I45OqmsLdm5DdKmR8KCC3lQupEOWboq92w46/
t8EDug59U7uNroL/cQL00DRXOU7JLkz8cZE4lPVQ0tVTpzhNQ2v067qvsgKYx8Bd
RiC7w91uNvhETzltJ3nWn89uaz6DdLvz+hF+r1UOS8OEt7xeAZq7Eho/WUbaidF/
XjuJBt1H58M1+Q9cd7I37/7hf2mTVtneDd/LWHz7ur0HdMBzXRNdQkQ5Ky6DFj67
4rQrWDWsSxboeHslCE1IROVJCUMKSkH1CKs9bl2VdqMMO41ogmbfw1w5zJVCg6eq
pX06CsfIWFRw5xYSRb1E+ev6YaRZprG18pYXXmvziqUvAR324KowcO894yYThRCG
bT4GcesokM8bYAG3+a5NHBr8xfwHI/Mc7jNz5KCcjgYWhy/g9/e0MXg0dp1nSnOr
pHx73ob6ZCg3fk+GAgkY//2OpC/1tzPn4idvtlKXLMVPma7dSZ2O1JlNcc77tkOt
B3m00TpUsd2AxmhaPdFGzCq1WLbShX5bO5wP0tPqpPtaeaUVtldecqlIBuSzsL3F
ByMDk533Mby71jiop/vtI4yk7x9LYXCrAtNxroYyHk3bi3oeY4kUgwZT9Zsah7wS
qn7KcezIhCL4igw8v4h8CsOTi7Sk0hmUeibWmegpr/QeK1Tf4aqsaj/TJ/s3+A7p
ZeSDTWddb1tLNF+m9viMkhBD/iiLzjby1g0TF5fylaYFQt/6HgMTTyDT0oB6q2CQ
sWcpDVkudV06FoYTSzFeGpFn4UYYgrMrdau5kp3Ln02Km4vYRcb/zEc77S5Ic8Pr
l26iHojh1jrZ22c7Fj5tUZVRGzJq8S/7SD8JL8A9IXt6/HIY00In5LTfjEDuSOBX
pznvcVHiIyFSNqDaKw2Ve5HLIg0OYjYvIeX0K6l+YE0a+SPdQ9ZTgIhy3dJ4G+Zi
9nBBGE14P0etQW8IDghVlWT5spwCmsQGyot08usYHmW0227AiQcJvA2FMKZPtRjg
cB7C61LWZiLgQ6JoWBxozvZpVHtuDGaIYDPHATHg7+eA0QneRyy/mPT0zuYmiMvn
VOZaN2RwRfpHxvrfSCbvz3F/25twwcMlDQWbJ8YJaLuYm07ymTXXshcvsZ/RzifI
iNU7URliPj4TcOW+OkvL6FbJk+5p2QzhfEyCRgN5tZ/IhDglAzF0xhrJ5+dBWhHx
Gv5HsUdlhzBLRIdoUcQoTH+x52dAiwSDjl/e3yqqHgdfyOIKTVr0V/KToWZuXQCo
mU4Onq3QZIoyAGgR8WXNKBd+gLdcNKiJha3Z4aZKn+hLRnxvbQA9yQxl8+fYhHOu
UW01YgLrvWZ8DPczYxhJpQOhmdVKEIAMVdV6LvVpkOLy57TbVBGaaoshiol/CkJg
by4YUQB21LII715JKuh/lfDIvlVQxod6sAk1Jen2pQAvneJkvy2qcR87BVwn0XPk
yDYvYGN+EbWlgvt5bktNTY0CkiO3z60Xhn0HbY3PEPJGrawKiopfeOlgwBx34uvs
qIgTVjJi0DGCeP3up3Nx1DZm61JH14/hbM3UvoDRmyblaREFVhAsrRuWrCaCAAon
BkQKjOfwC3eQ7ePzD7Sn0GQ2kkvpSiVy/iCHwC/880IzUrI54X9m2wl2FKMuKo52
8IjbCcQqw4IqKarIREBv0rHrj7KqxViTPgl6DdsG4Ds6zF2nQCtpvAKO3xb1X1N0
aM34AFi8Ss7HmX8EGgN8H7Ep92l4vmQMAknbuR3InyZ76HGQVfc8NR/7wI0/0bLh
QxLkEmR/aDh68BvkoZHKWF3YWao41+yYHHNu6kZeelooJZkmCyrekvLP4jocaX2Y
IyukDjzYBBuQ6IUUI6ANWTWR/8el7pOZhMR7NERIDpe1ixx8BWXBEctO2SbtkSug
XDzInJiuUcR8nG1Ptob4lyBpNLzQAL5XeuqdjP7mzQfktihb28jIpwoEiMqcJ8WU
X57hPtJh1Nb5WOVYPAmZKSwsGEyxI+fdYYN3u/+biiELNvXhvElAk/RIgqoH2PTn
e8LZK0OvyJIay8aA0M+FqVlEaMceBU/K5cRkT/TT6vWLbsdpvqKtstmYCGsPiqxY
QTx+rVRY8ihUHsP1uMcSir1wH7HeRD1HgMb5yCqsRdSnY5W2laQRT8o+iEj5MNGy
SJ3E6vrsfh4V/Io+uVh89usmrX/MUrbJlPgj7jpafZdKP3YPgdyJEFNkS4Vb5DXH
jewX2KvZuH53MzeqAC1uae885iVXWTmxjJVYepLc4pNprb4Ux5WM4aFFxmYfZIk7
utrvTBWUa/akeIXAiJ5Ce+HRY68aGVHUmi8pmkjD0Qs6Y6mi2uctF3fizd56OFeb
yjsqkqQ2AvJZxrmfa9qzZrXgCbFGE71+Zu7z2vAALeW0E9EFHSFDn8FcUPZPLLFK
KZHrNGAQkC7tl+t0qdwYPv7YIAj03qa4/Uzye6t6hWwsj3WBpVjeocRuq4hCnWjw
0+7mz45mvba+EkAI1OYbRH5BkJWx8eKtjahGwCk6wchtREJTCSQQbx280b2iRtMj
YBSZOd3MAkzQg2FgSRJojN3sd+Nm2QNL7BCOxJq5vaxsfkrYVWZPUkHa2RJ3gxOn
IH+MB61lAm/CvG54rL4+h7mDWuTs2ktIiiZgZzGfUMpc0xkKvzBiiEnbEAlGILRa
EFvouANrqHBqxmGRqYKEvk+i6OE0oA0K97FocIMWiWAQ9Z5KnCug9WMbmwadVj+n
/AFYbpxHrvgE1KnKc+5EEVunSaiHHltxDzS8azAcQLRIJdMtOKrC2donc2d4oYpf
rlSuykTWa0hn+NBZWAwCI0Oe2yumIQGb9kObUPnZzDsKHTQ38Uahv9vv6bw2dVnF
AqZQQhyda++c77mfOZ9YWOyWwjlBEXXA8gazEmbhSND9j4kUqOMuaXUOI/iMhcwl
6A8XAiq2PlTJ2fLgxvVYnqLd2nUQqs7UCKodn6GTUh3xKr5yjLPKwpvS3VI4VEum
JByNXFk1aVZ2fqHk43VlqMJ9S6oTkDRfquCk2sRMFPBhgr5mIJY/JYrshiMYJKAW
fQGeS1WAFedAVF/gn1TfxMj8IEX6NsqqWgJOSaxfU3nskfKKj1p5VmA0MO848/BG
ScHs2JC+Qf+s/slRfqM5l5vtFcFn5fiEBt+8AQ99kCcSre6gNsGR0eAjV/T0nWJP
Gskmwz/4dXBG5P4rNjTffSpP6hLj6kVdK6UJ+Cm8jZhRJynsXem5fg1QxTzoiXqX
e+x07gXdzVI7tAK+vsITJf45FSDEkfsBhIzcsNfTsewJ3XapsvpR9izhH9zvsq3H
21LXWAy8sL0W+cum7JHsZbs4Goy1NNldZvp1lWQpwcKPg9Q5AbaRDQTvNR/wmu88
SYordfeGF2JWVBWNEYcZm/LsoAqkxvh9aXKPXJU7LGoq1h4QOlMVw2vuEzxRK0Z4
Hj4nyMGgrQBCTHoUf/wxynVd9HtYshbnoiJ2yc+zkAE6msVxv0mfVORYQYzAtWAQ
fVRr4Zqk1EzaU334GvJ91xjpS6WBSq0v10jBO9RIqk2UMlmpyQgk09t5Zr6QSTWW
1Rswu2C26fA3mnBK7TcjdtHcVF/wRzGK/vq1NtvSlLfhq2+jQ5wrDjx8Mxd4zskq
hQyflzBBJttDrqIYUvTwkjYJjm2Jmq7woNKE8t+pb0eSudPZ4EnBbfVBW29h9119
XKQGk2FtitYWk0r49RkLQ+31gHg6LSh+efviXe5A8HvvNXT+gC0hOiuIOtoXIZ0r
DwPKyrYLkNIFn/ziDw7IG8SiwjN0leoDT7i1aLv90DGeJRxm7KgMpCogpgmg7I36
dM4uMTiYKbDqZrt/jOsdJHSxdb157WcsOHDfGS7eHhUAhlT7x5ZpOWTdkKSOmmTN
5Om4HOQ9gIHrd4BTZjFj7zuzNvxgkRHJefsLZD+WVPvh0FwI07OWzjXuOlhMwcvI
/olV7KdO2l4uz2bCuXOea6+mHLj2SWgC0fWSR/XNVIUAXC19i8fO8GwfDTYtsZaf
ffs1kzWf05RvkaM623PzpKrZhtqKvF8dZtcrIC/WFuG46gsFocnae7uZ3p5/jSa9
XvHZWbzDuJro8cMZnnVRGw3GTjNq9LTpBvFbfVtLEVJ3uq697Q8vgS3MjwSRgA0P
Hax46Xt5Af0zSHaYMc8ABbJ3gvBSM5CIGs4mmqQbiqLDudI9E1lEykeaDXndtuqY
wSDDhh3SO+x107A/Scq1lyNBcPxQXU1Xt6yeTSDA3cFtFiNet+UIQ5SKDb7wwZhl
QkLSjAl0Exsee2uVcshjvbhCc4zSLDEtIEwOZ+Yd+iScqXAx4Zo/iZcSSgJua/tD
YDu96Sf3gwUzyZzMFhvWA5vyGQr4W7ItM1tonb6fsWYB3A8pr3yS8zECklJVpJYN
YzshsewOeQopgiTHKJ6H7a+rYr7i9jpCbejnA1HH21CS6pO9OG85vmBcMn9YKHlG
16y58TTXLnAKrP9Tt6W4KmA4JsPg8chruho1JICvlwQYZf25G+xjOJ5pan4axB+l
Govhsk9aKiSr5owtPQaxwBF92CXp84ctWtklQzBmEwGxwXwqRyTqsoKkXPmQ/8vY
56/SmBuOYgO1bvNMN9UaV39BX0ZzWv0KxqsudtRfOPhATkc723T6D4GnPTJHS3tS
NdKDaDe46K7FGAlxdvDavX4Y2m+8eb0hR84bDVUJ2iuInKldIdJojQC7tETAi7pQ
ipk8Xr5Ae6lpIRFNG28VJngmzuiayzEXadRtv+HNGK6O1poyyoUoEmxkKn+t3x1r
plwirN/qdKkQmQg+qRJ7/PcL/vXliDFE0tiwYnbWFjUgREhylFQbemWxfOvsodKV
3SrFjOhgJzPJyGbyh1PMBxuRt13ZXi3pG6QLtyX6IhNoY6qfantCEiF+YxeVPZGv
u1hRQYJmESayy4gUmh/dAtDcMO5D3+WTfhYMgoWOQWc2geN7OjFiqRnebttRK8bO
5gnyjg9rHyyNwfYXAX2Knb30crwScoTa5C4OJAG+gj8srMgFG9DOaKUPqXwtRvgx
zmV8THK9x/2CELwQutEVD9CbQ6XSUW267BrSwgo6QPOlGkvSyFITO+J4sd5WWYAI
lWXcojzFHf4PuLZ+5gSv45/E411yxys68DFolkSm9T63Mzp95ktCZ2SdhwfKtc7s
zd7IDKFpdWQDanz2yHa9iLMXJrP5xRqhAODtsWc6ISCFHFarJzrDTWe/8LVYbrp6
Xwmz7lKbMngkw9CSVxy23HMFh7wTlPNsFZRlMW8vbqc2Kb1jPu6T8v5/5vSZ+Mqx
8wMZajxN+3ZcRnDIVIzgvBFrIHz2XUe2CIau9FMHjPy/rP+KpoAHfr8SjvJXYX8b
M3d1I1foyyssRtyxMewzGz1qNexwNO1vZ5qTtP33z7MfXmjGxR1Y92WJqyPnyjqH
h26GchXo9MvnvWwGLO9ThoeXpnoWvq1nwVDbm5F//nMe/6hspl4SvCMOqRh2sY2Y
C2OTtz3uEKTsrNNlhJCPrMDDwEnuSjTeMZc8Hf4R+zF6svJvkXQeBSC+LQ7JND2x
dvExtUk1tFNySwahDCuGksjEojNqsVsYXVnNlSFO+EAjCmomVOd5eGqeJ99pLENk
+VvhCUgjm4okyy7rgBrx7ehbAXHO5PzkxROupyMkFDF4QnIED05Z/V4rlKVKUaid
0tuocO42pmHzPFDPlrgQCUcEj/6BRr50zKL359kknhZy0clTOZh1BIzV5kXxY4zo
j9bHz0s3pTtWPw/wpP1X6Xi6outanVkIa2ltqSFlc5vosCAmqFIL0sv8BvPDfPI+
AqkR5wt5YrWmbxCtFzteC5bm90866opCPyOxUdi1oTPCKeXVDZI9P8usTJ2RmPO2
CLSSMlLtfe5uw4aKeInGv4m1DYrPkxa9zIOquAsGUQqabxgKdOPJZERp7wxu57GE
XBL1u4qoCv+Li8GYHTctb3o7sPOz5kkxKWBYygiBd+NryirAZCcOJLl7RNV2FtqL
VcCZcbcEthWEP6s6rKUSaGHnsFj3W5KBvCjQPqqhMW13m6T8rpSEhx+btAkv1mtN
1r8aEr0GXYagEkzPpD5eOeZLbXQ+SE8iGvXqoVERmwpr98stEC+QYYg3hSWqFwAH
Sai9PgLcA4HNuDpNjv4y0bpGAHevcF4VmGu/mR+KmqUzItoOkR/qnV76PifhHmu1
xiSYOdO+VpeR3dghFpSmSnjsGN1i6aMOHtrrSsUlzY2nqgKmu6FB10/lKk082glT
xcs3z14OgHQ1q1zqcjaeTDHd9rSWgVIChNLxmoEwiDdIG2pCOG434GHpnlKCoGQd
eBaHibnSLTsIA/+8H8KnpavdHMT/WQrrB0QhG/12Xvcv2ZQIgoGR7EsNyrJx7eOP
5hjAYdGfMk8TZahKLpsT9R/DLyDMSVXj/yepvPAj6GRWiqmK6NGGFsJ9alwiDYQm
jJ91hW0/JCSHImg6/A5mujCfdpCatvyI39A2jdMDEGleLOIOt1UKGUVaKiLJtE3F
+jkfG3BNboCZCmi4aS1pbtWGMb2q2apmmxZ4me03oH9ljZ20lb2EDG+CiiafGURD
LoM9MSDwiRnEC2GTKRb/w6E0MGWVIr7YLLTjKIdwE8eXw6nFRwlchDAQ1cxYS/R/
gBrXVenCo2DHrsWGGPePwJLjSo8pf0onHRi3HZJztGcP0HRea5HbBN7WQ0XGQZuv
tdbEZXpbdZQ7wNqivnHxBTIAPxkQyLQQ4l+IxjPx2yBI8mcK/ZYsAahpgxtrq15P
GffILV7HrAzU5LwoiJADbrhaAUhcIWEBslkldRWeyFcxPmA+DziJVGIVvZZMIeiw
uSiODQg8Y5sCtKlz8NiSw4i8tkiQdb0cmDDghOg/hD34+n08386PFQS/d56Ea2RC
rySzX2R6dUijj7MBHPo0hTmgEVGJ+ZvTyvb69RGaiAOeuyq4+dDUBixWs5rEe3V1
dlY/4P29vQa+1tOpPE6c4yXktAZhsbIkVbHAW/I5/HTpxCMq0PKhvmc9ht6MGGsC
UrdHe1Lvd2eeR6ZyIOyouW62zkxPOyuCcSS2yFxqLq+RWjxEx8zRBNVxeEDFHdN1
kgpEczq/cpOgevmOj0VVFQ7Jr+V4fiyXQhf74juBnYfSU+USEtN8QeiJB0LAvIG5
IiaW/9ZDOuO02tixRMer9hd4Ki90g5tQAo8U1qdbprq1eYCkrhmz7QI3hw+w2CuT
DNzPYRcdTw6w552ni6jlEy5aG+II/iHg0SSjbGVyz5PG3fMosr/xw+bLo/G5/1m0
zj3OJIqGCQQY+nHy/RvCCYgnEKMQ2MGGshrAgmxJvGdDt/Nzros8aI77tpmSGu2G
MYHo2CPyF3rbXmsZltihvYZmMSTtSLspJnJ8yqch5yhZ8HFVXuQMbH88FY0PoID7
Nylv5zPfGFbo7qj2j0ScZ64429JxgrM+Jrc+Z/2iywcFSwD1xlm3OOOfrRnp+YRk
DbqzSAO4xBYriPTg6BQ+fEmIQlD6A4xey/Q7X48AXlD2z0vj2MxZir0QoAPhP4d1
piJB0pYFphfvjdJ0pFLRItAwQYjI38WLo5T+SmaFQP69gE+fjV6rW9ahaXooPYo9
HpfvNfLogjit+j4+y5aKQ429qLnnQyyaGF73lcNdV6PdRPemw67bCA1Ct0vo5Jdb
CHkA6OjsFbZW9elGY3ZSiO5IgSbPeyjxCgS17LQUhGOUqDxQ/qW/M8w8ezWdy+NO
UsrmZkMVCXL2z66657hdUhSv/rsy/Cn79dFE1j5YmirEIq65WTJzWCp/OWWhQIsg
w/nf9im1sOvYoHuMxkSiqDG9QHBo7oXdyaeb36tFJQF4JepUsR6R1NdQNljqYIyJ
D7+su10KYSC/Cq3N09pztETzC+XWl+Xqc95bDgnPjFvi5eQZh8nS8jBfjtVbxyJ+
12NaWWHYiIYmCwL3Lb5f/ASoGeMFR8HcAqxNQJj/ruIKUqs4637fLKdKPqzjQDlf
pYmxop6CrnGK1f2MFXlJoSKFw2cmoS9f8+d4g7A1WDBL7iWNiVM+Jm0gJfp6BIs8
YdU5TCmch4uytdDVgS89mFI78TP/PBdr0B4iRmEs72ZPRg4JpFjv+qvvfoO8uwAN
vTL42ubIzTZD/3WynQOiATLBUU573FwoBXJp3kGvhJCkdPHS/p8N+oduFGIp0P1o
yr6NeYO6sIq74wuRFTHRBIVWBoGjJLPB8VFoKYfHsn7i0LEDD4WJoWv2V/1SYMfr
TPkkN5RBulxCB0wme+0ZpJf4go4JtfnYqkrj3t9glZ89eFQFNnIzjLdNxTk5LrIR
wdwGlkjIcOXK4NZ9MgHhrBuQSb79hKG4qtCzbVJ5rqf1J6fbMuuejOG9259CZkNy
4J333v23MTdXSAOGXmuT9qa/7h6EoKN7m4IZ/ek5C8CNfvN23FgGJVg6lFumpeQN
M52cq+jNGY7trUVZdyjAxPoD6ZMvReaDyJPs1ygETCo6Krz0vEW/L07t2uCMQNZs
ya+GtDmzKsn1QQ2cK40efWZLzVWqkvWkbFAr3iNEwEtPXwH36ZUOSd0wkjJsVKfL
6sr9OMKG3ML6aGgdMU62sAXh/ln2MgGZuJsxf0kgp17Ovz3o9409+REg/AOiMqpo
qGeoFHYewWbTpk9d4OGLYL70CcH5doprpEJUtWMD4nAGizUxJ7mjgs/oGy4i3edQ
EY7WSPlGBXY02FPdFjTooiRBy1yvfYevG46K2Eeyr3XqxB8bADIS5tM2K2be7neO
xaIdtxQ6YT9cgrr33QVZo3fOu7UzNwAanMk5rGXLI1t61zhESnCQaciI/StbTLiU
eWBWnPgmVWL4zaZXZCVsp84UT47KxaaUjMJ8YmHQ4zqtT3NvkhVlXxtdqNsaSnpq
SKM8edxrCfexbH36Vo02/DETQ9MU9lZoqHP7FpLS8upUMfSe70xpqww0RWHjoiMN
zsSIdTme8sRV2OfYvFmnwEhpboo+kJwbsUke739n0yPMbFUAWvTcOCHQ9LDCJEpk
zcrZS5BAoqnwXvzEyPRu1wrZQoUMwhSrvM6RzLIxn487Xyy3yDntjqXzf4vGzIBq
H/veVGHhWOODhlHsaP2S1XL76r8S+zL1I5b4cAaxd78nRI2QXijyG7ZPSyBM4tc8
AbQR3z1o0iFaR3pqv08VIlr9OZTMXKZNgoCPrr6uCtN1vgg3RZhz47pFxGRJTe+w
v80VkO7Z+yejfZ/tiJpAdSpkrmYvrEwLfYJpBaPILLMElvgjBECDSYXdK/SDYEDq
USJCW7XCszYtCs9bxtOZdFSuBUrN2HrfrryAS11mc1RVPa1ZbZ+/Lb8nmf0YKyjc
53QDgQA8+ll7xF3xt+BjM5T7Ct08aip1ghfqV8xWEF83b0VNmHjo06FB0P8epnI5
F26oeNpED0Tqy39IAquPq799BAw76nCCkIwfdI9IfY+t9llqOPfBPu/b2ussQM/e
LGNGUC+t5TmyKVu4mX+6oXMB9IleQFBCGYOViLoOu4s3DuOHoqsJ5X8JcEIiBmuF
iNETez4bgG6rfEky5jloQPTg8X4Z80UdFUfPMAZWIWGsnn+cShXwfpJQBK4Ut/JD
IpLfvz7QYRyu4LyzzurW+Baek9QvdlT4axeNOUIxWCmHnXsLvf7+qy0dCWEZlpdg
kxbyQP+Q0jybVakLymBgWT66WGmTFpb1lYm71uI7x63ZX026eIFxu9O5G4AEurM0
TsFZPhvpkWLrbkOKCatSj7kZreJVfh0eh0kIspbVnQ9LaRnILPNOZjML3mwUiwGn
nlj0OTjzsUpTqRAqjXKCg4Zww0wezKg/zX6bU+vvCw57cc3JjaMonJf4Ilus3LVA
OLRCFGhJLgczhxauDiW/CbxZNMlmmjiYZkd1pAtqdqPBhRvYSVI5sBfP1VSApB6R
PDK4lWRlw/7ecL704WaaqXvgytu1mHLjAG2b9fg/Qj2/+Un6lJBd9txoIoYy2bmz
iYD+Dj53El4rwPTHfG6Xe5J3eaazG41t1B0YXXLON/mHiRup6+DHjNyFxOt2shG+
le/7GHpT5F69iw0l6dNmc+3hvPGpYNCiV0SH7heJzD67lx7wcTKk46J+SiBYP6Ly
cMq7RR0zjUsC3MofsHJdStwEShOYPHnq9EfkfHGWX87Sm2hgD/2Qbhpbty4ZU0+F
JLgM3Ng8r+LhIeY3exqScMRzQTRc0gCkZ2oU7DMyGfH8gcuKwEbBQwaP+OAwd7RE
0u7OTx3/IrZZHnkeedKRHkZ18Lc6vUwSgBYLLhfcePkGwK+BCcK7pZBpfEHJuij5
L33AGi6CiwXwg+Ak1pdp1A5A7ANDytg59jmw+jHhh0dTpjZ/9IqbHO3qNO0X8sQJ
tE29MQYvneJPSgeB+5yale8C8J0x4BBc8O7MZ0waMQlwmSF+50XEQF1oVueDtk3c
fUcUoOp0f7XXs/tB+wfpC+xM1lM90V8xTHpHPQlWw3nehcWjxlnlrdQnHdAhsW47
r0v7t30tq3+fztoe4mmtkZHdXhr6+6tsQ4PCDu7k9969Bv7x8mwElL7Gi63zDbBD
5JNr3dS7cfXBdph983N0jJQRDTqQxoMGFagzWutuqOm1ZEjeqFtLD8y2MP1A2Ixh
ew2df4/Q9XzoADlO6OkEbwkJNGPh/4KrChl5eQP4d8Ttdxq4rTVm33gav6YVURqZ
rJilXdi1ZPuYnh5qMb1OjUX/Ic+7BV9ZA6Rg/FYwODY7R7aXH/LFVPi4fYSdZWWO
97DhDyIZc9GHpRG/JLRVpH1AAFkctZV0SMHgIJQfgAZZKJ8NiGLZhapD/YXQTv12
XQtDkc+pANnP5tSGJEmze++M+LwI9L7alQ1Bqnn2A22V6wjkxitu6SKurpc6iIPW
zDMDOmO5riGKo++Z27rlynpNTmQelI3zTKse75OFvz03R58C0hLToPN+C5grzMBi
xNrWYSAK04FuegaEvJSWUlUoqj94nZq1bEltJWM2J6hv7KXEY+OP53edDeE9RXiw
SbaelWbR0hXq8U7d3PFe5IDHw0tIsyCcFp5oDDPX+iFcc+4g9Twf2r7l8b5UDZ4g
epzu8KRCrJmQHWOZHvTZmiOsmOQcjn9TWvkPB5clxWRCULiEfaE0rTGgLlk+Ww6s
7da+6oR+ktDQ8RUYEFN+EHgMIpj5NLOcdh5xJ6ZrOxgrGAbaigLvI77i5LvcMWir
wdIISQvXQ2iuZAzr12ThkC1VBTILggrQdSbCJwYODKD7xnc1n1fEbBKcI08I8MYv
mcdlfgHftw/VS88x7awe283Yn/rTfYGM1RYDMptGAMkQZFW0zTcu/nFLV7WU3prk
Isij5AMsJkcHTiookE4dpug+F72zKDkvK9kMD4upHkSHawOL+uLy/zoZw6ImUfUG
JMrz19kNXdS36qmGo1It4sPwKGrcxWtZPxxaE5awA2UW9nlM4EJnI6Bgc/tc8ACO
qWim4n+3yVZI1Khe8QlWhZ1F59+zvdQEWLappR5IJiZMvmC6lX9iC3CwHcRo8Yt4
D2x6MAjYbLgqCcV3KtZEMloF0MbOC5u4cA/aCDJJ2dWORhNUuO1PyfkQGwZZVZbp
mNbXQicYQW69SVqbPLsCx3cOThJH3IROpf/oJZsTWC5c+GxD6iyLYVcVj6FxDxcL
Y/mxI/Z2K7kEB/j1JrShvOBNm1V0bO8PSsHI0bFoe+XZz8O1IP++svIg2qpBknyF
rV184F8MMg4ftipS5kiITTJwXDu3RzGU7f7nixcgDVEVN1XmKNc8MXSbwzvUHnB/
PCqrk46YGq7GZipOcdDeS0hWmtcmq8DnDmmNxEgYXGH7F6RkEGZEWZZ5e/jc4WDJ
7iamBBwflUxWrDNodfNLZDTggkMbp3zci5u4xeUXv/6QTsTzR0N3bp37SJHmeFHs
PUNRb2MACb6YEcSqIM1fVg+mn1k4wLr4mgtIlJ6U4uXf5GpqGLykMglbCjlnCE5A
VTqtryLXw9RgmyENx0U3ENc6reDs03lKNxWhvB9OidfHw8KfD4o5brQgXT0xWBWh
8/E1/oy+tpV/utgBia+BqY06QJszopBZZ0qpxyZvzSpKpzf3nXiki2EtmLNuzgG9
oJTq1W1n00iWh43bDxfhfEoOEyWbgmYyUoAleHXusqgsfNZ7Lk1c7FQYwLcqhmZ7
24fSroMLBqxpOSEVTZPjguDLTae9O379zdzUqhYXz679AWtDd4S5N2BvfVZ4t+nn
7HapqSqL9KoUf5PatvWl/Y+vvfWJ5QS/b/iv7IPnCRHKCQfCGUtzsdnqmEGvHNCN
mHmMd4LEjfKjuGYeArtuXGMxnfE6Q4fwfTocZJH+6RMoNlh+43wsjYj3YmsGTuSc
W1zbyxRYLfhB1JYyB0vWRYTIhYyMWlDTJkq62J/qJJjoPRZrvgsydyw0njsvyREc
RjbCnE5LW4OK+4GWw2CFOIr5w/MOJJGxNO9n9x6D+LYtxIiY8vY8Esubb1tccrnj
L+2WuiIKHN/5DEuOiPAWA9g6ligz8qzYkg7rkh4PEvD0BuqXRPhMru3T64a/6968
pxq+KOjLnnnIJaGs6O0JtUrp+HGzzh03B7CReXOd91vUhhfyBv4Ue8krLpZ7nWbt
+Ie8lS4gUSKaMoxJ8CxtbEYO9H7tEXDlG5dA/Xv98QsEmtKmn/wniJIT1k4QYmQm
rBIeQpQpZ/CGoFFudKErbGyB/M7G3U2WyjEOQzjovf1iEqu6a/ZMJVA16Tn0//yG
dIe0mK2OMoPQtrlbfIiILqDGXVCLorLNjY3SGBUUzOzD6/oVnHOwkr/WpL2rcfCo
00z85dwbf0Cy069gyleG9bzyNesVqracb3aqS/0HwLfvQL6dxgldfc+Z7rCVcVat
Ar5esOS/4Nhv+yiJAFvvuC3RQPTH+8f90n0vIyMen61QUvFMwHFit/SNOoVwumBm
vfNVXZ3UPgT6bhOB8bRdh1uXfPNcOAFNzNZzFaFHVGyIzzY9jQfIqafcVLG/waUX
y1p1PbqTact9FHvMEBR5xn/BB4O4d6ZYEYkZtYIJD74TOQqivlUGym5jA7olCKEm
EMwZ++RnypXa0ksHqwIulGtY4ojT4gTC+sfLdfnv6KiOoYSlhpo5+Kd38OezDIQn
kTpO0JyEG46XZEr/IOWl/ts6Wm2ybai7rIozW+ZIUJOAMcHXqMf01zuBqyrimokY
ZHSL7Hp57eObkf0Wj35FLZ99fCw0GMeS3Oyo5e+N/P978xiQTiOh4eeMjmn74kdy
vfoOdj10Hk7U8AdebdMKDs8QrDrxgdIO0rBY2TssQAJrwPI4Y6ulcrtIOJ1ISLWP
pOsUSuSOtcPpFYydD7iwHYiaFrgWBVdN/4eSzz62s/C5GZVOm2Rm8T2JpYib+/Kd
sDkMIpXX/jIiuEUPQJz7W8a5jE+Kuw2j/I7idKb7UUSLw2aaroAak//g/V/HETTr
AhrYbVZiBVWbPlHJvNNPylK71D6QfCPK1hScWAlO7OVY5XgOJupsa2PVfrZVrICw
AhDnFvhr6ma8QlDdp/oPkeacMT562bZMt9cfqfm8xOaz1f1U5K49IcqS/8jwHi/V
kL3UosA38k1hK75oDZEBkb8NNhFE6AWX1k6FpI+xKotnqXuBJ3CnW6sgze7oo27/
jdW+7cQw5a4BtpNRToIXuYTacGQE+YE1mw9REKXS7/XI3w4TLmy9JHaVLGzgrdBg
j0PLD9k8b+zg/5uAm/z7ojk1I7Srod6vrm531uoPV1jmVYwLo/Kc/4WxiQWiOfNB
g2FfP6YU4oNTtSdvYhKfI1vm3e+e9UaYVhmL1NUNZai98jNaDqa4HhZpD9niZmfw
/Oat8/Jz9WADHGZ6xmBEOFwXYBNhq6QToEgPHC2BSeO9l/viGMPW/7PyTOlOJKgv
+zd39uX5JYAJM7tEbpcNWxNpcmlnKpI6knNSgjvu1IHrdz9gdABB7+PknDE4Ue9c
5ssoSBWU76NJTe3HqUH579eEuoGjdqAYkmQfCb5hLMkMIQzaXNH2gG7QLf/s0iwb
t33U6tP13XrLoElacd7XEMkAH1/gDU+SIEkjKsEF5vuT26LHUTzam0G8wkKXNN50
P1QkiKBe0dA4/bdaYBFJAkqVTq7VPMmTK6htgQ8SWZxwo6KOJSq+eBsvE1iLV0gC
x0yX+Vu/x68msEJInxuG0jLZkYdShfBw6jVR/I2T1/L5r2PoJcNTdzZG6Kce3SRu
SLGngkBktw+yyAbw9wHUe71QFR1R21WkqBTLOBV3umLy/hnGwmRDjbdl3xccCF4F
4MDzW5W0k3DV8PU5B3IOyE/sCEQWXW8zQqxz4nEnkPFlZN3YoCCJavtVuvfKqIzT
GuowkfEx18Qd7PMwOTgh0rrdjWu17q4KbzpyPRQdMCy7ci++LC5gQ0vk/wr8m1cn
kYPyEmE6BIQ6ovd6KBpbvQBbnTMPMEMGMA7zM3t++/sq5pSvU6PvBomLCeR8im9z
sIAEqa/RekLfuXVWQ4sSjVWZb+gZOnd1KCMorzafik9/bdXFjFS3Dt1XVSRqM5II
M1Fx4HTFqmVdx3JZo2a08B4jEVsxRxMrXdLSBuojKH1a4wj/2pFeVYmzR379aHlv
uI6bq7fcom25kAQ65v1iZphs43EIy4IGkQO32FXMZf+NT3oIYmMxIJ3WxGed3EK6
Z3flEbYpGbemNMqcselN1ykhJ7XgK8oh9dBqvIY3E9cCFCD2c8k6NzDpO40L1tqv
AEAqbj6rG9C2bg4xG20Am0klYJ8OzShQWRBQc76OVQYlVeMbydZmqTmdO0b4Xpcc
L7QVALvLdrX91LV3uw3etvhsy0u7k1/ARrxEibK0eU+RYM5E0j5u6UcJiF0RRUig
7kOdwdpwIIsWZojmzu8aqqAdINlrmXYa5ByQYU+42z040AnuzNNWpBvJaM8W1G8Z
MRq8nh8n5eC8j+uggft1P/AsamxWm+tAf/6/hJQpB+pPyRJPTnl0pa60CsHKjY3Z
SxfoSfsj98ohY4ASRpwLOJBKmO9fcsOj/Tf4cICr8NTGX9T5NUDLnCBBdjF5L8un
IpjJ70fYdr5kHCRkhpmza81F3sMhCGJfoB3LBShYTp06aFoa2yf1J83n+Anlqw9S
DkGPmX4HwL8M70I6j8P9jFW9nnAub7S/SpHm9mGo5O+hydSILmCAM2VcFYJ9kdTe
LUzeR9YrfqUWxWypO+nFWqbTlJVqNGZkemHlW7GHBuMI8a7tRqI/nScaoEg3M37C
vnFlVw6eW1IvTXi7tAnNvO+E28QgvWzMw2/rRqU7p7w/WYqF2iNu+lw8Ew1NBwO7
C8MnDBdQPu7XFEBUqxJCOhWkb1/6r4tY5g79fu9avmnavbeGq3oPz6dHd2D4GXQE
ioXJlNaPkE10/IzNYc1SxBORC4CW+GMaqPz41sWT0ZstCpsXh0IQIFa4xuV4+I/F
HTYE17GEzMfBjgUP8yWEbnrnUCLYX+n+opnx20bjPULAncAHETOZn42Pc4DGHJ4H
PRxf59SzrtGXT0xqiBBPlkIZmynqUP1QkOXg9wxKtrblcjAlxMZ+ga3RMzlYAXpr
p9nFSBkizEre02nrv9ZD7SiYpHPzTwA8Gh8hNytPCOuh1oefd60Gla76brisbQRD
17CyZkg+GqL7TS/1JJQjLmBOkloLhi9VOArsTm62hRewOrh15gHXJamcaGFSQ9u+
JEEiVTVGFxjVkp2c9Ou6nQmWQOc1MDEqeOiyvPfLq1s5Q9fS+teiSnzLWRG88hyy
Iq1MDxetIZnLetG59RtYJvCnZXlS48l3+1jmoDCe30SZmcwhcYM4dMb71EAphqAp
EW++XY530wLwnjFKMqJHs/N96F3tZF5A/IuyS9Pwkn5VAy+db2b8tOp7OHC2qSer
COFkeZ50bjVhXXAp4HBCKHc5TydC6186xXV7JE/cQuTJecKLcRGBM8KQJUxJu1EP
NCTtmOATuk48zJxr7P+JdBiRcLWRtMkCOyTno8QyCEYS98Z7puI6jiP/nDCKVADF
z8VHem9N9pUSqkNVTnQMxCrg4Ev62vugdR95AupBISxk759rNJOZzQDXL39Wcd0d
IqgwMQgod0mYBklKTiT4X5n7DhjKiCq36ALOS29BSfQMSRR1pZEZiBYQV28ORGIV
8f1dT35EdIbXBm3waXYeBIs1LcErCiZO7Yyw4IQFSb0zMUDRgMQDeqhZuImOKMNR
wdgjx4e8Ir6PdJY5mazqDFaBC8VoZgyoKVR4PCC6PdZJTRhsuWt+RsLae9ehtkoi
pnua87G5B9WMM9A8gO4VVSDZlu6xVOWnIHWP4+FiV9GXqtgtXVQoNqDsSUbyeufy
6gsqnn3eyPa9BAz7+yCb2lYn7UG+49+uM3OHDkWysn7IBWhutBPwkaOq8fIzd9pG
jdk45+2MWxn9V8eQQ/AqmmqLCbbDiZGMGo+O5CpgwpiVvdKVXudaKwJjIOC1q3Zb
21BLq1ZJmEux7h1tWzIas63ky/1d2ATVoOquwtOnWcK5zhoHzAD030QOFRst0wTV
XhPfZVxTPohaIOuUFkJI0UNHc01PpdbnuF5Ylja2XhyhybW0JTSJ/j0ENwOW5csx
41AW/NmTQtVXaR/RA+YlbJS5a7mvHG441eEClyYYb5ffGxwVBpCSWT0zOLrbWUBu
EArHHiCjP4JRPesYkQOiCqLVBxjDAxL6jdEOxPuhWnQmm59zCWQx+Z7lTEYMrknG
/vDqRrdwxsAdiyfIeGu+gnvdKYPEOVYFKFV1bUseaFTEC4xLMdEAU5CuwDnb4BAT
Zj9SNsdyK3fRhJ95f8dtncXWGYkwE9PFvCUx+1cQwT8k7jSBaWrrTF4yW+4N6L+O
xRJtP9QuCW1lOBgkaI8ie/qeXOd6PInMhG7BpZYRz3g33cVxYdsKvvIZiCz5MCjL
LbnPxtNLC9Ov51tcloZnV00mY3N8ZNxspV/lczbJTL0DWohoq9u12MT0szvRzQtZ
0oPVBO/88WK7+cdftrsfzOk0b5kR8n5VxkHEV7Pfz28uiC3jH7jVhR8TORlLGXWX
NdQ6R2cUUMF+2xHYSwL5n3b6r8NNCLeOwk3LxwCvjYhGRFW1EVDTAk27+MusXLaC
EAKLsHatoizEc9iBt6JD225/ocFPWw42/eGQsPwAmMI0N9EzMv87e4O98Dd8vr1R
OHAfdTaIRJ8uCFg7BBbFjqhjmQ2OtWewSpjncFXCGAqp70hcoXUjUr+ai8RswEl/
mXpJBwDW9E0JV6vKAp+SltQw0vf8ub192AePD41oP6bU1M8EGD2PoagzkmezWQC/
w7N1/tNHYNcsSlVkXrx9rmVmspN70VHIwH8IFv81AZiUWXT1ys27XVCk+hpHQN3Y
8HdhKSQmwZkzef7lcbKr71mlo8Z3HfiiRXP8ymxxE9j3ypoxnTOv9hCWZQRxqzy6
LfrlGsRsZojBTcwx5cgqZUZtgN+ewcEzL3tHycji6xXhjN61oOIKlRGB3VPsEwuV
yQj1lmIo7rf46igndBcs2DZUxIwVyQdd1mPTJ4YWAoFdhxyn4cJskBmh3A486zlC
db2erPoCZkTcEV9yRtjZ2TZOij/wn4AZ5Pk2kwhOircQ/UrWUnZ8nTje5c99JkPF
KQzNEsKbYc7QixoijBTmAdZPG8Nc9eUuOsJhSbltWVwKvyX7R7+Hu3y+cLHlaHPK
ZyUnd7X0xeb8TvCRwChUuBnZgCxRBLHqaUdUxo18dtFixIWauyywCDJDzOqTTOVW
ocPvveuqS+iOOetha2YaGrPLARn+YoQHpLH/mWKb5MPy7r3mqVMGS68X7mQYkcYP
brVmK39EODf0UZr6piFA/csvmPySxnsVTYTMB/wWtlsVckW6hDtc69UK9ZRgFe+X
Uo10SOpH+ITtkQkCcTqKvPmAJjxRdnVlVHUapWhh14SVlA73nxqqJIEClAPfguKi
3MW1ecNGvmZcoZuT0nuyGjqQ4Skbh3r6ejN2PcW8YhkxpcCyOc2wsCLOS96Ng1IL
B3PZwZ3pOu4PTaHvDP1zrB1ImRmjCOt7vnVabfLbcs2XIzj0FO85DoRqGWOXvK/e
xzBFb8v2RgCUbK25w26M51rJojQlvvLzl0Km7jh0di9bQgexk7IpZEfbLxhIpZsh
3cFkcSdvW/5t0CAY8WA3sod/HJxPafcX8eCN3t2Mlaj77yMIENcIGbSFPLd6nPv8
iHnGwWtopgkkktuiTbYNYiBud61jMoIAea81cZLRQNqf6qgaVkzeL3q9UairXNnP
08/5Okw6wMKCZavITO/fRF8pmXZ00qORhEctRYxof4C3EA8Ke6hoSGa+EeNp25fS
wNKsWmOi4RkAbCFduOvjtBNRUNMWiX1JNpPv+hD6WwEdgb0LYJkw7SbqxsqFfqp8
pLqZmak946AXKUdRA93ODGfJhKcYnMBOP6BZe1vDlxC8VJt0n3jLskpuNdUs1tXp
89+Wx3xXGvOdAgz7FIdvok0IY50RloYOrWc6ZzkGHfB5eE9ncOgAM6rsZWxnAyVL
3IhJS3EnVED/zKF05X1RkruYOAd6pvfobdZ0P/UDQ1RJEm8cU7WvAwwT4nF+hOi4
SAQoS8NIRRqZArAs14gqK/IeFYS4nmiMpSYFju4Giq7NXgeTAARwKGKnJAMSsY+B
HLbrZUohouXVs4bu+qQlLt6JyI8HtuofFAnA1Rmm2Wohe8DwJMgdHDBLU+EGY27X
NCDWx/o9nYYnxBKfb5yxMaU1na4jYkVFE5IgnIWU3w1PqYOPYJb5xZslZjvmrwjw
EI3gWbfj4a8fkp0e7443nykCk/x9vaSjGhM8J+cxhyOdLVmM/x0JJ/yiK9FyBUed
XpuoRSy1WqciX6mGGkBduK59+l23MB1gOhVW7LMqABvU0QTFcnLxlBrQSNX9oteb
GddzFdunIdnJD1/HGtWhguciMGTxrY++VDf49HtLY1LqbsDE/5nUN56jszMyezcl
dv14pWfbvsnt8qO7OqnoMq+V9O0IZS6dRA93Sdg1wW3c+P592Y0weMoeEhpt3hH2
dYtgMtz2qz+XQCfJ4mFjUz0lkXYZVrR58bHlS4B8aPoxq0BqjRUt7UFgTyz+WndZ
fbf9o2QSDCjKxi2TDtTUgr7RTqB4keUdefrJu3Uu2Rk+UvxE/iAMlvhNhbURxKZ7
qaynWHfLSaKfzjhiIVvS+uaYEN40cZhZKF7YSJFxzTlbx6LmvzvQvsDRLhy3oWkI
aD7noj+ftBx3QPlpEbDrB0jpVb8uxSGHPKwnqJ1Ou2gzNkSiglTxDv5bu39HIsGY
BE/7VWhzAxiovRcJi4aIpLFGKv3a89YyBlwTi5o8Xm31r9ksn64KECzid9QQV32c
z6mL0CwumLBvRfJlCfy+UMkhHToUTpkCeOgMAiWRatkFxyPfRSVTEcufdjWMfMRq
+SopITdqG1o1Ljf2fJFlTs51+VKj3y1Q2IoMNnl98K/bFB+lHunJl+M1yurq8KRg
PANI+8wqHKSTe9ZXn4JsE6ErDoomMxBFPy9I2JPEbp9UE0Oz4pAwy8gEs+rv7zcZ
0BQeFCFYYMw8S8E/C6DAfH0fQR0f+ad9HhAcbsttdBBGYcQMyTcZUTtgY3epC5rt
ZIKuykiM9reSZ+fbSOV5lkFsglAv4gD2mT5L2p6iEpCzmb3UfWfcIVWRV/FlsiYf
7Tw9e3Kvov2Fr2P49a7PZdS2bPtjnr5TS0X/l1AC6WzLqYY4YaZ3n7iA8dDlirAs
G1Hmi3xDpmjPJj/b31Ymn4rMvKKIPqfQkWDJB/FruEwaIjnsg35JGF6AL2O9PwHb
EbmfXwo3GcNLKkzw9oop70r6WgvCcY5dBpFTdi6M7IOxUB8pnP+4xGfO431GNd8l
mjnmS6tBcxkm/GP6rE4FUg1ScLDT4MQj8LAb1EVVmc+vBGaQYFcwp6Y5VtI2qWtW
59KKKNljZpgqdMlUTJh0J31sW5zOBZzhsOwnlR55qIq3pUFI86VDkepxSWRUawHZ
BqjEI27gvvn1Mqq3P9ctQY+se6tCzAFNV5wUdy0xWgJQWUG9gdKrtf+ljNHuqi+s
ERrYFLBuJTqqnZ/a6jLIEa2uumXn4wjl3jdQKoNkDvdlOYmBDz0NQ9yrpDOBITki
V6BRFLbBrR6pwgKM6Y4BR7eOD5O1GZxR7G1lQT2JMXrfMNsIcp9j5CVpaTBFquDs
T4yhtFh7AJRlw/QfOhvUm8s5Cz41YJ0oYMdQHO4J9tUBKNHjoltNnI5sm4aL6Wxt
CH9rk12WpISnuirFCsO2laDRUdEBPfgyOQU9Vp+UFrJDy55muGHv8S2CoTOsLASN
qiWYGD6Jg3QcDpI7V9URbpuJd2yHPvG8Q43puxwTPbp/MGNz7wYPyhh231uwLhYX
0oTEnUIgx4DaWRRaL4Wf9fbIXAFX2XWuKmk6ezOe2GaPCLjoEKWnnjowSDfUTvkH
NZvfPy6I3gI34s5/2NB7PckQzKMVk+rBz1nI2WwfYMbYN9GnVH12UgUU8vnoJB7d
0uiTiWkfhhzhdOZrpxN/aaGeBVxfya/L8O/gnrHylvbgKfIoSStNsTdOC6HsQaQl
x/XIudZUWQOoW0GGmvpjvuNvpWrtqX+owKtQrnS6MpFUZ1KtlT+Dr7an9lZsi6OR
b+xlnqOYCka/N7mVA+Gvbm6VMv11i9w8TvQ1KBL0nitLNnYWORaa0NY4dzBjGnri
xcSXQXedfxTC/n6D64G2QHSi/XwxHG9/YpaJVzt2lT5EUjDBcl6o7RyX2gFS0cSy
gJzZEKwb/OmK50t1xoWr8Pvfk3D8fam+ktZlwHuLGSLPF6yOZpVOnl2r11zEH5TG
cH/3yq+ZgdtEevDK/y2XvYcTd31COkl5MVfEjrPU3CbwkaTAn3xncCDfza2wjdPk
OMstzIW9SMT94/Y/xX/tIisn99eDFejgBtn5DBxqcN4uoet0c+50ifIOptA/ePxD
D6P8NWPAWAhIPFbEnuyRd7v8p3QYuUbY+en3iYT2yyHi937mMkj7oZ8RynOXSzoH
xn/p92Slr5Nla5FN++nBVHjBV0sx3A7MsL73GSX7P9ci9t4WUbFlNVyO/Lx9eIMj
YAqA66TUdryRdhjS1ZUTp2dEDdqr4MPMLNZemqIc5Ho9RDd8MiRoGxcu+LOj/vKD
237YjNeZbD147/xauUwQWPGjjWVl89pqeVthDMib1HMFK/7RM27oHympTOaP1Rc6
2a8fnQ3z+pOGDYHBlc3yvcJilZD6tcBVA+Uwm86FpVleEOHcw9L6VVus+8dI9+XB
3NNJwlcFlqF/Gqq61cK5wKcudopgc7XF0JLT28Rs5yNTREmJPxa475QsDbiooQJP
BKWdIFj5VaSF5n4Q0JctzyIw7u69Qn6tUZ5xWUZzXq/BWJF+5+mYOLqKYLBdUPfV
W6Qu2gGwyfCoCKmLUUR4DW/ySIcBekSDxFvtg3dBNpsTJeaED4qLbTzfc4dy2KOr
21eOGT8rokrKaQtBc4OFRjJTRvbeuD44dgIrSnKQ6E2Kn2qwXCObK3MVSmHfKntn
mBQ86xrCnH702FDQAia+zZdSd11+cam1K8nCJgo7kIRyLGeCcMj1W/iBec97Lp7i
bgB4bTFwYkAANquoOSxH6u/l7x1lu0xNhiT25xJ1oP0WZQTWsCsyV9p82nHemqU5
goQ8/GmqGshP9Cix3GTHy9dSzcNqlIf/b6JDBSaSZBeCUIj83Q8DQFuZ+e6s/339
wppR9ZN8mrw0Sx5tjmI44KAH3aRNzwoWWdI/JTa/QFjPFYqZWLVPub/IcnngemIh
DHwMb/jzxMjceA3As+H2JxM2oneB2zMHwp9nOC6QSTqT9WlEBP2UZx/3OPwxsX0D
9xjlYqY7QSp97FYxoJR36ShBoZ8oRzf9nr+jCy0BjINXoyFj0vYOqf7eyzsjU6Tv
bcr7b4AGDWu+l+LoLxDyGaTIkjUc0E1sfeOCREYby3BDBjVxevuBxjJD/DyXtQbH
Tk9apDtImPhjqjQLNvv4HtSbKd0GLlGfqB5r2dNHFfIEH5YaWfmUcpQUcnRNB3hW
ulq8oLqEVxPevs+msEc5bou1va2dHobN4ZJmcGwmYRituQ0Ch5jRLB0qfxiJAqRc
E1kBZ74Pnbco7LqcZy2UsPpZaEDdMZu+G327jk+V2zmJMQ7l+qmy2QKQI63HXcp9
o84YmUrEc1FReUstTRpti3MpJTnHvpZD0PG1+pPCQ2JiK+RoMXdm4GkFa7ROP6hz
TuXkZ5ZC325QfLWY5K/TTwCNgumhHX8SbRPxeurih1FpGV5b3Kp68H60m953DLer
mAndqM126YDSl0wDTTvm5I9sSuOlK7Y0MdAWbzkn25aTca+ftGgJ++T0HtG9ezUx
+1uoj41B4QSXzjAi2N3kIU3sf2D9NJjTg1Iodu8L0fkYs8MthV7QIOpCye8SHs/5
FCxz3ir8OhlEhw4sbhIXqyARRGNgIT1Jfb/C/IPKNUohHPWkIluX6GJ55+4d1V/+
ZOAtbfC/2McjmR0T9Z6LUxgTWUNVQf0e71tOvRxoHvOrmEFwFupOLJlqdrlop56V
J9CZMqXOH/MyvgxxLoyT+VyJM1tPMMjZZ6WVmpP9BFnRyADozhLucOI8pwqC+5sP
0uV0s33a/ZWKE0QaeAqiYa+ANysMVLe/KF+ue1EVXestWsS8ZO9GccUwZczemFgP
G0qCc/48g3Skuy+VJ1SRjhOc7utBxuvEpTvK3/Av4T0oACpEaT5pKwJo0jbhU5UA
PZ4scLjGRyUM6mj3a66Hgz4aZ7iYhkFqfCeZM4gmvZO0FraGfejX7hvOFh2HpCGX
Y8OHzeMSwNn4HqqfECUhlEFjiO9s9DgZZKL2NVqhj0S6fqhubKC2e7B0tFYZb2Uu
YjBtsIQAnYI9Depr8B4S5lpbSXp95/7r4IjMuAXpjR7s9wsZ7LI8Euj6isAlBVc1
mC0/T5Za0yfwf5/JXZIPtSK2Y/WnhuK35xQZVxHDDjkKVM3cBU7vHoDz6/u85huS
vERmbzPi5LvdJ+rNF1Ud3U+VmfynHSyMwBALz759fHVR0jD2y9iQvfRcWYp5Zs5y
MZifE0SoedgtKfSKKJQeJ9qi7K9XG/VC+AZsqWqjyq1Zdfs8F9jgtSjt70oOymBD
LoxarsJOW40lrkk/8kEoICe/GdVFcIbIg7QjVm1U6ZYshAj1Zs7q51hSxSTYXEdL
WvyDHbQQBhTXF+aKOoZV4Ymfiwh+UHuPzMlEgfv3HBGzcCLUtHYtcFVvG8uiqKJ0
VdM/IQQzMhX0BgKoRbrsGu7/LwnKLki+qwykwP+RgA9Xt4NNEsLvu11yRxXT+F8/
PvNhGGmAqsavXyljvxvGnD54uQQ1Ndk5Z4MyY63TbqeoJOkx+X7AUBIiJeVfq0W8
5iL2gH6QvsTSAkrvinTazKNnwNmaCmWaKPVDvWVHi1wDBaq0yNDhJrfHeFDoHCL1
YcTL/fKkdQHHEinT+hBAgaAGHDt9GA6VXD/CEagvuC24HDgEmZ50UnHrtIbqwLHH
j0W0w3HXfszjrTKo8UO39Ky/9c4utAuJPCCNF61kyxIaUS5QyTIjpzs+RIelHOzZ
m4ER/5RMKLNkd/EkjsyZPp3thrqPIoXkGeqm2XoY/veWmZgcPLCo+FDbkGEUTXPK
kMwNSEcgYnZgO8p0l5tamFXOcnqGHsInhMXvMVJnRJS+elFyxsDnPxKnsljgzcQf
3CDZJ1uaymWh9CyB2HCidLqFvgekN/z7bAPaOPCQ690KmkmOQfnChfaCMossA9DS
9OtFVakl4EoR0gb3ieDjUga2oY3oG9Ki8BsZZ1riooq4e6IKye5QX2YcoJuLzHxT
QcYUrFJ5IkTEVKgc1AaXk0xG0Zw8KJFX1CpT7azuCO9ussCDK0wnySVYAqQM6ANO
gxD0nY8us+fu5WETUe3oDn24ZgdJGpeVS4LELqRaV1ONteVF+jmsKVP6crwwXtGq
F4RgOpWbs+JfNkQU0S1ZT0cXhSuA6oEotE62Grh0RruwWx3iDtkC+KWY2qVbZLAo
cjISHj51sb3j1Oxg2n1Pqyg8slM/5+T/K8y30NuPAKQO2TWKR9RVJV8h3D7vXO+f
UCKO2FADtrfpXtT09313DYRiC3eut9fe1p0/tVuBLWGo5bpbzPwOIXvRU7BEwsVe
EyZ5URGghL57JtnvkcLrdJPi3VZ2e2kGPo2acXOIqeby+eIaPpvw4C1VAnyQdDaL
5Q0gngJ2mLFjQJVqkmzgRybkRd+LPEgB6gqS/eTDosqwK+1MyhbKLhSf0NOXJ7YW
F+/lKvXDhUzaZ8oi75YGvDgk7w7z9e3vjg6D8VoklGNWqE4+YQLXi6cYDF4EHkf6
yqEUR98tE1PexgBVbwomEHji1AH8+oPvijlk57TBmU9PEU8hJrhO9I8lF75tgQSe
W/YXD+jBFH0FMFCwVn8e1DKNZU4XBbVliRIAutwoAlQeYhLKqCfxTxswVVOlc+iR
ci6SP1RDe65rKh1yT03963HAEYx9GE1phU0pjZxzVLV4MosbdFJwvllchecLRrD/
HrUL2k4zqNHvlLhZ1tuAzUbRw8eStF4umpkyNElHc/XjWjvcg3UqajxJF/bCoGru
EO2JkmtcTkkutgl/JgtinJB5KbyUoiK8qh0kqs16tLvzhzSgzr/Qv4Py901gzKYL
JnZeBd3KeYfQp13I5UQ2KRtOEIC2I3VNo1wo2mlF7/YwMvd8QTas1vqnVg+ww5R2
atkdM3+YAkDLT05JbsUkTKU4wOmWaTjlCVB/RQUP4H15x2Yt/htT8uVxR+DOgZoQ
1ABNfkDRg9/RvL1Zb1EYPW6dG5qobaoLAZzfm7byEWRYl2tXqx33nT1Kiv+RMlcz
x0daMZuL99odj1VOFKa8EWyIyHWVxBUaMWlUZ1/tjICP0pMmdFEirNNUgiz6PsYk
AHtc1QzlId/Gqx1IcADlMJj5vC+OEHzSZBGGHvlJZM/+C6U89zwtQ73Y9iTYUMEh
NqEDlNVthONeZ/5Wz14qu/HW3+xcWlNIveNU55YcvqJOJXwbgNDKexTNgYLnPbdj
I0KEf7GLyh+o4mMQB136szjnGl/dI009YcXIvvyg7L6c4mtoeE88RmHiy0gzbGiY
JbTp5v/w+9E1S9uUfawsFUdmkZW2YphND6H6CkK66QKyG6y/ycDn4YLQ8AVZTPet
Q9J5IEqp1g1BFOVE++yLXdAavgsVUdHUTaaRxnFiQEqSIKXdnk9HP3XmSaakSHPx
aFMbNVqdTrPPwlz4+4bzUxKTW/H5Tp0qWPg+2p7Fn2kn0NULWdG2Y47GHvjJ43e5
eBi3SJOXMt9ZyhLtLq1p+q6T+jtHDAjernM4mJABBfcF+x3zOToEu3l282uGqtCF
m6Ufi2x0/7y2r9fCoKcobDekI9NVUcNlHL0g6mL8DjhvywCdTvIyhDXpRWvnlSjy
4nGfcadIczzfS92KoHR12FOM5BoGbeoD16bNoxLpLIm1s6Mr1fYvFlc/ixGM94W5
46FnA3Zl/ncJk/TXfcHCrKTyGZY3NQRpLVtLplEWLPAwC9bL6jWovEGROQrw+mg6
N4mHVbc4X8wviPS/DKyadmVBAQOIP9oVTQLqvPW8NxRvDog8j3fBSAZsF/6/Wkd9
erlNUh1F03luHfdcj3IFaFr/QCmEuYpsT246mnIZbBpbjrDpAcx05zIB1BGSpEwM
fpNhDXIszPubVyJOe3xAHgEu/yjsv8AxG6cYHv2LdYytoOnUdFxlCcKhTuDlHmUx
fl+fLksLqnG3yD8A+Z3fg7UTtIFsmciXTGWcO4Ge0e1Uf+PjMe+nCQnBhfqGhwtg
q1A9SHNkzgUA02Lax6TYehPMJ7gpji9zUtyUC/JtwWJfgs3ljzltW6Q4kRKM5imc
QAp1hj8GkVn4CLf1w37g/4Ui56q9x6L+RnnYsWpcPr7fUIxgUtofTEZgq4PW+VU6
iYHu3RbqaxwO7JHRmqPxqR5RVbsJCYIjjd8AtKIptofRyHwOU02HiU9ZnTQzhnSr
X0ouiLHNWL3+R9bM9a4hpMf2W6YHyq+5/IzCIDg5pswP1rnt0b4pwBqpeffOiU52
aj/35dmszf4SCM96tqJp+Jjq7PPblEn7uNo/SHrZg53+b6vi/VbA+4QP8/7ebDva
zcaSe9/YTpKdMI0vMCp66Rr+Q3BoXEL874jRaTYlza/e8VxviA3iutiu5RssUdxl
zr6xCCglNLi9IOENjBA9x0ybbUPBZjBsWsSWHV9lMW2oyJf5Ma313FVqIxZQHItc
3XdQdCjOJC+cz0/2z71cZKgsEEdG3pABH2NlDTQM+JIIeGyGKgBuhs3VKlXYh13M
Zxm1RYMl/+4EyxGzEBJOFMUHA1Bv2wk96cM7Kt0sjjkA2JJqFhifNEbY2v8XiwXw
3i8oe/KwAUVhRC60v1VdbJEcdKAPwBYAVlM+SZVEakkUe2qvFuMTsDtL/wfkKHhs
M/xlot2qAS7eozsEExYfy1Cqr5EqkIv4s9hT8mCIdEwPQgH0NB44a0IzDMcJEFfw
qWfK+myRtjmbhinL6ttky5VJeOMWxtQXElN1OWIKz1s63H3OEEDqVDb66Vnf6U+R
mLKeZr+qDkc8b84L2O38trgsv7VbeXee2RRlYBkPN0MtxsDTHO8ksMYVuq3/koLw
IByusd/AFMNX5HpqiYC6B0OKsp86RXi5iWIQF6knDIBpLcmW8Zrkj/dmOhhR8TJs
unJ0U55yzJJsOBa8NFtHpHATGcnbj/byBKWCjblU75mxleqBiq3TBESchCbkret0
9tren+uqoXVQJG4cnZ/1xKeRzprlN6rDaea1Rcy2Aak13aho39X2WHwmk2XI1FeY
XGLcksP0VjgXmja6wbmfJu54ypVXrv2gEUVS5ktSCVG2zD8nKyM/zC243MiIG3mt
K6S20JSaBOU33z8ODrsmoa6QIBSfVbupniv7z7a9/gnnONBr2N2bxJWnZmma6Tmu
vmvnQ+FUhegNRsAPMfImiBwQkw/DZZ+ButFgpyj1z1S8A8EtsOH/ukXnb/D+AJGU
S8JwjO1cml9t/IVMYlZybzfL5JKRy0A8PRYAOkb8hSsglaaWcFHSANPq+RjmTdiD
PlHyLPkcd5kRUNzgOZ7q7yl6j0qSkSI9gJKU31W99q8TZgN6sGUTfjpQ0upM8Pjb
eXCBGBtLmhdMghKU5diUYKxrRtaaB5pSnfq4JDdT9cZ9Zrx4GBwP9En9gqZqiHWD
6PtVRWgAa6D6luB55HGqqSNYdKsgep6vodP792IuXPvHuAawWMnjQBHjvEFQDanZ
GQmfslAdP01Mqv4u2jsuEKdmnZ3cf/8FpNf6X8bTUbtNXzmqW6zDOemuzolXanF1
KrnHlDGWxKYl6KJSXph75ppqdKbE31iKoF4xmG6kw4vzPbcF6dzUIVMCimxjohRq
Qmaonri8SOXyPItb+QCVvjtyMuViTGhwWk1b2wTbJKPkfbO6+jLJsJAB9VIdz3Ux
9tnB5pmcVCCShOwPxNJ7eqIcgyrslElQN74rVdOROQreqUMqDw0S9qZa7t4399Yd
Zafh6Gn+m6WHYrfjR/sUJZOQq1Qgu9eVtUkcBl/i64cSoi8cmQ8DntrNdvyaTata
HzvOXQnNX9Nwa6iuk+k1cl4aBbJFmRPP64Wgs6bNv+Dzn9NEsRhMm1p845cOlOCr
tKwR3fliDCMO2nb4X8fyjDRky3aaqckA0tnsxnFsDD8zZAdZFl3h2ybiDWvOhD4M
jlr0HC4VUQA8PZdLVEIC0AN+EKK0DVMoDasLXhBOa/YQl+7IdM8TUfO+/MLitOBO
XbAn1WY3xPCfirUualtRADHJmovuFIJa6jBIUwywySKECNbkUI2JSJNvxM7dbzLW
KWK4Uo53iIhiClFEea+UBtsJ7c7Q4WHM/wodxJTJtDWq2hB03JvYeL27BFodL207
nPfowoBoel83NtOY6xWAkwsbq1IPNdy8qdiv/fI5dbpBt8e9f7BiLFg3TNXcs/Wt
/oqkDeM5+ev3XuQv2YDGWcD7Z85hZMvuHnwo4ybtH9CShFEUfnk+9AhrG7duSOyM
JLs+DFxS2PnKUzmf8/lB09BFrRYdVv4rzq58JjWyllpQzNzsfkX6Ot4n/SWKqCnY
y7GUjDG5WJUJx9Zgd1EYuoR3dISioEaZkhErTkrS4IP2l5Y0rhtmX3/Tix35CzCd
K/ERCQjp8Fs5cZumHCUneyI3CgeUB3ODOBR68BsSeeRSzmmLEO2D8su2gYL6S8MA
nm0h3LJVLIc/YcdrGuWsyevH6ivC0Ry1QguLtiDBtlUQ7XmuiiWU1LFlJdGZX5oJ
KOTvRTr2XnxioVg+9VFaf6y7Qs1mB6gTYAxyjYgWijcWgLEEQ9TlVwoImt9uegKl
1ZrHRQlTOYgYm8qdyKofHS0wsXCLsg5twDGNxQpIJ7Uhb8Jc5BP+j5IzudXkIaWt
+CsuKwEcN5rQ7YFQJmL8WkgPZqGfBgCdnVCJnTQuccYS5jY7G4pMbHqtRXfMYm5X
aEe1IlT8BaUEchS1kYz44H0XAqzhaGqPKS4jhvolmyynkolBOkaBL59OwLpvrlun
85XjZUzVb2GQluTjtQ7W4hQea7Y3LbfyX/oteW6RV5rOaJiA45xxkSvUGOOzjZLd
voxq92ax/uaP6P4TuF77eFFDUpHhwRdzzy1JI/gEuTxlhXVXS3JvWVP8lJPyssgq
jv4xfYZZZffEyKXxRYaWs3Qt+gbyqpRWWZuktVRAgqm6CzHU5FPn/cX4LUbVDDiB
MvAFnTVHcwsLagvmmpcwRCHqKzKnlCexLZUyvRmCWmKJetvc8qzeN3REHkqiJg6S
zCnUegz5iqR4eoMjOpV6IjjAlHFsYcjn51Z4vtYpyqFinHxZUiXdAx8U+J1ThD6B
GSrRAoIHA+FFV7cIpbMVet6spLXRq9prCADdU5kbw2KzQLS4AqRkxnG1dX8EvdXF
ftTw9nQ2KoMrNd3GRKqCtebLcMnb03pyfn2+eFaDw2tIsXj3swUfkO+oZ1uTVWwF
iuRAxXRopAXrLyt9490axDMWi6Rl30AwieuBhFntRNc6XEAyuejL677NxIaxMPK/
IPFmYV7WLUBMABhF0s7fDHX+qscC8q7XOSY/8CcMXg+gza6CddjxJeJm8jDUeTV5
oc1Hr8loc/QO5XX6DftGDXpG5rvUSUliQFBfpe5NpjYm2fTVKACdapmQ1x36kl/D
o5VlzG+7gsTGbqCyZMKiXDFb15xg2R3+wO3vADkQgatMZg++nMdKo5Dn4SptRHuc
n+cKa3eJ+fnK+AE0lOU8JVTxpPFs2n+KyRP075WgOXOoUycrBQKN7RjlqfcFnTB9
Z+6C93uohKlZ1RJYAuEMUFNljHsUgG6MQUSxYWxSCsCLi/m4Ti0Ae5ExLXZ/ssks
u1aDF4dks3rhm9uzm1JpE+P0fA+eGPnlNr+J7UeCYtCyusmf/4lfyMuaIh8PTyx2
laoMmXLqZ6qIZhIG5nERA52gNtTb4Nn2HygWmW8pQ5x8QRBqgz4DOxAyz++W5KiW
SfUzwWMdCceabSUO/XmDBrnolcPzYsXo49rmmoo3Z6bBFF9Df/Ktjj3uy7MQWscg
kxuEwUEcf8iDIBhHktW0EWmCO2toptFlo4vzE+Ndl8sl0NOhS9XIwCaZsC9yWMLH
Sk1dWFh7g0V8kCF9BUwki6K0J8bUnGuwOcPMZTwHDD33n8fntQbSCW1Uyz62gLvO
e2PWApuZ4NnpAmaehufb4E/6PrBn7MnKCjt91PLfGfJMPJvrgy+eOQo/0mx9WEYK
PVOgR9zsyMGkYnav1KiQhm0mQ1xjV7R+1F/PhxB8AUmG2QfOybQW5PK1KP8e+X6U
B37iLBTY5qYR293DWNxGNnMzOidweH10w4IrymT3s2S3re0W/09Fkw2aZnFfOhqD
Y4AIJxgIGzYF9iEDV9RO+Tam35YfhJFhj2JVMVP+TCUWVeQOIvJ/T47Q3lFaxaSf
6rbv6D9zdGyu1GO8lyaAw3r+FqfdVZueDERD4KiCAFtEtTeqZHp/nbgkAoEIV5n1
BB1+OnaY+99QJNefXLpX+0Lz9yK3fiTQbOqTcPOsmnG7qS/3YdBqlWPqK3Xjjnfy
OupTZ467gwCmXlM6I7EH6Px7AFW1hTzd/CihWgQWvAErV0/M47b0KBbw2gglhLP+
Xs+brefEy237ol3MWp/F0QYbpemchYdIw6FMynfrOGOaQpnwHx3XLOzE1O+eTqR5
Y7bEiQZieGr5i5HYHcalr0++7DBdFV2X/8z98JHEl2m1rfBxytdfonQ07+TKo16C
0XYLfJvxHMvB9lr7dujKfwioV33iOcgX7uwWzkbp6fkzFiG7aZfLh04q3UZUzHO5
A0YAArDn9A1NhuHygQsUw8EvzOe13Ycpt7xjPbs2cvUtsPC6iN9gZyhcLupjOHvf
31UVbnSeZDdfcQEwTEm7YVHoi+qh87LZg2m+KRoCQCKoCD6EHnz7XtMyNcXEaq9k
XanRRZ4RHeGH1RVtjSejNqToZQaOHMQFluIxfQz6n5YfOKp2pTni3gRk1zd2GSKS
d0wsibBBJtBP8hLbBdmv9g0s9wyrfDX0xmKXpYtUnp8qs5XMM7Cyv+esYHRau9Xz
AiLQ+Ai69yzBNP7Q7wKek02dzokGz3oBAhK+8UN9N2b0XnyPuVQS6+M97oL8lo5g
5Xa02QHPKrV0zklv9r5atkDG5GX8c8/PoOoYzUpTp56R6oL030qNk/VhcikAJC4q
w03i7B3BkCx4NyhGfWl/JpFfnQSPjN/kC1xx02mpLQ4irOBND3/lZX83v+i6knIc
6mMvz3ZExpxaNsMaTSQYZmdjUmZFEV+1zEwvrr7RHa28yMvtQqmhT5hOijLdLbl1
///QZjUKII5996nYBPnR9P0WomL1YsVBCKwJ2gQHPxnLHdFqK1iMxRt+M1yq1vgG
9NyLkJZgP5RvBLZE1a4qXxSzOxKgJOMHA3TCRKU9mg8CPOggu6io9IkzcUlMKrYB
9rBEmb8SuRxuN7n5JVT1WD2T2Ktw/q3Lm1m/fnCfA3DvIZg2uC9ULg2H/cwY5xKQ
0W1y4loyOKAOWs1xV+rg6uzIFnlGjv/l2sTcoJiu1dt3kziK1tOzYLRvgMhL+kyq
yZ+l3k3pVkqS1WjnoPiciMPJyeMoKlyax4D+I3hOd9Pa53KhRv79Tc7G/REHbV3E
6Mpz452JMErlXZIPOsHc8FBS6dw3xwc420xoVax+XzBXhkHL0JNhhd48QltR8E0M
D3LWcvxPKj+CIQUbZK9VUAurwFWCFb5UY4EKLxP8wNuBiDjATt43YN2kZQlPDLdE
bi6cEksK7lrhttj+JTQfwag3T2IU9xVnK9BHNBSEDHFrg9ZFkCklgjKI/DV6rlQK
8VIIIdfKAYI74i4iebfYVUjUuX59x06uacqHKoxWkS0A1Q9zME7wsZMFc/Hp5y37
vs62qyFULTyAra+PYcNcfsBRQaEc4aOt0MMg0deSi0cHiz/I1J6MgWPZwvAhQ+kx
A6qj/CAZt7cJDcNf+9EGq/a0JdFQQj4isukQxXdPkxGzwtt2LlhwQ9sR0WUNIrHI
HtnLBwtmM7HECQXqfZTnC52ZSCtZTsEduuOwWBTo4fCFwEs6Z1sDpg+rTDBDqmvx
FY3fZMjYqP8O1ubWoaDUHIePofUSFN1IGHlpGtYdss9KRrftdwxjewo41WxNy6dq
CEBK9tr5lO8FbmHnLK1ULZBPJJiriVsFXU5Q5t31pnDWRPb190rW5TtTq+LAif5X
3isXC+3kDbZI+CmjDK+LeUkU3ex6H++N3wnPs7cUS+kUzDK2f10PAH5AMQLE1SZB
QcKh9wcU4BcjPQqJwdVSugYG7cCE1UxZpH3B538zXD5oc0EFrklwZsoBfek40hos
R2w3NZmUhSc6IFjhyjX6bw6Y/mw+dlohpAM/jfyFLfvyltIwnh5OE4mJq0/LSwmw
JA1M3D71fmp5UtrKLmtubZzUoWTTrxKvyektn/e4W4e1iNiBtxxqgRC3TiD6qLuH
K27iWtQJR8CX9K0+UCQaJZX50RZkn0zERfvzbaSIuX31k2Z+8BFzCHvf+B6zVBkh
MLV9B3SnytLWvqgXJ7WHMv0jglUnvj50oFby0gfK8aL+d0N1kCOXryXFNXeoxrRR
w8aR02H5BE3anhfUrYQonkgm1mB7/nbKV09HnyraNEuUGpkNShniVeGurbXHWGdl
mDJUKVTGIv5LiwoO8eodniwmc1u2gF0Dsf80eXzUk7iY54M+nmMrQIqdhcbryqcy
xnLg0JPDwySlK0MDDEBCtCfkXoEy6+96p9dyb9LTkmNYltchoFAPej6en7nK337A
xjG8JhW04b7I2GvA5YwHN6OGlHTHTCVwavApPHkXfP5cr767N0Vd4wWvzXpA+CRq
IxG1FUBG8Su5vlpsl7poHBS1OoAwBmJTbUJAeRMzwDkb1SPadsuy1iIRfRgEmjvR
8ohF3/IWGwOGcvM0HwNmkw1L3JDq0n8nYJzusg6wSr+T2q+n9ASyPXyJQ+2q56lr
prhM9+tZ2/YBZ4jTH+VXVKvK/2+YrXjSeDSCi/3cfpTU+HQllH6tFhs6czgwbk7U
Jcb9rjB/6eOAhPxe8LkiUdBwc1Awn5vzcTVn2YdiUZcqzvVO7NuPv+8JGU2a9yr0
eVk42Vy3BGvsxoiPfCFrl8BnDj3eHxQL5+SzkkIbpYg0xYNxGuADbjRDDKgR+98e
Y4z2KaLSXA122C5UlBKASKS2DV2Z9lHTtPLyBo3RaGCUNMAOzSmEJ+qAMB2p94rd
M9cX37x0YKbVB+mWTnc4A/I2focB7ciMs+7Imb5FCB6n6RjdAhe9gUZ00c+kMLw5
WESRzl3rmxgXXUwNIhVUzngaTZZrlAEuw6luLaeuoPDBxuzuJs11uOk5xtpsIjwa
DurF1GgR6zOpiA1W+apgCLeOj80ntU/064Q2V9RU8o4uO5BA7zcQz6VWS5H9/Qeh
4o0Ecb37aAXv275eBS9f7XvzMF5ftIEluuoZHMEPt5XOkANnuuuY0KPqOjDRBeZ8
lptVk17CgSjE3NRHbjQlC47hmfESBApX0KlTiTDXc8ri5qar55S0GNR/xp0dDx3k
gkQ6QmNc9I5NKTSOUwTDpKCb+qdfu4dbTXWu2nW0qJ8vMAE44eSSKjsJXinZT2GO
wsakggbDiXK0z/Vaac0yCChRRFyIQJpB/beziE6Z9sMhvI46oJlIgU0NRudk2Ikj
00sFEGLnuYPA9IJitxSNsLxrlCuxgbV/nWQLfT575hjvNE+DH3BfEK+ZidRBQLNS
+7mrkkawPBi/iacg+vimEP5unzc7lSAUCEOcAwiTEy/ZZRQjzrbddoe8bdXvn+DN
YWJqhQdfVY+IshIlmmemWWuupRzxK6GAMIxebbiomIhWBFBs4X+1MsfzvofuyAdD
/06dkgTqpAbrGRYZPNsJEW/SsIGhoRiOvsV496MY5GtkMcbR56FpzVyGJP4n0JWc
apiU0AgBymdCj6QOZfRiaZQl+OXW9b8InSr2FBDmK8C/ZF0Xll+mPowLlvvvf3WX
IAGX0d0ccZNonodxgMiZn9TGV9SQB+sIyqqgfxG8yw78cVs4MMI1XLSFLTLw2b9S
CkretQ6nbv/36D4VzekCQzbQK6SbpvNpSGLKp8N9x651aJC4WfZZHxAY9NYgRPkx
eMDQGip2581XyyFbSk+/ci1YXpsHM4llGhSXLL77lDAWqC1P46UHWJB9vKDSqtCj
W3G7ObA1zyZnlPJ2oGjxob+QdzqJwJQcCpNea2nScbandXjJGeRxk7gX+I6vqzh6
YeQO+YiTN9nDR1eek880tMDqZEvpBOv+cVE4ZR/rykl3g6UcWkmBEA8jqQE8aG4i
Y9Luq2J+C4uMIc12Encsz1d01/pPWUIMIYPvY/MHntdbWS4MLlLuAAy6T4sIyXAy
MSVYoAQEmWYRs18iSiTyI9gz6SPMHEBKKFYbCLDQzDBxou2tzED0TkjkiWDb0MPb
SkE/r4E4rYiMfU84eNSHXQvljUN/sALNdRtuUf0aCs7ZsgkylI8I6BrDbIYu/zq1
RMa1NxaMHzdGDMGJ8fM0Fx+Mz13DeeOpeU7ustmx70yAvEalK+OPLWXL7JBcTnY2
DPHWpxy87+weNttDZ0HxePSUxyjYlFG/o9fKMk0m2KeuFmaTyxbxZb/7IsDgYuzw
57p46meQSofg+ikRGx2Mtw4MwJdZlpJ6E7Yy4qH9y5OmkhQ/69X4sox38Ci1ADlo
gZ1zUYY5X3033jZXexmG7+3bXlgY38onXo9IqquwFn+DV9o6cpIJy9egCRF782hQ
yqqeHOppNemFlJPGUiSb0eID7iwnS7gAIDVqIm8dePsWnbT7qcfH/zM0J/afj7pk
JYL9G9DqmAauqlK/kzPqeR1+l4IELEORy7djP0L/yYwv4dPm6R57+NmIkPgS1y4d
VOUekgIgh1/ZmeQ6RO5S0ih0p5e5WQnjSxHGjuBTM8vXB89cq5RYrOQWBRvbGPtY
QS34efrbD5S/nzAPhA9N0+RE1LFzYiwTI5TR2Cj4YIJMM9BV7mECafmEH/BKCYxG
UiiQswSKym+BVkvhjXSremTUbCa0j83rLo+Px7JMNt5bGAEIacNRWsZVSZPqXE9m
rapZ2KDX++l4rekyNoCvLh1IyvTps7TKm9OMUs40sWy8/qKMwwQQCP8YjCWDHaXt
5EngM+yW2ix1/hmNz1EaCKO/9wFmsR9omy08t+XPRophJdq3na+w8wrd+BvljYrI
0KkN+3uMM8HkRPxrwzd47CxPlRQuo6s1vdIt3Y6ffLwDiHV5fz+yS+gB9m+394VT
PTAPXEZ/GERApwoLuvTOUg9/0GO7+K31LOVyRhqpVeQ9WvTOrSA3wH1dJKX4mqPN
V87mRTs9gB6CE6NpyrKB7S/MdR2njbR+eqqP8PD2qlRYyo8UHqvV4w3MqMA0vbum
UKrKD94+Wkap5eQux09AYE7bcfJKZ4Xrc/Lh+L62ehDr4MBzyEQbVgxdNVCvuM4U
o3Ta6RqYqsrlxyD77sv4U2oqFA/o+UGalWfEratZJzcxRdTj5VZ0huv8k2JP4Cik
RRIx+VK2W2ykDvRJFCpe/bWE22WGJEDUHXKPLtBoB7IQXewDE2xDpl9/8670nDad
kG5c++HK0ssQsAFObttv3TNDasbIqkpq6yzGYfI+goZ8kKB6OBCOIFfjiOiyAGmV
ZFB5EHNrvZPrdalHaNDO7MzOuU+H3W3I3twVTg/FRBeXQ6dralWE+mYP4xFwIr4c
V3B7dro7sBK6BmBz9Bcy+i1DbpM3cpWDvL73XWxPsRqVdrEkpXuYs+OPvIQQeKLS
9nWs+oyMdcTJ/Xy9ZUAciGgqh6/h9Z1Z/PSRGYZ3LDVifWfWNqJJRwVLmEGnT+sd
6RJsZCfVHMmDC8xuRaXQkee5euBqyZyThKOAtZZZFGqPoRZzNjgLc6Q+MzOnWXAq
WSx8wgBHocVf5JSnAIBNyRKMGEJtGWHwcgqki/HwJ7cXcZaxlGtQtxMujnv/rv+r
vrzv1V2144vNIMX12Cjr8nmNIhVN/GQY9aLICSnx/W65hMduMKNUNrAhVcqKPstk
YAJ0i/6fsKMe3kmAIVMEpzLVxCdpg930gVjyKwgs+G3taq1H9x/EdMQxQGBisz6K
Ci1xo2whEOsuUznswf7O4sUtk4cFbj+3HZtuNehyvxh+K48Ed8dhC4shmRHjgijv
GBmPnbdt0E4L+k1FP56oGSOcl2zODph/6AXFQWE/qknr50BXoOsop7Dq5zXT1/TK
MR6J93qYxNdgF5zke1OJ0qmmC/jhoBAX4sTCzCGl1WO+eArI4PR3kRtC+nBKqdlC
BEfNRC6xL16x63+SpWsquI75vqtrL6SMio/Vtgj8Ym8OPWDNS6GU9E1DvGb8tpgV
2p80M1StttRcNoPe69fFEgdxd0vPYfPv7DkhmkJRRkWyDMiU0x8OEEYdN0PuVPz7
LQxzv/INX+iVIokms5LQK3JqsEDhOLLJIMUaDVeMn0OgS5j+IqwOPTeDhwams+zV
HqIlL4WI9DuxgW2ZhSAQbh6fVDLaj7QjjUCsnPpZI6/WS2D9s4JdWJ+/oAeRnmde
dR7AeV58DAksSSUaDH9Qq2rqnqf278l25ZJN+D0q26sTpHRXUQLyW9xv4ig18tKZ
SpLfw1UwAFtk80D9vtWT/JcfHGXkt0AdRdxXBkNOM7XyEQQnrDbjGQTW170wN8oD
lvI9N9a9JT4I8CVESkpUqyNFdbcHYfcn+p1kYbGzr4PPlaDC4oMA5+2nnzrdaYjO
FZ/8Ivs6qX4UhBlgpRS3DzVzT+BUmPi4fgP0FqV3wxH/cEzv3gwILN+fmXZOLYT7
jJ0pCOZli2kRC0pBBIoApU9OMFuoD8GQkhUii96PZVbrJ74v6rVOlVJ5NNH0UyYM
8SUzq/E4gUSJMpAIbvyIx1DH3b4TUJKGsDHdtgPhImspDjey21k1+ClWkP5N0qOS
Cmfr/8qZmX/FYY1nTMKlv0PfWFe/Tn6B7ScEcsjG/6ByeRXl/hRR/7zRgxa1qZKS
Z6JXdMJzlEs+PtuwANccNQSfp/TvrofVwz104GQafxpfUtZs59R5bTsrdUXLpI5g
DUuOiOWKmT64yd6sUl6KrfneSkxzA9pfatf9U9onAUoUf4ssbcuIIE2LXyVFiGN0
uo0Cioq4BdErLhXdhz0QOF0WoIZpHXdQOBkdXmsjyPW8xjbVJEgXp/uFEBgh4ZzV
7wVgY08ljBVurL5GAPhHJi6OaRIzjHZ7BMob8Iekh1smbneBvngESr9fKp8azYFC
CCn/76EnjsQGl8oUTetm+wgMV7QHf5fAYFJJ0ZpgECJBW9kI1CElgh6xMOSBKb7v
d8dsL7Q9bE+31WjmkDBfjth76+ZkNNDByfP9bDwfI9CLkVBlr2M7IckayBF/Ltio
Tdg8s0EyufKFNe4QKDOs64OVJvImdxole8LqgIFrmX0YRzE1N/qemjzo1RmfpsPA
iikeTDr0VDW3kD0KKOCCs40+XC4JMSC9s1kXmMhZ6T5fkIRRrNOthgs+uObgzBay
LJuEyQJ/p4iNGYkQYubOJHpbfMQ3tMQH8HNjZkqqjdsRX0BvinWY4I51GOI0bmhb
OarAgoG/QsiJRVmm11LzIOauw1ZM2utQgsMzfSvkxgG+sNJPGglNynCeviB/EVfO
UmPo8OP6pRqIRL/rbKxk+h4zNKZrOVdZ1SedkDsqAD/d7WFGQWKzWm0Wm46EZP9H
FkTM4mQv2JiK17cuDOC/O+w3a5dgdYfE4Yy9x7gjhC1UkgUAnpw8tZy83NrHH3/C
yp2pENMIseyMXobUh0HGDD88yk4WKVCmjzp2wDAXxkuq3sL1vQhTmRY3zx39i3w2
30tpSUJk+J53+fSn7ja322c84KOEpzVFz6vITXPEQ+Rhv8ed5AxFlF2ijM8TzmR1
1IkhHaUCdDrw7Si98dRblYJgn8VLuYgVvJJ0j7ngCKPBvE9cFIR7KEwA0jCButSF
Quoos+RitF9p+PHTlYRBLJXq837i84W74AyZ53fN1k93dqk1dvr7AhVzXkzNrc2U
xkQ1gSv4vZLwqle3PksuuXgtun4yAwKBB5PJGAQTFAX2pjktwFHqVRWhPuQKugXY
MViSLplngAEFajIvr5uS234xafeX+vt7RJZqOpmt5GRiXgRj06DdUUrDP08w3ejc
tHW3MjAhACjqWrQZI9Z+r3Ii+O6/vomY0pMQPKeojUCLUl4vYTgJRvEJCCzhVNJm
0dkEw8wWVDh2SS6Nq3un4WD7+hVNTbQSnwmTuWxqWwpE4dKNyDW5nd+QyXGRo1SS
T8grQ/Rpas6cR0LCthOl8m7I9UFXfAIC9p9vxUihTYdFJkc6rHWj7FhRsR5acZdK
nr2ADh+IDoXt58JrLQPkz6/1+OLOs2CtIpIeG4jqg75aHoZRgFMapMdvCaOnbCle
lp81mf/weezTl/AmZVKMq6Vh/t35lnzN+BmIn728d6i46pDQUHcf4i7ANzxeBHJi
X9QY6lOC3kTEfPcZPyYADq+OJDCy1N9+oqZQ+nDFyWTZHPOO92RNmAlFZZAH1GFK
t1qewi9r23unFGD3lZReMFkpj40HcgtAjI74yc2JFSHhzUHSDbEqyCiNKNm562/s
hUJxq7LVfjkvGwbnADlsCQsnXtYRbKI3oeRw7jNhBPrvBlEdNY6DIYN2I1QNCqEm
aCSJistNHg4IrBqA2f/05m6121YSbQXrTozJ9aAfpXoOzs3Dc0EL+iE5oHXpUsO3
gzKINdQ96Q7kZMht4oVVznpJqJkmjJ9n2mXL4SbHF5egXLNmC7ub4NNKHvNXtbhg
6KqJO1Xs7xQstrqpt5traZwq45ewVYNPHxKotDqOImHKu98897TBqdqMznN5FXpa
OYsd9uKLpXaiTDhe4A6z2vGy3NNZePAX//el9nEUnHnkOO2JC8U7qPsnivPH9l+o
8AgJVJzryp95N9lkwkjvcDkTNqC8qoe/Dos7ofIcIV9tkhz3W15510NVwaarSFLd
eMttLJz4duS5hi+UTy3PBh/hicAR5twcH3k/Y9pklHL4PX4Wiq/o6OvilIa1bXxs
N4Sp7Vkk34cHulXP64o7ucnS+SCJvRbv0K34uEKqUWUnrfJOCvgfnyItWTBmBTCE
Ac8gQMUTV836/+qkuP8Jb3vY1imkDwAu/afPgGY+MEw1YC0DjlybBuEf/aaRADgR
2VXzmNQDnUxVRQEcmyutJhjeqrOuq30ya/Rf/7bvZF/2XnFFLfW4hTeTMDDf+CFG
idD9KX9TEqyBmExpq9SihOSRXL8r0/EcFgvKeJflNrjHUPa9TxCsJQS4apyUGIRH
swlnks+I+nCv3ncJuEiL1oHbAezm27+6iuq8WOthkjZV+8YV7uumVjochLIT9iT/
EvWrCI4TzTF/ImggJx30AMQbb2IzN6L9PfozEpgCi64J8cl7rhRLq4GxNQn56MB+
TU0MM7z8DGdqYyYqQJEAOTqOF18oyUd064sSl2NXPfCmAz37Tp57w4oqnKsXXu3E
2t5uzW7Nk8gLAEcmkzUKBf1UEcML6ypoHWCEnKSAfcUB1GutPmtGxkFUx4N6cs/W
j3DupHpHZ+wkcOcFnoSjYRn33Y61HxiqiW/aZQTcb3aHViJyl5X2Ej6EpRD21DEb
GJ1xyQhELXpQT8X/Evl0A+zC+nKkwy9g5gFKB+LCi8XhrSSpgtO2wsAkNVt3wRsM
VB9tpKYsFYQKamhz2SZG+UZJrq46129Ert/sSrTOrXyOJukNSJfqoD/Vd3Lt5IQT
q7ByQa+sbDJFfOpvZo8exEwdQQKi3RUUa4frBP9f1lzMqZJipJIAsLKRWn6Fep/E
fG/bzJyRBeLM7MSvB+gsE2IL2H1HagGXfAwDm5kKuukd+l4qMlKrKIHSC3CH4rkY
+be9Nyz2sekFnL/WKEIMMDnxAl6p4F9P41gzwfpOAs00tTYCKQpgyTAvs6WA9sFz
/6u9dy3AvE9fsPf/aZUk9fDzM6ZjVgxHOAdi/DOW5LQkDWY6gI4tl0MjayP8ffF2
hMmUwMAAOfaIUhIyE1Fq/g8JbpCH6eNdxqnaJjuTMAi9SvuR9+S+2MS9OSpJHDWm
KoJstPRAyREcaIy3xUIobLA5bax+70PoQnKZJ4OVrm9/UYZu658xrzMW0z1orEzU
YIgZjQVod0H90tgjnXSlHKv8YXnxEWyk+/ukCTEDsJzuirkDwZrHtIiwIQf/v4yJ
IG36scAeIOgfTnguzNWWN28NxG4cjayDcC6zuKwNVsqpYoIAeCR74UpbMBgV86Cs
aF1M81yGZeiltm4C5J7eEk+JffiElUxS4+7Ny3NHc1qOSEOruwmsDh5NwBnPBWBz
ak7+nDHycCEeMcaj3WnUHU1UReDNvCCkt/nAeC3KwY81XxQTQl5MhXqS//lfu78u
FsroGCbaOMGDu2TY61Ilp1tIgah6lOXHZYYv5Ba6bl9XwpuCPbOhPvRhXYXG4WBN
OQOmNhZpEJaUp6khc17JUTi7EumYpkghIqR7z34NwHSBN/jwEvfL0LgT0XCFr/qX
5SYxQM1f9gD5Cila8EmjtJTKefz4gWS4ZMBp5+3SAwMnJ6RMg6quv+fDnvQE5nRZ
aCmwuAWs1XlXRo2SF4MlzI6OBx+v1vTiQX2l/63hlengojiB1aNd6s6hS0II1hkg
woVmBc3ruKkwcTT7GrTcOX4Potavq8zDtr6wDLJUaNzDhyBXvC//h0bLktW/XeB3
iKKzrt87x9q2jV+lY7+bDwtg0uvRq/fFQTBHnMrMVT//SrBLc5di9HSY3eYGh9wA
jLKMSSThLrhGF35lszaq1Hq0t/UFVMOdfa/7p/Syo1F+CA7pUg25nT36bxRtFZig
xkM4MDgGA7W/P36aANFO0i0Gw0ra/e2YB3ZceYqexHzlSv/B3ZJvpd5KQ6MPRdHz
agh/Gi1tjWh2yFTnaUhbKwbIsaPUb2F4wOnHT0f9QLB52miM87BOu3VnpPyunzL1
3kiNas8sDjE5xQMrrJHD1sgApev6JcpXu96VfW25lq/SQj4WX+d61TF20COQEd44
i0DWCrG2XT4ebvPOUjQfeTo1NHoOwE3yfXBlQjvabwUKsL8jaf0m3nsu0rVC1EtV
rU9EFL6iddyJzYtlHMQI/Lo4mDCQ0dMSWJyFH2X7kD4yck4fZJllPNO+wQJwLj2D
BPPZY5br7DTRfFgdE4bDkW17adtNwv0s5zrNhS6Hx0qTHWDTNKTpYCNMYMIY5oZ2
MTfjtfjCeH7ZeDVuNxFV8VQH6UpcoDmbxT1e2SRcEBLNcXj1CnOVn5/zPFJ6Zbf9
TyxWV87eCUVh5vALEZHNN5LsvP/XjUKxq85euWKXLz/FwAGlNPPoBHxBnRmZRygJ
m3O6zYVe9STj7b8W0hvCV1Pqwk8tARLfQEVXzi+jlre5eScXhzxt7WLH9iNRNMwp
GSkrzcxP+roiYDfm1aPQjFXGpSdhZKTJCDkLwkkVORwybtxDfnos/9FGnp6GV6MO
sdIPHhGx0qv5ddyH3+HVRBbvTA1sUo5X1L9YXe5IJg1r14gtWnNB5YePAgNiDcmo
bQyklKguqDWvLre+ENBvTMkVzXHuNDBLwf+DD9J/h9j3BvgfTxiNWLPFWUFdH6Ji
4ufAdEfZGX/I9/SnvIAQzJXVYMpqa/5Rbo/cqrmciarkgpNtyfBRCL6lO61emyqS
AmlCbXA+T77VVAzuOIlwP3EhmUPFzey1Cp6/hozVhuaWGq2zfcMNCgFuKIwTdoVU
Lg6cyS7Mli34DMjw6haAKF1b9fCF09CYTZPWRfXlBkJtRJL5Tw5C1FC1tkDGecDe
vd/FHXulIkeGng1BWgw2uyv/cCV6dKTb/Hq5tw8gW7f5V7MzgDCWdce3RByQzBSo
aZ9EHK8g4Uhl/IrI60/FQ0JD6X3QGrDeiwNDl2JFha7GBPL8Dp5U/usqgRS+mHdf
ao9zLqIPEXema9z9lZcAitLuHwEUEsoRsSJ2O6dv9h80GSPMv6OenW+4jXtIZ2x7
SY7iBtiZNJ1LFn+cpKbmqY43lqxGMMwkmZO3F7GXPPHEeCOBkKgXa1QTLXve6r7N
hlq4JMytE9WYD9/mk9umWJjue0g43buYxQD18Ro3SgaK1Fy5dSMtBnAG1AW4sOFw
+QGLCcQCv1Nz8J5gbIvqF8Qf2voSoja2/SbNb9Dup+GCkBy5rEhpZyee1fVbqnuE
gH/7B6osNoiHpR7jBwgK92y7mTfH74NEDqI4eWHePazICOOLKZLzahaZrWPEtedd
N+qiyGMhmdvp6wNmAYIC5Qz4eZoovyN/J7+e2M82IjQW8RoySsOoYeGWzowDZvw2
SHHzVYjktibzkyabBp2Gj6p2Ps3vTGsWsp/zMrRRzWPIk33rtJBktD+zM1/U8RLa
b6o01yF56MzzBlMu09kam1Dh4QvQKDaYfLWyAwDS+SRHI/Q8YQplH+pr6zoD5rOe
yHbxrik96Ne/1r84w86COpab2X5ojmVfA9xCP/+M76klWaW4KwQPB4B1ylxYuHwZ
G889KPQz54x8lcyB0P36rZUdz1WOpRAA57OM+k/ULkZ1t/bSYFLX7R3ZaIximNaF
0M+27DWGiCrpYpHDPfgGLjDy1QL+Tg9NFKkmxk7wmn7sZHR5oAkwYTKgN8L/MLO2
DAqXoTQM4V7jNO50a0sga5RIbrMMvxdjjeeF7m5or0eSLTjVN+8Soz0EoGRuEIaH
sHn0UibkZt8Ch060LF8K73fD0B6s8WDdPXHxY8kow0j5VR3MZjZ1Ghp/LG8CbaLe
kDy2eqpNkONJnbeem9Se1BJ4Z9lP3uQefXszSf0cTyT0pAN5+baN6/ypax1DQqu+
+PuwveNu1UekgQcJ1xQs2VKYsxRyO3fk2UbTKlFFlRz5aXdO2+mEn92OvgLX0psj
I0eUPNqsEekpz+InkSo+oQ+uDRsdHb2HsphwsAZBVRNAxu0cAYJdgcyRnj54kivc
4yVTEtxJyRSs9o6mUWzdQzbEtaqhKp8gtcPurNARsX56GUlZcKuttsKNglHzFd3t
SYlUbOl0qCN+Lvke7bdpAo08AhkQqwOgUzMF8Fba9/0FM9mL3d5EaBm6+7unBKr6
XDySeicS0nb9gdRmzMnxIWu//FbgWXyXLHX0/BhJ7c7EU+BP0BhFpAo4Xy9QNDUY
l+UqmTB1/aVo0BO2B2QPxiTrUkePSLRwziZgnbrhC409b03BY8p3lXrSIb7VmsLy
UiBmeqwMOXejWVXrI4S95Ubb/bYrle7UCJXdSP/E1eWSWqgfjZ8MNdpw2MDmL2HO
8ldGhjDVzjyRCVXM+iRBzCw6LUShV3gmu2B/xXT00A9ZRzavdCbTBOQBUgLraRD5
Y56V0mSy2PnJDHGftDhYF/DImkQAj7LOFBaois3lIIHes1pHy0NRQ5ngHCjpk305
3ocBeJeTlfK9SDkkcZUzn002H072QLaicmBLCKdPTPjua/ULWDqr3yXYKu4SgyLD
r9W/K0LisM6ATz5hO7HbtpKtLrgIODCoRETVTraI6BVtwfERpH5WjCfGpwf5gKTU
JZOOIDSirNApinv+Iu8Qc2WmmgGYUSDVcluA3GXd55ogh4Jndh2meTvD9h4MTuQd
1KUFz+Kaj5oANC9uqFPKdKSIarLetrnxdzZgYmD1RNeoHhG6l9FWnaNwsdKGg2LE
AIevSriUpzfMf3cpSa9acrgFXTUn/AbDiZPaDlPIlE7KO2886cXtymUntLRuv+tK
0RxY0dARFHsS/cbxDQyrxcuMB2AMWXI/nOgc7X6caU9Od3nH5TUcU8RE8wkwPj7K
IpfhuSg+IHLjADL4WyXQiYi+n0MikHitvESN8bERV0lIxrvfpYwsbovn40j7F+EZ
euV/biyauaXWrcG+Dg0Gihosz6VU9iSKGcAVx6K0PIB3YxrZ6ydFcD1YwtDtYx9A
gLnwq4a/kqHZb7/ZPIFyEELedvO06j2iCwI+ilpPLEhNcH9prucG25jz1wz032R5
hpL2snbDY+9hdniMYPKqVnte9ZeZrdNiXsBNF02M4j0tnrs31HAmHBfwFv/2otnY
797UV3ZR0BajRj0fHw9VyChHhux9XbjSG/WF31TDUm+mJbqFL4Vt6YbWq5qbOWwF
sAsdCfhfjJhngMlX9doK1NC97zmcYHst1Yxcl+5dkvZJg2HoZNOTS7U8LaeLWyY9
UY0ZeXWNne3pvjstQiadGElpY3rMP5etogt4N/VUgnIgdbDOPk71U+H/y28bL7p3
AmzcBMiZSRCMnK72a8oM8HBXO1h3ZSjeg9EqW8zvDL8x70Hp30Z2tvY1CDk/Tz2p
QHqaxGqenJ9JitFEOWCwGGAiABtmKtYydyZb1gcJiMKQN9ONOeYUDWnScGifcjMo
2m6oOjx78EqI+ajmlzG2jteW8wuuzhVXmGfL8xjvsbY3wpDS7yF7C2B1ObC2rjwC
sbpxjwtzPlceGQTNY5AT2lB0LUwJdJLafUptP7sJ6HohZmbFpjVJuque+IGsDa90
6yKlT27TLxWfNSvr/iTg6QLzP74h2A9Jt7oU2A2Pp45wo0EfvBGpL9N1xvLUg1iu
bFAiy4x/MYYAhEsAaD/Ys7bCTqcgmaZ/cm88iH6KObN2UCny6rgdxD/4N32foGJX
NUopJXBa3izm2uscbSZSoCFI/fct8zfJpQe+SvdYQ/d+KluLUFAxk9xmtqCq7qNl
yySPSxx8g8dmyzI2oHTLQ5NAxC++OpMQMtMZbS1cgzpdoZJIXtNxvSZIe+ZcWEvh
njZQxNqH1lT4MxXnYM2nvC1Y/TE72V5YmnBcZRx4pXb2R+iZohxrRgmK/UlR1iIG
t5HPwY/3lXD6EFALqtWlzfNUpscSLPN2QoY/vSI30PhF7RISrZUscCo5HPHBUrjz
Vi/3E4rt0CNeoiA0m9wQ7TGOsrdiUg85xRJrA54WsYFXo8ERvUkMhxXht7r1lYIb
S0hveLZ3hMjfp5yp/Wbnf3XmofJB+6V+48VwfGvYjTnxnZsRW7OZWpUxzJ5Txmyu
FyXi4WUqDeS7IocKbB/s40K6iYAT+MckZ3VFyNF7eB/kmOTDUNVBfe0blgNtptvL
iyRSAU8MvQw9lN1HB2bbV7Ebdp6sKvSU6IOW8cXJAwktqXX36BPcii5nwI2ZMzb3
yYXEFO3udjlbyC2w2qR+G8iKTABipEmfKp31WpPd1/2595wRRJRJ9Ho+X/SqsPr9
42MNerI0k2VX8sEv04MbnvXNoE8ouV4uS+2maSZxlUaR0WBVUgjpCryW+lz+BTQQ
75TVqOtbg37ZQZgljZTXH8WO+5uRsm1nBIH1vQH5iKuo3qnOFmXkvUWHE9weu0X8
ONYy+RJqPozlMsmk+y4mS2nYSfugG5DNhdgRnJcKgimGqsnXPVV7qIOQNgaHUfWf
QmnP/K8Aqaklg7Pc2AudDUNUnSCkIk6A332RZxCdii8JSGI+vii7SGDL57E+Cu83
tLMurMKCAX1dnf78wd6uUIqUX2sUhMRGQ/ZOefakwx7nw8BkpDPqBdOUeakxFTLQ
K09+ao7fZdUed/6bQ+osIgg89E9JOouk6B5MZAJ3H6DC3PQE7mbjo8nn7RaAtSDX
NH2YQbSGIh2M45ONHOgnP5D1xIi35jtQ61EWw0HA4gCSRR+MHeZbTLBTfHBg81NY
WosS6mG8i/CjZ+ERR++ZtRBtW+ZtvLmR8rQJDmMJaALC5PvGA/GK1J8IzovPjop+
jNwtE9XaBg04bdcQpDStFt6y2Cb+WIdKtDYqe6+aTGGyGRCPZnYbBzZczOM0gLEm
3PJIrvgNnXOnQ7rrHFGS8XUEhHrditMmcJiWLFcY7Sq17c9xU6fgYIHIx215TPke
JR7T49KnTuKm4yOMqRo4DP6s6U09INWWp+GD/QS6nyodYW4y+wGL/dthh37mBYkZ
4igTay1GZBOJbFLKO1CS6yF8F3+r44KoPPiG+KqrZv+K+GffTypHEUpemNyOrH14
2kO/Ms25dHFH8N5YFRCEsffhXEucEQOncN067QkqlFGzwOGXXfC2nFZ5I7jdwtHI
18gZBKS8kuX7iqZhLmcOvlmAvElGqbTFvUEXLKzjgOT/LkCUcR6N8lk/KJ3opVed
dQtnrSCm3Tq97+CM06MSpBKZqM2+bvRa7lw8IdbamrC6NlxxCwzF6mCKHjI6a3f9
zo0vq8qOi6g6vy822Et6739c/4+tGU404dlp5o9vUoMabHUfV7XRUJk1lCdMir+9
TUuD5bgfiDi4WK27jt5KW1SnJllAiBxL5BkSA7KEvmbO0/ZMurXxJTBxcOEVx5an
ogEQvFHXu920intHUIenwduXs2PdELfx39xdS+IJp9kTFo0vQM3aDMAVWi5a3DqL
IGvFRcFb4qP3SmtYTXZRMSkBsSVFInDw5MUurPA9W37K6eZB/KnCIjtvg6OSRPK9
mKDstXwMR0XxJQb49KHmacFRraFwVCejEHTg2suFG4O/D8iREz/bvi1VqTrwGseG
GlZsBjT1DuJI0jr750yxnQ==
`protect END_PROTECTED
