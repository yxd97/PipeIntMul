`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hv2Qyg/jakuLxRF/9lkuKWlkGowZJ7+YSD9tpjZD+3Dw39pmANBT+QkyS7MDX3Yw
o9julUTxJ4oQzjcN98HXS8/p0A58UW88si0abR69Gn/tz3OjIXtw0NKpivPnlokC
Duvvn5weY31ejBrUh8jrD4ZTMaAfyrJmIVIzg7LOh5GleO1OuzPDx+MlSztUeeWB
pRv2m4gHYhx3781y63DB7MGWHGqhPY3fkEftLowC4PxxvdtbFh4U0CtI91iAawEk
+3YyxHDH2W6wewnlxx04fwVNgyy+HFB1YOJZdQJvuCsALf+zB4Fd4C2Wdwbr6FPx
BlTcbvSpzapJv4RDGG2ecTTbCCfvrILGJTqh0fKpKqI5Cx9HR9j2fw4WvAkfy9L5
`protect END_PROTECTED
