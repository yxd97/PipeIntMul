`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJZ3mvxG18cG6ELGy+Oi/pvDUsqkMV8AFdD92hgL9xtfeUnOD9TNf1b/JOx9HDGK
CrK+rt00qX1cckFB+Y6WObDkA/GS0YNGe1seNH54BExG2eeMZ1hYdkNrLhZhyT6W
EJHxY0BUJCFU1qbUQU7gTe8FWWH565yrpsbj9Xd6NHnYs+dibDpyex4PFrzXVFOi
VCNH/qLr4uyHfZ4QTF9JWkluF15dBuam99egSnNSdNKgfk6mcpVQMRO78TwF0Ibw
fzbxwV6hyM/OtqcO15PXD0LCL8cRZc2PTiavvw0t0pZA0g0EjyYLTMVD4AgvrVBO
5r5vrkrWB5wFpjB+aCNFrw==
`protect END_PROTECTED
