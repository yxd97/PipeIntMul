`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SRPXXmv0xBoSwN3n/pFmLPVGA/BP7n8JQRmsipHQTE+ZvlGxTAxdxyCXZRZzZ5JS
d9zgaaAHXXfZUYZI1NKXJ1N5Bhnq5GZtanaYFmUEdI7FuKEw54yxfAMiitJVpR/v
MqzXZS1y2hgllNXWDya0MfOZF+Ja4NB+TQeghhOhECspFP6rSsmmx9s6wIEzDvm8
LNQIEjQPXFMZ4ZArFRCYS4uDGw7wtMfwaNezaK37KObtyZSEgxOpLYL3D7r9e/DS
Fh/Jd4EyAzpJpBrmn2jCpEf/1aw4/GuQM8xtCOw5ObiQ0cor8xAGtBTZe73a4bOi
H5bVYA/W0OMctPEez2Cb5QPKjrWksbPwvGLvK1UgMQdrEw/PUsk775oMZ877k5mm
vkzo++G4WldmPEBMRnXblm1lFFrgP+guYBsWAswHneSLD8TsCUKirXNMUxBIYCzB
QW1v2wW35ZFNMWI00/sYIDicvB8Q4QqjUlx3yLPF6+FgecoiKiY9+DKeFM6943vz
CJAs7MJT4jZ6x+o71itnqAhIt3fnNIrwYinzq89IpXZd1CksL+Aqr0vP00EVcQ74
MSsb6lM78/aY6gyjPnc5xCc0SxK6lDGiVHITjrwMrbLH2MrWee4/FcY5huySVOvX
DYP/itT9yfagIkwln6dZyD9rNCVkKBgfSyS7zIrdjo1oOY+wlvERQYBBWBnHKtdk
6Il64F8LpUhGkzB6w4xmOw==
`protect END_PROTECTED
