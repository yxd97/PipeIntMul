`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fncnfg6e0mJ5oea9mejWBtL06ZCEiW2MbL+EAiXhsr99CMyK2nq1ZLdus6memdH7
DRffVqfvSdOdvGpMQZhUnCC5yQFjSVr+iUpFj5IkZquyEaCwueWPXPxx1gXuGVnN
5C8wuwWL14UXxvK2k3kApuaGTD8eukrXS5Jlv21PisigvlMGSC7dr7qI/OwUzH8l
+/0VHF0aTgT0TQ3/2Ai9x/V7Vs1ZNmMRySD8cQgqWSB0GlBkWXr5cGnzaYPDvnTt
knCgP3MeLMsIhNpDayR8p7x02Q4z+/TH2KzjPA0cIh7HiO07NY52A/waYsEg8Km3
R9S9FNT2TSroQuvOTKg4UEhoPS4f5TCiIrpg4xEgPtYrh/KbFwtor5lwecvju1e/
zXRoGBl2T321GlNgSIw9a3WP5GM+dBvkz9zUZH6EwBHQuvR9NLYvISCG/7dy2orn
`protect END_PROTECTED
