`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wacIh7Iph1tYXP0/l6jmjuECpF4opt2dHAEunpeol5eLPp9Ks8SipU9ha4TSbkJL
K8EbkJMhZU8mWfU4cpeKAzJAClcro8+K5SFhTmw54Ax9sMlzGpk7Yst9a+FD9ys/
YWt71ZKZ3dgit+/FPfEeGONuBkrbYRAdUFacK8hQS8WPlZd8OiOSI38hEMEbfizi
ockq97SLcBzmDqdT5X0Z8iz2YFrYCn3V5MR65286DtA4hYbP+d5eEB4gvYWq1Pra
FFGeRvBFbHW6iU/sN+bXjNpZL15lL1SKVjaB6ASJmhaiIGkZQYd7BJp5+26SBTmS
BeyQfOzuiGfJnsdPTPpqbxT/yQqX1SUnyPlF/bvi8PsuYurB5bNnq6ot/XHuyQ2v
78/g5xxZivhPI+wLi7dtNfXZY+MVtcJf87vadxaDOTXQR62sPvTeAUPOW5SJhrtL
W2kC5ZuGLhSUtu8Fc0wrlvX0S+52fT1l/TumP6kIn+TNs9Y0PGDEhNncgDuxIH30
1j/3vZOEtXqEoUHXbzqrqdSdhVi29OL1ving8gHUSaUejCTvOf6IlHvj3QlJZYv/
YM5AzpCHgQnlepFvI02u/lx4SqFxNhARTD30XTHVWJ6SC5qDFBn0dSOlTPAb4ugZ
jDgLsWfDK74Q9/3DPhKdYFxvdtPuaQnpYS6xGpX9kAmtFBROU0vMO3CyAFNG02le
/CBk3ANhk1N5A1ZQN0VaWV5uX7V29Z3WWZIxxiqJvUNJW5g3VjI6fKZpzLoy4WJK
fAh43GfL9FXKA67qjzzdl1HssT5NokzsFDTqS/G4i4MOm+JGSSuJhhY5i02Bakdd
m7p8j47VgoE8FUvHChgKUUlJSEt1UM7b2WPXHueu8hc+L1xhGuEiF9qaH0mukovs
p0iFsJcj22AFfyVv+yMUweW0iyK09IrJyV6F2U86YYi8oOOqXEZm3lWLoH3UUUOc
LCGKpJKq50V2Q2ffGuC98n7/9AZUwYliyIsYzBl6Js4+9gb7WHFARgtm71kIjzrR
KikGTTLaHKIEOQlTX4k4/wOGETj2zybdKm4uclwuGxU/0qAelpOr1o38rP+cNxr9
ZTSrI5/X7Tiv3yzWeYdHplAjCY1RYBuh+GeBHNu4tsatHSUR1foXFkgavkgm+CoF
vFrxVaLYTG5A8P6AltCXDu6DlYeFAufP7WlOWr79gzY5n0eD0i1KzEDJlhcxYnou
XpojKz0NPhYS3bWpkS9PJ3X8w4EEMSLXSANbljwISvN7ZYsu4SK2rIEwyPeGfgve
TPNRWGix59xZwJFo86/m/wo3AR0KD4kBuOZrKYF9yEVsqiYKaDL6yorZOun8FUFZ
tJ/YvAZm+3GefBTTQf1PNbMV5/t/FyC13TjeoeZqnZ5SKDyZtT7Dzz/xYSOUhi4t
A8dKE52TLHqVTwmufLglWBLWCSjdb0U6idNKzKYo0rvbpKNwuHpA2zlmEgF9RthF
WS2n8g/RfPJG9rEmxnOUC3XVjKyGDuLwUq4Mc6htTtGwpArnAu5IxLEBfb29BLfv
U2Ecc+Ys1GBGl3zf4Re5MEBdW/s3h56Bq9am9K7Gs/rvdrWEp6uoC1O8oO7N+5yo
jfVKe2RpwlOZBYQVEKeudq8IAfZ+B6sFszBPNaTNusy5WURpnLOMIjYsy0XSiIXg
88fYAR0k2xwUu5pC/5U/EO9qDoiJy//p4CTIQ/1HtG7gEb5GYrvBQfWsFYl3zLF/
uTaiancG7CE67f3oFALtJ7+s0OuXQpDlgN1JG7qW7UIITo8W9XZwKNkNYen7AiRs
jk3KL7GglYNd9niF8lGfq8UUdz8peIv0Z2qzrETnXiqedRyvt5B1TpLOye2kl0sq
/pnCVtZXha/FG2FID5ksEBFOh2rwZlNt1zKRRiD86al6LDVdplEgbXsooKLPW0UQ
9na7c5rSzZstQzmbN+MI72cHMpTp0qLehkXVZUrr0QrqufmdN3zdJb51E+zgC2Bh
L5wTRfKg5yOLIuNRzQnI2sKwgL5QscsrkdrTRu6toyO3vQZuWpaVDOseAMX4Iolg
pUpKw28e9AHrniTwkq0eve72zZCtIlw2vw3cBDsvVsGuPdSn63Qvrt8EY894lBYS
n4ludJSyKLf+oDIvXcs1aowl8J5fblUIcBuiHmQNeOj6QeUmSz0Wz8uYYdH7HMZ5
R+qvsOffbNYjCNXcCqbmAmRc+DANfI9LqzPewd9X9tmrezen3Nx57O7ZfoscnJnN
0el/RZo+iGO654AU797aJ67OQi5pBxN72c0WnmlSBOu9FHXm6OxcumqdkoJSFhb2
BEXv0CGCAQ1eoVzcGubrj0H0vlX/23vreRaiVsIiAr7nk9kztgvbnCECdoKV+8hV
sIXY7fV03M9pIEXmc7IaiyfxCJeX2auyKtOc8goyY8IdyAUfR3mbI2gf4Mkmi6TL
G+Ck+/cFsgt2n9fbp9EEJbT4jLlgVk08wLqSgUOV+MBMRXOpu2s4adiAIH6hc7+5
bLP/Vjg2Pnkat5XhdhXsCQsiyqrJHZ/ipmFHp6BCGHpdgyDPInhxkHXF5YztZuHT
vQSjbLqnWh/GsCvB9qt6erz1GYmbeiD3oyfmj0rkyCUR9MRNmT+CzGJMAiTD92KG
Sqksr5b6gAJOSc9TyhlHj2Zstb3X5jae7RXWGRgkCKT4RTHutLi8OvlmpuzkiNRb
CvQPqb/NIm7uV1XpuICnXrQcuJNxst1HNuE52xZeKaROl/IoG3XJNJd2TgwGEMwA
CzlDcnLYHZIQluGPgkF3/ZDQrCP8oxm8OobxDqZQqhfOGoVSrH/1Cwv6MdDvKPmD
6dmjRK8i3bn55AHzBS83k2iIpKZbONON7wG7qOpnbUi9tnFlVsEVcK52kawxNngX
vTplEuwW0MWneN5hD6N8Ycy6MWzY9eP50SMJRRUl0cr03gPp2aC8ZzyYRz+5pCh+
7ax6ObxUdUxZqAYqTn6KXLewh2WztQpTsVIQeYasUcPyFxJVcQvwqVAlA78HrmRC
QW8lMkF/5RWkBLSC8Nfy/s7lWN4QasTCIlM7BzZfQ1Tci2fWnhkkr+3u7T/+SuMx
47h9Ut3DALWZ5jGJhmuw5q5WjV1BYZNpvziiqSMKZPcHtSWnWJjwKskt8Tku0Qb5
0Y/bFfnHAHZtvJqPi3mJ7a5sFW0YPUND9Zb88+XjKRz2kZRzBJitGF/NZyLXuAmf
1NRbb8edxGgSDk2sYAbNOiD6B5YK69Bn9ZuKYM7AnMIY+FcKD8sMve4dX4gXgH7q
5uoLYeFM7vNnvwHcugvIvpw9bJrKq442LMtpTYilrQJQ+xI9mXbF3Xy9srisK3ki
CQOuspiEblJwMJ6PKXeTKU32Pxf+xuW9nJz7dIvlWr3vFsHNLLbA66SQ7hqpxVp7
7JAjFt3uhDWqIpQnDPKVldCF9pdyPcq0T6j9cKUkCxpgU0OL6Okb6lthzFhDb78w
QxTiyk7vGoWFNzVulIMO3KUJZwAVCFAGCYFkWx7ChOH5oDyO/pG706/AmwKs2hU5
1IORCfDICKYQgQj9pF7mi/jHeuNg9KLLSLJUPUzTkgwWrhVlCCY2YoZ1aLNS6iIa
NJy2vcRGvmZXtBMyn834P1/T5Rg2AIvzGVsaVBqhPfhwHwI/yvBnW4e/8aynP3JK
vN0icnwIzFuZmfJqKA4S0olw60L6fiUvNOyX6wdP2hSQHnU4zF3H6q4W34x4F1UR
PlHMjRF8HDdusB4ga6YYpdOA1Di9EvcsoO4Y3QSDl0qlIJWRgmuCkIqsVSL2mBys
aK3f4+rZ+YFGOmLjSlxnJqPf8qL6LCZaoD3wZougpvRty8aU66JUnDCp56Y8vcZP
xylL2VMic8PK1S9I/jfH3RAoIBns+mgfq+KjB0FA9oi/taRLqG5pgiEZ+vBale0M
pA3ofa3+Sh6d5YvqwXD4VcxrcwLDVcritCTHKw4sytrokX4EOf1lXRmAhgnNzvpA
QatpiH+fI6aqxo6Lu8hxqW3QhzP55WS+rmbOr2XFPlRFsPWIHSUVnqFGlpZbtJ7e
mdbDzX6gFxaWfMOSVFJgnSQ3+es/Dzx4LmZLfu2TcG/7vdjchbbXbhzUXhYSqqci
tpXRlEpWjUegglwfVUcUvzj7kr2pXIr40a4s2fYKCyEdAnAO5Lqhcez6+NVbIy0v
q5mseoytnELorNGRqhTfmxYydOvYdnQJI+JmsRwoFWjJ3HJGHHDEAdgbl6ATcQ7Y
T2lD5hHM+N/TNtA/wZu8XI/GiLw3PbJs6MPT3pRowXC+nsh4jWp2hx9I04lrXBeV
fGcU5Gh3O2DnJBGR9oDvQ6g0BI3doKEHecKxVn2V2yjqgWltHbUb4RkllhhF6S8k
8W3Z1N+qBc0UGkfiymzqyksjItNpTVjuP99jsF9HBTnQsbTYbcKdyvsh58Ote8yJ
qnXUV7wt3QlyEOBJP8ToXF+/pL3JLSTT9bebSZ6UG7dAKYGoSi8XzPLO5Rq3zgGd
S4rkCrVwxEzdea5SbgyVHqZVDVJEtq0OQJdmgBomiUpx3XQUa6og/SnZO3iPvBRW
zJEz4b/a4hvU6mMUBujThoCYZkMqCI8VsGToInyODn3EFeNkMaSwXxRakDpGq9ks
MUYJEfqdf7yQKlQWMn26Cv9xNSez+2AtZPIioDp9YX2efZOfkDP1H/YvCD8Gp1IK
kmP8oRK4TzVLZ9ioDmJFPLjDUCWQ8212oMe9Y5UHg0yarSukhXAkSjXYWLqAEsWG
zhvUHq3N7sQ3HtQKJZmoB30X0OZCmN9WRK/Y7+kIlw8oPCrcEVp7l0SMgVr3MsVv
wwKfwZZwWESQFXYjPtG5+advGjRwkUodMgY1obQA3J1W4eKlB6IlRsuqDftOnSF2
kF69zCsuWPsQlPnUcRtqULmUWDYucSsJQtJGiEYYTh5U30sAYHFO3swuq0bg9O8D
6LwzQRZk1Zsk3VYhwMBnke6oM1XG7EYU8FyahBJGc0Eywex1/O3E9Or2SMpmEJcI
1KByJMaQFCCQfg4pORXSVQPsSrSSPVvpsjc7OnbOMWLVuQ6l13tr7TM1t6fp5jrp
iY8hqVKrqsDW1Se98LkYbbYNgNwUUU+8WeM1AXJodHBVxeTV4JCSrzQ08k2BbZ0x
yS1f9AARmXOShCp7JhKT83AD2jKoPw4sD0Ff7A3Pc75J5dbfYkY4abxBgnGHRJH7
Tf0jGo2A4g+SfH6Qn8OSxQ91YOvaKbsNhTpl707xxaAKHW268MMclQEpDwoZtAFc
I+mjbwviFU4jIJnR8ylhx/fmHrEZnGE6aRPYNfcI02qy3ziVUXAlwm2NuewMTQEn
sl6KxP0katpGpkZOO7TyleI5bt2xtEYs+m0j8UlhXJPiqaBpmMtOcmzgTXCIdLA9
erdtkLVDqYcAdYHo8dtdxvxYCvQJ+tf5kWmvOMSNtOaE+X9PJvj0FC+HgoUUIBI1
ZqLA/nNG7KIganWtSABE+6Mi+3D7tyXTAKbbj44PKyIBmZfbrJxl/0iKyMwlghio
MblWI9mAoZ+fGhbcgL345nf61bvaENE9KbAfgq7l8VvYxlLIOKgMOLCKIAhAqj8N
CYswTP3u0EYf5ZW55hzV2dMQwexxkW9AMpR/dxq+lIM5UZy1FsVBrrXT8TCbNlRT
yxzoYkf8F4X5suiAIoI2DW92uJt2icxrvbAciL7WfLgxNff7ZWzFkrd0km2akUNN
XgRhK084DczflfnfafZh8KDUzcaSo0oae+MpJ7mb5XItrxJQTWx0FL2P40Eg2bOK
BV6RAFRukNRElk/hTumOZVCg+UyWzNo8vIBwngdwLcq00pSZuqkZu9KB1KQc5i4F
0tUYhViUZhYurhmjf033zNOC/+9/vsFevZzye+ENjDeOxI90/MWRReGBH0VhZcUD
2owYql7jUOhFGqY0QEg0/HbgOf2NifrwboUNcB/x/E2EK7Q1xv0UrZDU26Ggqowu
ZGnjrIEuKJgd/1UPcFsKXkUeDQTP4LG4IOJHaKL9NINyl/OjV30jLrjvkK04+sB9
5bLGf2H88qqU0DeftqUgQQQVfb+/3Vx2pXeuDQGnxzkmzcr5s32c/EceBdhyBlVS
dsrGYBuW3iy5e9wwA/ZtzRV2RotmRIR21AnR1zNI3eI66XWHlcTwMfUZOIenZF7o
BrEVYMPaIPAEQLGL3ak7pGTHtE2B8OXTqluV0z5g+yG7kCfNwzNAT3laCK2xvK3G
0g5lueXqCM5NAcEEV6BMov3p1YCznA5LfG8riMV7fT4G6ogWEblZ52ywrZ4hjcVQ
FMhZc6vlqk2m0tWEbimteCoidPe+HghKEEcPSI5PEpFa6umoyP6FonaDJTlWeuxA
4xFBps68eZPpn/bFdDBkaJ3e3ETvLJ9i/Tu/gAE05cTUBBEobBjaiyS1O/2fwjN3
fBuM2iXo8yxmGwOXXQhqurXX6TMV5kYVdVzE5nfgwtdoEjh176bXpA8tPDh65pb6
eCIuiFmahiW58rPI8a4Y93uEDvI2OcxYL6uqXpX4V4uph6zgZkfFXWuVj8FvJ8ok
9IGe4cqAS4wKIf2ssMDddN3difkVfpqCZ3ZFRA1vSA+nmuY5Bp2L1kabg85vrbU8
Axgz7UkUF3bOlZjr2lNIarTclE3VuQDaQZP4ozR4LMIHVqLFvR1OP/fwoijop6Md
zzqvq0RGQEjEnfrJJJkah6EFb7cq/jfIg80Op8W4X4d7wBwM/Rx7dvm2CaePL1ru
laPk3M0yXQlITXEvyxzcpBEatG3YHih8FrbvVIrF/cxdCH+6tR+LGri2y7S7TOwr
ZGT310z8LK7sdfXUVrIB07lmWtNw6PkB1jOs2bVEV22EMFNwWwTs1Yq4irSFGqtt
mZmJ+l/i4jz3rsbI90xZwr2JSW/WF0ieEITBqFwbOiuGRel5FpiSHdN5N425IZGo
6DSZu8w/u3Z7mNeEW2U8ATrgXoWK2b7pGl5uiO/USqNYplWcwzGVVx/eZCKH306s
gQfV5MGxX2zzUWluxvLzj/a3ksyzohI+hBCTCmSNsHCxVnVb1xJFrcyw0xQaL37F
X8Hyarn5D+Bb4Oe86vww1++Hbs8U0gBVORCXgQICg4nHvJxzd2lJ8XxG7+d8O9ER
mfgxwihWUjs8EnHqXyIVA1utrIZSY8da3tkAdNN0n5l12t4Uz3JXw4cObu1o80sG
maF30PvXxs1Q+gTqrPSgJh6VyVa4oQnEwEJv6l3vhwsIQnZibmG5Q9YAjTloDM7E
6+uooCEXfBkJUziwSwv1GpCE4eV4HZlTPDrVAbiS75ywwEGKsqqsHCgkVGUouUuW
8+11IUGDlbPl+ZsZc+hT77RoYT3ByRAn52+eqVO8WGh3pI9w/je8fileMGsE5fLu
NrHormJRY2MB5fOojwQj/souvVJ5AgdV5Hq1TpHN3Dt4s04/EKIvv/6rEu9EHtC6
bMTGW5+TdwLasnv/WVJkq+M0B8698I5Kiq6quntAM0HHVJxK86SougZjlE/Cz974
C+UYYkaFw6ccqzKAV2s3TEzAoEQyyF215a1nm8SdkIfvMZckJl2dyb7rNWc286Oz
jSD6jhY3DqZsgEK5nCMAbyyyQ6vYC0zW37PiezlN7mcWYy1taucAaC4ddtZPvots
y9XBAWT9Ne67iBdwE9FQK3kiPVRGkp5M3axg/xB5uD7BDd5ce3p73lscaLVcwLKG
S6GXjTkxTw41i+kTfRg9gm5H2HymPGrqrKQc/uhK+iHNvhtgRy6tAo8WGe3+bw7P
+BjrPLcplTrpI8+gpFIZ6zrih1qFu/p0NLeKGvXQYLr3+VruweXtf8TR7W0CqUGg
rWHscuwGz56npDr3og4umoCpMp1BWhpshLy+4jUetvLebi5uU9TZzNgB/egsN61g
1h2/v/2uf7myK/mh0zq97HAWfpIPAtXmWrU7mwBZEJax5tHGozRjaX+v+hhwkaAO
px1SA6U2H2tpdxTMy82mArsYRXxE7LsP2fgmCFYOp3GmW6yQo9OOzlnbCkGPdVu3
omoaI9z3jWFzJ8twvvVSarslhDBFchtUqUDujMpnU2hVEyTJZut8LPOLo1ShfaHK
ts0DSE7eueK7RyY0Qukrmd3xYNupyQl8I7D0i+Mhu3HvhJRA8ycnF0MElYud3z67
+HzjJMkXh7gAprCnVOImsAoyyBjDEIqaYGfXR4KhXSMAtJbpwR8a4zGnX3kvyoWY
pwzaNLS1oIfhwOgf6R3vNBqIl8KWSiE62X2/E/ULIDbXeOEp7vDvTtCpmIw39xji
9kNKvRlKzqkb+/zD/sRjwgACtinOlMsL3hBnDpTQAC7y1vFWxrM2aaJYKmRQW+bB
7YymK3rJce3cdDILPjkJ9pSPAX3deWCEwXVsNyg7GkdQP443QW7+7TGso5npA/lI
d0SW62yS4TlYCHzRo9b4JIyXhQri1O4n9UXt9jik1reNs2jcx0xffVGKwYA3g4l/
bThLTNTDuYRHieuPgNX7QNX7j61/4itXUyGk1SZvt6ln9MisdcxFifhpUTi2vTmb
yvVqVlw/hLP5MmhtpC0toP1XyZ4r92z7L9OXyDWIxrtT1qMtEPgt9DBEEPs6m1jx
Zic5zF6e5JKNZgnSSjJVtLbpYkkmErdT2hUpmQwc1LYBOdIWADOsqoiqhkMJBK5s
hdA/7Blz7xYnEKo4rEKTFh/nlF8zRshEbCWHfd1QCnjr5XvbpuhACGoWeH9DrhAa
ARFhgSlOZN1KJwlMGeawVmKucKyuDpEpoF4Yl7uPSPaNqgIWmYFd1Tw0FMPRN5gs
XLhJTg3mGGJbc7KGqoLthppcvaoncPZR2ckyx1/HFmFzwmE/8s63pgIHLG3jDs5v
taclbUqP/EQY71U6bW5OfDdjZKNLumI1aoHWqbND8Q12k1jQMh9xI4HXjys0JNjp
+4qGDV6nbrpNero1Tb/Os3BZbr0NLldWul220Cx8Kaj2ik9OEUkN/7CIdqOBIG8L
tPtUDfH5w26Bh8wrE6dsgk63HGQZ6JhmmHKeeHn6K1yVY41GyzHz+BfJXJPiqpeF
tO/YcP6+HuVQOsBgd8DrQczL+kzhR9ykAykaOoOaMGmFinWD+dFdpRGDnt6+ht9J
Kh8sy9GrXd/31I5Eu0DjHK9mpTJCG4PSY64TLm/JG/4tX1a1bc14M6zzmXSuHd6Q
h3L3bYQkP7+4LR7meRZ7F4xkaXbIhXfLfr1lpWAR2P9r7Bcnn6g7oM1O3T8o0f8b
jJXjVyzC0Dei7EaxyCAlvHf0/+aLQiwk0zgvrUKeQtOGMZMBe8PPYBFjs4HTWET2
bOrkpdNpwfRCJbX18Uu95yVj61ndLu3EoQMTC1066z1W5CxrOFmHIMq8Qn6bzr9f
5ITx2DEx8wOwprVnAbJ8aM4z9JOu7hXIWsJMnPvb9xQhicZO84qIZChMYtPiEuuk
tpvg6udOwETAHXcCuzNv0IRfSPYcrH18m0uGvStncUikELio8AyAuSaCK7mMQGPx
6PId+XfR/ieUoDk+tHBD9HKQQnmpua6kQ/8rh3F0H8EygN8uQ3qaxJ+CT5FuT3N7
M85UY2bmMX8GEdH7lYSwV+zc5AE1YBwN+S9ec1xf2MPh5lpQQ8DSEGdhzBbEOf4o
5uZZz08+/cWeTq2AKBNmSD++bB15X3JbXrQSX1GEsAK281wXm1d486qYBlQyu3Xs
x9al3gGUsPEdegMd/b7J12tnyDtK8iJP/RxR6ZCSd5Z6nXLB7Vd6piSHbRZ+n1zu
IJTo7fiLEagXuWOIkvlX8vmXI7MIUz/n849iXuhGMT0qKjuI5qESLOXhe0JhlMTI
1JWv+pcFnfiX7iBBgNrZdwZuXSFsShlfOxf7Y5/2Jc3OvUt+2vTnrLh5q+dEi6QD
373xc/Y+7LcAbmDttzcVcBEgbDWfXoJotaB/H5p7BmOV18G2UXtVXkjrfnzBmPNf
lfsw8KPDjJEnsaj01eWzR6BNINxk4rQtLc0/0sCgZj4dJJ1TTme7EgSOTpAWiFUI
/6Tm5s4shl+Qr9hxxFm8vSZb53nG/jACiHfwiV42dIYiHaJ5nd4z/6QaTnEYN/h1
Ti6aGbtMKTvRGmg6XHcpEEcY7AFiJS74WCE/aYVGHjp890WEJ9JYV9lnyHlxuDrA
aVpTURyAMHbFo6924DNd9IkPSisdfaEDcKnPxXECLBrgTVt6VUEjzkbwOqVf91ZZ
zZLWU3lELsEcqcmdZQeZc0MhUERmm3C2BjK1fBVE0LQOSo6IS8d0g463aw2Aa8R3
hQ7jJ+FbLU51GaFFB9u3/nYKDRUF2denR+LIrXrZuIB+moKfVFg2e/pIe1LqDKQ+
G8Dc/s6BrbRoR8jOTCQqMPwcoI1kTDYNDbHEUxmdle+CeOx47//H1tqoAtLH+M9e
XwOuHrGcEZGI9fzvKMzTXmg7rxRpU7Gi2wS5pGMky1iIr9vlrCQ/9yhDPAMxxxg8
nd2HUZvEVADYitIMWhYf3n9HKJgrGsMgB7h9pRUZaN1DlB1w6DX4Xp2hwAsJj8Ht
rp/Od98TfUleK2gW8TJYmH85yGcAjYn02EZcCHTtqCEyaBBIBKUxLu/oYsoua3kp
bxbW6gUvkAsjN3FVwqgMHJIQxAKkvIBibvshn24yQig3429XeG5QyvTkXZHFb3GO
ZGy9DFpj5ACO+DPNsYi83/QcN7e1rh3rSj/dqRtiex+tTH8X7D4zKX9e6DdbQNHJ
oN6lImifPr098mB29VmQGF8Vz5XZ8TylEpAJgpkt4n+3c5JiDK0rFoDM739qwnHK
uGP80BDqrvIYBvRf93svghtYpZEmM452FtWNc4Ws+ylLY1iHdG/MOkmW8WQVKHfH
VmI4DkjW85yffd+sAmE6zx+VJNlMnvjOeBYi8YbrOxBeeaJaon+Zq6JFY2iZvT/f
Dk+7lNDKPDg4IZjVxy9pQuEYbU56lATy1WAn+yj0qcJ8Hk7TAtESJCr2eqI++QFN
jL6M9s6WrheHiwdEkzKtZZcE6n6/0cAr8OJQmtZwk16bVAnBAUiIpubazJrwqQxJ
9x0sizb+aXMUUP92TMq9I90UJv7fdkjrKM5wahQX/oMfPUttg42NhBtFzc7p92Vy
e9dvRjBWSZul8zXXsyNZvBmxBSqPbvbEyFxlnNME/g1K5JqgVxeKchN2O9KKDsel
I7/jVgogRaEjkQ9cAG4htB6OElWbjAMCxfElTTmk43ZsDS2te7ks8DNFPL+2T3tL
RRF+fHa6M4U5v+ZWzr1486z4VFluMwXzHspC4JE7DfcP70wLNRnlsCVCalDb6MDb
uOT6xIg+Wm6ZSN7ZSrYCPs6gNG/8l6B/CL3q2w4HJYKDLs/1L0LHee7zBLy8rfB3
vE6iW4/AqIcriQsbCu0c+Es4QOuUHJnWegKuJKQiQ4oXPj7E9SJ3YDAfcLM2l8fJ
QycDGogT8GWmWn87hLUJsEQvWCzzGa5pKnQK+WD1zsC5fHfGm26lizJ3agc9+CME
hwXtKSWlBJTALD5jwHJ7lYgzdSb1rI7OFFBjSXwwFJ8UZuG6lw4TJax9zh4hjyru
yiA4Nr+vU6qVwC8bUGs+j/3isnCPYGaapaPz4ol3jzgEwJeiHM59m3SjNiuXVgJp
6sb7Aq902jE06D2ZgiReAaALXRpJNYFE45MKEdPq5qGPReASEtiQpokEeOJOGTtL
0yvlUr8aTo4CevmT+DltOPkDgPleJXOvX/nNT9E8M2i3vxYukQ3voRoVz5gaQ7TY
cIgfMtRDIK0NM1KbsQoruxIB2wlwqG6ATi+nrJfLycmBC2D65Pc7LJitNjGY7zg2
HRAJn5o6TcTzukTbxbnoohjpWKt0/JRuFmXzVQ7kXAUhq1MtWrXbtlXTr8SjxBN6
f9LqRqbHTqvvqO7Syn7Ox1eKBBXid5Uj0kl4D9wBxcK5n//u9mv9Y1sxTk0dd7rw
xZS6cQH13swTCRT3fZNGJnC1Cqxqgf6WXDOw9EZyLAVARr3w+VtQKOfsL6TYFyQU
AhlDXqgU7HgAuqoKRlgpMIKzeMfzCDxAw4NcOEyDW/mNeVYcEzGXkxqbG//7tH/i
ZPTJGMCv+zRN+4nU266+KGgg8t53ywVQEI28w8NlS2XhjEbU1tq46TtCWDRnD3rO
JFLLj2dSN3p2P8RYfm1fBctFZi6w7UwjE+1UBhUVVUcPyD9iL33s/geZq5nNXoRw
M+Y2QAC+KrX3m4/RjoigFBnnJjsO4bDV9yARrQvWppHRRlZJz+2C8BXRuyScZIgC
OsRVUGqH4w4IKyQWaJZ8QF4C3vdw0sYRKd60oz/CefEGv5SLpj6fgBD4MHhVC2mi
+tWqbpQKyKlQJoKR7kK8KFu/qDahIFOr4hRhMXYr1+TMXjfoZt0mK0fZUtYDPu8X
OdfPfyLQmRaGrtUDeg3nw7jZAi2W4l9l6Dv16372j6l8XVOM5NDdmhwd6WPDYxqG
dJjallS0t1G8HF3rig8PrM+9tqRA5ScsWTF+c1hbTD5U/MHDfDEFkeFeIlqhodMd
N/PFYGfdoeM1CQziJJSuGq4XITGGGwWGgxewn9ml2xDe5TtmGQef1BstD/4t1KWE
d/JTmXseqsK4xboq2sKJGj/A/P9BEwgGoPGD+SrYoZLSDf3xIQlgVBYxuminmywl
eV1G89JXRjj8TStCxKZadvYl4pqoYU0MlNkxghWcjueaJ2bhJhrP3DX3CGW2HwZh
9nmbW37p/G/a1JphnjqbbcZPPMhqvaURfqkZT4dfnBQOT5nUvlCxaDSfQOznd85o
UW/uPOZKDitKXI/xApSAkBcqQiLljcyDFg+SdVrUn0tndm7nSCWWVnfHl0ewzv5n
dfbHq9o+Vb04PsN073aiiOk4N7a28rIj43WnGynyKIm+xu9tkyrXbFC0Q/6l6p3p
t38Q77o2joJeNwTMd2fZnEblUoXc9LXhpwcJFFlh9If6A5123ubW1Ru4axdRZwpF
5aozurtsVXoJ9u8Eg5Sg6JlZ3dbNxD4YtR4t1MftTcm1Ara78Fr+faHVKouHURaO
3XEakZv4S9qwN/9J0kaForXCAQcDnq2D0K1cWsSAhzzC1Lwowp21r+fU+awR8VVP
zTeiCawXpKmjKhH0R2wG60CbDP69Iha4WpIXLGPSTXTIFcKNtwlMrhuvQorI7rXi
vpkITmYZQYD1g5kZaZ1vWuTVMPz2NplQ7yym2QOi2Td6JP3TehyO66aIPaLPf8Ws
A8r766mQaLzxJJoV2+Ho9neNYCEQE6Xl7Gy9K0NVh1Tq21080oBAmMi/L2EL5z6K
S6CCpYPCEWdI9vQuY6PGlvbAI5r5FBDxhdr487o5bhMpjL71qnT/cxSaWcjMDGbd
dvF0fkCHJbqpGmggKU5S6C9FVusSGYKnW5I5e7HSzGpWlueN9tbG2+4efXoP2kpi
4d5hxVSGWPYdpTp1H1T2vudFcxitbjMm97sYEaxXfL5UxHl0hR9mNliFVDc7lRIt
GCVKau7OQp5I1cuKc9meWRkfJ9ssKsTdyuJNgzDBNYYKhcxbNVKE+92T06dyALrK
YKKW9oe9hZynEuLiEoBz6cSrs0EYhQcoPedEhjyu6cUkPMHRdDpgLMsly80ZyE5f
K0bFx60WyeXoDoFmNEOWo7uX3kOL20ieh62eAmvXYIIg1jyXDDMWGlUIPljI+AKa
95OMNJ6RzsNyy6Ojc4SDpsX/ED8mfHDhHOOjPMSfatT9UH6Updyoc/PfHg3PpSez
QdnBB9/wMqxZFDTFSLUFDGwVDBsHKUr5fRWaXZWOql+vwHZ5Ss8qsgF8Yfbed+Fr
N8lq1NqebY/fRKHPmtpFaF4veyuu6YkIjunRhmroUAgqrW2tRKvkmg9gopzREPqO
2a5b6szTtJ00E3CS93SXJyljm9sFho4ob79cj9Pcve6IKk68oYre11unnwVIZujK
ZD0I2HaL0KdlugRs2yzOeIcZgIvpIWuZzMq1LXRQMXKCOj2pbAYbgZCzZ38A2KmO
zm3VUZ3lPGqKKyW+qcq5WB64a1h7XQx90H3dKH/25oGqdo27nMyU3NMpHWu3I5JQ
01tbjUjj+6IrmUIYVx1YyzoCMYzTbwKrgz5DENe1maKt8G43R0N88cX4CUqGsa/Q
KRDyoOWfOucQzCXEUzv1Z+FtIML4iZ3sn/PSghjjENc27fjGFeY5BJl5GrWgHtxw
oQr3HStUIGZQYILZRjLBuocdoO2rxg+JLQDSevxRHww/L9CGnq7nbCMsAh+BGTTe
7xIAcQb8fXIOpres9/EhQFdF5qE1GiMiBq3dg5PN6USzT4Hldb1rvoHm5PeABaoe
r+dt8U+huFL8+xyatrbgGFF6QlX3Blkj7X2sNEG+ne31LCYidlZ1ArNGO26Ml+Ss
coVxaeZR3tF99gmpV82CHr20yNy5iO9qBl6kkq5ollbgZd1yIHHjl4OfjvKLSvXz
7CjQsH6gvsywNYSsAQCbp0cX4z1rlFvRuJpwj3d/SNKKW7YmIPAowW1HOHKbdTji
6xE0q0MZYjmzad3U8anNyNaNUNuoc/3LCgVlsC1yyS3fvU9/7Xfi8k4UrCbKkzPs
IJm9MnPYyqoVyL/hRIyDA4N2gSIvFVqKpaLw5mCO9ZrlhEwaBzIwTvRHXa7siNDm
ZgR1FruYKFiSNmnk65BoIj8Ip46If1br2E9hTsvrucvgq47OB2w3WBiuFCbKxGIP
06RgGCL1o3JC6dyjpgovkOIc5/WMSmhTL5jPph7E74tSu8TLoMxlFG7ngwkFp8gq
sskCxa+xu5CsuJdyGhb5cJqUI7DosiXMp2JI+1ZuKn3u3mA1mrG79hk3ABpucvKE
8cVkx801MQu2hxADb4s7w8IPej+IiDXPzKT6lRMf2cE4uooy4Kxk5t8iehfy89Dq
A0lI47Xf1VEdC9D8V3VltkMLDgFtWR7HLi1Az44ECtjwd/bRIG9XSl+QIzy2bbWO
gF7N86RNnSStk6RYSjK8E4GxZDJSuCBZas6v+w5jW/uKgyTvR6rw0oaBLrLjY0Mh
uQDG5i8QZMiwFsOdGSLZMVGGLGOzz7oZl8pJjxbuGKSWaM/G5bYK7DoLX5biaszz
5KKL3O5icfwOsCgIsjgXi2s7WFQhE0m0yQSTC+Os77jEBXour7M51lNAy0HgInxV
/bkdOfNEsCYGMxzxPFtLUby+BE10sNgDpobLZ857DAvDuSnvcABmvCm0140lDU5G
P9p3aGTf/m7OFMO5AwQCfDJ9wCAWC8TH6K8dKWMOtrDknbiaKjmPoZJxxJbHZZGQ
wV6EkdviBvVlSyNOYfIeqpxXKPC28c2p5Ua+O7ZqeUCdMlxGKhMsS1JU9EpCHXw2
FynFvlj75aKOZi0D9hFgyQQ/+k4pbumHf79LnRds0Cf7T0qSIxgvEKAcCLkq18gr
TBeT6oqgklukRnd7jZnVvA2mpb1837ed/KfCL2Q6V1U4y1Vur73KpdEMT7JbsSSB
yWCC40g6z2tH5bAITX8s6KqN3hk52wue9LFBM2MJI7CNWiAQPpgoJIhnKniRiEjP
oXDYssYFxluNvuoFM5KTZVgFuPuEkpC8/FFNQtzDuu6YNwPtyU7pfn4qhe3ZIzot
3i5wKRtdIVJmUT6T2hHrd+MWUBdnneZe4NtniT7AKRZPMqCqaFj64fy2H3m2k193
H+zzfoHcwETF85EAbfrpCWkAtiIeqX9XBI4C6gtBDxO6awwQQYHAt3e034IuMt/b
9Bt4KrTjxyW1EHBHpqNZTWBZg2x4CnWJ5xSw9aTIiy00iHY1hW8Zrx0T/6xYae9Q
X4KiZahChB0TmVOA5xymqdU+lllE9QJ+8JMr+BlfbHqHYwgbsLl1jJN7PjYL3WVQ
3sdhSB8VASXPZ+JUIHamBsRikSmj904Yq35wgjMcgIcakWWgT5cQ6stjNYWwvZBy
aFVLKUJZZ1oXBgZCGHm70r/5fN+cZbf4jmiDp7VfHWkDc5CEXF+9uLv4JIppuw7D
+6Cu9651zSkYaNV0To6d0KryYuItLLS6rgNmq4xHUtgDVSilh6ssnAfagkZcOwVX
cMZVG92B0+EGSR2SWEDWpqDWOgUIZ6Rp6NBcMo4d1uFBi0qm6wcNQwdv+MSnmdq+
NwNwVdz+0+dQMc9zi2VrQe96oFQZERtAJmhX+hYhogoCpuuKo7gIdjV+GDpTEnGl
L3AjSTuRAfiE+VLHNWM1NXjxGfByaeXeM7M4Wz8F9X/c+HUjQw+zGtsA5HT7UYbp
9FW2nrcn7P8FhuPBhWJfE9J639FniESdM2lopsC7Nk8qZ+s02IB+h2DU4xKHVZwc
lJLJraPhQWe3crKz0xm+va0QerHe7kDJOm9MPprN0IXnc25q3nkknHtOdW6XrQP1
zEZ3JCCIypCJWQSbSzGIzsEhlpSTVR8AO47exh5djfH8PAaPxJDr0P7fO8ZuB3gf
dONFyskkYB2EjRwFjnqJEVi5XIZ8i3Hr11Z6WedB3NXHNhimgrsaI/0bNK5o0lTQ
X17jC+m4uqLO54dv3gc59x+rCDGiCAFdRDGue6ZhKSEFgWxZ2L4oK7AMySnNLs2h
5rd1yLsXdIR+xbSLpgCRGy/K+lAVNYlJkHWhjB/G6JzeO5XqMV6tbfyTIB023Ddj
xT0Z1pzeAeo4krSOqWFCFLak/CNhWD4j7hoePZJJjE6LQKF3yk2vVqvXNku3wUxS
x6Fni1JZeU+vIPhsY/Sqdj7rZdTPDO71BRxmyqk6YZGkrBRS0crWBqNse7rr5FuS
h1phxBA+1e7h/sCVUm2AQ0ZF9rzW0Y9zHBy48LmKI11YCxrajnnouZluFIDzjMYX
8e7pmhNtPqswDOhR9nE75d2ye1KCkXbu+dsW6GehDnULHptoPo558fr6pxkriH5P
wHaghfTtjf1nNnpST7Frw/sfscvG7zmzmKCUOlaGQwB0Oo4yOE0KjovGhEeZu7R6
igGgMIg8++ntVbgJbFxqbPgjUPkwyYawtCqNzWoP/OyWUmwbGjbf2mSfIBkivFiT
4pMM49zXagRC3ZttKtscp3wyAygm6DHbsRLWIfTdyDTK09lox2ciLOb7gUKONPPk
rNoEvgPtWQuq0pjgHkR+TTr+sYYH+WDc6E0UDTcMcosuX3S/7bW8lS6OgfXVr6ky
McsbXWhG8j5Z1eWUfMXwNVLkWZixIm3icetRdEzCtJE08lKppDNxvESi8DP2/YcE
RMFMFCobkjiLIz3yL6tnFmDJOjvBal3b4XF2VbxnRRaXaIquKg3l9hHXFM/jyKTJ
z5RF6VfquCpsBvX3j2wWXBxhZCPxXUlfcBQvjdve+UrEkG5NB9Jul0UcwVW/o+yO
sdUciPOA2R/LXU94GCYYnkSi8K5KT9rmD4A+IJnQkNl8X8PuqL8Wvs7285hH9jTV
Xl0sE4mvX3BstlGDw5Th4B2fnzm5L4sfsNruX0mXde8+B6JLOrOESz+66nx3bFjr
DpHLmwbfHuu/9lDM4v8tDhTpJKwcWTZOHp4QDcfC08fYchXYkr9d1aKC8CSPZVQ7
1m2T17su3rrMl/AT+Pt+giaI9qiA6pZCaMKhNOhsasonXZpM+Cuki9sjkBWTATJk
udbD/KuAk5ZHQNKQK3ZyZUyZUpx6/Z4AVmZrAqyiTc96e8j/Ta4S1Ch+Ea4+gz9Z
UCIzQ89YuguvGanVM02DNQTZYtL8XvYykTz7ewf+qq6HgUzvoj2E+zRC33tEkN4l
JNVTMESFH3MouHn2ae09xKrOwZquyD3eeoqndxwyIRhUGY25TxVZs+YNNOV61/UV
0OdgwVitojJvtJ2tX3Zgg7FpzafC0PqWXoel1AuyM+BLdIPJkKS8ubM8gbI/f4zz
DaKh091DG+eLElp3iBA7MhyqZez5hZG7JLBwAwNR9qzBN3T6B4FWgqf8wAgpyXyB
0uo/8f6Qb+0gg47HcAkQ8kNVO9jvfGntNgZzIQkEItZrclxu2W1B2n2A5aEydFMK
aFSgSTi9hb/T8suabfjUxDgtn+Zl4Vgh9FwVhnzkSaM6TakYH+LBziG769XvEdew
MoVDHXBZ1lAF1XqunFuhr2gFFQAxmsrI/J/0By5iWnLoTCvfjWGq/jGuDAbvFc/C
8612P4VL2WHVu/rt36qeVr9f4GGlKdVyg/j/i0cBwUOYGN+lgqpx0XQRigpObqsQ
s0tTjX3q0UMo1BXCqIjQ3zC+2Tr0jMg26eE9uHrJYHVSj9rU7bxeq9VFHYN12HL/
P6vWveI6FQmNP6aJ0QHrPEiMh84fCt+/JlXDhanuSk/QFFK+Q4F0HD4d+2e52PQp
vBIbvXspr0oErgTmci1MQ/iiM5jM3yjHF77WN0UhGeSym5FJLQL3OZFbGL+k3y6h
gnTFyz6Fp/uTr5unbLrOt0cByaKeuLj7sAvr7R+kjlEMb9CWh1C+buJ5eSVPgMXQ
RbzifpqUmYmt5859WnmdPVVMXseVC1i4SqL/+MVvkhlQbzyUdWB5rgfrOhsGGHFp
X30RhFlnua+xFYxN8WN++1+KI6X74aDY4WyyTOsWnsy/3oNdAKHFLPbLaeEJYPra
vBOhI+ZSHRgsbPDke2s/YSaoPB6mWcSIfAtkID71ej0uvI+XgNx4R+VaV6nq8iwm
+FiEKYsANqDEaiHhHGGm7/PEic+3X7H+x+ty5At53YB0RqOSAbD/M25AyX/9L/31
ZVZ9nhC8TfWQZPsZKem/QO65gtc821G2NLQXbJpGWUCpPARiCxi24T7imWrQj4Vg
MjkEX0l+fCCq+D1gBcESaWigIfG00ZHD05gcr42YAv8Qg7dJuQEqrtMrRuc6dx+A
VwKKIGSm+LqR+FnHKdFnJegRLAN/VPev52OpvkPghrLzOhcd2tPFrkmhNehnBP2M
3MFmo7KRQpnJUrb9hocIULjHr/V+dghEzjhKKy95W4qG/AcoK4kd6OiPXcHElIxN
aN1o49h+H2bQGhHGPS5150nSpThRbK87ciUX+NBKzU+V307y0rpBLeOTjgInaLZ+
2wUG7rFFp04Z9BQHdZIWvcqfuQ+LEv2VMz4RGYfD+XaNyiJBnlfRp7o/sdGSQ/8S
FtC1nDJv1eOlRBHpc5kxeMrMOmAIbjFumiTENb4HGlGbFFW+yX2qi///piPt6rkB
dB7SPMAZwuRSSMBj/NFARjl2odkUQOcLUBZhQgeXCKA8knt8cGRz+as/75I0Wymw
mItc5CqbPTG8JvB3xqUBGVANZEBpgyPBYUX0xe4UADZ0MwS/E3SB7I4JX5XjPPXu
BkqwqR4NgUErchxuUXp5dy+qNK3pgbatHboz9jSe02GOVRPnXBVADBqEebyM0diW
/YpUR9w42oguyvN0A8SIjp480I6KT8uThLdU7tW6AU2r+oRE2O9Prpujk6lYu5GC
69yvSVT8kamUku8ZvmExeREr7xRIRMHx6W6KHujkwUWXKqVAPgQAWeVaFM5H4yu3
8edJgENCBhHvGQxCnywPfBwFnlWoUfh3rmiNY1pieDH7CnXppxgvVGM0ixdZkAtv
W0bo8aqLyGY272pqvRpKa2uxL1o06L1PJecoVvHSLPYm4tsAynDRckVHlur+rhd+
8YG5Ang5wCa2b9KD5LyR0xvUaYHdrIjQTxy4fOUpbSQbyF2Nq4BA6U+rLaPJjOZu
SQYnPNdRMhy0frfJwy0F3k66q+o3pQ+v0Moh4s0QnaD96+6pFraJJtdbuKOm0IXO
8NGOjPklSNmwPKJJSJ8vU+m59R9Law70BuD7WD3Yh3tHi261QmMMwfM0uDSaHiXJ
RE/ETm9/4lgAOtwIymbcNnYL3+/04mUh77gQc/qgMMoLwpKYLUhNKvBK78LFZ4w5
b2KnzBvOQiBuRXtTdNF+jbG8OTAYcWQSuEnUqmRjG+MGV+4gYsumOKvAvwSa8c4I
6cN387XEpZIcXtoTf5os+ayIWbiazIefs1QnHN0AaucF19+d3mXuD7z+kOQU6Kkk
ZOeNr83UOcMku13En260gPxVe5DfRWfv2lPA2WmTzEuzZ8LrCZJ5UlfJX70/kAQe
ogdJez0EmBiFVtqsQ2XLgrG1kpTfbchc4e1+BsVGyjbwAZYUlq20GBAmf0VdLikx
ryRhYN4xDtygSliKnIEHv2l0L9zkXZSLBjbzhx+3oZN2LH2eMjU0d0u71Ra/zwee
6NxPwkwJrwuItGXbQNFATJB3yf6/gAT7jHVdJVJeJ84Kwg8KIEmrpYuMptVn/JpV
L0LNg/VYDLAhNZKYpi04it5Z3jWc9bo5SdYvZmbr+LQ+E6sKYEwYyVJd2M5Nzji4
nrhv0n4vmrj1T2aJX9LWr8mCERWpWXzfws13Y7LqAHY7Z2BKCTpFhUbY4Uf5gdtw
c/vtlpppNvgfpCxCnvBQlF2OcjrH4LuIKuoHca+9n6fDroTrns089X4ivoQW6TVx
oVOQKIPUx68fkBv5w0w052u+plSuxBbYxF0u0dY5D8RDyhnkd3qCYW1OizAM2M8i
UhoNT99zUs9javY6VZza6bbWNlpkp6G9ibR5nUodYDEUF8ArOs7gwvmtmYlgk5EU
8G6Mb5uF0BZiahurD6MF0ki2hklP71YJlA6Qc4WEG0rtr4xSNIZ7GE0exzHIYCt/
1nI14GjMCfF/TXBKSUYf1ClAgXuma4d0/VXL/ArJIhDmX/qwL1xjFSeX+zRK88VK
rSYjTgyA1tWSmbxyRbZevGVIZz+aiKKZiCfTdUfrYEUncrG6GsWJ1BUQFbPOCWZy
2O8uC6MqzIr9uQERbPB4Hg04awTdt02hOvq1J2pJwEjRe9tfMbFOFoIXsxDzDhjq
40BpdTMFl1iMLG8o3s8w19V5a8oMJq3MbdOoWfWJFywTDRO8uX4ZdHJ5S+yBDELF
BoNDfWfc7QKkNLLfV8uJJCP8bDoooLcOgFXgPzqOEu6e5n4sX/GhTynzbvQgckW/
Y1j2vAbb+9M4WV3moMkPONfaqSMUkZroYfGeuDTYrxD853iCYX7k9Qr/vJ71VECM
Koyh2W0AQfoJ327A6HWG8agHlnSue2a1Tzi4Br2OK8izMgu7q/Mu0xx936EgiS8a
8ZcdgoHPN3DBsyl8QK1wfv8Q482m+YC1meOjoxhw/zfRahMSzFk+Do390MR/JdJl
qpJmfmraL4pUKRgeRLxOc1HoN/IJZoeNBHAYgtiik8gUJ6g4n9GOprfEJECskis0
Ae2hMgHoMV2McmvJGRtmi77t558k18xPYa/KOcmyD0lkQS/FVnJj1KpIAdPFy8k5
IlJYzWNhmzKKwMQGR+EaqdfbyZQ+XU4nnnUf0XUZ8EdPb9UPvLZYOSik31Xsv3eY
NGSi+sqel7zzre+LMuvmFtDOPal4MYirtypq7uor/7vgK23g1wlLPJy7EyyJK8rz
h6VFMqZudoMtNVf0Yc/F5DMsTkmJzAgO8xyjpYim9rkFralaPCVTboXFYPWXTikw
i8vsnWn3eSkXncBFNwClNqa8GSXzlUCMV/8lFmnNv6mS4Hh5Ktwd12fnNVl5eirn
kmSup9LT096Pj6g6o0xfIWDcIuytU+L/Ao+21+zRiR0Vc9A3wytvQ+E+TH48RYO+
Xctan+0NafXtyKm2JmZOGr3y6IjmLAyQ1jcjt6jE58ESgxrpfwKDUc8V0xggxTtx
5QCZ0CiwYyp6GSDyQfevqcOTmvZIa9jBflSPU1qwFtWkj1SWZqwXWS/oB1Lkm4mo
BOh/Qzli2fQPFWW3Ty2+6AEIm1wr00g99r8MJV6WPu4XSjJXhnfNg9Ezwsfh7bkO
zx3TMB/GgvENS5U63Vyg5JwAT7uc0v0Q3MD8LEThS/3iWtMbqjEt/E+IVmBKNSQf
xLZ3qvCzLTSTlVcbheSovRpTDx8p01m5FqRirKJTp3hp4L0vzro0LglQF4VAoO5o
OHsnvQnczFcosJUtUfb3ypbnkMjWU1ZMIPGVIuXKYoOIWibjT8AcJRg9Og4DBIDv
S9GphGLEXK7XW8O/gtVT0478NYI0gsqg9fPpy5OAL6Gzh5ro1nTH12nAykLPfZG0
CRPYijCD83Rh9ay7S84ErmOsThM62Z9gV+HzxZyEydL7ejIRFLJJdgLER53wzCp3
MkcEDotRjlVRuVPdsvT/SSVotgj4ERbkfw7P6ookd9JVvbzyiqW0t2ksXoRUAqHL
GQNwA+bAXc1lr/Nn4oQXz2e1xBUX+c5sXnOZRz3h5XFmyoS7uipJc/SCJfVSiZ4x
1+8OGdbsu76K/HPNfWopaHQT7vyKQLKHvH7zTdH4/OVXA8l7o2HlNSRj79f9Oecc
a/xuTmCItwC2I/8R+hxqLk+4YYECOaGHXl8PtxbJOdxw8XB+loZTK7fo91q56w3/
9eIm6EWhDwekHw50EyeXQyHbjJ7aP2M2qPX/3Mb0sKK528mvWitiD/IDvvAI5cAS
98XVwiKWpH35b29LPv/PmbfQ5jN5i0G5+W5InbflTKP5UJIBG7NFSM64j4fctDhn
Erxidv818jwGqE9qa6qASEFxQ3jWzAJiMscMs0GHazYLsyGyH+9NnJkwhnWV1mnh
NpBOiDzdIIeg2oN7VmckmM/Y0qnVdybuedr4Z8sqcoJTkvMNpkCnO11gOWSHNhBU
KV4vvmTPf1PhCAYbnDpXZ++vGAfkVp+LWpMxmuNDEf3EOh8iz7iMGMhkP+EaYO+D
rIQyeiEXed/+AuCB5pNqPW5/AG+mKXHnrQUTw0MaInFUltS8YQ1CV3S1A1SUh7Pl
5T+NSyf3L2M+LK8bP4WwkFEFOzmyGa7CWe6kpmBOCooeZ1QnvLYWf1CL9f26isGG
H+BeuVagTqFMV5nanEL2vjh44mGLdEbKGhcFwu9HPbr50t010YN0gTz7se7drcA9
+3aZHPS7zW9h9SZS5Os+Mi9qNP/MVeEelqjAYeisxW1+Qzo9PgEJ+Sa2wqIYobZr
CiL4vkXZa9f/98U5/H22aNrcJ9wwnmSDXS51xgAiSevczQ0IYLUYs8nfJqDPM8LV
UhqCNV+WoDe+IzesHgla0Y9Ysx6o1ySig00kzI4mwhW4PMDWRwRPGI2OtiErVcE1
LAMN9diIml6j47mMaNpDiaxhKAY+xyP5x/btWBCT4UcUfnA1cDsYO2ZlI3314dcq
ghYdHsscgS77Zm1aajvdtfBoQDxNfHOPZsxUKwAj6tcotMm6F5ReP/VilIZ9X4RE
dhVW97TqXblpeVxXCflORDu0zvav0iwlFycAXqFDPLvD6ii0F9bYxvEFG/cmutfj
qG3mhNjSpdEy5ku5fAcaYdPRqZBZztZ2GLCExdB5sYuKl47df0gPMGMwYWrNVGPs
TVytuTS5Oc+RyQvGcW3clc0eFRKyqMFwVfYc1M/5rUysxtL7SPnnnECWnZ/wMhvt
O/fR3YmpJ+d31FrdifT3XVDDIV1xZgtpLhWdGcZHu3vmRZ0W+qklBFVvTXbMN0AK
n+YsbjgwSkR6vV/yNymrbb8wszIEHgxtqvpFyYdZ4MHQUGtUU+MuS2NekZxiowbY
/B+CEjhJ8lDmdLjxNvRdXmUTURyOr0yxAkvZkx3vgsLHOx5TcBONQ0hJsvv7CjoF
/I6yJulc2CIfJ/B2UbQQnSKstYMUy9M1hZPoZL5VSTSRFv1lppDQ8rQmIj47NVLX
ZMy8XeFYQ5s9tF1hjl2oCBQ4ohnminw3R1h6N+KBx8uSvVAs4aKwo/5WysEVgr37
JsYI412J8D4Rj0KopRwHeZXR3IV7AWV2BVqMxuz3NeNfAMrth5jNB/7T29EAU5Rp
mDH/sYS+CgrYMyOTLfn1Txb+Yl89NNyegOR9HTtFFF0IsU3AkoLPeyqlMhi/UbJK
NjY+k5shmBpU7dx/ezXgxJx9wOIGc66NJZrLfHQSJm+m7fKS2SIqqxzsWCniSTaY
Ti/LfroidE40YcD5tx4nsTqb8hRP+KJfn0FRnpQuK5lcQNNtiRdO+7W7mnqZeBxc
VxUNR864lfrneq2oXOO8ucJAed5fRPrFANBC/AEKaNaMiYN2/I7dv5wjOUba2RbK
TbuETC5WqYVxeVOZZXl/NNWLi0Q6hTz1BspiTi/VKh07hyvJVUilI69cCqYFLHRg
xjWq6nNeeHRI695HADpmNv2ZwoxYjN6bbOcZ6CntlAaMEfLb4XpbVJQS9yeK1cFZ
QlGM+yacc/WsbBccjeWCYDIctiE4Kfm1gaWLreCyE0vW+O3lOnKFgGjccfdTlhHQ
3LvZ4nKYnZcjzJz/YbncAFnG3V+COqE6fIbCKGtjjHGp8K9rrnT8NW0o1GS57fC0
qY0kMRkJKLnBFGbpa1u0X6/C5ILkMCQrsgX0EyqYx3ZDsQ8PvUcJloI2MOALwGGq
zp7/cV2lYUBbHylJj5QgoVCDRh+BFquwzZCqJTVugLhmGXxkYoZTRuEe30vstwT9
4Dot6BQl9pBfKJ5wCWkjccxu9byE58cq2v26FMAXE08bUn85A8QS0vNERBP/qbjF
8ycTvHbd8zxw5ob7rVm/Z32wrx2rlm8KAS93Y7DGl/acTN+QpYN7m87LwB2jfXw9
NoT1W523kwasZiRJDS+YShWB+gT7RTwzHTGmj5d/2f7O7n5ma37RWDfDO3Fdobn4
ewzqgDPoUzVZuY/3ihuh33xn8Q1mjYFnUgSxABiGSta7ZitiohZspG3U5jtCs01/
KDsuvVV3AWqGIT/Owjc3ZORc7ZFJfEf6YjeazUAbajhV3kSVeWtDUNOrDneBsHvr
EYCf/n3eL/UYmuZJXzBmqhHbtP6qYPLnIiTRaLNPNQRzlOBqO2c/EezjbSqXovBa
9XufqJgvRahiD+uEh0uqWS2D1syRoff9Dc5fPaDRuADq2QEO+r1PCp4cCJQM6ZB3
49xuf6Yk/pMNpdYs6lziuAjzjS1PROJcgXCSvjnDomCIhop/6RAsViNMjMF4AfJn
xpZ76kTHdv2NcnHc0skbdkzjWfunqdecEwIYOkHdUk83AnubVfcxWH9XGhx3ii4T
w7CaE/vQp5oPKIGSpTtb88zRhq8HKFlgCwnsljMkwlfH7aOQqf729X73nTMPdDF5
FoOrdDhowN0kChuk5qfCb7ER+BYrrldny6GLVSGeM7MIgZJTNYiQ+BhWqh/P8WfR
by6txNK359oF5gM2LdBm1fc4jgOnoS1iZxllixkyEKabzoHGqfTbDOZZVjIye59H
rNWhXVEdcp3jITGSC/VvBTE/sJ4mKxgZwNqjxk9+U5vj2wakcjosGB87SRpajaRM
AGXVX3pL6s/wVEXduzrhoUMY0PBhf13qPEVqjjZX4F0Figy9Ek8tzG2VeX7SJLAl
592r0Wc+Nd7QgMeqMi/cj5a7o3TAH9i4LS8Dlfj93G/VMjRG4WDDkHW3Kc+vYlSg
x1t6YVMcXnNUoLcjvTJnLBwiTgZUy9HZxBbn7rK24OWfepI7r8HwSy7B0SRziUxN
wHeJzgXaE3FJ50hi7ihM+HDld7dMOZNQ9Prl4NyImeWXS3ab6wU6fsmcrsj7QdRf
LSggVhnmqvyBcE2TUsGm/vCWp+FAoazYjfUUg28HezhhgulKwyK6imq7dc74Mdt5
wFQsa/ACIefLKpLIVQBvkGVc7tVnK4Fr5S+y269inKoEibyn7Q1L3wqTC4aOIOlX
yj8WBm/XD07cT7xx5AZOLXgP+MdLl6+1Vsxy+uwvM1JWds7lhz4k6n3k9Jkn+xW3
FO1k9mRE3OvEnvXJRjApeT5dGkJqBBGfSRt2mmbmTQnfIRz9cLTsfQY/csNpY8yd
OHDSTpLm1Cjo4ZVqoUPCXWukHzG5FVlVwonBYuCrCvyt2ODtqsOzXTmKfaDkfIuI
3yhnEtUJCaQYvEzG3xXM4WCiYooLJfBMVfaFfsqV2IeaLDVmxChQ2tFJFtjbjsKI
89771WH5hL3uTgIDKDbrXo0OzM8kW6imhBsG/ryy6Gldi14yN5Iuib1JaS4/v6eY
mW+e5GlvKzaFJWuDCVhUTQcDGcOIRtrgP8kebIz4kkCP7nnsD1ky3jkTZP13xj43
6nyBb+9uVJScHiTutoC9SSGCzavCyLqGu9fw8yDjeE5wYzF2LlHuDPrSMLT21BVH
kv6HQsExlhSPZydytDKrGEgyKRdh76u2ChBaNDdQnSFLzI5D43xWy/g5N4YdQ+YS
TXeDTcKqhZBixl4gclELJqNx7q+QSGbDaDHLuaSKu7DKJLpdtd7dceMkCVhX50t0
tpsDoCtD8DsLF286JYbv6gd8Cmdd70XaxXlCXRNcY6o3dfO+owGzk95R/QIGJ1z3
YZktgFPA09Sa2v5VlB9UDgtUOecRDJUpRV627Ro54G5PSyJ+fQ+21qXrepZPq2H+
9GxNWi6h/slwXwLK3YPXtpCC4Yyz2MqqY3C6i52F4T/cWgkTRo37g3u8DEvZDq70
uhysp+IpSGaFHWc9LrnKbpg06eDcdkIxEau9AiixxosbNFM7S5E+GORdQWtxt47i
b7Gk2QMubet1uAUvoXWUq5Wmz6B4uujAXWCvReV2NUvzTWHvbDEsO6vCkNiUymPB
EQE5ehPLUBJQy+6MktpPd7NZOT4Us8cAB4Gpt+ylvuAv7hH1NJIBCkm9o9dQF/dW
X62VzitMB3Y/FjIF8qeF+WTGAHa8lNm6QoMmn8ZhinmDHSxvipkGHlRNtlxywwBJ
+DYFekOgtnsfImSVhHfsMVcU3jadYkg2/qmzUm8AhdDEdhXRtGskO2OqNe9HYaJ3
nAxnS2fqb1RJvpGNgsOR/zmHvZ70hzzywgmakw/s5Wm8bgib1AkXxyWfcM3KyB4K
osVX7HsBTcgvNPUpywinogBzjIRQNS6SoXj3yNz8VijOEiuvp7OfmHghq6x1Yx4F
Q+BfAIVuMqz1IHiq2jjrI5vDDB4Dn69Idpch6Kww/8ERCAxYN5QjBnyRUMm0xQ9p
dp4BHo1Z5/Dz4DQZgOsqDmw9ERtAzatsU7H2qrfxVwHklX7HKbbZWwrf42VRUvPF
CQz4AaQWV5byjhBx0GSWFvmKSXfF4lhmWrm6gaa2rdCPHhAATjPZFmXz7mLBIhlH
phwc4dsX76Pof+z71Q25b8VEL59B/2LGrRnc0/ycI82ktY2sg7xGc9Sux040nJ1f
j8sseJvlz2tUcsnlXnE0k0gI1jQsD1qIGZAY2WVyegpU/1qsrkqv1fOr0YK8yJgB
KoRTY2xikdrwYkpbWV4NKIoDelVszNMQFaul7Es1PLStLpAk7V7oY8AfZUmA5owS
RIFNEGV9XPTt2oFKTwsVFlw+hbGGpPpEjmJ3Hz81FC7YIZM+ssHG2x2RoIqT422y
uuSRq+DZzBjY5s1MH2jVrxTRTmMvVefdRtU667WEHwt6M9lpoC685YRBmSQlavby
9y6Brp4FdfsJKVFtdvOzruislBSX8xPSvj7z8AojKoi/EQwReE9WVxUWf9ZTSWW/
zBbkcd1I2XAa2DddzerqBrXvercZNNVvLjrjuv7aQKkedznuXw2xb2TnWF+Tov7t
I4v0Xmt6b8NWeX5c/6HTwrAtkDxSWXgK6OlZe+Pt1+W2nS6c8roX+8bofhikFiFh
8H4VJyp+ouCVyMDmE11XHgtL6fs/NpjU5pB4nQyDGQ/wUZPWHzapR8TJo7CQqtiU
wxXkh7IJSKLPQjiQ3SSAUTgDTxesriSy4dZXL9K/iGuVhU+BujM0aZLHx8IBxrRU
fSLSkkkgfdyCUaFoZ1PZQ6lKlwh5mHB0RTMnrD5vyBKKIQ2xHLCIo22nn+mZ8NYx
wbzzY4leh7SDid/74ZwxlMyWO93VxrojyMDNVvgwMhZ++0hvNuYjwytcS77GXZ1c
j3WNUG4F648hE/g3eA5T2vfbxoZ1S+Q2JznQmskwxnWSGD/xCjTj+KCUwAmELh7O
wSBDvqTQcKBcG5VC4zlgPWdttSDFW9iUzX4BSUsMXIUQqV2SLshX5ePnn+tyW3kk
jqYqnTVPlzEaP11jDIIf632H1xb+RPZBt8ZrzRGzBbDTnWp0dykK4uMO9YEV5rZe
pYsjLk8HpDZbMBnNRiiEAmUwxv0kEpU6dQ7MzJERhFuyiyc7t6LpOtSIqKoH4PSH
LbbV4+OEoj8o3C1KBSVdWdcJYAvHRSHlQLfuibpKl8tbdaZ/Sj57YHrvTGZwsEQ5
aIU0eQuXql4QpX/8EOx0A3JAO9pY2kBzPZm1aemjgR5yfkL4KfktQpOJmh39FPPG
Aw4OKr65psYYs3PNoqMDEeMA3BkAEEUyuBPIdl5OGY7tRw0+gxw6uwfKfi5jEA7M
ZM1uWHNeeVfXXa8f/dV5A49cxFp8pFjn4+Kt2XGVBrqNv9q2UQqwNGWfkIhzYOIF
Djb0/ElyQ5ecG/dz+C8oQHAjGCfleCrCI4XqzUDewMlY2LD/FTW3S9fy0j2vWTOi
b9hIswiJlkKG9WwMm00RYNEX6Ckk5VJ9uT4P2RiDGv3RBFSJkrxqNf+XigtB6/Xp
HtoYdALZg+0W4KB9I6TBU5bzGkzHBcP71RzPTSFmY6UoevvSiPJPuuROgQ5YgK9f
GBYJMESv/cIUdyWB5DhJL/veuJXX7P8fvvvmDy1lT0zDzj3XdiQmS3TfPYiUlGT6
FLT/tDE4kDfjGXaoXOPkY2jVrTLPAKOA1ky8kTFUee8hUQuA2SMSmHDvd1kDEoP8
Q+nn2x2UhHCtzj0RSs8TKXtlGI8vPa/M/hw98xzxXOK7Ztx4IIDLBkdmXItaHlbU
sVl6VCmfekM29M7sPKzQqjTqb8qG/S3Vn3jZV/w6fjG/fmTJTxp/va/c1oRqCy24
6pU2kxcewKHd3b9luRWSUgjPezjDp7V+o0nT39HubpwLg53aygXrfNeo4GDSKYku
4/+3joKf+QCUmc0ztjaHxdV4ZPzPlgtGNz9Ro6+jxkHvpS6q8lPi0Is25UotK3wa
7jJuwWC8oLIw/Op5qp7OzWUJ8UZbYg8rX2jDyb4sNggO92MOeIWCkkFOwFQQlV4q
Gsb1elnCK8FDsG/tt/h8iebsJhZ+HxEddwA4QnOF9ZGoreNsRjCvwOYB0vcW1kNI
HtifVzar2Jz3G79i/pHfwG90RyRBbAJP5zZa+FTcg561SnQEBeC8RtyrY4L0vO2i
60iWtj4tHIK5W3pgsBAKS+E5UMz9XlSoxZXIVILLOs/736N/Sm0Avv3ggNzUdcXq
WWi2yxx//m+o69WbKdV/NloAbWuroQ6CzNoOkxzPCGU9y4G/3o/+HBCZsf5h64gO
bwQvpYPfjGAB4X+87X7/qkatqMAg/gw3XZRPpsK2qR9Up3/QxNMbmyheQ7igao/l
1EYP6NNwdBdaJqFdHBKSVQQhz0qopN0Qxu7AyAzxI7rRkkBnWkc1zptyLwzG6DsJ
CzoD9TORLnCQv0p9KNz3tEeF0NCq5ItB2PuqmUwKpn6O7qeHX5Z6JKkEaMlqOBg0
rXPZsMz+DAPfmus18hzgdpVzOmenqowFK1TMCub1HONMj1jLR/QuhQyu33Z5C2Ot
Nt+QsvfAYwopiNnsu7x5MTKfQeu/vVPjBjlmH6F/5W9bqKtqE0ZdShnaGYEqDaAK
j4cTSAyO7xg2LYynpGIr+OJq2LZCcsdjHG18egwfYukrDgrZsstQ9BFmy/xs0pwT
f6RcBiqqFHUQtyUTPa2w2Ho+0CnYpPFvOrb3z7tEfbYbWj2omYIU9XHJaq4fIJYZ
7e4Eh+23DKWyWbkoQcryhXFTb3jFvVX/bTj+pPkr1IEAgabkp/iEmY2t+K1lHjKY
IOl+TfYe3XqqdlEvjvdYxyj6M1lRsiNftwfh07zPvWyjqdK6FOReOkYDtUIl8qOP
mKkabdHRcdnz24ZztfWSNf1k7XKZe6CNfQ7Sd/OAre6hzB+m56UX6GXv0FoQ7lgr
d/Bzqk32S96gTkWzOtUGU6TjbM4TkcdGglXLMxFaKJIAYLDXs34PkEeQ2prAqDCg
DRLed8zycjyH8YA9zv+6lliiicbLEZuhRv7O+LwLWKFgIEnRdEIfJ1JmOOJsUS6V
Bv13neDlp5pWfBKinL2KaAG7oujQYp4gBQ8wUZM88jnjHHErIq2w9fEsMObO6/Ml
w9jIZhNXNZksiKXarEmR0GdLW4yyu8SYAFeUf3HKEgIDyPYmflGfSVjDR7Wqms1s
kvd+S7DK0Z4rQpGHdZTqiN+se14ud8MMaTUAwaw3UgZzHAPdfDLYd2Ar6XkHrK1p
GnTromsaKeMOUTmNOoQyIt5x98gpYthHcOzlj0MPipzKIPgcDOKhkTBtxfD+vd6e
TP/I7xgN1dOrUbgkH4AcbHcnF+9lItM3u51d+DqTEHYUK4QinbVASLSyMrCAIAe4
mlx9aFrzxaxbHPfv9vD1b4wl4nBFqeMPmM3FN+C/tVL+76Zp2klQyYs5yyrtjJjJ
4lhA1W/R4YPr2QnfsaTVXtF1kVspJXMxC7rihq7d6G0VqoN1T1xLieKMNWiMtUmD
uXP5gicDKqqxDbj2OhAJojtlh+w+yWxYhkWGTxkaQamVQk0nMbKKCPDZLbrx16EG
VHdZLUUbBopGvM/2IkLTG9FtQbB/Bkw/LHe7VWQ08m3+lTp/6zO1OulVObxb7VOA
OZz6gbdqmvdQivPEaMIXMuv4OIiavPSodbfvUOWkQMTRM3iWVog3/iCbUNlA2ppW
pBd6q9v0zKatfLWaTfmRMiPnF/pKA5i6UpBIl9epuVYbJX2Y0wXFU9LUSXgKaBY/
ZvjrAWvzXyQVvshlL0BxcPfFr/hayd/EQ79AcIO/spvWk7T6SREu5+fZrrTFGwqV
fERybs2rWS0aoedSCsH2eZg68F+NaESVdwf14Eu1PrUQk/UiFyLKvVaLx56kuwWV
KIzaiTdsU19mX/7Lz9syYArMsJuAUQTIrpwUvvQwG6igggNjspHEvxDQU8gmHFNj
FGaNWYPd2zRjdNS0uirIIcLjR7rZ4U8GLBTU7RxQY+mP9Fg0LehVfqzytWCtR+Im
zasVrcpcIhf2CAuGTj6iTIxZrxY2k6sYKDTU40Sx7xmOdMSf3e6/NGfzFQqdDH/8
dRfWRG9/cPMAyG3lG71kMM4syuSj7DhlfoLHCAHW7XImDTdgJEqDpei7rbLqPCc5
Qd4A4RaqRlhxOLifR77X2L9R4GyihY3TiE3f3EAwhbs/6yM+AhufS95h+CJz9TFG
EPTPBYrFhDnLWCO113hquPLNdtlQVPtbjAmyRyKBqgg6lMNyLNCs7qkmMOazG16y
N18sz8pNMcRAV/w+jIgSZU48PQ0tCv81RZ7bjB2oMW/O/jqF6hqb8v1tFI9w2xDd
hcNj14Klrx9iyYnkii1zt9tFWlue+RPz8AJAFvTrc50E2/p8cxRbjuPs0izXxmf8
54PHhNj9qg6DVlkBVOgOkOtuV401TDb4CUfAodn0CCsGEwOVpcBLpvAO9SF4/R6J
JC1UIRwGuB5sSUmDVUjGAyYRT1GizEe8xtYHkvwFSZl02rlTX+URVD3xm/UsubZB
mH/4GHirYPSM37MyaHXf3RQtbZQEj0IKo9aVEchAIdx2VWT6mv1TrgFD8PlToB6b
FX0VR8kEhfIzdCpd59oONbcmJDeCtTCfzP2nyZcKqFG6DA0TV2GmGZJhiIrQxkOp
Y6nFeZ+X5r6nAWEJBJIWF/BPzUcVAbKnblHJ+QYa6XVCnrd6qvdzI9ihusmPobq7
8rJnuDoiqwHTRrlrfldzuElKjeQuq9eGniiDJZ4sCB4psZgoQfi/rzC3k+BYjbYY
ltDn3bx+vGoyWESA4da2aLODTK9oXkRuv965DMs6yAGcS9WSoabAILgwIzYiQNpK
1m1nvIk1aJ1faU4ozwzqwUDdBpBgjCbgoDGdXdOPn0MbJ6YYXkZpGNF7HbuOlXj/
woAXbEqxn2BnC+K09XN+9vsUqGkYnSawvtTuoYYqcvM4Ag/K1A4zVSdPQDwWb6dM
hkhICfhrOuuYuP1jgg9DBasIzrdERDm8m/OCWDfU238f2eHVngMv4X4/v8iGRym9
USexQXxqkmnS7S7bTA+wlkzctqXV6ZVSPXTVWjpjoX2ttz0wX1+zc0VbSNH3Nl0k
YJbpZtjD6qedePjc4XA6gc2FzfFyMYn3Oyh3SBGceKm05x4n5ycdHQZJwe6SQKrX
ihi2vgJ1GGWnnBvdLstlxED532RRXROJsiCERsE4LAC0hjXzeL7VV/OmjThl3pfk
vUyK2ZmukEUoMTdjGvT4ctW/XXrSTbIxWsGuSeRrM6u5K82HjJNLfmXdnU+xzygy
2nCznHZXgij7qScbXDnRvVtj/lxHgx6NZbKo7VN5XSNtNm1HEB7/jeztCb7ATRfY
UtyqXkWkPSVBnVlF+GP43DXsSU8ry0cioJpAR3BgnO4FRJOpJYIjd6QanfXlD+/L
OlEERlyCAseb5p5+ZKAl4bSlJVEipzvcnsngmdzOYOkK0VP1h5VI/wI/oGNDURcO
sGQdVc4GgW06M06+zimHHYq3w+NIOPMT5IaSMwxpdfGtP34UcPTvaHMaUdQfRf7W
Zi41yA467BX6jOeexWjc9LbLnpf2hbrzQQuAjabC3gTBz9xu4TBguLgHITGB5XBY
g8rH8YZDWQSR0CC0EFHFLAMmcRG0MO1DiOHA5Arw+h3hZ8Ryd8CoCfL2frtb5UXD
ZRzCv0D6sqBZOxXtlFLTifPbhnBnBHGM7tmw6iSRsdiz3KW7PA7AXpoD0uzIhlQ5
nCKxmcoWYzts47IHHVA82djqWtJvlZfYIf50x7vMG+Ljn3w0DSJxebbxxyEhvSaQ
zwUHoOV9NZXGVa9B7VbGZQiOIYjN+oesHfpK+NQck4B/osHqciyQlDw+/Tylh1L/
sE0xy3eSH1yhbHHvHw/qzyRt+vkK2kpjhrJCu+7AXBa2ioBITz1Ij6aXIbuGf9uE
v48V8q29HM7fuGERJ7ovQ/ZGYGRPaS4fUU/uj0Oemgn2cyAFhbMXCIir/E7g62Nk
1DBNg8AJqK7ZQfPjRhREVhABpzvMuhtNq5vkTNQK40HMaPoGs3L9FdIgQzthayEN
3ui/kFN3gAbmr1eq6Fl+6m4eCd6kH8fP0x14FliRO5mCngz67bewrsfK/AnkJA5c
+nh2p6/NEye04lG7oHZGB2sagSytGXeLXAhbMQy3yQGrZJPVGNv7OzEMJ6AnKtyB
WXfthM9mBzJIkz3keLPGByiDs2tJdzkf8saLsp/5y9uG/nDHRwuex6017LG7ho9m
wO4glY38T9+wOESRkakIMH8R9ZPvcabqRdB1ZEbNMSqWQ6hj5Inq+0KqGQFBsedi
KVly9g5oJVTlEqo0yuUGHZeqGeRlZCm9A4mQ+p7oNFlhLeEA1NYCtmErA5PW1zLO
FUiHgcOaFV8Tn2ZBq1MzEbs7vJENKi4uti3x77Xyy1KtndNwkKJPw4phDXVMawSY
20vNapVrudFrY3i0/KRZRko8g35gOsqCYmOzCrjTdgyot/Qtv7rCu03lZZbvrIAP
rqPAGvz/xJrnFxzM1/eyKkBbtUhEoisMRp5Ya9aFogmlvLxxa44L6OMn4BR+gPji
cUmPlItrwkj/KgPdr4yEwy2gDK27Ba2MxFSVvJnwUBkXf78jVbIfeIkGBdg8YnG9
pIFjN0UYnatCybGIQEx9XvEfJgPmGYjdYFomDFYXctuJxPcfvc9ly4/S/ljFoadB
Emxr/ylNWCTRfjXuJtb4PhM6xR+3Ytj1Z6u1Djec0CAAZP9wgoULbRvFoP86893u
KWDvow7uCni4RjFIEcrO2QEs+cfVDnJo/HES1O+T8sR0UHG5qF5gOtPGRk2ZrEUY
DbL1V3zp9xREQ6MdjqNEEjOFnvGmX55o2+SN2Yb3XlltnJNFDchXY5iWn/iM/55y
qrJr1FCyqeKZHyj+2wnuNKPkM7GrHgSoYU3yA4AYAgJxUUuogxf5TLrm4k5qJuuv
b0TFORD9v0QHomZOlZtG6qhHQcHNvJwS53cL9eH6c2nOJh6KiZcx1zTxE9ikXITE
ycIR/MNWUoN6YnNr3lKL2XU20paVsIpg13/CBq6NHy+PiRyYriQkjmba010XAAKB
9TLAmVFo9RAAY+XHhsCe+SPuathBmO6lxUM7jhaHnpIxykqKVvVjb8l8kWFx3BWG
flG33VaI+XEyyIonM37wM1ewXKcyM0YYN/pXw3Rtb6eb5X+RBI5eEFAoPHcjz6M+
H/iGbUVa/OAcfE3olEwCKrWefUgTTITb/1wKu3+Rq4UcFY/Gwk1lsGnpDeCQb/O0
nEIfrlNEe944//zMqjJxjc1TdWrb5fYN8J/0GJqBiONMATNaLqfCoCVXLDxwOQYa
7daEH1pdI2gIO1YPpY/+8KBKUpG33NipGFFTpH9Iee5A/J3S+7s+hYBZjH97LryQ
C0x3dBthU/JT068dDb/llTfvahcCgL3AtRDJKpiIkFiJ0KgtRHlKpkesS2UkvCb1
x8+RzX8moRuDU66EuAXjQGGQe267jAvB5S4Cjl+QE1vDt09ZjoEaF/4TESNPS/Su
JFjIgURKC2ve7LeYSBC/XpTlkhYtYcCUPObm8/D70ddLhn+ra1zyACjKp04rZOIE
MnSy4RAsSkavjKGE8vQlH6Wdr8z+hCzpa0nskH4pqMCqItoxuQBQC3jVChj2SXU9
Vwy9E1ynqj5Gbjm5cG/22ecS8pVasPCF3k7l5SxsMeARaZ5+e9PIGU5EUrna0+am
r3pceTQ2YBb9YmmTOQaCO4FoiCzMcbDIxDtI28WNF1L4c72eqdmxxalK/HwlOGJ7
HXkLMIJ8DjH/CSW5SqOm2B1oWF/6RHIajoKShG34iXL5lW6NMcNYP0dU8bhu4ZGw
RCvVNrx9c0dxFBLj6tR8Htev3UA9DDOHvsUEMg2GX5hUYLvqx8OJhHFXK449JPYX
A2iDDAcvikx9YHil3fFlr9kAGLcWdbYTB2b3cpbHyEJNOM7hbe2O34phUFU8tkQz
9b4v0PfllbRwe7R2EuOZQcAzWNMSYlDzqPG7BOYnKEDTW51PxoAE1+7mluE+J20Z
mKAfhG1DEyTgDN+5sSi61uZSYqMmRRtcnyj/lYBhN+FLi3CAtCVSjCqV/8ox4vhN
10MvaRkWdDLIFFcflEBtv4Ckw7Cl6BjkxxPL29gmc2Kkd7uju0KlTMk+mZu2ilN4
VoN91q7Xv0zyI7iLoZaNwDt56TtafAFQy+tBtFxQPEjN6ZaiPFMHdh7fSvpNIHp6
zss3QLUuTrU59u3V7Xiwsy+a1zhvVyqWDxUEygfwRPpBvfhZxNs+nEAP7XI2UrR3
J4zmwrKq3lo6FGqrCIlZOAwgogSRQpN/vKrdvr42wc485M8k+BjUfaP3O3sEU4eQ
hwJasyGrzC5vZSAEJMM247jphSSkbM3unX8uQqVklYS/u4qOP4t/e1jPgfvoJXob
mkgwWCV+FRo7LbUzpNU9bDhYcMzX4eoC3Gp+wrxDIWt0zHvwlHBNj7gmfxqqDDbv
7AqOCxZ24miAyeQrXFOKssYXSc1VX0xDJbYR5zmfSIVLwGg1wKqOXDXBs5twBdM9
cVwQAYOQ0FC52KugAIKquRw5xQ+bl6IQYqQLqmqDA4xGHWzUTZyunljpZfff9Kkc
UlqWJg4BlOO2nNalW9VYaMpvGF84jGN7uisgaCKzS3SZBOmkWeKCJyjKH0UqNtFq
H4rItdS2rr67EpW09gfB0ZMPaMC0uWRK08h/Qv/dHwdVSmIylWe/rwXyDub4otaG
/drAL0DKryMV0trX7Sz2NMPbiefI9IX7GzttLLCA5qLiVsoy3Oe3kNMebCOPox9o
MYiXmlWCtD1XleAbW4VF/fpUJiroLqOVaQLOQu8jKm+UWAYL4k5L8OgVJ4H4y2C9
gP8zITtu+UkX0XgxzPcnZMyqG8jwQIdKvHGc+/D3JpBaIANN6eOOtPBHxEk8ZaYw
bQ9pvYg3mg5ZTzEB8tx/uTg+rJ/37U1HwsJG3uzYoQwxdx2AdJl5bEzgZrWiepLn
B+Rh1TFqpIgpyf6q7wS242Fs5N6v92u7lmiURoAtKZ8SiXeQFjEJKwj/5NAjZQKQ
1LJZERGXOiPFfFUOYqjzvBsWcim0DnA15XSPmvDI/ehyUm59TBTjVvX/p9hDgCSV
KQ0d6wrSSSDYBSHCDyQDSE3QueumN0w0O/Rj2fO28ZEO9+FqHH5TH1CpBxYlz7sf
ut/rFliAr13wM2tWB9MdI/C1+XFUe0ZnaDwlsORI9gghVUk/xAvuBDGxpIPwl1cX
Olib8EuS5x3+F6A1loY2yt/WHQwC1kF9/Ho61CNMhjFWsVVumZJpAPzir82QeRC5
qpfXW086kh1Tr92nX4XpmaVGOfDWL25Rl0rMNTDU/Lb+6ndiF5r2NTnC1BqRQLRW
3y/bM5uRUUsav0s2GnLAk/twbQSOcaPrPND4Pi2na8spLIxyxX7LDPA+MwOiTiF2
C+vll6sF2DVq2RaYZu5xwSDJzMgWYXNGRjfElAV0W8sIQcHw6oPZyTnn2HDMmoYb
w0Pm64AlL5UhzztTEZiM2uWivCl2utMrVw/2wSQrT3wh3Cl78gjd5G/T1NqOTHMg
tBWOlHEpLO3d3GIYuUlRM6h2MqAkIoBimqYYV9Dg4hPV/NaaBwioGssGvqOkCJ2l
uOxIp/44z3Xuf/v8VCxBSlOUi/PmesMNiGgHBNa8jVSsmH0SuXqHRH7TvhZQSu+6
hbJCoX9Gw/3GGQgswEPG5YV0xkLYj9vTpj0UR53Dk5RhZWb4ltCf8s0Qpy7UauK6
mAUBI2p6wUTJZdB72b35RFOMZljLoex9bfAK7IWzOUfi8a9g+gX1ffkVQ4FgPDd3
HQOIltk0cQHvkSb1QTaAIn1rOBSefXqCyr8DVLEs4SC3dpqcBA0NwKXPjl6M4edz
cxQbPGIYeua8LCGeKK7tmgRiI8/3kqKetCRwT33uteuBKhoF/ZPcZ1F0Mr3Y1tCt
NdnqzJujWZNCEKzQhOona1kekSkM4Cn8gScvNDEUwGjyjHQ5+15i17ucIptWCeNT
BhIKq2f0YESVIFHav8+L8sWyrRYy32uqfDxbUiHilysaipZmuMs+KzQWGTOXvAa7
j0YhiiZvEk2/8HmKGh2polq4nToQodyfWuo6cdsLZdiydzbUJXdNuKvIYXkptdJQ
62KoOh3/Hxx0nxVwMIvcfoAkD5vn+hGrfpE2ugCb3+3UBOGsCzEYi3jnNTnfaqVa
xHDwlz5bGqv0hmd0X6Tgk5swua4+8MjVYHva/z5KFnDiP6hCJer44euVtgs0tN1z
zVWl2KNjTcpvZLjwTTAb3A9sNxu/xJX2kiobXWg8npaAODaSiYERpI8HXkPzvqL7
TyO4sLiknG4OrISpFl8BQt6p+maTaxEtEHe7OJ3KJwkfIiRXyFd/ILFt+1ZtCgDD
FSoJOqGtI0UtmszsHW17PAG4MyEjSvRb09BN2oe9a0a45tDEydvQ7oJvFxKQG1w2
XoPUVNecPxUjYOsOeNSTnEwU3wOIwletSe4krwr/0LK1LWNO04/ejDlD7WCkB4s+
5XfIaBUXVMBf3/MwQNlXIjXtI4MuUCDe8YJZDAwZmBdL27oIty78UQtmSb8CwoV/
sbtJa1nA73j6+DhuTDcEvozfWWi6ipFuf4wf64+B1LyweP0ENlPfeS3ImAv89NYT
9aprZV3gpLLwcDbb1E2+OjBOEPSxGWQ4j0PZIAS34Jz12iMUgmMvMN2xsAQ0PNIA
AjAU1jHgoe2dypppW5Us9BEM6IrvuHRqm+zhw0GhnHBTj5DkM6q0h/AuQVpravuH
YZwVHuOtJafm+l5LXUVKivyNzB66Y0gypB5KBTeIBt4R3kv7EV3QXz9TJpc1MChA
8MM915+RXP4FGlArarTcBqgiM4tW+NjpPmRrSarciFqU0g8SzBq69snKvljj2M4N
hTrg70QI18P2LBmHCuXqVRtgMicgCya/gOWsRAC5BNmEW+7SivHBDgroo7AzfwLn
j+4EJDGl62rfyIDyUQ7QoG+OUTY5ZoQon2Y8aOvdzhtUxWYWISxONF8jfbTzZFo7
TLAyTXlgesOGLHeku5j5ulCbNyPJ+Lqp1pKvMfdeiFllNzL24So3QXk0Dsi9FvI9
IHKnxJMGEackfQShxerCJWz86NaAuH8LDas7uFDrd9rGCJNU5LUHk5QKpr+O9UZz
JlYiZD3+1Uu8m7myfXbf1vJ3Llwd0ZgCtwoM+TjakDrR3r5//kfp+4uNyikN/Gj+
XXrVd8mcQ3uMrWb9YCA91WlKsrkiLcrdwGqNQdCnhJiEVwgNbz2Xvbu3fsPlwuCp
QjuUCgzsrs6BMD/Q6kml1WzuO23TbvehxXFMXtlisSJOyH26IzpniuesTf8HVUI/
/y/MOIoZjXMdzu/xIfS1JUUYQZdgWUd94h1Jh3dGcS2Ls5PbvAIATXPPVVR/kkNx
4QsK0rclEPbvccXkRryTI/Rp3tStwyBqYiRDo/Jw7pi2r12W5H4b3LKmWy8HxWhO
LnIh9izbInb0pEmpAo57rJGUu3X5CIdU3vk6WcwQh7G+v8mG3RD3CquKJiheZBZu
jFJVLBqXvLNGq3E1dlAqvbf64YK7w4Q0v6Fz0BgPejHcWNJEE0FefVgv+WnRX6n3
d/UAn+Rgx47hCUnmh6eeD3iEl1lkh2QarEW3dLgoRPo8m7pR0NdjFEPdNZwMM8DE
l+7C09+aQwazeFDQGG8ZQFDSfZU62VPEtDnkLd8ucXkbzRAJU8PevE5rVPZ7WSZL
IJWPn734oCpW7RiO2TYsCm0NPwThxNoI0fd06E7Nao3OvRYQ0cBWsY3j4hv9Dsod
4uad0sSRLie7pD0VN6X1NkhGV/s2+W2NVZRhqJvwe5u1TicxLgwqSELUILlUVvw5
Ao+cliW7CZK+A2vkQ5wRJTOdKRS10Qmb8pFfOh5HC2F+ah/tJnie5xIdphdzBH/D
QlAV9UdDODr4jb2uTcFkDg1PPaaHPBYxe7GezK/JS09lGLOKGZ57kiSq2hnctbxN
SBkyvnucUHHYtNyagowjsZz8gFB+smhpXOkZSwrPM/1vyxm6/f2DfhT09P1vnOGc
65vHEDQkYTctoe0dxtYN8i/daceCHXKOQ96L2Z1CLIKzh0HWrB6PFRnshv69aakc
WvGPb4KioBcVMz1tVRQpZfQrQG/ZrFb4o+UD9O6Wc3kLMhs1CXq+IHbfz/JaBBX9
vIjq4DJ1u4EQ0nx8qi/VgpUTL2x6DakU6lwqKXKfcAUxIVCpA8rRvIizr5r8NZXK
pjHG4IQlJEWvQE30s6EjR9cixYejB8iw8hcnaxIEqwp21cRB1pU4wTJhheVGMCu7
AKKL19Wu7n+cnulwldu9xv79h9/bFRTc86bnatN6hd28FjRyUKcU4oJse+5q3H9k
7w/Cx+OwTXyxEOg6e8kgyhGeVwTqHlPiEZMTtQ3/9EEubJ4RRVivF19p7sW5s+qn
+8sZL7Ow8/NV8YD6QU5yGMBy51DOAyYTKozCfYPpYZbjR1jDhWIMRNd9Fhy6olnO
J3VF2O/GduIjAtwZ27gUFIWcelcMhBciJ/8bSI317sOSzEGkCPhu5m8EyXQFLhHh
g+tA3+J0IQXv+0yN6Au/A1xr8ZaJaTLP33LPRj0prttl2LNV682WhdV4hkpqKGNf
U+UzRPbo34EUSil+jWjdx/aDnzzeBZqj/O/uoWzPX8r97fFS37QSCpVrZjykVgpj
Q6tfgbqGo7vTGWdB7M8A0yHY557c8Osh40jmY3HLKoVuAhsX+vgeNjnkO8Tdcdzc
mIdggIWawUg5i+HWMpap3O2QIxzGB3NoHkTeAX0cZiXxSBHSGvNcxS4iXAXmdf9B
ZdwJIXVKyWDyWV1d6eVo2cF/2+rNZ4JuvkFw5Thfa13osVQpaM7nxNZ13jBseYFy
ILrcL5mdG7bEs4wvDmpG/sVO2GiUqocRuj2+lhA204WgBJ/452S2Uj31Km866Fl8
25FGYaEbOXky8nW8hflCk57wOUK/Mnr13IJuzY5F+hkOX2IP5aRHGnPGgkiSuLFM
C42uIL2dhriA8YK0Z78by2u/2cQoFrEDcY1elpWhpDE2vCDkAbrWrlBcRGL7FCN6
wLeqAlg5X7VXaeTdQBjx4j29qimmxEQI1sWKjlb5xfD/jjbaSjQg3daxHgO3CWdz
vSbSIqROzqGfDPtriFF+dg4joao02gFh2Cli1po/rYEKxtJoSLYCcrHeADYmeiSQ
AW167l+UZ9hQCu1/EaqvHQ6ev5fTv3uVeQeHeSE6u6Mrg9Vw9pboh0yzdisgHuly
Avw5vDDyCzRHoVmenDFC3WETUZ9x6B5J5Hrw/0jh6Y9VGktKsOt1fQ5GCJ/J/I1z
rDeWoPhyAgy+F8Avn/13ybsaPR1yOLU+RPy2k9xMgbDrZ44zXzkGVmnyJqDgNJBn
ffRJMmO+ffqsoq/zQ77tRwb7mx290gaT9lPRQR8RLGoCjsRG4obxybogo+DwcNeH
JyeX2+DL1iAnyzVB822if0iU17fYRtLDrhpdqUjVjIIX7qIrZwmHSJ5CuBWu2WVw
AuYbQZat/MuNP3shjUkvS5ZqCrYm1ZhD3xdq+eYwbocbZ908ytxCO9R+ijlwP+SK
e+PhMd4KrWqeILjlYHEH4yZVBEXNmMYwHfqa4LUIKU26zUg8Ey7oap9o2mJ++5ch
wLVxaY+5kKdI98qO2AYYScxzvS7LXxqbAjXECYSB4YHwX0mxBfGtI8UaiaDhXGjq
jgtzp2t6Y6cFf0t09/UBruGR58MCG3CUx4OB9idB5ftVjBIf4BbyPFCGZZl7dMJv
jFBdXtPPBJ2jTc/1GybY1e0N8tCauE6AOa3a39xohcVLnRcg2pKAavITZAOt/1kK
MDomly9ZpjP7/m/3QSUvU7lLmBY88fAbtUicsKiT2MAaV3jy7IFG4iUe2CQrLo7z
0YF4UqyD9r0YPvTN1Fd4seR70ero7qP82UMBKFI7mBGHeJ9ND2mugI/2PS9UZ6aY
iGtGACJANDia9txTek3M2cb+0V3If4S7aJCf/bROG5+vXM+YRlDJXxPKTgtYSLCf
AvC6jbYf6JV9NgcdT4KykAh8FIlp6JPxhH3ijPtxuMdcYeuaDdqye6guIk1PLTOv
XEMykLD7YqOA+zEzz4umnvIuPHtpRRALjmGHwJg5LTf6tuLvAAnOa1FleWas8Ck8
iapMIgiwUveJLZ11Nh0Oy1TjfXyTmR0T1zEG6srtV3/TvnWO1rvOpn3PnN5fWFfC
qa9PKvkzINNmHUoVK0Fi1LvX8/TXotyQ8Uj7/RnWoL53luSM0MimUxFTuD4RZAIq
BB7mJb7uQTnX5eYJ7s3Fkyn1YFVnxamZ8OEiywq/lkUkvZkl6YjrmJdEA/sKEXvU
iZKkJNHoZXVNQFegU2aCZ5nsDTVY2xGR4D+TSqKW9ifPV6SSwsSv2Vvr2Plcoy+c
Zaj+1+ZDkyr0t7Dh7I50zLLfekvJThxhsVexRay85HUMb/aei5eISbUZEugKCFET
IDfhhjTmGny0dwOMie89PEG3BpALVa+myX2sUQp39A7yL3FgqfZTSlngMyzAsUf5
nczHZCxjY1lSEE15DZlPeDlI76aIZdVUAwR5kQ9xHzMzPXQkBNT5OUWq9JI7qOKb
9I3C+T/M+QHse6senYfwkQyl1RmUUeVW1N6aLunBsJIrpiU3bFv+gUQhKg5F6zu1
5ca78Pc57dn12ojcHV3dE6jtYs6XtAMXh0+RyVx+9HyDJUp/x1wShEV6NSBEE7RN
SUb77CfF7ej9+vpN0pTxhX+Uw40CXdKhfuguISINSud5vuu2JZZSHzqWx0kh65Eo
zuPHo9aL/2WvwAnjameJMzU1VO/N2h8qrqLPKhJKGr0j6JX6yKXA0zotHqPomahk
E8QC9oZakV8lN5YlkbTr3crgt8OM61RLI3ge+BREUV/cV1iXcHavezMDUfbzsWUU
+ko/erz9L0Tx6Kyse+BAFF073wFqXzV74XtOIFMFL6b6YLOpbO6SGB1+MUVqCi6u
rAEG++zP3jdCzgx9H6F44D2UCJAMASjZ0i0oyX+B2KRHQ4Lg2MCHWWNmcN19C7Zn
R81Xrc6AYIY3ipOUpAZAy+naQwnTBMm9nPpk2bsk/BCLlF8EAZCS6BNH/42kin6e
FkaeV39V3m840Mlr9BQBhZScNaIt0p+3u4CSLAPu5TdDl/acbathDWwTOZKq+S8C
joyDJERNiw+u7QhA4jT4w6Veeq+Fcg9aJx8IwUySxyZvJtq8CrsgwWlzh0mk9Tma
D08L4VxIuLdXnTNLjWXw2WHNPRaAgBAV8pEFu/3wUYtPSSr2S82cMasSis/QJ0Me
mIL7GR32Y9ynDPKC5eUrHbK5KqR3Ix06Bf+6uxV5QkhYRAzacrVCuvuRUdhJgXlG
WF4lrsjL/8Rnk2Vt2Ys0HlobB7bKG+VThxDsqHBUjQq0AA+d1DLIL7GpCy6BMefV
YT732m/3lOsK+PfsUjzk5WIp7QXrmPVlc0b5hpI9Gi30hdtbLp0vLuvv4EvRHItc
G/gQG8PVnJL+OA+qy8v+vzhsy/w2NAY4Dd55D5QZ6AgT1RWoLm34y+WY1BLQwCxb
grCCfuf8zvNEMdnq1amdKbsOcjutCU3oRYTz4w1Bv/ceyJwveHXc20WA9VXFiUod
58P7vCpV7DsyD53NAE3qA1Fz+ANnCsOh63dU8IpCTpYv/b4PSEbQMZWOZmjiVqj8
XvfCVhRlue5keICP0k2rcwcQT8sU27shF5roxnNiMeLweTmm2olwNbnG/5BfC/uG
GZMdlF1nSh5CeqllMyaxVxqAgxGaKnl/HH5RMCkHfbap59u/39GF8lIhQewQhG5b
WMkSrKRGu/amX1RgEXuKRKl7cE1GXLgPw7Ac/RhmAMDYUfq6zMnJQboRauzQeGNx
pIfbqPugaNIjGgxp/tIex5K3ct9gBEeNmltj9pr1l9eI0t4SjiLP/MahPsm5H2AH
MUtC7Pc5NVk5l6L7l1OZKiI0Dws0jX9Yr4tuPpFj7toJoxH4MgZ1PCGYsgO/1dhq
uCVPVqi8x2Pj4HuD70AD0u+pgLVDfRDEF25yuPj3a86aLLbMQassHuc6DSSbe9wQ
2IMo0HClD++HjCeNx1A1BADMsqVHSBJGpQDjTcajlpUdc8h8k+OA6gCeGCnHn8vc
`protect END_PROTECTED
