`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2+Zep4ZogCeOMXEcJeeT/gJxBFTXsLrXs5j1JPNfHkU3DS26tGWpRdmJTck/CJX
8nF06i/0013dk8OZBUHfccLKbkrq0drhclumlOF5Z94X8zqfRTZdbjAJ0nqiv5Qe
JvE+7Kizc7SKH2Q6G1sNrP0jhUdWYwbFBP8uZUdpcZx6Ws2LglKdq3qZUVt052wM
sdWgnJc9zgd1AMdriIgomO2XdTdW8voldoFxL98IGKJp3Sm5eNhlWVwLVXyPcsuP
PBAvT/z78JQ3oUwl4uAqyrtLKQP0/rftFO4C6FKP7wYAklKgXGlyNRmwl+cCCLsh
u8XeIukjb0G+y2cY8hM98k4exruM8yp2sVvtA/jozY6YjwAT+zJL9e6Q3hsHDCzl
aRbR20baZVBt2YMct9ZclDjkY9q7YFPPE6zH55Byfzicr7lyRqPinYZpgocVonKy
RNjgszytIz4uajdACRTKPpwrtyxoSeOn55DrXgrOZwlfaNRfpAncvy2bL9XDMFVr
FIfHpWQu1T9mc5+bdo8mnJbEZZWWlt2YpCJsjSDiMeySp4gcyf4X7TkuUfs/pIfO
Gk/qolt11UntN7ZccqHJRf/oFMCrIwfmMwI2YA/KH2HPhWWgdrfappdurA+15lKT
KkzBNYW5USvUNkKYJyx+XtQ9hBQ+ivTRUxQhP832LuY97gcjGeMQK47NznjYZO+z
tSQ/7XKrZeTnsmhIrWW9oOWsiUZCPhOWGw4QGWHnrgGWWLYG8wzXiVw3x+TYiUa7
A//jFp7yIHwXx0wi+39PQpnW2fdkfbxeU0aThmWErV7AHunQFqzVSARCdFSiIoy/
F0VAYbpqfDygijKJ8MbvSqAV8uNvds1+awT/Zmk37yl0+o+Khz7/JnhwrtjbQoD0
9ez98OZjLFTEExhOofEq7dfnHKc9EG3rHMcGeVEEmcf7emoBgnbfOLOaA1xwa3c7
5fJbHf3Xf6sk1CW7JrS8lSKhz4K4oKtt4VYsM3/pcmhXSwioZwqusRAhSEnKWUl+
bjM/w627sSIWTq5K/C6Q0QPa3TuNcShMGQANqvo2vYEgMEjuXeoyoL5HXAPwzQ6a
7Lsn9AaexdtkKwfjJKMr1P1beKA1pT4rA7EYzl8ZYEt2X3o9YGawKa1366wF1JK4
TszsIuvqn00svCHAp63SJjjwx7sgyM9J60sELwrv+pldRWu/ZVtGiInVTMElYPM3
ZeedhPEvcyN3a7Tpgrze+kl/FM2XjX4T4v2bVmXxRfEItGpJdt+mT9UPz468YN8G
bVQT89NECddrT/Wog/OqW43e08hziJu/pJrGKBoaDJJSgABog4RhZsm5m+XyDNxD
rxjN18MWOHZenmS35p4RsbV3OWuEL3Ui+/1DaZo1jDCmIqZna+PV0msYmv4Ovohe
vMi5Plp7S57GYmVdzO4v0XTeJFOtKg1AzoIx7DbucP8kezDTZnmsIjb9zzSNoc/W
dYeYY2C7k6PvcJt7PVXs1stH67sJmU0JBWo9+aKXaMja4cSNcvQkWzdtIVUvCrEW
l3q+NE0PxnYsX5TbiaNbUwLUgDqlRetlAqEZRhGbTwL0URVL+9kvhNqGGNw7ro9q
cDIxGpjVB5Upn9x5bYhGvx2VhtU9Z/FXY6Sj3H7r6XO4rLL951+gJZBSGDdnEaxo
FHsVKA1mgWrwBvT6tVz5yYGB5T6JzdcYI6ggwfg7Ir73fFWZ96F7pfDWo1cmMaNL
13GnRCVPshr8JgZuy/DtMkoW3UonhK4M2W8FYTkCPUV4Ew/Tg6GRx/OVOIBIiFIe
k1iV/EAK3G+fjRZz+VZdw4LCbvCQMWV89QpgE41mJ0qH8yHlyUXKRph1U1i6+/VI
4okIg0B6JJqo/PRQc8XCcEH2ccHhOqdUBiftLfekJyjXT/j3zPo5ypXLZueM/qnT
kmORXy6AYRlMb0eATiI4gRTcd28zQQbKrPkvURNB7UvkSBBPuucUs+NPT7jYf9jO
OsPXY26+FuIgP0KLR/Q3hCh8SJ9OYwazZSGk4j2ZgotplCldulC0oAw2eXS0d205
qj6Bo5p5w0CIixvUlKkiDt/xT8/PlSbv1LPYfEhLmQjaa1YZX1hGnZG86gi4ZPxH
NRmM7pGlj2btQi5hEmrbFSTv7X1tzXoQ3CpzEZRQL5I+cCt/EPaMUImp4inHb/AM
i4SuYnYIL/9fi13lkGVB0XaX5nigevgKAn4ERIE7lE5M83XbpOorzNCksMAr6/T8
PTPJMTzVQOQx7GXnfTZyLCWcJg8z2Xm7mUv0Ltkx+oDwffRuW9k0wRBeskwTOczH
8aLd6nNBIgGCX2xamfMumf/T+RRrQs60epICtvf2OG3JYgVhdBgy1LsAAFW1shKk
YlpIcSYlNfPe28s0W9UKT7msR9kEDowhxCr269dSHz8caAKAIdRStOvC25VnR9Tv
g14PhkoQE9iLRWJZWhUx0dZAS0UK0BWsWzP2QIKxILC+zrqtBT/OCEBejtHpkglQ
3ISSJQXzPq7uqCWyVDhUmyQmuFYzhKeaYYE2eqJDvHRnb5vcg01IQihuSUggJKle
f9X3PEFNzWB3b0a5U0iqBBFvXmyoUHLnwo34FLAQPpwiaTfMfBDNiP/sJJ7juQa5
`protect END_PROTECTED
