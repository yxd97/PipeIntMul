`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VlCWh/bkpMQ2fO/IUoy0h4tarjVNkAQLMSP4QHuGpWQUS/bNfM/GfQaFYZt6jFPW
CainBeiyL1NvX69HRhMxQZWlov7R7caf6Xt4wRIBTR7cQLY1XCrXX04tWgOWeYxC
217zWE6euMaZ2t8aNF2WVWf9UdIXYNLj4hL4OTwjFc1GDBtzLIWRviVypPoPvMl8
PtQ2NxmTvqsaOEaPIshissPgBGtMjFrwV/lJ4PEp5SG6vG4GaOpIHrE0uKnZuDxG
1TGxYIpwvX/lOCm9WX/XbhhR/+aiiqWFTHnhmi2ap7ubAebYL18c6e9Sk074IkY3
Wey8tAb5kWqu3fa4y0AHOH7V2FK7cmE1iSGOfCt4Yzs2EPdZlYY/2QDxnK7KgLS0
t8VXZvcCzbKgkcUbkwCpKewrwfpHpk6vm42CQD2lK4kDRL+z0GjjukhQGB1AWXqx
DjzvyMghBcAOTAO2lOgpTL7UCZQVZkY3NUFblIsGWzIeV6BXCmwE1LDrO0zH/ppa
BeHgVONYEwsbuTgkwDcEA5yjYtB7qD6BiET05T1BDYky1AdiM/fnFroYuOgggzsR
PTgUZdJb7BLikhiwPwIpoBR504vLtGYcTnY/+vcMgpP2r01VyfIVrg+bDamSKATp
kVRq0KwfPndqRoxflDrO5IaI9UfseYtZWY3CvKdyKBG/S3wmRlgrUGqxYERwvp8d
m3AsOtU/8rIMJeAQaE/dGHXanMAyMd7lySt6RgjmCRzd4s7zer81KEZQTnSWKOnX
antyBd8bNhgGCGIFnic6Er5cjbKADi9yH1T6KoU5y/9PNzLTV2umGZVmkCK2hYew
/d/UKAmQNPoUFA6iTeIDFCXklZ85/53vl/AeHCOgP9p42H6qVj6xKwiVHVQ7haVX
86MHZhEU3Lg5VTlBql5VCwyLIv1IGx5Vj86gYw82o9QP6bm9inBTvW08GiC3YGd9
6VazVAHyj/dn2+RkIj2S1A==
`protect END_PROTECTED
