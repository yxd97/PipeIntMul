`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqih79QH/iU02+1lCtP9iPvkTELI0aRsSOk2MT+ta0IhwXv4qVUl/Bn0OIp70aEz
Pfz/qCqk1gG15IjYirrp2kWQJmOqxx0cSQFHQ6eqnlMzv0NEoJemQkKmIt5uD+yE
MuFtmh2YzfpnuBntHVj6889dqXImRLCE4hZRUWrhZbMdpkZIM+vNxH3PeeAHpDW1
Y3uUsZzSaH8vcaPQDlEHBNnM+Nc/wQsSopx9KjheIaRvEJw/rQPDVZ+x4u4vihjB
46ACxMsJxg65Xb3bMLtACw6C7Xu5H4TXP05ED/6MtZK2ZQsbcZHSGBDv79OInyfX
qIbiJUzev9adVI+nzrd4AHhxHylgtpfrCYldAWFjvYqiOmGmegc9pvBQO2FBn6bo
fx4QYc416Y7sTnvvYEdhuc4FGg8cX+bqmFha0A22FLOmxTwwKQlAhnz4w3GjysLQ
AnvcIYsYjFR+aYr57w4dimBHFgD0GGT0DEHlK8aVCc2qgUQSoaOAbt8ih3NTJ88Q
Nl6qWNgvYobgNsGXjkoLEEFF+3wa7gqvQ1PriYvTAUsKWqbPnuacAIKQi376n3I5
o1uO5hAdhJywB501MfstjJveu0fuS6+3Yk79vwbhoxOdrAA48J9rrcU/t8DQx6i5
Dj35R9TbOP5y+LpRyL/+0QdPhz7YBclZgCdt/sUaN1VFwKziLvjOzBRbdDNTSV3e
PK0sPVWPlDg2oP271DE6qg==
`protect END_PROTECTED
