`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVTFhTCBLm0lWGrvgjfRpXtJKKBOLoSw39vTGd3/6x4AS5XS5Tkkq+Cc2UOcAhD5
IFV57Xdkom8cP2xGP4Ti8zsG/k7XYp4P9MeYcRi80Hpit5OMIpUvOgwXeoEw29yJ
B8nko6JuxL4SMhH1uQvbgYfJ10MfhWi3pTu4Xo0YWYL8ko4m8cw077ioOrFeSZjb
cjX2FkKb2MpryIahB2SNPwOiVDUOCUzGLd56Y0PnMkpoj6Tfi8JvRuO0IiCnwCAU
Lxx8QNaQl0N2Yws7EoI+a6U68TjzmbRg+OtdM2jFOOxzLEwjbt6s09pjDljrhjZb
+dl4Si0ZG1EORtyFOjF8iaEkSo6xOXNX8W9e0nf2tf6tu4qdOuFhQgun9ZgY5z+c
rUKokV35Y5HAnCgQltTJI5EDRgA48QcoeoKY45h11nDf3d+00cpN3S9tb6zXwNF3
ABHj9FZyc41KwmPSVfeWBSAM+J74u2gFlHPHXemIM0VaRnhC1I8ycL94t/CtFYxn
Qb44txV6QnCgjM/luLgnLLFlf82ymvbFHktbS0IwBAd8/d3Mwydy63Hyl/qByU0h
YxnWTx0o8uovIZ+cwDnJZd2tvyHGxIDfocv+Jnp5IqyBh59IThIMASLdd85UqpfR
83gLFpHV0bRhZ7gepMQ2UxlVU914kTj6icuKRG3f+aQ+M3yxt9qWufDZSsDV337H
dLu7yNJXRapNNrtvextSSS6ug/0qma2/rbzFdJro7hYN/XDgDHOS8jXLcbjbjCz0
BOdLfZ7Jd2qAY+gwgw4m4k+FjZ1WBnztzKd12FVbPQZVRWtIyFUL2OIKM2SeoBLW
qM8DBr8gKLwSLL30nrz0WHT9AZ2aK2/HItxRshuLqGDKcs9nCTOTe+fWNZDaHl+t
4Gsh8PsqDP335iBAztVbGTajeIhzXmL1zYc0gdzKKNkOAG8lEAiQZkvuplK8zJcI
M2I4VI7YaX11F8vu2KPt8PMBVNjjTAfHbqnJtt5hXE1cm6EZniwxqW4yeU3ftexe
pH51Z6iUp+D9exb3FzumCJKm98fp3eO6L/miBb+cldJi4zSCK+55pXkf+iYa1MSI
4qVvaOS3kmo+ScDXIuDvgA34qkCio8x9lE935hJ/CdTCc3zJpblCOpTJpahi3wl+
UQtUHQgyEK2bYgrZqFNwFOu1qCaGekH9B3AHsdtZxHfDJY8BJcP72FbOz+oYoz9J
dlZzJR4fYMxFD1XVVCo1Mvv48TXyUPcyZO34CF0ECZJLbiabPZ+MDPNku3XitvEW
d7gnkYi3XAZvFX2HBULXuZvwV7m/9c9TwVfU1ZXXvC+aATtJjCHfBJp/6fEolCLR
y4aYGq+Ubuo6yVxAuibjGVMHaVWcfF4cEc+Ayv5rtfKHU75HmdtbZdRQRvEia8qZ
fsTtMN94HKPqFbtQ7lvMhdrakC8hW9dPYmf29l1macM0dpKxSM3Abcbbmbr+n/lJ
0n7dnJ6D40RI5k81577oLLgCx7sLESzACCxZlaFPAzW6kNQgh34fjUlNM1UofRUU
ugCpNYVJleLTwEYvm0fPjNoG9XBp2xDDX4A6U8vRaW+eeYojYI7AxwEM/uU248tN
t1QPJi1pj2Ox5I82zwXKBUv/7fj0lPW198AAOdLNfrFD5mGhX4td87Ru3++EPjYT
55Qf1P2X6Hv4TZnIQbczLRtv8t39dMi5PygV2MMCje0uufD4e4t4NP+shgD6s2j4
jwojusVTnA/FGQ+ehtgngfWB689M19adjXU55rZ2sMcaS3fFf6WHWatqgxGS7f4M
GdiiUbeZo/t0X1YL4u1qnpLBz1C0F14wT/JJKUeTlf3dDgXSfCYezRT2ncNtsJvI
KdnPSoZOuQtQQmsMUzs6t4wHwHS71ucOOPNJGe0W2P2jDMeBBL47NVeprUzrb03x
guv8cIV8EEoRjtziryh6yMvLbw3YDPxtNYJB8WSgBOx5KB2Z/BxY7ByLohOiQTaY
X5gBA1xumHJO5rePAsTgbyNbzxhnDCsY4+hS84AhBIDY8SwXQjsUTA6PwTud6Uhk
ZUhDbTrjZZz6p7GLEa6+zKa6v5KCzmhynwX9i/YnWo+jj1TqInnqyM6uVVMGqADM
BH1/t0yJ2xzs7CVUgJNmqZXDiBmHmPY2dCvXbPd3U74nmNCC2LPJ8VtaQ90c0kjN
a5bDOsnKhmsohEmaPA9zHGf4MJyRp3qDNLwNj2wevt3rwvYomzsccEK0HZmEe3ub
hKRg1/TBFnzLq0NzEgFR1qh1KBb8XQStW6cEdPf1+Z0vGaPqgYzRWGHTEgYc0vTq
qYiYxAR2y7tqIw7HuK73hvijnGxr2vVtdcxgy6gF5D4lPZYb87zgYgu8L0B64QhC
4AYm1IloUgaL8IOrOvsx8HDKBSagEHRdmcF3ZOBn1ukmvkpJTpIysaob+bEb0sY3
CWROTlxgpUQqCSrPddgO9gXOAXzstwGka+fVmqhnutD6djReqVHByJ6mij47Sn3q
lSo2b/v/YEfkeUmgSRCoMWm0W/Bk0CNMNGfsb2JWX7d6/EWh5ph6/DfKo74jOdu5
gRO5Xotm5pRPLnhjv31BhswQ7e8DX6ndP6TQZzCvcnPh0zJCcLvyBbNfcgqy/Avo
mJ6BSw2JW0/1LPF5IX8qhCCLezDPa5xwoGK/6oqrivLRXcif/J3+FvnD4PDUc+FO
DGjWIIE15BbI4RtZtbRpdqRk45aj94ywaSKH/LcRHPWe8TKMviGZgpp3s21d9FKn
PAklaLg3xFb3CwzTfG5HaBd5ivYbrmNVBr21xqWqaQfcf6hV9pf/YJJmoWlcOcfl
mdajwrEH/14zSznIPjgxr3PuJ2ZZlDW3LJtz8gwsCey7LgEi+WSYSZd6+bibt1zT
VN/ojEi+r7BPAQSXJ1qnxnzNo7NnbiUsrbZCGCeesk3JhBnWEJq+fBStdKVpnVGZ
0prZmwJxLcG1A3Z4irmYhNMfxxToHwTKRONIbGCgXBDVO5G/2kyqWbJoG3gNHO/A
3ZVAtBtW9VnAkVQtNr5Hylm/3bfQi1wIjbxX1JmIpVMQXW8CltLkR/x37Hrf8KCj
Q/FZMWU2ypaoIoz+y7n2fFnrb9wUIoCe1L63nC+sDh4RVqZk6vH7gE9pG2SaXVGe
tezksrLRf8yBsvWmn+FhexrR6eCauqhTjrK8QcD4gNBr7T131u85XP8MCNv0d06o
yfjZ2HeZBkEG/nqrMlJNsO+oNKLf8+GasuoUuXkZNcaQcQyFYLun2uKCZF+RKNo1
el2bgJu/Uxt3ejExYyBXG2eYn2Bg5FyPf5gn2FC2i69QOHznXBW8rPtIFZ3P9SLa
XV7m0yJiZV5iCoI8OqHGZrL/awYXYVPIpJSmghD3uD3eapGMDfCRkH4xw135Aikg
XXBu5S54c6NJFtjljK3IwXeFAfI51J2z20HtTRmzid4xMaQgUEEBX1UwU7Xfr6eS
Q3+e14UnTw6TfgOptUcun6f76n3mWnOqmyGqsMMZwCaQ2rIlbPa4lCrNjmUB8t4w
J91p9oOD0/ogcORRCEi1v1S6I4h1YC9XyP38m8HIWz4xJ7gsnQA50vY/ulk6OtB2
5c0BeEUKx71xM36ZHNYQDbfcY2AZf4YHsl/BLoOnDexcbwnkx7DDIErZO5BrJ5aY
j2p5u2k/JV8pSEy8w2oRQtjzCipFEviGXy/eloEABYDFWF1m10gm+mWQPIOJ609p
cOqttCQyNHsuBDWtw2wOARymOfEQgXotujl34g+VMTROHz3b/Lsa2FpciP4/uLLy
tkOnOA5TBUOaIozH6iD/3lwlANcxbFeratCIqlipoCJN3Rb9TOSzlUB6Za+UP1pU
dNIIUoCnUylBYER24MAQ+AIc3xlmCttQSQG4EnTzU2Y2CGtX6cLtwL/WkMY3SPI4
0QowiUma9Wd8QqiJVu0wDTKn8c0Zod2BEwHBdVN47xE8g7p6NrbN07uz6G+jOonb
8qqXz1norgDVqVFu4b6PexQ1A1dQ+kKD6jGGNK+ahd0VAuK+B6LIrioPepaLt80r
QARHJzgBetcLaRp50Mg+OLAcLof4XVGrAHNB4AdDz6IsZKN/TAuWpANnRSXT5h6i
vFbr8+taadKe23VXldS3AClzCWY5QosrvmJmiQ/w2eM7kVwcTD3gyJVlSPpmKQOL
GJ16zOhG0Tm7+20gv3wNsLmQZwlSV0fxmE4vLRpa/IY6cbPkf2RrLNNAKM9K14Eq
GD3xWPmwQTEX8WlzaJW/1R2RFermUvuknxEoKnjAAZhyzlyeFQ+8IaTDNcpZn4lK
//lErfggN1Uj48Vdu5d7hHqMqJiUZsJalATmBOqaHABN37nk1stu+B6qyJboKlz2
AQYoAt9vXfNEnt8kdU1XgriQGp4FLoQz+kq8vqpyQIYOJAtSwtPfi6R4xWj695xc
5wC17QXJzm4vDgjvqP8ISnccudsx51sJvosuwK9SWe1nCVG2weenzQ0QAdiZlzdU
IntMUZrYy4vCfAeMx0nS7VSvf2P30zt7AeLnbtxR7tCUv6rJUUtMZoJhuyA2cxXb
ETy5GBxPEJkK083XsXLFAYx3kGjE8sMGfXeO//2sLU5RTp4yn7wf5boIXUJq7nhd
lc8lTg/VJCRaO/IfRgx+o48BAm8OpQV7pERu4Eq0GVfbdf1r9S+mEs87E4yKd9vS
gLQYCvZLdipgel7MrvfGpZONsD9E3TOC3dd+qvLwe96wqN7wWAZ1/M0BHlPCepGd
zA5Tt9rmYNO8YijhHR0JtENiCtMx8/Yj2yIuIPPXp3uqMWzhp4ORmxg9VDuibo8w
gFZdeMeJBXwo9Tn0dzaIhJ2Nt7lBbuW1ZLYQ/63pgtVDGJLWKjhH7qXH47aFtmjI
yGvrtbisBRSRYIM8C5qpTbw7hNTZI2ngt4IdZ7wt0ZZ/zOWyawcCbYdJvYNLuz+Z
ZWFom0Yv8SZu0ZyGC94NlI9xlfEANo2l2vWtOJf9gFOmlTkaItoP5KyvUrubqku6
2FTTvSCD5fCCP4Gy+Iyw2CMZ0YIpxQ6YfoSVnHb5x/stmF29VnKSgd5xagJf9ECC
uAyfkoVHfepnNX7xKnI5GRLcNCcKTHgTfZZ8CbfhswqqSzKJ7bsM90e6nUwgNMTc
y2I7ZMHxkTsLqzrN5IrgRIv3iNuGT5sNImKWPkaGHfRZftuWUiXmKz+jiYTbjiqU
50QqI6NNKhmcnSXD5Y8eTL5VrorHd5PZWymv7mXNa7V2DY4vqlWtiyRF0C8vrhnB
2CPBEL7VRqZ2AxAXFUSmid4FevEkLNqpKi+RIZg+10gQL7dvUot3d7dfJqqoWJya
Kx/h0PGk5RgASX337NKcmi+7jxQHcAcSNym8jexyWUszKym4UOalAJoN3RMjCWXx
+SiAAj1n7uxxWtM4Aj2wizQm3RhoAoxveypImPKb19gMnT6SK/R4tIJ5xI67n2J1
HOk7JgGj/DPMoxKev4qru7ZwOcT5A8Cg8qQM01qjB99Ji5V9nI+MAVXuzV/Tcgw0
H5o51x2XYkezddvDqCgCLZwOb1KiKC1Vr3M3/rQj+WBWa3zqwUU84b38jaNX+i/U
T3FxzQjY0SfGkfEt+n16jpq6m+soMolZjwOV/6yIK1FDP7w6RUeK+ua8R2iqyTNf
MOGsUV65t+Plxs2k8cAQe/nccWTNbZ/cNDFac0NkI46xvVuRqV2DDNTj9IUXAJvs
wnqmtB4sRPxnR7VNthQ2Zm6mZDf5maD+L0eBIj+C1G8cd/F3cyQXe3Cqfak3F/9h
QdNLgSOrHqA9YCkbKoGfzWMbpK5PjjyDYzKzHrugq5JyZhOnGDgxkIY7nsRP7Vdi
3boyns/SN/ua/mmeZ09xFKiR2NEMQYsuiuzva83gnOBrI47luhq4OBmYtmMCMURy
wmBZZzOGvuOw7z4ERj8XVSRTwvQp/NXy3ecXGDc/pUFeNZHvbuRpFulNYIgg3slM
8FrB9+4yBFsrS1V7DnptB/tXUDWPUf4PW7IxTINfjHkdIV8PKwJ5pGjwfVQiaPhY
ACFLs2Y7yIJ/UYk7uXy9hwNQg8HrYDRAkN9fCIZqh+tbXA32bslPswdqisZaIy5D
po7MmleBRQYV/SwqTwrLwvQhZqSc73ZHYdqUbYnXfkql8rQJjXgne0c6VLbgaLxW
kiS1SkZgpv0YDJrqns67sdYmn3Mf7a8zMBWMZ6cGxRcixjrYDWzcTikXPKD7A9gV
7sAeAy1zwOphn2MOMI6wnNf22Y/V69qdlPkS/c3/qodnziP6BvO4vp/Uzj2G+0jF
q4qT51eR1MhNxBB0WA1XYc+TEiQVkLBuqj1a/I4TvKbrnHWdq6fHAiDRs3tvwhF1
PDqY0bv0NqD7i4F+AVehzdt/e1jUh69hp214RWm0clOq2ipGMJsHWbJHJ8OxVA8m
ruqQVWfEykuMLpCsId87oe74RZ/GjcKxe9W63CtB94wBsBtNfxQp0lbeDhGqgkVz
fcAo5zXRWvVGS8VE7rTriQ0ZITJqndtlyYfXhMu25sFMt3sB9yAkKhgiWncCVI83
0Z5KnuWkWVKckos6BfAhMRm/HM0SLzRNLhyiTiZJzq+rUXD11AQEWJxPjsX7qwPi
EUPtr0wKN70zOTCM4tegWqOEvQICstV2LXzyZqW52CzrI8x4KgVGhVC46pa9hEH9
sO0KKNJqDJe0BQJZv/xszPqO21ZSk6KTJy4s9BWhv7H8yt6OPshx13aLHMcvnNSF
LucI4wNhSlrKil2WC7C9r5YwankrMV97bkpOT9uwe2jY+amaEuY+lpp7BU84JSIc
MV1tV+b4ei2RggzOfxi7bqnPSSlHU5g3LR903JPdQhTvLNRc84hFOU7mHaEj+q1q
Ou522Ej8og7cNujCDxkOKhkQHcWvURN1t9226ySVXd8bF0IzByo4hitpy9t2GFK+
cAgI4SLliEzTYzmnp3F+93Do2f4pb3DL9Kqd0yvw2Fo57lAWJ+6LeaiXw+Mb0894
ikpTvZBYSiO+HZOX+N7q/EPR24eREex+7+0H6YRtjqrMIvLfPhoa08OXI+v81qH9
i1YwcASL1RYZ9JwhmgyUPJqG0t4UGsUNOYm14+4w2fjhMM4P2AVbbrjhJS9EyFzP
kwQmMkQhvz8lzty8e4fe10GV8g+ZJy7ZTsmWadeQRyUbaWw83FEPT09uQBkHSv9B
qW0L02x9yz65J3RYpU3ani28KOZ7XArWUkMf48z0o0d97/FbeDiCvupqbobvy+WU
h4+bFObmsejB2a7qdgLsANNGR6Hr50uhBFsk30gcSh7K7FdBp3AA2bu5W9XL+iEy
xhhu/95bxyiW1BlDjI57F3ReCUIvc4a0J2rzS3gMxk7QyYl6NYTnn4oFTkkIGz+9
HYzw4xDMzFcToOe3a9uEr64X6qitpf4vFGOwu7wdVkSGJeAdWYdvXCSEYZqj3/BN
9OEyw875IxzvvsePxjbK9NnIDvox+Z645UmcWkEYF8cwi5w8bYK3e+fszkLlUBlN
gCD1HVM3WGn15Mx6mRBdhLf7CZdW3K3/KyhMxdjo1hr+DHK6YLgY3e7APqfh+st1
9sKtKR+5W9PJpMCEcB/tEWfrAjyPA0qR04HGjLfFSgDoCDm/Vqx2B00wOxOzF2gN
lvt+qhbgpAtv4/7M+++fIX/I5oy6WKe+LI1FeI2HhV97nXRcDpZH5ccUG/MZi+AV
MU/n/drunWkhYibGsIUB+R6vuFv2hIuNj19kgYLzjLlSmH+NCdcCX3EglFzq7jrE
HBHZ9u1INBYvb1avK3vJ2qvcdWeajwn6A8crs5OitSMcpYb6zaVKdKz4fu6quzgR
77QN4VBlpK9NgmVrwF0t0L9oQiU/AZCvVhuJ8whdsEbCRiHVnuqc4COyipdNlrte
w42cnVT32SHv+82gjBPX8fayubytkMggzXxzXteGMiEbiioZJjfm5Fclai0HVPy9
nHQJz7OcfQ3l7q45Cg0kbL0JCvl85IEkVoe/AtP16Y8MZuyrqzScQdwqQbLDFnmy
wOmBUnKONsGCNIFAeUok0ss/d6gqn0IpUjgCg51ETMviPwXw2Xz3G/qFze47EOVS
rDnozwfEvdlKhq9e+mEkZfmKB/EHiVtHYwpNdJtgrXWlnSehd/a1+a48xvogNEDA
VJVh0NNVxe06iegtRc4f3ScFJulgWQ00uMKxUXYOBFbZIC7AywmfVk2/Gz+1vz2M
9tSX5jO2KbE14f2zjM3rRncvhsgH0eKCHmG8xytJlsQRm0wDhIEXM+U2VyIyPIyN
aBY8HxjzLlAI84bhwH3hMhm+NhnvqJNo5xxOrRTgWv9BFsTBMrC72U8YvVD6no9n
s9K+VmbKT6yMDKX5u7yri5NJ+miL86rJ5LnIfCY8F+9cIbV23PK94HH68W5XyjdN
sjqDwy9t4FHzn46eVWNzejEa92jaZ238KSdELs/g3oawePvFZpFCn2BRZeTs8rFA
bfikmJrPgciJXX38LrOVeXw7MBlXXdue69GsDKQeSXix39lNUjdJO3ozRglpwtdH
5aRrCvZaH2FiW62of9vKe1pN9s2/U0eSVLHtSKyJrP3IwD8uhNDHxUMP/Pfeub6V
R45DtJ2N55YachP3435YShwCwzepZD+aR3rXzzPq0taYZBUEs8V2czAmtxCUCGFD
NlFR5/Qej8FWyGzJhlijn+BfvsEGrqI2KLPzXUD54XkiKRF9JeMPMmAfeZw9CQLQ
7CtA0mjWuFvsx8xH1k1dF/v2pmnSlkv06nKnmFheuL03c5shJwOA9KBg7gFsxq8A
C8lgCPi6kufEY2qkJTPWEolPCtDKH1kpy9sRz040R1fhdmoEBTfUIzcSu1tbllO5
UAAVX3wBiO6eIYeUzTaG8WkciJ5+U81o4QmyuGInB089RDMK5vq7DE47L0EwcUFf
6jOgEvNMaXunZgo+zJ8LcX1ThyomWqi0WhX+ci1JvwE3B6LEm0Q67Z8UBhfuzSu9
iVLwAdURSIQNCHDAa1zETyfPcE0Lid18t5cfhmjGFu6K8hvrj+VyxPMa0SvJeFHo
Xw0LDNgPAsuEFlkS5cMvqZ4SErCGZnx16UICfPqVMimefSvirQnB3nl0dq3twC2g
+pIY23fOMfPHxwpZu/Q26/yAAs77J7+j9wAF7V3Km75JAg8ZtO2+R7ZyYZkOhhxK
jlcbMPqH3JULIPbkrZjeDjWDhoE6emGVMRTCmUyzCPno++pKLsPtrAXEK00ubV2t
G0yzbsa5SqkstJST9J/o7qBatqGSBaoyj+PBktSGsFGwrPpv2peL1CZ0qtdHJTtD
Zfdt5Gp+lSWaSpaoCUUw0LqMWcV4YnpeeyemEt2nHFiRenCnZNCy/KSRjADW6BrH
zt4LctyWMxsUACEeT/yqoGp1sdLO9SoSGOyUvtFa3AmUX9Bi6ysPZsZ5zpkAtbaP
Q7rWBjgF2vtqQdh2bv8QPSKTKGnQye45u7KHXVfVJPcoSaHcrC10lvhrsAv4WbBn
ZpYqlaXs3TU9pD/yqCpuarLF/EtL4+7K71kR3qxIKCPeg9AFX0HAui+DvUwldnBJ
YO9HXgZHtcqbaLamOF0kQYIPCAySKjq1xZmMGVmck/e0wCQJ6kcUO+i9f3/MdP3w
JzQfrtMDd4FzWFc/JerpP8fwOSAMgfS2UKahTLbiXLf7xVudcYim4eMOkQVYhOj8
3XCEC6dLdduqLhcJ61SYZmYCMS5ZRu901ZGBH//AT38bzpLGDqRD01Je1n6CD/SY
xK32e/4rV1d6OXT8gN2Qwn9mVolrzwRbY+RB5MZpG24nY6ZQZuSbo5s0DQv5Fc0H
8ir6JSWfp1BP7tvkqsXwtcpQPv4cZHW0RrSmPdG56g82akgoKL61P3gWDc78ZiWL
fwXM35ux2LyqSQix2RWcq/Pt6Ua9/HEwFhA/GV9zWyp9mEJXLbvCQQVSTTl7z4dA
LV9xoKWYJb/TYvgZEVuMVUdvWqany/0hqp8E2X2yABPP7fnmG8S0h47TUwk+d4SR
cnOGdbFcbG+SealGih31iKPTuIOueNvr0fzjbNyF8+0nYOQWXQH5MJij5HgWffwF
3LyQjyiv693yEh33ZU59OIeRgVb4nKrr5CTt4Mb1P1Mj62J9DptiuI79m5nJ3GBY
mDJmFzwDN02QPQ2zoViA/O+cyhfvB9rfyawkHjFwgQbyetRv9DR8g4vbGbSlEPSj
+6wDROlUwRI8W0Tv3kIFQeB/LNJYJFoLj7k0QYaZTrjkNtkgYQGd3D6684yFDc5T
hExo/aTamMvu730jbvhP4CIVF1OFuHL9FVlWvt3xGWDZ50iLgmVrLanI9sIjomeb
SWZUDTROwfNSSP3wQlmYyaRcx7RbT+U6ixPTwLxVs8kIZT9mFq5kcjqG3Zbjmpc0
6aGU5Oy2+NlcyDPBlORS17GFvdI1HRWr40NLmnGpHtIwOt340QtV0+IxwgUa9BQN
KA4NANxhNcmJeFzrxD7VuBYiDUAGTGTriHOOOWLzDpHRIYW3GNoMZaZp+DfZ8lAd
wtNIW0fg3Tt5KJXH8FlrTmDsMOuxK3Bh6eAcBfiNblvzyDKDrx2y/yXttTAMun/t
VBBuWQb1wfK2MYMSqOf5hXMS5lAGBXYjd+YNHo3zWNU0OwAEYdgsJ5rE2kZTDVh+
IV+wIEeafrnz188phtLbSGQtgun/kFTFUkzr96If4gdI8pRYg6YWTL1RJYb5GV1Y
j+reIZdV+x6u+ng4Z8NccwfQp2G4jK/claL6S1c90nPO12k6O8P30GiKY5rT2QSG
aTqoqsNBWLdRf0/K/CaXr5aGupSUn5YhqjH4unFzHLXQZJm2o7lHn1WnEcwhl56H
fPSN5GR9+5JwvW5Lk7Konw33wehEK7KmGNf4AjQOXBJZFzHxjRuRfAjYIjueXZRA
vqIZIhPAG/I5vcDDPaeBfPPfq8uT60kp+YDdz4OppS7zMQRLIalmha59mUiTcND1
8LD2itfmMz3mYbe2RxH3Bxw0FTxNaQu56k9tsvEWecrg4Pg/2kgPGH2wQuyJ8Rkr
8lj8Gv1MC5NSaBuIsbZa5IQ3KPpK4oxOnLbx+vBpmclRohHNFfTniarwSJ+4E0bd
k3Ba/mdUF3FYp+ryoBTAuqZo6LjP9u1N7Ii7iAHBgaBf24p1m9B6BIJJsukFnNYL
kXhRA4o/BvMY5H3PXqn7X/RmbVXuZcpDb5QNLa7Ofinda1KfUKj7z5X7QQXnL3Bn
8roaHgHn6ZMKvZB+9ClWij2M3rhoOYShtizwwFNSuv425NB4pM1egMnql+A/fXjc
0fHF2v2zzEVD02b2C0EHOyXLAYKBlXh/Owe5hOfRP665XFHU3NMOlDwmpKRwMNah
2ajmcCKJ2fxMjsQ8ni0Joaw2T+YyPBLSVywRYDu16xaTJsie75JYesoWfArq8xnQ
+H1qQNuXrFoWXRmsDb0Tka3zTzeawu7bPRRYUfYT15rYSFDf5pRyo4vithcml6N5
MLQawdlQBMjRl9S57EWltlYfE3FvC7RHCThj+J64qLevmKOqr7I1pvKGCg5jJ2m0
6ZifJHPHa0bKvZtYrAxKx/Vy2EoGa8H61Z/LEZS7Wp9ZScSYMd5ooeduOdoIzDfE
YWSiF3corPhAvdVgZt++MShBdWC9ke6qesIrbokhsyCfhC/lXzZwMH2aDeDs9/LX
6bHe8cJZxYPhzs5merTQKfk60VEpLeCo5vJTfk14PCKs8+jm7naY/PqXnovzrDcI
ztRkLO8Ot4t2+x7XpOAlIG/H6m8Yu00m1QpRqJ7A+vypU72mqHU7MgglFMhyQsEl
6z1zHI4SfH9vykt9SfNWIpT7mg2SrEd22nq69CAwWUMI7IY/yo6iag7cCksmii2J
EaB+uNdRaAyFqJLG+SgPg/nmRxG4tF1lTPjeIJnyJAYoWPFUp3YiIZngCCAbaDr9
Gxu/310XdeE5kWV4CBu3sbtz5rxN65VzbbJPssQHeE/eHI1pxvtiLLd5nMFa3hYU
Me1S4YmOVwd0CTy5oOdc2/s6nJo48zXtim7gUg4GsYWAncENQCwJTSCI8b2ddDRz
d5mtt0UIjlBlivn5RXbB+B4CQZ4JQaX1HEZH+n+pIwCub/40ffj95Xf70PIFJ8xj
A2QFmDmn7ieavuNlMgLzY1HmibzYncC0WHTCZZdAh8zfMlx9QWKc5+5DTHED50c6
s3H3E6No6OzfSSGb+FzQDkPy0bqH/S4PB/26jwsBeoayZoiDS5fLc+X28LRr0VYl
qUamekyxaLjgxkTIzWDVN75JPqA4TA8b1oF1oZS7DOcpXQicnHJupmM5hFLxjX5p
t/eiCJMFfyxvMJi1EUWsjhT9aXIU8h5Y3W/vYlBsTnEMd6It9gHZ1sRX9Q2rjTO5
PGK1+E3uQRMmcuvNqH8nenWgkklik36Q14R5WCSD4OBAFqGvRJ4dZzd+fLQdKh9k
MO6R7tpYv0NWj83B8LroRjfAy9p9lqWNdl+XSxLloyX6YQQk2QEcB6JI2UPaJC/u
qu+ljWFr/G2RwqwjLBGtx4FMb3o6s3woA9Wbxdh/nrhmA5Za2ylAbydRe5Wn5Zv2
WnBGFDKp1LaBlN80ehEXUGyYTJLI0/SHtHW5l47Wp97qOCXNK1ucTxx/0tU6vfD4
85CQ2rpKx9cMea9JATD76fOjkMYnvCYANG8JBynJpfK4E39skBHaQ9mhAYSM8t7D
Of2KICWcDNSFJ07ht1+pNEnjS/Lh2KHJvUwFoLeuwbMMO4cpZd0lfquJA1tZM5LY
PX7UH87s6OY7gpk/JNRjP6bm8F2OWbKz8YyWBp7Xmqax2wu1HUHDEatxSrPyiIkJ
uWhqaBqIKTdPuZuyGnTXw37Uw/KlQGHnqvQvpSa0XNYYNNdyV7hvhSHm8i9/UCD+
tkziAj0qd1B/LaLWbtz280oNSxVMbocAfF/P608lrmh5OknThIwEIh54+R+iYYbG
u1UdiS6iQKiwcIxYEeJkA6SWjNRnBLGrNzmWyaNAlINe2v1q6ua0pCsal3hFAGK8
ytS0LMyeJfrj3DDXjMAZ5iuYdr0Oj6PiFU0U/23FTBCkTQ0CEmEOrePL6BDWPpUP
Qg5x8J2KIWY/3ufcN8+hKVKiQoG21Tvtjcnn6Gd+xVcRnkMpJYqMPPl0MTzKNZnN
tX0ERe807VRTrPOWf79eAPTlyKu8TwdfX61IDAjSPs22hFqpTdi8gBsMYHip9UGs
HD4D3FZH+z9vunV7y3vYEcKPKGLAcz+H3JsMHSrZq9WJfeOcnUfm4285mZVWpS4n
vBIWojEsEFMyfgaconITeJqE3iWV2992hvrS7kjOkySz/wDv8uvLxNiCTMSUYrc0
V7/0ZS0ik6ZqoqzF5a97fKBarM/Y1e8IlzsKeU4imygPFIbTZ9aGitpJ05R96Aj1
e2UzS9a3FbBLFOGZunwy4ZzXSTFbERkJ+kpUHCUjqgDP5ySL+6MTGWZOBeKSi93e
9jugj7CsH+w4Q7EDxubw1KNycyryjdmeafK7B7ZSdefLU4qLyDm58lVO8VSloMGU
2cqZQxLdc97/6vEuGV4P54inLEx+p0HmZ9Cf5qi3dOQ0FNoVMhpTiOGJPVExVFYq
tLlzlPeK2GA5kxibAxJa/auEy31g9tssUm6PhFRkTr68QUuIFRaFyDeVe1CrEopu
z6/YIO8dZ2n/ec5FkPQAlfXQqrPdK6LSkhPCgsXKm7hpc3QCAAoS7EV6LoN+gSRk
xKI1hBveXPZUTLyL9ef8bL1AfsnxOSZWQwTWBs+i2ITOLZY1auyAvYaQaFjce1Ij
UAw6ksPst+VkjkfaDoD1zj23WLNwuaLdUoMCZJi7Ktl1G9Rrw/T2VsYCVDM6+Agn
mWT7oNcmmcVv+MDb46oDfhQOjkhhxDNJF+p+YlT2DIJUHAGcxTUxy7yMt9NpmM94
bUL2MrY5Mo62JGayrSeRP4hG3wSXhiCkXcQHPqzZrJq+bt45OqMAJsIuR3ldDrEu
9y7JHEFip/BOLrxrwUoc/JcdcS8M/kgZbbjAPWfNqZSqk+tJDTD+x+5yzUguT+SE
IYA8e0g86eBxSA+4J78Os5yrh6zcv0aJq7cnn0liF5fBJlxdt6ZucF6zNoXpg7Vk
k+HEsvLkDfKmDhZ+M65QOmPQ0C95/VSe8TImCy3UOTbQZJuEBUzS2vLazXa7DWPm
1xrFYEH1/dPP2db59a68HHydfTP8t49Q7JQoD5CuNPFCMyoa8Aab0XiypCDWD3FY
izFZ0rwGHSUdUrPWdpVQ4Zzg28gCKtbc4GdjxZ9fHYQUmgcY/gtSs1hvKJG+tTBd
8X/bC+9gzV17wGceCyJjfEn80i1DnGqpjBrkLl8p19mHwJnq1XFRpvM5Qm3Qq/bD
Y+2Ky5VyRWnWUHvA6WxtvLhSuj894xcrEwXNvU3QmIk69ZWuDqmu8RncqvwwGi1u
hw3gvnPwZgM7kqGJ9O1hYwLY/tzZAdDwWweWgPNNjm3v52IeRsxKAfcYfqNFnkdq
MH3PtQmyeHU1BcX92ZfGGV/QrtQAFnHKEjqCoFj8FkyiKa/E0XtmgThICGqpjMZx
wrdaYrosXvZYFKeUiilFtulkshGMF7A43/6mn/fzn7vmHQZtO7q92rQQMhA+VzcA
lWxz+P0F1PFKJ+vXCQTH6Q6659Iem4SgR0Ain0+AHGtw+rWdP2eE0WDG6pAks0RL
wf0VS5Fqy0ASsdHRbYfHTMRv6l2Jy4c99hJYFzyQiHVjnrhb0Qf3E48jOk6G6Yrx
iSFA6NpNXwDNSO1ssWxuorSRDNDoKuROjtvmsg8ocZJqhICTcVoy2HWAWV3BZq7s
FMkNGRLeDq0EKNgRxFA++W/eJZU1kLq4IkpJ7dkKV96a656oJb7HfySaZjsouxL5
bznZ44TqNl1bITsVjSnIJ2bOmU75qOTRgA+Snn9w2NeQbeMH/PgbrdURnSbTDGHz
LBZzboz1PttpdPI7SsgqwOp3dr+jxV0PwRnPltdD4Zrc34RejKLaZOVtvxTaW2zu
F+b5QUcDU/46SjIwn15m4M1YzlYeD3k8xr+BeGMfgAY6Id/GeJSToZpMXMSgUjAb
Cmz96RherwzxJ3R6CeriT8hcYMlkXye+SkJOWbNgfHJ35tv09801dSRNwXbephRl
dUOA6JNrve3jBSyL0WmRvkl2Elllc2MBalmB/6CcpDj5VOfrNAaY+8cvlojgy5HA
MWhMWi1szH3yMF/733Y+zKN57SeI5/0YFfO8wUmJm4j5X/wDGUE0LTysyx0LbeLg
E5DHr3qSz+iiVdYmOnyGwVmk35hn2nBh3Iqd8cB42PpGBfnCAGCQqgu51JgpbjqI
oXURM612F0btOakx8wFYCScB319Hosw/KRrIhdaEksOzpgrwAGcKX7ILwx4qXnlX
skkKxHNpr0sLCdo/YFELR5zlTWAgHaeoraM+EFEX0g5SiKLj6f7L5IlGam0nJ76g
k+tz0cdy1AiiyUzqOkaJtiNZs16YncZHVjOYrdRwxzSwhyaM1oAUGRnj6PW3Rt0O
bRfvqcvp4Yow9g56s0jBdgcJIJ3ORZhZjlOinXOcTwb6/ejjNaYnJjrMONnKsiVu
b9XhJpaZxNX2PKpoNxPo9BbDgXJ5u06pfXRtOc5/oey2DnuKNZZ0Ilk5DEUzBij3
7j9eakhviALWaLJnj6tM0j73QNx3Obxo0sXKQ+xB+rZQrlgnPPAGnKltpABbfIYq
dO3+ng3p23BScU8srlmFBBenzEFsInxpVv3bldfIPV4wlOXye9TjwZ7MAVFASSfq
cBTXyW/HMFff7i+8L/Lb5yaPaFD8mX47j/vHVXAhRhtOABZimqT0jWGkuhmjjLeL
tCTpMwGQqZvsys9H6A//+wtM8c/Q8vsWqd0VwRNFCRA16DrOrxKZeNN6ivXiDEpW
FPk2s9o+SCWDQaiWn8DFzmNP/Ekb6PRjrzjiXAG84YQ6BlhKzll2B2Gw3m+TtORy
d8Vij0nIXpb3TfDgn0aMuqSjcke5pQAPFiNaooHE5pc1kTGFTgNdQ9Y2/2HplaKu
Y56ET55AiOSTbNRF5txxLXmxov6QMt0z0hQpwF/lN3b4JCcqNA7Si3Ks5vxG2HvU
fl1I+pOWycDNCjjGK1LrAk1mh5yEu/eEDu5ftrSp9+kR1M9+/p+v/W+lROltUhHV
6UZcOxExO9rr4DozAP64vJL8Xis9nCC8PJlGSGM76od3U80/lcL8ZXQ+OkK81pIh
FnQW9xEWdtK/S3w1DHPjJbENPmVdfpY65FjTBG/+6WwYpVfaslAdtpMSW6rZSOxV
IPJapYMCgPa00Y55kTkRvzYpJh6JP6XQAUrJ3APoYpxko/mdL6CPO7eDgMx4Wqu+
b03fuu1KYD2vKhRWVyv1ABJIiNUwRa4GywyA0grwcpWC6NHIDS4fs0uJFBAB3qcX
5AnRpuF6Hps7DD+HQAjJhdUeSKNNWf1tlVk8aD+GDhbOGFmqEuFs9KE0wysyiJQo
nvu1yF+bQbgEua5MvOozTEcXr38CqqBlgKp7G3cL6kJAUvuOLriwbsCBNv2lUDVh
dNgggKIpVUkmN5g7YyQxBX0gnoa5EdiJwtHskOHMgaOQYsXwsxDhEkoE4kMK7sps
I98tSb0Lx0atxMX5jDw96XEkRVHKn3Abu67SLLlc95AfTS5NR54npdklc/Az92FC
h6My7oA5XFL25QIeWIi3eZr4X0V5gev0209yW+SsiNItanOkAKkTrcCm5iN+IhT+
UTeCoWp8l6FClfCjfSIUK149j2uIhN/d5ZnDuggtQjentm/+HvI/hhTQrTm8WSyu
1KeEolDMVyJkWsIow8F/Yl4xjcjB72X+aNeXwTbIPYItins4oNsljaLujYWt3tUb
ihfyjfe6YHUOggP7apaw6c9WpprsqxYSZymWdJBnxivK2Hk1p46y6NtGKiA5IWWQ
sd7fz3yVZqyIHcXMGzYDUjFL3OSE10uLvBCKNIaXOck9VVRcz3TxcPPWry4/8qq5
T76qDppCK/+H9+2IsQs++MANVPBhJtnsFnKOGkbE34rUBIHwBBw/HUmoIyR848Qx
IFMNDhwQmImHebKnup8qA/K2ckRh7HYVGmbe5KIa/2Pqwdrh6VEdmrMWxsXDUaLT
Ws4h23dLR15Vlbs6cLjOlDsu0FTht6bbgWH7Drmb/pirhmSaxseXZ2XDVIhf44n4
19NCWocpA0Wr8a9PLkbRCxklZMFidFItTSYaziNia0JITZWyUevkMEDFeCgR4Lvy
CzCWkp630ju3hlt1UoYXhIi90oplfIhzaghcDDxcK+y5BxDlN3oYrnoI+mpe50j9
mi7VYI+x/hvV/QGYhMvQAJCC3D2hk3WUrE/5LlzgdzFIN0JUgK4QDUXTGHcW1zEs
hbbF0pSLC3w/dJUiMP4XORiu6jgADkZVvjUXRW7FthbPmEcNl+L9sOCoi19vuvb0
JXFOhTm/OjpUp6YfaNoKF5dc6Dcp4dfMvZIippcL53DkvlnRpnOl5W/SmulYC5I/
bowXPFJOROFhNjEnhPZjBIPyGRBTwUyQafXOOGmitVIZvWbrdlYdyj9Pjo1W3rnk
XVhb+DijDOJMyes1NbW+mtVq1UwJrqxq1csxs3fxRobZulVQtyNHYv2T8LSg8rci
z2P1fiLdL7n6D1x4Qq7qKFgXwv/57IB5APzcPEl6D470unoy9/BU/+Fq7U5aQ2TW
8m/7Mf5nbWSdG0F/qjNMtRgvkTZHc229C1GXzYGUG+6W3h+lPnjBLePbZZbvVtUo
1Z8OV2ruxFL6HAhHMQ4uD1GbVvWLmwyicOm1lHS/G3CxQM91xDY5I/WEC5vqqvyB
MitY/X8fFQRtB/wgPl5vd/yH49wW5qrcjYqHfDsew5Ih+G9jd/ECPh/3sCuDOhRm
91Mx1NrZiwO5G2bKOGEx4b4tmlsSeZfWLFAmWm6yHatx/mNXX76DD63X+RIaiGZM
xd/uQkTEr+L7GrKyOjw4usSjDH/5QsbzMEM2oEqqvJZ1zP+zzuLCUe0OHwy5BKSu
hPaoCsuapm39GpJg6cS3kflqLuRMLmrXIrJwOoxoPpcXO+YL5kHsp4QGvuKJu4B1
e+Vrcb6F7BE3I8MPk7u8R9ucIZLHBv9WHx+Z/nVLAGiYd6sp5aEmLXJhV/PGTO5l
EWvOZ7GNkZpXgPzQnoTPHkZzTabfdnbIqS2+s4rELXNC5YRLudN9/NsNwdD4NCAe
g2KUqobciSjrBnVSnf9OZJpDbp10tkWgnfGH6hgBgZ2nlIRwupW1UoAkd71cAtfU
PApqQbfQgF8POh3GjcFLOJGHj00ehKs8g+67Xp8r8aIG2FBmNXVQipKXuYkhSMS1
9mkxUtilpo9ORMNSHP1aX10oO3oTGbp06lgvkD7w1d1l3VCLAR17YT+FsKlpd9IU
Op2RGXAIy7+6ibqjfihHtIgCdpKsgqoLsI2aisgMQlMN30opHgfeVU3GNEi4x2HS
MiwEaJcz0TLEMqjGm1u6Imr76cd9/0E5CoRhK8XLpDHJ+1AwqgnjO1X8AZEjNl/M
wTXCThXE1NsuPvRAbpXKcTkHOiDHJerZVp6rReDMSNldaqi4IFKUf6XSFRkpcTZ8
ClBZfhlUdG2JdMTdgHiRheOb3wJPxgCBzIJxfh6IWpP6qyuNqf6v/u0u6KQK/R75
Qne4PifRw7e4hVotp1lItIC09ui3z3QXbUr/JX6xs1dMe6X1OB/DZXbUrk2/19VZ
3S1UD1TVudx/xE53VhFmbJRvVtChxGvGu05khgNWMrzmvMOJEb+NPn160tVT5DJc
iENmT9wecT9WrdfLvX0lOsDx8ybUR/Qpb4QvCiRJKFXpU3bWeYRIP4+l+9FUPeX0
JWnsAKG4YvdGP3h/SbQJ/pfJoU/xKiLDRjl2vaMepgyqBV4TL/h0TIMZE9fE4exl
TV/jC0/ToSyMJVBsxRAWmANqmuqlm9MKto5siWSbL2xeud6jgagd/sdpTcm6PLHY
tECTBsszKy6kI8djr03B27WPZpL6M4lglmx7A0n1vHX8EvB2gG/C2nBhiqCA3t9v
Kkkxb5yr1lCKg25UYOV0V4ln7kWes294DYnhOkbHpUqeV0JgstrEBeiI9mLZnObW
O8X95pyXNc5sN4CpumOwBdK2fOEwcOgfGVA7Q90XKKgrfQ96rYF4ZVaYlrWLk0WO
4iM43Q+Y7sCQGr3CdNAiPIc8Qa6ZgHWMfFF5eQHd88c7Q/FAn8BgOjhzkctpj0Uz
A5MtR9qE+wdKVrViFMSlepG04lv1cXI2P8HrC6R4R2Ou+JYBjlJx+hLS6oTG0gju
UheJ9uHYKbYR9+cQxnhrrH+tUz+iWkIAO2+7znQyaGNoh40Z/WSKeFP0ZXKNheGy
Qo2sfkrnFZnZMYn4qLGYxFuE6wPP850WohHg7xsImJgLv4+Ew8x1hKKSesHSLtnR
4JVIMLyRtFdrggiaKAaQ7EYgpDpHTK8L8QqIerzf7Q7KL2C5mqC8jaUv9K9w3BAN
0jgtqI9HQYSdJX6J4zDANg5NZHmqhKmTx6haC3quNb1Evxyx/6Rw8xihm4tAPC1o
JNdtUef9z0DfgkfCaqRPrwfIP7Bp59mGMDrkooX0/AZCjoLeuZUdnRZK18Bjv2eq
jFYflCrVThZXwOi6Y5a8Sw4N38KcKng3gf7J49oHVs72U6cIJI2OuFKQXUuxm4NL
x8nhvRl6JUtSJ5/0wcd42cxxmJlS22wBgeTz888mWKgY3bgj5Idkts+IMMjS3FPC
b7Bt3TzrDxITLayNQ2utSUHy2r7U7yhUhqv8VQEgDI++pIbMg9JwnA2T4xHkskqF
vRekTozLykWIHWk9pJT+wLnMQTlrdV0F8PY5QeziVdbQEs1AF2UvYJGaCoFHtzvD
x7e8klRyon/BqqyQiP0qebrH5i53yqet25a5H0k+hJKUaQiRACSWss6uk4A+7DvO
DrZKACAXJDPj8wzlYKaUK+EvC3StfAeASDEeFjMDKo6yXCN37WUhi3QY48IFGWcX
PrGaTWFhMDHYKfHLhYYfu+oBCGVXPdjUOH1tRaiErjdShDUIhJ2mi1NCUQOW+oYh
oCx2su3KdOSTmiePjDtD4BWE8mqdubS2Nhz9POdbGVbVtUfx7EWdcDxMwrwFtxlZ
N6slZTam/N3WjvS9ceJYVOLYQOLLC0BSdwDpDnipfuSksFS3vVTmSCv7sTI5oC76
L8MZrl4wUevaIb0A0c1OgMcw/yZ0zGLfDrsoswpwWfsUMOaWJPXL/I1aX3WYKG3v
VX96u/V6oxHSCY7XzHlJsMILcpqpak40xw4ESTwxY6Wkn/RiGdSdYDTd81h5BAQB
no29RxE5wA3MpIpCgXBPJfbmxInBks7IC8Fcc3J7f1bu3c+FrXNn5LsYSIjyaLVZ
AiAfj/tdYw704vx5xrLKtdUEkNHhu3cawoAkxT8fDcA=
`protect END_PROTECTED
