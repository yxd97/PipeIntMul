`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c68RCZCv1fJbVDKWdo/QZVR7oc34iWeHB3jBTh7/3vCRfHQfTe7NJXvTtN1R7bfa
Z6sNMrUh62Q8wIh81kLGZJxlEFNe4s+h+7aJd8Z9//Dgf6AH85dPaG4Ep7wCKIYN
RhXB+AS8kuQVhV+54cX0Hu1i8V+NfmcKsVE2vYF20VGoxFcZkAp+SCiYldO47Ahi
L3R661poLIm4e8qp5risxpkckBKiNTKp8ICCK3TPZG9nWY9Bdmnn6i9FxsHu2h2w
RK6Y8UyKJ/B86mqCpZJMcpAOmzw67z0L6u+LMPLVdxXURTx89rEWewWuG3rxSBCS
MGMl8ultwdLBaZz6+d/jA3LvI5EGAXUJ+GRs4iEhs9UgntVKpvalwobNldbUt+Fd
hFzgYXuouctNAzWiCURQ3BMVFY+Wnyu/bEgjbBVQL4bgbpmRjAPul8AXQOkchPVt
gVFZwCANLqlTESAbJAdwFBojVHX75Q04uYH7d2jIBEwBUcOrImXzez6WWDi9167n
`protect END_PROTECTED
