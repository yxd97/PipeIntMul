`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ckQEDjUeLTyNXXHMsCh7wmhvVyKxNyvU9MqyDwuJRi0jNf34rqesMwfw3NNVFHBJ
XccYZqaHwqo+NwkQ2la/ziJgkpt4PfC1+NmRXwh0PFnTqpJfjkCIqAGu386hDA1Q
PurGbePiv2ovXqLrgmp2/6wv39EvR9BjLahfJ5HiDovjX0Pw/nEEhdZnMtQyIeV6
gJTSlbU/lNmI+lyYfi829fZlhJCEnXiGmclPsL7HhDNQPA9fgnhPjgpii1gfpZge
/oFbsaR7GAWSfjQ4KMyc92pg96wbTFExUOiR4Pw9aObnsJHAaJgzgyGWXt9HRKyq
imKka4HEup0uHEnxv9+XCzN0Nhgn73kuksgQESb7Lwy2nA+gJvhimFcDuehnIsHu
6yqcKHDQRMfQPdKRxexU/J0UiLkLAatRDwwTo1+MgUzZ7OStYGGqsCZqRo+/oi5u
Cl+DJDgzy6qB661ZStuYXUI0KxMaIov9aQgYQbSI4s/0aQJzNb1Vk+EGg3cn6vCO
jy2zfZCd1vK3VUMh/8NS1A+M5mJHgRSUhzyghU1FoSKoo3+Kz8lFdq/4Fe3sHxNf
992ec82HJDjo8VLSFx4LM2VFcUQWxg7Tq8/Ljm7wSQ632Eebt80rJZrh+BCjjet2
d7hqyufqD+H38YVcBXLy4mrVHQ8+/vXwyt7EtLH7MxqQvg3NCEoLJrJuuXGO+Y/m
F1zhtyIMo8q03FIOMxn9SCucqoWsh/LcfzJe+51r5L6Q16XxcySElyT0TVvV7ILx
s9ORlD780f93JEFtYRjRHam+4MkyX7vLVxe9/7XpTs9U9/i1Va/nmo5SLglR0zbo
7l4iQSYTZxB0bIjguwQwD7Q8PM8mJ9jsqOy6PhqZjRDhD5+eQbPfEyCVOG91bRmv
9CwwlQ8aIhj+A4FEI/rUabIhw3Swcda0n80eaKyKoiBiCImi3zWP8VlyarYdXGMJ
BtmORWUeyPMNJ76Oj+cFTQ==
`protect END_PROTECTED
