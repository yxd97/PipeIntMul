`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8pKwipjQOeMvVbGoGbqpVahoHrQQoP+hYR/Bo3ASS9y5wQ9QQg9Yn50pz0QhmiEM
ZZfsAWJY0pc16wJa5+xvpIoMCA6W20E73kgyigf4AJYmVvDICzumSxxTx2T1flFb
/s7yDIuKU3LrvudnkXPw2CdHiGD9c5j90U933sQshIKbe/gCtQv0UUh5pXJzbAtm
bmbhQr5lFHrGw6qc7Eqy27qRWCUdTA1u0qDEB+USUpFb8jgJx3JiJTV4lPD5TLIU
cL5DQvCsQz539hpWWgxTuDpTNLpNDVeOTBldNe3NdCrUj9l9z4rBCh7Q7VmOD5lr
wrvtlMIF4CGYc6deD+RJ2Q==
`protect END_PROTECTED
