`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvNO3y9y1c4xppRs6PH7dZ5gNL+2NdBmXwkj6pMlHByTy1YR6GS/Ngnq8i2oiiAK
OwC6gd+9S+MrpNS0fFwuzjMxDrE1s84Hnm8vQpxjNbsIag5oSv408YSAW+HiVA0c
HxAwDx4B0Xvs3tNjHT7/O2uBb9W1yscj2CGH2nLCm3rt2MNdKXImPUIYtSWeTA8q
7bGuHUpFTSbthbPBHP4InmaCca5ftSdgxS4weaVhzoXHG3pUL4JbnD2sxo3X6SKh
61nEkmyLYLC1iH+0L1kkyd4Hc6cK1rUpB34kSJZm2rrKXXz7tyoofplaVIiDRb0e
e+MQQioTEts4qPAlxQCAurwUBZmKNQGYyNpU/BOu2PaY8MAJbyJIR5Yhp7YL9sxG
QALcmfIU8qH9fQZh7cQrT2FaC30r8V1SS1SS3DmEDgIoN9IE1iuO0k/KjdZutbt8
mQ3Y4h2p9+guDNSDV8RNjTekSzJd8qfJ1xICcbQLVeXYIfTTXjpwnOVPITrIn6VN
alnb4sMJ6exGXaLkdYeNakuNsBL6PZ52WqDO83fS1dfc91QzgPGQfWSvl3yR0A5O
s8hWd7oLrE11XU4vkvwjumMN/wdvsBOzFkjQdPtAhCApWErNPIWtfDeAFsKdXpSq
sGpbxQFRlLJUC0I7TvIP6tsvc/2QGA3Ng7cH022uSVw=
`protect END_PROTECTED
