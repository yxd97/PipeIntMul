`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F24KOtA6h330khKxkjC4kvY9//baoRvhEhVei+Ok3dSkRq6RUuuzJxDq9qFr4yHX
6K+dTZvzhK47xlgS+0aQ79eNHAyBV1Pmt4GceLrZbkpnwZpXFQlaXXZNrn31ifK/
cgA0lKf8iFrR0VGiEfE+ZRJMgMJ/FnqAqTKtsK0UTRCymyA6oTsW8XPqVNj4lIU0
w3v0sozOYSARbHmW7KRn65AHQPL6jpSaEhbp6ZCB5orNpOHcvV2j5F4JDwXgXcDY
gA+7LNpNrB/m+FYWWwavD2PWWx2D4MysgspDMVEEiCsVV/5TXjUtSQVYrQFoNi8t
8OKIM8mQmJ/w9cyPBure6UQfPvC1VAtfFFrfMedb9NaJom61XY+29BJqaWxg0XY7
`protect END_PROTECTED
