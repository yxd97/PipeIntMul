`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WXj2gdqqTFi97a2JGSr0AunWQq/0Tb90UxBCM4Mt097UrLsM4FrEAp3wZeML3WcJ
xSPZp/rgyZIYCTOATmHc5mstEW5TmjPON5S8+PKG/zdiJwMO6JTzrbRcAywQeULM
aNnw1kodXUCUyM4AgeFAZUiuHoQObjo1g2rvRPAhad8qOSrwTgS2SIysHAcuEWZ3
LWKnXzZSw7VWqxmxHh23ccW2TubJGWk1Y5cqW7FYrVWICqfZUumHFxbCWluhHdPH
hoU9pi3jv1ZfOna7n2JUYbnU77x3pskbh6porFFao5Kjvwi3tJlZdyGAyJnYbSEi
fWtxPJY5dXhAgrRtUK4ydf58Ie6y5slFwTOFulyJnKZ5hxZVqjWAOL4tINCiZDYW
ikqMuwEyCyuRg5GKxc1Dl4NifM6/T4y11KNmOfwgmulz/mVjtyd2FWyCMEyzmr7z
`protect END_PROTECTED
