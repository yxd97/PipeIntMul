`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KSeHYmCSK4Iq8QheIPklnR6TVWfV8yGMLu/F8dKjpbw9+zjRRqDK+2u5O3dRotp6
RCVIakbDNRtCZbiezBQX8o/6BVuje55o8RtjYrTXyf/wEsN3YNOC12E1WBERsY33
/jnyADeQZniMO+eamRDT1e0f66wGpm2xxMkVf+CzduLVudyph8QDUaAqx1OC/gR9
dqDaHQc9BjKJOw1hpwEGAJAhTmNtkM/WIHRwKP9mgJuy/1Zlzr/0d94M1gWTT88Y
mSVbNNxpoTr6+FNq8d97upgy/AWXls7L/b13sc3Z0zKheLygYRfeQRHbZCrXMSTq
M8vnSI7NJ8uqDX1E92lddFJTDIQxNjeNPcH0gzwuYuTlh1SPvJ+ue5Hel9R+ehCZ
amEnIYREVpaS4VZ34svMlX9LdiI2zEeBwPjrMPaZwKIUeVthepxQtja3K8efSgOn
3KaoeyV3pNKMbJiIXGuJCTSEPPzvTZWI0H0iggRU2OHYD8gKrM/oDEsL/pDeNHRb
Z6CV7zbmr8A1/fj+RqWdCWFOPMzloqfzAvIPoncx3dDUTjcD7Zsh+9Mn1P3YYUPk
iFQzIZwM7ieG2PaM7MmxcYB7ZdDbaWon3AsJolmwbsCvQ80/j62CUyYOkL2nYaar
3tYVzcGEroDrsEzBHQgkxhjDRPhSI2tbJz3Is9lODDYf1XSkxwTQBtMTrHz3BXCB
Ii4nEgv0Ra/ybmzHkKAumKRnXKVw1EORpe37EJ96mxpOUeU4wVCijWDdtemu2WBP
N8WAhEjKAjmT9mekCIYRRM6FiIZt2C+vOjEricF3rtPEO4impeFz/BG2BQRFYrm4
ToVzoucAwgSCe68UjRemHzxJTiqvjNgKv/GFGdNAADYOx1rGFHuLFA1ZIiEJCDpD
GNgA3hL8YxIEdE+w00HIghV5zUSJRz+2JyOhEvAzbSmyu014kbZNEFTvxRcKcvJJ
SXZ7jQq8aAFzvy+hm+CgvT3BnKagjiclpSRUP5BL1aqgMlxFcrnFP7MWfHfJTEMX
D/tijVcz/me/Vp5aIj1oI6W4DN1r0oZXXTXvk+bddngMYcY7FByjtw0hYjvfr0RD
Ej7BNfJOPZnIn12837aADF1HC2cJZ9q2pfGaHrd/WuBAi79f5wMNafZRZ7bffl8R
TKy9UhmpGBH8lF8bYFeNq4a5aEPtXzPNToumSz5LbEHy7ytC8UfGKaQMYLvOd7w9
ptdvISNfEij7+MAIYYQBVLMmVt29GrgrBMxoAPbjqH8=
`protect END_PROTECTED
