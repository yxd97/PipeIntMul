`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Qw6dMSDiUT0V8w+C7OEWGaSRYXcY/HYbAntg3zgFv1kTCLFzDNdsWiRkuPAbYUv
oVNckVu5mnFl16wfncV+JX58tbfoRxEcm9xopqOl4Hg+Vjfs6F9Nvio//Vnjch0L
PFX44hsV8xV0Ljl1JvJKcGoxMy5489Wy0VdPSuSTwT0PMJHEzw9gr/Qe8ZuJVihZ
HcDzuCNo/lwdgKEDlosBhtmLiwlZnrQZTeGwYTyoH0ZjhKIuKM6HONSIS/qRsTVy
6HbiGWHaUy2iX8N7aGYiv7Ifj0Tr1BtfGcXDUOqgemzbPmxQE1XKec5m6Zcy5CQz
DWgIDIdIqLX8JdFRO4yuEuBvlD9/7VfGql4uCgaL7aICoEhKhGMpGupfge3VYbH2
u6GHmFKpAdXWBJGXMDvOR6nv138NzeNtJZtnaVg13FHv1zzdqbqdeMzZ6NcrXWbE
ORTb4KkleuXi4ca7yikz1p7bOb21P1fhf8FOxyHWV/Du7wE1RYfkZzrvktoGCHnd
fCLOerBwov9gK1glA4Vf+Jt8ocscZMJ2v37dLuUw5rbg9etCX3m3LDYhGkKvAoiF
KYOq7jws8lZ7i2ZY9ptk2SVoOYe/HbcXrtjw6fz0iejKIOPrEixmrN1vnbu6EKne
9Ijg9chNiClGt74RbH8l4FeUg9Z5QD7fwHiadltCo6Ol3el7ZAyLqO2Mil5Kw+M3
yLVB2DfCKXUvcuXI88jPfxS4Ybd4E8ImZLjW2oIYbs1ZR436dEzs9NgbM42bHs+c
dagZKpzVk4g7ZK5q7oUkE06GBPSnt1sQ8kOCkhUsb+FUvaTh6hiyIbkKPCp45LTj
yr3GBW4S8tvV49MjC51B+vWLUXV+IjL6YC3FwU3bwTvEHPt7APeCMJkZt1lDwDmX
Mo/hODm4GMt7mD/vPXAqky1h95kg6TgzQP8yiqRq/i8lquZRvdRIcz1fHJm+Sb5g
cVi/77Sf1PkqVt4TsXEIoZ0tk7EnDPJNttrDkDKWvZ1+KvAQ2qPL4p1D+u4a0GH9
A51AzqeFgHgso1KddbUNlntuIDNZUQwG0mVVVRF3dJzetlzUB1Vl416v3LYbnu1c
bz2XwgaRKsmxpZ7NCc0a7AunsLmV4pKXMBnafAFmPei6Rg3Thlda7fxyJWS4PLV8
1C49/3X3J0EezDgWl6yFBmno9Il2gKr3BTH45/cJuBY/E1pFx/vJ2eT/K5B09Kat
WIqePE8CXfPptM/jlXW+xEiaWjjKccGnAt78iLinemxUcpfL4ncVZx8y1K8N5DzO
Nkeo0TG3mRmNTov1q5QmsKZMq1iH3J5EiJrZvIDYN7ipXi6ipTTO3NopNwtf5laU
44OZYC0QVWqEOfiOE6ps+w23qYO81DlMRhHDbKp+2um14jd7g2DfQHQu5OiMAfUs
ZQtwOlt3VTh+rqPTDp6Yr4F7sgQKLcc5YiqrE+pxeBOLCIdIOqt/lDE8L/ddYIJb
WBhY8MvQJ8j21wskHOZXmL7N1HK+JfT4CFol9WJb5HvSobSIO5ZndNSKe1hbfZDG
ipl38eynEVk/g74CYb6VHxiRvR/yZIHlfZPbdSAU0B+rllclQnEQ3H5FmMklI+2Q
BbO4AAaJQuqdN/kXnBcmgClT2pVL4KbByxYqbLlq7o1/1jz0yeyRtVkqxq8w/t6L
Rx4iuQHcexObwYtCqjA9IXn0tVVDzuBaoOoYOs5oEjWgI8iiKopvi7VXaAM+jsJp
uuuwS+u5SVnoPKQbqGstTSrrhAC7YyBz0I/w0/ynWlaOOgZN+G/yOWA3oUdxz2mI
DMihER4GZZunsUY3Tyta/lrnVU8Y+teCC6Q5oh4Le+6/tMpho48Ca93+mQAn6SYM
MlAOesFg68oqbBU07qrx7mZVSloJFRMCVfdcCHf81CuJOnxsoMnrAPRTJwWG/rAo
vazoywnfZX4HglplFTPlZ1myznAI+KJhUrL3smXGaZIcOjGrxJpcNOtwHNz/SBt1
U4Ly/2pKFTnbgUBHWiuzv8J7nXoMKVNLSMprQsmYChSRGmZEn5xG/9TYxfR5zb/h
D76iTEQAkETYFtE0B76CARbX9WHo0nvCbztqw0uFfZDjbfG1w9JZPBER7PL0m+9Y
1G8wCYWUlVhqBoMVQg+5HztVLYuvpO7q587ubdkdJD0=
`protect END_PROTECTED
