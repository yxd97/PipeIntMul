`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEIRcASVgk7NZeCZJXHG+p/P0pb8M7NLNyGcoofPRyYlfneutE2tEuhqO/lLp0pm
FSaOFaeCj83AKqr4o6QYmXzCc/F7r7k8iyh2Wq2mSGdiUx6DfFgjf0SopeYAZM/0
6G5toLup9CoGVOaYeJNFvFJdHovEsND3Oc8CoeQtT4lCxo8ytm8gDHrO8jrR29SU
udEIpfHpN+F68kK68QnZW0+Tac9p1h+qF1atCJ5uVAApVr1XRyPlxaPi4ndb5mXX
67ioolsI4VRA+aoei4rNS6i7gFWEJRbjeUslPLV/mR3x3zQXMRCyoMURBCZuXI/L
iMDGDNrtyeoZC5tTcL4iTXhu5AIKSWRyafoqUwnmQAkXN6htKco9trTGUddLhNBA
x+1OxgW/llerU9Skx+U1WlmaWUtSxBOtKevkncKOCFuffkwZFgk9gTNTekJuyrL8
E+oM5+p1z2AiSGlR+FkePZrcm5Uzz/yVcw8cN2QNHORxajY2HxXaJ1+bCKv5lo16
7PWPxgnX4ZUPTkpadSowgD/UzqRZjSG7Jry1AyJq5i+A/Ej9us52ue7cFjiDXGCs
SVq2Ul+DW5J+1FsC8wTxC2CC+DOp/t6pz9nNgAk3zNkpquaRD7kL+trCJsO8ztXJ
49EbOK068sQwHLUWEuAhcRCXwSue5IroElzHVQRAWtE=
`protect END_PROTECTED
