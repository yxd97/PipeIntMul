`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eovHhjkivCIg3ZKlJPNqVfkqgtSN+iBMrjetEAd1xxq1KbNrgdFyH1sv2+rW5D2T
u9z/qku5H17FReGJs3VgBJoqXuUpDt54xatjKw7v7rYKuQUtYHmxPOn7VSwZo4ZU
mllFScLxkuNwbzDdiUXP0avWlr++TNFI6KVBc8PSYUHs68ccmb5hY9eDLvd61X5h
A7ElZqTS9q+vfyvNphWu6Cgh3tFTf9HDzrrGkfowarqG/dH7SASAyv/BhtpDbAWT
Xu+4tmyn1yL63QSiUEmnLBCsUEJCgU/EpX7tvYdSNq39BtbTnZQmy362lkvp/GE9
Na3yJ1X1GbWxvCCQIacRlTJlBYEwNkjXCdR8fs6arUGYlpMAaF6B1ZxrGuxHLUMh
VpsymoQy1WADprAx1EujZUj0dSNUzt3VWWEHzTRLnd6IxFZmsEvEaAYhuSReQ15T
TkoAEJhotigxjuryQ6npLGIFnSzjxfGDfoQ3WA5ASEEGVyGfFS+Uzw2GG4vXqJrl
D6kRlCgj91Q/ycyhPErISQ0k+OQKAK/U/2YEw3frvbS2402jxdXTEiykZwX7d2/1
0G47qB+9sIQChk2WKV+SX3M+aSnfPAMzfTq72BMgVS54ILGhLB541KptPyZn0jYq
LcRB8Km0+2f926R9Q4YuI7TZzd980rgoEqwfVnvoOz1dowlDM7axEiklB6Y5SFZM
P5skRg9+CRmGpa48cZt4gApGJUiwuZwdYhO/33+wrqR3iL8qN66oxDIzBgB7Hujg
uX7cE4/1Z3eKkB3oRAExoI8qysAbThofRRyRlWlfNaw/HKsdsYfP2V7YxEeZN7eC
mzcK5rv0FDIbkFx7sZ3oLPYGMYnRU0qkVacxC6IDxIUAz/kzKiSlMBXDO4h8kZkL
9CiaROEEyokbGCOaLEpB0xFiwsSXWglpX2yzgfQNrL0RoEgNcsCUJ8rvolXhxtYj
JClL4QD+gsXGYdLeppqEMFGPFRPukzFw3JPiIYscdwpzHPHATCeDLz6IjBZsau+d
BDF3D3K3mua91WyvIDu5aGhSoZhz1iHniVLvpngaQl5tM6o+R2sMZUF0ij+wYEKG
d36OE87pK5hNoYNNb23aC7iZi9gQvPcs9USMPu0n04seeT51kQ6eKuYsD0I9pkZw
fzLFv+0fnj9+i17kgFZ7Trg3sEYuzebdUsCvFnkbHXGqrhMBVtYW4tbCl4qSWrLn
6BVJB+R17ZJE4NabrRYYmlMgo54/gUracBPT+WmeqDTkLGQwOvGeKnhoizkGq+PU
LQThfAAKfRYjkkEdeJLrrzGZxSujtBLOan3MuS/Jo1GHnk0dwm96k1KV8dAvfZES
c40gnJ+UcjoKVIxByXpJnfDa+qINbvSVFjFCWjZnlefZrn1ucojJyTOOmHY7h8vb
pgqZ4T7wN7m9edaGEPVR0xki3NsuyCHqaSHkLQUe8KE0wdfEJTI1IfW4hoqTJinH
bbxpr+KDl1H+qnVNNQ4OCXWt+3ccC+HvdEC5uATaIrQVNyZ95z6Wj3d7U8qRaDxI
aswzI7GY0xkEPxt2V/sK6bhXVnH+Fp01bSk7/zFI85fyjoCI+iCMX3C0K9vwcqI3
w7/pAQEWbfI9qToAMo3mp63+hiBbDmrS6uAtRWQID8Ah3Tz1oscFP11KapD2eFVf
h5LYyqCFN5hs66V+6kF4Pplfitcai4YLbaaS3WvaQK+yZuChSgojJsaN4Y3we8kc
Ndfr0XX3CXSvIiyFDazct+LyHyCHRlYOOJioBhrLDx/Rr6m6rxkrGmGlRMuDj7AG
aFQZmwV8SBYB4qgJo1Okmz6Riyg5GObiM1NPoEi5U4dLUWVwaRrSaixVyEI9usZv
T8y9pbUKzyzs6NOlK5QdIEhdGQCyKTdbHKIuoS2zEq6pn8svCNMk+FI5Ee/NMVw+
gBhgpBL7gUYgH1lmKo7zRRgi77cOkl3iqaz7S1T0qzX2TKF7NTxuyH1iPwzFmNJa
efhJx7PEjkuntjZdLOF+OizERCoFF/8MRrC0EBjWnSLM7nx841RDUA3ydBDsRV03
b7BOdmlNWExGE2eTJ1RXqO1xOnUI1kAM/LVqyV8/UDuvpO9qXt9cPxohk7aiPDnS
ullcZa9+0dXlEtPRBqXr+bU0t0+24zdmo0nVUfD+r+wc6JWHdFWQB6YPNarc1NtQ
yA3mFOx5pTzaWS8cXyks5xeyM26AvWWeVihHIX3GiIggR+hFUuYEsxNndFIzje0J
aai7ZUIDfSFVilZkI/al7ZnFmyFTwjRkrf3KIlf0aJw78/MwbDdZLU/FGGv6ouM7
FDHDriSEMoENDx+wyx0EU6a80t/pu5Poe+AtMw7hFy5iSBKIE5ATvgmr2e1DvDTW
YhcGOYNUImqr5GYX6G7eA8mcZ/99dVKn+xERqJkdGyuk70ppc4lBhGpRvjOIgeWv
0ooeMSMH8kxlxfkMXG0HXOoApZXdXE2vSgcQFBWmJGHOo4w8SMKbanUY1oFN0OJL
LqTIOhKHtomuE7arRPD/qHhmiMk2EZNSzrISn594qS8yZjh1K0Vw9t18fhRcwwBe
/pDF4psZH4AXO6H9ZCBOu6kIhsZ0MK1vpxa82/Dqc96MB1ZY/1SA5r9p30jwB92N
wBscHBSrwT5A/kRfhvBVvCt3r4wh2ul57FGve+9OEHNLcfYubKQDTrknltX4ncSp
qTEfXc+3l6bHC841TDfQB4ZWcFvQRDAxhMywJgsBlmcpBc7Ah2dPPRklwtG0vFcc
+27+0CGBg4G/LrvzEl5wR+wZqGnikpfcAPORXhpDWR1fijo/e3yg7ZiqOFT//vC3
ARmf99KP3dWXDvAaEm8aUcvn6IXRYOEUk00q4NaCORcMx4Gh0lqg3appd+XeY6Cb
ysQrGRHg5vqAKoJEDxMr3RQ1YnI9fJfNqi6m62/QgceSKBsgGuHmnbeOWRbiuRdo
M28OJr5PpTUyIFre8u0+4XG38HenAg5n9gnuNgzbCKFWI+mB5NR5HQEST0S1UgnJ
5ON7xohk3307ETNzIOQBniM4pgD+f1DckwQS65lXsU2ZIyFxn3dJXY7aJBz5k0tY
dtTUWLA9ru6nDSTpsCDG52VBLlOeqOJj/luObOQjz28UtorU90+Apxghhz9IoqLZ
P6cRryvDy4hjfiWqZYyU26U/ebSoi5TjZ8LxZW5ux12aWI1hcHSgoU/6waLHrHVG
50rZ6LCoLSgqzCKrBK5lUeXh5yzhI9R2ZEklHRhHPsFXt0QZ2VWx3LvCqqdP390R
LEcgQ2F/eFSXFCqwIfOHRQAmBFGLaYP5VG5xnqWo/S42C5z5/3dFFQvJHG13aRqz
467XOB2gwUwqcpnMeDSE2CJVwml6plLuqVTjWOWl0NTLcjhwTBbru9LJm/vGER5b
EcO4JrcTFzn71cCFwo1tbEX+JLtl+bWVny1tuFdUPeh/FCpv7y2doNHNURBPH9oX
PpMCraMXMCacWyETzoAbXYuA2kq4YEyX2oEyAbXOJUtA2U4puQSo6b/bIV8uG0e7
KQ4YyJeFYgoNyqxzbtk56Us0UxFrdOKjd0akULDrA+fIlZrWh8BwnfGoV72Q+64J
EXW/HOIo2F+npkbPODgVe4K7qZ9HCjjImGb3Ezgck9UUwb2mgroFuBVefPDVDDub
iEY3B5IVKfDIC4zoNFLpesEmnguN91lPhaRHsggm110U+t7U2tMt6lmM3c0hcM0A
AvevCofO+mup0P1b/LUIRft4tCCjzXa0288PK7gx2VynpcAlQQQ8gdbxHtn41RNO
2tF1dS64PakjGb4BiVWU+FNaR5RqdrzLdFWMQYwJO2GUWLIA6pV7J+pXEsctqtG/
+ciLbufcBZCRVdKyn3DCXSxcP02+yuHIQV2gBPQKw1jyPL1LiSzU8csEf/mJytd0
1rRELfaESDgJCwTgAINyGvdvCOZIcL434S/0kuHv/HXf95epdD7+7dCrCSrHDG5F
oZaTFPPZFJdxcOfUYEwdE5Bzf/RRJrcOkxBREBK7T6TzkdYgibaz+mLU5whgtOI7
SQk60e20ZEWLmBCib6B6PMwwraKfxo0n0g/CRzsBmCVLYQF0ovZlccEV8Vb731FR
fdLdmri/KmqoGYC4P7zHbjnSha3jHl9zdBiDyQlFJz/fSC0QP+JwM1m1op+X0ExB
g9Njw7yZ/xsBFKLfLe+h2PTE81TXH4Pvh6ErBHxcW6TrN8BLepe5sDIGDCLYERNC
VuOL3Za/ZASszfkl/jyOBY5NpyBj0jL7BkRPA0fyvV5CcLac3PKyKBDeWOkw53h1
QmYUv+vnYpVdUEnuVRFKTkMGD0dxxJayWmSyY8qLKlK2jdqxWYgMNU70NkBQM81y
LAOw3lTAFfVhlRxqLvhngLW8pzIe9h8P99sEXfWKzbrxKu90WOP3VWBq1hSl5Ahr
OZ7TZLElLSAZ0hJVGRcLIO+bLyKNi/Uyly3elJE+VRmht5D+qk3hJBSekn4LY65S
sj6QfRI5+UajPL1l/JaDQyFRdxPqEE5QYlA6AkLsgsJE/jnm7MwqiQHDEBoRDhXv
U/6pFsDGuujVAhRto2woaEPZjC6iJm8mqaarPkQdQ4qwAWU0EHVn0OsT0H7NUtHm
8JpmlK6WJVaP7O52BTyQXD6dSocGlxqckznqi+bI8naCN2WU90xBe1FB4sNhtH0b
ewRyC05ZX6udicO+MgkSMzzYMBoVCpKAeuFs1wUpVTidKfcr5/BI+jU06HAHwnE3
aoM1ca09gNkWTSWVtpQBncUlIekk4cF7EbHSpRnpkfqvD+It1ZH+RGNkugKHjfEL
LShHcR98wxKeYpVnMCRuLMxHANHiLkHRl2Itl8p6V8H5eUg2VhrqY9hpHwgu+MwI
Iu090wWI0CmFjKoaCYBIKV5KpItwRrgSIE2D5URIX8WGAuojJIoTgQ8hsJuSYbvV
uahTaGZo3D3fq2NDov4cwdhWLknXIvukUoY4bpGkIiprhCahFKfGPeeGK2rw7td3
lrjmhz4peMEf2Y0KrZIOrg5Wyf8Va3KTTCieckq3TOAb4vWgBQy54xz5Db/DP2rI
zp42NPIHN5qH6+Af69PoFxagt7XUxnu1OdFON1pUC2DP2aOCSp5UDt10GCwNrmOb
Z1MUM7CIOKz6zEm47YUz0MtN/q4hCxn+VRlL6zDGmqh/h31ivcEXJTNsud9TUWCz
fH8otcvdKSr48LwqCHfkFJpP1n76GMjkwdjHTo0iiC+MKGJKhhpsaiYmQb8zj9If
diI4Z043nxodPZnfkHo0R5cQV2eTy6Y1Zt+JIdH+z89R3DhUyVVfWdK/pIBbfqLZ
8y7nOwPuEOGOhVyJefyW0KZVRu+cUB7kWT1PQcOvUkS3/tOc9RFNGl8y3erT5oUZ
rUt/THOT1Jhjh9liYKjQy7W3Y7ETL5GplJMrN2R6LauMQHSL97aLJ+TDJXe1AUH2
X3LBRWUjnbEoeQKenNcXgFPGlKvcr0WTHSUQNpCrnDwKdqPZHGbAb36/xHUiagRE
gAw7U+eA+F2QOvZQQTJ7hWEaopNeeu+bNwFDfAhAlpQRUgYAewMKnTN6Ks8WMo67
3AHq3uNlHYK6HhtioNKrhY+DbyvzQUVFg5xARFWrjrIBMbBjnsEf+SYjXkEghJ38
jkEzXIlVZWN3OA6p7aVd3ANBhkC0kM8fMepH3UR0a1zTFHLpO9kCxIei5lsCtWI3
QeF3YOQd3r2n329f4SvUD+tx0eXEhio/idZjw78e8Cvty1+82BEBZ8locdf8uRSl
JlhAMOw//+U4h74hlkacFB4E5nY+NTmxA9cNAS3ciUoqTOxBQeyk46fodVVx+DdZ
+A93a9RtOLqeDzVC8p8qV49ivH2ho2P/rc3HZjGZVoiD2PZN7liYajdSK3pFEv6u
N+Xd8JDtk/qcSXkfhFHygD1RqS9I9mMdIGgp4j+hJoHXPTRugt244D882oR39H1/
Jpd5SLU8Jx1qOMyv5cUlvxK46Vqdmc0Bl07W2UPRRnK/SeakFJF/K100477z1mIW
4qIOOVxoxQV5japTUaoIgiCw6S0+BtAystrGuiM5xHJT36uUlEKDuKDAXL5juc49
GH0CqsQa1RbEip9aqWCqmgSczqArzztKR8I62AT4lW+HeOYdcTwrey/uxeutWY1X
6khAN8lMDEpwVyrab3mi4gRAZypvDtQ2GWEGE26nnBWJGyhzM3tEs1A3fP0Dgtd/
MlC0VyVOrD016KhT4yhmHIh05lAi7cFOiZVbNU9VtIOliQTjBNcDJtdei9tQ0HxH
ugPLeSUT0jFMBUGFqRJZXHbrjRAklzufxPJx9JDng0R6xs/jXvNFU2j0mX5w4Dn9
PFr/6LOrjgDzrcg6xQPCn/Ckzms++eymRCWp1Jrg/xZjvKsvkoLMgKjj/dbIJxJv
73az1nOhPe7vMLio1BRL4pKldW9yz5pzaeGOzaLGNpgUQD4obOOpIebwe3PY7wlz
8ZrkWVyD3qrGy2BU5o4DA77LLMVnPQOeKOT+eFRGWndTu1V9gOKijAq1LZjWkyHk
zI+6PUhUHARnj3R4Zz2aloh7qMu53g4Og900MMaOJelbOtn3OFIZFTYtdeAXpfvf
9OyQ87D2rI4NFePNiuy+nHktUm6TQwL1EU4DU75+HuSFhIyZQT0qkyqy8Dzzz7bH
617y8wsm+tZLsxVSQrbxbUZTL7b2mLcuAk0JSuQMd/givY1IQtCATPpjL9rrHxg0
7Zqco+sSF6eVy7G62TCMKkJM88LTce7s8XRJlkSuBqpGTG5pelM+8ZPZbvxdUYkz
uiv42YaO6wF1rt9gg+9YCfEhRdzHhnH1qNKQCMG+Om8IHUKbA+LjVV4CrYyyJDoj
wtdMWd6PR+vEZYillwemoqB1PjbwzqUIhNUQ9Wr6Vg8yeXRabeytHykvwOyK8lYs
VyirQwLaUXfvzfGO7duxkO4muqsOJX4ilHX66H9cMaYKzkFAV4GV/xwTU5ZOC4Qn
jutBi4KDSLfSrTRPeI6t6g92tql3nYWT+MFfv5ug/QMvynmobul6pO7f0Z415240
swPYFYZjuyMrctM3kAv3zz+qXmozjrN0dvluD0+rDgCWXyzcYk+BGPVWjeYhVs6C
NGy9QJR1d6pqKKvl8C1iGWO48/D6C/hp8r4MRXLb8s8NeHTBF3HE73M6hEiPNfP0
ePRcLnIrmioN+rKLQSI6OnUx7MpNZUVGBb6o9VR0O2e+W0jOdv8GnNUf3+zvbPH7
Gp0EOnXzHUrEgjUSrZLUZWTF7rfKg9H1XxINMeWtioys0zh+euayLURTOsb1zyGD
14a+4RuYgHeg6OSXRsf2sudfOyTosSTSErQIFdXS+xLe/N/4SV69CIwCSnXBiixi
JrBA/70AMJJyM3rPop5+SSij3lKyXYr7jepKIpc0ABZPJUOqK0c0gG2KXw2u+Q7K
z8zWWOWlGejr+U65+n2bBqFIe1S7y+pJLRxiRkjREiQ9D/HysPy87YFn5uL0o7Zz
1A0sPXwNE8R0MWdSx4CUkB3HOHvcTM40sg5exQgfbJGZE5GffX9OHkEKRcepdjWL
CDbTAbxEz9IJqi6jLoWld2p/3OXbbSnpjHp2KsDKXTE8X0L8XCV5l+ssugZJP3T2
6uuIX1KCUwBIJYQ5rXmFJZx0gREVWgsn2xeZRZEr6i0/8hPOquLRl2dUmtzhFKTJ
bN6B5YJcQ33bZy9KyXbYZbOqovUJJ+p0X7meGaze4CDBAfWx3C8IFiqyaDMNSxrJ
Lol/EBNVIKcc6R9F8P0iGVeL/ZmuahZrxIJTolnszKyfCHI591UQx0fhDx0sKJmK
Z91OgHjJ7dRUV4n1Z9/CP6PgRfhKQUoLaUUIpHzydLn9PXNg4gKeZgJUf0OBa9UO
hVjhdNhn/V8D3FyaxAifNhof+wBzuFI/xaaAW7BVO5iHsEZV0Az7fEYV9i6fAGmi
EDjyxJmRTVCqFc1sw/I8u25iLsDORbIAU0IAFNd09lZXzh/OisND9+apMb0uL1NI
rnBtzkk00+naC3UB08fzofqgZvsbo/4lNnG+wa9yq0/nMhdmJteMqbimyBPgGVtE
BTEDkEJIZ3XHj2o0l8EVFxtO8K9aUFYEIvsBT4QAYQ2UjAB6h8boun/8qWEY4OF6
CtaEjc4JKD28OsymW0GQR2EfCNOsMxGpXuMZqaUjOJ6CVzvC3EfIDsU4gL5oxAR5
uKGx11MslN7uXHD7BJhjSA5XmrmlsrH/Qv7JAFTXUhpzeJYiVs7C3vP+y91FnKih
2tHAwTUm23beCfGZlINH5GUk3deeXRWovkLrLYOjMNAH1KkuhP3NfnyYE2YybTLX
QMKAVugRdQ1hGUzmptdz8QtXwyP8x4k+czy5eZd1OeJmd/MZacArHA1RXxtEMmag
cj4Ph5PiKufoT0QkhU+t/V6uN5ZDx3u9TaAwl2Ep1hFIcgz3uSD3mw0OtJ6J1NBx
7qTqU57wq7FIEEflWM67siNHJaOKM/YRBw5aZSJSp17YO5j/uhxGRzpneg12ZuUd
7mVao3vo8t/IXzxxIkEw94hiFnZqI2w84GjybNFW9OEC9xy3t798hMIBRQQs7RHK
TnrxI6VKz3vfzDzX4FH4yRPt+nhRG/Z5KX/J9VxKMIRaS+2DVKc0BkDT+6kIxAFv
lQqGy7FYuKg11RJ9+jVRKo55fVTbaDIhaXkqDcJeRuiJGfGEb689iLbDdEOCSG7L
3MyGtPDupm1S3N9OHAYk0G7s34TCzKrqUMP2LT4isFuzImnAWMBqVZ084hBGtkxk
9zWwdupWorqAoYCDu2pG4Yx/CALXpYEL5cBS0kmV+xLvEGF/ZrAcmaKQ+pGMwyJd
lh9nuzfU8QuC2H2mHHot21YrA71f0I6xv76ryG6Vuf0H5UnYotuYFSMDKqt9DZNK
4XQVRKcDaNFw7Wu82Krv49eb3kr4luNHNDcnragVE+CR8skc3RDropwryQdTOs0U
oteRO49SnLn2lFQovLcleZ1zPU9WrdRrRGJuF4f0nmqQ9pHZMcoa+iqzCylNJA6y
tcI7ufI3GbqWH6C5VlXlxAXODTUNNyWRXpkU3R5FpcWLX+NtUAB15IcXfdbzGK49
aOjbjM7z9NlC0l7tp3R+JVP6hwXntc1+oZI7oqFhhkYgGJff3TbwdXNW97prSYli
nt+8pJd3SFNeMZmQQyImtqetK3cVtC/pktRxApZQ93hqjUVfaxy+cihvU4G/jDrS
bbxB45szxvYPrRl4onvtjMAD+Ln+97S9hRmSNwmkjxIUKY5x8xsh5Bt4Zs7njafV
kQA+h3f+qnAPrpMSztAA/UH/1iiBCVfRQTIHbrM4bXY73ra/R8E2qpDR/sAe5lJk
jP+JSy4GVLTSMMcxB9K6WoXYZVExjlnOzNAp7Cet+uhIAx9ejDZ+w7nDutdMVxS1
HcZ5qvTDfdyCKTh3wyoSu4UKIoeP1iGhYOeofCZIeP5hAmcEizQdSfImh0hJqmoa
2fT1QsHIvoe/+ZlANsRcOtsbRSmpx9f9KdNyCi1FX02VtAMvC8YoSdJr/rbnXaqG
cBBTVqwj1vHGfKA5P0b7uMi5llsrKOpvjrDnzxKJdP7ykac9cMHC0B+7J1y9Ifvy
AmTtEFUiUAq0tNiJ/m9BadmLPpzAxuFxpwXulE7w7wRiOD6mdjnOiAA/PDkUromn
JK51PUTSHPQbzU4Of1qgSG7uMdyvV/hWse68LvH4sB64NznGGGMvW8aM0RbytTmL
Rmuo4N0w+asJgnfQ60BO4p3y111f4MmowgrFzXrLQvT9JYoIG30s5Zdo4iBhAV9p
XMWF0kWLLAplgY1PRMkOfupKQUUJyob8+yj9ezCkWu022frc7GJEpmYd2dKOqmTC
65vBttdlV36Kmq6yPjN3eqJeLT3PkuYL3Tm0Lz9VVpp62c8nmf/Uy1hL1lVNTtvF
DrOTI/RmjQPKhvH4hka8ftJI826GhYSLxk8Vya/kN7OTh471hw1cOIIHcQvV3r6/
dRi5Dh/jq5ZJRxPR7+8JSEDscn5x2iPET7dD6MjjuN6obgiVcC78vXq3zZnvHORr
3Fl1hU5tnN01rbVow7E/G8RIzyOKfPPfvhvWD05Y2m6icq5bj6SMPvzqDOIhXSm9
olqTTHCGq71k8CflAlpERVn03DPCrWXYp5qorY95DKDHdNS+WaIfHsZ01f1NlEZq
GlYLXtXS09s7NK83wqizTH198267tcBldpyZYyNGmKUlkssaEDoHEkHCBLfyqWRE
01DPAyZsx9yjXR9RqeBm/ztNsIzCu5QSvmsT5T7ZDzhzEVG8qWtKDsPF6opBcEjV
nqlYGiRW8pzSgZWIKOKs4kLTFZZnH8oaqAO0yU/EdA/MGIeHFGVvDkSrnbdCzGY2
PAIBfQ8a61XomA53k3z1zQ4PFx9tutxX1rVZcC70oQMh+gWFJ2DR0kT+8jEXaimy
2zskri+jt5r9MLAp/5nDhz/2z3/VpjcHDm29N1Y1Cm3yidufse5yoOuo+oft7+xa
UYhizcX4Xl0Wl0Knp0C3LGShvhrTvsj9FwjgzaVu2e5MTR3eeiT46uXhdaizi/7r
589iqKd0kqdhhh+r9Dd1XVQ9E1Ar+kYxo7r+BJo8c5yWYr7JGeknyRxXky7N9qNz
ahnAcXE3VZtiRDawyXMfbp2mgUprxEd1SNO2pmtvFcm+6oKHe4EAV1eWG/tNnXn/
7unrPR38putm5D2Z0EUaCECY0DkDDJ6ZAsE/yC3bl291Fo/oHB2kfAF7lsu7d3lF
UdZNSIBFeN7COBcG61hgXCH7rElmyatv3W532ywenwEVoGQRGFaxNGZOCwpdxlAf
Yr/t5GOXXBQS0yQQ9Crnxnqwsu/HCmysKZgJZtVY05fiWpObPPdpVpWfhPCavQkJ
nhDzcfN0rc2kepYD9sheLW7Cqh/+ehTu60UiEbDsn1vyDF/NuJAjE5iWHwou5dYj
yto4SUT/OwOccwte+rJoEvIS6EQqn5r8rYoYzkRZ9Eh4/Q5geXvCPHxYoCtYYR8+
B8cOKzQpEwCpqABNosJADzA4c7nljPJ33XfFKkG2NGYaHTqV4lAUAYrL5/Tdj3L/
3VzVVh0/19UuS249A9L2EW8x6+jvvuIT5Y5h7DkuE0P8Uki42jtV25V62QBbK/FJ
0WTxt1yYzq/Ifekh/0STiVgziWa+GIHPMqdozWHFYquAWBFsV7n6XUUwC/bnmxR9
MP4zqkXR8W+L9NvfStE+CC3SE+XBFq8wvi6VQAn5ETJr4zWGcVh78f182/9lt38w
5VwjbM9X9hljeTI53+mQy/nbq1sa44G3rxm3mq3Xs2xpWzEUr+ACPrc9NrADuOIc
aKaj8HqNAcHLhY2SEfE1gAy4D0BXve3T6s4DLQMbxTjs7Ie5CNVZVQQE2xdvjaMH
DAAUilozM5/4hXZHjmWHvjFfNEsZa9Dd5F8n/+uS3JYsHxymq6q+r0gckiX4O637
WcMOqkJ5DAGqofwvSI/usbnfiiPjiydQF54uFtj8vj8Bi7b7taOLXNtFxB5C63RG
E6kJ7kpVf9zyaRZ9CBNJZ2kLr8X84OKnSaPOCAg+nFLOASZn1hzoESLpZlBAvgt5
2h8X3zXt20ThMrkvpvsFAVBzBO2MR0esLtMvNMDCq0UHyWuh1Rw2+0bWe82G7Jm/
/8rNUneNEvcxut5xYIVpUyvZzafMhWcAOoGQJ8I1+S124gdM8qHpPHXtxYvv+uSb
WmNFZG3u5oMHeNtgIBUPjA==
`protect END_PROTECTED
