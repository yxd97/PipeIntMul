`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J24sYKlaX3QpZwLFL9/+yrMc0ZWVS3xaAVmG9t2QCF7lk0jloiKpkjjUGxK8+Uuq
uNc31YngbDgtkPzB0EOw/Tboaq8bGRiGnc+sv7KB7cKRwNnpkFfWLIuynl3fTpT9
Tcj3bbG9pYlBSCu1StF0RR+/uQZmLMFmSeENFgvhGtK/gNDBxedpfkydUjGT2+1s
TY1PxNbfQL2ZP+PPsCIwNvVYvOXD6bHfBhMZh2Sgev0NGIuDop7JJOuGgbdjA/kd
08Me+cEYLl2oHeacCUVzrHreFMfsZaIPwU7+27O8H+tGW2C8FN9RSzBhhe/BcfpX
Hj01cLLv2PzZ4YMZ8bp3Lx+38SPnEeVhN5LKvwbUXzvHwVsj5vquSVIJDzsL2yL9
JUqHIg2BOFNnzoFfV71qdUE1nefXbTk9dHTjG8B4BnTey9K40XSqOmF+ZxEGX9tu
ZpzKCtv43BW75wICRqWvTLCVphl4Lu3EyuRpQ/A6RulwlndxbKfuaEDzapAWRsFh
DRpMg3aORs4HOGw2QAM2FxJOYMUWV15ZE9AWjBBe1UnBDbJFiQFUcShBjzmuR/++
gMQq1SvZxE7cDgJKtwUHOGrRlj6mH+QwOB8slXuyhoLu11sCrtX4i8p4AENoamj3
DUuufD4X8MAd+9PnGr8r2LqsqnoXE43YkUnX7w4ebV+nxuIWvjY/x8nh+vOZI9x+
fHFrjEO0gjuK7/Dmw7M3RJXUhmRgyPLPXLgrPJO97ePkMKuGnYDmdH3bSKKtkrqJ
WpOTcYix9htFLCHabnx9YuZ17M/rOoZV09uSEpz7vN1MDkYvPJZJ3giC10sJkA9i
uOkbHk74vQQXm0dDLnHpEK+ve5oJSqIlHYVq8ByT4k4eYqOUuZUGi1OEXOX6smc7
S9P1mItk2vbeXqGVxkFbDWehEBboiO5ZPaDAA120tWW9dTZz/vauFWx2J6ge43NP
/G6gBQDklnJ9PH9PooZxEV+yFByvVkzmEPYILJzigzQPBg8NnpYVb8gOcaklul2o
rhrhMUMa5lxH9lCaUXhovWkoydOPFzv/VAGrszPYRoihldA4b9eZVurdiKDD7OcQ
E8cNK4C41NZfOxSKw1Flwd8+6wOYaO7K2te5usGVgXVVqqCN5xYSPW67HxnskIDc
Mgb8gitkozOwJvsD4m8QcbFtHDQIuAnnvcwbUXaJXcqqkhbWdBBfVnImruWbqLrR
1u+u8AZ8kaV92kPUegcMi0L1+5RZPVMebV2lec8h6EHKqdSuDUO+55cdsIiLMPYs
5IGQ7uKc2q5D5rRBeKGGsgboH66rCO3n0D1m4vHjnZmNelQc81rB0kSzIKOiWQzH
mNuJwwJfECzevpem1sC/9KvfDNYMCKmiwHxAcpu5yo6SyYKI2Fj7p1JGroediVxe
ER2ROVy5gWEF/8VqH9adH2WIrCNOTgPzxKEi58Zot5RrazgQ5P6VEQ3Tt7U3LLnQ
O1h9n1vrlecqK2yyeoVbONurR3jd0JvQZiueINCJrSSnAy6hFyM1kWn9dqcGCJvc
tKM+gFtY61wOpnZns6FB1TTQJvyHktfIkVzKKotYD0b6Ib6Xvh4rI8zNyf3Twoxz
PhFW/OqVmqutZ36tU7W80fGSVFxkAye6FuIaU0N42ErW++jAQULPcIsiLR4MQeDe
dk81k1o0N32JPT+Eei56xDtn4Br+ws7hlp7ZRqYyirJPZNxFNMrf8R+93OxuuTXa
RAd/IXJ01uunfMSuQmyplbfbRz8yoIP3hXsl9dxoZDHOMUQ2ppFkdKbLUb0Ro9hj
yCU9vCFYdMpF/RHPxcRP9EvCRE8mLm8iwGRoNGgQo5/feTAGU/zED8sczOseRv4A
mPVPQXXl8Mq9B9d9O1u3Jjgxe4O9XZlN4tK8++BuWN+fvcj+RaPGgzaihQUEeY8i
gf3V0w+YydPM+dWUhvgdyRYnF6dSnYxnKmMjuFqN9fe1uIFmdPlqxSBvDhv48Psp
kRxQu0930ArCv5c0f69kyAFEA2iYxEKcnYhQFd0AlMEzYT4KHZ2Kcrz+3oE/jROG
+3/e4toFFpdEU5wmR59JKsVNaFXO37VUmvg29EDj7ZZQPJiHj5Je9xDYIYsgQ3Kn
51TpZ/lAfyWOGBYf1VX4r2RMdugfoMlxTS/ajqxeaoZjPKG2o2h+1oXfPSJEBBSM
zN3+Ptr5GZJ7xaztReOi2Tpqbjj3XwKdfWar/B6xz6s=
`protect END_PROTECTED
