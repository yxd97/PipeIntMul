`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
03lzFgtmz6rQmtBNVxbwAeojSqgOAwgQtrtmfe5be+zBcyiDb/gG0SyTRmVtlZyR
xK1tyAeQeWm2BPazrwSSYBXABBvlH3vpsbn9E4JjaXA3yoKLyw9h/sgwpDtJgusS
M/jkm+i/frNspTDstITOaD2kEvYJgSkHBhY9+oT2JCICiOWyAAoFxEMjlYm6EyRb
mmiZijJwx9v0RW119ELYVJk+HSc4sZpEHCE+p/FSKcO8bjrxMlLg+ePOnodO4fhF
iz9OYgrUyGZc7+VOksS/4A5PjPIKVyHwDDEMBWauyyqywo0QUxp/ZBYXUKS1aPzG
YP4U95FRaFMq8bjE4bxm4WAUcit7hc35Hb6JljNk1ByTp8UFwv9hP09EADG0eHp2
1vKnRUtw3oJIVaj+QTq8uLmQo9PGijBus7Lo515gPAR83IWFjKz7+I7R7UKDK7lc
P1S27OHH1OAdqt76CWHj2xE5l/+kgNE/pPY3fQA6bCcKQ2XUa5KQX8oT7QPr04Rz
cB8A4ZPScmlsjzHZ027g9KrKHFST5qPSH6dcHk6bQ1AGF2FpN6VDcYa6hwq+3uMG
a186let3BHYxxdUJE5Rqo6BAJwtKKUDtRtUN03Ok4ThZxFDeYeEVBjXcQ2njw+kQ
0EyOwqzpFgwKSTD+xqDLR7vJQlrgR7HUpEEzQgJF5z+WbvdpZXCzPgPRxkSY+MSP
Ax7TalGXa/UiZn+o/+pKHMS0x0lFlyUXgiQ66lAXg/c/NCA0jZviX6UAQGtbNdND
Xon/XeSYIvBWLK9RS8md3W1O2YMnCHlm2ScAoyRNaDoTXdoTKRJngFNXkbhwQxxN
LXECO9pxF+Ln+JQXxiV6Zv68GYFkx6zee/TMC3Z1JQVKnI77dINFUlwmPkxGpQSW
iRDTtHLlmmlrKFraMMk9FdFM48RVtO4eDlCPonbcfTY=
`protect END_PROTECTED
