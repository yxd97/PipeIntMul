`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PjtTbCfdvLmaHvAWcslgaYBz6W7Ue4Z+PtpZ93GBEgcdk1KkbT+LFn7u1igT0rj
7WA7vzb/Q1gmVi4hkKfpVOd1v3+Jn4UQRxVMGD3ZfHLqbtmU6rzR8L3YF4jII48e
pkSfrjFHrrIN/svOJ7Z1mM4pAiZFxT0NCRePS2D0c/inyq3ouC28x1jX1uFzpCib
dLpUPpmbaA1ZnljPv20cEQ2rLw4FofgMWk4+oYvbf6JqSSHUr4dyjdTdMixp6ktI
VxL2ilD7C2XcjCys3sFr8IbtrWr33gxqikkfucTa6hawlXNv/6YJvilwk1DTtGW8
JaICteHPOa5mJRFNnCu8CZhyvBQkS21h2YjQ2ojHmxdufI/pRwxcuKaOn44xG1/Y
ASWFUGUiVumViuo7dFcjQhJX6xuZCgCHPj8uC1Sjy5/Z4gN2tt//odOIn6MjzXkG
PLcAJjbaVqGc+EdXq230y0VVnwiZ31j1Ab8eOb/6Vyeo5xQ3jHnNQ93qUHBSDAge
sAdXsvf4c27QJhGOq09mcsOnUvoiRoK1YX5vjiqmARIhK24jcDBGcFWQvhJWIERT
A6P4oGEmiqLETDQLWcNtukdtX3x7YQJy5XNH3P8C4LHW1y+o2yNg1gih4m8uaZpt
zRYCI7btReWkr1PUejxZrhAAxcQCt4P1yJOJfj4b4vjbGKNoAnSDHMxSgEfMlZv9
AJe0h/2eTnN64aL5XCx/QEzeS98paapWcjWcIzr2GEQs5Q+Q5+082d6SIXgk3zFi
ER04oQALoYvk7Rfh+jmTZNDsT2Y7iB+LCl/4vhfcWpmlXDzX5FwZztiuMKSSdgPJ
we/Ipr3N04XECIXX9B3SRnkr+GmJN1WXNkBLhm6vaPiW4MME9v4TKBDsERLjxW6u
aZ8WExYFbSKaUH43MMXYbegItdlGZ07/B7LLWJky9o7gP5ArzH9YXGc3jJMUwvF4
a/q0ABBpDyqCMBwsQH8iiTgAdZF+BVdBtE2vkphCZypx9iFQMRTJVwAa9cLN05mN
IDdqKS2o90mkiFHTdoRMEg==
`protect END_PROTECTED
