`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dXw8W/0aCWjLiSNrjYWNW+AkGgc914X/mBKOUvJNNFnHJafFtuxrue6hDT7D/tGs
9bNWB+WIGaaJXGyZgLBWDCi3u4HfpxNTZaMfQQEZJHSKID53xpL+QzpK6kvwu97y
QzEG3V0Djc4qdiYQyE6YQCdDW/rygONoOFclE15za7T9c6Wv7diffqghzKRqB1MH
adVP9Hr4WZR8H9qsEohlfxQ8TntCRNPgdms77yAuzyRreQRuZb4mwwgWoICUBjy4
jBEfhr3rB5fYTh/mCi/ccCztr0z0dbJGZa1bQRaroAwmrprpQ2exrDurxNDpuWfg
dah8PShchAp4qShXgZh++Q==
`protect END_PROTECTED
