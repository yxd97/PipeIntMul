`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QrrB9xufUIERXMwfO8vd7itfdsAt3WVjc69mGmqAbDY6Uq6h6wIJ3H3C2jSuF4SQ
ol8leDIMeBMZd+9eLlHNRoKYIV4oGCxbwjrr0Z+wRVQW8klpMU7w+oNFcIy/MReg
VsDLSeIpRrXcqfsRIeYV8a0r1FW/UEz1X+EG+EsiO2RXlmtwctZ8J/Cb2BJX/8zi
TqqmfXJ2ZoDOnnWo/kXBW+0WsfqDg5F5PfcvRk6b9URrv6+EozUtFuKEGT5cq9tb
dvyANH2cygALrnHr8MX4S2GW1+F0kwfF5SQOXJCJ2/rG1XiBhA6J7LV34gNCqiIO
QBKmPJ/25wFppemAeJYLQFypmZuBoHWsinaG4WCv17nwWltMUm166J5ZQxRf9s+a
4oAfHLIeR4wkrObcAi9oZQDvy3Vys8avgtzgdvQYN59/BiZ73aFujuKvxA3YH/8V
ZTffm8ZKwjSbdpSkvY+3dI0uUu+gsqruU/GHYp8mekI1Ohl4vgm7Fn32q7kfBI/+
F/ryEH9yEpsVvctJ8zTqVU+CsbtVqgY6j0jEQQy4QbOaEI+jiTxu2IVpI7zyVi6b
`protect END_PROTECTED
