`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9rsItPlJTcUfFhD24PtrnaU67FmrtNkEuQBqCOWgZC9hKi4TnSR0v6W2p1uskku
CXvqtSG7T41x2Zk+o/hSA7WmShlXqCIoFrRSbhuBk0nynps1YD/un1su8JxVKsFv
x1MDjF0gCVOP867SM5nBw5qip2VvT4E86d6fb6iee2oQRctQegA/zc1pSCeqlVLW
AO+0z1VCQfrR70VdymTkNg4iexSooK2tzx486+UwvdSSBdR3HvfsNMNgj19C2tu6
kCfYdt1KSMIRKbpe173xSo8rYHTf0z2j5QwpEpek0v7L1V4eIRnXULbxVBTb0bEh
CJxmoNoy5APDOQJlkS8PPgR2IJIU1swFbKvI7b1VeZTGtyA9/tfNIyT8qFR6GUIA
P7LYzIvs72EyNI9VWLDpNaMYd8OmRwcH1AvbTxFnmuJ9DGQv5kvCKHSnYJY+0L01
`protect END_PROTECTED
