`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gg1puX+p4HeSY51UcsGLstNyGDt6ZRw4sp2VzqoxPHZfycWme9nXD8e2IRop8iPT
4G2wniL/L3su7kYmIkqzoen6jEQXP9f+ZhwVtU7CkpInJtV9EBnboIRT8SL2TCdF
J9ydE2Sx7dxUfN+eaS/YR4+ZgMS5typ7RT9UgxwZ/7sCgvZsLY5ZY0JPjd5BYOtN
YJx2jBFlwOh6EHT5kFPfcy6BWhI9MYwQmuNojFiMZ9gHM3tjCFkqYm3Or8CqKGbi
`protect END_PROTECTED
