`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aS4Q6AzZA3+qTLoj6Ono57bnTGCnwkZRZhl30o6p3BU2u1B6b0i86T5SuKwhpT5J
/21VUlkFNE2RXlZGKCVqZ1eTVv5NmBhmjd6BKomiyYXz90SyUPNQq5hDdmQnZTyJ
NJUIQAuyd6jlYZtytTeyAHpdfTOVzgWgAJMuQNnEWlgNVYGyt47E09Z6S0IxSXKP
9QJCuSsdbCxJaiGArbxQcZF2iTcz2lmYm6JuYH5XB2yIB643BLm8UglzQhGcdmgI
CdYARs5jDnN9dMo/Sevq4+DEFZdj+KftXqI10vf+RMaHdLo+PFnwbHEkC+h8GH3g
q73Awy0hbvcH4UTF991vzB5l3N+4eCI4E8LyOSD8Vv03aR3DSfrdElCYllNNvQb8
28P6R+HIz7014COxlw5+Bm1crZVbuAn/wSR2j/byYjnxGE4sQ69pTRjcRlWlg2GQ
spY1msZtJt+S3VJhLrStHjoP5hNix/kDeDsYJws3RL1DS2DDUpFUwMm94O9uQQf9
nsdtM933EQQ+3z0+tHABD3xKPtESN8OZopo1nKUkxW3wZj89Dat80iuf9oa/C/FT
xmyoiBeS543QZnJwbnwODaAXr82xXhWpj0sOxHWHvDgZVHsNJs4Kk3/ZGisaWx6n
Cysjal6k8pNs8ll6paTLK6Y3enxFXqZlEnwR1QVkeVneFYWZb6mZkYgzh8060HZ0
EV5/Wj5OibZ2foNuKolEVJN3AYDtOGgxnC37RuXA6hSGfwlp9j44sTVtU98YWchg
SMZK2m7eeeU3ciwyCwA6ITFj7KbUVCQssuXxzwdqSTgOe9nJeiSL4RvSs88V12qC
kWh1arPe6K5XooeCDZTkl/XbZ7OvVYGV0VASXqoNr0k5TrmgWNRew2znfUpMmUXp
eInIoJWqSeU74fze1IlQZpJaeA1L4lybSGeKKAFwhF5pVsNxd1+qNoyHxfqKxQZG
x3kKNyiXU+dIMdxXt94A4VSP+w0FdU4UvmTWaC4JRbXPYCahH4hai6aQiUmthSsI
`protect END_PROTECTED
