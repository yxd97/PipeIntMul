`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pt1l5RUkauUq0c5iiFG6w+cU+ly2B7eOqNLjzU0vNGmSXKY3/4Waod/P7+11imB
FiNrDG7CWdu3UPuwZxMbSAwglJNgXYqVsC6D2ZJ3VHcMZ3r1w3EFn7LDByUqg1vT
t7r6n3gTGq3/BR+7Myb/X+wfgClsQvF8MYDtsA9B8HwS0NZqrS9CyfD5zRbsXv8f
mdNwc6THYebUAdZK54GsmbwK2lEahOmXreuQXMSDw9GiT6lT9Kbs37PMGyLvQbEE
6M9TWOUASA6goY/5dtV77V1us4ks+rLlMtWVqJe67KEcxbO6v58CymfzwJ52Q84c
Io0FBOQXDRepCPzbzIeCuA==
`protect END_PROTECTED
