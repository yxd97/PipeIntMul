`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGqXDvzTGXOLptXvgmMCiVO1/WkkWQtqTytqfHhLwNv7liBUzR0asaqeDQ/pVtgl
gkajbYf+LV49RSn+Js4ayKOi3HNBHjBD7yGfj+kDCZKleub6JBc9baZVmyFvO7th
raWuklfa5//7Ln4SF8UoMB6XtYz6g+/6f8yKC+q0Dy0AlwTds7V7f1qy6vsbWXe7
ZAPLln59JoL+o2Nsi7xj1L4fhxdYsX5BAUI3u//Q/Yk9szh18UqqqkmkYT01Uu9L
epSFylNw9l7V9xbOFC5UNZ2oIijgr9DCPmPpFdjikRqngO6Td/nVCRESpcx/cCZf
JQ2l3sbFb0rXbc5UdIlUx0wrZqTdJfHNw9lji/oWS5dNizbEnY8I/adE9WG5luZY
oyFdXRSQi5m36nILFJwN7N0UC0uHqgChPJielWeTTTpKVp2efBWVSH7rZWBvnnGU
JWxRanlr6e/pZOIiF8aJt25aBwnVg3KRNUCS/2d+ItdAmhDaiM8Vn2w2eCzPwUrW
7PUq1pcUE3eHLLzWo2bo7/1Qe5JrBgzJvHoxh0Ic/Hm2J0RwXNkgLSqcr3z9Ja4J
KVu5x/d2AtUWiIiUVm8yeYdJktonBmxbUIXDunuiOwiheEdXAjpnfZ+O5YhJGOoz
Nskyg8ZOnurrdYuczyFiLEU7+0ixfvIwa3a0yMGLpcwCLhoPfK7O4neWCpv8WmrI
Z7ESeeJCV+SA5bfjEomBE4Z7Y0Ne2vm16pjj9eQmhd4EMnxOQ4kUH2Ri/OQm6xUf
cjFRFhVQcnjItEGI1cl3cAofh6WPxupZOgYV2wYI50m5ugqmDw0ZGIuq46mlpsOn
C8E6LLqEdXLq7kytOOGLQHzqqpjqpUjS88Y5JBwEoKgJBkNqqmQgiYKf6fSswXjm
V0NQmUyLla+oYpTZ2gnGi7SAlStYYUueHk40xcHDgKXOlux0bGUQ1uSAthPHsDTd
W9wPripkTw9hciGVrP+Im1g2Cs7h7kLTNMrQDAirIieVrFBEnrB2PGh6BUNrBeCZ
54UTCatNv0cWA/e/cqs/iziM3hJWeONwxvSE/xgqks1MNbLTDohfqhChCXdPqJvM
gJTLzykGocWavCxd0znTbiYVnHxr9enh2J/JXYzDI53i09Q0gXQFLoLWiIaeUr++
hhElfZRiqQzI+In+Y765tyqVLOxDSckYro5VEeMxUU2M9SDpER2sgYQ9QLJymLeJ
l6/wQ16ydN7UPr8Qm62myBuYfP/TIxj4/7vDQSbMJK253haid6ZM6VvZL54eXzsy
0ZQ5p8gEEyp/taUMHjYQ9gDiKv7C9QEbXCvIHwNrRg0pf5LAyqVMUBOOZ6juhBwc
zpNkHxYPLDyYiFHulFXddjxP/ZjDTIXiraHo3ren5/BJwHupMk1mm2mthTJNqfBN
exeN0z6dT1ktPrEXkL3yfhJNrEOXJChA5jaiW0q6W5NtZqUbu7jz5BUhmIPL3yQ7
45f3LRIc2QXkJXGUYAJQ1vlJX8a6Wq2HfMrD1K60aWi30ngyzreZigpAn0vPGudv
cQu1l5lD6ZCNwaxz8nBsVfVJHNy+xxuODeHk2SU/IZmPzVOlLBopiyVht5URQ3ah
fgOfTiwDBbzjLnxThbwOd0mTlgIFvBANtRU0qg3iGHWyF5K2QlISNeRgzWShcOy4
VawSjGduD3cN8g9u84QM+u+Fay+M3yKKK0gS5c85mYAcMEKPTe/FG1JgLr2sJ82y
emf+ZihG3F+AGu43v4V4P3thHfuJhBEs1eD5Z142+v3amb68phQ0h40JWDdW852V
UtyUiBTC9stM856qUY1tT9vYxJlstgK3UwP4k+/Qjpr7Qa3Q3itdFanAaxTL3BNP
9CFBfLcCoVHfpu4hEMCfo4H+4f5DusqVABxKUC7tCpafXnb7gTVYBxBHxlYbkr5u
a/FRZptTHuJWBXk+wrT+3HoDbU/zUHT2j43f+fYvwfeHp4Szd07nKhamUWWejn+5
kK/ArZPQGejgDzJLoOMlNOcz03Cc+WwFdhIxMKR8CdSF7RJ4qE37vBBiszHZLQ7f
CYMJWYUTWS2rX5p13bnj65mk/mfiaPaa2BlrwXQTcOyHsdrLoduUyM8FEyKgSpHW
9nQvNILZK3lnKknmoPr5DhkFMLNLqW9xlwO/kpMnrko+3IEnWYmavge3PwabBy2G
KCvwqNTyHf0kDTt6U7zKHFZ+sleZoEYsNkmyvV3yoGrHPGS1qfdTeEOhekapN+SI
LFsWrb1huewuSB+vilGYdXaQgksEUQy1vSdBv6+Ho6w9YYGyOqSv9QJ3JdhgdfJH
NpkFWtU4E48LS4LUcBYXHhRlLEvYjXaleGS/OeL/DBD+T0abGgSvqjHIawx9u/kA
kdziDXhP2sXSFUeOFwHh0CZh+ngZajnZgFfTwR1X3ugfHvM9tifc/2kuk+faGrhI
mbslt6pKgNYtJNDrbuY2X/4iNkfmcr02DwJdWQtATAJBBn9hYkH8j9y/CcOorB+L
hthmb+VTzYisZK8EvYE8kUQ5u1H1ILkqrgD/ajF00j6km3iSGQglHObOT9WugogM
4XBF5DlSpKXjuVU+8CTkiaDbx2A/eNdsR8ijf0s1fjVCNrB/TtIgQ7+ltQV6EIM1
xanwg2IYLXVVtL4JyRfupxEHxtyaDRJD8lgT6l8ib0MuYzjkzFS+UNW7vvKG6ZxZ
ORwmjOZ+EYuNIwiWm05dKcYDURJyQe3k+FqG12CUfb1FLnfV4k46oxIao2NsA/Q3
zZzMeo+achjkxhendotrRWVTKmhRD7XojfKV7rviDqFEumVTnx5tu4rkitQnU+F/
4yAA9OwUKOR5KRvwIEYNiPxtquFrHKSij2kAhu39kjtfwx6YZ3DOco0CRTYVVzAO
uaJbFgLe9xIScqNm5peL5BiZNc3RIArJWAtZu8DxhT4nahWLPZltXfcMw6YvR0++
0qHK4nRRjxhEPfqxuXkOgwrjtpstFJSmvdOAku2mAk19kCj40V6osFBFIgwYxSIt
1On2onfDTwkB5XsVrlcM6ykRtmNUFkZWPgFQCwzs4fWGo+swYsYMJhIxcCPhoLbK
2a31CGcFTJYUUjDUF0z/+8Pfg/vXGLLY6T8VdJ/cGipjfrd2scEmczo5gYdKwR5I
VAib+MlcjoQELnlLoJRsyA7qKxXRAtkOcCSG/3wQR40gPUcor45V47LnJ2dVXYIc
y5zn9HdIpWbb1+oShfenRqqtxwcCCgG37yhVn4swamqd7EL8oQhtrZXHkRdI2oq+
lp+lQMqkEQbvkKTLC+pPkpdhaSg6R0TDL2fUjsVYSmANkDzkcIA5o/wd89uBCRP8
0B1gNCm8vreNmzWtUHdeBVp1BqPhzsfoaXDk/KauMLVeu8fxYCGPh+aRtLjov/ls
O8DIkpSPRQeeAT7oJ1yEC3x/1F/7D6in2cWlRMV9zYJA16hp37UR1o0cbsREcbQi
pEnr8+qtjCWVv7EZSwy3JU3CoxTWUpOQuAyh50uIj6TJa5WYkzVEUydpW+KmSmMm
1RwIufoSCitarDf17do75SyIZXpIy6nutz+mjX0kT9CLNmNoDlyzVe0B+hhJ8tZR
UNa5qrak7fpJ2kFkUAjAoIF4G3otb+R7pRBb6FCm6GPUCftCbCNSVdBKVd+2Vy89
UpESATgqwYBBskiBCyGOnSZEJQj7tcisuu6pC6ys1ARTklDWfiUh30PPfrrwx4+M
rvTkBPzsNuvxZEvtKmjL0Q43uxamzhbCpSDb8ta3Secv/IuUln/t2WOCxXU5tFo5
FA9FoCSoFhWWQi/PcTcElz4HPdr+wcgLjBQ1tzAlvLpkSK1bolmi+mM/e3bzoTzY
02yTRorGUM4PjT5zXA08Cyzlj/mYnhaKZ45wKtIA+BBcUZ+lyAUlEFkVGPku1Zji
D7Ys7/ObhB/lKBnGRnnj+AVv1/lf//hkZ2o3azhJrd2STOYHaykfEw237AezN5np
PZETxVGvj5IerElf9nKepJj67aC3ZXVKmjMTEuEcF7y3gBPmrjssC3t6ovINCfM1
ZXrJF4qraYYLWD2Y1QuwRzIfi062IX/K1QEJsuUF3AnKoBVP8kq3htMFI91CK2I5
f566rzRIu+7iNVHolwkgDtU6q1aQpY1DxJS7Iv/dnktBVCzMfLN5fbeytzhMfkcd
oHDKaFIm6o3lMCudu+s14QLuSROGL0TpNwgLFo7d6r+CwNw0iCqCmBfOtsgCwwMf
FlCuIXtAT/WB71HA2BF6xqECU0nH7PQ07rOA3/aSxT6rGz9btJRjX68ujXo0uDFt
z9hiWwnGEIhL/7SsWymzut2EtSYy1Owe1xG0+ntnYGeMcbh2c81cHXqz/Wkcs8Uk
2dQAWHIcejfqwTujAYuEtgDZZvaFm9LWUUhOCCAz8/nlRPfZVZ29ra/BsluILmuS
XwXh+icA1c+QAJiv4W4xc5wrF0cnwKsh1U6ayvyTgSLwOIQrV70odh2ON5hSqjwY
0jKXFK5Rk+zYhUOAVzqaiXkHnpX2beYWTtqGjcGaOcXSObNnzV1ktIQSB5D6UBqW
GsQnuTqZ9fdv6Utbumu8SOjysj3LY9yCk12/ypmpl6KOG9ZyAyFH6K/YjvyT9OS9
Y4veDl9/lvRQSXXZpNARVMIjiuqdtzEAWNNBdDNPMFVY8E086ls+0zuJS2/+/pRn
EcKO9Iodt4/FP5JAB3FQ4csz6ZZ5pFsSwSHELyKlFsIN+u3goQls/J+1gu7wi2+T
HnwmzpeJgklnarK9hoR+ifkQHDyQg/6cFtajvHDFk2R+Pox70OIpXr48u+ihdYSw
`protect END_PROTECTED
