`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aV1YlAd96EpBaFwd7oe/ULO25Fo2slpMeCGG/fkfP+kOVCrVzaCPc7x4osGoA71K
Jm/h5wKRPAFBDZAFVxnQKDoazLazAFqhQLdx6y1cQ0pWRiCvJpN/0qPsSqvy6Jm8
KwVM6e7Ps9aIIkIrAaGUA6fmIDdgJesGDE0UhQPCy5EDjVhQFiYFzBc4al8PGzKN
YnP2GBSKxuaJQJuFpwXkBWLbutY2ygTanD151FHVJu0Qblfy7hK6mwDCR5IeUN9Y
etlCMHMNnWuvyWW4e62S2ddrkfpIZiakTRAiHvSS106TMzh/JM+mxbWEqtUQBrQ2
BdSdThJFsu/UeTq2I9IsXB0srgdcnqFgCinlqevc9sOH6Hk8sS1ZKK3NP86b4gY6
fq4YoYSVq9SSLtRNzHvxV+l4j+OxD154Qe9f+SDPqv0QWu0H/W0z1ZVw0jXGqL+Z
SJErwIXrOD23WkRsmE8ub/XCiBOD5Un13W2gDeYI2SiT3deUAoZ9/vShb1zSdRxb
xG/jA8zWqH4cgKyfZ9HrQTGAMO9S4NlVyHYPIfSBt1DAnWLvZE6EUpJ/4IEYnhYk
TquRlmPQDNug7qokpa7FZMuLT2NzoF6xo2gvWJTGeLE6AdZQ4w5tb46LQnaFIRio
YCZRG/7mQ4OTq2JAjCyY4w==
`protect END_PROTECTED
