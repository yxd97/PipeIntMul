`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ssVdtT+LUgZgDTyP6IZWkFHUj/OZWHJPz7sb8mDR+HWCgrVQbnWiPgygoqmhVKYo
66vqX5mfdMlWAPC2oIvboXF+yZyPJ3yQjBftcogPoDvveDth0U1toy87xcmMdI8p
wi/hz+Pe5GbnBiXoOwO3a+LdKyJCNG9EW9IySmERJ0EfIKPElaO/pHX3bgyg3pUK
MM3rk/xEG51LL6dTm3Q73/mGdMbI9OmcdmhaxY319esnYae1LFH5iO4vxng0wRBT
Xj6x6Bgl5+Kfi3vzbosoimzuRF0isrPFc+A5GVT01tngIgBsbzBfPGKKMOuqNyVJ
G+LCzeiLHJkSkVWUqUEQIoM8NR6a9zRGeQ+Z7mN6PC6TP4hBC1rSWd/tZvfIYnaB
cNfyLEh2UZ/B8TsOXLpWbrkY2HR5aS2aJAlsO+Cb6eM+auVl0FPxftzzwtlHfJ0a
yqKTCmaNU0pi8aIVBUEA76BW2X3CKVK7Bj4tASzk62F/mAur2xD57jIMdiiNnnQf
BA8FPmFIJ2KnyLIaW3FTiOa05XZ1KxxiEWhiVyabBBqIgWZbz2VFlG56v8zAaCnX
ccPUGq6E3kDYWQY3yhxammynmfMb7t0SXjAsbE5myf7CyEUqdoXYgj78uaK7o5+r
asy8SYZU3N9FRe3fQ/GY6xnefSllk3j7Z6S3MPxnSKVZbUu1ocgVS9DK7Mw/qvb5
CMQ1gxUySi56UaCC+wnDoJ4UN21mHvla+eMFpKOzDydknPlHLYil9W/xUeQ4zs5U
yzheOq0EYv4FtowJ+9hmjOtCFEAP1BSbPZgk/wpn6BF7oxw5hpQr1ZkG6ElqCngg
+bFM42A2bouK93c3ISyadg8R+8DcW71zBYsY25eO3l1rdzq+MzS5aVK4FsyHp6qH
K+dWrlSQCkxhdmJgvUa6NMTICWFqxtagWOWu6QWit/3OUPG42eFnHsnuve5u/4vZ
OU1QGUtVeNDlSZ/PYTvsRvjJa7IdlkeYwJmp9IYo/xRuDnPg0lEjp04rpZc1s+Be
nvPrW2lkIujPBq45ejYATJFPPSbfhAZmE8lsXXYjXMBWWOesqsvftu7bgBj0a0Gi
UyvJX3GLE5k2uZs2pK/7HkSSff4GpLoPjH2feHwTGNa9z34xcmWvnXeyrxLpSRaQ
iBpeP8+QGlcR3nI19r8XKP8F484NGMtiDC1AeHtVblwk8MEiGvpWyQSAL2v1LO1M
ZHpvVjRjnNaqSQ38usUuqYb5Uu9CeAQj2GpG+uFUBNz3eH6xnS3u4ooeaTp8Hg8l
QzyD6EgZcJZAmlp4pK6HrCcvyo5KGK6/TyOMFEI29bg4Fg9iUy1kVpMxBVGFjgm/
R3KNRcHMp6F6qtPFU1Uv7ok6Rf5rk3u8nbPXWS2kHBMrt1pYn83XPQqOJgNHmxx4
oI40bHLdOvqN3moYTK9MG+ERqiN4SSFR7N4l20fybeiBt+2sSZkK258tYbE+rk91
o4CBM7DCC5pbMX5aXdXdWN+phiwTfx98DN0X0clgtBOcZ0TFHzEj0BsKfxGbw33t
qHzIh6hc+DD7mvDXXaAhSf9DkqY6dBqXkmaN7r0NEF0JnisxSI2xJ628gWdVpp0v
FS0lolUeSwu5BxD6hsHbwBC2erS3U+b0qsCsBbfzWQMP8f7mmPdb984ALVsIX//s
BIN+ZhPm7f2Ryc3QSz+juND6anFfWzAZ6nlLdvJg0NwPwtYBi4XX9fB7Y/A+MuaD
AivkJGetfQE5JkVWppIYhKXchw40ssx2RJnEPOvxFkbAaGc9WtRwqh1dn2xA6j1n
IYq80C0rY8TIspZGwpWjBta1OY4a+sfM/S1EEwk7NzeVgAwywsvHSYm/EL4abs8a
4u8Gwr8wopGmifLkHrm0cI3WFa4KnqbFZNrQ37GnBlBUl2rtFCkKPLH+5bT1LPcg
cAEEwxnVWnpVjzWiBm5y56eMJq4DJ160hpFhaDR9E3STQmWeo23O0Woqti9THbux
/okRTCmFy86S7/KBZkrnghv7jQIgrMuYK3+GvBQrG7UX3LX0aLJTeNKjG5yw9nGe
qbq4CxW8DtpQ50DgC/a3JYjSXBuk9K6s0wY9NeBpPVGrxXJUFyXTra4JN/vLaOtT
/tcfZEX3KepTWtAB94yABPnI7jSVROsahna7xNMBw+wSxthzYET82s6cN7HFl5ZG
fkpYIFzpYyZSA0Mf/NqcAuZpbBA8/4lNJ0lP8mNkCRmtBzwX7veqe0bpFQqgEGto
OGWVLlw7uR9NQIl0obtTIudVvEtt1CoFLCiEzXG/aOzWrV6VC0vYbyaGx0E0UVUL
6Zu7NlJKycfYEzpi/gT2ccFwPQMYv2neA6j9Cv0hd4gEZJEiE+oPIcF1OPLcSjs2
tPHJIpLGvEioPkAt+SwwH2nxn28YbufeMCGvkrPjf2ckyGGu6A8XuMJhGwDZp5VV
bNQ+kBGIwgZYR8cn4sNDYnfQzugyVJoESW2xb5/JFuvKUvVY/joqJru0CaZjwrQX
r8KChEv4YXJr2Ppqp9WMlgAD+wkFarHqTUD5WoihWUn4sYBHrTlP4BTERGC54/oM
rv6ExFKqHABDfLvAqRW5A1wHZtDcF3g8P32Dj6vwM8CZ/OX1ue053YXwqF2VW5+B
bXKUB3X9FlBSw+ijUvEaTQVUW+8D2c2IJmdXPE2brtpraHYBgfV77G/OyZZPaj0t
AYYksw2rm0gyDgNxQxejtI5JwHnbpeO/mgBRR+/2ChvKfgrsukqnpQUFASUgEFYl
f4/L7bf3bbGvmV/WBMMbEYfxHoYVlR9R9gAdaX3bs004oE33Ew+nQF4GnMQBVFAL
Ycf/3SE2V9i4xVIMJjfQFjoWdqtEQxll83Yr1y9P9zjTrrNG8yWBnbHY+7BRcg4q
Ya3th+VADHm27CeyVCXXeidIYwJOPatWWy0deNkBfl5NGUwUYfLY0Azs07e9gamW
hJY7XrvwpOsjEETPuq/ee98oNhMRaCxoGAB3U72wZ8WCq3OBSwYE8pWnwbuzflfd
/7jJMasxaauclMmEVgvCRNv87St0WgyWqYpTFyvtXf0aJS66UhByqdjzr1f+yLCt
66taR/p2j8614v6XUxTVcW6f5VABXWc8/7qP3hjT6N8LNgEu9kkTswKxcRZKdpPi
CshGKvfSjbnYy+dZl+FNkI7LiLcqmjrMuKKzMlpnX827qpRIP3rUFYk2GjJhu0ol
K447pCgKqT394dPEn8GprXI4LL3NyOe9F4a7Fag2KxlmkTHeOo8EmhRjuyzVlIoz
avmmFzZS3/1TokZSg2WpMdi9QLcMCVfPO4kae0oA8QkC0q+zCQw/GU3q9FS01suL
U/44xBMglP1dpC3bGfpn5DHUws/SbqZDaGE9qBzV9M524weWmaUMMfVXLOi/+aZV
tasGII81C2LyJ3cS7007k5oo+7LDXCsr4fxzspbmOxnM2GPq4fpLuQw+Kw3RsOvz
SRMCIHXFlSyqryeEvVijfIZXZAzXmZcN+enDEUy1d/O8yAiVS7o2XWYdhBGYYfL0
oMUmYgHgSRuuQZg+GooQK1FQau5iFYkTS3J67ru55FD46nwVFkh0davTV/JIsZnF
o9NwUzky/A/USVYSSmQvoCC04JC5vISAsq5/spfu3Yh8WafXnS7Ka2f/IUuavrHi
bh8scu+1Xe2tO2hys0wgjUY4yHZROp7BNoa8foanmGg9DfkxX3bRY8+qviJSMQZa
D2mQ45sz8yz4I4vGu+9QDZ4f3AvK6/C32q8F+mDUUhZD279nMUrm8zcNYXqwDFnL
1ESrsAliWeBqaMx+kTrLoeG4W/RTElROdgwsS7fE1UwT3Px5wridkUll0fJiD45V
reUdeMwoyJpRxqQIDDGPlOFBmkvYa8M0ryLr2IUOL1oJIoKR66R9fbhVpq0ivIDl
UjJ7fMkjm1BvhoVxOEVIi87EeqIXkx8YwW56/Dfbzh/FA0k1gsvl4tU0JsEKRoVh
Oz75hL7bKplQIOFY5lOep2XBZBB8BtiYv9Bq7yaGqcucUYDmDNH4qlx6WCZ0UHj1
H4bDuG0aFmCBeYsi0EyfU82RUu5yPzNaR6itNvEBaVFswPmPhH8KdfyosqNLAac/
xeJkNTF5ZNmiOyCI0m5u+JxdC7oawMmZ3CuCCIHC4hZMrTkYBBECvU/tmB8JDaV0
JwQCH5PFNh1lk1dLqmzMVgEsZ0+2PiTsn5iyax7SRaxjrAIF7fNFrb2uPBCZ0dzN
c5a5d5q9hzP5FnCzkmiigOjbHZkp0D318+bWrUXrUSf3EIjsgs169X4vRTAtJvSV
7FnN7wm4fxzGQfTf7FdZh4RtyUXIzQaZJtFgcHGLkDf/C7fJhx+vtXl3F+rTP6ZH
E6RR2wBOrGnU6Zb92UBJhjuXLLaMfb6N6XrLR9zKBVn3Wx1MXQB5gW3GqPcLlMYO
0k9xvr9NhIMjS5TWANaBScc+oweHBrkw/uGAK+J+9GnWeT2NXl2sP+LuQhiS3Svr
YP7tDTh0f05EPYV2KSm7aNJy4ZjCNM1wzqFxxrXsQbfI8YP5CJXiGWKGuaMjIKiK
Hj29O98quzAn4QQ8BafVd56fG1uiRWFSMKOqobslIzz1236naZnaatwzkkwSh5KR
LgTk72LPl/M29NEwTZNxCo722cMq/y/opAVwZs9ehuE30LIesiYXCyWQDiY7hs0L
issvRFTdpVyU91kPVseH/lasQ+TIOjZL4b6wtmzXUoph7TI9KATdj3ppcp2XecW9
MxEGKFUiWbZS4cDpjXHOafJujK87UDYP1MIMkOFf3zQvLkx50N3/Ev1A/N5wiAC4
BtqwUGlQ7dxKidz85XzXTNnG9ytNwOuwQXb6mLBrafDjvHil0QNd6y1PVi7InuTk
j+AmfblAuocdPg+d4/xFbbXG++34kDK55CSRoIXhz7oQhkcJXXTEf3v3XpGjGpso
a9ZRVJbblAnkMpktODBO3qDiDirhqS6tqOrm0NNqNa7wafvLhNx7ycX9M6phULLe
7t6uttkPlUawCErJWrYLqBNLeuJbCUM9CDvA/ERDcsZW/+1pWj0c40gvSH5/RVQ6
IVukRDOuXw5WevpZXaTvf4OypCrl/ss3ShU9amVCtX/8aFMD98SL477ydFOmnL8v
4M1Fj5wUDWqbqeKYNamxVIRRNdTpm8u8ROzg9TpAmN1FZuR37ehesJV7cgfKqGEi
rH27su2e9k05dU1/FYP3ktqBSqX/OAj2plr048CqGTmSvpNX7ur+exHIfPsldord
+tlgECpUVHfBTBhUEng4SBZkAnKN1JlZvWTNq/dmsFOcMpAHTYMfUnjXbL1fqlQU
8LEZXRCJgnkyX529wyx/O/u0BBwIgArC+GGPWi75T+F6Q5R0VMpV6Sa96xCV+I4L
y0h4pHdE+VlTktiYepEE1oQMFsEIWW8VZP1LX6cGysrBIZ4rTNSoic+xc2Deoklv
ILJ4irLXV54O+fgRix7XQAnssjSGAvHK7bVRc8OCkgeh1gUxyfQ03i8cKVSPtf9y
mKyDdm8vJz4c3FuGg7qVR1ImrJ+iQ/Ubyeqe6oIzGa5f0oL7ghZmASetIOT8p5tl
9tlQF2pusg4x6AW3uokV85S9+D9T7padfEeeagajxF5mYoC718ywhFq4X2s2Z2PK
/iPwR14mMkzo+TcWXE/uJ4PmI6lt192eg4xIijhdPZWGUqAVZQfjT3vx/RNaMlaH
P6VfhYlJaCiIDUDJiJmA7mkIn+vDOwcRGLRQsDUht3mj1/5fUg9inqQRwv3KePeB
KVKCJhQOr7lATkqJKm8UCcCH0c8Oz/c2pQEwigIxfTLEqm9aIxoV0G4dLo9aU3EZ
EhXuP2MA0Hs9bDH7fxZlB9upGuQlacconvifjWA9TYS/oXRQ/9P3UwZy4aawqhn8
D729t+GJ1Zmr0p5TOndLd1xYSabli44e9yu7FZiOeqK9AZxGYN6MUBRsz0B/sIdZ
o+Cv5WTCHgkmXmvTtRfSRvCMs0aRLC2E9+OflBWFefzXbg3BKwUkEw3Jo13JlV0W
X7PeJWzR0KlxaNHIP5JWSrlLcVktb38NhAFcW7k1Kmm07wDkLfWSOfKiYhNzD1PU
CKvL1dlfSaCwyU+KPxhqyHoRiUUaIunDI4BhUG97x5Ues++Q5aPldFwNcy67exnx
5p+FYMPwdh3nq5At/TAHzjIt2kKPdmNQ0j2BujN9lzCBbi8vLNMMRh7YOtTCHHQp
+RY7L1rFYHSkJ1BB3I166novkIQArFWZsFRICMm6/jhoGUNTI+dBUkN5bEscR4QV
FDlPhamXdRufHOybaSJeRS9C8GnmnuR+aQ2U30xzO03Fzc2qRLL3rZFGOYmUwf6S
X/2OUHqSOXiv2rDbHNNu78+g9IeK6xfEHg2leEZgs1BAxyw+hAi8QdPOdGwQCGRQ
Cd6gGrA3r9vNDRUZLaYypGqkphse59i+9WAuyU5yT6Wy8UI/IXKm/vHqgGZqDBif
PTBD2rf+QuPhfZC+b9vhY05S6aqjoW1E1SXJDK4wgqoK/UpA46mSKYgz50vUPacz
Y4RxK565ucKDz1p3xO1xZPGHEr870I666/VgggCBZPpiF7XZiR3SzFPTa0R2rGyD
Dq5ZL+ss6alOi2eGcb14ZrS68ugvIwCAO7Ndm3C06i/lU+h0zLhjI8IuqQTLY4jw
Mg7O8c459fGOYBbReHyNWnnZbv3yWlk7FjmQ1nDS76kPhGkYR0JFmOnYCwcQOcg0
JlrAmXoQmfCvj2IhDYaayWkVtaPGHO3CgA694ksDutyCvphYz5S5A2ZCezBw9WBT
g9WKI99OI5Qtos8Vmf7VCXhGokSI7VY183s84xyrpP+ewhL7gOk/LakIPV77tGMO
cVxz+5HTLkx1y+7qp26U8NITwVoz37/sTIWxjfhUxPl71e0NJEmUmTkjpWeaAUWy
+FOwsXq/LOOtYlJCcZt6nrwIFaL+MANChWg2kNKnkeR9JFL6drw78NmsRolMIiDS
KqiFcU4LGIal5p62Cdd+QnngD6rpX7q/O2S8hgrtBmg6qGRdK7i7haVMJwTfaTbG
wWd4fqKih9YU94Ybh3aWiexL2NhxgXiROVBJ9x5nvO8LY3DXCltPC8M2h4IEIrCU
CUUjBoSTlDOd9UXJzci4jS7cXZzyL+WCb3Uc4cESpyvRIWgVbowhywItZES4p/3s
IwlhUG9QGoMyWZov4PtdrC1U4w++HwAGFCcYziGNbNu576iB/xOfYlKwZ2ixxn67
IR8LK9oOy9eqNFItgYKbWLRyMx6U6flMRxECkGbk37hBl0K6zgEfH3x5qKgvdc8z
DBn/Uk0ZOyy7W6vro7c65fQyRH5DNgD5+X0G8L54cPZ+tjnmunM+igOFej4XWYOw
+Ec4p+r7HsIu6tpfDXtiXFzOzw3gCrjabeMIuO31ScTida9MkCoJycuITVqvGwhb
Qr2akSkE+4tzw+OFx08RpQPY5iUzyS8AOtL6eOXPZXbJgB0OtUbbmShDZntIz5wT
USqS+N9xNoB2Hp/8T2omtep14dhQe8oonJMhl62+FPkADkroeGbE3HIznaQk5tpI
j6aaUwCLzsIncG+0I0kBuOFkZ0884sfknAcw7drTwxDkOvQL86T7GDz4upJ/3ldS
9PpgVPh4Y9xfwd5g7r6EPbOuKZZ6SY0P6NkRDFsbcZtHXcThlTBK/rlGFv6+MLAF
4YToJbDzOYUEU0c02YMHZoZZ8XpScMY1QXpJp0J2yJKldhvRy8Ngag73PBmYP/hk
kdVWQ/rQ+WneSiEioux6us5AUjRvo2Zy4gifAnh6SXrVYPO1LDkwNrA6LsYBZ9ni
cCEa+9pbbsTJw2lpTUGvGozNMyX6kjSyz5sglDr8dia0moEJ14yZ54OqW2I255L9
Gxeo7IMzTL7Iv8V7mfQE351maR/vhm+5/M9PrSRqFxCrkGVe0wMO/ydDAhC/ULeI
vxtN+l3uY2IXsE0o4F8TqnTK0yObl6H1zNlK+gm4Acbccd381MLhOLFqYP3IWk2N
gs363ZUcj23w1/PlQ4djEo093wwNzbR4kX/UQzvzQU1Ontoin1Nm3S+QfGD2O/Wk
8zOvPlO1sa/rMTTbsFHFlQYpjqZMyBylSaip6sVuJAFl4N4fgTG1Nk/d30EkV6/r
DwxKse5eRsPYwEYeXc+0DFVcHRGQIDVAM1c5XLPPfY6WZa7ldnJaZjaqSbpHrllv
9AFGerpNzRr04rBTrIb7oOUnyeQXcMUhiuk31DyeAV7HlDYG7Qkf8RVPeqlQc7da
TdRmRuxhOiqPEiUQ0D0gIy1yI8hI+BtdGAi89Z0fXOiWzSm7bMh9rf4bOj14A8W/
PWzXwHPBmu8XG/gko7QDCC+ifXPspC2nN+3QEGIqz9M0yY9jLZ9lcL/TjNa7Dvnd
6thaf3+6Qe+RLASIQGyqwMwLfOv4pOkJmXLCFT5LAnciwlKl/XdEh14Gcm0X/qQ4
6Zp9qPmRfSa+7nNdkf9lbVBpFeqNvb6N5Ijv/UPsFbYqbDGsbRa+3VzU24vXFhuv
w7xy3koOon7QT4S9ihBGjzFfv0sMpprtwsTgCrp53Ronohyy7IN0fBFe+HgSvUeL
zdglU9FAXyi/ul+kIkHaGeZDvB+U/aBrif5BALLXv7DOSeRSGTxcswa6DcBryC10
BbiImyFMqtuj/Aehx0ia5BwkGDKgvjb/p93LA6wfbdIFSYb4cWmnc7arUygCm/st
CR1zySB3ieU6cfZrZcBIcOzYB2kAufJwsuFbqvh+l0jmG+IpSnTMHLfqEVOUFsHl
Ned+KYFo5FqGc+LDB4Bb9jNH7uZHYrZ63P/AIHbrUcjA8R+IZ32CsxxEQsrX6LA1
LX/EAppTJcS03AlVv3cMMTiTXujGr+R0AHGRvkZhqBQQrhd+F//+bHmzS+U3Tw7C
F+eF6dBItyxDzz5aeNgSLbDFNQ84uxrFZsVc0w/lVoQwboHmyOuM0YAAKGTDNB3a
JJRSa0fc0D7GoYRxjlkKX2++HMuUCCccltzmsJ1wyHyECPqIhrFhuIg4Nm3o8FSL
JG16RdAXZZbCWKvh/tS9RJAi24mlFTtY8QucCuU+TaJTuMtvsl42xM7bZ4S+W8lm
69EULyNphmIog/VFvhUA2B9IJPzsdgLKpEvv9WgUa5UiEA5jP6kpMGRteQMg3+h0
LzUc0OoaTKnKvHDvLo4xJm7N3B++Hkxa3+Gf/AJbis+HIHr9JymrGX9cOBaUbJ8b
+8TnWaEgigXn7lExOpc2z4ZLF/lPej/+ptLcYZGshgecYMT5/MF7qfhO3fLheBoe
OgwRE0qYDVTKNIFJEWCAiU7bdcvLLVoSpg7234MfT6ZUe9VH1oEbia5Ij4thz6us
Luhxww8mdSX1xVITqnZ/MUabGeOT9eI10Ickz7gzcXqd0PE1r1bQhygFN/qCSB5E
8BvG2j+8zQGXsJHU4X9UpWU0EGks/KNKHqa+AdEdisge1dGTjJbkDOwvqs+BgIbX
LBgMBwyxfSOb8wDsX51UhHTm/vvy/rsBCGYdg5mOXKlF9lHYI15MQh4kl0WM75LH
8QB5cQu9scnS90qctEH79kxORAKR267+4io1kqxsjJEsTWuzJBhaQLiTXYwgrxbv
fpwAuZ3uMXu6szFtPdQ3WkfoG4NsxQPGMWD2V1V61YRzYTmVm1y37MsfyAjabur/
D0Hg4NuhP53PkBSZPqmNUPPk1b+VJdvZ1r5AzbCC3FV2AL1LF5XIf900cXb8KKgf
WVQgL8WYtpNUBrgTtSHHIYrnq5p3Q2CHmmQCmN/lIgo+NyeAfGjyQLiBm8DUQnod
otwE/MCw7E87d+U4ozQdCgv/DTRNDsO1ySF1302ijK4nBceitS+Y7lPI+juIPT6X
rPKjffYIZDhnfSpuGoFndhPeIli96bkhCWtQdig5tRSnK0pT7Yyd4I+W0j7NaDJL
M6ekQt/eBoXL9d5bUfpqLFuzhRy0EiFHNZF//cufcWh7XpiNptzuqOopXjxlcbmg
lsxnRWZAKBzvSWk81rU1FpAMoqJPnawZ+QCV5Ll3IbcurQKTLiQ3bIZm1FYo92Ad
XZjcTRXFuZRjXbLKQdnya8vIDYYF6qjTWQXr2LwYSdRaXHtNNEzz8Nke4989k+t+
A6Vi4A5AkILLoSIkC94PV51FXn46fehK/PlgGBkJ1pb1hiE7c8T+ESQCat6PLJyE
yYmIaH7Ai/27BTaBNjdVYlZ7ggBFNEKWrXBq5vuBibEgXEr+QPrdxi9RP2Hbj6i/
NfMVkTM/lP7T9ek/q5Kr3XYVuCBeX5WvoyO26xFYUyk2innFebA+Dd+S+3mWnHE3
85LhRtf8W/Gc7o08aYDKaZRL+yTsbn8DQFpgiFhAe2xh8cWVcQDy3MBiwo0LyCbP
BSR13eV39BGZjQmxoLCALNokcO87o9iUJ9nDONg7bcRWGaU6mWt3u1VO3+tMu5t4
TIj/zxitpKJnnkgPeNQi+pKqTXb+t+xxgNEILsAXb4L891UEZ2T/U8mX5IUziK2f
Z1Ej12/wjcRiSUJgW91eVzUH2AKvuby96ci/DHdWmc+zaNEY//oh4m/TbRLb7mPH
uRLXepF8YZpHF8sS6YVdcF46QriDsJ/NakVaZLlN0Gy0/Nf7ED7pLDZyK/MlcWwW
n7x6COwFjV9jTWGjestYUVZQTKSB1SLtCZRziUck3LxnBVqXmkT8k378KWZkf6ZA
7hjL4P8YFkoZPy+zMZ/W6tqLYzalMUvuyV2FTvyEtJMsiyU+fD/B/UjOR6QYCqS3
O6hyroz7hBRx+ZxJiiVp0MHW0PsLXDBWCgmPmw0kUDfB5APjw2KwD2B7joR2mi86
PTigNE25Bw4b/smG3Q8JL2W5F32IOuggpzuSjRZUcsY26pmby0APxdO35zSHMU9A
l0MiFC0RXoj3WMTiiag5Yj3eGGl0i9p1bo7aPlnTp2rYBJdP964w1h9SRlHMFRn6
0swDHzCrM2W/VUQiT7I2FDCHJ+0VvgrRLZC9KFyJcxgbwQ4xo9YylDI+9HDEkOH/
mEFmXP3G5rrbxQ2TcoEemgqU+cWB7mY9tfdshXwe+ku6Jxdk+RBZPeqWdGq9xYz1
icXhdKv62jfPS7nBapnk0lg4Zcibuwy37jQwDMb5H4wyJBPctHx+LYEHKt9L6fGN
E3QYMwDscGT5nG5pP9/5ZJJWR9LDfCip4my+Cg2f5fHw/9uez1MARo0hs8yx93wV
zR/HmLhUg8qW9KxPl9QAsd+EJRCmBd+SMw/wYdNhadSk45oX+mDCLfXtz+/dhq4H
2wSpg5AvJvJNIN+Zqb46VXlF5vcokImJGjrTW6mauNOBKkihdYjwCFWOLoLO89f1
D97dj0OPocvzyeuASTokmReE3TW0zSwi6ur6VdIkRlS1KES8A5JlaFAr1LXrBLLZ
wtoU7zY2GCNHGR/l6WVOHVZdrUpNA4GTKraM3u4AX3ko0DUleGLlCoUuHktpXqMA
HYQUUWjhB3X25zFkPubpwJjrIUB/nVsR1mPqaS2EnYJGQlV8LqHRI033IA/J1LaX
tyzNSKM1Z27H/OndMFr2Pvv2pug6wGcbXWBkd6DVsoHspg6wjB1eelTmJp08RiDr
F3A9mDaiQMr1T/g49BJNo7haRzb6eODUemZ/RFQtoW1G/AmGsmqQh7Bl18gfcld2
cYw3HfewdLZqIvq+T7WFmkZJ8Gl5vNmfoTcExixw9U+MbQ/rPwjTPu22QoyyE9AJ
AnRMWFFIcNlQUTIwFGtqtvu0wvzaVMyzX7KsUMdvkPfAqYvaxkJ8kJfWbF+h3x3C
feCjqQcrfHvVsLPXbS6tp6GPrDb5tfrmgmqNxaRS3yBgvQ/xiqTlTAKYhgUV0lGW
E9ZXE0IEHJI7G0w7SCrLwRJ68oD+LtOSrpy+JLnuVt1qBu+S1u1RWpWHGF/xT/FQ
BeyT5tXo4sOxv7acUVGV2K+NJAgOwnMMAy6/CoR2WrTgroy0Tzr5EXCovZtb8al7
fElO1Y1dxZ+IkOXIylG4a5vchNqgrkReA7Vd8kdsgJC/Ifc7kLJ1n3BTwJB9lWYH
Hi3OM8R9EZskU1BFGVGElgJWE8BrHw9wr7cbTKRsruX01oGPEwzVgph/A8yZyIIg
Q4F88Qwl9RjhlQCvh4rWcLaKiGjJYpzsi/E9ieDPpYHAyJU+oAFln9z3BhpQH07h
r54zegAglhP+o0i6pXcVzSMsWzD0C5xMIF7A/xlt7V0iqRm2+amv9WUjW66qYVM9
2czydC1M3/vfGQydsUFKW9/vT/U4wXjs+qSGqtwwnU71+INRjTLlCrLUqsriUMR5
HDt62tT0iw/bzPV7mgNcvC3jty9BxX8HaDOUsVow/caGImsuzTAuC4hj4u0dQ6d7
8E1UBph1FUnF9c6P/sSFgcGjnFz3YIB3KZyrWKC446KbcWJvZ6277yRmkKCMTPE3
J2wLnilabvhUP9gl5A5HmVAj3WOHhFc46xP4myje9fC/SOqjafkgb8frD26nfWGX
Q3YoLZTVNx6fAi3BaQPCZGc8ucgBqfGbxDWokZoOKjy6YddeMYVRFkREvAQKIFeX
uGZZ1GeZPAZ4qLx+qBlQbYn1INw8T4t+PgNYS7gB63YfPJxcBC/DiWgCYqB08szL
H/llBASH9t1SO6lCDVl+PAIE0wuthFlKrk6kIfbhKk0N9izXeI4SrdbqMbNjKCMs
/wUKz6iCKmCSUfHj3zwtco1ux/nqkMZulMtXVBYaccPrZ836GV7FZ8yRkoo0lEdf
gF0+q5oIR1tGGiN5BBBRA3kdMRz4RcVPpN7r9NfVCy5NEzjNA05UKZN1ss/IuLrZ
Ewpo/h9CUD9zkYiw8lVIlRrmCA2DWqzPUZgEB+bvwTOfrjfMNfOkgXRRCNeK+rBQ
hMlA6nUyNFiJSVC8oHv9n70e9jeF1h3f/PHFWJwRSrPgxKg/dr9wGDzoQG88smIw
irHyNXkkl0sKUUnUMPsUtTKjWBnsH+2I0rRNPOzXRsE/MosiCl1GiiqSkJk6sfTI
/qN0Pz5Vog5ftnIfBlxl2nAXX2i/dCgDwkwuRRO4/7b3QUJCRT3sEFs5qei3zX+Q
QmHbDsg9HCm5RUeVGJY+vjdkKXAu3tYaE5cBBvAN40jxV4j3ru5aCHNz/v1rtlXM
XKG0m9ewIQZDdCW0zftrlILg+xE8trBaeth0eiEEsoW7IPFnGnG2ylMeTRL4rAFC
aBFzC48o9QzpTMXs3txotbdt5jO6C5UYaet0aryqA1PMiQ+qxYkeRFvrQ/jrdWyl
vr+BEwKbgQxNG7UQHWf0oABHBqzqWGQXpXVAyQjjWzUy4r/0/j3CSzhfNgdSm1rH
rhCl1Nwl5AAIXjRrw4QBnoBZql1PR1eHweUTwhx93Otox637sK45j5gRTndiLKk6
5iDP/k67BZd3eq9eT7v6LGbSYcDZTS92Lis8RgoX/W8tpDQKqRTRxf2sK41iDc9N
OPkc+Xa6oF9XqgFaevq3Fbd3GNzCIAG8TgPPxenMTuNJIij9V9SFKviGBszr4XjY
eulAGou0rx2becvMSldRGTcyhwaKlA9Ni2WUb9ac0aj1vg9r4IKwXT4kQhJsen7i
ybceCX+zCju9bJvTWD9yFUlGm6tI63Wx0WyrrSGC9Q/LMY0apdh2nPyvG+vJSHYo
bvDYsZFiNZSjd7ABmN0PTROnQuZeNC1OJwyeSogL8El/vWIzpvgVD6HJVw8GHD+H
T9ZF85ipXrXotzKjHKT6Z3Q/10PhFDcdtTGS6TvtTfp6aWj8fyb9AvvlKE6y6v5x
87FPwFug0MvSI7vHrErLfNhDf6S39U/X1+q/2IWNdHlB5BmhI0jIEhBPYMXngXf+
JX2/ghlrFqZOoNtNwO0x7zybPoBjpJ80+JAnsTywklaVpqUZUQmoa69W5yIksbCY
ksv730dJoapOBqe+OQZtT9x+NmirC4hnSuwJ/2TzsnDZLTTh5/uYU4YnJglxH4ip
aKnPR49PBO8K3PAFGCa8xfmanolr3aKXGFmvMIR3asmshx8fP2kzmv3aNNr+NpMf
HKFgsA87Ri20mIYJ9pXti2cgHqJaQrZ3dT+u8sd8yDOF5ZUiV+J24cNFpFf8Z1Bh
m//fDseF3J508xEC9FuntY1H5nh08k7n//UCBXuz0e1n5MhwnI7gJrJqg34/lc2F
0cfyfMY3PtdPrybqAipFkFm7kgVSGuVX4tGQheo2VQC0Bc/eH28n5J2UiZg/o8r2
ZcYP9zdXBB1wQyIm6LAyyRY4U32INp0Bi+n3D37Ftqys7KtV7Hm0zXGRSkKYzirm
O6w1cA1e53jFiPUVLiXlLlbLRBF2FN310sF+Ofkz+EW/V/itJ5zucMoObBXDg3OY
G8w3XMRr+z1uBxzIH5i51tIpHjZXSxSsYdNM4fxDOj9ZRjNFtcttjV3PwxRyA/Qe
dOR9UudUB6ifOZHwGy8uOU85xzcOH53V7tIDPXU1ET9lgYwJ0y1cWY7vKRJ8a2Nm
DYuqMZsZ5/II+VgvzAuRAW0swXx5wH9EGLajALRQav/97Soho6gnwcKwgVbM25cT
IJwTvFdcLX2ccigaQKRx/d1HUBV5aHvFyLORO0kCmFFk6cZiA3MQhWAA8l04g5R6
dOBdwWRHcJ85JSPXm+TqhxxD4d27JkviQZiZijxny9u1drv0PWUTWNfd5JHNIgT2
QwpVyYnY35gWCTTpqIPD/rBgJVrY5H7PEOxv2l2C4VOwBRvBYMsrfWPmd614RVex
I3U2zrdQhNT4tXT/2ifZXsardwSrfH1Q0mHrFnkwUj9ku2mxo/JdQ2H+Ivo0nqEz
vEcVyNhB1CuCQeiYQLLtu7cSxhvaKNbzxEpNPHp0skynhCJIR4YFeGg0EJBvCxrz
V7wRp+eSsUXIbpUN7UFeM0HMWfvdDrn1qGJuI7BNDRhhaBEC7yyQU17Kskm1hyVV
PByA9YRjErjpiLyaceBZZWsgNdJmP+yYVIKod5VQ6eetQgcqFE2tU8SNpkongnsq
RSKVEpU442Uxs67VTZGRGVm5fxOMK/AaW0WANyKLeHBQF9h62hSYdoIEy7SOzvjS
4Kw14P12YEc1ifctbHJaQlMRnHmc1xjHbwW9VqbfkwgyXz/LHiZHJMsZ2+CQ75vO
FxN50PYGLf03t0Pk38S+Ps6XcMa29jLl0KN4j8sUB2wL9PCo+71cdyKm27A24QZW
R4BlvGKMMUJ9OxsDrQS9mYjLJhG24IhK/oC4mzjzlxnpMQIskrM44gWynaaLUnX8
qB7ZXsQNBLK1RUDeLOzRmXx0E2+S6oePgQPuA3jdgq9/c9TIy1TMm68BaBP7x+yq
qBrMkXLHEtmD73EfR5UfW68denoih6N/zgJE4CemthVcZHgCnMjSYyW8YYW39BWG
01pZj7HILcSCwTNbX/WFPa4IEj4ig5sX+W/3xXBhGp0cNowEiDxBlseghkj7XnPV
jDzto/i04t+ojRmx4Q0SClNBZTkvxRvuGS8zD+ZSVNaL4JJQYESlnB//XUhX8F5S
4Dheltj7y1I4sbzwHxjVGW2Fy9rBlpxR4pGm8UYgYMDHR3oAMILEyH+B3BAVS6G1
lXfdq44RL3wYLxlFadpyc6HGX1m8K6jA/R8D948nPtOp+pOj6tkubutl+Qyibd4R
4z2xVIv/IhF4a5FXlTYDAbuVCTFR1EP0Mq0L1sIJNxD2ASpnt0qFvArLxWwo+J5S
T9Ni/HGtBRGeYpxGuqkqOgR7lVAjQoChAGG8EQPrwlenEzzJdSruZr0mVxCvL9+H
Cbv/cZaFpkRtVdUWpxib8wK6QZuDsm5me4Hd0QJmSFl9BvuF+YZ1s4qrb17qFoo/
A9a7aFejVkY4cyWgukWmVvns0UH88VnMhnAQeqUsuOqnN2rJUAAcRmA9K1FJ2uCa
kRhgODwjlLy275POn5F5njYs7kOhH38l8dmB1N1kkesiW4qYEj7vSZanaj1HVmJ3
+et2HaFZ618f4esJAAwlEQW7E+AqBffTXUDTdpDIdAeL5yJLScwSZfgBvrqchj5W
jo8unC6aKtlJHF8HLETmLmF+dfWiwAf+GjSjfxvzOjQCGFmJaroVwmkL9fpso6xW
xkUorSQqy3VguWyRP83XFL7jaTxbl6wAKCiFv0vWRCjjW97+uQCEmI/R/Po0xbca
+UEQzdxBt6BSoUJgQQymYTIgwoQURsPNokbKCYFL6cR71XcQ3NLN5+5KbXycgtb/
aP5jFOji+tsi38CTz63EYkMX0cZJCPrjzBx6oWaR77Bf79pjjgGgq+uQxTPN4Min
1+3KxKikR95JbXyUwyXa2Lyzz6TO6C3atGYLk/2rNSzpJuLhhJWLXfViYejUsqYA
fzWD+4JZn2QTKqN7WBhJilRXAxiqob/j3Z3LQbnwsvRT9wtrM89R9nNWHraRSIbL
LpWRk5G5eW4VugXDTwUe/JsKgFf0jRqbs5dYF+31Cus8aaXtIFFTfd+Cx9cX8s7/
KysMvibfBYcLCtdU7QfrmdgYeJ8xepjw/VsfXaA/6/P28mnuMzEdQO+8vCkUv1Oi
RZlqdXOu/FSLGkZpqjVex5/K1oScbMIw0OadUWQxjQvivnRW0atmlSDSOM5g32+I
daW0crOFsy1HX4XF2DnBHYHwIlOwThNfw6F1C1w+tXjXh+VLUsDY0I+2/8kqSghK
vKYJW/XdnRea93Rmbje2S26XNnTUW/jmCAvobIiW2Kjo8bxxzHaANt/V1KDBEEzf
CTkcugf9vGXwtAEAu+e+12jKb5zVLWR9dyuYPyDGjI68m9dr5blmv27nFZvLaN5q
kw41qipRM4gJ8wJ5JSV+qtkQMvTs+iHWI9qpfaj1LbCuDM0sNW7b95xGeLsvPTkf
fnZ0cKAoU/bXj3uJblYRgbmOW3GGa3N+Lvqq5HWG+Cs8H6X6B2vlYO1D5AQsjBGq
Rbhe/nMrhip4dUSDkdsq9coba94CqHzrkpI9QAk7ysrv7f51Wjm/2SsIGqv86Q6n
boBK9kLQYKS2pcKE+/9LLBVBCc2r8RsdfceRZSjtT5P6KM5g7yFmHSZc522GV7QQ
Ef9Fih4mMT+TMTYW/RGiAAZQO3r4PMiViIEukCgmdQdirBIjDZSjMyISMdum1ZWO
qJG2ZSV1FGSaWQEoE0gByBtv7E4N7YD32a97G4sl5he6NQVgWFELc33Zqa5tb2TS
C7tRbsRDfZq34f5fvyHsw9cE2hHv6R66RyRYpOyEKNs2xOfYbo+JXr+dNRNXMtpW
WewMMEHmbjS94pfkDPpxBucKdibuc6aUp5B7gN3YtwrQQjFcThwG5zsqN836OjWw
9URvODOYUymlm2q+Wv0vXnb436Ml6YAxmxmfrbj52OphzAcv8i+AdVmJYHLGqWOT
FJUVvBzTKpvKtxwM4+gYPIDYlgGSxjCB/pdQy3/WRas5sFWWUxZ4cKEn4jDViiqL
5SpFa1AU1d7IZuc524OqKNOyZYlPLEVd4sOIl5zIDPPIMwO94BL1Ea6kMpGSAKvz
2A/p/T1R7eU3Kf0y439vxT4BgusNWGKsoDPf0ThKwhw5wgLLFMD2BZs7pB6OmUu/
m38E7qGEuF1BCTmzbqGFW2I0nmqFt1qsPdtUeIl8FkPQDOhzr4EBQPw96SgxFTOT
aVnHcatW2H3cirOp3zKtmKRdJMrq9LLn3g5gqoX9qaBGg2Qt6ioRQUEt1dNr2pHl
Phprmt6umCO8kvuSRtLc5qyCwM+riJ0HZkxLlTBzUN8fnBp7el/06TRbWAmLYvQp
OwRSfGJUpDZ/LBxoTNVHY1WYW5HCCL1RXKfENnacH08=
`protect END_PROTECTED
