`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EETL+033VaQVqijpnk0Ejg5qtJ7IwShNkNFnb63c5cXAHbBmrDi16gqqpLkcD6rh
G3n3SmhHvj3inxuG3k3uNVrFFroU6Iupo89R/y5m74fnPA+P7owI8bfXBkgXAYsw
TIg9Oq0Jm+UnR3hkIwwEBVkK60Dfi0epnlBe2SQ0hDrkHj7Cjc3apVS7ZQ/aAb9u
eijTdIpRDVgCVsIhPdJW6vxLMlf0n8/DW53rbYwoMVy/NJsBXFK/iUccQYXdPb6h
iAuth2+XTwagLfTF8infkEqSNRQlPnvZI1Auvz/UtDPJ4ZkH1zez4+yZdUH1fQEJ
/UYm52++jb8+AmS91ZJ5ug==
`protect END_PROTECTED
