library verilog;
use verilog.vl_types.all;
entity MULT_GEN_V7_0_SEQ is
    generic(
        BRAM_ADDR_WIDTH : integer := 8;
        C_A_TYPE        : integer := 0;
        C_A_WIDTH       : integer := 16;
        C_BAAT          : integer := 2;
        C_B_CONSTANT    : integer := 0;
        C_B_TYPE        : integer := 0;
        C_B_VALUE       : string  := "0000000000000001";
        C_B_WIDTH       : integer := 16;
        C_ENABLE_RLOCS  : integer := 1;
        C_HAS_ACLR      : integer := 0;
        C_HAS_A_SIGNED  : integer := 0;
        C_HAS_B         : integer := 1;
        C_HAS_CE        : integer := 0;
        C_HAS_LOADB     : integer := 0;
        C_HAS_LOAD_DONE : integer := 0;
        C_HAS_ND        : integer := 0;
        C_HAS_O         : integer := 0;
        C_HAS_Q         : integer := 1;
        C_HAS_RDY       : integer := 0;
        C_HAS_RFD       : integer := 0;
        C_HAS_SCLR      : integer := 0;
        C_HAS_SWAPB     : integer := 0;
        C_MEM_INIT_PREFIX: string  := "mem";
        C_MEM_TYPE      : integer := 0;
        C_MULT_TYPE     : integer := 0;
        C_OUTPUT_HOLD   : integer := 0;
        C_OUT_WIDTH     : integer := 16;
        C_PIPELINE      : integer := 0;
        C_REG_A_B_INPUTS: integer := 1;
        C_SQM_TYPE      : integer := 0;
        C_STACK_ADDERS  : integer := 0;
        C_STANDALONE    : integer := 0;
        C_SYNC_ENABLE   : integer := 0;
        C_USE_LUTS      : integer := 1;
        has_q_ce        : vl_notype;
        mult_has_a_signed: vl_notype;
        mult_a_type     : vl_notype;
        mult_width      : vl_notype;
        incA            : vl_notype;
        incB            : vl_notype;
        inc             : vl_notype;
        dec             : vl_notype;
        inc_a_width     : integer := 0;
        decrement       : vl_notype;
        a_ext_width_par : vl_notype;
        a_ext_width_seq : vl_notype;
        a_ext_width     : vl_notype;
        a_w             : vl_notype;
        a_t             : vl_notype;
        b_w             : vl_notype;
        b_t             : vl_notype;
        mult18          : vl_notype;
        a_prods         : vl_notype;
        b_prods         : vl_notype;
        a_count         : vl_notype;
        b_count         : vl_notype;
        parm_numAdders  : vl_notype;
        rom_addr_width  : vl_notype;
        sig_addr_bits   : vl_notype;
        effective_op_width: vl_notype;
        a_input_width   : vl_notype;
        \mod\           : vl_notype;
        op_width        : vl_notype;
        a_width         : vl_notype;
        need_addsub     : vl_notype;
        ccm_numAdders_1 : vl_notype;
        need_0_minus_pp : vl_notype;
        ccm_numAdders   : vl_notype;
        ccm_init1       : vl_notype;
        ccm_init2       : vl_notype;
        ccm_init3       : vl_notype;
        ccm_init4       : vl_notype;
        ccm_initial_latency: vl_notype;
        add_one         : integer := 0;
        extra_cycles    : integer := 0;
        numAdders       : vl_notype;
        log             : vl_notype;
        C_LATENCY_sub   : vl_notype;
        C_LATENCY_nonseq: vl_notype;
        serial_adjust1  : vl_notype;
        serial_adjust   : vl_notype;
        blk_mem_adjust  : vl_notype;
        slicer_adjust   : integer := 0;
        reg_adjust      : vl_notype;
        pipe_adjust     : vl_notype;
        C_LATENCY_seq   : vl_notype;
        nd_adjust       : vl_notype;
        desperation     : vl_notype;
        C_LATENCY       : vl_notype;
        div_cycle       : vl_notype;
        mod_cycle       : vl_notype;
        no_of_cycles    : vl_notype;
        number_clocks   : vl_notype;
        ccm_serial      : vl_notype;
        accum_delay     : vl_notype;
        accum_sign_needed: vl_notype;
        accum_mult_width: vl_notype;
        rdy_delay       : vl_notype;
        accum_width     : vl_notype;
        accum_store_width: vl_notype;
        mult_has_rfd    : vl_notype;
        temp_offset     : vl_notype;
        temp_mult       : vl_notype;
        temp_accum      : integer := 0;
        temp_mult_out   : vl_notype;
        predelay        : vl_notype;
        rubbish         : vl_notype;
        accum_sign_pipe_rubbish: vl_notype;
        accum_sign_pipe_rubbish2: vl_notype;
        mult_signed_pipe_rubbish: vl_notype;
        mult_signed_pipe_rubbish2: vl_notype;
        intO_rubbish    : vl_notype;
        ncelab_accum_complete_low: vl_notype;
        ncelab_into_high: vl_notype;
        ncelab_rfd_pipe_select: vl_notype;
        ncelab_rfd_pipe_low: vl_notype;
        ncelab_accum_store_low: vl_notype;
        ncelab_accum_store_high: vl_notype
    );
    port(
        A               : in     vl_logic_vector;
        B               : in     vl_logic_vector;
        CLK             : in     vl_logic;
        A_SIGNED        : in     vl_logic;
        CE              : in     vl_logic;
        ACLR            : in     vl_logic;
        SCLR            : in     vl_logic;
        LOADB           : in     vl_logic;
        LOAD_DONE       : out    vl_logic;
        SWAPB           : in     vl_logic;
        RFD             : out    vl_logic;
        ND              : in     vl_logic;
        RDY             : out    vl_logic;
        O               : out    vl_logic_vector;
        Q               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BRAM_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_A_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_A_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_BAAT : constant is 1;
    attribute mti_svvh_generic_type of C_B_CONSTANT : constant is 1;
    attribute mti_svvh_generic_type of C_B_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_B_VALUE : constant is 1;
    attribute mti_svvh_generic_type of C_B_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_ENABLE_RLOCS : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ACLR : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_A_SIGNED : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_B : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_CE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_LOADB : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_LOAD_DONE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ND : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_O : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_Q : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RDY : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RFD : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SCLR : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SWAPB : constant is 1;
    attribute mti_svvh_generic_type of C_MEM_INIT_PREFIX : constant is 1;
    attribute mti_svvh_generic_type of C_MEM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_MULT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_OUTPUT_HOLD : constant is 1;
    attribute mti_svvh_generic_type of C_OUT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_PIPELINE : constant is 1;
    attribute mti_svvh_generic_type of C_REG_A_B_INPUTS : constant is 1;
    attribute mti_svvh_generic_type of C_SQM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_STACK_ADDERS : constant is 1;
    attribute mti_svvh_generic_type of C_STANDALONE : constant is 1;
    attribute mti_svvh_generic_type of C_SYNC_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of C_USE_LUTS : constant is 1;
    attribute mti_svvh_generic_type of has_q_ce : constant is 3;
    attribute mti_svvh_generic_type of mult_has_a_signed : constant is 3;
    attribute mti_svvh_generic_type of mult_a_type : constant is 3;
    attribute mti_svvh_generic_type of mult_width : constant is 3;
    attribute mti_svvh_generic_type of incA : constant is 3;
    attribute mti_svvh_generic_type of incB : constant is 3;
    attribute mti_svvh_generic_type of inc : constant is 3;
    attribute mti_svvh_generic_type of dec : constant is 3;
    attribute mti_svvh_generic_type of inc_a_width : constant is 1;
    attribute mti_svvh_generic_type of decrement : constant is 3;
    attribute mti_svvh_generic_type of a_ext_width_par : constant is 3;
    attribute mti_svvh_generic_type of a_ext_width_seq : constant is 3;
    attribute mti_svvh_generic_type of a_ext_width : constant is 3;
    attribute mti_svvh_generic_type of a_w : constant is 3;
    attribute mti_svvh_generic_type of a_t : constant is 3;
    attribute mti_svvh_generic_type of b_w : constant is 3;
    attribute mti_svvh_generic_type of b_t : constant is 3;
    attribute mti_svvh_generic_type of mult18 : constant is 3;
    attribute mti_svvh_generic_type of a_prods : constant is 3;
    attribute mti_svvh_generic_type of b_prods : constant is 3;
    attribute mti_svvh_generic_type of a_count : constant is 3;
    attribute mti_svvh_generic_type of b_count : constant is 3;
    attribute mti_svvh_generic_type of parm_numAdders : constant is 3;
    attribute mti_svvh_generic_type of rom_addr_width : constant is 3;
    attribute mti_svvh_generic_type of sig_addr_bits : constant is 3;
    attribute mti_svvh_generic_type of effective_op_width : constant is 3;
    attribute mti_svvh_generic_type of a_input_width : constant is 3;
    attribute mti_svvh_generic_type of \mod\ : constant is 3;
    attribute mti_svvh_generic_type of op_width : constant is 3;
    attribute mti_svvh_generic_type of a_width : constant is 3;
    attribute mti_svvh_generic_type of need_addsub : constant is 3;
    attribute mti_svvh_generic_type of ccm_numAdders_1 : constant is 3;
    attribute mti_svvh_generic_type of need_0_minus_pp : constant is 3;
    attribute mti_svvh_generic_type of ccm_numAdders : constant is 3;
    attribute mti_svvh_generic_type of ccm_init1 : constant is 3;
    attribute mti_svvh_generic_type of ccm_init2 : constant is 3;
    attribute mti_svvh_generic_type of ccm_init3 : constant is 3;
    attribute mti_svvh_generic_type of ccm_init4 : constant is 3;
    attribute mti_svvh_generic_type of ccm_initial_latency : constant is 3;
    attribute mti_svvh_generic_type of add_one : constant is 1;
    attribute mti_svvh_generic_type of extra_cycles : constant is 1;
    attribute mti_svvh_generic_type of numAdders : constant is 3;
    attribute mti_svvh_generic_type of log : constant is 3;
    attribute mti_svvh_generic_type of C_LATENCY_sub : constant is 3;
    attribute mti_svvh_generic_type of C_LATENCY_nonseq : constant is 3;
    attribute mti_svvh_generic_type of serial_adjust1 : constant is 3;
    attribute mti_svvh_generic_type of serial_adjust : constant is 3;
    attribute mti_svvh_generic_type of blk_mem_adjust : constant is 3;
    attribute mti_svvh_generic_type of slicer_adjust : constant is 1;
    attribute mti_svvh_generic_type of reg_adjust : constant is 3;
    attribute mti_svvh_generic_type of pipe_adjust : constant is 3;
    attribute mti_svvh_generic_type of C_LATENCY_seq : constant is 3;
    attribute mti_svvh_generic_type of nd_adjust : constant is 3;
    attribute mti_svvh_generic_type of desperation : constant is 3;
    attribute mti_svvh_generic_type of C_LATENCY : constant is 3;
    attribute mti_svvh_generic_type of div_cycle : constant is 3;
    attribute mti_svvh_generic_type of mod_cycle : constant is 3;
    attribute mti_svvh_generic_type of no_of_cycles : constant is 3;
    attribute mti_svvh_generic_type of number_clocks : constant is 3;
    attribute mti_svvh_generic_type of ccm_serial : constant is 3;
    attribute mti_svvh_generic_type of accum_delay : constant is 3;
    attribute mti_svvh_generic_type of accum_sign_needed : constant is 3;
    attribute mti_svvh_generic_type of accum_mult_width : constant is 3;
    attribute mti_svvh_generic_type of rdy_delay : constant is 3;
    attribute mti_svvh_generic_type of accum_width : constant is 3;
    attribute mti_svvh_generic_type of accum_store_width : constant is 3;
    attribute mti_svvh_generic_type of mult_has_rfd : constant is 3;
    attribute mti_svvh_generic_type of temp_offset : constant is 3;
    attribute mti_svvh_generic_type of temp_mult : constant is 3;
    attribute mti_svvh_generic_type of temp_accum : constant is 1;
    attribute mti_svvh_generic_type of temp_mult_out : constant is 3;
    attribute mti_svvh_generic_type of predelay : constant is 3;
    attribute mti_svvh_generic_type of rubbish : constant is 3;
    attribute mti_svvh_generic_type of accum_sign_pipe_rubbish : constant is 3;
    attribute mti_svvh_generic_type of accum_sign_pipe_rubbish2 : constant is 3;
    attribute mti_svvh_generic_type of mult_signed_pipe_rubbish : constant is 3;
    attribute mti_svvh_generic_type of mult_signed_pipe_rubbish2 : constant is 3;
    attribute mti_svvh_generic_type of intO_rubbish : constant is 3;
    attribute mti_svvh_generic_type of ncelab_accum_complete_low : constant is 3;
    attribute mti_svvh_generic_type of ncelab_into_high : constant is 3;
    attribute mti_svvh_generic_type of ncelab_rfd_pipe_select : constant is 3;
    attribute mti_svvh_generic_type of ncelab_rfd_pipe_low : constant is 3;
    attribute mti_svvh_generic_type of ncelab_accum_store_low : constant is 3;
    attribute mti_svvh_generic_type of ncelab_accum_store_high : constant is 3;
end MULT_GEN_V7_0_SEQ;
