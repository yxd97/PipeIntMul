`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LE+VT77HK9KUA8mGxVP/iMLrS3cyriuc5Ao1BoCh8/0cpuIsXwLqjjkh57s7W5yw
x83+G8q2yJ8xSQru8tHpcTa6TSsHXP65dnL9c2fsC4iN8rlhUi4Je30OtZVRbRon
wEiMnpF+z0pehRBr/3U2iIbMZuVw+NhngvhzmN0noVuP1YLUa21XjdyomQXf1557
RnV7qoVkXVur4Hlq3LcV60L94t19/JzN8qj5EYFloQ+QTYZdl3BpKkWBUvD1jy+7
Ly1LHEeAcgH921TMSBVJWQO0WV75aSqUEji0n2FQFMX0Uyh24LtnLw9lYu1Sv8BR
zkmrFOhe+7+ee6CFaju6p1etZxz+kBCsIoSqzA+wck5P7kdeIW8SmVXs9Sodukb6
eGJ9964cO4msaRoOvQo2Df+99FU6AEy+z/VAtSkQBBd0VW3rPsJsxCsH4IKr3xMr
X2i6KVxzDF7+e8iaRVNLutYOhdqJBhLtT6SFQPwccPSk5Rx9SGy+ZIlRB0wC90jh
d3+USiq8b7XV4jc1oOyMHys7u9G2kYr0l5ZKQ60V5KLir+/n3kj99GQ8Mf1lH8nt
eVLS3CQmworFlHionDX2i3G90xU8S4FF7sluUtsUoCzFVSksvY8BFvmQ/JvTVakB
CcmOQMi7UY1N5GmbyxaGxFSg7JSw2yd49Hz9WLA4zrYgLeGYSZnJ+IscHHr8UoQj
u28Gg5KiIkiz3p5RNbZnxqjWkDG1TWrxsJjDYUiYJ2YSv9CdEsKe0tt8JiQlfdE+
OPN/eG8/6zSx9DJ/2iA4cg==
`protect END_PROTECTED
