`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qqRjRBk+Q/4oWH8ULwmdG0/z28bpShnCiD4xfREv03WLBwVUdWVLgenYLO36V3Y
gLWXfQ5qP2cfyUHqfGjvi/tJRQymKSSRXYAd2HqoQJdQPvC9pbOwniIkMJMbGLzx
/rO+eGzMreAI8jXPrAlU8ny5ivHZn9H3yzdUYKYx+rV0B+HXFns+s0A4TlD/rkm9
gUGXQ/40lI8a+fe8aGB19l+JBeB8uBKa8ueKnkYvCGWv/y+BIdzrV07/Z4xEkuSR
`protect END_PROTECTED
