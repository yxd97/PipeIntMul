`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+vVCE3wV5ZDmpX0b/BjPaY18Vfr8XwzaILOpRXC0jV2JETUj5ads1I5YB1FzrmDr
RM+r53X2qVD6SzYH73yEiODZ5nRXygAxF+rkhJXH1jwx6pfn1avS7rZj8TrU8Vzl
vwiLSPM5haGMXlTzCsk11mHCnUFirt4bP5El8YBE4c3Fwr9BYpCtwVNE2D8pXORm
eRYqm/2/eT9WDLOj3Fasu2XA0/8Q/O1g13y1YGjzyhHMeARKaOv9umv1i+KXdn1O
jbXn9aM1jx2fXpKFEEYraC3fclXmWsyxt1jzj+bWGJSay4v8uyGMuU6CBlpqxITl
gj1oMiGs9Vn+UPmJRfSxQ7UM15ztSMbD4Ng/HqQ7DJpmnncFW+mJLYEXFLbTOVpx
bZqRLQnwGXQIrDf4N9SretZrHrp6xBj5nV7uYK+XlFar7Awxfx0nwRJEaMgzfaHP
Co8lxqk/PhcjmhClyPfLmCgaAsJJDiGtpQOkbPUdTDv2meA/6OKbAOmvTGJU0DE3
cy+/ro3xU6wiR4LtfQ/b3xUFTOG+MYu2e+uWl9xsDYmaiJGDcXx8dZjFonxlHY/U
SA/Ga8Si1IMZA0yKgq1H2Ahd5neBvvdEkoCb//JX8iA=
`protect END_PROTECTED
