`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/QVq/crJ0phJ5/MRniazIeS+kUcifV0fysLMJ5fsqkjoYjmpY1feTAsN45OcxvdV
5E+nQalC/NXqF2oYrf79vl58wrRwGxy/uDQ+6FG9Tnl0YD0C9WDsR6lKcYPnSvC4
RRDA3DVJ5+lZWYGjRg7OTcI/FinhJVshppuXB+3blrXqCjeJLC7YzqYuJO0qHDCH
cRoyOQSs3yIMejiiWji2S1GvjEL8Mrn2DkgeeSImnSXeMDRKy8NL6HtZp6ekdAB5
O5ZoAjLRV5hFpQHnmxY8Ur1rVkKXfYz/M00XFrCpiag8350HIDYDGFVP+haCqIO7
efDntNIhd/Jz/tjj0IU8WZ8EWAtYUfU33SNB+A8Lnt9IoyRBHz466wc3Tmw4SX9s
dr2O8o6onuZZhz1caADktybX77xOv0ZKLemRAYoDCWI=
`protect END_PROTECTED
