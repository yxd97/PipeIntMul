`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9d6XuybgrvInI3Jf7sgRxid+nShPAp86F/SGmh2yh7ofOSYTorswHbSZyZV7BoYG
VyPjxpqGOlq072Mot6+ozhjOTJd9jDFGReU5BpKHn4n6fELpzs1AU1K8jVkstEM/
1gnMsTnJ+9Q0z1RgCUwq3s+Pngr7xZ2g3TlWoloOsB4BUbc7AgkVtIMfGO3J5AAm
GwqhxaE0J13LO4323lhEIEyV6DriHYSueG50/vci8PKmbdDFdGbu8QUXWTX0H707
fGOLSA1iWlfTDfihBWpxzN7owlJDV7se4dihHlFw8Vry+iKBS9w3EHTljylV3w5/
6OiXTicXT0lVoO0qSkJzPfhW6Yldap1nMyhOYtgH+6e3ANiq8Tf7UyZaAOKzEQtd
Z5qTF2yzuBHFlhI65ht5grmjPyMht4GgOrpK2vBd5I+l5bRKyJBaTJLwztjRJAwb
Qrp2ZArIvhs3L50trJfTHXWcqWum2UFokhuj4BxXGLnzA9fXeHycnU36bl1QcUN9
ytyZZSID/7U71zFjpw48oqDAEFVCI6JGuYUEJnBEzvAMZwuJI6b8dONCNXSJPTb0
dfWp14FSTiJKtP+H/1hnpATLRLFVGU2dMTLgZuEmLTlHSPWbh7ViobqcR9H/AaTe
rFdO6T06DX6CDCSLtljC3haZcjjmWBqfK1uUYouxtY3Gbt77jyLvMdyylQLgV2eG
UfjTsUCf7v/oLVyfw6A3rA==
`protect END_PROTECTED
