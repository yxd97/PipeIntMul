`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YgUDGP1NgBdIr8KqFg0CJRVWZm/K3tHNsnGATn/3vV2Rzrmcb0ZxiODuk/zWllER
yD5n1iGkRXZHyJRD8OEIM/6t3P2Oq54Le6g7z4CU+ScDqkx1jGdCZvOyZ5nuGoJp
i0TIsUHb0VP589vxOShouTAnB+GaYUf2SJjHT4Ri12our3GpUiofDQAqeoTL7TvW
qEoI3oqIsA421DD06XLWBzRcbZe7ZzoLodtthtrenvRqtNbakSuazdppz7bo9SMw
p6zWSLPGMHdK4Ym9dj7dD+oWBd/ExVns7C7QRniIx56L1ILewQg9DmF7f0E+c0Rp
sPQNW+utq9bkDNq9nK/jVPTR/lW6QweCb5jOm23ok5IC5LsUF/pk6qAAhaxF+Uuw
+IApnHS4LDkTSRG4HheHK4KUjAil3HFc41bz+py1SNllNqPmPGfHLrOm+afWlylg
rvK79qWa6CRpZ1/nbLw0PMXJiU7HuBouWxVGDYDX9IBRX6rLi7Qyav+rHwt+20dt
smPFTwOFFw6Mj/DveTZmjoilE4G+5lmsa/O0IG89w/sV+HBrFjyO1Iqm+DaJeBOn
ci8PSoodoEZP012eSyjlLcUiwpYCL9VRKJrTRjDIafSLDFhNiFNIZGegCHW2k5yc
44Nyrp/Ypa4c4dGbD9Y09dg4gFKvrWP6qDRFGeYgqe21S87MDKsSJG5J6yG85Hb/
bWDAEazhHGtknZdxsrv07qGZDkv06Ad1fn78XGzvHg4cuRRxVfxqWCx7VUvhdnJg
rTj2CTDzd/vnFOrsuD2q6zdcwzufxOSpdK7Y0GyDv35nXwqawlf0obWR1nIOKMrN
x6XDvOWa2QQOzX0KGuTdle+vtv91rql/5dn/qSQxTVWSJu+PkSEMk9VAi/wsZ3Lq
qLMPgD9St6+HY2a6uCDCf/ZrOYvYImX3cwWWc5NZx01GTDA8rg3UWAVhCSYVK/p+
45UQOpAfIFD7gNlzhjZGFl/2Ac0hvWGlmpADffzUp9b9QDm2ilJ6U+XaBq3WV9tj
O8bvwtSdaOhlLRnCsnHweLDkAsPK/G42+kGA8M1AuDtz6ydpmP3L70qC0y27Avd5
m+VA7LxrGvmG76VCOXFgfNWgh3L3GHk+IBCYyrZKbmsCeDVTQjUvORM1ppNf8rXy
9819FwalaNK18S0wEzAczNpNWAszNVhwF5V6sZHJv7G9012PHPOVxYLY/+KeYgJQ
L1PCd+lfUhaFpqP1h/I7XccvHtDkRZdkyUEmyBsLhLWtkpPdi0SyZiuHn3yWrZPm
Oz9A6eTlOloadJ7Mn0wWgiwCzkEw27wLJeeeETyS/0QRH5A8rXeqFQ/Eq3X746ts
B5VhNexjcoAkhrhFWU0sZUAdBcR4LyWNC8ScrvK9GhhU5+tG9Bw1EmxUh+qkNepM
qbVPSZLAyk6fRGFJuEAdxSENfd+vWJy+DiieQ+uL7HKdDvMKmCdtDuEGwAuigWSg
ijeFoDWcVdP462wj79qq3ldhLPlc65IcKwxesK9hXoOiaGudpUcGJb/pBVj0WUmh
ffSiFeyf2peTZ/fAj5A7pnzWAJUX4heH8whJ7wwGFUQDwMOd7fSclWlTAXCA4rIa
Zyv9O7ayZPJQA4KZyO6mNu4nAcGuKJ18RykpAycXQInJpidhwju8d8cvO9IP6ZY+
+MD+fqIgFI41rSHLRl+FllyF2GV3GsTMJe/TEdwHFB44yK4eu8R5rB5JyCcgX3dB
Ug1vcgZYSZS1z+5LgQeW5mnxeiNDMI64lnUF9YEBd8TmmOCTxC85Jmsk3oAxXTKO
nhfNpKcEXDEyVei+bS14XC1xU6llODsZpH/vjyYblXg/vhLGOqVMTZ3qGli0Xktg
WREkZ/z65hdp6yApBsANTqyVv6A6CfA2XxKsbdVF3lfGrU2rwo4zFu0U0kiyh360
prq4FzZqCSk0KuPg9xdF54r0wMpRCGp0NG0Enx3WpADQekCSgCEaBG5rctC7Are6
6jtKyIDqVehSyRrG0yQp7EwXINI0jMz1sUcNKBZcMw/aPYqV7trOlfVZlx5b78lu
AY8bWyxYSb0Ov8v+eyND/gpQy5RXFD/b6zUr2veVJRZIkn9SAvkkyca9kaMgDMWF
OR/5iaCh57+6A1CIz9nKlm9kSd2Ny7blQicggwcsLzYc3+ezmtcimv6pzIXVSp5P
628eXkDivV8ljhKL9+mzQeQJFiRBLpKOYTiCXFpSEq5IY0ExiQ5iYApPfMd7jBWB
lRpRh/tuIluRnrLDtTaAfd0AbnAH86CWq1N35m7IodXEtD8UvLMaT3RbNojjfhca
1IK2M8gtEUHnIuiSSN3Pd0Bt8/CDtD64K7dAtiuoOLu6bu89RiKEWEdqb+lDLQId
2YARlSBEDa4I4edJZBh/yQmDd4xm4JND7NPc6zgfWGRKGFEG5/Dv331QhBC9Simg
eQoWBN+21g8yg2LWzTfHB/2vdwrLYmbGit6wBGbOiRqItWhOJOI26QqXd6SFwERv
KAZDFrjWtLeSNYNsvXar1cW7B/1A4dPvkFaVybyvPw+gPHdUs8VsPpEZ5NTa9Lug
QSW+WbHq0LXXcgv4jAF1TFJgWikZOf/WCfUZ/cJq0zfemcj0PV5iQJS1TonVKfQb
1i9aA7Id+QUpU5XkPQ3NqQBa3Pg+FP7sVQkuu9Ps+3JrmDHtsj328gThhGtVK29s
Qui9yxwnRl40m83PP1Kn4pGjXsaxcPfToyReBi9Jcb0ed4KAAPyWKHLfLpm18/Er
Hgk/ISaE9lu/++cpAWGJBLh2ggVqml+z7/0xrbhKASAgOJ0oCQ9u5DC69Kv93529
HJxvp11T0xTILIt2aCADmq5ncIZFwFCs3Fh2dTiuywTZHxfoX2vXe+ouutxA0fF7
FA7jkSG08pah74auqJcCHHL3as8NdrbBIeuCsCuij7PGyLvHI3W5NIf3O7oSyz5n
I5wKl8Ma62dApl95tZW7c0TLwWGqF14mPIWOecea4HT/NkUO0SZOSm47KctTGpNG
R9BjeyVCLf/5fx5rUyU8QRMmJU5PeJVmIc/7CQmmuM4KyCo0DZkZcfjSU/xx1Q4u
F1BYcC1kLHC3b3hdrSt7yS00lRDAxdmFQrXfeHW6qMqzUH05dFRvqPmTNx39o70p
tvwlJ16umR9CZHtIpBWOoRAJj7bUvMAiHpywTDF76SGvupFfUiw8vojPsZ8NfkAL
scRE36YQleFt6yweCjN9PE4sq5W8m5RpBb0lhr3unBnucl3P/5rnWaa7f/XEu0P9
gl3HcNLq7bmGjZH8PVuRm+zcQkX8nYT6kZ77xaqcefOGC7CqO5nyeZS9Fh/UapYG
aT1GDiBFNHE6Zu2uM0CaFHJiKRz8dTyqpkFWyGDt29m1y957MDug4QGYMFfe6W5n
FRvnyRsL5gfPqSguwM3WYGvbkVdUy6GmKmdHNw2pZc85WyIKuDFimewgLQ4AUvmt
x+XYFMgAD0aWG8gYsHqiUzlw6yVqwQftosw5Ks/h6aVnbnyuDswuqYaj/g7u80QY
ECCeU7/fXQ5mZ/PC2aV1zpAIoihX8mJ+4xU5DllNVaebTyBlc+RhTH3qdLBC+O7h
R6caerQR5zDfPJHg73C0QNJSV3uD0MpXOoOB679Bf3LER/lcSfuW5yx6yxUfEluJ
2FjsQUJlu+oT2i8f8jjE4iH6CVhjn0uX0rmJqqiVx7MLRML/P+2p63QPzDV47/R/
EEzQ2zJFh65Yw657EafNkAqgw8f/67r9d52or8R6srl0q8gl/Dqkv+J7GLyZt/U7
IJOskKtIlCrggefjauSV1D9z/oh/r7O8AG1m+DxrP02hlA+dQzF0MZNoR2M2tcjg
bLAOeGTCMrtKi2m9U/G/C4UsZMZ3TnoRxbsyEAd2QJM/DqbeRRN7F1X4kr7s9+UE
+skmglk7fQmvpwJBYlfyR0GkaGWwkWqnfqJZU0FDMhrz9/Q+jg859otP/M8c8/Yn
pSPqoQZWS6CHX39uc5ZQ4lRg2leXev3lTpyh31h0cKz0+EqXrbE/AdJaALLLsyJV
pm6FYbdawHF/n3MGebW2c4pIpVxhQEckd4WunBWioEylWPVkL4ay9EB2V5IZgZC2
kT4QWPYSRZXslr1u2YMW/GVO5D8eFnHoxffwhl1obHGniWKFRUnByBDyFbB/6YPa
N98nlJw163E5sSzTpv4T5HWqVqSr6za89l/+rdWQtspPTPueYm/Y0H8KAnNIPlxP
d8T8S/hV/nqF4uvG3+6H67eNFDA0LLT3kbf0EMY+73pYUkUuJi+ZDckox8ugiDXI
pqSifI5PDr6rG2QGnxdHGg==
`protect END_PROTECTED
