`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8EL01lQxzB3aK8hAFk9Ld8aq38aAxCijK6PFqyFuLXKDm8BI5AV6XD08bQOO3OZC
+m8OHW2I6xr5UKB/ueHIOg26c7VvPdLLCAV0E87MhYvcDEVjcokMA+CVZugL23u7
7bEX9OfOLsYhjuGLWXbObe+68kHVf1VbzSV1SIc4/nzRzJGRGSGP/IZ/wbDUUJGR
ItjGTNBKyFk9JxahhWx1/zDV+CkTsDasDdT6LLRN+Xba3B4A2ak7R4oq6QpdG76V
0dBSh+kMZMcyuFrnlABpRIyzqO8uQaDNnWVXoxz5qB5hzXbIA30fqrFYC9gxNdDj
HgZRyuZuSLpDmbGk+Z17Dg==
`protect END_PROTECTED
