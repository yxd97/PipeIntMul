`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eaziwuJGIJVuDXk6fzV1iAi2d3gThIVv/Rb87HWC5+wk5/U8BRFOfaRwaZBKvFZI
Y5qnAP3kHwI/ctIaedjW0XJ4ocoV8wqfqt8rYOdrV+bYDnsfsmbggglVacwzzlij
VflS//ndgJS2yKX/4O6G6IWuOoWGqPToydBcGQbgdU4zkRoq0CHpJFyg2BwPMxmp
CBuEH7WF+/FcMmKnqUeulOCsss5cKn8YJKbcPE5qjks8XXqbuBvLnENzi+q82LW3
Vi0fXx7rGlmwVJVDVASwXqEhNr7mJqBv/s30PcZgrtOviOT4E6jdujVatz/sld31
EpFerry0TaRlYPGFeGfKH6H+cF5wCz2kbIoKJiC4waByvzLMMYiLTMMuTzYReih3
fXoN0uLKZjkW3lzJGUUpl0EyLQ3pQugGEqo8wi1DJ2IJykVqo2MMUPBJxVBsZgyL
4P8RjX3H8yFUZeVykvKZYlCiI+hwW0pRix8GGthzVK1nJ5Fk1QsZhteTn7QKnk/y
vV7B2nJ3IiMHHV3hTfcJs7oOmuBqIkGJvdESL1HMToZFtt75OyVjeeyLVN/NgmHC
Jzdq0f6thtA1t8jowPaZwu/feFcfdUAbUnXJlWXwX3te/I20Cg3qbJnF0uXhyoK5
TG2j8d+5jjO9OTIw7vGNCgZaCW+CBOoadvD50LrfCuuaXlZ3H6MCVtYTVDs5SdtL
KB+fmpRxUK7uJlRnoDym/nObCRXVLH5vRwfwRHuKXBu8Wcp5sBiVaAdf0hiBwZiK
iPdDhaX58T0p2RUMx962dLd+lYcczGmfVP8EZ1fR0/uwzRW039R82CvRrLT83MoX
nekQK0pqIqjedAeVvPLZT7wRSfgSIRcuNtPAsixpXYKrgcgEOyEgjk89F25w2++s
gVcvwpKoex1YARmWLaXfJDMBkRC1CwfpWJHxFIwKJuFcB8Eo0BAQEXp4B0cyrpUY
QRhq4ogRObQ9ykXMVyulRF2r2sNjgsetf66iK1WkkG89mrsxPMZh5GyJC/5TbCZZ
vkaVigVEKV3GGT9CzzG7BxPR9zES0UA6Xo4Xe+d08K2o+akesdK85H8BXzHhVq+i
yiPk2DK7sfH+4wFPJ7uaXjRCQ9bOf0fjzdIXg7bUfMTyrBnuit37s9Q+sHiF+zMH
5y9vYNlANjjOqqAA/aA/QvvwBgqGYCS9ZK73O4RnL9PsU6MNj4JSsfyJhp4jWoth
vQ1whLsgvje3ovPrOdeGLuDMwAI3NszDVeJidIlkeaDxOPTidaCxjQkkfCnxfCsl
vp1nb9hMrQJHJd27pD59Qk0NYnJEO1btjuJER3+JTPU+lXts4Dy5X59OGYxdL9KW
AZAdiuVVrqJwNxUhhc0Oxw0/PFVXwEBhSrLGmWea7Rx+ByleSkKCJRsqdlyS+tqq
w4hj+ELtcf0K8eZpVwbVKJh8NmzTPFs3uzRcgJqeuHBQHhGSFEdDAWjz01WysbpD
LbJbRAXsolyJuTfO/W7w+EUW+lT8F2Vkzok7U/YNHowYO2KOJGyb/RQivGX0kiL6
Vx0C0i92Dw+icnoBnIzNTsHG+U1QtekWxAuc69IIGql2ApfMfY4FZuJ66ORFtTD4
msh+QcXR146kq8T26+SQ/+GemN8lIa08zyanZaCu6HOM2e2QUujdBd4w9QjI/n9E
Fqlf1W1I8Lvv64A6yvGLaj9sZFomN5CBI0SXAfUFegpx7YLT8DScAn8steeeJNiG
8vNWsJsx4kp88tZh6+r+Jnhv5DMggSy9SlsndNkN8t7U6ziHMhltTzuhLpLaj9Tu
Ez2c7AzYMO2EJy4/OZuFUTGXglV4egWUwpsACN84m1A=
`protect END_PROTECTED
