`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZvOHbtod2n/hcob5fsM9sQmJWoCHKJH8K7uWT2PR//vQX4YT9iL6KdloN/0CHec
K5Z01TL4Lw1aayGKwNd5/G4icsp7vWXjZoio1PqjijXo8+jRaRM71BF/znAmBwkA
9ctPVrFZJdmMleRI5PUNAjCUdwpUM3pT6Yvj2V7/Nb7T9Q70S4StWyoalCtg5/+y
NZiXjrs6pw9nMCGPlpsiQGzniWiN+Zzq0VGUb4zVr2hpcBv+Zv60/YXwfvgVWsCf
5YO0+bIqDO6Vcrg3l/OS7025wnUQzc+zy0fA1C6ArkmxMX6xFCY7ejGop2H95HNx
obwVyX2yXSlDi3aLaH4xN3xbA4NwmFuYyLJNS3iSRdReEVXQp0NAiDwe8XR3Jn15
Tub+JmsREdWChw37wUSYNc8+mYYJVJVAFexOwmrPwRyXed0gEz6lmMAT9TUxlr/J
`protect END_PROTECTED
