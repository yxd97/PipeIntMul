`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73H48jKH1KSZdr3KDAeR87Q0/rP8tXjd6KvgqQ/mppY1n0nA7Xam5Rvl7itOe0jI
B+HfE1f4o8kldOTRMCaxnajjNzPhwyRO3C9lXlpwzv96ENUQREWKWRlY8v44FX8X
q5MpKXcmz3gNqXK7ezFds2+DJ8T2ihYTlabkKSWO9kgRwRjrXXmJQhV89+e6r6Jd
0aAZuOz38Pc2xmv06kVeOWrtF0eC8GVWo7zreLi8pp6dxMNMI7NPAafYXZ80Ezx6
MKJxADYq5Kw9FNI/oAVHlg==
`protect END_PROTECTED
