`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JOS53T+5pQ1iC1rWlNty/mLYBTgq6pzx7MNkzMWbM1gRrNV8QnwwBuw4td2CkfoH
1uzhX4TTk3T6QgYsip02dpAFhqhZRWUZRlAZPVz33XUH1gbvHUBkwzwZd0DTzEWV
GPS6ViRnG5OJddfpNDtg+MTfRpE2UQSgEL5vOZJxkGY=
`protect END_PROTECTED
