`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BvKj4mRgOZIIQl7cpV4r4MD6HXTK9f1Fd9jJ+7O//yC/EMsjcExzx1KFdd2fgtDP
k/qLR0CCeFhIKv5GpzJHQcZppEdeINP4GrogIMTv23hQdXE2CKUK25wSq8+EfzTy
Yth4JjH6oRPTBUFCV7b2K8RpxSX99iGjfrVqd4V8+3Ak6Hv3Iht5qCn98PuGozUi
xGTSdXpKw/AsOb+11ycSWyJeVl5aVoJQvllbLOIWF+v4j6XUiaFnSIcRKDAB7bcD
X3h6Q8q82DV2/1ERcGbl0ZzPLynpISOeZR5keuCyFVsjnuIOdIL67z4+5JqOAWms
fgghA8tZQWTG0yx35/vR+AFWkVIh7v9+2TIoWe/puXNBnJaUJmXsxfJ0s3O5zYjT
cUmwAxscQsjMmXNNwFB1VRWCYB4htlP69+S/RQXXA/K54LniAeBIrRXRuyjhgeLC
kNE6mM3nhRRP29mMmAWHp5yeEvCMVXFKWNmXkAN8ctq+Gf7pOcL8wkKjO2Pi0Prz
+ooWXdSFAyhmcKJPM8+LYI6SFg9i6QbZhYC4VRU+GjxEaQID8tf4j1kmfYwB1mXP
8jr8ksms9q3dB9a/vSi0tkLvi1xDFjRl5Z1jbMA8wLoz9t89+iYWreSb2n6FH01+
CHQ634pfEPbk+yvPx9xJkfEU0lxRCHza3Vnt0o0oVfjRKO5lJD9S1nB5BaQIPdrX
vwnkPUxvgk1uqXnAuNaudVKpoWI93r8TXcHP0+TW1LLsGq4o1HfhSYfNQwz98gMc
2z0YLyD4DsoQP7A23xgD70dyPKYwyVx0jsqB8B8CBrZqnOMQAzqf8oNsmybJcC6O
Il0bArHkYsgUjOURsAjD9AMVOukej9wm1Xl/OWwthNDDccW8E1md0CcOD3+C/NBL
3Ek2d+M9HpNUBqK3TLZK3Bz3/RsyyBaWFH/1sZKRatvyZPOvQkC4U+eAlgoEnhCF
sDGMVXwt7THZLU30OiHb6fzgA+ggjrr3guBLhvvMmP3ccW3xPPBRyU5Kkm+KrAic
IoR+DFEJFTszbNov8Kr1vzyzZyRX/sTM3MaqZImZXDt8eaQgis/0naBDzRWf2mMR
KqvGtuamDJY097QGkyqGeMiKYJh6hAyqWEoKNL/sHYSUs+C3Nmyguy9PVbxjRiyT
nKFk/gNN6nNkl6M1Qw8NQ1j4VRifJib4Gw/GAFzcemI6Z+0vO932ckb7Y6QuGTIm
TltuHSk/RveVToXJ9mHXhbYSD3JJAoouDG+xJ3Tu5mviaqaYy1Qn11F7GdwooORm
yjDBPJ5neVv3O+KnyaRFwL0nG4HQlBWtb1m/D8jfM88SQh/bGc5OujukknpcUm26
EC1i5GDMcuFBmop9MD/+5iDLTHg0XEZvcxEF29sOvNX5RV1AfFlzZ7fAPBOUDSNa
7GsCDWTpsN5cisOB2kj7me2oqdSdMF6UHEI/RZV+4xCji52UDa3OEbkGZQ4MpDZs
w4GgltLWOuM9iw5desCQWkdRYgC94a7nT9NfcEp/YslGsoWho5U3igZhVSF5jqYh
Foc3ZhslWDRYmnkAXB9c6bCIqSl8R251FsOaCRF7hz1LzcVJA+PcMZriB1nvMAWI
/ET9nlCanBt3U1HiOfXQJHXkki6xJuXKb2pzb1z3wKbNnOSsrmFt8VsbgG2u/SnM
of2GlqYOE1XyO3t5eVljOUhjzg0WDNyGPAt4T65cVjqkQAU1FGIIIzYFUUgL4W2z
ZWJMMYAEU94tXcU5d/ozi5elSFDMb8PyYiwXkPbjpgC+5ifk6PUTMFKq8SqlOEn3
G7tG6ka4YXpgqsnUVuGD/rF/bTxkC6x6MpwuXxlPS5HZEJvGYSAVD6vYiNXK+IFR
bMYnW/FQLcif2xGaW5PYn+szXUV6ShM0LhI3wz/yaLOkG9qIB1dvd5wTUznIexWm
et/UpelfVaRfr1c3f6Dujzf9KPhq4bjGgEwLJ2Jb/NMdiJSSy/5/IzOuII+R+4Lb
lpLfcXqnXvJPWOh3SQZd0CVyIGtdLCVawz1kq/nYUHWMWPw44FSZo7j0yLz9KDq5
h+TTyjRNRtpe4ETLgS21ZQOd/IDzUOkqYGWZ1HxnbPO4z4RFtACpp3/5CuS8x/Yk
A9iGoCJ+zch1TZ+0Tdy8dtmTYrJ+bqcJ9fqYnaoxLu6Yf5t3tiaZWuCMxLIUlBl+
LKPfwxLiLAG8C67xP3Pl8dDOPFr9Y1elYbpqzHz4Z9A2BQSJjTpQPqCgwkOSc84G
8nIwdHiWLAi6dOhQNCepfHzH7lumD3bIl3/cJVhvRFqwIGjE8a8S1C6fwDZsSyht
4vMeYMZqVpOKcgFSH8d7u7vefVDhEcWv4KR1QDKdTc34TmA7QPR2AlsDp0sMqUPt
R1tY/ktaxkWeiEbGMXrMHN2tZlgLjaiqXpYJ576zfIidhbBRlcHNvGjlRT6g/5RD
/8X6Dzfsu2D0zahb0vGJTbGpFIlwmnsraJxZMuk8OSI4IsBqARRGu9vegniDqxCe
GLOxSbC6OQRTIOCbojtD3gSp2hV8vCEf8iAfwVK3hRAONgSuHwtD79JjdJfan7pr
DY8sOnLchTxgOAB6e5ReGrjP8B8uMDHiyC+ZA3lVaO3YxPaeOlhQZU2bcRj1a6Dk
dh3qz5UuV0Jl4PpO4VXVmT2EgLpFDBYI/n+tCcaiYxaPq94xoQhjkV/AGnyAVhft
P0gh57bRcO1nXtP/GqhBxNdVLe1+ZjnhSFpbBT3pr7pHwdF0rMNdgrP1fwVeCoTs
WP9DfchPWxFhPgIXQ+Z7YpbRUB3XQnnSzXGXttuNjrjdwc7iFTTSfrYN8wPIs+jl
U5SoIVQ6eaK+fPpm7FxujHUCkBoiC0AB9aWQnI9FZGpC3izjyjIHjIwHF9wXCt/o
ACjoLFSdik6QPeqbc5LB7Da2NGsFPqo6cn+cNBN862t+vzn/hGrgL7ULAkWjI85Z
7SEFbcMgLVJdz2DXrkkwblW7aGDOMaykF0FcHdJ6Mz9NDZaUJKJhrPquwOHLdBI6
9u48eJ1v4HbyCG32gNAU/nG7rwknSSOV7jv14RVMz9jgUkbYsFAdrisaPU027bd0
PTbp6daHjkGTiaVMeyW1Ijy4E6k9c/F3Ik/yN9YBj36kuPQ5hOMIFaabi7svtpGV
cnn/Y9azhcWUhNQIT7ZWM7/fTd6Fnnk/qbs+T+h8AqY7u+2cH4QXMwZTs2wqglyO
0N6nMAoePSUvwCwxC++2Y7uApRnoVbrzL0J6AaaQghIkj6aBAi8E3O8MVCz6Rvdb
B5cLVwk+eHsryGFfFoCd4mIne+esr8PIietBZHGYqbwFbzcOikhqfel8cm7xSIZ9
Lrzfakm79GHCT0WWQtsJ3F2ncL3CqppDkz+KJXWDKw/GNGYLszHRizw8/SzMvmdY
LDmfqzdGie3Xr5oJccwRP1N6Z0A96Lm64L5cEf01l44jgq/ZHmMKUenPLNTPoecP
1lPRI7brPf1SR+epWjQTk+J/CBNHjdqzAjfLayADiilX4uTZTAL4Uzma8LvzlMRY
ccu/6MRwChe+mKS7UsG37uVJlFwDyCz9z7u5iA6uMzE=
`protect END_PROTECTED
