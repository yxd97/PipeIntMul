`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zwi6AO3NqhEs3V/ZTz0NtV57nSw6Wi5yqw2wlzsVCae6WHoUCS/XXxTEy1Vq3kDx
0SuWyL1/mCR9l9O7I+loRXQP6GIV5iDgxi2bHbWoNoOe4I+oMhz3kEADqlckI6Ti
Cndwj4sFwy43aT8ibzQ7KYbX5fw2ntVPXAz+/8YL/7eyjkKAhqF3r+KL7eVpOAgw
aW1c/WOPHHqEqN1YJIoPkNm8vft+HzhFy6n0ULHNSamNloBZ9QtBghVyPi4dEz8D
OGNrA2FxhpOMB0IqLTNHg9NbdUfutaqcASZoiqVetAA84J5AMSVKokcNltntEbke
BaJZRQruTE/gacLnx02XzwdEtWpJ8blKp99PPS0kwq2sQR0pYcA5wF8VryflY718
3OSDKV4HrfxQHgqWzPH1MVO/I4n6KBajQYqeiGC7q5CXHhczV/KD7eD6SgwIzBpR
Mc5W+pp+XBF/0iZw3GLgY7Fm7MkqLO61Q4sG/02Pb2g=
`protect END_PROTECTED
