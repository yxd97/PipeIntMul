`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DN0EXgICg4uZTprFpej/6uwfFfm1LublRFpg63enHFgfPBOVSZ4u8F7+iMQW9sKC
N1ddglhytTa9+gjQvcuFBUqF7NV8ml+FzCGHAKL/kuKxyq9L5mNLvMXzSklxYgi7
DJ5LGrVQoz9Iaaoqh6JPlLd1pcFD7bDZcK0kHkfSoo8DqPNQ+YHqN/KIQrgig7PV
lFhHXqQnHZrzxERm952ySvtvDDlHmfG2APgzgwuuPFSh8BOPHlfc9bVmPPWucZYX
hNIpe+EhNnfB/HdOEmRvI+gAQ+lJEdP8z6DN+IcSXGX3dSqX/N3WXzKCfKRxpJiy
LY4dppHOEaSGp2Yt6nPPMFLKv2+L2bgrwe2ktBlr+HRbVtZOdjbrBfRPoloXGhFA
`protect END_PROTECTED
