`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vg+2qbU0jGYMwTRcN1rej0WF1WyJBc+5hZsdvsgaOV1DT42UTFdNB9Rs7MXDPgl
wisfprRx0zt3s5OGTy1kRaexhiw9rHT1LwXssig+LrKGH7ns5C53o1348/x9b/0p
tagDgQ86qX/xM2FZPCp/wQFylpdR3wE15lH5C3MDAr2gBAJWEhW2iYyFOtyTHRil
1zvf3g6ln+uFW1SPXLB/T5fvDr920mLOEmIoh96XIHoTzfvrO8llDpm9+cuL8UMf
+DhVXfoIEo6taxoAeLw3pyIKU0V+cTLaNkCI1HbeI80hcGgxfmmvpunI3cuWj1iC
hERcVQvkljkCjB7pnn/i/c7eMMZ235Irl6UUFQVuHu/NvCFZl3RppNQSdbadGA1g
AxJYZtTxh2Mnigv4QO7R5VM0HA+JVREJp3/oc6bfsq2BvPEIRDx5BJ81saWlIi/B
1FGOVZopYjtiHZFKUg+ukxkLzOdsvxl3LKmlBr2X5kWVbrHVPN9DB8+juukuVehQ
rvExvDV4S/esJAr9XDM9Eg==
`protect END_PROTECTED
