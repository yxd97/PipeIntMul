`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUOz3SGc3rKzV5jVOMTBIMi/a9EINHH2eXk0E6g0yv7NvzNv7MXFTEa75vLP8ALn
hC5bG4X4XMdumRAzKN1sG/XXEMVRqsBwaHThz4r7Gw3CTrZlGu9txE1sUYuPwvs8
H/0YRDSWEqz7CAxU0manlUor2SpCH9SOYHz5wB27MYABYoUhvAs4Baa0ZHswnb74
1vE2ax3PH9nmMLGUFMgTZ3ocrgbPKkJ7IGwB4anhpI6k4XrpUzVDmaS2QbRKe2fZ
NghDfwKSMfw2eHGFFv45bTgcckybqqWStGwTP5h9ZMBzdG5gy+DQwEYk5KKC9MJh
ycOAxW0Xo59+3ed7g0McDg==
`protect END_PROTECTED
