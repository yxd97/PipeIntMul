`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OpE+whc1CEOz45kbXwtzlIC8SiEsflrtmtGM9GTUVeQq8MelASL/27ZyCURSBsaT
i2Di8EEZolkQRXvCQRB4sLsql/RYepLTr5kEOlGxOGL7fCyA/ZJzQbs73cZTOwgp
7bSXTU4bmFlrG2WKfZAMtedley9p7g2v0z1jjKoCZAUkztPain9SVaWdtu3AnHmB
kt0Lgvf40+Ex91ArkLeRO7sfbOR5X2ikY9xR0ife82CV7s68oYP8Z7EUaV1juHuk
KEej2Far0g7wu6PQ1EnGw9yplYDSlG3KuLWoJji/b7WByozHt6hXIy741lVJ1nr8
xzaTSk9snOKo0QUnWL6wBgA1kx90AQPn6iA1sDQ2EWqBXxuRIw3QeikWvD4jwu6W
LCddl/q2PCjkQ8SFIOKD9bt709HLxXVRSnkzIerLXzNOiT6TmATeYph3HU93TMj4
ha0AQ3GFMwwKBcayIfdK/cpYlkz9Wb1bC1Ysq7R3mmgdSXmGKyBMboxYKQuwGB3z
uf8TI1+ilUMi1wZSoWWAxjDHMdBKk4g/Gs9Xai2lXsw9ViyHUxnMMGqsuKNaATYw
L6dJXd3rY/svq25xh3W3qXWsDWinEfhm14FQ4OAudAdXmgLXTfYvT/+Q1Kne+TCa
/p6DsSMZ8jUynqMz6Zdw1Dq7mWX+12hSWdXdNNk5xeySukhek3dca8ATLb6fJPlX
wlNl+2L5PTGmZmNmLQouJ3oWrBAEjz7LeqXahtd5TPFwUnsEB4BAHgdj1zcrxO8Z
bI8q2z3qYFIO5gE+ak/VaRlWmW2ud+c4Vhc5CZstmm6UZDys2JOwMcryRghQS/J+
58vVO6An0Wu3OQG9U+fhXOTm3BEBysIKDkgO1/xYu/OTP31Gtrv0WfRN4YEe/6Nj
5/eg83GzjxmGMhP70+w3u/vpNbuZ93nRUC4nFj1u7h9iIyTP4GhjQI0l+xKuPk1b
UyzMVWLSQlfwjdf92Y04ng==
`protect END_PROTECTED
