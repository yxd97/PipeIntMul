`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6eDMwt4sll14GDUPYeCbbnFst35fsWwaxkfx9Pt1MESgXtr9TuHgaid5JNN5ng8
XqyKm6H8VI+svR3DD2n+gzevES5vrYSPo+OudRjbzIfIBnhGJqkGFSnYFoH2fPJq
Y3KAR9Ya+p4PGAdmK3sa0EnJWo9ZFPpQgiOn0xp54jScK68qPWAZFT+kLWCjkGty
TtRVPW1DE6N4F7hfxigXBC7pWvKCvVT5Fg+VlzNMW+eDxno5mT6mK2zC8uR13SNs
/PaFL3KD1hAFYoQvfPbCn0kwlJmMdJ7L4mxkPfSrBtQaJROVyr5rpeFDt14NFfaz
2l61zn0JTUCd+5ebL7fN187QZ+dKeNAXZJAA1HdLCnd8VG2cyJncNcuWxnGzf+Ey
`protect END_PROTECTED
