`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6z+BjOsBmp8b/01qbCqDLXE8vfUagT2w5C4RmwgOhIUZuM4dkIIuxUKcprZIHCzX
KIcmppg5/XOOP2zcyhOaSqqletsFMpsy271VYZCF3/boV4bY/iej/p7pXUMs8m79
HDz1UolFE/Z+4ND7WTtBYTy87nF8dMBSf3A5MTJpGFRohBZxYKCvlSpbvHhN3qAB
8A8GY+SkHoG7DHBZb6wOrdWdZ1ea6Kc8v4L19IeegvH7UCj0x6Sq6nwPzuW7sCei
qAp1vGJi5g3DqV4zXgdROjooXRZZHkNLlDSP68QQjDNM7Is6CBrpue1RPlyJ7afn
y957h9GVdTdmBszyZKc46umhmpcOqjKE926t956J+7yiolL91Zhrqtjb6Z3IQ2iQ
ABC/6epqkXbqCnbPL4xSiXI4Omhm8pDOfkjzbgtHUL1QlJ8fejEl4wqArMwba+/i
FFP+z5I9IIJ8dkk7j2vQdIGyEKHc5QRPsL+oSSAzYWvy+y4tPHIDPAhZ+rqIaewD
IgihfFGA+I4BKeoaiqJSorgP8XRoxRP9jz58dzp7czAEgz1sw9kYoClCuBCsNEfD
raXCXY773OhoFj0ozDc8c8LgOTCuC3WLREqsmHIWAgiYGkyqJKGY0+1vnmkY6jP+
1yVkCLppWb/LPWILFlA9GbeNqVtvDU0NRuEKYomF/KMw0R8jkBpXVQHA9xmhGB/U
69qrqBcUrbLpc8+VvW5d1GS7gyVrYp9Pzj45OSFplLTafrlkVvCMdkeA7VzFsC7o
0ZZ4IquLf+MJu+tE52Tiw4y6jH76KatHJIFuYCTdYoSmixLqan7sJX/7F1ou84o9
VMzpO4kIbkTZhJ8Jws3X0A9VShwwiip+3AuSy8Hga+VmE/GfG47iz13nZ1gA95gk
gGqmhsbdGXAZmhhVIMjmXTKA0F63p4n2GGx9jY2y960=
`protect END_PROTECTED
