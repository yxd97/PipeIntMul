`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLmo5NRP1JtHsUe9l8mKXF5aIF7GlHxLWb4dZFyk0OKHgIFd/wn2LJIzDfBMjMDr
nr5BcdwJcyu0OEJPywvVc7G/cJfc1IbZoYWXCv2PG10YKwp6qVKg+RPNC3G8ty0t
O799x+yzZAkDdMKLL1CedEbuQ4tpj6PQhDlxUxrSFgG4Ww6CQr6EpH84m7hySI2C
FeeS93gwbIhWedU2cNvVc84EI2vcGHmMEGKBOWwnZoVIVrjnOxMrXxRoDwVQPU4y
YwkK3d8kNxYtB1Ob/mlX3cXny3YYHM8tvC7eljCp9f0leAf/5i6N3GYROQRN9H2V
RnTKipZyV3yEzWKGWKvarnWIh1YeXlzT0dl1cPvlfvM=
`protect END_PROTECTED
