`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MM83F/y9QYyLnUf03xvUUsoXZ/zxqFoGBr4IMjmKZh9etpls7tM18RXBEfbrBs7w
OTaGiAKbeDBB/wZrh4KaCwxWDuB2FoFwLSlxJ4TZnvUcduTJLHBEI73Y9EF4fa8d
RHDy3XrsmHDwsdd+TnRSMI9zdsWpnARyotOyFBmRY3VJDNhBPVJ+pSWrX5gRI2Bi
owGepgRovxnJ05o6qBlxW5PL2G9OQRUnoiF9oJHGtdUhnPXVC4+MxJPdqla3IXpA
3sXmN87mv59t713pioHaVgZI9qQ7+Ei3+li67Xm4G+fc81yC1reJoSBqwBjWIiHP
8ur+w4rQzu5DfsycwhDE+4MbXqKW6/c9Oz1AFJsMvPlxoysMRfZ3j903ZwTRy8hR
vy69+Way2hlgl36XLVH9744cFr1wM6yOITgjuMrfqmCRLQBPfhlTXzi3gcOAmg/2
bAPLvl/9wQnMw0WNTySFHWHeNncvg/xff1O4T+R03sO44PEgh2qoVIONDS7v2xvV
LDWmEdLYUc/riDbZk0/tuk9S1ZL69ddQugiu6xSgEqZpe0P25KbAsu6VYz1t5rvA
PmjrMbu7MGArIU+oYOtpB43Y0MOQHWhxUii+ItuvHiKblEVMswISAxHm3rJMjr0i
pPD4G+Tvyu/+wbYvgErmLY5hilPH7h8QxM8u/+lkrR5eBH+BPJQzCuw20x0dTcEW
ihz4DQ/X5taVIw6MOrVYpA==
`protect END_PROTECTED
