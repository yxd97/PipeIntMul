`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8nKUGS/lNCKlxPUKVz9HkddmS13x7ZkXcbpnyiKZc6X5b9ecSV31oxZOUJHogok
yGNTCU6NycLRB1HfCbqyvCa+WIXTwYkbVcusDRcbmQbjQ1Wh7l7H6j6ncu9iOOBr
ghvJOK/p22qMgwDA6Do8sNMAPtsDPti1IFZoIsq+sj9r9PQJ7ZOZzd2MSlsXn2Ar
AZBtgnK+jbjw5dX4MrUINwLJ8WDBMmcpT4bZSPmbQut9kx4oMUvy4LkSOxrFCT0S
Vo1G13mF6u82Cpjw9HRWJi+ITIAoYcEWDy5DO/0YmwA8Ipk+1NcIX/3SFPr+HmFa
mzufoDKJ6nVK13irgwC1XXkIfwFm99vkhT3GDrtd/9GMnEjBGALs8QsMpAaM5N6g
YkTPZpWsEIAP3PIJnzhrIb2Dfz1Q4NV4YEDpI19eB7ige7+hNL67pSzXT9Zuy/Uv
NZgZQr7PCVx1EQGGlNAzP9+EP3SAC694TaBLXskX0h8WJN6XltJ5psxGOXWTqcrc
QZD8j9gRf13vxGtF74ssTdSP9xw50nGumzf6qXkG/xIuJ6H5keyhX6ZiCEgtrhlW
TfcEBuZ4rxq8XblATceTIx0ifrQiY8b7COZlxVbZNQxxc0YPcCGmKylxS3D+D/gI
QTBscUcUL1AZaI0BdaYDF2Fh1De/wheQjNjCp1wJL6wLqaboSKI/4QpGhlLG/rcX
hxYRlGNZhngtLSBG9R76RG3asyFUTaaV369S0AapA4XfKruCbRvqbnMhMzGi3VIp
V9+bjMMLzrt+MNceM9H37lE0RC5KzdpFzzSHMsivNgbWBbtLfQEYIuNcZ804PYNR
UYdGG+zlDz5VjT+87yQDsT3hpHUKH8WqiRE7jZlXXze66uEmA9/KOzCI9wuAUb1k
y4Q7HZKP/qmHbKlJ8uenBb6YFJKn+R/oXMLyqWW1eN7uQukMj2wwGHRCXb9RDfeu
wp2LacbFQeZq5RD5K2ZYxSET3tRQ2mVqNkw9tHw1A5pn0JecKv0P+U0INXedqm89
fqu2VgTKIjdB/XHE8+iSjO1fdZ546YW0/bU2jbPvqI1x/rLjaxFEhkHIjuHHUSzF
/7oXnuGOePjQu/rPS2WBcbQb+BiQK5EjBt/TXZVT3hVwfyMvLyPYDeoV6XTOBvr8
Wymo0RW4YWqWLhVCpuvJzCVdj6LY4/RhURdxV4tX8U9l6iL7M95Nirxq2Cl7kONA
UA/UOOAaXveMaOFHNOI7j/2GK2rSvy/a5Yu1L9VXHC73CkAPJfpxa7XXxdjo51bK
YP+NTb7MeyPqTfO0Woir+Unlxuhqzr0pQC88O8ZOp5n+xz/3n8hQ5lWMpCh7VT4B
J12fL18KJerHMMSY2SaUXmJ0kappAa+Yma9ikqQ2pxA+DSVFZ9TNs8kn5N3wo+E1
SfvkuX3DKK9AdZX2JFIYtkkYjTTsnY/j3tMI+sNmDfNAHwLsLcvROARFVrS7Oju2
170TlB6OOb74es00kffsZ85Pn5tVHmsV2t3bb78vmdShiX7Phk6YKUICnBoWQeX8
/oB8eVZ1J2tdoG9Abn1B4wEIeNxoDlH0DAeftkpGfO43/L6heVVOOkcMpmfqJ2GY
M08AB3n8hCJC+dPra02j5RMUIc/TeA9I0VUBg+G25FfNLtOP9IePXpp6UVM//ltA
oaCQ6WntEBB/IQjggV0EwxIN7vsqNVeZDd0CVfXe3Q5j8zMB0gLDF4OtoDbU8XbY
KAQ2WghtZVY/jQnVzAy1ZitcKy+bqj+gxkt1XsEyCD6lmGqK5d1kwXYd4UkcGnSC
gwD0tK2uqc8yQAuFZOo9pmk9HSKkgAIgXUVvZJ9bsDGBTiKf8DZCefYV7i3gng8j
cv5i9nUFedp5wIGAFKU0PEyZhGz2vCEBbGMNSgg/YGw+J0uIBk/F29YxguocAC/L
udADxBop7AkVnE6NE09vy0hUOiJJxRT/I6S7VhAyCdriuKhQED+Hvvr9z0G34fOZ
SWOb2r91BA2IgUVp1GAhLi6EKap773HvoDQc5/MqPE3cuPqt1Q2VGtgWvQEkdciQ
22RRtcwAQ0H/a8AamhetQlBbWV30vpg0skgqUdtmUBWPZrM8IUc4aWBwva+NKEWj
oP+F8QG+jxtCCyBk/FlnJe4CbuKEJYm0FcXgx6WWdQgvJMWo9Ogx+8CC4KVWkcay
sB7U7xHSnnXP5zvQrc8oQI9La1a8Vot8Emm3abnGSFLNhLGSUiRry8mu7E3ea+Ha
/GQyn6yb9aMqOiqLSV3GQrNuSUkpfuPe/6S7cd22rPuHkEvHMMq6/w9f/iLODd7A
PYPY69E6j1sGxVhnGqPO3fs7dEJxVVshPEkXLChNwppvxolDZE34PIdBtniMKfS0
8rh+BdUsp66Kx2GQ+DFCvueJpR1fny6BcRwX9syaC6igA0Prh9NbEbRaUfHYkWwi
H3wEWGQG3yKiJN9nZfTT0BO/Xi+ub5tDcn1ex7Du6Y/LcRs3w+MJJyG8Gys8WgtQ
nJV5s07BNjSNsD6IX5sqj4V2VUisxcIsTpDLgsFzEdKWN9ytAUDdyxtCR2nC3CWC
e/pfttqcBDW8MDn955hhRAIN0GFmYsljF89+Y0JsZuxm8oJj5zaB+Dov0PrH/eVM
VeLlYHM8smRKp6WSEEb9sGZN/CXuVKIvUYsBDOwBVPzRQDhme5zqQCvluKDsUvl1
8MtGCnFglDqmpDFp5Rm4bzi7zRnKF/d6/PnpOvF5VIBiQFZeD2rNoQ5+f75l/Zhr
24WqzlENbSaCEkDv1xqawEsczhL840mIEf7yzsx5LMXB81xF6fiMkFdG3s0C2/iW
l5AwM4CbmErFIMYr1Gjddl0CXIJbwbGBL1umsmy4Rap9dMDMGTv65HQ7AU4gasPI
5e5Z8n70bFh95NXgjhzlimnZFG7ikM0x5VsAYP1s4yF8IHS2xBmr0XhkixvICv2z
TecX7WDyfpcI2waXgN67/9AGOrVANcaoGk3F/gpZff5XV1LCfg6d4w1fFSas4bjz
RdMEYmW/Zinonqzhwt742YYUbeEbbWJW4R60eBHSu0VwQLcZrGLLHDPCeqviuMd2
WacUePj+m9OUWmOjQa59kZH6iMEc6EuLoPCuiuFyT3qAWeJLEQpr/MsWAKFvQVB4
s/5ad/Dt11+g0HZFPZoIG/nsXsUcmJgDOq7TdXO7qrMFvtrSduegDSgxdnHDXBd4
j7ThqgXoy7WMbV5kBxDjiLrazAM/UI/zDh9bA3g5ZLFPm9DIjOVV2MoYIhckk/Qz
OSQXWWbNZDt30gHNUHwePcAzka7RHG0aBGcB/IQwDCrW1N9ja5hspySV7uH/1jCL
BdtcvBUibHHoH0s3VOqNmBS4N4hNWIIah8HmQHwA+TqWPO5ADhu3WU4sLNGAtQDm
9jpTeRBJbBWXc2pu0Scb9l5psel9P7V3YnCsFJey8SyOVB/lfCbhbVRH79bfk56l
dZd2k9DRKlPoE66lR3WRVu0Kr2yNoaggOjPiPkAvofPjVBJAZ5X0kyi4q2XeJmt4
lLKpYAVCmiZCqCXuItmqytGfQrtcic1Mblet4GP1uJrEpkSFpiXqf3NQwWSgES3z
NbDhtMA8xSkGapDjEnmiAESx7SUK88QRfarlINVNA8BZ/Z1yBfyUKy/eJ4cjm0OV
jKui/7MEbort+YdKEiVPwNGZob/K2gvV7t8E9W7GOO3TMba8xmvTtpLF/c52bJ9s
UKo2dHIVhVIk9KEb10Kmd/xuRVeQwKiCHoOnxs+rmJeDFqazFFdKL5hXYDx5PoMn
vlyNK0ogBLZiw+Dw6jhSMaA/WfNHRbQ2FwzVL7q/tZcc9DIvmnCKJASUah6VX/dz
3Cx33dcCXRbVGEbmrR8Ee7XKZt8rLIplvxkK6pIG2S07Ii6HLf5mInQJ7ILTYirz
GvYMSAfYPPfQnQvTLuDHgPyFM8fe/499YhQOtE8V9ZxDJvtjvuR0Pns267UmJbNK
0MpXxC1My3qPMxHtUmnpea0CSnbdc6Q984YhIdsTfZNkOPvtGPDovKjOb5ClgmkR
kNbLSOblkOlsMYD5LEhq6jQjYpwar6f9fgTseLYf51JuJ913XoL4h7ePaTq44k2C
fvw9ELWJTMeMoj6HbqK/GDVw7rmaJQXteZPgwGqYG+6FrehulWMspbMF6l5KXkq4
jYezugh2GgF9zmPwKlEuCamAyljA1o04bbFSmu9cOii+zFO8KvTD7JegmacZMk9B
tjyCrNEHVL7IN+OoTkolXyQrev0OaTusxisJ75ZA9neFAT2ouK2RhpU+tTQ4rsjQ
yITjIfg6r0iPTc0j/DkQEzhP8A9BEOa7/D7VB/KH4T6WfjWguh+whBwPShr0Bbk7
pxc+C2NubiscNemKR3ZYxhCJjS1DC/yiOV1C/mq9OVNN437hiqYwNWeKRctH8sTJ
VjV0j3hgOz2G3hzk65BOX4qK61zbX6awzNsKEgxlIyfxa/WG5JnEgTGEiLDBVY5z
56e2Ed5Cl5hCShYz5PtvKEPvbXdtYVOnpfZoXxBcKx3/bD1p499noFmT/0cbrAHD
fMJR5q2l/Ue3TkSowZQfmtRgWJ6iJXkdyUrRh+9h4jtEsVFbO8mwET5IezOoJy+G
zDevB8Z+UoBavBvJapW9xAzNMoZqVZO1c58+3ct4DOnjb1hfXE96uHYd3w1Gyxpc
p/HoJVt6crlEugBt0AQCu2KsfB9/WmEGaE5P7dwTtIZ/molEoZ2RjBtXnDJVqRAB
K098Wr0oN4wka+aJ1XdEJAi+7KXGQPdzv7b2IYfif/VQn8fHACH20cNFluRcCecT
HqbxxfvmjRGxBVIeRELDO12AOkEbbnElCbYKY6f0PK0xCWMtPRa26UHLxXLviyc2
LuUgbxVP6sz8FfFIcs6gSRJRAKYx9A3zPw6ezzXAtMNufUVPFvVhF7xvmKc9SSqx
syNzIkWb8DrI3UlOw3pgiP2mF5g7NH+sYMFivH1F9wfWEsQDHoJFFS0MTXK2GXvu
RsTVdjwtPZK6zGKvkGNj68/JpqFL2yTdpHpaNVpBsqEvu9HtyB26Kw8dEQyNawx8
ieewfYG5QQJC6vMxXUR4YgyOmiGcMdZ1HkNgMQduCzRUsmB/UkezHd6SYE1i8kma
m5a+BTjNz958a+jwAMNsdEXcYrFo6Ny0IMnV/q+jrLhJxHmq9JL37BzVeFMiVzs3
FiLR2EwpLdTkMPaiG/TcPgb5jT+4ifTFSRjFESR3KrNMamS0Stxp8cE7thV1b60o
R9f71GJWZ8M3deHvMTl32FHTLphXJG1GsC6DvXZcaSC1jF7bv2LBZFxpYBR/Sfdb
rDq6YQ3X487G3zvUWZ5iFE3Fp5cSuhreibsXkqGPUEFGGj+jlA9SPFAwjDgSzztg
9UIVCwsiHsqTli6pWt7hHPXY6oO0CVK1Uicz1sMyXlpOxM+syRCJT0jpp7pCxlPQ
8rce8ep7zXRo1IZvmewdMiI+tD9stARQvEeKbJ4JkU+IuJhF8ZkO/xpSDyGDMwTF
5AlyHfkKuJH3mlouumG92qchvrL6CcNws48EtosK/kGEvN7P2wWguziyjc8Uqy7A
qHo8hcb08FIEwEzjQ+VMPjC3cFo47aKsUToErMJMEraqj+0PpBE1/1cxtjKHhFI1
0jgsmgu2VrV+HEEtE9bn2nfwyoBa9ebI0pWvN4uyed79taRkfo+eQqjt6KEJGOcb
ZFXnbpVjHV0E3pkAqDT8OKUMbaAYZPueP+SPyJt1PXjxdgQv/hcb0itiSqt7AxqU
S7HGnnetKeZlib7xdikaKmqOSJs2h5a9ZG6KlxWQdeqSm+OIOI0Z+QJS8z7jxAiI
d+eF3a/j26NuPqtzhTTCCT31x38/Obebtj3TzeNG8Yptr8a1XfzQ+IkCSatWjGhL
BnHvpKlJa8DwIcKwZeonDPmUA/vr5H+TNEidBNmb01UpSCgthhjTOkOy4IUiyuh+
X2ci/IilAuCW1DKR0Dak6V68+ZhBFspkfAOF9PGLrLoMguqU7zv0IORNIBrG3v44
jPBdZ7OhCNZeZqHiZsRBM7yex98EB9iaBam8FfyFycyVF4cpDw6hwQcvUThGh5jb
iErn7oMgzkKjKqa/INZs7/zj9tJlcQDCdAw3trkszASiZKYJXOuW2FBE/sn8tKBx
V/TYumU/rSBxR9rUt4hZ8sNy/2iznb6emPkIWXfcekryXw4GMw2klijSKJdMwtex
4ae565iiqfleGfIc4VaF04ZuANWicjhawmKnS26r+BbKaIufAszoJ+CXEb+tJ8lh
GxTuI4DCy3DD0Z7jmLYnz88TRF/yCi40vKGG3xrOY9gvI0l1M4QcNcuiGNddxs5X
9U/d01yJ95iH4EuwpxE+gNZDDIAbwFS3OctgBqmBYxfCctdXy+Teh9hfd574rV50
v44BpBv9UaT1KzvMEVD0rLpTAmqsqLV8sb43kKwJTgotJHxSQYcxOPz3bYlBtzcn
uMrMmQg2DpEXCdCDMWxNA/d1kHR1y+KYJAqrIkNB30mQo9dAnfOD39nSnh2WqkYw
RFTeGhMo1a2EyVktsEXrItc3EqbSlYjyZAmNRZvhhvvSn+n2+tvGovza9ngq0Tpq
rZn3mnNxgnMOltxiTE7sWQUyLWaPVsAfujZSqCbgK79zuMn8ZP3qWRGRzugk8RYS
RVIzpm827SUEvvhX44d7pyS8co8mdj6/wp2qjhl5hfh8sAl9kpIu/Co4aqh0RVOV
esphjjx+rZ3iDZBlThVJZuiyWL+IofirfG//1ejMziwNmehK4zgK9hR4VT1puye6
Yw36e3bE12HFF0tboha++VEtFLxunuYyAKrmAWoeaFBqxT4QzjcSMsIrZLvqEMTD
DxeFHGEfxIG1Vl3uHLBgTHVhsEMEzkQhogSn3ax6lKrFzC6GRWL04SiaoDhohaLx
3DR2wBGhjvjnuYkOJiEOJNzjP4JOKWgiwdJv1fmqpyLl+j0Yg6UJ7p8tSlI96F4A
K1/im8ibpoBLAXETUlqjHdbxwp/HsigqWJnfJtAuk33apkHluh5fIm7IFevtIUfw
v9uBPbcJsR3xt1wDaxSSSu7u+WLFQmK99oROJ5FURIE40cKugn9EBSPQ1dn23ikT
n8BI6vKVi/+E0lfX5DpXUvb/3m5SbI94RfmFrRZ8DM4d4HaFBaKd5rwhn/OUDEay
WyO00FqtNKqq0junnI0GqGWp969xJvVo+lXNiN2hCNtp6ktl+/IcxUpQdlXUO74B
EION3l+c8idxy7yiQCcMXywr3Eu0sfR3Wezv+1D7zHNlbr0JZzy3nREInZTOW030
vu9E8Wy/18jWnihfbh+jsXhxqvzfWsBkqC1++J5KVURyoyaAPSurxT9dmtc4ww/B
csVeVXlC5x2SJS/6LELV8M741trLV7NnMMM4/BEeI9tzRARWqbjyYmdnpdH2cNvM
IVoXibQCoVibzWolpZnfcOYb6XsrN6f26fIxRBS/a3CHYcHRdUgiWRdEgWEF/g+u
IEEF99xr3LQvnF5KxA/9rU854ip3vjLOpJZ51qMRTo5hml611tJezozDXT1cGTz+
8Solkos0dtVajvXIsR/tlpCZGH9m+OXQsgIhUt+3u1Nl8umgZ4gpFhImex+RcfNl
J9e5Cpbq3LvJYQU7yV4SpWy7cmtyp6IV+TwiYA7BCvd3U2zyQBYznOnLHVb+E1Gq
COMR+7iJuwOSqBQ/k2wY+XuAES6v+NhEMzovA5MzyPOW25MHe01xyuToI3jsO6qw
4YLQZzDqoj0BG+o7wB9I98H52mUPyEHncQAs1se1w5NO57JlFbiTsICeN5yil2hP
kEhJiYRJ9l3u/rqp2BXn48x8f3dHxEeQYgAkp9AoDsf9mYb4Au2gLWfdxQ8kJHMn
QJULRrB1lCinNvH/RUEjQNGOCsxFIf8eOGVluedXJScG/4yCo9MSEJl6iAQ/jnaq
PT3cxn1VRMpigYgTARhgO/xq0uea5/dE9ZY4eTC8liTSrfDaDHxH+Y0HSslxIuzR
pzpR88N1Iyg6EHBi9HPRsf/aY5XRJyVqATQ1OAIwWdqVCy2K0ToZgewMQtT/Ahqf
7rlbnByZmaQrTUSZs6atmqdyqDCSSsp8pYwAMgwHW1hM37O2gKc8rzc0z+6PnZ1G
80dB6BK5JIRL0TgDCurm5uu5Vpl9mMiz2fkLIqFVvz61q3IIFPJoumVrxs0UwuGO
RgZ7Qar4J2her9zKA0l5N7mzVyQJ6mREO/8p8CiUojTlHfXfSrOpyg11q4l73kIV
IOVXrXpCNSJbPdeFm+ztwHGwmN1+5IW0onXhIxx4oAR3CB1KkcJrL/PQlFWJM9g9
AIOi9fCIxBYyk+0Y6VEvfl15ZtcWOfmk1ZTwWj6t9YCax0Vug7uY3Vabcpc4OHtg
o1nYivqO9bZ7qpvihrwoFyCH0MqRl8hVVCM+DqAoDEeJoPw25xPYQ+ZuSCR4krN4
BcZLM3A/FrkJKNnjwbTufyRB4uwv0a69dhqvPe/91+Vmo0ZH2FxkEwnsZNmbDtiZ
lCnO73j/C9Kpv5W6KTY6LFPraA8Jw3qR3B44aDO528JJgt5pFeYIEXnsgKL53zr5
yduERZqExY4tUJ8yEoPblZtVDEOoCNis3HRJDoG+Mx24t2zDYSjLRNI7yW4323dW
aTVuSAMrwOSDD+Jpjowlw20Zpro1v54UE/TN5cS5ItcH/5m97cNrih5kkuy4a2gh
GJrD1MoM1fRRqlbDNTpWSdF+QfB7o7cNthSvIjEp8x7L/5ha6s3FsY6Kj9+NTbUo
9a83/Vlx3Yznx1pJ9a3qejR5Et0g8aBupVMPpBnwmOB0ZqsUXocwDoWakATUNhWk
yuZETikUpRatnaJWFOpuqJbVwYuMpoNUj3BqWLlnEzN9MGRXeJmZmyFLN6Wxsc8e
z/bhhCS+d7c1wdaPlIDBGQS0rmqNduClxkCQqrCC8LAF9RbtSLRVF9o1/4eWM80Z
dibJTcVUES/tL+BEfK0FuPLD/PeALHNSl0bYqF7tLCE6V1IyBafynzRO3GLEXKId
GfMAUAc5POL19bzEuKG4yALsDpuouoWGJ3vmPmd444RIcqcchrbBI9Ru/2MmFoCA
D1TZTwvqxNXH9mVnHgw7RL4jrlg28L52k/7bYs2+63SfkDVY+xdo9YCd0m6VY31U
Oh2MXSRxSPUXFQAT2Q7I3pq9f2JB/VbiQoF0E0bQ/f+qEyp5UpFUMHbAZy6V1go6
Ogh5UFmkZZTsJ5zemfaNVAuOIR3yEkVLR6YuaCDCZcZM5Ej7TDaQG4g0Ckh4kHJv
GTSpAH+hw1qP2qvaPngjUfcAprnYSKwTe/ITWfnbMgncfrCobtXCAx4vqKQ6CtJT
XCYDBgTNoL7KjScJFs7gPE294aDy0z+etjel6SahYBOO1CJ2PXiQpQjfql3A1sTh
r9/peCSj+vwtN6hdELH5mmsqTeBBTdAQVCspGM7REPbkxzYvt9NZAaiutkHj3jr3
KruL7AOzW30U20S/eic85m4fWmj3+ufxlZKXNZ6SeHMOXCy5NlmmaVEKmOzJL463
ZvOwWg29cspcjz1LmNCnusBOBngvxDiDFJWJ4nhTUU7ikQLRlDqoeasezz8TrNCo
GiwdGIZXX5o7X7j5ssw4Y/wxqp2ZInyc4q1M8hiZxE97ZXQ7j+npS3/0XP+Jj9T7
rMEzzkVvIv2wTa27f1u+CREiQv886eyBEqgRSFhtT/tPEicMBnIdiy9VEYQUFrvJ
gjiUSYpWmLiB9VadqRh0926pPliEq904GHcBnmdfpExDWGdx5LtIUda9+nw6O9PZ
fv0LMIS2G+FexKCaLUQ8jFvRS5yu1ztHRal22+rRnhhFkCalwu6iw3qjkpce3kqI
gbRBmodcrx0BvGO0cIrOHIHHIjaaL0gMok4SWCJ+k82WCQfSpkEFv/ShHgZOp8N1
pZV0wjepJnH1cuTm4qMztLUUc/axzM1ko07j8Ux5rObaosn+vX+2FQEzadczeOuk
Xn7DeTvQ2X9BmI9jf/X18pNW56I4nMf7SHMpXFlC3To9QdqX7v4OZghGxyIpLmdb
mmHDmKKnX4icC3XDze0pir8sBuDvmCXE15Mi1jiSyCy2tLZnXwjkrx4hu+QAnTsc
5YkZ4LITWj82/bguIiagrUBw1DSVaWsTT+ljulTJD94+rzRxiehHgwADWyGYvfwP
e2u/wU+LPBYJCUiKnNz6P29sOgiqD3pRcU4D8lRlrwUnMVtSyqFDEm3zz3HhYlI9
uXecHoXGGjddXmeNG0Egnw3eLWB17h9tKQDfK/x9ENQth2opBDAETzJONXLUyR/6
CQiz55aMwOtZqPGAErvsZDfgZ9BDyLBcykSY1ar0K2gPP5aGPkK5uDXO967ZV12C
h8JpkapFohZQHjJO28Ht4uegycHMc42cnj61WQQ8UA3pkaWIVs/OHFD1eLeFvkGg
n2mP3Hi0en9q5JynWxsa2qsEXAtI5veCpHadTyfI1FSaAU223XSjkbSyMqYQL3r6
ks+EbvJ8AqQT+j9SZSqyNrPk0GHg2Ct2EEFwyLfq43TR4gz2HDUlkkUbiF0uoefQ
+qVV7SPdvb1pzuomrh7+YV9M73u3c9srBvbaaDFsWNvmd/PZRSgpa+sp6n4dYgh/
2mNsiQ9pDPn5NBzMAtTEBVHwMep8s+5Q33CcPL00jxb2Si4Kh/4LeZHBtD9+kXVn
rjR1n8juZEPJZDUKsMgOg63s1Im3Kfm+SMyrXPoEettsAGRzTXgUHkyfA980bqvw
0BNGJXWir5m3WEfL0qDJPAkEaAOOL6h2GEApqawy0ntA9y6u4gm6l/+DYZidNZV1
D0d5zQ/1cOrq04Lm8+VsyLo0ob18kV0sfODk7N0nUAe4xWWVG2jbvpiH4h4s06ey
2+kBoKETm2NoGtDDSac7aH5ceSyJl4IZ/krBk74P7AbFLjUD4AkxEK+/OYgZi/7e
kmR2+/Dd5YCJDmTZMc7c5qeaTzCS20OxvWKZTulcYznkon1clncuNgZOc+o/+c2k
/owp5kjCgclRtxuyB580ca/OLbcKSyCXHIvei3tXtZhl20vJVFHPCOyB/aDgBkQh
Z+57G+8XIRGSyXK8QEDFYGaQu+2eDLMbxoQfCBz3bvU1z6djO6TEWO42oJ5P/U/q
og04DMBtyE2OKKlLRqOnmReazNHDXGw2INDGuYf3JI71jsxw+nq4cuy6FaKPTB3/
UK9jZYj0kdgmvnpn1wRIhTDBEa82+4Au7Nk1HgX3yiGVgKx/ny01g6mS3NxGdDFh
Mb/yz1uj8Cx7PTgwiRbguK9Y7qoHuaxDz+jeSufW8GDcEI8RpHntfwqSU0gTajHs
Nu+T3CWHCEiM9ruGlv1JvP363Q2dlkBBCvkpI9HqJO5J6eab3wGpg4FxWDHPz9Fb
xu9/PFGDgn75rfHUDg4OOIHSpmTBN9kwHmyfGvD8hlxGt9imfvI801rGGdcoayig
gC2LvQh6chsbDfGXgXIyNXlR2Oy/6TD2UubEWGPwqQ5tUxy9kBRtlqE+HQY5lpG4
VPbmRdAhTs0CohuCcAHoVZsu4yzcdChWXTgcb55yRFr6goRjP4UCXxqRILHCQNj/
SIhaRqWteJe2AYgw4WoeYsqHnaqPVz+uI6jzHKGDfSlxkraf8tLaWXvBudRcWJaV
gHkcZ5GJpmdBGrk4XmZ86+r4LFaw2JVE9XANRGe45WWmu791O5IPIlDXOM8xO56w
GOG+9w0ZHEPwZk0rSqfr2WIhigsvC0nQpWJQInrzaKZlenftj1P0lOQ70wbiDcMQ
MsGz2HJq7lTqjnnQxcZBQZ+EnlvfltFWefIgG0SZPnAKD9MAk6uRO+2W6cl/p2Ux
N/qhHxgaLawkgGGcpDGFOkKTlBkLKWXGoHgYBQsY+b6OPEu/k7eUswdmvgimmrKP
FNwt/Fo+pGeyv8gfpqJwSLebKPpEckPUO2IN73Yc1pJpZVwmylwHRbk+9NJXHEoN
Vdn8Nf/LNMKeLUhP8tmjQR8VL+ooEqG4GnuaB3cA/PTO4Nk8Zfe80TEjoLIz4UW8
MkHcrSpDaKGJWsxiGvn7YRSEUCoXM+0YwxrSB78LnjGlDiB6qEejApdNHX8xl7N/
72QYDwusg5lC6CI+LM5wfJqjqpJdnyYu7VqSHbDELyNWItUTP+CgP7kUseTZzyir
HFLIZ2ZRIDK1IP9IurDgtGOpvk+w1SSBqJfaAT39Ni3DPHzJerhW+kqFfaP/eUNo
MJvrm16vGjJHQ8PaKPuDDk/r+7gK8zeY9aOl8aeK1t9+/r7FszKKmEIJlelkhRI9
djLO+jpW2E2tncMr4MoBHbWlwZkDLQUgtghL6gI+5ts+Edf/EneI0VdrVF7QFCXH
apacuZeLgcR+1NtC/4bb9h3nkOLPSIpi+vrw/8PntSfivbSkcbJ5fyI1We6wZFdd
5W+roc2v6RAABivCzOdBI7Q/ujVwFGShdSPo9xpihFG9B+piyo1q139NPlENlKkr
t9NGX/6GNNEK9Msfxo0cb6Y+5g0Mr42rc11e4KvHX9uIRMVsyLCXMOj+FUmLGPt4
yhbQZ1pAJuHwLl9dvVvMfx7HDlx+IDSfzJQZXd4VAucr8XDSmHYcmUoSK4jOU83T
OBPk86yAezleKJNMLrnL+gbPqRwmXYsVkhmGLvns36Iu+1H3x6Sxe9IYbHsWPwJf
c++nJD4STRS5q1i/r1GiMFJsmTRoiBfJXs3zlhwdZuaD4z5SOjmhjHnwbsF9thTi
l82UQV2+D6IIga5fzx1aQfR1uWntQnGilPkWS/unyo2EM7KAwQO9YmUxQdCl8y4e
mHk5V36RpQnAKxlwyswOjyvuVf1QXTjYmB/K9+osB3XbEz48ujQsxkjN/XkHBrCz
7ZsZvioVZlJRlx7uL0XgN5jqTFDlaGjoRPvX9IGFeA458byEqqt5plB81PSDOxZb
gECIgJQES+mOEqQBQh2WOjmLDqSUXsFluThMWEMhG7mbOsx5yWQWF+9rNFphX1rh
VyZblsN9ga15zgN7IJkv2e4I4O1k0ujkgGz5/SA7IEUdP1gfWERLexM5gOYEpvgl
pnhvYa0svezu9ODZyabfUu4zl0MJOIrZo47bv/VKVU7O7eedeb8NVZ30dGM6DSJ8
8IVI5+3hnv6+ZByVYRufxeqvviBMH76biR8S9clKGFR3IdmznVOakriBKXFnUeSx
JzLgjMjtN5qSmWyjYyivkIfSgVG8EjnSwCenT1QvUFxyxRrg4S/Z4Wy4TJXMjMTy
Dy891apbYEzv5sZAnFcerpRKjR6u2jR2FH+hNKqn6cTXzqy3hbASVEWH6kOdPor3
o49Mo4SfF78wmf1Riocaw1gdAvpJX+1LhRgQlhgXJbKhh9qACHm8c9Ir9/ErDT+4
0S2es3gxlJNqYE+YQVkH/QImBSAGlTaMGstZbuQW9CjBMOtZ99Pd//zactM1hugn
dX65hMgiqXvUpbWtUAWeFn8TfarUUMW3FcVINon0ECmPojtqDO6iXgJiNrggxJrs
jJTuoCRD8XqKoodergD0RUionBtNlX66aJpFM0XmpEJ3gCrJZ2Yr9WTfItPjvujc
6PhDo8v+kReQKHuc+Cyv8/mnSOrl8aSf//yVHt6SjCSJHnHG3M3/uxFRajOqqUTT
+7BuYnwL8e2AUdOD5diYXTi6qs6uvU8o8PVdAncX8WOESI7mGi6+pBooQYq/2ytt
g3dN40l8RUUV8uZTcIjTtQgN/xlhrgfTmHjXKbRFb0HGKaNAO2QvD7GxiCt6op+k
mCw7j+x6GlUV/biuVNxhoJH9p0zw+pV0xKvNl/Ou8QYF0jIncgEep0mHILTvgjqX
llccEzn5UdxWtosztAboCSkJrB+/kvhOyAiB/e/diP1MLVHYMoKihUVSAaQtaLWl
eh7rFGl5JKPvpg3f1Kr01mNG/mk9ohmMKD/YmWDfEqKzV+Hqbfsm7BWTIhR+IfsQ
6ZZxyds8Dt2sfiqedkKJ8+U8lZodWRhA74b69Wz9vG0QibrzyPzf5h+df1O42/fB
cdlQjkJW7uso59NIjolh/At+48HWY89gTxJK1rvhz/2oIfpXfl0KWBPT5KjB//C/
ExNFnckTLM39Kva/jrEWyAWDSHWChD1IMhUyhZJV4spOOmhMKv9rgvc2Audbw0yL
0tgv3HKgYgEF+Lk5VCN281EQAU+p/c9LPHKM4tRmVsC5RjqmA81ddn+YKig1xTeI
BGg9rcoYiK2gWwLVoqJLFM9mz2kST0qJR23UDJCGXhKr5zYN0SaWRubgwD+DuAPz
S4nWeSETGXjYs7w6grJcs64bbMLMSY/xNw1iOK4eIZ2DypLjFdtiOfRQNxyOM2tu
7/fl3tWiGfyfZ+8Avqg6GBtiWymOiPWeviMlxYbaJnpNZNUn/Vnrio9wCcQlAeoo
XMINvHfzgkO3CoRfvCt6DX8cmnp13MEcZZESgRJ7nCNfsDAR8fiQIGgWSNbgWZzl
CtdoBeDBjyDUtQzUbLLneLxQYjqL+o10eATj/dIqCmJBAcxaVlX67OgiD8rD39rw
ydgbhgwBlS8xwY5RYpLohpUC65ch5OqsP12gdih3+sNdoO1hVXg6W8LAVbY8v6pC
+/cOQkxzK3JX5OaJWBZwpvTurhjcOY1oJDB+uXpbfF+zYwSrEstyOiT9rCL1fv0C
d87cs8JFTsfVzg9K/q9BINHSZBddWdPgLtkCXSVUBp3G/h2hqCcQPHb8rTEmG9sZ
S1Rb4UC9z127Zk5VXavRtrkQzWz3vH15kZ8Pn/+P9GoFhi+NJZZjp5FodtqLOsek
+LirAD9equQfUiOLdSyzqH79iS6T60j5bmM8CIzgrfK5C4fSLjJGccRuoi37fdqU
pJ4+MSlFGZmGbkQMiKk8v5S8VVzrpTVgajioLgTLYP6LRvVaL9NvEp6oqDLcQZGp
CBJ5vm0g1FeA4whZMDWml3GJuhcW/GqZubNLhRNQC7W6W+YN4JNGp96qz5xVv1Zu
Ci2DlYaDtsxlu2C7/gBmCy3uoJ8Ssa/JPjL2d0TqQ2WDtlpdsumfUQ36lm5PxiDR
8vk1fROrzR4pMutTuyQyigqV8Ahx0iMx/euiz+uJrDJiIRdiNubNbt/jvbIlHhjH
KyvRHEGWgliV8e8EDV7luoAzrkWW47TAhLMs+Rr/WCl1PWpS1xhgLenoocgPBwjD
IrHJNsEnO5i7ET7VPxQu1VN+GIDvItymjLDsBMGL9vWJWZcPL1Ge1mAjbMA997hB
lIg95C9KW21dIvBHVD47kbhwUO8yKhDrHHHKKpsmM4KMle1nOg0un2TgbG1DC+Yt
eVrEMhPreM11bmWzxP0gMkGsJBreHlbnDRF2wt7VfC56xFzygBRlaNhVye9/kI5F
JuQtABTsxAI02i+BbnCbEWiQ64vMp0O27ifsokPGv/ambiAmhaqDcGCMXbRG/edi
WUL+nluRruIpEuK2ay7ONJsHr37mXRIk6NC4UNHtjzLduJ/mEKypcPgjNzPlNB1P
+1xb0MCpDsvfT8bq/wzGjl54wbUFp3QzYlG9RfrlOk0B3Xnyz8noDSa4cqy0g3VJ
nxwMiD7Ml6tDltcBxCGESlmWHn/dzbLL0B6cb+I2ArhTkA0/nicyYvyMdJLw/QFJ
YJtx0cHKPNtZn44qX8Ei7hk5BD5LxklPI589hNQZb6YUzq3CSNZKUSkptK8eMhF+
BqKF0zVN3M4L5pse6HgrFZQWykcA7+zGUkSg8zu/Mq66fMqMnsVJ1k3bEeOcKOnx
ZK+H20BV8kroBIKcsVWwFsvfxt86I5gjDfsCKiFR4G+HIJTc/32pruMpnCONcTAz
nJJOB0wTnP23ZTqgCe6EKZc5VEnHhou0MpEeVTSc9zYgYtbJeX4erFbtopK6Jhka
74p3okz7lxUC2qu7uUpOLnskfhFpVP0PWHJ2ENm6nOOBupxNHGBT2ryoox9Ilpzw
gxk6tl9oiZtZ67hp2M1Ki2stZx2kSJ7J9o5M83qtuXIvBRQ7lOpHovQph2/aS+Y+
PPPmz4F8RSaxhqWtej+zAYYCRxcpXmE8RaxydaszTHZRAToao0lBi4zUl/4PkFP1
voE3Vn20gvc/Ii+kNcS8RO9W97KUEOvjsk0onlvr1eWzxlD4WjsQ9PLfxQWpmCXu
gSkA2/K+T15xhZsGnRWuh0bvc3/tB8rkcEP/dL20delbIhJadmlHIXMQ1Rpjjz/s
iIaM29KuzODKOzNAtngpEDTa9TcixT11f/TkENBTz5vA7bHHTySbl1szz94DKwob
Nm+0YjO1pmBRo017DX1OvIUgXcknBSrzfRB4tx48A/8im3SdVMfkpMDKDxbX7oQA
poRWbhpK5mD419JgCwootdy3VHwxzQMy+3m+o6xtNPH1RRLtw7uo6l83/uI+5RD/
lPf+uU53KX41b+T8OUJmk44P4iSCSmYTq/qRv9WgHjN3+ekxCbVeHeAgw7C3A8Hw
w+3cjA1UjzinU+JLqsCxjOFsIvWO0xox96xl+pH3CQwgaKvwbUGM4lnXbkRwsWpL
jg1ouVbsV6tpfIzH5DWRgsdjSUAUMwy5RRH3Vj16swAS+zxyOH/DPqpq/tdX+y0c
C1g+8EqKHc2KC8RSIRqclnl+vzZyjRvz+bnEZmUJWj0nzwOOdHHPA/rU6EY0C8Fu
asCkWsecrTc9+irtjd7+xiHuam7z+LXerJR5/hHcRDdtkmFg9OVkRJZUm6NQ2rNQ
6PxLvHHlLIhtJej8JYqTnnw4ybSIurz79vkVdeF37HHnDjDnkySTLQOTFwlpQ+ME
F9IU4STIxRhEWTDFw+LZehulnppt5Tb+ZG3z8+cOshv6kh7CWoOfPw++qXtbq0Xe
D0ZWQmfoIuN7XHtA+8sI5aVeqqEkeT7zlholOEK1P1Iwjqx53TvghfIczcGQ4Bn7
7itozWwC/gPkeIVbUa9yo+amuiceR6lTTmtAr8ZDLMqxn6c6KvZKICJr7p5oqub0
3zzedEYVvZLuBkOoDqkckodvpuJHRekq0HC/5aytjdwut7VEIXSVPBo0wmj2X08M
FxS6FKNIczW0/j6uIfvKUvDLQVBMd2Vwk6AreCjP412fGlwlHPhZ0NfHzbTsrE4v
VsGZOiKUHSv0wem/zsBDksDfA3l+weIhID7EOlHFJmTgJYJ5Cnsi29kPvsuLtR29
NWO95uPDGp1MMZZqAxUIYgjQ89G95z7rVK99K4jXyE7BsM13ZmeXRdidPlL0KmLE
gHVzJM/1WgCPHLk8mUihi9mnMP5GS7erRpz0ogojPdfHhn/W2XV04I1v6GYevvjK
Sgc+wUKtAE7JJ++R4svVOHGjVpqFnAsebPEtDsmEtV5gi9BwMhjFkdiWN6Ol6MsG
F2NzO6Ng8TwahfthS35gCpGx6xcpmZC0VgIH/pXlDMrS/Ptv1U3nMIKwwvUXEzpr
qik/evy/42Vk7YBhqd2oSn9dq0MsqPicbPgMz6ufdxu+xZ9P7mfX/YHtcyE1dQ7h
5Apamf0P9OvmKJsczW+XV/AD1mvzce3lqUZ1mNqgy62JYHsw6yu50DP9bwDtHR3B
7d4ktAxBgbKSK7lOQP0ynJZC5GY6n+LsQHPygp9cgO71WmtY4KLfkZTqZFQVCbWO
3H4t3KG8cLmsoPQ7TwnhtRgxJ/MKRi6gC77INS3vK+i/BSakZe2shAtHoqzvLkmw
FOvrqvtu1KooTCyv3ojobgywDCOJjQsdnOLct50LV6GGyLkynC1RXvbGhhxqVOY1
BHMizOqR/zorlQsJj2aKc81Xkd4+fPCJ8GewzDX9PjU88bddfQN4QVn0Z38SiDmf
sl+0ycX2Zu7Pt9J1BP2S2Z6qAd/VTV+jEvqvQa+wKsJOvooQdDgF1comDCJNKHEC
noFandKqj4+FG6b9C6ynCmrl6rC8O8POSNoAjvYLEhjAI2PC4Ty36ENYcHE/JdrY
6ZrIitB5xUw9iHBD0Eu6nWwUvzFGLA9oqYq/iIuNV7o2Kftgt4KOuA0hfnz27can
dda7aHO6kHRtW5LJ3pMlHkM4k4xFShRPGOoto2GuGROi40DKQN/eJWVJAF1jLGoJ
RIAdlc7AKmjBw0qk2o27WggV7GJPu8o1eGFCy3C5kywpZNHga5PCvNWjXWBfiIj2
HbXflE5yxR8s3JVVHDrqefkoNfCEq3phSul8M2akIE1jmbQhbcbnGcL/SCy3i9h1
zclrXo8d2xJU6nQBCsZklcOeS0za1NQN0aXhu7fNs7d61XvOuWMxB3RCXSePa9JJ
1oV32EPCUulkhruvHnQzTdeKVPKMWCZyfAEN4F+pJxpcR3feiVgoG7DqYkS74ABz
cPowVozpP0vLiklSz6xl2pCoOwZImy2lGfokzWAhDBuRJ6WR/AeRGrh2jd73JFA/
Mc2KkANZzYC76xWTw6OwanQ4iQ/t6/HpVHXseAIlkxzOubsU64hOcZTGO/XUIhrj
JfZ57LKeK8LDn1TJNlituT3OAMOScFUtBkU4raQt3d6kveoL0ptbn89C7EZMBaVG
DaFo3cQS43Ykp97znMOIkmmiBT5BA+S77jWqPOtDFFkKPvQMB5laNa5tQsahtAG4
1LtnHzz8C7zK2amYceBwnI6cwv0J6hsrdaEvAtWtxcat/0PxFw8TIa6m8C67TaNv
bvJKUvDyPnWtvqa8fSUiYqCpa/5koixrMxvUkeskxtncH2Fqh5oBoKaSkDf3RAR2
e62kGP9LY6TO03qtAuIO54KVEdvevHRCtF5cb5gf70lsnSMSBRB8N3zQbGBv3kJ1
JSEoiQ+6mtNEGY/sU7XbqVaLwRHDfcqugbILLnLITOsHhphorDxmAvCGPX0ANOs8
cXpybLBAa/mSoS8UtYU7bCqtXY0WJh479Kxc0qPHJN2KQTtlajwwrg9IF8DUkC9t
6FigYXAf/HiKHJZbZHxpQRnCAsk+0K3QA6rs406yp6uCf/UJzaiATcXNv+eMlh85
x0lEoZ5/dF1/pXKfFJbl9aG/tQnmjpazxLTwU9We1ZPVRuhkdPwE1H7GL+pP7j3f
QEHckzrnwWCm/PB0dxV3rnWSMxRlmkqhw1fD3WY2n570CayBe2omy3Qiq0U9vHA5
ylvuntnvMvu2gOCtkJbZ8fs2zQZzDsviF7gEUo5lNi1a56zsOc0ykYs1BhXw+a7I
XIobFcG7c2zHM+tLwYuelRJ5LM4Kmom/p0zk0UOThGcFJDCaOm/mH1JFX/Vu3Roq
CuykcHqK4VWVGqongd45VZlmjpvz6FiM2zln9g/tSGfm/acluLuwTmjmZwgXdAso
kC6ERf7Zn3KSdgSF65wjoS+EeUsHqWzoNBHn1i8yEEHGsuljBMBlJinbGHEtfSje
`protect END_PROTECTED
