`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rped5yplxinTkhXhzh2sWqggg90TgmKXZl0+qtQc4fhIFkZOHwIU3G+6/WUXGFka
XOy98OPEI/eF5LpuR66HO3PEuVIu8muJmJarnhD5EJL0UH3m6nA8jYSaUShCJuI1
AMA8xbOiv9QYK18o5GrVOz9pvhsQvN9UL2/rCbqeYm+XAyTvQ4aVp0XbDwTQCMmJ
wLqyShN7SvFFUXvOPW/FOAgjs56p53N0tLAHlegtFg6bwvD+xZx7EP4/h85/s+dr
X1+gyrnjSvicgGz2g2EOYtq89BRXHVrWiu8ifoxma5TBBHJKy+7jR3hVxZwfTwFB
gxX8y6wOkfC7sMbtsT185Vif+22PwmnLxGAqEj/m7R25w9qQm9gG2sFxfxPfLi4I
VvojIHYJgMTmTj2OuTh7/CjFDzzFwx+hqQX/CYpCAaeWMC43W6vmPWkAWxtJTnLJ
QEEMykDap8SMygkZMb04tw==
`protect END_PROTECTED
