`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RODJwtRIWjMP7MzQt6JcSvm0CR/GukCvTAH6cEwPvEF+tSJ3g+RzEw55eUMMkA26
n+tXDCXKIQROxi1BVeuufdeK+QLxz3mbRBrSk6gkqPGE9qfkH5CjyLN+fJt2As4F
q/ew/NxvTmZ4yyi7vuywhItHYCFGonAPbeHMw43gg58PwSE7CRjAgU+9owRELO6t
gkSXuc2h9RfousWc/BLiNQ2bJx8b08yxsnvW2Q3+TM/sCoF1hM6MG7tUmu67jJPo
lkXAqHcVF3a2G+5GUwzMGCVLpkcZ3LN4bKRuMY/sxO3VgYSYcxM9z0W3+bNbOdWf
c9iTMXSJRtZkr4EtJ6/G2UrY0hCjLmDVVUnUvGi81M9QkWzBxu30xMDABWiFV3IB
urNxayjhh0iebqlmPpwhiClMtDLxRbQwcN7Js+suXULVLi7k2gs6WVAIS3/L9mTi
APk75PDX+/Tm/QZrT7kG1I+N0BxBkzJ4UyXBm0tgIpsJkELMhjxP6xGLBU8leGdr
`protect END_PROTECTED
