`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wN/XS8Za2kClthmS9c6ZfSPrbMDn+/lOxVO1Ui+bn83rAV6XsHJu+OfMDiFiO3h
Li+QFhDEf5B2rl2TcmIQBbSGf5jIPhhjr7RKte2oY19hEhkShKCRltK9S/S3k6tQ
xLsIQTImrh3CSriV2cWEKC7qh3XgJSorQ/tabOpbXLR2HqhLiUvSi9JZJ8oE4n6Y
+VDdmxOUKNYNEC30eRXocCZGc4RjCKlxTbsMYzbzHkbHKUW+HO11uC6bmCJBWzLw
/CE1rRoL2dwNprShBvxCzx2J54/47Q9ZAEqV+UrUmOI1kkaBeXMzECnKzG8pkNvJ
x7dzwJVn/CJ1ZWv7ZlpMH+8ff4wFXbDgbL7x4ujWi7euo5Fd2brSJSvuZKe2IvcZ
qjxecmxADAk0be+Mk1SUOACg0IQSUEjwaHxWqkZRkcPdfKRnPmUO+aTsTGX45C+o
xerCWBl1YX6vF+YdyEqC6jcbjYXQB3qhwlzC68T9ZJ2jdBmNVdKXg0WJV7QfKbDs
2tJbZVy7i4W03NUvveiAmLrTDtz8nH81YvmNT7GqsA4+1ppKWVJZkacmLb8R9Hit
`protect END_PROTECTED
