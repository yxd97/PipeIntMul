`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Soaf0AuL8WPAZJiaA82Z9C8RN+NIFyJNJYyEMwBx8XuPPNA6Uswsjc7uRSLAGjyI
7AyacdBtqWxQ84niZKfp2WV2g4n6ZTSj/Qgdb23oTo6OtAYnB/fyJpx+lChdr0lQ
mduoAOA8PJdOZEyO7uLS5lt24AMNXJOtDvyrfM0Niq3NwJpH5WHAYQ6HRd5A4klp
ueXc3shqFAuRmsDutmgLXlmQ/6VbWTrH7duJTovVpsiS/7qzDJhepWTWNsN3WSxk
Numo9+kA73u1dZnhv2DiII0kTitGjbWdHTW6lyN8mfvgZ1W57S/7NCEz1V+ON44y
pLkDvzV0/Jsb/5BnUzCltGr8z1vI//MYTuCjHKWp5+47qp/6SpiY7J7MWaaGpg+P
64QzBcwcijkCUDMyRTns3+TJDo+9WvOuZ6oh8wPJ1sz1IP9zubllOOsxE51YMYZD
QGb4FYmQIZhL5mmC0aUfXQ==
`protect END_PROTECTED
