`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zKHUKO3RLQQfkCnFwX1hOzkIs6FHzouG3O2ErNe4Nj8+F0RRKUe+3l4/vLY7Ucb
K6lVhwmF73iRI9emHYmTAbQq9xhH4CnB+Ip1nTiF9gd6IhgcD0ZbPcmwjmmA0cdd
cfkKMuESvzLMaRM5zsWqXS4GwrNobhkPat9KgXkTKCAxcg1fwl3ylVrw5/h/+9+k
eaAWOiZKQF6GIhyYB9mrd+8+6yV4CG3QsQ5MjXWOXK19GAGrYIfLogrwFb4G2Z2n
O4AUbLWSs23baOslGuRau6EV7jEmfF8qzez8vPuGJFp/Cqz8IIumm9Y8jx1X8Z7q
o0GRRiWUlO447jU0IRhJ/8FyOWdycRJkgYAQPGrHzenTbxOyZlp4xIhzyRqX/mSK
BmhfAlKgR0mq1+h+uQW5brqp5LdHrI/+zZUUtT4YgeATwFk+yI279dYS1DHiLoTw
Wu4gpImRkuz317gks5i1aeLNnp5pfyR4KF/270SQx8+bkrTacK8wcPi1HNL4xrPS
MfvVbw29AkRqFB+5eRaKcRJUYNg0+nJQLHfkG9JU1etA94yRHJhX3DRpxiSMUgi9
+kAWYwCTjwYAp2SXXBV0M7AbuoVOYkaldL/h21uac6Vqhjr5jadt+f7y7QvGnKMp
Yi393LfSyNGYVYidEtc1qKKdVAmFki+1wlKF0VuUQWMjkyJa0WbA/SdY+XSI75b/
kH+ehC/aWDceu8ISzSiO0Gt33AWFov3GFBAhxgC1Ednjp6bWXYYUZLtqoh+gfgCy
shKEQvD5QilJy3a+HcosaZrpclIi/allGSd09GcCta669fsWUCzRtvJZeigP5evh
1BckIyJOWkelBxZGbpXe1rw6Ri7AyfE4uAOxxEegVYG2OkDET3bV9SCdrEcETe9y
ybsTZ22UmjEnda41vlRzLg2IeG6TlOy4APjbP5FgPySvpI/jNt6B3rn1f+bWYM+K
TKe5e4bvMxWsfjY/qVI/XiHwlDbFnwgzjwzCjfuJqU3xBTAzZWGFRuBv0I7y+Y2u
6QLOFluUMoya0anWXTBNnqzopd4fk/nGipLGOd3I0DgFTmplLsbr/se8LKPPmTkL
uqWWCgTayP8TGqIlCd/E3QIgT3mph/kpX3Vcnv/EP0ZmNoShBx0ADBElxWh1X0yB
0uPi4XXLmF+dKooi+3EnyLIqoSfLuRcDRr19dnGLTwXyxH+OMoE/wcrUVPMd11TZ
m4m1CzcV/EH8hk8y79lZQySUya8/3sidOY8ZVilVgqujPlOMA4bSvbwsIBF51XcU
5lAxWoSMoZuph08CwiyyL4ErnAcIA9G44rc0UpTPXfUsgsTR73AWSJbtuAo9gHV/
FcddBUipwkassUvd6ytu600/0hwoSz2LY/CQqF4xxTvBLTF9UjjIR54F0/lk4/4t
Obxnk1K89uQYSWgGyAOPm9hS0SDdCH0OVhgMJWvclT23LSZxAQtqFfLM1YAIs3Af
T49yhvvq1fTdNtTmqKQy3dsX1Z3utHgtAOajOQmIcUgwyVPfruso7bKMIcOUcEXx
tQWxxs71cYmXLT3IGXJlc5ay7tdGc2lAXLA9YKI/Ftf977fnGIDIzJWJLTWThHWu
CRbTnSZrQLr8rhKGb5qTwlw3ZXxRqJ+sRJ7ThbDss5cfmti3E3CJwpJonQQ1TBd5
6EelXoPA7aMYqp/Wq0Vpcq3LCKI/1dT9tZDRZVO18DyyEPFVFaesRzF71zEOkAiU
IllZBn9GHfElxZBvBWZaHbhhJG73xOk3KE8f5nBUoD+8ewTzPQj+0P47swGG5T6m
9e2YFuZBsYtk1VsaeUbGi/dBr2Iqo56R1qDJ3Wt1i8i2KhDgfdzTjhVjIjOnJ4IW
5wUmauXAj+FCKNhBSTFywlF4ve/1leqGwb32T2OoyeVqXAAgWcxX4wpWfWUBLv86
indGvBGzf8jtaqYufIj1YVj3/SUTSmLhGEyzZ/QrtfmdeHV9bSbt5XQXXRUm7eBT
oEeEBFHNOjoyRvoRIlQBsTp9C/O6Ui66VtsRt40rnX9aL2RPQd8/dcEgEq/rcUSX
+49gEeK/AT73kfd2xZ6RjMPcr+nIpQnFj9M7iqXHRfF5IoBtOin6IqH5kyCh+bGc
GTBMdvzPpYGmz3kl3tU+YmfVj1vdZvqiYGSraqg2Cd3pZXUgA3+mu1I20e535Q3I
AL2qomKe2qJJjL/Ev1TODKSNrZit2xXjj2SM88723bGMgXg68n85128k9JiOSa52
RWqTp2trncgFcvlqDhVNAM8IA2sUVXP1ikCBm2s0Za4d9OdRfv7JJx6Ukeq2DNhs
dOhkGNUX9PkoBJSPzhsFKq8HfdmtVZAEQ2ralM3AzukW5hOYrFLQ4jlCWIXwzxhj
AJ6+LTLT6aGp+8zZPlg6t87tqUJ6X9jSbJ5B1E6hlldYDvE4dsOhiy144cFBvlCk
g6mZ52l0Ovz7uVWwq+WY8Uve1YBGm/VV9MDyRlqTvvEIVPoNJZSxJl//p0GrckE0
PWVuY/8MG0HKHzs7YbkhcJ6kkpQLyKk4X5T0EcQn4pxwnOkh6tIWrZuLGQQbr6NC
xx72/lf1hS3sPx0MLpGWPU46/cnyeMbkopOroNxmqoEHWzQZCklAE2eLXjlvaGSt
oExPUS/i1Sn30S1FF8n0Z5Iu+45+i3wJ81fvbyfgPgua6UaQv/UNRzf6SFYp3mnx
03BBRM3ZcpF2VioT6iN3NmY37mp+k9AIIR3Eft6OUrcUsEU8ZcmemSgbJFnRik7m
HU9RXMS0HSKqcj8pgrOiB5VXMvgehl+8JPuglxI90/WydX82MM/rXAa92Gw3qi2Q
xADh1ySwRoVba712nvN2VeM6yC4OznqFEkoPaDTPyrvtyTLubPAwc5r+Fx1DQa6b
kvgrfZOx4t2BlraYFfEN05PcpJa6BzfmfM4xheVvzM2GR23YgY9eyb/Wg28p/PfA
f2g860rOQZJYV0O3QHaska5Zz7najreA4yYGCHmMgm3ldwC9l6CnROII20Ol+53w
pUafO0shecrBqko3SEI36j2NE5ABzHIoKNVdN21r6aToTxRd354wrCJrNbzleafD
dc7Q81ceyAibXY7R2wPiOC4TOAerg2aCU7Nb8+LYBXIgz+q37/8ut1e7sVhfo85f
XACCMwvX4ASTXxJ8yp0lgEYfjhHSmgWBJeCzd/nBYWb+LXKdwNUMxKjf5udyu5Q0
rM1lsJd5yOwMmRseOlD185TX3tOBpgp3kq2oVT/m44HsyDZM5ZGLM83UnlJaxFc3
KcBvx8543ag2NBjXhYh9o6qW+otsnuJ5VuXp0MDvwRfT2e5gd09u0Rtn/pvI6DDS
utdcq+/tRTX0uS5hpQ6W1nmJ0q7Fn7Q7MAllBvGTzYCsO9MGGLxV2NOKmeKGFzMI
mAgIdLo1By6IGjA2BuNwZuv3/79C9AlT9yfHCQ7l+he4KbIYuOT7NaJ1OrxNj+l8
brXK6Mmx7GQu911z8C3d5X14+aAg3GJ2t23yiohW2N0vA/ihKqxCJEoH6b3BP0a3
tKsG3Uw5gXy93Im81O2wN70Ca+1rgGQ/xxTUG/KBXP+m63uGRbv3SoLrq36Qu4FV
YSYgpekfzmnmra3Km24O7axrWb5eYpBmhC6Toy1wrvegjPFcAwzXqLQxZn9oYjeq
fxrMrKvpKZbQuWLjKdq0Q552LIQQeto++MHxnS4PgCiLdwWq41XsxNgdkwzVKhAv
dZoDLksJraxhDlYlkokA2XARt0/c7G7ewyTGfonJKFmI4jH/3ODQBJ09+WA8Aqel
xWWcy5QLQVcvyZGOn3mmqwbRsKVDHfc7XzSm8LSQhrGXVPTRVtuzPIgOqWG5W3az
q+52+bniF5skeDAJeWRMg7gJphWxlJ7F/fq0HZOcxi/LUwNkwtdtF3tJ/HyEzJej
FFTOS+iPAYnMHWrVENqmhxgUGYOmHmCITWM1ym9Hp09rzb83KkWOYz4DaPNONwFi
s308U0OGntbl39h/LjrF+czSBCMgwuwvwnliqUjGxSZyOa2Wmz7MxcYXC/+CQszK
vEpJGWRocZ5//WvOVOed3TLfLC1XvAZJGnL6Vx4mknTLcc6/53PPJn7up5JegEzw
h4jny6PXzOx3NUXB308Zy4QD3sD6p/gCoOTNdpbbwWj7bj9t19mOH6BWjMGKKWXN
8+oxV6pnSxpkzXSDJM1IorxQADORJvDpIm79LdHYEFJru0LGdQKH5vxetI5oDlhr
BIO3XDlyoq/U/SPS/NF1+H5vuCVYVz4gUGjeXSffe0WPsCC/r4rvMFoFiiawOlXX
uabBZpjL4I3gqUGsYNkI+vDDjgxwmvnrdZmumyERJ0CC+hUxwkV5gQEu7cNT+VQN
cw2LALN0v7l6QN1mu+KezqdNwFwmGbZ/cWK2rvVGykPQ2FXJijA6wEcPPFhMBCpL
CWltuoBB3Cq+z1imS5upZ4Q3HYUpubVhC8aPIXWdLgAN/eVTzGrqxUeAZRQ9iNha
oraKa4NqbLGxX0JhiSyfUgEzlHBmehSjkysukufOYdreg3+zEFVNKMEtHEBNyXRz
B+856GPudPs1of9VafopjeIqm/WM3mH0tHtZ/vQq7KTG2zqxewzMQjE2mm/eQUfs
tDXRk2kT1I4fTZrofPWcPEQKMoZ+jyOKszcex0UAl0Jqdleh74bnXURrsOGQQyh7
XfXEeyLPatxXTw773LY0mIEh6xmepccG4uT5X7w3gQjw/nrk4TKXAeI5ZBbihCLG
25X/tgw7udow/WYR+lqwTCAKKaWsgh347TMCnJ/zvBv8NFdiL1bF34JsjwFs3s37
ldlON/hpBnDmcWYO+6FkNLCPPMIXVCPucfcJ4jq8M0dOM6gapdN3HEo/qweOmYtY
bpsZIwEQjBXjxmtWBbWR7gtU69hkCZMlpK4BJj4WVdOZRL7NPp018rQR6RGBzTCR
e4lVb5IMOqwtpsTMF2towzoHZ4om+/30VZi/BRnGLsdIxY/o7tzTC/0vIwbQ5hF8
frgLDQszX/Thl9/hicelLngzWFkoIUvl1nmwGRKWRHE87+b4wojpg6+P9aGjFZNr
l5eREWkJgZUlivWQuhpFexIHfC+ceMgnx18mdQscINSUkx0fbv4hlXsIJ3jW52bD
rNCxvKC7yUXYEcN+2HxevJqVQnSE43T5rDhOV/ZorZEW+loZEFGZVVgg0RRIzKDO
lguGway8wxB/tpxwev/UttNjV8f8HvX7unWnrKiOeUfL75rSE2dGpkoeOpTCAdgY
EmbU4dw7r9wX8K38nYAnbWeKZRK0ZSSqh+clKM6tluDPrY99mpcCtgM3aq3A3l3S
XynAqIS9dxLjVuzmegpyawSrY+GTGuTpooQ1TGrDi9vSxrnhuQew/Mcp7Z7IrpAF
ptcpb8++7FecK1nkX9beWSWH53ybztq0rqf/o5xsoY3VJ96yAHsHQlGOxU4eCaD+
aEwxinHSdNBCvXgmTUTR0Zuyrt0kgxk/GavjacVHFnGOzz/QUGTDQmC99GrOYZs0
S/1287v25x2xYph2XdfvyirF5bgteAPb016zf1QY20dTd9xtK0t11czaChUmen23
DtvA7yoALIhteXFO72DljuyvEjw9aP8uk9hze2SJ7N5Sf4251gu9STt8rLjjPxs6
rE4CHlksMt/NxC7TU+C7/K05RaWTr9wHasU6g8WSuV5MS6/SdFx1msBEinrn9vJ2
lt4m6nQNoNKNM9PmoSlWhfUOc+5t6KsIdI+TQ4fJkC27FHTF6dKln5gf9KQzvQP5
tAJtqNIZXE6mOKVcWvnq9vEafI1TGO3XypRNtARAMB5BPu63GoBRxmhSrv3Mctum
Ruy145GqPgrja/Xdf+w9aqJ6R9arn2zNCgM9Qon8yQ8a3fTWS/zg6K24lQhX8bbW
oY1Sb2VpsqF0ctOlW34xBWRSoeRXfrF+MZbb6g1t/gm+f8vT5Jug90Fi0lAp8YDt
OH7lzHdPpYzh4gVscc+zm+ihg3YIDMKcNOvJnMAWRFizOadtJS+nvW6HLC9zk9/H
RU/IzQDdfcoeS/TZA7+MtXM93eXzb7OwZZoVqmnzsMQQhnGN5Q3F89iXkptrfnhu
p7qWSi9KuX1b7LLHFuCiZA==
`protect END_PROTECTED
