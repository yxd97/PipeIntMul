`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g+vt9sedTIkk9S0jMmq/UM/WzSzecZ/b4VvL/uYIRG9evxmh+iKc0Rph5+CIZVRZ
KIRCoPbr0AKkkZ0HLFcceE3ZYRXsK4X8VUjNEF6QAZYeDKH9y/zIN8mmjcQFH5ep
QM5JnuIRM494EHOoru2NsaDoB7bbhErbzAuqloEwBx8zsW83gjsFVx7gzNYHFsig
dnk2OgFA+eYyvgnvMbm+aEh8eG65+pT01LqROsAvQTitgwAIdF4zcQ6jilWz66WM
FonvvUzNJdR9Uh2Z7kUYOhF9aAVfqH9RLlKBUNbA7HI=
`protect END_PROTECTED
