`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y7BC5SxzF41XmetY4gusr2DKttqyk/pvOfACDfffUUEzTFIrlQzC4wp6F6MsCvN7
J6dXbBavpV0Hr7inV8HnVOhrgqSVSMNpdNVvXi6T2Hhv0y7pMQTAyvcAVp1SKoVX
YYmwjAauRuTGzJqGZaX/uBnNqjlcmZEQ3e7DJ6IVYIG0x05P6x8FGQulDdfsS7jB
NZevMGGFVel78h+jgIZpDB68j59z9YUU9jnD58t9wdsjlIMSkLgIsARFgWpmw7TR
30AwQnv7IlgGtXgr8uHf4BP4J/AbKGU1mxxmRKHEFG9D+dXXzJnfHRKEfTEbnqfw
kuQ4TZq505Obhd5vilS9E7w9lej3xztVJStPi2GOabPLLaGInPNV3hSZZkGPIWt0
O8rFoax7JiGWL7Hvk8l1daJQfzOGJGxgPO35K7mH1189HxE/6C1ie5KNUsLsoyVX
Gha9Gzz/xqXkSSIMC6qSs/utUNJ2r4z6yfQU1VT/f4IQj5m3S9WZKfm1bBYlaHh1
pnW1t7z+xuReOwK7R7KJOoJme+7tSa14z4qbMyjS+evUcCPi/s2wN7QiXcmjqQRD
lndjhYuq1k+KaepgMN9LjAyODTIjmg651xLEZhCcA7npOQwWJGu0me84lsy8n76Q
GQECq+5xqIetsvlO+CJeT2SbgmScHb7j24/+3K1YW3eHAssokTfX6kEp19p3iX62
FDVxMwL2Ln1uSjifUTGBOk1SPD6s4qJrkD9x+bAhuBJCqCcD/QiLCdYXLfotJQ5c
Aa5c0JM6fatGWflUPNE3vn0yBHyjszMXzmiAhXUQnX0Y9/6s13+ligGus+qC/vmu
xg5JIQVSofJGdgqCV4X0O4293FzDGI4HKj7CoIvQjhwomv87udfdwZpjuK3jwois
xJ1I3GH1rqIPuWVVBP+jcJQtaB2A4RhBnHvHOEbaVurwjB2VLhb+ZRNVPyEAsv8u
O+cRf6LtpZmXj5OJ2RzQhpC6v6VRUkpfu6YD1wwcVpLVq1vQMMGGDGLcr9e5G3Aq
23x9mFK6Z3sJ+BWc4+l/762OuDyJ6ctT3bblnrbOnHEIC3b50vO6QhwId1f71PMQ
svx4x451DGfW/YHStwE7jqiglaAuqjjIVqhe3LUpLkGkQSBtqiH4GiRo5d9tPMFJ
9cCbaeaa7t078U5N+ikXyLAtNZtzh8miJFdTN24eChjBdeMMl4EnPQ5wka/5b2Vj
nyxWf3XyBYR6RCq8JFPT3gj3cbqeqHqyuOr7x8aeU8C6o5Xz75cUKn+tT1QRbRWI
rxSwUjXVs8vU8tBxnSP+8QpmJKbualsFpAGOAATJhHEXnA2IOf/2PY4t67WVH2Je
ZpqDHkeZYrfIMkHR/L2C/Lk2bN8Tz4dvDKhxtLCQ/NlrRYHENOKHkyB/tM5BmVi5
yL1jONnIxZZExwkHxvRf99h9+Tsix4gEtU4KWHmXavXs5sqgOonGdH2hyFtuVlOr
XvaHeffUUnRl7Jk941VmIJlE0HBrjbuYC5qRDg1dni8IgYp97ru69TIxLvTGBfeT
08MJN403/v87d5UkrPt7ZaUqH2E2s8ADO+L/4lccZLA6gm2ahSRPJmikWf29p6VV
iYixiXnh7Lm3TPH6TqISVbnFvKSKtB8YBFfNtiKV2fwxZ0sX3Mm9aTMM9+UAutgv
P1p44uizAL45cQmIHsI+gbYL6J7Bzcp5kAqlW0hQlR+1s1GQn8ylC/yLaGTX6D/j
8PGQKGw4VzVJY4uYKMpYbi1+ntACsbinkuHnkPA/3wRN0Sa8XyvS7JSqHtPwutFN
rIuhhQjlodhWQuWQIXh2FqLUnp9s9/bqoH7iV+Leq3vDSAJvCZ5PNeqcDnM/MJAv
KO+liEf3t771Y3h9arK9Iq4pTeVghC0rb6BrH2Q23WD3bJH93gtpPPSqnE0wv+BW
k24daFDRESmTSJGW3fmNryXES/7uLLaAvDBosGczUv1no2SkuJSdsyLpF5AS5biT
GXqUPs1MjLgL2v+nVQEHhGOETzXjmf6eMtGjcRb3pIFa2PDgTiyzVER0P0lVDvMS
EbCkTADckG4IY7RV+MWMPrlS/x5apBjfrRRVjUCUOerVV9oJ6bvPhssuX+9Yj/CO
az4SGnJzR/77Y3WDo7tQ4zPLTcD+p13XJRYGEDV6xPxsA1qbPno4o3WlAQwntq3r
kJxz7tfABh8X0m3E2LXbxgh4x+ldkMc/5g/0C1kv6pAbY93WFGRcG2Mmuj7jsphn
QbIptnJydmkPDR5amM42DFx4iby4PLbuqhemUhvrLy5NNoxqDKt9anSxvsL4YWO8
1OHTpkvTagAUDcQ0gJzu/gQopVcxzweS5Orr8vjU9wC317NCeUy2miSu+PhNSBZI
jrM3w1NZtmj5IpQ72OXqhgND5qGWEvO/MS7qxaiFAhYl6+sGrf0MU2+bZql/OUep
NULzO0BmnrpjwmilHikTPKMUzHetQTePbrPcIxGghVQZcZKV7xMjfD2IRWXiH5ji
Mu6N6ayq8xVAcUOAFa6pYAPZ35JlyT3W9ayQiE3nTyVtrweNbvidjVD6oY44ymmR
uNVa7glRdfygIcnoqQAZrrPpT39JYDmVt0WBEYIKhRfLb+sS5lHwYmZtOo+ysVT3
uj865AkzgxKdyQ2fpe7YueHGRs0Gk3av+gaAKhlwl6pwOpgikPtijua9tczlxAcv
F5pwhyUIHCeXYP21ysoIbs81YWI8aXrGTZJUyyejfhkPDnXgvjkWrg+HGw6K9g6Y
PcqwbIQmEL57DuwaaDOICYHpvotWsG01MKqHhMGyiTMHukn5mQ3mYuwJr+SYU41A
B5knmqRKX2nIiQezGSFYskFLgCBMTQlnTwAHoiJQ+ca3+FuYJ24Tul8VwSdhjEOo
BTmcQ6NhM7QQIt3h48L/q1q6eWgZ/b355myBdGOR6HsStNsWTPQYZU6lxkN9iO+Z
LM4q6ONk435PRPN0+niACdI55KjAiCcAAZrCFqncrzAgmPy9t2D/gp/eqSm28h94
mY0YbD3br5TIHi5EaSUaIpo/Q6DVmvx6mF7SAlCy3Mpdsz/o9xSX5Ek+CgMdRbcm
LJwVdd6FxoQh0i3ZS4L+fN3SL2zlEOlMY11V66bnqu6uxzjoROQLJwWhEpDUAB2j
SNXVC71DeX/hZQvUWzef6ke+6J5VZupRqKYpSdqNgQ/vYZtD1uxbGskwKLCuDw8R
Nn5maJDrONXdZQaUSuiujcHywGzUm0buHPG+Y1JMv9EDq1935RLQ0VDq5r+ExYDM
d9ElxuRtFa2dPWr1EY1/AV7o0ik7fyKYre52i6vaJhp44cQHUDlVHrYwAjoD1gVc
+/GbURzot04w0Aaxs4i7IwRoYOSp2eAa7vIiW7f+6JEcR0mrz4YOgTs9JxGxpOFz
9brFTYHtc/YAHjfhitT6ZBbPsWgNeBaaFVq2FDXvvvMZZK+LJTbFfBpYm0LRc3uU
7H75dqSOVyvontmkB7jWrsvYZseUtCwEo0VoQoas2cPxLqyaNb19Z+L1EBhUHRVP
z0LAiQKC8A6tYdlTvQ+YlB6LcgmXKlznOsTygl8ZL7VCslBCuFyywUalYRL/kG9Z
5B92uNtPLs+CXhlDxzSjTam63g6+Eq80SVjVDTyRtdWzd+DYsGcOSHgtL1l88b4O
1m+ZCJFmUSxA817ZfkQPPkqlB2frH9HPyEBNscJ6WHIZgLLuStWciXpv85aShFwf
iiTNjFuyFAELOBLEfynoFHMJb4FfrOQa2u64qB85bFVrM3rT3A3/WoUfaQTi+e1m
k4DaY56H7aoUGKZeESuehP/GSULzv9JXx8EHlQbU5gE+pvXWueLT+mMmYx4pws9U
wjVN4sWo8dxoJjA040oxGEdGlP9W39a4EGXx+2V8RNoBHd7kxTHLZ9GwiQxG8iJ+
hGRDzPhfkN+Onpa0C1BRVaZVzzVXoxDi6QLvFEyvUfUDDNw7QLYhKllMKLKmnaok
NrRxt/jGgnsYwxhAZXl7O+9L8WLLEE9llh+pLOv5RzFJXAN7ZoUSDhdgvtHSncob
naOwHFecWULxgd5WxoWhqW+wKUyaaKBefHfeZ9c9RR4uAfaPCZD5BAYLHAiC5L5g
YVeENQ2Z3FMAYzSAx79ymSsNQq8aEqmZZ/TdsECvjuyh3sTcOUO2mMbAR+hRe0I6
6Wz9ZjJInI6ZI0YUvXtv+n+XKZy4aujsmPVLL+Z7YL4ouNl8ZuS/GDMNx99UP4wa
vHk7j3xhbE95pkp7HaEdc80TZ6QUHqqscvRga/EmalhVSSR1wxyUJTf51+uJSS2L
U80KCu5vzh+844FQOtArmMZPDry1eX+GBsTuvXgltPC0jJNWGfSgN8QNABV3Z6sY
JY/9yT9eSZRaPxM0aB9uZvTXfzH57BmW9ENnDAxyd+1NU6k3lDYE23HO7A7b3YuO
bFvhU3lRxBQjS+5CkKtQW6j/PXIa7R+OUGbkTCKZHK1JhSQ65hSzOQUosKk40Ei6
7dgOzVmtwEFjQFXlOXko6uR1fskp2IUL2MTA1x78Bix/Ls35mbuhHkNd6yCdqDPj
t952XgE3n8n3gVP7YInmX+mS9BVBGZ2vSvc5JJpeaXy3ErvFFoUSs4SFQ2AuJwot
L9cMe265U3NtJtsWSTEqAGVMHIDld4BUTCHpRd1X4Hk1ze/9Fn/VsqgYVXh3BO9t
Vej6ao2ytwfO/vGPnMNr4UnChk1zFks5+wM4MAHSLdLcigiKfV5Mp3wwBIbfX9mp
TN7LwiZnEkTZLBvU6i/YLIuj6dKeF9Fsq+bPiPSBWmNmlfiM7ByVDt4Cd7qWBbOR
/5wYJUcp85dKGaVvMaQ4d7PhLab1V00y3EPdIxhTxyBwhu8QJVDrbpHsdYVQDKwG
z0dMVr/E0EXbRlrdSRDw1hcA8NJsBGiOPot6s1d+gbe/05M+C9uYFIjMOt9QkvZ+
DSW0A5xsurmRgc+4liwVWr7/twxrYKGWspDNZylt+okimrLxf84cmM/qLnV/c5lN
k2ARYVSl2OMLXF2eafJbHxAJzlffltydDqbaWFPB2nFLotMTVuZHLKgGHEs+VrRI
PcYkTqHh3OTvI4QT47M2eAEpKF2C+9yDoIOsgbOdHqYDfzV7eh6hXwcm64BGqjPC
bypzXtmCqVl9QLUga+TkJO4MFNzgj1l2fo3IsISLssPToBqhf4vzSgN+Npkrm/42
9BfiDBuONatpCHmxqIvY2yKCVdjg796BlhnGgO+cHDCNT39f60DnkWwpgwI68+Lt
nobMFN+16pjGps9WrAgofdYuNjZNFG8BHP5myoG2cybQ/Ch9oReWBSv5LCC8PJEy
WzhUNYEK2EDxOgbrkAi7mbFWUasZiv9IYr83Wb0ye6vKhAn05CgKZLOEPLj13JSS
clB6MSuNyv5ncBfgzrhLazeL//5XdAC4/kOd8QtsC4/PyHfBoXENxsUp1dwEkMwG
`protect END_PROTECTED
