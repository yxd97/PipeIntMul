`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lfzzronb74lGhGhNINu+eDxyq0Lhi/1lIyf4c/Wht51y/OQ4H1ifkGrqwYgydZh/
jhQOQpr2AHS0EqdGxI4qfUqwsDXGQkhMfB0RYU1mhIDR5EUuEmmUHe0DONvxlAHr
VCgonDsa2NqjawmUdym0tpj1dv57fGguEsNvRLziUhaLfla7XbmHgZlWQb0/51Qt
uYxB+Eu778iRxUf2dGLvnCLyAAwEVNVulvZu1th8x5Rf/cqBfnk4KG8quTdUs/Dk
MO9JclmPDt0rJmSzLx6eubHsfuqa7ol7E/CVi7KeGLgkJJSOPzkfHj1ggQX+9sGB
ITa/cQU1hDBKJi9nl02Wao69EjuI2N54u0SzJo4PKDsrxPsuJ5lhmNWBh5R8jg4L
Ml5ltJoRl+mCar516XBSK8Rf368w3yGCyyuRR5EL5bpb6aAqLk9nSPc7zPT7FoFB
yV939i1xRMwhIjCh4PIg1UFlGTSLGQsxZpPFwXbkO13LD66gRV2jOArK/1zg4Q7Y
`protect END_PROTECTED
