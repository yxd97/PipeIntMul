`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tRHCGImdKlKL7vip2ftGw7++cAwQ4wOOxu6hQA3WBfPYYh6UCMOcZXSYvkp76zqH
lKrTlDHCdveKe6w0XrbnzPoHUh0cBL9FnjLFozNz2OhNUcC+m/K77ctsHaLHZzS7
2AmnyBpuvBbbH7qUGINh4mbB8TyRrsH94ojvPNnYRkxRJcMzzKALzo5BrXn1RbXw
veHrAhx5lYLTbFYJ2m+/A1nSlHCGw8IXbRHQ4eklAoIQW+YNcJEnNI16LXkEZwRH
BO3Si4FnoVzQRcgANA15uj+6jQehtAhTV/kzVTgPqg3ddpShk8inr6EYZODnHI7r
54vp4nTDZzldOEMIZ1CCDv30qVZJxYrKTkz4XPRFwg2/aA5gvZczkZfjfQGGdSTY
gD/Y4BPWx8v7CdVcA7nVE/+7n/YHZCy4z3rJJVcv+KsNhSHvom32OJh4dVJyuLsP
bySIKXd2/Tsn0kUiLVrxuR2n1WRN5w5oVv1g8e61mlp3pO6whHzWxL8X8KXLin9O
x4VVgqTSGW70eB6bduRoQJOmR+AjQ70J93gCdnWxKF9WzEHUKGuQMmOhdhNleBzx
NDfgD9BpRhV89V6UuxI5Qg==
`protect END_PROTECTED
