library verilog;
use verilog.vl_types.all;
entity X_GTHE2_COMMON is
    generic(
        LOC             : string  := "UNPLACED";
        BIAS_CFG        : vl_logic_vector(63 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        COMMON_CFG      : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        QPLL_CFG        : vl_logic_vector(26 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        QPLL_CLKOUT_CFG : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        QPLL_COARSE_FREQ_OVRD: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        QPLL_COARSE_FREQ_OVRD_EN: vl_logic_vector(0 downto 0) := (others => Hi0);
        QPLL_CP         : vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        QPLL_CP_MONITOR_EN: vl_logic_vector(0 downto 0) := (others => Hi0);
        QPLL_DMONITOR_SEL: vl_logic_vector(0 downto 0) := (others => Hi0);
        QPLL_FBDIV      : vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        QPLL_FBDIV_MONITOR_EN: vl_logic_vector(0 downto 0) := (others => Hi0);
        QPLL_FBDIV_RATIO: vl_logic_vector(0 downto 0) := (others => Hi0);
        QPLL_INIT_CFG   : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        QPLL_LOCK_CFG   : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        QPLL_LPF        : vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        QPLL_REFCLK_DIV : integer := 2;
        QPLL_RP_COMP    : vl_logic_vector(0 downto 0) := (others => Hi0);
        QPLL_VTRL_RESET : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        RCAL_CFG        : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        RSVD_ATTR0      : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RSVD_ATTR1      : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SIM_QPLLREFCLK_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        SIM_RESET_SPEEDUP: string  := "TRUE";
        SIM_VERSION     : string  := "1.1"
    );
    port(
        DRPDO           : out    vl_logic_vector(15 downto 0);
        DRPRDY          : out    vl_logic;
        PMARSVDOUT      : out    vl_logic_vector(15 downto 0);
        QPLLDMONITOR    : out    vl_logic_vector(7 downto 0);
        QPLLFBCLKLOST   : out    vl_logic;
        QPLLLOCK        : out    vl_logic;
        QPLLOUTCLK      : out    vl_logic;
        QPLLOUTREFCLK   : out    vl_logic;
        QPLLREFCLKLOST  : out    vl_logic;
        REFCLKOUTMONITOR: out    vl_logic;
        BGBYPASSB       : in     vl_logic;
        BGMONITORENB    : in     vl_logic;
        BGPDB           : in     vl_logic;
        BGRCALOVRD      : in     vl_logic_vector(4 downto 0);
        BGRCALOVRDENB   : in     vl_logic;
        DRPADDR         : in     vl_logic_vector(7 downto 0);
        DRPCLK          : in     vl_logic;
        DRPDI           : in     vl_logic_vector(15 downto 0);
        DRPEN           : in     vl_logic;
        DRPWE           : in     vl_logic;
        GTGREFCLK       : in     vl_logic;
        GTNORTHREFCLK0  : in     vl_logic;
        GTNORTHREFCLK1  : in     vl_logic;
        GTREFCLK0       : in     vl_logic;
        GTREFCLK1       : in     vl_logic;
        GTSOUTHREFCLK0  : in     vl_logic;
        GTSOUTHREFCLK1  : in     vl_logic;
        PMARSVD         : in     vl_logic_vector(7 downto 0);
        QPLLLOCKDETCLK  : in     vl_logic;
        QPLLLOCKEN      : in     vl_logic;
        QPLLOUTRESET    : in     vl_logic;
        QPLLPD          : in     vl_logic;
        QPLLREFCLKSEL   : in     vl_logic_vector(2 downto 0);
        QPLLRESET       : in     vl_logic;
        QPLLRSVD1       : in     vl_logic_vector(15 downto 0);
        QPLLRSVD2       : in     vl_logic_vector(4 downto 0);
        RCALENB         : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOC : constant is 1;
    attribute mti_svvh_generic_type of BIAS_CFG : constant is 2;
    attribute mti_svvh_generic_type of COMMON_CFG : constant is 2;
    attribute mti_svvh_generic_type of QPLL_CFG : constant is 2;
    attribute mti_svvh_generic_type of QPLL_CLKOUT_CFG : constant is 2;
    attribute mti_svvh_generic_type of QPLL_COARSE_FREQ_OVRD : constant is 2;
    attribute mti_svvh_generic_type of QPLL_COARSE_FREQ_OVRD_EN : constant is 2;
    attribute mti_svvh_generic_type of QPLL_CP : constant is 2;
    attribute mti_svvh_generic_type of QPLL_CP_MONITOR_EN : constant is 2;
    attribute mti_svvh_generic_type of QPLL_DMONITOR_SEL : constant is 2;
    attribute mti_svvh_generic_type of QPLL_FBDIV : constant is 2;
    attribute mti_svvh_generic_type of QPLL_FBDIV_MONITOR_EN : constant is 2;
    attribute mti_svvh_generic_type of QPLL_FBDIV_RATIO : constant is 2;
    attribute mti_svvh_generic_type of QPLL_INIT_CFG : constant is 2;
    attribute mti_svvh_generic_type of QPLL_LOCK_CFG : constant is 2;
    attribute mti_svvh_generic_type of QPLL_LPF : constant is 2;
    attribute mti_svvh_generic_type of QPLL_REFCLK_DIV : constant is 2;
    attribute mti_svvh_generic_type of QPLL_RP_COMP : constant is 2;
    attribute mti_svvh_generic_type of QPLL_VTRL_RESET : constant is 2;
    attribute mti_svvh_generic_type of RCAL_CFG : constant is 2;
    attribute mti_svvh_generic_type of RSVD_ATTR0 : constant is 2;
    attribute mti_svvh_generic_type of RSVD_ATTR1 : constant is 2;
    attribute mti_svvh_generic_type of SIM_QPLLREFCLK_SEL : constant is 2;
    attribute mti_svvh_generic_type of SIM_RESET_SPEEDUP : constant is 1;
    attribute mti_svvh_generic_type of SIM_VERSION : constant is 1;
end X_GTHE2_COMMON;
