`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LU9Ra3F0LmVLm75rD5JNWhmsDOQ2I9xeCQKbzk6F5nuKQmoy7yL9ZVaa2HeFlMK6
JcWUuNZsN3F8TTBFjLI9pMyAcY3vL6eR7OpVK4hByjO/9Bz1ZKMK2VDRq4/xjCO/
AXqunNHswddFT/MmVv5Pe/Rq8zLOb6nTmn/QZVRP1D0JCb5Y4yzxAo+HVFB6mMTb
WliTws1/DHVki5ZANQ6mlQ2dIg8DYCWnkN4Ic1SvPVqvkifN7KQ3F5R9A43nWoEK
WT4U+w1ueql8ve6EUp6XaRBkyo0shtUGIPsBEW22Y14=
`protect END_PROTECTED
