`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NkrzuWuVOfq+FgUfsBnyTUiAfGQfqcxM6M9mJrKM6oz7gFpNenASgfdlIKIwkm/
jFAqe+87m08KwnOGgLWSElU44N3TcpjvCNcVLHqe6tSALf9P6+3MsrC0W74MPP31
zbHSivXqpZeH0iX0L1v9MsRMnDF1tIb0A5rU5W3Sxd3cxrNwmlTXO+yLko8YPHku
xuBe/1mpkeAgERyp6OPUGimWhB+NWJDi8cJvVu5av9LI75+BJv9k4IQVLjcIxGz0
DrAybZgK7BxDqN8ySl5Zv0r2pFu7T1FDvoZPRPWkIZi6UMZBlpxEnpur/ToyMHn9
l7hgwr9mDENp/zfj/Xm9Eg==
`protect END_PROTECTED
