`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+6BxJz01uMqLcklMXQJTq++dCjmOc2fXw+4f7yGep3JI+2eMpibj2zvL3sBn3Fb
h7880esHAbOKthgLr166MguEBLBznoOpqK2+9SOgRlqfTXU3JJOxi0poFsYpR3C3
WchUlnXPVfwvIj9Rmj+LcoStIzaA7WvYdTJX6JFapGyxZCfrPH4lV6eSHkKNYRNl
DrdT24gno15qyVr5umaaq4DUtaKOhpGBE1jG0xVp27l1+bxTIINyi9fom47ADrgh
15VrGOotSg1smoJjv+EsizX59nu1/1EeG/BwWfsoFaI0VdeFiXIpbXdhPjcCVsZk
kjpLJWPa/T1YMQFN2pdpKgPDA/qkxKB19gRZ9KgiXK6kdaK9+0Gcl0c5XBcVydYq
AKbH6qHatt/gj5QvvAJV8FhrUbxv6LXf9rHwVosoUTaLwCXBXs7vf1RAfJhkEKpr
apePjFmdxOoTV5Qm/SdzbGcs80rkt49GejyMzqyrSEI=
`protect END_PROTECTED
