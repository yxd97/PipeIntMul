`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZNojWzQ0irngvgZenAQ6EtUK0BnO65CJEh4k09l3t1Gs1+1mG640/SkMNRz2Q2g
GCig/ahuZOd9xGezNMKuAzQsEK1ct31EzEhaJnMvNI+FBEtrOu7tZWsFY1Ee0/kd
eWk/fAgJB7fC2iFaUggBvBAzslqZ/sxZnrTUer2T1CK56k84LKENJb087Tw7+cAL
syGE61Hx2CnIXhlifnqBQQNhNO+UAVq6BUjXFw6lREVRRz6r8NrU5a3Mp/FTRoTh
RPsgg1PYw5amysR8e3/VUxFdHDOkN3gJcG3OpzgFVXsyJUhMfxlHPg+5it25Jxl6
F6lGZ6sNzXNtpwjdxxMGURno4vTmKD5qFvwUpuQoExmRZhaBGKFoKMdeIXc3ScRE
6IFJzgKaYWE9fyRROXtgqF3XAQball3wB2FZW15vtgm2bbceAohmsa8OGa5mA+08
WQYotcmfWFueQhnLwXf9edLhN6PxU+EMgpmnHJW21cjDALv1tPr6ZlzNNrYx+0+I
ZXTwx9Girn6zs03MCHU/aw2jU6yJMIFw7nxw2Yocvk2vO9Fs7qVL6AtIZn+tWvFM
jEfQWI2lYAaP9gdCHIvIv5BhtNvS6oisVVUNzw2/SmiYnIn5qif0FOExc628HyOq
Kli2Xdl775wDBSFHmjraY+tg526cUufZnC1hsULjj3nRVvOWFjxwi/neCljpt2Oc
GWPAeUSqDwlQcEj/D6BTeO8KtnHv+uQz9awAVSlj8jX5OIbV3/mV2F5uyZuJU6cD
lrjOjI56VQOMeo2G28JN+ssf8U86b0WfjAJUXqnIYHZrggQSGoW62QzWdlrYE8Fd
p6Ve4i7uUmOyEkscgLTkszbFJyOIQua5LEduryhVNszXnjhHFowtMUoQj9gaoqa8
gEjcIyXZvBTn2A22nBxkWjb+WSKRpOUp0qGVIcbae4Mkdv0/J4KzOLH5veXkkPzF
3WniXgNW1sEa8Ac/BjkiMW9obJs20vDMSHcKPWShxBu0xec+SxW6E8EVzXwSeuTv
iejGGZuiFncG/mGkNqFKScC0WsCN4GSbWJ3q4XqsSQttUFINSgMP1C/cfI5w0ogV
vpd/6jSy5nT364h3L1NNUPLbip7vfZ1s7acgJ1IbOKNYgY22fmBsKb9Vpnz9BT8B
ENAU0agl2fuFmof+zaByU/YpqvKtztTHVqVfNtCLcIG8UnjpepL++oWcAGC3dbw6
3qBo+Eb3ZkbSfM6iqrAd9w/8OU90JNkhnKNB359eGMfgSG8Eu0lcruG9d3gSJq9S
vl0Uj3qvNqtirAeloWl4wdFYvEZJOWyD+wxhLw3SOvfDKYhDeVxWDX2MJh6XWymK
f2IZ5oCoL5nft/b6CeJ0zeERXWxfmjs/iwK+4kkoRoMr5CE0oqhViiqY18YRV0eh
twewELXr7kq1lkFs/IcjRvnkW+AJM/wA2Cr8VBypSjSXosyxsrIuUDgBiEcEb6R0
XIdhw2Lk4L0i6KtQo41k4GnlwEHPL34wn8O9NyZZ6nZ+1a9oD1NneWmCY5Pub6Gi
gmW85Myj1MWyM+4CWamuzQS0sm0Iy5HYddHy7m/FgNp4wTWl8ZK0YF36F3tC64lu
FBOgSKHEmrKIIhCsNcFg8KYRN4cpEuQe3mz6U3Khh24/KlnvaJAnjTHBoYjTnoSq
ulIfM5UPsYaKaCXchsPHAOBv6tATiR2K3mQn7GLaDTBB7JcmKEGH0SC513IWIfbA
Rqi2Mo7rl60hNyathCVByIPQpcdIE6F7Kf8M2wg4Oisf5jn3wlcEqc9DZJBgrD9A
T21znYQ1m4vzRhYHcFWbfvO2S5SSeJH5YKHgSR8ZRZAA1r5SCuk492HlUGK2UMqC
8mC/z2dXU/pJf2Rb7QNLf1R1jdByzLUVp6D0JmPwvSWlvGTubwDKLi34tHML9pjv
V2siYGE2VfsGgFft8+YesqJQxxEM5QbWrIi1QurVs3AyeTJ5vR1ZQRa/kaIPW8Av
RNw9LLDfQupqjrZzXKcP6TxdlvQD46WMM3VYoLoJlRiohu4UaNdfBQfArHKqiPYJ
LSvZTt2VqXx468RCcMPKE8DjXUUl2e+dmbk2TE8KGVOAmZMtnkOY2/YtPMwcLimw
iFSBf7l+MhsxBWQU2RQtm39GOZ8A81np1MdiA+1Cg+uwg2k2QIY68LhJnaKvm6B/
1zxIXeruOKTyG+Ox7+wWcI7xBF3c6z7yZkNUDTKNEYgIkot7BilYWENj9iax/8lt
VQRs+CFgJCx1STPXM9e2ZwKGY0mhcqJ3vSE3c6pDKUZJ+lheF4+/aLE63XyBSXZm
aRPS0lUwba4JIBikaddJYMvgBpFEAtIOH8rknAsZscjEMpYE34a09cWMcZyIWdOy
q+TCgWrVGCtMg9hHDbq9BdyvOhbRaquEQC1mTdvEbOsOd/0JJU2DbDwxyhhwnwZn
SKnn5icq/u8KwHjHu2X9DMTt8sa81jHOW8IQaxwH/iKN+1ue0EGHHQCGI0nXpOP6
IdVz+FugLXi0f359Jo1o1sUEVTnDCGqQz0MAtoQqMavioeMqfvzeiu6uER9ZKwvN
nqBqQctyfFIm+pRPs6EttiiUkz4TQPKXQ6Mlr2Nln+igi56kEYnh9r+s7O4mDBGO
9ibIQooG2pUFFCjFAg560id2VzCOazKBGByN6jAiHUXwoamVp5PHlrMB4W0vO5Sb
lU5ygYEhANd6pbjZPYqmbzK6KnV0YI1R1VY/BjmjTIGw8lEcXsVhVz8oR5bA0fJK
X9cMWRylycRubCpqnlgj6S+uj25mFWp8rKZYIaJViaYb7zonOG3cDKk2/vaM2F16
1Jnw3HHRxulnxbgpz8pNy9gyJ46yZS0uwrcHjNdvoCZmTK9OfL4/XOMmGbtyYQmD
ntRmGW5CSJerPe17OSzL0VANP8yjJIl3y6MIhMM3B7mAVKTdIFWSzcISEPGh8+mB
5M3wuWQauL4x/nkzWfBrX3Wy1YVfzYhweWGubfROqxhLCRVHJjx5W2OBiAcX0qES
ts4OkoVNv5+ZDqBQEQ3IgefA0v4HkBIwkHCfXZNvNHpQz3QLiZ0NNPxKGWzWAi3v
V0jR7GW1NnJJS5X3aN6q3pgGw3mp0dp7G8qur3NAGXzM3M17qBP9z3xnwgEFT2+R
VZOe0GBZJfmnaMk3t3/SNmhFNCPOncl+O3riZtcgojB4CdxUxQtoYZd74UGFzsbH
UKxRCM0ClreHQ4q+j1BLr2jt4bYyK24K7sl5djmS1OVr3zkLbKR9dLa4y6m1oOk8
Sabx5HB6d3nE6QKfenYOjbvcP4gEDxlzUhFT9CBlUchh7wcD2lwVSjeX25d3G4rd
k0EyvfTuKzofmM9qli+hRChVclygoGNHSwLg+UNeVUbtk+FR/rORyx9X/BVXO4sY
Ts9wAPRbvyla6vc7vJNVTY2fC6oYxOg3KuOv2ng8vAqQB5Eif+dV49loOAQd+IVF
vOiGwNSFgW/KgdNnfyLNWrqjJsnpv0rB28WSAAKrzZQrZPETk2LQq8959yQHxLXR
2DvOlg2AspkLVzH9rrO5VnuTl+SLxrgqA/abeZzGgJfw/t8EfBYaCRMf/ixO/lG/
kS88aUMN4ntsChQYnQrm0BpN/flgN6JTSIAim0wf+T5dUv5xnoJPzhR4gQw4PVhE
7LKXYO4L9wNDqMbv9RyC6Gv23pK+LnHJbJE7pAd4fQrgSvrHWwbGmctQFyUW9EWk
X94Dlm9eN5nppCHqc07AgZhWIKfamBWYW4dg2U4NFaWU+80FW0wPqo7eJXu9vkSh
ZdFRD/wcDRIdAB/HplOy2nN4ojYWdQk1Q6DmdxGIFBDPSw040x1fWVYjL6ZTIDwq
D8toSL53k4KL99Kl+HVDLJQKMX8C5s6ON8b8saCOYE5SZ+dq7tsAdQpg1HbH4zVO
/y7/dYWCW53Tw7dLjFrIk0dMULTggmZ8+BVmBtgck8gmKGn+jTY4NP/V7Boo4MC1
`protect END_PROTECTED
