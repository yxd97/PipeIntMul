`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XQP+bvKcPAx6HLgO4Of1gJcqpCzqM95Wd/OEHoGeYWi0D+rg6axyie/TFCqlRTvw
21SVxgSJG+AcrOKycnRphOzutq7E65PFqpMJw6KS8dAghdvscqiwL5+QNO/dzlz2
uIOoaem/wnaWNGs+5KBw6bQ+xmbq1rcV4hz2Deg4J2VS+/1NFm0JXOQT0PvgW788
pHuYRLjzWVtsBP5K4DfvBgdCSgJ0oXGrLvx4i6l0TmQtjlRU+HbgW9T2X918yzaJ
4k1xw5YNXlfG4wlBkBd3t1UkSnI4I1bc43ZTRKx+gCq8I7caYRp4WmmgrNE8euFz
2T4nGCf3w4aRNYLLJMr25qY/L2BCEcHjOd7+ltBaX6Ocm1+N14fFh+XFJt/yCwoc
qEmcAon+Yjpt6fSZxFWUjW8u5KK12LWmEdGZylroiGTqHM1Yv/zMYDNfnwjlGCVg
XFqt5aShl0G8f1s+ItmbNP6nz7EqSokcY/H2XWreLR2MVmPJQW7rLL9K95pmSN7+
`protect END_PROTECTED
