`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jVGnp5gTnwbiYHLABoV5XsZ/UfW3iWjvmTOOV7Mltk5pbTY82jJ49RAHsf4EQT/R
MIHcdWpxeSo/gynloerhB+HcZSvFsKV0CCEufA0xK+16qIhhjee/RWrosvF1xUpU
/SDjRBRgpp6rzrP8SgQo64Iq2skv8nOI/b/Dkw1k6sea2AO2YrSQlbSWibPpwpw7
h3Sz/MgfLFLnzIHiWrRc6tETPaoR7lVLFGee6zHtJTUPcy2QT2fuMjTwe9cwLusQ
7MTUR0JrnGZqZ+vt30YfyjQf5gm8cTCxoAaI6WscJzI+0bpvTPYL2bFBR/Dc/oq3
EGd3gSOrvpy340g31RCoMrCmGuUwJuALnhplEWneLRv5ortr34yxeyQxgFATscxb
h7Wl/+W5LZarrhX7d6/bdlCJn2uor6uTH4ENjk2eQaplNwDnRBaiZZoGjea8Quck
WoW+keRI9ydO8df4Qdy5ba0nc9UEWazblFo5YCtjTM2z9uJ9i8+jKHie0BJwFIAB
oI4PrfEgdOBG3RkXQL9+6mYVnwqZt8j0VZXssTzKeoWzSTGpOr6ygqfBTa+9Cr7z
jQa/c++Ucq1kfHUgp4T4oB2IEz7nceY9boQma/MOIrHGK41mfpfsCTZcsnfMVQJU
/ezR9jzzCTYIC+wLkB/g8K5EQSTLiUQdXCgCG3AhZG/x+Ajn7XoolZ3m6cpTn/Eo
HkaNCEXDYSJNqntIU33+o8gB36GkgdQS/pD/VQIncdSCdYnvVYskdOMeEm0fBTgj
EDZ3d7PYeWBL0ZsF6prlNAshpbDoB94QktwcOKMmOBAsJkDTObXg5ghA+EI3CgeD
`protect END_PROTECTED
