`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LtmmpudcHmSQFJHmKfiKowbftDgrnnk9XzD4lM5y5EYnZ7cAXVJ1nHwp+QEG/AZ3
PSzBhqW1nlnr1GoK9Rhbg27wgOxHBpgC2RIO2enRznWIoXsTqNHcYU/rsf/ZGVqd
NuqfvSbVpSLerkShp8ubAIvGb3yoxDLGEQwzJ1twMkp4MamJ2F/mI4iuigezMxsg
2pyExUTcwpq4wAT3HxjZlp79iboKa6tGwrLPMbr92cLQndKjDmOnWpoxq62fA45f
s4xokI0OSzJedpqbWnBWLWU/0Weh5m+NYJHxlCIWxv6n97myJShftHwN/ar56cVo
PILF9XdYcByms0zK6E1ZQll6gTiiPeuGq1ALLXKLAQ6xMhXIze45yY4OK4vTumKK
6cM3BzktO+qG4bBnXPZZsmhMhQ6V6yXtnEBY4iU/pCPIxg9okeerNLJgc4WnBYvx
0V53bc4sHE4g33hVKfo5Mkz7oJYmXDGaVj2/xGp4lov/FBtNAS8cXD/N3zO/whfh
HTVv/THYoLad+h1ww/oKh6gLpgnbbO8e/d1RJIvIULacIuRivZTPH2fNpSkOYsYY
6HWTqP0qEDeJMD+3IW5Z5nZl5GHtfiBhdPwYlxo72IiUC6SaefjJm4pWdab1ehc5
HWYjwurcrVJYvKST1fNIPP34PdPqogIq5awkKWbVKYkiLs+nNhHGiECuasNSaJJR
H6lwugt/wS8DekqXU3hTB5qDce8SwZC9nuNWxDH9UMSaUUu3q2b8RgdJs7nRgWK0
9StPiCZxhtZya4fIvidcEqc76G3fU73Gg3MzTq1rwK4lcGghNcSLy3zpERE675AF
gA08YwE68am5TzCbu8aE/QIQrfhYsQwmFq3TSWX9bTh1PsMra8stQd5LZAK0lB8t
DkO2uvlt98fGE1Kei8ekSgL5Zw+Z1LLilX+QLToCblWVy9cVExaxLoDx145ZAPfv
AkdN/E/LNkEAMenMEX5t0FjY1bZyeWn2j8JHfujkgMmQdAhL08BxTFM4rrFtQX9X
26JGpW6t6PsfE9d3QoIXzLaYe9I3YGaPl6YCBmAN1CAF13QGB4cZqTycKtUmdI2q
wfN1jNrXe6JDhyt1FoD6m3YjFgI+BTr8WaCtgv3c7mMfSb0BQlD15kAp5+gEcbMg
vT7icNfI2j8oWdp5En5G9YjiWTKpipPUlYkx5ifX+1hA2Mpb6qAujorBQYT0MFD9
oUyNT81TOFFwcUM/CX1CNWr8fvuTy/obOARLTbm5JyJ3fbumm566F0h92PQlXZjh
YkTtNOAFngXkngFiMdUfaMQX5WzjTrNp6XkgoHZJEN2kEMPsj/585RUv+GbwJmXJ
0k5kYgRUMf2NZYT1rWjxAP9eFZ756IWTgtOIWlYzI2EZZvEFHww2xh4raaBY1dTv
iPcX5tF67xdsGajo7b3cl6jxcir8rpUQ3C34qAImONHH7STEUIy6mQL+bWC0n03P
DOk5YzKJbhn6wUvwGTFakhc7YFcIdFXpTa4Sw2r+i8IK0Mj0Py1irG8L0z++nkkR
2HvOlfrw81YVchzspVnHsQBNKN5zDrBnRfebqkeXZoDMivwmnCQMwyCYNtfrFD5P
UkJjz/qThUh0mERC8raEwoB6mPePYrqyA3JC/Tz45f42NFP6JpgIkToSsktM0Sm0
tZn6LZksYDDjHBuiD4/1okg1GLkOA8PmpWiYNbHdLM8=
`protect END_PROTECTED
