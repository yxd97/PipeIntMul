`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cWllxGGw9HCdH46+/lwNPpU/Q+EwwUw3ysCmWC3mJ74encf4DDVOhJGdww3VBFHd
J7mXylLtc76b2cC7agEujbjXYC/hNWrlWnPuYwmD3yCiWkNaDnDzzfVVXAR4sjym
vtGapEUzgDH+B8BN4EuM8wcCWcFgIf4b2iEH8ZSohMIzSGEYIQncmkJ5B9E0hAy1
F85CvIY47ANAEWypQijK4kL0pSrM77A/OFfQPpydOFt7IaqVpSQN/o2H1VhK6yT9
2GC3EllNKu/2y2Q6mkIk0VvQuV6J/RUCtCb6HYcyY2OrC3U6xltd0ZMaIulVuAVr
J9NpEmM3gsLwbfCYf/ADYm4HrXtp3Kuh7BN1Iv/555EBb+MVWwFed+fM37yYFTz9
CGITyEYF1Crk9MrcT8jRuHpJnpTUyIuUbdnXQBQhF8MKntkTAy9Owj0SMM2IsHx0
1zaZG5KUPUoHlQF3BIs5UNnUiLHZ3+B/MK+tq1zzgXY2HnzSLkhJwemDil8hY/f0
y9H4W85DZ2URBHvyhXRwGOjXybt89jEPXfRe8JHS6lkZcFV8ysvMy3BkYfw5ENX/
H6fHsp+OqUMtHbeeQxde/aZbsFqXpXHu+Ok3R6T7vNUrZbvlcys4girOFBuNmqK0
4kNyIKI5qpxKkG9FyzD2w/XuuRHHhylUZKRO6FVjzyXHO7u5Uy2aHQn+pW0HHPBw
tNbfzxxPY1iqb7JQMB4frw6ILVSfUPIbYhPKV3Pe+tOEsxYVt2M/P9/95m6WfCzy
of2jkFZIshzhCfDdViOzBa8veBrrcVLUSgoaF6umr253C69IPY5UEyXnWuw67kKs
pzQvp0uN9n5iYs43NTFpzhXIJvaSRxScKe1p5RLtNPhPilBqr9XBxzgQZa9gsbBm
kXNccDfJvXnVk6oc2bOI/8fXNTJISQQK11mWQkzyN1jTXGox1eyDXvqfSoGAE8or
jgt2cqNnjyMlfGz9WZL77mrzD0iWfxAtG7IUqQ3yE9c2ID1DdDNtAF4kLuybsgnb
SJrAXklBKqFgYaGLCD+3P1NBkoXoiZF+7wsQAZAXjOyMY32pr8ax5AOfuJN+QD37
kuvnY5GrigvzMHRM8i5z3wu5DLfmumOCs0VKLzUOmyiruKwpwVMvRfa/lP6tlZY4
qsBU3dzoHfJzxiD64mNd/1RdV557OY8ds5g7GnhYQpxJ4XyYjmi75oz7LeWltSLe
xKQAjaH6d3NoYcyGox5V1VQ2+THnJ/+YzfezozOFQfOhQHvhWtAULpuGX/hMWoyq
G7Gq4Tvz3gkwuvL651TtUSWixdFuVxnO5F/2DCU9sCbTzKWwgR7s5fThy2pmeQL7
dWujMiFWuMg2Yb7tcXLlCHY79b+D7W3SbPxNadHeJHFZ42MF2uU59J34XwLuqiJ+
+C7nN+I4ZGyNtRDECMyXIIRDiY51WF9Xrd4sgWhQICm7KtwUeAjwX9Y78eUp07PO
QJqOGjgreARASpk7h0vqsHKr2GQeCYaeSURrZPSUk5NFpx6YzhfGUbM33ocJdwht
yL4zZX5rD/3lPnTW4AtbtXztKbfsTRGjG8vhZN0MbONHuDyAJFmDWxxkDuoh1Uq0
f1DEqmo+S4tarf4w7wtNiJCG+6ufxnNoErXhIqKTQPLFHsstMl7hlnZ0hLBVv527
b6moZdCDlSV80Ljy0ob31svTDgrw9/dwyMVhfC4K22F99DFcVsqDhRrfC+AD7LbM
IXVs8GAfbBMzkEBgf+85yTZYvy78Ua+46B4eR0C0mQDZslgIMBiAlKiRctNRDkIv
ZlMLN+DV7rE8R3Z7Ujt9DvCjuleIisk4elXvMB/HT3ga4oL+Ln7SVXVxGGoWTCtN
x0tOTVEjpvH0T4OlpkH/REB9KzkukX47+1CPk5g5BFbAKLAyAoX39/fAxVJSt8dj
ODcczNaf0RcEydRuiMfNWw0xjMw+Hklt//5dSp0dNdu2cEkuezI/2ZCpDjy1kp4x
6sSv0c5Mg6AEAiHcEHovb9u+ZR3TxrGphFPQMOgLFRg6eoOipxR07kz9EcQ10Cpi
MbENSZpyQs8uLiWBI2EnqslPAQaM55TQmMj8d3GKGhFE+yGxf6E5y1QgAvmRf79O
RkP+KFsnOS3QhbUqzvTTG02XeBaSsbuSXmJicEXlZ8wyHEQldOQ2KaYJy3sWeE1B
ooP79aUH+5UufV/GzEFgYmNE4L1oy7MuMqxwrBzYvlITj07h77yGol8BXp8fEIe5
`protect END_PROTECTED
