`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5NQ3FrMhxAsiu9cOw3vVEH9H6RXtfcjuV1EpK8hNfrErrECLbbb6jJ15B+JC5xcW
YGGJ96dzr1tltAE+XVrCOiDV9ZU1Qk12I9/BT7tQvMNygNX1o8NSXXNpchF7IdYU
c4TqMrTeUFvN2LG3HTs79N2Bzo4ZuVGxCZeuuqPEJzPrPwBDepJLtkXpyfjJuzXI
liJOMsdSPdRn7h/eRpIla30KvK8Fltqdyv66/xl5U80CoGDTO5nBece5bhjNvh1u
22tyg1JUqHYQNXlMV1B8UtWKsAJSk6oN/ne30JfTdhSZDYUljea14LtXAnhHoafe
i5HldD+FsSz/FpoTS4B+Pz+yK2phXSPkxkOMJxDtaWYxu/D6/hYgHCopNcN9ICCM
JoaPjxUWelw2nyBijWG1sCCpI/jHqc0EJgq79pGxmpXx7KfNlBJ0A7ga3BNEDy/2
7bs80ZNfFkyExnRXRzGqQmAO+9EivsgFQuVcXnDhs9whYYOpfQW4j0DuhoAXDKw3
`protect END_PROTECTED
