`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2C9DbXHkgdw/pK2oZgtVESzqrDAdlFpZ1tCUrchneAh5xH5A1K9/AWd2Lr7+drrA
b5F0zBr+FmryBKu2Yg0ANN+8Cd8DkvOJKEsEzvxg0Bx1KxRWD8XZJQ26cJ3kuWU7
dfcv2/5mqBxFzkD96O0Fz3dsENscYER7z7SSX5pGN1+RrxgOMvo4s9HxZkRPz3hg
YDw/F+tYoXS73SB9c/MPtsl6egertMW6UCAlLyDM6C46TaP+CUDRrgrwJnB926U0
TBe18G+J2IKf18TrcnTkPMDN9v3L8LzeJHoqTzYmSNwiuYxPEfyZroKhSdRRo4zg
zH84cF0W7aJ9BTI/IckXl10WiJkOrdje61Gb+pqFsLCspNse0KNg3F/psea+PF1T
+ZBYtMsKmvkew6Pmw4oUSetBrLGU2/XmDjjwyJocfEOWmxpO2lpUSkKJx/0u/anp
MuQeMW6DMyS+ZwLveIOJyWBNnq8uXDx3SMnxCkSCu0C0LPVutWz8klV0OfrqSMa9
FrLhmM8AB9tzE0i457BRgQ==
`protect END_PROTECTED
