`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MoO52uZrSGs/WpnwCAC7l6jFIwXA8YrRGLWD5JPtN1pZPD+zbBrslLCRCbhucW8
nXvPUaxXbqITOMKFFCrdrPUzm/rfbz2sXp2ZLueSMRv0JgFzZ6kf4HaIbyZXI3F5
owxLp2vaJ+ezYQmsu7HXuyZfwllFzbDBLF9gPJpoPiyn/gxTuTWWGFAmUnQfX/Tv
JLReB7Bsui+P/gaRN8dECr8Ozds4uvC89XNSRPOj7jaoxyNRCy1VzI9u+XsooECT
DGvUb8zrdVWo2C01SWkPyWJ0Y+4JLSUdE9ruibN6VJleqs+K77EhFUJpSuYcRIj1
U0xtoxZicIv1rY+SISAyo+8/NKUiSw0NflSS5cnwBpjW/zegPF0JN+kd3Vjr6pQX
OOaq4LlwWfb1baliKTyiYL378YCh0xzgCrjpZLKQvwXgZrwedbVtvy5bWemsYMXN
VM0sBnXW6XTQZ+qkN6rbHh07zg5nZRxkMqQ/umtxD4P8OjMWLYXtw45n0gsGeqzs
OsodssAOw93LpjaMMMOv6itPzYjwA5fZncKlnAUQhtAB7Qvz+0VL5Sdh/KPxU/3D
GbCDfc7KAMjoZbQFg3bG0K/vkRYaJsYT1fLZJDEinNxEPYiA+Njo2pPpMT5/Pxxm
VY0Geef/qBtV0eFi/rv4O15l8rzCOOzPC6FZNKr35NkVORI6HhaQRHphkAQs/565
Uk6cbarz+/ubFVLnrKr0Ay4K/6yPY6ZKIYMM0tg32zGYlAV00FFYeWsqiaTWoAen
syKlcO7+SyBuhngPMlRjZCyQQAztJ8/Lmc/L+vBZ7OSw3Td0654PL0VNghkxBgPr
VByGc5xaYL9otXflKtXolAmInXKcQt1RwhY9YX1iH/w=
`protect END_PROTECTED
