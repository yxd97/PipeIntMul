`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWplWe57IHK79z7ey0kqNzfm04wy6RzRDaOmat3Mui7miGiUkP4FS0aJruV+kMfK
MuxArRPKxgFPDgLOtRW5TMq7AHFsTXTZcN814/Gy0cgVePoQ845OqoOKErrnxVGL
RuWSPFLjYAKIpt76AHkFDy3Ytzonc0UXc3i6IUGzGy/19VJgLtsAPeDuYpv/FotM
KAwqUEU/qAOQFjn+tR4WUfH/65iDhCMt+D77B0HTwhJzBM7F0GVvPvVoWeqD7u6r
mlrsgye0D5zp4Yyd6roADiXd5YragTtK6P5qjxIifo3hraz68uJ2ZHE30yO+3UAq
ui1zJ/tXAEbZ2VFshQyUtA1EbrBDyOQLP9H0ES8icLkDuJBM7BPNRO4ekUv4VVwe
dA/x3R06ILohF9CJ4TKr8BeagRrjE9a66yerM5Cft0uGY6WP6gdakxVFMPKZjIYz
xAw1QtaYLOrGY/eguoIXJl87bjaBBbxXgLuUFSHrbwz9DpcmmCwE8Va8MjtHiMNz
Avi3gg/8nAfiiT7EtKZIe4Ejue5iD68p8CgYw/I5FcQ0GxNnPruHG3xFHDU5esOm
ZqeoosMY7LA0LLSxydELa9TPwCy+h3GzDXyy1wzLPq1zmGh9bhSABXZK459DgyMO
PcS9hWDHPMrCYck1GHs9wDfSZUMmlE6e2G4KnEkw6WpC/04BNaBIO0CiwekYO0cG
NqWSIaYl9+lV7gGHS7VDsowQ50uO/HUpwEANyGzoXDB1m+NYfkee38nyv8mHLhHv
E0gkC73avkCUwbXVl+Ly/KiH4e+M1gb0qxFl7sfv5K4CJLN0u8IsksAGF7gHpHhS
LZeVZfkxii7OWh/e5tIi+A7F6P604AR8APCrN0V39IRD1RyMJU4QAI8HeJdJ7li4
XOJw3aiDOFkZfYIqHCDGgKAcbliibT2fLnjXZiIh332MnKHdqe+dctSl1re7iQaX
cLnKs6ARgteOueHqnQn2O9IVimNhqQb+g3JGupX/L7bXgB9LJhRBEs5/vumZbMB/
VFdo3ItwNwE4RJ5IlwJ2Hf9XQbOuSUbyCWABVvTlBzXCFVM3OfgobIltMniiQBo/
jZfqT4o4qAf+6ckLL96MUaitVPcr8GsLSLN3iY2Jl6scFNVV6vNw1WeLBuUBRiiz
+schpjF1XYuANtzG8u/WtGueKg8tBAG3tZSYCYEP2kXAZ6R6rPx8YPJeP9UpLWdG
PqAOfE0J18ysHqmet4teO/na2+8icV801Fadsmf7EtRAT69lQTR+bf92lpyzK342
9OVrYtnr2eSZ4XPr3hsVhGxE4+DufiPL7D/HHLERtVhec7PjSRJd8hQurdFXFiVV
6qbgvBHqGPmJYvuf3+WcuWiHDd7ffXcXZY9SocMdGEqYcebx7SLS43QKUzIH6iyY
KQ1uLAPgG5CQVB9dvCBs+c7IG1rf+YwvzbwLtLMTy9/h8FdVZD7B2PBy4k2uY2jV
6NvXNTsA4CfdSOtXy+0bX3OMWGy3eyTHjuAOhocAaX8CN+WwtJfPmFjxmoPzgM4W
ZCGO0mPPLki4yQIcm1jxaP/+OS8qfu5cgSscr1HbqKM3kpV7hBTXSp6c2XpG9kr5
sg1yEH7L2GT2OYtgDITF5Q0sfwj8WNduUEwPUDBDX1vR2ewBaVzFVWRuyloZRk86
Ok4n9tWQrXTFMCSXUAyeZXLEICaYg0nUIYIEjZtk1S2sRd5JHicM9DdezRKY+nbS
G74pvU1vppa70ZNirGHdEdkON51EFtLC7q8MusZHzMiztsj5D6j0WIA3IyL9deZ8
zAuTfP1Syf66MjFDCmUOD0o2JAHfeehhn5DmvdOl3quc2Dd3L4PJ2MdbWCRV1bBg
+onLTn5osRQY/LrBEFqUKRGOavts73Gd2N3UbVzPMxRLJAQleElQuLZb9xKCOiBn
boYqMlbZlwUZ6ItR3fi1cznlOzCtbl8uz1XhPnJ1D6KQNOpBWto7ymGFnAe9dsIO
m/89HCwZiJFzESGa0Zws9bpo4FY0UCp4QUCnQX/ZCH49hMJeiFSR2O6ERZRXCGMJ
TQk90MNqSSFqnULmvFtA1xE6o6kNH5b3RivBKZdOzpReHiDET5jHrkqsYGPShG06
QkyNTZnVsthHK8lrAZz/1+Z8LfI4hUb+vmdH7cA6Cn2E67ne0jXjMaJbdtDFmJjP
EMX44JNcnWRG6+uSHWUcSbs9wvI37wjRy06eF6zXxoieD4lFMcTS8s8U9aGCyrcV
mp8y28Y2GZl3AwPnHYklGv9k/FkYGmAUSRxYj8FqrEuNrivwPcHSjQ6bDyf2a39F
bJzMj4ZgODIra6mJYrv443NRYS3UvwxVTUJYC3febP7I4mg50samLA/ty0E1vl6q
cVEcTwoS6pBL6ZY4Ta+nmdwrBF5PkhaGM+EeASHTdo1811dIV4x/hJ0nghOg2R1W
Z1tK6jWQOpvbkyGtWRGs9OcsdqMsytsaMnWZUZNZY/DMdQnW3pcSPs2IXQzq3n5A
bTBl9M77FIpBAbeNfedk9th2fg0h3s7YM7yWMexvWDxdPoSHsN09CIbGK1R1hyvw
MH5DMOLw/Gp78e/IIDveE0hpT+PH4TAq/q/up3hDtIsBq5BxVnvEJakM1TU39/3E
mOT7sAO2Sev23QzJavYoBlInQiRIfp++15mAL3xaiLvR8f6oesS7EcOjYZLTE0e3
cWDLNwAER5pAVRt4MoqPkA==
`protect END_PROTECTED
