`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+W1E5/VE1LPgMfn6/2vZjgQhIBC7+4Y4pwRlJvQ2Tc06i3PD4mm12EZ2Cbh2D75
DPIAaPhb9u7rcuvIYBT0y6iDBXHoH2Ir5rKbXAZZkSpFSbwYir/Z0ZoisVq/bjdi
fkJiq5L/jkCOTWnxwp8VB+GN4zS4HvMaABrW5vMWw2rS14Ah810ViAdkqAETnQ2w
Zro4cSj+Ef5ssWSgiDDkTrHZtEHa5RW5NwUtFGzUw8c4u51vh2kuUFyUeZOdBliU
+xFSau65VDbD+30Fz5uLlrrq4XwsG80pgY9PzwgkBXL8Q8LWLtLRjFZRiYSP84Fb
of9OfhGSVOgshDSNk5bgHx7mWxCZtCXxj7R/edfsrvpVyMZA2S4rlo0yDMkXitZd
sJzXrG1MyZJzx33vuJR5F3hGjHZ3ycimnPMfMfXbFrk=
`protect END_PROTECTED
