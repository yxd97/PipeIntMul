`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeNkP80bbKFVTb9kBRDRYdlfliX/wDKu7QOFybBYTXo7bePu47U4hpJLdYxWUfhi
djF6RFg0POldQrPDPLU5V1edxeBeG0ssunsKxhqqQhVeAkhg6dudAZVeU2j0Ufng
1jxIyf4krgcVS09MOWBIqz/ZVcHkRQIbyWugn2c8v2Z/PkXUr+MGh8//5i+5hgXD
sRl8VAX2rAHCb/xu9jw6C3eGJxYCqDq/UfCeE0VOCG+eDhyse5vqDIpSEvtOrAPG
LkJAs1oQFjmcs2/ot+aj+RqAtbPgCFT0/OkJHoJubJkRbjTYs3UYN4ErTXIh6jMC
c/1UCO1xcEB/U8nNXNiW4Dl2oohB/sHZkCawKGQ8SS4yrLEgH3dHPlQYAqeWMCXu
95ZtFbeIFidhQRYJ8jlYV7pQ4SPffqB3EUG8dd3ldbDa01ygzUKWB8eZgnRwb79y
daBsDA58N/xPk7z+RZ4z0szSmWxlIR/gstFatwC+DaxsmLKa4Ofg0ubvXpcaQW0w
ElxsKMe2CzAZJWDLq24n3zwl3VdlGbbCc0pO/sMVe+p5XFGRqcYBavBPJ9zzWiot
h8fS4UPVVuV46qX57cp/sW5KI/6swY2MSClbjTUZZTx7yt+Mx9gUyX+2hVauIx19
AdcUv10xRUqJ5wtKRbys4gRMJOhQ55zrhjnt+YDGNZiSs3iroxPga8Qj6DWkjxn0
1WsZvLOpqgKOAHpVgvQq0bK/n0QywMynS26hVUdyz4Dj2XsDBXck2HcYKQsZba7R
rtQQUX+1Q4dxi5XH/BSvT55slX8gGwsU7hqlyGoPDeQ=
`protect END_PROTECTED
