`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S2w/XUV8hKfoIwH6p5wrGT7NzCA4DZIWHjj7RH5lHXRidAzzXwYO+awd433etTjw
dGLSzGBG+ZHhNblT1qhFi4+f/p+RSLw2QtBzLjTxeUe5rl/04lAuqud7yyzacFde
st58ij+KuJS8ItniyyJtAy1KdkHftR+s0Zw24SUq5jkY3TJmnNI9As2ukdlPhFY1
yKhV755b/W77q/mU8jZyp1S6QqnlRffN1fvPXYVAMKlnrQdsoZjQi68MFfvqWy9X
XQtYsAqUehByp8vEUZpY+2az9mpytdLFQ6lfhhLNnf9jD8qxhMFpOjflE7gJMLlK
Qw+e9Wp3M3d6j3vF8+YQ8A==
`protect END_PROTECTED
