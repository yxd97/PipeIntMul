`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbqvYnsnneqEEE9VjdMmxxG/r9dWFQfjfcl5tI1NvKgYqqBn4YxusQ6qKU6ytT/Z
e+s92XxfiYA8W1Yo5wx8JkfzV3fXKPwvzXsBYqpM88pQ0J/tBILW45hQM7EDIjlm
ph4LSC+qlslZ5YwNxstQn23Ese9al34vR/MjC8J5BYngGUs18Uzsvav1kOePM913
WgAk5ujxHR/YFKNRqS6UVdJ8t842tS7uG/SQKPXlbvzW9zxp4n17seyhV9JhQ+11
tsyrEw/KO2YvQ5Hzss9O2IzgHQufVj8MH0KgPpJuRB/hZ8IxJ2/EtQLLH3mh5ztP
rdqjbeXDwDQCHO16azgpIfO12+EZOmNQCpyZm+9cEogHdnNh8NWMn/XLAzgV7Ur2
FAGbmIOJWhVopnaINBPH4QxAsE7zxxYHuJYs9FOCRmZEGNoz6KkG6aTKZp/tc2RZ
yQKlvaga5btj2gYNKRzOppHkG5EphYyaV+U5i7Y69eRDU8Og5ayyJMTjZgz7xF6A
66UwYVHMVsNRDzkN48JoWVb12cKr91RmBwZW/B21uCcGl60GNSI9H2ZzuxEzktKD
C9Rj3JPiUanQWW0RgaZ6YcWqWEFEGBqwixk6JRhHwQDxEjxGQwAPz03unnGHJAvo
KHUE80uaozQz9qXJmYVVp6snXYs+w7mu/hWaa7O1riPkHNHQMqj4Boh4dv5NqVFs
1p1dfHGNIAchRjmMT4qGGwdobDaDzanZnFXyNG0nuNGXikFz/Rq0hGm/Ebz3pqfT
UqezLVzagcAZ6LOMfcMMBw==
`protect END_PROTECTED
