`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nu6X7Mjo7uo86t1HC+k0TX+EsZUu8d5tQd1RrOQdcVrTN0lpVz/hA5exvQDWX6Za
Iitlid6toGc5mMKm5cv3day/Nl+NL586yngEc04kB0S301Dlr6PnMYKJP4tLIA5j
ojvEweBkVKJFvWZToWwoZvM/dn5bjZ/J675+mEa0LeO9xJ+576/tTOV5bJo5wyaZ
Ua56iYqL0/eNPTYmYJCRMNoE2VFDsh7SlmpIKYdPpcaNUh7gApinYveWnxs0wot9
YaJir+Qt4QlHCXGXrXbWY5CKNev0BGiPEPfvxEbxj8pA3pxHUhfrgjFnC9lU4zhT
T6DOv9g+ot5sa8mTaIL2mNGcFJf0aNEJC7sH41n/OXKK/rMy+lBjKYOoP2jzHlvR
i7v5+B+mDH5K8pXq6hHoTmUh6Lfc6N6Ffpxd8+PJ0BAwk+Xb5UbM4ohmgy9BzHHj
nQN9vFJ5ir2dKszYvSitTctRf4gH79+NSn43LIAqSChcGNZi+Jx5ZHxefU0ITepb
FM0pi39bbO/NaM8Ym0e90ZrDgUWPFZyaZ9bMlSqm1b88K0wLKh3w4e/m69HUiW2N
VCMYoBjJL5mr3G2KPkGsAzJl16q1iITSUY4eJ4jYD/wiDyPt9JOwQ407HVgcOkm9
Z8F2A2eIojwVe8Wj3wrV8h7TQZ27YGyv0O0Zvyd5Wf/nbp3d+PUMt0evi6qwLNSp
RZ19W5Hb6mFNQzeXH/OWaAzz2qynbfoIk88+g0xFMHHPrrjGbiFhkA9TyEl+xhW+
IR8ywyt76PEbeggcqwa0BEnVVBvJ4RZNWnvZTOsbZ+abX00G88vL33sjFxxgX80O
`protect END_PROTECTED
