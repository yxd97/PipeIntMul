`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2RN9i5Xn+pBtGwtOfRK9bsBO1LHE9kQ0UyZ1K/DMHnBJKomUSuS+GlZlSVSPWpFE
JmoUmpm8g/wQGS8CeadLLdB7ydawfJprQik5SWG0sLQXyqN5Li00rPrwaYP1wyr+
3Nf+Nt/gW7PN1aScWtv5hzWuLwxJLsFSj5SMuxIjmd9DWfCywhI7D8zFlrVISGPw
18OSQ7JM0SvyKqN/xwJT0Tr36TqRnaj4q4bBs2Evk6PymkWpeVPWDmXFoA/3XGSu
VRvmWXcwQ4s+Yq//t7rl5Th4qeq29BQyMhRssFh6iQc7LTRhzvDvqf2vZPsziEWQ
Epkdp0Boi0COzdubyvmiX0/2tMVvfPUaNA/Rby1MSiYVt65xvYWiltyKvU7/eFd3
5790/IVI46KEQ/FRaIzmxl4i+qkhdS0jp6utLK9Zb6TOTP5SiHePHQJ3ZBFhSMbM
uaZJ5GZ9yu2l9gm9QqKCjUWK/2q+e285oBAP9NhAZDQ044ZYWikohNpKfEFcX4HS
SdLekv9F71ooLut7h3SQ06UR8b17g1y5X96AifPn3ym5d4LIBNVdpl77WmneN+OR
Kvvc5w67/FLz7uGubHG9Sn3/YE/bjHv6Q+xe3pxWBPI=
`protect END_PROTECTED
