`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4tFlSB6SInsGyvHlHkEIDO+OxTeeQyzPz3TlcoBItd4x3IdTQdBwV5HM/ECbNPB+
jx8AQxDfTEUiTv9ksFu/C4OYg6SgVAbiZ5x19O0HlT1CmFnEGTo7pimjlg6Xe5Ii
KDfSiyI2/lZh3h/goESAGzseFpB2ToQSnchIfnqHjvn7LY/ioE4+AXXeO5o8JNbD
7kuBUXdiG3JeGohxOjdSxdsMD/dnsQdu/2xyxutV0Php1dRX1f9pZl5+zHF3RENI
AWcmvtJS8GmGwmvAa981Jv3f6XlLHsm7/ZlmWeniKx9JzLybra2ReDffM471h7kC
S3yPdHx6LyMZJSp9uXxtkMB+PL7AMjQ2+T2U2DhNsTdKVNUjqK+zfxEID+UyhnEs
wGLma2azJVj7+0/BtB2pPSu+VpOkfUYE0HONZBH4KonjIY2e0Fb6K8WrmnQBFe3R
HudnLKkk1KZKqnDENTKfFXTZbeTH80AgaqymF8YN/FLYHU6fKB/Lms7AvHXSTZ7s
IXPHxMB4FZ5juodkT5IYSjnjS/hE7wN4gYTfO5fNN9xoBMoJDA/c3VxvpNfIeUTC
CbiW80CjcbE3LT+7NMpaeg5rK7WQbvbCd9asuPsKNH2FWnUpEckgY7MFa5BboSbm
SJtvEjiwJ8LBehK5Ms7Y+YvdoAUtwoFHehYfV/+ViR6QNHgniqwMYSMITVGoXOe0
r9FIuOcQeqeDA5ZJIDP8H1hPI7wGTADeG0d2qM+Dyjfes/Q/XT8dNEGEdVj7UHvb
WH3BFI6xaBIknHcBeyT2iWyMkZEdrWeNjeOnx8BeR7klRYDy4dMKhwpI281BgWVD
xNYZMUZPB/7i8LlyWSXGcDW2La6oXrXM2vQtrOoKqXFYpzEUSdEERalXbfIbxJuM
IYPgpkJ9Zz6VG+Stehh0a28qkqCVeySP1eVTi+7FlNhCr5wRVCKhYsIM8Q7NUaFV
kj7wmq2WD67059H+/m1AsR7+2tU6WazZ/dcpzClgNhHNLuRmxMgzV7DI/QV+EjOr
xW+th5gnYv6FI6k1FoMCDRHAeU164G4bPzpOQYT8qSLGPwinK9v5PjmKcJQjIZxP
olfQcHOTx5kLzKAtunN5ozNDNq76eKT0Xxw8Vr2y1q8rZNxo/gFcm8SU4kA1lnB+
BesiKaRXgFSZemyVeCSTVDGp+iomrOCw7Vqq51W3h8Lhwz2ddemo5HikWKBy3ZmO
7S5w5WyL8wYE9ornDx9KZbEhc3rjjv9z8SnDmNCbMSqoMjDW74aWXsMs965gAVw6
i+UrJQc1PM3sTQ7HYVRMR75/6PVX4nOqT3xBE1bin2Ssbyrg0eOQTDbkk8ISF3B0
jy1FP3o5A1Ac74BDbIXWClSUHTY3oTbv0y3MVuNS/MmT9DufcBbMclYHNIh4wKuN
qDORt+jvSRbIrKOyubAWYZrOn1nFhyC05tA0zjo+kkXtlg3lA00crUzxAZDQfxhg
ocEBKCd/hC9S9TRtoiOS6/vgxLJkRATRRHECdxdxjMEJOEpMJQ5r+iQZ13mg5ei1
EqEtwJSY0MqmATFfQ3HnGu0FIBbZT2bjBozJHxDn3bDKgqDZZiuscK1j+N9+2RB6
DrNFZ7MuHVkX4LjZ0/hFUDfLfujgUE4dL1vzuXnk/bSbTxIc/IbAK+YDzyYCgW7T
FICN2zTmoxlHq7ayhl9svgcuSS23rCzWfpe4yfQEvmwzTANZhLv33Fn5gi2xelMy
O3ElBG5sKhnplzFInB4GD6JeIw2CnZ+NFmwwrxPdlZytec6sKZlh4cbzvBV2v0G2
q0qG8rNZ0WsSg0DmPuIzCXSf0aQf2pFK6K0OamQttYD+mdMaJvZSf3KM+qywmHSp
`protect END_PROTECTED
