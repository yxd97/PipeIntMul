`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3DPkoS3CddKsfiOIH55Qn/LDeZzeJZOg70sf0Gr4aIzA4wicWQJYrPqbMVAEeIe+
P7p4aNNZZ/nYTfY249ZS7MvuDWQo5dA7yH6i5N+rkx5NfPU0yWwbsVo+3P5p/Qfh
v65CuOlZ54QBgoujxx6p/d4vW1ro+zci1uC8n0iTGnPE0ax9FAddYm59P82VNMjY
Khs/+wuZ+OkxD1mb2Kc0dPMFiuYlU1ZuHYlq2B/V6WJnOAQTl7dVKSByyu+kT0CN
PsVf9cZTloo8iI/mwntPCHHH/087DfMXhuYgzaWvHaD5jy3L8nU9hYPrz9nP2IxN
F2MPZ3W76Sbx5d2bvnjtTAANtNg1bq9+l9a6BFjMr4r+zGmjSf8KWuK1mJyDpZIQ
BqDc6+dCC3HeykMhW5IQyAZjGQGt+a28+8TGr/YwTAchnuUru67V1jcLEgVW881U
N5VQsjr2XM/Zr2w1sybZOvzkHQeSFFZWEx/k5duzmUWdOceQF5S8U7oh6dQ+ep8+
V0Ei4IqV1B+rBbPL7Hnb7RxaNLtBjj0Jd6YuS9hAcrZURXEp8HBILeHm29A05L96
zsq62ksQUx9/bT30UO5QhlTv5Sgye75eb0MmXZ6+oN8isos/Gnw6OpPY+zIdWNSs
JOyF2WHM4My6O3eAOwofalOfySRflSR4t10SO8Tb+wi4zUNadgrleqrZyMaC1oGw
VDQK5FEpJ3oz1r69IV4bihxWv447jy6ZPNp+NCy2z66BNecagVm+kqHWYzxwcW0Q
lswxthm88Laamo0Tx0AXkiiExZlOFS6WqqYAgdwirlXn0KEDjfrbC2Z78KZyzAA7
7LL+1KNkxBM6rzo9r0VXNOPrSaqI8Xy+dbRqdv/am+iuvY1zJpkZSDxpCzOQi0de
MGBSHdmFQGjWfEEjenfUjnd+b7vjjammw9C0CYDZjdOn1mdxMC5cxwEzcTvNW4Rc
LPD+6leqO3WCjry2IoL27nEDpJaC4ceRB59Vy7RAh5ayVHOZWnfOnyHOZ725z+qv
cz9KjJwQHf7VOILyO1bcZKTHmFYY+/t67TdqQLSc9fp4211wqy5uQc6K67L5hCD/
L72tuzVH8dzMrD5BISGqZKdLPB4v0Cl+Frkc2T6s/Z+NP3jYuhfZc6S77OSXA462
VyVJpuehbxdbKUB7D2W6FhLE2K2cCn7mNsTC0+pjtRAib515jTklLbK6oiAc6ZTq
IFT20+tyyNlymDoLfdTlsQjQxrpGsh7zDpFEEH1yuiqAkXa9qbI4VU40N0XjNrY0
QBbhpgMnD1OQs3KK6W+ga/6valcCE1yhMu4D654lrRsNfGowIE6Ac4cKlYL8RP3J
2LL0MLf89nXa2BBILlAmSM3ZdSOGQrSDhkpy6HVHURhWsaLq9TpU+7v8YxXpahoB
bs1yew2GxQ6auxpCgTqQlfWxk0wedEct7vmlfU0nElNNrmWPW6tqLr7GHWA1GOG1
j1qPkynfxmdFTVpyu9khpQ==
`protect END_PROTECTED
