`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BaAfTwO8qIj/BZ2JmCE8VpRzfDhwzq3AAhGLs0tG0HjwXnmVa8CQMICymd68PfNO
ibkfSHUt3t3wOWkxopASQ8ylaQMLWl3kIZUI4rzj9AKqtRM7TaBs/bB1W70uFkax
5Wfa8QbgHNzYxHnZVhPweY8BbkspVHy8ErkT3/h5tq+v2o6JXWnncy7ZNz37VVq8
+fOx2J1lJY5YXtgR5Laz4iBaCL7l8DkQbIPZUzlLqdXJg91CDNVWOhU0uYt4j61D
J+d+oFXb9MogUul3tLfaa7XvIvXtDz8gJBWDN79XNhlyZ8p4eFaTTVV5AmgXATF3
QMXrgl1f4v+fUY+Q5MwLHzOIuc11KoZpaFj+6w+uI5slzt2dpAGqX1LI2YOVLZub
uiRQUgLWa7K225QrA728MtTujR8e96T07ksXZMLUCVLl2Rlo8sURxhiQooreX8gc
ie+HCmHhpehZFM03SH3Pu1xPp2aLqryeTMILnBeH5k0IghFTaPjwtxeeeUJBllqo
vOER1M/jmc5O2RG5dyotQZMv9/2DQumMX1v0rG3yzpcTdds/yIpH87LpNIpGgtY6
rwDsaQPeOj6X55JIV0GsfQ==
`protect END_PROTECTED
