`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHXj6jv36y+QxCmGcltGw0MwnBIWiQ5GU3PWzGQ5kBezq61HjobeIjLCv8ntsUP0
E+GnQ6f8nttthSwOAtJaGIRpteZajbM6gFpo7SoJ4yC7gKzl5e9AXB3HIzaZVimK
CAXb4tV5JqfjpNMzvSsmz+3XccrFbER6VK1HhjXAkdaLPMIswWJ8I7osj64ebjIv
AAjYWfIxejECGaGOSSFLnZZaog/Jm6qSfgJ5y4634ltpwt8NMUvOYfvACvv8FG0k
qANijCbD8b422I/fVvncPQ==
`protect END_PROTECTED
