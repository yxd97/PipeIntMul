`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nwdb0Wms8M3jffwwhLhhIUoSJCp8o8cP4ZRFpumGN2BfcfOLnQKRbsFEiWFdFCqm
nmmzXygHywQ6z+pfiegUND2VMl74jKdRl4H3WWVrdhbG5wugiWWmbbdVvSvVVGM2
2cU/r2d8T+Zh01euCP8HJW4A2uwRYbzUa3d56Ow7cWujebEFqNje68Y7RVuZ4CjF
snbcHtdWCRUn2yy4+Z2JqFc8j58SfEKXz1qVCHpO6o9xq6PBl4StX0EqgemtnqXz
sQpn6OEacUH9w2KPZQ7UMTnGUupWaLipqROgdrJoeutDOf6kzJNNtIB7vc7+qdUG
QNQINyilf+LTWi4L05wMddwWKJ49a8duP61dFvaAvDk07eT9leXnsJiJgoKy+gWo
oPxbZy48cgQHKeXlVTL4b1iZvopS9OPmrQmImZqsZPJG5NXy9oXPPNHMb+AhBfoz
OFc3gAMd1Y7dg6oep3RRKU2L9oQz35dMOs5I0lrbshffxtopti/ygY0Lwyt4GQOE
Nw2F7DNBp7pE9DcwUd9UfzkoE40t+kFcYmqaIjiB53ahQRliqnK2UhTpESsGmHnA
maE9olt4wTHlRFTN6z//LVtgcsMAE9NXYwutZq0uXe2GU0/jtfxgHgVp+W5fhxUB
cS/UcCfXZ6RFirTNdL5pq841f4hg9YA5KUS7cgyMOCdZsyc6DrUa93VQbfBonXSa
YxtQ/UIj90/bwhJavbDw6B5N4ANoeMov7EZk6W6FTidQ/MfKdLclcK02yvZozcxn
8AvOkbiVD/JAiKPg1UQJGbGYyu3OpqSl21i4/p5jXWunEwQ3ytY3qxQG2BWo6aHb
nNB6sYn/9iLbMag9oAL4t9NpUXeygpVoByo+k6ArtuHC/dEl0cJ+Qtb9zPSVj9x5
VwPrR8Pprv0DTwCVVaFmfs7R3npfW3tfjD582MM5mJJk7fEfWqT3Uv4LlkcLHjK9
LuVhWGp0NE8gHoQggITfdqkmwfHTbnQsSJCTA4ITX6POovYMLiRURqvtEbIL9IFR
zg7pvydkHevq+D2LilvoCbWCoNYlSdrdoj/eYea7LcvZyvfKM+slYrSLSa7f46ja
0gHzGaSl2F3pR5i+qHx0iO7sGRutezmdzhIN3slCf9JY6jriY2Iyy0wRIcJHDDcB
sF3tvxkOFf40LsY/6HLhWCi2tDsBP15Vytl4IJl4YlHzxgtg15mvcGibGa3gMYcZ
rkpf2Z3czNgbtsIBSVeHt3QUSgqdIxbVOr2/GNwx8BKB/GkRJgJCY78eW6f6Qor4
tc2zUqm81lQZJonh/jUoV5I/Ew7pFZvIcUkbjeMB9X/ACj6bOG4kiBxETrj9rGTr
Ho4waVfx+G7T9J67mKP/DITxAeJITn6lBCEguqZb9ztp6WLse0V9ADBCeyCUYuGQ
9X1Ip0i434WMmSZV+w7ARlRh0UjMLADZPo7v9c68zCwJWYs7W5L4BrRl9K+twq3M
MQmVS390Ec6F2/mBmrb+oIGtRJenVPA5CZWFMZEeAQjiIsuwsybdU6b2DQNY1o8u
IdqeflYJoiBdoqZcAMf7WKYVQWuMdQxZg0CtAXGKqZ9fVbOQAORy++TCZjgYmpof
3A0EZzrDgioSE63glGBrTw==
`protect END_PROTECTED
