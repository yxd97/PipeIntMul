`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wYLmrd4+vCawj7GJfErU0Ck5Zvwh3h97wWh4I0gdpDx5k4qhy0TNocZSq567x+v
9hYp3E4TwhuGasgYSUIbrT21+B+SsL/Os6Dfl9LryWDGCy5auGytKy7HtnrfqEoK
WjCVef49W4+F3DpukgPZAHK96sEarSJHDxUcprjRzdgjR5IgCJ9G6shmWp6Q7JGb
B6JF+Uvj4LtDiqvZJMfwkseICwYOxn7xRAdEMxS3M2NUt2qQVtC7iuRdZrsxmo7M
EnikSr8jsp4xAQ3Cf9u+tSlklfae54pwDD931waKt1mGwM1Mk9mPlQfzjOsKoEZe
yJhQvvjdaA0Kc6SI7CCoiTFTTi9+0DBd1R6+2G1W+wlRaYtm5czyFHI9JgUh54jD
m5tLOaDFqqUk9N+ojFGc/NTf1nZB/7j/y2w0yG6gECjEXo+OKQmIpe+a3Qo0Rl6y
isrgpnTwqa9MYaopO5+kBw==
`protect END_PROTECTED
