`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xL7PxZlXwYSrcrKwf0O6Fpk8wxiDo/UQ+atqds+F0IW50TXvNaSiwpDgTirKiFB
G/JL/TxPJFSM4vbtNZq5BQ6zeWVIAbYc1dUJ/JhblMB1BWQo/8MJMbAHk66MKMMB
FXGSdCIxnkpV4Hh0JwXdAC/aERDZBX1YBTGhJUJ6GrtcKLKev/Q3PuGH5gU+UOyi
3ATgXQ94DRAQnHFE18bjvoySYsMVCxSVLHNrH3iPeQvZSnR14jS8cswX1Zgyrb+F
xjt8r8uB/eNGRBzodIlNtBwuiOl8KpCNmmvhRy28LRYXpWAIkm3TfRuS2kMxDAYs
foQtgx3kiLEsU/pRl5Xxfhyu38dTC9u4rMOwc4Yf8g0VTwSX1whjuskGb07vcfNx
+X6bYvm0lcI58ZoYcdcDI7cqxzleB+QV71jFFfseRPf9NhMS2QgZRSvfMjM4PO7r
BxsP1H3QNd1Fwk3o+BE7PnKGzmRNBZek7zFm2PYLwOfxurUaZggo4M/t1vJBxU+K
uijVDEekAQhln4XUMUsWU7P6kfNjC2tBw2FZTl2iReEUFuLM+oxvkIe8+JO2/zaT
zjQNjsnjdksUfHm5UyXLIpI1QH2TUNeW6u6vNSe1sXAQweyks9tNJ+QDo9eP6DFB
H92kUP+MT4GwQZM0sWI9ef8Dh5CfTFqNm8mQqgYnARaEb2hEnwz9gnnEq06D93lw
xw2Xb3s/nty9XqyTY+bjs52mwiGeCgghamdpXE6nUInebcZb2GpB8J3/86LcZvJ8
UMR4yjNkzShymYiGP2p+sLV7zGvaNO3tHEEbhSKNXwNZYrEbRZTVUTovv76ex9QT
3NNCsteCZIk+tew9qkmOL1W3BWfS29CiWLiuxHVhZEAJpa6xNF3LVTzB1xzuCc/O
8q5pn+7MaWKs/T03brb2SitV/NeUQuhMPo+2dlH4jd7KtvhVW2CMXXpae8LZNNV9
VcvPrbgkHXqcjEEBo5SN/4QaNVyOS0Y0sk080H6iotJuxI1XK5+Q9p/pPzow4a6v
kn7lwJZs2Jus+umrN27WYg2vbgcp5uko3N+3agvv+GiZDKZgCV4YrqxzwxFQ1o1+
+d1EcuI01HurPEWJ9/rfC37IvLos1ynG/uQX3CQU8a5Y0wKioU5un91HjbpBt5Ko
dB3QLk5jDkGawq1JXriZ+CLQReEcHnsmWIF+fUnNE7biXuFo41eaOSnkELLwR053
HhJCJunfcL32waeYmc8eat8dPVEsdEvHVADmyEmW2BXxlQymNjJ1uzmf2+5zbA3o
AlmedJEGM1gP2ucHbbjWieM5Y0MljlIvPAw+lqs70MZpuXzuk1XNNzaI3RT4Q6qB
FShINC0Ej2VKwnQW4LZxu2ku951zUzRgWKnohsPtUSrhYoCNrBVCM1ehNliNCNXS
Or9JoBxdiqOsj/dBmKH3kUlslvEOqTfZ/kjjGQVkPI4tVlwkkQXpDdTa2u4Y6iR7
LnjFrVszLcEfEdQX1536eBJmZn8GIID0/fstQVBhj/Sf9Edy/Lkpo44gQl2PwGPT
5/RzaAB9VUP1LBd+aNwR357QdsarmYQO7xt4TdBmdNQfCAsuOJht18/G/OrOuFus
tzjP8mWnwYv2lXZdKdEYOxpvr2x6U599CIBuId/ttN3SbloowLBQq9onR+Vm1Y1/
EEwfdu25hDsxKGHATOP3rXZWGznVpc+JKVey/DThwaq0SFPo3dkIh5EwTBRppC7G
mmAQDPww1dPZWVhPnmVRJuBzkEBQV6yGUAr65y6dupa7bw0sOjR+K7YN3Ux7ioZI
10l8BumduyGoLSPHi1uMD2hXft3xyrd1AxgYWhkLt8iFD9QeTeHwbpUCYk7eJzdO
e/lwvUCGIZ/O3FeBP012qCxMQ/ZpNEG6qXOk6M5RoP6o97q5iaJvGZWPC2kPEPhD
aOdm7yqK6wPX8JUsLlhQk49utclliXAIiaq8Y/sMjuEAoBm0/IbvLRqZkafv8H2m
yuo2ZDqf9DM4kVmiSLrdMIXNZBinjDIRaVPSpJSjYz6mA59vj9/7vYPF0gWlEaWp
eqL0h2gTC1rqc2CRKIzr5atnZDz4yf+6J8Q+i7JAeWCdkUtXvC4a2byrVVid0LT0
eTSEP034cecrC2ijiA4MHfemPI7SwqVQrBzkU6I6nw7KzuR8BvG+at67iAyCQM7f
5gzjzutQm19oRB3XxAb8+YFf6i7+c4snjb5NCV9zgirCh1Do+TWdQstRGa9etJHI
7H1vel+xw88FaaDtSagZQWRihf+nicpvbTQgbrn4L+KZzsdCTD9F/3TthENVJ8hF
753qqJ8UF3VeSjiNqKJ8s5EehMbKxLZ7Wb7WeJIXVWGKD+2GFedquAwS5QUufbo1
EAAOTGYJ8bOx/Au/ZYP0IRbNsftLHE+TCW+3/YyJEqH2h041DpPgEeIHLp6y7svC
syvmGre2ziOYNJxhKPpFYOFwVTGOSktprT1P7g8QtrIPj4qHMBqviVTqnY04ciLs
ZRZCFOovDWwwrv74ZnO4JuHQJoXEultNnIa1WNI4cif39XV3+ayap/xD1+5bKMQo
i4f8oovnpYXx6+ISa904cfaN3C1WTH40sLyd643LE7qpKvXlIgMmQ/ZfGXV9Htq5
E7bJDocZEv1xOyHNohPULmkzRXjJhzbHbvgwJ+MMlVbw3AJjDihQckPZ76O95aOY
N6vhqpZxAr8PsREJ+xWESK1nQ90wOha3cEZOBPELhGKH5wEKEtN9cU9UpeiQW3sa
ychXIXBtiCdzYljQDLcpNP9LX8NTQuutYMKgRYzv1hwGHGIv9tTLT0LB87eIQiU3
MQC9tfnwxjJ1NmSQGVQ5qdTdb3ED5WktH+Jk/0p9gKTtNXetfx8sz9I0izjmBWNZ
AJV7eUPqBVieuIXiA19nGEOJ+EqB34XAVd1VACuyr5grTbJCL38QL6xio7zY1aSP
5MRybrBfxSqWdxFIAXCPLjRDw6pKofqgp5KJOP91NIocYDA+SAdElrQDwz6f+ZNR
9jNA5fw/vw2/ptMaIHTIksFTYlB31NnOwGgqtZj7p3ziWdSsZq43HDN0mpa3VfMx
rz2HEfBEGuDP+1CtFC4qwk0JCYazxv1W4+xwqnGNyh46wTiOsv2hbEc6qGJ9JXzw
MofWGYNStPjVXkrS0H3VewiDYPNF8d8G7VAPW+JnUvLNSucVtCTNleEGFeXarTZo
QACbkZKiBIH89zklv9IPgWj0dNz6NafJYVH5dfTgUG48Q+usmhWdDoBUnDu9BqQB
HidUIAeCOPd+G/BldybAXq5eiMbYrhmtyxuOPynpsj+/f56oHVnfcypyPDSh1lka
AzCGUcly48CoWogYiVyy2Gycsiq1URfn18uAWv2RHoaUCn43d0gA+59e0S4yWosy
VSzspGbb4sGcuKArfOvbp60qcwx6SBkAxQ8rwY0Fif4I/FmyeTX4zA73nLwd050Y
kNFc7M7sL8RjeSvhMYY7nw==
`protect END_PROTECTED
