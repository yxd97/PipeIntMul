`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CYUj6lYxOs/1YSSckgpE3ffG35nfN6IYXVqPoVcrvSn4w+XN3WdXhzsxc92T0kcg
619dpF1+to+aiB81pylN+wCE+q7djX08m9wcezkXvQBIABpeqhgw4hh+UZjqIJFn
cSJ3N55AC8zTsDGlVZo5wXW5RJ0AlutcEGkr1/I27QH5YmVjvsxBzLTu4xQVHhSp
CiItW4ZMeLU7itSCOKxo7P/+Uluj6JmwdAxP4W+QiMVyY7IY+4aL2eI0T/+izBdI
mStbZPKjW0NClHktcpSTvW3JgRgyLMc6xwW+ujoX1jcaW/lWEgvIXIa/hFceNtGk
7v2iuGv+5yGAz4q9MjWy7VRoxlS/u3GRU8zChkf4YAmYZn0kj9NBI19PLFnnTw7m
Ey8YqGxSx5BxgwzT/qNYOQ==
`protect END_PROTECTED
