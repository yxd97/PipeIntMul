`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4S7Q9HQGGn7V3XnnnALAdpWcLmaocSFXcP8FnV7bxedtVhv/wjt3q3Oz84PMyfB5
EDsBR5i8Q9HjtPvaQGoZNaI1qx3m2bTHN7edIgZkY/L6eDuyXwgoPKHgt16dxvbn
5BcaHcbBGg4JATCFu2/pv2wLPNlpOOtLPVyla+zYoVhJRE9ULh7IZ4JpsSJAjqk8
rVPM56Lj0m+Us0iGcC0MfGkdNAOZy6rx9IpCgbwM6+7ADKzdBiasE+ZYfgx5PJ8x
zBe7kdskF5bp80FczyUOPNfJQExpW+pnGPIPHSUd2aY9Pu2Bf5tlKu7QCjyBRo2p
Ptj2N7V0ci628sePNMXyDWOUy9Ij7CzsOzvil7skgBRX3HraDroy3+Ta6CLOebqU
oKWRzd/3AhdFIRVXcWKvodYiopEkGhuIezw8PZ8UHs+CBnWX9xZL0gaB2wMQje0p
vTbT/xRpztCRjfw0ICZiKy3xifU17ym/VTrkHY0WDb3PGfsC4n4P7c0R23ShNqvc
35NbeTK/RDIWpiVSBf0M/L8ZrA6D+sVr0eyv1e+7ODl/lgJCo3HALz/dQxaN/tWc
e4Zl0WVHxKZmboz23C/QJP05q23pKtgzeUS38C0G7lOecyjJuOAa+8ZJrNc4SP0D
MfW1jGMb8//bfNpPS8gasg==
`protect END_PROTECTED
