`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1CLDeli1bJfbSKVi3mCcBG+14wC4OuBElE7qX7bPW/4eYmHP7Qbl3j+QvGNq3yj
iYcHhPASxdvMoP5CMA25f4e/EpBOPo1NOVzln9rJAR6WK/WBWq7UYh2jTg4wSBEn
JUFsEmccqqY3y/5RR4OK2cBwTedW4wBUT4w0mnbgWY7Yy3G3ohYDYpOBK8v/ZVtd
D9qEmYITLpuZtREi/rX+UthWIZL2iDooMMEPANGUzcQXG4YxHzz8A+pmreW24Ubx
JElS7qGeKUf9VEHlUUKSQ9WLdDjCnlQrFXiAfN7VB/NLEKEyfznxckM3HpiMt9oU
Xa3lhpt4ofIusmDlwTfC6tP33aJvfWL2T02HhcwPlEgqYLoIOMlh3QjeQI+mMkS8
Ot7tarLYmYocplqIqvH5qozCWQHXUB2W+zvIoY7wLhcx+mUUSd2t0BjPULT+xGFC
F+Dqpma79bX48HAlbZG8/y8rQwTNJalMbrpwIumHC39oo4KkBAvfX95PFiQ5wOb/
IsRln/CCEHj+Nzh86dJiK1JUyyCdqxKxFLBBeVZZZnO3//z1mKU+nR3PijL54+xw
iKKSeMJLIETfsMVCJgSbzskjlNrH1w5TFayA+3WwCfAdch8eV4Q+SXcmcQJdjORP
j6IpLj6ejexgC1A3F1MRYgytk+nyKEv0LKWDA7LOPCm//bWviiI8xy9f+Zr4Es9A
`protect END_PROTECTED
