`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQsjoTgnuN275U7UY7tZHym87elUNEereWjwT+vtf20Qbtuk0AMEFa139jHolVr1
vM1T20tibARbUvv8pHaT5iKoZkftDLWurY85bOcoDHYbl6biWM+8gkauTKi9KEm+
DRthMWTGl5s2wM8FYjWLwMkUSFSis552dFGvKY7sRS8nmVGFDRuFFnn83fDTrY1S
oZEaW+/zjBayUv8u5q0CrjSV18AQH0DnpGqQlZp5dZaGEi+J57g71xz/6FfqjQlL
`protect END_PROTECTED
