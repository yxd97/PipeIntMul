`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AnniTTHK8drgxVOZ19o5mtOIFvtU+4WbEKXd1OZsoxvQPonrWCvEcWkR8rUYEkNd
FNZjmEuC9VUMGiZaeEvUrMiJn2cGoR5f7PfXHVj4nE+AvzxFYqYSJcbwP1yLK93o
2X229b6viQVJOetLVnT3gGDC6c94DBkjnFHPmPJak/ulFGwKwNcAVgNA/sPFGLWN
oYhRgjW8whIbqUQr10/f/wJEXnf5wxsMTYOyaqKABOqBw7soyRPJn1nogzc+Tx6o
0x0Pia82EZBQDP28qHot/J6UPFYkP222hWPKcJ+3xwOHMOYdeWiuHJqogrCcrF4N
+nTr4N/DEXYEPWGxcwL26E0ZzMZjWWjjzJ/JcH8+WlcyqiytDJGskLl83+Oi6Opw
UKQaS0JTTJPGkvJE/6j9xAc5zIxEvhY7NOz7mnqmhBcKKpsA2aQA5SK6j1s7JP1K
`protect END_PROTECTED
