`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbIjFKMgCBIH6eMq/AD87mHuAHjjGHtPk3xIWkZRy/686o3GSAJppt7DO+tjyH9j
jYzyNJGCDAf1/TRbrXf/yhirfKggvpYqS9K265tVEOWV2eh0vipMUIFgbs5I8nXX
wWGWplolpQeLSddQoBNjgjM7Z+JJbUdkENgnmVcla4JasoKH67oeJ1qnjHKXhif1
9qj3BZic8hEsoWDyaDPF8kG5LjjubBBn0q3XimueGOR4DYOqVwXrnptd2OJw1icL
N0ExZiwV2LUXJHhp1PLd5sNx6UT+5hGn0hY0KrqOUfngu6DtR/cxfSVuiBkksPzV
eEo70skTd+1RnoQvfm+0XSHvGQgxR97KOR0l+n3pFvvHOXwnqcSCE7/4KFqMMXoo
wDocqrLEQOE/9BTquKWKqL0FRfFwqmxr25nJcbAjxy/eCav23YSOv6V8vqXIubwG
hIjkJ7OZZvOlRc8kASXxkWR6QobP94swvlx52jCHFVr5M3oNHn8kQopS4PNvw4zj
N80n6fjDXMjpXqXf/ZT99DWp+f2msUEx/KR9p0i9W0XGuLjpOeI/DzIGsN+2N3aP
JPU36SohBIZMPUiFs8WMNhXAhW/MHOd5h2zeNIRRkauc2BsBdOCPv7DVee2IkszG
oZnBnRNntHlXSg64IftEky8Gla3jqPqKOFGTdcQvqUohW9VOFEuCDZD4NgWc/Lai
8v8fggwHY5yfRGJToWMVuSXy1NvNgqSYMOkU8uUfik5aqPmR6FpBKld0hidzrWyx
6ducPgDPmDJtAW6sedrH46MHbST7CqYC1jA/40KIjyPMpLxQMJtLtMAyYrg1+toz
k6Fc4p1PXJzKAhBPtDZDTyCkTYCD6kjTrjAUMP5p2fQ5IC/UpWKjDcKZMmRaHDpW
sWkMtRd/9OkGvhz2wya806uXrQ1HWIupMLJWHekVZAY8n93WqcxOADJkvNgD1fK4
nXQKapLv4lK3/yXMCKEfnl6hFZZAl9Gl7wvRyaj9oeyhalLUgkUCg09j0bz6iDSU
ZuoDd8RZdAaPLdCERrU0Stzgrrz7Bv9Ksxozzm4CDD5sLH1L/3VTrLNHDdHKxv9I
efNgzJfQkVQBty1Ua8SDVkEnl0cEdpGMfWJrYc/aulgxRXnMB/RU3Dqq7kF1XVY0
enAJbyTK1I/6m5uXMEouWLOE8WJk4oRUKgmDq2ZEPmq+cwp/a8WRtF9srRaqTmke
w2iC8axCR+c3AEgOmmJgKCAXWlHjZvkHmqDeVW5bEc1TOyrWN0SQ7MJ1V+DaOSkl
TfRQuuAIA81IPveinDjbCgzs8Tg/Z2thGoZOnihl8tVdDzRI8apWOo4Baws+vGm+
LXXEmC2j2CoiqqI6rjCmU31CMMVTpzzprabawX8wLDUrTWAL6dU+cySeaNysR2W/
Cudc+f2SxvwMQDAyyN3Bkkzl/sq0TX5R0tUq+MeVW7K1Izk4Hf0QVPlGtx0HievC
zzE+1MYdZVuqvjpu6N0aIFQW16XfiEPa0OgLXtc3lTiPub41Y53+cX6o0ykXUCqo
TrbR+GeFznEGQBMfWO7BglfpRB5x7Pr7L0K7HpyVZwwk2y4PsLOtjKczCkgLaXc/
lg+KvYO/RLaVZ7GGi9A93j0XiVvO/3+GL61+JphC5kgnrXCAirO7zG6PsaAVgVxn
chIngfJZo84bz+6dILVubYR0bQNGsKFATnJVrwU4TDM1xLFCLCGwxd73ddzs5wW1
pa6wY5jP/QNfN6X3Y5+wBqaMYrTLx2fvfjQcRfWfA4wkCcACorsw4Zk+bAdMhnEJ
URqbFLBr5lTKmkCEHxE8aA==
`protect END_PROTECTED
