`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Em0xKThbBuOiGAyRUTDbPwqgQgE3mqTur1lq32pNVX++TxLnKpLE+Lp6xVEaijTm
r3vHsEaVcVm8bkf5l0CC9fAcgulQoSMr0HD8JxVmYeFOo0g7yh5gg9urfLTehRqZ
OTWOAYt3TRfKqzWwhNTW5zuKUJwzDRlV1p5oVLTxeij7jzPuRL1GFXuNhaBeqep8
hN3SAqtfsJAO9f/Z6jqKcgynHKWuVq8F5WhAtdX468R98+EkxQ6eUFrnppXGWtEM
WWOW+Kk2uTQtMl82RsabLbD9Rbls3nx9EbW3CS9hkBjynlPLSC+TVoYnOlCk96dC
z9clSUkZy9Q/U/Ive4xSsQaZLG86wA3mwbssEywb1aIbdWmq1E8d5T1L2hdqqLMl
rhNm0dMkq45iQltTkMhiilQZsnHAE1Tq4VbkQd8Wu0L0cAUl8kkdAbvQn86hZZon
`protect END_PROTECTED
