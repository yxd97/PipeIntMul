`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNCY1McEUq0yXxW8Tp7fm+10O554Ga+w65obOX5ZtTunPvvjzBg2spxAZxxpZC4D
8zRJyop4Gw1+7WaAdPwf3Ya5Fmy9AyLECw0H53es1GAJOaxVT0zDOSn3wAmS7gsB
YgAiCR85rAWNYY/rdcmWZsl8t21q1Ul9UfKU8H/0F+cqOQ6XBXiCc2ZmQRw8He8G
CywBkOF01sL2jta7c2XQJ/If3BfFUNoQ+/K6d5FS04XdRE4A05eD6C0y1zNx99VJ
`protect END_PROTECTED
