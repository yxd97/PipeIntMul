`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70BCixmstSF7H1bCaEnji4EZePY4TbRcOiqY/UEsMhsP3cEprE9TpKAm/8316XE4
aprsNw6YaN7/6jFA2WpcuuOu4pjmG2on3dWGE6D7flrTvn9GiL5coZ2XInF5RCe4
GRXMQBYs5wB9GuxmSe1nx82fPo2lcSAHp3Xx5cj7QochcG2Gf99GGN2uf9lJdI9G
4vTaiCfw89z5Qlpt7DC8aDS11FY+FXUtkaYtcydLo3LhcNijJwYW8aWjnYWKvIdc
NWJ7RS0yrcazRc7khGW0sfzf2jta394sxg0RdLh7YDpV+P6xNWeoLsHZcwZvBzrw
+VrfhGBF4NNmhLJrSGPN6NVg1AzT8+EtqBmME/mPUk8fBAnHowzQeLox7/gjNgLg
XJcZD59/lGZU7o4v3o2daTajGGyXVVpLbAz3HIQmHRBNniht5ULKJqjZr7+RpYfi
0cOua+DOZ7Eq/Tbo+6axifLvthDv0O+2c/k1/17VIXA=
`protect END_PROTECTED
