`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+lXJcAa7o8OJYuAi4GpQ9cIWseU9l2x5wrJf84soGc6oPs6htTxgoJIKeCOE1Uz
fooNt9bdtFYszzPHxm54TxrZla54j2WbWKWWQ6z+hrVwN31rHtw+WEciZ0ODjyA5
RoW0VtLAK1wI2hkzkrvDkeFO8csHFadtu4ibBc/nS1tdiBr7kJuwn0Y5PzJnu1lk
DOXVUP53Mfc/+giPHPRcYqSr5tgd+i64JW6v4MvleSGSaNztPzwqpMB+BIE7ESAQ
qNkt/rzwC3MMwbiAqeEo4d12NcBjFerT10B6/F8R3q8=
`protect END_PROTECTED
