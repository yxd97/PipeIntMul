`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9PLySnCwnXJRNgyF3ewkedZdaQB8mDuxmvo06lh9r+iFdFxd407ywp/M/bijB83
M26SU49Zt3KsHj/KdoR7GWK3Q7JGhRVjXRsBddx+p8U20z6eWt6sQSqAL4ZAI+6N
bn27c0tr69dOOKqvD2g4YBTWe+MvClnBe/LlcYyDD+g4Er+XUc11+ShZ9iIpD+17
sJ2SdGLf67os0cWs/Q+YjD9Ev74dGbb7+YcEGHmPqgzO/p+FJNIb7gO7AEFmqrO7
FAStjg14sTB8BUko5hKc+G0WR+gHdupUytI0e3EppMEMCLY2Aa3FsDXjsxFk61gh
1bAKzh8Nl5JrowfYrkAVa48yggNplmAZOtCN/um+JJGxvAh1wIEXjCNJBtgYaNHH
X8Gjey+TqimXzl9fCAMFY6YwLtE8Vjm4c1JerwV8iJuR7vDsO4sRLQm3knqrbv8V
YpbehU1XJygfhdNRJfM9hppBBwQKRhPvT3YWo7Iw0z2GRyqOoRHIKhVs7HPhn28i
w8fuMsqQ12b/NzYygmbK75glkDeATq+biYcDJwNG/cVp7ppc39c1rIxrk0LY+0YQ
sOKzHSPz7IJNOlc0SVK7DRSIdJBUnhUSm8tCAVuOm21DB4b6Ph0TVRNUTcYiKeWf
IC+jlg6z/xMFT7VW9p61oyzhqG9Sl3k8fBczITpvy8Q=
`protect END_PROTECTED
