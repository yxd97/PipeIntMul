`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7hzn9Tc6T1UQHl6opKuHRkU6E44WjNn9v0vRFQ5jf99PjG5XWgpgur0PJpkZpIrN
SCsmlIsPy4QAGdKPZdfANOOzDtEOjZ5Lmiuv4VAnkDoxY/7menPpTbYlKgxnSoD1
bWqCwFMuskZ4GgnWVn4wexkjZ/Yj6Gij/ENuixJMYp2m7RLljwX9U8yW6WPqORAi
95LSp7dr2ulv+8sRc7iQzjn9YfQ9si2O89FsTdC9a91hnSmUn6duiMhc8e1y1KJ7
XQqELUGEpWwjj6lgMDTZIWkUFVGaOF/zcrOrytj5x5M=
`protect END_PROTECTED
