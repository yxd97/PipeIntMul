`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5WSK89jbPKPy2MgqaOeisGLtGiU5YaxE/yjff+kkZglTEyq2w79AlvZmkEoPfP2v
i/FKybbv0gGStp1ukaYJesKhs8sh/AVZ59OetiyaAhIPDxmQP/3VDvVsj/WhEE1H
jKsf6JxvaCBDTe9hf+igjL/JHbtTK2ngtIz2mci8l0GC3Dpj5w+VgNzfuwFhjm2U
zZ+7orctsTSPbAzw/rUmoGzBOFmvnTrsJfIZ/ISiovrIqnlydmVjSOL824iyHZBQ
3OhkeufewLre5chfYUzJhUe+o7eqt4PF10+7H34qrk6KX1r0TPDILlw03Wlos1Fu
SYRpdlh/96ZtnqE13Xn/mWFnBg6z2N080t8e8A9v6o7C9PKAcDTgC6HceJbS6BgD
Mket6qNt6PxQFHzP3W30DL92Ds2SvKF3So+RjYPpZ7+rrol6WLNrVTFFVjWaa4bl
r3YaBEPLIWHmYVXt2nhuozESkGr7oHxRbL4A+ZH4eVFvu+e9B0KR73Iff20oAPfb
+8QpS1XN7LN+XKPkKGphA5vP6cQMgotNy0QQ72qHpTYfyO+O3YlMe1bPSx3rhHeE
FaOZVcqzIDTIy3xViPFPAn/wmU5GQle5KrflPm60abU0GwLOCday/orXsZG4IeHs
RjtHCTVSQ8Pbr55oBjInlIkmLPNoAFT4bbHEEj+OFL3nj40kkojRNi8RWhUmoEap
DsVeWA0v4XqeymnbPkHh2zvuEA16nBl4isWfg+P27NFVYX3IXJiTxTnhXc39FoCU
/r32kBYIXkk6CdIF/IAjc3OWqPJGyRq+I7qhSu1JcRsTFhdgn/KbxAWpDIxNd3SB
UOP7yL9RBqbHt7FePxY/uT90FFqT6UDlAoe+Zcpns4XZgn1CyHy/+lFw313PkcU0
onptz1MUYwyK5jQQk+oSE/VLFTZ6laGuD9+tvWoZibvEb8r2V3ruubcSkmTHAn4p
G5UUC41tu3kLBAXdzimAldf/OWPeqlQ0X/PJCjuyFot8hO4dYhvncXe7QkjmioYD
`protect END_PROTECTED
