`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nM5k1N0sG2Ceyur4udNqqUz4SWY+Di5Ko4dhUT7wcgPrkWK0hhuFPg24k1OLz1fs
rU+3CONtwtRcYCCmGHX9hw8TPaYIegTOJoxATZqRvbM+PLR1u40Wh98gThoyP74d
+T8Q6xigYqDlIb4KSVH7vqBzZ1i4CHXU6hQwzxQw2WZkYB2lVHKCN2/nUAypO2Rq
QSVW8i8IcfVTf1ntMOF2r4+WfaaVGufyzDndEccERGcPoqxyAVsBIrXVUqqZCrWb
CO3FF33BoNwN+2DqwxsU5GVZ4F6kgXZB98vtVPDIAQOfwFqn9sSNB/FEmYL8pxfa
5ULXtwghw4ZvZ0JbLQjzYf0xbM5CR/IXPt1YiSy84TYj9+C0lutETXc79Aed8fyx
WS26Lxj5fs7aWqsEtozotYFC6UQECV5xmlpscxtedRyVIXwjX+ov95pJvovK6Ex0
YVLDUDvP3spcPism/uiSuOLsh1dtGrpAIFl7aXYo5GtWKyBIQnS4hk6HVNgw28k0
Z7KjHck396+gOntNIzOlvN22RVO4Abj8NA9hXczykpQ=
`protect END_PROTECTED
