`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7LIHOPAvw+rpLkf8otDyr0v1UdQfLIeebjfOsbY7I2hqXSv/Bne34pTgpleWTzKC
zdMWl3UyD20CUeAh1Q8CLlgIt1+NX9gT2Y0IUU0IeL7ufGbv8pjJzjkRc4moyzQQ
CXgotN92UONWhhB4/+poiKZ8Waz+G7+wrE0nty+31hzMf2EkrE5DbzMY7mtO3ph4
ZhhrDtZGf3+8gjjgm/a0xGXmjRTdkkeH8TyNIwe1EUkM+nVQRMmVomjuJkSPJJfS
PBZsYcIxB+Vi851SDhft642L5tsZSNEWNke823C90y+STZR0j4kxREz3tc4d0aAj
`protect END_PROTECTED
