`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mFGdukEfKRCTLHNZ5I7HkVgJ1UNYc7cDqtcWloRPUZYX1iTmgMrjm9c3iGkR+Bt
75qMnGZc/jkoRsMWWl88OWTY+lYWPk7YAu1fWVjJ1qyglnGfZeFih2YglrrJfdVu
SHzft87J64FaK98NywkqvsEuuiKknq2zMGnoH+u9mZPv9AkE88CiFrhX/hkdu/wn
fo3cSMwimwSqHuPqcVNaZA==
`protect END_PROTECTED
