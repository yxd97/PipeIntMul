`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
opvpUOn7xKjAhKhhjg49kAp6CtY1BxVrrGo/NiIZACNxSAaUemUQ4RKu7ms3aW6d
/rq+5ZeoY7yYiYU+lxtlZf3WzeSH3Qe4Qp+y9FJnAp3gyssoO9b6i61TBKLCGKAH
xdH3r5TqJKVzQOf0YFVJGiXgFOCfpFIUPFyo07XUw1cRNtmUv3QMlCC0uy9Bb7Ca
o5eqB9+lBKf5gCNjeHWfktSrDM5bOL1S6QENaI6sA7V98myUFv3e1iP9ayZ6yH87
4b4h70nTK4QjYV4p5zpSUUfdjJgzVaObiOatNHCFjRrbogIXht0HT12MKTWDTLvo
9uHYUtZ6lUeV+wly92G/mxHKywYmwwQkOOn/yL5OLxINv+JiG373XXyLTvgzv1Z3
He/oj2AsDy674wpd7cU4v/GAXtCYyoeElbOpxvMv1uI1qbldqSGZFS7HvJjTBz31
zwB0/9zw5No3daRXdLLCaVMyNboL8Zd/WEgPK4z6M8IuryjguysGutXep1Yw0WTC
ubKD5pvx0aCasXV3N8cXS+BR901PSvpl89o8Fl4J9c/zKnqOchF7dOk3A8ekBNB1
MRGEguDlnh0ZYaUQPIJSBQW/OWeYzc4LrEsIsnPkhHw=
`protect END_PROTECTED
