`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d0EGun6KOKhtHpIdUwcFj1YixyQrgvbQSBqljzUMqryJ43ghVRyhwlKkDlW13t4v
y5aY/Vvz4FrpqMZLqzg6iglQ5mfBPCE3Y1O0MrjzBBWLhyytW28I06MfpWVTB4Gx
G+BvZtrfONLXSVCYW/fvmcpMoPam8kizXN1e5k7VFUs995h2SgmNM2Nn5i1eIZHX
5TjweKdsBpB3bRXO9nJnDZXKSFu6gahRrsCnS0s3eYTPUo+C4YKJZRssOYfVmeim
h8EFv1rwTCEYHpInar+7Qg==
`protect END_PROTECTED
