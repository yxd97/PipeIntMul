`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zd7U7T8cZaFt/XfFUHf/2j5bKOhU8GVCsoEd+5NDiOLwVd4PstHAOh97Ni9TS2e8
LvTIVHB8KHpammQ05Rc5ehT1ipYMidv1dmFPgSn7a+SLTVYuHXYhk9AC38huTUsQ
uTLyjrE8xY7go8RcEsSTzzIe8iqHCbV4M9RbE0Nov/c4m+Dy5a29ovPe9Hgpnmqu
z1c96pNituojv++g2C/SZBQZudKX230WYX3z3toZRxKd8fKVad0dkeLw61i5O/Ie
dHeHTqwh/m3sWfWPJIGTWNdioQHTMnmfDUngNfQAxxenkbkREy9gRtGcU4bTba45
ywUmyNYPRa+zoEeyjohsZf+og/6v0n3OqqZTa03KumdAAb/kEkx3AGcrSz/L0E4r
NZpd//hsmIoGtwgj9hfHjV2BFqlQHvg+LVUI6lU1J9pMxCDFqarPrGr36GjorYa6
1++ARRgPQzmNvju5Mc+SlY6WVLdEZ8D2TDVGCMUM3xkpHsxblJpA6IqU4N9VHwwX
nNV8V3SdNtSwI5+TCjMTeA==
`protect END_PROTECTED
