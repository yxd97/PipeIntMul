`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GhdymUj2Epj2q9jDYndHdwi7Q3mVtpnpL8eq2X8+fPerrmoQ/UR4JYjRDWynXikX
FNNj1FKTXxRVCHp5HyuBFialmHAgHTtBmJ9TPLxcQen+1nECcfhnZJpUuzSlEi7B
5fpiMxjgb2wzjGArKJEuh8cwpyLR71K5mFsUj0TgnHCrync2Kkl8il1iZ17PcdeD
HfLFBrfqkTTZO7hA1wIiR0+2G9TMzhoroy8TuziNLMOusVYsrR2FZ/NEHofFuJa1
BjQDbQ0crQfxffps7sDEo6Au0ZeB/EgeB/r8Ff/yP4St3vi3+qB/lIwfSDm0WPsY
1hufrCrf+ervV273r4cRFrwOptH1MtzMk2xEhYyuAJxeYWpgMD1DuDpLFsLuJpvd
KQ5c+EFMgquSZOkv1X5Mzw==
`protect END_PROTECTED
