`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0CipDT6oV6AbfGIPOMdwDWQyr++cL7dN/A9NkvAS/IIBb70npkrOHeIpzXusRHz1
GjjJpThfb3Sglr0RIY5uNA15BRALEWXs9BRaPfzGHfaWLFQJUyweBFQ0giFTSo+0
lMGNtxyh+p+XgsSkDPnwP4TLY7VVhsqG4z9XR9pzsr9e01IXq6Xpax9xonErKG0J
+fAy2hRwmrO4nHTVGPWLoVVoeI45eNU7GC4SQ2NSAlqDd7dQiwO8iy+v4Mj1CrLp
Cqn5eHj/nbU+YHtwO6nMZiKd6rgl+Xh/QG5Qa9zDP+rAasItEfuVIK+AGTf6b7pK
w+74kBEs4+QFqP0hExmDwnblxEhZ0oxWlddXdur1SPHf92unnNghFpe2ynlIJjNp
pHsHAjnaRT9/sFdfS3a9mPIUZ/Z6p2Ja+IAhYl7yZiz/tttmzU76ORR6TPQwpgry
2k3I7+Z62/WlqgaN20J/b4TR5Nl8UJV67pL4RICPT16o2Uso+11EgnE4/Ib1hR7X
Hrm8pxqNSeGB6u4D1Ic+lP4OAQdc1RPyDyQVcySPVza5pXEGtcimRAwL7Y4aMMuY
ST+ulo/UQnJbRUWFqLs/4fAsoayQ9GID8VdT+ZkOUB9XFZDJsprkxDC9GrAIFWQW
Utv68kyDNc7Ex+P+Vu3WLysffZOZK63IaZWoN0aWQ4hlio92ntdyZkX6gUQWqABI
MMNAvy5veUIrPIzH9cwjO7HS3JZBsECII2TBLchBas8hFPev6ZhbvLThRsh5inGp
`protect END_PROTECTED
