`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
etv5d8cm4g2gDhHvZoWSXXr1tmKoXwOFN8GJA/QREu6YZaLHazjbhVuM6QzAZKxQ
9JL+PN3w+kK5StQZnO28W5V8k8nfUlE50++YJhuPyIfLUKYlluvP0qg2hRBIKkiU
Nrw1YxZymFYW5BtIBjpVKY3EvpT5+VNhPIfoI1NaUChQFRyrZ7wAWHWVDEBMRVOk
SQ/TYRlGfKRlbg9wGNoEKSyWTvydlFMneTRjgz66JmQrKef6mw7CNE/+s8cyvYnM
HYtiBpL4vBjcCNDU/mRaps/mMqNVP6xym4ZcZwfQIjb6OoHyMBW1xWD7XpTDyXLc
aXeoAeTpB+HW2DUdJR2N1R161W55y6KbtqtpqckLQyptb19POKNN3AOwzZDvtZqY
EgrsXzY8zqCt75CobxOwvgSuaYDCs1Cl/RavfdvkEF0=
`protect END_PROTECTED
