`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/wzO4F6YtEhsSxx8Rv5q7vpiF+cA8C9yNwciKQXQbJC5c0NpwgKVfLBJeSba2gi
Uhpbrr1T0oVvE5MlpCZTLUgdh4/oRxNMuruug0Kt3TksvTtMTcV0R+9UshD7lAHB
2Oq2mufFyIaSsf9ejTNRDsXoTFlrLoP8IXRq/odMZtosaiqc1dPRgMok8UPYHgGI
buyAtUD0UuGi4kGLnllmlOOD4o3HZy3HqTc18IdZNSORW6pu9QAVZq1CZfY2Fi/P
BQ8n/8izdI+edoLGXoz+Q8EkdmLIqgwy2vk/FW5os91CQ8smVSwjZR5W1t2oqD0u
B/yzFT+oZ442Epl8uwOVmalCk0WJuaGnaaUzyKyel+/pfQAyclwP1TnoGqFYrzF4
AC+i8ivJdj7Wi6fuGKrROYrIqdMMj1lsicngW9tuiOEuXYObzxTddFwqkVaoBnwp
mg+fUfYhqsIJa1WmQmZP8MdBGF8rhXJJjy1FGMoFDBU=
`protect END_PROTECTED
