`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I5s/UqaLlxHYGzg+qgWb8kfpWe+M19kcA34qFSL3i1HNz5+XY8M/kRHq18DT8lbp
1kbKpuk3vLveqWXxjFbZ0zJJOm2TrI3wZqVj2Cj9larQN0Z+WMQHs24VrSexYht9
OvEK2WfZBSNGLStRiTn+HgrSkDVi2yQcuu2REO7VFofcQRjjGPBLK8xG8yUey9YH
CVA33AHzwdwFbAen5DlilhGSGC6vW2rZ3m/zoLLxQzttELZ41dDSyxyUtaO8/PNi
d48s4Q0OhAHvsL5mKd6cAYnsS9N5jU2bBtxR5CDgjz8fHaVXl8b85itYraz+v4Eg
Jvwu/lunfA6YUfMUqx7x/IX3BPSOO4AE5w6YVGRSyywWBplaqP5XCNMtzyQSQmQb
VBbhaplr+xxmXj8YEqFd2Wmc9S4fUzjrbPyabpFmrhCWbHKyBv4XeepiZpgL9vIM
ZK84rYwpfqKCNelcfyiw4K0OrIgBBkUcL/JrpYYsi/JA+v5XiM4B4/Ba9Nnc6x1i
+pnuL9XIdFZF29RSo3Al6SuLssgfGUYziDEEy5ZQ8JhonYdk020AQb9lVotUNiXu
WBGmdwEjpEnWHPp97/7ndf97Nrod+XRlF6z1CfTr0PNTW+EQalijq2juepLE24GM
QjxwFPnVV7kqGgMGPMsvbQ==
`protect END_PROTECTED
