`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxbebfown1Em/sL/P3+9skAaEKD04iinQG+PzlC6yWVRk5MGzrH4sqSU0c/dKjNu
9mz6CqUQgNpFIkdLay6yNsQlLqd52pVG0IVxqpqkjuelIPlw4g2Bn7O7KQq2A+hY
KkQ5Z4f4RJRh9o4PPLPWylbGGjsgYb87TGS12xRhrjKoBf8CHjnCHgWLwGi+kuFY
XUBTSHEnpqf1S9fSPTWqg4Id5EzHH5XXNs0r8m43cONQKa8quige0Xl4yCub8Jeo
4nquJtqAeOeDbDcmwwsIurXqez+IzKfIxtREj2J43WsfaiXX3KgRaZUbiyp8ATi2
PArQDP6hJpYEbLUWQt33rGA7R5alqv9I9JvcNOs897rXhLQhVHcbH57i47B8gkCT
z22qxNUd6j9/7IpTUNWsUU5diui74I8q/Nwx2S1dtkobX6aD4Iq/Yt25qklSkUyL
9AyAO6ALAHPFDskUHIAxo+IjLv11wei3S1vawJAlO8FVY31lhpQ2Pl5vcAuLVPm/
C0wy/CqP4p5RiCsgXQJ8t45tsvMdwojvaidaiT3v9AO+xc83U13dh/Dvajvd6u89
4Mj6FHWv8Xohnlg1sdWVbRKCmLnPshyqUx4LS7LCm+Se/m1fjRHEjihtYwGnMWBE
z5NSVogEvcrrTPzQTLAFsXv8/krsET3XZ/ItmdjgGUPcVFIX9UEO5D/RYYc4Bhtj
978IwJTGeU1TPXu/3MRBKGq+Z3op+aERNjTYEnTLdXHDBPH2v+aKJDziLLOoIkdR
4HdrxdO7rsyed7OH9kbbdta7wSowfhgAnXRryt2MXE0qAj/221O5d/5LL+Kp2QXR
TgdaCi/0sx/t0mmrGDH2nLjsCgvouw+WuNKLhuJrZYCT7CjaiAVnMwm5J951QrUY
2s3H40qbMa4aObsWXsBOIMVOVr2w1nwOgKBHHXXYrhWxDvoxGJvM3FDPmqfQpUsV
qY0lts1t+unm2IVEAFPL8dXZ0jReTwSDWh+0pcqd1NbgWOqMapyO5KZmzDKcoySD
YUkhA+XkeEHBK4M6ZkbOsiQ/VmDqwgdO3DCDJgxlGIo3F0j2Cu0YUYtXCtyp6Y+a
7Ku1q0wYRvmaf3hv88MZ/MI2qCSowC/BrMFQQocYvLoCKyqWW6LfIGY9vdiPi7c0
PNF9TS3lxh+IigER+0/UskB5WC2wLieKCpOUK15eBGQL6/f8CHMpux8Bu57g+bxX
L7mLZOwQKYmgl+8K0AJ0mlKtfk2hJeDegD9GRAVcJ6CVZ/6hC1VB4d589OSsnOsm
2AiLvHb5OSYyP2peoO4p6C+1sWJ9YDtW6DLh30AukjIbF+jA+Qvpzo139BctOnls
e3bYdttRUIA/bKGMzjTLzeplIIg7YGd981IPa2O9Gb6UTYLqas7jIYxLbEXTv1Rx
`protect END_PROTECTED
