`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXNXAOEhmI+pbywpNPSeXPcR42nMpor2hpg4COLmf4odWZrs0v/vQz4l06xSfvaI
QmW4AKKniMkjDkUHG6hZb/UGRaQmHqYmPrBQnf4t3hEoYs81ZxkTrfW3MSFcNt3M
V7YHKTuFy8A1hHPidk3YoJv/Rk9oMfHpS9PrxN0zGfUOQCXzqWMBZendG/4t5wPM
w3ssXUKR8tXFdNdHUvhFyzlbCeW1BXAhN1w+Aox2uSJyU75TPHFlNuwXVeUeLmSO
0oAd07vacFUTeim6rSMOHFKcFSBqwmQ7xnDt0utZUCJwWCCdLdBVyzzQJAZiOt9M
n6nCIhba6+M0ZlY2Q64PwmyGcHzOuW2NmLCVXbURD/y/0rlXhFV+ycp1w5gmKQdm
e0dOJuPPTDJNOXlwoJ3PiwtQrdqbWFD4CABCOvVAmrLnEstYc84lZLHr3wkMTL7P
YqS7M8CgszKQq0tY/+CrtZWaaLhGDbpsUPSAWWh96Ircf76peg+a1dUH8iKcK1Xv
l2WuUXVOMYfHVw6P0EFe0bK58RoGTU+O4VVUlgfEQYGnNagYXMLJv62J36WeGOwO
eKZAW8+X7AM5wdHg1HZJ3b3cHH4tOD0XaDmT811y2o8lrKABkVC1wu8vAKoi+kUE
60bfBNYoM6+2/U5QmSnmkV3lHDueZpOt4lPAcwqhcLUXYkC/UaqLpeFHh+yrtbHd
rpCW6Qul7qZxryv3fhCe8ddyuuMgIfkRE8zuKsAQuCUWfMfemmGLS6UN/UFvA89u
zcRpxxy7RmCQky3D2v/5LqU7jUTQQXxYV3S4GEnlwRJ99mmyuP92FBrzYlYNXKJe
DiJDi0YK+7psHTB2zo3fdw9zSm0ZOMcct1z843Xg0sBSwfHQtlMrTguccBuZsqJI
iAGVi0PIHClK34jT7vFjbcMWYuOH6ZHI5bI0x1NewUALFtWBY9TvfXXPvfRtsNOL
wCCkvxYoWiip76ezX8HD4pzxTT2XbYy6UybbzN/vNtUVsfYbT94jKOtWTUKh9xOS
td7+ThtbJiOsprOKnLYdn5cecrtl38W/RIhQBl7mgRu/i3nT14GlpA+m+H+14FTG
eDgAxtEa15GDNBEFiPDtLCxifg1O9IvojNM66yzk8z+Avq4FSN7WRCuZ7wPB5Ww8
x4b2xL5b0n81XmnZ3TFxJGJFEwAhSkZsUI6H72WF0Vikhh6wnAsHK0r7WzpLw0j4
xfsZPsbRozYBimxeNECUALhxnjKAdNKCyLZmcatnTTb79aj3xA9f9bboNupmGovM
6MVWWrh1czTnDpCnQb2M5483JIz/lIdUbLIHDdnfXuUJN7kTpdfCpy1qSohYURZp
yLy7p9POeDXzl5G7eRfSbJ/jIa5le0/xFY5DU+LC5KFRTws+sQ7TUZsha/EXRGf+
APPKOL/gcxkZhI/pUc/Xw/cnjqB8pa+qJl7PsicClVCaW62US+0zWpS0ZinacRob
DljcmOwCnIOMMx7OuXBJCZMdpfAbzjtCLcjdL6eBYbiAsqkUJmaE3FnXXPvkWG8p
Tm3BpmSkN6oqWB7L8vZNiO6WhDz/Fc4jK8RpCrBmwlJZJ72yrLk0QDNXJBc2FZTe
qDfs3CSZqR3JvDtvvPN+glGRuDntfqu/ZT+2RNqFJKLstpjOEDTA0XSoYhSb5crn
+wwUYp1GhvBdO+4wTCjlXLDrxW8JL3GDRD5/Ces4f1XR2YlOyebfwN86+3pv4+4u
THyW6EhuLo7+YmCIl4wRCWh3cQqCUUBxgCu9EHywe6FKhVKMtbbxrpCp6Pbw4g8s
6rrUwpgyjtiVwWn1EDgCR9lg1bP+ngGa5/gejzZVyaRdL7FXyGBNF7iPWWGX7Jow
ZQ9xVvwhq7wU5a1OAGKq/FKgbFTKmpwFix0+AloQXQQQ+IhxspPZQvVmo8C+lEYJ
KPZ/CaHhj11ZgM9jqbzX+Y0UnjRalYmr3Ho7Wd5rH6RxJ6XaJortKnUML46uGGCH
PmzeKwMN5F07c35k4dIWKUOXS5MoHDxSXTcJBMl9N9IrpPKXWLALNbGmWvXlNhUD
bSkLuaztirXgVNgmsLg13+Sylh/lTn9WNDGazDYCmdI8aSATEl5KJq3YNVI0Y9Gl
HghZtwlJDFWaZL8+I9FZpwVrbj2Xv7PdMPE4TcoZLyEA9+nalUHfjJfto1zQ0mVD
bZs1FVwNw6z17Vdx40Rcshl3ZwVknul0d+lAztWvj8G2KF0lgS+zlxF3N/fxxhtJ
xW47hJexQFM35/XStXe4k0fA3aoHekSHJSSXfjRqHa9XbS8TE6p4yBqAz1kSHG8D
ecTTLUENzBjmvm2nu8FeO2NWcfThLHUN9khv9Vm1HjWk6h8cVakI3SiWCABzTVIE
vU+6ZoAC5E+z6/bSISGhc/KO39drRU36boBBwKrYYWUK5IpFqmSZAxrKev3K9qeH
wrZkw09YtQq0HnhKd6kg3yWadki2oDeLeo3jXEZbdxyAAHIn477Rgv2+F7EoUjQ+
J/PW9/4ZNvO76ytiXr20pg7XMoHAB1yj3C4pJCyqVUQIJNvLBROAFqWGU59VEnvV
Emg6SO35E8ZXoOs838CM+EJnIMtNZal5mD7qssK5lulP9Vz7/m2uQCrH04u2e2M1
cCqY5jPknSCACHkIlBen6anKBArFMLm7D0/rGLt4Hc2Y3D0efLyhAfAjPPXXQsa6
MFcaw+4vNxQIheqSZ0BgIQnxnJhYo31udzFulsTjMZ7Nqubf6MvgSQBXFDq7CAVX
QbcebrQKkHkRxB0bAKINfGH08jKiujjlM9uSlsrPNIMkn9J/KCNyayZUFNl7sA4O
c0dKM6Nxxf7oTFPvFk0H6ZR/OqPg1IySSUCR8Uux78H+Of2ziVbmWgUIClqJJxEo
uwWvS87Qn+gKrWz2iuShwfEAqfLWyiya/1wAcXbOjbCbpX77q614wXOYqWasNEvw
27xd7YH/Op14kVQ1sItKrJb2V6Yf/y2D4/L8NHbViJ2edTEx2vPgTdityNzlGieg
3+WNASbBqXfmF/9i4LxI9Jiyc1pFiqsY0eOFdxIkPKO8b5HnZfJn2zbLZWVzpg+N
pqzcbaVjBiEFURgvD3qDnVeuIzwjhNq86Kw8pVlYsDc=
`protect END_PROTECTED
