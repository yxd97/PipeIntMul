`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4oTdfBZo9NJOTm6D25GaYezeqIrZp0IV+NpzSDXkADRVQcKkRhPuD3gmmEyjLX8
D/qxiW62znY0KkH4vjUj5o0G6X0iHF1iGyYtLwimjIJXxFkAym7ut7BQM8R6n0wg
0FgLmyHFdishrsfyujI8gywpIjDzIFhYJJXlXVmCcUW7nyKc8e/McWON3l+n8Gnx
ERhmI5TDsRQIQENBvjF3VGHeouT8zITrSZ2cwHRnn3xg8S2LDzkEa0AcXqB8BBKj
qTHaRaLdpYYb05tY3DqCfcA8rhNbBwDzmukHloqtbTy1Uk44tMrb2kFK7CAJuYp+
EBjeBu6Xld/o8spe0ixD7WNMtLwQ+I88cs1fW6hEXj1et+5a7FFAQoxa1dfMfFzb
8W89XqsVRFsK3wdI0bDq6Avd63g1rMUWl50oAsSnRXWGj+mdR8H5iWFlqemERPlS
+xktKhX4Evi0YWC3epAC+o/thx5U6vx0Bim3x7KolqXmjcANhL8jmU9pijkIksUM
`protect END_PROTECTED
