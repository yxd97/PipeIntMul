`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olBqgUXRlL3ghSDVeZxwb64TYomzGAg7FbA0GHT3B1Dg8ypAF71cDDZgBL6OI1Fy
sDXs2KPJgX78m9M4BqUmK8twHSp32j04AN76ILRcvqtX1OmGHV5fwg40M8W+2s2q
zmQ5Q4fnW+9UXMGSga8eI0sA4NXyTIT5RZnM/1Eq31tFCJmVnTi3iiCskx9Fw5fV
eM34WZew7BcmEe+xK321vQLIrZBiHw522XqjhR/K6fq1/StKLroaBX9d1/INeYHv
vXRhVvwX/xZI97un0diPqjGU0dJd/5WaMC9ofdVr1dNyxn5anVsimcCAiC+qqAZe
0kYGaeDtFCCO172hmGQ1EZtIEHvTozAuSZtqgO51U66gEsvMAcozy+49w0BBgaay
phuaQDLwsX3cEIyFe0XStdeMfyqbvQWTkQ5XTv3WqF0+Fgcy536i3j4j24zwLgJO
ylGQHDEMEj5FYw2s6J1BXidX+VQvPxs0dKAqUEi41wCmSWyd2Fag44npgikW+meD
Ksrbxtg7q+nskw9SZLgrqbSAt91yJJyFvy1Zk6EZPuXJ7/319Zble4u9Q4dpbz9T
A/ik8mD867Z/ci9CfTUKJfCvH5+5qa25QHOUs+OUebdGSi1XrkA37G4VybwTw24m
OxH/r3bEDtpZCSszbnou5pVmvaniIxvpu+sH2DkqVRw/dWVtTcYjEZ2WNzC/0WIM
aEgYkPcSmbVrqCIBY6fjPBLW8/IQMT7z3h3XzGXQmLFIDLckcoqv4zC0p5m4G4ol
nL45Y6PyHfJSiL0bL6B0k+RMbrmDjdhm6rk4mhCX4k/YYa3iXZQddHhiCovN8v54
RytXSexLltM3TjISMOgZ2KtBh98MKQbNgKkoEA+kULOJWS7K9qNYdABY+GUiatA3
Vz/9MppL51vIRBsMJY7aqo7+0LcZ85zGrCUnicvZXiUCtUD/X/aecHARhD14Q8YC
4xbmhL7Rhbbk6h15pcFL7qCEe1+OjctKWSF7tA1J3uzHv598dLIWcLV5N2ouQBiI
2h+6PXcLXZGTBAfRUwDp/6rwbAxdSaHDxW8SDQtlkivnIgq2GhIePPfVW5CXSjcp
/Qp2Ge/0SiIOx5cc3j0RrnzS+4KLKENlU7d4ko8h+x/5WP5Wh9/qgv6XPzihkNjJ
ljgeHoz065vrEOBDJ0duGZdHsqwWGq2WUG6fQDACuXWHF0XSd5Zk4V3EnrRLOML2
/STsUtfwdDzBo3B0gpa3xSbGpJOIvatGFiDp3YawehyHDVV+KXQEAlqSxqcvAaOX
p9rZxzncKbEmyPa6tnJtJoHTpPOvtKUqonjpry3uQsnT4YSep0SzSaMN++jBCreM
bIIi6Vq3VWF9qx12z6MQtEbRZ+K0c6jHz7lzVtziYZ/yj/9HNFE+ZhlzndFHI672
fSlVusxf8/5uD9xu5DA0cCzPwoHkRkM+br1CYIaJ67fngNoubrO1Pm7169sKzNXd
WjZhdz8mfXpd4gZqIEXeezsIcaDUlV5arpnOvSSjV26geIphEyIUwa5IjEuc8QtC
JQWtuRBzqAgWZlRvWGpHaDDZKaCsr08VE9ePnEsJHIwfRkWmGD8KMtdzvx0fgt4a
+hkYRET2ejMNINhbTs+7UaRgzh4pcpwBEfHVnUZrEcww7sBscFu2B2mE6AbhRpaj
hNHJoAmkoiT8f/Eg+9VfkK+ywgdM7zjr9lRrtc3Yh1cuQ37KsTdJH8n8A4ZSF5zp
evm9cIiRyX/w4MUcV9WkVgZIg04mrRIpnGKlUEPbHQQUUxM0CmiJhlVejJAMjUxK
6mHgiIH/+fa5wzGwjfvKGGvpSsxilcU6naqQ/wmp06lYOZUwaqAceTqYfcS8mJys
HSrzQ/c5J1I/oIXUP8O3Qc7oseO2NZIRB5GnNqU+7tEp1rRY4NeUYpOaHxJ+utmL
`protect END_PROTECTED
