`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHdRGR5g5C+IkzXzVuueFihiwzlt6waEiAEnOdJmMTF2jjsrv2obJSh4xh0TbCR/
2vN9R34tea9Doc9pq6pX3j6fTqzY6iGwPDOAO7Kh0omQ+J5Il3Mz5ixx0oPh2fiU
nXYOSRCPSXOYcbzRBKCGab2r+3G41Xn7Bi36UQsbPXwY5GokqmMiSwqzbCDIVLDU
0P9bPij6U+NGQRXL0eWKQlO1Zuv1E3ge9Aq4lEbCASgEzT4jmUzlEt3a0X9amYG7
jSgu2h8UKIG0K42d14Cp6Ld6o9rQs8enQDRlVSb5BQg=
`protect END_PROTECTED
