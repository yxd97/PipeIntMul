`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCbeXVbwglMjUcLOY4f7xDNvhtKpYI+/RzlfWYQdi8Qu2SuOcnV3sNMFZ3EzcWxB
iyYJKj6iarRoZTfhBWbxpOa27Qs2xGjii8zM73OEwlcam0MBUa2X8qIDYGi7jQE8
/kVaaEDSW7D1JA72NqJ4fJuAmO9l2DyqObRlx3MwQZl9XtAsM0KgG/HJHopguz+o
DMYpqew/K2UfywD9/On0BnL9oB2wajh9WeRtOPi8mHHlp3fApXigcg8lLOuHqKPi
yOA27tQE2J61WdrVG7E9pvOmeLEFlopA6BgBjpRWLCPWRT94BrnHbbaQFdTOIJdW
1yf5E5dgd7TUBFVl3oxYAPmFHM+2/j+v2JZjSJ6n27WMR3OD1s9LSnGRfoyxdAzi
KvfbFpp5AvDPX1DcGGcwW0t0fJ953b7OHc/8pYvVWX8sXNWMggFKY75JUCndkWex
ipsuwVlS2o1c6lrMl3FhLm1Vv70Siy6zWEKCry6NJunDtc6pdSN2a3QrzdOI1qzU
fPBYzgLpn0y4ehMKJ84aO9zEoQE+QSpvRH3H5eETSCFC+fI0Wf2d3mI3e9V4Nwwa
wezlEIZ8wuX42aazziGAGOQwAjpYPTnveJfweTtGws6KdUysN517uAyR4sOR4FVv
30ISa5wno0TUXWX3rmAWvK9/reVVEFoNvAeqCjONISqxRLue5+29vwJnPv/3NI1I
bhdkHDKK+pxv7sQ6BEJEltyv6ne0QtpfATlsrSxgCHPQJsn/ARak/ZBmNN61LWzu
tFjvoCyl/0kOlFmYjkUZeXGiv+Qcuko1zw9IjG3eO5bxnah3PTK97p+Y57t0WHDd
hv9q1K5bZD3O40mGgZK6v+VbCOVrG095n2bKQa3TnhbrxG7lsk5NCZ7hE2IKD9pc
bxp/qek4R8N41MseZ8BeYBjZxuRlxUBSqUXLOg59pYGKjY7nlCd4NoPZ/ikqKyx+
9q+Xu7Op/wq2ziNNHsNw+rUy4OXPpNiFkWcJdnswqQZofA4dnf1Jk1eyjHQmaVul
/LiEnJ0Fm4Zs7adw5pdZrz/HlSbg6sMInVjukhxywUcp3ezPsZFFLPAkDzuoNcMZ
2sVJUamq0msAc8K53pPuzZuXqxw+C7DpCpbivF0gFNqdsMDlbU0892LC6ZkV7kxM
A79NKdk1vztTh9sMZt69Mqx4mqpPesmUa+7KgmpE5KsjX8z9U2zNme/aaB9DhR6b
c4vsN2UuC0dOdl3kTkddi7oUnvLtgsH2oGRY957Y9/bwYYn7zuoEyrg245ITnIWO
x1QFh5AsLkzz1EWa904yLcSMHVX1Lo6sYu1/LlmbkajLxLQFim7SNoglZe6DHZX3
XmucQXYLG7OApWcKngoWRXlt5Y5EKPN1qDAERzg5iDsSk7Agya5titNto4AcxMb0
I7uW6CJnvx1Gqu/2SeBlKBevJDUjMc0MPRUr6OhbHKEBxwv3VGrrvbu4w4RjxhXf
loIeN3aDNao81+WKhTpEoWU9L7MZ6AnZt613jcm2dwzvWpIUOXRa9/+Vpu0bhior
RGPY+J86Hj+xtZkutnpoTBLxnRgd0AaJeMpcPIL9ColJ+An7hu42CXddn98o0w9I
D1YTJQ2mnPF5vO3pmi4lu/+/DgxUc4Em04fL/viJVD1NXxNhoInCWHF5afbA3DFr
kmlJZ5R/VRGPDUgrQAmkkV3J2YIgjqYxjdFMbJcbdSBNKv19N5pg2kHpllktcDFW
HY0z9McUanG7Z0dhsajFp+++0dw/dKSEpJn0rpsNDjKKBYqvReiUtn65GRKrRPmu
ME6thxo9jYFjaR7NOmBpzpe0LCklb6xA8iufkB1n4IgMHmpJWvkR4jXPLJFtAxoE
pxuFAtUfIYb+Pm+msLpCdpM1txK6WbAE+BkfJblkavPlshVqLQwPyDfr712S/5VY
N/mtupxSDl6fglTCcILgT+mssggG30Az316B/5W99rmb2M5I0CWWAjaoFkJYDV9P
Ls43iNbEQAtdboM0zGYXKxVtjPzm7qHECL029oAMU89L9medFmCe+GoFAiJ1YzVf
i0pxKwqc3vE9Pqeh85eZWbncc45poorUzlESqsnpqaQogeYf8rkVhCKMVQEmRCdB
6/pGQt9Nl2KEyXenf3AmH1Zi8gg4uvTAdgi+msDO7/r7ljsHAoMWrNCxL9cyFlxp
aDpJflCZZqsrZB6H4voKb4VnBEsRaUFrhIu3dzwwlC7dBRcfGOCXec6GA4aUOMvO
pF3JXnqirXhTDTn825xbVB3Qzfrq9/tWOMZHaJ1STVhmna40Wf+qkdUl+6wN4Ow6
7mWbMVtKv/Hv2lYnKalyKZavPkrbq3Me0LoZ16D9UDak5NIOz9+RJRpid4sF6Paa
HPxzH38aZhVktLCmPGnv1MpsrbhfAqCTGT0Q1bzgceRccG+t5ztQb+RzoaABzX5N
8w84QfT7kQMecVndkZlj79CAyOcnoCbLLdvdMANU0k//POp7x6wymvcPNju19PDQ
aAzv9yIvNxpPZ9oUcVq4/8V+lrIRB6v46p4B96FUfSUjnA+Zi5SZ1tb8hkuRkQXK
XgS8nhvsENjgi7Z1ryr880swUe91+V5LDd5OisWCrfPxC1vRc4K6sTWtZWFsCHvN
4aFpbcOlcF+B6aqf8Kn0eMc2JiavuL2tEd2HoSNG59s=
`protect END_PROTECTED
