`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXB7tbOx16bUQxuvnA3iKSFrlXJbW8qibPSLgUW4PzoYkjWAUkb+b4o7HzlvFZ9S
/kFj5YPOftU2S04tnD4BQptMog99D0SV0CA4ZShNSJuuDSBcUz5tp65dhBdPg8my
iDnDuU0HO+IMwq80S6Gx6BT85B0fXSPzhTI3Fj/yi6CZPzEMZHNLm1s6Bli1vHYh
G3WbgMfOR2a2jIMCnlO4xb2FWicMCzw4R28vCQE49kVmWOh0YIIDMnkKjxw764U+
uCFqjKI1fj1osqCLVby5zatAtnfEtT8rZu3VLyMllZyaRHmuSPoh6+1fd/oDgnI3
3dHToRO5qgHsp7riu+YPMbWRjnaN8ryIcrrCT1fbCg9v1IwEcPSCFX0bG/HlUjkq
CAKsxUTaJDjxH6BoUAJRNspF3XpObhqQxbnsjJJn2R1sXKdUfJZqESiezR3bFc2c
NMlHc7U5AJdauuPW/KJmEA==
`protect END_PROTECTED
