`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85NSHfwxAN7nZij7hXyfN+xfX3y0m4FEDRjeWEPeEet2boWHWWMX8MW0+HhYmHvB
cUJ03hWS+EzbpDf6mqd6QKacjLVjVdIx5EZIdMk7THWu5JL/t8EtE8UBLVyPYbmX
9DVwZbWCAX+alvRl0eZhRGPXdBRVPti5mgL7qct1bpXrEqgQj3gyaDUEKW00HxG0
mNuNnMCipZZp7JSeCUOcHutZEvqDUM4bOHI/DthshpgGseSzysuWc71Q7+uxAHt1
GiY3vEl1+vtUtQXCdZEXL/kaJ2JSlT1vGgFAd1iQ7RDXRhSJXEtYfn8tujfJvTpT
2PscPYL+2jkjcSdL2qZUY2awighTZdQo7EUhQt948ycGAqPWn+mwTN2Z8nLfgQHW
W6EwWmnFIW+M0NNgdd12s7b4ROzcuCQ0gTI4/PqLhJQqFWTzbk+KewQHRj9Yv8oW
GGHjufFDtb3HqQ162ERW9tl4JQqXQOJMYyuWax2X/5b6KJQA6QbZ2ZxTpai5YR84
BpgilqdfmzGObu+oHIoGiFNn5vRLSsnGRidjbECqBOclniLnJdH+1SaHK7SfLSHR
9Bw2vPVcFKjaa7vAuEgFhCw/SHfX9mgsbcrmRLQnuqf4PHZhBopLu3TefOxq41W6
mUHdawZtaJxsowg8AJfvX/nRtp7s5w+gjjFKHzMfL7Jr8EJXEffek5IAaXIzFuQz
Aa5tcxIRMmae+6tOzkOztN+biKDFAt+C8+1GtfhOni2lVGI/Y+3Ks5Bm2UEFImP4
CKSKhh1VJrFtUPi1Cvc7hlWxAUfIMlBLJbe7w2V6t6K++Eqy6L+3AZwkGiSzEMi6
IDn/76CaDfw7Eyk1bmyD3UJLqKIpN2i7DsWiM/F3HM1bvNbETBfVQdeQG1PPZazU
gDKSIN3s3oWt5/TNkrHbyqnG/PEKp8ljLhiN5S8N1Au95DFTnvsJkruNLIwP6NRu
hMNb5bmcIT93nCc7AFz2s2RhftMBQtD2rswOmpTvml4eAiO2pyaiEn7DHX9ZQXcL
cG4tL3xaLw0Hh/SSykhdpw7xYRODkLgN9VxlP2SHn4U9G7RrruDm1SwAo+XZ6H03
oOcJ/QcRdyqftttH4rF0vA==
`protect END_PROTECTED
