`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hO89fidtB1memMMjaNL7oTnCESH+1irLD+7Skrn3ASH4GtDZdHIpyI9UwWXtUXF
LjJqNmT1TYFehs9/wz2e16mbEIK0os+eAxBAXavUjhuAH2UyOlR+niXbdh0g4hyE
U4VUyfNlt0hXRu3aOqKnqvBoaExXG880IEjug/opVbZmm5ld0tQ2+I0ZR6kJD0/I
PQa4z1Un3W++H3L1EZ3yf3AVoa9F7bPegw/oB85okRbxageAVeTeNNZd4EBkRf+X
MX88ZG8Em1wmWXW3btOUxpjxzyB6fMFHdQ4TendAiSQqOMYQxpSrL0/ANBp5UhIl
39Ru05lzd2ND1jE6iusDmA==
`protect END_PROTECTED
