`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/GY1q69Vu/2LXpQHo+jxMoEnLlegXyaZ//s84dH5pMRSiCshNvQVeJ6GnCmhvOu
LfUT/oW9c457jEb3Jug/Ya+SLz5d2bgjbM8XDrUKc87Lemkd9GMO4+Y2fTYmG08/
VVvUKsO+e32+85ZGU6Cmu1UVivMIs5Fs5adjQ/dGEyoqLMuKbq6u+XMySn1xiEeV
vMssIfitqxp8mdrLm/smndqQk2XeKHqOZRmOcflTuh2VAxTFwunnfOvAE7RVj59X
YzcIzsOxxpspe/UTpeTpsk99Y4OMt0dNgHmgjA/qQ7ghgnwwtAJ2aXWlNe4P4tZh
JO5LF0+/S8+XnBDoz4GynMDf1tUMirnZo8hrrhYh/isQVWsw4rGj870KnonQCuX2
Wr5TGlqIy0mg1coibNcLjgHd26t6s3UB13i2ncXuY3q0/XRCCpNPorX3Q2RrQoDU
UGZ2NDDgRE0rWN18Gho0zl/iMSsJ6hUtD4rdu8XGGrzIz+u785d5K4qZ0FIgKE95
zgnPb/BJbQstbx6OLQf0UiDwHKTA9ftgcY7NyQV+xug4HgB+421QQosIeLyCEbkH
cisXZJ/p21h4hezRkDMaAhIg6dWAAIgCQLEO1pq+axOsc2YEAeeJpqX0lXM5AuTq
6P2yZhC+byXZud2mwUGFsoVb2Tx5rnzAe9JZeWJQ6uCxNjT+7jW8HZ1x1dmPNdHF
jyuv3B7nQoh1lF2E2QoWq3Lw5M+3KVcPknY1dJuhjxfnqZrlDXicTkAAaiMoTfKo
NEI/g4uSiNCc8E8U3jxho4Z8FZM1NX93N34MMaz4kHCt1E4tmC1u4r9CB7Rg8uq6
vqAkJAItR5se5CeBH0rOpptUcu8wkHzESE1Qp01zriimE0ad/8svUA0P/0boEkV2
NEMPrstt6DmiP5E0CkCVkxLUbL8D2lBZgoBy9h+7iS+vtjL7fiRSjSga2T4wXysR
Vx5SuM430qFwBffhtVWi+h6pXZ8i+rIuAgtAtEt3BYSsC83aZhJNIvRwKlhPYQW0
VvIiYHnoHJfpGAiJJbE4cIaZIIhnXwG9DQtI8qCZPuxSTPSs+F/r5/MgaxAwCdnI
fxlqO0cIno+0svHV/IM8ZPNmDGMfPPgmeT9VJRtopvoCFTQCFicjqiS7Y4ncjdPp
O9GieJ4ft4KAo/Bu9Kfw5bTWvOOIfd5bYndk8mhYcEoo1zeDop+7PEfOxwWM8Cu4
J5O3GmVCA4LJOQK2DY1QjKk3J00jNuGYAQcNaUwpWckc4oPJk1LgHowoD872lN8i
LQihcku91+NrOD9GOzxRp0XqXcuia0FzBviAtleJeYfzYVShVGsBJyv5kHTIY/EY
+HJ8IsMUEKtnntmPN+V5YomIS718ejh19HWmOI8WBKZNINu/I+MG8ZChQbMCrvuU
9EB1lPGhjoRzEGSQNvfZ3BwsQ9vVco8jkE19O4vfxQjt8CzW6XYTvHAhdamjKg89
Wzt2O1htl19lAVURTbObLu2PivKm/iI6tptEQrhU8UKzVpkHQO4ADNZ9GEktQ1Kg
KNg4v3XhzBaT//25fPfY2djipjFumswIwgUhfHM5ujKj5uMmkxQNja3w0t4qwd4A
fAGtdbNosyIPR4zHu48CiCxI92PlSOyO4UbIg4is8s39ZgBg3L7N9ezDqlnYAyce
mFrcSER0cqkJKSrjokQhVuEvlc5aQpwhi4j5MHtR2ouJdcH+d2+i3ZGnRj99HITy
DWTV2fetEoX4GuNqh0ta223ONGmoHa6splsbIJ5LQsB1SrkrJ4juH9zKs3n5zqPk
axSTc3IFFBfoYwUXyCjOsXfbx4WVqRSj7UCQG430D5M0MsxfEW8pQTxyKOygR7lV
9+M1m7EvoHUcszYLk17rsj1JIowmWIgZ3gBmoBt6DqioGWINYNtEYjFEstqSyp5o
Qa9DbAP0DGlfM4trhov6BWdZwGl3mFz84ZDnlqZ2D038N0uvERXENCUFcKPflxEj
ugJ1pEnJsxHk5C95f8gyxdIuWoOgLEZ49N9Y0v396EGFhemTRPGXKpCxvDAe0yf/
fpYLmY4tVi+U4p37gKVI6USAfOiQkeGFk28X6BvpLv7FaqJr5r04iW//H0s/sB9N
adaq7wJzQDdy63aj15JosRxcG6fJH7ONGNhEdrw1sNI=
`protect END_PROTECTED
