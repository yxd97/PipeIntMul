`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7B85gdYt/kG40CApTJKplLWEvo+LKSSRWZUn7DWXU6FKylW8VZiGtj+uwK4B94L
wIWEWe31Qc3XQ7qvenEA2lHOB9E1dYpm0Hrz7n/chY1cZO0YFeUcE3sJ5E7zHBeP
sAIUYeXPMKTzk96EnlXl+q9p0m2BLtCpUP16weIdeXCxiQLEHA/9wupXAtyx521h
nw3Rlpbp4gJXOlm6WjSqGI3SdZLOeTmXihzy0EFm6qS7PVdIDb6u9NuCYP1hjW6v
C4/JW3vW6sRY9N4igD3CZGrv9n+xB+HVVK9YXIhxeJbk2TRdAa+ZW0H0ZL5Sm97o
NFPz5zCm2v/6mK7gp/IMwZOBwaD2vmW8ovaC0B1Wg56RJi23qqEKbV9yErDbCidY
YiOqtfw6zoFmPPwK68mFphsRUQIFrBm13B31nkQ0WWdl/7wxrzb7hniY2NuUw2tC
EHmVQwC+Pvi/z/ykXK9xj0uRjY/WOiGh5K9EKtShvQOqibjzJXTMBf+zkaBIl+gf
/mRJGdBgNKO2Aq0p7LRaZ6DbONHmBkDWhTgCW3MpDOnlAxaDrByN19OSoUuyOp1o
bd2tqiV7G6R4O9ISsqPrXD+20gPnwHFUE6m4MGrPLURiVmi0MZZvW4qISrNFu1tx
9VjFULZ8AngCeXh1WOmVtVIbcaUZaNTuUJYUhirTtDs=
`protect END_PROTECTED
