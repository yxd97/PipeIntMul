`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eN8ebDjBYxUxY6pweDQnpyDeQjGgFmAWCmT46cT0F3JIoiRoABwB6RTft6yoo/Cz
RkdNRJmWtQLuYeU0QjC+txMSnq2F8ZJj7fzFjZ1QZvhDAHJw0kK6J5GWP0CqxMyu
HSH/KYcjtKKlPHFWzPnxmHckB0rKKEHLb0Ry+IJioKhM62Vpq8GBMV3UO1t6boR/
wW/rjHOmTmnn9VBEftrSGCnLt1YUDDFYs4xiP2Xb+aTmesP1LfBV8wRpRyXdavVg
8G2oabNx2HeM5D/d/BTGvb43FGe3hJzoFmOXhj47hQnOhBCn71z4wfno+jO2cvLe
Usnk3BtOF8GJ/snsQ5LF6ncKWgJuRjN/Tdox2Yz1MRi/NKdIvACRxGh8W3nqxNj0
awSa2/agifT/+MZXFmoxqc3VVC1cYexXvPiV5DaCU222qxr5fK64uHiBK0FwztvU
z7P3+0+8ggAfpB5r5FtsVx2hcT/UqET3qhuoEwbMif97ExXbqTTgYGYjRYDQWr66
Jx2i7WSS3ZU8U3aRQVOpnWejNMyVQIgLJ2bSliPsmboDq8fvxxfltPQpvXbJbKS+
zBYkam0qn4hYwyhQxa/mqE90WhwJ+m9AfkRV6KHO6wriXU031Xr+YxCrQhZeY4A2
iRYeWxJTTCN9xaG0RkhgRQ==
`protect END_PROTECTED
