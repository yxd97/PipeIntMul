`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mODcLJtola/BrlBoYmne3FUghsPgNXBii8C2/yCzBO+vxiuYPM3W6X45BRDSXKyD
5BQIhoW92Vgcgrn46PcYiJNqc8WzY2+OA6d6h8pdYbaggYexLRlcc0IUlnbXAZV7
Xeso3rDlQ8fuFDmOw91OOusO4RHawPozcPETzbcCkj8E97epkmkc5pPplCiVzFAP
aH8nn9Vk16SE5yIDKLJEHSR5Yr5ioxSSJctHKHw3ngsj4+WN3Ocx9fjkZ0ICFDuM
xCKdl5zDdUP5qXk9SbC240lYWK4hQBWJ8VV2596arGBsbMUGuqps5EHZmeDybygn
oSqKQcjjO7S+JsKKWoKbqGTcw8jcyz96EoGbq/oy9RAx/NK4T3NR3O6P/cweLOHu
bdsDpacjTH5hRHXmk6hqNHysjEo3PbOcR3U3TQ7QrHI1qrShRNT6spvn263Y8GY/
DhTAO7JAwWwHRlrJZ4CtYgCl5+nu0j2UbFA5067xFsXlpudvgrCYy0lgMWCPHvgr
0dfz0qUjUOEKtY5OPqki38LSnU8dW49UUYdogjfotQHxME005/pj+1oaK2w1oEeV
9+hdoUwH1dfuieHUFrzp1pywPiAf7Lrj7yim5bQ38L6Ac6bldhSLtn7jKAytAINg
fg1sPaNA6THHE0XTGaMz+GIMHumHN7V8chA3/V9e1Az0tkl2oPpm9/bQHYZWi4Bw
Bw5x/e8ShEgpluVTtVbyfBOQKRSXRn04olZmTbWQra8RK9bdxltBMuvlipbX87Z3
+V2AMcT2HEfWXubgKbBU/bGCgYKX1MNhAxyqTrBHPeyFUQP6NZgoBa9LHowkQkvD
dM9JI3iHC/yRLiKiQbN/kYRe8ehuEk4dOACcUOEflc53eSayZyIgfLqk/giNgkyA
Rgtfht9DjjdEK9tx1RTjPd21gbVdfr30KDbKa2RENJg9gbJ7n+fAeHiqRjTO8Ghg
0FP1P5t/2nJ8z0LSeI+NmsBHCIKdsFAkyFex/2HBGDdVJXU6r9u+nbRQndHsOVXk
JV6FS9JC2onicGlLdNcNGODxg5zR/YBjs3ZJnopULRp8QbGXaZ5sbcltIYu8b9fp
v80mmoB+hFLqB8M/CwxJnKKl40jLw+cKK0Y95A9u/F/lr4Dz1nepW/DNxjDVknzv
A6PYjYwelzsKSUW6rLl//+ghKPVP3SiBqoJ2C7GkFAIy/GZgEF/Dytjo7qiY80q7
yz33FacGWCTl86NWgppeWv8PI9LAWifZ3Z79F1hIaJKxKfCeQy6ut/hZ8NJ47HUw
RLJtm1t6dOAop96nIog50lvWssRV9uGfvsQOqlfi1SCwOckyJ59p9xCULOkIXr+X
nkQBNVzFdzWJOZ3ynbUI3jOnqegjSqzo9YWEFWGS68Q+rF9qvIAxaWGSPIyUHuyu
f20nTfhQ9v9OPXNoWyL/IdjnhRQ3aeNnTMNCEtaIxRFhIF9gzrWZjQpcK5X/WwhK
Hs2pHAJj8j1fdQ0kUJDknNMjksS5PmRF4Jrr1q+VvEere7ch1k19oBLIA7I0vNI9
F5PoHSQX3aTGXYA2X2iLLW6NhiJQx2OzCbvjA0mGHdXnAMN55VioFisZbh1Xdrlz
kS2vRMBQ460fkCyw+xMvrp9+U63j7Kx5keUJkJdDmayM68B26qhNXBmJkQZr1yh+
fgZfukaoNIACh2Fp7PUBspKJxtL2BXGr8am9kv0P6Pe7k7LSsI6SVC/BF4ij7cWS
ZIXT11eTC8pZWsuFx1mON2ouXm86K2qVTH2F9eQjTiSD3aDzEGHdzqfAK+JawlON
YgqNCS9DpKRb8w5Gtqs5mH2BSAVIRqtAMASTpeQzc4bSuNcUtbTYRjoVzWlU7nMw
t+BEEI2KrkdYoi5odNIPv5UivQC08ysTJSQV65iRghmIemLtcj584D0y0Xm1F/hE
vJ/gwI7KmX1n4W0jFNMjtR5QWoM/Ts1CXkqCI0FrARUzR0wb02ay+VsKckhQZT4q
U8BiBAehdp+uXhiXM9kkOiRS7EvuGR9+E/pscdLO8KSso+9yT9q76wRU9mApNq6I
c0KUU7Rw735ZnbhagpDPlfEY2c3o20wumNp5UojkMQMvjtb+IDZIvAdUK4Xh96KW
KoR6L/KH4uygzZWPj/HeyApFlNMRgzd6wcZO63UGsN0tRA+3YAWSnVMrw4ei91Y/
i88gUyBdzVQwE+T6R7hV29uOUJ/XiufhOWYFS5Z//BFPn34BkKWsYtYFaSRfpFHE
geExCs2QiyD99pT7x5/wGkcnzX+FovEMsuM2EIwp7AP9sgrvEBatGYuQpJjfXsI6
1XrUo/xltN105nTn/qzUxuRUvg3xh+gPC16vvboRglk3I/C6/949+I8c5SyZ7Ijy
cKFNLkp22g1XhMHSJz5x2rwg9AmK2sSf/31rKBlYCJyi7yP+uTDe8O1kuXIT7l0S
1jxwp8WEHFsRQARpaihAyYUJ+tH38cMi/JFpqqMJhDwmMy2awmgLb6QCb9gdvYb8
6DFv1GvQcu+MqqE1nEdMUuNu6h1LyDov7cKuHu/l4WzsmJC2hiTJp6ewIr3G0EqR
ciZmQN/CxojT4bsTM44inq7Lq3Fr8vWIlcytSgBzweMgIy0ClMFI0uqWRJuLCieD
rIfUxFbHgXGP9i9cwHXj301cLzIdN8s7KqAFTxyvSCLUnKGIPbRb6H7b7/AUnq8L
sJpQuhdXtbTQd0k5Rb3Tbn6n1sL4efgilcSm2f8HdSO6fhWaembVzpJudSrZUDyq
q15PcKRBQNSzOyTEEggW1O0S/4Tm9YD8LRYKcUbDmFuabIk/Rd7wRdSak/e8Siyn
je4M4d6eeJoBAyDLaaaAqGaKT+u46l3eq4Pq4w1NRoDsCyXTINixAUzOgSCDXhOL
yGtewvSbAGGdo5c17KfC/Ba0V8iQnfd/ab+YN6fVXvpA0v27hbmeKLtvnZq4Vlj4
4H3bBYeqmeUSCnV9ASxr/rGukVrV4qeI53PyDyz2tF4Mx4KJJ1cH/mIT5BSrRmrs
TswLZn9GIantjIWDdAH3Vk++7dXgOi9WHu6xbXh8QvgjrGG/Hehsv4QAuOTVe216
WQsmnQxzgNjDLpXYp2/gyJmNMz/PurV7JtBbnlnhIL8jiO0NqyyT9dt7AJC8s9cQ
H3uSUW/OJrSPjAypWMiGyOJvhArrmSjuhiNx83ywfedX20bCb/MjpvvMCPat04VY
jClFSEJATlWL9leebT346cIDVgq8WSW1nwMyZ83vUTLJAC6ZeO2pDg5d51j5qlm/
/M2ycZcEipAwci2bvBZ9mXHos/0szJM59/CV+WLNuy3ZKbHC/scmIiV8awb8HrMd
XuMz8bW58E/dYbaWKeAP+vZimFjfibjZ0izWlY4mxA7S8oVyK/LOdzBZgI8Ccii3
CFGTI9TwEYvBvsKsIFVQG/3uv2diQnixJgSVP55kTaWXZuFyK6MLKgrp/qij8KVe
R2+k9sk4JGFNVanqFHP6XJBBdtGv1mB0N0vm3AZyqojV2S+NYhvzqdkLNmw3O52N
0PAbHDtgaWuWXS/UNx0gq+c2X+ISoi3Dq6wOttefkH73xF4WIzLn9j2WjLzVUmXh
9hxb1pF0B+v9b9l5NutwYLQjdd8ay6zTG+oHO0kRgjyjN18mFc/PeX+rlLzKkTbF
pS99LfxW/l4ksuz+iVRliQ==
`protect END_PROTECTED
