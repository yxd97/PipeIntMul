`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZvL8YRnPIZIPdos4X0qTHgWCA4UWKNmgHmWSro8z+I6kKyxbAzJnetzXcp/6/aR
Mi/gQuWtmQMbKd5ATs3jdh9ugsCJ8q/Vhw+SrnT8Fefnd3XzEi/NyHNKIgkan/eh
oJxHaV4SOAFHy70i3r4VlV+X0TAtI8J6lgAJ2F/BuJWkwsOD0I3qKhhGhahD0RCR
Q6meM2o0sl+SjcfZkY/1YlovANFqsO9NVHblBVSln2pBRrTthLh1e458Yz7EDuyo
rcUZ+WeyeQM+saxv2WYTlwHwumReFNVtusgybjgkAnd5S2hm5luGdyNrAjnRxuxk
K2cLo+t6oV5lqql8ZtmPtApO7ZGjF1G8rtBmMEmRmyrN5c1AeV++ukoOPK0X4jh+
PaFqrUdRmxMt5kjJWqUmga6c8LT86cYPcYaZCNxjzaxJpdZ/N2CVPh9tCfgFbbc8
/KTyo5goLbNg9e+YylYSxrOwM2QD9/wxlaWe/rFguNNkeUapddIQf8JTNMdWOgyB
HsXsG+xq2hU5MVN9F+Xuh1CFwN/r5/g3ny3HP4LcRHofb0nIkb/sDyNj4/LxXkLc
7y+f2tY0e6kh8K1S2FDdd5cltbC/3ky0lyDk+brku+l38l+3ro1l+zTGyr6WaxU5
+LgoOJzBDsUJfF3kXF6aAI+hk+K7yX/lKXj24w85RSzNh3yu1VniYTwH7FNSR+1h
4WSv7PAmohy4Fvex/rytEZj/n/aPzE0HO8+nExOOf0Y=
`protect END_PROTECTED
