`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RyIk3+AF6Jg0pZbHavm/711A/zFa8p0C6rfuIki+wQ/4WMMupqeGLwAmFbTOG6JO
XMgNfa3LL6vQi4i8+ATRsjd2M6vXEYuRnTd4pICPbBr5XOLRpmGXOaU8tfo/lupL
cpLXd8JqT8AnWUec+qO/VFpiRlq7riq2cGU1MOe6UXZUIsaG2UohNI3EEoXEcUqt
2WwJRTAJlWy0HXVNK3AwilA8bNfYUw8e3PykqrAXf1KylbKMplybcRJOqDwdiao3
t9WeIVxAQwW+CczxMQaBm6zUVkV+uXrDpsBQFNaVSFfuUb/is02qhP/JAg14H82a
OpzjO2u8MD4qpvLyti5o3e3cNTV2TJZaRA667rC0jZn41X+Ur8F8FE8iVinZCdOV
OLmarohSFqoOeN6pITTLdC07Yzy+6G1UbdHIwkUnJiV1KOzLeEA8RbVawF2txa2x
yTOLM3cuLzneHtCxCiPEDsGRs5QqXhvUcyBXBAUGg1PeKONo3aWw3TiEgZ06DNAL
P19tvKvguQrnzXqY6WffoQ2y+rz5fejVOvyzWA9isPKi9XBT/Jrg9H/bEK1wvzan
+NXTq7LdvZQ/aBqsxog29LnnlyUEblvLHALZQtelgLb/BWHlBXJurIV/AkFwjcOm
ah/rBhpDORb+j+efpwGT/n2kIVe9kY3xq/taBAcCsh8fUThoO+iMb0EYugOFA28N
01ZVYLF9W+XqlBgATGM6ryK1r1pXupHuIp7FN2OElIE=
`protect END_PROTECTED
