`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ieTAsZviKz/Z2XA1B1GLWO7fhp+SPYOCE/t1LXKpQbXNV8Gn8t5CDPv7pf4EqKHp
X3OPmd8et8IiWGAVzsxI6sL0aLDn6Ox8gnqG/obQAwVgQhqipHFP4JG84gD8RgSa
qJYuavWoYc+/RLdio6ycMOM9pNVMlwYlGjOIvNhn5ypMM88U7AHwCBo5axqYpbR4
f8yhQ7AsQizOZWLosOVDlekOcxcrvQvgms9YxvdfkMOr4/I4PRi0OtFx6x0ZeMio
JuzW6W526r5czhzLE6uJCTtoEiG30Yiri8UyaIu3QqZR88AqrYNNUmvPuQKsacDA
ws+q6/uodG7CZpCygugODgI2ZBmx02GTAKZL2jwS9T9O7w1WmNa2xw897ZLrxI0+
CeBoEcT5PO7ASPJeiITTCbEEEYl2PmhRf7ZWvSrAyuPmQbmHJIHpXHaCPZnn80Sc
ixBVOl4a7fho9FhebL7lkfzLGuALEjs/ZU134S800geTI/e8lQ5s6bjJ/7gnQ1Py
LGs182mSHs93xZ53DDCqZA7p/5VK6b/JHKWyKtOGSNgBOfURMw2LlHKw/POC+0S/
+W6DYhESNHKRUc/q5Jjz19sY10mKbrrWf2YFpesx3+QQbB0osJbLCyuTaKrdt3+7
goqtguzHAPNR8j8zuU7LD7sWGbvYS1q5N8EbJg7Xh0tCqPP7MUaaAVyTkzdAd3GP
qGVee48ZRRSVcOLrpISvG+Y2ngD3Urk8eupz+DkkauVbH0fFuUgXx/F1geYlp4DV
v4UzSf0/VjYtVCoAP1ZdO/3RvCzGECxYAUGhz+JG8RCHhVUpBvSLlVsXc8bKWfVT
K6b6iQG6UVMROG1hcJFE4P0eQKDten9LCD3C/PNRYFHQOdnfuW8q2xyQjpU0/UwP
r3YOZykSD3zDouK8ROhcgyBvBki7tgK3ChX+wDs4oDxJK0r6TYeKkZDXIgeAovAH
7BJ+gprwYBBYIPZV4XvGwF5T/cYt1eUnfk/9R6XHUl79Ul4DZ6QCbHAOCr7A9Zn4
UjR4zObI8gJBOmAKjcq+XfU6GSjEnMz7ywIvGGdpDH0H/zHx5eCMMHh6et0HnOh8
FYZ42IvlWalZ8vr7hBLYz4tMBC1+lVjtOaG7eD3SO2zCz/CjFZkbPISvlL18xbqS
Sei/O1RMCVwH6GmgFFwCUJtAokVAqHDYGCRhbTC43jV9Ss+XtsFIgjs2MSATOskH
RQcNO1Np2bWgU2Ud7zxgIXFDuNr1EgXdv1onjJniJcgcthR8GINczokDMmQ86rNY
NvAz1s44fCuzpzanPvm2lePojpXaw0gmtpjHfDIc+qDEdwSM3y+Ub4EGxnWFKSMR
WULczBQ004yVBJSorB7Exzbs0lzh5zGydZNQyIMKOruv7KG+UygmM4ygcJqDpq2M
BvZon0oadWZxENBHLQPTKE1tksAFjnyi5007ROM1glKJ04Q37cvNLDL/FD5aLeyI
+ZxOE+A4prnRywzA7bUobqPPcMSu9w3txCy/klMd9aQ=
`protect END_PROTECTED
