`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwTQQozDj1SV2aLM39DusMcLZi6R72kIV/DLeX/WkL5QlHAyP8gjmwLuAmN6j99H
+guM2bg3Jsxi8hDZR/UmsvvLDDttWLzAanYKvdJCUdpyySBoNjSIUaR36dydNeVP
lsbpyLvZo5G/r8tW2DtkpcwbOPCeNAKt8WFnDNPsxpdoqRch6klm3PFzsCgC8i95
gge0sv0PDgQZUV8e3Jonp4+h1SBOoGWfLt422IMl1r68f2+73Pi77vx16W4RCC07
JqE+sXmbty+9tWbdBzORWTuvn2Jyrij1Cf/gp3ydwk4g8GnnRpaZLgccaoI3Vnpr
yt1qWuzk/6AnKmWKpEuUJPt+rLZ2oDwRUBCb1SzqI8PpEjJordmajZKxKjX/NE60
G90ZRYmdefK1F4uawlIrun0YUe4HMN2IrqKxS/zlZKtKheo9r9YwHJyo//S47UAb
`protect END_PROTECTED
