`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sUhS23YvJslA4zmXWhaMSsS5m8kMtQkyBuaQXBXgzsENii7JGWQ0UgacpeRJBUjp
fQD87jiQjzzjcvzja7/4LkcNBVwylO1j2McigzV2wZ6jdS8+3IyoscCHP58blQst
zKTlL+Ur/yPO/2JT/FRf83MbM3XUlKksYCn7TRw1N3/bFh3j69L2ntb0IebHi1V/
7aDaCqYxwDYbQed6t736Q/Q+uQRBDEID1aMHbDQnTtuFfespceBzEL7qQ4i1jp8n
hG7W2O9FYMFCzhuoR1aRU+gnIe7W/SuXWpS0rrgkNzrEICe6tcVTJIYwIbmq/gf3
lyAo3yoBocqs8KCEfeyvnw==
`protect END_PROTECTED
