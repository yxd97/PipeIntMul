`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2V0jwwaBsxz4r2L1RGmDo+VgZG1sE2qoGPm+R/hK3fF2DrA0M3aQGQIY0iiBn7Wt
GF0jo+mVDhWYamlciLM6n7DJWFP/iCUGCksUagdM/izdWEIuGMBxN+CPWlyT9FV/
XLwf2+j+1eJKKeN8UAAIVYsm4WAaCGNbH0IRZD+BnaXpiPyqw3RX8k1S/uF2riw4
lYO5+Fzr2r2PqhGxFs/MLUiUmJ4e5Kx+5mnDc+3vP3k1AdgI82Ra+HVHow6SjC1T
/YWxBY6iFTlWbq3cqVKOlIpavxP2/zt8S5O9Lds8P68qklLvEaEM6HwHb+C4dwhb
NpWIr9EdTtWAtirBSzKxhX763kCmxYwsOJhLMbqlH0j8nQSlYwAiQD9oLe1Id8X/
0ymgnQd3V3pGvgFGJkPj3zYm12dH+6+pz+i75swS5k70Y8hOOYNRbLnb9FEsjvdp
6kjXp6QkckevZSMUV/sMwlD4PxfxayKocD9OmOZhElgT4bKhSyipNUDjusviHZSr
Ak7naSYPJkCXjpfcW0NHz9RysQRvaJ5Kwuch/JhKXGr+EIb9dwh463Xlkt+hgQtO
64/Iy7DdUdwrO9Dg41RYOx+apMA4+uKC00i4YgKAdLDwwSG9DWi+OYBix80OXJvJ
vyYPH14ltJTREIt5BsHXOzAGuluDyWAZSCoDbjb268dXipip7nTB5B+PELo9o2eA
4CsDcHrbC8wOKkVfoyBcD8PALlhhmV9fqhs83uwayom2H/27M13+8NZOPSeDnm/V
Q5M7i11ZLN2uE0uWozUHykkEc26TB2Uxkfb04RK0A3QB2FF2NU0nUL5Q8/MmKvXn
lqDrSBSQdljQw7oGoj+uXPfexB4DRXHVuT2kkXrK/ZotmeSE3hMj0zKwvyj9G4rR
9aTShJUMQbuRauu95hpmP/Nfz30whbAIWQCXqL2O87lxTg3zI0RU10QD7slBRvAH
RRPE8OW9RsR8Mpo3ArbBRkiFzyE3YmBXg2bAwBu6ih4VTI48b9AAaPh6AMMhBnmk
hqyN8r8yn/A46RTUtJ0qkXS/h8/qsA4EJk2hmC9bNfJqyWLI/4BbYFQIiYV9Fl8T
Mk8DX4Ix7JyUyokzebbDnlg1tLp/gtqCN2hMqD1UnA1USr9GekiJyjprhHHzk19c
3Nqr2jiNHRR1A49WaRylczNuG9QrKtB7YKiYsU6IYVKlLMWqOrhMTUFiV7tuWbsD
txHnH89ySaVWEhFEsYRH3ST1Fpy9e6TpY06HIzmufmY5gaD6AxPpVTokG19nAPPO
oSUUhc0amsbAU9t3PuGEaltCBz0r/DA58JMSCEeR0b/lCrq3oOklUtOhTrqsKKZb
VMN1j4Nb85gZqIYsQehcSgbgIuIYraStpwfjcPi0+S0jdhd5MCqIdHJE3g3gGe7o
pxla7c3UQ8jedhe2xh0ksdN5JJQGEcTEtsHDCcBAb8RfMbQjusV881RqOwOnEBqH
qCOmpLnOQ4zABoSIwBDwTrYbEg/TiB3zVhnpvmXwT89TbEJyHSlW5R2N03VnEFVy
euuWz1lz9dX6phhmobQZWAFkhez1jVHzDk4dMHQ60TSvhLIJ1KA/A9sMlhk0nden
0oNEKuJDGL8CriMHPDw8JsdZGAode/MywMiCn73PTTpjrU8Jjl58rleuQHG3/YDd
2/EoljUdIWhCfcXhByxmJ6tW9TKuOPGAEnvVztbf38liu7twCvNFqrix+SGgLmS1
obVAFe8KHXdrbaUbf/uGqzA7NycZDUzbZSbfw1sbzB+dh8hRipa3pizrjB43Zz9a
xJWPlMPb5xhBwLbPZpKulHftHGbiQf51sjtGMNscFlt4wk82yAgzi+u/aJ54YIur
IL4GfBPTbxo42R+oGlDpvMzMe7vDs8g5geaBXSnnfIfluTSeRdVl94mLgd5S3Y9G
/ft7viBZD4Oly0RzPqWGTNFoDhUgZzKyNSJ9r1L2Jy2mW5/1ajZx+qMlB4k4UCkX
6VQtdcXh1iRA0lFojbHiiGJD8VKw696UTYbUMlS5ajEVHcUOBvqggdO233fXyytC
3AfEz/vudklfkazf418yEiw1V8wDzRvp/zk6lU1mLa3wgQqBVrfGtU3qqxJtSB45
AbqdALH2vLgZIkfHwlUBvZcQPW0Mddm4BNb9sLdwN65c4PTNVFv4JnQTZdtW4EOr
xisNGE9LLXI1N7Qd6KqML2jmJtFIutSRCErKR3rWSiN+0pxRza6tTo1/32xaKZuH
Sn1Ft6VvcoEC14VO33A7M+LGl4K4V0MIUtB6nnu+payTmoYOIXV7baN+nqY5iTLh
FJTIP1HLI7A6imb2ENsER+RO2lorx9nXkPOZfnkHpzB87GGxqAvM81SaBC7GkjgY
yg3d2HZiESlErlPSJeZZystmJXINRtGElKUEeo5nk8E9HPoK6KfkrgJgQf2lcPYX
cFSXGoYBAm1Hd4aXGsgLbfFHFXMsoH/b5Gu148M1t7W8p/2Ba+kvNVtYpXI8rsfH
WH0CNaHERlZ9ETuj+9Aci3jlyJrL3s5zVOBfi34rxLsv3VVREUf7u8TIXv7IBGWI
FfmJHSc1ToXcpj0pYX+0j6ma6RUS/pKEqFU2w2XbdmolQ81d6B1AJeYIhNsS1b7x
epqmz69YLxk1iYsCmMKXU9QTn6WuzfMLz9ikUGKygJ5B2EaCrTA5Gp5WjP71/q5O
Xu3rywgM2bWVdQTgiZvL2j+kBPi3j04r89KuUq301406wJ4UnyF99TgTRW7Zyht6
Pp/VEiK0c2T0GjeeOrf/3Y53np3x9VXmVihi4vz4Jy6kbno44umVYLRHZ5DBCVHa
z2XxasbN6k7+osHybpp6OoWl30TOriehmprLBSvUE7b2jArLN7LeovtpAqyuFj2g
zU1YyW9FeZ3bL5DN8ko+l05UL3qmsqJJBOd3oNSkOFqlkIgsnFBmaHjE2h+dXITz
oy+jADDU+VOsAfYu0vuqmjPa6i7KKG0Vhyv9m/ZqrwSk1VS/N39yAMe+/AP1k/Jh
PxRDBq+2dBPjq1SHYzyLnD/QloFCirjzhIWkNKAQbmG00bgXT6g0folBryPlKZnR
`protect END_PROTECTED
