`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+0WYPcgN1Prdv1QokWR9ySIsRkVSJFFo/RvOsfkDLVbbkbGPVADLvvTmkB7F3PeM
QYw/PLX6S4fFWSjAY+jA5OlSqpWj+ypcMCM8Q9QqrYSHbfjtQOgOQ3qN0069d4Vo
SOXOsEH1VxLwSCPzCh+R4ESyQzW250fakElLXtp2IC2aQHMLR+4y80sPOhCQuVXn
dmF1QtuM2HM8zkNoPfnRhibowP0b6JGEmNekZk++uQ0d2PBt3F4KWjbn5ObDdJM5
5zep3xxbLpqsbkeYggCwrAUHsexrWoyvcTC2e44GaVwOf1VtObY+s3UklOcgMdk1
D7ge94R8JydLCV0JBIXhDDx++KG2q0Os1pcMt5Jm8oyhUEfxXEbVNWnzhWl0QrGz
TLjcG1OpYZ8fyt0BzHm04A5FfX9sAF3/09L5U63h/o8MKpFcsR2+trHs+KF0NHPf
UqOwhHFWnLCIB1qO+r5O5+BPPlcJA9aC8g547VYsHe+bxXot6DUfNCHFgXz9A/us
5KuMBJbx+4p04jJB9c+zrxJ1zHKs1X1KXFWjCDejceAEzd3jWpuPVeRyImbV0+WV
zPMzTO8xbxhy1i4NNLRAzR3rSjkVnTN0vk7HgfqEv/c=
`protect END_PROTECTED
