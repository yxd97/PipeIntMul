`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6d9kLLhOKlsP195dTc4Cd+rMrrb6uJgbys2GpAJmXFMsja7bTKqFfdg3T5JD8rd
TIdWetee2t6ngdOg1t42+CO84USfaCHQu8osJncObXVkn2DTz2XiNZPSEtjcC8Uj
0gIBsjbWBXY2Fa6rLTHfAxZYDcFwmkTZZcqKdd8PESlXlVBviikm81qLeMKBgEIa
dJX24C6FSU1wNsIEzM73NM8H+uo+B/el8VPG/oYG6SEiLg0Yaa/p9TLeoQMJr63s
QZKIGLJuCgb8wO6hYQUlmg==
`protect END_PROTECTED
