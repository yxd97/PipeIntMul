`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MPh8HzXjAC9DV4cYlQvSXaE6TyqXzUTrH7/soxk/UMFt17IoV6ff62I7lEb07C5Z
cLM+J/XSFjzQWjYhFtAx8oTzbwzq5uKsLx6ryr4Wh+G+jwQLz9i6I43C45aa1Ms/
+GULdGs/Cjrq4k3y/XqZYfSs/F0spMc90dIyeAVIHwG3pb7d+ruQrQd36cqe+vq+
plZpi66IIuJdol5ffk/K/dcWRaR3ru1QBJQODS4GTk242SLHHZfMzngmLu7WEJc6
IUHIfcBv3INJdhlPUdBfUt6VBiBxJ3dG4IKmxZniaHZ7SflFhgB0E3OGstdDxsA7
sgi1Da+JsFRPOUYW3JfIiDFruJCOrpT86/kEJGgL4c2EMre0YGi1wUbGCsIlcxfZ
+RLlonhoFi89w2vTNymGajI33o7MKJFTUWtjTldDkdA=
`protect END_PROTECTED
