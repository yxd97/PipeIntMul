`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rWAqaVW/CbG97RY/+w5il7UuWiJHcEpMEpSjvgPly6HhLahXkAd8iGtwgfyuWg4r
K4DdKYa5yQU6gbwex6RBiAadVqWq4eSkJjBtkylq959afvv8ahMRFdXEvKwzogCe
P0f6sHLCL9G8atrw0GscfOWHe4rc1Zta41dG2XPyU6X/wtVnZIcr7jgdS3qvmjF0
erUPFd7Nb/EBrVD+jFhC/Ulr0BRT7p7hAPbm+egxxPxGF1rUdbPBZMkMKjKvRNCe
Qt2ea3FuMpLeWqUX/AlNp3X2JnKxXws4kPEm1J7zP4XmU3806r40BuQYvOyD+ISS
qNrKLj8T07VALHyt5nKK0P5VPKCagbQSXpK7DoHduDvotvt1hAeDzPnq70rVcol4
YrYMvCYD5c8iyHUkVHg6JEAX+YJTRMg8u3lLVsG325AXqmzcOaOYRp3NBlZJqhWt
dMcTHCjS8er31mzw51nNMple9Wdte4umhVCEsd/pKVNEBKW5XU4Xxou2xvP+xIWp
3kVEjsTNvzOPBbhHOQSXb8yKW3ZyCx3kusylvFqXiNW5zUBrFJ6Xe8inYbx1CUl1
jteB4ogeB79y9IiFo7sTED9y8tiYAESlxg19QUlL3atrAMOsA9Hp+qv1syF3VYAQ
CnFTiVPsRwjFQvIpZcX6iu5HzUrZACgglFVsxzVlxPf3Kfq3t+yjrAeVkwIi1F3J
MEnjuNx/hZfJIzG6lgT0ZhByFTzwz+UR37G5g6lPLtpKGj44YYAb5Yg+d6Wz2MJP
gxVQFKEV1I/s0I1M7KmVZ+Tnww71lSkBrfsiOakaY+V1kQiSpD3al9Zmpy9Hic04
BZIiJ9IQ4TczhY93twwN9/NOZs6zMNwTMQybTJGe+03OxGEYDsLA7jNKL24Hxrm2
2xyW7zzLki5VgLCuuAa8yE8qYZxSbybm4nUv+KK8OpG2fKc8oi+ygNP2Ccq9L9T1
bfa7PtxhR2oeJx553gqoRrF0aN/ccBoLwg4N2DjvxIYCLiXcSJ2GSJSTz2LWCId1
SN86edCs6pIjMT4OEdEh0CUUI4JKbS1QnwiP9ZkY0YFw5Ot6pl4WLW1XbcoaMEIC
Bgnw2DZDNOhwMZUYxucPnndBK2vl2DIxjD2bxe76qdQFj8H86IZfeT1pMBVwRe8X
y9pX1XGHQTRF0FQ0BI7M4h2R/Ffz2JX/u864oe1O0nD1tbtZJwkhYmhlDA6Q9Ywd
nUhxW0MLVn/y2EHu/yLZr/xpL8Y0LZZ6jj7gu+NqHsz6tbi2rbDOTCdd8m6ivEcY
bNeANRZaR1OvPEkLmH6PjINz1fWDZ+TOVShrUE0/xyTIyWVox6t1nZIJvsUt4GJf
vdkM386FpbLq35w+1WlEKbkCkOUIMNvvQoNepijkJvPpNtOBFv4RWRnjp3ecAFjI
l9IPpGznJqdGaHfiyNW2U3OZP4Fq84tvo9ioQ/cfWijWXx3qJeO4aGBT1K6P6tL9
xvXPeGD0vOfYSS1iPao6d/EiNVF+TTUvqKuGtY5HX147985pJMezI2B+Tmv+ASSu
F+QdkVfhJxXFsQ/y6ZW5YFZCBAE0JT69p/QgFRmKUzP2gZ4y+DMd6QbsoQcICCKm
yNudVLh1iPxLigs0N53jt1pjZnV6xqJv5+cL0QlP6ZCjnYSV2QlhxByM9LMZY+hr
sujDmjXtqN38Qdg9AC8twG0B0oNRmcoxld9bR/in1C/chv8IwGFlLgYzL9q1i12X
V3++0FoU+USAgwjjs53l7wIjHrxQCb4LvMQrr/OzXsXDXVQS757VtHfsO5EO3x9G
xd97szTTT2olcBYLzWsLtSUAgTXjpqcQbtT7JZD+ZZrI3341Li9sctBN1qc+JhOJ
+oyimd0w+EHSIZVuKEnIAYvZ/TAyOKQhQwkr5K5XnJb+0rLSA9FaHMEX04PJxOnw
es846MvU7vkUQu1PQKJTMZ/O9qGH/el7BIuXuindBCqozwIM0DWqVJMH9dgLYz8g
QWFqUKR6sjYxNnW5mFEOZUPLcr25yQhin6PdQc/Bs66aRJF8bR5m2Km7Eh70PKUs
E+xdyMI9c8nlRT6b9n9daDJIZFgHKfh52IlzEBav360zJ7Ta/WTOoaBs1UlmkvZj
GLs91JN8xfw0bY/S+AKUIiH0bWxlytfMww5g73W0hgx7VIyylGOeemdLspTzGbO6
vqXTtvexLoMYBGITvGUudEFr7k84MyqPDs0Cc7LRYv6saIKZV4rUdYqERhA3k/Yl
AjRdW4RlF9UG+menjQXH2Z+TWwR+chxAaKEIyxwwLUhFqf8B93XQ+OAoGYZUtbkp
rXpsUhZfQCMF0NZ0vKWCoOf7lmz27nHDdzwrPqh6WbXoTK39gkmo5AzRmh9Trvcw
isgRPtUEKzfqJv/Dw5qrnIb4vdLTnZY8Akp5DUhX3lqDjj6Yk2WkaQiExfRkA3hk
sjL8+dh1K8drfXSczroTm5AbkeMHcZQIpVZo3jwZ0R0hUkPx5GDZhN8Xp3DmoJ4F
Fv1YzoUolI3PyWGAGhrsEVzBWAxDdvqi/kTh7gUQgrejxUNZEDLTQrrrO0tEjdnE
75P7rZm/evxu5vMP6BBCdgPmcCTwbbhHUY++hVq5lSGeDEfz6+njLIuPDRm8l/nk
L/1HzIQGRdkB/s3RAsNs+24elZpg5Z/9I/aY4Av1ajElJR17rTpKiVXjcX2rF9+L
CeIOnb6GGFSv0ySQP1CCIYKZ4xb4X2qJiXNR785+6icNSzDQsQbkey2cpL+j8y87
x9FlUjuZZIh6YPr4JpVzHYMfbRfuykQ9Q4HIgKwqU+0Gki0L2mRjouTY7Dan83Xq
r1aiwz6IcOaRW+kWVkk/EnHahKuCLlm69JFld7qJBRFp9shUZz+wOOB6af3iyrNb
CHvCZCAFA0ohcIiuvhsVCjMTjlDAK7pu57kFhBQG1A/1slnuAJHaZHu/5auT/Jff
EIIqLOswdPkEdtorvLHzI+K26iw+ETbxDSWuaMutxRBVONWrFm23T53bGYDFGFtK
KFqIRl7k32gYW9maNWOkfOmdusNjbIojkEQm35u5dm0ehFRIJHC5zeMneHFbyhdv
E8ORvA5cpYkK/JEIlU0aSfOXNtux+fE7j7s5wRyQVattBNuWQeeWh/KpLsGlZSPo
qEDVnRrNRz16+VVJtADrIxEZhORt6JYBfogBAY4uUSR4zOW56ovczFpq/uAqyzkR
JFkv+Lr9JNiuhuuGOMyWKf5hgSTGdDM7HG+IZ1lh+MpLVsH1RcBfI+M0Fry2uH/v
Sj1GuKop/wAhjRjuy8ctkWIF7q4RghlqFfxcpHmXK1dR7wFftUkuazN6+m3jvJ/x
ou69zkL4GqMQjflfWyjtyBgiX0HvYMxqvkFIEDobQOWrLRZeqjxTulCLNawL2kh8
0Ek56/su+IFhpy95+iA5IkD52j0jCd5iZA9h7DxfLbNBDU0maBH3my4/sc1H/40o
BPecXEjMpCh177XO7Oe02nCEv+/EO6eYzBFRnLAjfcTVNy/2MuCcoWbLLqoC26ZI
mulH4IDKxcYP4G/3JHJCBb79Wj08tLMljDlMNBsnci7yYcC/4LBFQhEqlc5UTbc0
dYDNty0gj5APUs7KVMSMWXsX8FTcv2mU7Gb1NuEsEMB1lI/LLCW37TU2bXqtVlp4
3xKAmewcK/2hzVvUZGifYacljBSZUUtmgbQCmchoCcrD0CY16CMPpYRT6vLE0nym
qAirOxy9pkNRXE41uIUX08szYJ5KYb1RbNFfoja6YSywLihPtt5rQpMFYkMYe2Uk
vJj5qYSAcLCpWHhRX+Kc+9ii4wx7k99OtoB9VjmOMr8Sk1FmMeDeYAT1ENftp3YK
s1k+0VUXiy4yxVYTD5KYPp5SzJKROOKO8lVlJgYDvwL1yMfHh0Wq9XUHecTpxnzK
fB6AYls8LCHewvl5scYZ3QryVgaRTeN1FtDiPY7FcYoR3uOurGvzoRXmt1LbBU94
7ZrDvMdHLAYKC+uBnxKes/pkihJLDib5kI5pXpCJ/AZkUEYt54YfeC9s8VgTXZft
WUVEADXXOZrtu0rWlop6jHU56wC6Io+Ka+n12F+31Ell043UENlYgLJZRZcn1eh9
3FRpKf0R1kaYnCb2p7iOn9ZmVZBmWX9Cd83DZJYhYvFQYsUy5CVK/wXg615RKl+K
TB8fiH/SumGM+svCVqO/W6NCKIeRi2K2QQWHVgKqp+EnQ9LGgvXGSEtfWxB4CVX6
lQRLJvt1OIds9m04m/1vz/uCM7ysi/twkTohJM1DstOezHuXK5qGzLmnySA6egpS
65c6yzdyjpJbtxXvGclrJTZmdW5wMBEF+q5AlBCKgit5P9QEc04zEBRHUCG5nmyQ
CYwkkwoEBxlmWKZh8+6ohwd9/b7CFmJWN3P0YB+u1rufz+9MSiKOOqqxsC0cjrcx
0x9E0mM/T3vrtch2KK+TKa5dmquBCoExvZ6VgJr4baAhZ2XGpgWmyM/R6Vaf5vUs
8YSVLXiwHpFLnUKfZhlLAhio6ZEXWmz61b8OY8KMSfuvIZW4qZ4c8CqgmKwheWVR
Jg7aOpyrXWehB5GmEcbsSrA3mPOKwvLQ0KCfH4gufTtHhUmz1M4E2fsxHLK1Y9MC
+WPNvimshNjhPiP1+NjrCvOB6O1cfrNVTayKEU56CKsAHsQZdHPxPw/cSn4GmuX8
9JMvDKTzgsB7XftQxgbNcllVz/dPvV9PC7070oneIVbTzemmdJzwKsdT71LpQt9l
gHiHm3R+FsA4ll+mNI681X6qunSu87cyhso1yQbPIxB7QNFF/+naYEyRwmBVkcBz
jhB/W0RPqpetHVD5XK4/SaUhO1Qs6mx+zJ11QEWCFzL6ecN4ceib2qBioRFF9juJ
gF3LArvXSpM7+ILouz2BON0QVtxAt4XmXVzaSSCHDyhWtGhSrLY8MZujrrRCsrtx
48TilRCn1O/2uC6OEMP9eH8ETFusFEuoLGFNsuvkB0X6qSBnFy70/E5u8QYYOWS+
uzOB294AzAMwQXvs/fvMZ6EZQJAeJxzdvsY4qrh7MJhcDUlS2u3Mig7AJv219oh7
0VWhUKt69WrFhBz6UArji0GNdpeX4fLem07+vqfbkarjs+tUZ5NaR0UE594Zkwi1
NhvSwaQbuFEovTAMiWD+sPuDtwuO5P1WOQgOsPeXANs5xTgza2/rj37WhwcyPaEe
P+wjueq/v94+IpSgxrNa8Jas4VGnEH2UX3zmfTkSPp+JmL5dnMMA81CccjQJ7Fkd
bMerDqC62XyBY0fwB5yXvAsyzO4AzFy0g+lHmBUCWhWz7L2wfxZK1LEda62jQLBp
g3uAU+czg+HbTr1WQMtskbDEs+yI/qiWiNJGrSXFAWVd/X7TK38ElK2G1bMeYAYu
`protect END_PROTECTED
