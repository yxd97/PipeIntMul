`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xdg6hnzVqK+/1Kv8tqvU2+vIH8bPRfD82Lc5IrEj/kZBswKtkipD6nLRhwooebyF
UK9l5C9sqOrrR6ZXKdTH4v1RJumEX1UpAGbmsI0hvsfp603h7pT89JbWpUwOr2ne
Ioqvz2/QlEvKVIo7jnRtnzL/NJZ0q/+wKzC1+YBMTuZvhKLe0j6BtBpUz2Keo/o3
OJMYs4zOx+w9hkmT+2t5zfGTP2izThgQ5lfl3TtVPxERYV81guGq4Y2KU9YuvfGH
hYZdy6YmZzdCXffvcie0mkEoBBcF8jeFse0ayed8j6I2Gcolk+xl4Fcq6M3aQFp2
iJ87Req2Vpu3LtkEMOFkyv+e5YGzZipwInoLFMLZr27bCYsVow1s7Fmu+EYrWmGE
2v5x8nnrhkAU7tBeTbbMUMwF3QXh3vsmQKszLSCnJxBJURDDQby4hUegnjGvx2xT
ntP9hO9jGRyPzoShvJD/0NKgBdznREZ2ZronprY5FPDdLgjT+umgGZ/t8mWwQug3
RBlilQIp25d//rnRziSaygc+aSjacC1yTvmnCXIAB1WWiyFZlUbk6xzsus1fsNpj
uJxMoZGWJsm2lBEPKvhjB/ELpw7pYSsihpBBkg1HzI+LcpuHTdCr9C0tPU/fFSyX
t+t69YSL+L+FxHn6CVM1LjJYMRBRIsekhYGszWu2+Dax3jU6ZD4B6fk23ULgIyBL
CDNwRPG0kC4QcppSDu7z2fEbVhPKwbVNK684NPS4Ii517+QnpCT9j+DVX4uwq+2R
csryjllgKdtdz13KN4kNM9w3TI+eXLfWnVYWg+kbt5PWdoh6UPKuCYYFQioSzyoD
GCyN2DADRNXXlk85w4BXwfhFB4PUTIpj2Dmlwka7u2i5u0/dQZqKskf/BFHcmsAW
zUK07ouEtbIIJemrM/DNqueApre8cT89wSQ6im1vBYh0Fi8+OfIwPlkm24gZt054
pe/fVEKuK6Qs4dJLri4Zw3aupo0biTQxHmB0RTVU4LDNiLpObEW+dnU/i3Hj9x/T
XMiBNksgIBtqVefW+3a8KUHMyBdDgNWWu+n1P9OJZIQxM9lHQS0FU71YDO5r/rZx
N7M7aRwPk9yy3srs9ecP2mXAmybqToRXO39sL0Voo3dEdYIodwLjRsjZztV4TCaJ
LsiL0vVsAxZWvJ2kY5hWwc6rtic9l3+8L9/MZdCp5fMjCeIeANF0gmDJiO73NFNA
yCKsaJmFsUqaYbEq1WD9KN/o5K3jHxREkPznUBGP1jRLidVLoANWClJ/yytYsA9j
rTgTVIpdmnzfLQ4TkxmkutBrPL+vwV1fnwEVeEdY1iK/FC2f7FLGXdRpAR7/gt+O
qUqDjY5oDf1ZcydBpxlGSu0I4n0XmAHbXWKRsEor8svwpAkmyRdZn9llJZsJHCh3
X7UdWAxU1ePQ0zJ7LqIVwqN0nTaTiwgqqmDWiy3927ESU/38Vj2ydQ02fVsb2QsP
N1w/za6lFInLw/fmjc0RQL9a4iRHUJfhSlMweaC+kXRd7ESdJ/LxOJHrbpzrdPS/
rbOdixlubP/M+VDF1uMznt3u7qmfyTA34KgvAAqRq++6tXwe55JS9JhTBHNsTogX
njFgLLTgPdzI4xnyGaDH7nbSDoWbR2uTDf/qBqBP4qBrSrlzdrPEqcr3ulAm+FxG
LAc/dKKBXN+fQ//aMvRuNw/+fahC0fNV+XXqMnorGGq6iJxjWnGcWA+Gr9Fkdjyy
6lxO91XqKp3SKj1rE/7P6Bc7UZtSDNHi/2VLlFRG8KJlh1v/WrWYWQHx54lY2GXs
fA65j7sCaaq7yDczjMFV7tCDc7/yDL8XfNoHQBgXh0CIv3GXWfrD89hAYTLG0d8p
qTlGmHq4X0abTvM65TVzo5WcSHxDrqyobJwvQht1gq/9tLDedJaZpbB9h0Px8opn
Uam89Ki0ifA+QpYXW1tC5U0aDmrpmBlW9h3yHGrQ0a1Iahb1N3GK9KMxTt/+BuDm
++QL1lH/YSlqlvPd8pmmBnCz/y/KVWnlq7xmEU8yxcmTrmpMTq93TtybgWJ5W9Zh
//Bt88Bie/fN0zFXXNiUnM2NYHbDsI0nJSXqclitbf8AT5LqHw0Bdiutcc5Y1Qd1
hqbprD1fEJWBSm2mMrl8uQT/rYNGcxOSkWA9+z/EGbr9nRpBspI+LHsQ1BACBl8V
ABc5vGIetfS6pxfwSXPcZWShv1YPUnSHt8Giccg15rZyd2BgiS4XCRsE1Y9xU7LY
`protect END_PROTECTED
