`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wz21P1G8SCrnM123RWq0jVDQ2xKSpDah9qSROyBj2Prr3ksEHlLajDNtWQgkRBDX
9Olsny+eXnaZONPV260u+Lg8tNxvQA3HrJA0j6bRZMDcRa6Qtnp3WolQHfqOepIn
Svfa2X1ryk2qpzmYhDExNgg2dTofrZp3wa1RR6l6cwjpZa3Ir08zOeKmm7I4c7Tt
X0sJpypEGYBTzhLwa6+z2oFd7/f51yYFH37Aae/5rWntqi5RY9pU0DRYZ6y3e46K
WsXRmDs6SEQPLiRI8HE/nlaNQBm1Hjy0Dgl5ocZ2oIH4YH5D27CChN4QduFNmKLo
d/5CrBO89pOIfpe+HXpkYAn7MkQmmMbRFOGMc6CziQdURiJnT/BxWO027OfsROnG
smQSjnSZpZhKo7mqX3T9arivWn3cqExtAGwL27Niw1ubFmqUX+fETzWzstFS9Ed9
ND54esTgg5G05aUwFkKtTyA5Xkm6iGqxE2iPISFKLSqW/AQunZswMmgU/+wgkDZe
OEY6kjZ5Sr4qyo/fVgKbrnOtVbVaN22KLyr0Yn/VpPU3Ys2pbhYabl6JVmYxQ5tz
ebZtogRToq3CFoj0HhPP6ORyS2whhCKoT2PKlHutfoiBVuwKSatDpPbYuIwdQ7wr
CX02azJJo04hwVDKBzfy0/HatRS4QLLiMJk7GcNBUcc=
`protect END_PROTECTED
