`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBl18IUg8XR6T3w18qxeWBYDzGyzypaxD1rL3av4dSNBcpuY18TME7Ay6eVK9EVN
EdY5NLmct+glIFCp7UfpU9WBsMQI61FuBBBoqg1Dbx0YjABexFTsOW+6/NEk188o
VJ9ljyr+UzYfnf2NfNK2GKIfv19yvX2DWX3FeJ7EY8+XTtZZ25pbYlx6jkTZSzcC
RzQxbC2yYoRHbMcuIqtvmspQJPvRV0Is9yybMVDBqhySXJHwDDB1ZcPAt4tjYaSP
qtm+Qr5JVCFnCmmRkoCzmI30qrtb+6zWlhcOqYUs+3/1WrPpArZc8hzBAe2+khAf
aLZEKXEoGW4QAAUUwrWxgxABpvgywLNdbpnWpuTG8cGDOkHJNMBu1Uefs/WUPCPd
x1QlopRcRKT8HwjReVwCvA==
`protect END_PROTECTED
