`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nfjfsq1yy6vKKjmR3B+QsYyI/Dus8YUZfWBtrpafwDcOXGzU07n576T5T0L0ah88
v34wXhO0f0JFgPh4H0yQhtud7Nu0JIrEm0/bYPu+rOSBrbQt+8EftZBPU4jTjBk4
KnYMAnu7eoPogzflAusD5YVLZlK4/iLkW964drs7l/i7dw3ITrsLzGJzRpApFmuZ
x4PI17STnaO0hi3whGMFNjYzXiz95GyUrTKTwCbB8JROznv+9ZnQqCTMMjxhzWxB
VtmXOSllkFQKbxUse9Hm3X0XRecKrhjpOnBGdSWO2hh8qvAdABWxrtQ9XVYHDoCV
tJRL//AEBPm3YJpZ3i0xWgQPDpK4eRJ6QjlgcWd3VjSGrrPA8oIYsP3BmX+jd1X2
6d5aGI41MgprAx5YGqKkgQooZ1y8kVSXdem2D3Gs5F18QWUXOJVASvNA0AppiC3a
Yi2V4BQ9EoYC07LRrrEWU1vviaiU4/bJJxbteuWW4S0=
`protect END_PROTECTED
