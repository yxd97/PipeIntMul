`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HXLrjqUOSX9zxFkOwePKR2G9lsRpPBwZDqeOZwIH0i6UG0FGCv+TII8mtNSXqRf9
dH5t3DKWU/E+10YC0lzOu3k8MID7uSpSz/5LIyMsnLw37+Pulg/68NIgvEfBxibe
INLSw2M4s2GEKqJ7ygmN93qGwiFPizfmvMbHY/46UAj6iMTHVuc704ygq1iTakbc
BaivPzbPh0fOawcxcv3rwCohKsFzolBGmCMHd2I/HTga72s2J8aJpQCIEsoRuBOY
Lbm5WEdF76kGQON57X4yLN8UFqnqzNLNsuHesMSs5cs38GL7LKpkhsL0u8qgVEEz
Av01RUNBumuDhorWM/7Z122l3DCmB4n24rjQDgduuhj+2ZeuZzpZBD+OcUHshVnp
V32hu7ZLnoeZeOiubSEAxG+MegDfPZgcN/YMoG0OndRE8UaQIiIfbC4/pN7HUrNS
Q4jazglnfaHwKR90TerEGqOplDP4layasslgrDKaa6T6jGMc9MZZhTqgJPiDbSq2
/CIF6otsYldUXMJw40QDkvPtmxxmxcrKoIYhURnTujF43yBpuBS/d6eF8Ug1KzQs
HwhHCCBUkO2FsTQNk9+IEpnouHO2zGlqRGKAkyQs+eOlmnrWz99jYuS1o063upTq
/UOwixcHGTrxA7dWEIWwz6SsX6EZhd7Evy4nDQ5YwKMLOvVz9Ks6jadHIhze6oQ8
SkcDkG3Ah1J5Fe7uACxksfci7NiZWiNkwrz5360uRLrdCi8NuKrVudv78bCVcAF2
OOyGYrBdbyDnpejsxa0VzQNpTRqwiRaO6BXNWRJnmx9lc44fZzQoLoMf9z7OnxNz
byhgMgHMFZTkk1SrHnEBr+jIeVEOfyHEUxVdlClw3hlT5ZNiHy9rc6vdCgLSe1Fh
VhpmdZPYq2MlfdIxvlFN1DR1XFyFgAvGzXUU5pjSq42RwbTaMejrzXYmdrdxhPrD
eK9DJEGSVCPZhj6hlwBIwHm/5cFvFJEYAalklbaVhjtB2OmYnMKxYDWGLMX7Bfre
ouve3vh4R9KBwKm6WgcIRL8+t2siqzrvP0afDi6IKWophBJVxjcKS8GkOKFyaJ2z
7ewBrgS3DMJ/NvaVonIHwlew3HYWRcrLu/Br6RrDD8gskuEQK366fmmhSyDDQDW+
2b+dpUf03tvaZZkGraZEB6PNXLSNZ8N5qblqCHxZLagtpFobTvR/0MLvUF4JPM+v
kNJ/yK8jJO1j7Mvo2ra/DIn3yn8U9V5y1SlITedSGFuwLQLvLDpRyVjah7YItqC7
B/saQ0H5hGTvMH0RcLEe1YUfasujCniUr67g6UIQpNY232PTCZym3vApa7VAUUOM
JIbyOqeiHZUglGqKIIV2TGeJSxg/NK24ini/Bgehr50TniZgawT2dhTHP4KZiCTT
qi8Mw/OBjMa6OC32Kx8c2RQuAJuI8x5UucPY/8jQyLRj9onfQqpj6OMBPYcx/9AA
aG/J8tk22OGWxA8JeEA8EO9xVxpZCbliY+VH0exLdaOAIEq4F4lCryWSK0OR/H0A
3fLWCeklaMXxo/4ILL8ZPjrEABAcDdilXWa+o8KTvCgki7qEC2LAZDRPSMVG7c4x
+45fw7ID02kXGe7r9L6tMHCfkApEjWyZHuL7APTpHGCnYDUYB6bV6n7pFsFTCULg
9LzH1pgWCqaD9rQ3QCxbQL8kqywBl0/n7VbTF5pwQGdxN67bE9j9W89asP0j3yKd
Dsk2nedhogJjVUzKRRU3qNkDYyjQPRuvsckAkXtgsWgiqdp9Ximz8eyop4niRlXL
+I/CDy/KeJBDDjiiYOkzAjOI5/mpBbgfLlTyADZkExmpQpzXOjTg4AiB7qMz3+pu
KSg2XjlcAAlkUwTJg8Hn6u6Qadr6/GyZMp6N15wN3o2g/b7BVK/IxYZSVhQCE99a
wlyw/hIx8WQfQ4vK9LwUV4Kok4VMbaeS3CYJiLfAisu/TcZHXYYpRfWPh7F973/o
HFtbHTj/km0YF1516z/X3s1qFtybE4P5K8/uiGsBtFCfaij78bFEiCaKX8RVN9o8
OombHfp829pe9KY+X7ZATeVWwRv9a48tUMLWHrgnQddNK5Z2AeZvo9r9XVAGrtSh
bKxfYlraFv3IENS/XtBfS+c53kYdQPaHBVKOmiPjzeMHXs4ZPmp6tZrheAkWPoY4
/Hp5iLrCI4gEs7Q8O7uUAkV4xAnHqiirBbD/CMn6TVCrCKYGh5de0WH/DR6mpoBL
hCguAOAMecnmQn3xgEt4r6YDw8mFeDkUHEMlTopiAlsHprJJ7Z98k/1Mx9/bbRj9
7c3NFJmsqzSCQFP9f3W1kQwbjQm8lljJU0VdeEK/OXL0k7oUEXbZcHCxyV7duWeh
9uffX6q9pGNbS4PZrW0/tl4OArIdcgfaWP3jwmd+ebdmCy6RzcJFhnDONRLxbT1S
qpOZ4lHyxFbD6wdksUxnkD4dqGpfobhipKsQC4DBU0iR847PKjTJs99HUtiDDh7f
UpYtE5X49l9FDQh7mfx/r3g144S2c0SlrQuFxu61OwxgB9XXDdrzLvolIvDk5niJ
jTYBtIV+ty4LlHVtQRkxRl4+bQo0BFzFyyaiuTuwu9iP6++TejghAc5S3kwl6Tse
4CCFoDP1X0pxOlOvXobyv42ADMCoXFBr9cWQqIZOXJoxzMUBxWZ7hF0KqdB5OM3Z
THpGwvNy/A+5PRDJoV/FSfQGrgCUSkn9oE4BoGDyE6vTZnC7YIy6+6YnUMWLPlTB
vqLDLeRs+Icdfn/ggy1hXWSZ/cVVGwrvzMXUBWW9IEUPI8X4d6H0rYxefqs3+358
mYK56d0zMaM5LO8pezKyK5g1F1TAHqbIA1onw++tfvku8/Y7HUHvtTQFrTJG/WEo
wbeASPFLC3KhCx+/DPTbJndVsztF+L9DS4bMQpkbf82fk3xFdXonydRs9uAiudeq
9H+D5ZrTfO+et6qvtjmEf8HBcazQ2BIR49pLaPU/3UQOqc1SeCs0sLoAVIsUaDwk
z3eIgM4lAuD8yrE/APrnPOY+TNCgu0EGJ1OZOALKYMW6ujOgh+cHoiLUsEYhYKsl
Th1PefnlM4drcOeybFqGurhmfHeamfs+8WJAQa/OEKXoOkv6vKlsRkGbL4x4BOwY
AdMszOR871ToE875+Swcv1bbsVBF8YB8NIElN+CABJleLxRzBf8MTAJ2wBEdMWzC
Umcy9hq+yzGY3i2Hbi3oegmqKR+D+1JUKp2+cyPgNd/ANxT0Jm5rLArSLShTFmLV
j0N6P4yEOnykH3Zsys7k6joObuwHQ65OH8VJGr7nDiR7+to0yVmduqfDuQX4oGXp
GQYJNOrSURwFOO+gyRiPQEtUCaSSE8gAEMES5JyRmaq7ljwPgANBwAKJ5p7kZw2l
lo25SE5iweB2Xe19WN/mQhBtt0RrSMQnlHWpCbCOF8xaC3d65ArRNkd47wURxEby
Iw+pExisE8gOXEHuXT2pJerrGdVFb/4UCi7CLVduC25QmsCZJDfQ94lmilJvBuNe
ERct5l4vhsHVtxVQ+WZSg05INHR7Jk4obBhegRyxvEfC8SnOz3l1nVdF+dL7gl+n
XTz5pWMFbFXRxumr8SSxGlKz9kVgDC/fsuzUY5120PNEYarg4Q9fq+XEgqdsAsxH
ueiG+rvSukVILY/6avEre/JTAnu2Egin0j4PSPffKNMBz8ZMk+5D70mHxUuiHXvf
vye1CnUlpdSavvmuRBhrq0PSa667jtGLrFrnaRuEoKnIWw3i0hMuDEcEr3e9DS7v
Fx5h27HUlLWZF85/VFfoYOo1IC+ymZmLfwDVc7PrdMWVYaAnRpNsEu8O+ZsoznfH
uAKzYUAkXUhOZqkwxZX23yacqHTHfHGYHHU15KcBuSSR4A75coPYNcYs0wH7DTgg
auH8Z+A4P00p8zozYlA8KPfYuoGw3qzEyPX/J9oyhtGiyrd9va/WYWzjcvRy2MYl
uBprWZkmqMxhocUAU0ShFrAgDSaWQEGMWMXyB0wm+GD20/rsLPMMFOVz6/s+iFLn
jGSjDEa0bTMDPb8JYiK6udfZlyWWwZY0ixPySINZkDnsfTkkTI5mQGmU4ueUu8Va
x6OuBOt6OQmGvPWV515xCygXPnY4ZVJLwv9zPfA7ntou5IrivNO3n2df0wt4OVbN
xpbciYRCeMpO+3tfInF6FV/7WPTE1/XmkP/8WNPSsxA5kfa9/2bAMLubezTQs+Mp
ymDU1XDts469LX/osY0x2bbF1MXHReCeTv2aPP5DZuVn96RPj0jQvJEYjlrohTA1
TiZqBK1yFLW2cx+cGSubeFhpRIKYllLQy8s+6mdxgVacSvCvZ09Se2XrWrShAA34
athO0/9RF0xMcitsJy4SlWUSWvw0cPWVFdi/qWLuAZ+yw0nUBP7SfFjmO4atiFhX
2TrJZwNTT/FSl+ged6BcwZ1Nca2eUnPMfEdSsNfubERqXxahdvWwple2EEDtwsHd
1V60hOVJ40+i2VbM+ypkqVy8ctB60t/IRC/Fp9eTaMTI0gZW4wLnqhc3NBD1u85r
17p7yh7XnM1DFWBpd2R11CoKY0VvveiWbv6isM3tP/ErrCA6dHO5YCXvi9sgZ+31
+vKudU4Iz5AZcH4p7OHmjzsm5zVsyeToctNFIaJZyWrXUCCeAaojt2Ho9zmCnvps
meLm55pmxbUagkhJj3SCNv4Jdqi85f+vvC8jgQnDJSk/9vHGyj6kq4mUOV2xVOOQ
CabH7sQ1ZWYnwqGeSPeK9HGVBc/QDSFouEiNPxdSTX0yk3d2SFBkRPN3WODUrHY6
Wsf+wCgL8Iv1qmM/f01pS3BQJ/E3ijbTgmufG+qXZUiUiZT41J+53qpCDNuBwgJ2
3DDBBQQsN8TK4GvYUHOGYLTWxgFWr5dw3Wc0JdKQpdvGBP6UPl+0H3G245FrK8rJ
y6/IlxLK5L9HB/J92ojZqzJFtAvZOGb1LWIBnEJTFOFxnHf/xn8u4/bhgV4tNVvP
h3LDG+Op7i24s3uV8DTbZ/YqpG4fpcmXr+ZRw+XvnySeWNZzIFg23CVJDCR1PQe6
rR+BuUx78cPiQw2rUJksyg+TfB7ESyKsRFf7ApzOEEQkd6jhwMyI6V+hlobXGB8q
uHtuAbne2MII7EG0baIFpo0h42s8zCt+Mm4chI71JEj1RvQo0cnYLMgzbI/Odea1
WufP8QbG454BgO2jVKdLJVmymoTefaMX5gbe2mB/DizF1cj197AQ0IObb6212vmY
gt0orsvtFzZHACzIhwZEM63klb5JEgUQwwanw2eP6I/WkKnYej7iAVbi4NUZ7CYv
ruVeX144DXNIK2S2/KkTBJGFBtFT0BAn1RhKAzP731s9eKY7kziZ6aCslFEPvfpQ
HT5Trst3nItFAQugGMfiuhokl3v8auSPItPDTNfUWp9zbBiMwBr9/MT/G94lGdf6
s6yzTj1SymhFOIvrRVOuKIVAymydlrcb57i2VsoyTwGHrAh4PH4nFzIdZ1Bv9QH1
E7QvfKFiHixZBPzEyOeOGlKSPWy+i0ee0t2CryBuvHsal/IeMvY01TUsJuqemsDC
UH8k1vgFI78dNbiilujRH/Qtb6pi9WdKe/ffZ8at+Q8vLOt5x1XVrl65yPxG6PN6
VgGc5uX7FsWOUWncOD48jz+IHcZbvC+CmL+gKflx+7fYLiWxi+zRq8j6Y+UpbkVp
oKLqY85OFWm8ZIjKaFxybXJ3WKZu16dH+WUUSI1RkNRfJFvB6dfR33YC4NoTxyxk
r1gQvHZwMybjKs90wtNRgC7n30D7tS+svG9lE8oaY3KYXsuF3q9/L+8eF4Mq89Ic
wRMquJ/CycZOxdKBrTHwAlDZmK0w/LBVkxpEDV1wjzmaKd3Q9WrxaLv/Qr7X8WEE
RIPLweJdO5IF0nrMVmnAdJ157CwQ5kLzQq2XlrOfyIp1yhs3AL51YZgmA9ugoGY7
gvVyhxhZLx8c/shhQx3z4KjrzaJIYT8d5s1eUnafcItdPL98NrYd1DMmTojsr/CF
hsSYM88dxKC+0fQyo3PrTlJOaJ6S4Zqp4I1tGY1Uw49pfks0AhYABZpmatg2AMtc
1dfR4VF2ZrCaKXqPzY9vhFsqFHptjyH+0DE7ABcnKDhl/AtH16hNjirGarXH2v6q
d2/w/R5oPBJ3cHWnFCuFyG8MEASd7IwmYLGdmE0C8samK77dzX6A/TMnteltOyiV
QZ2DtMFZUQOXnK4HeHumiaU5y6VS1c7QLIrrX8EarxB4URCRdsKzr/d4c7aSXf3U
W5kEkivU6a2M2W3lShwxVOxmD01Vn+4quMrIWtCF0IC3DhWXR+vx0+l72gXNILko
+ovze4aMXHZ9PXiyrkhp4Rd07VticEhAUV0PiGRDKZ3kfTNyLSQ7zjbGBjUbu6Ye
47Rvm2u3MKPUowVCw4FAANoLZzEga6nxm7u/MxwqACXCM3oP4MMiiyhgD+aU5NGv
LaOIuv5UgKtVIGYiDSIQ69SYqQJQUyRT5N2CzxyW4iuUf1uPhnrWMTfL0i0OwNb/
KTRMudX2DXZbdWkfaKuV7ZKLBncuV9KJqZjYLN5b/9NaHFEw4rfZiXCVmMJBIK1/
OZVMTZkfM6uWvQNfwt33KD/8Jo4/VWuKMwPJdGOk4OfQE/Xre2LZHZs3vJ4VxKXj
B1h8/2jYKbvnmthx8kXQjOqQVIbOW0fIx+nC5gieOhOF+BJu5tsy3ZzApZDrIy0g
a1a01PQhshzxIwEnnKAVsf55MH+FwydnNArXaCd+EDdoZZjSnaXDAW983RrXpNl+
9gj9ziNeaEKpIieddtvEjc2ivEDJtIIupy95Dih5C7npSGDG6LIfVIiOzzdjSwcC
R4kKBlxbYs0uSFWwIj9WV+eHimKJ4zYN3uyZ397x1L50YgiSszOMtBzuN6atT7yL
HW6YVdzogljYJJuHltlGW4YKOJvoAykt08RK3ni62o252rchwEJWaxdhkSOREiiv
XrnadJNkHXR0XP7kR6TJRZC3fzZZkzwalN3DQcxwh4tp1O7/lbgqG6YgqDhZ7yvf
V2mRxrQMLkhUZv100raB6XcSxOIo17+1rRzfXOoIRoFvZvQUwotQvXA8qRc7enHf
Ry+tUTRxKf18M6YbRn/1DDY2oUpOeNz15J9v0YHmwYYQhXdUEjajsy1wJ4gxLq1h
kFCwXHZcQ6jWTMBGRxu3zzJoc0CeLMumWexv+A7E5MArGldHWooY/3YfPEQsBbr2
PCk23qXtOUbQmedw7EViepZ2Wdq5WA9XSOcvHybv2EN1H2dCJpFqGEoMmwB5+yxO
WzYHXP8GMGWibCcAokoTpFbK1t5g6dLuJ7SDZ6q9xoS0V4mT/GCRo8yQK4oh0uug
Xo8Zodq3BTtyaKa8rpToSq0z0Nt2qCDyCnhYpWOTv8r70FOn7z8CLzvgU7CDJncr
laFV1sEBb+MYITSh5eky6xW2VwdWWr0Oz0GDFhyzPVVC7ohINebYIDUrbx8d2RoK
JAdwQXAoOashrClAGKLxRdtCuYaNaFjp6g5OkjCnjhUkqmOECPY1L15Vcz2QwaE2
sAZVrkugrdKTDfTzSyhNLzEMzKJm1JlAwx4zmCH1eNIXg+CyIk5Qcrtg244Kty3x
1ebPqhF/s1dhbsatfU+jMaKqBuWd0rWea1GsUCP0IvmKInAN3Y5UCaDBlGmSnRj1
6xaIed35xzPh1WYfElY6gbOSv6IhOEwqj9wAWAiaNioSw6i5u8JckLHCTuG0vu8a
13PAlvIkVgUGn+QveSkhsuXnTfsJxWtPO07RKgUafDYthB9WN8F/wDS3B98SHTZQ
6phucszfZXgK0FJhi5Bitr5fzxpSMSCKATfnq7q2F+8zc/t7n8UqcAcYW+au8AI5
EOVgx3l9ibT3wJHSAvEVEOtAcdbPlDZU6Jr6HszqEJLBDZGI3pc1Bs5YdkKwgUkO
K3/plrSl/qfjZMFtsn5T52N4TGe6nLzppYhH5RWDbxidfBYSg6eMFZZEyeFsBQZ2
x40CF9W3FagRU6clonAke6nUr7holcnOzrpiYbwq2KvzisOStIuzZlFAU1Hv31dZ
gPS/vtv+MOq0mtk9le89kTXw0JGSKq2x95COfqThsvbvswBFxlJMd1KX3TVFYefp
behngfCOBcMvr6zGsiujv3ljBH4iH8SrIpJtSmVMpPTilwie6b1PPcr22maj9ZrI
8ZiPJKjEgXU7numr6Yj7be/D0X7TDOKA5IIlH3JQCrhpQuQ5tFDvUB9Qm2MTsMMB
9dEcS9BHA9jW+zKi75+T4Rh0SHSIt0tfY1RP41y6RNC2DXAZBoRylTNOyCSKDjen
kRBLzqaeZ2fDar2gty4gjGQxiisExszyK/pP1dZkbiEHaKiW266jRbOVk9eI6mEn
0gtC+7dA6n+dWRVGMWnU1QkOUPHgk/NAZCB97C2B5+FpcC4WK1L76rOr8QpnSpf6
DJLCFtDxz/fLNgwe4/ENLv1TBlFUy6ij8eYUh0lj78dOarfM89iB2OshPvd4hdOr
IiTCxT1FtNI3d+TZ9HfHJJSFIMseICjJ1f/V7vxwUKWPgeXlg2TWDR3m/d5nho0M
GSQFkZsVAphtPGWIXXgXs3xTO5fw15orXgb+0pIP5TXHolSsz4bUM6NDeAPiiGP4
Yi4DbCDI9iTS7zaEydaxcOow6jiDG0m7UOW0QBR1qwZPGAFlLZuj0qMBzrk5tHAW
nDH58l9fNCxNTvLlLBrSCXc7tU5PPG+3PIkU5UbCqNfbjf6ZA3hJn7P2b2HlwWLv
82lkEwb4DIzjmkHFp0/Gm2BDg1RzDcuEzN8Ngvmw9y0lNPRbHNYvIY7XWJ9pT2oc
+sRrLzyM/EWkZF1ZNBIZVvuTnefaGRdl8UXItmMBL89eUddqvbSFBPbdoPtS9sOY
pTIV+EX7Zg/YnsiZ9Fo36w==
`protect END_PROTECTED
