`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzhqOecVEXJ/FtYDx5ZZIcYoOJLUFBVEcI4j92G2/0GwxCNNNpp6qTH3xYZmlEnA
S/n7rupzpGV364i1EeZndoTC14KosVh7Ll7e/L4LCkS4yy1/9aHMYrp008qsH+ti
JLbiTd27cePLQ+6IxyVtqs1Mfeya5zwsP5vQlE49wGZFjAn5yJ++9y/uPQYqieH1
yNMUdvOEbaup6nGuQxuIHAGjGpnuxGXWovmftX/6/kRfR6KFDBHWocztMw5u2Cir
ui/eE05VziRu21UmLWKj3f9r1zn/QUOrzRI/O88n7H3krJf6dVWPh0n7u2zIqRvq
bCRtAEb4sJUUNaVcAZ5gXhT+kaT13QB5Gp+OFQhbaEY2BwAfRXs0VkUQBHXmVQVP
dklC97M2cc9yuvDStX4Z7F2FbZXBGGP2m/ECBlhx0M54MLKWGrxozgC3bSrJUHZs
i6stRGgfFrrPqowv7UDwktpN/t3EExo51jHkHa6BC9I/Vt4lH+PVUhE9+fWFZpc4
dR07l8PSsplQwLT83oGMMWdAVDEXNE7leXO7gVgCE94tzFCCUD2m/ubfE5VD6xIA
OPruUJGNMBVzF8klnk7F1qzxc1Tc+2z2djzrg0JtjFaVGC3xAoeaeziMt6TzW3BQ
9ffW7gHh922heaDLmNsiJ2D2/Lts87v2+dFiOubJVKBiXnQvyNuvvEoSVWZaCiVS
H9zmWiLrKbxZTiF9j58jq9U4XscYeKFMiPke8MNHWqiarT3kUZoOwI2cJqt51Gpk
Eh1mK2JIHsmX8aBikLdynMbyg7c/Gc/uEtzk48nc+Zc017eiMwkW0aJwg8x2uYIp
m2pTpxNPc19FPAIXv1adbuCRHaL/snVCE/WgxzJYkdnUmxq02yXGjSkwP4ZYStbd
B6oAlaqHaaz0Dzx8a00QfJDG9a4maotOhev6Nld1O5iuPD1x1FjydKpokerlRmbK
SUPaNs1uZpVfezx9qUwFgIHQmu+HDuC/CahbFAap4krkIf0kobh4pD8Vf+mO8shz
4AHPhmE4hLFy7wUDypgnWTE87Qa8cRB/m6rxkf1MJ0j2zYAfTW9YfC2iw6KkplmP
193sVblqh/4qmt6KHklDOBwH4LYStn243RziCJvRzsuDiK4RtW+jjJT/ukobNakP
`protect END_PROTECTED
