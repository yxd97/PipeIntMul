`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GsYUhux/C1R8m8mq4dlmo/okhgsgd7UoVAwum/xv/9jUmS+5MuutXSMpZqm91WxO
fY1gK+UGBItebSDycdmgPDkyosXPiiv6j4pE/QThensOIkbujcq/JkWoF7GPJbv5
i11EU/zLLI0c0ARVlOBnsiP5uxIlACEwFAcmSdZ9LZ7euZnKEFfznJN5u6P0Gd/F
WFUdvl3x1BkxPsxJLJN+c5ELbkqON7x0/WU8TieGmzhlOOCMq8xJZVd+SOUJdVnq
lOWwv6jlTMIkfrcmbpQTqd3puP9QXhw14NFjZBz4oCzZ5jud02bBYXA2gOky4BpI
pkdJR6btV+MjSIdtIGenVQ==
`protect END_PROTECTED
