`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0i1Vjv6vI5mg54fruO+6NDXSdAw0zFleM1tynjLz98+d0P5TVQw3TKw1GgjnTn1
qeEkmRH2/srsuH7KSZsRe5Rr9TVwMDnoaTHqxokV6EkG2oMvzlswXdPu51Web1K6
0TqVvS1QX44Hc4XHI7P0ERR4I/IOGs4T6lrJZ5t1d0yJPDqoX90jMqi1+0DVIn9D
0U80T+FpttJX29uyf1sEwkOLHmQ/JKZo+tzt1arGpnO2OiX6eYr16K6R4NRQwewD
T7EjWuKZ5for9jjS0gWnJ//BdNPs1VvP9QBu/P6q+XrY7RbgWQ6SiXSIVrGHob61
U1xPcqbEJuMLrGvW/76lfyL/iWIQn0o/s117Q2QrpYsnKcYW1k28XnW+5SwZCMM1
`protect END_PROTECTED
