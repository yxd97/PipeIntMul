`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jSty0Lpozr3PUalWqvmmauje1mVl9GcSh4+ZMt5L8gI+mGYLTSuCMbS5fOeFnW6
qpNmKDKS2Z92up+lifRhfyPR/u3/tM8eAGesYpf7f6nuWQ5oKU4K2p9Yh1iZA5MN
SUFBPigyVLCkDRv6FC0KeAWoXn42j+5tGLZP2oxveQHVJUf93QMGti1pKs750K9U
lKOS8ACx50oudjoudNgvLFeeCf3KmW5rf86+KDoAkIJ96QPZ/HJRdEGYqe9v9LlX
nZDGgjsrgWEFf9XcHFUlfmFYn1huJRNAVm9BEci5PCF4GLTU8wIsyDqY7tKp5BE6
0pF2XaYKlAAd5WrBqnnfMxzPiyKFfpxyKhYqF+oV5TTQ5HTOaazl5OF16ST43TRd
FOu2eJGcLHsN26MAl623nQcF+Q4HAC4cn+3ac1jry8ldY4S38slZ10/lGlSHx5fg
rqzNk2AEdeCA36Y0p4MVwk9fkYlYpyyb9LZS5h2RIo6Fr+ynFjI6aFZgF9NcLLUo
0QOVmRv10LXEZtQ72zAdISxC0Fp+KDrQ9Bn48fdzSOAfDsQCa4vQtAN81f83s2YK
uLWxBfM2bTnuKCYGLkOT6CcZgvVzHQnx7eq9nazqEIiI91q2EW3zyBhX2NutwxyZ
aXD60AusF1mKKAjrxkP7suJb7eTZNZMoZ4TOUHfXneYVAckZ1nUbB2qAmiGWxshX
P1nOv18C8Li4eyBHolfd5lbBiva58Gp8aUCKo9G2yBaC2eAqCNfAl3u9779tu4XS
dYFAZ1VlLAIaIQntP5CLuDmQWeIVR5qUWY6hcsRX7js=
`protect END_PROTECTED
