`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y6zIHveQ/Pnh0E/40AzO7osMGISNcG4BUV37oCmYxhwg3JRJ0uryFWlPIP3Rk73d
HijsQixHcjh3PgRXRACMGotSJNsCqGT+L1jItJj4Gdm7LObUieDxwOWa1BfRA541
I0nXWVH7hTxkeB4X6HJo1/TxeVMCYKOAmcUb9BzQHcRUd0A7/0RWNyEZ2tvAfSHz
/ebqgJsDhmjK9WFuVutCzLZJo90ktnd7uy2Co0f3/W5wJi19aDIoPmfy5HAogWdY
u4GeoUZSqCLe8a1xyFv6OO4xXQnTSH9OEBjCNaWtlGnuC+RhDWCfa92LQggWn6yY
BSWLf0Xo4GPcNvAeNEc+kuPtidGrMuyQgmoLChooybRvW5UrXI8HEzNvgKE/xY5X
McWY0TihTKA01GSD8bUFT6AOSzZlrLN0QMpo9zod0h7iIt88AZBnZLeJLQhBgm39
y/X73OVVkvcKMQX8ajzUlwxZAHApT2QjVaxGlrSJ3iMca11g27cdgToINjI90ed/
EwU4ClN8o3/Mv/aAcvsA5F4lW0EyGif4BAp/doeK8KiUnnzfP+KFWj5LWlEEquzU
8udyzuaeiZRT8H0so+esAw==
`protect END_PROTECTED
