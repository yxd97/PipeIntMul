`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9Y/k47wx301uEYaNj5isXaDEjaWMtdre0AE9LclkVktkacHqGt6RM9Zz/SwFw3o
0C1dFI6UIWMAP2KNSFM9qLHv5+w+zsN58w4vvc2EhHccHkg8DN3NQHwj/iica+Vz
houRud4KAc2qgfaFJ+obYa2oKXZGEresUiL0y3RnfPhMIyTM9tphEWZ9BP4aTynr
HDF3qJU2XUqBVjjxvDN0uECijPG+L49fs6MDE/IzzMTKUrzro+rEpnNId6KsLE8p
yqlwuF/LE9amKJ3GEybvAw7psqRUbxS3WrqeLfcIpKCjIaRTgFHEi+s14uamFWtB
ETCdroQP+io2nMAyYVMYPoimiPYWEdJ8o9WBRVERscOYmk7bWJ5nDwJK78F6IIXM
oyqQ2g9vNIiZJfOE/Yvo/A==
`protect END_PROTECTED
