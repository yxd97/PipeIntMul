`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ika+eHg5+8auDCX3dsFiv9fcWnu+TyorrdmFD4za7r9Fpla3g16f0IhMaQrWe01B
y8kYZwXCcPvRP/LnMm6vCnTQSJhpYqKGioXPooow3o9Q2t91kD1pxjbUhZt3EAVH
dpHmagU5f/1oh2OzjaNaZMwuNnzI0Vb8olyyhFHFA4U7tBnsmMeJaSbmC7nIwydb
5fF46KJGyIWc+UCgKA2OXQcnIxS+dpCAZeGppvmingZuAFQtmmHuLtVId27lbSk3
6nhpga5uS5w88pEWsFVAJcE1to7akLT8tNYWHl3jYIdnOxEHCryENZgAKZLYnS98
YEOsi9PPds59zXGrTErkGqRIzoMFQbOmsn+sTbEWC8bq7kITK9xpn+S44q0y9gfw
bg7XG5/Pn6kyEkRt47puiJiTV7nMQpnRZ455fIU6COUGdH9FsgQy2402NdslE55u
d+Q61up2qR0ZeuLUm4zse4IN+eEFwhIJ6bEMRSa1DuAsCqsm6fLHL+8rb+vzB89p
ixM1SsUebqGYBNfZfjfXpyqE4dgmrIdAW3Iuy7YRW2dCudf3ia7iA92ZREJToemD
Wwo0u4CSbbXXGW8NrqMEwC9lFmEy3ehA6SbD+vqWUAs4mRxsyYPLkyABjrxzbSua
C/nLhPSUvPhgSEe65tEPIo9I6k5m48SUyeU+KIPHeMEL4zs+Dm+iNtoDdPPOoeZg
FHScX6bYnmaCACkmBFtWcRBsFHWzBvf/QoQFuA+PWoZVzVs1+ULLGcxGIIJRHgcu
AO1spsGtR1IcjeVJLnhPUGfff1L4LsZ7G61KKm3HmbP6bRacRuBT2zbOIEQnmdmM
rymRAyoOxQP7D7zSVvBFWg6anwGo3Espc2DnV6iSpUC5VsWhvQghIlfbqzZGL8nT
dTjIwuUFrYwXOVHJ3r3i4FLHVpScHDPAOFcfNoSZsimlswXRf/+YlOlZz5d7qJZ1
SCsXBRjwq59VYLUEjwcAKhkGnsEXi1zcKitlOZ7cGElVDoPdHs4+T/ZTb0C+fcKd
z2Er7i147VV3dqvI+SXzE5hzgWRdSnP0TyDleCkurQrnXCg4lX4yAmUkPzMlp0qN
ILv42x+CPG/CnD/uyzkjoAfeXTLGQqLD+IkhH44q02/cnv6WAk87B+qffKf5bWZI
T6yMSM4RqoOUO6WvVA/aX/Wu+SeZfwA5+P6ZdC2eipqnCK7259EyLnquIwJdeU4K
XWp4E4TSLLJQrBa3avX2p78CCKzNPpTcILOOMN9Wze5WlVtLR34OMJJ0MWU7ZIMg
7lGAmaWj8pSPY3fwxTOISy4/EOYRpu82hmyDeLzYp+MDs3JZYyPfLKFvhy6jV3Wf
1MZSwU3HWg6eXFjGujEqCs4XIuSsSCQZ0X4ETUUmQbsNItk/m+3C6udBu55N+BjA
l+ULXp2nENVF+QnGOdE9X7ETKqqJRiM9GxmNEdBG6tihZf1numCt1kp67zQGwcyb
xaO7lBiV15El2vtZxRV2xZWaD6OYDeI8/EcINurgvzT6yoH4r8wdrCrq2Se+HXJe
22I45LgFx9NWpIiO3QXrhUNwDL4UcERhNdpRXbAx5oX6ZumiIs0Oj3yFBab7m5Ui
XPY5DiSj+GRX58aF4uiNRPilzWDNuaVn5cpjmRRDq6Qlv6FS7Dt9ZwMtL7Gu8HVo
RZgVJXCWNtdMVNj105bjExZxe6qQ4lNWT9oAZjN708gnoeeIgL3bxlgna4kNAGFk
BqSGRLzr4D0fv2phPZyZix2+4eKSsZdHCHSDUDxdov5hL5juyT+q7SvPNrYBy4MT
e0lq9MsdZwtGqN6qMTOI4rzMSwsLTCss9cwIrJGg9cngZWOTU8M3pFspseZeKYln
7nlfLsmNSmso/nB/q30xb0B5suhaVaZzY0NIUwF9kitmpMJU3YoQzaVJuNdD8hf1
TD7LOh+KoKEOsiYCWLsOG/JpVc/NKNv5F/sV3EIWzp8ryk9b6LZerj8RGRpiy9XK
waHfVXLmXV38JL9yne2F5u4O+GXTF36scO+fM1PZeRVJBOTCNYNOKP5oTEbbbbRM
fRiae8j/MRz8IdRbcmRMCYjov+4igG+dQGyjWc2tkBUfTbSTOKEYXMQet5wu2Wv6
7v/vzGGmv6dn3okPEGZTTr95RFQBzBgmFEOogYX7AJJXbREsT6SojFRMTM350QZo
U/7adHbjgEIuNEX3PkatDpeTZPqCBCxc3l7gv5rNtMa1ZYgWMK5skwjKhBSCr1PG
y0emvaG78bOt8AcTAnmsDD+IdayfDDlukMwXoyaOzsJz6SKhYbdh0mC18goxjgdq
0Eoag3xiAyo7hMd7TquNdH4BoZYVZe+2u3S9+xas9fI9e+zyQxCKxpC5+93NDL4O
SC2eUCzJ5o2TXVXpdHEvNizLIfB/Iq/NVDIKjZYNKPcuY4UGVZxzz7Hf7wI+Uktj
nGF0U9P49TQZ+qdr/fMeGktYmtDahmk0L9OsS5p/SiFYSZ+YneUP9vaTNnJr8979
hRvNg9SW293jLzW0d0xA5t6HBJE3/e9+EaZeCnJWQyBHUwiQBnHH6gXBLK1G7B8N
ZiDL9tG3XS1802ZAFDO9J7b1jDovsYmPaVnEBkv0wcPSdLHv++QCBgl5U+JUm+cE
4B68POwLmOJ6NGSDW6BKC5cWiknCz3fwYb8zt2IKJrnK5Br75vQtWblAkHWvXF85
jIB22ftIEvER9q9uS79wIs5fRsAQYQ9WnCS22oemCL17uM/9dp3VcS4Euo9VudSg
NeRwBOn8JtkbwziBh8m4PCh+kZNhRgz0E5P8oOWGAHrtHHtq9W8b71XDtjeMRxI/
u5gvNz7ZsWXoPNuU5q/e7P64KQ4lhSAd+UbdSZYvQi1klZtUOYZeKhU7YQqE3TPz
7OnjDsAm/adUeZGMdxsiIbDBqFA2msn6MbETvJXi5Xyl/t2ng8EKKSDPW8Vburgx
ntJ8oqBnUfGzqbhzO42EDXCIXW/SZ9wXxlQNJGOEcEIbOGBgJVyCFdFcMaDP64SW
PtLiQQ8W1HE3jvQM2TZa8J4wc8Es6yFGJ5xhRZ2a5ofLH3uWzyy2vMqDkNrP6LyO
hGwWwDPzbwumQsmpWudQVVZBrmwqrImFQhns8TOUHwlvL1FsHj53hMtXI63lX2eR
6hV3kQN/YZVMb5oSJa2K/5XNWMl3BK4otllENEkGWtxaZZ0y66y0jOmdj1fN+gIf
o0bVWMaJ6quW+LYEmRQEhXI8Dvvn2sMc3/jBPPh6kEi+wCqmlp5lT/4+2l898WWD
OTkWWQTsXxJAovdjxj5VD1Jb8CsXszKeyizg/Q84k85dMaZZZ/Ei0s36yWfDoLnu
vQQEtZhFZynik8l5jhZHGhouva/ryMCy5nZhnx6azhGNfNcVfoxlhhqRwpVv4E0I
YQF7G2WpN3RxK3CgAvgTX7hav1RiXlT0y52pDN0wYGPe8SyeivQajgKQpJ4yegTg
Dt6VT8YMmfx3bV6nMShsWtmh/XpXZ2z7WZRPhlocJvqdjBHqROk4ybGx2Q6S3mQP
cTVZ51J66vX+7xR4i4DU0Vby71ip3xTA781Nz+anGbKsLabxy7Y//ZU3KGm/TZTX
yEWyHxn7yhmoJF6rF1ba9Q==
`protect END_PROTECTED
