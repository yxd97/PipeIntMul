`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0R+92o9qbEl92AyWtPw2F6wiAKu9AfA0dgC5cTvkA1RiT4fegMz443B5vwo3wL80
2FjOXh4stzBys6psI21myxXHMYmCAy+seqrKesINCU7RfCn7xzi5pyWaqWc7c07K
rUnwLK/DAiRxQxnz6EkO76gBsiOibGZlWvIubB/t6RK2CiwxNVdy+M5oh04kxXcP
MkKnrON+MMA0F3/sFZUEuWJtSAEPGU6gOmMeT2tbtsZ1z/nA73+P845B777oQXnA
fdMnKW392norcJ59BOV+dRa+sEM2gtspxCX05DDYD9oZkq+7iqpgYuq2/8Osth3P
GZozGv0b2jY9dRCC/jh5qpDYwWELJ1Own41SbMZ8/exPrkz/s7TSXGqqQpeaHt78
ZUF4IBKGosRo59nbb5MVMw02eV8nkC3MqDIu/1OJAsX3Sk13CQWhmzLS5zE3R1Fw
/Z1FJALL6dwSFujKxHFSdQ7JblGROfJqkvFX7XF2SIbcXTMDGaIIVYngPEFcze/1
`protect END_PROTECTED
