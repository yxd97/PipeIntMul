`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKroQ+QAR5nYKUqQ5Lc17ZnxYPZOf6cu24YT05iObemlX9zirPboT6yj9PedCl6j
krDD4hWe9uHjUrLLk+MkjX6/goz4/Qv+pGBZHZdO8eSY7/0fsPwv9paM8KjfOCiv
iXEqjh/8bmCIIvg0GJGM4MG4LW0V4qsZ0bivXHfYujzjPrRpzTG76hXSjFxRyEZU
qT+EB1B3erZfIMy859eZmPijLfBtQXqzZ8O6zGt3vc1fh4ebXoXxSrZA8YNOF4HE
SDTPTkrI1qtY5tKbrllFf3+i+fzbstRvlRHcD26ULl/IhxngWwEp3i2jFyLz6Atx
r7odZBHc27oNFyGnLXOqxj1ZA1e7TFbNOrNii4YFqnPN/KxDu4fleyElnD+8zou4
THT9Xnauu7C71Q9luOl16lxPSsENo3xX11Ctp5N7LH+Lc+S7okn0GJQZmHdw2jsR
wwWWNLbNw6vB9eqdxVbfRSy3xYye7Pu9tp232RV3yXQ8ttahnNcE6HGyHCSubReN
kN6FYJNHq6pGJMD3E9UrGSJzwEsDr0eQqMDlF+CXVWyeN687Cs9aBdFIsU34uK9r
doycJk6kfKV71wC1+f9Xy1tM9bI5pYZvzN3DIz8/Puon1LU4jzD3EYi19m6s6fUI
`protect END_PROTECTED
