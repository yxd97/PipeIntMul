`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YIjCYuo+BX9Bdlf+W1fcF+QizicyCu4YxdcD5N/GYmfkm0GW/28P3b83UViLVjCV
mRtDzmHIWxvQDy2t45n3Fl8/6wToRhfqkJaNxhv3u7nygH1N/kHrfW0+wnnjvwGr
7f9gWHrhr3FObmaDGOKz4nWZeljXzLHZ14V+OqIMmwbMFFGCWL9IOE/Pol5KdTxt
a34R3Dz7ePtk2SwDh6GxmD1l6uVyupfiHf96Y8ZaElxrnzLrzoK9N3VkpOSy6Qz1
ZZrjcWc84nWnYB4iYZDMCKUlATap/jGmhv2w8FPfpILqu9dSGimyyzg8UOO2LCsz
rnL3G3z08vCv7PGhRMbhM/LaIK6wJfotEi7cHw9osgJjQ1MraTHoGuHXovwhxJwT
VsgfmiopUTfbuUF52LmdyQoaiPsIfQBhJYu8sC3NPXUN0s06knzHn8/UfrFlKWKR
`protect END_PROTECTED
