`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RsFlaFZwTYTKEnSXyY/DiWxycXXl7xUSv33lcrSep59R/2Tk71pn6IdxHBeLSY2P
SQnZiSU6ggp5o8hB/7jDe/YhDW07TOPov4px0CWGAem+m7nxI0Ah0qglRi7X6ZBY
7AmSuS+HONJSUS79ZOpOF/aiyWYdSeXmvPRplLSMjE5Ucwevm69WOzkmUgMzE7MY
Kc3h0+G9vM7mH0nS+S9KQFdVeBBtFifM+Po2eHo3NjVb7kYRVsI4UDfbE8dITuec
nBM/BpLIYgq/QPuTf4dNyA==
`protect END_PROTECTED
