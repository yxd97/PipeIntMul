`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FoKGNDpL8XdPJoY/RSbqpCUh8xiKZT2r3puobBk6Si6J22dqhu/sILAIroNWTDDU
zINIO3t/1l5gpJtLLbJNI7qY3RpUhCoW705LbUKbFq2u+ShIF/BH4yNsDaoWhCgD
OwqAka0rx8Vs4fksZovOfynwhrQhgDxF7RZ8EK42IsmX9Ni0oUrI66B5zMnzeRi/
0PcQAGujXmZNKWj2zOEBr4YWfiB0/y8y3i8AvJGaPgg3ve5lywzbZTI8wuvn8JlR
laxVsyoZSEnEG0ulTeQsTC2+mAaINK2IMtJi2G3yt99xOad93R4/vzLV4se2z5Re
xAu3hl0dlyBe4Km6mzGQvoR9H1/Jvq/dp0vVi5nKbql7bJnpaylY1/BuxFn96IPB
tK+b3My6JqjrWi+zMGySZQ+4hR0hiQTCkxGcP+Zgm5Q5WFOwU1ZTtBOO5LB1aFRW
rEI1XMAvAhsRdOeOaacsm2gV3hLvszsBiWF7TsiZGYjAmUM7rYeu1fo+4oBNZVVT
1EqOtyFaShIFnSiErn03bzSESVs3sHUWx3dfF9aS9T5kI+wMqTOpx4cH32stLCG5
wnKznZRI4lxexuZwBS5ovS1Oe7E7RTOS/ONFzrkORUU8GLdpqBBAyKGqsVCbtMtH
IDBeZCUoqhtlGnMS54M3csYMo0lnbeN+GBeusk/MhJinJtX2fw5kKm062Zi/e7QZ
NE1Cokb0pe3Nv61G82nizE8neCdUFni/iwxxhT4wgHKgBrnI7guZUW+OvSeYrMHn
Sp5Dzlu2M1IJlmRSDKvkAtOgrTk6v4O4QSgI0tB0CkVV/uT9KwLk7qot3VvK1dHf
SbqUVk2pNSGXC3o58rgayadSd7fUfiPKacFqYsqJ74E=
`protect END_PROTECTED
