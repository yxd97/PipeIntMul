`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9epemCxD8hi7RBWaRvUtzEYYWZjydIA6/SAcfBu1VMoGpiRytSUwtdKFj4FYA4u
ytUMNJA+cc9Q7CCzFaN7IZVkO9ZnC97PTOwk+IgXvBwIgxHJvz/mNponfc/HyXo8
B8o5PyPG0jGlcN/grhr9Np3dxSdjMIaT8COK6/E4qFX49QlB4PiTcIRfi91LKGHG
frnm4bapVrHg/SVX6UPP7lkDGsNCSt2DsU+ycOD8zRFasegD8d6I5aw20VgcNBUE
oZUkA13wwkc0g4N9rSoqQwz+ZwMlNhbS1rSlc6S4Vi18X5tck21OuCTzKHyxoKo1
gN0inKCLXUH4Fv/f5MTLfujZjnLpCiB6BminZa+Yu1wBbxwPfcCnqZ2OziaYNWFC
/AImHcdFb5H+RqG4Srce4pQyTyO8mUWOWrdAwoeGEe1BYZksllX2XsVhzp7++5qp
asaeH5kRstAHB1wHzr/tIgwvJSsNKS3E4lQp7fe2+/JYzRMKGR9b7XC7l1wnMFNi
IU9MGOTvkh85sywz8Gc8/+dsDHmK7K4/9RXURq+l6Zb/dU4kVyJL9e0mLHxA4eII
`protect END_PROTECTED
