`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/qdQxQ8I9OouRxedVS5EDRTxrFJxqiBvXrxEWTWUfbXrkhIe5VoqQdVvV3PC626
PzF+V/KRuer/L0J0964N0D3RmBZnBkToKE/e8yNJoowMeJThlDminhyaE9VBJgyu
VnaV7v5p+oMg1D/xIbosY49Fcfew0rkY6hxmvmM9d1r3Ixr5P0cHjwK2YwzHa8tt
vlzB1yZ7CMTZbAtp2sfK8chB/bRui5l0D/j2lADx9qj0SDeqoO0gSfaIrUMTs4r9
5MTwKBbqA4oYbAlCThRvoSFuMBYwBoYRMtTCLAqlBlnOkiRHfDpkvl8NmMxytwrN
GThgl1FIKthHr//leDVCwA8fMPbpLkq4KzM/M1a8XcRFE1xsjkIBBpPA3xyVOvBe
`protect END_PROTECTED
