`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
stjNjP7i9UNoxe4q7YSGFMoJErQr7AOxG+c1FnRCxEgSP/RsIHgGUvKawE6cOsm9
UEjdK5x481MP+lO40mYfCico2TIgt9jlncePvaAbNMxPK0ew2XIpzKqYrDdnl3fO
du5ZD0bk3XHmWaJxz9JbMvOAIQNtWFVmKlviHufcU/5xGDwxoOXJqSHR+skINgC+
lRVMo/pAZxWObRDeF/QHOqxQBXABy7nv/fEqH5Skf2w9EWHvHY9V79E5wcS10ECm
LHHBVf5Tr4wf+Vq2aSBC1NXyfFo2NtNDQ6GZ17XXTbUT/L9zChHyJ91ZyOyZQrTX
0lWCjjFo/Ufcr1Dxx170ldYLDp9sLQaj8+hQrnGiu2HlJQM/RDkkHrzwyum/u/6g
neWy6sUgtdandftcEcfhPcBZJDkPudAK4LdShAMm0eA9XWdCJXzxGL+hePYuLKgQ
D6tZ2cpCI1lVb8TCUBlUsaAWyrxYykTyyGrF6uMsve7k85BW3dxBBZODk/gBvLk/
`protect END_PROTECTED
