`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7MTX4HGqeIXiUf3rQPVVlJc8LaKArCuuyCdw049YP+AxTrPD2f6lSFutVWF132p5
BBsSL4shB4XmugPVQdAvm6LxKKxwdg2cpq7XNpU4MD4QiOMD0IxprrnsJ6HC+eJ+
tyUphWZNj5iu04rSZjJU8ggufRjLP/OYYSjgqTgeJ7ECHQOD7nR5Y3Q8AJb2Ozw/
xurRsrXTWqZc6pXnXei4h0EARGTE71u8cZpQHLlHuYd2xBDBFGlyDYhjnKE0AZQt
jXF5FcZ2M0/DHdh1/Pl++hPJbcBaVOoPtaBYkgw5kQjzklrfmxwFej2W+T7eby9F
MueoHSiQOaZyr7G0Z4bVKJtBcvx1mnWeAjNMlU/0VqQL8U+HnNFs216Jj2f3jT9p
tdutno3J5R9Iu5QFTciSopWcgKvW1vWd4Jw5yyEmVlAGUoqJ9nEco97fXt48InTn
2medyMgM388zCkUg7Rk3mID5N0FKHwRsGWhR9GGcoE44qCfTBTqedT12+4xBxvCS
GBgev/HfkpbAtiBVi4IZAD03c8TpPmv56VHsccwLhY8yJr3YnZXZJAOSeEJlgrtF
vflmsaCSH5f6nmRZLnE//xTGK1bN/pLlGx6bC8qCj+Jh47f4GWfzL4IcDghhmLUD
CT/yOVxzeehvc5Ri7O18ag==
`protect END_PROTECTED
