`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yt90AKKcT1pYnQ21RfbavTHR4h1m0vgfezxW/EfbtIXyl5ous6uZLwE0HkgDKA8B
14njJSOK4JPoFfuVHqwatHqXc69I0ONq3y2XYYpPRiVfVzmMSB0y5yMmKoW2K0qT
v5PPaKiwrlosULCiudGkknHEdjvyI/ZyyD/fA2TtwYcFL51iHMzaC1em1GFDas0+
sLrkJfWA9ZEOMWhCUCBcDFLyviaLx4oR5CSdNQwF1sVEYVO/ZZjZKYCpVbv9l4zu
jqex4LieshEsdITuAx1BkRN74HMkLTk876UVb8jEIkm7KjnkTCxFNbltQlcORy8V
+cxDw/W84T1nUqGsETkY0QQzJRT9TB/WJBtQPiyGCWA3qPYbFFw38Sa3zwRjs5Kh
BI3njBnvcBSGI8wRHWVKJOX3bPVUOCG/L64nGZrlmW9BUspWQHf+qyzEnTRQEhjF
9ZCdDSRgRlBlOarjN4nrKp0WEMggdD7258S2bYs5hYVVUkD297cKLVysyMmevBzH
SyuTll3jPS13IttjPg8YnPVYBvjvno3pRL4jCrBQxJJ65B5DEIakYMyLg7dFXwal
g2u7Ov0hlt5TAGHzDnqg/h88QSKkyRKjoL92/7fudQ7yZLts4BwPjuYrVyBaZTo6
HKyOt7i1W5e7PaP4vBhcOKZBMKKK1r12ZGQy48FLjv31tOQ44glNJV6YnFJn2NDD
1g85lMDAxaemNSJ41SVYw9IWlWwGwKZ+JVfuhFNKOVv3V6gI4FcRVRzrWaKv8BMU
WxJDhki4xbY3pubnR91Fki/xDS3GJZaoBa5TqJA71IwuM3fcE4whIIDBoyztgkSX
vG0i3C14jWrDOe1sIa+xYuwmSXZArxOGWWxAlu/ph+TWyYXBOK6As/ZMjDp+pe96
W5uymT/D5x6aoTpCOvVN+i1ZEPbBW7xGUjZU/QiJCg8yB2ozjpokD+TkEgW4VHYz
vzk0pFEjLLLXO82j3nSFjkHgctfohCZDmKfkuw+2vZ1asZ5g+9/0h2tm1oRHy/XA
5IgDRJ5qgodkY2q7lqYzWkyowR4FBbrXl4IKod628urYuNzQct9hKj0xJ1hiD5uD
j7LRW7VwsuTvaLqGD0y7mSKcJfq8Ldf97Zzd/KfpG5ioMOVeh+Im0RHvgj211fE5
LhF0sUxrl/1FVq10PlulLanhCeROpUi59IxjVe+wEn1xhOuOCd1LcO7qr7HRLMAX
m1/kEKs6sm0X2usMRvCpXHWK7DbifUkJsh4vVzJ/RIZh8EDcM2oEvhHWmlh+dXPk
RYKPhvNSNI9+LtsaxjFNIRCVhkMJ1EaEiZvYnDaYBp/kJPQseeVWMasX5FH9LZ/v
/mOdsRIHiFlyHdTvOEDvSpsNIOOMakuSZjzJ1oRhuL6VUVQYQQqwqqgJreEoXFVP
2xWr04nDybEZcHGkeh/rFK8BDl70orm6MAsGQa7l31hs0UE2jReAlYVEyox/qVz7
Ft2/DMkRkcu+oHBw+/bzDdXwaOdqyJxN/CQ5BGlVpQnFZR6fWSlHJFNKKKaPnSs0
fxmcXkMMzfVwuMyY3rRgeUMUnz/fZhnXr/fk7HG1reN+mBCGIbr2mzcTG6187y9o
6aKMuY+G+w/zAhg7GLSmHQqFgdWnLoYObZORIiCZDIsiqr2Ecx7kdOjiTiAJ88zG
vYmu4VrrLhn6h2YkJxQ/CTehk8Qr/SqcnktYdZmbDf2VP4c+LoXS04qdppzWIOmy
93UAaPhp5ZSgiBB2RXhA3G3WQpAbg/CbKYfU/z3eqTOhc5pO4cTk3KTGkYQeeMak
igB0+7eVgC0oLAtlfHwqkbLwU8C3qRBMunpbdUyMcWIDcsE3urk/H8JXnaZbphnG
abHho9sTyNqnqwZz3jBYkE89PBRnGcCMeZ0Hkm1xGkD3ykYyfAYpaIzyb8AKMArz
fpP4qRU2MjlIisC0gANPcdLoYY5DPHmNyCfQTzkat6jY8H3W11tXPiqvRF/7rj4m
U1LJaAdF/F6xPW3tNM9C8g9xEgm+8T3RhSrpNqJyGKF3dL+dRBjRd8ZNRTSUdiQn
gT93scxNkj/xjwRjZdT2+dn0CSygHrto3ZSg8ES1P2OyYlVjNMtBHD8GIDxfHJz6
KfOywkORFyDps54KAIZWsXRiDi7AZx6VLnR1N9mIv/lE9dSRhSh+7nPlqy5lGFX0
VPxHCuhOb6BJvrtn9qVPl3/O7VSx2HbRGHsfQhcyF8P5JpN2bNKa4dA2zruyALGv
n957xKHolJtlBj/XWXSKHjiSTjlApmBumc5WQ98nK0rScuqQVkNgsEZSb+wxh7JV
xtQu6FZvxMd8BQEai9Vy3Co+kg0OfDT6VTN9V756iXn6w9FKLcI+xvaLa7o5mCAO
WSu3gQdgBjTJkRKfXVAn0yL3cEhgPTp9DFNVAdHkgsoj6/+VVFXbztwHrcpp2brr
hi4t7FYEfvBxQ3NB3teWmiFWywjVcdC2O1I+bAiZV2hynsTagYeD/07tM7fycw14
NbuybvTTMoTNTJqLP56kbunZRwpSQP1xLN3ch8ytCROjvjUhmjKhhPSQipWwXozR
7c7+PsuHK9duQBB3He1jmxBZDbm5RiSSoqkGsOa57AcuQbuSoc4PHOpHeYAzRoR7
KldYzbCqk/3TO1TGbKoUdo1IHGP4qoqT36RGE21dpPM1CWgdQepQyUyZyJBffQ0u
jAtyU+4eofJ08oIQTs9NnT177Li0MNv/M3pIAM1jCAqB9pWYX6P8AEXYVa8YKbxG
Hr9+tT1t8lEvl4QyOaz1hXGCZG8yHY6x5+cXEwgr3mjoLscINCzkpvok0FWul6CV
QVm4H1bWcqUp9F90yTwioltDDCJjcJp1VP9d/FLpPkUeS2Ccn+TrSaBqaYGRrKBn
u5MkSTrMsDD4RbCq/YO1xvxFbekjaJZD14KCm6vWBKF6x66Xuod/8+em1UTscgB8
pp2n1lvmDQ1bBIKC3Fn6DOmuzIYmd34f8YFn8wTBBQWP/0lYPn4ax1SGki7uSHRk
Wvzwhi6BGOytuI6DWV9EwwlX2qImhFONS83/UPJqtiPMaEG5QTukLOr4SDoYsQi/
0h+04oM3TnAE/oYGBti5kKxwn9u8QiAlvx7/PKqPwt/L8qBkNgDRJC8VYGb9HRrY
ZmKWIQq3YdAdnj5+W+vVDzk5uP77WygHbg0IfyZiEcakv4szeaJyMc6NNGLUtPQ5
F00MSVuDvOCcp9RxJfY0eixspeswMPrqbOC6dNCe1J5EpMVo5PncoF785vJT3rsD
0DUSImbN8lW1/QmlHEQqzNAisjvNzuja2UoIxbC8TicvGRolWDNajqyfSHBqO7E2
DW2MBQoOg7OM6Tel3XlUXAs/IkEwjwSV5kONL6Qjb871sEVcgl2sTaFjiVtvRlYN
cd4dlZ932ZaZvJKDjq+T6WrWtcOft0YgAqKZrHNAMH6bD2njwDfoLthPAjZG/7FA
PECKk+k1dC3iQT3reHDEEf2yZci76fCX3jEK9bJBRRTOgWzc+XjHVBQlA61rVGBx
mDCz7FCODEIJZ1qG+UpsDfd9TFwZu4zbKVGBSBlJQEH0I08BQPRuM7gzRea3DpSs
SrdC16KudC3PTB9UtFiLjbBA5f/7Vr8lNIcg99UFF+uWVb3dkzGkXX4u7/M0Qn1L
US8e8vxzcIU/mBm+JppVpDoOTq8kskmF7yCNKSZgZTukROTieWLa9I+pDu+NOZpH
qyrF3ZTLQeVll2c65iL9HjQJS8RYeoM317rkUm310M7TbOg41Jm+iN9F8qY14XAt
L1aXN5TvWAURZsOdZzpioYvre5DqqXujb+iDvURpmTZ4BurzrVYnKquOYqc5q/qi
l4yXAH9aFPL07aglNdaCkF/Kob5DTOPbnx/PXIf2qY8R4gyA4eGiPF/fiJNLu9EZ
xsFpiMT4vWujD0WZrYEGiToQrOUpV8lqOo9uxIU7jXPq1hPUGuNUHNhQSx2giP5+
i9LHnt1KRPhXsBKtrSv4akghZ0JAp5pbKTSTFSCPC/PNJEbZlR2Crqy/0b9qEAty
LfkQb67yOMRwFfaABsM/ITqg6VJfG+X6OZecvz/6/6dQUl+7wA9H++0Cz9TpZT7P
ouegqr5JPSdR4psqLlZ6v8qUpw1n1TdA2dc80W9sfflU58j5m/TT0YsmR3s0pq7z
t4Y5TgVZX8E9vqWLNSpLh0WuV7zRJUJoIiwysVlmwLQcO6AkTGFTsftEM0otxqKo
SjmaCaEdQipCH9n5anG4G0bjLpaPr1jDcW+tQxkW8XYOcNdIMLDvfbVMp4RhydCW
F7xTHdnTzjO2M1djZ6VUFXJNqspAlXoA4MGARSdGoajyNkqBCq/LEayLf6ZMK2aD
iMluj48mG0yqiZIanh9MybY72g3b+7hgAaFzVpFRz+WBfWnv1NbKII/ZHB+3B30U
f+eFz6aBOdVhWGkVn1lQj+rXS9mWdRoqfn/DvXLNmOz3pVpwIYAFth44rv3p6M9B
f7XsLNVsqzGZBhtJxw9dUR4XP0ztthNZzUkqATFSstLW6AouL5wiVbvPckhhmYSt
r7o/b6ydH7j3hLVRezmJv7K/hyo20S7M7/5TlGUZHfflI+hp+0dv2E4AyxzCbj+Y
STdYr+rXCoE0zUCnvBmUGAzxIMwd2GgLSOLzzYGaaiPNmyr+KpUVm3DWBeLU/ZAC
ars8RLnZvVQa99RtBEHwOq+PFN8sezVDWMyoQ8T6PeV8FiznQrgR+UHNBLv8g+jv
7UBXzo5gIe7qJqKQBWTJPrh0tnWXgep+EBsDCgKcQKrJ0r/JCfVslnkSH7iHvqrn
+ZLy6dFhvf4/el0Lzn7Prlxx8Sgg1n6+DRD25VRnVUiLQKDu8QayxpojOQuPXyqy
yeSsg9OJ6laPxqjKD8eyNI/kcHNXynBKyDcLeF4/uMGFHuFj8ajPemmpDVDeJ3Oy
aGTh5QOgA+qAmwSTETr7HfBDP+A3oVuOwEf5HGzY+OTI9HhwPLJ97LOe+G1JFOQK
mTQ9g43DeWABTvOnyQui1UPHXCA0todkfd+XQmuXDy/dBhCb9vDYAHMomf4TTHlK
rMQdklOhFSBhOvQXTsbRVqoGwD62kft3sy11hOJb2YwsXUXWghinTMLu94yinLfN
Fiw9LRZa1JxECy7AXUsN1lT9ZV9+BJKLVpQ/uIPV7qjgQRcO8Sj2RSiB4aV1hRDq
45q7LA+V4zLRkzPbvoVHUR4BR95iTyjyoyUWGJYksFQseXM4NrZWH1KFIXsIN62E
KnpLJjWUQy6rAh8mDzJmE6ARew330xiToRSY9+UQTjxAlGj1zhvNOrFrFMkZSkRL
G8ShgzrJH7XWJhNVHBkEbZcLX5BZfn4px47fizk26EexxSNU4DmECNwgiCi99WEA
I53TaYbsPuPnKAVkDYjOaLMnQ6gT3sKU7Xinqct7oyVRqmUjdgY5KmCbwlwZJIP4
jQE0bIvyNpJqdP0VQlmbk19GuRiz45rTkD+KrSOH3nV4hFeu3dDYtKUUK72cYXId
hJeJPkJBRJ4FpipetonNL8c/55LHy6NdAxxwnDsHBNN3P3i15Rzf6rahQ94skRQf
U73KD30O9JFeZ/6VZAlDUy7FyBygHIFXILBq3ONrwVS+Sl2BlzoDemGLzB1wwSEz
Un3d5v8kPkp+CNtVueRleYNbf5gde/1M9orfrxpDJNHXUobsayW6rRx5kBruqVen
0VaUCVvmC8pBreikhRumOjlBMR4t21guayZURojqEPNi7L7SLJYDIP/vXDOy3Gci
HKZtDKJUc/gRal0Dbleh+YtndUQhD6SlHrdBfq8fSxjLmdJKWvGKUXHLyksCRLIx
LuLHrIJCx8Y6Ca91K6+BfOOD82ArlXEBD86/1Q9djgjaz38E374rYtSZLuK7EPy5
rX/Qw+FlwWmqS1/VAzqZyJl6sSOI7tZ4lQhQEToVE6WpABXmKWIaT08Leyjo2O4u
ZDygckZu7lHdsdJKHnXD+EshmozBXE8e8EY1/U9AButBj6w/Cb66986T2zVqy2oh
S2twlv0MenZ/tKz05dsGy/Ty4njQ18mIrsiEQxf946jys0rKVshvmgmmRTnZhpXt
Q04msliPP0T+DPnuo9/ZB5wan8KILhq+eEZCuIb8jdXtVa7Pvw3/+j1YlOyZem7I
Eh5R27EYIwV8bCQNaYC0VnDVLZjd4KIhy/vKdPnln1qkx/GbbZN8R6sc04zbXjow
/gFQJkanQ0OofMu4WwltQaL3qXZzV1A7anbiLrEvzUEUnPlQTj6NhTcRKva6UGm5
mar7V8yWVwiNQTXEkageCtHs5v5uMaJ7C81AefMQz2EeaXlqMvWN5ogOiWOZBtiU
7AkxBnQV0v7zYGq8K65McgUVAvu7Z3gnKnLJEYZPms1aP74t46vHQbV8oIXblOa7
Q196nHNmCAxQ8AV0FhPjkEuvo0G6ygHhK+Xad1PJ48THdlUe7/1/DhijhoJKGrWN
3kK854fAtuoFzY3E1tc+fdm+uhodT3AbVt0TmlHgsif5uCMHYeYGMjPpquZ8+CZx
WpXDKV4JUPJPpFqynmMQkVHvWYUCS2dKoNvp2McT2SlBx4zUcM+0xEicDtNWHziF
TeALEiwUXJBVXqhwN1NU/VIkyVUxOHtvst+7uMQPhlBSGPVMMV+vHP9LdSIbAUS+
Jj361XC1OQYVGqG1X0P5FrUur4diHubfP41VGnDgUNdQ4y5bErW0xbVvlT5t92fF
pC3qOcaT6HbvkaJaJnIFY26n8wcrhkaTaefkA/+q2lSe/6GtYuznkc2VXXgnQ6DA
OBNIyZnUm3vrt4g7c0/6FObcorxh43MErfU+9Ro4FDOxkRp3DAdietj0R0YIVpNo
tnLSh2qViCWqWuEMiFbvMQl3Z5av/DaNO25Kxuo5gZyMJZfRdMutlRNTlOKpj/jh
gZg8WkQCVmZkPURhF4pqsJaw5wPb04F6mGUFmTDDgPUrKK4WXldJjuGrrOaSoSu/
bj0qd88JRo62zbOHX6KmJ2bqLL2LNMJX56277Gw55vlxW8GaKfJkY97u8oko6z9i
4ocOO+VdhwY/RMeAWk4jQX+Z/NAvQRQs4dyaggvw/pLPLe2wR3DSr8Xa4sOGOcU7
8Q39u9/RxyrMIXACh1Pp6gZKTTh9r33yJWtr1acqnG80nCGH+LrW8UKsI53dy7Cz
sBgfs84Gf9NRh+Fh5KbjMUKvOhNX00Zr3lpY7V0z6hyzZIKmrDua6jr8KjExr7BC
CIByydwN/KWq+ig1I0BhV8P52dAKB///VttfVj//7+l6ldMbAEtiJmL1P4KubKCb
WM7FFbfJKNFWp2OZy7klZNSF/OfV9RT5ZEKxtQ0KH74QOj6KzCuGgCLaTrFy4L/y
9rMg8SoxcGIfuIIsttbUgFl3d2ZzbXMCbVaBoJx3xkZIoWo4/37bJwmnP0kl9H2u
FMpnBB9UaP4hS47aNppoulAd7d9uxPiNgPVCHiTxjqy5H85dgM+5ZrvYHfBv5JyQ
ziPlbAYuZs0gAYbKGzu141XgmvM5sGWyIPbwtpe5xoF4FNfF42NUvi9Hg90ljFcO
IIzo9LW9vsJkMivwixbSOXCGgJCYu6p32M/pt90XHhcTOlD160PZf0F/2tw31C+6
TnaXLGW/TY6M1a0Jx2MByYH1WPFkXV/zNlYzDqBaIVjDtiougiaWGjlBkCXCrzIr
uemrMI7TeWfvSjjAYV0d14NBwtwupT8NTraxVhSIsY5NAtcV/d32X7fXVn1mlhFj
hVegowH0ORrUHILfdZV6XiM8O9OKAgDubYZi5+Nf+Tv483W3JgfEHOlCH0YPXiAV
x1JKd+NSrTVM6KfzUElBRYJ+lVlnkE2dG6JShMLRia1EVchhA1+2Hp5ehZc28Kw2
q39y3MNhs97OgW6zpFyy+g7lj9o3gJtAPbBLX3nirEIgADdy0g5hGlxF4BGpcFNs
09dBCZqKCckLbGx1d0Cnxcnh2EdF/mDHS9cU4ctuusH0StsoqWyu6wW1GoweAxzf
96Bx/iT8+CBOwUY2AqHB8nrjUWO5w1H1Vf4kKjNhmekYywmFH6hTG9v4IKMJdl6N
IVRQwE3G8iJQqVbsL8BR1ZQnsqnl2Fig2DDGwhMxffCk3Ro0+EmY3dBe7Yd5xRvM
pd99qA8onkHobgO6XMF1EwBufWPHsPeERwgOCRJbdDUBbX4r727Fcb+1etaa6f8h
V4YZHgAkjkABTWkLb8tTszojaPIYqVEMIJ1FxMfga6xr5GNQHAFUIisUw2LY28sj
Q4SO9G2mzKS6BI/hmctfnoKY+nGLWkQ6dJuWdp8MRcDJhiLHYVVNPyPwb57fkP4r
rrKfgwcZFArBc0zT9NvdgO2AXyLzDXHadc0oZNH7uxAaJEDeT36I6Bj/IWKODHW7
bWupB2DX4TtWoOE1/F5TCHUnctcFNPAlWLcoXGMIZi+Ib0LdzjVvi+OFUQqzGht3
IDLc5Q7kVF1xWbyfM8LujpqOO8YnCgNcg3zzk53ZI+WEkDQkQsxftQ+QTedj+0PF
8gL+LwT+15Rl0SJBojtsF7PXdvcrBUnFUOxzs8+HMP+8gPSY+4TIMw61CUzK5yBp
KTykXkfEpvhMkhPdd8fKNVjwB+0ytSTQmV4wYqsKiNOFEJ2LtUvrn4V1gwF+g8QB
PNzsxeeJCYglTwtnqR+B7DnjF29eUypyEhVdJsHLSOnn4oiTegWc8EoyFvzk9ae0
SIzuM9uGAaBlhuXiYgTC66+MvvPvAHv8xVcZ/p9shKJr8QYHxtQJB6r/+af/sW6D
vLSoy5qnwKVkyuyAKsvMr9G5ojcJ7ZMpqSRejx2eWKjAsbSrWTFVWpAJSGId+3ZX
b1qjJkRZop7ToLrlcelSmwq44c/72FRipHORX55K0tCJkgkRee6MVjzs7Oqapk57
Vfy5A5epwz044CyBF86t/3RzRnbjdhFl6vq0HxoofqqZ51Ruv+r/KmdM+zxs9jT7
NmsWN6ye9PpvDIh3FH6CnlgoA1P5wXFe/jjR4FtSLX67Z4AfqfgGAgQapDIuEVoo
0BoWR44tdBz1O/l1AZJE0YzkCiGFPlOPt3UkfB5/XgI6caW9OOrNZLCfcAH7Yxxt
plDfZCmODkln7eFui0Ze+xiB9ERVlqjPoi2TfIEQ1As1eQvlMlGnDe5kMLd116gP
s3r3LN1SVv4YcQYecZ+VpJNaz6lz8TWB2WcePpD5ki8g61aaQmEF57EuTlIYTtaH
iqFA3Zi0n2dJ0D1OzaA4oB93/BOjULev14FtKixW0pwWvUdR2idKcUQsztwzNgzs
ZfyE4NCmOM6hPQtnnr/yS/UIpd/GRcjWLR+G2MSjlWPsqjnDDOmc7J1wwwoWxfma
V/n970r+Uwmp3C8A4WryL/1XvaGOwIwUo/xqwsMHsvlFGsDimUtrIMDwpryk5yYT
xT5DFjh40lbcIuFrW+iU/HEh8VkTGlbzrsA/GkiJeY9i0ljar4vi3er4ObvdZogv
+G8li513Wqlw9IgA8Wa1SydeaX537qoSBZBrTQr24DdrJVE4/EDHd+nvPq9bPupT
pnv+ajY9LM8Y4RKFATc1uehes0we6/EKlfax0GGJZq+DHbd7K3C+I0bvixXa4fuQ
nCoY7fNKtmITi6+KuEuue5TIqRkB47fbx69W5SAno8xcAfsf5Z8hrLUY23nyihDD
USb+WcOVPfSOmJhINFOy+rVWH0cO23iJRw8kDxis0rWTn+iz9cEf2D7Ft1icrt+f
51fhpit9OkTPPuyC3Doq6khho4P0CBhrzwmNikFshxx5VySyEm/YOlATTj29ScVk
UNMQG+gQrlTKewC0K4uXspdMa/Lhyuay/8dZMfKkvssMA41TYgDHL561CJCUPrGY
12G604Oy+Tf0o6Uy2CcrNlMMQw3rs/E72fwlTdy3fbllTEJYwEFcLsTJ+nHnw0ch
Ovt9k1tRcUce9lOZRYwZo+4YdXXuMlLAy6mpbIQVpULN9sYc5yNzeMRD0hw4YIjr
PEoSzPyMtg4pniYVpJly45CzH6oXL8GE9G3WFBZiYFkXuYK4LqY4U6oLpUNuWIdC
yKNg/On/8RxQZs6T4Ku0Hm0tQnVMbefOIdE/enqTggxTOUCvxzwCCsWVhPtZmUb/
cDMUx8EdedTYbY86xO1RYWE1m1VbxVdQFKYjqEdhzSQaKhe1fNtuYJ5wZ6tQMcm0
t+3CDsTsF5dlzbzi7gJWUphbpxAiS43f8kxrhdWYZgIR2nFuCEuQPWSVyPr21dxI
E49YlP64p76HIs56zCIDPh3chH/NpajfpfYNKDsFfnlp6691teA2c3T8AeZU9s0X
T6jt3n6IJpgXs8MeeG4Csyr9v0VuGrn+A6BVQ+fYU5h2q5rAhGmkN8M3U7RFsbwL
43hsllp56Z0jL9x5BTBpJW12cuwXCOvH2Cyzhk9DrvMJm73nAYsMyhDumXT0gTTK
YMmNRoA0jl/pjJ5Ois73gOMRJp3jYldERRYRJpjXHoj9OvAcP9qCNDWLh5obaqgC
p0ZRkOyYBYa3Dc6XKcMKQYhulWq4T9TsSqtOHHu2KwcAVAPh8Y7kVwq9VtAc4ldL
guWpDjp7k/fHTiNbeCvgw6a4IStb7L90KNAdE2b1T8USAfIozBBErR4vaMSHptfX
pzpfOe2dG+6S2SnVdJM6bSBMmOlEW7G3SHT/1YrqsZ8q7xufZrmqbPpscL6HWadp
XL2xANNSNPGzPKPpe5HLw2f+NewFHI7PdFsiqbwvZ+8iJwVfkGaAoaBcmnzZS3J/
+kbFIY3xLNRKFKl2t/LPTLvNhuGVJAUVQdxh/suQGEP2NRCIrOj+1IyD6oAWefzu
/+6X5AYdIi9daZu5mfOVhsW8qfqbxCQfP/xUPngrL9JaF3M+CW9mSSpdwIEF01i2
5yvI46Qru2oODpswfLZrk71fGBAqleNhcuKJ1/4WAAWlX51P+WVK28C7DqugyrGX
KV5q2IMex6pRMatKYzxORHRIipFvVUV/pp+HztMW0/OzQ3J71/Fh9Yt/Udd+Bi7F
+j8uIBRKsFPyRM+75sgJevubNGq4Cxs2j84+sjwTE9pCd7o4wOcei70BUp0uVupx
B15Lq+ogQoChshG8AWbWJpTZNdftJliy116QZAzDnt15dg2T/U5PoqGIib9Gz3IB
yA6Xc+UvzuhtuTkeKtVrRNm8bfEhIBCdyK74UR+sKcQp2TCuSfoh2FKuznHSfcwc
IQtu7iwrSy6xLhvxmVCyIaj7UDYz/e8vRQUO62uUb/4pdPoEUAADuVg6GbdBKVC+
qUxcqz/D//gSyZ/6trGvol8wTg5slh77q7xAQrk6mLcmMNdiJ7FUvfwLp3Us0lqx
LO0abL3hqbIWmxg8GFp7k9HvAZbSf8oDKcZ+pZk379PH1fqJAk+Vve+wcBAX3SI/
qXPS0dvhBljMH43tmG6jVeZ5xrlB8RsQ2fltDNp+958bHYAju4HmJpW7trWNn6+Y
tvQda8sNw1OUMoZKUmulToJBuhOuikkOhbcbatcgfvrYbQMJMM4wuhTl1KswXrIh
wxSlJ382mkwivp8AMFRMM1VLRxEYu1qbtxXFLdu5YzNx6ZNaT41HaCANikTUlMfI
V4BI84vq23cXJwetH5T29sopwxmIlf1EmvjuKtz3KF0=
`protect END_PROTECTED
