`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0dmCeVBsttpxh8/luq2QK9qa9MnAg+AiE7Qj4Rg+d7OgAPiHVHaO+AwKjUbwh5yw
5XYqMT46Xya5/s1gyhxFeVi6lW/TCwqh9uf6+kxSyb7HaMtf7JK9r2HGacmcwh0P
PaZg7h+TsMQCIoK7ak0dbkvSUqx9ENYiPRO5UZL8tnjR8XAynaECPjf1WKbWv8L0
u1VkN3S7iuKfOwY52h2hGLcZjzc9cM0OfUL9cXgzH1xhAdI0qEedpw994N2bHk2U
36o0A80lYx26ZJnmmkln9c0NUt9VgCAqJIPPfhutWtCctUjsW1OMxCos1Wvxqr9Y
quLGUQic4KeiyysI1Qw83/WmTWphD9Xr3saint6n/vIGo1jgKnHQ6SSx/6bQwY8p
KXZqGf5xU3EdZ1OSyUsc0IunVD35u/Kbse/7GQBmmZ8=
`protect END_PROTECTED
