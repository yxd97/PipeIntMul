`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZSa+BHBR5pKoyFseljHtIkyxVlX0E6ERetpuTaXJ6l1V5Xh1wbPzOKzCLflIlut
GIk3aEXwwfSpwsQDXwXTnbvTOk7TJuHFA3tvasNx9b/J9L75MZwgwkiL1gdCrm9W
X4obdYyRRoWocx/NxvBtiC7mzvgkRKCV1BFYlpk/NDpixciA1dri2hUGlXFLnQjV
2Rj5UyEvczfBAY6F9UOiWRxsCMv2W9m5G6ToXRGE7wW5G5X86HbGlGZFTN4ffSrR
Bha1sHYqyy9WopSM+mu3fMUJ4PU5fC2ikHx2kpfVP8c/ep5isTLDAUuVXhaLbLcq
51hKRDsYBlFTLBQjskZLW0UJpJuWBmaljTVSKriXDGVw338pa9p13/3VWkk7llgz
Op0EU6a5QOv7Lgw+wQIcmB9C2NmAY8pGool31Np/1bZoQHvElirycQTPizAJE5LD
A+6sCr+1y4kRMQ3FjmqO5v5EfZC00I2ayjUdcTq0GQxJDisFDvMKStl1czetIDtG
S6TXOrRRarATl3ocH8sbvm55dcD9ZVsMlDtc3kwFV00ThUN51XeyOgNAArbOtZro
7HJmeGT1ccUioyhGiRyuKoXJsEJDEqq5nUHdiWFzGOH+Jn+oP8epexmxNxd5WB7b
QybW4T3iyLQA7Tm2vlPZ+6nOLnh2ePbq/pEWh+k6tTUSdkFP8TQxt9ojiSAsbfSy
geSEgdfiDLjfyRKAKHwsa3haXoo3yEPyLZUH0L0tNzp6ycLgTva7KNFeAN57H/bp
t3tGZx+8U8WYTRbeMcaGb4HSorH5OXxoI7k9io5+2gNXHLP/O+hEKWD9Z6xnCC0x
HMrkBep/Zo81w8HNoJeqr+Er6HeAZywh9nOcE7EGl+gtwhRy/okWjWv64nkER0I2
R8JVS4Adnu5E2WmTB8Qupqbw4Wk5BlbtHjm0oZt/GSethBWLeaA6bGBkHXMEFhos
+x6nTdi/6BUzYGAYn5XXL3/4wGhhP3qKUiFBI/ijPmWrK97roBYHR/Lr7nCxYhC9
6NFQmLRaV0i/MkOSXL9yjGeDms6zUQdJfXpIZ5eWMIqg9rbwwX/OrBe0954dla//
ba5xUhc+ilEa2hCGU8aHIFziiZvbDhdNDmG8lNwZ4JH08/jpMBQH8M3WuIp3zlWv
akMQwtS/2juiO0RDtZPQvVYzFACasqoFVIKoRBakjMvNgoOZbUW/1gy4jS++jKk6
+VFxX+29YkM7JQsp6d+vXWUAes3UT3iMWpwUSLDL8Gr+96GNYoryaGK9ePTnfM71
7z7Nxa3dwHGPVzRUeEHvQs2bynwOaZHarp8gft+4ZeNKn0AACVugpZmx9UFNqWtE
QobzXJpuScqWTszvaI3FlX5xPF0K3+C94IJ9dbwq2bBeQQJZXUDaJFCxZYpXt/au
FlM/n85aLM9ekedAv4W3SE+alIBuDicFWzcH/EajyJeklj9wPHTQ5pqBlPhEJzrV
azTn6VRuk11ZhrdYUe+608I2u0spK8zlVdxH3ESv14mRGlAN2pWtA5e6JhkRMPNz
lCUMNxbgqTxLQ0bx4rBaGGA4R6cECz53oyLC5U4FOB/JyOQZ/DCEaT7rffa90kVQ
fiVZi9nsYJgriSsd6QS+jnUmcyJe2HC2elj9zkrKOwDdwrkdjeBmL6R5eAqiD0nx
0qV+GSapx3QVZY7bP83u03gBddYfB/tULsqa1tlP8rb2WQmOzVP9kaDMxUvRmdRF
2QCLON9nuuTrQwLVM9YA2Fs+f6+1Mb/UJp2wWG7ldkOeYHhMmWjcJ5DmT57E/rz+
xwCdIAEubvWye2lDyzk115j6w6QwDk/Z9EMGa8GnGCGds+T46TH/nfp3keqCPq2n
Tdk3+HczRxlQKm0PORYpIym2POj72kmmSappHXVctrHS41QKKYS2Xb44SRhyZ7WA
rdE8twRb3jOkF9z3uWdBza2/SIIeLt0a0F8EO2mYcSAL699N+7XA4/fptdnKPJvB
c09BC36suco7MuBEcpVawpOqEvNtgFvUT3VOJvRyaXGggmygfRJuffDjlJgt4EL3
GGgFxXZ6PQwzGzYxiC4IXVE9LevsPCUBGWYDSD05Uj4zkK2ztknxSBy7+G7TW5Q/
`protect END_PROTECTED
