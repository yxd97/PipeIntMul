`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGeN/MgH7FSoXcWSFMAarvh5xCclVaeEziI7aoXixxBxhHAB3iAZ3OK1j3iUBaSl
IvQYfTy2x59/M+mW5nb1jby8kfmde3THunq42CEFYCwg2SVb1w7n0DhEKVOEmwCF
+2SCMcHEnyBioPZrFJFj5IUhPvCHE9FK0pBqyOUP3yuCur+zaie4nAi5uvJCyatS
o7m0DUQcFz0Hj4B5//6L0O8+7rvYtfKuPis7FSk6qxtRYUlyxbJjPuMDRau4Y8dq
I+sQ4ddS8Z6+FZeUozMAy9VYPCXT8/2180wQVj0NDhZauam0rqy+x/Pz6yyh2qQK
+AW8qdT4E1Nl2qYXiKXGqzEKKpZG9a0lGOWUHxvBSRq+pW+mCPSDNX9SY1djEhBe
45OmzpFR6Bk6+MegXinjd9YmNsoAdNbrhRuvl1Jm7a/zY4l6Zh3ahtNP2W0VvIYc
cvoU1lJu4OroVIpDY/CUTxaHt2oqJQlCzrn2M2SUbhZEfGcGZzmnbSYCTXxn5pj3
Bb3wBVdQ9M9a1ghIkFHugBs2FxP+1qeRCcMTF8qd692vkXLUj7NMIpAFTj8Zndrt
tafBHdxocX3j2DC9rcghQlvzxFI5wVlskaMjAGafjiTr9aiOkQP4yjxl8uO5quMh
OI0ZR6Rm3ksenfLAXVDnHPGBF/+GbN4eSeOYI2wzXFArL/KLTZZFOwxsaQofIf4N
Q9QYQjFwRBi4HPukfffwvLY+Oa93JHP4OzRAs71+ZKjM6f64eWBAoRXC+U0f+aRI
33vcpXEwdRNmyPO1N4XpIOlpitLDq+M/WazI8hPb80+61HcV8MHUWVdKVrmsWA0Z
XL5dR3YAcX4BKbjtgOKPef75Pe3XAyKGOE5PFnBfWOdgJx4K/IdxiVsMiVwzzFzW
HzPnXmJTI4k6XstTcxxDIdocu6XgEcvs5+zzPrROR/FdpCTNW/V8kPmxZwiFT9XM
`protect END_PROTECTED
