`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6anRn4cmV+5hZFq2jugc3yHaYkhlzQ6ZcfXU4e1CnGPynbK1Ett+50i54H/IE+R
NqdzGTl4azJbAqc4d1dOMynCACiV+4FzevwkXHHJLk1WCIrPPlnGuZlZTOZb1H6G
wkxq7SjeqTQzhTKFyb53afGOruNNIE4b12MJYV63VvDTf9yjMVwnU4WxsElatQ4u
hI7DkMfpzbvwomelD3g6QGztwL5hsKzZTcrjRAtrN1ED3pF0ml6oeXs4mai8zIfU
4tUJ6/jnpU50kxaVTkuDdOJw1yAXPl1VA9lvnQMpu0s5i377utuuEWrX/NEKinL4
HwtxUBbg1YPH24UeEsavRYGEA9L8ADxGNWiinMHdMXPL/YbvYV3HFywsTN6AQ9dk
c5on4R5UUkZJPUzkPktaC2XD1GK4piWSI5ue3tZVmWu7PHMwCsnoSy/bdufwzAd8
jG0z1OLH3OIjQzyo3hUVHY6qPKMbR6FKImte9GCKIFXTMDWSFs7Y4XpgWa3j1MFB
KAzdPBbL+vHJe48yUsb9yeUOhSphRnyprjGBUMtERB8rYGLXt16Lnm3PhNsuuDNV
aDpEUyzu+CuGVFv0+A5AMAB8FDtI7pnTsaUT222VdSJpw0A/OFCy/gw+EeeZ5dcx
XF0TjPGfwLWV6QA6XEcSUUMN+aiwHSMsoeJJD85dQWj7GHvuIb4k+cgdjcAckm5L
fn03UJC1G8CoIO/VVTYxm/sfjcW8VwvUtFvQboL0tYT45t3AJbp50tIzl/SPT5Ev
ftfoA0f2EM7r6JTG7A4ogKhxrum4rhzH34bKApMjDqolpg71MsaeJmIKdYyOpTjO
Fs+TabTchiJoxrVfNyTRPRBul41Y+6W4Kw+DVFF80v+1z2HSj36SqJazegNBrG+q
k2KEKNwIa+mOCgS41TFD2jPJx6+dRm/xLhx9mjTGgjX5GqjCTk3Nz0koWPYeencP
Q3Ex8P+cJK+9fAgTB3KAuik0JqMlaufBk5UGYFKrbZjdtE7TvXP5e7w3PMpPDEal
`protect END_PROTECTED
