`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AEyMWL42E+nXaMrZadlc+wLz23/if01ioWHzR/YuPkADAUzWGeP9GHCmwUtuiKxb
OoGwUEP6A43Q7MzcvTw4xA0GdGPPZaiNgAII/P/a+EACnHRIfsAsYRgZabd73LaH
zMe+ZygIp5egLUAHvfOq7Rmh0JZVI9F7Hi2/erg/STT9vQM2xrKuvSMdAa1X3hfA
af5gi7UjdbXA1S0lhbKoT1IpuW6Xw2PHxnmGSGB1+kgkTf5J8MREULAdPak3otoT
Hs+ZagoeOCKbT0YFIdbgC4G/86anW0dBLvum/rPLLhb1FqmMDqXfTFOdpNAuotju
QGOfNnxpaXaLer4PHZzfpNMc9829BhJC7+9VnKeDfNK1D2hTiKNyApBNWtvlzvLt
OJIatd3ZHHyTqfj6lbCiapmBA+Yn92egSeIS4cyiqUY=
`protect END_PROTECTED
