`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zEXXc9qWLR8A2THjvzf4Am3niKicTjMUrQxmDIb10C1NgLpgX7bEovxM0cy1jTYM
onIRqmUYo3itdarP1pnMebgSytmOUW4pCdqe9+N0aW2CdQz4crFKZHyhzyRaB1hu
KXHmTmiM9tE2yDxh2nt7gDgq3KyvNQx/awep4wJfLNOWKDBFM/xPr1BzLw0K7CIr
6gzBgpzVPIASJ8CCYGGhCbMhmnVwZdod/I5Y7IjtFIBV6bM5F4Xtpnfy43Si45IR
GhiPi2cOPTeuilVrX483eilqlI9Ed0ifzmmDoDmexHmhSJhtX1jMfCxW0UDdLjA0
7FsQfp2/UcPBCytDFED/sJtYeuWfAUB9egVsFkQr6bS8+kWfGA4/SIyGaDkpXJ1l
`protect END_PROTECTED
