`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gTz1yzJNhOFXmWVHOWzxCPaeJTeykqBHKdZ2el15qGFAMnHVmj3/C3AViXS+K2my
QkIEImaP4AIsQE9+FQHAHhO3YTmLWZuVj9AGghjZoMkbqSI6MOwd9t7ne5e+Rdwo
3yhYsyL6TOEK0IzNhPtVVTUaqRH014OwmCuT5n7h/JKY4psXMrqdQACrOsYr8y0g
u3wfJ+rBngvmFxETVVit5QFzw+YRbiJraCo9kmJpcQCVul38Gk37HAGX7eZINSkf
4CtoHZr6SvYzBrzcUatoi9pIwK0f+8CuW1psAuIE7ggQ+YZkjYdD/2MIH5Q9E2z3
vJlITza3qT25lbYq/NUxFfkYXwNkuUT+dIfJSDlU+m/Oz2Uo+eRtves9cnu6oWPe
cnx5gxYeKe3q/+fSuAotm5FcdInaUtV9HJWhcSDzk733Yd+hNjCtkuTGfh+v4ztX
`protect END_PROTECTED
