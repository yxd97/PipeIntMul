`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJCUiFKKaL1bQojBE86avtO3eJbi7U29az+u3d2GlLOuJ0EaYPAP5Yi7XVEUi8Pn
pTu9JJCrZwXU+nklyFzn3db1AYfReC8vRP5FdZwMpTrdUhUemHlUoALQs0KB6BjH
IWjkbnsLH1ZsMCnhWggNCiqt2wD5u/MMitkDAbbLYnBzJhWzAjqt6nPy58bOplUB
eyjAlr+K0PUReQXklyu0S3aaCvWJ+Vpy5ra/VNnLT8JsGrPeYjxI6oWC9uNtxbEJ
BmYuWcLqyywpsLgAkfhIS7f2NfUt0sIvxWe9VXgOA6MG8q/SQCdQtwftKPcE1wBs
CrjZyLySUxVyzqr/O/jAFH0Q3ZEgdF3/wdWarnK50hB8Q/B8GocPOlf3u2kAtYFh
ORxZD2af8Qz9U0LcUc7ImfNq7TDfLp/p/ni531Zsaw3s41bMY96r3yIgasuMfYyG
LJK5z1yuzubphl40Wpwe8o3Ah7RRARmdA8wH4YiR/aOrp6adm0TxX37zihPguDRa
O50J2Q5V8MMo/ZAetYYgmC2NIop4S2H+qRPaoWJ43FWRauLII6i2BCBGfWGJHZbj
`protect END_PROTECTED
