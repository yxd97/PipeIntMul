`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aeT9hpORj579QV/qtmH58KcCHLTVNsl6dzXe2qDiMCpV8KBEhfXPNmmc9uIncPmN
3oXMtivCsL1p0W/UZfkHLJMHQDER7BkPMInEXgdr/1y2SJryeolFWTvWC1BI+I9A
e+qbb1GGjYU/wA0mCmp9PzIFPVV9dECYZdFpKRUX4U/Z3XOAaO3US2cPz+lqDQna
l9f53A99s1s2e+u1b/qg4RwsJEDFJMvC9/O4x02avcwWsujqx9JjNOKBnxWGHQ+e
HqrdDmMZv4xmjqdCNEJ61eF5BssBirc59h71QiMiyda864wiYO2hKwUs/XyKptJy
9p8zenymuT1mZ1al85r8Weft8i+WeEhX4Md5tDpE9+MkQux0inXYhMWUq5Ip2/vq
XsjWEz/h9ZVkg/ixSMShcJ6z8orlCxigEEuwSYPftYP7y89zRqzCluJcziHufIAl
Q8nSmgFcWOUAAU4JznOscyCIOia+cmEup6yO+/hsDsaNZ8T3fSMQy00bV5BCAH7/
5HdlcaU5Wpi+EwT0XaUknJJT75b5+7DCR+pyVSpmhICL/fDVC1E9fXxFK3l1xdRB
PVRHliodAP8xAOc+e37qYHFRc1WgqbDDUVwKULmOWR5MM/QvF8+hfG5rIDHpPvus
zsDZgFIUdXL/yQOm2F+scR3UAcZKqjVmBCx/OCrwMb9vr3HyxVrTqlNorp0MKCHl
bsJBjvDP1SscDy4Pc74Q6amwtG/joG89h0JJFQIfSftU4Ga9z9F8daE1blZr03Fk
luR5nrCxg4IuT0FeOJz1PeUp4A/6YU/Tf+1aYFr86VbiKWAt7xcJ7oU2LaBSqVqT
5NK92ayV6nS3S7+CTW2B7cVMpVKoGwocFFGwnin8ybyvh+WyC45m2onPaL1Ch12u
a2FPDB6SycmCVEFTQoMF7r/webM11apF4KxGyh/vqssWgRb6dHa4gb8c2cjJ1XrH
Gv4+wNwseTMJYWVZVEPBJrclMrE05PDfjXkglduE5qQHk0pi/E0Kndweh/waqKa1
CdfztDGFq+/0R0E2wgrG6Ol3eL+QmEWSmAc9nZq47JAh7/IGDFrJ+OK/am4Q6nKh
olN9aPDvr512fyliz3G/LR8eVwOIeRe5kk5Dqj+MYxEjWfzCxCuc6BrArSi/PPHH
qPxZusUX8H40ticnLzlnmJ1x2heEy8UVvSs0KliiqBi4hdTQSjK5b44BZwOTt6oD
4vGglcScvfT7WWPcoelBNxMusUU/XwOpItufoWPxh0hDBcNZGIk8HWvo2bEoVSE+
eYUQRqaRNTbNdOUJZAVJUbHi3e1LKVSUQbNmaShkk0jCoc4yOpX0aOm6qmRreJT1
q18fZ65tGBrQLxWMzqmCuI/tsMqJLjm6IQOc5xh//HhtziKr5VWxJa+DXmnsidoL
iobaODNSp3pAWbkw7PpgpYGr1OCenpsD175rKipLhFmks3WoJ0NGA2/9JKI7qz27
FPMT5rXqT9HUPm3ptL5Kbt6ILinNOokAyTIpINmq92ORuuNyzqQZBb1zfrAIE08+
p2VwlZHeP+D3i8RUPLg0ii55ru16M9gp1AZmPUZ2oI21l1cwLywHFk1LtsLAvdCk
n7RYbdP0M1kNoQv6D2O+GOxP7SHiMqbDmHmGLRJrz7yJ0lWjBigvrSnAm2L13rGP
e7eKq0CVGBtGFGbx3xvViR2xQMxdX1SigcOJbj2UghZ+slaPwByHafjqDXaxUGCa
/VUcFfbGZwnM0JHQ02UfQU+jbUrymI6fnGQcIkY34QCxTOD7ZflpmGHTxoyS4agt
n4fDdr+YWksfAHac7xlWpH44vUuNFpbSYz7U7yRZRGmwkHklBsM+YGOzzvdLrilJ
pRuqUBL22FV+h6Korf5YwvgbVTZdHP/xcH5pL0mlPNoePbj4zIP9oRz+rtRuxJaC
tqF/t+CvWCEOGVvX5FhXaK0j3NGiSUplWAJprwY5ao07kdoSupcmFEfvKJxAFp0+
lBKeA4hCaqXFsQuP1FJPY4qZRSIeV8TMtq+IvpOOOtVbgI61TuBRtLtCW3tgdp7E
bIo9Kv8JExA6Uta6y/VZY3P1+yzpN+k26yNkuefx2I1TK0qAP3glDxYZ58PIOQ4N
erbiRwLctZffibykcE+339hmvnGck71YJ5TYCX21ytHqx34dBtBrCzKV69ajCCxj
Ebk8o/tHdpFzPX2j/RNo99URst+BvUE+5HPTKAgU0BEuuiyffCvQ54pLLcgd9DDo
ScQdG0qSE7YRhTU/OXCdR4+/evxVjUPd1eDfadUXosqrD2UU05mvfgPDLQ21l3+6
c2iH06ZIEFyAdRdFbwFhgxznE17MyjivgcpOerMnMCxod9efVu5aEcn+JcKAACCu
odvru83drY3f8BKp8mxyY4f50PRnU7LsXGqDLBhxLmMH+B80/xYbTVdlnIqidjxB
e6tL/X5vfKaw/F/6Q8Bq5vZW7fOqLOR//CF8GGabc2Syr1VPR9Q8NmakxF3eijSF
E/54OyO3RUEAunCOyDgVgo61mLF7j2E3CS2ZXbm/ubcW5PdtXLtHPRdZrnmMhDyu
/r/nVQ6ogbT9yt/TtSDB4K3it4PskBIs6PLsVLQUF6qlTqRq3+/oZZ348pskTT81
cVp1pEXUrD+OoQsasuR5z9kDPHn23wtDt1vaGqqC7DlCRIcOKI+T02PfPbW/JrDo
RBcNonu1OMkFLQXLx6AkHiUmuuDNKBzk7haEQfneAqJVNSFtSPrSUMDYL5fj2F5o
VPrmsFgtaYlFqjw4HQ5BN35szNeZNxeBkAVgyJd5Mrb4lQc/W4VM8nFTb3JKrnhS
CgLHhJJo+dTllxUA8its9kUzc5TIOBzzCrpRRU6IYfd1jHhN4rID7D6nxvHqkaIS
TymkOtLShwikrfwUhAXgJhz8mZkNFlw2IlrdsLc4U1FiSffvL7ib0FaHSbQL8ps0
gSnjtmNzP0m0jAoyyeb40neeiBpxR9vdi3Xz5MRZ7QRTioimw2QaHcQZZmopjsfv
mXKaZNiTbsOa2nBb9CVKC+phq9/WBkW2241By8F47lfqltcFtagkJue7KxOBJjg9
W97gYgk0Jasm9dWSSnhU+XcDAr9ocsG8ttCwEuvIHGgFiQm9ngVjqbQ4G9kCpC5c
Q2NU525uq0JKazehzjtklsL5BzEliN+3xYiY6YWSZIKqC+GlrtDCv9mjcP5+IWwm
6I1Cu2NVklFEsI19Xd15tjuy44UpLpWYN9IsbOOBl90D70sgu76sCZBRK0xxLuux
LPsYScN8p2BITtxy3wqDd2/mAgQ8OhN7qbqc1HjzDkanIhG5/FoL+PN0rTydENJm
K2wwb+pf/jxneGProJ0fY+N1tf/pCcFIM0H/Ca0FNF8Ed1A5iNabslfynoyHmHIV
zZgexZ9mYND273NiEgxP5wf+zhiS8GTpwUEfhoQ/nP+DhFc+eQftkzpXzyyFiSYB
EmJxKvdLMI9drIXafRK6fBT+O9RQVdWO46fKGTm0/79Z56FxB1KqK1UVtLW92shH
Vk/N/bnU1PXBpCEGHttjtteXlzK8PFwjqXhRrvPcfWHEHJ6Tfx6/pD26U+FLL/RN
+TSFU2q7jDAuniDwXwporcA/H/e6TY5O+HIldVDgRot3zd70UJwQ1CR4yx5L8+KU
SKMBsIZdq5wq1PJkBrGr2opRsPc+eN517oCrVfPCeWesMzzd641/5TOlpBstjo6H
KhCxsdCXln0bU0sRx+790l/sdsghVgOwAez7FXMqKu1z5Z7WO2Aq/Nq/6EDaFUK8
autraQC9Fl8nxyALOsi96STgHIEpboJSZ9NpARkWCh8qFwzfQV3cfeh98LsImWxq
mUpCvTf6pE/fWhHMv9ud+2IPcpov07/A4pq/NBwbW1soCsLnm1x8VI79SlDsXCLl
6kULIb2OCp8JyQYEr4Mmt4G4nmw6mUtzLIdH9tuiwzqWZHywo3cCuB6vXxVc76D1
2pYcdyq/6/U+E5dzzmq/VKvhxIEcMuE/4QYvM85Lt8l49PCyWjZCD4bT8Ypjicbb
xU0wxsahOrsISe/FvCzTyrYVP92GwPWfgTcVWIY2L32uiVXYRSRxaHO4M1+8Jcha
ddySyl8My+lFr83N766ZBwK1WkqJEb/n6eE3V6tr27eCfG7+Lp4yDZeKj6KXnoxC
gzxgKxu5YnxiqB6oUEpzAlpiXv6iiH/dzTfjITHJAQpkU0A4XiHbsBsVOI8YCPv5
m5OeCQXoDIIAabRmHjYdvHQer1x+3rqqArHIhfl5W6K9czl6tdF361DIw7CX+sBz
wArDyej+Hk4n9N5USiEqhBxsk5gaFB4/JTFm+5c+t4HBSF0wsFB/fNh8imErG1ri
L9Ecpzq+RJy+Dxu+ua3I73lupq1BvqdAy9/8GdOA1ZEHvdhNNG/vhNqVcQEIXFag
Iem9YjSbl/K/9N6B/YT/A3p33jLDVUtHEvLcD/4NfEu7RaxnT04BkUy6W4RE0z/r
zP5t0D2QRjK1hyF1ykTWB6ZeCxgTYvVrKyCvlKth2BKryCLaHg7PBK/Rezdcrw0v
5f2YQ1xsxXn/0Sm9iqKmRHGcKAIBKGU0Ucem3IcngOS+gC60nkucz1y72+zENYd5
9ru2vgy2IE/Xbh34wfsB9/inpWIXvUsmLbnIcURNPSmjtgYM6Y7uNtYnCAkQjZxL
GWdCklHcTMKB40yoiQRTGEZh6kb0KFABdn2uyaXI0cLDYQb0R2amQX5T1LBABoQ0
V/ksR/Af8LXPjNPc8IwPY/y+AmfS+2XZSTKtrU4xdKgPnjJb1U19MimolHqodr64
UkRFFkKDAqq9Irm98UW2oLvidMw0oLZkDyjXdEaLmJI8Ew/hMoaTltwJJIMIn1dw
fWSJYwoXwkLeqidhwxYJTXFetUD73oS/pTcNZVWXmFq6CfsWqiszbJej0+91SxQg
P/qNQ4xZ2jS2C2CARCfquPP8mke4eF4KS+FLu39hwR/SRIZVgmZk2v8sxPmQ0F+5
sXs+kN6R2A+1d7oQJy2fp5H6zB3e4+Y+7cJ/0NCi0gk=
`protect END_PROTECTED
