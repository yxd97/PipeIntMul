`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qj16WI0/OD/HIZlWcIk4ycIiavyhjd8iMoT8jpctDEbPIsGiR+QBFV5WRfT9A+dh
nkbnOZeR1m86gAz32o39FTwWuiFyIx/ymaE2Tgqy5dGAUHlQiNqC9Ypd7gyW5xbI
j1OvISYhEbILdDbVun24Men7J06oJQPGaEGJu+tecfsjOVM6f7RqsKvgPrcuxcrX
TZpDdJmR86vaLPouErRgEzOS8h3dhQxll7Jh/KToPFH2BxzvB2A3PPioJ0WFiNZd
6c4fHCz1ThlzWxPC3mpiN8rGTQy2aUZyal7hKezwXippEtjthaCv2HrS7/WveKjL
LzAgBPZB1bNyZnKg7RsoAsj0C4YmfT78YetaoBQL9RaKWpn+ZnkhJbbrZRtVYA7M
Hws+L8QdXAtnn6XAsnf89i+mz93fdHLTSzxu1AmMTeihLoLB3pZtiWsRnkVQy9t9
6E13J5RuiZvBpRdMprVPs4TA65vELywJzRuDaNVwGyIfdCQRcpfoMEYK/asevVIl
cls1ou/O71GudWVfDHq/HKxgA7JrNrTGnFki7ZY7TQckc5o06NU7xYHNguysHomL
2L1QGg+q5WRIrfm+0MAW59Aa8MvptgkV03U/ZhA5yRniJaeIW/cHRcpIyEyNqNqX
RfGQxSWXDVWk7hqc7SfMYd3NYZ1zMl4nsouqo29kiPZ3u279mtx/orBEoYo3hiQ2
DVO5l2+4FM4t2DvFDOnJLwmBnO6s4UFQJMkRV6N6Jj9w1MXFpKvKwE1apVREEisr
XAzIqxBYur1jQ+woNMNNj26VIMhhUjIVj1GObxLsEDA9wMFIaIVhtdMzScLRG9tq
Ewrb+GHm3TPFbl76kpGajU9Pp1ttHwEJInaJLNM166ZcDTognB/KPEMd1rhlK5Ke
Ae6WoU2wCccgY/jSKxlAsC6GHYKjBVgpVEM+17HM0U17jlOzOCdiDimOR8NxogD4
`protect END_PROTECTED
