`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v8H2Q/xuRrULo3GDb3RXFKZ3HX5BfTSCKUaQQ7n/tOqeg9Ly6gkHNRjQ1ysvkW7O
e2iFGzOqPbBB7Lv3ssOpDPWkOStDslGKfTysz7bnvRsjaRoPPRrW6kWKVnZMB/pQ
JNLJJCp9+Dl0ENnBQlHlmgx+Tcjzc5tr5Py2UBrTHuvRMxJaPRqNQTVfbjM/ZwXc
wk3Lof8t9HP2RjBkrb1zAtOv0NryMpvDKPgGq74K5YqfwlZaWhN9DPLEtIgmw0AO
BQ+0NJeDmH0SsD9Gxo+ZETqN/THwUgNvbfth60N4neViLieRLq+GfhQ/cvoNOaDQ
2rvG36DVlslSKJedvh13YorhqB1JMq1Hs26IJBTAknoVd3uUoUj3+ZRQsaKM5S8P
/h3FOjR6VMu1n1TMc6iautNVuwxW6Or6P7QBRiAlblWrWDHoZdENXoswPP2cB1YX
DpYICHzmdnPjIhzTI4gPFdNkb3KhXNoH1nvC6LdF7SnXHeMR3aBANtULlh6+yxwQ
PQ5qouM7cjWZvd/zepBNTvR5qRC8m2pwz1asxsBVqlJph/LXh92bba6QyYAsAF+t
ClquNsEo39cFjFlm7oPLSYHFfEF54NDV9sUH+cxcWhfiBWoenX9RCRWwDjktE7CC
Rkafrx/snG23TlPdTLF4uIMJbvlN9z4ATLjDQ3kSeHBHyZXY+8W7rqegyBhxPF0V
wo7Kwe+L5zm1RqfgF94IE7C440pLx8aiKQe7ottr+AaOlBiIW+5t9T5ZaS3FA/M8
4Qa39HTWFP/J5axgAagGPymHN2sVhBWN1M2ZP7YvJLxQLRvJCghfnzaunzp7/fcF
Lk7v+iJp/7gsNgg7AfCf8KpMmUsmrclJd4Q6L3yPrfSPq4olVLQ+D8yI15+Uxv9A
AsmuyLuyAAy2R/jMgNAz3ImPDm6XTMMuEWD2RYtJL0gjs9ET8FyNLlFdC+IXsA6L
z560lUAnr+mKElfOeTQZ9DCMDIhr8cnPcVnn1+P+IyhYdaYOwL57gX0/163FPncf
KEj/zzAxzT9dHOU94fGiKH3KxrDdWZe0WwGJ789cYDikL5F35xMm3MaSddEGTBJ9
vM5AeZdFqG7d/nUEUtGt/gZ3DWkQgyxuDhj+YLXwXkz37sK2KRkFZFF8NVhXlcyh
ii1lcGcKCbTnA8PTIu5yaNmUmrsK4ZonBtXaUiHKDalGSNV8Surd6yBLnn4eShJq
uL2SI5naaDAuZXPEKuf6jiOnVSa2uAtGluKGQHmtxt6pootVYP61jH7Vk1b0LOgG
Mbn3IXUWh7HBC/tWD2GRru72ZLFwpESoioSZzryt0s6AhDq97oH/gXNYXCD6lC+L
k/6Dyrszv51UB7VyPfTgAE+Nrq3BFwdO1fLY8JdTpmLgAEu/eGk4QME0Jm+gPTkF
6Gd2GMb57QHUYxEzc8FBaLENnt2nf3exWDzwRUj0JG6vDSS5V+/ve4J+DSmICJQ9
b4i3ovrwCQTJJlP/8eU/4BQezk5zfghj27rl5cm5wiybyMKJHPdbVZ3RAw3lkapr
HNoJtJSg5GskCukDgcWzwyMO8oOPhpULEpLDSRYIPh2PjSXZ+IHrr5YDUmRdONoq
PGKHDF63kmLDTv8SVW985vHPKKfCMeY9WyDrJspSUMsnP4v0xA7kZaYoU9Ao0rEm
lfiHO+WViH+UlSCELzBBjyvXUIdq5CIP9J7qhyiaKZd0dhu0oitCbxUsa9xtUYkP
e2PMLbgxS4YV3lp+4JhN/7Pq1UUp0TxTUJh+jYWJJuNXc1oNsPWgTMlC10a3PUBx
y5hJEFRO8FmMeLVkvmeLP4IhQupanj5jRvhHGcrYdh8FCUWmBaa8Mzj+emCwvPFd
d85gCLIwV8kIITEjzBalKfMlZZ7xBD0GohQJfpvzzJPrTXVdGpIeMOQluA3mR0o1
zj31h3Sc1DJLfe9EsNtYIKhJQ2vrpTjj0CDO2gUTEm96YcxhmycjIljnG1Kd06no
W6LQI70vYbxY4UaivyGPAmo4BHozDvYyfM+LM9MN+AxFK+xu3qEDrCkPM+gcf04i
tbpojZ2Hu+5sOvLiBPvePbTWVJPXZfEPS7nWZfzOTibgyBs0nX+5bwq2PCZIUVP1
SoCcILjANSb5j6kofSmNbZ6IjT+8ryVXkQJKUJcErnleGrdSYYlDwTW3L93GrLdD
Zh54AJ0/i2M4bSgQzq217X37QNmlrtzDfXZklyWjBscfBJsL4U3QSmK18ppid5tm
vcBnMn2G3umzH59KpFCWDdqVXDsntkR7RuTnpXqnsONJG1Hlz9Is9UHW54RRPPOj
zl6dLKf9zbd++FEaFjqK4ga49JYv9De/ebzy5dmFn3b9RVWC2ci7oiHBI4lxnnk/
`protect END_PROTECTED
