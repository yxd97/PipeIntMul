`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQhCjtHX/E1mWzsfqsj7X/vl5Kn79zkCbNdD2qS4Lbx/e4Epn28MqUSs9grT9f9A
h77qpYLrEaj9kip/5NnOU9yvSIw6gor9oUhNyt0krIavG4aVFZFbLkW/A8r8zLtS
K30nBHwlrFwSmES1/KGHFkLW+JeX1bCb0lXHZO1c9uUmiwxyL4gDx+e/UK3EbPz9
IW/u2nYsLG0GC/WznSUeOByTPT7sEmuwTdz2MA7DFN1xUT+/facxT0YlYUDo+orE
zwuipnnvqK8ilgCVWFLO+LW0U/u+0ASqsHx9A3Vo6qDEXCTY2SRkANOHsII+OVWR
UG1LsabM0Sp9u88RMMRYh9dCJUqEXIaxKHpM/U51B/4zMCn0rdSHv9w3ROGPA97O
0OmF5SFKZaYPD1G4bFrsvE6q9atDRDKHhJYcj6O+LCq6X1fzwb+dXS1j6dotQDyk
HKcpZ6+HSi/4/nt7OYWtCEzmKYCI2K2a+bKNHQlM1xBQ5TAkvS56AWzSpxwM2Wjd
sIm32cm+PdXarURk+30XWbAFghJ8UMB+vQTTwkyUPCYRJH3J6nbqNhGDumOR4gwn
N8lPTOd5FDpZojn3JpkpDcQb2or6SMjaejK2IuGYWzPsHQv7MChvoLp3wb8s1XgC
`protect END_PROTECTED
