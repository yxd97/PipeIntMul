`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cPi6+BhFgrfOm30JqLskfuYRxo2idcoN4tVvS1oN2P+kL7tPno1fFEHOM9eWMV9s
df3jYsD3qB7SfWrG5oxEyL+yyrns5QOkLG8iHMrZoAJfNJRe1E0UVOFA6WchOP+Q
3tbpU+oth/CV6hpRF7hHEsGAQ0jZFkutUXUHso2XqDptFlg2bcR0K6AHBrYcerXx
KUbHANNZXgfkLm6SAabxl/VEkffsqv+hDlUDcxoU2PBpKL/NTJEsqlqqhBWs/YND
dyn00GibwTt/SwWMtliAzSd1WzVsoe13XtkCR3O/xFeR+7PRpUNCDbnCjPn/5Xul
ydztAtN4opiogTxoiSgGooGT91D819D4j9vCaIJHlik8wOQermlveI95nqoP3A7a
x4b8aOhz0tzGe+yT0K9nXQjXWyEGG9r3rpjbeJ0tO1MUSKWCz7c6YF+D5xeCNcNy
igqfTEJmtsYrKHcEtGWFklyaane5lC+551ilVO/7Jkwpnwio9XZLCQyalk4lfzwl
bIjBg+l7R4f2GcT5nhoGVA==
`protect END_PROTECTED
