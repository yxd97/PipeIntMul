`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0e43N1MQcsrks7ewX8BmKhjVUoO5nNqzBhrAY982OhFIa9pyYQi4oKc22PR/Ji/
25Ws0jeECnqnVgDgrfuIWSfv0rkP2aSixMhbwxhzVguXcFOqLu1B7W/NxtGQpcV6
yx3Os08NJAJ4ZmgGhnduxQxkXi6mEmV9Wyk6v7T/6ylAtqmqrrg84z7N3c61zPNc
V39bk/6TRZfoRYvDmWQofnY0nj+iciId8MBfFXsrQYgh23DyzMaH/HmgsxLYLEkU
+m4wvW2gfIM9Utabwv+qiy58ZrTv+yfwhrPDLBws9rchPOtj3Wli+T+GT+G3eHIc
d+AcEuWYiaHZdzxV5BK53TNpatQx3A8VHVG1lsVgE3StFpjQMOx7bRHUl5zIAGRt
/Efy9ZwbsPfo0IVWfcAkxWB2OJreEBsNiXxN79EDdueyKMKi2o+P7f62/DL35CYW
/tg8EcgLyRorovd6lowDmbUuIJ5ic/2tUJ2YGZkAQMDyOsTcwCfzpXoKl2UHFeN6
0iFU9BgjEERFYMwkt5j84pLCK8Hduv+YUjCZJDnHLNhHMi8zaYBCpOqniWi8RSMl
nUTy2X4shjxzCfyht4TEwA==
`protect END_PROTECTED
