`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7YJE5bcW3aV+pN5A26zNBTqzmirCrGjKloWQRCBUtbAFwXsZS+dj0nzhaRo9SeG
2/sjN8RJknM9grc6d8MzvEQv9L8LxC2I+Mq/+lRhHS1eBIw5A1IMSIpxTg3w718y
lEL7/sBCvILOMPkmt9WzrVpBrVh2WnK2Z2FhyuQAdFLvYqHD7bskcuByQGSZjtWN
Wdx/zDfrNfbHTpidnYbP3TQXLpObcmdstNIaywOmhbxcRKckOg+hpq9FKIAgYahy
FGqgsIHHqGkx3MpvMoQOgOBoqi4wDu1NKQvWR3lKhuPTPZH/vWT2sSWKioUUVm0c
UbkT02z/9axv2AVYY+d0YofDxxxzejH90dW3qxsipKuGUYbGIJyE3MP4xlF1a1lv
`protect END_PROTECTED
