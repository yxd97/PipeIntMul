`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0KhCY6UtBRZuqeVtlNqxK8mPbPfogFRuXyFRFr3d2JnEVnztXTqlNH2YW3lxyMSj
tVEI7RAorrwxFM3OhtyZuSUPPHVQZrukKlcVfXNsbo7gnOC/MvzzgVlwHyXyNLpT
BmYnmTr1M8yXWV+pgQ8Oj//g72HhQxCYeH7wNM9ywbCuip++vCd1/jULRXvEgA+t
5av05sXoh3VgmH6KZfy8d7UtI5BV0GNwVbcsmrR5TCOlXlh5cKYGxbdmHQO3DfJl
Xnhw6B13pW5PXr8iszG25JMm7dJ0tpX2JAAlYAhNiIaR68Pfq49IZC7SJvA0Yj1E
kndZdxbJC3ojv0ImN2bLZDeB2gjcbCsm91Us8bTGXFOJRpYTK+bw39krTObV+Ft6
Gqv1XtUWTkOoFoVzaG/zjkul5e6BxoN7Je80jWgt99onQZU4DI+/JdTrEuyF0vyx
a7atKIDlzQ470qTkv6+UEesDN10a8CSfqMo93O0w/4jpxlmkkZFehbNCTc5F7crP
uYLEKBV3QD5HuEqKPdxqeTNEsf4BSZ0mbii19XyRW+1nUBNfmI5zWlub1fu8e29l
gzfRFhGoqMmr6bld/hqZFJmp1Q7T/W04nnePmqwYTxN441PI7dE9rNQYwdADsUmo
vnSB+TWT1rPRXD18S/0Z4QFQrHrcS/hzBFax11cMSQMqCblkKMI1aRw0qGk/GlnJ
23OgnSNaiFCfLVHdaJZfMGaZ44BK6dWVt/AbpK4cE6dAkwpxmxjRSTEDRrdJu5YH
/3adqNuDaeXEB5fTmiqGDkFGjEUGnP74QghAHL3/OFVXvMjnm82SXCtqMVWYvxC4
rLScv6ROdXRha5RH+qLQsg==
`protect END_PROTECTED
