`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOFvtyYFi8g1s+sJ5sFzQxrNurout21xeJQslaLEzv08bLbib3aeWR0lnjIvThx3
PwzUF9Kg2dsJVxMO4fDBUR4hYlnc3GU/37RxA92ezILFHxqM/0MWiDOxEyofBtd2
LHsWpwud4y9DmU9wJicNvB5KyqcpFaX/ccJ8E9Dihwno9x4M1cq+IN59MLIUat3k
rbca17bOfxkGEZEHXvDXpS8miW5w7iRk2w+UA2fsPu4AUN9xbCuDq2iVtB0l5tcX
Wb6ggKKsTZPlmI++czSn1q2AXY++4k6Iw5BQCUjCX5lFaPAS/IEl1Q62To31iJD3
I0+V3gX8wm+rj/jma3zB0v29vPtulc9IUC8+OQMyzos=
`protect END_PROTECTED
