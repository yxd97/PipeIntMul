`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x395dnXkOfGF82xSIIicYHDgmZqtO4GFyjnpyyL8R4hTwWQz2HrJLHwnqV7OTbW0
GWgZAFWVBttIttPdtaiT+9apWTjiLc/b+Aqk11lJzmi4NOAgfztAlu/FOeiHFd7B
fwsqnRYM9NPdGVw3gdmCrjvPVhw+NXWNFBuFVwz5U8oymJ+jCvEMMLyo5wXARHJr
KrM8WpPLKw/pL/niYywSSroKlfnN6JiXCFRrbPsc8INTEQzZcX+omys6RJQ5+07a
yQh8B+/k3ttStawWatg+BcUdRDc4vDd+nm0IzUzoIILJJdzDPPQ+QxAliMh8/c8P
fwoovubRa68qIj0+0VtlQKAI64KPzsv6A3i2r7BJuamkmrAQ1VBKwaAuRMVjC3Qj
SDtWLqEjnsaqgNTNnLIFCHK1BpHbEUGH1/Xvp7ifH7FWFiQp+bT67YHa1eOm+n4e
WfCZKntj4u9vB4addMD/FMrtB5rDWdunOGt9+8/IvJg=
`protect END_PROTECTED
