`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85Mkb94f8BEeYr1HyWS39Bm88S9umyPIWnFJT/7xtpPIdn8LaoZslacn+Rm/NTOJ
eyA8+n4gfv4AWUb/Hv/rDmPt7W1X0gDw+nlYb5w8jzQfpitS3aFBLvbXulfQaoIn
cyEvyXDtBz2Zy3UnojfCSVdjzXzKId86tgIHVmwm4DxZVauyoFIFIt5LrJ2/okHc
4gbFhWMWywjIhuvsMtNlmzZq/HQWJ0H11uBb6wnzlE7Nyaz2/l92JngDcHoguYdx
CRcZ4TdkwhIqQCMZwwvI1Qiq+exGebeVABXx/DirPnNd4IPKxAh5kUthNV+JSDgw
3aqB6KGk40wMgPyu098jNBBCuNa2IvonAtMSlM1gY9Dw8pWZw6vX4UlJR/4P7pxR
LgbZIedzz6YThdXFcPfDyPL8qDX3qSiqRBGYODriP/YtQxUtQw3Zk23/aYa0BnNT
sELvP5nz44XIeuQ2shmyEaoXYeFjOaF7xvThJkh+vGF0/f23cWGYuoMUGnv91PmN
liPeGwLGHdceVYWaAIKfqRWH+b1PcpadOGqV1XC+r9EbmKrkA8f6ep+KkxzQeoyk
o9Z4M0ukrkB+W/xHuudoIefC8WJ/n1leywQj3kbaW8jMEp5PuSZlCGBYIuZ0R45X
Ypoz6WxKh8CLzQsxXtiVGqt+cvX4912EvsQJY4if0UIt2kKkzI4sqhvkISTAfQsz
LDQpslu0LEljw36qEbQWqDI6G5BC6fK9rdhgJK9mmrTz67rELh5reYsspb0iiVHo
bYdWa/SkgIeokSQ+kbeiBpI/ef66enDxR0hic+AnyrJ7P780NS3kbV5ev0h+YGxQ
en+0+zhEad8D2N4GqWcTj1XjI/dDGIoYRlMBF/M0b969fWDS46WjDAmRWxC7gylD
FWW2x6UmZ5IFCaqpUZ9OCvUcWflG+oOE/0CILGLJkjWABu4tybFfVAKgLq7HfzlX
QiV0oiltCsakZF1e/fZ+DRL/1d/6U2UasR6hUYpIb+LPcjSNJSoo+ibBjua7XfHK
`protect END_PROTECTED
