`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4E46RFmAziLX5CLB6kSHgECqZvZIqcL+lb7en5PPgl7oHaKgNHYATwgxAKZTEzE
sM9bsnluNXxR+3Naze3mZgOdxDQiiBNO/VgJPMRBev3on/QEQzIsUJsB7nHGf4E5
h5qtv41LqI/sQgC5Kjo4xZiE91bl6wuO9mm3DoeSmpeCperHVqSsl02sTFbrxR36
Ms0c4MnH0PYqbndURDCclbMU85fyqJ/CEppCOq+Ysa3KQtng+zG1gTbZGaUUxXbr
IAohCnayLZk2LL1D+L7+jQ==
`protect END_PROTECTED
