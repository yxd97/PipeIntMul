`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcL1uBt3PUp1iZh8rM+9B5XgWNgsxdI/QjIXrAhdpDffhJ2BLfwhHaEzWURAqtjB
s220tS+O7ls0yn+dznwfR3wNxVyX/bK5Uby9AQFyENbCdCUQowtsbfMvGJE0tgga
KPmupSSAVZMS57muRLdVDkUlBRSNn40tvOjIClbxRPf/S5A+v0PwvsjDBKJnvJEd
axgFVfRovn7D7bjzKcpxOxbt3yAKJK8mesBr1OjWA43WV1+7uUxnxYY8fWj25IRr
M96rw2knFIWDsPu1pRV1M2lpxoGuXi5tuWCIS16bGv4KktznSZ08nTrKQ6ortEtS
`protect END_PROTECTED
