`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t4sXA6PisoK/MD7R9hWD1L6Jg6ASuCk/HMlSmKaqWW7IAFP4zPbuXGgB+b/g6WW3
cfho79gPDFyVjJDCb+RISoBWpc9xbt26rCgUb1H/Af35pZkCAk/A/xN3Pth5q4Va
IgMR6w+RTagPMPg56ex+majWE+9ODuVjkYJ3nZGWLCI8vsjPm+goP51lg01sgPSY
rg4ZidjHjW8/IKZiK+LAldi7SpioPvHOuBS7UF36vh2zvEeCp/N/GWJEmNasKMDK
A14PRkmC7T12W2bL6fHHIg4Eu897Bpnt1TIhvRZmTq9rl5DkBOzBRSFCV1q0czee
X1j259pMZKhX3cBPvgJ54g==
`protect END_PROTECTED
