`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UVfQMrpn8bZigK+pJuFpDfr43WoeJqU+72TEcvVrdBXLMSQJexlsdF8dq8hKbOm8
ioSw9BF8Pf7JmFHMmWITa7eq2OqKe00GcItC3LUhzkNL+xMA0PSPWlhYlxovRiYZ
mfrqQrYtSVAH2tFacm52zIywCenRrM0O8xHCgweQfHNUcOzOIVX21JBrNCJWJLa7
qPN9MmGfIvFI+yOqrisfNC+lRHqE/ru/mUv0jTB6kot89vvLPKJjmMfVHjdlOizn
W6rl8xWovAz6L5OmpscwPFBvhADTTNgC/Zv3i/1VpEZKJFa98o4eyfSwdL3CVPzL
`protect END_PROTECTED
