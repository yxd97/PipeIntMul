`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6M8tuhOISRzRcFm4lM0CSwziwI8D2DLLDgZ1ilFwTwoqFDjzvtz6Mj4Wnq7I8f0
tKJTBIsfxyHAK54YbynjSChHDQe72B5PP2bi8ry0JBcFD/l1ThWRYCx5ItHonhnJ
LM/NcyifDFziLWXmBbNBYK/E3Hkcg91L6L08iQmeLmOy6ebQn4o5y6tFauE0p3Y2
sQ+lBEFGJFQuc+HQpyhuSiiabkzhEBIp5r8IMP+uNN3G2nYzuOawwwtGX0+NM5oC
dwol1e6zIDITf4SIIMJdRsInWC4KN/pRNfAe4ojYkaHOKr0z6Kk5fWkxCbOV/uic
PRsoHcPopawpmc2YPqDKLvG6GRc+r7MG43TJKnTF6yxqy3ZM0hFlaHk2WKKdXGrW
JOAjNh6dhztHt5JZTqlWEYs+4KULRHXAo+xfkDQN31Bm64OIuE9tQpeqUKRHMrhN
0cWyqADpEJH1wZzPMfWoH6b5DxWZLbvpojjSSMqRK3Y/+T/5rZOgXKQOE1tYt1pQ
9VNHBUpqrL1PeszAln8vISWkvERVosxdjseL5hAbenchF8QTNOHYl4JGka1pMB2y
NbRLLDzG3fMltJhPxKFop4j4mQJ/OZvyMLIqw4fQQuTQqaLEAQEN/0bbjujfakbI
zYjoN/34jMk03TIGhS/5ZH/RTWJWtLZUdnC079wzUPiXr6DfSbN9OfQUd81k56y7
xpwyLm4cjPd9HuNQ4s5SuzkwjWSpl3gVxmX938NVLEeCJAeTJunxMzVqt7+W3fns
effpcECUHWobXRrc8JDanlty+l+0uG6xD94AGIWE6BqtQOMjOOwwxxFwvhDrSCyv
nMkO2fVqRQM28ozH72eDVgymYc4g2NKSFm0qpH/haKnGgfuOffKIQUSU5sWJyr3M
AZQI+r9yPVbrvWQvZtT8lXOc32qpUKre1OU5G0uqgKAtoyMXShxUp3tJs3/r73kC
dHazybUTpjKMDv245FnZiQw4ueyugzezKKLg1jkj7rh/EA7wis8Lm9RdnnO8sBWJ
mqNZVKeFR6+4U5RTU+TRyNjY8bdD8TNGzajxEkBSzTm0bSvZuXUaM0re/5Q1T7jn
1hR0RVTmZkB51FVE01hGOkPKEqJsOHRACa0tJFwU/s8me6sqQd7wekqGiuGgLSf+
oOvHVcFdxD7LbvtGBXGcz/aPT5iLodU+vYGxN5nysaly7LV0ZIV9hFONoIhfn9Z2
KeEpSO5jaS1ZmTumtIUGKUXyiqKDj+Eu8H22xoq0w6vLHekadLIu+97Q3XqeAlmn
3V4L8ZvutA8z3PgjPsO/A+gj8DOzKiNMVu3Dk845JJQlkURzW6FBp4Cx/1sRB5Ye
/xYjcjkAYC2h8PFOFBkIR7C8I9NU9d4mc8TsAobzym1JV8swHlgDNlFfBusJm5V9
+nylgOQolwRFG4DQA/aLAXFO+QAHBoboWQItrj7Zup7U/UUYaVWgsC+Pkg67qvUk
uiS1uAFq0s1OKg+Gg0VF6N70fjUrlZVJgLs9e/kHmKWZIr3AypI2z6QcwqrLmI8x
fM1VmQsMhR3xz101GLqkW8jRnlxGfbkLEmN3dbXLlIb2w4rWC9xyEZp1ma5gB1LY
ZA5ujuNQMf9f2Z5d1VKjBAqKKTVzqXTCOvvMwXpiUU7+ShMNFrf+tOnTSciXz5RI
jqwUR/TsPYB7CJz4PLlOEuhUfmDfzlbROVi7C6Es2NTGEwbo99mTylSTfNgkeCNL
vITvlJ2ZgurVvHg2K5RjszbftTkNoX1Asd802A04kepPhEWR9AaxC0K3RrsxPvzc
X9hgmyHtJvZgbWLwjzqIJs+nJaSC+NwzzE3tEBHinG4PJ/alNwTRBtjR0N7ZdYSq
0OlozjdGDMtgzbOIULgLbuUSYLhzXlkcT18O5+oxjLDnlZrZdjFd9tawuVOz6WHN
I1GzJCaMF6TKb1JSeBH3dMwF+0NyzyKpf5KpEdNShraqUjr6+is/Eb2ZRf5U3quS
cSsVpcgwMYo2Rr5Qo9Rbunnf4fPEzHyDjLS8AZYsQ3m4ymj+KgDfUF/mZKSg+zF6
BvdsDp1HhhJoISAnRm6ZKG5GeMjLyNKsZUXHkTl/C7HI6sQkbd4QD7JRK25twHBS
ZUewbgUxo36n9BaJ+uHp7bv6AhaLENprTeYs8aD1F7xGL/d/i2a2+Ipj/GNxeiOz
7SERwmSa9NcUpdOoxEzweZ5DzkQKy1weAQxzbgvrd4YI7a5Kl2IwQRx12KgsYwQD
gBxrKm03e4WcXVpH+PntmRZ9P0D4A0IYzs0KkZn6mbvdxHR4TnjFs6Di60nY7kv6
gjyBHgALBz5kFXupNurOhPhtQv64fgXdh5qwitbWH+h0oj5eCUatYp8K6lCoGbGt
nYv2TknnOPDqQH+dIioyJiazKQTzu0e+wwx4OVZ3rKaU+DqpDDVO19HGAn8wPF+H
sHwCWqlni8eblFKselrf4CLXmuT6X6WGPvTc1h8McU0wb2PpdCNmgTz+v1R4ydsF
L+TxJdJdWns+qqTVaKQelJBx9ykMqAiUqSr3szTd30ruHYdPVAx2sMPuzDdDtVSo
m2uNoOqHLFHW64CIfLr63YCtgB4J2efsbVfe2ewfBt2Yv0QyrlOh2e6xaEHjU7Ku
M5F5kncofpd3I8VOeqCvINivGdZYCrEb9xyQRB1WJThbn6MBg9XmiINBwbdRuj3o
4moBAjq9h2X5ZDkubdy+VGVKVodp+Jod0Cc2OEVKRIz0nuT6F0sdQxFkDXXcrWr0
I7pEJE+dKhM49t7wvjuy41WdKXew5nEIj1zycNd/7eCsIf7lHxLeB4pywESwocaS
t5FnJUgjHT+Qbr7FJKGICvyg1zMmJSIgxTlA6GXz3XI=
`protect END_PROTECTED
