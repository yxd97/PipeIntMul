`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UrQadwITLLob9kFfQhNJ8B+f5SITab4kU+5BVtUe75EeqcJ8GbfR5V2sDh+UMEv9
cimpR+eQ7/0oYBn3JD33BQUfbnMPN9IqD6vmCWX4ePZ5mo9jfOssen556RO7UTNx
yHtRF2YITbiQyOJIYqhdKKFk7G0gABzjZDj1u9qP1teZAy7WYbJuRrcmIjR8kPlJ
1E79x7esiu0odT1rGJ+70+IuXsOY+OTCoZwsjOyXfKqeW4+X1x2r7eVL41MulDoY
DBz9yEXAyBpXkErbHj6GCntkWM/uOids4XY/WoIhF+bQWfpZgatNX62Ag1tFFUHS
zgRjQ35WhV4KbVNPNJKFcP35bAV+6fdw84FIw/EjjgJAZx+PBsX98MtdCk8Ltijr
IE8KYA7feuPjquxJA+VWlYL0vzoXWdbu9COpYNPXOw/Tx+DTyC+E0LuQuUm4xzlJ
ktXmZJ3oRR306DYV8ORSw+UCgylG8eEq9lD6+uUzAkAsC35s704kccSfs+YATm+H
Pejf2+seXcQNh0sSCandRqFSqfQ3eh9PNyQO/XLsDYU=
`protect END_PROTECTED
