`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WS2QdSWgs/5xwbvdoLjrEz4sF+mlLFr1eOGVkdUxgYRcuLQkJ8GgthGLWl8EHj3Z
2WboVWnhvGtrht9frIRDAH8WIc8lE2hM92pukOMd8eEdw0KJzo5G3CSLOJoAQgn9
tSZMnm+mjcAT6875RCATdq5D1VXPjtmI21wIDxalSm/S6IMplH2jAtozfSjXK/9P
0/X8tyyPCL3KFaiCtwO4FY1nQ7S9CEgVW28UYe9UsakKMMvogr8BsYUJqVWe4Spi
ffwl+cv9ArsYHtXStTvH0gzqFz4P2Ur3viokqspJhfwKV8h4/0FNHz5EKNYtHmRH
lqJPujGloAuBQjmFtjgIoJGeAMe1RJ1EC4Z/3vuxu1SKX5hawvN7BW5wiF3lkqV6
TuB+YHj1aqUj81Vv+Z1KOBtSPaqFZKGsUFl5Y/e41moXpCWO2ATwrpbSENS6FoVv
Fr1Lzo8EOs9vrFk/4ZJKA5grftxQ1hCcRuOLszEWlPnMDDRIQZGKcx3vIevw+0PL
yihUsq4o03o0kCuzQszB8In6YxRFxPPdSQQTcP9xnrzug29/+c2Qkknvdnz3YKry
+XvJs5rSO4lQb+2dy/nCaocZtdT5z6wycKwEk5Zp64N6yqfBefWOZLZJU84VVC3z
5KCf91deFZRTETKAuI4Y9PPchHT5srrTNeqIR6k4HHXpXpkLbtc8iqoJiEznPZrh
YFLrebqARUPGGjyMa7sojWeJcafBoIuGfKEbjcV21m0VI00/FWQ2AEiFwemNZReO
LdE++MDmpdi9yIYcaVYssYeQpET0lrHazWFUlX++5KNpH7yRPxZNtfDkMc/8QRlj
gzKj5OHqYrZdHiXc15kFlUCLBszguO/6aRdrOggM2EOU0myzHO+5HWbN8ExKcse0
kVcKWFrJJP0Asm0uE4kDN/GDwOlEGPM6mcWbsxaoWTDNiCt/UAArlSRSEPc1YE9k
8AffIJiRlXm3yoPOFQaqHdyjcdcHGeHpkvivKP1DnXfruflmYUyxGiuFG8BZt3oa
uqIKR1QrDd4XA9ZukBx8kgvIxT2KDvvzboQv4jiXeSEGJcDUU4y+QgKINU9LpTRE
h8ERgtzy2TGhLEGKxYo9haCaAX2WoPD+WPiIpZAFXA+bQvo0aCZbN5XlHBB28RST
Y7naQS5W0C5uxS3MROcTSEkRQebELvjQUTWszcf2sHI/1+QkVBqFkcP7F9KaEnK2
kiZqS5O8Nydo41U92BdLWIDtP4X8lR6yn6Pjp0IqSgEZ7UrCe120cJXwkQQLrHF3
9ivbnzM118Srv4Ee39twc/7HK5PATzUkz6/4tyJK4DLnSvHkTIkHJJcGCbZsxvJY
9BW6MQyA2J2F2zAMXV71Bfheymu94an+V6WHC/kbdbpxGrJAVPksjn1azkkkh6mz
uii8ulJp72HIaKwCwayQvpDZideuS6v4YLuY5bxmExfSbc+O/hyznq8kWXcgl510
cQFQatc2tX3pKDH0zPT827n6b6BetwNzoPC6E5HjpIeKrxyEa/VTosPcu98aMU9n
l3znG1NTN6VKuzrSsAbngw2ooeN7UBOY5/TqWOgePV/EVuMHSyo5v1NAUmaU48Q0
YMnNMCet1X0ZB38PtibkwHpbgWyvlZrlxt4FBg/oW/j6hXGiqJrd3dk1i8R8HghR
ByNEpiQ8QkbXog+1Q5LIqyexDVH0vWDMWV52eCVcH8lugPulEOqXR8B6DxApfVZq
q48TFhjpn89V0K1Mm+FL75Di4H/3fzOlfm1uWiImQFYgTbslfZofsMVfw46VTnvZ
ofMWi/z0VNdMhjmYCSD9JfIM7qUDa2Ux64M7t+WZ/ZnWn0dlxfD/D/wJdwc60M5q
kTYToIgIJJlyXaZWZGRBBACXgG095csJSZpUy41rlYgvLkvGQpO2lbhfai7qqXov
wT/9aeeukB0MnW4ZJT5bw8AHTT+ukaOhBjPRzLmk9oj79Pszj5i7g23Vt0krOfNf
/guIptrUdItNQIn39ZWHmujvXp583qD1+DZNCy0dgyFUu0eLhUYTO6Q3DZG6tf2p
N9Nb3pXe3SOKGCMQB1A43pW2HJPtgeY+D+dUM5D5OzQN8Hj/OLzPK+WLuh9OLsCh
y1QJ/1M0WudEBFgHaRyAp4XFue8wlV30OYtAr4NwLpetRlqrC/BplUVfZbyspZYS
xILPIxU5PRiO5Zqs+Gndu2eQjcYl+Shgl960u8Mg9H4RDF+n3zkaodbPSUmeWa5S
TamaMn5pvjSngEByxP6tuIDXUTHpkmWIyVV4RzAEU0miVup/Us42gWK5JAGXc9zB
Piuo72xqqrhZHTCUWZI+utSvo0iivvNYSDHaD2+D1mvPX9bg6q8SrG/OKOkkpEgh
K+hD42c+yd7Y6rB0wjc3vicP7vW8KExkoquZQA/96J8=
`protect END_PROTECTED
