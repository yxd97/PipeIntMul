`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qgRj68M8tRxiYzUoRfaTiSBpvODJAXZFDsckiEgsf1yG4y6tcxcUDHwWoTq5hHoF
PmFfl36aCTLHH6JnhVaZWmd8YvIXadK9b6YOZYRe4PHJj/xJMHfBJscTSeLFYu9l
lOp4pu0NoR1WgGzaMyHdy3a4jej0yH/Z7d2Js4igcZjNQTXgdkL+KFZbfhOa8X8g
xnIawRlZuWSmfj9H+5N/P8GtAuvrVbVp2IBL4laGqc7/FUfsymOOwXVZg/8pDaQm
8mHQeUNAtgNvtvXy2jIAYPhU0/kBXP79FAJY9+SLrwCqNfpEjmNFDT9A3M4DnAwF
P8ZpjwTo4duQU57B0QDZ3UD2Jkprn2UTPW6cneXX8l/P++mDO45mHm/MCJnJOQqB
tkPCEAxQPIH7y3+4pjGnjrcVnS+iKI7lVdNnZosw6+qji6Lmr4qWDwl5LqVeW5Ll
wPz9FqMwXaSL/4qxFBHabCkaeCHd0JQMN0GXxZ02/n7r+jz3eLLEDnoBW8oHfmhG
DorB+iJkO37OCcK/i+/0gGa1XRs6KS6lU9IyRkXy4PxONoratPEPEvuXrR+WBfKI
BTP9HO0+PGtGMyk28OGoPrbWnZlc1aI/HVlHV25C3BazSsiap7MSaLrI3Y3a6FZ9
O8yPggEBWW1E6DwrBvkcCG2EiN/vZt/cSltNr/dk9KyljaHfpzCp510DVNo/gdDg
Dr614BO1fayAYiVtxaLB0w==
`protect END_PROTECTED
