`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fKqyvLFG4zkvWOz+3hb6nakUBDkwneHnjsFtGrpTTjzLew+Mj6/dsDoJlyF+/x6z
bhAOzdJKm12Hr9cMp4OnQfICFGmviUUt7aVze3jc+W6yiSJWlI20eAEDHRKqJ+GW
tdeuWNyZTcl8dsqEHlsQjhF/zCNIIIt0Mrop/DmHRK4BrFz6RAY5do0BoIToYEdh
NRkcOt0y6QzyVK9fizMHGyyi0rO4WQRQhh6/FbPuL9X6Lic31JVDwAwWW/me6tmQ
lkacKlJwRninZW4GHRXwgqzRdWkKXlqg8nlg5dmliJwyKLcC5XZX84HRsbcierYO
tYocXZBTrBIi3lEoUJaswisT17Cw8MZA9f3nHyFQXhyM3UOZoFL4QBiD7CdMMUqr
XGhpXbuXKEZ/mxVum7ecPW6oe2MDY5YWbJdi0yf/KITryx+qQpIaCBtP4Q2O5lYH
F11x8iABZh+Je1sNW6SvjeRN5+DSKx08J0YIPxvbDys=
`protect END_PROTECTED
