`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FlS0tHk3w5IlgveDJK+99FrtMLVvR+cTWzsugt3vOMQJtCC9Z0RDP5msxwHWrcDA
nA7rsItXhAtlByX5hRrcbajmw6b8pJv0KQpczU6EAWSg7RTdonR8CFtgWZUMJRDB
AUZ75fDXRJ3WyniA4xlfvBiKCU/Ju/0Nw9+raiBpdikoCAbwqPCg78Ak6jYq2vbd
kXFPrL1OQ/BDRaYs9Vl5R4jJ/kgHTmdmOm7MH2lg+RsnPo7N2hFk7x0Cd2J7CA+O
CVOOorLPlcf1E4/qMIWV5e1XXtnX09JNs0uyyTM+Rzu7bSdqlg5VSK5R93RoFPDF
DYV0umAXmeeD/RE4kpOchJOfmdvqaQZOjM36vL47vYaxIltfJh/rLUXUxMDyNkHy
Cr8NPgHK6hKsW4Jqj0SX2yJuBWC6AUAE7SqwXHmLMnDZb+AdiYaalbmYSnjYHF7I
4xapG+DCH0H8F7lJYc4+qfuFOsetDouQD9KHx6e8fBkcTARUtNuzzvbcgW3MxGZ7
MI3/lqqfg3Pg8EIGxiEABFNHw4cvCeUglgbmUCVS4Q5fHQWx237TqMTBBO4mdGOa
r9zw40in45Dzb/ndsNZ1cdM9YQS80cMA2cUTD21RKrpAQsgdDfNZM2iyJnjicod5
V2ZPnv0l3G0KMZWo2RBcMEWJr4M0fSOvGM4np/X93RX5pIW2TNDJGiN3IO8CnH1e
q5jjlKqy92rp3387AdQoiqqkuXk2IFZbHSQ6/1BlzycEqnzQxYsgFWpoqvoJp399
svnhToAndfhY5qPV2B4TufD2OacFJ3Eb4FqzO1PvJ93/mHWiFSDvBeFr7Pnpe4fs
YUL3xo2f9MXzLfcyzNA/8f0FwYXN3+5fYuS51lcivf5KkD1kVvXSZc+7r497CMmU
LlkU2eEM7AwLTOhF/nZhhr+drmzeR8ON6VK0ME6uRd7Diti48lO+WbghbPw7aepy
bHhIQGYFhLEabK3CDfH79ZkGhuDHcxuKE0qo0Ja9orw4XxslxUBSbPmaMSHB6N+x
LbwcScvlefvFB3jp6jzoIuA+2xhktRgVCE0EKcwZaqb43wIoIfxMv05lC5HtaKtC
++FXXtuliGm0V2HNRmlAog==
`protect END_PROTECTED
