`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fslaxrn0NTQbvJ1uzr1ZBX8bbw+NyEQ2WAK2b/rF2XOt9YdkvkymIU/b/KjLHUiL
o8BB/g/vdGfgWEBntGxTdNA+4myjqhKKVCo+5+t1YdVwWic4GqrbW6pV2zLIrR+E
SgqXe6XEIbJTBnckOlPDKu/muGS75asiiUxr2FkxWosO9Y5OK9AnLKtt0iTw/E+a
IeiFyhZn4uqI+WtVw5Eow5i2aA+K4ouVPFRcyOCtUoyd5xxtIyfeqJT/EWFQqDUq
4yqiZRf+N8FIHchOMvJiJv7B+3nT0R9VqT1JOHjR8HeRXEKvaIlTFDgcZBU+a/Ga
xqZTjXchUuT0tf7aX1nIQLm0TIO05QlILmS2N7d0Z81mejbtmYbMcbAYYdi7hu2l
nzma2wXBhS9IV15zY5pzWEiYryWe0WJFu8O5k0D6yrg=
`protect END_PROTECTED
