`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tiPnY4qQQA3yOCy986pa7j+3Eb1bK0oYb0b679B8LmCD+MDNcasJw+c+Fj1YTWEX
wCev350rBT6d5yvHyC6lAOo/Hcd/R1jwKtCgQ3f1drwq2ywJZa0jKEriTMKTlwSe
PR5NSKyr3XySwwSDMUghxZcX4Bgmr3xSfuBWqjwJq4dB3PoJY5scwuuhQtbSFix+
p7vc3ZAUUIRT2KieMrWH0pId22QdX+G3RPd/7gtbRKTsgWmTChniD0YuySvUsD+J
6RAjUxgf+NZCV27RxjGo1VuAfgJPzFkcF/0hYlNjl3yv9hRn2A7d09O2H06vZf5h
geOR6AGhX98khQTMK9+4GZ0GuU6tdmZ7bkfahNnnd89E9LRxAY9l9wjz82cCwPsu
SZN8O4tHJcJEzOrOxlCyFw1lKgKuMe8pdZf5AbrEY7JkGmHWjN2mD2JicruuWGzw
uRtAH35supGoyIOXDowFXjQH2PR7gnB82klB+3MiKYvRS+M8ItU+L+HoQnhXO123
lG5FHVDCBPVSsjybnaJ06W1RMMGE+YDZqHs8ZIiReHDDJFYOmV8YsSI1gfSc3GqP
QVvCILVC+elr6D0A0+a6i3SF8020j9TBRFKCjqS6FdeaMFwOKqU2v67LuURlet4f
5sySza0s7WiiLO4RRzGf8J4XHuhy4ax2wbDihzoC0n8Hnmo+Ypp+JE7StEsKOgN+
leGDpjLuStvZOCVJigIaDU8vHRPoxs03qaXfOqUnhoPr/ij/03XtsXgcYRzBlMjv
dwMU3oUjnIFVG+NcSLUYgFQv5AJH4DQ91UY8vOkHzMbxxdPis4exRgP2gZe4/j4N
HY9RQQdALlH14KeogUp3lDKN+Nh8dhW8RDohlYO0grjjV9VjHILtqltUHSOvJCQv
JkzZcGVWIs5WSadtaX3qduB7bg2gd2SB51vbo5k5mLbHdaaoQbrf4mEr6pnXjmu/
lCZ/ywboEysfOU0op3AankPti9ysUiNH41VY3GqsZ5PWlQGYuUEyBHevlzesFsnI
0QbLD6EjnatqIhcRjdLKe/TQ34lirkNUXygWLr4pTeYxPJ4Ms3mtXsmR01X6gL5F
FOpTx/R5R9OuXglyYCYDDGUGneMALsOoeoJtOIJPFSLrU83TquzyWtBUwv1Q+BhL
KlA4WxxknenhxALu7a/UtkiYs+OqODIrgvIUVJxSdrMppjHkTOzkQTpRbP8d7CeA
F2UQeN9GEI4MNG/abNoQYttFClM/armokFEM9vRTVvEGn1ds0SdbeLD6cNKwYiVB
jNfMmTWaAL2StLcWxWVcWS8PYSIZfM7rR/wnBLuUEu+qp7Ld7Svc9nazFnuTTnZh
ZyE6GFbtDudH/UFadza4G+hvyuy55yk17XJPp+OSd7A7j01JfSBRqGG5s27ccPG9
`protect END_PROTECTED
