`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dg8O/P2/POYCtvu12rzAylSatvWctywwAKu/XutFRT2LHPrx5bqKXV8Jhg2tK2Ba
gkBfm4h0IKwWLNykNq1hwdcn7JU3oazCHMkTVJ0K/63W4VvUkFyttOudvhsy1QRd
CdEczfj6gO2+x+ibtBEWF92RdtrJgR82V7aSLs9KVhH3OLQYsHQuiuJaibRQDD5V
o4iVz56TyfZMA4XcVsmDLWrSZS6bGbKJmGKkxcmItNqKl3Re35um9PwZnnpBFWCR
jIRTaNBC7+e6a3fWfFwzxQHtxCvw/nR/13Pp+TJG3P0Asntk8c/FktP/zDTa1F2j
VCcWzcCvKVnDUiRwmoMB9dCbkK19ocXes/O4ahiYqGj7SHZ8zt9suC/3DO1cluQT
TRAyNHMUYmAComg63mOpT8ttxYv/M7mrA7xoL6fnK1G2vu21cup4JXe4QUQfVpuK
nAVMtAMohJT/mvR58BzW3xv/cp0EP2X63nO+OF6PA2bahNVw/fU7i1SuGN67oN8/
jIZGGcRAvXGjNekuJQBeyjCrfKChinWYEzXUCf7/3N9ZOFa83QoC1FbC9UQ47H7L
OygALYcBpNspns6irCmP9eK8t9QF+hMZEykCFnoUPt/tlwEkHAcW+al0Bi+vu4+E
NWDP1eOick66umjnHCjM7VWk4q6NPIFK2CVtRDscLMJtmqUc8mES9g3VjOlsLkTn
eOM5490eVYWSJDef9bnXy72PDUTcqKvK37dfkK0dU57QuVnnGpFY3hq2rQzJAX7l
FmnLvYhE7zvElRr4P/hzB0sjHS8UAnS/joQTgfVWlsfaaBwAYcKYqcg2vTEc2daj
TVZpEji69WhZ9RFODxsc4iHebrCwXZFLjic1bkgXw97kgoFjmO+rG6squZOUyluZ
nvs7Lli8NqnsCHlp6niTdhGFtucGyqhTY2jR/CIpKigW/HoMlXJMqeYM0CE2JTJt
7QUP4hNzQ/SGfJrGzchLasnzZrAqn2st5eDv3CZhIrpRo6Lg2VEWSEEyxJDNzOYi
iVBSIFWU359NKe9LJrjYkZmuxd/3TPGEBoRbbESC5JxHuqEiVZJ1CGIHO726sI4b
S2cFV3VrVaMrLyuoA3sZUFvHYFufEj+jjxrlV5YzWsr/7FNGDVnmy0He8YWhTv59
a1PRN2eEI+N7/OVZvhWJivy1BnBPlgo6kXt17/POcIIigUreASHdBbT+cHsje8/q
JPlkAq6fGEljMm9RZkRGDrctizNaM6udplVOyZgwUenDjX7HVxt6yjNAY2lHJ9Hb
30mwlczrrB4sP7tLlR6SWiQOrpZJJ3NnqPZiGCAFYiC4kYxiaQYHNXBkKXJk0qNa
HMrHr1hjmimrhTP+vfOlcj0jeXdu0kxwhy+bETuZRwAkBmLETtINcSwmGukJZt4e
P+tpdEb2z/lslUKnuIbCC56gECsW6N5wfngcc4VNJ7d7+0sibJO1oA2V9BS8bCtd
lyS0a45y9R53JOZYreuL1ggg8SMJVG0OGgpUsExyBNs=
`protect END_PROTECTED
