`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2xBz0Z4xP68cJeb3Clt4RiUTDmJZkwquE0Ubkj+RigALUDvUeYdJHb9a2ouHZTLR
hFThmDXWZDjqUcI6OrDt8DUFnbwd+1JfCq7OGVcwMbKRfDenSR6Q0/bMI9lWtH+N
WRApUNSQXi32m5HUVMbIn4SPPlDOM64WQkvOY+Oa+YLTEQfLqoehsgjRUrdf9zDD
50X7RViyfQgGsWcXLWB5LAa0cvYlxd4UdZAlY8aoDLFaSFYnURibXxSwpH5VpJfK
`protect END_PROTECTED
