`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c80Oc7WsShf4AjIaxnqgzUQqcKqkXuvRLqiNLDF21d7Ahn7tND6Mm61pju0pum8o
A2VIssjdbDFGqmjlMwAkp4YeqqiuvQzZC2n+mKNkGyAc9Rv8b60NHLltdVUN8oa3
ybKjum6sX4V5N+0HhPL7cQAm1Qfrwbnmy0RSqLSZHzgG3IrLEXbLJD9pVp7SH3fh
lU0Sx7cSDBvWvfRNB5If5yKfiB+sPVruYFRBpRMUHKC2jrBZZuwN3Mv7weGlRNfK
g1LQnbEHq6wAYZuXmFFXHwbp6cuGtV2xRFrexweh3K0gIZeaZu74UkoRa/fMHJEg
YEHcH7Y5P9E6x2OijAekKA==
`protect END_PROTECTED
