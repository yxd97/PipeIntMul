`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y0gqjdBPiDgD51jdnAT8y5XaqFWxSSns9Csiys3NedO+5jYbLhrIaNsaq+b7IQGA
pTXq1KXcZydOMIQxsFMztzSiaJTXHVVTsait9vFvTDnsgLBf1Btr8TsEesbNLbE5
flI4BQ5drpVTHgp7IlEv7kbeTy5R500wtuM0VKMsd556FunD5wxFEAYpCbtBcnqc
G/Uys8SfrFHl+8u5xbQCjok56y3slkbx/9aUtVmREmWluDkKYGFe01t/x3TV+JTr
ES7LsINU62N3Lez8llsJyCuoaVwE+smgnZHGwSJR60NE9xKgCMsDQ+njOjRiJMC8
ASg9eAmUjtO1B1Q/ZUO6zjgBYlwYmIRBw4xHBgDyvqhTfVqqC9oHk9craAKaEert
SDSBFi/V6v6GK119NJvaeRzFOWy4igCCJynhrQegRrTIIhETTzQtyYqHL4JFoi67
vwjFmzyBQ5djv0pGlWhrSPBnOrYhuXO2RL1DgN1J3WV4XL+u4jO+k+DzsHwTJiKD
rG3tYanIIcK+vEyeXJIgWTSB+wE04x9rechgIvCdeh3iMgw2A/OqSHaZJp60/Kpr
J/Q5bEvzpygDtnf0UGRr8Es7pY89yuSusQGBz5er8jlpfqTi6lilwGp1/MOq4VgT
zXUJkAL0GbVXzVRUiWDJ9aeJhsfM4hkCL6Ihhu1aJeXQRVgdQIjH/Xe62yPnm0dB
OWwZuueJbyBF+D0bucD0BQF+zd5S1gEj47j0ixJUmk/yB2JtFTDEK1YODOOlOHVN
+qxMC287dRvGUEe3m5vQQPhiLgehoN20oV9fHbP3rEkRsoGnDE7oDTPv4i/Lq4Z+
/QzyckGN4XhVs1/uDUeHJoCWsm5njosZzrbkX/DpeFatfuO7+JZXblpKk7inUSUV
g9SA5ua6gfYF1WmYXg9QTNmWerVj9BHztoMFn96xtJXQ0ctsYPs2OfMav3AXv6nb
XRDxtVksAYg+6TBZYaS3DGWQa5FOmKTpUivdwkmpbUNxdsG1hsYseA9hE0Y7Au/8
2geX/3s59bU55Uk+de4bk1q/acnB5cAurkgVMsxf2HPaRRBk61J2+B3SlQX/1Txt
yw/J/td0D5AWnNS/Llc8wW8Ubi7PAqJtD733cvczOscJ13jdfTN3skjJhRzLnLvM
3bVO4M3srPsooa2P1itXK7DPESJVV/U77IBRFarykgjyIEOJR1pcrKpvtq5QUnYm
Mcypu8e+e+bny2KHw92BiRydwsHTon/DWNQ5gWzYAur+ePNRjt1NCyPIyVp938Qx
xDvE0DXOGsrf2WR5PKMihmUyuQAtbnCFucaUHDNyPqmkZt5msUgaofA9NZm5zucq
cTjWcv0jj+QDygKsyawukyfti/lxuCaX/P0gT9wmLYugc+IzHfjVQQBxtzTK0e4T
0uR0lB42N0uCmk+DTHXCKg3YwCdgA5sTOCkHYn4qtTGYbjV/CVHNK5xvgBJ1Dmnz
DDNHsUkoCGDA5IV/OjjpBUgwcXv2CG+XDDdwaBPdgQeucKgDRe3gEOibnuyniTMk
VHmVG7RYy+kZYn59UP7lXbBhEDLcy1P6oCveWH8G6bKWhUH7LLOY6/InmZMcFHZC
lVxPAxlmf6OFKSPDSDA7DFuQWfqzjxFsqaHaxcL2AOJBve2PnBOYbIhkYVvTFEPL
sXB9jc866+VYEKLKConqajSYsZKG+M69o50B4g9YeJDL7sC+Xp6N/Yi/WjCSPPXb
dXrHXXdP8tqnn6SoVaNUY4TqSu+BnpjDjku36bsAqd0w5yZ5eh8jxzy/kFRbBMKY
38JjrYL6R3eKO3rlfyxgzfW6b4I5qZNtXK1nmYZDZrHIV0/RwBe018p/gsdbJhwp
MPNiLQmnTQKQQ0LabiRHWGwoZzlhoGlx8DezdX1RhcXtFLGdnv1WEHumdy2P+UZY
JZ5EhjUZFAkI2DC8Dja6HXguzRH4JQNnCOMywQPfXSJ0+OBWQUmAE91CJD/DF4KO
ximQ1IGk1zomtnoOT47vu49GAGOZ/TOGrSiyLpGKgLmL83H1CUGOJ2ZOuuxNDpFT
4IGUkd4nk51eWxlusD6IXtgXH7lTOA08XGgGOzMEFfZ445wVPhNbFcsMoeAbcDj8
YRKySHbSJtpCUHLU0w7mhhb6jSyW1KCIg4Inn5rlIa+i86Al3JxQxuZI1pVgwSYy
MrvgLKyXyz9orqD+KQL9MHG9pdF0rByUHJIrAIZVvz8T8af9dGjdGSU+lRpvg54U
m7BYz1WDIgbNPyPDjLZz0qhapOrU29vV1TOprHC83R6zeCNi07fkPhN+WbJoZwLT
vg7r9ocf0mjR4zmMQvSPNgxEyf2484uispup2IOi1utXLVfLxNh06EE9/mMibxLf
t6BcyLb9To7GeOkELi76YUHzxiqsvqTYYYAu9tOUgqm7MrEglIuhGy7fBC4xZq/V
izsmh/Ds3P1SHIwD5E6mskSsLngctFBAYCdBGiMBGcoOlxL8ymA/Lo6oDTuBCsIa
I3jlcLk+G6MD7dg+JwuJ1G0b2jWv2+3lE80UnlmFHFf8IdobXWGqZy7RCv3nv2zf
ivHtQntBYdx2Vtgbd5xuCLeLW6blGicMLVSFIeuUwFG8gWKXxawaIKyF7Js3KXOl
K4mDTtLq8YpamqhAzSgSFNySOUOGhstNcCn/MtYFrnjovdjOK8Mg7Cg+ZcaDonKk
hr9uT2kgVSds3QDHZcJ/4crOBzj5MUahvWpxOCzdSpBWTizaJKv6MrChiIZt1462
FhpThfBl6U7QBsN1YwKt+F3lFVxaDvcB2qZocwlIQWsaEQ4Lx+CwWKOVnm0UWl+6
Vc3sATSgsvE10D2XwcVzDvQAu44MZ+eneo30GAbj/2dzCFdxVuryUOmvjVVcewkI
xZ4WzQWLCWD8W43+fcqTaY7szo0nMKW6B7F8R7hFynrwWuV4jcteNY+8tn+vmUUg
KkqUQiuePKgHpUn1dGb47C4QOtCjt/wsa4JjKs3DD3wvdEHmTzVf4bX2HanSy/J0
aEA+AXSKrc9MGMSDRiNQ38gcTVvlmKGZOz2wVxJWTydCr6u/PmtGaxsFfZRRaywq
rPVjJkKEk35su/516ds/Xo2vpm95Jfx4DHUsCwgVWqFBcWw+SPjrsxgqgX5Np8vz
4lIh+ubVEBn+/S08zhOndPMNoRaaKRmMmlIHuBdb5wHYqT6UuaDQHyI7Vq5b7OD1
9uAjF66KpymO5w+EjpzBc46/iO3mwHkwwuDqWPIgIfCPasdS1GIQ9dZaQSI6NpvO
tN8xDUPnWJ5ZXphHZSRuPJUQFR80EF4LXPnNiS+6YDjRTCHLpLX3qdTzWuYQi4mA
Fxw9mssSqyz4Q5UcPy3+PwYfd4iniCbioheAngK3mzzwtNFZjKYFSJidArUDP7BV
maEogll2ry6gkof7I/aukbM/4rGuW4kHG1ijNa3GIOPdC1biDwzCbzt5rH4sAl4z
aUu3FgemoGAYQlrZplZk3ftQgP2IzmqXAnvXSEnbdCSF4XmHnsl5F55v6JgXj74f
uGsg9/CqtpWpf61E9DoaHcQ5qsvrZBHO6MiUSuAQnLUtgaxaV4ezta3GjP7LQbHm
JC+F1Thmqo4oSDTdeaJKo7IevW9Zx4R8MsrKY9QK+sN22ESrUVU9F/F341wgcaxz
zxfNOeMopU5KT73/iJa/k5e6GsTdkPqGUabwP0dpNR84ajJRDcGj5KW7OKLD9LOJ
jf1iJkbBMXH1nD9T3+2C/TBpWi/5sGmdDYMBqu4DD6wEWbPI2oK4i6VeSzA9wJn/
lrwSvhn1vz2xo1gPvoBuGrAfLOjWwN29SdcETQTc7J2lNSyYwgrN7zbLjNeSUF//
TQMlUJ7pv/7ytYTidLpIp17gQ+Wzeq8ntSdPfA2IQ6Up/+x4lYg7mJul3QzTDWzJ
nU/J/EsJ8CMy068JlKmxo/ZG6L6pgYudtuElJ/oA9Uo=
`protect END_PROTECTED
