`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fAsv2RSSQjWmTGFQcKLT6AuhkptLpAkUpTonuEZfYiCbTSutB1QeuEec4glou1ja
3JW7utrCXI3lCg8f70ia4ytiEKvBKE2CM8gEmzD7Os9/ARlfPV2mOa9y5SF/UP9/
YTlmadmuHKjmx5OLmLDziXUdHBdBxKzoMp01NpEcDxjfB8b5Sql4Qk/O80J5dinz
IeEc4RMZE4x67rG7Lu1g+v9aWmgA/shwU56U7yIi6YeeLidMM3MwQevVTnWFxgPS
NCQVALySb3E17bzDwXli+tpxhXVTulhTad3+YkIEvpwM/KjRaTs7tYCJbG4qwr+2
sco93mu7UYkne/bSrP6mRw==
`protect END_PROTECTED
