`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVSFsi2d+bMLPoQQTN1tI29/4s5Zvxv+HgjMJ0YVT1mvP1Ef3+olbJPQGmASFxbk
3moQfvAxGeLGkNmJQZLF7RTVjTqTIdPVjmlhCbirmPJFcY1Iu6iDvd6X6gRVs6Lv
TN3WJbyWpUflc5DcZQqmB4tmfAJDVPwRcceGYQgpnWz7cgjGD9rvef+HVeCkGNv3
AZYIUdUbe3HaK6lT9rh4QHxsAJdnK8f8ZG5XFzCQETHwHykrlzs/Y3XgcuOEkfCP
1bO23AvGvQ/6g5cxoIzaWiEh2VIrsg0DQHEVsKljMVEjNakMvpZLso5GT6Nk3VyW
EyvAqRg8+J09a7GOLno0aCTtdYtOOA/oqMv5tdXNWZm7YtdilZobI0+uOypTkVxx
hqVc7pXNmK1PCoeF/033YlAHZHQDBYJYG5ixS+3D9wuM+mkEgjQo+iV5j7mGDldw
mAoMtR5CPsIeaQ7wYDxPvGV1G5j9tESazpzHNxdiQPXqnhF8aoG2F2bjxEszRQ4f
lTV8m/9zYCjDxgZqoEHwC+rNjsgaDZyzwRvbfqKH/7flc+bq6+7bEVkoKW70pxLe
43TmQEWM89zgUrBOLtSrRiWDVMnY8FpwgzIvLvPY7T+WMNyriq6jk/oRpGDS4ba5
60MsJTt8CeB5bWr06rPIjA==
`protect END_PROTECTED
