`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDzvFZ1BX4b0k9d229Rd8VyqiIYpxR3M5tn0AP3MR4BvXKjxW7AALw8eQCpICyzu
u9CzZhpJghzJ/FROzhBngSxVY8AAvSXFJso8kp4oba8x8PmAE/2EJ4r90T0aBCVI
C22LVJwvaN8F51FGImRtPm7SokjT1IoHsT//kco447H7/kCx4UGprOTG5fiIetjP
gmeOJPzTA1O9Xwck0mSda0pUBFysZd3ZMkWw7oxTuEinzn+hle02BAX7CumRuKiC
/9djK45yasFjRhoiLIpwnDCeJKIpV1bvpyvBb1wfOJgp563ew2H2/Sr1Tu4yHIi1
TTXzdpcHMNpWKgsvT/U5fMEbbhy1ol8X/vMyqW2gaMo5f9br4+km7b2vyd0dl8Cq
/fCbV+7VhMXEmXgqZEdCUpdZ31tiFMkWn6+PsW3MjAtFHWtCr0gI3nbunFrKwY1f
oJwnJ03YO1YpNp/wzXXhxXyRlZnYh66J6AYeWcllwC51sZ8jqFG3Fc1q/cw6uxds
DrQ6eO+MJMjrq5cc5koNZIL6HyHvmCrskaO8WZSvLCwLrk2LVJYcHI7Jy7ZjVzu8
b41gzCwhHiQeOEcsa7OFw9IiNhFWyPk6ljadboAX0v4HWENHyGZp99FNDeQoUT7h
CJYz4HHM7yn4SGk+7ALgdB3tjd3uqXU/Pu5XvoYP23kbNcaaCxGICR18Oip9XiBr
BuLcgf19KMrICIPyZQxAwFfzxusXQ7ty0uglR5Eol82nxmWA6Vkh+13NezDrZNjT
NTvA14o6ZxdUagdYut1HYkmmaGHWKsY/muLLxm8zVYOovArUMpIGMTPGq2gbkMz4
frIBv+TsPF5dSMnHyvxoSbYAYxskA5S1W9HcebQrfbhMWIW1aMnMptg1lDARo1Z4
6gjJLraSqqr7O8WLMZ85x99IH3FT6WtVQbzKFBvT4dJMtb/9KSnYpCOpvbtjsLNf
Wy3r/0ARcFHaKhbfEIqOvkPd8grrWfg4mbP7aCrfsu+IV7P/H2rSX8yUEGRp3Y9g
S1579u8lDQkwx4ppcxh9AUQT10k+dQYWM/WvDpUeBroT9DBqFlw1cV2sEvuqZJhY
P9/kxiqfw3BW2EvNv0Fc3snfCv9aQn4piupwT81Ivxf3Ejdv8RW34+x/55domYzP
K7fYbIHZRbxbR+iIcfAIi4XuAv4QulZy3KvLkfVqA8tGdVFfzUt4zie64saymyxO
/eqJbe7zW5sMB4/4JT+D1aV8OHQyn97paqjXv7r4I2K7J8fhJ+FyVtpxMUuiwO6u
UwtHu4YDkJ+P/D41BBBv6QIlW2YB4Zegh46qNsGDXO3NTh7x3ox8TyABjwVue6vn
z4uf0mmY/VC5f57FXOZDVKNn3wvRqzc9vvIOYCvLVLEJpc/FpAtMWwCDUmsIXg/d
++3gD6drUwIYJIdP6CITbz21IoiiJ2cQwcbFTd8uTVZN8Uz2Lkqwf+/521Hj8ZH3
zFW86ZBf58Lyjkg6P/8msu3GSC/0suBKrnAGEB8+bZdEvZjMo5iWxNdHnndJ5xtz
84X3vuJxCZxttKjaFRtV6mTjNydmZjr3HoCxeO73xPlEHUfV+LdWSp4HLAF+9Vco
dSOM4ZG9unW2PrsY1XAF8YXzl0D+Ki4G3NDbbrzvMk2unMq66Sdg9iSggy94FBWa
QwesxNyabmqw+egkJO8+80C7t6tnDu6MgzF7wiMkOlvY3HLJZ1atyvHE7DlSFzDy
g2/gCWQi17+BXxr+zbGj6MAe/JaaEDdle6+4aFNKpbzP7CIBkVf4SYgIb2brkStg
BoRNvj8nYLooLgQVi6gaxpRkZXiX8b3cs2iZt6/SVEAFW+Qm4zX3fY+ygS6cWhHf
4VJfxE1ahU0CLVKC7Kw8PWXpLruqDJyXy+b801lPu337LY2L5BwgevujoWXRt5Y4
8PXZ8ui6rJCvoV3tJxkRlcGNJLun0WJMVq7uLX36OHd6cS7bm5XO/QC4yGIjbh2L
+RMj92S3C56yoRn8gQ8YedZwm8Fkezm4wo1QtdYAAalpKnsgS6uFKUJGQQiiGqBz
WYEjGmobPCn0hs1wlETxDWnUg2l5UuyrTWM6ilSmAz3dIus9sorwH1WReeDWHHJ9
kyoF2wfiuR6zBOTUQt7i5fInm/4hYL0KCc+V3QldOiBK3jaSOTZv4TqXdwtkJCZa
tfNEfoXzJVm7uTemr/41Qz+qYUDbHvHbOECqw+uOIFB6unwSP0EoMBlHJ/+pZte0
JAFGFiTvp3Qy8Ze72KxCIVLRmomSL4qrjyCwR0I4QWI136xOiLkebzjT5zgieeHw
qy31v1C+rQYql9Hc9BsjmAiPT0/PnCUrmUhdwWhZv7ZaotuMPjO6NRqozCb/YWSA
HvO9X/LxGggIx4Ztus5HNUvOFaN1UIIzrv3eC6RrMMW0ldIi4BgWR24uxCLaPUCw
CNsxrdkrm0PoK6JlrX2k7pc67RFj9QDqVUcOnUDJIstzwdUgiTbU8EFTaZmbiXiW
MQC+rcUSrptQacM7uzD83sZHGFrsO6neEcoKwKyKvxwH98l9Ibs7jYliAVUQc+uv
vciL+1qHcRMPUVF5Zj/rSGusniohPu2H5tA1mM/J9OsiwrlTzVqursykBRc/EKMs
lZTZ8ziFFFA0iTqkesO5Sd69PjYPyXDzIF6Q4w5ZN4+Z9UwqZUnFM0H5plXvEJsQ
/5KZFb2onkcbxBp2gcX7IYOmyY7i4uF6UnH5Vlk+IxEQOwCKDdweTAmgKzwBb7d7
ITOk3jQBxCeDt806tvdoZsTBv95/xfGK9j/wVTCgNvWhMoyqkUkRNvKnc2Jbts1x
hbLqu+Tha65c4c1lzUPUPL+MJkasTa6QRz4bHNKBKWz6+i6YInxwf05CxfotUwdU
hAg9VM0Z4p3DMP9sd8kmIp/qZFfxaHKelyx35YNMLHvccLWer12a8BbKVwxim+iG
ByWnMnOVViHwsQvxuuoQSbg9uomMGAsM0RL8eRH0SWw3j/0/xz69X1mzUKMjEhgE
zHv1JGVhe65FOz8LTMaavD+XuBFRujL2u35Wdq3S4AGvdR4prLG9U05BItkol8Da
YGebHDZvvK58317m/A2M1NS2fPlo79qKe90s79aSACg/4HZcGshjg3hleS13IWVN
07x48JRegAZcz9LPKUblvW6So80iNL3w+BaSheDP2xXI8prcufyzkGyD89sYmvHS
PbZobKUCw775bATHpKp8UyVRZdEg6Hhq5kfk3RFrMbksMviTFsL0cpIO+eSaDR0G
gKs7YyVTpdtDWE5wV1ihFYsA7bwlt1oVdt0n+NzB7EP5FL4yIDJEWbfHfL1Gh+w6
hjDU5V3CXmFj5gE/xLYxCmvbBVmFjYr1wWUJzyWq9JXJ4cM613CoFNCPO7Glutd/
lI7Wwn5qwZ7PzBYGeZZO68j79YpHUTfMR3J1lzMZ1V2MnPGqnEYHgFCdVhk8jpEF
VkXK0jX9n/IIWyhPo57PoIYT+CwDSC/JRpIQxUkvsiFxCvi8hJkAgh13WEoMpXOZ
l6wg8Z2Bc2euZwG8V8zkzltm7HYE29UD4dg3oEGkFUfVnQJIEsKMzQWk+9Ed187n
ZQ6UF99lCqAITQY7Dv48Pz/OFtoB6eIjS0kiRmIC3gUByesf4CMd7dV0YjH9Y0Qy
Hq4vShYN+YqZ4Sf/LBOxmhxJMkzIg6rcPHctkNDWvpNPiBCa9rEf4+tlX010Nn78
bOyZzySZO444Rapz4mlwPM8iMNQk4DJUqgLR/gYx0Pg5N5i/PRdXbHCm3dZSZXT/
N/iMM0In++8gAoUGHWsevsYlpZgzh+58SaxqtpZDaiwb2XA8+ihWDBTv6Eiyj2F6
kKfFBLmGbSe79bb9d0E3mIukALkH5Bk1XrxFX9zbmI+2kbWh3+xrX1JMxGNN5KGI
zwii3wq8a2opk7m023UQhIMEF61nb8USP0PF8S2qTopv+1PqDLPV2RAO1Jt1H4DV
2WLtAoXz6f16TjDbMMzx1vRwuyi5XklU3QrhAfjAwK/svxpXi+qsjkKLPZ9xQRX+
NhikgWMprSmqigPlokwpLjNYFwjX5zcY8WTs8n73cNX1hYbPirYrCZGs0gN+gYKL
jRsenK0jnEr2Oo7c5/7hFKygEtDJ08516+8B9AZYHU3IXx+TQg7mZCYng89sn4yv
TFtGMYcIEhq8FRqBe81t0K/6huJLC/2nsoTUxSz8z6hXQRwBUZEKxCFjcs3aNlVh
cwUKWQFWbo7QKuh9vzpEYKXe5TaNRmxtpnErFH5RVXxvuobet/TWra+/KGPN61Ep
2ASOQuwun+s40IcC9oW898kkPumSxf+yD3sDdysQrVPJ7J4xVxqKNdnWDRXwqRnm
a9yifKwIA0emhdnMR0LBPX6wcusUTIqLPcnOtxEuwLMbZ3qLavhGkR3JdzUaEQfk
aj4kKIoqoTV7gT1lrDwq3B58faLeeJrMaqv0SwrdgWfpf5q+C2MkVzGABrxrn5J/
k6pNCiQSTZ6rvC3bLkwx+DGNseA3OwHLXkfAYZiInzRBloY5G6EQ2Tqq7vwv1y2D
NWnw9gA4NpAYSpsO8mRKaKPoRoMCdyCjyGPTLF5wdJM+MeaCzVPv8jgdubcq5xWS
9qnNSiBQtZMewrUXwrS+YePVJDOk+4xrwNgdLfBqjGt6MqdYG/68+CSAfKSZCw16
yvW2mUi8c9ynDmBQ3mRsUOHP6R4v+ZJTZ4J5mhP1Y2UtnojEOt7nrK0y6i1/RUoY
kz2KsQMDs3yrZUQxFj928chlGjkKe9UNitfeU7j5RILN/2JU6Hn0CIh9x6bBItjM
hM1jv2W8EDOIbsCE6aRn7edT2/+MAnLJ7WcljMOH9/a/S4HQIDa182YXrNjmjPVE
bTalfgX41Gu4fK7XfwWr03yT7ijNN7qo4wGUha6K1YGKMEjvYexV2KF8WwNgxxn/
xD7vZxOhFZwKTz/LR9dZ92oFP/h0SqH1422JKnj2INM/QIn2uPOwJ0d2wGWDhwws
S2znIJlRbzVrjDf3XdII9s6+4Xt+Kb/vZQMRJbQn3lcthsDCYQkojtRXC5Ju6dvS
leyW0H0/HydWpHNGxFLvEVtpOT2i/NEVC5wDtJhgqTAWbPTw3pMGr+xz05OefuRC
0tYSEhaYKNamwpVxNZlTN+QyA8SwYNYpBGLhVeulydo3vj67IOU+JAH1JzpLUZ8+
E54bYuRAFV026LXuDxT2in28e01L/JN9lprlmUrYJ/zaAw4q4ZFskPP87Iw6KqOx
XG+e3Umd/tJ2UjckIlAcQwCccm8zwkDXoAngAbFNlkASFcEVf/VV1RAQDHEaG/Cn
Z2OCBUG86kit4+0vzeIF3ndSPN4s+Lq8ujg+DjKx0jSy8gsj11psNAli2j6spW2x
oslPxadE5QSqPBFGm27GntZJagKn3QyrQWYt8EkUZIvNfEPKZ8xfYsxu9UBtNI4o
2MqINQEb9YNob/f2DgkX5+MlPgy/LdqcYzTzeDR7qzRw8vGPSDB4x+rSmqB+l0pv
sF1wmOi8pq0No+VMd0NllDi43sQWPkp3LkQyCl4ucjPLdvycOjnUgvqILYksojm0
DHcjrtyOBXs4j4W0B8SbBf+If8x7+kTrlGIQ8c9dy/rwlDkcI3PKAW2X+x5o4kwb
bUQH9o5SONUh5CgUJLo9ClVSTwN5tcn8OazCm/l3T5LX9bupaXD2IvMF/AMqu9Lu
N1OLeRmi5Re+anarS4sIHX4E+dbJgDxYQyDyex9hcAUqLKYiEQAvXtyj4efZuhVF
dQHGbVvZhI7pOGEzNirF1plpvj9zqQHzyEnQ1x7sr7DdmOV7OE/FQj84gF5C8Tv8
Absr8mikqohbGqtwjpnlLhcd36xwyNR9o2nky9chnOY9oXHWMDt+wSB1ISySzNAA
bA2oGVRA9ZAXQ+Kr0IVQyp8y80hf2wi8Sl43ZKKo7YrDuuNq8+TJEuzZCgJO1TGf
EePDrfGfmPVHPtKhHfF7C/oHtO+aupJNzMtHz1ajbjE/HjqJ0lpICseNFsTYFV3O
hE5W+DMQ5Min664Vnz0gAOF7zS3zFB7c8a/52joI+0b0N8z/l9yg4pdcS+/GGg5d
1wpRYVp17vrJooSIKjOHJzto6NHOCU61R8CB8j5YkqtjUddRDJZhxrSFV0a01MWK
DLw9bwpe47HbJm//1eEiqYdqWjs+rJv8167NaNzRV01K1k8scL5VttOxAyQyvuuS
oKng5yNDNpIiUPSUdDyfiyAov3hENt72uUbagIhobJEj8OkbBs3n7RWyBdej90bU
8DAJAD9KymIkCvbu2vpfAciLQYtVMFrSpOvBoZDTdg/b9pN3vN5lBmC3Atsf2BID
s+rLTcZchDegDEUzm7swUoF6ffguKu1Fg+bQGRo2yGvlmWb8gZO3jpYv593H/khh
iHUTkJmB+Mb0J5+DujdU3deZBYnmlUIs2w3hm9z8OfykT3y9k3h39cPP2GIu9/qF
C5KTuhddfwT8p6mvDRn1CtqsWM0+qmwB1jyVDPQLaby7EaHJ3xjzGc0wexFVXB8C
ax54wqkL5nxbkoA1VD/i8b1Ud+8XOmV/Dulu3dVzkSDbQgT6iHdp293T1s15XKnr
ZsxSOHDcDjwFLr4eDrfufrYoX5e/ixJ9R62WanYR6XqttrhrRyNbmDJ4oTkyFmEv
z9eI4E9gHAxa8ZtUho91g2+nNV6TUAWF/ojLKtg8CtclZlruJlZupOcoM9zacbS5
n3I717iIP7kZBOv8ImxWy/gob6xy+X1ro6XkuyBSTW9lJ8Ta3+SqeTRZr/lxWquI
tNIAtG9asBAS/OMkpvaX5BTnYEXMwtm67g4nDYdK+3xCBMfRNj7XZjY9YOpDsi92
6PhF/MvIiGsNGt/LGlSR5KamIIlDuToNKnkdlEvUSgtH05WT35rxQ/Fj/mDS6axI
fwv9yI2y+94/wsy8nBpAGMNfifReBBzSo2vnO5kEKV48qo0ZisnJUy62D5ia0u9n
IhHQXTSeXxnnbAn3felSlrwU+9gwfnBeL2Ptiv52pGd3pvYtuTdJc/Su0OE0muIu
/zHMCk0euxjjjbIM6zk6Fr8gBq9y+vrzdR1jyb5lXWXrAmdUCEoP/FRXHOLBTuD2
1ag5Tmkf4/abjaCeV1dRsVXjtKgQxvn+1PXPJe7IXHEg6CVPlNvsApU+82s9PE2K
G+2uYs5pRgJRpH4dT+9Kc6XKuuy2iMUtmNOlAc3r9QhHtQWgTmSi2GWlvUBYdK1y
xzI16GWKjDacra9wasjv8KdJ+ROUwzzuwo3wf6pU7Oq3B+wuMQr2bHmZTRRKMphv
dpbLEar2HJmKXvYGmM4j5ThW+vOrXi+MVG4IyGS6oC5g4ztUjznn0lrGCpKWed3A
dkVLZVfjjO16V/+Rzut45BZIyHUVJTVDFKTa6SUSp+MOJJ/eCF/9/qTgs3S4qVLF
HKxqB7BH2AUiAXpE3NbGw//Afm+ZD2qF2KPkJ7Bd9hBTNMKvmmCxM3OvP1C36uhM
seYRqiL/StgCZrvF5PCGo+qqtDg55mmoCuZK9J8IBIAuYUaMxxuHwQf6iDM14gNe
ZkGfB24PzhGF8WY8sOgaK+1/5IdrxPkHjSEckn8ev4UYe9rRn/Cg/uSbY1EQspxa
EF9CeNfbBqNhxSpd8WxIWp5gIJ/J4kMDHstCvftolVE5D9xmp3GG9i1T2Fqv/jUR
4EukZilHK7END2BBNpXHOlBP78gt1a4ddDECzMIUU+08xdmjnrB1aihOWty+Ahwq
UvXXAza4HHtTG0/zZ5gs/Ck/sem/IHE2Qhq2PEzFr71onpX1r94K5ppkK/RsdXMO
qi0sH/3ILqnRO5olGUBmwgXSgoLtEMzFNvK2jPrjRE5DKnyLhvsgJC7NJaGWnysM
pxRmiYqS6bVapgPVzK8FQtNdk3ei7xZXnvT/bUULcChgSp1sdckocztDfF88lAvI
BUzAAlwPHPp3zKG18MO92jwzEBGRptIVaEgDU93CGM18JzNvIas+5Rtjfg4afz4O
Z9PEY1wY2gmKnQYmzu436B+sAlsdEC5/UCvj+Kz/v2S4tLudD0bb871Rb6TbeFfL
WdCp553d7tJkfWauGcnR+b4GANoRRwVD619WzVvBhExlN/Q+S0mtJmuBnAiQucVL
MG0E+GdCFjPyxjehNfy4nP0rBlSqHWY+7pDlS99Io2TqfxZkaNCI4F2KcnQTu/Lt
ybMpzSMbI9lBWuLTfgPgAqU0+kmUuvlz6UAdNEDLB3acHTxAea8uu1SujmPDVDj7
z57PA4i1VJ/URupk5Z01uXzs2CXXCh9PP9ffwg25r39shy8ifZLivEK5IqJ9Dpop
wZO0eIHIiUcYB2pfRcuIx5nLKGfiPVJOFr+T0dE1KPLW2oV3rNktbEZYdqKqYILh
xITasiFUcDXCiYW2yIYFBII60Y6S6a/MUD2UkawX+ftIQIwbmHmMTrBykHzK2/FZ
L5EKRJXR8dAP9k35EhJcBWIpijSVKNpFaFfVZhk3odWwJYCOBXXpxlzJIntzPaki
BUcOUqo6H0MIDAawtmxOhmJpl6WuXO/pQgr0kOyUC9R+jzW+NO2KeJ7ylYFxY0NE
cT0yjxboprTqZ1A1a98X9PsWMlXUNP4QHBOb0hZIKegcN50gETpHdiWMSPgScBr+
BMjjznzlPEFWDBZ60jWpWWAN7vRuHeshuPeTIraTL3Erk8u/ZD5spkyxJYneTmO/
cn8APO9Q+b75GyhH6j6F5lfaZkae1PnW2ZUUEWiZTDWLYcvn8/lYqaOJt9J6aq7e
CWN/et8n3lhl5efsW9mg7xGtvVDCu94b59B0VQGfy4pcMlJ99Lz99kxP4DE4A3m7
RiPKhNwQHh4OptkJb40StcHQDaY7EOl9DxBsRUAgsxrnbOd9ErPL4QwCdsx/vX3H
/CHv6NUEAtoJxLvwIJeb8y2IjZtEC+DE3KNbLPV5tcsy+78SGKGTaL1Jhht+HJ7t
zHtjXp+M290xrEBkQoy9jslcMaQpls1AP8RN2X0KqBJLp6qb7pHSiDouvpUpF/yy
9GUgpeMYztduFK388mHP+gqPPFWRsaHwduayBL+TCDgicCM5M/DJKUB31pVKM3y8
Sr+GweBv4LilBIXx+0wlT+dBtIg65gkJaiFnVj6RGYfxyVCtCkFjX7N+onFeqOdx
5PH8uMcASzie0hj8uDkZQLAg+S4N8hzYSfTSHHFCazJB8GKSZuQO5eSyLgY8uv0D
SdO74Xx6Cr74TTiir0R6F5h81pTfHdqDw2spulNXTlYYyRxZ0YNYs+oebrWhRTdY
bWKIxQVqQKhFLSP24Hbpfgej4nAPpQ3mlsMKY7kdrQC7LL1RpiX0ZPmy4lEAPhW3
lVQdSOteJsDUZGEXJ+RhpyL7gS/eMS0AGhXEgqZr1nxFb01jqtNWkNCldTkf/pLr
99Bp3/5UmZn8Jg31gdmABeiS6bAo4NJoIrfXqW8ZJRYXBZv6x8KvXzS5ZHzJqpM4
`protect END_PROTECTED
