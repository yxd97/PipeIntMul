`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kzcdLu8p+KZEzxHOd1VJTuIAQH9EGhPYaIgofGMhaP1VJ96iUdCbJygKurdFVUby
SQ62MPx11NLVd0APt4vSfA6yMwbnq99FppYIR6U4R2jUYS61RwIDAjwLCESjhZdP
NamMacRWnY+cGdrWXuImqBIvNen+mlTsz3F6e1ADw2AsIQ3PQ06CI3pIFmEh3+bB
GKyRH7tgUL+JEFvQDg+cFQpyfT1JpQ0QErSGdwHGpEWrrVusiq6hjPYigqPaT9Fi
6Fx2Ba8AN3T3oBLAkvO0iRluOR6Chm9mLwKK+CHsFQaNFvOxfHxwFffqympXKL4C
oOJI7WtSoDWbc4w1+yE7y5bJD+eMoOWmbW/HtkS6tYU9UGn8vUQFI5cOE4lJPuzh
l1lau741nKcvDc6i6vCrjouKttlXbOCaDQBZtP+Ax5p4fe5yU5+EwOQqylc+dRFV
tK58GhGQlO3I/q9vaaK7fOB627N6tTU1NwUhzNiLP6FyNf00jB92dPr1WNFSHtRp
6S1Myflu4rpnTITUcsf+TZm36L4YierOL9Z0JRqw/zsuPSZGWaKBpwsvZmV64pjl
En8yrAvxcBR/y6DQOel41x6XyHEEEG3DqK6fFtjD7c6/JeHoYC7qB3ZFrMiEOQPd
FbzV/+pPW8TbD33Jmb7Gl44am41AG4od7vsdEdskwtHBvrEmh1vGs/CxnN3TUy9D
R0BSg+mwK0Hstlf/pvo03KKkhGktxlnO4xOGJkxrdVvyrQk7HBWZL0oxxByVVfRb
xsODUVrwK6DQN/GIrRoaO4NmEq6ZlIcyfM7jJPKmvoPVd3gRC5Ks3S0dL4Wb3vqv
QGyX021om5iFADGUoo1lzepLIpM2SnkFNitFT2dC+jxePUuPj+bYFXHYUOrl3GT+
6ndfxefUMp00sSjy7z7vk7Mt1rXKKQz/KzyUH7moCq3lGRPhk1Nb4TfIZNAzyroN
oz0Opy55bf6Ic7fEC9r0qCzIuTA85ghPjMdLAkxYZpb4U1MzL3WwDmLjc8wm686x
t7EVomrLIULsVicUvKqxVwNejzVIY6OvZmbs8Vpw/AsxRLmd2DsqL9M7aLgpYZUL
E1zOWDR0ZSTOQcxRmTkCAAj/CX40wCsbqRXolXJWdDjbvSdXZmc3cMbMXJimpvpV
o9NG6tR9C86ccfLtWCVdbX+V3ZRUowVMc7uilbiKqbtvHMsbamD8dPsaUc/sYeaj
x50wUb5c2cNvazmUJKh4qRiKbyq9zdqdlurUndCvG5ewiCRlKS1PlxDWGBzSIxcx
txrwy0g1HOCSMCBZ4nO46EZ2wbuYNOqkC/kd4h1LDXSkHWb6vlVUZXtVWCs82oaA
4u5LIlIBgEZ211qIaYOP7vqXz848DHu2tky8KP5OPOqV7Fx1AxhnYadpmCqvI0IR
bioHYEVv9n4YrXx5UpyO8T1FEk0ykvYsMoQtfTVAFWaCWbcKm4IKbJnZX4qvAKX4
KzqoG14C1+xivNKvSPPt8iWnCSPKuKLsU24BQjiBEGVlzNRq9CZ6qs4S6oTCqCHn
25Z4QKkOdwdey7YgL3B7Hjoadz38wzMTEzZBlmPP1p2WOlDukRNw6fdFljxz+aCG
ikBmYkmmZO8mEV72WTUr/Z4wQQz9QQlIj/M+zUy9ZSzlPxiYzfylpsG194FEadoO
VWf0mxYsNGLAtVQ3EEL3O/PDiRCBN2Vg9TAPSyCxeE+Ke/MVsJp2EpxBI2oUpA+l
JHT5qv2kFKWhxB0GDARB6NTdL+wAUhkJnIY1SnjI6wPB24Hl1lSgVhosKTqX+K45
YZhF3g4eOo6fsLvl+rlIs+Abw0mq7cmoF2q62oAlmtLMYNg3gdTra4famuhbXq+Q
mxIcOxlrDI4J1pk6qC1osnWkFOpJjKbzVgfQEIbV8kFaNkVccVwWoUJ1INuTXuzs
SkjcXTYQBRoBGsfEin1W6bRxJRBafFBVLG1c12R/rFY6+VKAqrXQzTZm7RBMOxlk
1vADOryLsQhUw0ARBDCiKQ78s6KYC0JbGoDG2CnEf3kuF2sxCrujkjkW/qq3q1fQ
y0i0uaFi/OD+REg7OQ2JsVAN0geEupptDZBPlDBQqzZRdmxzQv6O59+0rehFd+dR
bt9RYEGbJ0K2ALaCZOKCDxyvzpGN4RoWd8Jzu0/BLCQTp/bA4AItCfFCeWSJ/3Sd
mxeW0EflOETPWnQ7eksgLnVhIdzldKAtkE1lbv0P1MZYgwOFXRPdjSJSOiVGzlgF
BBwRgdPQr8R1n47KZZiuEWyzIKwWEw8342tSU2BOpIcm5rPIsXCwqPr88LVU+9ey
88qQ9Cy17irj2pH4jENgnzA1Q65gEjT0ohbKBIf1LKrkx/wQL0gJDPmE1641UVdD
N4vgQIkrZnR7G50bo9ip7di8DLiacVj40nyXMPhD/U97fgiswidEih63pzwJ88nD
SnZaO0AqHG2AWn4ptEFXl5578x/XH9jRpLEJxVjafJiJ7nk7Vr2AL+fBGhZKU9gH
1So2dBLJm8AhaAxupmo+5x9DfWQrQbKiOCQW6BqWmyYYbD1MnTz6sLjf2wuZRXTi
FWMqbjEAHL6P9+J1bF4UACunKH9X5Fn8H23IxjpbtmNcFlxaeFxLLJ/YTG8tEFys
dRQTevY3svZkAl7GeVXed8NPZxOrKuOZ2jUIK0hBLpUdv4IWlyvt5zrxHI0nOvZD
SyKBkeux/f8jjlXNy/wK4CIFstPnT4Ggf79GPGUCODdVuEZepv8aMepjGHADMYJ8
pqt2sOu07GKbxW51pCvAagw3aK78oiXpGAu7vqEMpfiYmfVzpptegdhlmy26xY16
2KUryKdegjJyEt+mQbDTz/JRg2iFezUWDsOovyEjhiwppOe6fIi8MHvT2W1SD8OV
ya+w60TYfid2kWSuPjFG5FFY6gyGo7tJqpYLxSS3eR1DRpYraQ9i9V89/WU73Xdj
aktKOcUORbv2B8SbRJ5aGTxrTGZ6H0AD8eV4ZuRsYVsCoVpIRHkhsTSEO6eIbSXp
Uzey7/3/ZN52BF4lFWHc9lod50+kegr/EjuPKqwRcEk=
`protect END_PROTECTED
