`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkj9h9uw7tgGevAvPXMw5OHyy8fc8uy24yEswbN2roKyI7kkdW7A/FsDa1lb0Jwl
Q8sisBMEn0PHLViYcd5xBXBU+EWpqIxas/5wgFEwSP8ObnYFp1OqDD7wXJTiFamb
nGpmDqxJCEISYBxVTFxvxcMpnDgzB+08EwsVj8cbhvWNwvGcLsZoC4j8Db6CF3bE
uTnTGrIMbDqFzrktiCb1BWImP5p1HcItL9vc7fGvt4zL02Yi2d5lpPC96zgpHd07
Q0+gRym4FoU6/dXXX7ivYjhHTC/rqJXl/nT5Z9ifPTwq1AtCHC4gNZknVzfAgLeG
2iMqFM6Z7owvjLhNUj74tyAqU3Rne3TO6PKIAE7hY/BWmpwFOsW7OTQWf5D4v7yY
yhUVCjAyxPxv8sxqfsEPjEgK1sece8+GgS9Cwxs+SwN3J+XlpvLkTPW5xVdnKLg5
oNId5QocZi1vpBGimvxtwtZ9uuGlaPSSXV5vlriS8tFAtLdcivozNVVMh2Ny79b4
Z5ZYa/qYb3dBpoI2sdSkyt3f+03F/cEIY9EsB0cUNcMVtOhGRmDE2gV4b1LNfp/D
I8UGc4dd1UTZ/axI8czfZhCugIeQvT6zfja4ny6BseU=
`protect END_PROTECTED
