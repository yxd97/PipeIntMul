`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QcPUgQy0tH13gv+YTpi0b1fnT1ZJg5YdXLig2WBi+d5ibQEXNVSMWncZ9YA7w9aM
iUniR94YHtwzlwocqHYhKhcMgCWrdCydyJWdQAxFBExWZ8a2Ga59OWxjwPhlsoTw
CHgEfIeZKsh1akLEB3wuyUTpGrYpUv7YS0DFc7wHabkyL5UsKHllwlf32NI06Ph+
MX/xdXOpkMo/vv1MsNoPtcClkVXVYrJEl4oS2u4AejiOJ1k+RH0YazdIddvyTFHH
f5oCf0/uc6nsCBt7wTu6bqNn9wyBiej4QHQVXsc0aukZE4lQs20tTBAFnJ75JZh7
fcxG4p7L1BFNro7uE1FERhsnGlhI5togK14I4r0NNYCidagezHsSoNKmdURatWsd
52UkLSAX1ikEroc2tYV2LKFbo3E7cjXNHpy+6RYtWw9v3rXvfhzRdkjm06DJenc/
`protect END_PROTECTED
