`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BV6/WIfkUAn5CuX5O3Cy+g2ET3Ff6p0CYw1p7N8Us40k83gFgb3M2I08OIQrsba8
IL6NUWSb4HslrERKVxXpcwIO2aCreNCgJViKTa5p5gqynGYHpZeyV8DuP0DNfgt0
/9BVZsY42o0mJ0f5RavyNKVWpzFy7qOmU077K9GumDriLG2hi+Hy8GKGqbdzSHka
AVORHSxvO80ev5Xv+XzpTnxPMP/snmm/iJtvbn7IqPbDZF65wbxJBhz97Zp2pmz7
lhImjCpwoT1g9A1LCchAv9C6qOAGpMkm/fiPV1nboksjOsKsmpw+4zG9ScGtpVYJ
MGPSYHHEBv5wZyMWb0F4ujqJQNAQNRQf8BKn9bf2ryV+r46kSbHq58MFjVNwbB01
q8huLEOusDKTZtFhdUe812BdynCVqjgSbhg2mjSYB8wrfUUAhQ4Ljhr7fm1n/l9/
jeOpW/IPFY4w/aaIheWnVtzE4xvV0l61r3dwzmwNzOw=
`protect END_PROTECTED
