`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9eMzNX68Km4SD0goS4XNKtu6kYp8+8g9bj0CXBv76XvgPaWXMr/6A03c6NPhgam
GLYc2R+KNLmcs2blcsOeA0/DRqq2/rxjO0CPCv0JL21UBeo8PdkemVOnNH3ChT77
XcEgqi6GhOjkUVMuUIFx+wRAITJ9BOkvFqOwFRDYJwU5Lw+k/+uKqan1WToS35Yh
Jelxo1oD69YtivNVvQ6F1QyOWnfazMxGQI6I45MuzPrk96p6NHt87t80rLRW2nKY
oVGg5Y4bVZeAE2YK6wEP/XoZKEBDQgDjaoYgywuNqeZCgEHRHpkxSBTD3C4UJuNs
qxSNenTahfqu5y5HrGSyei/qmlcfXa3jW7kLI7Y+KcTZLPmZn63vBPn2l8xMZnHP
S8Nn5jLTvMc1prXHyKlOPcVcPHKjfm50Zr5UvrenrJ7fB2nSL0ysW/IBNseRidmw
Ed0dFoAeLtBONh7DPqsYYBkJJ4hFqo0kgEsfHATUVTTWwHqyGlIFwo9OX/csaZfl
Et/46n09XVvnYwXmfvK9WfmkRIkp+pkrClYJfimTIzdUGcxHZAumrfTPRU/RbLvk
y+w/0vD0KrKeETyI6SLMkg==
`protect END_PROTECTED
