`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4CGSjvIKATwwecxT8j+/SAbh34ZwBQKpv9EJKlGkSA9ScC6Kdrf3PxoVt5JJusoO
2H9dZSruJQM1enor9itWFISsnyTk5R3oR4sS6Kw1JEkF1mFasLAuOTpvCv61ILze
g9xtrA+fQFeA+AXaj5cctn1nahqQbVqr6nNyM6wI6RheN3NtMNf0mN9AwLS7Y5FS
5bE6fTvgxqHHpmglBzZ+23HcgBkw8B3pxvPsGwRnDBAJtnge7RH5DOl2ZTt03M7B
RguXFO/csB3TwpagCrGTGw==
`protect END_PROTECTED
