`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzKWv/WYl+XVvzihPDTl2zxV4RLJxlqcozh3iJOi6ALrtZpdRM/wGjMhncfbPA/r
28oktPVTZa+djh/38MDlO2juSxDk21KAQOFBiL4+9XNeGGPKOoUteaGqT6UW85ba
01Fsrj58qN4Tfg8fXQYfkrDt+CHfTL+s3POmPo3sF8xaw0C6Cyj8bmCIjG8s16ra
0s/riG/FyyGnVinn6ry711Pl10khnlY6awyFNOyViJAp1MgUhU+AAwEy+Tsd3gME
mr7yL6syKa4VpRPGAurBNXu2IPTCAbg8HDzRt6ztIPbLCubXKNlVSRb0Kg9b9fXT
v7jZEOaGHEMDlfAaeqcotg9sqUug9kUNgZl7kLBGQYaEJcHLOLx9L47b0sY4Tjri
z5kWkEh0xV4BLzW0jf3X5ew5opajmRsbzHII+mnNhwpeHbHCzxNoWnqAk1YFpmxO
GWxOMjWubd8DGwfpvQcJgwSvM5ZvwrLe33zZO1EqYIq5cxP0KeziseEoHie9w72E
+5uKJVVzRVpaVv3QVIjMpmyHV+oOMT4BLCPPqvQ/2VmmQsi0OUkMeAAFPIhP8wWN
0uFxye3Ie43A4ClFzh0SQsHmwVada5OKEsu7LPk/4Nm6yoYyZ4MOHe/v45T5tu1L
4zNJjCaFLa8a4lXLFxTJydjTUACrXlyjSvsGAX6seDblo5Ho/aCT2592/FmdcIGt
2wbS7lM8RvWBGvIS+TYP9ZC/gqIp/6QLZ7W5byX3v+8LU8eXWeIKH7XHFyHtQ6k/
yuidNU3rJSNDzjoUeJR2iR6Fis9il3YAljil9aYY4E0OpJ7/DPe4dmSC9DVd0R07
BuEVXav9OQs21Az6KhCfLA==
`protect END_PROTECTED
