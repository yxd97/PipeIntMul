`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F1lbAStylk14c/yOkDMfkO6rgfQggGrdDbNehj4lnZK9JH+wmbskz93v7ljtXdtl
6Vfrump037pCBXnt2zp9B8cYkdQF0NRqu1Oq5jrTK8tohcJx2tSHf0j0GEVOAQL1
JvP7BJy2Ah7DDwY95KIrsE5XDa11OAchVRtw/PzH3EqDo7oePHNw98LIxB/Wm+Hk
tCSGCikOLKHaXL3wKZTpBO6a7zabBGgc8lqc2rlR5p3I7goIVMrLv91RDMghT92P
8/qv6y1wwx4sV1AhmyoPT5sRxd2O9KhJ5DTfle02VAdue4+1DLG2YmonmynWqCIW
mppGclgfyRdVzXN57qAumRHx98JKrDCf8czJNSwsSGci2Q3woPIDDAdKHJrHs+Aa
jbz7XeYNCob8axjAMB3kHIo9l0clGXeYm8/ZK3I31q9qarnRXL7ijvXnWxmFLGUB
Sd/PuBKQ8kCsLYRPMbTt1+gtiH/6NhQ/cMIOaxThnM7UEyHdIongxRn1LlKeuhJn
L7DaCS1TNaCB9ywNhXF/0k8afruLVE26UMmwv9YT8Au9Yu5ywMhy/OwpHX8EtHSr
Ke4ZJ26egaTLiX8Du9YbcQzGfXrPTz7Evx98LAPR+4WToy9oUN42AQT2YOpaSvd9
j9ko0w4mOhqFAunE8Iz7xeIT6o11Pt1mQaBQPGCHEDwDNH3fCfhqch6D2Tul+xE/
L7i1RsJFeDzuWRzcfwo/netDWMUCFPWA0Ejz0w/YeMbwNFOhLn61jNuM/HOiUnxT
LVzVbrc/q9wq8lVY4tb9JhaYUyXAlsmh32+SWfBc4LU+W0TgO+DCkVedgcTdjP1k
/IDykgOFDmVJrT8mHuCPnTk0eJwYjbki2Ztp0yway2A+04LW+aR7UD4nbnCSNec2
ZrzxunWuEGDr4kpypOwMFOTR9wfyJoXkK8/Kh9Fu1JaBa5JCVAdIt//g8TqmXxyc
+DjveCxAvjaQBVajHnLXHisf1l7gRWEtXaywa69ijgw5C442HUUPpB25uywC4+iS
AxhYdbptcPfBEj4jUMPHBWDwFNDECAiBJIK/dvInw+HehrOwm3U34ewBjgKZU+F+
FmmWlW3qAoW9Uh1VucmeXGrOMuNQhFcpSB5Ye+Diqtf1e/TvU1WoHS7Srfgw3Xkc
NBXcDIfDx/nCYMYd+l5EVhtB/0mgPstrEpziYLDNuSRk7bxLiogrRZmj0z65cdJw
CHX1o/hnm7EFgmhyPfZrmjqfpbtJWjlfElTk2jWAxq3AtYAQCZB4Xt/TKrCn5xKX
ZPraO3JT6Uu07w7XfZAHQs3Xjh7DpAfVCxjuJRpnJt+bsNKJyzScW5b0YekstCQb
zBgTmhUKyHdkoIFBli0JCvXS+kNZfUT/Gylb8IPMJNF3H5x0A9J2LdM0Sf33J77t
hsOctcD9SktPItoelAbGr91klvffYAln6gahc6MxQFdSFc0CTaZ+e1ZW87O7edt0
wCz13bSmmb+JoZ0s/4+ngC+fe+Esg4Tw0jY2Q0BlglxZQ6EuMkMQ3X4QEys7blBs
2kztwBg+NMxceaMHnMKfMsC6qwhSdqr5ekBFHjvVw+sNgYU0GK4BWEJS/s8nIvOn
dasl+XF1ugztw765o9MKM0v7GOR2ZUU+Zy5MnMtDMOCXxETOukvaRA3DKvaCIFMO
BLfNrJ0tNq9CBnkJoSBYXooDb9X4pwLIopcCaiHqOyqrPs+isDa2v+++uofrkSBe
cjVlqezxJnEuv5pjoyj2Ymy01Jvba4jwQGrp0JQJIhmBEX0kC2auKlqtpUJ88oM7
mCClpwgupVuhzzLujueCpzWHUalCuvo2GGbX29r8VmdAlyXJKYkmlg6Gl8tAOtXm
gPzZfZulKd9gVEVTN3CMr+XUHggOh691iCRenRNo8gcjNxrkECHEp+qsOcPR3aA+
yq14hSx3e5W8tXsElBhgJ8L6eYbprKXiJBOusPFaWbqMXEOKth/M3XWfRDvlivEg
BT8jMS7PVAkEBNRdPjP7zQviuD3bJ8Wkgs9154oPfzY+NIz/H5vcjE5OKD5W8/4m
3mOo7HUTJx0eE8UWA4QmEBRmO4F1AEkT5BU+zQSRW0j6XOEbcdjyGtuoMCGUH+tv
rXMDUCO6Kmtnch6l/OAuaRoXNDkiq6hhxDlriBVVwDvI8epQttj1/qdyOuz9b3CS
RdHBYdPsG8FgcNqi7ft0LSAv4E+uWKDin5a862cOiee/10BoUiM6xRRdSgojaGZx
3GY3lQyQL/ptNVVKvdN/dvIQZRcbt6eGFvvdX9SfXs+7yK03g+54vVyb13WQk2IS
Re0U0vH8zNHgN6tA5iMwGxuGFRsZh76468OqxRQwtp8z4FTgNk5NaIcLeYrypmHE
GoLgeaVq159ScKLNUagkmO+X+iOPYZNRKlNC49wjkNTHDP8SrHJQcvGMI/k2J15M
PG+FW1WvoFf3ainkI6DPpqGGrCFaxf0eiQkALAbs/k6hOwtIdKYB8LPgriwYsMTQ
RYXWuyoKtaVYkulrz0fYCsq0jXJtm2LRQMj7OABr5l2nO5mEm1alYeM8n1GLj2Vn
LPbOWQSlCztlHbrgi9ehcFFuCMhRtC47dVt7USeJA7G1AgmAF6kgvfubhdCV23/c
RdKbSaTGz75V2GJBkR875kakFpCvN/nLIo66v2lIdiwJ1z6Tt+ZlF+pLFiFwUN+b
uCsJVmeYQ6PJJY7x/racjhbqWuPtayIIiG9MOEwpGAJ4MuZ9Ug4cK0GZC3rJEhYo
c/zGcQR7Oi2rrBxh4I1gZUviLl+AbTpRCgCtW4Uu6RZzZqriUth2wyJl7mo81wHC
g1/8Lg464CplrhNrU78ivHGD39PENTNW+48ee3TgtdKO/AdUxVhYTPDhc31BI6qZ
SbRYgDgxk5+VaM3uFIbyk06v5+S9rqBXOZ0VMZMWqyyMZZcUYzm//z+fu0NmgHhH
+acVzc6shthxdnX2bpDi5Ty8b6yZ3SYE/XBynonBqe1csPc3ucp8v9CfpoydcpmT
72ErYBBXo+k4y1n0RQ/wCsouGDP/e/CFENe/XgkkyOf2A27PoM6yRwyqnynv+X6s
vMOHQ3qDO0ckBDlfOP/eOmqyNqElKxvEg+Q8OTW3bh9MF4b+6YpKV34Ma7o/8EKp
ThLwXq4yWP9cyF3pOCcslfmu3ih0LlFfp9DsJAx975vjOYKezyYm/myqXtr+j+Dq
GXwVgpVzHlUCbwoxObRdQKvZspf7kABF3XRPVSXGyM5bR6jDadSVtyrFk/fajQl1
V5xx2lm2GRKnwI+6e5qCIyfBTbVNOPYcREkgNaFtAR70xGihzAo3O7ctzHIv4VBw
5xzwEodNdm2ZikmexEYWNodJaGhyfVM+vdriAoFWY8dPCee0qRqbKOkbsaBsFmMR
lPl/Zx4x3totwFyKS0dNGBazAhHQz9dcqzGTZ7s6uP6/jjuy6JojyqhBoY/Bk5vv
27HFIJheYI1I07zRSbpJdK8ezkZgnwX8U2cHgkhohLT/N3mEo8UVBh6s7zmA1l6d
w61vpiNh2BFlUL6MZvIwxmRVvEr2FuDbxCK0mUgV3KTm0atLCv9+N3PQ4XsESAYq
UNJeAvLeMJucUafMJiu1vHzJPa/NGW099Jps7CwAW4a7zJGq+HMmof/e4C0vvIep
Oc0ZlLqk5Q+h8+eXW3dRe+/Cvsa2NZLndAEMtQGkRiBA4/kqvJ5KlF1ytEWGQghc
ew4T+aG7BTo0w+q3dto3fZG38TWdSNGWEGCPcVy0Rqf4cQ2cYmbKXrZaxr+9cm3q
77DkvKh0rd5gRjY/Se9jyfAKDZBzt7itlQbVQMh7Sr0YHnapBRagsMDcQBqkmCTE
dpJ+CX3/efZ2z5O7Nrh8b0yECG11FXVxohgoB9NlsCM9VNm5hbp1ts/bPCoaDWtx
YQpH4i4c/AffLnzTlql6FuDqhjm91QzvkTQEwq/6XdDFf/4vZvbEZXcjZCD40ipN
e7jHcLAgPxKAV83f+ez2JFUDvIH02EfGHJO9MABQDot9hhUp/hTXS2dJDv9IEy3E
S7KYSSdQRIKaGaMCQQkWPaHppfNXydjOTwPZPC94Cg0tLh5+Fr5h1MCfWAj77ShI
x4IeeJLmrM/NGivOlZ6RFxY2hMsWd4wl8CxKvmZbr0OKVTT5M/a7pLUGVX3cH3Aq
1BilLtfdEWAJoi46F9+RlHUBt40K6oiPe1mi0vVZTcLmGFQ5P3i4mel4omXg+3x9
yBiY4aux+McTDOMwJ5QnjE6fi7AkEfrK+JRHdpQg1DOKg7KmUBCctNDQ3TJ+eGQD
myfKXPGeaFnEJoYI0dN2uygBLvuyLvtxfUp2ZFHMNN/PC9FWkMMHZjIJYV/3vhyM
n5/06m/n+2KMk2IPKQV7XYuUvxRX30mPO+csqmYUqMY9gJeNbExsTG7ukk/GyulL
BBBKaBrqemfjL2wZZJImAKzHhvK0aKItC99C+tULdMcAdJEPiowFnHsEMde+J3lQ
OoULXjMIWwbPpxZ7Mq6V2fyb+8Ci9kuUtOXjYl4O5CtMipbQRntJOxMGnIKupZ5Q
B3RclpT36sSIKoDlyhh2v5YCn6evp1i9fZJPtXBNDyvoecIq0fBPK4hMlj6/6+fj
UAeqJI5UHKy+rTCjR8U5/sDgH7JIxG2nVXvXpIq85sSBOJDAIIFVb4Mp/a6UgKyq
ueRCzy9n6KW/IzbMdMZjo58ndcrp6B9gI5TFNxwVy1qSYP/DFYRPnRHdUrrgknIo
aWcgu9LtQqB1QdCXtE1csWQQ26Du6FS/c/GTEnYTJNd/lj7fldpE8Xbwa9Bp8iEy
ZpSsC2pjuLz8C8WiimDxRiCLRZxdTDm8hDFfHaByF9ycXr0xrn0mM+6zLaZT1eFP
eqEkT9TJQ8ra+O22XT5GhDnhzQ3eJxR43eTwa8rb0J2uTdsVK7rcH1tDv+56Ue5t
bIH5ylqeOZot288C7Xm4Jtd/I1dT1DUwz21ZfJx9Ywpeq/QMOIbUv5XZePuXwhK8
UeHRTvoTgESpZz/ygE9ZHJ5MpTg/bwlgz/gnBongdUyvQVZ3WSiWtrYtMSB5ixA6
7LwrcRBMLNHzVh9hshN1Yy3yVINb09ban8uO7BxnC2rVm+HWQdStITZTSOQsdUTY
icxT77MRDIF1pRh/FpktY+guP3IST7BMhFjs4gVtyjjfeppB5gOK6MmSAku/n8Zg
0eNcT6QlKPMhTyWf6xTjYYrUp3K7r5/A/27BhFkEMAuuA7EM2UcAjHerjOhx7fN/
8TMB/SAyaUO27Lw4YNCPmK/JY/dBgTj7j7hUb7CQHoEE0ek417JWK4RwwkVE1mnY
I0TECPjztJKWXV4Dl4DnT/R7ALBchEcMU1HR2tm21tk8M5MspmMBfaY9zw0wKVw1
NkRrFm9it1IrnlEvTCA434yQOhmixIAprV2OTZfZy0JEU+VBjYqfD6rLkXhXuLX0
DcDHCo93gB0dYCDpJwkMSpAtDvY/Cz41vAfuRD57gYWVwjunaSfqV+uX4jMDSBmI
L8oWQEPWE2jJ5Mi3Qo/VQW/KlYyFsue2zyqUOUog/JKE2pzdP8kdB4M43kV7W1Aj
gbv1nDP7ZS6CNcm3nfjXEyGIAgZ2HJGSBbRmMRpvtCb4x85f9Tjbc+J/k1fj0ofr
U8cTuPq8EK5rJFC1I5x8PmjKeLBL4BCYWSniyfS/Jrb61FKZIokVyibQ3BGJN9A8
dO51bODTVHBwTYojxhZpsqw6HQmiax/JkgBLUnl42kAWsmAxq5ZWxO7i47IPWpcD
1N36f71qnrEOJZGwvTVi6yUboQYpNkyOQkWkO+N9uRzoWH3SrySwQoG9CMAdMm6W
8dozTu8EwOUvGoz2c978PVS/KbLD/PFfRxClEtfcaYFKVbyW7sKSeB9Jm5RJq2F1
GMYrY1oXXBIGhUttLlNJ6y/NUudb9pS1610Gukt5jktIJ/dB9Zr6F8bTPs6mwN7v
hNTq7CC07uFLe4g2Gh9pRdej9kPScPWHgU/8mjijZS0PROCQooTwobyFXXa/ciK7
qEwcTRjI5cqVeF8YqaNMhvqOuHtnjCJMooD8ajvBRwHobZslkmQpSRV3ULfY/N+D
tT/WNgItgFJ5cOo5+Ai7SdA3FjRlrNpXoTn/SXNhv8znySJ/0WT5lr/4EcKxHynK
ZODyg2s1mFLwWn7JZU/rDNzA0iUkLzP/jrdzN0KKj2vbpTdciTb7AW2XtGcQuio/
LHQKQX7y1MFoGzxiIYAMFbTpKPjJCPIDNzCJVmYG9CneuxDEb5Xx9nZsIKGABO0c
ep/NbWyvl2Qm8ZRGo9HOuBEB4CCUywGiyBzJRWZbHUffc5va05tXUIVurebbBNP1
HCSACYUg60/hCgOZwuAQvl9H+ck3NimQejtvXgpGnDHGN2DuK6pHxYfMuoa+/seP
68fdhK776PrwmiFI22PmKUGhdbZHNXprBSqJekBHPd3xyuy571+lhdR4shHf+IFA
QPzLJf4K+tkRXTRanei21bYaON9CAW0UDUTQXiPGcTCT21BBT+irc4rmu618Euwf
3FEB2WdFC8kTZL/e+ZLAbW5uf41UlAwb3CPZGBKi2QkCh5OC6CQQBCMebaQH/O7B
3vDYT93Ro23b4i2ayRZpuAFsCpvsBKHyIwTeKoytNOAQHFvr5zqH6FlOlbYfCAED
L8/yTCxqZPQZNleMtRPGxN+xfsM/4/jCJQzj0B/JMJ5JC06FvNfQS6RIqHy0uhL9
RnsflLvT0cJ8YOoqnIb3M95+FNkrwU+GZcb8lxPDl5xLXJa/sXCK2ZMfgNfpJ5ND
v9LO18MmXEFAqwuEeZjzUlFHhDo3Y9e8ueqSaWvgdNH4iIWPGJemIZ94eCszKzHJ
90fBFOGtccOjn7Nx0LqAyFjpEjr3utIYpzN4ixxZrWlabF/hUWOifVI9AUQlFzTV
eGWKLkb3G/axUepV2iu2W9NB/d6MJLb5LNbdpTSe+9hgfRhAbiEhngzwM46kdZvV
eqfNK68/6BgJnBA5Ul9PO2V7SMrp2YqtFrNb9m4fIgGFJTq2zA0hpPI00qRokAEO
1Y8PYEUhRpVfeEB6b/HAe81uGjWOtwJBIJof2VekFs1ry+D6nwsMC+sq1fwxjLr3
N7uN9Y2neEwpt/udHB2lB32JL+DWM0fhZBkuNHNhc/jbnkzn53cl56XlxGi87Ce6
uBaB59ROPRl/iIFS/VVgEsvBeJs7Tb+cvZGaLl4uvupLkaeWVJ8ot5jvfT8dtPnM
ZqbwioO5tuVblU/M0y1X+mVMnsX47Ok9c/YfPafkABcR8xP9r5T0RTOo8eyS22Pv
Jog377o4ZJTcZ9SSOr71COWxJpgcgKj68c8tdLHv7UPoZAz9uiBovErgceDcWzAQ
7pfFAoCOQRhsjERNVvOtFuEfK53xrKzqTo3K1muIZ+jUqPyjkmnOpM0BM23YYkrH
2x3P1OfJJq2uZhhHfHcrBf63Xjt0BskIAyP0BgNgpZSlWTxZdr8VLRlYPk5p7Tmq
eYksw0cj+aGpY9FH7E0oOJyyGDVuin6RMl+TfeLqQSSqm6/GozPWpgbbtqrGhysv
WZgm+MMkLEnkJ4ijxryDfDs4a8pKIUhLEiHNYfagCHPyTUoPGHy6YnI2Fbj4lzN/
jHx/JnBPjyf2NQlxTNkE5njVznV5zsu+leJ36uyboI7hznjvJ6pYIByBTPU4XfR3
HeTRRkedcTrV7Nyq+sT2BHUEiYyNAmDLOgVOSRQxCgbnfLKyeSsghrUMzR3Cj8H0
CNHEnv48e906NtWHMdW+g46Mc8YqN9y4cIQdfAdqpQb/XcHSshJgmtEpwcOxmgvG
u/eK7tKYfmmR6mytTXsQy2nrRTeY3HliuAnLQ5//7MOmmQfyowJhbJsq1D1hBxrX
YGm8ngmIxgQpmSA9978vZ8wiuOyJ2Jmz9Ox7RSZlPKvEUUkceiWIcbmbyyx5lhvj
uoJpdiEKKPmPM1PgZJqI4tffXX/ExF02VNbI4NcwCp3hRKxoPP60xNEnxaRcKBWs
XjHtSe7kMq9CeifapTSbeIpTlU2E7Bgo9Anj04bYElev1tWiAO8Z+z6sU8/gm8+e
BAlWc2F9QZw9xDu0B+K0Aw+W3Bf/D3fV2o9u8bVurRiiu8GxhRsfnCPdB4z30DJo
nyOwHzQSw5WW8npJ0R2Ki+4dsK5I8m8WnVOZbp0b0VPLmLT9bw5NiCQTyNXF2WBl
2QNiVQYoaYDPcRKFD5+WkLjeFlnWypOk81uI3fB+OvEXLtg08RtYny0xqtDRu3Il
T/STgd3K9ZBtSAWPOSz2rlGocnmPL64/uzc2P5HCgKQkeV/EVwx5O4BaUFuJN6Fu
ASmAsNfxxFLR8v+vRycEjif21PI8qBjL7SeqhmxRrAiERCdRp6nqktcsrETTV4aZ
oH4Rvz/qrZHLDoDEhv2NWjiZFbKkMSlIpNGNBCrLUGKISqGVL0N9BWPG42mbboHM
nb7J6CNK+w+5uChozleWvBjv3OYM1dhQ/Y+RPlnoJBinARcA8VWTtFhkf28f6IJY
`protect END_PROTECTED
