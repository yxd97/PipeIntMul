`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bx2xuwdni2X0170skAtTwoF6GcfFm4XCoIUXGxWZejyPftLH3dcBYy3Q/eLHfIRw
Or3hyCub+iwyjMKq2pDA4VrYeH5Dx/dzPA3dI8EucE4IISgWXhOKa4Eh4Lq1hxm6
GnFxKcBJQeGJA1EOi2ieznXysXbge4pw/j+8nHqEpvIFH81onLh0jUtjuO/quI/t
VjFi7MaA9C4eruIrduFN3lJsG3Y5IXrQ0/wFCj7r/LQd+eObJKcnrtAvcePzBx2D
6D9pnIiNokgvT72fOMCrFg==
`protect END_PROTECTED
