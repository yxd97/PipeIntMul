`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czkj2OBSbjEJwJCEVZZIUqu9pAU31VRkPBB56iapnTn+YApsdWECLEYtxH6aINI9
urqQwuM7PFkawKlfL23KZ6KwxJqHRGHO8pv33/fPkwOAGffczRIag+j/S49aorGL
8X3Y9f6ZGamOdw7Zmk7Nd1970JJerjBXn6HDKoyEf/FH4bvp6cZhyXAyZrVEhMaa
SxiimKyjZfaOgKsQjRHv/J+YZE+6IX4j0utDMNv8suLX+VHI+anwsDSzB+bNbuPJ
Q5bM4ojsK8n8NeIhWZJc+p0vtwcIfxg8ShBssghBJacQMoiod8FX3i5vhcx2e+bv
FJ5Pn8X+7X7ilbSPmz8V8MWMfMJdcOFZ6lYCxBTJ9r5LFEYMA7YJDkkaYT5BPa+G
O4gVvDDARebijeJ1HmA4riNzQPRYu9rfqhRPPD5wKyUWHGkPjB6g3ekZdBDrrCkX
Lp6/dYi8EYr0YoxSTSRc4aJL951cEC+EMGOr5oD0MOw+U1XD99aPYI9fjU40gs1R
LcskMCjmK33LriJ4mWXV1bIPmbRt/3K2Fp/samy7keN4g6i+jwB4Glg5XWLZCfOF
P0/uek68+yo9l9mI9zf4GeUe9MUAlKNMZ4sElak+SPvCAhIQk49Ado1fGWw6Q6+/
QL/AaFowjBAbLh/fILkx/72PkkYG+fz9Rst7gdBy2SKbRWPe5XlexyZWWPysayPN
ZLcbr+VhfI/5ALN31zzV82yco+AOHEQLV+2FHzQ0eG3C22JKg8faRCuvq9pWYwoL
Sar8HumNPBIyfqPzuKBqblaTZMh4uRS0qm+J4YQiozfhSsIuCTWCVdFTNyvL68qs
yVXubY0HX+rYeNJkp16jObjhAzYq38JuoAz+Bl4Uvb/pizZooWzMhpdlNSjJngHV
b3xLQUkdtFP7zVBlDwxxCuOjwePhsmhsqEZQ+gHG/dvAAINTpVFh9EpEQs82jC0e
GCTqGRdLQXZ1WLx2GaVPu9jM8RMHGIeVd5JyIzEPTzVLQ/NEDBINFu/uUzZrYOCb
3sX2Wac32MueFKgTQYVsZ3LPOm4LmyNQt5op61SnUD3uPDqZQ1gB1OBi8tKW7ihm
T/h680FXoZMYCPh0A3VDBLvV+sbnultgy1w+ERIzubanHjO5+4wXLNFhzFowEVeD
6yDpG7tA6p4kqBPXqgyJpSDozgPdx0E1N1RGFIxoy61yfcw18iVxTvuzz3GfwcYM
T1XFfuxJQjCHz3ry8g3j/VTDXztFmMYq4ZyEemYfVKRXRiy6pF3tL8naWnU0QtD7
KFcWEfMxeMlsSLrDARUXmzTZoAVBu9WhKA8KSFVsrR+LRfGAa3hl2Vsw3p/n7SEl
H24MXmKFjg/2OpgbeQz5yTkZaNXjKCmYsLWvFnsBCtY+BHbrktxKmPjYIChHvUCz
37wgcRvj9TynDB1ZEEZO2mOBiu18g5p6NWq9gp32kTe3V/ymUA2QDo1ZYv/0vIPq
quZYrkEUZH4ampvy+b2qA4MBySzX2iK55zlUOc0C/0227er6xdjYn3XJzLW3Uyeo
`protect END_PROTECTED
