`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+uPfup7br0HWLRgHX89fFRMLVPcDzTN+qwQFZ8L7jO5xOfXs3urQhX9tiETn6yE3
T4/U4LkrY4pn3D+5tDW7sZKUmxy6skG1sJIAP3aKIPLiJNE6ekc4BivGEChfGtom
oC5so6VI9Yi87nQi3RwyIIIfLAfySfT6+OHFlO537e1m371isLjiW2awYCafjdMb
wZsEh/ayrbUKi/Az3dVklNoyGs4xJUG0B45aAfZF1D+eJBhMoW4dEGBuXtkN2dil
2wKGCSYPo5qKY0ubdodvuVBiJnJIJvBMovcNud3pSemDFvQMvha+HndAvEH1JmSZ
`protect END_PROTECTED
