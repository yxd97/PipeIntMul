`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y1ICvqQZOuPL239/i6G3Rtwixb54YHH5JrWBqUNwrze7ETEWaZO0zSnIBjJN1QVT
JoHrb6zGPDmeDNUT9XgGv7jQem/1vSjJ3BqcDX7Ev6ehJu5hTfgVPUDF2tqbjkoJ
zCecMOqKdusUpLi6qpHpI0AVUI3ImiHq3+JXqAYsSK6RlLMHmCpU7VxzS88Ue8VM
MnhyVwN3Xp29ghTLp5CTlYL1E0keUpcWwAHk75fRJIxKHrZj5oMJQBD1v3od89IC
TQSBPv8guxEiAzwN3jH0up2/F7obyCHtTxYkJ4IuilLrQsOgzkDY2X3EHSwjHb83
KAzqGLea8N4TQYet/MnpHy+F8McKS0VhdO5b7+seAGXT8DcvzGSi9e+NIsTlhEV4
7BE3Mda1wD8O623peSE/1sEHZX/ojJTbJwSf2J0dj9jUHGIr4EElPFdqhB4nPMEa
sznkRlpJBODdq5tQxzl6MQ4L5e6/OsqvaenZAIMS+z42yRzzzh8BIm3yLA1hv4JI
kTkON08NJ3Qbsu+0eRwC62Q13davOGBhwx6McYAnLr7wiTvZyLcaTBG1VXCvox4b
dEvSAuCJ2vn+GA+zzoM1v1j+Mx7HoRgTCweWku6aiAbryAkpK1AzYMtTpTV8gMaC
weUtBSXHomyt9lFCKnxRCpZGswXPxi56P0JpUmOpr2s=
`protect END_PROTECTED
