`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncihZ1f85AroyiavmvEl3KOW2BPKizxZx9BNYbHD0FMS8xLCmmkpehz49uUAMyfS
rdtFafryZ/jVBxs/ZClL90LQPDEAy7CRng7SFapBtACnS9k/Y9vYzMhelNjD8Krd
8j/Px8OvwH8LOWlE9Jfvy7E8es+HnyCFaIGAG2jIZSuIC+ApQ8Cfi9gQnKP9Onw+
r0fz0Ok72H/1HAWltCvM70pDY/JufA1YFsymgMF9f8k/VJfvHZYUZDmjShyDopev
CYpVO4z0FAv3AgdUFPtbLJf9YHXfUhYv/djCtTpBcGZ1sOoawphRpQBgwTtWBeZq
qP3Z2cM/Gp88eDHXYunhkvJIg3WdwsrPAPLJ6N0MWLxqLz/xBkammeDAI6NSpqw/
`protect END_PROTECTED
