`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGfkp7ZVPKK/f0q3RJ9ab1CDzTSr/xNbrMprJ2Del8qpg8g9velO1sDBkI1nxVFr
4vwxSYFRMuoDtr3m7LOE0VD9WqBI5Kffx12Moq5orzyHKrkWGwzitgs/iHFOB8IX
IlIdsHtZgWsa4g7OgNfmoYWQwp0XKyJzAT+PVuJyRQXWWttXQwggYS5qZvrO8UD5
4ieBUHUIts9MLrXjhKjUS3mpIRkHW8K7oW8j8uwfo5f02OgQYT+aZWkP5j+AtmDf
sqX43z6cCHQ10GbXfJUEOLlb65KM/vR9jiSVY+68lJ7sZMR359iaJtjIZORaB2qE
B1Ah++zTgBsZxMWTwo75C5f8QwzqssfB/X3y6xiKX9u6Byx3h64IZdwZ3WQevIbC
QTh9+w/BzkOGD5S9mER0pt7GoBVFE6Tqgh71JtGLUx0=
`protect END_PROTECTED
