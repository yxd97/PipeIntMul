`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vf+8N9LCmn+k+JzFMDUXIzwY++Whz60CFBfQoLar0cXTGh42626WGhatFe+ZrqT2
kunYdTMW5OwqgwLF1kO0nq5BJCsChIYntzpBr5lCRKZ5aM7+8l07ESP/GUVe/c9X
/oy+ydGVp5q+unulmXY6u7Ppu9c8oqPYnsvhupsBMyhOXUkrF2DbfFUTRgNB3sPN
sjrF1K48Qb7a/oyddG+baKiJtulVkpTriPnRM/8RuuRtvM+nqVPyHNb7snwZUhWQ
nNymVnLVzMM1TNPKloxeN3B4O+bNjMr3InDdg3Xrw3b08NnQuHuCTg3J+XkfCGI6
rsntnnYh83m9RXtoss3CJACYoolHJ243Xh2G+ZgjKf8U4SFLD03P9hDAiZFgQn6K
rUaX2eLa2epKfAvTiUKHJ3zJDogc7e/Waz8lTjuFoAXXLDhdhTraSqsZHXRgYKCT
BYnCAKFe8d84HjFWMMGy/1oBYx2CYvcL5gCt6DlGCY8=
`protect END_PROTECTED
