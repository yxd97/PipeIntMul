`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5elXF3zjV8cWu7a+tg9DRx/xDgt2762ujWkr6KDPmrAlx3zGr3NNxFO0V/TLk7Kz
av31YsPN2DChv6MGd8Jc9vHqMXlw0l6ya6TYqhtBPXSSSZGZsSutr/IJMLS1QVeT
SIY3O9Oxaqxkie1CBSwo6ClWAVR0ortHeB9XrbUG3umx77tMQ0FZvRVS8sh862HU
Qz9t69L/EFhBnye4xpd+pgX8ObRIXL1kleM3BkXn/tYr/z4m+DFIdIo5PxHlse+b
YBsLslHYVFydfveJi11IWvGQ/0mRri5Q1tcpuJASbTvXg6VmOYrKJcBAuN6RCEdz
WxZ/Ahd99KnRu5tDTdeSinmio2dX1/L/2LRvhve3iDbounfkMskJeqAPj7n0Gdqw
Q036024DEWTMN0XMOnEggK+aHyxNFP7xxmGAmlKvivMyQR+Pd6vfskPTZvVcIUUa
pMVGXIxkwcyvymIvy/yxkptobTTb6TtUVFkWSzJlqPLTrrUiUmX6gk7epmAtmy1w
OCOLvO5d8Gq9GY1QaWuyn5WRpaVQWtPndpwjlTqX/dBw0S3lT1MZa0nnA4EhYzN+
qvS4S6Z3qu40asS9uA7SAWfy+hrzb2s14vkd4hzVlMuGtedsDumgkSGW+hqYWPY7
8CpxG30wL7pQIZtuVk9sIg+r38OEqiHZUxcO4hfHmF2Dn7jgYphsnwjc9tnN7Rac
Rk5qCWHsm0cpX47a1VBm7rtZyPKDZg3JVbjBg2kMlHvr6PaYuCK2w/Wvyse2VFmK
JxW/XH+/IzmdKkadFsPJBbH1KBpJAEEE395vQRP52krEhc1waI4bShDryFujo8dJ
0keiXs70x2+tW16NBkLoYHrvMvzgFepu93zTBo/v6lxldV3Jv8UZULM/fJkappDU
rUa5Xb+Ty1to2u1CR3Pw53UqzBq++8xSS2q36Z8kRqer9LAMpRhIMF7yV/C9hCxK
BaFf+XW3rhQHQeB649oIsOVYFElt5bdbdc2dPDXOA9cOBTDanE5Fs5qIZSlvw4sX
g6J4hiZ8CSoxm66FszVuiLLtZkgHXp24DnDMYIkPLBMA6UnN36VU9oFuoCvvsWWI
CnYT9L38mmGgo9fnEiY7Yow+o/tVkoQCVCb7Yd8nPHt+Dv0MHIhVMzFbvrYBMiw+
5D8K+ykh7JjLk2x0NgBpPg==
`protect END_PROTECTED
