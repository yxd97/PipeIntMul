`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6nsdkznlSmS4bNwYqTEPV8YDZUFLw4KNRQ8v86cac/E+VIyO8r7plA+AuniWgwBA
tXkqo421YScEEIbdza+YxWP5T8JZmN3gEx7ttH6UN+SQ4EJqWlRuUHOr00Ozhrhz
qVqvB5z1XBi2Z5ZSwAgzGnQpAL9Wz6ly3pDppekgY0tQv00MZ8n/eCO3M2khtN5S
UnkywhGt7x8i6oJ7BL5waizXNrJbWIwCXBSIV1SisebKEPLGCZ69qtOm2SOjnlhm
v6GPwnJsHxgXgBlpmoEhrLA9zIc1vG6inYhIcZ5GlmbHaYO6aqOJbuQ2WG6KEQUX
DFXAIwPvRh02nQ6BBCqaMyvkDiWagnnKDCvLZuJgx28IgU/knbSXykGQ61tBxljs
/xtfoAv6kZGPMBw8zK3eckV72impj5UnmZWE3zPU2/xfGs5RYO0QqYytk597RnIN
SnOYiTCdCHIwCVzFN5sKmWucn+3jr40INl03DrRfO58=
`protect END_PROTECTED
