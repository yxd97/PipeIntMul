`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DsIhBPfJ4r/COQz60wOyUN2ovzpol8kbqqXCGDOH7zDi6TlNKBx4UgiGQxVEK5Qt
stg1g46JY6G573xpsnd8DtlqMy4JwVrXAYHUN4hdllDJt17TZf/cwfMY0NjqMgCE
DyTctuOihT8Ae2ZW4vxhuMW5HDmYS6X2ZXuW8Mfkaw1yIvKqKEel4Ae5YSgSeu1U
C/TZpsZGc+J/oAOjHQU3lb7kXfvbAUz3aqMBKIXOVgJdQwmbIb/YqIpBp01GeKgM
waT7zyZBtJejATdOsTJ7NSkkNS5mpOKuUYmmqn27zOmJiZDExCvsyAxoUNK5HIAj
tzcg8CsKnE3yObvSwwbkcW4iMPrY63ELEq3shR1diIGV1o5SsIuWb3fZjBwfJsvS
RqSBvJfL8YZ8A/qH5Uxp6or7wbZXm1B3vVjEoYoZUxhm5dvxxPt2fbKSOmKi131W
Oh6dcrWA2jACG01/Cqi1bNUkgk9ovn4g7spPB7OHkPpkNwssTjOw0/Msp76x2E1V
G9533jeU0/vNHaWWR3Y2K1F74W/h9GLDXNmxKbDL6OGpNv60/67YznRdLiiCHYek
Cz0JadFCQFycuoZ9mL6b4g==
`protect END_PROTECTED
