`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TgNBUKcOI5mBySEVhyq1OMvTYQcIDQwj+kHvF8sUQdWl9bz1c830BBhI7E7dwhun
5trUe+uCylwe6ngS3SkUoPsYyzpA2heQ/aS2aOrJTrYKS6M4xz7dW5ULryYlJI+E
wUpt6IzRGKJrLfGlQPt8CRA7slRQyZSM5zoNPMn52WCsV6Zg6HNW9OlT8v9ba4Sd
A1lwPMl6kecQpZ2z0x1seSmnF1wEyLGcLBV82RMYjoplv6hj57psAGGThl5zkotb
4i4pXb4veg9DDBXokcGxScHefLDWLT2mVhA1xi+xGd4fsHjvwQCahgLcTASJ3kAp
V4+NeUGmnO03knXXtuYyctSlPF1U/cKnPMLo/u5b09wxMIjxCyugXwAFm+4ITiSM
Yo4U6+FkhMyeeR7n/gV28Q==
`protect END_PROTECTED
