`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KOnlDw2Szj7Hf1Gk695iPD+zMfn6qNsThX8j0E9INedYW1bGLEFAea1Dg6goSVMJ
ROja8hfCqTicuYmpUA6v1JCkW/FRFyr9un1dlT75ntyjuiDtEuVhfJQZft2YkDCy
0QZlPpqcI+qx9OqCV3mBQz8KqzC6P7aoDohQ0NBCzE5UCWAKC3pXpqaFi0luaUQf
H8/ig50T/scG0k0Ee7DrVoO7tUed/TUC77h52PeruxihasCsaTAqYt49a8NJQVsC
EDXiJMVo1ZdwLXL8WyVe/q7HNRbBE9pgTe9+sIDetzO5IZC5xQCnUlM62Jw1hwl9
mgmaf6vICyVBtLfOyD8H05lePdiDlrWJt0IDyiF3q3ZZxoOKvSW1dpTQS9y3G9bF
cQrjiEdsUy1Rg7E8xiDQ3oacWy9rCM2LlFhvmioRcmlEk/kM6sBnv/A/dVTYipgC
14z2y1XDuOzN+DE5d6X9gtbc+okRoPWwaPiH7IbecYgSlHuK2sc0s8mM2sb7vxAI
XbTgXWYI0fdI20NZocbWJA5pidQ2HIMTHuZjjQpbVuCOSlfZx8CxVUQuEcIP4jN1
5EDCbQUrUsckOkU0CAmt/9dTC49vYEx+w+gw8VSRicAIpX2gnUE14yG15KSsUNNm
NIjMkWahPHgUYZKZ7mFD8r2Bb2TssjF+6gGwvUcYrHtRYKPRBSpkvBqkTcJFJvoq
4XUdl3rARn/MwVwfqS/e89A61rUU8PZqblH1Fvy7Fz6nLlYage8tPORZ39mORUW7
v73avRbyqXUJM24310Yg9njCX3c05TuonhZU5cbjrINyP+qNFwZXDEx7L7+xxl3U
kpYxyYczM04hqpcxEPVrCC4rGB9eFuegYC58Fd8Ke4pMDoU5pLuttUwu3FuYGALR
bH76CRjt4fTRIYZa6x9WK9NuBpRYIj98wXg+B9MNbgXXU1/w2J1nX8xCdhCvWs7v
5UTEeXtV+nFlf6rDL5d3MkKLepKXeDS413fqb4VTw81KixdHu7WNwrONu9eTB4C9
1WhyL0QtKI66k7Orw/kKUotGu5XycujghERxff5LZLf3QwkT9H22eSxo5JfhV/l9
VTS5D2KPJmuEdK5dAgHgal/5sJEZ4mNMO3kgIaxWpnHZ+cWHvmkXlzo1qZgbW9o5
DJVi3PxHx9n2mr4xQ1relHdsE+Nt/wb9h2vIhSCiNqdTD0/67B35ZoISh5TcVVnD
`protect END_PROTECTED
