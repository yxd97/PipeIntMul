`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVY4pCNXbPCBE4HRFLcynhdTj/TOd4uOscDVr1t6dtmOOp0Ubo0wiUpYPzd5Q3oc
h/5Daw4w0KbsjCBXGtlM+MDzhmqFXkJUwKf1fT7h6UT0XQcinpBKcPa+mHTzmd8z
QECia3M5KlkxB5UeZ2CcuejhLcsCcDrQAjF7w11voMXvTSiZXX/xodZGCMI07K8I
Fr9H+mVefiKUsuxgMpvYQR6AZbhQcYQO8nw09zoPlZt+KThfp+7XZi1WNbFI33r3
a1JqGjau6RMYipkwMwqfrDn6gOohquGcgFrEW2Of24OUK97XAiDyfkNII7S6pTfz
3MypybEYZYtB6+NHEuB4hyLFwopn8+kQI7TSwuDz8jVNGcGIMbhrQT5dNDnHfAat
RdEe43jbpuiqYx9Lso//Eg==
`protect END_PROTECTED
