`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5lqbvPJd5kbEgEvId890xEJBF3eofeh9rbbxn40pd0+Q1Ng0dujMvWXbtwJ7DuU
CMd7Vv+M+0qty5NIKeeoTBhKS1Rih+BDKSAqH/N0YdiZncBKLEhOxWB8ZjABYiIQ
jxEJID4vc6bhTqQvU7gXxbOw2QytgkzrO1aJ5uSz7fl1XvZ6yz1XfFqgr7jgsn1g
rST7GrQbMH4YGMWgU0LR11dy0GFsoGgh4Kad4xcExKucXBjYG66WTx5st84jd5SA
NxU004vqg8L+r3z5SPY56quq5rCkD123fh4O/UrH94BUCy0eVMBBsmwCgXnUjbG6
KTVz1VLlZcQqBG3si85DZmiLEH+B80/HSzLLR2xlyV1+cuCBD6nT5cs85bgCosJ+
DQUoPcC5wsGKOlSQHLZW8T/WhwtsItRRBrA8dl+JNUp1hcOhiX31f/TN3HKqVGkw
ijDuyI8qYDGPpbWVGL3n3h0f5dunYBVf9l9A1v+gCTJjsx/b2UhQH3I8yHxQiU+R
Flmq/PGCfSTrF8XjyMqn2WC1jL+IlVvQZMdiM7YMimufwtrB8icm96vVl0YcECf9
gF+1wqnkr3me0P23ssEH/oLdgRbEm0f7PkScBsfVgRu4woJmnCYNz0okF59tKYlX
rQtyAadmuygtBajoTp8xrA==
`protect END_PROTECTED
