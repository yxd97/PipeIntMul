`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8w1REXrj2hZZEgdHHDqbc+3ruHpiCEk1jYrJHkfpZCddCCU7rPaDYY3EczyZTwTr
YFsOiu9n83dSaJ00yqY+InceTzSD0nL4zL+gI2S7/v5lr2KmgGlpbSfR8P8SSoA8
Pgu+Zisbd2sRqb14+nfOsMgn2WfGlyH/U62iSx/3QFomP4on75fwG+xiCBMw4YN1
WE5M8PJSdnRFmbCs8YQJC23/zRD9PHxlAliKoiWhtd1eqTfjGMfafdz2wA/37Nnc
hGZhAusAmlZMUPYzoCSkbsspnnCeUpgkpiLqnU/fub+dc5UAsDmWSgPRDjQ29AAc
UKxiy9dNS5330QJZnPb3qnKm+bEVZZ0hPsKD+E+Xm1rdvPEdOFHMWwH4c1ZdtNE4
ONGhyoqPkNH1S8X4ehvWD+phbVylUmgJgobmBBNyiHhJnFXV1sqhiNqZaqUTszwG
mJ6lAX2SvTeO2FkCUly5WD2cFZeXBQaRK6jsCKP+sAHAuIZw/NLr+j5uhjowl2ZG
i5OZbIvzq2gS6RQJ3ewrqhBbsMclkAlLkuUGhLBt02OOJ5rBcmcVxPmnSJWFYGbE
SecV01wtzc5Kb0x6l42mqI495zWm/YuLzFJvgc1xaEhRdd7QhVgdIjGtPIkwStqH
Yf7Z8ZQQNdkO8TxU+WdbPLi4HS3/4HnTP8L91mrAhXI=
`protect END_PROTECTED
