`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mEyhCAfVvxqbMJ9+GF1mJZGYHpqeH7Ngh35VxdHIEPIrIS6p6n2kZAlZ6TVNHvoR
28gdfsPKqhoR3+iajny0pIb2242WWFLeXYhuEMGMik1bkXSoUrflXPSTkL8tprq4
MNMj+4TAjKNcJdbJCCE+Ke9Ic91ZSQiod8A0xEIsq+lEeiXDFEc+JytktTC4O1rr
VxJYKwrHTj7yI0pQvfVu4w==
`protect END_PROTECTED
