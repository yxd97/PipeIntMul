`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OC1x+iLp28Km+JFuH1lDS33I9i4jhdDEASy6BtipLiMEGZ4ZEChGW/x6R/+sH1ta
iwYU4LFKBA7wZ6gvJ9nNBx8KMi1gt31NpNPy0ImvH7Chy8bWGgduledR53ZAZmk9
KGhybk7eMzZmKBn/FWbHAt8sYwzgWGIjfKgc8Yrte35NBZq6Zvr01RbG8KiYt2cf
itaBHBn2Cjr5PCEkXUxjzG0UtvSESKrV1rPtT7xEDaaR8DhaSaMall0GxytLg93t
j3jziNhjv8LcYKy/GtOtCaklDfFzYVcQrE69BhI2XBJmtFPfQB6zZOxD6HPt/Quy
jQ+oJLRPFOSvXgTw9JRHYA==
`protect END_PROTECTED
