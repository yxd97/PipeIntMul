`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJ2CK9WFnWZydREMrjJBQAkjRojUb7pLDfjN1plHefDtnM4SDcaGx09YeNmITTfY
HOsWL8reYSoUJdIGankFXQZpZyEoErnpxymYaVnXtUSFNRMJBksAD6DDJDngPkhX
7W9m5Qlhr4psltVzQFFwmBCYgwj70woYbp/tBqPDK1YMEvxmHMxZ95hrYY+PbW3h
na8g7/IGbCorTqcUpQFB08DuCyV4dmcAywvQuPOvkXqb6u6TgGfMtfmP3OUWFWNt
a6SudZBiJEyx3OksFGK5NZ7t1vOK6GDPaTlrf8TY4MFoWyXd8srIk91NbBOCvdXo
aBXyJbWQX9Ng175ejhfLPcrkziFUCvGyJ9I6bIcB/0ODxHIH7HjW3UNa/TYgsggI
kLGsWPmQxUDtrtV9tttpvAXMvaX1kaAj7rs1U86vqe8=
`protect END_PROTECTED
