`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XajnrJ8PHWgR77FPW2ISRibAX0+iYpZR+si7OR4Yif557gjHK86ACcjuVMMEGHQ
iJmN9NG7AbHFjGfPDwxaxCEdXWvlcB2uPAF0rT7MHeqQ5yiGbD9UpxlVIMP4iqb9
h4PJiHueM9Dy1aM4lXTa/Lj9wxQ/8vpOGVyBs5no93UEIzAzAaRKLaS2FnbKWfKd
63fSHXK8mTRZBoLy832Ivj283aEM72nxxR0pdoUss3vX6ysgG2H2WvRHvdyP8hUh
76jteA17aRaHRvqae8pLMn8GqJd7vuFzsQrml2HnSV4QKbdVLkrqFt7D0gRFZyLu
D1HoXl0B2e/qKy5K/cbvhZZy06/4yzuJZLGzh8IO1w+XkKR9XhCbb7SQj0130q7y
oWHruerrwfOT1ZlZiEX/1U8BsRH8iLkvxfTZrCIx00xMfWOiuas5EsYrpPlLfs2G
F7bxxYMJVFQy6pRRv6vyNeeXjny0RlLZcIvnoE6B0hQ=
`protect END_PROTECTED
