`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZFTaqaiP1ZkOibye6M0N3Tt2NqCe2siIHa5hD3gBaYrYzF4CSjfr2enSArOKXHLS
oU53V3DUjBsWR8j9cb9mlJI7mYYxwzUDHe2hp1OZTdvRIvHnQvf1xdn/CrEPfYop
YUGHLsbuRBUjtP3y5DplseKeJKLq5A6+R5HRbQGC3/GdzELfTtZGFRwtidVK+V4h
xHt2y/bs+ZJMHC4LlAL7nSgmUWEgRBsRrLrEDHaoGglb90HIohy/QcqjSJm735Dm
fUi3rhh39/TPvrpUdpyysiKTv3kLiIMRpFtlFbaEbPRfFV+Tkqy+/o0ja0RdV1Vs
vn8E9qL4ROEH+6NTreCUgrPe/vkekFAVXnp+nEbRri7FHB6whUE++focvhAnRtgh
avv9nIK1Vq7n+9KgBqml2F+YEV+1DA27HYOxeAdozGCxZ5CU6oMbcfyuur/RPDZ1
LLhWZWnyNOrGLXWx2HZWK0Ch66yOEQMtZmKyX1G0NwbV7WupgFSO2PdVy/pa80+O
pTq3ObPiEpl3Hwr0Ql9xzB6XjTLaHDZPC3YSsoNADlS6f0a9VnzHvQsK1jiU/z2s
D2P6Rl7t36kg3+a92pNLOid3NKbri4OkozEjYYQOUF3iZ8X5ldoiKGWY/O6ExAAN
vEg8913MpveJQTQQa1cBxkMSzp4pcyoUL4wrAl8Lu/I+NNE4u1NYEBaG293GX8KQ
SbFaCggNPBIs253Nm9kNWh7kDct+aYWiuS2/Tn9/2qPfMTloS18x4TCaDG8XhH6w
EXzqZQMkyCcAnDuGqP4Aig==
`protect END_PROTECTED
