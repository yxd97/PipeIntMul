`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vXSTASZfZcmWtS9ONJt6JBHsJKRO99hazeitSwc9Z5fowk0pXqNFrM6l7EHGrDIa
uAIqV7CwUrlHd2HzQ6MlKwIGh90Wkiee0Y28Fv8SNnUSrqwHrOup5UpAHM1bf0BL
JNzg4QSgFsC9c4U9Jc8RQnKgjaBujCrH9/kwwc8xBfn/lV06AjnMXXOGgGKvRpUj
j+josJ4VMisw2Rq/OxMu339ZyAD4ePvBjG+I0kqqkHoh49Md2EkWDXd4n9IaXGHl
5sqXOFgoIDzkLm4WSfTtsYjwzvTV9ykEqROpehDQgb80I7RNqVTqX27WjvpWTfyQ
km2jR0BNyF4Rj3MZCM2DOfe0d5oZJTXMFgvlcojr8hRh9x3wwsqdhDjtQ4yGf7yp
m22rZgl2ml8QwwZN8ARNb0y2AuLaiu3eH9IW2hyDAtwNfn6RgMFXIgkx2WPkbebn
zv2ggFq5xeIDBLCImyd+/wysmL17JAZ78FI3FIfwPj8=
`protect END_PROTECTED
