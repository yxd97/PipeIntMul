`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FEoOGkerkP8IkCDUutm9AXMV3KyraTfbuaz1N0fty1p6rcCkQHerlTABzLOhfixr
F8Ht5dqU84xXSbEb2sgwRgj3FWH45IdITcCH1vNgTAJ0/KSltGTvvoUFYbgGfRz1
jn8uxMlItiTHwpn5Lc2I7hX8bh8VuDbthHHAUvLbz1Gb8Uf50yAUTQBvx3DyPOfl
B1pAVOge+0imi9xwBuxRPJpFrvsalFIpwpWdWXsbGfI5/Shhf1uVf8i1M9exEJZ1
xHXJGakWAUxHu9i1X1uIMBKaGXHqOyVWDoTU3dYCd7k=
`protect END_PROTECTED
