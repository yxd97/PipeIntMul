`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YlJmcxxlSIclaMW5nyc22UysTSpZOuA2xtJkawJlT5wmUn84PqMNpOJRlXndtNp
yC5vZ9viJ/wOlLRc1HS5zYJMAgSW9YtxTI+ciLD0fLkQcJiuVeG+MOER/0BrSM7a
948hb4fy7HDHH08s9SPiiFOE0+Z/9iN0LQ5YueKh/p5lq35taAE/Hwx63EaqBCWR
I97VQGj2yySJEXcturYIhS0SVsjk+3G6SYu7Rbse3qbj7QemZs9iG73BjXteuTnH
XzLxHenqPWdNJAra2d0Poo9gWbEiAmEu5K7gzwApdnfotopZZbGljf80fCPap22v
lUJOwtk99XhbKRfJQjvpwNICUd4UbOR0SVrQs4O9SvhHeGmd4SPOEu92qVaHaZVN
4qzfrm9NlxuCvuMCESecGu4kvJIuIRxnXEW6SkJGaqGx9YZa9f7lgNZcuNyt21sJ
S7zEAfHKtY2/48TbsEBJMIV+LWZXXzZqUPwd3b9o/w0eJ0lcWX4Ljk58e8nxy7hP
eCIYV4NgpYDsXSmhE21FBLG7lTSPaY4+2uVS8xR/rYRc/KCEVhzpmWCCfHqlbsQ2
+CqsiH1sS4aB7WDiEePg2nQcXbIbVP4v2+EGRTkrIXgpIV+rzgum3va8YRmrqbwG
3bA46VJAqIqL467GvXSPlQNNBmZQnPRq821lSXgV3lLpWFnHimrFhfgUXGy/j/kh
VA4cLFdp+R7QNS7QtDrvNe7yl4dfiKIKU7eWiQz2w6ZR8YTcWq0o4We0EODWU1ii
m/6dGS4VrZCpzQXB0HCU3Xr+sj0kz+SB0jnrX08YAwsxFN9t4b4zwuMxeJCWdK5l
ei8Odp0C+dwiOEpD4xxknBnS87ljuWOiHwz6sp8ZW8t1L3M+ZlP2LSm84b4TggNh
Rkn7kQ9SKFcdVlTsjharSMSZCH9JCyy5/zd1CyBtzrWJT3Mvr6cbwYil5AgVEZzC
hlqtnMA0/dkHvpNpJuC5UBYDglHFuTpsqyvTVtDBm3vaHRHKGro6HrbryfiIvfTI
hgNcohXXgEPmqY4Uyo6WSdFz6xbMgzKOyGZlMFwvge3uAgvftC8ueYBXh8TfMnDK
jKl0j5t/UfxVd7XeDYKvOK6K8MAWPtCTj6E0g3kRD8Ph29e+AD5Sf2WUw+kkiBlH
wrTrJ353jKSQa9aUjIhz2otcSGlIkz90ZUC8S3JQD4vblTkhgEqEJkamHl3l1qCJ
yylnj5IYfQ/yzDPHls76oyQ24qhVi93YhLTp+oMlQbGAG+d0P1Yusc7KEb9AoAr4
YKetiy6O291A9UrfVye5dbSuVQNc8m46NGkncsBLjo+VlWyFRUVhew+z0DFnoPqS
5O8lkQj5eyma4tBvXWBD+buQBBHV6tfSgp30cVojt1U3K5LjTXV/lOYeOXn6oyHs
GYQMO/mTn8OsDSVu5TtEQgM8agRf2vtTh8XG+TXr6oZcIbULuYNGau/fiuIRXaEe
`protect END_PROTECTED
