`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28TzDsqLVfbZq0zAGg3ArOFce+ytPhXRvgfnxwn4+R9cv09Bjk+ZKRPTQDZ9j056
Dw2mAHNgDwafKVMRQcXn5/TYNsBB7xdoyz1dL9HWT1KH3CBBnQpBM1lcNM+G5BSO
gBuJ8ZNRmuXlgm2knIwwr1Fi2Xai6abU5HPWRSeN/ozMAs9U1UAqtAkHvK93b0De
wrU9wDvcctID8ZPZx5VHHj+UcJuBllLiHw/vsp33AaZNP7ibzM6jLFNgqlvoJxxs
nzGjRdl8b9Qe1V0RGSGKkVtP58+FWkb6kLRioAX/hBl0yIf0Gsax8QIoyGFnpis3
DrWQsVTjpR1V5fUQ0UiKi1P4XNJdRu4Jv1ZCl8wVpWdyn4z4sQNGKjgfHa9fLH0H
WAi9if0cswL8FMdFvN+xcE3EZ8JnQxWqwWohFX0TKbrFfvZmwoFzz9rpjwzD0PnT
1Fi5tHVAe595yHvGU+M5SpKTlkIl3S62jLFwXQE+SbVjKxj2Cv4cqJc5/liL6de2
y/qgriyIRDPXnMsJKZNO6KGFKtsT1MLjGcdT85jFr/cAZrlsFr9/SVP0TJ858ZKZ
Y5uctXsD+ykCnM9g5pE+YXRcytbfe1FnW8e8DmpqZQWjUeT+h+Nbvg8HOeAmhctU
Y32CkS9KVyc2LL/+J8T5afJ3jlrr60kK9ozt7Q+yTXV6QTz4922sHacVyxZ5egRJ
7azhzwMnbUm30hl7slUhdf8Lk5d0ZYx+dxgLv8nxEQI=
`protect END_PROTECTED
