`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YYH6PTsL5ytK4r+v6nWfPW5CjE8MUwiRMUMVJUHdmso6ojB2HvMgdwTQ1cbWltZ5
E5U+vnVfTThE1AkvZt3CcDh204CbWAqL75FTbc1tc2BqT5+Av2iYzeismcV3284u
nKYT3WPly3mF4VgBj/FCUs+/+yzTdzzQlczwEEzRmu8PBTPHwTm50bKhH599oa0W
sbzuNuC+6Q46bn4FWEBm4nIN09M8PD0Lg+gBSkxqPuL8ggy+Kb/3CAZ1yoKbEdcI
Wku/czOFt3ZS7EPgIMAk0SAnuXnMX9chfo3C+Ce0ZkSJuG7nRA0TVnrJLACkNZX3
v6xctX53WrhWgpyGVv8TjzUqSKNb8jaMcO/v7jpn7X/J4ATcTcv3ea4EtxHGNPoi
Ypd2zQKSWBh2z04JP9x4438V+GkszzaWK0hb6FeKL0mR/xpdyC7DpMkgnVO94Hnm
G01Auyda9SHBoWzMclq8Tixk5ocTJW5R9k/AQ45k9h8=
`protect END_PROTECTED
