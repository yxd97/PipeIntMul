`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6eRBcgIaehZL+ZSw+0BIVsA93F4HI+kKLOsOLJ05w4efobs+x2S+pnadqv8fKSNW
mf8YkF262sxwS0oXlaYz4730c1n9hjgKw4GgGdsnOJ7JQM9/bjSyFFdAqhIoVyiX
13cgAEzR3S6/xEHkUd4VkTetLSS8H4aFe7yX+zkTg5YcwDbEaBJ8jwzerJqewVIe
cU9LH81Q4mWRzqWT4pWwQ5LHnb3xGZH3VreSCb6EYsWwyAUvdnfcY92LcQr70UXG
RHvyIF26LW5Iz8n/Tb2wtGZxCSEXukN8XDjomNZ8KIA40+RgfLivwEp/m7ee7L9q
zxx1+0smiuP1nqIQ7fPqVyh097D5Fiye1suQtxeDHMNNS4yiUQOgGUc3U8wK95Gj
qF2vupnEeyl1SMKwKD/GOPjDKyuwsjrU3ikc/JYT+oEuupLN9CQX9SwxCrWPDMdW
zr7odq9VHRCG67JtEwZQ2PtCnWj5wwXCnJkRYeANhDDycbDlYL+ECEyGxSZLJAQb
DVErvINvHh4JQ+7BZ1TJ+F3gA07jIc3aiW7RkCRYgeUr5Q78dPRd13xc8aSjcr5N
qQM8CnMJnURU2xkWSdx2WeisEjPj4qL8aplviBjLShzo3Fc1m0XJ7mxewTHx1pp9
PeKU8mTcED4HfjnPC2zCZw==
`protect END_PROTECTED
