`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jfoIxyKsVSnMXq5zEm8JzaTjlAKEEkuycznIeertenI2ttbw30+DtxuDw5OZbm3+
uUg58Q3ES0iyH5eVy7AxMm/pRj9CBOpyl1EBWY2ffCYmhv6l3HJ6h0wGISRu5XHl
UCZyFfZS0GqJLfRtQw0ILjFTW5IIq9MWSZk2tG3eG4gUMCuEwXsLrM8/UuRNhwBL
mV7L2QcbhD6/LonViDNoJ1kF0GbkF9umqfbY35+dHoMCxqYpEy0NoRORHy7NRz6k
quIBq2npMklPLHdsbaq6mOqQn53Eze70bWdxGU+FYGG4ZkIHLGwf5QJKxpjpjVVy
ODpl17dcf5nxlvXT+HHopSdE7Eh9CT9tQcwUmKyjN84dIhwXjsA8s6QCqfqzacam
kY5EOA3O8/Sa7z7RsMjL4n3NvuUIJfi4e5UuEoq7OJwkHqJSBbbqw0vCQVlg4P56
Tw1su/+FVmpc5qL+TgYVs0pNiPhh4XJBnhJ5NvNA0d0=
`protect END_PROTECTED
