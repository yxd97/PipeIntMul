`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nh79aX3nSkluEwZeiSi4ZKA0T1b6GlBMI60UUEsVPSIDE+RfJKCluCUESgn0/P9o
j87jFPQXo3Srf7cQRc5wOZv814ya+gWmjYi3DhscNNGyCsWpr6pRzghiIbZSwXD8
GDMe4CEdGXBAsxSZhZL53Un2750ICxCMdI0A6y8K+Pyz5ZQZJlJ4kmhuuNcawh+t
ZCqyI85+Pq+elJl2clELB63RmfQckpnyj0g9q4qrJ1eY01Dr254iTt2H/wEEaM8Z
ekwnTSQPrjmExROTztuZoj4MHQ7RsIX6isngbb4DNvHvTdiwwmVXVFF9Ff2FE+O0
1XJn1d3qv/sdWvxOIRhFUIGXibz36FNIIdCxwcEK8KulAd+sH6WfBNSJuZdTQ3se
YYv1Umc43OIIEJfyCpQjnuXbPBMm6M5i/ue+dsBUrQDX6Jo3UWgJTeAMNPJB3Scc
0U0Fn32De4EgUyBv7496SffA1e6Rp72RfVsjYn22CpAM6ZngadfNc+oSN8Jmxrql
6LDTj4mo5hm0cSZsXkTcwa+TYiqhh9+ykVcLFSnLNKLQ6n2CN0F3kOGL70DsfwrG
AZbbTd/A+L2F2Z8qnJldbaENA0jm+rLsTQZIBklSTmqF1d6f7sbw1UZiu+tovBZH
ap8jWd8qPLvqISjhTS8SrIW1jskU7EMIan7Ix+Vxar1gF3v6xpKGvc9EtzpTJcl4
`protect END_PROTECTED
