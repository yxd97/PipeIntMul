`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Auq7HJBRUGXcLf4vvV8qMkTx4fZgQi1w2ePWXVFI4vcKp0oMzfVZlXSMYqQxX7o
NBNZ0pXePV8oEbs8zk0JMhPhMjP4Js1DX5pHkCaRcsJzGvXEJ2QvBg4ctQDHq7KK
dJElQfpZ5txiYuuJGDlMSgKix97nCNxqqfsnnehULVIgw2U/TIHBk9pLsgXwwhQG
pEI6VQh5iLQeElExdXsSXy7AxDZan52gkXJmnRxa9yVVWmJyqo0Ia8mTK54Te39N
Sjg4/rVvrfAj/Gexilo7xCKOQCEhWp02oIIDVCzd8AN/ktjPrEWrqgq9vfX+we8q
r+ez+s0W0x2gOfmkeGgilw==
`protect END_PROTECTED
