`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubi1n4+fxgb7h1BDyVGGUV4tsAG9mSAfcULIxCGWpCRdIdK9XtSQ90FgQQ4gnY9i
9S5hWkTwLL3BVI67arzgy3Egq4USxt2CSnj0FEvryWnr71+RUvnTnKhHWsKMhrJg
vUH+O8MwnHJPY8JmW5MExKP3AdE4crZECSuUmsZNEwvGujAYCG78fWO0eytocJJP
HprwTlQPor7BjdGQ2+X1ydtH9uXb2FXFAvBs6atUbQrtQwq5LvAnsWZfy5r+JfKl
9kUERdLrO0Thdz506C1ZRlan1yO43SEG2JgVAK871LXA9Fs1xn4312qth0LSptkF
7kNIyAUGpek1h1QC/8Jt5g==
`protect END_PROTECTED
