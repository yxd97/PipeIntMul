`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mlah2bkpo+98jFx5hmyHEm8PAV0JhU8gslJNhgcvKhbCGtYNlLs7DadV42o57IK7
HHw+T4WFNBiChmUjJPKQE48Jb/6YhkJFVCRpfJHEXlurl82E1Vq5uMr4o1ixsVIN
mpTUZ2Pb43XGzKK2bSJv8OncToHMt3BcgMIioSBWLH7HSHfRJUVuTb9iYDPJpTCg
n/L6DGLigB0C+jVLD0BaW6YPO/5ROB98/L8xxun3/JAuPRYJIk6YQSemp/lQW6Vw
5avLj6876RUXI9lPTWkYRdWveErb7HLlqML5jCdzuBJhI+jkYfMqfbl1TJqX8HBs
G1Eu+9aQFImSSjg2qarAYiD/TBrplUumwAtc7uIBWlfbTjPandTnmgUPHaE93NvK
gBkKMJQ3RG16gpYKcPho+LvQ28pa6pb27tTF/ahc/Xn+VFbDvYPkubX9N8sepX72
W9fkQS0psLgKHC9NjrpkPSkEKSQH3BU1tabSVPLF6BCYAM8pdlvyrRtU8qIHhd0D
DjfnlDMfENadgBVsm+OCjtvnYX5H7H3D69l8ggoX8GdJL5+jDmXou7NPzYGlZxpv
/8c7KsmIUdHvuIJ0ttQaHJ7YPhi8rBLBxDPBfKz2w8o2Mk3YvNuTJ0Pw7pVDlX/r
TfRjk4S6IQItuJ8X4QHXDzXbd8CdgzjmbxU5EC24htPWQ3sz3aHDzlzi4Q1qS0dD
JOfpSuuRpNKpeIneXwQFtkLciB0HTFyp/YO/5z5h9S2+v1pT8A4FbFQD3l2b09bZ
fIp+8oXtWxAJg0w2y4/iL3bBOcI8+hb1cTIEEmkEfg/W/FQU/Ub/nqFvDDhmdEut
ZCjK6CegeQYvOxxNEx5hmvpFn4cuswX8P6AOzp0EAqQR6Curw2vMvg8NRiWETEb7
GcfraB7FG4EFD8VU/qjL66s/pyRVMpB8pg9XEdQDNYyAmLhEzRg/uYFKzohfx6iM
2VJOiwhBs5/Jq1xMsyx6WSKYAQhwdZmmw6AREdJa2hgkTaeAJJ1o6dJYNs5W/XQA
FQOB6XODQWFdJEeGnW1kwMMDLoqccFIjxrM6KgIntOxGphi107Veft39KrrhV1rI
SMisIaUjI0Pzz3GqICzET3pFeI5N4FcNYHEk4qIqJT+ZwlO5+MdX+jFbK1AEMOF4
`protect END_PROTECTED
