`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GYxiXQhw+93XJCdrJXnnt4uGRagqOxq6OT4kMihLw4sFDp/HApD2zFWXVIlhitib
yiWAp16bmCd1Xt/nvTpYzyg5dBvogFWYzxwDD5+dno189Kj55qmb4n8VH2o7cF1I
RIw8fb0OwD/u9iQtZMsl+Q/+LptxbEDRbe+DE6ZoAIhqXGYWU/fSKgpewC3M9qzP
s0Cw/9mfnbzGdKo7riIQgFQahEIn8Fbyq/V8dmM6nZ/dUsj3CuwjZqr2urmbMYGy
1TMt3d2xi1v9H+I78daibUSmtH4X/jmrKH/Mn64gcYCuAtnWp5hSLSoajewi4QUi
+FAXpbtdQDwCLCoAmUBuQV+UL6XKbtm5jsIMC/34av81oQjx+FuEnIi5YMTnbyfn
`protect END_PROTECTED
