`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7iyD8FjWxe8UWcem2LQvmfu15x1dQKwVRdwuqaXKmDclJIqjCVIOB6Obv7uFkcq2
dMSVcbXeVHfttXq85fS75pwfiHDfwmx5qmmpd3GQ12rr5Bm+jwgvIk0Q9DlrwAn5
+IE3COyFnJ0WCZ3QUdJ5ql+6R6bFqcksbi/j+9LRFKNnbYfVcHuCXsKYrFK4Sbsm
q1mTxvTHl8MDyw1PS5zLHp7AzM6Be1cWpDLoL0oyxRRlFw085jdrrVuOX00PXArh
nyD6R45qd0ZbiogM8AA/VNFN5N/7NSHBmVw9AVSyIOybwh+BmS4w7sYz9owzondA
k8OraWdjtAmQh2FijlnjERewghTBvHmxoaYmakqib1ps3lI8MlxeTkDUNRqquk+Z
vvZ9QsAhhFFqfxsv+o+AsnBMqBB79p9RBg6b3mS9H1iNFQPW0mpxTohxukpf+/TT
nrIj4ekXKdvpQnvsO63WjP+5KfQOVO3WxmX4fJteQT5XU6StsQTIuexZWPq1i11g
Wq7oui9Cr0IpXpRqTDPCbwy8QJnD2D7AvthezIGUrVSekcL7OCKUD9DOMbzFJaON
yteVNPrryISPP/RgCE5lb826neWe/sQG/DNMwVB/qNZyfzj6dCUL0zTBi2KPTQYb
5TJ7ITNVr+SdJYM4lE1b4uFDOlxGU3UHOagiWFE7g9IY2wlk6NPtP/r1oxDpRhXu
3MQtJJuRDdErgf/JLXKFnjU5IdE3igtrGlnfudJLe2yhAJjkcYuuWkJ5v8DWAX4m
wUImV0KCtVmSeP2Dd4HBWs06I/VacrBToMlSKttuIjAdoAxtYVhb3E6AD6WJ/dhy
Nxtjf8BKgeGu6D3BVkSqLbh3sD9ZflX2rK7PVuGCiXiBof2yOLtgfNgEi63YTJdt
3jbqjQeSEVWdPn/q2f/ObsE3BzANn/7/ClyQZ9iSroZGxyHC0i84pb5pp7XNVdiU
k28pLDpkx4cLiyQ+7O+OUOqCeLnb1Owe/YbVHhMJZkOF1lMtAz3LKeJu/6kLs4Fc
XVEX7GW2N48FafY2IxsYhhWfyd2npUMmA+dYXGBcvJjU9d+wru6VMln0oy2+SFQB
cDh23+YpDEUMqZQxzeWGj9Gv3UYwvaPx6FBiG34eZ99rHiaXvgSE9yEl7TX0WdZd
KiBFec30cOy/C6fouTSUl+VxCs9c/cXQe/hW+cLyJfKkDeaFTD1PD0pe3v6jD407
gk1FB5rpEZwNNzpZOfLfhruAds3nAvOd4T05i3JyjprYRg2mg/VyPkn6sZ/5Cnx7
6QAcwAUlRtPVJMkXIyTZgbuLtpkt61YJ7lFZMIUnBwlYOG/iT8saV6xccftydFBz
YdQOklSRR3Dtik+Y80FAdD2wAeuG7IoLwyXLQUzTbPVYwTGviD7gzpbTHs7y4Ztm
milEXrwO0UiKhZugdUKCTPT3OdqspR4xSL2FIirt+QJJmRvLjYKzTOiUjVbqndHF
qReMePxAIC+xFfh+sHMH2fUqxJeYLWOo+8R9h/R8g3Dzf2Xb+0Vyd4l9jxZrlMyG
NoaPiaPE1rogUCMTISeEITjZoeMztJqfE6FhtgAlbEsQTk5dunCLtZjNpo1SMFcB
DyAujwREqCQjWqsXat8U7UF2YRmZcWxLppWxeXpJCH/2VfekzOQ4x/BRcyiGJBwN
MYGCa/YFi8N+bvnl8o4A8hs6MmkRq3ZhzbgdYdV/attdFiMlucfanwIOfspdqQfu
aTHuXHBTeKUEDudRlacvINKLnKyqR/tjWT4Db1ddr8819n2j/ueS7Ksn9IhmGpKa
Ds6iDCorvBU4iOKemLaRYodTw2oUD74dGmTCq4jiwGb88T57XSjS4Mqbk74DjgtZ
fxmVXoatKc+ZT/jXr368fsNQeWR3lF+b++gnacdefmT9eBY5FRLqRHlsw0AMxg9s
k5i2w/EmjI++JTdGaRrCCQLF0Hzo//XM9Ei5D9sctmUvLqG8CoGybslDDy7N94yq
Ho2e/5g4hvoXNcjnYAsTx/37Nzi/DXe8i59LQ7Gb9OiU8/cs9QRBZZtBTxk4xcPj
vaumT9+mIrHCzBJuVjQ7YPcasmpgFX2EbbrH0SD+7zt+sVFLPq39yUBrN44qL43I
v76bLe+OcpMm4g4+clR59XmMjgEyjwl5pi6W/Y+/eoLNsBQmoYmPbYvSaGYhifdm
MwGLoHQDmTCeY6TrXVyINzu5vhrlW6tM71M58tHapVmJ8iyj4XDT+8pDrW1X0F/F
3rOqxelyPUyPJOwMn+qHduPxDKrDxZ7MTUi1iYP0JeNd6p7ZtNvxUI6weVNJNecB
E8URQiRRLKcrsx5N2gVZT1VF5zhgRyc0xRrXHWSB2VkSJX/i2Et90IwcSQVQyMDb
igjxofA+MvItgvDHYat5AmUFf2K2YFcvK/yacTdOig1NJRg+bP85jTLJnfyX8aJH
hzbnJoRabRNDjzjsNQYpK+/DV60nlIspd9wan67PquEAsYuJkShHccCu3rO/tH4h
wxgO4ePef0J9PkIOAz13Pkjrt7a7nPxVsVA/Yf4V0LAXcYT8dYzqGzDslGXA5rJG
wUfWqaEOWIxnlKjoN8km38wdxx4W97AX8CtxD4wxZ7Kbxbyw6PwwOBmjRX3UWGuB
y9fA83Zb1weLr9g22rHAZq5ETUMwsHyHgTQiMShyRusa6DXa0+Xpec/QOAZ1R5AS
K2dQXdI2Bp8OXVVibaifJM6sbERkMbvBihqYaIecqJu7lVlcMfikTXMCTMif7H9q
s1pRjMnapmHfqPK0RmdzaU7WTFJ+xKn+WLRMM6hxqTrE1/nveJsHAEjWtIO1jaJN
e8zvvh7gCJ+Gwjj5q6qHffuoluYwYV2v08J1TnR7bQE42IGZRfdeLG+YGVijSkHY
pvzUOHvKAtERVxnI4pSRBoZuSMNRBRmquOUqREytJGsIIrVVdNquc408QUwxcj3D
RRWoS2+w0fnGPnX6A0BwrbzGXLX0VhCkjUWkAziVkr6zfhYBJdTstfDliMH0aRj2
7anK9RLiAj8kjOGwcQX9n0j1X1c/T4PybM6qsmhaTObhwo+bboyCk62Eidwh1Bsi
dsyqjzJYEMCYIxJ6h8b6KXf1OiV4Q3Cqxna60o01TZKFMOyliFO5K1LSZRIDLEd9
eiWwUtBs0Jrc6KUfePZz6Ky9OZKlzGyNs1CurKii7xGzSttOES4ie0c6lZDI1SOE
quttX9kRQzHz7oAIks/14juOShGTLdZmFCVoncR9aH+dKLy0GBUZoQCRJRDbcz/E
U6rQZyz1jU+wCR6vKEMnJv7pLsXbBrgRyEF/a58hUAMUNi2jviGhyui9YqsUU3lK
KwC3u2R25ojL4tcgItZnPtlubbbbuduigoWCvsHBSpaI++5G5R3Wmm8kwzpodJYu
ag+u6a7gbiRz4pEng1LTGy/laecsVFGDs2yJ5x8n2iPaTTySISaA77OfVilqvvw5
wIQ/ZmqPD2J+gl212gdz1L6d4bwmLj+CbKtxJyxw3pLPbgg/N4LDsVyIZUpFEuk/
/H/BfvCzjhviVv8ffw6O68P0qzp230aGYRAw93AVnBAxycJFl1aAxwvIQKVJ+97O
iaKjOa6AoCR++pf/aOY3Bg2O68eJzMlYvIBv1afC1L6Vfy5jt6h6BDK7Gu9+qkDG
3o1Objn/Apm9AF3Ktzk8SVSZtRx4bYvqvBGgLwRxVkN/L1a3wy+f2rCEJkPMsNuB
0MYnD+gvDYqTOxc9JXbYH1DyaK4sLUYFsGomQ15+We/cqV/rsRNpybQCiFHLajs2
slhfXZd02d+SW4Zv800aEbPyFgaDoVK0XALgUMm+ToeSx1gk3kD+rVJavmOocawd
W4O2ywybYeVfb2049U+yWarns7encOUInFCcIaFAWUlX3yb06nK+c66L1Jmr1/cd
zndhtf+GaNysp37j14f3LPeMY5TMyeMDFms3fgotGStjUE2Piz9A8c/QJuFarOKF
QVanEgOPWkLaL0Afq06/KjcZHaW2LiScFRidu0wYDQyuWWOxLnFq8yIv3ah3Z8BQ
fFmPhwfIyafW2cWup66PJHcOoRjz1hD+SHHOjCJ/PPoFzVH0VrVQKLQ1qr5PWT0G
zZ7Ek6UCbd2rQwwIuOYya7/1sLwPRFYNqAkCdo5K/qExChHjw0d73RNNxJAxvh6O
AowMgMB/Y6hse/H6A9hlifDVR1gmY6h8SJjSSRzcsFjUhZUv6NLu/Bq6QGW0gEYC
6Q447BFqqOU1+NOEFweQPdrzp7t/MVjFwVVr26YvJ2W1ujWAZuEV2+myJ9yqpVi4
JiiBBPA+XmYEkbCUAx3uvfu44dwc7wdNjB0VmUE8tUZ70/6UrsCRaAdT5/GQ01RK
Y4O9B4/M41zAyS64UaO0BMG6RK4Ip4zRlq63RVb9MiPd88u96CWd2sM6c/vFbtCp
dI1x6s+SC+fxHbKsF5YHApB01pZlTSTIxW6nY9x2GSyxMr1DtlgoQBOicvXhjlWI
VulbYa5mypsSAqEinZxt+O+bveGTBq+MPbQFP1q1R/mJf9uHGtRwvXu4O8yuaqPC
os7X6ZRSMaYOs2/ooNd/+xfD5pHBczQT1hsgj/ll4rhjBVItmwESAJcLRMRvxhiL
I9X8TyBym13zv9hrP99OP+XNTmWhXRCOkCXtCtR15NnBLMgOmdwdu2oICSad4m5w
69/6oQnjKg56/3lwj47XXcAjTCcku3q/qPgg3ELYx+xOzglqp8XnksTiLvmPDt+Y
BsooozTfx6aQmddltjjArpD1oOu1L0XeseJHd8eyR79fkYPcI8mcnT6uX/MRdfDU
EkyBrYZ0+NqCNSJwvhfhdXuR4Mk9KBDmVzn0D0apkHi/DO9/Fj6x8gxbo6WZXp0S
vgl4RhVi5MjG58PftDkgh7iQqozyyIHcwSuI8MuYrX64Jg+iQt+G9Ttp9ax+vGmu
Bp1+4XTBktPC2yC+e8ra8NkySthggQ4WJttqKv5fLg3zDDilkqiobuYTr5ZziqDM
k9hrGA7BVrQApfDK26JGyckfaFL+K730frTFpkpEOliaCL4FokuKEiuww68815f1
01CST/J9UXJxAQ+wBpBoOYzOoO6PoJLqANYR+/KWgiRT+D9bO1H0xhvjVITBkhpg
DaS803zOMT11XGYEWLADX0sbbKxR1VdZ7ioGIA3jb45wTecdn3wQxQZ8fBIjdWOD
FPa3OOlmrDacrKKGZUhlvTleon511Jclj+9FTZvfHm5pDK/NyvrCJN/oX1LSNAUs
zYiCmt708+xDn3s+Zm/MkKfhxGnawOx+T77gR/PGmdcge8iFK/3ju2awOXksMjDD
TJD+cOFrNZwWILCgUW8aRJlrpK++aQAN+7wqqN2gaO/zK9mQzlFbbXid+VydHohX
HiTEeK5srBaj1VfZBcaNCQZYcQS6C2THbTZ8Z7tM3yGXS8n1CvidotA+gBZT84JG
yuz1dYZ+8PIxzRTyldtCBbgUeCrQE4Pn2Hv1MWL8kBcN5zTyWGw4kFMh0TK2yeGS
uFU+IthC2uBFk+QWAun4CLsloYiRkTaY57CwwKdjz1X5URvRWb1msKQM5Elvx8cW
JmDpi0Jb+WmTBPmbF8/MLtcE46Lw6X/l6eg8vkVHnFrIkY/seOufnitnKiek6Soj
aejboTv6GOk5ZcqljorXONMG5duT9HZMP+3LkEZ029TErFu/87GWwVlcGwzitWl1
VzJLudWIWbgE1quouxUl3NQ6Nw/eCPFAnSvXKzZSQeU9LddOadVyKn3zJJd06n31
Ih8s0chpE7/MiVs8qwb2Nkr74NMaDS5Zv1mxnJ1Ht6Qk5NvZhCAJgvuUEgM//UIl
cISij1OUC+IGgZOrM9oMAzlVF0kaUcegF5wc/0Su/vjYsqky190KQ/SvKhbd78Ew
08xhKdcxqkkQxg42Aqa6iSdGYS+DhFdegqUH08Yankj2qtEa2c3tSihEtAl5t2Xj
Yb5BFRW7wPJMTK3PvUniWcmjcjE5tDUHUnPJbrVdHARvdZgdtLkiNc6IfoB6Am3p
+zD1CJNIzWnrE6AwPc6JJn846YQA/XCI15yfhqXLzz+CCYQh5mfKPImaJD6aMuml
okcTvNBDxw962+uK1Bt40zwJsodGUK+7/8XMwLR7d2dw5zlj+zEGR/xB6ufYgZlp
JFJ4Za16T5/IyZT3KcSQyjYC0MBfZler/qLQCkUntK1ymdo7hiwNy3HFGocmn79X
0kDFg7up4WUaH/S76Pkbi3XMmiaa0NVqy5FoqjCdzybUk3wsIUGgPuRLpy4uWOj/
i2zG2i6j2C0hiFBoDItyWX3HKJjPGj7ijkMYfV9QD4FZoIb11wGnMEBQgTh5XOJ3
DTFU4CfYJmM8fOtM7zBk+lEaGNj9q7Vb8w0I7zU00naBvXrbP9NoiRWAdn0ZzvSp
vZGpicLvF4fuPI8t6mq8JqMQ1/fi0iCBG0JVFZAaocVI1oFOakVLsfJCGpfVqN0E
u+OYbCMMZrnXmphiQUMtwXdsnQUrn0rNyPnZVfmlcurU+FhzOS5tn8ri/1/Ho3JG
CTjAcMMoR6bfTxSyaT2rq9ruf9qPYP4ZPbz1w5cM9ivDs/+2Drewqeo4U8JEeTHu
nKCCzXaj4hzykkTlqz0F7fGqxeid5QLP5nGxwJ0mg/6kIs6Le+5G6sVUIvqccw8P
RKrVYR/0lKGqwFhuLz/ggwKmjcF28YaJmDzUIo2iQI0iBh/W9O5Xte8+k5oPqXjI
GN579CNqsY6MU74ZoTwIc48M68y2lrHT/l+muGfX/Ir8CF5xxvMSv6kb+keTEil6
kwPo2PTEzWC92MXma3SJA2YsPq82oGRYihINe1HJUZO5r+vByggVmHTZJg1ZB0b9
3gnwHVHyS7HULdVqVItN7xOnfSQgi65UPJzY2GjuoBGL1JxfAhy/8OmAKK6troUg
yKJVKRuC68K87XywTPrIuxr5OPhs/LLV05ErPXFDfSSBW7ZP0CuaZcq8XUvob2Lw
YZmJZxMNiuh9Wi2rTJC+MmsmoYyi6ml0I5rCM4FIUALF1euJM+LyDdcEJJxSa81o
8tl/OzejTO6jfN/2h/Jcsl+1TvmSkDzoS928gobWmaJAP9hK4SEh3KxAkB/8yy8d
vXth/a72BaEwQgbbww/zfTrhESyI71Ev9n1E77sMFIcZ1w45PYKS/eieKeCsVaYr
PQok1RSQ5q2YPESpwSJ6ls4Hh+ZAHtmeDpd+ecUvcmZ3GjcV5oVr/NDjOGMjgE44
W579WAdzWCvFfCL7hnB9WbKWEm0Q2tNHfuESd+ywu25VpOYaL3BzooyneY6i48R7
nqgJ4JmWfqbxbT4AGkWjptUh5qUYMQxPYFNXZ0CC3Ecr4YHWCGlIyph+fnJ1CkTp
g0NcpPf03GoOOSJxme02hC+fTrKNDJKApLG82npVV5HUN7A/QMk4X8BtSwJUA7GT
LEZ16M3D5pvozrwW7rxQ8Yj4q/yaxQJUb97j8gj5thL6eiwq2LWf8BRJi5Zg9BQt
hJXCGfPjI8S4ZmO9nakqxKBUACnGFzbBp1AR2g+iotYRFI0s56BROF6mTTqgHfvO
g9Bbj37m57Ym3TlGxYZYqgm/noocj8wPWQpbr5FmfOfM6das2wDoluwHnhrKk7Bc
EU81pgxTE3OI4o2mtqeRqDmLxLGa90bS/pynC7TpLpG2zQQIwpStMkGp/pMhOA/i
gGq4YmFRilRRXUkH9kTfN+y88g/l24dfMeuJh0H5vOLFUc8Tv/lsBHKrB6BfAb2w
OMW6tQNPtsw59GX9tr4c4Qge59Lopovn4/oayztpGZk80Ih/MVx5xJ7Um4N+0TpT
Tej/Uvvl2B2jATbXzfqLS3jpIpPszqkN4TdvoGth9zeX10PIP+XVmufiQY21iqed
UY9tH5N+Vf8WfLO3SB0OqBDWZahd3vXbiXGA6KAHNK6v4XU9+s0ImXjFjM1J084q
mQqEHj7BlzclT3A2jPVXoWn0ZL1p7N5RLmNHW8oS07rB7Y/1VOiyZyri3lsEgzG1
WqYqj6H3hgxrsZl/BS5ItshtEyCDFNRE828+AfEr6c2tdaS0SWhxoZAMNCiEmTeK
uzFgEd2qKsfLMgNtIqShOItEvElWsB7acanhjUwW3KIztjaSidhV1Qe/zbXAORvL
QYD76caDMyrm37V7Lq6DT15360Bn3JANUYU52aIfW5VtKUYq8ipcJOOgatPV19hV
OhqQRvRdYZRDtkrDSHMe3eaEIVFqRIIdgnc1YCmOKQBKLHZS+rYxnUkiAK6TnHCn
XuCaO0+dSXpNh3b1+M9EFhBpMNl4Qx7TwCFhM4lmoqESelNmAS2llDCwAdzPtvBX
gQU0kSi6wCpw0//gY7m3+5PZJyGSHVL7dcNZuZlBt9G94FaExhwlOwdYgPq+bjUc
7b6u32Pww1kXpzNhmHQwo+9juMBBb8Iq2uv8o/mAapaPAzkVQM0nc1OUS82pf810
cZXAgWlXw7E82oqH2tg4ieA90sLslLC/6Z95fcFrpanxT3UrDVUi5DXD9mVvJZQs
7U43yLp3IiykNX4RUEu80zarXBaUkgK8IRTXhmP0pIK90qHuOYDzM2pEcJjSjuDu
KILohfqB+t/+AOUzAbrC6+hbT81NiHxwig3rOD80e2Ocmt1ZpkE+DaqARsUehv7X
PPKf0VCHzKe65nKib7zZq5TiBk8SjAxTJVmms23/+ikBP+goiTcamJ5odICzo2nw
AsQgDYlmTem1a2GkR+jYAQEJBxrAKqvJ1mpZdY2aAocDqKEu/UKRFz5cajENJ9OL
dSQxD8l2AZiJEb8mc4CkNun9Fylko6ECovahggQEIyCrHRkk6IHmaCQQmSCN+lX3
Wxx+ZAMHHoL3kj3UbpFem4SJV8qtoZc1DmhCeTuEYqqOQy06uae/trFwAx4nwyJs
xfq/UPjpNV8SvCpwQ8ueGKDzDQeyx+xFuCtcTHkCNdjYmFBss5W6i5h1AHh3Ala5
OmRCyPpKthyeR6yoL1uVSDJVis6uERsVYaPznzPL8BC0qQOhLF9Da2xrnipoUsJ+
iVDos8P9/IhkSmPoutJCUv4ch8Nq0Y4VifTsb7qhqHvuwUyxOCkfFASN3kae4clx
Z1p4v4fvWqI5lXxCmOEkHHdEHVv6ljCmPOrF+TVcu/iifpVwK5hVCmRa0GjNMJWK
+cxQw9iabNpAdTazVPXe02kdkVnA0+gfBV3/3oBSEFavSr0OyEJqeIaUlJS9Ot7z
SBBy7rXLiBHh19C6VnjERUVFecAZXZ4BG3+vDk8ejE5TY/4DXvXxaekLoPALmkAO
5cIOkVdT20QU6k7rTjkjxo4TkHKDmyKgZaDAEQ0H/779kobfW8g+4tfxB5MR74Iv
U9y+DU4WYzx9lFqELUt6GJ4ew+vVmmUGuAA26XVPiw4+W0tFVgvtrLaf0YzwdVVA
crsV7AuSdL0SiJZzXwvUYn2X2jZSsDCIMty7aX24tWkH4ymGluxC/ajr+HZ1ezja
FDB6oYCukqB6xnGMbequdk13uBpG6QVEd/b6HJpp61dw3SoMD9wZsnh5LT26/s9d
ANbL1OFQ5t1lFvM2KxvQQKPV/6EDGbYjW749bBWvCwUn2SFDG3CHjPwXoe5YaoV3
YVCeKj2KW6haSRLvIkUaREYjc2cPENAJZ1domVVJi8G15roH8rRgBpkuhbq7PPR2
neV6MuiPWYm/NgEE2IN7Pwt8UWAbejl1mufP3QQq00dmhZqeF5UJHKAEtvTvN4Kw
/JLi787vgJfsvwgqFZd5ykK9CGXUphJrWujT0cUFG5IGo8CgRF6z1A5GFi352P/f
d2GS+e0RVR/18nZfKJgsE0zaim4FVJgH0Vzg7PNfJVI0LNukptDMcXyUYCOv0+5p
hR1xggoSn/GBsBpUmLP/CnFG6XJGpoj7AoAzlwNv2QwzBzQEfSHCt1ic8jcbo6AZ
VPh/xbN+ahnkhpWmBrwFmYzyXgfxqN0g0soWJO7Tnj13XzoJ7NcO7lq3qZTyeoFZ
oDLJ4DqOWyk2F6Sw4GfEFyMuTTD+fOziBLdGqVtPKBo/KnNd+tXrDI4ALBjO19FZ
7Aps/pAfhmyCDhFjPUeHQ4ylA94KF7Im0u4xYwcmrHdCoodPtk3xiMeOKep32Dvi
9ofbPpsWP1MMlTTUfHxOiejCCZeUNlcVEvYqv62DQF3lq/BAWN15ijXjqBGqVnON
w5pRoyDB8xwIPn5VUaIfqfiAvU+WPkLwNbQN3kSkP2q8NuKkL0nNTPlDNbBlIfOv
+bB7MIyeDa5ieQOx3kUc7d+AMi6THq1xnIMij6SsN03maBqZa0ARtbs9uaEVi/vh
X13c5aM2k8obLYVocs+aAEU0vNqd/Gm1Du0+dXekTEhc081/dfNf+7ngycBKE9jL
5Plr7w4ssUMzrzbWtMA0riCq2up62o1PoSFQvYZrobaX/QiBUQDv1OkBb3ZoeTT/
eNS8X1xc6IifqJGraiHbRCTrPpw05nqQ7gVXUdl+LYzmIA3eh+nXbB0ezBNpizBg
eq+0CCbecOCWepUYOLNGSzyt5GD+t9xVPeTEN1Qht+RSFn5SHMhRGK78CSLDPaXp
zBYqQEnLmiSmEv+i91lJEy37ByscNIhhKl8JrA5ONfFcjd9rIcp5G+wFWbJR1WmV
TZw/aYyxY5jrZcBQLsR9dTZggj6PgvTpHs/NQbIO8Fr2OJmBviXPbhzLbtoYsTeK
wjmqihXMO0/v+7YL9xn+q0digPW19BMcjHebL/BNdLlc+wyAvSSdLKyhywao+a34
mYGZwl9VPNP3E38g0e84x4T5QOs/aQ2pt1MG2P4igjiEEknZNy9szoSRx+Z4fMFt
d7dZOBkQPH3LRtKXAptTqBbQrY0tavb4bOoPWxrpQC93JrG/ab3CRHp00jaoiDMm
bS3+w3/HIvP8fXq0SH5+27lxn6CTLwXO2TEm09GihjkQqnBbXwEM9Ktd8Arhf5EI
d4nOM4JqeQOxH7sZB1OzhxhPPTclQZA1eF7cvr7vxN8kdSAWxi8kCcs7DJ1xt/+x
Y5utbFec2u/XpDfXzDKz6chGU8il5Vj3JXEoDS9kkkbdaigvKKgcuHYSUJpwEVty
nAXWeHMPmpm6QSX+AhMbwonE6oNExR1FHup7Fd0CCNL5U5fRmtvSxgcI+1KHKmHn
ysg8xC4WBK7lgCwu+lBBXnd1I6cuZKNGA61lNhFPdYycevvOctn5ffAgG9MK7KOn
t/wjgsAk9FQF5fXJi6t0M1H0o6F3xEPmVPF0bnLrDG8eKLnyW7/4pBQ9qMYsMmPp
9BqWW4ut5asN9yaAfgNeh82xBpoaoFkLcBqkuc0UE/RkS0uirW6Yzd3h0T0Xn+Z7
x9zvPbxZ6nvmUjzQpBZVNHeIBwH/ke2v1fwgDUnohsIywiyf+0+MlPALWhqedkJx
gKpDqKLbNKci6MmRtggAsrcYs//+Yi+48cBt9GH/4eV9YuUA1niTyWURI5wqhxHo
FdmLw3TnVdGe443aCGoKYl4N1b3lUgmPj+9sEctjbD4l2+UYnWROSy0girypYrG2
rxz6H5Uz0Tm93hxLk7eIcEag6yPC1HFUcnsH0fUuYq5ddzfFXLJbb4YNmTAREET+
1HeFUG5gpj92Rp8KoHtJAnNYyiV5LyensFzcqlnKd3vur/JkVTiNhWniFzvhL4lA
32WO/u789r5CnQSh9cy1OmvJpGsxh2HI1PNpA6Zr6V1yBQQD3uWkyEuknfGcdHMi
+3Yn67apBXZYpkuBNne9g7/ijj582vOUtxe0v6zIF6j6bTfJGdFePMW+S9GQ+vIR
EvahFr6GSys4gEGj7NyyzzHQNloQwNsd9hAUX6zJrziae/9EXrf3gPxanHSTCplH
OEWfp6PRsCLTNyxvTNTS3WIhKmCx1NPfjF6Ilsaec0rjX2ZmixCDqBwpbSoPJSgm
aWbvWQNX1er+WCP0AuQVJWH8oasG46GgXbTZF+XmceX6/NKQsbMtxo7jvX1gaL9p
G2CFcx1XN0O80PT2sFCwDMvxkpj12ctqBRlKyQA1Lt7Q8ZsMifS6pg3Ox5CKFmJh
M2eASRrkbSoYBEBo3gPQgnCpsHsNg8dryFp2lhZ/4LVoxLZOM8NJ/Hsy+TkniJhG
1DoxnhE5C2Hzr6jSFZDqQoGeC1M0x7Q1k2WtpmCDgW6QFinJTs++SmYd104QOhyT
c10FR1hdfbstUvyIjHweHPIYM4uediHZ2KekOLbzygxHqQkcB7GeiRqNZn3j6+gC
fqF6FFlqB9AvTyg1F4Q8ig+5o6CVyr/vtpb0oLLURIQkHzGtGRNXYzTTQv8SYMoJ
Wd/YkmvJYHOU0nmwbOhjhIhSXvTyC1fxr/colETabrREwghIDg108uyqOxVjf3vw
spGHQnfARCPPkpIdeH1UBaAjmbxf45VMtsFGtqtI2wJ2e1wzKqwx05NWEKKQgDaz
iQH+5lNomWtmT9CRuIkM71L/GhDuhGZ29NT/vrvt+rehHTbvmFZc2Rr+rqRlnucj
rS9E12CCDPPWk2bYG4JLcCSMIEBqiHv0g8icUoh/+64ySr3xUOZ/9ZQ+1LqK+EXW
K3y3nPRP3YfjiiIG2xBjDb+UNhopHV21f0G1Z+plwSL/7VM1R0kq8gwf6rOjbrk/
urZp0F8O7P5aXbXp0KkHGALjYcmOjEkER3VbY9d6Kl/xHGND/BlGmvtJBQhA1Kxn
ph6HtHB+L/UoieqzqzBujjFDmsCu813VRZ5gR3yqNet0kkgs2Qe4Upz6gISlbj46
KlqsI65orMKp+UUdNZrrE6K/mfsLmp4rwrME8O6yHhbbX29dy7XF9FndjVw8/QVX
+hxmTCZ4PP+VLKCfsE2my8pQ932rA1MzKjaTTSznzfdF0FCzvyCysj3VA5ZBjcV5
ItFhY8mPXEXEsZpfaTuW2Gje2VSKIdr3HO3VTOfAriQhrR5f65EqnXYQ368xps0y
h+0c5RnbQRFF9DaxldXCylCSTC2Iblg+pUQK/VBzZjefNk+lXlnloQ7TQGSTJq9X
FxepL1AnwTU5Pq10vYV9b5QHhQUnJQLR/2uDWBuod1cA1RXyi1gxBOfprXguvgqa
fIcu+yrSLkPrpSB7NRDcj0DEfAZ8Zww5UXwIBJqitZqbFRJo+uAs3PS4W2GDWJ8y
1YPSA89Ijjl3YKkG5KXgvUZI+1P4bxJ2q4AoW8FVwu/XbEcWTgu9xp77E7cyTOkb
hktven/IPgnk8OOxhcgMn0h9IjzJ3ZQ3GQKSmqEJ9kZ2kQiBg9PsN2KPDipnQHQ3
draJxmPZtMoKN6r95ixFYcKzutmM1HeObPAiS0N1wgRfmBTWmT/uqGFNq77qhx0I
IiXOFGj0bcqbNZqEwkSNf4H2tW83VsicjX8QnqEIKfkMrUhxwfh0ENrDEk0LtDSs
adFOv0SqsBp1ek0P0raLML/TEDTZi4iofuydfoqIgKmiigZlxg844zpNYMU4qqjr
d8eZHhVOMw742ISK/jNM4SZM5nTcGvAmuyVJ9DKFsktQUm5+kR7t72s4oCcbdvbp
Zrz3UL0hm2CYURxcWvfmHENRPwNL7MFGjsEMMIMHL+zCZ8/MKeuaQqXoSETQ8ULo
IxpHAoVRcRNqKC+Gc8Nh1+X6Xbnr1ajLAJALNFeEV1RPfyIs5Z4fOFAYYDCbB60F
UPWDFNFn3scHmazSrHNVamyi0w4ULG4mqDLAmLCm6jiKkmem2XGY5nQsmRuMhtxP
DT0a4MxLnCwYjeVvHs5Di2SBgA8HQOUftdG6fcTdLJj+J8jUET0cgM43dOqwNOoI
CspKL/86AOHX0ep+cTu1YpS7k5T1BCvXydhP4pp/F6PfirWSrxCKmmui6VY3JcC5
pUfW4A+wAQv2A8o8tzVOdZa9eD/uAYIQHMTKi9UogJNcKMunkOwcDzvpSg5sUOC+
DNhOc6rDjUieALZARuCjTlwksyoGKTMtglfJNQLFRSCfWd3YSNwoLMIjqTVUPnAr
fqxNSZpjY41r0w9Gp8NFCjb6mrMlM0TykRxIujq5qwoKz8SaeRZxioia09bLOJWa
dIUFhBi8AySgT2TuTMfFoYgVK9YYdv6xX3kp9Ozel3PbNUp8oni9Qybrx7YJZDCp
1v+h4qlWH8HsR53+dDJRYU4Uu/zHP0PPwWmcSy9/03SxDWbWq9t+c6+wOheIAqa+
YCG756LcnWxhkY5QODA04UVYsVjqHJdoOb42vgsl7UC4P+LA7FEnu0vMNOejBVcC
KoPDX2TbULkJRjSvm26lKMjV1YDPvR8F0iwQUpBPxYhPV2f2nbifAu+kcKx27UDX
kgI6pqL+fn48FR+UpKHu4BW+Q6BB32AYNoMr9dxAcTf1VBVbyW2R688P+ebGr6N5
NF5IP4vue74dP65bplqdtol5g8sUUlWdzmLsSFvs6L4mBy1AWMshtmxqtIix5fK2
+dDHSxtaWey8F+skwIfFznJbIxpg7Aa63TMz2gNcAbkYQHuBJTAiiHfmMLa/TUHl
oZTWC7w0KdGUkR2/5k0ZyhR3FXd/XXzt/pfzhOsc6so3PtK46dEkqiGomy5J9EdR
5Qa4EteghcJrx0h4YuIO8qxxE9h+fZIq45c6CGrgbVZNoRSZOEKJBYSpZnyhedcD
lEIRKBMv5FX7RPskR2IbAUX9jI3c7vpmdQ51zi+r3DOpofSED7aE+zF0p2g/FEpS
u4KLSmTKA+Qb3tMUU6ySqHZGLY8GbZMaQl0MIC3JLFUTo9Jq1zQAE4ArMiB/fWkg
VF/e/jaHOCGlMPdAHH8v6XLRQOVX2mr8MwW531IKVaLbFqsKeT/r1VaFYiBGXfXM
eWOKpGac+q/5rn5FZ9PWIhCi6HYMupsivseG0LGaPONtPndgJag45cWLg5TsmCnE
BH101MlFtWHsPadikHGoN7HHeacT1JCn8wCM34b8+yZ7V25XZPGt4U6oJT0Fhjhz
BIinCRf2hPfjvp4T0XdphLrBsxASM7mEl+/U9SFtl+28KehH9m4iDJ5vy/FqoPsW
m73TZUyTi6zpI6flTg4KbEtt6t80FxwcC8O/P7YW0/G1Gw/FS8GKImGSJ6Mn2NFf
h7w+PXbxSBePrDt198zY/HeDPYag0VzEEQ6DizIZzJWfRgebJpOOvuEdwJKRGSGs
jJ6HT4D/t/W2MMtY6uYj4r/gqLu6DzkJq1j/THKi8AeONVv7oNoXFbKPVj2nLXlq
q2A7iESvuHuklP/L/4La4mMdjPMFET+MQC7TXUyeQXEUJGjlUAHphuoVsSpy6q1T
EGchawcEH6SyhwmxFG2R3wb62uX9XjW0sFCu7YLFfZ9yVjnP0c+nOizZuCB7D39t
AnFZmdNGz4hvRALW+WN4iVVsimgVpHg2VxejKBouKoVbxDDPL+g5g+Yk0LxY2kx9
4dNLQZEesaxLGMIjFLlPl1UZQDU7R3KhFzOGZ6h9+LHEmJABlm5a/QuZ4Rji5pis
e7KE7sZASI0CrrPzda2sNUOLTR/Ueg4dbUcPYABbqHjASS13rBY416kCZRBHi0Qx
ErmuIx+GwCQW0jXHwvswkx3TYLwK6YlrnD1RHTVA4kQuIA39NZUwXyShwNep/Srl
aXmKczSq8+D6KjBzkgcTMKQe+A4AQ7Mmq+TH/uuogKlUSLhahjNkOLuuTTqsRwcP
qyn6O57zeGuXnSifR0lcQTBJCrUdcvrfJ2lWH/6X2vF0Jo8VWCITro1xELYA5T51
u7xlOlyiPj5wP9DSdEX2f5747P16l3/x2crnyMu4vGEOFzaLckD30g/iQlUL62Z7
S0Zfm6L8IBKQtmi1Chr0Hp+2jXhF0SiUGAoO4+5UVSSFep27fqFnqKdgGuS8FAwh
KI8a02W6yTQ50jf7nFqZ4W/Eo3Kz5TuzjurJ7qFcPN1JTykQH326xVOqzbv6J8Iv
Krw7hor94X/8ZJKXSh+TqMdi4bLWAV0UL63BZXoxuftv5ftFuEAijgGa16TkZeBM
m5U/gdzHf5SimPiRDj/r5VGJ6nTRnoEIN8xcpOx10LVqbv7W9bGsSVKJzsHvBFYu
uM5kCVviMtoaiKa1MJ5iVbdZQLSK8wtkZMfqkdyay8/y7i6nLiaGWqvw+9r3y4+3
CbLUBmR/RcvjxIZoZysOyYDfhhxGg9amiwEoL2KNrnsXEo11DJUe9YvO9wWUWx4a
ON89c5/bGvJatSLtfsSeK7oEbqNHOoFrQURXfv7bz2lKDpjU9A9o5+h8lNbdbzNc
EenwKPPd4rNp0Dk0v2Z46qeZ3lk51Z7n0JxVolLyxcadEkOTRYMNfMVhplepXTMM
MUbDHXiPq3g75SS0VrCWjsTIbAy/g+c/RNnhfWkzR+esBSterDzzPnjyn8YJyF5Z
FNo4EIn4WHf4d7RFFGWFzBc49OBa+57wGmpQtBSZGBDHeIaaMty781q0gQwJj8XW
Oxg5I7F3sck1pH4vzpLrJe5DJbxpwCPbHNKH13g38GIqbTzC+fL7ILoKPTrcm5aq
UMglfZaMQKXCFCW2PIhtb1geWtRVzxpPnLGygyfqhlZHhhszgRghw4JrdR9g97MD
r+ljD33wRKnxyypAS98nLD66KiC/m3WoS1T9b+kt4J4JGQywvqwcNsOSqGijDwEc
BhUwaBlw59wVF3opiYMf3+HZY0+ANPYutziGDdzP6xKncNrYTL9Zy2sJPbrl1cBr
3WgBF1qlweOHL3ZykpBK3kjOSm5Gu/siRlCQ6+zQ+jdXjfnqEJ7E7NSlKfSfSNv/
2h1XKhC/j70o7sA6nCI1vrwzboQ4DuPT7KMaO+NAfeOKuu+yYBi7ZbSJ87TgsBJ/
aNGz6jI7jrMsAxQet1TWHePlpqe742F/E/shcm6BM3WA3RkVpspjJ9y3NruiM/Yp
KJLY8FUthm6kZqTsJOKhiWPG2USI1nz9/tEQbsiQXm8ENX2y8EuiMuzO6l1XX+3h
TNDXmoeL8hL4sLDf3AYyRMeEquADG7diBIixBbbp3xVzNeqK3KAGzfX774ZrXUOg
D5Y66ukJpLcc3C+W6QHTa6I0s6/ajMHIWMNDmyv0PP8uGWqjloz0Uwg1Ez5UW1lt
zWGGIUMpwuxVfpKiqS74cc1yNCU0ELRmMqNKOHE8ci7SYbzd8TDUEWzGdG7/wylR
Twp6PCWAYKuXDufCh3jFUv4fxj2VIEYtFQ/ho9FuFe0=
`protect END_PROTECTED
