`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tvdFb9qd2SPWXOwsp7xev641Lk7/QupMhRsNKPwFUV8+rUjTsw8KzzJBfPYk27AO
kA73uV+zF8M+i+AFDFNExsZocUr3LIXbg51OQN5OtNyHVOjahBVoYrU7GsQvILOY
7eqQnIwuiMqmoCJkcao8p8G7rjKOchKsdtCjM6beNJqEL5hZDz8YWC1bask9thGW
vtnHE0TP/skBI/6orMp3xREzby/xuP7YujGAJeNckNkiUBrLsvbE6tkNaVgR6wrA
PcNeokZQqbfgvAl7QhO2WD0F3N3wflFmLxyyWe5hDSagxHPUWXYt7g1Yk+4c80Ul
C0b1omBDNrUIOSRlyh6R3+Lih71aSaxq3WtnTMGkN3QEeSitYBsA0OdOOBhN+ovq
IF0Jin2kk3Bl9zFqVXArHJ7zpAkQcZTlTljiopo8r/Cu9vHU/dQqenHIbbSHVDUf
JJ0avXkoAgIzk95NN9Gu0r5hFxmRAhgj1FLo8GeeiBQBEs8wN/FxBHTdtadMI0Ay
NjVSrVDyLjkDkPjFXgP7A7JBOS+6fThYY6OfJ333wfi3YWw9E17zTuxLtcHH6rIV
zZGORcZR+9H7K0OhHZudI25c1ZwT6W7Ot8WB3RYxoLI4lUo4k45zyrd7abQN/RbE
SnHP1C9SCAjKUzm34QGQcw==
`protect END_PROTECTED
