`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndbWBRHzecYnzA+hPks17i4csq3ZaJg8KQgdSH7x895l4Cep8fKHqRiujVY0qd+V
kpHFn7QW0kOPUEeNo81klh2OHRhpprEY9NDktqfuQQczDTXhLqBALo6/6EJEZrkF
IWgt0UI5hC4TsFHlSbhrsZxYMCqYqts0hXNT5cKhJmpwP9qxtKEJ1mvosVvtG77p
mWoFeQ2810PaZidS7x84oQ5DOAHTp3EWo6r8Jz9NWLjxJsQruOm8WYcgbzoVDpWk
orjEa36Ep9Hjql+FBhCfgCX4lleFtDXRyNDT0hixd6NnEGM14uUEusZ8iGvWxTOg
asVWgBnY7tRK0sopo3BGKaWvGdxl6LVbajqEGYNf5xWHz4SAyPFZKHZ8m1JuZV15
Q2SDaMBD0nMNDWuWDzIq9xX0uzq3Q7u/yoGKxStburgxICQzRrV+xCPGOyLT2IfV
6wPuqoTVK5BmfTwhI37M4s/t+7y5gxa1AwO5kKmjSBo6LytTAmMOM6pD4OXeKLeI
Vu3Y//Wdu23IncdZwJz8/yuUgGeHBJIkHOHNXcPLMB3H/QCBfRmum4dfgXB2pLRP
j4GUB/PDL4UZHkA1CV4aAZqY5A55LdOSnH9v1+V9s9u8Wd9Cjt815O0NXEIwbEox
9t+VbZrqaDRhp0Ic0nfXEpTKQcDiJgYzTB8W5A8i6qbXR1IITBt3o6VmH/sf5u+N
OsJVNX35d/5qK4AE8IfV0vH0gx6gtybC0m+k6C3AWLF0vHi2S6jiCCO+kQ1L+9Q0
eIBwvg1MsBp/fLgp5jmPqw==
`protect END_PROTECTED
