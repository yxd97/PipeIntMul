`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0mgHs3s3mbQ2A+A72ovaSEgobaX2PLRT/aNEYJTYoGIqtNJRxqR1f/m7z8pc6MT
oxCmpW891ok1Basd8c9JsRL6EB2d1m08EIRrpf+PO/BUwUtkSFaMMYUx40i1P+QQ
A3x6eMyGNdCQYwawcTHHccilVCw4rX61oF+Cwm6xlPuG4bmC/Vh54H0i9/lItodI
tu++/I7prjPFV7t5HLf9PBNIXZCnle0S05LqtoL1t9+TPh6TsJz7i6BTlIhN35jU
DytaawbWA1JuJEwWxe7z3WdVBSfkp/JxlO4gReNIlBnpX+HIS8sZKVd9+lS6vMGW
yurSEWCrHTiCcEqomZUTbovX+1JoCAh3eBkvCQtssQmYhSz3QyJsdDNQLyZsd7z3
ZabZUFtab/56ehqMKy8hSxaeO15cuRVG+t4d3veXyXX1CZUbprSXnIrnK/pTlZei
8HKKwjDO6fxF1uH9eRwdWqbAK9vr2kh5DA8YuH4p1hkmHtai5cBR+6Yj8Z10LofS
`protect END_PROTECTED
