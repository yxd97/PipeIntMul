`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xK2VuBaoM8tCAiKirwN+p34JS2lzhqBt3NVSCKCSUeX8VrUHbOCbkQMG8qqja3pf
0nyCYOOh5Hbv6J+dCpn3IPQ4l2Yf3fCla1YTqwXAvkrUEIHs6i2fGk0XsNr0ksH1
U+p+dp7LDiN445wovqpetcN8rHIxSQAcwmFFdJ8UMd9l4HHgr+hAuDiIVDEF2w5k
10h2Vj0HjabCak55iMHEH4s/KWS3V1N7NTfDiuluiCaxTMtJdMcD3HC0MjjMzBWJ
Xg/s/r/aJ3y6rS9JB4kXx0XjXUO/E48H6t0qEryoFlu5QEO8xS4S6TqCy5Bj/E1U
iXCDzcGDSoCjWjnNLNwpqRfjXoMlDCplAtYbZhtL3d6aUyXS4WZyi1SFFnOwOrB7
UdLDTZ/rYqW7XGM7f7Suu69Y4xDDgPd9MMySJ64yGkjbL9fWRLWUA0dmnctCluYo
fi4NHomm36Pf/FiJRoWllVBnpfKm4EanzpCbk0J2pWvKxHtgNdZASNdEg2+oc7DZ
Yw7xXa9BGMn28Y32Mkq8CjKM8hiPLiaCgDEGGpT/hUxVXrcVLoYi0QsIy7NFEKlZ
0sg9ad2qxdox41wISXa3KwXTBQTkRN9AkzIgugp3m/6bFmKofCzCoxp5XLP6Bcfb
bFkrYVo/SbgGOvYAUpLU7KVo3a40UT14SgH4LF6vLcZNiw2fegy/KYp3RgFUdAc5
ZLcgdNBHnwpUJ97EDJggQO4cQ4Rg41daoe+1ViZ0f3JVDw/cqqo9SnAQVxeWdnxY
qMGvL0J4V5e5X9yv6n0c3D3ZR1XMFy3au7h+Dqt8AaA1wJCEDjuWFVHZdRCFg4u2
cOndDAa8HaCoj1Lfy6azAyV6kw3PMDZJYas/mfLbUUjJISSTqB2XLow/CCzLspYi
8DG3YMB+FHh3YwoaAhnUMUM4qP8QVAoJ76O19MZg7vfNd8ONKoP9ey9l6wC7oOk0
rCtwIzngBsseafRsua6cRchWXQvH9qrbvjKCkmK2rQsCaE8omUR2esD59UzJiheA
g6zJ2NbyRecz0LumJcCJfUrTdAf9f+9zGYMzMIRUGf3VaII0t8W3QpOx1Hseaa0s
HhKg7AgIJdddOloCResXGVlfmwuvXkTTrr0gVhla6ki1LhcKZmBX+BDuRzNsFU7L
8p3oXSyPe12kB82SuDYpTwTIvKXDegEx8ffSR42P/Yc0IIm5g1e1Gk1eDHPeaqaq
5dmKhd3ytty1fmoCaQ+uZl/i6gUlNpmVPe/fBkTM3oMKBNnWJ8f+aVSH5ZBHyDcX
4sZjU5jY5bAIbDUqWYfNsyAulifTchilF//v7Tw49v0BVniUrSj4O4I/hAnxLNsL
QP7A3UNK5ycNUiD9D9PjRSIvIvJcVQ4cNqfkQqdunUbFetpS0FIpRGepcBAzAL73
+baaJ0XCdyh1qefzBqFA6mSz96Yp4E5jDTXgtzm+RUPvwiagcQErKm0eCD9j1QBi
NIBJe/0yF7vnwWhdAWXh9I6tcP1X3q72QgJaFPaL7V59L7BSoL0OIoaeogCZ5xGa
uHTYmncfe9d2Lt0MStzHb0RQKDM4mr4hhn/5QRlCdokaVJkqhclSlGHqNKzq1siF
VE0/fIct0yMkCHF+QzgTjILmNfQO7cjZJ86IpOBcSqBNjxVLKJ9q4WuxJcUMhR/R
HP9fc1gxf9jjpJNiFhxW7cir6Q2EfC7KgdvkCkYq6oIpAn89xbWfDPe1/yFiSh1o
chR06QifnJOgQdFfW9+0BWKuCOEbsiQFa50HiBS2nLPQsGxaxTdBtSIjv96w5jVi
0WgbibFmI5X4kjpqTFZrE5v7viktAtuCu/kiOBItD5jdc9CnqdpIzHNigA1Fa1VG
85WDyeUXv2qp9qR46spa1u57da5jusi4iVnU0cA4IYci5a4Z2TY2m1sZool0nqs/
OcuQzuwZjeKXKShstP7ZlprSi5VohueN9utSsqBuR07WCLnletJY9WFCTJuWO2m3
tYbeijYLarrvr36S6C9y2h4jFvRePAjx9XRi8yWPOYudypJT5gQ6E9N5kY7UoDXc
TPKhmddxx5/rbazYRJ8uN1JSXUjhRle4RusuAobImht8qwKTQkxUj8F2VATJ9Agi
s36mcDUwVfIfKzUgyc0lm4ZxOkjk0N5tFLjq/ZsNap7hY61401aWryvxMjDHUUfj
eTM0q9wU7YgTrdF4s521XrRXmmk3E/CC4nTygYiI4BmzqUZSf0MXi+JeB0ABgrts
K+h50xz1XxZ2PxsRpk9nKUmZ0o/WXmnwDt8AuuLErIgVlmiOr2mLK2a3dCY20scR
mItoyE07OpfXtkXcohx3SeOnSUB3V8LExNcmNcQvTK8rZyPxXrGAsMS6pfkx43m9
/3R0NSU0ERuR0VUhzKuPO0M83CQMTiUqwBBH5C1YkJNEcLZMDI74+5LYeP4aYYk2
xnXwU2PaTthEqV/GIid8vj3Q65WYLr3AJA8lDxLN8Xtu+fc5d0GKKj3YbLtYXKDV
LvhjnitJmoyHNtKTemK6mYZ+GZ83NxwLQmRI9zLbXsOGYJWJD6vEY6CaSgxFuWmC
+vFQcKVVIeLp0jVyGlztFli1uId+Brw93LZahFWN5umorUSBceGM57yU1c7iiNyC
7c0Xzs/UiiLM+VGGwaAK/sRxeRlbpOloXBuxkILWdgMqgm29FkD2sdthToRFwggm
B98mUbAnHFDxFGEvKCRYAj2XJ+iWsk0QYb++bwuqJghSvByYRmpSWDzjaP77SoV2
m1x1JnleZCcp13bdGF9o1Vy6GqSfJTCTWGvbjLseM7Ajqe9uo9dvHMr9mM5SVfPQ
CXGzezSukL4vmICLNoASDMpwiMaILjg9K9cLI54GRnhqBErXB82HHI7CS66sraE5
fC2ohmNh77SvhgPRBtkMbfPxuk76IEjELbKv2bypHa8+lO6q9RBMhMqxuvayhB0V
g9LdnVk9iziO1z7RRygt6WYPrGJxsZH3HbgpAvHit3nILKnUb0WoI+AXeDKN2FJa
8Qrf6zMBdjeACcoto3wQMfbx1evnYebinfJc76dFPlwVfPRom35ZVfP42zYVk5Bx
pK3gIBMJEAlk+7Umpx1+DGC3umQhVRnNFmPr+euF9drWN/nvAcIFSjf4urqvjsp5
nhdjmMSGg0Gb5uLJ7cemXY4yHbYDt1KlVgptdFH/jZdqSBf4zjtiC5cCpbt9++0U
lBK3d5z/wJCNtMbCBdd87rApquJKvaW6ERt0ILy0ocK5WRf3LjnZsGEY7u4P0Dro
JId9GZaRfSt5I3ePXcDED+1QLorgUgiImLT83T1crEeGR6uQboTRa6TkGkXuTK3a
qL8HFLiK5hx3iJDxBGLQPDFK4Zmhzasf82otfX4VsrjwWUSKah5DVMFUS9HbbppR
7kiFIv7v66zxmehDwCtoUW0y8susTwcOzTKphDkdcwrzCMAl6GIYVEz0KgEU832K
WFmIterXvLcXIOZFwvP46ETXcNE5CHSrjqdTEKdkz4k3QvCA1dnKcr6RIqMHCWr5
3T1BUFfwX3rprTMppdnc+I8fTYI8SgNzTNj6ztG+PWTmTerJ9CeyYncGw8lvsZ4g
MIrdOcKge6+uPSKW3LtuPH1cvQOJzQSwy+Q8vkmMmengo8WKHCKb/+DvbqFZ3DbX
EDvCY1PxfXeDqD8DcqyjCwrig9q2lnT8Fmra3WnZc/R7uKBe1no0zo2v1PK36Bq3
Engd7l44xY6Vnzj9Oy0zdic9Ds2gzJF6vpsnQEuYk78Q60vTn0HUN8u1trLtgzR7
HWetrYfd0nPb3OjfFj1GWUBHCt6pYZ5Q5bSRHFc6vEeWl09tXcXmpJifjm0HSq4w
S/fKf2YXVlfRRQDizeIdYA2n4sdRMqb8xSAPzijtANY5mviBmy2FaK1M2HvloAb9
I6+OwePzYaBKbFa+OEv1IkYAVWEdunehyp3iI2O/00Gjg1evFSjEVYT27dR2H8Jq
XDBxcdNi1zV4TVKLMx6zz/iDb2rOZl2o8ZVY3AsDwqSvRXoRIhvUrQNatUVNlwqV
/BPtMFhj2q5iWio/fdbN4c2MxcB1Y9MNeaY1M5snzS92NuHtAjihhEbiAo6yWmHi
NfewgT6t34rCcSygRU6EwbvrN1Mol7GIVwIdWzhgOBH+xwsuErZHDpOw7QYFjDCG
tYMBGMWk889xIk7cQKrJV8ITOlrYR9PqFyfYLjjM5U3Fs1cgGLPrP/2xH+yRVLVd
giQ3B95m04yqCMjLXt5bRLAXoEORjHpmJyY+2pO/4KaPqMlrVnix+yMhoviiJQBC
JT4l8gFTDJDho7tvPqjx5ioqJKC21R/qNohme08/WHAuIaAhuVjFqfjb2ruVYq+2
5P2QL0+o1/EKQ1SE/WmpXNYd4ZOEdrimITXy8sgoQSM7DH0lD5ntKQr+vclZ27ya
mhnjNTMxX8HBJc3NyEw2V7al63/GFMuzOO5vuZhQkzjdfhMsYbee+Nsyq4ZaJziX
dMUoUIn3A4PJWLk9Ud2NkhFK2FoLa8C2Hi7kEhhIc0VjME9z/z++0dk7bKauCTnT
1mQpmH0jquqmqDSIxQXq7DL7LO+66FbEuabPdXK3bOOl5xr3a4CF+Qy1BpCJdR/+
VQzt9dMVDvzZBMcLCKJZxZQg7iqHSP2geDQiAlH8Esc2LGF29UbblwL5IrSMma1A
XbaOp3qCu18oYSwPztiliWUJC00NK1Enj1/8hYLV+5qYIMv5vyxPFqGn0RrSB9II
8+8d5PTu5WkLXn/hx5qmqs8CrGCRZo5sWznXBthi51M2ZfuUC/jYfCM05GeYH+af
9Tcoi/5RMQ27+xRSpddLsFzjA4heY6lx1VFr1IYljB8aJWTtLlosYieKc7aiPSuG
LS+g/fqtXCuG3DKQMNTz8cM7p/8SXGRfEEeulVnql3VTBv0/raJgp6I34y510S4B
a3WAufabylFS+1O+RhYMhbnB19xKOu577DopL9AHj1NhZsIGrJRTwDGkLQsfTffY
lxyCP/kS9NLavXVFttgQj+hihlverqDLoakj6MqYv0u3/faxGI/+NNs5OS3eTU++
7uM8lDf4i+id/H8zrGiNgi3v5nx8caA6JUJOfWLg7ZUvuRy9FIjwkxqBrbg7t/x3
XKe7A+mKzONvJ+wHr5RuE//RJi9m3/HJXoLzVRNb5nKbJae+T3lmbe70EgliJifY
5y9fuKBBrC4r8z7lEyLPpThyrTGXZIPDMHNDhEUtkne4J6+3e4CYxGNK0fvjOhpX
vgsK2KSH/WT8pAVRRiRg4uLowCcS+AGIVc5SPFTrnsEPP9cJfEc+/MbXZvKOalvo
ETM//CItb85MMAFlxSQHJO7mTbVcPuf0eBndhZYyErZvhnPf4jOULyuwDp+S9gVA
P0LTxMKvF9juVECfAHXqs2R7H412Folrw/nukIvZ1RfjVzSEvtHsZZ7wy1lPdcNe
EYLVIjrthLPgCRwMreMmei2hfCYAEvXpohoKSVGh6EImRmt6BH6bcrGrAWX5O8LV
CgJ07LYnRA1FeyupLVDWQA51xUPIeNFytNo4cjlz20V87K8+jfdQ/u6I1KakB/Ji
Jy7wG+MPJ1DzxDkmWijNzlf1d+KaydQyBMdbBHfiajyKR+GHuktr9j/4/+j/297n
dD6WlrR4H9R76ppyWMibMBPADPTXagORncNEPQ6sdtxGcgOjtjnFWYeoDAmmhJHf
V9SOflwN99X8FG8ZPwE9KKaa8GFdTjmOP3mA5k4XGXffiy4MLqn93P0dUT3D7Gx1
MwltYumgjzMTsrhG88J3MooQqmveTYfuXT9RZ2kqLJBfqoxZi+VNInJRGCMudeh3
rNnQaYOc2wC5Cfpa4O02LoSVsY8HLIrgzcOStK1CdEHxBE3EN4BxGR05W18upNLK
WivOVBc8yM5FPYkFG3E4zJR0YqLJoKELuSV5Vx7UxYpsqvMsHJlqzM6bxTQ07hTc
luhqmt7/lnhlswyuK+52/R+BwIY2wlQpfUkgL5zka+GYgfItyYKqPuhREUqLdCRP
KxmFWEZF3sa+Q0JcSg0CaTue8/qO3K1PnUOyUoWzVqys1wqakDAwb/5ATFxNVHmY
OX3PG8dHQDXc0FOGHsBLgfMyKlplCymZnSGCJAPE3COWv9OqTt2PixSGwitf610A
A8OX0eDWo0oHLqMr7Y8SIT32BjvYvF0p/8csIMgsy5gsaLDE+La0rbS8OXtKdvWb
Gf2/0S86KA6Nd/33isTKTAFfH1ea2UqvPHPcB290ol9zE/yS1IlOpqy01Qqj/EBY
LEKKV2i9qZjyKMJBmEASscAUP7C/1EE8l9BNb2M9iRrAinpLgvsOLRopA3Ro7tVf
64CY9I2AGf+21RKri2U7+8+yKFM/Cncsb7JmMdhiLZkvPEVBnfZzgoaOK/DpLowR
vV3TUdddU6px9OmuwNCmJ3SbHjVwHP7hxi/yr2vDpYYwiP4u5QNLYso4qEZ+mAoS
cg70uV4p1bjDZB2gMOIdYtCPuD9SAx5nNgLCnCTgUhPiDx3vYPddUPAaDkBlMLAr
3QutpqSgqLqSHcKq8kRdADsx7LXG2isw5pTFYcnCRdpiH3vps6tfQ+8dAl/ETQUj
L1RQM6gf5ElQ0biSPVVg+5B0kAy7Hb0ARBFqebTp+pXELvwJZrHQiDIV4LZa4BgB
4FSCi1VO9ro5JeURkmAI9aZckJvgjYKDhHvubQ/xGf84wR0ST1jLWeLFZ55cGVtG
rX5Gd9U2S2mBFG5iQNvoy7YuGHEsjiEr4uek22dpnmOnbfiAPr4w82zLgnn+nXDG
XbCKFrhS0IWXmbzNBpzTo/nULD83L1IdAx4a/o4LW6GPhnd92whpFARg/fsNUBaW
7mqAhRY5ZlLM6iZr2cFALPy8+csXPZFrUN9A8nOfoLE4ryHIatiUcsIrPTtjNAF0
zH+zIFpS+t+OW58KMlLEhMgxn6oKP7Uh5wSCBa2kdEWmykdqicim1VBBUc8KtN4N
VHFd3sxKtpBUsRC4Vn/LGjr/kSnu8iIjBy54er4+VCsNCbrVZM5gPELQb81IdXsT
J+rxx69WYgoVFAJTgB/juo7TX0RwB/emuBMjP22Wbtm9zkEQnr3s2xDgEsQ12BLA
aLZ1YloLzSVAQf/rPq1LAsFqDY+1I4KGId8xDhyFo0rpZwgMdae9JSRL5bNUvPNH
iq9K6TKEi4l/RhpvfTr3nP2EDulpWsHN2KrexzDbuSOPnBqCk9k/ypIfsm+QqWVJ
uVj0rrKPI+nlMQbnY+1mgLLhcXl2SYzCswpDd450N2w3Dla5QRbXlAk/9M1Yo7dm
7GTzWS6I48qrf7pi1/kYPwlQXo72df8Dd+f9MiHXt3N1MxdylG0OYo3wsTL6+sGL
dRlm3DcBL7DQm3lMLKXa8IewsbV7OfEF0SOWnMc9w2YaQkGSLJ3/aAizhDjOdo0u
bvumppSe/kAngjLxl/mOxc0S71Psk471kgHsHfcSaOY=
`protect END_PROTECTED
