`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOuFoe8alkzOGVmnFxGMRePGvsK18yD3dPn5Ao+m6FptXfEvHCB2cfw1qkQcaqPG
jkRkpo41S6maTqY03S5YNcXPACcYrVK6ziwwajt2el1JiL6Yh5ILVm/o9zkj0LO1
54ted8xAdwwatE8GWwWXJmK/B1f7YGPGs/qPCZQyJCf4k93U351XQarwNETe49et
Pe+yuMlT3oxa6bFQ6dbahbfNqEF0A3Wvue8hyoWugw96ylA8oupxrCQBsB6w5tw4
mLSHq8tz8gLLpMFTa4UGS7jX9+gwz8J8Ics7/APBSn2uHpqcAjHGrX6RlcRtN15I
I3A+Qq+P7amhkHv5athPLtj9OCLuBcn5DhqnUNCJ9dJUzU6qFn9+sXTCFJFagpFk
5VUn4eq2CU4jHktNSLBnMkm7Lg+bkdW5MHfUAOEdoLfr8Nahbim9g1j0geud+iyq
ynZRLmE3VNGM9/JpZXPeQ1zwTNoqfoEbfsiWQjhNUyrT/POy1ZYvBjzvpfI5MBR5
`protect END_PROTECTED
