`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ygxtuIjJSN/BH+Egye6pjCuPK6k4C8Hl/Uasb7Y1scQetAqqM3lD9b1QvRj1Aa4d
kGCXOb5mlBwPOxaS+YCdDtk32I1hvoREll+5UMpWocWx8wUvp2jbT014CC1pW88m
PrO4q8y0PE5nWTXIdmo7ulB/1xW4JuUjTY7VR+NeVkSiU5Uscj5Vci2j3o7ZK1an
oG47X9TA9YviQfPXRF5iAyctr9ZPlklVabcZzni9328P4UQ4LxObMLbwFKTu7mZX
ezM7kAS8+xwSatqSBXU04Q==
`protect END_PROTECTED
