`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MSvmEtzloSuqD8Y3TNe4o5hruhIUPN5DmM3g/ueqkSaDSF/yYEJy6a03O8WuNxoU
Kq6VMINgBA0PCcUj3Ecp+EeBkG+9ozb7pwmF84wjP8HDZNhRNmWfTJ1LLROcxo5k
nKtl3IAr0FYiwDiR01NwXs4mm/TFqDBBXHGh1V03kFM8+DTgurbrCU6sK2RU6eUx
1IQErZsIpcjjSojDfwaYnQOH2LyGT28mWa1XNKFycbL1KNCE0j8m/GPfSCJiczda
HHJCz4jyT3UweoEec0V2xMq2CyCYHvo48m58wa9W2L9FuqLNvE4xaG9XdPih2h5R
CbZcOWHE/y1aTUMVg1qafk+I+W5LybW8Gtidqm11+dbbjEYfND33r1WA3A5E79U5
`protect END_PROTECTED
