`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R412eG4ahQGumIVxXCkDMOGHPVQOwHxqg4jXCJ97tJkFseO0FF2hGAfLpV9pfCv4
w0bHdq5EU9zM8UBZm9KYfb9k/7lZ6O/OJG5jC89UCUVIhItrG2a1pHMD4em0kbsu
eS9XJCYJIeZd0+4jB6cg1ZWtS7yexAIrxNEBnHgW7qDwWAeVNwSt2NurukQJXpGM
1qsTsVg7eakiVw3bpPCO2aIy6u0q0OOtcC2lwVYEb05jaiIsDa5Z9JL7j9DQQfFs
tEFh5F+SseV3ttKSELabMhXfo9XrjfrixVJSDNdMDsMoCg6Mz8SCFfx/2Hz/L9MY
JXt7s+YIxR0Uzc80F7uMxus5QHBewqovgoNZMVn/WYImP2FiHaISTquxmFQoXDmP
lX1L5WV8MQzhMi8prK/+HerWNLr3u+3q2wHGj4X8ayzqOuSs9drUJlrXrA8MO7N8
9Z0DlPziKy0ufHVbSyGGLMf0V1QCfOWUhIRF8gKV1pmiGJheRkvQxrDHHD9tlfsh
lOiDPnDzzS9uz6Ablqi9Gw==
`protect END_PROTECTED
