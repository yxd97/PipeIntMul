`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Pc8UQNNYquzihTZB3/UmTEksWzQagArI7Vzdmw+L2oEDMO20tGw4KLkqiTC6vHF
nZ8dGMKHyGCJuOlfQ2G6Kfz7Bw9LddZ0woOW+FQbz0Nas/4aK64vPphtILmqOICY
2j4GeOZsW+FsLWbhiJFF0FOOekP0SD0xdUy96znH30TvnxVWyx3LRmMISjQ2EN7A
CJqOlY2hCinSPsGkVuoHczZh4bWM+Ewn77ylrv+3yV/qDS//ySbKh3HPCdPInzxC
t1yQve/w7MI3+Ro8LgelCC1dVpyOA9wVpOfZpOm9EuyWzM+CCIpOE4Zk8+sFrNxK
yt1u4h0fK6Vxg1bPPiAG+CYuycoJXTN/yh69kPbCmTmdgyIaspNuqHxyVP6VAvVU
TONbpt2oQDH+llXRNOiD04PlnsSuxpKUkbBlnk13aabruvyVUY5IEwDQD1Msw/Th
B/jkQOiPoGr/nOFVbNUlLvYo28UBsI+pcDEszND+iO2Xo9riu+7GY4FJ83t+a27T
3+7OLw7/60Cyzne52zPwpp8xCcC6cWZTDtrryXQ1WpoIglFtaa8WDTbGMWCLbp3D
sy+ukvFugk4ID/1KuFR8UuL2YtlsMVaWmKNB18Hl3cp48IQSodkqFJlphzJ95Yuo
2oomDpml6yXdlg+msEwyK9MM955avE3xPtDbtxXzbViGhwjIraTC3WnH6Jb0VcnN
oBff2M4ZlvZ3iUtmH53bFHwjLHXWV0RmickdwBcDGFlDeACTDC9OHiVK/EeV9UtV
dizkf0s+cOEIr1jkoTm43DP7iVtXbQS8b5EdQ36Gikrt+NYX4vQEf6pDsVvc9h5o
/I/cJiadHocwvoMGyY/yyA/U1BLcytNWbfMhfU9ENs5a6N10MJVXTV/gsmIYTjLF
TfSUdb58crnimu6gYF1qxt042VwufosUnFn1+xfmc3os/Le6HgmyZsIj8Dsckv8T
5AoXyq+2++86wqYmdybEwDdwAyDP16UL+H4bF++46W0auVIl+T0SJJlQkmvoSo7g
sCHGPleMYmYZsWGMXCy6Rbo0ZMJ57S+wS/LOVNomDhw20geb7ETMdjIYA/iqfZ8R
`protect END_PROTECTED
