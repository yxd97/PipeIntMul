`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0vxJ2ViXlFv0Fp727EDChpAPtapBdXACxp8+u+54BH31VGurIQDfRSUWhEtXcM0v
E66VNZVu59q4eQqWCMiBg3ItIjpkQx4Q9WPpJNqCyO92Ff4yrf8YrhylUL9cdsr1
bcFXMvBn0UL7NBaRhXkW8cKe0R7HJIo2ssylu4VM7JFXoN1A9/+5jzMCl+s+4CrS
Y+44nYr3r2tD3INslNi3ac0+50A0l98E13zaMuQmd4XjUoY6zRTMalbF1sGH8Hpv
q/56hL88yzhQnWtmhh2/CK7q0N1jBRI7w0s1fghxypyujQfp2+nsnA46hqCc7nRv
s1/CMT996BjMDtg5iKLqvQ==
`protect END_PROTECTED
