`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mEgHOSc6jkhxc/gj4e9pJJtc2jAqiURWcjJdhzI1/8sedgu9wNGPIgkQCFRw6SL0
YuCx6xckHvlhHwriyh5nDf41v7QoGCwrY35cHFmLdAZhb0+NAqjWgHMRqD3l1QP+
URnAdK3uiX3c1M9TmKt2Bn7gZH4WiDfle9OL/8XUz6N8QN1KDFxjeUN2Bdv6jui5
Gvp4svmy1QtBJ8MTrI29Bdr3ISggd32fqyTlQKTRwGWzoylSVWE3QfDEsEIEOJE6
4wWeemNHidWpd/itq+PU9zeiqTeqo6Qvjna0mHoOx2hT03WyE5rSZzo+F4Lda0Db
oC2uN3rnZ4VIOWa53jsZyVGFaNB9Yke4Pr96QHXtb1KPnY9TzeU0E1TYFtI+1etR
4XeyQDj3uPh+iiyAy7Ixq0hduM81FUH7BKEpwPKewZIIDc3MhNTX5NSCe/0bofJz
zLmzQQZO+1XxzoQ7UQ2G5BU6EmSRLSpfjteSkWulXtk3VVLoYUNqZJ07A4DrsPMD
YudHDk+CsdjBxAXO3dYygiU+K75cIzNwwv5T6dC+j13+gM6YZnwR1fd5wSbnCnOz
2QvFuTMDdLnmiMDdybeHbZwkjx1kIZnMhUgO2FuxusM6rNThVC7uSkYLYzsP22UP
fo1/uVTf3SuGir/PjnSAiT4IKWGTdr7Hv1ZbgiI1PM0laCApWe1PcHJEJqyPfMI3
xBGcRrPU4sqL4xDaXtDUBQYm+bxubPIwBC8LvoDNrwCiqfAQ1I3U6AzQg2PFYijJ
gMhbO6k/zQxmmrkWYg30Zz2HKCrvadVkwwM4L7kkfBPYT9h5Mz7Mqc7qfq5pQhWo
WBJXamVaslm4Ui6JIyPwI40kpPZDiHTf9nW4SEWbMO7A9Kno6pgcPFGMVqUEzP8D
LbqMxwBSeM/U68uaECTlVYFAEM9pduocXMwowfZ4OBnsZrrGXdGPmpHo+tXGWjUp
nkPBKzPplIrrcFZTqXkiGuIaywJXTA2Azra9PwhHk2Aw4Gc9tjtfToPxk8duMe1d
0+Fcy/gTX8TxI5/6cZTdYABi/DK+ueoCxVXkOR/K8b242IIs9FUNnMa6nJ5yQV+Y
DUhoJfZb28pPyKA1wO46CRZ+Z8nkDhcCae3ZikHaMHMZx9XhSozoPK3J+pwKoKzf
NZbKOdKMiAZQ4M8yejIcSqwO3bhcHgOUFZHjraQBSuTkRn1xyGySZucv2Q0NsBP/
01NuIdauSgiBFNoq3nFU76d/6FmlKmSZqWO6jZEdjP2pn8P4Ozh/M1id7yHtsmiE
T9XUR2Nx41oFQ9FEhliGkOtU1r+xVFhbOCqTnm+TaIA4kP4vjvURJ9dpPHzhvqoM
nX4yyIEm+9FsPrtRlj4mAtilubg9/u7kEtYJcryp6BN08G7XOj3XCNXHB/90d55d
/P2X4UrHDSg1e8SBOgwE2yO7ZfVoJ9nY7a/lkuTDafFJJ73yhkgnU6BBEk5vt6tv
FkCGxWqRvzg01KjkPOdxX9+omyViD7C8/0KI3pAu9szyCZhoE/eKY9sbXDmNgsVA
jiwxX6HhUIvrHnkNrfA6E3RRNrLir7lGv2MN7rjnEqocFmf9Z2oDbh4bWfwx/bzP
PtjEyawkCaaGjB8BWmvur9XJ203FKrjV2VicXLnbv8+eU1Galv9jpMWlViAZ8o+6
oNvY5Lc8+68/IPPzuWHvqSGrcTxDRL/OA2bjcF9BsfynxEjXKRAlLE3inVaKHZxt
HGwab8q0btM0wpOdpH4Z8Y4Atmvfovoq59f4PEXCT9Mgbo394oizB6pR0Olm5bfW
prFTYt3J615yVYmKezlcvLyfMr09mvxOO2jcFBgfoja6hC9aiIS3vV/qjS3IsVYO
SMbaEo3COGornuzuRZa6JezeGeYPyIBpQgj7pfk0eke13QHHpiVnQa/6BLW1hQv+
CMDEZHtJiIpNw3HiJhpAHAftpI2HxUh/9oypVTijXglUCM5sGprvkJ/96eFhhyf8
yLM4Iwk7KfJjd2sXeyyYJhKnog1+pWfPRf2Hg6eKtYU6Xxd/vdw/m8v2Zjv+KjnN
qvoVHS4m7tmkgP0iBXvJpK/qB1lBlJNooXgO+WKInY/qaPrD7mqe6CJ9U6F04sZN
tTXQnaRU838j8dQ2L7pW6g1vBiHR7mvnwGW1to8OKOUYkygg/wR0Ski+nsjc6jdV
fhUY4TnQfOreSAHQ3uzY9GPK7tJTeEvZLLd9roM4LE9fDpfoLu2yhjXfccucd1nw
Xc4ShPVnXEYsQMDtxF8VTIOgrIVETXErbv9KAA/zkgDve+/L13skbwvwY8sOS+c8
HIVLzLSW/gXzIApYpZ+LldWVZz/9xw55WFqdgE8JryryU+aaqpL75tXoYmlx3Z3s
x+9p84miKTsjSEotKlLXbzBs8sANd+PifYPaVV+gq++E+3xl5uFaQSQbhw68iEFu
a12KLNSD9N0AHG5sb7GcXjPRdArrrU2hhLEtEOs5otVa1j1jYz5hN3AmEuoiIk0H
tqiPG2Lvqv3egYBhsn/viL8JiSj8w+mo6o8kxOGsMnmu0IfamdGNG69aNXr4K0Qq
HDtwuhDEsohCgpPP5OTmTIrginqNuU7UM0o6w0lb6kWcQpNBE0JPFj9QLKlSdU+E
1e7O09y8ZW/aS/+M3V1ZVhz2U4sMOdOTk8qZRxVTvAfwHdOQ9K5OhlWe1fbuVSzw
h+aeVnodi6OiGmEMPmqqn9QAa0sNHpCUjJc+pP7rlr6OjSOOEFvyrNiRXb0Z5cyw
d2QZqh9H3oGmpXzbZ9/mRWO3hatSeHhdL8XkgTkpyWDWFYeyPUsau6PPfU61oFLS
KW64GoFbh6tmoTA6vRAemLx5x25D7RTJgl2o5uvGwXdtqgadmmUC2+O/rJqFdj5F
eMI8rztnBMYGIWfiD4aQsGPHicz0qBr8r+euJitlug8fpfHOilrvQti/tMqwp9uE
GvvSy7sRRwt+kAs9KpVeciNRhmus7XsVAJWQTiCKy4ueWjNc0UQeUJBf77ZaVQun
6oVyqe7r7BddPdeOWZF9aDJ2dOqaa8ELzoPRmYcp/FrTp+n08Y3uopLJHzYaQM+q
RbWUG235jzjMLDznT0P+3JAVk8MT3STCVTc1l7GIK5w=
`protect END_PROTECTED
