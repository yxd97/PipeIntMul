`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cq0JNb0vN48cUhn4v6zu8YAE6H8ieGe2OPpvvhDqschfGdCTuoWjeLvV93GfIn8l
sYg5m3DtqZeV/kcLA7CC55KFttr9IcIOGuPSOcwMVTaF+QdJM84e0MFRgdujlYE9
TzxBUr3x++0gZSzJepeatNHmvPXdMWH3LgdbsWPkhmwyqhrl48f2aSFrFttSLRmS
ascY4B/8hxvNzVrkc62S9KyimWNN1wc+4MCuGutN/DQql4Mj+mZpu0eYkOY24nRZ
ISxLn7wdV1X0pSHUhFhqdnHnpsHNYZtlaUQNC0vS2n6GOQHdowUi+63/kINmZ7D/
6+NAccOqqGts0Rovem4XQg==
`protect END_PROTECTED
