`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/urjJspTuq2FOFSFF912Usfe188rZenHE6nSTtC6vnvskfi7mqQILar9k36Hvk2F
BBnm9s5edtSyCWJ/qzOXj5uynMpialUkOGAocJ5qDIfN3Kpv3o6B3zbiq7rd9ylP
ZVsuETtJI1U4lG33p6R++xOyEyhKE1jMXSBkj37JP/cfchomOjz3v4Ap/fbzFSIS
ecqpXun6ese2SKABu5kLcpansktBftBbuu9GTjXYMX680reAFP0rBxsJxlqofG0x
2Fyh7KUMtjWTlJhljUTA6l1bXNnjB20dQIvTTidfw18ovfOlKIbJ0+HvubGf9aFR
Uvwva2u8dYMGYOnUUdpCf+vc7ZWtAh+QxBvZLGTDtpmSiIc/38b5Ihs3qjS0bGam
vScRgcEPXK6/EgmOGIaNnlG9Sv2hJriEEEOq44LDPq3HG3m4Ufb6HbWjB9Zzql1I
nqv4q3BgEb6ULfXs07bauwqvvVcOiZ9MSldrdWJI4JUtkFwLw3PZV546d/4t2aSo
AdwHnxQWc796OR7wPcJCKihCUBx7hc/l5+LyB0cvh6AN0XJvFsh8FfOKfHCxnBwW
rgwCZAuy+twSNtBOoJVi4WmY7D3C509KFE8GD88+PlYQtq00S0+QBlV+K5dHgxQ/
`protect END_PROTECTED
