`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hlweOebb+0a1GVGytkvVqVwniVZ6grwT4rvHTmzbFkGex8mIwK1uAQg48lnFt2Wr
Q3qwv6MbQnC0MbVtFbkRSNiQIxmJdRIFVWf8t+zm/0WDuj9u+wahn1LlXCOTC9rS
Rv0pD7Rgv7MgmULpf/Rh6aBAkQsKMeempG4ZcjD3ymkmSYS3JLfPL9zfC+esh6sK
wO98jJ/atKngxMhRmuishbNtk50QsXHP/tocJw/ViWayTQiF8whkjUIBbvFp1dbb
qm+fC+SD+spPdnV0du6a39DV1lj3MKVDCNc0/WYRcaL8QsuDfpk63gULUQCEs1JA
xrbjxeuAob/s17uOkdQH4vOKY+kL0QYq8knnSjR2NWcadfXMYXHybw6WOke/eo4A
H7L5PSX/aaOq1ZrYM0J9oYEQM/0JleYlxLVxZXCTApEwz+d7zwNf/b2JPJiouiA0
zZZVIL/8Uske4CnBaAKqILn7YaxLuYv7LceuOeEfN8Tb2vz1tBJaAH7UUEkmZc/1
9WhRPKzNk/hw+8JvanEP6EKcwXDo9XfAhwHoIkYjs5MEpRpWsFxkANPtYq08a3QR
jRJ4nF1Hwe1dUfUQ5qgpjoruUD22HwLX34mozEPH3cdZ+HTVWN8CKQEpxXqAOkon
wQXz7EB4wZ4045vT9jApK3pUEleJDSMDDhIJwVwAn21Kug87NrSjs9n1hbnGqQrt
2hvE1poMqsX0iNNtb8OjwSZTQxCT6FQimczT55m5s/3kVMEDXvtSOhFqFWez1b8Z
ZAqC6coFw9BEFCfZx1MByoY1epyXf7FnvzTFDqjQL1MrAO1G8CocL+hFRhk5oNmd
p817Si4qu8Tg1SM2wwX1vr54fcoJotgarw6phUAFEreY3hBZaKhmlLAVS0b9anVa
mFK336hzncWLKq0vnmNHM6mT3z9iE4Nl/wcRQ1DJPvqwA/0eyOky3mG/l98jo0K7
QPG9UjTxWZuwt5eeKKOuDzY+VkF5LQ/OxUJXcyvgSv0F4UtoviCdYl3m42nC+wqX
wavLBYfQYJWEWcEjpm1pddQJ+ZTdXKiUXqpFebNIPwWp/bayRBMoB2JtKYWAJdo4
DtWYKTpIQKULr9caxHuBPkcTjjGzlykhAEEMdHuMOrs/Z24aCw6QT1kks5noIhjJ
76a+WaL0QryI6lyzUajkpDMQTCgX2xiDyxPAgChDdkAM2wDtUpSNJ1e0Hs7D/StU
tJhwJtdgqkRPF0LJ4WnFMDhaMYRD9gYdisVope9eRGSLqvAn8tj+vExRQ75zVC8A
/C4LrPc8eodmpw+wu9DepJKfVi7HPECXM/2q694DwNWdIpoyKarVex8Ur6tqdnVs
1HJCroo5QOUa0tIpn3n1fVmissH2vbVgc2SHVziBC9iTLLmbGqc0woAbh6wOUNC5
cFtXYHQ4MpvC2LSOpTpZZYxzhud7B7I8fkEQtegZzhKF9RMbN42paGwI8y8uFdge
z/89oUzuZrkeuM9R2mvteUxVUks9doOI3sT56ts5ZLKjkcPJcyef6E1feGSWBxJ8
nSJbNrLrhlEXwI7Cbg5Ayni4/lwmqA6A2ss1F2maxqFpV8KrE5gow6JdAUAtkBq8
fLTeadgjsnH0xzm6LwYJjXc+KtiwvOp/LGF+ym3rrg1bR+ALxII+jbqtAgK6B84V
kcp2/dUWF/fDa9eQ4QOqBPPDaia1tfCCoBRMycT4Uh2ia2WlkV4Opre8X8g5BQpp
ekz0wxb2qx6kAktAzp10LelLNFuUsDlJ1uUwItKYwcfUIGwQixnBU/HS2MSG7eap
dR86PhjxHZT623tGZo2NHpFeEWDhecS7LtNkk5SYFo+iHuv4vGBAJI3jhF/T/AXM
T+Fa8myOWlmH9MH0Vt0v/ur1ZaviB6vxrpd5AiZrguO0SiiS4TPh6XVZEWgucFAJ
FNnEjh0hSLJCDDb3z4dIaQ==
`protect END_PROTECTED
