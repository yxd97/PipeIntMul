`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fH2QklJN9KwGVj6sLiIrf5YnUFvb2z9amgf16QO5pOIqHn7phLsSiXF6MEE0of1o
IZrKWl9hXSDpfvdaLRoMItGCdBVmH/FQorLOxCeqMldgYQpeRVc8WK5qU8nmkuDQ
8Nngz4we7EzRFs8M6tOCGc6DEht+wkr6Qt3S5xmiNoWVAuA6wCMPIoSMYhKF+S0G
g9BHe4vguLzINxOSdH4SvQSFfIRdxq+3Kt+hhkY/onNfdrtxIDcFzMW62nrKKqPy
obc4tVikuagT7RpmAr3ib6nJyGx4GXjAIiiRnYltDaDfRqsmNKpNDwprVkb6U8aE
4maVWfGCWjJkYOjr+JNiyU8pthFngHpkrT7MFgMxfhO9Chd1ttFGmhVdl1uze0S7
CHZhx/8Bux5KO4IHzTaMAjry9kgXakxUmboB9Z1ujY5Qsipk7CbJB6WEAmEdJZvy
0G8BaPiRB+1sNaOZVTmYURuhXq3HO5z5r46YaKseI6WDKLie8N+t42bcx0+6FIcm
`protect END_PROTECTED
