`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJRiTD/vmehLV+O7wdHcntCo6FXwisDDlwIcD+ki9eAjywVBRtum3CXPoCWV9bVc
1BpANBKgUoMVsPc7WiUqAwlvDJba4Sa1k+nSvMVfQmNhNdNA3c/eUAj02Qr/Ga8z
PFaOrru0b5sLz7WV2O2skdA5BdMjYy/0n2jey/VjbAtmsqiMezVFpuk75vdbGn2K
ALtbeCH58rc1M+4x/X7zZLuhlrEj3m25GO+6a7pqOFD8Y7BNh4bd5z7o4YqahrXd
7T3KZmPhjC5VozUexcQN8JS7GGbdh3YgfE0pwSDU7AindrIgfJvPVoZA3wNIzcj9
olzME14j02XKNnIVFAlajg==
`protect END_PROTECTED
