`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7tFk+AHvJdZfp5EumrZT9Y29m8g2KVkQ+PlQIhBLoSjHzaXLVT064HpWss250zB
ICasQaXz9ChxJ1CiIEPLrr6OLKNTlGzWA5/r6ZYls5nmie0TumOJAmEmkaykO7zS
x/vh3Gd0rbZP8Mv+Kgb8nwIqqdPrAyCZPb05Obz/3GcTml2i72yk3OgJLgX65BpO
hmmP5V6urPRcoReKu3LQ+k7zTMklsjY1leo8kj8bdfTDrGEh781AHT6grjymmSee
WqUh4d3PUGtvUB1Rq8LBAV1diEbupXt+I4pQx20iAB4=
`protect END_PROTECTED
