`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+d+ndTAbyJyuPHycKWtOBpd+mBDHUqoqRDrFE/7gflSDOaNBlnxuFr7tT3Cv2X1X
fF8SpvbRns1kKm0kh+EOTrjmFfzDb58sYnTPkhfm3fhhoodaOuPoQ471YhA7l5Ka
gmGtkdVr4YRY5vmdeX2rkd1c/EK/VeEss8Za7mOKigJR2hgjrDr31YeEMcfsDvmt
Pkz0Xj7ekVaoqdKt0ND8TUkTkpRSgxDYCX1MqFnZRrlz+3ZFSy6ysJFuxcWA+0o+
KgBqUwi3gk7Z5M0mRE+RhsCf2vAFak647HhEZvXhofyAPXtkTfFxprPyuD7G9Skl
gpWq3L5NK6zbhtf72a2TqEz0ktaogjwxDvv0yc4yJZm84VtP9xnC1X3XuKNxtxhy
wg5woCCg3sn7t5UATRyNxrZfZvUpZwmHkZI2P/E9eRx9ycHOVpwE8U6lZ+RcZ7DT
z7nZN3H8dvDJ5MxeO8FbY9lMOj+OZ/MV/7g4H6V4unfVUpdss5GSY9ZpeiVjs2wI
4ECSVmekrMmXsPIgujVk1huMKHDRI9l8HO94fJjVJP53Pw5QuDrZGIKjO7q3s26V
f5L5y4GAJ2S9V04B7XAEkftKOKP/e53lrQGri9ZVInM2HyWDDJydsGigaSYmN4CU
cKK48chlWB7vA9A1YWeM/uQ0SHp5AGV48FpT0eoBlhlqwpFk1wRZj4ojiKticJca
B+KVGpymxqFXJG1hyDgv7wN7HQNN8cS6fIrk2ulROhmrgDkIFmqEcw6A2dXkxiuj
Y6kc3c8p8D3UkAPiqq61A/C8mfL37k0RxtLvD99XUNIDl2g7lYk8bCicB4O2AZGv
5iwsVJxfdMBex5hp/6P+o8PFwCORRj9jvb2xXHe5ZRtiFMFHNOd7pz/WMu0B6mM4
Dk5niEYOZrmd1Jb6mTLEMYgByKDIcFfxpJqcL6kCZ6IN5bEbF1AcTto0quCsoNfI
mFFnScdpMBdSenkYhIWAX8n7nCm9jZuni5gzbD82Lf6O6wu7JA14/vJPiwzdThTX
Gi9mITmY2+WgmxIXcjBtXqY/Ze8ST14jwWXrH+lGg4exM3bLJPDFVoCGl9VxZgvP
YQHsx3c0JA9STzPF9NbkvxeAP+pL38O57OQkiIT9c2+I+P7XK7UAhj5OSDRfYb1V
QbBlp5BTEeV54G3VGeVcXSb0oX4rFLxPNU6qDbOYmzQUbgELZ+u5CJrRwz2Rlfda
78SoG2bg0oV/neeAiei4I9KF+Hy/RfdMv3fHGYyDOiZleUvjuq6uzlILurOigvLj
BBZ99cuTc+27COPmisWi5DxIq2yzRBN8bHZWSi0ySQ/5VR0U5nrESFbkV8oi0lsI
3T99WSvi9tynyIcS0VQJHDa5beNCYnx51E+HrozQCcvft32wZJoKGiC15KpH/aFk
glwnldTVjkIOrvtc0ALqPuXRKxJKyptY8YSXJbc/JbiOid3q85yDqqCGBhcq0Ccd
VFOKYIwbJp4GATu5sMPdgz30wQ8hG482BAeNQPqItyYlZgMekGIlJBQ+ONIqtQ75
Hm+cQQaDERYyYJyZoeefwb8wVfdZmI3Bb577vZnJnkxrMDVVrekVRif2c56Wo94g
+bw6+lQ7w4KTV6kHQCORBi96hKJkI/pGB2d/NbIaZCsxOv1nqVwe9KkRaqLpUMMz
NawioBa1sUQoprwzSKFQkks88b1cj9ke+ONGp8EJ7YqbHl/Mxz+cGV+5XCohYkBn
5DOfy7LBngKEziNTzTEqfNfworhZqG9Bmd5/uvVkGg8dFdJSlP49sIRc9B/XSQ2e
HswG4MG+o18d9CzbSEzryQaFZRLqI6QIfyMcdESg3upQx3xxtmfxwI9eB9HqnrkO
OGfhHvdVdt1u0/gbPSobxsg5oBvbNuRl5rLxeS51CmAUPa0I93+xZQDK5Mrfrr/R
yO+eKMht1/MqnQPfe8u9fdwG7WTWwooW7V/QxLG886zqkbT6PmP/66FRQUxwDLy3
7wQP27VhwpaUqjslc4ozHr8+zJaTQC5+m5X1C42GWHeQNO8r35BnQa2h6aErSWuq
x3r03iTaxyjpg8TBYQXfsIwtJ/SZyMWeJARxh5heaY++in0n0v/ZMVvnVeuVd4hp
bJGVchZbkUFbmBp0CJSDPZaPlbGHsC8ACf3z6zB/yX/oNb+G6k/lY/8TGKzpmGP1
AmUWGuZ6nVcj/Q7DZ/RXpV6ryNLpSIcufG6O9Bi2Tfqw6UVoJBlFxDZT58f8RM0z
9/6d9dSUx41akudabY9v2voij9Dk050jfzLSkSEKGW5cEMOKU80iSLyGuY9CIdsn
9GVAKKt9Kn/v7BZfEAjkdQ8JbidZmtGruce87+E26xvNubtWRoyrlElpO46Jr3uX
0mNeWkeS4Ff3NNfmi6tmL/4Pf7KtyBrE5Zx2wNNMSwJQC8sTLg3AsikiVplgZgrD
PEV0SZCsUUstqV5w4xbG4SQrssYppu25HrmJQ1gRXsEH8UGadO/DJXUOOW+CAOzI
pUo/I5sGWORfeMmJZZC7CjV2Tzk6sced+ZJYnclcWZPFt+hprH5QcOeMx+0Wzu1t
Rzh/jbkZSSwKz/aiWSbVGgvPMLMHOj2I+EvR1M3rvXKawb3R4IUos015pQMP6DP0
BPpjIj4XiouJhRtjZ0xmD9M9IkdCBaerc2wWmE1jBRBberPTxr+igjpKUgfxWFea
c0m/+Fx3FQVUdZe0qxWvMOXnLMjXozDDaN4OxZMV5BNTZ8diJukfgr1Gc1DSilVt
8cLcJmLcE2BJS27rUr1ry+Y9YlkvKj7Aqs7goYZVIsRPnsnXaXs4x2igyxtItahl
lrZd0561b8ykLlXzztodPY/nauRiWS1wCdjtEfJB81q2Xku5mfWx/ss40PSWb4fs
YCG5sKzlkUhnraDbvYHye+R8wpg0xkBNqyE7bNQL90yKlQBEV5wNeNeRUz5U005q
5uydO8SAyloWtbonu9FVXzmUW/C7ejrnW+GYd4yH5I81zzhZyLchKfq20gQoSkYq
Lpa/Oa85qm+VyFZGqtNQ5w0UvGKnrijRe2uzv5CThmnzhPdykWLicrKDu8Fgo9iT
x01i+Kfah9pu0/UBc9T0SOwvPveBvYXTMotJCl7plXqrG7BRhDXcFklstsXxymd1
/y3w45yldmciHa2h7Tnhnt3Ek214IYOIElHRUsPqPamxtxNdOn3xQN0/utbKtJUZ
ap0HxM9MjrS4V1aFp1fNUeEgSWvn0y5ML4cJasZtLx06wNFIYZ2O5E5isKzIPxGM
XBHGjzo82AoML306kiy0Q9zZga5M87pGn0y61ZXnnxx1n29B4hOjSP5li0IS8FsE
WEVoF9mHXYbSgjTIEneZckY5F3aBDAUVKaOFB7zcOwH1KVz1XzPJL3xJaoKHJWc9
X+LiPDFeUWYIJL+eGCG2FtY3ATX+3TCAQ3nbihDi06418Lx2Az1K0WJytw8m3xbB
CPNRErzrZXapSJ7C52DuosYiYINO9Yp26bE1nJnVgcFA7xzyAnRoL7EXVJnJ0YDP
qVAqY+wMK9pt0AcwkDDEY7OIGIc5JttbkxBVylfaAIHc3T+k/FNmyW4HrGV7Cys3
a5cVk/oAPQrk++oFD8KF6Z/CXhMSVuDw26L2LBpQqf8hhJJiR4QmPgr6DTEFmxj6
ck31zUqT+rwkW8pA05uT9Wx8a4vfHGBTZacV6j+eI0o6eYvCFbihV0USNT7BdilI
jqbgOeIxVNyhngQrMZ1UPX9xQdAK20zGdiTTxoSSsNcZFPXFv5FgCIARLYcGhoWh
FfDOhbMVCwE44CLJnNTwZ30jiBZYp2NZmdTDgTXb+bGjmki0oXd3SC+B3FNXKpY+
Yc4CjiWgOqFIm3cPwh6NHFucC2xK62VwHyJSPJekA8Ue+9oJkvhNarikZ/5aRHp5
ldOrVSQk6uzeI1rPcAZZOsrRkdA0M9Ynpvq1hKabQ4WLH9Ffsjp0uKfUC6cUlyAv
V/mLcFxLjVPe4PhPDaIsTA/WsfdIrlvExO/5hOJV65qIlAX+ljqa9XJzku/zDF6o
UUjYfRLMvIFqMTNpmIEwaasMC9L3BAk93TxZAOYdX3RVSV9LPnIklRB2v0ALIAR2
mPRvFfy/n/nUoCu+lEaNAc0XvwrpqksY5UnIAY8R9m9nz4yHs4wTvwxeqQ0Slhx3
3BZI0WWPHEhehPKABuXf1tJ8GqGIaPVHVio4Uj7NIZimjMPwhYh5Gt27LlI9/o9T
IddYERAk4D8v79AGgFm21Q==
`protect END_PROTECTED
