`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cORKG7WyOrN0JIc2t9geHxKc2BpBO8xWEXeDMHJ2XegcaVfCDl4OnOb07y4dHxOO
WiLyK2LFCs9PsdIhQnCPd6/XxNJQK94aZUGcOS+zPgk7axyrA9kYqQfsm/vYc+eI
YY13npkd1NuchQ3+eXXmkAt1Z2rQHHu04VPqzRNbk+AS83uEaHzqdN+E5FQ015aV
Hq5uAtvP8L8ID/8AfrQyf28iW71RPKH4/uxNlkuMYl+RYc+3vBzO9GLPkRqoa4SX
RCvWT7M81WEl8Fp6yfuZUVQcaZnbktR4OKinDxq/2od8So0AhtOAlE4xguTnwBRS
2vo+2aSUId/ecGC/oCrQ04KpirBmF5cmvTsCY7QHF2n6G7qNI+zcUri3dpoIX+oS
wp/JDrVi9TczX1XCnTYmDjaLtJ2fbow08fV6rseEV1KIYXCGtPZsMmEWZ1p0cfqI
+RlVL6/FGqMD4v5vNqo6XfrP+PpEFIMlm/wk8R22VVo7+wH3l5j+jv1rnISrBi1U
`protect END_PROTECTED
