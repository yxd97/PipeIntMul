`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rClLLB9vnzP/rRdzqJcfj0lUHihunwKN575H77hDApg6IYb7boKrsBMJvH8rgauW
iZaXnuqrORNJ/CedjiUCr826RAiv/EinnSefg3wQkQlo/cyudG/bnz5oGb5Ld2X8
sw5cGEybDM3grd5L+rYzYxYXILza7O8kKzJzyXEuP+0uzDqcSDQEkAGB65iYwwuG
KOJAnzysBzgKxFck05mLp6hJ0VUh8OqW3Iwpb9A1brA7110BysxzcL1rwtI7qXvt
DklJsarhXzeudb1Q/b7zrxufb64eP0u8BugHL4tXB+gT6I2WM9ziZDugpFOV22Mp
3u1l8bH6BNdCafQhTrFdI9+KEqiEPTPKaUdcZDPytC3S2a7QpsbgDVKdjvrZYTh7
ruBDUQ6xx5Ay5LXojDqlpROqpbJixMeRPqP+8URWI7TbbudESs+hmToVnhch5CQj
EY3bFv1uns/8IItJYX1uHqttWaLE1C4jCLXqqhgkV/47z0SF3rj4/fZVgZdbGjYI
hS4X8G1nqmeRUJevxYo7LszdPYreWmkvr5zy4CWfvh6n/TZcZMzUxkXvn4a7JNbJ
PihnAYiS86Z8LsFZD43mXG4FqM0snJBp63mrmZva/lvhTBWuJD5w0b+sqS2CLM3L
aXluJ8unKeXTnL3H+2u9h94+95xALm2TvfQGzRM0eVFOyadZf94fKADLG0LkWZFq
eqZDrttapaNVppVwICl4MSIVq/y7rZeAFyh3fEXbZXqkujFaKT1JJDB1LbMXD5zT
SbY+MZmDNAz+TMbkliGQTjFDqz3YEcX1B7orkRnXVv0l2D6NRT2rAapQfxCIYqKW
T4fkOEBaBnXa7G3rQKW6IiqgTB+FWeFz/zf/FyK7GMFJCCCQcHIZ4C7PWxurPxL9
TO522SdmUbsp1M/1BwGOZMrKzHMO9IAzjxZgRCfhNmeEa5qMW+Ia/GgpVXwHZW1u
5P35Rd3TZz07w2EKFA8jfJMjC5cVyswvZFm2zBhCL2AHznoHF1UprX+zn6p+7EFu
dEcP0gaOjueTqs0b8iZhHg==
`protect END_PROTECTED
