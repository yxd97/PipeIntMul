`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSbe3dBcZfeF9CnDvSfh4ExY2QFv1WYWYLvbdXtCgzWMa+wsHKcCswacqCwQ0LQV
oo0LK8p2l5IlaGJfCQPlZuwDCxtvNa2XK/7pIEkP98SAV/NVut7pBPOL603BqHRD
F8jjFNMVsmmP1pszgb5K7/lFhup0OYWXftfQxwHk39CYojyZOAG7+03UDaUJDJfy
77TovBC//j23XnJvGhoSL8bggFDofHrvuan54K1HcMyVnIHPr8WyNcoa3jQMDe0c
8J4QjqlZbsxNtDiaY83KIAvle0ODtIla924Yey/QzxarO/bhky4IS4j38Q9IimtO
LXza4dno+W2bMO//aJjXAw==
`protect END_PROTECTED
