`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJKPrmpgJktj2OttftPcxbIU7xXfrRJXTZDcrCyhwl+0R40OHBDPZLV2h2Ucc32s
P2S+koe5mDj+L4WHeFm92KxCaYkFnu5QgawcCIChHAi5JI8K/UqfWIU/TeyCWk1v
+ihMS5TuYgLWsCv6PSKPM0J/v4f+RQSsRd3S9R6KELsGn1TLdxtxDzrL89mUzbS6
t6AuBVj/BeE1xwNl6FuIkwbm90dRxgIms2y+TFar67MlLkZUD0sn2yu3isegP0Lr
r/J6FYtGun+ry9o4B0pyVXMcVCIztQq/LISzBTZBS3dTbdq76+ts71KCnaSra6pl
2fPzMPowR3NAX5TqpbO7R7pbIaGqM7FaySkxrCh4LFBYkXi2Kq2+iiz2rjFpzY1e
`protect END_PROTECTED
