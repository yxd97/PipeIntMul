`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5wQWaIH0CLVMNAa5pifgsoZXYGdYB+wHlwCwG+SAuFq6VD2mfXvbgWDt8LpxRm8O
ipVNkhFVxQapzRk497Yt6KXEW2Segn7SFiuPN5bk/rjS6bTGKyL7OQjLgx+TuNJo
aByELueMEB3LJwNmgnobiHpB54A6GEn1X9o8gr77paPpCh8qp5wZfaS+0ARy8p2B
8W3oyGkx6K03V/YYkvlTPi69ji81A9kENqnVa3vZbKuF5Ea0J77UBGdp1izwQ8PC
fLkUx5fx85EOuCDG0MFeCsJb9fK67PlTrLAwY7kR3DuKZmdGPfkUiElVlWEBhPZI
gRKC+y6sguxK8vX3wGAFgs6HJ/R3wA35GBS476A3UprU916hBlwv4S6NLQj/bnow
VzldC1lNUE0SStMy9ecy4VxcbIhBFzPuFHj6oYTuJDg=
`protect END_PROTECTED
