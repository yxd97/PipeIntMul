`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AsZHISpsK5euv23sCM1XYOGUNZcqNiuBNA0f9Zpts8H9Wr/Ht2pcZue0Pja8qIHw
eZtI94/TB3Rlbw/lE3TQsFA8aLTvU20JmFphCzsUrEaBgSx9i+nM5FNh8ypzz+kO
ElCFgJqnYbHaqXRKVQiczRMAWD3oPjut2mPCq/oTz8rEHv62d10INgKxC9ssC4yQ
VGVdUZFNqAyA2jUTBJPlK0ev+G3ungUU2M9JHi4ndX7rPCaKJ7TN2va6mWCXsoE8
DaiBb/xhY4UTlnzNXAXHhRv9v1aq0ltMKrAVIxwjXQRoHOz4QQBHRg8nouqZlfTf
5SUpTJfDmsZ8hJs5VrAATY51gh4C5mygqCgqSuxQNum2ZjrL/fCBi1H2KLg8XYqb
pJ8HA/4IpUrFT2YeqmuOUfrnN23aOliU7bKx+AzpTNw=
`protect END_PROTECTED
