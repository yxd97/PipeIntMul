`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifxJEay/3BIZY7a1uQR2QOu4U6+YyqzJdKTc6D8bfOI1+gYFGrzAMzEWgOe/wywn
Qv7YiI+MxaULBhLwfY+jHYkkSsHtc8495bS7ONqI+xm6tWU7AhBGVw+1j0hqklxo
13zecLatWImAgsKqzVqxDjTy60CmM9Ha+XS6uhDhW1M3ArklmgVLlmSqC91QgbA8
yQBmJHnKpiSD8RBBHvUICfhqSsYfgs8AHT1BN9B/J+yIu4gE3A+um8CoO4VlXbg8
gM3JdZpV1WEh3vtydJ1k+vt47QbTr1I38SlHuDKpfPNql7Oy1eMunMLNPhdLSKxg
Kl1to+oPUA1sJ1Nv9k7kfAxaj26bykcZkP6BlpfLD9RjapE529XYvPgsoR6EHWg8
N39NC6Voaw+sWV467KULDPqA65090rQ2T22aJL6Uzzk1gh1e8SxXDEKeYTP/DzSs
ur4NwFH71EvR7+K8bB7miLvlzt2tUYmDrlxV6MVWpVPeHC96uKlcJDLQx2iUQ+HV
Zt83mI29N8NHelijBTEq4IgUA1fOlZjwcbXXkFylurH8ga/cCTrTyS5orAE1U/ea
PIwNgEEyyeBW1KEPWwHspJiXV+ONJD2pbTo0QPNah5QEIj0/leKV7Y0Sq2CG5Q7H
DH2srBoyRFFpMP59smjdLg==
`protect END_PROTECTED
