`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlFAJWTYhvHmjFg7PH0x4Egi0sSMcKcy2o7WOwTFK5bzL85fVZRYMqAeLzJC3tU7
pJeKtSIH5Q0Xa9w855HTB9eC0fMjp2Fok3LGTzdHSdOkkhbdl2QCv6IGiY9pEVZL
OxjDHjVOgd+GM8cdYWLcB6qv9b2mfEHNCvQYSeENzH2rP8gy/Sx1XH/nhJJT/RLY
2/8+c3T3cOqGTLkN/r9/TgAgcplNsFvB70Cw7Ggz4sGDp4RqWT0CO7NF7+M9T7L1
QOOzI4IbKS6V8CQLxL0HuBp9xYkHwd8Pn1LGsvOBS2luaIyb8xSNekMtE093fLgo
LB5TXgpajX9vYLVf8T7YK78U7rWV7vENoRKByLMpuJ5kpZazFohZwyNv1nm94zBP
5+2LZxAYY14AgQiDh2k0BPZr+PjlLaS5U/2lmrr1xaPHVXs7JA/o36EiE3Rh63CI
tG1UHaXxC62wGCf2zMfZan13bdnvdNTyS6WnCNvDKS/Eo5wfk0N6wKKw0wxqUzvl
5ZIRLhamsPB2Kf+Q+rEH8nuoO31vNdxhUyIC+KkgCCMX4KFVSG7p7nc3aYYg0Bn8
KAhMo5XT5mbpMGDxZ3sh+Ir7T2VNrL+v/QoyJSXZEVK5jqPV6UXWK+NFozGxrVVU
JAZuGcNC83QZtWnVQmFefxzdJ43HLbP2Oy5bUm4zqs/hXyLRzFXJ8APihrlDSebl
E3lm8Ee7nlxKDwcGbtDtsyA4Kh4im0+2LBZnHTkUZb2ITlFolsaZE7g7GwoA0/YA
/9Dx4cWWBPmwNj88VcWkG6LVJzO79AEE4PvEwOGGgM/kfdV/i8zvEbdwhSFDf+U5
xCGCD68nn3DPzkkfAIlroTo1I2toA/ENUG7SLLn90CeMXXd0JFxRpNpA9XqQCMxg
8z6cGst4V9mqw87mwn3qUD6T+VpEJTlU/orgN9gd5ytaHoVry7ontMx5mo/aXy07
YraMaYp1Xi4+vpgctOwLLQVP6u8w7qwSaZhVEtXPceLHx9ALCKhMpkRI++2It2rb
iM1Tf4X/d8TpyWYm/ALVX+EU64JsJBrutn+4uM/melDWBjMFNv4Ry1hmZIAiBFZC
toZRrPrBY6pheLiJQc28KZl+3gmyTF9QLqO1KE1LPBZ6yyWtptOrxldiqMVQyrci
CmJVK3lW2I1puLHU513ws/Rj5kCl40tu/8770/2xqPCH+QrydXc+mULQl5NfJfQo
V5SNzYB/Ru9UoM0SV6QPVm1QGF9IsmrsFTivFqfXBMqcVJR0BgBkd3EqPAxWaora
Syz44/EAa5oGVbEuw4ctbeDoJx8kgY4VY8u8tqumpZsD800QGeUnN5TJKWaUObuq
udEOWheZBJqaoTOd0QBj16X+tPni/LJYgs9Slea8HybKj5DTACvlxahGSvC5XqEX
`protect END_PROTECTED
