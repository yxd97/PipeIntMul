`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dH9zAlTKzVJNMe7m4Yym+A3xlrKVVIihJ1FiHlNYv4ATCkf4U+s4uSmqmB78T12g
JWs84Hej+KA/CPXsrVUCj1yGPMNG6/yBYbcidfr3I3Xm5PvL42sCZ9qnd71O9Nm9
wazGvuMBGWzuOdcARB85f9KjKwfLzN1JsB6J5DCNSxg1EuqxZvUL1ys3cZu7GkJJ
UBSjkl+eb6jktnPHlaQkpkEFIXzNLRd01mSQqtcFjwdi/B2KOj/d3TtNkIt5Uf7P
I6lUmcHlL8jae37IEen4lrZ8vciq/xY7dXrBvb0awa3uKj7Ex32K/2jdBXls27yp
9FK/Yu7Ff8jFvhVU1aSRfQ==
`protect END_PROTECTED
