`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fzx7lVdnXJ+iUwg+LvUW9g95Kaw0FcQKBiQL6gKLRjkLmNaqiR9JTE0vIFB2kLrn
xCn7ov5hrJEE3R98ovax7UAB69LDSBw4mo3s080lXLQG4OnzSfgByQbn9e3Ut/Ak
4aLsO6cAdajnDU+geXfCcZvqVeMczgVgVgrr7LUKGkLlNZPiziKuCzceGiqooJ+L
lb9RV8QR1ynH2dbcTkOFQv8A+jrozrHNLE1bG7+lgnQzRIz0immrV2AetdnVT29F
ONHDIJzoYfmTymPG3XH8vu8OPA5I0H6oqNFRXIgBHXS2+z/ADt6u2Fi3BmuX7yp5
BdCVIiuFrvhddEVCg7X1z9+x4kgiEO+QGPFDSGDRun6WC/T3D8O/2231kFC4AwMm
E+05RB/JOZknUCu0JorLxP23jwgA2g9A9ITfsirKE7ig/Vrj2IjO934MDMaQ/iGb
wvQgZScX3S/SVwxL/LIJ1VB17OWB2EhFHja/20MO/0obF2ZsmevZrLjbxEvgDzLU
L9rRQ2qFiD4TCJfXedRWwXib8J6hOyKSF9RV4oDa0L6MKwzrj9UaTH0q4vPh2pHi
`protect END_PROTECTED
