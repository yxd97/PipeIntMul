`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0jz8NC0ebNTPyQqA76nARocrfQI8peKzK/ehVajT7g7x+WP/wFrPqAk7HIxFyK2
ixhOYK+02BN7Py3bAoE73KzDIdKYYW4hc9wRNk8J97ypZg/UTOa7HtYYU+P479D0
AJ1UMGoRHwCGF0zXizgF7ZJCTlwsLxVlbzoJVOyfkb6Dc0tuVKvsD4fiVFecO5ts
Noav45GwCatXD1n/woWPJOVBwGjEIgxSOOPie3ziIh+5WHn9Z3T82reIMakw0i8W
u65XJhrPT7ucM5D1aY9RXi6TuXtaDxkfyS65N4R6MyL4ZPHI27WjQELcqN6ntKMo
cQ9HC16U0wdl0601dAZTlwJNl+zxbYUZAUqTRjRdiFmBlTSn6msZTKPD+/gC6wzp
F6yognaCadQydBJOjmjl8FC3JVGssoLej0zcpNOO8hBBLuOUPFEqJeKRA/6fiSMv
jniKzHlxVztfp+NZvjcnWz3qh1Xmkq1HjMWbSI/0Ib0dvfe4bO+4eBqPUoButUfT
wHmatueYGyffOH5yAJJzYp0Y5kxkXmLM2G9WnXjnOIeht0LkpWqbM73Cz33MWpFe
hzLu61Zv+DNcLJyP5VkX+mmkP1t+Ke+S6vvP2Pb5rIOwXlCmOkDeD1v+NdhtXPKt
pYatyqOHrabcmDJm/AmLOID62esBxzX1VqjAw4suoUI+n+rE9/zFMt4ef68u1mO/
GlA1JrHkuAtuvUXebVCI1uWCFuQXDuZXQjtO0l6sclQ3RUB89D6ddR46fAJoqHwx
4tbIjltbllVPxiN6bKldDkv2Vbc5QCIY17h0eM55YFcbs6x46NjkVuniZSVpZGKg
PtAG3h22o2HO4aeuXurdAz1ChjynS0gZi9Nb2ZLpznTc2Woj5IBL0BdgAJonUfaw
xG9rbwiJxrmEhxqNdwzJ+Dgn8HFZLDeyZddfGVQTOMrWBpb0E7hHJB9YMcwekc9/
Fg3GjdS/JradaTaNv05x9i/xDZv4A62UbOrpCES+KwNHFxJ6n4xxMpJxGPI6jkKe
TaxIZyRaSlHnX/R+8sAq5tIVXgLUWuBgEmItuHqdowrMcQvBniXfMut5C2MUzI/O
VCeTf3+wf7PeKEjaeF1TrRo6Yn92TQaglukuWXz6UaflMvNiIVuQeimENa2Lb7Td
BIVA26T6DiXMyCgpJzNfYVRocgaXncPl+zSb1uEHOBvB6+cOfGSpuzo1+9q6Kds1
L0yCurboUp1LZwBvGjoQY6/HYua19tkAvM8d64aMjP4/xnctovBOAdZwNt8+HWGD
TQEl+V+2/ajtDIpKjaU9nWd0jzgbKlVLGaiXwgmwJAV1Csuil0FHGjdKMwTkRRZG
AeJHQCNufdp+w3txsgoMVt6neeK7DNJBQ1XUIW3NbTGR91djaBuQuIgvfpGsri/A
75XAWPxoikTSf/2dQ8SPjz64nBSh0ezAEoH16ZO8VxwiQWhD3lDQO6aSqTeQyUsa
MDrqTqXPmk3ETDkazkIc16TpgfHNBkYVXR30v7tZl5/EFP+aeV0dEjs/vQDF4xVK
MsanneVDqhVFcKUrHUaHDbWzTa+hVc2puiWhdMPDoTIFFUQZive7CvQUxWmn6iHp
T8UEyZSjbtNG2z3KKQ3szmAZ5qIajWK/Ff6CIIhFNhEd0Lu1GKy94xgWbnZvjOfz
nhNIs7XImDs4CN7V8ghCahJzpaPLCEsuuLRIhn7aaPmBMp4z2IesGe36f11AHq6p
8hTlL132FGDb1i/IhVomluQd9QsMvNkCwazr3nwybNXk1Wp3bfQmwcMECs3XJ99z
S2vl+gpAeFrz25zg58wloMcJK3HmpARmrKOxeJcfoJwfBkvDP/H4z26Otk0LRPBW
atyNWEj6yXGDuTblW8jJUNm7n9Zc9imAIBR7SMZYuSqR21FCixoDLCLEt8/Esb0F
u0/qJ9jptgWBJ7SAz36fS5LjbhmN77H6oR5E3CI6wEBWJVjwN9LRbVVl3Vk1Fqf1
/EUcYZNZLXDOmmp3wsDnpAOLjdSmyYZ2bvonPLWguuFFc9+6QVqBeEM2VO6jvL0R
rAxHxc9v7N3t2y2Xi7MjTvJmOF5DyTWalfg9L51D0BODngUmUYOYdMoMBdMX2J16
qHkSIThwCIpdEdfo1G1TJT0CYeC1ePigzvWZ14mGx8gurWED22BZ/psNBKbvOd/S
buPv2PTGVbETA9d1oDIQYS6eqBzGyhITabY4sNFRx0pvG+icgSzu0RpKrNrfblm6
XK64l529394rVFrWa8WJRa3wWJ2BeJOJUczhVJ8uM7WSOfTgp9xrJJ2dEs7D1B5S
oV9oCqEy+FBp2h/foSHUgW2wq1UBsYqPCs5uk1m8Q8+TxyBV/9PQfMU2M7rpD/op
9V34bHXRq0s/Ejtf9vVjazgg2FOb/VmrSVZ6O+W6SzXymPr6Nmmj+mqAqyNuHK2D
xhaMg0YUARATqA9ZHW6ZE45KR+fJM7ojm+yqB/wJ+AJr1RhGCguDTF7wcZy24i1s
VyWwXkdULsmLIA8GjQ8Srj+4ADrb3mdRkTBSPhksZN/9FgJ5ARr8XpRpc8kFr4ej
JD71HwBCEb/6weVjs+EJsyp8r0+5mE57fg4X76b3+IlOryOj1CwDPeZ86WnBqLAm
+dC0k1v8eEfkxFMwqBlHNtpftcUy2CfVPNqq6qXSKCUY/zWjbQjoFAstrdltO0KB
BWe7WZZ6j/hrBcNUmOOXfvBHTzIDhwQ+HjWfCMC7/Mss23z/6OXHpEHVN1VSWoDj
TK49RzpS8mwllZy0i3UX7CMf5AalY21tgLmFcgG24A1JNZrWANsvBPSpZXgO1GhB
bRHi3+zoCJeZYKtpPypPGehRwEOF9iB0n7DkMOpVBDDKEIitoYR/QAKTKD/RGmck
ui4H1aJtqxt6DHWTAnggVzLzqvmdJ3bVAQQb/l2s28IqkcPbht2+DB0wMFt6rEoc
8wmtgb/Bp0bVlgN9tspuojLlFking7MTvnNZ0oMjWJnxrDduZrI7zozG/b4wfP/S
Y9OZFoTfS1Ue9tjybbns5ZmKapS8zWsFTs8StXvgnLc83y6yxMxAGcusLOvI964U
TrPLFt5CfiNDqBbX9GxSpMEqEm5oKrBiedvfrZMXGuXSLcKz6sdsfd5PRcIjMige
G/eCGewn/LO7INnG7CXRGPY2+zRWBBXIgZrHlIC6JzOmFDNafT72mQBQMc4GraA+
e/lE0R/kXdnqdPCerhEkr/HYS13fI7mx75uVhrfYmGx/MrUQ8KL20fbpUisPkBBS
qny46XxLTLlvPXvqSrD92oDAfBYCpDCE4NkTEOw1jykWnz6CPXhJPAsPsDPSdA1k
o6Q/Us5yrj5BMX5wUkj0fde8GzXSq34BW/uKS74B1+PqaGRQQv44i0LiXcfji3w9
id8O487x2aEZmFjagN1P7V51rimCWRlGadw4rxgt+cC8OhprVxzgr1w3ky91QD4o
gt49ECoNJs3SKxIAJX+6ppybQr8V0Mh8MLGcXUAcp54dlxhsfquDubi274bhr77f
lwfu9dT9DQe71kBpohEB9wk/rTHppyT5YufF2Lt1jidUKYys9SEu1FwBu4jDArvB
RNijYSSsHN70CYHODzDYpc8es7q/bcS6eunWgSzCs6I7/YQSkN2QYIx76lA7IprA
2jc2zOTT9ZExkcTFlnSrNygvmP9dWu1ry/3QVise/ht8ZRVzyObDWsNEqNEKsN6k
A6DSPxJC6sa76ugNAw5PSVsfqWS84TM8W0hOqeGcQE6oNI9ymt/zngXigSnCMx/2
l1PjWCZAog3tTyQ5FveNLw0tT+fEMr9DSh83pyCgt5GaxT1HWxyCkv1oMnDhgJZU
7SGOkzIjyatbSwxyC0mgAZQ/kmUW8ye7WLOU1WwQZCcNw3JzMZasR/fobF9jQOJv
fGVx+JT/83XVBYVaUUDxnDYBRvYu5nU3gqS0ZLO4k8F/tin3c8+ThXJrcGqxbLUH
ZCR37aEsKpboT6bq/wcYcOXVxvEeNUE2iYs4Y/ZcKA27R57YWVMp0v6A0DsBjy15
D/uhEuZ3+TbezDZoHzH8/620p1a9bcq0pxY4hs56MAkRGk/J0gPGraZxHLchii9p
atWVtfmGtdMnafdcq2lvmccvVM6SI7dQCygvrzswjFQMncYKUoQLZzhgz7ZVtf0c
A8d4mlENr91IOouNgGwHDvWUjESJt1rXTeWgAZYja7tgXFrZcj96jH8TIGJZsf2D
47gq7KfhhgpUQX7chR8dLxOh8mACdstIRcVCwFgEoqqN9NLxm1CvYDGi7cVcIxyG
wo4LMrWyjXVH10DIb4fG0yewt7T+q9eTRbt1vflrm+E=
`protect END_PROTECTED
