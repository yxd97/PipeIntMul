`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ei2k+37lzlPgleAuK9Zev+qYoC71zyDgCuIJ8iRF7APNaoO7GJgA+M2AAkuGUJmo
GfAUTInIY8cDmZ5TY7yZGfveD1P5F9I9Xw82K8r3DCDgKr5+sMyivMXwX7evPvJD
uocQkBnzdcxQnJhHhbPlcIMmVG+nITI+DnlJ88+qJSoC1ZzWxeP0DY5PhTk+pGMd
2VvK7fAe/MeMilltdZR+f8yrjfs7lLWNUJq3rJ+tCeeI1NW8Lja2ivOK57kQtVxX
TJJNzlebiXWRGHemWDUMKMmM0ZW/8+9+Hp79Na3yNm+oovF5+MMDd/sxw6LWUCPQ
VEQOwbTLTVYK183emH49f8G2NI+qAMUzAheT3swVu9Nc3R55KkGkvboYF5d+1qi1
3Kf7BjOYROPZse4s/niWeevReamnIVaXgbGyP4pndM5XWDx3xjWaT28NwPFNuzkf
OdnVL1/jao0vawhM5mlOZzbn/ailAfsC4U/oTQ1Elp2Mxc6Kbc69xBNAzSowDf6N
Blhb6rezvU2JqBwKC49/2yt50xX4gHJztU5FsZokFooAgbbqDdrOC6miIJEID70/
1Jhoo6EZakt3KQXJFYhQK/kBjWQMDWHMZILytiN63NY4Zbe2xbRUoVC/zWho4aPr
UhVPqVAsjERB6UouzcKVJ3TCfcwxUD3wbKi9iZKcIDcbmnxDaxLfcZS6f31/slAg
iP3QT9SxHNCNS1atN8lWf4F5kvNJ3HlGzFzthbfZAXEZbOjgaqEoCMoyuy9G/W4r
tZIJpi4MISH/tIenG/5rgmye/v16OxUryUB3CYtySHYxtumCuQ49GFsj1mpFOUeH
4EdkKwdpzOSOEHdSOCScVRt+MmPSfoGpf4BVgMPdr1jbsEeh9cazeagDRc1hNzL0
OmSJTpN///3ZF2cuwh1JBzyMluqs0v4nnHWU5NUpvB1RjOJoPp27JaY7EmSf4hYR
e1aT89q4NxlF+t3EqRHukyx6Ok0dg4IAhhnAy1jzihsffI1HssEfsZNej2UpsTkK
/GuyM2B5SMgfqv7XqXwkls8v9s2fxUljRR/WKhlaQ/NGW8Z0xD/a84zXK5HP0vjD
QDO9xvXTs1U7w9xUmkfOxKG4/4hg4yrAfwIsfYrrL9700q6xfkTJ+a9yCLf+hWGy
9eyZWXsGf+NT4A+8dhOQ4PSpDDUPgQdAPWDrxYyLFM5cGTSrJj2+Bn0VFIOsynwg
SzxCSQDdf2NMD5+IBro1ybVv3scCtd/HrTXBBLY9A2TiKRZ0Bx9qa2a8gJ05zXH3
GCWVY4had/b7FYZzNX0qxrBjEWJz4RWwaJNyXzIIrWNPnjtfjSM1OGeR86RjUbxO
AMKZSdyt2U4gFqQez9TjY8k3ShsJiJ0zhHr0vtVu3Tix9dwaez/TnJEY3b7D9ZLI
2xjm/PV0U2MZLyD42JxRlJfTgc3/DZk5hmHXrUIJEVEJ8gR5pQQnr017g+07SEQx
DRYL7ofkjwJ2Lo2034kHwIyrgGdxgvRMtNj2pjg9pEU504x0AKEKBQjngCWIz3d1
7D5J/AwapX90o0AkwxK9p1wJRUcnCxoKeOKCQqlhtbUQroGl7NCmEfL8fE7enLUk
QbkmEg78XtFOkWyzFlz2r7u5NQZTGxvXEcKYWNUBlOGp4/hhBmmKjt3k7MmalTY2
a1Q6hOHm5fFaq0O7E2bEl1Q4iv68iNfVQ/uBrqPEJnpGx0z+/7uiEVjwRkccJBcs
iqcjfXeWJ05lqhI3l4c/phFdPisRnYpNk/GVgCEP6Q2rbZkd1p62HG278R9aoqdB
yLTPW7WGtasYfTKZvFJf/FdpF0Q9yHxg6gwlu2KdXHz+URdU0/JQb3waflFfmhbx
IgKBz4p0GV/hQCYw0IAh+/ApVUWcjVorPHKk+k6qjL96Kb6jHYct6A8xG+w3XxV9
n0v2HWtZKzh2EyTqZ7q0khlJrADudwE7Zd9bX2yS/CIJPQWr+CASjp1hLKK4gTuc
b0WBQEVg7jGTZluLmuoJM+kjhYwF5uRr266vIuiSfzRj4C+P/4sGGseOt3mZdGtJ
mNJFCiHAgl3X/8YVxv/yY3Etd3VjspZ9qZNtbJNclf3mObM9555Y7UKRGsMHreBN
LmyTUrOk69U+ywS7Q5Urn4NzD/JsY+YInkMrGRAv0yKIBzWtliwIgq/O1KhKTl22
ADW9+ZPigdy3nz0rqRZxm9GovGjNz+Bk0G9dIhjmww8esQiY26Y8s2/d+avVSTyj
RvxCBwwLXpNK5Ay3B9EGXoI7z4wFSybD2S5AYzW0Ob8dIjdGAsCJ5hpr2E+YtJtY
lqDgXIHkaMeJXmuUh+o1CACHw7UytwMtTgrbaOsIQzQvfDOEipWSyrvp3eOuMy9B
IkTKGWAEgjJjF0Sjsbg9cvZdkiudSRYXsQJTbdO1Y7/xkRPJu8lBud7jvPW32tnh
cnOfVNkiEMTQK0oEXPeyoquUk/1apqFSDmZ9N0tp0Jg=
`protect END_PROTECTED
