`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmaqV0sqUpP9wp9KrovfdWE3AE/n9+6ZNx+nSfKC3z+RplJTx5MHofX7lsKqzhYZ
XM3QG6f+V7PZ/cEvv738s3BlGWLFg17yt82ylBHoSDrU+/P8UXr7FrrwHxDIX5MQ
wFqx3JOCsyDSWFoRJJwn7OH6K5Vry/feUx/lhA63q1OnDGm8RKVb1HJVEpygHRcq
QhBxapwKc/pFGrB74M7Ntt8hoSxBY77kp1MluLiRp1e6IO50U51xxF1Dhm2iXyep
0EMU8+m2xRzFKtUhKMHbe+IXivXyIhd9rIEpt+dsK+3JJ0Je/0IHUXwaS63GcR1X
nY9S+rXYgwZss3LT+4RLqw==
`protect END_PROTECTED
