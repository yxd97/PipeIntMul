`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P05qe1x6a0AKil1oMEVD6FzmDmRaZR8aQL5D+6EUi1Ztq1akykZAA4HZMKt5KlvF
wWUTI52G+X2L9sA3lLJwDk/zekGIGbH9UX/HgIjXN9kHlz+hiTgWVYNng2x8t60Z
fMx7nSDTT+SzitTnw0qbM1Y7qh0k24j/HJUT3fniJsJbCZRLLumXABnKgAzvxx/Y
G+jcukCVRQPkvjjiflfODfUIyRI/YQCRkWjYOOwdop41SnFLZFvcvC8c2ck7ghtT
uHPkSEUBrh0h9wwPdG/ISl67CGqYQuIrfD8obG8HoKfz19wG+5Q+CYU8Wxf8F04q
XPcxkLouEtS/ba4/4FJdybpfkIDdDi1pYDAe39BV6HhLCjDAQcgNCPyX551bos7z
UTWFi0EmTJCR8qvHNWak6xnZM7jmp6cO0LpWtsLyy4XbbWz6DKnUlYY6K82k87DD
n9Xq/Jcb3biLaITQQgPQM3+cN1UIZxtV3Qvw1WpIEA7JrB2x/PhSK9yvR5AqY2xn
`protect END_PROTECTED
