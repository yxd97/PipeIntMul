`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jcNTp02fEPr7v5qfjZU00STl5rxA8cjJg2TGh9DcWnec6+qMADvVUsUcUORTsXCe
K62tln+Wbaph+IpMiGX4iR5vyxcU/FX27z+qTB9STeIoLBX+mNnMqWlOs/Aw6zYS
PXqOuAnJOxXj6QoENDW0MtjxT8LJeIUUCFaLHIvOl7dv+5tS86MJ+2CjOeFbb22S
0WljZzIuXp1QmJ7tWlbzBftXDNm3ZXhHdVOKIW5n3G8YxhcKXbCep/kBomOuTF9e
hciozM7Nh9ra5Cgw5lk8hbyHB7M5+wcRkW3JBZ3ocdTTkIEETFsUoLojFOb8h+GQ
zUzjHd153PjBzY7+7rV2enzRNwkGLmE/vl3FLYe2QyuotDrxkBXGOjNeG/pcRgwK
Cq89xkkReLBeSiqPTIGZe9jiFXmpZp+0TTBhkbgFQaO805xZ3OOxH1utSVb3Lj2C
sZq7jQeXg8pr6ePAF938gMl4bry4wdhwm4HJeE2pwOeWADnqiF2kqil1wa/DiifY
`protect END_PROTECTED
