`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
myJclSGrhFQGfQ9ZWMECtGEjhvlzs8xinYTkLReLQy+Wm4yt3prCHsNlgPvuaED3
7WOHVkpEipr1BLsU+UpiRmNAPfYCcowOcmsBun9zSxhumj+pjxdSDdolez2RNnFz
DUzn3/B+F5TNZ3999cRboNmnjSkK6zbAi6Oi+GwfzNprxqIpRDLWJGvo6Ir6aAMz
zWr2KqDWl3tf3b1zEdx0i6OhoDKeo3/NCAI2DUKNmMdoFVXsjiGYAN6jCdkWsdCr
ok2qM5e81BdLLrfAuiKNCob//59Lsd8daUntYOM0lFUbzD8RPzyMOLaVnzePKzSU
jcuQtsFmD6FQeaK1igTUdCyPnahZhdYJro1PLiR0THwuLByJi+KIqbxmhwR/M3l7
dN/CjCdh6ApaJMKDQ/pHeKD8ma8t896VNzil8GbK1kY=
`protect END_PROTECTED
