`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HiTn/tPW+KeIHEBO4RWIlgf3lRcNXZZMY5zGsx10mPNxvF7A0IpMhdsQ+jE5VqK4
Mt21fG5sKN64HO/r8ZzlKqakN/RIfKbzHMCGySEQtg8l1lLbEhxc1lNJAXF5vkoV
DyZwm55ph+Mk5opOapIfkcwj624daAnsSSX3yb3Dr36be+Q/6YB3EgzoJ89eqTI4
IUz1h46/Iii87OIMbqIjDTIYDGbKr4dbSGUoBU7pcpU3jEM4/0kr71wujDrQgnRW
p+r6G/S1ruHNzkBb+f06gFx5Xd/Jm8Vw3jc52OhPbMrv5Q0Q1LFuJgQR2NIylc31
76saz8w3l5BO2MxmQM5JpA==
`protect END_PROTECTED
