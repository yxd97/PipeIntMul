`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oq5SD/Ok5N18BenTTmSeSZwGcdP8k0Mavju54r/MCy3opSZc+iVF4bq+5oyJO0OH
dGr6sl51r64EmCZCoYUtmkoWdTJ9wqjgGIZfHYkx0U/O1tKQ2M4i0RJuReEJroh1
fio7ojs07Gvf6AXVnlDjd0IxHPhLusY2d/Zx64nSya52f8ZBWKUEYOpAGfZEUBxM
E584q5D5IPjfneKLvVsIeN5BOdGBxcvs8Bji2tJQdwdSPcfqMy4qs1D5htj5Og70
/1cWpcvOwYaFh8WUBIZEsFau4I1Pu2Y+8iPegjVQqbIaua7AhhrHpnxdZE+5ert3
S34Tiy41Vq51IipRkI7m5eeq/4Hd+4ViWKXCh/tt7fgGXp+QlLl9cip1un6xIGm1
OXUVdLuxaW8PNijVrkDkW+J0hYkjPx8tu+1piQUppm0W5ZN3S6FcrmojFtScJu0t
0GQChrdQq5k8Kbg3KVPurb6Ud5/gPCH03QMMvy35ND9XzMVugwtYoqTT0EhOgeXN
oJxW6hU2eP6VEONj7RacMd2+mTP2smHs3YWhQhcxAgj0ynueIhEkOj8WNXMz43Ws
ysS/HXcUqz0ioLi9erQfCdYSXJ7FC/OsUKzxYywc5Mmc0zPH1KeSjmWCWC/z0rjT
PW8odsHZN2uqD8BcBhlG61EoSFL31w+zO/wRFXLCPCdSsYo6Uz4wOJ6YbY+A3s6G
CPRv+xBGIP/1b/NUgIL3t1qjMvfHWmU3EmR7JU9xbFwS0LJrS9/HLDNo8qmRH71W
KQIk1gZ5CF/9HfnoUuAIRdZo5hsy1JbpTgqiXpHipX+Ijuw2zcAcXO1B6xgHDv6M
PwaCSfaNlwYyM7oFBizH/aDvdOh2z9LUbHG+Rwpf1iLoSKkEVzNG7j9aWpbJhjJo
8t3ecbpQynh0HTxjapGD23rn0eZqcI8bRfsA0dfaKMOdYEULm0zEbOM4WytN+r4I
vHiXA/OjVw/XJVFEt7sWeULj3dg7YwI5TdftDYMqn/sefZQKH+IAOasbr6NGFmGV
i//zdACALhgMGHRWAGNDLmDhxkwgv5+tDmTd5cZQejjI132IsZhWrSmY3/BvZ9kJ
VQA5numAoDvcOr7enXiT7ofrQ2Ll+bEweC67MQJMwS2QAIxMgvaQWv2Sj3ICYZ+C
CbTaR8cAnLh0cfcIaFbEddeBlk2ti3ZUH7D+75RWOnifURLD0s7QDyZ/ABcZCbxb
k6tukOhcBho9HD0JHwPdavLl2car/t6NS0k4ygAVhvh/aNWbt6qHmCnDwfsmYdp7
4Obc1hEVSOqGHOV8sLpuQqPgi8OWYJIHKNP0PmL/GwWiShGWnINVve0YlgB6L8vo
cKjt6JHZ5ziVOcerdso5O4/ibfb6smFiGDsYdl+RmzMss6+Qd89dc7hN52Xnkg1m
ISF3KZP4Aed4I2H/EE43vRkj54JJWXU+2YNnvQsjzXmveWHWo5CcDVV2iGjspFbD
2LSJRyN5ByhCKF5LVoU8pIGiDZTBSXURCz0TCcDYEd3C0U5wKl/gMVb6X2cHPFGV
+IC9p+ZIOk8YnDv73iRbnKqI3/QVC2l8W7IJ5+8mpvEsbBc64IxC9DOiapYeDABe
YoGQW5Y4JxK4xu4KEl/39TiNf1Ui1SkTEjC9DjiFOoe2CZn0FkBYmGOptulP0qZv
SNLw5b2bjD+yhGf21lxUCYwqPVS7ZwY9rE/SQLZpxdwD+FZcQNUHLX+MSwpUpgGL
11LKBpihB8WtpRkrZbVrO+7KKUnSyedl2yYzVvvjpV/JXcGmgFIShTZwvip7UDyl
vApSHb2V2quSlNSFbVIRbzoGGK4Q8zw1zfu+JcG9Vc5QrZrLDYtZAysEYrjN3tuF
2VpjrlGJGSobB/gMMrEcZDrdrCIoTKcB09ZlrJX39UnyzEaHX10LsS6+1+Qy2uv9
3PygiebEOFKGIDGC8x9nLMNvxAr60DmrxFk2lkxx+RcmnUgzu5OB6NkkvXuRokYo
ZpdnTscDs10pynL6iFqS2Yw6tpBvIlC3Ocusg2IQaHJuAF96on4Dkl3dDgpA1BQB
cTtRGO5pE5qJGqc9jzRO6oN+9qF7bLaPgr4FXBGrP39ATyNrDOqNzMfQnNp+pVDr
m707IiaJRQL+xTeuxsRFdMOMEsyPR6Osxr3E73aS3yVKDwkYXB8Z/en+6uqyHwjF
UOIY2rb9m1zdQteRVXjq/m85Qgavgff9L/cPwMRzcLMjkhxnozzjdkIWPVeZDPKq
OLwlCmgED06w6WQIZPW+s3q0sQxqkNq9AK//m6CeYMtmBmtuIoMCtm0HFK/jSKqm
AS7Iuc/TrEFMjhdD7SF84mGExVg5DZCbPhobhpGDuLvq/4HJeDpKlAPxdYYiqKbS
+Y5yj3uHx0Wx0OR8vfRZq/jk/IsAAlShnEvTQkPBAgExXv1Yk7bYTUMkGE/MkrKG
0P+M63lvmiHQJyx35XO/ETpMYfwrBMCtgvy7kLXrETl7j/hBaFsyPWULHQfB1sac
ECVYX1kmBgPeIHHpU8ZUbp5M9050opY4dZY+QfOlzOZ8lDBsJjwWsLVibX+y3ggR
SYzOuGVOcEHiGFTtQUW/yHrCRPv5LVPynspsP3fiRpfRtQZzj1pWqQswXLhDZRGi
SdmNx2DBH7w/CLrA1PTgDOCn3QNns3X6t3+hvYkzyu03zCYVmTjan+4f+ALKAkQG
Hy72B/KlbOqWsHGPZJDtQgKxUb3zowug4mcO3fit7H84Ls4E+DZPRCESn8tj7oUT
KH044EqMsXuLZmUw3iHDZH/gWVbvRK3l3E1RxrECut+zvzJEsYEI71IvUDQqR90r
A6qgENs5UFADoT9jKBFY3r0jfHzI99BB9jw+OeNhtCm/Ev50U7gh6DwAd/zFIxcG
M6uzkdBsBOGgBnkdRN3qAm/RxvtXUKuRFYPueqrNYe7QyGaD9UTGyiUS7DTKCcQv
qLnTJHoPqxVbhHCU5bEO0HCKGUpbGWQ5ZRzLO2aTOVM=
`protect END_PROTECTED
