`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCjWv1VlH2jX9yP+o0Bm40jPbHkEIQRiIz+vxO3mOhB+kn3jnjMeYZrbgeCP3Wva
2V+RqVM0QBqnI1tRIk9sGCsG0UbjoLt1GXz05hA8odD50nEz/sFekJRybPJEjEwh
JF6at08ENx9fJZH1ehR6F7GaZHOWEVJxBkRCbA/1iqSYMlOvoZIWs2acU4TzBEKK
AVbIcilc1wxdnPwLsna7+jsoTwJJrdK+tbc6G2dEgjSXRiQXcVAwlaPG5TWJ3zMm
mUnTOLnTA8e/imRgfOwgyJS281DjnaDwy4qKLdUDf0XMvoPQxrsxYqwzwRRt7U7K
XqYBDQDZgFgSwMxFNzKkurBzlOQVsNGlgSZjlUmnOTeoYAZaxpLw9BJQ8fJq4EX9
QF1s2TlAJjLh2cg5sChJZnfS54RG/waKrD3X4OKFvcUCYbROy4ouXk8CphYGnwfb
4dD/r9aP/hDonBsWV8sARnaxjNUO1CUh+3tFCn7ALVAWYIlvbwmR7G0bE3GGkWQC
`protect END_PROTECTED
