`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nkzkbDr6VuTjrZjWtWv3PY/fdJ/OXNZpq90O8qzEJmvAd2P/LzD7rRRYbbkYupsh
cK8FgV62pkWR/9Xt0CCYx0IY1+AFGifrpvflFbcFJp1hF5V3oHK7uEM7CfgotW0G
KkXEcpgU2tNC8vWMlIp/BwB8MAVuVz6gO5VJVmbD2jUwzRUW2oWLw8aqLZ6v+4XB
K0nowomZ7LdDRzq91twvhizcg5bPg3z+mj3eX/LMkuT5jgtgOTXro+Rfdnf3kbL5
ReW5zXq+hQKHuFrMY7I9Hgk7/tOBHeJHO7SwhN1U7iaKiayHSZy5b8+7c/jmyK7q
E2rWi7W9tUlbKFbTMGFUT8FMztK/INlSXCwcsln/QZMLG77KEUeJtVosmtaMyHd5
XII2S1x9LIbKH9ww0yKRxoHLY5QUZbGcZhQuIdNLevU6kfPRBNwmoiPDzJryGNU7
`protect END_PROTECTED
