`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/3kpzMznVDIvfMYIQY+kkDM47XiyD9oWLzmirD0UioMOTnKhB4OzjGBznuN8lId
BTabZdusV72z0r5fO9rdCS3SphgG1jcpn+ZwpJaxtu17cfB5YhL+24+joSseluAA
PXNE1qB9Ab71YZiaI/k45XiZXMkIGxTqvoD64JNYoHcSlyo5cVTOBl7rM1w0rXSx
QIa2arx4j1WeZm9x1HTMwwoRTvXjc8893OlqEGbtcYHIrnnq0YvlQIz982Ns0ssg
AovD/E3HuRTeeKBTY1J3NfzUohPS65lp/ZXHSo0/pXtHVz7giccE9m9fCwlCKyDJ
JTiOKJAnaRiyl07z6f4gsK+uTap7c4hR8hDkH2Ahf/RlkzDUPBnz7eeoXQO9Ue4d
qm1f3mgcEImdXfaCtCqjxwP72545vSc0HLR9IODXk6PNIXZ3EgDKViSNnzArw3pG
sVcBq37q64oJLABeVf42U0C8gnaDE3v0lKFV4U76lw1MqLmey/zCqggnw54VwCb9
`protect END_PROTECTED
