`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HmsSv8IEPaXAjGba0cQcvEnqbstnBlFJuFXpyLpELo9TR37GCyRJQbgzFiYcnz3E
epfmGwtvdC0VpJXfsExOYmwfZc3+By48MdVDMItiPs904SqfFM/J4O25NKKmXBwA
ehTDpbpGMU5RDiX+BfB8dM8xVXqMin+b/cNCcSaqdYK3tJjaLS6squ0K+2LeK7fE
8ZoUD0yzPC0WCfKYNfbEVNnimmgjb1/YUvuXRMgqVnC/5HhtAmDi8zd4UXr+qrNy
wXwJOsM+kM7PLrHOR1C8qaOTDM27W3Ps4GKlvnrFadY=
`protect END_PROTECTED
