`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70YD26X89Y1NFOaN9vUyPUW1A1A0fe0mQ6P22hCGPPph+83QGI39mPUui4hkhwPO
9DpQkrE/5gcX24USenckpiiVuLc2tVawnxfc132Q8LBTq08jUy/m5cAUifOqKO4l
JWUBsHo3iTOu4zlX3LYCcN7iAUu9nFGdNnjG8iThKYSDFlkHgQkvNMVfl+HhRvaC
lux03l0DDBvBL+26dJ1co/hcB9ambjzbXZUp9oKsvfsLVmN+EegXMl27yKX8GyUu
imQcyKj0jZWm6ASNUzddB/mrOo5rsB1qUxWiH1cj87j8UspgRCdY+l9PKg7xAp+z
DbGyYSoYtoF5wo/SsE+kzAVPiAeX5+SZbBm62UIc5hnJQi9X8K+CEitFlC1VS4U/
UF0DjFeF4zjFINCKosbuyvmb9m5fol+WRRaxN3Kpw/4yfOZivHxV1hI0NmdsvGNG
yMf1KdjGgcldRCpYCKTBFZ5zU260QyKxFU/WbiOGOhLn7NpKydIE/HtMzKgfyMcF
`protect END_PROTECTED
