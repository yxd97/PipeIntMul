`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzuv4PcGIVwadXXom4RI7fLJz0TFhKa6RPs8MCylBkX/dDMhhsMCBp11i67wwRus
90d6Re9tgtazvFJhNoYfU17gZKzKrOcTabuiCu5y41GkktGeWDasGJ98v1+ohYS2
ZC7ToYLq8OBXmZwFWDvzQWAi6izkJfM71Qz99zXeXmKrHc4g2VP7mVmaKzH3e6uJ
Ho4uWijU9q5HElGPnWql/B1qLaqwh2n26h+n+erFxcGi4EqBiFVBeKBZgAiqTNQG
hQoj1ogwjZ2Qz3OXNRvweqyjNShp3T1TbH2oxZvA06lwq93P7HJmMFyTE9IPNc9O
Cl6sEvfPJx8J1Il8FR/N73hwiKr3R2FlV2piKgTdEFOgdbfG8ab7UsCGp+i3p2Ts
`protect END_PROTECTED
