`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BsLzKcXLg7VRPdEBcoWdF2uzgGrWQNN7R/UhiZwdGsbVbIsE1Gamcd7rwJ2KD/4C
P4rxdkHew19bb0NC5cMLQKLjrE4KQXsXMgayZ2JpjAS5aeebbAm7tkLK0jjQGjV0
flbRHhk/jUayHU+hPAyp7ulRSmYtEG9tSnRha+C6Wcm0gCiPLnGSrJI95E4NYULN
vdsSmiPr4dxW5j79Nndu2+DB8Ah01POlfn5WXZdb9jNW/PWxIpDbxMoujISRi9tU
i01rZhWRjrSo0oVztCoTApXxn66YZApYbxyY9kzPGdI=
`protect END_PROTECTED
