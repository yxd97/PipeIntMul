`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SdUwbwIiXQYiOiJhz+0Bw8EX4QwdslPxUnRLA2epLVyzvnPWqAt8VE/ksJtLDi2F
Co0EYFQPwygS0i47rLqk5OI91rluQKV0rtbORRvNCJQgc8juhRRoHQDGRLZy7/k1
iv6La6EIPh5+sRH8ulUqfvve65a4VmIFK8MufbjGGV5djtGdWtTyOjrs6GcxlX+/
LUBxslCqb3cT1AjF2HA+vMW07Awy5jfpxQPxq0Ci3tqckwI6lsQzSWSMUNFVCyrv
WvC5T+7sxrrjyQECH6bJQNt1wPQhd3aDOcFCjg8SjXFK7Fe7BJAN+7kdvLKn1Oew
UDZLMuEYTu4i5aS/xaN99er+63M+CjyvKd/MzlqlAZLn5pDyElnVTEOmkXisDtmP
ppHCEKZ/Tnd4mcyUQF6tp1AaNZuy12ko+FHT170AWbBFiP8wY1miCH24J8PDFf9/
cNndU9GyqUr+vBxMyNmNiHiD9ymrmt4XG5+BHEctM3/rPHXLOymYq7yDTksDFPlf
5xbpROn/X5BRMymuawtJrTW+NQAsMZkyum+FOIoex5s62MZAXBJXI9q0y8qEGVuM
6NKz0xlrNYV1w+nNNGIAUtyaP4wIJAjK4Tc/moVUOcfVVPDVg7U58JMlCCEx+wtm
SrPmJaZiQ51XGs8dNrPk6desVbWAIHm6TSEeGhUignI=
`protect END_PROTECTED
