`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SGnmXL8hcdbjTkuIyI2uvNyc0FFmO/ruvSBGFnxYMkGCUANk6ZstRS//JgfKzmFQ
71plja8ONWuasew4+Zrv7oYogUH20CXhTJccmJnzVD1xfngnQ2qrI+YP74Fa44D0
hGpxyJ3NHIZdsHCal3cdWpIT0YKIgMjGH2oeFnGsYVS8hsMkxQaN0hFbGQhnnQFn
DVoLwC8cQ4iqsQphh41frFerPFIyHHmZUCTbQf2lViQjN8QY0WMkQkfutVtAnuOn
/Jxn7T/MmoHBVXknq89AdMfbLK+UFhc9AtqANsVW57PGi6yykGzSfCJkaJRRWpnG
i1+fk466cnMR2T6oBaV91A==
`protect END_PROTECTED
