`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GYPgYbOGBIbXtlkkSORVJBDJaGkvnidKQK5OBtJi3NMYWAn/ENIEkBlxBlxialaW
8cl9Zw7hH85SVOCS4UNsmMVYLetBQf76bE+uuMFHEYesOA+gv2GAlHt0GRcKsBnZ
duK1ciLlr7mnJJbANVklt9OLUJQVgJq55fuYHW5bpSLv2CM47sSe1mscbJYmtU3h
iC3FCVmqQbDn8114PpoKEXktoOUBTKIEc5+nfclFXn0TnnX5UxZANZrYvgLBeW39
CX1HGDfhsYR8vMwmG+FpylfoAlmRVMVTgDDA+L9n1w7tfmQWVLgfEndRXj6aMptP
dmmKPd1F+YEWoL9o9RM75W+v9sXZ8Dz5+2+RMNK/AsBqnPhonZFAW5x0wA6hoQ6j
qvY3c8FzVbNNCoOY3TwrYrbOAgBQSkViqV8OHYl3px8=
`protect END_PROTECTED
