`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FhVGNhetgIT+7YAMmYekytsAdOvqWVDpss7DK+M8NJf7CsOePi/9HLxJS8F+Amue
9vwN/ajniaFKMbMzPhyk7/FhF+jMLV6IxU468YiwAHKFJAS11mEzqoVsqlubryee
1DjN9ZGbdlANrqs595ar9SmZ3FzI1Ug9F2EckthU2axcsPUsa0HlxtotdiwZ7s+/
s5+SWxr+TjzH3RN/RCSH4VzuoiU8f+R1ZaaoXc8ItRbiEdgoNLuCjcg/SM76XedL
MSlz5QO+B7BsqhvEBkZKdqgzEqvO2HsC6exjG00B9MZinjLn/b2NCFAeQEUY+Ll2
zM2/e9JfkoExELCgAtV8FR/rme6lLTIMWPEja7IzAiUdgTrUj/Sxr/9LIDDOxGtu
Y/LA7ATtLV6FjNa4MCrtjfZbhgYX+/S3h0pJyqStS3qYkqU8NPolCV3KOp3Bb1y7
TEhspiIWXrnOXwk9zro5MKRN1PMmw5OGyK690gaayVqBjzjyVc/zbDZyOqTZS38M
f58qWsFDvOQeMkZ5avHjgXv/b/cTHwh/tWcq1UvvpMIV3smNdjY1ZH8vMgU1cGRz
aWpJCo98hrslkuycbtdlEA==
`protect END_PROTECTED
