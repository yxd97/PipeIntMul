`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
krjSIHi31vEAYPcwgfCHNZcsCFs+KHq8mK0v/9TrEYfc8GvEyNV2jvH7HcXDSK5D
uJURI8iZgfE1N3I5kV4FnJ2rhKD0PIkjc3iRIpw2btJKk6zjCy6z2jTlrIF/Yp/6
8eFbTeHpU/7mKXkwrJ7RBj75OJoqVxURHSZ/zBBbKBssj04VLXuXtH4eVbgi5qe3
qpk3N92uCBrV+Lmp4js9+3Qjh7v7eI+goHoliTD2bDuujDu41yV9pgCbTFHlaL1r
6L7J8un5Fsz7q7qqYwXuNwu0TsdwERhdbzTyzG9wMXNpt5FF/erv1qPAnY4dy3PW
sJLkDWbt6Rad1HtVTuwTAQ==
`protect END_PROTECTED
