`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VhKlbEFAN/G/X3VmAzdntPyavO7On28kmhvRrZrsKrW9iK7DN5Ase0D0WvN4i2rB
nxPQMxrBW0daVo6K8dN3HUoJxcTxWmyrF5qgTtY/nL9hGrJGsc9yNEbTw+nUMOB4
6y2Qu2Z3mLJvcGDzFwvCmncWJBT8fgu8iC0+yjf0qGGbMMNSSXVzAEUN7DxwX4tN
ndGyM6kpbmlVOlRsrc/AB8Ed1s1+TYt+Af6C3XYRYGIDwVKw1270MkwSvBdPsr8n
tpml8ExRVP7wDy9jOkI4RtUiSXlplSpY1TfDODMxxGrDAr27j466ny9pXPP0kHV1
67mA1ZTwoVvyPDATHGWnhrKxzcdVqECYsN8I2QLERxSvE3IYqLyqS3708XXVSRC9
4m7tjjh4ZOYqGU1Y6mZOItW23B1NhJ9XgCHT9oinMDiw9TiArqavEYMk/PHYFgG0
D3pCwJF6MUgGaLrTFMQtYKC7VM9TiyAu11WUGB7Uh+0=
`protect END_PROTECTED
