`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8R75NMQM0TOz1XNFo8yWjoURJTXjRHbjPXNAAUkAdiIOCxqHMN82c+NA2W9iibSx
j+kzRWmq1GHpc3WqDHERPRjdrKJ9VUoVvfBJ2C3qT2yAI7ATqBf8bh5MqvEj9vBb
0Buq5bdnO8jlhmxEOefLnU06qHMkWra8Gozqe79mi8oo9C3j/CXXN4d+uC+iUhIT
U94/o0zUJI3omD8E7KR9igbaDu8L/MFckG3TWMw+dMyLvqWRlLC4vC5+ZdABUsJw
mCn4LYHaP2sCJ5suehFnrGwiDsRgnEGLBp7zoYivwzw=
`protect END_PROTECTED
