`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oOLif8pQY87qyaoMPiVSBCbTwbCsPwEFbczu9GxeXo8kQxjznU8b0RwTwM9D/TiW
aG84rNcqIWpDs0J/gEAQnx3xyVGkPIxmQr2TjTE5nvOchWWNIqtxsM2H6jIyWvsg
bscV8fUDi3oy6kmZGVZ1lPYb9xh3cx52VD8j7lhR/oCHv/s5wpwzrzSNE+ajIhB/
yT3kLPTYi1azpqd0wgUp1x3VlYe63Ozj8Rx2sahnWsggobosRbQrCuVWxEkx0RYn
iAo5MAWy4lWP41JKzgjeegGSkp/oVLaxZsuwqDV5Y/cT0Oo8J+vXBiwi6bWkvT9B
tp10j8udfLmMsLIkYLNHK3I0hLxxYnpQQVHHJ+VxQ4BXL41JODb/bXCPi8/D6rJs
Ox+Uh9/LawqbUARDG4lmFg==
`protect END_PROTECTED
