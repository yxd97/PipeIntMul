`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OT4kGKqbvI3esq4l6EloWBJoxlaZLEF+29JHqYoRlDjRmvYwaY52KFVqThrOyeH0
QJN1zNR/TO3ie9TQKqqz/5oMqHjswyow0ig8VZzvCScUbLQBGhc9063AULt/M+SU
gCZIXoEBSGrTPkKL0ZpyVZzHSEEezD4UCWEwegG0AIWXO9hikO7pFMAtCGFPvHoJ
9l5Twow2LtXV02NT/xrtgxPkkFGmlXVcUfaZkaICtNQN5WF+wGPHXh/ZmgWWEH9Y
aWwxMXedSpdZA+TuDuwv2EKySFVoyTC5KHdrN6AcFe3s+8sCaz/E4BQ+GBfeaIzz
6+Srp5Y0ekSLfQSrqpTnNN6ZNQvCDYDiKOQXgUCG/L8fxrXBsc06fAZBLFe6XBP1
N+vLpTEkuMvS+TfhDw2EwUKWlohlE654iP5yS+5d6VFiQPZVn2sK1/ppXuGGuF85
3ztFi5YmoijUv3kdGpFo1JepRA+8EDmK8uYTNHljc22i5m8UZKYw57aggDCHcclq
9BvFTfMsldkxKt70LucP4UoEwJ+bWfSjolWbaO3YBz+/rEVFOSfwcDzQA4HJuJJF
YbX97/kxfiVoJXoGkuKP02kWk2Zpfxp6LJI0/kBp0QhN/IlH/LrHBrZzDm/xw8AS
9GsdThJPws5Kn8rEljo1RifXvZKN1pY6Et1iv49tawES5N+kvVqZWnPUHDmCrK8h
nYsrkqbOk/l+1si9guncfomIcSzevc4qUeYOvqMTP1XOcpr6sjUe4tXQRbAs6+6X
ciaSfMn8URYnPjRnoz74P6zwtwGQfeYXnfur1g25xz9WWGexEg6x+HJuLd0AyqeC
ciyi4dCgNwJSteVsPqYXMMl83TeMMvDrGgbM140HOXjKP7HF8ZwLdj5b4EpWxM43
Hnx4slEP3+bMBvQJRf+w1i6G3I4ilPl6BH47t/OekKGch1Wx7gxE0Tjam4eFLCqD
ZuDIU9RVozHuPDbvExxJas+sIZwhJ30+ZqvYtHOHCTP8r7uu5W+PBMwCORtJbSvy
O8UF8GRp4pzOMmDzN77alQ==
`protect END_PROTECTED
