`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+MfYMjM12JdgVox+WR02Ducdl7BjwseUPO7QLkmoXLdxnLXP7+LdqwkCSMH2bUv
q6DydJe2JwX0slJRAEq/ABoRo6nNA2jFmCcgnNiDWY4iqEaXr77qCbEdojx/RgPv
iM6XWSjLbxVhwty7yY/KoF4qXbDj+u+iCeI2EsSt+Cs1BI5VAsYS1G3RNEPITP7c
p2nc7huQCUNG6wx+NIzKQAI0ODGE9nRwjd7b7VfmWiEsVj/fBD/LLYhXaHzeSbVB
QQ735G3aHmNz9rRIA9k+BvRFw3oQ3Cufh/StxyqYvVieQWvFl5m2LmVwVuaXQcR7
tkvMatYHb5j1vZQct/S4QFLOVV+LWTr9LXMuBM6bPArb9Hn7E3vrmMsoBxpCepBT
5Jb3h1p/euDCVCI+doel8DdnMNtWnjYoM3NTUEXPYTtYSThoKAIm7fgu6pFIBrkD
3WlS9Dod6hLWmk4EQBrLfI3oYpD8PeqIMydzeqcn+U4aOp3mes0AZZ/2RA3bG7KO
mHDs5CMgifktYlBHJS0W8OsM5lW2Bome5A54ElgLfuU8HmDGflF6EttRw+dYYBDU
OOCbIiM4ACrO38J2eh1VBlQUr9/+df8CKcG0W/+rTZQcsQu3iwu10AnTXNBfnOxw
37sv+qOpnhlP3St9w/FJ1NIqh3F6GDxrX/Wf/PM5xPI1nhm/9akVeNTsbzdzMTN7
qcec6NZRmrBhcibR3LlMkEs8r0hOMerOoBCxmAf+nBiECm5GSlyYychjDVffJ9QF
qeQ59ToBOurQDN9C37tx6gRNfZgHvIU90c4SKlHS3xQilr50eRSTjxko0Eyp+oj6
ToNpRabs0idJc28V4HIEIVW0mK0ahiQISlp69eONifcemSsmGVcn/ORKxuTMse0V
B89ZOSxS2I+QgQHTA7AEee6O9fVNe0MnIEGU2DTzKDBt0TBC3j4K3zq+XgLx8Uzd
1G4Bznz8p+LlBs2hwGMKcHYBabhYavRGoTjZaTJ14OrUDvGrc7q124qRH2Rtf8CG
6EXazCc75BaUnINuqQBCfIGcmAziAl3+g8rRV4d7AREofUQ62hIN3XGKpK2Lpc3F
0JfxFf8sDcTpc/5WW2gGJaDVJKct7XToke/77i0jsFsg8mxxcwhw2QiZeGQstkye
XXPBrqE3pCgPdGNY+ZNHCJdxLqhflh2aosFJQqqi8f+GlQMGlvGHw3mDX/y52uTn
5jzTBj/E41JdsrwmCL0R21jNPwgVa+Yb6CLR9pxMP2nrCCMsrg+EDbL0ZaAPGo9q
MKYOZs1oOi2KyHkRqxJrESN8OwPDniySgcJMMJaD9zZRI3ed6sHRlzU1QMKMrrub
pBppsAlkoeIE3T5Si1CahbhkCYQIb01+f8dUMzCyOYKzcebyC/Tik/YTVxapdZ1p
Qiz0I2QAncHxJkj9t5v/NiZgjhcp51wFGe+w3XxtYn6kvm4w3RDgQjRgA56eJvFs
7NYttqAN/gYsWl4dlHz9bk2bwSt3UiNUvvBHEL0nI1k+YOg5ItZow0v2Fiy6rNWN
TSJX+Fp3RjjvjS7KLYCQn7gHWEksyhk0I8TleZu3wnGXd8NlLMf/sxITzq6VnpaR
S8+s6IQqZzMKgK4zKZWj5IYXL0ehWwOi2uriv0XIbJTUdAH4y7YP4d+EUc+Z2BtC
+sMm0jwAShKJQY7FpURnDYWcNr+2UmadgJnlCoKfQjH19c0h5J0E9JKKljAph7Yn
xTQs+AqpDZeAtRP29R2QRKzOKQEEWglfiV56UT87T/1U186fdpLqw4+k2lSMRHEX
pZep1NEMBzTY9rUixpKo1+EWl88NsNGWpr6Yee0ohlkZxN2rMYR5yafbVAGZ6jq5
8UouVLzOi0cregcV47e1DxJyPBFmb/2bRUSuslxi4N4OIHfmNXlQC+AEHJg8xNBv
gJXyKIKiKCqc4n0IlE1bzvSoKeuoP2ZBxnUezpLKvHOAbts8/if100k6WOwXcKnq
K3XU0CChMYwAEWwR7dm8CWoxOZv3MtqUnLbtcIPNK0BI+P5Uh2Cwwyni9YuJSC0r
WRHV1383big9OY7X+SUTwUqQETWLVuN2JTF5IQQnr/gJtnite3y6jokY+kRg/aky
s/cGjz7qpfAAbTITA4ky5ZXQ02iMVc0bK2DO11/6AeY1qWgl/+zV4NzxHyMdDUpm
3kahncwVyx6D5R5Nsv+ZJQo6THhIJ0GJXZ8JJxdPUkRG6MkVaIdmPWMP7XXWDXyR
DnK0dQC//PfCrkD/Inc/SyX8Q3dHQndofcnaUJ/TkihXmadfMZ0raZENs1Q5/uPv
FRtBMc/8RGJuJOQfJ9Iy7q1EOetTEjxND2f//fCxc1CBoNDknhuBE2Y2TViZ7doz
gmyPsoZfUFwvOBFLiVgiXZqZ7qpkNACoWnjnKwN6s2aCqFWTfBU0jB8t3WDRzyG4
QvpUlDcsVgOY76o9hwOo8nFbE0vDw4uokt3OcyNqLqNB7YVBpvRHqYzw8SGU6YJ8
iHb04oF/9w7MdfWCKiGhjkYJyc/nqhjuJnKVbVmqIuhSaZJomwtIM6Dy2UXjBhVo
sAUgxjmrro00UrE8q1ngkX5TAKnLwUE228MzSxpJGqsQbzN06uvCePADpLxiiHkx
g8rmaX/wV/vPt0q1KAdPs4jk5OErjPEyjemCtt3LO8nnEbt87wsvejr0g2pcxzTI
4QEuuYBBzBdCJNMoaXJgmDioLSofq9eBpCEXV5cu+lmMadFpD+Myyy/UWJN7M/Pw
s5wtL7r6I9gpcWbFST1vNVpWlTndOFoImGxYVUnVi0g+6A4J+AomANTHTAd/kd+t
1at2LVdiw6xwKI7RCsngVd3CcAlHizg0YKtsnF3XUWgSBlOC8A0VhUAEmPfBM4tT
3YxFoWEQsISwaZyTEdfckK12Pl8HrEjUSwonWauZAVvcY/al0TM1s1aH07qh+1Tj
M4ej2vYjxENV7CwbaUKN5joJEeYg+cNlOLplcZ6CFXU4Ea9bkVD2gLj7ZPmCx9+j
77DYIhASNs6zWX4scK+di6wgLrM7K5ktrtvSmzF/3EA5Txjjg8WX2aA+s0j2091r
z5/4ha57zowlYbAK/+uvouP+7oUp+NnUMO7FybCCzNDznp1z0KuoDfN5tspFp3pS
`protect END_PROTECTED
