`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
010TG5gh/gY3Lxmc01razgMnzXXo8hWCPtoWEAuqr9fwulMByNqmlEBY7kror9b4
HxoYvIqHhNe2SXC72OrWQ6JxfQk/D8quqSRqn8+kFcag41kbfgZQnBh+NQ3brlq8
vebmlkDmMDpmjaeUGL5Jm1GwJ4QMd7zEfFDkzRrYoKZXigN7lWrVzih5Px4Jtc3E
55M6LnVuHIjWYbE/F2MenmJH5mO6tDY1E2DydC2YOskHSg8ZHYoMUyV6fBpxKfdc
fmsHq/Cz+Q2TqGGM+tq7YIoA/PTKkQ6/DILTmSPEuS1AlCLhyzyI0Mgb4RNCvkyf
PCEcDlNkH/7McuxHEAv3IuPecRIYM7dVpe3LZGcVReyTa4ebC5NI03NCDcnuxDS7
j2FJhN+y+ixMF7exAwBDI3SUiKuWjwZYFJExQgAlsaj+NJuHd1MbDI6Nq4o5nPqc
LyOd1suuClV+pv2AlDxlPQCQExLzqHe2VYs6YlzwNS17D43RspSPobuCyZSTk6nF
9NBkRpBk19SLwfls10JFPtS91Q3dIWps79HoTT2JPdDbikSCFUOnGHw31TX1jwXf
vAXYyp6M9wRXNGnRNX2E2a5PfZryGq8smb56gSpy91jWPOVshikE53fyqqfc4kzH
KmMwUVyf+yoT+4Rsp1sOjAexaY+wkFWRil0HMEkCks/pfQ+zCdTFtkr9jN7Pf4/9
xW9ce+du0JOqNMnteYNtVhj1rFrD1HWbQ5Mq95ArZvjrytf/fvpZ20Tl6AhG2VF6
f4leKPmvnd1B5HUsSA0OF70sVaErTWVgAqWFebYckTo=
`protect END_PROTECTED
