`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ztC23IIZaISqh6Y5MfFTsxpbzh88SSYBefyESRYD39hCZMrnDNarCx/uifloMvZQ
V5atQD3RU1u4NO6hnYqbU6uZyXyapIVoN78iYg/f6QvD+/trVjk8Kb1W4dxxFac8
CV8ROCtztYo7CCzIciPhr7m0JAQ3TKoldlwpWDVK7uWYz0FnFtEQI0b+FfjuWSig
LQ+cb3l1DYKZ+xNgY+K+P86YxOQ4gAfX//rYO46Cd08dhGZy1cQjvl+eOgMzRJlM
EHx9PjTlnAxmaQouHtJQsLb9DZA6lGOM9Le7C/P8owNJxDJo22Y/o7mwyoFX5LKl
VgwOsYZEmnmOcVnMgPnoOfJOk79YlrGruGTK0XHAG1Q2AQwSlLENA255CxEt/XI9
AdrrnoTJFA06aXJIhzJ8kBIITFD176B/tn2nrflAFYIidO83b6wBw9lGeRWKfRR8
miob8bKtnMjCxeEv2QvnkONQf+g82c4fmiZ3+Swmbse5Iu4v57AVrlCWHMLspqyg
dGYM07F/xkyTRcB/W7xTMIr9Al6v/SULSrdcljFygVDhB/CNwZ5H2uyN5A58J4hO
6W5cQ7wTaCeNu/Bh5mivz2lrOlNu9mzReIFcQsRZPGalbCKI+dbYn/WuRriT0knG
CyGqtRAjnAsAHJHhiuDGq7XvitPvUQGcp/sc42culU7u4YsJAtQjHppt7BoavZ01
FFbkKbNo3aLt0kBKkO8pBpHsfPiaqOK5DCPZL52aRN7D17XEVTp4UFhg/4GQAKPI
P4aWksf1pRR7oGx2zQqs24VAE1QlTqEA0/xd91yRqgpA/7NAKMhCbc2/U9CY+mp2
US2MwhUpmYdau5EAtSy0A2GTlDiI7jRMSsKpxnspbo72947+rZkaEIFlW7uu0+VZ
9XukdNfB0AgfrkFnKyV57MCO/wz6XsAvdmfVZlUMfLuOopeXFjutBIsPdnVJcrpc
XFbsySItgDhVEpvwARSsOad++uHaF4/BVr0qW2DKtmD+xsJD59eAilncUbFpRiyp
feZ4+qnYBhSUyyhp5JfVPEv0SxQ14nG2k2CInF7B7FDxBp5oFWGvKXlVBdYXWEMN
m7wlqsrB/WTl+EZ/HhaQMyRi5/V8dKNsW2lD5OhiNSiDaFnSThaAj4XAEflkrMg6
GVreAr27378D73Lx1duDAVmLtB9HOJ+CAEFvf5/oF2RJLTd7Zy3P8KgXObRn5Tbu
Azw8g8mg3OmTgmVtYyeYo19guq1hfmvAkwyxhCrShWrWW4yiXXfDVx/++ScE6OKG
emTRmI+m7aRYMjRl8L165ML9nJHnvnTxmnK6HEU6xIVKZeHLcWOP7SjjzCDM4+WH
UdqGVlUgrcD9qixtefoXlW4bFFbxRM2cN2/+fPWFUZGZNSe/rUnGKP5WgiPlhYGP
RvO5sKrYnYgHAa/zonjBYxoOdBcLKqhzwTGeO4+sC/gBW0tVwEDvM65Ui+T/O02e
EZaXqYp8x5yoQwZ1g7JWLy1H26Vt0e7gkrLJWBaAxlSB8qZ231xjljY3gTwrwZfE
xY2eD50gxHmz0HH+l1bTxPB7WBEMTRaSZYzRLttyoWyVo8jfZz+lJk3Rlgsr3Kqx
4XfPhYxmjNF4IXmXbvmVTNouLvvUAfhMzEDYLnRLBrGjcAH8Cqi0omC5WGDlhhtN
aUNv3awGcf4k8EtgkWqt8l2IH+1QXJwMdoVcmNLb9UOwzNtXC4KiWcHWsmkxBQmf
0L1dILAIaHyXcOhGOcNPSrLO8zR2GJmPweSndabjG90MxeMtZLTis1koE82hSLj4
wGfB8rVBiNZ7K4fz94jraYN/17GTMscZqibDdOzAzjk=
`protect END_PROTECTED
