`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tPiGVTlJMVzF3DU0mBy1Ufp5qGu17u86m8/e08qPYnKLmiYgpFVj9jYzTLMJlnEG
ftzt1TfbGXULVIq8KAL3QcQ6EMjG0m/KYFXjnlGpVgPuBBvsuR/efdxlFPXwJCPl
i3AW7qGDYFvb5CLUfcgelN7aw/OC7tXxh5h/TfyWoOnHmV8JgADWwpB99JX6coKb
IAdTsViUS64KvxykQJIIUztgYSNbqcrAzSJ/D8n6MAcUqQbnL4JqL26Zp9JYsVbO
BGn5y4rLKx8xWZS2VUievV3vePMk8ubcy0n3NlsdlPcJbQDXFRw8WS+sVy/qgkXJ
FkDpaLApbQmT9czUxNMbrxhu3+8t8dzhbUnpGDyuiFWe6DPIagrpdOxud9/Jsifq
6wIsmrV2JWQ6mksJ68Op5dYSk53gmdXZ1IQ9LkaVim+IUAcrJC1i8pVPm4dnrszz
/G0vEddFbnlDNt2nkazjRAR20R7+2zYMfOEOVLrS1t9dDv1Qre0XiNx4vSw8IqMq
hZK23Uy3vNvnHkrkf9V+w2t/Kup7GQfxGoZLHynDC80ZRvBxdKWKLzZVdzpIUbQ8
Dn1hJFI/47d4lLuVE/beJ7kyZM83Gig5BLVRWq10UpuVc9tExDvmnq1l0Exur6xA
XW+c/6bUHhOc5TAqxjoXVw6CTTGNN22M/JPBg6b74fXvbHHb7SMOpsSAsnMjVW/M
4XGS48wypc0NMrDPis3pmhnO/qD90Zf6DLDolvvXyGciXx2CdLynLotvksiGLzyQ
JmmP9e1bL7NIsDocSWSIy43tkrygKienDpZh6fI8oCjI5Xmc1AN8ItkP/UEoT9T1
SXD5QWfcF8zou0mUxFh0oVX9qgCx5oH/YyZWpxbd2AdgO1zuLKFujz2fr5YcSHpS
FEhxyUl8dZH4esEs34hCv+Tjid36Nz5Wgg+VBzQJ2b3jnLYorCFCobtTPZpdN/1N
1EvhfVMW/j+B6FkL4Njokg==
`protect END_PROTECTED
