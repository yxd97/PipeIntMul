`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/fY405/q70mZUOGOcGMx0GAEyaWofAye7j9Gu1WN1rEEwatU6XTzDvNOz6tKCkB
wmsyCNequVpb82QYho9V7dKl8BWG56CkKc+6jvuu46XMA7iRLi/G/6q20e0CNcp+
P4gvzDtQ2zG5/mos+djUt6s0JJhzlUh18LU6Cqi5qGQVB1Wcqu4coG1TFVqZrzhk
n+pqjQg33Fm3SMb6XhcxvAYx3fdAg6fITuBpisNv6EmkqYN0g9okVa4YF+yDZ5o1
JrCQw2oIRrWlu5ahKPr93OjwcfTMqFSPKd53/9NOdv5rvXYBA9S8IW+e6Vdi7Me7
ZOZD5KWZ5NaIFfbz5KPZUhdVK019QD88M8X6LQxWGBWBSe8WNkKB+aVYcUUVmynN
`protect END_PROTECTED
