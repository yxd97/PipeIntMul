`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyCsPe9jWYdNUTF6yJadJUfvCOofQRwwNkgMRTYFAAEmJLScghQLVHJNyCWeenxR
2YJwn0JcEQhUQsbzA/wJzcScKcdyNhrFt+lOZyWoc8GFb6sdJu1pI7DzRoafoIQv
PF8RFSpdFq3Hvwl2IoeBrljfn1r3ePcpccBkh5nX2rl7BobkyQzkQeKcbrFMqd/5
VIinm3U76SwC4GYJga17X54D7myTHsTb+eorJUtbOyZc5E5VVT14SJyEjf8D3wg5
LwuoCvxxvf2xAEyU0oLfHzxN5CMa5MxH8rYZrbWzKzNb6j0by0F07YuNJiIIQZLX
BC83I719xdxJgCTQci1QaTrpd7LKHm6vFd+VeeTdEo0iW0LkHObgNaqFLtgLUTAC
H5RuZqLSQQ78P7MzntiHTXX9K0Tuiy9eSO/oXQDNK+CoLb+M3bfd+haUT5SRraoY
iQjIHqQegHh0b3JR1lyTBz7uF8owo7UzavqFhECbDC/qvLI+tnPCTvCOyVzelIg/
`protect END_PROTECTED
