`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NOO3irDsFDzY0m6AKdidj+7jAWexfl3n+VdNaqZ7WmORXQobiSLRecavtWg+mfOx
pLSl6A1vp/VjCBqS94JrTogHSZ/uG8efeIogPthnpiMtVT/BBHGnw3oteT01xbxJ
GfgWyeeQsXGWRUflnd0u2efq6OzqIw1vPFDZFAIbF7UTMrMG/we/590x2d74T38m
iVKMkjkhOI/ljBP8uu4Ougt05peZ1HTueQeSduq3zwZJ9aQjUmeC6DW2uKJktHdY
HewR0SRSLRSYF0xFKZJMo8xG9lB/idSqMIBihq6SseWewmTdGdnS65SU9BAWasqO
y1uT+QuzD+JRD9Ql648kopEb4NzvjlOmX4p0rBHObGQbX5ZkZkgElhl5MZPVakzd
AeODhUBLn6PIr8SMvP/mf3H0o4dfDjpHOngSSUBZyAOahCxtAxqVG+1n0lr2/EJv
k/WaFEJR/IHSnS5k2R3NrrYuNjYbEN/nOKEBHWxeQ7W3wIB9M+u0MhG1ZJWVxIfq
yTOLMiaDBaCY3cMNCSK1T9iaHptvGcr/3wHPhZMycvWJOntacFlrnq4ritZzyD0/
sO3gzXA5oX9H7/8mdf6NtffLorvr+RIN3W+seeN/Gkp9UtueDCOag5Ckq8w8xBUv
w/ngdzYky3LacvBJonx0dlYpKdTdPMWSEIaBn59o9Ul9gIfk4xs9ftiNU94KZVgb
`protect END_PROTECTED
