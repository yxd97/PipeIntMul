`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rKTgdv5pYFlOO6bs33M6y+H0y8ZuAZ2JQxZgzLGNWHjvHNTXD6go/Fvq/CgHF4I
4qZsJzjHnBbR8Xohh0m44tehi0HMLCqfgsFSe1ICJ1Iajn0jz5N+CZRAiUqzPpOL
ZMd9wCjXmN6EnJHsMmDfkD75Xj0j2Rw+ask8/7ObfhQXcpDkoLGiwQi1geSw0DgN
ZydncA4eudXWUeM2iLHrSXxe3afHXmF88wYPxcfXcmcMkPvEQ7FtNBpsdsCsGZOx
gqvFkky/1U/u4mphtPDXaQ1snt8FfF/OAKLXVk1KB+NmZPvJTN31LwGBkxU2OIBF
q/qY1wZS8kg+RQtxKdB+PQ==
`protect END_PROTECTED
