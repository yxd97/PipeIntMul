`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LI091wG1kV4bQjbl2VJAnd/846U74X/UEjlwhbijsxccEi7u3aE/172STKISJgRQ
uK/UeLPLfrQ1DMIFcLXgSCY2MBbwL0u0/sHpGasjQ7yZYHht2JW/PLniRZPCsUWr
sgAlmQrhcelYRNijYjIxJUsKRy6b2G1Vd7vdvT8FbBB18LlsgAT5A6/rq1nFo28u
bSWH+4OUbRlEGz4iubXw3erRBZGVfnbHzeSToqYuOJsKupnMnaa0ccEDCK4EOseG
02W0RV4OOGDJ7dmUnO+5SybPIGSdJqOD5E7qRF8mFiSomnZF9ATBAzniO+da697u
ocJtbm06/PJsw3URzPilNpUf6nVu/yQrfyXofPr7O/LrP6zVm6Wqtk9M/hYOcw1O
q/H6lD5DhNCFX2xNTg3dXA9bO3/+Umo3uZgw0EbZ0Unf7GTZ1ea8iKbFqH5ehJpT
V/1cKZrW9eyGT65mpJ6K5f1gyPD9+59yWjLP78/btwCxxxhVEQBEELGtcwsLJiuX
6EhSQ8chxWqBqwDrF1ZEIEUzsNJHavo4jTd99ikxMfk=
`protect END_PROTECTED
