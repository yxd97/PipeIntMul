`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2KQp67Ve+tURGJc9PD+TZd9+HIIecxgbC7BPkPErJkBul0UGjsP84nqyThykzxji
q910YjEvbt+7ESHSnRlnsdaeBMfU0blQkVvzS9CJU+vC0jOmb3mxfvxYKHzMGZyE
IKZnmD85AzrEy67GwUObE8ymtRVVUj2JOvPWDfsnFgf0TBDANMyBZgwJ6TBuktN6
aev7v/drqaVpyqzFWXdNAxPN9qjRxDQdSAD67XkcSVdUutcSP0xB33vyo10gFSFZ
hCsWAz6ucBSqvMFV/LZ7XZhd5evLbDLPeZI6x8IhWukysioBkS07ckrovbM6p7lS
5UJwgYj6aE6uI7DMZlck97kplzhKx9hmb3Fcrst/inS4eQYzGVhhKRQpQAho0GCl
DB9bPeHmBY3kd0olOA9k6g==
`protect END_PROTECTED
