`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJAE3E6JyxPFQpj3whzAryC1EpZEtnnYIriH68aNZ15cQRizAXsMuMl06RW8o/6q
mtOzvBdyld6zVFFKDdfKw2OcxH1gLAvj2peIu2VTY8Y6mdTqKGKDLzYPPEUZ2zvt
uFS79PuWbHITArii0nPD/K44FYtjkAEiNr8iVIJIKxfzTCvojGg25ZcsJiR02OY4
BBBF+vr/5rLOLtkE/EHU7T+71yzwxXBFc4TeubfVkmueldHtPcpPzwT8tAWqQWJB
7C7qdsbY95onWWIabamo1QlsPdAKjtBQsDyQDR8NaLlL9xCrTFiLzQ67YRvIdE2R
ugP3/O/LTzG1iGo2yN90UysxwtCXfOoHXcWnMVVosiBfDCGa3RQAIy5MK8wzySSv
eLzSBp10E3+rdBss0KrtXhQhQJTxSh3DdofDOc9zw1o=
`protect END_PROTECTED
