`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bUZTRe91Mf/S6TY4zWWVooMroJfCs4SEIuoTNO0MQC4ZcH500U77XaAz0VRlzdJn
7xh6pwbSxUAU7VxWmepZ1sdv3K30su7flU83nofwAs4PBxFqe0uzzenFgIvP8ias
w/4pK/cRS8lIaXSSG+9PHvaPDv6+J7ayNqjkI+jpqZ71qE1zwblVnP6ycwL96jHV
WSjDYcoF2C/cBBmn2ZN11IqP/qtqHXXIMUgkaJZaZrXgB2YbQ4z4AiIKdVn6x2ig
z/VO8p6q9bk1Zc90Dy01l4VESewjEfiYv6vRhrqM9hZUO/O8WfSuLEFbAHtW7Npr
E+COQdUhlHpR1LAfPOjI9A==
`protect END_PROTECTED
