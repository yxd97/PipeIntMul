`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QHYyNreG6p34CarQhph1qVhIkJr00GEU2rCEY7loxqxDUd244mv00mHvWdLnpIxf
/gLWFnAK4HcPI8CYA8b2xUq0/1PdJYYSDZea/XnRZmTM9Ik17ynQbuiUBQpmWhNc
2+XsToj3HlST0wjFrqPDXxZ8XtM/bW31TzQnmxYPeFQ+FyI+RDkXZc8suXXAbO1w
q51v+Qs5v1TVyr978VKpV8ViqajZetpta2OaG1DoeMXlYrHadeNwvOkJI5j4PcgM
rURutxFsWfnQeoAk/eCaenuCGSNkVyBrimJgAnrF7MV5xLAI5LJMQFPG/TJ/l9Sj
cVCn2W+Lhud40uCv5bBiH4xbD06QJmoWyaKLbM7l7q2eaG+NkOyqZNbwwKiaRTrC
yAwCDncozyEZplSyp6uLmrSuxo6byoZn57nkIbBbEnc=
`protect END_PROTECTED
