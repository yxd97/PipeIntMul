`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yxuq9kKrxJUiBibibPQ7j1sd75kiR3wATvZRwazW2DGAY67E5j5SZJ7/JRHIQkMN
baYxgFxsiYUrhXeoTxOsy/IpOeP4EX54601r+4KIbMlHmH4/tmvP13NHDTn+Q/Fe
Y0jNgSx3VGhCNY6A1pjy94mQM21O70iRO0UM/2jqrlhnLcYgipjg6ruroMjL9ZXr
ez2Zatyspv2Mt7si+Uslp1dqh0qwuNPQO//p5VBH4qRf/YoyXBEhvxHUCfrDQ3qI
EoAxrSvkkdq0n4//Kn/1Om/8cQ9eHEPjlYYu1LS52kn66ClrVO3RNf9kQsFRHgXM
GW09eax0lPAStaQ11DG6BlxedPU0gCPTgmT69fGoplxWskO0ttoOxQrofXgtcB4r
ooY1dcff3mezaFM0B1i0B81nCf7dMFO1FTmEpj9Orzq5/vTe2FleaiyX+Hjg6Mbp
MPX7HFfQdaXxcbPCEBrODORLuZlWUkj8o80uoO++P6ZlZJZWh3iIFr/Na97VAkDv
Y+XetWZcAIVVAmkIhyUcrGXzMo1RduBm8hWZw6X6iyLZQifCXVFaJSvtZjspIjST
A8DY9wElM/ZqsFapDjCZePmqJ/JwLoQynzYYbs4bdz/XT/qsFIxpTBcaUFf1Fe1M
U6Wrb78Im0pyCadISZWkEFo1/FEET+FpBMM/u/JwPZY=
`protect END_PROTECTED
