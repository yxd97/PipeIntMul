`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZDwAA42l9zoY/q+qpp81k8qHfWJpWRr80702QnuoaySM33XCghZsNb0mpCF0Mzq
KkD/kv6GxHauLIvELtZu01bAPk7YJf0/dvDkFRulIFyeMvw3iz2v5nsHGRCGS++i
eORoQHrK8E5Xn5OZYJ84mYEDOrc8/r1N0zci07AXUVuxGwzCAz+txSE8pK75vVNn
E80Xm9tAlUtIwzuHUrpPBoaRb2wovRU/sst5Laqlq7etabRh2aUf5+TyvGrG4roa
sIAko3Nu/ZhqaRZNVBdjDmsZljQN6uW/ul/0GQoedhsYhNW06xQsX0Vt69A1ns8k
AtPRVaN3//bF6p+s0GSfHqIL3o95KiFgljWYVLiGJ60OAVLb93G9AvDIyjDfS8JT
uLjXRbRn1IK2tJRXAiv8nUxnou+FPCPth0euTpqOm/UT8zYfW0Zxw0uIwuEias3L
dQieFmspKa/vKEY9gDztu70Cfwp3O21nqZDf3Asl/10cs3aiuXitRThYF7rs1IHp
/6fjad4Q8ZOZVMD3tZSB20dzFMP4apaQbV9w5k3nugi4SKWLqDJ9yLXnpv+LkpL3
xbQNNUxZNMNN44KQ3TLBxWJMkI+o3s9AFt5EhDPyKbQBizPzGV0c2812DgOmypQD
RRlv6ovS0OKYzVsIKl+hAhD7ITBFOjmxlyVg+2eM7lfEZML26++Eb5PlYQGPvRhW
p9iCV08UJ9hguicjFafD8cSh0npLzI12xDXIffnGOD3WkTNVp7FyXNq+R0SNnsLo
maIrGvdmb3NbHLTYhb1P4fVGQnvZthwthGay8N9665UWPnH+Zczvb92cToyQ7bDf
z+fo64kCLUaKsTS3PxJIItcmJIrbtc9nc0Il1eJOmyys/zSRwSXD45B36DO4Sj1K
AXzDssEMTzGp5AeWAuiuGBXxU0WpR8Vb5jHKH83DPsKgV2PzB8/AtafXaKByuFJZ
RGFBH3SROV+6UBIifWGBdlAZVqKWB84yewcu6Z06nUJHjJpubKkVLXSES5Jq3aJE
LAn8rATJLqi44OkikNAVroZ2/Z1qQwv+hmLMxXrLT2uY9YJDzt2snfV7BMa8Mfbi
hGSxPIbF+2RRbzeHgwHmcQavqO67riCcE1pOS2HJ7+3J1QD8DedJwnZQM3X/fD1v
5Y3cgBQeGQLl0oaIAmZ88BYdosCxEe4FIZlCsO/tqjW6ewqN4j9fzaQvW8wzXA0/
ZWudAkfJFzkBhKrFSYc+HyIDsAr3U1c+fHPxK/VshdcPepMjc/DM4edEL0hrNDjW
UHEQWeb/ndympG7K6NHDkjFotyVe+xGQgsnCje96JpY4FGzA6zG6TDMBbx/ZJXv2
yK7ljJETbBKwR4JjjghrpHjNKWokCnuJG0cCBynnKxYVDeFGSKTrmJVEJfI/KrJq
7kAiJm9OJ5KD0MDvRuicBvhEP8l4rh70pB1t59zsXR+ma16ls7wZM1oiV67pcOGu
3/yW6X+EY1TTaucRlYbvjK4Us41dOhWyxOULqQSoxaYT1S7bz/jd40sttsWu8ltS
7kx4DccyP76bUU9jnunLcjyN0x53sPFLQ4dnxGILsozZzyKO2H87DdYJUEJFluq0
WpK30wy8CGup1u+asr7WizLCVfvNdL0HyxRFGaaQV000ansD065/eNc3XB0G/SPN
0XNBXayaNjILoOZszColbP5L/vUFbjkrQCnpThmrEF2Z8kstqyT0SN9tTm0BP+1D
ytG0Qqmv9U/Pzz6s+X5vAA==
`protect END_PROTECTED
