`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7MNkIHTOnw/i1/2i36WGbQARHshQH666hX6DXZtRarzly7aKNU/C0FDG1QXmrJPU
g/xj6lnq+Rp1YrfBL2zwVSvHqyrgA5q0M6rdZBUlhqBie5tt+1sQ1vSkF2DvZBVT
qn7ux3cQElFlnHFFOhIRrNyYdQMMG14w6HhA7N22eGXmX2QNvFP5k+yPTNOqNL3g
0G5TsE3ssuPGPsu/2EIwReuEdAXLrfJrckWuZM7EuOa3vMCwpuR0HLh5qou0GxaL
6eqbEmHJQ74AXK08lj0axQoJpSyV4LuHSDYKJTNE9EJl2w0pWppPCnoMdaXA41of
LAq9v4FFCnsE8pbMIsgtzaeEaOM4d7c9m28CZBePm3CIK9JTHS3kVdGWCC6SQ70c
FrGMKUpAb4IionjGfe91Y861AmSiMkwtxoGX8EX9X0YO2TWJ44xqX1DwNY3nacFl
y7cF2b1V3QJ3QiMGczLC+YBfLcTfmu6QVoplg/gMDOSvw6EdFxC9aIh4bLRguaC0
`protect END_PROTECTED
