`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/3bMEhAPyo7Ux209S94Onv/+kxh98+7T4F3ApBsNgLN6Wh4OyzdCoMbcBwF3R4h
R/VkZI2TgZuLCy/wuYBDe/evbytmh+Hf1FXKIIWFio3W3ShAOullPOYQ4Yidtms0
WHclyvAZXkWpvRh9ECdrFVIHX2g2Cf7K5xalmIIvlyGMcdCYdNQWNXS0whB0+9JG
/wZFRQoyrT+7w/aE7w/EzCBX4YJ/K4Q0IhNdn2DGPyWqfKjcWwD+awIZQd54I1Uc
9iby/lZYG5wYCr7O3WsbYRz3++4glFzOyvavDQIjfN9IS/+u9iy6gu6bpNWanj/5
/4Wkrnn5pa4u5akYpElODOcqEBOZhRf/JYOR8Hs/u6oZzQU7k6VyeePp90kzLrFy
0IFdXIpAdqFbsSSBFoXGgeFqQKHR2ajf4h7KxeZ2VjfwUmHqa3wziSGSrYC2BUHF
ZyJJVjsMizopJMFYbfqwAG3MP/PMMb1yUyNyqLiDuZxlZ3Ww5bccG/4PUI/Yfh1k
lPzwWIjuCzIC6ywQND0amU7TpuliacqytM6pyMcTMSs0Beybw6tgc/39lHOxC0Hm
PvQ7ilGuFhFI48LvS8Qmu3b1H0o4fWjlkMjDZBKDhL/Evg9PfnzbYvdryY9o4Ejt
P3RR0k1ne20zjiXewiZd9eLDuy20vK5T8Y7Tj/NwXn4nPB2QfPgumtzL7yNyCiWn
kZFA5N4PHfKQLu6gNjmyHI9AUymh08N82wGkLfyuDWw3SXL0g6vMcQ6Bjx0VzLfN
IC06CJZ8jU2P7T45Ma9WLpAS4NMg/bNtYVHdp2zfNQ13P1cYCMTAHWPSpNkEgY4u
Atli0KJ5hg8MENhFC+GknXUG9D+2yEWCy2cqPYvsPVg3D6PYVb+v5ZzIQZDvVU4H
ncuqDslXupJPQFy2K6GPmyJcQ9cx7HIlL9zR/P/lZ3PmweSYk3ZtpSi3frr7dM4a
Qx7b6/RbZRXuklFzFmpeQrzLJg1tI3DOHEBgZyiOYTINoMao45UsC5EMivDnPxTh
l1snIEkqINxMKcSlNeSSDO4mlk94Qr+/vrjTuspP7h+g7c2Vxm11Nh+j4NBhvrV7
ipagjoGGFvAARepn+HrzCeZg35uqmpSj+T4+AT6aWwz95jAMl+Zmkay9izCV/O6E
QF7nPMN0Xx+fDY0ywWo16IwOXTfa/WPjoDTjEPMs5vyZ71XUdFOi4JdZwG7yaEE/
n9IoxNZGhUxsp/6gUUh5zJ1139BCaT9uYgnOTvyz3ygwY4Y4p3wOFiklJLsbNIbD
`protect END_PROTECTED
