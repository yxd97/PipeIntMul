`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTIpfUdLL9sttxCXQixSifZ0B2sYzKqwdvtvhMQm6Hia9u74w2FJSNew11GuHrYC
IFJSfDBBioOBeGRnapdym4CQCGb88qvBLUZaQu5Up2v1BwWue67B/5I5oB5S9VuX
suAFubZYqS7k6AekaECICCgmUGHqAvFFA5myyiiNE4SNiFcOCII+MP8Cnlrz1CrP
O5RCEnk+06dy8EiJ4v4RvRBjyvKf+8VbM7mrVrBAlrxC2ljl9xR63gqYe4JnX/XQ
unXnP345x0ZZw5pH9GW/wrRCcJGQ2LdyVjcB3ur96dMmxnaTgT9xkPogM1+BuBtp
jtxCB5O2ibDfy/bVzFjulDbNqnHltHuVxWCtPqEiZgLe3DUNSL+3F5rjzspRdbsi
L/8ZyzXRCwDaMR9PPTXLhRr7S7qEplKOzLRZt9j0SZs42jMGJLqyWph9Zji4z1H1
cRnaIIvhH2vlbYyGirVc7kNy2gjCGbQ+yYgo6CT0CIF0jn7Fiq1ivHhwJes88aSR
aN330QIsr1hr4M+c6JwzTfDmg4GD8g4XHfjb1mopJwbRQoKrdQblraucaCBmwYcP
`protect END_PROTECTED
