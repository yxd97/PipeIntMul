`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7AavqitBdYoA/U6uXhFd6gsOeLg2Q8dHdAt1qzgTXk7kZI7dXl7YXdLkgLtobrI
OyYiC66at5ZD9+MZRHwTu6j5CTvqqgp4JH2/XDQ3MygOauX1A1fThmxFTD7Miju6
MWXiTlUDfjm7k7kJscFGG9H/t60Fm9U22qj3F6i5qKjVMemGe7oxi0MmIQ9mBL8X
+A5NixvZ9HUfWABvOie+Gzzw4+vG8oTHHzVQz9n5+XqQgRXF3UjkWJokUJiBVRHK
PSmDiL7lF8V5mvqngeEnhoJswgmnCPbPOOmJ9Sp1mRXq7TuekqRpg72na6LmFnFC
mG0gxKpECwg/3MBNF6IvKKE6bEiEaeRo3px2Oz5MiPsmtgb0wpiOQftdSShQmJ20
jFmIO5u9hSxMxorOo7aNgkDY/+qzIT+9inHQ3RhbQEl2NMuXw5S0tpKSMVYU98bu
5gTj9D6lWxztDsUpPunAhl4ecvGpF130p8t1zsbOFvUJcUfYhtxSY8pe/419IWJG
tp4jiBEhxbjHL+eJakm1ypyOv699WSuoWiLhqqOM5MBo86mTSmAq7EJSeDBrVkvS
p6S4/vOpqentHJh7L9fjNX5fskT48jelu/WLshWABrUML290mucbviB/PafIvLZK
Nr3X3YcEokYVqOnv++zU2PHXwiygU/FyAhaE0qas4owmrA+K93hc7xxw04NaPe5c
vSlvmhqmde7vkXyWSKGW2Q==
`protect END_PROTECTED
