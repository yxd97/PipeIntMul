`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/dtN/N1uYDwkmC74k4fx2UbFI1rIegHVyK2bKJV6mhjDA2kUp1oKXeTqoV5lMqj
M0nh70yPBfQEOKKiM4xyxwVpTM2+aZ+uI+GhSKXelclh6oMqiQgDG2H5AjQsNOyR
z6U1yHmZlSHP7H1DQiJ9SYQWlYJQx1Yp0HY9YZY96WemGk0+7DrRiOftvdzw5yW6
kuQFqktJn6DjcQimSPQc33L+H0hTxQO2+LFEYKzXNf6giCTmKqk44LcXx/RGOAyR
Ue3iQRBicYafHcng8+N/VDUIXg8ceth+4dHi9megUoMaj2whE0jOCS2jqNUNlQJx
ZxCaaMq3I3LdxVx4tCEFZwd1Yc3KTzVZnpevZlCG97NaofpWqY0GPSFl2fKHJPt/
lZ+ktbqvt7B6ZNbUwl8Nks5wVuPUNWCnFySAU/cDiLuyyTjl/s9pRY/zpAVbC7xd
6hrrfhMmyoHMsGApzgSqfSSp19NW44/5UmXD5mosmA8BpCKTpn/X7OybEeZJWOHC
Nr+fCih7VLvbahEB7JEcHQCVrM8DtXIK+vlKVb+teXnBHmW2u9PAOLdNwB1v1kk+
+1+xYQHW9x3s+ZYbMeX7MIStDLHD5c8BLyEhbPu4v1JjY7MfzCqp5hWaKdS50V1g
dDIdZIeJjY8fTYFPIq06YRgOr6kw3QEvUqZ2vRp98SrfuUgNidQ50addMkSksDQT
QbDJAnpe7qbZ+OVgvCf54rvfCONrHBOcMOEVPh8phr6RGjHV835inFtr05YviTiG
FrQFE9ZYgqOZivFljUiYsYU9h/Bq72MSHAGMuE0NhIqTXEsL0YWNtAOHfPdb7sWe
4l5FMpaZyoYqSqHLCCoTcLJkrKtqNoCrTG/ke7KgEWMhRZoMn/kxnbdacuUYDzXe
6vL9/rKLLSdEUKx+F2TTlpd1LvKk2FXgRsInJD66uw6DhbzazOfs9xpHBRp2MGJw
Ifv0erkcJQkb1WHMP5gKv9WUozh0VPGSoLXHEDNeswv2stSt1Ru4nwuDzRy0R6BB
Ac7YRjZKmnreQJw92nPGI2Gcq7yN3AF+zxHzA8Kj/apW4fi/Lk2hXL73ZrcZduvO
Z/anJBxoZExyCfim6ZCFE/9xdZI/fWrF09mrE1oAxY1ItXeJZSgAXClsuN/dpMoA
uanyss/vpAEapMLfb3235Qv4+lFtmEMCMmlIzl2xELb+eVAcz0nTwzyCVmkSTvz8
P/VQB/8a5brIkOj+h59kDwYSA2siUMNfGeL5b819Ba5lq/t8LnJTitYJOFD+Q0pP
mUc78nTiqhQEuQ6akP65QaIYashTeRl+o2tlrzrRPNvugMq/dRUuMs0en/R6Tzvg
aITg0hJ1vjHN3IHmEj/UFWV1MtXSCnyWm6IioPSakRKfidcVaP2nT0/IP5CkFDX9
AyLRQeDd6gQEAjpKHlZNyY7Nanx/rdiCw4K8mm4xGQmb4xIhE6DVYH/C82Tn9c65
lRVp8k4GWyK3MbdLEeL0STuGKWZcC1wLj5FVWRyxfIfYuGy9OeilnbpO4FzlUVp2
N3iJnzUjOInICAPRZnyi5ZpGwhAC4H+ZpEW0pv1o2TXQ+rGX7p6vdxqDWgHekVV+
H12Qo0J6yZscmWVK6Ls3565rN4s9G1X/NIW4dlUXWQSW+WUJyRXpVaolm/FCoFTF
QcFdBd/Q5MY8n2vGT/kEbVKBkU4Lt3cZ/Q6X9wJIRq41kiTs1SetcH1I3UFYrIQD
kfI2pSkmyQpUwR3cXVfRX0cWqd3lTActNsekMSqAUpsNZuNrVffj60vFNnB4+0m+
xph2CGkTRKPgV74ovw5DOEqJf74jxX+2UBt3f0Pvu80w+eXRtOypRJzRrvJxOvd7
z/9U4egmnpBuhfBBPchBTfbn72ZMk38Fdk6KpWdNqUCv99/pNIctO2jV9sz7l443
9rW79mjI0T/I2yy9G/TDa64/EU69PeRewNk/Ss2aeCQAwQqMK055PWll903kqBbN
xrWDkHGMN/p3MUZwt2XgU+fyLN5bNjMAheT25oTAdlJxewXo5v+8v/xfj0lC8b4A
Os7hkBLyfF0ZmGu8wOWKePnxmdWu/ihLcw89m73vxokiBje1i/csc4mtlEYNaAvi
vZmPqoKzrESl7YinvHo3KOoW2HAd6I6FvtbT9uUB+6tNeSrysBNwnYEwovqNePKJ
xUCZkPkjDUVProCwHs/nxYJIsc2nh0isHlVVj76AfRXKgS6eSPBaaDmX/BEV5FQ9
5YJat/1eaHxNJx5QmVACPsqrIhdyqET41NJG2GzssMdcPFWODkgopqC3vCiGUIpv
+XJgNE/9RFP6llf3KjaNrahcG815G39FJEINrauwlN2b8BnI9SBWMV8xCiaft4y6
WbUcBWXeXnYfwS8XB4SztA2jsROROc1qB+fcx2bNnSq0xbGdutgYr3fGoyDcMb9i
jbdKCsM/7d/ByWN7q61YRtH0NIMxx5l0n1vk4VW2Evaa4QvWAXa45nao4J2mnU7d
Vrc5f+MZsnqA82ynT18sijMW2ae7BtOznqJWQQZxGPHW9i7AZ8T2pLxoV5U6AWZs
Me6FoTowsNV2aNCY59pmt2059vk9Dcr791jV4DzP7HPb599h4OfUHb7gZOAMfJcZ
5JKqAOLffNml35JA5tZA2nJ4vANc5ASW3YOdHj+GxyIq1/SFAxeU8Otmxigrdm1y
PTkcyMJJHgnD54wLC+bYGDNRB/fpaS5mY5BQSYh16da+9sac0v2EbmXKTBEXJ+6y
+DbTJ5Q6IFF/v7eAblf8mBMywRAxix4TqkVtIBAur+f67O1RF9QPR4YV/DIs0D7t
ixcTMpKvx539rNt7OdZ0MnQZab0zdsmN9SUimZNIhBsEea8APq5kPvCQfMbDp1V8
BKb+dEfNMwqCk5fHEbh0tDCHfY5ialdXiJci9DBGElf/J+mgsGHa92aWd5as9aob
bpqvEWl2k8jAVxQhFjt3PUMDp8zj2rAqC/Xrcz9nbJnQCEnJoC+Y5KzwQVALlIPT
fRazgybzSXmb/3c1PNv+V+5vk4PclR3NdVPa1KBxO37mVy9CpjpBbXf/IByy/uv3
w4V2XKSHTLF4rskmedatWuLy28lKa9HSCWUDCc80agxubc3rXzUTaB0PLtRokO5k
rhvlr0ms+L/Vti3us/WzRyi3EJuL4Jgk9UwWVSuyF4lEk/5xV6+z9xj1GnEtXDwW
r/0GldAr+MvBZjaBN0/UQx3VgQaqJ+vpcGCKyJj7hFYtk/RDdB/Fjy8YGAA5veeG
C+IBmsNa7VpwwC3hMeW2UkKn444tCGzxjSZhEchcwIEzjxfVq/9oCBBtOO0Ym4sk
G/rg4GKE40ad/sJU0+/9KjFlk+uR1nkYXIUKAORmLb2ehky8cKqXiA09ZO9XjIJE
zCC2WTfqdTkC1XWs7YRK9lU7kyzkegrtyWfYU4gdalTgACnaadyWjwP5VGixAmV5
MD42keQgcR/83oTe0SEdaSONOOdMQjOwZki84k6+qMhilVlFwApunNsZLgxO6drd
/1eP9OatG7dEamStqcfKSSHi3nOsC2ljwLHbZmXUxEUOZ6mN36McZABO9RDJAlsF
wcTaTBfF5FinspJptYcKuectG2nZJhegf2IvUwhn7qQ9KKVRe8wGGzd+YcL3gz5V
cS+QprYrFlWj+Ap6ZD00GtOQrjokazBKmKBvGEk8Ix2aXKq9BrsyVE+QfpXA7TGb
wfkL+3qA5Kskv3devWApgQ1//KS/eNNMMd/i1o/ShVg+Yd+alPhHX9O+IHfwZ41f
LSHIMXxEMJgi7sb3yupccrnHRfxe0ObxePPwFAg2hQKUg/QtYyNPIb9XLnsCummO
Ya9c394Awi722yAx1nT7u6kMCgit61epI9rC2g8+5C2ZIjSqNG15tc1/E9D2V+Pk
N0jmL4Z3ni4njN6qKjqURpNIQ0rWrMq3V0nR2XFZaEcUtV9BbWqc4O9nxGO30a6r
W3816U1wkWzqbRdq7ID19uPgh3WwvF6RLjBX2FvN3yguOfLLcfrrx/RH2se257CH
G0tGnGbSCs8FVV4ueEltbYL4GyDic+34kIQg+bY/hP8/igBKlML9EWH1lFsmW1Bt
JU6GtQYDKgvQYK+Q907c+iuWTDIzE0cCHeG2K5rB/pINqcy18wfuT6KTl0PEhy/c
TUyKenCjW90nHC1mONztWr0FVGgvMfvDsklYV7avLDD976FBzEtAaiQcvWe+mVMT
gMiHFaMMiB5fx5ZjTLI6hgpEfUK67LkKz7SYb0qv7E/qRthwtsImRzRUhoh3fa3T
COkkHD+l8EV6XrWxv0RKXbzozydCn/D1rTL86dXamAAvKlDtyH9S8MOlY7mzuk+c
aBqMvsXEL5O6AeIsYYG5yYx3IENzq5Ix/3h71tbsEFZYUa5gngom6OfRFV5f4Jc7
BqPdY8KE+GfbxavCTtuqCU8jjvaROsXRM2EkysYwmgKc/kvJS/tptl0UBpAD2Q87
diWUdGzaad5U957IAPuiQd+ROfUkotZEsVjCvcxa0Whnd/nyFW0qYFoy998w+bDj
GUxUUMjw/FTTvqXFG+CaJdlBj9sKXOwDBaZd+MEbcSyESk2BmFKRNMG5BbrybqvI
qG/bZPV9VYgoxL0lN24h3UMYr2b4NkP3FVuJf8dLyxPWO2UWUasYFvMqjbilmrUY
Tk+KaSwzDiDCBPOS26MKR/xhC2hSpiZNnRX5jZXWzYrLtj3j07jt3QjMkAQ33ZHK
0eQtoXsMD6HHr5lrTfhT0i0wZavb2C/KaGKVEjg+a5ZVmxgAwnmewKPh5+8qMFny
P0AbpIPpKvPrwKydaSmgDQHZDMP2akt8jDcOlvSk8Mm/llRuu2E9a0VWiguZDKmT
GuxPcurDDG7k79r5cNv+HBVtvn5N8pBHNVrAtkHMAWNYDxglqD8zTXGvsrCqIQvM
UzndcjCWWcKIUdXIgpDqA/8qKYew5CD7ucGg/CRWretgGbAATli6IyhkNye1kGEH
b3LnPW3QSyBYm5/++0WBi5utDSN1CCQJlx8ca3pT+AB6fMqnon+CeiGaoNwl7Els
lvdAiW2KvupgJfzj9SjTJb2EsVFpVY96uFcvER4p0dEHwJ/57LA9l99s+nbuHeY/
9yVfpb4f4Go2Iq5urCsuurlVK4bIdhvJC7PyMNwJdXfBwhl5/J0YDdAUKseJWGWy
d9d56AjsDjuSWIaNcsyU9r4sAnfR3cfR+/6EAawrbtvI6UlM5zKwoBGU3DhEYni6
/M06fnBgksZdJQ/AeOrNGtTOgBVUH2GMlr7v1eqh0Xfg+o15f4Ls15Wjh8BbwdAM
gyGj4Q9kWDkDuxk7oGugnHjp/lIu9+U5RYOAoZupMJ5RtNz8Oiz8lY6CTdYZs3GT
DqQxrd/cMESD+k1Bfv81CEFQgHUuMnkRxgRz37FSPVlKdHy4MqojbvI6upq40/6V
vWVWt5lpwj72yuWYCmu1F9GGvqtmad00aggege/7ANpdpGeCvv52zJHEX/jRuCWj
fOmUu6z78BdEPRcB9kEoW51G/7j+DbZEcg4il0UcO5rxFrAUO908Gw6Mt1pmsZe/
6jwofiuy3H+vgKa36ECOm/B5gSjn66PB0tW7oowbaflW9zzyPuPMdaGXJGP0KzLu
LRY2+xFIgLyisDTAtaV3YsdFJ3eIiCeNrnktQL1Y2clkOuT+Yr6py+e98BhXWmxS
C9HAQXs0oFhrlMb8kDVqUij/7VwV4ZwSUWsI6hCqllnsizBZ7hv2EnrYrI5bA83A
RceBFJGH7PLbbYt9ztZjGVipkRq/Xq/yQ4tnh8iNy/gdQZL/WotYWYY6vEkCotq6
ZmuDrlSYuQpYp9y78iLsc84ryRR1zu/iv1cqSUlz8+8twDYrHY2UshsW6CdjVexF
BhGIUJUcpJn3VRHsTe25RnSUsYgyEa2Yx+v/YVYPaiENJgHZOn4rti+Dt0cY2WYo
1K9kX7M2LcZ24j/qdCzbQa8mPPRXe8z976paGZRM5TuZPNZBrWYGUJ4NS5k6hUNi
Lf1jmNo+eIpfcpQOwnEWlUAjuesvnnt7wH4zO50+lm9l+Z9yVBEjaDrNcALxWPz/
RL5k34OFE3daJ+nhqV7jEQ0vGGDhfVCeuV0tfi5CEuiJAR6N/yhX8CO8srgI5RgN
wxAgBGoZ+YZwzfrqDCpCMpipxBZjaiq/7wbgJGiGXqxlqVfLbtGVEAPK1MzjEla2
e9jZvKw+Kur1HxyIYdDywzb3WaebMGFuv2U8RI3fQVPhSlQ4ybDcbvdyniR0Ej1A
+99ARJVpw706c49QAGImUGy2ojfMhB7nLHNW3InSi1pjeAyw1ypC7c35W/3Waw9Q
PgYUuOC6cTXdvhhDw9T/dr7MSG18zlM/5ws9QEAF1ryQBpGffP/Z3BiWuUgPLGt2
Tp+dNb2+f+G9rEeLCMYZBJorF30r9i+5Ggj2zrZnObYcOXB6kmKrFDHa5UUPc/TQ
Zd39dvF0AxyYocCnLZGko7pjo8hqySpAPT2c4u6IB+pmRzoGGVxRm3gozN1GdWEy
xIPVWU3D9yYyqODxsleyzL9LmyzMyChfFgLPbqBlmn7vSFWy0Yzai7/AEtUijeqJ
a6WbwDjyhOb+l2p5Y97abZ64n7hFBNDjV1CqiZviEWj0qa8jUvGbafrhsJt8J58Q
cZ8ymbd/7ySLhJr0A2VskB/jknGejGBZ60fmd0tE32EaEAn+4A+gnaxKcKrv0G5W
OZmToIyd6mMCtFynXq+OzIgsOoqyPqsr5I6VJrs+RshuoQbEPY7zPfnlkTfDU5gR
BE1LcwX3uEu3MrMWLBgprRtG3qAlSKg7ganIwbyh31khehB0gDk4WM/ewh3L9maA
Ayy61x6g4v3Ui7P+j/V+uo1lXgouguDxD19wMtgP5GVjyM70mUsovzblf6QAhOOS
vj09vGcOJHN/XlJsbwfxpdjZ/dcZKaC334ClRHjcTuzqBmv5SvmPxFCMawsvg8s3
FyY6Pe5R76cezBW/5COtMKKC5TegThx1I7agWmr20lxzMEXTBN0TfUoRNKBscZLF
TuZ4TaWVUlLVDYaMh7v7hNUcR7eoyugzLzzK5cTYmQr9fLTC/W44aThGfcMR5fmG
EWw37K0LVPGXLY1Kv832t2SCdRT7HLRyk9xIYlro5AkCE+Td0q+rWbbWtO5ogGhm
f9NVehrQx2KOSD1wxWWLieI5ESYlIeAfzPY4ie/r08L8bowwczqS0GpqBwfvtNGf
UiC4DC0SvDQt8K7o0eXG1PnLucCXhfzUm32OAM/QHI1rz97iAvgy4U0l6DefCsqy
xaIGtn9ISReor5zBjkd1/Aer+ViE9nAIaiKlg4C+t4wlfmmq8upmm9eclW5kHiht
7brmEVssnvaqyrPKftMLCZ3PYGWL/BrBbJsFo2RDCzYop0meKTklwid0A9zaekNk
Zu1PHRDUe6ATLWwS+fUsmKE0456iN4ruSn/SL8+SQ2d+Xsa3Y6o7i8laVL2z19Lq
dCySGZZ8Cs6GykHOfN/l25EJexK5ieHldt0QPJdr3WLVuv6DhAdooaR7AscH3QrY
fFeMOvNpmqiZmKA8kFCzHkdYPos37nRh3/uxrjUhmDcnLLlqHa0eep19E5/GtSSg
GaADLPdPVlr+nIHdiQC02YiR1dwhwV7sVnTNcq+shhtFiR0FO0GhNMiVNR2fLOyo
G9jT9CuT7iZiAKVZmZ/L4NoejNkfUuCZrXa0TSC0jyRvV2o8/RzghwIuED3GQAdU
F688BnB8P2EmupmWM6AKaVavIL6mx01gLO6GNmJthR1cP/M7EOa/qUx5wOxgQbqC
u75tHlErdD7A1DIIpglsIoJApTTfC+Us9gZpduTmqzJ05AwI+dCNwr2wJPXqBFTP
e28qYh/cflIp9bs7Ko3IJffU33RTgEAbTZ/N7mL78BztIr3rUohELGV3JviLVYo6
+a66ufL/RlfxAvivuFOGn6j1CTs3xqIszgXYocgjAYyqusZqcc24Gxmtv1BR2puf
ELTGbX5PQhQUO/LswalhaRaXbNCyBM5fYEV0D3bUqqXXYR2L9q743qaFICB0KKVn
n34l3LRhHXPARdfynTaT8Wdfd0FmewV/bllWzSAnyD+FSLQ5MK1Z6IZDiPT10kGH
uQa4Cl/P1J/28V16GsfbX8v2bszYIWY/1U+sL0h8zH9nC3j0LL2SJbBgsO4CAuzM
ePsaypclRBWgzPJ0O6D+AyY2fxgKl+tXn4oSs1TpmxU+Yi5i84MmIJHDUrzf+55P
JlAOsgrG0lwUOJSnTEPKwvqYiozGjCwbNIJ8yPKpwWzuFQ101KSieqd+oWiqYSz+
jdnDJLgQJhEPCqaqcAgbMOuthVVoPJKy2rZQ6OhOz7CRH/6+7881C1FaeKbZA4V6
n0WrBeKaASjvBiQa4xSXjarSXTHNkOgt5xBXtY91yWXD4+otUvcA5C7Pw07fMLeL
O5LxtFMBe8b0bae5hlhFC2h+vtfdcJk9oqpRdE//4ECSSkFS5amvFgSaqwJCo9GL
3sAfaSGmLy2W8z1ZWU3J1v852hNj0CvR7yuIMgwqcHlGjy+G/S0luFEeOYlfw7Zk
WQixz09/tqImQgdBtMbDP2AnQSqFT6H7UjdSOcr0H8w8dmb5iBbimp8SmYkZy4Xa
UC3rr1mIreb2i1JkYJE/Xd5qIquuuydWMhoAz7kfEU/qxOvgbbJXlsoCkxQ0h/82
vchMZN5rv12sYAo7tqcThvRPD36QRDTDdSPydk0xFSo/lKoiFYeYqzS9WaM+OPtU
uMTKhINe9XRd2BdnfpqHJ6ST4EuJkRXSss/IzmzYYS8YRLj3EKn1J1N6KajAxYeY
CxlcX5FVLtV1GdkfholWQN68yvzwxzbEhKllha9xu+l8JO9yQiS6+GmNJiClbVEt
rpwH01anUD58CKO5Xem8eBwt6+yxe9Osfa0QMZeVHm6LnNBMbwWwEcDNk6IuQ9r0
j3Bakl/pqh/c9ZGWKQ+vfhegAduHiXkK9b1Z3yWNl5PEzDTSreKuZHMfIvNgq93z
naTs6Tjpq9NWtCR7krFWB3LD99RjO134/qutbwoRumU1hRVN1gm9IeFwHrLV6mPo
vLrmcC4y9f7qlYrYG/wnp4KdMxeJ5C6DI5lVHXN0lkJ3aHUKXL4PIHOv150nhV5t
XLpoyPlYpv8wms05GmohV2qYeGiGIrZxpcJYYtGmc6hns4cXAYr+9N32hTPJ3vJe
g+ZCUX/0MBvkp7uba8f5fTbXFt8OojGt4TqftYUx/czxDixtOBr+FobpBwWbAVzj
O2TVRQyHoFoGbZxb01S9r+Jsx5z+9dHTBLHbXwKAoMnq0xtSGi39sxR4dYAESubF
T/+FldkASvbyvAUb10m+b5GbHri8J6zy4iips4LiXtaYociK0PDth+KQETg88Gqx
1xaaU9lR1iynv3RydxAfwyLNiqcmqX0ndBeCD/4PBdZbGYAATXXZ/JLDQuNH5jwg
PjQJH+n08Waoch/xWVGKqoCGzkPLyfqw6VC02czWjbCPBE3xBQml0EfJ2+1Aw3em
SpXCnd8ac6/jW+p/o65/rNwVdp5/ce39yFHVp6a3KZRiVXNWpA2MvVgFSF/NzF6O
sV3186TfLSNxVzqY1RbK61GM6+Js2fufADmCV9y4Z/yxNqgpw30c3HSbF2Ylh2MJ
eRda0SJreHJFzpoRFT4Vjy/JLEMbejcUInU/FwPPbXvi2lRwzBGFrLrCDKpG6w88
Wrgw1zNQ707WoqC9vKNSEwLxkazSSP2ZHFMBkWcaFWJux0sXoosXghbEURADjP1q
H906iu7MvpvYIePWDH572mx6RzP+hjFwX/g1eJxitmfRapoIy3CeJQxLQcY8MUdH
Uo0pxF3IjfwHEr6kZKRjNRRmeQsno8hPxtrJ4SNAWJafDNMd87H6ZB0ZlP1Pxfyz
RQumPRFE3gFwWT+Gh5Xm0+JQEJErqXzEG49m6iP1vRvI/3Ik0z4viJ02Y0oFsvor
E15yrUBcmAql6qGrX29dqTPEhOc7szM/92UgYqxeC/DXKx1HPwLpNoc3Vj3I+zHQ
AP3Qq7qW4I7gjNItz96z9QOIi5Njkg06B6aG9peyKlYi7A6qeECYBjn2FSTaNGWe
qavOqBZuPLkkhBWDA+jq13Fj8HegQHeUcW62EKPt2uC0e2v/UOooUp6EJFCn3R9a
7RJO5FkV1KfkTrQFJOWS8oJV2yL3rfWoB9UhURyg/IFUnQeldhzVOJWSAb4yoW43
LRKU28lNO7+e4JcDmgKSjIPzXKmtAge4yISvWty5+zp8x2CWdI/GPqm1vWUKb6RL
0HrL9pVpiTc3YPyQHSzaZvQe43TfFnpg9XkiGBKzsK4S5a2EN2UKVXbl+xEaDHnq
o8qRbAX2fP6v3LrT3HRl8TuUNDOqpXvlD/T+WJ1DLqnTWIDZy66gaDN+gAUWkOYn
+xJptuyG/Mkicj1ca+cGY4U7c8lDlefKzFSIffMRngzPHpYFTLozrjZLihGaNNdP
K2+GbDanEOivquR7bEMe+bdHoFdt5Sy6v7n96WtHofId7gAjkUtQgL8R2W3BV3Za
IeSrvAfXXzejXDGXxhhA5Ifl1VaJFOw7YxpxRWloVQfPN63vO6NCMiJERMYWZF9k
nIftjrDyg/NACqq6Zaz4oTmr86cUvcLKn0dp/W/zTzlELJfQ+ceg6YTQhuPB9swf
1e65icCl4KxlMQOaDwcEtNoduDLH5Cyuao5c2OtIsZWsvhCQzSAV2zhOmDOV4Rp4
JRmB2PZgHkuF7XuRGqT+uDI8VxqWWv/W0Dnp6uUFa8g37V07xxaFYy4PGYC83Uyx
a6rmlGjutRfroTXxL8f4SQUkqDmOW1KzK5HIVS5FEOAma9K06x4tiF3sHdnkSDAJ
dSiSggMoyCTlqPDavVevurTH3BeG7Bbvqi/2rzhpjXX7jD5nYPvM5sw7ydA1PkEC
8H3NPun35v0ckl1dDtEvFCVIA9baHqWqIPmkTzCVnarb8z19RB6XY0x4qux7wFrK
BLgQkqIzdjXVOTBcZF6wDEf/FhN8mSMuznIWedYllf7EUrPAFnHJ2nU/prsbcOl6
O4fZRgDCWR67dap67IFybAeT/3IalRJl61+ruOO1+jZ1sVqZ1FdV4pXNd7+yTsYW
Ur6Ss+FMrgmjn8ZdtgM+sWHcvaL8jzv2llYLA+I19Nk8+q3mR5O53vf9kDnW0PwC
/0UVwjsehBLrk9EUnrAqC7GE81JnzbrE0uIlbhUyamxgEVaFK7+Hq17nMwjRL/b8
e8h69yd01hJHEgqzZE8Sm60mhc0ec+s4AjPS7ve91aJ11EH8yVmUufTKjeNEl4IN
rGBpAVA8xq0JseeKfJ9j4iLXgqlikOHan+n7D/hwbeizTGnfjQn/gSKOUy6Ls3v4
WBrNAYpJZqFkV0Un+fG87q77ly1Mm/v1XBRva3w0wtIw1QzTcZOcksMcc/YEOIwf
rtC9czIZzmPLlFJHfYU+qJPnqsGLLoLNvVoH/pDfZ51VvRM9+qJhIywUYzhJPBKX
dlcITq3gXBrANlcDAL56FXkJOBYptZNr82OcgjNVwGlmlF49tij4ZS6hviH1tH7b
khqusD4En8wVSp3+VragMj1hbybSX67nNTke+BVTnoU7RzCyJzaFbPxxHA6k2OPq
rmDs0QaMXYU/8X5EH+s1DjsygA3aae3GIL3EpT/4OYmcy4USHVmDMlPLxByeHwPX
tS+s9c3ASZCUE10OLRWD3SfbXTLSGhTMBVi9JLefC/OIp2w9+2CyQm8H9CQVAEgt
QBd+XfKMy/YxkEaA6dk8vKzfuDRmvFdsY9awtsT7v8UKkIWu33nqpHFT8oYBnwFa
6npZJ/iKDB7RJIvqNZ4+bkP2KftLpfR9YPy1+c56VEqC37EsoVTyp8QzkHXfxGBs
Eb61VzyJ54wjtqR/nMloRIiAn0WxKGLp761FhQUp4XPUMtiYp7TpdRcF6oneAwgU
mtEgm5pTOJ0kw3Uytk421S0ibvd9uJgWx1zjAif/thJ/ItBhlrCZv5DLlMiztGzx
j3A4XBoFAq6rZAogkyexFGLNY/ytWMsPl7xjgB+ncXVAI8g8jUaaxIF6TpnMAB00
1CT9u4l45SBJK+DzOXxJfWMOSwP5ZrD8GaMjJ5i91M7pdz5J5akkVTARqU504AA0
lARdRjkDdckhJqPv7rQjmK6zrOIaeI5fxUa+9KsMbvJxMIGbQRqjFRZ7CyzUp6m3
dnGsMrIF8+XIut/1bacKSIe35Y/X+nl2daih/PHhU9g3PRrri37CxPoN43VLcWfs
96OVJNdWWLU/Vle55TK9hIG/XKjl3dkRzSpJKOVuQaVZZCeLdmvdti5KbjihjMbu
GmNwhgk7MUIUg5pBDwobrYMfIaQn/iEXggggOwDnSk+ENA/pPjiJtY/3hmrL/rvU
NgqfMg+Uo5lZrDk1IbwWZ5hr4ebZ5SI24oJYcuiEAbi9uWvtu/yZg5lip2UKgtVv
kczNr8SFPhaE1sYl495Gi32ApUPqHYzSEJSXx01JUjmLYjbtPzjJksBzvStADSo+
d8JoI02HC7I1BSZaMqGQuU14uOUf1G9IuuTllv8XLxClpp1gl7ZHU/N2pSwH4Oq7
BU1/ff9b3U37/3JeB8QNxcVvwoGwXBLkLeG2y5EZv2cZZyFOwaryx9QH6HFUl4Lf
JGm9gIPxw9gE3D69OGv1/tit5QalR1clf9+VGv5jMD/HWYcWzlrvr7yzyTxuXqDs
zHnhhfd5GDuTNEgrkOaWlpW5Mmvd8mJDT1EuwYW46fsFtegddvUvX36c9P+C/v+1
SfJWgf1E8WYQWr338mc2R85u7mzwDzq/UZJWn3nx2udIdYAeW/iG77WZhCSfqONg
pILABZe3TaKe4OGlnAiwaEFOsykXCPAjs6juIE5cM9wsSIm4fMm5xVfZMKxqw2SD
FnfBdHx8gbBDDK9hqvDbRTL2ewgoTCxuoAwsj9vCnH2V3hjqeR9BR9ek385zusOn
bO1P/pCFS/HVvwgGNUD85km0v25da7pfQgNS+Si3a7130eIfOaH7jzQY4GtXBesX
U0Q3JA1iaftNg/BlQXvq5Yb+Vv42XxygG5kUyur8qdfpUgQTkoM4wpGYIEfMQFa0
g4dgdjgW/V4eS/nTgINB0aEuZkwbOpB/RI9PtpREWpRyo0couG8KDlCQyiIvy/xb
VBukO1IO7d9CtpgNrsMyv4rjTPZPkMCaAG52ZO3D35x/sP1RsiACE5vTwrmrYelu
6a0lbkLpIm94sNAqY5XkVlcFMcSgDv9b6agUT8DZjsiXDnRJlkrHekWa5F5MkCk0
5laz2y5NdQDVlKWrLqGJZ41mkruLRRB89amDjjWPTYAu9rDIfOr6S57DsT8ynQxu
e/VJ+qazMNmW9BkgBMsD3qgYBW7gJMnoYuafds3N7qIVGIoo5Ocu2FlNshTV1zGw
0hD9dY+joF+Q74optRfa7WG0fv2S5YRtSEFMbx2aCyGZK6ynIqoIvB7UQwQlTBki
/3HEsVonTmtBSTchOFfRe7SgN+ChAiInywWIevP+DHboxAfFP5vRPogFLUAmZrSy
KehTiZ4GfGGlXNvYE7pre4wLmLWCNjDK6g6+AeNjWvgR5o6/S9ZeLx8ktnJyS8DX
iEDWZZPjc3SWvQ3noOs1bHyeA2Paw+dFwa0VBg5dTiBi4gqKfrs35LGPmTh9iyAv
uQYpbptntcSxlfnWcF2m3fMaO8ZMOIVYJRHdWlqm9AIdDC7MJjrxveAe9SZ7RgrT
fx1YI2bqWDXbHB5Y0UlHPFla3BwXTjIaXVjk/M7pTzQbWlHnjEjDjMwez6elMO8m
yqO3vCK7vNVL/R3lR/ws+iX3W0CndIxsj5BbHwegPYA3Ek9D+XxTXZVEfOMbWPUA
BbNLEmvu2wNy8o8o58dhrMVhmhJSZOxXFW5IfKFOjauSyOIiC2psUsKDLSLlvjDc
BVd+sp3oQi+DcLnqb/YPc67/YlQgSWiRuY7dakMblEewWmtfXDec0GfI2OZ3oVCZ
q5lFhJ2ZQVccFJBn1xbMNi0VqOgJbNhJ3NUpwVlZP6KqfyDaQhlCnVQ3eTayx9ta
m01RbEqzipKmWgKsAeAZWgP4YLg10YawUjU4hX8r0vXJDusi43urq7HIQqiWWJO6
nYqM2dYTV3phBuuQ89Kh2Co8NJjdwkfi5o++SNkYrpH+tk3WRhlMals8pbv8ourx
Xmv0X0tsVr/FoSDtEss4wu0xaTOhBVyJXLETkt+WSSWlWRsWcXE/hQeTRh9lM8s0
Az19fBch2UmjNFG2XTQe3JAfPQvsqX3BNByCi5VN/tbawXHhus422M4z5kL8YWTk
Ifl/imaoTpSzwnGLY+YGPk35ZsTdxZvAhca+w4enb/7zvYXiew22q0lU8rvV+hzW
H5BOmfNnmLY+Prd2YM+rleQaITd6e4lLNswTwtXi9nArYnjEfIMXql/ut1yj3sD0
7Em8ty2/qNuzCXm9mRjJ3KAd8DUgfuXTXLU2ugQemSFzArnKmNFYXk/TQyPBNysf
hHfG9OfkbvJQ+Um0ebXdg+WB3ks0B8+klq8u1MNXvkMWtjwDFFwkxWf+wpsQTKMb
Ov1xyu2QFkvN3iDiRoOvfuzxBXeEW73epqRBNsqwKA6OWC3Fko8wrSg/HhsExsXM
bRsRCuQTc5qextB3fIcgDXHmUvXRcLGi3bdeK25eUsO2IoUFzboBVSkn47cWNFFI
AcJzKO5BYyGWw496gJ/Tu2/OlqrejkrTimdzFYfEoKMQf75RUDNFVi+r9EdvjJlm
k8cxhdOqy9CGp67s3Fehe24tJ9A8BBgizIbpkcqn1RZR4NgzpopBy5VY9qPwtQx2
cMIRIifzJ2p1kOX13/z3VBVuozHteIEtrvgy73SlpRGVpFosXumei3ZZqfUhxHT8
pUdqdjq99Fux28DeK482NH4AahV7lv2MVcK0TJO1/Av27CexAQ2Gi5aTSd2kldq+
wF+yd1ly0SRHiVq/quiWdgO89dlpphF0K2PaO/ahU9HQGdJuW3eO5tOtwZt39kUA
EJwWJzc2w3Sjm41RNfhxUu218qJSQySCrK2WYO+cUPJtnmLlZQl+QV75e8zWtXc1
gROa5+ExZkBT83MNEyrCffCMkMBuzvGrMHYgk3+/36FxRBVwmhwyC2UtRrqkh6wT
CJVMJnEoZf2Le56XAWcujBTMja6R16zktSEmAaa/sat/WaqS4n48H82TDhL7Ed8I
XOHqMQPCd0lOF8wwqCkBHokpHDrUGgSdHh7MMtSpiOrMdaUuomkWgAdZHwFKFWgN
XRJwysvJf08+i8Q2+mc/LDbEbD+220ft8jN3RIfPoObBoG8qQbNG9HVeMMnVPLv5
rUFJhk+NgbhqMEVffscmBIDMakC3VmxieF6CQbmuWKHzezg83oBlKYVmiproFol5
CDCryrq41t2lGcygFhFSgP/tNeSzc4UI7M3S5vVlxw6QbChAwGPMo7nZiPy/G3CP
n9pnT3440TOAtMiJl05wbFx45AYRjJ5wN/sJGu8KTyC15Cr8FOBIJSEtdKrv5p1y
o9OwmA9u4ftlcj3Ql8MN8hpgN2m0Hu3X9m3MZZZe/yHUlWe/oLRheBAj0pEI/UD7
ZFne8Osnzbf2gVRjYi9KqDxBxB9EAeiBubMC2uoOG9LMy6LP1+2yDY4fE8hDGD1l
L7x1VPsguoTUlvQpaeHo6hfFlJmUxWe7Q30v+yNfR0xwWVkMg/6Z/a+DQV9KzXrY
J6m9MwyN/veGmxfFXyHwHFwumLMzGJtf0Tw2eID/D3eEGIifx9/iYOSV7HBQIpiJ
LSmVCDkV9JEycH88ka+ZFpQyv71rRUmrUGBiYfLh/0MMMFxzGBGA18NCrrT+2gkx
v/TQpG+sJqmmEKH25ziTCR7x1tKkvnFxbLQcag0vZQjQw24KB5TJaaIKbtgKLtp5
nqek2QewUzlaOsTl8dYPgFhyDzIDASho6sHKVxXqOkmR7mz8myvkj64mlzY//rys
IYpwMT1hWj1Lz+pyB45BFb4oJYYzK6ssrClg23TO40JVt9CaRVSFNXrRye8JM4ed
rso7UULqCuM0jyaCQZSCOvaLf4t9JVLAsHFyt8mV64R6c1KlVS2HC8wuXcftV7bf
Ajs8ea12KcVxFZtBmr1nMK10LN37qEiVVNFfDMwAeb+5mbT0qPzoL/AQRyN13Rsj
FsG0NEGEOf0wBrskz+g4BY3U0y3RwtD/QBQsWAfoWULx0qmcMWpYKATEgaM8ZU4/
lG4FrvNUkVMKMdPhQT+AidTdkP9tcE5kYd+ltxs9EWQo0Yy9c9/68flFn627MmDr
iVOoumItwAozymBYFdYODZduiks4W7S25EcCtNbOTjg1inHw3AAdpm7em71kCIMz
ocKypghUBzhbK1zKAvw5FKoGXWz3qvbZ6Fi8vQYpZPedyqI8aCoimVp6ZhE9Uypi
+MXhbdSemB0kQfp/UEeTcB82M3/qr/bptZAaacxgTggZKri52D2/v1BkWBCFb/Z7
1IHPDys6IDr6onXHObLjNSrSF+y9Vq+8UKuG4wXhKZJ4D2RkZuCFOwFAAvQtcYjz
lLkqju1fRl+zMp1Ehh4806pbA7saCWIIegaV7yLr5ei/h3gIvtHH+pCz2C8OXqBp
nvBgN97RaMCDt3r2pCKDPT6qBZhcnS40U1ZhxmC/sVMYWXEZShXWhu8VDD93dBdA
Z3NZ/ur8SraVPDMfgcU+cTnG8sNV2IXzjvna1edQNzQAbPjkNn+cwVwQDR12CRMY
TzPWqKtntrbKxIn+yR4EqgQYB9wusFZIb7SxOxHWFVTWnqPLrGgpn3urm/SphwR9
WHAMLVIsBkXEZip9R5EtlZ/ApPCSrJiI1ooeOhYsttcX43w+aQwtolKrUO73UrSI
7dgHhYjizMtozJ4L/0IaJoZmR3E+AxzwSri9HJDPxIFJoXXUSVczsFNRk6bv7u0U
lRjuyGHgCarxBb9l2+3voezCbFob47cmXW9c/2y6poHmiSCtcbI26KDgm2wiBWv3
7yUMDrXLnNaZ3i3oXzDmGDUZ0poPZk9H6YMSGCSdgWlvYe35DfgklZ0R0C1wdIdb
mNE7TsyFHuGLQ+Z25CLBJFYSSpSvnZvzHSzPep32LLK5VdbNNlxk22t+vpkk8k6k
hrJfGMI+tny0aWq7fHuN5DqXibupRicI3fBIGotYdQG8c6PGNlLvA8vpxEjib8g8
4J4ss2EI0WQPOZ4WhEo79dib4gaN5NH1GeM3o+yXrNGiAA2rbuYPfh2CFqITUyMh
m+YQ30VvcJpYedQ+GlTedDBfVPXWpbItfX4U1N/NqcZE/Ew4SUXoSGBi2POOeQSs
Dnpp/Y/xdVXR1epqQNcVa7jp1xijP/0l2viw+tqYCmrldVRr08Rf/bNbwRBvyaMA
zGfzPIhKzkI0sNBpjpTWwq1vi8cQbicVuMEnUyHxz4ky+bEPk5uL9xc9wp5ZyRzW
sg5LYx75ymleOKg7oXYLZA/gHqa1FnKq0B4cCWAazxQ12nLA5cb57IprEywb9zKO
DnouVkugi6345IFFzOB6AcurthM6tN5Jt1EWYA/Sx/NyiguWrm0zbym2qsWG7ZYr
1XAnEoVS3YMy88Q6nNbkpD9UVynOobGQswyOnWPxLj9F46GhCCvSj8MaXAGMWzwy
vU9wNDhYr6h3yIw/v6mfrsENJPEpaCWcm96kBv55C29rgwkAS3LoYSfVR5M1my/z
+Mo/c+G6Zmroqg5WhiTqAQktg5qTR5br8A5nG9jLjKfCpjyDLQcZqMRTAG/lnWvE
tHHiEBys2drp3UkKFyJbx3mx8O6ZCRZ9bz+B0MM0/+1B3zH7XRYC5kHgrdHc4h1z
fgVrwj7AwP/88xpfz2PzIFrcSg1U6n7O9tJyDfLbLQ8QuI4byxLDKyAI9WjUsoMb
uISjeYvyh/oc2vLZsqNNBidLj78+rQSMeFRjNV8euBb4h1V4o3Q9h3QN8jB+3BNV
0dsPodi8+f2svcv7JMAvO6YyKfavb6a2dlIR5T6kKlqE6EoVTxDrAHqK6bGQeEYH
etl8CKajw6XtP5jE+yckkh2tnL0hmvrGdN05FG6kbfsc+ObXYRco2iCZlbKIWVes
evRqH/1m+LpQXwBt0m2WGhd/75JAWxU8Gw7STY0lyXhdcnSzQGKJ/SrTh5YeLIKd
dpA/QDCIvVI2hS35sHKgdZTgEi0D+A+iSRJQqQVJefdiZjFjiMA71a2ot8Ips8ou
zBU29bd5hibfvjWoKhxdM0qhR1MJ+LlMfdb5slDRXMmhkMw6/oqGqFV5cO69vfBt
AE6eVSS50ZzQlxC5FyL5dzGGiX9JGkiVrB2L5kMJ8K3LIsA5xPqIR4kJbd3uf1JZ
i01U+0XfggAWcQAoSPwMraVYOdgnU3C6/8XUgPlmg9uC3KZrUgsyxqi8NLU561aT
CuGcM+xRrNFOYjkT5WfxgLD0ARd0l0s01HsM+iZsU4TyYGh3iJGGikXACT84CJIY
F4AtnGvwpaFpcfoMfZ255UQKwQUznqbfdlQ4Ezffx5hcv6sr2ny7fdbeoWF8++Xu
BJjtPDMeEAeejBy2A+Go6/IEpY0N+MYhDc4DOIiTVy0fw3i6xXHuWRsPehRBOKE7
c3wUM3MmaFXCvZBIXuxsN2HL+eGecPCklNphZINFTEtm/lx33+CmYZASEGXzHe/c
r59puWOdXuZ3GRUJRZOFWyemW4Mqk7ktkOEb/OX53n83s7O2L92scF02clvxvvwc
Ep9LjH2EnzCp5WCS3IkxJ6khie01IxjD+AvM5y657jmwKMH0C3KN+j/lG0lYq3gl
Kh+CIs5uP5eUQ+ceC0edQeN1AOC+pd8vX3tt8O/tLBjrAWSILqfi7YOTYWM0r+IB
NLI2LXlqiYfUBfTwWzUOYNegMZrpZMd+rnFCImRr3gktyntuEv2czqbMi1HNLw5K
DfXLcrM77O09A92ZSJNoG7nTHTfFSYyFq1y8Q3jgjYPvmfxSPYYBHKwFTcu0ZjjV
xd0DJZrdpvrxw/ouyou93YU4oqm3wFBFCr2YKP0+malViUCJ9NUcvTormT6o0cYj
3CRL1Zp2IvdmPwaoFysV6f+wY9qQ1S4rnOyN4WTf29/D2xj6MXDSlemVkf95Qo/n
I4J8d8PR2QaoEvFFdslirxk68JhXOx+cv7t7uUm1wLK+8yUpcT5136supftOnhQN
NF10+2y58uUCz3mzjZr5kJTEpc3LJOYeSbP7poXjiIm/0sZ5bt9P9KzZ6VtAKB9I
TPFAEeUs40Gm6580+1W/rE3EAAupD3gK8lfmEADL6kKfk5aDlGSG6lD/UT+KOau9
X8JXOocc/qUI2u8lo4GHh14vAthrmOKpDNWTJ7KqWXtsp9LCApm5SGpyEHB0NtVp
RMBgIdh3JZ65JCt5j3lYv8n5j1ePbwZi57lU94ztat1pw0IbJY7wwq9ivx3lKXlx
QiXV0TqKE4lKWFnNlsNLIxfWdJ17DbbuO8lKilpN+ejjj1bRKOLtjITVNMkFQQ76
8nO+JyHHeZq7p7Y1iY7prHuUZw953/vY9uS7/nvtIOJLD+IsRSsjirVgZwnsm6id
mmT9WkqkM9FMQvetVfoXRo8EjqgoKFpfNk9tFdoQDDdq2g/kZdgj/MBNfwSWwg4w
/RJJdD2eVhZ7s+khqGKURjZ6cJfCIyHBsWuxuVZVPMo4RZhPfz5Bcxmy1DPPAoa3
hO32lZtmcAGb/CIhzxpCXWfeuNsHh2xIijuNzyZnNp7u0Eo++i4Jd9GF0m/9bvUs
LhMk2ByTrVbDM5Vd+wT3am25UhfvOR2NOh5MmZgrD4jjW1jUUrBk19AgK5MHMyPE
AGL8f2wumsaz2k46FJJZA2z15EJXtcuqFgy/RaLKpHpa20IiEg+9XoXAc175O5KU
S2iMyGy0yyAC5ZsJ2JRY5jKJE/W4bG2XNI6ONcSET3yN+nLU9xEiu5CwsP55LEe8
IqFNMjMpsOsn9X0stp1zA2MkO4oBvx9OG431teU0+LCxayoetP9cbslW8eaxLlLc
nhIVn+0BEzIxPfxhEfbt6hx1lhwCBaLi1K0Y6oUBZGQETnCjDIM4wEboYIzKOGZX
7AziA0d/8NoNygEiYOZzuZez9+S4Zn8isEmB9BnMZWYo596X7BRoK48GGu+Abev3
R1OZQ0CLSqnwyfECxNOJQiUJlM+auCqFTkdSv1HB+uus2Jp64dAi0KuM8peC/78K
EUAH5tw5DodwraBJxJdG2ewILVylYK5I2jWMgLfAFA6covLYy6QHGOEC8UOymhz9
pdup1CDzF/cmfF3NgMDTGzU9bvpRychdGcPP5WUsJnFDXOiQDW0EqCrKIR2H648X
SuTqfxBUO10x3tS75OhuEEfoh3Hw2lcD3j2D/DVxrKwB0Tpi5QesN2LteVnOy78t
AaTQN3aP02YKGv0BZlSvbeQvXUvsXtaF6PKnQ7WiK9FNZ+JB5WmO0teC7Z3V7cHf
5gphtlMdVCWlOLKXTJFhiGEXutrd5mTRfIK7DpjzG2SutNr+nhSZlazKJR9xlN5Z
Tjs3yRKf/OPaeU8iYRTfOi3B9AcWm/jJAtrWb18Eq2WTWTUCArJh6XEa+AJp15b4
dNLRa8C82qsjVCC9eKnbVH2Bd7F2RVo6wZoS6H7dzgU9y+72Vojf+6tZysQsRYU4
uBsbo0uweAiYHRsZ11o4mtB2KOzroV1z2P+r03qOyp8kyCDX530JIA36O1d6UBZC
Gd8C507wG9Zrm3V0NwqZDlBdOgf2bdAJ8iPsg8RtMxwLM825w9818VtiB4x/1wh9
F/P2RDjcd5Vqv6u/G/zrAFjmOx8dixfWR7bT9ed9xc5z5zhGXM9FNS/0ToTfe2oL
e48I7SFsG30Nn5KU2lX1i5EL3yQEjIfWMGsoZlGyxtXn5EVd+9sVUEzj12+I0Icc
SVuVfPtUb3v8nih2+AOHFlBFI33kuj1D2hEt0iAW9sBbI/Il+gm99DW6CYNLK7k0
OKZc7ktbeMNaBkbbhINNHbuY/4La5ZRB+2dSfrJ56cFBzBfQ1K8cFreEvbGESQAn
ijx7catgpVBBobQsDOmdRdqcRlkbQs9RXiWVmPct03b2+teSlVaG7nHhqbofq/x7
cBTzNWc2Lqy6Dfmd5pXfS8woQGQtzF8+IWxP/0dhdWinRXuIUjAEaP6Qs68HmPnH
EJM+4eb1hcHpvM08lnhUriX6Hr7HuKC64+M6Aq+XQmPnvmrdhDd8lWmon4mKb4t9
Q3gVnnST5WSv0bKvHCokmgCExLEtuykQpR03NWZeZfU/tnDY+0474tuF+Y3r/dTJ
ZmBtnaDzqCZj2rlgbAPHZtEwhyx89Jpys1MRwnUn5eAcg3bm101TjYF8Sv6v+HFA
opgtzftD58B343swsOn7e3+6+AJDfWtrU076lSoQcRzZsKTXSriDrYuHozL78FLn
mK9XojeexbXilpkMZ2CWLCQ1mRES0/HfG5Y4kD8Nku2J/POGpjCplDk43GUmm5A3
W2go0wo+9miEkNmOOFqfzoG7ISV6qmlaV8lujfr7CsXDWTi66PIrJQzCgmYAHSpb
cmQGfpdbwT1f/yJb4fC84SiZc3VY2cwq4omip2ObW+B2BEm96UlywJVQTk0PJlFi
S8bKcH/DcAl2qjOY6G9QtT20Uw8wr4DPbQBq6wj+AXKjI8c68DJLrIb0YowYsGgb
40JV2ncF0SDBmwqRik9Q7SoGaVNcFCqWxUUNuMVX2rl7YVXUjPFOi5X2YShtqFAN
8Xc3IivYIg1Ed5O2awbCXCe9UFQ66OYXYVCGToIGDw4MFpwv+SSeTW/Agr04t0aK
k0DSRxYNqUXEGNiyXYbBQIqgELKztIKwyqnYF7CLY77/C8cbu2+5grDPNr8wLznV
VSbF9Z8q0LyjqUwMDz9iTn245pBZPKFO8/60ep1IG1yhAf/RXfbg2ZQfo5WLLHnY
cErTNDQDGpd2vn6miWD/nmHbXoKK0PiF8UuFQHeG0SUdWtS8ANdlk20Z++JZ/zji
+MXPQe0kfmwYhayrfok9sw3lMHRez0+8lPjWDaVDNJPOmfkDSBwmnjcd3+bXHYlS
RtbY17zq5MckIoOVYxn2j1MGgnWj533WKzp94g2U8e5cShcUCTDjKc8H6OpEdajE
+8+f6Ol4F8jrE5OJklJNN4bY7jhcccybgkASS5yVt6fU0CzbYuYeRYRhKG3KPh/B
DOOZ2A+zUGYeVeu8hnJ4ykYJ7U62Ei7UJKOUnYR5jZtlIrzSpM5Roof9Py7z4yjf
NyOrRax/jC7Gr7ERnRZ+8aqclcn6DnOPeHtxtmAimXrEC0GuYxpAfIuFSylYWI+T
vXTercg9StHf4i0eYIki22lOzpbx0GapVRuXXF84b4KSyua2Opd37JtyCkfFQrtK
sATblS0JreYxULKFlT1YdqakrRHTz4hEokt2yWN/l+F11JXVDOfNaXDG3Pm/TYLc
gVUlEQHL3X2hgA3Ns+/Q8WvNvnKt1q7C/yAak/9Tfj+tyy3Mjz/DMHqs92H135u/
KR18TyxSXvaEw63tYMpgtDgnDUzVr8l5cBb1teGuRid+vEZia7dEwVdOvedLHfPo
RXU3Py/4emp6i7M8R6OhzroUGVa1I3zEGVwk22+q4EdpfbejjJGjdIewawZfIeah
nM8IczKo8H0tfiQu/hx4R/l8IX8HwVohOR0rRr97A16r9BXKqYwrbLaBh6l2fqVf
YI6dMYPnuRuBAnNReafrFHEICWz9iFzW6dZMrRUeBggTrgzOvxGh1QUdw7FTKhuJ
MYsuQsilbzfAl3NeRqJfgkzCYc1P9k99tUo4GHzfGUlUHXpKRi+HooNxQNixSa/j
Mx0eUI90L3U0NfEQefTHTsD8tXRv6co3ochXHRtaUldLL0gHcpgIFWHdJs0fP+6E
hF33I+pj/sD3Q93eNmuc+WX0d1nuPgWtG6M+fAB07R+rql9ZfH4K7xfgQdYK3Nuf
u66omzaQF5G9Q3xfMYRyjN+4T4SSKB9jQGj02/XKaJ/6GgNRfaKgP0vaqaJULSoI
imSgBXbsglAfexdBVYX8bMBbL8g4KUTKL3VlvRAuAi+rgXPfBg2/tlp2iXFEDCQD
RJs4ace6XWCoH/xr7jB0jCCc4B13vLvI8Ry7oTPDlD8vtKxrSa7X9Llh80JujTs2
oFkDGPN4EmRSHBugEtfUhIKiHRohn6YujD0FHyDN1AIbK4myXRfYYGSkQtqtN50k
zkOc4PHSq0exnfcOm1JGkztyAKrEEx2ya3vLSA9eiKr4jlIca+vQ5MrcWpjMZybm
vvzDJM5Vuya2W35kSvAiYNUsMyFKhaWJDKVJwx4gsXa6gOLfYx7+Jfr+pD7aiKOB
3xl2U9uv4QeutlErL09Ic3IsxSafRa5BA0K2KuF2IyLhs+HbGI9pODs6V/DFRKrz
FrRJ5GzE9P2/b5mqJwWqmsNFy77pebt8p3b+D1wTvnjnD7fikN/zNoExt8kaLpuU
ajblkeN1CN3I5TacSotAyvEZUhqRtsPb9fhXxfwcQyB/3xSZNTmSskWgkDi+tlqS
Q0+DJYhJR+4+Fn0aKAuzsOHwowRu356KzxKYjMURQ0Hj0/MXbbgSw0snv83qsvWU
nNqzPfQLkbKisRfkZ8MSn5d+9fk6U0JrnpAT/qHxJLIa6UkiQIGQZSz4sEh/L4Yb
lHaLD589q0W5LQaT1wU+4WQl0ILm+r01gbnymrwi7YHDc5WeY1NjkHP/W94po24Q
MQA/dpaSaYSq7hYoIURG6Dx4edjk69Pg5IW9BmX7wVPgKqOxyTfZgQGzywq9nbM3
fNZctA1Rqwg/mHoTArpQwiE0XS6/wxgSiVCYqiBrULZ2bnIoRc6XyUSNX+GYPnZg
lez0CtOXHOgfkn8MmbIt3P329TeQ1g92A5oTNSgK/UXZa6QrG4VntnmjY/UR5/Ro
dIGSWqnOLsjcfvlSURJ12ye7d/0gnsvzaoUnRNNFX5cz7g7SrehRX/UmyWNgczPA
w/z1QjgfKEcb2nEQtDdb7LDiuo1RnbFajb2pe17jsKoJ08svWPgK+Jgaz4jELBpN
zudBplqEwxXHQubvRaB8nDrngAKatqr+vAkLjr9wNSkmQdunXHSfhviz07Wf5CQQ
lniEfY3Su6olbNtOLKkVgrTFhtpPkilnGQ/k2oRnVMV3mArgIZxBruRAHX/v7QEr
wnToCKzkyt9ED9sQb11lG3qcOp0uzAR4h8YukSwjcRmG68uUPzthaFLXo4vdiCe5
vXZF8IaewgNq3Z2h9HhebRVZPKvugc0i9IFUVIpiHI5JMZLPRsRUe6io9z+GC38c
x23emdg+aGeRATz2sFFmI+ol1ZkRaEyNjPwftgGbLekFqRd1NHoA8jQnPAz014Tl
RHbq3CWZ11Eobq4XTB5PlBiOQNd5cuez3FNsaaqESfSS8KDHAW8PJLujPzf1UyH1
3suji7FQ6nApNWQObd3Ifl7uR6bFDNSTitIXD3S0NJSdwDrrSibZPmy42ZPqRJWP
6LSGbJHszHEKLmBrIMqyu8NMzFoT0OVLBLqS2CMPYEsiOWBp21xHDa+MR1N/8ZRw
vlUPYM/BZYc9WOONLYf1NhUjJ020PhjPzeQfE+K6donItSN4sxHnDHs7whCkkOID
M9hpPQPr9ctPMi+H9+IO0U8ngRDsgrEi+BcA2316piQ4a8ayqK2+Q+zRojDxuahL
Mni5k/vo6GI54EI1a4aIzGPCorzxirXPqRnGBUMFKDRxEmKnMXl7DskXk1zwBVr8
h3iHNb/hCGLOIe24VRiwhDE9PqSV4OLcUf5wcWFCDWJelOCz4dQE80xTJTggChHP
ixc04mLO0knc0TMOlkESOy9HfAsf3AnKk1mJTCGQRM+as51XivIVoy6s3ETbQPUk
0UZQ3u/EjQBzPlEoW682VPMsGrGRd2E/q22SnFRLZRKgTg8noSC4kH8/JmDdGHE8
2uc2gNZD3CTNcWvRf3kvKrqnYi+bod7gpjb5QmJbN8Al/a+0PHuq4aJjL7sKOgJf
PkHQbJmEuUabcrm9NgfQrwO9s9TsdEHxVGsaDHcXiAnXTqSc0PjJDqxNe1URbSL3
mhH1T8/MkeYMD4w5O8mwui4rj3D22uga+RRud2XKBv8b7y8UOB17Z8lF0txTDntc
MHH2nV4J9LVuHHJA6b3NqqCrDl8OIK7Ehmd8fU0TaAT6OD4vjgijfkK3nypk0t8r
KtTMhfPn2v/7Fb8Furh1qGirNkNhg91wDBnmBh4VXctpuRH2rrHU6Ll9UUsG3RVp
W/dD6Ra5NOukTkxKkY6L+Yodjw9l9CvaZ8MTpGMOBOhZ+q0IrkoFdgI79lrgOJWS
z+MSVqJTNxY3qrppVgYwJ967eypOxl0jelf9HC6MUEa0oMYXAROey0aE6oRHNwej
yY7ounP/oc3+qOPyOnAuUxv+VHPsR5BS4SYaCVXoxLKqudU2BKXNUjqJrKLqZQho
lOvXqwjTU1F0EwougA4urOThS+MoacfTdzay+9SDsWpnw1LNL6tkxU9OKEpBE+4G
Tklk+gTN0GYgGDQb7mc2hv6G6BHtDr8vaMIWvS5S8yLnBLR7Cf/D1bpQFqW7393I
FKjNF8ojl2lsh/ANH3HR4wvSY33LTwy4ijv3FNWNe3w/nacuivZZ7TQ/VhgqPwWw
QKDHwJ6pHJVAXJFdSqWhNbmlVvDdEFs1J/lWw0sg9AhZdq/Z6r3YDrv3TeHr0oup
U614fe8UaGOZ8UqfUI14GBzTcThREb6ZIIA/97e38E7bpZgyNeXxQEtSZub76vw9
P3FbyLnYvRW2d8vgyAYcuRhCBNI3dZz1TfCSwCzaartnJuxbv29YoH3bJq1T9m8H
paPpK7c7VwVIpp8N0KTgk4ELewyZ5tzkRhYFaEtsL60s6AMnihtRinDF33kpYuki
N/fnYEsab57CoQWQs5YUR9p9VypDMY54IV5rC22ZHNdW6bqtxD1u3glLCH6LES2F
9uKyMnclcFzDIFajQ1GjFWep633+VIoMoOtL4g6C04tcS+tjnia3340ZGcDgLBLS
dNEK9L/19bSxZgS6+GHhxXaOpvNbq6qpEVxM3wc1pNzZc1Inb1M4zr9Vm4kyd1Vc
wrxpVec/gc3yuSE2c1XYUiB7Jh4qkSfe5FfHy22IT73/5/w4pY4Dbi/JxB1MxhIU
xqH5/rpNx3eQFal0t3FLD/ip4Ns99MvcQm281k0iOwwbqOkspM4nSPkv9e5WImHo
9jpMwVf15UFNOCg+18HAt4jvrFvAqMmigT9KWu+BhcGRHD8l8rKxCzdEtYbr/nHP
HHVpPX2RbODEd/+0q+WTFD+I78mDUSUhriZxYE1WlRlGmuYnv9xwE8DDQP+/AHMy
GlMqS5G/gnqseZQlth0E0iWCYoVgTY+DC5QfyRWjes1bQk/bcSY9bA02feKUkzqa
TYFbZJNN+jDi+f7u8JrtopLGfGyuV3fmZ4+47P8xq4AVoUoS85I7Fl5/LGAAo6nJ
p+zu+7x/LA5ucQOaO1drHzFFF9YjBVuL6eV56n07K6iGf5m7W7DBx+JcHztSQkjn
Dm1WKz4M06gSWuCEcF7q/gO6Z01xZ2ZVOyGRp5yom+r+kf7hNzypRw9mmKCygJrB
bpcq8oknzUtTXfg4tewWztAitXUiIXmbIgrHM4tEiOG8B/dg0D6Avah4554KyR0o
L8MZBwDbjkd/ncOEhd87nLF44NNG0EPcUoOErtIzvyL02SzJM8MhzJcChZQwSWq3
i20SLtbux/o+wfbRpm9PlK+Q8rItzhFs7caKGvmUNQ6uu0yAYwZjxQyzDvunnuW8
w0ZWTDUz1TQzG4YubzQ8ohC6+d5Dc6+NwwBlxjreMIBMA2b4cVRxOAzH36avGtHo
HcxM9TA1c85xWEh9JmukZYaDuVlGskXwSstm7jjk20MQss8j+/jQYIJc2fGnH5eS
fF3/mVe5u+lR7cYMsXMhzRUeGVQUNBIlW+ySAVdBeh3nRXPEdb3y65MEsUvbSZla
irchtrs7l6PIxOShamdE2sywiLokSmi5TidbChwY6x79lRNBYxwr8XjgQcX6CUzm
Zck+tsuyGqI3jND7V6V1ndYPqA6igULd6JB+d/ZG08FF8RAds1OffIRitforuGr4
VTF32f4JDEKCLaM8iyOGbdAVh021b3TFtsknJw4S15Wuv2RhJ8aUvAwztq4kBaUY
0thO0NHVKmxUx0d760V/U9hrenG34hT4jDY3+mfCJZU6a8KlxvkH/dJ/RhebM00a
ROrYCq7XH+/ERuBLuoVw4bc28ywnloMxaWOuNPPnwW9hWFu3KfU7Uc4XWIQ6WF4l
5Q0K6ryAkxMQw52FiqMRGDY09uCl2AuVNSw4C1VCXK6c5az/3SLJt97Qhdh+w2Ml
LWreO3iZpRzw20f6vh+wAiMWt68++rXzSXNEtlDuyZzJpb3VeEMklYKaljJW742/
EQn7FpbsdfIyNb9pSmNYtMxaJMl6pkVnAl67KNOoH9dCaUZ6ec0ZiD6K0YSSi3WC
/Wz62CS76golh13qPw1TU8f9LaHWI4Mm+A2W0wRBuQuagNcqbDNVnAlwosk1ZsOv
Va1ImwOaQHkQa1RH/n3dNzIGwKzIOwTpCaoPKeexAgv247uZJIVvlvumUbYgCES2
eyG6Mb0B+OK3b4VAKnefS0RCoCU0P3Y9UR/vuBFvyHlTdFM7ppfU0nJguCfNRdcH
v1k4U6m4s9Ue4ELB/Zb4tHuqc8ve2fyrztj35xPkH9XVHniOrG6NPCh0uy9KyJsu
EXO+SAnPzcq8uPQnP9yoWmpq6wP/rwSRJvfjDK29NkwqEt62ol1kW5Y24VLF80VC
YNJlX2st2MW14nIYWGDUCkwZe9GwfcqymJyjeK6e8M36+7lHw8b6Jexrh23qewU5
wkYCtwbbeyiUgcrSZMRf74eQh0VZJw843OOKY1P9fAXVRp4vyC8pyI2QFHx8R3IA
fYDICbexIQJFjfQBQK+u4Xwoy7GaPOGoU/jnCr8pvSSCzYfImD8PXBpit5sz/dzk
6lBYS7kCJHsKJQoL/qyaBts/Oq9SJqMno/uK8G9lnw4THI9gdLFLC4UT8TfrvUJo
nm9CjkwEnmM4X7ihpokAoyZu/flKpcihVLnAL7ApJKBDkCiB7qT5anFave4XQsrk
K93Fk8eFN+Fj3/V9fJf/ldFvxmEAym9S+IW6Cju7WEf1aHoTTRB9nTrDEI1RwzdT
zvWZ3shR0w9s22nFcbrn/TAf+uQvQAxJaVgpPw62FmhH/iutuogF/Eb1dg1ITGBG
7/mDis2S4CuToNHrD1baHXkxns46elNF2hE7fNDlScvcyI71gDicJdFrULlVVhPe
FSSbFR+tJkiWm83+5oPW2AUQO5ydOM87kDn7fxW39MQUWxaGMFOyzyQM1N7LgeKh
IloFsOjsf9QVAq27SoUWjUtiPVcna6W4wM4xsPlCf0DkJtEpKrfkBJylEanrBPlq
cz6EwP1czyGiSqX2RuILxvsrOmrfR9dBwQJ4HDj8xT6fejImVb14rv6Gw4QqXr6O
NSo9aLueL9TGJoJljuGa34/w388vJV29hFGXx7XRP0sfTNPRHP/WQhIJcGebN4bu
+Kd4mV+h4RX3w6Ch2AbRIJMMkXhapoD10mmWZWcvYIhjdc6yzVIiXB/G+CvjWGao
SMxynrErQs8MMwBbMMPZH3SU2tB1Fg09FabgDJWncs5LExemXbOOhHGSnHToUwp+
oGlEjo7spJ/5y2aHWhkB4sR6EevrpzI8BjwOKO9uw9n5oBF8IjApfwVfJn4SRvXU
dFRnXcQNsEcvQGBGVk62dhWSXJH53aOixEIsgxpexKD0sxn1ta9MZP6VKIcr4jBn
QzhGDvGYF9D5zppY5h24gKddIKyCkS4kteTBGy1yUl0u1LoNGNWTnDymduaFt3lH
6HdcQpIFBKy9G0SNWzYNi4YTX+hKykXB6zf6+LqRuUnGNrQMxrMPOXnVmVK248mC
q2FEs5YJfwESYj/lKDfwOhCJ+cnX4Qqg7cl/p5mQY8OCudJdyTFcF8uS2yDW1l9v
t9BVgu79mI6h0NTcn2zyYH+9zlGPiO7MTO0VAB3ubELv1/l7D3hB6AKkTkglFOKK
zjG/qLsEhXtocM0GZ/ju+Hkmjlyj3C7bG0xVvc+LkUVLczlDWWzR8K9iIElxt9ua
NHXWzRn63lY8goo831Qt9FhtMCvFY+pc5JCm/H53yOeUcwq5syKQ5J7r00+IyfeY
gpaXljswiMbohpAktfoNykPfPItmmbFmeLhtde5jzvetKGihkzSLczfLjGwyMGJD
UUpYitqCvoe/yKMhH4LHRytOGv9Z9hV09scfgT1g1OQYnP3Hsl9sacsyHbbqgsJ8
yyLW0BOIKOUBIvsr6gpLdkLEWmiXwXB5DCbOFazQssvV3WsGGuT0Xn8TLz6i/iiF
ONQAybPJnjhpqPlL6E+ZyTbFBT/STSruL6qBPxlxKnLcHuAa1XQRyA5FmVHGG7dt
vTWCWzyWRCbjkDVAy0bHXpF6xeik98kq1nHwbhyUlnL7u1ygCMFOJiMbhPRA44Kk
yfMS/xIvezHVM6iSSnGFoE9gOdnJw8+XTeACJ/i4Dg8zUQA3PMKKFesQ6LmZ3fcE
Hpt+gFirgT4rYFpPcfItVotsLgJSG1pho2wlV3hduc09Jyr8LGcoarqdqESvhDuq
ap2+laEAYZ231xOr0e04HHA1WudPnv4D5tndCK9UuVejj2NC5EFz9BFT24ir6lG2
LO8ZJ3gE7yC2o5gV++YQB4PulXLR2xdLZyU3TJgo6/jzOQ1JFUP3p9uK6NxLoGSv
E+Y307D3ziO9ryogkEgFwGSsRG9D489SnayR6vuGt/vtsbpr4kfrHZjJvWA4uMMT
Qg1CqqZdAh+cKFgNvkL/kTMPJxzJduk6m/h1i6g8Gi8338OUOxvn0nO3GNcwd9i2
FEut1ngdwk/FQEk+O0uLhI1vD7VgaTg9NEF9Qf8Pv+teCGtDXXoKBsAbzxVgaf2a
VqixYIbHxCbJtOOicezQ2Cl5eF4EuixPvojAMJOyxUrl2seso+yEGsbpm4fTZoFa
gVyZCftmEbnqdSRcL0Q/z0xFg+BFSSZ8q4Tg3B0UhJcMb2K0fg0RBMj2fqP06j6H
3PT81laXMYZudvbAqGfsLV++6azFMb32ybKZWKabGkd0MHHFMS9k0xaJ/C21Ln7c
`protect END_PROTECTED
