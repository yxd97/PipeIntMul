`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufGb9A5ig2PgTuangbLmDNyTkR0ZS+utFiyYQptL4DtatCMf4UKx8tq+nT4wywz+
FlgUxdPKesyuMy9/NNGHEo+cpbcb12cWcgCw+Sfl1j/sY5GUGJLc+EFmrxxa/C3Q
ajiH7mNDIInKbNxekTHoRxxHMDtCLJXPElcZmidrK7iNOddwUG5xDkGy9cRCkG6R
4tYztL2YO6yheadvV0kQZtNP4Jwj1F/cEUz0856su02hT+oa72m5nBp7FXZXWysU
5kdLX1EZ/WvUwODwvXBdcXTj7gWPI7G2UZFd2jfcF9U=
`protect END_PROTECTED
