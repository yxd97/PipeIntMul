`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dcIbd4j2yuvKf3YlU8cQvRpJnW0ULPYQaWi3V/NpXe2eW89jHL9hFXYLHQWndgab
xbRREPnhNgd/YDzMCZIwxCRp1S+ZVr9fEHvrSwujKAuNVMJLDq2CjWCDjht/hpEI
dB1bMuEiEk34Fu6dsX4cFjtkhlcux1U3Psa2gVeDfBKaVXm3guZfX6IJ3P7nRDQn
brHJWGlNcuMrNeseDyP3+meCCPTWh3ziSOjHfNdHtenhWNDcnud6rf/4vkdq5VNp
1HQOBsQ4ULBxoAsq+vDWUlaBf1X/rlvfPzcrkZn71Kz4VdaztGYKUK0IwZKNXlw5
Or/qL95gB+KfGP3cme3KNd7Kq0ugbTad9BNnwQtBvOC/PAgw7Lh7peeJNDgvXqwP
xjwOiE5sC6voL1R0Id5vAPFZr0XbNjzrS4oa7KmEaBGRNcxS0UxOSIR3FbxJa4yA
WYgfGh8zoCs9L3N1sML5ByceS1HYnAdROxqmisRkEzympu5Lw/96Qtq22lHS0/V8
DJ7crDh46h1YXISePuLxYxjJa6cY9MAidt518WDsGGIHvpudS24naxZn/23P+0Cu
SANCzNl369MafRNU11fB3kgm3U+/4IHza8lN57u4+BzotqBLBbxcKfSupktDgZBh
l5y56gB3cY/FsbKdZnqZ16LsZafXfcDQ3hD4zSze8ph6qsLQLLN3QnRgR7MySQ5J
M0VM5JwJcnqWbaoOc7IZIIuKn07yGKRKNaZ2nswH4gXLcemHoX5RuJ8pkKjZkCts
MKATgNI5cxeRCC8KzauPns4DHgIxUpdwQvkjiVVCMiEgXXweFZD1uXDUsnKBlI+v
+H3WoAiSQugur9GyTLL4Qvv9w1d0QDtJzZHew5AU+8LhLg8zwgwttdwOHllo7x/v
/94fgNaEBzHPqQ1MZWeE+grt3qB64eiFHm73gBHTd+B3Xom2ONBhviQzdVi20XlV
nOp8lmuevfSXH7iN42pU4MYrotINMxs4joX+9hZ8hawLoKeBRIXwyx5pdrQPpVz9
XR0CvpG0VgabpECWbMIbKipqDgH+Oh/gaMU7dqH5S0t8OowDOoUwfm5gQfLLRvwK
oQhlSlI29S/YfGOK0Ruxgg==
`protect END_PROTECTED
