`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
edYIEW+hZwSzP72nds0IRZLivuDZr3xdhT/03AgLy8ekeMeiB6VJWWxR+VK9CYyx
huq6iuHV75G5So7CfO8eqVPBwIek87EMz0QQ4B487iZ8McnjdkX4izK/whnaN5Gb
xB8ZR+MvtL7jAT8h5rcbu5IuKEuGuXAjnpPiqxuuJbY7LcbzhZs/eINEOcqdp1bJ
n+Ru8lyrgrL7PUvHbA+FIWEx+7zhU9+E9eo5TI5bPynTUbO0ue02YkMV5DFg0pcd
e+uXc4iEmtDSAW9HmbqHW6cYCFcUNPq21vJWWx96kRqhOORCTfu3PMA/HhkfaWQb
ocMKBJDV4MCzTYhZf6M6ijZ1OgtEQx0BlgkSv0kQIy2B3FY366iTQHCvT6KnINDp
k5WvFHh153KtXXuwRiqeeZqr/RMZN7bLoF2pcGYrtRK293PSE+qwfHN/OMS3S5eE
M+FPQ6VTA5HZMGEulBPENUqMmp+jTjln6bxusr4y3T538VdtfYViyD4haRjB9YRW
z1ywI1QmDXkjamm9TyUJM+0Brwvr2Bh+eakZ6uGqp6vI+acVR2dHl0fs2BvHN9f2
qNGBut4FcDNuvmPphmSQnqnmkCDjcZQ155/tFjm5mBqXPdJzcOpKMTVWoLIrHhSZ
ZtDA2T7hkZntH1T0omAYBT3vUQYZfKRTIQqaejtD4RoPKcSK5VxS4SOAdnQ8b3b/
oEwTVuaGMvGsfNGaeM8DcD0M1TWscWtrOvlzbHARzZwownFUjeuWeBd2UEdpKPzG
7xniXCZSN+9ZltSRk5ydMaoZdHaFJquVVc8QRmN/c8sUoEYxaLi2m7tuS14ygheA
dueLZ/nGOW6fZps/HbIrb6QwwtlbwkTgf87W3Nlztp/QeUhYLwgD1YPwf97kBFqT
Qbs1zNlDbnHcSqR1afcd2nszeJvXQoNllbSehq0SylZGRfj8SQIQH0EIJGUIyZfq
ClVR2rrjPp7iDGB2hzVOSxqsIA442tuhVoavmwuBpe7ShePTT+WeYG/enL24HIfR
Nwi8dlLck49C07yBcfIiZwr4HSxaSIz7V1s7sIq05ZIt3dD5R3V9vD3DpnV7nB+B
A8KDQad0o3YNbkSPkXtG4YEhxxJFWjp8rSnNinHDrYxnRWBMPOH9M2IDHs6CB0WJ
J17ItBiwX5ipT7FotPFJ05q0ZfefAAR0jZW5PVkKKnQP8/6nzAROWL1MZtRN/sbf
Tpx/2AZSYHz7ARle8f8f3d1yKQgSVRl+EVnf0Z6LQ+uYQ8izdLEdBM28TqFLqcDz
QbsnWOWtgzlXtDjjIRIxC5/djchLP5r1zY1amSCgKMg/uWoL4swbMtU9D2o0/B/W
mav9yLHJ8+W3DxTY2F0mJ3CIJqppUiHFVt1Or7KCAsuycJCBCqPPQZsNKwgp76g5
nlkEOrw43vcwQaU5QUtZEciJSZk4hQ//JRoRv56vuPnSHqqzSDzAga+c0FKUBdMT
`protect END_PROTECTED
