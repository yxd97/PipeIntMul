`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eKDRPiU/89wLWnpjc8Br7Vap/PoYC84U5LCcFzQgcwIOSYgs+9FIKYOvl0qIvHqm
1u2pgrymvZYW/bCK4W/jRKOvhCy/vPAQC9MpZnz2NcnHtCuDPAUFouoFTvKGtfoS
K4IKcsPqswMkbfEv4F36UNmkTE9mqNdKjX+MdYbIaBHVxVvDSL0fEMwY3P+Hnp02
wmbCQjkwfr+tkYadgm8hsrPPVb2MRQoolW1z6l5lxBLSAucgiUOyHsPLTQo4PYKL
I4WMBYLTO5i9859xx8BYwBd7NFG1zjmg3NUH67AJwmQFy1kFd+IOHerk4VVxyz2s
MBVi1iOGDDiZp2yHKzfnGG1VPv5xWXT2uGhWXL1au9Ub243Qjhys5wnDScmY4i3+
K/J9moWXDa9t/0VAZ9+v79GOtnHVgrA3THxhomgInpvT+LJJAs3b5Yf60ouNffnq
w537xSjNWdk3EccgCYzJYKFTseA4pDhTMwEODv903kmATdDAyGpWENRZrXR0vIkL
w8MRoi4hJOK4VQjoFPPZliCVwHvGad+cnfnPNeJ/ANQClRNSXunvji0mMwCQw7l5
x9HjLdvTrOQmLh7ZyKam6PfPQ021M1TNApOSoNM6GLRWX7pR4qNiTZPceMER8Tif
eaqjQDrUezJk1ClfC4GM0O4JPps4QvbSMFTAeU+vLe7Q64CcXuldgnd2QaOo5yTr
4x2dtOJMIPVRg7fwwsJVOO9jxpKlen+IXySHtQbR21cTmpg/AR5K1xUKCjQ7rBOf
/Vpu8Tz21cpQEy/wYqNQw9CcVvcMZGHcezPPDmlIUGrirLLMB2oCsM/XU9BxDsTw
n6gq/SsGrozoZunpe56abirpeIXltdUIhNF7b58LSX/6+dhwLVjAhdv7rqxedrlS
kvqIcrDVhgnVLQMSbjMn6R1hDymy4YCD5g4KU5otoxh5Cnz+XzfOC6yZFZXhUno4
`protect END_PROTECTED
