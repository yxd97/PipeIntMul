`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYqeX5C5oDVE/uONROeLvWgKjp7MiqWsFg+wkBlu/4w4RCioo0tK6hD62huPvg+c
yoBZJtAAq3lbfuYIM777iBbwRCMOeMHUX5gyB+8ZeyVzZEE6nsHUGJLm4xNOpzfw
Ob3HOWeWaIZTOAajL0ZWZdvDzJ5Zat1RydcRtc9D0qH9VXxhcuQqV2fuf67PI/D6
qdlNAZ9W7qsRUF+2s0ECmZ66iwlRS9g3w4fheREqr2Vr2rOuk4yxOsFcxz4Q0NM2
JUBkI/p8sMlpwgY/eS+MC0uDaN31k0M6u39ITAvCNVCbagHsAx71Afty6UCsIzdC
r3eX2YnAT5J8BmPZIS74jUa7ZS/NPSUm0TNK0DzCKt90z7PNyBhOmCI1ZzCcWMFt
AIdBs1/UHh8Monk4tQx1CGzNgl7P5hZMUfJzcAUnZg5bPJ0cGK8GuJHHWe+ROEMx
sjdtti4a8gptL4rz/VmSTOQJ/aMaecvwotCGElBGq5l35aQk+VyKOr5vLDHi+nSg
`protect END_PROTECTED
