`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YoYBi4NuFJruuy23rJgMg1LaSyOJFJ9Ym45+KLZgoHbC882EoQQwyluhSUvt2RHY
ThbkyCUDJRFwiWXMnZBJqujxLiBpNM0vt6J76uflMR3FQY+LeziEzKQlklRJfVg/
Z18xAtRrivxXFUlzTNcrjnMcWG5NgezLyItgmJRAIIr/tPYdo0trGp6bsGrUPHSB
TUO8cuwqSDie5jTh6EGZO9ac5aNEFqpGYPk8Rw+PGScYpHv4p7Fy8PGXYWfGlJLz
mVUcSTJQfBH46OdDMcR806P/p2BLMqcH9dG7w4D+icGQVUtGwqowpMDt2Rfa3L5O
zScI3cWUN/8cu74wF21NSjIX2PaOj8tOPsjSteBUAudrI9za7yNbVVYvVzVgjjsn
0TM33DhlMu1pi+MFZeuFZVlTfMX5qaHF+Xr+GBJU62hDbyKgnVmjyd8sZSct/LJX
KDt2E8RnvlTmUSyAg/LBdJuXArlb0kXE7uOQsDeH9jVZk52ZyJbxwe9AXTgLCvpm
CXBdG7zR5TBu4Rd1+7IqoMJWEZyd4XKNao3v2Eu4MS7Kp56AgxuItKok5av1pAaf
f2DmcqCJe7hzWCVebM7eg5FE5H1/jJYmGpxtDLbRxF8eVtg1RnPjbyAKAe0pKyLx
P/0iyZRTxYcb+L2XHUnCSi6zAlBDwgAsfPL3V+Y/HmGKvKjv1L2VPfU9Rowzqzbq
1s4JzcA/Tk3iykt4oJymPOf0E3inO1Qd3alpliRB5o//NO5Ad6GayMSGDyqODSO4
eurmNfPGrPma3go1IiQEg6Z9DhCx7tJTikGjeCp9X7h8c36V5Hea/e77lAluH+62
IMhzxqXnBMPffLCOcTYSjh3UfeMBL8XFyoePh9aqWWXBpq9JS+wbPkVO+MIfMRdr
4xHRGREkqTBV9wAJjNu3gH5/szqNMP1N8akIW00uatbw/v05nQ+/Yr5vC490FXjr
cZjXV7ty564ko8fUs5Js+/prQjvOd+hijkvoliOPW2d04QefdFt3DX43aGRpLuSj
RcvFZbu5840IwbAb+xmEsCv4nde36LEW2o183YKeE5S3hQF/Vyoqo1+xwege0yKg
b3RxMvNufeCxpUZEXkOtXXHx9sJ8jSgWOfIUvH0nDzxcXDHybm3J4F7WQhneBiL6
zxf4UIMa1XsZREJB9ytmmQ57gqpqwFNWcwbQBtbhOWddY1VVkGJqmVKJgkuwfRh2
PsM3c770n9YF+5Qbx8j1MTUn26w2zLdaQnNYOgGj66sLxzdsL126lzu+rhmdSb51
2BIxqswmlG/CS+odyFzYQS0jXAY1ejvdduaI7pb2gfRuA/oNJx4QbdtLk93e0kE2
2SAECEtOJs7EIExxFa9KGOKax1jsnVrfnRCiofx+VwMQgWF10uazPDYkrhdcnpfp
3TDl7DIc5yvqx9pzP059GmoCq4lacStsB9sKZVCEdaq93o9hK/+gYdqoUk94EqWE
+OhkR/onxGcFJ6HNlOsEtM7nqqflePTb3KsmbC9yUBnn8sabyYirJwQd6HqQzIgF
+KYr1utvPYa2AVjaHho5lrqV9V+mHykI9HB4z+MIouXaCjsVSYXkHC2a+Sd302qw
lnUa4VbXYvZCYl9hMifibo/oSRzMtBN3vl4sXP3cItL0/Clb0kXd9dJToQPsL5by
j0SPmdCPhNQpZkgakIKZ1MsfLD+j+vkuNb4gVnSwY+MCI8pIgb5m+tFGq1IjPtZ4
BOsrs/tzoCuUqrkoRV5mi0DQg2BeDWRGWI1xflvNv6E=
`protect END_PROTECTED
