`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
otNTiiX3lIAlsRD83kjUWKlQZZAXt19mPPIjwNoArarO4WMLLLrpRCk6T31H4RgM
n3yyoVjbazCPMDpLd9SlrIpEjeGIb06vBXSLgrPWatvGNBJw3FNNqdSzZfrVb33q
3tQog8ljVeae8ylPakN81hO7Wx8/KY6+LOMksYmL4HCgYBe+UAv5F2hN4ZX+kv7r
wcSYMeuVkCnytdo5j0NdQ1DTQyg4tYGdWUigfZzurrpPBl7Iz4I4kH6hqZ2omKp6
zmjZBTuvsJYfLKBW3vO8HlW9PetHne+7XbaPH7nefxyjJl1oKib17j/1nIxtcoXb
aQQTF3sYWMB5wgBsH+L2fG+jqCb6CyZqhRfUXf+CfB8=
`protect END_PROTECTED
