`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uATsl06/bs0ncBTZhESmFblbs3LufnTc/yOTC1obsm9olwIMbwNJfGLAeneoU4rp
N2UI8MOr3Ymulqe1GNRCMbW9AhEaDYQqSQesSVUIBLQxFWjofjd8iphGnqMKFPHg
aflQG8g3qvCTAnqSgvJBvu+64yArnksO/ST8+yop+9L1xjL9fnGN7Zu3QnRQ84z4
AL6hHajUclxQHaORH2PNW7HjV1rvUnHTml9WaJq+cj7BkoBCfA3Zu/sWDJCQQ6s5
sVe/NvNZFCbznOMpK4TDRfbgp1mNkvY/bpHCVwjGMuZ8ilpuN7XhsIdsyAKre5xa
Z6rwKRwlffsc06+0WuPrRqCZeLKXemegqWL/5lqVlo3CHoU82wWa61nMBbkp2mT7
ricodeBCe3/iLJAGVts4LixQmbAVBUFYMUFyNJCRg0sg+47as36s486F/d7/fah2
GK2kZg2LhH0VFo725h1g1FWqZ0cwSUeSCaWxZeB7vuLajdYKfHCRQLG73wYJbaJT
6PV0oRyUHHldDlyuXaDgzQw26iqBJMfU5rGX4ULo9OE3q/NQsBisfx/tTpXzVrnY
2BH7PE3nMbxEVLftIUdDC0NYC7OIArelaQ6H02fnhcE=
`protect END_PROTECTED
