`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rco6ClikiFg+2SR587kiYFWWlPFKwmZOywDhY/KtJMxlSOaDkqXpyync1kLfC95b
CwHbHSP1+15V3kd6A/FgKSlxZ+tzsnb0uMAaKSj3LmKSEEBM6DgLwng/YpZCKknV
XMNe/LGGdu07zgzpM7FDKZkV8hpQMF8mWJ/mLr3Vw+fgaL17oZy98zIXT9Uj+akV
OaXuRnos3SwZxSF1tB/j4ih3IvThMhmTYqdpqYfuuA6cGa+5RPaTZdLbydRi/JO6
e9dk114HxHNwfgSYvqEXz/IXtaRrBuJNHzTr5Degf9BXF/N3LbGlxXiy0FZEtq+t
db1r2NblnniNgI9wki/0/Clm1b/NVTNGH88a50XGZUd0iE2ijY4TUUsQvcvoIKew
ef4QXWeLu5oE9ZCodB2XEBHbizjV9zqM0LbyHp3IDBZq0V5lX8fPQcSP89rk5Hhl
giNz0kJhuMgVxEbm6fMqqcnfmWB6QI3i+i0zFxtfZkh+zM3q3n45jHC4kAUqYNWx
C5zy24tIu/ent4hzLUlapR7Px6D7q3ApLqRsREk6LKNvVsKsLf0XYOJf34orZAp0
fy+3LEmJ9O5H4fl2CA91bu29VH0DFSoZyEAT8S/DRXlawh3Ke8pTBkVeEuQ53EiT
wRveDnF5CxcAYpcL89duO9eURnMLJABNm53TNuXGWH/b6etUJHX+SouZjey8dKRJ
`protect END_PROTECTED
