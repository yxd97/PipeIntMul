`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9V6/eqAG1dl3Oqxa1j8MzAPHPZsZL/oeXQ3r//yBEd6R7plSIavvzX2nu+/iLAG
L8PjMVluesk5JGr00vev5BPLhuiUBeSUuspe0GRnw9rrVIOxPAbwSUsxKwZm9wVJ
hRkQfONwuQAu78NCRkmE3WwSwZl5TkeroaUOz2gNbZDecOF0WCWMmC9xA7zoLQ8m
h3KgsjfYrGR0ZC4W2S04lx2nLWpH7ZOvY/X9lN5VkLTXUD5QSlrrO81BnkyADYwd
FDZztnAE3jYwtGXyFH2VrA==
`protect END_PROTECTED
