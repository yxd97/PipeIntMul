`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
go1MSLshALu/qLRE0CUrG4rUID03QjpUtb+ekIpXm+V9GIwvh+ZLUJVO5D5H2Krr
A4Z+6iKpxDRf8Rfayj30Kbtf8kKjALQFzAy69qxLR9OQBWuaGXNEuqEljpYubVfO
JMu4OZCVKDhISGeEMWae3vbBW7eCSitqrJ9TatFqn2BjXcZFxgF56YvB7FuG7jWB
57s482KOyr8yJ58U7KzVgl41yhG/7PlxggviPZx4xs2AZOvVTlJEL/y12xFQmi9B
NWiIIuwY5GnUee/fdkJ7Kg==
`protect END_PROTECTED
