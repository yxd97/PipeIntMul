`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oEuYpFtCekUqm/Ogq/mWnVw+8DEzrDJtkyL3brEYo5+cA8B5IXJs7fQ6PmaeHqug
UrivtkgyrgeMwkp0OVnId+4s/GKMZeLUyooGhzevNNTF06n3GwzDOCZsWaPHv9jv
O92ewDgP0XFCT2lXeTLfam7zCqWcKfAwZC0Ae/3kRKlZpUB72cKYPq+4TY5W142g
eXosIcSZ5nXWYFsG3eGySdeBslq3i9KIsZg3Sg7lg3cplJpn/bNSAvz7doVapNFT
NYgOyfruG7AaUn4opx0mgBMlCAWDy2c9/b8ZQdq/1O1dI4remcSTWCv0qwFE9lip
bavELD/lCZaHSWs3Dzqh/ZlizId51DDqj8nTMpoXqQSuU+v4JXAKTOaRMVx1T5iw
`protect END_PROTECTED
