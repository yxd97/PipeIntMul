`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/32FEEsMGllABeDOF7ao9EFCCkA67oIRny9bCuEYpZmIEoU70qrFS7RZ8/lZarP
5yCxvfnj8uFEEiSawHoIhQrbj9VBKiedjC1qgv7DR+ZM1ryOiQOKwhVEA8SguWab
KeZwfKVCHzvKVqBBFHQ0RIul//TixGOw5NswoaLDWTnctB1Z0prymMwn4pL96LsH
laKqCEMB60J1dbrN7TmA729x8bI8JQHdGH6nHK6zE8nr+XkWUk7qgt2IZH/rDzo5
QyvwsUYqweurky92Kj8Kb1/2oZ5LS3Pi2PI4MgTkWljLoAj6pD/v0RgoVgGoqW6i
EpSElyOWMRSlPcUiZIahxFQGdQ4Xo52QvLEBmVZ+LfcMzYvyeX5rfL6EP2d2vphE
xmsmgFIgJ49tX3UnXpFwUwJIsXtab+H3bHojRPBmFQyP8zqX61Hi8Zz+7vIZ/Roe
0w7vs6gvBaXNovYY20H7xRdQ7BfDMlM5BDu2LFfFx5Yqc99HVPZKY3wO2lytuGAT
NSn9ZhU8nyrqgqCSuXCHB17XvCH3DwRhIV3ThU69Hqz9bJvyBYL3FTioClRSPv6t
ETEtCeWpIox8KIFDU1XZtPY24kBPPd6KaBrNvHq3r7Qvn2mGu0hfkCQbf04eaC3O
sOnmgk8R8b/FnTMIwgAcjUWN7TkZG7O0lGRhkj6UaBdMyVjUj0h4lWHIm2sGEKqr
tSabQYgrgp28+FJDX5qxKUdlHWBMuyWGYtaibPsPwvcqaFvUpKRZkgTeiq2aZCWF
Eyc05Tv2MtAYEz8iPWaF8DLYhavXpPESNt2TaQIR08RTYBJn05nc3ml5puVPkojx
8hpVgY+8T9mkpSFrLe2fQVzLzxSY4GuVYlYMeoaKvA0qJq5qSFvtx5HvgF502SQQ
f+n2YQ0Gvi7j3EqUPW41/R49FLIOPiJGuldrZ6cqRtc3K54QQyWoET6RbNevttuQ
lUnQHy9bwRetEa69mYSGgzPq/RFey/VBogQg0f+OD1+B8Pglx6gda9mN++Jgtl57
TyOTq1DnzZ3INLXQOLXGu8w1uuPGLwYxFqND8CPa9N0nkCbpNajgTliRN+ZFlbuH
9lhKlZdQaSKpD2WkovCEC4RW+vaneBJ+Sr1CGhkRFrjTO6dpQaPrVUCVuYPOkdrf
EFB9pmBNKKuKKUZxtTejOEj9Ho4XCAByGk6Ebfj+5k8Mo5/j9jFe/HWxH2qEJIVC
WFJmV03Kw5IbYUHNOE9jF/7K6l82Rsvo5vzL8TCiRbZ8BseX/1UK9F38zChdsPuB
/Gm4Ur276EW4zPay6VPTmzI/w4o0Zqn4zb9BMQq3QiwsLo7cufc/9duVLNsNb8NX
7DpC/D/9eG3sRN544jdTl4HLPQl3b/4iQBLCfm7C9Xzb2HLW+wTZrtLphP91rxq9
+doKtwca4pO3/FajNGrqB9PZ1WBf3tRf8YWiuVLEujL1N1k5L/dkQt6hJsZfxK/h
QBwtK4cMAKpAg64LT7u7CaLoLLzQ0C67+6TaMw7XikqhyPDUPj3PDwDA0P8U8SPF
ym/P3tz8t/HWicGBG11smEiCWufaPYpQeJaQPxipOei8BQdoxHRICW3OyYqbG06d
F/tgPfvR3p4xuBKdVFOMJ5KuKjzQ0MangkoVn7WNwaOgMToPjLq6S5BkNmqhxWy3
ZiUtkPjWztN9glk3Hvn6kveM1HrnqbaOcV6/zAqvvhAbPjt3RdOcT47ESQxplPKW
ffy+6C0Yz4qvddXTSuZm6pg65QHdb5JW8hmv5mydxkJ2/o8xibeNirf+XqJuTBBO
PXN84z8wx7Zh1mEqifYmzuQJUvCVkU6a2koYIMrnITQ7nbyKHRdtqmIVi69BqT0X
9HpzfSORujmG0lCXAzx1Ml6pW63eGOk+9UKnISCaBiK1H8LYv/Jym0zovM/y5ARJ
j4LFReP/cqYop8faysbOKg==
`protect END_PROTECTED
