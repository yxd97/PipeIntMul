`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pjYlfDn+S6PLmh/QSLN8ZnbO+O17QGjvrMAYRIbo+BQMn4wAHLnQY76qPyxu5kvZ
7JVMfzqF7D819y0ambnn5+BJU+4QuK4zQdxyK65VSI3MLoM1NkWHwV9QdPYMEL6u
c/rel5sGOPZVlsLhMWsxl2yIgGqHirwoBiiUr4EL+yb/srmGjCVlBTzgN1BiLaTN
bX8G9m1WI2k/z7RVUyreHU/jozS6EbVtdPDhALrkouIC8/ZndAek9XJyC1bWQ1+7
GrQjIpfi1YNj8zg5HlQwaCi3G4VGj8ntySik6b0ayRQ0RN8ZHxeqFKyPEBS6krNF
hPtuMGXfPMSxgsodWwYexFSfQoB2BX7o6KNsA5Cpo6lAxjxzP7IAXH47I6oaHYbd
3Do0yeLNmaTQhbebK0mntg==
`protect END_PROTECTED
