`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QyUgUTLe+LM3pkGeIT6YfBoefLW8no3S3NOEm6rwA3OLbR73cttzjt7VlzsKkc4T
C+AO+iEo4LSGQjgZmV/vS/Dcr/UD+FZqEMlLLzhciK/FOCt596B8YUX2ulLa1WOC
ECJubWS4iRK5f4mXGpbGOOTi9c1xD+GQlWAVlGE4RGJ9tQ08FSiZh682ALO3xGpc
li0MpbAWFukVKDpmLNG4rLsb/qTxjZ7dX4OSa54kitjxx+w9A1L8hZiGSM9zOMVG
XzKB6FQeQe+xYUvelYuu5yaPt7q6NQY6wAyCKzQt4CW10IFGgNLoiSWTSWMIQsiR
vRzOvGxvnB0xZ+VvkyU3Z23nCS02Gn8n/2HLOokpQItksQbi6+YmIpIkWaaNmLxN
20WZ84+hp+be5hGnVMSOmU4nAwS8FKDWhIRiTENUO81nBGNIogitM0NQmaIleJ1k
`protect END_PROTECTED
