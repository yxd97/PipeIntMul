`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBENI7wKGt7JiuJ+lH1BC6xk8ElrodTlGcPc5Cp4jNXF32fjx0202tGkmB78PEnH
AjNKq+CZ5M6MeWmFacH0fnSWQUGYhjGlpZ3aJyFVTNUINkyxe0+JvxlyuLz044sJ
XLmJdPxaVhA0N2H3UC/KWjr9v+7bhNRvQ7Wt+ndF7jSYZrk2Cowy2ZoHJEQJxxcQ
9yqJBG5x6w9RugOv89yU4CJzvC8cB/oqCa0JJ1qNl217Red5SozJAeq3yGBOs79C
LuOEKUEeYVW3+i1K2nPz/sgIm+saByRs4dDPMD8dKXl85YsmkFO9Uuf9V4LpJHe/
4UeVQIUO0PF1VV/Etx3qZx8IdDV49O3rEx3aliozrv7YNGfmakCyksUhrq50xwSi
fiPAORhP6cbd8epsHE3tiUz7yThBR4NEzMwGySyltWg=
`protect END_PROTECTED
