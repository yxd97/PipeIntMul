`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjkM6xsBvhrBdwPaftNK7KI1h0axYWoSBRRJJfSHh4xv5SSMe/IlI/XcH/ifH0Uy
G0EWNpe6iKPFt3EvbrvVsXfCxwtXsdvaz+28QBUj8u5NEvkZdEenHUIfuE+uovk0
pXEuZdQ2JC92IiBb38bYGkEm7A2QJcWfkQ4o/lIbJ4RKjcs4vctW+jHs9oRodJ1G
zEkvRLUtrpDFe0+M3qck1BSQjGSxd+ixO6rd8/91Ahduo0ZlHU3WT0xuACOE+q/H
mcMk57dGNMt/l8rQpmNPpGR+cZHq0BEPjW5sKU8HDYU=
`protect END_PROTECTED
