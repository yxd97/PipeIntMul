`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0RWg5qGn/TcETJ9c1vfHJXCve0eWQBlCvOuiYLmsjjeVi2p3Z4SVuEUBZKAvQNbq
aJmfB4SYxaOCnnsXCmtSfo3jvh+jHyIhErs6IkJ5ESSHt9+QvdRDNsnbsM708SCQ
2uyLhD29YlaMejgtmqcJ6MPt8gzjldvqf7XoCy0IdCMEGmYsh3RH1E+CSHyYBzNm
RxRooUApugF44kPD4u+WlgsACAPpSILToORMOZDrfAsiCgEF3E/JV82PzX4rbK+d
zaiPsg2BEcx8mQlxNbi7sKg6Ex4BbegCB93Xyef3CVmLwgQ2Ec4LxYcWAhVBmRF1
8zdwm8Sf5WUVmfKmi/eu3UhCondFNgWKd/NHulODuhMa2Hxn3gGg4m6ALYRP25nz
XwHs22GNcPO5zB3hM3safQYzlzTznQrfsRVDlvwHQBPOHU2rdkR5hmo5oKyKr8Vp
MbDQYOMwOGfmhPRKxwmDTDLQKZze6wiaEXJRQ6wc0Hcp9BFzqVoGIbCkmdnEh6Gd
qk11CYZhzbkU4ui1y+66JKwj9ISbkmAg/liy/f5TQSRQOSrwCfxlxm+KKEFLBpOY
X5pR2xnGugnjHRaxA7tOWw==
`protect END_PROTECTED
