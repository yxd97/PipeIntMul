`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/vb+VtWlzppQB1VMOSp0WdJY0AWWhvZ4rMKX8a56xxIM75OZzCzw5PQQnWn4Bb2
zojVjQljDJV8LrHgz3+Ean9DRgtIxn2ZuOXhVJGtT2fgdoO70rVjkuY1TEUL1C8m
zC/32GNQzAdi3ZypnlOSSGuGpPBXW1KIfFQ+oOs++aQO6NBUUbMm5VYVDCGoeogO
mZR6IZ4CB46NrUqbqIbMpY/4Ehk0DhNhI8KU9vRFchjXmTGql6VdZM0TWcU3ST9a
GeLYdZnxf/5nV5WwKzfIn77QdXRWn672Jme+CDaMGbvR8bwm2ESwDJWbrZVTW3Gq
mqk6FyW26PwTxLgc4zRWkH5+PC4V2Fm0c8tYRfrTDWfyjVDSZQ2ViQmSzzihUU0K
Ean1kbovvgcNoE5I4gsIhJZkqQYSMDQV2+c6KPuCnizltP1bHNEu8DrRQZ1FA/su
xyRGjoQGMawFR6YfKVZ2KkawrV2reigrLiodb1JsaZuw77s8BrMOJipH+SF9hdle
jeEwFFuMEa0iDVDbGcbN2WytyGOohg1IQikp/48efQr6fNTdXOofuT1JoHPE5G4e
A0MfsOn4SpDXu+2KlUzprujxjbkDl/1Gw8rvyTV2P/WZXP4E0KDP9sP3L3LN/Sdx
Mk30whK7e1SyW5gqeseZhg==
`protect END_PROTECTED
