`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQesKO371niryevxDLIiDmwbXpDskeqLKM9DSM7BkggEigOYbD65fRjd4KHnVDmM
JAjccQYQ2Xgjv/Gfrohe44By2mjXx940LnYQDuvWRCjHsNzPmMcG6OP6/6nUPG2R
byWn5jWix3df0nqNtAY10TA3iNVNcJqYSzcLPnDyuoDe+C8x9mM0x2I6CkI08TYm
HxxKQ4B+KgXSfP+t/gxLRP9qkcPEgStzOMBGycwIopgEE+8sufB7I9kh6WZLYHEA
85grDrhXmEYr10lb3owNl4JjisWI+ckcCAvPtugxGE+mwl/LcfChQoO9dMNsV0YP
N40c4irmkMHF0itBVia5aj+G8yFtzTtFahsly+h+LvQMiSxl4zDTJ3bxc+kw08LI
A+LrSeCAqNSYCfAeuVlBcw==
`protect END_PROTECTED
