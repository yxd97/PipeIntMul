`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRD9BWeHzdw3Gs2I5kFKBNCQTUQVu8UyDw7bgQVIRbK4fcfNycfCdWHCqaYusRFT
rpmPBT6QqHNhyxwz8ueAGmIlDbaRDVZPUscSQB+8H/3dnYy6AoRU/ElYYaRUQtdw
pIjzuK2sIIVtRMEsUQG39zdzWWgHsGi6RHR2b6jsDvCbyVvyinou+VhQztikigSr
r0o+hXRP/tYctA79PKAsYHgTrtoHNHx2mYtNJfH9H+Q60P1FXtkWUcNIISQz9zjT
Rav8hBD+J9zIVF4ItWlWDYBQ2Kzac2e/BV09viXDjWE=
`protect END_PROTECTED
