`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDDHZ8i4iOUaTE0/mE1lhFJPBhp9IB5hB2UJh4V0usHB+wYqhIzmek/hUN5yBk7T
t5OVAZn5pO41ASHARHCvVbnOil/xbHDfsOT5x9zv9jBgmNPaJ7Goq6GsIwOft+TE
z+qO8gYs0e97bC8c2+K4jFpsL/EztldiPPY/DG3uKzgoD+FYt8WQ71jXjuYXSsWt
fT0Y69HadqWJLBUrTlL+sRgZ48sl7QbGa7x1XRdUAKbU058zAOO93t0+Hc4qwGy3
clMI+wiFiqkCO1BFakGmW5DFKbiWTwjiLKakMvn5nAydp3gO20Qt6NPkrhmB2www
45VVy29FNQrX1e0fdEBA8sXxQhG+eBml/JciZyjQ1Pf8whFAXF9THS4zpH/TNcdd
dMie6iiW5yBxeHRVI7Vey1YBYNttD/AW+8VwwqcNQvzyUGgi9c4xZ+jF1tiAguKa
u4bO5reJipjU95R+Xrv5XoGCkk2I7Gci7EXj8kXo9Nw6qsS/QNewiDMfWAH4rN+k
lFkp+P3MDarQjgayaJVK4bEANAdyUkorF/7S1joLF9A+smicURaDt24SoPrKiqCN
78gcvqd0SHPJYjSRf3LQew==
`protect END_PROTECTED
