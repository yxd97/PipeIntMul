`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HIzRWJnM6VWTJV+9ApWJVUC8OfI79i5jAU0VR5YcLN0fZU5ubiCiJhWZbWfKpJ6z
A4odlbuD8oH/UgoXmI9YVTy3BRVysJlb1yZ3NwKWvL+hUTMVFhAbkeCjaPb3tovM
tZsRHyKHUuQFMMAOmEwalISRTgCYgI1AGz1c5ZT2FT72nuWntcr3bro8k5geTG7c
b0v2c2j0/1BT/DEPlbbizJol2KjV8U3h6AVhBdXohU12iYpMnTgOYzrg+e7xzL2E
5b3cdpYt/UcdMCUXJEFuKgGV109fbSbsNmwa0/TuF/7rE2HqbzxgQyfFezj0xaVl
m4hsd/A7mdnrmsxfaJCBHgUCQGT1bg+Iox5E27r/XlZNM4Kd0+M/eODfaB5Qb85i
sCX5rTjw9K0Pr/erke5errLXqGRvhT7zvaZ8FJyekvl3KCm5kJoGN1A9iwqJ+Czn
5tVYu5iFq71+j9E0YNyqleM+7p3DI3mAqarbrOmeNfqfJvkwze3m+6foBQMDk6T6
08sTKaDVrBTFC2hDaDIWZFjSN719LmfQKE77EluH6XTJhJNVKkffmus8IxA5PQp1
dT3acHl82yj3aGafFKayWI1c9mBztJRdB84Tlkixj+swxzSoc6YW4EF/FOlH26tK
KG7X/FFCKVwz8gns8Aspbs2dSme/6mts/u8pKrbq2qy0IfIO7tPdTIOSmgwL/QfL
KQ+NchW91SxVs4BvIXH2lrfpMftCvnY+/vSiXTHUKInZguVu4wg0z9FTWZ5VaNAk
n/3zAWsR0n8EMMfONtaAcFaVvZ2hEVd9Ammr+/am8XdlA5KkHzCRSOnkY51qHVXc
dHeEHXqM52fSGx57yVAKvpM8mBluBb4hFXA3JiSZOBFapB/YJxLBMm3Uxt1pq87n
65OJNWC1pqi2A8HF4yRo0LOR2gHA+aQa2g2izJaBGPdMWwIUYVtJStX73fXGmZ9k
+HirK2AGLTjL6XAy3Cast/RFKvpjnXJUifZiLa5TT2ytf/yb7IB8KKrtrVNjG+1e
DOytPE76MtaxsdMLyT0DcKNJcEElsdwos0I+Bm7Xr84yG6fTuU7GXDr5oVLpwD+m
X/Yq89e5Gh6rxnQiVGs5vx3AQM1WLO4XWP84/YGl4aculbNQAQ1S0I15OC466ARP
wvFcZqhxKMXkSzp31KOToUC+YfGSj1zWlVr/dbEWlaUN2ZY0kO6xQQw+wBWOEzyG
l8pEIaaURwDV7aQooXKXyaDaQbqiDbuYa8ulq1lR3d/mjt+L3b8WDyMuS4c2eW7n
MvJtOhCjjJuUoYgWwzR9+bxRxm2FGqg4tgqliI/fPoNLYeV1ywWJ137ESCeCd0JQ
2PuvyzdVbd17/QZOl89KGJfuWHDo1khBmnYs56iBpEiqTF53Y0YNO+EOZB8XmRxa
WNYQ/8Oizhgsz5dEyhEUW1zBGsroKUDB2f27ANzNMdl5bov1UWtzwoR8OiVul5WQ
LuKlmlSkBag1i3LpnJ3OduYgyXkUqQ7+wSdAi3zOdOLjh1Ym1im58uxOMVrWLRIe
ao6hcFS0wp6WdpMjygKEs2L7qSmkOUZSbCMi4uut6GGzbO/Ma/0H/xKh6cnNEUFN
ZJsOxU7WJowZXLQqCQuBXm6Ly+NYgEf4vp8vlHY3UicCwWQTvhJUkn4ex5ieSmBv
tUs1Ds9dckG35JKR7Vt4DEJqLVr4XJVhyBH1tfaaXjfMLwmpyJv99hah2nNRAaA3
sK9EKyYFDfOxbun8AUiAIQTFRNk4qAF5qeln71wObvlUbwF60EN1jGh5HVAemIoL
RCxrBv7TW+PtWpweML0RWzO8OmR97UbktFwIDMykN7Z8o7oUyjBk6xMFVDdAngbV
Lpx5G7HoOiyK874FejGnLVwBmu2uUIslc01GaQ9Icr/zepAks3AQfibahrqMoXzG
0apk7wX0RhBw5Qeubz13mvpToZ+ydzubt9vswUsY83GciBBkUnj3QIEQsiTk4tkY
vDp28Xms6D4O8rvFUvoVILWj+af+grNPr5heNsvZLgU5goBSRp71b92zP+EZ9k/Q
+ckqvKpoq16Gz12Fcl2X7xEq/NnYWwFg5uBJEAOpAYkggfU+c8A1oJ2Is7+7CAkp
mSujNXc0B8Dv/4jiMrJJxFumIbFmPwlBCI8q9RBs01VqAZe3EIqACg9dsiGEycZo
chMGwjb7Rkp0bi041/UtUGL0D8rltKfA3kJtio7jFdeaJJhwn1vlseMHag4XAWOK
FrLvm+vk40AnJnAGjGT2Fiv5+lEJCyM+oygenn7ueqGLNMF26KR3NYzOdMkmjXua
p3jS9jsxINDM/JLqVwdOaV9D0TFyZhcZlX6SoN236VNkXRH+1UO/6ETtyXbWWKKE
tW+hu3tUPVZ5XZhcbJr7O/Ad8RC95r63+hVlDeppyqs3HLeqPv31/iZxIWlTS7Fr
QZxQxYe9aFupANXgwQ5KOHQ/YC8kngrXzXtNtJjnHCI3QMuqtLuVus3wxwn3OVhc
d1hBNWX/jwx3ydpGmE2Tzxs6Ga1qyGZlO/4Z0teV4jlHwiU23E+S0HCqZyrzoyy2
NpyZE8dQrl612ZW2q9YKUaokXxAYbYnP5nOHIwk6b3lJJH3FJ7JEpEq8D31fk67n
teYkx/DiaUd4pKHoHL4YqZdI/Sor8rWC7xWy/Uq+svCRYgNUpztsMFXoTJQSjWVN
9DpSczpIilWaawDiqa9Mkz4IwT8uqQhztkvyt9BOFLtLs2cMZWW48Z36ZAR73PCj
H8L2IKaJEJDkI4ixIYvPKX2irdtBNgPI6JqFKJZejBhGraxvI7wBOEo2hN7QfWKv
BRE3EuggiBkQWv4LNKsaaXeC+V9/geTr0fA9lGwLZ5FyOF+8ZwMa9TsVf3YkfQ1N
lU2V8hh7XsiiRr8U5MkvqA==
`protect END_PROTECTED
