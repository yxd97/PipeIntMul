`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fJAsUxJZs8mnhonivXz39aN+hIoheRBTGHbdwFQfr8ngD8Z6TM04l+P1AilLeKM4
+xE+6/+TXxNKDOJVyDEX4zIs+2xZMllvf/+XepKYgrXerOS52CzXaL7aFYSiwnhT
1Nt/BOfhASZ4oJAfVIiyQAcYh26915FQE4zbXVNbU+eqYE/U1Qlp/kbZU1C972bI
cu91Wl4a4cC5v23iYvuFbY4AWTED/tmz9gMFLCYoPH4/v0XUcOJYM+93cX7Uv2fM
EdBAh+1o7TDce8Zi9s6A3OBfYfguDFJ/cSBcGcVDY+2vj0pDi9tUYJF0qb1DOwZ6
LumAJLEQetciTsZGmNJo1g==
`protect END_PROTECTED
