library verilog;
use verilog.vl_types.all;
entity latchsrcpld is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end latchsrcpld;
