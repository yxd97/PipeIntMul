`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5qhdxFvqWOYn1ds2wnEnkSRCWAA9PTp12OyqDrqj6SVcrGsVO8GhF1JZvdHKhxnf
M7CFcM6MGTwwJpnGlanrhYMyZS/0hc5eYsmW/mfOWEDRq+lSYZ9/AiwGQ/V/NrjR
4y3rxYTQy/MKn+KTTzozQ4K42VpH4Rm1HvgYfz8airdWbPk3PibMmmhqEl3tJi49
Gxf2YGXAeU9gmTrxw6vu5lEFpjjf/a5LgRqiU/+hyChyoO9+EENg3wuDbY51zhp0
EgQkFTmX6dt1oxPbE5IX8Jy/KTNuZQtU3CVWQcd/Nb8RfaK6BE+BUhPUXBTsQHOE
S906GDEVDhzz377gSxvvmd0ytRL2tQFN/ez5j4jJ/YJQr/GEA2U5mp3mJr3adPrc
wEU+4z91zL87uTAzdnXtqBVlyANzae3EFvZ5XiBZyXs=
`protect END_PROTECTED
