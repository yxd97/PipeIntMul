`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M1orpeKuMkYNJn89NZEnxj/fhWF3cVspR/q+KM1h3bfch1ShQ54EcuBUX4I287Gc
O9yT4Mqinjh0e/qCS+EYXKn+OHvh5Egb+FkDoIeabsrFbSfS4eXPouqssbU8nEPJ
8VQyoNpVF7GUbvXu86tLaG/g3zNro+Vd7AWo/78yYEwdUettRjEjqiGHClBgjZW+
tijoihZri+y+7OAo5EcVzaF55C0GJ3e7FCD6mIvqgw3TQ+UxRQspQznpkVfLP/Q9
913uYSe7VJPLbxB63SjL6ZH/Az2qIOjSyCLcohCz0KwUPzYeAPSWeYLtkmJwMilV
KTYhUoI0TfAsug5be+Ucgbv4XjIpyDDe2UIAwfjBNlRHgJXtxgJXXy92O5q9iXky
pTg3JVD8vmHnslysC4mzcHDOb9mBQ630R/tvN2v8hMaKb0YPasTP/Pm5M+39LQR8
rHGpdoD5eyAtQ7iCoRkzSIiBgM3Ody2s3ybDbyq4kIYtBFZSZexT3E9AtbPOI6mW
`protect END_PROTECTED
