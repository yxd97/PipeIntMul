`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eP/1bKCk7wSDcPlOpWaWKnLNf+QCsNQVWtEdJiq3avcggwIn8iPCyZU9j2jWOkgT
SkwaDA85HHucB+FE3TBOnIkdFPzXIZHpZPsiEMWtSTjJgdstkaEKz4t6nsDRrXme
2t2JjbgfopuY6pSAKR9lX9iN6vYXbnM9w+PSKBG+1y9k/D/Sij2jCVttIeR52cyn
Ex7KtPQzi4Y8TZHFHznseE/hdL7VvxSMVHUhgnq7ECMqUPmY2VwUY4i/G7pKvJ2t
MIJdHFlAlfY4PcQ0VW6pIty8q225BUUuDHzK9wK6wU1b1Agxd69dbytc7eW9dXwq
fgQeaJNi6b535YP3iFVeMeSn4428O/35y2JBG8gIimft7lU2OD/ApUtXA2EQeEw7
uUZuNNxYKSYs+aGsnjNjTk60FdpYUvKzlHSFhIVONuA=
`protect END_PROTECTED
