`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCzpFqqVfALWGYfq22pT8tZzMcJzHL/5+mazW/0ITCtlmj2uicPrp36Vx6QdS+PT
0JmEBxmgKm4gQArel9vN2rPlSVTDPv8NQRFT6FydOfs9jB6EE71DOrbTqQWflGLN
7+I8Y+MAaF/Hx1XRUGoQzhTJ7l9LQhTdZOsgJ1aiRRZUq+26PmNCd5knHZdXyNs5
HBGy1Ma3K+e00w4+DpbOFdTfXiXWGuWkJRoxcRlwWmMJA5bxFD48ThkIY7bcUcK+
4I4QJzQQHYa7TX+ZiF4gDYiqhg3cYTLWC8+Bk6s/yR1+cawvzB/nsy3JkmJGXnXz
KXh5e8Pf/e9Znfa4XN9Cmzw0MPq16MMaCxlbgIhrtrth4OUKKYuufJzfnzCXeg/2
70iGCinu3yTddFRDaaew4XUk+gTE+UHzfzwL4dli90GTJ+gaYCZdENHSTC2rLCk4
87qD/vdXBoogtSTqel9YtL44X6WdbfVaW6TKQY1S9WKi9tmS7mqV0E2+76sCe2l/
NqpuiriIRKxnnFtRYOsQ1pXyNoZY5sK8a3KqThClJpTJxCwi+FdUZXRmPrTtJpFN
LtYYzMLhXhzG/9z0hfEO9zDu3ojjqFjLkAl+549hrwcMISebJd2jUsLJhsKyVn5n
2q72nVqss0eEhrd0M25ZFTrhWCi5bq1UiaPe9WVOjHNYG3rYvzOCs7vkzxY9SZVz
6wVH+stmSAUOySim8irCxBbRZJOUakfOhPwjEG7G55VGs+M0EfVX/HtHuln6KchX
bosU+dlmDyQCa7jT3Vncc085nlzXQm1V2pTiU9xG6cfEBbhynrDXjpAiVn43xP4M
B2QlDNLbxet58Yylcvhl4FTxoZb1bYa1w5Q43GNZXM5Lt/EvBkDGbf9v6Rgnu/TR
4j8l/JyfZMk0T8eQsC+rB2R++4aqfrWCnsxDnc35s1nm92wQxXwVHK9csS1I2dSr
xRZVkmNaDhWE62S70HufA9RrPwJqWs2Pqf4EMdG39xOE2AvQTbwcYMPcE5mxYz4X
J+X1e4+wl0Hi+pQT+48QB2XuGc4cjnczejg93+Lu+eAuU43PAi/U9nvPZ966hRYJ
6Cs/W2GdDWPWxlIrS4AtAMIxtJMgg0KMajl6wzgXOcf1r3kT+mASyTeY4xDHLBd9
NDVRi+yBL6Sn3zjy4eYerSqAxoaPUu/XyOalqpf+CoaRh94AaGcH2dHF9fe8Xe6s
0guSapuiQgx3CiRl82kRgcB1OQiP8ZUzpyr1Ccn/jNQOvPTuvHPdFvRM02dusSVX
ud6PKLJG7DGUBXMFna19Ja5/CPpsWkXzLtwGvtBdLChV8qoRzhlS28vzJesGmMjo
EgaZkKUAMNoctZwHS7YjKrpBQtRFhtZpvlp5s5urT+RmLhpRbfRFuR3gNL4kQMfz
ANJ0NOM6Dke6to5Plm0K6dkSNXwxvxgyNV9GQXKI5ASmXr2ASqW3LIPJV6YgKPz9
4xAq62IlWzq8YvWUnjP7P8IRfpOPRX85RE74NTNuaVPG1cXE8wd/O4GwpS4XDWut
teSWHP0e7n3SZdZtcy8/bKX93TgvyxCs0CED+hqo4JSjnCjq/+xEdML5c4L7YBz+
ZX4WOX72b+fbaOSQ+LbGsP07pYcf5V5Z9/+Vg8gi/4LIIluLOjHI7I2KrQ6adkwe
t8pCedi3JrNJ/xKoS5se0pvVPVS0EiZp49wb52IyV3Q0mnjlQWjlzd2flnpCgFCb
fK9285thaH/1FhTIijCwYPLPm0dY7O2wrQXeBmjOdIbNhoQWcFe9kGgTFS/NgoWg
LEwvrbsVusuu9WQjYnGyBJt7e2ViW6hweW4qCvX+zL40CVZSh21gTbRkoCMjuCLY
jReV6ineR4XhNEWiwIPw1UWvsLPxvhzUqQ/iZ0dmmP5WT37EVNgZioPLFxhXE/bJ
/HBEEFMALq2hIsAm8szHWIxOimOyaYu3ZWKv+HuhyHdd+6x4FW08zDK3oFgat6nF
uxwdTBUJx0+W7JfEfmJsl1/TCuQ0KjU+r9myTmFmx31biGHMUJg4JEWsyBt4izNq
HzAsCBKcvuLDlcExpQYt7mCT2uEOKbzbPEzMhWOtuXutG093BygUvSFGN/wQezPl
/69plz4pLRyGjWIeOwOs7anYu5tl1T4TUua+iabnIchAiMFCRE2aucxDtD3tnCX4
zTyYWry5cBJBsYQ4fKosgvl0QliECo8FQUZMDqy22ICNcTQCzsHA4AiPOaplsVw6
QGihJhVQ0rZm//Kr6TJep+W24tcHQG7uCBnAWvHROHuQar42mWp7gdtNtGeHWzMi
cqlTfkSpwRFDx5jG7E3uvkuJKd8NjeZoMwpE0gwN6KfmcvTz5u5qmA47yCP9yRSS
soDYH8Q5breZsNohn6cPy7STBIoWfG/h3mF2x0St+dfTfweQ34zR8nY3td6urHR9
HgCBowlk4eopzALllOseOIUGAcMYtyjeJ3oaDTbamkvNLk87lKG28FNDIwRT7hU2
E1ntficyY6TafhhopkbQV9C5YMMwpJrpW1XHjZNkX5emjG0bLqD1x+VgLFgFDn9S
t3pPLSEB9tssNccv2+VbpZkkQCIa9rf0JMqufnDohB83UVlDmnjRTu3ovLaBc8Tf
gYLLdySfhvRmLiCOQNhYV2twfy53o8AE8Syl8RelArrvz3g6Kc2JOpV+eoRtKFx7
Xc71qTxn5jHWHZxUroG4+OkCxHPMtYGH0FS/N8VcbkAUgr3pAiUo6xmY1jc4iWNe
jKdUcO+0Qp0EZiMPKqN3CgnkQpzxXT2I0Sk5dkCsBde7BcTE6R1ujp40Z0Lx/vjH
y630pyWYjDPovF8oHThD4dJ/tRUP6uHCQFCsjX53UCX8hsMMjD7ju/al44j3R4ye
5E37lWcLMMowWXQJGs4oRXwTALUOH1IqUpPuL4QfZvSjtL5AAjJY+6yfbYL3xqvw
HRvIp81snguWJMLLGcyTnWv6Rl2KCifvd+WVCzAbdnIYhN5sadl1ag9Nk266NPmd
lPE2SXD2K+W1o7YS9Dc8XizhnHkg1/ySkwsx17E3M8A=
`protect END_PROTECTED
