`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ql8iNLu3SRGwA4QMfOyIV91yJ6Z+mUIeJ5yAFcibZppBmU75KRljVNrA+UzuErXS
YqEJXF5TjnpEQhGhpmtMXdVeVEoB3zsGdiPnpA9749MVFNaZ0rT9vXTArcVP8sbz
q93AhuHLyrbWKoiD4OGjWhzf6cCRfpaGbLdnqwhOep6Jxia1mZ2Rx2WUUKK1669Q
4RGOREW88TmsBu8ufX9LSFJyvlcINvXNE62DgCad59fERWw6qoB7XglpnFhpwGjo
PP4JQ5asIv8JOxCV8JqeWtE7anGNAQgvO7EwqDR7axeNhYFR0nXEp7j2Zx6l7U/R
zXZrE9wUZ/G6jDkmgkHvoT7CY9HvqRXfrTZ6ikx13VZmKFo9zNfgsxCxYxce6zE1
f4+XQUmnkLmjLkPY9Ft2PxqCOavtNLFAKEhXYFXMgMYRgHwwD7TEDGEiCkd9ZSAi
KEhDWj8pwAcKQ5g88dY6Ds7znRI/brcij3CNFnCs6ilu2t9SdYMFGFWhvDpju9e7
WGwQkQGUNyEfsAhGKWf9zuAtnw95j8b8xBq/E7ECG3Di7u3kDjaxyQ8To/ekbMYB
G2ahkBM5yzH6X0KWm7MmFagRZhy3rrBkoHGynI92Jpmfn89jEzkAFP0U0R1EaW0t
2kHWtT52I963mG4SEp0YGIjuxopUi+tncRDU1S8952mBtXtKM1b7UurJuNriTwtj
TsS7w2G5iAHDCBXsgvfj9i/fuTv3dkcXf96BZbE1nYp7I5eKmeL2Xpl0PcBwxxpc
JJRrdEq+AP549C6Pa+lR9umNzdcEfviC1y84ZyX+9oVBbevqUzAo3I4oAaQ80Sub
uVizi9SBs+Gr7KkTaxkGkENaAIrsc2JQmA+LgEEAS+0i+Tf+ZEA+PWNiriKMO+TZ
Mg6/UrBAKiejNldvE1WG+spWOe8ZemMk2c/ySU+mGTnnafhJ5yuuTtU35TYGFiWh
loeRfWqnbQposeOZGBxswiA2gPvw/V8yRMy/eFnZYVJkQvKniJR9F61+PKKnXYXh
mPxY7tv+Pf8S9g/JoaPDKtccVHljPW7vDPLuFLqK3ba23f2CJS2QvoZqaQGgHF15
Wd+qy0uUj1rdf/Bs3zYiX01If/TxKPiSqxyN+C4GQl+9KFByCGbtdL57zr5viFfN
S6VcD9BCYDGzWc03Zgnpc33JNji4fNMRg4aMxQCpONsPKxtXrVmjkAqunYlji5SK
cb8Zd6rBzjKMNF7ThQWs8nGk2Y6JddcNSFe5uK5PK4Km6quwKQ4IXgDBZrtNSRP4
VNbuXqZexweOiEvRoOsNY8xMTPU5YTjTgxpZt2qT0PDXOxUqemG5BP/Tf+1RiB8R
JkbjOlPk/vG2lFjhJkbqRYiw3UNuLjHE2Kox9Lp4glSF9gqoqHGagz9ovt9Z4A78
IZanOM4ItDdRDAilYyPhSJYnJEZsuAjer6si81d2dAMs+mFAjGeyl53Ajl94368U
LiuNB50D6+PwopFUrov4nC2MU/ltDiSYa8T/7qM7T7BvgGWz3NxccQcji9Z3Vt83
fbWdsmIis6NPeWfl8G+UjysTLNZAVhBOoNJVIGpGSrwIOnM7CaiKhWPVaFQqrLjV
IvitsY9bOP7GAAgMryTktA2Rle97uFBNqGgFt5rXq/BEXGGFVHRUoIMEP9hpiVD3
Sgc6N7VNMkt/GYuIWklf6sRKqVrb78iZuTLWaefTDYr49gBGh/c5aEfYHIo5wcLg
tjZX3GILnJPUQWVSnDaH8hC1ty54gVzJXXSlu+aNG85RuWDjXyH4NaH1GsL17B8S
MhI4ZpMB+mTUak8y4vJvQjyVXImLGNs5uCFCAOtlHX6cVJLiGbb2xP99gaTg6QFl
mZCIz8iMms697fjm2+SyIWB2ODMNlLuN27KVuXkK0oFwm5cg8mG4AvQADy/et2dK
wRGkBPMUhaLUTMmdMxzYQHsQMqp0rSqlestE0NEgAK8PNQd1hCWnmcSkK57iA/Tg
we9vNyTroFu4E0mE9RrGvSkJB6IYQq5edlqlJw6wYSnlMrQmqPVQfebVTb+i+HrV
fW/JyZuKY21MbWtkE9PUWIkl6/GmOPn4ofwLsPwncknlWteE8QiSWgR3aj25vgOL
bOSz2m5eyFTeSjRTFCo3ZhrVMuxKPa6iYkz4rh1/h4B2qcSQnUyKms3YiLNNM6hf
5akVxL1DchdfxO5Bo8ZuR87f4qgNteyUN5k42TgFdE+T6ANe3bzxZeRtQnuvmEUl
M2OGlf16aoyhJPSM0xOqG3s98QZDNUgKGyQHfVMXgr4ehoA0pHX53+yDFZWkJ1pl
EwEuhYdbXTA9y+GqG1n5m3vLDIosTKZjL9WUsJ7l8CxyUlqHHnSDmNjOPpMHuncv
mkGxLs9gYAV6qxVhEqEiXLO8yRt1cHspZF6kVqEPjs57y+ibIIYvm8/hwV3//Dre
mO8LZct31bO3hLT28PeYMtK7I9RYWQsz3Qpyxqgy7MPe8Ayj4tqNbCXNImkkEows
e8KuaoIs7ZRcg7mQG4ep4n+aXwI9XHb33zbRwbRUwCbXrClS7bkvNchlHN4tCc7C
VMCBx6elXc2uH+nQPC1bf2/rB2O+HvszdOuP+qZ/+nAxWNOpbTQN1oIVcgu1wIx3
bi/Dku16SQKKuKjYwZed9X4r0qAGFjhU+6OMX01jr4bQZgIAlnnJwk2kDIXsq5Vu
3ERg+XsDiQIptcvOrjDX79kcqSu5pov9WDY2F9AwIQ8PtRhW97IlyN6WMaW2LCek
h8fxrjMA3IDZOSYeWC+lHczeXUGTP6ygixM7gUTOG9kddB8lu1WfjtNJiq9Fx9zc
WwRlaUU/5Jlft85CiEO0YvtEwegAg1kjacbhuur0b6DkSh0fYaXitTYNKOxnxSq/
xikYuWjGwmZTUpOw485l95apGeC1i7/DVsadpnbHaEA/Ua8lVz6/A3uAfFnxu2WQ
/EULfdhYBHScabU4u56z7A3HgUQ1GYg1FDF+LsK/phakP/ac9yH5sCxYtiXLBO/2
vEhHGjD9TN1k5rXOd1qYJPsNrEVcqMOnInkg+SxN21GvyZy17jPABduS8Uaxu0zJ
hz/ZUuHABZhFDoWhi8CMYF//avPogUFR0De1uGEkIjsoy6iH+QF5EeSP91flJtvv
UUYaILqMa1XEGrW2hWYLJn3gMTT+J6ykneIWEDcIg2pPWjPb24QhIuztZKkfLMZr
gD0bnfHooIURM9CiGcgNpfPYtIaYiN8XOggvFrjThBxdLw0O2wwAiFdq4A+C54Gp
/1LyutMDB/K0yfX2FbJeCfXswQou6UQck5ZHtZkU6ZEvsE7hG37KKK2XySocpbvr
Bdspn+tJx2U6KHjU55ePga7myzBYwzzfgO6tM92Nh4IPGATIFUOS0oZK1JUH5YJp
GGyJxqmCOIZiY1sAWoNqWEvitsoexZ42d92MJUPKUMd6c8ES1kdq74VYHJycQbfO
67zGL6MPbQjjd45zbsQ8ccNm8v8t4a6sZMs3iJPGBuvCBNw3xBAF9LbmnlD9H3nx
TlQPD8RxdqskSIivc6FWVseeULy1AE6jPqYBIx11A0VAdGOZ1Ak6z/qs/+GFNjnd
FLobANE83f+aTJ0TKbisQqACqf8lsDrgRcvby5INuGY+e+g9jQCVo6sOW//CLEvr
X+8xkNunM8oSKIBXfBaKEwFMzY0TxsBTXLh+0oDB5cCsoFRRSOkyKNOVzZsgTeRs
x+1WIGTxEzeGsfff1GcDkVoiLF0+S5soRhJbopZUApSMBx++bTiQappBQ/9GWMZC
frAVFp9P/N4ZMHnjj810nXTZrKrgnqZyxSEq/jbc399M0v/lUeDNfVR+8jlgikNY
D6cPTT/kOsj6/oUhUQ0QBLQkccY4M2RBlq8gXpWYwI0jeYQCvJL9bK3WGYC7h4XF
FakwER7CxGUi242Sv5XnMIf38AD5l5bqqlFh3NwdV4xZUETCNkXTL8Kgie14axqd
atDn6jvwN3EuyWYcD1QkiM5XDwRFe4l0njtw4VNl+ovdatQ6LbtqalRJiK+VlNf6
aVlipEI3oEGDUICz4yM9Q2GiR5+sXzEbLvXilXsQPX9dK6r6B30CEEtGB9HKqq36
uWnJZeTtbxWjyRx8GeztVFcFV4wXKMeoy6Ut+unbso7PPJx7qlWt4QVZ/9Qxpdrb
qsaEBhDW6MFxdZn0sTPoTbs/n76I1DQEGF7oO2WlW5ClO3HE1MXWr8gIqI4G+qs0
L5705jJjLDPQYMSxdL9jXECEA5DotwMqybcsEtkW7ZBsUNIA9eewq4FhQGFwn1j1
nx6aEqE5zuAOuejDRMYRnBBp3/bIb3SGhZl7r/MQ6HmCZtm0HkP7k0z2lZcI0ZpU
kEsBCYmLU5WiOal+ucK7cxDvRxpKfYpJa3Z/erEqGl0fs1oZXVeSFW0qON/81LZD
NQlUsFx4VOQ6aU/9nw86NRpcf+udVY95AgYv9EExOviMLQB3+54FG+g6If+9rtWl
Mfyq7SSYQpNMi78FA8E9dj94gcpALAiLvTz9Lzs/zwBOfl4yOGTJjwxtK0d3cJ6a
aGCdxI0VcsEQajGGwyVFIc1VWIIta4hGpkkIrj1ZI3ZbqAGU3dBCmwMdLUyC45nq
owchsJYF4F8eR12SQfsh3UCYcy9aA5uYx5zIhPtzTXxO3UOH8GicQ5IbOfeZSdDX
5e4qz/5RXX1SXs3BeswyoxicJ0G4j/pFlDHpATML7J8nWkge82/AqPDiQDibqni8
Llv4wYkJMgWjjMWvSTFHUpSyvYs2r0Il9iYfo4MZd+xaQiC8bsA+pB4YTEYQQUF3
00mCNNSA/LphCWq9ziCOKGDi6ngzJZQ4+zwRPOSKAqKRmpJ6vHAgX76GR6FePrOc
jAsHNutDDEE/znM0KBbbZ55gFf1YJgSFeQ9GAT9R7bq2uqmvhryikpDpFfLWIhYX
FBsrSmzNarhElBnLHriBYD/3z+8wPzjEuslYRuls8qnRFWq0+cZ4F7F1ADZGKRZd
K/ledP3krG3Q6GIMTzoZdLidIEALysakZ85nvLpo8824u+txdIGtWd0+TXaCnXGC
lCD/ENvncv/+zowA0dYauF3IvTT3pgEknPtN2A/TjBh6V5B9UzgUWMgA77xJdowi
ZBmId9an/jgUiTPdMKnxV9UTAHeOl+t59k3GwTiy29GoufaHN8toBT3xeJN5D+i1
brXMTiUhxsC16XQrosIFFr/jrQXjgSh/r2SIfoWSPMLvQ/yjk8WlDz1T7KBuJ1yS
yBtBEboAklJFpnT7JaT9TcmPAbA25S3PReUjUz/5/X3DY8/1fAAQ6qrrnTRp5hLA
WO0vQ7xfAiVxNhvSNJYFIL7XhjCozeLfVcm0RbKXaGRlZ3NcY78OFDbYzBbKqFm0
/rvLjdYdJJ11Y3uejJUvHcYl/jvUnz24JbokLOR5AUklj3Y5Isld0K4SMfj60r+V
wCTmisxakVgUyuqCfRdlrGNGK/jwChttE6tNUOalEDlmVj7RQ5FHHy4b785lSTPM
C6ArYggYv1UWDc8X24Pt6XVXKqQPIGdCtjl96A/HKL0MISlb5pCIttZF1/MG4TfP
A5Kt8dNfYmUs0BiuJphG306kRy2cdIL+3qlLbRkjY1RbG+bwvQIPg8HiAj4Sr/g4
8kAnGhVyq4TwtHo9/txVZi9fqA2YxMfpqoOH9RTuL6tO/Z9olrxcD+fMwGqiNGdJ
AywvW7KmZZnH2RYZVIiPylU90GdCoWyiw3td0FlU4OaKw1SL1VNsrELgh0wOMnry
i7xLEWd6B/xyctRovaREkvjSCFM/qMx7bY2Ow0fwfVeyPYKjS6uYuYPqKwLe0cZB
X+UpcN7Y8Xt9mwYkC5Jp5qa0CHea7+u/EjfoEa4DxSHMY6GXlWm5vyY6naey6yux
qwTkPQ02eeP2gkgsEFheCNNewCQ1mRB/SiACes7uAauhPU/Di4dORM16ZvTalcdE
KkEauiY8BJS8A4gsxJiLo51koYq8bYeKGowxV+Hpe+7C1GxrpPmyFKijKNzjDVJq
Rn/WQrO7jMVjlyP72JqQ3uMI6K+tnPaq+57HIVIai3zU9GWqiSGqs4cp8hiUm9f8
bR4N+8sjDVBhYzjy5mT1PB3KwbL4dSdG6TZeMl1zMU8SwtbY09JgDdShLh709TND
6BL3236+6udLpgtgOtf5xEVw8VXUWgUY/IvS0X55GVeEN+xPaOQE7jyTTkH6gwRX
MNr8G9Pt30TOHh563m1wuBg4zH6THhesYGshQAeDDn8o6z6EfFC86Ff4A2c/fK23
TujppPBH6IBZPL7b36dLgYzvAJU6Q+l1wzM8+EAXkJ00KY3Yp8MlnVIIvgS44PdV
N5kYCtB5WdrTpe1zb/6Cn81Fo1XMHYryYx4D2hcYrq1v6TZd82qySw31p4/tSFjL
oWVSaHvZjYj536ODVU4vEyxk4pM7IzLueZXx5AncpZ/M5t/TxxBNWr0WjQrjRw9c
mhqjgHyv2NG5gZcmOI7jsqQ9/8ij4hEcaAgxDzrOBc/S3sSkoHGkXJbUinzhAHTX
eq/OlK6hiqaPgf2ID4ptjau6yVuuOrIWVqMQu3IoYdjkDVZ1CRPXDFz26Lw/k14Z
XuZLtIEyXSZResWFoZ/lq9mTiEvK5LP8Vq8VFUvP2W/Qq3qShB1I45W6cR7I7385
qJl6e/ENYZNlyxJ3WJPt9U1m1GEFjWqxKaL5tM/duAoKjKg7pGmJUmUaur5LjAST
5OKMCzAvhpC7/tEBB+vp1qNpdEZ9FlITRt+vnKFLkYgWjanEUMG+k2pUtGWTjnI3
3p5QGNQRgoDQoLeMqS4iR4pkh2n9BsXPTY/NKfsMVE71tLwVzuPGGAV9GYv4L43T
UGiXsMQqok9TOLMCtjA4mdhSY/6tZRRil4QHHnsSmA3FE/ICLqHWo+JLZrL8f7dH
iMg99euzNyHhRK4MbUsyTyURZZsdHVJD55cwjAdHdrSlD9+eroKTU5nBDXQKWZD2
RX8Fwrl/bnjr7qeCHUx/lAiivNeUdNUpx0QY4pndKxP6sDhV4sQgVvMtwzB+pY5W
kNLffOdwF9/BhjdxXvJoe/MSNiof501nHjlhYhg0SjL8UrglJuNzsFhLIH63tTbW
74OlNq8svaIWotFDULf39Oi5kJueB2Nz0403Mc/UdobLEFW6HSxrQAFDXf3mC4fH
oLe1EMWR+FQvQuewaYS6vhSVmm8jyha4SdONPljIdtcYYjNPnEtyZSeFwRp2DzB+
Un/7hgQVCtqn0pC6m1/8twjCrYlP9OGQdOF4sqmzwRezvAf5t04nmQFYkGIVcRoF
QVK4eSiG0BKv4g3TRCeYAoZWefs9ILbu5fKPAIPKFMyFLZd7o8Mqh3nrWLqnF1yM
8gXDODYJVWuEB1YkiO1t6JBV9YyQysLj2vLYE7B3BbjZCvkNzIihp2GcjGA3rLyp
XheIQegil71gKDqG5lzuNBRIDZbV9QcZNKVLMnpTSsFO8ByrFkpFbtZaCQTVm+6v
G2PUuRWihvHWXCgoO/uwSf7u2XehhFpa/GQC/UN7/OAI2BqWucy7ZpkDrDKf3EGJ
w++FO3Qq9hYjEP3aNHb0/kOdSjo4YFefcHx3HYXdTPRFVP/YxRE6NnQlEZFP4pIZ
PkFrQCytE+vs3Yk4eFGh05iAMu4UNp1PDJlR4OeLfvK7IkHp2gceTqVrWABVc9Yt
VAl0Mi8mBRjgmDsrmCs5vpSMqbCagOhJOthbaSD0SSFBOQkQwY43oJ9yd26JVrIJ
gnBpxJseKkqKM2UynTyqHmncUcz3NGIBZyzussYnl62Bx9v586HSLyLALg0FIhkq
Wz6zs2axOkXKFWtTGDAozp4P35qNZ8Un5c2nWiTVAy0Z7prXjrGspmjvQhAinLep
EGzlgWai1azDcUEwSi4AcfZG75b6US6unNX9adci1mnm54Eqcd7isGDr/q4Q3jtG
8GWB1bMr5L/p5QIl7xYgxH8N6rwzHWbtkJeNPyUg6Ce41SVEjrMCfA10Sr7np24L
9FMOrZrD3v51bXKcqPVx5dloKtVJjfjwD0uv71cWszdLCr/ntejGy0+kg/g+mhNu
Lh8offPFOXuFou/gCZJ/wB87PbhlKRI0B2fAtFySz69YH2dJqR2+z4KkUUkCT6r1
Ev+zXaLLn/D2MSXbxdQvunyOWAdRPTHebIeSXMQpn81ai4VooZcaqHo+UAYqwNtt
MxTM1CTwlM9ONS9KIShjersBsEZsyGKWQi/Y69uekkRmEO39i30EI4FKlEkTRvu2
4y0TRvjmIbEbO5bWjbI0fmca7cIEm2vQSQV87OhY52wN4IHcStbuREPtZj8OkqNf
bL6MOoH4eabZehmGaYr1hUHbedo1a2gdUN+EvKQyzHeeJ6cXq45FT0JnzHuFuBYr
CrofZmZfcgk6QKrb5bmzP6uqcFD0wfJd2abj8zA/nSeYDH7Iqs8ip3ith6km26Ul
stsL9uVX2hFhugVGKu+EPtMahuEdJqq4MjgW+MQqyunzx/otIbPl3OWTFATlZ3eM
EU81xd5H/s18ZLH+ff3yGztFti8n84qcbnnFhYBNpOiUWZ0rYzFgmUjKe0nBmDKK
8hHeX1epbdGhHKD98kVB8QDFubd0SbpypLXRTUbXH8hDbMsSvTn0dnBAGySh/fSW
DN66LNFPOag8tuCcmqGBUHuvGoA+PWcwXsaIR3SgoHfvcY3wyMeAvaltsR96LNbk
NKMuxl1EwsgFFknxBOr62q/JfFEmXOsHqte1f7O3YX6baQ2TPKJJ3Ewn89168HNK
ZhFq7ZMCkYftgYjdNLEpEOkkOtI9xFoXW9AAFp+QDVFE72a9NcmCX/w23dN0w4Tt
vPHTsQr8u5mObsaYaLHODFcypLpVqs4P3EZ2w4PNLzVlLqEBMS+CMXSXCvObIFce
2K44MGMIBjwqXnrSX5SBQ1NPJnijLiEAO15La8tE4aTT1i5h0FcUCL1rKMcWs1Tn
a8BSq0tWmVcl7Ti/TKnhVsIWM63AT8Kkwhk9GtACLK95AIIR8hKJDFjlE+QKJc8t
no3ti/MMJ3xHFd9vGZEHXsrQGdS0dusglFgA2h319dd4vtU44lD5b0ptOim50u7m
DIaR+N10M+BgiwUTkHKWLAuHL1Y7VwyIFCxnzDXBs67X69Si5jsxaz+h6qOdkK/B
YLbkYv298U60Zvm83gLfnyqfgA14ert4YGst3JNe2VVZKoqYlN7hbk/Xt+KOOSGm
aYywJ8hUHswmyVpymqy7Ih6ktwhhrBD9wBg6GzkRhJWVRlGzjpHhCPkIQTudE4c1
30fU4fyxMjI7jiVcu9qWRbB94Hh7yccvM4N60voYdkq6GGQ7kqdg08/qF86bAhD0
8yqzLwwq0eiMlXob6Yks4RYAPkvzLVhcrld/VM82RkGqeLN5W0rJCQEht5aRPEiH
x4w0skYeeA7p953nK9iGWcnvC4LDGY6oQ7XxHcdhqGz3UA9p+vUH5gM/suD1Jnlv
+9Gt2lv5wU56yyo37oo7gV0QC92ll+qwdMgyMKzOQYAWMseyiDZa4yvi01T2hWxz
a//TcD6T0BiMKOUQzM4BZHqjg98SOVoejN//zXiChPJ5Nv20bEcrQX+R+PG+lO7P
2iB7mz/VmEh+6lyM8Z5cIdqTPw/OLvmPqISgaQM+rbuS0AL/A7V8B5HL3nxQNcZx
d6vMAqytrK2VEUW0e/csevTIcdbhLkucYyTlCiN2jHGewjIp2Cen1ITNORj1CVwv
Kc+kIdy+0tlu0hPiwDtK9BdIgO2LzyNLs0eahek3gKRJjBrXt1DMLUnjodK4BD9p
g58nODdcoiu1l3ni2mmDYzwGZ/PV+TlTCwbzy3vFU2qBKHxy5Bs+Z71POeFAgK3A
O2jtGIslEThCIyBp1VC+XyrYqkFVCmeo47dSayUadBGRV5CpT2JZyrVyKxTwBrf5
`protect END_PROTECTED
