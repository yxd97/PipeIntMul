`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUCZT8E5cI3Ca6oOv+jQIFAkag1PPxpbbSAG5brrjbQWjfGAOZCxQZMEL9AD5Nkm
vnF9YZCXGwheOk16ZhgEvhq1H0DVKGQUJlRqA+StFFVkRvm8BueBX0HuKPW2J+L7
1V+rE4fW92njHcc/2FdXIkc1E8yHqpZWg6q96V4mlJnsPkdgmT+HJMWmrlQLRCjV
TvOM2bENSYZgSIeQzrklzPoY5XpcjQyvJGaxtlk9AiIb253K6CANKUt0MKkidcM3
BV2NE7GbY5q7vh9u1/OeZfJNqHHtQEa48TdBGeOwuI8roBaC1wEunIkcsWXCruZ5
oV5lMaFwRSElj66O/zoCqtrYo744RNsoQQ6iz/EKB8viMigFADvA63j98d+TB2KG
8u0lV9L+Nc2morshYYRr85PrYRhZIgcvVsWKyUTJvbOU3NUYwXFK8jwO0YNOVmgM
pExfUfxBR08ecyInBAgNtHoGE6c46+iSuEgBBIfcTG5UwzDEbOe89wbCiSxr9J0g
gOuMTtEjEyR2e+4jwRv3oqhYv+Y4g+cO4D0NLEiG6k2jJTXh2Q4E13RVNNco87Xn
O3kFTa7YdKXvZB5H7wbHRvDY3h2aU6KclCytDXzxGStVHa8hIaDYfQiRmsLVOTTv
5tjiUAPeVT1ajcPcwpqQIL7DpC0/PvDXhW7HieNo8/dtNq2Wqfy3uUrL7cKiImPy
YXo6Ms3FybNLm7BK0dFkXr78pO8XsBMsSxQm0aJa2GvdeCfwZg9KGsitj4+VqQ0B
qg+oJup8TYnOKuuNVXpw+GANXv1HkUyXIsaR0nMl5fHg0dEpOUs3sbEvmH0+0x1a
h3Ra3xUS2uwXu96s9HCw/Co8z0a1knVG00S2rH4KjGR9ghSV71hn/hadkU1yk7O5
LqS0pZXptAuhv0M6jy0S90PD9kcFvz4VpZpFTtBxI5k276rgLUXQBleYp/rcqBIZ
vDo0pr5JToUYBbyLuH5ZHCYvRke29ankDiy2pTXaGZJTTM8kdeMGvS9zobulk4T/
WzA29J96r7sLe0329p6cTxjmYmKfIOZRMQgqXLZS9VzK9bJYQY2EzCrwtRgHu1kg
OeKEIt3nPhZbLoX7HXfg7Ivg052qMffkusnUxbtJvypWfGQsWBijIH/XNK4S5/Sa
DPcRj+OHZZeliOebgN+wZjW5QCYFJlLFFbiivyhhPan1In70DKLnO3yyKsgbehxc
/JY6gqh5KaL8u+rJZN6/DU98Uc60suw6zLGOmigpUKGoHcf/696W/2KlETnCeDLK
vcYKZToNwFXG5Lw5hUV8xLsr7Nmk747WMgWfL/N4aSKHNqiopAAdQn/JkirURaFG
GqpsQ3roHV+dVYwzxOP68hUdlAw4e45SNaqrMf5exDRUlCUMH6nsWQjINIn5RnRM
wIpBmOOkdqpg0X0OrbJwBelijvhw1co5u+Rack4/tIlzlrk4sRaM3Qns/FCStBqP
J86k8hv4oeYR6jgA6epg6/yywZVgc3GuyUB3e4gbOqMTvjlp/7LCxtmYJLlbcWsO
WSJHS4D9kHQjpJS3FIeB1xap+TGLvDI5jld5xsH2ZyqnRuXVxUJcVHkwrmZLK3uU
+kAhbTzWBUieWRGp2HEiLjo+kzB6gbLSeTwF5rGlQL8sfELiqfm3/gR9YAQ9QzHL
iwyScO1lgjBXI9KEYpxgY1uzFMTJQ0/5eu52tAGzdhjQYnlROFz6fc0OtX5yFBCB
SUl07f3VDJyHc0vtzibhpMegTMUcdqUSH3N6hTf7DumPyv4HOtlYkourgi1D4BI1
6mdb9868+MNalyzGKootRZZEhX9XGBzZjGW0c6G1C09TAqpbXdmxYuvuZt07iBOy
zs6Kfy6Mp/i8DcTw3HyuIcy9sXPeTSXyYAH6rBg8L1i1Bj4xWfI1aGGGEkrP/VwY
V/1RjwZ4SM9CwmFjKKGT80FFS9qOtJXIVk21c6w8YOPtBSKovdLeYNyj99c1MJR9
n8jbBMFK0RRC63BHGlmNm+Cx0gWrr4zn+d3inNdwD5HnyiWhpWTaR5AxQYCN7Ljq
Jf/CwyZeb7niMAFJZKHYlEXHZQSMls0zHGKIc2TreThuWUTb0qF3KQbCvrbC0nt9
rRA4By4guVl5EUVluuG2mJCy1Kms8zMiOS/aD/7RE78AwK/VwoNwyMvwFk5OuGqn
1n+QYRJs/kO7jiP/MlDj8bucyvQNmEJL5Golno9lAatbMMnEulWofUhuKQFJ0IAw
QqUPTjpfawlIStahlcPZkdxUH5AL4mmkDTTcZJCzkHotCgBao9cF3mZO+dyiR5IP
yfROKGwBXePVzTSvgmP+3gI59QWrVUMvDeQils/CAbm9AGVxmtXrxL7cvID1OeHJ
5d0TC/vTXw1Nug9l9QK4jcgQS9nsDuLvx05Lw0qaBP6mR6YkCQAS9K97/2nU8leZ
Jg61jPvquqrcGwckS7qVXw9g1ejYLHa+rHp7+SSDQER/5Aox1PiSqeGWc+/h9kkp
epy8DnwMYY7LScjmH0k6pKJ1gQ/kN7VNYxGmbtyGkKg=
`protect END_PROTECTED
