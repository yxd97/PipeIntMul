`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3HBYOeDhYB8qGEY5OV0Pm9ZFnafjQjoY7wm3su4qJkHzdrXOJtKHawNhRjOySyY
Ix2dI1yjscVdr16lToshR8gUhwFGXJjHwISvFLBc2EOkNwwfSMhegb76cRNyVqKF
7C7T7tyG5kGiN4FFdYeqp5wQVwh7vXWfQWCLmj6sUe7Qvbwh93hVx60Q5WHv8r9Z
YHUDBTfDJsfEOWsPMpgeucxTEopqod4vytIS1QG1/t7Q3L6Zp2Vqm6JLU9+PqT8R
P/9CBh58/FM7Fpj5tOYFkGf7iyevtkan3ZvOuk4/4qqoxYTWC5hmyGxhdYxeIuNu
EBozsoYUpplICyMhnr7GX6Fn2xB9TPMzuqijUThJqys=
`protect END_PROTECTED
