`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GC0IroKLpfE8hTOrIm4XVfxKsxXVp2O9WwjhG5+MirMGRE0Xhk4IFKdiXF3p+NcF
+Vq4xN37zQ+vseoBTOtjBiHUicyqYfStnoaavW0hzaphrfBZjEZTrq2kHZKbdC16
ZVtmnB0QjH3ph/tUZ/NC6bqzvIowMexAyLdDMjT9hsdvv/5J1T/34xASvEJjPDQ5
sFxUK9Hm+ms1DDh39o56UWDvCnyzHLTWW17tGYO9kFVeZ6y7protg9jPEMACX1Kf
2Pzku3phY0LrpHQG8B8TKxpo5OE9dAVh6RI1rQG6vUcs1Jh9mwkhxcb6mw5KAwBE
Mpy6Tj8mmwCvSfXyqZoH39evu3FwOajGqWvexvg4JWET5zoZiXpv6F6oHBTAPeta
bkyLDL5ZK14ieVHpG1AX/elTDJWRRo19UhpwG535mzQkcdLT073lum2JpoW9nIWL
YZa985Pc3XLi/RiB1f7xTwLhV3tFmeBJHPADbbPwVUMd5LGI5knsNmPe/VA15BED
J2LTLCUiyVRurTqU1gkxiHcuJ11+ii9lAlQp3P2R8Nvt6pXZYUT997l9jxQ4THdb
THs4nDNE0cNig2/qLJOZndI8Ie5WLrElIyNsYJ4kbUxJKNmwGNwPX0G1vDm4wZFS
2e3wayPEpqof3sL1wIRgkxN2GcPP7MSGQWdVWXHla5L4askkVtMNF+NBOga80ObI
lkaG6tLraCn4QB+oLl/z9D73y5/YZcEt7I7Jt96UVMQ=
`protect END_PROTECTED
