`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VjdPwYpq9Ydq3Yo4Hzhk8p/CySNrgI/42DFoU7cwKMyChVTeEXT9NoX8swduO2TK
O8TbfSQ9osJTOQrF3jZDVOgFcE6AI9Jryff10AQ3rp1SZvANXZNz1IS4spyte8wF
qFwGlfFuWO5/vZ5qINON7XUqhnXqSvWrQt3Bk+4PUSh+XjL6w3Ex5HtPY+BGpgRx
Ag3SzMwrr8LGE8/NJ7hV12JIEu0OD1Cb6vLUMy4thUrBktNOAhRIRFrgde/UnvPi
LfJ4/ryAXlRR58UfFr+h9x5gcVB3vesIAWUGxvw24+o9c9wZCo76y5sDGPuEXVRj
a60raxMvo/Unq0aui7w4AJ2S2dlo0gh7yesr5/W1awd+b+OmkBnckRLakl38nzMW
ctoRITXqU0JayJsEm4novNq5OB9QfzRqd8wy/AP0L/xBeIhfZhZKdlBYsBbfuRBi
eZLeuBN0aoT8ndRStlBK9Q==
`protect END_PROTECTED
