`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VliX/yYdK50bA+59PF08NlqPa5Ho+m57e8dzKgDCyUb2sYrWq8J7XlMeaQGERocY
YUZbJYuJVSueVVWwxHP34P2EbZz3krHFk/G+EEkfTX7BAHKChAZSoLhZRp5QzkAg
HzTTghn4YDZ/xoipf0wkFdwFwPxEb2L5oKSnOkpR28rVjEG5Cts/nScs5diIfYYL
3rEDht9wJoUd73nCunIC1n4a5laAn7gl4ztpWds+Fen+TzPovfsCgjEGLbB5MBQe
`protect END_PROTECTED
