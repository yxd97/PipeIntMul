`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JjWpbhMaio58+2fek6olNdwjVLfU/uDn458zGFRVuU1AVnSF+ocH04KTlw+k2CK+
MLTVoeLyHIC/fuPYwPjAiJPmPUUq6V7tY2vtSk6oTKC/fF+u7yPt5pPwvfBxYNNV
Ywg/9zkbvN9Av4lI3aZNVxcz8Z+nhi/S7zg+3iD6/u4j4WUu75FNTsXJRYaN6vXZ
kCk/6S3+8KbmNWhMlXO/IeVbjAJ26vmCa1PABv8az3HDV25iUA/jg6lUcdsP77Yj
A7xEhsO9mwJ+a/pWWBBn0FiurIeakVcs+synci//ZXIK4WoS4/w91+mX3I6qeXL9
sCbmRZ3aqNUumDF5P7t/5/+41n+oGbePX0iIHKBDPNCrbW9HMdeFPQgcDb0ORWF0
OCd2SfEE1a14exJA5EIs3Q0JuztiMTnMeNW4hM6Vht1+qVgfA6VeutXY+n9+3prY
Jw7wDo+Ep5zX2ju4Iynul8XqR9sKPMbRSTxs9+/uENSUp0LsSKNVnsEZokb7PxhU
/dY/T3tv3Qyjc7iA+cp/CtmT/X2LINvr0Q/gdgE+KDEAshk71HsfgpbrggD9wNa5
fZrnvTahUpMZBjhH1rfG5zXKf266w40+U2DArHDKgP+Hgcp9Py2ITtLHwrCNAAV1
NY/tqeoelyaQYKym2b1EDMWAMRHGi0YXJm78ySQa4gAi4e9wFVf8ryC4tkeS5sdh
t9QZGbNkEKTVBEGQJ8WGQ3+QV1dpIPQIirjracJnlqc4aBZXNbN+cPTik6WAEe4L
RLTHOfpgVk1JvvYwOaXTzZ9okYOVo2Uvjf9iThQuKLlWoil4QJpxIFs9CU2NxZES
2d99/e8q5HcTHbnR60gHvUhBjtb/Cqs4i7czlGyAkYuuK7aLsNKjHj92zO3MeITz
b8Uzhejj/+KMSFm1Ae/7p8xXhZeyAUi8CLK84Va5Bm8o6c0/McxVilJ+Mwnkh1Iy
0bQQ2/F94/sOVFVNW/QqqlbENoeuOrEG03hLYOVrmJyYwdoux8jBtAWp5PfIUd2m
EKUn6r7ngu2cg0K089z+0cRbgS8OisXr1/vxkDbFBjGvhJT09JobBmyvhxGSyRui
oVHHuZ75w95uiZo0C6Sbq6EU+QuGnNyD7C10MSmRtn1Ldlx5pCICvAwifaiN7jFM
50ytQoNaUhMaOQ7HKZx2CwFZSK6pZMSCD3LRJ8lC9jIUnCmgkgFSXPe93QXBMjsJ
Lvcjj2PnfaLGGPoppXImN2Z2+GWuiW30RQZXv0CNiXFNl1GLMBGZjkWMHprKJAB1
KbctJOgx2WnpIsNtBSasDrsZDBbDH2TlhFgFlMJnqwPwAiKMN3S4cGHHHJega3sq
M4VnCt7UkMsBa0S2L2cVJe0OG4yNHqXx/qFVO/aQkOGVwsYGYJknM4bRLhB/s+yt
navlS5QikI8eqlRQ1UO9HjqigJ8ffJ8gGQTOl3rGHxk3bT564A6/L4eQIawjD0dE
ErdQCcdKA3CwgB1Tj+x0zsI0dEZj19bqK5HFAuEozoWQlqEkmQUMkKQoiqKRzKtL
PbcPghRInFKVNvJMK8QDS24P/3zlNc9pRp0zruT1XCOasAF8pKS7LHLuwoP3G5dH
K5RaUUYAU/LltbtG0ATgsoBoEb4muMaXzPWrxxCK0ZjV1D6uXR0HZDn1sJ5OcAgM
ibfh5RHOmXDGbDSBRihrxvK/JZ1aKBROkSrwez7hhpvsNji0ZozDKLLiTLQ0Ffpe
m0D1kQrFBV9VdIlGyiowJSwPzC6Y40of8+wdKCC3qS+d5rfa3j1OgBHSUq5e2EE8
JxpdWNEelnBV4jo5fZlOSx0HL1MiPT1ii4la1S8KZbPuB/WHzF+JYkFE9bh6714m
NFHfJiWX4VVn97bsjYVbxqrKO0GxsGmEbjhob+s2i1Ys6wX7t83TlP0wf7qxTYAG
E928dUatgElOWhP9gf+O8Q==
`protect END_PROTECTED
