`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yd7dUVsGMhLNARBYt+7WzN/P6XnRBB3KkYjDEDmI0zuJwEG5LIkBXYGMj2fEhr9f
invAdZ/oiisy3W/ChLwm8LcxHFQY6RiFHKRV8LMi4u3Cnr4QD6bb5E50ZSwMMmCb
5LDfmwQX/O+k9MN71zyNODUMA7C8FEnrs4+m8exj99vTIrcNmwdfwjB1E2MDZI96
maw2EJWDAmXxNiXkUCb8Jp3HCuLwcSNKnz1xjzLfVzRdYirtAGHlAKO+fM4OnHTD
46dcb5c6q35Zyr7wgx6v9anx/3YkqtzquTUmxs9esXImUmNV0H51Z0jn2QmSdzn4
FujuyXBMkn3a17t0o/x2FmyeoL/Torbm/z99PmVM4Il+dTtgCuxDILzHBZfb0Q15
ljiVjJNiyr6KsJjgiN13AgHRXNAhFl1CWb2g8wi9WbJnS7CJOAdvxZQhssQ6P/JJ
o+fd1acdGGWRlNjeinz5GF9O28T2uEI63zLA0pRTf2J79Td6kGaHprIWZ1siPBAR
`protect END_PROTECTED
