`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T48m1PjHIp0CGCQGrY9C5hoA6OycNhvxxeq+edvC/jAsqOFsHwoCNemzGTFMJKpG
JXlZYnI6OXQBvI//rVrk+/TQzB/uEA94JsxpS3E2U7FcR8lJmulwKC+siML/3QkF
7YXW2hWGxlh/+XHc6sUmMKvwqbiqw6wIfyCYnX8zSqA46An3v6tPPDMAQWSnv+vC
0/dmZMzQxZkC+3n29cdQEXaJiwJDG9c3zhrzW1h5X1FzWa6hNakVPCmUutVpyoKe
8klHOWpnc8me6xXkMGQhJGkjdiCe3dd7OVVjbMrgQiM/0y4A/i7JWhpZVdGyuDsj
mOY6GyyzDvLER2Hbb6IGk+VYEayoWCr6U8tO3Dgm4Xqn6AdEs8K0DyRRm/2OVkRV
WAU0AVXKJsBpq/2yW4oZPTveJwYMenq21lgOQugs6UaomA1l6BrLfwRCJ3fcldbK
`protect END_PROTECTED
