`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Cf+I8Zh4FJgx4tZbTRmVx+4fBetMP4rdS+zfKZvVWknQBtroP2NJV+Gos0+hEJM
zlUc8AaafhXxrgWgWAgN5mlp9bhSLNGAba/stLrIP9GgWBKvauJdG5so6yCoX+aS
ySQukWd6QuTlSXipZJyyAVzq7v5q7uEzs/UV4D74uGZ61ca3NAyvg0NLAZbOK5xb
u4uhC8CziACouPcilmqWwBf6A9hMdit5uh61VUA94VYKfCl9pscfXi02zm0lx14e
JtaFfqXTsb+OBfmVSC/T7z9cXEY+g+NwYNxFrWtjlOsb7cQuWXsL3ALOLX6OVa0W
wYfMgLD2wMW/S87AoiHku2PJkwamP6YnSOAvNjzude3sZwG8kgqHLNunuCa0LCnI
scrJqXMQG/mZQfHjo+hp+AddNd5dp8/bcPaj8ZxbZjbcLGOZT3pVe1T3LKlaaqPo
+jvaLIXC55j9lbbnJa6vLEyQpOgNym9dGTBoB8XM7bGKiPMmiKzHCiZzpsafDHHG
N4tdD3ExWmkygWGLfkQLYJ/LH5mAz3GNju3E4hRxRbgkioz102fkPYiXfM4mehpP
vohfmvo4oYXADbckuS+iTg==
`protect END_PROTECTED
