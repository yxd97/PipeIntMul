`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Op/1IIGBYR4Zp24Tzfv06DGpHKt1l2qrE+3yIYjYukPQLbAGrgPBOgsg1xCpS79Y
9l5qtsdCW0Bo3dNO0ww0yG5aXojb4NPxQWGR8f0trRD4IlahdCpK7phQpNDKZ0H7
eYHZx9ZNlyJRZXCmqvYKJnyfm+4KtKkHIiY/zd8ThckS2whVeTmFYAndhJWlMnVO
OOownfQh5uczSosafDMvWbAdAyViCtg7+Yd13hXj84WMc/zHE33Rv7I7XUjcydbc
Km+UxmciIgDgz3jGH0X8dOagUlhMgtMNaVvGsXkJm2XBEhxu3nezlgOMdZjxCcIs
XaxI8dmfJy47H0LUcL3s5nX+ubJkx/MO4ZgtedEq15y1wXc98SEdQ7M2HiZlPrdM
MUGR/UhIdOlSezFsxZ+LKMgcUlDWn0oYlP0e37a1CyU=
`protect END_PROTECTED
