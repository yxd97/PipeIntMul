`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EaPjqQRiQ93BkMoG3NQVP7BreEKGs1e358s4fr0im8Oa4vjgILwDrpayC7ztkiBm
obakHUDa+P4v7Ppvr1wtS30HXAs3UtDSqKQMsQfphith+vUbkum85UDMb8LGR49U
QoyiQR82DmAjXjf3kj/fCH1OvXEfFmoLurRnN0ku2OnAro5Ol+e+35eHI8ZlisZr
59rDSlR+9SL1qBMp1WZ7PevoyFzl9CFqXd9wPhEdS4HLmpiu8IoLmQtb9Ke0ON49
voccZjKz+C8eiLGDWZlDDRCrFfNCzX3CdalL6+jlLqgKqgAmYeRojCRgztju9caC
2R0px+AKTmjald/lHNjhWnZ5kt1oacUeOpmw5ekwRYR0BqBh8P5v14CjqFKyySmW
xxRyodNZoKraoqMSFAU/7FhYaX6vGNzswTKLtj8cPILKtc6N0AhLugZEtDVI3iLl
dv0ioEZG3b559IAW9LuwBZ+n2cwW1e7QyuIZU9DjZ3iT1XyTAU5paArSaEoLltR8
e7ihhN9Pqya45nrcjZkWWndhTt6LDb49qgpRb7euwEM7AhB6pr84vQOswnLG7DQo
4e1Lx5YV5or2kBS+eCUPXAAd9KZNrksjWoeLWw2aheECucjdeO55BPo0niHr6TJ7
IdsBKBO7jfIt+E5SglR8CzuDDdsS7Z5YvZ9S0HeIjk8A+OMeoLPHgaE3268x6X8k
Z6d5fCqvAAHk/PMLHgSNoHVUQxMRKxL0s0hoDQbpWHlGkNtYaLMsLiiGvWDOPmwI
IPv46amxLd1a7KIf714DafSvMd3QCu25dtm0vs6qX770kPJDNtcwpmmTslBmV7WA
qw27tkfANI01udVRjLZvAhxvw4RN945n0b/DfMwnEAwRx3nMu/FKqMuUsZn9UNm+
tBHEW+eD31sltYre9hHx4EMuYHg4xcs3fI5yMgdkDDnAklNlGF1OQ5BVfG4YDPwf
UDoZX5Ka4jJg30Mo45choy1MuTGl2j2IVpOIFQQQJEPWEu0IDwEIbUNKvWaV/lJ+
raKHDwMus4/wutEOX/D+P55CPU78n3ARiBW4ADnj9CVydVKMr7snwM7q0X2MHUJT
9P5AXaANnxoGCYQG7BEi57alDo/ii8v+yaN07JUrUUUPdaM8i648+UfKCUssrNRL
`protect END_PROTECTED
