`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a65A/UIGes62jl0Fin2m44NOmUiatD8DD/SNPehDB//A8HcyLA8axTfxocnS43HN
xpHL24LCPngRfd6xSdNvqAYbKXZEGwF0IEwIe7OLD6CPeM33+Qz6ACMfzSHVnwZk
a6XpRyCSTH6ev+glNXe9dNHtGxJcF6moPufk0CcewJaBItx1U62y2nPh+RerSIYs
zIDNPgetJGolAfwAee/M1pswsZFK6Vm5A/O+ylEpM0LHZoJ4VyuLm7NhNm/IMYSc
fBAuaQJ+phfPCN8RlHg8h0i+mKozO/oEi+ABmJLbj5snP9MJTyP2KSw//5j+DW57
OiTIQ/SuR+yDpyHc6y0zxF71RUsFI6dE94FRs//xw70BExd4LV38PkHYE0T93Sxz
wkHqBxIykYn34Gj0FEPCVxAvYjJiNbDmpipVD3lecsLYdYphfahl6y/vk96/l/16
Qj8te6maaF355gzg9+27IrQuWkCqNcC8UNvGOretzVmmbv7qQpi37fplbRlMMXWv
5SDraA6LmsMDsPhGPPZRNenMyycz6nrJWC7zMvysFCqwqwpyPsOxws7S8XC+Ld4L
zxDclXnKLPqLT4KGmx6DrwXsY7P6lxO4F9MephoXiUogTeG0YGmvAgI7EIiaOQ8z
G2vCSOFlTuHMjgEASbaNhqyw20JESRGIW7yIPzzsas1cQoUgD41O+Cz+yYT+bYi9
KmhoYHqEU573Z1LvabzoboONrAnldKrHB0vl2sLxe3qiGcS5M4YAugqGH5AdxboK
yblJ4WigUMnRyDMmsCj07lf07YuLyzMMXdmI4rlXfhMTd84jaHAEEO41HeHGLNev
9dkwzwIK2ZllVztqzR8LVyPRYbPzU/hMVmpyVLNygzVELn8gkcMyqu9+02Dxm7qo
PJahaOVLgp4glZKYN5fk/4GtWGj6WmnXDvJ9j6yIS8jBiJ4c+BB2mbK4nVZIRrUU
nbS85NVOqKCdLvLqTA1ueLK0OkV66MUYyrw7at5gyjtNSItEpfDOW0zTMM0jVfOt
Jn4rKzewbj7i5sP7kHyvTLToA/5qI1X74NGvx2Qq/5Wj7WC9JGiY0TGlDmA4txsM
LkeZi1WoJZip29/VSQLxw8uVR6zm2YgaQNx4MP+p3Bc=
`protect END_PROTECTED
