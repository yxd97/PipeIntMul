`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ybboRY5J4gGmPvmUM129SgTRkHBybdlT2AF16qf1ICsCJWg1LHW8TfQVaYpjUZgz
uXEJ6LZHCQxO41xmfsrwcppr04ykDLsAisiF0i1i1z0s5MDAOq6/Qugi0SKeXe28
dUGpsz5N5tJUXoYuI6ue2rGp8UtzkTngFM1K4iXqYKJVcvZLohj5o95QdJJ1ElDr
Krf+swjcn26aDykw/7WizxTdM+aOKQ2BUJGL8QO4Uf2iil/5BhaeDBfBHcZj4fUS
wVQbSgxlTaCBfgr4x9RQyx6l4Q2Nd46vvh0X3HwJjCBCGlVjulx+emL18uX791FX
M65qJNC6fKqdLZDqSrSqgvxu16/AR35Ep6EU2J2dmZJ1+W/ddsVGjWmcNYL4M5vS
abOkLpee5fOCNLUNrP3n7QftLCRS4VLuiDnb0Nt4GI2u6U1m5tWB0wym3knkLkgr
4I9IjkoAB2fDkhnoFqzwiYBB3xc6kYZUJ3xkV2hK0OIuiDVoN/gPqE14LrbngqGZ
UXLOq10nkOQR+5cKkHu2VzkGmlMgxXRSra90SVf7BXNPUYApwbXXIey5PIXCMuqV
jrr21kz8XcH+Vz92n3aFng==
`protect END_PROTECTED
