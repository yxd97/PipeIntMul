`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vKm07oTPDl8Qbb9WFodAG6PHjREyxeQ9gPp8laVGO/3780+LN9nwUJ0Sy+SRue8r
mgKJm9e8JkmEREjP8/aM9ztwezQ6sx5FD3B095t4Ji3Run9os83bgO28G4/ADgfJ
jNp7t4WC06TCb9o8gtPwLBLxRUMsPoZMorTbdip7RYbl/s0nr28CxHnCL31RHFRJ
UOxM9BXvsL4FTtFaLN5eE44q1dXA7ZcEWgFIzGxj2bLwK89djws31LkshiWHhjP3
0oW+KRMx7So4+PPqz73hquDOtMXF4ZUG+tHb1MY/CCiMJe4CUMNnjaZNhJ/xu4mG
FKbhkE9tvD3Dbb0o+RY7aoWNjeSfWgqN2Dze5wVDDS9rQe7+S7q+3saI+kiwkJCC
tmefMe3m3nepAny6hfLl56lREWJayuONBdu+7/eToHuuBtFXx9GA8TUmjYddrLkT
iCowtuqByf2AKG3CtoDOjEffNrNhapBAXhAGRXZgGhZeAHeIL3vvWZQ+dxjPZz4H
RSFHwMLd8fkSK9E9eiwTR5d94vpQcDH/OJ1k0nGLzdAek2zvElkzE7Ihxcg2iRDq
bMbTpRlpK/XMGfAU4hBNl4PIklxxGoKQBZNERteO0Dk7CZG5HKk0rA9kdNem+xhX
F5XUy1dl0HIMtNRIQ+0INHN6kPyT6Ve/b7H3yRmbs0/UeheqHNrVPeUJyNsHSg3H
CG+t49h74mA7AGtptRFTJj7eKLi2zfHQbGzSrijWhv83oIZi8oeJ+YsOoXbyxlu9
kOTN3PD8tldTl3SaOxYwOnsTW5Yk2p626LhDBc3s5YwHgUkDxt2vqM9EkMuT0mVw
tWC3VL+FJIFrUFktd4mb+C+D3fGGY1PFbNXS9BohYDFlReW5Ss5ra90vufWnv2fh
RDqUiYJ1WKGr0CGzywr/2YieoWRbWhhzeV7KekOakYFpcbnNAO+CTNHQqVc0C2rM
UWgjntf0CN47ZSaOOJ/ub63RAa41jMjF7nDlVgUpiV910pjwaq0TwcWyeIGhkb76
IW01QMSbccch9xVD/2bG3e4U15SALO7v0CP3Mfy8qiX9pmuzE6+A40J50Zm2U3WK
fn4mfhDhNpjOqBK1RlX2s9jqjHOMo7EzTsUV/QMW5VR3WjyxKqnxDo7cSfOyxQ37
xy1zpvzQemoiGkxRDSN40GepLh4/+8WRDx5Z215xqyOFqhFMLKNeshMisW/DGM3l
zR5oVmU9JB7nZNDahkAW1wNbQxrDnJ3A1DBWxihckFnnq82JGnJHhOK/XZzzHQR3
n6b13AkeVAr4Sp4pkMdCFVlp6r8t2IZKz2FzvHp2Lq8ZfR6EBVOzoesyfa6AvPZS
LOsFEZLArREa/PcU04V+hAPbcefp/HU3Hs+Ixqi2VY0gSSk3SEulwLOKuJGA7m4U
WzIF3KxgQdnKwd8s6HV0xTR45V3F26M2XCseeNDM+AD82oYXh2tCwicn0kguNwHx
Vcmx2EFyNZXUPrynPHWA1r8SrT8kuJ0RzwNJ3FwHdynf8HkVjM1lrBdr2kbsfPYs
hehGmRvwp2BoHM/mj/R8Bge1jHr4jZW0TQDf8tkhsDdOW6A/o/P3qBfP9UYuYzV/
DaytaKnT5Fnqo2/w5kit+kjzcR6Y4Ilg2yzJoUm48uaIfpq7xZNHo436EkXvRCHe
ZrNDw4yUaLN4xqhNbLJ9Q5wNrisLML83gLY7GLYEChO0Z67fpfkalxMD5lmveTAu
0zzASvaOvCBIUmO8bff2/xfJCxVE1eQ6rE3AhpHmnmvNG50Ed2hecI06mCF6TaBo
AsLiJ/b3LWHBRAiIe38oSjtAaYelpHJSQmuNhaxaAjASVkyHL7NA9onmkh0zSMOi
8iVbYA31P5BMBbxLC+4uCIMTwNQPjLEX3E4CfD4hr8EzS7rVIUawTEA1K+Lwi1Jt
60NhJYaJ9uUCPz+UAIrxiGTUZdlT768lx7b1zssknylcfWSYV4ntifoYnbteU4Qn
AQfeImGt5fyTA5c2I6Vi4wIQnuIkns9dUeUNB52T94lo2IG9LzvBL6LIFNRoG6Y/
yJdlc/bimNmtSFPTgiCmn7v2Ce5g/jvfxolj2FYX8l7/5Sd05gQ9ApegBmnxl/OR
MailwwHrdAh7xNRxlu+k2L3TcG+f6HPX+mz2hI552Hg/jXrU8xZNNUCcHkrS3Hjb
yNGZ6mP+8ZgvS/vjeBIdlNBuh+n9gywxDlXew8eoIZW9+aZsbNdnw+utW2hS/oDS
CWI8+Uv4D2mMxWjxhIW9m1M8GytesoKf4pyv83d3xDoWHdyu8ABYg4W+vnLT6VIe
Jp3Y/qjjnsXn3T73FkrCzIrbAiiCK5QjFU3sCEB7TabMUDTdULHh6gIaU+7ogFlc
492sJ5/WWvoDziFRo/CRKevc+wphCVeXQiCRNPZs+hzJcPqLoOzW+4JYKOQhdt4O
BKlhwTUayLT7gu+28f9b5lfARRwBveHC5L4p8x5Xzy6ut1hrPtZSWWXQvowIkEYe
MmuH8AA2IREYCW8booS9YAjE92vyJfoMLXas/nLinEZgCMdWp1KHVakukCt1bNFt
GM5HFQzL/IORvZ7R4PIeHJ77PGZO73/9l+kkaDV/q8J16A9hBZbiU5H9ewA2klTK
0VbHrTmRwfG9qMTbh9x8X29gLGYEX4nvRhrJGOAbvY45I1l2zwJxQg2w4qXEOSZP
68w0q9d3VYCHUS8Qs7Q3Obzp0XkHoZjZXWRc2qOG+x07+y7PO9fvvuImxWPYlEWG
xfW5OuLKRCC9U8jD9i8XTDqhP4kIJbpDSLieckKzBYCoH/31GFQ/I4OYINkOqBfw
YbqS+Fb3jy0/8xrjiv1w9PYYiZ4vDD0ZRxO1Z8ZBPXs/2IDHvlxEJ2bbudrGixkV
TyzaM5X0ufeyh9YMrR/ZZk/gseQWr7ljKvIqxuYko/ihS4V67g/PVZJK8ngVSBAR
M4HY7ooLJFOpF6A/scDqg1qGO6yHEymhIkBaWJDQVrwFrfztkukcY7I7ZxPrmh86
V4boctTIf4Tn/tceBMu+nURbWXOBt2XIkbo3qbMy69MOav6avmWJ+RQ7lDlrqgDH
sWaHCm7PR9xpuFomTe9LQvvb6+ibuZDkFypaVLnXpteuYIgYpdoXOUxjIzAOG4lj
gvM48JBLvrU4UHBOZ6LlTPf5ExO2ZIZoGi09xeCTD3F0QmU5IHDo5zoZuVfPxw8P
Ko0d1gbzyxm+6TEGiHSDc/JYsWa+1k6EZePVggAoiE2Hrewh9WxmjW8q+8STWgRh
tcp7DFLLilTM/EVUncqPMaUJzrR4tUyvMNM9iVDCrMd09Y8Cl/f1Q3in/UiWaOGk
GPwiIpmZqmXsEorGj8+SmnZIPHyfxM2+9Wq+/PSR8Cg=
`protect END_PROTECTED
