`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdQBol0mDEtXp/m6BbfJtVCOHbKuX42T7oXrDJyOBRh5NVHvfCyASQIIPW+4/WsU
k1wNkD6I3qU2Ep+iHwesHfevizsoiJxzuM7NRrXpnq9kKpUulGtj8T/ro3WP6ZI6
Gcx3gb13NHKPJJ5C+tLNc87/BxTJEKml9CZAAmWqWYKtL0BEsGLidNWAKTiIks/d
v4fPP0JNJRCsvdPvWXB0QH9S4fH9y0fbwGEs9bKolqqSdyL+Z8KKUPb9ByYMFaUm
uuHC8WaPBmf3FNxuZ6uweTQOTCJr1gml+3RfoGWxe93PYNIQZBKAvHMOboj/slxe
gVbhbrNdYv7ubwQaqHbMD52Ng7P8odSo/aiRCC+qevmnAjFaO1le+o6I+pkuePzn
QXzuz8xt11E1XEiuzdfuFY1gE/fy6c/961daMy3uGxHvQsOvitPCY/AC51IA1JYl
rnrYiaDIVZRPfatI/oJm8ZHKaM2qfYBIqnNkbaGGf/TSDQRPga9On6navndWP+HV
+nKyH6QSpnC0stJAi82+pcbaDHZ+cuqd0bPGNRH6rspUXoPiG5jfkI+odoMAnS0z
ng9xvFPcHDYQCnxm5/bBCIfXJB/FZn8ye048HPlvzRWwLFAwQY03BLVJjFqbAoEI
XFyIT2UfRoQvbiUUx4f6b++FUvHgwPcKKLQW5+SXqXo=
`protect END_PROTECTED
