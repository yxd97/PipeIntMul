`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Px2sdqPEXTNhllfJqCDoRtvZZvz+qWyRZiWnr/gmKIM3cC/U1hqNL5o0hUUDsP0H
bKdaVSS3AO9oHLaJONmyzqFUEhkVa6MI2xqPQotGeVDcoAjWpw8IyHzC2RSON4n5
mZibJ+UFJ5wVBPiXyEnbTpv522hiezH0RgaHykzFbsYnDQrWAzA64o4QZk/LI1Sv
J0sLbGSNlirFpfiZIQcE3cetfcOJQBhmOzsHqAumgDNs9+VdIHGx6DGusoh/WkcZ
niucOfjtrGrF4PbNE5ubK/mkEPTWbK2muBgY0TLzwbOAIFW4YpRHlG/OrhaslMdF
x4BpyhSViyLso/YzGROELxJ5wPZvGxu8nx+furOC8JH0xJRJ+SvgoaGQdCe3tklE
LR+vBySrViD7elAESbX19sNw6wEiYbgq6835YZftTpZy19HCNPhhRfpMCRzcIoze
G9nkBSl35pHM4TJ7cXx+tgyuGg6Al0kBkNNwnTS8o6CWseydzyQuDsA0mFaqWBhh
Fu5g/jQYuiid1JAPjpx7V/SE4yujveH5NVF7QEOA6wyneZhnFu4TVPAHOv3iD/VV
87P04pw5nlVHqbOsHqd7Kp2qexrT7Buy34UXSJ6vBBlcr50gqCbqLWGDYcvedued
ZzKTcjS2o4cVnx//vAnREjKwJF5WdmaySv2aaCRcia4JSdE2VI4J0AtAmUig8LtJ
c/Hv4301WHkK59AXCQZuE6RQpscumjUkMmO4PRlndmemI5POWn1LvdZRSXfEcmqY
ljDM+OLaXJfC5YSbu26QnvKzgQ3QSPolPigufNCI1EGgZF2lANEKybOL9/z76wNs
tKM+GLpnsgjB/SM1pfzK2zOSE6gyuQsQ8Q3UXSnpAmFSZjr/vl9N6Pb9Ok5Gvjqp
`protect END_PROTECTED
