`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
80Xss134WKaeWwKJ7eHGdHs9OVc95ba7WO3VmPoPgRgsH9LGMpASG3CP2HA+ErLJ
YCVfZf5Vi+Feydvtgu+653X1d8OxXOEZRcYSxWlMac/MILwXShjDxRrFAekIs0gs
TLsPbLohzRNByQ8C3Vimcn1XS1wvC4rlvxNbvl5NJYtg0EM2+dGYRiWdbAHBzJ4H
E5xIn9V7dRoy46pOvveOEH60KY3c9lyZD5J5Tnq7/HCd0kyFle4AYp7aUKIFbGA2
`protect END_PROTECTED
