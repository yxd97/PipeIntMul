`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/H/nuXVOCSI0s3D+GPAcD9AGVHtdAa0cBPhtkGtyDtLvGJCBn8nbq7gSWyf2WkP8
IlhTomNs80xhNG5D9QgX5yJufYEIWoAhkZr5Gc16KCHt/oqtinEbVRH3u0Cgqf+B
Xq9BdzQz1zBH+ZiHcm+5nvVufacmm3NaP00g9+M+5TFu6SJhkpef5Rn+xVCpCtTd
5goHFicFYNBHNooTJ3DlEK99p9kH4zJxStw8vL51QWC8FlgtpUlHcTE1/OJbKPW4
bw08A/SVRsEyEWMoJuB/3Cp0Dl85flJtD6MH+8Li9fSXfLIzEQW+PH+b81JYZql0
ewjSfcy9EAfIrrDgVt6DGm98fw+N/M+9kJQ6yU1V7dgKTaIB1NxV/RiTZs5WpWH+
6bvgefzf53LM5o8at+rgIjX27spg4V0d32hWWp4R3lLF9kX6Ds16puEG/BQU+MZx
13yLY3Vaqxu91m19QreRYkirioL84aAsGJ+7mH4PekyD+TGvhDhpo/Sv1s7d/pXR
DEfrxzzMnhP7Gr9Oz/J8kqKv1FbY4lwkbmhPxemw7p6c3aCEZSsg4PJV1I/FvwGG
8U0GitXm0/CvBtyXuvTri369gLmKnf5UdHU/wycFT9eIPban6UgVTrPBa8neJF+I
yP8+skYZX2XpitpuI+gOHoZtoRwQl7Fw1d7b9BmG0VGjM/MvySgX/rg6v9kKcX0S
EqooLbQbLa/4t2YMVJqVfAhwjFjgOzlXYA3+VpQOxInI7NS2P4MLsh9GLzNCFBT7
6yzcafsPReNTPibEidSCdVLHhzF9GrECNIWdmlW/9Z7v6WT+zYckVs9MPEnO5pNj
4qM/pMzDEofiglfnOdKd9LC9fPKmZIBHwvLUOKkBtk+NCBPoYX1qc3jEMGXukf+m
SCTlETADkXrptrBZPYXriDOruGG7sfHN67Y3DikQf24NFCOju29RVw7iB1ikjO9h
FyyzTU71+rD1NuHAIEtrmFf8xsdkHweYvcluYBKA+/mtrp/XZhrf0NpApGvr2rEY
+axsQRpegqifle758dDss1BMUUG6HlbWJORhrwQosMgbWU1PynzaKADA2kadJRbF
Pv1BAsj6/z+JPVKJfyYdt6IAm/kzgEJbbLNEvvu5v7GgGSsvqGIypyetPZT8OM3c
Rnl4iXJdYP0H0Rv7xKey6iQ7j9uboVXgn5SO94bw861+0wMyoUyBDeldjHYXBKSo
DgYFtpdIjgpwjtriIn+F5KIEt9QYX5mw8zPKKSW66KPl++p4Y69EduG2qoSTxR8I
ghBmBOnbpQfIu3Z9d7DUrdWriUbt1WFBU6/j2tFqDwCcedpDoFnac9iRL51K//OQ
tUgB2IJJJajCZJBbv8mKo4EzdnT8Db3MKEgH/XDrH2VyYioSKX3LheotvS7XukM6
YaYxEvtIYmuwK3oNDTL5mheNB2vuTbOlyVLhCLOS2hw=
`protect END_PROTECTED
