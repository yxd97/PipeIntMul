`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgioY+ENV7ewT2i9/R3Oef1R2ayUWHU1QOOyvs27kc3pu0/u2+4yADohscc3QrRt
YFgEWkpSqAXinaQ6H+xXqYIHTzkuO4AprbnN2ZAb9onfMwbNkHidUJHw9XmyeKmM
7LA1PUhw2p0Dh8C6c9MQCVIzj/5Es/ZdmLPSxPVyTaAwwoRUDb0dgkBwSzOjqG/V
I5dVrAFD4cuqgSKOrgNef0swn5KeKMessxMtp31AKnsCZ4a8bwiXZf9E2KRf2EXE
XAbrl30+XPCZQYS1nYZvkHwEUq5wqnv43FV0O9Qp5QDVthDGti9BQiDUcuuS3vaF
WKuvnqQ/dKcX0fPcrrQMFsUkaUZypQFMIvwByetE7XyiRd7upQapHxMy9j4Q/6Mh
raYQzogGWpGFBQC990kG+aC0pUaY+ytCgtt+Drkcj3no4Q8nUVcNfG6isA39rFGq
T0hl6t6Fv5D/TW5+SXjnc7Qzd56gCJ6X95D9EH+jwD6LL0Vjz9FuGa6+hMmyf+dQ
ahV+H9uZ1zDezpp6IGtoypQVVfTal4ab3hMoRKkZN4ak0Q1khf739csuVTWWloik
98Cg900/lhb6ZzqLVj/ck3XrEZ3tgbA0Yj6DrMdIrMIE+fBIsJfCqqcy9wsGKyoD
h4q3G1U21b5U0kDOnGEEM3Wie+QGrTs1NLDlaB5tqBBGchnwQhcnMCFuUqEFvDEE
M0v2jyLG6k8h1VdBEfralnQu9WhtkATiyC75lxygtpqAlpY8PzENo5XOxP6N5GNT
ZaRfIgLZsCe1fRcW+JV/BG0gmAlK00iJ+JJCL8NVsAQUMssBhHXLZhoEXafVj6wt
xqYFCgkPOb8JoSfo3vMPF7WXO3LY4rOTEMMOrONhcUciklsWx9ICQI2H9xdhFS5N
lMYJTDzDCiJ35OJBX8W5mbtv0MmmKcu/ZekpgTfZvRKEZ1Qu9ZwWMRCRERgaaA8z
1FeeUfCt4eg6fKNITwLigaFhwn/m8Td4T5V8gBctbRM=
`protect END_PROTECTED
