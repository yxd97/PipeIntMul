`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sep503cS/rpbjMcUQJCXuPV6+IbvKANoTBgftLJyDE3mvr1V4GuNJdA2Y+X63YPW
UIB1em4YaeWe+zMR/cRPUmU8Hunlsa2s6/ysyx5c+BSH2KL7+agYBE9Ai9Jqz7si
iGxO1hNSl5qzPkGDGUn/l0AvotqWrZPzGam6ABl1DzkSGc48ocaw+xIIDEPVrCEw
MH21jnLzj1g38Wxxs3gD/mQfjv1sE5xC4uVNpp8WBjEGNPaaER6Z4AKpOMBsvS1s
VxaKZujOH/3nrbQ42xvFqPEgdatMqnHELLbQiA1N/kTUiCT6HO0vMiWCeek+CXRF
yIKR/H8PZgvpYC05oooUwBGhrx/U3AL0PM+E34fQi8zqjCljDg952/plnwKJOfaF
5zH+ZzdFSAG8EFwJrOlCwI4mdxB93kKHYtsOALwe0fw04n2Goc/KBPuXWmAbfRoj
ZHiYDuRYt1JV7juu8CpiazgSYKc5Phj90Ew9KkjKB13/vO0tR+4iXEAtt8sMD/ST
vk0FApT++vec0qVij/mnhcChNbnrYIw1s32vfZIuh5dJEGb/3sphk+LGtCkwPsWX
L+HD9wwc43sNxWNu2it6FH400v7ym05gDaob34FHEK9s8FVAMueheZu7Qm73kicd
oxTQaX9Zky6i/ixWvKdUVg==
`protect END_PROTECTED
