`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XpbA28vZ0dUdO040TMoiZ8t8IBOiYZHf4kI1SDrDa+lbv04eVsGJFskG4SLpAL0F
fVZ+smeB8gkoM4Lh8e5KsmoqWbYLNIzkZZAoLdPwjGQnxgazRdeevNlm6CG/MQKv
DbXA5ug4IED+YBEfSkxEJj7iPXFn7vJ3HOKyBjE1bOPtvmE/43WTbthpjnXuzZ4+
uSe9UkymrR4um7mQRQMOLG7VaY2690rW8cm65cVA7cBxW51LnBxTOwBn9rsHi3r9
zM8J984rdOdNnpHkF3i1XlF7Ae5DU4efYTy7GXGW3tD2PPU2c3Iam3TUWWqA1SYv
J95r4uHTm4X8KjknHkxjLAG0ZSdWQNAwQ19+CxktLS76psEy7GE5wa825dSqDePd
9HGO7gndONG+2hvMBG/7ZCnMtz6fO+Ezi/8ksxE9stG1b9BNYfJG9z2bJ169uo03
iYNxRl/fNBfipnH67cA3zKSy8TMJDKtepy9IK8xKcbmn0Ek54p/uaEqPvfYKaTGU
VY8kIbebwZA0uZFq/hcrzdIpvVbn91ua4dh2vfCzRulTBc3TRaBAZZxnUd3HVdnO
t3HATqnHCRJjZZ2dC3KdLuhQWc80cevZZGhycqqIkIzTTd0rACTutm1pu5F2vhmr
oyiVCf+vPCaT12mleYV6erPiqPt8kZG6aYDyTVAywMT4om4LWHZB5wEZPdk4qM11
jatciR0fjL7A/onqpMPgsUkg2mhpPW/dpHqiPIw5UrZa1lBw6FQAVmEFAI7VD6XD
NLBTpSQEq8T3KPkuv98IuTiBrGMnopDdp8hW/82KTxSlE1JVsmJcdpXGX/RNdMgO
8A2KPenKsxfgExIDikhxDlu3s5y2xpqW68F269+QNj7kTQwTfQi73BLfnz8jvNxQ
u1QmjhgbyeniM3yUrfFHfr2tg08oSVqWE3KfXEfQxuev85o0Gr5o3VL+KxBuevX0
7HvwnNE32CkK+sOUJBALhWNE3fvcrk58tcDS4yORTLO4zkwb/rdcbiz18ypWqg9o
v8/YdVfdU5fDWrYOZi/vFTJcw2NxEDzo1L+NjslvCm/L8PUZzfJzLmGLmrHDxA1W
hnH/RloLfu/J/Ga0R8zsNiZifiy4IZnbINymo9SOBNTkYGsG54UOgTXOaikLsvqK
PDEYtFGxvE4QG0a4c0WkP9hpX1WaVhn3RuudElKVqarthWYgLzLbO7L8T5d8xuFL
8m0ZbBUJ6m6Y9oY4xGpcN4pj7URYIhdGT7aAvbEgzSMF3gN0yj9QLZNa3Jy4dbB6
IZYjZIpF1fHFEdKh59C8X3vAEX84UXsMv4IM3MhInI1RtHWNna8XT2ChJKHnMTpY
oETKTHsQw1aNsbmQz29QPTYxzrCk/nm1R9p2IDjuR4lABPbnLTwOoJC37fhrmsxY
pvHfjA8v7sACBVgrjC2A5j51dKBwGOeBQYSa8jJZdKKWj28gVmxeUUVuRhnoVdJZ
vohLLsXv+0BOtFpsKj6mh6/9r7Dy4vHPV5n7kRHxJrQPAHOqF/h+49Ih0jtVBL+r
MwAQSzB1fiVxtz36GtJvXhK0vIS27mU/QTkZcuM7A6r5Y1gTaVb0l18Lx6vL3fRD
IhSbKWMTjIw3oYP6TDVYKTF1iALTnnbE5FV9uf1LhwhqjS3nw0JcyD9Iz+0/OV1n
BrPhiJGRylY3SDe3gvvLH6j6oP7/XxCMyAAlG9v+g0Ce28ddlxc/ptCL1guuF4Jf
dZsj0jCkZqUf7TsAcmm0eBt6l/xw/oO+hVzOtkCP5F8lrj9YFBu+1kbudsxtw2KE
km/Z1OFEJSrguCK0qB16kvS1pbkWV3bervLkNRWo/8sAs8zZRkq+lXti3Egt8Tw2
Qk3Plyw+0EjHWs10LBtkEZOVoHdkvhEy+gkLvfqTXD3cc/Qy/I5qaQkDeg82u+9z
9Zg9BkWslxx0FcSZqAq2zvIJuJDQzNJN7AgA25uK0uD0NiH6bUlmUnyCee42CN8Y
GPYzINeNWH2e+DpiXiLUQVCtCPhUwALmjnV2w5MC1WrRcr3Pzjqb4h6l+LdA+idy
5m/FvRFRUfufjDdlzDWZZmEV5MQxElTc5wRDwvMtSH9A5oP4twfvgjJDi+6bgAax
s7qtsWpd4jg+x6RMWGzhl427gmG1RsRNCvELIxwVNBdkGUL45uK02gDYNgbC45Rq
0xsNuX0WxN87qdmvsJ4aXho+tttDOmBpv9LTyXCKY9TnHgDNkNIy5sFGFCa9qupA
kPXYxRzlaEPJ6mgI79xQ6zaKvZW4epesEMtL4jXJzwfvxdFaVgW4sKCiuG1x8W/u
skk1X3SbUZ3BDQ8s7At7RexsTz8bv//qM6JRPAAdUDVdDjRDEZXT1uLhauL6p1s/
/X4EIYKlONTZhqzWZ4AWcqpw8226Fjbaboy9m528X6sfI8BdDX+ejl58mzr5sJcu
77zhdhl8EZSWEtepUCcy7MOtYDnrO/JCXvzNDjFMYUIuCbsovkxr1MMNb7B/1ZZG
KSNF1AUs5KNfa4ZxmHK2TuMzYel1kf3xJOGF9r9DxOJYQSI/JrrOUgaF7AQ0sV0C
adfuoTyGvNtc+1+FPH75zEOaeBhpjFRS2hiuA88rZKdEE+ppP19PISq9boRnFAa/
mscIhYTbMnWwGYn3wjPj5wJ+M2ilaeq8mDjmyfJvlareU9gZRnyQjAcpEHnwBHWr
cywUeyY1We/sbewwlkZZ/zWfuNPKeLutYFuJuqw9AEYCi8JS6af3R0QQ8GVmPOkT
O8N3zQfj+g3Xjqc/bdAK5xjDOOycOIixnqBpsoAedV1M/h57kYpRHgU8NrjRQ7w2
KiGXhpYWrphDlDaXjVllKmrL2FaRM5GUXoIHFr4uwShac6tpt6tvhjUyru/0jZPx
/RfjuhNvu3hcf0ducA6LW0LPpSPrE4yCqBIHxvK3w9Mf99v0akPVHeEktwS3cOPi
tLvcoXn9TVIjSKGWNkEEne7x/n0cai/54JpuWY14g5wNdNH+HrRgWIOo+C1AJYvP
cj7K48vBvKPHTR4B284dx6bE4euX49veevP9ecmNa7u3OOYQJKYuWZcN6GVDfizm
MVGYqnqYcRUjzW15r2FP3hQr3HICyrRj+T6xMhApNJ4400tZkRCkd/D5Dsn+o+Ik
HmQIAXRz4s7GHvkV+kB72IXZmQAJHO5zw5lmjXSWH+WgZC2T2N4UzDxQj5bM0DuT
uHSp+brD/sNYGBgaN9Y8zxfPh+L4vpNsRoYkTHVtfjc82gswE2GUl7PeCNvm37wE
ixxRcKQxDdA8GY7EwP5raCOdrgkNpIR/vbfjXhQVdt2Txch87rRV0Qv1K8R8r/An
hueLoHzcqqr6XVLgli7JZ590USEcbJ7dBJWWFjI/fV5VOajCoZNjXlcFGigq7X/P
wqOmSRAsfL/LN/CdnF5ZJ3ucN3viIDEL1vtzm7bJIDrRHF0Gj/BwvqtPEUxXrFMe
vRJMnSAJWSCuIh1tNv5zp6DVVk6BB/wksnb28q3lcY9ztBX1VuMjX3NfD5d47ctK
zGC77ZTAJ/6KEXf01NhUdWjRXgvmxNhJawnp77VvuB0ui3upOTCg6SrRZe+V8yKn
LMzIZxyd3dcTKCcVoogs9nyOKV0eAovUP1uEzvhFjjBcJpSPSv+L8H5YU7lpmfQy
OX4f/CUjhFScvJB870iPm8PCtMPxIWbAVt/vQp5ysQRoCoijzlDFw+VrcYNaoEs+
75baCMJ64L6/tY5YJ8znftK0GWjopyO+AER8G38fGJquxoiwcwcjr3c0g3gchhNJ
b7jRbiG3hEyiFpmkaAmyIB93RRdBhi0hWFu9S6+zoV1PBxkUxVNmBvT+d3HfVr7j
AJErvhlYMoWf3rMwxnKj07/hi1EVNCYwbr/2/6ng4Rp2I4+qqQBF6xNnLtaXz6UQ
htX4YK+OswU7JiHCVoh4q7zvJB5sGF8wQY5vxnihLGk6Oo67TdIcHfrCANc4w4MJ
OwWOHZfOtW6PsIByqmw/T5h4Uxe01b1RokRAhMvIO9sTCYcrTxRHDOZUAXoj8tCP
mvKY+H5oiitjxlyGFpME96hM5720VIafelkV0l7PTzevMk2Y99KuuPdFpe0TNbFg
66d5GVK13o2nd5c2MGqYlvnwc7Ne5XKSY8bZqOp3qJSTGTuM4KQecJyv3R4dJ2qo
zyVmXegIpMGRstJp6KIwr3fznOOFTs6tOExT18X8i/m9eZgGsztWfgAinNwtjwaL
DaDBYCjtZHchkGrWFVF6m85EeERzIWuertTSlmx20s/ZTJGy1Td52duqMaw5f5Gp
6oyGCIxg3TSglmU6PP6IILuJ32VnHIBnw5Jk7sKZEz8tLG/ARJVRHHehB/SBy1CR
l30dC+Xta36MQ2z6DaOmSkkEq3vgfvT93sjbKX9I0tDQlxUUW1SdbnhcyJROHUFf
jPd8y1CaFb5XxZs15d77u7jcG1G8gtL4ep4NyTW1uaC/WE5hWzHjkuTuRaVDMhVV
phpESy74YmlnZH98bdS6SyCCl1xkwwoyp4RxIqLWSyYbqK1/DfEHXrbGA6pKPj3a
fnbRxK7R/ituGvDP+3knQg==
`protect END_PROTECTED
