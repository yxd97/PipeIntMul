`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uUbQGFBZMfVOq+aixzdevRKxcXsJLWIjHwUw0Uy9iA4j8xCsSOCzGjDuute6oyr5
UBPnI6kLiCYQ9rsXDUTqQ4xTFrvkbtlW9Ad246AI9fbmDFmwwgfyplHX/dy1Bg8L
9p1YMQY83c15qVXEQZM21xx6EJA4gBCQ2McyR4L+hE0dv3tClitEof96BX4gYXgX
sbtqR0dxVb3Qe58KovdS//emjmcRIIHq9vQslyyw+ikTXKyngeGAsh/sFvj+UMOx
bzqlkdhxzs/6RnRA42dDdOiLGWeNWKCcn2NyIbwk3QAWHlJVSN6jqgsgS6ql6kRp
FNoH0PVYEvz1E4ghhHXSrswlgoKWnT7lO03xPOPkAO9B8MT3Y/G3F33mXtDdxhZ5
TLbuAJuJx4tMYMZBruA+VGvZ4R3pE4VB2+2wFkchYNqSQY0wiBHEtCZbyd7k9Psj
FBlqV5jp2qo1MjxJk3e98BQ0WjE3YCW17PedMagU/YVtKkHByxpX28rBpMpe9b8H
XGs/SecbCtxArDsIfdxV0aqsn90QwQwpWgORG9YTlBscPkZ0saNXgNpLi8bylwRe
/eswp9hI2YV6Jz+Q6sE9nA32UsUCEzU6Otqqd37yu5iW3dCeOOAA8wS/KE1X7jO6
Shxihhw9YVvcV+21ISyuIAQce8cr7WxzhhzDEWn8jJNF4VdqOVLGNx6765Kc6Hea
fX7lst/RDDsi4onfD10WvT/rKM+QvSpspG9FkaisoWtc4v0TNe7dH89LC3qfFsm+
MfjSgn8dYK0J6637z/IORDZmINHcI53p43vqki8wAoF37nF6ueNgk1ix/lD7GL7S
5uDvTvVTIDtTSHJhxWDONFun6ht44Ojvvoi2Y7cpIphmtaeUq51cpFfV4LOaRXe6
hPVTVIJ+9o21IERea9vlzFn69LW+jKYLlWy4XkAaKVWM5NBWS6sJqJDYpt4QGfAy
zrPNSbZECc+ROkB/0ETF+qkopzu1QcWm9peMWHtb5ZXMJtwOLdEUYsU8RV4reAtA
Siu1G2U6MXGjnwb03xJVNNbEfHE7cuFKUG4H+X9KDbOccXRc65tHShZpG4SZdFPm
DrFI568e71yWLy/FPlvwotvGioXqBIa3HDp2+8IHkqtg1zC+T0YDBAOMlyljQG0e
vx5UGX561FlrsiIom7T6JjuwbXnxTTjX+v2bvtARhmXD9uXjwAgZuWfXXkIFZ7Y0
3SYKnYpknnJGX1nzqT6V/jrDqgVP+/HVF0JefytIDgMP1MMNUoHmwyfbjByGGQq/
wvY6+kDQFBfNF6saQG0yGNA1f6M4lxR9CK6jHtlTZGCYjkBSssgo75GP8ark5URh
iB4LlOB21rjutUMxhbgwuwpQ/qR8tWloVCotodILnDw5/7yT+tTqF1aNBtXynLBO
q1z1SSR5lAS4raV8e+xLX+jPlxRlKj7VSbTD9L54xtugOmmE8TfxE3dT7GnIC0+I
w9d+vNCNKuL4033X6w9yPA5b/Ktkmu6c5k5i4tFLb2DnNXYFXvGUNqeC+JAjcf3K
gPrCYvT55BdafJK/KqYbpKrGoHOEKsbL+9D9ed+ADTP6mXVuMHVzR3sD0BhTaFrT
E16lJ+B1X2r/7oIbna0jI4Vai4kLdDN3jxlGghTnDBgIjHqI9a2RwIJA2ZuuyKeM
aPh+B4z/39kTqqVLS7P+p8LPpcqeihBuT6R92fpHq90KGnPvLtvnqR6me4lngrwL
btytiVDDJrszhzxIoYmYdZYcZ3ODYhjDV0RvZmWdF60AAzw3jLW9NzBO+bElRmtz
u76UxxdJ69hAhRg1zsm5qePXawolc9KlrRbt+uEzlR/VIyC9GatBzoew0nuq76zI
lDqHHwlDJsmyTlpk+kIHxaknsE2C8CS5RIzkFt5urOXS6FmitX9Y0VmUeHysTv7O
8dmbPOv+s16EzOnyN3zmSFR+RCONVkA4AUOEpRN0HlDMGg7wOE1xXq0bNciUE5Qv
CYGsCXZkcAKQL7MkwsvBgWtfB2UL2Y9REG74zC1U1jQNeJLrVC/t0YE4L6Z5uWS6
XR+JeqbT+oDHTE2ikbNNtUn57pEdefVuZROrxB2X2kHlIUKfxKEhI/qlhW/Gu9sw
gzdRrThd4hfboGXqOBDj2e2MAytQhASCxiVSlrvq2C4UhP/0NwOhiWAYnWskbN9s
JttrY1+GYxaPeSE1mBAmy7+W5WNpX/yZftFiNr+ZEAKdpbQGtL1QiaRF68PetAfW
2pR2tLrKURKEZzMB6VBrrJE4nPcJL3vBvA5ypT4S6Y7GiI3U/OA7XVjh9+ymxIH4
TWhKbs11tWqWlXP6bqW2UlXjCIlqnzE5pv4NTv9oSZmUISMgot9xeJIywzarA4ET
2rocyYq4HYBKOQuujzrVdYlTSCZ6zd3m8zTjP6yAuJ9LLciTvvPSn+GPZurHc5AS
F46z4tdDLaQCbeawyrNcOEXiZk0ihLaTDcudjFCg1XN3k8xppGY+j2jhm+N4M7pm
YJy8D3echEfq0E90NAUeCH/STV0H+Xk5jkAwbbG5Wvueo18wHEtwu7oSDdJ0l31C
nH79kHEXwndshRYibo3/IgZYAX8oqapurOmtScpvKH8fgwGD2fUmIJPhAEe8+oF7
/VAYkLoaxL/wgH+O5Z8NfKNOy5ZZ4VRedRsHqaqohauDFFvuw9W2sTBces9JfMPg
OANiD77/XlHUZLyiczOtWYmlQ4z5k3UKo76AS+ssd/1GnSmcwsfgY/e7VMEu/4jM
zum4h2C228/se3eIXvgjbJc8YBc+7puWBTXNNY1kyZVt0PdvY5VT+TjNDzRYe9Hb
/LRunWxMD1VVsreGRnoGRUb2UF5un7PWwQu5IsuYloI0Spq3WD5X6jkVyYTUviAf
ZlxJdZ//LMB66Uq+6mafAg0MznpRV6wVnWXitFVeXc7xFibIyAJpwlxLClrN5Z2e
62TERcAxzFKSm8yHK29kgV1nTjxsNYEKeUgyI7vlYzJTRIv8mIDMLVweag8jSXRV
DSj1Od9T0nHm/MdLxUXIA+kEwq2A0Lgr0SDtVMFVWRQ//W5LY3tZhIPsH2vvNW0W
8PYKvn7tkbiwdbY5AFXEoKGrjlLNm9q4cTjhrXbZO1bjgLBRHnMYwEAF3JbKYI0w
Cj9CbSlVLAnNKQ08W5npdN0wftuw/tNAmxuQBCoM/d7anEnKdpUV+90vNPuF7rqi
IO8b3nZk+Maqi5OiB6OF/8iJ90ADJByADtzggISYwucDtjuJk3RFudeKmbKO+BhB
yjI8p79o2+cx2Bo5pPW6cAmCc6OqesWK605ZoeimINh5MHgwrWMHbl5vUKDF0z1E
Drce3pyq7e2Rz0sibQa5FA==
`protect END_PROTECTED
