`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5fqF9UYR3PijpAxAP80SGncZzZ7uxAn8TcUB+B5rbKXtH0sXNGJO76yuBwBEECzy
n2wQkFc2VhxQjbAULnhDtwYhsAL8GpuvVzZu5wpWc7SJLv2t1A1GR09+qfLGJU+t
8yfVaxsvRdHW8ITRBk18RC2hmBe2h9bVxN3KbY3POWQov6AjSNtj/tB9ztmlL7dH
FxPFXEn7GY+ZsxGpxhMHWnlI+r09kbY1cCih6ajabeoAZ/WIq9B0f0nH6VdOEsWl
Ue7YSbNnxiu5+0J3tx+TRJbNqOe8jCy0z4Bi7rc0KyFgQjUCf9UyWrswbrLJYKXx
`protect END_PROTECTED
