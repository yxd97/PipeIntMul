`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RX5PzYdsxokuyYW63+VUTc88J7M7/UGxVYiij27AsniXrUllGZT9OPtlb8aryJPp
D943lUzsz/j6/Ts1nZYQ5M1jMpLS/S6utbHM9/jgF2XGXgSPuD0QewVDYfjSUQJ0
BD544YZ8YoNhL9tKLF3UxnWYE/auW1r21YCG2SOyRWwrQlTQlm5eMCuy8k1CDSyF
onjtVTV8nubSvEa8TjNaQqgT/bKyTAJUvjE1Vf4AvKKvtrrglGRylnelefCKAGmq
HWMkDVWsYX7aBuLJRmNGqt2FI1fJFMaU4e1/dmgx5vbXD1YDoxfIEEzbqwms4FUP
MFTttB0UA7KS7YOoMzoFEzuyn120DOAOoOtv5XhVU8/Qj6BgtX2KMjxzZaTph2gW
wqGk9D1xz/E5a3gdfk09AzvypwDqEci6Av2MYLrhq7Vw1gk98IG+9cEofTUQxXxx
luXs1o0WAaXfYyDivDCIvt09Ct7S8pLOzgMgnLnTp2MoEnHNeitHC0G0fhlpOO2m
1ZubIqTIGsVYio6cyiLAQVGKwACkkQmlMe8uhTqERHlf2UTjieYh04GHMM39PGEo
MTTyHs+xPqKYiHANmzsnLkOGRq61D2dT1mhgwibQq421oqoIeRDU+8Z/zl/HoxLm
5xu0G8cRfSo7LA3ARW1n7163L0dw3yw9vy2G1vG0WmwRdysEnnSY3o9zqx/oiH0t
v+QzI+IkQ03e8VDiG01YILSzkgrooqsXMbRpn+yZ0LEv+brrOzegzZrPH0qlOJ48
Icpeg6M+YBrWkpwYKick+wIcfu3/+ZmWIymmjYOlvR7W9rSfii4DBF7FhFZEoCFZ
opxVWUb94D2VLuYyj5ranFNFmD0pc5PX+Jl+gLPsfZ64t6mOuGm+fBIzIpIXRuqW
C7Qsl+ifbIyuOiDl8FbJlNJwqO1svMqqvLOgDbZHmI3G6RO5Eynj72esUB28hncw
C3HwzeboOKXCH4oJmUzAVm7rQv6WfSyirOVtOqKoIK5OVm3SG9DgpfNTm/Qcjzcy
`protect END_PROTECTED
