`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKoFTbcC6cq4ub/dqxQfgNCPYItKVKk8wVFVVPfeesTGODHZrlusw1yYVlG6yKCf
VUPV7LXuRWBfMHYtADCBNSDGX4YCMEAVaUA8iDdE063mkfNpMoh7rkqwPtvmyXe7
p8C2p5w5gC76XYnm6QmzDX1v4ni1wH0Y09BKoXgeIN9AZA4/FXsKUAhvLLRQdVzB
yThxnt4+iPu9JjTdJihjaM7ajdPicc4JlWb+pBt0K+KGpaW3kRkv/3+02S0QNkgs
ELtPR2CyVUEqc/I1PieC2ZWwellHdFFhI30c9CdV84voN39bHYWlS1XXBQZ+YXrr
2RiWgOWMmXxD+n1pmG0Fog==
`protect END_PROTECTED
