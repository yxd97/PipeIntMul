`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWTIjqRw8Cs4XK/lluRD+maHZ5zVoQsHqly9s3LdhXvFevzSTISimNa7EYxlNlvX
/quAj7YMCfgSqYnoRhu02DHARnMKUKFg7TQj9IAZ2S+/n/zvNROs4SWfyfU1h+w0
7GSXpEOlMPLqptCWreKr4XVI3+samH8izJcskiZVB1MeCNNzESKUm7CsFVQxUuJy
M4sU6Idr/75AbUwMxUHEK6hjO0bOeQ0nWD9sHukjAJJXwiQHaGcosuCl7TaTNzN5
O0X2/bP4jtIzaMPewoaTYG4Rh4i/i8tqDz4uhTmW4iRXCpC/pb/h+P+EfhY3Hzkr
efRBmC+rnwhiqf8mAXRjYAis+jFNXz7orA6HVP899yFezbGznukiC35xLeETGh6h
epOIxgx5VuNlgHo3LBjFl9c87vMva9I99azFKMlS+nU=
`protect END_PROTECTED
