`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TT82AHVvbdK9K7uGtmlb3wWMyw1VRRGZii82szAkeqJ3VppqRDQxwSp1qlOasxYa
vYKRhXOV4scgCKzxOu1t1+WJFhNm+3pOXVK9IOGbE3CNAoPWGR4g55gj1LhQYHsL
IK8zPwxYP0MkSO/EYnp5iBJ88O10DUVOgLoE8jYsYYerDi7JXg8c01i4bp9o1GgW
fzjueChO0Bp9USXsZee8nQmwi+SEUKK+bosdMZ9pJIxBp7G28ZPyWti96aMnMkTh
1BGbMmTdy0Lbb2r0ykw2H7Cknb84wZJmO6bp3RINhvOzib0bF4ibj8b6/wwmAMpb
6U+GFMPTcjOeAAaT4k+EaFBe82+pJsJo3fsNblN941d0lhLbW805C9TyxVrm8qv8
rHXMuYqc0xyXOrZZScmt4uqiPcqO1Li+r1lK951zslWH4/5hiK+SSxEHxFbMUAD3
oVCFYxgWqG2HjvN7odjZJjmFSret4YgrK1vfzrXBbptjErizTok/zah/5g1tbXwn
+OR+I5FE5OQMBDaqbUoItspiG8lTSlhfH1CO7l0HlYDCEu5IwHkyZw+HyIqgVfMq
I4T2I/k0zoCdWE4glKjUCGtnqXXx3ojBMqOAp8AQeZg934yymhwqhf8NSNjVxrSn
24YnmLuDhM88e/+2OGk0dIxBj6/jI0awZC9nEMoegZ9DrfFxScT/TLDYkED2vZ/B
qt4bV1jQ6Zap7mGVKwLvm3qVYpuOfFzw15Jr1HmqCIJDdeEwQR8iLaEBeR26ourA
tdZVYJLkUmSNNwmsxbdpPlPiv5N0frrZly0djO2S+azXhzjmO53Sj5Y1Z5oSTiBI
tok3sgJiZ87E3SfQGd2wOlK1KVKyhZy6dgC2FweVBrfwLgq25Ok2j9Bi+D5pEnJD
fozBZoZ5cb3DTPUKeFeZNv3Z56s+HlOQNElABVS2fPMZLnMOyPS07+e6vkxYya6x
1cqzO4X7vlb3rirw9VNKS1VcUSbQxQACdXdOwR9AXAupkb5q3ihlPygdwbvOlfDn
+gYMwWlH0r6fglXT2Z6n7bLq6W31lKmxZL8SWnuW9gRtewbQgAV0wftGUFb+iFEX
mtkeTpRMaLf73kywX4RUDfq+nEjoFUBG2Ir4mQlIE4NeXoe5R0mIojQe22TPsuD0
J7KB9e2K9Huig6TDGfvImXR86lLTDCccISRSfoNdpX0BNhRmQn1P2DZ3PJDYlZXs
VQly/O9nClCMhLtlyssGuXOvURG8b1f+MX4EOlRKOypICfJwErKQfXDtho31rpDw
G9cSanLse+DKFK23xMuq4Ha2kCnCl4ke9FqW7Z5AMqcCSraxDHDps42mjsP3KtYP
7+jzG0BM1VrlvVfxdPHuamJYT9DLA8vHZkwtBF9GDjdyJ3NDhSlJGoH5L17EnlIM
gMuwT6BSQPE3gfhebWBFij2gh1Y8jsLyNk+HWzKvvDBaMWNgutrOHc6/0IScz9s6
hCNtFrMSPuCu03OZuWTjLMgKpzxerXNI5FSA0Fg5Ti+CcOXbLHE/GQ36RllhXXLD
fd/VFd2p7Evq0QoDjie3U2sfNh5KULwxxR5pBQ4fVdpkhTvK5D3/XsMdjr0JcvbZ
QfRzkxssxmqjF7XCJyHCPOIu+RWHzK4Y+n5W18mqjKAjxH2SqxCfKxrubihBodZv
fSXouts/+yFspIoCKXdXWxe6Hh9up/CffM2C74jn8uua4yd/YSPlAauNscLDAtr6
/CzC3oOBoK7WigLBKxrONvP8ZcJt2LSWtRNqrVeasmTQVah/t1d4pO0ggEM2OzbN
V5Y6EwGhCfWiaJyKugMKvv6FdEEIWJCijqYW7cJx+WfaKiiuakM26n83a/heomnf
XuYkWieA11e9+wDkXmb1F4JzWDgX9vbSMHsXyvcNWwRwq4V12CGQBMZAW0lIvSrq
kpXaIYjjo2XmCebiL8toOyH5i8puOgsVldi6BVwROXZKgIMLVAj06o5cFy9M7zug
fflw9DPPDb88NYh0Q2tliwspUvAdKesmDNlIPoItP+rpG8bPV9iwN1MtJUr/XVg2
PHHmc8ekSCHDVvsTA42TbEBKhA4Q/Imey5eozVleLChxXRO3HoHIO6A59g6zXwAr
mNJniiko2aO0U+eqI/xOdL1Zma0JJpS8lxahyAr1L2wOqoHe9vKWaT0Z6WdoNJfU
fbtx00g1jTgZAyoXF2gAD155ZIs3C++AQdyWqlO960EOs6mpaHEFtNnle9pH9JQ2
1PCBygRZ3MB8M0FgttJ+ozcmlraWtRjt3QixfLTOsBDp2VV1Q/UskNXhgLVnb8om
I8G/8uvpgmiN0bx5mg77t7b9STtoLUwcapgjeYUEBZLMhMuwai71Dk9BtWXcyEtl
zNZxUsQw+RDnc9tN8F/bEVv8oQgIHUeUncsrIH6VovYYC/zZ6hU84tjw0jpITr/m
YDJXFgzF4zkkdMbJmI8nQYVll2ipaaDaanfIfhRrThs3TMiLPreSd4AIgstSsCH0
O8W7ghh8YtJow5qcgCEZnRacgpsKECMhsUcqAbZf00eao+AtwaOL1MWQcVYbHKZ9
fLvU1iBNnw6meUxMnUfM55mHI2Qi6hqdWqtc0A3v6L2MMfqR7ZhRymPzWuKsKsUe
lWRKPntTb7rp8chLIsGizkQfE28JgFjExGDy8QKyA1IGouXDbWQtIlZ2w6OLV6sq
QBN6fsvZwvqgsotqtaSDgiLKlFIVWOM+kTMKwJNDvJKebUbBn0QcZarnV/g798HR
NTZlS1SJo5/gRZkirwS3TA6qze5klRdTk1J3yRX1BRTDn3CFQbKdzRlB+/Bwjq3H
HXXF+CIo7kM7tL+OmRXHbxYgf3DnE5ZEMY1s4dQxy5LQNBezJnFmTS78pAU/MY4b
EJIAtl2wXnpp3CYSTZQS1ryCCS6MPhWXNdWWo2G/cQ4Dr1itmGuP/0zUSRJ5ct8/
KUAGPY3+CiEoL+K+UmERY2NPcTrEXgs3SMe4CSMwihVwfV23OOp1JWl3o+NVB59w
agPjZUGF0NgZpHXI5kp1pHgkWBAWrIjrqY3L/S0JudRqZ4AQJIl6VO8IJsGnVtSx
rTAgdRQ+SAdAcCcU5eb+ZdxAcpXYtQrfzIPpsSWURs6cGsLvTfATOhp5z5Mu+oVB
A+Bms+aV0y55tNB3WoLHPxJEK9HTecdvoitzwUYu5aqS4SWqtmj0HiCjXZzt9Ucy
oiDGjC7Bz5osBQX2P3O7V0jZMGnuqfzuMGi8Dh4arRIGhsn9g3oUqbSXonrLZDZU
GobmUiQPdWvbnoi1ryx6SN2AMM3y8Ote7PVeSZ6qGi82g9M/KHw0LPqORaNGb6s7
bYs++0bLCJ07zmtuUF7/hBWDCO68m6xBmotKmXfeqfd4r5NxhfY4RXJ4HrSrzcJO
x0j1zFD9k9dCfMAqTCCkb0PnL7Hh/Q5UL24WsJrGujrlT4t0xU1a9KkSdvRDEfm+
oOUOpoXL2l7viUAleV1k9oOqD0ZLx11ZvJLNGhLqfEtKSrw3K2KHWezUac9n4c/Q
tY/KTREXvGQC0gamU1hTelJVO0aM5OWt7ywiHQX30Y/WlE0MZwqTa4OZf5qI6tRn
80pne/StZ6BHXVUWdJPe7RC0o6SCTko+wDoR65wRbCP/YCU/JoyrKmx2oZQuQckO
RAxEt08iSSz1aGW2A8AOvZTD0B0EIzt15xSxt+iiKOG4sJ8LYJraSphTWDDYpi3D
z/jzjeBF4F15B2z+VUWMGUBDpp/NyblKS+7Vwb86zhNV96R6iPvdAkGNUmNJ833V
eawniyPipDBdxU86hmR+TF58dWO9r4N+P0c5kj8D/TnwgziFfMuMXAVmho4FMvcl
FmbrcVHp3/eN8Tj8JTz7DnNkv8an5qIa7/+S0QUmyK+mm1TxJXc8uDcBOYJdcRwe
FR/HOVD6IAZGKVU4iyW3Aw0aCMB6lFkQE9TD0T9ADT4HJ80JdHAT7VnhygCgFNdH
+cWPm5U9XCf7XjHEy6Py82eUGg9KVHcpWkANpTE920lRYWbLIjRbl94yhk66amJb
CUvPWOWbEdFQyRub5U/2SM4kh0YsfIrNI83gSmT+lPEjC3025IUCS7bNTDQElbrn
4rsql0ariQ/ZNI96F+lOA5LDCJo/2ebZr9K3IlTyLDvtrGoZIyj0i5NqWyeHVakn
MdH41J+tQNQFkFiJB2NUxwA3/XMst+I8bycGxB52VcAv3LLOR2Q8dwrEbiLwdGIR
3FFDHV9BG5nEqsOqGGtfylJ6KvPKpxxfz+jnWbITUMKOJkiY00basxhJkCiWvw86
s2B+7U0FiWVBdDibML7XY1Jm9tmbGOGgTXQNXuRSdrtESGiR9IpTM7rkVRYyZTDk
3AJIXDJtNv7iCDHkvgxPqW3vrp2F9zmYDCWlALio29ZcOulQbezGMKrUvp2NN80a
XiYxq+eIs3C302/vJQ/DLQvbBWuSxHdnoQ+1Of4hR3NhppbKlzTLYgUnHWqFLSFE
ReFuFhW7JHishF/qxACQNtz/BUCBB6zDTTezbFznwS8WXOrfvds+a4xlnfjb42J7
zgfISGRWzRDLGaOGmPVtwvUnA3tUie0qDHLDAqqjP5+m1Q4x44mE0lDKuMhPz0ib
GyW5Jj41jpumMYF3RgOkvmax5P+FLMhJn6/YCSNI5ptRMx3hnQAQMpksDYKSm91V
OYuZsH4cgWlpDyubtaNEHfW2WJkDDOSxG8VHTiD2eozqbHVWVBI5rxiTsm9vCJPO
M3Uipjd05hzp/qO+X3Bs9lwJrcq5mE+TyaXN/uFlqsToQP6CkbPTioQq4h61LLq2
K2/EDC+LlGEcyF+BiYkJAmil6oyyUnzD0d4ohGbNe6iL4OpDIbEbjqD1b0s2agdh
tIwWnF9R8qSDhxBM190MjgvfxRZfIOI0U6vTtwek0F3Nz2O02BxsnrcGF3lgrwzA
3EtDxSgnAX+1xIpu/1XEDNWqNoRxG/cvMroSt31oQLKLIwlPRBElhFJN215IDrFh
hLN1Dra9LdRDw85wSKQe1AHP2uLjSsqJpwo0ebkLAt0BIgPlnl5sLQUQeVKxmtC+
mW3q7dedPebbEcm7HnGhKWANPGdk+R4lUVhrEusX2I2uXeOmqe2SHmIgwpOaxvIs
5urq8jWoGMdyg37n+HkdjWTZt94c4q9gMN45uA1X7BjjkYbExZv/hnN82pjq7pAF
+7szQJWQfzvr/WE53lvnRyIHaK0HvPBuwkTwgBdNDZMUoyB7KhXebOvLBfIFbTW9
gxrvOD7uTu1m1DJX+djp5WVN2FTWr67KLQO/G0phP7zDZ3Er2nn41KCeBJWen48A
b3/z0By2Yic8U0MtQrbln7PAzIy7USLEHmaw4QrotAqw+koLzMfoyu1IjIpGsMmM
bKgIf2g7Y6FaOSJMwZGTOHtQ7VPmACiFBDY9HtnJWBebd5qtNmEX1m0dz6Ix2h8p
nTJh2KAIHNv8aRnwbRWy+LFtoWJHtjGjMpZeRxylA4zNYHA3ufsUGgLNEVe9MlYw
5zLSrwXvojhwCRAILkAgbYS06k5Io/azfONebSJ2upNx2Zt6e/mhJeOonVdRvGMl
1hY9bpwW7UVPn9mGjQnB/6qVJY7M3F3bbiak3+R+0PZwMOotxkxAP+ZPFfP5Ty8c
DkWyQrIGy4p/RXCze3NXO+co4JMVt+fiQL720NJg4rilIse8EIj+UmLDuyWBhD+a
3zmQEUnjnVCgSpfDYH/3H4R5JPdFK2e7YlzwRqBbmUUM7v5BzjHQ5OtJ65BAVAYv
qbjuMrPalvzYSRZ0tXhAe1GNj6tODI5NsU3tLKGsogN5cJLNStQ/uOajUAeGK2nO
wMIly8L6M/IlExFvzYM5cAiHiNRdyIEhKZaCdvVtT/XtdQB/sC7RrbpyQluxSTuT
61Es5PfKOvvYkYCuASQ1t6hnjpsVW+w5aoZRm7Q8ZfpZ6LZzq5t+HU0yaXhaDHs9
LszKLQY1D523IodxC8wMVK14Hw4ug+CDsZNrX/PdTZXP/KPwdQIC5slmDA/jZHcS
jUR/4tUb4P1gpBqc+KCUbuxiERFJSd+PO7HlZ2JdgH9I8k/tzNhMhdz8aJJCzrbU
mFbBn0Dsh8lVyVeEr2BRfveoMIwc0zdGLoh9ZzT9flkESBtfyhOGIgH/sgwDfZNR
fjn4CZatHN5YJ9+doE+EHWJmu8dZgRxIB6x/4NXleISIDkn7ajalu3mLe5FcLvep
qdyVdCd2Nj/H7t7WPKpgIeBQ8ibMGl2H9oxeP8KOg1S2tPGDjrwIe/vdLqsacmU9
W3vf87EsTGKjJyz+x1wY6WsQrAHOU+cCShpsF2/odzyAW8iNlcrxj/kGb66n7ZUL
S9PxUgOfB9AM3B6uG4hwIyvx1TSJEq2LK41VLI//Knl2PBf0zo9foYykuH3i5zew
eD9jgrYHMl3ggXk39gulnmJu0M6bKvnprp0jKJmZIUHLrLeRVdk8ajkIeVqJ6tL6
eITwxJkh/dal9R8+PwCIC62jQc1ZIGJhhZncY4oQsXGz52F9jRQCp3lfsys+bzh8
gOpMwWmTK+DzwxrLT7sDvrY2wjlfEVzZcRJwpgaES4dvnbRTDKdhpaCN7Yva8uOW
REWcAR4MvhAdkn5QFCoI4+4DaPQCgGgd63h0OiWagao=
`protect END_PROTECTED
