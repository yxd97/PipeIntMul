`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xg+gFwZ6ONZXIj/KDP9dDFK1/3fDCkC2yIqLAV4wMzaD3RfmLJ+RThc93/1z5/y
j66mIM+E37lD5DYNPEiyS531VFuswyBHUq+pNROmxqgboOH02H1aNwnYzaK/u5g4
S8EbyRmMrTD1UvtC5OyxQyUVnBuZnf0mCtjM1QN1q/wEF0X2AdVeXUwY/ovznrKi
B8SAszZZF7UHCjtBtHCtDEDTqFmowEZvTtmK67kjZF6ZAmm3TwV33fHRRqn1x+Sr
f2H53Pl7zC2lep/lUN8co44bh/a4IQbhf9WzQFD4N7O1zdHa5cT+jPW0YJPg3CMn
ZMNECtNTxQBGG5QsvXhJwjCXg7RdpRjbk5zHdrsEx0fkoXyfZAQrEpl4l2hjDKPz
MHJ4g+1js/KSbMBx4rXd1Q==
`protect END_PROTECTED
