`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cEVK9fiSehpRzhvuDCVarRmwj0GDjrmgVX5+WV8yNJHq44WxR1XfM2tFrzksNcnY
lP4oDK81u1CbKT5oWNEE+I0kJq0RBqCZXye6EtLXDThOSf+ryXMV/35jLlyLFsAB
dewMwaFwmgW5Loyfq/+lIUSflszu75bJHIWpEEpAVxXr3qX+go/mRWjdtc3wS5+8
v/vQrzorg/p74ejX2Xrmf4vwOmSNBzlj2Hh464UNFB5o6MJC0oBwE75jsOLDwT6O
hwsyfB3smk8OFrnQVkMHbw==
`protect END_PROTECTED
