`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7D5xNFzJXoaTXdGKnqchHznKPMRsyyhXUuGL4MbndHt6+wbbklo0cxRZ8biJ7Zlk
X1YHpiHsZAwe5OlsbvmIFG4MMRewX1JzUkvnlq3iP0/jw1XzLxRg/jtCXXuIYncE
tXx8RfwjTqhdk7hqJs4kmBSNN68JC4tT61xUPYMPpHhOJdeBoGwDxyFb/qqncQO9
jiV4MFp9xeBBnzDqUb3PC6ooxVU8FFXI+WysyfpI2BopNg/Ed90TQtM8OT9hUmOm
VfLMbLGTPBNQLLn9uB/6AGc8VbT0iy+IjMu9jJ7tLFXkRJalB1LA6WCqud93Qh0m
5vNzcZJ813y1yRkSTAKy/YqDRuFK3RVSe/BNQ9oinJwwJ/uFycB2OfrKHJ9PKkge
NUjhQ/vizB/v7Xc/E/WbaVI28Mh/hpR+sL/fb6fPh07uJ5AvXOKDvqaLXINwnwG0
1R+ofOke1WtrhF5gGBpHYzkpBAZlxLMxIN45+wpxdxYcQYpVTNPUbjbN/EL9rz75
n/35gfZqkJaG9GMyzMxwH69i0KDt2KYS/+5yHM/lLjAhG8vmt/giPgK/MDERF4js
QEPLupYZUOwTS8b/B499LSy0Fbn4Rg+Qs7jWPOoDMKISmwTr7CB3puCnQiPC8pgW
zP8HO/vC6UykaWhlj/YzxOWlfrUcRUqLKJLO9uIKseY3bi4aZnAVKPRUlART7Mar
iQ6F7Wv3fPVRptTcWvEB+gPiun7ZqCV2iPpqK6TT651Ik0BDe7rIQkMDx0tE3Olf
A1lbFDjuL235ywNAsAHV9p2adqFiyArXtzCvSbJyWC7E3/97XI+SpGXFRkolVdyM
2QGBsbK5jTvEDrzhjBqaaBTiH/t6Prg9uuf+LeZV72pID48uMY5zClVe7X7h+i72
yLwKpgnymCfKbU4vhzesDWnWGvd04fLdl7hiqTyfKII=
`protect END_PROTECTED
