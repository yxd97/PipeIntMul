`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e7HnUPuQMOwg8qguGhNf9afAnASx/2ak3pLUZgRTqz96lM9HWNALY9ZWnKLPzOpI
ywTe7V9zUMnnrjy1KGDNj045l87c2pt0yqCt3sLkIhhi9h6+toMSbuB+wn8PfPMD
IS+V3ggJfSlOYDbqXHKV3ssqS1q3Lb7x8AE92DCoQAdXdtSCB3pLNprfqODdiya5
157O5mngKeuUl8Q64EsZJt/FIZ5NWnAsxoJrsgSrppkQT0XYJLMbBd7IK7peZ1wl
4LfOXh0MP2ZpsPmQKDCaHY1DWa0Wh69x1HJMqLbwuBp5CvFg+6r2ijiyPs6uyBu3
V6jaz+YCPOZV49Y5Z3leQBBghWGtihRFw9+Pn5KwJ53a/OXkxgCECYL+kfSpDzu3
g1LFvWl3WyM7HZXBwyZcxvuS6NHjKT7ABXmqxIwyBl7J9RReBJqmC3If1NwPbaHI
ULoHWPBM8iTsOKcrA7MTHqJ4lXR+qew1tCRW9108Q2q4dv/AamRSu4Fd/syQ9Gvu
36OtgRUj4jCHrfzveB+srlb+IcfoeF8jBnJtXoqaatg9SIY57Vi5X9YeNUZg484D
3+HliSP+Bdm53wjhcRKicaY6uWsgKgTpdNUKYBq+O2WKYOdn0/A1iOazzY3stBVU
mi24/puswFniYwgXY0+dObNuxh5PTo2MgdlBIIur/4uUQj58UN1CG3zc3IeyzcaK
`protect END_PROTECTED
