`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e8A98SpwoEp6LHYt3ek+Tdcvrujy0EVShHG0bk7NWFOjjstA/g8U7SvdclvRAbEE
w1cDBh7BAxQwV+LpGFFqBdS3lUDH49z84MT+7npmFlSJ5s/Zf4StD+PQLqUeb0Tq
w1CQDO1A2KzThEimkMDoFmNXhGFDVpgFtV89wuS0ZbAt6CuX3S+DuEMJlmE6XB2t
FQ87nMO4e5Tcl3JGV1aSPkB9KdiYNmHM2atKOVuceQMWdYsIKuxBGcvOxZCZJW4D
M0GPw5kygcOy08tN9ax3kNJRMDsS+UoPs3/YFNdH+JQm3EwdQ/+BA9eIxW4JmPxJ
hz+mSJ7aSuwUgotgiRM0Gvx7lns5HDKLaoRsUxfrFluVoKgTYZ+mALySJy/WaVWj
QUSec8JCpCBdmUOgtkLUdQzt0hvC3e08nMgU3zjqPXMOSeEFVPc2CNCMVt3Skv5J
jBZHQlJw574MXCiAMLgZgZBhkYe4dQOfwR5gbOd/WVdfyWBZIlqa/qa7DmE+C6ah
J3EcbvX2bHvyUBnWwSic1A==
`protect END_PROTECTED
