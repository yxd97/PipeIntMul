`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lR6KdrV3DtQLeHX3dSBvMklbRMX821YKyTXEArnc1PV8ePSFE1nzS5QxCRQfmOLi
S1RLkbiFU3HuIOahWZVZrmlDF2U9tU7MC7nue3hlxG9Uu1UQzB+aWrT4AXZ5ofW7
5nHylrk3+qru58tRsty4HYVc6aDvSBJhPqrRBaaSGzJmUL1KUTAKK5Sq5s+LA4/g
n8qKnFsD2WxZcFealie1odM6CtMek18V8/eHluDGnc2f7rX0pyOpmAyW/R29TK3j
HrJnPNNEzjWYOLQj0i0/CaITNoC88B1T2USgNoU3cTsSuNFgzbm2tapLrLvL6Sl4
9rd4Gt7vmHK5cWhQhrWejXbofBTO/HrAgOlIz3IWlVsaRDB1fl8Xf2LUyeH7EGCE
+/wiNwKvRCo9LdSrBEYQyJEq62mYF7pNx1w9LjqiZO296dAO//lS1uwcUoYE71hO
vjibn3w2/8LUYg6koCwZY9cP2GU6vzFJdD/xIrMvWBZ4M2wxgRShMW/Q+pK1GbQ7
`protect END_PROTECTED
