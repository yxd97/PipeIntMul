`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pfbbDjGBF6JSXp666Bqr01Tr53BGOFB49nY7CNHwn8DDuR07HT3AQOPw/DFSupwD
ucn553gHtp/9PamcOFuBRBgvbehNGtQanakO/xNNkE+271QzuwXbVx3lzzQ44CDK
BZ3btN5IY0Mq80hR/nyn+6JDxgmpj7rj1GkD4Ry5z4clYiwnLncqDnjc5dt//EWG
u1sFqoXchvHxwjpRexqNnMMa7pjAqkmq/qUdpVujcAKDqJaPva401Q3Xp+uZr7d3
iKFWlKzmysUxJoTR93O9a0nyydH3zVIOynF7kNkqsKTuiYymUsPqD/cIpM4eXtn+
WD+As+UYEdETu2TnYQ6LB3jk+ex/WVcOtl48OVjJPW6JVQded1bduNcQeyCK8ixH
NUJzXzCOksBsY+LRNRGAspg+fze/t9Sykh3pgrOR47TmQxOiTXSkhl0N/CH/Ych0
aNUx2WHppaFhJpSdQ2h9j/39FVDpu0bjrSsjIG1JVUVG2Imz+v4opEaevdYbQNyo
VjBvGj1nyvl3zZDyjDg+TdHto+iP4az3uqwzUQFnrfRk+XK2ddjsZlHHqBCecpzS
nJfx4BOauHfU7OuSBHXJnOrnYS+P/B4KnIze2zpRCTxZAwZFlN3syuaA0CA6quf1
imGQxeReF3X3QUOuDEbNe7s5mkWBZ+s+3uiGuIRHX2uDmi17VTiW6Z68NIVDzSOR
Nh/M4SenpbKK5h1/Hv7ByO8j1eNDDi0W/E2Q6fpQ5C9jsbAYUM/g644B434tfGMT
g7Klq716QxglvyZk3kCLHmuuWtl5dlxOvei093jBoNLZiQmfhxQn4A6vBVJO8rBg
b28iBqwm5becS3DuxnLtY7LAlwyi9l1yDX6CubKA32cE9T3HCRxVViQqIJaxSrUD
kx2NJBIUdJy8TcIfLaYLkx6izeSPuJyk3FCI90puQuo=
`protect END_PROTECTED
