`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lJikhtY5Ej9EqfzSMrqJevf9gHYyfyNrU8h2Egfh+QCTRHjs46i83j6XT6i8HGAL
a+0+dxyMSIqUB/lcIpDddgcihvvqdwn6Ytj5/WHuLDk8T8A7HvKU/zzbVEfuFfTy
UIlTOpM1q4f5Y8tnbN11dw8r1ulfyJHkm//Nz9fcixvblEdSIN8y8Z3kmChUl/cr
yIYtur8abEvhNZ6x29zykHOkclbDA0dxuP23a5fAiCzreFRD4aMIGERRW9y7aQGu
5pThm8Bu/IU9n2F5pDPPVsl4Uqmdkjy/9LxSU39q/XgTLnoIdnALJW1bI0Qmy85B
giVeGUikA8Ma+Dq0Beqih3/vzB7Z4IheA9iDpHQByneaR6DqhNssMc7ZdtJfF3MS
7R70LsTubtcB9MW0YmHWgef22j+yVGtcw7Kxsq1X1FsLWxyrRCt/5ZjYam+0AAN9
`protect END_PROTECTED
