`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwAr9GLmyVfWjvFzf7NHlIhyLpcuwu9+3Ywev+V9xzKk44/kIhHeQ2FssqOtnDHw
PytbdCx/q8It3/oYQRxlXJ+MlkFZtc7ynQaIUIytkPL4j7Co/GpaWukWAwe2V4pK
KM5IZ4bBBpMMWSP5kp+FSqXew//dioADbN3Hd8YBnG8F7uQw6kXejJiHBUzH7Axp
Dt/p86xWcGB6POosUDDl21lp8A2m8dw51+TCt6eEKte6+q49CbnECo+vaeKEteS+
3wQYx3Z0A1CVeFnYWvNPT6dFj4SkI7lavOp2LwcT6wavQs13AUPud4XFZsmy3EVh
nL0+H9PUfMiCJeQ5Maiov/ec8AGqLjWh+yPuZdpbp1MCx/hY07wsgo7aNerqB4BT
RaySuOZ8CEXy62xEBU7H6NDphvpIxnftEDYQ2Zx0OhY4pE7HxXINiCsCKoaJna/K
t/PqNFts1DLZyK21BquaIf26S6fqin10AFKMkM9P4kU=
`protect END_PROTECTED
