`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXWM7XTF8C61mh7anPcilj4J8XeZx+uo1hjXqs8CTTABLdX1ULUbqm5DwSd7FZ2G
Kf596tSezPfiX4lZcGSpI/ipV8/Ibu8woFb8zYN9s98Pt0x7e4x9B67fmhthoKxy
8pwRkwUZTHiwV8w5wZ3hlrk+0xioBi5X83UkE9kdhKwwE/zSugJmSmucmosC1ybL
xJ3jA+0cfBeEkQTApO7TsoXUOkuMUSiEbLY7s0lmZb472oEtrU8gnm+rYcgztWDu
fWCGJNa90SZMHvanyNUAQLEvN5AXSDSr9V2LLLC95hZiLSdWB3qVeJUg+A1brXhf
SKAAmZjeAugSsIfgW4X3DBa3suD/zzcGbDg6cYMuj6FJIYUq5pIn6QS9PoBk52Jh
SGhD8iey/xc8Qf0IhyD04Fm5aspXO2ogGmXEyx7aFGjt/KqceaxbVkn8sF+g+Ouz
Ai+74IK2pJuYDFexZ68XGPI73EYbk/8B0oaJFwBS2kt8U9rHwgpJRIU9wcPpi3SW
0mPza0ov9rsR+7TE2xvEsb6IFyAeB0+gag3trjOyrGw0f4spno68axMCcAvO0/g7
qNeklsUZkQv1b1Tb+D9qqI8TjBp9qlgy00Qbzps1s5PzhF3MmQjQlQY4E6iUtWmU
U8vDrXQAtfkERzQZVgqMDY4MzYOKalh0LmA9V7IMSd7nyQtwrKL2rM6VurAAwEn0
q5PTjpz6ideCKnhoL/Pgap4nesiSX4fwG8db2bduPcTRHAlLEmlDRzsYYyZR6uqt
SPscHbuwueffcCyaGgFLr1h7RVR8RL/QjwtoARiOHSbn2IzwB52nHveb+nHxyuno
tnocGqWOA+//T69fStF/leUyS0MIgT4kHRg9ieXhuXaIvq4wkOSajtnURhZCsQ8Y
JUepSJkZSp7GYj0ReTmMrD6bWvrw7XPc2RI5Xq8OUh4rCFOJak1eL87i4guyJa0n
jqPA3wnEVeah8V9n4tKj2jJom12eCH6rXp3zXIEu+XXcc6U/l/nIMf6VsjIrdS62
`protect END_PROTECTED
