`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiIQYn6AbLoo8YuFX/G+YbYhjyzq0JHHLPzVNrUMiuBJ27197rgi/F4KxMjECmIM
2z5Y8DQqoLEOxHMOwEYqEY4dxa9NBMSln1Z/s2FWNiUogG29EdFmzVDknBYU+/l8
YfuSyUWm6fDRkTn92S9U4kvMOC3OPusoLXApuy6J+64cL+24QLg/FFjW7HkqAvFL
HZ4rr1CNDTeuIU02w+a+pkqEGgykwJp+O8MkrmfGPDyOdqixy16aEv+HQT9C7KDT
UdFYKzBpVBA+8ZCnVpg9kVnYalCezs+iyCCn47Qjk26U5rdSmMYrulbaKP4wFGZY
f++NLpzX6NO/cK0mFN7XG+aDmDczvfmpm1/pf1765tTKYm+ydXZxyp1YRC5c1xuK
wr3etbxkSQz4eE4At7aNO925hekBnMKBhVksMepwr3V/dGQxZ/eSV0lJb1hRbzdH
`protect END_PROTECTED
