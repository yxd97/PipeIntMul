`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cYm2eNixrnJd0/EkyQFSwmInCd6l/3npebe7xd+IcbFSHBI4nvPo243aeFfw0JXW
rg5PcSlSaVEYS9oZ7FOPbbHNySuP4cXUqpaR6IpZY1BzLgKuM6605RbvrmPE2iUX
yfS+XwEwfwsObW3mpYxUtjbSTVqDvvUeYRqKRl2veq3xIg027/eimNcMUiNys3tO
QMKfN6CXkz90mL9nmcyRBlyFgVKYlTe4XpBUdgmhQFcOP/BIyNji9A48mOW2uUKs
bYEnDjbZWgCpnSjn+FV54KoabTeW/w0Bb2l20JH2Eds=
`protect END_PROTECTED
