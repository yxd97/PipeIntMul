`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9lUc3a6WTYRSfJloIjNymP9FxfQweBAC3Iw/ZdLWQ02L9/uvZduJBrphhCN1SfN
8wvvjBv02mUfzjHtNc04HNv8Af6EumUrxEoY4yCmZeLR/L4ne13TwwVRJAVRWcJH
I+kWmhh/td79zLXGY9reCOr+NHkaZnJ7vO7KbCwq4WQ/D/6C4CVLIS+PXASm+j4X
rVxhCw/r/8Xv4hJV2/eK0uwzarjNdF6EKh2tanl8KrAKHJh+wwrHRJGn6woiQgwG
AJ2lA/MgPXxYQLsD267P8w==
`protect END_PROTECTED
