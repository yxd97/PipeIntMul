`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkDpNnOQ9hlVEw88ZFo2DpdCsPYAq5PJA3qsqV4fCcnnhExxPJXTV62EoyII1+TK
Ujg8gKJ1rfJTxEj8Y/1VdrPKrpc9+fI1MzBy5a5Ecnr3UYqXt7CKQd7O6vObIg6O
r48zAtVFcUrWRMq0iHL8AfLP3sYXb1mzOCsyCifEEdHa8GUube/3+gPJMarVCrXA
BsAvaGX4bxiyO8drJxiz+A3FDPMbEFdRmwKVZa1upwYb3sucoOE634hL9iK1LXy+
0OMauOY1B62FiXTEZPQIIK2uaIG48S76HXw2M4Z+OmbCtJxVHuRSEGmk2Coqg4MJ
gYLomGzbw1MJv396Rx0NacDDRo4kKMxbOK+h/IlAglDtNF70PGxAoLyO0sCMbyHt
pM+9Sgghmj1e65dpMMqLG171bVqdwc1aYYqws9wHV9DO9PLJHCjZBv0bak5/AucM
`protect END_PROTECTED
