`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GI0ry3UHWcZPAPytOZdIWLQInh449x9hCEyFUnVha6jHBfdgpQi7CqpM5WYLgGyf
6Q78bn9pS5nDjPzViiYJEhHQtpzg8wSjh5kfihVhWQ/Hv9xzpXLoTr+cA2PfrqWe
HwEXq6tqLHjy0fu/po9A+YINygdU530eZKhC0eFRDGlmDsieEbFtYjML54i+jWYL
9C+QyQ1w4k82Ur7phdscAq2H0hr03rD1KuU3L75W+gcsA5hmffw4twc9zJ3r5D8h
pB9BtWwZ6DXACy+zk7gVIHtGWOH+mZjw2uLjkiipN0o01lRoR7/7gFJ5MgH48H+1
2YP3N7/LqnWD3aXJgRtp41Vw9WIcG4vHKaHwrgBRJ6LEEbvNV4rnZP7Jvy2Bl0qQ
iSsHnuP9KKQnrw3XmdeBMPVgR6QPd7T2piX3bTe4dDgUy0ErTx52HUxG2P9TLPhW
Ydn5TJ3iLLRNgbPxUAF43VSFOOtx54wtdz9zuaCFc+ZVkFTkaWfTvOnR4MXde6XK
JRgSJ/E+oT0PvONUUFl9H2VP+1kieXE0w+iCN4sHJIfjdbiPKhpp75yV7VimdY78
+nNkUxElBOERyNZ86l79UVwzAYVwkCKRxJ6cg1QcmfIcWyVvne3TbljYQQ/sazQh
ZquA/99zySiJazfquVQ8A+Kdxotp83iyQeHdk704ShdPL27qAuZGu1DhqaOgUs0P
Qzeygj2kCSe3bUxfoXqOLyZP6V0TW9f/Exy74nHuZoQL2npDskUMCAq4NEDqlFTh
nvc06MvI3FOw0OOVw1V1WFamdS1wni/bkSjKw0wisKEAT1GopLFtlsTlg5WeMqh0
I9dWH8XYFisNIqE1PooddPiz9yFTFgv7NHPO0sAgpl8pgmXeerJnes/yz+YDg+/2
m1txxnf6fZNFm5bzxw9Js+VaQ6xTYT1KZ9vHRhq9H2HKRp/ZgXuAZK8g8rHqlkgX
6dRxh8Clxgd/S9O+rKK14vdcWtldGrEvNJ3lmtAiiRX/jJj5rcBpfClIwSc3Ipbi
YQRhJlYNIXJp9qsQx2g7URruONH/q0C+Z+PXAyFt3zZSTtPKIkXjh47NInjQtFHq
SWUb1y0VN2wI/4GRFpC2XTaazSoayiIeppO+xfuGiXgWG/pmvJsdZvLuF0CJ8KYz
fEtv3kihWGbMHHFQyvkchId1jvEbi1n5Is29+jZm9VxnelR+HRgY9hG2ZGXwfVZZ
QVF0mOcDcJaoX+yaEbvoZYIUD624p0VgWDVbuKvX8XjDfajKY9R+0IwWaeXmr6oE
b4j6Axqd8ISHVHs2wvHGlTFj0uMpedCq06UM1z1pjp3o+x1GPK9ojH9LXyI47XIj
yc7Nn5jYYkLGwW9ZnekxEB8TX1ljFdbhAuaNC64sqZVZqPm8e3+2Ds861X9146r4
W65bsa1N5mXj061mMRHed1JNllA/5HqiFOKEY1qNJu1VAOICqMNlW7nGXZ9k4Mbo
rb/FBeAKHa0pMrldNYXoI851Zorb3k5CKLCLPikxZQQbalHZn1c3QFKBvd7x0i8j
BicwIQ4c9+++P16bv79y/jjz1XxKwXLfJ/oildmtJbzNF90XONZTFdwOzEW371AJ
DNVs3gV+c3CGiIWmyvQ61IrK5T3d3WRvKAUdWAx0nLRGhrLl1E7CeNxYT7JhBhEw
kv7CEVGLU8OGneGfY5zqyq4Ej6XMAQHYDB+v6EzaKCRvKKadP6Ua2uBeCauOHhzq
XsJpj6bNmrwWlycL4mtFUdDjy+ot3vtA3igWR6I1geS58b3GktyqhCXwEAK6cuDq
6ovqEXYbCZMcaL+8dXVDSvrDg1mX9l7Dr+JL7Z2yzPutprx94jikgo7S9adNca+/
+GK7CTRdUqz61VHkzF/DIak+UgSOUgxpYKsPY0VE2xSMyIAgZ0CaJiDQYFJtxw6T
OwHu/zm4lvIWpXqoPpuqKFSa9cZ8ws9fYQ78sLQ7hkxohX6vNrP0D+e2KhYIabso
RJnehPO2jo7LB63h7vtd9NLKnZEHl9lAvjlXRvBe7w4HKIbUH77cXq/F79tZarO+
UU4JIgLg3TzTOc4qOTz2jT+6mRcZsuw7y1/NWwFBv6SJ2oHWkD623BxfYL8inQlp
oYbexXJtcODD1mHL0/Fw9RIkoBHR4X4D/mWOSzeLgfySMKKT/hZ6eiGymVhtPaW7
9oYfkErn7wcFVC1yToQDMiSGs4ip4EfGH8fA7bZQbU1YWPTzFzCGfrcQguv/qylE
eWjriMkMYY1jYPxgHjm99ssYtCCOfMT0luTAliS8/JPFxC3P5nPZmkCQfG9oTKUd
Q2s894J9PXR/ndhNUF42B8uS9+8/IB52X5Ni4Fe9IsTiTyrPvfO6iwccovoDjpPN
fttrgs7WhvOHft0mxO0Ox/LB9Nk9Mh2AdJE8AExrmM7jpHqhP8dmDOXZHgTzSa5n
ccrmIcWXOf05aDga3F1Pmrh9CEhr0kNt/+CwbrJxHi5P5o+AIUvfN61nZGItRBlh
sAvNRiwUnYp3p4UmcOg5dRuEoPfopMEIZvQh3so3kgYoy+BH3wbDepDs3FaymXr0
wAwU8I3MHnq67a49WktX5DC4G4uclbtw+bipcqoQk4Gp+D3WEqVZ8+WbbyeNgfis
jo4HiYez1OQ/3bndLvoju0ayDIFqeFMcpwk7iHyuCXrp3Re5Lalc94SRfj5jXYHL
NF08iwtMsuWpzUd31rCSbvxkRRxMVJozg5UZLCI/orF51hjA1f/IbeQgrloCwH2z
WJn6RHaeWRhqtUv8jqva0VUXenQ77btmVl5kkSIxtigjnqnw/9HnRbidd+oQYwIM
+mT+ky91XMpIDChFXACPomqTKriT7KEl6jOwfZQPP9k6rU8WwkfO7R2oYujZLDsx
CuSv1thlNFI2XPRTH/QKIzS1oBGRKuwRedq+OWWhaHcblr74jD7YpxrGJ27Sh7lY
g1sA17f6UEJq2QzaxCv4AQnELxpSQ4yX5lDPkcHWAJ16+2PbUH8SSshxpXnHIq2W
/s9yTUa3/t/PFCtt4cuq56nH9DhtKbrqW3dAqZLYI6OYRK/O2An4aAfEbmt7xUWb
oLfzqai/hknTPKWg+S+3zSYzL9a/YF2vHJLEALV5yim5lCzLQJFjLa+Ym3/MDiWE
8Y4NxW/C2Xv7LX1YEjZ90M18Ea6yv6c5jnsy/86O6sLCXZ+vhU1pKfliHsO0YQRT
ZIc530DP8Nr680/7/q+HrWTvEqIBnNQv3sWDXThRjfq0ayzJV7nQ3oMNu5NXb85Q
l2sIUzUJrewoRgxIoMBXGTGgWjs25j1iWEpIsFT7ENMZq8byO6zlHkU2Wqh7SAvG
njSQ7LvRef/LoqOq5W2cVyoXdXLSqma1Ey3vxi0U+yn1kxpw8pf2kWTpDXIG2Sbv
XXdqP+rL45XoKMT78IJENEml9LB9pfs6+sYHNPAbyd5EnVOGZ12kATYJAyHqbUZY
lBRQs5rZXg0udS17eKs2R54/BGXFVG1gSAw29odCtWCfD8V0pUfiedCJbDVRoGv2
2age7fApILMXfQpY6HGz/2zEzl6pZxOxqR+jXRIeUPapxCTB3gdMQIUDoeCjpMCK
17PmWToZnXTN0Eh/ODvnYhSY0zA0uZxdKU1qiSzPCnXn1bKoeuuuVa6aRbAONi+8
uNVIA9IfFgIGb3fRWrOM2echac6u91H12dzjtLCYRZZumjociVYGhBfdmtnTIaI4
M4pzP39gxr4rWxr00vOS6pMGIhFx37aOptBlKmTukeTbrH3m3TW10/Vjmvr8kYXG
pokCQmj+rXCU/42bM9fcdrRSsX+dVAvtI887PAl5Y+ENbOeoI0QqxeRRbjcAppYh
+r+RtHmphtutyoNWOmezVfp8adbIdr73/uAm5QPFWD+a27VlHB3gT74I03kNV0TC
IcIexOCAaTx6W/mRgKqopOP7Jf0UAmSD9gW0cfLxAdFkTDdNFVIp/4Uy2p2vqAlU
wkWLXahLHqzZvQpWRnnEY/xOFLiyTcQdTJvVNdO2wk7+vYDyErXuITe0VJ2kvLeN
IDSJA4Pv7SqyThbWMN1wJht1rvFMLOhvDHB7oZ0SOhTCe486NZyqf8GvwB/NCOe0
eorERAJJ4y8DwehPxma8reRmhLhvVqn+xjpg10wLEudmRoNESkNNaWCrITtdy+3k
ZSxd6yVBjAdNQPJKAYxtmFhjAIlmNEU8gUvD4trtnIk3ezbQ7TK4nEnwY7SfqFA5
WIzY1TS+AOeY/otUXDeAcGlX6I1q5ZuKdABTRDw/OmcuuNWfl5416NhGxgeZRytR
vvVbuXBkAFO3WOR9a6v8V6mZaSJrbBxeJvZfCDOnSmjkCECI67FAoBZRSO3et5eK
+4RtWfvjxLHothV18RRSLZ3zrT+MpeUROGS/uAILHHUCzBn3Iz4eZyul+jA/OTmZ
lLCPBjPTgAKbN9V/lrdYBJFjCJx5rzaUn8PEF0Fp9HMIMpQkHwYx8mqObtxNbL6K
mafwuzEFQpUsK/oy9I80hRa3AMh/QKEgTd97oL/wCnxHOUkpYJSqeqr6bMaorRj4
Huejz5BCFIOOSgBkXc7Ry/uOzZVbo+7h6A8SJDLoV20N070HlHsr05GFP+Rrmu4J
hsez2A+XAENbycH2/PfPkd2i+tq0jGC8hmqT8pz+PFiirq9LKLvSJMHi/C1NjfGS
hrbN9lce26dQuBO9rk6hcmxHz4YBneJIAf7zUnAZ6jYmhFhVp3JRDCOEKkEVzzyE
/BK2Wf6UN+m9rzSKlDG9Ug8WlxsxqvK5te3Lzx+o0GfzwoZ7Wt5H9n9Qcw7e6/qp
J9FVpiM7uj9b2BEXMCHV5KyW6T0WYRonIlE6/Wnc5uCfmbktQBvDiJW7KTBn59JF
SlQXh2YWn5tKhi3Z82Z3UdkoWUT2JmJqRVynsiPU1c4dM3bg14iwDFTgegkXyVRY
HOD7McR29PgqQ/bGp77oXU4+XiPno0/mcWbflgku8vjTauLOf0hwK9SpFM32hKZt
vJRC/PjNcyNqhsY9s8WgeRxrCgiY2UGG1yYTrSq0pJZ2r3nXiSR+5G5wUpN70j1U
A/JFpwtcJ2NVQ4dxqzDiP8W+yJQbZ4i3bNwbvcQQ7lJPr11/XIdwuybpVloz74eE
mnR7vZNfyqY2lMv2Ft3QXZlxkdNvOEltChfi/PXmlevfI/MSD6uXBMv8TKjh/ofp
KkuSjXxHZnUPb399/B5I69bgJoshy2kAdh1RoGHFhZdX6KkL1JaHv5Zwl2MHC/8M
LyvxDekUjp1/hH3WnOONWvZRGb1sFToDcXEu657z+2WWMp7lso85E7x22hUH2ypI
aIGPExQwl9iDYEhftNFkNA==
`protect END_PROTECTED
