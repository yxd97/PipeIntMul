`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCkBfFgFdT8FpFRpn8gN9u6a+5gOx8bSdVEYPqoy/wdl1Q8QIyb+0pqkq6raxkGn
GSpqpoWY6/4635j7iGL7VvVQbzGAIoQx5eGVxgfw9HPTJuF+IiROfn1zSFEdb5wf
sTiejUEm10qUc0aAqjjYDF59CXBqzogXRNDtjMqgbcVlxZVQglNO1RNHPmL1L8CN
wkbyXcj6zc3230FQbT/k8XhO1pscB1BAUQQc37PmE8DRIHBvv8PRTTL5DLyRfzcu
Z4IE2t1kuP3ah8hbiWkC8JK9XaZBfrPOjqeBSR9MZBS3OQemJTmY4YMEEPevzELo
1pzpnmGmilU1Ij+FZyH5urd+jbpiE9q3mQCLs2PS/S/mj00SWio71EJiErbfzxVt
XMSABSWYBVaK2CkRzxwyHz29lcZpcwEiju33xNsvf9/WN2lpdQehlpJnRMtK4IYl
4tvBLSjGfm0sFbthfsFvGQKHKxJZ3BUSHPkNR6i+awQ=
`protect END_PROTECTED
