`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7bD5HUB2YwxQmLvI/TNcCWhAUIxMJiKF7rbl5Z62GX+hdmFjv4B0xtaa7zk+OrK
CC3uMmQQYZOp9L5knyiCs1qvyYaaR7bztVCJUNyIGMK7PePzkpHsOgZkAH36J8dc
y4DzBouy9uw73jQcLjzXe1nS05+IjKlbkdfL6un5jthJcJ4poaUw/02rxvTkWexb
1jkagkhcsl0c3yXWPjdRk3qlnJdVPTI3sBCHjg1T2by3DO2SuviGWuVKYOT0iVNR
/hDli++XLr0Oh0IBGo3KrxyHNs73550zGjIM2YYkvOAMDD1FA2d51AAHrI7CXbT1
7TQFe5BdmNaa2PBH6cQtjkLVeLXnP9MrsHPnsWRpUOV31pcdC51KvWQfJ06O/GrH
/HXunDRbQPUGxppGhAHODH4UyIvBZAbrteUJYUMJBDuQ8ufj5bPHd/09NEcHxGOI
QvmtcTDfyV/WnxNBxDKyiOJc0b7/p40UGmqMPxM5AmzEZ7TfGTg6/5GppoDGyMiB
Zb/ZBAm//tgNqovs3ht6Z9nyZAREqhCBN47a9J9iafpy1ZpppHzmfLRdkgyfuluY
vUWreH2jLEd/EjqIrFnIkWFkahsJ7g6IA5WNKwcpkchDElqJCISiB/uNBwiKFyvl
6GkCVvEFvf1jho0gnilU4A==
`protect END_PROTECTED
