`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zRwzNbHCFSc886dx5jCxq/+akWBjdN4hIi7M9G6rBG7vav1Zxa3DaWLrctUQbutV
o1qdjL4+3g/5vuYp6pJTolJ1ayqX6aApqiMkPl7XLylXnrk1BUQW9lzjEeH/kjD+
Sb6ZHS5khWcYt0r+WOXuzZzFGqF8TUdvuEtbPcoz2OWo04VTTYUniIyjz7BgCXLm
apOFADfmI4iQPJ91pnEsE6/KjozHeQ4Sg1mRf6m2Ag2bcMLJzlY6amCyCQkJqpLK
PpMCdjD1d5zW5EKDhts+kn6nwSupxaf48PTWQgm3b2NTlH5UkquyvzhF9DNLRdkc
tSjJA++eewOszkEN+byZZfMICyVuHJQO9AU/eMzaVlQETk3d0hFhcoMLhIjILchv
CQO0GO0km/ht0iEc+XOHZg==
`protect END_PROTECTED
