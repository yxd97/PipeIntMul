`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67E36NriWczJyCLV0mXFZ8oSBcvR2+yCLnsJQHBg+BLPT6ISbV1m3PtNoiB/04DA
ltz/Y/N//D9lxsJ9LhC/OfcwAeG/DvcA/5BPx2zwdo5HSVmXgUJuGWUCEGzOXKrF
oqIoSNWqoL9RAaPpq4IDBecD3qDCc0uw6/CHC/0C4dJNPKN35H+k5W6tDOLm60JA
T1qB24kpVwaSlNj2UErGmhFaLiBAOI1+ibTetSo0TFfDG7fdnfHUFR5kObC8VXOV
V6LwTgqzKegM4R3lguSlXMzozLtkJGvCx2OdGgYsAw6flPrVh05IzqV9RkvCOdTj
O3Ws584kBV43HOCEJWZxPjR6bHWM0ns8qmaADtDNfrzwy2GDpH5EOwAmEkFLZQb+
Zg9Qh+fY61KPJJoB+ov9BKfZ1Spbue9ZGLMxUdUQoRW7BUbJmoGBBnmja2i6qT3l
AHrGdbYjkfPlhkQ75WJG6+3p7VALbTtKXl5afDsFHOE4x+b4fH88uHcEO1PQtZ8w
pncR2mVd1GLBE2PDpPGKqzDKrr56IFbK5NYoQ15CFc7uLCNc2RtfPrtSXKbw64x4
s1FWLc0hrCIyl1clJsORE+U8sTHbVPifMzTIKVgDFAEkZLPhCDbubiJytFG3xyyG
R817S+mu7BNb+mHRuynVWULpBdbUuSlRIpoY6RbU6+H4uurDuogs7o8IUlHzvDjj
BTD/rEEz8L7tXpXK8bSU31oK3aythfEWHn1f9CSKollG/ExC6akuMIog/3wYMPn0
SrDwa9fouGUKhw1hFOrMYbPUsYNQO973z2F4aeSvQeq/VXltHN69UlclXartgaqQ
E6nUcAYhSjqbQJDSjK7bv35/9GoT0f67uSw7LyPxVcK78/Ru1wBOBJwhN4G5w4QY
UMJ8fY7rVwby7P4fW/B+b6YrZusCDE8aYz+dDN0mvKPFNRXSYPqscVuFn7oRVzpH
GOavKCSOp2GoQ3o/mr0vUfLPgPMnS5dOj8o5gJOxtmEWjlODLPKp91BVtfrUocpA
uJp7/+1fUPLiUEUnOu15ZxMjNmtG4OexnQZohCQc9Ukih6FfA7NTQphrCv0t9Z+p
riY0d1mCuVlpkry1njT7QlQBuAuUU1BfgCZqzJqdQYgXUkyGiQ2AkNhelhhgtmcR
OBol/6Xq7Ya3/iClPz0URHyuqyP/FsGMP3ARv8ycpSZVVSL/xzQeAjansAhduzMt
jv03Zb98OOvsQDPPmip/iY0kMh2ANblCJB5vJZ9RaPFLjvBodzGGaEzgy9kgoD7R
VI6FAKiyac3vWfPkPcSHAiYIeNvgN4vUFApE0WCxLEU4S4MG89KaP6K2UZQLPvi8
cOeinmdAC2gdPY883iJcXhb/QUifz51aLBLnT+nBDKYCgt8E8xeLHAUKVaCP6p5c
OG40tynOixmJOc8lS9uf1qeuhS+tdU/kMx/yk7RXdYw2Q897wlHfJpt+p/GO07p5
C3Ec8A+7deKn4YXbrjMz3Bo0pH12+hDNlB72h97aeXRl/L1j0Xvnkwm2EsPRWyV9
/TonJVczwh3sjBMwTQ26prXag6DRzYUyAULyR18jmVvGzeLGsCSbJhyjECJXIi06
RO4enLCA7mdU929ziu1hxPzVvfp9fpBv7cDIqn1ZCwcM6DOJbtSXBp1bbdO8UzWq
xizYipyp023r+/pWGbq+UZRIrFW5eZnEl+BSNXs3SeO2eda2ShQhqdJ1IjmB5NpG
/Sh3NJfwCkxpwVITY9HFoEzeHIlCbYcHQwfTz/b6p5KAwRv3r4wWFb8CMSL9O1Ut
wmZNzFHciHzYhU4Ap72fmBX2MRQdC1SaHxhgY+qMOm1cysllLXqMkMHWgPvGfWwC
nJp9xYPa+oYRoF5//A5trcWdPWhiCq+RgQ4VTBsZtFseWo+ja2G7gw23dzTxyy3Q
y45CbL9sPP1irwjDm6EfLLDam8aYneDhP4b/ojX0GQjvyiOjA0h+RagMs9mZufSr
qudD2qO7tMuwwMtqlhccDh3uWB5+QJGx+7L9+FSQsEXmRkMV6h3ShQomnQwfA0Ep
ek1EssLKECVxo1wXnd6hoUn487MjetcjCXwBPu4HAywtdSmNrYgi9hNxSujFBZvV
3IVswoySvD61hueVKXtwsyWIQpdB7CS6+TqN4K1WRo9tJYkk0MLDlW6wfyQ6Juj/
4e/+rxcBvFmFv5Mh7m/D9G8EPxlFXdzvrjjx4ZpJ6m9DTaR04Da3wpNwFq/1TszO
gvZlylBGUx2wPAXNH1jM9BfzhInyZcrAP+Tw+df5xoGfD9V+Xuu/hK5R2XoxIjHI
9bfbNpQQ4281805U7of2BBYvf1JqAqt1O8yxtxbC/bnpv4YEtZw9o3I3YoBFZQvd
m5/g4qic5QdlEbdQljhrt42YrsDfqBXUHrm+DjB8/W7FPTYey3XVzn2ODJ94wG+0
9X8v9qam7DErMjSm/KODpJos4TQFTRR03fMjURVzNhCKcz89HTmQBhnYPENH4v0n
cLzoIVi6gIeuNQs3W/p6ccSEYuzMOsEldF5VoOOEVpaCBGvaXjiFm8NJQTRM7jPi
IYOJRka4S28EitqM2VKZNUaKeJq0qjE1U5PXw+4IBHIydg5HxKM9ekJV/6U44KId
Nmyg4wA5eTKdS6xUdob/7LWRBBwu1P+1Uxo0hmBljtJRqrF3sjp9RasWOczFjKM+
d/gkkq9VOrDJIhX1u944auGITwddauX1Qvt1+ehTRI7l+oJJkAGV6aVeA8yRpQbT
govXAWDwlHYGlJUkVbxoKTfh85Lw7r+gMrmgKznWCmnYrh30F+UaW4YkK11s5h1U
YY/UdHsv8wkxMP2yHWmJJNKkhfoGktTHpWFEl3y3RDbtHXxAKTlMXNKXjUL+B8vw
rd33cZ5D/EKS9ZD04XygviQCJmTbO3UUhc3rcn9jUOrcpfi/H+bdb3tppbDLfFU1
6y7zgjoVrIJ/cy4A1dept/qDjKVTl1MyeFM7R3s8kBZrTtDksD1lwBUyG2ix6Tpb
0xIu1u8Q78yGdUeWAeBUn9QRYa4Iu4tAFuKDwvSuWDtiXXavl65lbkD5adlU+XL6
BzSwGCTRPzTlk6quGag01F7k+vRKQX/K/1+8NM+OLTD7CVC0dWTud/RWhJwcGhNZ
S9nnjQuFqXSAVRLKSExrnaPfbdP3oZ26Hx4RE8Km2KfWE9WF8eDjaX74NXp+0jpz
X5plaHTWaQ87a8LzXrQbcWBPj0fIS7yJ6LTPBogC/GlDnvn6cUa234KUKrjA0IrK
sMaA8ITJ9y5VldiJ1SI9QqEECJz925+TInNeE6RSbIFxDwsdJ+/h+y67WIg6oHLR
+NFwYBNhq0joyh5lR4gjhpG5YdfdrNDXLjilKCDvouKQ7sfufZlX+uKZnmVrFOHx
zon+DBb7TFAlCq4fc4d9i1vswBMh9NDp9fJrvJoFoYgLTAuw5DpTPMABMzBLwlrh
fqBmWm74WY0lG2/9TLXCJ2GRE2dwBrZoW6OMSPMMtKWrZEOoJ7X4VlvdFDhwzh4L
ZOA+Pk7TGpnsrBMxIYAxxnw/RwFWZMDLQcCO4HQDqvr+MRkpXx4xJhz8sN+YRqJF
1Olc1DuCpLZolhOISaE9ik1TEvn0iQOWHGySaAV2W78b8Z0SNTO8bx0YeRPaoIWt
FEpoqhPa0ZCmzIo15IBFBwdEDSvh4YobAg2Op8TcxWV957qUOYOmpJahSH4S7cIU
FI8uUYGGLjk8nV5BNJWT34tP6I57l96zkZq4x9+nt71XBohgtt/JornxhE+5i+t6
Z341GJhW9pjiBumHA3XHjFD5kgWbbpwkBz/8N/Ejgudg/hrjQxl8Nk827XDqnMdY
FMpJXWKyOKNrE+JPkPUcgTAl002wsTp7cS9Q1paiEq50in7gT4Dd91k3SvNfAN6V
9q2w60ngpAcrXl41ozEuzge3hqy9bzeF3pZCTVXDVpl31fRAek57QupERMmxmtUF
CFApaTG4VQi627eGqNZzgoJ/3j+RoYSnsBdhpG4lLgk5KYNnGG3vJ8NzFfdE6WYA
Q33RPvodMba6A0pRj9+FNu+bKiIGkPcszNkdD5yTOfwo23FgmdS8pwLH5t4VqUfZ
XeO+1H7LTU51Xqv/wJUKReGWfiIli356dL7bgL1Wc360o7BSUAyxJbPh3M3Y5EKT
BgqeOu/RdGTuR/PfBtGPSZfvGn8YiHsc2qkLuijAwCLF8BZa0bnvDdwTU+gb4SBn
H5KjKsSZNLvQ8ej9UqHmNoivjSWIiNJl2k4RWBtEBmvq0w31/5z4kn+GrOy4pKV2
vfyf6N4FpL04HjcixJkFBs5HtkUR+rweFj2F5O4IAJHLaxaI1ibmCJzRSAkV1a3e
1i8W2zjBPV1qux8T8rNNIYaYA7pczPYSijVrIt0ycePrlGirX8cYBGW8KmCOy/pY
dn3+SFctLISb3hEUgYmHJSqJNdkXLOqBy/lwQOeNJyBzzezVUWg8K/je+3g3Ejvb
surwQT3fyT+Y/eZ5bDP2CFAxeQuYXQ9yR+SeBtqUbTLaBfzGSjiH0IzTngTzwdHb
y/94XXxRWlxD1FbR26tdBdJKCEyOSkhIO4km462972FOyq15hv/znKEkUmZ4J/YO
oDUOpBGfTdIafQPhI4LlePWbo+bYwefTXNeA8OW+uIiQcdgL86YHHZ9eMyZiyXS4
Bco5IeMMl8hORY4p2IakjmR8VP243nVxd+fHghmv67ladwUzP9apwSatxVl1wIAN
AQQYi4yZJ7DkN6wwpRBUOrkJvSO9lG6rxwVhbrM2J+H9VaDwLlJTl5z8d1EeVpiV
ZOYaCxcXPmmDPoCExVhS+HHSt+U8E1YSVZwVsIcqa1Ea5U2rr3/MpojciKUHlTrY
HrWFMnhNcX8l+hzm+iweFtf3WdKt+uaK57F+veviW/AK+E45j29tauBT1qsyFtin
t+iGU9zl7vO/vbfFnt9FXsgaaJmw67EsZ9RCYuk9EMBM10Qkbd3TVYJnJQh14x88
vm+XB2y7L8BZmLM4Laq8RtS+s/CPkOgi1TGPV7UYD1JOmwu554lDrhrhZgvDUh4s
V/JksyxqMeB3a45rd+78B+b8UWoH+NocKnd8bkTArI4aj9P3z62SjK0xyCrNMCdZ
RpGzyUHPDPsuWSrX6IOJeADkNmpDoLDkG2kgKuyt6izKsBCOpKxn60Tpk7lAvF3l
g0AK0Baijg0t+XkKeRl725wStHnQCRAD4PeFTVA/AhY/TZi/ACZqgaVl7whyq32G
XzjQaovmPZ3mmVyREjvk1/FO9t1+FwhlvxOThen2TZtYbF6VR0yf6TzeeX+L6fqC
5hPyReI5IwKZh/eMY4iRvjCYZXXBJ+0cuLzWMyUzxQCtpO6BbuleQUH5wjXWEFWO
+Hkf9fy6YVI0USHF3C6dqNsK7MBJqGANLL/Q3MARfQphp94k0Ow/GIga7YPrF/Bw
on8V19a0j3BZ417PIxme1DPxgLxLVcpGgGyamf/5xp5IYbQvI72mq+rEdrhZbAu5
cKAP7azHg8NGBhnyQ4nnt5cgDGKIxUtAGdJUSKmDGqM4dQNYF82WaqBZC+BBVp+n
pQshDlML283E9CY9V9qTfTH6YGYtRRvKV+nhDC1APSIJow2IjQ1B73EjpoLK73fl
7xiGGqOnp4YeouiXzCpcWGqP9sdDzZzCdTZ2QlTe2JMdaXOIM00Yps3pYOfOqzpK
ovHrRyNKi5DMd8cakBP0bOwKz7kSLbmPTkkFO/lOsuvN6aEmCqH5csi1pNOAujDz
XRJG3kHPj81uMoDbOOrWRQ1zUVC646nIOaFUyzZFf3//m/fXHn/v2jQvaDo/ubhb
jI7obKw32XgdnMLRgLjkRuPDE5D7s8GlPnMwuybucHOP8tPrGNVC8nmDU3UDJ1Iz
zIwmpCcwXGp2p1voT4yk0gnBNnY/MqzqOterAY5E8D7IQILmTpTdreQy0EQ6/I0O
XceLWfPtMGkjuikjkFPYsT/EGkZ23lRFeTEWS8LfZReSeYOHhqbainpR1caZgVkv
OL4jbjQtpRZmIVWtGHZwgxl98X77WA727fdq6Py9Fg9awR1rQjUd0XQyNApYpOEE
jUb1QW0G9zGCKSTvgxUHduxoNoK2UA3Qx5SXXC8Ci1ha5a7MwtfU5M71QQdmf4KL
KMqaCcv7Yi2aFTcToVlOqM6Ivlw8RMDkD2xGV9Yn9BPZxbipwnFOb473mBtFysh5
RtqlzD4U1ISCgvmGXFGe8ZXyRY4v3Rtlw2PIEk2agyAW+o3bYQjRM/wo7Ot6nULH
3abNzhRF/J5HpvtAR2+us2qQVTqpVcoI+tqfnKeFnWBYdsDwLhx42tt6+QnUgGr+
GMe37gWuqs1piqhrrmjXtAHJ29n8NtswieJpa4rSK064oy3cmXvWUGqb6nPAO7Dg
46B3R6Ledr8UY8vAsYszcXBAt0Qevp3ZSrIEqmdpp/oC7+F1UkfP6b5Sa5Bupuzp
eToahS+vDn8RSd6yCYtzMYSb1/H/OPGAOPlgRN9KQwrDkcaeHHYKE8T9mg1j9dG9
hYB+rK+AblqMWKW8i85OQdGnYEZvOPT0kgLY++cO30jzq0778oEdT2nKGySRgZnI
JSgLx8fm8ZpDA/ny897nTUJ+icNaQfmwLYaGiZtAcWEI7NS2UtRa2dpJQLsfZ++A
sF5n9zV30R98oqRZSZ+8QCteQQyUqxtXmJm4nzlwR2IPFoDEOPGSV5erDqIm09YK
Oq6d68W8hKIqrka1t31Mg5sockN748utKmfrV0nSZpdtaP3w3rtiApY8egq/Bdlz
F1CavGJhxoaDpNySVVxtw8/3VoyFoiwPwB8CX3CBqmo7xR+HT/p35dI1w2NtKe01
bv/DUvxLdc8JtFq0dOnmr0pu8GAxo0fJue71dG1K6F1urt9V2XIBoTpjafp6m/v6
dpwxAhZiPwXpb3lHSHS07L9U1BYpOfox++3TyghNzkYliYMuHmhW55FrBGrAjier
MiXReEjtGqqsRh7DxFP7UEDN5x7s6Zh+n/gC9WBAmmFmZ/ELmp6VImQ+jTktiBi5
3bbC3xEM5r8sK4F9vezbjc+hPZlNXj17TtVA8AHa65dIh0OFcF2TmrbUZpOWyVtD
qsxB6YEPIHrOAFu2VqFN/VrxMq6zqXVSUsSpjSMUTYLEcKecctu2a/5oHIJZbB7/
BKRmxdYiiQRIphVjZsfPGTAzas6TRoxJ/aK9RER/zI4/t6mIB8JgpjQGOXxXLcKF
42TuaHCCzTxuGCdYsn8oo6856xJkftw62Zu4X3jvk6v2kZe3rQGoW9xt6pdLM8qd
UUsQX3iAD8a34RrychajeuO1C0Js17bxDdaI/Kc4lcy0LxQvrAHNLWQ5Kz6XYb3T
x0L0BQ8NErqR5kXIVxBtLfnJnUbdvkOyYB10hhLdaAdLlH2Y1E2I3TkjismdIBMk
Xb75Mvi1PCyaC4h19JWXuXRkRJ6gh9er9na3pZFl6zS/HgEafX5xt1ESNnyGp8YY
C5Xuk2S3jhkfmxnfFB/6JeE/mlmLhGBILKH4Cp+L6e9WmKBOT9ES1iS5XUEYZ2Cn
UVLXrKDl6xYMcGkktS1RiPEKUPy95cFgHnDlDclsx19cOTcTTnyIlas+4GeGLUa9
berldwdSFJO9cyD9UJ4pR/U03yHXDNCVy3yX2mI39aHwnPHPQQPBkrVkwnb9dHMd
/4+nocnVbzOjzBD4A5DpeWgjqeEhvaPVsGKLZoBkRgfwjKPi91+LMP7Du1k2g7gE
Qmxq1wp/KeHbHHmZFoMmvv4x8EF0aPXl2q498aYTliaD2Fy60gXzeWOKNeWhCR7U
QJssWXQck7Awj+OCDC5weuAHZp1AqsOd8e0uAwxksC9jrpM0UGNorCfvk9lg4OsE
EWrDjf4nAG2JEw1h+m9GgidxzZp+uzlAcGsPjxyiYeBUEt1OCu8lbfO2WoIpWbKb
i61pnPLVGfTgwWJ64WpRUNmA3gyjDi8fOhXuL9eElGyTxx9D6GwNGWPdsI3U8RVa
OeRDfLvO6h0rzbmdbL0DBB2YPClLilADCkXemSsbvJ9ZxdqvvBYgJI3ftXbk9b6i
TvQKxkRz4bTrbJwcAq4g0uaOAhDSHxsLZk2+WQoE8jE6wwCPCxyA/TmPvIOy0GFN
331eZ5qZzmV7eM0D5cOnO58XoL7UBezXd3XvtpX1fpltxQdXYigBWtd3dS3obfZ8
PCYf1Gt4OSkF7K7+LqQztg8G5rsArV1kNe5JYeAu7pu+5W/AslsRP2EdB1yBXj9K
XY4jhWMIN49bB32WMPIpodWjMJAGOoRnVZMdW4gIcvxVLzgzmI/E8IcbnazXfBGD
dxlq2Q2pWIcbQ/9ZipgC7hS8H2oneiCzmeN3MU9GTdX5TNfX7OIVL8cMGUatUpMZ
Op9OMA4v0GqMxbaoJAyKBqceYbDpOr2GE22WOHCY0wk//WKaj7SbSZ3r38uuHQyI
HbLVGfq7B9kov8Z87Me1gnzSVeCvyC6t8qY+r6Y/XCyRsetAxWRAkywpwaxwtZGZ
mi2L9NvhhEv9eA7EuB4h0rxH02PsZhfstjH8C48rOKs+XaWlrn3QYgI7uQxOox37
Ftwy+8ELQHJA4eHLcA52JWPeEtMEgEuFF6UrFf1qUohntZcDP09KWek3z/bi8ZLF
/bRm3MmjMYG78ZMS745t3BetZliXns0G4U1G7X8HTDOlapEsgt5nm6WynUC2M6b0
RY/YiTKT13VoBPbkOSrp95z7AKTaUEOKpKRJvDXjexc8YTtb+xtq8uvx+qD9QiFd
h2xvV31Y6ZvgH8NUeMBCi73pLINJwJnsF5G6Zi2aVlAlzXpbPOzRii8HECsm6sag
E4pQDA8JIgXPAvT/cisBeE1R+6aLw6DBXZPnmnR010JW3XCjQO+a5+FuevTN+L3L
FaLesseOH93hehcPrRH2dX2/zZxJl+tImTQMSZpDBlSFpUYWxq9t9O/1u1VOJgeP
TXHWRzYN+k8ehOVZGn7sZAA4AbBmEBbx/tTcdFOM5y+rH8Bs2TMOdAa15fJbKxA3
jYhHXXWJmuoLUCaIn6fX92ongcH1ggpisRqi4lp3iCahxzqewBAhD1DIboe2iEiQ
lRdyQO+xKsfletT3CTY1wXv6/FsZjKZJ7wttTgTTf9x5BCpvRMCJ4PuDaesZg/nX
8U8hRAjw+2qyOjmYMHoJvoE/udHAIVjTy5Ge0nTJmNBo7AWu4II0egsQ3tSH3n0b
jlC+xRQzXk1Q7L/3BQZXuWgrbxPUdAt/HSCCtkcIQZS21DeToDq3Q84z7eIKwgU4
FoQNBoKbehsnCpi+0LKghDvWyBxfJjZ+P98u68eEf6oOvXmQrRt9dzABSNuc7+Je
DFZZ5LcWw82p+tWExevC4E8/uw/wHHWvoVBn3O8PTEYH57eX3bNJY9dsY2oT5S0c
f4vxT+LPbrwAp5e2oBn8XOuabL1RcZz6nnHzMxVpPKYaeHKFDrB2Oz5In/AykE/1
3ua3G/8g+mwwPIL6xXQvVdFCWjSfHnSkWL3Q411EwYuaU0DFKwPwCY37IKIWMHyS
5/y7ipXCECZGg4fZ3QjTzBNXJheaGWG04Wo+qlGv5qjXikdpw6xY19//X+t3gzJj
Id0CVy07oWCaFDa2sj3cxxZpq8LqKlknwaiY0Qob6pILoZGuqQlSsbfw5OWc9/82
x7ql5DoZP7RC+CL5kRplVzOgR06hZdFTk5H5O32zx4pPFdWIGoMDpsOkFBi49c78
JW9s26pM57J0ipmr0E+H/b0iWGFYc56e34DLp85ECiyPt/rfKKmmqYc205ClX+UT
FlpoJ4GlKmaYRcRG7fp1NnQAgpe1cKftmognYV2MoOJuxB7kjJuGOh2dJ26kN/0G
rlL6+4RssygVmANMDy/iMuEMWGmwCFVKdkTjmW92N39JU4Xx9RyhT2/KZ5Vvxyga
145maisSPsxD5sLZNN4Se8PHnn5AFvl9GKdsAkQhMIR3nJzNdg2lH8qxjE5cru/9
8Vz5IsgPpPuMt80xm8VhZNesUfAMdXndY+psOvmSPC7hRaVLkRDdRoDmm2D8iVS2
LCzSfQqHTbUxGSKT3upeWqhQkndud8cdxJvgZYoh9Q4+6vys0T3zR9ug1Iqcp6w9
Mtbz9o1WN94Dxh7M61dvDJkkR8+MLF3KNnvyuzAbA6RbDckIoUkNsCWZV+tJdvcp
lw7wLOzLO0UGfKHKTnh3/hxONQx1Zu8qQ5aT5fQkTMMKTeApPR9wO6e2qepE+kzT
bFkYW079eEKLL8219eM8LVIf2wzMncyu74dmPsfRyNciY4gZ1YLwHkKHZq+YVCkx
rMKWIqrKwwue6nFLp7yGq0wfgpxChwy/WPJ2VatxhtriSlplcgIa+THb8gXyc8m3
Zr56mODEud5u+Gu+BLtHKScnoKQ3ZdYfKXqQMCdJnXeo9+K7Bs9+woeIqAs14opV
/m2QmppzPXk1kUZ6YcxVH3RgNxqafbHC8FS8fGeIymVg/FT9VwkuMrKmFr78dytR
HNGrpFriUv3J00C+ihAAdSn02Vn0j7tE8wth337Tf20hit7A7+VZJwz6wPH2++f5
uN9OdfTrWQxnhkLdyokPRj+D0KCKV6RfUtjEiRkxwkQbW5p+LOY6o45cnWyHzPr/
P38X8GmmqHYnWbPzevDajD7E11qBTvHHyz+qKGqnu3PIYLIP6auG9CnjR91WOL4P
Ji4DWdvu17LyKthDG/EzI7NVx/Fyur75J9SjBLQ6Wvhzmli9HPcrZJYZAHLV0G8g
U3eEx+Lai/FawZ6utF8Gcauugz4W9+InsFQCc+sC0cpkY2M3U4aIzBDB86oC5wSm
nQoWIXJkWPnoYtFd3uAaj3s9OcqJSApNBGn+kobQEouiMGenFPaNq7ysOGV0e3yQ
GOeZikpr4AimGBRJhjIdOghglFpGcSjtkRXUUHS7ah5ti8IMiM2v7+nsh6vzf6sG
PzhYJjHVks2mj5aEkJWy5OuFCqboVe1vm331DVUr5SYM4AwZewhMqbIz9NNGsZnr
qNXicOLzpDN1j0NQJFyudWrx6Gpe2d9kPs0DP4cU/CiBtK4vWCs9gslNvXi26Z8c
s6VTr+qq//Us+wsyyBEKldnQG3pMRJiohCgEldxLqeToUiV1wCe5ZrNGf3nlYmzQ
RA1N46zFB/2Otqj11TVgCePtL/61w5Nf9d3P8O78ISa3lf5be+x7T1/OyBlvIMl8
KAlWamhRhpjAPNr7Q3sHgomtforQJw+DwolK4kpWkClZzLkHmlnIX63FOPXpr2Yo
B5ogLTRdL1Kubchf7VRITnkvRlA/EpQ2piPozE9tygtRWhlL/nvRwGTLE2OO1KTE
tWb2Kw+LnU3bSJAHCtjUR8CEDSGUQvYv31PnS7bxfoHW23RJDX7nkhPtgwXFNl8f
k0D1FwbgxDOSkb2iTFzgF2eJ9dHbwIG/kcq20Qm2VFIn4adChCu4wvaXHR3RXhT/
AUuX03rSjQtwCdpdM/uEt42xMrnoY9r96dw62pXyP0lkxp+xdrrBnZJHZpo6Qqoo
KqFY9Rr+xR+dAkm5ekQCAgYjKxgCPGJUCeql9aKtqja7uAJoD5MldQ71N8ZivlAQ
15/q7Jydhv51t3ldbf3xwYvW27kij1Y4u5qM628p98Xkidi3+oOiu2gkdosa8Thd
RFICvTQJFQVtB0NiFKlxOauKRmn6z2pS3o0rHH5m+QOqPNH78LpwQzfLP4S6Xr0/
Z/+MCSkA9Lj80cCDXBrtdn4Q8jGtaONoADcLZy0ppmcpr9vKWLcjbVdud2uGE4lo
8RruqaDib3wrVqesMehOD/W5if9/0HQTHLxTsRCrJwEf7X4kQjLNr/IIhGzK68OQ
i3Rwbr9JJtNrvcUYD+qYXWW1B+Q3+l2o0Ozkd/Dh0oEenF0WUT/hSSlZnChlKmZE
laYoHHdFB7mAlftzAsg6H2TJIv26Rvy5M161v2jR7Tdly7j3RzecHVmC20jlivHI
0wrB7jUFqpzvR+u8AvlPEgod2kVmmHFoZslClI6wF9NPlxGtI9MTvmaqY4ax7lyb
rVnFld1NFYHMH/6KMYEdMtDKHH2QiQbNuZfO8Wyy2E/MnIZj/p2pnM6/qsCuCjs8
WxZdNSVYTo1a4jrUbMsUmKTc7up2/0gXkV7eZjAWO/mVQYvIUk/OzgLNWL0nHk5u
7sA3avXQR3EUwYhqZvXbh5NgG6dXbiYk8snlPdzJDgyKCi2nebLuq9AHmO880sXZ
QMzQfeSw2cVm+5fHbTHCfBpgsTfcIGtHTZQNFt5WjIuD08MQpe8GTMipmoL8vVkU
6NoHlPcBqsNt+an/uEwvHzFpB5UZUA/qRMoLb90MJTSz3nVj9J5CQqmjXmgd5MFD
dZzEjFV+Zo5U3c9YLDEtBWDgQ0fl/cbPorrlUtZwzTzZMzmN6mSvbTO+Ti2BRDVK
n4OFaiOfT47Fd8x9PrrnvfxpDuBIlBxmqbWbB16ptLw/MWyzOhYVIN+IyU91D6sL
pFqf5phYjyfSIitl5p3BKuUt4ViJdXbNlkYupQd+E/TFUZU7J4RKw3UClD0elYOq
eYFVka9J/HES4oKNwd3IdHfo2dVF6o3uYcsZflXJ+dpt56Xzjn6dWDoS1TBYDjSA
/+vOSWM1S1bE3KZKGEo32RY3g4w1UTP1AF1GhB+Kt7o1jPv4A7/6J7eE3LvKn1YI
3HOxMrF9q5dNEG3GlKg+pL7YZ8l8IYinKk7/acoMiUiu3y2WM0V8Ou9NADU0ewkl
JUIKc8wcuMkC8BlHt/P8Dzx/yf5Xzq/gGURJRQ24cW8sMuBQoTWaMsyvyoNHYyYv
ggADP8Ydii2BScqHs+MX5/5sRi9/00CRM7P15ar7/tKu7WmbQEe4UzQu6TplGd3E
Tr2VmAZe5UQ4dKnXPg8kOSwSgcIb1rfBzqQJ2df+D5Ti6JX9fap1qiGt171F64Uv
MtFyk9BpYnWG4Kp+A9SEuX5IOJg27qQ8V0gS2bfN9wBR+T5D/Hz5SvlH1Ei//76d
pwWYkbqoKqh4w7e8dzO2b3oTRpeiu5TQMFmGEVbsyLa4sdzaFG3Aq+RWDrWx8F4W
dwLjHNmsUH+tH6Uq7Vq7gLLXfXtInGfsKCIWOlhAfAkJN5VgyhtDyxcoMJM6/jd2
XDwPuaPQNrMWlVMX463JGKit62HhCy+rtvrAqSeqhO86EYdT7P1kz/cnCPJkhKfK
8InLzXRVnJdUHzK8lyWicZlLV+pAO53Tww9vuK0OO7ndWweypgCzkHaeW5T1uV7J
HeaXIxj7a+ywhltu+e6GDGbHBp4jMqCnP3kHM8SfXvx99h1bMUOBBgTdNWxmgO4J
XgUwzLxr+ZmmE0o23SgLrBlRTJJY4obrKU8Ngss801B97tGV15WQ4h7QkEcvt7Tc
tkqHJuQV43NiuanLRQwRbmhlmJNcbQLzjbCcXu7a738wKyiidekaeZjyGbU6Uwb+
R0OMudYhwXTdD5gVgBk5rjcgFjTtTAf2MelK2pRrLjShK6+qsIt5Xl//dgi7bQfq
wjYtBxDb1kr1q3c8oYoBNiHb6bdobgINuDP1Ab5PVRMt/zue+PMX0C1FldQZ/V/N
5XFNmBdg41S4cGDK+htHbE36CX5eIHKDDJMwOwLZ8uOnltxzBtbG0ibyrcrlwcye
Ka6hsPRdRUxOoklPQL3PKBFvLJKjsCH2WsmE/13G7Woc4sTb8fcVmylF3SKIamkN
74e1q4RmqxavV2r8bE34wMWXW45GeshM+/A2EnLSSXU1YdmTYCRXyWHMOQz7zdou
GqX29Nh8HyGYe8+gyVXWYdK8026d1XJFQjMG78Xv5QIj77etzkkTYHuozUU7sjJw
26gXS/9cIFstOcl3O6HvO/X6XZyTHCvsGg2qPk6CT6L12M63TLe01WRnCwnkLMGG
JQ0EppD04/+v9EjgTJV7E4LWT7Fu/KQJ9XiezmL92CcsHfeKtgSp7/OXFyTk3K5C
vzmbbFDTWEnpz/aNCEZ8dUxbzTW7G+qSAo126dNTMlGLDUjySvaXZkxqejZfiA9p
FSS/M/z4/hOWyDAig0lPLlgB4LYFTPy2CZVja6hqT2KLE82ncASMKy4qU9oNstdc
G8jhsa2xeG/W2gITxcOO9afTAq5rB3Qw463AIhcIhhhdSoP5NJIW2vRFhLxGLov0
3FG+fsBCQFS9Cu5CxyhtZpz3rPiG0d1o2CerzFWJJzCKq+D7w2UzsZlKbgP3ocdc
ebSnxY2VOz7I6VB28WrM6hOLVSKw/DtO2YmSF+ypE2MtFQAdKC/P4c+AOV159pcG
Bky/bOn3IJt1qgnkzQMq+C631l9nBqLJbfsZvMGVEVCwYr8UC1K7/3qY9uFH+qsJ
aeGtpKAEwt5yMkbrcYM4yhFVhojpZIQTM3QYqBXWeMxWzmlDred97gN2sAmZDU4Q
NMoj56Z2BcFT7IQXZhP1KjnuSlilpup0NHb5EMs6lXYu33OQ/Oc7Qpb8kNZSGUnF
X7WiTw2uKpq5FzDqzdL7KAHcVt4O3PCG0LWouX2/YVD0xSe9SgEHziNTmIi2vw9S
M7qNWLH9K48W6pHj+J797126M1w8FuKCInHSDbtK5Ink2gazoG/WUaiYbf+VELau
aytQYD98YlG9iktf8cv/JsYZ+FubXhm63jDhdB+drqwB9X6dF4fjqwWVUbkEyHzB
D0kiTNzQHV1eMKrCB5SVLg9n1T3GP+Gdu/IqFgUSxC4QgKEXw/q+G9CQWDWVhL+q
nxohrNnZjkAAFqtA4xob18ipk/4s2NeLYgfHqWcJU9vdYy9nrOEWJwxC87VCpUMX
y9AMIW2TwBI5ZkPFlyKSXfej1egtDka4Y2Rzgh5SFvfm3asB1O4UwGwh4K+FU51P
XVtYLGkJp6C7oyONHjNk+u2DoXnDOKxxvxlQGfrp9puEVcSX1UPeLlTFjkm+IndI
swCrC6EYeWV45R94qyLkA3ZPTAH3iwjhxdgoF6mYDwERajQ02eYomk79QaOcu2IP
bd/ukRDOg+a0n6t19o11dfj0i1y+iiQlil91avwr0oyg+XS0KQ2F9TojmHRkQUQM
uZJchecNWJ63OtHeH2sdAg7bGimH5Vg99rujGjKw7p2kp9n6sdOZJg5/xCvMLoNW
NaLC52MJd2BYw97rSA/n3WbW73/oz8J+0PxDYuwyNMzLM3xSseCmvd5dXAO6LyuZ
rdlGSJBopNX/NyC9PTIDKZzvOOTrFTB4fBCybE3YGTFQDiNK3tvO6XuOfyhmC+Iy
FPCdj87xxDUCk+DU9tkE57CCMK5Ex8aYfwVGZP9JljwD0tDEEWZiivDr6QgPg5vw
BqagGCzwqaJVeLJDgQq0FMnw7aszNA0QlN3q8petEnnRmg2GL1sUZmPzOIjY64vb
k0X4LYS1HeCc0bpUpBCIzWWHcZAI6zL9pAp7LSh4IAe7d4tXjFcXigcV7jTVRBaJ
bRIVvzI/7HImZx1PHoVdpMzQOaUo/KeNvUYBIIftZrLAJ267NMBrh2MMlX4zjW5B
PSf04GAMsGAPQ5m+ww4VaRcTpjrw4tODuaRAHZ75bBl+Ozjn/1kOhcM6iS9rCkoy
K6OhZdFAPAheLny3vcXgWZgu+B9sI5LqtPc9nIRbcutoOjGhIGj9gpFwuK1g2bLb
uXS4/LdJJTt7+X3ymPLrzeXZkcKc7YD0y4v0MIhvzXC4Gwn/nrwj/R+Ea0CwvTzX
ROIGU4C0zCrYx+oLY7n1BLdptIrHg8XKtdgEcfOzYXo3a2HowvtwRtHIeV6nYNqq
bgUKiuFwc/vyvwIOuT6K/ICXG762lOf1XRnLcyBttLc/MuI1jcrgrD3dXXNAWrhP
GQtWBrSC111L+YCecIJpfKpXXrLMSfw+pe6gzzbBBCUCIZKbQ7AGtZq02ZDiUtUd
fxsgwya6dR78S0UlZlmnyxd9jzvqYT/btAOl6xlNN+BhP/EUinTux7/cmUhmIEWV
qHqAuhPluMrUjkboD6Or8eaFtJ2IbwXFZlRrD7il0zlVqyHlnZrXuGDTnuZjYGnL
jYjzY+HBUKm9W+D19mK2Vk8hxVWe5PgqelvuF7v1dLgm9BArfeYOibZYVsjiCXrV
Yc6WX7f/esRz/l+tWfQ6KcCzpw6ROZhZdc7o8+teNSBj20ZyKck+coKjmJuCF2/z
JrgkbAhg0rp4bGs7BD25/gXOXuFFLC/31KM9w5wP7PpFNpBvZiyOnaGHI3WnKRpx
jFi30HJ+/LEEoi4WXjINl2tMn9E9MxUB+ioYR0LI53cm1rBPmVuY0RAfyIRuI6mc
3N/XGbIMR9cM4JLSB6SR6sHGfbfoqc+i0EY5ck3pHDSI2nQjlIKDNYSMJrJczo9c
dZkFJDJtLEybKvavo955vViNZpvt0f4AzCK0Jts1YR+o+J6DaldmjhU24tCefF/F
gfzP0N/mrCUsY8klIew4u9OhN6lK44dN4/nYJF3ie+17QUaUg0P6gU94WgBa8RyK
xnI3X1PQaXHdas8s/YpbsNC1zeNB/x97iPTe6xsxbG56TAJ3AMXYni/qMIzUdcp1
JrtSfi1Fi9XWB7ps2iA+VpDrNeTkF04aeUocO3t/Y1k+ht13BzenP8rCk4PBYwjv
LIXFMBV1aaXqnelTXNU83r2MxoGfBtWUQQ5b4rgFpvsCjfv9xtx0RL9tFndjiIBr
AV9/02Qoygca5AkQvBeEMHe4auB8NxGGef0fIBG2aHNgJtpG9NOW7SClnCr/8bHZ
Wp0sSlamdGyknMNIUOkHvn28LdANAebsgVXX2r4sOhWWVh2YcgZ1BWTxrb4lqK3V
/WcwtieFe/aKh0xJsySyZds+Qy+4n5Gr2ZafyJcUYWPkV9CnrKXMNiTCm/uOWUm1
T3qp13Z1UYGcCtp4LRPS3AfeRk0qvAVI7tfevZKJHv9ykro8MjzyKJRWDeDDh7mq
lIWHfS6jIaSLX4cU+tZhgfuuVOqWMhlNGCvao8uuBl4g3Z/tTQnYK0wDxIMdMo3Q
n6dr76n4TzwKBY2U7L2jNyi0oYc2cczYblDsQQFfovcykyDkoqxfWkIlQnzMY7Qc
pAyP3jkZycOoZoivgFHzaNWsp4t/eNT/mVNdoAoIL6YSIod7yiM65hie+XzPlKfB
GxKAWkQ9wY4nNemijX/jhOlNd/tY2fqS4WmhNXLysJPJPmU2rB6nMiJMlsXIFkPc
FNG9Hd4xA50Cd2M+6ydPaOhSZ1stkDbUCd/WsiNZpKR650cGO6+H80X60G5AwzPd
Oj7DYFjK+AuuMKEbOzbFydPBL1OB1BFmDSp70JrNYi9pJkkKsADZ7BAoXKp+jpMG
AzD0HJTWBZnYnzm1fjIN2jahlinGj5Svy4/vP5kgd2A0xgwmaLoRL8V84Xwrug8Q
E8Z9N8jVtulGuSRoe0S4CkEQ7PzqNWM/EZpKBjgqGH/cMmBk4vUzT93da3gK/8i2
Q5eFscxz4aO6Th0VtLHunZQdZ70Pw0NXEBlE/9QCgm9bdWCL1Gw260ptDJitXoZL
ig+SxJb3VatVc3pZo6+u5yUEax8oTtHQfQiqXqq15JwG5u/ftqOb3koqQhoiRFPL
16nGwn2q8hr3M5AgOpE1PFSMeoYCEWQwJgOOtIL1ZLDF0G3f2yNozCGxSIMPaedP
/eYt5F9Tsd/ndzsugV5wh1ULL3vZGWxfXGFN5Ffv/QqLxzVXRaGJeB6ZVFogF9Dz
Ez7BXk/txiSjwLa/8jMG6t6CLTOU/qr7LR9ff/DDDPcuZlY8Y8NjK341lRmI2io8
KdONThla9vWTn+gMOWm2Gs9AfTA7dTEmBhOyNyaWKn/XjdIkMSwkqqAtZm3zjYZk
6kjybi/lTO+Q/BnUBptKbmt7TJToHyLcGcOJ093w5w38g3pY++HV2fSJ0nVegFCN
LvH7GA6DJRknC20DJeQuqY4bW7t9W99pIIbo9yjF2k9XSd83BaDtuIaYSSXcfV84
U+HjewvqK6aHeQmzDSXNFitViWUcnfc5y0yXYNpWF/ByzlsqAqm/qw+qg2NZNSQy
TgqbbRm7VlG65mQSLicPxQSgfsoO3MtYo8sBHGXiKXONVdbvlGxR744+5DHbb+fJ
xYeQI6i8AXPUvB3Hfw2s4inarTeYEHtGxLRUpus4sDU6hBVoa5MsgVMnL5XGeIKA
g412etQJ6XhHr75Md8sCLel74ZIe/fEG1so7Kxo6hfMwNjE1hB+V4hLh2Aak3Yb4
aEC+CR0H+8BXeTCCqB52L0KALU6lx3DUBGfqL96c8oftNfbZNxzr2i2ZUe2ihdw7
jrqGCFaOMYRmD9Klvuujqna547L8OUAIYGriFQwrij4YwDOvQ9LCNoyAgcexcmA9
FICA/ylxdFQjAO1FgLN0vSEKAmDIMexAsuUmDP9N07f7ekXMMBkAEKqws5BpIRlb
HS0fcNyln15J/loPEfeIlAVqjIN/aWSkvqCxNND/CBlZvK9NP8wNRWqAcLgd4MRC
v0NFZZyzS6zol2ZUs9gtRydfQVz+5U10M3X6QetCZE/SzzsUI8Jtczi1HZIT338u
BgLjiRwy2/fkwHiwG2MBchXSxu0ttoHThKXyCWgh5LcRVv0vZJEAO3/6E/otVPJZ
nHetkWhM2pELbt15rmtzcgHAIXRr5EwBAoJkv2+cUr7+RhdCcHgrutGkV4B/i44w
vBCXydZ7h0lF/PXkAfPKE3jxojfRV42hxstftc0oeZ+UsPQ+4ge6rl20nR+vHVOr
cxkK99EwqoohOviOvClQAYFnlw9SypK3RMD9KvAzB4AAc9eklqT6/ATRpDabcYOC
A/C3+qLpJm3TGM1gXvfn1cX3cRDHKf3nWjhHb6c/2fBXyapNMaLOp4L98eDQH/LW
LJhtFQ+rDU4R5NNJg+mB+RiSHJBwmnGRgxLHyhu0KjlCQPyyf1kP2zNhCVp1fIwk
gKmPxTG8bquHi5xnsNl+oCsSFbZQN9jiBxbmZJ8ydOYPzp10EXFIgbt5solqyNYn
vRHyyVTWIPwA54OE11RjVTNwK0JSq6ngsGfEAK46e4y/BwarGFAmvfYEvML2WWcp
/HknwcY7ZIQS8dqLNiIZhZhG5reNuvYisclzq2ci94busOfLmoneip4oDsyVQUx1
RWDL0W9VD+rwF0EnyUFY9a7UAsbf5OOBUEZS/mVy3+JJF4oOr4h13NS9NWhzMkRM
BBwPWcL88ASA8Ynfov3AGMHivFjIh2rJbVOQfkjBj1/3Dk7a4807LT3EpUb/Xc7X
HV2/7swQAbWwyd7nm+2Dpg==
`protect END_PROTECTED
