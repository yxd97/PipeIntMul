`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WhEkbTIA1UuYyPyHO1RcUhju2NsIGXglmXpolVj9mzsEe1l7ixApwsytbjstx1pb
IzrDsPaUEKlhd1dAzsm51HYefijk+X1R5J94hOv5AbnjMsA4GGBKc+6yjiVgl3f1
nioxCxiGWbVZi7n9gtEJI7oMtXMu0kpoS43u+Q3hRJ8MvDHrrLxTRWVUxr12DWHr
R9CKVM7DK4uQSML42HEKOVF3eNxrvzUdE69vpKtaLxs5KtjL6AufcipvrQyzPwPj
VlJ47jMdssGLoYYEUUu58f7U2oZjWbJkphOpzx9Mvn+a9S1nYxG9mVoEtmM3MyRM
bF5jQIYLyorsY3AS4rMP1mD5oPGtQy8hZYjvW3kresLZgQSlIDGSI6cr9qF9LimD
ve0el/Fl1nTMcD/NVSEr82t+6DrfDon6irD0WeGZzXf/pGDXtNDOS6LW24k+6Wkx
VRZqhQ7yxGMNovrr7NbTynGE1tgclEj2RFBCgCdTxR69JCqtHO7COY3W8Lcv09t5
FdP4vCKUUrY2pZUstiBNo0lKtIsoCONF+KvYdDu/RMGw9XtlRNcfJXZhVyPujazG
rlo6UlyyKJwIJvUEJ/NH+KBT6ZhvwnMsbY/fJ3wLrj4cQQXIem/VQUDlFgObrb7J
vnMzsw9MXZoqrugnHj6pW58ns5al19rFXvFvxw0uSSN9oY+MadU/3qRe3LQbyYzo
POtRA1Bv3/UR1EwlbdWsIJaYCOl2kDYWY2b2MckbDBHuNZ1jH0inuGfdL8Ccvu5N
L35eb9ZxIMJR8w5uicUjcGKJKaMd8w9VBc6Yt0DLC2BFovxBsOGDMggRuwAF0npQ
Y2Bbl2ohmkei02xX6EBXLtZVKQebiN5FBfRut2BDCcmCPlE+xTi7/lubvYcV4r0/
vU2dUscJgBM7kprV3z896E2Ij5Ub0gKg7UCvrsRXNEXWq27GrZanCAcAp1lEXXoR
bbnDEZ6evqHk6mih1UxkA+7pqRMiHf5Q/ieDux2phSCq+CJMnEgYxkSzqqDOL862
WBzIsfL/u/HiiWzhnSvuGmub6YECaFZIv2mW3cWHF9wUrsP7dtmcFtsGmFwwGCuC
Z5FA7MvtCpLuqNzziULmjyqnVmJSHdyAcTuNy4Nuz99z8nyugamkF5vLLOkFEASi
sJnfUKVpAA4ktu+w+fE5pWXFXIO+f9blrHykp+H4npohnEm3O9xrKSfryH3XkRff
RdVjrRFFCjNTY1stfgX/ZAE8zHPP9Nu/vhSmjwynJX7xpvnJD7a6qZuws8zPCp3W
vG7v/N8WxPvUzksR3kT+FMoVAa6Xx1KQmfjDwpLG/o/aoIJZJHe2qOsXxrM8jGh+
6y2NRvuyQ/hlGQhav1NruQVU209837axZAKIjJENWXGfP0/FYtc4kI3KqWQ6C3u1
+oIQ96SpxupwQs26VatQL03brsTjt2YsIkN+egkJnRzoP7WP8YkZL08kwo7DXruv
vgjD/Oo9Vh2QyExL1duZU14vnrvhIoDCzDYHpGQdl1kcGydAxEC8fuO1d7lKw98+
Rd93ryGGvowPm/zPr2fieyf28M9VNVW73VoebFCkKkvawBuqdqf1FaQwcbmeUMXO
cb4EyjwwxBnKQvz7T69YTgrJ+FQxRXjLGGSiR3rLJiAkBJyj8RuErwyG0ta76kjI
isJfrncSlyXtz4IY0WPjqP4DZYQo3fLwMXanvF2tOJ997a/3wWAjJOwKpY/25i5W
0uKbU1b3j40OPQFf2bI3zujbYJW5iGyZwAfBRz7P9OQo7s2qnNxxFg4HrzZZsUGA
ql2Z3CSPlw2gkJYr8bnggUostZUtOtGzx1Y4SwG8RTiFn84wQP9tuRPmVZk1U35a
VICOGrk3tYuhk52NDIHqrMvGeFwTrJRTivvAeFjVy4+kbTQ8zGWi7o0im4yG8KiB
iOeoLRVGrRsSAkJFuNEiXveOlP/SqRqtObpPCr7uGedllXO9VhF10bYfF07u2mO4
p7QiEm0ar4AzmkcCzRzMNd+SX2GyJvFl0wryUZrVL3TLKYO1lpiBAMoLYRodr+H9
50qeUEZp7MbwVadWGe+wqi9VSwdZ+7fxrQYNT+ZGJY91e6sCp79Iy15hGddw8xED
6R1LHR6wrEU0jd+iX/4WSmynz1N3IKrDCuSSHNuotWSCjEeKTdH7R7NdMI4osLge
0cQtmj3SJqPUtAoWF7s+OrRG3oIhQxYeWm/zmoqbpDxzqt9KTwPT9Ho79lIKBflt
lW/F4kxIsaMCfy1N+NybeHy8SBx6iaS8tt55MtqjqhMVJtPHSJp3YK6gxXJFjXTh
Xx4RxDv7WQDP/gYCxd1sC4kXVhgvQzW0nUl9ybEaiC6CEDc4ReKgHySlvCAfJFt8
1jwH/aIKXkJNNbA6RGGXx5vgHge9UAzBplmA4nWx5LPJcIh4ZkfwVmvxj+mEpa6s
jmhjLTHMHFpHsoKrlssm/Jnil/CTRk7nRvqvITLbhcJUxR9x2OiakznNuyhqWvPi
eLGKhwqPn+SmwVbc2hyYLt+rYQv5TtWyxG3PNrE6CVrL25PqVTIf9FLhV3LgoKWN
mkqX5dQTm7LzuquF/4h5MMCQKuCGiO1dC/ESRlT+XTVCvmqZTMwZeGq79k1HkfOs
5lhh++anbOzsmMc4gOD1Ur8v2/4KSiEGLcaogcoSMvhaNbSLWZgABysgVRjJnBVQ
RwrzleJPL3JJ4KPUzAC/AokChBmQbgrwkbWdhkKRKI3xTLiY8MODXyHU7cGXitkF
jkEK5d9xAmNw+y2ukpSwUrfOndXU4er+ZOd73FNgqQWkFSg7ppJpSV5U9rajh/ym
0g3pNPAXxXJAXWc5wHzZS6aqk1V1i9hrnhRwrMvjsYHI5b4VoUZ+ALfgthcYipUx
scqktIcGC71ZG3749ioo7E3pohNTAdTGDVNqSk/RXn6/EjPyZU+r03260STrrOSU
ExBeKQ50QWdTOWmeVg5ls/k9s0g1ta0uGa+actsCyZGhMMuhAnInNqxN6ANpyIKE
NLk+97hvab1XrJphQBdi3UoHeVuGmwKp1x9S2pWr994c/IxU1zvZO0ydAA3LDGl9
fdS0mcGaRWDAjfKTPzoXTOIen0qAn60niZ5c94lBOs7K78KxXloUP93wngIQwMXj
hurVEGHKl0ufiCsTbbB7aB1UdqcCpMVp7jwKthLJi8tnDVriaDOv05UMvt5SsuE7
W0aTE6KJTgyC9Om73qzVgdVWjGaDJTdfB9kmmnmKaEE51QxP7a0o4OMRk9RYPzgB
WyCjWXplI7q0UFzJJjg+ElpqPA2+Mfsu/fXp4sXwZRUYoLg5CgITsnv0GoZdA3Zr
1xRb8a2P/vb7uKSfl1iulfIasYEOnZ9ggDseBuhwBCUqD6hvFYaHyh3+0xTzvk24
0BOvr4AU+AQ520Q+SD2RYgm3URSkEM6U0vNzR/tXthGHQgy1MDNpgVUCIJ87IRoS
Cy6xlulRQJwyt+N/9jPX0xOVd3nQSsdCAjQ9b1TujUp06LOXHafePx5+mKntzqGC
9ozIvuW3/XvhLMv3TZ8OoooRIV274zfhandzduiBR1i6wk00DFaGagD5o6EksagL
i+TVkZjqDEsgTtZ07EAmaG6VZi33hblkKbXmk2J7Zyng4KRvhbT01xe3cyR+5Kc3
8pyPn87mPj3xl+Weima4SUjJhYtIGFLkRp3XvyjTay67sLpbSZrVxyiHrFhLk/i5
8xW5Yg3KjdZuvD/x4wi0WeW48I849VbKonDJ6jbT0j9XZF8mAUNvZdtgG4/2VeJK
YH45ck+FHAH8+TV2GIsT/Z7AwYtnNx/l/A7nTHe7cU/wj9Z8rYhcQpNtXWbl6wjO
MnegnWbpvPoK6ZQU+Qi1YVoE8d4cVtIbRyR41CibqzToMq0l7obhBK2a5x0q3OzR
ss6a6wRKPwWBl2rFKOixGs6OKzg6KsFOPuFWgc7dEdA=
`protect END_PROTECTED
