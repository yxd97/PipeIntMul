`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HWUyRlQA0NqDVzBpwl889RtuklO0Tz3LM1Zd9mNtFWHbSzqX+NFZu63rYeFm126x
E4Dzn9I5YrMF1WrF/65yS4Flq5+GLIgYVRkWEgEwIXQOZ1STMiaBXy7v7X1/8kSV
X7ei+3Ah/oOhAtOZtICZUgmRSbs/oWLtFA4I/7tp23PwKHFQ/pqt90MjTPHE7UAM
Sv0THatNgN7+NtB2p/s5Yt9dHZGzKZrn+Q/PgA9fbNUBBiXFi/bC6K6ylnD2nGd4
nXSbLzeJwjP8gjf4hvUfi6/38nqv31OU8FtT/+JL9YHZTXAlW9Tq9X7tjVgZJ/Pc
f0Klm0YzGypA6rNqHVs5x//MhuEJxPf6PFoum3Aax5liQ/GmXYR7wGzhgJuFKH3Q
`protect END_PROTECTED
