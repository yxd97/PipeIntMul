`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FWZwVXA1YEIt/aVJvs3aytAq+O5D7kbSJ2YeFgNu2bbpBRwL+aoUBdp0cPMmkSeT
955+EuRCTXRBZFs4yzx4JtJVaSXf5ZQmbTQITTTgWbIqJ4hfGmk0ksYY2E2zzlNh
q2aezqgFFBptYQOvMvF5jHRVeLuGA1zc9cNMKuv3T8w6Fk2IfCTNOY3ADm8QlX9m
q2MkQdy+tmIYj9yk00T92aeQNgaiwncLyuva7MaZZx/tZzrNmO2CwoQf93W8D1Nt
S9PBVWblEiNFUeoTzO0OB+Qhyqr/7XayFtIob9iqOA2stxeF+/+bunZNdmjUbgNQ
qTsyK4LfQytc04qmYUwz+jZaqWl5ONwkSZ1WLEINyX9rjuAt8nBQWpwSaNmPLFFS
0bNb00NPfPfV6sP/92kafOhbxIPdA6wGqyuReBRQz9x9cQlVjBjQHpDWmbKV+f3z
jBbwhp+y4n86qhcAED98BJv4wJacBUDrQ0S7IvEO0EXZ+Xksyfc4c85A341BIJ1+
2hC0nzZbNWYMdogGccaw+ZlJ8IalgM9fw3qeF1+juKOzMFHplV6kYEBVrK/UfMPO
vm4q4/23x3HlgDOzZ9lUZBacuXj50lnd+FlNNwWmcA9dfoe6uUh39DWClvADIRcU
34QNKgB2yVCTs4cF3XAx+0uDXcLT73f4K57B6CwOL/uhBk7hDb1byz3/SDxry7pN
aPI3QjEgs0hcWyNiSixK9ayC05kLTTS4xy3bUTfCLfvswLAryyjVGfloiSzZk220
bKd7WsnYL9zaXZqv30GnmgF/hDL4vgpa/R3UisLzwkRpnDMrdLzezQpgcwthBWJv
`protect END_PROTECTED
