`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fXHPy2Oz5joEkv3BPzweoeTX10NKNHcM+MJrESqbkE9iQUIIBt9Uay8s3IUv6XA
pQZwj0gmsDBw4oJsnToSTkzBDER9We7PRD3l5c9ZSEux1qWSbD4kkQhB7RodKRzl
tbuyLXBHRAH1LamavkzG7Cg8xK9HMRJ9B3euHE5JR0wtwK/0OW7jgaolXi7Jbt55
APjWO+R9us5p57u6DNU/sWcV14TFJ0mLS2EqGfGWkvmcEHRCLoklsQX+afwdpdxQ
NE8WDHL1QRBgGMMpSkrPwyLVCuT1dapi5qfbnhBOvOig65w02PxGBgwjdfOl/zkS
LQtrqYay3eEVl/igKQO5DvPT8ACUDAgxWo+tyJTK/lMqL45JzJsPGwg1CuCvhZ47
cq7voaNcJy45o3Fx3IXPW4Pkka4hMrLmbaDCWltw4WinW0ka2M7piiiKRw/EHON2
y+6tTjLncqEmBXuQ+wvoDYm87MnJgy/WEX9yQHIJB8WVia4fNXi7yvCRxZivLGEN
L2F74qbzl/GAbEnLXxvKPFFcwePdg+YHgmotQW2fPP/RSRIrBR7friJ8EJ0NQz17
xNxfWWrEB2Hzp8AWM8P9WE8OmNn7xhZmQR3BfZvvuszQzGXjErUorcCnwGl0XCbq
zAZ1RqS5teSVdwutnSoeLY1gxslVyBUmHsU3w7+bUR6qw53A1jpbiOG/7O4TA+5s
rjP6n0r9RiQ5p4VMPJB/zStKNs+yT4h9nsiqgdn2+X95aObIPbQsq89qK6MLtFii
cNGRTdcX1LGZ4XcLNnIxrp9sUR6C503XGtqbJlcB0+u6UQQfF1ZQMfZWCuBfSm3U
21IMjQYJ/4hdQcGLfYmgkDBaFVJQrDpF/0R6JqjI2QW/0GAF0FMRwrdsb7e2Lmft
sSkgkn27JnfOsUHajxFv3i4kU7AMFbxtQQczC+4c+NegY65if1mYCROBFHUdFqwX
82HF7izfBRI8odqvvJH0mX0W4IKSeuQWKSxKzeYGdv+EpX0T6vpdUHz6Klc3qNmk
goaWEi2KmoviAsFQ7VDbe2d9nX9jVDWO5xX+qeO3ORc7mgjO4l3geUH7QSq6x7GT
8lIw2/MPQ0K0JOVpZEBL8KPFKeP31PY3Bd9SnM/tJp+daZLzoYPLZFh6in16S/EY
OTt776NfARpHIu/XLD/mbUcPQaN8xZcwI+S8ksvcAQRNrle9oRPNyW12gneDcl8+
b9Dft3+prY0YipgUbsS5ri3KgE2YneX9IcEaXj/lZim74aQHgz7l9be59sh25zBL
0hI7/MrkBoRJ4sjJ/p5q8qQUyo/0gymyZe3eoKy2/59YZorE2jZcI+F9/jOOd2bo
d43sOW2G0OUAWvnnI6z/5J8L7T3vRW7KIzqbsS8H9oF7SMitnj1c1eHEzUvXvwU7
+29dtSpf+3qeaCv9Jiwrx1ak9+gt9x5em7dGuE7/Us1a20rqYbiYVNbSQZwUI2W0
jOEksrItSlB+qyEymCQHFgT4uAurSnMJZS0b3NoXgr/IxEFBjhUQOdPMk5LSyi9O
gDINEhR/Jfyk1ve5I21GV/zpwQm53PcGW6Mlm8Wxx8NML1hp5MPNv6euVUXW5qAJ
jpO+lUVSm6f2U/kgHhDxPOPV6SfRVanwvrw6qp2NIqfIAi32ui4/1+sUF3LD+lOP
qMB9eYv1mbyCgMO7CU7UeAn/sU9R8/hEYh0hcN9+Bl9iB7kKEK46/6UqiuS+RykZ
qg3YdYkBBx+JF7cfFXkh4bE7+QlskwouPQlfMgf9TZinMhJHnzxG8qZuXMJSWmlf
QymHv/ibvrHykypQG19j8hWzXgNz2M4y3+DXDEUM+T+2D9KFeU2NiDf/73wtKPUf
qEjX1noCtncpvx7I9s/izf/nMEOuabNF4JqQHoJ6L7aYILtniDwJKPEa6Gmw9ifa
KrEHUaHSSEX37yC8WkKuHvbCYu9K6IHazzaoZ38zIaPCpdwE+uLNw5ilknkX5vL1
YREAOFlmbwDUppp6qmc7kTPFsvboAOAUHox0R5el3kFUQoh+tqVXfxFhP0jGJ69D
zKNzIlEleMV79STWUpg63oO/PxesMEM/HHamyuerA2xDlXEo4mtPgUi6BWnbsqaM
KcSU9vy3scjdp1JOHxv4ummaE0sJsowaCK9D7aZ2wL9KA7x/vLD2TeLOawlSbI4g
s0IshKMz76wd70tGs25yCdleVakFzTxyDKJ0vQGiIMQqb4uwxyoSY0pxtccA1k41
0mGHtE/yX982kTuSeOeJqGhlClZiHkTzTz+w52bitacVtzU2+1C7qFFlUMK+UBQZ
ToRYhuLdj2GPRK5a2jelYgzJqTdxr1zXs4Re4LGQZRvh2lGU2fPXs07nmRlsOcS7
aWpzHmnlZrDkgAbS2QBIvR4JBrpVsBKEo7LzQQgJnsqUMWrEyp4sBZgoZq2oyWqc
DuUJnc0viLvfS5hkpG8DRHZcqCBa41ps0UkJvGgVCMqLRUtqWK/5LQkAxGDboHvJ
bcYJXUOzM9Uy6+pwQsR4NWWjqtJqZ1jVdN7VYrTpE5RFtSE9UEd9BYbBF6bUhfK+
U9NmAmZFthVk2XUnRJHwNAIJlqXL8E9IJqTpq7JWsle9PTJbhcknvc3SWOAv0v6K
9xyG5q3MklBJh7vHWoF8qwAhxK3S8VCZxXZLl/9egmB1ywtfyoWnOJfLvHwHJyAS
amYUIPCgdUFp9zGGf9L+y5i6MTrnQuC0WLvR9UbCyyiClPUwm5MQwd66z3cbt5O8
3Fz4Vkvg4dZ1ITH7WrTWE5QL7tx7WX1NLIx5z8jzDjGLyxpjlt2JdNI7tCv0FFEG
nX3SHEC1RD3SKKPID633evlcdht6rvk9jXXT8MGmokAWqd8Lghp/M6cBwF+NCrI3
aCp1deG6CgVG3hcC4C+P1JGRIwvSaO/Axem8giwyaZKabTS9S580c3kZ+t1L9382
a1do200L0yqlTtofR9dMOsYr6Erq2dg3ahSVUmOkq5Xc48u7eONrPgwwzoP0lYRT
7pIVHBp9gNlrsroJb/ugDVxtSjMOEK8yx5dbZdVwadmUd+lKQfdsyNyJZwpO2mI/
koeP2DMjYxls223IwvRGpBoCL3IClo8k0JyjmrLiG9VuCj2UZ+632SVeriT5PDtW
D/ch/8zHB8mrg3kBYcv78VruYsRNtt6I+qIredpTzMTErqm9RS3gIbT0e6e1Ffnb
qbWFTxoqWMN55sR95fnZH1teMB5nSoccyhQSxqpr4IqcOQ54T1gMKkRNrm10Btq8
K7/fQ/hVAu7bpm+3QewiGUsCw86G+BkAxOj4x6CA9l+7tsq/s9xYsTaxkeHf03/U
RML3g9+qmZ0BPLuH0TgjsMyKdNPuNk/RaeZ9qNQYe9ygmaOhYalsh4h+wU3tXyc6
nhzxyL7csG8cabq5u5OIy7hpWE9eRTPOCE6YJA1YjqG0R8OrKvrpzODnT/ktAXsW
TWZQ3SKuJ3iZfH3Wul2tAzeoPv2ADCl3vDeQf5NzJbZtUVh10LarATQc2e2DGoUp
bOLkHeW2C53TRGQbUe1/Fcyz8M9M5Ts9jmETXv+YQ7SWM6c1PdFS2MBB0mnOuNQv
LqmE6my42ki2Q3VsZL0zAyowRa9FqcuSUTeCqaa2/IU0aXliZScIjYdZFso3gq6T
t3SpPOnNR+IyDKtZ3H23U2VepSxB4suhTe6HW7VhAjX7N7DVHpuT01Dee3wvPbBk
TFzjNMXGdcWxrPNyZ1RZQAeYkza16x13KK+L9BoEI8D5ya/dFxXa6Ah6EdsnJ983
6BUDifjmz93F6wPPXfkBwdnxRc7iMGZuuWfLJpZu1GYxVBVU8SvEfS7fAVKgoebZ
FFF7dFzlDgiP1jRwl1LsPhUveO9AXD1kSSTOZsA4HXxpJa0BCOSJvkpoe1dIv2Pf
O3brApNnyuQ+d9C8GlkpM7LpbbKMlNCKqXDIPco3kXaWRUxF0FKz/hX8JCJqtQQt
Oij6ORbFbP6Xpxp/BGySoEk85AI17lSDgeaYwdX9B8LXSQOCOyz5xIguWKM3L8vn
ndNplAV8f9uy+zEiexM+Tc1hIYemwaCB+GYZR0062ifUNM2SzoiiikS4sLAuS25J
Lk6javNS6pxvHqLr+BnyhFJT5M7PSUkKHoUlRR5Hi1mKhkroM34JAniQcGsBJyCr
ZuwxrMIMJRnswUTLrMw/mMU3wwJ2JA+UENk22TCklO2AK7wO+p9oCiyCHJRpdDDb
JEdkW0ihu3kWuimeXZHaT60e+rg3Vg3d2RQaVlBhumcJkIBncGuwdlm706fKv4OK
Gw3WgoZfQNGRmsXMLxAHJbQ6iKr9h+hBgJC1zzSWHONYnThNIEqB7h1lTJ4kwmaE
FHNo+RBl0a9Unr0+/XXMsj94o3FK/r8Rjj/9H6yYfnQw3NmfWNbqWTvljVgtEQTB
p4EEdRZOLMGn+ijLiBrpqdonA4bO3zwxxpYNUW14r5iLIvJiilDHIVV3BacM18yb
fdoQoOfaSGraKw0KJCfHhR6kigrvP0xvOJeK8AsBS+BbtdCqwCCTCi44NBJwMl2d
FKwI+1afGKOzYqZcw7wm4T82ghXW7glKSPsPIMMVYozN5t7M5LQ8Apm++T5d4l81
0N/LXlDgdZFmxZax3NVKwnTb/Br4kVLtby3dpINviVP5FKyoWLhqxDoP32rWiszM
UGz3BLabFc3KqzcLAK48XY6oDagKNB5zcYm6MkY6UgwQxb2ohHFDgLDOEO0CWXCI
Ihd89M3x0jEdlkNuk6vh/tpIFkYKqHNkh34YF8QlHmybp9+wnIkUuAguIQmT80G7
DmDb295sW7P+Tugm19JXgyqRf12qFDjUYCQKIk6M61WlvB/jLSAF+pE/+Zz4nQmH
NVwlVKtGphLjSNgB+XbW42ZtQbIHxPPUTxaf6GMrBdqS3I11twQC8yoPzEAcCKop
AHcGWSDJcp/XcK8tUIKIORE+KIePTFmCg8UuCPm9CtAvZxd1TPWKWqmnW+Jtnw4q
XyYgXtvldN0h+gFaGOqTIbnvRzN9sc249eJOfPWAFchZPBcnLXN+RpaIkOGDpfr5
hEZsGqza8Pr70K6tGITGMehFzXIkxIaYwolZZKwbH7PdABO7Z/xPdHlf9tntqRuY
xuD58r33Hcx6r7VBmHo2ugxhIZg10nQ418Ohlko2LqkUGkx9W6TSZ6P+xmBHwgEr
buCx4SpVlEIIKKnMyxCSNqdLTyPpfgg3Vg0JIFggpJnG8TD2hFtAxnDx4rEXXjJX
zt99HU0/tryuT2o2b0kiMHRRRTHo8qwCddcCwD77krCQfM4HtPPlHIVNiKgYouoR
bMUdlZvwAMbyaJI0PYVq84RiQwlW2jMiZo370zLB6LLj7vdZpuXzCWb/CE0XUWQu
cdJt62mspe5PMRnAkYmWam+feN2Yrxvcfrmz9vCM5cP8GJsbcHGsIuzOENiYR405
CNqkT7WFh3v6/EoriMzXnxm9so1RKTE5XzxccEonyHfpb9J7cV8m8AefmNOGW6Jh
EkFTsxPdWwteTul1pdguCpkOiHH+dpEAROOIhf0mzb83yNixu5MfiuTyuNG2lthO
YvHRUPMoAP8GSGz9v3TticQVM3wOsdp7spzPLsY/91C+c+4/ld9b3qxINDDDk2YS
yrZ7Ico24rKE5F0V4vaMVnRkMh3N4SxCldh0b6f3qJ2uLdfBC9oAfx3c6qOUrYbX
kLsQ5+83VQoWAYg+83tvD6PAzpZlp+RkwY1CdGrX4fQ6F8sBjfjA8wdW1lDvtbE2
ia/mQgAAaoNNrZyVl9hCGl14f2kDyubnLrFlffQPSadKgFYlPc9TaerQI0QR5L2j
hOCFKsAtzuwLYwIEFcKC7D9qS4jOHfecLG9GnANv2gxNE5tAiVpWvtzErnj2pHUU
XJH5ktErCaQAxn6Z0gXFH07oEnUBh9zkqG+DW583LNZR+rv6qX7pv6P4RWIL6HVE
jcyw03oOGB9qQ3SswoOopDifAb22ss6c5lobD4Xgt+V3EYe3hb/dW/1yPJ44YJx1
RwCVe4xXajFKpNo59IJqRIippraID0oHHLMLKSRFrHKUTeYBBZJjwv4F6V8Ck7zg
4pxtAdc2KW8NruUfkMF8gbq7/aU1xeXV6vx8gIPsm5Mjlq0dc/jSjH0KR4944ZTM
SyAOcJrJNooUlZyulg5j8KHAlWAw7OVljbagBXHkW/1+9cu5cLsurmCKl8GBgVJ0
BSNF/lWgy/tGLq/T6fKfU7z5lQki4oEnpmn343Q147Xus4GX2wbRAIzwKGfcNAAJ
u+57TgHmj2v2A60M0V4kphIqnJKvvzMG43yt2NZW9ukCmI+XzOyIJz6qq1ydk991
cUnPcdhkcPu63eiUDzo5FwQsHnJp2AfQBGLDYfX/B85DSU1ZwVYt6tL4lGU2c36U
NjsnE6EJzU8xl+oabbvii5oFrADlPsDx/ltO4aBlCxMIyj4/8GbhKxaA2Ud8soBC
pnHDAfQyfXMHf402TXo/nJvLVz5wHhDuVOqrzA/2oJDXveJC/83LZHJv5X6tJMft
2sEZq3pk+BWRlrVewG8ZmFkd0vzSnGI4nzcTBWkJwzGPZe81ntZNBpc3l9mXrQJn
FtxKDfppS3LksqXO6pZIWeooTHthExv8jL/+BvZBbyLbnwDhFnqZBfvvPfmYTdzg
GhAZ/eN/bondC0AHjsSzXB0ns5omUkE5uz55Mm9uCZteXXTfY4zSuMmDdDoowXoO
RTeXCznztSf76bPlk/1m3Gu5JaDmquT3xFXq80V+2/MxiGmVepceIZsTKQDdzlle
laazwc/hml+qCLR6bQfbvJj8Wa73Hu6Op+N8F9f2qh6hepPg/EZe6eXfJswt9O1L
t7DGYe850ffOn77QvjbTTQwQNNHGHizn8zed2tZAVQeSt8AHXfgm7eLsEgPJIAvr
WjXylL8vSHK3rRo+NcnBR4w84Eic5tvn/LmMEW3OO7vXuhnBn4nQPQFUg05ahMCw
zGOXUoGPBt61veLaI7PgbQv9A9GRpjhXB3zqE5h3sqDoEG9NKnm7fc0FcoJQkjmL
v0nutjxEciT7+eekloGiyXZUeq6psFCV1FL1b+dqheBSX+k8KBdutkjxggcF3qM3
hD/on5Iqq3QmMnm00vLBWW3O/HZVi16ydi9g1cqKoW79krTnsK1PEbETtJvff7NA
9QovIrjqCR16bhrcIVkwylG14jLQLvlezugZw1ReqJlus8xHKid/xfMfNbn8F3FT
RAzxmUIBnJQXj6tPw7th8Gh0cpBkVPoFZPEiWztFe1soeBGWKO3GeWup2hCmoV9j
vgdqT7fhYEpNw4uXYW/S8FvivDlw9DE0eFolscjeaf4jAGhwCFOJIpt9QDRW6//8
6SlCrBz+mVw57yd7YkdDDX7MR0qCc7jppQRRXiNm0zLR45Npm8kUZf44C+cZuuoY
nTIiwGL4Ee0kJ01Em7GwC/KFijU0G4S/ZesY4CY+IlZI9YiHqGCIYcJPrW9+iwa8
VQ5A4EAovfgnja/hGy+ZSkrmX6msweIbrRmD5IBJCj0YlE1yhMitTV9UhR/rDaEQ
2lZoj3NtUr3fvWuLMI81j1Ofpw33WwepHaehtZVxg3bfT3YYezELhIQiH2Vb/7uR
kN56G5WsoxVBdRYMen7BP9ovdnJWN4+STs3Fi71InQTuuoTUPJLwXQcG/t7PGgWf
huiuT75la8O2dK79lHmNy+jw6QeGmoQhWe01w07oNzKalNIogmQnzPhkmWpQ9nN5
17EADNCejkwlKfHEkQvl1GfKmfYNojFkazuSO/TZDS/1u+UWKfyZq/1HpVH4p6ZP
wkRimIXmyjp2Cf8BPQJjL+f3mXYE1ZiayKf43AUJEazT75xHIeTJE4oMhCBr+bQ8
W2pR6kkAlC03IHndu/uUwZKE2+txRxkEwM6Xa37O7Y9mfskifsEbuquGVsTnAdr1
sF9KoLsURfXBVxQUjnFHs3bsyYq6/WqWj+GmPCIr2yEBmQOxwKlsLT1HD5/UBqnQ
KUBZnE4clMBcnJUyBLq8mrfbja6/wHj9Npf/SwaMjnbM38v47iHuwsDcGMROak20
0GlDL5gP6yH81lGXIpe0ivNuUWcw//MLXt7HeJMBXVKIxVmxz5z/Le52voYGqMzg
so9bA5kCGVm4kKrFLvxMGbDjgBmHjefNgRAVN6WZM2rf0h/OHLkPaXP8zEY7fTKH
DBnwBPSKI0buLPn8pKX8HaocadJ+tzVQ/6ySjosZeSDOkZtp6ytp/88dM7Li9OjI
EMLcSqbkJ/5+M5obXE0Luk8BJmy0OE5N7LQVZoAdjg1vKRY/Gz9icfHJiDyug328
XFps2IQqEzplYCXg2ODwb1ICmPhpETL6NB8Aye4e1t2rCI8lJcEzg8w4QrVZy2xi
6yA0mIHDlhGbRlZzUclnKcDnR9sP3E7RyGa4yawOlBLSSJ35NQC+cC0RmCJLamMn
o3ACgx/ELWc8+X9dGTDPYXtplAZu30sUP1cterpMzkK2qURH/De+wBKjzSiFafBC
8w9oUMKUAfVtY/VhZtqpXd1h/ao/BmnAf8hpi/8Q6sH9xHN/bZxHWb5PPRohcFYf
aCaWM8wIojR811T4hXwiLhZEvBYRR+MxdbS+KtWJF4FAVZI4EO0epLEW/zCK+/b3
vP+Q8F5onXpxlUq5pQr5tm2wn/vj7JMXF7L6dO+ghfwiWsu1MCHspw/Y6EJsc6Ig
yVKC3BTCui4RXUdfszNeqKT4RipxDU5UHwGOYv7rgUTzhzuf360Wdh9XA8oRSHqu
zt5lXPr6p6guj/IRgIGnmKINTKBf5ktes2GauM8XnoIBaKZNlWGw+DH1AzrmIDsc
v06z2Qu+lGBAl5maE5yfEe7JSVJT+64LQFYRsQx0R9gVBlG5hWjPER3PpCnY4/RF
aaI/a/6FoIHcbdammR3n0AVtxeDTKfozgvBeEb7nQGPnCV4RuGm3h+mHXXoXcOPZ
jUK7raRSewCWesj5YPVmEG1gvYSrk0BPRXAH72yL1gVMJUr9PS+rbCWg/zUGVB68
zKX3a0vT8fnGjdCBeWpCg4+/sH2ZeRzta9JXFGdDBvLMtQxA0WEO26/4Gh6GLfLE
O6j9ssnQ3PMuYi2Q6PHrpuLQivwJSwQNfOA+sy39wPO285cUOcSiE6/QQU3t2fvN
ARU/Fipd9iBzXaJsnEoM0GLIwpGuFDUlWQPs62hydtAytYaramtSZLjbrTfobeHY
qWsXO/LZtzonfT0yDViM2WG6oZ+Di4s7FxWEFQ26iUcsqXjT2+7KOOWvnkB9i2uL
tPImCzNyYkLr5ymOfUY13cjyQyRyL4hmBIWfF6cBJ/+xrwpCBGRvkzpuAwUKCBc6
hzMUn3vfP/mn0iQwx4cYTg==
`protect END_PROTECTED
