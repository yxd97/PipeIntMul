`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h1ZfHFzxjjwIXHYd7YszpC6bDHrClmxiKUYCSe40RvvRzRr/++0/MeixW9Cmprqc
OdGVffJv0ASHF3Vq8Xo+263jatyfKieNnsi8bp168D0B1xKLLjDtYhMrTk4h0Qw+
OB9PDc8I6OMggIF3Bhh6Uv39ZqaoH6BcTSnuxzFmhataJvCJWCvU8BW+1d2q7SAX
YHP82cCfI0C6gDklrlXdvvKOHEOY5XJGOOuW3VnqfI2sX3dUgMMy4iHOR7TXb1K1
w1d9QorLmneFgX0YodnXxEhL34C/BDLCEVb+MicJwAm8W1VCeSCS5A7HJfUmsbkX
k7I8tjzocDDJhO3i7yDaMcCISK/8J6Zl45VJU8l99hL1xmQt51gEvHodAP6V1J+p
dp6LAMrwqiBgkemXoRjLyJlE93VAiK2M5ZOvJVrnn0jJlrVH1M61DO3Z+mdvkTLV
5rTyJ3cDc2sFSnxJjsDsVan7RtgR2aWvJIZTIxiuCvZ2Bi+NIs85GnNPfkNc2/qN
Q6kDT4ZY5FsHqv8FJuANzUxOFxbzbfLhF8vsulAIq747QlFq41xdm3w2PUEKA3EQ
0gu0+6IYNCTq6FqyvCrgPGUAh2vguavAwCjlOF0L6bl9Zw3zn8+B293pFjouSPSi
M4ag2Wp9xwOXAQYb8r5kD0+OoChs13T77uGtE5WVEY0=
`protect END_PROTECTED
