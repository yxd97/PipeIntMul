`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLxuwmUbTNFpXsX7DJ4n4L82EVJs9SneZX0bTdDL94haW5W6WFGNzjupPX21t1+1
W3XAShr7IqdPH+dI8fUQ/pv6/5eGRGU/TMyzNMhW7iWiOkOPL62cMCGUv8ghM2RE
NJQgLV+P+YdqDbGYD7hbki4M/9hw72qf8+bro5tIu61I4a+gYhGEp/x2QvNkuv9Q
OO+CXcXXrvJ9UH/IoccochTV8iHxoR7TZg36Z01Y4j6HrWQhA7eFpXrxioOocdzj
0YbA6BDXE4eHKH+ruuwW8s0L+8skwNuvFf1aXI3QJWuXzITnUAaj08jUCk5d8qtZ
cM004kG4aLFCJP2e1nHtguw+01E60k8JIz5mRwXcSJw4pjYJ3nWL/j48oUWjWSac
bqlm+qxjY7rc4UQFwxO+nimzafeEzGQq6bt9bFrQ1Z6y+y6lxfIgQXFaiyPgj/fv
+c2oleKP65n9ZxDGaq0UwV/as26t71nhpvt0xGlZmyRtfrtyApoA3fDKqNfMxJTJ
3uv5DAhg+o0Dx4RRLEA6xJVnJ41HQyP2CjiGtDFKUNoxFtGkcV/BxHQEmqFxaMQ9
bm2ulhgS/mAENqV/wQbaaJzDxBiLT3xKww8ndgtG9mSP09DfBMEKphZCRWqUnsYV
+21btVXjEq3UQaA7x3mJzSwZshrARL1zNKmUKT21dZBnIB5MdTKKrJ7leWDfuNXS
rvMHfw/7RfQgABRHcHmmehwA10OaUlUmT+yiVHBMSr9lggdAXjHfnXyg15kykKRx
5JjFwBOh73IDIty754LTRhQGp+KWZUKYDbkGeVW4srQZK4nwhn0M0Q76eZFcWjZE
mNiJViTLLpwzgvB8Yez4k52xLNZd0LZv/rMbkBfglPALZb74F3+BMM6FD8Pgdwqd
/rRop814YnsMxEiJNhxLc6sAZNHWmkbSF9tz9mwjGrKMI0ewgWNZo7lpI6paP9ih
N3lnzUt/mvW3ubZuQSPeFWkrZpYCxfERATkf4S+uIYgXjrnF9/Rn5GmeT+3TQDAC
i7N+x6a+z4fzE0f5bmgVBorr7lXqwgH2GGRfkLR8q8h0wEbSOV/Z1MxQpxwdF8z8
TPEO6xVxP86nLHQXXU9aSXw5n3l6XdgAxwP7r4DmUIo6Tzm4hAtDmcV64ijpTbjf
0KaPmvlvbS7W4eQzWfoQ5QNB/a3vB0nhjZepXuETzAeYm1iYTN7sdTDYz0thh3l3
g21g4CVDtuiZaBUuEs1x+iMZ6ourFkdfuEvIpmMMzv3agNoeOuwAfxw10c3QYW9b
ub6Z5g8flwsWaCl+HbkiVsA/1mJ818MhK+DiU5IM9y38ue3NHo79v0hLrC6MBltT
L8GgCC/dheUlTyVbDgvSmzWEKHlohYsRluxz3i/o281PUjch+syC7DN5Tc7lY7Tp
G2A6cWFCQ0Fh8ouicaEnXpG2HMmqm9+upQGRhbf1sUb7rZ/S20Wi3IFAhr4Jri0r
7pEKK5cVYJS6r4icQijs7juZTU7P7B1JZ5H9gb7zQuLVl8vgca1oE07DLU8SnSOP
UHHIlMpgSv1YkmEMt8JGcV/DakGmUuTSHZ88SKMfzXWTtsYwyGDpMX+5oRMtPobU
WTkT5xxski6ktPh8cKIB6y3NEP7EeafVhMYKnEZaLYMl9GgVOi2PRliqLhUdE06q
N7GiSMjIZxbWRd9LgZd6HhCmRAsYwI06PzNg203rX29sXZbklOn7XxEud8oR0JEt
96VLuOEMhHUhQ27MLCUCnVd1CvLK0xJMoCUt8+6s7MSieEJhQYOh4/TLYdsKhx0i
LKF7xgvqpeJAAfzlUGaPZllx/1LJvIQUZdQbclCW+DHMfNQZD9I3X6A890n49M/j
1di399jjqms2+WfhfWf2uzPsdHqDXWlfS13GUyvMElj0cL6B79YkYDFpAsl6kiLq
TjoY8OlNKi1cHj6A46wbaaulmRcRPSg2V959zgYDPMiGyB8I5nVT0djX4e6eD1FG
nAglrT9PxgZG17DiOnuvsbvCFXitz6dMzGjHqv+gHiWM+fV+5gDRRBkyKSaKJyTg
x2pgegR5yuauvE0i5vxlQJwmltVbTmq7QOD97kQrrNcyEQWwHUpWUnH5+b8u3oRi
tM+U1ebQsrk+4GavlQbpqUQdfO09lANqTnU4dXYIQ4OEgcDH9RM3VVRIYLJUDFCQ
65u4+G79WYjiFFIC/3zLyvKBXSh4s8bRQ0UVUhAdARFXMeteIdBsmQVBHva5bi9Y
vWwDxZEgEV9D/zouHtdAvki5UfX/0XZtbgw6Pdf915gqkBnoIjbf5N1AEXCc09Lx
JDG0ArpDf4uwxX1ENe0EYzVte97lmWAyXDZ1tMAwMe2GInw0wXvtJgm/OI29tIhb
KzLfwFcNHVO8IK6vyfDmtDP036hBHl+r2RkIFfwWZMJeFuIymFsJ9QfcUFuwfBjg
39nK1y33+b4axpePHyVWl/VMRspl7sVxO5+ThPzI7iGU+uQovD8exL3eP5EdSmam
+n/YoPn78vs4xREfSTkWo3wW+fafXnikRbq3HdNJhwOOXiuyMRim9DHm5fEFR/DJ
8sE40Pi/b7hx84PHrmi43fhaOroMxbUliUQGHqMv8Ma2oQ2AXc8enuBV8FN2V9ha
67tLeic7bpbaV+cA5QihSI1vWb5ERaz2h4BlB844IS0OLFZS14xOesbCcM/BwK8h
`protect END_PROTECTED
