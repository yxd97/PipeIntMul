`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HjJ1KSacJBGweYcxyyR0AvrydSD+XYJiRQTWoZA/IgR7EKMydP820kdukN7EhMq
ikNf47kBoaKY7noyUtMqykrG/HM07xYxlJz5BSQKAshmGbZgqX4nG6yUQuPoOP6k
IbVWmFKvDIgFNbwZNT4gCsiULUEau23Te1P4mt4iT0GwwkOr8OvbU7mzpffHOOrP
Z0l9rM1cQX8mntPTqN6iWbmobbcwlCIKbr7FjoROIpphnnAYFRL6v/EO/thUGb1H
H0ZojrJXDXJKiUe2d/W4nw==
`protect END_PROTECTED
