`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZU9+i5fJ6h5OZ2lW2ga+/ADudIJlgyjRYIWt++wImMMw9eC/mNtrBnGZJnnBRq4x
M13/C47pZY3VahCO3swvOKD2P4ChEt5lqx7NNdTOjzjgKW+8YIzKPtC0rvQnJJY0
I2F1MHh24pFDczYv7Ii706IoHMZcjtaCiDPjlCwj6UgveWjNl+1EQeH37xWh5+73
6isHP+IvrCHldnsSTkifa4aq0UZGvQ+L5JPsW5HEUjNR0cQqVqZaXy5I82hK394j
gzoq9+mJueXfifLZfxMeN2FZkNkRZbVHTwYB7CUBG4N7FJQewamatOiggwhIVSU9
dzWgiDDumJDYZUCaFohhgCTs1+c9kAqBPYGCZIjBAYSjyHognZrclR1B1ofr8/h5
ZbmkyIYgFZm5YeAhuvYQER6v2EBfrZ2p5NW3fsQT1S8YhBaS9lB3pql7+eyDA4Ep
eOpq8vczA66A4W5ntv9XT/Fpe1u/0UamsfOKK6DV4/88H/m1KbZexGztyEiURd1l
XEi6lc2jeLhDt6T4a4unXBI4X9UIqhW9aaDvu5gyqjlXakJ+duMcVorTfl/6NIYr
FODQernf/zTmVWpQK7QPY+y+jjS/ocA4Mm0owe/+3Hj8mdIE45L/h0niZp5WnY1q
zQunpk0Pprlc5RawBPgxv2sIFt7MvTmZfI+5EAMI923nC6GW7qpkHWpdM0eQ9ltY
N/hgaEgr/EsVrA1wz+KpCOfv6YrdPUwXgLH9rqBMNL7PzecmOm0hgFzthJsLvs85
xIwo6knPDcb76nrhQr8fYZTl//P7daUHYpPmleuwyh3fYYtSQSydsopRT7ImG0yk
DLdE9VYsWZW2onJJfbK8OVo1y/uDkT2PRw2gPUloOBsKFv3mzzKJALFV8/XR+sAC
8KPhuwtZF3oVD56rbHmzHg4GvacSfhr2J2has4enxUDeq29vjWJBqINjMSQSXbzA
qJBo947v8mmVQXImUHFFbEsi+wNDD4ajjFXMsYsrNeGhtrqeeOtfJA1SLPAL8pEb
dUDOz20Dp6yxVNQi8tXb4SxEoV8XtF410eZsLjb/qgQ31uETd1WGnYAdtMV2iiuO
Nb7SxFVClOgs7jOi39bZbKLLXpF45pDYohxKCsz8cvSf0dz+lXVEA2YoMVg28HV3
daqnh7vaJcsOO92yUD25PINx5NnTJhRfT6QbJyczVGHRmaPr/uXqweODzSP0k39H
DoGwkOIjAmqIz7Ov0K4iHvpvnc/0pfreJljqz2xpqaqEYbHVf4pKqHeBSNlfKfrF
FSgsoVk7gSasJeaJE1B8d8qcBVcqZbjtCVfuvHfqh7lF4uzYQYdjXZVmU7h208h0
8D7S82lA1lqz7vvAU/MU78HfKlLfuzyz94zSW/5dD6kNgJSu/ombFD784HKy6OZ0
Hz0OFyeojo4ClY8svopsXy3ZWa1Jfd/mObDcBTJhDY00GByrPrcbtSXJCTQEaWl5
rrCopnj9/LogUZaYRFV1pKJKkNoijSI3n5QsctsUq7Y6CokSURPmw3HEJTmlIW5X
hQ6wIbs2K4moJ55mFv5F6tm0Di4p38t+NBJp5NwiwbnxKKCP84yqDbUXkXSYxbzg
/g6hso3/IUrt7MNcQr5TfxS+Tf9VpcY4mPPjAk1jGZAbwe1pb8NE3Gdv6wUhebPO
plWeIp7AR66G3fGug6ZXNjBHFDTwgpD5EdyODMlbfuPRpVnQ/JIMU9CdLuFSkOcv
7skO7F+vd28UoeHyuoi/kCD3kSAvV9Iv8JiKvGwOarCuxN8Q3AH3oGzsQTm9VqCV
y5bfRFtZ57AVcZyTHiK9UF1aNWVc+YJqbw9d6UUks2dy2P6wQ5Z5kjZ8iB1rfcnA
lk8hEm5Myn1sCGszPd8vc7FiTPjwDnOkTkt7GxYBxKKt3UfupLE+Zr/BOyJ9RyZy
6SPkPSBvR4nEGLo7B89qyscOGcwErIHgOWpCEQeiFa5fFudXTaGZzBB3T38fzHaf
OzsCMkUY2KalCe663A/hwmT6gKHq//HGmNX0lkkcKv1kOVbMJ5Zy+DnectZkyPhb
n27dkPjFL5Z/amaYj5HZb9m9stLnEzCrDiIqLZrvPlYarfTKsYyYJe/HJF+gFjXZ
l2rnuwBLc+rtict3/+WRcv2KTDFsjNCq7vkUBYp4YuPVUPHHdG4R3chO7Snbvvxn
o1vTFv6X5zoYnRbEIsmn6i9Q61IkIT/bHKZrQYCg/G7MgCPTSmpSq1YlDCaIJDyP
sd9ujsh8VFl2EvAx20MXMsF5SD6fTyiDggqL1ZkuGqJQm/k1dvUJPGJ+60IJhyS3
i/5lnCWD6bvdupR+Gr6mA7Dbca77ccQ4QIllHbEp6LxT7Sou83ws2cOdTOGL1ObN
dlJapFy3l5+Nh1wzY56xnlvy2PC8XTTAIxvqYyRbOtY+YX4aStY8r6ooywCRWhLa
hhwyAVgHOVf/lFhUvlvRt8KVnhNG15pF4DE9xzldVK9Xq9hBAmP96dxMZdeqkF9/
FmBfqwCoLDgAZwnSgQDMqatfySFl+mqbY4UcPACRHi6IJbopByi68qPJC77nsOph
2MEVjfhfkWXWU6hToN7h429B8cK9a4RGsTJ/gLrtKvik71DUBcnqkUQvZCR4x8kc
SZ2YlWL72NDidRSzTB/RsMmPKjkhHcu+slsbA6yHooAxwgM7BTYFzuIRE3SBMopN
3lCUBIkKGIUefCekZ6qHdkDHv2ZIuSQ6w/CnvhiXxeYfr/aczdmijGu7LfLV6Lam
ofS4M3MeNEomuLBUjJvyZmiFjkLry+WhasnsBrsPizRfB3UXlogqbBKfq6FZjKQH
VlAHqMEnKWSP9YdKpO9lyZh7HVRnutnuUNgJMcB4YsO6vjyVoIKkTJQW1/vsapvR
12dTbOll7r6vzHWWW8IYfmD9TJ/TbF4HaRR2XW+mh+gjFGRWbZ9pSIeZlBlpb2XV
PmVWzJOJDAWQ0a/VrkIdYlJVARj6dbHeAeKG0mWhucnmY42tKrNqIx0iijS6/N36
Oc+ahaapWzuUp3wdIvYURiawDG0g2QrxIa1uV3z/NPAXhdBn479ODO70BxrcidGZ
tdYm4nFNk0p2FmqZ4qb4mgSX8DDomlpFqquTuJFiirWbUhCvJMn3qPFRcJ18Eyi+
Kwx/Xwu3h74Zfo3J6gkvNITstQuttTLT3I0xTNuYeCrHIfHVm2pyYGb2PNVo63Wd
hjYAZyVEJZHLr9ggqFnX9QdF3FPkS0wKkDcXbFeLj6BIJUTywC3Zajr1Z4/pjCDX
1BvqE2g9raZN2tXWi0sIV6XmdQC+YskkeDwWZXw0JdJYti43lV9qeorLr8xhgEuj
QYQC4yxPZBy5ChjjvO0CaZLUYkx872zw6JTbeEjbWNAy1tY10IF9mDhg2Z3hvJVY
ZAsaNB7NDBRmZgIfD9TchP6hf1PIajQ69AOE+zmw24KaYT3H09+qaUf/9WKKdTmJ
yFYbSukP0Xy411aIRNdZCfsNEUIxy53kgEzwVMSaWU6md3DB3nFBjz08+DJygaHY
iKAdKWNCkKMkP/nuir1Lrn5Er/WG/Emeu/WYmQcXOAI6rmX0Zc2wZddYeEv2Ziut
XVWWs/ZNmP+eH1fc0zzIULpLwLux0kpxBRva1C1vhg0jOKp7msDCKs5GrMjhXZ9I
7jK4kq+JtCpnb5lM36fH2q1ar1lxrw9ukjQaWPhnTcCFn2X8zkVrPjGfKgO6nK/b
CkhoWhEPM8jtWhZr4ePZhKEIhCtxZ+M6sa4H0VS2u1J7Xbp+J5OZgwFNncAIuDtF
bgmJvR/yNR0dWBJCgoWXxGw2x44gbAjsReTsN+RuA6ZuWsVk2YFBLXftnFudBSrV
2iCLUGC9t05GfVRfiunqUT+fWcwfqNK4RlSchMvld5PXQSE3krfCyb7yMAa85VDN
dk89cu+vGKdHuZORbcKqmPFxyrbeRaYaSVWACT5kSjzCugBHGKQFfTJtEKuL3KA8
EthRlckgEtqy+b90dVk/ivntNGREEsURCTT752f4+YGeJaj/mYeupuW9mfD4RaCG
jUWTnpPfSkQaA9qeerFOJBPf6l9LyHNnBgyQa+p1JTV4eSCozhd2qly7KDMFxd5L
`protect END_PROTECTED
