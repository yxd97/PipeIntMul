`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rb+9ZznEHmkFEYdI7KMswu2mYfvS/WOCURxjD8xwf1uAMY8cor1tUGnxTf8qMws+
Ou1bZ8auT2AWj4/6dMdtFVrzjpBW/TQpCPdInigx7V0obqUQ6ezuDoHSHOcpHIbi
9bWJv7A4o04/306MbSXYicFMirL2vfYJzvzHF3WEv4WI4L6M66920YK0UWJ82f0X
HRnLEJvshMg8nFd3tKGnzwjSJEl5IRcVnBom3s+Eb5//umCrqZSEQ7dxYMy5WsGA
YwFlhTpL3MUeVPzqmMBskxRVuglbALKpS8FlQearY/9+GHJtk8EA0j2v4KMjQfOd
mpFJsjIBTvWSNVTH2d0RMyNoERNPkCBleqGmm1VudjGow/BVIFF2gQDt6bCKhpnF
l3eMu9RjfG1esfl9TeTEwFSWlhCBdUprunAaf8e+KQzAc+tsFN9tPIlhu5zJuyxE
DL+Hxl/rtJxYLyeVeLyL+wC5qskRwSCWT20rlkfT710Kl65IQURSOTRqXLDNxPjt
dXQ4UIVNpyyvToR/OKvZrDua6IS2nO1yjbiZZf5iDm5OkTx9Jg30mka/Bj194yUJ
vIcFokPKf3CmG5RkHgTpQF7GGSmnJWqbR5fSVhuEOcIAdqhpr/uhuy0kVjNbFr/D
iqSq2Yxnftj1V/6qzZOFcxoRFeGlJIper61yonAAb7uPrnCG2DeH4LlsBnCE+G6g
c2uCz4q8E1Gy01NyqbCUKfS7a44oItZqDbRZfjJoj6+cUKUaChpn9Wj7O47iAaSa
oqDK4E1MHL8H5GMXhZxjK8/OUZuh9eCZQYvapb0avJkSQ4HXhtPLtA1ZoduTEiHV
pL9C0c40D33a7NuMx0LFDxVqxJun2fZ68xo1EERsHdcXfeHSEftrY69RDIp88+6f
zIZ5yjxhhM75aR7Vi1j8DjYGmJZmYoe+DTi09be9ucAoPhRsFh6MYxUVN60hwdQ5
hRIyU2poagIIhIEufuiSDqPAr+gjMRvtJs8M0N83D2KYNY613IUmA9B4s+LWyqbk
qK0dD59uzP4nbDjRC8pjMsbHfLm8C/2lQBl5dLfwiTz4apPwByau7UiPMw2U/w9p
FBaI5+CYkb6+zYqCkMp9nZTj3gO9UQPYy5WIedKvefcRsgZNQpo2v/975M14JSaS
SLpE2SS5AMhOwibxeeOdn9waqFBxrTurfxCxG0Je0PJfPtK4BJ7w4BAquUBd2VeT
5ionTTzwvyGla81dQsuobPRG7jmAkVMCs7Ky5KVi7cPdh2r7j6LLWZZ+vrmM5kmN
K6HRYJmk/TWeWwmClrQVupbVxXtae//eidDcouQqFcEXOSZ8BsNYfLL1lBoTj0DH
GWtZS+KUTVRA6fOLGVc2PzEOHeOTly7WMn3lsOBJlmE00dpuKJ9nU+dKq7/e+WjL
L5/Y5ZeVSrz2+m1hEzYamhe14564gTVfsM64Bfi9QoUCiZHuq16WsjFkLSwAUHEB
U9hAoRrxGWn7wPZaXwKpLhIvvdUvwxJnmqHCZTWBX3FhWHklS8Rz9shiE628xY15
WQSYvrNDPD/KLv9OgmKPoE0OhkbUX/d4rkgjfdx9AAhxZgM2MtCoWQcbuRuduhaO
`protect END_PROTECTED
