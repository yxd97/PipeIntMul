`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UyTy1cQNlIKdg64Cd9R8LX30ltkSgssooQjMhq9VNgmIS11XlAgH1D+hJIW+203U
TbrpVfSyEdr/VNZOkAOfOddwziIV4Pqpbd5cF2zJNhUhgMA/VelluhGEcsRZLuvM
mHBlVrMEf+9crnGxEAWyRZ54RIHjm+rXXPJRiXpIbOJ2VyLWm2BcUheaCJDEGV5K
FiK/2iHLwwGqmAkmwHD7L4a6DYG5cVZRHfN2bKA93Oexcts6x8mFx49lQxtEPm/X
eBtxYtEy/wwizI3wHwHAEvsE+XT40nIXu4/dPvxPbvo=
`protect END_PROTECTED
