`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2qlHBAs4IJkHSEyXhI1H6MH5RWENTQ0+jPLpVOSQbUFwTrpvXhYlHyGXUAGHpJmq
4eb3sTn2SGv0Qk4Q+hjb0myG3ZBLLPnphLqmvJXSwL78bjj64pPcXmuY9nuyedK5
+jok/LAJgL8Lv4EDjqhr8ZnVw4cj1299nT410xqeLVZKMwHotu85s0BJBPFwddBD
mkc58cf9J6vtEKy0uXLPUU0hjzO1MKDV+ZuXWnkf/zNzaqJF5ALF7NAq4t7P4pVT
M1kCvU30b0Qxl+jqW35FgGQnfmUfxK1KYMMdzCVj82AGat6Eo7VJVcek7APQh/x0
+qXmw5ymhW+6GxgFWfA/macYdabb89TjZP/NREX8sxs=
`protect END_PROTECTED
