`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T12dC62YLh1Lcz50ibJfKXtR/Oh5F5YxD76favXDwJKoUyJfV4xeJCwZ/nuuzbGq
jYVW26vVlw+LilS4BY7UT0RUl/6bIn7ErRhYCLfb3zVmCYkGURtRgw+NKvaXp6MY
jjbWReJSYcx2q/P2G4k4tLm2keeFzeKCKlM2VvmBDhtoprme5cb04/MkNvJNxeET
b8VViMQxxPgGebNRpTeWt9Czxi9ffrr8oz9TsAbv2HwahDkz7VoJTioMCrNRkz+s
c4P4vXmBf1h8XhXwcxeB4ePVS+PPTU+TB8qhbuL5I7SYk31kXURFEj1RNeWmAoSV
fn/otTLIG9Dvf9q4BrQx3aC0UbmkYV+S0otkyrxbp5G/3c8BEWRKnUl+g8EjnbYb
P7tRtSpK1Gk5TKIrqhrJaRu0HsDdAX0tgqgVvUWnpG0Jl9xEKLz3hJY9gfsHZfIl
Zygpmo7S+Wj4wSdvf/2aDcxkyP6elSHjn8EY2nIuCs1Jqqg4GpDdT2ajwTTtODi9
IYS2tBYqMy7B2Vo3aQawjGP7eVwCTjXNxJSmH5MpS9ntux9RqQIlos+QcWhsuFeV
P3TxpYH5pCA0s8B08FmUBtgP4Wn7gPX4r6Cp71RfFT4gAxUAErSDSaoGK8HrfHXS
eQY2OfjzRK0yrpFw7YlP2hHoVzpcwJ3zgrUWIS6XemhnFGmPbhdH+bZvWNXqK8c4
PrJQFiqMs1+OSLOcz70EJE96jLMoqAzRlDdcQES9hxkkZ6GOGN13s4fRZPCOVATh
w7XcnV8JPZPmKpCMMpCNfw==
`protect END_PROTECTED
