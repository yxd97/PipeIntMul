`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZkpXTBX34MZMkafs4CJHiZztImaOVspqaQS5P5m/LqUkPL+2zGn2ZcybwBunaEx1
orAcM5Vq+SgDrPidXX5H9fckgso0LOpZ1mxH1mGKwxpjU3gqfcP1hMtrmWQMViIz
vZBOCRNJDznq80zVMD5balhkuesoBZOtJ/fagupwCWDg5utXcgSw7KRGeTDj83uV
QEaYX02GAVqb9pyaUBeXO8KOnSV8EUz39yp2kUjSio/eIVrQrnl/bcti0qtT3gAE
n9T6JEmlskT8J7hX+h7+sEAj8dxSuvdIAsD1KQe5kcl3r2U4GNBTvEPW2Rkoudmz
eoagh0Or6+c7ZsEsOqziLvdira4GL5lRO/d8gVtwto9yFq/KZkrEuPPDqn4zmYrS
2RXu19CunKjC8wqlWt+dKnHx3IG++J3wBkFpiHiDDnDEk7pBg2hcnZxthgVd8Hjq
3RQhQVRuegO4Y+76QUc/AB3ufPYeRtDfYzQRzF3N5VwGecIGxUUhyLA3NzYlR06b
KUlpVBcZ8ADOx2cwZwE1mT+F1tk2/ibD8MikMcm5mJZxOl3Tnkh0dkRVayIdf0Eb
BYwjIl00VjgkKyhxXXkJ9Yu8+llqjr4HdAXGOigfOArIU4LpQZT3Ptq4vEabf8ND
BGvMz1hl7fiJFUQQY7YVqfSJh4lGRN+qilNF2MN8UryCKv1+sK1pU8L5n92o3OuU
B3OxA4G/4BHweD8xnbEgoMGwFRbD/TFy1izpkg9f8uzpICdr9kqd6jDT0eygLOrT
`protect END_PROTECTED
