`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKOtl4lvRbNRZBSn2YiZDtC/OYj38Cg+MHKnM2Ymbe8q+vZWqwK1vS71o/0dq0Dz
FHRtAvNWAVtzriutT1PxNjdbvcfWF+4NZid1ONiiuGu2/drRR74YjoGLgTpsrTMd
7kOqqoztYejEtEaP6+264kJW1VF9+ZcgmBbeSDgIiZ2xNj9E0JOjCuH2I5saW06k
vkzkTSVNk69p8Y8KSj1BpnmugMcnHT9ZaQwBxEq8dPh1hRU4DWFCATHz3CN4l/pk
AWcvUb3YBT/SN5UzmN+49LQAl0rCw2YdpNn8NDzpOtn5+dVtmnkrR3l9BZpiZKmn
gDevQWWDeMBqvuHs2G+djgZfIG1ouuiTLtw4zTJraq8VElJwWoWUJEVY18RlKipY
7DnHVEHPVd/qn+90vGxLM3BR0jf7/X6kPQ7eh++j71Fsp9h9IhuWEiDEY+j2yZxi
hvVHOYg8FgdPLFrlNHdz5OrTuCfoPN1A5ioZYD7/YoeuSIUEiTa4QAt4W6iTFSND
SVdVXPAY6VqyFC64Q8zGkVhRfj+g3g5b5+59RDUVMP2RPcLF7ZuSTOObyuuNkUiA
TFgiB5VZ0QnkTPjAQlTk2g/7lYnW7h4n1qRE4J+ClMpXqyxtlLsNYeQ9btBoe4KT
l8bNlLyPLkhT6ZvMtN64iAiNMATzf9sDYGJACXgv3v/c/GthorH4xIas982dWsae
`protect END_PROTECTED
