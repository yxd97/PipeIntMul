`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZkII9Gk6m8jLVbHqNnm2jTnjXAoXhg9L6e9V6cRy4iYbMSA/7IdiUIfeVVG/o5Av
cVXuMRzJ3yV3EVoKmHFkEUAFndwmusrJZKvZBvYCZefhHwWS8R2+p9Usi94znd0m
+y8+aB9aSm20rV0Wy9HJZ7fyshoh6SpVlJvWpSMUf+0rd9fK+UtkabEchI7qF7BY
Rl6VE0Iu9FBbfs/NERDzKYD6GSMoapHquvcKg+mCbKfdRqRxWlLfUbm+URVKvQkn
0Cp9GuISJMS5cKLpRAZPunXR6HB9zUaU1r30tmfaQptFda0gHs4x1KCoDlc2Mf4o
kUTOHWjVHgXgnBNjrqHt8fvxMmKNcrflmTVxGHfZGl9Hxui4evDUTQsJ+x1xt+/5
jTuI3xuHL5mdLbDisPhAPMFaYA/MnIWXkQD8JIlMkNPHR1WziwkhOeVDtHMZ8CDB
OcN2Vc7TUQhWpZnGQXKihq17GuL1kMgwqqNeeweg6ppvIEkd1Uk8u5clUASNXXjy
xRRREHKm+/1srrkmTPT1dAztCwA54kiQX+LmkXKrwt8XGGX4kyvIBt9P7yoVOGuW
KbkjcrEFzeSy7HutkT8ciGXIGPYWXfRnT25RevllVefYGO4hvl5dILeGDO96yCLV
OBipo26gD9+Vy4YRH+vMEMN0o4wDPCOeCphfoeSt5ir4FeWv2H4iRnT+rdGLw742
rFXeY0HBsurGs9i+gwrURgmwl0bcsXIVIt+Zo0/BdDlCih5fVHnFWwed/NvkvGHb
YgN10mIvnM+JpnhWqPuWqjwQWq5UGwcLw7xSBq0WiTluu53DAqmOLzKSHzj0m+5k
QDi6DKbI2WY+iSCHQOdToS5w5XQ0/OL9zKBcK6prqSS0ZuUf1/0b1ciBN+pDQRQe
FK0PggzzBnWoauJyCk3FBKJDr5OfnzpcNojGUtP6QOk9e/6PP1NTX9bY6R4QPtrU
`protect END_PROTECTED
