`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IdcdtJVk3r+cl8nLG+c5QfhJiz8So7OkyCB0Fv7auzRCtPiJ5V13TdVdV5FW7NZl
1EisosgqmypCQyPd61dR9cpncl5sifhreDkPIDa0nj+dR7FWiHRiq4S177g+N5lp
b8xHfh6DU4OA2ElEbcKPo26m/jwdsx3YRBCHbrz0ZK3O2nvhzKPGIqMv3z1TLc2O
eLUxl1NJIvA8arbcSWiXJw55/f0XOT1X/Ih4fJzEYYuVYkW7cPd5ixFiBrOshJkA
HR2f6US3OkhsYbBMDNZU79C7SIVcTUSWQ9B5AblZ1WqemaoGDkHMaOEFvYek9SuJ
a2Xam6MrqxZOyoSJymxVb3hKNIUzdL4AoLAzf27r7Wa1xM6jF7bRIUMTX9Ee5eQ+
OteNxuBbn3feyTJIQiv9I0xJKEBuJt39jxnotGvmAvBALo1QpyNuDjFHHhQ6VpQR
kbgglE6d1BLOMgFBl69kys+Nfa2mJSRpscZMITQlGJELFpTdJPGbWcO+nl9B6nB/
MSspHP6tur71o8tvwCOM6tEffheXhjHpw305kNxtG7495iCasQqiEfrqo+c+wbIF
1EBlcQJPUMhsXABBOgqpDCsCnR8acyjLTs5zVor4cODeHwhV0Neh00sSXM0X6QnG
vLwm+LrpnMrBV3JFfVfeyngmWmZVrrksWvAnNSbRsApZrMKvo8x44jqgAl+6bJTf
VMMU3zNqVZH+zWGMNkL3esTqW4ry04iHdlil8ZVHzJcBDy8pza0e3bNminXoxv3x
oTSAR+UhqYSo+rhv/TkfcDK+T65dNKRRs8mkMi6DytoJxDOUcW86BfnAnqIbbkM8
OP9o6eEHMe3mZkdlbO6yB5TiOws68BSlxwAL3LB7K5uGTUxU9VYOxq/fS5PySSow
4PW4v0RRwkGRCC/GgxlI+glAAMVfhEkG/ROnAevLL+r13TJ5eMG4nQdKdknVD1oj
zFn+3z0H/cU0tEbky8ztY68eHDx1vKtKPWAN1nzgATA1TZRMWrE/rDgZv979Lb9t
rnG3PCqaQJnyfc9KQxM7nmC5NGYUVIWkokH0VW6xcMAB4EGB+KgZeBNkCMslij5Q
A9oRAsq0isWMBKzgPPiiAuXq+nspoHE44dqjC40MFoFQrU8sjynJneIUAGM9c0Pn
DGYsnZITfnnFT8r57VaOHFPVyBnbZwQjD1dEb0XEtu+FlHG+7HUPkeZv9+XgjPCX
v0N2ojuXQZ1ZPcZ1Fv1iuQcBnNcYT2b9m3zE7u5FicT3ybW6bBINvDtttZ+hjsX3
Tyu7khGoynym3tplxJlWedk+GNVPZNmyFW9MYiZ8k5KDpZfWa5Xukcob97uhv294
/bW69q3tq3zygyGN9ymsS8s2BtmrxxLBoVF5aKUq6OqwHeWtrfuUGGbfLnImP4aH
ZxXmVSQ4dSoy+UFUXv/wgq406JnCsjMPmitNsgMxEJLbjk0pzcDXWQsy5oAOIxjX
vb74GEOkceEL+Q3N8N1YGA4OaVjyxd5ai3nenSWlq7GI3O+ymu7Y2scZAI/pnq/w
UveJAv1dYIqiynmyvp56bXqWIeRL4n08NbKQRAA+tlv5G6yH0qitu3HvOqEUrg2a
Cbyhjna+SvHgvQlgKm5yvgupi8uoUJ/phx/KHD1A5EGB1EXblXI/BSaNmcxkILFJ
EarSbG5cczllQy2T6gPRYn9XG9phmJekZNiEiQs6z21usb1YLemeReCjy/0Mci8m
H8N5/rMuIFwug9kqu+rFFEnMSzQfxT+lIjJYyer1i3qxUGZSp79g40LuRnLYWbE8
lgjhoEnVqK26eFrBJSMnUg59n5TWHg/yDGbmTE4Jq29vWiEwvpi0CKbolmCjUYll
wMOWDgTOJekbHWU211Iu8mHB4bHq9lbfKB5yOC3ftf4eux0Wj6iX2uR2aHqUaaFt
wzaR/KNPw8TzSJj+o/dvMvA7zj5BFLQL81MiIe1UfliXCRiMvAG259Qin2NohKug
oUlb7tjkllNKF4IAvneHs+eAQf7faSUzHW4Skt4rUtUZYiqcjP5KGBS+XcAEDTJR
tc9aOxVRafGoRVgiqpftcuxJGvPJ0gQWXIcetL/DynWw75Uu6bCpNGpa7PgocgeH
YHG6XKG9zhESFNMXZz8VFHnupT4bcfFBodVNCZWtx35+zzpoPA5nxYdM97bCBoto
hNCJAzYchlf36zWTMl6xPsysphQBKh0Y+HsbYt8nK41bpb1BIDFQNKkJLQgXoCFA
MZFCtXfiXNLIB7VXOGw5K+HG3iuPPmtrMEDevQScCxaWuCsuLJVcECdvthmHCYG3
pU6+7gXS76EbjU5gkaVfF/ttxPwAN1BIisUqxfa1ZHUREqz28wwnU62BnpbuHluX
vtmBkQQBLLApwBNmujGMZ3+Nw/LfJ7CT2hf2GPcKOcM6Tda7T5Cozs32h6AHlIMV
h/IBZWdR2ARs30/2Qfc45QeYtbey4w21B30bflXxzETq6yHeASlWcQ+sA2Q6I43f
d/F3nnkWCzeqmW74m1fZCpx98UNdM4jjXUU/wdlB6+Ghr+3GKlMtl6CXa/CJYfMM
jwD5UBqvzhscqD6NLfYjwFNb8TA04sNl+fvRX1ft/b9hAJAwA0UkV7C7YaYcUKEv
2RCX6gTeZorneQNQsQt0PjskXFG3MWN35msB/b3TWesOSc+Rf/1YASSzUhc3hHeU
44vqyKin9WAJjTQ2cST+/j66tjOdi/qH/uSujc0UoQKhTYANZwmn/uAT7FMqP2N5
zBN58vUrmCwwOtvYYsAYGahcdZjc/ne3DagP2u0Fz7AM6dJSLnDjh/9tWfMRjLfF
0aVPd/21nb2wA9cqUKmhtSiKXfHIeeKrMM+cfB5aTGwII9vSQLTV0FC1YXwsypd8
HODc2jSzrxfEybOOAngzxjE55FBnzsiL8+J5s3XL1SYG5mTjapzrodmRhQlVz443
sb5XB4PL2pymek3ulxA4frYS92ALOPodoP6GJ5hQ8jopmTwExPG5+EGKBOukQiEf
nZWRzhyeeJJmT1+UsVIDgsJ3C34pGvIM51JB2YIIbMKCcOLg8cRY2225sbIu4Ynf
MYlCxZJ+5HijJR49l7THLAYKWoyi1EPdfwyQmUtlUTmrhGJYLz6u7Ga7MljLGxGg
ZFIenwH1gFE++XamVQWw0jzrh6xIUmA/Bu0BPH5t8iEFwT60wNLtAaNXeGsh68y5
/seKdWIVcjSu71aX3S5syHCI6wl4S3Z8PfHOAeJqnZG7NH/NYR9a9Oto+9tvLKZj
pPew22TSWMI9ZSbcPAA/RoEfalmPdWTkbAxhGOIhHNasUlIcTEyxx8EKk513mRMU
6v73Vez0nVoAWCUTW1bV+TgYaat6FS8rxOiQO1sLE4S9bLgu7U8YHEMfDT7HxJFI
e2fcGLH63UFS5BEW521ZP6EHw34fDvVqegjdUNy305mJl1M0Tp9E0qsN42WMVA7k
ql2OmqO6LVnfuO4nkqbZnnEoHr+cimVRR0hMvp9My4hhc5upefewDA9mdLh5bPGH
xCRrXSjWD6kuwQePRDwUK8XX0NxSVAxBIHAY7Qx5jZ80JkH+9DjekCRJa1qvu+Pg
VZF2dQ3O4/XZUxX8TCH/D857ZjzfyFl1pNIUih67PUdr/vuuOoMRrp9tNMeCbcxs
ZjQxel1r8vU+H4gtrAJqgYJ+GEpn40p9g+bYa1/ESTLsdpsFE3wR0fpvC3fyNsU4
z9d+g1ADZWT7PY9d6CQockH/iCkimT6C57ywf+DXd90hmLeXUBOl/seLLw/kRkS5
XFtcRbg3ikA6OPLt/5WKPq4X3FPsefie1JG69TJU7J2u9/fNxH8h/HAFg2RnmHk5
C7FZEbuViW4MeIRlnbQX2T4l3hKEDxOHJcYXFbEjdh3Cd3xyYcP5zzuG6vrCFpDl
iuuwKgvKuJ2widEO38eUrz0F59SaY9y+LSj5nZ+UVAP+2EXObbYjZ6nSpQfx6dNt
3SvlXVdeoSER6z6yp9uyWSD1ojIEqr3QXwgNBsTIPrRGrzswn2R12wMkMjIT0WFQ
o9XW3ZvU8ZUC2IWuis6QAlEZZ8huT+fwqRcnE1jIn3pNI0YUgJZ73BXIXMVRWYeW
Gk/tLtCbKZGk22kF432xV1tayB/rWnV8DapOm4vF2HS6uysKdq7Jd73/XVBNJwaS
nriHVLZLMEvd5URQkLGfUPeHxZjd6d+9BfEqBuW8drjKqcqhxlWVVK8CbM9Y2qQ7
f/xprojhjG9ZAdk9PJ/nlJ/sT0XxVQDQhr8FC2fRd9EWLoj6Xs3W3Aiujx+8YOUc
zLOOJMefRXlxEyPEPI7giw3e+ox5gPvpOFh3Pj2hsBrkSgKvzqDVq+ZHQQ8Jx7Au
YhFePhT9DFgXCOnyuW+g3TxP4+cLe8q9+5VEmH3ECcvyc9OCg46sxXeTO7mGsCHW
D+g7iQ7KyzHUNkUfmBiVKQp2nTU5U6fzCzUG1H0s+XJ1bF43Srv6PmFs7Z7dV7EO
/LxDLJf7NoG+ebpH8YECOM/T9Y6BC0IcHT65XGiLoWhW/wY+JBSEaOv4a65sj3OF
fe6n8JsC6wDpkc8ZncozXN2ptfaZgxpfsNGy4wAJVGsD6dy1LroqbAx0L4JO/uaF
7d/jUT5kPtVJ0EyYuEdyyClL+ybzKHCmE34NDcBOze3ny5vqnyZ3Xb4QHqaNc72g
ACxEQbCgdrAD+kkFdD8uXaR4KnFImWzXwXIhXmRxpKQJL3NEpsZwCCHV+1DYtxNu
2WoZFuvmek/IREeEwzPdvlrcTjgiUG1Y2RUVbztVPMg17NvUvkZc/FDKANlPorGR
7J706dk/2Lv1ax6Ex5/dfxHu5SxSqFgtqxvXS1C+iGLOtsEe2n7PTGnm6vkISiz/
PcPw7waIZh50kqTPcIsFpIn+BEup4DOzxFVRs2H/7ILmEtO3aHurPBTvtRGQTBpL
Hl7B1rwTQqaknNJdf4oM89bdf43GhAnD3bjIcI+eY1/4zRngUF3J+8ce2m1ByV4J
UCheGwRKwRF9v2hCZGB03Tpk14YAq8+OHssVBckF8SqGcxoBCVTTrN7eqenuiUF2
nI8gvEVUAm2c2UvhMaXEdwRKJRJtOXsMItwNEUjn1Ernx0/Z7wPIhp8m84favTpd
u55iiAM9P3sgh5XsCLKKez6yEfF5TGzjDBJrmv4FpXa5fvTiFdmMEQZBqgquyHjS
58PJDHOPurP7lnGVdYMpKr1pm7otNCjxrHNNl7il5+fPtruzdNFbQnmhrKLbDv2X
YX49GgGh3niXDjzYYfLSdoIv1dItzHFHTVY4OmBiynDqHpjNWY72S4PcJyA1xD+c
NbD4k/tU3Tguvj1TRwdYBJx1UlPFiGfMwMkCINt8LKz5XDC9dEk9Y475g142zzLX
RawoXP9oBKEb6kI68gGt5dqKEvzLRlC1ZEB+mQ5gxAMEJBmqj175plXOPxdp+PXV
f3Edj1kz/mAo7pJSYmBa49ie8dyXZH16+g+jBY0vTqsrP9Z8xg4prrIEB+nx6VBY
1i7OO7UETn5fcEBOv3zw9z+x1dcjoTbuEzZP+EuNDPBxUJeclg+XvhTdYbkIpSA5
o1EZCqBVmo3Jg4W5DflfxBBy1SUApro1KTqSubEhrStaW9QgaQHvTIpwi9Oj5msp
5W8ksqUT9A0oU1xhVxgmnCmsFNsFbc8b7saRmEiLpqKxK337zJuZhpnNceQAMxz0
9jqQogqD+Y9RLecXJcbh2P/EURdPxYq7EUugLtzZ0p26S4ZoZy0CL/b6t7uWfiNp
iBzl9c+T4Nfm/RRNwTdtB42dR0XJe4JCXNEXgM8+JopGBbjXzf9uVajyF+2v2/ku
BDHi92FKpB1MgaIgsKFFbYdbEwskaLWR+mjwGeMrz++ZK+fAD9nK7+1BleCj65ms
dE/06SIBaiZnETr3B4JqqMOVauCfVeHoM+60fTb1e74gS+oFK2/+GoHaG/1FOi4S
hpwfavDuXvFRnqXs3jNHj1xmXayn5ErWHwXGrP2bqZOnbn7SNyWV73L+5ChIRqM9
gn/Gy6lzIMxe52AwVQQTm0G7JM3Vpba5NHC55xgiT/YM+inYv9+VdS+q2qxo8oQO
KcplGg6zQUh0UlqipcaggztIWle5mS5OfrQVBWgz2buaqZTZjPtmDSPGPNxoxgjo
yQbbCxopeIrWSOwDgbqq26vPOOOyoEDlW4acFYddf2upW1KNvVaEf1iBgDTOhPjr
flNWk6tRd+sCReCXu75hY2ogNTw8HZDJWCeXGjN2c32F9wtJK2m+OTWPYs1I3m5R
aeWlcSjkiF6zJtfcVJsc36jXLtrUykw9wcxj1TiSJpJjvz+oDPgBq3gR1qeHgkN3
X6VzpdKn07/f1n9x5mzVtG0p6Nai7UJOi2p5Di1vK2ne04uJJTO971Ic7Vg1QAEc
G5O7oIEpEGGLgAxKirrBDNVyxqqnXDO7fvVGROVoGjENNi4iIe8toMWs9+o8n4BF
aXMSqkoFLV8nW9lnQ1++0Q/SOBDewSwKDN8YzBIoVwWL+KzZNn/4X5ilHTX1hQSH
lNPz0Q8HkaMxwO6ARtA/xrwBgr2aowV3HAXso7vBXHAvdZb522Xua+yB3JWOPywb
D4zqNtvCCYN3y2f8K8Jerd8D9cxgdcv+80GJX1oxt6WNU4mb9MWPG3w3xd5mXnaL
Yyk0gqRPjkV9rCECKjoDFbQDvq4RJWOZ4iWLD3Dk/DmXGfXW30oZGRCJndVqPFv4
Y0GJR9ollnsl4XDe0AJgmmKHC7h7cGI3yNB0oY1l9krjBFPiMTCT+kJTs8+tKZGR
DC/3hLmuF19lmslQUdFhYGh3Sl4D6SHDN3vUTdhezrxIg4LbhIXz98nq9JFk27K7
bZ/LQ8cb8hZWkJV9+9uEBZSo9lnY3YtEl73uljH/YfptR65aQfy72bKMa6icvQ/W
Fqe4YBxCDBUgKq9yX72leHyT958S1h6ECmlw042igkFNjpyDpRVGZewOjQ2iuKa0
11952tM5Q8DJDdZfO5mojhqRCAXXKsW5Q+smMiAZ73TcG3zmBV19wayz4rsDrQe8
93+T1lWKVyzmsGoRRKEWJYCGHkjrYzMVku1wHVKbKXq0SS497tX8mYnoyq/zmrWw
MIMFaKm4tI77R6jFHN3iWgeJ3D/Kz8lJXSGna1aPIX33fWXm8w3Me+0/mHFmhoK+
ga2B+ZR6NNYEadTGM6qy/Wna3jCeobnpyT+zHzou/O9I9obBIdKrzBRzaiJ0kyOT
isCpCCczR71rRQTbVdEHKRU43/pS4TiOqGiAE2H/hGya7hEE0dWYNa7r9bI/Q1QC
oAHIuTkK1lyu6aesmjncA8vrUn6CL9bIs7v8vseKWrY/7J/gCSyAgC+SvMIcXbCM
9pTVZnclJeCzrZ7jX+slwaIj3kDVUPV8SZVpP1n6C5s43WTg2gGjfi92+HfOd+22
PgqxQ7sKFY6Gxq/6EDcP8obLj2UBz77cinlQGfQ5sSSQ/U5ZwQYvVMBt4O50OBhY
0I2PXjMQqEZPEapwBTIzsMdp4yNiQmxNw9WZdOLar972WKhs3pBoKDezuVm+UUBi
X/lpnxOosVySCK5BTATT6TcoOCWeOiM1Z8oe7k29Y+84TDFvwRnZkg0X7rCsF+RV
yEbr5jGKRziz/QqDBktIgu4b2/UgzRFhXOcW3LSDlmD3OvUR7vdOQpXB92U8+AnG
Mjkve86JEgz8+6rENa6pi11mDYBrK2WThATeHDUEy9SloyjLXRtXL7S7Ka0zsAam
sZgTp5fVgxAimqQPwSh+yqsr7cAT7eNp/mbq+HvbedeytP8zmb2BJBJqYLIFbEdv
brrFHa2iEj+ydawIBu+VOk2xqjzDOX6dz9jwrgBaZSyjuKYRTryVnEEyT3dYri1j
7t7Ie5A/rYlcbznacr8iZpQbAl238PqCe5gcIHUdTH2Uw2vnFdfSa/dzLZ+lNJDQ
lMhvwcWRpxsEIgJYwme2IkZHxogwKAXPhkxu6SrArFNAfWkvjiO/S7x6YvqIbtXQ
gHGA3vgVzrau4d7IUZ8cClgr/7fkLcM3Vg5RoUe40HQ+oWfVCe/4v6xbCQPlIg3M
v6sltnZ4bv/xe2NoedefB83auQnCG/zkS4XbVLgbv+aMmJcw9Ado+aW6vpDgp4rD
DAu6zol8vu1H7mU9L/7/l1MCDHhjGfY+gwairTS/3UxKWRyNywQSRp4bbpKuWM4t
vVMoTm4HPt4SiDssk+3CYbLnhqq/YLZXNCZTbxubJ54FT/w69jsfT91kCwKWjuZV
qg88NXDUUgbv9T7vqCAqmLtF2xnQRu8aOQ9yrCAsh7Tns3VYx032CtbhX8Rgl4vO
L5j4OLSy819kqyeRcJxU9yJsgHY9RCX75mJDw+pGGy9Io5X8G/LeTDQ2wZPuVrDA
C8XmRF7HdXOB84VHfZsfHfNHp0OF+9o36AANPKWRgceJDhRMz4scTyRnO0vC+s/W
+9esOusx2fUBdQ5IwnwdhLUYn8vclOaPWS2D5l1wcvTC3w/j7kvEjJMJH7ret5S7
GGQwBDQtpcHsDk2NUlCZ20pnnQ3Swsx7nAC4lu4nOjU+2PDOxX3B8k/P/pgmnjTP
Cck3r/7CpDCpub+M1QIvDnR+rmJS/I2GDh2u+8qC2kbwYBvrqRRCs4GDc311hjUw
U3w2E37RgSboic9ixpyBj41MR4Qgw9CGWASZiI2v3sDA4Hta79yQC1avICQwZHn9
9RzN2Ji2rbanihr9ki0esFZ+3HpumoDmSEirhlGyb4EV16T9lAgp9X16eghxh6Ey
eFBHo4fh5HGMY9HLkzsMOlVUTedyLYgPa+fyPZvoTgvgibh7m52pHp1b5wwz2yfv
MUChWHAHekYWktgKd5nC/za/aausRu8Cjx9VwdwQEMkjL3LKAPFhdxCx4BjRxpZ2
el/z2XYlR4ZWrCwJKj4Bs/BTzBMW0/qzNRkoOh3xvrG7HGtSr4eQFX5WvzYCF77v
7awxtBLjL3CSU4ow3WJanLhHuIyxe9jDxeWCw/Glj9IkYoiWwBeBTpreU4BBX3/s
GLIIH/7GB2SxKIvaNCDkHpLMlFFWdGl398FdKHPspF4J8fhtaEv+XMJEB/62L5VM
djM/A7vN5E0pC2XCdpBtrOeNmVmrPX3PfCqBX1OhjehCQztWdZcQaw/1u5C3J9Xl
pPWQ7lSJXPkZAns28IiIQ70NXH1R5kYpONV1jV69N84tktL7jnroHBdcpI+esE+J
EnUoj3hGb5I2dMWqc9ayzG+675EJUkk3oJVwatIRwh82vQ2NmjPlJl71u/IS0qQJ
5GUcVS8No5SH2vciDGQ69cIbv3XFcisBiJrLXaBU7spBR0nUaNNH2xz2ib3cFxHl
njHq0C9ADZaCa5gvpu8tAUhYQ5QlBuXIX8amllU+LaC47/DnSyfPvd96Uyd7PDAE
/fxe4aKhDusBRnFzMzy9+bf3lgtmNG07cVbsDW0x7c2C8iMEVQk+faaaaiQ3SlSl
SLFfJXYldnTPR01T6g1zZFTMhHvd5H7THsMTtNuVuXCp61ecsaUxsnI730ePJMHC
o0VR3+gFtOXmoapsWldvAu03ktGbSDjXDh1zBtv8fwv55aFFCYGdI1f/KQEnrHK6
hzYA7/GNEcVw5IFee5ednQFT/fA83av4cIr1gGuPl23uiOul5DaWioMsYolmXftb
JYFFLZa5UstdqCZf/1CUjmWFP0LwjTFY9S2QgEmYAFeuT9oMPpcsIFXeTt30Uxlg
bPNnSAiuZCQDgvQAocYI89ezkeSsyUoWHBJ+yWMjTvUOPtxIj8sItT6YOn4j427u
5PrEXwjVZJRiQqllxHEE5SS+Pf1zurJSKYYodpAPEH7doyuMjK/bRwwxoDc3uUtY
4566R0oe86Ebw800s0x/WFCwlf5qhnA4VjEgYJh2k5mG4fBVX2UW4SqI/EPftCDf
thO5wDIIUVf+wWlryGPY1OIt3L/c+2Rrw1kdtNJTS1JS+IhuIVoTPvEl6LV+1Dn+
4TdvnTSjVLFog1EqkFZoOmJq/Fedq1E/MMwstY4sa4EEYQNv9LnVCdSgyic7C3Jw
8DZd6crufGpGWmwXDZi1Ntgx1Dk3fEKH8Than7MimGV1tIDN/tUQ7iMLSMT6Q9iF
Unu0pqmuBkmvcibw982Mkqn7Av10jZoq+oiyDpWFj83YlJf8Gyme67FeUyd2nVx9
fBAHk0MMlPVmwk/p7AOKPjWYk7UOYnQtPCPnnCzwS0+NNSxs0zQo4FaiiFu3SCbs
0BMjj7u7liMGTXUNMh7/7KCASqsWlh12Xkq76Y219YVPLmzybxUYwPSq42YuR6TA
q9eFYv3lu00JrUvyArfmhva+Gs8V4P1qT/OREGKwrRM/fECwsKOtLmwpZsaz1uCQ
5KYGro2KKuxUrH5W25RmbXYUb2NEhhRbc5ZFoUy98HzPcLTBEJTsDKacHYWxh4je
892YL4q4LpOZht5FIxzi86z6g9UcRsqi6Z+d4AkugGB4dejYXR9x7ysE1VpMMGi8
KM/iGuUsmGIJqZQ1OoQfnDpgChyVqM+k3+A/KQs1Lqncjmd+2yx1GAiMJZUlvw2/
REyXmR/Tk3ON/YCcmHhobiQl4e7kSW5iILOueGEz7T7vnXpbz6KtvbVJ1v0Wy/ho
+YpXFHu+KG3xerUKWNzzouIqJJ4I6Q3xDDcfPVRH0RtGV7cgaPcZgXbioDp1uKuP
FxpXfxVQTIgH2g90cfxDOh/cPyYNzq8zHIulmkUqP8l22NcRySNEoIO8pw60mmeU
GQdQeOJJnk0vYNwvmvqcjekVDUWk+bgvQHO0pMkgrt4hs2z3esxjli+1nu5jQkaK
NQEHdwTaGxk05Y5zL1JLX5CNDh5POMAi8Nec/Osk1nID9kWF5jSuCyPiB+cG13X4
yhijDIU4MVU4ZKPzuByCwzoiQ2+JTFs1bqXJWTPm6uSQDpBRzWE3pxZDaPEcls9b
CDyABabz3+ugY+adpZa/YgPzXEfYyinhPezyzoDEvZguY4h3NK2FqOtbg1iHgMgJ
gGH7cOoo2sPpIjylg7fQj/3IVZWVDPMVshSv1yq6eztfF8iAqwIzT5VcTC6Bi4qW
GzjgyQ+/HMowLveQWprjO6AnQDPuxG1sVNKTX+mS/4Y1Az1EOC4yj1vumhbZJiQy
yHdlhcatyXStdm/r0MfCD2WUMR4UG3YdMv9wTQlzaXW44mIQVt1iWFFQOHmbq+qY
VZSeT8KG1p5Gg0dKbFlsWFePlC492ldiIRU9CLfki1nGM52buj4F0KGGsIfmYvh9
OOC1MBMhGF/YNED5ifn0VMk+i0CbZqHi+/UPMGzu6HJBFK6kgYzCn4kCIVxbysA8
Er3Q5DUbHUOhHqG5fHkhVcM1Vq2wa4gV/wgOVV5669lX47q9vaogO0uqB0bVB0yw
SWaDLJLmzRZsIl+px1NO3f1KjkvWAd0LyKQUpEGavQ6ZuExViWoQzbUBkxJbZtpj
gK68gJvuOXL/Pd42CmvnTNo1Pixaq9accBkA5TYoB0ruqVgkpsRuyK9+p2acGAxo
uTZi3EEing8n4rHvEvQbg6RLMK8Cv50xzX5VwfyOlBkia+VGwYQ4wktLqWRYH0YT
/9gUTBIIUFPHn7nwtLo14fGWFxHyUYmReB23OSYJBzqIEbiMrtoDAZdQz/TmB56h
MncNsT1/YeXvUXfQ36vHCE5scoJANLfEKe1dtBtKzlE9P1TfdnfTW7kjXYRa/P9J
ddry5mDCFTlWsiGGfTwgskYvSYNbKKd9KKNKvmU9xVASb4E9fvhCM3wGGNBqOgYc
2jHrxHCPrmJNBTjinDM4TJIlE2fPVw72FvobAF5a9c8Kyyiwklr5lECF5Qm/RX5C
iBDnbm0himwIxjMffzTAK4/YEVr1qjDhOmI/Tsl6EhmQ+wjK+iT87nch3m1lCKDh
BBbfYDFXJ3tBQM1PrXNM5BSXwahXM+vcB1QRiQWftm7PL0edRi/F8a7E6QMqk9aU
EbCRtEj1zSv49IeXIl1jJm/StkGQ6J/5/civ7IjRdyrk14y0qn0/nLfuZvmuvN5G
hUcOCrAzn8oIH3yCcn2KVTPy69uv5sNFEDc5QxwTviSIJ8eBDR9ZR3EvkawSuKOX
FQufsYVcJC5G6jNFdBXGCtlOt1lN/YR63ujzJjQButM4nRDevURO6gLp5Muc1Suv
R+x/5XU9kKx5xIfBEfz52xgpviyQhnRQQWTfIPDRF7TdtC5860ukWiy8vAjojDzh
83kO5h/bGbVFmhFAVtsC2sUsZDX9lZw7KMLW96diAwW9ZRKO1+Ph6xExa5QFLzA6
7sItLC78hzeoSOCCp5gK3VTBtRhforAm2WNusfCqbKT3VexXTlD+BKiCUmxJng7g
1KbqemGw4GZRK/Sdtn/KGly+wJHpxlpKZVrKcAXZxCTo2QdEIfz+ohd6WvyGhOJr
oyeTXbX1Zblrx1SKsOHPoIF3qxGShpGvGu68x6IxJtKRtueabMqH7KCD54hMfXTD
+8oKzUNPcImWac2BQs6lVL6pwiyTocBi0gdywSjYundwpvf9mn7EErbQoGm3+IMu
tZVpSn1BP6OuRWcE/J7mGcRZd1bxaSB+CC1+YuuVxb/NsTvAq2yOUthkFO4Rme8s
kMx3sJhu05IRs0hX0ItQMy+Cgp0YXgDE7fbcvc/T1JZiqF8lAoP7PD1htI7WGsSd
WY4/D2ETZ/Qm20aq+Cwp3rlBM492DYjapnUjPSb7bTIQd8qNBNyG9Pkc/OCkW9O+
pPsENGIIy9qidPrLuXTbtkiQi+daBoGEIdMVrjqLYDaKWwj1QatRgF7ibA7fOBdz
jOfaI4ZHpzMQQOznPx52XkKUlpCo1pLwPWKqpM1dY4xcE/gzZk1jOdiiArgYbJT3
BEfH8cNq5OM9Yt4MFV0M2pgYQ2EMaVPD7u3JeypJ+JlS8B/+F0oaIfSfZLllDIa2
AncFp7JGfMsTaMFZ/Hl2NiGFBxeNnb1paCeFII21hwg/vqGNtGmfnHSUBNAKSxkn
BaWH04D86odmmo33JrhUbDqML/htngcfEExIzeKKt2R2X/e+IbsYzPVFT/hpMtVe
jtGR2aLzjeJdOvqdkep72rBts2knswYdLFHtCbPJgVYtYPkaz4IynydNtRRQOgcr
Ar+tOREleMX/dgz+kYy/aOu62xeXt4BX3nKaOkGwosYary9mFMqVLLnpcBQeGy85
xTbK+W65YPj1tiTCV2Wl9dzcgcKja2GxZaEDp9J8ItIB+don9tYr0VtKNrs/K8oo
TWLpGkUONi0wDWVQsujhrbqd1XF7YZGcisa5x6nx6rxoMOChfH8djLOKgUZN7y/r
jKv8UwmMoz0SsLYKBeRvdj82s//UZWFcrVNNE09soq2IyUPeKYLYNXJf2UnAzjd0
FA9EAMbjbvr3lLs86ujPZBA+Hs/wDuU5mNGtdQqtk7juzfTmcVjA19M7eY7ZJx0i
sagOq+89K76eOLxiN3h8tWsjSrXxpzZgUMFxmc9hCvkZ6wnLRTA08IBiVq4NN0IS
/8W4B10bQIMNywPn+MKLDhW8qcCVQeZCV8nqAzgBe05290IyVWb+LnjKgLg7WNSt
eXzzQcjSIIvVAf5IJqG+PGEFOnPZ9+jZiXOhwqh/070yr9046edsTXRRWHeMxkFU
90/j6A8+JxUCKuht9pSwNCrNqgC+JrocaeCVy2uwg19rULGkSDrWqF0WG7dFLv5O
aXlSH8Z6b7wTr51qtJzEqvLP1dC2BROvOVoYEchsEOejPXLMyfcWb+ACAypOA2d2
+Huzg6c3BO9BmXFJDpcNnrE8JFSS4gyXEKTz9ATTRT2GKCLUu2TakS783yNFDHVC
nNaqrjCncoQBOURjYDl7NTNXasJcEfpk62rnQxB5G2kElfJIYakM0HsYAfhwJmeN
MbMdh9F/FTgPtJFyii1g6l/X7NNmiJrRmYajsWGDZL2CaSXxsWO6g21+8FQ3+GEf
bV0kIn3GAnDScszAzT69UprD/hvE0FY328agK2vwvZybuLpDNzN2PACI+04X3d47
bW8CG5HpMvAlxxiWQPTuUy34PzU0SH/kLtVUrOvZGLg8jHU9xFcNL9+1HdrBJQ4R
IZJ9KCoZ/FT1Dlqz9NM19p0ytVpdb2978Fj6VVbM8fvW+Fgp+DH4p+qTjudxD9qK
oFSHGAxjEa8ovLFkXT4o7SmA22ioL5We0hpqbb6SHsPvnAcpjQ4r4gO09W8dFfha
W78VY3+LPbZGupz6L6ZOP9W29C5u96/LFumTF2qMMtx3XFySH+ak1OfVCJphNLbo
6BMV0JDMb9kaVvtiPjniZIQ0dXr8OX0uFfKOzExI1k5Q48kMCFAET8SULvgBHwK1
IijTDGH3q2uYVe+363noUEzUQ9YrCVnWC12hEVOu3yT65cVRD5dRVuSb8KzujWpW
1dzMVCZ8s/Y2cFWVpvLkW+Am2j7NacyYnkzSs5/qw8jY+oqp8d1Mgv9wsv2Ly2am
6foIZbsj2vEbwgRSbrV6NB9hZZ0rMtyDYhwWZeNN1gC4JBAgiV9LUTnjamLGkE5G
Wy2Yvtscei1TcX26HtoXmVeDWQ4aG6u4QIRw6t4cqRJ5lI7xWP6Cz3AdfAzDxSuI
VzEAIJTOfIf8iLTns1guy9vSyk/VM2TH1MU2BSw/fpVyz4ZHFe2ZTvPxjvfPTUcZ
jCLbIWjXgw4lSCxpgeC7yODZA4wFx1q75klBLBWnw0ATc6m+sNVMwAWER8vf//n4
uHh/fx3w5KphBdgsKyQHOq8iQRV+7jeOY/03ZMWtEJ3dKy7+WnnSSqYYJaYzRXe5
wmqyOljluOPWm+ymTB4RAbo24hzzETuF2vei7kA6ky8oWV3U1ZJ1T3z22XmLawX9
h01DZ29PEkfqoZSH7XuTmOWW3pSvNQms5QEGl3NWMdSru/OdkrYZdHN/bwuKkFoT
fiRcPJHVL0xwtEgWoPLHhty86yHEvdH78qQo7UBI84QruXzecH62wlzz69qWcMJI
dUm3I3ExDe3o6b7NYRM9hrAfAUIhHKYE+X5d+A7fwZe7lD8hks/v5uTwAm04U7mR
0tvK+thrpmtBuYHipjwSs96s3r2QdBx9JnJucn0tQBp1IHF7zE2uCP94X2zW7HHN
efZI6rqlWik4ft9yAPtHAbRG2Ft6msizObnf8dGt3EWOsKe8AgPqS3cqkndnEA6l
ad/ltYvwNCSLde3OMu+xIEFKofrbkADa0DCB3pLPvSop/MNcTWI/ZQiRVKcl5Kj9
5q6PH6CB0GHuxoRP1RwFw+rEDgWEFHqUSH5tQ3ARcK9tcTBcLhSIj51Llcylb/bc
UDUoehMSKdMgdKVocSb6wE8mriMcEAPp2hj2q515lhtCkirrwx8LeC6SG2GM9dLS
mVaMcMd9OeMqsa8e9E+/9f2gc8BZT6r+3Nfz7N4zf6bJZXz0Jv/Vok8rZeN6nron
jPZbymKlHTSe5a6liMnDdD2y9katzKQmcWGafG8p5VPcg802cWxRRnUAtrQjUVq5
MemXALYFyRNAg0/WYK1n0UnJiSws2JCuQKmTaWykLLHL2BNWO9jYRa3tlkBjVQZB
QtcwvngCxmslkktGap7aGPio1htwMx6TrrvQOTu0b6ZZ6ia20fvfa4pZuF8nO6xs
HTsRS8mDqNNbzl/s1p4qNbE3gqbGwTHRPHNcyd+85LSnKghv0G/tY3tIkhzT7/6A
XKGEokCFiqGrd3eU3esjvBWay2nGrUKF4bZ8WIW0E1HuusEJiRq+6z2MWBNTAhvP
oqeu5t+jYYsnw9McGb3VgKz2C5Rm68N+36V28LJSTpGloD8rUFx0JOyGcONGKuTw
uC+9kKHMbKAWbvjy/QE2zQxE37Q9+nrtyuPy0SR3yYgqrZv89N18Md6mdcbjhOFs
pVsmdfXKwVSadcUF2k5oSgJY7byaJ/NVKEfgD37FHjd3033/8eR17O1KokplVncp
JlPTx63/mqQ/YFK+lzpt0gcnW1snEetGvIZjpCVR1MhV+kjdrz6eMtuPbrg2KRVs
j8Cm+hfREHeMKq0CcbDauBckA+U+fIFIpb0UV7UjlIogSNTyuPpJggpqWTHKf6Z+
GQ03V+X/42CuEXUL26Yr+ec9RMsv3bxueVDWLkdihWG96qg2gKm4L78rV9GI24P1
wjDOK6sdLmSo5jDqFiOBcJRYmpXko9cjkvkRV5vlA9mHk2ZaqevSlFqNF53lt6Gw
YIMWUjSbldzWO+4NQT/e2yyk8K+DDzF/R99B7RZY5s3RULgsABXYWbvO43xWPeJP
qUMFEVASIF0j5OeVfIW8dkRIW84IvxAc/lQ4wVyYSVAvLH+mXIW2hytRJt609sfT
BXI3hj9q1yY0ImFP1HIIszxNQnIyorNTvIbq7e7ffj0aXvv5faAkMbQGMik/xBkA
qwQuL/2NJqQRwXf/nFN97wCMYp5oRbjNX0pwWIqnQdnmXVSs5+KYMdUDAwuMoejA
PegjeXvlssHLGalcxoxBKp4pegBScjGQVEIwk4aFjq3w1Q6kADZTwcbkbJ55bkJC
mjVJh7q7RGF4zU/A60IvOMNm7TtYrGGFpyrh//9/X0bvU9rLFoOzek6pxGvOWUWC
g3bAUhqX1yext0fxonHFTfHRhxPuBLKjfkLeWUYJ9GT+T8Ha29zuV4BpCD97oagB
jyzB8jJ4XME4fjqf86E/G1RI9jChlFGQE8rJyi/wingIXkThPc93sXrGiRD+eoac
z6qLdVrhxxY/Bj+YD490M8STN05Cn1pAc/DzMKerhL0+hTvDKFq4W3aFRbjDs01F
MUHgV2mKAKE0RrvliNlTQpHSPlvkcVaF81Epe5eIaGwWA+oHUSi+nJp0n4lpOoRn
qtzQO7xCrI+4Bl7cYJA7IlcSWo8uqrG5UL2FpQKz4tUsLtageEfxbOo3WKL2/ytQ
2tBe8mbF+QyYXaD31m+Ugj9H7HYOvNIYoTF5D+96IjtVjY/tX/5I1VBKhFx9nTDp
O8IGsHyJzPnMQyQY4WXhb18E/IODQRwsu18rmt838x+ETOXolwpoDta5T2K2Us5i
Aq2W35uRfFhlfPbOAOiqfaLC4xOv8JIs8cXrZ8Rxk3s/qhLmyIe0fe1Hv900tHVu
/LjnhRz6V3ngUnHBahnJh+gq5xK0jBcioxmA8H72FYSH/8DArrSo24xgwvTeWbk1
CLY60qjyM9L5SWkEecgpmebk7WutCSFIlA5Qf4OOL1z/mR0xLIFkUWw3cKZ7muDi
6Wzqear0O+OZ/Q+F1b0lIKlt/uqH7PR2pvOpGZjnBI+OsejesiETjUU0Nq57mbeT
gmxzmsjwwfWOMVjouc+R278PqkQ0ucDewJ/w8bI8ow5WHvOvKCpv0vIvFLnB+96U
tNfkVv2iE8VBszqoUxo6AQ0Gf/wRnKG2vYsUi5hshX93PNAplYiUSlXF1veIF9d9
gDhr9vv42ZH9qh4ijkeF1rPTPaC/94/vAbNxD7s8tZINZziDqKyw8rL33inPyOmL
xhiaHxiFwk/XK6O6tAfZXpXjes5nzm1u3lHvepa5nqKbhPs2NEhhrakhTkqt440d
+vfmCk9OEiNjZt2CxJpvBppKFjidMwslWJbD1N5OdiwLyKd3O5p6zrn15JThparv
/4LrFlaSXtX9jC4JIe/ljUGiTmOsHm9OxGiMFUlzcxFvZS810f37fXHzOoRtmT9J
UJklfR0yrGB2wGOJgTLmj9RoQNlVBbeubytZOPtyM8aQSsxvn7C+vNOY51qF3cLp
gmxlpLEENIFaBVM49Thh4iRfgDRZ/WA96gKs4jlQqTZj5NpQZlUE3+0fzy320HZ3
X5VdMV7Y6y3/KELRCuhYavHXem4ciXrhnDS+ljrzLNDA6f0pzxE9rGOvmxjcPNp9
TmlDkFVogDbGwonBGztD6OljDhVadr7HrvRzr3vO/8/nBKmplxwitG/a6pSscXh3
sSpLlbMy8hOJw3eLF7iqmkuGdaMYPM0B9VC1et+NQbLEaPR17t5i3odvADP8iZQp
divnVlAonB14eyHdqPCDOvxsaEN6Dj+Ob9e3RLZhRann0weH6f0TdVI2zceiVbcp
uByQnVNpW4r46+Q8qa1/kFFyv+8UtM/JIRi4i48DANA7QNKNf+Ik6CUVT+YsqWeG
9hfNghfZ7Hn7TatwL2n0R0JB3/4RSIBSGjFaLu6TGCLhpJBQYAIeYNAcqvMF7TSl
BDlLl7PMrG57VGehLBbtBj3N+qyXBgPjf7sSNshDoMB5A+8NUOhHHRHWOsk7CUFD
dTm3PzVDKg6f+VH99mJXRbLxilzTUzWffGzxOmFwaGwaEDZFk1YUVbQQCS8iGaDo
AOOgWiLWGRcsDiQrFBjvL1jDvquwJdWZUaSP+FOUOUp4gccJeiKv1HLtPgDSNvAy
B5E0qh33SIjnSPdlF/UwKVLbXWltmTrWzeyRAqACqtsYjBmC8Ne4r5DBzu5VlbCD
9C6u+qogJX4FuzALWbM3zOW5BgcPHfkP+jacvsc9irpDvhrzuUs8yaxmiWtKp3DW
+21xi9I0SD9TCm7mC3M0JbO9tAbUrqDIO+XQ/heGivk4y7Jn+kppyr1EBUprQenz
IdLjANqKRtdeA+2gwRcqou3nGUG4q/Y2zBHhllHFrfuBKa4n3tRNaGpBblISKYFE
1sLsns8fpDlUMcVdeRzA7f93bfo5dO2x2a+bHc24fmC0KTTw2x/9Ux31DWFlEBPT
4sBkLBNXgrB+gy30moQT2yUfUWIpTXOKo+3bMrzl1YNEJRmepdU6zFyfKBafDm4/
a/gWAOWyVQqWSuR4hA68Bsv/w8uQx7sQmxPp7Wn2SFRzF1g5qi7TNCfINEV/C+MO
WXwQ1f++HI/6ZOCYm6T3s8i15lCOZxEYVU8UlsYrhszMkPq14Divjf29ovrr0mqB
a/C6iu8NKwav6LW8vviM5usAe75VyTOsJj4QY//rZWgFfYyXB8bm+9dmBM8gbwgh
/uGG9C2UM4VjWT/bfjmkHc1UtuDfW+mUJh6Yem3SFEKt71ykle9vhv9nnLulShIf
6GvEoXSA+43+9GP4ryoZp7RqVufXUxXufaF2KWbiWH7iZVNvLzVHtewNbfOeQYVg
4TR/KExbxJzaYzqE3I+Cly5ptK7sfJmgRYIFvpoDQGI6PyZesbAMiaRFpQFjFI+s
q6KYnt2JPlLViVFBX9k7fj22mHjDcATiV5ktW7FE47FQsPpTSEVvgzatudh2nIGi
v9IWlz2oiPDYoyyN7kohXTqye/+SIYmDNPx3JDBH4Yb7Bq0Fk00NkIzUD4dH1btZ
qV6jTbgBoxhROlcW3Pn9Sl1i9mv/8dfL82Gf8wGDPtcH7aV7kJaXvR9AqHkipL6z
HECWJW9t5qfwbmvc250yY3K9GTwhdG+doCKg30RBm4xBkI7X0f2XZhFMIUE12+Cm
hrfXjFc94eJHcggJqr9xzUCk/bAmISglZY34jdpiELHy1/r6fbz+z+RLVoyUMva5
RRJ0qXvl4aHPVr7CyN0IIziAS2UIRGDCbKmcNhsSC1iSyXuTgiIj04SzGOysjM8F
3bR/tHS8LiBCyoUU7yAShAQqc7s9YXmRRfJA2E5I/LnWV0Fqnm4KoUQfw4k1CBfN
6qzdYbHqnp3U/YpnYXDmtOilyDQQrANZvBqEX38NZd19wJQAVoOJK80DStgsV6e3
As5N1KPcAxcxH0RPtQuQ7jDMDAO6U4NHwY3rgNAbKKh7S+6+FN2UuKfpBDCLcYfL
h1wn5jAYRmAEsDpzzk0RKYKIjS+XABB1CEoCTBd5U2vVyAnu5uHpL/lFCQsPg2ld
8zDW2mLZ0F6moUF6YkPyL5Ge4G1YuNhRdpvnMnPZ4cyI4z/a9YrBw+noHtXR8iFu
Vp7sfdYnOQjghdANkQyNtxm58j7Cag0AWWCT3vfzZ3IalEN3i6FAgJcAZXZ1mWow
rKoJsBcL4fMdRuoRMIusGQjJrczwNJ+jihzv04DfGFhxWeOGOX8UHHdWakonROeh
ctRUekDK8ycclaJUoyzX0916lu16a0D07mJT9qiZIkiUtG2LPSjkVL/46j+bz9GC
0Yf3o/kwCDFI1V5qYom5cnyvMObAfoYc3DdZz32ncqagLM3m7kLoOYaD+f9dzxpD
b9d1E5cebrXs+ZQAdhE/H7PEuj/mLFYUWmQbvXJ4FYo9zAem+yijulf5JJUY7WSK
dXJWM8n7vbdKjrt3bwIdR1eeZwEA9ls/tOefcmfN/SOopJbLco1gXMGJS3I4elkW
eEg7vt2idKXZDgRYQkmN6oqmilTKfYtukUKtqy6zsUHZZgxsvMyH2Rsc/ijU/Rhb
K0O6dmsDsZZw6orJsfeDoWVAhRZMtwu4lA4+bSOP9sxDyycx4j7AKtntpFSyHD5I
D/Jp3hpDSkUZHCjTxTJo85Gfn7W32nC/xv3Lp5WX8SMWvzK8X6hVfkctOSYPp5wV
2q1d+1QZJ+fwOo0CsY/Zcxp8zoXXATjSKqje9m+hQEBm+JkhWxADp2UrbdM+VLF5
yjtFsjfhRcokaK8rlU35MUJRcuEhfNGHqeLqtOoWY4xP0h8DkanmXlMd/r0nBjk4
/xookGg5AbPdOCqeYo2CqVDw/xU/DOxebF6xtNb03IzzNkl5ZqRn9YPwRXVS2vfS
eGSqqWUhjKGuYkb7YbwPEvyvzasp9283iNsC9+s2uJEsEiLY3eoskXkcFXLuJ5Py
pVvo2vMb6q0sEXfAv6YWfsffNPeUr+3I8EzFNVXR+L88tp9ZHe8N7HDpmXpBGVby
b6jp6bXh5hD6ZkbCNa+KMN5Kluu09LPVgkknovYs/Ckp8N3VI5kMIOkaTi10h9/q
E2SG/TXEEgGXO7h6fqeAa/NVK2hOaIdv5is31oTpX2B04cN3s9V1r7En/mEtRW+E
kzRHe3AWRMglrEdpXEKHcSQuHQTBuyRF8dKwLyLNjoN06HFi8ngu28gZjYMLmlXd
s5lUNO3cPmvglsBLMXnOaRs3jkwsMCfiTxzxZSv8RaRGwZY+WuIPqfcdVfGgTX6L
qieqBAw2PJ9X+dLNidnRXAGvIYrPydnzUJlVmhlXbWQbRDu/QC+IhIIUNd7KGqFb
/stiyWYyE+QJ/NswLapCmeY14KcRyuYMbdCgAhrNhTR0PBu5OjfKq2csWK+jiUb8
ba4h84oGrkLt7jZDAKZAcoJln+RHLyhFFK1Uz+BYaOeDMCMz5UaPrpn6EGNRvhGW
bu7dI/2ONEkHp3Klk9zja3Of4qTi/oN88mJL7JTtZGK9RtTguoe/qRU35WsR7jsj
ScPdC1oAZ4x9wtkNCY3p2b3SOyriB0vjMpVsy729TukAbo6LiVRlZPL3avS7oj75
/86cMD+iIdnmzB/ZeBy2lfuH5lx9LIkoCCKHvOexBFB7BkWbNIpO/48jRjUCS+Dk
WfDeZrlu6Jy+YF8W+RhHOqqMXKYzo9Ec3eU5S341Bq+zuK8j4VfwK3kZMkE31Hg6
BYnJjUjuO7Owko0xC8tt3PdJXXCJYq2sxKXcM4So2Ezc5P0SaefqF0c8fuG9N6mr
gmoR8BAPN9DkF7sY2JQdqF91/YU84UMoEQAOCemdk66nStQJ3nF3ky2OPrHoxv6F
CWhVJtA41ja+eJUzc99Jla4gqSaq6IjiGDJ26JVs4qku9q1exdqIX8WSNF8seU/5
FNj+BiTZhZ7R+FDSLGKG1wN5P5fMZw7udQ55Y5rmbF/tHvquIFbc0aIKeEHUu0Jd
kxGn0EEi26o8tVSpqHW4hoCB03utaGBhV5qpZufwwar0Ah7x/BpLkEiUaKZNjJzv
nIUPf7Ld1nlBTbCxCtfw81v3JZSlM+WaBbd1pwUi30bQLGLVkH3s/9czmdCKvxJL
JcsGuQpmeIS9cggjNphcPqMNsw470V150V2Im0LpOklB+IhLSI/Fi4FajZ3T05Wv
qA0nS/7sHTBMuhsKgVnTVK/QJNEHlFeJ8q2pV/DK4NAr+SrTZ3ZyYPg57DyUDa9S
bVX9tFjf4mLR0BoosqfjMz4yOq/nGzHlNi0VYez5SM0NUT/UH0NIInNUdVQ8NmIY
MyKRbuan9BBDrEphbXbFXSBkJEezYg5BgC2kt0DqyFswzmWwor2aQVWkAjf8cBsR
ysDYw6XqUUVSk5GnFX4nzXT+jimlo7mMabtFnEw6EEr967WW/bJhuL1cTZQJ0sZV
H6jA4tqH7v/X6n/AZXaQoZGcBNggwJFvivAPy6oG+ctij8/AQR4dyI3yLnZCuxAr
MUF+jfn2ZUTINQ4gK8tHWCMMB2AIw331/QqeNPJJaMq6p6bDlAIdFRczSkv70h6K
37mYNsjI2knuIf8kEyDWp48IpZOzAT6ccRwGnItWBxJ3rwsJylUnxAgGbxv0flzK
ZVlunpplcMl9J9gohu08J4xL35PFqEPpxzxV9ke0CUFxNYNHVqHZ/OaHSe1B3I8e
6cK5yygUU7tSXOb6lbH4aXer9J5qaT5AgoDhmqaFd+lJ69mMH3+YF9O8Zey0NoR7
FKhHCI9pXgFhOxp0ni5HfjVBdeNRIeeCEyLTyX7zHcSy6ykJib0gtsSaZLPg7TaK
EMlAK3+in6SWmtUERDUwOhbMRJW8Y+GL46kX703loIit5EDUuSoY3nIP5Z8nxWot
/HMb8BlF8l4HjLCVXQ3RkRf1MmHLYnapW2afhjvHkTvxqptdP+Loxd0HQnjYeCgj
a/AvJzYVY0Npt+D2DB/KvM8p0xWo4bc8uNBqkvl5LN+94WfOB/nKA/Nk8nkD7FkM
kNKjGEcaRnQPHujIcXq9UTA0B3UFqYzbOVLcxdDUK1JDR9oyrtWY5IjuMimUksvj
30m/l3p0CzEodNWrrrAeslgC88BjnTKGhObaiDML6EPsCluLxnCRNKh6c+a0FZlw
yi97lkN05QPRKL6gyVoOMJA/ConHMhtMkxGxqgqRewWQflk6RwraPLjBrQ6CTbGv
bzdJfa2P7RmaXg8vE0fj3f6mLS8u4TrdiMzYz2E8sHtyE/+fMLVrf7jAp/mFM4Uk
yHwN3X4K7tUpO+TG3kpjhIVIdLxINxb6ubzQg9p+DHybMARcnfgzxLhJKz+aHuDq
PwHwORLwRnXWkbnHAZfLCjySHEUgbte/YxPUlzV+LtfuKhHdtEqlcRUli1RwmvV7
TuEhHbObUnqZGlieNTi8/ykwbI8RRP8RuHEe1jliSQFR3uGA4puEXVbnH3OIr+40
GbX1bbLHsg3ogiWCmwRzJvVmtSXq8QxVCA4tMiDbcE1WZIYv3T64LAiTWOeuVdVH
zNv1HnzrOWJEl9rC90MN/K07VW3M2WbbQmnXctdqvR25otr0UeGvFEJH80jtCm9s
dLjNkQSI4rDNtjQHoVMTZTI4KNx6Q9BYG2VO3zJn97PIoHpQUQsXhP5mepQARbR5
rDy64sTK7H3y6zY74jpnIZ2Zas8uzGEHm6u9Bq/57dK9W9JsKkI4YHd1bkt9Q+Gn
8uH43i5lwkKzAiIxfcwxCB7wU8804ebdarXj4jYk51UXXjWwaLrjq8wv9ZuckU1T
06Y6+COjAfjYMY7LhoyUmVmygkHXS35zYdbRpVTSN2fhV2LQsfO6xYhz4gK2OUZe
U9p3wr8ITgE8tRcgZdgqiyPKZ11gQEu8l9+UOByhUPyPOdB8sfsYwZVlr8gpdlrS
zlpn7wptYPDt3s16DCr9S7rVDqkz/ja66uadSbUkDpFw8RoDa33yxYgc8z1JMxBi
UvncAv8IE0uayYIwC6e8Dnz2SBRCXq0GHY0qjicuCd1SKwlx537raLz13BsSkqKc
/VMH+1yhPnwQhTQVAnyeG5S9Zv28qt+NbPx0WKcD/cTx7PtRDMB6vWVIGrx+hNms
LjysdBhHvUbKXhlISx24vqJL2g4aKIt/9EQnQmIYgmbipb1cwJ+ufNONNvOeWpSV
5/XXVsO5XeaT7F4Sz5U2yrCM6UNugHkRrwC6/uA0WhzvKzlA42HagTH84jQOpunE
6/ZeammbZ5I1LDSvkara04o/93lmwF4qaaouXqL4DrEgkBQH5p/+N3zkPdbIXGvf
`protect END_PROTECTED
