`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SCbuO5Jhww34rd6PJckspZZNtCYJt5KuPA/FjClW4WTEXP2Gvona39Vj3JjsGu58
Hol9OLAaUD+562gGjzzQKk0BGih9vN3XD68rV1pLzAcV90lWI02HtH/HUtqmtoNV
o3KjCWKhJ+qCnpDg+KhTIM75p2V/qH/pNfmKOCS2lhHsPia61d161yvDTX0bY0hP
x78/1xqq8xsfbjxqaS5KaJEW2uQyV3VJ3l57fJsEFsdyFCWcKRE8hBsfXL2MLLNQ
8M5qUDFCq6IH/5jRlT07K0tvQQ8+3OOv/RJppY1LYnSMBVJYeWQF4ibaza5LUGtM
zhsaDwVqsUkZ1W34IuCU2RAtgvFhZNBYDG5OGSsuC2H2AL4dU2doaVqET20JluwQ
m0Qiu0/5W8dItewNEXpNK3tg8vvNbhTK2bUa674iVdV2jfQdG2Yk33BA3p2mXz52
1xNozHFazBF5owOiD9knvsMcaMtJfQJW1tvwW5lzTdpS383ACgcEV9lQSU5Q/a3u
`protect END_PROTECTED
