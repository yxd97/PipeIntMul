`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Q6yfSSeqffPaGOKf4qRUpq0GKusaVlh2e9aQXeemUh+1DwXxMpvatdU4JywbGZQ
NM7UhTgNx8NVeZisbRSLvr05oWxEGxAQUmukzmm2oFo4DXToR6faq5/dWoiGMy0e
bL6Pvz66rt1UNZI5kDVwMUkpCN7dWTfepln368tyJxCnbxgL5IRpxiTO5e6XcZn1
kTKDqNZJjiOb2cFWDPvGlLs4+OiLd8L4cqbPKD/O1aXPbYYplK8uqKaZKpP7Cyq+
ZpXgflHtx5lzzRgyGNJ1QWooS0SjlDbArQdgG4ye5AELDoxTvSJwVOgUC87bpxu3
gDvcTr+gIu1bQXKH+fN7QdlP/WfFr93RFWygH0EBOJW82WuulRzRuFnt1f3w8eIl
d4ZCPu+PhQtu64D6UQBymecOdh8bGUvht7s4b1Z8KFtPwidgABgsOP1k/VWTjdgI
lgk+kEywKuUL1xO9wf3jAdTAUIDRoS/L4ku2LJUaeuXhveylL5EyjsRS1e211YZc
HhDwJGakoHrfCK3a5QvgpoaEMD0jzSwo0XlpeBkBMHe0tTXNzNOgeZwQ4sGJHgMG
Up5/TXqVJWTD93nfiSih1hZ65wTZ6Ah7uvthrlP4OWLgjkzmha3oO9OW165t27Jv
VN9+VX0czsv3rB7ah5fPthPnbQyC9FKkUV5zsIitoHaUxwZaFMsdOBcQwgUCklZE
9XSt3T4EPQXDZ8F9ZVE2OAQ2EKbvtuFQgI5t/MEiEWlgvyF+ZfbbHTC2AQbiC7u5
wxxUmPnH//x9TJQbndM2WlgxTBjgbLJPiLU36h47aBgerroha9vq5SmOQejeW0k6
4+AxSehxZFC1bqwHpICkdw==
`protect END_PROTECTED
