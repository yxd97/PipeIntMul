`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bLZviyIbJbd6thBvgwwkxm/re1J2rHvK33Bj2SvhRIGaYrb4DQu0VfEZpjpNp4wG
gG8CJIrnr5ujnnkPm2S3R7v7icIO6dY6G/SQ1cAP7QG7QiiUtAStfGOk9Yt542pe
gd68ShaAW1lXN5qqUloka45EW5NcL8XXD8qZfFvMv/6+01jmcF/2/IvYV5MV/YO1
HJmQqkkasLPd9GUEosLersP8HiwtmfgNMUDnaptcyA16jHayQl75P3J3PR7pGpis
kwFbB16Z9WrWcd8ggAHWeh/xCFxHAcEDAMEjC1QmuD6Z+VcR0ngILZHS8YkLhMFn
WE2mCR7n+gTvCAsuK0lsyvD3AA1PNBYM9ro88DdYH2AezzRjDmHx5af0iosEDHo8
FnlHKUW0Qe09S5vA89suNIMfdXzxvnCyktaKW/InOXP1Ac+tgK5SqKAdyhb6BIIh
q0euhuCIGAVwEVSXCsAnplCVb+4YzL+MZf96LEL1FmgxlbHPKbDDgW1yl15q51tP
OiuftEt07PjVgC8t+2zM4BbCU1UciuZdPeUEFLlLxjNp+dj1kVhfoBNRbGSRklEv
JRnbPbMnnK9Tcv5NNQSxiK6zoYAdt8P4I5zoyTz19JYElvZ2F8fhq0+A/VdwT7ir
0Nxs/jf1DiU9FaRC4WCXnuUuj7qJJtlhGEGVIBVW7rn127qTHbD3biV0Uu0IH3g/
B1uOETcRyFccdxa17BLZoPYmYEZk/7SmwN8ox9siFx1hd8xs3c4A8f/DYa/TuhSb
JCD0fWxsus9EShKVI7hIMikj6qQX421Kv5vuaJ3sYE8vM4q1fvqikfrqjrrZsV4X
ALmQajbMM17ILbFSo+zDwlt3tC1ls/KJDYA+XtLOrY/Grj2/oRNQmIKgZfXNveDZ
7FccxcM3U9HN5O2hb6fROqy7CcEXji2nfu1YZV22lFc/598bIfMPChQay4P0o05W
R1S8qYmBEPFGv5L/4sSeRxNXMwoQ5eUpsgSD00a8n5N3OPCDgY0oTOP2qM98btIY
`protect END_PROTECTED
