`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wOb9vSiox1TyK3WHGhCOumplwOMFpbbmIt9zafJ0CsqeYaUyTAjRF1NI+WUo1k/P
lei8A8Ahy7skmb3oq2PJvXbNaoFHizxShKxo6FBVs/gIN6ObQmz87NusvJoXlwxZ
5HeYyUx7rH73LYLSAtBeK39BKClM96PnaSrXVjtJJoJ44ZpaOMSNvJKku+8UtruJ
M9uocbmlaeCWvxdCQV9S1B5XOw5nY8pn0R/4MKyiD7/OS8UL10UuD531aXaBqLNq
fToiRRlnm/+9rqydAqFgzT42OdggSjXnZQuP2O71oqc3I2djw+6a9S3WOWRImBQR
Ke+4vNhuZfrv6irKSbPak3uB22Z7o1ZTLjtCd2TWblHVfIO7xvp61XzbT9ToK+Gp
74ZWBuOEZ2OmS4OHvri4UcBztqTQUP6Y/EZiicUBOrahl/8e2T4p+buc3XHzyOvN
qyJF1jPh1EgvHutOWp/BiLGMa9baBCVPZTcHN0Yh0h6Epa9Bhu42j0/hSNORsiuM
Q42EjqoqEeMVfb6nOHg3z/worpgqadAfvOYeA4mzQHVfMdXEkCMr6yIQjIbTIdq2
FyXcMKTWyZ2IFh9/EVd72ldLrEcShkpKJuOM05kCm6Df+pGJ0/Y3KSylc/9+7Y1T
TUON33h+64dF/GOllytbdw==
`protect END_PROTECTED
