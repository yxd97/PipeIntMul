`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GmnxFTUfbxsZCqsmJtzqYtCpYxIYNCTMPVuFij/0aa4twQ5cSIKzSUO6+dZWZIHc
817Yvafuznbt2s+kb+K1T/WyB4WvFgdtw3kW6o0Kua4QMt4XiHtjmAGLptEbm5Wk
qmo6/7YD0coi+YeAv9o9MmrYdZj3hKJsQf3tgBwk3/gAsAaDfGJbdAqB9TKa0/VE
1mQBBtaLSoTZ2IsARxV6TagIzu3fatfBG/BUIwivunT6onsaVvbmKh8Akj9RQyhU
82BpDDoQMriCSFqHNM6QdkA9oFrSYuePCleIDYuOWpyToFi9CiQVjB/1tsFTfWsF
b39CGCU1micybDf1vNdoRxq196P5N5WB+UnDnS4XBw/Q6/ICvWEntKPvdaUKi2BB
FRYMP2uYRtO93kq21HZ9nEIu8NHIenlOEURXkDWP5B/XNe84tSDn1UgOZYzN5dzo
AZakpMcMQgXFMQffc+R8H/MbldfRn2p2uPxr6lskKmdFVb6OeoC6ZZ38RzHohq4Y
1q0PpVboAikBgv5ZelJLYU8YFxbw0du2TdrcZfZmxOTUyPXcRErzott0DGH5trKE
C9bXTCE2rP8u+YLK61EDzMTBpkDTpmxNnhp/HOtJZWKPTve+qyCymJvd89ELgLz5
Ypixw3pbXyaxFeQNxKUMAw==
`protect END_PROTECTED
