`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WezGIRZAVz9hR5xrWQc2bf74fKsa5WaF+zk8vK4pipnUgoQ5yRqlF5JUcl7uMcvG
ZpXCjxiEZsFRPPgANU6csqF7/8oyRdXq+hBE1R29KOAdBD6dUSRg5T8WKEKywNC2
VoU9hssHueHJHx8k+8YH0HPfpePml7qyaYLkF7whCJ9mJkU6D40KgHzGNaLSu8sr
u2b9liyLd9p1IGgwiD5JBRmeOvcCP2aswSUrMmYj/R3GTZdfFFijMa26GZ2WiRf0
a/quwMOwLL1IAYBHm6PcRYvJBxpx5yAJqnprJwiz52jBFvz2fmcNFZG6+7mBytpn
Vz0qHajyG7BCxRY5Zog5eGS1gKhorPWKjd5v/OvwXl7oVWC7JYRuGdlpxMMcVOCt
hVNWVphzEXO/qfWG8BWLlqNyPbmsrDCcUm0rGvd1rFWnGRZ3t5BvaLOw5+is0dUL
4eLIrEodgTWfycvcG9iCixfeXkJkGScDwxo/K/+ZIawuBRcPU3mpJgPsHJhGwJB9
gnrp6X7mpn1mNzFqqVZhvT2pDo3/s/JlHJX3pvNHitz5C4maYcbtDiF1mDl80Pqr
0U4vBV9LyAf9aVgXlXMpCN8p6QAOPsbUXo98qS8hA9hOJTknNMTEQPcOw9hC7q3i
OIHdPRblO085LwThqcb/u2NGDlujw289Hz0oGUSaqzuxnjn4yzWqugQjtWJNXGbG
lqfYnV5orOyARNzGb61dMA==
`protect END_PROTECTED
