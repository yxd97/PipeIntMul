`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnDxwNyvEv+yF3KRWEoE0ez3bSvBrhFGIMwX2xq3krMSd7phwB89iYelC79gOty6
c2FXHzpN4s4+yQQZ3gS16cbeNqHuPpaMycxspnRdVB7By6izDw1ClcUHnu9IjYqY
dbos9mV8WhOpZK0LM4Du6fZwK8VpyePa2zRU3XUneDK2t/0swzvYZnB7qUuKqoLw
l5n5fCKA40I2nSbrIjKoqMncLvEs2m4wnvXrJHgSQm9PheAIAB3RSCSgURYCEhso
VvNU19ifeiICbSE4OYe9mNDmQ4nPmPGrTFW545L9hjQIIZrHEhjx8uAKmxVxu5Xr
kvrjOG4NqwYzZQrt5Lms0xrvCOILcj2TycplsiWMTNQc2ceJ+LJkAXssaNI3pgZm
u3TSJjxkPo1rArSPEMjBixi7wEDtvCscdbz5WEMSsV+lP+BGEYF+CfYvpUWgBP38
`protect END_PROTECTED
