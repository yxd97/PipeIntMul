`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
df36kHL5mudxMkYOi8cx3cZL+AVOYmUGNzQ2lnDPpbeHSu1uvOGNH/XvknXkujOO
ntoxCr9s3Tiz4fq2FOwMp1ghoXgtWhqgbXtuy0uOMAKWKghsUDWKAxqzQWbocehb
Pc0O/aqvvyDlVxF+kD7k3qzBHpEzxN2ZtMKoqFx1YooHzehrmFb9kEjSTffcteF3
tkoYTvQGMSIqiF5oBamHCv0fr+rq8nEMo+hVYIauc0PrkUEUay2zQuZqXL542rS4
nXM1KpQvRZxvkIdjzUCmITNGP9h+E/lFic3QZJv2YTXeyWpTUk3sv0Xe3ngpl14k
QHypR6oupNTDSn4L1om7qRCas+/2IN0rfMcrMmc9qVRUw+Pyxy3KzIfnYc1PQypL
fxoF35sjqOrNKuUnZ1n1gSWKp1NSWcgCwAHD9k73+97YuIwF5uQjTHup3RiEP26g
5qiwA3Sv6/Dt7s/9B6O62+EsgP1D53PgSgLz58KWmVtvipDlX2+CQNZm7bnQec/7
zP4/Kk+cToUtfW8CDtxPIOq7Ak1O+KEwtjsvr02N7djbTD5eKaIfD8UsGu4uDRux
xqlXnxeIlFnHZYxq665SJO6FWah6OqCxzUyYVPb5ovCXSrMP6mWUUHOJisYiBQrt
h3UEyBFtUq79y4ljQ1HBT+g5ela/lnrAUgx5q8M6uSpQicv97tPL2mFDGGeIosEp
Gml84bllRo+KWWyalCITMy1/uTBLBMRxm78giANpmVF7IWJzoNdDiKCPii4XGJu1
IbvgULKaJQbiixaql1O9hx/5xvd13bdd9tVsL086uprUISawzoCqihVFKYXK3tWH
cYdYY1aMXwAuWLDzcdFWvufF+Ov78myRKpvtrra1EAqipjoec7KesA+QMk0aC22T
NtnSm2FxalR/XaVlz8p+bU8EA9MP5aXACawGUAR4WQalY6lq5PRpHJXVQCWsNWVQ
J7MulKmT4xxSpvlvHS805R67msfCJRds+3EvKy/h7XyH1b3cB8lD2aDUYvrk2/0J
Lo3zCdF3eGi49zSmkj9zqT9Cudf0Y8ZKahWouTK9he13T2pwK+Y+oxp+uqNZYcnO
Gk5MnAOsRY+SZogtEVTMzt5LBa6xyPtKR+fxJakxRCoPv+ZfbWMSWHf/luPQWBGN
0eLUQ/nu3Ui9c9IoKnH2Qt90yq1zwTpjkbhGIry20+FYG647taPmRBFjRF7FFU7f
Uksrv13QJdorHVnGvmx8gGhbnRUqa21DTD00ANPjNBGznz6Ypk2w6+sHIMmAFXPI
AWbmi6Q9wKgL8BSf9/dr5wRJEg0utcEa+MES+G5z07lisXt2Jbz+9azWy3kVSMP5
zsgINfL8xj+CBU00eTNiJG8bHmVqVrbE5BtqH7N36aEH18MCADHPEqtaKXoEf0S1
6wJa5sjXVDG41AVjT6hq4ZJDqqRXW9ccjTLsu/YAeJy+xS1EjDHjzfUWLptJKnTP
aqC1q7jPOqW26EngF7hlBuBMm4O9UqHMNH19XmJD2VKClNc3CFhltAMLknu4O+gU
YNIbrB9CE/Wm9o5fMI9DygkIWnKQLeLYA2AyeDCkmjpsT3uzDq6uWq+FuhnHhU2j
Ncwi02dxPlse6PZX/hbG9g==
`protect END_PROTECTED
