`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K1UXRA/gqx3p9ZzOQtgnlOIOinivfVlHQfukmgJakia9DzN90LY1K61KWyz0riLi
E4nLpTKJlSOdHbcuBe9n/4tngUlzYu6ZCCXcodIu8k8P7LUY7pPmpfXHgyTdNetd
6O8+P8yAujolqOktPoHh++2oQKV0pCW7WcineilQ3tC5z0oeM1dP/nsE2LJcqGCP
QHlzexu/g/bAqSAuJbEjagjrJlmhRzgsMiPbou/+ku9t4RqH7ygdIXI49vl59f5k
43vZ1k5OsiZUFrk26M1sNfyxbQ5ogmVg1fZIeQLh74MIKyht9apZVwNFGl1t7rpj
kNjnOJGddugln6etBrk5Z2mYpXacsMarmMLkYJjiBSo3Z3aOySBYrk7FLse5y2AD
98HpwzpG7M5lea4J+jwbPDfm7T2x/C28NX2pDXxS7GbwdPSrdGX597HMbJDIUEyN
HGpgYBzo9djIyX0asEhNkajxxycEeyuzj3VBn1KlhZ++N90viPtK7WtBg/4wOm1Q
mI8LPVmj2gRJ61v5dwX1nQ7l+QEugCYOmxWRMJB9BK/7ojW6iUZLWdm/nBymfGLC
mwXhE2Cww4AUMRnkG4xExKXcR8SQcUtSnIv/YDPC9L/bN9Pp0u+j5CNpJHDT8aVY
qFad+BCwo/2DDUKCrU9k0yy5W7iSqCW6dQ9wvtysJNaaktQ6AoxQWIVkiiuJ5mgL
VeEZwIKBebX6yYMZitorH0/IjGJG4J1fWn2tw4gSW34=
`protect END_PROTECTED
