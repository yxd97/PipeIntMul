`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OGdYcY+BD+pboa8hv5Hx2jz5JVksURJYvu6qhOoCSTb2lKOBU1KhJExYdp7NQwNz
S1k9stg04gR5VRyYxeLdkcN37awpCcYzP3wBur3Q794Zyv+8PNoptJ8/xjqYi3o2
wu4plwsmtik20XplTBckfcKMsi6a8ffa7jy+tA3e5pxngFlLLkxRKqpbd4DKImI4
1RjVM8tEXFjJjPP9oFEqkUlZYUOJyuqGwGuZZTRSUek8MsKTlo/A/JUbJotQ/1dk
FHpVLhT0D+XF8W3pwWlp+PIYWtwK9W42R9RHtzeZQW1i5i3/Ewm50HWDcUvVq9ZT
CVn6cUAYRP1xthZq44ZrYaGEhZBQcMUTa5kwn/5QKsjnBjUuj3PJKpNWa72KYzMf
xD2VrLYWduUivrploenDu/e9f7RYaJfXv5nQJdib20dH6dsRphYAo7JkxxPUZj9w
JgjhZYYV5FzM+VLw57vDskqNNUiQvK4YjlP4r4wuNTI=
`protect END_PROTECTED
