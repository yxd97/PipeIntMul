`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euF2Y8S8wcBLAXJdrHrCP7vg7Y0V/R7JsoNRlm1nWiiWsP/rgKBl6qlcCKwMkx9j
HOh+1MtT+yvbfZVr8taeYCyekMaOdM624uDCQf4lboYdJXu2BvSc7cXwTVKwk6Fn
s0QKgp7Tf+SkwTVgLr8mLB15JU3ngtJmnpMaYMEy32Aw8Crl+6ondqkm9wjaqFAy
zmRGBAkh7blNYNvrgDnguaUxid0Yf1onaUOpJo7CCJvcTGj99Agz+jj5AABLdXP/
IhPBqsWyOzLD+18EZgZLZTK69mfuM8w1rvXHE2hzs4wMzKawMcnXSjYVW9sOa1on
YUnXtA/3e0z9ufNy4aIR1+32iBdAaGbohGX0tX1AvtTZUaNOqxvSxX99F3ke4F94
s4AZ5F/H8+2MG3tIe2BcocXehp2VYpDiH7dfkQSnOni+v3zczBUyobC4fcf6VMBX
IEEAI/HNSZH4i3lIrvBJIA==
`protect END_PROTECTED
