`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jVseyDI7r7KT2mKIA0iFRUbR3x2Gpvesu7E8dbdfsnRc1rvJSMEC1wEctC/cT1d7
CkbaZeDiKdcXKdVFWjYtZnUf231wqJ9YvYdI9nvYR71mcTZ9sUjY89DT2naQD1G0
SeSi6HtY1ols0KaDqqeOXyKInTWrbJGYi6smeiaNwnRC8KuO3Gnc7gE3mKulfvii
G1HVX0X1T/plkOi8YcJpf12DdGkEqtBfL79ml6CmL0rQJAsmQZmBzAqOrdeRcgDt
stt7eWUe5ygQYjIDgUQi1xykw+jjW4xFq6n418CaZ8H3I1vuxzKlvQzFSJ0HOsti
`protect END_PROTECTED
