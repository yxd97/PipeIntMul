`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yzz2rqIAH9YxrV5ptj4Ea8MOXiIfR/k2mj3Yru22t7rUHA//pjBhulYz0sHw0i7g
h26jNGoZsRYiEvyWwjazPRvCFv+ocbqOoPHCchn77ZMJ/GQg1+b2RpOzj0NFUtjw
0bbHygF0enIBzCKeVigWe3wkHEnTL6jTBmBoPkTuE86NBpOyV0p0iMioFjPRch4L
Bd6PeAs+3EvI9CXkYj/cS4RDe1djfZQTSsVG5M6NQNxCb4Qx0ZwTW9r7TEuKwOut
QpGdguy05oiBQ8hIUrCfup+mVtSPvvMmmojfnuNLaLC9SKQGieqcOV207Xj3k5gn
XmpEqo5jOrA9vbwL2eIwcFNrNmFfiicAaSj58QxS+6rp5eohvJuGmhgS5IpRO8vT
G/0HdauIqi/xo8Fkc7uLUHxvOWEPh44lZLVX2JXs2Y8MdoAce+Kh+iGIxNG3VJNC
kXVBV9b8gzATVBiKgTf41DcT0yzJlnzKftdbpCSxIgy2CXOKnX9kM9aRu3X08fxo
PTuxyHrp2f+rU+s7/pJUjtB3cbHP4pok6CfG9y3TwIpKrlJI7gwDDPvw3AJ9pfwk
sIdv8dfBbjgu62IS0Ny5O3IFrHpi0x7v7XJ4fqfl7vsTdQ7oJPAAx3xcR24MlLLf
Sn40Yib2o0bKVbdj75hIbr95VK1fAUSAe6HIYlDj7vCTI6YFwFHVkjc7WheAtArz
8wUnrZ4P6t3cnlaLUFEl1mNQnE4B9BxQ8KT8GH3ZQiAHDhP31u6nLOH0YQVxwOmt
Fxj/EeaXNO0Q4X7O0vPTBNQFu4EgKrgx4FQS2JATnpWfhfcxHhr9GKlWAJ/F9MeT
dmfWADK8FKQ/JcOassOfFw==
`protect END_PROTECTED
