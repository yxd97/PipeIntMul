`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yfx7YX7VYireFqPHpUTkA6jwMNSlmX5BGvR5ONspcWs9qMT5ALt6NhMjgRpp0FPJ
H219YrhKit9rUfqYmQRmteOJYBwoaymVTmZx9PkSkCsQarcfn8/yWmgLW0GBSAVV
zhFhErmbWSiqc+nKQNR6Vn6fc2Ek5O/PG0QboaRsv8n9W4HNYPbVv/9CPLHhuZMk
B8VIj6xxjqM9xfNzZotj20SC8pun3na6MfcjxtKo6LaYPBonnoRiidJmb7zsTrB/
9wUm8vArsbkY/nY/BxwhLg==
`protect END_PROTECTED
