`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QuMR08BYUyHhro8csh3jzv1AWIv+9ax6ZB5PLcMVOabVNanu9OuumCgHp4K6v2z3
4rgRy1cGe/xlXGUMy5frkfZqaBiAeDsH4ux4olxP2GK6FsPjBfHp+CFYnm1XqWxu
WrjkpXv03/Geu10SWB5lpOkFIKq5Ud3WRzHX/Z5wPaOqwcdz/AF1YJ0zTX3icp5r
Lznk/Nt2yOc45yjJT5LQKY3fIGwzlJFYGX+SaemFm7ZaekmwrybuuJ5SBh7djlMk
aiXQA7ynla1jtBEiy6UMS6rt3uv8P+BFO/JMrRvUvb6cKMn4Ycyk0MpOL8b2AzzA
ZuX0MzNTB6wpYz6GJASZv5u9o8xbi28FI0YCvcRNbwiiePb1NYplZatgDpmIzxC6
eTfYru9wfBNcUXweTMqnYbBLcZ5Jm0W6S2332EjefBI=
`protect END_PROTECTED
