`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjHBsYlfvxl6QKWXKCzSz5v2vENScHmR+E6KTOAYBVTaEPWTqmIFMnd5GtjMOTtd
xkbDDyBRZ49/+H7qE0Knmn+ZdVBmiBTD0WQSLHkPn1OlcgHp/HEYozFkHrkVOD6e
Z2ay4I9hcLrgz64Dl0u3Qrpnf//IqKc98SHXWdXXDuDFoh1/wO5YOtEIhAqyfRXA
outs+urtRprJh6G5xiV8BRHV9kGhppceHcwkxu7NShp6L3Uu86jjTSItVtfKDSrL
TO0BA6YvassAgG5KHgRDEXTyO2aXVBOHI8GHsIzNXPhHllf9GosFRMwC7qD9EMTA
92PvI3++HHLhLdIYXpQ+5wp/npzH13Fa7UPIABY9i0uJAwXeGyIqHKEziSUDjuum
MzEFBomh8nWi+3xZLimtiKW498NUWbovZnAV72fIVM9lO2XOmtQRIWyBK7GMk6HN
lqprasbK5FuFbsewLxiiI3OQaSMZ24axxHXSkNvBO9sN47YLGMgLthcjSvBozQvI
hXmXE8Juvj158scRxoeGniEpFSNdURWMrXij2IvNMP9FIqUjzAapFww2eiF+EddJ
`protect END_PROTECTED
