`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cicFGDt+w5dt5WgnYaO8p+rjsP2fm12xFHGqe3Fm6UALorj/slVNCI2+gZlebT4o
WlCR2THrMuYy5ej8m9i3Z8GS3VRYoY1s8XbgeEowKDJ+iYl7aEQ3N6r6L0ChkUGM
DNzsy8p/22LIhhbDFuFlHqhBWhnM+DuhCllP7yJar36W0EvYzbXqJtC+iAXfRbSV
9+s6bKehG6Hyk6r2q0lzjH214CQzWG3V/1/rWHRWq8rhsbjN4MPIgulI0BTj1jJn
PpkBELpKbLbgTC7+ixrg7lPD2Ck9XNF/Og8oD8tq1hgyGoDb8s2Cy4DLBhT/CKJK
d1ThAKDXtmHgxskErWFbtFQ0dbUaPURC32fYxraRJ9TFZFEsxv6kxEhSKlwQEdkX
DxoKA9amRfJrf9rLhCYUyRAQZutYuSE7zCkuHCrxtRP00skTJsxeJGv92j0epc7E
7hISu2asvSKGWzW7MQHeVZlyO++ZcJQSYcdOdb5gqz4T5p9AGDqMuzkPWfaH5hOE
niNE2ijWMvX5Aw37HV1VgMua+cfNCLlkuME+GQ6daOPjYWJtnH3/J5o9eAdOlg15
`protect END_PROTECTED
