`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+33ROlm6TNLaeaZ3ev3bTe8x0/6m73NNEtGWss86xNRgj8CeINp7UlrzgAqhnmo
dZRNne0Q3Sv38PaCRv8YICjx1D0pQ9scVqOkB0IavKkxZNuRVHXD3GFJfS1SO72/
TB9iG6Dscat6WlTtsVH12Lm/OObAiVoc2ffssWbW2x08QVMZhaoRoNArRkwVin/s
uCOItehT/i3eE8QtWfhdvnBYjvfDPh+/24/8KZExt+MZfJ4N40g+hNDtTp6NB89I
USLG5FAjGj52LnolgC/Xi6BTqXUaU3uMgl6RM2UQ8oWkqyu94FIr/jiPUASxu/gD
UD6rj+1qjMt4/V8Fkfqq88Now2wQKuXhdlRjTq5z8bPNsXQaPhHr51XCzbrQmY2O
X5cLukYJ8WEIlARYm1zimg==
`protect END_PROTECTED
