`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
reTvoV4ApUTLkFroBR/RjCVl0HDaSbp8JPeAS2uU4d9FG0JgEPHIdaPoNsKymwOv
gw6PQAeATk4SJ3bHOOlLZflKEf6q+0N+onylki2RlxVDsaC5+a53a2I1mfR3AwYg
AVZfuOT7k4O3kMuO+2d1PfWCvBDtPH01fd5vPlJpUYaCSKIJDpdqySIW9Yzve4J/
3JrKDaFkrWy+Y6WwDswtRwUyQ9qK65Ytis1EU1fRr+kcp0P/Twnr74ZZ3Jf09sak
2tH3jpLNznEx05lMhmocmXeJF0wDm1ahXUOb51LJtGtBgXjM4mhSg1klYCFbd+1m
O3Q9BaVJljG17XlesiROZlse3hAAmfiuuWMn1oK1xDvvKOWgNGAhXNfvQghrPSow
gLxy1WtuAkWLJyqtMx5ETt3fBsA++6EjNdL83DROqnqCwVPN69O6avY3Qta+bKvv
rBNkXHJWufvGgfELRZrZc7T3ehmhZ44XVamNEAvQBfmD5S9TZUWJMbNo59U+RHyn
H0Ayigzhy8bu6Ibb6NX8U5ZGXr3GoNohh4Llt2RVirkXrSVOlEC76GDfei7ZjAAo
ivhN4Lk6UzyEHVb7f7WteA==
`protect END_PROTECTED
