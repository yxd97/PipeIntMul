`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WzTZeQO8TGUjVKgDLpREoVQPCcgWgxaa/Gj52W3ww3uAlXcNcLk4CT2HaM8/ii0L
Srbf1eGmT/uM1MhjDsSivxQwW3C9n7pviYoAxQWbA/baOjQngJIsWy4yvnPvJBrJ
xWABjLF+EoBJeiB5myJh7IF261zB/q0hMU6LDlAtn8Uh4xgP1q08s7nkTaZdYV2S
fRdS3eGI5n+xSRec5S/Vcj2HXfdimD+cktLGMICxcya5M1H6cWfFftnUGP+CagMG
jgsyUAlRSBFeacY/C9pcsTU5rObNUUc6Hc2opaPJ1z3EspHi3k65DfRbEgXztoio
mOnWHTCtNC/fBG1MKbp936JJg//1fHd7jsOR+oKP3BbqXOfFjwILoUK/nbh2w+J5
ER73nvvTyVDkIXMqJGFISIVOzdAd+pFHEAq3I+nyTqVY3UP+tGolC8+rKlwhCW2j
D/3wapnd6573OC663K1ySTsFCELwYMrLSzuxtnCAzuL9KYBTeaWxL2Sa5LiF0sXR
JZryMcw7HtFhVHmWqA8Ap9w0Hsr9zwCY+md0H6Vv/KjiOuJgcpMtJmPoeaIBz681
eoKfgKpxhIQd/F9ug/cwfW7xtmQ4wniXuAUf3hXFNvfVCmgAjSVedcFv7fS7ttPu
uCZLsOTFMhMcy7+kHUX1hykH4Ip2GOLke1zT/E9gxI/R6O78GXcx/9qdKz73ALsn
FgxxVJIJOBz/lhOZ/qdOAQv3IciF7g7GpjGMJLTCbVJ5g7T84ehUstT6e1H0EQba
R7diId7Q7i8Pxn//PDWv+A==
`protect END_PROTECTED
