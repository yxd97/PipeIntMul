`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zfyh2oRh3Pk81vDnxts9Tqa4DCEyYPCU4wolKb+MyjLef+PfLBm7SYp4ntWSXEHJ
ULDaFMZYu20DawGnBR7SKEo3MKKIBvxwvMbX0vZwfYcGFpDIiGhy/F/s57QFuzGm
O5Qg+HC11fnJkW9O/krFow==
`protect END_PROTECTED
