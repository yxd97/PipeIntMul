`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l620rzGBXAp6Dn/PbvPYXa8Y6X8sEmfW2GaCMe0+eAtPCQ8c4CtdMOEd74oFbwPG
fYwGRxlXZU7YhWWvMYkgfRpevpXbBX1X4WYYNLWLQqKS3oiQcrQzLPX1p/qW8v57
F1S9tLgvA0heRV0eG9wXT3Z7d2GfwP3NxfzNVCVqANVP1VArimRWusIJlG3M+/y4
JvrY7Edlh2OdG6ni+96NTiTFLsaoatOfmFksLmlo3ARCgtFM/Es4sUVtER8rd4Dl
i+gtYEJxdnresHVr+5G5NYcet2mtTeTWmLDRxUv6MFoXihhglHv/y4pu2qqBDvXL
2/kgGOXyxFDw0/wdqzYO9tGYweczfe+DIPLaJ8oGgOhQZVGw9pRbE+qVj0jhKu3F
uPiDmlIUrnZk1d5xaQrcZvXfQMiGRNFo9tciTce4P0bUYU0tHlsmi/AelkceiZbO
T7ZNJmymzNPt3npi4p8aabNiZqy1OXUQHv3+7zDkFQxvc1/U+Lp94IWbDnqq+qyv
x8vIX5lJsKgHsMkZ4f+724DmAN65KwajHWcASRir3sHjNXjjnE5k5CXzrkVrIDzB
0bdTekMJu8cmJN5kuAGxpPjdqatWzvPR+/yMd7oSZb3jJWxlE1qPXZ5evQmqvBL4
Q+yvtpO5SLTG7O4+oOZxPr11UpG/x9t1jXoGw3dto5Zouq6oOmn8Z55QrV17+/5H
vgNfGvMKrAujMHB1HWePawsl7HA+SGNQImChxs/DU7mjsm9czdJ0L7zMgC1yUMI0
b6RkiU4CG60ecwwNUmJ7SPqWbQt9n33wWOwpfFdsYYoN4Rpq8ZyCnOgeyWal2rk6
xxrGmYdHAf35BpIx8ucl2yd9v4W2GRUzY/WDryM4omdeD3tlYnzlgM5v6AmqMqjx
QU95IfwJxUIgnU2aqL3TrYGI/6LZVfGmyUB18dpzteAMLAywy4/p4hj2LSSYV3nD
gUunNBH6yjiFMzdnM1PV92fYxV4tJW/3kh+yHMnl7BGmAx61U9r/vDeqIgCHygmj
p4c3TxiXgEBIzYzp4rkkcBl51c9a+3kHdtK1etLntm1VK1IN2eTXuhSjoC3a3qUD
hthgRnxhAlEBi4AknJxTvHhSLYSzagy/6mCBF7E+AnrfH+saxxuhrCiiIBuQ1mRN
LrXYDKhbfsIuhBpx8F2Ty2KBUNu6p118pZcvGNlqjwZ8VtrNeSGRJIPKhABMT60G
dVplI+jWlBmZklmPQW8qbOZoU/s0bBB+jNFBVfBgzDLsWbmYqizRiZuuzQ3cDdDx
gpIXd7t2bbQHaFI2nC4/XuFTHEyJCFQGt2Ze048Tjza+X0MCgyZJIncyBCizzWbY
JKWT12ieIy1dLfpWyngM5nRvNbZlssGDdGPV7C5tzq3u3NInbOCUMQ+nKUSXMEIa
FCK1SZ2EN7Si3VkQbVpWRbYniPq2knE1N+refX8evWlgaSjqHpkqcTmCM0rAaVXZ
r79hJR0eJFmJk1k5CTCcNYk5JvuJLNWlZO11YhSM0E62CwL7w4XFjNs24W06vY8D
zFfl+KJf69fBfh3cww/Te4azyMzrQ2dYYicSb+qdnmksURq+5H2qmCiSyV9Li9FC
4xm+E18C/lnt9pqjniQFvISoBtA4hXW2AZ6m3x9Is9/DqKFX+k7U7KCdl6Pg5ZWK
rzjCAu2JIJKyUj5gQgXC3uB0tlMLMblhVpm0IVGmPXO1EHENWYRFp9ZXbWjQpzms
zRW/YLxjCje7vvvQH1wq1nzHC/Ef06njqXrNaV3lFIYzPSft9gvdHVrONfTKgeEm
1OzeeDL++sw8e8r539DE7O+lMC2qzS//IumCFZ+u3KKSCr4XVHitqYLDLqu+yL4n
qTCVQeXzfpY3u1JuS7GvdaKXqaK4qB0JAHTDHY53/VVX3m1urbCKI/5UWYBSjlnj
QGj/QVlq8hmBM59g7gBwjXCd+FHDvW65EGjWa/3ZxC/6JveY/xMAJklu6TuQqsT6
9ql+T6G/HW+iS0N6RRAsaKUYry/f+NsXVo9zPODCpqlfRT97ESQfxgNd/1GfSbeb
U20iY/XWJRyQ/M4dAUNYB6KNytb2W2s9GqWOTp5Pr/qp4gPXGSdT2laNAMiwOXRJ
wNtTbDiLQTX3AGeACh6h+Dl/fx8ZWyV7HN1/hFB+58KBmUOneQ5zPpwFNhN94SsZ
zCVGSfK+cwJJy698CKG6nNo6CGqYqSdgmLPRJdArkRs6TZLLt7RWwa4/UEZ/crtr
QXZA1Eqoh2I+c/kxkWSr4PTqPALcOQ/mQSfKWhTo8cincthcmS9LapPrpWt0Njt9
3fh1FV76j72NcwYbWSaYr4EqLe+TXwC1ThZuLrGBW5OHkYt/KI1m9XrfALeP9gOy
8aAQeShHFOamAMslMsn7NGLRROmKXenCmiZiPXrFrVvmrQYX0+7jnZJLdkqRmgFk
uxPtxYaAFTgaG8vqra4XwZbbE9R2q1/6qTjhsoWghTCclgl3jcI+uzphXnr3HPMw
hkl3ZfdU7RgLyVYmE2TLG1LrQrFTP4cIaBMlYiMXpg9SiJBGt2zNusnZZQu0wk3P
tK7ImKlUW3pK2KVi9nSpctCMU5hzD+jawdpfEvg30ldPoRPK658dGGF8xoB/t+jP
DZfco/4MHRvM2X8mgsBjpXlYBReiCcnb1L7G2nimOH2o/TN7tnoWcvEWmqBYhUWe
ujM/X8C/Mpo8wck3RcslFivmcukwx1ATzOZzWEODC454+NYvj9119o3ibNZFJkGC
bkqwTm1qTuskP2Ej771f+Lk1JjdXQrKcz3dEMWPGebzgeHpTt9Ghs1tFe0SipGjo
g8wrK6tGMjK4L4CK/5LjVsdbxer8r7IC0I0YvFucbOXVEF/Zs0UntskQe9RurL8N
jEYhkazY+yz2n7hBWYCmxzDrafoTgrN83tbbZuusxMDW4IOif6ZUKNwzYw18N72z
JwLIxe1bcKu0WxVERnZ27AN29oYl3u/PFaxSkeFl9xn9716I2hHi0evmmR9ivqir
ChInKOU7moynalUuSjMq2Nn3v2gYCPfJ/rwSD31+0Rz2UIBt1iUzu+l7TV822FS2
4WbBIL6F0GZJ0B3TPHfeZf7zE5lNU55M8jzRHnbpJ6NNvUuiS7QMUz6aAMIMhePu
/1Rin48WCORhqS+i+preTsypeC5Phnl21lX5YcgO0a2kbbTY+H9RtQdvBrNQGtZn
Hl5qPqKhq96FTcMvxo6b7xcW750UJ1B9RjHO4D2NkspTgi3dTlczeGNbmaSdxFgq
JhcLvx5yy3uLNjJPXDIqL0iIWEeRrIsq9CdxSPnWa1DEc2GyS8/fwGgfHyXk1KuT
iHXhT6C7WIj2YUPl7VNUABjxIdfEc7R9PeS4r8Hy/BaQeHDbia82BV9/Nw31P8Cb
0Mcyf4/NYJM/OqDxL0C70h116n6BBJo1573dptcLFaW1hUeRYrvL5O+nvV5mydlk
+msP2VwIiZVmfmvBnfVOvGtHT9lltkAhV7b3Itw9TSH9rf2njsMpvrXfD2JZl/NB
f1JYNSlaF740WpRG1I0+HXcIAEmcB7aVIq9RddsU77TdmW/P+MPjESwBEpdq8HJ0
PQcbSp8/58jvOHg3/1DmFTJttwmPJRtw44Gs67R3oYjuF3sgcdUfPUKBEvSrRIk3
55t0DOboCUUxRel9AqU4o2h32WvI3+ztq9+C4UscZPW6JAK5L2+1GXQ5ZwtTHJLf
UqW+mgU3WlU/7U7d7F3xleCW7LAfCI3+vZ1pe/bECmJlWfm57ETKDkZphQS3LA/h
0XN4Ox4AGWaV9fpwRgmWI+/29HvnI7GxLG29zW9vkFB/pNAkRToJEMtmu4w5rNve
d+CIE9+BFllcjv/RLOfYHJQHxBwdHvT3YS9HAQra5bb9oGfNPHgWdltwO88OrGTK
8cneuxL18sSarOoB9Lf2Ovrb6lRKHMsxbBufMX9JVYQOGYmH5hSoF4/qkejy0lwa
6snmVHc4TuAk1JQCuZapEeJXHOggVGCCj3uuyZ49kMvvoyy0akxYV8TiOrJXBNQ0
EzCLwZC/sS+asSmCPp4oc8ZrL3NABvYwrvliYRcGvT+2lE1T56XBv5ArqS5+m3xY
QQBq+sw/iIU7/osEQXU9N6fQ64Ky1/kummmwbqNCiQvrWMaIo1R67I1q9DMJkYHP
mgqvmQp1+uonwZDd1RHATNMz6G1WtwgVHXeSbwucds7ZqbmHBQ0TC+VZqmAyXMVa
2qYAvj3iFcqAmfyiTbcIx7/cOYXvGnWSWNwDrG0xISWL8otELH8f7nPm6b9QzGal
zutUeP6evwAcylVLBByvz7oXfK7Mrz7StqzKjIXcQGAwTBjLBov7Fbvr1R+PDsen
Z/01d/kc9+b+BeU3dYA+VWAUdUGOHlx56QW2Ui5o3ZItJ0U+ZwhPw/2nJJ8uEQXo
CjBfexKsDp8RzecuJV3FZP1BSVrarUUy+MxV+RPMoP7GexQUJJL03gwIHABOsjbg
JgOpHP9KUCjsOH5dsIG+asrobucA9ruuIO0g95AjGSrMGUrYs/GN8sPhbhfqVxOU
3dhmbxgLCWHOCZ4H+kSJSuZwaz+tThyZ02Iu8JzVvELbHgHbe34z7/fDQo6ZcvHw
OBybsoklrCZ1rnjX7Z1IdoqRXux7h2dKzcUasSLhczH8zQqfev3mEFw2VNebiNF3
oDkE8oKqG3DkywQ6js/7FsE+9a958jo3OTdnjkGxqEz5j2B7lvbxrtRugSJyNeW3
YgZn+be7VbRah+A9wlMcnWf6Tl3mUKoQl/8uY0qFoFv0h58N6LK5eygBYSt7Y3/S
IRhyjQQXznZjhLsWBfIhaEyoIfKiCmuZdgRwNCS7THmakW9atwwf+gp+NSpGBa4P
Tnn6nbMOM9uTcuLZTiOnKS4ecbpG3pG3Isr8PLon24W3gDCRY87/kf8JeZvwgdMm
GpS8nR/RlvtGyzRpb2QcC96rtowuN+L5rNPUT+wpmdylNBfxOH8B/ZgVe7em2ag6
UtWqCcZ9N5b3HWQue9eW43/6gTHIbv2NbKl7+dfMnRbcteA9EzoQsvvbJq2WaoC1
/rXp0OkdBzezTOmaaSox+yJrscr/jg7dLjaQS6BgDL6fX4Jn3cQbIJORgjGHdaCa
i6CfjU9g18D6cEVXZVL+/EgFqGd+RBOqRjjKNuupv8G8nxaYom+Kj5ZWswQVuM1S
gDnRmI3ASOvjJkl+vdPp01lsYN28NmOOD2MX8vfHTD37mJlvZBINqIjrSFJmCb79
ixovsKSSWDP2Y5mV9nrWozpOy1Qb7pCD28AuMuU5BRVViA4gKvbm6WC8hI2Mtkfb
7Qu5CSvoXlaG0ccUWhi48jgHqq50B1iXCgcYBOsOPRMK0qCQ52t0hxf7nKy1hDZv
6KOAYaYZmler3S3+zulZ/ts25lub71Z5u8d2s24wRqUkGxbEbmNOYsCHX8p5svYq
3g0yGT60Rzl5cPzYdYDMh1mfgMzLIxDH8KyGRFjOYxudd2GnFrjxiogqjzgRrB4E
1LryaM5xC/sHNd1YRx7t7nxshq6SsgU496GSu8mPdQxZdq+S4pUn/8xLjxvdNNXY
OBa3bn+5CzlQAX++RhDkr26b61Y0sBRnW/aabCXrjRS2JmrMRg4CG7hAQTxa+o3J
vGVUNsxIlKVe7DwocbzfEBWmS6Cdc06F9r80zipmXnOtwTF2liM3BPYGzUIKAF0R
Fpt5ZcX/R8c3IIxFKNCF2TDy5qqtsIkax0TQmQ6ZPFBfOMPQoVxrbGWqZImPZXRu
/BWXQ8THo/GBAuXmVwW+tuwYwZJA6GNavw/4gK1r67adlu7QoGMScJQiwMVJzEP4
xferZ9+veXNgPdkIcK6ETjmdJa9OLS4ibVH3wc0UJuY8KFxf5TEpQubH1gNWcXtw
mCc54LLZIP1GmPkwgAT1SUHIoTYFzq4K+NcHvJn8B286BhFNrqQNOC8s/TU3aZay
P1+NW72tlhj3IFcVL/GpsTBD0tLs4xQVmmlxI7FazJ5CPS/qSy5mzE+GlbjTZ6Ot
Eo/LG4YRfbB4oyVAFja9I3jMB0/fXwnOHHUR2tkRCd4NnRkzdg89qKy1hQvLQTyw
alDc8Y82+vtToV+ymjOv7YI3KriTpdcRcPh2kHtlsLOHa2PI1z6EJ2pW+ygNmQaB
M7KPfmSxgJsWjH1ki9G9Z3DYLdK2CclNNTXzK5N0Nb4Ms1VtLqlk6Tp5yX5ZHYsU
mh7hZy5kjsmB9TZcjpNyoRlpoDmiD6Egb7q1GnZhAW/VlG5v/zehFSUiFkdb+S1g
FsazCt+Fj2zs5BIo+HG9Ly9EZ7Ixx8WZyEHSUET/sZLdNQ/5poO5jTYKrOH/bfCG
VOHHJpJMcwb6ripUbIk7jyPX3NxhQsLotFZ4ApjiQAXjbxj3Dgof/bHTHP1h5QJ4
Yb+7RyMxUNM9SZjoB9Rq+Miy8spoaruUOfOO+0oje+fKDcRxS6NBnkgbD3cNOMWF
Y+gxQRxx7CbydiB//IkDP6mjPe/jf28ulGgZ1WcpYZjtUlQvhIOyBMCCHMo02jjm
ix5oOitRAb8j+azsGahZTfAIvAGI7fu/kSluLBD/LPZ1fAm0WBVZKArD5zuJues7
j1B5YxoiOgXhMPPHRwiQhu/xlH6zRvqq6e05Z3q47ID5xhYOQcAEvWX/hvedhC5Y
784yKZ9kSSXw7NF3zEV1GHUdHyN/E0zQgritDkUOn8aHTWDxk/46nGzjDQF7C21k
riBXh7rgPXtK+WEwXtU3FiUonH0svbinF79e2uT3JMbQr1bp/r1EpnuifEVHJfN2
bzGfDLsvB1vauwM/ErqctY+OOi4A4SXdGJRw8nv3CTsr3Vf11f5bhKXPDAjKXfM4
iohzo94lam0ICe1tF8ZiQnxwWDw1s5DbvHavb4KBOzW6NCFIADpwidfkPwAdLRvQ
2iSFhBId/uzC1tuLhc63b3fApYwgSn1/sH8VQL2VM6tEZy3fIJGmeHYT8den06tE
Bz5a1pTwOdHuxmB/KAL0uPWBtrk01dj20Z/Ttyxbre9Fhp8eiR9MNtKEXKuFxq2Q
D6arcbEmfRbNQ5fI0lGBxDdlOIjKBKzHUEwbjk6VNoqzT3JQiA0VhiFLpBZuBdA/
8ZBk773jZxE1BmK5oX37AnkbBHdFPLD8ORH47ZNE0M/+4nA5HTmTEF4joPRhCEkS
uMOmKmKEXDxXdtbO8cb9jpuhvp520UoYLOzILlBhQv+jscJHVyCJFEz+StoWvtt9
qHp9JCHZGg/WvCWS3QLsdJ6dV/YQwOUnHwKiByupf1AJQavlZnf5mZ5tfHBTjO7b
C+M7GgiXGMgPI+ZqyNkarGcDmSbhpRF7om1EZxqxHivKxzXOUKkrKN4k0K+3KxTS
B8rPYFzYd80GckCvvBLbbNtjaMmP28kWv372EhzPVNfb1W2Amroy47KVCD5MI7M0
lY3b5PRBbmn+MxyjGv369im7IPgaMRfPPT32EK4EvUddr4YFUFRPkuZcN+JnTMVo
A0745g4NvDojW9jELuwox8AG2izQ+sUuCoNxauvW8Iqy2draP5Wr3RkdpGN9qOJd
HZjvO7Wyawz/80mv9JeSYzSk3Ho2e32GSJXcPu7OO4AzOyUWeXadV7Oe38lo/cqq
KkzXjX4tmuBTmPB01tytyvyDNpVa28+1UQ1dloJAp2/f+86S9+Q6WI6VqXAh7bTZ
YutrSbOyAwYHK9dtbFw3NPhqmfMu5JkVTemAZSAPCL89hRhnGAZ+Cv+Qm75aIoMi
t+S5h+/sXXLgKhLfqkDbJeVccsE0Bol7OUx5EU97fcSiM8wg1UOIo0TexDMXC65Y
thvGDbMxjaIOhneNU7prqTGDSHmLCaWkRkxa+uuvUrngb+a9T35ORa1rWjqPgoEP
bv8rfs3bSLoTntrZI6buiN/Yo6BXsZ2OF94LwktRP9zdoikcdxYjh+0BXsT7NORP
rro4rhLHrVcnl3/x7x1GmsaDBgNlhV6UK8e2FVgRqz7soOWdwzuB8Ar6EXaF1wUy
LQyfZL4bh6nuaKAsV2/72iuieIC3DwaCeZ0RkCgkqOUBLFoil09hbzgXETkByY/P
ovjjs5F9UbkU2O/oVwu3B46W/pu+hoox/m0iwwWbaqfF/ZksEJOMy22cYveFwgSp
RTV7NaFwh1U6aoMyaIbat9oJcRDEUqg18+i5WpF5t4NXC8D7rtxWBO/v3zyWCxmF
S1vj+xGA2xlKai9w+XWkDCrYugq8z944m0+/Ny8EJnGwNiqKx75BbRh52cwENV2Q
gRXVXNIjUgOvcOdLu8HaOMWNaK68kfBymXchrDKRndIQkESxsC1EzB54U/89yaLU
yi/SL4F3KXBcG0udgk0nanukgtVNm865gLxWriqM8sjL6ZyGw8IVjgKmKyfGFvoG
WseOOItQZhPWiVmsSm2emigoCcxoWvojK7qZLx90pzzi5ZXMO3aXuD9v4MdbRYtU
rjEw4c7XvZBaPbomnpCGGUCX+LFMmf151FdtKP9nQVWpJEDYoOJK3k31jPDuvVWt
/bEfuXpWv+DrIxMryggJBTIYOPKoXEme0F126QgMgRJFnKszXP96c6Y6fN7Xxqbb
iAUuiEYHjlm7i3uCZE+c6HoJfboVHTwZE5mDl/MhdUT/CnfeilKrQAh3W/jfe61F
ecu5H0usm4F0mnuGGQERuPqLyczTPM9QGPc7HO0aU/14TVZgeTXOlPxB5bEEH6IP
otAtYEDFrbid5sPM50T7TIzoWuCwrAtGwF+03+xHIKEapJLBmu8VRbqqfVFT5d1R
sPRnVZUxn9R3Sb1JL1I5zLdY8x6DyQCUTR3cR57QTfsNvXxMtZsAOkMCwlqUZK8c
j6nzrSnniZrUEfGm+hWXlSWMIJdS7zqhlGiyHyMKsuMuirm/Sz0mjHJrYPuGqLi4
GwH1PcMQHN/F/KeEUjTjZ7jEQVwsHZuBV7+rqsgPLBl1XUi65AyGLRYFzSegOiia
m8Dew7/Q/k7E2o+/f8C1IopUdcYjD7TD1F1+rS/mrwFy9qXPTXbypsxLb8MZuiOB
tM6ZfPBg4DywQoFnV+pTfPQdgOiCrPuD7sC1eu+aoAKJR/kn9FikRSgHXikz/IvV
BV5l37USNYtrUdjIjFH/+aQzQzm81gs5orpaDazUesuB/v/qlE95gfr5KTg4jIAg
F8mKd0CFmCyrfrm4hIoeKpN9m0nE4xaK/cvGkWsT+8nqfhKo/4L7SuzZo1mZg0Yt
tjO0PsIlINvBzQY0MerTkz3Hb/21Fj6fU9ObKl6Go7cEe+DGmDQ6F3dMnLZR72p8
AYniO//iRQ6Q4uhAbW21eA+VCykiNQZJhIbW5rd36o8MEjNkpxDrJP9RAQtgvAUZ
VoEfvUqDsHECsEwsoxhwenERR1pR9nSWzHcTFEP6jeQxjly7AfqfG3sAaqfKqBv7
56XLN/ks6EiTxKsFt/JG0CxtVj4Qpl5vZhUCsO8mBksuYu066OUPHnT9LKRGhTkr
K/N8dy7srrkaSJL+U5OaGA==
`protect END_PROTECTED
