`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Db3T40FdXZpfcYxlL855rBvtDM9MJIXx1oXKvGWnUSmF+DMUEbqjFqxSyRyWUDRz
png+iUNb2Wm40uMMh+zznVAmm0GeVD33kVu1DyABLa2o0WLpR1XB3rpkAlCDZca3
B6tCOyWQEmO7PyQGIjH1GMoJ/N8hsGoJZq5A0hgyQuxqhKw/In+CU43/7JBSMgi8
ulALIOkfrwwVn0yuaY/TgeWEzHeB6RWC8OF65ZHSheH8L3rKZSDHMZNYzrMqMEqt
MA7q5TvLcPhwPOeTLhwE4DL0ji4NjQn5Bd5nJQoUJeLkYd6baEjV9Ti2C6wYCHc/
Pedar0xzhqkcrifhi1QprAIm/nGZSYCilBT2P/y7NesIwtBAiGBItcrASuD5DOxm
iQtUcwm4HLrPO5AZGwuDjWAUEHpgx+47uAhRMshw7Cj5qz9cLV0Vwas7hw4Dj8yg
ktr2wMHqrOncm6tm7XUzC0KM8vvTb2e+ruEByP3dnwAVeuayhduCu7WvLpyrHqM7
Jn5yHbxr9kDDUycIv2tEkQtqhyQEmmoMPZe1kMAc+NfBUE3dm96tZ24JXmKujGc+
5F8ywT6QM7xUIeiKHZhH4Ct9Pc312PtzlDXyyjgT2djQ+K/bqVIfdHOM4HmRg2lg
XN4DLxptDAxGrUd4CkwJsvGBtuVCgBQVjanuVr1UtdPHRkkeW/PAjsQES1iKZin6
IVtjya5hK/xejmOVHE91uJEH1Pe40ukzYe5oii1/F2qOmtasBq2fzPzAWspeilLV
NMTVXQZ8tI233CsCUBNovnqYTgymYFSmnooaWmlDay3YeiA91dm0CqcNdDzqja6d
ubg/p81ltbZlYRvop5+03sOONKDuGgPIGeHrRGtBvs2iX5Cw/CUArcFyHQ3TuQUu
ANn7fx+RuY5MZGHhpRkiNFznbWtut+Eg/uWnDFDCPTcE2r0Jx3Fj8I1ImTV7amgc
T0quZSN0jyCx6XujuR0ssm+3IlrULwFUpBoawOa7so67cyU23Y2L5Hmbs/89F2vM
VPVxQ0NN2BPeV+O6IxdH6PA/8c0RcRXVkflYZo8GDW5jViCyZ8fWl+TXUE6AacdR
jKwkck7FT2DxHrSCOWa1XfcEV+RC6iKi6LdD5hnUD5jQACurts3n9eJWvBQd4OAh
46RbpTJ8oLtXSkMeQVXFnrGUCwqzQolxFJFL9ML+2T8atNSM90A+dC1v4GFeIJlS
EOZShlkLN2jwcfnVaa3ePhCrlDpffOGmu+f1Lc3eHC/JBpw9faR9O64p4roXhEPP
5jrKpHalFzW07i9ZvaPeOvncQ4C4e4Mv5QTLSyFrFhbey9+a0Mh2a8ROmu7EyoUX
+zNBD5DyivgzLXFKmNSA4mvFTnRZiymwcg0r/LKLWvdFnWoEVdtRisLXix9HW2V+
jzFvj30jlUBiaS0KK3OX6SJDD8cgbAQjfFf9YWgS1iUDwwUOQCAouxmsrwqbvWpd
6N4/tXFjoJCUL48YS5SbDmugLMbku8IC6/WyzV7PNgZ5Rs/rxy/H9ELUUP+SZzgG
blNKDG/gZK2u6R35DDZ6edNxVdA5FIWGaPA0SbT3J4niupN00PEk1rld5adlnrG1
pAn8o5djGFbiRHTaivGEzWvDUiq3QYTDR/i9VD5fvH/57fkK5GpdsRvyEZ3bMF2+
ifpDMHl9kouoYts+LKHqzoQuk3UuBYLuCYhzDKMJpHGFD48Ol+okWR+RbxoXmU16
7nV3kSDSHEyEPbDcySD/AHWyawpW1EXGY4Bw/6ciASd4A8kzcEiXUzQ/31yKIkNA
IXW/QmRvwazit33teDdILJ6szxRcw2WBaK7FC98Szx07MCgoBjV6iKyJ+m9xiRDz
cUtczyHGg9MtEM4vRcSHGkFLN8ucIsrpI5qnJBpcIkxMPBspIUR6P4hPNwAtTH2w
bEqzDOCEAT7T58T95PZfv3JC7EJfrcFPHpnGN927MpLZTWq9ZBxRRxrcwnsFt0v4
uLMnXzx8FVtbtMuHJcItbY7JOsZbz9bddGmS0zcOXhWT+A2Ra5rgkCGyx/rDD1uc
ldBEXH4UbTW+223KNmLDGkFbW1z6Pi0qLmDwNP0P/ZNAZHWuv8R2lE8yWr7EkwR/
ZM5NyGC5Ybn4cUEzOVHG/q6DOG7ye42LRknCv8rDQJ7FsnmUmhTKtF3l+NSkFYv/
TlbP+cyRiBaeWzRM7CoEcVkP0h4bLX9ETP7EKb1d2HH1vL0OQBf2vPHynY8MRxpa
IB3yLZ73usG6H7McERxmza4RWyFDHWk0Mg8jwnp15GPIOW3fLt5I0bX9nIxJj3hZ
oyi+mD/EkeJntDlxODJLV1b6XPGlDrLu/NijuLNFplP/C6JnbRMXyrTEWMkR8IyI
NuJ6qlkZoUdEIkg0cWbHhLTEVG03RJJNf6c7/xwk9FQFzAduENLbYtNj/+nKtS4G
Zi2koCl1tJ5+dHsM7YKK/+kgnspZVKThcesKMhaSL3F0mK3LKgCUYJhYKtP+q7z3
qvXjPgGvAHExW9RhMeoW1L4HADqTW0MgtdduF+RU6C7zAlVQ6BxkgumGqrPG2XFn
oT0v+h9i79dAxS680g4IzDAS71ZMKOZYTKxirRoIYoBv6Hfe6ElUk+MuiyZxPGMB
uyoa7UgOU1vq9KVzgzZJVa7V+4VYAzMlPK+kwttGfg9MlHW9nXCPk09mIi9b2kpo
xiOoh5jmmZ8uD31+2E+Qrm/j/SEf34jX2BPl5oFXG5KsUyMkslCclkdORqhZGN1k
6tdqH9y0uDDvefmfy1I2vq6GU6nog7/re7bHZlFYeBrErXqPk/zjoxsAFqVH1hbF
2WLEL3oXZBm8v8VagvB65+nH9oD3cmz56L06ciUaWhTFAKKDdkY0OxiULjgGx1nE
d/Ffama3xHyd+tSKTX2iO9qigwGZ/045GJMTTwL5F6//KFYzFOfx1VJRnXDQeNHN
+3Et1hzVGuaOiCm3kssKHQ==
`protect END_PROTECTED
