`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M//hQvJBbhnWch3QAQELIS0E6c4z8UW8Jmk7fMj6smeEJBhtY28vLmAd4YxelO4C
jMqrb5aJMYYeHlscwJLjVNKPiE0WM3BaDB0i23kA+YqC1vql8gf+IXyzfryWnb9E
uNpmONdvAMVdEsurzKQ4ogT2dYMIa4EwtmjRuyUMrNOgLWNxP4iTMjYSkbJqvzTO
BuUZd+8jlTgF6kZI6Itmh+YVjbRth+TqKlHIoNrTHMN59SRyYdCjvRD2f3cbRrUN
g8zjaC1r0S/Ge2AcAePSXyR61Nujdu0bTtlAnm1Kcm1o2MK+328+HZBQ84c0tu8S
2FD1Mz2tTNRB+i433kUSfEw957V1lIluN7fif8zGC3P/e1cqVWe6mKrOKC8Ibp4p
TiZvvZvmyIo/WPPRbCBYPWsvqQULs03NEyQd/e7MNZ/ZhtH9+kESxQF4TrbekHD3
bon3QpP37DoBW76x/ODFPLDfofxa+72U85x/kR9+zIuHYxcedBF99QBQKJsPUMwl
mrJdPL4+Pm2QiX1geXbOvvhy45mrOpCHxUw7MJP/jOhvmDyEOYr4dPDgLaoUtpvS
20LoCSCsycLzbKOU9sqvxsasiTOVq+L86mNDMQjo2gE=
`protect END_PROTECTED
