`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ybSWaOTPIzTIL4/pKv8VAdGjYbz/5W9RXXo+peTmPtbngMdA2OnL3Q4eCDN+wqGE
5GmcSF6QwXzQN7JozEUYuBRgSxS/RJQrmfWfPAtJyTLfT7nUDlM1xTiqvLL69rsh
ekDMJbYWpqc5KnTjt8jepr6O0ZFrtPRS8YPYPKqDToQCpw8Roo3OsziG3wj53gOV
Mh0CPYPyOMkRa11lV8vM9gp9B4cgtHk2CTEJL/kv5Q6YcMZyASvAiUz2/uBAvLQw
nP7/fvyBt8hfliUQmVRgPECwToKabRoAlzjSNnWzgcL7Im1FosOuB+rDXPCwTXQT
`protect END_PROTECTED
