`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+L+zTY54vHYooI3c6nIu8ilHTCLLWlZOQrw6RQafSXmCT3eWCLlDVTe4PfU4hWe
QehRjD009QfHdoQP+ag2TxMRV901gI9wKPOPqCrlbAAMBlfANesg7jd5TAOWhd7c
QnUCMo3pll0ux1epwV+Beb1LK/lCdXTxhmReDZj+RomQLcIobPdNoJp2SF/abiaP
T3O/1Woan75MarKAKNHl+t2tMRKi9YFPNhihwox8Lt0VDI6FlpTL7ExlPieiMA3k
qelUMjsfcYDC+iFoPxXoe5KU1xXoT9hB0cqxF0o4IFkm8gGAwqquDB2cGPgc3QVK
IX2ue1Rzpdt7xzKj/CEACzvz84lU/XFNU3+ohhQjtLUHSf8KYyXXuLk2aXb025dW
nnsz+yvAuJiolE/tu3rQwWUDTDbjgLlsvboHVB1hQao4Z5W6u1W4G499yM2NFTDB
vF2pmgAEKBANxBa2r5zqhA4iWuVOheZvhJmzz7D2jmq9/VDL0lxGyUR5Y7PbXuId
`protect END_PROTECTED
