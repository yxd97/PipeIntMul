`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTYH9y4fN/sw89Vklsl3AtVmBTq5c8qOuB+ZfF4xiZTLqqS+VN012vWHCr491t1C
xa29OST5wNWXF7OMKjBAoygoGyxNs+uwkBK+QSGS5cR5IqQxT8fpOrYculp7NNqL
XHelpacvvFtSbQl0guY/ithbOVWEFm/Orhgc3ZRQx8fZwahz95mD025LwZRv1UhX
9av2nMOG0JZpQmaz5RSJHIHmrvLSKmky4VZdRPiLXek1FgTdubbJm0cfDQKONb40
ikxXPtIU33Ejyi9GoVkiv4fLkgHBH2i5bcjH5+BfT7oZ2GtxCPOSzqJ53i6SVShD
H1habSAjf7pVcp0XXPxS5g==
`protect END_PROTECTED
