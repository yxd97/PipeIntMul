`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iVDmW3W6IXLazmCAfJIu8uTBrMs53JY841oVkSm+56YxVkHJEmkoZcP17VOYZNo
/xc/suZEroAyzEKw4hb7JjEhrbK577RxECrQXcVHejr1WxXf4Qz7kx1IwdDghYTY
Ro2gB78MuxWsmB5i18OFaSpZVHg3PVGRQ2z1RAX3dy0fqzBiXYwj+aRs3mlZyTyk
MN7UXuTNgoInh/6ukvircYiZBEaTCcZa2PhMTFCOqZzTetH+XVre135myc3P/p1/
qbEdnR8NMgvndbkA9c1OY9gmhZ/Qd6nlhbjOCA5RriVF5c7foVZsrz1nI2LoLsoN
tZKJIsPtIPbARGRUKc3JyCy12hh4fNl6pDpxMXzopWQHntY72zI0bsn8jwyDzS4v
xPCNbqPD4SKWnqQIMPt8xeFNWyQYSH1G3fA1IFnHa/M=
`protect END_PROTECTED
