`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZGGqmTi5QrKhLHhs5BLyfo5ATR6aK1Yx/dTm9AtS6Cm6WqHl/c/WVtJe0L54bDh
c/6KZQlq7QdyJLhhAraWxF5r0bpWDwQWyhUYf1f2IPc0i9XXSDtnSyFyQoStEQ4V
wmLiCGkE9p6+ORYxJKPArVIkXKzr8dH+f1ZAV+Kk+gJEo22uPtev7pf9ylUAAS1J
S/Xt/BzksaA9ce7RPmMQU+L3hAO0B7pSIA8mU+cgIscaN4Rc24rdVC0RLt0n2ZWQ
YUSb2APmRrBcTvPFdx3WZp60A/7SsUs5aXyljBOo8fqJLjb0cAm5ywPr14EsAWTt
zAZqweyz+2EE/Tar/i8tsOyYRqBcKrx6nQIZOonKlmIVK6baIQXQ3deX4mgN6ee6
0nn/lnTJGSDgkg7EldmZdA==
`protect END_PROTECTED
