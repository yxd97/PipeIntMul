`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IWIpQcDXJz1Jzt11OJdZwc7oDlyIXZ8y0wPU6pyR2qtaMYKiQmmNASdbhdPu3Nyj
M/HJ0QRPwx2ITPbaKq2trC/t47prhQ6axoPzz4/uR8ibGwbUbBW6u4Av6edaL5oc
d4TVn+MyVfESnQdetceSbDO9B5XRua+PE13iDmC5EH88CGbREoeZIbHoJoGcPM09
8YcDMEa7s3I4eBoT6srM00JjDums9mBYhM1isdmR8Vp3BbOsvFgXeEqlV9QEf/yZ
QotMTvMBWEHXdlFRgN0UgA==
`protect END_PROTECTED
