`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Ljr/bGtpkrtCZYYNAe19c4w2ZEgjqX56r9oOm/OABN3R0h91JKvHeV8K37vpPpX
iXMvNmPd/Vr+83sf4MEedCH2GsBOvMm+CiVZ9sHy47y3f4ZKpotVZfPaKYKnDPnP
EPXlOxpU5PRgt4kfypXqBXLeMgpVLOZZxRU7g18P4QXSD205Or2aX+mBb+fs22nT
RTSdozs43cILC+i2e/nSX/3kdPcO6if/IyFlOcHRAnhdNOPS0NKUAjvIoHBvgC5O
wLCHBp/ZqkDnW++/SNC1/VnaGaMv2nqnaUQ0s/MBNHp9NPSX/wiFyrvkZQeHlgRB
x6fDWXYjE8jq+AFO0yQTUg3bW3GptGXM0/5rf8bWtEvSP0VzoMW6Anj8sPJcNVDI
ZdTdt1ZcIf0IK9JYav8my2z/Jco4eYOA7TloPotinhePXI5fl/Z57N9k6Mn5Us8o
gq2FuwM1KjSOTq4LXkVPvnhAV8QZ/U2pYIOSF17wY5d/Uab3fRN+khuMCNM3nLWh
dUExkRhCzH73vI1AiJW8RZEYmCIjm4XwzGmBtiIAXsCEL58nzVbsMas2HPfbw4vp
nh8YQC0ZK8bA/SgmWo/NFG2nsbNtzQGcFMkR1yqDato=
`protect END_PROTECTED
