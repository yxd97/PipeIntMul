`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6iVB+q8aP5gqLV6Hi169EWiHBRUiNMt90+IJ+YotwVYTyoBgG+0mnBpWL7CeCOOi
P/WxdKkVTsl0SVNn/KysY0P7glcudg1gE2oLj2cSAgY0OTCImRBh27+TjQBJ5IDA
U1smIYha/F47g7wwAFXsRrP4WGNj/QLIGTb9fsRVxlGd4S6vP/hgloBDUnB6A4jG
h/YLPVmLerNershE7WqCBpnVzJKjQ4AP2fOVuIbuUfoL1O4uTZJewMGrb83bqRKO
jcczNAVy6khBMlHXF6CZUXjt1kcyp0xq5X9nmJWLCI1wDw3pwnQkIehNDvYxTTrq
d0ufkXENSCfj6qbYn217HE75QGrS9F8Ku22TbNBHXgk4Os9UuktC72/6JVUPtdNo
UwhRxdE/3mT6qO5E34FeL/ty7hwIAC6BWiAp2hkajuXf3/V7XZAFloc81TYgnfbc
`protect END_PROTECTED
