`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7sAnqHSeDxYs5AslHBG4FW1cZqUl2rwlSTo/N7zy0RQMykfs83LPQ4QsOWn3xXmy
KficjnkEdlZC0jbghDMawDZ9P9eEjHrfSu2fJSTM4Kdy13Ue+XcPCXm0z1X7N7bh
bsULKpvTvzhxCYbhQOU+uL5lB5ZURT0iib8YA9S1vOQ5ZffqSk5dLqzYkeISviF4
To2XEawyWaqNrXZSnsBQVV5upkOvCAJWmurszT2BIdjLfKNW/u3B9tG4eursZS8l
JdVDHRbKsNVbcXTmOTu/EH7TyTpa04ulblEJOulxnhZB9+4cYORAgX3mE6feiVN8
boOH4PYFpm5dbWtEDx4wukjNEzWEH4uRm6G9p/knSRXjnRvO35Ix/F1kWL163+yl
yI/iECLgtfkFOwJM/SUCr9fhy4FXJKWta4P/CBXBiYw=
`protect END_PROTECTED
