`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Szkx9rZlVEFM7wwSI+9MftEV9h4iYHIlZnJ97ONlCggE7kDDdvItLk9CS57XBKtp
QUWJu2g9XuPKYN1wWwRTv2RmkwV8ngHhCk3yOqfmf/WRrkS3XmczF+uORPKM9Tyd
e4UxHu4b6MOFKrrREvfuR92myMMGui0iXTVDIlypN6CTD9MDl051/g0Mdzc5MOW2
LCDu9IdGFNxujJbZf1WYVc3nnBpmKqteY0T6Jg9EhMInzwQZFEJA/oC1VAO18KwG
eF+db62caDBK8WtLT60EqapnZcxGMtQzOJyJZQTi554OReobrq+FZq9aNqzCbJky
apQLwIYpUUz/v4EizBP5tA15OJ4fcuKEEYzo6myE1MAVFQlPe1mMbLvTcW8ztMja
PQOzXqITAYWRK/aXHPckqqYU63r3v/+RBsmbdAhjXP/rK3IhfHe2Cblu0Bhuelr9
iBIx2cBUetoldHyCw08xbBsGx+6wlY4XUdEX26su6sQcE+7KHKUcEfnAQVbhiuAz
edGGUc0UgHn1+qM88nkkzUd531gQv8IyQwgT9xOao9bUnO7+92zt+DF0//uHY+C2
OyHconkqEXQhZ9rfJ+bM9nes+KZKmTV6+2fhm+ka0XhplTqebIzFn4odUP+PxTUg
dxA96PHYz5Y+CImk7ZlVmFcNE2NJCybZ1gQAbtGOM5C0pcEUsunaM323a2K3Hj3+
l3PpF5Va+q1et4ypC4+EA+fNAUV8mmb4LHKe/8cT7NlxDyz40qQI1KviTqUeFuTF
g1x5wSd76vYGitIdpxxwXA==
`protect END_PROTECTED
