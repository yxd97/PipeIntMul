`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2yR4wpqnruZbtKVbhKZ4//mmKIsRvXxFPbZyQoPxpfc4eqR36nesX0+FX1+IwWD
tSC39HG/+eJfzK9fLj+BbT5U1iYqkqxaNkmZkC7I5C8RmV/PevHFptlWt/98cSnp
wpMIJDRMhKV2CeF6+l7vA+UqqRvXLQD/0rFml1x3MKX4lIdZCIECYJqX0vHOdPZ1
2mfEH1tIsLdDzbbdWHs+eOAQI33kvbj3cDNvacZMAFd6XgCA1MK3dM2UQt19v/0K
dhSln0ObqVGOEA/p41SB8QN73XBSt8lOQyNdaUXrTu+NuP3JkvYZ9OzP9zIzjCp5
3jGPqigzVaLSWt0LWO8ueidgZJk4yj6+ZcyZY8nWu0Bs+B8lbVNUrSRLlcswprAR
teNHSeqhPQ7rmjS1Y5sID1yyHh8GaD7P5ZHWMRIiAItv4DFBMrOizi39IBX3DGJj
u+1XL/OBC76ztraUbHnrMaJHBSyI34rtGd9NUR3WE6+XnEXkmXo5R2J/TyDZya3d
ebVz63x4jVKRQS+nqV/CXqygfFnArHiSJNziUpa9BhxqK1xAHTHMIKIF77H+Zm8n
aDKfsvVTOlJ/tUb33NvJfcGnubBo4S1vI5djlyMzYe/sxO753hGG0/oqs4aiXZqQ
au7i8Jc3M4uv8yBGq4DIPFzDvVbYOnNoyqMVy7L74uYwKIjWR3EinbcOtoeymG/9
CpyG4JlFC4WWUgY/C6r6OGx3JvH7Ojym+ijXDQDa+cQ=
`protect END_PROTECTED
