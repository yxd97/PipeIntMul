`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j57/zIbiT5sy/UXCiGGlXvYG8qgWZnRL+zX3LMjp1o8+xj14mYV0DSO4xxtHdkAR
Dvz4gVhcO2u4tnCUE9yYCYhGwOpCxW7CmDeWiZtbWelJUYjftF8M5yJPKS25fVML
M7UjloPa6ztRJStmakbu88F0VBENAJfgk+Jb511FqZ1m5rJTNHq9KWM8Tj4tMdvs
hUNwN0vzQT6O7CiCKaRJ/BspdEgwdBnOTH3iwewPAIMU5czpRuWdDLpGVyJB2NuZ
4suswJpDWT2N31RtgwHuXrwRwE6/rqMol3PvNvY3zpv92RvnfCzaG2yjuROQzLI8
0bbgFs63RYKWFdOEqqvk3XfzdRuDidSJ0jitgYV0j3X2mmdVLzMWc1X7izBzYCz9
2WE5JhWYwmlNDK4i7UadeQYn9LwSH5sGz3AKo//48eoX2wrA2HiQXujppjcTCiXu
uUhrMnMoAnuYlJVlHcIHuQ9R0MdfYxia0v0qVUV7uLCw16Q8Y/TYg2a8EKQyTAf1
Ju1whBmAtdr1GD56uBC3rCmtBlcOROAUJVug5YUUOgt3JlOmJB4qLFQD2vOMKBko
1/Kgmi4RFIat2MwOEKjbO753fDTV+0ehyL8mgVD6aUA0my519MsElb2hJSKri7qw
RBtI1UZDEtW+e2u2TR6MKvmMt9SIISok0ES+e07FG++v/y5LjBE3Ps421yBJcoAX
s+rRD8gxyl7XEUxoRgJo0DKJ41JJLtwVXu+vuYRVWaFkfVSqr4bUelPkFWQKGeKw
Vl7xKp/sDCMfPGrRGVIYkGIfli8AdeGCw9KU/IL4lLN6OVrk6WCsvRPgZXx8BNRg
WH4972aoJ0l8iMUPzaWjQV/79sa7KD1EdGDIh+Oc0GBJ3fhzu1EE/oyOXr2Vuhm1
DSwtsqD0pZAJQE+lvJKAjYMGVZ5Go7rF7RxgBCJ3ssCf61YRw30n6R9sq1hc1YPj
l9bOjXhhqCajNb1w8QI95JDHQx0LQxR8I6bh+nmb7saLdQszVEXoOWDxxW7UrxzN
vlHtUJxAy8xcJhpg6yaLA7fijyLkE4J1wg2kZPipUAh987kHXo+okCLCw8kBOnVX
Sdz1zSMza5vk9zKZC1OjkuCE/6dPO3hLQTaYvsSIaTc=
`protect END_PROTECTED
