`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cb2RpMqPw+6AVbETwvhPHjSV4VfhzXODeHJ7Pi6V/pgTpBONriIQNtPEIMRHmmHi
57SZ7LbAya7rPeoX2R2yNYTG79PdVoWBEc1+cTxxjkkPZgyWQlu5PPp7EAb7kvHa
ydt8Wx27jPFBFyXMZy2OLkcGS6P9xIIfT9ULs0VgA0uTRbQOtX1RSitoJqnrT+cU
w62peImieHow6E28iGoMzHQGNwsgUTK2Syo9eVfwh4lOoLZmc0nKxxqKr3Py4fUk
MY5o+ynfNRI9iiuw8FcwKw/g0cIbbS37MlOXdAUuOxw=
`protect END_PROTECTED
