`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rI44hzYs9QIQLXMNT6GhU0edvE/1wlgChYO6gSuunmdTVOR7GK0H25AnTwN80aP
TMYVdt8KP6bMtlm+d6+bSAzm9UAxizeTzzsuu5eCnaYKPPbWgnuB/Mj2nqXomTZ+
3vhnIcMTabl+RH0FppIm0F/a/b0BdIG9ZHnUtsLORqqwMnQoqX1qoKB2jKhe+qMW
86r+iHwi/3x4mPWqq0OzvsSbbOMaY9kONRrhDpNKTQnOjR2rofny6eg0XofaLM1y
QFWOXePF31GUPbClg/f8Q5DFfaSJnnH8DKy2/hx9wGY+SNUsZHnrmdWGZPna6D1N
bkEnKh3hq5Utc9ZRsRsuIYkc+MZgfX6zSyS0OklAD6Jy3mTzP/8vmNRE+rwOCSZE
XZn0bP2BSdPUWEXX+121h7hXDUYTVlJcvmnKHdIU3GOagwz5woNho8yW9B9mHPU1
ZzbpSEG5bFL6PZsRCwYWXIPDELuu6qdZfsxi/GX2f8NJzVZwAYJKp4lk5LzaLfHc
o0IKcTuh+oMT7d7mWkce27SbEQzKJYvUTPR3a3MsvFX33XpVskwa0ZX3aljt0Wyn
7PntDkGNSrY1amEKBVVyx/1yRHsZNaLnOI9VCSwHHJq7zsKp/PMLzHeAq0GvrtR6
q3k47c+ibO6rnuG51V2k8IlA5skjWyPqy1NUcCY4vuBwiMvZd1RUXNLP0fo0SD+N
kGoreouXEh9qTjexJXf7HoTJHiNDtzltuORNiPu5mDGj7SgW24zx8Rx0fug7mh8I
pL/7nq8LODdPkzMxpVTqkq42TbwQ81774xJIPed1JErT685m/EHyFZoxb9km8w84
R9+1elYtG/vHRnnSxNN9E7s5rdNacIAr27Rg1vbN0S2F77cK/O2LRi3j+zfYF5Sq
k6lKX6weoNn76KBVT6xeZMr41okweJvft+/70mrga5Rw2QqjCVOO+T2yqVuUCJL3
BPltPiHs0XdaPvwT9IDZao6TaJK9sxLLHoaX07LPkFIW27SRu9caLXIOT6n+IYaD
NgnnHvLv+G+WTDQZcd5NUuMQlSa3+VujthiYmVLc0UW8mKgm+ZX9snr53QN82gm6
8BkU1BBEYS7fO78qVqpaAwDqT/BGvEJbUf5WSTMzfnLa6fpqhf/+XVWtLrfAGOMw
jGtbFeIC5q4F0ge0E97tvN9/Kjm3axe8lJ0LAfRDNnat7vFqaSAgp/Re566VsDGs
NHMGiBbDBxyXaMkDSEOW6jBz2fPlL/0TvbolXfj+VBX4FOoRzMuHv4fKIAGQWvKi
cP2M7B6iGIwDrjHJ0NCigZlLAv1j/9364K46khwzWzZ70a4z8k+YbJ9A9tz1Opqs
4lGByFOOw9Q91yNXbXmxacnXz5OQyhDrztNl21WPbnJvLRyaSmSQGf+Dp/gJBZ9q
sVzUsJtogqx7xin+H9wMgyZeecB5D7zG3cUHga1ZsFpPDvuRPGQ/4xWA+aCVY9tq
zAytbdfT1Vx2EVs35FncDzlyZkXyC+UYt243RbTJYQbotrrEd0IkKIGVus41FHnZ
uNreMbBTmhA+0FHa1/sBQeS4n0mo3A9drZ+BJqPUxF0ub9/Ho9jAL2hJqGF5sEwf
5xqhE0gVw8xnppTMHBgqSWdPe//fpoF5s47QEsmboqBSDjAoNza1LXt1cD8Diqne
D+Eod6msz06rMumaLPSqkf9mqcpqIVyyR9svtNHzA4ucNrYxwjpY7mDi86COJW0e
y0XuqyYVbCEFx8V05UbiY9FLajPvc33jFPM1un1bw4GJIgB8JTdl30EIfHMLJTPb
DTb8leP6yNgH0oKyAeuO0VxrlMHTrKfVh6Kjy0rgoOQs9qLn8nYpEp1nhT1iXDx8
SaYeI2lg3cO2LBXOrva3bome58vvHlFxXbSElGGa8PrLlYZ+QcCYfseWCyVQbNRh
ETYb+bGEbmr81UMOn+JkTfYBjDOFa4uJR7mpHQS8OIvyvmnC/FaLaVKbmWT4sz3F
8ZPpak0ID754gHE2FVRR9C8dzOCqj3PR16P0Qs0EVtg06GwCIhAF4sRk5kWR4NAZ
qVIOzNV0Fw/852bs/oA8Fe1KbMnnwGkO4E90anmvzGsxbfkw3cuC/m0mttZY401f
NIbn6aYmnPN76iaEr+rEUAoGVuK+x56YyzoJiM/IM5jvhmh8Ci7PY2NadXbstjfS
J4wlluId9eVA9yK18OyOz+xYy/xys/KzfU6cEqX/IkJWT76E2cCJIGWwqQCyEjIG
gxk/LoigHmrmPHv1swZ1Zs4lUv6c8la8i33++ID2Zo0ItziZ/BS0a1/RVtuDfFYx
swSvtO7xIZNVt/jz6mxuqd2GB9nHry3tBxIAorcuHxAexgou4MedGehJ2pe0qgQZ
QmFoGMeidIrF22+RDxaqY29xXxdOTdT6abZwqo2r4E4Qy9jY0PENMDfF3sqH9hMD
9kubk5M6mLrMDsCIyLtefKN0nw44c/3toepR0M59eQT8NEBQ6mi0IiUac4ZwXxZU
xv4mmBIxoRYPdzY0SZ1CtxtQlDqjpBJhsyrvfqF4xMaaZCOkH9vkgmUgTYEJHghO
6wXPhplSRmwDey/dtUrjTZlideP2bg6VhX2J4LLm+MuKDen2SOqfm7PdZAUD/W0h
d+Q4paFGd5yUrhOHePk8yXBEK+cEaMnMURPH9QjF7NjjK4Z5aOjNz6lNklFseTHf
PVlgYx0DaOeRf+JWiVEbEklLGgfoi4KScTPxIi93yHaFyXkY+HNGSs6pCvRXqXK0
RyDZuyo++wBvyMOx5omEPEZDSG5UqccOJSGLwjl+UAQymeRwN8VDAd7Ukop6PqOw
d6bEoal6DIq0GqyXuc3GXPdvu0FOZPRaDABgJSNM2MJRq4ntpb4DjPGbNFb0sifb
1Br3poT5BeknXOtniNg2wFadp+7cLY0GcUfVP4UyH6ppjJUnwqn6QFlShQ2rehzs
icl61SS5wL3uiCQOYvkuSqP2BdGqxV6oSEKw0gsvuZDKkQvGAazpWBL4mpENC6uN
tCM5CWK69wOXbmEDqm0B/FFZfcZt3/cI8DPRJ9z9v1G0HJzZcckKOh+6ZTnJV40y
fpWFHFINJF+uKh/7bbvaeJY9HeoxvI2MbXp964yS+CJ4GC8EodPVndELe/RHn40I
LvRTgZQTqj1WyPpOlTV9MxOoW7a8KeiS9TpcoCbCTw4Su0Wnxey7znmcnv6nVnKP
4KZB+HSD2wQxk3JKr45cAdz0K/5z9Cclw6yAXzGPeP+22PC7gM0iFvUJd7rRJ3U7
H/bv3aVLxrnckUzaKno6Bz4Dg8yOxUOp4T6EMnRQooHZ9T8y6UcY+ws/uXjyth6K
6kNCEovgnwIH/bdneeoKzgXt96KGQi3NnYH/nSTt66avgEK6vTSnsa2hvTE4iLDj
bNkZyotsR9xyMM/za0gg2rQfguS0YNlSf6HIV/m4TC68VNCgq0T1JSJqcaHmSrWy
2zJKVFvp0B4rTKKHe/KFPF7jKDQpcrUIrW8ngAaiS39pgvSv3BKW5oap7bx+XEF8
qxiNidq30RKLeyRwd0RpCOaARW3FyXnNdKnyM/O7McZGcASk79iEY9EZMSDJyb6X
eR8G/jhxk22gcgEOB9lHBi0x065JuCH5c4KBsEWQygpRLJBWvK8nws3bJNY7qIEN
eTWFRUaRc+SkjZO0PgrWPIiottnq70imccrqbdtpZmzeEXJfyy9bMEKfYM8cshyn
8KGkXstU3B/usEwWzXAd2Er4x4XIo32WxaqfpNkcSK6vmTugPubLaXEyLGyy1cSc
zTEwtYObup5ufShRY6Sk9R0o2tO+kffBhB434pZj1H7Alv/16m9I0wXLscT330T6
6MRURuG9NrBtPFeU+EONYbtp3QwR8rEue1iJuvg1lhRUvQVhMQaeONJD+f3GjZoF
SwYDcKnENiwCXuYoQ3I9yJpBvsclk4GeQVT7nJTYP1mzf9JTssHkRWPXHOw9NLG9
/UTyakFmXQu3wpfW32SxWU6aXhhpT2jpimA5iIMHTmbPJ584xwCMjGnd4Yvmy4XP
Ndp7Tubwy5xErBGGdXiI/0BK7pBpCD+O1rU8ZPJ/ZkaofjSP0ksp1ZUFuDJPTdIr
SdUBSlhODF3l0nRk2DlBLO0zLNBHGl9vhryTwIs7aDUw9iy4ljA9cTt6YdOtG4YU
6Gf/zpnH8/dY5zs9g8riS75iAYgjxjVWOsg/bEkSg186hrZRifumOQgR49LvfZLy
YagOlVPvPHcfoIJ0JGOncUSuJFc2znNyJ/uQRWqlDvJGDZmcPz98XenTJ8Y2pPOI
xJt5Q5k/3st4cv3S0It4dgNp+4esXNJb+6a8xp0Ln/OxPS4MiO/4k7g9bBt/TC73
`protect END_PROTECTED
