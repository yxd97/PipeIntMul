`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Lwbcac29Zj8ukbX1w7rTdZ/Gr8HpE9lyERYrOnYndjQdtK6pQNCdZjK262ZvtD+
QFMg4vuL+bdPanxp2jRGBhT3Nkv8kl9iip294BEPRiXIlGos3Sw7d3GN6iYtCAP3
Py2wE0yCuqvBy+ljLfzGWneGTXq8fA4FCns+8xkV37VkG1DFc4XZlqH6hwg2HOKc
bsod9Vdghps28cK379PXGZ187yWEtWkqGsMxhQbjLEcTQW2UIDs5techU7wzW4KE
2uTI4GheR0dNjCZp3W+gByiEORtOclODVLg8ng9+F95hY1rZCki4iQmW9VVKrttD
I8/4vrupk57T7J8H9k+XJV+IPExyRwIyWENwhP+OiE0nbwpooC/JJHBbic/rZTYO
ZmJ7a/6akMbD+WpwqY8cvHc4F+ED13W0Cm9zA3AOHoRrYBy7FgkmSL+MoiJaZ0G5
b68R7Y3gp/YbxpWHSazsg1noiG3xzrhJZXTKSJIKyj5CwN8MXDzoM8X2iLvpaf+j
24sO6fNul943xFjdMNH5lwrZUFYCrMZgKtt0oKOjgwiSpoliC1cCp1PaUsX88GhD
jAt+OZFIn3RdCDN6rWFRQN8hlwkF7GOWWiDn/zfZyMIxhNNlQpbWQqjQWmlGB5hj
6fFFOre0Kh9P172P9Z9GYHinzoAK58CiEjH2MLY8qVMqtktFazEKlZDZOsz1mK2/
5Dwh/fSVUNYK7j3e1VgiFpoYWLSrnRwZcCVrl+qiLRI=
`protect END_PROTECTED
