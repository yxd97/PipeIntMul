`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/hgJM6b7BSggUX2FVH8qaqsAfZBaYCodiltwPKD+ZoFpJHXfid0HO4T556D9rwP
L3rADPIR1KvdyGK3qw5a+P4T5gesjt1cq462UOxtrsXo08S7D0epaKLBEZYvp9AS
9/fcrmKxwLrfMRgl7aBEx8E6sPvPZgOlCRRYJCKEN10vovmcqaYUH17IkPHeiznm
aomAyAmbozdTYKY+0Lceq2VJw7HUwzH/iueb+54mGJSS8Fenca2L9HfHyUIJVoi+
CzMiQbP726mlWd85bCMHfrdbxNhQg0cxrtjMDY6fqC1odUEe3qSc0s3J4s0SU0vx
wvEFO6FRfzs2yTpBVlk2kEPA/vpyDncVVV9/o3KZSoQ=
`protect END_PROTECTED
