`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtKZIBshd6AgscSIrtdawau2lkEXig6GoVGMLSQT+UVzKdrBzokDw575dqksTlDB
zXdTPsMlBf64hA/c+LsT+Ahnwmi2DKwLCU3N6scjo7rPZTEWlYWizi2zvTwzkZmh
QCnMie0JrZBLcMjiGZ63QbctWfTU4aCApgJqRzejkFLglxyoewJKohhorVL6GLpz
EqvC2zStB7JyBRjpV8XUxB9H4cOJtVIZQWQf5oAWdv1t4QZq+6v6pb+2+pIGD3XA
SxOAREHe758/qrOah5vCqSeHE+05TJ/a41pSQG6PXx2zHHqwaTjksB4elQEmCVq4
4blSYjW1CC9bBjLrk+pnnLpNAIlmO6K3YF1nmoq9K6Q6dJNojTHE3wsj3QprrCyC
csJMUFpK0JVR9RNdwBxNsiZOhpGyMuIGX5NpwzS4qSPv6er69udu062EZ9Mn72Dq
UvsnUlxQ7RAU7hy4EM3DQUDFd6/lhIw4K0rTtv5w347KbI1tRoozm3eZkU23TeLe
`protect END_PROTECTED
