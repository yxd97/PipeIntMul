`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f5/YmrkX3zfDC47JK/6fj3fHwQ0Taoo1r49xce/Xq8wmvkWUzVWQlilvxfOhSn57
gity6HVE1gLJr8CLMhpEpg2PVa5vjoeZR4gElVyThbboOxSbm+kSjC6foTNyThnA
ioIzQRM3884AY4AtZK15HVXnz+NNTFD5lDeQC3bMX5v1Mz0mgdaPxadmnf2tLeLY
wR1aVx0lXObTcXElIBOycPJWLjU56C6btPU5spFSv+5CLaiYNGpyFL3NpjeFI2hW
wdDCgICFdHSag0ssX0BfMre5ugKqlTeJL8hU6radOuQoolCwm9ocQDuWb2cNVQtN
IHi9Q1hx2c0k3j4J61V85HoFZhl3+1QwoG/BY0q+OMKjoXBES75U0wPbNefKG6BW
VErA+3vxzZ9LOGDxJy3mB1fktbBKeNKZ8H3pOpi2GC37XNF8zLfYadk1BKzJrDBh
k5NknDhnt7vImIBnnCmxjzX6lSUOlI76aLFe966LheYNPord6CUBeoGfKG2kcEx7
d74MHkKTSi3RKNHj2fUSulPPb+yyy6NKx3Oz+1JxL9ktCgNdMQ5T5u6SxOsF4KMI
`protect END_PROTECTED
