`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I5r7ZSmiG183OTy5KWYDrxBbPf8wgk80f6N7eYIJu2ufxQYGNktA1nhNvp1XJ2Qt
z5335R7gjzMe9yWFSTGIQi4vspmeF6xvdGbs/KM77/TqruTKHfDY+Z4gTchN2VQp
l57OS4ES46qSSv6jErbhsSwzwPKvjflmjQw/AG4S67ElSGk7xdjbkT1QFF5rgrN0
SiBavu2Zyr+obVBz8CNj8A2TV/EKYlvXS6jfB2dvNOrqns16PyoU85bMt/F2Z56B
1Tl2WVobCPNdxgW8CvEmomQExmf5GL8t+Oi++lcnvrX25t2KxjlPreO89bWstR7H
A5mqw1FsbmlC9GovncYYZ5LzvizxngrwMSakxdQqakIBlcHwHYGwx5hQaJdwvznn
`protect END_PROTECTED
