`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6cW1sPyZbDgW0RngM369QpzbhpTtqCE9E0Ab7GOFT/KU6QxZOYlXJAoQeK0Zna+T
VnkVCJAP6ewBIUhB/5JlYLVyGuPDh6TJuWJrjLrW79YUob2mnOg4r2/UyALMEMOb
YNhCP5tUkAC8KkwiIC7PZNvWwZWi75J77gvfjGnQOlgQdN0icobIvtUlTePTXS9u
jI8jBZXK/xZE8Nn8IWTviq5KvqPgLehoRFrEidKOTv88r0TCylF+DAfCCNOJ771v
BwMq/Vs4oP0Mtd7LpHY8tpQ0dFIp5W5zjShBftadK9cwE1bjuQM0mClmUblAriSD
z7HFpe1bH8bl6FqgPhFEL38wZWWz5bOEfNqXe1yM/Wu+Oz+5NaRH3sYBrWuITtBJ
ERwpSpMxqS3MJ02YZqqNTALOPYD/FgrhEx2pSH8VCxauKkNmcZNcVMvsqsLdGhgz
`protect END_PROTECTED
