`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kTmswlk8JMav/9lWg9Ois97DSzUJMknMeGM4cE+T4szqUqJVdDbr5ZuuMtrmXwCY
qKMZYJ0mwvghKf/Rh+gegsJalsVz7l1daUIH6BwpvXzxp8hCxcG8q55/Ux2GZGfE
g7BMyMQuz4OCx1ncBb021lEj1LXc+Er7karNersRNd/Xab3U6UXxDc+VY8D5oDXS
XdkC3KLUbA64dbtwzrkJm/GWbd4B2K9CJooMBFHMhjzzbLubr7Eh2RNaft47ymD4
09y/Pjwc3YZ+VJeQflO5JIJrxHEg4oRwp4dw2DpZl2Za/FPX3AH04FrcLNNTU6tH
L/yE+2mNhgb+6RskH4iqG03pql2QgI6Z8fipH+epFsIWx72oB8I7ivPzXTLiwNiZ
R2Q8cY7cPQP7wod3ASgJw+u8eXjOUWcr7obLXINTOUFk+sn4iTbqQfXq0fHm/+Wb
g75Y721AIsv+OxhPCO9blA==
`protect END_PROTECTED
