`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WtBDcdUQ4Pceek9GOww2fOpBXyBoMG3bMbwUdVMHQoVQtsbHPQyhY0D/q68+YcXn
Qpl7QF+iKUDVFyphLvNecUDBNyhDRqj4Ig/fL+tHvCaj6d7ixLY5kpxP1XSXO2Dt
BTjlxU2jYlORVHReZk86DKRuSmxtXMOF1YwQhlfFfne90wWrWLCriQxGzMU90Nso
hTl+Q/JhxfQTfJJqx9O9IYMdC8IaX/qgx+/HvJ6s3NTUmiAUtPp71cipXQbnscMO
AZ0qnjRP4MnyiJbgKLeT1NjcUg9m01miL94atp+WWeJhnAgWx2YouwrRvs55hGky
6EOs3ibbw3skyFyVS7qAhdLGcETdgexsaKX7OtCEc5t7gi+P/WKZueqbaa5CwDqg
5oQzBi5lZRZ1ny2qyfFJNKuAtYVinO6853yyZ86GSvGOZozAhGAhtWXDwZ4I5a0o
KmPOQoz332x8eoFrDOEECSGgCzjlcyd3PfjNyzZBtls=
`protect END_PROTECTED
