`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MNc+NfKZyi/ftI5a88Qf4V6yBytdvXJ6qQxsMzWvnzH4LLVhJ+RyyCFMChuPgQvv
CFub8zbUQ1JfLH2qUPd8cj6ck0Ed6cJ1T7eREmsB/pWM4U7xOwwqGza2UjA6MGfe
g//MtZxkwKIQBk3A3bk6aMtYiGru8tVBSFhygFYndE/fqFbA2p65M7uJyFEGDtMH
+47otDvNAB62ZSmXeEKpGwWXCBtMAcDK5pr881DPi0Nq9EV017m/vrUtsyeEDH2g
NdTHScpb+2swEv96bY4ZiF3OxFMgADhfl4Xgzwer/x5GK2M3eQhDtHovOZoncjRe
cfcSVbu3TROHfHsEZRS2QkvWKhuhcP60hV21Pa/DI+l4+HFD/V6GDvE7s3iyomqv
uUJFRH4Wf9itbKPNnUjp+NV1jHGbZ1udLIBXi9hkqazDefVcofgU73oen2SEQRBU
pWm3NgozHeBr/S6VnZn+01TwCXil5jSrh8TKMeBMjhrNQU4/1EV3jBiDo1/AuMQs
+aQr3nBw0udap0SZ9WWHJvy8DbRc9xabhdq4A5LP+O1B9IHTcNwu5wxpaKLB6ayt
UlMw8V0BX6vGhXIm1cW3PMc97EMLRNa2MmgkHV44IwRmzmrPNEtuicd7kGJF9Aqp
++Okd3wUeYu+xrTqo9ceiQkZ8Qa7ysuo2FkQrNgqQFbYyfPY5R8aLR1A6rip2Obx
YqakS3GGm2HOxC2vctH6HYgCyLi27gTK2SSD3vFkzZs=
`protect END_PROTECTED
