`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmMyZZ5oqfjTSTP+lh/rO82KIbBTtjeXkZh5+u56FipGty/WtZUdms54WYcF0TXP
GpDj3ufNYSV8V0Fbd4qAUH36cSZaEnlgAchw0gLHKqHjTy6XzZ0ymbAAQiQBamZN
/1NVIy5qmY4zE8drIC41GRdHCJUujSor07vlivIuIsDH1SEi1/tgvu2CTxsrWZj8
UgvTAy+YKm2vXy3NZnEZDmer70PunLZKXqLjjJxToonuFnct6pj5G26KrbJdIWCX
Mu0q1+XbrkyMqFXEQbSN3poiO0HWWtQco5zBp1K5WCuPU98mEEI//gre1FWnlH89
Xykn1+TdY8DtpGMMjnyTMJZMl+npWQQiNiYSPbZZ1PoC1p7x16rYdseOvhiykmJ8
dP2SSBD4wNpEgUvyifR0i8vA0gDKvxbjf9oKPGUiGnwEewJ7sAOc+j4JUyzI4kMZ
hMLIeMnRnykkflxi9/0jW8MkfHhaSFdH+1r7T3UNFzZeC5Fstu+3MH1PJ+BImP39
ueJAfKQZU/DVBC6gIH7Tu6dxurQ3M061y/nWdBSjZRDGwffVLJ0T2necrZ4t1Q26
H8KEi9AVRHpHlpJkeldT+jRdExVTau5eOpWGaIG9ZgYYFCJeE1D0sKcjpVK3KnkA
I6Ts6C9pjc9LNdru+SkLG/zNiMVdwJA7Gt2/fMFegnW58COrZfSFQVR+ajQSp0Tp
NBZ8JoCzxV7UdtBuI54ogr/NjGUkFMDQJEQdiYMmrtiqp4vIWS3t4ndzAsxJEX4F
UzS+Le7NFzoG8cMZMKdb1n1RY+2aTepP/+cNGubKuVwY/yx3QvgAzAPG9Y39Kj1x
vilrz18z9OM/VH9lDcYGi87+xbESLhX3VIb2fQTiQMyc2tAzY2Nf4n1hnnks8d1R
vwM8s1UDvat4Swy0lsJdRNwjIk6HQ/KOnMwiTtzYqaUHV4g8SokeIDrJLY4LM5zC
jv3zWVA8bInngKgdta1BUjYQhRsPIGCHNKWEEWFFXIDo1eXrH6DtXh8Vygf9YckV
7FhKsNfQcEltxNl4myD3j1ly7gYoGGupwxIHgZZjBHKFRtIalfem8ujsEbNf2d3d
ufvaSQ8xBHbP1rpPjTSngeC4ppTPUov2ngSYp5wSMjlSW72wwLGCt4xUwm4xGsKi
nMOJNuQ68VNxc+Esq+/ASBFHUJTYahvd37C9JYGM2VxtJRWzuNUWzDuwNhwSNbFe
xz3G/p9KVf2+trEN8r6MxFgo3+jdSoIe9wJgf145LLrhBXFNP7YQroXYn067RoYM
hKd0XZ5v/fSrIffauXaY66dqtYyU2RGHB9yhIFs++B3s9uG8K/dIEKQt8SFqJEKC
QpB+jv7OVN6P6SUB0mOnxbG9NPhonLZgIJJkstJ93rRecfIZ4uiDVoAed6Yw8ht8
kJu+sNy8SwK2GBjvQwcQpiZwTJ13Wd7gtRnzK8GBMqRWObSPkg4LJM0BXwyG7QaG
ZJbSAaXoIogUgRYcnvq0wkhf9qOJVCFh/VpAnzkMqHUsDlsAIS+rVU2+CP0ADjH9
yoHkfNhyy9bipXQI5NYzsTN6AfRIdN83GBE98QBFraPc5MySJb6zjVpjA8dCrHqa
Rm9fM5+kcyFNcTGynl2pL2RSKKEs2bon7F/CvYCf9q9OA6v1dEwuD71i/HiNbFm1
yX+eXsuFe3Jpt30NZFGtRH+BFYJAtxv7pzr5mwOGRVwIzn+ZUu99G5AsRI8EobY/
UxdQ12EMZM+fHddbfcjpmQ0N+OeI0dEZXLfxn99u2RlZo2z2n+O0g9pKOJFVlXXZ
C3o0YgZ//N4W8PFElTcwLaTidxtqwEGzRvvJtj/nUtcj7hiuHwEJ+UoZ4gQtnR/a
iq8NUuJC1hwOL1n2ZOdvkjsKs+zbdcqGJ+vB2mAHODGGE10sIELWCjZDVMh9xx4+
UBUKU4c3MeH7tG+uRRoeoWptuEVP/KIZrsVtVrQ5M3Z9Kie3lsl+dIakvuexiIZt
/R51zTfkKqPf3tr2vZT8OKfKWo1FLwYyjI0sormuzaladNFz6UEGqxBvP3L3pGnk
puxQBnAsZKrdNHNLaiWFl9y6s6zvh7tk0Zt2TlVqQlWfMJAsScrd91TfpfM/3EYf
bMRO4im6Buq9CxggMG0ZGXv1rfs1jy0gk9Kn1CXh/qesiSKQaYZOM1GM50jwf2Ia
kYkljO22xGiUH20cc5jA5pjP9TA3edKOVWtVM0MvDdAqqemkd5a7uscWJZskDjHy
vLLFT0/WfmWDQ4FjZxVVA0az0FZrOET+jQd1kfzbSZbhLb9qYHC+wpfFxoI9pf5D
45eMYnACBMJFFEhw3H18kkun7c9nbyiH0lCI0Cj1PZOnu/4fOFBYrM9chlNfdbTu
CGLflqMpsTcgW+ZikV8Nw15S+1E6SjzJYL+UwjVf7ktyDdRacoqTeR9rVUkWuemH
5Zd3Fvxwf+Q1SOAbm8HyEDDjXYs8p9Ix3W/45rmdPj5cvRB50de8H3lahex6coVX
HvmCHGYhsRsc1P0KU0GSSS84tUiuNYTJctuCkbuW8vFYQra4WyPNYmxAQPfjRtHR
wrPpjlJGbjPA7IQ5jgqvmWXj8ay+r2I/LHNzX21jYe5RvIoG2lg4MWRvM03F60gG
SEpZlgCHXJhUbywcgM93nrqsxs7GCRw5L9Ut9KrRXJIXJ1ne40GQMdowlA605o41
VNZLVRUszcY6YTtZcznV+7Cc+9RlI4cpk3OCVjUU7MY8ytrZBdMmsf+fad+4m9ev
Wd1rMZwOx54roztotBmtswEpPu/iFEcLfTXerziLaP4KeZfrlm6OMsUdX75yX2sY
sKyWh6hWgb2XkoGEr4o9xDe99U8yL4GH5YQ08D0/FfZMLe4FGQAC97JTeeMwIJD9
fycYv2LS9QfA/4RiXPYjS6OH7/bi0Dwrj7CRRR1sTzkHwi4roSrTiatGZcoqqJmx
zUBYI9tU42mzSQBlWSo/DSVQYR1s+XiI5bFiq/Aajt8PhERdxthw+v+f7c6eFqjr
LvLSUI7Dla/Zf446njtzFt73g1F6Bc54u/N7xXJ8sPoyCUdHHxkJuXTSr7zSz4oY
IHsboo1wmBXMxmS63e9WkMBfv0MDMqLXFLRoRswNWdtpS8orLtcbXj2COJ5rktlS
TvM7JGQKGbJlAYAys7jfX8S1z4ZPVwmPSR9NbBT62CkPv4PZGznxWTL+jxV0kQbR
BSOJKFwGgz1ZqWfvRYT4u4hksB5DkWOgin80DcrSo1GTsTtUchZNpzeGV/YrU817
vQikP/wR33IkfSEUmD8Ljxww13RkWHQiXPADTTCeOU3npiU3fhRPlAl6kJCc9UMy
i+D3JufB3u24O0A3YB+kiS5TK8oXrstBTS71wgMi7ps9ZnHIV4CZYrVNkJ5k2VKY
q07mNHueTrn33lDXHHT+46ixNnJA4HZ0OjPK4Jz0UwOx8OV1lnhefJ0Iw26D4vS2
5gWc0b1LyPLXMbJP424NCPTDOfGsN3pTYEK3uw1ghbMlJWXiS5HMGyeF7dWO2IAA
Pd9U8ntCjKdy+vJh5tNIHlPGsTFzX7TGLhyBEbxyJ22KLzzqSQDUNwZl1STthJOc
yA2kKfVkBI5XZ9IzNVhghhdtVU5r7tyTx6q36vdwnMpFfzhoGBP+UnfWMKXE6y3c
3sQnCvYvYfh7sawVq4qiBPaiodpffRdtTuEjw4acQpcg1ZbONFdCurPX7RH1iX0Y
Xs2ErieMmdhkIm9Ntkgv2ZJfuIMwm6be21X7I7mp5JIuisjmO+stGqHGBnPozjum
L+qWyV6XGXPDEjRrPgh6HZARoCtagpI7nXxUzwuVccqzKzM2R6GlYyyylqQ1/yDZ
bLBCMMqnXZsB3N90EeyI07mjXBBIQkJf9tUIvZv82FLzf1nKs6kRGysW2VmKxYx3
kyX77gUj6edQCfi9N7nqQbw31IRJelgbwvDpDUF571UGaiNzwuxPULBDNs4DaRH1
G827tKxrICrbWALJ+XxhYUEoOEXiWCyvVjb0uHBEsjjY4eWYnGjJvlEvoXxl6I9V
7/iKCdsVCRZ/g88NgoRBciunYEjt/mOHv77HPc0+JgoOKJTfzNLMuOtjgMlufPEF
npIGLJ6b1B94aOyQwiZNFQ1eO0RjE6wMCSzcDJ18tRKFouJyk97Iqb3miSHppWLc
L6umMd4DKf1AoK+22urdGK1cTWmjoAeht8MVhanlhxpzbvTClfq0qYKO0HMfeCUh
InNX/K4MiVEh0mPdy5YXFg6zLStTXSbjF0nttoZhk9uytgW3bih8Z3JaRC5/GfWA
+KFQW2Leo0TchClGn2um1nG7LqCK/zkcBa7quShA84BcriLPTtESQKritmpCAe1E
pVS48KfojL0qZMwnTjgD2ferYks7g8/biwpN3NdrfsID3a7vqXNzvqQ6KpPKyjDe
PIUhKooW914NZpLOJoaVFXR/4YgYgnTNn6pI6qNHusfL3vrmhnhB8pR2hE+N0yB1
+jCOzy1Jgw3z+oRdp8dbfX/BvDO74DfI+pkjnvi6r4cYdJsTY5XF8liecEmfUkXl
iTukYG80YfekKkaslCfK51UDuGomSNpmRbzC2pyzk9y3ywsnhce6jo7HAGHHq98K
ZwPHpx/dLXFO0gZGoLZ7mCcazYDuRHW/qC+IdW3lGIdt7srZz/wNZ3TW4+BG43ep
h1XnZgEWZDhh65vJuTwiwCBN3Q1yN4/aoDOb4Ojum/OHlujPGb11CwW9+mMsGccx
Quci72YEf0RVjCo8Oane0XiUNORP6omEKps8xiYskXS00xBfTPFEK40gLw0YPtQ2
S3HutusKY/Rz8e0i3y/NnC4aue5RBuaXtw0jh7Ru/rey0e62tWGA3mUOuz6P3Rh1
aJuB7xRz+yvfoI8EoOuj/AjvLSK7UfPqc7pESnceH7ve0BNY9cgw8Y+9hw5K5rDQ
ILBJDCM0ssIeEHYKJC1meeny9Y0AtsicEausNN5RbCSFFSvWKn35xbKkB3VFgQoe
5d6VQLkuuLX6ULZUYtck14Mmk2hfFh6D2UJjKvhvdJKQ+nd4zm41+bQoOmo2k/uo
VLllvwnIkXrNaDslqw5GICZ8fGS5W+iAx0VsIEkuWUx+0equV4pbjyRvfjatqkMW
GvyWl1Vg02hbSHFSLml00Q18LJPOC4mHnjQkTJv9zOO8P0i54iuCEGDJ1xE0VuWz
PdAR4+G/TFB2QeigJV7JsUBfCKpjmhx6TKxDF96j6ZuAS+UqTXf2M04UEJWP6Awq
c0nv7/fke786JEDktFIg93YXdd4R2PFp60FvRpzTRQlw/0dvMeiGbEkp1DkmMVWc
/29cSc49T+BnZsfBIS57zf/IxvgWu9qu+smVJ4sVAbTqCyWUGx3rZqbOg3SMdNRm
NS7htY6Z0BJnlSdaE+zRB4WMEtv8T70kzkR+UYuRb2gvddlMBesaSmdt7RyeuJ89
QemvuyXBaj56YcHSgJfQupfktyxuFVavLCma3FmsjFBhwEv6iKDpAS/t1x/b55eT
X2vXjJSZCMrU4rZU/p8o98noBD+21jR8ngFHJc8n17bQaxqoQGkdpOmatTS25zOn
0s66LCaUTX2wiubt+NCY8xTmgbbqfpHJ09dw4WbhJNydzZA6ND9JNqWSpvdP+BsX
x/GabtJDoApyuP2ervmjKRPm5e1cQTJ15KPQmLIX9Dg5XdlgO1dQDgN2PGDbBdXG
qefzWW0ISU8ShwK66XgbbhHBjOAFyv5Cc0XXlVFF9t2tfnjNOeJUm9a27BIvT8V1
P8UiGGh/k2rumzbhoQv6Kn9o5yyubMyC8lbZV0pG5s+HLjLdsMIt7Mn373XyIZ0i
Issx10Bc3JQJEKLBUiuicaWgHu6I/9n/gWgTLOH1lRJqY0AXn7kB5iOYhZw3/Fae
eNk+qiIxvyyj1iKbwW57MwRPI7d2qITCVyO+dx8P4IAsK/1Sa5y6JHc+TuG/0D/n
d0X3EMgEttovg5NGlwXPHUfIW+7prH0B9peRLa1KwwRa21PxHSMiESUJ302n+yZ1
7cuK0hzGSdNKshnMM/+9c4lKNCJCwQaViiQBuVXToFdT4YB1wyW7giY0+p8MdbR1
5fZTTqI+RNlCUYExvpAOiyMmtmEI/WJEBpWRxli9YdQ0pF7zMAgEel2BasOn0bn3
JoUdvcfNOV2jsDR7vd1k4d5WK7QT+kE4m4KD56lFPGqAfwDfGyOIPVQkQvGBffit
CmblfFiINxNZANWf6T526Q6rbnpxBjH9U+0n+T49kF+8pX1JGmQsBS1EiEEUB9aC
QqtgkXHr6S1C3M7OEQonySolztjbD6CpYXeBtHnAWVh6gP378HYnlokDDaO83QE1
Fgm1gUUAr9y0uhh50tZKKFx/IKxYN1dQJlL8424k0QaD4qPOBq2DVTZqzRetck9P
3ehi9VzXFy2S6h4RFepeXTOVhW4aJ9sU8YRsSEMuTQ1dW5/D+COE57w6WhZXHdpE
DcLdyskYUAw/kx7hzGBz6+1wyvdXwhIrPZBf9/nQ+6vdStVp9TBuyAyjzfag5VSr
V8X94+VGiw0xjOVHLkNuarqJHCq+Ks05fqM1rPziWWMFeBVtEuDG1WfQi2iJc13t
n1Ib35z9u4NcvpcquVNmi/ZieqSRAf+mYEfh4la8DPD76JY2H/DxKHCA3NYUArsa
i5KxcyigBaOedQKk+sCC78rARguXQ0TpTZbO2b80ZOPNjsHRvvzWISnNsutFYUry
ExbbEOKTh4PJYCsJMaENGSFjWX0V03TmJrjpK0K+O5QpGvMuOuZsPflOF/hlot2y
rheMBuRcGUAYzlVu0y2K/tF1jviVNdXwYraH9XTHDqkqTxyIReZNk0at25NCsN9r
fzROm3aLhEWJd5jycvlPP0d9oGV39Qpt5zoYpREMqoQ83/vClGv+LfXTubR79K59
QKaIPewHXxP8FIF6Wfzukt4zKQsX5U/xsF7TloTYubBk7nP9YNkhf5dvP+cj91QB
5k7z07FMoqyuPcURafkKAFJ13XNq0PhL1Rtpu2YSApA8GTFrncJTubMI8GhRbQjg
DF5gz+RCyrAF2AToC5R8FH2PQ93vhXlszcwHm2VjJ1QmN9baOidmwyYv+z0nhzv7
QGiY0ONZ0hXWPIQmUqSKV/ekzRM+e7YpM2rhZBtdQyyMMnCZYCa5AZxVZkHuBrRW
7rGKf5eODaV/qbfnx6EDhRPiu2NgLrYsXXybUMRm43EzXHK6I1Pf7IPtyKvHtZVl
NMI6iSZYOvOdBjy0TvR0buc1ZZCrqwbyeL/LsjYXIFtr9djplVsr82fDojnx4cF/
kBY/vMv9a0aqIM2MFkgSmjVgomr+dXq2MV/zUw9J4axk8irHK2ZKrlsI1RRwROrk
zkXxHYYu12uAw9zUW+nVDqmWQJVAb04tHsVvydqzie2js9YFdC/hyTYHFO5Sym2l
1tx0zKW+OUmTO1iHsTRUKtJNXmsryx/15tSVwLq1vaQZXbue8RolavAAp28+lH/v
QTV7NV6YYbg1gX6Z7YS3jHulxa2qQ3UGZCMYvZwV7gyt2HmVST3MFDw7WnOlg+6e
w8kiMXGRTO9FqC3K7zxxR8A3ZCRS0oaB9FBnC3mRmw/Uc90MGBFKJjB0P4jD6QJo
DcgfspKmhJxDPC+HEiGVOcGd5GC0domdxeElQr+R7PGBGB1aSqFMoo2iqOC/wPn7
MbfSeKNmIrjzMWMrtCrl109Ag/XjBzTuF7X7pAimIWbwyxV0PWvXxBP9hE5wP7cg
iGoUXaI03BXb5eWa2x6XuS+Ri0PzAeJ0hKealk0351UADFXrZfN++23JNwYr5S0k
0bvANkWLR71S7b/fLEf9mriTPhi1eH8Dkaq50FYufvHO4JLc+KmdJsW2MIv1DEPy
gU9yABiCq0rn6UNhzQCZHiLeq0NOoZ6V6GnLsSk7gmZBfPl/QVtFIJqOFQgWsB+r
61kQoDeLZWyATRtvERsWdtMkcyT1nyHpz4AqOlkfccR1hE5mJGUAWkfcPDEWf6yj
yxC77GEgvEeZFrxNEd2cVTH4JZoyX3bwHge/zzVdvbWrLBHKMdLTqS1FfrJKx5XI
tJhhzMOHQg4TU3N5M/mLgKxXuZpXwBYGt79CYSgnCinzPzeQ9KwukQrcI5uV9epr
Ap1DP11YdlJ8rta/KQulZ+Y1wWvE9DrbdSn8zgQViRdm4/s64Q4OjZYYQ0Nz5vOv
8nRIInS13AebpNiqe9dA6I44w8+xXJJCbnAUrqhWX55plGaEoSDpEQu4aca9AYG3
Tn6CeP0pRZc7EUUrIP2LUX+be/geRYQGA8b4KmLXYcmutQ29LgG4xSAR+Kwe7VTU
13pu9HJ8deZ6VIcydEHekr58ENG89GnkitrRSlobEuBuQ8vU1/fbJlVfLLLBBozG
2s2fNojSYG3O3523yZQadJC5oh6ZP+yHM2+Gzyax+u9mZW6nsOu7//RFR8QfsBkD
5h7/U707XV3VHqyUBmrEWR5+NOwAWG7dXdnEjm29DcUzAsAYoz98rocsjQ+96XFU
sJuTxmCB8WljBR9YQOSpCLOswzDd6oaIVTl/JQCdKX//0hRqnIKQTDBdPQiu9YdW
Lo1z1TjEJZOn0H6+ukSbMCzLARR43VhTYN6FyDlTUJTgF7J+5N+KhdXBRGKmvMJN
4lqobQo68M/9EHO4zb0k/iyFkEJ3NAH2KGqB8HaY/vYy10ZJL2G7Jw8nHKfg8x/Q
T6OmvEyTwf8l9QXXcn+gE2xSywhFhhzixHgAOBwKKGCt6YFmGRgMusZLTZGmUGqD
UScnACZrF6zUQgWSupTpK/UsBLF95WdN+rgPHvc8/LSB/KhHI60P8x4VlUTKyEmS
tzE5wHd+sF7YuxO0/l3oOJ6Wklb1g2bsbASPIdD0vgrL7pR8DJdqePHMfIuHQNMo
xXhgzduTkacRyu7nrNsPAMdAMY++8ntnxFA4iSOC7s1wy5zqwy0d9nifDbqBTzeb
I8rsFL917l8V4gdEy8Ghy15si+PjrOrKFSCBN3jZWEPFaYM1ieizET/arZG5TVkB
kC4ZWaN4a+yG3taPKxpklNWEICSxOWoQo0M6BzpvRsowrEnzlMS1MpPTesTmbNFF
/OtoXpBPDwSBhn9+DAD9IRGPNeqfYpAUWyjnq4zR15isrxe+fM5Whd/uQ0AZiO7L
X7lzvJBOJkSgvoS65NcD8T/1ZBN9SAnFgLcV6vCNyHh2Ho/jnq9Fzwtq6YC25Bre
GNQItXmu2bUWc5nrJEXdpK3Y+U0kCKqn3xsbF6kVUs0iZHRkDDB95puiDBzpsPWI
XMF0ijesOsT5dZq0aPEyGa657GheUuEJZ7aXKuHARhVz/8zirUU3iKvVGuhUjkJy
dYnTXuiPy777lI+TEInnIk5diJstKpDDTISWpSz3QosqVfSMf/p/SxHJvkZrhklL
bewFYrtaEM7v3ZLiGcQwW8ywFZiad+/1jS/lzr9v0GlV71DcCnvFX9s3r7TU2ATn
XfaS/owRhIc7wHm/OVfT8htNGNh3+lPXhzF8waaLdJ/Vb3ndJoAt8w6lmn/2Tmr5
0+FQ3ioVziU+eovAH88W9JJnX3peKnvcyOcp7UoJZsYdTCXWKnRoH9oly1dXrYDl
bRHGxvBLLGnBwIKaByg6UnkDoTV7M1ynXnCH39KZDvEu9283/noaOBtuCD+HKr2g
FJKI9m5Rmeg1C4pG1LPAQNAxCygMdTZ/Cqfnt/KDCl9j9rxcL4bygy6V2nEIQuh+
YEkLAfWkHjTX5a1GorVtPcOeX9UdGZU06DcKQkiYmIw8rBt/cKhKRyJ8829cfjA9
Jwbp6y+LEHrJ8tHTPE1kbVO7njZCrjbAwHsKwcKG7vWGoe4D3IRZ6HUjIArW3LrM
kzYf7kMkpVkSfpx8OL+barAMD6RUFtlJ+D1GAPHzK9fC4ISKsoV9IXu4cfgNAX5A
vcheIxPtzPwVcCwDaeFs1MZIbDhsrtTzPv1d69n8mXAkBQZsRASRfLDwvV3MYS1h
s5oROq9IgMHkVefMhVRYttJYxjBLMhjWR6EqVnUAT68md3f8rCyPjIbXSXOU8UFp
ppRRfMNJUH5QXUFDO3N0NmfwxZnemYNaPE1kP66IFNpIry+MurrO+GpmfpZremSv
wTlWgqjo8ITwTnNM5MEKm/fZ+VvZ4XrfuTFcmTCnkh1ASK7dPQ7zWtClvKWiS6Ua
C/8+AYSH+0FiqN3/7CSB2jqN0kdl5hlIOL1Ru66gd/hOaRQk9FIVs9p0C/QDPEOM
K/BIpLWGIUI/VUwr4Ikd/g0+HgvE/0yiJggoB8fvYuzz1ldT0fp7qVvqPH2H0dGa
PkI3Cdu7c5lHWNmJinVIHFCEbyV7y1SlSh55xvvJdSvSpjoIVDhjWnnch49BEx3A
yi7KSJ3ZezQPHAwHtG3Sqhr8O0PQyCKhK1kANLNT8G1Nxs5YjxjMR6AHoT2If3te
nA4V5b8M7YefUn1K87TmJlies4pwPf2hy7PF1/tZ1g6WM97U5Zg6gM9aMkNn1PSd
SrdwjisJ570gbogAauosQ/CbGYFQ9nQ/tB1+pYHIO4yWaCJwuIzPRRo0Vgl5SATb
NuPO3B8nqK4ikYClhkNZ1PeHOg+NmJB5yQBytYaP1LR38N2ILYSM58ILx25iYvvu
D1Ob6kGUhs+3dsQ5QsTde2vrGxojLDVZHFwXOI+xkDfOEU4YmHhI2hF7izVfnK1J
m9+9DUBnjx/hp1nTn9/pSj47oJYUzFhSgs1xujgQ0o7SIyf/DA3Ya32dIuXrODxV
g8QkYbeWzbjFzvCgxsYG6llpkqtadmd7cESQPjjMoMGb40eOdtGqXAd5GeN3pgU2
RfhpF8qZiXdOnxRiCh5IZX6UvFT4OrwcKAN/5onQUC+SRqqf6FwJ7cONQYHwrJ0X
U4DoKbQlWt10N1T8ZNxsYPWVWzuz0cc7dku8ZJMYd62uIJG/UZNgr7zg6G0kGCpB
yeS7tjQ8UvCjH446YOcoOgVyTKepM3c0UnIVVOPMY26S7tZHLjwMwBrtcYyaBWUc
x4/sOQyYPh69gaJKZsnUxbWxlmANrv0f4zu8Bp6lZzhb7aKqSX6+Vd6JU+r6/UYl
sELrIXrT2W2PVN6npJLYARELwyE6xucOJ3cKPLyT1hBwTWDP0PrgFiArhgqpMwlh
uQ/HzHMFIS9V55mGqXE5HG3KvhpXgB4noXP6fOhblcNz6jxYPpGuTSllqUm7QRBU
EWZHophEpwhddRwV1MmdAJDxWRIdQ+B2ANSpqpbeWrelQxxDUSkjKRM8eX7uBoni
a3pCP4628NdSm+okqctfB4XFTpjezrEof7UlcSVPrX8XCUqdzN/WP9Nvj9fHIk+m
PCCmYGvmXzMX9PP1gGIYaW1uMlp0ebMFqhwpcRQWMNWhAxSKl6Qv97H/z3Spq7sX
bvuvo4/jlkt9FlhEYHiq4YRKi0iMT8YLsB44x0Zkb1yHftt663yh0lIffrG2l2pH
ueVnLeHFjOAMe4tA7MC4zBnED8Y6x3RKovCZDNYRNHjsJACdusv/yI7dBXAAOL4D
PwxuQp1E2l/Nz32vrR/QkFVaXmcAgPIHCYzXAfi75LBuRnEFoGJk0mimDVTiqGHE
pfzONfdekcM57OFOLvNhHTWBuDnfyXwNnmfjXJjMjQSL6FdVawpeTwgbFHTJ8vKs
2ODUGAMzl9sI5So1TpKgOMq9rgKGJJtYoT8y8ODQ/WphoxcAqcmWTUaqGyv3gSft
lBVBh5RGa0IGMQ3ml1DIAEknMq4AugA9BrbYtiZrheAousXAMDZVoWAHN0NohDpT
INDrP+ZyvI8wQO50WE1r8V1fNGO0KdzsETu/tv8nbzbPZPL1doiH1Jvod5oN0K2B
9FfkeAQBKQSXd/kbkY1XKjxlbKceJ9LL1O9QcAocPRtKgiRnRPY0oV5pQXMm84cb
Mg1EV/m3Eks9ccLk0BVLGDwIACisZhwSKqr6ZGB8nmCZ4zEonqJ/0E6oUgECjkI2
c5B9Q6P9CgZAEG5nQAgSUqWnsH/tCKstC+oMAch8K1deElkqXrExvsofgkbB7cj2
IKlUqX1obcNR4DTScGjBfAhLuTWqKWxeKlr2HtKm7HgPG1w2SEeRKedxHFivK6vU
/GE/A/8H8poYdGTT9q1DDL/ASME1z6zbvyZ2fJSH9lNXtsPr/8whKBXomIonvKuK
0ZsWcYOB0SLdIq58AdlfeHkMQhX+e5LTljbO75CxuJeyrYcdKVqODCWAfyLYGcoQ
+suQ1wGhgQ8iOvEo2c+inROePyp1M0TOzgIPqXhpsDH748zUi3VlVfiHxoZM6u1V
fGBsAAKVHu0r+fsglbyrgltuVRsmIYpsiRMWVcroeEgkls1hSfY2MSeGm5NWyOJ1
J2IR468Cp7/UBBUKVzMhJA==
`protect END_PROTECTED
