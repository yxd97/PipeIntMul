`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hL6444GB0ZAsHw85+EsnvMgCwP7oYZXaScDhkrSSRrvwmSVo2xxmJOswjQFNuNSv
HmlScv2e62V9Ib6DxshVKd+aDHb+dqVJ4wGoWkOmPV5fQXZUrnB3SgVKPk2G87sk
RUzH8o5J1FVzutkuNfLFquX/TgvQnNII4yxpfoUJXctkWVGo2Cz5memiyaDPFBrw
f+ixOYJUTLaCs6myS/YkBx7dSEqsZ8QbaSZt+QAAGmJ6gl+dTCc1jJgPjGavW+50
WQB4wKO1vQ8K29fJlghD5E20vxYePDAQlfGYA/l87AfX8UppEjq0UGXjMpIJrpDp
luDoE0/VoMis9ATVKy6C2Q==
`protect END_PROTECTED
