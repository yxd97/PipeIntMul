`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qj6xQhazRLCkqSlalHgIUzh1e4Ha3gsU8b0fMjFqc+NNCz84Y4m0PfB4rN9TxRd1
ybewOQExkm2imAHoKjAuv8wzztvQ5piMZeb1SDboauYMz6vCWdecgckI35wRLwEj
K8jRRMR/8gKf49xie9nJUNisWROKRwIPjWaXXY0ioA/Pe2OommqlJ/1ptQ/wZQnT
HG7D4hW6/QVbx5ZIa4NW+fRfxUYli60sLoD/3y7o5GRFFqkm3ql7mWzm3iCUG2Qo
VyuxO8zz7w8j/DYsSFPrK9d6qD57suwyQH7fN4605XjV6qc91zem1e1/NLsjbZnH
6ZlkWfXVdOxZxsntxzwCifv7YvD7N/fO0DDTcbeexSVxRFxY6f4pn2uAcxIOK+8E
K/OnMxbxNiGtM8LjVpyqhzV1it5wc95G3eSvftnnHZLmiwiCv5NfGWk398cYSa/W
k/TDZBvZAdxjUglRyaaS6R0KpnNhfaD9maYl2dC9v5hTFIjrWWMd5RDbFwpCrqwX
0kqudsgPoHYe2Y79xI09xYR4W2Yp0vITru76VuDMlC8Aj8LndErkC75FPZwiaJoA
Rasju2sAV4hTQovH8Id05xhDoyK80U0N+N/mPNrq00LHMeiS6uMxteNE2xOk/NHj
OzEqi1SJhmq3i2f/hK+Ads/H4ffFrRsiksTEOxrYmIC55AjAVp05qn33JAXa67V6
fY2KQb1TEDU3oSOigsozi7WTeoBhHXzGoct9q2/oGQptkkCsgQrmPGZEcmfX+0Vj
z8ddyyrFvpNEdZt+1/ecm5QoIa5CFsoSSjOLGnmMDHnWLJzAowZyAqvEuPNvLGff
nqwSmBQB6vVIaUnTQ3pwJKAXYUBamkDKCq8ftgsgENFPu/JxNMjAcJCrqeyozu/v
wLzimDdf2Rv/Y9uzFcXW+qdda9+Y3tLZChsspr8+2D2lonEOC+WuqauIG7cy3LAP
fKeDvGwMTpR16xkEWXWIZtYRGCWKM2TkqwV7a5jHwWA5GF0A5ZfrWp7M+B+FUbEG
qIKaebei/K5sK+hu4yHr6rFe22xgZXE81BHMdYfJaNU0egmPD0Q1nvfjKmdq7sTx
rr0WbsufGHaEP+zmwl3V4ivR9RpdOJ0agvVd9kCyidzCMGy+C3JcJvVNjkOAD+5S
Q6rM1NnpXhKe/xP9/T6OrrCN6aOuPNFU99ZZyOnh/ZtstZNXyapeQznixcE4FSzp
nQYvvQvKUsrAF//NRUiVwsP6STJFmJQH3bKj50RfiHIruDIUXTUvFr9XwLYYskWS
Aj47IetBkwcyf7TJvp8QOlprgpSqwtdhaN1DIYfBC/RxT4Ajq9DbMMrpcq5GnoCg
7Vx+VLLdACl6m64Vx5XPfq6XG2GUh47osrniiO8N1vL+Y/uJ58d4xauQ5pk/ywEq
9cGFkxUsIgrKtAWSazZmfSNQH/Dx7OjA17n/3g1qfV+t+dxaLghb5lP6yADLwWuX
Sph4nmYPyvsKtpTylPMVFGm9D99g/dWZkuixFISjcd5dKGjEDdbtqush8tvzy/Vj
e+hjVFaxz4uRvcXZL84b6kijqLEuEeqo+0HT3MpwDe/vhzG1X7YnHn5VA4QFt8D0
zeNB/aUscIxe61B5MznqvBTgNPepWSucAzdIw2nFFIyR88e97V7KvkpAPaR4Utxk
7TVSGEsOfw4jU96xxCZUeiQyuZF5JUkcu1p2FjFkyBJsqtY9VMATK8gh/KjzTufX
csKsDCTJHco3Ojfdn3EjQxbcaPAp7huLHk/DE/8TCCR9EtgpnjRuFhId5a/bw9yn
bFKujt+/nEhltyZcral3X1m6rDoAbIPWyuhtIGJk11RciTeG/ipfzFObZln2PMDY
FaXgVt0snE6A9R4PpcDpg8VkhMA1Pa7bHpNQ2lVsjTurpGTwY2V2htJ/WSpaiiqY
5B6nLbTm+4hlcCoE6XjODjcy9+mnxnA01qgwpuPJFOQAKOwDqCgPHPr3M7VnjAPs
gZC79gBTNZJd0FBcynqT8bFowlRAU0iJQo0kad411sxZcfEFr+gsPh3ImqguT4Ol
`protect END_PROTECTED
