`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+HUvQtl/cyAExsDfvOloXdIdxLhi0LWQfYJHfoDnfOzhVQnjsmUWq30e4EfDkL5
riVf+wrzU4tBAVmqe/DfGOy/WMB0Dh+KPuekLQcahEzFGmoLo6aQRe5V4M9bSZwD
ljwWMGQOwMwpbRlDwDseeKJoQkYYqoxkXF01LCnA5qW/W47MhzF9rJaDaoKEcv+D
QR7D4bD0S1Mwo9F8gy/27xVhfPFjEEvRl85fL1QN2BonlyhBXUjJaPqKq/3SvrNx
ZCaDlHes9GTOXCPCSib4ZTy3ItOn3vBcLFI0ewj1shPSMc/4jeRz3ncgeGKDgTRw
o31brKss9q3Xrefwdix45I7ak1Hjy0zMjfOhWSIObEJ3rIycRsZNFgtv94qclA0v
PDhpXh/6l2PKASJqOz2SD6B/X1s1W9HhaN6DEd8Ui9Y=
`protect END_PROTECTED
