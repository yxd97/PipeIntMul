`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2tAoAxcL5QssJ4XiRf83F+eRvZ64Rs5mKRgKvSQ6FdDj+kLQVDEMknJtXWBBqGsm
AFv8aimhIZFXLycgiNrjJBVbHdC0xeSUaEq3QcCp9B4GnUrERQNv4Z4/VxZ21jzA
wPn7Phvl/tsPPJCnpa7eRQDwWSsWrmFdi8JFRLCbxxhtSZ0C5drwK/tmShm0AEBY
r0bqnKwaltsbF3U1XTygmElfTntg+FZIh1sQaNJZjccUxgFUrt+JgtliVkilS2qt
Y9sx7D/Q38JRxnDSxhPc69UG/XZNueFU9oxBMWVg45CXXFvJ6xJCnGjwf7nPWT/f
hMqS3J4CamsupBxBTN8B9cUwKq3YuZ7Nb69oKTei1gSxj2bvSz1AXptjXx+gJG2M
f2oRBoIl+K0zLYzijwg2GAr/f7pYbX3cmOphKcbgSrxgeNY0XKzdj5ed1lvK8Rlr
5PVD2CERlEtUHL7XM2oEj0PYUtL5pfcDtLUcqJSj/IvTQ+XZZSKSnXHso7Kfq7K2
RpJ0fHP1iwtKJPQOabA9zQHM38Q3ouzGIz+TuuFZMXeBiAT7FC9YmUAA2zFzcKUu
Bwjy05OuPbtx7YztjemBClplnvXHE/sH43N26newrN9r5RayhcVY141Rd84htLqx
OIyAQEYrnUbHJw85qjGfzg==
`protect END_PROTECTED
