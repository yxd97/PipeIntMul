`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTzUOSwZqeMjCu99j2HbRYETV6F3HTOFoaN/W1zjQw2wM78P4Cwd5fVRBpp8Mj6K
pf4rsGyOAwtzOKOOSELRM8FII4pCkenPsIv+AZ5P2K6L6M6djviA/yz+jnTUkeCY
p5+U2500QcSv/3HBuB2ryV1UCmV1ADZIKbkn0gC31T8YTXVZS+pmPgrcJZJ3eVsq
q+jAIiVis6/5+i1KYSZWf6GxYWsS/nvCVDXqXDyWtyX+Zy1MwCoC0rK7DN/skgP2
lJX6i7JBceum1IL3GR/NFcAEMNz7XUTJxPxVYvpq3MLCouWU3Vx+9MSmQaaH5Z24
XkeE9Io4D9NUB3rxBxN6Og==
`protect END_PROTECTED
