`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2vx8pAhgpynzJsdgoH4WnA1YL1gGvgFlJmC8Af9wXb3G7NrdSW6WBr1lRWv1l5uk
z0a2Iq6KurPljwhrNqlxgSsKHL8WzzGvZWUk9EQuphmUnKk7YUelSakQ3bpCgfsE
ZckxazS7CvcgnyrsJl+yaIqi2yPgjS0ozoEoOOaw1aEfi3blHJqtOArCqlyXPZpa
wqwlgZHoTZtiHJSC/8LMfgDRA43gf716+ce4kSvWU1QJciGw7vDa27GCCtRA4RXh
DxQ34qEDCaGVkRW/ePgTbXPXCsdHJJEzw7XbwCfjaGlea7JppG99Lo+dOKld/aQ3
`protect END_PROTECTED
