`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z48yetVaQCV0zkFw92iZV5xtZukgzWhfe1dLaUT9LLZZbRStfcYHLDvuP9EsUQ/v
etoAAQrRTc5zgQkl6tWoJK+DDsflTkmaYUzJuugPgztt4whMmti01M4sgt5dclSZ
KqDOdebsC128oO6qqb0aoc8yJbXigoWsUL9hcofh5IPPCPSJGpQxpVtqtv27Fucx
QrkJADE9UkZOxObw32f75VKjnYqZaPwZmQC057pniJ3q0N9NLnOkgXBj8mA3VXUe
PyEWEhRx/l1gyEgISHlSSR6Yd1bt4x90c8o4U9mEL7YL/tdEqJ+CH+9fNqo4QPSE
EQG8S1/E1mYukPf0raIOCA==
`protect END_PROTECTED
