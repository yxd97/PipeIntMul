`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkJfEz1sAqfj/nGnoQbeWlYEvFLyqXHTKjTh6ZkYjlekBcrqZItPVAQhFbn1h/FV
Pphuf+KjIqVD2rDJwcrvAL+A+RxVQGGO68OLV6tm4Xb94WO7lqPm/45DCfa6SEvt
d1fqvcHmV4ggSeqCuQIfEmTzU4clqVeNiGjRPB1SqjFKPzLpeGJjovPhYdZwZXNM
6pEPeryaE98Jt9MmKUWE6hqAmC9Mbgj3vyLj41V5eK/SDY9wses7+vnvPpNIxjIS
j4dNQZ8Y2cjaJUkgdpwLVVHM8kJolPhBDE8rsFrE6ogju81R10IeaF5pU+aKiKZ6
`protect END_PROTECTED
