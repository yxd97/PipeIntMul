`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hA1aOGBvm/n4Ms75nq5TFfzCthF+uqYwJlssj0QDnQ76nEGYcwV6rP6oitKjw0im
XHyn5stAvv0prgHwjREtuJ7j52995i8btenkdYceRsd98hohqfHr0gPJRZZHfpUO
8As8Vddw5GiX1c9rJlDl6/eOV6vDJRJgEoXbCAPmjla+je2qZvlWo+JPZWiR9CDZ
ji+F+pLUkVv1gGlnWkDrxc9ZaiMagpV9MBUmw9GxPXywshZ47+rG60dMY0MJE9Dk
JdBiCL+eGK0UMxkPU2u97bxekYIwgXIc4JM9NNBunxXUDkwe4NdTsMSDFom++ckH
`protect END_PROTECTED
