`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHZlBYpFo2Qt+XqjNCZkV01v4NhQdRffrYd6i1qImd0c2yG3BNlX8mhxoKRBmWRF
VEvJ9CcuFccvPUOC9+p50P9WxqD8a/yo3UnZxWwGDf4swSbMKphKRQLCkPDhhyrO
DkgqQP/O4BkGzAJTExCvc+5VLerLUypF+ciAAGAAUL6uiXIR9ILIl4vRniSBTdkw
aNXUphwGEGCFaw3G9zk+TwhI33L0yO6on7NzHDrkdrhlhDpwwpLzYp1qatSBfRwf
SLZ2Zih3v4ax28hsPJIHjw==
`protect END_PROTECTED
