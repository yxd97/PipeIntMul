`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pF+2hVZjYR/F61JGXXwZCN0R1uEkHKu/VmcLcbDOCvebojJcLrnnmVWN0xdbodhk
nijVgyHf2EnYyJwHBVg7AMgIifsV787fFZVQ7FjF01SiHHH/UktdDAh7ThSsG8jy
j5T9jr+BAbpdGm3if56mLFpUUQfTNcIyrt7Q2bKJS+D2BFeTJEMMLhD0p7W4LoTc
44mbgNUCwOutML+qHacOazOFOewYrRazUn104yo/S7YMXwCQE7S8PYbMkmGYji8h
lBS4QTSV5pv7+rW39XgVRVHiOOhCyN8arrWuz7hJdF4CYUR7tHyb/3vN11pJftIh
SeMMSDQmc77AOlup7Qv2SE5C7hqZPARwCpvPa/c7HdXVfvosrYg61P+tHlrMp0rh
UYuntWjKCtZxjtnOwgEtjtOsnv8yAGsy8jKkRjVpJlorqmT5RHxUh6l9GJZxC46T
EGJfAKy7mJIVO1+xtKtt9G+iYldm+5Cs7bWv8ceF8IUUSFH1lztFk0GGYGHwkpji
rXBQvgBU+Bbshpee6vGW6nOmJ1dk/xmPsDeZC9FNhlNtb3cc4EoNypUgdjWU/2M1
9P7Ak/4Bo4mPXVjKd2ti+GEj6teyphAXoaW79mfO8crEynm486r2QB1y4jfQLAAM
ewclG+xhDsjfBwBxibFHLBC2IUJfwfC8MPUga+lAnf8gN4uvVYIyiO6hvbS7A+/T
P+7tN1E2R74R/pQnDegZ0VW3Pp42sg5OJNHZ0DDfH2mFDerbKXV0JPP0tGcy7JCn
c8V2pG2VbMi5/duk+OmOJggBTwYiEAa/0unRXbHebh9+AM8ixqm98dYCpJaMtJUw
kVmRzWY5qC8PwaZWeD9+AVO75F7QVIbwH52heIOJiXZ7ns8iqJMUz41CbpZc1XfD
s6AZamkBVGBKohZgj3G+wJfeKcaMfHrFDcsSB1XplycAnD3G6PRWcqN4cWlqulef
K5qCYvoAHnIx79uG1Y1ZPJgmQo+Gy7ovuShmVrYZC/EdaEVk0/ZkfMSZ6uRxxrJ4
C4fOsz/jE/2eJCnWJho6z2ihCdDyjV5sjKRqPvCvK2Top5MxQxLuZfLi3856xhfO
OBhRNEBQR/0koJXgfwTtVILq11hSTPKIYKOJf23sP3DFLZH4iiU0kb+AvoG3EJil
c+CIzLcAJBCsKFl7KR/dfDZ/r16zmiWL/Y5mXokvuatzMTMBnOtkzrszBJMT7aVj
zfpP2h0GmbSg3w5EDkP9Dxt5RaGS9tMO2rGo5b8xEpXDXbXXoMTTyaOl2clOjWNN
k2rFH86IYIF29Srbg9jYBf3+qOQd/jBOjoHeBNkqc9kouhl/ZSjcOB7dEz9HhbKf
JgWbYd+Nxjvmtju0JCntXtM3emH2JdLjAoGZSngAzZYxIflPafK5YScclQnor1AV
ShB7+TthRX6GPrX/hWAsXvumqhexjaXfXRscojiyxzlqiIdqis82Llx4eMsOlaGL
VyzhFa9+V7RYOZZCwZTtYUe2BMXd2QdB0zELWkWc/k9zptl2XJpL/PHW4v0GGmX4
MCb5IHRRdBXU3CxALs0bo3c74i3QD7Qf4l7oLxmYAQyFqL9wXvb6Txvit71unMYs
QqvWvKFttDt+IW6P9GbwvXmGusl+89AlJ2RKOWg3MoLDH+dsQsgCtvig24Z7YkF8
pk6pPHwaeazHHyCzDQkik2A3b17+PMZAPRRs58qacXVC2M+RapAM7ZTxkRZGb37P
A4oscijrJZ/3Usptm6hGkloyDTvDkzK40fedPHh2B9e+Xmj3ijoXJFnNrkN0Il1g
LTP539u544Z383pxJVjyQRtvwnZYAtMZzFjNtSn+hLgV/m8UQXD+AHy3U/yIgvFY
4CltMmKIqDuuNrn1KpRJtRWYP3g9vBYQGg21jNxDXGNJU52n9wo8lknelL8NQkH4
IqRD2+SaCLaueyiNUE4S+XLBdKP3zgQlG7znxoZiSl6o02yugJ39A95MmmidLd3L
RFfklvHQEckcMuL8Y3HqzW2lgNLhR5au+KUl9rnFLWyT8BeFSU7+daocugBTd2wa
rkprVRmaERTR7ls1ctv9OiDSbsgLAqDRniQnWq8dQhFFdu4CdhR0gwt1ZKzIBHHY
QoSZCkHSSCzBQnznVx5z8GbZS5Z1GazAMM2QedBH+YSrouPQvVU9uzLrcX9pcjFf
85L6CWamVKMsh88MmjVcxcl26apIdG4nhpCNZU50kUsipTjYk0OwWBhz4L0fXo86
MWzn3/Koi85H7LoliH6svNaRSK4CgTb3O/DHvh1BF0pJoCksjAF7On6ATLZc8cpc
VGhCTRQQkKTKCqXDmwqGs0UccmlHBXWQ0ryNHEZoIIVleNk+cGT+2BZrO59kM7vG
KlmIPL5vfTh440oH7TQ7iqrBY2NCgyWgWmGvvYMcVm4pB3XW4CmMeyJJ7OPMlGCM
97TRwu7Vt4g0ptZ8zhQr74w1rFP0QjBChK6nV/KSzX8yspieX71FuF23bZC7a82L
a4AqqQjjjoFwZBN22cl8QQPC0eZDHX8/pkEVsZ6u6wWRpEiPpJaRNF27m71+5LI1
80SZ1A05Up2sdexSUmzFnY7gSYvCgLXEf8t5uOEcRXK2DH5K2ECMv5FAK7M2nIzh
2pdFk/zjR4iuy/ycnLLptyQnEFy/HcifB3EOb8/HKb59H1nVO9cX5SL2kWLBuC08
T+8rmGsPXtAsAqJGSKzjhLtU8J6rxJwRBpauPMignp7p4s0OHEkxBEhH7NX4ckh2
v2H9wAk5rjRPuKbcRxtfWqTeLMS/q/9xLxWnmgOApm2FSjsB7oYKhSRnvqplVUc6
qzojrFAFyizcF8o5gYUkRyTbC9Pz/zECu/GYKPYUCjbXArDH9/Aubg4U/aLbjFqc
tlfz5e+jR+SQu9BtlkyDvG94rv6Zo7zDRnUM28T1a/w5U+8VsSfaiDQ6GY9lJ2kQ
uUcQwOS8v6hKDyMyrGJOs7a8JIWbNT6nc+tfL5N72U82P2Ted+7X3bBoFlm1LIHT
CLgrYkIPuNWmnY09L6oEPxTzCkEW0cTnihuQiC/q+vWNa+gOtMwEDVlGWTaxdhpN
uQYQoU5MfshuVdT/oIOYmKy95E4hIGDa0yWjPz4fdRdJmpo1U+9ck9qaca11eydV
V7ZMilPlUKy8tgDwLM9/6E0O1y9j5MaOaXHypNBnSjlGBl1eLZFXncrOo0irgD/G
TNe4i6o4mHgloQ8aFt6toEBUeJifCJhL4z3GeSburcgKJfFlsHyb3CfC4Z9f2Med
hbYjGcgZmzS1Fcwe5OkyoEGNoYtrgnOJBSZA4m3cXU0kIcOg89qXkI1/IgFDZKhV
sXS46O0SSB2Taw9kw8iWz/k2sBAbz7Z0uWZ7sDaE0rTDbcOWSIA0ChCUYfjgtt3R
yBFL0SFsJIodrDKGuXap67VHHEZ2JSjBVXMr/XK6SXG2czdku1PbiwRJ671V5YOX
wDI0i816mOX6VGaruSIuCZFImz2oZLQUqeLReWA6z0flIHlX++3yvtiuiBxLJx9O
z0c3lIc37kp/I41nOAd6X+eH84nsAlk12kkfPsfkdyeEuXBzVqURmDLwhLCDvFZW
v/2UmJrtL7La7YwouP2GefuMu7U8z+KWpgfMhVae2eK+84Ak1V7WxAjx89HxCARh
HZ+rNzRRafwHtRnA6kqP3hIBIWZxj05G+GVMx3YTsLT47kZLEp6lILwtbfSvQsRX
LNAOT0KoLh5wMaurWVJlUmFJMnyiFzWswIxtJ6yF4YC03MZPwdgjTA4rtywSSGZm
HU2duSiU9P2wCP9UpjyOYXKHjuOLSIu/FNLuqQX/ea8i3nOgXmxBMYpkyeAcQqU8
zDpPUp2FBFpIkXOFKyzaBict73iDqifjQO5AwuZNO+DvmasSULRHcSbsNjfH4Zne
j73flzoB6hFCK2eI5RnRlmucdZyjXKaqgHBIdU28TOD+Sp6OFDXjvwDgyy0zlttG
klTzeNdvknXYSkBFsoHFPyHOtr5f540fglZuRJCGO8rklvzFcGEwRXpJaGJ4eKQQ
OoxO0QjpluAsyBFu3/l5gY4xckhjdhKptNXtTDprFCoxtTllq1nPFHAapN8Xutvr
sD1eINxKYf5TY/9Nv+I0DN+0vMvPIQIIEchnhQ4ysGBRT9KvgIYhfzwGn6PASmT8
oQa4T7nezlrccWOzNtHuIkuynNpLY+TKUdvMavoerHFSFCcrtoV3Oyq699IcUxSL
seZel1bUQBUoHDjXl7w7TBRbvZb+xiZ51hAJXUI3fLUNhlXzy0DC8ocxNCtrsI/0
MAM1cmop9tScrU0PGYkgX1k40JzHCY+nqVI99k9dsmkgoryLr2bvfqhV3XcZe6UK
MyTPfD3VTHx5jL2/SbL4P/hoOpNZWtVvE9NugL87xE5irENszIb3TngRAOwPwL8Q
j8IGF7XwwCoOSO/EI4SWfaXgHbOp/9jzTUC8AKJhtqPti+PnAcvrlTPXRZZKHD6q
RJVgUvFaD3xHfMMuDR3EqBKfzbkKT04n240wbxOCwB3ehQn8WEBeSIPaRsloKj1L
zyo7xDEaR5UH997ntvVJk9FlDbrOXvZEQr0dii9y2snd/CxaavPBSq1IW3JanorM
+a6FOBJ/DnWxargRYg7Yiq1LNEHrPFhSGN3AbdrGaIiXiAkrcPJbwqrkO/OcVnD0
3biKEWI7eBKxb3b5odWBWl8pg99HxsF2pFx3y8RePl2uTeW9CVormZjWvJ4l6bij
P+k4U+MHR0Q5DWWW41hxXMJjNn1MZnUN0iF+inC1TS6PC8Rgep17u74xYsJ/NmSr
gSfUUzG5fsD1YBbc61AY6NgBVyAtGEVi+0JO748aOuiXjS8uWjoF1KKTwA/8qqw6
eflvrB6Bck+NCz0lVADVogoffRu42dKkW0ZLKpW1nVKhqZKXcbMWoceIG0j3++3/
JWbDk2YL7d20EnisgIFLdYxJjf9CQVLMV+tA4He/EVO2Gppyah2DzygC+UpPw6Xp
JgKLcKRJFc9EvUQw2VTSiMUk+YUrE3LXorOYdc2lQjnClBIRYQmVP/6YYCTVZK+e
drEf9DhEsZvgyKHoM6+tjesy9KyiHZ1p7VxK5jumM6o2yJ5QyQuOEdH5v+zDc/pa
HUhHBAQjSDScazOq/0ZrYo74qQv57jyPr4iBlk+wEHdqoyKTy/asv+CMlxsmT36F
5jXK2OJoC9xbuGUWrs7GOZ+dSl2GOq7bLdvN8/rmyueCnsMGhDXoeqMENpj4zC3h
pHQVLOhgWLd4na3iQinRSA1RsndPxVRCAqrNtOH4IyXj8lLT0F/DJCI+KcmMQIKz
UQH59fCibMRTd+hnV5Gy6waULTft5HLJA5cdwJclhxogQOLUyd0K05PeNim+WJXV
31tlkty/OPHBZ+ztB0wesKzqbzXRNfUUGVofqkQRhQDWMulkm3b66O4PyAPjRtJK
ZvYH2WZWHSXGNzBZUfqQxkQ11j6Tj/+2VKmnFoyMJEhWJRBfG/wT0kbISXptYiJa
LB53/L80idYytfH5HIw090G+xeWhTkkmr8UmzS8FtVpvuCVH+ktg7HA8+FntuOXP
evLjJPZamjMKxA27v7TSf/Dmpv9sXraYDR0EHWjtIHSQk5sOANFkLXBmQ7Gg6Fbg
TsSJHNNJK5KHDe6qyuv5a/5HS1WSJp1RU6HFKM9N1Z0nvmmcxIEo5G7HDsipOpoy
hjjZHuIt23Je45Tv5+/0mCqbnqyHmnUBO0+HLshmmHZYA8Y76aGwZrxfhRXwh2AY
`protect END_PROTECTED
