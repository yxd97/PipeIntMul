`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7KpkoF5DKW34YabtpZkTi1DLvS9u1qn4brM+9RvnsWWuU8lBvnbI+CC7CR8YvaT
fDcRNm6p4JjWfjGAga4xEMJA+CrA8mo0ir0IS4MMdNipVOzaMIdVj/aYoomRtuYK
zt8ovr4esi5mdQTp2Xi63b5WoiOdyxRnHeSQ332rUsd/L1vNeoyD9WMEB4VYVzfj
h/F2NWPXeUv/bmJjN+7CtAxfcGMGlncJz2QMNT2fr4VsV/URgdNTnMlF5xm3BZzz
PzftrGsUBf60L2Y38IP92g==
`protect END_PROTECTED
