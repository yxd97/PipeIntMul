`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1v9lmpcxx2MYTs7hXK+R7o4I0XVjKLBoOd8D7cTLrJ9w/4na4IuxWqnZol81/jq/
KbbPb6fsBhSrCIpbrgv/u6sfLqjjHI+/sI6wNFxPqCeaK4eLY/+iUVkKdcLv37c+
HcMiHlEJEamKA1fe6pBpb9ZVfK7ZNsegKCyxrdrkaqlelMiaMjnTja+d2h5yz3Sx
UsheJptwtwbjLmMaJHfLYYLkX/hoVITwMnyxq7L0LI2z+7PpjbbaNH9pPCNnm58t
3Qmi4aK9IIL9qtKbtN+6fmBmF1Gq/f7jGGaBptvSKUgi0ttNSTXKTuXBPcYBgMQ6
Fblvc/9A2lzsFt1pf1tjEodm/kSBrn9gmLWR7GkB5VtXVgQtYoPPKLkhYr/q9gyE
iBRgba/sC2kIae/peC0Giw==
`protect END_PROTECTED
