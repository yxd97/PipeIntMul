`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mji6KkJpinZrft8c7SSQDg4StdPxDYcfuwckVNlplvVdozZiItUKqgMDLepSVeWC
t9GtRP2gdV31e8vLA5fXX2dTR1AkpKqzr9AVj5F3E20gC/iE2S1Edo5aW07AGD9b
6OBxK+8i1Mx5uPOYTKRNDGiQyk8XjGrpHRkLQWT+uc9jZj3GHi/VBeEXtx9MtXln
kD1T3MBtqDAUHp/W3z89mc6Jo83T+U5MCOB4H2OELeFJsRxuq2YorzmhoWCm06zq
xBlexHwkDEW7oYFILMpAacLK1qSvUYg0bF+iYlUH/h4=
`protect END_PROTECTED
