`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxiE9/VjqeOTS0tinj5rauuSbWODKMbbifqN88u7PrACEeJwBOwk2DwUoLfm5Ati
2rVC2+1SoYSCVp4zcWmdl1+QdL8hEZbK2dGh9Ym4Ck+vpYwQf04EM3hGOBqF/xoE
CmQzwJHZSFtZVjAg6Hc5p4MwKQEUuq+s7+hi37GfDFccvpV2koYl8FvY6FxFCRQt
Hoq4/L1uWGlzqzwIgFKEP/zAGMTdZ+cp24Aja9e7gKvjxc9TPXDLwOFA6f3VPG7y
N6RNYBvoBrNTDeRisz/WNN1RJe4uEnVzgYHpHsnwXLrWsPL4qcHPx9nBrluMmnTD
iWe25uLO8eqgUt1vUhCU0XChL2dVQS9Iw6PvV/++9fEU+L8AL7Yk/cxQKQt8QtLC
WclshD/tYi7TbOvvtkUqcBJFeriIBiakkuorwVSzfEFWdGr7XAxVCidYCP0ebDzM
96oIqU81UHtp44F3BjhOe91jyldPJnh4B5yrpoVzEGRT2au7F1lhUSe3YTQWclCW
GHxnlSlS+8PH5D7Bn6dPKc498z2tz8Md18P71vljjgjhuMx9V8NyBBvC+5P9Ecdd
pTY5FbPLo+CWLhk+PqS0sSFKB6/78b4/UW0Qxix9CrKlecDpozEo7aXrjp4SlGX2
91JqLTn2ZpRH/PLNCVdQxaNnZN2SCiuzr8irl8W92t8vl7o3/QFv59HXKrTojKyU
XX+hrmZxBLQgPmtCWBJGkahtthNwsCm4DNKfhKm003EFvBp8i+xLZbWjvqRMgslk
3hzKJrn1HSQV9S7Ir1OWLXY/DNc6yWaN9gEI+UXSwINHlpjrFz+8x8UTsT7BdSiE
LgHBicO/rR47+yNeFUs6LQh8tjVu51+cv5EFequif5CgoUpuLqN3lyV0Uh0vL3DU
YEbDpImv94/LyEzsc9WZxjpgWdLZSuGQzS4mU521GBraoLMzKTX8oPiqssd8MVzu
oYI1sH37zVLTdLZ4FSR2DpQP1xLpLJO/jIyLRIsKI1Nhja1VmXXC8VBXxEFlcLGo
bybphn3/1OyIKCz1x5UcqgA2ypTL/JyCgpc5szfVmZUFewlPwcCMjjU7u2N4pAjr
jB13I/OBXSRyPkgUtBKSGLgpcTS3aZcJcQI0eZvI3HrKMurcKCUvhPE2B6NvWjcs
m6VepyYlS8DZqOtUmCeSk9MpFUQHyMYg+x8R6lW3nwlz53PV73pv5+4Egt46a2I+
`protect END_PROTECTED
