`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tnjt/dnYjaeQlqVQZ/JBvg/vGziQq5Z4tA0iEuTMkUYPyDLisc8wBko3OZymXvIj
bkMMjsEuZhjzkVK436BLBT7DDa0iRATkwQHro+PL23fNnpfI5B5t9OW4NXM1zjmW
8PbZ/WeYJJn0IJgDpvtXycKy8ycEiRmJBzP/34glf2XDaOerPYHihGCBawQ0M3wv
UqBXrRH5sLQ9j2Hn0/CpTrEEcFAO96bLyRSgLxNGl41npFEXEZCRQQ205NJQ1AlP
x56rACTIBvgiGEazGmXqdnhBBuz/6qaOxVo3m7n49aAKcEBc2o0tbawVQ4BhLTQG
Vjt93it9Tir13zHmzp0vvg==
`protect END_PROTECTED
