`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MDcYxkhlgdO0h3/jdsDw1CHR+/UraGfADQAAXFKvgAO0igSn1ayCHmc9zUDHMk4S
cX9n9glMrzc7KMuaR/YxCYip+iFdC/8Uf79IParZ8Ipha0k6Y023qI/j4jWOGvi4
2Wt/8iIXdiEzaADFwoOE/mETvs5+dSq1FLEPTnmZ3IPeZQDh0HuO3WEl0w7lZ0ZZ
HXSFTgrQ/NcENUE0lp8dxHcLFwuSMeVGpaa1yks8dJtiUaZJ3459KrSwoscNg8y8
0vOME9GNiQ5bpWFjgWnEkQ==
`protect END_PROTECTED
