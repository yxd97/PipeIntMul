`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9w+fnYNJi7XJGXVab+BKQFy0fUCjJOXlMXl/iJJm4lfqcN4ukx+1axBTGJyg59c
W3AUr+O23Cwi6W4PcjW24hWuhymYLrcR+Idaz5UDtEH8mQ18OYx3WXqC4azyLQSI
vKg90gWrdotJC7tCVhjqWbDI7z3OZ4UKX6ikjumuhundcsJH3/q1SO8XvlwdgpS8
ueyW8ytcWyKEtRyZSeZc1USXonYMVayvg4zYEg5kxY0zHGUdhLIY3lyEDvtnkvmj
yeurNZlxMHVfDgJI3Pgl5wsv8AgMt2pgDgk9BPOifxP5j0i11O0Rz5z1kqwWyidZ
2LYs3UT5p4crZuOSjpKlpnGWMzguWCPd/JKXHd+vCOmOpkD+6ooELnTdaRA0hpWT
bDfCrtkSDbVy+6V6ZXSU+aGQlJBdlQCpc9PXcrXEyIGn7rpir/n1YBwf0KdxR8RA
T+3Bj1Lcxp4D4PkTK1o3RQfi575WgrQU+jqpRWTKB8T+A0SVadaj12I2EaPjNl3A
4eBV3jL7BbClTQlyVdUqwb6nEZxXJALWjCiayWs1CS1UMCsiuU0Cp8xpJ8SjmRRR
7PHir6aoBKgFd/+ykHivJA==
`protect END_PROTECTED
