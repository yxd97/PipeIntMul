`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29tQiL6XgFPdRocv4VGkZR99mDo+T1I3soZebVEc0/wpWaKC2tW+f6N0b4WRYAP6
W46GP9qPGk1UB/9gnX1toVbSKHno8TDsrDt7vokwYIEKtdMyC7R0aqJYq5O8LD+Z
azhGEotjYYnaIF9kchftBne3wh5LP04z36bl+ydBx9lzdVCSjHn4P7lohBxLW9Ru
hPe4ZwBcVPkf0VgoifP1+WImvYubFtRm7uBkC1ncItWTrchYFCIddVs6a677r84C
Lp47mzuPxqrg6+OdWhWsak/0K/KBOuNMaReis3S8/Br3+j2E8M6KMxnFXG/KCfuJ
jIVMdbD9mQERySng4ejfIfMDGiFzPgD0MzXesBRaskdaRc1q82yBTzmmv7BJL0uJ
CJG+qRacer7UIUO93l+bXyOdVJmzliDPkIB+isRhDKTdQrWL9iMErw59CUJ7axGG
0BkX+HSSCrgqdFrvu2HQ7XWEwV3TwLIA3Zt3W6Ev0R2nbo2oi0WOwcI/nuOKP2xL
4YNK62CANm7xT8MQXyO0ticXfGmA5Sxin3MwV00oKfgSA5iSZxjIf7cbT9hu4Ioq
iLwWmRToVotpI6Jhq25e0kPCEyYylHtPrbc1CVE7nrweL4ia713ILM1IWPLBD9CL
JkQ/Jl6MJfDuOvUrcdYGzknpxPJlp4TSBy91g9/FPaFkyfMr/QFiI84kwdWwlFZX
`protect END_PROTECTED
