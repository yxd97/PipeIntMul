`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gi0VkYkJgd8cwEBqrki1qmPsZ8dOQpt9odmglX1jnUoutM8uZxoVyJ4cupaihaDP
YfbrYwmP0gIgh2ulOek2dwVKDyarPo8b7Hvz2pQBi+HA4V3RfQ0OMXgpqs+IZdPn
BFV07atNqpyuGeR5MN0rKP2gUar/ToM+YSVTQ/yzZlryBVE/q8DrVND4q6aS/wd/
6AFF04RHdrlYTWHCbUSmUfd8D4Y5uaMwSCg1Rc8bwumTMg4364HXwdyg1fhItoN/
YhkiQ7VlzcmppTMs9JGpl08MQnq+ZUHGf6uZZhN4f7T05eyc8H8e7rXav8WwNdK6
+3tW+9J0PkfrJOXY2LP5k6adHfmmwxzsqsl7oFrzLhvBTRPhGuE4093mO4WgZgWB
zZkujCbc/axs+p7am9+ocRb93VtoesESHjq8pCnYe+OZBKt3qsXJCXoEVjvRgvvm
bDHcXUNL/OTIni13jtLF7A==
`protect END_PROTECTED
