`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2czySQhG9grYMDKZotYuDhgPkB6/cLcIWy4WPdEtuCyE7LMvH23a3gn8QUKCHd2P
Gygn435XmILl2gpVLIrEBSFtpGNEaWtfrgONRsJT5VFNJ0oL/uQHDDwkmvG6AEqg
QXBe9SvSZ72B+tWtXwSErVm8NW+LWpKpBRJ2WQRiAa1Eew/AJwvz4DPBlgR1Rpki
fwMbTxBy8rm0iX7GErfeWtGYXNyZ4pNT7wrJRzJtw4ZbqOYKeMRWVevwGKLyUWWl
rPBPRpAOe5mGBkz2usIfDZcZgAYHFhNYCt34TLiok3LVgYeuQ9me8ek9rgQ6qPM9
`protect END_PROTECTED
