`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5JJBgg690KwCkSa5vfrbt+IdnySskyTutdX276bNd2uhEoWO7FNkYiztkNyrRMY
q3B5VInSGdNQBzieEopVu0vaWDsWkf5Bmuh8up9YvIUpv+wMjDeqmkqSo/t/Fp/S
UbcqRKwqu28IKxbLaiWTeyxKHc0/Ujryd8uqSDVBL4TYsOyn7PgsFh0QYPyOZBri
aX/pBQQiLVGv+JrshTR/ce00qHxd6eHXZIpdCnlfCcUKPeBUdToJ3VRg20ciP44M
8gHifL52PfKPDdAtLhXcG28d21N8K8lJCRKHoFRnR75CgEgZngs4jMljEHxbc2Nj
bUb8KsGC9+fqGbs5eRWyd5fcZQzyie6yy3eiTPAok0r166vtixvD7Dl2J330/67u
VTsdP48/Q8LsZT/TrR/3IA==
`protect END_PROTECTED
