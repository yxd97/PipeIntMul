`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TWou6PqSAPdE2XiBizw3RC61dtxDAOiQicGB6Pbvh64AxYbZYBkORXs+AvdEGEsz
a03aYiPau+UJgPEv4RkynNefMgoqVr2S+6NjYdw8YzNNNARlykaTOZrvTfLSrrY5
1NHNPreo1MmkmcW0Qu6Q8U2T+3qQKsHPxS1i93jg/OlPR5lBlIyprldzl1MKJgkO
Tw6juztdFiy2b5vr24ZDBvNXHTaRN5UweiZTdZ+7+tHO2xpL6iDzqY3XfhKQU74V
+KdMiUi+i5Gr6Jqop0Snng==
`protect END_PROTECTED
