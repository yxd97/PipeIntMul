`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4C8VFFtK2zTw/5fjbc+G3jhKlGOWKbB2LQmLP+Cz31wW/tdshKvsREiE1f6aY39
Sgk1fBCRXEWEqF5E8YOBI1D5Bpb9iAX1leEMHOkDZei06WpJQZevsQAH7O+R4F9c
QM5g2zz5jE5nEg5LAdBRytEo0CB3jMmkX994gC6uOOHT8ebW+hbyJUIfAm39GLqn
PnFmGUy0e3k7HhsyIJI3CxV6HULVDSYERk81GS5kFpigkGawqisFbYFSqXhx/87T
/PoR6EEhF66JJ0HcIFRXBTgUav21ColWDhoZNTfX4BIRz8R/SmMDttwI+ONmZLWW
gUsMplccaFe8SV9lI/pV1Ppl643QCXtwuGNGrJXCrut6PLA3z5Phc/ffZio0WLsy
CwO5r7FR1p+HAUvgnHDfvc+viO6eUPLxyI8fMMH4sxRp0mCpJ+Bj0BA0iWgG7/qB
dFdHSfsUuFEqq28zeStyuSm7pk5vgn9nouo6gF+eQGwoCCBH1lGyVcTjn7+qFl9a
6Z4okFtKQ4IbTWlFdgMm/g==
`protect END_PROTECTED
