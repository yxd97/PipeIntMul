`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CqxhrnVybVmBi16ZN/L6anMF4KUZXMZE7+4OuzjGjnQCX/nD5t6I+h/AXMYORDNt
uRBVnDHAGY+gOs+Upge07NedJ0RBMOuM/HQ6t3q8qDI/WQ8vgkCqN1ErpqEMGhjS
J/iHxmYeoWVUk885aQlf8WB7fTX+EGoIhAtnO2b0PWl8mL5mCt7rOf6XrdCngueY
ZWORMHRs9EfAAcrbMSyviy3gC4MrNXrUw9Rn3V9N/r2G7BetYI16wkZS4NCt+g35
EEIPQ3t85J6IkTv5c0tvLGEdHF5AvukQmhzy4zENFOqg019Z4N3eGkyijkSsEXvG
YCDNj0cRsaQrdEY+2CBFlhzqrWDOOS8/3TVmT66is93nMMAdVGwji5XYZ/qmg0KG
RUUoHsgO6E07LzWmKPgGjkps8or8/tbuzxlRUpmTKIy+CO4tKUhuPbfLW7tR6iwV
mjR96Jq0prrPZ0vfPKNqYsmnJZq/AJOkfVkzAY/EXZl76wcown4XqUXYdnWQgA9t
AsYBsZdLj5doqBK46NBztEI79Eg5qQJHjVXaiZ9buk7OHXG55ecUiYrVX8ZM7Uia
vXJJz0URIzEeyCYH0CfrvzHlONu9lnM32GvJvret2JPOdklXe0N1X9u6VN8SylS+
GbzlHvJwNwNVIXBB5XUvRX+oKgIsmaPbgXUjYX0v3Wl0BNYp4InLbTtCzoE1JSlA
g2X0DxOzm5qvhtjZnzTeUIC0sRwGw2HGTejW9jkfLHevM4XDL4Rq6IZ2M1meTZus
F3sCRYermFcA4MJ16vzIChBIScZxMeFLDZxVOnFmqBDAPmTmnhWSlb8JWo0GnM8H
UzF+NzPzaeZ7yhLuWnJbF/MSr9XxJZD28O8F2UKzRhL0CK/jOvsujCWYn6a71RZF
qFcZjh0C07hGM5uVHZkQ0afWb2Bz2AVw47wwkolIasqBOzb3l2bOWaSZcvogwlu5
t0fd1fjmlR+YpEaJhO4f9Yv80RujHKshIJrJBHbYydHfSGoiWkAB+7Ud7vlT+0go
z1aUWVeIlT9tGJjP75bQsGJ0+NMAMQGf3PZzQZtLSovB8/sSC5hWAwtTuyo7ifOp
1d575L9yUyO2+rM2jFccl1luoW14K+Ua8kn0zfnSyH8WAZrNbZ/TN4Xc7J4Fna9K
3jnI8UG4RtzXmEbrvtm3K1+rOgiFL9Af6mSnzBfdLcEZZ8QdBiuDcuNgRxcFOFWx
20G81x2vqfwjM92wrOVt9bwhDPY7lvza1CUoMITWkocBGQb4nx2pEBlEqvF3/eeX
+KvrNVSORf/7ODdm9B6WZIG/a9PrDXwf+xMqoc+bZle1rpLPeIpkuHeTmG9krqtU
W+vMHizXLAHEk+eEdmWkkM+FbgBXOtdpLcQdfB7HGR1usG/pTOEzqwJSkUp6ZgAJ
mpiaO1sc4GcUCeRCP/CKfAwPfdVbuqa2O8wRE5VgjMpnNKKQw/1ooCH04TYO5uh6
EDdNL5iDMKH0+ZnNLFhhu0YDoyZHYUsdKat2JEUTqjcbaMp7Hnt1yaS7w8wQsRAG
+UYsRQavT9LwxXmUSug4oq4WFXzvB2wkSk6iDFrLyp9+lWj0QsuYHZ0pNhr7uxYy
VjlM1I1/zut/LVa9BPmZ+XiOAhMnFQR6hyhKT77NN8cNiPMvbv1gll7RHysUb0TF
ZUd1CiSyKlfpuRDTkpKkbszHHng5Ygy0NUJIFjaoqx5JUdXN7d9b3o7YvaWN/kzI
m6GQW0WRdX2q6tgYPqwWS5i0N5vecCUXWL/GpKNkpD2sQnNWNC9vl2bGurWeE+Nl
5dmJl1NPqdEZ/qAfCF0hioh5EnKpdOE7xy1J39HA0xH6NTU3E4mDGH+gyZkow2/7
kqRPLSgr0II0mF28NzUWTRRaktZUmzXVh9QdxdsIaYmUiaYHutnnM6yV/06+vG3o
EoOt99fmzGA72RCe/b0sJyEyD7xSd/bwfGSl9MTBFSv9lNHpyuC65Y8UhJ55subi
9JcxnmWFW8HQk++DT2JBCF1Q+OPJ0cSv01tVrI5f4ULh0GlSc4tL0ZtY89JLTkA1
QxDK7RPHRw7AkjDkH8GGF0EtyZm0MuWq9R0BjxuV7E+vriefmsYhH5krxDm4rGs/
xDxzUbuRqBDEdcEeVI7VForgADDJVtOwsAZOIghPs25hqrLUFTBEu6l8n8GIuTVi
SVSsyTNL8Tg5WH7FIvmWQ+r+/JcBztOIUG+aPY72gZo7b9bBigpi9uCYN9/YI6Tc
k5VmTzzZQ7vtyLBlgWfQdi8OSvBjIIxW8vIWJvbSj9/t8dJ0duSSQnlTtR/ShfWf
ODln3wmIndBz7sW+puv4Kb40Wd0zTAI2VlF2Mm3K/TGhjh/HxSG5IFY+BPC4dlBQ
EXTz6BrzA1jgI0XOpTiqxLr+tY7xHFKV2VjPZKD8gaoidqcAe8kc3JFajfOU+8Cw
lYwZzkEP8Ghb4g0FXyN8TBy6RueB8z0Cov7GEnMUgI4plm5O9G1yyugxzkqt2TW5
LBe9uV4phw7BQ30OfLtL6XUu16hyOEm0opO1++JUonoUClmKuNStYDXDOBZQJMQj
yR1Wb63DMMHgU9xsLzxMikXVZ7B+0/SPNgguY8xVwDGvQJniOGkaxLWBV7wzAp50
+gm90DCJxm21yV861nwqZK2HMRgZsSq1JmOqK5qs/vVY5qy6zattCCnCDye17lD6
qBMMPGBW+UxCI22YVoQmuwDJP6/rpH7dVE/AsaE4PmIsx9bctWkVWPoAgmzxpHCy
IpM5peECjzbBIzE3J4035KloevoyDD14jYESysp765l7RdvPYNlNXXppvK+CJfwo
SzqfeAnMeZYS6OL7NZOJBU4DTLjAeL1aWqY4WxW9pobdihtymwFYsl5FTVz4h4M6
RmY5g0TWinlXGed66X1mc+8CdglDeZc+KST0tKGuiIkz8bgATppzhu/W4ZZ/orPU
kQHvGqWnO+nE/KdhP0iBjoQ3dCm6QE/G6Evr4ewwWWNrjxXE0MyJTF+0jLqC5V2V
ZRz/+yfkq3oKDzxYTnZqEDj/pllNVGvZwo1apltK+gwgcy7a660TnTI4WTCQtPrd
4/5KAWFJRO5E3ug+7ZMVVNuovvbrcQ07RZrSrJP6zhmqaJ6O2aJTU36FJX1fvBHG
wTnIS6yQXYLzL5UjRzrLRNrGjEfxW5gjlsy/bICH51XUzFT49Oe8XFl/OwRV/bk7
z/LhUB+c3lmoelCJ5xlOoAPPIFG38zfsLzvMfK065OFu6E8VgYwr/QCgYaAQfqs2
I/DUW3Z4M/GR3D6532ODTAhN1DoPSpule/j2LtqN60ZFn94hK+mMD3fXBvNv6czf
kRKMZPMIPL9sgxZbC5O9JetCBvZHkDd4Yz38y53hjmQY4sQjiQhiYKleoesd4KsW
FOVXCqQykKD4e8VynMT20KGpFJEc62TE4wX9IEkP8dawCkkINoR6F6/OrurU2J7Z
M+buEZ+uvhuQq30QKwHJS2Ug1bYg8Jg2zIY3rP+GRZv3UfDRLEZ9UdCpdyb+DYZs
MePv+pNQ6a0ZQK6eXmCeMlbU078bckCO0zjne2KHb47DJ/0zWeJ+UoFSfAT1NleQ
psdNEvVMGQjnHiAIoXbhLqoHcUSY30qd0b52/qMRHvYe2fLwdwoTrZgP9QfmCW4J
WVZ9hkcDuPaJXH9WFzeMQmxV5Dej9zYgaPQN4N/mu/gEGm9Qvbah+sGWLPoKjyaR
v94iptmQd6F5UDoT3JU9rTthxc3kroEUl5sJzPb/MJkmPKCUSdRF6SNbEAkwMSvc
To/dmc1H1p/5N11vhRMdDpzKLCfNkjVMD0x6i/2BnsKmpahw4cQIdHzOUgPe4Rr9
Pps8iVw7kBVcxt3o5U7wTWcdVg4Tiei/KQAeDhq8m230s9ErA4O4G7sk9v6pb9gX
KNEFxm7k1PS2N3E2S7J6CLLtpAAAOUnIJcfdSd7gSgig3thqxqdYsKLl3I7Q0BpI
ZWIlZ3i4CnitFtKVmpaCwzzjHEe/glFSSewF3Pm0hNQ0F4/jwmO6Ydin86T1Fw7I
jgJGuw34hfvHaI41E9LT5Lp3qXkKd/osGgcoSaMdGQwRYQVilHZr+nF6JY0J4DRU
p83TlaLMf1FvS366jOR2fRoFYJTC1h8U/rPxY5QeXQ//f+AjQM9K94r1QXjRbLzG
JNIIAt94znoXOfkGKaKQgSxx8dHxbZ0JodJVYT+utmgyfa3ODpVZThXG/Eodh8F+
kg4TlBu/rDs2I15Xjsp8J1G555UDbgGh8+vGL+9DH8ON5jmSRMwxQw/nRpR6Y5Ru
HGvGqxxOFav3sXCdRL2Z44+LjtSCYX+jiqUOxhinuc0A5STEoNtwNc4XF7peeA1n
kDrayP9FWTCybaR/m8U/yF7qcFv/Y9E5be2gjkQPqIFgQBfdtYITo3oa2QWVxvPI
vD7wopGyexi8AW1K/DMLRA==
`protect END_PROTECTED
