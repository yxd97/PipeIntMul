`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
grxFiBh85k3W2oOgRAcBK/8vUSAaCgex2cgfC31SjXLM89TJapwK0hlBP5VLsJVl
wkTaBq7u3xyEJW0YXAh+uAqY/WJ43vbLfuc7wA/5AelQY1KcNIlA50bK9qt1Go42
WRgjZTYexldEZjoFTsG/4pLkKYmo368uElpbMia9Gl5ipyvmPCawEAzGcH+fWa/I
S6f56zVheQHBUsib6IMCdseG9fp2lpkro0Rikf8ti1FpcSKq4dB32BU0uQINc3q7
JX1pWhbhi1DPAlXmm4kMdcUQE9wgkd3nnbcXRvc3A5hMOeO3pCnzcElfYQtXOmPv
ESmw3U74P09o9V9LayWgXVfQHXCLWBqfpp+DkNGK6152BOXXgRpNhvFjCaBBmBYL
oyopzrUtzkciQw2ju6WR9N9m+kkV9QDMeXyiG+uuUzV36wzxuC0IH2ZVpP2iR0F0
BU+hqup0j9J1LlQUDVcQj3FUT+w5LUknJCed56URZjUpA+ziUceyybHM67+r8sV2
RQ5OqYpOu/Ghtoo5H16Ksae4ENbSOtRF9Qet14rihKBdBDAlJBkq/kcnWKS5SVyC
cvQLPl9sdJWbafO8Wp/dH+l3rrWZfzP9tKQmpkuTwB4AbE5KF6pIwfAxftBw1hMc
6ZrQOEWk9vlzaWaTuAgSPMFyC03iLmNRAVNMHI+48YKwQJcLiSXE7kgV8ziOhxil
GTbC5v6SBz0QrTG0xIKGv4bO4MXDHIr040iLL4ILbCx5aBSKOaQEIxTnUFL9u4EK
OtuDzTD8/5WZAUqhxci4YDb+c2nBgdqOoubUsIBQzvg=
`protect END_PROTECTED
