`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mBCqmGaUmq1vIo3j/pX+JICsBiV7fg3xjmPd6Vfh0w6iCrkbX7rT1z8YTwL54nXZ
+5Y84yLUcFQ86op1J2D5BjIDxdDrYHMboauX1UNaoGtyEbkEXbEIJogX6RrSxddt
bVVRA+k2oy/ZTKH59TRZ9QyJB96Kezv40IzOwhmJ1jqI+aOtsuECCabhkaT61iFv
TrZBuzZDqgaorXM2pSBsThBhnXv0mQ/u+Ig7IAc7Oqv9ZATgT2PAfnrrDWrlCt87
p2XCkQhxqlK7puXIBmX5UQ==
`protect END_PROTECTED
