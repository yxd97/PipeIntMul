`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epk6d5cA7H8YPnzUdg3YI7HYyG2P03WAaS6ZrAZxFZ4hfb5qLWyKjxnZxHRJMN1T
unFxW8irYc/0yH1lkvws1u88D9sbp7aGolZjWrqnRh4yWm6vjkFvAur3HrhEB9W3
8gM8tU58nDSTCHNUVXI/eOe3FHprN5IRrDOoYGD3CPsFCH32JJpYjEDCGfGySoKF
0RIAA6hYsVvaZvC/E5EV6nkvg+3bnuf+yPuYhL/bhFCrogD2diQ7xDozYsvcjn5G
Cv44RKKHIApHEE0FEZ/W3UdKTd+pzoDvmo1jZUx5itoLn756+Qx+LfzZFKsutDHb
onbkdAUTFqa2/5h8KkJT1i3ezcwAPF/ODqYvSWINvvwCC6dGlmGXO9GWzSQixkhA
X74yCp3AgM5qFgUoBkYRhCbQip1hojk93n2CjV2LmXrcZLkCUfX8ZvpH5iEp9gGp
mh0qgPpa3j2rY8XnaaDe+smSq8dtnAYNvk9UTpLL9HNa+G2a8RHvmr/lGEGe7+r5
KpaCjoBIRGMD+bEQ/5TwaZl8kYNYh9dVNjZqJXTctLSuhgU+Eeb0YaHjIcqYBM0t
xeM9H+WK7bKeEkZt3m7rBE/oFcLRc0U0XjHcl4esp1hhrGLjPm7HZz4/E4GT5Vjt
3JoKbgcACfIFVA9yNRluINwkBcMJ8ZXV99DYMVD69XlV7GfBh8OYm5Ma4cQgAliN
e0iyuz58RA8drbkgFz2TMJmy99eworVo0th/rVz/mtHYAThV7wiMtnXYAQq+O1VI
4FY1T6EEBsFUu+5KCY/9jA==
`protect END_PROTECTED
