`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQLlvBji1WGSNDI/7LqdNplNGPH/qjhBJfrbP/p11z7j7i8MiZL9eeoy5NSfwjVF
M2f/sSrndJ3GIk0QvWcmFT/Y7U5UyuSRWexDpLCeunVDaxx09TcyEZtUKsw1NHDj
ZL2/y331XgnitAInC69AeXuPxD2nU8pqH98Pgmg2R3j8nz2aqsM+MsQlNqYFfKSL
4cYQQx7EEpdNJ3+RHXUHeAhBGcq2I3Dk9LgXIr/NJzN9vLPgoMN4pEjHVAO9nOWg
SrNIn1cidm1jJ+BdLIQapwrT30JUkVr7PU4BXrtbXL2vF6WgTxJ1365sMTpWhPUf
RDb5I265TySSfXPj44zoWvVxIhyz9VvzEy1pP371zqaX2SBf9Kd7228oQmxVN/T3
grTtYStESFYm6SwUH+oCOYLAjSv1o/xHl1uRLOG++8Qrsf6dwFNaGBhT+p/1gI0o
s9PRWZTmTkeuJ1QViGsB2A==
`protect END_PROTECTED
