`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pjRNGat/+oxmZiOjr8qkttGxhBwaItcfARIp3ezy1xd3uoJ/4OkSHu1qKzwfScvw
gb0QM4ka6H+vnaZCyymZQnhjeCnwuwIjna5CWBSOsM3mC4mclD+h10qBIHpT0wVJ
KZ7AyadVIx2mVZUXH8otxdww/6ZON4BE1ux9MEa/jU+GK/ZE7WeUfVwtTBh53aV4
qaneRz2+sj9d+LdoSdfTe+p+3bKGomhmyn++VNe0sAHHcbO0vkKhU97nE22WTSBG
CBiZLYiN0++qChEjEYGM/SK98C7NoTu+JAT1PKklWSJbhkldf5oM60FKah8rCTBp
5XVy9Mc7Pd5NTBNmSfN5GihNv/E4xXIBRrsuYDQ9MdZ2kaHMx6nTyy7uMFugEGg6
PFf4UH3L6YD3Gle9r/JUciLVt4QjrWMtYebyXm7d98EMHTLFhHqoq+6Aqr0j34Mx
MAhmAQ39J3bAwRk+z9M4xFs/S4C9XLyXQuPASJa7/hlMjB5A77b+yMMqv5lXrBB8
9HjSSFUK7DAFwloHyJP4EHURmxQyYVaI7tiBE/3w9pR4kWI92k1NGMh7Vnul+Tby
nn2pfZnoflg0DxDntCBhbXMlSVl3rtllUeWBDCmCYRPddrUxIyYsenLUj5Ku/CV6
uvC5TkaEA72c4/Rj4o7QczmNFp4bx5+CzqgSoi20v0E=
`protect END_PROTECTED
