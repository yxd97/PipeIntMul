`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cn0zE7+zTLn1MUWpSRkYnYnAfLDoC1FuEoBZOwlIjqgCKOxtx7gtQEnBEJBcWKd0
/CaaXIZdO5vPpgvawUjzc53aW+hJopD/uUAPMIJsdc1JjkU9Zkob7huylGKotP3+
wcF9ZOt1VRRRK9zttT7ac/cUTYMdEEq/ulLXKMkGZFFS4NfqLt+4Ek768ZzRxq9r
vlPBVucuzPho3mjr5Yn4xw4OzezEYj8yViiPDpeOn4RYlJIFq3917TSpC+ATnqxy
WukoWFm5NeQx0/P1BMVC+qA0Bp0le5IjcUC8WX+eAW8feiSYWZQ0esDU/Kz/4+Mi
rPE6KXMVXVI7qwv541cv1TY4T4BucQHJDEtlp9KyO9KVHxsPIz/xTLBn7HHatx01
Lw6qUrhQLKJi3T9IfM1350X4OER58tocjk5XjOftSnDeix+7WxMKsoq9o09lWIWr
aKTouWJtmT08TYLW3P9B1w11eSTOMky5PWZpXXsEHYulUO36w3TqUcKr7yHV0qJg
IN+r4uMRUVVcvNW1dKp/BcVUBR/ppqKt6QQCi46uRAQ2mtVPf59OVQpN/h3j07eu
/C6L7M3tuX4TbySPZ+c90z+sgnPiMiEJluOLNCiL6Ub7C6aRh+tJESx+THSP2KV7
L0M+dsnXgdjNpmY/p82+2Bc7y6R1e2kOQNBthzFlsR2ILICIYQjhzu/LnDf2LraA
xRKQcmQdDTTAtoquTbksDNoaTC50AugaMXA9qKuGx7Llm9gFQa/suc2gBME887Bd
zVubmKPtKUWu8PzZjAEHIWZwkFmQQnaTNO9+JeiYlqnvJlzo/cWldYqx3X54mfs9
5VCdSi8n8pBOyy1riC2wJW8n1j6VAxiAdI+ZFFtwsKvWHTVsI+KN797q2QEMGQDH
s3vljljSfug9+cOEHAeZbw==
`protect END_PROTECTED
