`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EX9R2hNS4q3BRtf6VVgRMuNI9DaQAoxbV7k2i48Y7iu/DJK0hxVzsXx9BPpbvjr2
C2VyRMonl3VJR6AfohhgUmbm/aLNcfSQW4yFLWRV7HSMPCuSeF6wmzyTyt54jW04
YEc66ivmgbIxQhfZ/3e4NFFaK/8P9kYnAo6qssDCDAGRRgakHdvxqAWRUyBXfd+w
85n22hS5egs68OGwEjicqbF70Sc76oIrL1ByD6/EwoJuMBLzP3yFB7kGNn4f0rld
eCTmnuss21yFJxFikN3DIeItYsQBgo3a3p5wPMPHbzzkwSjFaqo05ZpWvQ2RbW+u
Aei0lPwZcItEQQeAcZBr7uS5Y9zCYL1zf4DI8VRXHyWazzAw1mnvTBO23VQyHgSl
AA5dY2DbfUJ3KkkkXMdeixWp1vUVqwaSpxrg2Xab3oYdX92YJKFoUA+OeOEeArQk
Rzn2bW7h7d/F4niQj+z8NaIBbjt8u6IKlyotROKlbuPcfGsY3ks6zgG774ojVPGm
z8daSL/3bzTru9wQtQdBP6uf+y3AKVbeE27lm4MLI2bZU5mmvXVJLiBFA2AkxQN0
cbtOYP/gbq+oRgZBj4nLMqiYNzH1TLEmtFYgVya27najhj7nb6m7+D+juk420bJA
HjCF3C8Q3g0ejYz82EbrGzYx8P+dLpGwhJUAEfEIn9kwyykQTHi5LZiLAH1z0y1g
YEXe1QUWfT7cNhv3AwC5S58VWOFl1YVaFMtu/aUOH/QqH9aFWIV/zsFRWmmoLSuX
Q6SaxlA01Q/agNd/lPZkUB6zmWpJ8iQhIzy6fScwLQfpnPq+00JUourqieJi/M0Q
jlKvJ1XI1QBz69ETfvJXBXkBoIug6gAcR48fSFlvSbSVbhn79mBQZxnwcwbElfjG
ylFn6B1rNby+kSWWypor4mSNZ/DGPcJGRhRVOCT1/O9HrESqxH+UAaXBqCaWXefP
21/XYraOhYHBMBQ10W1LhFk7Guv1j8YXDFlUNCCf7R0ji2DFQoCSHLeChI3dDMXx
7+wj2JB3Z08Fd+pTS3YoPw==
`protect END_PROTECTED
