`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yv0lJAaFhVVPxpdHruFgofYvXY+tAIQc8qZGQmrjfao4fkbvHrM6txQ8io+XkJna
y7IOpMaNMd2sYiitNMtnIB9yZKJl4VaiH2xQYTS95e2crf1z6lRX72yz6ujTddbY
NR5a72HH1H82yQr5Pgf43EguwX2oGYjKlpleXD/8xZBFTxBdB1Lz3jXqvXssoDxe
JnG7zy/8BKG+tfGQwt8JtpEN7AGiJYJczWY22ooCDwJC/nr+dSJd0qrBkhxNrZ9Q
fgw0WbRhXt6NxtHP1oegXHOfaqE4gWOwBckegTMYlouQNVXlJqNADv9S+ku7l0L2
o72bBrVT9ArQvlFsgpW1dZct6jkIWifLPslvIaGjjWHeO2SejqO2ZHA47kDY/OPH
kXzpYNaxX1Y5NxNTud5WHh1yXrUa/v3DzYbAND/2UA9kM3DRlgcPMBBVSAPCpUeA
rpImft3B38CXeL+wlBSALMM7fJlrKHJ5hlQ3bkEkVgWvJSTZVGRfAgtTEArNKDx8
w74rKYvM/5RGV07UaPs16/Rxyy9/Ow2tSy/8k7LNJfyHp2n1PJlLfOqBHaZKlaKR
AFFKZdD+S6vxX8OM1+d/sxXc6wHBgfWykQxKXwqEKmCUY7xH/okTA4bja7XAZc6H
J+4FkBSTLzTTHNmvSFyMRxWONhG8QazmBmnSZxHgqt6CSvOZuS+F2U/18mNObRbw
dK77t7cU+GuQ7FJxWmwnWVVVsBmnpI/8y9PyTxS95vH6zmtooP/fBxwpBIo9mzg3
Q+MqAUxBOL9kyjtMqhZFVjAN5a92aFVXOnV6TWe48/j2+nngjrPgPedRgGaN1C5z
eXlwqH4suoy1D1mcDeFvkH/RiaBmAY6dx5LlhCdG2TUCpjET+3nZ9E48Mlh+mhio
r6KqxxgElwaiyaT4t4NC/k5k18/TXM3eWsTcko0QSPFa85PYntLP/444wYwQ9KjP
CWTUz8fmbU1k9vPEBahhvLa8194Y4NPe+gSmGfByc7Lil2hYHLzDtBiz9enCVhqn
xO3ah+S1UaS5uHJEXgH7URPPtOVFSlHjymLDArkqIXLEmya3/S3jIvELj7VskBQ9
dh3vQFqyPiIOonPNZdMz+5tZKjgzr6G5s5x118MX2eW9D3Yp6200Jsn6lBYXbNyz
/LrorL68XgqRRU98pluy+0I6efOBvIIJGthRrFrHyVT/7GUOOW6AHaRXYhx1bwSW
yAEA+pioU5wmPerK0jT1YVy1tqRNSMk5tsqYXno2VMRSxLbdqgIRgFQZKEOwTN14
XGXiwVyjKqi6/59q7YpkGiGrRi0JP6eOesCd7P45Cj32hUyd3ydGpRUMopKNsPkt
8XH2rPocS2KtFfmGytRlCHeKUHjDrPpyaZVOGbNuQEaKyVfXesZj3Dwp5uEiNmMV
OKxQ0WOmTggnRBY6zkXhdA+kievFRPF0jrlBtY66MzPHgYwiNQSJJtaIqwcArS8b
I2NqDv8ONufi/nE4jZ/wA4+FS0gNb/D9a3nu9aMutRWnBnw7FxUFzO/bVUW2xAH4
n1ycK8v6a+7aA/6vhWx3aJdBXPaiCFjIyC9O2XSkGtoPlWA1ESdEN+wbwY2vlYtw
jIgCk/X//0njOzcBJWMrVK0ua72gBdE3rHempEy39txU7zo8JIiTb1SwvJw/iXsI
JO4VGMSKOzTAU9eyoMt/ou8pmZKgfQAvNPDHjpPrh/eNSXLSl13cg6KRu7HqmEwE
Ay5m/bM0X0ORZBw8WnEVtoOpNs/lkCmQIGWuGXa0z+i44NWzAJ9O28vLSNPlbQWM
20PWN89xOJ/kz8VVaxypvhrYGfbOmWlrLf2lc3cHqRUev8ZBpsFdhzNMp1BfZWQK
Oxpn2AXz+F8dqsPHxDvOTd+h4CrEjAUqdQyjD007tRPOZN1BEEm9Mf0jWTEgJrmt
bMK/cBrozAUhOYh7L3Ncqjtb8AR3w0UvCErJfr2E+ZoYCkx22Hawp+Fn48lqecu5
kVVYWmivq90772d9kf2v2iIhXie9qzJqt9v0AU4GG41NgxEXYLyZ7uIqSVyX5Mld
4y1Z2rw3VaSQh00IThLgidRHsOiBp6/i31Dugr4mWv6lEL+K8VjM1CQZeZS44MhM
pwsokE0kEn+JiC2A6hwohiDtMnJoy9zKNHyJq0MTfTjUwniQe7c+bzjXfFwC8SD4
kbxQyXRerUC+QNnCJLd2h0ZVToguYtT+vzoVvJS2E4R5JePFz75TU+8BfPkpJpnO
A4Sy75+iCcl+jARGa94w/5CaJOt6b9VkKTP25GZtsz+zg9sXMxWBXUvXA7jazBbW
qswVZ+I25D9LGYtum9FTwCGWvYJNhJUWUQoUeNpoiTLW8XO8lCaQHvrm9lUgnchI
O7KdudDZSaPDh9s16fupF32Z9X7UkQTi+r6tjMSoa80OzMHCZ2qLslwGDksqdJOW
fUTgja2/9cMJrHctALYrn3bydwKPzG047FJubLumxNbvMR/2v2gYcnK3z8igOTOV
BtaCK6HwaIxouEu1laW97VHM+JxMP+lZ5BJgANgVLiCbceQSnWFvmdj8SMtfBqCx
hPQeARonPKogy3ASoUlUC02A+9o4fWD5KNnYz/m2BwUwbSxhpOgqrcQnCHyOjB8k
1PEJ3u6Xz8/GhqE4RU2O6zjSm1nbG+wUW9f35qB0xlvkxB6BDDBrsp0FWYBjb1Xj
AN0dOLpqla9qUMZj96u4hZT870L2PKJbRbTQlsntEZXnWK3cEQZ2RI+L+1HEp7oA
A9GS6FNwtiqsCzavXLKeLyNOP/Jw3M6XF8vACHrBDDQmyA/rjsfK1y6Bvk2Ep50t
iWCmtzdfdTJ6nHFhw4BQV9I15BYvqGH06VewL51Jps3xwK63GQQzZbfnafdCTbxm
VdReXbSY7+YzaPdp2OPmR1ilRfv2lb8OKJdL21NoS0ti4nJ07ATvRlgmHvZLTG0S
oCAawI/Y+Ntqz+f7QQ/WqA2qwQsf3Kthu4kxXYdnR3wBqhDpFDpyjR5iPYkPzBP1
AIAKadtN0ZkF1lBJJzixtfx0JPmf+LOJKbIeZXbSMRLSL52aRiwKFuE12YJNvutq
gKZgMGBpWSn+QUYRhWE++AKMKaR8iLVt2S2MOTPXT1lQzsOSNY90FtwJEGzRCpRO
LCvuvgsuPp7eClVt3kyFmIwqLMMzVp+dcaRuk3acezL4U738YEb+K1sEDyyjjMnC
hVdR30OXlaNowjVjBt4AkkiGfeQW5JVB+YauqH1WS4nL+F+0rfHFu+sl0zzmDJLJ
bye0oWcr20dTllQ5/iuAkQVEizwag+2nByBPnKqs+VMTTRDpdVMnfzwaerQ6ZAg9
fptGxzmVDV7tMBz89tj23C9k2MfxOaZjueBpVb0TCDgSI68ISwky/av8IC1p9GBU
bRbh4BmRxXa659fp/9Q/0QaXu3hVL07L2yf1E3ayLPv50Sm6AY7TckeZ++UtanGW
YIn0tkWU9Aj+MCQ9nIIn00YNg0DAtdQt1r2jXuo1JTPy0X0LfpuV1NK98SEDn5X5
0zcWSGcEBgFPZn4zrNKvFOEFBgebmjHvUlAjdik4yVj0ZlD1mIdIZu9QmMPc5dtN
JaAc5L2bGucrbtb4WKd2tMLX29xxa8Ab0Sv6F/S+DnHONKqvekXlDArATN/0Jp2/
FEqtal2s4WBYjerUpHme5yj9jcmpWHUeIvvf48lJFS8GwcifS7KaxhkAz2qW8Jy5
af+as/nu4zGvCEqDsC5tpkCMTj33uQ3aKMsl7T7Z+44EIrku4M4zVEax/YC1ZBdV
OLYenFhfZ93U74O934iiM/tA5Br8t7VXcNgujUX/otyyl7ZdNvmYGdPAnnBlB1GS
gnlPk+ev6t/Wq6wPmYxJ1y3371MutJTVl8crdqBdKY7oatfVXYHDxHZFWqPk0Mzi
5sqPreIyU4o/ot4iLUSjw5DCZSQ1Rm4+WMvRfCADxQCZUO0yXxs2wOMYyppofAqa
P6akooQqudLovTXWSfAnWVtAkFObuYrTFY9zL7/1WUMQu7D0Tp/FWhZu8x1IGx26
ZvQ9CD0WnNBlG/w+axN5M0O4ZJzIEPJpVdnYO5qqdgSwIvEW1xJm3bmysXDwX2hC
A/8DyBdzlCyj/b+sZ0AvTSP+Gp4ZR5KdZnR4Q9QstnL/M+woOxzQWfFtJwfhaLmJ
K/1r+iybC7knyVdp1puPrrevQO5n7z0mfuNn6xI6SlEkxndYa00TXeE68dJxiqoY
AB5HTBOcO9xwOhLgD9wTyd77smqt6HodS40QK2d7eG1l2YMKWuYt5kqG7hsB5a5b
D2S9igTRNgnc4zUHSbsrBF6YIGxilN3+aOPDHHucDAeD9kKqbBc3KU7VVfD37qcP
qcYXYaeBPClH347oZbW/bhL8gZ36BsfbQn5/ELhc6sKdDFaPQ37MFjZ+XFBs6rn1
zwpaHe0eOm8JaWetQE2UFg==
`protect END_PROTECTED
