`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bdU1190l+bG+8W2/P3ya2ub48o3wRLN7PZOiHcQj8hfKU09D5JKSOYHvVpiCjz4n
A2Skoqz5fvv9dnsiyI0UquKA8S0ApMBo0RHOmHwt5TusrpVv5s5X3B7ddlkTPmlK
rcADKzg5tjhypmXff/AGC6dqBxEFHR1Fr0RBIsfnPqvfH6sYFAhc1Z3BJAzj/Hlw
JbfY6deFvuvJ+iOuqC4iy5EtyN1J+VUMnh+lIy8udVOa/0TWpM417HLmdPxcMEII
kJfbegzzWS6ci2CHaoRQ7NcNuN+EqEXMKQOiYoljtFnKtns1dbiNq1IYgyswQbv1
`protect END_PROTECTED
