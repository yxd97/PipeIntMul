`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZxopkwsRjQCKEUhJ1SEC2ojbl4mxq9eIFTGuoaWUDvXQqXcSDfzKWpdnqn2qUgw4
xOHg+6P/VsoAzvJcd+bJH7f74RBKOKZa92Z30H00ksgj7meFx828Ghs2ZGzHzXzs
WuHWYmB9r1J+76inrmv8w6WvQwDS9Fk1L1lWZGOMslKvCg2LknVlvnM9kfIiniev
xwJwIv61jsXUCYmLZeCRaBIfb0/4W5XSYIYVFa3FVA3eH9UMRjYG2bh2T/PAb4Mr
q0FCOodqBvYOFeH3nptPFkiMyn0/53gnwh+RZZzlg83yYorzxbL/rsYUthD6gOui
fzGai97Job2P9NLUIiIQFg6TW0FI5RD6NOD/zmxI2MEewETXLXCgG8epixSelxfl
mPO4kw5CIRroFrDfmDk4rrug6MzdpsgfTMwBbTjxNzigc6mTJF49pX0m18HS0qgW
YH7gI3Pi7nRnEKe6AjuUH8RVetkQXS5rwpCswWWvQY+KXWAOjE+tujPkIJ6jDBhM
4xrNCD4Wx3jC/x/0GJPLLvYhHNVY3H0FBUEGEOhIdMt++mMNCZZ4BSsAqRUCRKSk
edsYCpTv0CVuY/HoO3XPdyk9cqfS4AEc6TWYwdj+XIUpV9AOGy3f8Oa1IUF7kpWo
yyhP1NG5JwF78WNqd44y2y1eaOxhDAujV3WU04chVrTXdshB+qh+HgBusuIMNld8
9KfiggXxZXp7Wx+G0yN/6GF1xbAP8fgC5S5i6Xmy/gpw3WIWj9D5nZlMVVBsqb/2
raWLrwEIfrdAdyKG4rxY0XVs6KqQNgskBA0fHrOYLwZ3EerUov31zJXkz9P5Ko89
5EfKxknLeal8eAnIBJ/LFiT27jgg++LBksv1R2vd9NUYR2jy83u1GwCr8xPAWwC6
S5Ug+badvX0KCLQn5yYmtw9hVkBGayUqKvzLMunbFsBnzjMlVmdY/zEwEd9BSS2y
NdkiHh+ma0x+Hx0py4N1eyXDVGOTOVfeWaL3UoewdMLn8CyQN/734onI02yhQen9
1FVGoo9dqlg8zAPYdOOzntf5oAvS9GXF6IMoskg1GF671X1kF91FK1hUom+TAKUL
pXgJ+jJ8mMniZ0z6V8BJzkbo7QllXscUDOLbmgR5K3S9JZeWnlmJcG4JGjAC/kDl
4TjhkGm6JYFQ/6rz9bp6KBNO0y0R7KPg7K5Q9nXKrU1i10Pd2rtyIjRWakxbfc32
g2h1Micg2dvSiyPqEVufABmrM1h0QJLNpMCJbNIPmEXqbPOF8oSsLeVQLyeTepVP
fW4I81aGyfoUanS6yTzeaM0wDswqYm1OlsisksduKDrtitrA72eQ6RGb6TOYNUaO
HyOieNCCM/YgV6ZE3huMPeFZfFy618qP/kKfXAepBkd7RCOjbXYHpk37IBSe1irc
hgPKVWVhL+RYXJthZ9PRdVGebkGIWJbssQB8tmOn4a2LuSFgQiof8uKznnZY8NjV
N+JeByxfEpFyxwYo8UJTe4oZ54JN/D/efTaOPjXyiF3mP6tGI/1TQGWa32vKoZQa
Ir/lEFEtqoL4eo2nOiCdWFNWyori3ucLbuqc034J47njYeBjC4Ht5Dv7pnuz0mZp
GwYrWS9w1kwLqL0U040QyMFTq/A9BlcNHH7Z9S1yOBFEPS4J23NVCWGJPhSqK5z2
Vx7tMy4Oi2ed8UdKiHuOT0Q079cWx/NyrlpCC80lHFIS47AlVL09lQHiWM8rnDUM
bhAKtgRQbTf6j1X03er0/XeRNkCIcXmSZDVPJMbs/6Nq1rH0m8lEHsY1wI61sYPe
JXfm3aEmdBQ8cN//qxafkBiLYRebNP62XzBFOllsP5I/Iv8Rnh3ltezhQ4iEOTDO
pdxfXPB2zzWOTqd8fzkZooMGizNF1Xj/JIgVF7KwFXsg12lWS5j4ZOm2M41tmQZW
94MUcMSTZGsPoMCU/Rz2A+pm3rGfM5uhzI+oxLur9cBQVBTnX2x0mmYMDDYRbcI/
ls4UkCL/swXC7Hrge4Z1p3fujKuCG2ig16+55ralZSTC762hwkDVAeY9ysC1NCSw
pATFGehwDJzJ5WdRBsDqlxcjIq5Uc/CckcR1yngZgzEaoKF7dodHLQNHvQoThjbZ
D3jMAl4BhpAY+sWlfwUxznqW9Klq2hgccT9xpYfyoA8UDcn8IAH7mDGx8FsoLa9O
1CliuFSSNN5cZN3azIeapdoAcGXONpaCKFDAbe+yVPwrRY+pb82vx6VAgcGj7reB
i4bDzJfkN7NVUDk7tnJcdORvnh/TRObboT7bWkPDQfB9KCS71ZZJ4L9c+oPB+LN0
aoa+SwvAG5tQ8m16wM6U2FmXjzeAkffVBk+OT92JWo4WVAC48iFcgAykn2sLZi3L
a4i2CmgBXX2P7Lk2qRE9RLms6YRFvA3+6Kb66kq3kGlPHCx3yOTFanSdzPaCZs0A
q+G5HGK59b5EWP38tjc/F9flLsaCNAdsn511VBz2cV2mW5URKcCYN4bKv4XAeCFb
yDj+19lX2VeisrPbYzLci04AB4Q16srDA9iYeSuzlkOlxCuBxcBf4fPBZ9UFbXYd
e7gAAGh1oYzyRUyGxkan+scLwKRl5JNGn62aC6jBTNMXWCa5PU1cIzO0eLUOxqpz
lgtdTfr7+Gp7/uQwNP3oc95mbejsI2+t9Xcf/oknYFY3hdgZAgcp8h9jn+g0zFMU
JaxriXmraCoMDLCyklczE0lIgEre6ae35ROv7x2k6zH3N6yd8bR9z5NjwRYrLjg1
IR95FCU7/gOfRnfIYTAqaA==
`protect END_PROTECTED
