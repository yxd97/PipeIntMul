`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tek99o52fs5qYYn7qdILQDIVz1vfq3Mmbv39/s5NlY6DDA5Ef+Wou9jk4ADWLQB3
xagDN8Tn1tVWtPng3/hsKGFmij6s0vUO6TW1Qnav9sFykrCXRSMU4CwGbmnUr1CW
BZ2KuqQamrVF4sZh0tnr+8LgqryV7UT4fKyGK5sJWw5IZTXnY9HTR8/DeYiUtfgT
PcsCgpXU7ENDYa4bIcmrXTVHJUuz5BkIwUrDB0xuHs4GNGohNHnPKR7ZZDud2dmm
Q+pCcB5CWjD8GQ1w/Cnfx2OyxoPfu10JtZLh1EGEmCD+QKCbdYujyCtg1dm15iQ9
FmHuyLwAwm8xUCMY4o4kAdWG/S4D0SVqFjwtvO4FCuFOQgwZCMeYJd3+fB3dysUw
t9fSvot2ytodxMdHysuvChIWZf7/h75GVe0JUike6cJsJvkiaEdwGI4eiFGjEZY4
P+rPXAEWWtPw7OWgpQs68QYM8DrsNnnkxt2vns8zZeweIOMi6WoekE05M+N8vNvp
`protect END_PROTECTED
