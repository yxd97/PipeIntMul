`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OK7iB+bZ+AVoDrtg9a1NXWg8vnLJHU0zLwm2SQEeFXk5kuS+AdrN98Eqx4atixTn
3I482Lwo+KLqEmz7SP9XCpghjg/hgBSEYZH2+h3oDHZsQPogzkQYGqtylRnaPTtv
ywi0fAUB/w8wFc3uqYUQpAAeChpOqY2Sivn5d26n1n50G+1ZewPVfJHQiaawKcTq
zGXS77oiYOyL3opYdnn3SPCWlDYYcm1XqXfl79zenDMPUHLrtuxV3mNof47bSX3i
c3fqLvnCYMtiF3/0Z0vUblYWIQ5MhqQ9HercBmMD8Q4jzsQ7aAmyjBWxrm2s78Gc
9amIkgZ3OnsrJqXe7SFCMjlojG7lrk+GZ8IHfF5d+IqrTzUlnozZaA2zWiMQu0R1
H38ChHfZYryILDUu/HbFUS0DqMIQh99KLCKTYeleWDjZ9bGGmR/nUrQuFsjcPYRj
o7hAX3zEeIjZ9D9V/cnq00MkTVkXR4WZMATe4bChU/MX3hfzZSOt6idO0jdZ4RBh
PjdufdU964RMJurlwau7Es0wpsNBTxcpvL30pLJG+P+SwF3k4YKgtuDTdO0shaa7
4bkIYMIKiGUTjfg1wrqo74PE7OIhjYldL+sq/Sy3yJskcqUIaX/zjAyY8ZFP7kSU
rWJO6TyYe+FLxlECdBpisbfTQ6xHFMxNk+ciLVaR5OBFGsv0prWPB6MNA0wI5oLK
DLv2B2wrN0rAK5aneomc/+yZxkOjhnEpizjdBS7Nb7++gn7folMMZOz81adiAsJy
DxEj2aneM+IB+40u2GOOTAJPY8JDDQT+74oFsniU+UA=
`protect END_PROTECTED
