`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzQqeWmb4RKdRh7+1yIlayR8/MSpw00PGPntbLIY5O4vqqT+eXHAX94HGV0bXgZV
bSJGZZSUf9kMN0YxYIyJew1Jbk1gU5nssS7rIlCjpkbqEBKAQKnbbP6D7Mtf9++E
Sz+TExl28Xmqb0R00l4BM1Peu7kORqjjgyXm7qFOrnVJGXzqHPbUly5Em0N1GTaM
8ogfInS+kChklHzM4cw5Wurdi4j/y3Y1Ic3k7RWpOoHKNqAmaKhV7My7R71pn7Vh
ZKKYhfXIE91i2hG96EQqFCsaioVlz31SSNQ9iHWLWyTFCDpJQRzuAOHa2IxSRViF
VxdQmnOB4iq+m5kkTpKW6dUdg8edgXDTwqsrOGJIvurMyg+lJZcUJYKl2oIds6VR
sea5ASyz9dZAN8tMyPqdir+rBNRpclXAbWXqClXlNm/1E5NuKDyqOczr2DgR0aJt
mwBRca5zLLotpPX3IoGFSlK3R4ND0UNNITxfW8aYU9Kkm2B4EYcUm3SUrnH+sJL2
LxQdLXLxpLqQuCOFqBtfUCFkOC/ijKmMxxFvXarr58hfYAEkAUTEXEhF7bO9u0lM
`protect END_PROTECTED
