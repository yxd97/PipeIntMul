`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4SPbMjKsoTA4GudY+z2qRtGRjWoGtn+nt+YB8eqy20BfUQ4fx4z+znrVM7bKX3/c
rEt4HnWKLhNdbyCKzpwS+wZ/u80ErYTndDGxU/SSXCQKIcGtEYQa8EB/k3bfLwnr
UYghlhcjJhFhDVHnA69NwGoE5pTfGzKfr5WNGcXXWzoVRA7d6uzFcllxiiZHXBK9
vMK8s96dAvoSO7iVOH4rS0MA51munzefhEIE/HMhovSI0MYAdtqN0Cbls/zfK1nO
9yGV+i0951hdzpQIEPcYUKe8aYVNkbC9waf98reJXoCUESyALFUZcNDiN7gLOQQH
PppNI+KnZPVm9QN9L7dcNjZnURCkFtbc75uY4ZXjstUPhZgPde6KUh+OO6X5acdY
sYM/6NDYNdbSJnvFjtk+2aZHPSXOf02cI9NMhD33kxgahRQ7X5qrDDOxEkAx2fWS
4qdg3Dfb71OvWPUP3aiiWgwYll/Lx/7C1wddhaTgv6xUCvRF9OocXkogJJkvR2Gk
epJYF2QTTj5wGcffbKisSrr9r2sNb1lINEJEh8gXyR32qwsecQJkGPhrBda9uhSy
qjSiq8bin0hqbv3mU0dWyD72L0CLGM91ePYX9OTyDoKhmaYlMJpTfHyeKIphXwKg
DsvNpZmzLldjSKK5oMepVGgfgDgG3R+pPe4ggMjBvqg4kN4rdJij1HBEgCeAqZJg
cEciJ3QkJamPlHu+2psMAqa56FBPtjWNT2giorMglWK1CnSgdnOplBPhroVaqCeU
fiC+tmRKLjEchCuYVyi1y3iAQyhwii912tIi8vciP1wlXXA0Ph/ZaVS6dj1KlIoK
3LAQaYYGmZC/cUcvpI2PggXu6rz71w2NfqIP0wiTlzYKwhIUlOpdUP2u5RymfNcF
1YL0QMKnWlbz3uhslqOIJr3rNXEugUalk5JgLpnet5yjCKO7m3v2RDZJ+rGUwTsE
Dc6aBlSKFEEgIt8KYS1qG8JEUoYRvw+0sJ1uB4VJ+w8=
`protect END_PROTECTED
