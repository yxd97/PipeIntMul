`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vbKzJ3hej1h+aO5CVc7nM0G/E/KXo9I+/nO0D0WuDonh6/iMsX3cwYNV5m3mmnd9
+vSIbz2015n1uYUsvbtwSxuziPdtyTcrDZgXT6MydtABc0T4dj4BGq3PC9I/AhpW
TpZP1QyvcmEoo23j9fSS3E6wAd199xpkAaYZpwlO5rpdYBJgRrfEoKR1dw6fXjGj
mvReDaoYBQhE+9RhZvomt4lxo3mAPejuBstAQVdxWDyucFZt3v9LTzfuXoqA33Nd
KJHAxXXrziASEfMjd83/efJ4tm0TqlrZAF2DoTgxpjpk+J84L/8qYR0tiWo95OuM
BubpxyJXISp9Q8aJGEvx/zVSNr5qd3rMj4lKCUmObDEtpkzzrNDzrS3nFURuGY+z
pQoeFKOlpGMBYjLVw2ETdvw2ztkzqwD8y6R9P7RGHR7Oql+bO7pKNqg+ttHiDJZ4
M1MN0+vkecLhYbE2aYZoQml9M1FvjmBl/TgpmO0wqk+l9vTWYAuveVm08baNFd6p
goQPMLkp6L26zLe8o60bHIhAlyXBuGgsCNEZs3B3qQnqq1EzRU1BZpU1QjZ8vxXT
2Nk4PuoJKMoOu/gPPZ3eizjOuzfceyS0BHaLClH7LIyS6Jlqnaw1b8d5VfiE3kOK
EKiKnMHhUChb/kO4Eon9ppXxVWfh96D6g8kLKX8WR81lt1I+PDRPA/G38hx9zCig
gTMVMYMEHvQ6LPcTTG4yyc6265gQ4WZv4KQ2cjYlmnvuXKg3I4iK7pXlxZaPuKFc
0ak5heAdts6tKLW3pPV0VsB7ziP7DKkPPMCNtVnHVZLnw10nayA0AaSoEN91jhap
F3j0jT5t2t6V3N7WYIQ0Jo8LVzjxUEWmv//0lDsc5K3kfAZt2kIzOXsU14H8w8ti
DR6WYcRy0dOItpFuIHai/28pacVp/D56Vppu/GlJXaULYvxxkYYp+syRRJT2OV9Z
cTXKOeSAqvXh/OMY/pePl8ogojRe3nUziZEesHyCu6rpekeUQ0w6a0Dbw0UC4i3L
fu0H4wZe3WjLk8H6ao5Npi4RFLxkcOv7ss1ieF60Oo4AvfZ6oU2E1wid7EfgHC8a
u2OvZUurH5WqHKFvKjhusl0SvbFeRn40ThRfHrmhdEmo5Dq1IPUrF8CAiGOw1xw7
wl45iLqWfCdYekBpGe5ycxyr6xBqDXo7XTR6oOJRA+tuOLKHQeob08VKf5XffF84
9vqHDQBtqdkdkRBjEOO6LMF0L1pNROLZZvPi25pjZZeAbRQ3gxtHe59oUaVrCnPH
0sLLN1mspXJ0Br2oImsQgaxHGsNnqGOmKCD+jAIc44C/ZjcFMTgy4M+FaJdvN7rb
N3im6RugzX7jZhCw+rFTBxHfAnWr9YQP2s2j4a1dUm6c8VXawS6xuFvl6DgyFkwl
n8LpWPhKnZXLfikaEnQ1bW9CT6cc93YuAefpwkW15/n9gd8aEwLlfOTlnyWX0zFM
OBGKrgqMdewhCPOtt72eOYrsr+wL0Dr+C7apMsUJ6/Bs8XLoKkYkgqOg+mw7OXNG
X2u/r16yWWm4R28aFpYG/QRslQkMaqnMOv9tGD8KKDAhavccYkM854CECFPGIp2O
NmsPHuGUvYIfgOT/5YUD/J98fX+eJ+tR8cQzoW1HW940rOo1jaYEQnYBk+OrTFfV
jof4b3qWuXCSTxWtwaJlhWkfdsq3QO832UoZd88MbxTD/tWXL9XzcQQ1JHsaGmse
Ia6YN1g5OEW7TnUsEklQLQp15hv4O0RMi8ZGjeAul+qVk3TFSQi207zmiv+dnIq0
MmKAfOOl7rf1GJAMl6iUwSEspIOVt+PQtbdri1z6oDEkQmEiWhmU9zeLxh4TC8uK
wYvfzYyjgP2qum6USJLfE2MzygUzXM3G+qxCFR1ueLiNQdN3wqsl/BiUR2DqTtH8
lfPB5yjRhwLD/Fq2mddXDkL022Xz6IXRjNyQ/J/ExRwLjhV0QymhLHY70u1uDCBi
/+J6qQtCflDWTKTBSfBfGIXX8mU4L/5YE0/dAtJEFJJqxFefLZR2ZcQ2k2UBDszN
TPKRSWc9x29sLmvs3/LkOJvSLFuDrWThQUQ6gu0TcRGqKjRtYj8EMLdenfYKqHgr
BqulOHTBCS7cuWq9mikLWhhi/rssy8vuzLEc7SVZ2lo5lZ/He9p/4JNv6tSpciZ1
Uck8YfCKVaoN8B/LDP2HphDZl5V87Pi+8pIzSGO9IcSv25KS9qGxQtuKmIIIbD5r
AllonljO1mmJ06p/PuwLNZ811y/lxQOO6qPcudgXSVB8SaOAEtrz4gv4i8OLjFKJ
zno5WNQGKbohIa4QA/gz5v6PfkMb7J4kXo1MPuLaj68TZd4/i7asigGz/bpEep7C
vzDKCBTGiUYY4w4iImhpi6MXlofQ1moxDqezacT+4PfB//ZM3KBjgJuHVdT72Hqp
jYLdDNolK07hjEShkxXzf72KFCJn80oLRruIXvOb1UL7VSLG5dpjiO1qpt/m9nUQ
eF+vLYBiuN6ZrzIc3SmVqqEmXPuSoEEt67ZuhhiE+IFmtiGZPohbo8vMJimSHWLm
/HI9QGCWY/Z4I30BX0FoKKq1/Y2A/RGgg9QJmVK8QTmYWx6k+FEntZ0msDJyv63a
m3b9+YlA0ZDjFZpYuIeOgcROaERC1roF6yDootQ7mmlXDdM/VtQRhNYRPsQStMpN
xCfyQP05Ghwp8ZcyTJ/h9yeW/zo5ZliuVk1ufcI2doR++zUYiR9TheeLJIee6xmP
05GP2YfNCZ/piWgMmodh6rb+vwaA8vyk2+ofAt6a0t3rmJDyMWHXLjbjg89HLNP/
MklfiHP3fTyDj4u+7CKm/+7ym0ZI8iHr0DDrSrZ9tJSDN5REiZ5ugd0q/VX1lwBL
lwHq/TqueCaxWISfZVWwhVeEsBzTYG5W/5e0KF5jMoeFvL/PQP5OdoUdXmRljWEI
8JZFbHGmg1kc/PHR9BerVc9mdvkcC5z4r9PcfoEj/+3gEp/4pnY5aGdpcTi4rSD+
L8vnYso6/MlbASZBRV4JaWjyKum3oU4gTajXEeqa1LAzeiYm3Rc8hMquFCahVZ/Q
z/l9yRYYUppE5FLi4GSurf2YKNTSKtJwia+Gtddil277UsXp+8aPTmJB4aWHIj2v
HJuAjqKn8cVeisyFY9zNKBQtq6OUPcVcohP2Js7YpJCrT9P46U/4O9SdYzlzVxm4
AmzEMKotulWog6M52jH+C8sJRcufR3MI/CQ6an34swqhmVm30r0dQqIl6w/SYhAK
AqeAu+JQuUy0To3V6BnSDQtIG+gaB5/Bm1dcgrsL5lXZwyUz3QUeviNgqDJmclRt
G8zYxXroBr208/9ZeG5S4TPEmn0GqbMY4cAPBSo6LEbxiU0dr+P/uwZTJUBNUfUU
HNQ7JKukp/J1PLJRFYplqYE/rmgytmxv6LYjd1wP+jZDOhKaHwcJ7efBYfkSruC9
5lk8RtXiBEqyWMtgaytKnlHaDn+5w2ihWzUXS2WlvKMnjbpw+6bVHYLee8/8NmS2
mfafiOKID2bEndtd6J4yza7ntqXruPo+BHSEj9Y01pQOhrmEFoJlvAym+E8XdBgj
yX+GuSJ/ivhsLlciJRnaory9h3HCU4+N76DFGxsKj17CDHGzWnvNnxXiOl5j8341
5Sqy/90uPGBbWW5Bb4ehYORucekKXdiiSu6rB1Ku9e+hxuQGV8R/lbDNZN0aujT3
EonTHBSfYzS1YDiFZ7a0h08Uvk9MWIOAEQ9grsXNE8FqaTh2VWbrcM24655rhPeg
ed1ENxJicXNW9+LoRvOUsipPDfA9z3c3faEwtgu2820QT8gDgvT9Ay5zZ73htgHq
uxwcwlrwvI2Pf62lAtJ/1F71UGmxU3TcdJiipfHDgySi0wlgXa7FBssSl9q65U03
M2VM8vGMsg6SXq9lGcb/iYFcdsYQjtAITRJeSp2DvUe2MGaKmiLS9wnIOH8uLwQd
c05tsJqEMSYqTvetMwdgQm7cD5CLIhjOBz+rFoxSI1EnyBxX/10UOqEiIUWRwvB3
HrIuqgKPpICNgQLIOwTEO2Jyb+5AKyf6rWdqPGwdsGpKvWm2hW0GMdcQjhQJxWj3
2mDyijWZm4Xv1goe5i5dgter8iu+hglYcbOhrolAHm+1JHFeUVTCAkwTYpkb9GLa
Sm7mHu4HSUt+A8VggKN6VI7dQn8JHMRd0PHICMW9s/AmZ4aMAyP4QG4Ade59VTOb
js2tUxIv5DVA3KQrj1G07jN3bgTNk7fe2mUpSqROUePVg0MQFIYWNqW/CCQnLI91
qvgWjEZi+f3wmQGY8YjUi1Ab8iKLaW+ZCqKlWVpqmP7Y2eKZt5rKVquEyj/pbygD
53yupM3SVPO2mL1RHzKIuwTupDKhPWmvDfY+XzSVYiQtYj6tfQtUbWcsiXfMM1YP
nzMAD9WEyulWQPz9+y0Q3HK2a6IVprCGbA/wQwQ1515XOytNDJcgn0PNImFJh3Fl
LPYjUHOY7HT9qzpbrPCbUVUAXLZPM5sVB/TjcmnbAUPbMzglPcoJG5OkCMhpbFLc
ZtNxkWkE4F2Yk+eZNx3ILYhkrcWDdw1NjMfN7d0fDYe4Ci01Q6JNfijx6H04fZJS
9lsy0rT3nYfLAXGr5EByYs876GIPavTVfXsrps0UGtVMnSSvUkFHcvXupwerVbI0
FleyRftBnNmtjtH7XN0E04FsU7M7mY8hd1sXGmpphp5yRO+zJITZebEaFPA1Zm52
x09h515g0K3otNyFLShGGhBYwrE32ry9kzaJ9WMeZRdYys1q4NMSvN+6D31+aJHW
Uw++TVDs4vCKENJ1bs/RNYP6YOl71bFLaGFcCZNJpH1zmhOlBXb2xyfzWTwv9G6k
q/iBQoUEPCV9FD4Ebk2/GqD5xCB/QxKyJkDIQ5xImjTxRLld4+/yNzUNyfm7d4Rd
Zbk/x0jSAROaSRMZyNyYTG1khaNk5GJAG7WUtcl1iUk=
`protect END_PROTECTED
