`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdojUFZARTLno6yvG7ING6lhygKegPRs4b5rfTibJUx0Ilo/vZuSZHYhle1k5mCU
lMiV6rFGmC+TEGsWqy1SZdFPCBjcebc9cnVjVLsld0eVPvoP1WpzkWvotN73gFiV
B1avEPpWu45+qKKPFl7gt3zExIdxleQscYhoSpkzT9y//jBWwUWS5YIhxpLXsXbg
PHqyZzl/epg+F0Cft8/zci0wV9RPN6rfPk1kRSRCP6hHhGrQs41V+cuTUt4gAiaa
zzCByxLmf/BcCD8lln8haFBFEHxfRNK2u/uNZJ8OqvCKm22gb1Wk5TJNA2ihGM7v
7di9VGV+V9NyOGf7rt62m5YVs5K38p/RfIA1UzbQoxi1KaLyn/yD45yh5kx27QBj
Nlzbjgcm7UexaWol+zOhdwGpfKRB2pnZAl1NWp58dtxBvUG4jouY58DY2aHGsceS
yeWROF2OeevEakMQcLlZ1H3//AqGksIZLzYEooLjG7GH5L9ADxWBLZCVEK0uHa2A
xTIkVmyLoPTkMZCLf763QkYhNSthVSO/Ofh2M/VrQVY=
`protect END_PROTECTED
