`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tMkG9DHSe1MSW/d5e9Pzjq9gEC/OqAcTc83QW6CyyAXQ2DQ6xTFuobvkMimBzZMH
RdDPfu4AlYT1JFvyN8PvRfHFGdamDNOQb+iA/InnZ2TORuuGX7+mKcZPjyNaJuh3
9ALNyOZ8Dxe8IWgOT3m6Y617vTBLPH9yo4hC3vMuRMLXph6O/3WZQ39ENqA7upYz
ni5U8BmiRHAeyeeSzh6dFk/UiW5Nc+L3pgd+vqioW2j5nfVhgXSK0HhEZvmtxyal
`protect END_PROTECTED
