`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8qjfqqYMOFJdE8P4EQQCslc5W5Z2c16m0l/mH9tsE1VVV1awSGXVAevEKJD644R
a5jvebpWjgaj2Q/SYzv7M16W8hpxeluQukFZQQay4L/cMXhwLyRieUkzs8bfaq3I
61ZYimPIgg1+SpBfvs6k8FU2qoenURFIY12FLntw8yEWK9D+zMkcNs4vj4PSQqdN
6g0PtzXJcoOgV4exbe+cYBa2RPCCPBe7sGcW0YJUMBZK9GY5Mkb7DJUnu6gMtMHp
Aucsy2qXTJNf6Vrqts2ak2+tMxbJ8GyzlEfM+oi37uSAI0A4LSK8c6taGn7gG0SI
bYKV99UculvZCuBgryMbRgOmpO2ElG2VF8OrctiGBEMCR4etsJUNDqOJFl/NmaKK
r3VRzpw5B01Vubpf8s4O6KXxuCZWYexhEiNRvksp7YSRNYMrv59PsYf+sQwOI92h
Dn9sQQwOc1GGd5wduchPS/bbcdxiEO9EtSNp65tgwPEw/7s9Prb5NkLNyikai6Gw
9B3ySJ87Es2ui1pG6jtOwlPt0Yq78X3/t6Q1iAPyluZOX/MNWCjVMGXpjORqpHej
VQ3etQIF+xZSgPWrkEg241Boi11VtS56Am0y4Pt2i+pGMBkaQ3dEeNZFrT9pY3cD
W2ZrbxGRbxBx8LWGbp9f/1E1D/YPf9uA5CF+LTQl23pZNdSaIKlB54A+XITXObNU
c3JsgPwWQBlfWxkPbJR2xW7H3fdKatbgNJt8WqRSzzGGIFh4NC2aBAmMgn6em+/J
xAh/P/QmBowYLvsyHqDk+XcvJlB/SJkwMpEaivumoJy0B2s3t03A5r3gHy5ZUoJj
`protect END_PROTECTED
