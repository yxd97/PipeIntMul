`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3BCtVkcRweS70uXUgAfuGAMqGaie8d7J2u9mUnevdDEJwxUH905ZLKQL1rOj7Di
6WId0lvmmKlactFWHN8ucV2v6Dy/wc8Wo1MTM+VYTwmu6TpjqlJ3Ncds05elZb7y
/FZpxuRY7LsVNOcuHHNMRAtiksGfp2WREa9Vv2+ug6XiFjkaAyVC4aX4GwTFvu5s
39I1Iqw30+A+CR552ugINHDjcmu5P3LVBa6orN9cEixPfVouYkcamnmQvTnOgXCI
qVNTAkzsqAirS1Dczderb1ZNXukVv16+5pRnA01kZycEj3DLjULNm2hfYZBuQok/
XAZNC6PeO+uWXk1DRiTGbZzrcveiHkOCOJo7JUI0vJFvXgHACl7iiDu+A31A0iLD
GnOGSXF20wRsef1Qm5+MQybu7Du3YXMlUKk/u9zFPgJ2yroLeXaAaW2p5t0MFSEN
SH4ou9+tY0a/Qvr1ciiF/3/bbtejesI1UOP71ZGcOLUQk0Z7nTfePllkFSItEeSf
Os+I6f6KlVCUnKEZaCrmgLoQMmkVe2Pe+HRsAxdxAMVaVH8Rb0cZckY7gKuDXoia
H4/ktIXSsq0CiduNy6I3w9o/hMMZEdLTMh1lg0OuCEIy9fD8hbG8DESGCEFTISdD
nfvcz/yOR7q0Kq3ZE3C0e8RPIXUibtgYn0jfvvjN1u/LH2ojJ64YT9e/DjR1VXPs
G6WUC9tiGiGn+530qNNwlGIF9rLfjH4uwONE2cFknSaA8p64wBQHEDRylZVj9qnU
qasHEDxLFiYPEWEh2KIRlHSjAd4qwL7cw5kyXyzcn29jaMHNlURSBHSvQevs85zN
MdwZ/ABfAYOTNQQNP1hyRYDe6thlo8g6nOnO80/HcasNQpVj9oSIHz7AcavS/gO7
wkngq32cmVsNyadAanL4iB0DS2TP4jRKrRHyiZEc9syUw6BgTDMPQZX9PeFW9Rhz
`protect END_PROTECTED
