`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZqQtGoCkpbwpTDtzG0YaYi0A4WQWLIYE44gv3aLLXiHo3JVVxcadWuU2ihiQrpO
C8k9xffbNKH8alkkHDa6Flzz3Y8w+PjReyHxUOHAYc2C0mc1O29FoYg9H5TTTgH3
jgg2NSbN1pvbU30lAmeXbBP8ufw6jCU44pQJ4aaOQlvHiIVxpgOO2Ya9nMOgu45a
d6PgHZzdw7A5Xk4FzoikinfoqkT76/YDrGP6Q3yc+XrFnc68EOCrtk+22KUHhVUS
tPKBvwtbwTg9irxkyZWXTgF0V9jWs7KOqKnu4BQitKScm93aBApe+ReQUScFgTd/
mQDvDHP2xwjaIACH8K/9ZOAxeBLEIe2h80WigSNMBxJ7K1iUYjXQr2Iw3HIJWCX9
K8cl3aotBQuwSv+az2q+nv/vtkLvt3+uPIith7vAf/BT7jdGS9XMeZ2zB1deN/4e
jtli6ueGSgIKsR8D6+wkvrq24PExfRJohPEH0fg0thQ0z9H4FoJrJxowKVUJ8fFn
`protect END_PROTECTED
