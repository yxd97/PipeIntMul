`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYbxtQnD3AR39zKal93jrkvOgKmwibJmagF95m0KoIdG2bvS/mYRaVKvsm3LhF0v
ArZElihia+CxWUKLjyoI43pA/BdOvVCa6CHgykF6V7JsLSAVnyrwLq8K3PKzcmxi
ljGIGYRX9b7FsL4nmjbGtu73+u1zN5Apg2mhJxQUf21Iu8LHhoAW8+u947poYPhi
D6Zn0uaDzJitT2Pnqd80m9XkrIrqMELNen5Lrn0rn2ZfXiQosZrBgWuI7q71sKoA
J4KCfR+bdt2vr1x/3uLn2so2vS7gYkueSzRwNIvX6U/ZHJKqgdOAAGURMqKZM+fq
cDkzA7Tn82/WjSeGH4z7qmkD9PwBCBGZUolNxF4IKaZ17ClO/fPSngW9Zzr/8ryU
Ck6faFvAGRnfABn+c3H5767G+oK5QRh6lZ5P7QT21KSo1gmsEeR3ERVMPKym5emO
Mj1oLGQTGINVDIc0mxO5Cjru2zPrix1RqeYnOWQiGNWUbdlQ5grjci8kJf1+FfKA
w7IepMg9qYgRPCdNtscuIwAICFBb1G6FTdKfffNe+cHSs2PUy/3oGobdTME/tYoI
HSwcTW4uy9Kz7fcEaUFTtmHiNfptc16b4FJxrmzKZghGTAP2VvUZVcAEesCDQSUV
JOow2btj1umBc3Pvu1DuUhUbN5KsDv796tY5Jx30EOyiZZN5MBDpINaZ30dMijat
Ta01VNfiTehu1ObrDmKGq2DGHVAzYZPtxAu6RvKejH7Iu4+e/JS1GtXPscNn1WgP
EMwCskHbXxWXH1fO2q5hJL9CuD0vs3Kngb1mxN2677tkZUeJqbLfg069HAY8LAqk
+++I/MV9RZ8+yDNjpGX2nPmmsBpAf3+8HOAkUGcsSDGhaVX9QAna/W0HbvPnzoCs
MCbXM3P1DBX8V6m+EnTZEI5WeYIgo1lH8GEW0zlWFEAamxPK1cWzzsiyaDKdzgMd
cX6biE4CVZTKGl0jbuMEo4ode6sxfDnBGdzyGNmxKRBqRTy18lRkQEJS3aXCkv9h
0X8IYRd7JEs7G+yxNwPhdRXp8yjA5+cP8h6IRaJzUheonPjRxptx5qfimu+wxyF4
EjtTWgqrWkEdW/24x+GmrgcFfdRypDu5yn9YfkiPL0ER+b99GhD0qivc+QsYnzi4
7kSFmL0zYwo924CAP9EPgKG7735kasgevLL411kbMxwgCHv17zPudel15via3IH/
Z6PhT+hyepjk+doOhRTHUX+WLYeCR44sVQVhbDlZsK8drlS/Mi8Ol436y8UNHOIn
l/YWirfa4ngqWWEb4YtEOi+mAK/YAKNZbbFMu1PAjliKsD24Ks0B2MadHxDtA94r
FpUg0TeY1aPc0xd3M4OCYTP2fCe3JlVhkdW7BEuEslRAiXgOVMzRBDU5PWwRCDR5
vM9hUpj5bDBIA8BtRoF4uUF0vES6CpqRjaNbPDsZ9d+dCQlLExWBmInxXk1eB/pB
OsrFvJaBzu+3kE7nw9UyTT22v/EMvnYF+5p29D3nrMKFHXTk4Mb+i5uVDcOZFmVP
gTvularT8D5JClgIrQucUtNflum8C3OIoK4Y8fsF8dquiDl5vYHYsXYXc4PErZ56
z23QFhCYwMLumO2tKr24BmdVNzzQ6so4jbRURYoK1rZwWntCMUiR5LAhz4tv9qhQ
plkDmYn12RMlW+6WM4kfarFZr/16rYm8V3D3HztpTv+MtS8ac9viurhirVH8qce3
ppUwdKMzNjsAdU4iJ7ihn1gIhLyrvZpPaHl+yvP6LcSrKl2w741U8gRnOf7YpCxW
VKQOoHZPoarM9ygIfNYE03knNWBHb20OLSM+sd8a7LSAA9HEbzUynQdc/C5COMDh
roDY5rhCBxgb1SH1dYKcCOglSd4tn6GnUpNvrCgRf+BIqouBKYKwvnTVrsjYxs12
1k9fKk1HeRgaXnfbjIL4fPvxFliMRuNdGyPT7pn5NIWavCDvc/bTU79CkfORvudE
tWlIWi1VfOb45XmcLG+2FcgeSf1mIfxjqkJWBsQyA3jJFe6tvEY94Qwv0rHjOLxK
8UeVvFQVU8BKCbdkWwzHlo9JGkk01CJAfvt9fdT1koQn9UOA6gH+iR10bQKV+1BG
kQqCFKeRCU6YtAI0CCiBZuYwfTzuXr0rVnOzjD8sub1y77bZya2cYNhsljLONqwO
EvXusVcByb3nw5eCtMMsFeCNW16zNf/7EHadwRu+LXEGzoOKUJxDgLrCWWSG1RAh
gbtqHYUOjrbAmfr0woY+AymC72LGT5J6qCS1+5j2GPzRABK47+sZgFcHu8J6IFvw
uS41AusReVlOxKRDDFAGwSk+XB12Xdje0KuuCZV883guuVnc2+thuV8HZ859EpZv
rLQ+bFooVuQ5OhzvF+bg/qlyb0nw8pFKyHAjvqmCjLSFS6E7AgFqzwtZ/m4QIL/z
RoyMh+UVtNDpUU8P5nRuSYqH91kn/gcMJ2130Zv+7X+36vdGmBFA2fSa0Pkcald+
16ku4kHEYaqJme7vucccjnDxqE9KsxBeALpuMK8Ksop0YnAOV+Z6X9ggGGmwJ6eU
exjB1Qu+TmFPut0cpg6QUO5TyxNMXHz9SzD7Aq5HEfSj6rVAM/bYt4wVuj6aUWwx
Gt2Ko48kbPqNnYUWp8yjvc1aavytQ6972rzjBvs4/F0ML9emqv9xKNNjAcy7dR0J
GlD4d7lD+W5b9PkVzlzWyBkfSVd5uXqUvlwjG+gBV5dzKIJmVlEwsg1+YgC4dXER
//doCmYt/vyhJ40His5qpWCK7E7kkUpcFII0T/sKr43qY6YdDmlG124i/D+IJCoc
RbQDyLjAhwFzE5ybiiyNyl5RBgGm40GprLzbWGLs8piG/MOtx7lXUm+HjnzyTHVx
yzpUSXQAsLAxjQJIDOLNxkQ1EpOsCDOyLD/H+xKS+dC3ncxxGMY/QFAI4le+/5FO
xp8wCU0MB5m5t4g9QouDOJptNREI7O5u1DyQh5/BBt5oUrqqjeZaalGHNcDAWSla
z2MHwlW5f5WMTQUJUVzDturXYmoB43iqe8idvlJatFLt0+7MNvqlXYemwbmZlFPr
/SWvUIz5uOOSSxEPT45MhOEaBoIF5o1A3YkGexo3HnZcTCpftFdO6/17lWdmKRYg
qcYTT89A9IqwfW9vuUnDmuNgwBYbNZNe0SwtHnoEqzUSdeBbDvAkpjSL40P/uhUG
HwFjYQ8hZN9FbAAgKJ4Jb1Da0m/5ZtGVrvleLOs+WW5qJ6WZ/XY23rUoTWE49wmm
4tPqVlvscmQJfDxLKkjxdnfSGPlOKCwURNjT1yQcj9EjxBMf1cfhOZGnxi67gyNW
GEFb0QY6Nwp6GzguIE88br7g32E/NtNbxMygGiQgNZs/mP1dgo8Y9eC9xY+Ao67b
2UUdOomE1s48b2A4AfJneAQWoDoDdtKo43UQPGN19I+Bl+6uj9Qn0H6iB6d0cNRp
N8S/QU5isaee3voNcKKDq0hjHOulS7bJ1IZfWjsyT7t9bcDcz8GKIfOYnS55Gr8o
r9p1eeWLv71nx/e9pNmteP+XaN2bQZOEcFdPr15yoFQJqbAnP3U8FjEJZmuDajlf
YgRcYfKY8ggzi3SaQKgYVSv2qHHOHpmuLKCq8ye7lRUoCdr00INSb7l/Fyva/aEN
Ibijze8AplT6/jPKvrWgFjvb5D1R4wsHTiL9ECQq2/aBIO9ZCH6zCnuFJrHB2Fsb
c9YpwinOqzEW2h6AITnCY9KwMi4OiC2c+QSqpWukhz/JGc4W9o+LB2m0GXOPSr2r
`protect END_PROTECTED
