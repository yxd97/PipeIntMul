`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hgswgpdMbRXU8ScbPMSBk2pYM+sBz9qrKzGgHYrBcKAtpzVKJeiJrr203Acfo5fV
9UbhnVO6T+NR6dHCAZPNQt+oGPR17QaES8AG63ogxahSExtDUYch9qBg9AMBa19n
Hx52EFjOVpnJfoqQi+eSTlOupos8GSJIa0ctEUKhYc3uZTPVRf8I64YPCDl93/7T
Q17RCZkELBBXsa+iLP88qSr8DqyfFPziZe1w9fzgjlwX4PbEE+m159lsJL8XIk0A
T3JtgNaTMGOC/MQRr+Pn3lZRgp98KKP0wfdSAbZ+q2qTKkRnz8Cw0VOIJiSuTMmt
`protect END_PROTECTED
