`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZm3rqqT7YX8YI4ylrotqsb0/V6u/9ll8ClZQ29hxhI00jlDVj6XBvTQkTurZ3LD
nNpLSNWx0cynmHaJYvi0Sal8bbsu930fCwGRsJR7KzKA7nrYm4A50ZCbJpBDBC8Z
tmeku5ur00R0xbVXuzm0yQMiqh0TGkv7OXRZFbgYVUEDVWqXVB+ToKzU1n1WtCpv
LSQJBvIZsR5gHdNVNmDeJCqHZKnCPdANFEJ8Z9+4I8DnUDmh79AgzTit0sQS2cVv
jlw7DZ1vJ6U74yXug0EQwWKyjleuzUpstQdPN1ERbpbUFNNEjSa+nBb22gIgq+J7
rExC0RmWEDFnBbG1bD8xAswBiTtwnAaf7jTXEolSCJaXkaRpmMSX+Nfbs2SCUg5Q
RaOppUrRNS51Aidyig0Xev6e+vZZ8D6d+VrBHHh+Qb/UyV999oDG3t09BoP7BmHY
`protect END_PROTECTED
