`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yK4KVr6P1X67p2bIbRC6hohKrsyD09/D62rs35TBS8EYtSv6c58EBqyOhUB+aMrb
nJEPyCCQGCJFcafNjdSDBRnCRaJF2MDq+37CEkuDpYXYKWqnZA5XaThZDdqfbhXL
0HQFWnvy5f6bSt90MBvoaYpmEEB6Hsb10mjdJMy3paXSW0Ht9HHNXAjjFNypkbj8
GKHzPp0G2l/2ekyWY16aMDClEVtcSWqP3gigWDkyOrcrASxw4qNd9+v0F4GcqQ1S
xceAA2FBvEe30aID/7nrsxVR9gar0yWAMwFi7pEpWjo=
`protect END_PROTECTED
