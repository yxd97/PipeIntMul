`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l8veAfgoOnT6vdZnUvQFRuLzT5IPkZg7T9sX2yUayopuwEnPR5avkkTn399to6Ce
AXlZ8avwHe3rqXhX3Qd9f4MYUHt44V/A46znFVJ0gntWaxaABsFH7r0jwCgENxdQ
Hy6C6SDywwsWGlyTmL4K8bdrL+gamV0Ce9AiXY+YsCu3pRMVzYwuv/zLR8N51do7
m45/89Qvh+fwtsuuIl5y/LxBRvPhExzTBwm08BdjZWzl2mmj6s/i0cTviXsyJOk8
TymY3XWB4tGdBFlJvHblW34R5y3cIXbrQrcg3dslOBiEa7y8PzUsm/UtkoGV2vqr
1KpiralqRCRy0A/PUZLYi6tKaqDSLZyZj7hzWKtRWraYpC0Lm5ZUYzil2cUvcqcL
z+8fjoNLDQTZzkeoFbfWW1rf0A2fmbEHP3zLwn7CwTYHXjx1vc0alNJgUFexomOy
0xR1qJO/btqDm5qSRt98uvJn/IoTDURjScinwHOFMl5QIjmnhHZWK+Jm7wYPJDT9
fIPWPAo3l2VoIyD+tlRTR+tXiG+NEIZ0g4Gh/VgUWPk+UrNJsKOONwKySyM73jBP
7DZXnmtxGwf+BCwg95U/ocijIeWOl/5fvIFtfHbWoXztmD6W1mrt0zaAk/v8VC+k
DHWA8sz1zAHlvVHlY6evJVr+AzW7Tp3H1hxoqkssjUl67EsgYURYubO/zE5hcat8
92F79EMr+qifBR4DfQQB1CQ1d2e2488Aj+pa1gN5NquUhV1BRsbDR3NBBzl98qq0
Uybli+QAQTjVRoWEnH7Zh/+/PrltGb1PzxsGK0QjjcD9r2lA6BswLWrVY48S3B8G
MODHyHo+ZvNEdNtYe3QxztVA4El90yxfBaVaEO+lKLdO1CagH9M7z3c07RDs58j4
JkZ7H0a+Be7OHPltOpJdmPS6xQSuU1K165kA39ZDiLNmCk1nSTLfdm+UvwRONKO1
gzSztIoMubwOBzE4j+6KRMJyxkglRPxvADRvF4NmlwFU1zWDzy/4sR+LXI52Ce8v
PWWccTJ2TJ/YsyAHe6Nn4N1SEpShXnOAOGKd/K1XRu/Iq9zo1nOoJdefuiSOpBe5
U5JN02JyXxkNn8BEEJV9jokUVcmQ6wrwNw2Nh3VSz1rC0AtSAGzZACNFyt1dep+2
i5vywzGJ5toR1mU2HkKPj6+dkgO2fwThADcEfxpKtiNwABFrVz1M36t07z85/mkO
dUh2ektLFRzRiqcMFHutKbeKjljhQgnU6sUgfEEcdoBYPk/ccCk1+2P9ufg9H2FK
D1eC8Y7WheX61nzjJ9nxpU12rk+MF2aoeKEZlBpTeNmtV90VwgHDz9Ixyify29hm
Yd4yj43MOwcaDWA8OLO3Hgmid5UwCo4ghaQvqYyDaIaavWu6+jtaavTjOSjjMe81
LKiTQC5grIvP3DAQ+N1tp7M6YGuBXLCm96IL5CaFKjfaF1tVsIyDFkPHqVvOxL5S
LeHBwCFpjFU63Yx0wtItdJqqp41pjhdOyoFoP/HL7VO9sAtD0Krw5iK6YrPRclo9
bUBdH45JM5jdFVFqrnf5vSxCUZGnwbcW1/UtEcFfx1QTOjCu0g2m8Z9a4hWtZ65G
MXOcg3RcOQ8WBFiQE/W/6H+zxbZmCdjBFCHSIZ5LPn3B4A4311EVKJBiNC/aWj28
lYw+aQ8ph/N8pRSOm7SNToM913/APTsnbLEEHTHDCRBdE/hTpVDzUzazd+f9qDSU
IjfSdvyMzh53KNey04M+74ubqvGDWI8AHoAXpIHYLZ+I9KHZOKQ/vN7Jxg11j8Xz
6wl/mnnn8nxXS/BkFEpQz9FrFXYIe+1HS0PyI6KVkdHFTPMSL6Qd/AvIiGryLB56
VtGuJYH0qTTHIDY1uPFVlkUe3eo+cK/CdafafPFBf8sRauDmP9ypr9/lmBfJbJV8
/HBgw42d3gFye1VfBriviT7oyWqCOPcVtrAneGTKn0qeJeDmXXKuRvgKKmud6woA
6xx/ZcUJAtH9hGU8UUWwavClSchtQcA+r7ZcCxhiBAmvmZ8MUCI9OfCoS2+U6JCa
yOIp2YWsdKJu0SKLaf9AYd+TaijYD/GC8196oPU1dnazWRlIY94ILPpZgm09WBJc
b88PmZ9CfQ/mY1eRq4C8/rfnBBj2Mao3XTUApfUdXtNIyIvwBf8bSQNt63eXuoFz
qG4fgAgxfmLW8K2diUYtQ47+lFrifHmGWzxyhJTEzesDCFnAt/wftbDedES6e9Oq
HRFhulEOeFtlojkdfBSHp1VmaHi0H7cQm7ZkYg1bjVBGhUA3OI7DZMsx3IUN9/2q
X4PA1uPwaX4/6bwK6hv7Lc9WDf/3S8TWnJds8X7x+KLR1WOf0C5k+XRuJTzGU8RF
LHa+HH37OnvGsySmKAZpde2A1hFPa1Es7WuHnAkZ17Y7dNWCnQQNtEGaJm742kja
2Jr1MzO03HYqVndjTlkgWMXij116vX7TMEkLz8FMnfs3xW08SLG4BSns7WIEv27k
`protect END_PROTECTED
