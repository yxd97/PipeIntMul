`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fpOBnWGomUfvbYmJazZxB0scwjt3w7d+rutZ57W/aC5NTU7bb3vPWhHdI6VPqPNv
VW4LW9B5UyXfr6uSBvDND58SGr2JJFEwtGQxvFEwdw9e260D9I5GuwNh76wLWQ4K
hlrj9cGA8zjoqR2GswH47SqPaLzoDGXUfAH7jVWx0HOSTCicX69F/LYCOktDqtdA
MC01KgL+ChETdkX5jwfqq+aDIby42kMOe07n490NeX33N3VNw7IO1ZUyjPsKq3E/
NslU11xgthD3+v/q3UIw8Nk3H5IL39Q3QDnHjwzoNpsrwH01ndLt/DpFaokVOsZi
t0cXPnbVdn+hfM3LEHAxHp+7o0xbq6KJa5dIo1qg5SdweyBRcUIlH5eMC8CgVW2R
o66fjHKP3kaff1V6NfWmV+ag0t/c2/18g2aEYvyTp3Xtu6WjoIua9PpywJWt2c/u
zb9G9mKxcREZtGVg0WgYBuqC5Q2cUiJthCZ67RcNGW7zcG/ObKG4+2/iiEQ8+b8q
4Q3iYphfY/IvbmOIVkf3GR4qMoaTq2oOOvp4VoqWKRcJii423t0cTDkXZuI493nT
leqn4XHN24p1lOZN5o78ErmA3zIqNpRv/bZ8dsqOgUD271SBmaP6CV4qLzKmYUQs
wvrfIK7OtQ1m+KNIID6BV4LDXIfe5pEIMRHMxaViBwKYTYoYcWj9rmNFyQ1UR6HY
yXUd4GCvh/g2d2eBWyG5rHSZCuOc6qOffNqMdUDUkiiu4UgMHBt9QU6AonA8epwF
KqGXjEhYEW9JnmqGPM5QV7wlTXGaoPPTcS8DNzq9i3aeFxZlZ/OhyaB6E8P3eInY
vRX0mTfGOftfKbz6zdrvIum7tnoUmk3z1jyO7UHslfNrFFCLvuhtNgs4E6p/pmM8
t1q4ZTRenSiDyBMhqr57HzhPlCzWh5TA3UXVUJz/HgpLSqHKYgryBg0ocXIDY6zd
IXcu5cRCodvRO/ximC3TN9V/7CRq7LAFUsOXB/jJFE9C2fcXbA93CWbMCZPa9O7P
9Iy+FmAJYly75r0J5bEdmgWOlmQNRLP2aoG7imqHDTrFiV/9EIpJrLmjc7hejnAw
xnuMfFBKemb3dqvyrcO1FoIQBwD5wieW0eLQ5UjEY5JouXL7QQvuW41N6WU0j0OF
/MW8aCH7xzwdziIR+hAuvlTtw3gB8mP01xT5upEVx27sS9mHZw9JxVUMHHY8smjn
Q/IFI3GoQnZBw5vyX9lfqERVA5MpVrQd3a/zuwp8tWp45Ma2TduqbTrJnIT1KPw4
9o8ibqd4VCipxCFOPxOEaINBY0nfhD0ffav3DCcNIqMTOkfpIRJQCWwG2F7dDlDQ
QDTDNEzN8G0F7lwyKC/podFST6Xf1T18kg2kYNQnnZB0eysPm4lDsa8GHfweBpOf
B0OqLtx+gi7Aa0NpoMvxmNFDdrZiSJ2q+vvfbS5PoFU/NnGjek4H6oP3rAFEttRq
1O8fjm/OacRgFKG2c4C3fj98Y5sLSwyYVhgMMDIgs+xIZEEkwgWbeAiidrQxCqi1
iRyilBo+srhYS0AZWD22QFTLqb4HcQLTLIbcokpVctvV8orGamkDglXwnsamfurj
/yje00nGTATLp9hnX6oUZX46tEOF9CL7xBYWhPfNnRAYitgx1Fn+EOHPmapiVRf4
9LRzRInPwLcpMqevmMh+Nl3tCEs88W/p8hRRd2Q57FKfG/gatMDTCMoHYGT5nSLM
37TubAyxCXHnSty16c9LHkFR9ZVLC6JgIHNj9ieUQ/3APiBGKwOSxt13nvMtEHzA
pezOKC+yQZqkqNPKWw3dEumFUoeqLWm01DzXq8GkDp1PFNdy/khP/fggnreFYO5r
wqf+Hpgy6H35ouOOu1wEDxL53hidMPl+q8E5s6F6KzDZgUvYB+XjSBi78ZW/gtqO
VgIrBGgxYpBzV5QPoL2ofR1c/79DO0SdBobAchKAVUEEeOjQz2faVHcr2XBYJayt
wY30fqsJzdM1YNTrv54hJin3rpLFc73SWRrSqvae4P0+J10m29bTSZObmiGX/9IF
+Hrm/NbXP08G2dt7tf4TiyLtsXsHNZLAObWSESwFIxJ/xqoyiBhoWZUkE+2lI3Oy
GoL7INprmhLUj+jUzfOCswq5REGN/r2PeQ2UMupg1JlVI0tP7H5T4C/EKA+xrNn6
NPeqHZPKfoqDiiJYQMFRqZFgrXWJh38/LQuwXsSzI+RurJ6ihbDu0p39ZjW2i65a
TnxQ9OZSdSp6hDKgavwf9moKb9KU69le4iK0QUFR0gU3OMwG4p+DcrEh4X8vh96D
zIc/wnzMBaiYXpQ5jVlTZPL+kweQa8GLbWdEGca8T2pqGzCyjj23aCxY925+O7+A
ZqeLgG4Whq9bbBoFy6W/xKBqWej0Oij0jF53cw7JE1hRO5suqD2l5TBlyiqYiGc9
kvayUcqA7mTzwjSiseHbp45LdF8yFO4RCdegQFA2vEEs+G5IqKy5UNLAkL4qnsV7
fu3cDDkD99PyV5Vbx960sfBX3i7TBbez4aY1WsfL44y4OogOR3bEOr7A7Zc7+xtb
fs4m0021aJNJskgNxrSXQ3B9Z5a7Y4Nh/1MvOGRhXyH8oRZs3+/U5jyl1IOpvACW
I5jLtsEE5uZcwt7O2a991Cvx+SD2w9Zw79KrtuNWdCX6cEc3KyAGTnpFEd39IXc3
PxpPXiJl7pyR7OEiDmpB7gfjO+j//v40qxBbG4ErPWpDZfbGh7xHyc7Z5raq3jON
aV4q7B2zy+PQVOn8XrwzPvo9xz5sNizCtVeciNcSNBjh9yKWymmKXqzwYbWSihrR
DyDPsEe+xFmUo8QsnqWHdUwuG+fWB6Ti5FM0bfgEc4wYErucvL8UprDHg7QipyOu
qy4Gsbj/tSKCB32rHCGLlgk6/QIRowDi6yHCecrST0eOsxtC3XowOUc23uHJK7MV
wd4TRfGb6nTA9YcPyA2tglIgK3ncMSJrQxkgAWOCFO/qTUQEq8Hav3Dm1DJIAzjp
fijLGyBrDGKtUPwosLkfG7dw3qPzxUgk/Ra+ny2oPlbsxEr7Gw0GO5LKbqCz7az4
gLrqq0Xcl4QwIkBn3+EjnFQIKRSIXni7IZ/zs3jtnIFdlAnxpGM9b0RPUsqcxpNs
8kbaZtDiF/oeU0m0q1RdPGEbTop+jTMkF7u6l9aWax5XLSxmYrSRyGko8VNHw93z
ZgchjdKS87fTJEGRFonXqZPI3uMiOQUMF65gA03OQMRxeGmaP79mCNJEojOIrXBd
iitm87bs23s5iYiNeh5QLbq2In+VgiaBuu05ERHjKHiTZIRreAjLeE218xAWQBye
936bdmI9CDFzt/SOwyrPasd/4utkzmOa2h024x3B2pjdYUVxzgmt1DF47tLgFMyq
bL0j6UrlSGgCKXaJxhjJdqmkvHFuTs8a9R5xFz5Iv/53b80snCUbgeRKBOIS8NNX
Qom3pUb/7Ap2pc6JwJggILuexwjTJM5EaxkiI+QShsgN1d3UI46hIXgevb+VSfGb
rA6rumKXY9ry2LGbNdrpmJ2tdZ0fH0ZHDoBq3VAtwBQtfyYtBGLEVKDPMzOpWaMv
P4B8LpGm85Y8bmFedaBsiWPVnAOVIvV9/WiPpWP3p3tkOYni7kYQOUsdgRr0icGU
gUmo6lw/Bvk4QLEbZpNWN3YgoYIjMNMn+9hm4ajadfTswz88uQcpfT1iobpt43n6
PpxVH0RAujT4GEChkWEHff+DOSqJTQBJ0JJuLOJKO5a5Bk+kXujM79Q27bKZ72Pt
/x78x4LsVbL9W4HtAw/EdjJ8x8fg/2lqN5TbzzUq/G4ztptwSTEgL1IRg8Z5Luxf
21Xfa+ZbIbZQkSBxQevfwSIyBAbj3EWcEaOfo21h0CQdh+R+7YA3r/Ihk3AlBr0n
tZB/TH9pDMGdEWJAhhwYJDIIlqU2m6Tb+Bog9077AkoYbMkflvGI0cCtiW1oKU0O
memE7bfnhpaLoC3LIPhMTRlWvGm1VanEksO7qZvxZPxSPVRLhv+VqJtEH+f8ppD2
zo7nENFw1X+tD8gM/HgbYn5oM2DW/D7q/NKDPXi6uk0qr5Pn7J4h1Hu9SXWXPTSE
15AQWOEOqa+B/6FoV7/4syjG7JAq+rlzcE2cqeTJg497FO9SkFHm8qnhyZYswl3p
nYdIe3Q5OLQ8agcGoQD8FTya+6fd/bcsWpH+f3NmvkdA7ZtsrGbTNPtT9SS0S0dr
25GDK4B53F+h3PAKkZqO+JaJNbbToFisdOF+RS3pAgMZjyy8VCe6n5KRMJIhctAL
m8bLoc6H79KJeVNeTT09l9ctQs78rXUZ88YOy+sjarzbhe+Ws9FbHswaVuh6Yh8k
JEBwRYCV3SXrVkwA06ueRwfucCp06wdG+JbnnkOsocRnUk4ngqsLcaNs2RRk6tFV
xAQH4TYOBTJdJALw8Zf/a1+TTFzJlO5BCTBc1lhZSWmmewZJNraRJfVXkcuuZpf3
P8QfbZSu9ITqmFBCe7GfnfgChAo2vPSoPkZjkRd6wwKlN9tkrmfv/q9bGYw2zfqQ
ZqRp505K8lV6QltjD2p3BQn9nDLSe7f8kIn8EvGGlr61jVJiJxNwy7zlde76Rw7E
6RMSNjNQ+JgVzz2Zyd5AckAavPbQW6xhzhYpFgoG9Q6mM6TTM8iDeYDQpPRkAiZi
pcAZ66N+LP6n3t4EtCzNrgmuA7qx9wVp3UvyfvqfC26agUaa9ZAq/Q1Wq7ROHiDa
mIxDL2sSGJFSvT3VXK8Bm559DsC2HPGFPxD3bdKPS8O+2RoGWIeGXi2fkVnpGaoN
Hbalc7OL12zQv/U0qzP7/Qq8Cm3Uo497J1OnedAhWuH9AbGvroz8lRtyWGqAfyYr
UVV/OfPXDaEVqOVoM74EM0i6zkeJNR0IR/nDalK3lzVLW049pueT0VE8Hy7fSxkx
mLhL5vTXUWy3qQIxuT1T+z0FkzA2y+SRdC9Q8d0IyxpE1jvmwtu/kzmZEqnWJYv0
q3IlVK6pfiM4jiIWhuJeaTStXWoCxxtYYaStztq+LCtSiQoQH5TLgwOGjwWmPnGU
uCW6iaviyIrirUstXNzaypQlKtKkNnas0bgl6w+AzwHZ7HhBjSM8ftoWx7/HLq1W
rQv5FKvLr98yEACFFc43CPnsqhM3JHuk98U8fGKoOgA/GJSL6RSUGoVeSTcWssBK
d2eebwYQ26zLv+vDSgHq8xf7x8yrsv/Lq7EwMfas8V9jm5BTLNWPeK4XdffmvYyF
r/e+LCNTy5/EBjKyda5/aBsUn0iv39Whgt6uIQvsJGQrs+pQD69Fsqei5W+kx6Oy
ZhOsliMWWDgNb/YjDgZj2nd8kAiORPfltVMx3GIY381pkxBh4IgDOhfUnj8Mtd9N
KM2E+rsRIDgBIWbz0HulhNxhvhoMEHpADU6z27A13tkGIRTKxZ6Uj2HZPJoHi+mH
twhKxC8TX5rz2kqAtGxzPmcDEViq2DI7OSSypjDicpQs5eUQM1ZwVNm2wtisvMmd
KvlaGmA5k1rT+hrzUf4/+v6DWn+Oz7aK1Fm2h/Mtjk7OOj2wZx3OVMlc6eabR3Ny
ZKp7DtJ4vonHAY8FoXOuvrvfApVKLfgON+lmPKpRBHlA5auW8RpYmZEMQ6P3WJ6t
jOiNjpApB/AOhHRATHvR087IPTPLWZhgFSU9wwpVqZrpXCXqDWfS5ptYpmabo+Ev
uML2STLs7pnkffUuc6kcsJFvoefuUG7jeiMvYOKQakTNNdhSwmMINFKiu86SP9YF
qMBYyrMhP9tZVOp8cqWqt1Zy/r6p8aSQTfsb0bIcJCXuWor2m0EUj666+w6q98pE
RRGvxstqHQI1o+fCmN7Q6M7sMtW73xYGMDkRQ/+RBv7rBeMK/Db2+quxTn4AeU+r
gZP/Tm0kEoG7+G1wHQItjUpE7YrMPQQP+18TSkpgnBkSBdzyxnQm9TV/aBwE6W0c
uVz5SR3lOh00Fr5YxoXNxQ7zyLCM59mIpLIV/YzMGZQNOehxKdq85nJuckoMuMnd
v/BucjTME31PJUYCwd49HL+ShkMK3QpntVraRPoe4diVPj0u/WXgw3TCWrOJnjZz
Kya8Fb3COKmlCY8K89plTY1bsOVV5zT67UKXX51daN1iveK8+FSj4Ezs7iXAdybj
S5RjOFH4RryIFsM2rERqs+3+FG3imCG1B6LZDuiSo/JQSDxDfn8Dz8VeLBQ5uiE4
PzlKGEefuexHfXFM/PHt7ANK97SFH06daq+2bBXT22sQ5WAVqO4u98Cc4uxS/3si
qx4y++ynM/6MHAiACaQuNQ6FavFCHf0Rjpkr9HC9IrW4G29f10XGhXvcVvN4Gp6n
hhvQya4pZS4Z8nV29woExoxUd+kWBPgHg2KSJH0h3qyxXILmeI9dnxVtmEP2yE1B
XKCSHz4UoVUl8dJsqhoSHI0Qqjs2QcbJzfR932+IWZfP+QXbWp6wUoLTUw5JvGij
e94Cs+EAaYVVy2IE/TEredG0IprEZjesrLlAKMwLlElJwRT2M4lEP7rHlIq7PTaD
LSENcORG13qmKCwFufpeXdrwFDYhIBtzwcKOpAEz4s++GEj2rDgjc4o9ossNSUN5
MadSFCNQQkrRNEGpurAH8td4yYZodupO1LYt1dmWUiRJPew2l7q1B01Mg3gXo1Xr
uk49P96RYIrk579C/Q6mIqOLFijQ1urLSCZn+YwvhaUa4CIRrgWmQ96DZl/WSO/G
pSc1TYjz5J6cIDlMgCnrbmMC2kk0szIGrwBzIW5tlgZlwtAzPoxLJ+6kivmi1thT
f5DPGD6uxS+JjT4W8v5XgnV40AcalP5N5/oWmliZGepNVXDSkVwztRjPCNVd0NF/
LxbjARnkpAUq09/V0LCnYB01sx6kNY568hzHQuZnl3h5HEcr7e/wlWVHhyNFkw6t
iCDzfMQVWVnOSEfCHhliv7w0jGiSX+Pg3R/scKdOkYX/YX8m58SGs27Oo/xYeENf
3rsWftkxPNfLH+3UTgOoJ9nwrDXiWmBFqKnb67jna/kf2XjnDOC/Do4jR6dVNoPw
pgdxU4fBZKX5feMLR8vYrqSxbShtxTSdjddV/mPovkUXV2wifUPEv/S6v/j0T6PL
ml1a+YXNQe5tk1G8k86gD31n6U5Mt4ZiDHQFwtcqz6/+YJ3ZXNCA7YSLatq2zSUx
F5PQBiHM2hiutIx0/zqwnmQOcUP7pBGj+4j9uqP7neM90Prxw86uc1Sk7VlTV8GT
/a+DAJetYjsD1hthM8r6oOjp2Qu8JI+lRNIAk7h79LDElgt/K9CTatzfxJl3yIZ5
x4/KaI3TtJK2Si6W01Br+LpSfZS5of1isdNYvD5CqAO83Ti44H720FdlxYVFQeBj
KABPo++zrbaPbzbKKwKioLxEFaP5OPJuj3kf3mxao66qkR16xeIzQ57V8HooMSqT
5Z04zQoVPe4dOCKs0hGEAZk9o9t4X6ZW411/s1p8OG2iO9RSSDu2Oan7sZ3MqWNb
Zfo7Ym4Ef18w2XU/AxonDfF8Nql6koozcHnddupg4TP1XBm1Puv5dmSrcZr5nz9I
Y3iTimGrFQsBWWJD97sDzXec7z/V533RQbjXRmcVVz2OO1CUs53CXsDtQVSseSuM
Bri1tfrmURAslANUE4FAtYScJAWvMmZG5s5mr/LlIpkU5rrFUY7K+Nx6KYnSLccf
z2kmM3AjuQZ91rkZpVCSWjn+1h7bpMSHB3drJdwm5OYUliefKCTOS2kPjIc3/pwq
KMBYeXTowyWnXJ2F5cPm1g==
`protect END_PROTECTED
