`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7bCyDrGd6ySJJozB6KJUX32MqhSL7fsNrWwA4U2Tt09ZmV8Urwd3jGp3Q+oTFJj
Ikpuu4gAr77LTRTmk7ZkvJM7aebPUHxc/9hkVDo7F1SIdqCOhJD5A8iiaTsxCYId
lm2xeqzAd/MsipUFZYF9eaXT/LinxRlfGLw5WyyDrVuJQEX8CRVf5614V2v3jBoy
rDR6+l3C7vaomItsMrhRHOOgwzQpneatmfd3USWE7e4dGNoKLefxbg7K21w+QHKa
KE3X8qpUuh3E3L+Cn0V01CA0ratK1mEvw1eSPfyjB6CbCNT80L6aEUGI4MGUktq9
VHoEbSu6L+utS/CCPgqNQaZo8XU0x7gwiM5DiQvGZkQPwgfiGO482gZBcXfXHHee
jYmmT+aIg2UoQqcH1P2DpgtDO4wkB5vk2cCintskoBlCBzAYM2SBaR2OtwuY5oWX
JLEaKp7wsSuPQBwo5FRhjkacNqhEZ6VaCG+yRt31VCkCq0TPQBa3gy6SrdZqmw3r
l3Mj2k6L4akVwJQ1pRU0s6unOK9X4lxuev688oV3+RFS/H6A6+NbgZHOQ/FTL3H0
PFTEvnV3Ibes8vwM6mQxRwjN/Z8ze6EEnLjePWxNUF4/DhSOm87Tu14VmG3nzbAr
dnaH7tkt+/zXCr6CyHACRoVelzmBdG8OB2nkpgi+55UKzeY+H8nCXjr40LgW1GdI
KjHy61Z5NjKYWamBrsK4SD+0V056bd1vdONQjUR9yIf5LLSNO9OqGLWINv/vrWcU
`protect END_PROTECTED
