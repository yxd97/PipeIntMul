`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v3B4s6UTXUV95aZ2s59M/cA96zmHEfpcxZHjgx5sbsRxXOnBupWJvOPTPpMfLBal
WKUqTsMVxfpL1dxe9TZ1uq0glM3V2nHXpXpK8tLsoq2veOLrmH6BtX09odfPjMit
0jxPNQrIs6zTm17hdxHV49DxdRCsoLRSVF1aG6hQD4/Wl04sZwpiw8Z9Bbo/mpsB
HmLQJm8Ok/3csnZFKDLrf6FRa78yUaHfKtIB5O7s+uf3EJHVf1eu6xzy2jtyIPip
ugayPIK809GTTluxkfhrEgqMFdWvAzIrOpqIEGBOQIsKzqDkInAtt7cBi5DqkRe3
IzDAydtTIUozXACa1xCDKemeXR0lLjcFQW5oOw0nKEkruAsj6pIo7gmg/JacSQ2c
ytSj/+wa2cj25zDIzIYwByUGrlXSDZapcUsmd9EOz0ZAJSwFVZek+qz7Dg3dG8Nr
DSI3EID6Oo2jJpQuMZ4uqtUr4dGzgkYV0mKOPzomsChVLDUCR9Dd6GRaFdyJ6pr9
mFy1akEYBwBr4ZkdqrBDsjpPLQ5iX0/rNniFS9O/1qzKL901tv7HOj3e2WwD4IJ5
oECPWTzTOnKri1OhWMHZwcCqQqQr5RGhYW+jLfm6gGk2NBSym3SL8eWMS31eULMW
84lUo+wEWHHnop0r/0HDTMYOVACsVD11MMtAvvkpFLje7kQ2kI5E8qgnknjj1US6
axoAwm1Q43514Zqvj4QcE56Qm+NgALx7edH5I9qlncYqtLXr6AH8ImEeMkFfJo6G
IFAJuVKgPteMREUw7YQ4vNTuFi1otmYODKCtCjXSzcde9Vp1MPtuSL41D5oZqtXr
j2lbea7R21R+ZjWfjGmtcycMwvAG19rOqzRx1iB9ZjAZ5aFKhTW3PvHkC2Loxt9E
eHAHWN8m38FOGeyxE1paTUl/G+DfbwHJ7FkZDA4UZ9EjkYCwX8EVGtsYTWaUeaWE
GtKuKaplQ8zCgYUcBybwe0c+ZQJ+uWIqGwqZjegOaby2tMkozTeMZfnjdSOxMQef
if2BOL5erLOQeSvPz1QI6aV5WyNB1YjYJDCeZ7ioOmSsWiqoTHH6ES3daPn8ohHX
qilkSAomwUj+gk+KtN/EeEGagklJf/OcBYYwqfxsgybvGGDSnL9XyEc++r/gUIiC
YiHKoa1HexmiEx95URI1ytXVypCPU7+a7hqRR6kC0jxTM9neP2K3O66vKPGk0hak
9Khq6xjhocCPrwHUihK0M7a4J6/X6cOiraO9mG/7a7UimOLIyP6VUEDSEOGLq2El
AoNhLnAVFcbdwpjnm2RONA5aLOrd8lix0osf2p6byqRjWdYx+TwRyWTujocaWSCF
9cvoXqqyFecBUG3W1K/Y0DlJt26cFaMjAZPz0hvFA2H0LdiLa/idPtZVF2NYt6PS
/dPTlZ0VHu6WOytmkP1peQq5wtMsRGE4mFzCBS+12LPo6/Wam1oHorcT5WcVw9NT
PhXXU1p6NasarioSFEJTqGFPCqo4NdR5s7AkTnW1vBLW+HbHKaqsdzuT2SGsWFRD
b27YoouxwTzEO9B222A2WQ1iHbmOvfN3r5/zYdjKYWlQSg0sm0AgMtanX97a2U8g
WBIP2n1Fkw2c9Bm7oLnW/vmvakUTtDMCp5KdU0UWpm/T9iOkAD1KudhP9Iznb1Or
X+aecx5IQmwHnLGEnXqFQAq+cCcsB3PgDMC5vH3OYBovFU894H3xSekoEHlJyQV9
O/33jfl7S3DgLBiPlqVaGEyO8ETVgYy/bIHcl+NCZCaA3HPYB7hnVawNJJ7HXjPI
CGnxeBJxW02xCf3uttkvB9hEcRLR1IiApueozu9qUg3zGvMxre3Nyb79UsDLyQCE
fImXqfAqZ42oXI8I195dSR+1Q9KNmn/bvziySn600oCb8oyqoZYfXpXxtXMAd+va
XJn9v1xSR5joGwgVzI2JNd7jqdDOW82iN6KOaEqZ+jNNuENDJDEob3q1yDeDhjaz
XLBGST+hl16D+P/ZPT1+/7xgcuu34/iYHd9vM+3FojyvYbpII2k5NYaan5PAYja8
mQRi04ODE0irWKID06/EYQXe3f4UUpcys0Tuu4YBYrzpxYYUUCcK+C7Q92fthrOy
Tb0Jsa7xBGRMLrt3JDbBQREgoqeGG1kS18Jelm9eRpWSC7Ly6gxeVTAO1A1e0Vba
QGBG1WD6PKNv6/IepHEWNSTZNcFA68iYGiH1ehvigaL8b00+sXa6wEL3FD1COzZe
dSlnASjGrZMUed8HiCTUzew7Dhxsmrxh6QDfVN8lqrf9BPpsI5Nj5BPcCFpgDLfX
P59AkMTXwPpJOI3/p5wWcHv7Z0wGiBC924X/hKesC3uVv46XDAXewtjQWGjl1a2D
vU2k7AC5+JgE9spD0IkeZBrTHoxDsaBR4ytvX7Q4dgpl5BkRUWcthzJ8nevmiJnK
kB+CT4I2xjUDpNrgKxodH88Ex8B/E4PabGiWiWQ6KxYzK5VphB5nctwJnJkBV7zW
2Xj0N9dPua3HxtUJYYpcZpdAOZz34LePAfCjOOELZdKvi43kq0mKnspEcgTRV6gf
p7Tv0LuLyFz08HrCm9Rr6lRBKNOfg6LwzYsv98+5lZf1FUmwKAKEk7vThc82rXMu
2axssWjzoAnxE0yW/BgZiN1A865ri3vwcPgcgB/VMQA2pDSXfB2tG6XuBi9wsVlk
BNlBnhWqf7/8gspl5BpghUj9mSBxOPprIZ4rgDJV0R2iUjLoHxN31rVzlIC0OH07
bQPHRQjOuHOAUkFWhRY7QS0mccw/izyp/sRBj5SBjyk1dRoI9GbK/Lvp9ySz/7mg
2sCkz7V+a5SWj66PjjE9R3VkGi0BOEz+13rxLuuWQsCcDIuPkY+RZ2VX28j8MTPp
qQC+B8fI9qKir+14uzW4vKr1v7yTrGVS2dJA1L5xzTOVh653piyG8q2J+96KdwI6
VVfDaHoAIwlIchm9vjkJ5cqXyV6zG/9LCLcAVLGBOzGmN0xtfXQsq9cEoiBBNw3Q
D3AcFnO5D6UTy30M0Wfb5P4IfU0yY1fUBW6F8POaL6UQknqIPb7vbRe8I4SUP6nC
N0pRpoRxoNBOzOMkxFh2jvNbF8jjiVoyfwRz9FfxaImr20SNMA1b+00rh2QJ3v7S
Dm2VvfxyzcE/QN8Twh/VlXTJdA75Zu6ZWfuzoEHxjdr/p178EVRRkwjFTLr4Mu7x
Q7iVbMefxdds4sfxJgcMku0VNN/dp3NPXmb99CYcm0q0EU4Aj4vkLfG1KUXCqt5y
EDD68ObKn7uzLh42WEwsRw7NCNLuks2E9S7StJ2CeuFH+n/0XJhuxuYJV5PoD6Kz
kkn1zK5zNds+ujRFBEpj4En/6zARwDSZKvQPYyp/NjTmduRtIxPzX4/yJY8THaxg
XHVJxy+WzIGqhdUCMweL6fRhTrkBZTALC1Yj/5aH2fzjdsPtpYfdFTowySvpx3VB
ceJjqtyMLGLVbnodfqsZAnyJB+3MHt6oqRcGUHBQHpkXsWPOmOMrS9c1BILrJx4q
ZGzCEVH3C6BWf7OqaKTltz/E7Cio/AMUvHVgFSqutdnQhRi7HQHAH1ygoCVsyhow
AkSfc/0uFEquJZ3a5EWiQvc5k6hq3cqhOegirKClEaNpj+zhP/xo4NHIiOL5X87i
7twlFFWxfSQF5eyuBfCWkLrXwo14ZSNDoeJz7fO6i+msdKoxB1Xd1Bg4tOQzUqZ0
wP17Re78onlDgLiQ2p7Mf2mw8x2nKyoenX/vX2yk0ChIyxNNZu8TL2G8PaROUggg
l11LMgfCKtVM68mla33VD2XEpTKa6/6wVFngxhSdJUBVtBX9tQ335PO2yLc9C2/M
WEmH0urmi0G6S2OwNl78ZDEIZe3P7TNS09RcByY5/jnPX03FuQZz+XJU6Gg1KKt2
QJcnxCyPqJz00F2OBIEVMJR1C/1OskKEaGsMnifEkSQEccz2mC89p37iTUJbD4IO
WbSLC9anpIm2S+AeQPFSg+tWbEK+4uICc6fxC5ooQ2wfzgL6Xc3oONXJLM3TxBU7
82tbyMZGo+OshnNgECFw6MqEzv/Nvn2YyMDeiAI+Ft4QvzQDqjxcAGoTHAl7KFnE
eILJl8wonhjkQO+Rj5pYGWUrE+2HALaTVcM8klwsqBBx5R/JOoOGpSHiCL01RNiO
f1TfwI/23URxb2hcN3i9JGSg4uwaHjca8CGCnF9hgReGx3FnXdZpCrW94Ai7+Ihq
jn0yIaR2CB+c7nHB3YNaWzzfa/CKeRCK9JboHEhdm414Kbz3Vrd+QwRliesB85VA
`protect END_PROTECTED
