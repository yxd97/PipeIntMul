`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8L612L8qC19b5t7SsJcfDrmXV6MDyreL7Gk0P7hWvbXGvZl3CdSNJ46NuCJ8RIs/
V5v3mU6iMc30z+6KKaytBJZanQNeHtBxZTPpYg0p/rLS4hUtyNKCuI52LeyB/URd
kuRNG1yWyQRkPhADxJTPCH6zZH9V6hQJ0q7QYfKYMf0n3Zag7FfjvynQQVDATzUr
kD8/zQagKTFNNmSCh2ZII35bUWhFa1nlUAW7qrAhicO02QEL7Mcc3FZWlgH2q+rz
1AGii/VDDzcbRmh3gjV9WgQOTE8Sn4ex8sS5W+PTB68u5AEqRrKBf0EjPOR0pNdF
ghxFR4N+Seu/t5MsalPqKzmrn4B1eNXqoMR9KIr+yYaWSgQayaLhNuaMeGOkpRFJ
yO0TIle+kJT+/D6BMDYPD6T1Axl5ON6ImWJZuAtRkZ3Rao8zIY5wUTELhXC/G7ry
BXr+bszZGVRK7zhZ5Dy/FbreLRrg/TQdkwlp7svlfmQR3FGZOyJBySf5jpnmvcAm
`protect END_PROTECTED
