`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPMelFHkq0dM+BjigkeZten4Nol8P+SPJtLyJc72IWy9KfsqlSMS61WdINloRTjJ
edekOepXTWj7dO1B4b3VAmlvu5xCOmIU9ab3YJJUPQCUD5PC96F/dSb9HKzte60h
XaSZrcfq5nP+1CZrUd3OI2W9DUEN43oaXPLcgKdTIUQhNiR/QXwAety72XqW8U6z
3Z3T1J5zX9PSpU+hat4HiuNkxJcPJdt9G8EJ+AmnS9YAtOP5rO8LAA+U4eYGkawv
i7Bez1NupbyfAUHhn2fiHyWJLucv7tjzfmjWD2bmQujtPVRNnDm4EAnhy4IlA9sZ
I7GR2tvDE8AzKqioLhRjgSgWu/Z+biYkrqC8W1Uvy7WfzIMB+0/bgfN7GXDEUiaQ
7PIYmKw7pye2N9eI4oodVJVTWPdTKJjnz6IHzHadM/OTuKZjbEOKNkteU66VFVBb
I1wNrGrNM5qQTi0W1SFNPouus/8WhlvLdHgQ59p09oveOrKOdpEoRJtcGhEpPuSy
`protect END_PROTECTED
