`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuaGamqXGnpdbmrb7lNGMMVxxd5qtrTCoxR+su0eag6O32HWwStE+wGq+j0z3D/o
2sxkGlKZDZx+/12JgacUW0rm+ITbqwNp2lb3nZbTKVpQXNUoyrkztvGCWVLiOJQ5
lm8mfFkU/dLeoBe+LdKXNZXe95nNbtE39FhWb4EWTrSI8LPwrAptmT35fj1uyZdo
mGtuZ5Nrva1ceXfvNN8uU/cFuKWDM9sHEoejE2IrJeUQUn38KWBz7SknwgYpTzZe
Q6epufKt3JPNHwisuh6XYdT6LTGVib12FH5jB4lQZPOUZZD+w3IYYeb7j0Am5ioR
hS27YSrTSybcfQwZW6+2tVCjSMwqbg4olPa+Ve1SSVz5mPr24cq1K+cm+NPhkPIX
tU4WR9U2ZPPIe+9aykq+SSqPcGxXRI4koBeU8J/9NBMJiGfT8nHnCvOIe3E+bQpf
3Wu9tiIjIUUhC+yURVmyGmE/9AMA6jKRxehevQudcqrnS/lEVVjRsMIYd0XMkqh+
x7O0hkUGzTgOlzo1HquaBrJnXHlqlfI8EZTm6CbG5NMu1I7sGh3gwZ4ZhrVdwBkH
MidC55B0YGJeoHc0T04AOCItH2LO5KTvcfkmMOszTl7LUS0fzTHXeRULU/S6OOXb
VJzmzx5h7aaiKjlfMevD/sBUgcpG2tgJ/UqyUNa4x+psKXEPMvm0ZiG7vopia+7N
36VFsd+qRxCdpdi//r/u+flFps9ria1Yh7bzjwnspVzUyWk7ybhU7nja4QwCgZ1s
xHF8WtKBeZcoOqShgBaXA/1AmSZt3GuUGx9GCiGJFIgTvcO9hOsolTtQy33pDbBK
sDYd9Oq7TI7yHK40ZCkplmuKxc4ut/u8gVqzPBhLQAtCv42bNbwOwjqbJ+388DUs
8bcH/jW+wZO+UoHN45zGQsA3PRI6d4OeO3twnV/0Zh7e+KhVjhQJBLyVrQmQLppW
PebsLXZ0KvYy4Ia0rLuNCWnlbjpiNQisJcmIG/7KjbnKVAMZHKQZvAo99tZ7ogBG
VWLbN0QMovww2Sj2UDeTCpJSXDDI0ND23U7l7yhu3QBgrKazZGLxLn//B7kKUy/h
uQpaHXLDO9zrVBN2cMqC29jx/Ku+uz9YWcVW07iHoGxkiImSRBZwzsGv4+i32c8N
N3D55HJTCiU8SrRa4Mt4R+1MOXd9NQ30NYb13XnavGycWWzuqdeEgxxtHiQ4jBjp
68HoD9qsq0T7PO6KECY4hQGAMQ5JB35j+BoKpytEU4sWICoadcqPICY8bgN5NGbS
TFJ8v7zi7tOBjB1dmVv3Bebp32ji0/bwzLiHyZty805IkGlNGgAfWMrCOjHGIJBC
DVS9UdZARuWbfQmfMO7fihqOcCfUq5zgaoySKaNlVYczJDA0/WkmgiPi+Zts4kuI
neKYYXLsMltx2C8zJg6HyX8idXzeGyNwlUddCwB2IJzJFaBx2fmK4WXQ7FmQ0t38
WfHOX97ukfQPUvC3UGVbZHW10rYLEnBvsjY8+EMzfTJOKMCI41NE6KPK5JeDbbB5
3H98/BIoJLcTBefKrzJIGKCrvJADl6XZwiO3xCKRPv1i3+dKWhFBvd09UEb6cy1Q
swCKtJuAVPeFtJmzW9XGuhtVC/POXlyb4pfQMe/ecJGQ88439oco/3YIb95l1DWU
Xot0/gGJlP+Aovu8WYi188+YqwwwOOgPblz+7zQ4PPGnoIQzezm7iwhOrHzR0qUs
B3wwv+W2XiqbTkaQr0OAY7mRckMuZTcYOqekB2DY26/z1/RxDXkDRg3iQJclvhAe
Yp+aJcj+rcPL7/eEITrSik8twvgRwpSiuolkaNy2Y1Rq5prVaOCSPwG85RSkTDSV
xdkZDeqRObsrLo10ovmUeArI7OiDWwBixmUMj/tTcD+c+ky+FqqEFk13PiYWU8hu
j4qRpo6G8BinappWnRmLwA==
`protect END_PROTECTED
