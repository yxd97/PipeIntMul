`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tz8Yz2/ZYi1IGV4vJtru1LfzBVl4bcOE0AgZDEM7Uv0bPD0+TKbLQoTBkQfQ9mYs
rs2/p1LL4KCmrDT0GzJQg77VjGJRaQ4o3Y7O0l+9UOqslVm0pQflhYwBpBo1agKZ
OdX9qPQsbXT9gzg8MWLnzIki+mi+8wTLGwOyiviwAiSy9gKW1yle+WeI81qx134K
jDrAx76HTe3rHt+sUsb3tQ0f8uLaFXcQ0GxTtJFF+UqOLMAUt6Z5UAnHasfxSioF
1gCQfaUma6AaEUpQt5AVe8Cs9+zsXiKuRVYZJnidQ3yC1+d+CPUepdfrqEoO4jm0
KtmnwS0p4p6Jars7tvdjOqhm9wE1pNUdJ03PDdB+KDn1kHVHYd/2UTJ+41hx7Nn5
SUz532T5G4/9Ymq0RfPNSfDW4GGtAN+/oKasoSQy8pjVjcK98PcQhP/HjRvEloZs
BEBHcuF9Vvhnnit8t0Wk8WjqyWenR5qSlnXvJDvJ7Rem9NgSJJ4Bffw0lLKjtjc9
fhFX2E2sQLEQMpFLd468y/pGwwwIOUTybbSwlNLYqVAha8fBQLRHl73MtKrTVMK5
S0Xsjrpyzphpefi1ElgPzKakZ5E/Ze8OkRw7Tdx6BwOp6YO02jSX5p8k5UJrYKO+
YjxJ22Zqu4mSxe5Qx5DESvu5ucYLM0NmqUts+BYSWW0gKjR5DgjpHPX2FQHBBrfC
SETIfyHjQ9in2pB4e6uq/fn7GcoOIcLNuJzDYKOvaZOQ8WCC4c6JhQK/qyoKqRoa
CJLaDCyJIAWbpFDLJQU/c2uOqFFwlqGiFq9YaxiZdTRGm8gh1n73A/L/33G64pZL
QbC3lWGZOKzCDxp9nVySb9+FWhc/pRbaeLFDzSOmWoaWfAsFy/aIYQzkm5gtDzqU
ALklM3N6t1IvSXuLz8MZam0fP91AAjvqmgKk3FGpxfXwJIVvo6NwtZCUf3OWs6wG
M3uOgE/v20g4DbB5MGPdU7oeAwZSdnJfhMGwlwzEjuTdPAZL/VDpyI+3c+qGPv0Z
/VsSwZW05/lJESYUlodKgfad4AMmBe2cBJshizgkwM1yiE9++1PDMJS85ljcAODa
fdvf8lCyOeACBUQCOrpnRdPQQRCp+pTt4Sb71B4MGbnKomfHfs+PBMv8KgxOBYUc
V9/xFi2t50+BqlriBlyu/Ms8IdaZkGcftu9o6e1mC3CdZJZQIAvPDWIxcEd11+fp
q4u2DKKLvTmqYBaiAjr0atyE0r/h5x/57yMN9FBL3UBwzZvibRvke05G2094pvZk
iI73EbvvklqmR1I6oVG7UwhgfBaQH1n1E83kuQo4NzX6rXS1NDTGuZggav00uJH9
ijDJlWRL6uT3uwBNSNc58YkQlKsEKsGc0BD72eFCEKHbGYuUNQl/u7vV3RDEiF48
oKp+ZGAbAiZkBfY1qHpSb7YsixGMgWd1fpcE5hJ9066mZFIzHqfDHO9cgKO+x32m
bYbXBMH302T4ZSZdKxoUhz8PhAxdGQMcHzKZXbXTQrHrI7/X2huAPolAb05yJC3m
w7rDET/DOIEIsdFUV09F9/PiWt/pibW6VY/lgTH7n0QNS0J7HRX1SunGUpNEOv2B
uh7zqDjxbsxuGl30O0W96Uftg8ATHEYbGLVXSalr+GWv1uRB1jnUetzREboVjuud
zbGToJyB59tY9sn1Dzk9cc9mxmBzTq/kv/YHQUtXiNxoThJaHA+l+rES/HZXIK54
VJ8H7iFlcVHaBhD71W4pzt4Y8AJ1wHKa+Q3GCO2AwXGu4R/IBKMdbLSysoHznhJ4
BUwvlWsT3Lj+rYwUPylhsmGoRFg5DWIUTanSZH/7EO3x0I9wCmMrGDdWiGMD0beE
6KULPzzWXQgpLnp1uFKpJSHVWA5+cwgxVOVcXrhFfpAm+Zr5A7ze1agJg4H+LQdb
RVabfTqK7fIXvknY72XZYUOgE7n/vL7wPhljVae71Kk3lvhK2+pjtPXmYDDnH8x0
VAmBpyX5JE9klJyKQfW0+Udm7heaG2YnJaetad5CoBb3MRAjiws5uFOsEdLuoM9b
k6uqcHSYRCjaiLdPW8h9TJMf+M+5d+BoqutAdakreQenhDGe810Hi8x/0D3HDbTE
03y4Zgc0E5XjQNaG+ICsNpi9r90tD/UEHcQXO9dRsg5nVtJ6d5OuRJ+8a0zxdK94
+dWCQyzSxZztuwT6m0X7sW4kWVytqwKk43jGIRjtSqvShkhPqeQqpvxthUJB5Sr3
ac4+WLMemoXb7VJqkoD3oIJJQAzmhWSD8bNnPV9Bn0+swYW1XYcMafwq1zchisjp
ASiYl4IqQZlJMIwh6I88AfLZ63Aj0E99VM6YWnhs1l67MNUHAb1nGXfUIEisu3Dx
/Jj5x+rB1B+8/n1jrjKKyAoXb1OB6ZNPGKfPYEBaVWnM+3yKb/924T+zCU5kVrvF
c1tMTqhu4kADydPsRyz1PAh+e2Jmuv35UkedoJ6GhrKJ/Cji1DpcGlnmgwvFDJaj
9T/GRThSQXUNo9C0mdKELxUc7va3T9GzHl7akCM6SiA2T49qapXhzcI3qWl/wogK
0E62zKLflWu54Mcxyz+gHVw/rPNJtnHHtph1iUrfx2gsffARdpZVnAE1R+bEHy83
gwv7ppYUe2p4N0sDVkErTyHvWriIxsjr8BH88XfgO5LOgPqntBltVSGivtHk0blE
Qwpu+aeViJ+qByu4+wycRVV1ovSi0wnSYVDBhXQI3JROyI0MGmsq7Zhxj7DQVR5t
dwFvUH1UQyglMePMGfG1EclTPlfuUOEpdaEYJDfarwzGXm3r/iiUZXrGW1ycfU2V
2poLPWVs9zMgKC+/WfmiWgB7Vw6UQjfEncGTfx2aLpXXMDt10SKAd+JhBzsEgqfN
KmiBzJN21BEIgePohbRqJC9HP7FnqQBoiw/Dw+kFDfh8IuogYeFWMWc9+RDZbBML
0yeb3sYiHAkayy4aps8uJFwfbv8ITixloWj829NRgcf7yFaqhNMojEPXiZsc0wL7
AzKoShU88MPaPGrT0V5qFT6flXtPoEfj2YQBmHgfsmucWnydUpXodVGWYvkmvJas
bSvKJhDR1AnLaMBmo0/uQOxihV3kun037zokOrI+0TVQ21sAkQzhqhXr0xKD5hv/
9qvqdHdbFQEWBx+/gTTVASpxNv3nYqegVl6F182fiaoIDTLq0Brr7ndDWNKDU5jw
dvavgi6dwdDmsD6xAc9pnIaF95q8T9uukHO3x2RqrGVhMIu9ohG/IBaCX9Drte3c
/jUQnAY9Syw+ZQ4/RIiy8yAad9WPPqP6IweBr9ZkMV7a8k/AI/2to5NoiLG1ilYU
pk2DaDy81kozytZSXYz8SP4Ha/E9l3ppyhAZ8f6WIo0pA6deRvw4SQOdWwGMdcw/
04oyth7wBDm6nlEa0YbEttykwMdqjVZznAYkYkQ9rYF9iDedv/p5ksRwqqULoILr
AkSPLBA3/B6Y5Ll9zbOwCd86HOpbXcfJfcAd8aW/l7dkV3yEsgwCll6ZKqbCM1ft
Fkro1K1chf4Ax7xqDwmGI55UK7bRWtKkV0NBeUmRaiYQ2P9Hv6H90v0Q9Cx80zhQ
gbudrhF/mPhcJ0RU9z0B2Kq9t4ypOclyX8juqUfX1LfUzKM+uhU+d+c94zLF4RiP
voq50/C2NyUDJUX/HRvGE+DLGV41DSonHU0C6Jt3MH/aY8ClKlHtEC0D6uaNUc+G
TXX8ekRcT0OIVjxJSX1HjIDraaa033pIhyHq4qykOhF5HqLkd9tTk/n/fhXSp0Q0
dT1RiQySZ5Ni65a6sSFChDY/lf6lyc5FS/yJ/fNQr44pst+kfs1n+UBXLVelFDWx
MUp3vwMn06yo8dqgsOnobysgo2nhU9EaUCL6Eez9Cb6AjVkolu2onI/11GTfaL+s
yMrO3fIyrgytg0A+flmrurjE5s5T6L3mYurmBY1sODKPd2c0G1DnNyZNT1cazgNe
bVPq2VVaFb1e3gg6exXpYEZ6xKPqlF32xdu/tIJD3Bc8MEGouQlvjuQYJ6YVRUFs
qUH+To841wYSzko5Hyb01n6oYX2UM06zcJg3kHh+BwRhH8JZUQtZ/hhzQ/NB4bCU
0NzGVAqzxglsbBP6B6LdREUz//xHedZdfkPiZ3v1dwWl+wQ5cQXFELDqS7CuX6wp
p68FYMgQAcvO9XNJiIeimw==
`protect END_PROTECTED
