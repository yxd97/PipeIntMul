`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EsGbLhRZxPegejl/2NOQl9VrjujJOPEm7QGAXiR2ToVE6IRQx7Yp+drjGm9LQ6xK
S2he22TGhVCkU8zjB5f+dCTxLt9ap5y3hdCcugrjJRNufS3sib+ljDlgU7tq3afR
GIUH7xwtbCqEZ09xtm1lnZdzkfIXVg3FnGnA9yVjAb5cZY04p/6DOGqHRBVxb85l
mse2v4z3M8/TjpyrFkdFRBlNmHety9s2q5kR59E2hXypIV86MUC7Sn0HeWcxkzk/
dhnf3gYQ7G/yBdivxGyzLS88mAyJCrY6DypxYKwc7iAFvKJtGlQhF7IKJEiFzeaa
2DpeRaWg5ixp7IbVUSPcd++fZ1oMkjxGaejXsyGCDAbpVr1XlRbwUINw8lvvQRP6
FP9sKa4DvRtVMn9ytmjvi2ocS5kpT0FUtOz1gETzvfxaCnt6UjWiC1UnmrK1HZfl
1/CyR3fsAG1pgWou06naNxNQccap8lWbdfNdUyAkAptCh2zB6UEwE85SRopuS9of
3mMmBuZBqLdNGiYnQuYzFkWEM0L8IteUiGsI0wpiuA57TFz37DLZ4UAb04mpFsIM
x9iygcz/3uj64UNLKqy6Gj2iM9UnhBnUmDIV37ovJ6SbvjMg24xROez5txvFIgnS
HCqykRLPM8WubsrsPWijA/LUIYhCFrOVT4ZlkRG2TwBCyHIKZUuA4EcDhUTy0XHl
sUfUU93jO578Mev7h0RwRRO3KsXK33MqlTRiYpcAMCJ6XFp4nNTlJYBLWkj17QOD
s4KtZ/R9tatEfX5GEl1nLNmgYydMs6maQ33ODqpdXUiGi+LfDxkXdwwOapABcIuL
exHczkBg43YP5mLr4pgw/Ngr23lQwUmtSwDaakna4J42xE+ezba9rS7RQKJ5e6l1
VbERahFLNery6LEiOA58UFHGOM+4ejRHjUD5gaR5lROi4JGQ9pC+4EeAaWtQjtOL
0Zlej1CTtjhqRau+l1WDRmqY2e4iGF4VOsRpV9nXwBe8MK500JdW84qw24AyTCKR
RzdBVsYb0cWkgDbIo/pQIiw8ffCxbxIarq5rchCKl4It6C9wMIiT7oXFDu42Zsfs
Wi+pmZJwq8xPe5TSaxp0Dc5vs8TknBRwh8dMJSGk180M8ZBme0z/YmBfRJBe5NT4
taDnYSPN9g0YViT4A2jqyIMsMOvV6Zie0q+HtsP9KAVbCDRvi7ImPvdj6C/5IUhe
5yxqmqf7vwtwqw1V+iJedfe+0Pt+nrAjT8RsdozpNqkEeH19aiS0HZmBYDYaThY9
qwNH+PuYLfj22Xb6n/jU7e1YcwGG4Gf0lVY6vS2DbCAmW/ysYU3tSoG9LLQ8/zZC
kAXTzEN6REYtMEI3mZXXdhFmkV1vxG0nk+E82xW1h7ibGbpep0a9P3ieAokR8+Td
PD+xWR9Tsk8X3gesSH9+C8QM3h8ndpTUqvUhlslDbeyOf8Y+02OM/aAnWHqzwfQN
ax6wujZEfLFPv0ahFsaEHqgtMLrCC4XBEQZYDPz5dVCZd83+stFNh9GOLhaTM8yn
wK80O460graVdPYSyu+xz1pdsUw1oAJcCed9r5ygUNPfkt8nWDJlCBYyMI/HVKzi
juU76MieHID8jDBdz5Q5rv6FbsNDs08MSR/VuU9uIz9QYwmGmPAOqZASBwqct6X9
npg6rSfuhc6jJCIEslsIyZouoJBgJJrrxWxucCOrQi9izyLnXVS4E04kZzUmVqci
EIEr9ZYrPS9S0Ria4zUHrMlBLWQOITvV9ekNHUfT61GDqQwNXCH0/TDB+dzxzE0i
ZdEiPn9cSITyEMo40TnzgiYEaLFg2JGW+L0E4G9xfRDAR/ZQgnlC/4AyE3kg/Q9m
PMOMFNL27QXm3JnE5whK2a+Kho4vLbBWRk47HQ3yzr1bbuSo34tczx0AKLo1sqY8
1AjLEaTWkD6nKLAFLlpdhu3sdxmyy4NCYneeGzS47Xr+WPJDBulVufvOrLwzfDrz
MfcnvCJ4F+wOv+E56pXziXQ9eG4aoqDZi2h9qgRWnLsopcmEFjgog3vPU8MfwTcM
llBryVZoNJQNpDgyAhMgTS1bu1qJJkBnicHdEHGLL0uusetvbmo+3PwTA3RJ2VfY
RAYWdqiEvxdvEN6A8Nd3HIOWKwn0XEeuNCUu95LVlF1GEJdXg8zaIqCBv+ABPmbU
ITJPZNpCCPpHQmrsmSEvK17wSqlwJyeR1KY5Lw1WJG9EjYg3dEM7veYZJT8zPTvD
hbeP1E1dYcgZQf1dVF4I6qu79z9vuwIEhD/rArhZzoYhnjDY/GO34MmUacmCNEa+
Zyu9mKdi3s81Xmm+uOs6HNWDOPLK6om5i/dzPJjBLFmufmRSjDCopcExzQNmxcUu
GXKz2rRe+DeZrXdR7lk9H1/yji3PMzY1GcLVGpR8XqaxedeX6at9xkpGtCP6oMSE
jZXffgKZrsvvNXwX93C4n8vj0KXYYZcrmR8i0j8jXpYiD5jwrOBddY/+pJ6hZQsP
q7xs/eTKcAw/nXR79sKWYSV6PzTtpjk6VnZVnn7yfjzlTQRWkfzsAKDg1Erv44D1
dYZxSeFhvxcofZOtz93gmjAeRkYGKp+sVsPCz255coWRrdNEiBRGNxRGGwD3mh2D
1X82AJ7Dr21phajisaKyxKeaqcb5QLUt0y8vfSTkJzivM8rvnlql5WfQbRF3uWSB
vbVGTvtulQO31FHwRpy0BY3ucJoG0/RZrxUjVUPSHNp5AZ0Ro/VJRB92vkGMRCRT
BvVuiXJJzjaCBxCqODsAhV5+Qo5mweOIqB5LayOwNdPk17CjsRlzlxbbN+0elDoi
0u18vDg+irNd7FmtmJf4pvax71OP4f7KZXGAkJ6gOUa1lsrWC0GghBZrcvbGQMKC
Zm8YJZsU4ZE7PmwzgxKgIVvo0FdIjL08nJTXixQKllu8zJ56dJjQN4tXXV4xu1G1
gkh+o6RPG7b6V3HXtdmofabVL5PcuZzkmjtCzHkcIOlq4GmISg19VoDTinD5+nj+
U4l9YFqLgZa+57Xx5cODzpZkePIdKU9CqmrGUu8GO8qSms28x06N8OUs5YsprHcX
kQj8BZ+lkvkqqI7RN7oVHQuc16cUnV7pWuk1naJx6WX8qIae2XruMm5cR5pqrBbp
bTjZC3sfWj0CQJpViWY17Q7o9X5BJdDgOUEjaCPm4+bmWO3RdV4ppnw7fM1cEjsU
w/TO+ezHgSGc1/TZdhYZ/CCo8A8YCw0jwAm5vuZjGuPFtoKhyBaleJX+PQRwmSK7
ujj7cGa+kiwK+9I44fE2EOphcivIpFiBCWiUO0vHXSkqgOIp94MCJ9dHWUHVOBst
eqLvdYg5B8K+E3TfE6EzRL+ZUZi4CNhqbZnTJEHBIJrkBOEVk4N/DWpSMMDnl6GU
THoIoSEiDJR/V/8gey4wv9/OA9JxW5KlLYHGjp5trE1FvBYNltqXgNkRs5KJxQis
FP3Gj+Hz0V1JFlQ9N1oj2eDpwINQXNze3vs3k/aiYqeaccRM2LEpIpipG3kzOicV
gXxRm3xDWSc2zKaAWkuofExWPe9h+1XrGdy+tsHpIy0OAo8LWt3ykK5JmKVcQOJo
1IEsM1V2H+oQ+mNBiFTVOWQxaFVxJjLMvcIjpg+LuVc=
`protect END_PROTECTED
