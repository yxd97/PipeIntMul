`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p/6cbEd62ahMHkfcdJQp2BrZrPugxDfFZze+KFAa2lHrK4GIYk4a+hv73+Jqph7s
A52a/cjDLD22/9VxDBgijKQm88AiCSQ7PJqDIQpdiIyL2o3b+9GYRpdWln3/+XPv
RUUnh2AooaOx+p4ePl2AG56wvBUwE3awbodnsM8NXIbs970JxawP8/0nFtcaD2oc
VaC8Ydjdv8eFaA2JWv0sgwiOP1+csm7bV7jGSF5Cp9MtnKbf48GXmjhaxIQwBqCT
k4epVHHvSXeibUTTOkcsKHXA2vrKvaFJtMHpBAOlfhk=
`protect END_PROTECTED
