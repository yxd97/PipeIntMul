`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+XCbQ+LiCI7kDT9hWItEC5a2HdiLt1Qw7opkcqyZAVhJ4nkvJVaRGUcaClQVEme
UqbVjItDwjV70p7yM8Ao9XrJGtCbyr8U5L8HBkvT3N09/okc9ZdcZx2GAU6A5l92
h4etcWhlTyA9YZpz+TD18o3vDlBoCG9g15fLOckwF3C4T8b5jwqNqIbYKmacblhX
4qj29DvJBfdd5ImkkNHjx5dCwgJjc+JsybfLZ9NrXsCvQ1RfdAQlcDvCyUeLX9O9
aRoKs/o3C+p500sRnC94TnPJCp9ZuBJgUmXJi0vRfO0ZAQbDdBayF89UJOYW/7hu
m8NscWsh4Kx996XjT6ks8yv7MfoPThDLGETBa/J5Pbw95pDPIwxsQLkdnzbn/SfC
RBqXJJOBIbYKEkd367LbIbKDWpqaPQL1MusxXtBfp1fg/jDWGFRNWFn2T04+asxh
t1kddDauXCVPFUrGfjZBbv2zHHrej/zrn5khuhbKuTxDUAdfgVfapEfEDiMnOCFE
n3j8FqW1NtxTrgFk/axQL4a3KuoWC+6MfrBL6S1RDy6bi9Lb6/Av9xXE8xjHzs4r
3w61Qihw7HgBIYPHZxrrsJXLcKIYWca4TFpzQbpjSbjs5YMKwAvs/XT+AafWypUc
MWGYlpsZQOYw4zaggBOpGVMAL5lakMljTSr3FVMM76vYrjRpANiXKi1u6sUNr3WW
AHfU9VT0oFwq68BAtg89ekOBtUeWiwo77Ezlh0O6flY=
`protect END_PROTECTED
