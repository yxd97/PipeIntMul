`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pa1hG4SQGqwrtmHdqppO6/yuVhxJF18gi0DdAwQwRzsmirHUdy71Jks6nWETVU6R
71Ey6KCdiubmn7YM7LE0/DvQGXlIB+iHOn+8YwAPoFZGSIphMtsLSSQE394FBmOy
i6haXgPzlTYKxKkWYaS3E7DuWOzUbQUjuDbDK0eEJcXRg+J0pIPHaNhdIQ/sAsiX
DJWvSqZexlLR9of94+vN67FmGMpoYHm8sr7UPKaNdpUyxP5XLbtMB+Z2L/nSEl0R
3WL4XIUARTP4xaZmsBSfnT6C2frOgEqceI9sbBrv51PU9tPmcEy9KJqW4AASBKIr
xA09rk6EriFq/JmVj/F2+5Y/68MyS5Lr7f1dweCIRE4T5h2vQcHMZvcmMigp5YaV
/iofnKNAu8U8YLubvExhs2U73MdtoXazc3RKOVl8oCc=
`protect END_PROTECTED
