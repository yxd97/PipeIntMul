library verilog;
use verilog.vl_types.all;
entity IBUFG_SSTL3_II_DCI is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUFG_SSTL3_II_DCI;
