`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mx3h1vTIdx1fMA8oV8WA8/suk4v4/T+aHyCYmNWXQvxVfNbcykb/ZPU5RsaXtnZf
CkOZ+bpOLsnBkwrbfgsUqIqEHXTslNgEhV9dcrt+bGdXjFQhQY9uDzs9WrOguLp0
+jDQL8jsvFXzyoPAJiFPC+0YWQGtFB+H3XfKkS6NGTrhqsIzpQ4g2bkea+LarcHs
7O2bDR/+61Hk40ZVViUGh/WbupJ2+qWYYWKUPQT4evCbpTGKsWVNAIzYvcuY2CC9
jB+BRf8ZXLNDr8Rq/RXJvjSUd5Lv2/tc4lWnEiu41q4XL8hGyrJ55NicBdaagAUB
z4wnYd6ejMU4TRZ042BycQ==
`protect END_PROTECTED
