`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NzXxH14//RWKxUj105CX/4XGraO2isESMWBSJnRZRvRd/+DMgycGabIRGSl9ZcyX
UHGSyKR+Ur9myNcu7sod4CwPlzmdTyV9swoICM0RAglS///LqC/kQsfev/y9gbEv
mKSAWgbYcL8GiEsWoI3tXDP7CiVZ6iZjAzYGyusUEOJGsEnXzFyoTMr7v+QClDEK
heDqe0qQHQomU1HGMYZYV4f+l2wZFCr1JP4N2p9zpfEsOxNTzsVbG+A2Xhx7VerR
1B2ZmojWYMGGcE94OvhayUaN7ti33yofkYdyS9Uf4sybhsdMiLURARm7dEw3TO+d
4KXgDom+4yN0j3j8wr9oYESHMDu6GiU+W1glTPGrwZSXUYy2KONoyJVYldem7goE
V++TxhiN+azRhPfuwQfd7CADMmugjiC4bYCnMqav3iI=
`protect END_PROTECTED
