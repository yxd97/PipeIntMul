`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/yn6tQo8NbkOU7Eci8POxabjrVmBEXg9HYroXIOI9GBRm+fKRtU0ZlmUPy7j5LyM
/uhUtVSIGDG0QE6v3nCprAqL+Cv3N2CdhTGn3hb9eC+EEbtq8EaGUg/stweuia7A
TT3jwd5YI+Ke6Q/pTGhfYFxid95CS7DIH8kEwLNIIYUTZ11gVENQObjzebK/vKv6
+YUjA/e9bS7+taLgDBMQO0pvGlGseFPTK7LqkQyDD/zW7CpdQPYc8DEcggxOa4zz
+0YIydmc43tuo6PMSGhnjsH+etLVFjz61fsgl12crzyDLesYOKUHomHrYmL1ZgR8
rFqRJtTiinlxX3mIpEA/WELWr8sLxtk/OxXbUhrlZQj6aO+j94RSbQcaSEWQN8/2
j3VYZQor/Nd0a06HZhZpMEadOACmvnlIrfTyBHGjn3nAV1p2CwaX72xzi6q5PJRS
rFjbmmrkKYZ38rMEZfPsNvM0L9f/9FLrIyC2l8JLz68=
`protect END_PROTECTED
