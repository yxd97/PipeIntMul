`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JmzIbay2NhI0Jpu9MNv403rtFOVuoiCCXzV4X3Au3bQqCw98s/D7G3UYCnRwetPD
Ybyg1BypE7Fsznc692z0UbcrC3txXrMoFpfEu3o3tuLY6zt0Ebtdy7YZiktwR9Rg
kiX5S4nRZyoLIA0fhhzsbPRrLjOFYK0ZLjY6uGpI4PXEegvov4ovnhpM1ciNvs6e
m6z8gHSe9/54H0WitvLpn54NoAnmPeP5mGh08uZYRxfXw9AqcRXHEPQDEfyua0/m
psKSQXK0q8ich3z2h84+fZUXL+IheoGcb1NFrKrKI/FVpyveKhWfeoyBY8Md6wsh
d+iFN7qRMKMzm4vHzZpV1FonGZBSwsJmqGVP7IOudrzPpNVOGS9i2au96w+pz++x
fxD0/vTVZUiZNCb7lWda33d4ACH3KT1XolS4iECjcSWjl0UttzJvS5rrMzNYuJEu
ZyTF/Pbx7j+Mo0VwlSlNpLAbFf8N1MMgIW/JbSg3AzNtf5QSUrRlxwrF6K3NxEq0
XP/lGJBECZVoxTK/00eNy+ZHaWpdqgW9sHpVQwiEaFXn60vgStEsfMS5LXKCeXVb
owqju9B+BJtrOLD55J/AuKaRyyrkqJ1Kird9jRFG1rt5IY1jCcGRnEeETgNi6Tmb
zJ5XNweduAN3HaY0d5d2ij5yYBm2Uv1G7c4pvcBgg3+glyH6n4mpGwm+t3emOIUZ
9e4L+AD1zPj7q3tKE/SlIJ87vj6hvD9e9LvQpK3iSl7xSlu1zX+pdivVhSptA10m
KLXOVjeYktfWJLQeMw7BVcVzzm7q6ifG4kDq+zdVkPBfSe1+ck/GPKC5BZe2p+ja
8B+xqReh/vv9cGpdbXoQIzLS1O0e/qOTG6WkhXNve3tLKHztpZcgEfNOIXmT/HwQ
bvJWIkAMAWzHFkgxdQjhp3iwtNvheNUorOuvXPGpfcWjxTlcUn2r6wHIJNcbB4Q6
/J/otQHRvrBZhZ7VBPDUu7L4fk2fqrkvUuTOx/fT+3Ul4J8IrJV2DRiApmmyP8H5
I6WFIgTmzILC9hSYDj58qfPI2/dW+T/Hnes4gGg3V8WXhL8K3koySlqdZ6QbHCK5
bUbCRz9XGMUlILwg4uKmv2WrqjgNGVvPW3ebDDxMy2GsjVJ9ErjqBxH10QFLwsqz
xS18y16GxcImazz6SmqspRz6rM5Rm4e+6xIL2qYEf/Ga5gXLRiIvgVbgjH5xIJvn
ELf1XeNL7Ah/tepzzUFXY0wm6WmdOTcNyU23Uz89z26Ti2NT523KQK2rRNBOmupj
tzu451/U0lS2ivW4J5vLnf5dTjMAs7PQF8TDdSqh1kPffLCcAvlO1djUIPE1coj1
E+jQQOcEyh2EQGBTphJs2Vdin07OZs+eHPplq267G2TEthrUEHMPVCC6jjAZxoxG
1pEFuPxG+TpV3xAV64Dc7rcUvjfiy5izkQMfiImy65invAJxIzkaAnNnQcAEPgn6
RhwmsXaQ/xx1QuXgM/kQzUwG3OZ18F8gQQR4fdpGolg5Oa19v5Y3v1cFfBSEETxL
AA6/Zrv3EBtm+Xv8t2/MM4oFkkvnIRUSrEaug3nNHZ47M5QFKHX+lzqiJ4PxyDcx
T5+nn7Iz8oOSEhTqdyRA0LpLwJfnEAGAKd4IBI3elzhuz30AD8+YYomdS6dkpXZW
dOGeDIc6LYBIJ6cvqPrqkxWOkUWe+9a2Z5xfM9O5rEzv0/TTJLZ8zCBDxRoej1Cj
gr9vXM79pwUciorHTzzXWdHzqS0PGQ6bV16y/6TJQRkOYKnytipQJgh4vTmUs77z
1sWhCv0XxDLbcXaEwtToAq7B2E2qsFl2D44/lN8lrwa70gd4tm3y+H4gZBb6rSa4
QUrk5VFaBrsxa8tepMURyW/rRw8EzlSclESd5pyR6Xzw4sQDqQ9Ag9Hx8gxQG7V9
x9rHKooq/P2ushj6U5Q4OS/s7kwny75sInkLaRUPR6enYVB0qpfeKOTuUYsw8bkZ
rTEyRWKjpfqUcmWEHWAEQWWA5UOGD1n28jyL4BKrrZQpzVsBWYdK8msqR7STllOo
Ej0nMwWpRy05oKe1+ncXd8SGUdhSOGQr+hHlJ28JxE1OG526Y4xWM9dlDmNJpZZ0
zBTMBA84FuMLf/VDP8UyeSwFKvszH7V/pJe/nMpSt0Hx2KihplBHk2ztIinaLoDb
zbyy7ohfUMLaoLnB5xP8C3FDUkqVfgSvPHYWM0o8p5ygQDac3hNtj2/NBJ0M9C1d
2ZOFb5M8aGRcy2paaPZ1MLScukcspeYzEU7HdSoiUjosBl42HqZ0fGBBc7j8hmCl
mGOYadcef6WGHM59vp0Sa1ErnsYHgo/4xKGUcVZb5BSewUK24wFgD8zTMnV9PI8Z
aYhn1fKqhnruKVVWHS6TeL6JDGmv8Vdkdl51uT9k5w+m9mYeCnKe9zy8yWArBmPH
DNfTScfekXDHxBHR5mgRvoldEDMCm85rLj/bOZQw6kGNm7CyaWugVcqhRp4HenrU
0DG+u6U8CzZGco+m0KZCFS+KE5PpQDJuDqJIEe1tsbnVoguNXYCkHWy2ckymfM1q
jopeTsYlhnek5y65Ws2EQAn7agr6m9zhcApFZmRoFmU8n4OFITpaw3DUVGw99ni+
4SwtfaWvChZKk7/02i/EGlgHu1nPhaZwsp6+8DesTMBF/Oiz5i04KwZycDrdvSKN
hAQotQRyfWNtavP6IVHcNCOJBCAkKftPlP8XKbduU98adHP8/0qrHW0f+OmLZkGO
bCLC69PBfJN/mAUY6IuTiuE0nMgPdk20mov3MNsPmldNBsE5SFIuq5RzbtNpsvpk
VwxJTpo2Biq3Gx8BF45TESuPy4MOTAkxfG6RpBZ5Yslt0r3l3oO6F3MGQYYEpq5H
Q4A288DwameFnoc5ApmS/H0vKSQ9tJiqxbL4DMGQNmSj6rU31qP5C1K6f4hbtjvY
LprXTqjNiiL0t8iGR6uRbWasTSL0A2r0Mc3km1NnpsRkF9FcbLi+nZpK6qQw5XqH
NxA8NZYBJR9Gfk9eNGLgS/qza2TT7p2yxAbnuXA+MJU3HZ/NRDtdsxYo05oJWpFx
BOcMwICauDO0QwzWvOlJCPVqmj+vyjCH1gwXN1Mg4IHj/WDsWdrCrXPZoTaXQSIv
MfYKPn/j7C2a2xmvShA5f5p59geGd0ANrgjx/IWJ35cDVko8qtMl2Ln0pzPAXMiT
Ji41770o+zdd/wlvPGA6lWoMdUlahnhnBPV/dqQMk/+VY08vmni62s5KJWMENkal
xRcCmwncBB4bgMQRaejTjOoK5gEuqTObmTupgwdI8oIf//kuil3m6Zn1dsWmlrkV
S4QYqDTP/71DQIvHlYN34YwEtRo1VozENzoDTi3OUtHcntZkO3ZlgRftSbKOPdiF
IOq6OzQI731JIW9o5zhznsFSQfaCnXK2/UGdZjJzhkwoSzU22qfMVE5fLdRdOYhD
NOqXjXHrFWZ+H6WIlq9+9ooOzbapoenWgQplf8lTd5O1+sfkxPFePxt3XheoXsYD
z33L4/pU+z6L0NJyYOJIBneCHu/p/cR/KvWom/tSeeEU8KHHr24ARJB2lsdgen2d
0a2I/Czdc3lurS9riGCZXjGZYLL6NJTUOM4ZtqBbvfFoVMdcJyM8pRMn1xEOC5vQ
0P08vfQRi9Zfyku8MkNReK+ai2MPd9xNAEPPyEkQLCi0/sxgf+wQFZQQoJEexzRW
QpZPW2KWDwo0PUD2uj9sKCkFWZ9yh32gyebX7VGPxpkuhbcB2Auubf2kR91/IWbE
QqaXKHJJEMjSzGwtb3Om0QwDbwpBeddRYM/+SE/wm/5mQymXUe5YApLsuRkDYdZs
xRHabbAFGu6uJcsX8zjvS+w+/tu7aupWHlj8zWoIgmMpvg2MRySq2U50dddm3fPN
euUf6GRUJb3cB/nLd8eOVxBlt3gf3oQCYqOVIdkbiwj4dpwqi4TnEFzgNSjugX9T
sMaQ1EIPuNkaSLmyjEOnAe8hUWTafyQaHwXFTqiVDJGU/ny/qrrLU3WgwWojhmfk
5a0qKXPhsmvNGXIdzYjoaAhBr1pwyOACxcYt/jmhs8bBk/G2xAiMOxfbnrWWQ9Ms
A8IIFtNsAnY9o15HxsyKWhcBqEmcfnYJdtEKBU7W0fjM2dn8IgJzA2ey2sW3Lc/S
B7b7Q5M4DeV8TtwelWdNXaS7YlXPkyEBw3NIOq8T+KaZuuPa1pfm+puN2rU/4+Sh
Px9ZIUfbIwbHIKXC0unjVdn1U6TNfjTpobwqvCikkT+kTdrGP/CeoAsIObKgOBam
o1BSBDxJQjjVw2L8yk8/WqDYj4SlbA7szP9sXsVMoQ6AVFUM4Dr34BfB0puUOA38
/FCa9Sb2bMGMqaJskjW2aFZnh2bNxZ/uFoTZQMlvwB1+jzT8Z05batDzC6C1sJ4E
4s1cG3GiGSTpPbpJmgF80GvpZNdvBMefjG4ElLylQPM6dtcqiSee5PlWx5LuhPES
e7+E5112KbJilBYd08dgyFHmnMAxP7IyJLLJVrLTBKAxVstqeQxj8IAtNiP2jZBg
TVuN7lffPZx6HPH0qh5jYKTI907VWv9KS7+KfxhdFL/nXPvS2AfDP06lbqp+1aT+
t3Z3NUc5nE+/SsV2HxpYsOeXNtZIIi4/5BnX5Ne6blztadKFVdpwHk8FOEVCdOK9
3s5gI+GgljhyFiseCLQS6zzkVm1YrUDQSdcUc75hWRgQV+qukqAzX6WGe6lUi1Yh
jqLOLDeh03zMxhEv6d5E5YJm2R1V0lRooBQntXt8VfmrySNIz5dtwa98H1hRZ8ya
KBpOXKSdXw5KRyF8v8yb5jVJ5gQNXnWL7OhealQIfoo0yYGd7A9DSoal1EVnvodm
SUorD86UglO3THYbQux/g4Vw+oD/TMMPrM069JSFUm94nSlTToqEUZQFX5L1pF1m
34PLhL+LcIR8eR+RtrlITx55lO+FS8eVxhn0oLmteYG2B7LM7qGhYsqTKhYC9csJ
ijT/uui6IzO2RREzeFhf/bgLM1WJ6al+l1+tF9DnfUoSjsMo+GrppxJQMWGQ9nxg
mudisP2ayy5jBOeEEjKF5E64BQ4qLjMgkWo3a7soV7+t0SKHQcT/itkGApVh8tox
Azpyf+SISlg5BVEBzKxFxALd/QWXlpY4bxL8r9J6KzNH4Mg638RRKAltLGMmEVh/
gVnUcX8gYtSe+SUNlVHLuMY62ZhP9cUk/4K8clX+SA7/2KCgBddZXAjAK6HXT7Q9
Zve0pLSXNf5dTS+PVJLD0xzJOwZZ4PuFW7T0efVlnoBBzcrILjhhZFCYuamF6FIs
hecLa4OVe7Sco6kOt5C226hKn/CgROjKJHPeYW17LDSSn4HbGnEVW9EeYTeW4V0G
F3Rvy+sgPOrzMyXesvaxeEcPnKLMypevcUzTmHk5LTJ4frPidrmuEjuQ4sSGDNjn
1OtHdacg0GkDm9Y+1UbhqBpM40mxGxzdzmik+HnKql+5SogE2GOs6jbUsY4sr8HI
w/YfPfwSqLU0SyVgs9mqSx9yA2zJM/Yvk/RKavQziEJj2KPMl5eaMdt7D/W2mJKy
3cE30ujSuLR5qy/j6kRO/iMLGUAm7iFsBMpWulsX55K0KI9Ot8k7tfXZRU81qGhf
DL/MSop0Z3VxjVLKRpyuPor6Y/3hJWGOhu54owq/sEClGZn+SvA3Gx6Rw01qjtkO
TwBSxxxVh1cnOjvRVE8Qy9XtL9yUCHpq5BIxHjm9o/YPaDjd3bn7Nl2CVz4lqIW0
K/kpFvA3XGWThQt+2bUP5ICD3Cq8hRMcndCEdD9q5IR3NQIc/rQWhs5oE5l9Ea5e
CGlDkGK7HsoBHE5eFZLUK/Au9bOw+WZXxUsQ204ojAGFFRkhK5J3MO1r6IzxSNHl
3VNjZWfJkarUkQRcJc82ZYWNXtNyS47gPVN0c5HClace8NzKVL/ZCHqc5oFlC5kn
/45T/EqdeW0BoI3RZfQaQdk+SBjWQXJYYrBP142n8JKoxkJ/u56YDhSK/Yih2T+/
BbkdfxN8GEraiSos4QjDj2Tuks+mr//UDTcpoxFk7mlFYSFAQQXEEJ7oFL2s2pKB
R3CY1G8I0Pdep+wTaUXs7y3fQZ6ua3QyT5gZCTHmHp85lo55e+PZ6Q3MU2VFzFNQ
vdlrKvlraOKfDXkTPyBBw4mBDVpvYEhj7dhB3N4a9CfRVVBKsgxD66p2vbh5UYU4
ZIvisdt8tTR25TxiXctRq8A1fM2Dba/gb09xU0iJS+2MFQrt51/jiRi1mioKSvEH
mcLARfCyMqnmNhhHdCg5YxJ5EtRIZNrFFdGrsFoiW5Ts0v2zbe/Naom9JgpsXPDR
0xkS/b4d4bKM1azuVAoTKjBwbxiKFU3gFlbUsd+9iXFFv7NpiFWWrV6fgmaEfMac
NvJVAr5xNE5MybOXEa0k76IEXQWQkn8qjLqzCafs4VMW9llCXZixk82tVJOjgODi
Hd47bXTbn4KBDp0S+bFrtxA9DZ4tB+b+iMC0QN+GfUdXpCWowQjl1KF4CNS3ZOVi
OQc9EyrQTTxYNiu/CyiGs4J5qYvmQoimCYUO9LlJyuCopPdOXWp35RIqsUre0/z2
4OzY4CILo6xX+EQpq6CQFyY5FgcU2V7CE3AAX3HMQWevSrfiOAEEQBlt3xO8LxuL
ApOPPahXTgpg3tM4iNsLEkSpmCxXMww6WoDXGv8ZXt5NzLF0Sok7p6Lr8vt35+9o
/Nkmp6AzfD7aOIMWKDHUHbtfepmuvsShCnqvnvE2qGqgWjeJKNdy9fuz4pxx6K1U
KaSigDVW32Z/aYbxLCYhf3nU5LgiXNMi9JP0x36qgwVaQVRi6adfSXxX1iZoxE5z
gZNyKG+FJ9hsIbxuE73TQksmEuBR9Yhnsan8B+lCjaEuCKKaDsEDJon54pc+atu5
422Jm6/BKor+mNOMx6wSf+eHTc1gHWD/fZB1uYCrPoiaA9OHBOH7uEZCE/GezXeW
oq77hVZ/iK9WtyplpdGe7baT3oIKNizZp4EAF+PwoYO3a0laqQN2+IQoBYbXS/1U
8CWkFRgMB5CvJcK09wLkmdCK6hbszNlHE5LmrKzbmQ4sz37WwBMvNsWipQ8uVonM
oc85BW2VBJcjJH6nTgcnVvFnr7I5hTR2T6YIm0jJLz1dnRxt6t/pgdnl8pwH5YvW
E6iDipRpysu0kitcUlDUwukYc3OC1a8aQmQ2XblvtYZa12qoNRifyIjHIitsS1nT
a6OzpK4BZ9w5llVeZ+vATFzBosxba9769VM78jE+YQEzgrSwcK880eZNWt57kdA+
W+i6/NVQCkv/hkbg/nDIK/7cgepILT2KoN5ZUs/BW26MgTg/iSWLNFC/lKTODCw8
2InxBjoCIAFSDQ9LPLAtHjgxp+yZv9mqxu6kJjVgWtJDoeZPG2LQ02dk7AWMpzkX
VN8yNIL9MF1n8WO3mSUtckC6HnPZW/0mss9Sn0MSgH38nTTRNAi1kgS8JW6Cq4hq
xPKuGj1nvPopYsW6CqXLHaQlj905I/fKOasX4nYozuJdzyXnQj26F2BYq3BHiQEC
52GY3IKAFvaAk4fpI4PsXnj2zSuqurrjjJoNFjumn1RUPxBMJIhnGeonPP/4inz6
rMbHfUW/AMB85Agb0isHC3YglEBl9XkmBDotYJZIJx0hZQK02kqXEek4Vbcm99Rd
teqh1HXWHkIjHEjA29pVE6V71hnXMxPy7G212allT31Af8qEBXZP1sUwi4wsffCU
si1OGpgKxRg3MNUh1pGbYPH9x+eF94dW5/KTV//kEDIgciAKo4unIuD9zE1lFT3R
8TzBINVFVoBPXN/BRLIV3+njjSb8OA1xN91ngX6gTuMwSw/DD/sxaSPSO+lAmRJU
ZLP6OVtptEXin53lnsPj2Uc0p1jDAb1RXDBkj7ieDxa3sQ/gQ/7mPyLWngx28IAv
UL2tro+D1EWhOQab51D/LEdfw6okHJanuu91ksYHHHhRZ4o8fnMVl5HV/df0EIKs
LJMQv2LLbwUHM1lou8tV6UqA/LHdSOfjVnW8ioY62kE5kTSCjvhAJ/PvYqGtdxNW
z26hdoeLlZ8iR6ZV58U8qFzbjA+d61ZZpG2rLscREiOcvEPBq7TnifZ3I8dORNZE
NkLn3TqL+DYMpwLFCr93AXIzqqNrH7/0Qi1Mq4s78SJozwk9l/zZZPnszKo4tJnt
jFwTepBg2ugYA/GJvWmpit3tQ833kEAezGDrWdbZGvUF46BLn6qyRRpxfYTrEnuH
X3fwvOi3KpOi96nRxmIPcjXzZtx0A+1uy0O7LetfLSyP+0OjKz8f55LyWgaeErCN
+7S6Cf2ddOs7sZiV4UjRgWQxw3QonoMA9ruCHRgPsEFNxXpowRiwGb07yvDVjQWo
OdwJGImuKpyw5H4sH199bKknPFtTG+fjlDlNfK7nCBJrN7kJKJwXAwf815v2wghW
c5SzmDVAx5kTR8k4QRw7JqTOs8m7Q1aeSt2lhCfml6QBYRml/LuTmBH5dvzk+ZKi
6oT6eWX/xhv1E3fMyjZ2WXxc7NhaxmikZktH6YSBdJQmFsVk6k+BJo35ZN5JV0pc
pKJOiNW6OeRHGKfCqRIAfrmawj4iD9TrCNDttJdSTYc0oXDHMWYhO5xDitJkLcIt
YJIRUJRh0xvSSvSWGi2adE1+klihtWopxB7N0EzraGqx6exsZsnIFyrmuFFWYjrB
9LazH71RlOTn7zovUmrdEEGbsCICdomE60Bq5cI85uQsxZa37YSgTBqeNP2a6wJx
oRw3xB0Kugbm8NtXE7pumXyaCbJ7TgfELqUYdj5q/kiB/LP2NG8Qer5RVORwLTsl
N6K52xKdQHKPVW9LcmyTJO3sA8LVRWt28W4wqJS1+zmH6snf0rlwAF/ETNfiY/hL
3w0y2ehZlVyucVMyuOSaQmJJ62qWFLj/qCJdrWbo4B2COQRC6NDSo0DdTcj91O8k
FaB+H5jmlql3A16IMDy9JYHBm0uBbg0PozmGVZARWTR7OiyC+KgUCNaPKQM7VZKv
idGA8lYk3pns4o3Ot9gfVcyq53CSZyYH5GdIgV7ew960ywo4zz+LoICDin/izj1s
/X9tNDPZOhdKwcJqv8B/R6PmS8w849BZla+HmrHSItoe+eUcK50Inu4LeTE8BJ+G
/wkWCZF/Kb5oMwXl9yjylkI/GMvJ0/oja30DKCkQul29Wip6pBvbhuMvrhJ9xml+
C/LzaM7j82C8qyr7mTt8wncQ2tsRLZdRmJvHlXRZMTJa36ibTvhJKx5J1JUTqPfz
bxR3TpwClnjX2zY9M87OsH3VigvlzSB4JuvzV4U3fk0SJzfP7yR8Csf0KO5NqAL2
IuezBixboal9pHwGZMaEd8XCCN1qXOyQ+9CHGvmF2AXxGtINKwuNIQonEwCudnTC
XURRfmPlgMEkUi488OBCm08agekAddfgY1CPGugWALnfz/DPKJHaO3Gzi1Ssp2yB
pfnIUIfPwyKPCQPUUUXHKdga/KkAU7YdvpkUmK1W+14gxsrki9GFp5HYt0JvsWuj
txLNR/cYvSe5vnt1NAToz039o95XQDBmXYExkozOqs06pGkZtLY/0L6GdA+4snd3
oUvJzgr1VwEwgC8th/dpxu92dZ2XYom4q+VXuGebr9pIaiXn6KHOliwyzaR1JNU1
Xq7xLQR1sMOlp372XaTLOtOltCFfPxMVU48dGn5dRamNfZSxWN9pfeiW+0gZ5Iqc
DLMyDL9sSOzwLQd1V2/IiVws2kvxX5U/PYqne2RnxYsUkpLzwJq+3szxmdZAYcTP
6M0qOl1EprkaVCnpVjWzHTQxdJTRROA9lRFDinYM4rbbAnH9Mv6Kqb8WFnGJfqsM
ryEnGUBYFvWmFl9Sxm+lP8Of34IXLNhQvUjYxa53Hn0hNPvXETshwmaXZ0Nxlf8e
Ms21sDkEqJ15A1ZLk7/W0sVo3njS6xF54JoTaOBGKbD7SW4X7BWB7cl1n7wvuBhP
hJ+616BHm3vparFnFSEvM5cHD/Rhm89GcDaGLA1msueaY7/7SiK96YW6OcA9+alq
mMte9xM1SZi7TWhm2Du6MvLLir4E5WY4/JeLnOEuSMO6X22GnmxVvIQdUgLedfNW
As0jCuARW8xc2Kf+DQ+KnmLezjt8VNJ8jY6RAdBQdnHcHO6+L6vKwyjRgVj975wb
TYt7PJ5U5X4SQ0lpe+4UeSDHUoSuFse6wsFLGXFWaHRb+wbYRkPmctY6OuEjnjrQ
QnCIk4sX7G1aK3v+GgMh2xOHZzTv22Ey6IMEbAFaFI133uDFfyzFKBU9ZtB+PUMZ
qPMTtgYdk7pUbx+2loIUFyhfAG1DFTML3mOdcmNMb36LbvdCGVGn6T2TSxhspfe8
ZRTAewDIgMEOE8GURqVooya0g00qyyBvI70HWzkl68FNbigfODshbbTTUbqEjgrQ
ehobLK/Ua313BDWf0gaI3Nbu8Jfu18zdeBPaq5cQ9Wq7Cgk6G3/Sv7kDkNvTmuwA
AcSiGPqP2In0jvBXFqnRb6i5VnThPZdVlp93nNavtVlLLSXCHPcEqwfnjS8wkMmG
FoUnNdtNK/ji2lj3N/xFViPoctC9/bp1wLn3EA013iFkUOJfCuHcoGgmtDqSIduk
vBP/UKQydsUrzDihWLQNeXe5sfGt8ku/5c8+Y5B+9L3LNYvjikmRniq8OnLVrAKW
1oXk8WJIaC5v/hQQdto1TZ9QBdih1WA6Eh9Z5wdBdhCLR3a6vnOmas2+Pn9eqPrl
I70RI8lq2ab9R0cZuku8keu5TlT5CoCbifBgh2evajgH+LoO6626YU8utc71303z
Paoh9/7yDnv1rTzqMJu2oXuJbIFiA340rakYToABtgZvPcpVL7PEzIwQyNqmq5gR
bgAj6xt8aY3TMqmLVvZqqVyHul731fLEw2Xkm0qSNeLk/wmvw1u6louW2USX8wnX
CnLv7evGvCb2zzFPdE6O116OJpUXLSHMzUJ4HBTHS4UMhv5VfsUvTg8A4CoZI4Mu
bciZB0TwJrO1/PzEDzWDXnzmBKGtkW/RPMLQosG0NcGS7CP0oYjTOHfKt+sOXuli
7SY/8gjq21JnW95OcarR3BZd8r9Ieb9xeFRaiuUbzYP7lFXYr/6rXRkgyRd0hawI
NhcllKVj5d050XbhpzF9QjqOOZIAHnSSd9RjNHToc0bAjpX2rgsZOO7GV4nCLVu0
LKr/TaP61y6kQJhqK8uZsxM2NnfFSG/yVrA8z+9EA2kBBu3AtWBCFeB/6wFYsS+A
CGV/c3bn1pgbeA9pzoq+L9r6jQ/psdvauuABsFA6rlJ8XuhLp879UPtqV+2uXnOr
V1Q5tfaBqnw94Mrwg60g9BuxriM5mxhQzTroVJ8AUp0I0gW+6Td6/bTGPf9mZj3g
GDDRjjJpQrJWMYRCF9JJqj2G/vlZtC+3uAReYeJmPrOxM8Stciaa3JDVCIDo45r8
hzd/yKz7FViYJhWg3WyM8baBp6CXrzHwrxbSA/52WMj9bF8a0TBtudShfeD8F/iR
e8MsKn0cLqM5K5CN0uTjVTR7RlI0iHveLvVqfp8AtjdfI0+GPzHB97sFKdEDmWyx
jn4LQkQuyaPW/nedWtUeZnl0hQF3OM6Vg861ROBTZpC6J2xo7CcsjenqZurL0hZh
B6w5DYxF0PXiohVEgTFR9M6LG2+r5nOiEObQBTeF/VLCaxozbjzridXOXogTaXyj
k9cvLx+w/yflR4oAenM8DcIX/pVN6czfV5igo5UCZLRXDhqMmk5p+uS/cIfeY6ri
tAN7BCigN4xsD4DDUjbPgTRNGyAA2nIk8UksgXZ0X+vy+UXn0GpauKoH44ohhftC
wQ/2W6J2EZOCDf+VurcEDU/VXkzNyQe17KhHkfuwzWkUt+4zKp/AKCc3Ajq3aAaM
ylLHs5/KeUhbDnllllyfGHVpXIPgWJkFBcc0ylz4PcSRnkg6wMxuG+Fiy8h2QWE6
HEK2QJaFFloS9Wg3rsIIremUgmXGaKeGJmQ7Mc98dkS4tXSeM9s3M6xIM0a43aa9
8PPeyBsXU4s3WPjKYHUlT7cHdBr/k0pbW3w69+f7JWnHOKCeE0SL0Lpgwi7QkZzb
SOad7PD9zpJ/5uvvJiLym5D67DG8BXViZy70Mfs11jkZ9INUnbX+hvYDwb66T/2U
D1TiOBGK4Pw8N1+gl3SBUKOpxKvg16dzEXIvN3tEXP+gtjzj21wm/OoGorlqZYXh
4S2fguPglZXmtchpz3TRazr6+yHd0XlXqyuyeiAFPNCtBhH9/NKBuG31Z2pXaDlU
hKrYFg57Q1PS//BzTuSbVReku226OHf6YI20J3q6iNepy/IVnWDp9NDZenIS0glm
gSlT06HeCVP+KtmqOdb6BoDf0iCSoqqdGYhfd+Q26Y/57Wi/Aqk1rWb29NGXd3S0
5/qTebqgPr9HoZONZyWwRRdfdPdSO9eekYLcgJkKfCVdGN569E0u265aNkWR/08I
cuCzWax/EnmBnWDyqpmlJwu4ZcmX1VWR4MDMgm5p6tgXuDsK5TZ9jFDojjuy4Xq5
pw/C1k3Gb08aLyVxdJIeOHx+lUgOGQZG8zr+nWD26haGTnYLs7muwwuTJgl7lAEE
m09M4QIGuu3txVQSl8aYP2kiHW5DFODakQSq5Pw70grlZ1DKX9bfuKWE7BAoFCC1
alHPxMM5/awifDtSlLicf9NGiYLTACBmlvEO7A5G6wpQLWl/tnQia6w/+S61bSLS
L23uoOocnhaMXRFt+tyXX0tHsTr92aD5QqJPnv/posT1jOjDuMQM91tXQDTCamy4
R0Q5t/rWL5EuZIJHkXkLwyAeLYT4qXs35EK46IJpdOX7FOitzfggJFRCZN3UKQOI
JWsDtNabCPgMysinsXd7yP3Hu2ANtdEBbIX1e4xaZKJ5Dq9Ocb3hIv2hM1+TlafT
QfiFO9XLbQBf6gIZIfuPocdZkXQykcwdDeRWGDoisRHztXLFH95KTfDcdTT5Jlxc
oFj64jtbSt0lk0blwP+mSVOYnmFtRE4nUTjEEoPYn7/Kq8f0CZJkeSc6Db7O8s2d
CG0W7cJSdfn/Ivmtp6e6BvogRtoiulRWr5hFonM2InBhupDSMYFfnAUcDtTddV4F
/rPqVlDke8diWMx4JUyJyEet3X6asTXmKRg3qAlK3nl4l7zUl0P/vID0hFTGZ3Kd
e/vjAgQtyVaKozYXHmq3nzRlg8XuXpQXcKrPJVbVLB9jfjWirwFA4/ZJnmS4/wGj
hPvIZ4E//S6jt9k+bV+xtZk0YPpaEovQ1pimzrLmCtkAETr7Z2qV3M2+A6vVfPNL
ZbIX+eG10M5Kp9sb+AlI8Tl2dn8+CGwHWm2vzb151uA=
`protect END_PROTECTED
