`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D576LBSi7sVQVrDK0s7Z2h+DU4V2hOAfQP10LHDZg/VDh6aTIB2XNpBOBH5d4eQ2
Yk1gDrWeffoJ32jB2WKP5bouZM6sU+6G7fsHFRR8VawZZk5DZVpJ4rI0N7LdzU5g
h1jmTMtpuwds2TA/YqHoD1sTyfj/2siG2KS9Obxd0eFDVDYnxFp/iwuuh77JpeRN
l0AaYLuomo5YXA1SaCo8oFKNFSxgLGiNPrPIVNTR/CmgiOS1Woq6AWnu1cXK4yM5
drEcQXpSocYn7frgR+YGZJbuX9rbdV/G9uSSDGXhklRDEAPmNyPr9/zNvB5kJ05s
SU6ZJK4YxJItwtWQ0TFQqaX8G0VkEDWgYa6p8qvcrUs6sEyvk2MMqS1dFqEP1xea
cIRvHkRrNH3QVFFEosGuWCFhvUlSgCcyaebMtM+HsXZIg99dg4GAl4vvgIYvmH2H
PVozJ/WWRa7UlhDI/OHnFLDyTE2Kkk76csTtQQWfZi4Di7b70J4hyVGJYIFjReDR
uL5FMvdrEgDVPKPyeOI6nw==
`protect END_PROTECTED
