`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8x/3ZAd4jKfWwRpvRRnRLE2Yu867/XIhTeCNDCFuDEhmtp6YyomC/2nicrUOWSWw
4JVuTVgcVyXMmYEX5ltKzHl4NDjozKaqe6/lLVl6lReWFcHWBNZffn2azWgJm/y0
5WwwDTdxE8WMh4Af9dJh9tPtihrUtec5WVpTBl6N+IvJ7nZ9PUAPK8FVXuBbRnkk
Itl4Xei1VpjIKUlVx8/GE+utnNY2af4BqDqYb01S9BwWWASIptuy8PgDb2Sn4TLb
6cibLvStq5D/omm7Hs5wLtRINCt8P1n+Ds9sAqQSyb0GGucrsOIJNek+7gTSeHMK
JlLEJF49XziizsJ4SsX0GuA11ajzNaYjGVNzYB8X1xpK8YsFb3x0LE3LzAzEb5rh
9JfKfDw5pD9uRE2Q8AKa8pPVvI7Y3xVKwESFtVFNyD4pRTzBufFrehUIZ/gtKcQV
tZsceIXCxlI2SQ3LOjKwQAhMy3EVfpbtV6fITmc9QRv3J/ueh1lQ7Q0QPkviMuEY
dAhGPGXNm3m90ORWMOP6gg9meM2IzKwRo7qD+sKYf/U+vb7WpG8Ite2n8k6hp9sN
/blp+u3or2I7iEqqcWsZ6nYoOAXN5uiohMPFY2zB2UflwdC7XjLmmwgLLUqnh5Jb
7kypMgOzzc+vP6Wtasyb36LkkxJOLhgrIMrjdJB/TutkH7dQaGefGVjKdO1WYolb
VYpKVZGweNNgKeqioXLMkMXpqdVR1FYBvYTq1HpDqNwr32Ze3/ROpQoHyrTwoaWl
`protect END_PROTECTED
