`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
udQYT4qfPQPW0aCZ2PKJMh82XWCYrrJbq3E/TvoggRAnaVf63ROe5pBiBkh+OAaE
OsAg4HrioK3It8k5dnirqgZJexpAey2paECBdFibXZllo6SA2WklIST8lbeNubWI
VDFQUU2LSrYYKjsYZUf3QLO4a2w5eyseAHjzCgLxPvPOuhBqCwNBketODWMbahiX
OjRM9XKwTWM9unbxTPBgW6/rXHt0lxrnSzv+o6mErKpBjSloAcaTsJ7reMrMcwYO
cUXF3rjs9lrpkE0CuS1aRUrmjTRJeG12BlQzKiSkvoENE7c4gtmtD5Vw8ATdznYY
zXTmKECYTWN1RFABP3wdf7FacnrakcpUlArHj3RTVzoFWyEcOF2CSvociA8U38ZN
zRn/uJLuxNpvCPtnndU6rSCTklX5+e3zTQWAiAIkrj92GCyzvMZDDZomcCyvuHgM
XNdIQRSNnwwiOZcHPM/QxPhiJDcT2i8qKyt3IV2RH+c=
`protect END_PROTECTED
