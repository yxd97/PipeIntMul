`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
off/ACYEAIhYCNX1wk0ihfeJN0IbgS0SVzlOL1AJBmhLM/8FeXJw0+45eiMHHZqX
hW+gHDCgKLklXEuNb9XwvXQNS4bRn9U4PoDqfY/1zmLqu95AHGlq5PUGjStMkXsN
v3DdfLxZkazL8W5BwXzumSX/G8P5lmbaddTR8fD6aPTocE2lDkWECGNPq6Rgzatc
TaA3Ul/NPyF6B32qdn60cM2OvafwHUON9isxkEJteEoowT5bfmXdwS/cJodR7if2
nVPRKKEYRxH5dVWCI4PfkjgUfofeRlaSzABc6fzoBA/6XNiR+UqowSBpsnIVm+Rg
jGrNZgi/+0dn6b1adQzNtOg10bJvM+xnDIqeuqwNdy9LaMeUOTWAp41wFlSTDS/e
caUF4CGUULR+6IIb3Lhm8aWa1moB5vrmZ+fTMF9dNRVjQ3Hifu6acwTgYgckF6bs
`protect END_PROTECTED
