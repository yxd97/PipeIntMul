`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yb6jR9p0gURQGtTOYJh04dlhj4Nlf3ISod51Tm/69XSz1VA5suKtsGUdC8k6eU9X
lS59wQS4F0Cn4xfsNDn1ejc4PWKDn8RAc28uOb+iunzno58Rm14CgO+SsWy8ETby
z+ybJ5/OTJ8SCsYe3MNMXjFG9gNfL1IoGMT6PQC2Ho2Tc1EN/OxEY9oW4Dq9NBPa
PaOvdmqILt5Nw66Y8NdHu0/u8tMJAUKvFS2Z14gpEaE6J+XzywHLK4Fhm2z5bCt8
ZTedQQVVrkUZKYhMF5I67Byw761WlAismGLiYydcclU1Q6FkgZJomDK5zzelJS6z
`protect END_PROTECTED
