`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xk6NnfEEmelKsMBluiya65BBhxV9anK5ZU16wjvSTx0ONU/LMEJTE4kr9O9urctF
IItOaM4AH9g6p1ZJjPkqmnqPG40p5+0rvfE11HWAHIlWt0DR6/KHAdHTqzvua6rs
UfoUe2X8OKPy15s44ULCh/lgg3KqvGuZd6vhyJ5vLqDU+KpOlojhE4RfeiH5G2tY
Ao+5AGt6dBYddjrmP+k41Mp5+cA72MW2kLDXhfUx/t2qgTi8yOcaJf2eIsaDSoVm
SRSlNPvkHKyjp5bsHR6lrnlkhIsu5KQqzULTia/lReWkQNTCM8EGH3sGoxPnPFgr
A++jsE9N5IcqQ8JxxTA1QsdhW9DzhZ0LeofZmA3If6zcH30v3xLStgWsQ+fl/dNe
xw3beCzI0gQuBB/7oYisthTh7CEtJKCuCvfCcgeVVch9xiJ+MpSHs4w0NQKPMUrh
l2AW6Ztf0CY4jZuTU/EvMtn/0ZXQV1VcjA/2eLFbXEkFBvE8gZoG24IgXV+PO11j
koIY+9iQtDJCoLmxFIiPxuJe03VRc6RHmEmckarCnxA41no7P+YqT7kaojcv/XSQ
XJkIvuSOqJiS/4W9LTJdetsV7x4LH8FYRh+BLAKsWh1CeMdUurlfXpccj4iIH8yV
waoZtG9mSXpT9FcqYODTjJZDgjP+gS8fSpJNEgmAfQa6WySuykvaafQOqViyoCaX
iII4cdfyxyMzGI6hYMx9PHgydvlf8RIA0/KfmmlxdSfPWrUnfKv7G4M+4jabMfwI
63naPFGvH+BB59unt6gQ9fAg5rTP5Riflg1crj92kUzbwf0/2qQYTQ6HVAY5gjEo
R+dgleK/g6N95qMMKAGVsAaGzpc5znzhPRtRLjAv/Yb/0EPo7rSOmVRzBKhaYckt
NtE5PpC5sDSHAdnTGsHBYuwME3rvNnIYrGyMeQomBcU=
`protect END_PROTECTED
