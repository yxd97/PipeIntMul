`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XP9109Nvc1pzo632khILEKstt2sjg7EBJeK08EQuQG1pv+Jk7fLdLQgXLbExsQVc
LkhYquPwTV5q63Ezzcyd4n6yFG8duEuLjz9VXPPByjW9l7wExvikNO7NTXTKrooI
NQAK0ldkoHZ4MPCYGUH/dSSpbZeHs2yvTyA17uNcDFfO89Py8CFGImUFDwstg75m
c4dGIIB3eLnua8wGlgba+L7z6IHcF0IMRMgql9867XLP0c1dd3GA8v2GXHkm05vA
QsPvYczJoSd89R3Rqu21wTtAG+FCHhkY4YKmDrDquAHAbC7JtkHzM6VLW8Pp70D9
R55PLl0Iv+FtBM8h/v1+6LYf5Cjf+nVpsLJHJIzq5MKjfsNci/bZLQcy2fUcPIxY
A5M+wR9yqMCTmLHfeAmD3IKQCVtIiIc02HUlhR4hWoF+5rj48fC/06y7XqQ1UXvx
NqkB8TAPldfWUAEtRQh7bOoxObASFDm8NcEt7ohk4m292fs/HaHogI5/9L4oXiXZ
lk+UVg+r2SHKC/BIeCJi1Pqo3meeuwkNbuO5lUCGVdXVGZ7DUks7v4+WIBaX9VRo
ssgd4fsuZ12N8dRaU//qrA==
`protect END_PROTECTED
