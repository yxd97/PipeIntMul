`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/MexTvrxZHYr+6GnsDY/j4rRkbmGEt4MwVkrVc2KHi8P1lz72U4/nXjTk8RMlq2L
XEYyUwHVLOdLadfPdKD587iV3rChWbQUFfwBMSIFX8YhNEcTwVaO7eRRPPRSyaS0
b/cwWghVplka22KqqJm5XZ22p2mj0kwJF0/ADu5fjy/+xGQvqwRpt0A0mlCsixzg
7TkFgRQEytM1Y4lJTFbwbmb6WVDC28NmEeGGJoUU4NIorkzjQ3lvF1tsAkyGWUaf
loSk/FusqRsjSMnl1RVDtQ/ozn5KKpNsHAa4Q2GVg9mK8lwJI91SSE4UcCkIgH1O
O6ObsvDvX0vY3apR2V0imUNrOVdAuWCrgY8fSnxuXl1mEaacC7uBxH4+XfByITI5
QJBT4AlEjdF7wfrwN7uGffYHyWLgCHBSR6WU2iccOPVP9tHrDDu5WCRgZc5N42r1
luObLqpJAk07T2BPXH/bx7LHrbMmqwDcyOJtW3jipw4rJnJn5OkcuAbWLUqT3fYd
7dGxqMptVsz+7jn/4kYVygZ+qTtStT25leZ4MZHB7cFO6rz7RIdsAD2jZAVfrQUH
QTI+YR50TuH6s+C63uNjcTqaDNcPjvuxA8PQCroowWswKmHTkERzbkFUSFUX1jfk
P81J1zGavuTUDvrnd9aJ6gwb5Lul2DjwUaMyrjgiYi34pHH09Q2419e2bLpJcDU0
Sb9pfHiFyO2jFJoL7n1R5uxCn5y555gOJa6U1TLc/aeFG4O2lvNvZcjyh7Wzj1xX
d9MkWMjixcojDm/MKAcJopiNLACgNMC5jgNhQycNcQjTIHvpdkM+EkrNbjQcC8u0
IV7gwiiItMHuWOZR7Y6BjkNz74uAX1C2I6uMyEpFM70doOp6a1IJN2M6teDQOwdS
sw85/ZqH1YcPUt1I3KSj4F5G8V/tGmH4Lzh7NSea8GAwupn8uFa/zZClrADgJfjw
P0E4R2J9Q82R9OLuYvNx35Q3My6jjY/J/cYCQwOXB5g/9rCPbvPMK0Sru5oE4qYr
JBfq1vjjqDvlfwr3tvO6zsFpZMToudEAT42/AGvlvN/LFxoSjaVjhRxWc7CYL/VH
10b+LLc0hvVZByDynsdbsGKNvQA1GXwFjVlolLszXYnhnhYYRVPD7HE3vfbWnsQt
l9Lu2S5skIePCed4BfqgY76avq7JyG8/OkiQtNLmYZwieYYBJjYaxPLvP961LvU2
rEcmTjUHdokcB8gYGNGUPtYH41maV3/Toz4BuEWI7QucZU3IWDHdLnt80rxWTLRE
3MuPQYhcblf1J+wTlmJCwylRA5iWHShCVxU9YOutwsp4o1OQy6nfJ3jQcPafMTC4
qpukqCp0NI/Gk8I1VvLar0/HiehiDTYzD6w6cwapooAPpgHCWExQoPzUkQbKyWjf
uWE5YtnSb5kfSmnqmpu/uEZxGs89JL3gTc1Q5+Fr9SnFjnJALA8qGds2UGP/UwNX
IgRsZMNNujFQqIUyDPzLKnYJnKQ6tq151PZcdi93uCRx1OpQ8m6I4flhFGA8ae0z
Ux8AWGb3impQNJ1vxfAGMzZ84GaH65LunbUdhLb9lT+goXZDEoL0PruG74cYuGWP
gJAAXqM3a4el2aWCQCXZmni3BKEislEEkCkKCmgAp8eByUgXqOnHe3lZIDKLQgt7
bXlCWLEPGb8uDmAPBueVqLI/vBWetwmI+R/TTEMKC1udPh+dl2QdfZQ8yDCAyDqU
FYpFKMerGdiMY77mRZe+HYZ2e7+GE79TJhG3qxXtnrvtKBqOSmlbOy8M9bKXRaow
iykfxBWjjcdJwbMvnnWNeC3a/st0SLd5yn8dO+lJ6ZEQ6n1t05V65Zeo+ObzEkJA
rm4Dpe9FNvMMLl5znyN9qki2mbchjg5xfcg9QgN9F+pO7Iry1hsbsXsU5zRfdMlh
gt5qbBqWuxYd2oSpWdLUW6Pz6dBQ7KK7CKLY7R1dwY4EQvEddieZicAEv+9ZtXn9
j+AwkrYSfI2KtUopPu1p6Hb9+1rR2DnAuPmw3wvU9FSINb6qnwtI0q1sDJNbKPCY
q0546iAe/cQmTCRqrcIYa1+meioOHRsyE34J0UQq+AmY657Q4yhj8MoLTDo777QX
HuvPR4AosdprSgeLpaCA+dED1m0aYM6Lsd8iNPDO4cpK1ZaFvjUDMjWCpAt1JEGn
Vk0Zf4/WALnQ6zXvuKXK07wRUl9wSgZea/lz/FMEKQ4vmTimfrXe2RoH0DM2e0/r
eSNFV32WY0W734Hu9bZY10tJTbEOOnSTxauO/eiK/uNUrWNxWCW8mVj71cz8tyU2
l8KEaGB+ktDa3v22w16Q5Foa8WAnP3LySybPQWk1PuqhLrhOMhyFRuIaNsLY7vbS
zIxk4jsuV28zQs73NI8+MebkHN3saxcA0Ypgwq0pGttMV+dV02C4tgR3ac8SbfR5
d3s0BUWEv0eblmT8m/mXB8E/epOPNEaznEN8lZ3tPfqTZoDwK62YbAttSLivbQAZ
pfvN5sCQyHWdtZIYqpnae7n6avrsFQSrxyddpmLEPfl0CSjSnk+zotThtOrlEn3K
AWs1+xNQrZJsw2s33H/Ef8Ox1lH9H0Tgy0JhlI6DYtmmt3Uvl4izr8djxSZJttSc
w+qQX3WBe25nfLahoVij5kZf085mitTAfGr0OKbxx/dKZ2KVjCxJq21M/E20PP51
8uwu9MqsAyKNWtXdyqauRsz1YScZA/VL3rC79djuryZRdyx4BqGjShrMPYEPM6xT
IFcO545MB+Y0a59t7dT1WrqIODfnvKYEsyIwK2vGXo2+UCWtmAajsv7kzO+z0Q1f
JWUe48m/+m9pgl1OKKlBRRJYb9v3bMjKBHMp5LLOu47OYrabZkbgEQ7AyqNYGTsG
OVxW9CbK7YRfZmzMakvz2M5K9hL8yD0raL6rRqTtXShUnJNHhsRcwDmq6hmkvJ6A
ABLItj7P0wfx0VRIESgn4kY+S1VZHue1wHklfAIRFZK7NDMui5BFIgNnttkh2+S/
LpJo9dxgS/YloL5aaFHdZXldqmJ8v6VBeb2Bjo3POy7bDDAXX+rBBt8nI02f3H6F
VNPRp1wRVfk+xMLKmlR8XlYzq+4g5/mYDmtE4GjGCVHTaL88Ft7tvKh7QW2vvGyR
QICWq/4mAdrNFohqPuJzMPhgfS98pVVfmjUSibVvUKmZG0fD++sg/kG995WaF7Ux
z1b9LqUUT1iBuShp6APGskcJMLmgXSRhJ8rPwYFDm46jfVgJkLv2S81XV/3krWsi
tuXryexTmL9wn8lUmZ3BkNBrrQ+VTST13/YGeJRSgTFNAOsAbuBXWpmi224H+j8g
fQTc/lhoMVBKp1x+CU/KRzgeOpwEzsMXUIJ8FhlCRcXdrPOoSaLQCOctsYM6xvj9
2FXonfExSkh/SZx9moZ5ZTiT/oKWTdsc7adH0gQxzuATSDYbrgDAH3sBZktqniPR
gbQQofZzEw6lVvpnchAeXUMXCZ7Do2RN2r1FhogcjDjWFFaur3AY3yYnIAlyR/e2
FJ0RXxUcXPaTxq0rC/9HF80866bEmHjIwBiqp3W3WqN1cXXUUv8afh4Xtj7MLd/u
K6o30ICacTVMFoczvg0G+oyGKyt5HvbPqGVO+U0S71TwXwTBlnTHPR6uY32M95Mx
4VPS6MPBWEAZt447V8g/G4GjPhxj6BQh6g7hhfV7r4jclkzX71FHCOFyqPura62P
Q6YH6CLDmr2A/gTGABmvgNGODoj8sDoBaR0XuIQtFYtJfXPKCQgkzv5bCBSt5BSK
G4jwOpZqDcGhqzYpVnoOLV8tF7u0hHHYR7fP8iHKNJnebVdKHlJoZXA2pN+DVXOe
M60seaiVeV6Iy70JmTqfOweU5aJED/15gkdTOVcXZ9x1wWEX+k/U39lvFnNUJsYI
7V3mllUHsJ/u/gsWT0AT61rymTY2IBa4AvCaVTjANYcyREesIcpKcRhmH2LI36qJ
mOao0iF9KW0Ov/IijGOGIlVqfvMkawrUd1ICoLJz7IHBxJdt1TIqcrUgV6AS+Rlf
uYdo7VtAKeGF7tj1pEZox2PGNeWooN+A4awB4SHApW5ggVPRPAy8Zwm1Y8jMDXYg
WKub09SLt23wlHPrOo3cYzkH40G3e7mAP6yw3Tn5ZfLrzYG1tS2LhkhSuHCQQvDA
tNK5ku8nPyEmcgdcjz5VqJztzlpf0qpbG/fdm7bsRnw2RgYxy5gaPH52Kr8t1IZe
tt9VLRjg0wMdH3NoSmBAn7GTR4eCpaveHkn7P4h+VN010CgefjxWopqqyqx15azD
yniqqEjJ8b7bR+Gk8SAvGokmrQH2xZ9/HwDAbSJ9hvZ2MrIEiTYwnnYCWAVClWHK
PLsY8rpUTvrBoOW3vP/xlFkPUc3QCvzRF/0zXZy92S3FtYAgXeBBOwDN+OP55zSS
jZGxWDng1oqG3PUdDQ59z1/q1G4jjlxm+HmlwTaYLgeVioQ8Ikx0YQiG1Zi84TK2
LF+neP65NLC72E3tJ+ld3OgIu5227rkbO24SJSHGISRfZ4BKdpvOCQG/opZBxZ5M
khpUJfMBnk/udOM0TG4PaEnDKnJMKVn83zXsV4Rjtq1tVUNpE68hyzjiYZipegf0
kOpUuCC3mSeMpExOg71PnbaOH5CzLEdYlOXn1tsLcmvOo+wQ1nFBOg1gztqmhFnP
jEfxjankLe4Ihafncr8AAO/xQTjYOYAPaePUWCXokS6JcXimMBYaVDnDgrVbd1iu
LGc/vjKs+kt7c9fYc3qvpnpzJqEwMySJCAJNYTIiNMjyLtX6zeTr/dKCWCelbNbw
MwcQOzVbhuzXF2daek+XRapUkS3HwNbZsSZvlgeVCEkpq69owqLPq8pLF6+KEh7+
Rn/4ui5aY7K6NXnwoE1g26QK8g43ivWSXsdupgCpbsjX6oYvRIbk5TPMk+0FJdcn
0BGtQH7dWkjuQLwDnHTlJYwT6AIOqbzkDyJLEUneZBAhlixG2T1esqzuiERs8eWt
bh+hFjZeLBKZhtqcTaejyyDwcxYqfdMzH11ibtzXfJc5rx3u3mEKVQoCqdliIl89
dltIQY7vn1cbl8nSSfF+ALuCUCWMg+0ZFIRd8XvVeXVkXBaja67PjFhHXjZYnXC/
ysk0noTZZDGthIxapg7L5mebAav9D8HrP9Laq4ouE6q566VrQ4mi9lhGGQDRk/Sz
/2Ivv2ozFh5JOvogueD4N55iB0V/jHdb+TkPlUV+6tLo4vJCqs2rca/Acv5xlG3x
okqzIAaN4RRwmBRJOYpCHKNuLMSPVwkJ7fr/IQzDoajJAuEa8wHMraZES94SSARP
ykm3y3WkGdv/29Dwf/jvUSiacNUA5w4ksRYrNJEQ5+4KDdn/RC9otQVsvkCMakGE
eLjqRPT9gncx8oWvF6un/k7OVXg4pPmBWKr8dEC0ZRZGM4aTJiKMwp12o7T8Bj6G
pUWaJOYBkzV/9ik0KxGT9dEIsZZhXj+d32OGTpbOx2KzvlcUqJgiGI9RTe6XQ1L6
TVonJ9Ykl9Dm9t3S53kW785bri5XJEfPoJJLmpuKEV1fR8xYqsMiKXxgCo4ky3zI
azL4dP6ljfa3ajYhWrmgrRu0jaiBQxYDI0EU01fO9MlrHvQbqvvAjh8b0c5rpLjF
+3hU7Exxcs8kSbJRbpCZR0tves/zuFRAVsv/+sIZbihJQ/mrE64bEcbxYJUHqM3S
7RAkl5cxHrNHR863jsydLtpUpmYMlpNXNRd/Yv2BaS230N7L4LDQs2TccMYDxHZB
3VSiBCRvfyJHfGrGcE9mXntDNDJIZaThiM+zAN8bILDB8XecpQ2VdNW8/YnT1GvM
9WqCw+TN3Vl9o1fFkrCdWp8cjZLYd1c4ZTclT4uyFPwTr6bJkEr47d+a/m785SoP
yMzNwiYSNV2RNbSuyJmW+BigNfIeHlX8U0rleQDEOsCz1fHRhEYXn/8b1+/M7AvT
9gkmpGEq80LX4JiHAvE7bj9i7FyDxlM7DLnPiBPLUNsA0fmVxSJDpKURSjlwPINW
0nCrlnx49GaQ3woMWC5Xqs/lBgD+xTy6DdF/AMOaDNUFjSSJXu6pLdA4uXAQqj15
Ppi08dsqLgUoI0xPh/aeXpywOgeJqDkGh/Psltkmty7kGIJQfuZGADKjuVbJr6MQ
MKUzCxVlKovJpQaTaUK5FQzCvVnnMzSB2L0oE9QGGSo3gOWddSd47Uyt/ZScyYUo
jNvsUXwrWUa8ocyagwnZcW4kE1Eoh/aMr7sNmbqrk93GaZf/HG2IJ649uE2vvyvc
Q3GyZZqCAo05QD6rnNd7Iz8LAKW5jmq182pn4LbZFysmxGA2oWcY8AyIjfhfJuyu
KPglE/LOGDOrvJFvPB4bOCsQtWsg8qLTspkFIVATlY8onkkiyU/FVl76QPFowYQt
yxykkvhDsFPG4AESOnODLXaGQHdcZa8zT303IzdA/zM+98eeqy0jIuEyZREjUsx2
aSG3yXLqgaK/xpGoZVleAenhWMJ4Jy4TQF+Fvgu/m6a8qzp6Eir+EcZzhNuQwVz+
Wj68vCKGT197kpYuomGY2tff1nXl4Q3Y+u36thCiWF5PYKbPdZgbLLeWobaLigx3
Ra6xZZsav8O6iCz/RbdCTxVCiP0PtoOYlRZRG3A6AZCBiLvwxgMhaMEf1it7/QMb
e2qEwYVLrq5CjKeSD9TxhHG7S4UhU3zK6TdH1STdaDVATsMX1qenic9jNuelHA3q
/58xMZCTU1LEKOA5zzfKDdQdhKTmK8pdWcKt2T7w3lnTl0ZdOmJ3fiD6hCDLQDcX
hB4oARsgSO54uTravdUiTeXkO+vMx7ZPm5fLzMbvj7anRhAXZFgwhc+Ba3HqRSj9
oFT0JBBV4OjII7dljbjo3EI6Ri/0vNutjnpHHNU3viPTt8skSBoA8lkPhLt2Xrcg
8e9x794IGKOTdIasHemuSmyiSNmWZ+b84BBtiA87UcGdjduFFebZEIZdz/B3KPD8
/7/uprb/6V9d8OQBZtTGZSCFoTFlULWuVBKe4E2iTVqtzHw0342BMtnZub8pWORt
a5bLlSF3+wmt4c7MVGPWoTcbGhdwJvmes2kOZlUtZAyxipreFXLolXCojtbatWzC
MIEXv3gO3rr9rA7BL7QtVRw6Y/pBjtk15AgfAqaLPfy5VODm1ln4WoH2qSIUBPse
EeFXc38dbzXyqRFyOj8vCTa+6i5U2JAokg333hpvFIg0fVhpwViitIxe82cAYR+T
/8rW7V6/gwV8qWuvoTvLBCsE9r+7xuiawPlNN2IFXm25cNlZhcSB4Qcf2MP1LNgo
Ys0ob9gBnoKzxURzB+MB5tqxW3VCXHswv4deg4G0ZGryMFsVy3VaLqi7l4AQGr1a
WmNW47E4fr91JLsEbkNova2FBA+Vi1sNXkwTfq0a0yc+17y0ve2aTSadq5QbvY74
vwsSYJJKX1cbvSirgWyjPSeKW28D7oLoDD8aGPBXl64jJ7GfMxGQ5R3juRsIlhhe
dPGMoJABi0yrW3VBFEGcy0rM7Lq1MPmv5M261/xf/0UjK1bSurRh9xJ/2LbSGnDz
glq662xySGmNR+b/oX9fiWaZFCDgz0c4xpehuIy1kfNyQcCWLkaiSwVQWtEFpVnP
k3GC7KsK4CU5JvhDN2uJ87eIVD6jzU4umWfW5h7nou37c8iQA9m8ZAD+EgAwuyUT
BUaZr6d9OJmEceLj6UcpPWhnDhFunnjHdjassKwR94riVomH6Z2n89y0R4SOCEQQ
Gme9yqCAwRLQI3R7ylRe19yG3CZWO21Gt3lJs2EybXyIsfeFOC0tHSnw971ydr2f
4Ol2xfe2WMnWxG1MXBMxp+6ZLaBc1WRbsr9NxnVeZys05M17y76pRwqtENRCGvNu
NAnUrVjmFRR3OT7kuNYAncG3ndlKRBzJtQcIUYSIsq5dABRY56HCOvJaJkiNp99T
Zwr8qJ5vUwXkeAzUAiINbd/+UG1rWvT5NtcDzL/bxB68R9aS8wslFxeZZIO0emJM
JR2mRGJfUD+17LOIgDnPtzNHIg/dpw1cO2QqsXhsY/V0v5XM4+nxXcBnFWYCZBY0
LJtdUr8yKjQpujgX8e9RxmqLLWCmLH8I9pXjs9IPqdP1rgxOIjbT50xBkXY1yAo8
stp7jESmhHzMs9SNvxY/o0YfS2L0ofx2Bgppif4auKhKaSThjK8R3T3bMhEy6wxM
WTALK2tZ0SCwOyFAcg0hMqJEix72fi96li9TJAfjYj7aLyO1k3UTx0ZcsHoF0JqG
OjZY4F9Ka4itnxtpxZvnyoCKV9+UOvmfH/sj0eDwYwCmh6bUXddYfiYjTB04vgcB
V9qhr9ITmGpHhma/B8moiFRWlznnAh8z9ts/Gc+g9FdvO/eF9UJEpSSz/Jqa5qYz
FshHP7LFcL0GNLKt83FSScTA6daJVWB0MJKVTGSyBjuh8jhFyBMWWrCERmfKUW5G
mhf4iRRYuULd1YoVf8MY2NNBJj8CG9HCch4jn3AvlJUI1ITR7w2GQlF88hM55kQm
bpgKg7rip6QqTczL0MRxUWKhGW+dvNXcwZ7dUn+Ad5zub/2syBQ+Pb30QlcH6S9e
+4SncjF2FOt9Z11eZTNGkZe/qqMoL8cYHCrLGilqHbwKXpHyX9wUB06yhLfz1R5I
c521K46muPayzG3ei5fp3OA6VQ7OMQWP9wgk+B07TwBxAvaYsrFIO/wNauRvjeuY
ioTC5XdnboDv5WT0saTDzcZ6Led6YffId9+UdWIP8YK5hZIKmAQKvw/mVxV6CPwp
lUF17M+DCWi6EEcY5z0VukYmdx9/2x1DqplN+OKoD0h1xFdDj/3/l72yfP8J/Pv/
+QnXTzBbqOU23b3gg6cvb62O2XZgHl771PDK+1RQmwAwiEApkurkUou9egvsxJzW
cWmZqaq8Lh1beShwYnpEQWoabB75Xv33dNSBCys7vS/Aj1dVTIeLlXM9vjQXP7zE
G+NbT8v9CFhgpBuir6hF8tQ8DRRc/KGacF1XYW4emYJEKlFJYGPp3vUUquXmQoIv
q27NULPiLilBpcryzKWmrcQdjLZGnNZLZzni7JCOdy81pZT6usWhwbekzxReJy36
QexMotEWEGX46PaejwUrpiuzz+kN7kjM4p8+7YRhLq4xl8EE7YrBo2XpmDclOAYh
il2f6UWENPH8KibitGKzyqsIqT/zeQV1HA84y44iu6MH4jL3cz0OIHSPipLwOxAg
5UbNEV+8dwRJzPd7Ef/Hk3LJ13Bek/+ll+76uJxiLlVKTL1GK7vPxMgoFqkIfZtE
K2pHsiRbQF5prqKuXFTz7xnrQnbUnAN269Jo9nnyiac/G41kl7BcS0vod65ILhKk
fnhEbl0BIOeeLTcQzQ+TkuSeme9zMAH5UrRhWr+lyaMRf0GXjbn+wy3i2lW1rnmM
igu54MOWkMAkra4JqPSF9hLzEdCMjAmUz/6xvOBGOEbHKnU5cQfAoISBJ3eI1aFA
RmwzW8XiV1dRYvqxPG2Sel5kCHKD/l2a8uJMCK7tx4Q9A+GZRXVj2XvyT8JKDmUg
ohDeIjhm6V4Nuz07CewGirHcJumq3qx8LRLO+gz9D/Oy7lf6ikmNMcwF6YXNSCDV
iwcSXjd3GgfjssznYtx9sQ2Igk9/OenOr3XCmZ9BrSG7piBK6f3XEAYw3O/mokfx
yGF8vLQLkgibqyxF2p4tiXXMpl6JFs+CEOmltLApUsSvvFUiWPgOUYCCXaWlp5zx
l1G9SlbjY5uoa00Cuo6dxkQf9YXn5+UZlLszv3Szsn3lBxgctmPv8PMca+u/ofpn
GLecc32MZs/Nr+oXpzUFL8ri7Rp1zJd0JskDAr492su3YFUiSVrsAywFBzaovpoI
oiYquD8JWSqhidteAyYYivtdDmrx0g7wuIJ/o5Ul/BwM9TIxa6ONbIAkvgimId/i
vIb8zlsXepM3uNfJblbsDcSV87g/n0hERVlh7SDQ8+R6b5ncm5212CpmLqXs2671
YIGOfve5AnVItdmfYw2wV++hRVsGhBiTqYUPP/jjbtGEkEYkMjCMmjxNmPYNbnyO
dwZIqahmI8mS91NO8cwMukWA4/rgdWCtRGVRzzDJgOOjl7+1oDRRoBDggh+wm1p9
6MatnzjT58RHLMVdnZfpwgjPecKue3bxZ9udupOXARaw1ViGJWB+Ax//XHcxMJ4J
nxqsZKR6fJs3FvRUNKy6yJxR+GYP9DdER08KF2zVixIBuleQBDknuNktVhV2gd/I
RDlBMD+eAgA3W3GntjitnEHAPKXsOA1SIHTMg4mtXirhpNR2uLb7aQCTlaCepDuG
`protect END_PROTECTED
