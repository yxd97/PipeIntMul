`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6gIAmI2rx3hgx2+B9BZfIp3IVet2ZcEueFdV/SRV66Pd796DLVBdOeRsv1ZIQPaX
1JU+C98+GGALWCJ1yJFSyD3yZolgry/fJoTAltBsGXP1m51igpzxQerwABhT/fZs
XB/GYQPPo5rphTDCcRcnB+uF6+ZH8hm2tz/Fr5uTWwhR1baT3WJ4jaiGOuzhOyX+
hnXpPvSe063ekHO4oeve7yZ3GPMiNwVW7c5+3B/Y619VObUZY9UlFkqz/7gklrFw
ey40wmlxbZhsjAv/xzfzpov25lHNAUn1GF3uKpxlvN7TbeCAu+mww5XKzAHl3D28
AWpaRdiMIL1+7XFi/cRzpYx0bN23N0ygCKP+M1YJtIQBfCFH0NOojWxY7St1mLWV
/qaHKrcJMBZcvry8TVAwhw==
`protect END_PROTECTED
