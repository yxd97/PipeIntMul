`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ON9qd0L13OCTPxB03LjTjiP2UqpVDWvJvYOlww/6gzDA5atfTSA2OkpSsc+W86VD
GViiKadXuznpHk4Du42esENlpJg5sQTKUQz+N4Kv+Qro3RheVoD2HGbQsqGrZs97
+dRb5cpv3xJ86o8UYrcv3Lsp7NUkDJGjQPTuFyFhLZLipYHrjhbtg3Kr1YijywsU
1p+G16U7oegwK6wwyJuHiADapPEeMeKTj/5Ecd8jlilWSbi0GmguZuRrHAPIcw5Y
Czh1FMgLhlcJKi3zCAlP9eaTl6C6Z3tpBxsgrVXMr4RzUiixPuIvsza93X3w7NEn
/jxRvN5qFBVT9CTn6lox4QoJLUjGV0ydW5UpFrb3ECC0nGT2jKrnjPODqDn+wej0
`protect END_PROTECTED
