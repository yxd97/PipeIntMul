`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oN6k+Tgh0o6lqqh6SNd3Y4sfIs3CA++D5BxDVkT1CWXuEHhqNdrfMq3m3TRiZYWO
0GcZ/DOQDkiUUnn+FRQ15EUQPiKrkRFWYOU1vb76tqNsq02MT7d9FbctliIxKxsk
83APg+fVkxVwouosx1GLAZbOziwDrw2FrAqX2ttqSSuptJO6sa3YQYCWNCI9Sio2
AV5wYnCpMHrZiwJShmpBSXHouRu39vZk/fv6SIL9U2CupxDe4GINTgU52OHpRwts
677sxsSadFq9vrbbc1THWh28ycjWN/qjS4xbHjkMqK1HiSrYQKo94uPEb3z2WdBH
Nn3cszo6k5qlz/fCViwurgmpXBl3PJCXoRa7NBWnHRESNzhiKw/r+VR+0AOqJL29
`protect END_PROTECTED
