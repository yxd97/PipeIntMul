`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPddb9wcLZ25zHqIgUAekZzznzmqXSw6Z3jvEn9DfBXsFU0FOEpxHQgP0AK0MXUj
gk4bdanxZtFcX0Lut6auHPBg6w0EruqQZwpAmkIN9JveNj/sI2cSLm9hJn+xfrnB
LLlGQ4ZAACP2yNBe2OwORxlIsrVdo0hIqfq83XhQuv52FHts1N3Ugq1UU6kwh15Z
p/IVEni5Uo2UFFyFW1ewNMYhbn/6ZaWjOUfX9Mv7DDnyHCTjlCfl8db3krJTtgBL
2J+d1Nz45t2lzNDCQZokGuOKsFzHaK6PQC0Xqwfyga0Lm4k9UklMYtfPFvP3OV80
B0+3MciVTMot/jiXgqArDLrKlC89FURMG/IKYNeBddBWrZu5eqM0yY8Z9pV7XIZ+
U3l0A7t0aETRNTo+iTX2jYKP5uCDkbQDCrX7rN7VkkEukUh+HaPvNr/UK50rMDq5
`protect END_PROTECTED
