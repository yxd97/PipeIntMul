`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UYsWDU5gNdoo++m+JhAXSoUZndeLBYTRzgijUH3u1cB9Rj92XO3onaXzEuP8DXQv
02t3sGT7KS6I9mEsGKq2a+nxS9uOpSF6VCcc5ki0dPpylizYEJxOhAjtM2tWEGpB
pHa8ioky9Kdp4TCpbhTWN8tnspF2hfSk2XVrS1ndmFwyPVCY3DOZPIDAyxDZVUN8
tFmMDiIBxo34XWhOtWJO3yLEYryTf9Sx2Uj4VcNebbQJ4Mb+u49HlmPFiD0j2Ode
1mvxHVWg5hGON2O+LigNDdJQ4AZ7n6YMAXmhRDwjVGRkVGEX8CoNl+e3pYlZiKPE
AP5C5s19d5vPInCsdmKDruym7IDGlz0+3rxh+pf/P0nqJHretmP2RKOJTGxm1a7o
T1CErwdB2qBKu10ItM+4onpeJHFjR9v2cF9v55FEY37rZ15dsG4sBYSOSkk6+wqV
9rXEvJr/nKacrJYuSkUv7IKTkWjyG9rsAna1R5T9jolNu3dMQyiNRpuSGtgSWh12
/CHRYKZRTQZL9mMnX133VEIRtI6bfZUTF8/bkZBu28gvpI3dxITuvHKhjfT/lJ07
pYLJohTrKBESwfkkxQCUJ9Zz2XHorrNjqEHo+ZYr8qwXk6emGdgmYVCY8MVBKuyH
Iz4H51Y7d9pniDQljct9YtH46dwF8vFq4DqE5GW6DBimnXFOxd1xtHfGcEblKp7S
K9ODnauM5hDVQh48Qaz+6wFOzSblNqP9480jUN/iWhkUgp9ibUs+x85LLeXdHwxi
p/SgG8EkFYVAa/czPaek7w6L8bn3+cvhwceuJZzJmr59G7EnVyI8hHjFpVauSUKI
FQ4+EBOB5PIQvuFXfKsN4sN33vzP/FxzCQaHx9Hw8BnTIlKAE4SopBNHkFGCQP3a
wBdlynDUu7PZl1fPgp8SJXqlaOKIG93W5/GB+Lr5KYm/FR9LerWxcbm0jUTHagFH
OUScRONLVif+ImigeaZdre5jKVzOhxPKWT9J1dP5reGZ2DZeQZJkuYgrvDj6JjcK
ppQK8Qp2eiwprIPmeyc6vJ1ykJodiy8lpicnKmIjVMMdiswRhAopO591z79Vp3qC
acS9Lw9KyspFiy8G/Mv7EXBuagfVOKRUmsKEL3t79ypUaXV2WZDKfySo49/fQtZo
CWIzlJ38yjhKywY/x+hHBwHn4HzzdbFPwYfB9OSL/G+UbB+yvaYtZmSdR1v0qv7L
TefnzDvXqn4R+5lO/fc8mg1xZ0i1gFrESqx+E20wxewdlBAgczkVHsSYIPYvjOkV
e8LVexJ8xttdzfjrrkkIo4wEw7nsg92gtoiPoWYQT+40Ka0eHyqh7TkBqGfm0OTO
Lvigu+J1kIskrolC80N6lVCcIhAQL7jSEF3KSo4EbmExgBFAvVGZVrOFcrcJ6o5d
p2iLZmtPPM3riWufWl7jppjcB+j5XRreK1H45HEzGKQY8ZULTiUp/pbEpTejLVlj
qaBiPJYEWjocccPJRhwWEmSxWM+zEyKEDo0LQgBzsP+OMM/Ny8nyBEyquf9D32Yj
ewXYgKWtNoGbJDlbTfWuD5DnXbcoEDJau7/jPcZ0BDQXUd8O73GZA53UKeTHko17
A5hLOBxCOEUqHmQ4+VMWWyICmkGxSkg97fzWdLxBFVnntHJcpb0LffQAvpTTKT6s
EQSUIyrCIwhMJ35us/2QFxaG3dnpjEjaoZJNSaqrj8VXXeENlIsA5jjtEv8HJfLe
bI8RXglCRUjxTMCYEBYqDhkkh8NseaigAlDM1SK19oEE7m9XxClvG6dVjliqCozY
HG+qSxkF4UvYmSBZDgv3qV47Q6LpGmyuGL9M7z8W7zWH195siVAkiVMxoLSsNMSg
ONPy3WzHe5ulFt+dkfdKIGKTp05zQ9KEWmrRAPAOweUE+1ItQ0fvKtolwgYwN79h
k8pbSgeXpCCwMNWBXwfJRVp5uWdAenC7a1dE+4DJ2rKaYcESFa+YZh4jEMi05HId
cv3Dd5oWMTXX6ioeQ3UPCU3rWVPOGoyGpN50ImWFpJ9o8r6HadgwuydT/Y8xJZ3Z
wVWe/xJUL+xN/6CdU48rGU6eJlNMZSLEW/2U+ZWEkfCrsBqjhZ+Z2MDKqhT1XLR1
r4Y2T2zQ8ZURmInjMc/+wjd4XXlYBXJgzhpCPRh6/R6Kz6RwxhRkp8FrKlVR66TN
nSuPWeQ7BbPK+Vqnq1r6MTSNPFPTN+Dwny8h/anJjH8cZbcOhAiZ9bUQ63nh2kVG
8dMl3a5mOXH6Ld96/cxJxPHgf15MbLycZQmHGE2rZhHGBsunyCBxa8KjGRzwIOLJ
34ZdgLefTLXaPTtuRWsiq5GQEOtmgZQQ8wADdESKLG4AoYZs5nySEJ0p310wzHFI
u1ghxBgq+maChyZnVUk8yVqixkmZF/X2lVBjjoCnP7kotKhXotcQNiHFu6k4iLRE
Rq4DrtO5F0oZegoMNiDKKplNGfKBAMlWAi8S4cqdL727h/7ckA8r6y4BhAtytGc5
L1noTOw7JF0eTghBQ6RYT237P8EP1GfLN4n8mvIei8Vy/0eFGhsvLWoThqvNeK3X
wO/jKEWkCSkdaVOJYdV6ViOFKwyU2E8hVWuDIk6n9txOIScuNuFuyxpjfpeGWGSR
TPO+LqxzcGJWk1tXf0amt04ZJ2peEaGJSdCa6BMyZKBIuL/ExeYGpwwrS4knHOLM
cALJO5XD0rX1CJvdUGVSlm28HiVkaNPgousb75vzC2mJ6XfwIZYX/EhzGUnF/ihX
coWOKFwzg3zfqumuY8T2wW3eIyEaUWLmVxRLgDSxnQXvAClct9d+D3c2MYZkMXsx
7L/iR5sQvB2L/kdWk2+p0WOhwVoxL/TizKF+T10ZPrVVLkJCsjl7z6l/SfAz1R/d
yv9vWgtIa81LRtNJyGDayDvqSa7tC/epNq2cM5dByfhnHA1zp3DpSLpnE5n6roum
EJzptfThU7LrEWIcnOVHx4xztq8VTQLKqFYBIn8uLuPnqQ5Co4L4LbviDw0f2Q9R
qFbIjyIGiiKzm3jt0qKyANd3tjjOZ+Mt0YWHjfK+0b2w4QN3pXwH/Hy/TqwNP72X
INghSqbuqNCwnW9o2Wv30e5MvYzm1LJUpbVKT2jkhmNYNxohb2KeIs/eDcT/F3n8
vNQ7Ie14Yt7D59GHlH+LC3Dr8bWpbgMuKXcp6TQVjwER4j5HFsyXYT2RL1XKfC/L
vMlZYWc/hwnmfuHmpkZqfiqWP29HWSJ5dliRSDtxrrt748qwV6L/bJyZKibeT87k
RqJWbjEyBtTu8kmhUCx2Ow4R5+C6o4G7xtQ3J4ua5b8UExbFmNSBr6UXTQLtcd7i
cvjXyXyGgV4SGOhYScw9L7I/LjfV4WhndIXCzaVVQqc9t4Bm1bkb6hzjoLEgbj8E
ZUREXLzXD41YBiN0q+zbUfz8W6DaLMmWfW+M/hMXomQkEmqrpqYmPVzSqvjOfm1r
vtt6Iceh7D95hV8z6/jlIPgcp3Q+J1ffNVHooltjgsIJx12tHrBxWNOLfHIknOzY
xVVPE8VqDC5OJuLHTdOmfVFfD89GizzTNT6YjDA9susaz+G/VHMWMuVBEZ6brZn8
g1JQk+RQW3ssNrv4eumF/wNTYXWIHIrdri2gqajT8He6EknU8+1BoQDZmhxzobzT
pGryD14q0qawgibiFm71q+25DzyBArZo9bsZmVYXaIBvZrt4AsQfQquovr88RCFY
WE+a5mAuBzl9Xc0raNEDd3voQDbDUMU1X+1GUEnAXEkUZt+G8HpcHp/CpiIpA/wl
veNPf7Vj5WrOUkw3EKH/CFv6qzuvmQct7uYj8TaS/T0uPvwBhHmtGrcbfw0l0Njn
cjEnOgZHVbNufjcZPtlVDmznn5T2RdWPWT3KVCaTrA+Cj+bIdTMhVe9TwamFR1DN
Ir9VijIi5vCQqcOTUxFCzTzXw64jcN3jDvi/wFwmvCqgpijBc1SsTzenju/dXMnO
axaC/d7irh4VGMfShsS6+cRGepYDu+cnNcSM4fdGKfDr1h0xCE3Ak7KM9OEBp9VB
p9x+L9j8ZsbK1veupSYpNAtDzi0vmuVjzMRUEWCiR0xmnhtpv16NhRv7752JmzM3
t16AeXBNypMwWF+XaZoU3yad0kWie1/E1WsAHAMKVo7Z0lq7L7pGw2rbgCTh3HQf
JIPRBfU5xAruueLpdXocWF/hc2FltXPsRS7QWbfz/YeV/NYRiiEQhkypuqib2Npx
OSGFJa/1f+M1HJ3nAANQoOq4G//z9xGDTxC/9Z5JKoiRpDHupFFxhZgRk/iyHpfZ
9sz37TXc9LHvqdVXTghYS6aBwHQ88Q0TwafQXsXH7LCYEC8YnvOlQBXlPAvIz3nt
BJU/KKyTwxVxkmUKZzq+9UQIpTDPk1wgRDJ6ywf60xf/gmeZtyCaLRxh/DQgZsdf
FiFWNOmZe5q1uCxbW5hh7GSeStd9rpBVQQYlgg0KORpSYJMAWWaKbHDBiJGiUzzH
FYJR5uoyojV/aFk9peCQ0ecSPoXtOpj+uw7qTj4bihjrG0SAjJmJxXM/LmYc8WJl
8mYAXTnyojrhEZNflXkCJP11RAcPd03NfQmOBFPdz6N34SuXIlwpZLeFUWAccC0T
QtlkeHAy5z1nyHSoYaB2IivlQAKlJW/ZsQbYJ9r3HUl6YqdksMof2vVqcEWkDzyK
lt465bZMCksutea/xkQocqe15oeKcafEfBQpdHLEvtdO+5TEgfvvhn3WGLlI7Er8
qOxMAj+VeIcioIFqqZkctswW7Wf3PvdDeXx+oj49Zq+ULca8SLdNluS1bESc8/oB
6wsaN/d4LSM4wh5CvVwjlLnb3HZoeDY5beIP2pttc6cwlABt6w/rahJZPYBpkoNg
ValxZdDoy5xc60Lw7dnhCc0ju8p89ugP4fVih8CsqsbcpEGszwmuEmB19p3sURBF
5/Dw2JWojGjx+ZiRVUXp0KDPm6krqruwyL/Aw7t0JLuU45+1c1cLOuRODCV8oMhL
seH8I9cf2KFnFRCJGNXC5Jamr5dRL6LJwGKu0D41m9+/JR/guveCqbHb9BqXWJm1
1H+7xevcIrMihUXeG9CuPj1yUtExD2dJJ08VL80Mg9xIFrq7PGYu3qOuFhy2LtvZ
Z+3zQabJmBfaokYHxaakXjJITJEseesl5k57bNO27aYgDw9CsPAljK8gN1HczBia
Zyysxs8q53uekzErCh3t/Jnj8jLUB8JnIfY2NzOSoUVK/jCJaUHi5ayS3Fr2SPNy
LE2ApFyNPn/xNPMWDtLmL0QcBX+nxOwGdiX7KCXcY4J2zyQJn1ViyFynvaBfzX7/
mTvJxkfwVHVqQfUb2887+h07qr4crZUFvzIt0adCdTIe+QuIxUBkkhqSZiwGHScC
yskO/nZZbugFujB/SitaJIkLOuPdCkH+3KF1O0oWa8TUK/6vECNS0eI3yUdK8sum
vqKT2jgVycCSVFWWYiJeF4bxyXIOBY1dop63otPZ6h4GEuUsExwob/dMX4IRQUuL
oh/Nf69wePepIvYhUobFCUycjjk+xfwJUjbE8ACOClQJJ2aZfI5eG8i6QyefRr16
MU6LYewfcxl69LCvZvojk3t5eU0QKJ5D+5KdDul24DfmfICnOMIfXU26JRVx4Xe8
aDaCrrVQWciPrNuKCpfMQLBHG8r4xdhEydYdriSnZLugvBeTwjAU3D2+JVxpBVq+
icFGoxSlM52k8dk4TAgDweah/qrSUPq9noUl6//+vZ5R3dgOy8DNC8BbQ6ROE7mu
T+mWlZ7jjn1IOUrMclZipxZFV5TDGyzxHHVsHOmfGdTkiMEjxQK12b9i48fWVFwN
a06Zwh/aGihgIc1GpW593ztGx/EtvnhqtgZ09KX4w8L5GG+sOJdI3UeLMdTPrpVX
pCm8anttxfSRK6QRbAap8/wrv9CexOa4U/YVNHlCtHSKYZGCUvOBXJbRWw/dm7Tt
s4R83R49WE+TavKhJt7ppJKCepFMUP5Rd5Lay6V2m89MTgKBQOgHHLJ8rdSKeieE
0kjvzcMWKpESNptI9+r0l/bs+bKWxp1nfbAv0m7uCYFQfSY9vLurzZEMAtxZCNCO
y/qEybMBUz7v+gdf3iDq6OYlRIF0L3ZM06yYSf3Xhjl/trC5TiSa5T6Qz9uGS2+P
xwHpjOHGVshmUBGvLbPUCZrYCXxXZHM5rTxibVEvezcM0ov7dIrwRsLn/s23Z5+C
XQKaQAS76fzvl7NT0HCFVkTxUY0QjKsjxLC794PzoJ0Bmw0dI4FshTUcJSWUx3X8
r68jWbQ6O77abKuQfBdOwKBBVDBFj/9UINYO36tGCy/0O5wZWIxP/z7Huvh2yi6a
YCFs8OEVum5HkO016P2n04cxd2+OQxpgeTjFz4cYSNczbCTuJa8WlAmDcxCBzaMO
36ZUvL1Xd4jJLFVORobvlFVCZ7J3/p5krRKMMhpjjDvuqzBDqzQlmFSEKL5koUMX
qS5J23djKauGu4d2X15GhscyW9wEE+/Ekj9RrAw3o72whB10v5PYn8GFBVGIBRKR
egnrSAvrRrIxgFpWkIoG8+Ly3Zn+9r71d+hqlITFxXGVNSzMmDOnOwCHk/OPrY9R
OZPzm6hnQMsz3XpNyvyMpO+i+eL7C1OzSmDbrBdz90oszpmAGoQ8PHDk/4zC2PW0
00ey7whXwluSLMqipoqyfv684HYyOQBmwhRfTmzjNoAm9QA8OIqeDoIvYzKxW0Fq
BqLB4mo3GRT6d9zzqvKQla0yJ25oK407rs3q4MI8fbPQuIM7yLleYzzpZwWv21kf
aEYyedIoF0sHfmXefsBlBYpkkJ0C0GHpmYUBwu49pLlSMPxViW2wxGAF064v5h5L
b7adgB4KHGpcUfB4pZlQnqTXgRB2DOhZX8f6M1YDKEGk+x6zubVIuyQ4vBKP8yt5
t7pH6oeFyFT7wDeJuD7oIWggJFrdHC7fq1Lp8ntSN6aFaIkzkkqet9xdcxESwHI+
xHZSRURAbi2g/yO1kFsdDnau4u/zbf22zwLiFps5Zcuv2JO3WLrkqspW2DWVhBC8
7bRLqNt+0owIUwaD3zDeBWh/nNy0mjVjDjiFjSeAvLh0H/KlAY4UTesmI4edH6Rs
yTnjSZnIHNfkvMeiUnyPIIZQB5AJv7WhSeo/SZNKpOr8GfWh1H9HTM0pjD2wivz0
Lr47W7gVzN1p6/RrY6jmgtxBN0OCMIArSQO3A9wyLoXOGuQIZqALLg5M4aPnSWEs
KGkBacg8vBzLrnScCQi8BBrJlYAMRDHdfFbGasADQlys/B2D2rD9X8tqwvOPZC5h
j4cEJInq3izjwFPpFIIEnPqraRmyzh8DL+K/E9qsBTheORAOx+Oa7WONnaz35ODt
zgC9bm3MWkXU1RvETnoW5aaiIWw9VCVCjcBO2i23YWnJksQkNit3JdyeAbwe+4TO
e8mNxNDyA4+613GXt/3si9Zy9uRq3SMetiP9oAEafIF9dwESHbOxT2LC6D9lU/Jq
HHTPxaFfTNC70BLg5W+Ts8pAqfbuiMrKdKt1v9Nn2/obQBgTpFVT+vZOQIPTj4HP
JIumuJVtVfmmZHJ4NBx+IsAnZ+OJAGomsOzfzeFG8UMJKYkuEuRN5CeSz8XIWgQA
qFMK7n8LaftV93q5M26HmSNXJnmQeu3ybMKwtih/VJmyPFa9veBCw0Uy9n2i2r8I
0Xe6zWatzVI+wcg94ZEPRRVZmEzxXUoB7a+TODSm1jTCQi6Qmr60t96Uo9gR0nk7
Yc+cTGBWpC3yspAHk2Sf1bsKsG8LZ/1w861hTzkZYgA49AGg/b0q9aCEx1uShPO0
v/qSA0PqCLhfSmFMlyLZ1QpKndznMQuH7PvjhslYT1bHm35j4wiho6e01Jyr5WaG
UxqjD8Plwt9Gsa1ZK5zAO11m1uWCkRs7xyxfO9GMbPBDKyR/SqZ9JtOuDMNgMM5b
Q6KnJmdDZXz5H8CT+q4ZABfwcgxkxzrb+unG7IxFt2s6wGuZ9uqlVW1tGryVhHhu
X2ISPc6Gdhjd/+nZr2E95vaKTfn/58dJHWLOqX1rI59NvqpuQp/TlKmrF5B5OohU
2kVbnIUcyLP/XcgeMSUElMfuWcMp35KGGF/2Wvf1L2ZHvgqlfMTD0Zv+NWxVVwjx
35rjvooYwZHvVtHCw8xBE4RVgbTqVMe8XzsMH1Tp04O8Jym7n+gAMypgIR2PSTv+
+U1kDh6mUBFrlaYdqTX+HGkGkXkQVnAXyuWa3owj+cajai33jFDmUDklNGlIilku
Yn2EYHo98tWUYmbmv5n1LVEW3OkCvizhiTG8Poi5JMmayJXSbLnvhWdE8ApD6AIS
cNw086UDa6i+5weQBxV7R57dKbIVbLEzcC/skxnrnm5WBPHQW9QaDT+fquUiCkVk
WnX/oiu8053HLlNr1soUGZyBwYMifkW2zdGhR5sOZBMs7NWWN2j483iX6UEFQk1v
hNWBiHnK4GIPNn+qz0ufObSySAZFy1gt+1ePV5oSBO9LAc+IP7nawY47qVYsxUL1
P2MXKYaF7H17tfo1MMT971Z4Ixtnbipva2KcUVLeLbPOkffpCODOu8qZ/SOUxLIq
7cwcZFfwQasVWjlwqdmVLzyaXmNN/5g4M0prO7uX6Ho0xnpMRGhi2ISNi+CUsIdX
Y//D3vN/IJUJxkI4pui7Mm5eGAFBtYXwS2MFHW8pABi2/PH0/wJq0mWRNVCZSPbJ
Qf7W6hlS3THgAg7wtPh5v2WPim4Sjvg5Jxxyim+j5qIBtUmG6spb1v4NFIWHhTwv
iKHmv3Abf4dEcwBJm1WwDg1lmeWnUZ0BEuF3JtUKxck7A66ZzR5mjuIsN33GW1vh
OP4+dGHy2DQfLDHZ+T1O+grmZM69oaUWmEe6YSyU+a0B8KleJXp7pUxQFC4gwtCC
Rf7XBLySlJ3NqHOo3fyFaA==
`protect END_PROTECTED
