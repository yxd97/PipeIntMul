`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZhhWOmpPUWJSXI1bU4f8qOkz57xRJraIyP/na0ubUX/D/zXUOqgmq1pvnHPwDvs
Kcw4gvV61j6qyNVN1nwowHueDC3OWs9U/6hnGzZsG5sTq7Q4bIr1JN1N1YwCy4bq
2yWDKbfTyqONHkJK6OtHlNyxtioF0jQLypTQhehB1bZL0qqXOqk94PClkD0ilrjK
Rop4rz52/it7oTSiOC9IoOGFEzYHuzUUhWB1L5ItkFlnUnaiw+/NxIoSsVriyct9
3JMH0zRhm53fnf4jZFgbZbHBEItjqmJHgKuID0P0gJy2D7wfLMeL0uod8mP7Y6Wn
vlpr/lwbG/j4GxUrc3gJcfKTgUzy89hrG1b66MaEfnpGmbBtuoFK4w9koB5sBC+Z
NFz26sbPSesTGByYqCJad5qHK1Xz4mJRjXaQYuitCjo39H/o2s3tRS7gy+Ldp+lx
1UbqVTzBO2iwknEcSGGk09bU/DCbJjZgkHNgXkuCVF4=
`protect END_PROTECTED
