`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vC2ISVMvDHU9HEs3hZoe+ClmJZzEW1/fV/BprA/0ZYQogDf1sMZIBmQOnn3+OuSk
o+V5WhwTP1TARYx6aUL3oDszmBsQhTp5uj267OctZ7+zxpbC7jmX8+l6N8TEtC+6
bYrSrOmBUK+JdnQrv8/JoLNZXmjRZ+Op++B3MRIra6R/1TmYAfd0qx7cR2x7aGeD
9twGw2jk5UCO9ihGHPNB8Us2B5i7JDZlZUqSWKSllNBGQrGmzREY2DEhbDe0bJQ1
61GAHVie17b6hpKcBFlx2jyh8TEXDm1c9wEVXDsL0ivoD0zIqeaxzopPOp4wpuVo
YIbRTc/i12JzbUrbzeOZcMznbTDW+SyB2s6ukUd4r9z9tLlmy5OsWLZeMO2daTq0
iM5oYakS8Ju321RXK2EPElw2RSK98yCFWxZFOVdL9Kk5Kg8P5nnF7pz+wZ4PmoAK
qQmNsVAbbDLzy7qC1LtCEtMUCbPper5QTQRcIan/KCNo5TPo1Vjj2I6hle3pfMsT
9+PpN3Rs2RFJOzL14X/OMDdehL5bzbhKlA0pqOlGkRxVTzzikkXWwaVgzWHJurhC
6g7YGqxQAsphp5bN+zlnBWU82sr3SpVXio1uOK4/IXG77XXckftAflP1jh2Ug/+D
mA//PmBArj9zV1cghhoADvT6oCCu6iLsZjM/20ylfDWtZfg9dvYB+KbSrtKcXHT9
PBOamRABfw013BR2+m6GJpQT/HVHJkZ0o/cRYhjlYOC2FaVPt62P/IubiaCdl2Sb
1/Cm1QV5Xnq7R9C7i5TrHreJtoZZ7MDJUHj//b2PqZfo4a7r8tukw8+ustfr+pB/
XmdzNy/LuNuqP/KnMgRJWDgJ2nC+3Y62VD0BrTWeXiHvfqoxfV9aIQ0N4LYLX6gV
JNM7xhN6FBI2oG4zSy1qEAvNgmBL5JqdFy+RXRrNI8+0Zx4yge/ZLKdlou4xRUlv
0xQaIo+/PkENrNToRHTu/EfEUE2JWV83mMKZnpWAmaHSItodSqIMYW5UQ/457tcH
8oIWxpxaXxeExN7uxOG7BHvdEJRe7MNYVAKFfWJEx2Q=
`protect END_PROTECTED
