`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W2vAdBAMZQFZH+rORB9FPct+DS4sRjIliWULwwJGxrOneu4EO9HzsaXeB639Q81t
pv2tpRMKTYDJVUnAZtDJzuAQs7ivhAJveXvUgB02EX7aPUkledyYxG3YiPOaLSBX
U3F4Z8UK7cfQx1xBSe/a9XwPA7NoX+6e0S41qkSxtdlka3kqfkAzNevaqzHlKi9N
D7NmZ3SxcAQtTSO0auzZshVSjmbDI3HLQpzefDYTltU/MbOq6Ax/f1ZG30tvkqd6
asv8O7EA0xk3kNf5TE2nafV3hqW/B2e8Xk24CVMMo5jOrkXpsnL38FP/85ZFKRLs
8D8xnvAgCTdg878dfbsVgUJqb8GowsJxlYJROWk0AYWAHtR8435Ctv6x5OfIsJst
59BfOzG+TdqEjVW5rx+CRs55SuB2xKvMLoKxncrbvdC6LaDp7ilo0ZYNt7uIHq72
Biws0bqxwWWg1mGryPPNJX5+VWBYNxu243WFv/gjNNVKmfB/UOsXpaIK6rWxFDnT
75zxDzsmlqlno65DTKKChQXRdyCtL/j6H0adIzUN0mmY9TnEHBrgpSDVWqti0mvK
ECvFyOgnJvAf6+uanIHudQ+RddZ4mvePIsOwsklANprt29nnJhtcPNwpCs1yo/vU
UOzrYRtQQY1FY1m6FyAjiPX8R8lgYjeiHSjj/yZ9ZNdgj69VdcVSmA0a6Vbt/fB9
4Gn7sw61oHimkTZA5vEhHn55WLlc4eZ0ZITDESbE5X/dGw3+eCxqe5EIrTE7OWgQ
wh4djgiXzgPWzPnLWkEMS1oNdIvv7xrYKg2PwE6OKENrLIj9GMpH7F5OPXOxYd5p
j1JXzLdB3lXk7cMswuhCQ3wRm7EZJmun0GcO08GFBa8SN68hCfrCM50o/IIK5VEn
44M6lZoZn4KYYx5q+S0gDX+31lwdDG7PExlIQZmgYAVzHmIwmDcxS00A54FEUyme
e+AYcMnm4WLYL2wK/YDoLBDmpsnF1POHgv2FpIbj4ygX8n5l/4e5VuF1kcEPVsYs
Nf0+W8xjjIKwcvwIUtlOBqz/9hx8lvFdbc57ythK4TYgexKMUWj7u6n48CNjNgqc
8Mn9xQGAdMMh87qIjHT12YeUe1PZndJg48sdsd+PvpzAhst18doiwrn9GUExCQvy
ZxpuUw1NlePwxMNzJ/a2OgwTw5SHwR+vkV5Ux4zhi2Kd4lRZLEYqvZIUgw4+GNah
kNwOnGaMfZB2Ow07TgAd09c9y+AvVe5F1TyrznDhRXUnmWw+Yu7JGo1iKZZe+2Vc
MdcJFR4rpMOQpkuj4HDwIWURe0uJA5s5+0ctcQVNdpNDIJjncGvEM8AEh0bMPBgj
5PtBbYdxFBc57Ipb8krM/C9SnAIhfXD2CpEMUF/ZAe8uLcIALcrpMRn8u04uEdF2
D3VfX+JRT4Xxyw6mQ2Hoh3E8zk2lrC/z/EL7l7PHFybkOzkzTsulwGC5AqaBKhcn
w9EmnnC/3bv4nkGg3ZY0Sf5UdGoVpucD3+F0ipF+Ce3LySb3GKqLjMCG4xSMwKhR
ToqPo3VR5+ARvjh4zizf877BSsChshxSj+teBvMYQUZKKhF02ERGNVF/b7eJ0QGu
frjuNR3xV1kneFxYmdS6UpttAPzK6c1bNlCznjL24mSWfZMWUo1hvJTpmbauBubd
iQj0mAtPzU3X9e/pMaeXWUExZj3TnNpqjiQayC6Bm1c3lZu0ohe+wL1FfyvTpGTx
FD1w4s6APHpQafapnFgF3ueck5pUHv7K/axM5pRrX16VMRIt0T/dR56ktlA5feXH
RsixMfflTQwL4YZQmSR/lVlCpiekjB19OmVgHBzaQOeddVjUIYU6bbSCqxhOs8+k
ji3CQPDYLbfkE9BHci4i796/zHbWwc1nrUbJc94toYm8DowSGLX1rQ65pJPHX3tO
8x9Z1CPiJFwv1HXtIhplnQd7dDEfNaqNUJH2h7qDPxmLNIP/SXrqrI/OpyFX7Lxv
oTlbsTtuMVd3uzpFk6JPPO0ZOmdeUysCJbC5cYFpny4jdeSNw5oRzPZDfeDNKtAg
xQ1ETbTgpsIZJCScARU/BU4s12ERbYaqolDjYZNS/Dx2GZ5x5Bw9b3x5NRi9lE5T
QwtsEFxNyyA/mwRFeNkvr+dosPUywb4Vw2QEFvkEUzJgLMnL2haxYt8dJ06y9IFn
eCK/S4ecURE6m4OHCEMEPAb9334dZ7UeFgsrUMfADvYJhtehr7SXRwZjf1VFiHyG
5FUc1pcS+J7UVTwLf7l3J227/3mpd7b8IxH1eaxA70m1f5ufb5h1RhbqnFhqNAjn
S8N6ADgUEElMgN3csiYSpuNrMAuUFiTL0mxW6KxHwgwLFTikFdzhvU639RXtGOjy
B0bLTsSXPh6SIvzN0p4cCrZW7c5xUAYuB2gUao0SFj5u6rMF9a4EWVdX/xxGRxqk
NgQ+oBMtBC0SPYyftqBhXwze5w/7UkAG1tysVJjGvp5di9VUSyOya9fEV7fZxIvH
KlLZqmgOfBG6uS9HHVUWF8GCCuO4rooE6bsTpICdro/hJCODCJEsg+AIVt7jh3RM
TYAQQkH2jdgUF/aP/0ewjN3Ymhm8RKFja+9isiOwCG6brXxyKABY2ZkePhiyEqvG
SqOoDOCRMSOqBFYofiRJxqL4qgUHtQXEZtAk0LKqaQhLW88/TSDnRcq962lxs6Zk
nHJocVE+SIAKU9vC5FVRKQARWCCo5KCnLI2FV6vjwaXQh1PmukE8aaq+Lf9a/2Wn
R7X5bdhPLMPiFtPwsNlhwmBpdh9CbtUXOWuBJF4x6nrCsNjrGjRjeQ6jxPQtpOjG
kw0fxJaCUGDNUU7bpc+6hSKcP0f6dCufM2e0b07QvC8Nn+2huaA8FIR8F/PJAKlU
jkFhxc3/7oFBw1GiDVLJOBWlht3OV7sBCnWld/UYedl9iRN8JKl0NpWEKeiJvyH5
d3G2VUrmWecG8UrqMdrI6mBScAXUC5BK/zyvs2VRX+xXm/BcdybcSRk04srcT7lF
MQeK/SP6B0dUyAOwKldNFcryt1DEUNb4B+veUiUpotUCOFsBQMPBM97enOPE+Tph
vUjKn9oHSaJVdzuAKU7TXUAC5rkL1JNdUJaeL7OzJbiL7T2aQhv47KF8uMTTU54+
oxIs2VMlRSUFnf6L2/yA4+MKGbFbixe5Vz0tPVyB5dKLfTrYr+Djynphi2XFUv7M
Pzrn6qPOGb1KtcJu95kMRrvWluIcPhauZbOXXv8yeO12Bh7QP1C/chHqPJzm7TMx
xeMrEtrqTYlvTxB1ksGKk9/zKNRH/bE+iJsaop0KdBAYyJ3bmpuAmGRFwYRX/qaR
U/XosneKv/Q7Bc5Jp0CMc3SXiDlFZVZctYux4EEFlgtjZJgjUYtbUuOLONIUD1Dl
GIvcExJNmLvXHGMToPBf6mNWaGwgLMrRzlsFKRaKysKR+yEloEPxo5rwNnwAb7Gk
Iv5FbzFuiLQsEKuTZ0fY7RYA0ZjWMgdiy3mLnpxvtaGjbV3DJlYk3Ez/WbIuLrhv
jJrwBGqO9Zz2xezjJkq6SAdTBdZAdUMeDEmn5MCDuIuw+hKoZ6diAcr3pDjXTnlR
nyShV3lZXDZ9TZohTkUUyGd3iszv5jb+duSyvcMDzNpQhgH2Abl3Yu79wu/3HDk3
ITAKOBd357vYMIq23rzUixfZSYuImNktN5oUiwdzI943fAG1sBds6FjDZLpjJC/h
lgdWxFmP6om9Ehfo5NLJRDV2HIrwxJzOxOVn0SAbGsFs9/O99UNN3QppjqqSJFOY
i1Qlyc6Z0epZCUJW6tNYDAD6yx+HNx5ODuAyWJOgbfiHyCwa52HztzbRtMkfRm/C
mMIUgwbrpiZY3+Qi80u+FsJFGoY5XJvMccJrj4vyHXV+/Gcdg7JPpQQT2UZxl8MW
hepBTA+C8ERc91BnBRAmq4rhEkp6B9qSsZINMDR2jDWT2pZ80HLxrhn+yahO6YRR
7PGjXPTz89AhgDy2WItsmAz3pMG2uv2tQwXonVsg8gIvdAR8W+Afa/nyDe6yFDm0
OALR6wWDCXPDQQhN6JGcNBB8X7aBG0N3YWwXzsTvAoiF4hTUJp6fO4LkE46jIibF
FDFAt6N8ncsqGnrjwxJ8LWb2TphErdTQ33jDXxecpoKd07fhX5ojmaGJhDT7oinq
DKfyecM0rsKs0Kxoam4Q/L6GzzuzRyt3e9dbf3YuiIINZJT6KUSHKjjho8O594Yj
cG2LweGCOA4G2MWGks+wL+qKi7datGFVVNSSdkxZFTTjqVdc501rFs5CsOplS7eK
cjqXTlN6npSH5NihC73cI8rkRX4LJWnfvvUPmcgVBdxwVfuqetaeK3/VI0E2gLUb
zaE7Oyl3QT+0Dcw5R1AmU9OnnSCzxXR1pDbV/mDRhKAFUbezZ/YgRFv6px5LQRXu
MSFmAzscYVfFbc1Y8ovE7llMegmm1o5KfB7r8sKDH6xPWTOiwzRiUBbzHKa9j97q
N4gCteGPgjEkPuaMswpCVqhvlX+v7apNnr+VgD/cdW82IialS0XyOiS7ooyQwYFk
biIuHDqdxJKVFzqWr09ZBDpxXCGfrZgp9UKCvC6uSvASL9CYjtxAmG+8EjRaV8JU
fQRYtr3j8ZHj4XfdjKhr6Va0uqzWKCi6jDgKKhvRd2qOauh0gOW4bpmeqAJkIDdQ
HNAnRXp4i3KZfBPgAtjf1HGNC0agIv4dJYiKdeTi0doZrEgGUnQdLckg2s87i+61
HW+GBsOIEatVAGVpKOqaDctQK03nYkLLhpMwirn15IYbV+XUfGZymA7Y9fUdA/3o
cMBw6BTu6iJ76XPMiDXuzhGnKAtEceZap0D3bPXAIArMct0vHwcjnETttguwUbho
Z9DTvhiiHRsc6mFXqmAE1HK+4kok86hk8qSZOY1pshrsGdPRQWCHok3hC1yUvEM/
loIW4Abl0ysppvJHncToIaFWd6wgIXPh6LXXcq776gHWRXWZtTGfoSGSGGxKsRK/
PtQwF81nBIz3tEaO2xfvwz0BtjWfdXnYyF+yaaVuMQVIiFAqkK0tR75DchT32XAj
z+VvvQZbTzDDeOHz/P+k3BpeYQd/Ech7G2s+rH7f3PBGix5PKPKsCClXZkbZG3ne
boq6Mk9eXW9O6U1MPDdeTmXzej9J5iJ8jHAd6okCXjML1vaQ3srUHKY7yG1q8cEj
5SQHFr8DWD4aSUg6x+VQ76ICLsCqWySkVmQYJEuitNK5dZayOZRLg68lUVoTpWkl
agExVQcqCMSzPsvt8uZv2djwO1YZYQxuGLABTsD6WwUI0AMaKf0gBBibFGnn/H0V
2VKkm08rrrO995VEQmn0/s2R4F6+Zddq2/bcCnrj5VtJFcytqhoUC+P85nA8RLo/
njhHCEu56bF5Rb4wjDwLgq/76pUXHo75FPah81qtIsRL/iN2Q184AtC+A7pjDnFK
6cvZpy9D31vgTvP5Ql1HcCacFP1qg8vVf66DPPTiOmq1i3Pc5wLOm61fyHPZ38nq
wm/aerUVNrTEvIc0aPAdHALpM3e8q3BsUpWkuQjxrrWmKMnO0UzpsATT5YSsPjui
x+vsT09O3b5DHVibMt1IEtKYCw5W1X8EZxxBmiG/n+xwnFTCWoIejPlsru9Bs6I+
27aVfMc4gtyK9zTo/6WCxYJkQEISmacg6+3SwWu5IM3B+jengi0HNOlL0pblvj9Q
LaQzfFIquwtvPTKkkTwE40JstoT7PTXFzwTpQqbpq2jM62aA3bTfsbDbnIkTpFlf
r2D37KLqRsNtuCJr1PZv4lNmLHV9hLyBCUmBdgdPDzf++uWJcGRU/IqwBa/fz+m0
ltJ/iATKJ/u8Ia0PBDzTuRUCvZmjkrz0hgE97fsNfaWaVjrdAJUUrWgFDvzWEvPG
hjsoTNpceqWW7HHyOL+1+52cG7irpjUUp0y34fTwiCfFJqGLqtVzP4HE4kuQzgeF
yQ1NpFh2HwD3/vrgqIqe5NgoQ/G0QoWMjFJlLqfJFUVC6pMa7MX7ae0ubYm/Y/WN
2OzKPo3XcfgaofQyrQXc8onTn7A2NyFIcaQ7WtEIYngzWOS0jT1SN/JY7tww5iEu
Ow99gZ7pKiGW6uvWbLPqL9R4d4sQGMm3dbXhQIYEBY856v3lFTsLPCPk1lnD2Evk
x98w0uSVyDj0OAc2WUtA0SNWrt1sqwvGHc+0ppzlGoHSygkGqsqvVi2FIi3gNQ8d
EbgAkMl7poeP7FSMktdvu3/4r1vcOVpZUBOzvu7FLjPxrM0duo6Giel9vpZWJEfX
+ozqgvKFFrz/S2TE9MXKBn8v8woqo/luHU2w0YuPnhSRz0XXRIRaXu/hqg0E7leg
0LfttYxjmNBMpCi2NSUeGcawRsKx0aGwiLHP+ZSob1z2Y5oMfkZ1/1YYyRRKEc5X
NgoMwlBKLAwVq2YLL/j/4ArhmTSkhj5S1WJW5oay5ZK19Z9iVD8Yrsn4lSKgv1zy
qZH2psmx5WD0KkvaT6oqPD8zhS1y9lTs2o0Nhsn1FTutSZB0BcF7+IQExQzN/Hy9
UND5sWhipJwVuv3ZAbsB4SpGbsqC8oqnDB22VG9FWW+TBreGpwJIK1nYjHxMfWH2
wVEHvFjUi9x4wB1M7wrEWQBSOHzMinvoMovpRoIosJKmzwmJ0ZvBXVEwXHKtGxML
wVR6K14T25vwMLrB2L7Asd/M2ra/Xlzct+SM0GAoy8rDj7G7BtcnR6VxsEYuYylE
CmDaQbfw0oElwD+MJFTF/6bjPUxDyrje1mFWh7y0G3zoPo1rz3sfSzhMQnafDt1k
c6OMb1SKd6pD7z1RkCfP4kje7w6jobnmcG2NjjfitokdnMT7l2zGhCxVN3eS49lj
TWmSJpVgjrNTsLp4xtYMfnXbNk7dclt1xvMtBXnN/I2EEdouTfTgCDpIdmcy99us
0WRMnrDq3xFTvT2vUuk9/Fz3EMIeLRZiU6zMEwiWc8tRH1jLItArdj6CCQySRtQX
J7NMPjAQqfAAvfiJ1RlnfYaEwjHF8MSQQrcXd3qcd3lKpFn0P1S7AHksFgBPWIbu
MZH6xV4KwN+d3WvSakWsvu2gKofbQeVev6qDHQe1IECmdBNYgdwldPy2UDW0zlQU
d8cuXWPOn0Bk5CoqpLi3KZhhm7ix+33vmo01dsx/yDZG9bc3UBTz2kyCoLlraAQD
3OlA+BAFhC6VRVSdbtTy5yW6cvk002PO6n1aI7ptIHkT7FjzTmgCt3/vtyWAa+VL
apxsYPcwmygWHipeXdONXe+UEPFd16IB/gLk7FqKQchUYmAOaBarq+OLJNchgB37
B/gr7O+yLp2E/522SMXKmiETfXqMHvvGaWBs2duFARSNtFDtzcwHDhMowZh+Hl9e
fbWldJtt59d12bHSyqf1mE7Hb8UO+J28wIkbRhOsiYv3UKRLuAQg4pTTm7QlWfvf
/tzDXNGY7i8RSx7no+OPuDJWJSvhWVXQ3vmQQQ/P/W6msd0pN4J2t7DWv+4XCRjq
6pMm58lUJZCn/OFf0csGgcT5nbPwZjKRzakmBaGi6c1Rwvi7LAgAFxiDQfaxN0ww
urigyizfnbSvyCUBEzD4DYSRf2P0ju+aweTT5qJiERkVwDAhMZWW/zScHUVMYnB1
K0qreBbMsDOftutSjYLtDc2O1Fo8XVpfTkkgKQ1RK5wnNrQnnDDsZex4MhrrrLdY
cP3PUcCVXFGLv2gYwU8DHD7l2iyshdPX6HzGkSUKGYchkDrVv2H/KenY9u3JfrzA
J+jUk07NoCJ88H9ueWxWGAXGSXpcuNU6LaXBz5jyPUBky0waSMhO7a+bNY5GKO+B
Xhs/NnUTzFKJ0xOHLPLEDyNWvFkbDxLVzKUHzcHQU/2unSe7ZEJfQp8flvh1jFjy
EJDvcqCpK3rTCrTdzISC0JQbgPFA1ed/38N+W5+5Rtz++KEeTSeliYA+YoT+2ZLZ
z1PLuQDPTtOJdeH7caMlsiRIvCR6qS/DIIPHRzPBAtDd4CQsWYmgEM1uDSXKkXj7
5HWUX4sdc9w/aIzI7S/CEqlREzK+DNukzjABsTGCSujJnAOiN8X+TO6mnzhDgXLD
mJMJ6re4rmU91Gf1ZCdKp8+k59Dvk58qm08B+Wj8l47NtFyxqgy7L791X+c4kunC
97XWJreQxT4sfFoVfCJ5vdMl3nlMwZLZIApkZMNk9CbehcE3gIoHZGOTfq8GDuUH
FIvkps1OeV7dbCe5tJ8tteiEj5WFdaAZuDXL0yzzw8vbLUhRECDDj2bkNvIL1ICc
WEfEx6wfAua7lryYNgE2l97cRrbjutAsA8Evvl/aAoeEViqZNKz/8BgSVw26bVLx
vQfa7OK6iVdqPnHqYABl1ANvHXZKonz19edUjLjlJ0MPmrcqplVwg7rxg9udZzx1
CWN24BLrA5y8LDql3Z6GbFazQ5LEpO+cbGEk9KnP/c4wPBL60hv8ZJDdxBTpTlMV
DuRf5p1WQjWimSctJI+bXN6H6XgsAtyiNQUdJG0LK0GzrftOmueOO/sP3KyG2yBC
e39kuQyyU97/Ctp/IO747cz+5gOJlUuEmQqB0Je/0zmCF3OhqZnSyKjrnLYRkxv2
SCnJgBUIornK2euAd8Mp/IO/JfuILjGSar/pDDMocmz6LxtlFywMOQoVDPp9LMkN
hKjSj/Sr7MqyV5C+lwOQ7Y4CscyLuIg8aVUr0iOKztHD2f1I/X4bBaTwoNMB235W
C0fi0msuNbzTYKAtEY+0TXwJyF1MvcE7sA3XoBWgYnXoLS08ZMFwadB7VW2ImFiJ
PeGviPP4Ku7ApP1Z2VOL7T3Q+JsDVZSUOIi0/sYUdcN1DcViB5P1NyqIadG+mpfA
RC0S5oWUcJb8JHoLVvQA6VQPdohClBu/u+JKQ8wG/1w6xGuaVWgsQhnU5nVtxfKm
VL4h+DxlHRbn3vzTd3zBJyd+THi8947KK5OVSr9qduDzSHgUsOrOZkQrWgjcLRkT
GSM2nG5QQEZmvINHcHfmY9Bsr6aaD2wWRi9f9VK/Eal3uu0pnoodZAfeM9SU5Eu6
kgdvSgBpSOVfAjM+zLxdoOXuBfxNpMGB7g3Tt8QTdYojZcq3Mmw0Gy5EL/Unfa9x
g7IUqKq84qukeUOlTb6qnUsfkzqJZ64ZeiMeB8kXjf+2YCkXw0yATBnuXuzgDpgu
0XElBBp0B5wFYvJ0xKTEwydV4R6aUK10PWH6ysXEpupfMpTrYNRtflNZGci20CYl
WX4S2mqLU13co0fu0sCB4rQblqb82z3Xw9HHH70q6b6YhDeuI+wklYppLePWRJh/
LQTU2uZhoIk6BuWAzi79odAXNkn3bVv8UDmrhzTAxXbGaRhV0jRqIWG/mzkC7Fvi
1qEEf4jz8Zffjrya1Ljyr+17FtvazLsMvbhyV9vplrNP8/UFnqWTYHCJcFBUyGzz
b1Nq7Fk/KIy4L2bh9goDRXgud3snzQPJ3ZM5aHKnNLJAzWPosMxoq85gwQSU/VTU
PEkRt40WtvjQPLXxPuUpXWtsPnVpSy73nTYnqFDIks86ylcgsq8a4MjqgREogtpc
Fhw4vhjkrbcEmSSPJFqR9Efe/psI6CaMYnIFdrJSybe/T2B98JrOYi/7RyV6oRnm
6YmrhKZgbgXf+iuhHZTdgx0CMPiipdiPKE9kmbM4YgJuDnmzAAAd1FPca5RyE0Lf
PQvLmVPDw9wbaU0R/47XszIEi1P5/rn62ve0Obd41m7RPZet8++UFJesm0NBZLxs
XAGw86SdNLhtBXAM5Lzy5jxOXsbX74SQGRUD02jdzrNWsKn46xUI4I3d+b1LJG1l
CGpTCXv8hqqj7A2vPXXGrCSpFFhVvCUxSkLdiuAWJQTdABBWHSYmx90lflYF8Feu
KSt/HvWd6PN2AIo0kYB0Dy2idGixPIj0DbCwtrhbc+2HHm7NAQHorFZfQHIBGgdr
Rln4+vwbMIvrObwYEJWXZQ7S3Xx83056w8Wh4lYM121G434+8MRsjNMv7Pkpqkx1
UItaNvFvnO702kcfF8NZhBBMd12I6JIFibqvLdc0IFeoBWANfGIsglM7sL0Hczxi
s6ua/GFkVzscNnt7hHcv3JBssNy4KuEsufVy0alk1eHJjwPXKzEyczMh+aCB4vKd
ox15mVBee9Sflz2HMkf38vy0L+IoltS4aDynfcklDdXSkARgipvoyEA6naw0ehgp
KH6J4W2YREMTUwHKeEk84hycIyM6yCTOG0/E5wdbrja5OMjS1C5S6NEMvId0F0O9
+sc5Bzr1EorEygg97N4hbkowbgwflQEH3sVsPZ5T96ySOXIBOFtPsO+xrZH8Su7L
5tj+0/R4JuDATaQd/eznan7866AOyimiScv1+Ser7i9LKYjeKN2n6OGz0Bv4p10F
YJYkmrveoeYFYoH8TNDZ/DNnTE1UaeI6R75AUobp1LnByZWqVY2vB47ddfnbvw8w
tlhVDgl4XBbu+r5xtqr8drWcFkIZ5Ulnt/GOrJl6nN1qKPz+hZkwWaefnJHCfbK9
rcBhoR+akuklUVl9ls+Xmjr2C+mK9N4Wyga/4thKx5TCQS24D8XICwE2fXRxnkpZ
kkDeKSQWrCp7jxyPkF2LHVIw3vEMR7j6nrJD3pYvmPxJP+wNPY1/eGAlX9lEgRIF
8bNCtigX7Xowa0A/U9prU5gUE7xtMrHFFN+coin0+kqo45X+ANu5J6iGF3cYOWzw
iODom0MmQp7hIHXf/XS3QFAwdjDHPuDVm7Gk/2Nqrnz44l94HbYv2Jt3D04u/fp+
auNhhvYin4wcpJQ+r9RHqDx5Tr/J31eOQXhKFOIxAr9fiRMeOaNln59d0bibWaBj
6vrjbBipv1XFENr4r0iImFDVOVMojv3G8OzlD8WDz57Xbkv3WfkanGX7qmmHBiMT
QwJcwA1TLFTC56oez6Hc2bF2Ql7WHoMFtKv1ysVfhJRufC1o9bLOwgRXRIQA9nhi
9rkvAxypgXmkHXhxo6FIekGXpWZwaBvPOW8wEwZHVcIzUrZw676t9uHt0RvzFMwa
CBl/KJQoPqUJo84iybQWVl2mVmcuj18dstKZyU/nVN7T4Y0+dsy+Jr8UmtlZQEQ4
X/sPlza+igpwe5Ps6xygTJvNXQY3gmc2mEuwL13zr0FITZH3MDCMsdXN6ZNMR6kn
9IZVQr3PwRs9oTT3BwAn/itJ0M7RXHvzXtcJ8WfMj7s+7OYe/mcj7/lWJ570XElX
swhvApre/OVg7ZPzwtp2DIMXkRIYTVjftr/0DUZF3iDlory/bn4buKAJ+PWvyV17
EmlAMI1bTdJZdORMA75KLhIonYGf+iZpJSzF9s2owlXnwoTdUiECoJoWXNDmDF78
h5QQq1OvhzTrDtjEu8k40MtpkNlBQEFFnWxrtJC6dlz2zJfOR/8b1gtQqyLhdGJn
tCgQ/ZE2IPWa+ElKE32RvUvVm+w7y+9BaSoYrXoBC358ix/FMD4aZYRMPOQgstNa
oiIbng4XmjHXmwn0Abl+rnVOqNjq38v4Yg9Ns+mTkjtzIpGRVyG/MdZzrlmeX3N0
xLA92SVEnV0ikZ96RkJBWKhQBkffCtgUdQWBk6pYbLBeh5xtPwTaH9/h0vfMaoPD
YfUqi+vkXkDeCLwuKr2lzQXGPYl0mN0UxQB5oyZDrfL2hVCHjyz/0hkDDVg2KXOn
VYEJUpbf1uPYQUBSeUodZon5BRDK1VvSG/wJHpeTMmO1Nb2cBOumpkZjY1mBJf9n
AO7xKkNzQIrqtq5Ko+4nzJ9dHgH6aRJ03wOBLFY9ijEFj2OHcIrqkqpaM6L1gIMG
Bf7ST6LgvlK3+s0WjtVGe9/SXPNxVrkTRD7xFktuHL3vSJTFlERu4eWPTbCULTCl
+jkDEHlVqrsjJNDAaGztv94OCrUIQxXDXAEIahhu0xZP6IyJuiTOWu9hzVXLMDFe
LodbXIa720OE8TX4oygPkyltVlXYGRHQpbZwr33IcVs+lGeolocjHDXVUZzWdvW/
cDYK4x6UK9Kdo0WN7r2LhZqEKVKYHZz9prLeTrHRevHwt7YgvQPsHpxMyFTFAwq/
wF6Db+8Mm7bloN+iT0ma8/Kpg6gYmt5QCaF9qGI4nzBKu/wLOs+db1Tb9yiCYXd0
MTSl3sCoemYcGxG/WTOE8LMwYoqH0OHwv9a0yic4AwC7iM/fUA+5f7HNziQ+3a+3
kV5HofzTwqSIRCjraA70TfR2/kHsrl7kp6MwsInietmK2jHUByQgW4j3Vd9pKpoV
3lfoWnqB1Gy2mr2Oq/yF4c/vdiGtKHWwl8bSGT8MWViWB7AP2kcSOoUs4ePqEWqH
tFSaxL7FZPA3qjn8YLT+v7e+/Iitc4kFmQKLxwtdGRluFkd82Hf6HxCXvw6jFvGk
Ykb6PxMiZ59rGbzCNCvBwckfdK5GVcGPtANk8myIeNJtsMJmpZA8SFX7nP8WXVv9
onjHAGDwzJf4JjsFLmlzJZ34W1k9S9pXDzsTwE7lGIVfWjABBej46eyCjjbty50a
CXrFBMFNo9FhkseoUjqAaqSUbOfrXWflJ+sQmzl2t2NniIq3HeUFm8UAzhYoFZGF
jeyVyMC1ALxktmcwHi6Nn311iBgZM9Nrk2QGCUhPy84EO8nGaJiTckt5LRyqQrJ8
lodhG3twsitOmKAlXNjnQsOYEOU/edJU0MPQQJWZmbkIGWSvUHUKETXYehtSXZk1
CKvVOMub+DjpccyUflueYMNzGlRAdIgIHQcNef93KnGyDtohUEPQba0e9ZOh785j
FglqSVpKr3yZE0FkMo7rAfifXPYS6j0bPF27pjZtrHVnSQmY6eaiA62cBbNVjphG
v7TrztNw8ANzn38f6giwpYe8MaKb0ftZEtSjmTKa1mgFHDuCwjU1T3kjciLfHRKr
ylFJuh4uCEcpm5fh1hA3STNWaDHG8Ie6sjv47k/hs3TnwFA23euB3RDrnHtDxeHO
oNdHN0SV85O8rTCKnjt1xmGlE63k+9dmzIfJZVEDJ1ZGR0xEUIEzkf7r6zuk+Jq1
HEqTmpSm545ZygyrdkLSaEy4H4sRXUHT40Apsqi4P7SvYb6AqBZr5alrenfeccQo
Xln1GpZGYeAwJuSZZ5UgRSzgaEkhaKRtlu/y2XT47vPei1xCkrGrLych1yT9yTE5
nN2R+5OKaqZcKGdUITUvgtEKtm37v2TCcL22Nc8lAt46mm1S/g5KYyzvO36yaUzb
xBd8PHVvaFRV98jlQOniFOrs4syxyvoMF9WovaVAEZhwJIqTX73CmEQCd1dKwobh
bRNx0Mc4lBVPh6KsgCbfTRLgLqGQS3Ijo+Lohyle+W5q+VnUBHRQMYFeIarxgGWB
VkEIc5niyKEZ8P65xYxDZHNZlolLfng0BRHUlTBPm2/bMD1iH8mLGCFslKC6cJqx
9WW5dTAx18e4KFBVBqlcGxDSZse31C4FrxcAmRgq9IlLlvnkz76MmTIk5XOnkabk
61Kn6n+YoUFQJppfIv5CilKK90B9bYrBedLTp6tFXeVPNFvz/9Yt+MiF2UeQAdyt
oCNyOIShOSeScqpyue2uJWV9UUdgzeTbjVM08YMMTsZhAU08/m73fseTNOYU6wIL
6MiUnQp5jZGYZYCMAXtIbs0kvLLBN5eTPdfZfMsM7YR6yCbo7mJ5TdyWEZ7Danaz
/Z88HoQSuHzReFBpUGYDRibxmp8uME9NJwdZD4RRbJXvHD+3zVJ2Y1CsOtSS1IIX
kVK9ly75hK8Z19/wZNbYU/C1Z/mSB6NZ/pb1SMRu1K88S0Oi9c4UUfkL+8+8i6KZ
hIVkXyG9vIrIw9ucwRh9wj81Iq+1DiePp0C3MtX36dnYrql+68Fc+gGu+0W3AR2O
l9XNJ7FO+I7D4oYl86pPgnI2VrEYhoIkecIGijPjQUi4VulLAL8XtjvWp9jG2qTv
bidjQXdTYNQ9vgYB8jv2We6VL2nR8kW3UhMR8HwM8KDdH/Sufs0x/usy5KPgahPu
gkoU3xTXl0cdYh1Qz+erho/OxlFHROhx3lzMO1vUXhExOz0a+9Al6AdhADjDVEAT
bDQRWkNn8XFhILsoFB5XoO6pgflF0Q3pr6axy+mCsTGzMHbrHI5f3qOFJb2JxH16
AT/IHcrpN6FeqFg8Y8wpSP8QpxuRxrH0UWIPYmlUQv4VBg3bee6F5yBmakuN/UCL
hlv0dtGnKxl6a8KDRa8VLIW71kiCVUFQoKXmuQRYn0CZTYtEcE+DcEZzU7Ob0BVm
dsB/OqrDXZi9yVAfPXfiTKNjH6KEGBHPcuGozeYcokG9rfpfpfQHiHU27Wy6g9XR
tXJFvovTa0sLoF+GlBFz56sii7UAmIOaoZrZgi4B20J2jWMxi19YjOzjlRo0JJl1
kON5R8cfXIcLZmYT2MadLsNgFUH+11fuo/0QlsScdNaU7i7WsAu00VuKaTCGVFU2
zQSLNODD9IVo12vHf1cKwLSk2KPY4fpS/dvdTdCsq3mEqhNXHwmZi6JWMeD3A9SW
iCkd8PzZ7boNWNUni+E/hwpazeCX0Q/F6yYxR/KiWrk6krlAfVE6/u/XM9V9ooF6
njr6/y6/Oyy26cDHTzRBJUwRCFjGKUur7kg9qMVtTTDviEe/naIRgMcYOHZPp5kv
bQytYUl3jFTeD5CNAPEelX0YC4fnSFNQXthrzStT8vvABc5ur48W6Zunk3Al5blL
3dMEhufQZ3uzeHYZzHZjaK7HSbUGekEcQCAQWGFbaKMI1Uf6/e6Zk/dc8gd3go81
vzDyVjLkuwLwBJB9gTf4EESien+Lwu9ScOigC4nZYdyh8wKRr9rvTLZDA+tW4YkX
Ypv5oJx1oPCpzlyzw+mStW3q64JwTlT0s7Fv7PaX0tMwYqQRXqzdFy2/w3AoBt6f
WISFtbM2qF65+GjwwqGWYFUV9D4zwojjKhrdRKkTkFzItvLA1MpPoXNCHvg7f1St
k2V3rxyO7TCye25B+XiqLrX2CLhsEnBAH6PYWGGb0vdB6FvY9PfZgmOiQKZvWA0q
abLCFH4/EW6VYLU+ms89g5Gt2l96B6XuKnHFci3R2MvDCmgEbVYCbo1iR7BEbLM4
mT0t9cG33l7jtMKbgOQB2W5Ma0BRhJPs4gSrRwU3/Pn/Gsmk9jhkjZ3tt2fuhjjd
aPg0tmv9/7UksFHSlk0NUGaTKj06wNr+h5xuJlvyZabNAPTIhE5xXKSFdm0VTDXG
F5aNGTN/fhAN22dHJQwdMlrc9TpAoINLTGhvGwrYBReulX7HmdPPPBIT2Pwp03nL
tAEhUj6ieYqOgGeNAA2O+Tiy+AGMHYSAn0EneRad86NnzjEiyvK7aHeyAtIT6G+i
DHbCUIfS6cJkEKA9fwAoqu0Vk4RnCEuNQMfmIQgLdOreRkoeGEee9rRHGg1Nxs7f
MRSa9blSWcZ3y+yDKXZ+P60Y7+F4J2lzWmWhcmDISsi8nYswJAgEqPNzAY7A8RqW
f9ILPje5SD5o4Mqj8nw2cYIG/HqX5i6qnLVd+Svyr1H6enWotrSxaJRtsedOf4Rq
AspAXJy9UrXMBnhn1hOBLlCSgU5yrxITIq2LMP973GWAzO6JX01FFlmMjxc/PkwU
BS5rZku5AslQNUYrA80UkLaA0Ks/CjIpt5tx736CqRU3ltXQxOrdpXIu7dojvMb1
sSlh+7msAn0DLd3zVYh65I0jMF3MCQoLsBP3EJFWBSD1oQ7gytjH1UXzm6kCyUBT
uMDlCh90d37wZsQ0LCIk1oVMpB7bB84TrBpKRzTfKbErIYXfHaw5kDKAEXUHHQq5
Ezn04uAcnKO1u0idiKVGAwaOX7apz9ht/cHY5wAmFbFLH/0/xBrgUVOIuxnARB/I
PGbDMoRmQog6lVcyb1yFnlEeg8x7y42ISIMWBFn0nykV0nFvOfcf1WjxJ2UM8IW3
1MUBnsSkjD4ZM+gNP4srBC581t6/fPtbteWval4AnMFBOqr5/20ynvQvmH75bVDo
3uBzDJVtFCD3uFoypyVnwBi35o89sjMl1hUuDt3VMSvgETC1BroTpAVwcuYXSMDb
hPbUWXNYYzPd/+7Ur0TbwPLeS2UHclMp+1Y2iZFjUAPhKIT5ftLGVsYJwdiIL7HV
zCQxgKUHqYpZEDc2UUxAEMrjiWMVPHEtackZ21bteb/l4A/FX7YjELTgmfcDiZHW
F3sQ/X/iXFamEEsSg7EOiUWrjbemPdwdbKKXp7jNLhPwJvckhgSpjED0Tv92/Uec
fV97UztDMcjEk9DoJ/w2MBKMGpsy85eoNnMkKOnVebLMp+YFn/s7QhQsUzqOb2rC
i0gf0Wg00oVd0ghUyw8RfrZFZ6765Ex4FtoGJIjyLHDylcmWbMDxKvWdcjppQ4tL
SlyZaAIwnebcShglMdILEMXYo7LdzE/hMBj2rrMKnwnA/isTwEcWvSoIRkVCLlhs
YPwo14Na1LgtUzjLlTOvg1ZARg2Qrp62p6sXNtqM/avkz6XRJdkj/HWixlfh+ZuK
OfI704fpeEa3i3+NiL36SSpVlj8PIs8/Y+0N5RHgx9H0e6mdnFSZN2nT/H2rZydu
5bLTmA/24JzhxOdedMNIiZN2kroAXkpH0X/fpXWpL2rNFjxmLafQL1MeGbWG4PP0
k5oMn3JuxCUCfxsD6gSJA8GlnyIXfN4NspJ/SuMJK8vP2UACygkhp4tSJD/n17Pu
et6kKOLAPdmNv9QU7Ck1pGO6vpK6OxV4a/XvI1qCdl3oKLGDgHbuCTJ7eeCAKhD0
M9Y6U7GhQoJKXieQeFzZv2zZYW4gXu+Dqut/2OzStm+P9BfS4ngqFlTJPnZSwH0N
cgS+VhWt/VUkYJjhuTNFzzGRODJ7crDyEPpAbNBdoHzaSGtWPzRUtdJ0V8wz8TpB
G8NSlc6+nMpr4/eqd8C1heoUdNX9fO4ENZPWUYJd831bCxXl5mmvaOud5JaX/tRb
+n1zY20qRlTc9ck29/bas0Rl+UsNvjYykvSab9fwYsYp3ODo5jhWOisdT6pRUiNM
LypKHtbSCne3QjSQvvxo8lRfAiSgR76isEP3+vmgl0Dhx3/PCxNZkW1cH0P/JVwo
PfD3nsq12FzpA6e47J6z9VRaFXxYJ+cIbPk0nL/pnakLnX51TKAtfAf3Yf5wGmu3
llwt+vg7HzMnmTClk31o0No6WMuPcFgFzx4ZMjnfkfC1hVw8TGyTT34OAoeEwdbX
bNv6JoqaxyeTnl0E8bbQO5whGRiFcEe1HDWCsopkRTnsPX0F+56pXwrneNqcSeAf
zHF1tu7ZKiwD0wIKvvwESCopGa/SkxPZoCqiWKPXwmcpxxLVB8oVX2Vz3IigF6Db
vUPEc6VcnOKJBLhmiPgzzmn8wsGOKQWDUkEWK9QFoAZ54a0W5OTFJu4tAMxnKZme
VSZ8tQ9QBAwg79x6vivh/EwSENeJS8x+ofYYZgDmLrpFceB8oOmsgVP0kNakO1tS
X9SqCLwcZydtB64RP29f/70AGej7f3LIWWrFxpti5vWFPJDqYXi4H5cNYxRzqUHa
v2V3W47cIPwdELC6aSnoKmIOp7prlGrnEZB7Pt5KMpZTumzok4SPZUHAFBcF37TS
EXuTrmWO6xyWcJsWiBCODQhKN2bEUOZugX/hvOkoU7GGUJWEXk7YolTQpE/gxWXF
gpt6zr5VQBknTGZO/AiUEnDwruobrQbuiPN8RWmrT7A=
`protect END_PROTECTED
