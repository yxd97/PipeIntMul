`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6yp7NqbcN9VW97R36KfVJOPIyZ1hEwpbKy5LUh9aYrhDNOdZCJk43M0/OLsGZPsb
TXK14FzZQNQ0Gw6tF7oyH2OuAAM3L+Y/oUq+c3X0SvzsBNHBgLHOU0Dyut+T1w9n
2n4lqAEhsHrOvzRSWk0hX6lxTGAnzFko4MeCI7t8bi4KWQi1MAavAJFmEUFVoVu2
MlCcMs0uciGpmVLP2NoKl4MqJthaC69Pq4NLjnWD0tb3IK7PZqGQEWL5vafvLaPN
eIWxWktEeVLYT1LOOzUwVeO5ry8FwnN3ce3g68AieSrlRHNJe/3WoWAhNERaHVt2
nnoyan5YnYTLTFsLIyyI6lI4JW9G7nZAOoWWfWD4Jqgc72sFOtIK5Ll5nqC0sSsc
wXuG274sz0JCYbcNS0GReqZhiBUPM9RUQ1p402r9GrFbvOheqgYtLGw3l/5jHBLJ
3eFgvwZSI1hr1pOw8Qd5sp2d/rmWPrFOM0Q7u3qP3BTIEPriN34yZyifLTN08QKV
9XI0XwPjEq9dCK2KWV1siDWNR8XXt4v44gqV/y6AG5EvOAtv8OYM/AvNny7HJbz4
YUMkr0MiFUlk/Y4V0fIfVGwHTqdv53qa6+j5AaCpjeVyGPnpM9ucInzRwqlzlWdV
TcYjUUcWEf0eI+4+FK36jVY57PeW8P+kEvuOY+yiImTXtBmdtsBXrHZuH/pthUGE
hLSxYPfoa3EF3JhBt57A8rmX+6gCGbYmaMJ7RhyO4QmDcxiZR8gYQXV5iihM3npt
1zYpEJv2DaxnxUa2p7PKZVRUaiJSERvpqG55o6UzCAdHnTBrYCqfPNG+JEcbzoiB
RFupLLT8aHGa/7iJKZIyEG7kWEJ4JVwwKIG2qrRuemra8KHNsE35NawJC98qS2Am
M+NwCQP4l62kjHAYFUc2lWB2qQCSvOnNYR6fXM9c7KHKSP7Di6pw2cgsm6vRsVF5
T1nX9cpJgkHo0jN+PfT1SOv73HTyAAj5PENW45f8jam2uJ8FDxROKhWJfGFWG8cS
8M4MPlSxcdiNgNaiZIQmU0TdYk+LoBSazV8ArXkd8tTRZl3URSKnFSkWGzE2jF+R
dm3CIYUEIVu1/4JWU7fQvoLnKAUxqaAs2E+JV69MobImjtl27u1wjiAglNe1LJBt
YuJqb5323sKUnldh9uJ325KBFv1rsSi4+iAuGQKkOKXTaTPMmzUNSAfz0i1h5LK8
RLAPAaTFOdDtR4Y0EjvDIYuo6z3zxsPl4A50ClChBMpXzyL9I/Zt7HssdCT6dTaO
AA+7u1RdRzqAYKHUNv6hvKyAEzifHaPJ6/8idi9RxJN63hu+LEwEjgs1RUIUSA6R
GPi4jsfNuphfDc4xNB0HdqhXVY+ibfkkQ+UWHc5RwObVPREP+levJjuqdjFj9kUa
aY+VgwNObinbc/Nb826F1XGqbfNKjstF2JQuBtXC15iYUy39R2HzWZajMJJyg0pf
gS1yUv5e2goioYY9mfgdNPSRh8WcmsV18Fy4h0n/e3HrR0nR1akapB9KYdlBWO7A
V7nwTEbI82NCtxMMPWcA3M/fBQMsxYt2BoWMnYxAaQCZe3A+MFBpwGrqUOrUiuOT
DZQRSM65INoNYuufeL30cQpeW6gfClN4IK0MvSXrloK3IpPAtatlBpFCbE2E2Hg7
p4QbDMZ7J08Py76cBW/BVBRAixmdAGZE95Zz95c6xcDSdzLJw0Hmf+pSxPEtDjIO
iYpAMSo5ErrkAQQjd9c1vZjp8BbtbRFL6x1/gg/vQ6uw4ug9hbwqYAv3XGphpX/X
eoBIB2wBIJMgyZ/cdgxr6W8nftFIhQCioVVBLxg414DwfuPfY3dlWIqsvFrFoCZY
u6jvc7aht6wNzmUJCSrN9ew3dsnAzrEugLViXOpWV2QVYhNDQQj+/8AZ8zLRDTgU
nuXG1+f3ugfbg1/7YBvhkE4pNFaVLc+MdUqnuZ1BLrXvmdZs6CVcGxabMiqOOINV
w8xlzyp3Not5yeXVceu3U3aOvxVX3N4saWSgFk2JwWsJjoldUuZPZIPIJvEZn1Vg
0qyk9+Vd5d9DFNTe1YeFdVLZDxNFFdBOCsvUXEvvxLW8DtiovHcL60CKiIgkARv0
+atYn1h1zQWl3l7YI5xraqMYOxk89krPU2msWBO7lo6y2aQiI90BkysDXXPhQAia
siTuZJ+DF6OyCAEdPKkt1uThyDdolDldtzcI6ABzmkWC9zxUB6WpcZ6D40HGXOyX
wK5MZgj0SDQy6yg+VOOJx8eAu28pmsXU3hEDWMldlHTtnKVymS88usfsuCuAfcSv
FZTeMlWLgvNhnlfVNz3Hxm1FR26E7q2OTQkJmoA8/gnmLiif2khzVLscXyQLTsSs
n3+fXOMcM5NIDOMZowZIRcog7o4pBW+PMgumvZSI5jWZryJ6rhCiwtCJ3A67jNxv
e9LpD5SesLDecuiDsALcXPqdx1R4EH60VxT1xQSqXhjbIAzl24MCR+NJQxsT+O0a
EEv/hNDb7+a4kGee3TIDA/R9oyGxCYuOGdBU7NfYBGNiKjI3gLjAty3QvRVm8Y9x
EW6bgsdxYZc3jMVZ3g/WSOfTAxDq2s9Ki699MpBU3bd/KVE8Ji9SOdqlf3mnDqch
KtH2Q5hjpc+3TicPxZwPZiVDO+MEcrnIdYUOBbGj6xX1+P72qi4WoAcoQOFzm61t
Eq6FDe5EZwbqV9FwGtxBRHxUwXPy4t3NArJjbeNRPucJYs30Uu8iRj5a/2W7Mm1E
t9hhR3lZv1V/LShzopTTwxOCL1ImihWFNZRrHtUtfVcBFCjQZuE942Cqf5z+3ol2
4HB/+4Dc15E7/WsiYGQ3fMPKSrPR61K+YTizrJR5BmqGuE/I4um7FHuv7k6+3CZ4
RI7kGxBrJcOKKyuXpdlgsAiyJ7fvsX6JQAJaBcJhLJK7f6RRILa+Ph6iyp9qaO9C
dFAjjx8PerC2W8Rv+Y3HX0+nKYQn2HK1xEldxW3DmrcKi3Dx0+dfXGq2pTgFXJDJ
S25hTqMucH+uDvW/6Cb9LUPpAr7/cpIfURpLn+wVD+FyIG1bhgMKWAEwT+gKHs3s
itujXg4sbSF422vaqtJt5n2dlAp7Odaa0RV8fpR9Yc1CpgRzG1YAk+YyI0i39AV/
z1fBCf5LnN7EUQvOFDBSSVx/Bv8uMB2neGK8q6HvESG6WU+UEL/3cn1m//6P5fE3
891AtVoVJb+R3NfTplsT5H9s7WSCBvhTocnE5A4169JtE8yGLVOu1e3b61GKmwd5
tOfQh97XUEZ4I0W3JJAViGCmTulhKZWygl3+uhR1rALQby42YYCC8iGaQNDZcvw0
XlBC5KFO3s2anuGQw3PhGXkeGVaG3b6o0Fe1e1dOg/HyFpEO44DDOLtii9F4OGJQ
isoIhRixO4rOa0nB8wNdQbRk6aKMltvkD83e16IDc/bC6PiOvWlA6syg1k781xnv
VwzPpPXRJT+xYf+gPVYlDe7Gr8gB110+g3knieniOzai2cD38SZ/jjO5VsYBdiXl
pwTunQxnbEUyRUGTJ6P4zeLohOjB8gFR0RlFOvrJ7X5GsEmU8JGLDvWYwIRrKRm7
f/yUO5RSL1K1cTvAjXSLvDkWRI7YIEyWEVjc73+UUxiqaZpzdj/IYPxOmJiiP5G1
lZBzC5ZZMJRp0y2bELPyHw6KGuiS6BP1iqzg6IeJvp9dtkZParQw5TjEp3jNe12K
uJJCGYaUvd3pqR4WTs1wNfn2olcki65UidQN60wXfSARQ9frc5QzHNtTQnekHUwu
cAkJvj4bCckXsLvXiwE3Ks7erqiQJ0ySNEYWCXF10TfPQwTrMeHxANqTBxjQtDJh
60/SxRXTxsz8SnCDOyQ6nTIkZjNo9mtYw0Bm4Tepnw/bPIKvND7ZiNQLVAAiutKJ
uZv3Ls730lsx3ZTBTpbZXUt/a5MskxQtx4AF2z1ayCeZ3PePnv5OlrgGanAuYJ9K
yhhxsTQPUVQOlzicSM43+5DzF/AYpg//0DrFxLpOS1i/T+kmI6AB6nbQbm//fvP3
uHQ71eYJvfLwYJ/DRq2ypHdKFZN3y4ySYsEWaPvvuJt3BgpNqQh8Du3geSVHLscy
yFkvfMqVloO4GR2RduOeRN6E5Ba03w1zi2pS8q8KdB9JD3XVvxh2dUAzRm9/10CZ
PfJPvWq/96Kj7K8lQTZx+ZOS2P+5Ti7Zv310c/Z9UYb8XP77lFxtdiEMBeXIjE3U
+Ocz805OKFOdBcQ5QDMno6GEZE0RF55Sen9WBczpHQiS18OzOSkFVFYaATWKJa4t
Vm76Aa7WpavX+Xq+KaxlvsjrUO1RaDFN5frZgNnB07Gm191U7DwUvUDqROYmZkxd
MYxlBsvkC+rlPqN2wVwToJMlwRS+/809EUs/oFALZHz9gljMkdDiVCk+D2HjO6NY
nTD3+aIG+8sYTnVOEVFq91DwBu8dmimcnrLEI9In2EIkQZGHmRG1NLmB60SFmYhn
Zsc7lP70/N2QiSIzt1i1WsUOsZx8d8ll5wYmP45en5IEkTByFwPAphGw/Q1JcxDb
zJvRB6bftRkUM0952LGtT3BJiXELSMNgFixSrk2tgTTrR6ka9RWbxpsOpqNtyfT9
DJ/wQ2reFVgR122R3hV21cBEN186X+DmjcWwjb0ifj5S8oRPAJdhxFImff24TRhM
Ny20X6pDW/8IDFGzQETYLWQqj5ruhi5n04hPWzP1auVcUx8KC9huq9xAF/XwIZX0
bnPU/mK6v6RL2LSdA/QMYrUx/BmTp7r4xUztxnGmhJHC2qO4y4PCA8yMY/1tpkrb
exrbCtWVx+RNOzDseH5cfh7Feh3od+NXztKC3W7X/fqhrV9mU1P26qZRAdUZZdgZ
iuoVhxFSeKmGb0XrEtGPcO6jQhVO681UVfZkRhtzN2Cg5PkwxC0iaBTnQZ4rEm1e
aO8sKT0z4+yyhNv/Gi2xW5UsNyC6vzBlvT6OqbHpLQkcmFVBZJ7H4T8XJvMwExMo
iuea5M6q/vkULALX4Aavld6tQ8vnUHlSW5Pf+q8qzfDsw50VfetVXvut7g90Sfv9
4kzaEwl5QTlcFFoRPn7rBXtZ1y/yo5F00a8ehVeULNG0ARMCvNzTtYOTbhV8Q9bx
9j7yZYfEQy6P0XaaC1i7K/PzOdYg7Vsp2WMJr7/yCbWa1HHAFVXN7ho3RmwDc55M
3cc/aYabnfUAiCdvmqddCWHPk+qy1IZAzHi5LGjkuILd2WLmUliA1PC/ldBhTzdO
PrGqFUhp4gaSp1GN3r+rOoaxoSM1xze3MIF+2pGnY1Vr6e1nAPptNZ0HGK0X2u+K
bZUi0rMbbZTOs4H+iqd7FoZWnxcbnj14DLTvJdc684WG9VfL9uI2SOIV8oILxbjg
TK6rZaHpII3BsMfn+cQlqSP6rsI9U2krX9+yNBwf6AxdYaUhGjsGR/peWfh1PQJe
eJ9L3j8jVuGvMBl/wukKwY7cMXfCm+k7PVc/+4GaaMUMO0C0hqn8QUKoyAO3gNGw
UE1ciLSE5an1DXg7Y+7v+H6Z54B82iFImcQeAT7qeIAkHm2fPM5ayQCvgdAnJth5
9NDjRfrIowJEz53DhSBhfaTnHxBVTjgrYdaWXAaX6q4r5gh4YZflW7PqxO4OQFwz
ntNdn5/LDlXIxl9qrI+9j1LO6AgyaBAlgTYzl2no22qAnFwNZebil1lwtAKM/UlX
SIjimFwrMp0oDd0dIeebE7XA1gbkF8z4noMXLlDXGZrRjFGYF3Xp175741QKth6R
XHCG0Hv7n5P/T9j7OeN/Lzq3Ua/aDfCcN0m/8WpXuzSRiUBOQdBpw2vehFraYGi7
TVLGzZIjVGY7WLUIlf/h6UI7XZgpQw5bb8dC/khwNC6R1vRHIKiZlGnQOuE79ASw
nU2pfdNgZA/MXp5+PPUFBnZz/huSMOKZmRSOwILPsTUJn748RyuwRbzNDSoZ8nZd
qhYQQSURaR83HR0rkmzlxQslK78fuDxduUfeYGHvKU+/kRpEb282ilJv2yx3OZ6s
qHQgeW1glBZjfAh8ug/1biaPv/VmPMHplpmckPwDkym7RmgH+zm/o9iFDdPou6xv
WBQKhVIUGf/g80sopO/+j5V2jGuApWawac8DrV+p46ah+16myy0xY/cBfDMtCquk
rtr0V3Y73/8FD70LayG/9BxVBBeud/w5gcpWMza+gNLppIUI/Z8PuESo+/bqWXGc
mrWtCxI5H4T8sepkgk77TCoqGFNBxW1lECRZaaqIYSKDhDwarsH09i0LbP2ZmRXM
6KyjB7yzYsg8kC/hI97lz6MDs0S24t/Ey8vKZi42jcNLukaMpJNBY1ysI6NDBD8r
WGwe+iJyB2jgO924PS+vjiVAHKnFmZMsiK7OBGKhOElXQGKi8VKUSTrfyyTXZKxE
J+6hlCbrd1LFJ684oRTj8lhlJr+V9ZO517DXWkUSvp9LMYsVDP0H/J551LJxEhTn
G2RzF8T7tdUjZim0urN0gm6o9FN97TC6wDODtoMOFLfsz2Oy8KxKPrc3A+g+XTgv
/XfAFzhWFtj5OqHmEgbcaSc+u6DkHDLMde23Ljz0+5fvBWsNdNvun0hZSmiCHw/3
EHj754aePQmoDEMH5SlWjVZNw40AbUQ5CIMutOe1fTnYzrdoFtMkx5JeqYtIvB+e
CzNOUmIt7QxpLgdtHKinK2L5s4H7vXOwT/wCzF2rRpVCQvehz73GpF6Xv+BFdAEu
dDOg8AZO7hhsDHzOvalFGo8fpT5N6GkkpWRDS9WtrRG2EK5ssZthAqO4QLVo5oXI
//uS4tC0IuFzTZMcqZiwDY0tTULgimPg5QMHSr/Db9GC76AkWGFMZZmWqi2jbSms
YdqIA0dREmDY8eiXVTejANF1c0i2rHCZ8/dvphtPIB2WP/K91430wJVGMn8LjaPx
h6Mi5idOGY+mA3hjFh9VNKDRtLMOc/kAa4cHaIyYEiI4HXKtx9hGd6HW83G2nRwR
xei0OY3tW76y90TYvIBi9CbLXsh+9xF3MyXJAetUrCxuDjeR8nC+u1BFOK9SDfyw
LOke1cjNYygo4ZTLNx2UMUYSzveIW5HzWT9q3en5g8ZJOPetE3+igI9mzBeqwVxW
Lmt5In2iPExdz7ikLXBhRxzfHjrdZtv8xJuJpScpg/uPAJs24fUVgtFeUG67sIi8
R4gkUe6iKNbXaYVxhYqHysXGyzhUbllcH7dI+7SMrHta0spkvekAHxfqxEQfIo4c
3uaHBDZ2VObeft/lIUZM5zwiBea2AjuuScBdjEBtBTtBYrWmjkRepp5q4nSskVaB
JbfQRQ/scoyY1WiG/5bSEI7S/kPPw/hNA7hTnALVO5Bs3WOXpIbknWp9tUlhHJv1
3rvBeytHLTTcZJSRRJgkyVD3pyx7zDRfacc7w77QxmwTkld2lVn3bRSUu7rPOnhj
4TRQN5ZHelMUvQAp/kqWxNOPX1UxCnBCuXNvbprSXYjs9CTztygH1okXGEQRt7Py
rS+H6vRvZsIfSyZDmDX9MxDimrwNdAdHfDAVJtc4BsmHrzZhaohVe8o0Xeckg7pi
koTKl+QPFlWFp9XxvlN1mpiFj/XVcwkdrDmG7OjS28l00cwP4QYOTeLW9z86nvrT
8lWsfi87l9qhmZLntRAfpM+wDwK0qyFi1E0u/7CFI3yuSEqkODyCPjhOxRhJioxK
ZU8T7Udt5wbsEs5ACCBU+BYP7ANZaJeP5F07UY9Q8CUbdOwMABCTHSdADB9JYbG1
VrQJtKRcWFIxKDQ21aqRZXxstICyhS8OSGmyzMMsuOSgeo3wajYFw3PQCFPUN8Fz
jQygJ4Wt2UFXbUlsxghWa2f6wys3FxYUas4ZvU0zZRqvOoz8v6aK89IJTBRxzDpJ
grwX84W1qtOPnfffi9Won0OK+47skrLgKNOJvEW5w7CL0adL/nHGHgxs3i4icUX2
j8OACT4VTW9OKJwfRpDFJCHroc2vIXiTzUvOUyvyQ/KCKvHh/7laDhXibLXagHU9
bq/HXeBDJuf1lC4FfN4A3xVj87c9tvCtxikkYbsI27a+S/eGt5WZc7T6nLAtB26i
U2MRESXUgXhHxexJmmHNLBA6e8k+k4T7umuQAj3MGNcQbTrMzGEuBfVAMzbal7iX
yvqsG97U12epT/WsHIgHOqw6zOepD8obsCSe9vCiHsehg0Mpu4HMrVYRlD23D+Tk
0m6Otw0x1LMmnmx+aUw+wUgaqKeV+Jz6hLoqDIAwtlLoR8lyK3VbXqgKVuOeURR/
YbJy8HfBp1ey/aXT2aTDmlGRQXRbTOTi6ogzm5jW+OadjjAqcNR71k8aY7dQCvVW
lkZqZjjy0nBujr6mPlGPQTLgyBkud0Obx79UZCyzsIr+DUMXwwkttcmUnfhRHiNE
NWjxueDtECp39cgCiABfhDCJvQbBAe56LCuTFEwn2HVJqI3rC7Dd2q6kD5Fpobmx
LVcVniEpBRfFjLpMjcRVOZZV5G3MqzhYPv96Kx1NVEOSi0bToFSdnYXhYrxPtYqO
MsdEjw2gj5wQ748WDjIOnmuLDePes8D2zpZZjQSassiD4O/jxUTtGTSkSH0MjY6D
D6+iQNamNVvZwl1gUAvBUr5ukH0DJaBSvw2iLVFn9isoECiDloRueM3nfnOfRtKQ
CbWU+IDQG5wOhjnmhBMMmzd2ruV+zKRUvoXEHDWKkPRaSEKcz0OSZ/V/oiukqiYp
voL3gywGg9+b4o52vmkHB2hHjeLZcIfGpuDTGHEDWwJy2fGw7Ea3P2PNvsZ3dUCl
Bw5dunv0HyPGmSwfukp3sziPZr6DLzhA3PQ9Y6Jzx3Z7kDTs1s1ayiFVXEtbXHD1
dQKNYw3qVKdM5VCZgo9yyDbiWkDMPnUIteyGvLlmZsMCoQ0dFdlazPt9nEDJY2MM
pfL795p/hWhUW2UptswdIo18kR8OoFC043gXyNt9Yg0P940NdFQKbtyGRxIT+pLl
EYe+Vof5U7waDaNmDpjxErnsSIEggn/r4VPKzJh5FTPAvaifaNRssm9PgJ+Hj9x0
BAACwcbFYexfEnNWrfq7i5lTmqdYnFSG0rpIlYxOAOoONuMCiIDdD2BYBgdlHtS+
6U150IE13KZm0EU2N8uknhAtAaQvGwB5CpUtH8N26nyYYb0VrPy1XbrBlRpab/2f
cwsvuvcxbQzY2tG3T+trmVeoHdjoSW43zaLokC38XBwjHno5/PrBjPmC0Q+guhSJ
BDt0J8rsHi1f8o22syCM58X91ntYJ3gakH9s8AqEvP7FhTcAginjIR87Uq0CK448
7J+eHU3pVAqXpbJOIzZW8RfAj/HW3/AMGFsbjAlhWIIdxKSePu0xMlxxykb+Otaw
wXb/mdAL68aR6wL0qmvQhF6retYQoTIT8PtcG9v6ZyWgYs6xGq6iUHRb8eeTnmSs
Q5PF2OtjUGuBz4wdj+sjKAtjnlrXPhSJSc1j7KXwlbbTT107utc5I4y3ikDWvdU9
vzMqt9ZqCN2Aitus3sZpDspbwy7nk22aSdPqk3N0uH9DJjTqwZJTlT4ConqdHONC
00DBhIgjJQoTPwMEKssztdCG37p1wS6VjY0vP4HzBwlzujN+cEpewPvAscuHrd+8
DpAjVKQ9szgPhjzxmLW0dlh4eGqj2FnmPI0xt467BWC63jOAoSdh17sq88HjeS6U
lFx5nHqC6iWDlHl1ZK8T/RlVRoiy/iZvwgXS9M2NJ9FDI7k01xCj5z1ZDkNgCpik
wa/SsA5G77P7OD5SrZI/AlXG1BRB/cmZKq2/85ntlINojg13fD8pQRL1onhnrWvM
ss0uGvF+ZCKi6y/Ua9+lFXQRO0DP/dXQ0W7agISlrxMhZnUSJkvwXNL5N5Bnd4/U
f5c6isU/+mEcK8FhLdq9hLmCmsDfIQxNE1IfbVYLjvjjaX7w7ggHAnNi37/P7d0b
4GxF2XPu7J1N+cxmyFTO/KRzKkuey0zJvgLxqGc0cW5JBrsZW0btZ69A+ppkJUzt
5nr0/6oiBXps+Dsl4anQ4Nxc1lFewfmIb8I2POHKD10KW/KkUZ6zNFgEhwFzE248
GrsFkPSWH4WSIbxLydQ41hYJhhM9EuGhAlssmYLI1JIDeOf85pzCoCj146GjA5hK
ZL9YJoM2YpwBWzxFKLVdu5f63weIgQIS0mgkgDfieHKd0NYFaQCoo29KWwoBVFai
qKP+5nFBDSVjLla8TqryRc+ZoU5COS97BFPzRe1S7m0gVIPUpRF+oTZQbvSIIcBz
TPZWdaNiPw7dI/wEqtDBKcR64tWADIuNqEfdi+75diJpcpUT2wRU5Lo/VcoiPd9H
vx12xMSqDM0kaLO5zAk9Rwq2ZxxhpxLwlmGzj/E3GpffW8k2uWok/CCGCvcNzsBF
HdvP5E04vLz9BPcjRXk/QJ07qry6aykjVP1TlDH2xp1dsaqbuBPo1i8UW4iQB3yG
mEZF6LFiReHwLx5Kh2S2/Q6hGs7TmtYkn30iRF9V+5AJcbIrpklKs2pGl7N+jObY
uOu3WUf6Wyjbf7HQ2JMbaZIEhXD96oaWucvJ1wXG1ulfQ1pXblL1LePWdYziuSqo
CrcVegC1I7a+kfOt59t+58yaEMxN3GYsxlC3pOkvdDdT5nLM0jsx81cjkDqzbHOB
ExegwH3diSSZX8cObpZgTWdGcC9KSgchZqZ+wnQeQjmiD6418JzZ0ragt8A3YsnZ
wPye8oDTPM8fV4XqDEaxi+KcUEwk+k7KW5xwOp0W+I7hvIbE1xQ+aIwCvuBUxIaT
6OzrHf1sPEaQmEFaFoTzsbTjVz70wUkxJVrAR3nPssLk9eMksbuet1IcoY/i1c5b
Frvvhq1TxNZw5JJ0kxbZcH+Pbjt/+35YJKLtKzE1mUGHzTD+ygV8m+ovlFqzgPKD
mqajwapXupWHgflHXseIQg+TJBRabLWGD7mq/FHiby68ScGmyFGqnbFj1It5H/Ka
wJSGcW7bjG+qIDFnIO0teVddUTIvEDT16UUXrjdbxJYGu174nkmDKEn3bm0xkvc1
r1M7dAPNk/AosSLOO60+Rqu64uSf0gbRCdJzzLAmC7Bkk/TB/KdEJ/bjsCsempmO
MOFUiWKAcetJ9YTWebo1dxD7cCpdsot2spmXhhV3uR5jRMKsuNqqUI+4r168R+JH
8gt3e9jFgYEzxdiLpwpKe6SLE0fO2UqiazQSaHO9rAnYZaHFLxDTwi5ftmdXnqxr
Y8cyGL//uKGsay/286Qe/0WnJjZmthdpQqq3ZLpgtYaxmdFzXqX9BGrysz2bCwSI
+QudaHCyXaaRm0YdJ/b6LAfFhtZltZsiu0/Q2II6Lk8xLZUN5QzeRluf/bBQHZjz
gINUvdNM3scbYfVH8xiJWtI430rBuBLbv1vFyW5J6GpjFn3f3T1q7mqyFepphDXG
FrhRgiSLiQMYfailBslhBbH8b9myaQZIGR2YnR0TmAyrFkkroqasqVC3Cw3afr6w
PGEGvpcCE8bJSxzdDbahehPngDv5pURCLgWilbvhaYeuG+mxX4G0B9trW3u6sgif
ZVllrCx618T+V6LgaIY0P3X21gPvZBbQzAlPKzG+bYTH94pttTC5WRYbYVLwp65z
75fikwX1hWIpCwWClIEzyIyIRC7K1nq2+gOMUXifrF0F5694XrbmeLvNWHfvPg6W
4+QDh7DUNeX80mhyBpxZASPDNXPSXAS7Qk8c1LpmGVPUZRxvZ2OO9hFYYo2KccyZ
AAk22pgiPJHcc9vZ8h/Z7YgcU3GPv7naOpHCQ361nBOjS/0mhysamggXXGBFQQSC
Qt+JaINjqJYk5cQFy79FpJQPSCYzcJEsLKdONLQ41yLNj0EjS+zdBQVg9B6r4Hs+
7QpXcyukjFmc/JRZMbqXAjlyCjSvAI9sEwRyNBS5XdMcjYR5UT4BQP4zsT+sDpmY
WOUxyLfl3ZI1ao7nOAIoaVoKUnqS4+RzsvFMRMHmL6Zq70nNo3V+w2bsDkU0xuuA
nEj3F3FUvZNDktVbiP7Y/N39A5J9HJAZNXY90DRJY+5ETeBs1qxiUmNc5v+JWrQV
SpzPwi2+U+9bvnphnU0ipJM2r5N55udIpUEce317yeBsTJ9iKquyigrZAO3EIbjd
psiR8lxwg9lcdJjxTc+mb1jkh37oIXjPdCysjnYQ5suQSNxLxW1RwU+uqSpSj5Ls
7qCNHcHU/HsDBhcXYlviI81b0AAHF2OagvtqOylOsBbgfMW4/0+CF5iVEUrAFGdO
wUaPSfLuZB0VnG3ZrCg0ckBRyLVDpR761T9CwZTmPgeouVY9oOXkMSxD1uzFlBIM
M76jp67BmM8s2uz99/VJDMTXDLyWVvmWSIfI8zw59cGKsQSkG3oR7vMul/RpzJ5Z
mdTyV+k64AnslH35Nwn6jJvkguVT/QJgv52Mx4KJQG0ECUH/aW1DcmIYozpeZnOV
Jvh8B3tPWz7mF51aUh9AoSFoqbemspbs36FuycOhMrrs7xvIH2khe95KwgaRqLtm
nhA4IpqyJZ1jHy2LEQx9XY4tFPKD2Jn9fnJEErP/eJCF5JlRbBf7miMt+s1AZloS
kQd40vsYeFVQ5WUJta8p3GjAhYfCeHOcTIUzaRuqjqbhF75oEGmWSOVNMNMH8BEW
6qiUloO7EJfjGYUH8/9g9Uy4py+RoNJjwRqcdz7iNooqzWHVXY8f3QoDHoMXrqPq
bPpehlIDRQNbkpvmqb6VhPYfBNusfeph6Q5Bwc5gKeNbiufyMtvc8vBUHZp395pE
uPJ9DmmJacOLTSpaVXg0I9qHNNg+gwV19OKeUwbsFHY8QIYSSuzr4MMkx0hb+fky
yq6W5SHI4/9KazSEznZmFO1bAuR5LXB/eDCbqC1BnOnZm9jKgDdz1cmcIamzMUVy
L/SXBYSu0vHo+Rx0IOICV4d5lp/y4iDQFL+MbtAb5Tilt6gMN9A99JNcCIkRCTEi
v+m/wwdt5hcVeLO3tlBD8FbmHpZIX00QmZLw85cYKfogIIIucavadojsKkCYrwzW
5IZrpbvfzzzWHIgOvOhbDly3VAPuzzyeFSBGPJ6ePXI1VJxKY9l/fko3S2jkTUIJ
bzK/PatVLgWGFnn5+5EmEkSRXTtknDxLyWK+wth93qK02gEW6REQfvBsBESL6SHM
YBsI6TIDW9rj368Oqp5aoZfCfny9DCEaJXTR/0thid1hoXX/JMZBPy6VuYbFnIT2
PJzZjzajbo+Xf5FjiKuU3fhIK3IDI7Qq6eW4M/K4GtmG5EHb53MFAQeYoCBCh5o9
fB229/Yj+uLNDo4hNVf+HnHpIjxgpTqDcKU0GLeecOATpJz95abGr2W/xfxz0EQf
N3vSNBNyxRxu58oY97yQYnE1XDCASufc/iJmh2aTCPxRH1zx0nXqMGywd6ZaHTCw
TPzGMirskfD5pG8YdwO5qGmISBx86nMdyCFRQWoC2aaXnUXUDTsmTwmXoeQYwPTP
KDcMgY/kXJB5PWOrvmKiWUDhNFwVVu+xLHz/nvcX8yC4t5yBiDBiBPk/h9+huWHE
lTv4wTmOJ+Qf8r5ehexaEMhIpc6yqjnFPrCtvGyU1l+edezgN8+oycuB59yzWpQu
pGFg/Wz13mLJGo7LN+YRoE7t8pRlwK5w1n9IuF1i+/V+XbxEbnVjqucD+PM803uZ
B7Xg+lK7Tiuq5ziW/Gp36iQQJziXc8nBGlMEAEZcg/WSdSYJ+lYah8Wy2X8//P1q
VPY1n5IDWWlLAdK4gC1J40FaRqyXqI20+GrI1ITmxlvefUEDruWrggW+vQGnEWRW
SJI9bz0TAFeUay6R0j7lrMIt9G4mPA5n5LPwI3rvsWiD6mON32GiLNTOwplwK1wY
o92DyY08LoOl/9NyFEEkBW8xJYZA10U8fqizjq+zId/genAUmlyPUUOp0PQMV9Mq
Z+oCVgPKZBfO85aANxgtujvnOfDgMsqIM9gu7OOkzQ5MyTd7oAdjEgqZp9Z2k5DB
58L2PgKCGnO3z99te98Vf6FsuBrzzVx0b2OJCysovGJmfNK0fLSpy+f1E65FA7ja
0/mUKHaXUuypFDQioE5dW5GU3Fyc2noXk4PNE88Y32ns+hbRmk/BxiWs13FAm5UF
CGmjWmyVpPXHbPbcaXeTrqPSrtm7YlmNH+/Wm2t2YQxOz0fEK4qRyQ6IjjDnN/hC
5UhUCH1V1cjfB4KC1zpHVf8+BXmSqri1Dr4v8H1vztKcX7fNQyZv/YfTtxe7ZLCE
TVYXnfS0t18bhKxKVAoxIXSyoyLQe5S4LQNBu5pXuuKpPkk44b3KQEfqvJh133Ze
At9AIvLyP5gaI++8XgyIZz9tMY3VUkv2x+ux6ChLu2/WRJoLRxklghQD8y+IbaMl
tubttkNIlYVCtuh4dsbg3di0z5lQ/0ze+PzR9xq81dbiHuTmO4SpD7TXqbKfCj3Y
Sz+CPbq+sAtweqwKbVHV1DwoNLEweQA+enWrhtSTyn7glmu8HDTSTt68DD1tR+4S
lEEIxlPJpcdkO6suQ4nMB9o3W4z5fvE0bSgA8pUfkExN6GsnI0fL/aJUoZqmTz2L
yYJLPNfjHEi9lhLUDUOmWBTihVjW66ujZg0GyhOFTDXJNAw3B5EsukFScY7xKOZc
ztCRQc1qwjoJ/bezmnpfAsFR/ByXyYf9FIr0045FboHNZJr/VpDcbVPENJnGor6v
3KlAmR23TWf087TwRd6DQeBKSHdp5pAYMHqJdQ0vklWX/L+nDeQsCrCVcMJNksZp
bqzR0Nk/9MCAtTcCS/6G3yfGpG/TEKUhxA4RWiuFldSZox51GlYUMlx1D0ALz2zZ
8udoMzb+7QcupB5OybuUxNRH5OhG6FMf2Kd78O5vmjkmm1RqK0xcUTz/wh+NlDSM
4y2vUo4T75ZNC+pNM/uCF4mFIsQPOIfI0qRr6iVL6qL4lJhbid78eyrJSzW5lyMw
WAEatsQMab5p+IAVWi0WYC2ihea1SHlPjfe3qMko7PoRPoTbD56s3ZgsuRzcShCC
we3ikxWCc3ML0r06Qi0MlnnkZ0dzorMShnNFEv2VL6vUXmtZGS7hVtVgAzJnnDqW
HaKKnJMKTUT8Px9caM+2ZSmKXEgjTXHkfoBHZdDEChnhlzqukxWba5c4sqTwi/Bw
eS0+y6W+dEF+bMRsMAmb+SJJFoX8FFYxrltd79NZ5+UOWIRagAlhaKEmSrRMmKz/
6C8OtOV9oOmgKbg/x8k7iQMtlwubmdnuqHBGpIvB4fmBithALfxm24AYZjody1+L
NRvg1B+4KA8t7E/x/IVRsymBMq6zvl/8Y/MlCxFid8Msf4aD+5UIcsmBlhDfcQgO
RU/mQRcMFz1HeO2aaKQpssQR702rIi6w4ikEU+rjrayB5yD9BKZfPUenSMa0XWfS
22FXOiKHKgX8gnhq3qQ7JOQiwz1WMUZqJc9fOZfWiILMup4RRbnHjGbPYpkhhOeI
YuBvK+RFyOdciMpKdKrS7MfBejndLz4gWQBxl9V3oIHrBCyBXA4ElgerqRYr2e4O
FnnlDJA6WIfFgtJpKotlnn0VP2U5DvCnuTidXSFJWK2jJ/+KV/N3+rgfMOeT0/h4
fLqm2s/2eIjIRCCuuE3JRFfmYn6tzfYd3cmI99vFGrSJt4VkGoQYtWhdgONYxh1L
E0f3FAnaiMR9GFKf4vPUGXxufrj4PH91QB7TPIKlrtG3c4HzocQJVbcUr7gkLgnl
dO2tu9vlE83Ar/KXJOji7sLHjjZRmKdo/9YoLkrZDFwfRqHCW3FmiebqyIQeRVrt
BQtULvN5qMuyNQ/CgjB9rTCuFzASQlFIafUQyogiixLR/4DHUXIjr86SOIiZh5ID
vh1+yFR7/Cln3p+lJtRfZnUd4GE1vgY4+L92GZR2qDxS8Laa0auW50q6zNReQpA6
yDOA4KnsTf513IT1+Vip4d/zbktNLfA3H7iQY0J/HGPIvZVamGi9Qa2Zm68Goju9
EesRE0ErpxMRDvuFcygltxdv3+gjDqY31R3LggMoTpqw4ypglidqfHfXvPZw1Y8q
Zj3IYJ7nysjah5EOpOr7bdlW6aOekdpzjE+3Y78GrJRFGaj15o5KCfvU6atK9Vic
HmmVqMKvxnLk4aY6gKmcReT6GZ0oHsSUu4XPiuR9nDBMPBtg+QEZEo1C1oro1iAu
hNfv8yoiW/FgQS5N8fad8ZeOQnNk/1hNa8fEreNp68w8myf9EB9iMA9RwoqsOW3x
koxfGyTdjFTzLaFq94+lKT8C5NJKRLn/wUdz/dOb1tIpv8DUq6IuHwiWQypDNxpu
KCWtN+fEcnHAwJJg2fnUbdZzVDQ+BbsLODANfyB0R0LpaFwDvITkkJAbfu5UFPNE
ouM/XPJF7aFqtRkcOrpPIcVINdJeN2aG2Mj1yYVSi0eYiSExD16rTzCQYHQ52TKs
Ec1cwWB432Lzq96FfB+4jMY5ZWYB/amkP4lLi30c5dVn6MxkmRSKEXFRPIu1gspP
QQwb6R1lOTqparaYSiuTmeuOSO1cLG2xZeLEqfxodWBcNW5GtcfjzoPFW+MDEGZF
tI0NAGePWc6JYN8sY82BoRtTBEnCCq5Vat2z+1djrC3mSBGowvZLbAUjA09jVZn8
jVjMWDOLRaanptkxXn3VhVmppRET5qyXmfNKDuAVjSvSif2yy79S7WYHV5W8ViH+
E+XYjxoleW34EHNonTO/Md9tBoLxMnZv3kkehvmjhliSmH/8MuNtfttJ7wSgsU+T
BOg2s7NgDwke6i+TxDYzdnxiru30LrYqm1CWPDehcDl5TnAhNMRBjWb483dBcQKI
zgH2FakfWxmrG1vcByfE+EMW4qc4jKjyzyu1/PUbpE4NhO8YjKebR6g7kYv2Ry6P
BOypzaJ9oHWNPu+3ygPPND+gW70sgC3/khPb/HtBrn0DHjOUDLlYAauB4HVlOxqo
DRMonC3+c0/BFBtS7AJ+h0hkA5zD3jZahlTvNa/6b6coudUDxfkpuO9ajPnk/E6B
Me4ahmOkqZLgNhEa2zUmWUNWv3rH5u9yuAKkeKcuWamdC3Yyvm1VAMS8CYypi9LC
YrgM13aQ2cAME2OUlyxYloqQvgmSCnpgHJ5YGFQDfavN3bvKCaifHKEHKOYDqy/n
C4J+EK52OwKMKSkremVIBvLLOhhX6KeLqKe/U2bOWANTo7t+nDz6MDisc3aUfPuK
XtkbvkP2aveUtH+F3c58dl2REpuSm2eNnnBxrn3npeDgIo+uuj5FCQmIqWeig5EB
GMv3oC1KAX6lhu6hj5VHxArkCYwBvTZ2gW7x8jr6khbEmVwm6BwJbF3c1pfVyl4y
eYChvRblITvr/D+JdICK2JTSMs0UtBWeZSSXIKyWR4dsoWZ1TryO7SNBCk30Q1BZ
JNvWiAzj7jB2M/TCxVRF/ahqKQWecfZrBShrp69kzG3xkmqA4N4PtR2VW8t7rrf+
4OiIdgOxkMMyhcDU8ldiKcgDTo2XVx+Gv4YwKznlhwzjb3gN8zI/O/HtcsqrpewJ
QuR680dmZ1b2kbUloQk5jjmCzD9HQSZdKtleQk2Dviv/3Sq0gGsgo0WfuaxKwEeC
`protect END_PROTECTED
