`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ke6zdPkNyTc7ZBYQ+zskhWsnWWZijEkEIf1eGTX/QVDDpLALRk3wurAjqTKYNBmP
pffQRDGXmuEegSRVCSZ49Q9PiUvKQsI8x91d2HxIbm24xgkAV+ASc56qeLh6WjOr
6g9DpcI/GJfYHtZ1wnlyxPEbbM/UZcGKDSXYjMOnxNq1wty5+zPxUaQbPqeBmdGn
8yZJXdCrTi1m3dxLx6/iqgycQoIPDwRD/9wLTumdR7nUK9z/5Ey1cBYRhl9/1jJl
+s/sfu0/jEn6HmP0aNe87CAG3hlw4Ix650VryvTqtI2Eka6BXERw7trKxWrutMPQ
D+cTUOVeGHs0mNFGLAcz8cu4ZRlO+jzpL0cNoiLDvgcmMaFQ2AIWJdbMzENTbPzm
N3ms6dnmM7JEBTEZhTEIapyvIQmt7uTFp7sUmSW0lBZjK+wvUAAy6y82jKmbwkS7
xDwc3ZkcFG3kpDoIbq1MMpft4/abdRK//IPAWe39wemT6XXrFq8MpkdBj/fm2Eft
r4Pvuw/XN5gOV+DZyiy1ANiuyqo+EXs27WUI43fvr7qPnA5YZRgBnmUN+xu+qYcd
RYvyDo1AeJKYg+AIxiI172IgVS0iELe8U7SLJ5KFcoJZ9guQx8wQWtlaFLp4oz85
+gEPthSVHtpo5Px+HmwAKXBzZ1+FzdXp13pg82JBbjsuFr/UQmSMDWkipXniOxmu
4Qn73WPAc9hcpUz6r0pugeN7tdEYyHirFEwAxy/w0NzcRqBifVeJj8DFPEroGm8f
qS3pAfMgyGs90tJ/L4Zz1qAy4fAycyhEOw3e6Ffpt0lFfiU/IxwAkKz7FvwA5rkm
WUInyM9J95ah5hjoG+su7GZz5HKJZq+jE9AXYrz8Lj/EoeTdkAU87YxHG6tiD5GN
XekiEKn4uD4F1TZFNpYdV+QYBpLU/hZB/piOUpo7D1Sz9VnhEsTG1TQQf6QOARhz
SpO1sLKd0krZgPadUpyGrHVmsLmWA8wzu5ead999mEeubukvytfa2DnIhy41eaKo
sd3hqpcfYdkBBv+QmA8o4O0TBNEVUIw5qPkg2lOP/R9eUEINIhyeXPmzZPCd1SmD
XvIsbwRBKMS2HEhZLDUBtEjhsj6wbotAIaAeCdclpqHpKMjV04xkNtZJVQ2TkZn3
SZ9LQeBbIKo+q9/Fs8zOcQhnWR406mFaPKnpZ+RDG2h6yqHkQvhxt77BvaoLm/EQ
MLtHRfRN/SB9x0f1/zVLgR8CzvUSr3saB9BXyG82EudiMO3xly8jJ0gYxbHlkBzB
Rz/sqMewNyC80rTfZrkS03g/QvfxM/YxQCOBv8tPcqZkHVV2n88BzRjBxxdhOxUf
ZEzs+BMFbSECkfbJ/0MQwnFIwrDPabvxvVkneyLiUUIx5FK3ABP6E4RiFkN8odQD
9QHfKlJzZb797FhywlTcIbH0bj5Np81dsZI4pRVCmbYi1+BJTw2BRvpClOLdOyaf
LxzqhgbmvvSqYdUZ+Xf6M2F4PHwdwifcNyoQiG1+sR3lD0RyeUVBIMgm5n2475pp
5aZnfSWu+d5F/QzJFYzG9Z7VgXMs6uaz4kNZGyMz7JlpMR9fbBjv4HgxtMoGyOXW
hApTqVZXDdK7XZbhp7iiyCTa24Y2tg8ffwTEEeE/SlBy/K8at85C5uAIqCzgCEvl
0qH5R7i4nHdxsHX9jsIrRDfDUER1jz0ORJ1QjR8buJ8B/B7ZnYoJH2QU+y2xCuYN
qXUqSYqC+RLgbKfqhIHzN7o2un+TcOkiv/mfJTxWeMGCErXK9WbCpEg8RN9oqkqL
UigkPUkq15htQcYwxsbYo4ZZeMjlxC435cDuWIHd1RQQNKCqDGww1q0qrWJtq1tO
irNdVxuOknAvxpstekYjcBzgw/Oc2qfF6mzVihpWNt6/cPPyuP7oHfvdsId+3Qfw
gxdFj/eDjw2ynztz/uMtu8EpjZCmDjWVddMByfcqt7z6+rA+slH40ZKDSNJASZNI
WKED5HacQFp65iMmUsI/fOUm27rSrLmwPCOORaHltMA1hMa7mxcxtV0IhzRH1jd+
Ojc/rqfYt9Ki+OVxy0QlBCs0NNBBb2r+OfLXs30CdQHraV8K2sPJS5Gx4/h8sOsO
3L3bkJWT5jd5DkG9SC7rATIlK+fxTUG9KRFgMlbk64PKOKQfH6YTMntoVREPja+/
zhEr1i+oZfgrdE0QGWrnFvQG0SJaWp0sbw6ogNcEP9Lique16iknfIIygfj6stGl
8iPyqvgSqQA36JOiXM2q6W+OkGFfVhHfHtDKzCDdWEYZW8hycf0dWaEI/spiIFfJ
NePCQa94O1QgTB9Msy9uEKMzaojvfx1HlVnbKkKZwa7CBBqdTSWWDU2ECEvONLFv
tx805+Kh+MGKbER1UV3VpPl5r9X20NBw7aAJaIsSxJF6JTsmoPKNLnXaiNutSNYw
DV0FWmXR7C2IyuSb7s2X919NyU+N6RgIgjDjTtIllMVilsnAZRtNd4H+8e8UGomJ
PeBjgFi8zStBF9VlMM1f2aviOtIJXEdnMW0ipvDtfUnFXe2i2XwqFWH7xOb8d34f
FKtZ5Xi95Pr6zi28siT0tRCG1Fbf45Ge/w0csO23B1vAyblQYkZar6M+q5kTo8Y2
o6HXzErSJ2/Euf0ffW7mCc7MtoJB7Xq8yGGUt3qadorvPuKL0wjjQKuzItayaZqT
dv853Wnb2uyBDpY/pqWCsVKWq4c7EB6CyZYiIl5ph8HhTNqKnm/ZfNDxs/iC/J9d
AoEIo7KjQQ0/PHUNjW0/orfEjZ1tK5O8DGa8qJxlqP1/MN7UF8kWa6viT7kIu/TE
E0phAEz4HF7yKhMFk0S1hHGoV5nsOCUAPbwDT6loeydcqbPI7q57XZ1GASEsrjKo
BZsHv7aJpcYIpasXyUiV/YreMiOll1zT/4XUW6CfDwBBbXO7G8OVIo0iGL7akzbj
r6KCJNNIiCksDos9vTcAwkaFiIRIK8Me0RzEi5w6UaNLGxXZyx3BejEUexYyojEb
7PY+IZarlQWMt/fDe4CGAA5XcLVOqgCbwvJBfu/qHse9aQJqG1ThKo6oONudIk4c
xcyBo5M4zqXvXyIAPvuUXbmmD46+oeE8FGtGmL1lT4w2kaCVX9ezfD3uEzltwvqD
+OXDz64HAzOUvkMxcaFPlvhusEpJroi6oL8qUxqNtcuoGpWhYzHhYuMYfAjx0P2m
xxuvBDIyl009mWQSFL6o7wC3RGS462f4kAbkdqMEMTdq4jPQh6etqFy8Dbnl6mFI
MuCN1U5rmYVILZmAcb1u4a7Mlo9WCT6j6zSwUMfUJnIzTu0CqrYDw+iIK65VAH9Q
u+IFgNl9I21RZ7vn2qreeypuQkTzjEvXK69LILCilDwa1tg7M2Ns4hUdPxVlEUGP
4kF+wA0XXmPkmR+KQ19QRHvTsynfPWA15sKJ0XicF5Dz7MTz//B9Xmvpn1++J65L
k242rjHF4jP1pBJgQE3HjUoGJttW8KGpsQIeMuMXi2qNmUog+bfiHP7Ro9NJfis1
ef8hnBbQeyEiMzTW0dMerZ+y/XyWLZq7jVfnDM8CcpnO5Vt1GJ2BmcUaEbu1qphh
s010Q98IB9tEWSUSyv0lAN0iP/VjKRoegz/U1wvaT/nLLRrGaY2QgQekI+tJgezK
8l+P5kfsuKX/FLHNUb4QWd9sQzdgc40SP4WYo6gQWlafJyr7KdCklBpwKaVniCoq
e8SeOzem3fJivPB1c7zhi8KWqs9SI6n/FQOpTnVg9XXUW5LwFl4EpIRgwRVCGH2J
NMoMTXXdWHMlRPhM2GJUwbF1RB9hl766oM7Aoj4IK3/xjuH4XWP9YUjwScxHyMYS
GC7ig0N4V8wCbqVD7NN9HCd3neEcHAygDEBKOrloY4nD+kBDcwPZ09mNzMs4heKQ
KUIXCo+zpn4mtDlWG1alEls647VQQ9sMfia+TyNx5RVbt4jRxfpzuKsHPiuA/gMJ
UxaHGi7gVRMy4tQDOLPf5KyUcslPFSjElspOV9kUP66PfW/cD54c3ZkAtjaHNUyw
+RQiJBN/EVkjbI5MIIehH6VqY6QLMvQMlUt5eR197/h2aookUMjHKAT8YIZddFj/
+rxSDP3G75ikSihrPOcB1q6KOqclB1T7UPIrDzinB7YNxfbqBRW+wpvAgBJDbWAe
KDb1Quqp/XbAu677oM24qf4nGzQmlpbneRrlBc4TH8wpTA5Sijl++mj/11qJ2IC0
sPYg+pBpqYARXaMRbJUnEBxF4TbL/VDC0Y3i3ylMCzShhABSt+OYS2uMhbn95hye
+KAFtCkA745gGwRMHvD/OXaiUb2Il9SW2O8BrG1PZRZApYxqyR+7lGeCSFlk5yNt
f8A324660X6/4QLxrExelc8su/2gJxd5nAbZttSXQslownOeMNRThffupVfM4cTK
M83RyuHjuFkFR5LXDDckZNoYoJQhhUad3vl5YoTItWTFbJF75Vv/3dPcsUxBVD8L
H9wg5KYssLH9GXwqSMlZPBvJv1RHJPIoFTcy3Sc8/5Sm6Et30GnjqbCocokcuDcI
+xgiKHao3pzhLHXgYVDcU7/9Ubjmg1VOiDscZS1R/ABcCl9amWjijsWERBYsN0F/
9CZrevuGVwbCK1BHXrD1VcN4U6k5rwUlMZQrPnsr01JhcNxIe0Ti7Zq0wue0OfZ+
BQz5jE02m2f3QGyiQhrdke+w5iuyPYAM4Oam9ODLNdWaADkZh9R9CBG6h7IXIGUJ
yCTXjxqemHBDdfl2CD2Hq3NGmSd9IjCMxVjfsQ06vArwjsbZfmYArNDs+zq976u9
DauC9sWtxo+SPB8nOSO/8DyNbMSJiD+MAw9pdhqrAnZSIh7xsacqZ+o9J+1zjRQj
MjHUDt0UDqSgnKjEjaP2Wm2rIuexcPjTpjymp+IX8TljO26znKdRAG9aYBnU8TeP
qpefwnG3Lh2Ueur6uD9zm8ljJcwny3IUDQbT0qMievQRLfY8qcYlbgj4b1hSK56X
9JTmZEXhatU7+13gumz1sIc4ag5EIr/rejIfXJkCaD8Vm/J04yrHWhtgRiJ/xsxF
LXaxqH0tHgcsjGYuiHiLX6z8Y6O7J51+A0BB32a5OwYtcN2XszOvU6Nrh/K6vn3y
yqNKuqz1vs7b5ciEzj7aViausF8IF81yb8HQXfnaftnHTGznzr8y7mD6gS4Vx4fj
xz11Ajx6eEYiIgfCpufHvzwkEZps58BgxgaesZOzasw77F7R0KPVX9VeMlSmSnF8
IUMMEmVvIRz5GjXEV7uGjwAQs8eYu1gSj8+y7qykVvbDX1tn25SE7vC9bHtbca3g
opLFiBx2D/NEtec8msoj5Hfw+kMnnkkbBGh4r3AfZMtygtJ9Jvcqz0tR+euW7s2J
US9UaNxrtSb5U5XQiBNPH6n97VxllLNMWCDypmVuFjurUDXU+44wfkbhE4aBJ0g/
MnqF05mdY3p/nE0z/GzlGSH0Pu4f4sDwTPGH2LsjfqD57IjsofNZwB7nNAn/76KJ
i/CIZAwp/s9HZThK6nCAy7iIFlEQGRekqJCg3g+2J7M2GY0OfzNVZsmDIYOn/fVR
T9IQfELS3KTp9X9g2OnsiAIyO6zefXKVbIH2ATKeO3wkOJFtz2bB/PRPS21Jwf1X
2uIhiiCzs+ccQLPd1g19L2VhBHotAxFChs8Vfpl+jYmEeTgEDquYy9ECF0UAwym9
5BkMmtUUhcBXfTvBIzFcKsWEjfPL4IMzADxDOeGLQCFfgQsOvnOcW1sFPkWtBvO8
0P6JYgARAltcs3wmjrc3QqFJaeBbaCrSmO+VppiOgVU8lXyiIwhr6CzpkjVb3kpz
ixqACWfkjZcnYQkJhG7uTPxEx/QRbu81nDy7dH4l6X5SUKG69HtA/rXh4ESLib6D
BHU4c2WCt+low9Qfy7ngLbUK3XXUZyupT72Jfcfph1Kaqmls2n4vLAHzAIYAjwVZ
lOZkwKJSrHXgfxIXxpKojyPtxY8I5EHTTapfhx95W8/ir/hUPCDXHZ9JFlsu/fIW
o56T87B2bXLrUJUrus/jN7Xz7txCAryH9Q//qS3OrEgaO0cN3uk9SWCZ+S5N4Ig8
gQf67AhL2qqLiT+arna94wxW39jsbSZjG3PUY3EaPSJ3GY90IPapW370dQTGSQeC
spsF4ubftTQPVybnEMjxZm39ExE9RfKKCrsCEjEAB8qpBAErnRXOjEzZlVuYvwHg
js3DkJgeviQp3CJXlhnHjIrm/ANhU9HmNxNd1Erbr/HY/X6TSILnHgKAUn40Rt8E
yGR/Mc3DpgWOIlZBke9ALjYPShUJjWXmT7urxXR+UX+Oym8RO9dlivUxvaOEbTEh
yiPrkROEvpQs/RsOebTLqzzZsnZ4lZ91MQ8+i3pw2uKdwiCItnrO04zwsalG4M0x
e1OwhD1V0Zec3pY+XvmHDZiRJ6QvcnhBDN8rz87rFf+xFY6KJVvjWr9VKJVmI1Q8
bj5nKLhPZdLoRwl7LPhs8Zk5QX8VIkWV9e542D7dTPkwO8AXSXv/8cUr7LK55v6R
GVV5rPIhJF6iUg/aTyO7hZJoNFbNA6tpbF2k0j7xHl5ty1OZirsBvk6MTiMXMaG4
3ANLHMxfEpHAuWJTtAZ5rEiygTe1Y6S0J07qlcLugPUpHoYguvGnAmlxKlJSb0RK
0BgBbCbtogi8DoE0YuYwAxEvL4Yo2aduzALM0GsM6U73vGShNdggAHNydFxhqhCN
jLiE1NVrVizyvIpEOTocFWCaKDwXeHVn0UVirxt7MgarG7stzH4u+nA2UPSa4CnG
0SJhcgEEDVXH8591qQjTkvOmPEDCM3zvryi4Koe0M2uU7A817+y5nS0VWDMRTsF/
JgpvPS1C6mlq3W3lQSZZat+8mNKlu5hO7MFb//Sac1moG9TFYNzUaTwPVTW2PnVn
6P8GhZh1twPftP1OO7tp5xqCerBQ1r8ztAaGcS4yVz/E8LdvflAjLQD+cuyai2Nm
UjsGtEPQEChY9GuLaabvrVBbJHyO8V2fo7v3b0hlxMd40acKCI5gLKw+zb2SkchR
oh83wzBfxgt/4p2O5KuoAkgKcuXKb2FgzOuFbOondfy0Fp6pY0qnYpnwJH8Smhf6
B0h+HLfkJb5OXs3FIYWEzGxu0TLjAn9bZATE+djRC0HVGIq4usSqax1WlMIeIQc+
RSG/L5YJ77dJ3VPfOEyNaT+WgTaqhtAlfJreNSTcDs8=
`protect END_PROTECTED
