`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ay/A4ROH8N6rvGTpmtQcWZnYJqPTBc3GHkrlihadQBIiIpqwJQTyedjDNLOa0jtH
3fTYx98Y66l60qWWR0aEdf+nbS1oe4ixOmPbF1PLqNNhZrJvWySVEMcKaaPIjKo9
EPeSnyzYYUO2wczZB9n0WH6uiK9UAXCHTqa7XJ3gtsCODA7/FMr95MVfOOxB+ETC
LXD/bBgKvWCAHrGTjRA36ZMg0wVnVrxnsFbpCXjuHDZBPgBELZKpFLoJct8bdxRA
SapmGIQEIDjHbOcS/2ywIjZSi8zAK9dKeHhF25LJF6esU4LEcLf6dIC6ekfomq/d
6UoPa2MhZHjQjXCsqJ4DG6KSZHt2kSQTXGHvl0z1sdo60z1/8dyjiPZQBNhV5fbA
zJ9joP2MSXqj6gjygPoXApwnI3uqaR1PcVwrQzCcTMvN9j0tyzpt0/0ihIoVpTDD
rDYmXRr4Ct8XXAd637aPmZr7P/pPetGFnV7YLMxlRid8Z27FqHn3qA84Em1Xc4oM
poPalObKmf+dBR97cAEYYW94PnHj9JEdaHgskejG+mzVbDU4XbVhMTNN/RQA2KTF
HVxLfJufuo3XkOCDE/47VHHFm3E3E9a0/zdFo1i+Cwtcj0bKIQt4/wYgG4SKsKUf
PAPjboZsIeV2pN2NxtPEcGip0+ye4NHnHVP+NwlBD/tE8D/BL30ENgx4YT5Qu2C2
608D+IvGv+IVmGbjR60xPRN1HDHDYIe03fckYG+8NWl7XqYa4UKN9LMezv871sTj
TvMILe70bbGSzcQhakFECA==
`protect END_PROTECTED
