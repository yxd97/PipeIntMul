`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWtP2gVN2NY7gtvPbimrJ+oVisNRfvq9QUBFqtYuXxXWGo5o+58dt6c9s0xSJeiP
EvXcm1z+1JOGq8jBK7xXcEtkdmg49kvVwBJY7Zyj+top/xM7eVTNkQRVVoJYugSc
6tGKMq6CUHf+8Qq92YnrDrroFigPUykfBa0luvR1njwSZrB8ucdu8+gW5mfjWZZr
Z3BrU3rhT3sCrMCsy+C5bWOeLtMj+F6/MPxzI1h4Wetxahb32ju41p8lxRriqG5t
CQaK4GYv+jrzQ1Itja3bgJrgSf0sIYS0A4ku4iaXLGg=
`protect END_PROTECTED
