`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQwyX80QZufHtt5TObs1NM6cIcoCic7Nkg006NC9WYkF35pPe+OcU2T2rvpQMTd3
xyTbGEV1zW1u9VaxE+8yda41Nxxb05SFD29juUCHx7i9wsVyjLWBVwtrnmcWQU2h
reR/gcjZXvG349jXGbaIhTEpDS+WMYLxg6tVbqy06AD8/RITK8gY24MiCOUmjhTs
KvR1U4m34XCzQpFnuCv9jUTh9K8lIvn1dWNEdy3bh1o6emTOXiMTzQEs2hHtPoKk
CjwzqWTUCYi1i6IBSUj+dXDIVkXRIY6uvsQYAbzMr6/0GszoW9TGTZpoYrJZ0/VG
9xFihO0G1UaiWDdk/he3w1Gfj8TSAsDle3GXO2TAaH8XS7kDk2/hRG1w8Jgw7zX3
ozJx+2eI9OIJuqLIbC1YyEpMr3IYsbzPXU+wTahj+pJVNUCudn6S/5344nUZjR2T
VzMwhXjPV6p6KWSQMm2dHfyFRJijlS8XcVqTNaKzRtEUvmoeGqUfE5GsSGC86lA5
qOkQD8CHATYR10gQqh+0w83TfD9FCnM8hV+2w9SaN2ZfLX0HesH1cvBs61L028Xo
LXwdKubEgEGVBAwQuGoTdkeyqe16ma/3N+d7fvAPLLu9Qa6ChCaf0F0xfZfvZ3Rc
mqedAHhnWnCpaKjR/nZVAKHFuP5fk5uJPCC/fx7BtMkZUgtpLLFWwlOCcoqyOtCE
AKrhEU2IyCQTzxO90PGA5sH1T2y4vAjBpsG5eRBnzwgMa0Qu6ZqmTlXgiNfMKH9G
S50oG1/0WTlU0PdOObq+2gWfX4pKZFs2yCaRl84i2vVLduu1NC0+or5iwOGW5Pqp
F3Xtu5u65y7oaHGddznf6pQEBBeSNoAtcuORIZuFMmq2JV8lDVEu5MIT6di+6FL3
sFTwlPU6P5cNijUiTRB0pHu2DcPG5EFvREcpZoaNbQzZqbq08bwxUen0oLND7Nxz
lYZIer2UtsMfXtjcwuUnNJmh20J6PPo8yeJczduNgDf5BLC5qV6yZB3c2/XImKcp
IvE4ldM6G4Qj+0hxOSmSUWlY5wNE9/CRGsnbS+CLaC25J78RFUUzyCbdznAuBLj+
UaJNqOo63aHL3/yPnpEKb4J15wUQCPlGyuHzkj99nQ3rYBumJmLC/Zp9DLGdS5hg
EYQ7q/nJQwH1VNc9+lXjLKZMi6471zRRozAc2hM7e6WqCbzSS2S3+K7SSwJbqvZD
S0phzQYDNtqQpVQ4lND49Xtsjg1GC4LjqcpKEmXktTbdqmVevh15cVUpf7nDIbYn
kw4FhHQxfHfRWayJ6QdP9FsEo0SFFKHA0vPaOixAx/s=
`protect END_PROTECTED
