`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EtVXVgWfLw5h3EDXqlpX6tt8DKcbm58nRqHwzvNSUBVOPUGZNThWYEGWNtjwZMN
GwoAQx666uwMsWtxGtWLOjpnlFd9wm/CH5cclFElNaLhCwvYAEcDGMJrDrqdwWaw
RjI1+AtkJnj+GOj9ydP/hSFwTeALGkb1KN2XoEoOa9ILkS7JnwOlnPXLkhs126BR
0y+pfHGMKuhn1/q9ttei4X+qyQ1zAezGTR3dzTGxVOspk4F8Ww5IwX2hAPqCNTP5
Lu4H2t54zkI3iEBpQKVFg4y7auaMkqfU8BdSdMlR/qB7X6QfASl4rK9/i+ubn5be
UaU4obTlc3wHVVOaLsalwskijXfGaMah7c+3BKZIfCGmajoIt/12b1KEZWBSi4/9
TtWhmyiqUYpGifqz+7l+EqbkQdKMnBBw/dtrQPJhZGmv9H+iEl2W4JxPKEKac97N
Wmq1fWfa/xcjnFZ19CPc+Odvw/zstFb42FbEWkcX+L0=
`protect END_PROTECTED
