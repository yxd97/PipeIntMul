`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVE31pbOg5bkXCeC9c5izV5Qlaq88Ifh4/HBhWMiRdbgKviPZwVkLOnlRPoLbWKS
PrebEizY8tJpbJY8imLnzCDqQ34fYahKNsHkLhwEPvOj0YHkps9jw0Rg+SctG4JJ
qtdip/M9UALc5GE8Obyz1/E7GaorqfG1PJJBXsulJDRVsNOOHn91Eg27CIJWKiLz
LGWvtJzXL6Zn9BojDWiOTQTEtJk3m6YN9YpRrJLncxN9FBdmtwTnt/a1sDGC2moK
qVgZ7lNH8fbKeTO+frcKfnf5XYtk9jqYN+Sw3f9c4Pyf0QNEQR+PIxKoiyV9lt3E
6gWAhrj/0WHnZBalclvymc7ofv2noR0eGMx9N/nUK23rjOxX8uMFlKmEk3faPCgr
b30NshOpELPSUPBoJyhZWw==
`protect END_PROTECTED
