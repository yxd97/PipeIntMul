`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+q62q4w8/GkMk7hiFc+CXMrnBXBUbqzqCLPY+a6aSj/uNBOM8W45IhJ4JNCJG+6v
TLS3utEnh5kvAF6JqQ9be64EsYOYPK1FJKZfzavVyzSzzivfT4M0aHikaAIwcm3S
XXcqlz/nselrGJQPtzudtTBV2WWNEbuMPl+DMuTTkgMscohlYPdU8X+emhIAVh/R
ETLaSxmklKYSLG2qYSWw8/UKJ/0/5+pjcEnyS0SKoVvEi2sPxXuqAlFytePM99Nv
nOhe9lr00YCj0QMfEj2iocr7kXXw9nWK0oZ1ECMoeAjVo2qaXhtNxHCCR8z6+3Y8
/JyMIZ9rrNpUsI/NmuZRWNPyYOdJrvVXnPghO7PcKjaDCEAm/gAbMWAUaC6bH+un
iV89dCTHzxN5OFeEzm5nRHBQW9KPkYNaS1A3gq3dFHbkrzhbzLGFvHe/h9M1GBc1
TgXXbNkFkofSxdO1NfW0sz+tpu1RC64OVyyB8iDWS3/rmIUeEINZwbrpeWbrFpjI
cyhsnlmA9R3rvYz1lAHMpxTe3Y1f833D1e1sIkI1HmluxO7ToIO2ZdIQ/GShQz3O
9tpz9Vvi6EMxhvKbh9TZPJICF8wIQ+7vaXvXld6u9rOzoi3R6o7zWz54U00wOqXP
Ip7OXYGqnjFT0V7pfjjkN3bhmUtH6F0TlJoj3197GXRIZdSWupDRgA+9LBGkFEkp
uFY99XINQj1t/mu9jxvIA3Pent+8efUAopQAs+cfME55qBpU26ANhDlHD9N4kJ2K
NNI2/ijSx00XvcfcyTv7yT/8q/KK7XpZNPVtQ/HnnWJqIld+sutCvHo6eAShCax6
ICzQdZoCEzQ0XWZNLAcfAVsLR25ep9wrvSxbLfsq8+v9lVn8jPrRcKgXvpAIZpde
AfWhHcedvZVFZgmM4MYX4dE0zVlS2f28uRm0UTPh13KJ5s/bkGbu0hOWkelRkXzV
WHeC4D/FtjMl97OArdz4j0DUkGArB1z0c0sB46DTWU4lLnAvTpF7fkBpdFq8MgFc
`protect END_PROTECTED
