`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rPSmvzl/UXiDR6H995jnY1w7H/42Q9w41hsgxdDcLqLUlPP0+w/pcckxItlPm6/
t3aWbKBUtOcx1aeBZ/ss3TPDD4IF3QzQCuqzklSkoTb0J9Rik27rl44yjBeteTOK
oe20xWI4xIyUE6qhTMmhwplyD20Gr/NZVBFEJ2vuRQQ1ktoxOeR+jihbdsakK6cV
8brBVQPyibMTr9oxmjLzkap7UGrmeupcaeuyG2Iu3rxScosXLLiqOSBXGTnYxwZ2
H5v7Cp7UFfR+v+2UuYevmA==
`protect END_PROTECTED
