`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zuVAKeR8oDzGXgEVhVT+MLi5ISrG56DXaagDxBrn3bPUODx6tSy45QQnoNXwgsXq
osK4HmRUG8evyXx83oXCq8AcKBt1Xwl4eyXsGRy8DemeQUay7PypGMN74ni1pmJa
GsDr8cDlm72RpwK4i9ubLnw0ycFuYuVUDu9u5gl2RtmZuHbn3urN7sHW+kiwtc5a
rOZsl1VwwqbnvzIrzmlDHPfdVyhaFSI6qdRizp9oFfFuMqt3fdd5R3bioRDc5ODp
T/nfDd9Q8tha4eHdA0SR2O+X9GfxuzGyhxM8OJftPNZliPwS6VGT03+cPow0261I
C3xoUu0gu3zDta2znA+36HxQnhjF7A56LlEtqY0cmfpnqMQj0Gcv8LCeoPGXiOFM
51sS8sr0yo6oRgCb2yPFXxmYBcGkJIHSMZUKj+cWXh8GfH4ofjvDg7x9y/OCKPp6
kQaCugpKhRv8B7Eo55CMjpQWfb3Grg0RVAlpO01ztf/8yPFHZuig14AhyGi5FB3Q
MjSuzO3lVJgysiEtN3Bmgg==
`protect END_PROTECTED
