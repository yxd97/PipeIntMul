`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I17mL4NuwZ+lTASt6C5md0AR4/w6HnCEd4z9+iTQ68xywnQmswHSfs886zme+ERB
If8ikn7Higi6bHO70Qi4Kqj5CT3ZR00giDv63DC3U51p7rT2fq8pLU4zRg+zIiww
QwyCMoVgxtL5dIYokkE9oaXWYp3/ge0wK7jtdzyMf+iwm0XGvn+Bhj/VhEsleALX
HH0m25+lu4yoa/NKOn2Q2hjXhNbWdt1m+GoHVeBKzQoaAjtRhHlUBuC7ac086w5T
Qn234LPcm3gEIfsZEG84p7r+XSO57+f2PACjdmrSKbz/oLmHkalJTjUKXJ8nL5Uj
86L9+Lxm21JyTCzC2nRVxzUXqGt1XpXyEpJ7lu94r+dMNhnQS1Ex8XQehafauBEk
f26J8Dg3AmKX3OvYsREc+Q==
`protect END_PROTECTED
