`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAv/Kw2jepBsgSsYkiP+PtFMMV+fa/9jCZ0lBYt+hPd4rtHx5Y5Z5CVabUK8VvYj
Y65sYgROku5CD/MRc+Jl595ecY5uiyQc0hNCOMWJml5SPAGU9La3MfURXVoXkF8D
cbxJ0XiJ3wUB0YD/3wcSH7wV5MXoJYtClwZoXL0qYWUbTZttfiHntmx9Sfhw8tKD
GY6ViHLYOliE051HXc2Evh+WNF4N7h7shyeFOkQOI1ztCO+Gk7Ln68SrXosj7ORO
X5dkBPknX7BckSmEIbkwzC/3TDhb3S37jo5UWxQ+o5xNunv7trXcEfCjab/hKc9L
slOE9QDvM4SSTH0lacedxZxsLciD3vrWkVEgvxJU++b7WlCiTGRUJkmyfxvl/491
4PhW3i/cxY8+5IRPOB1qUL9iwm9tgSRy/vFqjBjuBkHKGGKssbg21zbdW8jzjOny
LdKJCI4BuPySNT8sE08tqA==
`protect END_PROTECTED
