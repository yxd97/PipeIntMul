`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
blb5o02M4NhQo61ZGGxQzVuUd6wqT9M46+xhkj+Bkf05+++DTFyKJTTggwUL14jn
kkgMx4FyHYkxZXo0JzmBzSdgl0gkMomlbllIm0E9HjvBZRQ5TIg2TqVsHLTZbQdV
5ErG17T/auQPXRgZyOxXzet6E6ZS8e0NwBoaxgEV0N0zoLp4zBJv3PmdCiK561zE
sqwhA5YaII3cNK1P0eMXjieri3R2L/J+Pjixcd/nYxAUrstFSV2yw8ZBsFxm3POh
LGMqorMBDJxacmOlcBFZwbroezbmUNJ/vo0mqT+qvUodePsErdJZJhf8onwPvTlL
xSFMfC4ViNxmtfVmcmD7EA==
`protect END_PROTECTED
