`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gFvCeYL8RcXYnmDn49piJifRx4QVm4xm/3kQtL/Oe8qCu9XP7YXB0oxogZOihvGR
m4r303kbHB9L6j3WA9fuyXeUrjn+i9PoJsG8CKDI2rG797flXhaBnV0wKafWnQiy
XBMb9PrrrTo6WShbbFxY0mCf7OANzTF1nxWISmHnysegFLQ5qKRynvrKWi0B9X/6
Rn2yONLReIba6aODbt7Rws3WcKnkCBgiBtP8DIJAo3jRu+MkUOLyqYSkFg9uoHx9
cK3TPUwBKW47IqQjTSrn11lS2PFrqwE+aLrptau42dgfouEb3cfBI9TZJuj/q9BZ
jnrNllTCfBNybDlCw2dtZhjfAfAsxJntO9RoWBBLkdpVicmE64uIaUqE5C3D2jro
/iLa8Axr/0pv1z0UWFMJFXjN+vCKM4iyiEAIZo7E6UbBmVKShhsXdh1eXv0LsXOo
yhZsNA/Lm0cKSnz+gn1/+uOo8EOI1ct5+awmOMa3ZJ+gETr6kB9WkfLysg6+wNdC
xFpO8SocePokVH3EgDQ8A/2dlKwGQFQWrTzMBvxZyq11aLuI2ohjbdlzBXHqdki0
7dMyONWj0rlzzHC8S7Zq6o7ZLpVoUNzVmTwA2eoEfyX9g91248emnM74z1yarviC
UNgN3X2hTca8ruW4v7UA+mrJfqMPDbaMcWdmtfYIpUqMLGJNRnXTqDIKYnZck0ZL
Iwb+073nKJkamGKRn/0RMA==
`protect END_PROTECTED
