`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXhr/EyTR+vdi+J4vGfKU38YNqQy8+apMLvgNh8pFMRyVJwXvjq7ue1dIV/KPHNE
uvYLdW602LvJM4L+IA5c2OMMLaq1gd1l4rS9lrfxha7MKqI/EBmuBuMfltVueirs
GgmPWtD4CWdXSvuh9gdChimh6TmiHWRn/xFbS+laKF2GWNwcEkFE5m9k1w2H7eLQ
NE5Cf2yW/7mcBXtZWUtnxJTucZ9gCgImEnSSvTIZzwCbUv4vGa4MFkOK+s6eT6Fz
SrPnfGBxWZl9xtY4pR8GWbBknclWqHgtoStUhZ96+oJzBtzNQG1I9Nrci8i/erKh
zd4Wvo3nUbygcpkaVyJAR8TseckVExMgT4QL8Z3SC6po1ktUOLoaYnJjOqbJEUF/
vqt2Hw0GB4Ka3qPvIY+b/6QAc4lV+Jw2sse6yV7qwhaTlnF35an30ceKeQh3DQGy
sI2lSkfJ9YTmqF7SsxZvOO4ZLpAlI008/eQxHP5zByXKQusChj0Sr8pao7Gnjcwe
Yqh6NfOkW29ntHGpNU3s/0d88Czbj186Ss++R1GKWjC2L7cyuePFhWuNRGxhDBSB
nrMmfXCej713TqnknIQJuYHSz0FlpaxbG0pSKt5hrAMewbRCNVwuxmU8adZFQaN9
T277TUz+xKi07tOFXM0iL3QZuf1BIzK0gaee1aFIUp0/86miRsWpgpnxRCft/ZVy
6MKS+UhGy1aVumjsACcPjU+ecvSqDGwh0tQqYO3Um/HD1u/feDfjVfcBIniScHYJ
tsG6HY78BbC3bc1tWgbKLYf/y2Ti+TfMyPQvpRAGYfUFQ/1FsWeNfZb95po63Uq0
nbN1GgEyfBkhxO6+7PRNnCQpCuWRYQ2X6smmhg6WJhoMEEiq5mssYeC40HZnBfqI
n8M6Ub/HpkJue1k5iBzroz/AxpjHLOdHYup9C76AKAazw3nm9+1Cq5HIYiPUBKzd
2JpGussFZrU2Ih3XrOEGn0uSridgNKajU5aNHbMvh2o5JkBlHyWRfpVNR3RqIU85
atjF1Q2TA3JOrahR6tdgHr5r22KN05sEbIxJ588wrzAR21RbJf+jZ+kxs5A7gyKj
MZXRlUJJeIrXnoDUnqF70Xpcuo+FEXvZ/jzl+VdO8r7DA44P3xtB/uVHske6qMrj
KrsDvCY7q3B+8PMt5jIlrmXXYjLiZ418ROc2ngE7v9VJDO955rNlVJJbGbgDQaN7
+YvSdprpEMYz8Is3KEvb6b12fWmzC8koRZigq7A/wDEXm5UrJhd32IQtA95P9udx
YAHFKBrIxRzLJVdDN/SrLqZOQG9z7qMkiFf4keODEk4ztRQYyduyPj8uGuNbS/MM
Av3ZYfdv8tvSbJ405NYGFyvM2txNVn7fTNehMWAszvFsEQbHK6hwzbrG8sKeaHCj
kdTfkfFDzVcNLa3JeSR6OAc/Tnva97s6K4LLId8GMCY4bVJBh5QbBS1Pb+gKf9Ry
4vJkqYPXen75ZcqJSxzdHDMCerm5pPv1YIVtx+/nICUNXQZBDGfVNeS5gPFXJTKe
gEG+FbqFUGksJyCM+yNDJFS8csx+QWzHtzQuOvanJ12juzKTFHsC11skj7MNnkXY
8ObwogVNgwLjIpXAX3ucXppTD5DBSCgMkHSDau3qh+X5ffAZgI5kmB3Dv5TvFftW
dN6v2bVMZdP1zWN7OY50HgzqDB/yUP6TO5uuXl6z9/N+bfN1pLhx6Wc39gyGR87m
FnyLahdy+oqt8H7imYDw4nEWV533gRrSKuNSYB0Yq/vnnhBNvQ0c2tpx/kW86c8v
cIOQ0I1Eff5Ah5Lbydqm4abjhOm3WoXHuMzJuF10THm8Ujum27Oe1tQvPBhycOvM
rb8dabsUKT82XFbSUiVDjsmtLEhc5LcyIaXfXvc9QfuB2eH+PoIBrUs3NsftXum1
5X/m+5yJ4LCR+wKRJmw8jsTC0cmRLXruUcPsS4eibKO5/nAHrwFlFkBoeiB/A/iS
zlbe3jhORTP22oJNwBQxYP2HVgUt7b0gV75R0LajnIcZ3eaR/oeXtd/uXDQ5xTIb
PSEqeiJCvyFGPTr1+gutPvb3rvCz0S7KfK6KgiBBFNr6iMUBAOM0xIp6CmM20l0O
CCQoUltoZGztO4RJLoqJFuE5tPGGfPmCP7scjJeMRmVZiwv9Uw+QoDrw6r1cCtKv
7rACumpRAb2ymN/zIx5vkjbztu32s+o+6Xw1Vh7/6n47me0hn1PmowDCKMpzvrsJ
ej88x7EwUNo3+AvIuyvDCZWT5cP48zXwj8x6Ytk+mTVo+1alaZZ7tZc77Z4Xvq5a
+K5l2hJtV7Cw4pj3gembuHaRD/P/2A9Hb90BJ6GooiVxL/qIRFmczwhYmeK2m+ta
QdgUjcSciiV/WY374OLGYC5eBXm2HUD73AKkI/FPwypu4CzKGyYPgPG9FZPd/KuI
tB666qqGtEYa1b1Yo1jF74XdEoY3EHMgiBNBdY84dTIB7ovu4jJZOUFhbT3zJaSR
gG4+wviMaEYLAm97VaaML3WC1kDDW/E21HTAlEM7MqJalyHNVdbVq0Ykk3JloweM
URKzSH9N2+dKO8mDg+wwMZE9ErbPa+a2sPgeJrQN1qrLh3Hi/kAT/aB7aPprKtKg
w1LEcPyFFLMT3jdw+ja7H7IDwThjcBV66cSHAODIovGCgPyRnYNIb8ZVWpPhJ8QN
NL06/zXvjIhaRKI5lo0JWN3YVrWZ2+fiuuib4EckE91barLph5fWrhe2g2xwuT5J
n/fDe3LHMipuWYWZzVMa1Qhy3d/+vamiD/Mh9+TUPBexKaFFuwlUkDglumAlkeNC
8tIAq7ZB/+q6dL1wlDdvHSTJ5ZY+e9XDKefvJi2pO4BW299j0YtQPdbPUQFQoXox
G+NjsP9yVzicEKEqKuq937QFitbhpKwKFBdzpUpM+v7V99riEWCP2seJgFUmgZIi
LD+4uTaQIcjChj51+3P+oi6jnmzD08AAlSMol6f+ac63HCbl50tjOZltcwl3WI/E
pbsjb4e8q7Evaos1AzYwyxiDme4WPlxYQTMHYPDNMzTSJGL5/aAXZRpNATEVMnoi
vy5CsgghTPz6JDycyWHmGKVIuUrwHI+rRER+36IM3U1eFtbQFUz8smia+DgaELGt
XTFWx79l9MvCk9vGC0XVDR5z75NHjujG9L2BVckRnXzGbC3dGJViag3k2WsJGiAC
kYCocicXXQCxz3KCztIeZRiFNxYspDlHH3bR6/8bgUbpTWZFsy1WZ4tpnCSPQ4zu
f07ehkJLCQ+LiodiD4ZX+XDb/g/nnQoxmx8r3rTDPnHXrLwfRhahEfPOMZN7U+aa
OGWpkcnZQM+livnJA/luO+/6MzT8F+HyqDL1xsohe3XkFnUifvushK+Ta2cC9K0r
GUYZpxKsb3E8Op0As8CPR0st1r7ioclUMLWcyA8fREOOEc+ZkWXj9drj3NaVcf20
ICDoLry2oKuZNGZ1B8iO9OEt6AkKW6ucSwccw3MdfMGA5A6PlIN2j6TTL2CucGJu
DeTih7TydbIpmPIbX+mpgwGoYPjzkHEq1cYfpEAJl+KCvBbMAHsZdZstNYhKhjIy
y1c/7yrP+Vr4cOOjs5HvMu99oKCbAWs4rHSzd+nTLhnIwqcl73c+cWmvsICog+aR
0NUhFqj1aFXOnlIsw13ziYFrwBjnl0i1+eUF2vv2HKT1u/GGAxughEltkTnSols4
XkAHgh/xjQOG/SVuUIRltXCOLWr4Wlz7vYICx2K82VT+4viId9YUzKiIfupKkqGA
tPJT/OC5HakPZGE1tLl6k+7xSOXIHuRNDVkBwWy/lkyjG8NKPgknKI3Su33zvvGV
Z8RA42eBGZA3nqPjtboGSmi44wmsSx3RNbKOaO13i/LkphRiG3nsMEdBD4U7ljmd
q+pO+nRwmXApznCl7IrXxVX6vg/kQVK4yEPQXCZ47EsJvCTJMmfIUk/b3M2OdflT
THv7iKOP0Z7h0SjbMK53mW96hbaGbb10keVxVQg/VrjtSkAkxJxgniJTlR3yV1m0
nP9ApSOGwOo2FwcI3aXAUaCwYVWHgOmRKnCfhIE6KvA0j1MthwHTY3fa4kbwBuQd
j9qYTK5grOl3YNJynmXC9KDri1sgnMKoSX2fEbrZqlg8XWzlr6czB60wy3FRGuL0
gXy0DP5ocad23SVIb+Dj7dOxYTsE6udKmOa6uqpDWs00C7Wpr0at/j5pD/Dqk1ae
SwkBHc73enq09tn5HqWx9vJdI8dyzAojQk/lzC7Ry5m2yMQkJ0UY/IymK30kK9yi
HjOrFRAJ9FmRTFlhJA9+vep3PxswGg5CipQ9+n57h0ccssDJuDmP7KvlSjS1e1Jf
Il8HM6e1LxHqm+Zbt4F3SbIVunk+BRHaWPURA81/tmHdOqE/SuzuLZuB/pXanrm1
Jp+Q3aOgMC3q8I6b2hewyjEHd/CV0Sco8w0HW52airwtKYgrjYyqV7gzHp1bpS2U
CFYDN+nP1onzQ3gMErHItgwyqNdqa7DwgHEEApWcFIsLspVdsFWOwDnXuPc0j2Sp
SjdZ3mm3OPo4wWrFA8pGIa1Y5I2HrXWvCUCk42prx2jBkH8Ny71c8M3izRLkQhhH
inQqaQYafkyBNkWiYDp7E9Ij/LOZgzHutGfjUsSF6jsclug4jO8JHe7UKCFW9Wxw
Q8h07qfPzU2e6AedBCWZD4HqcpZ4IChvXeXFqCCiN2fSArhpAta7puhufvz0+l4y
/vfu3brQoYTqFa5qEW4oOXcxB2EEb+0s3NWwaaJ34LSWajDk4vZwJrd0JJ9lK4ul
d66a2+IBwjrORlgaq4dGlJKVvLHsBOl/oYP558z72lTyUOOu4NFwxODN+RzB0DjS
AWnl3br/5A/tOVBJwna+jUxMyBCH45K9MaddhRS28QImxch7lyyhElfyiIT5jBBm
3J0RCtm0c5Xk8tdCj1d0oR9O+9hpsHT1urecblqrtGtd3OHC039TuJtu2Dh+8kTp
x0OWdJUhWT4aPFhnXhERb7JUxRojR8SJewUL89e0y3347AcmDbZT45V6H/ESnXYN
++RBYRTGsta22wfCSu+vyB9mvabEVXsH08+AGSo3LTtu45l4Eg+MhED15s1DKt8e
uRwiFQICQJGF4MRsZ9SYeWjKkURChCKgSaJ6VSf/8y5FJoB2nvqcuBjsqOw8Hi70
3VInjy2cD7dSh10g5WylnnjMTE4O+OCbUyuD28WOsKppDSZD/bWzObff+435fYDl
hbEZ67MxVYHZFlu+tBgrD3+DfA/pHGyglwMCoUDkjO8AhBkwZV63jhobF24K302A
+IMlPzoltajMvTFJi9uKk1lFBOiGNSCDFnoOQMg4zp07wwVkzQzu2MOwqYUYLdnv
8INDSbwUpZWn2piSo7E2iTg6jeyF9j8DU8+OU+gEcJL9YRBuFD7Q6R6hFtNTPQtH
Xzl0fBXt0OVaXRlT6ogoEhPDe2uFFo8iVYZtZU9lL1dohQO/oLfgds9zGils3194
O4RPMXvZnWLh6q9DOWuaMqm/+ytADRMWa+GN3URsXPyOq13Lklf7NC9yH7JEA0iH
Wmy9d/olgQhOE70B/VJW8yX+Yr/laV9qa1J8fhTlCKhWHNV5RQuZMgcLwvkZxTGA
km0TprVRa6wV7SCdxzsDznRggnACUPk9IxL3tUEcib+EyCVhAq4o7+fKmGPvAw2l
WjhOQYIPvD432hB7R7x2dzpkR58WOQGFxlsCEjDcqUEkdzz3tNTovNKeT2QPhQBJ
d2Dvkz3IjWlsfNZhYWqm12RQE6T823owplHnQb1FAJqxmupUgxpaec+DduUHfYWM
gtOwhqB2xD/Q/ADdjmtcuGmG2E6J3jcbOXDfz+qVuK/EyJHfDZi/6nrLzPXKCnZC
ZXtOYzWgs7znv02Z8x3G7xBS/2btl9r+Yj4y6dNzzBe6nLP8g54O/cOorQK9IUpS
rmEWc1zdssNfestj6si/G2gQdjQCm5ZvBCZHzUkVaqiOFzvOuFE+uZGpbQaS2/NB
0R80ig9p8u6/cHFPh4ANkA0+qgxXcfDk+kAyH0liwEd+HOFVAZEIqqcIJTaZd8Xe
OZfbj86JclR/aymqSomPWtCSHq9D2zf2pvjZtD5dHoDfhjgaziW9M114PYQH/tYh
NtVJhpCX2uFJ5qk5ey8e5J4gTM6ryAvrBo8BGgGOWllV35ha/1FElQzFCice7nHT
or/t2FPC33OIM+hh2Tan4Sped/K3BEvHc0FbQVA1z4D1GVOeblo/I+zUG8dDkWaR
JWRW2mIvDCsyunYI/WVL7lXFvPOL6T0EHB5wTBHrIkhrS9Q3kFoOcKuIzjoRLUuz
VXjewFnrHlW6hAy/RCfjoORL6NLPvMTapxvv7L2U84uDyWlIwm3zel4OFjm97nls
x1Dpgo1/5DuuhOc0oKhwh/JJsPVPg2mjbcn8zfTKxJf2oLnc8H3MxHYE7y5j+OTI
MWerO8DP2saiu7fkw2EPPF/RCBLLk0IKHKQyP0KaEoEHWeLUoWhbjyorokT7xmd3
/vfnkYxYBOMFyz9c+nUe2vWLtSt/k1JyVSsPzwQfWGBtU5dTPrOz9Oqc9hnYF1yC
7OXUsdWBtBx46yYf5aAV9kVQfYKuKTFoilJv5Eb117wD5d0KyrWwHcVjfB4zutWY
5qtL0b0SSGNlwckhsvNjud4svrClA+HLw2n8+Upx3igj+Lm+v+xYRavmkDUikG0/
QrHKQ3m7GYDmAcNkxDPALcIJDcOTFcybME62C7M6mf7xYm1PhWp+gX2XcGFCsV71
/fGoDOlqrCfSr6rBQawsWqQxcSbJQPKdXG+4rxjtzZ3BxnwvNhNi7lUpyBz5M+be
PMtITPw4ECTtlBqI0UybQAAIBvsa7ic+rxad+kMs1ZCW6jLE7p8UUl0qEyvrQXN7
0dZSIIroavDroD0EIL6llLFDrjT9Zgbr3J1k9fSuav5zU2fQPvQOhIcLXXGoS10S
6M9eCU30mrGAau7XVuTnxOK0FWZOZOTeoLNnrZz6R7t5f/9A0hUJ5cA9gVgkOJUE
Mfopem+BYcNcGtG/p1b2AD18FpcsOCiZ20caMMUbDGTf3y51pjvV0O8kzDJhl6yf
9eAFkN5S5xEPlIJUR81ziuUqc5aDg8C5u8Aq68a/RBOIrY2Dql61yGbrztt5dWT4
mvPd3iWy58J1uFyRJdlrEtc4iNlh4ypf1ZXZxc+yoczgX0bBemC6QwSXT1l9fVms
a2qLHP2PcnAyP7rS/MNb8iodmMq1JQfJfOLIT9Xqcay9NzEKGiN/COLPi3rnnaVb
V8KJiMb3PpgLhpOqCCEIBWdp9v3AmrfbaGEIooWJR0JOlIk8N/EXFSXCZ4OsMvkh
lPoCcSlVdkMd4ql8dK/tG3DrfGVibPd/H+/mWBPjBFTDJGFliwqjf096RdMG67vk
bpa+Nhl7yw33tYHunHpDuVjY50x+PPYSKUs68C26cztt9lFV3qkeenqKA6I4p98z
ppTSMz7i7tgwXPZFgtn+X5ENCV+eEcw94Ula8S1B0NXz/+maHOsVQg9yv+d1vNPl
fLzJze3MsG2fyyJfXTerPCQKVtyI2/IUuPX3CjjzBTL3BbWthOCsH9ShB1Fs1Ffe
LUeAmwihSPyNkc/BbJkhV/SjaxRtxVeRvL12RTf6WWIT8Vb/WRBJWrjNcr+hMeO1
6JptqVKTFBG0EJl8MzTnXFb0xm0CGCgvGBjwHx4m9jXz7v2WycoFB33UAepAo2Ic
aLURP35HXkSkxgA6+ER6p+9M9HQmBq1UrGhpvef3+tqlGiYULu9R8q4V3Cbu9GsP
lSCr0xjVsHxH9Z3FwXOFInVo3osqxEaUg7/k1jmy5NujexOVJ39caNj394l88Sq+
VfLBqJaKHE/M2VDG7TZ5/V+Khx5ygGUXRllTCVDv1jZJMO0vi5MyOgGy9MbxrGjM
LuIRrlpuzmBAPLD+Wz6pTcBX+BC2AL5FMbgOX/sT5kGoE39q8lpnt/3qgRL3d6+i
r7Q+ht7E4sVJy7KRjVptEFlIIGBUl/WYcnX+mwK3Y7TVbk2a/sNwaPKUqd/+oamU
4Q8IaKAXhDFpphWRy+o3pKi617NsGATiXoyIvZHWSzv90tY50UXEdQzTjR37G3T9
Su+JDcZEblNloxx1jHW5wNwrPaQX8rYG3yeyVbgxOTNfw6wgx4ldAW7J5/cCxpFY
JN9nsklC0Ddl34rx52mehL0ft7sNbjR65vtzkSimQ4zaIeo1nJWiVjjAFj5bjBx9
/wCQfU9DmhP3DMLz/O9ue9eGrfmsoA9Kgpq00trCyHue3yN3xRu/vzVvcHgZlrFJ
D/LsRfK2e5+BGA87zEnPcuuCNCkGZgD5xMKfUoM1x1K7gNtGnxnD241bOn7K5po+
seN1ZLrX5uh9KzzR8Jd7ogQNygrMFWwdjXT6QvA9k4qHBVBJVWF/YuAxQV0isfPN
dqc3efO2LppJMUG5PUvA/iSnPhh3+0ofQgUpWAq88FWDHOAxIq8yKl7+NvEwyn9Y
qIXWMaOuKeTAKO+OXUnVTgRnnm+ZR7JoeRNSDA3ImRsjibBeU0Vt4Jd/avEOF+VG
h9Ek5FJmx5REdYZQ0Z9qFlYjfUZVzIxZiF6HRX7vphcMuXG4lDH0jd1HCm3rKO/z
Hkix1pR/m8ImkMH6sXLAHaqp7D890yShciinBgqN/W4R+0yF/dCqqsp+K15FyliO
cgvRpgH/yG7owhnY9kaEkzZcHsiUMlkZ6BCZM8BegioXPs5JeL3xMLfsTtSUbRj5
V7xOg/xAuaGuliqyo3ko1w6n9Uk5tW90UWj3fuO50IjjFH5Ppxv2tsaf+B6brPFU
WDpkTRbl8Y/JH9EEUYtptzuFLzGFtuWjncC4S3hULSkUM53Hpcpg2zus62Q5133a
Ncv/ngsRILnLR8ae5huLhv+sKCfMnStoCQuImifvsGH2Q9+F/YUhU6LxQDqjxKC6
/SVF8L+uPv+JJHM7qFXih/m1Dsu2Bo/CfHLjwah746g/DU/osl2IzwP4+iOHnlrc
a+7wnTmNmW1NHauIhc7TA6PxPw0o5Yx0M0Q2lK2p0JZASS/RSML+UXXeCKgEEFio
ndbgVtzv4IItkv2db11xgPMOF2/3D4ZHaqr9q6PTnNk7z0QI+AXdzCqEJBtMbQsa
pln1/jr0HsbJUBQwvSHnTtHuZDGCr8knyM+OUzx9vs/CsQBClG0VQVf8NG56k49Y
hBfgGmot6+20gM4OloYuHZGUi2KwOFRn43xXYj9sbdFXRX9sGmF5NQzsy22G6pPu
zD8kJ5aDQKvUjFXITLxIDhnXtCtKcg0t6XuT3obN30U262HBVCrjdSUqIOtXh7Yt
dzTlDwVp9uAl4xgwZatcDQBihKKX+EUcPWmp3DswnsmJchYK7SUzakN5e9SlrriB
H0BvuhZfKc/gEZNQLHIyGjqUEpSu1jHKAq7MqCQ50rZzibGuIdRQAL7ku04owH7d
SlKbyI/VmS9uBnKy0eys/dg2i/HunfmBF8w3Y4KSJghkllAH12tC+TMkKbr3qzpZ
cskFHd8JJue8OApgU9BpcUPRJb0Jq4aZWitKinTIORbI/7SGdnS8GK0LMG+yD7Hd
OBCRAzHCuUvM3NkanjBWv909zuUWd47c86a4ydmBKwa9SkUWEuQuFj61HGBYH6uz
JVjUoPHT2seOIOnVU1f4Z3MPSNiOfyARAdaxUMxbYkUKc3J/mwYET06rLlJBV613
FzDZgYaCuJ6QEiIxxiOe/5sIT0AywAxfjS6KoYq845RMXf9kvg9diJ47Fx26+z5P
9nYJ6RPytncB+C4RES6A1i3qDkCtGbqw1EZSEpM79EU6LxMtwR3m4GUsWBJzkyxG
rKJOazB/RG2mBc6zpVm33aabD/LWDwYYuWfzVE68VxJ0HxuLovlo5lGbtwrmLT9o
jxPcttAxJQIZk9MN/NfjUgnJYi8BHMoN7iW1WJtwRDJc3fldvsOJl7H41l/ZczNW
PYLg/cnvxctPXXB/gVUgaQ==
`protect END_PROTECTED
