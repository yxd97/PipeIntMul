`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cPv10u67RTD9B2iWlT9BouUFcOaPNDHIozSiwE1iMSiTFx+Mpwj/OJ1WmPW8/BlR
W2iGBumQBd/WGqew45q+IDcPq30Vpy4w717TUM6trIDxbT8JH0RsGv6oS/gsEyMH
W/nbHgXhRyD0xpxSTp/X1Z0isy+VxiC7zkIeOxx/d/Ifm1yMTGs6NVZpqRkPkwAd
8YY3VAWVlDqKStknPIU+wd11G6cocVz8Y1CFK36LxUJYRp2UP2YmQPXk3BDD+g2V
gWTk3ss1S0KyeknovBzDm2R7B8y6YFXtOhVNR0D1r1mQhlunu4D2+JIGY+pyXvyH
WkpQFj63fEphGjJwW+eD7EisnUFQucUrzhVbpUWH4o43Gcyi4MCKXVHC3B8TGke7
7OJh5bjYzg9bGvSg+XpE09d7aWrq+68UkdOJtIv8tMz+XFdDCxtRgNKgJyKIxcsB
HcQ1bYOjYyPebnTXhVlRsX67gyILs2IyexGkA/q4kp1xHIDIXOXa2GGbltLdUJMt
hfvXtqeqmMw0K5d2gQkfJZonihDr9vwElOCcu8xjGe56HPVEiNf+LRZkcG0QkIqz
kC4lWVq3MM0osH7yCP9FJpLUD3aAGlo6MI6FWj0PPGBUHWg3g4VC1PqMJl37HLot
8YZHgTVvgv8HYl+nkvghr4f42Qx6DdMv2t6IeoWGmLz9+d7ikjrG3IE8J8LpyV5q
tnj/bVo0RNyGMEc9eu6dDuDQqMpfcBNnqzY/ZMkiC4c=
`protect END_PROTECTED
