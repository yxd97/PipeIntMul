`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWRCTSbb2ZuLTU9jslX+1uwP2MfDxZcGZnfcucE6SKSlm21wx5lWLReLcwSTTFlK
xRnI7Z5NTXSVMzLFTqGxggKnzNm8InsisJcgOPgGK/VlVeUHwbStmVTTKgs0MlBJ
OZ8xy0cUwlnTNhsr5gQgyNG7UXd36q+5GkyAT08KEcIS+xgxZKa6xMv0/xibzx+o
yY0okp04xUFhJydHeOJSv+LKAbnWLtqVOB/RBU6smdmUa99G73wQCOrK3Pci15Qd
phTOxNpx4q0JIXaycKUTlybLw6m6TwP7fZROpEMpFUDxt00CRLsbT3g/0ejjWIax
g27BRxZjxwrQCmNbYaXuVBasd1dX97yk3woTFzbrnWsy8yZxSFubi67ELWh8LEz6
RKRhrKDzW9Y+mVQ9UnaOIxwCPZdyXlgv1De3t4ghxFDSAhwfOKsrycFw2VXbtcBL
TA0LfrTtJ/TqLhUFdVbWsxdY7jG/aBaIA+TRWY8NzQ9Y0XxFdQoRV05OaygWqKCw
cUS3H03axlaM1XURUkibVbFUzSoQ2nBUkR1HrORPWd3hibKAzQn/PJrc+f2Ypspo
MxDiyfAaSCt00NiqYcGRFsSpTxFbowMFbO/t94lkz1lkIfzNUxb4AkA6loON+AA2
bjo26tLl1c5bWgC2RutYX5NsS1Gq3lCUZy4yq0HbFBbkFOztnQFa7plH+FKb6CNr
RIZEl5udd6ZGHPiZ5EzEC68VCCyPpIMz1sKmpd9anmC0IAHTCx0yq3/JSIXEi+Hi
JvS+dYhdsDjId6EIhkXI52cX69cz3KgzHBySH1dLnNwYFDqQg2XqDcE90Svymq34
kHMDrMaSRMuOks4dz5IXsnU5zkliczQXBlaQQB5rPxJDzzPOzYWoNyQIbiF4/Hqw
ukBsq/DhtO5BGg+EWD5Gv5APyfIJyeDXTw3CX4fvZ3QZ5A9Qp4/EnP80QnGCruP8
Ruf/+Pa64fq1yB+Hcn/Y5FLpGYqWmzj+mrXvbAO8lhpyfH+w0ppAuIVphX8x50t/
PYJFQC3jn3/hMiWfOsEE3dz0Zy0QevMKq5NtDOGuCCXVHgnpG0B3Q/H0l1YXGpeY
+riuK4imfwmDMxDroNK0xhK3tgPtCxJ41LrHsfZ1J8OPe9gdbz++GkLfO5vW3RPt
wryag9G0sCrsAwuIRGFkRe4SbRDAGLGPca/JUy5kkzDncdblZBsoHD1VHBlpo7P1
fhU0I7LeiVrhD27d2vZHRazLNxNPODoqmsJbdpGorOjv0jqHYmPtQnIb1ddwJJRU
e1kYysHI24IPIKlPSdCFrJ3M1wGw3u2fYxlt1XRP0h49eqmDCjjXzgt/mCbzWcXa
rToPSja8ckICGJN1VTR6mW3KSU+jB5my/451o3cMqIx9sl4Z0eSgzTvGOzxcHheM
W6jJs8J8+Trux7ldSdxXCRd0V+gsUAG1uPjEdluWrqoyw6AeDTUW/eN7S6SFNhtw
+QwDsXA2lZJMcD2OhjQ+d2JlKiiiCItB7+fB/aJJ5XSr17JyqkP6xIyHgYpBOF+X
4vjZUXqvExvH0X9kyagxt6byAnod3Nq0Mf9JaxqIUoNaLpga0RvJO1d89IULZrCB
Acev7dq/HGFoBX88GZiH+pBMZ7Wm0IMMjqyB0hjeZFyNAeZI2D6h7pCLBI3Vi+cS
6yCkGQWWi8KrHLv/wal9+ZrkbQTBAQDImKj/U4x4IOTuFvQrf8B/ifBSDdbNrvmY
FXSmAXzuiUBFCvOKwOWvNmBEivMawTh91I2MQuIRj3Xq9Ts1ZIvlVDLd+/snYtAf
RL1bZamXIQOVfy41P0hBqRpJbYhwzMky+ZJaPUNU+RjVshqWsl7AerzUnD5oXqC2
b/4HLCV0p1ZsO79HakYEdo+a9fgsIJbgKXTwehq+g7Y=
`protect END_PROTECTED
