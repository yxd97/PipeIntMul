`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XgMk0nFJaKzpY0C3aEtMJG4w4scdwuDlyrmZKt/bQ8WmYFFGg0/dWkZfFkN0DF7
JNGdukpD66oyYkjC4hdKJSSlsSUrFFnz14h3e6N+RIOI9RORHOScfhNHqlq0hvuD
lXov6l36W1duN4EfzrDLMZBbvOKtDYbaE59Xx4LGsu25NWVYXYTcH39Ys9oBxC8w
8gHRQsQeuL9mQLbeBNOMvlx+tpkj6PIR7nZkQeNt9QMOPyzh7aAqzfP5UwT5TwB/
XFFdg6ecpT13hXvfHx1RMt+DapweGosTWDkJ6jb0+++21+nJK2t1x2bvG6w/nKCN
gM89/ncUzR3DqR4yHjHSEgI+VWkAFn5O3eDr0fLw6ouUb399QUx8qDwUkznzbemW
rUFVvh4cOgymG05H+e6FrmOQ3aOtK8Rlmil6invNb1bIHQGvP3q6BROpAjIJtX6V
c7OhkJNr1PEO+UjXEO0D+PC4t2FajW4ZzZNY2gbFwARgOCQBwGd/pr+7uKrBP1pd
`protect END_PROTECTED
