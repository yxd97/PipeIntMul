`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LamGQNDlIWpYbBKaj6MAhfb3OqEgcH5uxvhXDiNQSyorsQJlxmweelwLD3X7v/Pn
IzpbI+9d9uYWz3yR/4IrpZxTlUzj1IYhyIE1UEuUIbNMQqHrCAojrjmi6rb6I4EX
B9PH92yW+pJeLsQnEBY5sugiZeUoYfKhu7oQ2aw4qw219pxrKRJSWsK9YgbLxgU4
UgOTgkhXuC/6c4d5/Afr4oi34RyHwPh7iP0lFc4/9VjKoyU99UwV876iVDkNfqEI
YLIYlMY4dOZEl9VNrGmMvRpa2nH/mZdfNu5clUBxUe08Y+2wwpuagv7+QhR+gvUt
La9uISYgpeWX2uEOdHys8cSNXLA5eGgbQnIHn4AhqZmz960y7c1b6sJqptgPLF2M
l3YK58Bzu00rvNJMQqxC2aUNdsIriwNdUVQQ2YoxOeM0z2O1i6PHP7nAB2tGnBkP
JjF2PGoBfkHyQjt/AztGJi3gSfI8ZBgg7wYjpLJAK8feN9ON0rePo6pbaLjuizHI
yxOXZBu+CD9Y14wkrPqp3AshqbqqieHkgr5o1tKY66VMCLmusjeIiiEVidAsNIb2
U/BD/MyXj9SFxk+WDidGG1ftN7/HBN4eqWF5fVKEluDl5jzKEJZZMI6gktbmUGlS
VvwvvXk3Ir0H8kWoxc6KmgtI6xX3RiHdoX+Uyj8CoZExAYBausrbBM1RfSVCkIZK
YdDO4z/VPGMQT0TRkh2cXm/aoqE8Ln17YQ0mAYdJeGw=
`protect END_PROTECTED
