`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Un9sCRYAmUTKiUpSdXwADu3/O0xplaZK82p1zdHs4dMF8x70lYFSJ+f8V7lsrglI
mx1oU46GG/07DbS5DEDSsKTge2Xrc65xwcVtYRcioXJjPa/XgOC1+1nbVW1bX28c
Tzslbcy+jQAmiia6PcjhPjJkM3GCG4dr+F7RcRKtf15ITWhAi/KKoEs72N9Clugq
zqc5S/UFFeFhPaECCU4D4lHKpnyjydbwXYyh4M3/H0amuQRuDL4YdtZXHtcQXDF7
fNOUwi0TWLm7FEy2o+MLqIRc40rNBOHkDgo3FhOx3CSQDBzsP2mhvrArQqbO4zJt
jfq+lf2gwHMct6ABhewzIWLX09G4uxJXvc3VsdDKl58+/P17rOIVtO4Li+4i2RYo
I1UIqtMtdx1NWdL1qOJmfKuFqNu0yNlSG6xXNdHFQWE=
`protect END_PROTECTED
