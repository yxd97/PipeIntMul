`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+OdreZJ9QOKPMVgK/JAdqvHrf6g+TTz6hMIaNsVGIglnJZGLmXfKX/DlmLeprySV
RAsrKe3SyDRhb/QMiZzByEezJAzQjSPL+8oOdsGRgTGRLW6iYRp5nl+bQU9NI8Vk
TDONDJFukGIrBxa9ORLTV6g247883ZxqTmLbFh3PWvptyMJEeuZxgwbwh2DR7631
aNERl4vGWahSykIRdm3uZR+KAjNxK/FreeCczITRlNq1/ufb+RK6UDnxIzc5mLtA
LA4QNhiKrmry/rQwLaYbNstBmsKH6564bkcoos6JwBPi6r3zc+M+e9hr0eD5Oql3
5UObyYtV6TSX9UwIgJ2ojZDqwA0V3go1ax19RfY0Pexkf+lmAOfZ3+EpwjetfMu/
vYfl8ep0byuxrJ1JafktM8a9ovSwnnW/XVIjRh3OPRlj3v9O+hSf1dUI5xwnofPi
Oz9hOKA6PRZeo9FL/+oLvlo8vpcjtN44l9Zk2ccLT51jw+cziqY5PxHxMmXSgVo0
9Ea7cogdeWEANoaCtWaRe7NDbKRvGM4KGdGmowgDC32O7ycOL92KGEnw75s3QS12
w8GrYvNL7W+QZh/+NviysFMdDWOUojon8uqSe35A225CUcD5NHICjVK+9C76Y/8z
ey2DDW0XNXIz4P4Rml4uHnqOUS2R8jt2S8T79EnAK1H6PELUHEswCKbw68bpaThf
wXaT1YlOEPKl3v6hDgo3e/ILFjegd2K7yJqkBaemIfmJrPhF3PHj7IDQj392wAeT
3gwwsRPri+XLy5sMzum0Vahb9k3Rf5+3WkbALIh20GXxLclprpsO9TyRL9qrwX6w
aB2HbmRzBamN2ZsrIRSnDPUBEDE89Hq1A+gYLwAcAZVlGdT4n/ZWXxONrc6J1D/r
H8D4XHAvhYD4F+Hm5jb8XDuhKmb7+Vu46RWrGQ0ak+9swsQKEN7UZsJenVQmntJN
yMou4ECvOoJHZhvjcwQu6BTUhHBZoUEqYuyWWcvBsnFYBMx81YByLoLWMR1gsliD
qx1H6C8QRnt8iO/B/S7R3+RDLXTcY5x35CjI18vtOsf9h9sryM0TdfnTH1gV8HVC
4egmwt1Y83ClUUjEKHgsQ0eN1Cm0+nlrGPI6BcBCqffV2SDf+/oIKvUTpDPaIIJG
tKV7ttIYLbFkFevUdgII5nHFSXJ20H19zF+aR7DsljMWq4sO+M5+ALES4No7aNT8
misz6baRkuMAwjOJEF/0ePyYNq+wPSrrdxj2VnGEFhap2Nvq+D90lHvmRdjKJwjH
nhHYEiwn19kxdUr5z2PjjeLOwUETqyNLhGhi9g0x0tbOpxx6bPzVb+6Jz2DQc+hT
md6C3HIp6ZXSuK6BBr7RxNPKOad+ge1PkLOT4nNrjxApcq/FS01meTAawZo3p+Ag
O3g8GKyEFyJa7SfAm1nUoxOQWOSgTIJKLrEzpwl9GrOqTFh43zgfeziS1xFSnpOC
/LMfoIS5YSnAPvEQhqQRU13wXOfZH8AjcwOFfoxsJxyt9FxaKKZoQp0+qTRf/yEx
IW43m8shhaflhDkdMAt0OCnYJJCzHP9d+dwEFNWw0y470TmgyXk3IqM0DK95pfqa
i85hZbxoc38hOERKqbjFcIp18HaYl35e2SeKmwcNRcePtdc/AppsE09OPRphz8dy
McDpYJGFN1FaKOYB3NY+cWTDkwQUkhGG96h03fLiRPLbWRhdULtZLr/7ugg3e0N6
ZNIVL6cNJOumQDo/MsuLP1OscZ01qDBTM4PKSctcwCKIMon80Ya+km9X8gYypF+W
QeUHiADOYsU04Dvph6Qb1CbRN4njh7W/nlCbl/+6kSEdh6DbSVlk3K7QIoIx+C3q
2T4LHwN4+FNEbrRrwKIzgjDmRnKmHLOLz/AOcz2ct9PjaVNEZ0ADXLVqL6HeONw5
VINmo11co7N+2jGtsxW2xO0LMfap7ezOLnE2Ab6U9uKXEdQyw9li+r+A91Cw/uMa
A+ayFAhbN4CWiTyWYnmBfOlFK2ga8fTfUYww7TX7J4Qvx3WL31FleEsl6Q5L7r6F
+avQY/Rpzis5uIv5udS0MACPj6JxH+uMFWHhYPX4C9gvQJRuzPLRL8Shq1oNrmza
7rauMUH/AOLoS8ZEWSwdjKvdEClaC0G+tRQW+9G/XBtN8VKLezTjzn9s5KFTrohk
/AFkgFpc3pgmav42rDRn4GmYoxuNQljPj8IUdaLRDyV4h/vJt/ueOz11gbF97HWc
VrYzB/X5MdAf+oPDyxCm/ixdlvydAPbIldrm5P31GE92CWXXrrV5mqzXwsPND0JA
ZBzF4/AGyXr3GCgCIWJA4yWTrACKCD7PhenymjED96q1t/06Jaz/F8SSeCV54GHc
gg4cTuFwMus9B9/NwyfKLzO6VdbNLwOLWAFGVkqoaR93OK3ptffk4y66doI2FiyK
NCI9WTxeXJVSUwhdGIgfPJvLuxw80WS3ZY6SwJ7TKyZNpjqEg0+qYXc6xJo1l+5z
1Ubt3lAy2Sggasp6YtfTYFzAg8Un1Oc5mxqIMIfVqGgnU43aNF7LaNivbgTtSt9D
8dWMxFRrA7O1xmjHd5qc6+yTJgjEn6S7cE77kpMiAxVTrQjJ2i5e3LwxxX3gepCB
fuK/MwK4IpP2FvsSS9KAfLeytta1EB1Hbq6zraNapqVsetimveNCSnWFf45gyLEp
ZSjFVhj4P1wk8K2Qp9HFKZ3E2WRvxSG0SztycOBVxAEWEycseT7NqIVXeeRZGdl2
hGa9JPq6s3myNL9CxPP1l9vfkkuOZRjoNlWBKXcgktdiwNdyvCmg+bWnDYqiS4Am
gSGt4agKhUhyj4PYYUtIj+CNuMwxa030YM6hCRNW9kD8jlgKdMqRvwzTZJ0rKPyj
mEZ5/pDs7nXXpj6hBX0FsuUy1HHURYJ95H0np9iJyF2ISQI5dLrkZxu0xXXu5hB0
ZuodUmxnwbAzs9oRt99Qyw==
`protect END_PROTECTED
