`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D5pqA0LfsrrV9j7hKkTht+4TNZzf0G5JevJNomA5/5dYphzcbgBqp+Pktchha9k7
YS0XIDGGnxaD2tBpXYg1s8OXkepZNy8nppfNPSel8qd8zPaOFVysrhZJHxZGQmoO
vqsz/e2Pwk6EsOYj4zJurIijyCS26U0/ed+ZWy1Pz8crWHYl997IOANB4LSZgMhb
G39CMppktCf0oygkN/PUCs4YKOGMf706plhTZ0vCh2K8tObaXLNTl/hI2+uLD8Ki
Mo95WyKkwvZX7Ut1w7V+hag3ufYlzCQp18wpqdfhwsvp0Wl2LMKGTt7B9GANjtG4
XmDf1H2a+tD55R42T7RctV7KzIfjfQs3/hXaE2EJzKbQtOOmS7T9CtTAlPC2isRE
HXxXmIBAJFnuyn93INU6qvifRSidoxRaIHxZzmxteVJKoxbPq7XxdTZcKqhD8wa2
1fVXGqA1k3t2MNyM59ATQHYEUzzfQ6Zkv6YL4MIlCZqn9dH3befSpcvz81oSiHTQ
HlLgi9O+dSmLVJS4i+dJYp/y/8Wg4Jy3j5OW9BIwSXTARKv3xOYV9XNATTQcMgDu
JUHrT334ILxjO3A5gBJvu2kCDOZ45E93hQj0OCKbf+e4Zs5NrmILkpoPg9dGT0R9
0XNpS7vzvwX0W67YssKq6CRV5m9Y0F2Sa15tMDuJEHimxgDW/BFkbwpvkbIizGwH
Bg60iOtWuOIZNkRPXvMQvJlq2mTtM+ScAhz+nxArBKBitJAzknoGnK9LNMSyWblW
bEhdk/ObVBmOupJrRAqtqKAHpqT4j782U7gZI1LR+NYcRF/T0mEcZSU2j0N3M31r
MuGZGQpnSBRvgmKAGAnuPLbyINQ7cXnb6Z9FCYucnByviIchEdioxCAl++xaEV/q
iT/hTwEt5l49lZv/iP9SbFAM70Y2GGn4Ed0V8sOkE+EX3f0Lf+h84vId5jf3Ipal
Wk/Y0LsqcK1iNRshkAnvP43iFMAusiylpivtVEFpAWGLP3ddOOqYzLmGPDZxflR2
xbMM5EWpXkjRBing3ziQvq0VcrQUDmd5TO0p4j3nXDhgC4zaC2u4S+/lhJo2IoBZ
NIISMfoTJyUt3RoEO4CbKo94BG6j7imWNpfu1DafG+DlgWqSISkEwcjj9RvkDXJe
DAwhUuhigZ1YztctpiWjyIvdKpyuG/PQ/YDcrSkDPWM2HFuo8gILUnTbv04ycHFd
z5u9UJE5iVDp4RDmgqB4IgagpmTZZjUrdcPs8PimNSuulohsAT1E0Ty8wei96au+
CBI0nXxOB4Vnfdn1fB4gC5IPAYnJd7iNI34+TtOANGK58s+inPtBkJ4+dAilQ+Cs
r8rEG/fhxa9iAGr7e6xEhPa4HTrQm6NSYr6fAqkeSnN3E0St6Llz7PmDMGwiK3xX
hcX2QdsC5ZIDicsy7Fpr0z32DkeU1xsrEicQwE9FETgduo02y99Lgan0KxWe1aLe
abjpZNx1yk0IsmQX9MgT5x9nCbHKy51wJEnv9kdz7tiZ9Us5Jt6Q9IU/Cyp2poYN
HJIbioHWbO//Yx7r49begKKkrkanus6XMmbBGNb0/nf4UflmPsVO7RnJeCOdpK2Z
PwcwoaaTpSJ/oHnEeiS143rh4DQGFjOSQBLKB8EI72JIYbgO6/oFk04b7VztPkyf
SanrYTUHL9JGpivQxgH+LX/4dmYlXWky6muB9pGFGjGlTCTLoB2in5KwO1e/CEHO
bLVJJYmLdfoprmXXjTmncSN2yj//NDupLjPeQPjlCrPIDciwfYaHbgm16HZyVr+P
55CK2LrZKhA92GM4IciLxkDoMmrTcQxPglqKdNuKh2EBJzb/9K90y+B4K2eR3Rm2
38KOqCAT7wu2iyao2YV/l4hppDYYAPUlYhUk5TfC1KbnN47xodif6vX8thimxrNR
rD/YpQck05z1QBmI65oTtmUeWgN/r4jDA78Wnr8wfh571/MqpGxMbv2/wsdCTOWf
J/EGrBl35/Iyd1U2GtVi/B1BZMUu8IRFflco9s8mMNiFi+QT1VInXQ7akzg626v7
D/PLELum91qLtiyJIJRfJe+9uQVKXQO88NvSbIrUr0Lx+b4m2XJrfPk/X/eMjsJf
WnsJE7dvDESl4LjC0R0H1KX1AIvf2LXYYLeTArqwu9lkqqr2RMJKvui3EE/VhPdD
e4ekLIQ+dHDDnI6l2NeENbMqaTZyGtrSgRCxVU56XFhINhplCFdJZ/h/KvT85Q/w
l5Oh/HNNyBfWkhWn3101vhkmfu3tRZMsDsuiH/hjMi4kGPygPHD20vzu0Oxw9tsH
bVs3j5k4DI6ru3s/ANKHcVSpWFpz570S60881jMHkQrO1Gd6mC1tBEy4CSv8Fbux
8KJkFy9RM2zhncwH+zG3EoUOggzyzni0PIIw1qIEYEJwkmze3QQRHrA/8r3n2yGD
29UKp6+k3SJlTT4xLhBK0OZeHUencalWMLlpq/y+Vuxf2hJrqk+0amRxnYN8X8pD
XStpoCwWW93hVRQ3J0Tj5HDN4mk67WEuBIm0GbtKZL+Wm17RyergBjpGfcZqbM2D
U9Ivmj05E+ME+OgZS2sXdgIDVWuoofJtp3Kfh9qk46bKHIImdrnXZbAMioFY606t
58PYV4q51up6IwEfJy2DOvzNm3o+QHRLbPJKBaU/u8XFoPQdFjI8q3Bp3MA2Xlrp
3I+g7FmBZ8GI6MpWCrusm1FT6b4kDWfrngKNDYguEEaP8Rj8PeMEGAm5QxdkomPN
voCy2gQBiwfigBuNI6WYPdcIwCqlBYCBqZ9P90KHLyI=
`protect END_PROTECTED
