`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLW5bjIIe3wKrn+Tt0TvfgwBuDG/VNEccBwzbE3bLfaSDZqB+1IR/3/vKjF7r5n3
TP8bDLOCXxheIyeFOWVF+bPUS0r1lGzWd5H+ZlnDGp/gqqedPZa5w45E4FuBgkac
Wn1dGzvOOrnG8vUCkNUgyhDmWR5h4LU+sM051AJOQUGhiXwZ4/fIVl/Skwyf/oru
Hor3B20AZCcAxjQcUGfIX/7yOnES+FZd58w78v8FgGlTC/Fke4mih02ZN7SII9m8
CamWG5F2nSFQJcgBVp+jy9aSkZaUmuVGFg0JQv9AQeG1WpzqZh5dWfIA804fA/eo
65Op93ZjCuufwLWHw4IhkGfzGSm9mRE2szDtZQt1sJM6XIEfEDp3z7lVCu5w3AJZ
j0dEFaGtgipdY+d7r7aeAzUvHO8mcjGXo8Ku31CqjRxDMw4ljDSGW+g/jAEeot/S
fe9B5NxVnAWoF5Xnp2aaYLSsCPfrvcK98EfzUwsV4ef1B+1GmTO8g5WjyXtXHE5h
Nryi+8lBQoa/dKT74t46CHG7OYrhVU7YKk6ws6+zj276qfFqLY3GsyoIxITrTdd0
WHZBusorzNVt/hbGBuPrW0XtVvSxLZzrVLTF4xWlo86ylMk/bX94yTBNfAQvlRFY
5Dpa1NATO1wLPbytYqNlvS6Loge45+Z2a5XAhG62fuvCgvNkBNlwCBqGniWTLNxq
c2Jf301zxVXc54fxh5hckfZ2f2RbXctjiNn8I2vQ4pz24AiBDhDLbC2bqCjyzbW2
Ol6/FfdRsEyvDQzFGy6AzQ4VFiTbp6FzislMPbgmoPtglBLitz2firl2nnKo4pBc
`protect END_PROTECTED
