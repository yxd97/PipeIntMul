`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5PcaQ/n0RoziYVJe7SBQeIOlVtjaTCykNu34eyMhhp0Z03pbP4jPMhEkHa3e1kEG
OldXG3oZKCEAK2+wINW1pQg/FjSuUA6bO9kTKGJ3xJjNfDDR++B/pFOWcIIXXiQX
kFMvwtgPocNIhO4WqVLUxdTjqu7aUki/TAcX65brh/QLN0wrcjMhYjEMkIWJI7qS
JfYg+O4wzb19f005YAXK1pDMQg/DcqiybT3wpIIy2qJLVF0pADXe9ozS5t6matt7
q5eQ9Dkq4QprP1pDfzdqM4W/73nDSm4QYjrnHjPCx/t5FBsAQtcWbpOo6DGWQIPr
xQd3olsPn/TbaDEwwI/PCR1Bi8MvaKNRs11ySzhZgBlwmOwN+sd3V9P1XNG34ti9
CZo0Oc38ypV5xaPcjpAMnhgDCkNbIHn0boCVIhlEOOiXB4ZENisgJ2FHYmYG7YCO
4CHHEBP+clBTM9bu7jRekIpJ2ia0jAJ9i7NSh6qWP9aUjwY6R3dxCHGcmCjuouwJ
MAdaHpZsRzR2cbEebLkIzx3YhSof1xFWsNKbmja9HIHd+oGebuM7tf2ZZILE3Ams
2KiZQtmB9bf2KNyCOG5Pilc9JBXWxf8kWvdZ1GVAJeM=
`protect END_PROTECTED
