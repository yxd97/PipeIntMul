`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Yo5IOI33FFof0cGTcQdGkE+/cyTuPo7FN9rIvzaK4XUZiBibh4ZX8z9geDw+PTT
f60lVRQ+TzjYkxJU/790SnZMgdrPebp8PZLVvA/hWMLf7lPhPSf3B8ZYdXZG58rl
uthjyzTGVXOA63DcdNwvrw9TJoNSBOef4acjbwzsWVWugk+Zpd2lNYERczR1tFz7
pPzv9Zpi+3l8MFxk90MqGohKzWwk1nRHBFmD3rFj8azh2hwgQwXXbUussuRWsVcF
VPfyuP8ggANIjLPKfn04gkNuMQ/USCiz3CAKLyVorB1FRa6qDo9YzKv1dwlrNJqn
+BoFuV1o0hk514FJKjJYM41VdSy59Js4Gh2MkgF74yzf/2IhSdmTnDwHz+pBEyln
+C4puuWcqw3FBUOyfRU8oEGaY5GFOoQvdEJqIVatSvU=
`protect END_PROTECTED
