`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B2j6HdhxLjFjM+ktKszMbRKAk5f2G/dQ/3p/bSBBwqDpW1BMt0VHi68D7ANaQQdN
su7N1iO8kEQA1nGaD9C424RaJWVceh/E2NvY/vCFzJNJULhwljS3/d7zpiel80Cu
SP6Yybk2DYUr8XCYST6XaAzm/yUsAyyrF0sq4u8vlT+vmxxCtMwV4S6w9v2cpwVx
cF/qNBCJpLhJKL/r9OybYYmWkj8DhE/ts4JbF+twyIOl2liYNpzZKFMpvNj+Qwdi
NRRZS7Q8YdnBBd1va+zjrNpdW0Fj15bTdUDET9bC9vm9vY/w6h2nZZzG1XwDNdxN
WceKKchtQloYeXy38Sb6QeKO69XGkiKOcuhr87EkXsoBaD3/PiR/lrvUBwgRsey8
Xb1Q4qs8VNF53jerZoFgt3rWCw3YoA2s2wUAk0/WbzgIgCCUO0tg3eSCNsc/XrjI
Dhoz6vz/R3FUoRDlgrEk8XmGegvxNPnB4oTtf5fiPR+f4oPNXa3W+qedfQZEFb2Y
wKsyin4Qtb65tFcbGqXB2waTlguqC+r18t+aaL5AvplVzuB2qUUXydHvQpDwR8Yr
ObfHPHzmXBfAwG9a7YKoXQNTzix2jQalWUoGOto5AmssMeyQ+tA9UCiegJ32vXJx
tgfj+ZzCO/zhwQuaVpSCz0EOa19c2JfSrbbMzdwwIL0DxTCOZYykJlwKIJObfKhe
the380Xr72dbbC0j5k4iArpt7zbb3331q6HWH9TDdD+dwo4GEUftD/VGI9ERLua+
8624fCvlzApwcFel8RZ5MJYvwpDp1dskwbYV9bG9mZA=
`protect END_PROTECTED
