`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5a7XqYd1OEEMXt6DW4CwAIWQyDRdMHIEZVlDnCYL2IQIsdg3DO1/MPjl45lxcwgA
NPDN6BVHy/24kPsaDPNI+kxYLhqe3JIT1zbWErmMO/gStw4HGw4ewXLaXSqKOYJ6
nLanjLLC3QchTYZZW2M6AJtx1GdPq6glCCDkSR2tbqlGsaBVQr5h7deOd3FaaEf7
sTwfuMVv1/Dmi81Y5Y6RRyKnUC2rTow2LBgyLKyHXlV0nDXPHEFk9meOUu83blE9
muFXJl98W0yTRT30ZABDaErua4DLKVinu/HqEsz30D5Yw07bxo0+G9Vhakm1ORZU
i5wsD4P/LBPTYr3PRnkmV37Yw3OBRzyiGoqVDm1LatuW1Ufa46MVOiM2rZtN4ZJY
WDUvFb+9nnab+izXiydx3yHX/S3oPHDrAg3jHANRclU=
`protect END_PROTECTED
