`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UKhG7oPhRETpoSAxv67ND2/xdydWlrIWfpIZxoLICipC8K8z3NP4yo1bZjtwh2+e
WbUdx7Q09tDMhMpRZBZLa0lmjE5ygoj0JZNVrAvm0SiUy2JHLUZBss3YGO7CgFsf
TeejV3XexmnDFlDPTun6LU9reDoWVI0kwJn16V2CXBiiL9YArF79YYtbYK2JaoKO
Nd+FHs6OU5FmomIFHD48t7GpCEnxzP89XUfqA/SrR9XAzJqJB6DVm3r/0xidYODT
QT7TJXULmm0dzT1VMA14bOXc0JAvshkdNVLySePL1GJdr1fn9+8y3fbzUs6l65jC
QnBkMeTFlFWqLBd3EjEuCQ==
`protect END_PROTECTED
