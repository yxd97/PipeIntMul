`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1zOwdUe3XmBO1XWaKK6MJ/we3H1QvNCZkA/PQ88K/Ue4bTNWNWXBZwXHTAjEO5a
Y2zBVtbGqBvaI6+35jezl2u+Z1NSPOXkM6Ri7mWff1E9k2B2gS2/JYJVXS9c0EH3
jbspnEojikKGbirq2yb9iI8jXF1Jw7wzCj3vbEE6ZXsSwFkv3bVpe5LKxtCwdLMD
YKwLReYseQD8VgUdGF29UIWzUdBCEpCpZP1IP9FGAHqpuUmXZUCs0Wz7IeJMRRof
E6JMmrfUF14KB3YFMBXzk0OchwqGbxAXdEbzgLWCaSgjk5dJQ5tQtAmWB0cKJZlL
iAphBTj1tMlQzRa+qj81szvPVM+xTSgJZfgQg8ueQcIwrXlVynZouC2nEtMTyyT/
d1IYQGSGNxLKzD2S5il0CA==
`protect END_PROTECTED
