`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCVjZZagW7hH3yhvIvVOyT+TsFFWvfrNS/kVWknVu/GM+luFftRVxj05KioYQQ1C
+G1R0zpX3Vvkd0+vkIQDwbu3Qlm//C5DpoCRjz91w7xnlhc9qaj9Xdgo2C4HE07D
BInsr0w/FEdQsk8IgAjf/gLTrhCxllnoLrAisPsbIW40kWmDpeh2sPL/lPiO+jMj
fT7lZqTmYgADkgRzYrRKHUKCyQfvgb73NgoV6dSiBR7jPu2oCf8eGddmPvN9usQR
rHmIRigmiwc+PWsRuMMw90L2sCNocvA1+u4XjaKNRwk2w+4VipjWBXQob1kBu69K
SMKAxz+93lpl7sBx1xSIQdFm+xCKcv07KzAAFY7Zm8JxztCxrKyDuBLxKOnCaxjx
dATg2/fjYhbLCNXXQEy9xDjEfiR1/AtxcBBwJLY1olVrsw4Euy/Ekr+lNU4BgEQO
`protect END_PROTECTED
