`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R3Fnv1H9IRuOisz8irHCi2U5GcveeZSzex8xOlEx4McO+pKOgbTa9KNnUU47Fagk
Up3c2Mi2n2xtzRpUqf1w3MuFyPaC7oekPKml4Fos5CwoWSoTk1kPiuJZLdij5vsW
yu7pupyz00yZzSATOVXiOywkjlRMm4Vt3EDKP3Y+focA0/x57wQAU9Y0SOSkVGCw
LXeFXPtPSzOchBHGY1aTS7dZvvkENHzS/tQbi9WNAjdG2STHiTBvHngkvvW9av9F
K07PZol6S5M+9XgqwwlQ+Ez4yhMV8nYe2kpSjOL6X6y6Guj1VN4fGBJFVq1TRrY1
syTKAtt+nvniKICyeZMqsubSoIdcIfZIrWX1yyMsI4ShZyRR0aP3YpmxEMEZTSaq
ghYf9Mz6uXGLNPWx7lhrQVzZEqlAeQMcJrVMhZci8oFSl+OyXjLm9mSJM6toFfbz
2jwVRiHxgzItic+lbYUQmOSyxIi2unGWPuLLn4v2LzaxysgEJY5h2xIlh0S1ufYO
ctOLFASWhKw8n/YnGNSv4WaIXstDC7tfCL7k7PQpJVO0a0eOX6GM4mVeJxksbKsI
RY795YG0JgJNz11HX+uzgbpLQZU8gR++kSmPygEak33OX2fmjmaYOTYsG8He20ao
pkaUYSjqil6wmhx0PJsP5g8b8puGoaG4JEmeT0r1rLkLHduLhPo6hKMAQAkJurdr
LQlYM5km2fLlHpME8Jteezepw9Y6TIMaM9k/DRG93P9oyiB6Jpmq8xmiJ15fFAx1
2OYSD+LNLX/leK61gVQqmsoTP9aEtPI1SO42I+ySo1bCM40eQa8qTd5NCyRJU5Sh
V+6GOI3YOy+1lfTEN/VJq+lBL5NlAy2O1/BMBOAmw5UN7T2CBB4oZ0GBDhX1fnC4
WQJKbtTz+wBZ/m06cWRpTr79FDb2LO5RtBvD/Yl7sL1r5NbotWxXZgXK9o7ayDql
R+5Rn0mQZgqn0AqszFy9SwMINwGka66FSfIwD5uvvMgsUUx4amMA+1QCM35s2dkF
OtnA5gWJ0bd23k1Tex2pMZvqFl7+WlGMfF9Ak1qIILro8OMfGiKpMEnETbiRmVyS
WTmxf1YbQ4Iv4vlbVcDLivSDAotudKrlrqEmK15qUiAg0L8XWHUtjjxTzXuyiIdV
CiYVtwe/0LZsoTVSTqf4RWpqT6TC1DDHEnJU2p5HictFw0XPY745I+t/RPhzmOnh
R+uU98CMKW30+r8ccQQOLIzlM2L+aeMbcODk1uq1YLiurFbPd2coWqmyuxJVMIgQ
wzUWPP9SPT4BspbHpQttE2/yRaZ7wdApMw4VlSuK6Li1mJnZE7BWqp+2asKTvuN+
AvtXZtSZbmWBwxCAVYvOugVR6F2c+iwAwDK/8Bp6Dgk6BFRXGJp578LH9+bkXMH/
+0wQjwtEHCYNcZwxyMNAdBYVxKXAYKaTEUuHYILbhttZZsOVywBxLH+LTa/g1XZK
IWDV+lVQTmpNabCg9BsVkOZm5ttrNBfQ6O2RotfqSFMCFqJjFML8WDn75+vG6mts
lfbzCgzuxwLeUZgwik9le3UKocZ4lO1LOQbqtHwLXFTIGk+xGjnhPHUMfHXbuMAj
ZkmAhNr2qdfvG3wCbVZLwR+os+uWkA1MRT2HEtWzHVHRO5JBXzMRhEfnuZMNXnXf
AmZ9J4cr57cyeRFp5x/JgZ0UGCojc82aIJ8ObdVTxCjZU7urSUudB44HajsSfHkF
UjxOD8aL4SJ/KKqNga16yTf+CqM0iO/i0n2K/8QNN/2gkzH4f2ySz29ZdGDr/RgR
EntXWu2DNQcKusafDY5EvaVvZbESVGel9yzCJYWXi/ayXT8F2F0pJFeDFG5iQCiW
yX22uW6vNfEgebmB1/jX8oTTctWieO8fWTBHEUp4qTbA5N+UaJXkufe08ROmwAv8
lP1QZzlLsoP5BCuJzmJ/quStVRtNvdaLRt0OV6pk/yg=
`protect END_PROTECTED
