`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVnpXeIGar94WIjbta1qIHkereIcECaQLPOQ+iqX2Eq38mJ1TfPMtFFpDkurjwr6
DbUHnrn8Nj89gObwIF7nOB2f6gK+MfTzlOdTBIwAtwFe92jqW2CJrD5saiOCm5TX
OOK5/97PB/F8oS/wGX/XovTetvsJRo7mSGuZi139YN4c6/ytqjDhmM/Co/CPQYQC
wJGjd7wMegBKvDiROb/p1MRmftHtXmM1OaKLPVGLpkHhcZ/F6ljHa3tSe5LePjBM
ZAF86U5ufUMw8FTRShXM8ZakssEU48mBj2yaPz4syuFm11Lq/AVr7fxPXepvjyzm
63PNTgLuGKRTE9bJionZ3X+HVrrWa3hRu0u+SUizDscO3wL9Quh/oKNU5uNow2Fd
vFpnr7etXRVQYHF0IgPZnjHrWZgIZS0aHpm5KetZBhUtxxsXyy29eY/+0PN1K6k3
TYoV0++fDxfoF1wNrdbpa5IkVszm6IuZfeZ1YgXGGSkembKLF7Un2n8nAQSDw0i5
wpUgYTWo3FghzDsG3jwnQXCo49lwPEqhXrUHmvej+uFHC7Xkq4BkOUABrO7x1+gt
ZFxwL8+x+xxWgDhIzI7c6cP3IyNTyaIPJwJ9ox8TRW5HgxdF4QFBjjsn0iUqZz8z
r0x3zRO9bzV7mUOpt/ihTGpQ7LvD3XOcqMChndoRpI7A0eWQk9F0mvfWoWYtbjBM
rsLT8n5DIBQJsePM1CVx5tbetXFbKo4j3TGybt9w6bigHfasndP63JetOu1/eN6s
p/3ZDX87+vArg7zldOPENWp3Q7iz7gLlVtjayRMDB+cjUwU2V4x/TqXAM5YvLSm0
nFe69+6XmB7CCvceG9IPNOMnJEQ86TCPeewGDMbwVXSUt1PuK0t1hac34kbp7f+S
+8GozPmkmNfzhxYd98HDTeQt/cDxfYtQhzzfCYsTNT/3l0bLQ6lnOqDp7Qypzawk
Mp4SE8oc4sbdL3VzXWj7QMV97eiBo5aBXZItrUCxMCy0KMuMiJnn5IJd2/UGKQ6I
xymFTPueIcmdRFJQn9P8LAHAsDsdMnNrCU2hZNlD9FbcLYQsY7mt3oiSZ826z8/N
PXofAgYeY/YeoAAlkh3GmQCP+K3qGZfgIfXoVABGOKxOhGklC4Kj8zrI97FWHoJM
cRb+5Pwl8QKfu3/TEtQfwDOD64N9zCkee1/PRix5FpQ/SRWC76OYnYYFgYIRmfP6
YDvT8HXV/fPNuAU+TAEZf8/ukdu0PbYWwagHFFmj7T2A7omWmqUi7+C5TmUcCok2
dAHirdznJES0ZGbn8Uvw3bmqSYQiF/2aGrGTyNwwaH4xwcvaHHRb7Ux/oH+hsPlh
c52d/iqrrDg65Iaj8yvSb2zbfp23Lr5lYbvEiyjrbvPbOXHLclMkiknau05IjY2l
NGe48+1jsfw2mP0OM6SJfKHr+5Qgt77Ncrgv/ASwzB53OPBVF0h6NZM39nI5J6jz
cMXB8wWDPBZSRvYMZVTh/oVrnTobm3jNxAVnehSfCOP+nqfz8/g23z3aDAO8JO70
KgzxRMwpmToaBplX3gdklR1uDe60ZxRkxDeJoRiPeYsNSsrtnjPevyt5UvKzOC1T
csDdwXwSOGCub3brXGKT6A2h3ogQvsCHBd3GeYmM92V4cP2HlFAgWoiK7mUhF+Sz
c11O7hHPOUmWtjjgi7CGdggHe7S2HIsjtLjpgOesS6uIhKwiB3pO1EZ/Wh2ocn7h
LXIEZs3j0jn1Gsi4GObgcjLln7sgPV1R6nRKDQRpM+JhxX4eii4RS6bUiLNhhaZw
JHD16zqqYlA4AyhN+K9Soe1YP6uJ36i7k3TLo+Y0nYHTKU+EdgyycvoQYxif3V6v
EjhdEGd7Z/7JG0voQE4DaJ/Sh4o7152l6WuucaAxxHxoQAgl/s2kGOKFOOa00Lee
`protect END_PROTECTED
