`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WLjy0XcrqVlRpCQ0nEuwf4UPntHIfJ+zXlTAxZACGgtNakRmrbbE4vfw9CbQLleN
r7i3uZ1c7jnqHWuV4wEeLC/PikifymEyNn7GGK9QGHIAQd9C3S3N2noAdaQSpJLw
fvKCPnn4HeDSAXChUV68AyNoFSPJaTX579+BOke/WT47DmEct9SUHhwegK0dtb3O
96rr9O2sbvezkPYwiB/ARtqxTLiMVquhabMIrnov3/TmavIgmykEaW5yBSQyfath
79+AM4hihjuGq1z6DF9r9W+uRIBG8yOfVm/gjbIyUzAlZc90Oehsi5i/G4PQ5XFA
mNuSWAmFZUxgwYal8Ge420fUkwJOWpDlQ46PUGmSMsvEF7tL2Ov2zG23eM9MTh1X
OFY4u/KD7JVMCEet3xnYZPzU94ZEwRY+2i2RvRwZKkhhjDO+tuoGh+1g6NKA4B8D
DEhnX27lgfl/taYIbRy9cHFwoeFTzhAeMz3csGkFTec427Pg16GNv7QpBSYUK8fy
nYfnNLkuhBlOBQNoMxzbsQk9ujEyXi6FHNFJFwVxClKyiJGxZaUK3CwKjsB0pFnK
LJMiNTacgsauDHgzH16AgWs9MD71npYcL51eR6mKOCF4HPwB0WZYpv41jKmiilZv
2/Yh+E4D50cHBv+3sVnJz2Qw0bq9bFciqIPCruegiVxqmz6umiXkmKBzKYnlCKNm
oMDKDn3fgXDfnojf8Cs+dA==
`protect END_PROTECTED
