`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKohTb/lvBmHQQ0W5CrpPWXBEXvg2t8inbp1ldWlzxSKzjeoSr/RBWYBSIeWfo1h
6mGiKRkRuAV8//5NnfGtxuQAQOVDzIGAAZSEOHils5xDtKCHRYVA+sk7STk2wnod
jPb28TDYb34JCP/ZTUH5t6HCG4xuITiCJYQbPY1dvEdPX8cf55JPd2Tk6z7ia6B9
DqPJI1z9NIPAnh4bOJ8W4+rwijEHY4o9EOi01hPVD1I2KFphNUluKMpFt/DZgL5h
/P1kwI2ecTkmKcqq+1b4PU7SYDs/fqgJfHvS7J9DNEcrM7/1aFhabIx1oEx05dRV
wMjnzLS0JOhwBUI35PyHc8CtJ0TkUV6URqVyWo1UqecF3qyA7AUH9w4OI2BD9tx9
wQl+xp2DU5021zlWgeLcMTsViubrqK30BazqgdmRLpLR6Q6jDy63+Wa3qFs6l2cr
8GxXCzC6XEJWljnj1/q1zy4CXvBm3RwaHtQSvpNTopLsqVCPqq651oqi6sofbwYj
uUyQv1KAexlTWFxrJ/fEnSz6b7PZi64YSFWlGCnEZDe7i+hnq8GYw4+KtLvWR2EC
+Jx2OQ/Xm70+kBWsBy5cLJ2rf8YxIdwuv3DCMh6JXlmwkoYdaSnlMpEgznywsW4B
hrLWKuKCpsS8RGSboLybo8j6PfUJr5VFof/dcUWpytT/ZnjoT/cS77U/MKnZeMN6
ntJr26BaBUdRfJyz6zlalVYtazR7cgRb6gjgAEBgb+vH3w8hVxqiV/oZmyTPOJm1
3A48OU3s79zfF4UiKKDvLZ8/S5d3MvneWctdYOGt47tjaX+WKG++2ST6FDFMHyia
c2dvMd/xvMo1VBU6r+PVdaMXJeXoWv+LjtoXHseba3hhkdx5OPjmbSRCxIl1YYVV
n7ljPQTwwAx0R4sH/i00cVFN1kvQWrI6n48tJhmzBigSNRvZE+H0+CpTG5j45hsZ
FppO9xU90DkAIeWQ1DIxnWfDLrZM2mh0D41kEABrRvIhajcaQ5/JkHPQHhgiVGOv
uPth6rjSEjKd314FxquRcWqpLtxXH3RSLjpfN4+uTpxJIXCHivhQgfN8v935IeQf
Dn2dZ5NJoTPt5moqROUjHYusFSoMtir3GyPAF+1MvFVw+47MyBVsP8AmSlY49gGD
Cj8wbgV8pEeQ7HVSi6Ci7U2sAYJ2Ntn1e0zvBhHwbW4xM1yGvm61dMkg4+I3bxl4
V6dYgfwZS5NGX1OGgnLuX/me+EmKWFYiwrFsj156ZrZ6F/QXNVK9tlESUCjq2/P3
VPGm0lYGt8wuYGAcLGjn6l13GoupqmvgR8UABv/MYFEZJl470+UkiWg3ASbQll9W
ELRxS7Yssj7ftv2ONCJuBrmB4DN82qZRIoF5ofMeSLaDbe0K2IkCUWuEBuPIkDfJ
UmsvlTx6uR0nQI6x2TNOOV1ObHE0wL9rLg+vWHID4XaAdH9X6VDFKLravjE52/SJ
ljXJKxavazhczqjVIwaSiGQqLmFHmj5TD+EHDijTfYcFLgrjHIp2NX4/RcqZ0QtS
aPVkd5jLfwWGej37XKyrjpyM1/NXqPkdIHavsn2JFVE00LnhSqKE5B4OFRztQ3vD
5Haq3K5URdirs2Qsa1SVGUdMLZjpS7/fCbWuupH/U7AEQZZJlPCYo06ps68x8t6L
0lqsjlnVRRgeLm4EgOS8sa6NSXJCvEG8hbaiE2o6PJEvVHkNRmfyLXfxVZkLdRer
XHuh2WC7kKXwDbPgjisTIjs1s+s9ZxDH4XQjVMO7ViEtoyptL/pQf4cOxY8yZnij
7CS3a+slMU8rzhpFgHwtB0C2wP6P0Z4J+OGTVMJtPrE5KJLXiw22gZBhqdWCTjoL
FtEK3m55Jrpq37xnzr+eeuKZnYLrUZyYAzaBHsKf+cnZgvelQyBgHC61xDawb5I3
QBWwWI89x+j6+7CslaDclquT7pY4jVWso6vvTKqaJx0a2l/u7ipXGAo9ismmrjfr
bWXmJ6c+zCmxA8HXiVoS2g==
`protect END_PROTECTED
