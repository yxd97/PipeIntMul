`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eENwig9bi9wqKp3xw1AAOjT39WvIYyJ5bv5TvSmsjcLkSMjtpeaHNs2YrfG93llg
yMmULpx5N5kLBGqB1u7rtTO/+A/NH8HyGzVj5DWD4eOKhoNz1ogDst7R6tUD1Iy5
LbAEjieNIr3sQ+ilGssP6c+FGf+0WUkDwL/XMQa0q3D5sHxIB2FMLNVKDKDFr+Ug
Hc6QK3k8PhdHNTU2YyVUgnNZNcRMcRbdhSQ9q929Sh8F5pCXVcvknZrPjJsZx3T3
Tv3AasfEijyb3DBfvE2ZCi41GCTLwM1UXZib8tOGlA56HRRiiesJFW+EM5vZrol0
LAaVWyDLTSKUnnYdU1RkdSHZhndgVVDa0qr5qXo8poUGjBxj0DXqEU+5Srwgjgcr
QZE94kzEoPV2WpdmUg/UGfYz369nxw8+Xcvc8mQ3pECrV89/DmgAy7jVKh4fhjIj
01enAHDxCymuqR+BSi3pWNsdpJeTzhX8Rgs9rxb2LbyO0BSE2IZ0FYCQ161TfhYw
YUIlH+wXBMAnnf2EAVSmP0itdQsKa8BZwllFV4X754Hycp3qp4Fqh4T7qKSHlWqN
hFvh2+F0QRZXarfu0c9vHTGG8xwlUYQMTOzRiFUzbEr31epKoCoYLuAnlP93VVQ9
A4QW7go65kLOm0jOgPOC50yfkfcnOO4dDnThDpKTaxBER8mMlWuQlP9eZKfS21YE
SfEjvUPzWBrUcj+c4bVH6NzciqYUjb84A+eB+V+W+jXuz/xFfpZCI8CNdhgC8YFp
5DvR8besd5ESji8nLtbIUUjVoVeItaUyzhM7xlksCHjG0iAHmijJ5QNqYIiPxFaz
2K9qDHHI1v7ibSZbC1tuhbW7hteifvcE2m6vnLks2JSxKaBVMxgsenGdkhcXBEbD
kDKjEl0Z02I2INfalz46r+bXGYQ7a5MbCnVhX6MIGwFefX6pEzeY0/PTXSLbfMUf
FSgzleJjpSFP33/CHOJcE0y+J0SRpi0N6zWmbtIndYhGjlITYRz/yjBOLqG7f5N5
OPqVyfGpsp8IayCg76wHDWichGmqLNCTWup7AlTcszE+sll8mgfZKkSCZxHASlWa
sHmVEHGRlMpf3jHLlkIFvWil3uTGX8J/HcxL8dmotk6kDO4oCdFb+HdVPHchO4Rr
sJHucBfcR/CUb/lNXInrPWAO3vo6e18J5EixTXorXyJ/2Etb7bbuguS31O3ybiif
NUGy0B/AOfULidKYjO5GUowGgaiqb3lPYpQvJhRM6Sl9dL8zYdvkM8+CSiNoeWqA
CiEOk/4WnlPegHox9w2qL5TLyYO7/cJ8Rc3P6AZgzKJy23JtB3x3oUCyCn9V5Apq
sYzVDLCzrm+XEMmOoZO8XaJIscegwdPqRKBm14DFBMUmxWDMT0JBGRoU7YmpocAF
ztXpq+9V5TOqZXHrkTpHb0mxXkbsKs1uczVGJ8t9K33ulUnKSF7WU8d+adtFlkTU
pxM7rS49cY3vCVTSbG1GAmAFa1RT/jdy3d4e22BaFUDNzKaekCYHiwDb7mbumrax
7VyYw9L9Akdny4uLZi+hhW3ijjKeoKKH7wHd3Fh21xXDFCFiEEUgalvpAMC7gTNu
ajBPy6Mx/WsH+uKOoA2kuH1mfjWCj28KuBxXwxSj9dgeuLRwcTgnPvtcf1hPd3me
kQu7F99XWP9R//9XyFV1X6zym+mqNu8zoZvZxhQE4OEwXmqQmc6Rh2T4EjN6GMAh
1S9GBwSjA7UdHNt1fH/NrYleq5ZkeZRb8bTTEH7SiHKSOHZ+ssznDJWstuoDIDQI
cG6Dg4/2GOwb2P2caAT4d3HcMV4UNaY4A91pbHzWAHt7rC2y0kvp4+LSon8fcuJ2
E28tJHNHNlDg8yhdY6vZeh+xq47LspE91+edKijXDzd+jMWBegbtbXv3aGikXQuc
y6QfE7gm1jUu0h9WUBDApOdh2+WDYEz0gf5FWkEXAZ5hepUh3kr0cVzObRuR32a9
QUHAg52Hna9+RBH7VcHKdDA6+u+wfdJnCQtWFH+ogwBVdovsAUHMenTVujW0WpEb
5Rn4vmRO59OXZ2kunIj2AOyYqpXv1vCNhWeWBr2cKWxTOv1amcoxsb9hxc01TDGC
bXUKA8Kg8r5OSpxezO3lETlBzRx9JipEuu01jpNUoZnzKwAKkj1JjBqOf1CwAK5u
PG5d6/eXCU4U7GVGuRAspJK6AWNVTdjYZWuV0FzVXrLuVeg6QADydJWVb+iwGPZ7
X/nP+7qoysA4Xj6Y4KQVtXM+DqB2EXyZ9e+Hdhy4DJcQkiRN9l56mEPKBFyssTCc
UapB83APjy/WHLjgG1R4l36ut+lkXjJQqoWVlT/OzAySv+AcjLpjAHueHsSN5A/X
nVBVYOBymWJ/UkMlel3TIckp0G0lH7678mmhgoozxKU5mednrnGcLlHfLrWsw86q
vYQcUe3dwUuoTV09jS6V+7RrsvAHSd+8d3gzNdU/2o6gAkrRU5qSL6ZHx5zARAau
3mFUEqg1FKcaUXyF7KSrLWJdqiEBhum/WtVozNphAvVp/iPI5Y1xAUi+xk7wZnTq
CJFaHRIjeSalXRpH0Cnoz/Zsl4czO8khc0m02XzSYp5vm/75qVhEaJN+X5A0Y5Fz
+uPMR+K89fS6J1mvHhw5xKmouftilK3fCUCQj12E6oeTdyjqW4adRHO/lavsuWRD
mS1+mYG13FeETSlyTZ0qZoJ41Wp9OvH1Jr9KNH89nh3u7tVVKlJOAr9HfWI151u+
gV0GVaorPNJBUizfKwNVSArin0I6G3mvutMUISS7FWzi8oLLzIurnEwFulYfPupc
OwH53eC0eWeiPsFrd9YGtVKXIWDRWl4pL4aWSiP/PxwizjL6tt9RIGdIsYpyw8O/
4TaFmSaKYY/dhxfK9HYKmDjoeWQVtQnmJRHRKWVAv7cfWNzf1Z+MGZu1L2mo6sv5
tcjkuAcadginWe71e5OPmkLhMRWhc9UjcxbPnzfeHlGDWC4XgqIhb7s5IdL0Vg9z
LrFhuLoBDD0whGF/DT47toNPe8UFe3MMMKWmjNnJPjvDdx8+kHP0WoVRWmmvrd6V
T8hqioKHgbkC3QgUxrOA6+PN1x72xuJGAZmSkW+ODYn0NILSFB9eqYVjrAmZ0Ehv
TLt0MT0099LnuS3amiKjCi5MJL4nPUTbyw18XgMdqbHWbQm+pnJ5CG+jGm2sFPSf
/sqHXiof7di2BbMgfg8+UiXehV2OMI16TUfZLQ6qUna55rHhL3Fij5EPhfrBdVHz
mt3EUnRyyX73OqEc9UBixnXYE7vxQa6sipcJSxUwVAy0bMR0rtj6vSfhcUKIVYDh
fDYSPKP5ApMeReqhfNcmzw3DvlRsg1+Ew3X1XCJTEM6JnVL5os1Hn373e3br+CeX
EhkLe63wwproZG5dl07ERgZD0R4oQwPMbMMbaRdxvU+wzlzqPsmN/7lVh+Rzppo/
e+cVsNlbGF/2zJglFGzBM5gvNW5eDmNRyJ84aChOCJw2qQ1I5RsM7f3up/cXcyL2
h/WMVWSmqTUg2eQE8Yz5aDju6g0bkVBLZNv1f0CPRfFtmuP4EGcJb1rHTSnO0p12
0fJOM4r3j7/utGcBYIkE5GuanhbsbUXX8kd/mHmd5QVPHJy9tzj5UZAgTrd9llU+
P+/2RMu7RVdFp8uIl+nDx4614j19luWOQcS7r1Q/wrpQ0CsX9qRZDJHGzI5yZvWJ
CQp5HMi884wVPfuE5VT65mGgMRdQ4P+S3JdP0B53ZmRReKIjO2kTHTlMrFs/NIPx
jewcC3mZrXWIWIJLbOaONALEJQVREAj6/NE+u8k1THrZ+Kx1xH1rNIKviogirVD2
sXwDf0shQLNmooLBvoRIY/mj9FGJ3TKeMAZcFj8v7UmXScDzpZ6TD2yM+0XqNsPJ
PxKhvk0bEv9lwtxv7ZSNoDs/tVASCqEdcGJ7w4lHm9G6LgyHEtj/gDhZpPHZlUnT
ouPgRkmfmKrQFEFVacGTfm9kZuKbO5Pp4s1afSnd4vyjzxdkLtpykPeDS1Epg++8
wOxP9/o7Mtc5THbGBZm1wgzrOYFUq3fVI9OHenedEHEqIKw1/ix23TvtMIME+tz/
GR25bimjbE5C6dIlivigCZz0HhCqZYZEf1gjWx23PvWIcHqq9M2kfl1WMOk/cj7s
YGNl79LvB/kK1CqihJQFEyhxivrvSZEEELeShgQ8GXHU5YnLxFma6CpiYSnK+Ww3
yCCUHmptW/U6JfMJBMayGIHVEmMSxRGaQebuW1FZ8ic37HOF6SKkdqyBsxvgK0tc
wdvcOp7zYZegXJCtzMXQZYmMz/wZ93wwPvM0uvzWLwBrbDSmX3GRdo4bsZrF5IJJ
tNrhKyor7VRmK7ehCeN33aV53LJMdq3ScGKGYIJF2Os22l/zxFNqWemIzg9vicYX
BC/Fi7eiYAz7AXbrLSR40xVFOEqCocBesYCK5h5SgWpPtVYaPumqTigyW5GQ8q2J
Fsz9/ARfjQFL8oxIGNFPati69JwP/B6xtoQke9rJ3+uylYcviMdMws3kUumUmmHK
IUC5dO5xjgd7R+rwe0JfWtwIJaKJfsX4ekZUxkRYi5Ujki39FsGfDbygPYncT8zI
yBS1Bba+i5xwIDgYuC2PStNpPcx8bjE/3nlmtZHt42Hmp1EP83WCujiVLENRw2+s
QPQlROiOw/bCP+gHH5D8XOwNg23LDgJQBG4lPW86WZ/h4scFCxYK2OseiNIbApTs
tMX7qfRK+IsnPSMdXEt3mQPzrzPAtxbN/MBHmrjhyKV79779nv5YZRxfHMgOEODo
X5B+CZ4m69LO1RmzGo2SaPPkma17aNJq4hs84AlyDHxGmz/QqkY6LLASID8IjSE4
szJmd8+U0zFSoNWhm1xIHKESq2lawQz4U1mcOJp4S7t1XTLXnDkNZsqHSzf5weHh
hOXrjZOofeu9I8FnOv71b5ppLa7sWwkmGRq4fnEiJU57eVoMKR4sSuBHyrcTgNyS
ANW7eXIEawpnJFtYBkdQ6rr3eImwJYqqF6KIylLp08ApbPi4nCjcAeqQzVfNoxJT
aq+Jh5GkPDfJ9xrbOWpcB1kjnlIDdbzm6roNuHVN/gTWQLYBex3uDK/zn0JJY48I
uHwwd77GLNzpMhGYokbjj14gMbX0h95mZN2y5YZmSUegLr+Jia8gUpJ9vuO9NwaK
1mVQB9NsB5F3lX9xFr1k/D1gRPDzYHx/lsLeuEigZNdTxf6je61B6nZV8LIbyAnp
KTV1A79zIWzfOgXFEA7GAUNusMDpaHj3nIwNtjG1wcIDVwFAkFLwsHqsTdwNBA/w
r78VniYZ3qlnpR1py0Zmb5QqBPeMLX/wdjTbsIJlGSEAlK7s6OdnOqHAtZw3tLzS
Fd+5IwJAiUI36YouflUS1iiVOiX9x4/F8g+l+yXy7K82L4JzfwJkLsD1cUJ9dxAh
SeRdkS0kbLBHGGpqUWrPMObRNx5CMP7UIqCc5q42FCF4uN29rfDabujCo/fQvORV
pMItsMmrmwW0Q4ZpW/vdZgAUxxnssYLCWB0La5Z6KYtUjkMEB4/Y/Kx+wfAQT2iZ
e24+JGO5ooQbXi01g2I1xITjtwcP4rdYsJbsIvnFAelYa685HSR+505lFsEeVds9
QbK39GfP09VK6wkq68Gdbj3b6lwtI8vM7rdzq7svnhcSdDuAgXNP3lH7cXmW/4/+
nX+Z6S6Kh+Zth9MXhqmK0+GgYZB3BfW8UGifRCkBgaBtCz2kFSTWUhwOKvgmJ9m4
Z0ket/Rya1pOdNWshFbbaLjf0U072d+WmFP+GZv98L1oe8M4K6XVZaO6yljYGqur
ol6V33KRUZa9KtrOkewXUcSNgX2QOIn80ClWB+tUW6p0ouN/rlj/Ic+xYZnDi/jI
eTZSx3em0KrQ4EyEcNAoYoxrg9IsmnrfWhV6L/HZPxLmAqduDE2X4BrsgRUN5II8
5YAkYH/+7sY2wPLlMAxYMaxOWN655ivCzVLc/QecD/gyHh4wAFiSOBXsAUmsPnXL
3jq63YUrThPPfrtKaQJbruraBIVdddAk/Z/Y6Gk5wpi4d8mqzbbJNdIl7MuKx1hH
XI9QBUlSKQ2FRP5vMFdIy6xiHGV9uFyClXeCMGLHgnRV1ZzmmdswXHo9fNDrZn6a
e+QJPkLv9EFGEoP4hszcbWXFxYn2R8Yifpmzb0U7WNDq5iKLC1rPtX88+1nTSBj6
IAP7FiFfffSAL8ghDe9LNvC0hNfU8e07ZlnzQB7siHNl6RC3KLXwYjAa1bFGw5C7
lHPQ9IHaJbnRe6f+9Q8luMpdcGW8RJSfO/2xBfLOnfkGOmAgKtxmDA+S3PNN2zkg
/kerRwIZb+1j1PIyFMeFolmhRM30+GjJdxQployJPSozSgPfAX3eWvwRjWRjQSls
MWSHTAUO3LhsB7D2maH36uhf531ay/jyolAi6G/5tswJZvzotPIsphpCfZEVNmWg
U/y8TWsXT5G4+F+8gDatagk/QFwuonUZQ8G3/xiuI9of2oFQspD8VeGW5OU/7CM/
37CLS6ppPLGR932tzYPwosGtNaqJsrAmpIMH6qJ/zlV1kXsJ6MVhZ1YU9N+FLb6O
P5lvrVI6zSWvOok53zyqMVGI1F6QGpzvPxFeS9Wiz2bKUbPNux0Z7fd23yn01GUX
b1mM/6qRSepAALyLKIhfN+LrF+bt0LVyBiUhejC38UKVuvcTczBrmaowy7/YAWXE
5fpckt80E401kAQ5Fx+5GbPrM5qQk+cRjUGB5rpSjv8iTKgxm7th1iJ/16GZF6va
nfuAI1wFUTEG36ne7EbVJcchr+9fBFBo/rsb2qtBhGV1mGZ3IHOiItGwstasXqdg
Ec0PUIRJqYFv2wxP2wSld+Ecp1c6NeiQefK3aK8iO7mEoXqQcOobi22bfwlaNxzi
qfWUAAWhQEsJbpbZzSqDIVi2+89i7pqhqyynAP4mLfJHvAGiYGWHkHNpWzw6rHNZ
YoczXkRFuCUkhdCTyt4Jlqw81mvXuGiR03BqNzbF7WHu4uWw8myqPBzobR9GTacz
9J7ISPXgpvQqbxDTBCELRM+5Tc6r1NLmOkvX/AUHvIf4EnUcRW4QqFHoWfRO2gyU
+eFVUm5S49Ga+KUH36RxCUsDbLbXbTnWrLELEHwmebb1z1abjsvny77YgtQQLuk4
MaS0k1rJYG5MaMKY+zmRoHzOdFePdOiVBihC3DlrAeolj8fqF0vPGax37Kyl/eDV
9bxIyyob8EcIQeEINUl5/3ktSMAKekaI9kNTs939q1D4FVr6t1lNnhkV4gnWJ5J5
yAnPimO1fYfIkSy3ZixqYR/hUTcLuewZihPqk0KB0C+WjHVwYzzYOsYBnhx8jFeZ
72opVdrSe5vKgGfGwZbjbgCRuZ8DjfrgfK3hR8PIIhmSnp3EDWi7qNqBOuK0c4nD
CfLmuByN61sNmKxBGKJc2eK/IbN/X2X6XIbRKO7/xG2Bk0w/ar9vddqW0TCdAxwb
zeLP4NmFRTtYB5o3Yka2c98cyp5eX8YeUs9gUKSRFYCw72kVSY92+1qQLWW2rGdT
ZEdWbPT4wilL+gdRpU4Upg2M+AhRihBJBjNnTLvKEBgNtk7G32kVm/twBoLurz+r
4IsDI/h8R4EYMVP/DkPw6ouiew7r3mXj2lW6oxC6zzzkon5GdE8wNqIJ5ayPs4Y3
/gkdIO0KWlj+VcTx3Wosc8kRUGm+qp5NCWvxUDAZKymAP5PAaVHF6R9O3+DyFMGh
WE8WKLNHmf63dXCJakylO4Ny9tcczN76r97VmKWHTQ/dbGatUE0L/82dFS0XCJoz
H1P6egiJWEMRTkKuz7e337TSTOluJXOmHcjoZyuGbRhIYOp3MXo0gBk4VoPSwvek
Z/yVKTF8E5NmgyQGi9/eHS4KYG2r0Hpd9RWnjJN31bejBF8RvmR37ueT0WlRsGCG
DzK9i7NAH+t8A9wuY/QrQ0E4nkzICfusSrfF0ZqtcZSSU1NOp9OBai2uhuddOCrc
kLBkrm7r1GxTmL6vgxuX/NVd4jkEJ3dk+eUwFkVXYrYUDRIfr4tHJW65vkFlmRKy
QrxQGapyCDjEausqkavL/P5GY0LnjVbcBTRAPHSRFYPTLr2RD6o0DWF4NZZfzGsU
fd7uh9nYxz+4W0yyB2Xcfj5Kpoeue79Mv+pgyKE/MBp4vEoa3RIhfrAJKpfo9dMQ
avYvjkQsrIlhjzp2g3lYcY0zNshGC3C5K33kfGRfGBjj9yMHvH/Va7fmuh9tHyqS
T4ufOLCcgmkuH1uiJYRYoKR36hgN+boZfIJK/Jl+pK2P2rxOkCVP32JpbpenoqNF
EA+aGkXOoItb5gQueHleQpskH25gNwHRdichU2Y0WaFraw573QhDDag1WFM7a20A
VrqRZZ5g/i0FphrwCdPxy9N+9nk1JtaN2Szfellq5HB0EjOlVCttxYPUCMSVsFoq
UIH2Efdc+ObmD7WIBU0piH4XsoSCO7YNCRjYmQeioplxHoDG0rLrHA6kfPMv9QYr
AxIWm1bYv5kU8ysq7HrzLBrcCD7crIOOqF0cXK6sP6HGCEWiqKCipoJJE/myVYg0
oqkmQrxcIYMkECJWh1/0gyutKYDi3VUbveI8IZWJlxPkdMQaaHvX6azxDMTVP33y
Gzsqu9H6N8j+X89B3/hxEhHxUH2ogr0XubulDpofy6+BktCP79X8SsFPI+jEgvAM
jAAiH1uGDpB3x1tEIDGkXwwcyKTV2gCqKrx8EGPpWgCKW9dRPHomcJrHsAVMyO/3
hPTaFbulIxbRg0O6UwcTufnwSiM7glvrKS+Jl7yc/l5hioj+K/1BnneA+oTCIvP2
WsjvE1BcSctn/2KfH1/Veh+kcnA8GSos/IqT4BJ9Kxm5lhaVfbLBuGmvxb53vUNa
BeMSaZZJPJajraaCKKiUm9fsFD+k1WqdzNu2TPCCn1libPTy56uPPzLzLFEV3xSd
knOSEk9wdtjUjDDeJbaYHSVT4hYo87X8i0k2oeqnPanSpncLeDfuHghVz4Si8vhQ
XxXKmQs7qV7MNpTsNGXKK/CZAiP+w72G8U+b5inYYvviGN1pasFaNASUS9prW9xs
5yKfBqi0XF4Js74qyACE9hlYr8DZrxiy9pugXB1s/VclTSjgqZ/IvMPLblYGY/qB
59WA4OK23tVZOrCCruqxAgAbbBBqb2fHNfpGXV/RYXalKpiKJXic+nDa2kBf1cKE
mlNU7JAfygWNluxZYCVkx75F5d/Q46VCjoxHKo+Z87nL2wIOBTybc1RGumqvG4Ou
aab48JSQ34nGBqi5I6SPrtZsePbll4QvBBiT8ImcQkvuoikB93DCM3YQq8bez+5O
xyKHxmE7GGrRHd5UJYMBaLIJUglPSNrZDH7g+Shn46vAkTVR5ctuoKgFZ8VJGu+k
u9IDig0/ZqYiVUdJNNA76ANwbDPuKvEO/7FXTCORWVl8gnEehYFjLcrrwuPm2Zm9
yVPKXUbktbt14BJ7pvafjxihKxxdWSEJEnDVTvhY6iwzy16zTc6TqxMqSnm9fi2e
fgnuPpMNAbYidhrQbGagAD3BYi5ptdBq3a6UqqVBBkfpr7aWe3Ca5bOpDQxcqLNH
1D+eoMrIcpJW+WyF4sdXQvBJQ/zLb0nzFI5Db6i9bgOyqjSz1MQmXZMaBeK/OMlc
r6fvUyPblE/VIf+yz/KFNcbR3QlM7rfeGBZkxjg1UH25WeS9FMi9MWjRQG5q+PNs
S1ZVHzgMPB/f3WBce7WlcEFu+XIaLVl3aEKtQYMcRYD5FjjqVCusX6vflG1oMHfB
OSEICqOw2ZxbA6UEUIK/3XrOmlKPxSRmkLGoOAVRcU1sUsrVGxkABV5zqh+qwsN4
2Bqe4JzqkSzfeJkqkAGymNQm2KQJ6z/jtY7kINZWQNz0jOUV2oEf8NiNt6NrPo/V
oPQ539PBpOVqC7e/IFKZAXt6HAvKpI3cLOXBi0GNT0qSYGOKdo0V8EqyqByl0A7X
m5VOeF+FPW9sVJxm2Pdiy+nRAr6r9YtMYyMpryNKwNyu23br5Cf+HJ67PpYLEZtg
ewF/KNjbhejVIFlRlWZJWHziW7PAe1g5NwXL2p3XQ0pcRVgMRJ3iNtMiyemh3nrJ
QhfVAm3zAbi1zrVZsqbLWEZMYrlw/FJMPJ4vvk8s0Z34Mb7sEtk6EX4CthnpDXBd
MKkpI+6Etb6Fo3NWkjJNGN76IDWedC7PNZfdzHB+1j4kPzO2NTwj2OHSJRpun3il
Gevs5dC/7hzY7U9/R5iKXS5ehAznUIyfXpq5J4v0f6v6g15CH2OPsZd+1t45iojY
Ya5eCxLkkaOB1ReQtmGwQpxel11GHdDC2xNcnkjksmj5fpi4+JBfimfUxQ7SVR4i
4ZcDo2RG9ylu+M7gF2NQctx5Sk7BJ91KcEVuwTxgZDbNdrnG0bekV/Ec0ZoHmiN3
3/MppAEJbDA5M2gTO6EJcDvajolsOC4N+TDXvAW40QsumU0gte2veKz05Iicmh4E
G9wvbYUtsXy3f7WEewWW/vvHM3lJB14CZvx1MvtrH22HR6yaflKlPCtSx84JEpKM
7raSSyJpicdaJNlZaIZgtA2sYQ3F7V3OdZP0HnwqunHE3gshsrVjDuoQN9Mr1b5k
1Uxh5FI0EhVkAUi6/o5nj5YAdqotZTu0eFKPv5XwS1SiFBcyYvnCdb9G40Q6IHxd
DNcpRJJLLRiONnj9ymbPKlHykb8QygL3CBROa1bGGUZFZUlgI/c+Bw1s8u2LY1Ji
nMyIyT7x7Hpx2cUDyD04iRGlOudADxDM4a9iDplxv9YGEDuQvvNC9h2d62fq5C0/
JoBUQUiJNap8PJYxtumtjWuPVPKoqOgN6cQ4xS/XkJXCmJhvsHpIIXhDYf89cpOU
D60kuPQPhKAqKeWAPTTRc/ttBeVa9YWR7AsN6B7RvF+fmbtMh3v49O8+ahrRzHn+
VEH9dvhWKiCTJIJHihmDt2GWWTi9SM8X43+uYaUAIjq8FrmrdoDXJ6+SsQwFUj/0
rk6sJHP/XQ89LbSC7uBO6rZhhDhswwc9R7gyYVhnzR2U344b9Wefv9D+G1cFzMCG
hBC3sGHbcb/sFtg9spY/2uFcE/qxdrcXr8z6Jo036qdorbuE/+xDV5k/6RMftRSv
1MSEQlZQjVshk9pMxsRYRkivNpOTupYeXFhyQk8EZmSrXlKHfqQchyKJ5FORT/M6
W7Y/3MJC4kLNMiaYO9sdjXOtDl807Y+E/v4ld2sekE5VgDMchWkIJ4bWJ8+nDWG4
5lgFptte1cEfRNZwU6G1WMr/sCeBMAFxNbVLxTN0ReRMyJWAXKKSc0xUvrQSk3bH
RNLwB7JyUUh18dhjxHj8o/44EXTa79ZJBgFC+OipXrgDsI3+17eu29pMWPAqnN/G
FI0BPsPvfBbod65UbDtRF8ytAILL7ys4kSntZUYtdodVK9bFyy3sg7w8Ney/NJ6C
D4nWmxLCcikFQ8O6rHsHaig/dP9ALVt3lEqZQrD9OKXrPgzH/x6aYRfsuW0bEErl
lMlQCu5qmV1Rmol9VfJXGHsaIz+hsOEZ1z5ghegykrp4W7WohWl3FSefS41CyXfT
/y8EiTLQqueeT7S7lt0kRAxAFFhTCgENIMycZ7BY1H/Rkza4a+dTXIn4P6yWVsF0
ptt9SSo4inwrqGBngkgKKWEnF/AQAiYZlTbfE3noS/fo3/HuMOw+HG3/PZ29r2zS
nZ0w4O9wqWnxSkYfSi63X/JMZrJAbB+p/kRMv6k8VJpi6mxO/VN2pF3CPd+U4kL2
hDjh1Lo0931iSeLQ+w25OLpskbfztDSKUrRimprpCeyuIUU0XapGLCH5QfpIb2jD
bidLF5tcpvJcG9MGKFv/BrGJkT2hQvvJbvqeE/9xJn9ErKnU3H96gsEt/Zd5el1U
/kYDrOYh80TpFyexkrEPqqPH5l9BMP4zfsjYg75LqZ6gtq2DHuOGGqu/RA2Qs8Ne
VI+XIUTM100s1wGwqxN/0C7w0rg/VaqL9T1/Sek2Qc0AFDXMkr1zpm3WXbrSMdUX
U8+wFcgNffAEXSk/MDX+3sOTvxLYV7Jqt5vi4v14hevPQoR3ZMfTSE0luKf24Sm1
OWs4QpN5uji3CUyTbkbPxJe0DgwF+oihS0nxoXEx/ws/Gy2EwFB5M0pCQpO0GO2T
Z71v4zw3KUKEw0bVuEMu9itZrGcgyNs4EeHb1Dz29yu1/gv0l4eqJbgjqtn0HZNW
ppqAx8fQWZj0dpc2BACnEvd41pSk2ZAvaXpU6ThD4leNE9Xi/0ajIbZKE1tNhhX9
`protect END_PROTECTED
