`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Yw9TuzUjSiiJNoqlx/x+ib/mnTBBmQmwb0ch3x9s3O5fqdGOmSW///32IlbXjyK
X73D6pP9MJEX+H5XvP58xQXYSuNMaUF0DscKfDshc84Xlv05rIzW3+gnFeKzGHKv
Scu1q/JubL+C6IbgLZQp+c0luBJtUIB3gtoQtq4FlcDNmI2QgUQ0RwTnrvGHCXc6
TDOhof1TmOuZkCFke58I1IMUmcUn07xq1CVWP4AdWx+IoLQ4MNy2JU3xA5n7VWjD
ZUpZSLzJ9H0G+PSdEl1hkq7gmPOievQdNaROiO3U1YHPjkc+9ff6dT0OYreEu+9u
x2u4G0Tyt3VUpp48bN4QWOxTILjAvt6zE4PODaTy5sd2SsJDAnLIbo7zKNnYAae6
CO4gUiuL6hL4KUq3JNhrfZEE1KxiU3+1SL0gXttUPsOl99xiMIw9vUoTV36/h1a3
xh/0P9XruCD0WKSELKEo4y1amtXhTEdIIxLdaTyqSIbo5YEj/DGjYWrT15mR3dar
fnvH785FBXt0bwZCkHNbmRaig9zEXidwix8Jd/vHQ5oirUYutKNpGcg/ICj2tnuI
QD7FjtPrZMpgb6B5hbJIkvz32rxdq4P05VfSic5y7z5AaNRjJR1WuV877WM4EJ9J
GvvO9keZKzVgysCI2MR+I0XP2eW5AWQqhE7QW0/sclhS5IUCCUsDAjleDN9flhz1
r+070gUs8AJyr9DpjQMwUYrPMyKYpf4Y4AbM+2eRXZRztvSajNhhve3VYtys8A5A
i79/XI/4m6XTkU3GFcjf0IIeIt7W+rFUSYH+OXZSAWEKOgYgC/ZcDuC/13xkWREC
20ZZaIhgW0ovdoQgUlmDxGnVHFJojyViAKNhTKPTHMP8v1WsfAM7O/G/LL+vePG4
`protect END_PROTECTED
