`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dq0TtHF+dtQtoTiRgEC8UmeU9YPUlSEVo/FYmynBa09B/tdU0SleUge+1zm5xdmq
5IfZNZdAFmZb4RzL3/+Nan5FLH+4ACTTxSSjjr/4i6n5p1YPjSJDt5/tfYVuvK5Y
JJpL/W0HE8cnfOkvEQqFYIFZp5Zwru0VlK+Jr32HBgG3bnGO1ALqLfAuFxBjmfrA
GWHe77UU//B5FVTHGlNuEyKZ3DtwaX3TGo/pEO4+Z8UE1rD9v5Dv7GBd88mxBFX8
0HOM2LRJ3X2H5pujROdvqsOSKeCjbMPXmndeHVhl0cLpBUkAJGGERBfJQ9/fAoS1
THSggIkVvBWv8L1Hw3/mUoA86L4ra5bcXhL2x2KgfeyI+2so+wlxE6j2GuXfKGX2
/DXDja9gRr4Zy5f7UjYqi+OV+upt8uCeQxovbEpv7mdE1mTtimYTO31aU+SQtbjL
tI/3rP/h4JdWvm3+8JJwxA==
`protect END_PROTECTED
