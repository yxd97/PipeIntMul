`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g02jPIjCH4dNXIh8GJ+LIgZulfMylxqIcbm1djUEp2Yy/4kN2GV5YOU9jq7N9umz
J7hu1g/9qbezSymxPTkx1yt1t3I4OO2Ifm3SXhYgVvElX80uXjsAjQyfRib2nJaG
fwtXygeWuxWFwF0olhTNk5IGtmnDv95hgBNNQ0d8KndIJrafalJxI+BbWT4QeVtL
upyjhzs0OghnfCVWGYW4MclnkZ2tj9bnfzoQR3MbWCodIDawac6tPUbtFI8bpaRK
w0rsImHMEr5mfCGES0nAUc8hLHc/wpx92V9AfN8nJzqSvvA+VubuJ9zXIqIge5vb
c5HCCLBuStN0nyHlKiLjnNMN4O0Uh7nXoDfV9gjYmyfIbV+oG8IocxbcRrTdeEDe
`protect END_PROTECTED
