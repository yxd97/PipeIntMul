`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1O8AjoeasJEQFevpF+3sbeL2YbML7ynaVZ1sN8z7j0YbYmcrkYMo0bVQhciFtWJ
elFpZ5746U5ApEkjXUOE2ABkKDWKayJW/IODcn3/Hql9zqgyhXBP/dbbRLBN8fUS
DrGUKPWybz666+RPG7GUGKrkULqC36yKhaVBn69Di/jpMglVRmGM+uF+Btno0bEY
tvwINmh60qucZ/6lS4YzGiM+zmEbekrBIK+pSJ70I7tRpbAv5Bsabvx5vaj/LC6s
6bJtcXJ60ByG6Ca9bwRA0CvcXBRjv8lSIsCO6HrWhuyDDMDTJpE41vZox5HoK1Tb
ApFCgc1rTNaWPDaWd57Su4CJOcLOXSd83WgczbsC7Wp0unSXuHlwer18pTF/gObb
7+IVxxRDStNZY2jUSLhgGi2fQ79icOf0tLkeiQwXy+k=
`protect END_PROTECTED
