`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evD36ge3kbP/PvsAa6EUPI8o73C4Te1kAO9xJ8OyJYdxDvlwNPXy1vmonWgQBPuw
dMZa6VKLpcc7m6Py2n2oj/V9CZGja9FFr7gsbsG7rOHwupPzuaoKAH0BH+rcfxWb
s8wQdYcg+AWEVAqnfQM4UbeDltGpTQBqZ4gEt89S8NGijeWsieLtgNwi+m3mOVoI
sxlQHXhi1/VwtT0PWuYWEj6z4HBIKK7Y3JXbrKO3dl5PxqpCITopG0oq/lB8/acb
PyS4Lnyuec5vcOWUc06fdHJwoeZ5HSSEGoxE5CMZ4PJ7s8/feL9d8S2rzElvucrp
IZUvOyk8uc6WqiTKe20JRR+l2LJS8WWHZ9XPru0ehgkzBlatnp14S2deX9wLYjrP
1PjMKYpfFCviBR88M7niiwRrK6wGYlF0FD+C/vM7AiP/LumxrJw1DbsALHFtEWn/
`protect END_PROTECTED
