`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
snlBQP5Mf0Ch7QXw4Zaz11CZ7kmRea392lFYp9uDLeVZo0c6UWKGxusklxs69fTw
14mlu7UUuMVnIPwHTvsuua5xuCDBSZMAi3bRqQLdxm0IxHYGePiQzIVkd0c05ZSg
9XU8ekw7r90uGm3MbT4Ep2mvgsyDpZe7JpitinRnTLLFpfM69er1wEtpeTulOXQn
kpl1kakysDshySFY0GpZGxuB+LmZ8Phe0oXTPWlpvn8jeDhjskZgCIpNhuKx3/NA
wVS07sCbyqELxqZ7QYnFoZaYvsmdB30GLz8U08dBfXVnGVBudkmRDWAKyKagkpzr
XvXQyMsFFhH1Ju4KmwUS2gjU9Zx8L5emBhm8V91is0H7Yv0uidyi411QZTfktZzE
KYzYVrm4KF7exFjDOrNe6Lpv08WRnMgg+KZcvlgXrXM4D+LKgdxVjBe1ninwXT+7
0ze8NwC/oY/at0gSaR3IGMoAuwK1f7i0FPMblTvyOOgZ7bw5NFbQEMJjN3+og9ab
e8tXfDUdI8kDKbSwWeli5PZncdwJWC6Mkxz980C3nDVueOH4sX3R7vRE6mCcf7Xp
zzKcsqBYfQAUtdnUZZUtyYpslxAd1DPuW+aBtko3RykxqrifYHEjq/GXHlWz5klD
xjub0RRevBW1l56xXIMDiiKVhqz7OaZjAJM34ceyJD62oUjw10QCW8V6PYtL1Tpv
npWUeGrm4JGdzCGJU9Yyy5VflzdI649qSDiMBtBuLHer5iggKVawTZJBm6wjCHGz
ZBrdVMAfdFadUuZ26YWl4w==
`protect END_PROTECTED
