`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IwwXR3ed20TADjBZulzr4tUX+Ie/m3byhnBV/RP7zFPZN4cXTOBFqHdzqISoAJKw
3FhJmApdVsbsrOCR9L0zPLnV6+4wpe0vzKnbGIjsOd1ZqRwroTY9t9K/QZ+oriAc
VmhMncfcf0IvHX2bqj8Ut+Zd9YI1XaFUAEiGMLAF82QIGAntla+sXvS4aBFixhy2
apapAIrBjPBmmexyxuuhkjtmoZaCmIXMlLKp8XFA2RqTmA0mu2QVAebvoTwbHoil
dTraJ4q3n5kBkQSgzmGnnoqISKDBBvQ8esNEybrptjKW4ukDwH5cgab/daByTRtc
CvAJjcFwjkz7CsJxHzOZk9/HeH5cHr5Z+a55yEvhS28nFgMjR4MJfDcnp+dcs919
AEfAp+FSDL+lOiA4GKdlus9rkNuwha2dS/Z8mNc3NX9cEEBR53oPlRq0OCygT9jY
pfMejiVJX1ORZJsRzvAYLWai60cZjsmZdwmsHfNfTpeLmHQYAsVrgbWJhlJlccAy
vaY7FBN/bt8enOI3ika+7w/o7kqwTV4aIy/9c7vSDlfdYgjl8+QxFiv7hhlTgciw
TC7KL28mQOD+gm8bH30Y1doF8Na4OPvXOUaQ5nPb9YUDKUB7zf//DDYMDaV6mB7t
1NrjbebWfyxEA/nkvjqmJobPNEOg8qaCdftdrDnSvUceW0tbtj4ka9qndKhQDCNT
Vr6UD5ln2ado3jOaSG14hscppWIHmhwPrSGe/wy0RY5hFCKsj1QS1CCn4LUQbpXS
XVySq4Yg3CSFJv/NCXCjI2gfPQkC5Z81nXFklR4miwNTUIKyDIxCS8hfPcIMIZRQ
FkWigvYnJi1P4eBJESG+0k3v233idxWNU/BcXGR13jCzbHxcH2unvkpOA+TJ74B1
aYoPg/knX6kT2qx+4FURdPpc5u9YaBotee214QQ9oZ6T2Q0f0oC/K7/NspZzoPY9
dp3nVza1tDsvLc6jdZ3+y2rzbp27gfTtuu0k+7jyPIKsXnjVyodXAR09dIJbpvah
ezM7f3PWFR9c4t38IeIe3KhEc8mHJO33C8BLc245SA8qecAHTQacGziSTkeld+W4
Qt8uqdJrfLue1WayuJCe+tDSFyG9N66/OrM6e8w7lenn2r07vjC7qI1EKUFvh091
yqPS0QfdXz2grOLyDlOGiqHqyJOAzzxTZ4XhButUrz26bcsvCc+AbZN1DatB/MEN
4kqMrZG2ZDn9x7tgSCah8V3l1TpWOpMYT96sPDvMqb4tMzz9U4GtSXevlgPJchHN
UhcIlW5FF2wMAHQk0COoguIKt+WepKML74i8h76dXiUwASgARK2Hh3PP0SS4w+JK
cjbl4Oxg32964fOTGfCocpzInzqE8hWWTNYpTT0b9sGUe1AC7QkbU5Ls/0HxGTzp
Gwuy8gtBMurkYZ50z7PoxUCrHdWM3HiF4Nq/7wlOIkdxaYsqxSN/sKJPuH+bmYBs
bivt5lnX8TrSK0MVS8Gul5jl79XJ05FSagc8Cmy3jtwEODMZbxYfSk+J79B06uRA
vbO2ubuuAkxLu6/kPnvCM8o6+HhbMRufdvYi5EcKqrdz+mt+bydCkAvQ2bBSmEbq
9hxsuZwPVrGFRPsPIFDv8zKH6mmDlbcmklvfkmsQVb31m3VqJwZHfKfVzROz2g5b
hgzaYbGVjaL5SdXVTpkCgE88ibEPTUHCjDmA7MJzMOn5WOfHGWBf4o4FfbyZBRSc
3IeU4zy7gqMGLLuwWeizYGVaivGW4u4sEUh5dIJf+Lbe5W48uNfiluUQd7xJnExn
WkeDWcCXs/aHhOoN5y2g2nmvtMEexKmgso9jVlTRcFWfFoych0YtPfjxHwWhVxcE
byVq9rMsRKOYOVo73c6G7+vKmRPteVSIUz0d58TWHMajgEjKdBATaOLDamSdH122
25GV/3Gst8jKSR9BjTO7vKStuJrAoZhUeOHVG4olGiN8HMcWHx8vjYVzI5de1QmM
RIAa5v/mPidv5PG8zkOYHiBOiOLZBwo7vgc2Cv2RwqIYmQcq+ecPQTgxIc2BtzUj
lyqKg81slFM9J5wzUsFu2PLJjqAzIB16tRWweosU3JKMjOhuFSOlnXq/IJ2i/M5B
k2pOSBgQdTCmQ7xhcjjHIq2CqIv66CTp4o+5c0dWYSKe5xPnxW+lXmpJkQRSDWWY
GREPpXMQNGRzEMt0A+CUtAJ8k0x/M9nb0UkYPDA+ive6fRKmVsJQwbm0CuvwYEBo
QjaQO8Au92a8aOfgXocoL0bVjEK5Ljpc6YMKjygmfDEh66whgI1pA0LK+kLbbdjK
XImAf6QasUmJWQ3MD21WVjBpp1/CNJ0IdlWPsikL+HjTobRUvLOJNH6R1c/JTCtI
+eFoU1BnK8E8uCnkJBVRfz41oDo8lwV98EIHdgfPpU7moXjlStkyZwx8b47lW7qL
5YUsoxVUA7xcypi/E7rUmRPAfnHT2MjvpU2KpGidIJRIInlPKdb4mFW52veEtO1u
ZZv/8m+9O2Ppfn7j5HAer0Rt/u4TOx6KEFVWOqsWA2vF46Zz3JrsObpKXDHjy099
PSnHT7l36Wz5L9CrGF7UNafJUnyePMF7Pm4Fas4ZvoHZEhNKxFYmAWEd9of75uXR
WQhOLEF5q+3rWBg401V9FcqZCeXzXHjHrD2XEhRDCLDPnvJUd155H/UuD9BZLM4X
8lMdYjCHwdxA8ChVidyPtjBxeaSsnDnaPekmrQ9BTy7mzB60nJmQQAFDnLkt+ZsW
iepbquwhV62ERSq9NQKwh0JUKni4U2nPUlednK4DM43GXSvl/09twHCR+9aUGwHr
6H/z8HeMQ+8BV0NPp3iJzngLZtZecETm5Nt2jZMhsvNkIWyjA/Poo3eIRhtg6vX9
HuJPGtFawoWaKun130ynArJT5LGI0v7eqC7nnPudIWVm9DbhbvjHOnSP6OwBRB6T
YpUx9SiI+0CQTmn/5xicv0PrerCvCafCe53ot5ipi0vCB6pRMmOlZtz6ujen+Zab
7/RrCr9RBwrtPcWEml42wZEoG7oHX1aMdbe4626B2CptweR+CBw2ZI2meGOy9v63
BwbN4TN5ccgB3CffThOts5i8DmofxU7b6O7d9eyncDbqO0hu5EGZNCubIBI9dD9j
BHWPbKT2JPTyqUf930+EzdE2IqJQp54AW+6JhgqJXjZqwXhYhiVeJRo53tcJsDMq
P+7btnKPzXkhY+Ld/AWbYiayg53n1oABgsIeeLYGO2f5h3N/sj7+nfdci/JndgdP
sD10Vpo8mQtbdrhOlEfT+4hNNE3av6BkMbJCMMyNJMdnt/1U5dJSmiVKOv3VoSpK
y3LcXCwUZmhvSft3bCjdbgQ2fkUBma3HA0bUy4j4/w6HPK7uqqFEGF2gOb8+7kkr
zKMtZZ0LUEC28Z6caSoe6UIkYFKgO1m8RZjRv9/jPZfk4s9Zv1VyKGb0oLRgfKnF
MUBEYzJCjv7PD+tzc3WkZJuoaHQswGbJwanwvJ2uJNerLuV5rWIcdrhGYm2FSUoL
p02DWjQe8Le8pIfXCcgR6BjLtnPCw+X819ZqiLQWDg0xQUa8PNHE6jd3L9NtHGKP
TTG6VdMOpPdeasFWW9/GU4Uw0wyhjZNwrygQ2U5a248Qjlpmbnen+k7kftQZQWne
Z9xtsIf3y9C77SKM5H0uRWbKVbQt5eAQEqEQaYqXT3o=
`protect END_PROTECTED
