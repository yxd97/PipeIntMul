`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqJo0sGvQMgowfbnNp5HrQRCoDRzpw5Joc00HLJpPH7J9NfZjfJbzy/kppFIXrTK
agEXLbogTQzBf+e1c6198KAfveTzdvpRDBzwS/P/cVgALvRMWk42Qiu4BxYOf0th
GOZaCA1BhXXNIO+m3m3x3UT6uhOxy1HMhZNsFH1FC2wQ+T2leGtgcgpLCZbP93Ry
2+aggDugTr2xod08rD1yNAkCDgqF2gIzB+OUU39F/KCUNU8aZuEnAiuE07A4Wqrx
hB4T1dLUEexL7hrQDjxjoDOl/UHrOWncZb2Z2uGodREiWfRpSsYFvkQvdXgiEgBj
+hEmS15agujhJc3RhxIGUeP+UTjbC1lUs46SRsQtJl8IKc+QHLonTT1s74qtZoCu
HOdh1XP3x37ZQJ/PQLA+djCTgIC5rkw6EzTTEeOCvflKpugtLY1Zo7guf9vdcHkO
xSbxGrDvIn80oO7Ue1+ALzo/PKXrpqCL4jrwtxTEHPNwDaMiDDGsPRStw3U0ZS2Q
0/1PgvxdnPGxbP96/RcfSJ1f8GdzwMhdAixDAkUa7vNfBiR1F+OqbBz1mf9HKMyz
tIEfmrOKGbHbM89nZ3jGakZQuV1UjdRc0YYaH5nNgU6dMYasGe/7G3brIXGrors9
17npRRSGNDJ7qSeI6iCTuof2ae2B8GAdigjYsMKXJLeszhJhk7kw4pU8slBihD0c
L6OWGVnzzbkGnI29cayzmbCcy+3XM9RtA6D6TViYBuA/K8YLxFnVWKeC8eB8F/kE
j42r6aZVpIQmXRYSy/KOeWPYhtWYL9GiUDklPWJOnGU=
`protect END_PROTECTED
