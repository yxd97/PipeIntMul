`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRwG41bBCW0LUddr92n81g1xk5edDCZSOP8igK0qKmR2KrEBbp/LGzZFZuG9+fyG
+PtzlLxk12/gP0LscBMnUp6uSuPU3+CXHB4IShpQGZZK/q/XdtJxgn80wUDJqiy9
pL//fgojhcyEax7nL6UWVsXQfotHYQnyljyd/cKfVhGKvVLfERpq6JDSr/v7lQD8
73krXhMTXreqIn6b4xX9Tqlk4uGkDNNtxqCuru9TMM+0Sbgs5XvivGVVzvNLVqEB
ibKkFPi8q0BIUBF3TU5RUojUkF7We9JTpLV+Pw8XOHis2u5ODRA22BhJ2iXvqONX
BvJLQzE9ViIG3g3bkJYBvHtq0x9lZqZzemh2abHhIOJPaPaVtNukSbTjwZx6q5oG
CinaYi3UYCKnnc+JzDM+oODmNgiAwFNxRXoJPXRZtfA+toJsUf45Xqjlb1cYh9Xh
7yn6qvBcuz5VJy/G5dBM7+tynITc7+/+I9M0ndTGv6tLR18CwKG3TpmF5Ztuy0aK
uBpRJhn3bONO9Rct8tNuMkrdPYBoi99mW6h62pSUlvpVakQ7shrVywuJ5gxJzXrl
FzEOSitM7NvZqqqDJ1/3uk4ssy1qPVKdrhfVmJuXoGGN+aQb9WhJoBf64UrtxV4A
wu/Ol2vgJJvf/7CzaSpKBFddg2ERmTSQgNH8uCek3i2rgaVwksL2FvTzIlzKwheG
MvLQBix1QDF0iWaKy5kM6mynzf0fGVdCRB8fa7/pvcZnGROw8ObETRO69BVKsmeO
3gViWw+WWrFC7dLYuMmZVkvcmhXn+GPBgrptDkVE9K/c/TN3pvgQ39M4U949DrjG
ZzjMa4nSZyiMdsV/rDBvk+8NnzID+ehiBawU2uNBA/zj22IPYFn/M4veNxfc4WTE
uh+dwfqeR/WFr6cwQH4J2dwjnfpaFAJBh140MDkqvD/iLYdZFKI7cVTmysV/nDp0
DSlViPcw/e89cr/BCcWVrk8dpsAZy5BL1DTZRcENlUfgJfsIOWlNmO3W/LHii8cf
siybd6+OyFzL144tDsxcuu7dPB2JjX4JaAjvUAF0OSMGD4nCL6htKcMgDQ9EvkSn
q6AOIpWFv05yh24H8ejVCajl2Kh0d6es6+Njh4ixKgUrQNqzbho63tYSd0icXVFz
n+Niw1Mcbof7kdImIrX5wPDBsJcqbpEWhYahBUM/pzFsIryAwuv4SQ7eeYqwwSNa
y8+fmDJcA1NAn49kGZey4H4ToPKdjdGPB3fosLw2mjaZ0tHgzv40e0kCDFb2MHbU
2qa2JPVh115CS2diGXASQFqlICdB1UKatmqwyCp8t/Gp08wcQUqYmf9q7Or6N2iu
F/AKrVmyB2RPGKgp5g/XMXsLA2ifTSf2tcO6nMKx6epqndvhkZjZx5eM1EoTW/g7
DMAPiiMXYFv3ZqxLziViUz2+5uVHvDMvRQZaxecEZgmXcIVQ9UzdYhSQovqAbJvm
CuSWQyivrUoHBvy6ECreTQVwPECw/ULryjiiHuQT18qZC87VAhAVzAB1ZC+kR17i
sHCtfhBO0coon4kD0z6dB9g85OAhPnOETnjKpNUV5eXGoklo4M0eHyHeamcM0yJL
yLvWsaKH/oeq+3XkevSBR9+WDqYrdKhWC1sO5Cbygc2RRsMHXE1T1V41NGS96MAH
vUTwg6yG/E2ErySCO+5f+J+wvG26Hhcb/XTYiKX+imM8prc8pZV23tgWXw6UdO4N
dOHiR9AcxsKEtejKh30IqwkxFJAlE2BAco2oTxqtoZkOT2OgHcEKZ8SjyXffs+c3
o2MPd/mQcx29pzkyleZh2d5YXP8SeIbuO7kCnrKswC72wOikGdGTvgrfXuIuqfUW
srIqDvwjwequfBwZ2t6mXBSfHVrkdKpxdWVsmmKV2ZwsuFq4yvXsKIL9JvtE6nXX
PaDmv7E4SsUIEpISrS71bM9wlytJxEnu4G1FPjbYVp27xKQSP9Di5+kNr8jWCvEY
gBrVdvcEQKkSRJSq9VnbNjs8o3x9rHDC22gazBPK029KW7vDilfAQGKN0Q5ICGgZ
wY28ooYn36lzVqojn3/w5ZLLO8CLE1l/JmxUoUDrMWEeuwkpZApGOjDlFShtHHYd
ujhNyjnE67nQhqQq+P8NjgoXi4wdWzVtbMHjLKItF81W+9K3FDB/R/N1wZ6QEb2j
DJmusrGvq4gZUMDWSonmDr7fL3xNc1EWbeyspghonDKohwEGFPo/ifQG+LR7nhNm
1W8JOS1ptaD8EZSxIfdK2n6GyeWnCdBN1sd+sv/9ycvsdRXG1Tqi+d787mikutVi
trXrVdKnRTrPQ8NTdCQaCXvU+m1nChUaFrl+FNZ5NKhIT3nUi8zasqjKuCHxucdO
WqQayT/+dMZCUUFxvzGAjkC8/nTPKlaDt/KEVMrg04ETU8V8r7GKRw+HNRyc4CiP
LtKyQ+GZprFm1hIvLdZTaPNzhefRsrGvabs7OlgKzeO/lcv5o73zr9x1sNh3Nfvj
EVL+XGRtkzrhDmANil8lfymu4EOd5ZM1AkL3/e7n+jkDYv4q1RWUQ231g19euco2
xwxlIVARoiNkRaH2VeD3VfASNZ6ifJWIVMe5HPzj2ANv0i46yYPF172rqwFCSYs9
U/WPzyfCN0e7gAiIXKdzINZc1i4ogMf2J1qIC1O1joK98T1OJfsXsrgJeL0xSJRP
QmgPJRaHl9oBqiFkhTP+S3z2uMQWMkPHc1yLIvfkCfDqrWzp9vQ1esb5hPM4CS/e
ccuD7iGzL83NNaYCrEjHK3voEWo1DFwuEh5ZjVmv05A4I9WZ3BPDgYjStpylzOb2
SJyxqHwbsWI8cVyjgfvJNegBr9j+A0C+LdSzVSBvUO0c9XHN/NlrLdrCsAltvnDB
9tGMoBSQ+dq5p2K1uz+iRnYnns0UX3ZShK6ovIK6hZ5nt04B/uLxczfBwYUx4isL
PPa2Q+s1rynD7XZ4vH8MCfkt1epzwJfc0s3kiCveGE1A5+OQDtotXw9ldDNTm+UL
9RwOn7CA2R9aM9AMqpr7pzZFq48wWGrz12EDwiE0JdT82WVIf1W56+9po0ablf36
odH1384Lp040B3tYRF49Jl73/SvZKA42aFwL1uHF7tGy83RkIBNy4V865hsPb3yb
Uh7rNfLYLUOXWex5wBsyJD0vSdR5wk89WkJKyRryIjZjmF3+mMz6dorgXd6mFL/w
RvDA71OQkdq1AwvUFD+AYa9tO0Jiy8d1hDQ6RV91ZFvF0O5Z57mBA/umcd63EiN2
G6TZAIW9nriwy476hDlvJyypike+/iTC/lKGH5dAwuH2wKWs4FxHacCOe7l+pEhE
PtMdEWYWk6YOloH9C624QmTgZ7X6kjjBPw77CX6U1buGyuXH2brw9H/n+AaehqSj
KFh+VRGLt6rADDubW3Myylop/4e6/rSH5quexRdLA7UlPvQpFZ/i8BQfPWouXplW
m+vE0BeNAcp4+NnIqGa7qy8/sxADBj7/EHfh8rv48ta8r87nCNvpwlDe9Jt3co32
XeYA6vGsdURld5vVeoQjxvVGC5i+hktcfB+To15fAK519bunmO05yUllRjKLOa/a
J7LJdD3pKITELcE2EqaGo38Oe8RMbUWdRbpPWWHWMO5PMHbYU+7WbHKaiaLe8nsb
lhPYbfsgUPMjHkyBdM7PztAyKRX3/u8sNKmDpJqNnT1jyl7Xp7aD5Etc9/5pGut3
s1/K/cQmvEqH07azNiFMITYqXPz8C5ceM9VomHYHoH2V383uNtoEcCJHS42jdKCk
J6KYfiYA1ZEiQmn7/uYt7xem+/Cef13PV/O6qIGdaL9fkGT6Cvp5Jmjdgnat780n
+gnCS+W4xROwfzsSYsHoE/K9hWF1AoIyp8I7AIgpxAxOkylcUiMlyuFt/3dRPiZJ
A4jJbyxbF2Kkkmp8PZekqhp2pjH6F1N9uc2HQgJRfD1eaFvuPmRfI3MQTYKApyFd
g3D+XCut4eK/qxk+Illj8GmGTUlFroKSDOayoF0Svd0E97g0sCkw6PRkZ1zrhGyU
r0E97GFDoZTLpi95kNz2TCtw93crGAuKj28AFnHYxKr0NrSvVH7xUWrwkeI/VxCH
7KqZ3HY3OFunJtkTXMp3I4+FRT/W9Efm99wJhY9Y/WR+7oQ/ZDnYCRiPAuDMCE41
LHll/CU5lTnioOzFL/kBfyNk3/b+BAYrv1mEgHyeGUiL6dNSPLPP7K8UydGT1mZu
QngHaDwntHcuVuDRA7X7eQT9m2KIsopci/CtNBsZCXQaAoYBGepQ1U/7VF1Nl75S
rHls7sjK572+7N2XEFZ/AiQkF5wImM+L4tai1dS22AMc55ZWMcc4abNLP5/hPk8L
q2jX9fSvxu/1Dtqbvyk+ezYU0broNkdhlaS3OKAMAarADGm+LR6cGGrVh472SyQC
wTuG8ASjmdX6839yyQdcjKlqw105mWs/XjXGrZ+dIPo8/pR+8IjKttAmItyIxu1I
YeHil/l8ambLIgcxbeB8LKTLQ2Qe9NnTMk/h6yYOW0nKkKuU0D0sYEPmdOx/4duz
o3ri4nt0XV+sM/t+AL6y25m/+bIj72hWcTaryWQ1oJoVgPnZ3AtQBG8jcSS6kjz7
AluQzKYZmvdkYIgEjh0Q7s0m8u7C5Q7VK+tWwcsytVe+srWKJrNobf5Cg5JO7DHt
JdjEp/bACmhJEVB0YoEpb3PaKtOQHrcSbhz2PbRQPqlk+IQUSYNxmCfkfcemqRmr
MKGD/6ubXUS49gZazP94fJI0jZaF9S50iHcKKIawX0LFF4pC+69pcCVsKOn3n+9W
rwo5tpmUxog02YamoxUI8fXxqp9/Lowrtg8Z/t/2jHKjYxHuh8HEZXWaOF9CjMpl
JZrHBnNtBnoex3NTlnYOGCi2nXETKbmud8g1Y5yfWILeoqbnAk9W2TgqZ0fr7Xf6
8cdueXTIEhDn0+CYz9DlDUTiiN7qnmViO/yC/yjYSSIiUF6zfszyGyQS9sUHS4AX
ab+wkuGk+HECldXndJGWFVM7gUq/7rM5j1gu+mydYhXY2995Ckv7gEQmiu4G6E9s
ZSMgzbSxecpUqEftlO6pqzH7WeUpo0rf79j6cFSm+dkzNbqjSj23pWB1uWKk+E1M
BfMPD3W4sGhAlhXBErWYBhz+GdvaY4BTAExlfCLypu9gaBBCffaFLZ9PyTBVOw/M
WZcU1zN2a5RpwlJX62lwVfewb8crRgxg5LS5TEjOaMnPrY8870cwqEzCRcTHoXKE
SxTst6yvClQyvD/WE5Fwus2sa8DXB8nVkizEu0yg4fPDfixz7Gwggmjjse3vxGWC
2qV2ADQuDtBC4uGHVPv18gIK5Ndu7SxJUOkdpD9fTci+LX7/SOb4Lsn0LcTfcsG+
/jJ+a0qX+rrhiFROD2Cj4JWkNv7qAho7+DUu33Bld8/P2YBJNo9SUpKFKGXKoxCE
y7xMCMx+hUX02U/I18GCTBps8sJ1eSiteijL7lwWptL+fZ7r8D7hPsmAF891w9Vd
I0rKeD3MNflT1CY4doF8DPayO2pKlcLB9KSoeKzdyOkNObtPKuU2B6kMCEnlmrYs
et9Wv6CcxnL3UixNL9yJHUuHSFgDDK2npQqPMVEAp+KKQiNKM6Q6a4spOecgsFsf
Nccu/p8wl2AQ2df5QxCzPwHYoVNL9xS7VbMZyRi8qFQmBApy7SAsAL6FQZxRQxHp
7nRribGreHI9EbInacgRtWt0LwZlg13Ya33xcPoRwsS4ng5wLTAz4e5UV1zBo6/F
SiWLhzdd//1T2wcNnZjaS/CN2AOZ1D5UU6m4bzHxbCCCqgudQMCn2DoAxTuNaxNo
9yW5VTls9po6gscBft7sBZB6eix1iFsnwGBaD/HYR1CKJMJSmu2XXtDexQdA4xag
3VhYM2lkwBWA5LOXDDtAwWB63CPP3KO8KSGIZp6vA6WVdCT2bDpvKGjqprGLogBB
eWO1FxNcgsHKFdDBfj+6bzrwi1m4Js9qzMlQSgJYANU8IAniH2qf3ecrmgy+HrlD
z4dct3ZVXU7iBmw5irIMMWLbH+qKkoFYz17tpCFu0q7EOt1ZaW5QoHdUUJAAMAcQ
C8B953k7GCyR1D1DZ6kehgBxTY3H2jrMIM0U//QzEeZ+2CaYuTh0uZIIlBEzZBCn
SfMjY5nEmnYH+/bVhec3joAFrWBvESFosQep14SV1J4oB4Fmj+Qx9gwPlSVgJ8Jt
WsO6JqP21SKB9dFrag0uqz193hBot0YVqG2YvP/yqTwQkotg/Cng6JoZOOi4ay1Y
vN86x1MgvaMI69sggZsv09peTeooohOzNcwjP8Vo3JhoDbi+em5lQig5ReJEup8F
GcelEcyqZdmbDCijXfYwFwAAvVqq38+XlkF/Y0G+cKXXv+NdpN3WES5gEDV6RsD1
CU4SdAnt52uRI0IEqEmmpLza+n0Ak5sVqm+GQC8Za+oNYSeDXHCgmARKChQb+3MS
sJiNrDFxqR1UFBGkT8sJbr0g4+MsV15tg5WzCM9FQHw6JOL6ZvppTvGeA5fiUmJ9
vRHNhyJqrEs5OoCtFoY2pz+wAh3lZosOLITY1AS4VWc4UkAhyxdx+fjXJogxEHsv
a7bIB1kTbXZ8ZuPc+ZUQ5utiGB65c4uGzvJyauHKDvHaLxThK5b9eSQSd6lcAk7u
+sqbXV2FKjNU5MozMoTHDbiDXUJig1MsWy/0RasI/bQzGOeowvcuf27EZT92OOTP
kQECGz5HMJJeC9OSuVk3hYwAuSf5q9kKgQMHEVUYNqG0TtGbPVQe1xXNRqpx7ddf
Da52R5bGP27OBzg/VzAwcG63W4BPDuTD0gFLH0lAxcst6sPEwjOtfZLYrPJ51bN9
XSXLlV7vbfKe2Rgsf6rJjl8HBOdaAN9U4uNxyN4pjD7vfUiIbqUllcTgkmz1l+wY
zB7NT0BH7G/iET/+DGilt8xWt6pytSXJXp8d8B92Iro1h4J/TaDvgpHyPYbOHrIg
PkGJmgn8NNUzpVbTnEGF5d2+WgqGu9Xijp5Wp9Y/Ld+Kax5L2GjVhpCupDILJORG
zGq9Iuy1eLQaQRawih5/YIWt9ytKVyS/Rg/y2sDyCOsesKKpZEIuo6v78N8Lh6AW
+CTII8CWo3/nM3WHufOmZxm9qakP+DWn8f2caca39IOEtirVt7nAxwAglIWK+iZE
788a+wuC8K/4YHjAQpxry5VIXPFnP5EqWEeXst6tL2aWydpPlpW0Lzk2BdYl6Yd0
MgP2fMDpc/H7wWsnf13zAaTUC7QF+ow0FKCsUQZ0MpmwadQi3a95GRL3Fn4ovbjT
Y56TKirOf+pNVdgyw36JC6ooq36euLIEIDNRLs9fP2I=
`protect END_PROTECTED
