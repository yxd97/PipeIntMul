`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/p5AZIIbDDXQq9W9dihR6E1lZfDZfsIkwzbM6x3zdkbw/BzX9i/VryldX/wj0+QK
ti2fcGXkaLVQVVTcIRFh3xmyrVlvLJpk0SjZiML4M/UeKdFDUUbQk37FaZwGrRqF
MdePxyTqoaLHkkoLV4YUFWcUfYhVulrUFCAIsk5O6EudPtlQce2CDq5KJEu2Ph2I
BKjIkwIMEDb2CPpLqV52PlmwPJ9b9rLgKifDjOeqmeLrbmmX0/+G3Cct90QQABzt
CpgD7ZFQGQEJ5t0df9KyHLC1wT4J5QFnZqYl2UNKjPlSJldeR4GR7H9T196ZZ0Xy
y2ETPFuyWyiO1hxCoV/GR28dPJd4WMjxhk2bsRC2O0fQLClr2juvJHaaF/iOCkDb
PoF0FKyiDAI1HhiO9RMrES017ydWCA3LUPqLcfSxVrmOGC8MbLQzdVg8rbYl5FwX
/BgwudfVBZUQesFLrXY8XOFUZqVrTqEMtS965D1dSXd356BG/z5321PL6pfMzelE
mFvy5pdR1UQME/fdXCtGZCTxw/GMpD1qwDeY+Pg1+0ErrF+dCTIzGJdPx+VdMQuu
ZXVa9TBaW88rgTn9LpIacqd/1Yy/NZ4B77OWVsAgjAmt3okbK/dVt7ybKghgNvAI
J09G/MASkckDx41i8DSHnmo7je6Y6IeY5xvA/7V5PZezO/v4YifSH50NLwbjX80T
Zcr4zdkCI4eX0doqEjv+pzMb54R5lmqyTcgyzd5QI6/vHPGG+m/u8P6x50gSPDN8
O1Z6PYOMLYIyAocE1IK4jSJx7LwCFL8ez0Gd5zILkpfiWcOyrUVYSoAnRT7yB1/e
Q6JXrTgBC0NcNuDerrJ0hSrBq22Oo5/d1stmkTgUQYy8rDwhZchZwWkP2Ovzjsq6
QEbCbuRBZ3CVKaC/ofV6SJhqpALQOqidLIePcghHRPHba0Zt8cIIEXYNrosj2hfA
`protect END_PROTECTED
