`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdoCAaH5FUt2x1zpRsqi6Mm1091tPP7qFY0isswgVJQKrQOX0N0yzWg43d0ONm+s
eNcOVG2EbWK5xLr/5IWaVjp6X42vQNe1/z8Wbp21o3rs9dazWKt98ffZ0xhhEddo
BSSBN57FD2GKn+8SNaOgHF+hTryCCFnufzUZwBj+5k81TcQmthq8WE8/SpVWP10/
RDEtiK8Rm7NJOO6y3frY9NpOK0pjCbW+xVJoEL5gqpyl/YI113L6bc/XF9ZjoEKV
fQgUKd+wPT+ZgT67daH43QcWOu+BGAdyHn98iQkYDm4fxzhdiRf9kNqRYJo7/aCm
`protect END_PROTECTED
