`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cl40jBs7fPs8gwuln8XB/qCFI/CeagkfOqgJaWdRApTsJIOYWamTm22m+gKVhJr0
qK5omiGdw/FOuYIkMMF13HzkFY+bzl1iX4FnSONVUwUuTisVxWxBAHs5X0ixtNF5
Rs/JKiddG6oYFtoFksVaqe6tY23AZYSzic4IgrEDTzOePyvDcAMhKR3OdHmacJt4
ulCY6u+NUeqmaEV5G6sTngQTtyoxl2eNeWF9ygswI7MvD1wdyosGu5jPV+kMJM2c
oVTW06hdorl41JK3wyY/anBsfz8ggZf3peVKCxcPYCNwj78HVbiLr3CVw2twV575
JKjiFfXh0zJkFjTpVM6UD62vJteZ5CfX+eMdDrhm6tYH82AYEZGiuqxSyNdiq+RL
qAUB9ATIN+kNM2kgA4w3z7JCb3ycoaZSbXjp7MFVVVBhSIYYv/peEzNC9bMG09Fu
WW8qYEYgCQiaBYy8MzihGT2O15ZIgdRqDa23Cuedl2P0uO8qQu94YvbQJQWniQbq
X6GkW+r0/VZwBb9PBBuPk4xwDigajPsmFXcobaNqmXKQzYo9Kzpa7h1PMbpBREIr
ROk3TH3QKOpFSMQhFwq/k4uqBJNTHNYHKbkdsbA/QczE1DLA8JW7nlQTQhFnczrS
KNDjSuOXSt6lWc8urB++Uwos57fBPxAYqr/l+ZZsPxpfR3TEKXYcKJ6/abwkc8N+
thWe24E3Uq5WANHTX/AhG/Wv48CpGcHhrQ7xi4odI/eeDtZHyCllKWOtGGJYewPx
ySexV2pYWnbJe5sA3XF0v8/1IvTTeVPx86+f2NI5Bu3xf0S/RYvzp9z4BHrHDwqE
OUSTdanfWMAEkFMbQaNP+alBdYHCEsKRMu5uiQWGkLneLg2mk/vtewb2Zq/+RmgX
fHrNvguGMiOL+4+BxniOJepma3yaB8mEQQjriO/uxje74jbk6I6BN/xXAyaXmlnC
krNHGPpQGm7/+p63Yjllb4CQFy8ShgSyOcPOOXI2TvK2OuUD5jUm2mvAlHadsWCx
U+ae9Ftg8RZrAUDx4pYeAz+77txgYx1OLdWx1sopA5BSPTVBzVvDcNm3u+ZTzNlZ
qZsHlBo8vhQCcrrXjbZFs2z5B/J1jN8VSbvPISjGyrScUFjkXsbZ8HS97qAiCMfT
KABdyqmsSRmnrKlhYQp17yDZXz6gCT11rcT3s07Ln9+hV5Nx6LwW5s+r0M6R9Wuo
jE94TaZH5LEHQEmYsOev7791cznO+A4Sh9PXsBzbYUFaBojp46gB/ddx4eKXmc03
cl1XCIt2FFDcAsgnPiRaRHnv/chHH9fWD5l6CvpTTm+J1GYeMBHRdvXhM2UlqAvh
vTCRhwvE53uAyQVPrgQtyyrBsK0NGpVAMomj/JXYKQYQsfqOqv9u0/5avZ+fYd2J
kFZib3Eguhtb6ol6GYDxozdSljP5XMtyBWyMao81F78uVNbAcR6elGEjvW7Jgxrx
6jtquE93LIpM3qDlA2R3LK8n6pESiHXZZBooyTQBLuCmh+NbdYYvoNz5m6i4OQqi
yvjtkpsSTsPIdJCzaguY0XwwVodZiUXgI1VvwcfswIakcNwbM4IjsngxipXdjlYw
tRhspzB70v1NmSYaLiSJkfwU6pNf+lPtXAztORGgEPGrdGVe3RmuNEu9eI9FbWHY
SXGTKOBuJFnAu8vQt0NyEVKM/ozerS6N00SQfGLZibQWxNgcmurlJTZlm8yzv4DK
xHXM6xcUvc7rblhl3wKiR5/ivYK9ppPSLZ7Y7WEZO8pvbfn5to6m3N+Z+GC8wI/U
BpO2m5ZT5xKDvEtrReR5Bc9WZsvSydRbwBlwJ5l2zPrsyWAxSWcga6oitLSsf7d3
q5UHuNMml4ARxM8lLE2wpxH4CNz3DACkue5U9aizTuwt2aBL4FR5u3N/2E/nyhd2
GKxFSvMxKqdc0SP7fodEoOxCUCxjBIx47PP1ZLA9gh/WivU7qFexizqSrfe67R27
Ndw0W5MV86aQesyYGEep9holU9TBWBqtqQV9s5/T+4VamHxFtrq/KFEJNsBuUJdF
tkkypbmbMFzpTRmllglWI+B9YEn9uVG6vvKOXwRbhp5WL1hFDx9lS5JlCJSsG1RP
OpIPLpG+df6dNCAu8x/VNp7WsgQprhoVRvw1mTFUPa5sMt2o8r8mZTZu/Z8XYFoI
juanGCHS0eG5LFcKdEl8qP9CtJ1sdiHokfn3Ogxel0Nqxbz2hEbBI5My9XsCn83B
IyiBpDVGgbf95kaOL0uUqftSWYBFkPVXYmBB0ShgVz52rfv4SZOkXbV+Jc5KVB+F
XtIVTGETLS/1TBgxJhXtawQjnu6w/93S0v+3Rr2w2gDOdryNjLuF2LBVX5qae8be
l56A8qBn56oG8gqGxU6qiu2m1DySzH8SfAw8qO/OTwVtJKqpnyglxUTbhlrm6PCF
nn8dcaWKlQWplQOy1kg7LINwNHsg76S1mv4ayXyQ/i2RgOUoFh34onEFw1ZeRLjv
gAnrC4WMEfFABUIEf1CSrFUeq1VAQolks24imNK2ypfKki3tTl+8ON2LbbKgvH9e
qXrVIpj1sp+S7EZyqmxKFcUHpFK0qubUpU+rFRryUgpqHM+3UzysUguuJ+Y9yVeO
R8ekpI/CFQL0S4BBx/g2D4p4boXrqS7kr3e9WIrnrY7l3KYq/hsyh8XYK1fsk/74
5fSiOz39eWZj/GdB4r4OVoTH3J/yFVHwMqut6aCTHyQFVvkpOR+Bq3HsB7xW6cgb
Zx4AiwVVMQimio28mxmRdqLB+k5YuN04wN7qke7abpMKgJXiT5R8LdUcPxDlODiB
psS2p5D+qA9IdXD5RmccYLLCQczq+XLYsKfwms69n6y+plEUisFhiBgO0MhP2GWY
BEcyISQuLKeSe5ikZd1NCc+SNk+1wELHoFlNkIluNiqf0NxdiX34QYSu9BG4qolk
KXA8Th5uEUxTVvkmBCQlUn6cFdkmJ406xz7ZGPr7q5X7mgsUaG7MeJviJ+HNzas0
JS+8HdTog0TVOG918vD3ysUUNnmvIygsxY8cwKcDo63+/cNtJnXadGKXaTlbLhGn
x8bw+8viTY8/hRCvuqPB+4NZcm2WUFpwDtvndiZUHdDXZ3679QL+hmdpLWu3sGqY
dFbXcBA5KO6+aHGLzpev8LAt3x6/z2QXdnUMTgLKeZa1BRnpZKHlTCIMvqw/oMqV
ENm9yE5M4ISdaVa2l9xCt/eFwNoZi4eqgMS3Saf33mmLev+QxtJIuJSpMKLcdQFy
`protect END_PROTECTED
