`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0j+qyDD2OL6m02QxRTKAXkM3d6U749wyE2NpY7fM8u5JcLatvkBhtB4X8QbjouQC
k1RO9S+PFaQBwwBM+8VQ0H/HRNkbFPOQl6kxYAXvqniyswV9IZKFPQeUwJ6/rePi
Vh7jZyn2RqGJ2qbaUmyzmTc5rcU3WlZ7oyB5tKAT+xQffJO9hLwxzzpw8W8F2fAh
Ofsm2zCD6tYIJm8bRWryHWZEOhWr4EkY2LaWzjyN87SwbHumdeQVgNKoDx+q32mZ
eablDjwjjwjsTWhah9CNgDoffiz3JQKQYiLjsIM3gf24UaLOMHRxRribgL6PqBzK
rXlPQCT6utgjHJfwHrBMGrnsAU2M5TAzm/enZIc/nqormZm5Nqm16fM+2Bxqbgrb
`protect END_PROTECTED
