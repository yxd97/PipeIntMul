`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wS5iWvdPqIkXtApDoixj787RdAUKxgGFS+O05BhkkGrhPBrcOiH4Pn8A5vMNTTJ6
UgzCdq67vPp/mLPBo+ROLnC+2YZ9xZzF1EBNYOl3YAtn9FmFO5plGdvZSYo2pes8
y0VgVfRhfhEebF4OlngCJhY5xqKcgCX4MZUD7TAriJnj6JrrSrWmY84FGVcipTqI
VTgSN0Edb+voQOlf5umdd4vEVlwdIb1eM2waP44INzAx+U+9F0kCVKyjlY6eKxYi
99EV7HOAALHOj/YTllynKYIu7OBJfCJw34F4squEHWAldqPY9Ck4Qe1mn5QX3IsO
3j1rDQt7Bw6qBB7CfzsbkMwnyQYvJyxc7Da7A1XFYtKT64axjFK12Fi+2UsS64z/
vmiEB5i2Q5lE2QDxn8ZH2djZeeOmDKXM0HkUQxjNPlDIhgMMoMEfDmr2Sl6PuPOZ
`protect END_PROTECTED
