`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sf2X4juJe9SqrOfAwiuTE+fzswF7VbEVAyMnpQkyFbwMAd8nxV9pN+xVpkjSIZCp
sWEJaUcotyZhboV1si7wsR74a3G2BiPDbaVr8xh5AyzwZFDbZoZ6mLG42GpUxKnF
E0LBqX94AQqdo28AEAE82p3V5vyaUMUxwUaScYuw85lsFK5wB2CJHmisaGLys+vn
kM/iVJEjXuw52zwel0vvfMUZ44qYpj9pA/EacXpOZiRRBUcpY+dJKh8WhaJ0X4Ap
651iOc76JEB0pu3wqsQhpNlR3wjAavaFAVgQ2g2b7UzcfKvXr6gYISER+7SqNEfh
PlRQGmNSlp0MfOKb3UOjhvJclsJala6ZvSSSkhQcFIrJe9PPBXmO2WzPZLCFBAGM
otQQzjhh4GXUphCXc18ophizNb6yVG0396VJYuBk4Z79hdv0x0j3s3XPyhHyfWNR
kyLg2OKxIaqrGfdBhz4+8Wu0aetapVDE1Ah5bPUfpqcej6WUGLDIrrgfSlU4sAxW
1QCAf859fd6CCiWxntc6v5po+Lr2M9fpIcPdBsfKclY+EIUsIWMJfdpp9m249EcM
RmodldUPBN8ioYAjno1bF91jL+czCvSAy7OkzjB5EYLolQH1tSLApnaHPR+MjBII
aBY+J3rmqUiAZGuzrJ9U2r/jDDuxaO76t3jJxfza0Kn5Pj0iy3pKWr4Zvo41bxNB
ZeSHR/IUbj3+jt/jTuqUKGeRxc5QM6Sw/aSohOlttUxVaWFy9TyxRgQcmVa83rj7
`protect END_PROTECTED
