`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VpStArmTDWdM5zbJkPH+62dB+7vow8sF8haPx5cGdvthVVrrsmwd7kW0Q3XeHce/
WfZa9vlJZRTbPA/quBCoHt80ijuo3OdJ59O3byR6UIsTloo1bvqCVyRjbepT9lly
tTOtSEnbkycyc4+5GIM2RPoTXqavwWkgeMOD+sAOHXHQ2WXeubAzehJXjm7ohNs2
OvSXtLcRGL/Qpe/qra83eDbqwcAvoa2UBhB2vTpayMNGbve3s+XTPVUfvhMGhly1
34o92FxZo+0kMCHjgxsYUhTpDqazW67rLgNy3dZyPGLq8F7zrnYHsAjq8chgU5rE
zvNP2L8gJDV8YDODO3R2xjne6sIWQomJSgjzrNQ01dcWSS4EpBPdBUF73G/KDIl6
eFwLsLo8IvUgXg0CNDP+r9POFsTHCedq9WZsy5uBQe5BfoPXSMBeVL2PdN2yc4WL
`protect END_PROTECTED
