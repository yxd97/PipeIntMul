`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5mLvOpFeUJ3634Vnz7cMSl3tX99hieIjBZJ68Oj9n9ESjhFnLULI5xAVNPcrDpdz
oqx19a2YPyH45Nm0q8Ejyf5O2YwcNAdJjyUSnTvaP1B/QejNJ8cKIEv4ZDgNryB1
J8NyUnn1crr2gWopAc0Az+LSGSrcJPOcTvry1GUBpnGIDL/xvK4/FTZlhHVDrKrc
9k7lNo5kXryu6VBzFsAevlITxrKHOaQGZticnzssdvOp84LfmiWOjvnuAfg0D6yK
blK+3BXaA4yFXqnD0vk+pA==
`protect END_PROTECTED
