`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
awN7/MdMbyQYcgMmm71PNza8Blf4vl8dUOPFkDyX2x7y2JAh8lUGeewnSmp7/IyX
WiEjlbZOBHOKFAgLI2yBmRIO+BQqDakb9yp74R0oHlogijKGGMTV7chKw7paAxI2
MQo5jVEzru9noNumfHDza1w1u5lynPPsKC7uDZNXGSFfJTYDtn3ujNdL1x4QbMIF
J6qzo4y6NL9Hd/BMdyX7ZJut/PDWJ59HlNUCE/t+V5iEAfu1oxzK2XYtsuxyRwtc
R//dRs30lIVEGfm0iSPjhE2SDskaIEg1HrFrV9liXNJrGkOaAgOyPxM8cQavY1+Q
LMXkI67NiXwrxBwyW24Vzwr/cKJkBsyf4JivcoB5XChpIpJe0QKwYqtqKqj27xTH
kbQFJ9zwy1J5NWRxnj0iiw==
`protect END_PROTECTED
