`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kOd6H1garqcr0LhPF5NC12S5y0D4oOvUQTUTd40F72pmkJ2yZRhKkLpPH3rDoQvL
RMHqSN0DomidIUMpUR4fGsL8t/CdJ0VL1md85qljfkiAQsbgZJxK/0KMJWionUGA
B9TR8XurZmfEVh23ZS6S0LwJdaurx4S8SvxTwiv9lRGOv8ZEoVKmV1sjcEonsjz1
6LLa+NmaELqLCqJG0WQ/nz56zjSozD1j3JZvsNJuIRO+kaR5A9ZNrPRTCjp43rH6
C9AjSU8YMsE4j7tfWLnjgTdS+ujrtXQoIBxoAa3JvWjC5Q33DdlHoVgBhk9fvR5n
OGPaeFhsQAUBg11w7EKi2CQYBUlsnziYX/UeKac3Kl6PmvPl8l6feqlbh+f77EpD
NMmOX2166pMb1JKAtpPtRg==
`protect END_PROTECTED
