`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4yGEEgVIY0msdoWKb8luZ3GXOFFSAILkpFN+EWsJS+PbC1SQiJMGpnb1qONzvSe
4+lozprPD9t/YrgXs18Lvrk7UGPokQ6XO3go1RqxxGdtiQigM8FNhVch/aUCheN9
5rUA9jwQ0y5E62PrCVab49+XGdRFmLgIYHv1N0f7OMscBl61skgpvuZgQdF0lgBk
mNj+ADwNv2EbSi27BrCVlAizMScF66Eh/BXP0E0co5jiwJhWI6siDTDmgQl99ixg
QjDzVomW4y0aBO2a/hZQOEYjHi3VEP65sBnlSfiHvN5agVK/5SYFTtH5+9Vl5YvS
enRx4yVNvTS3C3wYRfRQZkXB30wNcQZELgJE9xA5tGreTZdA+hV0IGWxRgNCKLEq
WbHzEYJAV/cPM7KW8iqibm7FLFpME6OuoHfOSLUxHz6rSZTNQmOtJKc5NkY+78oA
uIOLQDjt3WNQ7aXgo0PemOzKejX4LxlH+1ZMUX84fIb4WdjmHBz5QXaT/EeNspP0
4R2rnLViV4ZrzP4d89X61Hs2Nfd7rpNebT9bbQ7gFfJS3qUfLDLQWvXmdDTy1FZk
t4m4LpTSsyzDm4Nti1jjUbAw0tJnUzwNYU6lCKx+9YQQgQzqNupxOqnb922moX3L
CJi6CQ76NKWHkfIL4qi+JHL32tcamEP0gfXN+zXDjuR9slWXGxmVsGGqwOg/Hbub
OXqAn3jXCt5eDGtToG7Ene/RM3hynRKXrPrMJ2/qmulE3xYyHVHWD3ySLqXPIXO+
UuUQQYrSbv2fWahkRAi+mf88iR2VsuRYsBDWFCwhdS47sUNFsPqhOBYltJwQaO4U
SGc0poNqB2taHIk251RlsA==
`protect END_PROTECTED
