`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Au5AAxvm8g8vVanPXfIxt+LpATcOJ50nWlSjgZNUQGc3MoXteJRzNcGFMGWESJ+s
56xvYxkgVQC+EXsqhKwaWWwz6xeSXPZ79BGxIfQh9ctMg2XULDUQiKE58n88SV1P
+vTNQoXbRfKgfdhYXXju5I9M/RZg6jFJ+2We2wg+iSLdYAEdHqGVEkaBEoeVkwZ1
Gv/+bDnlpzLT3Hkql19rs9mNlq+IzeV42E2fIs6xdJvUE7DXNklVco9SZvLVa4A+
A/eyFrQXvwBMkkaeIC8xXE0fBnOFMuIm/TW2ZBj0HmrL0EoQE1hsO53BpmJ2heRr
WlxIM0mWj4HyfxZk8HHSKKvwf7Db1+4F5xed4kpg+O0PSrtPgOIA17m8U2xVe+v8
lQF6FwvkYa14PUYsSuigCJxKBvpOnLq8B9NLhUZ+oX4mY6R3OJo2eUR9jyciPObi
FLah/qgv1KZTupNp74CzXhxNYmQ7whbeY9qX7RIV/G+9rehq1fXyRwa/5sqB4fo6
sgnncNds2Ws8HkphA/GYJ8jn5rRWNFWPhMCYQkqAqsZRi6WBXkdv4B8UhMxBRiIw
n8E3dwssdT8DbV0JPfI/EWBd3eWsXlXKDLTs9Is5XOIyhgU+mxpYGPn3blfq8zE6
Dpnq3tf+G5dst+V9F5w3XFzNQ0yIFjlvO/64eihf0kRyr4tcoKqGtG3N2DVQLvVU
K9NUUr1cFq7PJpBVdR0lpOP80XtxwZph4dQRmtWG74PfndVBEraswppGFgn1Mm1d
Qq6P0hBmA+P6zJoV/nJRzZJzBkvGL7gi7QWEssKNDJLeD/ynS9fK/j1CMFFYDPLK
xeD/9MIpHGjYwTH+4DrkP+EJLigWyz53/rb0ueEXukjR7E2kBifDfKje7eyD+ETt
/mUoJMc08O8pgySAXIAZmVRP+PXG1IkIViRkKsc93VhbeZRqjY0aPS4+ZSkyyDJj
B+LYt/zwWSNXwPdAgoaajpvOjMQnUzNAUgnAyrQ/Z3kUnE0+cr/sKGQVRqVudBTs
ZoZPQhd10G4kwKzBqYe/+QgzzGEOa8jt1HVzOznNVcm8W4O9K20H0T2xvlk+8nCr
Ot8LQ1b2jf6zERBS+sys0uek9ccAhG5fn/1mgA6il5fr19zKEiloWKgc6a3iEsK+
85sXlio4DfMOiKY6zGhJf0UXGz0znSVIAmteG26dnC61jPAEkCIUCUuMtAb7ki0w
5vqAMs+KQnd64Aqne0rSXFEiNhPIUUqwbl2KB44t0SkuJ54zfs+HmyhiOfkDrBvW
WqpYX/p0AJMGrPl0RLSlRQFt+XY22RLYjlg89XWDlQV3MZ5foNuTbcfbYZHsiStV
`protect END_PROTECTED
