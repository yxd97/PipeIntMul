`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/3EcocqiakIWKOvBrEHrPBzV1B8/0ejsNzeTmAUm3tYOn/yfGS/aMMsqB6Todh+q
F5vjlMq0PTUP9/19lFZ6PGAYYJfKGfW+nzuB7ZQL7SZst6wVDbMyQZSQ5mFJx+cR
hMIf1a/kMJEesMNA/T3RM7q4B3ZxHK5OYLxsaLa5lPe5QECJprOpbOL0UMcQo7U4
uqu8TCU42Dg2YAJtprgyLc0CzPubxo/Nt9zVsPdcfeU=
`protect END_PROTECTED
