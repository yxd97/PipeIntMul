`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqJHzIIOMxokKCHDN0/aEzY5KOQFFUsdwB7p2yH/+/9ry74H9uVr8gCkVE1OFGE4
WoPR9o2G3ADk55NuRQm1Xq5XaV8xQMJadOEvMg+N7ZrPSrBWJwppzAvwB4wUJKy2
P4x6l5bSbgBkENE6rCe64BkbrRU8j2rgT9aA1Mmoo1Izcr6KmcUBQlxh+aUmyuo/
QMXYC5sx/cmhYidcFD7ukVHwD6FfJ3n/heYdXVtaJ6pSezD4guJ+3xAzWVOTkIHc
zR39EevXcP95fzxX6KsutL8vZRADWatCXhIHORlWgzWTb4pcfJipjg4tZINuJT5c
qPKURmRgQvyGZfG6snN0Glc1WzU+OM9AOIpa1be33rB2JTCa5Vfo/IzafmkNK/zQ
QVSKbDqfuVJpxoORuEbznoij+pfO9R81iBZ9mkcpSl4eqDaWFsy/2yHz5oVCsSpa
lmd/MViv3p0g+KkIS3NEDekuWcJfuE8YR59m7FW3foM8s1fubrjZDku5jHx3E57K
`protect END_PROTECTED
