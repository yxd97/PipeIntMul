`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1YtLldIFvesVJPAJ+CAukO5dyN3gvsUN7Gh3bkWWZYmVJdWWMAdXxPBjZjC88hn
/dBBdNUFJpQBB6aEY05WPBfClVTul2dRWPy0yWpRfB2vqgyGP2LspoOFaSCPOBFG
6nrX85mgJAbEC7QD1m/BKdnT/AxGGeYYo8Zz+e/Ue6BxRAeuPj51THeoIbtjWNaH
UpODx9gYcagINGsHvihMVygTTbVgWcdPb799TJj/D/xgFjU62kH7W/7RqGBn+C7M
LbAbd3rLeyu5ZXDuHrIRaYFbF5b4PDnq/ySbzuLzYvW6c6TH+xp7FPHZtakw1JDQ
IprjvVTXsjxVIn6Wz4QnQX7WX0sKvIGiy6XR8zO7rAuFNZ69P8v272mUssfCL2Ii
Qf65nUtXjTIZ1H48rWGLJ+U0yKjiHTs0UJU09nTB57U36cwPcDVpjH7YfeQ6CQz0
oJzLFea2gGheOP1kacrOaI61VFR/mUnWKT2RPFd1yePjE83iXMV6VgaH/xq4Dxla
KNIPjtKCZ0Eo1n+tmAe98ItVivNCA/EOZtQfJoQj5sCBt1pQBHl/s+CCHCUH91Yl
vcwWxAXWmaLDqO5lR1mHvih1u77lf1Gu1FoVjEtt75o=
`protect END_PROTECTED
