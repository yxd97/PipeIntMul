`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCKrQfNdDAMADdTfDpWYRHgN/S0BFnJdmSPVf1El/Cb3ou1MhoPR4tVXjQYH43AR
uxGMkfSflwwYAhU/eF8oCmZcYZEPODd1uiffIo2916YMKeTMAWXYWpQqIGjp9wiz
mIfkCjH23i1BtKdtCs5DuV1yB7QeH1RLGA5sGeYj4Rq77RjR6pAFL6R8grssGVUl
zPCdj2xcqtecyfE4s8X32bPk0GD2XWAacDtG0L/N9EwDo2u5qPxUz2MogvuAQ7XD
GeNC6RGR8APHvi0Hrz7tancaEmzu0lpc2sWUggAPGOPqmiFJiCCaWwcXNHP7sE0G
r15XGcRPR5AiqarSfwhtypa/9pp2kBuw6hc4liZBTRBM3NmHevAEeIirgfSo96R/
2rHAFr541Qgc81n6Z9RU3QZ0RX8NRdqVbmQKv3ndgDlMO+uo7GMzJn9u/xjI7UC1
VwSFWMVkYUzVeKE//CXGs9vRJd0yJmb2DWimlTSejynDnEuEQCHdchVXpvgMrkqU
/bK9phdQ9vR07Quzi0MAEQGN0glApP3tw2foiP0NLYjrno0Z+9v9azc1eAHYdk1Q
p9vmsSROn7bRRZkURb8jY1rEL1WxqBCvJC88VGqPBrz9gqnQ5Ps4hTDrs5UirTuI
DjMAZLZnG2BxYdTCvEJpGfkAH0rOhUrgox+6qslAOSO3AfY+Z+VzfbgwrKHPcwHB
RCJGRIDIHS7tLU470olsfvSGTYSlbsrB5zHfUZVBJDHV4WC26T7N8jG8wdSSkDLT
bq3W6Q9CDaDW5DCbpCNmJMObEPPaeRxIPDECc+H+GeqxmKeDrFxvSSEp1aoZvzKm
vzUgjyp+KQ3NSqqrE/Vdn+njCoqxLAfRlisAlBB7aBtsM4Mw2TMoyq1MPhIQmjyj
b8aUCVLVIjQRzGAruTQq1sVJiTh5uZOhwxSDxr+3GALTn97MVO9h2PqTauZsQHPp
VSTfKd2lL4v//8TujEIa/v3AH58W9E4dst3ofLvy10/QqcJmPih+gWFgMlhm5b/w
DVZVrDmrIYoFUp9l4vo7OokCoM6M27e7jJtmkzrrC/dY6jraWthveXXPbowYBIws
jU3g6P8qLwyWwo0Ze2TXeI30DwTlIfh844syPgu9c7m3QRYhdlCkTjp3qsI3qttK
ZYjsHRbcB/gg85DojSSQfBjsenSF9ZXBXujVXhBf3RGgl6NlhUy/g8z+/d37Aqn5
Q4Yhq39gVJqZwBZdUWX2bFszt9f74btQWADELg9d7zUOb1TyNgioHaYXfGQyPNal
VDyMI7MQ6+QjpHA/Aswwzco1/gz2dGuL8VrAiAhhtDxgIdwmKbKkN13G7UUBluFV
4yX5D+AS1EXmILVejjqfCwpWEMDn6VMyj/2FL4CGg4EufH9a4qR+AstDEauwmaop
/EXHPaP9f7w2JMjvbgdRiNf00WnoDmNfEi5kfq86bgeugl9t3wY/gWzZSaJLbLGx
m5gUs69l8jUxiLdevBC5ZlLgB1CWd/J6FF3bmKydwvWq9y5BOP0X1TRnWlZP7AfP
2Qk8cLcO168aDdCjB/KnDV/j1DHYbLU1GA199eHWdI0bG/PSlHDsuy/DiarHj05D
teJsBT0D/ginlvcHlK4m7ZrHx+1eCvhmD/NMEr02PIKM6UrOaGevnkUE5cVjBvyS
VrUwJP/tteBR2MrYfYcBL+X8xyrCY58yYCnw7PO525ilK/BY3FPWNKb2zNlUptN3
sUVfdCITrKz3Cck0w/wubo8khpD0yoSk23oGYxR+J2bRu3pi4TktCzlfE7Jwfceg
iuyAGYsVgvozB9euAlbl7OL5kWOW6bFYT4MDfRtEjHLoKdIUsH/Y09ppPetOjJqZ
Ic9KV4rjAtTWDpNbJNhpp2IBJhR6Gq2w4uxr4HMollsX526QsppXcoAUCJT7x9WK
O6XIIa+UHsFhYq1wkffg12UNq9nCEMOv6bHY1V13Qv5sDLMQHXGtVrvft0vIE7kC
v929LIhy4hJ+RwyjRACvQ88kdu+s9x7BOe4S9nuuGQamWZQSxXLkud1nHl/oKnzF
mUQEdfNQUEXYGGOMBYh67MLJ4RyhwqABjJIupfvBPlBYsfoApykJmhGxQKwysX2c
GXfkFNjRZsrabGN7COXb/8/BKncYdJYNN6AH2p4jKMenyEeZ/wqd8JbnG6ccsOim
p+6PcwNXEm/WAlWG15pace2xLsMionDqx0eMKbg3RnQKZ/KT2POMOtCZxCflaH15
LHoQpSqypSQB4r5mfOFHdusSMyXmMOOJ9RlDy/6byk1unb4j0BH1f+nkspf5F7dW
pEau/x7mjsi5AfOnmn4QyQZZSuRx3DrckLgzOOjiVH2xsJ8t+BvLAPOwD0ZGygxf
FcAxk/6TaffvUb1FmBCva8cLnqkkjJ3fHAX2kRAhJmWSKCUvcie1wcVlF8GFPTPt
o7iAZR+054VbwUyg/lTTKrrubxnqMa6XzNmc46N+XI1Y2pFfHrqONLoa4ICIV0j8
cvLkc3iPTTiVo+k6T45ETvEm2KZGf8yuz7LQ4yyQqMl3NxOwwxdTWj0CjkM+48P7
vXrwP0X/xUJUIP5Be7n+NGuMxfXfJqAjFuvJ4nMsIbCsN2h0U9BbIMEVmtulqFuV
GSKhzLYSx5bUiQCjV5CnGibvzLxy097BleUSTUO6tAyA6EfTsXsdJIDYUNVw3/GG
SyXnjbrdexp+Ju7+Ok67I3YghYkQI6BH7w3W+zqbhtBkB5KfAXEpV10yCkrrf6aU
VxA9qN9esCo6W53HCY2vT7NiuXZmQaxAFMXHcMPTYyueHwzNCquOZk8JGN+3mWNF
FYgZhI5Mp0zdvsumbky4Jv0p47LH92tHcvVUhcQYx4OrTUQKeGsJGY7JWvtyqCz5
otFWmpqZ70aXHAgyDupRUgMzer4+npvOI0Ct+uLuC2PEcCgI92AH7ipUIzGNKLnK
4yDW95JT3wd+8y6a9w6RLvnW5V6bGz92fvnnG00RFzkq8ok149Tnf9v2m/tLKlTL
NcKRaB4RJH1COyl9BGw/djaPPXpbu3r2HxBtT6WbZQk/9K7TEqIpD49iM4uYyBLv
wO0bDXk7gsebXghKPAsqxls2lfs72PyyDpoJPImZz29IpcSI8xNEK9iZwWF4WAl+
zTsVxBNf7pe3Jta4z50dxNi07UIofwSe5wDHhMrUbGHZZ1QxJ8UsvxILRWrlKiEX
oZt1EscGm0dwwkE5D4aBcZ3Cm9YklHMG2IHlHM6uPYddpGnBu6SE3axtRxOoKef9
Es2L2je9diNen78iO3ijuf9rX3G8ntwKd6B3m5sMTUibK5GVDRZo17s68ZVDOm+Q
yqEDBr9w1kY8Cnc4bK/i4ngPqWZbnpSGweVhUQqsPdBW5pKcTqio/7DJifAcGfN7
BOsc54Oq1cEXYH03q3w1SH/bnasCC71Z7sC8czHmJZgGHct95n6Dku20fvXwHN2+
33kiZQlWpZ1oiOzbi+WYSfEqPtMp4W7pqqi483wdbNxQ8e4RgB9z/iD15moC7pw8
xwBMxA/xEUB+2DWHAxxY/njbGun7pzWPJWoI6bpegK0WF6xv69hMt3LEvWXZ/B5k
uHTRX7Y3gtrbMRQ5QlEwds/wrtN2MY8+UIK8MJNckd6dRA4W3wqkW7v+gffpEWjB
b3xxZyIONcfyT7BeeI2N+I3W59S4t57lC5oXHxwh0T8yBu01LifprwlMjRklrMve
KJneJRriwI/3rFoRavEjjMFXb9JAaGDYm1Pob+yMRSBoguossfd5gTguA4iGEtrD
31ABBjdnhJWMtEEsQ2udM7uI43aU0SHOgBrNxWjt815vApkTvqwlFcahTTezpGY7
EIzpzqCJcWZ1/GrsnTQvlvjEyal9+eSQ8LUBWfherJp0Y02eNEArHATNk28FLHPO
xl2SvqvUN0YaMSwVXpHkKI1KdpNVSoH3kd2jPXqeT5tNyoQu5/sqEx/N3k1sanE4
TcXx3smR+bCY+RwVnFPzS/zpmjURGmsmMhmf6yqdyINjIeZLxcDUdq2kj+lSmODp
f+FditHGGVrgUU2nmeJUkJxmDWyP3oX2lRpNYTXbgwMBgYIQERLqsKwYmAwyeQ03
eyv5vxA4JGNZY7Cj1zruoXLu+fJ45Vpo2ZAGROY6tl76kBUkoAbPOEq5cUuXPaMk
8OvB/49C7pFE3QEjhYE35XM0xQ2OPwwKUGRqhfSvX8WUgbihBaN+Vr+lWuKOHbqQ
sLq6er4IxADsjnjBD89ri1XjqTOTkrzK2lNMengEnFEdOAKQwXkw0T+DS5upcRH0
co9NfYP+8TpVoElRTMNnjqyal8Xrh/Dzqgf95kikSIpEkgpq9Zb3xaaB/CsQOuTE
hUTna0qgvBzcdudoSJe+ZltIppqichP/4ubORzJUeaZAGNY0Ao6td7Babi7Yz0Kh
P8VUJ7Znz8IB7Rfdz0kmIAXgQ2QfiVo5VhxLGaMec2Po6mV6stdrFwalKzhnIBDS
MtUCRK+WNpy/7ZHHXS6PzLnEm5H8OYtIkZze3mJK+P3iDLsFIJ2VGFfOd4Qrh56o
+vUT5kjRuTGHRjkDf2mo8e7X/93k6J+YoRVKMGTPYSi2L8bzm65D3fndswSym4Kw
JDrrJL8bAhHAxbeQ5VCa+CD4EaHrX79viNlIHoeanL5Tp0YTjeJE4OkQ5dZFAXFe
1fHWHWxROg6ND3HrmR6Ut/SeE81XrK2URSra9Y28IP7cYUwljXMSJCWeu+gALqPp
45RrTcOUMBLCiRkb5fAV2Yqj2aDRbWyRPjmS8Mg6AzAR42wYYPlJwei1/LLYfJTz
iVvW4A6eYjNr8f9rybrRs6ZykX36nLgoRMO1w8z5IlRHtSMI3D39E8FxEJLkU2lr
dZmz9FOr29juHiYhEZCoPPKPxFXuc9MWAa6cYDK7jHv/rqwMATo5sRFuVjq+bjzL
r0UnZU2oFaq/vSqTnI1saMRkSMxpdrtudW/xBwRr/ZQni2UBFbd1ybRcKW+rNYZQ
0zl/WO6TF16KSqmow3JozeBVrQnznDggIq44SZzJkGNNRNtnN4j8EJyhL8UIzBK9
iaYZOVF9Jj+f0KiqmrNjhhO4NG8QiXvaNfWLSnYEScZJ01LwQ2+0qeDqgcsvyRQm
eVkVQ+9BnhBuTDJfaePLpj8G/KfD1JWt/85ZHb00e2a0GuvWaXmocYe2ZEN9Chy6
WGYkaf9QrKtoYi4jqu83rlNhU86LC3wQJJnpAb0F4gplxwNIJMXIn61W1cbf+yUa
VoOz2oK8BNfXrexpQlf91Edrj3VnxBIX5maH4vcO0+ye7v6TJkyFqjO4oTZCErbg
GcLNE3NAblAtW9yuZoDyV9KFDjAhLjIwj7dKNT506CmoxjUR5kxNM0VGKf6nQ2Uh
4bYO/K+6DIDVZtrFGBdznwH8QY5Jb9dZPHa7t1PmmfuG1rR0uj0ble+QYIAfbsSh
1eth/iM6MIAog0xr6SDmOnkWENH8HxO4TOLY0FCDE5MRfuV48H+dfgx8L9gxfsn8
GO7sWraxdbV9Jy7vjv44ytayS8nx7RVOTDWZOhvb904acTYWYz8LKqVQq2WS+Tav
pqiNu0AMS+JCEY2caThJdIsFlW1VY9iPPB58AAC6+6EgTCnzJWtX2UjUGwmfEXyo
O4bJNgWUlrcZB8VHSAtBv3JWdCqnkMAvC9VSTiF9whB5uqSKf+KtNVm82oyAGVZ3
zIzviBzGUewVbdLNZeCO/9hrNsGetOrMt/pEd7UQDbbQZB8A2k8uZ6B44qysADp+
v7yAyMjnqI8uJ+rlQSnBohAyGrnqTqxDFs9DIoC2+b2tSqigpyrgIyJO30sgndWf
auwATlzF+4g63FBOVUrFplfrsM5u9mX7gtuQrXz/CA0lAtc8BDuoVNYyWcw40wjL
lDvqnBzbjWCNk5TLdOXHt0jyf+TLxgfY3oEbKZJ0eFtFrE4Kr/0ABte0Hb0W9WPM
6ALAUJkleva/6I28VWavfqhvRRPmbUAKwItm9Kmbd54AbL/ll7NmAp9hsSGBs2O6
idFgyy53dkNjUO4NkiCu/dR89FPEh7uh48VXJb1mFLkEGQQy+xlSfi82z2VwVaDq
NenOMWjnky3hi6N+/4gHEQcbdUklDMyejktXMmwBZ6AnU6/TbYd7yUdfRq7hrv+c
MoB58waKhezCHmqpifq3doDU9YwwuSQWYYYdzp6SlfjMHOQUw+QHZx8QQk3r0kSY
49PL8O3xb/C5E4OsYM/Rm/AI3MEd1OKeUTZuZUgMKT35acVKsDtNH5zvo67WomYA
Ss8dnKN5+auBut9BSA3fTMTBJtHMbgT6ykp5Umw8Mic1nXXo6zDApufcjHZTnw1b
Nwvj1PpBIILIeVwev7EjzLeR+Fa8r1jwFi7QiHA8xyYfiP4QU3e1rvKQCQoyEY7f
nCjU57wUpkDsPanGSQKozHsav4aebOnb32Mv4luEc0QKbZXGC9WJE3uv6OigVGpN
LIcEzAzKbqRobPbSQN06fAv+6ZYDRAhWV5DXy1Eb/psWIIkvwUsWchfI2I3eFaBz
nAhKcumtUAX5XBmpauQ7TxjTOTaKJaV7MqhMPmo3D1dh/5z03YtZzL7v5RWVQco3
T5GnazaryrzTVh3MdwZm1SAJPCTY6r44wSCWTPo3OqzzirIR6A4XuWbAlWSYut8j
YFC9TOPmm6Fy4/IHmHxdCE6nYXbIgU8GSmaMq4q0jWdtwnsCJ5QoHiQZOA36sDjd
KoBzL8BtklGZRYuPHOfshNFRsRNbiIb3d7Rp/Zo9mTluMdA1PzWN8W2em6ZQ+oDo
O0AjUc3XskhNDgKNbaBGpRA1t3CE4J4wMyToOHaKEBVEBV/Fh4puwhQVFA16DOK2
BbOIECQUZB9gqcQtG8QCE/ex0FzkB0KqnRBiKGJeaLPrndNTt8siPzLLn6vuqbrO
laPaPQ39o8D9zZq/gojM116//ycioSVRyBsC84v3KmE8MLoJM5hxTbM2jlu2rOeV
JQ3HFAXtNHvOYCaMbXXQ2jBV1eCQcYDILi+dIkXz00AWYUgRgR4oaFQj/UMZGcVs
AAr7QrLjHsKx3o7lEbqBc3LGG3Ul9n4UROoEpq9J0Txr1hYAXHnem8eIfzZrRk6h
/WG6JolD4HaZg5q6wU959MuEKSwzuc/FXH+ZVnNyLCrgl+1XBxqM0Ej9tP2IN3eb
IhzYzSQ71uLW+UouUSrMz/Rv8R0LvvtHeOGj4D8hCeIi0nnhxN1gU0lDYtjkvx0F
KUmMyL7wU1IHld/f5mw2Wqiv3wb3/vFSDVPP2XIs6pcnDiU1OKyd0NiAZO5aGmnB
frm6m8NUDXUZ7N8c/UC/yKiCpWRIyeX5yzYPxP4OgiFD40KcOXBmbPZKVAPpmSmK
v6ywa9vRJWVerxtcvoNHbCuRf1ADR/48UxHIkrITk3vDA3JgLOPhgwupch1MA2RK
Tq6NVdGrePZzeIgZ2U4sakg/Nop5x8O51/NKV2xPYqQZqNrFV99uxZijng0FBIKz
FxW1cLuqrHteesr8mSY51Ei6AFmjPGosSRtAbfDHm/lF7AFFuy/y0hfzsoRbnYKz
BHH81uaac8AsMQYBZX5nTeTDlfk9MdjkbYnvLxz2E8qOPdjl09AWVFm/Lubgw4iz
dVtnMX011vvvfk2WC2XnWMgYlyiBDhwFCtZVNZLsogj8u6QryteZx/VY85Z7wbn+
prRbvbui8TFE7oViQ/P601oGZU5kyedfL3lvxiFZyDd/NPVPbGdefEVpPYFPFiIy
K8TrxQYtbUkHLHqRlnEvnpZrK4S07Xp9R9Xvu5MOzrTp1heLqmNZfqKhrFAZY9O8
vKTdXv3N/SoID5TZdGYWroin+N3iAKYwL3udTMUK1HUj5aHWEWSP3pLDSHaOk/f8
TquT3nbYyNHLg1q+OkVaf8/Zv/Bl50kIWScLjnHJx4LuAl/9v3z3RhT94LAV0JLo
th4Y0hxWJvRJ4DCoxMe6akBm1NkRmqNnApRuIDMOhUipue38w8yc4xTl8I1qK2OE
CmPl0x3AD7oYtlxVs2Me1Gw/9IWocc+gqQVZP7R6ZMSerSY4NLF0hnNjEHEVhhwi
wCUMck5JGcb/9PdaTFCtc5Fu3vuYlovu9epY38tfg4unA0ay7wXP2gdnFe34f5aR
DBDTgBw8ruK3adimDig1jJAcxaGeyVxZ/amaX+uLpTjExs0BZLyV3hAB34+Fjf33
Ts1BBnEKojAZZsyLs34o7beawUiPKo4FsiPY+J7Av2BawVWppvVUofpvxVtIvYZP
9XqWK1cH72nKRh4PYc3uPdEvEEt4Zobjf9aoH97isFNsIJ7q1JX1AJPsZgOqo12o
ZAIetywcml302u85HUX1xTbmIYh8kX3vuleRcQUkhB+D2fsg9GDtBIRpGV91AIUG
xENTvqEBpakHxrLdt5UJeDWm4bj6ZlQ7ODPW7Q+Ux583p25WUVApkZVy92Ih1yo3
No8Azv/UKFKBq6eYxlfiaZ1K/Q4oHlcthd9IbcIGO61K6CcJx3JlPX7fGx0+GvKQ
9+tAONOQGxi7u2/aqJMRatYbfvbk8kmbygHH0R9UnelnzYLmlK8MOtn1D+0Pc11M
R/SaWCROuc950IYQdHcpMX7TpLqpj2DmrVSMLn5XTrqsNBSXjbCN/TGYw0BjGoAU
MFphGpp31Sd7tEtRWYku2nVbsWUdLScOBkPA4ewVH5CvXy5mCooyBQz4XRR+MWK8
QYG6W0NR3wuKrsRv18C2KC9wjCXSFdWf/+k1NoCmGlytk9fods6FPsnqeQjfbsUZ
zU7X5qw+Si5hcq0qr3Nd1c/EDEFcoThFYXST1fG4mw88vh6T1UM+BsFCVFnh1MVp
ASICyCiolUAH5A5cSeSP9Y7neZNcB+WbahuVYYjtksBLO8FUZnTwqf681PO/XH2V
EFzxAuT6ZCf2+WEtKJB+3+TphFUTzsOIBxVaVYQQiz175sQbG5Iy8oQ+/mvj5cuc
FrmAsUa+I5XlAyRg7mE5vXdh6XijhkUEQTxiWovUrwtepqh3ocPaybFN4jfLqivK
MwXb5qney/QwdfTSlKClFcxkDgBxHNPMprmkm/1DSJBNy6+jRInn4LQj90bG3zGl
RuHliThVm6tl5c06X2/PddgZYKdNpPRMah0X4bDAfOOlDuVyiTlSPkQKdeNPnGte
ZG6078HJTy/oLQe1bmcTr7XXlKwqkvfDUbEo2dZdCjAJ6EOgO67wvaRwA1PmWJ+Q
N6zBIiLlxOvH/1AN1HeatbEHR12pz7PapilWV0Bf9Iat503vLF4HOn+dLOzM0vO/
RdMgVuZm4cEh0lwOL/11HjQ6ZCHGrxRaTfE/8KUci7QbdKVWgvtHcRdL067paGIQ
r5uzKv8X358a/xgi/bpoFkQIItH6sCBDUfMF8o3G4JMRxYGDcrZItd2tFSqQzvMM
NozxSiNcpYsMSiJdnsXPrwFvUQjedYGy1/AeixUOrP2L32oK7tbcdYOwSWuzVFDK
+oJMC+R/knVb6r48Q+CIxHaNcYMzsmGOot/3iGzpzX8Io16jmVBo/yGtoN7u1cm3
ZHZC17YaWNGDL1wWi1lxeRpuWn+FtyRCuhWNR2mNvOqh+GYpTPwKRcc+utK9oDUD
J3AwthRqWwdGhmfnKV6dQ9Yx1y9BMnBSvfY/0jVlrlKIFKGYKaVV5Yi6K0cjq04I
StYDkyL4KbZy5g9U6g56a7m5hrxuAEscBvdGQOvhKC/mb64CipTzDWYqPlfjwmuu
ebwT4CH1B+J/8hrZ92lm7klydEhH7boS0NpnkDgzInJa5nrs6H5x0JgqAsqoSyVW
hdKRIwCEW7oVkOQOjMUC3F6ckdGcu9dod4VVXwFlonUDyMvAgsaw8gp18vWXoE0w
10yupQv1k28hQrPD8q9QdFuVti0auAdzbz+88Q0Vyc7dTJ0nyi4Bcuw+J5KA3Q85
dLhvi83f9h4wfxO9ZqA1bNNdPpIpzHROzXn9B13YyxVqXN8cvcawow6zBbVb06UF
iPtwwlbp8WWtHqn/fOF2OAL9lua89RSlqxEMOoe3dT5IA9bP5sbuY39+qjuH376p
hvZqqmGcIMSu4fl+6dPyFQfO7pH8f54MPA4m6+CmiLa33A+efc+xq8q860UD0oRq
JYKYJX3xRvVcLRw5+d9EClQkWFx8lwXYwW/R4mMdQpzR7A8GOelBks0MclecoN0l
TMxPzSYCEoIQUZs7Ho5Mlxoeo6dEpnIXuanTZIDaHAHQR51TyAkTtObapZlbBINz
Ukz4F0U+nU/VwnEE4r+x9rTg8WntjI2qsveRPU2Xdz0er98ItLIXZQKhYGqMyFLF
ORcEESEZsMZ9ULftuFLjeaKl3Bq6WM2s4jPGR5iWL82h2Hl3/WMAVW5/R8rVOT9w
00ejkKCXe7/913+S9QsdYBhs7dk6m+/O1WtOvgXb8UgVD18YCxvJGv6rKpLTBzB4
D5LXpeHi3UHop3ICQaqtaG0Oe7pKfZUdUaUSi0OUV/piZxlHQ0Osxh62LcfjGe9Q
ndok7zKr9q5Z+pypt5p+WnMTw6p/m18UTW43qculKyHdznyaeZa5WgGvB+YD3BH7
iew5jRmr88rdCuBOZgzn5TYfLYrkeYZF9JUHisblp5+xDSEoqJZrAl8mv27KY7Xs
Gat2whA5ndQOfq9CTpz291mBsDI2lkqtery+8jAGR7bNYOeNVuHBiRbfkbwF6EFE
F1+Vn+6rHEhVwaldjDOGEAH5NsApxMJQSvKK5T3/zEVX9BpN2odLcxAaTSR82rch
S6EV5A1glcZIGJVRM8TlRDbQzZN90+7bTQSxCgQa874KBiae2itfGqR8gF8b9DhT
vRkD2FgReBrWu6htx68H0ll3hTyr5J8OoMW6DOAgkb0uitiWNa7lne9Jt2pMZtXI
68nheLdP3YOXXP98kN/lKOtXglTPq+OWvApKx94ktxjufdCaTZExlhI2wxInWDFc
GKz/1zrTsAXAfkR0s94eugkY7k83EEEF8zd352jl+NI09nAWmW5kxv9DIjkJKfEw
a5LD4bbD1HlQSQcLyBjVrITDsVPj6TR66t8PNGrUmxdRFTsiaJjCxnTSQCF/swvP
aWu1UYdT4C4MhEGEyDQ87tR3U/NDZJWPq6pCbfuXtNYM5JXwSf297cWGpM06Tb3h
oZfTDhcmLhixzWRxeeixuLU1u8wC6SaABTLyIq8cbyGUmoIfHbnNR3t1tb/MsQ7v
hQ+eKyvUvtm9Jj+CEeqEc93FlxRz6qPA/mZzst/y2WKGSy1XP42Haf2AnalkHWZe
3fjY2QpHH7zFXsqUJT01VSiCpCdLQsey2OwwpPVkmfRO53z+fzZUzc9SvbnnQBtK
KT2Meeo7nNeWbxLivDHQiYRhLMtVEpV2hNs/5IxnlHJu4pfdw4ocTR0FXUdO+HuF
BLqL08AjGLPfzVmGiOkB7ioLVw2hv1dz+/7ECVr2lWCHaMCW3NPh4eHgVgdU2LNs
eAiBEh2HKFs/OLWn1rb7zEltagqDzSbHDX7d4KAlMhGKFvtvbcaNcxLp2xzM1lcE
JoaOw0ey/Gn48xzF57Wjl/mNODG3dCVSXwfaeSkLEvGdFwCBhZZDWpyvpDbsA4CJ
V8ItfPor4F+0Fva/Hs2A3/pTr6nsHbnlbsF8jnjly5qktz7GNK/ehkTRvz3k59+r
vskYsNBJgA7VUu0NCgkmkyRX+Q7wxG9aqnlIh2vUKiHFx7N1/7SnydElBm7e4w5r
T+Gr4VCZlOMxfqpi9LJ9efoqpiC/DefZSJ7l7Wnwbv/EFvlHBjbB0EGyMHBMwSnv
xDlIWeEkOSA3VW/rmeDHTJ1eulTaHhsFu9pgJF2E5pHInOePp0Kq3DGrld32Ppr/
BLMZk9MWJd6drJ5pEZZXKWBbtCZNYQXY+tZ36jyUmseC0ED7O4K+h9a0fPkvOlOG
ZVA6WMdolkboXWO/B7eX4jIRHVyL2puaLUfcAZvIAcMzLoP7Bo4Jp0qnkzbseIXa
taVzMyzHCD4TUnpcYHD3Jimbm0S/2QD3+7AkDCVlyXPle1zQI1AaSijJeFxjqTDh
tL+aCAvkQITfagqTwVwZoHZo1KtRC+asCSnahd0YpCjXcvcEXn5Xg41xwF4cakSe
eGxVLn5TdSgZhRYe8SefaUDuN4F4lEOkWdfoRomKSZsqhnN9RfAW+cOCIuS6e6JY
HPxdp7/E2uFMGyg/agZlLM2xcrqttpeyfrCMASlF5LQtBROO59Jrr9YIiLwjyd4i
o2bWCFQbSvzeQ/nFnQzlD7F3cyJPc1SZX7RUprP+6UIdvmAaqdjlUg8Ld2p641kp
z4X84+aiDTJFmNli8GcXv94LUcA2Uia8Sz2pLb/8cX62AlTgG2J5nV9+tPPr8vUk
ShWZSmxD5YPvB+fQk6zC1F4afYekv8ClzSYP8l4Kgzh018F9chYLyPp/HQufwsla
KpcATcMqfR1N/tO7rvG/rK6hUToSSiErNlASu/FxITgJeucQeEJWhD9XCbFPsO+S
RCDFvMAj9qlALAYE3yNq65fknSacr4BiRBOFU9q0Z9KzE/DiLLBJSn1Q9WxR344+
PlzIagX1CRFzbv6vo57QDltfM/PTyJNGnaj014Gb6jBbWwzrO+eyYxooEbQ6/0ch
pKAayU6xNAzi2ku2r0DWfqEiLa0q7Z4qcPv98/6CkG/MB6jn4cHudJCk9iHiH2PH
TYVcbKtk0TL1arDeL2JtB/N67uLmeTdGPraQpxzL130RHWf4LBS+ew8uuH2TIO2v
nW95eBigjKcw1GR/APTJDkMqNh5vrFhVEeg2oQHYuQX4brLzbf6Z76I1pooknblZ
PtL0SFMB45UsoVHPR5y80yRTvLTzI4hUeO4qNTf1DmNUQeGDSEsrxa4KocNGNRhQ
/UhQORMNFyW7IjcHvghXbOb4R82V4Z9PNgCipJpKTCNGkKdl1sNbqV0+FLDJMJLv
UyqrGJh0L5JMoSE7/odo3qAi/T+th0eZpyUcvcby1tK79t27P6exKqBaaDuaUdvr
zMEk7sDqKzMk4ofDo7my952weqAOEJRRYWn4acSu64HzBBaLbQjWeLx0Dft+GY+4
leGSKAMQAPrNechCHTsWm632hKICh2DDfFXvi+L3jhmm+lDaWpOCpWg6Omsnl+FR
UAcO9A/2oR2V10kzJlJJE2kvamO08zm5X0ZhUh7sUugWLuxLqQjRERypt1FAMQ93
WgmJgSn2sodV2Wve1r8idKB+19MNuB6KycXX78HVE5Ok/YPEy/0Tt6kB1t4J4D4/
nE9l7UBRoYR0HJSXVKrOpyQuWVOvvcl9JLuF/PnhivwS5sm8EF4BuOdCq51t54bN
Ojk3ugjALD3K7PVLGxQOxJ+/QCul/BGCP8aBdTYwCEpAeISZt2rzYzxjgLBE5wef
D6et8sRQQimoBv5W5nt+zzWVZw06cQmuooFNymk+vX2V6MqYyzvpmnw+Lnf45Ekj
7LOAhxJED+DkhvemClT+A0/2i0oztyy7BUMrszgJ9dWww9Sf5Ck0dBwvqrtd5ejR
5lasawPd3ch7lOiFCg2ovEwyHzFov/aM99e3fFwrKgAkG4+dWh0H3YDuMEBeetYS
7FU0hFV2L3iKpVwHpdRKrBICP2KJv6S8msmwfya6LlGv6t1XLc2iSenZ2CSSlWpv
AETr+RmMAPdhmRIo7ND93NGZSDGD2Syb1bjY0TGT3r/1NKbpumyXMweso2lCrQ5m
U2M3xip/2xi7FiD2rkSnL3xKCUWrAA/DhQIe2K1HOvrJkFiaETX+EwWwRAOaMYJL
djfQxKnGazxk9cMqF/L9Jcjh1O0KpvxAi9b4b4g5Bo9VqK9Ye2OgzzgMXQg9AJtD
vHPT+Xi09MyEZMhBhOVFi+ii36Nmwqb11xcN+ExaY8d+Ou56cGMaLsoGRbWfVekz
+KQ3NHhkmrIO3uIOE2me3jG4lRd6LZBttCUwfWAMorvmdAyCvCrwCaYGLwXMSL5C
ZPF+90L1bPZoxKw1CnACar5N/jGD9Fb7KKPk8vhiCzrxKe9flykkCCWaLFkGUWBB
WTD6rmD7+0rutmDnmuoFBCRhH/+Ilta2cIm5cDCKi+RUbbNqsgQqEi1ZZWpM/jQe
t4/hb+QPy6HGb0U+0jyl7ycrGDHP/EXb8inbvTSrle72+QFdDTye674pRnPqpz8g
LzBB32GMhTX0z16NUzV1BU61Ozur2PcsVKpqAM6g0hgF9Ol04Hqun0EUfipkr1/t
CQ0df3F/+6YccDhc8wRvTexHgLvSoV+AsU5+u8unYB0GN/wFUiD5czEp+wwaWdCw
bo4W2bzOBGsijIkGUHhEU9sM7fGjIAkbp6qiSMKFNYj1dJHFkDxhoi724Nup7+m3
CSm78IGxsmfy4gEo9618hl0H1uS/oqs293c9kc1GeBQeON6JW+wSijEFXqwxnmXt
GFrPWUeDvYcL/z5hUZvijQ5GSJ6hQr/xYq5z4S7mTg/BhuriObCx4JX6JcWTRVHi
aFZhZgLVOqXcX2j6VxscCJQdrCRZ3Ust221dT0aH5xoEeCV3E24V0wD0QKUM47Mi
CYdqx70EwLo5+bVZuKj5yyrlQxXUlzLUQBkALyNfFU3tR9hA9vUhUelKouaeYMYl
3hUxuGtjPxYBp/R7k4sQ1gJ9F62m1uAqbEXHSHyj5E5iDOcXMEuSY55cUY4QA84f
LAKH1VfK5+uGOhElHQW+vwN0cqaS6eQQ/DL42UWH+a5+pTY3WT4yBMzAPRfuFlpS
70owFV7LYQsDrFQmJJFy2iGPn9FIVaYSSt+5nE8a5OXV2FxGU5hkawI7ZfuRQggm
PHD5LtMRS3kKH2z3xnZmesl+LG75ggkpA5/EzOMlcOfzOhhiGNf2kgJBb0g0fiqO
zXhO5klJ10ublHezIjOYlOuOuh9bWYOsludxzpevKAOJuXi0sOzjTZBRhNsgXRrB
JMLAew3vbq0OuI6f/kFZTS07vT+691d3ZnWDFwpgsCDwGILLBy6SSeisYx7EHsuk
/jGrdbiXuP2pU7Mf6xs3tSPh/d8xJP1lBRWTrMaATRbQqoh18GZ0z/bhNBtFhpme
nTsjCsKzr+6O0SLWFpGLRUGNIBDrk3iuxM9YBiJQzsGD4N/Hu77M9jUT9vrk+uc9
tVw1SBMfaYqY9GsqNQjnB125JH8rw1+1/9oRZLXLn2IeFh5bHTtqN5uQtdyaEewn
75T2GGBA5a7iSmTmjQ3TYcdvf6K2NshIftwq0C0Qa6P01IaCqg1RYfO6NZHVP0sj
/Ij8XeTOwfkQC9Gii0NwxN3xXcIDrorrBcAg2m0ns/t3mlnZmxciyEbpVyfs6HLx
+m+Ijjv2Xdar/0i6lumvHWQ7lPUMc8VWUvDvk8oUq9RB3ymjuhr9ap6V80jGQw06
skbNZcisVcz08/nhYrugoolIS7TSFajLxtGfF57JsHX2+VNGAttb9c2MgonBSatY
ECj5nL2czMf3jzto3N1VLLWx3zJhyEYqc6uCJaVPf4V5zTCFqBlh/5WDmhgFp+mP
RlJocgl/22O61gP0sCTKzGw3leDgozGwzu78pYYLmwsaXaTV838C/ZNS2Oy7cMMz
XZaP5SDdbsnbgKEuuIEaHgmlaRSd9SEzZRBWhehUuPPgqP8gauyDExECjF/dWZIQ
cIRjSFCQTJw16QQTccm+9NGAeUdbztiRBkVuZQ7VjP/IBIMwAHFLhoj++BSJXaAz
Sa7w9xz0LpNxwWIam2VPkxoktfh/8kbUnCJRD3w2+rS6rZ9TyekeiqMY7lUTZXHZ
TnfHQgMuE217WQ/nQix/xLi35CJdQSxalBmemBLX3JeqeCltJqiTKW7X1EtHJB/O
dXhldjYlFV/iMsix7fDOUPny4/W0nrJ42NHaKeIuc3eCuWljxG7hBbem5Mp1VtQK
RI48nU203f/Y+rzcDQrSuuKHtkc5k0XMvo5DDe6ZpLxiQOahoXanJeFyH1reqmAi
qXI75gs0ELzjGNWkF9UUHJASsx5qVz79Ae74fm7rhhe+R6Nt9DmP+GLM5rlw08Ve
UzZ6JBbcyDHpYHlfEugWah48dmiWZE8yyy63zXViT00/wIJI3qTFaDiGFiGHqr5D
yHrkARzUOIcT8srSwZWkiqPUuzYK+TNchsQfUN0NXwfIug6IjMyjiL7Drkr1be5m
UME84ovUnqE+116uUb1l8ZQdfB+q/2ob3SFjBT4bN9ICocStq9uuMrX7VXh1yQnG
okK7QZxb3EgSD/QH8C88jfe/s6w+Wuu+40NmPjVEf0I4jlRQuQZ1gLxX4N7Qy8lJ
Z5FXKDrvia5UN2ntR8LvHzZddYMJJa9N46uEcxwq5lPaLUmav1aTNYbYm/vgrMBW
NhQwYphsG3qBn6Qpa+6e2ASvoW/S7dOgfaGzBx227C36Qzz6ls5hpnpBB2sKBkLP
pTC+j7tBMCsy9v/IzfqMM7JATmAGih4QNxUylR7zdOCRruDFogTwHv1r2hUDGrfE
G6E7szwdSmeDfc3v2PB8zlLbA/WhRTt14+0Y7g86imzGwAU9rZhwrdCbwWDQ45DH
hHKzSVJQ+aBIz+TTYKQqvLngs9yX8J4YdRkySHANMBgD0yhxeAgVrtxRkiEvbYqo
T4pPtp+LZWdx6TTb1pMMWS05CH0yw65R2XEr0wPmDtXWzR+WWNc0TS2rE8PM9A7O
MyFjfWd032vQxtVazUYTG1RNhtIGC2iTSQXW4ZSr6LJKwNxnWvrDkdngXiST7wzx
6Ho0ZtzgBz4JlXw+LOW4ArUY+Z3G1pW148DDLj7JfjPvYWwvCJbbEzbT9e1nAj3R
zQU7/eECvV3Wk6WcQs0V6XojVKi4E0zuqcQ6+egNOhu5Tdcn/HulO2MgGJ39+prE
EgwT38KT4ZlVy3sE4GHNaGl0VKsifMMiVHBNd2zUuNSieumdE0wAGZhIhlknOlVm
XpzYihZ4lNV/EdUIuk5t1MZ6ZxmsobRT+X4JCSyo4bdDRG95ToB31R91lRYGcU8u
XCaw3egqcsAUDDnquF/iQ/ToapQOCSqp+rXhj0lP03FmSeDrfh8VIH+p0TfbgnDr
xmxy62S5dNttVK07YhQ4M9pksxc628Z2nUaBex1yI/LtHR8ge2oI63qVf8SRAtIw
loj7udvXesKVXg+XOnhxFbDtIpqlrcDbbkPB3JFO4ofWAlUPYRXs6G+BlFSaHY1Z
pzakWVsrCBFScyy6WwrQ7Dz3V7L7d1DZn6OO0XRSOAd+gL423gcYnGfCj8i1Jcu4
CTtQVlLoFIAbzHwTiLY1Bki6jfSRdRAABa6qaCQoD5kWVQvK9Wq5e7dpq5qI5hKO
U41/sseNK6JualKi1cTkNJI61GzJcordziWDASSf8vRkwo4JvN6Fls8vWVpEuh1V
MpZTsYOiAfQeVpf+j4Mg5gYwd/iZFeG9wBDW1krJbpcbhRZWDi2RvLEvOtFkUQop
Moaq1iXkBDWrqIS/fGrKxX8Xxkufzq5LS7Emw29uNytC49zKWFngsKt8sKomUCyw
TetgODq6cChfvcLCr9fp4V3HXZ/Wx3IWUiHn9z2afad8jdR9uk0fQOwqNv8Z7TgV
zTUOov6YySVutkeq7BiCt5bw5rpdKSBeKKtLUjR5Z4U6lMC/6Lp7RuxuQ+CIMuGT
jvwfpyNm/rYcziPaF7AbiE9zxHfhgFLiXGivNkkgtsHPSIW13CYzl44A8J2Sj9+3
UyZxegrSFR74oyQBnrsuig9GSZ47ioPfFpSD8BgG1V/atQIaCCltFLli+xPwJxiz
aGQZMZJUWC7jzCuhbP9EkmyLoArsCedp0/v9by0gvT8fhRz9W5ohTnMIhTY/Iat2
d3WjzRH2KTSWm1JH5pLe3lZXA5hO9mXDbHYOVV2qU6z5ZdXzb8Tf507E1O7jrOOj
cy7CqMP9f8Q+ttC37QgDEw40FdowpykM4eilejJPMRzazjFpW8Rdf/abUYOxFn+n
+4F4hFSuLwvctr/In4jlUHswLPgMXJedM3dSorQbwoEuTSixgmxJqchbGqxezRnG
b5g0HeHQCJjZiBiQKMxTgMOwMLPY1gGr5HKBimLlBUSh38JvI8ggoyk857UTwTty
h9IG7kNBVAE/KwHaCT6eva2v7Sec06iR6ca9xiqgMd81VC+DJnep2gTs17d/y/1R
yO/tlYzfnFJzxIIiQt8VS1OUoGRqUE5gsjQHqLJ8jRcwL4T/iZTAGVDm/vj2eEAt
kgTqkm6JYOtalcT+7XKOcY249tfIAFrzbxH+UGCu+HWRXNVTmdiiUd4hCE5+0izN
4TGmD4VY3c0/LN0Yz1pNXowJPKUJ1ZAVsW/1hydMgcNP1e38/Q+brFzo7120WxKJ
rOsst67svnGZsXUUa/Khgl3VK91jFM6AsYGr69rfdgQ8lFmv/IAB8V+rXJvDS9hg
rvFsycpwDIZOlame5Nzm+4Jglci0HCFnXMBLilraW1yIhZwizI/JAcGnUIoasnCm
nZaaweoSDQXuXJ10dmXGE6NpHSUUCj+udr08WkNybtu+SIZhffZbAjT17knxHkVx
GJiTFasPBeFXazQgEJMjnwazPjcbsFuNxPoYWJvGxYh//oxki1GpvafZJsQgJh9/
7kcVT6PBwezwtIIPeyh7ejlXCiM2pRwJQ5ZINbfv1BV9T0mAR6whi/ncE+eTsC9/
LrXPTCmzCumYrSFb+5SDD7bHf4flDNHWsZU7AZUe+J1HAEiQnax03Usl/AWPOiMM
duCkF7Ghg+uvtOJ7kEXI/AI3UaxrI/i9zqweKq8WWZ+mIDE9N3EXArulaFKq9xGQ
BU3WoTCo4x77CGQqAb1ZAEMV7awSLmpz7AYAQvimQi9QPOZrxldrJqwqDVslhsA3
vxyfJpgRpCFzbU6xy87u1YwrYC0DrEhk4UJSkVHXik2t502U+ONM7yENeAAsx52b
dZXnlPUm73TjMRVSWA+fnPeLp+Y3Jg61nIX3auSuGSAGZFMnKrYJYcDsR7lc3pNd
aYBuspHJiOSU0PH40Uj/a2xwDxE/14ozsVR9dYv9V3Zy1uBvX+4uh5YaOC0mgfIo
YEK21Rqg7frSOvWwpSkEQfNCCJ1wSZdVc71ua9l+2ERnvkiQf0G6Dgo661bu/Mt1
kPpskP45dpORRUu7VCp6AIU/JbnoUugLgQhEsgXthuCn8m9j8Osv7d3F2ozG/Qva
u6MESWN4AnfjokazvM1i54Fxxd0IJZyvyN6pYZjkD0F0QJ9Krc9Op+xwIdBpV6ve
UlbVq7qLAv56/AjPvgbdR9phCZP3zo7376yOnoyG+NcZ0e6tO5hYeTUmbcnmNvFM
5MRdSLljEoPyIFaBIoOG88BFR+HTDFnQZtfqXTi5g+zs/ldDFmOGt1pWJp6/ge+E
aMIo3bgbmqChg00vXT4ExWiXK0ZoqJWw1eqITtp7il5cblz0/+6ozI5h1KgDlOxM
H9g1pt30rWRrsSn+cGY/8iP3fam8IxJp4cUzSUzZps0kZa7FsBJIP/N86MRuxEa0
+pR5GGx2BdZshV/98LdD1/uimSXzoIIdOJYu/rXirmtfVBT48XDEYCQa6EYxsWVl
puR9oQTIkrQm2o6O166rTaraUGdj7RR4Rc4Ue6e4WcoOOMJrcKai114FF6cx3ol2
muY7I9s+T7G7yQMyfmGTATf/oUE1G9KytVslRWTpr4jjnybaFPL8kWuxlqahoxIT
C5lUcENnXR1MB98U+z0M6UldB4hyl0XlWIYaRY/uSkGTKM5qk2mv1hdnS6xniA6g
PUT14KOfTcAV0szYR7at1J//IzlvWsvBBszbl4Yf+/x3CqfDDpOe64JCAT+/l10G
qdOxYWcttO7hj1K6ap7v4m6J/+kAL5+RVvqqaKq57FV2vIOxpRdZM90ut40GOTau
kPXvUvPTmeeiQv0k+EaaZTEX4xpNrdT48qRhMjnJSfDpaS9zIuKZohPCPmgRBwIw
6tr29oppEwqsVF+frs1mKtNiXDsxA8dZE0LUkXx8nrwDa7V2eAKp6lFutVJKzPHo
VS5H9GYzn9/StfwOIH9o7M1vqGOr1GkGTAqVJVausiOlGI2ClJsLfFGmXdFUQIsM
capID3wSyoEPqU1OPL5sBf8IBGkojMnVMimAt3KjYpyShOP0knsl2fgBpBp3GSCB
oTmoY1xyCETk1Sn9g4F3YJ9A+terC3gStN4iTLXxjjRb+CthhgIbWkiFM1RZgSUq
DM+ZzQzUu4qVQCa0rnppFyW0PT9Vum7BcoOr1KCTEXSTKxIVYIMShsUzl+mTZpcE
dRuTOIlCmq8showfakM/ZAfHdaOqiJBItxJWyoHGDHoLdpI1FUMM7gVrE/ClABy2
wax4fp1VIsO8xJhQRFsKkfz/i5oH+ZM3Wu0loI3JMVqWtZyyiM5fv+T7BU8J7Zwi
B8rpYhhzgsAOhnX40XSY/Ojs1w8dB2VZurY8nTHrX9WVIzMT6uENhc4tvDaBawrT
Tk+fAOvlm3yVDkiekRR5AScf8P/6HPXdu6URfjNbfqV68RMMR6NW3ShCEMyBBwjn
LfniVmyfrNI1KnV1b/TfmXXtsRi3Vx5p2pIAOSnGWWNPo6ExxRfcGY3FkBXK4+aB
SU4oBNPWp/4w1VzuZugNUsWXqnDV5IbqwclkYw7ro/5m/cgUC2w4ikz4syFIyFdz
DEsJmRyHyxBpf4IIgPSjeHdbMWWoycrulNaxVxnfmGUlH0AoJdtdeBelmxn/Kwd/
B8dJ5bXaqCI9YnLL4Kl7m7DCzKQSjy91m+Xi8mdehBXMEzzNOZ1+Hbw1y4ymwOZC
YiFHEeAatU/u2Sv7jPURMFeT8Ift94/ebW6OGcD0TH6WPK+gn2sQ8YuU7udooFVV
YOUsLu/95dW0NwTJMRD8LrQGSrkzHBohfOZK6MqxW2vygY1AVHp9lW1QYxzJub9c
6N+YlDpwJer0dbkrDlEbClEv/wBgOaBiBZX4lllid4n4eCzI7CZZrV14QIQW55Sa
+Bpwu1nlHPSh9VHEdhy6S7bcUEbQPzT/bbggG4KUXsaOdzkegdvKiQ+AL8WQ3noz
iLC+gRxYqb8LfccRLDIym6jtTuh7tFgI3+Vaw6jSnKnwi6gf/VRULMu73Rhz/IPg
YSIK71XZ1MdOFpgbo0CmVz6ThmK1BGt4uVJR4tXYu1ryBZlRMtXPGDrmCHVi0D1L
bfy5nwgHLPvyx5D6layvbN1+sAaO6bUn6B9z6+mvNVA49N7ZyKNnXNWCxmnrsrRA
32/U7uB4EJCNcdCp1rzvwZ5/GPNd5Siagzdul1LPupN5Pxf8FX5gK8yD/2M+dST5
vPwPTQWRUcIiUzofIq1S8shulFqq4mZhAWQ1rQZIz+IsdnDXUg2o+Ak0Mm2BrCmy
EfBHGLgxujbyqMCvQ+yQ/mjmCfZq8/Mj+m+CUkGZeb9Zt8JTyCvYQ9gR8TSQRTzO
R7+d+x7q0WBeF4h6VQfNbk03BZcmLuGc4/3uw3HC3igwtsO9s1QNSpA8jLONsOtP
Mo+A2qJtoSqBqExsS8YAr2xXoUYIT0DnYUzF5c4UYY1hdlGwO1C/5VLFyni4UVDF
UWDUcf2SJBxffjqz80s1jnCS8XK9ThriAb1pHIzGj+MMWi2ixu1V3xpmiS/YHynt
nV2O2Hc6B33ZuTtdySxiMXhuJ/cNG/nhqMaTwzA8WMI9RBzcU4sOjm/ywYbNvagT
VSeNFQn1UxQoak+eRCykxa0D1uklvJj91bxAdua6iypZjkojhD3QPNKC/Ew10VHQ
ukULOTGhRyv/Cid2rixrck4BDgSIiztobB9cOo80rKszziWGsd27Wri/lRp3nOzG
c7mCeAfkZQcUIq5ex6a9Qi14zrcehroDCR9AW2diVkG5WPLEnwWm0dxXnWP/tcBG
XK7nrsVz1rvgFlAO/83RCh5MKSyl5rspAqo2+Pr/yM05vzmD6w+2cRJPbxSnOuvg
QY54nJ5qdRNXTs3t8VXwip7II7/IcseORQCf7whZ5oF5F9tHSGfiNugBezt/x75C
YuZjjgwNZy7vCA++9AE2b3mvJhO6vwwtfNZl4js2ykCDUo5pyP0yVMq2Fv3V+BSw
p5/3bUBUdDDaizCvbgmTPIBuXHJUmsXpQjJK7RLIp9u2ZQc1a4C76rPMA97Dfnxg
kMtYq3dyg7dAz+AZpzUcsfbvPuoKCIoyNvPTl9HZwLTYLkIi1fd9sw7tTVmTbeOO
fZTfSEZgR1A0NxHfWShlFZSga2+tkz5y3Shi3yoxBsO5kn5a3eoVqF7kF6eCWdb1
7JcYHUHbbyUaw7De93tdBm8OXZ6AexjP9QhynRCrwd/LdjsWBycoz7709ixlJy7l
REMhkx9XpLZ4heVLHrgk49hlA8Cgdr8VMTsbwlTtZmd8PNOJDTa9araF1JSAt5mA
K0bhBc21pshFD35UT8imuQ3iztRQFlOdpNpPtMrfuIdf3meeZiwUpfESADrAUHj+
WzRKgzf1xG+y0RLJeVbYp63BKrTwrrsuqm7I2YzNWX6KNJoWwavgp/zo+aq4YhQa
t5+pjdjEtDOMwfgX/nY7pi40Qi/4ypjXmXoDIdZp2dZ5qFIEdPpAjb8F0+BVIt+A
DpjWjWaDvVNKOVkwa14o1XYaXiGVkgeIFsnQJRfjA0e066egQbCXWV+vZlCD2PW/
jnN8JwQ8klsoxR4hX12sCGNP5FXiF57LINHM+oBbdYxaZkA1x98zWNwxrwvoM7kM
D7qtJY+BH1qiKWLyRlPOJ6VIgb1yK7Xz5PLCT3xZWZIXNaqBGrVbplHcJ9A45pv8
TQM9BvAxPd8BJfbyf87xr90/E/JPDVCJ1Zd+bA23M7YeHY5JvVzIICGs3MU2qQp2
sW4FxAy35OvLXLyBIof/4XGqR1hEuk9tAbaw4x7xyuP0Y8BfsaN/CQYEUnEAcqdp
q63E9kX/jZkPg8fz7YIWCj625u7YvfnpBjf77g88h52KPlSHN9SDVhpQfWvVeqCv
aTZShAHzdfatf25oZKpQ8PpfN7+O/nVo3peldoTYfhv8/m+bLXE4TzQrltFyA0zN
8nuACziNnMPM1ECJ5KYglNKLpGC9aI7I55EQhrfKO0812geDIYRfNiEILpAbIrUR
nqa0EWwFqZR4BiqBekGXxPATq3UoVDxi+gM3lFcet3hL8NVDiA8hxnCdSZkcu7nL
jNf0h8687zLoBromBlQ68BOrq0QLl1mh+nxvawIJTt5qak5zqGI5zFj8ms1eva7c
Vayj/DkkROIkXLeHW1ToNBC1b+5t7nc1AKIENQtB2fTZSLDFApppAX/KHx1TGc73
BuFFxh76vho33ajf4GVlc25ONyseyJ1vAaMM+1xRSJ8PXOJtiVDyzUZ1vE6DeZMx
iNNsTmkRuzuI9eqlZlVdwFJx0b4q91VW9CdpyBAD+DHmDlQADL8EWvr0SgQ41ojp
KgTg1bvN0BADEyhUHkP7cpSgic2FSkX0OZ0eKpAHMD5ZuX3ti+VN08iU0dPkonVy
zjgqUtUk7AjK6/4302Jcz+aEexnDrqzvosHX0N+MxLrO1jwhJL9J6dotAhHH86pn
GcSZYjZUa/y+00s0KRuuwhvc1F/5qfxoUsjdJSCMseIwx3r2Y14f4ylUVVr98mAr
UzaNcDaYWLK7CYoBX0PhJe7f5g+vlsCyzuHjo3G/+f7xd3hI6u52Fe8/4aWTR+Oe
ditZi1K+xgraUKAbY+4Zl5p9zGb8yKuWvWkQHfKs26HG2p1j8QHnMVNoY6zrnBT+
/JlTyqlXgUYPq2aY/oRLb5h9p5wrcaK9x7yj7IQRQ0H9ECiTDEg4RCbi6cC9ZUCV
k06trYrc0vGoJvrIEmUVVgLI1xXG7IsxwWY6RCteh1+xTNqZCUEgYFhfHEsqgdGC
s8BdCD25+2xfEUjLinW1vTBp36xsaDNkCF4yLBOK6iPOzGBeyPp/7urpl2SDY3y0
wXDtyX3EtSayHqo1nJ3h6lbDyqKOC0Rj+ijcJHrA6aU64MnxgTB6g7RnKbUY1pdW
tm4KaKevCYBFQYk2BzZ2HxYhtbs556LvbSeNho5KnQfpjZnBdEOeWSc35EaDLP7l
/192hxGwAc6b8XNsWGt2aB3Bp48HPrQJvj1Sz5oYzSIITa/BmGftppXKwxSudkJE
Tf5HCXM8UZfdtHUBM5KwIJiU3ZHYbkvEt2gGVywa6KXcWmtvH/ki+NKFiJMxEEbC
CAT14zwSRuDdjg3N6wXeFTGO9sBQGhjAilELZJCCJ6omD0w5irKZk+8rFPrJ+EnI
jBqzA44u9NONHYkPJRgPLEJK+JHqHq+rV2dF6szCvvQzpHXYAqXUO9/pk/YYWmj6
ssrMldSDdEvFI1dBM0bLciYKy4+i+IjvxGhlrh9dELIo+OBBHyIFBD74e/Rq9FYq
ououYiCTyddI2NFiIHmxcmuvIfCOrxoWPS+1jHZ0Bw86RC4JKDkoh+8imBZuwGTD
/CCnCpA24ELpFaP9omi53OxodSXy3v6+dy5iqiHGuX+/XT2jFHJczzzrzTCy8RjA
//sng7u/oSToafTSigHujRD4nGQhf3eWBZ+xWxDG7LxL1bnKn05w+cDfRFo6teR4
DrjIHjavHsFdgonSCmhJRBnsWHSpGVLeJ44RUa8fI6yBpgyHvaFBoL20NthPjVYT
vWQZfBSgcl76keyHkCji62yIc4zCmLtk4tmKqr1RGM0OUUZdTOzpKX5VLv4obthz
56THpZWO7sWXr9nykmUW9mjAZZn8ed+6QV7ESBfr3cE/gN1JhHAHavL4ALgjF9G/
KVhF0WMk0eSrif4Ak/1W9yMGBXTBW0UyABzD20eyXTewHkD/OAM6sOV2N0bENI85
tKCk914Lu8brJ6gA8z7Lhut3DhiT2uUVcWkIuzBFC4RnciiFAmp5dFNYgYGjjaf/
4xX/M2aodHPZl1n3NiM3V2c/ScEe2mJKh+ldzhNewFm5bAGa6ImSrMFz2zsRH2rM
r86wDBt6LXjNEQHglQNw9p5JLyxsSmM4SDo9Bdfr1HN7OPu/1MunXN74AdyxyUrh
2XpSkYrp4TZQ2y8qaq58pUp5uKGH8fAK3c7XaRWVGupXsu7YAAvv7zs30o1xejKB
C1RD9o2k9lcsFshbhRROjH2Hhw1DqIyo9EVUBrPfK3rjtRQ2Prh+9HJXvpspme4t
s39ToNBjUZ1lKRsYpdF8xtyn6yqDayOMVI3lemesl1+pETHYl4OrFwRGlWKLsR4r
89Iq1e3gJksGQymQmPjuc+BMMR12GawjbLiyOlS/2Wpbdi2PvTTXy4k0NlmY5aum
cgMDFiwqCFSoZybyhAQNBa4YsdnqFPxqY0QKX1wy+Lcg3g1SSAHuL1ftDt8ql7qX
PxO0nxN02IvcBlUFlfEFab10LnIUUC8FeU/j8HirqVSbyA7s44vTQrq/dVq2QdXK
p4j7ycIWkRGPgFvd8ZBjljfaSTepvNJ5mhurNEMLfg0meorrgSj34zVjCSrkG4+r
xrCRDSU1zzXI+vYs5t8YPXeVMG+2tkXBnKK0r9zm7C/ki2ZJdI8hIfJr/JgV/1ej
OZP921e0d1mk9DElne+84c7r73104Oi/eKWsiH3n0/DH7jTZpzbpUxs2Bbzu5nUK
aFtpp5p8hIgIZ2tDDcUp3p/WHRfkqyKcov2B0tx7bkylhiIouDZOaSj1UbPP41ww
B34I+s4U3eowcFcxLPYHneyPBvlFzx1ablS/pWCE1O/YDYgXjGk0TSwFdh5cW3Jq
KajnkD8eQCDkXBZ6/E34zyiq90/QFW1/XNVizt0y5vDJFJ2e2AzGwyXVNN+nLeQw
ie4D1gdW/hUVDSYbEPiOLDd/ucHT5foFXeS1mB0Y4AQXl+rkrl0Pgk5gdBqTaQLi
lW9alGB5YRGemHjcoYJBi11f9l/gYI6aqGGBWIpDys8NGfFyc0zgwiqBaYnqsILV
6YH65fvm4R9pcNT7pfiky37H6FkKKUF3Ykip3iWvZpAji6PCUdtcPKgiLyHiQJw9
WrArfMXrDjFjSDns7wf2AsMjcNE7bKaYACJPtkyZOOkGP8PnHA7g80nvEISDYeUJ
SjybQvmpWm1rn0oC8ljmbn2JAO3ME6nFkAKskpNDN64D0vLOrPL6kkPRVCVvxlc3
40C5m+eyWsqoLiKu5tvMpqw4qxzefGrB5P2t2UoNrg+NBlDHNdiyzfAamUQ7E3L+
HFjqgVqE4BZcB9d0cs9dWzrwMa4Nu84HgKm59YkY4cerZhl8kJIsvRKKQZvtLKWt
AfkFGtIy7/CJ9igm0OOt9OhOpwrjpjL8SeDfyb8rvbU91kxPfvrqVSADEWs3eb4q
0RpojV4pMtEPairSElKz5+IBQhO1JRmnfsBAnvza7qDwv3seqjkg7hhpw6JNawO5
z7YokTyuf1jfc8xfU3XlxvdQapnNLTtzOdymBgL39zJQzDwtkJRF+5eKy2cYAqtN
cBBXLvSgInSPG4KAgB6DoAvAwtLqVqoqFsEke5yXj/Rjqz0Bfq8pkumG29if3HER
ZontFKWE/p5h7aJmXzhNZDksDOGINe/KcE2i5eBkKJKWXoIugW65REhpBfX7OBrV
4dIwF82PBOcSnhDkvqaXMbXOPNQLpoWpcUOXI/ACRmUwXU2u6vMP/NO1wOP9Em+0
QRUwhsBN1e3JvEqmxSBqKtmIGVtbU5mnUpLohxL7pRvu7wpWbzOI7XS3aP9OxhT0
bU8ixl3UYvFmvXKj1VKvmzFFMzaBO4x6C0NCs36RkF5ItBCArNAE1ffj7FxS4pzL
GWq8UWIcXEIbWO+rH9+0JINi+TJ1SAsR1LrWAbe+u6x/e0SjtgjxMExq6DfJ/Xfk
YqVeeHkJ6nvN8+1H8qy6OIPCVu+CCWlVpulOsp9mA2cOx3HNGeN2+GpVojJVyPhW
XtOfy1dgTIyTfT1oq66aTzY9udmo8SE9jyWQjPcCJb221S0LZQlZZxXzBKtrrTlK
Z1SWVUKsmGoNs1GlTutCw73F2r4iFZZSa1lTykKpVbHHvAccZnnKYr9agSDfYJzc
pqk11EDZxraR/SDP/03TAZz53N/dB1lCkb5eb0SsSeyel5eS5IPyd7zOFxsax5we
xQK8k3u6W95F6SOYS/Eh1+gtiBO1rwfzFivdyVxCSM+HjJcITCC3BTuAS8quf9tq
Gfg4weRjhtQqUaf5Ak1TfqJob1bKQtl7ufY/G79jbk/0HkUvZWLDQ5lIf7jRwB2f
RNgcH6/6+hdWidrn8Y3PNrzrpJ6qvFiic1egMiMFTlQAKSXKDUtuCzw/O7KLS2Mp
Q6mb6S3iTIRgsopkHfdFEqPYVIVotI5OY6cJo7GrVWPHwpiRaD4o7UGM8U7zOxaR
dOBRWavYxQBHirK3aNxX/wUTLek8rFRXWr+RVcaOL0pofSsNfzBTRCBrp1kBr2o0
P/pLO+MadiOtmHxuskzYA+siGXLL7TEMdNjUw3+URdHgN/8mCwot2TAJ9iMGTFNg
/4cUfApaAnJ6BzTSVpNrj6an5kRYdH8Df6JCDEVMH0u3g7X1+SiyL5iHpqzrMGY8
q7ItjuUGqz8JACx31obbNDNVXk9JzcI6p0o0wIYHfmBCxJtkze2OFFyXgpjDfU9q
dSh9bCqT/M6F3TrdWCmZCMmixOzwhss5kkIsem80mQZ1Y0FluPPfAL3aneHuFI70
xRjtW3jgmThXvp2ku6tSHSQpUQoAakdb50cg6hDEs9BgsSJ2UqmQFMiDWAjbekPX
KHXLMq6UaXpJOkQCgsaGmCJzE12BD3JVVrnm7W1Hv7YxDHsLeeDvLcmgH5e13UpM
4ftI59iNRs5xdM+QHEmn4hvQyLMWRMx3e0KHX+2B9HYFe/93G+CauLyIJ2XwYlx5
jV+2f4kKLj+PAnY67bcqwlwP6H/vJDwiCKzGhDiaVKaS5OLgyqmyV/HkSHgiXbYw
PM3q6u3APU9w0C2IWKYFpeJRmtHYwKbheza+dZSC1ou4LcM6bJ8xgPlnt5eGHyVv
3Bw5gdCXRa7x4ch9DL5XpoyZ3MjPYGflzvt2/ycd2pkyCUGaHjgn8ueUG3UlpNbx
z3tlWLfkeCq6SxoebD990ENJ6jAd5IS9Txg2LKoN9KEyQEUaEPel05xetnh0qk6I
ywHur3myCgSsfZPJhv6IvnZ8y5Q3hvyhoklgMuP13wakgXXysdKz2t8Cx2tZ9qeT
5OUUdE/3gpUXl7EOMROkHHm0bKGPg9kWRo5LnXZficA4Ui6ATARlE4Ef8Xu/eMA9
qFHq74/xDs+i2kumnPalr0t+6fAXNZ3jbWXq2otinGd16Yr36cInsXKY46XUBtc+
0agNJ3VpfwHQmjxW5Zpgjccq+eijXr/zzIJinrqB/jal65fCX2O+I20OKTQESEwc
M/QrJnXFOvvjktLY1vwzIxbgOMrsvrmrVe0adg8pshST3x9FIiPo1cFDiL8SNtH8
7Y8psgyIH8Ptbv3DYXegxd6eTFqEtTX2JZXfeO4mQI93dinbaBSJYym657eXiw+q
wsSWMxqya5MdBkbo2sKprf/BSA/WJFA6JOLrphJWq3xmbdr9ZpO6NHQnfJDrCht3
71k/V/cf4l2CAxNqnMb/AjDOfmAKxZQxQXTfS+N1CR38iERIp7xjzHf6z7lyQTeQ
tBZZIOz9TKHkI4XbZhEk0dbim9tQjxFqtKdvfS18SmvYOB9RZSRSaG0y7/l6hBlz
jmxONZ5w1G4FsLMFr5ZGf0pbOXKYn4N2bQghaKMVeKwmpi/FwRHgM62LPOKsLsb5
wdGIRiMpDs24tcXIHLyQW2dm57EXZNz3q77wTuPAjw3RrIN6ndaAK417+t3z48/x
m0uP5xrbwcDJWjWaOj0jt0oBfGg37S7q4aSG6hOq9WSbfTtnKEMp5tFzzjIbGY3d
/2axtZkBka7WHznTu7NLzkABmJOa8wYLleAnpAtwwAj6v/lbeHss1AU8rGATgLC3
/KMgu38jkreK4dt44abn6fl8MggL4nsVuO49sMxXTH+mBzEn73T1so3CYUXBN2eN
dZWpuniatfEPnX/SAz4Onp+O8XXUQHcY7uQl3cVeeq9DRwtCa2zthTrTknzwTfuz
0y0Fd7UY2Ehr4yYCDdVytrKELyS7mx/m4lxJO/4cPtgG9a2X2gPDHJBteSDqpTcS
bBv7YNJs+lzl6wzZY4M4tfE5KYpvNE20YLfA3vvQuGHrfKfSwwcecJGiurAJTYZ+
LSHVmX3kxjOVKKR9rZcR5NavsmSbaFnOkT7DJBbh0qvu6JHz8WQg6um2gtkmx6rz
7Uwfk3CigcNAfga9gR4bELWX0uUabVFbxB6WhnNWVcRZLKQlx9lmm+F7i7c35uaB
QtJP+GEJ2AYM13MzRNggl3hpE+z4yhPyILJLDyeSzJRpQ9mM0dIs81hJki6+3zCj
eFzxTnVOhyQY0pmdyvV2UpkclzmnWFAHm0xmYx+4rIn6OKriChIHFCINf1sra0dj
iGL4dIV2r9TAw2U7VO243rFkXM8ZugpYEpODfpS0wxmYt0PrnKcCWxZiY089djM5
6OYZuxWAwP09KwLqmKwvAGnZFsK1QA9vM+LJ2WYXl4w1jmlfLllQX/+QiuVdx7SN
pHHobfFcya1lw1IPq5hS5NkQYFN4AdPlB7otLgVoE3Qe2UisXvx9fsMDMrOYHbge
pkAXw9w4pUeaxTdZeOU+d6g2nyK+Ih/FyDekHhS/QpB9aeRUtHEO/En3cPt0dC5z
ufOE2OBT+6NxWXGF2aHrLOLSIxbJIqIGZeltQBKDADoqizYJU6Rk2mFQtlZFfokM
grtiyXRxM7PCw7nq/8nTHBqX5xcK/nl3US5+4seHRMBNiCekxbNzz4ulrSzooLsJ
Wzm5ogv/qCQNtrnOjNx7pFnbN+hQiNQeW5KYWIMKGBTz5KSsHjkJdJJMBeFvk1l/
ZYmbzLGQuXLnpmK6p7j2U+OEy6xOrQrUeuIlFSbJD2I7PhcGLdcW+T9RMJ5lVNNw
T+WYznP/2ht5S9xjcRQrWYqNgHCF0dadLZBOUFI6kx/aHvIjtJRX/5zZj2NqCZNO
+oFqSMfgaLiO/7y4w8ACuo+RDGTSRumlvZblbynpvgsGt/sfBZby8/WUEVfo1kzS
fNP7zYih5jxCREAvV/xVB8UpzTIjwPwa4usdY4J/2AKkooe2rMkTfEFDbVCDmT7A
RI8tBXeQXhaRUvvkg2xJFZLQojLBv+jVToiLL1dPKB9omT7gzlOSAxhS85/du3BQ
Z6L4oeRaA1RCCQPBopxxS7+ilNm+qFM7kHx3d2O0iu8GEztfNbVJKuyrQkrlvFdz
9DVDDKONDkeyKPrLrKj6bUrTntxjbwUK1rmR+jhCF3OjkIS94Cryk6NmebgQdXan
WfpyHeI9R+N34T2ACZ7om5E7wt2UaQKgNGe6xbfpuWO4ITFwS0PRCRduPsY5ekgZ
nV3dfBaJiy86rtnX6FcCwHPxeI0I1ZdD/i1nmDOX1+fxQFiH8QjXlyogtZONjPrD
1ACHThzZW9HhFaCfg2AlxBLB9mcRrYTQhrZoiL6Kez3s28WoLyfkohQCVdfPJWrh
J5/ezD7n7769Ikh+4DOfQRJeUmxjjxJvIa6U1jBRm/pf1HFtgJjbc36DL39TWaCa
hYCjwTzhx6RpfZ/lRbtt1AgYrKduUKCXLPXeLen9xCuqWOyyX0dxhteUaI4vnTiS
ov1rDM4xweg3fWhs2GnX6OQ2JPcfnY+vwlHV7y6659FpNdiVUZSiwydHmszu1qhg
JcmJzxK8aefkqQUr3I6gTv38dmvFS4KRxEKuUCt7fL7Dx0D80QjXtUWMvyZ06inf
UbGmllu/7POB43F0f6NWUm7A09/nypTOHk2xefF7YKZydVgAOKyyaFof+9ZxydZr
E2094jtdCfKDzI3BvWZcFcT+hFyRAZULzzQRPlwzbNZXG4nVAhGTPaGxXX8sVnYJ
Wj7ZNK4/Idl6BV6PNfqfTgrOyi9apEF0L67q+ufa0jLLvoFS/2N9pmXH1yWb0nrA
GjsWs52pqseyhNIBMd60jFZe2/1+dtXGpwOt0YcY/bE+vXzpuJIHrRRfIzSxZdsH
9u1T9wV3qgCgnM5EMU19XVRUrR2zLMyKLYOxIJJqAC3ulWc20+bUbOXvBqjUAgeV
bNI/QKhWwtNv0Mx6B7M2WZ7/tKyA3Jro5jJugGuGM9rCdtES/OXbK5J8bmy1Y+Yl
Ig9EtYRXcwgw+w+l3SkrkyLDCIolqy39g7AztoDOfKAnbh375pNGjUlXTxWb5ps2
utj6N421GTcW/9Fa2KkrkxPnhZcfSH8H2T9mMZt2Fiu7XsqiP3289qQ4esMBx7zD
JWYuUgievuLL3YeKHTteHcHbANOwMGKhb+PialtDcid8oLQLcQU6QybvZ9IZGUdC
BpF255KUo/cFMywjxMcP8bzAdmGOuNWDNJG2oM3p6a1P+Rh9YuchWM1ZvjRqSN2L
qYKKDoVA4FoOGWJH4M5MnCETzQe9iJGl8QvOuXwPDSSK43joMWGPwKUsYgW73OQQ
9gpTg90F9btrt0n+PcA24O4UjmdKrIe9fPj7cfP5YYeTZxGVyt/lIMm+pbOLQ5SK
8WO75KVVp2RJ5JyS15cQj1b02mMcbLUZLHF2qSMhNKVOaQJTk/3s5uAlLyoG4BD8
DeOAGjNd2OBvmtI4Z4nBm5hUx4Wx0I2yQcZRer67ikoWTOew/DTlQ7FE7ehNS9uQ
wbc7htNU8Xoq6XtdZv0zHqug4tUk2SYvb2nUSqgjYKWdifm+zS33YPACZqaOdDd+
RpjmKNR2cwS6tuArjLdi3Uaa79gM5QLwdQoKEdYFrohP2Hv19VDla6tj1b3erIUK
8/d5E/xwrrbs+l7PzSl0U/QVKMLwMmy5QYXk6AdTr4hNQQN1sayuW94cnRSudmsJ
A5PGNeiB1bZZjZqV0s9NaCI7c3w6IG6lyYJb7uSSItKauJuGYOYma8i2Kd08JttF
7Odupj3xvD4/hK0GHGfyUXNRd+cE1Gn6soN1AZYMooB3NvQJiPalp8uHjnkAiL9Q
iysz8EhY8+Y1gRBVCtTh8uvFHbiyFVKP7iBMIFWRMenncAqzPUFww1wAgLOs2UEh
uI2slGHoV+ix0eLA1O+S8LxmKA/3OGaGBEYwecI3ahoHI+4ZMkbXcnVd0fSbmpBG
EXyrU4gElC7d/oQSHpfRV4HmZ0eAVurql1+6t2nErs1kcbZ7nPdxsPRxYw0YIb3A
ly6kj6KbqkD5AX/5WBbqgtAlliiRzhcrKcGstA5M3ZQFCkqn56z7kG1S70G+hTNA
8x7vaIeQcQBbAz2JfIBHc1tqBoQcSYxXNC1GEv2z9qMaX5XlwGx7/OgmeY6oA/LA
s36wn9n6JSyWgBHZhG2oUGVFxdmIZA8T120HeCjGWBCKD3SKMz0OwAIHZTloXeXH
F212aLH1eRAd4PonKuK4QsS/gsT5k0z4gdib85jxNZhdUAuAqH1hEyDjMtcqJXZF
y0DcQk4dTYL3UPqzs7HTC4O9ec5qLXaKPo+duUS9VscB5xCF2mpUo45bJTiurjmf
i8FxNzCxEpk4DUeP+feH0mB8zKO//5gkhswYq90ofolGkqr6Odj0eo0hDw9d1sPx
6L1F/oj3yNtcKUmeg0jgCOVs8TAmQWd4+5gfm8OdcBZ00B5UoXd3QjEbbL/1W3vQ
HYgJXrLX+ZBX6fLURX5Bs8vz0d/rKVIls1DiL4YTpOc50He5yoc+dK26cSh1Y3TQ
kIP1hQVLY4ZCH8RceePggoZU3we3Ehz6JODCL+1AbtLwhLxwWvzp5tmE70RNBJqx
+VpLPxb6nfjIvtXjxNV2M78X2qQ0RUjPyH3XfyVrh/8h5Rx/WafIAMKsCCwM9vDR
Ypbpr4/cyhuht3mWBZzx4MD4Txy+Aeev2DOE20j0v8cCLcnk8E0TpdPQS9h28LeV
+wV+S/3KoOatbMV+je0KOYt2qDMBz9dGbdng2eLr+Ir8jy3iojRZ3ft77tpBxcWJ
nVs3d4pl/pdzwG3Th6Uwiuc2SU5o0AsdP4kDJHvuqva+NPTsCT1eK2oDp5mj9qiF
+xGErhlPM79fjyPreiaWwAQtEYVkAyQs9eJY7ZuW/ickQkcDylDDIVtEFSsFjmxI
OPn2NW+inDwXhJ4l9QR90hCEfNpu47aKkt6QSZksK9nZHewbZ1yRDCzQqq0aCxCi
Jqn7pAbm1GBFAWxvvcYMd8rkvOjx+dE2/lJO2RNfh5gzA64KvuEjbNnIGtycTTHY
Jo/AwwtnxG921nTv+WlttgLCC0a4aKOBPh6Inp+WEyJBT0f6xv63wnloLdfwjKlf
tp1YZwM27G8wgokhW9NTfMOg0gBKbziNqqk23znA9t0lt7NJ/tpjddfNlnDNTi+F
zcAiXB7LZtC/O2oVtOUzewPKFKQFGu7FUtafOFEvJtbBS1dUtvb0K2TqMsOfTT92
bMweM7a6QJsVRKC7wNMfi0Ev0drQQLUqdBW8F/ZEGDnvey2ndPi9qURgTyet+TFY
O2A+ayaue15yaJgwfAtGZz2ml0nB+SqJrTTYC2mPWyZQAPRr1LErhcbGqRFRYd+O
ZA9EFsyPjwN9JyuyzB3xjTRs+ZOg8RSP6/GBe+yQWB09v9h5MYUBTmuEw+bQDUuL
3SDwdQGIUYCjpn3xQqMjs32rhoawDKP0CzlzD4l8n9Z6CNxItfJ1Di5Q4QLXmu2L
xcH5E0eS+UOuOMK3Q0wtnM1fDcPL0SHrmPd9Yd1cwz/nhyEZo/zmVZXowKNKbNF1
je0mXkOOiJX7/vdCtf3xWabI6BudRsc50CqWgnjGEdDELiSZtgSF9IX8ocSKNuni
KDVr4XqMCJ0fXQW+DWhb5bibBU2DgPIVTeRyQWudMcIqcJN0knMhsT5ENh8gEMDJ
AarBwvIASIxa5eUaJiEshU20zDateVbVJDopg9B/Jv8/57TycHb1V5kKowcDLPL/
IDtRBUN8QAJjPVIwPCsyPWxI7MHh1NqS1A8p3cJ1H00e5nUMdpt9oNuUIzPvToIz
wJ6+OIgaebBJBzK4JP/0dY+VK7L/yuMh8x/Ngw6TGoSIVjLq/7FWZusLtVBtzm3P
MnDEy+4SsAiReajWP1NbB+/WntfWtdDGMdpEaORLcXIeykBK9kbdy+SjDEvYMhhg
3xc+s/1mlG7NCI7E3qVtC/Uxe9rHKY8WwI7oZsAI3Q7M2EbN8zdCaz0nOQU25rWt
Wk1dZILXLLOSOKGTqEHDlH95EfiQzKKnhbA1tC4pGN9eNwL4WoHhbiHyZ1kLwCjQ
EML8MUxLxjHCJNPdhaJ2vptyVoNTgvwVDXpc/nEwz4xl/oFa3LpZqT2yuoYiGzRf
ODgKQ6uDwv3L0zrb25F0ihL5rhUBu2OJGZsTJYvJtHHuyWbro7EIrWa+IN2BCfLM
P2rKo4MbxAE63mCWcSKtXwIGAEqFyeZDgNdZjUgtRUBgJTZz8qf6OUwkDlNl8VLQ
GzD7DKN1gMhC+NbEZIkDJ9eHJrNXQr+quYn8e3YVwikPyIZY3HIrSLZ8VthCAznl
RjWRpQD/j8WJfIAVuPhFE8ZHkRv/6QOJSHwLAaF6S29GBDKJ9TQ+j84VvTlNoN0+
YaK6HRKDxZnnVab85j+LQ9rfN9pWfaUOpkNeHHnnA3wakFYClbkklXi/Kw2DASmt
AOiFtrSsYGC+TNk2n7XcXmgpB0Osy+RIzsYtLQEUFEweDR5fT0BWKudK3Sccu/lR
JOP4p2vsq6Pt6G+fbsJOBXct+J+6qMZ0xecRN365OAG926gW0QXzQlArm8N3NdED
WuZ6tuFczRGi++iTwH0pQ3Kf7vjTluSotTzkuk33MLYiZNTdByd0icb711YKfMun
fJjdptKFqAi5MSzfhbITROFjYafNGMfEC/g99A2BKul5Si0bhjPXYpyHAP0Ek7eP
Bd22lIczo755s3pmDoJGFgNnoSY0khBoUlNPWOBT8SC0WFJNPrZJ6FQ2ay3lov8+
s2cZidsKXi7no4N2gVdPMP+neT/Ggh/7VhY1bcWBvFQrc7PU9DV9RjG1Jo20BUbf
s4mg/0PFqqMCy5PZjP8ViLTm/CTY5CitenrHaqwsAioKVyUMwLxMx0rTdC1e+qUy
o7U7oMmMjQS5RTaNcztGQ/H5+ARki3KqD5VGrOKk9zOMiynksi20wWUWbvsOmJ3m
Hdmt81KlBxdxr5erKwCWBMW6BPCpOlmt3fwNUeAjnqeZhI9bPkshkiCtz98B/m49
M8lwJUihttyMkIfhn0xsk3BwG742XS0XtRLB+T3hqwfjVdshCzGA/p5yogEw4IBy
KOFnCMI6HDOQfzl+Xcq3kH8CFQ6B+7/QVx1RsBF8QyKS0XjqCm/ksvlLa9ib81hs
VsN9+ZkeS7Ht78/b4fIOVo8cOLWhtPYC/L4Mb1HuUcLuHheAGy4ReJEHmqhtKwGG
Gs2ShXn5vB/W5f3MoW2bcEgEP6CZZVVt5MyTdaj9yPeG9lHzawdkMu5ePMEb2hOr
sD/N4lMdnyo9REO5XMqVsEUnVVjEQaaF5rU9RDQP7JmJkMLpt/oaJIvj0Jb/rqo5
z9U9HTxor84qq7h2ZRiygt910YkFixp8stzPSJ5+YSRED+AnHoM8OmUfh8KFU15+
XMBjdDNipJdaKSvgJsh2jTF1vDu0RAs091GdsnTgrZNRV3BjLM1UmjNf4NSi1Acb
udLfEy4t5Lfw1efobQZ2AyxTn9oWCH5jDQGbKA3LDCzH/OvPyJuNwUqFm+nw22Wp
ix+GmMg5MYOMF/vi++NYsWeeNJ2W/I4FLrK3ymjwVmxnN2Pdav0wjWgmEjYv87qx
bD9z/yNL5pHv4eKrV61UNzWn2K30Ta9QoHRllMqhmac5R7P2kgb1e6PVeoHaItdF
5hg2SqgVfbuOXzx960VXXGXYPvD2sJd8DjVHH5GEM6OepnB2R6dzRfuqRj8Xk+k/
IUfkolR8N6xSPsZMG+JhcPMwMGGX2YizMwxLg47A52BpxMkSI2bCM+S515U5Ci5E
c05eljGLejRZ4GTp0iutvNL3lIYe2CiXKuonoXI6Sc3pyVsMgzpACbIEMVDVfAu2
qij2zDs/HJeD8acPafnrKjPYUgx7xW7gqNk+y3lDxdPNsBrXofW5EkuVczWQJQ7E
dsbpS9D4j3/Wx4OwfcKWS63/lMwhDUqNP0Rjzl/70G8SD8RMD/AIH8yDAJX1VB66
S9oApVfFr8RqTVXkBQMqVBIfVSAOC9WK5D52eh649p2EEslSxXvixqOoTKoy46Sj
rykO3fKWw4Kh+36B6AToWVPSePkqFaHU5N+xCeVirfaGXGmSmZk0RIniMiTBDJqh
/OvfCJb3TUE70RhLcgRwbp/CMmeGPvGCEKZxvBc6mcBfA8hiqI85v/0Fqe/Djx4q
GhzTNeJQBoAzxNVU5YkG/bSKT6KydhVl2iYDWp1gPmfEvkwAG3nZJo7zFiXX3WZu
QEUQ09dPT6+Ua4NY+V8Ri+5TpCTgfuC7Rhd6/6oLQ6T7avLXrskBV1EH3WmLzKzx
r245rHB0AO0Cb8Sw/CKciEIjvBPp7Jk4sZ2Li/wArrPY1SNmle3MNl5/SgeoHWLK
c+mIASgRacwW+nCaNOYyqzlObrZM9OmCLK2jMqrdrOTQZqDvmKfIqna/QgQUBr+D
G9vJgJM7XxEqnSUuv2SE1+2f6VKmZLU0GOjl0Ku0AM4GZsTuVY17JenmLegV+xHx
jpOP2pWmXJoWBSiHVpfgzvokuhYOtAgQbPqmQ6FkySHCj7C4rL2/2E1Z+P74gSPV
USXMniMn6jYPQM9OipbDEaOalxL/M97sGv1RsEgvkOnEasdFqUnKGRSAuI1Mo+ZB
16DE2XlEwLqLPkOPjMI0uFvqwci92mCzF1odIoWCjPewfzOQ0SDe51CBZZZjx/Nw
SLiPwm0uwqT2H24XK8r3CqjzLO/BpX/J4CEotQhJ7vVkuXjgrpFCKkRJMjbW2iBL
mS6bvKVbTjId0k9qqRf+dwCpyqDSwD0Qmume4Ea6sq9lQX+GE18ZVHGWSQF5WyV+
Y21Bsdir3BNwI2sGRh6KPTu/nQMhP6HqZVPyTAfkFxw27TRFR00xKaEXhAnfmDRm
4F4/WDeuf+/Cj/7hbr24u1WIIVmRNhYadwTpqeE28v6fiUIaadOX6hweu+jrJgZl
22ibPA1qeitSEKoK2EjQY1H1kh0uM9SIwr38nx/8uGTmDGrbDK+IY5XR0X1Bnvxw
CPi/6FSIqYUjAngdY95xT4SEolA8A4bFz9jNgi4KN3vfaXEWRIa2TTHuWFlB+LUT
wl6sWHBuZSjCJM2Q0mqFD6A587N4YkCrmCVD/BvB/OuyHBXGlzLxB2zb7KWtHPdz
mVEI5TxCNAGGe5hu+kcjiDwILyuj5hPJ3+WYQqIb7QukYrAr2XOpVPh6uhzEnLi+
C/uwOehpOiWH45Cbp8hKzH2t0sPKH8u6TWHC4dcIvEF+XjylnbDz6HAyByTF8OJc
sXAiTI/saCznp6LvLFv4pEUPoADahDNbJ+CtAeKmOY64RZNhfWEUnryNzt6dnF9z
4crG0R/WNZX5bP3DNOou4H0UJaFZsel1eTm4UNkkM9fLVSL7D5chYuPICsRoy9VF
ZnYV3FMMNnp9F6V5YS8Y/mtj9mPK5R9qyqDgjykxvlf9ZMj52ECUeXFq0vtE8Wis
BAKuEmfHKkUD3xR4tcBuTpq2y0N0dOCtaBEudVd593xXd4OmihQPB04oIbWCCOnW
BvW6KSW6nZek1Whx1k46T7Prkd7VSJ7gJ57xt6fZZ94sAVhPYmMSR8xgLPAcrShe
YFxGZogEvd7bhbgzXLGhlA5S6zgYtcydnZIALVvG7uaGA2D5yF4HzrJkQW4vBmpe
z6NaJ0ROyNz1pBV+2VHuo3KmiWvEVNCG0KbctTbMqu/MQtE6BWTlQXqJ4zuMjr+0
QBGcdZTTihVdxKvhBqZF2kzd46BdeLx9gZ6FEViKoRVY5Cz23/71TO10e6+MODCi
FsUBfdpj7gNqJ9lBCVI6+BOuuiYUVQYiaFZxsLlvz7EgzWD28GoOdthCXb58/pPh
kVFy1vrwRBvsjxzrI9KO6pFPJ6ozZeGuDJ4wSiWYa7uwyXJqFq19Fidib+pOjAWY
nPUip4VucA6iVgKhvzxtwoNAhxaOUDJDPRM06ZcBtv9/BGWTC8pDl023oNd/pfCw
wP9Qf/zQcAmIwYJKyJJL6c8bkNmC7NWNQhL927V4pskrXfXzKp6Kan1FecB9xjQI
rLgiHdl1hnNHk/eo6LWKV1RJaJWgUNUuJ44DejF0blUXVvV8uizKWi/E202/jneF
QhNDFA1R1FSznZmIdRz8W48gfDQgshhVGTRqiwK++wXShnPM8o2AIM3L8g2QHiYf
sqHgydDjCZrg9e2wbIxFw9ARe0jC9xh8jU2u8KEB0KlghZS6ngBbv1h4JCHeyVrQ
TVxZgsIwy55HCtvzMa2cUEbImdZ2epVLufBp980+JgtclXS74kxCIOQDcFB1EeMn
3YLjYVx6TQfTASomO9mWl+3pHorXtlFG0R/W8d50niFoUqjiYvVHfG1W5iZhorhl
Jry8qyyzoQhM910SD5y301eh2eDTwjn/jhdGf5eQxgycgq7ry/FEuwgGhMT9niM+
cvKqpfvuN2VycQ+Q8gsgYDCWHYHlbVrvB0SmqghPLyl11p4D3UcmWn2yytvTVD5s
ZeXSPPb7sOs6PAWVHUJ+6cTvXRdHAXLMAJyPrs/HhCZmw9jpbOpCdtPSIpmOKRvB
KArbUVTNqRN8ZT3zAHFiYOXmYJ+s0pFsbpX7KT6t7sG3/BIKhCzgsmIcUYrmum1s
qMRYMzYyJgLH9tnjPTaIifNWJ56B5lAWWHuDevvqn8QI11oO7zG6pURgbRcuJ81n
veNykURb/8/acJWmAZKl+t5xGuAjsniw2cXsrpZEj8JL+SOxnAGjH67jaPV4cZO4
/X5WGMMcC5xaYu5YMbCV0UQswRXh6vxB3h3BtVRTr+Af54OUB8ZuKPjSdXlMtRrG
KA8iNyFtUjOijsq7XA/q5dLxiDVMmnWkLOC5vz86RVE3IZzh1V/FgtlDdjEi6NQ7
J4FWG6/AHuVQr6HIXNlXfEUvVtoHq5lRvUIVyZbvC4oUcL9HcLLX91dsbqCcI57Q
HCyWsErrGsSccwFBgMmazGdXIbwQX+N3Cx32OxORBtzWcK1SOEhJkk4D4YDXf5Qg
kYmi5h8ET8LZuC0up4QjQ93kAU+NYoD3C8eLOQcHGCK/yECZJAzHtB4E3JlR3L56
FIuXdYE9kuMTTZOS1TbeTJmr+X4X6UUFsdGp4+LP7/KjzUYMeN1oxYkn6vnNs7MR
wMhoLsknUIaZxsbpLVCCxUr5IMxI+UxkaBpC7qMUYhIuHV3vP5vY7yLXiLANtnMq
zxMW+KAxy20rkqDMrL/iAA6FxFAgEDHWn+qwR+yjtTlcKw+aMUmjtzBuD/8m2tIw
VMzW/ikxd4Wr0LmHwzOUFcBS6dbv31236FCe0pNFXYtiXMZd76Y2gsaaSVc9jmHA
76fPIWHr59/0gp5DNXH226Fbl5HeV7z4JZpav0JXLP+XKfwWBC8NF2aHlleTPjIG
/miNP5SxxdB5sibL0nhOdZEpaPthISmfKEOrJSj4rgooHec52c8MfqMZ8b7bzKsZ
ve9IJnzLiiWXbqfi6iC3FaH15MPqn5XL/VKAxbp1AfMRQF9NZLVW8nYL+j8vDmpf
NUUlzjecO5BwTsofq2MEecANtiF5zlavi456hqCNyTS1ZG1UjicpjSfN28c7OtQg
sJO79Bk8ZeNFjAYU67pNhIui/IwRU+c9s5eAX4zVZv3T3iIXOQiwfTt2oqTuJCxs
xeni3Zm4AQRC0BGDo1idqJ+mU3UtdQJ9Ev0zJJx17UAwLMeljcJAvjKG230fOnj2
3En3fe6OVi5U5drnxA01w0WrzKJbCggicCPVDyU9uT4RxGnZxnlpYr9YSKssvitf
enFcu8mCA6Wh4N8Yrv9Y+UgARW0lJpefXYREZ2tuACn7SCzO0azBbeP90jS3BIeo
UtYVSMbDZgPRKIZnpOnifEekfC3WcSZPrXiGROk+w3bQabsGmWO4Y9Lf4VRxUwF3
o24yk9CSngreUT8j27k0HKWAQv3QTgRyhAXgLxeMBqBAvcqbEkuA2gtcu3kKQZg+
y868ZJA/HJuhfkM6l9emcmXampYM4AMducdJ3xVFjEodxyD5zQBwfGTIC3peRYW+
qLZDzgi55/Ogzra+LM+o74lTfEQVBsBTo7A9s9XZOHEm/IjJ52LsHBNVXFoaK6KE
j7zCEYKAj+P6BsjcqVW303riklRjeV9rkfm12WgDEr5hvDIDylh/5LCnBKBMMDMT
AvBmQftliY/srK8vMpsg0Mjq4FN7taXCUE1d/2ThmcSKnAwIDFhne8ySrN7PQsI1
yfH73wAYIA9TinkiuvNjpjIPqG/CK5JZHCeQ3CbXkCJ1tnutUm9Z/L/Zn/7IHCWJ
OU6TtXJkBXImZjcxJKDCpCQl09oJHJi97z9PyLO5ZmSkFNM/q6FvzFXnwu7bqHC+
v2ilAWjHIfwFOavVSDgasd1Ul/Xi3isBUCEGQ4Fl8ZjPKPHSlvEnNzy1YTx6BbuD
5v86X67irm9PBaTkdjQ2/foHk7NH3UQL4QRIrKZW8JgYVAbL/GYBB1bnaLx3Wfnc
/tvzG+V3yjCnYCVK0t7MNRaWb5urRQG9vzqIjl5RvyN0lKjc8cqvAnW56MpwOqaM
7z7dZ2zUKBsP6t3vM9/PrHey4wwxg1ZAaAHAj280u/BBVfkeNUEyJD5XJLHY+41k
B+DOKnzjUjZRdmYwEl3G3x6NqsmEhLKTICIaPjCkXwX2b/dm5qTiRmjBipVw5NqP
FjPa6xruCzIL4n9glXJXxuo1xRoei5s9XVmithkMwxz0vnTU0BXsfpdZlOSBQRfj
r5Ha4yMDz9DuN4uqQZJ6lC06y38KMHBt9xdDlPYTK7bB32kpb5ITnMVFuuufPwZY
kTFXx5H0IatcM5hcmSkzih6jgMLOGlfhF+NAD/+rPdoba6tNDTpuYqtSezORVhjE
yKPnMDhY9ej58YTtu4v5/OscOJ0KUaJZhbXVy91JbzuYya6eK1v0LbbNaFXuE0CW
8JAhHDfX+igXzNRy3iUCJsrkhAlCMFlmCzdbn6oqtBECf1d5LdWoZ5XqxqBUA98S
zh5XLy/jert7buLoMR9WbZ0bwbZwj4tq4fS41n7LPdKYqPuQ28h/Tie2nUqpON7z
o9KQUHKZdmuk89rVnApRiAA1fW4qPGQGzrxsRhuTe3I45NcYbCsOMcZDL2oz228I
RBMD8v4DY9gQrANt/S1NpENJClPWQ/TKfVCdqKpm0W6otJc3XURRRRQsG5blVmWz
VblUvt0RbMdhGHUClr8+Lt5p4pDG0MK/37SoRQG4kF0igIXtKJ6SY3gUqudkN56b
b6WeAsssiA8cGF/KVUi9ZsPIfvPIs08ll9LOg/y9CWQh2xLX3dB5TxZhk0EdjtnW
a+RJ+Znqa6/BhQ55pseTUlUkmjCKO2oI5T3hueIL2qdjGe9eSSY3EsmIJhK159Pi
cP+q/gXzo1iRbWDR5Sdq53QwHjN870ta8tQyXGqsSLXIvxYbT1dZ73yZy9dcffNV
uZ5mFvQwP8Yap+Dltzg6zW6RZC1KnraTWzQnp7jY4pmYXktVRCT5JWUnDvrzYB6N
AVFhbNotxtActzd2Vu4cZmxWQzfKtK6JEoAyF5IZwP/cgil8kyRBgxigMN3c/Ivj
+9a8vwpViUoSqRNHsfcgAV0Pu/0U0UTpRkeGPFs7aSJo6gmnpb8yUmrdwmLS71i6
A4BoRcLPo8IpvE0OMdNWPJGGxzVopT48sdCw1Ut1Ui/POlJNYOeNPat+VlaQqwj8
tYKLmKk/c6/Puj2MdgNIiFoIxM1q3MbDnc7NPjcfmLITIRGj1SlIIr61T2yevojA
krppo9nMvvR5DZ67mBWN2x9GsMbuSl06ACHMRKg0t7d8XR+eUgqA9q+Aq5Ntd2I4
zyoLhwoiw8ORzEy0rbAPQ+YJIbHKTg7gXOUWD5+AdeMQIDLgcp/PdAQIt4XI8jzR
sOtugDY+FW5AtwXUvKhfuosPAAjKnhmWbfgUajO6K0BrTK7jFFy0IFyuuMU/fGGC
UO44hrNZk8B2+aBYorqdElUMVkatfZN+2tc15KN01GBOVdUo15iapWTEoPjqAGfF
uQmJknBpoNkjDHZWMIcoTOvFutMalsGTw1PW8HRYsBFv60hHuiq+Pw/8uGh24Y0k
UF7ZBCbKwAd5TyykhhFHHzQvDn0KOmJ0dNIHM0Zu2eetVUoepb0CPUSJ3g16CTnQ
heVk7C8NvdNedGkm6ioxjoag2LGf9nzfOT/vbXi67YgYCY858J+SfSR5kVtwaGrx
//ZYSmVGF54YelnerkLhR2nMlv5mJZdeFg79KtRmxOD3MFN5IxCoOU4qi4+o0aaa
VC3+Mn5RsTmdg7eZ8Yt0okK38bD8sQgdciZLUj8UuaMy71ShYgszMCkOuNROCEzQ
VRh+E3ANb9yvEBzvTCUXPA+OullkGz/aJd69LpaeE3yEPeHlBv/lAhIs32crJNB4
6jcN7sxK0uvSmN/TKAGiuUjDKCrC6zpwTVC/x4deUFQH2ZYzmM/k1zOcY55qHuZF
HqlbO6jrL+cmPn7t8j5cmcRH7eq4swNuUo+o3aOW0nNYfQrXrtb8xrNRf+PXcrq6
fmelk+Zunn4vx1qnqa0zXn2SsQU0b4GI4dOR52PoMktV9w6z6GjaQFkhnSxP/PNb
GGPU6CTkWToq7K0UaIiwIr7p0nUFlHp2V/C/JL/PSmNDXTeeLow+AJI7IkRHCEqT
TLvggD0QaGk0Ose+/iE2TTXcI42+wAF2Z5EgRHb4Y3njH4dEdqkxuO6E8ygzOv+F
GbXtpJosAHQQZnxjykHvXZe2DgqNcHR4KYCfWdy6gP2IST5C9Rqzwv+73RSBiEnH
WhGxlSik9JN7pF6VEwQR/u+G4EzA6GRuDgKASf7BeQ+pLmZhG+bKQ0pu2g52KwHo
sIEifbelVTFvk4m31h2dgDfVCILA011ZdyIFlEy073qSY2reGMx+DP4RN7O7XCxd
lSz2P0rfmwGwq7LeKJ5Un8YWUlbCaTuxL8vVCW1Vy7hsg3slDl/zQIo4e5zwc1ET
FtiUw06NXK3AePu4/t2VCXVIuMgsub1lhbVElR5nnC+Tdmr5zj6OZtX18aY1Iwlr
cUeeBQ8k6bJraJESx9jCPrftIM0yTtuxqFNqW8h0qGzVGogyxKp7JTHFPV34iSPz
IEDpy8VCQ8LyzKKmjBd1aaC8C0vHoEOqDy764EcTFUxJ6yDbh1k3E20skOAE/so2
la9yQzLMzBSLvkQcJq/+o8ylhZIqOLmDOJs6EnBCCPgTYiJTdWZqu+cXA3OLrQ71
0rcqGbHXhlOKXIK9KcacxBVa977bsaoNbdEphs87Hdt1za0RrxtMwCZBS2oGo9Ku
a4bnX0k8GuA29aRoeiVIZKIV0IeCPFOl3q24wVZoSZ6B9XWabv/J2m9tdLbqa+t5
9CnHpbmOyh2nCixENo4KjN0uKqx3zoHn3KVrLV3IZt5hNXX+gO94Omeskwa+348p
9E5cqq6UYWBCqcrbL3T7gpIQbuZEsW7M/4mGUaqhaeYLjOwOpYEHp0BrLj1oGZxS
08jFCJHnY2knE/MozTZUa3ccKRmLcQMrP9Q+dlTqVetr5LfNWunJyjwIECOC906U
RWtUfQsHgjS/5g98eV96P7kQ85MQ/ViPcqTsMFYTzGyXDbzVeoJzbWG/0ifVlVvA
vq9YdcTanWuNANNGImfXppQQOCrHj4t5QEioqhkpdw2eSbc43xxmzwKT5oSL7jkP
zRdImUnFyftwLnhSdw0GqYAyRw47Gx9XBU1930mBRcpb6WUzhNNyXbLAFppN8gOM
c4CGce6K0wxzjPwVPN6k/wOChWKT4nFkQDvdYRBnRb62qWzdjjaDfAo9abEFQMic
BQ1mLI/kYh2JgaCMBXiONCe8eT17rZFV378P5FqHjGjlY26u9SS93nBuqmJIHt1S
BNpKk+CkdrF9KbNXrisv2aUKRgrlsGwf7QDnGqKFWdPgG0eCajf/m7IE6vY+8GHV
4qAVE2aZ94juyY6MxRqT74qqTJVpC2g6137KaFaU6Q8T1JPjvlL00ES0YMo2026f
bNvF5EmwzDUhHSKuTXP0gEtK5zQ28FE+dzUOfnni7u/HdPdZGAnmQ+MNW2JgUXXr
8rO7EfLvmW1mOIuzbjvkB69s6NU221WEo0y4jXAwhZcMvJkvXD3/yDea9uoC3RhO
Zd7o0xS9xI1qXJZ9d667bozBurmo5+rTKc+iGQq2IVGbtk5Z8OvuTy2e9K+Au31n
42nQaJh7Z5Gaf3Gn59zqHcycALrWbjAGDwsoy5SZupq/Wa2IxtHPHk6kQYPUZGQ1
z9ldPX9oqJ21hpurK5A7L5FSvtI8iu4eSkkGg80pBp9GKdngPf2WHTNGaEaxIwxn
U/+vbh/OA1w9b7jN9jjlaBfovywzhWrtujY8Dj0tyjR2oug0PQWIOi8EhyFG0XVU
Dl5Y6/Fwr/ZVRriOM90niM23ejyyBq/tGJg/2GEVdErJJGgLAzoRW/v4p6RiXBcp
z/0PaCNEKd2PC+FPzECPY+okTB/hgIGyv3zCB22NGHd3R3fqUEDjOK2ktSaHc1u6
7U0hw8Z8Q/ocQyedScAoiIqh/yVHFdr/JmDtlzXXrOqygGSUz+hzSIMAYNRXy30F
HZT0TPF3Yv2a2S3JjQaZT9CL5s+hyz0nXAZIoamAOGGzw85m02pxWNQrRNggLLPh
1/IL4DrhbaEg9tin4ULbdLHaHhdrA/nCIvZtd7XQpYuudyTwijskdwQVZWCZGBjC
WFUxc4sERemGgSFdezGImh7PIbRcwXKrjkIIZu/dQ0ZuRzcCSX1LpiZ6caaGg5h5
L5DsAaRXTBxPJlfaVGH9MmHSdNXZ8bcLJ6OQ3bz+mWCYK79D7ceB2HL+8O1cCgdJ
X1Pl2aL754kMNM+qyJfEFbYX8q2OdVrKPQc+5D0fP41eAWobmV+9QsRwCxWxLnsP
blxRDPfWDgSJs+KMgWkKYGRD1o6k88PtKxOqknGPtlgMgSfwLniqKPlv1oD9MW3i
HQ+i9DknRcu3goyTK6Hrx9Aim7mJ53qpaxsrlnJqGgyauQrgdue/EBN3nwkpd4Hk
HB3tzBfJSxlwk3XmmgkxWbYmkCBug7/BfS+i7OSUWEb4jdsve5ZSmG3nCnF0cOdU
srQqWGXDHHukUEqJEXABmh2egBywLrx360qHfajmHyYW/+iGEcXsL/YOgZ0IUvyC
AQx4c5sCGlZmrvCbEPgJM1o3l8pdPuZXrS6bQlFGiai3a5uemI4nt8wkRIBk+Wha
c4e88qitPqtmwO7HbnioljkJNcGEqJiHqlvJYRVUVArfD2CM/dAFp4jn4izFgk3H
T/l6MCL34HIoOjDeSOz1UO4MlpJCAleSigc8fDGTzYg8VXBn2tS0H3naxCwDpg+m
4iYV9ZGONNp4I55kkBydOZi4t+MExyq57Ou3VAZX9N4adx0hk3unILn9H1V6sT38
UK/YEv2R76O1RDT23lF9FR5QDBSaFga/JZAqiYGbvSTjiXMHzS6cZM1TgijvOF28
zjZcnmX0QVfr1jPeUZ7YdXHQ6b0IG0yC3Kt2XeYrSR8n/n2ylSvykbUr0vBfSDhj
uf4nGMjZax02+xs6NpwdBAeYsyTlqHB+zCts84eDcNicNFALoGLlYoaKJyzdFLXN
++GW7HLbllEZgQ4ruHDOKlbez+ksiivsB3XtSQvSuJIhH5ESD18iPO1uMIwburya
DHi/MqjwzzlbwjXk0aMoJrqSGZZl44j1Gs2uXyTDcPZe1a2OKSpjvE5xAEKLbt6M
mzzA3EnFdl11l2rcNXNjlyVOtCsCJ7yLs4+05ie6fq5b5DiYoa8hxlNg+/v9U/uQ
W0lvBWRf9znEKEPiOZ2idXXKMNuDdnUQM+a6pHmPMowVT8KauNceHsnk/cJ79HQh
v3K/JhcH0HAonepeyo5v0rUCzaf6AjbEoGUuhbCCDkC5mYd+ZoE4HbyK4Z0pbp7q
FOsc5mGmJPT15IS+iWVoBceecobaOt+9yItuxpvUhXAM8sZrRXuEdaS3M0REMC5/
zY/CufIdyzAt20WXRgKq5JvqRvX0gpUnPJCMGEA/MvViuiiiUWNLI+ldv29uSoPB
HKrkbJUf9x86sK9WVwu/Pxvm/IM//nLuac0ZvYvf+WaYZwfD2Z7NNz7Fak+mpY1+
SwX5Mad/XdczOSV+P8kju3c1QKpBegbcKP0MfY6COYFD32l38riBPk2fXY6sA5tW
cQ5XL/uoX43bmC7RLezoLoZHr7CiONAXubkj9SQgd2D+FS7xL1mwTS4QVEA66obd
pa8hW8CDV3rkUS7IvU54TDAgjl8/TM2devIJ5CY20XQYQApoL5ODPA0y1FLh44Y5
Y0mBQYgtj6903FUJomM0mT5LyRaIiFm01KjOOMT6wkQ+R+GsOZY/5nh/p87uRL7d
BNAG7xcFXL1RvGWMeEQ79F+/nlSM5ZxTo2HgOb0BLyij+GcamW4TNYB837FA3j4g
dKzdOnczJBfcvK5HkmvrN3OnvXyg/dLGWLS40dqdlmDHYJd667lb9TiWGsSp8M6Y
xr9vaWLPB9rurB0PTDvNqwIlRF8MgUvveoM1STUv5Q9X1Ywt3TGmiOzAmYBek9uG
yWvBxbNKh1XZMH2cPZ6lPTaEmqOjXlNOh3E25OAbgJ14f8tgPzoEMLBBDhTyQjsB
NW5XjWhdiHQVmqQkJZAN8rq//fx7HLC5sl4c5pawqNvGNTHT6OyZw4TiZQXTYYdg
AkpDJhapy8xr6RlIiwuDpsC1HyzH1ccPrNewUfkkdgsg6js+W4JezKE/7OrrmKXj
lU/Cl9zIJUoyaGUvKJJ6wm7xwhUQmh6sYQocS+FO0QRN/UI5An7H4EQJ222HXmgi
/dadWgN5DnBMUIJhjK9lvdRddwloA0NcAmucj6VeOABDwkYRA/WsOd4YrdigAbKV
UnKdowLckd38JPFARCpYPEJBcI+03GyykKCTwjvB7AByOdzkRmMIry41mImQOmkZ
gSJtHsaLoi8IAaOKxSW/dWQQLNvKFbOYUufpidXTj/VXSFepkylKCcFTIK3iB8CR
aqG4xAULjRkdNY9Ts/EEGKJ48JPH//KFkTEs4t5M1gDB7Zs7vuENELC9nhc6l/Rk
0018KIdmItrz6l7Y0OHcVdPVK8rttNNiKCvLHlmjeoRMQ8hPziW0N+2Jo/Uwn3RK
lFDbme+CHljG8c0iwTYNjQ5oqCRjgiIfax7Ne+MrXhwxPQZNmEUuVo5yFZfM6zMv
YKNvim8ZDCEwImwuVqWlqKbc9tQve5wEWUF/GAHmUX63jpy/sLQboTbs1NJWh83c
qpGZl894YumEkXAjttaJ2zoSmqUejE7P5HVp620HhJQ5uNyndYfzd0ri5higJ5/j
sMtoUmX+AO0kU5MvidTaBJ2RMXGFCD9Va3IonDVVExGcCOwTOH726x73vVFg9UqN
TufeSzaJQeEFumKC68UQES16aNC9C90uZRyEYqnRBc6w/03sd8LGUqeLEZTrrllO
ioFVkjmPVvOPfL0AqquEDKTjLrbX5VyZkzPKHhfsnvDEA3FIT+csueekdy7mz9Yj
0GNjQaHDicRR2tMqOuzzo9gkWyFq7xesxo0jRq6wolNqBCX6oCUNCbPXbuQcFcvX
51IywHVXKPAmytbrDfkU5enkQlVr+mjmZxIZf+6UvlAC/5EhyVYmHfFe570B7Utz
k2MOz6/IzZTG8ktHwbdV4ZrvbbMmOwdUt1y2BusQrbm3f/91Kw0/i54IOQg2+QCg
wyPLdAqafzVTTOK77eamLy7HOX7S+XvHZVyfhpWflkcsNhKMDF2r9LuaNKz8VijZ
0UuomsoVG6t6tAiZVXeimKWVWrr8DdM7WYul/D4ik1LaraycduNr+an5+/KMZWfy
ooQmIXydQw6Bw1BylpqWAR/WTJIXjO9yr3jBFA1vPB53QaQT2/VVVIULAQAKSmmx
pZwYfAtc0dPIYYSir9EzrsP8aZMhUgTSDpe6r/jAbY/CYyeOJKPNUzPXuanmol0J
+02hM0nw2D+QYdYr9IxLhujE/+AJix3DrkwPm/08flNzpZ5If3H8rfTqMRO7B/p5
r3U6VXJbf9Ec9htiUamyZ4rCqZgT0KqyTwgfCGH1qBPDUc7X0ZWNucCwuZO2pJae
SRONart8K6UVUwJdLjIpz2tavkvZm05mW5ejaYLbHpEy1H7O1Zea44Sge48cYXSP
KmeO1372X7yJCs7Ry1QyHYxsFZb0dHXU6GRKpZTxTq2QqIwKyHvagBmdJCCdvc+L
Aup8a3KwxfPJiM6Ti1zgXa6aTKzVUvmNiAaSw7M6DTjWgAhRJs+u5DCucf/qxtxC
0oOAiiIDYPJX9UhogI6V3IiHunUbjuMnEz9DQM3EVqUOxIRBAONhUJ9tXehqkNcB
6A3OkvZfz61FGyR9Iy8HiqPefk/amfIpSdLPSEeBoPijO/GE97WF+Di5CghrID7D
6qkkw0XaqyBBXLOIEVLY0N9R4Wd6VGpsDcFturgRIWdCqonEKlAWytPVc6AQlnTT
0RgtMVD8n0ffknpJKXBNu/1e8/DpR85p020OnJa7aCgSCxqQ3L13Ze7pTaY4iQzq
u2o/9g0k5HZSgEFyfWrHcI7su9RX0oWzesAMOA9DTudUGM6fYtMVf2hTdU3sA4AJ
F4wprskABOkEvVwMZ/h0RiiYhTsExz2NPVYOloRnKj8pDshJu/e1ETLRa5O7fD9n
OiMyY3gc4anq9M1Bzl5vwlKQtFCS1Wl5uyUPAgZTt0lSQcqegxSMtAOGRnZxO6yt
KVQ1xgFwsQxnH0Pyf9Xa3xZKTMoBEak7g6zrjtVGyyiGZhW4pPPxM9zANbCWQDor
SW/xcf7Q8/RdOImnM2v7+wpbOeFL0yBBe4wB2TJ7ivWyUG95rn2HYwXVl1vZLBpn
PhFJPqBT8cHqpozLQk/BE+iLxb66aM41rOi6bu6shIQP1JJ+b/4HnYUkpEMKYFmF
nuvsVE9RG4fYQKY4vEQcd7G8Fxo1KyrMJ6NSMJCCgdxSMlp2pqGqCjCeDBvAt17n
1e2eSrvIRTtZlPtOB64eF/TTugdhfLTXYauKgz4C+5ebyQ88x6ow/ltdtVuUvL61
`protect END_PROTECTED
