`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9azYpEcKA17Hzil8RhClea2tgov8s63rFkCttV1GAAB2RRLO3jz/ZaYT8QZ/BYW
vw5+NqVzx7OaW1PqIWzo1jTLyFbwpVHgd72QaIOH/8rIiAFViL3FGO06rQ+zJ+WF
467Ldum1JFkp1LSbijj9+p4iQZLNSHFdi4KGm7Dx5zGd2n7Ozxv7Daojs8XYWfTe
rdPNanGbHBrgDbfAhRuIXVXGL7PhvsDiOXgLf4JPaHuHTxMeq3giooupWOabzirk
mokcOiuQRUok6aE6h1V17dhsb4ZXPKvQTTmWkZtdDBENZ68+Kl4t/mxiogeVNWPg
KGMiWB8PubuQTErez17WNfpAr5DWCX+XR7KQfR90mj+e8JKkbaH2CsS1GUKVtXjx
XJtLzWZqwqqjdq7ES26S0dl1iClkHLoY+9FbblWe1dyEuH3PtTAwOupnfuL4N9RY
`protect END_PROTECTED
