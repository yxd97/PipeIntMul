`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/IxRDrnXpPxWdENBiE5t4G8Kn7LVusqJ2Vx1Ba00UGJMFTKlarlszt781QbSEQBA
SGWmTmOy91bQwwgSJbizr9rVGY+e2sO21ob0Xa3KsIZ3hNrlEMwlecrwW3koAIDu
oa/6EVBW4R+efP9anu92jA7rJ+7DJ6szdtc6NhCaYaNiyis0jTEAc8N0kQQ9tRSV
Tk1hrTLda6d7ZP5WRbwvu/9zAVJhM9vi3L4NvUdJiESDJ8qjyyxxiIM/dWoKxtlr
EAPMBCosKo2qAI1XqX4dG0aCXkIdiRop3+wWAobP1lEz+XLS2K5Wt+5CGcLMnTaW
SdkYpBmZj22vxPOfRXMDgmZ0ul+ppCxAao30+JZFDkiq7ZhhUgTOEHaQHf0lZdfb
9wuAePoi8ZnG2rCxAY+WvNuzyit14jGaMvxeugHN85MdGrq7W/hHyKpfr5DrQ4kl
6+Id81+JFyO5hFEvXojPceUcwwzVitUW0oXizwMVhFS06LZ9dmp184xTXOzF9IEj
nM9X10+mWIVZp+BjiG8G/Ctv7G2VycedRNaQF1lZbMMrb9+Ny8nllryjr/TAGNj5
ruFv/nflzkM/mQLBhMKA+u/5mq6KRySArhgeSMgmXyUhaveBvh2VjE3GNTD41w4r
sOs0y7a/NS/ewYIl1w4VYX95z2U4aJjYDEu19lKZDxw/kQYtHk9y4yZzCwAE4QB8
W2SzysdxLx4CqsBS2wu0TAkQOBsy+btFtd0aMwFWtHyHTWorWwcjixuxxm1ipX6R
xyiVBJBSKuBeXnZU+hVQ8Haiyg/ptLjv3g8y+M+lDebSWQC2geYUMB7qBZJxECIv
mdTaBo0IvjgHtbpltIaZ0EtqmldRN7FOZ6NnDc1HzAV355lEKZykQRcbThW4c9vO
B1x/zOrJ7tv4XsH4VWiirdlXUv69driCF8HpB3bRZ3jWIKAnO09P3wUkE4ewfIR1
i9Z7JuhfrKhyYQEFgJEfFGAhMy7fWwUTIHudHvalHoUl6lyTZGOW0d2oThShgsPU
zou/VCAGKJs2XsSvI5UR0vyYposOJ3AMPsZNrWjsu7uAvah0ifMejvcPq+6n4CB1
rUcSv8RNjOCZjtad2S3+17KjolCC+iwYezVPCQGfEQThbqZOe9eNwuRvo/D4LKC+
EaQJge5R4/vNxgZXJTH3REz0Tz5lf+jdDe73s2LhDmmuSfwYFP0V9L5opSnuf97m
RfiL81faDrk5We34RlYbRH9MM/6DdHuDV5dh8qaU+OyiW8XEQG4sgmoZbrwek3uD
DfzDR85SsKKg0lp4db0ra0VIwMZkp0C7uyf1RMMJ6l55o5/KWDCERPttbGk5wT4u
VKuc2mjIcB//Mu1/UQyv7hoZX2Ly/a64QyyJlwCQE0t7gTfBzZE2uN9b5L0uamcH
0nhl8PY7AqOc+WiGdUmxxC664M02ghGtc9fYzLxqddVhWP0N2Hc0yGEPhLgNSbuB
KVQdxdFEstS89gFQnBf2jUN1KV5rKqyE7jcegQ24g+Ja828GLxdwyoyJQbFvxG6e
y+eZPFvLfz7SF2Wbxsnb926HylXUXdlLCThX07jTnjiNhbAtVwaMsQMU49fuC9vC
SOeBgeC2Drry8qV51a27REGUMh571iNjR3I1DtcIv8jpjaD8Xr5Lqr/zWvzsr1iF
vj8EFymQfVGulOU7RAJAnB7QOjKc41u1ldct9zRwwRPXiGQBUCkUyFYsor1TpLPZ
aoodt/gaH1Eovu6rDLyYeqlWXPVs+PpAsAGQqxiiIk2u+5dtkWFSBtRww4naojQe
eu+P/UOwzFOR1UlClbiEw3V0GsDWOqsjfbn1RjHVSKbEx5JLbhwgaye9elHUn4ky
yHAfl4cw16NfmqQlO0Tgn8ANWavP57MIZMk6GWYk22512EHZ96mHYCj68rBZZP5f
zhsE7HROQ1NwfiNu6p/Gzdr4QFhtZua8K1hv8Gx5769RQkfB/snvpFOva6f50Cp/
aepme5VcKPxhpredzX6SLIpv9cpD4amU03/yD3jj4Ymx74p61ppCBGATvq1Yo4t6
+QXISb/keNjy1KqctPMJAcjcPHWcf+JzmaaMDB69wmr7v7Wn5SLrA/PRkHjvxRco
LtjLB41v/ses3fTS0StC4ZCmPFaoQwSGCjLMcL6G4hD7ppx4w0YuMx2Vc5TkSz3s
Ieo53RL3DglMS3XaxF7m8G0+IztsWgAzdyMTBN+Z9cxG0CkcfLdJxT0SWlkQF4Jo
FQhVqV+eZL1Dz+DSPXCmDeDsq0Ft1M3PDOgC8PEQrNhX+JrDG/TNXnBKh+AIWqOW
AYqdH6smI5nb5dSHpJDPHQnabaKBk5ja3P87wkb1goML6aM27rm+dq0h9HVn2o6+
sR9tl8sFScPt4dwmyUwyLX/0WchlN1o6MXD+ObzKBbKiLqBf579VobVXEJcWYVKA
WH5LjSaq09mY0bZM9Jn6aHmqUlm/fkeFc2zjmitIZMu8o0OIV/WB1S54QQixwKZ+
N3IXbIE+a2oEd38F2ihOSdNuzBX/IpwYq46ScABQZGOSGsVO8MHU1eT7Ptv1UC60
iXJ5JqwdmOOuJ7kBgR0ojVobF+2gRe7EEd1dj/PMyGkS93VU3S9xyCHsPNFmFkDP
mUpIUphPqhFwfyi4DFlagmCKT20s8V6npgz82d0CSiXxPLieesC0vTngjOkjTpAN
+mdUDzSW/au5yt9JD7g9lULqMBjNcH5yeLkyYOgVwgiCXX4vewAuwy2L7n2v8f9U
GsOR3lQXE8xJFtmEUb6D7aotvlTrEGdWis9buwK05bjIMEJpOFWINB/zBE6ryrYf
y0p44lxXN2nDs8JQ1xnirkFHpJuHrabfXJg500xdUWFiKeNRSUiJwarh2F/kleOz
1aWOudfuPmIph+7L5lXvPNTCkRb8vK/VLKYSnGjJojYVES/qd7XJ5sRlTucj2SlE
1DNW3jcQuQg8BjcQaRwwgfjQh2VYztEQkbYO6MJW/GmBEzI7ug1bC8UokQNJvXx+
er2VH0L9EEp+RZrB6Wd3YQoddbDguQcHyn+LUv9UXPNq7VXyXc1lEvvwVved8t/e
1coQf4lzCo0q+pLRypAfbFDYqUj95y2dSqMBzOTZCYuigYSGbWdm/+v4Tl9nah8o
kTajQrImqtwE7egDTeAqDyEh1VyF3R/kk7UF7sSYN7P+31pBvV5ynEQZZPXp8t+R
NuxOu0JR5YnYAIbiugkIXyes02OQPTyttuuGogNBqJ03F1ukWednqakbB4QKXQqW
f9NcxncV4oR7Pa6jg8SX6XHcB35HKv5pdGCkSW56Ih4YICpOPI/5ACj1SZxXaKO5
hdhlakxNbtMl5ZxTgRVcKkso11y5SqrcPgPLbt7GJgxWwY60q149QVFDHEHSHobj
9tL/4i8DGGhVdMI9v30wbaJwsgG/bWZ+tHa6WkRe2pG1xLhYUT7ij3n6rqipxePK
3FXSPhRKfm7cNWg8bfgMTzE7dLu3qbOlM+tRpL7P9v+4yAIBSljuvQiB3jdUh3dz
nNG2s+xrCzzgJAfhLrsrBHvM5mHzVYnekq/xWD2upbPh8KzrAaF+SOGMIqWhM2Oj
NKvD8IFBvNgUBaBkUFFARheAmNPQWoKNKM3+mLbk5uXWiyzBseuquE3eeont77GC
TVK/y/uJ9bBy3GMr7I2WOL0cqsbJZaVrTB71Z0+UhxKtqO/VuJHuHkWEZHjoFOrj
texK+qPxie+6DGX35ojWmuwfgIOAC19K+tzz+Fru025djAWAH5/WsK3CeB+0v3tr
yrWlwK8s45av+y/fKk5HqIPijdUo/eqPltI0afBWhKTQtGa+j7V6Zo5OHc97LytX
QFlW7g69ub0IfZqfDp/3p6Y6qoEt49xYvTsshnG/p0fVrfmDH2uAds/gQbkilxd8
4N5wLmmyAyKJx7Y0SZ2C0w68qL+JbzXaHZ5YhCbnLsZL4l2Bv7bbqv10Xq2HJSFd
2wQQuM7319iGO4B2B7couFMyq0pVG0+HctNRwoWWpfro40xvV+FjGI+4N31ndiaW
s/A3ijsNvYV3sp1NkxS0QLeNI7wmMpxQ9eVHJB1ETGE898IO6DD+iqrPIIOlTcBM
4ZBAdVFLZmfbmPtkazLajaR0kdFyDdF80LSzcG1k5SE+xKjLT+t+CgofDrguoOfD
07jIX8R8cDxU338KK+IQE82XuWZvBCookUVdDJfVnIcv+6ZDbsjdTXTRNTI6ja3V
MRtGAuZrXXnnwQ7U/XOpWibqKVXSKFwyhZz8LhuHn/HzzNzZ3pKnnG/z4uFA6WYn
1zdpYu9iZgRl1/IpbD4SZomQnrpwvOyr6Ar6u05xHHTCyMcYNJzyMRbDQa81KD27
yQGpjhUUIxuzJYspj5O3sByoEBzPE+8uPeAnFCMvweGlOa2sTtQA4m6WPQbcY3oC
aP1UrPShcuM05fY43P6Qq+ctqSUrheybxfzm7vYFZOTHQNCndRPKnq6ms05/c61r
XqiYTun+7nHxqPYGqXZkfK0usxf19gXycDOkDkt+KtFHtGQhddzTUf43DvC4XeLY
yKho4kEqBO1IvQmr6xc/IlsRcJHiWnM5kUyPg8/MAT38rBoElp+t+qnwrJgvSegZ
7rJeA0gMqQBmFlQiA9A5RfFJ0VwFYDpw8xIBPE314ezVzB1Y2M9zAxHX1w38ZwvQ
Xr2dSnx3uOHJEcNyGZoiW+tyTcYWMorVluEuuCzaRr13ZTJA5NVuAPsy+aXug8XT
WKVYYKHiKlvQYtSFOeOdqwJK8EtDiOyoHJZfWOFWzOWHPgWxxu67mwhNkLiDmVBV
ur8zLMq2gPZhjugzE8AtLFd8Hbd+1w5hEHdJgAGIL6PClM/U9E68egdCa8Lf/c4/
96TQmyHgFsdzK4APNLg20eitplok24ueeborxY3yBrdunXP3sFN66cgl3fHEQ1+Q
eO012y7qaS1EJ3p2M0MYnGGPsNBJy1AhtfNtxySP2jAE6M8zSe9mbpxCq0h6x+Oj
T56kdRK3la5dLLtovSvBfgo+NAPoddDqls+xZINJQxi7DzB9FUvvNYtaAN8qsS17
PYv2XO6AY1N1TDUxA4owmFYpqXKsLLgu4sNdGGhayhMAMHAGPMhJlwB41aGqwPjo
hNtkNNZ3ausEZ7XoAelbbS7JbbfYuFL47cxCXhfU9IjpleFJz8PSE9c/O4V1reoX
k4f7Tz2CThloserzDt2OlKz5VhfNx/kGzU/MJrgeO9bTPTJ91DMSTpSujUEpBPJI
eL8jEUTnprFUYx1ozfSiDsx/qZ7nRvOQvSaRwl68bwSo4aDpVNNBwf3U6daLVe2h
y2kbMra0n3qfc6xqQ/gMhiNDf2M7xv+M78hS67sxzcA5/oCSS4yYvJ+dGfZyRtDh
RLhC599okUQCwro/ekDd1Nfd/x1fThsRb/UG1BMeZlhbIGUCwRc8K80a8uk0nGHh
n1MGxbfxVCnSvIHEFIGSWEMDerkXp0hr1Ggp3yc4vdiucVSQ5YvPSf0nVM1u9Rp6
WHbWZ+RjjFXGBXScRes+kWdhp5PPup7D4r9RWL4k89qfBCDwves1FawCbye662Th
7IFP1muvRCzBr/lGOPPIFEl8xEe1zBfbhhZwEEt3HBxTec4GnWWD/R74QIowzXfd
6wxNcDjFCE5g0pwkzCE5Npb/AmlKFSheZliFxduYhTqAqQKLA2woRQ5c32EGXn03
MjE29OZBrdokiF/bq1YreuLLndJBM6Xf+KvIP221KIg3qp2svdg5DiijmJfyf9Qi
lhpft10r+TN+FfgqchGT8XqR432yvJDRifiAauBxuhTU6A7WfnljpgLgCGFcAYbV
ZP60yC5OrIwh6EGjOhTr0Xy5h9d7Ti/8R0pQmQx4B+FOUt0EUbaQsKIesC5+m59f
o1bZ/1N+MtXWeEnBILDrgKxl22qOcPNnnxYpoXmxp998F4smiQ7gb5COutZaP7dj
e2C0N2daDgu4vjXK0E6P3aMHHAw1n4sMs3IQFS5e1eNFNxqHnMPObCvXLn20yNi8
C3C14ALTakJNrxXgux1k8NXQHeLih5InwMTuwe4LZeKLyWI3bgQv82DIZSKbeVnL
kfvVkIFrE4VQYlWPJz/NoDrq59DmOP2voV8ldzB9utWGLp6l5EfYadH9eS8Cq0Kh
SfxuxG1ernp1sWwqjAI2JTHGM3mEGGvdshjo8+XhIuhOLcY+OTNFMOBkzckqphG3
X8Qw72elXW+CraA5Po7jAAqsnjariwQ9a7BvDm5bzyQZMHoPrhQRXyrTjxZr8Ybl
J/+apTOEMZdqyW8Kzm/GQMNMT3I27v1CJ4I/jDafoF/ifw8skT1RPrCt/Vpg3VQa
brgf4LLQ5ZxBz1rnv2i1P540tVKE8RLDBxSoUhMu3oR2c29E25jgoDqPB9e6f8E3
H4pha/9RsOVa5P0PmtLEBpopPSb07S6ON8pSlYJ8bevUVHWGxixXGutoiemHLuae
HPfvpzDPob45GI55buvkaZ+As2uKFJ9Hbt/3zGQAjVXXxg5RRVHy7g2qJsXW3SFb
x/JUAVBHVaLN+UzVib0o6relUBVqSOVSG5LwjfgLLkU2KwC/MB+tTVwpilOVuInI
eEMh+qE+Fq5V4lsWVcoyjS0PL5fkcau0ee18E7l0p4N5xYxn3BiaqPb5Cr5P/aV2
/A1B6n+kyYr14OYEp4W0oKuth3oTfK28wxk40HFhj57rJfKB3qRbREQhsxereMn5
VPa5rGoz3Bm1aQUyndlEjxvLDnym6TJt8+fYr9j8BgonTDYDjpjijAYvCRiOSLjN
BLYRsFLa89ida/0GiByCRFiBqvyrA85uomhTObWQCUU12Xf2qX4AASOTS3VDiXma
HnIeT6y37ycwjzTPTe1WKbd1RnGUnDE2BJdXDYtBbX9VfVZA1DVGkMCQkj4138oY
sfO2TgUHgV8PsbFEtGYd5A3n9VUG6CWIoSW12WY0GDbHV7t6DNnuhzUxw2MsvPjc
FNHNnKQX9KAYpdeIZJ7l13V4sagCoCI/qdTsyMIAa/itxcy3GZ3tq7DHlFn1yBwM
SJi9J9WYVO6Ly/bOj5U4o1U7IsJrfdVzk5vXSotKTLKM5oL3bcVyrIbSD01dkYfl
4OI62iQOuKO6pSvainPth+m5v4hahx60rkNQCSyCNqgdJyEzpNM5gTs6r8nbgpH1
sUn/co3VPvtyU8h5RPSbF5v31shHCEnmSGG7uf7MbZwJOGhqg7cp7uNtuwDUPATD
U0Yr5ZnGc1K2h+BrGhTqAVaFZAgRchMlXfS47knJrOFhqc3t/51pHgJdN1vlqAf3
plojZNByGqUtuSXAF6T96/pJfqiqIkWRkR+8Wk7GYGMJ82iVp7PJhvD7k8uvnQub
ik2nHMVF9c5DB3ps0F/Bm0mui0Gcu04l+oWNa6inEB/FqSQd6ezDNpkdzRwEf/5m
gzcHevL12sYTWMXT62MxRMvh8stPd8zUp/ThlimrrKjFKH72Ly0pOKc/DOSgWQRw
MlfSUR+gNhs7Xyx/+UxQnn6YD8wyuLNTmlJWqADPhiVj8ekoOa/daKc3bnQDucof
Xn9ddovi2R9a+k0qsiC7ZZa7oP8Hj6bSU/uCL3LDMHn/CU5tuF3KJxbnQV2QKzoO
BWhO9WLA1dip5yZQVitsnH4IHb1rEOVvT/x41vDJ1heudthxmuXIHqP+wuHZTFYX
4TJx999rC/qnTBUO1DhxSAYmW3b4jV+Bx7BoWGL4yaCUPeaksXDG4vjfCz+eMado
C9xJVXph98fqBSN9Cfqf9PH+861z5T69BB2EJCwVQmDD/lfOD/ZcqhUX5A8pS1TG
8hVpGVlRQz9sGV/Vw7c5WNTlC8+LBsesvZ0AX9q1B37LKcMKSNwITF+720B1s5aJ
TAEQPyvd+C3fNjOelLOm32hbj7qP1EqU6v2uwuQwO5+rGXEFuvnJzgbxKeJE5Rfg
JqF97VrMw4OZQVw1sIqTEZAo/2FoiAsHYPrU9gOnpzpPDRL+melc0Pv1SUTQsfbg
k8GGWJw7wgIc0odQUImZ3dixk91WQbaeObZikLvnqnpYYr6oj485U79aYJ+N0HCy
gVE0GZGvwZ6o+dwfHvstvmDpG4dNa7Fhj/oePNT4KLiRjOHlJyuAAKdnbc4mQ207
nQw6Q/4SiNFr4gwb+/j6BaAf/yyjHYrguI+h9RDKUjG+PjgeiPn0zidgc90JTH9O
DJ0zImINvE/t9ODSe133O3zuax/alXGS8/5yU0xChALYaj3bh7KOH5+DkLJ2g1ki
h8LtmyjRI1HwC4FIDtGhuOEYPqZuRz4LLxS75twaXQ4XPI0kA7NfKblp8VorUqt3
U/29sHJMmZA7LrHuQ27f3DYLzr0YeuDSbejISe9f8oE33SLCg2ylvTTgD8UbTxAR
LpF7Q6ARTI2x8zPZiQN20YAlcV1jGBNN8cfKkAudaNm4aPOUWQWcAmwqx1Dy0frS
sRDRL9wExj5gUUKK8wBxn6ijBjg6JDc5kmuIyr2mjp0/ZUyPz8sIhyJsEEyroUkm
AV0IR2NKMqIuLJxg12l+Zth9WsjozzwsgkaK5eB52TVS/c7L62oALaD4aNqG6iG5
Ri8arH4JY9Wj/QIWQVj/ymDkSWmWG69y9hS/vGI5tgANi1JPm2XDUSN1L0WFFfPg
cc/DxohVe2xP7MpJmdzyAF2kPpJWETwXYrzTetwjdPjy+4NNmHtshALVvOOQCrxw
6/uKO/xkMoe1dMNjpoxgLH0byuGfJ3EuZDpJd7pMHPVJZ9gTW/3yfFm+DFZoN5+d
afZleqQeJ3Jz8Rw2QV9yMpcVyp3cTNVW/Y3oPLg/2TmrhIKZ13z7N530IM9A74Ce
4QC71V9v2Q8Ua4mYqMIU4Qtq79SAz6y2OmXc4QgNQts6diAfcS5o4WhIA367utUC
WKrCxscX8gqd3Kvje7VU5PAUVPHPqrhsY+XZW8G3um+ugw4NuXfGiel0Zm827KCQ
oCAWaQPv8Us5OtnhHBo73XuYJJYnllK0WZZEDWkJoUx/lyCjm8vubpcQnIeWDDeR
NsnbRWT9NtuIPecOHIf9Lr86Zlt9KO+Qmit1MFc1Z4gjp3yH251Zn+lEtRqdLoDz
k7tA9dZfqRtB24OTfuNfgp3suBbEcxGXAY27+/9VzPg/dGL4u8slzTSdFa6BsHrF
QvGafy92BcaoQiAJl6Uje34vI1nJPLA82tP9VYzqs26jGXycwWVcfZxcO44ut66D
d3HVZjht6sX0U+CA6To8/JbbHqJnCacL3YTMLuDv3Htw6ZiQV2j7DorW3+na70n5
BTch9r1/4CoEUQZPQ5vOnA8OjRWluwI9JIeANqw6ybCzIFlq2hULuWi+az/59fAG
8fw5klL9T6L0Up4mVzGmAEJ2EDgiA5ISkIpD/BWle4XOszcOaDvyVoDM+6sthn6q
FAVt00eCRncYJ9pQhS5QSM7uT6B/yd8TNHygaJWBL65Aq9uxOWx57zpwqGI/ywO5
Q5e6kIwWDPEnkLkMsgW29nEXB5wKnNsa5jHYvErAmeTaRwcb0wNRV9+6jew6XjpZ
GsUwG2SSYvOEhhDmKfBX+PCMDlkl6lcTLjhL8qBAqZMAb+UnI/evkzyzZALV+Rbs
ENnKTo6/1GTmIiIDVJok5xKPSfNRAKwlQnbnq8WVFnsP2WK92Y2FKsyTcwUhdKff
qexudr47miGidLvvsSR2QYv70b/AGeiQaFGFZO6Knb4xCmutrL3hfZ7CaZeRm/65
0ohI2cGmnW8qXw81UydrboSXdKO9oNrr1xzf8r9wSY/FmbwJdDaqzbbTDd8zPPnu
tI911snu3/MOzdSj7J14xCYWjmvCLO7IcgIPgJMJnMoVc0Wwmq+pW9SGKdKLUXAO
WPCsusqYtFUl9qs3agNk7YYxLM3cHKD+WDgyORYi1kyCPvhlQwAa+W4FyPwVlRp2
zCTMIVL8zF1Z3CK3FXnmAmCjChEdGpVe5qj3eZ+dPlRQ3b7gxseOqUepx+CvIACh
5Bv4VBMdjqoR7rPqVAWwvqvoqjO1V4TyrNWGHYs1itEDrLwu+rkts0PtvPGpvEaj
5hl2/i2kkQR2b8BYXgZskoO8vXm3GAJW6LTA3F1m2eXm8PKAdr4g/kJH8ltoj3x2
ZsiSdlVF6RZIkc8X+2PeC38lQddj4DFEGWL3UmRuBK2w3CrbcUa9i8fC9uIwvj+c
//qNaIe4Wok55ytisMk7mms/mwJL36a9JlDlJrmtZYqOMeIDMXmeeoMBOhivTSgD
/FOiaBpab5bRiLeB6Taba7jD+9Pp6cHynXJh+er1qyj/58WQKRXqRAQbDSV41O2M
5nb6AtHLAHHpygSxrDvpvCNjT9/mL+gU4N9N+hYRiPnyXJqjlOJLjdLgvrd4ZNNI
9CG1OBWYWWXbzx4WXenxMZ4dvwdkp/csc40ngUEtzUiL1gyED6gE21U8G+/MnJkw
LcyQv4mU5t0TGV/xdgj1RvpYtGKgd0/7u9wPZTzoMoj5loCGCkUEnvOdVEFUl6mL
PSfI9S3H/kLVDoUZXdYEYCqyao8tOiL+4+XdK+lHOrYl0+ewTzlHZJqrMlBOdf7A
zxoZSpk4ZldV4w9xrcS1GbU1qlm5ZEPsY8EwOp1TVJEIeHNu+mhvOM88Sv3XvZ8L
j2nW/HVhFOuqV444MmDVPWDM5xQwMBihvirhfVPCSqbazTurYXS/u7SklhnuE9mC
s69eBVSw7jL+iu4Ch4p0GXjtNr8+z5L65iUCT/T6jikpyv7LA4U0270E3Wco0veo
rPK/2PUCfSbirqwNHTdNlTa6RgfAHaAzAob2vq+4GSOC7VPpHX0XK1dm9H9vi/KO
n40Gi2gmMs20naobNy5dl0jgul9k+53GnDZKbPtDdMKLnWN9WdBK6EKz2PofnG3o
ayP6i5RlYi/7SkcTrX1Z0+GmjQkYbZodggVocbu0jUSmdeetQOWJrRB3in9Dd6Tk
4HWywmik8vtK4nGDKcc17LMFAugpsFlWIeUorOPxrXaPNUOMOxmfKYPh+6VcrU+p
i72NhhjlSVSA5atNnpTG/xmRtyYVMF4flA9H9f4ZLttKAtO0uAZY86EM72URh/mC
ML0v71R6Atz+RQ0Kfv8UtE6pKhJzJ5dWa8WsjIj0IcROE2t0Z/wFfHEA0Yn/PxEv
Qe8gwxvCTmBUDQi1IGxrbYTM8ArIt52bHVk8L7gziARo9ImsaPDiEazDBNdwR3/j
Ocian9hNoHnpZWMlK6EFp4Sl3kl4wuav9wTcKyW35dQPWguA3NGsCgt4iKedJOWr
nFGK5QiRAfub0t7d6NnnJDKLYvqm4BSKYRuy84Sd/yg4092EwV642eZzo2U/Wfw4
lsDZqNJ6ngKDfTVUqrYHm3vZWlszo+uQoNALGnTrXIt7kjUKKQUpwSGgyKT3BCuv
e2C/vqew9VzJo5rN0tQVEsHDVAw1ooJhXYJ7ODykSx+aRLLNkYYS7FopF38SIIhn
+5OPb/eCGpHGqHVEwM6Ev816MbiPD3NB6d9+CpZOtPpz7YdkA92QYLm3QfhwUaLw
ecFpYDDG53y1V4ZwxUJuoShSkTe9XYKONgHgS6VY3xN6Jd4ZPuP//47QrVKCpzX+
Gqe0JeMGglgVix+zK5w8eLzKvmT01gm3eZ5Z4zLyJMjPr4wqROx7djVNyRBe2MHh
nlR4+HtReuvLvTmipdIN3VgsxetGYGENnpCBOgDlnH4bVz9+XHi1nETb7mRdJ6IL
SnKVKu+tR0v0EFxSwkI51hjkF/hYU+dMElbG1j4SQFWTFlOtEvJ4DtNLhGWjAzdq
JsaTvjfRn+UezKjazF/xTrD4w6FtDD0W7LKwh3Ebk3S8BAWyn/Uk+3r7ZalMjAFH
PeOOOOacnaQ3x9kpwBVxVSMHUMOUH9tc4RnQg3Gpo0hzd4bxNvZHxRCNXu5lKga+
KBsF73cXAgvIs8feoZQzuZjeT33rEiTYcdDQmxPyJ/dkY5OKjZ6LkldGDcTSLzYZ
LY1/fwX7bVQf/5SMe5dmgtDx5PPPYImTXJSPlIFzTkpPDBNFR2zhqUuJEJ5uCKa6
ArGV+IbUW/euQ40lT3XoLSaN0CT62oTQnSyHbsqhWcZvbWUZTnuxK0tXb0Hy25Za
iYPQgrOeg+JStbknqJu623clceoOeWvqLXuqryKww+gapWRZ9O/UjIW6Qkempr/J
rgXjvY0yLKnAj5/T1T5oHhDAgeg7wfiYpWUU9XMj1osngvZ7FD4s+CnEvmGZ0OxY
YtSfmurG0QNH9day2zI5aKnfRN3jAvCwk5yv+wkyWyNJgtYb1jrwW92gzy9PIX7F
ntui6kVjR/xUQf4u4ol1nfOb3evH4ulyXUFBZXgOWI4MukgWON/KiEyxVZ6W4sjB
KBMe2F9bu9rVmHJX7S/BCVUe4XakX9LCsqlzEpxM0PYo4Vcd7Vvpv/hH2ln58iVd
9lJHJxptfyz1SnTVMmVx96x2tMPskkOVWy1QZcR+Hoeex1bjb1RSkgb2EnXP7JGl
v26GKSTJvQ01gnRIEJyWTR7Qr2WViEbLesCqK5L89oxHwOP6z5bcEr+R04Ih5tkm
j41UyGfQ/i+Pwo2PMjZWRda97Vo5hDufJrJZ8O7ZLv9BuAaB2pAB5oivXqcZhRhu
Y19x2avZY6qrn/sJ8PUUjBMMpgIGZ32AORCDwGHWhkP8gsZoMWEGC9XQC76OS0OH
SYlf2qymvzyV7xklbq/7QMAzC1VgCEn0Elo5PKQmVI+2zRCJi4o9PBg4BF0rZG3+
doV03Ogv4dDl60A3pdFZLQsteWuzg0mI28nAgFqOQihfFgMcib9sIiUowypedV/k
3HZQOOz9LuzgaHb/GeRJS/Ztkcg74sCY6qqC4eVYZOwQt+CCZBSYvZyYUwKWs6C4
IdZH2lK7alS8jOVU2YG0Q7WqoPOU/zWBXvOrJJJQ56bDJeD2VyAgX1SJBsCl4U+a
xAMsy5A9KiUXMm4cbl9XIjoPzfs7g1M8hMDHFV4/FlPNl/5+kX3qSa1HUV8P+Js8
3HL9yyeI0TFL1eZRdlzfcBLBmz2K/4BAYGo/U3/0foVbachADR2Lk4T72PoayMWr
AtY0Af5bIkSfnkvBaj1HvrGCkDMVOo/yvQ8TaYbOv317N8kCeF72PUN3osJGsQTT
5rFcKxd/X7cMEBO1xYGFmbjU3gCmQ2Ax/cJkVB6Rm5HY5yC7OhFcfQd5mgeW8QT9
inPDbxaSRxo5bw512CqiXgZX8R/a1LXpIxie/rzoo5+QUnVqkg68Ags53dqfwZVs
6snBjk40iUP8uNDxAFHsjgjNk11qRAoz+ho+Ifk94KbYFAd2U+dkJdGqiatbvhFX
XwN8MeIricT9CcGD7PHwC0HhrnYZ5HpSIsKkF6iJZ5TmTFPnkNyLIg9QpxRv8QeD
7k7DqWNAu5miGdNBza8Wk3sAHDjLM/ZrK2xn47dXrmq/9Feo2alp7awsEFpZuvDU
x1KNXyQdoDEVZbUkuZU/+st3Eg6qnezeNdD6alCkuVbZ+9BGvma0ze8PwRajzjSb
1ujVecuoYCX7RuJefD3mm8Uodh3zfR+zjgBpWCMgQjOSa2o8DgcYOz+SACQsFVn1
b+DKNRuBYD8E4PmHJu3+G9GFJNJIhtKjLCqiT0so/Df1JeB90jngrooFQ7qdZ12k
0JKX2hr2pCcs3TpqBJz6/j+cS/tQpBcqsXZmxP5lDNfDyi+0ztNJg/zZlNhLISTO
Nzfd1NK/yVXNk4cagl67bTTUe2EujZrtT8bcI6Jplta6sU5EYGB8wCNQwgjyZpOh
KMPmrgj6EOY6YZs3fU4uwX7jPEH3tuwBD3I1/wox/J2DyXuov24CMnYSHJnMTV5C
swBQHocNpivSPNuUXE12S4g5wua6t50YhCrLf/WqS6XApRKy00QjLcOHuJmJ/NBk
7diyCi4f1d3sZW4ehjwQwAyaBJi+ySYEAExDq03/ZJAuSfraKNyIOAJtc8KPfov1
yHtXf8+LugTbt9GCQpZw38PUcMLSXaMFHGiy3MBIdZK1X/DS4c/0GkX9NrUBYPIz
5GKcABPo1ehCKWkj+9It6gbQmztTK8CvCHDeQuwAs/AlLw6mCpkWduW1vuRCaV6X
dJhap5utCqYkUgyjyzf1Y65VrU1P3mm9+r5a4kr5SWBNsuSCx5BxQms7Ts1vfrem
hXKXGxckZaRKZd/9GJBPJA6Us3WkUjuanDF36cg7lkMcrhTzYtPjRoRcfljQ7Fj/
WFOdeOFHNAggCwb6EtCq++3KESOSnkxEnmV3bixOiYRByExW0Uw0DOo7UxtR/Yio
z4OyeQHQvfRNlvuwhudBH0x+yt2o0rUja405mlAuXvgJfRWgfWMYWE+YUo8RVPQm
8azWe1BpH7xoYJFU24QZyjPw7cg8AABo7uBV9BHHzDvZP6Q3U9LE+eCLS0t0fnNX
+VPDhRRIFOCblE4pHD8GurkvBwm+nSlWe1ySFxZn7rrIY2/tzfkQBC6yApXOUn37
3Zh5jaXRicl7hct0kztMPP+8wWrZvhC2br/FDaZK9U9G0t6eGYbU1tUB6uyGIET4
CC9m3sJbKRvFTnwKPnzpVOJRPo7L0rJbmtEimhFYcb3EHx/vXM9a80xQezI3uV4T
acfqZztwklpQ2oU/PUcgC+IcKyvi+UQVyLsAtBabj21vTMHviWfhEVRBbRZpq32E
fU8Sb1Z1qJ4qM37eZI7EL2qxc6ku54ldwkXrYWnmBVCIFLAlQI1AG8RfTBGfFZQi
qJNF3NgvOrgVPHneC5cEfdirJ4ETb19xkaggJy2tMsHtHNsZQSvCaHTQ1PMELV/N
IM27wbRep70xIpz+sYSzdMRgPAoiDjEWDivnKjLe2jWA+53I2oUtdG0SxPgWgPSz
tLV66CiYZuyfjuvyQ5V4Vm3gHrwwJ0CMdrB+27cabce7kuxyPlapt19SyUEZkHrb
GraEcrp6IDGWwGffgtq1q2FwAYJC/0lIcab5Ysk5qBaToW1kTbCCRzrgWmuZqJUR
dE5T+h0n0ndi2lSXiiqDkXegiZLbXNVd78nOlsoLjDoaZD1STP47WwShUiG5p72y
oiBVqsi5FlXprmNU4U9zNvzYpFSwRvcUaUm5IxNBuAYnRm/php/QRIOxzh34XY8r
XdcliRD5D2YZjVB79BX1Eli3VADeRfW3teds20jxUerz6+z526kttGKcCneDNR5Q
uCsuwXN8MF3jMZ/CHPb5EtybZIEEFj7gh0LEX9QaDkGTJGakX+Y2GH8oTo9vxZpn
aTKNVHTW1n/R/fdNJ8dHV+bQHQXRbNqJM2dtyKC6Guq9nGE4alwp4WdiA5dxUWPb
XAcbsk3PT7PIHDZSv6mQ64gfu1Fjs4lX1UUivXXyquO+GfdYv7u3WmMd++Rxp2lC
ov/n3yMTjj7lw2tDpE/Ksg2wiJfUOfuxVxVt5aK/B4WtCuPi5dpCzj5tqVlN+dUG
L2rL64RUJqoAj2vtHdF9mP3DoRau4LdJByRfS/QGunLJfVNrJ1OI1YoODtVFUWd1
uBKrd+PhufsvaqsoH6bBlxrZU944vwJ2saBz9nFROv6+Db6cvSTDhtm8UJGW8XFU
1kBUqvbhaX4lo1H20rGchAJnkhw7mUg6Kf5NsZmWe4mP/7/d5LLWPM0gR6Af/vzC
MjffFf4fZhswSbJXFeW2cwPwn56EfSEl8WHX0Dx+cGe+QITdhsQoG7pKkvB/eZqx
jF/V1Nv5pDqZDNG2nXGN2oj6OM9KjDTPkgXhL1/ZIKtl7ksFMPgssjJfigeFui1p
ZHMMZrMJwzp+4z8UZsOKxyrDmFj1LS6HYVDRTfCAFs6mZFpaZ5N25XLj2LRE/hgg
pxjmxvmKpTDzjtHgwieL3yjkJC/SGwsWTlBJkflgjAuhzsl+nDkb0JZIYkrb0btJ
m/3WJmlRyS6miI7uw6RpvcHGROZ/W/taLGTxu59SdRSV+JM3/DiMN6m4JNTOZ1v8
lIuRQhpg6tWQtT6MvjrpI2zEwe1zISIeUefdFqH+yrwsjPsKmg13TvUU6dR1ASzP
6MLw4jp0xMU6QHvrR86litDyaykZhG8SRagBQxyVIiZhvaa+D6KJwMPJdRk4cYV6
d2LA95hQiAZkmh/gj79LbOtBtxERGmC1XCnckg24jrXVdIZ2BRFNIesEWhEthtUP
5ZyWT45giONU1qWKtC5OxI0d8bFAjVQsuEuw2caTXS6yvUTAd1x3rekAgPSsFJx8
F9WIbdtlBGpqiNSR5gdiDIfYWg1wwG5hMl5tG/EKSS5kGJ0Z6VZSfk2STncEzX2w
qusuhLJ8xnpxnPUaVLSRSRV+U5MblbhJ5Y/caJYCt5EdBBfxd/9aKdp/Pjer6NRP
zY+/tavt+vjxlm8tqhlEHOnpWl40wZpEYjE7xRIMAXVWDN0KJ/bOZ38eCjAmKvlH
PtzwQDE7W4AzmPeEdz2/jk4mkrrYQTyzLSZe+mkQW+uUt3MHd8+HLwfJioYtpSTU
j2XyuzO2GgoOi84ackiLRhLVuHnXBs2l4SWavNxvLXXpt032tJzshtj/JUQcQTKZ
gOvycv5rMgvLgN0WVEhY0Rfzy9USFdpHH9cHav2KFgqA7qqnnVOiifKMuDHF+uJE
rLWdjqYYKLuwl8t4VyBN/7MIPpKPUYmtmsRrEuT0X0lDMDD+iW7x/lj0RgrrxZJz
0n6z51akoQvyEqrJCLdtFaSZOe1BnwYG+nH6hg7Mnw3PL2UW9XdRODNv2WTxzdfN
TQq9WDU5bBXjyorHWIX9laVK+rfjyTzCj5WJxkUIu7+m9CLzS4pke4DBV+AxcWRS
VEx0zVqvPAu6VxPephi8XmxkRRSGSpRpW4Y0TXAhX/2wbs56CQx3EKz5cGbY3lKz
FJJ7BBox+2FIzbgYzyYrAK0RUveobIBXSfxmIGZ+VUJDvZzrKxXXw+eK8k3rjCf8
wXzf8EFNKKNy4twm3Rrpao18HGKtgSovIuMKZH4rgzYab+Ci5anZTbMWRspckG5d
tifjUhjsoIdl2p1lRV+WCJlvrAThJpEspKRM0qNk45ByQvc4g7h5JvT7ptpLZVNl
e4s+sMv/4MajJr4KVXL8jTrb2lbjkaOLVHKTg700MJClyswEBoeD8MRsSJhCSunp
2C7PuAwE9bbxPV2LC8LngiLTeZrTU7SO2qdHyRMvC8kL6X/RT1vk/0i/0x1KjgDF
p+f6Dtf7YGhMypMpBvGJMiYAtPqRYOcCqxgyd7nzfOTbIUbl4rSXCo9XHQ/cXuHi
G48NaNMAWhJfoYk4lpIAZW/3jwlt9x6eod0iLn5QId8bZfJxn+v5t3eX1J9fJfw7
i6j2WECWVfbJbNE4CLoGy5LqQ3z+BWkPd1Ab7Isa1ZJCsXeD6jXw4dndRHrnfC/v
HOl1g+h2wvvQHn0Zpl1V7l4S7kw5Z+3/dl3Zt0N9LvELpEQoTAp4Pvotw+cVTbPl
aqfmcvVT8Vc7Jv1Zo0WgGSNQpMgdrO1sXS/1oIFnsTbDXjHW9URDLC8xXAtTQAvG
OfNmtr8WPlnKvYHVkvevZ3d8oQO4ooRgcyeP3LbUVOvIO3Wr8bGTETOW8YZpa3dt
t61fkmFhf6JzlD/SqLrQofMqugWGUH/wrv7pFTseld2vmgapGRA1ZYkXBFbUYmm1
BToVpXVIE32G95laMQ+9MJlDEzXWv9hdzipMEiZyQ4n1at+6gKMfDBoXva2lOjEa
Ao8KGOXeNcc/AST5Of0aXemrzPzLrTRliJo6JOYDe8doJcmqckYO0s+Vvt6yzR6P
nloHPJ/EgRI+uDYCAPAkjzK+b4aRHxu7NulRQ1fn29ndcUAyY8acj+QCUeEM/Ln9
iUiaAJu0AvvK3WwueE+jfvxTDXQN8Mdz2KHl4gwGEoY8sEGUlZ2CTZ1w9Gb5T4ER
i1RWQBmVLreFO3V0hxt8MD3u+1TpBr0/bkSAJNQiPBGPqJr/yRJXFj7kq17Enhlh
3yLgYRwB5EW8Mod1pN/rin1bE+06f5g2wEzPJV09LF6Uy35rqgX3j6PZpYIlsWKX
QkarQhQmXAQHGtNI5Y5nNn0Dmbb3PzuxtROJ50yZl5jZ11HPTz4Ls1/S/YdVXNWG
GccCMBMaGdRVbF4IPvI2R2Otk/w7kBM8AEf5t1C8mZVRj1nBGRQbkVyTRe0qcY3I
bzn5wjJFh5ZFhkjjz5+n7zAeHaW/xgIVYb3SdX+RgI4EwcVCmWnVt48RLa+LU1EN
Q91yuF0sKdDFI2y7K5Ok17savkUqo3dtTR9o1leN81gIktZskMtyiIHX+yrkCAnv
Ndtyx3ZZ8IuYHy3TZPK9oyj51GP3qhV6hCkg+KwzQeS1Buk8hfonYGXmTrzOPP8/
gpbeVX0zIW+kS1vGvoK8tCqZwvwLwMJr5ic/ybIx5YS6GcdjtTHrXrphWJb6ynJX
9wk7BU0lc9+CSrH0+sbihiBAMskWNU+pq3Ho/eFJnMGzwNYocpQcxnDKSn0KJCAV
26SLx/nyrHHVnjvw3lMb0a07Czb5aijTi8N3mAxH6uRdpWISdBd2M+Op0nvdNUPg
bQbe4mghagkaSSnZ19mD6ZLrI9NWa1BBGqE1Q/FGUFosvEy34ZH+vNIdpi4aspw1
cTlEROMsQGRKaEZZVOjyXch4wX4h4r2H8kjR5TmukMJdv7+QqA7S8yr4HEm2BZhE
ffUkzeV8oGwtARp6ujrREm6mli+ObiDfGwxZKyQ1w33bRivCid0UKt2T5q2RmW1f
c46C8+qOewDD5Q9qwLU7D6y/7MNNgGIJoKpNQVPPCesiSpojHsdaHncp0rPnY9Rn
oo14AZBTGUuM6C7zNsRRWzs/wzYEzMLmaGtNqKthELExYR03D5pZq9zgTdAciJfT
j9fCJtBJFtlGd431qtQm/sU5bQoy/5vxtc8OElfO94wxsEz0JGmvnWd/gX7V8F9Y
yTTJzLQZrtyiTi7+XXoqfJQHBTBI2GckjqAVg68OMISLbIsPLAlIeupkbFxKRV/B
r2YqWlzhqoAKPrdlnPzuQMPUIb1DdNKG7+dZ8Hj/E0choDQZwolFZ7f4fDehjntJ
i3AGB3JVclodEdhyIrNrrKdzlcXxJn1NxgZz9g5eTqkvEQL9L+xKMa+Ua6wYI59d
8ttmEU80mXV+dtVl2/LDCwqvq+fNpLE3OR8f2tZ8LMp+AQmpXuumew0XDNpB3nod
G0O44wU9Cixt/sTueEMqo8VAYjnVNHHISkZw2U7Vj/jVVDX9Pw80v807yWRfiBHO
DEdINiRbxfmtZRvRDGNThxQIpzn9wfbrBze1XBXSPhbyeYxWNuRKwIdsQyGMBNhO
Nv7B0R3orWUCM66TOs2NT1nvSBL54XoQ9UvhBtGhnQCpuml0C4U9zHG0LDVZzA/y
K0ztJOCThGa/QF3gfRbv2+1SLtVHtcZ9brfGvO71jNVMl84qCTCHD/o96BlHS7Q2
S9O2WqANwGirKqqs99UHUjmusSZPpFLcXu3+52XKmYR75mUG4r9DRAaREjaQd272
DYrAoQe5Kbsrna9mIru+NKsGZGVLE9tSuAdWjXVi4zxNy5xt5t7fWnFjkqZtIAzW
PNQjN0DVVpvkQGfm4Xqs+uCVvhZnqbYJ3DCZs0N9AL3pMwO/aMI5cL6VmN0Yf/s/
hhwH+od2iGJqmJdyAr3Ieuazq1IHr4VYV09995kMxxYT2C+I33jXj9l9F4AlF/H6
JmYSMnHP1wj/heWQ78VingtHgox7GZ66q7DwqtAdg4vj5HBtPbwu1yEhi4UmNVZ4
QERgR56Yr4hp946pIVtLKRV4xmZ/47PAXsoLwqWTPqIMrqfFHqjcFO5f2EJ+sk5z
Ri6Im9FGSrry4uSWUoibYoiD4GxKZ+Umvk6868FMO4F5WfrKkmCpDTc9SdiRmn+f
48vNYUyAmtY0Axt6FDiloHexKYzLXg7EkcAVe4kyf+OPVvA1OZZeD33Du416oQ8d
/Z6WiqEfCV0YrC/FbTeYtffo5IHw0fzU543xWxUBTAVkdXr4LzwoQpTZDZ6/FGd5
lijfqR1LLs4vdRZ+mPjxhxAp8FnZuwWMhP9TbMNoIG0pMpIs3yOrUOKm/f2dyCAD
zTjDDKUVsYxWG8R9Ryk9Mcu1+WS6QMwE0gI4P2f1eee867AYDO4fv00CMWPJ1Wxb
uUAije1bf+CpFkViDJEu5cZaMCH1qTgfzDgwa8psAilLIhcCo7Y2wBL3cvjA8mmr
98d1s2D/slqibgU0kkXX1cDH4yeGlUj32nkdbKL/CQ67COnh6RPf4doCnz2lvhYO
MgE4ZfelfGc+qc0kGKlfNj7A9df7mKQxmiHPWYSeetVFuBCSahJz9WlLxmqAjqYT
wjtNhHm1NZBOdcyvSZM7TkB37lmn1OII49tNI8g3+H6nYefe1xpUPZ/R2rF19iyZ
xq22xuRhMFiOX7brtYqjs4Sv1gG06CSY8IkmcPfOOfcUlpe4bQ7PjJMNaVYmpCgA
4zqdF0R0OFvj7M4hYtru1MSibXnfsYW5KXaMkoRDcGc0aQMIp6YHcOgKopGnIzyz
xQpN2N7um4gh207HFlC01aNymY7ugDLOEWA0g7E9lKTTPSMj2OEZkWSg+DJTY7Lm
R4hZRbgUHfbBP1cWwXKK9PK29UgKmNhBVj5P/RNkxpWrxOFnLenLJHBKfWFaejkK
gs9+QHrKTaPIpJ9HPTb92DsOEN2LetcGZ3s6F9uz0pOdfCJe5jj2WnFBDMliQ/I5
i+oYTz3bUSwrnZV62Us0oyKmQuhX98OuzUGpD64VcpAW9MvnYfL1nSi5cdQ063RL
RPYp3Ng46Tq2VzzE2TyZLvNY6BPyUywKipeUkJ9Pv4abVenBMWkSheq1Te00azDF
Qyij6h5BWInM1NvfmuzPtVrPzeHF0xPq+L7ixc7+bCq29X7SlSH4tjckgdRTWf0Z
bfqbti4pEnA51jOGvUVRI4QsWsw9OvJjgluP3ZSA5R/lZHq0v+H+TznwxW1u5xWC
JPUcUUdEgTaf7SIym5ze8DgmxvlXMERaWRh+QOfvgwCC6cJnktDk/IZTS9rpSVit
2MMah7PLOJ4rVCZzSwi0Io14kcYFHV5OZ6qY3zO6vRGHKJ0NYrUWOpPbm6qgvQEA
UgclGQwyD6kgnB/2oJ214slhYzrOZU5PHC2tF+j6mLtZefHiX9lRpShacAW7iE1m
UQdtcgovvhawPxo9uhRm6Wl6ZxWF+puvCOR8ljPH/28qx8Po2MTR5EOz8bJW2Fsz
SRQSSTAKbiX97tQqItv1P58spFokI0sLJ70LKtj1IcBTvzSr76aqds/1IDmpSKRc
GCMYhUfa1GIXyHfUEcI6OhKAkPGu4ySDFMskellkjizD8+VomupZKJ5T+58y8gRd
MK1JJJUOa7hIWftvAHsYBiz15gdeS2p+bCq6HvByNDdj/8uM1IdSq2Hi87HHv7cC
wxiK2i2csVhlwIJd7sCaPcFtjlp0uQFfHnHsW6Vdm1RujxAd0pzRnhtiF2CN5VA7
JtSElocafSRNkV3XL2KexhXpnXtos0YD4EvG8w4yCDvpjDKPv8l9zLOqtS/Bi4Sd
sU7W/2CAV9lYgx/n3G0igA5be4Z4WUtHgTLYh+vv8XHfVNI4+g4BPu5AHQofYf+M
t0CADj5muf7nv2XJTI7TR6xLp91r2x5gMaFTbSPlJHck+Ml+Ewpx2OSKvTw0KHgk
VfrcFXBfXkFt7IGcm9U8tGqphQ/17iIOO4uVTf6oWpxVSE+V1PvfXlqW2u9xBW5b
68B3kn8YKE+pFWmU6TvRLfauB5bdoNtbe417G3gi+iAkK0oB01fH0CSZLYSD2ith
8DeezDAeqYueupB4Eh4n9YibYV6+tru1C2CVosqBhU3bd4MwSWvKJ7CDdZt03nHC
aAfhTQksPs0iq9IF7Boy00o/6/Ft+82gEpiRUSQjCngA0QZun+PuXKejS+zQjyNX
RouSfHQxJs4z0zfgzIwVR5GpVmTAMGHew4jPXB7TXbVeCgtx/s9WPak8zFGUV5SL
PtSEM9voAIfuV8zjiJZLu6QBeqjesm4yZx5ErB1W2B0C494T/NzooLxMw3zL6ntc
ZSRfP1su1qBokb7L9ho215TCowaRRhHkHXwPdBkH2XUmdq/QjleRSIDWgqgQWe0c
UvRLWkN7Lc4xVpIkYFmLDqntFIf8nQrG0pftDI2MB+WirXI8ayGcJmZ0H1Fbk9Xo
N78a2Q56dWP9ydnGbLTcf1tbpWE/ShiuZpNwWJyWLVkaeQVXxe/HP+pk+XJwpyoP
fsC0mReWmKtnTnc8Myn5mH2VIxC0nrWPdv1Epk2mgBTOibcdErAnvHSW7mnV5a7h
rkSEMPnSpr3s4UR9EykjRujreC3sH4i5W6AaK9qZYUpdqQhRh0hlBKq8fIW0E4M7
G/qaq2KNKB41D07gmMGJdd0RXSxWhd3OHALNFPohoPYKkrZUmXWs0y0C6kEQBe1i
ndQYvYntDc5qSkOKkkPZ0/zjvf3zEx8ypau4HZaPzQzHUH2YqDV8GQ/G9hQBW1ST
E/YlJh3/ZNsuD33FSpzdZOBptokBmRSUHtOO3H8aYIniQ8UV72rSQFk8RWR7pMa4
VT12EHK7bejtWDoUaUCukLCQBJiJm0+K9+n+XwZ8v4IcxNHc6Bpv0RVM8DPHk8go
IpUddHzhsdgB6wYYZmvfLRaKpgezm7OXq0UrMpzdnuLYijOEeMcHI9v2NjqY4sFG
bvPIOZekyuqrK3xCzaO/N3w3ltIkCfpbguk89xDZrujReRZhG+EOs1MUu2zZN0ub
+EwLBTwgxSQqRIp+y9+j7HaFCryb2KzRUSI9U91fnaQXi5SY40w/B88w+Sid9eTI
nhXtSmlAPilbrQGY5oCRklFTxkUAPfIMuVpyiXEia4ojmL6QhUSGDmTTnrEowXr4
VhTwknTwfqb/8UAiEG8PrPgaqW2UPYVNC3gp69f4KgHR9xWuv4/xBEpPx/+dyIJO
9UKKpwD9HE2g+BNkZhxMWq/+iGJMQFXv9zQXA8+WnBlaD7LborSLjfjKvBUnHuyc
Xc2tRghwcCC1PgAMvbGO5jqYYLL0cvsXf+1qfaIrcN2uvPHGBGpMu9dDM0SJA8Qt
SFimLsgNO83ZCEPyIX0t/h8zOTs/EbmfkUnZG7xPqKzI5kqwXf6XZi2Bb5zs8r+l
Q4HFHsPEWFSi+Shn3WVIpgvCs0jleRTRCoMZxLdS+Z2YARxao+0Pe6k8Uje6TXY7
NrU1OmQDciSzHNdVhiFsR4Sj9buKeODEg4RLcar3TZv6mzmVqbmGilOildVqRyxa
tvYA+LIKOZOtV+mAZw5dWRwbKrfClnya8uYiH9KyLfzqHXtHCgtIhtfpYnHfGq2d
6Iq3m+e41SO+yd+sqGoM3VOR+pfjAkuavta0BFu07X3Df5ou6vnL36BAqX+NzB99
ZYh+IEJkf46Vpyug+W7Bm6o2ohiCylvceIN7G6jR8C5UFsN1u5vCCS5PR2ccCjYi
860GW4ukfYCALjMr+2Fam19qRAvwGPrj/ARaBIqkKdh3enZcOSvblQ3Bw3+c7dhi
I6i/24Rluj+3VQjja3vhDvSbPMc7s0BlangclEhV6dbD9OPKr5V3Oao983XzoZx5
FA0AKqmGaRrosUw65uunpY5v1RRg0TGOzrfJ+Ox8JkokESRYp6K9AtV/Ij4jatZ4
dZjXXqs1/EpiUwGI7EClZ/Fngcgy7OpoByitZBXS2S67zVdLrAORFbzJR4vYOzno
Q1my6YFZu3fa7R4BS127KDPGhrjhQ75nrql8Gt/0Mwv6aMrLiu11Ozn0Gz8O+4rL
VwU3PzmxomyxrYCWnkcbuR4iwh8VzxWy6LsTqIZxzdM0A+8LD89gM7+F4nd/gsI2
JA/IflKHAWiuGGNYb5LObfhtKuElkwYqlta8ENO9mCmAinIt3y/a7A6dsmpcueKp
qjwYwKkSOKRxjcu9UxbJXR70nUzcSDVAD3NXN5WTuLMguU6Y3Z+hid3kf7J0h0YS
AF3LvvU/9Qi/wLsznPK/YmRoZS2mGKfoo+L5IsqwFEjjlf1OeTZFAuE1ph4iqWkc
z8fVkEvl5cTDs7zsRl8uHhwrkqZCIVdThnFiPyVzk/6PUatdSPypWsMtXe9zTfWT
DbpsKcQoQX09YLpHfEF7SydXzHqImA6TMTln8pT6QxSTci9w/Sf+7PNjBhTFNLxb
tat1gmt5PlB/kpKvdNSnd8TwaDzm71xKKbDjKPCaIyDKr8SgbuBouwgHPsvSSfb5
bx8TMutwGxuwvucknbn8xDi6GVq9wx98rWdIJvgSfBJap7gaVmSaYQUI/YTAUFF6
wz10HpMGU9STDGXkAwfOyi+h/EUqsfZsby4s4RI4dxgAhpxbzVpUgLyPM8GqKIdA
E3Jsp+RxO6E87jBrBhXKKhB45E/1feehmgqNbIARyGVbRJMIqU0ftD1+FD2dDBhh
eZvCErZ5NMG8tmJU5zuRBymHenX+SwzKI8qii4p6ffaT/LRsn+unHYZvsS6HeL2L
XOPKYX+KFrG9cs/8GmK6ZaX3mN60OEChSlE6rlZ4I9fjxltuBp6mQJlelu7KJWoS
YTzzu5opN8sMHqj2BcuSqCpd3QnJ0u9K2IeE8Xw19cOKjFQReVqL4fPJO1Lz85BB
vGZzjFLdmjjaZw373oQx78ls9gp77z8Y9jBp7luYXRtN8Hl3/06T92TV0p0g5Dr4
+D1Fe7ftgkVVUeYC10sDOYNea9Z1neXrPUbMSXgaAZlEuoj/z/I7bIlXdzY787Qr
T9a1VY77pulwIZQ39bo2owdwWvUH+8qjrRkqqOoY/ZydLw19WmLNu7auBaAIgMt+
XhCyQlJsMmPRw1vhD4wdtlbEaKMgZmle46VHB6kNf42+PwXhYKagiRkePJLZN80F
rJkGhRiTF8sa33f0qVbjILCh3/btE82FfArV1Hrh+tw1iMh6Dsy0rqeDjFFiJBAt
l85FlBYIRVxwJLNoVmSZokdr/0XY1Q1iPNUdJE3fCJrfWj5AqmO2IZgm5w94qrX1
1Ov+SBGkLTAfLCjRkkz9Y8ZsTJ9XYlZ1EqxN1qPmSq8gTv+3+wohxG6e61X9DMEG
1PR3b+zMq5GuXGmFY5VHUS/hXQZ2a7M5A+J9rHrPxo09kGANxtbOtSdtxKIFPTFk
nn+gl3IBYRCk3MAXQ2cC9+k68BPKLyqLj4ta/ycoE9/rFxuejxeu8tg6vkb0OjTG
1Yi5LfnwWS1owzOF8mbcP+4/hfJhFD92HexWzgdGo3R1e/DLYf94ANz41s/D4Drx
oJbr+1bivGrLH2vgbkatgg5lZZ9nbRcuO6uzCUuw9o4Qv2FsJ3MYSUZkJ+C/axPJ
38fW4gBlyDSyQj1yZF3SR8Nu29yXW/0yHhlTtFnzH3sQO5V9n4bMShaiueypcEGO
xsVG59XKk0or47LPzJj2Zbn7dYvPP4pwAbqgXN/ibhvIMhn9kRrCqvzp8E6Rp90r
SWpPaUgQHhQfkSMOSmMYidCaGSgJRxwlwRB9JO3UeNrxQtEZp3RFno69JxyEWPT3
lg+odk5qs2Gw6JMc8ADZuDU3x2EQA6SxiYJ7/LSsh82jMAirE028lYJLx97qldku
9sNK0bwk0hzCGLPZT/lhiY2XjDk2aG3KoZYQqERuLA4mSHdMv6ctUGoR2MCBlPmy
ImraASnpCzMCip1HLczaXcQUZI3iEs0FGzWKE6ReyQE2Xs5mtbD6vqdft2C41DVF
BFSrZXx8FueZ2z+/ogcygInHV4kSeRbSkjpfpRMF8PVyNZ656ar8kEWymdrp2joN
MMFrxN4vtTGRqVKxsb/a7r8BlToq2Bd/Wi6Sj8NWBciWD1kTMQ1giDAmKkUy2v4V
bHPareUBNgk/52zdyjGH4RDsq085/nxuszAT/ZZTMkEbHnAiySZ4iS3tPDG+0a16
ngBGvW1kDP++hWFQCg1ylWYlmYqHTn3USZVEruNjk3KFgasmnU9l+UyLxarLjSKM
hDo6eufgBCwGqOWX2yQafUm4Cfy4xvLuCbNu72ld2aVWs0z/a5QFvhD1QmPE+ZvU
lPAtpjvD7oM2wUsI4TEJPydEfAcqTAnk1tZn8K07rzuyIk3VTk7SYDHCtHkixz/b
8dTu+n+uP6c555eeKDXRHVqIGPXgyJ9bPW172ZpHHPXh7aOTIv6PYKBXwwH08xES
ubfZPABGqsIcoM+z5ulT19E2Qb0sIFWB/22VanbhAtHeQD/uqjwfLBUK8S5Vmjp7
ILyCQ8kTYO7HNPurlbHVfIHq/0HShKgUzDZD17cUtP/mj1W/4qAGjCdxlLbq49og
Vxq/fmxfkxdyh9fg83PNmp0DSZHl/286snoNJRNTvRqdk13RAOt2kiqNxDdnksap
RnKjFPjjwS2CuFZcPohPva/zI958C+Zi2p7OJUdr73f1v3wi9jPOkYdwGtEr5/MW
9RRv4Yq7vTL/oL5A1aj3Y5OH2A4iQRgOfAKl7Htf47r15rMnk9gzKvdRikfZF+E4
Vg7lfSXrarwkOAuWns+VbbbVmdhUBuT61bo4vDLnO5dj4DphSEpT/CYy2t1bOlAB
cNUyk91EL9S/I93GmhskeTDflRWm7rX8MX+qjZMlYEEEOf63N88F9DcVVWvZlND+
CdhyZwk9QVIvemdRpzlnTxUQCOVJAA/YTQrCTuOz5OfktJ/ql/WXfXMzma43a1pW
HALQ6wPQl7VTIBYdHtd/qj1YkQPFFJ0X7YylVw+8eXfPtTOh1CHJvlu5TTQOPrci
amYcGOaSLBorpoZbG++SoNbtr8tRICop0XCGzmHIMFsH5v/yB6auDBbgKcAnPxxX
PwLZ+AUoV3K4LXcrtFu32gKSPolCAKyEKYlPTII56I73ndSewCWL4OCPhLeD2nZx
80ZhG/5M0HIjpptGrj2BYz8wokiJL8XcQo6oO+ownSzU1GMSNPq4h4yGrsKhG3XG
6uTG2UqpE+3a/VhzItBF2wFbqSMcmOhCLADMJ6AdGkZVuvWDFS73e1sLF+fMCeSL
p5sSbZxB5PzLIV/ys6r7N7Wta1Lq1hLmjU1VFbJbtxuEVheVHI9Qi/wt8ayHwbYA
aB4ZlbyjrAXrBI1zr9AGPXkhSxhegXaF/DXgzIpMhCpOy8HemWSzq9+d1IFi/xdw
VNC6tjM3KYn67egsyXfnY+toSUlgUwYERT6eyPxAzT9ur4yfSDC5RT4420qoB1YK
zO3YMcpImjKQ4IXjUtl66D9hoC11YkvydtUCHprKsDeGFKcFvux58APv4t1EZeNZ
BRsmTK3DjbmkZa+nDpxdXss5ONWdVwChty3yr5QKBUZFVWIFk341C8KdjFv/IKMC
WSgI1z51J2nGEvS15zGvOyDCvZacXHFG5j1dgKrXHEeQ5t8ZiyHltsKk90DCXtgh
uFDoW+J1BKz9A84QqBOGrtD3uO0vUPLgYgo0pW5Qtrqjwu6a2ABy0F8MkfvfQNEB
E4Wz0o2P3gLkMNYP285sGXoLc1GS2QTCgy6EdUhNPuIcEoO2rTw0qAqC0KwKAIxs
GbH8ayvxG4GXLlHcfTqO64rdjO5amJfTvskU318S0cJnJOQkoCMBUOYBjAjmmxZP
83wz1eGv3BjXgF6N1xydX/YfkRxhUt/5Uvpmd91MlZsZcRuu/KpxCJsk2t+ND2xA
PV1qWlAlCE9nA/MR/9VZ0tZcmjjybSw7TQlgDgH97cpmooHEKvaBqHwdAnwNyfyg
VT5Ul5xDaDVliqi0DQYwTY1bZTHDavUZ0JV/0jfFehKKdpsBCMiuyOweWsIZX1CF
yiMq18e++IDLMos+kpkSQ4jwAWpuipP0oeqE92Rj9CaL2d4TzqaO19jkXOd2p2//
RzfxPaJhAwAI4r7Duf1b7JtNsLWJYEqu0iPy8PNlnLY+97hbj28oO2UwZM2uXMFb
2wFCtkWB+VXuj57hunn/VJreFHkP/OHnnfbEctRtI9bHflBffbSgzTzyC1uE97UP
X1nltaLSN6Z6+6rL5ADfXkKCqzuZJfcx4x9bMtFhYg/tOJrRqhpmbLfYBDkTEph1
dKU/z2E47RHS7w/3c2Q4FbgMMsWix1nW0/vYqLVA5j4l7+nOdrrXdWY3DajNvt+a
c35/6CjtreXSdeosl0lHcR85WtrOHXabdsVgwiv8T1s4croFhyq0cDrL8sda9mC7
9l/pBFdMRhS3y3A0QhzZlj86sdd+dn9cYD5dau4nPkQTt5IPMu4ZYsNEgc2fzZQP
FM4jvmMDEggZSjZV01WEoUiSJ83tBPslzAN8+VzrwZOmI1LvzDmKmDRjNXYc5uiz
w/UeEwpipfZjK7hmDiEd4bBYn2kEK6m8eElFjpivZ2VuvZjVJj2NWQ6sYTBiGAG/
wwiGOEvEv55zZbmZXlVJ++vj8PT3y+Kp2SyDJPdldrLh6Wb5jVD1MLMhONv5mGfM
flSHGVHa08NyZLAeHP5DNnK0824tMJNkB8zXV4ETwEFIz6eu8BttZtf/YxfXX3ld
wVnsA7vKJJC5T9Z9wodDHnllHyUl1rHZg1/JNkItnmQJhDskNSS08nzXeEwf4XTS
Q1b6HSftugWr8l7EqDKrYV9zT00AiVoj6iI6hZ4MfuC/0YMDnuBTlLPjfmlcVsML
JF0f6o0vl3UXw1/WvtbVkw/3w6lZ/Sm/1nu5vIQe2BVTpL08l9vtlF+IiMEKy89g
IoAQ6gRhD3qvrydQENXYAYgSP+2+aFO0WXa+d28sVmma+N7278dtbmujvqnrj01s
F32Jhunl1oxyeYOWC/xFMh+nlsGb5dJK2Qq12msZuz8QFnl8kIz/BcQAHUr/4F4u
MigVzW1z1oKyA51mMNnBgww//5kCfg0RV1PYWarQmDm3YZidkf0LZiOsMi/vicpX
7OfRVVLFreKFzxUxXffMUtHJ6UQTXpm1QJUPQnOvKHTaG2Pl69VUGCVh4vNtQdgY
zfiJGvtPCbBxry077nVZG15+ta7mgb6llnpSZcmPwffi/2C71FJv4eCRohnwcYIF
RiI7/6qsz94FVyYc160o1KpMpGS7v+ZwrfpKDTwvr8vNFWwmjBf90TRwG8VjZ484
4pI1vSnSB1XqZUu101jicF6ymtFCDOsjkx9D6Tt/FA9iVGyRpAreEspTxI6OPnnE
zd/rSvAsVBmbOaErPATChCvVWG/2/qwqbrP2JcFDR4h9i0JuQXe8hJBZL65StQ/o
+4w4hvYidbD2O8UtvJs8QKrKiEbPN3mCa6KCQMaRZYmzfzZ77Ui0rbU48mVTHqFM
qUWGptP6xjlzFc1Sx9Icqw7eYf/tb8EsJSSi7+0z40Zo2Hh86txwxPinhzYfM5z0
8AMJlqxmQpTTq32465k/cZBpqTNgNVStvAFItWfLZJKzGoeBrZ/5tm9ig9ceDx1w
mq5ErBLPv2+eg2mrZesVHd5MfdfbAtbLjFegceEThrbCvDY0o5gGara4EUEy1pS6
1a3uG8DFRheN5/C1nJHMQ6icufXAV/KxJkSvTCJebIkuXN9/SffiSeHZwiwK0TtR
k6L9KXjseiTUoOwvN/IrlN/tUmZK1bSlbWwcQrJJ9gJhwPxXqu7CdEDap82SSJnO
sul+dYvWs9u9tInbnCjh/CBlIwcLqm+p3nh4WSDyDlMomd6+4eTjIG5QcMdHX9vJ
+5QD7uimAseMuPJtTQxrATAB0aUFBf3r0qEgT+FYlvAEJIapB1GLuNjWRSRnWhOZ
z2a//CuX+Rn0I8Af2z1wVQr7Dpg6JKsuQhxofVxuAI1XF29wRTdctl5UoG2AEWcC
QPQw5DLZazIsDDAJJ8uyq+InQr9ojSq6CNaEG7vZAdviAzTQLz8ZlmmGuXCGKMLa
hyOikaGwNDat/XRDtHGNfaICNGrfTE9HKiOhwW2vDAmJC7jX2hqivb0flxUJJkKJ
UD1+2lY9k/5iDbCBAEgMEBMi9yskKIpC8HleHvpS4OxjKj6ZA8+QZ3tfXVxitVu5
Wq2lKAr/3NwN6L7twpoFMwBfUN+KKvD/3b2pxLBHZCBWaZFW7pElBbaFGeGF01U7
2K8V5ECIoaas/8g2iA/p3Dq8+VXCprfFvaJD9Sc6es0B8RVV8GnWLaOnUBvMMjqT
ozljxZq53DkkLoXmizAh9CFOrGvBtDCNIq87zJSiAuJI9RZ4vFabYfx3A5CK2zBg
CM+w3nAHezwdnxOSgt56bo4mmGTb4i61nrlyDQUsZihX92jL6JVFb+LT4eKjQCtH
25m2Z105yO7iwQ5W/f/7FlXwxO0F8ckIMllhNmR1Tb0+dEGEPUrdC3Un/q0eOKrG
+YFnyOgv6mM8z/Yat5+27p1qFklvrMK4RLgmwcYSG3DqXuEPVUTa8u1ZYUStjgKO
9FsYYnow9sPzLZXR6L2dFgCAJWPMphJBtwSYz8Kl3F+n6LolA9C/15uuV1yit6ZU
HXuAZ5D+wCuOqDhKzhPGejGn58xvZqgj1sr2+/xECAmXH4sWZucSqsvIU34Y1YP2
AEZWi0sfmzbx34onpXjEKOIJen6I6WZb+LjvX1Z1TDbR3dLtDnPXKuFA9Fszvysk
f4+rYgt008AXQ4vH42c7m8lFP5tnNdhwbfVYcgC2vOwcZe8LoADJSyFPsefpOag3
Cuinsu6lpnEBwJvPHL8txRCl00t5rGVFRAfQDWCbBf+5oyMSMQ+9612CEsLCmHjJ
FEjIA+tv13kSn/2dgnLx3A6sKTcU2pqqMaNohQ8PtdyIduaavKxaajvXAk15Ob5d
oRZ0U+TAxsBzcZNeMwya1x6f8eCimp1MS2vXeSQtF22G7RLmwrTUXlozBkmkN9sV
4L1Dch5c0aLyvU8Mg+th6ejOLL1xszHuLd6iit2/kZRQ5xSP8EhWXdadW/dNFgho
APiposOaSzYLdb2yDrNTZg8PzOY4FYdVMvdtAXcrrcP0NlW1goJcvhFFXDWqbJHV
zgDk5ifD/bztfcV9HQua1WedQZjdJq+CdnQmIrRhBmtI89BXBtF1ZLX/7TbqxHG7
ErsWMoBqtCZqUxsU0HGBPYEBAvLPTNBRQOS4wBux58Elr6au0lSrvniptQ2is7gI
F5XSWzCL8ZWkpG3k8ILcj1l1flgziUU02DwUshaQ6H+OroUQcoSXSHvaTEhTQNrk
z10d6UZ3pYdJ/wP7RBr4lGd+F9HEwkNGwzogyOA/tcAmh+bJ6dplldO+aamj71w5
C3jVeFUMvZPgPP+GIHrWYl1LVa78SyJDK1pnCJPazYzXlr94L3dFF5DX1O0aC5QU
JPrn6jo0ckuBJEXILqidJxCf9sxVr1fRgpuiXtfA6Q5oI27rFU80vXl5UYuOThVR
54yNeU/+jD//neDISN6DZlmWbvLWpAXADE718lPiPY7FhK9qgC3dXlKAv4NND0i6
gRkApYgG7NwUEKsPogBHmCZ6hCVQmQukaqO4YfPkF5yqTzMebF99DoCPcAmmYoZP
dx7auzg+YVxxJ0geQaYZtw2GcQBMjwYEnsiuZJw7MaycWDzVu9Qx1+Ye3dPMz2Qh
CCqeWsolh2EfGyXH1pmvgvAqIFgKL4bkZY7corKxozH+WlwZixOkV9KI7ASQ2QYx
xhpG5dr9rSRRgmLAp9Z1MEMtdZ0Hf2SJ/NMHSPNh37RGcsJB47dobgGINMBzFGdn
movEfQ8oFvfIz+dxch+VOlq3iHxgFapCJT5DNvDUuZnd9x/QnA4H35qEJOLFjzrR
FxBvJRlF9GZQlbpyVI4SUCpzAvmXfV5jJXLkc/zGVS4nTcDjbEFxD+nQ+Z7o6RBO
C+TqsYQlbuJ/U2SlzT7XESy1HVEdSHMaH5BMf2/nMqmuRclvX913xclGvd5GjBXs
fUxpREUwTBbOF5cjR934LdEEYJ/7a9PCEe31QRxQopaXgatz7K/p1bIjbz35D2Vx
OAYZwwhDpYl5KLGM9lEwLcJQMyPLM1Qp+lnvgSMVc5xmP+mPYck5PUxHjWMYG5js
HQ5/vXSUL83C7K8YqbvOU3D6ZW3ZdlPKyrD88qBqnznw4uZpxWOi8ODGuczVmpuM
I0HYvQrhIaWkO9LZIGJwRFaCZEZ1DwcfRctlqEc6oEPPvhOypys0bTrPTwKQ+9bm
PskDHL5w1G1v98SUIf89pnYacSHeDeloOCg83otq01EMUHlcN+XhZSKeKExK+Tcu
JlJJk/H6pWcVERTkxFTs5qIvdacmtVXZP/mKI3oyr0nzPq+g+YuX3VOWkBxLCzT5
Hq7nC3CK2l2610G5rb9GZqJCT7Fj4zwz/3WRMWQs2XgXuCdBxBE1w3aCY8dqhcsa
0LiLkBPQ+PSdwY9fBme3/zy1i0kH6VSXLoAj5FW4GUd9xxYoDTFw74aRAp0MLvKt
xFMDCaDt1A6I+uH+yXwJZ4ZPmTn4VxP4Nia4DQBZ3d0hpPV/K39aVVVY5dwKUSpV
DV6qMiIYiw1QnyW2ZYmANHI2aAIuer0MaH+mocwBoUE90HxKGBD51GxtY1M5wFsP
IVTtqbbhX7b4YBXwTmIqrwqi7xfhVPqC5a95ddRTEOxpYXnAnnxxCD+xZd9wWrRW
HpDwa5JKbS+IFfv5St1Wuv7U8Un3stD3jikPgkwuezUpokLwHJBMB3dis9YirBww
/gWiCULem6iXcuCPon7E6ML8PTDzOYedLo0rMYL4vYhEazKXSHK7ULT7haBzkNcA
fWIeWxWHsOLOxAOK6KB/0dusilz5bxVFEyY7XDBa09t/HQAeV6ilzZRB+lN9xT7I
Nq43P3Zhc1++IelSG6t8278vohSU2I4vZDheyULZSZdAV297fowTv1fd0LiTGnmu
HMwgWXXh6qsunjh+qSNiM5HpSgbKai2N+/MsNR7lYrfHmf/cwHNmFWfMCrl+jouM
jQufVdqCSYZw88nscdLnMB9W9+4dbuHY8jLo0sWH/O9szMqQfKT4EGlXoJ7Dgch1
LTKld66KorLWYhYE8gyg2GD/S42RxoRBGTI2pjO5NdQixOhGSO2pst/u+wB3rW/f
CrwVSsIrvwZ548jB+qRYb2W42/lzVLFkLgRbEDJh/PE6Fi2J8vzY8KUonJy7Rhss
Gw2Cf5Ex+k2rakOgBUDKufc+/aN9j8kcONWwvcqSvPpml0MSy0FVUIbpcM9gCw2K
ZBRDKmJ80LYhkmSToHiJREUeTTazd3ZDBiH8+Gd/UM4bn2jI9LEe37+fshPEttMy
856zV7fsjPOM8yv9MQxIme8yBrljEupD7Xc6FQe41envD/tYyTRIzAXfhEpnGGpD
5Y90jcaX4AJU61ihFWyOO3fYgGYRMl5EwbEpkytHKmpjRi55JwfU4Zm/1pzZBQYJ
mG0TLMjfiFO130JpdCO0VG5cdSZ1ECa0JcISJJFhlKf6duzZMuXK9XPGgLlzEheY
ovkg7hCFsIO/dWSqwzHbu7wI6nzkKfN3V9TR2baDHdkoq/hmUdgOXOWB9RR/M5gL
RpF3pwyhOrZhFvT4dGClAfTJEyEf6wVW5wyhkkVIiw3cfhj9LSJhgjCWV/HqcC9f
NPEgTXFs4AOoDfGRCb+ik2vM76nGV2dnUvCm9QWeQzaV128qP6S6PYAV5yRIgMch
2bLV1VPIosyU26mx0uWEZvPssfoogJ3D3VEx6sp2O6MTj42zjPa/4lB2DfyvxpIT
MBbZseA2Fa7NdhaYS9D5+PDlQyu4LtoxYeRK79Vd2Eolz2WIkoIrkuAKKZ4797Ir
xrC76mGvfcw41ceX9WXnxKTYaXxabqUUi1ynEE7RvoC/qusG7PtYkCa8OR8LkO2S
kkuCE+/2luqSqu60bmu8rfeQpWr6xWMbZCoyMROtXRrawEV+Rwk3K2ptW9zHClvD
qfxo33rTOYY1yTPzsE6tRbtzzYpcDpGYLQZPjDvBXgN33N5MJRffDaZURJhes58d
61WWgpoT2h3EasVSVtfDybzXUFpUkSrZentQbkO89Pv1ALO4kXMs5XBhXo01VBIe
X1y/wJ/nxDfrCYalkPh+vEuZgi6YI0BzV1U0f4V64Qo8KDoeXqx2MPAO31SsHOVa
lB8Bu9MSghxpLhFcnbVPiiqrjwBG9F8cd2B8L5iU4N0bC3dEqmxaK7IEf9zHbPm8
2bjqCqnEuhix4KvvYvX0oDUKgpUVkvThbQuEA+b/QN2IDBH9WR2Emo3jv4Wtbylw
n7gOAj671W6TvsFICMIm/ESVvvMFBIDO7sIoZuHDOWf+625VnxZURgtXxV+IOQEH
TeZSnc64ufZAbZwLZeAgo98Jpko+siNhykstdEXaR2mMWziMlkRGC1FF0FpHTWHQ
g4bNQ4NpURkMb48aAsbjS1PIPTvHWlqEguXHKBAGkUjzofGHOJyx7tsOH2v3Dchw
Ib4stNeZu5K3zOf9DJ5wCGw6V8smEs23kXAKhF7Jukvmpgw1+TAfHzybCYY8r13H
PiT9Jhzc17j+Wh2jNsE2RgdcHh2k8hFkYv5NjHzo/ZhJjadTRBGZ1x4mLzUt6t9M
6C1GLYE6hQHB5VCYXAACPm7siEFvIhrmai0M+EAsy+JLRB5EolAf8cOYIylbehQA
I4gSpMiiRYAsCAO8YuIo/D6LyUk8Kd0L7l7omAAqPBsd1Y+wuhg59CchuM/mZ3ct
3GvKAhweiPcrbnoz1Qlu0s8eydmnJAIMbg9jN9apaY+jkNL8kCmMvgWTQ8yTpKRR
Ylpa0phllqlj6wx4T5eFcLFynUaqRiX24jyA/1jHx9Ig/Gnf6GreaVzjs2/F0skA
QyuI3GYQIeiE1F6xA1AG80vWBNP5bG2L5OSLxyy285/eeOXe7KkQ2I+emGyNsBoY
mbWvzpi01Kpg037gD9zx/t5lcp6iCYhWT7nOdOyi4x04PPCWCMbnG/ZeYUF+7sTC
Z0MxbRP5pwe4ZzmzXlRqdNkXsHxYuNRknvGMBqgsDv7Vq3jhqG8nj97UtvPvBXO0
qGdxo8jlULOjITTneehFNrmRokr/GQwyZ04orjxd3eJHDdybn2esUN8PeZg7JLVW
N7PAkLC8betz88JB5ZC+dbsPS1if6fJygfVQF+DAP2D857U+QhmuwEpnKIt/Dp4T
fWm8yyJim13dzwQameeIcLgP0nYl+AayGfQ6o0Nw2A1pHY4zxPVUC3Tqm1t/PXT2
Mus6G13XoWWcG4ebU4i9DqO2p6GvfomNfbS/1RVxkvnoDHMIhLumvd2najk+cPWc
SVwIItqTzrO+UJvPNwNSsuI7vbfDd2IiF4tXWeqRarp1YLzt429jp+Qrv0YpL4pF
SlyZH28T9RX+siO+NgsukgsXZpiZOrc3YKlhfCaWeaQ3LOQBHCsHMgqQFoKsHjZy
+6ifzXn//Cuur182IAk8X8lMc4fzd3h0vXjwK2TqTh9PrB1TPKpMgxZoeDKouJTX
GY4z4kgxxB6fFELA0QuU/c4NeoFNaXYTfH22XWJunq5WXXO57f3ktl1BmyKbeGjc
0/3Mfx116ObTs9I4XMAHTyTI8rW8g8j4lHHomBiWIAl7luRvwPgyFyWbiXq5pRLs
Mexl0SeDB9UDJhY9rGeL9AJ0ulHXVOi4pRMyDGBACB30cZWk2IxvGt9QJny7p/V+
8coASHhWKR9CP5hN4VZA+yzYLsfaVmyEZBDSVJZaxiNH8xAIghcaZBf15fqHegK6
4zb3WRXsZztSWf7AgIODcRXF0dDmHwe2BvEI1/qG+42wpQlYGSL7iJJbP6zZusWa
4uuhAE9LywbthP0Wax4UF3N/QUlpwZLC2qUiVmvTQ57puA8O0qpha1slkFb4vgoU
17b9zBq6oJ9Le2KUpnZwTDHLJjjq9dx9zkT9Vq67gprwQcQyatRzfKbowNrZtUbR
HU+ViCnqsHxtpM+CQtAnT+0KaTq8U3mUHGbZcEklEX0gECD9d0FXv/OZev/YpwYT
xi72mEgFnNjDMtGQJP5fHoE/ro1m/VH/8YPS7q7nIDNjNQYetr+fiE6Aq/yLI9PT
CwQRhRaUphVHsQQp64qDCLf336aSBPwF4D2JKk3TWLt+3GF2+q66rhYQdWd2CPiT
D0ZYwTm3pL27G043EYA/o19aXeaZdcy/DQvjmmzmjqRgsDPlLKjMfDvcSr689IuT
NMguBHfTd2TAWJAyy/Cr4TFVqJiC1UnNW0wRc8sXWUt8x6zkD+BUOSuuE+LhQp1I
lWH0pSXqjYW2ZE6tE1bsRP8rgi7YGTm7H2pkCyb1ffUlEL8eLSACslVjAmxnfB4T
y4M9ou0tcs3sGJFwfNsmP7RVBh3SjRCMklgfKgyvrWXY3Cf0xcGaARI+fRHURT8d
lzEbZeMdaRlVhKXhdbBQcuXzjj/am7uRyijf4kddlli1PyHrMaJhCpb1q8hDmVfb
eDnhDJbvNYvLmVTQ1fae+u8SYzg30+G6RV/pmelVrbGhYKKycwBggdCeZkBNj7os
94/V+kZULGz4m1AfvyJZ+scFrtPTCaRL4k3xaMe03cgp57wighyeUCUDeH68KPjR
hEpoW3SWwmk181be3B4m37ns3/csBmZDVZRISXyTMMYqkV9bjZExCUpxaAPtZCXU
OM4HNk7U6IZqV6ypGQ0cQCu5DNe3XKQ5LeDJ6r6uX53BTyCES6pYaxl6rqWH6oEq
eyKxDeaAEnbk0aao+n1qRjBVYpd9GRGwf1GkkNio09lSonMQdpgOt37r7Ln2ROJ3
4wP2wZ1F+SmP3OgZx/nDM4sZ1UOX5yY7bkS9pZjtjqRtE7n3ws+keOIGwyFFvA1C
fvrt8i//1gQmImORcFmhJsSvQgMS3v0gca/vzi1KlVnzOtHgIcwGovnM1xRRFfu5
Tf/jt2hXyuXjziy/sDxCKWbaq0zB21+wtln6WN/lrC8tjrdyfWUTS/SJgbdf4VDI
RbVg1ciVwSOiChUIutNpY1qM9o0CQrIqLqmTZJmCZGAWIKf2Kzg8WwhUVWwL7qna
JBLXUpz7GpJ4ookDT0SYYCqwbvGYYjt0eKnft3i+5EVxJJo1nBKGieYma+vNp6Sf
KQasx5STOT9e5sxT7t29uqPU+4sBgeobwLDXtUjsvT8LYBWvqFiHawb4iP9v8ivo
pUIGhY3PJ3i9JFtN+k+5zjuPeNwAk6rRmF4PPBa5U08E5DEzRMdLDt7/Bq8u52Cl
j4g7hBW7o4aiL1LrTQsIh8wj1niSXOU/c8jeRLP0GX5XC87qXSf0JYcr2Ghh5FV5
sgB2r1lsvcJTAPZHAajw066HlUhR9doaafFvY5AncaMTxMuDHmDz5CGoneOa9Cee
W0pIr2Z1jS9EGWVZcj0mNBD2mhm0OLm/a85CKkWkyNjyP/dv9ny036ecz3LKUjwZ
yQ+BgpZD2b4HQsr+vQO/4KAQcSiCawzPd5vslgrNvtyNDufNlaqnecCb/8p+lq6Z
UBqwhWMlNutIpujMzSS3rdO0XwPV1pSjm7M7ZyEnTlW0dC03VyAQianJ1TnQTyZj
UbuMlNXirYNQyQUkZq+e05K+O/ot5V+Y8gJID8KFo7fqie4TRwdabzefaBiYOuBP
0XfUCYu0/oD4ToWHmTJs95gJrd9wAHgDYAvJk8XR8rlkSQaJRDpHW48kF/RRZyJI
4zrNPw96bWdYx+niznFVD2jgxLRnNYBFTYoo9AokdPbbBrHY7Z6jNgziW3iw66/b
F2jxuZ7sWtAKuzyhtCGkQurrAqZKgh5eMSVsxY5bY+X81AoL5LfOQ1MDi/5XBQWr
kD/gXf7Eny0xZfoVpkCCRcixgbKIyibAMAMAHVw5BmzDy4aYv5/UVXxaVk6G/5XU
ihk51Legzkhb1bXHehLRlzIyHCqurRyFUcmSu8awRMbKLXxLDYF0WXkQbOvcvuwr
jHnWt3EHZm05bsXjLFXdMNurd/1fg3ONkx7L6W4eyNlBVzVGHVuBvhs8L4W3Vlsc
swNO3ekB+fCP8++XiXHabPQM7nGCa+ovTZfY0wuVVPXv4k2nstTUquxep3pXkSa9
SIkoBJ39yAHqyJ8+sR4hjLxRB+mrwQF4PT2oxwaCARUuVejAnHEnN9ZPT5rFeEhA
aAsz0uZWhTqmqPeQRXGyckY4d2nhdzGaPCxx5QforfcQJoUWzq4Xvt9W4bpjVAIw
KJqcA7fb4qaNMGZ0DYvU5A3bmDHO7fSRjL9B90VikvVVbYKCna3/Jfwl+0FCMWO6
DRVDHNfdDIfeynlXev2QErpCsXMhNmygoF6wOaqFtWJqKkOX/cqpNkJac6SCdWxZ
+6QmWeHsCjYVU5J6B3kNEh3NSSpFdXl9Mna8nJppEVOYKs8HrgBpxyC1fn1tPpSf
NPJ+B5ym0vdYNWpyyoyQ7yLzQJN6sjz4+up4GaIry1VO3Rd9ALO28Lcsr3esMxdU
maV5Lent2tuv1DcjDnYdYOgzdPDzx295i1Xpmx/3x6n1KRm/gHoxygZf0DUvn81d
4+QIp/hBz73w9KdrELu1yOv0NXXjBpJ8OcJsF/tqcXcWCLLdYGevqVj7c+DWe2zU
Yby5e9wrlXLvijR3xgN07RHGCwbSdRqmy2foCxP0OGtAkZw9h9Fq6iyc4ZFHTBrv
975dMADkh2fY+83VF9e5VKtxSF3vMdlz4uvBv4vwDnaYCL3+msBhJZsuQyBrnJrc
u8asqQ+XbIxhJHoYTOTGHk62xjWQMWhr/TxxutiaiQSgu7dxwtkiRFt1994oi5xL
RzGBUDwPGtK9y/pmoip0nDAvuEpTsUoxI2JOvMf2xtU5bI3m1BxT8lJVg9/H4omU
0jKiECVg7Nt6sW+AdzKCVtEDra2k3dUSOF7Nb3CKGtJPQzPZaWosglmOk95PRGBk
PDvJKnZpnZ5Yb/vYEYaX07psp2c51+0bJ9vg3u1BV/KJalh4dKCzNC1FJpVHe3ll
hHKIOM2GlG3hCIkfvvVm1wN5KqxbO7Y02Ni1h1bKhm9yfAnM8DGs6KJcquLcKsdu
HDkUdFVyTewKn5jqrOZfZQbDGPRzZ5CEOM3MTdSz50K2VOJO7xdYGTbt8fqAo8tA
Qeo0MOoVbWQvVXscCu6cz8naLYfRiH8Fna+PQCK9YTsF6GA5/afrEcNhu/p+zozD
p13FiHuBj39rGrkCSq50jz2KMp7ty8GrindSujXXai4d+SukMHB9xZ9AE9me6FRl
dqaKfXF7CRxcQQYHyOmXt1daopEu+N7WfikltGKiSHtBcwSaUOAepmS0lOAEXlll
m8pdMeS+OA2InzUNySnPnusTS8fEwK2nVM233HFDvq4sRjAan3lxJ3FNQnA4lGuK
issuS61xxwXCGWinvpzLO2aJvSNT2PyI814PYcqrgWdXYOR7/7AQL5qv0lZuGVJX
cQSX6SibxkdxWPf2sgpiQpTRyZdSWKZI8jc/moEMrWX4PxjlyQtKT4yPt15gBM+G
1FVPW0mu36qXmltwRLX8LIAVH/38G5lKp2vj5nZLXXqHZTryGLrxsJ2sM08efUst
aIiXOTpdgJN6cmRZKAOrFfPtOZvybx6Q2vrkCsOqiWkMoppZpm2aU3pBHyhFZeF/
mxIjwtFGrwd7prg94KT6KuQmIYGJ2O5moIYiuMC5us499DiHzBCtvE4JdV55W7rV
frGDkRnLkrAeqYJQM9AniMobRy1SZNE/2WyqD5wvDT7rDkAmpobXbYHjwgKBxKi0
4MSHWBooBeseF+R+clycz0XRvn5PDlFgvgc3ccYEZ/h1Y1msKJ4Wmf8lMI8jFMz5
qf9P/Y4NO22QkQivIMs/CYCpeIUWEBI1iRpyzU05QCzXvBsLaXj1QtNakRfYB17F
pr36qZUMWVlE/hW81Jfj2C02SKXWLqccPl5xOZSiif0ffDqNIdbuL0mtAMaE4xDR
EIxo96noejtyd4Z7BdA5i6Eme6eii+HdCgfKYf6nm9XH4VfgE2Rky9x7c1EvthPE
I6PpJFcoHVZ9ne+47pE9j+IqgmNbxnPoqc6sXe1jbmkUUz27fMeihDnyYtwUoM8n
emMIA2C1YCgUX1HLpNARL14VYMwDlHNhyhlSSsdW7LflvO7Tm9VvekdfiTybtSAC
2c3MMtDj22xssozGEQx3TMuZXXopbk9hMfOCp2JlsQNgPaAgM3INVB6AW33IPDCh
rQl1ah+2jYkpBhQpFZIb+5A8EL6QO56KO1qcWnWFUvZjwXRnkM9GZOkkRWEXYk/1
sHRm98VJpOc0Vohziu6RbRjLVGNgZX6ZScseAWsFE25pzXJJdxWyro4UxUaPqA8r
AQCzvyJfQQ5aEvhEcx7E8po+yjZuAvPqLCLbQZ9G+YHapehxaXl2TnUS488qbz5V
XhzV7THw/zTAMeeY4j0rwqYm7+KLCbxypFp/LT1++XuFXKqKZzS+PZuGGxeaeUih
9caqjq/w32HojeeWTGti550bytYpXGVOXbpH7qHryNiJT87kKRoDtJsSMPR/cGO2
HAFaNtr0MkEo5JO89AA3c8i9kjiTKgwdSSN3NhdgVRu0nilfP323Q8bGacH+TGbd
FWm7SXL/ezQPiJWDxQKej0PcnC+2RQL0FtRxrhGaZwF1Ak/4GI9aBSdkGa/8gMLk
YcGcKobAOCOOigjnnT1orc3Hz9WZ0hL8qR7vVZUFVfxNgUfrWTrEM3KEqUXdC2eK
OLWXKjnxuyk9aQ/h4GdtrfCeNQYYgQ1/R2iLuWbYAJXIvqdhlQy2EDBi8f4cPjHs
fVcRWLPspYNCzDghiEvc0v13y8QhwO2w0dSFVVsW+audYFdl1KeTBTOovRwnAS3y
wUP6iwOJ9jaQJdYejfTbqYRXyRYa01nr0gxxCOUnGHz6OXdrVQVB8AOIUTqTb26Q
cvs70koOJ8g1pzGIDyTBhiLWh1rhd2peDLnVY68vCf0XMskzp67CK7skK/TTQuAh
yi/JqfvoZZrpYSy4/meJRFm39l9W2bDgYMCMqxgAHnUFrUGLTneKUI+AOfUb38Zw
2rI2jCdvU1NHn/QYh6jTUxdGYiDl6SZ2MdL1d0TMlVW7SKGlAxnLuYq2Q4MuuWo0
89xLIszbC9Vve94CWrY2xMRO7eNDuy0p7eMLF28kq2+w1it1KvFMBeAVSwfHiPr6
PsJRq0Rv37PYIfLAkMSUE1EHdlCXHNow8rfilc0RPMBw0sPn2TbexslIagzDWhkC
Pe57piaHNk+Qg/x+hHmIjrOSxC6GlMpp/3IkPW7k7ernDKcQE78TGnNfRI4E5sHD
OrurI2pmuc2ghdRPgtzSv68CKjD3olftzQfRk3ADxtbSo92r8vvDI0Wi9g54UxEE
oeE/1awNzOBvIj/pRaxBQqlhfaEXpOvriiTAclm/OJBEzW1MESprdstrPzvt1yXY
lM5hkq4n61VVfHYpn3cw2IAdH08a3btX0CkF3eD/gEcW734JNYsDe/m/W1KWhCX2
cjqDJ+aLbUa2C/ycHce0dFFMroR0vwQKbIHogQXo8vJupXzn5vw73KKGyxza7V90
PVEo9iHExKPtTFCymChZ+rh9ki/TBhwZ6nGL4ieOrqBPqUzViTyqAkBvlv6EurNj
sCH1hpxSR7cRO0K1CX3S+jgvyKBGoNxs5XlJLSdfyF00iassrA8ByrSRNRHrlBjY
v5W9CCjL78wYVUqOoD5i+WENakEI5fo3acDaktdL475tiCHIlFTcUndqvisN0uOj
2g3MD6NZ1S5XsNFvcIavJl6+BUIL3HnM3vAiVlMXh93uCkzLtC+HrkeCz8U3wizq
bjhdkQyow9A7fy2Stz6aOjfZJO55bkIuYUkl+Hp0tzp4rq2+ndnbg83O+4ijBb25
8QgPGMJIN+4w96H2kyDnXWGz0UKkvfPjNH6SeZVUt2/Ye2MsQ1aPqFMMTOZI3l9c
gKiKhmjYOrAhraE6Cd6OeKkGdVFK4gKJ8vgCDhSAzauKSWqMsq/a+aSBraue1zY7
ror9vUVIQW33EmwiOBzI3cmpvB4ccjvVNw0NZwpW9vhgU8q067mDZceTDv9CM25n
596d5HNo5fIzi5b9fX1Az/tMHVVmyPVSW8V5HgvzibaZwsKGCeiTZqFqbiUXHHWZ
EVI3oy852weldSh9AxNkoae7vAEdgMYL7L798j2v5hA/xbmZOwxQv/BRZe95lJs1
9HcbOfDsPKco7hxu07vPU5V0Aeot36+QTcDe+WVpeXmC+rI6NW+MkmYaRMv0Scxt
B9PWCSVPJ8CpSY12nv8uai682IDbK/NJyyNtGQLS4thSWydopemXs0cOAdMTNY4E
0HNzEYyi4uqI4jLPHmYFcMx5IE5hL7CPmYdRnHWf25fq/v6vHm2takKbB80iQUQT
tV+d2l0YzCmPvArgFrQBbY1de24BTCc8yUPdlexXzSjbw4lr1MhTkudcjr6wqdoo
CFslyROZL0zIXmwGu1vnQM3zmadKl0ct4ywzsayu76jbwhtuE2OUd1rHEKzJzEyC
EfdIr41G+QvWfYgXTxJOLWMc43DcmR98SNcCZPzUzFQQeU+yvcpyASRv52j0B8ij
ZWXLupNnDaG2u6/V5TNUSLe5fmyd4N/FlwvwD+rp1DYBOceNdGTKwdEZ0oc7rI4z
5lbj8nuvrFuOfYbPG5Uds7A0ym/K1OkxtZ6v+W6t0MfFW0rqafPBq/uTvvN56C/y
eRggP6h+7i5y+q9GNT4jFoTPXkHB9o+snjZx34N2qJfG4o00EUEP8Edsdt/UIOnk
C1fVbSJg7WzGPA9NlRQQ4mLylUuklVuZY5SgH15p7jT/zqQiigxXmt7gilCjp8Li
Xmo2R6BrVTiORVYF+UkbK8G0XsB1rVAizHWxgCGGRRJ8MoKi8OlcSqZh8KmyXENe
Md+bN+wCoyXH4RBWaukvDLDa5Fro8TX5AaD7mh7MnVM/2Cep0xugL0iEVk4BFIBj
vg/5DZws9ZSNoCUipAmUW3ulf8MhY3Z09P62uxvSdgu7cU5dxyL+RWG6Mz7Yv+W1
+M7CzB0iMnYTVut0Mesiq1T7ZSE2mkPed1prUUXZ7iY3PverxSavQBv2iQ/wabIg
BrFeA6XpFawwITHlIweiFdVUgtUcd/IMTW4ljNjvdDrhQUekcbh0ocWJ0y311Isp
pdfn21Cy3hkr2IOUDXvacJm6DSzQIQ9pEDPJFyrWMhTpSE7z0njhTJtyR41Qj91B
29qmplfF2KFQj6rJxV6d4LpQYn5fwTf38h8a7eLDgMAlw8prH7aY804LceO5Y1ce
49P/l6V05clkwld0rrzANZqVH+6ExyS42BV+A1qbrJezzSGeBacD0OkfdY5tCuz3
rcMErn+cPFZ6hYNCVUkxOB6NqqNcR+fqvgm4iXgxPAsasUl8msNUmoFhz0tw7301
koOMbb8yzICPwAh0qAEF/WBMC9wCXvs7vBySutZ68KNkn8iWglEOheNzlakb/H+J
+N7zdIxplMFJag+VCb+NYJcag8KbRoFrc7MoftEG/0wlbIPwLXkTX0VZ97XUo+qt
mm5CMTQuJcUmHxoiDT0sRG/W8/EPG3XFUdRLNX1ncaMivopJI3QTc+qdIa27Tz4N
8VlahP6Wfr0od29bsSji/wRrxHhNz2+GOOr66mxnHdIy/dKASy6PZjlp5DhF5aLS
s5ePlHWC9rAr676aihJdlVXShIw/JTpH4qt3SrWOe6JmQLlilV3f/Y8AvU5nv89+
I88vU7h9966q80eyzo7KJgECendE7nQyLYLpu7suoMBX3bKZMDjIiEzWRBd5T+v0
oUwVoRJCMJtnbzOFjPMDswbZ0dyC1el5tWVeX415hr86JjCiE7iBVpJeDWfmGnsg
KA51VTC58h5T860PH9tz+ELOZL5dnRG8sb5cKDuGEA0be8ipSUUxZmtrRCQOU2ij
jK3RRBGnmehkst0imSUrfwkVPDv90NA0QYouS9tIc+hMr+iLrkcFhJs3wAHXZ6RE
ZHyICM3BYBpRe2agqKFEGTWFSTAdEG6D/n0VwPteo6ggNEASdvre+YmcVC4R+QJj
8ZYPw+LpKh3srLkmmJFtEc3n4FnHUOI3TRVZeZQ4CL67xoji5wLaeXpTGed2DuaH
dt5Fmy2pxYr47cdVnZgogcgBfo0MiP1U49cHB/mD0IU82qSSd9ZRTaShr5XLzMCp
pp8yEOqgcdKvJXSQeqew0gM02YQonlrdod7llFwSoknFukzEFT1Dw+u4I0ZLDU5g
Ohf/wChXYBqg4TBDfoN9OAay7ze1cugimtGL7kWF90OH0j2uCfbh3XILBLj7U0ug
4Xht349e8Dxwdy+S5UBH/dl9d3dmajlVp2Et6zAYuSyctyyVSTKiHK15BvYwt5s2
LDIWSeHqE/SKkYSR9LTflfkrLycEpvM9gZ0Vv4dAFcp2Tb4Bpt7mBq9ZB6+pJyjx
bhV+48hM6+NdHoWtURBpfXYp8aLEDZVjlh4hPGfyTOVSZB2BJip+hzEovBQJlmQM
vnNuVfsmPoHZMfLtXrtXozpGKBwdLhjeJh3zDks3iwIJZPownfa2eoQ2pRi3SbFD
4BvXI3H71MQ55LLoPmq7OMKThgQDm+eXlmo3KFDeMC+U+4kXSXMsvRdUif+ZI5jW
U1qV6EHV+0+LVHuBwv6/lax10JGMFck+n3YciZY3cgfkmovCG4y7sAsWjwlURcF/
Q4HkMt30HDQP6c/V5xe08r3eeG02dBZ4pluKEJOrNzPej7zhsS7woS49sQNhgXZa
TiNtQMg1EkxQGPoKzuTbk4RaHV3tn8yOIUa7mYe4n3J6ro7YHyHIdxnq4ro/gsVS
CUdn17UYcYpT0p6zD6IgpF5ZstmNssGA33GX+J+WiQggOSCZQ/Xx+UtvB7yk0VPA
L3eWKsQINhH1TYR8SISUupHjy4/j0Q/zsWQaU3NoGohr/ZM1+Yjat5U/nMOOC626
PluaHiBcuz98B6UkPs4n88YILGPm9tjVmP7+EegfRiq+L922oi52TQJpoo/vBGB3
aaBuW7/JxhB1dLH8HuS4Rx6S+Ijr5qdE04KUCyoby/HotRQ2YWuzSvx/ask5C4Nl
I60cXpgaQMJJAgPVUINhLVm8fYAxN94PM+HVOk9XlDIwydm3OlzpO9L82NKDY17g
0RMCTbmmzFQhCxvTWO2TZBzSepYqyM9B2G6urnleMooKtorJrWiP+NNIQRjIMtUG
VNbQd0/ZdNR/HsPdjmNmvOhkRFWSsfegpnusBsRoQVM86ZyemDYUuKQxiGbqRHo+
hUU3md1CAillfLhsZQeLrnslzPXs7HtZSt4WqERZhxnuuFB2jyTxXAsUdADvrHE9
sadBjwLwK2XnTJfftc7DMCysxmpPhM58vV7yFIdqGWe0AFFKuYslHmm/V+neqGrD
oFx+i2Qy8uXUM2mwk1bd8ReLEqf7BVDcgT5d4uYH3q3yrIeXMjOxdR5f0TRA4iFr
rDzzrmUbPuMaUG1OphPtKLXgn9Cvy/bRiJ+F/6/FUv747YRYrQCfL/heBW0MvnIp
tSCzoqDCkKDe7+EITJwtGU56Ztqoq2ntfuWwp+k44DOVYNKelOy0OBveu47DLF6W
QtkO2veWZLE7p8dsXSdR7j0BslpIETQ2wUQUG95g6ydw+6sI3V9uBFodmnu36xGz
CCn4cCiRIGHzXdZh5otSBCOQkE6+2Mc6hpYGf3QF6F/gp/z02PaIjrrMFvLM5nuB
BOAdB3apaJMeE5SUwcJ7Zxtw9jyAX4OVDmmQnptlEfgv9reTGUZLWuQ7+cR99YaG
lIi8A/loHPud7d+5KP3y488sg3KN5s+OJ4rs/O7CDAKAhuNHEXu5NIIvi3a8lyCk
bYs3P1ciUplD1bLceNfmgA2X1mgA/nJRNBjFBu2L4dtc0wPYGPi1jY69ghQYw2BL
TtOEhXLmq5St+o6fdKBPEjyALxAJZLqKdv0M/Jw9ePwtnvudPlrYmhGp7+cnBu+/
6PwWVZzWU6AyG+K4Jebq7p2YX9On7kwD47Hi4e1LKk164d74aOb2ly3LZ4FWEjd7
KfVDhhWBIhIVTd/6NWdPxkXhNwMmuxUQ4Fempbnd65hJ5smLNeoSXnVrbL4cZfym
VTrLKssXMe/qE5lP/BkidyjDWlY1A0+6KfAjAy1TjIBSLNpsjdqtlfmTPD6iYfYv
4tN7JN/ElsPhL9EVPRWWum5BaZ6j0R9ROGL7smH6h42WXlcgkLI2EMz6pOQkhBWF
UegKQwlIvPVFMVojSLobwr18tFVPg4XYczyOvsBLgNTFhbm1PeL4mWFvF32V38B2
3boCC3wklwxy7ZGxJwrJq6+ePc2O2XSneXocU92JQrHFq7WZ8W450eM0NFiw0Fi9
1rR+JA1/jcQLN1YJ1cHea/OMHShMQ6X8GuuOS1wn7jcpDNp7EJ7uYZtVvQKDVvBu
F5Z3SPckuT5etGPJYJsSbmxVVVId2EijE2DnzOxA3LFZT3zcPl4tggiNGUcmM2le
D62z8WOvRq81IyD0q9X6E4eNw5zt2Q9IrsIYi6NmWt6mybT/6rrVex7rhr95l0D1
5h74JDau0IOVRM3XGbYwJxtbBvAr24KIp8W0HIIUnxL2/ShwCftCjIWd1IAfaCi3
HCNANptl9EsJ7St5dpS8+BbC0js/c9jkNiGxTLoyz1V6C4Cdyf/HBv16gFJ5wZFB
6D62ds0qYBrJ3ZI48UVqfAJ9qwPJfuvuN9duKNBjSKV4WGW21coVATMQoy00PRO5
vvbi4UL15sJJbKQv49CaUqARJeEQalnlDuITHQTdApTOfVFxGyxR1ON6i+cp68NB
7Hkx+Fz6vhjTvdGBfXB6FSjqAfS8mfQ+hQV9bKHXeHiF6jl9KaXKzG2Y/HJj21yu
AQW1Ouhu6PoPXAGPsdiF3YVsAX5y7zZ8UV7+dbu2Ee1rt+eNdtqMRjloAdsm/bGE
+x4AEtHm4B2n3trDhDYf1ZXQTMa2QUptNGpYX/uuV/sGd/CzasUlzph35FBI1Tbo
KE1y6YqKd+H0EU7w9EGBP6tEMtdbhaEWiA1+61NQ1ppQkbPZFpMowcklP9VkIXyI
IecMw8evsutR+5drgHd45f4mNBqKLf4JsyD7e7gA9GH/MDCgpM0WMjhtinYYSEx/
MClhkpe/uBdio4JxGaOct8r6uTp52Z1EbLeMVnlLasmHgFAfyR3LUC7dLmkTB8i1
dlcQixhtJB3PDMB5tm0ieBLbJGMBJcnMA3ltIU1DkLF/1Onx3pHYhK1mh4wvTFvY
shufJiquPCxMF2K/dtHE6GjV85lsWOKIvuVAblmfMC6F/XGq5rLDiFT1W1CEgZJu
YxvPOGELsuE8PmIpEguvS82xz5zUmGgZ+88snG1EE1KfwOV/7s30hxrb2BtRdmvo
MHHvdZ9K6XSfjonuXQ1JqGez7DE/O37iNvMorSzr+lrzWf4MM15h5GHxEp59D8Ur
v4gg6wQYOKGAvzpwoAzbuDZVGBzuMZvCAsSpno/fZBNtYXqpnjzVjvzY8kv7Oq7N
7quXkEdqMLtnyzhkJeGYASqw0WnM4xs+TB91hApKkFUb6WG7cydYHPAWYK6z2JQb
x254+b/CxZEOW/0ghJsp4ex8bhp+qelt2X8UN/lY97puXZy06tfhrprXnwRGV2dW
DN9O5/tBLTdDzK7EuYXHic+kvqqylZOdHWl4AH2NxxbEh01RcnPkBcp/1bFY2cTB
f3/iAKZEXL9Ap4Trb1ZfD8YCGDsOpf5YrMaVj+TeDTpVvBq6IRv3I63g0UKIb2+/
zFbgbxcEHPvEzc2SNy4fu1EDEx5udadSV87IwheQPaFDgqwtpbw0KTxohmykWJnz
WNsuqP7Wd6HfbgXxlKPj2n+svTF2l0KJwRtUO0ckyWF661i8qc2/JMJUmKSjflSL
QX2iYXxIwtXtdF3YseJcgO248t1vjbODBp0vX/JklegGQSbP6casF3Q8vc4GrlXw
i4cvlt0k7yIGuv0wYnCaa18J7Sj0WuL5K6bdrEItIJn9WuuMFqN4x8LqPSNQ8fBr
FsT8yXMbbLEBtF1LLKM0xdbhfhcLdHoTkwp4NUxxQjqjsjFxoq7AUDiBwCDctzzV
/r3sY+i9mz+TVzgT4YZYXybvlb1MOR/CccWxMbyQWkgmX1yv8OmojyUszfAv75L6
ltZ8f9W7Z+cL1aCYJ49qh/VJb0v1T1PGCPNX5PR/5xPMId48ASc0cmixHL3TrPwO
LrJDQRgwNmKbTmXXS/KxM2ks+QKE5en1K9uzfGI7Tap5Gl6f/N4mGbzLwHZ6ySaf
E6p8Zt3FWlxIoqbm4Kca6JYnJ7YaQ3YHiR7F+frUPFbokVg4CehKAPl6PWA60w+5
UVS8cn7hgx/QgdvvIMMaeqNUOi6mYSelRnB9zY1ZvzX2O4RffsW8hvf/BaBz2j5d
46g5bJeken3mimcrpdxwV7vxzClnrreFq3rtqvGPcpJEzoMnQOm2hgcoSERRHLpS
kgFZm7v4WWvtlZNzgqCfN5Tq57rMlV3No8tVi+/HrMxtws7jdbWDJsV15Lgp4su3
DjDNT+IcKmxrAPXCnbfwjSQlVjzfL0tTqAjfEi2+Z0gRdoA4ZDgxZQoEU8T82Cc2
Y+/wxsxX7O1Vc7dAeU5slVkw1Syfb/t5trwXCjnA4OGMC5is9/yddiGMEH2nELyC
MrBwzDBY0pUpJUGSL1cNQhhgifhNA8W3HP5vA3arXKdjMeBcos9ZbAmLIcmgMUGF
yWXUJD7PuDwg9TFV5dtKu6sis+JT9cLGh/yl9HmJwWJM2cO7LxqPQMfo2jYY1zLb
Hjq5WcLAe1B3yYpe0aOz0XwBTnQPr+cYUEWkhdQ+KyHsN32Yo7dleo7mV344l+8t
hkQuI8ksvMLdWdOiayklfatAsKTeIImlZT7i19cQW0dHYF9yngpnR9LnCKYcwfr4
3WIUdJjpOOrxXBKn4oNyicrlixpua0MS5f+EwzgukrBnuBNmc4Gp6KzK7t2bfiVD
1jXIUPl7puqoZolHYfzlZ+gqkrPq3wYliy+GcVcqlzUgko1iIPWzaBALgfcnCkDP
wEVB5xq3dJKWBa9vZ8fYCZCM/E79urbz2ByD82XYPAZzk1hZ+/XKdhQATF8W1All
GFjRH0xgy+soAfJIKB1H6rvcj6Iir02eWAyMPMHA5aNcLPAGqg0MmLCw/9HR8WJb
if+ZOpmG8T4s+mK00XU58nosdynlKgZbf0uTLIs6qc4nY+09SFUi8agmbH6frHdS
r86CsPtGO3NhaMVB1c99hHab+qnafUW6eHzT1LXIEXC4SJRGTnUW1nyIOHAWlr05
MplVcN4tcofcUUdZ9BVw77fYpqiy1EyICUXxxR3y5KkVF7+JOGTGSqV8iYJGm9Hx
+MNbYlEVdlamEIBQ+L0JsqKrlPAhpULGpAqFVibXv+jni98DkYKE1XSfoOi8e1o0
yH8/C5IVjCxTmyNevieKUFsh5FIsmwEyrJjV0TQsOwPeSvTu3QHtGJKN8MnOiZBy
4fbnnLsTLp6KR41TBorQI3iHBt2zUGzlyJ7FynJv+zTKgLAqEoNgeyEtXjTusma1
7wVRGvcN4SeKIDxJxD6hXvQZwa5DYpvLFO+UpUm4K/sqjLwezEjjL2/oqqUKT198
PW+3qaqMCyRXIHsIkbat4stBj8YW0qWGPI9tUJYLpTamrcZCARs+Vjmn8Wil3y8/
SRXakJjURIhiGY/nI2lFclNqqTsUw+o3NPcnxK6kRJpLwk/NsHYs+5Kx9TSjJwy1
4HvQysMYKGLudHOuN6/FsGy1P7AWWTxY04rtnDyuoS/Z4GllSaiqKdCT71IG56z4
5wxzIEkEqAwnrGOsZrNgo0VFl1RJmuywh5uqyLplBGa1FXNxOnyH2PSaEdLVRZoT
fW+BJhS6CcI5wTDtEDT9EuU4U6TT5dNdh5Pzb+EQdqWr0/AS34V33Q2wYuDktXdE
dnjtw+ZvoIlLJwLJpTcCbLOq5kITb5fjnApdGHN3QdJeQjgPsjIHSqka8OVHsmLr
9+9TeIgwlsGUuGNDYSzylOVB+ha2tzlRt3/aqI/pWOI8KcEGgUWJJ6GdukfoDoME
m313oL/45TXRe/mdIScu9Zz0vLk1ARDVkO7gEbLCeVmkVX5ujjdna5c5T3HAAbsE
QX4hn9G7tlHp2339/pnWrPDysIPlWW4N4tXQVYPvvRbqAK6kF5RvGhEC2Pg7Jfnx
JIAriBeIaXoSUW72u0I8ZhYdOCZAAapQWrg59IGNWlIq9gC12wF9EL8xL2J/LJI6
/qfORHsCGB7WnOWakLlJqzqmvQowPGXYmpOUAHEp4JIcpV3q4oXPd6GahTLbzoCu
MQ7rXcRvX69SWZV7od1SCAp9yvATiDfbCg40jPrIeUFNuDJFo3GVoGphJQSOc+U+
uJLbYJ3YdHlOsBmWPxa1qgr8FaOoS0P2SKwhawD5ZlTKwhtFodKkiAW8aqqeN4e/
t5NAmE8hmd1uSuTsYU8iz/SWNnt/R2YclgiVyijZuHgXo1xJu8I6T2k+e8zJFRmn
0cT7gGOpBuUyTcP3ZnV40hrahhwatH3pe154YeievdQ3kNc7nOxTGyEFKqF/kwKF
gX/L+mCMoIdF+UHpIX9k8iO7RP/SAD7nuMwhLdB3dMzVwUbw3nfaLPagxMRzt3+g
8KYIcfp96/ojdWH9EB9hbgqb4e3ycW8Qd9Ms1U5d01zQ/63tvcxcCUem9eA8O2WI
i/5/Z7Eq+2C9j7khPitwxKeE2MtBF6tJN3FJvWOzOgWYrWkH+moGGmfmt2DEDs89
HWRy2TmAVpZ9wXnvQH9Mc2wUZcFbMJtpuA3sB7pyzMnhN9mCg9PfjDmklFBogSrB
piUL6+iRjIoKf7GPRBkr5DrtHT8kLH85z0Pcb1IEM0JxUDbH4VL20HYS0rKmyk0L
kDlnHiN/GnPaPJBW5HG1Rxz8oSt5X1g5lGudhcs3rlDXu+xbxgqoGJI/b+dEMy1y
nOxQFfmkiqUcso6cKbRtBPKOSfLXDiaN9hSBinj9HrMovfKoEVZuAzGJeVjRwePc
En7h/YM+G28bslQFBts76nn0dA0F9KaEHY/Lsd4DZpeJhohqH6bylh5SFOnOHvls
ypeshZJhOb0XYnNKDH6Jss2RnNZtGNXnbkNj8zWTpZFke5f/oMri+Ehuy1ZJhKqY
rYANwRjI+qkWJaUV0V1ZZQXqdfaZ130LG4u5DieD0gQ/hRLs4Eppjzqkf6l++eCC
lCRtEXBdvozLQNz+5M8XzFS7vyVBV2wpGMwoLGtDdgOUuB9UUMeLj6PGtY/eCt/x
K77qlBI32RnmwgLUAdhxeGm87hvz4vi14nxXfq5Tjw/W1YK9xmnQAVWYWQP5Akrt
ltO2nlZucAuI44XUSy7MlUUCB9dpOVYxLvl99P4/fRMhOnqJ75m/DAub4ZTZSwby
L1Pjyx+V3j+91TVPUOq36koHE3Ji5RTzSx+yfuFb5MID14Edo+rL7i6rlJ4QjJyG
Z0qew9g5e7uE+ifrZKIrHFCgmsGgTZ/60zXdNvs2K4RKggtXD278219JVUb0MEnf
/S3c/ahj08spuaAbSoCjOyEuJZFGtz4cY+b60OSvfcKZjyPhDBdPsFrL1LdmJDlF
BQVWXcvWS/9WxzCnI9R5zDDjsu5di4+DpizF/PPi8sPRSAjExdPeTO9a8+qUCicL
WHhTg9Z7Obx2d6Tlpv+Rj2lHWaTlFGgH1rNd+tXLRwuSA0+71zOn905I8mIF2iqA
gfarNvcU5AtME79Z1aI+Wen/rxw0coYxNNbUeTM+7EmMzDVsVsC87Uy/xqiZxPkk
kIput/hSMrHjcHER+kKt1PHyRwx/3zjVdgWNN80glk9iYvPhp9F8n3usrbfGbkeK
g9CpCrIV77WJ95q9ULL0nE3aqNhhHpV/0OMYg/E+3By0y6axircPCQV9M3WMhHiZ
gah+5tsq7NZyTHiNq3iY0hq8r3cJ3GVMZaY7nBUGj8pfUD5SpwcMaXWBDkDolk3U
ZrsGH9VgfyRgnpsJveocjR+mnlu/XffKIg8HqTbcomzUDS7hBHH4Bgm+On2BMC+q
UfkuAbg854Ho+wMLpy0HFgVubQJy2GNVAnXDm5JZePotburCEfJ6227T9+9fr4Qm
XyEmqn7of6dQ9pdHwkAFgH44chbzYoVtpZT57csVm/F1VhmtEtrD4o9PLHXIcSfH
lGruf2WcnicIOCpVOrKA9HEW8uzYtH99t5N6FEStcA7NarvtBLvMLn5yKSoSoU3A
aPZ/uP37tJeHBHmnPwJ5m/quqhW+Jjp+Ick3hdbRtVj4ZFJKj0/hKWsKIYi1Ov4C
5OCNVtqlQnN8dPIguPcX/VsjuX3GE6mbZp7HdwnHIWpLAJm7oGgCpJORF2LC2xkI
Z0p2T5QJaNRPW76LVts09rxmiMhGIFuUaYHk1PxzdMTb56FR0YaCcZzL7JnbIai0
CZZCP/o0/SkixG2iJctz7KzV5V0NwJ4HWVS+EwHS5uFvM5LkHhzyRhIKM899Qj7M
Kf1PFf6jhpDT+O32+M/f9cE0i7i3pV/Tq9UBKyZcN25Y1QiDddI7aURD3Qe8uQYN
J+E1JgpFn+ZI8jq6815QUanvyXlUcHuGpLhveZfiv9XlNIWCmQsRaqDRcFjs0GXx
E10sz9Mcrt9LUq7z76r6OpLBT/l2pfG66/CQDGm5DwA7fdxsWIM/cbirfbyWPCoc
gmthe2nQ2NhmuJU8zwthRpiLLEjkblC2ns4YewSZiI3kFsb6MxdKDWNpfnEOeZvc
igwNPtKiWj0zKxnf9Mkr8yTcfOY33em0HsVxBJuIWewFKDvU8EAyK5gTkWCWrO6+
JrQb1UdETGeHPxUH8jrqUfoDXezoanvZ6AalptXdpPVKO2zqLVdYaaiDdBVWvZcB
zYSrfC+De3kHZPo8UwVVN3ACDpmeYLFOC9BHcGS9OWuQ7vCSL4VpCp+4gmVPiC7Z
PujM4zkxq1puBKhhaa21dcyZGwpmiZZlY2hm+/TcF647ciZAl6CMUlMKvRX58Fkd
5sbl4Zvf7x1S4HjEKdtWSQuYHJXPargWcqQbWx8UHkLoXeYs1Kfah7qr0WHPY6HW
MjKraiLTIGflPL6ltt7JB7R+eD68NaJ8HBGNcNeI4o/IQ1a1qltWeCRDfSLs57Az
LRj+OCqb6IrXnQgtOjEcIxn6J46tFCXUh7GIuQVD8ycOVH0Jqch+2ZZ7jwOtzyZG
C0nY1KM1VoRXurUJu+BvCHV+RZD0zonMtgavFNez03phfQP8ldN4VIl0FvZOgMb7
xOYGy2sYY88WJG4Nqff2/skgs6AZ/q0IgEP5MPlrCdVJPJd+Y/A139vzSYsicLl4
E9VLFiKYSi4rNIliJ+YGnOkr935ISwmGKGu4AyWFSJldY1RapSAjX0en71absuBc
rzKVYgHMkOiCf+1zDqAaIK/7XQO60a4SfLBxCvw80NHtNAm4Voo616J/dkgo+aQK
QdH+7j/Uj/PSHZ7x2YFsItg3WLRSMhUo7u9byTrm6nrYEnQF7rMPX61Zi+8nbyv3
DFZoAOeKNUFIReBgo4JARkuKY+BNFIM5AC9LOZ0KoN6Hc7fj+FcZhauFDRD6Ce0r
HfoUiUYn2+YPy1GIC0e8Dzm3dabsUwrT5w2fFU5lFxcyBkfDCEFRqLoLR8xneb37
ITj0d0zrobHhqc2h2PlkmT0wi00vwSZOkx66oJQV1kL2x9skjwV0JkCsIIXmSSfa
+XziDWmaoJiVgRyYVgLUi/A12EDNDlIM+qXtraQE45R+0mRR2IKrhVYRAPwoH5rf
kPRvlqSQJmZflyYkmyKo5M7X9K+vS4r3HZgg1IA0jOYrtJbWN/KD+vCu9ekxB/xh
+r/u8Rzy6KMNhVX9ACY0Ub/dpPbNWvpfHdduyBY6Ndxp6tD1e/71lLToaQ0XUE72
DmwmejxzWKwthXJUkKS0g2rqc0iu+4eMHp9ALjpxN7K4SiHeZeIPcxSQmdCeRTel
4FwkGn7ykB0/ke+XnPJEW4ZdylZE/wr2u70PnCDva4tRVoOKedEmJwhTA4fY/8sd
9LrwkhCMegDpfBHs5CN+QW0uOnCAQRdfqubqiD4mGO+LhhZ+NuovR6X9hafvNjzs
xqoD5QW3H7weNzhL/m3SUPFepoXu/y9DYml/1nkKPQNPl9dVpKwwohaLN1mDyXz6
9PFg+vqt8RQOEMKy3zYVSTkEgweoubeMIRFNr5Mcauv9A28/A3SzYczM6kY6dIBG
1TXWLBRp9QFi32GIFYMgZmU5p4QwUT4v5ayQrjrLZz18f5rQ/ImVbvweNkX5PQGL
V6KRWfPn2iFTbjH4jxcbLinBNzTDmMnZyaBNyzBZukqzn71mBlO6qPajIJ7mL7HO
W6/FTz++n0zSEBUHPrdsVAbhfGnb753Si353rixXIdjdUXXAbc0VLpph+JIepWe+
G0zCPtyFggmX26OdSlHBWO3/BdB640oxX/bZC2RX/puNPgVV2KLrjC9JFDr9U/vW
L7ZrC4IIZkIF5ulyo/MNK7eLhPnG1Lq2F/jYjSVCHYBoYnaddjQRcaqYQbl/jaKK
u1obub93altnn3vakMnSrnGpnBVBg4y9r9CC/kUJiL1NyjQlMGF29TssCbUbi8+g
IHmm2hASIT1c/mRmNPaUuIgm6utNqHZHCKQ8ImRV7XIlU+WJ2elbsT2WZW6xmc8V
4hCSjJEQjzSy3ZJofBnmS4Iu7AwW82xDU55KtdHJ4TEM94NWLhOz52o9UundXdYj
Wd4EOctZfOgHc822vVb+ADugK0tk/8SBz7Rn6zWn/s7NAqb9gVMR2tsyU3wYtd2E
PrWTZ9h5h3ub+V1ZCNycIxSanIkzOyfAutIgs0c9UbJ4gWkQUM4Ow+fp87KSU0sZ
IcKwQeOFQ1L+ihcYC7+hTbJtO1jLZEFqNBRKHCbzUYBA+uoqQfzmc6+s0ztWksgD
kj8tzoJ1iqF9isztDfK6ZZoczV2Tswura5qvcSSsBUdcmh1G0cc/RIG2WuX7Tods
ZdVAqVImokzJy54EG6xhZSXbVEzQLAN6/fsGDuuipfxsrDo4v7ynZF4sAOVTJ7zo
UdBnREh7oeOmI3m9pQt68j8RlVf9NcvT0npjhZZ8qL+o2VCo47CDxPy76GkYxel5
YNq41ypcLb+Kyg1ob9Ny5r5P1lJ9mAHc0LSo91uJfOPmDaQ09T72a9Bx3+3VblrO
a+zlhH9HI02F9uJYDDejgIUtGdt+eaLbHAnMZuS2rdeyY11HNEl2o5lTtBHpgU/d
PJvjFtxeaT4BLykaWoVGTa6noUgucuDU+sxfXqva0rLU+f69/3sl4l5xkxIe12Q9
hWxXxp51VlKvmuPMgILDU+OgR2WbuEG4xjDpGDxQkq1nJx1kxi3SDnHdl3MFEdao
Ed1YhqGotwrfslJ3Trw9braqD8r/MvqPzXDkEwFxUAFeFmkanEsQFC/SoP14CK2a
A4LKKIrfxWU0oSHVfoHrv+V4tJ6YxV7JSgOoQ2J8d/wMPhnHKc+ahuyNIcDw80+R
xLPaTpEETTtS6qBgbopTJ4noIYKgeIs+OT17fi4iFmxEwI/DTDQF6RttJbmsSZbX
yJRlFgOLt0wxC1cxH1wTPEJrQQgSfCn2SWzqHdmkZ12Vbg/WT7UYUTfefsGXblPl
4+3PyjdC6mpC2IKY98jAgDDtbkgSWFvpmSxKSm6iPDiZzl3cMzIF3cdTCslCEMi+
2AzEEf5aMkC6qWfDRPx0J3fn+krus2R3/kBNo1yP9yq6Fhjcs551MwVpcptVUzAg
By0kQSzxyNAqEPU7rW8NxQpw0CMxvAIAhuGi3qu8EcAp+u+hSyW91Y4Kire4H4BZ
QysXzpGn+yrxkWHTTP0l4cBVpB8zoeKdBzjw+/JKbWNHEFDc046naidcTp7tAE/+
3VHIV2Ri/CawOg2oRtWN7lbeNhosKMpwnnjVr8fL0pTkxwtjECdS/nOESwEjZz2F
mNkJBSZV8/SrGSltXFP4niYIlayJ2ONENHGYbsV2fBisgXunQl3RuL3zS4bWcWFR
ExxgomJOFctvL23XMETdo+4FeFn5QNyCGZSLXspSmrBZVFWjWYNX10wSatMSWDuE
tymxQLsO73Vxa4WQjhkgmvBHZrnRFimlz9vy/zxWcHilmmT6hfOUYQsw8Y94iFuT
VV68hCSeqnQqWVzYzvmKvhoRium1UjG8DcU+YO/52OL5zhyFNxWbawabukoA+vM0
sppQ7gAuBnX6A2yYjOL31jm7HSISG7xGO/UYzZ21fShMs/Cj2eDUcsooQoocXWjU
1Kyoh8H7Gb4uXPDG8rapI4YVNrolDJwxoB9AL1g9BDJkTx6eMtVV/nkpRdN+zYDZ
NI8t0clTzz69cqg4Z+wSheaLPm4fZV7JjTfHQIU0hEM9Ot7ZPYIGoGoMBocLRSMy
ND/471R7A5FD/pvJpkrklqQ6vbZkUlT6YEmG/GQZfphGg1e3x3OHesZXHn1bsZco
vzjQNWwCaJpP0uMIE/GO90iRYBYNj0kBoemkSAIz+ku+lDeJdeuV1B+oUH3jUzBd
X7UWoGX3FyqGK+IoXe3UqHbjKCMYnttocuk0/SUR1VRIoVeNsE3M/SZ2dSX19khz
QaggYoZ1LUTipOy6F+5dVCoJx6OG4By4vLeGuyfG4IAzOMMFJFpru2zPYo2a/hW3
G6A6P+Q0ZvR1ftHTXbdpGGNtYZoI0yFo8gYGmVcClRZZTRHK5BTaysywskIuGRXK
W0QQndbmWu028dHDmZYHU4wDyfVEeZxYvpmBrZgeXI42azLiHN5npj8Ds5yPjfgO
CMMmyJos2t2CZ4WAilQZdQjBCTJlR7dktNhSF07eXWhC+P5WkR/9hEpX66Leak0l
3fK4MgjMWxaOh4/NDJgJzl4oY4JyOf+zAXfNo0ZEZN/1d78ezUnk2xywadpVQvly
TiW5MbJ7U+PKNmu6z66FULjNaLdLdahMGmtL/AkSPVfiszxvLf+yH/YKQaI7k5+S
I/Z5Gj1LFlYCCNXjOzde0vaLfBq4ldjGrMayKxr6WX9vyI9rMvPSUOpGlbqmoWBG
ZYdUt/8rP4HZcoos5MXtVMbpfoJuHRcfBePNawIXVXf+rn7PghlQHpOcGEdImOKj
SfKKaJrEcUpdMyyAmY3sh8eX1AyS+gua9pGKA4QBVnv0yoCmVaaJPB7x2r8lNAcw
lN3qu95NZ4NUK3wB6FLm5uEd7inq8Eerm+hSq6O9BghrH7hTCeNGRykpuV43vglS
BSuXABqU96Amc4GH6LJSryjAVZM6KfmY/NwAa0PJXTxxNPN28B0tUmON9D1aU55P
hViY4dJ2R0/62YqClJlqf017DC1KpmzB60YU6aUSVT+G+SEhV/NdmaVQz1WwQ1Tj
McwbTi68h6SmqUi338qCgohx8RpeaEoxlqoWsS5ZebDEJdac/7ZcjEC9EwV2bM1k
uZSROD+ZuBah3e7Ql3mXQgHra87W7ATBoOY7fUc+mUHCdc2CAkvuQWVhHUPKbYcN
mYRT8FW5Ii6LqZ3V526mrLoASDPOg2FAQvNWC6ZdTEmHL7GPeymTR4I6Bt1UF/bK
Y1lOhfCaFdChxrWZO4ew6wJ5l3qNr1Wpq0ERqIf+DvxQ9C+o+rcaGDg6GjZoeB1t
fdbM+FGIco5UL3d9fhOfT2K3emZAn/zK5f3geSitIjn4x2PvEON+5AobbxLV3Wu3
ODGJ+hLfcQCxb+/cK//ydvf7v/TwvaUdO7cWP/0ffPUz5RmctEoLPWom2hjAY50Z
htou/ZSBFCwYBjqtT3n0GyuGAbIR8BlBWDqJplAaeV0Snm/MKzCnnikwB6CCPCNq
3pYpkOROM8pKeEELcL2NhEi3m1Dl/fnYQWFPGXgeGgduAujQ8MChiLfYKLRNGKoM
8NlqLJlE/HkMy7cOC8LitY0Lq1x20vwXVUkW3KFuNM0zKA5l3MQGS8sQf7QMWz39
QkhboPWOlVWsAE+wt8Lax4kJVUYFeQW4n4oPPi8HNSq9b619mfFyVtxR2qZYFHJT
ZKGP0Zxd8cBWbQs+KG/HAMSOBuG0fVO+G4/jUjGeYCphyJ/ujJ6bwWLXY/KJ9Wq8
BzWaiHsQeib3NGE3oZKQrg+hkHe8htZosU167fJHse/i3cfn1C8E8wpl2BPaD2i4
0hyE5fcnqc3/I8Iecw2Ibp5wRMLDWSckf9mxs7qEi9kjeze7IZtuK8hb06sIayfI
hUbekTNyE6SS43Oacf4f/pClyhwTeHR03qdJ5c8pfUW3dhX7cf1FSXTZa7s28nY9
M31nt4rr8sGH6ClJVicMfloJLHh/fZ22qmB22QnStXOxxFBwWZhhFvu+gfnYNyBO
kv26K8KP0XfRiHiOIsC96JWAcJ/VMAbuRxq4GV8Bnx5u2iFAIZ7d/vyXzuCcGb2z
9ECW/KtoU143zmMLNaGfcIdIOJGrwG4Z4zKT9EfsmczdQVJvTKjg5/SQsb5ZcSCw
X3BDDAjlaIdMq8mcI+edxnpy3V+WumFLn6jZczXXkk625b4EQF1Rwu1foib6hWWX
v5grACDcP3OVn43i8bOjdRHa80efO0XJ+61n+hyS2exClTzyW78scfWTiC0vLnPi
heLbSK+Lm/VhvkJmhhbbRXgvXinoZn7u5hbrmjLvaubq6a/Qf5dnLwL9y506BWxS
maCSA6W40nmx9i+TWGuO+3+d1I8i0ekrp6pkK+UuqqigwFYvgom6MDZ0eVejtXUw
slClNBmjwfxq/2/A+QExGrR7TsfomAP/zXOBA58DZBcciFsmtMw3k1TVlJw72Cpu
K+DAbpptH/FHlLUg2lyE2yP/E5x5MiATEHpsi78nAfTIiWo+Q9Azy9qXbdvNPufb
fJS3GpKFiD7sswyCd82b7JWAC+Z40W42sPGAmvadbhdWB+bxPT99wvEfd6zcj+0C
+mOFAZiScZNXT7q8fjv/hAE3gGg1jDXK7vf31QM4V3JIKzyS8emwdw56GH9V653q
VS6D0GoZ+JkWgqiRdYoNyefytQc3DIzXxzunB84ioknvRhYanvKYg31q/v0D+0E2
6QVVQXCOwC1+klXGpGos9yYi8r+6PojH9Z6htR/LxVSfGvRxRfjdEHUBSpC99rpw
Dm18qMi3wCZtar3Zm4Jt4RIRRSk2Ytqck4jZA5yVAe+nazTH+arTJZF5aMeJIu/A
9mxcXTmYdtpokoI6VCbzud4SPFzZAzMvo3M9p3yRNf1Z3yLBB6Y0pJLkd7eelZmr
1b9uGUv7ZDkNRXnSVfO7DhYv4EcOyYwFGlYk2IYgGajXgyKYFIar2P7n1urt1Nxc
68DzeKCxOGvvUnaLrtsVJ2bYGxWZ1LcF6trJKBc7RLD44zye4a7Ld8f4+Tft55Nx
lDWq/gqkgbpC/gAP7YStzpRluBLkvbEEKdSQg8+kCpgEkVuGTv2BTKsMe+3/EKK4
Tq6AQukd+iEftrOtvwYzrjlbUKNzOd5BEsYJQq3y75DSWqMudpmF7IEYigtmBWdF
kUSM03z0j/26/eVK7kIaUGpYwVtYj4FnbX5FKdBmekRk7FTSKf6ZjFGpZkEwhGL0
tqkdcf9CNULdToxHBZkDvahrQ6gDzBuJT1J60cAQbLOz9JMeZlgwTZgcj2/VGdol
jGgy1Z5Cb19m+gX5uDkAkkbSBpO45fiDvCiWU5UTFdN79M8YTQwK4H4YQB48mhBf
wQMR0lHxoS0Dfd9pZ9QkxYFZTccmRuwXcyDvY2QhgemBWT8vBFq77M39vBD0bo/7
4T1A2IZ9VhX8x2KQyT4qnvUNyetglCvjLNUkvdTnPEBswuLO8ixuKF+p9/U0kxlX
UPAUaHY6tz0aR+PBw9EmnD+02Z2FRIS7YqwZJvWISe6Z5W9z2EIooK4ej/VqPfLi
69QrUxYEWUIia9rH5KB4m/78oJS+jl9emSwhtYsqH+lv+Isxbr747p41okT2LImr
KTi9Zw739ydXWTGdz7z8QnlzhgkCHn2zVVCsB6ajBBeiw904/Oj2XpVaLBLU6/my
dItxA+Chd5JEyRLsBKHrAQiQw3smBc25wYXpJ2zMJTx15Ckf9o5x4JX3JuWKFomW
PxDQARvbZ4TGQw5Pelu8VVY8uPVuvot9oCaHoTGT1Pc6liQLkA/YkmhJZwoJztwI
tg8ZViTC1xPpC0Ce7yAOhs882sFbJfQ7NdS7ZPT6P7hL8LWiPCoQLwAPFkct7V+H
LPZqPg3yg3PmF0CxTzewJ+gwvjPvDOYIcsnrMD0hM9D9uQ6oRwPGAroYjmM8k9te
PqspqTWo5ToF6Zp2y3CMei5C0HZljgG1B8fl5ue2UCkyn/l7If9bOKTsgyVgPYj/
vF/zS9UlK5g56kpHbWIQQ9vNskxpNFCga7NqWKbhciMJD3ydxrhMiDHxDbCbB66l
P1TcOES9GM5CjMmlc/tPZdEeR/HTjtXaur+u2qttedbOuqtHLrGzMkbHA1gM9z4/
fSw17CPNShShLHfka34TcX4zgcFzYvUnhm7s0EcpJ51v3AEEGDjnwAHJBOqsMQLe
OjQ7TfGMffcmXpqGUfZIgd+nnC07DsmpKClQ6lM3DalJRbXVB5sZhOR3CeBi16vZ
qnuhIPRq8AqJKILNxArOC8lmmjrAatewe+FnvOR4P5XptwphyE387gqrN+0p7t7r
EFQa6fS7CR9exnwlG5Dg6+Ucg7ZPGoTntvfuIewx3VX6c4JtiYMM3pRLVzTMmVA/
z4gruyTGaOCaZ6TKldbOyRJ9/bAeYOlF1DN7IrxMW0jaFLDoqOO0kJ/TQ3OHJ3MQ
kPqMhfzlf9qCLmnkLPcF6EZUU+a2PrhDI1Kz7TX2uyUsPuhWS0Fof9PgI+MXuBHz
rKMt93JSJGEDCInlHKe/aBLLq0gbRwdr607Sc9rdSttni2mszCFnCI5w/ndtTiDw
P83Hnm7xjBFuQyJ7LKtCZVTN6D5kSA87aE4jQIoVnRnTM0uFeQZOw6cnJ9OcTL3s
dc4aGbDbjyQvMEfzh96uRfsETjUTbqgey92Ao9xnbSCmzzYJQlNMLmMaTMzK5/EZ
sL+EpgNXBVzgRsOzzVJ+hB+SXSwKAskzKH3YlX6mBe/zm/Gu7rXSDy/282wtSXuL
A2jWIZ4rjIutt9Nk1nLZTvjQ3s771399rFERvpxIORaeb2V0/l/pEdtCJRLN/K6y
hj+5wYpOnLlSjIvpkL9HUnjhpyiEJngnKwyLdQpXSaaJs4jf3eDrG/Yz0DcKGxtp
Fzd6jNuR4Ibs9++SWzNzBt1zKBnhElDWXvJp1HZJNgSWYj2bGXpQ0uHuaesXBmTq
5NQcBB5OKlr92TQYUM4jBpUatRc0C0+L9k0B3I35AwbS2N2m1gYbMbVs3qIpWtgx
YSxf8j+tL0KtFWe9eZfq1uHo/r6r59cHDo23huraIalfSkYCy0R8592Wd5R6uOzt
jP78zACdAr0A2vJYs7zAygDIX5zexcVE6fCrJ+g2jdAh2BRsFj0W8Syq6QHPKZmW
QybUH9pkXN1vAgqWmIZ0F7c9c93pJ7RztPBVnwPVSBzeOfJ9CuKzan7nOraNqWzJ
PBu5gzS9S41ULGPuYCZYEIkdM5WQy+uVknrjZQLz9QVLMdKTtBGOrNcqc/3rmTit
pSAtdonhxNoMGsKUT5fp8ZbSl/7OnXqRBFxqw0SVe0/Jun6nZLk6mOzJKwLWSZL+
xqBTyP1DMZRDXR4mfwqUTpwHlZ+Bqed9fQfFksk+hpHNZ5A9BrF9R/g8vsRu6p85
bvd2qTEnhNx3KRypyZoTiDL4vsQ0QiVxPD62BmcU0ECZoNcHt0g075NGgtG8/VCP
xcMj1yl7qrxmywdJlnSIg+GdF9oRyHgGzrim2c7WfVN+BgsYEWh470Vy1h2VAmjz
U00mdSnbzGkX4qum8riyr39dYOTwPuuONPItpAvKpTI+tFpbwNQw+u/j26m7eNRP
AB+O+W6bxDvdEjz0PqGDuno2aFO7CTJ1/q3WlhO+Hpcc+MO/CTfFiLyb8elXdBz7
RBFBspWErzaxWQg03To1jOIplPJUq2C40Tfn/2xu00ndtGL2DekW4uXam2+jkofs
1ovT9hlGEjNlvGklkBBGV9+eFJ1V9+UENA/AIi7beFv8SmxJwHQv7DNnMb2w6GVo
pqjeDKxkYYYUDmnZ+uqpM+Iem0fg+GJDmDC/usyDh16gBrsGvpPylLS1/XOcut7l
m8wNqc7kqqD03pybku6g2DSWErlZq4KqWmSO3Ez8/odfV+8iu3bzKJv6uLvBrqM7
n5EWE1ipBZVTpgsrpCCiaPTlHL4v0emSXmRBHoDiDqeoa5Kp2o5F/lyhy129sSqV
i5HgfJnKKtiRMhdI7E0DbwA1pv9mvsrFu47iEDtsAuEjXG6ubdS7SYz95MEJoBAl
opFOcmmiOMMx8Cwb4a5apwoYaVxkxOfw8DB5MJatZ6oJ5tDs0+ponbaazsx6cHl6
vPpQu04i/pkWsykNj1vMO44rJ3Pad8vO84l8frjIRadY3PeX+PSPmFbJNUMV5RP7
0ziMP6GeKrZwSiA22xsR1HRn07YTCTYK1dN723Sbj233e5tEiCgGqGF7TxoE6dWu
lObgfXlhNy6Nykr6zuZTQ4/j4Ztpt1PcDzRcTpizDKoaPa7NcBAfQCD2CFl+qxTO
NffgRyniISy+YUCo3B6zUkDjk7CsuBkJjMN6wejifZlob1Ea/6l08kX3BT8Bs+hn
VoSQO9+GEq/8eMAMoZtU6H1J5NCkiiLp8OlWyX9TJLGE/qN0LO9315gYvW03HkwB
sQz/qQx3sYDl4FNaizKqzQA/kh2F+1NBoRx1B8r3TeqIZ1Wjj00tcd/V6P4RDzHN
CTa1ntCE5D8TiPLXyIMom8Zr8xetAgFhWjCwy7yV+3SFnqCwyzYdQAAt1bcvYQLy
G6Snp4AKnOyZQuuNIrjlGcKTGYZYDoESNn9Ml4uV0oSe2Yswka95tx4mGH+QT7OS
/O1x7ONXm1tVY7gDczHJwqXSn3qKCTPOmA4/qjx8iQOYfqBRUX1iJhejM1n/Guyn
I97Nr8+FBrwjVZdlII4f8wQLZvgzqJP3QQsD++0RcXRTcPgQ/6J1+2GBhpA/qNvw
bnKIJPZC49dqWiz109O5h6Lh9Rm0qQu7AIoc+NGZUjZkWwBnDP1SPrhYj8Sy7uVt
SQI4IL7WaGCpb16tcl7xK2r2JxUXWPwyir0MPDEvMpyMGYyo/pXZTZ+8yfNNUA/R
tacaWpqDjsg8PMMcvCbAv4QS9mlZMgXg0AgNhv2wZNdaUqmNTTFsoeQqGOHKV5Iw
e6hN/AvsW/qwY2Ioh0g/lXRUTxCdAS1GclZX7Cb77YwTsSrh5eiTA1hh9jo7ugnK
wX1KwxA+aBav/UdF36cMuVyG3VdRlsOnkuyaU1VjTB9BgIKX/NAYKFgpSrdnnDbz
4KxLJZN/0W3AZomzNZYJhrb8XhY4F9KHmv2dzuhbDjSvWO3cysHjeIklvYlBqr17
PanwKfhhpIUZjNHQvYY9OH9aocCSK0qc8NA4V1eV2KasrPzGnJ7BmvDFaxVH9xYa
RC+qLL2VWnWCz8QygmazDyG4GmUJxHCCIXvV95ZuhWkn0NbDCgFGjCLuY63+NHyv
NxqggtrSJd+r3Y6vszzRzvUufiEKp05QVPx9CfMLKKsunk+LHd0BcbbSF7rQzArD
gdXRwZo0lg2GXBG+6Vloenwoi/FWYmmnLEEcPiXMWn+au3PBvqibLRVXpqOoFAH+
htIcO57x3dGvJjMYgxQl5jLYRlKJ3E64zCDHnnacBt1U6gzJTFbhYM+xALyAIAW+
AoLF3QbVJDd+mo7sFAi5PQuOj9m6QPkmccN29FFEONp3aDutahKZvjNYbYjV1GA3
TFnTYsEb25c1BD9YCYqOF8JV+AXAO34CxnAiSBHVS2a7qc/wNhQ3sPjwecC7npjD
mLO/62lslPFWqzE6i7ZRJzMRqragCN4mDYdI+W75aPZ/9OLR8y1LIsfd0lv7iZkh
ZSDGHCb/rC6k4GR1Q5dHWULDY0IVaSL7P/wXzDURBw+89PkDT1IECFoARhIgLwx6
bUOCxf8aTAA6t246hNZgeL4pdXMwKV2cgPANi/lMbpePTjBkb1MsTcpAs1DvCXNI
ZtF8oEtK9P7rEhAORSJsUqcPq3nh9k1829xxIVToBum7HWlJNsXLCql3QA3knx/m
RdDmfSam8x6vGJgEnODf8FLwoeQcrt7r/PojSNUBryY4F29lnWhBlny7aEQXfFeR
6NLEHpnNbLXX+1u/bDrsJoNYLZiDWuK469x5Li7CfbYK12Ade5RJgWaOjFa7iNkQ
XFPQ/XDiOtpsl8raeyvpnPaGRdU/V6C+1axSVcKFA1dqjNRHeiJVIxfwOAK+nipz
ALwKTMwJKsN+VtsvBFO/NJM3NWNRSPm0IacbBQl7cnTbXNyUerSNf7B+/QzLB+gV
UM2YIaFDts64f0RXmNX7HLbH4VAf0rZzM1MqgMv6L82r/cvOqk0icrOlNgpzT9xr
uPpMtn6xt3SqqmAE9P9VydPERx2qpDAk/dfSgt5SoHCUtCAhIa+YC8nDk0aeBe6S
Z2mMpJU6KsDFmpJzPknrQMB2RfdloQP0MczbaVpJZcGZJhpgLSlve8y0sZrf0eM8
a+NEJJseDlg38rgl88ixMo3Lov2RGStOsNXVKGYXdxdDphUJFVaROEqzh3W0c2jB
kzvzX6v1/LWKyWJ1eNWaVcgyy13P47wOVg2442defnQgOjKbvKKC3pxosZrQaGOZ
qe7PKtH6pFq2hrKabM4t37Sas75OW4tkcKdZ5fZod4X4q+t/IcnjL1fFY5/WgL4e
SPP7Gpp0iYOwle/svshoi2GFyDIPFaONAXZaFwseV3XwPFbDA6B6EaMoAQfGvRxq
QEM5M2B5QwwZAgjpRdOYjKiPjCZMosTprhiqetha4Q8puGq4Umjgwgq7t+XswX0D
Dtmj/hORlJzUxkR3PQ5jRWwV67aOTIxkAZoCIVE2cmAFoTC6owG+toU1NUTIGH10
h6UjiV7fkyGzcvX1HJkWNCNRHZPsopO93+7LKZliL4Fgu78KkQRW1fK6kQeOaAHv
cu/A3MY/bu/uXUN3YDNPjMkB5G5x0xRvoyaM3TeaS0TvEuf5Djx/XN8FrWw44Vxe
JrJ0+5GGpzKeuO6dGMcsx8aQ7q/oaGhgeMUrfwUqmCvpMwezzWkmfWtEsipHn1RL
68lmOD34Otn52MQXYNLreHobXtOYMvbG5zVPk2KDpLuRtsAR+YbIzLmkzOBAZv0F
re3KnLUa3eJd6VVOep2NR+bAIyl8G2c2R96JDw5+BB+RayLILx5m0vjs54GwYSGK
ND9QzDqLHUYcVMAJMfabEwSzQD3+fXjWA3zEtPT4qWjad5ufEkBqLVFOTGP8IlK5
bYIJRo26iuSmfYnO1fEml0rg0CVFqAkWsqrHdP/yi4HdKzB1sXT6t/AjDzP5JZwj
c0JhbgLnU7G+IhNzZMOz74vdHGgtgRVW+pWpX72pjcODA3FAbqDYxOVYQ8JCUDnO
izPPUXpesHkxji7A269G26C9kpg6ipRmcbx5VIrVqBuLrLThNRbG2pERiFcvuaBr
mXFvAHugbiSsdC9/7VYH/MVcCCdAxijxrWIjM4aG5UhXBGtd16Qgd01RJ7MeUoNS
p//ILAlU+L/S8WYo4VpF4ltC5qoF24MPH8D6CGc6Xo4qUEO6fHKLdZ1Zzd9fE9IP
ByDbDjSUvs+ekDmCirbiYkOYZ8I5jmQ4hosR7WvT16h96fO43I0RK4owLRMhUPLa
LcFXWA/S4Zre2K0GaQ6k4BxBg5SSMXqx1tGEvv31AAA4XvjeTNf0r8dNAd+kJJr6
kkaBVrHXNmsoppmOnSVlYNPs6vhhNlphNY32HGXRscDIvO6X/1xvWSjM6wM5R+WW
seWQR9aAlcghGVUERkFH2T2QpG0x9Ql7/7559Evo/m2YH2gdIXbuXVg3hkCawLh5
GkjwCpBsmmVY58iAsUmVukgXqTggO1G6jRtQggpPEi0D2RMMW08mJf5mAn98Fnsx
xfjU+ThLf40Fm++3Bkkx+kfwkdIyy9uxEXArVatQc83DoA1G+baOOAnlt3IlC2aH
JjIEx0lyx1bEjNxZHOGG9J17pAD2lqlt6d90r6L22b4rO+7U0HOLP3lkcEBMc4ER
IFD5qo5TVI08WEElYRnwFRpAjJlCILTDc00JlSWJEcidoNdoW1iCidI4u7j92Dau
wE1AJ1GYMGkop4X6KdbxCQsI/7NBjaQcW87FLMa5FnoOGduN6464T02/+tXtuKuV
m0MDAOLGLtZ0z1tlC7YyQLnqFWiVlPm3xdae6EdmjHallEN6w3S3/UcROO4tf+s5
obLhwqMtG1eNhL5RtIboXbqGowNxrSr7nZYPoopY/hEOzUzJzdcwHeky4fVF1Z+g
GVL3nDOq9YPQ1yraWCwhAxbJdfwTG0sNSRfYUKFThBRkrB4b2lt8vbRERwMWWOYY
O6wDWPhk9cqZelgNCBfQ+UrMpVyccOe1URjSekFm9iC1JufwsIzbACy4BM0Bl9wT
1Ar1OkkQ7viEIUBzio3yMiMYg76XEWnVMH5FFzAFlKVD5lbuhucrYwbs7yfa2pcZ
xnflCZvl+mHtE1piffX+HCTOC3n6qQa9zputaOqFrjPdEz61wy1I6jvQ5T4Cu00E
paZ29LLElY5mdbB0kVVGG0QNLkeXD+vZyLS88pIzjJL0Raq5WULtLA3gVxiyTz+f
tENQQxXuXl/f3ljBypntoSrlKc9n6sI/2wb/5SzGvgpuJwe6BqVMKHMjYA1xPIwD
mdBebhqhSzwsTYIl5jQKNyGxt5GdYaFtrF004JsE3PetuXdm5gRhT4uFJcw4fe2+
XTREx/SxtQA1Oyq0BABtIi7ijfYQGstNlzhg5fbrCh+EHNyMj3MCkdBcRP2GjiQZ
X+SmUAUkLi3omQBp3ORJrg2uJ//j1FuV75Oxao5JPIaC/5a4gR8hYJWBl49lQEpu
b7P4K/bWZkCADX8fo/aB9AVY7HwJOFJ5ccWOPTFZ5RZPa3LkLI3ssv1pIA19oWTr
D5ErA6wSJFGLvQwEF8woW7+0j6J9xevyNK15P4e/+sTZ4zu4T9Tt48/3ZETmMKwI
W6I91CaDHW0mw9xvOnxoAx9IcSnRzJQ0Sdl3sjt57p/kR+2/4f6CRv0JCo2uy/uz
Ef8W9vUB8wTJCSb4Dxg/BtJrQJs9SHCn/OkZXeOYLguo0Mq8yYgnGgIMiQZfJtvQ
KnlBoHaR/5FVWSWBq20B05I+wzi9uahf2XZ5N6NtO0470/9FxyLuULkHE/EEsd15
HveIQ1nlABXPJmqSgP4uIAFxY8n+Ulc1ve2cN/KKD5Na3jdQtV3ImGUuIwKzpeAf
Zp9Hv6Mu9W9nxnlnxU1ScAi4kQMrV19a22xQKUf3ek2ENuIFtm6+edsXungmEcor
cJ6bdN1Z35UMDyO/3nndE0GuNRgLfYDeSk9Yge+fQGjHOHXLxB2RBPvLGM+fY57B
hIUZoFZITn7SVsQsgRInoMYr7kHz536wm0NbkU6FLKY8kBSR1pVUOsLE8RxjL6jO
EnSqgldOy77rJ7dbGcfxHlEerLEzGW0uPofiGLv3yEp/T2ES12XFtKjRNgsFSzoH
GQrlG9MXpP7tvQQD0JvYRAKznYwGex3Vo/PhRfWOcAYegjn3G+Dz1qeQ02e4TDDm
+WylHxGJnxNf3o2EqiLmO0jfB7ygG7dPmLimbroYJC6wfY5A4GnSH60KwlDijXuZ
pWtgHR9F3iO6SwlYDHpUYWWNuvzWJO5PYt9DHAywDmGu/mTF6+hCvN61ruZtKCvn
lI+oIpKV4zCZymYEbvK6Skk0VuHPDUhyN6djF5zP3sEY0W0hrGDwrLsRWB+MIfNk
fDFp8VOLUqSuNbRFr5sjmDR4i3KU/8rBBruW3rp4hppfMIpse9QQCaFuOpCwbTeK
DAZ41N/YRzPrC+F9CsfRZi7r1mQTj7x5Qs9oVV3vtq7E8K5/KhyOpREgvRQ7Xpno
SaAq+6lKjnN1ziPlYQnNN82ZcVZtJ0tynePHwKH4JgS/OtqQbx17SGf0tIQ883MC
GMFAuzYj2bO5lfgWBlSOzhovefVmsba4Oe/M4C+j2MXntE7MVFt2kCZv7L1XFxEW
pqMsuNalkdmkjlb5aq4GVDyZDEuq+5PP/fuP26bsTKe6XA1qOrbs4v8RdFECYR4d
noSY19ZKUWUf6W8LAPf7RkVlp4j9Y0dwjj+EQg0eukCj7GQ+oxtV/N9cS8iRZ+M5
3nf2iaoDWkyM8rJvAQW56SFBdfQ6SBOPd1vJLWRnpLwjYgQ/FIvTvMdtxl/569/T
BRIt9kQlIKbupQYor/P5/vHGDIj+x4ku/sYATpF8fK1CmyqZK0bzHB3lYwcXv9sj
lrAMaud8ZEF3F+Sn9Udp4J5MCVYK2RLK+f0CO+4PampiRfEXOnn14pbTOQgnbJwS
s/SRSMn9Oj6BBuIys5H/KGTZFxNPvgSNyEWvY+ndF9f76xKb7o2mZlTi5Z5Mom2Y
1tDJAI9zEK4uNOmJaqcGnmSgVfFZiMDLdqlhvu2FHW5aWB/vAj5EyBA60JZHm/3o
BuGI8r0SBl/JfnC1a/EQwA4+c4GocMJHbFXOtsmKXa8uumh41FKc5YsNe/ueRHyN
/jAQScAUEvZMlLOIPE/Pmu/+01f4h5NfGtqnEbv6uQCbpPG+Pflyc0JoIuy0bMU1
gISe9Fg+Y9rJCUZBJNIte2YGa1m3gJnQ5KUVvFZjKRQfaXBhT398kl3bbgiPYd+G
U8cpvcU2/mT9xExbjJN406EZDN5Vhd/fu9D9+p6QqAUgvSe/slu+nLWs+FyRD0pb
GNwYS6DEFCTJRjr4eUSoatwjlP24wGwtCrW9v/pi8O+K2mDxOrVXvPsVivV6pKsW
6Ql+KH1TVHdneiMWpcOjbawp5SFY5bvsAbNBX+JSL6Aepfphuvz3YKHQ1XFb/pX2
1B3PqibwA3sy2gkcelKBWlYzC61qGiESH/H/cSnb05xMa81QhZATImDXaTG24hN4
hS0V5AdKXD3FBL7SirmOpI3H3E+7uzW+4opNQEdpcmO6nho427dnt+3Q68eMft0m
ikhVYfO3VkcXkp4nUBlmY1+CQB5IIYSXXgIIvuhx55s2Gz7B9cWfAyJ3CiqwD5Da
Cr1yPeHA8WXL9EA7G3U1FC3yr04zSBj1oWTyr/NBqqpcinXDIivqN2tnUcD9DWnW
GUjZhVZVoGzfYAqhHwNnjVjs6eneHwig20mdOVSj+2vw2okqfT4L1Bp9hr475iaZ
NS1emmEac+wKzBmUQXWvGB8VQaoSwA0Wq01iIzjNA9E+A2QDGtFcaMoF8uTLuAHN
skK6UaFK7wwqx3aSCKuddT8aLfEazMGqxah15WDppaOYD6osX90ZPAAf+hxoLfNg
1CQYK1YU+Wefjc4UZoQCPINGkp8MwRvn/AthxmFIetcq65uorlDk2a3+Xw8zXIHN
GRMRlQWZiZqRmI5eqnEBQJ+3T36Y2bOVyXxGsdidbOb3HW4GkacoaFqjDV26e8oj
scBjBg6vcs+BahgMChzJQOi6+nzIJSwuRdNokET5LACxdjQLesTN8QYa7qwxcK6N
6EhzD46vHxpE6KaahISa2phnO7Vv9rx9315G2aUUDT0ZJ37nl7zqWjSNWfc4oRXS
me01f7IhpVzcV/IJp0+J/bn7E32f+pVVoqnohy0w5mOpVJkFT84hHayg1740PONo
SL6T5erAm0GK4pyJ61xuG7evlFfvJPI3PsatdoNpw+ObBrgCyXu7OSceBZphlTfj
WUvzB2f6bdND+U9Tuvc/OD3TnBUea3Ohgo8xmxuQcw5jo7/50AopIdjq1/2SnvGh
HEDE1BbuYWYFlKd2Eo/gtif7BU82zXoNTmwqezXLda1pT9bmXJqpc48flUrvwihn
IiD096m7OaeLzyi4saWoc2QtM/6YxPfhxwDNTbAWZcazd/h6iQBnaB5g0ytiFghL
/sucN0K7sZkUB5IkXiyvpjGjVD2g0cnVZMGwCnBATgBV+C7I7wTfygS0LCG3OV1o
qXHA8og7qrRnCuR97lvkBohnZxsbwChYniC6rmkCXOeSA2m4MwUCYVrEc0bLStCI
0RR0mtPM6HwAXcod73CPWd9ZM38Nitp1sFcpjAcbNPUqcRF4RWxPgoB9WGmitKhQ
w6K1EiGO2BUtrx33vFFH/j1Umsv14dsAN6mZowBNqHvsh4XOxPAu9mdCFuuFs+j0
ve/eoYUNafb0/7PIRjX+AQZc1qemOEXMjozheWEnUKKSTmAiGFW5e2LxBBoPQMjT
yjBwpubQ14vfdBNpMr/Btfw92FZ6mP8zZaP9rTjOiQ15HsGUtydpbXBoVmMHk6Iq
vsH8eMCb8nKuxDCh85/X66WAdw9cmA2f85Q8tgDxg4ct0bN2UK1+RC5Zppj0pjma
0PGnv78CmpbQvE7u4SM5wQyFVnBYrqRU13XirdzvImRuduxkZtvJNm6huVYBzWxG
b633AMMMZ4tUqx2iGuiYYbm9oljE3RDSoh5xJ/Pfo279KRRMMXfRSwg6RycREd+l
OI99Zb1TFcA/VGjFJFSoJp/7sfff/EsNlyiMlbDtSSE8AxJqVBC1YByRvzaYkn+C
uTEfFHhomCmR+kOAs6ikiDQe/QkQCw6iqRpyhSjnuyBE+BvQH42mQoVgpUODPSqy
XPklYaN9xX/59Kz8SaDJBxPbsoFpg9t1qe/+l6d1vSrOvxFvM+Y5CzGI1AzEVB98
YJZBI4iQLtWg08ccx1LwmAumKdZh91Zt8qJMbq0kN0GEi2c1ukKYa+5wqM9U6rO5
Fg1fXEZQygNaRS70bv4zuOBCAlKDETRkN1N1XGHAm5teOTEFyhdMIuG3cxGPisM0
mex/m32vicCDE/3skxvjozhdZC4L+VJFOiwpppGe17sL2UiD3hT8vWcepFRIKhQI
HDelAq90NKVSnP2iZ0zes9AGjNd7exREBe3XYq90OpyYT0QWrx7t2bQLOtn0n5da
7v/XA4cxrr4gRV9NL378b+6FUcQgJidzvijNcVd6KV6FfR57Aa7mquBTI7W4uLhF
EYNcmv+1fB28GeAsvDt9gHq3vGkqgYE3RJ4+5PoYxJQGz8ux1R9pVErIfa3ocnO5
h2Y77FJr9NdqNxwUIJT3GfzxA9pJLnUiDt46NPC+FBv/xR1akSN0DLuC3FC88r+l
jrnkGlM4rGdGzKMvQYJSfJu2ue5lvBKtaLUEj3/rT7GfQkOyPVVKOi/GdNs4gMYz
Cu/xj5skn4oYhwr6ywb/EccHxMDvBs3Mw7BrJfZREVD+MtDTJO86fe+ap2uDwbRd
0DltK8VEe9jos4BTjtsQITpT2HQuqUYYpnZZE+QMqPr+8PwMzPaxq9W9a5rUAsKB
3KvBKYn3tltNOmEJ9YQb/k3MmVCCA0l9NcXpEaBnzlkOGeq1NpilhzG8ta/7Kcrn
1i6R6oMHNtac6fov8I1i7G6kfbkEo8+ritt1X3TZycduCkH9LepEYkIcNZERMcDs
EsOrpSsZrFjE7PpffWPBRcHfqFb8uCCNxBQLDwOHE55607mH0MNie7QcwZ5w0efL
ojZduF2xBzggJeiqruLFPATRtkfI8/FqgDnQ66pBad4pjPD5J/XJUiMt+1Tma7B2
0g3nADYNefxsmN0g/6DKTDnnuhmGBB429+ikB4NdVzQ3PcjwXZWIfNvaHaGUdcCd
YNLUFeRacyM8S/xAgZ1QFhLcPn+ur+Uvptr6YGo2mq8ZUiiW9YJAI5aBepzfwtub
WGZCQonkGtweyMSTmUL7TTDtMBDJjlEDgGmdlbcG+3AuKyOkjaq+9K5Ou3MUJVSG
YoSZDZ4s3/dkCQOT1UNMi8wArC88mwhpLGpra8AIJ5x9/U64g9TzB0NiLLIiheCu
fldoZC89UcTjwlCDMNJ/ruwaSMKzcTjaRIiaFZmzLy0MHKJAXGqdstueYHbtpH+v
WaZeG5oCIfoiLayrmg65CmKpxcVTOOJ5kJ+mWs+PSixjw0BevkYgvqwCT7BI0PX4
tY9A3rLWfxj2fn5WwOzgKX6i2arfEXlYMyuEBk8YE34Sjw9GQPwsT0jZZbbKu//Z
ENZhNJnzwHvVTbO1//rD9KozJ8Xq2BgPC/S6TWrqnN40q/rN7/XMY2dt/pfYNb25
TgxkN0rwV4QR3d49uKNNNTesFinErMyVy4GsXjG0MBE351WhM22AHg8Esyl8U9ar
8AsdryBrDq9kTNIPxpVVdoDywkgQUt/98cvuDnpoXFYnPEdT33REZK+V2LHlv2gT
fffYQsIGJ+bTofYJIqJmnCaTn6oRhtvbKzYPZu6nWyOK2/FzhGCJZsrLRbRlKgAc
Zk35jhDO6cnBoK+I2Q/AokApDWa2iXvv7hLsC3iSvsqOerD8tUwL/N9ZoWH0SLB+
HRgy+4COl3MNhFzIsIu6N5x0oIsJSNKVOoJelVTg02U3qCqBnD7tNOUm9VKj3fnk
IOZKi1RrTCmFbbeHvcL66cT4l/DC4QYVS9lQnAeh3MK1e0CnHRgohCMvyXFF2kf9
livZ8K174aoTS8X85KxVeGbjvusIoycan6JcIdf/eJhnJjVKljvVMxVhvMow27fs
SeYqEaqwt/JQw1oTspsO25z3QUZN53KXf0J6H0AvnjXL5HYckHXs2wXMkJ8QLncw
mvrqh2w6G0+3hjmeYsgRbnINz+tAAo/OJJXm7+zsvr1S5rgnpE3ziAs8mnEuJkbZ
9sKk4DgVHhBAQU49m1vVwdNN1PatxbCx3Gs76kXa8POgyK5Ah418YrOy27TpIOUF
QZ8Sz44rP4CPiE4TUGUEx41n5H14EjV3FgNrVjEDpTP18ofLOkg0Q5UIczxgTq12
sdLE9pwvwIDuVIu5S+LBIf5DSkJwlo9MKcj+ThahFgH82wnmy4REXk2E6Lg/O5TD
t3ZCx8g80uz138zkNTRs5M/ig6SRuZCrwcxxeqwZogd2jTH1V+WhEMF9BZHOsSML
VyE7DJo+uL3nJw6PdG0Xc+9nY0mcG47DXHyUTrNSQZqhnCFx5R0r7ZqVPnOotkYD
nudwzDMlsjYFHMMTMt8WTgBlVGvbXB2E84R0Eh+RdEzi24/8l1iXNUqaNQ4OVKZE
WJnEx7xmqfn38HwDQohKboyYEYBpfmTpArsHFK5vIxRfYT69vwnyrGq71mPK4rd7
UpcFqnBNm161QbgBpCRoh/xoJ7ZM64sbw8yueRmHECHu2XEsrMbHwD+JtEq6l3Au
+iwcWHNm5UC8qh3Q0hS1d4swK9COOCEK2XodWKADs1u8gTsavlN54oqec0ZgkwDS
dyv9YALp/I3rOetrT6oOyPSIYtHoIW8D69W9zHPm8LXs92AYNLFxzdJBZOvC6Q9y
Jsis4WpmEwXxskGnFRGIP5onARcyOToGCsrvcgpt/1r3sh3hn9AUNB2BGlDr8e9G
jLqdk/TXbXtMA/ZTpFlQwBXC2D/GNN0G8WVwhTNVikHoy6WKnSpYd+AZALyk1kaw
yRQt4orlf/CgfxAVZalNQKZifNA3w6ViBGzr9uqAgdJnMPNO9lPcrLljTAj3Dht1
AVY2b6I+9wsbuWP2NOfmnT8DXOjPrP5JSqmQT0/XqTf87BTOzHkk+lLtrsDHdvfX
3LQ01+tosO5hnAcwNthDr/yYBre7FpouYhPHaVoEL9G6w5h7XJNTPMw3VQYoRTkm
4LK3B08FtypOT1CLjuUnQcTMh3Wcapiw7siAbMSuKm3W1ngKrSRSHskpHWkfchiK
PdkG6BzznRAGllKlDeqNmKNNDVf8nGmW0neLpBxSbEXkuc/H+BpcpAOYDxbeosoE
3AzQvFZ39LAW7avZydRRvXd8yWOtMV7JXOa2xS+r0KolFBY5Rfpspo3QeubIgIFJ
fdVrdLyNOL4q5XGxacKktezf9RWDGJrmxzAgGhpXKD9T8/PpsOwjZPvRgmWerDls
Lj125f5Ub4JPAb63Icch2/J4jzbFJJhQbYhuX4QIWkQeOTFeVztjTp7P3/s/ok2g
JuYpqoWkM3m+qYrTHNPlWHnZOIZHGpNfuaYA6wN6/0xieg5csQb0Msyf7SiKBkv7
BEI29tkleJpv0WVaNExevcmEwc61fVtj2aOZKEde650sP1I3HchMvBeHCCLGR6WT
2pdmdSPg/jJlazVDPOZQmEsXDUPtYw5BPRduo+i1CXyl71oJ6c8aKbpSZJo+YZTg
flhBZhb2iKeA/G6+PS1k9RoPyTblEQaH8hyoCZPsHom/zfbsVuTf8EwQGtEuDf2d
OdDl8nGJTYin1hptbSRRBPgXn2hzkLDeYff5vD/EvrJh/vpPWUjRNE/Q/Yw54ogX
pDu8rWnDq/qpaqlizVVWelDlxt2SBU5NGigail1/cpBbgCxECckJEIBEkd31Hkvg
sgGcB/Kj66sywbEG9aJMxLTf6zrKD3g9HHbqd68e53WjKde4LMDnAJLzuV9YNshS
vy9ja9nLxVbBaU9QS8h3zc+U2XLgsecEzaxmif7rHh8wMPddzjz3DmGyg4q6o7V3
ghgT3c6kBPrBzCo/8u1BBfNqGAVtJ+SQC28troBukHIeD9AN1BV/kZB4btTBCr0l
4dHqeh2Gzm0sCQNJ/upNcks3FOgr6ox5qgJSbFNnTmtgUfJAy2Du9XKqRvuO0lqD
zcQ3uHrHvDFE6+yEkzMKH+1lwDrneYztXOy/ZbHzstPHGY4g7sA6c7y/yRl98wcy
Lr9tQtw8PfngaGZVAi9qrbhdJKKpCaFgtyGjlV5KEHiWtyZ8Nwmd5WgpwzwQGOYw
wajdaCRgotdM/duGXSHSLgqImntbWwO9UBOmyoZpJVGQhNON/bd3abANII228ems
1+S57bmTKq1Nh2QAIKYhbAZIKDE5ujAqMcXCYg2N5yGgeFjz6YOpNNjzNsIjmtdd
u/o3HJaIhQpMS4YX2U+iR8JoL4joykkOnIvKm45Li6dyWJnXOkVbvSQeexCWlIOC
H7mJGZ3aJujTvfCPe+iODU/1pKw7OZIWLyryhyVhMGK5PXlU7sKUU0iYsoU8LsHZ
tCGlxDznWfl5pnMfhA72QHGSgriGhbpFpdEhq4nXBZ7jq+JEC/xKruepK99f7dL9
HJaraEFHiTN9/WZxSgk82K6TZ/so/Sx+qTlyt5dbAMB2HWwYGwzcBPAq8YNknaiO
/C/EfZnivmR5o942Qnk42p++ZPEY1cSEG+SIClbEgk1hPyNgxZBXNGp7Azxa1By5
xjIN1VKNjKmodYst7tIKKC8h+7QcC5O5tVSwcvudMRFHhww8Gg5xmnS6dDC68aTg
5OhAvvu9EqvcfVNKvgDaM3dXifJRoDgOkZ4vXzi/Y1BZr4TkCcgz0StKb/jlvdvm
yAjJBJjY4/IXbRssM61QzxPXnvAlHh43dAQlB3HM3kuWOGmAQLnuVPVmTQjw9fOT
Zim20olmlk3CQ4HE6kT0inx4JUsKG6vvb043arB1BKRXH7PhF7SLU1xXQ4tkj4EE
oyavLDLW9zfW/z2n4Nc9BCiUGrfvMdIrYl4/MNKBGMXr4DOS1q4sIKvsvtxsVIPN
Qu/SIdxqMQfdaXgrR++XMh87ikxzwrjd0ZpUkS7s+xBsR70RMHws5F0TamlAHndI
10zMWHTtfQly6EvNWqAxH4Uqzk/DDw1+VevQJYY/G38igwj4lLxtfmmwOpAl5E8F
2CJacHSUco66FZlA5dAt9eO7dMRHNNFt07TR3ZGUKRSMaW9dWl0QIWfBp5feIyjY
i5a6YME/27FAnyyNoayShHGYLfWrtzBHe9tmh1yE5cRcqKqHpGG+wBksiRKrDyso
JLHRZVO9090zNK7ZH3P4O0JdSfWeb3hA2rSk6shU5uA8pIFFf5xUZcahRCaAB5JZ
iPlJofmTp9q+9mCOleSdaEbu7V+oecmeu6E/zmCnMxeoCvDbpZFFZvzXGJ4pJTP4
83xHuCx6ZI8+G7QAeIWvRV21CEJBbpgV0AvhJEyq6HFXwpTib9tVEnY8cJHeFdfl
3zCTnwO4jZdGJy4N8hev2UdsHEaUgjt3dfnqCZebjZAtJjrVIsDeDAX+cPhDmN0n
VotkagKurbV2JfUcnDHCktKG7TeJokMYxLNGNxlsrJhfKYsYHvxgYnsyb2NIsXG0
L9qWMyuOWJTmYqXzmS0DukaGDLiw4h6SenTwOsGA5u9ukb2pyHUK/E/Cy8TG1ehI
mmZH/IaXibiJbOZ6HtmYw4nhTCOaM5I7hJUj/69AN2xXN3Cb5/HHzIqvEmyDINp/
7FJgu4Zlsd9lwf8dsrbZAVk1xu13XqWj34DphBF5qT2GyUqqW7RzNadnJsTv0TZF
g778srWwQ9wKmiaD6Lx4Pe4rWYL2qniY3iYEqQwUVbc0cCB42Co/xb+ZnehzgDyq
JzcTv7RiPyek+XW6cbmBoMfWC/zic+rbC00lbT7JFHguVAXoIJjZd6ZcYU2a73Iq
/Q/LIBK12AGKhD2YqEUbzOHUAfiElQd3Xatshn9QrdyldzqwOOSSvvhGz8KQfmOz
TyCFRZd5AgI/BtJOTEpRRsVkBpNSsT0pk7K1khtDt9gXUWTbcdzsMtVmGykGjgiO
Twwyr8dcPYJBE7T285i/5JNu1UF2MDlIikECwTI5AQyGUNpqZzgAoWcMHT/xBD0G
7rQwuQx4E18Wps40lZLb6/1GtIwG4ri/4p+qzaos7Mfua+AY/xEW9+fjgAb9BiR0
5qIjwAHpAZ6AmQ32cWwpmzWc8+zqvcX6poepMoFuMRJlQUfTu+ZhyTNn/dswA8oL
tJwPLJAYTte5tHK4/hkl+ngrB/8t1dk6fau0zzcvdUNb6ieJVf/EFbj2LzQ3i4Rv
ljI+jqeXeC3IMmuRwhankHmwQDfxn81qVGu3kxPVPYNEW0VC7Lju6fua4+uY2g4S
KDYStxPAukPkilFUraKIyQaF/DnWvXYEei63TtJ8+dJTQk2Ba1zZP5fFIludGsA2
PMslVGTFlEzODgqDc8OBREbHJWtlBAu6ZTrOrWvsJWGCvAJOJEEzNGGSwsNa2wPH
1CxsaroHVOSHEcW3FYPqDK+33pm9NNQoE9Wkzv3mrLMT4or90Fhc5uOnIr41x+Zu
rj9nzke2xCkW6Pkx62TQSEDX6OcD6+zTFQPQesf6baWd9nwvD1nRGaMKtmUR5Al+
gTml3za7hODG4+PghEfSUxYdUH1bxzvGquCeq7DKgwJFAYwTR3Ker1h1mQ6+uFCS
HFMS+Qu1+NgDGQrxWJaDzZXmxwSfmSNioZzAr7EzYvFjG3LqnIloNYCmDp/0aVBV
cYX53wVBEMSp5lAnApSG/WJFlcvV0UtsmgUN59M4mzu/OungPb7KALOMoNrUmmEX
elWM5XgOwdUqFJfjoGlzIv375roLRdSCYOvUaK1wupNsBu48xh/rP+u1xHfRxanE
jLhHrkgCE/7J8qcloWRGZHhaFIyIfLx1y2ziqhEMdAOIadwdoPOzd9HK7w6y2G1M
jfNs84oIJFQYgybJP3LhlPX/A0PFMqcXoEzKm6qp0lkeAG3Hicv3bSbC5A7y5fDE
S3LhteS3yHOsG+sze/vSve7AUD6UeknD32rvbAnrrQzntyGgJ3o1/ez686u1OvAm
HzLKmKeo1Sl2NaBZYkZ8hwfqcRzGZdTPrzO2vVk9r8btPmwRh4y1DXmBJ/L6BtCV
wJSulnDvc48jM3z3zkvQcFzJHwXc4n3m/DKdGMyhrJXroiuVv5o4HaCz2uKAONq8
lTLcXv72/Ntr7gIiyH+yey/J1Pl1AOKO95TALYr93eh1rBCSYjDNHEU51hcwn0Db
YTWSsEjmULSXzKeeKq/Yc6r777yALf9qtvY7/0MtF+AEt4uDbdsQWnXfYVNq4h0j
hXhPPiymAr2K8yamh4dUXw6G3UrPg3rK3fGLGCS/keR+Sddivm1g7d8IOUfRDG1C
p0DgMz5SRiy5JK2gCkWh0ZE4cu9fLuVGsh1W/BPT2Tma14N/iz93OqLYIaBWuHRi
oPb+4MQmoQcrO6FP4vkKpxBDjLASYXnrRWg4gKj9e0N08HqZnGo42xaWa54aylnF
qKQ0kUnsmYWsg5I6XUyE9MswPoWzIhsXTALaP6P3FigFTUWFHpn9PoMXRYAqhNb0
NGtz+xeV5FtYTJGTOScYOi/3Be39kCXlkuLrpGRaYjyjVwC/0LUPDwS3prTJYHTO
b4yj/0gDjPeqQBJxSeDrStBe/yGYeizCZNstPBYr1yJE0/kTxfYfLXminoucAEUU
mUgqDBeHKoLDa+Nnay9CY/BpdbieFpiX/IoER9k18qSq5lc+LaJS7yOQxBtpfA/U
JqvO/CXARbzh7JFjkjlWaKumAxzX2fh4WNXJz1JAw+qLV1Bdp0yNf+biEwzX384R
z+nncKu6I00tN9wZw0zJsLv8JWL2d2H9BP5AkrT5VJxUD8OFQ1NzJ7MtPeQcpKux
qozZj0nGS/fAMrM/aE2Bv/UcP9CxZxRsbYZsPBXhjo99Tw5XwGw5ktszT5md19Md
qZBYI6o1AMZXbHg1J3a83bN0hSq65opNpPGgIwLqq7dgFVxcWtvnL7B/TuZGVbAI
tx76i9RNPJvpkM5MP+KTurc2BLSoqhMfWa+75SI/ZBVWa7TUY1nA/W0uVFGjovJF
r7RDAQ4XCuOpFToYMpHcioWMT9WnSPXen6tH1hk7XZu637niFpWOjSreZmfudVeD
9L8TsZcXZyTxfGvpivzJB98pbM7ZB+EOCD8MuCrrXbWInAYECZsUrVt0JW1mXNSv
FfQ8moDU/x70IyUuzcQFUKNoxcE+npGd2stAPlbtZ9yD7aOpfecXDuQvCKpNXz0b
GeNwpuq1m/KAhoMX/dd+zvE78Rj0K46BHs4IxQxdt+M5aXzX/22bu3HNh6nbsU/w
OO3sCvcYKgvlKUnDzprER7QhDGIyTtx2AWMwPCLVw2GC4wIZb+7kv0L5NR3Nm/nr
Fmt5vi8Pmqx7ob+T0idnBUY35tGpMEGGP9yefCLU3HglNXlYPVC24T6oKiKdBoqX
xzq8qV4ofIybtZwH5NCteYbqCbV+U3rO2ynBvGxQiylJ0CQ4/PwY6VvFmPCXujQq
SaYxJreIAUqlNHJtcmAKRb13VT0IBXenqEHpkTTcsM8O02wOsntJBiQIFufgAfQg
Qa3GsOXn6o0qeWCFsO11rob1Ei6/61qCUgc0kt0zMuUmeHiLS6XY9OzHasMUUjXb
AtDWJU/6zhbG8hAUGmDIdfjoe0amLyb9sqfV5Bc8rFjTlped9RgGxPZmCghOMouO
2D2AQPZDoPrWn0hgPFM7GoGPHKCmKGqmQfN4l3reUTH6V2zzbhvE40FE4Iko2qCI
kPZdr1Ec3i5D+FdLElfF94jWOmhGSsRU5aanw8RnEwj7dwLkC5UFYEStF/qUvezs
AoCdcWVM61IPn0bspfxIvw52FSq++ty6g9snSK94mmdLylH1SoVmwpCHvg4VBT3W
pejN8DW9YqQx+F6iKwsM6dsEyETFTkyy9k52Bv0FWs57MrKul0xLFS7tNYXWuM+4
5z0NeTxG7BlDIBUxAA+nbTR/VV7jRPOTZVP8laUT1rWCydTOGom+l7jW5GOnusnS
F/GW5SGia+QfTkYO89o3CNyDB0NvEqlgB+qfSJxO/KOw8Cz4EQ3qzQ44ngSSb48u
7bSblXrwXfXKI2bV0t2GlogdWVdil0KhGDziK6wQeq4b8YnuMYejOaoLtzN6iDBi
iY+Pg926owWcMX4KXgnB7YJK+k8PdIbpKClnAJKwNy5/2XiPkYGUfMqLDMvtWjQ/
Zu3t2j/TUM3dZr7qiptQXGHjQ2f00SLAx/WTsJKVIR5hE2kbBWVWOwpN3XAfVm4u
OgGWgf22t/Bcm1jggMEqqRLObbFQU1spiw9LXwhziQWhT2ebQYBwc5rmKDjM+dDD
N4KQLPMq2+IGFgjGLv63m4RiIRJNkHa8+6hZYwTYsJ/ruJpFxq2b4aJFtkQcINCJ
SrTrBFyATj6gXg74FJAsHbQWnG5apLNyY82D51ElbUBX1It2AQQcQcw62/n9bWTC
o9rc2+HSBPyBIHH+w7tL5zbxTdMCFclo8Pyysu5psAqz6cNkHMCNdz34HVztnzQw
iz9idUUu2LY6DaCJtm+oVkKMDnX9zgRubkktN0lTMVzmtHbvV4D+TCNIA7oNYXBJ
+QlCc21TvV85OXDKDJYyuC1vjvHjBjTynIfNQXP62INOc8VL1hx16ZWocRiwjKwA
wkeMDpzv28dCKN0UwKI2De1fsTC9M9WuUW2ulMAkdZfekbbH4fb0aDrMF6D/CifI
lh8Ljeh7E3gERgKTd50xCETLsxiTF3Pzvk441vu0VemXBL6Yaq7EL4Qu+7okr+mg
pMi+EW3QuVPvBt34rQkZ9sFpZcONQ8O24Bbf+ZhqzvuW9R5jE4h8kv1SQ6SMvNR2
HgB5vkDdg4/DROzPIl4xuaACoiQ4FU3c35V4hEGASkoqRB2e9++pf2QG/Q9zg8dq
GeLvAHJvxnrANw3sHWMGMeXDVFz2CtT+hm7izPGyKY4eM5TDvx7ZO8v2kk/vjYFK
6tVE5JJaZWTJ7Oc2KoQeGtD7p7EaUYbe2O16NvVE31wDcYEP1djQ19SX1mHMHB2M
g//yTuTcXj1DhLRkLvyHTartM2SlCg/bJ32youEQcmtFdA1kAsSt1zDU3o+mpbLI
YIi3acCcgs/0cdHrttY3PundxpR3B0POgJxBTZapWT1xiPaY2giG8S44DZYIsdNg
MI4hkyMWqtlQ6wKtqYzDarFHJ6dSiY7kGCIr/ISQz96VVXgz2EGVtK3AI2dsyGhl
zSDzpoWj7xm2KhGUiOvXZtYU9zAk4bpGDfWul7MXo9yv+NL7GY56uz5YQW3NWFEk
UbFh8MmGmw05EWMESLiIgpbk6pMO5xQQeQXV2Htz/6zaVadMfSxf/AxH87XmAO3s
o0/zfFwX6GcU5yUFM5lKXgUg+xPEOQTEQOAL+IpfpSakFQSgIUbjL7d0nSlcfd4a
CBnl+sr3GRNZMaU9uAQNMc8Zy50N8P9G8f5aszJjz2eLGzrT3E+XmAWbcpEIitkd
sZdmf4fdRgT9cpkIzRJbRBeAyqTmv848BdSD5aCuihAnwnQgSIrAqZIFIiOiMNFz
1KzBelZNJzw2D9bvMWWHQ/KReQaFjnPjcxqoQnqFJSUXswUk1E224fudpbGfqHWX
ObRbjjhBjmkoCCC+ycVnHkUACqnZY7NHSn/6XdjIM9ESNAB56toi57CnM6WcBQLw
2zajZ5ZvokQYcOZh1m9FHp90G8tN91H5RnU+ATS8QsYtOSzzlJVj8Kg3WBY71f5X
DEL1pBo1zIICsEH5JEAbCKWzer3meLss353gM2XvQ6qSgYfcPMRlkAPpFSJhEtoM
sOVLW/azK1MJD5/mCIZAH1cWXKHalzOd1LuLiqZYjwFYDRvU+piweycnegyhOUO4
2oHM+Q4J4GDcFCYy5EuMpkj0UrFPEEFYFwnWYloXwHVa9UWeQ2BiP9ao5jZ64ZmC
DSjJMBTz8xwYclOzJ2XfUw6YpR9aeShlev86J+E26ozvBUTGE6SlFMnH2qq3wO6g
P0L7y0nrq8ycusIE/N/JwH5js/dVlKd8VFlSqqMQMJ6NvmS3m4uvtq8K4KgPu4+F
2rSyD/udjICoKgVSchCcnCWLDczTbtq0o+qBN2nO3gZk4bkQF+OdLLVkZjnagkxK
mPDxuDiuJu0yGHkIWnArJUjq/3Wk4Q5aCQK3mFuxteu/ZJfYN2mxw2coOmkrkGcS
0lyAm5OlhsazTDTGWIF7yPLs9o6vLvkdxqxw1UrVi1UrltC7cn5VnNmGv0O0Yj62
JkKU3rVMVHT0gfR8eDNWn8Z1HUKvWWfwrrjwW7UDlITeHYiZuaU1LvHwWokpwzgC
CbSdnAxUVl7cuyI8T/aRd1usLMXCN61YlU0AlRAD0702O2BVf3OPg3RXkNJmF8Qz
Amv9ndFIINejgaFzxAjWN2K7vsC8vynt8e1jySZQUvC3ba4q+S5epq9aN4tSHyRV
+DGqV1m1b/D9har17JuS86npNZwe+U2Zrimh2bdhb+E+meNxkD6TrdMtd/z6HUW7
CI7ZkO5BmtNQx5v1VeCyasFAbYyCyst1GMmbyw9LjxV3GYrWpOVW0v32frOBBo8Q
2ONEHm1YvKDJanm7BzARul1jT6Mkncvv4raH34za5MUVkuYaD9WX4gZB8j3G2LNI
CYm3/RnwnrG37tTf1t2ub7n8QaJ5ReReT+aTjF7W32bXicsdySoljXT39h27W5ub
lDrIo76APRdJmBvy0YwZax0NTNDZc7VfO3dKCbgIQomi4iQGXS3tN616R139yc0L
TxcDDwc5kGP0TBHORtGPZKHxBhAH+lzk2Kf1btze11qXjvl1oliZIH6wKfrj8RQn
XXtMFnY4XNMQfDCAvPDyauJGq7tsPYUnCNlgwKrL/Hd2Z7h6WC83s7oByPdzQrm2
2Bg9Ye1XTdJLrGKxYPxk4RPv9aAs+zgzV9TnrlFJMOW+WMIkJcBSj9aSnfSxq+6k
BXpAz7qiakvhwhVojaniAIXd9VY8WfGhCrd3qjaB45rtlgJqIWUwvp5VxxpPn4nh
YwunIBAut1Tqvd46UYmZcO60xtYKG9DixGcosm/t1Y5N7sXjqQg5A5ucYu8Pru3r
UBzzrf7T79t1bJTLHYHG2MGYJQbujiJATzX9Q869FmYX6L0O1H3+LhRAmaKAS/Fa
aeKo78ZhThZdWWeGr7aAKXTIGcjmUEV+SyWUxvTefAK/rXbW0pm2x6QjDf1G6e7d
a3Hl3YaYrm1miQ4WilEwBCAXx6saLMiCMUd8+BhbDeg3NLliTOUMU9ZvjDaWz6zP
6jTYDoE10ARtJcekQZGjNBL3G0yFiNvd9ur2KjyW4YCXFxljnYQo52pAuPjBKsWI
YKdFUaJJvt8rVmLIA9VL0pIgGdSjd2ocIE5c52KsXDBlxotum+BOc9vCsgK7AEfg
zwFueOAmt/+W8YCW2B/ENSNP9Fl5QSyigNO1Qk+e8YJT7oXtFQkM+oaKZcknwgxz
mXKX86gDWx/qhQmKITju1bQSdyKCXbUnpKSSY9lRVv4Y0utuXLzG+MBc2i00lYiy
O9TGkLkpLFogUILFq32XssF3G4v3FL9I6BL9N0bukEf74d/poZqJdAOCJWToiU8a
DUxXtnj8tsikrkTShxVif9TBBXwhNcvX4g2LFHkCqZeL2iEE84j/1+Zggy1aA0cP
+nEw/Q5Wc5a6HymHsgCD1jDCwNpUocaz65geFvqNGDeIEy12yAIAadoWAY2x0xBd
WvUErOQIH5KBx8ytKeGSk+j6oxWmIrRNWt83GtTjt4WwfjjL9beWtpJroC6WQJA0
MrRt8Z9yWx0MS8WvgvC5UvC+WbajwKQJIfAKorW4jtf2Xm10gtFvKt9NtkkyzTWi
DIDo71JDzYGYt/UFYp4coghm17yoL7YNoa/QLAY15Yo2B1glL0KY+sL4FfpdG8Pr
jbS8ApJqWIoCjYDh2NXNbDMewchovkoXnE/wQ49QqqfcMTds35/GSt6gL/Zb6qgG
QimM3pdWL90rjV2C9YO9f107ZaebNoLa/ujHBWAVL2f3IPUfe1Z8WKjml08iwOdB
ZUqjAMBn52BTdKtBXfvOUklKnRc0cFPKpWQrxSV+fyEwzc55rHpXiXp/wtS/EVTp
MxizZdQY/ck+eY2cYx6EcYpGda9f4W/XtmQxJzvWz/Fc9DsS6FWpxyVp5HVFMuKS
giH2btOBh/zzIfYa3Mli2yEMIdyzO7TabkJ7Tj4dWjSz4b2b5xaUuG+P4SIPM/lk
bQle+0o/DM62pAdD3fcj7eFSihWHxmKBqFVQLWOew94cDov8z2iHK+0jcgyeT79s
7WlLonh9nUS6lqx0F2pDuaY9tQSSd6RNC7nRYkXV+3uTvd2dMcVh/J75h4QM7Jsz
8BJJvk/uKzKLZl7YdwBPmuRvtM0blkhkoSBEE7iYGaTo8L4BirVM/Ka2LKOUL3/L
nOGQbsVb481M9GDPbAtXMOrGwY/51kvIuA+mWiTzWNHvk0CN5/EreqBfFpsVDfZ+
qi54eKFsWRx7at3pVHcH+iHfqYzgTKnooovidR6U/xuyR9szOhko51E5k9Eneigz
54cVSYA/rmY2jRupw7oMoOspIyoy0SKzLIFGuDbIFKHEDQgwnRCwt/btuV2QkgIi
WAMBAO8unF5ykcS85OeemkBzLQD+WFyRXX9l+BWM2KAQt0wejU9YkYQyDnTZaRSc
ONGA09Ld6IU8/+JVDmS2clx9LpoeUXr5Y1W1Jo4t/X62mX/cLlInpEfaqlt+iPG8
FqNfjHoy4TWvFwKrex6MW5QPTJc1hHR/yk5+gNT05Cp7STNdwcVZRtuPyXFcGCVN
IDCCAAgml425rv06o45v7zkyZQLueP8HfpbswJlA8kfpJmTWCZt/zpjsgtU5SANa
C2SOunaw/bKiJUaWZPY56b7/BNZAMH9Ku14wT724cMcXVXmfSyo88NisTC7NBuWn
mOUs1g0RHxeR2fkRPj7XMoSio2z8cNa76e/U28+v6EeRsD8YEg2ya2VRYqNYACId
zyuBrDdCj1x3Fk8hvyzR7ZJlocTcFm9Or46RXdb/alTp0WD9GU0865I1cl4qj7KX
LdqWtuR5XbO7t01Hv1zliO5lglgphIabdGUcBSUm1GyLID/ZXtaDzpp5X8jGLfnx
CMcEgRSVlM0sCHI5uGFxU0qDhaAs2ygisMqbbNvgP5toj8iRD4lqmceay++JhJbE
60Ou6oea8+XAwcCcO+av3xuV1dLme7Ar39rgZK+LiDadG45mR08zEwLb+aaldcFC
p0VrobKKWa3gfJ0Xo/doexVmt+0UXpvLjTZYjcDdLCsiV5614Zewt5vtBM3uQ9Uw
r5ABPH0/Vxat0TASHqmyhcL8F5YehJuDtTr4iJdhaL//HsoygxNiuGJMncn42ug7
hU/Of1z5CsWzu3NESfs56cxmuyu657nlsJ/MaWR4z0uEku4HD90ovt6h36vjLzDD
ynktQ/g2Cx7KnOWcgEiUtZ1T9q5mXf7Di+qBoWdlkHs/uemxF75jjJ7j8I9VVq55
QKVjUNvh+695vcuKzHQZRlCR7qSkKUw9ZeLgXkf841w4JW/qzRXkbRniOG/14yT4
iUXXLOGvBcnMSwuTbTo+hnKhJ8oW3A7TJHKtPBeHwuvIf4lVicqXPPSKfqyyeWRr
/lV4eSCLAOBR3KBIqDw0hyn1PQ82nUqA0jMYFrTIaAtM3rif6GzToWpPLrfJZxdP
j2nFa5m+wbMYujiwwvTFIatQxZiKCMPXh2WL7wDb5ud19fxDj8hnhr8p2PKIaizA
2IYGUWUelVVi84WmVNyVZ2zM2sUurKGAx+/oIMNHibd6xfLQcsmXL1SOh5DH5t+F
b3i/h+5unTszIXXafh8DH3uPsTh2QkieZuk5BcBiYeL534+WINMgJURoFH9mXK/B
qU18aWOwcvQSHQZALQ7n3ZZ9coTZW1kK8ZNLf+vefifEo9QInQB1XfrJaLxye/E3
dhIrxY/EZ78J9N0BUi25W+5YKsyWPNRo/FvMwc7F8m002HnohgoeKS33L6iB+WSy
EwvL1Jp8Wh2dP5dh7BEwDMMxyNl9w89glL7Bcf56Y+vJNq8mW4Kxj/NVcV8+Bpcm
ghmmNHgBq9lLfI+DrwvFAh42tFWxFE8kcVG+dBB1td5RGp+bYUkUzwRRxEkT+cCE
P6vDJBb4LoNyaAXm2mMJLGSZI9D7uXYBQ6OiJ1pZU+vd0IKh5OAuw5ExCi1nab2o
fYSPF9/wOLi/7qhWwBFr1l4bnVhmuq9wkbx2tHZ/0DDSBRWB0ai2KzsbLm+kK3mt
F7zhWzr0Nmya8C7rABnowBowwqWn6jJC+kJCNDRZ+fgmLRfTQWvQnqbTZDZQN9gN
dKu4dgaXrXah5cvMvmG+47elsqbr1ujVsk8uzndmMq/q14NcWt8Nb0Hqcs3DTE6t
bKFGoFW5Jmc8teLjjK2yvE1o1+rD1GTbafOK/veym5xpugyATm+MFWVRkVrf6kX0
IpdLt0CvcAJio8Bz5r0Eaa7YjIzi7Yo1OHWZnYtjjGqLZz6u1Y0TyRfkKkUGtLTX
DRrqzjcDh9NXa92fWoc8rvTD/jqI3rg3mFeKOEpq8/0zF9R+QkotpFoLKeOCnsOD
m0c1rvbA7XucvHzEURS06UjAlcSCE/dOhmfX7NYnnboeFEMK8CxEPpJ7G2HpOWi2
8hCai1PVCuc6AJoFB9ivD7GVr0rXA4zObdW19HXIJIQSdn1f9d4EntygKRHeCxzq
JSuoLzGOTnJFTY6nHO259nqxHnrS4Oa9poY204DcRQ9dqVQpYvEJ0YKoLPdMAVIO
FvoDttKAZaP7Q6T545pDDzeLObCqvkqrYOlRfSlfxbLAffTobjbrlTMqnyL1f2Nc
CFU2JC2iVWfk4n7w6veYAmbDs98e/etHIe8EjYcQcnQvlJ6R6IgLBWnBYh2slSWD
yhFXmuPwoiTXIalXRU06+90Lr3qp6jwaDGtDVRiCNxR95spR78BnFjvIw9X52qjr
uSXo8wYEankN0+ABXFJ5M1d++UaA0miottX0FtNHUI5Rdajqun5f5ANMJOzy8TOd
zFtlwCOEyT3DKUvQ7ueIDRMp1bcWaYVJJ3AHoeMC6ddCHfTMsyA4zOt/NvPasB82
2KWkGZbxiwmF5oggWkiz6+J9Cj8onAgB0bHrSL9TOZpHELVpRKaVAEXuIDUBq+mi
sWqtHmrL6lfZBGU+qQlPb+MNQQDxyT9VYIiIa82JGZpqzXH2BRK/HpABiQ/K99KI
s9MsIRUde18z4mpuXI0snmcl1LUhIQEwegLQEnlaJWSXmOFmeU9dKxj+130A2mQp
yw43YqQ3OLJBv7nPV5nufQ==
`protect END_PROTECTED
