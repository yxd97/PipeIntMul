`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mpTsqVm5k4NQJtBQhFVU2bMFeoY6U0+3EItE5mUnqO5uRX03eNFEDyHah4/JrNHD
LWPlngSphCjiRIHtjFccktt12/jgzoUQThbZg3A7GMGdNEG7AYhb3ebhkm5EptLh
ho5NARMPZqp8ptRMY0mXHsR4xtLdBJDnW7tyIGqC2n1Y2wy/1vMnGw2FNCjCI+ix
W4KX4eNvfvvcN7PHQX0BXcR404nxHI41RWHfcS1TFJnVQbYJkUkCX7sKkBoonIHU
SOQ0YrTnCjYuwyH513N2YRADXKnsAqYz+hZGNvkfQPtdTVlJ99NDTKuD+nGvHRso
Qstfd4KB1K+mmZgUogB223Y01JYkrqukpUrXBAjGdyAzQp0MZ6nfidFlGYCdG3V3
xDzB/vzMbzHzHQaZw1Gf09hFjOMuijfGMFZSuvCsFWVgpX+0s/e8YoibJzTtEdcJ
hDXXESmzgW0gqwHKfcVEdunZCXCUoKos0B66RwE7DnGV257n7tWz0AxnKg9B/KD9
15eW7QAUDeA5XeNl8MjzFNvENnmWcgGNHvPglyiCrjAEW1E8nt+hRx3UBbxnjt0z
z4S66fKE5lByq6cgBzm9e/HxUh9EvrTQmUxPhn0GD+5KSaItqO8pNPv2E8nzVRcc
LVPYnzx3WRDo2sEoademvRu71bl17opl7Yuuom6HBYnMtzMpiweaGAXBEnZaPyy+
51CyTCSK0aLzgifU6CidAN67FlcMrRtdxCMrxxnUA6JXbInQ9ml6oObopVUyyk7i
lscJ1ThmMEHvINMDaKbEvQ==
`protect END_PROTECTED
