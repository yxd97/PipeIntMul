`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMgAtT2dEOvPw9hjjDxQ1KuVO8pUXsrpZpb1Q3rHMrSKuBkXMJe5CN1SR5f5ZfFF
16iKFByop2Wi1PsFntw/92aCWNH0ohgd3YlxgAIDsEhNoNEw+YsKVcHiU1GdR9/K
dg7oIkESI9+PuMhqP0djrdNz5fdgRnchVV4/rcQPemnevmQBf6Wwbv6I9D3OxzuG
GlldCypA/8nsLvsPOpGEpDklww3K2H7Q1IcFeFIpwbBAajg796+H9T3+GCEWc1A+
1Cj7lAaz11jWhOXnqzUhdnYJE0ajdViyDizMEroklb1ll3raqB/JUrMGeEKGOo+m
VA6ItucFtlTfsc7LSThPxl440SEzAbBxO76LY0EZTx2fD0p0vPSyUGK3iRJYnq8X
uM1gH7WhvehwR0Htd5XR9rIawbo4cU7/XSnBLXldEr1J0cKHZO7cOYysLHKnM2aO
UEoim1Nq1WVtKiPavFShRT4jm+wo87m7BQI3bDCOzhs3O+pFiR6UE3JzZ7dUyv+K
FsCS80X+PZOASF7cdq1A0t/Zqw2d3t5qEjOTcR1UUVUK81fxVvV0QrgTI5Jc30FL
3Hl44OPs2AvRQ5Mk31QnhxKko7NBtrEurGrh0ysOhrSdngCY6euF4+9OKuWwo9l4
h2Xqc8GLaaHdZC1jPLftoHx4Pt7SXFW4Z0aYIUuFyM4dzML1/ZHxRXHgBw6jSNL2
ZQQubaSBGhiAZDIHeugo72HUHE0kGlpC20F6mpkijppS3AKzWXfPLPl+nUn6P/zM
aPdvhlwripxtvToYYbqJ0RDl9reI8DGvuqAjPcVFPJXy3IRp8BC3gD3ZJ6SI/gWa
DKC8+f76KN+l2sGFX/TEaphJDXCYX90thEbbBAdB2gm9ihzVQAcS6fHlT3kEd5X+
7OVN+tc0dvm/WGeKawSzlKw2xftTAUaLS6h3PlabhrgMglJRO6qtjhlPfN4ilw7z
2loPMsyaux6sxjOvTP59joXmzhybZoWJSxruSq6HU9ESVIyQUUcAezvoDlJbuKoH
ThGqqhn3xWIwFT4Avusg8wBZn64XXY0nrLmeHlnzweSqeNyEjp7500c0qmOr0tye
NxI3YGpRsKYKthfxMlROWoMjD4QyqAZMotqB18xJT85bhL6O1a0v0UeRNxxybWRO
xvw6edjwvLZKJ2V98cJKFzsurAmkmv/TnO75+pSzj3oODZ5TVznGLwCrsuXr3OW1
RhPAdDFf0gpw26zjU2fQpPjcl7CK8tOhZZ6kWFTNt50aMDSyBOYv16Ws6/Wb7xAx
JA5KKv8tzKKzNasfSzZZn56BmV/thQ0oSZ8d0H0r4BnsqNeIwVLaZ+5Fot83C5aX
50mwpFBF8mn+VxijLoQB4DkdjKkPZSC/xTa0DkK8Dplv6P70Zrj85P8Hcns0u03A
w/KniUZUmdqI3Oe720cOWBs6U1/urP54XY3PXYr8JFwXl9AXwtlUCtP5rnv/cgtT
GIK0O74hFbnXSIG0wemSz69YOnTu6qLteW9MpTxiz5Odwwz2ZKd32/rwJEI+C2LV
8Q66n+NMefQDlyjJUGTEZ3AGm2OMLl86GAm/pKgOS73hkJPZ595be571sIssHVE2
NGbG0M8zWpvcJQ/7+La3clr68w0YsdA/jw+6XLkS1Uv1WN+addyV50a7FDNEDRSl
UY3Phu0zJBQPn4d2fcG4BrVN63V0TFnQfEny649rmRbc6o/Bb82eKazsXekEYAzx
XudH9XI6li/jIGTkL/oVsDRVgb5abcfCKvPDz0AzJLArXanWZ8C1yGuaW3V9fV6g
DQ74aWJFWCbdSE9wAUVl187XSm9HcRGpVPQVoNyZHxdITmiSKl9unSpqrZrYZrDC
RgkcJFrkZ9c5opxS5MlW/SC7GxVzn5PNKc38pOz/2CFb/sMjG51YNw7wfiV4qUzA
rzZAkcK1cG46Fmy+EFWtEdrIOYWdc2qlpeCbICUgyJnp3/4pt+yR1dcw5XuuNVCi
1tbXMsMNy3JPCMkCKMoRNhzwsXIZtEug6HgyY3uk7sgZNOqOfzHfXb6yvFIWwH8/
EeFdLSb2qVVnzUpzJj093wuTS+cF3Y5iXhbEUIE7tXRL5C2clDef3IwxlJH8lvdf
5CxtP1DIngJyr7GvaAC2h6y5ornHIqUTbpUHQkZA7sYDiProS5Sk0l0mjIxeVrjT
2mWnLvVQf1JA7aZK41GWsl8/ZWgwkOn43WEa3GwUq//Pt54SClUP877e9yM3oYCM
378f0ZIOEwn5IyXTE9274z+0DlGJBgOCM7gYLtPyYfLL8JXIgdUf8Xlb5lLxoLfT
KuAYMW0AA550e5nY2bAJdNDYJniBFXP3KiEjAMrnvpBBVm2ftS2pi0VkfMWYbohN
j99emaUnGxOprM4uQVbtRkOHl0sR/wqMU5DzeeviH/qisWvP6cIf0OP+mHnUW7YB
vYjzNu+D9TZQl5jGiFKTSXUXqVLJmI0MzGnIr3/8vAxTqA/EucajtHFZtR+/S5lZ
gqu4GdgNtNs8KNiAQbj1Ut/6KYSe2zEESHS3OjDhfoOHMws5dxOtk/ayjRddcRku
fRbYnnVQbHUpwGDKELAOctekyNjFI4wKsRRhMLt2/Mz/lM9YcjhEvtwqJSUJLjmp
hIkBgl3uTg34a0o6KMRSUILw6SSYxhmy6TLuhnJOTwvEjtKdkdPsq+lZl6ZdQVrG
lDb82s5mGbHW/6wdc8Wh1D8qhAsKtZyGF3BBOPFEB/mEU5AsQjwJk8ImVOLGg0/z
/JAwoVT9YwSAJxENM2CRfrmHgjYDUR2g4gR0iKHNwpgWg5NQHTk6SQUaw4c+2iz5
oyS/soTYw1iKtZZujva/HBK2RnbuN0E5mhbKyXo+ASpdlR7AvsyV//9Xcem3MRLr
Hq73fHyLNeLy3zZrtV9WViGnreot6IXtw9idYXez7uzcnNf+nVi1nUREFiT7rugP
H1ii0RQaY1AcWQ7RRxGZOBjM5t7zm2lyW9qJdsAvR44AdB+Bg7ZxlZWRDCGi939n
dbe+znK0/RUqfse55JPZ1ZExHZLCLyhlZ4AhzqPhZfV81f9FezY7WCilqUtn6AiI
cxFWt37+HjIJNpYaSWoIbdwlXmuvYKil1USmC6kQNJCTojDEVnZEOX3SezPsEQa1
8TkQV7VNpw0qXO+2w0tc+A1ACe29s1oKWExPj8LiS7iW9xaL0QKohNp0MNLarxfO
HBDolbot8aLkCtYXymwjaCdBAC9PuNmADWTrausX0v3LZlm5wHGSyq8e9d173ZKu
IkT9dju5elP/ZZBB/WADzgw1eBV0eLzoT6gqoArM5XW3nzcVeyad9qCrceHi5oBp
mVCT86sPvdSmagrRMVVLeLywdUIGv1sV0oiyXG9CdJ8tKkCa8NehNCXNXpxc80+u
OlFDtkuGglFt285vtEL3UftPGS87XAvy+paYQZElaLMHaR38v7uaDbb6+YwnFaOL
cVQydTcOXWbPqmiArHqiViDlb3TgnwtUFl+Y6wtfs+wk0AXJfYblRvpt3lEffZcC
ygc7k7c4FNOP/BsuuHqzcQS81HBN3vtw+oQ0LECASF9q52P19oogq4il3ZNxibx2
HmEIm5Xj4J5ZG4qyrf4QqRgclCnBshgrrxXP/96dG0u/JB3I2+3LATfn62z5QaoD
CLoGelc7rPekSujcybYLkIUj72LOn56OyVsCzUNt8JS6JmbQHSqUD0525UIQeRpD
EhFr8m5zhVhRoyMY48UAYV1CkoMsG7hEcPkj07WsdJwiRZFEORa/Awt7iD5D6NCD
+aPZkxbQs6v9qtRe8U5lQqVaDtGmARzZqc9guh8fCy/Lzg09VyLu1jzv8xGEj/my
MdD/c8Bc306/qLsEz5r7okwoTypReN1zCQVI5UGsUeLs+scp1Yhi+14L0YB4Advj
5B6E6xhkL3ohilVREEFFu/KljdFPXOs41+wuxY252qwtt5rNlTxf21Ue2mAKFhLk
z9ce8IXBgyfyh4C1WEYcV1i+5th0XnslLog+C78NbT4ph78vg2tADwzUUyjrXM+3
Rmjw6R7ulG+UhNU2QgRs9gIhkVs5U5l02VFUGtMAPfpWqqr8TjkCBaZVMPBrogfn
1azB+4cNRE8+ZsIk5xMILQHYWrOXR1Tcrr6mxolvYYyygRNSvOAwYeZEF4iLAmYa
2OkutHX24G/fV7WSsup0jO8FmkQJpSGGQJlAc5M2gMwC0SvtRa2PVLjCSk7ThsP5
v+dSOG2jFqmzWDeK5egdQzBQt0/1Gd30zxmvelEF6FVRbPr/h18dyrJZUhXqqO+j
gzmkE7dRA2aGSfsW5ZrlIF4jQxpZrCXk5dUKTBMD5Y6a1nPpLbqaspaAusyGHSOa
NJSxtBdTPG0nrlucO4dQAZrVQgnBNRyb4qm9AygP3VDwrJhsOnzj4rTla0Zo/bZv
WbTvK0lA6hIOg1UFuDPXsRfvhrNLLi80iHlcEPqCYZukrcxICdyD5mL0JYnHsIb/
IR4+DnmGpQ+HVToi4tjUr7trmKc1Qsmok2o/JZ6rAmlkbeB/4yhb5vMYUQZbAE29
RkziIihu8NupzYj5dM7LzISlZDFigyQqfmUKG8vZXe+5I1XlmQrRCO7pUhkebdqM
eISsqpjPcaNM5kbBATZSOt5V4jCwvzok5NQkJL+70hW03gYr+7AW/k15V0m1o4SG
jO4/R+OCqEXwdkoxvXUVFPT0tFxPz8od06gS7p4cZhoovvOrVOSUsrpPKtFLUxM1
7sRvvKHDPNKI/L6w2bjUHd4b1KIbR0rnBucK4fdO89RdOZ3fjAP7Bhwb6eF1I5Cc
Os2S+0gTTmZktqRbjhkXYqauSwTMcKRZccqa5A3lYUe9oiAny6huK17BuTLP0pPj
IvmCTY5GcukSqIBGOGVxC9v1zOB6vMekV8LDf6cYAnJ6OQ1fcD3PZaoQf/fGYNsb
xM2vGUW9xjWRjjolIOuEmG262kczRAHratnoPlBIcg1M+t3+kLZYs86ZPooJCh5h
tn2iwfGi35H3HcmtjGrLMd/wLZ99sv+PhQYjlc7NIaO3AhVQGMX2YtG7YhZvxR6C
94BpSg+Bt0PFANLa+nJyFoAYpjeeJP4+YkB1WxkPQ3KRrxPP7il8lxeMp79dqOgw
K1agoGWJBLbkNKpQ9d7Q0nqB8kgWx86YMqTZvP8GnnEdY0RLBrfWSfMle6wzEDs+
d7kbf3xsQZyDbzmT/vJFl63ckcQb9UR230Q8qEvJhY8infXNNmXDeeuhr9Lwpduj
ycozkfwL9+wUsFo7YBeDbMQ0ohrDTFx7NgR8Ew1D+zAZM0qU0AfBrNaEjfZCJHwe
A2s3KDeuDZlq0qB6KyVfL65SEUwpHMEwRjhtIeUgFa/bqPD9730GnilHfheF3N7G
JbNK67Mc9i1CzhNGgrQKbGnqCyDexFlZRp2qJC58aSzzsWNCuz0TOQk+rWI8Iygr
P9ZV0mUQx9qIBSItU21/l+7uYWicq2xVDocx+J88wbxHcTiHv7hf7rR6S9mxlQQW
YqSf9KCjLr8heaNqbp4SYRd3jeXkuGgDO69eYqKWY19YsgMEL5Z0uYEVrZ4OXUiR
l7T/EcJsRrbfQIMMHvz2c9ZPdhf/SirQMwzwIKDDtAN0+9u2MzDIrlQrhFPlK32M
j66HHTrdLKK7O1ariPZjw13qbiNvo8gHCGC+KDBIom5h4XvGDhJEtc1kHeraiU3C
MsqaINsAIv3Ilt/NCJDd5i4656+Ik+bYrJO4iZbuzCW11AUNk4XZ7U5G7LSq9/Tx
Jyl7NN2F62ELl05vuTt8kmVqOEgWV39dRXHjgs9V99txusGcqgXJ78Vkkk/S8OIj
CmJvRRCWjKcSDaQA8B9/U1KREsjgRCg3O+y3cJuK4m7DAeKYgTcXeRa0OjhDqEwe
4fxiHfsEjxMwDPaMEwchZfkbB5tB3SjQSBr0qhTprFDQ4XvMmjHvC+3CkueN4v4N
XRhNR0UfQ+N6oc5qiAnGI8chdC47mNRS8oMepPLzGOkJTNWTVHRAK4zQRRoAkf1z
LHt7dKCkCwQuRpQ1bPyJzaNr0ki0A1CIbQydzWFSn/pI20pS8dCtLo3qtA4kBRP4
/NHsLf9Q8+vDDAkTrEb5oy5GhdVgzh/qCQ56ARY7Tu3CaaflcVh5m5Ov3a26Jqxg
kCJbmxkRP1Xs2iPpX19aX3HFXp96NNhwKU6XWS0w2eaIcPb8QKiE8sxq29CU4eKy
CtMUhjyqIXBV39N4xkB6o72EFGG7Q96YePhpy7BgOE0ZKLDfYmkFDh6xd3/Y9f+B
ypbxwZ+MilyH6gwPaShxnQNDpIA9kE0nfEk7SdmRmlaIYT50fbfwLgS0jcm3MFHe
zWWk+ngTM3nPnYGrsWYg8hB4Ud3Ptg4+MIPJTmXjHNV41zw+fwMlGtWaQK0kzTZ/
S/Alcntr9dLgzUIjJc7aGoKFoQbURO72spYGycfDwAsmPosXFHbWOUwfaKBqCMPw
5PyEIvx5FRKEboYdcGoQAIVuJTnMdV++f2G/Mj51ml1SAeSLYk/AzlV5RchSbRMw
PNc/fdHQA9g5sodEToetLd/o2fctAOR2pjt/p98yI3Q81lDYZM26YGnIklilgacX
MBcS0TFF5bjpiMb5jStWi3UcjF8W5N3ur4sBIkqsoV0xzldEk5g0ZOdZYTrm2/JN
Xb6clF2IVhqfrMj1dyvnKfLklCXmOXmp091/2P+ZMHLGIiP7gTM0w+nFCOg/1YEU
PY5fTr3vuBK6/0bRDmxy/To5CnFppZblBvIziIJIcmdAkFkYz0GfV0ICYO/R0Dah
ZrTx0D4ov+7ZPPvOItX8NDQNZ9VAjY53x6AI6Z+BiA2XVuoK0yRy4WGIxdG+x/FG
1//sqYpD6/9PxD4lgqVwcU+uTsS+Pc2ZcMsNf9IiHvLFguBxo2L0JTTguaCnmLvp
4CxdBoownRC4Z/Irkmfj1UD52zKnOx+RWXHwgaRsTivHCXv1+MiGtSeJIdyjXmK+
C+NYk5I9AzjPAgNrcE5tk1VQcDUdmclhctvp4HhxfhBPEv2ub9lMZYEhkw0Eot5D
LnxCALfPWD5QVmvtGiAiBCErL8cyvpMSW+NuMLBk7Jt0XzvfkukMJJ3d44XrfrVv
SSpc3Kodx4OxDH/rSAB0Y0PNHhb7oktfXnSlLqUH38Kh5xcYNalg3cBUM0ITVRig
vyXPXLDgv1VSu47CQv2KyRw+9SD0qxKok4SfJlmak4pYRhXV2f4NuFl69iHdglEW
Y9hRvzFhTJ7McaGmg9wCkzFTL4++FTimCcU+IssKXD9HftLhqcAUXvi9ty/c9856
NuW6clAXVYA6733zN0KJBU+D3Tpk9X08PKvP0JFsPoJGBuGA2eAh8rN4VS7I9/4+
jWFpWTeNpwyAqprR8XBakl/hDqyFvLIOhk0URzaNovZvGIXuNr4SwWYBcWNCWJes
XFus/wLV9xCng5ZRaJuRNJpu5+t1ffbWDkKrTpPTYBOR6jRvLOPzXJW9+6zbSeY2
QsUzTByyjtBQQxUeyGg/UKX7i7+Q+5Q6SrGS8MtFv8/bCInJnBcgkcrPMXWdMfLu
xWjt4bKJ4Mgu7X9aBymyjMjaszjl3/T7QAy+TZ7wY6KM51aUuawOa8Qn37cEqlBJ
skzzpPGWRATxNppCHgwRcK/eCDffJTl/c1UA3VLZauwjF0/JkW5g0JYPdSAxeK8o
EoBTfvurki6Ida+T7fxBabV651g9uizkwafPqCAuBh8jTDROBB2bf+vd0vVGbzNC
M1qsYEV98eQqs9L5qnalPHm8WR12/e7SmK9aBGH37C0MUZ/upFhryDBF4Xd2OyWm
cTvDRMm0ijQ1aWt0nB96xca+dnBEKmO/1kL5hpdn+lq/LBa5V+A39mz4eAjXC2bp
do20dVKKAFEQqloIiBBUc9aB6lS2HylsGzjFIjN5Acp6RO+Te0lDabpnQJEkIJ0b
013YqKYIAFMBbBsgn1xvmE0HI5DqZGDAqzQdv9E3VwlD9PUEPR0pM/Pla10MLFS2
SoQ7fneZkM1OHLtt1HREtGIZc39MoWi0iC9Sll8Pin4JZ8VkCRyA0/s1CqIJ5Q3C
wP91b6yWsZkTDHf981Vlc03j5MLErtosx7u9tgo02ANb4pN67UCUzMt2k0nJWN1x
oreQmZA/Xgx3KgUOSS3Ogxu5MMlgnYxX1Qh66eVyiXIR1lGQxloM76FYsJJ9fwzs
/WZx2bJnhxjIrFnJMqV+2h925ZX4VdWXE4/2gDDaCjAKwlL39A7ddq5a5QbdmkEg
hosxtxo5NA6O61EhfkwGUiBk6Md/gH/xNvRHoMBzGIr1Pfsv0pVUcQnrpl/nURQE
HvXYGCgYK0dLF0cigFGKZL34TQYcl+yW9r1IyGx+7EO3Qs1D4viu2kGV7ZDVvZzh
FbBTRC8WvMfwWrxWsT8rkJUAC28pXJzMYjWG4YkJF/xzjhBItDWWCUbNaewsHMs3
oWrKnluJtDFSw/MLRBPsgln3Srzd5XVeNwswf4jY1NAMDdmw5DGNLeFibEYHCEQV
xP867lmZ/0OT9tWSwOdOMH17A2C/8is3WswCdhCnY5Q+icPtllxzT4lDXTITcI0I
3Qnpc7wGquXf36jq3TydqDJJlr0EcEnLykRAlHFX69DxSb/JN0NHg6e91Ak6/i13
Acv5F8TqddpxeHPKoweJHmkBO2UTLdZwqKiZG1GFisKH62i55VmSCTqNPLrC8K8w
nitnID4UymFONvpsA+8bUW7UQR0bLdAEnADuw8tp+4eLtFoiqnXkW1mB1MNPbUXp
fCx0RV+uxq2ew5DpXa7pMx719sSLY6pge9lJu9/A+2iX7nZYkoyo+su0ZAD3MuFa
jmK+oJinrcN7KjI2KwgM6cSwWTYz0PmOTJlQ8UUE24wgoLI0uxRt+TcWDEh55z8N
/OagjlMMPZXKSv9i4G51a60TWPgROXMKbZze36rYCZ5GaTXnIpgPk3MBUmkabo5+
eGi4zJoGSwRhqMkV3yaLOG1D3G5+5qVY2lZ6Mip1ARbB7B1bMKY6eAGcZbM68TMb
XgZTnE3wmmVTIQcCe0fqrSM+IQ5rumQPiR5SncfujZbMR/KXVkoJaES2GFT0gzrb
gU5cpg5wcuqBm39I7nq4jTOeKvr47e0MjIt2VYEQ4s/s8TMg1gH1ZHjEd/nmoJay
gQavSxMKmc9W4hdfqfdjYHf8RZkfth8AB/aG/t/5muM+BX+QiIkt8ALBG8wheZ1I
yMNk9N3jH48lKAHd7AV+PHNeD20AldRp8fHHINGW8zq0VrOwQqCJ3SZXGZxS+eKe
ZQrMT3YYwf5grKtjQNBlBPuFVujh+geURPH2XfRVgQg6EmErCCz8+bjXLCI7E36F
H+3OVqHU4tiHXbpx3BtW3RyU31Zw8v+Y1EmMg+CgJ5cG7UPYjxoXxCO+jacDzdCt
I2kMPo/459BSU2mBDngb3wdKwg30gFG1IYdp22gx+7+57cv8pSxDSIt8N48KDKLr
3zzI6m59V7I33mRmANNgoYHe+1V3xD8+NSQYb1dBxc4z3WgvrhInyROuSieJwGq6
nrwt4v7j6vtqFs6jDz9+ywZUz7nqy416Cf+BSZmE7QpQsK2CYwXlRfc5ck9OtnoD
DCSvjHVmk8ZYZcYfQUItFNprtDqTjA8RPx6Xy5K2MrKIz3XrXfoki8luuepccTZd
1W4U6ckRRzI5YGQp2sx3cXwo0XtH6w0NYVrDwo2p8sQCeNheUTa5idXNtfmKGmAH
kbwE2Mu7L5jJW4iGDAOM3EQNglyJPEhN4NH4YEseD6+TfTNL84R8Q7tMS2mX57Xs
pflUfm5pD31cdZetnVw0u2U0HAXAtuWosq0n/zPouLVQqDoToUxw6OAdJAOfwJVj
`protect END_PROTECTED
