`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+z9rhkw+CmMQrNv1SAk/fw7bNP5ZNBEfpi5bkmtlxCiXaTXH6mr4VVrPNu1lBGu
Hgr7sh8udgoiC5Fbh3rE5RitxNng9BkNGlJoWrxfJQ3fCWThIRjOLl/C7ib0PBQz
pkfANmkkMiJ4R2wONgpGxdXMNUhlvt17tHUl7K9VgHP1b0nCdC/Ixcd/KHji4Hpe
99bKt2mlauYwreB3XxLBqr8QlD/Yocj/ye1lYRSTBCcLI+p8AM+x1POs3DZaF9Pg
Kjb5mDAz94HIHvTUjAYfVh/DXEHRawDHpmOT89hygkUM8NYD+m5jO9MRxBkwxu1t
l87c4CW/9RUjYbr7v8e4o7F0Kl8Dh1b/z1Qsxgn58pHMcuzPb2YaJ6GguFeHf6nD
gCeTpeXFOv4maZY/yc0Vc0OeD0OqqaMqzO3g0TbZVEDzX9/CtEV2tMwvmMejQ03O
Fm2DKlFr0zVkuuRF9r2n1IVkIdhYAllExE1MJo570uvGIpx2x5lBLRSLD9PC585k
vFLv2AaO5JaqRQTTJILU2TWi3oIqnDkMGFQuFAMTPjWgrySjmkBkAF5/Q6WzR12J
Hp3EAUQS9Rh7FNK4DltCpgl3GFT/6B9svniAQx/WRiCNalz/evgQzRFZG3bzmDeE
gDHi8AJTPDF+D9Eo8P9wYQ==
`protect END_PROTECTED
