`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sm/5vhbAw4CIdDbUowDu6OV12fCcC8zBudDsfiSltkIGzJH9Uv5hzXgNFbwzACbS
YNB5iKuvlTCkTY2G1orbvH+PnU6HbVc1gdk87wcJsX28ARngO1Dxszh0yRPzAf1E
wYKeNRybbq8Wx3VWHXxZbo5d5MDvCx13g1VkaZjnY+Ui3tTG8XchQuckCMotLx7f
AaqFAvzsPIVnBDULqWWWQHB9gbqkaMzJqbvzE3zi3l281aD3McY6xhnqfv3qwElN
qyqHC0+HrZ5ljCXfyROtsW+GY8WsN8hm9P4CvuPgdqZPLupJGb0B3O94xPemCUsW
Ot5dxaEqre7UYt2ZYRyMI9maY1t0GASRyM26hQHnC0oyPlXousTq6nPYAWlJanvg
ciVNbP1Llqf9FZ53e+iPSg==
`protect END_PROTECTED
