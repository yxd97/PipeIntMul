`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQC2VqdzRBDf1xm2vdaXDaI770gfIMzOT8jjtxMDx/gUtnMYAieyAaUwwKMGKW2d
NJpjxuzgP7TEv/s9BZZ4JbTf0fojR0fHqclMV8pdeuf8l0rOK+0BA/6MKYZwdCE0
uISC3SYONSkmrjjJSQLy1PZFP9iq6J7xHEwKZYgX7h6g056RU7Jo9cwgCKdDe151
a+As4VYwUNNKs4CMNfSb5KMKhvLcI3rOBv0WXRZMGbzGHvMQALhC4qavvtvVdvoZ
WGMaYxpSIgFcN7vsjMoOUlLD1+slYhn1qF7ybzKQFhmWQiVnUSFdtix5g/p8DkYL
AeB+BwSkoFYOexXQIgQLME9vWn88e5p72gaMVhqAZKLoGrCnqHARGEHRhwsH4adm
XeIj66Zl1dpRj3NcnM/XWLf3xiM3IIltvaJwGUEBBqqCVvSyD+3L9stV06K1C4BD
DbTKoVhuC2SeG/NTj/OPCoMbaaAk/H3kRj2HP64AJXIon3/xDFLVxxWlQI0YY8sp
kZs95BT+HJ/8ZAQa9lVlJmRB/Iit0ny92VoORwD10Cg=
`protect END_PROTECTED
