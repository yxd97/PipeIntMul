`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/tTypU6jpJrjxD2zp45geGxFhvwhDCK2dZQfxs9dCSRurIas4tpzB6CLQsbSu+X
jROgD3bBr47uBpPU1KtJ85qLY3CeceKTrQrbKzCBtvLvWHYLkHc36psp7OhBp8K2
qmn24IHo9NkQtQbx0nf66/HJG4FQfqNk6HTEgt89tP5OdBlhN39TQkVvKOarVz2+
DN+CrdJh5YFEo+viaxZoE1MWohoAWfvR046UG4hP9mnBFJDurrFInCagbZKMgJT9
MCK1UZMOTvEzv0ZSTV9siDSF/Vzfp1XPQyz/6Cwg3Eqxy/mxWXyhHYgOLcaCg1xn
E3Yi7IBqJTtEsaeMVrQpnUSPX5nAQUg3RWXK2UiP8ZR/LRbcdxczC2Wiw6hpCslp
XEM2CPw9Dz2e/PYd9lRC5QRTucneenhp5IjCJiUZfXg=
`protect END_PROTECTED
