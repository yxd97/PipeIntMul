`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WwntbCbZRVnjb2sy6AMVE6HRhIfcVDWPrYDz0hg+RbkvoT4yZN0vNUDFZhfltoZz
a+Gc7LUjZiJLcYjdGLzDwqHVL9D+4xgAkvWTRGnUu9Gfla9qM2bteujwphn6X3Hb
ci1MZG/SF3J+PZQlzt0MvkpGstldBWoqeT/CVAgk1THiAM9vyeLff1SNgfz1jh0R
7GZ0/A2nHOe6hwVei31BjKbYGRC+jSexBZRb63eCfoVJbPi3SLZGKm6uDiGLxwBE
5/99/OQ2PqsNKzngdY24+9h+qUbUj2Rk/3+qX/FkjFIh6vT5hp9fpaRWjrgMoj/h
SBUYU3OL858tolnkGFG+M+oHVZXHdU2O78zZuuUW17o/cUiYMf5JjNGDECK4GGf0
22X3iop6LiGeVZPkFZr2N/gWRUwQTzKuPdLqEXIm16ECzlYTqzKb286r0mzs5xt5
ENBQkrCJH53MsMM6wUTXHEHQRTEeUeXz4AJOkQK6XXQYR7mYx2EzXSAdVk6XUjcz
3JN2pqoxxKidKN4p67t6hWQLjQwIg2bAl7jeDuysqUI0OXcmL/C2gGyy3SXRcfN7
ufBLOKDMG0FSDGvemmvkJd6A+HbyYWTG/uv0ybYpClaaM/6AXg6yG+aHTYgvcHLi
/7ynZH4Ch6TM0agCHUNh2/LTMVe/h+fi5kwTU82fIusxROxh3VZ5MqhQvaPaCgti
faN2z3Xr2Tb0JIHETHCphzhdagwyTpnW4sCBWmXIOVN7UcBWUCQs8ejqdNBBWfGd
3Q4cswtX5mkIenowYqfszootJLpkvBtxMkvFgY+dWYD9dt8cf6yFTRFKUTavmJdO
lcaHnG64ktLOVLB2gibpJ6/mTYYlHfnYCEpkRGIsnJhkAGa4dG5YF/PER2wNQ8Ix
LGOdoWfipX3nPEKdWhdyOmD3oa2Ej258lvZ8gs+l9tSpnzyEKKaWf/jJi6SLw4ZR
YnBa+dmkEBtZ7LKOlkzuDeHNh4zfUCnWn4kkSx/k2hvyz2QNRF91zOrApyZBs3zj
LSdgTeTW8GaXYZb0cnFW63GMIGpL/1fnhOkdPCHJu7NBjLSSgddCA3kcxPKdFIDn
vSUGL0FPq1o++rVXUhmqoW6QBjnPXDWaSKRGQOyDYYwWtWwE/aFLtwup7WnZ0L5W
3tWE3GzOaIMcMTho3+SVdyjEDtrZAEoccnrzOxlMaBQIC+77+r9uVJLs9cIB/m19
i8sCS6nNVR1EcJ24yVqVQ1D59+I+GJWctmr2dl7g9eq+AG+T0xrAr0MFJb7hP+wV
vds980lgQk5bZTYSUQBTnnIAkPSbCQZLwaPXjt+7z7mYDoWYr137cvg88qMkZEh1
arl/sjK9xlYybjdInxC5WejkJSzdg1IlqIasCv1Jc7jBKLsWCjq5g+xzLlCiAeYx
3v2dXj1k/sVPn/29igQsibKHWPlhWoSKvDWU4JDAWimGvoJrAQyDKaPQEfilEdPs
`protect END_PROTECTED
