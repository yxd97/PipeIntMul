`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
llx/CXkqr5VBvOGGzAAhtfjZ3/c1rBOhggESEXEo7FoSxh0jlpeCMYsqdLoFIpul
T8EjOwx6mmVVM4znNRfVyqoVuv6hO1AXCcTWaLqANpZLbHXirCXZQ8ZTlQ9BTr75
HkGSM14mXcswY0hzCQRPsLNNkpwkxDGsa9IAgu2oSFVDUJwDJlstRXH4+meD9In3
49DC39LImSpoizGZ1csE/HV6RLi8tpvJwlepl76NJZihqH5+NT5U0NQ6qIAuh6nd
9Oz2EWpooKJoMZ9Ag7JQbAUSKy2M6gGKcI998dhIWQtyKjVtSK1tU1AbT7gl2/Zh
zQrtzVSbAm3DFKbW9R32r/0SOFloh7XyXUeOC03HCz3cV5L3NYvDAI6BSN/8kPUZ
uB5m9ITvIO/Scu0Aa1MX6heZAG68p/Iy83NemYOcR14YkfY1mJ5+S7t7e54Rt2Sb
MWS8Oz9FGccj553eqU+KVRiOOatdFfOf+Ybw6hm3zRHRIqbFu6ehtC3Z+3V5s4+e
TrbY6amgCrY0wDDvBLxKbT/akxdxAnHkYTxDl2FcLG8boe8PBZxuTbk4mfB3YI8d
w0LYFZAKWkBs1Y+FIyWHOoFesmkbGwWppNsSA+37hNo=
`protect END_PROTECTED
