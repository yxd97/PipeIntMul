`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LovJdxKAAZlgR75QJv5UWiF6Z+sbg23pCP/kOVfCosjDWMrPHHEW9HJLnsx4YL56
4Fu3U0nyQJogJqF/jo1l0EOfLr3EkDy12soviaTWXYa3AN0z5xFNL2pXg11UBgO1
eHzh8qBCqRosyiVwAO0UxhbEz5t1m3LfCHQmYURRc3EfxU+UOioA3NvpulDpXo3M
lXWd15Gs1dAqWI3bnbkASatP8Z2OT4CShHNnzRDHPEEn1sqB1XJP9YpzW9+omokV
oo7lkeAG2jo5gHa7v6UkCmm+mS1cqGYxRrnuorQfcAoaDdvT2YnQEQvQoBzhiRgz
CuCfUL7sQdsTExfwMQEv1t0LY1f1lV5T27ZankVib+o3tP6nbmeOaBN4EVQmsVV6
G5bZTzWrAyZ8WXR/rstuCmb1hkRFFzQZi8kFP/Zl6wvP7dn11psPFa8hCepaa9tP
lKXg/fJQHrF/3CIcNgX4r1qoU5OsZ1MtM2iAmMHGthOZ+3BLMJUe99uY/71L4amM
huF5uBXGMiHtplzBPXCJmSsx7wp8mV1iEqPa8mJhXL36Y4HQJE89kNVF1/DzE/gK
o6XSLKld4K00YZFF62DU+Tsd8khYxfeuz88obFV938KxHbc72kOIbAGf+F1Al3hx
zIKXEY3Ob98kOipKeK9IFnrSmlHdRpwBgaCoMgH/0eOvevW85NPizkyIF/seYyKp
ctrEhP3Z9k41NhCMSsJIMcxqbBkv+uYvfVCzPU7DuFT8GdGM+z/zYMa2nhAD0Vnv
UHU011mI9PVK2Yo9L3KKloGhdXx52fMb61zF/13niPQGlNKQYiJtz1WFcVhl1X3l
XOWs6/2rhnXgh31AkXnLo6NZqu0oazfI+RmlnBvRJy3THKATFvaQHhy4iCGhDax6
`protect END_PROTECTED
