`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vgYzI9kgPwMWkV/ZWAE/KdzYqlLV15VzLIEYWFksRLsMDzQzxh1Ly8Dv7zdqejvD
FKxvRuparPfXVWc3oaQF0hnEye915CnZm7CphbZvOt6lF/kJ7Fohd66fqGs/UV3l
NQaB3ecjcXNQxxkfq63YiSVvxeeNu2ehiC0P3jUS8fMrZ4Iq+/sLklZnxLe3njwU
o1DqfFrfSs+HARbcEr/bbvP8T0PnA5eDBvQvNRyZU2oIqEWLRSpw9sALvfYvRBEu
2q8QlzANGvQ30wga9H00HpOhRkTRt3Q8DJXCMevCrkRYbcxhblczhspfa42/4wLM
PW+1SuJqVkAfgHfw6C8QenjvBiBIU8m8kr0lY1mMbDkubDOia4+f9Q4EVo/z2VAb
fHbQI/BLSgsrI6388MlEw7Ejv59O+CWBkZGbl1uSLeM=
`protect END_PROTECTED
