`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FmO+cPQb1tgvuZJcfdXd/zZU4etwdhob5gy/4h1ov8DgLQLxGH40UiF8zoIt3xty
Pjh1xnkHA/5VllSQgYTPuQMtmnA+gtQMZVof3FGEpMX8rPyWKTEM3Ng3xoe+FlkA
hp+QEcYYXVhxZoFDLQRiAeK6Tup7BP3WTeJmHSgUDZAP0sBwLXHDQmhXtezXcmtu
L49nEJwb2Lxh04egxAav3L74NfVMw5StzpVGrQ1hhExy7ChpfaV/ax/lIZ+5WONz
8IlytMaWOgzKgElCeVkZbiWRUH8+++m3VDYj+09ucOoNeVATZ0fLrnjiuLOx/c7P
Zrm4x2egePTH8yHm5fKkOZ0XVbLOGk8a5kZc6GrecadRyMWdbvVs0Z3mjtfYi5CG
A8whMNgaR6hsZiJTBwNyEPC/x1TJNpMkrR6fZFGYriasIlfOmp+Q3E43Vasb6as1
uaMagkFBdbjxN1DSfOf7p4dz67FeGay/OEgvS7kSklwYni42S6g2tXI6FPn/iTea
heA61TnQZHQ90mXXqmId9pSGYQ9dUzMafSZA22sExMk=
`protect END_PROTECTED
