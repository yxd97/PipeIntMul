`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xgLef+uFlFpXb44nT7NiaUlGWVdyEXGJ05ggC8ytX1i9333Rl9fNGka3AGW5tRI5
dDwEDpHNuHTzqwT6xXYoun0kyfPssrrFAnr2rE4JDObrVcs0QXkgXYU/PVOFfCgy
sWd676e0H7V0Ww9Gf//tuBDPJCX+/P2s3S8lxZubbhtCyoElDi3vb6poDLJ0dKNs
Mn7UZTzL15hnZWMdYrkESOoJTv0qvuvpU/1ECey4TJ5hUDo2BBP+oGznOfNQjHlk
w95IT/9D2Jl+gyDN9zKW19L3ZVH+8BRx3pnVpvBx08SkCgS7iToU/5kQVilbyT7v
wutyqduK7jGIe+Xzwspfi1HZtDdJRh6QFunaQwxpYfVpvnQR/Kv3EEo0MPIOu9ZU
Bdv5Grrcfjvf3QaGcuM3zbQUELuvUeKhy0+UTrU1plNs8R0gn+eex6nO5sWVRsyQ
`protect END_PROTECTED
