`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6ZMIXjiaBRuYXhhoD8fALz59SJVJ4QwLriDkPEqjlUXmYCXeqQ+MlQyBg62OSDR
HAxU26m6/X1xGLeJ4OdIOacPrdTenGCzSw7dG2arvEyDYy57RNUECTsRuPqattC/
ihf1Ggm7Dgz0SzrfhEhSO+gstOSCQkIkGErn/SGaLUBiHeYTshz9fA20CnYLqXxS
230/7i38GeeGhUPLTW2Lu3ZIKQMreYBz83UaY4usoP3k4QaUWM0eM3zTRqp+j0Z8
flXmtsDyfSgLZSyrwTneM+Sg2aKjDq1vj+kE50QX+NlSLY1SMI/bajCgo+bqDCJB
Td/KutVODOeZAw+r1f00jGLPMG/kpZuvbUIORd4bWIweXJy3hZxamAYhOmXAEoMv
tQBncVJ/7cN7LHlB+i5YKI/C3E9ry2Xo7D4+5AHJYrybqq/Idii4WE+VpSN+lIe7
fc5YHzbi1rUEciAIUwALBQ8Q4CIhTmWYQc8IrvMB4CM8WGbN9OhVOTl/fAdhb9aB
Q961ltvtjQomlis9m4H2nTbZuzJ9Nkuxt6r52M5eLj3SryGvepTqzdI7zP4s58iI
D0VlXqvcsShWgg7AfUl1TzqR2tg4i2TaoNKh96pjRoIPBHJ6ro16HCQKL+yJFVXA
wEv5bM2UNzLVJ6UifMp2bLsHHAFqpssP+pGSbE3iAlElJhhHY2etFukn+btP9qrt
QO8ybbOKhs0dh6GZOOurCyleY3axoqPAwb5eOMzVx6QT3+BxzOhYbHOnak83Ep+g
8P2WEDj58E3WBRG2uUzb+p2Sl38DTvMPtoIBLFQjVf9ApJrwGh8QJDxL8e46c+FR
nrMp0v1R4wKTaoOh5tqMR/Pz5W+SAgUNUbeNhGWnedAz3IPmAQn3g6/O8iBCgPcD
Bn6Uv7w+DdVD6KG8CnwcZw03s3kcFhM6V/IBftIpwWjFC8JNzyxZgxPjgDYWtewh
NabVTIKdlXgWG+LhER+Cy1GvuZrZYoMRHObfcll8g3zfCDU6KDJWjqRlRvIdxsGH
TMknftmOfIXvN/Z1OOpIGm4YU8IRZ0zOosVLklssBpkSX0v8lExECJQo1QURsrOw
O5TLoMy/XOB8NTkF5eXuq7n8Ujse+ZVB5vdKkL3w1YuFI5XTpjhD7bqPz8VsIGj6
aostFDWpwR3qH3QG82w7kya/2Vqlv1JTRgoAFH1MZcgpvMoojUQqsaEzpeWa3Ygf
zZ0Np8jI8sU8tJQk+lLawK2Qg50ijwLWkZtSDinSlqXesLfSwDvBALLIPb9jb7zQ
`protect END_PROTECTED
