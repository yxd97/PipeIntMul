`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPmllTaRYKauuACviNo85kris6I6ElJVjh3w7yyuGi8EeQM035mrhrjftkPsJp38
VWrhDs8CZyQUj+qyjjcqWXOD5ACQElRUC6FFfX6d5zFFrwID6ppCoczWXXsF0Hyf
FeDkbfmV9awv4SDCLBQObjEwGsD0THbfLxT4Rxd2bTSpyQRmruQFxkugnfV2KT+Q
BTG557lffVU8gY5zG+Z4R1oee4vh9rPFt2lY6LUUsC7z9yN01DfxzCwJe2+bJUo5
jDadZiHzcNT0a20NLdm6mKS9DeT93STjV2LZYh7NkuzY7tsgVifUGh+gOVFsx0Fg
NP/mEVTb7ARAbVz6dzS1zyYqCiCccoCOQqs0GJbe2wFEaZ2KNT0COe2Y8f118AUG
vSb/lYuBmLmKHYQpdp3yRZFmKXtyBjJlELttsNQu+wgpF8p8Sfg6nszU0uDEH/GW
/v63HVfi8rZT8mAdkGnYPKjg2fws0B5uU82WQAaqqLdFtpltz1/LBfRchHSPa/RB
t/fqYOBnJKoAXriz3NPsrVvUiX8/nxDP1I3r03h15mNtyqJbMlgMQMxmqmeBe2Na
gHBdGX4I9/04klTN8T1IIEJhdO5fJ+Aoc6ZEJ3LdUHWQTq4yx2oHXHALC6ZwILsv
7UU0/SevgS9Dm1YQ+fqmgg29gXG/K3XSwkKkzdTzB1lDzf+t7BrKiB7NweRwHW7q
SazOhKFFJTzq3UD7sxeFe71BUHvjuRcWzAqxyXL8xvEWMgFtx1mmCGcp6evNGlkz
nDLAmSYf0rZ4h9FzqXl5Fu0zRJY3gA2qA5B89T4EBwGdBOEhZ3XobnBUVbqNs7S/
jmOAG/Mt33QzkkweG25jxGiAUNBRGJYS6Dxueo5mi6xxzsIc3HVp6LgtbRehKU6Q
0JFIJ4EmNcFCT4L1jGqxvtGbf77uMgnLWtUMb0SNfb3qxIasLb13VdvvgPliJCoW
40h5CaZUtOEvWh0fvmtFPd0th7TB23Gu973aaJapODnM9Nl5IPW9B+rEbqn9llhz
G4oN70E2jtciqKYGRGkvBFZoMxnO6HPfszWw2AuH+mgi5iorQJiaXdbKhFce4ijA
A1wXhKxnAEw01UsYIqRH4q3Xcp7bqpYANUNDoAXvD8BreroYKbPEvP0I4X7npBQl
FR87+BWVbE8FeCWDGPNJSo8nyAWuRxBYtA+cRtrfQ4PRa4VqeFd1g9fVFSDeM0ei
sBO/v2l/zLQNdV+0DOwrFTHmf9MkxTOykONxKY80piOlQ1SSjG6Tbo44Lie5L8wE
9JfHzlHVccwj9RR+WwWETlBRbrjQ2LTLGHx1xFsFMttWh3GdtI3mQ9e3f+dlmRVz
8NyJnrvcaJpbyDTMB8JQQNI762Ty4UXe24fcl9Z/NaH6RZDFh0nIbm1zDN4TSzmk
TcKpM0YfUap7VXseagSiPQ4FZ3OR2yqETswsSYs2RO0Ie/tpz5lgn1ujyA1lzsH1
u5x4WYU8WSSRzwY9Vnecirg3kyEbTBsVJs6vf9PwlVsFmRbjmZk9/go6bKxnnXzp
auNCu8OgRMiUB+Org40cyvKHH+eX/OzMWvEbBzyl4N8Fn3U+BvaorXuDetznd/Ws
ZeXQW/pO7wdFwywuXMJ5WRMI04SXuwtwDlux3r6G3gdk+ZaglDlWdZlRZBsJM9qK
j+/Ckf8v4qYUcZwjdNmavLI7Fs7Kp5No0g8kKQ5hY6fWa6e0fMqJKTYdyVT7rOS/
N5RyE4qK1np53AWfD/YwT1W/ylpEHBz541h/PiGtCsHc7b/IWPp99bDllKdqaM8E
JRNQXZQi7TXeMP+5X21PthvyOQElIdAc/EYmCxweuugG/vLZHkwJc/BF9f9eTEAO
7GUE/RrNkBabsS3bEXFqXjICnqcH1pKBs2IXRkB2DImcEmpZvezMnDPLynrCHRW0
j4EtLocoqwJg/5IvssVTDwdjzfnezXPZAXADKeWs8vN7FGkGLwZpzNZY8itdTphg
wiTNyRliv5h5XEnQ8FoZxOsSgcEem1/9xCsVO5+vLQd7BB1AZpOusWAlxJq8P2kq
QXUOWAdHPeWJTLqiOv2jYetyi0qVzJ24rmpf15zhCxDV0rEI2k8iX76GOkBGXiGr
UmlHNrAY4F3mh9Gq5HpkkulBjvtIDBP0uWeJt5Z0U9xrLLbqt9Zh1vISlncRF6/I
LAc9TOQ5O/LGlxR/+MHg0w==
`protect END_PROTECTED
