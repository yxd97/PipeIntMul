`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VM0CzBAhppT9+Qxh6ccGMQz/a4gxO1tzGEOIaXH80Lr1JaqI4IR2GRaub7UXlPRu
EPqDve9HytAHQS9H7emQLBfVKgqA3QK9RwKNBr2m/bN2zi8yyAr+3mZ/XNUaEW88
aFvbwFoUcB1VtKv107OyKyN/ui7EPPOMwLSPXcgb6BdULF8c3/m1X0wk6UywRWsF
e0H82VhdQ7dqAeZVLOwocdX90SCjUoJBdWmZCO9N+9s6H+WTKnroQCVI61VNOFcF
WOY5cdfyMxNxv6t/MEYtPxMj4KooTg1lYSifk705BgZtKqyrUBAZpN1AM1ij3ljQ
QNJCJDicLE/8w+HovGax0KkBiU0ugvrFZyGe3WAsyqxDnX0lgCVklpouhXQI4J8A
Ou+NkERNHQXDK+SP+0b7yE8Xrfn/i+cq0zOW0x8P81QXR7ReUHomMD9p/OuuNfoS
O7K91adAywFFa831+KxJ+w==
`protect END_PROTECTED
