`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcIsZw2ZMrmV9cCpinAWtJrULLMP7l6/mLeY18ocQAZ5qjPNhpeZxL84xc9WSvbb
+6fA5MKVZ7QXiN0kp8mYL+XoCjw27vJ7yeju4XuVYFsVtVpLrnTxHEtmn58JZRuN
TnSZ4VBJwXsdn0yQgGlYN4ct02ovz6S2YPrO+dHUfQTPCvUTj2ErqwUaKg4aqDBC
+uvjVPUkF9I2fQgg9SIcBvBLnBGx7PRumaABe60vsepaslM3hfTgFisZ/5+QbvO6
3JvIo14YsixautaKECEMUA==
`protect END_PROTECTED
