`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h4nuCmPXsCRhJKlhQn3bzNlQep6T0YVlah1ozkc3RqwLibaB/YTc7RJyI5G23uJY
P0ekUTC8j+9JvhOQzYOXxhj8rYmBfBpk/40Lz0IZQ1zTUIJPpjupeMabdyekmfbz
5MOSvWyxzZB06dxdxvFdNJV8RynqpzKWCmlqMwtHSI1xBlBvaMnnximQ0KJ+A3Ng
4EdsRsGHRykvikQROBJ3HeWJFyHwIUUWgrtf0hmk45dh3m0FVYD/rRRMOa4aICfJ
agjG+fXktYQkT/almhyEhlBYGUPYTyD7ZSxaQ7Z9+zsb+yHH+BmP3jdfYcR2jQzC
6v5gDqJZVGoP0e8j94TQpq/Bi151PRRTcfzrvzdIrBn2Sj1/TF+TiWVyaINJcnwf
xQ0CxWU8p2gkmeX6B0+lcMpUwBGL/vYoEPOz2YRvpnzm6TcvH9DuzF4NvzGKt4uD
sSZ/KQuumE0+BVwI11OvV4J8TyPwVAnUX3Me1vfp94IuzBIKQD9EptacEqnMGx9r
o/yWBtk3wVGPW1sMQR0ZQyQEwsbtvFgFKX5HhWTN7AIi12jNSdW1KHdDqUzfBLYY
5hgNsXLlPGTHMUbW9rO7E1/cQ3RxInx9iVSPWfBBJCEvTpvJxxrvNqHNZntI6gIV
`protect END_PROTECTED
