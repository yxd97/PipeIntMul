`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHhtkFCoIpwEkS2IrMnVRMglEqZVimILGxcJ+2tsP7iqNJ+AoGnuN9WvQz09Q13X
7/Idx640wu0LQFUUjoSjW3trArg7mxezTKvZluMR6TJWYdEXRGAHzI4UgryxhSAB
s6owD7t+XQAye9IhR0qDM8IN8XE17rSOv1scIy9vHUhl1BFgp264Upyo+/sA9e3E
3b+LOh1HvH4YMfxhUePzHPc8/qf6mHRSrpfcBY2c/YoxVr8tSLa66LRDVod556mU
OEjzEWwXM6x0YaqLLLd2pYSOmfBz8dH5bZ+D7nO1r4f2XD7XlMpidjhzQyS4xuRw
s2/ryfpSVRdTILlpEuM3F48sH0hUo6SiOtQwKpR0v91Jqje1q+F7o/sBp7yD6lOC
3xeSV1AkCbx/YgQS6x/BnkuSHU36jgDL3iC3wXZILah/5M9kuXVz8hzU5Ts8trvq
`protect END_PROTECTED
