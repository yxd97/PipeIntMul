`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yYmIlKdQzXLYRqSXHiXZJbdbyFnWghqI898tBfH2xXuc1WQkXdqk8QkfNuUgJyzQ
AL6+ZgOj8G5f78dpPZ6tcGEGB9ZwDJGXXk1KXt+3PF9nfMKA6z4qChh1Pk94QK7S
OH8GW7dkxkWMFUy/XVzb8NivbKzvMv+t6OlNMY82ojGwRaq+QrxmHGqBRFemQ+UD
ueZuSskjhcccbkPJ8ZnABKw8G6nuSC7x+iZz/L4xq8nbDrO5pT14jSO8msFn/L4X
OYMcx5AHSM3xXf8zQK4rXc4uiU/Xyow9KDHNTpijGIry0RpWK7IRkDFVQ1qGyFlw
CpXY6QVh3EAo5EDC9LsPDIUY6BsSWaGhUx2r0v6pbuFMXJNntYhlCUuerGJWO/4A
1ZG13ipfINo5myafCC22oIDeXDS3PH+RtL6dFKAs4t2f45MxORfzYrUYWgBNF2ny
aN7QIeCEU59gnK3tJnehb9mqw0KMWUlJ/SOwQ/oYz8ePJ+Gw7LCV+pIdG+1Q90/p
qEYApxX0PZ85UdTBrMvI5378NsWGKVc5uvaeyzUjBODJCb1IBfZsdr1KgNZIrqbg
yRB4u4SzKMAtzCJ/wBmqLRkDHt9K1kTBpEBxyR/jrbubyA4OOK1ny6duIYn+OuMU
pqER7EstdzVPB+nCuhNSyGeZq6RuX08jyjATBwzz3MF0dFkhm4Yh/tiqh5UJuKgB
3OgJS+RNMcWk9uLwdgbxcI/BPYmBEcdjtmp0E7sOjM4TK9gpAe4Zn7SFCVdJ0PYM
2kWoEBiSDDv//U+4rmGLNxrlGKqs5cBnp9/5oFKePz8/Nxvi8M5BPE95O5/dLcS0
oFKP76zqBhh8wdP9igJ3dFYQmGGw7xngJ0h9zz3Hz7eYKc9Dmaw8pSqhZzN9mh0P
nGnaDpjJkYaSkjg78U/AtuBdH+QVPlpUGllhQoXeCvg/+4pO0JaSWqQMurPo8mWK
YRYS3MS6BBAls8swvbrZa/fgNcgBYu8zUX8PVilWYrIaliQOqgh0O/DxbB6Qm/oZ
nDMClqKjoJNJHaYHU5rlIFOMPD18zfqqc3OZOIqlemwP+SJhFrxs2bSkuayWPkph
Jmpe7jsQzgiJhRZnU85y8xyLQH9gXe1MbAtwNQBwQM6UQAewQJYfXEHc3dtQRbGz
YAbMKNaBbLmbT3A1z36LsL7qRRjH4RYoGFLP1EZgmww0As1WcsbTE3LymZ4kRT2w
GO0SQRUPBUB0gTI3Uv2vhbq/iA5HrQ8+veOtEnMXuQ0nqcxUfv6pQrsh2NANX7vF
dsAkkHT+s4BUIujAi2qekgN17seAQLL9+MRSexipuqjhzJllwyLxETb5oQCV2Fxl
U2PjYURTxajfXle3T0HYhy4ClLViL6G2u8WNzG48olptHen+rSJS3ZQLPI4RlkCR
BndOFZNOVeCdemJXkD47rwKZ9vrAlxSMgNoCoA89MPgvFtuLUArGWOPNvsVYJnGv
wUeJsTgg7lm82y8LYUkYLm8vmqlc9Y64zZRUfUpuFHSw7LMUjZ4xsFYVcQPot4pK
XuvwaF8UpldAH+PWm+uzwmqMjpv4bDdCK1Jqsyh+quIReCYx76OBILmhmipampTu
s5HbaeF1uMwUAeu2cL6iDuuG66cMyF7PXSOUKq+oy8bcFfiBSyHsfwaKf+wipCuf
3TPbPsPUGcizi13AyACmj3nQikwPiReg0DFvQQiJyJLkLilqPrsceZ4i+ZgI9x70
k+oR/1YRe1G61FxR5Z5C74pnWPw183R7SSsUbU8YiQgVWCRIW11xFMgONp5PbOuF
XOeiom17W9TzEjN0a9Z7sbicVSiNd40TeTGOwwN9AIze7CjHD1A6xxPAbhvDQZxd
6FI1aJkRHnTndvC7/tGsWjaYuY/2xZ28nlLVc1Wr+ML0PEOKBR+GjgkhQJ99/f+t
Q4jWjG4XMh5O5DrQtSD4NhczAQT9z+eZH96w35/ZMakn7N8AXs5OcAaNGWQg4b1D
/yi42BdFQAe2S3V0S6473HzKfV4uFk/0KTb9l4kzoT/l4TWRbHqOomOWTDYzIqb0
cC5G/tj0fsDcbaW69tyJ+6QIbDjklTicaKbqYniib+F8Jz8HMG9iXlqawMM5JHPG
Svu66oIsc1UArjpj5Z+YBCB/C5d+BZrwyQvETnuiHFrf3vuKexRCxXN29GR7uZ7c
XoxWI5/Z2517v8OO/FAGPaSQKth1LkYlwWErmnXAilDqR7yFgJvdOfcOP0UDaDxG
6pCuOnr8JHRuZXWSn5v8VGvBv+Ia2VZ3Y1cAvF9s6qMMLy5RtWqJb61Zp7z8RfG+
sJkBQQXExGh1xcetY/xDSyXLUk7QFsW1g2OrgOyzkgvQ2DlYMIgkdGenQ7OXhWgm
kzGqQql6eU5CPgJf5drByj4Dz8h5b7TBqWTW8gByuJU4CawJAUOGnC8MqBq59zAU
FzxXy8PEsLvFm7NSXLgML0Y8O1eLEQ4U+Fpx3UsRI/z9n69glAcIkeZCcIQUx1qr
qFgUbVGgpyHfTrYTWl0rU28+N3bIUXKptUtxiht8DGKzSsLtUsdJFVC99MY0vwEI
vBuGNlAP8NyEHFywM43lq0Y4lgJldOBy1+3M2at1Qf1b1AoXjdpb2tOVfDm22xQN
f+E+bDPzO3S5Z00bfxbxv9t1qGLGdDGx7iOUprHtNS676619PKO1TWzhwmh4kKrd
`protect END_PROTECTED
