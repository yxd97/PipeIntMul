`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L7VxEsx2wL2mCxKdBWxDYvnUecXyNeS42mEsuj9qaUhKdBJ6KzzwGUTFzHPerJcH
Y/I7zGkKqVsPPZaVp+EbGAS3qq2qfo42HHnSIWJd8zbehEIRRfBhg5K6gUOYwdUn
zsap60/UV2S8ct0OtFUYeRGD40k/WTEMkTPg4Sbn26p9EI9Tdir0t4XBblX4/gPa
62iFImH1Z7SncmOs1cFSp32dtge2I50OdZe5zS9puF77GuAYGV/TKdv+rnHBEIOA
GpkSPAFoHORVbPITDeivSELEtWrp09dQfcOXFSSInqGVPYmUtaICf/lvcuR3QW1q
tJxhu+jzoSAfrgK+ROqDgDnxht9y2OgdcPB1RtJV2k4lZNZ1agsKS/qC9oyxC/7f
Ik/55i4VGES59G1aWYj3b/MJsIyFEDydJwEBf/x8aYMAn/0fyjHez2oHHVO+RTPX
VnlB2+LVsVl2wwRXXDUdbSaN1RBe4dLHFOdvh63pE9jiaLUjeVe4GT4Cs1zFiBl6
g0sIV8lCjIPLLDUMrzigCG2682PAuhZcLRSqdRFkrySMMImD21834/YjzigCvVs2
UzWtSGPikv41nEOFJ/kktGQFzg19M6ARBTH8TmaY78W5f5rMx+MOF2eL8nbVA18P
WDoOY3BGq53ht9NvYQgf15WYm+UB7S0jGCOcZmT+IY25g4NNE6jRrRcBXGjWZ7x5
WiXM1US5/ut8kG3JKFSv5GGehh6kWb8eV83sbyZkJD4dznZmwSz3f4IayXc3Srps
keKSDT3nngc1iEuCmSqpJagClFvfOffjsEanpOmSta8LmZ7rf7ad1CSai8kuaDk/
bDwXf09Fd33hQuE+v/bBrcNp+OOX9K97ZswTWWjeujXxuBdGIiKTfr87QdyPE2jw
rKclqSrEGEwwq8RdDpYhTlZOW6a40I3GuWTQHY6H0/V3/LZwsJCZSPJWMNDuW9Vd
+KSJlJJgBHTDGAd30F83x3py7SVDd9eRu8oaXYKHDSPQQskU9p/5bOlqW9XsE41m
zOkGQgILIhmy3y+TdGiYw6+gZJu4KkHn+yWmaV9VXhkmZUygFoIs4PyC3Z7zk5+I
ynOl/TiY/htCdGZuXn1E1lxu1SWb+p3IMTM9B+qi7uwnS2nxQdl0N41n1wAndy3n
MoD/fP023a+vhwAs+BujsmLjifj0CKU3d8rFmOr3Qc+vVwLAsauzurMkIrsNMMh+
5thXZ3AdUfAHqGeYxZ+dePgY5Asw+jRvMJP80ERKkYdPvsmLxqbS41h0dMLF1NwF
nYXb2WRZZKWgS90bPFBsOK/qMc03A616TagIV5TG7jao3VxaG0XGV58u4L5MCZlE
4vC20enJCEgemg6QrNCUXf0TWvFaTITL2HsyzZL+JSqwJYj8V2z95S6J/8/Xqyzw
t5tDA4brPGMAjnR2gTtUdEbJgvSnOUohcLH7elkVLCqpEJTfVglm7NgI5PGHKbsK
nAnrIDf5GUeRkoHR+c6m02AbmwXoqZM2gAEKqHCACAIR3pxkSs5TSI3WAR9iSJ9i
YiiLnVr4WQFBOpFpHlCNLVGp7wG2bg4P1AyM5RIiNxBvG0LoM6r7QcKhaQiiu4l2
6DsNxxpYfHpw/vAdP6xfGiRlab2pM3IWSyEhq7K2pruHQ6EutzQApvsod2bLrnKU
cEctK4lm6BWxGlNcDTZDQRaolWrOABlDlVZ6eQpX2nsJDatMBTNiPCEek2yIXYSk
S+BFRPz/W0tnDmcoMLhkkLHrfQ4lWd93DE4lgNhxfiOVQpSQs5M6hSYikSo9Aj1o
LpSA6r637dQMRG3CE6+nNnuUkXy1MjRtf6Ve9JIQCpkrfJdUCfPAU13BiAigL6ck
Wff2d9MlhlWjDh4ce4Z9CWv51GKgh2Kxa52U6Oknb8dz2hYUtl4qpLFHd/DKESR3
mUQZ7njRDPaClHvwsuIgi/6GX9XcLw77jBNahGYH4GcRvwjb6jR2LpoVSc8BuQdU
DPWsybY42mpYzyEyuaZ0eRPQ7cIxfY5nwwz2wVpCah491ppTE/0LPlMDT7ZYtFvN
BHt25NIcTlIzsjzCd82XBxn4lIUYYXI/jmmcub81Aaeg+zUHTUlniv241BsKnhLp
/wUFIbzJ94QMFRqr9bMt4A==
`protect END_PROTECTED
