`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fKc9h5IVEk55I4HjizdrWv6zPraPNQ1iC/C3OKCyNV3v6Uhd0zplDgSeNTHvov5J
bRZuipMK6A8iD41BsF/3H4+jdMlL1DwjfezKHrtezuXK0vg4bwydTkcHe20s6wPG
plXWsl88PKuxIszzb55t3XYD2Z8hvrDH8qLFbIhiB5wkkQg+nwO/jOAN9f27U6WU
HObHslY1QQ6Ly5BhfJwMF7S23oR5gz9QphsSoqfxeSS+n1BpnBj4JYDhkUkky78c
qOQeu/nYOQ154p9nXiANrYgxbtITcNOCbG8U8wRzy20et2eaVwQPczK3hCo3bs8S
7gRb7bxm6WyD4ch9+pf0XCys/Pz8lrAW4LrLEpSMbMSr6saH9tnEk6dlshnoLtbZ
htYig+kpQ08PHx4xzeHzdSuL/vKszkHbipgOlFytyP6GmGUVivtNOc5piCNBvoxu
mwiyd7fN0F7Jpdz7Sk+2+kVz0bjinO/dHrgQQipu82qTyjia2Vf2dF7QmMF/XOnu
Dis9/Vmzib45WNLILgl3Aw==
`protect END_PROTECTED
