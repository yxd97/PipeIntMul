`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCgY7J/17p1P9x79ysqrRMDLfpOCKa6CkuF/huloYYaTcbcG3XInLkY1mRQNUOCe
g6LI407bFecAGskFdL/QdsJ9i6sQSyJ0l9k8SwB3zwkyhyBhnVGMB7jj1L3kn0Zv
+FuTIdhJirGC4AvSi51hMQIY8kGxpsuFop8PTTTmKvHAdb9W58IeXKEuY8vrMXiW
jp3LF+ryg5cFDVWrPc2FcnWe/XB4zOOZrGK+VVdkrGwFHHA7rEt2g8i9ccueh5fD
9/5KND4Zuw+3QFLxbYZA9vmBzbEBtyjmnKzkHNiuJW66nQcO3lC/3ZBRiDvqqGx8
7HPl0CoXZEsQapkLezGHLA==
`protect END_PROTECTED
