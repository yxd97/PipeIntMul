`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqiAFQuMitxBytEklLB/BQ0GsLhX4Thm2jagJT+aLiMHLhpSm9Ug3GojVOgwc5Oe
B7y4HjgPV5MltWj3jlXuaXli8BcPlWc9DX2ow5+6SSwoHFjmRvNi3jbc3qoXlbwT
yTT6Ar7zZgaOvqRKyjobDbNG8BKaTB2FRKmW3lYnAJQUv4EBns72eHYyVAaWwA2y
tNndC2kZDUweDeNeR5CMoNtfNQmVJdHP3vAGgt1CYYTB0ZCb8IIs+832wiy9HUZY
FmYae5lnMF/dby3GKRH3TXQKEP2LeaLyssd4qrKgoRix5GFfhmTcHZu1hwJ+NpE+
RjPvesOFRu6gYYeau+OzP9AizXrX7PziY8IPOtSKYxI=
`protect END_PROTECTED
