`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEHj3yZ7yvJAENJ8z9VknIE+BUpeuVXN5JVTjnCafHnjdNsEIATXBNfe8kSzRL7H
Q8oGI0GtUYObmJgVTsmMEkr3bx/qNtmhRx3uxAaATFj+MZgpsMvloiqQQ5TJUdl7
v51/vXZ4VIH9z79WZ1VbJK91Ab2vtcZC4+kYGPH6JeCE8HDzv4xaiBWvHwm+Gje+
C07y7Smcl7Sy4pWQReJLArfiZJMZJcraJchfJGmR9HdUQ9BanyPsLJUmbu/r/0l8
VfUnrAjkARy5Fw0qNKIE4Jk8WxY72maot/6ARo87y+T8dVCY46ctbZiXT0QWZaRh
NAkNUXbunEagWsR/eY9Go0XtAX03LrT8uwWl9hY4M3PCp97RtlqxIOvq8B/6Ew8f
M4W3UOoCoIoxsTiwSbMnKmwDXZ4EACTgW3G1JjusDqjhwDWU/UMRtLVyrjV5jRqT
LxxpcLPMXya/3UfRR06uvxAzo64vC2w7F7Ax5IfeWmXr6k4FMMzp376xpImNnGah
5qycxL1VK3zrpiYZ2WNCeIy25WQs7OqBCqJN12Pr+h7UOm317kj8PDJ1iLXemiE2
PmWe+l9wgnAetVPgrp1Zw7P/4CU1idVSjtakP+kEq0lGfgHNEdcwPXj3KbQGeW5Y
rBD9C5aoFsyYU/EVgFADaROHr2jwvJXNJk3LMFWLLjb9uBlQaoWEEy8p0QYCI+Zp
H3bRMV7/M7BMmgCY8lPuTl1RV0WCgpWuxBNnt91SIaWS6MEj8IgApygKPhf4qrmO
E4X2zhfSKifYJ+dHO9S3wWXsXmnAh2kRdafFEL1oqy6mJghysGk4yi1u9cF/oKaa
WhEH9FzGzXTPtVmPDds6iMIznzWAsiFoWpcHrcSdm2WLn0csAHFF+cfSgcNHQu1i
7U0S4yMKT6xSI63rDtpnVt2XDFlbUnTkf8uUuA1JI1EfwVHiqueQQlMR3gAkE1dP
Z5SLKENvsIaJwf65dKI+siODsf5JE2dkMuOKF3XksMIOCncbiLHnr3pWmEeLjMQ6
msHLYrZAp/iPheACamBtMghhvvh8kLROUr6IgP7+8RNx94f7VMC3TLhJ2F9zKenc
oKhUlEO3zurnljkZH4u+a+hXrMkULf/NZHwO0ayJ/eS4irogHFPlxYvqft/IaP3F
F9UcYtM9D6sv9ssMow6neD6mqP59cCMBKmDQ/CthRD5WpxSkwtTsDW0hhUrbIknV
Qk95PXwEU8Dw7DYy01ilbqln3TkSxpRJZXPde7q/XI+4fpFoiB7mbPBO80Ad1y+f
YCpGsXqQ24Dz1ZTOozyj/TjIFFoDs0/bwOmgbz88MZYXPtW53zk9NGBJZXvcmyKk
qsS5UIW6o41VRRmvCXGUEXt7I6no/4ZZ0dL/nv2FkJ1Cx9OQ2hlvfSws2WEeIlt7
NjjXnuOTCjsC8wgfneisLGqRGnwZ1rk90ZRi+YYvFla62BJ9/Fs94tur++BpK1dy
RbkpFBirLi9jrCb4FFoWo9MMuB9gLIOvlJ132HZmJbCHz8fir0wGvoqWRlhFSDo7
KQUh4DjLa367laNEQ11u3wxp9UY+CwLu0sTqam5LVTL7qINVKWPn2Z/Ylm5Xla8t
+nJKUdopYakSqM0OFikfoW5EavSdgfY4APFTXtAxuOXOoPf7q77Zsl+QZKqw32mq
F4v1+UHdTWGD71xV19NqlR7DvsV/Y7mz9Hg4YgFJ8o7xP0vpMAN7C0iJa++Almje
/STttEx0g0yn3H3T1gpWtvNSkf6I8k/R/5iurF1QFC7JPsUiFQSUoyzQ31IOOI0z
+YM0qT4YY0WhedtamXJjF7IsLboQSZdgLOxQDRdfwdpcF6oFALuyxb8XSgZrCOz6
BaYHxLwrscC2EmJpVBY/ndc785SfZ0hdZlxdaa5BIP1jw7hiEKvnTEl/Wez/P7nZ
4Fig0jqPEPjIZwLqX/bgpnofdtVauarMuqtCcvjVYwoB+RWigu0gBvPqMzwWpZbq
YL6A26wc3AlOkgKl0szvEgg43cop13wUseneKMPq+MybZmFYT8b4VHTh9SxXUODN
XPZIhPAqS/scP3KIBoXlFkzDxw0LsXXPBIhwvuknKtlvjkHdGYG+pXN4ZxwgKdC9
kwcqUxbKrSwP/1+g8uciKsRvGT/QTWBau1wXA7xSIUj7Qfa48WGHX2UqYy1Qb+/B
uPPlVswjkTLOmfzqsQaU30opfRasFQaNk5vm7gE1QYIVrrPqe+kbTSxdObLXTqqz
OeZAzTifuCig7IPVTqlfWXwWyM2B8HlFMS1ncUcMVGiezSpsi+rbd7yb/9Nj8r7n
fR+o3exATLvpaORuggsV0jWugfghMvhio8pDe90z13xqWwavd/jBD/ZOXmroGSjd
`protect END_PROTECTED
