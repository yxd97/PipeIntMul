`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B4AUIUmx0BeM1t0D14aaei6ZJPDku1HMmTkZrcNH/a+KT6Y7SK/MB0PeaiJzPhlK
GWAc+OUx37bDNdg8sk3tZG7ZPTqt9tMNZ5V/kvcwFgXKRk0W6rGK5PAXqQNPhRY3
CHCRNdFingCuFcVXAveOYO0Mc7PPnbt0cbREqgFhG2Kd7Y8fsKd24F8y2gJWiQ15
WT8hf91sb8HoHSLlAUmo1iwBIqpjYSOnUuXIE4fTx8F4sdOkhqE1b3ZTqGP1SsLr
9UAKYsmur2jcW1BapZZmF0kJAYoyKmOBGQo97CzdYEsd2Wgp6qfFEqRjZobVASkF
jqEOau9ydu6Rbfy5k2kQBzbUIyXUWKW3pJBxHVW2JXQAksYpdTxa9JrB7kTaaObf
3lc+mRFF2LYt0+Ft97hvaiFVUGpmUVo/MTogb5l3Ds/+VoakQzgzqWI803SKt3+r
tPzYIhx8LmqHPC52JsVCtoeukk3U/thm76wWUrmRIE/pKXEBxApfGoZ2kEJQRifE
KaI8Qnl8NUqMKz0ZmwkjmYA0BTfSIeKYOwKiMu56ytLu1f4HoHafy9YVjBB+9n81
fAdJlN8RntiIyf8G8yWZWwxEW8QFHVzHzR4h563DG/hhhwCWJwfEOSPtPDTK6dQN
zwrHkGIWAux/DxhuUYrKjC64XVn1yYe9jpLtxWnOAWDuJCeKHRaTZi1ewju6Y+he
xyHQEZmOLfBdKFVK7JFdZEyUBxl7zY078aWANDkkyzeCoE7vSYOGQAQyackmqCCB
qvTxEeabLiizuSGgTsh7U04Z4aVx5iWigG7c6heN2QLLPBMUiVgbaO72L3gSSbKC
FoQblvu3UbrAXiYaYC2N02fzq/khZRsTxhUrc8CDYs5VpGgdoNSy2DUvvDpSHvIg
ceBX6MI13/Yqzm1fvdmcxwNs/Oj0amRhcJNwBmnKCMqDDEmkFHzz9aAo5GKEBQXk
`protect END_PROTECTED
