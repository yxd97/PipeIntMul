`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QS/mwjiJvU1JGQgrXfAN1O5QhnB+61R1eYUk2zGsIX6D7ThR8BKnvDH/iTsy2r5u
9gOMWiDIUzavH9/7sqZUXy4c/V7mXaF8V0YqNXVgj0Kq/cfVGW9xFib7C6GgZ9MC
QjesD2w69N/rT8R+xClCOdR1KYmzHJo0m8f32Wyj0dBlm+GPGnHsDoIY9zPjPTSp
rSzzHB07pntpuLX8pvuxSN3Q5yTiIPtTXyLi+kf5e2Lr3nCGlYSI4g4XcaVGrOaj
Tn0JZxOcHCZEnMrUER8JTSiSrEkBWDcVnqy68m3qzAFLLdCLj3UXMhmYOrzdjOtP
gtvn87EG7soCQ9OU1MIoDwIUxW4phRjXKmxrrbBKER3FoaxiSRZfDFUoKMn7FF5d
AdogyXHige3TX8i5yLLHsS09QmHOLhX0vgwW1nuRAYrGYeI8/tjhmOLHlHtcnDBr
aoNO700t1BPyDkKvLb3zGaHumi1MksOACGQhNwBBLTzRUKm6M6x8LSmq2LcsMtZ2
o1J3RhDewum5TpkRMuxlAAsPPbTfUGinLI+hE/V/vJjZjv8BvgM8uMTwl1mTuf+/
f/tSYZpsJ3KtSLwgI2NlOGg7YyExiPBanZO4jflOtk3WRg0Hahf7vByJQDoy89lL
PEsTJpIogjd98t7zEtBwnG0Nk3biFwuaqq5BOb1Vwk+bF//xoWFejBKtdWdhYw7Y
l1d4rMeXmTVVZxdXx/5Nf22vAhYhlRIaY0jZSeqGOgWUcjdGqezDUojE3NJl9g/B
ReIJ68JRgQt9zoOesm6Ib6X+iUDJ3N/1qpt/5HTcFp9fADc8slHCcw6zbQFIy/Fd
TKxPm7CFg7CfiNC+RHNI+n+mYhma7QnGsalmenGC0hw=
`protect END_PROTECTED
