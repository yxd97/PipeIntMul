`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CqovoBDJeF66BejNpelGF5rtgtCk0LHAcovhIOoKnOOtQCzKhOIfx/zcOlRZ3EcN
FRleAeWW5KDTnGB035Il4FkIFjeNodtQSZaxPb1WiKHZWRGBbBjRzwlHI3BeNfHm
JYMJGITm9+oCWXo8VDcrNeezub3iLrUvE5OiUrxEHDbH6AyST8ixqaBGy1P9o9ZX
rMR6Qid0DMyEeD7+7Mwub65jhtnJPB0z7Ce6fcbD1zQE5t19FPVdRIrn4Ip7JlAg
+zMpQ7WJpKY2G3NyPZhLMEmq5C6eRD5CGaN0Jfkzj67l0fC3MmeBT6rqJUjij+Jq
c4etFujJxqeXuXgZ5oFyhg==
`protect END_PROTECTED
