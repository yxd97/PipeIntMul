`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sh0zUirn1BaOMmM2PHOTYc7cqAI6Rb6Rz1/RoORNR7yLULOv9WvL/22gARICkWnT
cykwQsTKGVoX5FnBGjUMNeVTJIgVYik0nlOJCu4A9z+feexKwISxNVL23YlDgt4L
skp8ghVYBTITrCuHn6NpO7QI3s1qYNIri+6CwbeHA/4bChROHVsFJ7Wwr3POIe70
XEdpTLZxJogoQkltd9YhubtLJmh+p+lW1FcPi9twsQAayqOVVr1gr31AyPEEYEw4
fMNmMOJdoHF9afoWaTYwuDcgDGqrWawklE9P4Y+VgcYKXbihhrQx33Jx+JIOlN3T
hnj7gySbzniSrdNOu7MZe5yA+Uu13Mj2M6p/uDACFwBHt6QqsDEuOAiZJo0h/7q6
4R5VJPtm3YBKuHej7IORy9uznoHwiRNnPqucMGqQgNcH33HTIvvAyOhufy8VOin+
w1cuAjzNbnkqWU5ukVykyUkVVb1okcXXSo8CWVai7a8OF/odYqGsFI4Lqm11dScc
6No1A57Fke1BzpFD6zgwpu31hUz8iH0Sp3VjOmBtDdjDswvyJEBX2rKoGloFMvie
O6h9AKBuBCWSnSMLegG32JGmLMQCg8ov4wZ7x1Cfu+lVv2tZTcYwgb9cjgdjl4QX
UyB5E6xuRdcionEobxbvYadNtbQLXGpRludhoZvL7YQGQxm87xao369PcY2ywo8s
/dVpvciyqUhFjs/iWJmSjDkCagSJzwI6l4fISELbM7hQgEnVuO8BiViWtxYdXiRx
7btV12K1J9O9DlxPDCvGAch8lxyYXp1nA4SaUs75WMGp5wSvaUJn3WpyqIRZ+nnj
ouO3oRzbIsPDz5VpUJcfTWxNhVY8AjxlCyfEhdrKKyOmB1jO4qxpTCiNZJB+Zf7z
bPOkJ4mCu2phJsar9KZsa2SYb0Q87UXqtWPn4GN7HQr351LfWGk2jriXMWuFOKg4
3AG11Ro0ZhkkeyPtTCEUKuYBMMEfuSOO79lfRG78BKjzUPznA7vtDHS9bQeOD/AK
OeKSFJ8y0lnO+fbw5Oar3TDIENzegxnr2Hqb45IVppwlkblrYipcgyProf8eq1gg
C6HxNlyVIeQVifOPHVGsm+aM4RBoUJ6zqyex5cOI1tkmzswVmTa0hnHdXXrI8XDt
EA/Y9puCydpSGbqqTY1BAP+KU2PPHgEJ4VMAxE5PgkSb+Ob02Expo/u45nC0bBL9
NhdfRZeN9UwFOG+SmoQSkylEgfhRbxU8PmOa2r5/zxHwEx+npSgwy4VEK/g+VYe+
ZZcb2Tk0ZKfapVPkhDy+Vs6hOS/PBGZLRPyII6dLFQOXuuJ6h8OwtJHeqJLuvcQW
TMKblU/5pyprK6d38baMn+kHUWnQpQM45degr1umhXAEl95wKeWlyeFcliUiDBxk
BCXotn606FAOSb9Bh4/5+PB8TRw5hcQjCvDxqkIhhLv+pa2XuT6eEkXVPKaR0+Wq
ZAFicl+Sbvidr3TXpua/VwRJFMCH0FHQE9PPzD1SFOjJ9UPnQSQn5Zda/rtfZw6R
XwZZxVqeQjhMRb+LPldInoIFE17KbhaeuuIYQXfnW6XD1N5ghPPjR+MIDsTmApbe
5Cir7VohILvc8o4QonagYpCFhjY16l3UL9j4yg1cE8o9TA0Ir9bK0wi09kc1l2L2
nOOge4cU83NPi5BmY9pviKbgku3gKYSPzdIroX4+0u97l+K6K4tQnCcaOYvkKSW0
kVdmakyVoNU+KkHfDREHI9e3ooYaQ+s+GoyBdOSZ32QPDLqt6DV+hoS60Imj1B4q
d2dTHa7QxPKnAaqJVrW7HhcPzXip8VU/hbxaveP/PXE6FNDtYCT32ClQ2zPQMZpD
p8e7Obzokbs39hLhMyyEiUNDTDa0ACgfeVCGSLdxmORqMfo+yKdwN+K+PWUEitil
ZtQ40bkt5voPSLazZ0EDX5LQIrVWh6QL88DTG2RYEEdrMZT9TGv0lC3vtB/Rrboq
cmLijrjTEdSjAB4qcoRy+VLPWLS0ocIEeOfv7bdkkuDl3Y4TANbSxHXlP4cyMXUC
01c0gdsl0EMSHAPtw61Wj9PXm7XCRlyT4KjqmYms+AJVBn+HE3k4a38JpnoojIgQ
4yjYEvxNxicv1JEhi+JR7ZGQF+ffu9X/Lyr1K+vGiUpmcSiC4ZFVC2TT1nBO9YzT
YQkozgQPUzjjKM6TcMa8vGPJ5gFa9zxA9xIVx+8ux53nX1n6WSDCgwdVYCgVnkBK
qliD94qqHeL1O1BZtxskfLwYZhiPvTIDnI92o3bj62gFhRHtmIbTIGe0ugvcWiUV
`protect END_PROTECTED
