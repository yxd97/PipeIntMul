`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EFi7Wuf5S4HfwO34pT8fsiOI8I7YZ9VKWQ4y9V6Vjt4NRC18c9fFHDbaKVxJPHdW
0UENA5LhnIVdpm+1CSPnrid1fBuibExXEwkrzmMvhZQ9zQCieJxnKd7XLCQdhJTu
/pNwIuQtN8cJBit/ASAVM9SDXgG4azz0yac+LROMOnF7jWgsGpQZCJZt+wjAjxuY
IhivKKBUeAo3ETPAamlcS65OaTdDYVoLqBXDs8vNdFApom9R+ZVppePoh7OIw4bq
M4ienpiltEu+RfdtxsuRSAcLNtNTK9bQlRuORbGNOPDdGfpmA4rE/giRK8H19Xq3
fUk2wKFdiA4oS30OWYsvpSGwinSERCnvrpMv6Cxz+o4GRsDjN5xK+0l8Wd5WMnHv
BMk3+i1moASHzalTG1Sm3AnC2anIToAuVA4i8F7aBtq3dl4f1qws7ovhl8ViBmDQ
Q+m7ExABdY90g48rDjlZv64BPK1XSmkkL7ThhDF3Cw/TDnpCBRqjONls0PYs4HEm
XarzAl51NNVzVLzkGEKfFjswlQeGeCOe9ZlH4zgYw+geANKduVWwz2WrLJ2zInQF
ACoDCtnI6mbBs5878DuuDZtbgZlML53+gVF7amYtXU3eNpt3IbWumv0sobKjBYyH
iYhoeVPGgf51OyQHAukszcfbEwtkQa9lm5OS9n87fdvk3+RnI1CgK+i+NnYQ1ypB
zlAUTegL93MfS9U4m1BVVEtmYgNITaGyXiNxwpmW/dgFeDKa44+hL+N/1XSYTi+c
2RDDfLCP2ZVS8NXCMhlnmbu8mk9vgfCf//y7Qha6XwCebSlEcwkSpvIg2IBv3fMu
vd47KaLErC98lkO//xdGnnNUYbTBtJvcEOScwBPpsb8B8f43LJSnrMIYUJPux1yc
rdWpmaQIV6aOkURSjXyAzD3rFOcJJAjf3NgdBxJfOelp47QvQEf1iCKxLgjALaQf
gt28ymmTTeba6pvRuLmbKp6EYjNCBNYu8uzgQud/evIDQIYZdgqWKknzTgIPyruY
uQJXf/LrPYi2wZJ2gRHP9I0FHufRY4fEoHJOHa3Ia/QWcC1Br+d6RgmPM3AIt+FO
DEH8h9Hglp6C3oLtUpCD0CWXaXVwv7+xfMK96X6FWOIyF4tmRM82+U4iuRP+7Qb4
CzMhv73jIXaFDCnDuJt1wtxmfNJOH6RFlAk257gHR1GXyazz/7ukwUJ4SiDJPAxg
wmEyyusUu+llfGB26lpaUBsp4+83wobD6BLd8Z0GR0NPDPBbdney6+djmmVkkblI
7ETHks2v8Q8zqjK9KvctGKM3BKWTKZTJ+UlKf85wz1NtODG5Qx+BTh1yUQWEbRlI
ZdhcUOXj7ndddlhgxCbPwdBcsvSNd2pYMeh86GsKD2XM/+51d1Q9keitVuDGyWUa
welxiO8OAZcGQkIGlNS5cXd1cuzHp3fVkRJ2xpk2XOj8kXLj5rFHtzFaZdTXHvUi
58YCIxWlBmyrJtBDx0aJiAoRkhBoJpO1NLcMEsBYDAPl4tyDyBvy+NS05lJuvbFB
2wzQ4VAMsOgM/B6b8WihtLn5JdVTLyzMQQw+Hp+mrUMHun8duPA01DHM/L0sFdGU
MkoKYMsUSeHlH/J0nc20tWKktT2Utb4WdnTEEP+HTWeuQ+ztGKZpxx79vCyODyPj
`protect END_PROTECTED
