`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UeUgwRM8mr14Gm7Vo3N9bqqp4+HaHgw08dkQPAFVopfZFKv+k54ECSULaqcpSCk6
gTGepvpZ9cgEVnUQx1Hrtp9KCvaaT4Op8lipQcaY1djmfgyElDrYnik4w4LP2bwv
mOrP/v6MGV51SSDzIiATsgT1Ef0Tt7XhAQvQrtLkztMm2nNzCPEhaUd1vccB5hNY
WIpXB5QnHBMJGidXRQtetg967WI2S+PxgafDGqJedfDKJbqIZFiBY/xuiWfZJXDx
`protect END_PROTECTED
