`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tPaB/agdx9CmK2nnqkee+BwzCN0qSO+sSaJQMYpb3l/r6PXJo1DR7HMuNxzboDE6
RhKVl5vnAkTJ1bPvoN7u6APBOHVe7Xg2hcoUx3fCwpC87vpizId9D4vgvG/gl8xo
th3zQtpvwH3w2uoSVXw92ORQhepMExMRSKQEsK5GMhyfyHMRcZyyElGN6vUOnfiZ
PoA3oG6qNZF5+t0u+IDoDjteBfXiwQS+M+0kJEwfYCRaafOqMqn9nr7tcQX3pLQr
3huZxzRdGZHbmwKdXN01baAJA2yQ0oMt2CjpvQCwG0g+5DnN+boADxOf7ofKPT5h
wnOFdxXEHr+8AO9Z36AzzA==
`protect END_PROTECTED
