`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yoxvO4GMxoJTxsXBqogyyppT4ea0cxksq4IfLJmQBUxl8DodqxL1C+bfNKZp/CpS
e07+MxLfENFm86q83ptdPAO8ju7C8Mk19w7xK9qh+bpZ6cRsbOBKhtEJKWfqihah
atpXdUni43WofTc+rN47zTUgRu7yj6GyT5gp0nSy8tohenlsZjsR0JcuPOlAk6Bn
HOXyygStOhU3qYAPxEa41Qwk3ZBZ6yAeF5EfoDHbB3yqKEnbQ+Y8cjs/pgujbr+J
t5uyO5idv3DxUkE/DRFIwcXISLXJUEXXji8Xjaz1Z1av9AiB4AdAyAdn93tkWYDb
Q50gUDnARY5yTpKo+2aBxspDaUteGA7yRnyzMDAw5ztKyDdadwtsWw6qfsigh1cX
D6CI6SLFUED+4VrGKKI7oA==
`protect END_PROTECTED
