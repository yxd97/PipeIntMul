`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7hKm39X3nMX4PcH5NYGKLec1aK59HuR9dk+y6ARyk/pVxsOpx4YCFA4zeR9PO2q
K2f0vyfshUknOdxUNu69g6L0obhGtekp1FqwQJQtmxX5mx65jkTN7JdOWBxqEjqt
ENeEKsSQdZ22Z9YlDc9l7Uf92IscbzsqqRQfhBatK/iL0fKa32rQDmkLqwZ0AP5x
idQYmv68ZLlY8YzPWdmp/Qx09SBsd82TiOKvtK63uiCFtA8Glp/o40QhUUNqUQM6
HqxTg8HsU4e0GD68m6+53SDfSb85M1F5WsUcxCPLQM/5eWHH/tGP054dS7qlHWNe
ITG8pD5M7anDbls5UK8W5rcSh/exDmD0uHsmqoSmbbXuP+kVddXVcRbZyiAGBI3D
GBiDd1TUqxGBXwTXSBi5CKMZzLCfSdXToUUT9fPS9IHO9FhsfNnFj4sb8o5mbkty
7PElu9QvUzpDVX/3+n9OCyVS/Xk/0m5blDzDwzawxx9rTsjg7mTDFlBQx4PK7U4k
aycKZU/F3fJCME+d5/VE2Syr23GiHq0VZeHT9npUjFRtOKbs7iMNyO7JQApvp91F
qZ4K3fCdGMLsGg5gFlydUBEcKg0tMpbRE3h8KGHK9kqfJh+or0TW4xML6IE12WBI
tRn94vAz83bpEeQQ/9AA7g==
`protect END_PROTECTED
