`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FtOHcKTrEDwsBV6oRSyTMhHr8/zTun1WK6etLe7xxTriXdvP1IQipX5bIbbHPhnS
zvSeBlbFk/21JcmRG1LOudSVGBvHIv9JreomKfpQI+eNuHn2/2XzkqCULh8yNL1L
3vuFMMryRe7aCkycPj7miVNGQoORtB4u7SxvhMcx/BpyeL70nV3m7OzZAQjYWfh+
ev+uXV2/nyrbCwItBZJ956ikeYJhX46+HXw3QBeMDXyYmYLYvjLtqHGdGPUVtB4l
gMsrlvhqXpsyhE5JbfX6AFGzE9nCZEvFxQ5LmibF2/4IHbZpxE7spKrqbm2rM9Bq
/1618h8K8QAfODDKxJc7AFUKI/SHKqdqjtfPC3nEZzTFxX8thvl6ZsvA4r8VNDd2
VoEeItjN5SVqj2HcIXkeCGEshGetOP52ohne0qtbqvZrfQvcur0m7Roe6qmCJSn5
Cvq4c0G46gsL7nh0RyUE9jS56L9YnEAarPwTz+BcT5ln/AklogjShdflJACpCRwG
K9h3sCMGk7SaPJK32//InVSzpTXV5BSJBt0wvG0HaovLgs97sKrND2osxaXfzhmq
E4V9dBemxz82goPp8FvVS2XXjS/WUAo6gkwgErPSniYYXPBLgMWdg/2eP5M+43G/
UsMw54T0am1wemGcNdh9FED8IV+9gHZjoUZAQPosNyfCldRgTRXSxxknwnc7V9cu
l6jxCm1Nz6l9CxXCJfIU3ahUqH7gc9mMv9FFfE3if38uDqSh4M8nr03/wh6IIxZl
P/xCXKDRrPDkok1Ajh6vGxTdkKrBz8CXRxm1TM4EsW+tE1/4EQERNyuPI3hsn2Q8
tPT5DW0Le5lukJ3CwQmlLDld5Nk5V/fbX/gFq6eR/Yzz9OM11Kj1T2jKKScIJrn2
cy6NK0oWleJ65C7WqTv274W6FSdgCKBLTc0nHUanso68ZxV/IMQqY9992NtICZV+
wxotm18atu1eJ/8rXugsH8ktCvMKtQlUeyTaDML0SZV6G8SEolVWVqPlsTWbNPqG
ywEqOm5uBTfq9UHu0tfDwyrtP4kcWjAAvryhQ09hGS+PeRDf41o70w5LM/9IIhk1
SRtAd2RIgtV9XuMU+yD+ZyxoZt2pBaNSKNYt8vAfoZw6CeGI7/B2xwW+qmd9tT+Y
7mmtx+MlncoCrRSq08DwwtyfuZfnxg3Whz9AMkqKRITxA2DqjF4umj0coNVp0Jfe
LVUf1JEmUdklD1G6JJT2/25hxeCV24Wt+1tZNmMvnx1KKI3OPsp3AeaCGxyqXY85
o5nSelbULYGabfTY1Rpuxobu9TDWexOoR9h4sF8YQRaCiwtIDd0fRvmPqoyM2+W9
bUrQYdrKZHzakkVf9Vv3TLiyjttM+medfWK5RCzZInHinJui1WEXbKQbCYiYAfEs
AXa7eY4PqhniH7UqJ3enyK25hGeGSNV11j5fq/uLcUfYzYzjTv5bMeOZQ/o6rC3N
EfRBQtK4PwyuPerYzteQDtn8G2+fGDbNRazrXHN8S+YJFFXNBVA+PuHpkweEVjIq
oDJMyzY8mHtDnDnMym+0/HV2MTZJtVQ5hvGcYOl7zhiC1kChd+fHPFtoi4FSb83S
ntfTEGl49SMgGG6ld1QL1pVl1i7yQAbqkKSCy0p+OcmKWjJbyATVsOLhR8wF5x8a
Qk9DrtuyJBA2fV9/K+Uy7m9NjMLZ8X7RAYol5Gs5q0lmCnzDeaGaE2oenTLFuNep
seVp+QQ8qMCQOosCZPNz23f7J6xLiQav3koPi1CNmo5Y6smu5MS1JfMGKZZ/AGiO
xrUANMP0u/uKXlk2H9MneY2V0Np7cnxvbkRumCsHUCO8YpCQDwBYIbig2Me83Gpo
etiYNmk2uKvq/IbmfQzcgLnLXB4AlchsiglfBGGQ1CAGv7ls2NUXgmUkkfPB9V/3
d+XFXd9mLiCwuvjxlKsSH3gZRL6yeKZ04B2tMrWlH+lFn+4Ft2nW+RKe1yitl9qL
7vpUUbsI3u7SC+6QBtOkIjb6/ARMLH3G0DAA+IW0HTRXlaeFNuRm2PXYf0Fl1Ubv
+FRW9SEX5lfnDqFXKfwSUMB5jNzX16rvlV6ONuKm092J3binblCiIwoydlET5UWz
lC2Vdb6XBkb4CuSOvCe/t1q4fHZdBnj89OYebbaap1tPJO5wu5T6FWmbOURH+tZV
Iux6nSpaBt66gQCyZLvBdk3H3uhIFBq0e62VNuybaOuBWJnFRjdykegZdkGvqqpi
WhwaMTbQBoNRMZ5cXQ6lG+q9xRQnY1W05/MEc6QKScjeo15mpz1mkqKR2aFKco1J
eLfQVSmNCLesPMkmdc/v5Gj9w9S51Z3BCGZ2DY9DTDZccv5QOuxNCkmp9uqtoePJ
LfNd/PtofL/eHIWZoQzWIUHa4nYirQFyJPCicMFFiN+zZJO1E+dS5fvBr91MCE/t
cT0wgar2q+7QUwBsOu36S2QO4LmE/7xLALQOmLWCHSudrVlcJIFudLUAQgQ9qCyF
2G5Pav3WRD2AJymNt7k02j1QXXMMKibexILhEYuBkiokn3bvww5fmRb7lRyPR62N
xrDOEUySYHKGqUoIrZmouTs86WJOcu2c5KA8iCnKhOs4lMyx9MERTQ2j9kVmy1cT
TCSFnNupDCwL3X+gHnVrTTZ350+rRKtyKD6bjI7geW1K6wCEzV+HroZ/MSAloRy0
QiRC6ExGcmOdx4sjSKfu04lhHHkuXiADYNOVitohIBM5d5Vd6mKnuItBAR7OveKT
tD/HuEAXclJ1ez1bWS0igZYqDQcZZvtleucttxmrea/0uvhX7N4gt4SJH6k5lH86
6TK4bIHVPuc+JmkAkMNtO41B/2f3nf4i0D7UtC8w4kZjj9HJKcvYAdD1WFM9yYtR
pndWekTUFNqfSQkO5rO9B0xu3uqL7IITL77js3WyeYc1EiiRkGiLq+cBaGv/u1TJ
LlkNkYptlCqSlARaO8rnolYvC2MO5YBr+nfDE+vXqqmEVzjLaMa1RCW1irqjw0Wg
g/2Wd2dejM8z4h3259PfA3F2G+SkK1Jhy7PnPAmcoFiurSniv/rBAqVjwzTcPyCA
svquOh5+VAvCy2CkabpoZh+7aybdLIRwO5fxQeADT+KyFkipgdKkXL0YniXWIlhO
w9SNlEWGQle7zq4roK4DKSBwSuS3UyJ9G6EIKLpR3CCfHw/Mv7HwJzE+6/WkfgWS
8P5/mi1J8UTGQYoqMl6smns4vMr4Og2CvA5SWsf5hnU0p2c5xc7yyKi/TMycQofL
yJIhfWzNuNY0lqvWu5J+y59Ju7/QTXlUDt6j3eTAe5iBavtmGevPcjAaVvlQdTRJ
3Evo7Hbc35FQ5iSf4Sc8Gl2hkg8rEFpOEc+gvSPqMysOODXJ1chs+yuNJ36PdVO5
8oSFBG4PWYnsMJ5olOlakOzLQou8/A+qYlCCWKpRdeCK5vnZwHTVlryBl/opLv8/
5OUcrsNMA0yVnMcnTuiy2RrY5EeO8oVdgbNLFA7gudHuQjORxLCC3ygpfWZyOYPh
/Bn653yqZyi2bSmRVNs28pLrh0Pt/VZF+6SFeVm8IvrCZmqfJTN09TKnaB1I7v+W
OcrWGyvR0q5iK4IJOEF7HIhaFlinNowjA4jTEDa/6Q8XKY0ROasyGp/S2H8oto9g
/KXxGj0BDrOMDrPMA867Q00vRfhVKm7ozHNqd6hHKFfdRP58QkGEtmKzkLciJlgC
Ngcw206u7fouFd1Wih92+7YbqQOE5d7Z7R/S7WbDTPllXp5Eg4y4Z/G1B8TTMrp9
QLUuHd0o2BTsXdt831qyjz+7dAGBbi05FrvC+yvKv7OFFBVFB1xUNJrrL1isluGe
slWVeQXh4Nyv0B4ouBf9AXu96wS7aMc9JRfm8DCB8dSjQfSfB/5JI+Xf38z4TQ/V
WkJUdC7ekt+tppP7rcGWUx0WpPSEMNrKrvX2i+R/gaecKt9Nb81QBaC34NX42p4p
4gqS027VV+co3gCMvZlSuTbVFSexnx0/G3ahPuWmZkA=
`protect END_PROTECTED
