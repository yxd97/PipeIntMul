`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ek7IW31ftMM/38T5DAGow3C+mrq9CtUaPGw00tpDeHwjZWkGWspGnkWyAU5/q9dA
opk9gaXndKulJCGfF9wVK4mrIY/4apeG9CDIEgmq7nvI1J1qi3vDffpx1OJmeBDu
e3ApLgfr3R7WSbIJXo3m2Cz77H3RQYooYE5yCnCUX7ohOZMTWtTQY79zbijCiUOT
vzOhhMIcRArLI8gAig8K9D0TyNO86eIu1za107o4rxiqca2F1V0WQrZP9VIKwElX
95ogAkXE0N4kX8h9ljQWuqo735OmQ2SWcSCMdPMMMibZlQ9SB9PBtfVt7J9dns9Y
3I+eo8/H0DKh9BeXxdVfDrbQzo0STv5SReJn8yBjn/U+TGJWa5mhtbQ+VIENcPc5
D81BDi7lvl3YVyl8ticxukGEw/A9QegowaAq7orSVHEhV9YNW/WzWtaat6KaGZsM
tFhvSDDic5J02euotNUAdchCJIP7Q3BM1ZFDrz+uMn+rzwxNF49589TsDICIeNdI
US/o/lFLsuvZQdDyj9osoeeRECYQ5brewC3ICnXraV0fee9SIf3+K44yj0EV0rW7
qOt3FplSxYsOJ1JcH5B2ZA==
`protect END_PROTECTED
