`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ak9+F7cPhReUSvf6P3e3aSrn4aLp/BrVfkazwYvtIQo5//iZRoDWkrXPwzxEUTFq
lJJywTZq0IReT99HuHayFWSA4T+73TiPNYEdBoIx/O8/TdcIWZI41eVJ3q47NUh/
Il1oT+fL4DNpu2F6qo1mtDMnHOBV7fqUYE4IgxHnzmVb2XjncOsGjh4RmX1d7dcF
GlQO8btCVLUKZixViO4y7tU/tkQqDunaIm/uD2SpY7npWTo8P6x6HjDnsacJN53U
/gW0BSfS4qTmwAJ5i8hG+223GeB5GvnKMCfQgfr3V/Ev4bW5z2sxOjAePvcLXYVK
fzV6d5tcUzQqw4rGPAEWnhVOclfOA7HaCpveH0vZSRfbtMGfLRl1KRC6ioNrNOQy
eotltlnLLAsl+ZASyqZ8reRrnLYmv8bqVGwOIQCjCuNG5Xcrwkk+rdOLzYG7lngB
AA1VAiED8YZWTisaLuLkWomNxSBW6iTReQf4xZJA11dGPWpLL2Db5UPdy49J8fjM
`protect END_PROTECTED
