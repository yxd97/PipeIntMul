`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsXsDskSsBB7DIG7fuVnMrJAvnn05q88EMsO5VOCSaHulU21xz3YHNW732k8jKUr
qvVvbswDCQzr7hBhr26I5ss8Zlf5IHgxiIo4THBT7MzMeqTtrNDDoJXB/wskYv4T
2gWOFogXpLGlwjf3m/eDiIBaJdP8Dt9zWmq11bbphPbRz0A+c9NaV61utKKsZ4nj
A7/PSNY9ffNLVE0fF0mAQ2cWq54daMUKOPnqR8R2xdhw9YcIZMwMLGVsW8ynIqYQ
0TmIkiYQDcyfAfbrkRD93XmqroBIb5f0jTNTFxwz9ni9YPhgEPfMSEAxkniAWkXg
96ytUgthIes82sybSNoWGQ==
`protect END_PROTECTED
