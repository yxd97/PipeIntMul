`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvxvSI/SUo0MoI86jkkeacy5k500NLLtrnbbh5csIZWp6qRknMArDF9QBimTDmit
6DfyOvTQ+sVmT3JToOLzrf1LTjNhIQO9kp2S8HCDR8iAQSEFCwV2bXLdlEGJNNFn
ghOV7AKxvJKqSD01u8P9IQWNTfw5QOmM9fwQprPqYYpr+t34FrciqzAvSaQb66P5
2uIa+VbWXhhB8Q1LMDYyIuxvwerUfW8m/mXlbBhnyNdd7cJ67u+uvGeaU5le1yT3
LlQodwu1LFAKOzUBO4ZJO5Gr/TnJm3zwl2ubUWZRv52uekEWqQbSOmJ7DJbu6iHs
`protect END_PROTECTED
