`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIXRl0ivHVkK/Ck0MYpf7rAALDthLLEepD5yN8Ih0D8Js0e9cx7LRfXTdNQNLDTs
o1uQRzOa6TapdOkV/SkFtW9xShsqv7+Dm9SH4VWZDJYokN4hLgdyrwMTseP79u//
LYxIo+wfWUeMQHolYEZo+taWTUyplmTu/0ptywFSXV8QZD60CJCoYjjlV5UPUz+W
X6v+eWRgPri/TKq+JwnvKr/X7Gjc1Ma0u57xCjZbmwqAiXZ/QlNkisvAPPqPsExn
JtMWg9QzqV2tNPiPLJMpyOFGcUplaWcx3ZuF2/6L46lL6AxvxIiYJ1nacLzYoNMa
v/Cd7bfwKjJdUENkIAOaZvkH00Zu9Zhzh7KsvTACGNYUDqaTc9LU8+et+akpNpDI
IplfE3kG/UGRnI6aSJImmLKMv+/o2ZEWuG4yuEgN718hn2NFbSLSBOVw6iMkIKHM
`protect END_PROTECTED
