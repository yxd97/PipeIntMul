`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I8dCSYAJN5WIjeGR6qll7wYGlJQzotwcSX4mAdYml9vMq2u270s/ri6pGvgah49B
EYVNTWeGfV4i8bwZFfT54zUMXHcw/D/54XlwWSi6UVJBRlmvZchDBEo0IzumPANc
Ihh1JNEtxSlFZGv0N8ouCKZu2Xva9lWZ/74n5nIVtX+StFi48pewxCYWENjGMfLz
g2ep7E6ebl7JXu/BC9WrMluioRu0wxkr2bBLEyN3suLhMyCG0U5zqiy69wgCD0iA
RVrEJl1lq26vdzG2yl3R9045fJbLVZ1VVxIslpsIPHLsEhGLLmZpMK2+BUQHKVAf
zYDCQSxaFcshBuqrgrv7ciKLIiX2tQrO8nH8Hc8fuKwhzMA1Mbv37/6uK+59G01N
1XT3zGb3rQKaB8W3VPpkHNh2xRyxN3YSdx6P6Odp2uEiPGuQRbu6oZHapLUWkIrT
S5kJxCpSxhEvy7QPV8X6NI/rWBA5JKuPGCZQLsK9xXH1X3rQEZ6kRQV6z15Fk6VP
9zTdDzNTEKEY1A5ghNoXB7HN4TrUUQlq4si4A5A8wIjCCLeFUU+/ONshJ0tHd55O
wyoIYvvzQI9KZyGNLK3DTB7gXN/LYpsWEnPOA11wAV8NDYFlqnZcItVdCTu5Xspj
75mIKRoI9aJcM5tLaC2ipEk+vvBTYrzktAHVBU0LofWg6cJetnQXZY/ZluQUahDu
BvNO0LQW5SMwuPbisxMgXqFKsqP4p/K9NTfi9i1IA+I+OgDvW4NArTJO8PuPYzlN
5EopkT8fy51oOoQ6Dh0FYw==
`protect END_PROTECTED
