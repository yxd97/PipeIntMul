`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SDf9eynu0DF9iHJp9g/1oD4ETkMpW67QgkAQyzt29c/tExMrEq6OawUqEwd9K2Xu
KF0WNZIb9cx3mU8QzE8vDkQkz5LUdy9i7KyuH2sahY+9sWf7rYuHJESj9YaD2hsQ
2SsrWeGG1U4gz/X+EHgpBjMbLbSfVaTwFCZgZHZgZZsGtMr6graMA2AUaKuxCc/3
0vYpWrxdeCGTy5xQvX0HJN8ydoazpFMcMqAva1VtF69sqvukng7OzeUFEgaxljiG
qeN9zNOwMzicHiKYWBn10XRrRI0Fkq1FfBRStEfISSbtoyka8vLuqB80wBRuZfsT
JfLAVD4UiWgHDfyyceYRgg==
`protect END_PROTECTED
