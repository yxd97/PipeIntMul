`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2pq86DqEorwliDu9kPZ6UTmU7IHZapDWAWvUeMUwOls29sljA3DVFQRN1Pamrqb
Cp5ldwuaQPGktYDy/e4m/KMOIknF8OlDOmFKixOD8XBmvhkwqzppwv29gURbxwbG
HPyeXEZBd3R9kE+IRog8pp6NwoNfO9QjuRrDjmy08ZxCY04SAgU6JUCviU3Uq4vr
z0OLwoW0ZGUyrQ8Xrxgjpt92kg01V2XuMgE2Ep6YlsCUAasQnmfGh0jNrCNmKB3Q
8HAOdOAGpDvfY+qNXewP6p4l02dtjzH60q2V27WB8XRlGGYsRAQRdv1qLxOAVopz
bGekVymrOE8ZNP0jXsh6+jht/wpJ03hxoDuipkIji9ERYoJ13BVdSfCILOYyocfR
CsbavQZI3EFF9NIgNtB1MpdAMqvaB3Jxn/fg3P+DMijjtTDJuk+6r2L4U07l9EY9
tIYSlwl5pbBIxOsdih+Bkxl6lHejzwDatHBgWMvzUrok6j2vDx4g0kCohZnWx+tE
TJP6ZsHqQDsfmikJ7SKxvH3qObxeiZ5cqVqelVw5x5SWijIuxWtB9MotRPmgiqHv
ir+ecTXRmT599B46U432C7P+Gf3X2JuGCoHpyQuB8UVtzRltpVssBwTyJ7pQJUDL
F1xS1NpZKvzUW29g7WPLF2Nczl2eDpsmPRSqEWVEaeMHkFYO/088YayyCkkGkwng
QkPQpwmkqw5dyrwtYEFBEJMWOE5iZBHINi66n10ZJMTsTa7pHMTFcqWAjI3AFoHk
0+GmtA5eGDi/HSNVPpKB9ITRUOOeeCX3r0/vLrFvybRaGfgtP9kAU/NfiCNK6Q/B
8ItFa+j9HBonxdMdKMqMnRDaLtLTlMMxAEQherQWYL2Z4GgElaQQc/RMIyCrwKuX
4s3dDpCl9kabSDhFENn4mWj1yrIHIHg7NAxp9ajd84IxcZAnz5Gy/iSMSbUW3qgV
vDaFq4Bzz/kGa244lorZV5VnuuPR2ADZchArLiHKaUhnH8Vr0AQV8fIU4lIBsunO
dNn0nxFnSojIojCJSwsyJqqRuxEqBmVAjwJYK7xrWme8PY5JrfRBrIURH/nN9LJ6
2JywJwgqfNl/j1tI6kI9nKkUoK+4ydzVn0Zr7pikdqX8PeqZuLvQzMhtcs0N6hCS
aV7H/E4sKEbYvgWcYHmKrPv8e46sMwwH71allNvzNd9iXzRG+5nqshqZUtfaqXRT
KWwvpuvtGEgB8SbJdZPJBe6hE9H7vo7bw3ov+A614sAAdS/LlQkaXJIqTchj/AQ2
EYl7RsRuSPAhdEOF+8roq8JvvxQSgfsB9QgfwbJHa7gAWozyjGL5OV9yDNCttM3T
QVQIcQuv6OwbyHGQaaR1BQ==
`protect END_PROTECTED
