`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mcDt9fK/77Vr49rnMufJajMbySRnj3+q2xPXM4ZWhxLWttNG+jnHPZzIQOCimQX2
krRgaBIGtpiMARg3RQt5y1kNiSrvcMOaQhvHXz9V0w3Gzoh0HQn70G6WOHxgOcwE
XG5ZZsg7fzpPTmIiQKocoQTYqVeALzBDpkOtudKp3Jc+KDn2Rb6CKD0M4QLBjl+U
NCje82KoO09a3o+xu+e+BggAsxIH+0LIfYLJkbhpLwr7R4qaXmxOAFEattF6w1Ls
mnSFsHnaBR6SiRJ5FvgYsaNLFSynxBzF2Zmk82Ya5/52yT33mxcXQj0bO/J9dH9m
5D6BoT16wkEg6sRU89c+0I/0AwYsbaplj9gAjoXNuC1nKgQKopi7UJYlLU0GEh2g
jygREcmKIz6KFmoeCxw3sX7N20bz/sx0nEF0QpPp8KRzR465ZF7FgMgozb8eiNNX
`protect END_PROTECTED
