`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KxDdq6Vjn9Gwe0VzKgw3i6CobMI/XvieqhWkiPZ8Jjz0tThizAB5CwtZwNwxxIZr
OonB4zNGFGxfD36wGjjL5TbTidevRWHTBm22X3VOtidZdMuDFoaLMtNYXeiRAGv0
aK8sva/YEUOKcozOla12Pk5k5AncO4fs6hWGPp89tpK8trkU61j/Xtc9ZcE19ano
u99qNyBLG9tiILY/t7CdzawButjC1PivBTSjSOP/fmerZwDpSm7jN6JAO6a6a+0j
DCopg2fTIZp0XmsAeZag80eZmjhtNtZomOy9QQRu1C4rus325c0SGBPHPUG7mfs3
Wmdn+1Yu88a3dzOEfCcEq5L522mv6X/Ab1nLlRXsUi4WMByY5X2+tU+ZlGvgJibQ
FpW4XHd7lTwgXkM8DGAXVi+yitAsDvgfJztXGX/VzWwThvmqPQ2XibgJjzFs38Yt
kkVhvKTn2zxeW0+8AiteMKKlTLEEtB9H5Hquanu63QmWPcB4+vIvKD8WRcJKVxoy
8Yg8wdwvkhkzWS246wnqf94NE6+tcD9f6PmuUGzTcuSrhc9fRisXEni3a+VD4iSe
HTJNrxxyPrrm+tWpQxc1ZeySUcmWesUzjrv2mu79hgXr992Ju5KCEKhJx/89JHBX
xom6JrOVMzjM55tEqL8/v19o9VRdA4RRhPLekmKKv/hg5IZNzX3F/saSB2/KKPgs
I86mlWa2r1icbRdQwAo+xCpHxl6o/PJ91M+wKwBerOAd2A0HlXX2cyvgbtMM35KY
fRY8R5atRc+jEhQxbEKbsRuV3POdXqB4l4LC0ju3lt1RuxkbQNWdnkXeRH4ZxOOS
59J1XDNGST0ECGarzF/89/P9xjJ4054gOSoVVRrIfR9+GxMfMwr8ulCAnIbgSKvj
B/tgcgyYeVDbX6sNm7vmwRib/a94M3FTO/v2l8Bznvs5teN0PC8q80QV7cB8/l1Q
XbVpOJOQGnyIxATi0gThT9lBCnACosZbN05+Ee8YlOm/wzpi3zuuspujVRyLjfjv
8RvrBZpKSzCN4xik4f4pt4En+MT0HodTyYhR+KVQ89aqHNxGjcheR0nRu3nkL6Kl
jYR9noXLJ8sYqE9cTQHr7f1F1Te1n6oS72VwBC2N47FxTvuLE1nU3JszqUZbhnXI
S49d5Oa8DXGvSk7KJi31LAV5KLVGYiEYNPLRSNJoUri8hifhpIK017RAAQ4kWkJp
Eb1/ukWHyiJnRtskjhYE87QaDAUs03/fbwMicNzWeGPawYQ9SiKOqZq8akmEwo0Z
aHo+OejM/vU6zMq/d/KfPJTNAl0b5pe4vA7nNmldRFsjX4mQssd2AN69dl0uoNAm
uEEkRMofHwLNec9sbYsia27uckWHReM4L0EjK4NcYp60CUfZ4xOJnD+xG5aHyqsx
9sKo+uH6nCIZ//sQZtqxDIxkN56H7xafX3GhXj/z2zsVLJrYfnKy7v8jPImFinvZ
pnW/swewsv2qkf7T3CHuovckvAd6NPl3LEkRYSd/7tl6bWBkuw31ti15niDZbj9I
VPBbuNFTeT5zjJs2lJZcEAPiZ7xiVt1s9h5dgAQgeqKFhXds83IDlmMjWknVrlRt
ycbk3ojvgn5veH+lx2qJlzZhWm/zVeGm0qfF+0CninGDIZK3FgGPW5eqNsVj4FPX
pW7ujNZGrxw2wshq+mDU8LOvM7lC1irIOOJFDD2O6u1AX+1F029n9Ja/teNDQkyJ
nPadEpoVC1S8c5GJJnRuS4609OXupjckKIvRzEM5wvelGtwb4TNxYNoxIfjvqhZO
prIYm4NmFqOhJ9kLwv+PJvJllQuunlm7rUSwYF5dTEres60ojJ+6NmRXgnnB3trQ
UW+ZBeEi/Q5XUaXTx5eWCFLLs3CJV8hmfZvQEPncK7aArnY8VD17TWbmW67oTi3M
Jdb7n6aWXyWB6TXT0MNLpP12vr60qvViaaiXkCrWhkCPSmwPfzCmQQGRfzsTZSzN
86SuzOe2Hyh6hqsD0n77vS1/mZzm+OhKXs48YR1hT2eIFjarBzWqltCpWoi4iZs5
LaqRyZTQA+1tGHvFa1T0fPloorfwrfmUjJrpQVEMrsEDAHClij7B2CH/QPjaWdkS
ZYrYFUNLoEXTUjX2WaEWSiaSi5VZvWkodGJ4UCS61LBryGFpo3KwIZdnFcheGk6b
gTY6B3FYclyeUktJMego/aGdSxOUASvEUm/G9WHWQ/XRJ90rE2RjbEknuuci92dn
BAZ1eDMWuojrgUDke2gxApjv4zvOtFdV3iTNBN70QWpNGCiYh3C9DOrBt8lxX8MC
WkDE6fuxrI8YVAxlnYxZzhVVWxsD9gBsTXgaNq9rtpAS2ZXfumAMGo2Vc+QwggZt
eGFiKvet6diyK5wuUhHJ2nem1PEgIRH0ctt5+iskVGEqpWXbI6/4gJUBqVGe/miq
WC0AYzObVJ0xOuBuiqzkEEEplg8vGa3ypLZ/L+olx7kEqEdLgsfG7jjGhBrj1gtR
b7D8nmgD2AwerHWUGTp04NR5YSpxQjeSPRzkA5bvUTwfroJIU/xPmpl8MwK7xION
1To8+p9gSoGq6ymqJnj6CAQkulzJKXuFZMDFZLQSKqCbSSricsFeXkKViJT3kSiT
PEyjbVCseAhFrEEWw3mTDg==
`protect END_PROTECTED
