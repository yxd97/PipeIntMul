`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mWdKF/mfocFMF1cVe4h/rIAO4kLiXHDuUTphEC5KBESBAPE9c7b7LtoVJVlpC8vy
0sShTXZjnILSGlTMSsCXBoOHBPSTBAmUGmvAS5ZtVDpdniJ7zkrBgEVL34p5+fox
MiACIObNO97Q/5x1hzuWuEkYVg1TuMWDnUzk0gcptsQp2qt1BPOUcw6KdxKFYHMW
SHncEHvw/2O/MczbtaYJDnaLiJCcchtQPXSOX0qcK5VKfr5VZ8P1Azl0rWhKtEhn
pMae6ln7hGRz6KPOCHIbMOFN1cZg3f/299jcAJ2pC9uxddOm4+8f+LFIJpmAR+6j
FFxBp4Uqfk/O00KqxLdy+a0xy3pcoT09gYo/sxieFuoSwjjqGpxHOb0Q9uaapV4d
WbqkE1jf+n8p5PUqmNgb9+y4gDdzYl3lf/GkDsmi2hU=
`protect END_PROTECTED
