`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zh53VtLNFF6zOoMZCpol0slKkBRfhOQl2+CUnSnrnC4Y+hCep1cHp+4jWGdPIoFF
ujRIhMwaEceDTOGitM4MgXEN9RY5UzgjTakBq5N12ecy4dM5JjwW06egSHXoQESu
znnM14/e2fSLMGVhXm0ixBSlDyKLfIEbclH8WrqbjFDxTUJNxquLKC3gM4Eb91Ma
NW+niI7Ey4CZir6RPslp7fWsNAq2o1cOOz6/mQFiMvXCnVYRXfGMAY8LRTX7b+De
1IRbKaTQPPFO7bbSd6+nD9QEjREp2imli+/5sTfbuuv9mGwLfGg9vj9lwvJ6b6VF
uiKIc/Pe2TUdcKxNZdZW+BM0uj9wwVPVdqU1+19+8sdEqXQadWcRLQr3rl6oU0OH
I/4MaSUWxXChMM9HrSmadDBYc/o2Asx5pR0fOPh+HFIzILhshFtepnuakoaIfUfY
xH3fQyykP86g4UNid6mE9bUZ2l9tsE97Dnlh1hOzaeInsJqbx5UzekzzgiOvkPwN
gcnEcndDMecYOpyoPGHL2smiraZNfWtTJNfHb0zgydRlb4QDcfKajJ37oqdDcrTd
eLNhjPBFd6EnNrlv1c1Qkum0hJ5tJd/Z/L94wdkpVVIBhdhvJrtj2QmPylDH6sg7
CfrllCctK6Gg/zXDImeiTA==
`protect END_PROTECTED
