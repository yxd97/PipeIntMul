`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F+WD2C3I04UVLU2RXJeF2tGhzN4+0NZ6ndV1HumaM19pkpiktspkN1Fsz0oYGobz
RTQjXuGDw4f9pNVmslSDPpFHXTNpPZMlX8A9sRduj8p2G40J6zQWoGjSxPGQAS3O
e+HNiDK6MSZh9f9BH5+VsEMkkmi6SJMbDFzvfLf7eHmcuLDo7WoYZEqe4nqUp8lB
vyRv/xu/eBPmeBFH49eV0GiovGQxxjeHA1et1MoTQNru2D6g1wSJ6Rr7UuXnQhZw
bbREoSJDbFODilXgA1qHkPRTuQ+sggXgwSnIBO3BzXCDKVrVYUgOk4AsS8yzjHUU
ZWTgsHwV8xev3odtdbIYXnr6WaH9tB3LGW2okraSNNTA/SvXWGVh+5LcqT4m5OlW
dY6yDqwfBfgY2qxsakPCCQ==
`protect END_PROTECTED
