`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XASKWmHx36mySGL15r5f148m3MWSrjPs8foRRRaxY0MLolYGWGnjZfbPfOCtKjXq
9ol1PKW3E+G7Mqv9rGFjx7kzrmEp8D/hmL2lhSaj5caZ4kfHBtiNqlyIsJS3cmdm
PGFrE0UXGrh+8AKd+FjHWtukDkIS/7oAf4UbwVRCfFhFBk8OGZc/5UnzM6F86j2g
VAMI/J7Fw8tOpIQE44OsFZONfm90EY2wgwlGwHAch0+JLqaV+fZFWqEQ8kSQNyjH
wIVipmNH3uNmIWuqPv6E3E8QJzjWxJDDI6H3YErRE54=
`protect END_PROTECTED
