`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vZ/OW8/WJG/e5R8OZ+SsRS5RhuHe3lSnwWlUxWZrpy73laJNsbRqrfZirzxIVqdY
IfCG1W5OgFKp3SQoLE6YwCgF/2BKIw5kIUmLWqVQOsXcJSXRgMyginAQuh+IcP7Y
EDGqO1vkOhAbs1j6uvEps8MKJH/K1Gz2BO6NHw3bDO65fFM2rSLJKt26qoLXp7kf
53gejOWwHfb+GpVJp6/jw4nORZ49aZwqsmn5GRP2QY35EKnyprwnWVn9AHhlgrgh
nseq6a+7af3rrGLNJWW75kUf7d+JXUNF969c+Io+ZkBoBsHrQsQq5v9s8vAsteiz
B0s42pfqCJz5yyB04oETVQ==
`protect END_PROTECTED
