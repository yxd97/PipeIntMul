`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vEi2tG/EwI45sV2Ykbwpme77mIlnEF/KqGPfDZdBbKnU/rJFem4coK4hjWCcB/x
slphDe5Po7gi8k9w9X/RhGV68+IHBzKG4XBTNvfwL8I10RjILSCJOkgy8BYD96hs
LhZcg0DFiUEHexEM3iygCJY+BWSTHYc0l8AEj8iZ+u9b5jcz7Q8NhzQhjriDVOk+
HluP9UNUKtAXedqmtU3Vd8AiSL3T15hftYi8h9Eay2LsgB/rjg3q7Hm13SCXEq0n
D7y7jvCxCSkyEmV8O6I5Nccg9yiUVZcm66GRN1ulpVk536LYnMD4O6rC8BhXm2GE
tRP9wPiOxglv6iTnuzK3K2/voH1IXMGUYOVC73pqFNjFUGhrpghs6vEJs2hv6kXh
ylZWOYhjPjIVWlfMx9StPTTxRAi9D92ZPWIIFYhM4IiL9uKBCEVLNqegRrZbCue4
`protect END_PROTECTED
