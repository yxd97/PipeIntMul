`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tt/uPyYff0uASJDczB5YhCrR54Fb29EgTshuAW3dBCAgb4KUyIiGu1j4o/dUOR+n
xq2huQB12GcN7idcjeE2y8NEqw7ZbTVN4lQndrRAuAevny9nl5xT7728ulSMfGuU
68+GkOZJl1RMKKtu9kU5qiCto8EkcPCAj2T6edE/JkaiQOzngqvzwi58SB/HKARF
04uqkBGwTuldCcRkrQZfMPakmkccM0n31SB1SeQFDYqqONPujJHAlMgKZKvy4nhi
8vnsJxK9vEfnWBJEpT0YHb53wC4TgA/Bgu90XbGBVTdbAuvsPAYWrhPtA+5en4uo
ud3rPce+gG+bDUeeeQItTd/lEq8rCoC1Qu4TnLFOstTXzrNf/dQlvuC5uA13Bj7D
CMfQvVwrg5pv/h1YVX6KZ9VOnV3xfcrpeKtxxDRyyOrzjdF8jCNsDQmo3a5D5Ffj
zaXMd0I7M3JPELT8kn8OuNXLJg43iUYO4lsS8y/kiiNLzQQsTj0gcW935PZltO57
fGCZe3M8y7p3eGzM1p0zuHfUIPKVUCQRZjR7Qt/NjY/2f3mWpNBw7jzrDocoajqs
FvSBvVCQsvAbR3maimay5y7fdaecwd1h2NIyc496sy4=
`protect END_PROTECTED
