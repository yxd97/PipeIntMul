`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTFkiedwoRI5Q1GYMm7BiexLWTDNkMk3HY1X2wZ7dtvKKgvGc2gkI2McxOWtbufd
GRAIR71e8rtzCdEP/bXiRCbTMqradlWHwCk9naVzLCB5k1eEKXnfQgQpZwB4HVV1
sFiLU+rPYHwYY9mkLEHz1gonFEn8ktBPo7IJgAXLJeKGFl4WA9v4OA7uWwy0bh6A
LOy6ySw2qKHlB5rkQjMAYVwqvRKybgm4HIQ5QZWzuPxeV7hBZerK2QgNvDV2VVaT
Vd83Knmq0Y5GOubZs48CnVctFf4TMK1x7WwD9h+0RzW5rg3clMl7pgYXkVK8cDBf
nBTnwYRPfNzjxiADlG6hrQ==
`protect END_PROTECTED
