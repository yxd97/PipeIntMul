`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OormKkX1u7Z+TINbAwxWyEwN2oUcuVdAUexPn/cM1lXDFPLNXR11Tf6xkoMp9FvG
3axLZkwCexnFgPHmUwoBQjHhNGMP4mbTzk4oRMQem8lAuNDJWrKdQJxPKqQPWqSP
O60qz4TO4iclCGxsEwu+AQ==
`protect END_PROTECTED
