`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxNxFJ6Gg6tqK8jbGdN47H7AebIhO/UyX02bvJHSIfdetgIPXnIiBRKbIvVs4NSA
nVDIvQjxwjEAp9Z7mCSHHXNVlNvELy7y4lzOfWMBN/X3Fpw11v+1xDNzsFOgWIvC
aWicR4+GXrDcD1xS1hnwMEN9IYKD2Rc/Rpvv1J11CDKhYRGOkxj5rJRfN7xGrcBq
6puTjgONsbsTQ2AWqEhjhxwPqnM/gzGSWRa7G1x3iMRaO3J5PFM8bNdTcl0GGgxc
n6+wyxEG/PAmcx8fRCHF1Xx3nbwVbqy6AB3qoPVg2Oo1E8mzqQ0qXIXvReaG/Mkc
CoKF5VEn+hRo5bnka+1mDT2CPdyzwgDVjFOv/0wVOJ9aG7XYYfe01McfNt68lfaZ
R3HqJf0pZceeTkorQKXhC83SVwsI3WMAjSny59rm1nfKYZqC1l+/lrFZjjPHlD/D
r0RBk6nLgf3jBrFRM6QO93I2E+BoJx0wryU1W1hAIN8=
`protect END_PROTECTED
