`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5oY9rVRkl9Cp3QhjYXNXHWq0Cc9HMPbzplodgFFzv0LuRx8ge0laWowOmNFBWCMH
TxZlA5jFkGMRcE2SDlIWfymgo6vPDCn16bONGAg48vEr+5MchG5NiQ7t/Vs7dS2L
ifNBSPYyQr1QneQ/F39xVldDMIR31vgpBGwVQVIVS0H+5fRzMHL7B7UDHClJkSC4
OTgCFkCAvp8S5QdEHwNlahBDMZpQsPbv0xQbGnAzaunXeqSQS9bTWG9D02Zn6gIW
iMe6rc8xYQEvEsaEem+qRItlzTEM8yCMZCg5Lac9dbS0TRL7/P7RCUbd/BrVcBtB
bJc+haGMC108xST23vFRfay8+JCMBmP8JT4R03qwaEo0m6m+JIQDODHagaJ2N750
0fP/SCyiWFcQiPYM2xOWJahgJmpp5h8CIian1eck7lY9EHJaRXe5U+NgI1wJVnj4
otG6VDtao8Pxsi14oIwOIFHR+cT1okzDm3rWVkNJeKeL5MPq6V7DLw7ebDi5yGoA
DXPyIyIbKInxyAuOXV6RxkyDT+GW/uyNqqK30ufPTZZQ4kHMhqKPRD4pvpm4Dg1p
g7cfQo4kDUr+4LzICBagF+ZT75rkuGY4QUvLDUr25FR+ncggsWvY8O5J6PY32MIf
LTtY7Hvh0/SGStN9NtrdZ1jwH3UwYdNhydEcv89Zk2/5lmkZrq4+e5yHdoUacT/9
tOn7iypy8CCmTUvBJjpOWfQHwLe+cZ0ZZkU9VY27eFZLR4bIhXocTI5t1rrwVchm
3NN1RtvwNgG38UFOToAk9DagPUKfCc1qWnOYgNxTODlfJ8AvJM7qnS8flRQm6ULc
KArtttNqdNEts+BcFxrpBexBdV0T4xy8TbTVXbl29B1Q+7LnyJ95tnoCVHqYTGSx
LANpbnGUeC9MZMEORQxnjnMqYSAdGzASt9fRH4Z8DCkGHV26qpzkKl7pXreO78ee
6vNFGbIye1ibpKCHQfoJXHeEuzh5ob4ZZ9Mq3R9ozjYbnDWGwVAUS2iaOQYlrnJ9
cD0Vb8PGfvQqd8Y7QMzh/LaA7VfRC28ZyYiwPmRCqQM+uzP+gPz0ErX3zhBuk+gq
THDJBGMJqn5WQB45WFnHeQGIRvP1ycPDgtOEGz66ojtGnf7Y7B6ThiwkTZsh9l9N
LQURlsawga1o7Y8nSPIJEukpmBFXuC4LQxdtll1uAmlnp+9qMd0fEajr22ryqaXM
0k+P8xRfotLqKAKGCG4M8a/+awxcZMY671p7pXkRMvhLBVWLOYLddZ4JMUej91Qj
PCkCT5yrl9M7eCPoYdx3TTIBl5776QKSvj+LpkjVKr9+rVp1NTla5xu9ydLl+1S/
`protect END_PROTECTED
