`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmiWewWyjUXHb0fcwktP9srEWGrfHtIwEeZ5BCMC5RMVUd/1mlMiHl2c5Znt0GrZ
qUiM3xSGIQ3r0pC20HYEUzrv2Tc3kksyLZWSgVSyXnwS4RHJQfJcHyHMlNuKTCrv
TcSCDogUIPON7qq95DiivCO1xRNL/S8QdvWhzYfytUxf3by7F5n32XtmnH0gJ0yX
trulRGVeKgeb7Vt7WsaHYLjZyGx8BlvXqu9Qo5TKcMOx3PoBZOVSkQrM36WeSRs/
/zcjnRs9spQ1RBWlMcOFcVdYLogWOi6zo4TZaVhA8NvgNFgDmnFJe4JRr0eaC1hR
8IxCEw3EfrU+UmrO1AsiMeFlj3A/co3n3HUlIaHgdwgE9iGWEWnYjXpyIfz2Aae1
ZJu9gR/Uz77vjALOf12qY/Zr0E6d50WHVY8H7j2kUK18askXf4mx/IjBdPEXA06i
qgQnZrenIYp+QXv8zMGDjvpfh0wB0phwYlg0H1PPaiS/kSU3vOqF+yViUEiGgmAs
eRGfPeoPSLbHx7m04xnlSS4k3USySd8/Zwv9dK80cU7vjOJtohAlGh/2/mU8ZXmY
vQoTn5mGGLZyqkN3AzgeD975iW+q5MZZ0JjV+uIx/wFVWISTXIGNqGAIpG+1UWLH
rqbV1srqYyiAicvyG800+rTIXjSqHZIxHXUr+axF3KquEXM3r0aXdwDk0TLMzInu
XvE9E1cJXxcC7IXsLjs6JmT2lvMnXB9ta9jJIHwWmw62Ijuo1kobpq9vLGDaNGM7
14e5uSYaadkzeE463hDauAL2LEr/UBJjPzR9HYkVLjJGAJh9wQ3/OWkxidgB22Yn
qQ8Iqc9GKheYqd6aZH9SbboV/GF0SeLYRGVHqBMh983kP7YcElrLMyTk/iX0mN/J
co23Q8UcgNuhP8kqhTc4JFzNt3IOiLRuEy/Ha2Ubgbj8Hcf8PAnRepXDtaWzPPqG
C/+Zl6Jg/6tG/rTA6gEbj6ZTLVKRYKTPm/NjksZZ/SCX7hXvNXwQPfgsIgkzaZOD
60G2Pv+IGmMzXfgKgMxKY4b5IUlvLexLw880ttAVCY2zIsuvPLQv6eQXEJc1aPzb
COwyj5utpbadbspfKY4FzfONTVT1KFVz6ApEHadq5zYNBkvYkNqb2TIWR9Rx88C6
HvRWkfGjuVlxHAEwAz0PoZtTeervX/g53pP+KcKcPydafkHtQtBzY4+3Kp3hYPaM
HD09y/wnJV4OI1jiNhqVn767c8IKs5cvJfT8nVIRVvnnUFWdxT87nzFakni5wL1a
LLcVF3igStKU/4+LbHYMdsBX3mW0Vlkg94LKX6wqskqdaIGTSC1o3S9Lu4KeAP6L
zChjR/qi7vTjjkKzEN8o9/Z9s1Ndudr5Q0XgZp56XfwB0rRdPm5Rz5s8792mP6as
55aT85A4uRCr2+cr9/vtGfCeTov9TRs2vfeoD6gl5aHV3iWiG7KULjpLQ/NCBMgU
7v6VkBIHFkI2x+pMyMVVanez5zVYrGjtFjDjQkHBJgzsiWrrG2SHOOlmUHA3RETv
+Nbz4Yxoo95sV3HZBEJ4dxjHLqu1nb6sItCA5m2dFumh1zoahglmK7dqD4Io3IMG
I40eeSc4MFIARV/vPCoYXCgZOvEIWvTSSTVAgF0KJxnaz6c96ut59m+azgCJI1mw
ygaxEeo7OQdK+amLTLNihRfS8GvueK0xkUjhAECIqNL+Nnxtb/XsKfX9t8aDq/U6
5025UjiJNRi7kI7RfYKnyzEKyWVy5qPejwvfEC/fuWKt2S15Uwqo+k3Wq6SsGdkd
9QRnW1c8DyjvcIBJoC4AbdwJe1K9KcRfPDtCTb1K/AiQ9R7wQZ0L7rZgfcX62pKx
igt54GfsJmyVzG/wvG2ltDI4VG5AHIe8QyUCs5G3psbwv8c/Bc/AJk5JogHiV+a2
sIEAoSxMaqJ3Amwpo5Yw7PsyMATOT8u9s73eLnnrSPP8tZnBoR+Ov3YnzxpP8khi
wNKPHdrHWMBHjsJudrJpvrJvarpfl4nBInqS9Sb0PdGL/qYJiR28jmkbyQmB7GkD
A1JRQd1WylzkirttmBlyL7VADoCSZHuX54WA3EuYLuRauuxt1zKM9SsP3z28VfJG
MLnhpskAWxvaRIUBujsP7wziXwONU711HiIfsk7G8By1kc6waH2jhWOSivI5aaio
Dy0uQAloysjMEGb2gJpBA0cIOcPo1ugZjxw28qygO0/FbJ4QDbUltxc6nPxyV0Qu
eKJCnJ+rO2r6YYRuTBjuSZKbVzvCqMEIE88CHV7SVYThMDysY39bro1TayEZnJIu
M79Qgr7hUk8NxH1OVCM1gPxxKfuiiecHauCI4ZYSRqcr+SbgerGCfIdr1zO7y85a
KJjNc7kBwe3t6/VRc+WTptC5B38qpOgolGcrPOY5r4VEjxirscuxcAvw0OotaCIr
wS4KIKS1HgeCKj90V268kRVK0+yVY7gOwyzXcfCKuiYw/devVqIFPtlgExnBt1mr
vfhmUd8Qvnp7AM4pjHipMQ+440yXI0LeVH29f9axeMbuNQaNZ64k0bMzaoJr4JnS
ZMrZexygwiFaJeAOBZCF+ZorDlVrR/UVp7hYDroDa/XtqZDPgvNeLYnUL8savjXb
ZwLDBfqHCnd9fAist4iXUBHR2xYZ07Zvi6aJd/h0HGUYQr2yH/g63Gb1BJQlUJMq
AuzlsGBLoxRnKGfUgbsYz6yEcZibkqbIrVKxLof9xHmFkKXAljkmn2I+wgN5SIM8
G4OM2t6VUPApJ+hmaOk4luCjiDLK7kFjfkPepLHUOuVbq6bEIFEyTzCSDQjBRPf+
y8Al6ZrdFosK0nO3nSG+Xe3mRTzzzaQSlfVXuw84ThbELRxT2h+TdxLaLiBuOjIC
cLZiFrCgm104rR/meCUoh2e62eVu4M7kG0lYPvOWQ/E64Tmid8mQPMiOUPyPsopa
KbPwF8kTEoEnb+tREz8/fWuMuz+j5lz2sJIMnPpGPp/6a3R4+iEVb/wPzoSKzk9F
aFEigdIpZfBzC4+vcw5BtXg8xP4WHkGDyGDUh9hsT9B6U/Zq9H/MsaX2slsGyJCX
UcSGfCTvn20GAZUn+VRi8oR+FgMP7+Fs6rNmFF7v6f5htPpDF+8XtBIbOVvxoBYz
SWFEccmpookV9hg+WznID1I43X0Tnyx9KArupZTbmyOntkzojozL8ln6eSoLu+Cd
+Tn+S3No2ltU+s0iBlX8XA+rd83TO+VFOPyaKVUDg2ELyMcqjM4XunGG6JbWEseM
`protect END_PROTECTED
