`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7SCKG6uYMVvl4OlGdJaRWSGPNi7D9AmEKdNEWrnngyWqVps4con6j8TI8BR5EFJC
sNYd97Mp3crh2ZA9S7Ra1MhVZ1yadedE4OUTEjrua5WYcO7LPU1f9Txwx84xeoGQ
6bi3KOjl0GEoIGEj/0jhip+WQnI7H7cyBg8/UlRx5v+ObltMOClr6EpP1efbD6E7
Vvl9omIV2kwa14j8Y4S2kz4KVbBqB2btFjx/nEAuKOHqh7Ye/883XvtMLL9y7WVi
HUAs6jX5XUMQnrzxFmydNsQ8Q0PNlQ6ozY8sgGoG4eMeT1x0fTtrgUHq6v41YFQq
LXiS3Xl6VajYFep+hB4Z8ASLG9I3JU+KopJ1jLDZN9/63F9N8Y4DNdYcrzs7yQiW
RqtiDVTw1sQI2m1Xh8W3dyB/qYzUoRNY5V/uHPyJU96z2yKot5E9lF/Lgp917geD
87/wb5dwINVAsq86QPYGvMoRVHo9ztSUVPYhSmf8mqMoJShmpHpuXBfdYecqP7nX
ElUncngR5H96F2BjgFYWJgsb02wmxlA2XBZC0PeE/96V9+hYs51NwUS7YPA/JayR
sxrZu802edvaLZ2Gn84t7nnJOJAUkkrkf89lkh3/+Se6BWzvO3rZr2EEG+sVtjhU
/BvNH3xskzE99AMKHG9TX2hgSUVXYSQSgXkoujJe3TBuyCMh6kduvNd10tGzpsc/
vFJdUYso9viLR3CoxOPVBoUR6d95AUhfee03Leb5kIQ=
`protect END_PROTECTED
