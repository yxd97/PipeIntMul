`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMcREf5NE08NMExR/jx9mndo4GLcTobBNYZ0nfhDu3A5BJHZpaxnWErJGCyELIR8
yFxSckKZr0kJgb/sjBzzL5HwCmwdKO86v/qiqeWu3jubUA4c4we0sloa0bucZSBx
WqVWCIC5eYZg3nQPZNiaXPZ4UVeMxejme89P05ypMupUnBmMCvqkB7O0tespF6BC
87rFIChls0eriNI7Afphuvi+zWKoGULFWvyEFBumxOPU3ZviW9IS/85odLSvMUnk
DUPaz1F7bAKmKzFp92CEUX6z+DWgcWCob898VNbEbqJc5fS2n8GMcsw5nnO4jxae
r0Q6vJEbHsbJYCq8Pv14I1I8paCX+bTqxpaFFTq477Ej+9QQJvasFAzhrha5AdO+
NSeciHBTVPGqLfajWY+C+y2De3PfJz+qZ8yh4DXNMD8lvrfolKYqyACdsF937Qsq
2aAWCo+qUi5CtC42sOWLRKRYazcympVPSwXYPeHn3itUFSBc543c2FdG83bKbq5i
D0Yfp5Pntlc38mabx0onrm9UTFcCw1T671nNM1+V0UAES4Rlk4mm/UGLQ0ou0v19
cFufMJ/NUdl0fq77SSOzTRJnd6iW170nZTLDVL03TvISshf5nbBSlndY6Gw0q3Zs
vXuPTpr0w0Fo9xRKahY2SL7/shvRAhzwHJDHZU6ZHzX7NOsa3tgqXxfVKvMHRWuM
rePoXiVKBL97GqEEBu4kin5G5Zd/UwrJ8ZeaDtWM4U3l6INt0kJ0zlMTAVWM9sVK
WaUj0Oj4zePgq+cH9hzt/73KFSY5t7oEEljN2mQNQR0/Uhk0pR2lucwde1A84sRL
vAfslTsGz0ZNz0jzw8sS6W7EzNH1YGzRBUipHzzLVFXDloh1054HTBzF2nVhHTcZ
cptYUfV0zj9NiCWDy+dBtEL9NrgITD6QRHVTGQPZ8DNTzK6qukoSb3op9IyHWB0b
n0MTqLDuD5EwD3xHMun4/jshrDpPsZgk50khppx2YqI=
`protect END_PROTECTED
