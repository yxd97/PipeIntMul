`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bC2evXLjkbKx+950eti29MiECDzU+/3lV/lWQco+8Aa1E991QcLjRbewB83Ke1+I
NGkFDPdzWBPrGsMvS0eT4KeQXKDKetTich2o8H8Qzo8ef08W4p9/oXoMMTuvTxc9
pLKtmwsuQbOHqLrJT9jeRRCrH9oK+8wGPVLZPACCdrhBC9hPKJBTnBhwSV8FrAdc
WjCgHtdIW+3Q9YmnBjFSpFBApJIwpQV05HId63Ddxae+0IZOFnIBb4ArMpk64MkS
yBD194d/DB6MnAny6OnY55SkwoCxaJjUiPdY8+wtv+iJsDkQSY3GjwM1ZrIz2boy
c7OpaTJny3yF3NLo/YQ0jokm4hAY7GjwEmI+jqMRElTLkMZOdiUsk0mjB5YhYa0B
/JypI8E1eaVyI39PxkRCUESFT2VCfAsdTSAqyaFViXfBV1f3gqTB+6CvYFd1Hx+E
SRrz8kwhAPNpifY17GfR7KqoLj7Lj/undQZkqgHV+TIhUO0tACUjCwBs1YKLzlve
`protect END_PROTECTED
