`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3OKwIxZBLjqJSz/R7VbzYWmFnNaTeOF/OKx+K0oFz1aEikpCkdyndY1OkYFcwa8S
Y1ChdZ56tmNrbRTVvYdIH/gBVe3qPujuQ1PlciuFcp5/mtjyQkc7WSdnQwo9AdWE
7PTdmxaxEMF6RN2NsvcUFRyOit7TgAQMekXd6v3wg3A9ZiB3SXheYJq1w8A5fql+
yspD2WDFUgcbGouXIlUi2VTAULKQl6Q6m/E6kRW6/+NbzjkmoxkzLsAjkBtPLfBd
jUaXB3pzVC/HqkpD4pjboREQlXT1tTw4UUd59BqdJBUz571hUdbkcwjP4bv8X4R/
GbNqztj+w+R4GQqkGCZuzRk2BbfeZCd91sfT2YULedBZd4HcL6qDzwhcOFnPOvIf
QIj+K+W0Xadj+oWAnUGj1Wff6ci7Xyu65rcwHTHaAbISk0F6TvxUcx+OTv43XKhj
3C0/f/nqkUOYk8FqU35IS/rMDUAeh4E5jRmZ3Tml1hZnNXWtVo44l14D3k1dsKaG
nCSrfFTfUsLPMqo3ZzmGTvl0MyGjNk91K4GNuTB/jBCPHiMhSgBRNZqgBTnot91o
BqLhbkM16HLnh3r+7dCJ2lVuWRo4ELMD1RR2ICsGGEWPBXYs9E5cpU3bTdLv73la
`protect END_PROTECTED
