`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5HAyJiUa1OzAjh8ieSOR0YjcZfGk68pahZ0tQfHQfJ8Szu+I+muM8f02gzAViMG
W7xtGMwPmac9L6nWj8H9rid6hrsJ7YiC9C3Bbg7xjxS6dtzjl76Z+InoTfyzOg7h
6BuQbnJazNoKrH1ZuZvXAZqP+VcYVAUc7vG2U/NetOgs/TiWGT1Mx0Pq3nnNqGhW
06DqW7gLoo+vrQ2AT4a3rPrEgdcvRyE+K+MNPiKf0pFBgZkS68Y34rIWeSXSlJpo
FqVe4k3ch6Ch5xQSoqLdow==
`protect END_PROTECTED
