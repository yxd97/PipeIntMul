`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34guftLhfgRYxcVEGSLXgJjbxCnfHMPrUVb8kDNnv3cJeQMeaZkMiH4Gn4QKNBBK
Y0CZMkb9cmZzge5d6R1k0AXgTy3NkjUvWu+E29PQi+9m5Iu2DaW+rhfr3pUpdIHT
T54SOopIFq4VdSY5JHs4ofXYpf7mG0TypUNeIzIbWByBmS0w4evFOppXQNns4AXt
Jiw7uMZD6AqHifRdM7312C/bdr9n83jVoBLHnzfVXCVQZYNyLgxBjeqZ6OXUlf12
0KQWYLvkF/BhOtUTziObdSEE2jHFmw0Si7VPOGSQQow=
`protect END_PROTECTED
