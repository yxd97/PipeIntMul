`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHoYWvwwQ0Z52kF9DDWSxJhTFwHP8JiNhIwEqdTH7OYhxYhZLA/qEKTBlIk848+W
VL/sAhe+zghUjdSX3whubr7cZO0ywEfTKXnqo9xrJ3NVmh6WS0lSIkTsGU9/Q5YB
GklqpuNtvFwHOghT5RTKT02BBDlTpQoT9MISXgSWxcZqSmTAroXDdq7+L/NkmC6j
Gnub+BHCo7c+6E3WiMqSkutkv9XrBWkAdwXbtl+wCXvXAQZtk8O12ASEwnoyJqEo
K1Tggbt95DLTBPfBwnDbHRzYSkWkF1rRT0nvxcoFA0iTja0U1+oTQLin7PFSCxS3
ezDLcZkKMBVqdWDwasBNJeV1j/HfEtKFP2MQGsYWgjcKHApAFxjO5nXU2Sz976qx
2VJkYz6m/W+hZRkxWew7I4fBjndWsowE23n6IuctxuoC5dRbFb6BZGz3tMb/1OVA
sBFlQNHVDyTxPG0aSB29lQp9z3bKLL4buxWQ1lhy8pYEGSvJDD++c+3NIuSjv4Ls
7c5884fQuAKTcM0xu/Q1a8ncPtK5Ts3JsiVg6nN7YOX0OoN85Zd3596vBVGvYy++
0rPwdPzJ1w0Wsn8CDVneOmMTWRMQq9Xsd5djwamw8gQ=
`protect END_PROTECTED
