`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HoLz+3DX5ggKFdSfeuLPr91wx5Wao+M1F9t6P7b9pivJP81FsP3pZNnbOOiobJDd
D+2EWc9BSi1tx7/w+3mSr1CyXfYh1Ei0N0LppdaFTV8dY0CV72HMPsugxZgEAch3
DoKIn0isV6hlsztZgGpwWFR1hZeCpmao/y52f0mVoHEI4OAB/cgTo6XOHqJs2/hp
K2QOKoMjQXPNNuEOWE5b6rin/lmyTrqeZJN07pyFn5gosZwdfBSQq5/EOVRN4tZs
YQI59h97ymRjpaXZKWsACa3wS+CHPShhQFX9YkgBmrH+2M5mKVcSJPq93pE0/YVH
t0vIcQIORDehIxJVpXJHAHQVF+F4iMLAjNqWvLEuMAc482L9Dd0pUzeR4VORYJI4
YjewZS+YFk2u6zSJrv6Urw==
`protect END_PROTECTED
