`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y7nsGVERaiP28hHRFBv6RiADoxtt9GcPoWwyBTy84CB979EZJCorUa8hC7xiWy/P
f3c52pSNQJNE8kuGZb6q0OeJVUBrLaTAbZUnJAaikyyTHFeu7BKzMFTkz93WyqgC
WYEQ3vAS3aZKZeoOOqaT2p/JblKqwf2BCunXXVTMuY7BXGonse4B9DSNYnWSkfuM
Ye9Q2U2j+AtwjjzTjnpYDQ5bN7c8R03YaRCMk/m09Vdo+N6jnRFFz27HolQuKqvq
/iOlBSzjWocLqiIqO2OHvHOZLu2vCPVsqBgEtIWmOmz7U5QgxNK+pFE8uXnhMxqf
P5SwkrfQK6nUUHbn7mMirpPXRAVauMQS30z9hqdWV3ULUmWAnnjQ6NA5kVugTVey
VmvyZp3NZueNBtvavzc3aQ==
`protect END_PROTECTED
