`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wl+XoCHmxtHlZTYfIFQZKcJ14jyD9UA2aaJDBpA/NJeaCQCmychnLaj4bGP0xyVo
BCIAVgue3RDHN9uzzs0cubc2TpNZ7a6aPESnBhTIp5d7uMJ/v0yM3kKcG6udGzhT
O+V+QQSR5UmulJASphlQwXFxxnGZy3IQb0luzgWz9Y9fXEIBolpj392L122g4ve4
GzN0pqgxqJvjncopinAKgIRCtbnngB9QpvNP7qykAn1omldOW800fB6eOGLuQipV
1SS2R0nFZjhvHaDD5w36UfutPuYshttZubSN8ItKVAylcdY1ru5xL0iH0Q+q+g7g
GWm0zlXxyhACQQX1XRW+7cqU+ZCOamKP78clW4VyXzCoQDNHsWmDWoeh/AB7Y8o1
lM0LsY9nCeqrJGKbC2e2WDkNX6qPMZnFY+gsOIeuQjwQN5vIwBLVKAE8vZx0atwI
mtMImsFLoj13XwYfqS9ES8tjDM9ii/eUm1BPkYnF98wNPHWzb43QglTj+HF5RBWS
jF9s5vlKopfNmjQNKhsILJZ9gnWBNScsjYZAv6C4NEVhMJDiOLkbbVs5wfPMaAop
8S+7AHRLeuYXwFJhKq+UnkiQrRhqkz84eGRw7lSP7LneeAkrnhxCo9fmZfPJ7CQ1
bvdZlLgW5cWltp/HepKouYTPTnO6HMoHfz+OpvVrv+CgHjkCgfR0z9q5Hz83al4J
52EKRfHo7Fgq3u8uvzRPm6hmuvJWwL/Efh6AhJsSoHGDZvPHJrHAd3wNy5/zPgUS
gXwuF1QXkWIrTx0K57qvJNVRIbSwHxwzr1v0UP3Yg77A+UpMYpi/pYJk4OfU8le4
yHyuIbFcwr3TCt3LGjRmaw==
`protect END_PROTECTED
