`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sf7b5SJSv36Kf/PgRAP03Ct/KpYY/RipgAypzdWotwLd4dNEfFc6HcVtG4+RMOdw
/5wfHv6gt8VP/hMJm9THFtUB1dYlAKXU5uLvPeR1VYHzqqQHEsnn4M45TSeoeb13
dEHQwcmkMFrzVk2iau951ISxKpPgIjYMaCsTPmOGQp3ZcMhoh9nQsopTjhHzV/me
PKDeLAxCq+dtsMDMpG8Y74KIryhLHnbWOJh995yzXRlGhU37KBo7X8rsZZooPUz1
on3R9oMEo3z7HM/8GUCuspX3ls7KrA4EH1arYIfQ7ChsGSnlvhnT+wPYZODkAD1I
rCscaDpZDq+Pk5SuUlfFcZnoIKGbYsaRfMkiw/aR0FSRycrygpdWpAuxecpNj5Gm
skoc5dM5/w0OeabEQT5IpzwFeQwzyBXPI/oCnl9FA1vMEAopNgDKp+/RqJhBVFP/
yDRcGyQqNw3/YST6Asj2qQ3uWRpBtquYrka24NhuUuC9WaA1gknXQRMVihA37hQH
fMyr8Morzh36j2QFMZhc74GBVeB0v0r9jHBypGlBATUKK1mn/XfVAvQUcKnR3ztG
GZ8VSs6K/XET4fLDSvL2pjdx/Bz9VyqRV0MHjf357UQrNGtvJE5agIFcz6TW4nSP
qlOcRzcYAn/hfbT6Ho1qmmCUt1tNbzQBnl0UeguVQI0SRrrFJyXleE527mIcAWne
A19xCmM8jYivYBcENAhce/9PcnGBuFclkCI4Yl98K2Bg6QnqvqSNSmU/EYwgMpw9
6KTQeTSfV4IgrXebiSTC6g==
`protect END_PROTECTED
