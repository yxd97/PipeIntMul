`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ofS48FT9qfhfWuUfQEbuCPIrtktbJkRIPWEIdmw2VZ+OoajVmyLxOjwoJp1JEM2C
Xa6LmfRuEQnIE7shzyPjvrZWIwfpIauAS0uJ5lYjYG+GtvjP/lyr03HspUz4aDHz
5KSoflTaSJmSYxS28DBj0Ax04MQE9WUqsmpyy78j38VpqtU8r2pIXr9SL6pW7MyY
+zy1hyyb4fyJQse6O0bUQtjy7wE3EmrRmoW2MaxEc0Rqa/X8M7oJKzLpwnlOmyfs
tZiqfSvTAjwVnmTVsmEu+oqqqNkwwltRyFeWRJmA2D9Cxqy3oMIhuEHNN50k2qV4
ALFV132HaiYwKXhMqMJmPqt8jp9gyX1DrKjpDkfb/+38bNKdk+VFyY5Bu9iniOs+
3W3zi5fRGj4CwB58Fb5QjWZYgTBgZJ+BwAj2+xu/9B5IUWE5LcaF6/uKn7ZsCLzn
plVB72FL7ps0hKU8RHw03bcTVXbm6pgOfA0Fj6kqQOR5hopVKfYL3vRkYsXH5QWH
PZ2B29rCLjanlZOeFFs+m7CY1V2ZgwbqRS3hAUIpryfGn5fA3uL4h80FVaEvHevB
0Qq38kN+ElpqxuOVkq85ERZKpquNYEfRMK3eb6dae71CA1juQpc1+YrIU5/zWW2J
l8ApC/w+zW0hmEgaZh4rDMzhd1ueyDZuwENIfj+NBW7OkbWPFTMuyZPJuHIiMisG
t//a/1kK7ddiaeDjBKz17CYO2vuG8k0xQP1frb/5Gmg=
`protect END_PROTECTED
