`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDK9Vmn85/+rqHOna42UBBpnh7RtuzY4altOroiJ42XT/P7Bh61w6vKIJ2VA4Fs5
Xdulh+vn7FzdoEcJFtNcoKmcUJB1hv97HvcDDutWFDDZn5rqtuUFTJHKn+H712YA
JRmyBYyHzMmUR3tIYDWNbDpW5VnSUY9H3yBC19CLkOGmddbER73SAjG0iW199Nr6
Er0pO+gYEI9yXDQ7OZ89fbC5eAIl4FrfDPZiyN9QATAZ91OXnMEXl0qVItxQrDTu
z7vYHsDeicAVgymfgeWdieE/L09Ykp90g4J+DddSHTJZoOtjoj2WLpwHGDjQsURd
InRA5veB0asZZIKlMstOBbjxEajQZGUVK01ijrZ+kRPUqvQseoKhQt1bXS2sw6gr
CBjKXsPocT7wMTiQWw8OFFypPz6/X6PUodUW0qu+mrLe3CkOZxUxQbkxYOwL5M1T
QK4f2vtNN5GIMIDWkt3zuhyW1ty2g8JEXjPoD090APuNn9V66C1EbWpb6a665TQm
BL4ZNfgWspxD8oXWvJT3bWSXn/9yCJcoK59StbhlPUZpEjh7QcFEex5zdtOAmV2o
X6N3Vh8m8xHBsKICCtA7xiHub5pGvNbIFDPP2gSrN70L/hhN7vF7F/xabPNk9mie
GwLYPPyHFGk1cDF1Kw4KzMUg4gvuLYPHCcD0I3ngWg2ibnbatrKhJ8R1AIGwEifE
11s1gIeTL782PSxjdbjMWksXg15b+8EX4of3PHoNcxMNAJMn3mPEZriDZwW0DlRp
u9tnuHp1yku3QpeF+XeUkLgo/8jzAVHS6EnxwQc/phwzlQ2OLRtZ5K93U6BpFQsA
`protect END_PROTECTED
