`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NNZ59T9/sviNXSP28XYHdbpMDW1SqNGBwYPtw1dRn1ALGX78sb2Bxaaj9CWfy9py
9Or6es2Gr+1Mw6h4wzaSR0m0zAMHRLX5rdQ9atCliPJ7R7cCSirKQnlqSHudbL4j
nVRY/kBWvwsH/MgtLIkw5svwhZpoCHYm5Q85bbL1DeHMgRfKQspTyT0wmkiZeoxF
Y4zADxUv+SZ2XDrk2wlmMLpcLerBGrUV/xgSXQFQ5DinHXc/XmlvaAf4ZDQARHqd
QQ/sS3gp56nkzCb4RqbDTD6nrwzQjdOYMmLrepRos442gBrMluzPznYF5nwYUo65
Fp440TR2ebVS1hzzHY2J47NaOKcZUb1k0pPwLBrX3Hcl71IiXlj+StLR3qYjYoEN
zlV5ZtjCA//MQzh01l1b+L7mBrvQ4jEbMUpK6+ED3LloiSlavXJpCMRMQRxsXYDE
fLXUihpE7CGHdMoDB3/L5RieP+Pj3iOa01AEYOlH69yZ/WxklQGmGgypf4xjuT8v
MGDV+sGpP4ix7T1hN4jmBkhJydAyzl2Q9/45ltl84ITRSxbAANrK9XxFXuXnLIBu
pX7r89wigRhB1O2t3gscqjKorqUWrxGJJyrXsyQL0Gw=
`protect END_PROTECTED
