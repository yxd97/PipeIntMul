`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vUciwu3PqV89XxhMDbI8qCQkomPDXuk1CX+EyxJe1tk4NakFE/XS3fN/ALGXAfr6
wUoi5vMEbGUSnyAOtPF948B9IT8y8ZnKL+Q01ejFv7xM3utQvIj9weiublMjaZmy
jyTsUAIOHyRH0KSuGCL7r+zQWK6LykfSoIQRIV+AOmYXpmhrMxsKiZpinV/5T0VZ
Dgj27I5iota0SwBMAK+tbiAkg1Lv8xoUCmEzdyHAA26KBPdyrY2DdPpn6NOYCvEc
qTGK002Kz7ghbE0xlon/KUhQQRQfM6rRQM692ocyr0vgaJoUHm3RRJyJSubJnpIf
OvnvOHTcNsYTF/yWZnb9yyFLcvMof+Z0lWgivwG6/X8El5WlnFqV2v9cuuvhAALc
IOj0Hi0hWLCsQcMWnOXztEU/t8uFCooQCWTmrcruwYMNGDtQoTefkMoiLNT4Zgpz
VeTL15YVpFxq+oArb7FyrfYZH5nlct2iLC+TIuAfvLpT/NlaqIg4FB58MK9ZoF27
p5+jM9IexVkvk3OSiqo2q2+JeLu0CAOMTvX2EwU5oTZODdMF/RkTj2sLJNZGNEim
9/5O0IUP3EZ807/H1ls/0x/F+WFFlsMF0ajWIEDsjhVLG3Suw5XOrGymoAVbZD88
8rVAfvRAePba8tke2D9m0w==
`protect END_PROTECTED
