`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ozx18sA5cfrnWlIaE4fhPK+lwqjxJEd41j9y5mT6yo3IH3Iix5ioQoWu1/XiDJpt
dT/p1jA0WU8U0BrhsG7PUz0VjyS/wcW/Z+Ki9TdsiTbTasIfaOSrRl0gsviwHuTO
mcHOCpiCKMdRcYkWo8JWbk1VUlU3Tx1vMm5N/glI+SlnGsRLt2ProwgbgSrEefMq
Kq+R3g+BFBkpqqheoeo8fq2n24LFYmq0HoYxOJTD6G28en4rf+QxSyC4PDhaNwkV
LGWhwnt4HH+Y+NG3lwuZufDSWRcBSD7aQGo3n9DVf8QMLB6cC1zf63G/Qs5Ek3Hn
F3w/0awK7x+0YGNH9EPweNoKS3jY56H5wlFmSnYgDsf+cvw6yOe0a1YhsCG+qrEG
WlehA27Fk6VucXUleTsUQP/NYTkNwPbNT1jBhOuISrBVzuz+QSPR0tC8GDqxSunS
IQJZr2gDaONMk1GLf+rt8GQh+dASRjzZMUoitFU5W0PU7IuAuNRUiodOt0q2ZHTq
+3EFV9jRlWxHKwBH7QVU7mP1knQki0B/UrrxssWH6o6RwLXtOhZMToW/tcloSJ6V
HucB47QP9QBfv8rP+7fyfeEQX4tQicF5kGwveO2Ge1euhJ7ElqlKPAjIwkEy6bp2
MqybwFSFtYk4tYg8zHalB8b8fc6oPsViC37cDKVo3yuBrLcr89cK8I3EIsltGwGv
`protect END_PROTECTED
