`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQfISUsznJWqyF0lgTdvk8aIKHqEDVZT/U02cyTZVzt9mlo0YIfPpggx7y+pjXwW
p/e/Nx4yyaZ0UGvVxjooRukJ66uMftJW8rdfv8ybm8fXOzP2g3YpLwCPe5rN1b57
/qrVPmbMl2qIc+xjn8Sw16ZYRmTcC45dGpGLQ7IMUik+rOvIugstwEndf6DnmhSm
1PpFvM/x9EFwN+nDfWitivKTzEmJLYeiVAkakJzVprDFe/83+46g0EgRX7QKitHs
v78uBSIgX/d+PBiVIuhAEhPRRwinEvr/APHtm0y79QFqYAoojR8N4g4sbqeTgn/H
k8OX1Qjvk+jy8UHKV+uPpzN200CYhgRjaEAYCn3ya69JxYGHWBr8hensOn1omEXW
pnIoW2ui0g609yLL1c3tnYFWTjlvFlhq+PqhhT1j67PiBikWwQZb1gVg8eqyyxBr
bCW0OZxUmmjcHGZ9SvORrTY8eH8m5asfafqSiZ5KJLHHvoXtQZkQiz8Ccmi11BUg
jarUNjD7CGX1Ght0Ls9OGb2YU1rjBT+ddEjiMdmdG4Vt3UZvGxysqgmimzjlc8nH
Rb7i+po5cNQvzQOZFLptsKJrRtvaACITsRLxM2JUc1gO58r9uwRJcM8uutifyxkv
tqJmMixNGKF8jxejtYnPiCHM03nRKSKRnKgGdmPy0pSmJF7M/XQIlSG5INKvLKYd
CM3QkDxUJg3ZkaX8hqH2T1bdAsVj3m5r4zLOdQWMQY3/J5OET+KdnmecM758yXkW
LfH4ZVeSAKeHF8i85DABMk9Bm72AlAWWUtNGH/I9OdqoeizFrgPMAO811JoxoFn1
Lmmu7SLhgiek7iIJbztTAyqhnMlO+ovaWTHhxtOx8ZFMp+bhWMT0lBlfNiehMLwq
s7rzP7nzXKELoLcu1S3Z2Ayrz6lizLfY7zQ9gXFFuyMgNQRH0c+a6sf/qLE64AkA
bx2a+aylyDTr44oJO0/a7uLxDa0gqqLzbAqpNyNjURc=
`protect END_PROTECTED
