`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JnLOws5hAmLDy7BgbnIGE4gOgYA49hraJjRKaqZP0kjaHRjuEWOLNqGLnlPSP+mb
EvORFhh1OnBt9FXnxDZiMR/cI3Jt7jbB2VhRnYMS7mYxG3AiMXi7ceb3HL4uJmrM
ofbSR6DiBP/KfCi1SaCeZ99jwzkxWEoWjjyguKWXgpRXMHxCPL1D/QxMaQzgP1a5
IOurRUcTviERI34yFL400Hvqk+TLF9MtpoOlcIJ6yoMCGlyYfVdeq76YO90D6RsJ
HGYF9rjyRzHYpAwPHNRRpN3Z8fxdh0gt0KYUZGir3x+xAN/SxREWopsDYiJif0N4
tXo+tDkw4Q86NmsrZplzjcIeyHkLwS7F3iKJ623w/lNL6nvRitwiOwFpvMobtLPe
ooBxmqLK59Xh8irVN0bOn1UJfX418UbZQNuLXb6JomN5ojGUooU8cbT6OBgeJqHM
Ze5CYYcW2NIKSTD/1301I2LqBiHJ8fOT0iWokDTUG4gtDvh5cgOyUDCSj+UZbdti
MHklb1DrSq07adHNflLDJz2QOWhK6SHmeIzDlsUmzEwFlQYtCY4JmTXGuQrz/PEG
6OHuyui9F41n1BIoyCD7Hdt+Qo/m5Wu1PV6KmvFnV9vlqQrKCLcdgCpeleHA9n/u
jvdXct/ZxV/6zA7iXc4R5A==
`protect END_PROTECTED
