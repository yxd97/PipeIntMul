`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yGce1m8bi+p8AY20FuDwCGpZhySKorMAgdaSQwxcrPsw68Y1pTiaNDs/ChEOctib
5zTTATqQqESsiGk6OihNSFYNzcvmUMEx2glOxpJe8Dj2wQka3vq3XMLaM7rgSCRy
GQV8CAaRWrxuG8LTeePiYK56faJsdxz9JHL3gxkkCKFUdVrxIBLxOR/sTovyamWY
8l0qhbZw8CkXa/iql7rn/rQNYMD838VANzIP5gqAZGb+nKf39CQgGaNRBAR59GCB
YNyCW/se5HWJBXefKp5gTOngxgwGtzGrZB36QivHO6yQaKNbdEr/In3KjkXWx53V
WTfFW2U51DfsbibT1UOHNooDNH1bs+awSJcf2tjcIYkliQsz9cLW5Fm2O8Bz7SCv
zZ9bzzhoDWLXxS43DN+DGSOWT70NEpmrTEUSnPnWYJdVwPiefdRppHfdnL9Ltl5W
`protect END_PROTECTED
