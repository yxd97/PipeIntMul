`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/+tbseJX7d9zeX3KMV9UWp08vimu6nYuNYODXt8WiNNfPELxwRItwe+gnPPAz7x
HGKksXyAeZCX2RmB/CbqHORqqerGyNP0C8+dhPSMmC7v/ZGpOuWaZg5t1xEImlTE
srVxJli30LkMjCxy4o1diN/Nl+4Ki5R5Dp/3tUafcR0KFMF8HkSMNqw84dADF3t4
zt7Hd4klRU9URZvTLr3BGA8xb15hj0QMP9hmaCvo7T0ahMLZ6zoGydjYJKdXEZmI
GQKgKCWTPfWmZR5ENaVN82X8RRtDE2iRuXxVwS+VRZZ3ORtADIDB1qWdscKOHoFo
pNrARqRiTDN1BdsEoFJcpd6LMzIoKF6sEs5jfGF3LKp3gG0Z6Sn85d9+nTDUSyEI
KYWzMiKtnUWJPFc50/O5A+gWTWL9YSoAhlf5yQL6a5DAnVirgKN4mVd1tPFtMhly
DCGGVKESzjBBLruXDdBuTK9ulH/uN3NPMCkIxmOiP+rMsDL2eHkIS1WWtQCrA0X5
RTy+OetQPhFSIQyl0KidS3HSTeAGwA/sCpZYZLl1zvzhEye4vGUyMxxYDeVFK9W6
SCiZr+9LpdLZK687LPJ40tzlb5g+wTnx/dym82mxiIZkQXMeuf/tD1kRUEe6/Is+
DiTPXjfDoRdyccb1pbLwDq9pFVKDc1u+2q8SwRp1MQWDnI5CNVugsPrOxdCYNiP9
RWyF5cmUk0IaGDKn1uxglQ==
`protect END_PROTECTED
