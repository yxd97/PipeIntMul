`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CF4e8qG7elED4yorh+fgDNmlMMkB8HYaciTaUk8BU4+MJF7QRKQzj7T8sH0vxjF+
0x3tyBGH57U9UQiKSR8nx6I5q+jcATHxtu4BWO9EgO1Rz8Ph0iPA2Wct3wMD6j7X
mTdvHVXJ4rXwZcFdwtI2VJf/mH1OXQhv6+JnluAdlKwMgGHBhep87QLQey3UQYHP
HooyzhY7rcQbIcw0k/l6/1GdfFTYFCeWnwCvXZym+Ou/merFokxJlzk/eVXkpQt/
okQdBUKH/SXj6pZ/mpgQ0uPv9D8ypgzGXGhdal7XCjPgg51V4Ox8qnRDDhL+w5Ks
PDGfbP8rT4JTlV+IZdzbHXHYcg5rsLmxOMEECA5TPc0ma6+Qxoo9iEz7zs2TFYtD
ev70svo+fOwi/WeAjGGvwAs7H9QIl9qtchXIfF7763DeoOrbI+jOd8LQrnr5XcEZ
n9Ri0fDbQZ5js+8TnyMY6D9bYBomDxVN8QRDVLZVEdg=
`protect END_PROTECTED
