`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vozDQ6YyH4zDgbZXHsUeRw+3yG5DGHsL3aBCyzdo+jnonhaiqGvJXnYP2SFyChJd
OHAQS5mTizUI4IPKKjzmYEkuat4B2Aj1GBI8aniwetO39VTA+HdpthjKHG9kSoJJ
8MskRP8h5qiZwMKKdLC8+fLfCvD3oAmE9qp8WP/M5xSXiuR1MqGmx04kwwz+eapW
x1MIS+eurAynauZ8KY/7ThtxNSz6nYKW4Wq/BS9CuvBH+p/pP7sm3FRP26JpnW29
Im5aXdgEgsKf2Q3XSYiJS4wvbbrw+YwixV1F82UMJoYf5I2osIis7iIjuyHOu5Fs
FMNCUYzx/O9BCcmOb4p/7XEiXj4gSNb7X/YBxwJgIoTh4crrKglsWMGGDv+k0KZG
8PZS+V8NqA3tqMwMepw37r3g+DP4KOwC69acq7IJSoZuzDIxf2njcB45OBHLZChH
sXB1hU73b9FI0sRSOQ/v9guzxaFXecpuxSZ/sQabiYbLchlFvk1ZvHXMKFEXYjjp
qOq9pSQww4Xg7jGOKOkBXf3BKQRGS+NGMEQ2WGA6TBJxht+CYkdUFbvKpXHgsiPX
T3InBa84aNv2mmYb4c1fBkec/FkUdxL+IK/RS7Ywla1DQeSbQseMQiNCrtKZISnp
8ragtemjjxAjKOGm2IZbbPkZ8ZFUmcujXYagTGR7yuk/tRhOY7OauGhZ4mh7meSV
2pfPlbuEEhuiV/CuGgBNgYwiaReECOd/pglUC+//AKcRnKjradsvDLR+LP0eIuyR
qrAbxNoiqiODj6M1SJ4dGw==
`protect END_PROTECTED
