`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lu6qv/1ubNQFQCqZXSv4XwT9itKhlMRI2Kw9MM0mAHBM1JbvTaMaZbeph3ZIWuxK
42vL0+q/MWzR+HFKnM1Fwa903BfaQ9zlaRXvgnK8hPB/gMOrPonH70T+jekzbrXD
nW5LE5a7hMNt1JtmQSSuQFwmY30Saj+1ZiIcUN1sJudXUqlLC4B3Mg4O+QyhsR8Q
6JKs9OYa/cC9o4tU2r8EXcX9KoEsHEvm+JLPTP1Yfu6imaCdX6DDbwqPEBo2LHjP
rrnLQKz2pTWRDTNw2y0NX2QQmb2PtDt3fhe+01/pRnI=
`protect END_PROTECTED
