`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTrs7fOU6Eql8NtecNpiRO9TzAQBLejfCRpfAkSo9hyMe1OU3Wg6PJHQH7z0DzVW
iyuYf8gB3y/0HMSldhd12d5AACbiv2b87bt744DVWnZea7qKl7C2NfIRNNurVhGI
/xSbYp9gBPkcDgQ7QOIyeoJYs2qoyDEjoQBHzeA/dnwVaceyrm4eAPjIy8kwz3TA
DxlGrZe/Ks8BW2S0R0awTtjVvEdlMUjEYQItn+jlYpEUhoVFxOvAXAzF5N8bhFyj
ydWJ7uiOFj5XUR3ctHG8pYymH4ZJO4NzGJo7gY1SSZaFWJgrXDOz5n3xGGpjpGDk
RbVst9NQhmiD98MK6VW2VhafOfBO+vNiBm6f98GCscDleoNP/PcuQY6kiJm+4GRP
HS3Z1p+pRv3aH8lgHrAf//H/HcxJqZl6j25KYYtT7YTuHRVTNlPy8SRYbH0fiLkJ
5b916/Qz2gsYAtlKWcjwQb+drb8lG/aHktl01FdAowV0TkYTOvF6/vWas9KUjj/x
GV1snqtHqSOad2nCydJElrSL+yltXoSVQ4bk/Cj7fD4lccs/QwqCRBlBmL3W9KCY
5hJkIcuJ0BWks83KvR6dGBPa3QsQoYN7GNB+DO7YP+0jYNkO9+CrivvRH66RzsXy
FBGzDeiwB1xH36eeJkJufgSYY73ejM6pVSvWHMHkt9EK+6llvS4IDGyHU3TFc87e
PpcRHpOJnehI/2QEJD6lEqRBlMYKOkiWZdcRAXx2i/JMmuvl2E8EnTgzucxRjbmX
yfoVnQZ7yP2tszarqIDzJIYMFnsYW0tde0o9QyC5dgl1//N9JiB3M7royKbpJ+4v
CF7C1+SdpZb11ORtwHVaZsJtsI6yPmy0/HgZA2t8vxLogPeEKD30g/6LmnVPylhw
ytGHLtLt2/o+9oSWvfubiddOJLz70aupcqXcq03VyTsz91c7QhVkKXEVw4ElB1dN
Lujt89EfP8zhvWK7k+C7qzntE+UGTf655+uMAiSYTF1t1EQqgcRoHQwK8SjJDSK9
Z1cJ1+37fWevVAbs1WPpLs1iwy1w3mNvuUHErHahEZzM4PuZyOXG7SNRsKUv+DRy
GZZ6FcHAIVhHR3ua4X9/yVViASf7VYEjxB1RA9PCnBQYHAOgI+k/qxVgpRSn+3n0
Nr/NTyA72hAIvaCHbBvbN3GfTrBtVe/QsmWwxcacF8I0IMXtyvti64OsPlc7hDQr
D4yzWU5eflwvd14ES8H11wNKj+RzumPJ8JO6ySgnOgJGnwLCiCH9zzLTSHRt8LpH
ZZtPYAsRSm5zIav09+d4WoJJqfctWiidYwqOQiGnNjvOpHg3PB5GVQSG8whd8ngV
RWCbDYaYCEQD9rN3he0x2Z5cPBA4u4rkL+RbxbcslJyTj6tpmpdQ0ZnGKLStU84g
`protect END_PROTECTED
