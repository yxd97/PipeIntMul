`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQ0hPRFQnU0Sbwp3OvZ6Q6AxdcvuXmdfiiFg8Rz2Oi8kMDX1muPsNBy8Mqdl148n
jPQvPlCckXorbet/05RibuOfI8gW95j3kEdX65tlZhlrTPdkcOM9F0roswMo7Ro+
pQmGybp0Ai92ujMmSj9H3bwpQ4pqzDO5zi7wvVXIwQzOF0b8ds2PPBuzdnMqeV+c
0sJWId3PLrbWd0szQUZ8jG6GEiEdTnxb8G/8iMnu6jopWNUhswC90Acdt0IqrnDg
IdVHjF8rEPcEGnm6/hl/sKJ2OaBhl231kKPZUEeumA5f/71r25+4qBTz1A5BcaIl
OYRYd1UqQV4/ek/LBOagCZYg8yr0uItEFt8TggPCOQNJU27smYJG7jKnNfp4SD5w
7ENiIIevLinbLMFi8GxO2F9pcWavBB/LPbw06HEfLDVpJLh4tGcF8HXsyNUzbpY+
yz+z8V93Ip4JJyfZF1COpNWBCxFoTy6XexbiV29+xY9D0wxtZl77rQ9xBZ4fdh+C
`protect END_PROTECTED
