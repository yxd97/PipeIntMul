`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jPmtXOzDMwBYHxsY1DrU2mSHgYZnXINlMlLywKn0dyEZmC/FRwIS9VO0QoNvaUop
zgE9A2RewNCiqk2AQFFUvCuUqfZ/Y2yYMLXeZtoXRCtKKv/r7DfsSSuXIu8gX7xm
a8exTqryz0Bl2ndfVB0dbtVYdf6IS7ztT7I85ImektwsliEitqVnGhTnaTtRrH/u
Gi5T4Nz3hnSSobp+qSQbKVS+S2l11pz8fK7Iaie9gMsbs9maXY5tHybUJR2bqpmG
IijVqcWolFAiyxFI7b5S5/3FflLFdq8He8ghqt5A7L8q4pSo+fDPfcddqcUf4TMb
KE5G/EgjkWlJZk0rvdJRhOj+IXmMyoJtR1fdZknCeQKzPqX0mmE2p79M5yaNYgKw
pt/Ly62W22f70O5YkT4NAgvuP5E3OAWmUmdlPTgrxYU=
`protect END_PROTECTED
