`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vVc9eI5MkhZ+xI55xTYBrnWWbhfpD4sh4q2ZO4ggmFznUr/xsB74OEepUSc6oYDr
BJqnUr6mrdbvE8Brhk6MrUOJgOl1jEWbK/FabrW3pBR06WwHOKBmxkaI917gBa5p
Q8ccxd4gzPMhcinQUAmj9SbusMiKdaMDfAddTq4AGwB0vmRZQe3ZPJEvCuBq4jWJ
Aep7sR7FJutQPcjL3xkITseduCVJPAe3UiWyfd3A1R/UMa67nL2cl4XV7fEKZnED
WbXT9Y7vMjaOSxvqcaEYeznOPZKTMXS4ElgCBGRYkp3nKFlrjldV4ql7GlQNHvZT
2vH47hHK0ItRCGpZTODhZQ==
`protect END_PROTECTED
