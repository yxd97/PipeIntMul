`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAhmu5zJ1qrxzdX0NqWRS0glKtjSqxKFG6vCf5kDvyYF0ETMymgtpl2UWu5TV0hX
CgFcRzAZCQgKPNkm4nrglxNXYdG5c8CQ55Jbcm9Or2qDL9OgO6F+0p6Z4xdiR+oo
duYStG2FlA9Le4wZZ90OtUkLcrz/59A6oYQh5gT/wbGcCg6eGyflQvtHFl4ETkPU
Cdn3+zjOJ06kg4TGIHB3rBuGdJq8LM03HCjePlN+0OQaiqrIM8iUtaJH+IgrjD1K
/hNYg1racywDIKWXk2nJHUq7MPCJ+OqKHvJRfYRomA4itXMI5VUDyytOXIj+wjbe
`protect END_PROTECTED
