`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vWInKd4KXq/62oR45XYSd/UdbvjyaJAFe7NMp+lhvgjaU4R0u2S1pmO4BN+g2na
jhyohsNNHvocMEEcOlVoxqfqlgmDJX09Fcud1WSOnKTvGZU+VcEqSbA6blC6oU4p
98oxr36okEMXAu8IleWUsTtiBJyhl3Ub/tjudvde6KfNxxcX0psNwNJd9OrwKpXR
awNoFZbUVkGnTzDO+OYRgJNKeHkTEXGmf/FvNSWTHon37G7LsPEaDcieXpn+y4Pk
nCRrDqowzyPdNvcnjj1M+T3aUTHulisbzhjbdi/R8lSabJ+tMlqss3LXYPlua6Ho
xNoK7KHs16TFX14wX8Zc5gLasOxvWuiS1X7pKm5GV0zYduoBNEt532n+kSew1mHQ
tEMyS3rW1vJkejAAPYGRSJjwwJe8QeMBfaM6RW8sziTikRMBJvzh7flsVspvTcWI
M/KxFTti8z4SQYwlEVFlZG2237JpcdFQOzAkYiwDaGiPwqn5BB/CAYOojXFAnH2Z
lRkCzxz50mfp5Cw8HgMN+SagAvFWPXGyR10F+IPbaJBzMfh18e8r2PZdof2UwJ0a
+aEv6kDmJ13TM+8cibMJJaA3MqZ9Ge16Ediz/MzZxWSLVkycQMM+sD9TPnEYejNB
/7U/diEsomviw1YSo2j3f2ThZMPo2GtMNdY166OXm740dYGkbtwicEcqiT5I3ddx
P22oFzxEHRCrM5fMllMuhR4QVoNLjd1V7oXuZaTiMwfw5DiNTAYpJN1lc/8vhmRT
DoMrHG3Gse6eERH623PfxnvUW0Bqs4xbShP7CPFI2XCBvxpxWz/VXo5X+YWX9PiL
PibwNm45She4R8tBqeCO2osWuemUJUm7W1H7hE5Pj3JHrkjOdb06TtaO+Arg2PtK
sbjkuEGXJW6hreNXzxJmJG8Y7OZANGlHfvcsnpK8nVREc+bf5A0kh0Lmtknz4P/q
lEg7c21tzrIrNLoT4ybJAg==
`protect END_PROTECTED
