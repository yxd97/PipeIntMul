`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SIuDsyDOOER5e8ZK4RDTyGPXFi0NSSaVTm5MOG1wuMuDmJNkDyVVxRBLSygatL6t
tpVwTW0BtOLts/29RmBmwT7JidgA13fsEXesmU3mgY2NBRTVczzlzljG8BAmcWkC
Vl6Kb4Fu06tlQd5qg8cCR/jvUHgJ4QsYq5Svgmbp+ZTQ0zKdF5aX42BTmVn1lg31
xxDwA87AMUOEGnWFK6N3APdUz5+x3bCq1VTfglLNaoXWmgu/oOgDDd4f76fHzN7h
rx5uUL1fnGObxEPxbI2/mwB4ryAA8UjPonKzXDh5q6bO4A1iI8J24ExEvUVfvNGs
THOFA+TfLDCHjd57Yd6J00t1b4ctkAWvbRuw3OqW6PCcP8tpX7qRg5qQS9wcWSrc
teLOs4xLco0tCf3XsaIyD14qbO/yJYiDMfXCgfZO+XFVJAbyerpKLUW4PUp2NVw1
`protect END_PROTECTED
