`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8+bDx/cDffiX2vC6s77VQiG3LW/sFGUEh+oCD4ASEDZFk7bHo192iHmr1OVz68S
2BclgD0a0O+i533QnLwmgstwnX+CtokPqOPP7RAwtqGlSMUntw6+9wWD1p4YEw/I
62DJJHsKaDX5X1DoLzAuf6pHQHBRAlpEaPJppiYSCOrgKnFISKx4TW5wN1+vDO2O
UOFsGF/0nnSRvA2vLBda/ao4MX5HJJafa8egfq9249+1q+Gm8v6cUts3EbKSP7Pr
wKVtouxNigtSRjtakorGgLamLQ4cD0bMoiYHAr2YSjNVCX87TfFofGjmUjugyDaC
5f0V2B2Br8hztq+FSDXCZlGwejRCF3nohvALajg77gNwWR+rqw0IFRYUdov2xcWR
i4cMbojObBWVxZEohSt6nhR0b+02wZyLLLZlyxnxJpQT/VTCE9v3ozjiBrYJeHhl
lhF/QWq7WxJ/FkByh+4p0X2vh52f6UHxNNB83F/9co14UmJp04VRa8Sinr510FfH
dsKKnSW7NPFInoWaIoSeAtrBCWMAXRGWuJp+yBtIazVOIRVyfvuKQKuEVxZqpMMZ
pj6oIBC9kd25ItnDHr10PzSuaH8ykf82tf9y6ThrfHD+H0nA+Q+etnWzuFnr8itU
5CdI3iNm8UDsiQGdFYhggA==
`protect END_PROTECTED
