`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wWiDQHGkzQ3+zODWh1yjA1uBG+PM0McN3TiJoBVdhvVE9FMoYyRjPVH7sgAijirH
LOoG4vsrBCTxp5F4pLdc12dSfEVrdHuetUTA2liIZQGsFqVnd8/0YSD/IBhEDXKP
KqrOnqeuZyyKgduFY4fYwSYtusTJzh+2AxMhMXUH5ZhMqYCSAmp8aV4GAmz20e3G
qO/q7uDI2AfpkheCAEphGnED97fXIwtvNNhvuHAOHq+jMfuEjct1hIwhWtXqezeh
TG6nPQ92c3F3PgmJ72G4R5wgz+6atyM0dSD2moqWCl9RqLWULsxQYzi2BsJThOSI
VQJEL2a4bSndqHS91QIDZFy0rz6zz8vwy3zBwSUXmCLobc/RH5YcJPcP2YCOf3Fc
yr0M4wn5twtY2VTbn+dhS/T2hF8KqsIJ7p4+gPe5hT04pmZ+8XDmhlPoklCxIBlf
OTMu44N+epv32QwBaMREceZSdF/fhWl4ldAh4Yaeib3bcfJ6tKkLZPO2PBxi0PF0
aI2q64X2QEUs6n51cCD3M5g8ZzJC/l6tF75GpJDgAz0=
`protect END_PROTECTED
