`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
et3zR5WGlFYKPABCte6mRXTDj4VADFrzJHKxjrZEjZlqI7j8RzCrBu7Nn1K86zAh
mVEj0xIB0m3NcRJAqQ/9gKiWf+u+RD2LF+tdmN7KptpGPdiam96aqlzHCqrJ7w5q
VQWQy80/ETR06ZcNnMqUg7JEX72urXP36E1o5yuKsbecoThxNA2fZTCjRwMFyNvk
BF20TRrRbqEBSxfervT52sY8VpTBzxprccUjINb4fiMJ+e1uY1zJeFmpWLSeY6li
OvdIu+CTUxAWR7tDaJl5x4hmqPFhNGIt+O85ZEq7h7L1pC2rA6PcjoyCNYIwiqut
GaumggrQZxDD4S0V852bYXk8Wf8mP8GPIHcJBfQtkg63WSpe08rfPI2Mop3e9+FM
J6FC2Bs6a6E4fJiKFHQ/6r5xl+RV2d4PJW5SoJBUfSs8KYDfFi1uxihW32pfjTPa
TNybGWfLsT6GEdKxjaZ+UdcReCpZ+Gyh2l5K9GkmjceUq2pgexq6/Y9rVJplsoTn
aiubJHO/nXgwnuMyR4j1ZrydpLgaZnFw/+oOuGTAmOlwwqPSDHudgGvpTfnHL1AE
`protect END_PROTECTED
