`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ADtLIdXTORYWiOrwrRwBLqqhvzSHSybFzDhmOXoZy6v6zbI9oTVeOk0WRdpQInJ
6uxi+wJ/UnPpcLw2bLtTrrRbpzX9bcVPpCmD/gjfl0rrnKeY6doe5P3bUhxi8eFh
XN/I8UOjGCppb9smCLFe5pZSC+CQtwLxhKFvSH4nLXApnrrNqq5Ye6UQ2+nGvDR3
+FG2BbwRDeuJSaLWGwYWDSrLs/BSd02tx908WHNnBLCwK7ZDBExVL94j8cLF/2YV
HvTBhvIJkXjWB9ZskM0+aFyKnFDSe0qqLjB5bpR3vxAV17vEip2tmqAGvk3MPc9J
0yj90hpNW0x0S4qbUzmZFnqTKN7obZK1ODxYD+1gqW3hf092Sc/2I95AjESW3NRw
cEcGWcl6Z4dXvRLyHE3o3V/qz1FrPRgfTMydxNRC/p3/UpZ6zif9DmrCYBjBq6JN
w8N6fGdp0NiNP+eKUjK+JU0cJe5x2UblyJUoBzlyWXxpnVNfzr7jXAJVVVvOELwc
PEXebDdzvzU/Gg1oiVnjn5KRlivIDbfBeh12YIShLhamo59mF5lW4rpTFMUIXqS4
7NmRB16hqLUABwfNFMFd+P67vXFKcuzm1bVXSV7mkgKLNGYG5pr1MVvG23qOkuLJ
7IV9+VX74MJGTRArI5PUomKDPlEuX6gVGQaAetswRFrr4ZwCVZxQZu+H2t7R3Zz8
ZrNCNKLy59K8YfLCqUN4GMTGF7c7p7+RrhDcKvI3/xjCH5tQnoy1J0JzBRm66iwx
`protect END_PROTECTED
