`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
esOwncJiZyFWbMd7Mkhoskt3MfE6cmHul4Oisoe1kaFGuOxZ4o3Ihac3eTHRqLhQ
X/QQG7NULy1j3j+rb4bBwwE8pO9rG9QcF2incybVZSpOVULWUrmtcjBz+ptPiLFN
j/7GBtIZNc8wwe0Y6iftEAeok5czh+LPAlokdvwjyDeTuvygyRuFBHqTmtBAv9EM
ki44ZRSH10R8lIfl5osYyZDybc9njq9vcaBl5/ysQ4SAklnXpwZ8YyXct5Pvt1Hh
NMIezFIbR0CWZQbXB14Art5OJ0AaBqo6MeWq+WxzTUltH5gJHc0aPmb3Wlvi+8eO
btHiDp95oij/pkVYhstzWg==
`protect END_PROTECTED
