`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VqZn0oZ0L2MsfYBVH4Sok63g169bGWlqvXTcjP8eCYtAHZo1HSarVy18+79h0B0l
2LLqEQenSVY2vbmVRmECaieafHhO3Dr77HF9XE9odIckvG29TLCX7UcCcBfk0ZtB
FSVjEVXeLnihgkniW5VZeyPPPhpMrAferkd+Z2h0H7tl4X0QE5/NgOda3XUYLR4m
V/7tBioHmFBbuF228ArMDU4sZlulLm4ZqUK8dnd1bXmAqNbauNVViscMWg3jYNxg
LgmR6dUc9PQfFH2kUggeSiBljgL32c38njFKYbc/VngFb5Npxxdpl0YkkcfrgGvm
+x+TV6eBpGd6N+Y9t2rU3pxMytxKFjBe+B2wyfp19L6KHoAC5FuYJI7f7Q0ph+QS
aa15gEkUQCLvS5VvYPawf2HscdE96CQ4/uN+eWQc3gJKEX79ox6OYi/97P7w/RuY
/X2l39LRhC2GV9dxdL6M9V5Bo6ybvSVeD71qfAYML5wtdRkc1FHIAjGf5YG9j7DO
1pC7l7R1tCAna9sNCiGBUgbWIUXtpoye8RWPrvYCHXdBzFJjOhdxa6hl6+wXLV/C
x4uxt5yLdTvFNd4Xeu0tJf/TYbiJ6xDSwfJ5hM+Fw3P117tATjZHYIY8gUw8pX2D
qko2YYNQoyyM3Arho9RwCoP6BQRq/U7U8sLLz0FdlstN9XnMvSYDcOCayt68Oy9S
GF+aV1fhtzhLsGvMJftEOhJRsBrh9TmzZxremyg6G7fdD91ckIjkWA3MXSpg9oJq
kZIRurHA0oWvg+zpf5WIQvTd6pwgInOm0ClP/6+u3NRfCbey21tflFaTzREWQArZ
FmhRThwKRl5Fie1SFoYpPUYDL85lNWtSwLr/rPYz4OqyBODJdRGY8Y/jbYCpeH6y
s7sCrVsn/m38R5CoKFUMDN0c3sC5nj6KaT6ykk8HcrqIIyIZ0bdvBuDSkrn4rFUH
`protect END_PROTECTED
