`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C0jyH5zIzId44xUQjjp9lm6QaaEd92oNrxzey8gNk951sbmGs82dgKvfmfqtH5Ha
tHmwcZgEKvy2qdH24FQmUyWuhC6/pFnc97TPfiNK5qC7hNrjUBX9B4cDiiGYME1N
bOK33T4LZzSmZIskWsmg0a5/BG1dkWcPHLyh+ntA8IufnZpkNheXIvWMbVww0iAQ
+wakr9sauAwEy47tVLrGDy0LkDdl7rCe76pU3AqkpZrZOZANUv6Kr9OFBK7b+6HF
OtdhGjNmr/t+Q5KFEUAcMj+ZvF4IH5oTNxKk4eQ0uxA5bKbbkgUdvGSH/aprR113
u4Q+Zaz/jbALlUMpTJhMbjrqutAf39wHg6HNvO2vB/6+ZQX+oyfcbVawRlfw6hSc
o/EDQgWP870vVf7eKB2K5HznCCD+YRI/mqkvaLPv2EABrRIfR1XTMq/PojDmtHig
3ZHfIpHAM1rSBdRLZzvgtb/1i6dpwImsuwwTe/vvTTISzq7af6AHAsM8uZ/H72YY
YiBt/1rmxESRuzvrkuJ2W+ywwSD5GLQaaGr7TiNAHMXajdM9ogC2TAGRiiB/KOBS
H/lIgCDLSRGDx+XvgBhpDddS+jJ/4MpVHv1oufdimZf1HkNV2EJPXUgwj24ftJED
yZQ7FfkIt7/Q677rwy0eVA==
`protect END_PROTECTED
