`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4tkLbmBTHl/cE+uC6cn9vnagSXITQA/LwMzc8bbScUoyfCbmpZzCfAFzX57+sKHw
fDKq+19lll9+a9fuU8yhVRbtSKd0WkL8rtA3XeGakle68645Am8WSq7WtgVSxz76
qBXBpbkHl2d+YiMr2hNz0Z5zJCqsgZPWPS9rmUStQkdYxGJ2niiCZ6BCO2Y7fuLN
iz+ghHjPINyg96x8ko9kkxyq2NL1kmPr4Jg2G1b8CHmRqYCcIHorNuwGgl6S10LO
oPITRY0x/YxPV+jWA0NINPamX2Rkx0hTgbUN5rfy3p/W5NTDyCd28IOiZvDPv2v6
QEfQkIjxuls8BWkXTnL3Xb8OdG0PkgtfHL9VjqIoYoP67hFihPGjIO5FHe5dvosc
woWNBnKbB5epO68Hj1ufPua9oQUPJJVuYA730IOWrJl4ub/XUbWp0a822B6C5Rma
S9K6nxyL1PJl3m1vlIzKq9HJV30l3SiuHvJ3YXPKqGgcNwPDT3XyIh0q/5If2SP3
CZoPPurZF2Re5HCSPCVCSv+QSni8eINNLdjMeV89ew73m1dF/g3Z3AyUMkiOiE/L
eaPoeQCEVOUoZt/vJanH2qpPICoyBpjmzYetWaRZ7TStlP2qrTdNsdJlXmJ0IBID
RSgxz1nTt7HrnfpFeDrlpeRqDxezyQgFjdZgdRyDFX09FOc077kgr6In84fYTJjy
aczk10EE2H+RPnkEF6uhFWZFf8sHRHiOA+9oaKJIY6h6axNWZ3Qa6jKviwH0MRzb
ghmvMK2bRtKev7atmnQRc5M18I2kI2UGjGdEK4GlltnZXoOOus5Ttgv5wlQs7yot
IEKBOaYehQSOn2nAhVi8Uqrbc8vLU2dDOqNz3gUfkmeZiZ+pJbVvZDagwjdzVqVB
maSlRzkFGcIsIvUPnOrwq0Nxj/rbnU91egye0+cX80SB1ybGkC5b+n5uB0R5IcUR
i6+ILFTozkjJ+06RSfDplQ==
`protect END_PROTECTED
