`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xsaQujR3bIYOEFFF4TysMTTdTzNnzQ43dBctgY3MgpPtYaVpExEnAWo8jx7aH7X6
Ve/5V34brAx1hwgH3A52iNNCIwpemAOteMwKlga0Rha2LP24bzzANJgAE977v9rz
3B5Mgrs4/rWIyu6+dU01d8wF/53VKA4rqw9S3ZrTsR3MQRlZhoP5sWASahV2ovqt
hMnNJxSGD9MSAnEar49csI5xxN5mfAo7iY7QhR6esRKXXzDVC6OyuYTLcxiLhCAE
e/Oami3XA6Z/00x3fc+KacTptujLbc8N0+cntH95y5IbRMVB4hSZs7rwlQw/QjIn
qi8XscZX9p7Ry+tqA+8Nv7liWlavltLEh6ubA9wLT/tSgFT2iNMC51zq6QuSFh1o
tTlO8RNsbj6RwMS/WuZi1Ds/4xb3CNuDswihIa1pv3ImIgmz19W/JogQv+M/Jzni
BS35Rx9RqegBQ3XPkeB/z3npTPRGQEfTG6KNsEj93ImSUS4gs8CH+YkWamvA0O0k
S0M2gUPEGpR/kHi7fGafRZDlJhQrBJrwTCbZyJuu8Ks35ljjloD3ft+MmF7CohKN
EBAsyWa70NnY6WoOYctr4uZHweKL80Z5kW96AttqA7nprSzoPVAO6P7lPj7Tif+k
eQ3iFgDVq72ZuYLc/4lDHw==
`protect END_PROTECTED
