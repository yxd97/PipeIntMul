`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+7xjx5tAy0vG5924pceS68+R1o79Z+ueLvX63WoLl9Yeg8GaWcds6FmgoBBjSFv
fDvY/wjAMgOAVQE0lDElus4bYpRQZWBwzgJ+MrlIUktvBaQ/maUXmfnXgZB1k89I
V/HF4AfHed6T+147Z45hRpzRqk2dc0+FqLAOTTUuJDewguxVyeoxAl3E71xRX+YL
xGkwryO4qzZnZ8/gJdE3/PI+iN3hE18CDV46hy+alX5FZnvPRZeRoUaQjJqazmyw
dkB75dYnEZGyBMau/PNmOuk8JT6pfOH8/Zs75+mKqJyJ90PlOtx1xerJ0pvikfck
qZ0q6o8yPpKocS21ZIwdKF6UZGnhxRl0PNyj5leVjzGRvQhTZW8hdJ7yS3oFHz4A
rZwyi4UWxD1e+BxwES3nON+xPTF/LsuGiN7b4V6drcsboIiaXJYxUlxY1+oOymQo
TevsTLKhNAuC7dO9ydI4qsrs+yqtipzXlRWZHFCVSrPbNuJJgIwqIhSktYQqN6Bq
r92ZyCzt2MJJ9647f/8dRysYEzG5QRKYv/142bBV1BFE8fTTPRNTbrNxFeQ+hzQi
0S7bU3PziUqvibtiHQxHBEFOhA7Voq2K93fXs+VAcSLrb4osnXynmi2k8xPNCoAp
gWU6yoGwLnrZfi6c7OqXqQ==
`protect END_PROTECTED
