`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7hcYYlVV1e+NfhApuZx4KO5qRyxOnUoi7PYDEJRFY7U50UYJqpKgt3Qk/6R+mtTO
BbqiIXYJBSnDM5QY1ARTvc0GjHnAWnqnYISF6aNy8PaeySqnXVUThaaso/sobnJA
TwOuUVGqoZyVkmaQL2cg0P9rQ0Ue06hvwseuCPlb33VRfzKNEyWz37Tg0E2jT7ts
y4A9DLW4AjdiR82V2bg45e0gdy5p27DNUyXncYSeiGvQz8N40ibWgi6jw4+L96dr
43rmJKU/ZVTKyWwxJ7hNFzKE4YvEqW+f3g5VVtS0uDcgutTuLZvYe3rjODBCXZbu
F868wMkHtt9t9jCD//f4dA==
`protect END_PROTECTED
