`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OOc8HYCnBO0YOKBVwFlzvP2cLjhhAboQSGAUlrbVVfTltay7UFpN7PQIc1zFb0es
PCmhbi2z4r30S7LAEDAra5QjmyqkXHFNpetCDi1yN2cJdvbMpFSLQZ1z0OB61vm8
FsCnpBzicdcQzg1zCL7ZtvGFxj8uFyK+EAsoaqqIPnGhqgeDGKgL9rXYZmcQBYp/
GR0NeRC8KVPEq9G35RrMIDVb92hgmqYirTvNxotzLTN0AhzgbALPqacfo8Q5fR8+
AXdsXvzwiH94uwe7v+NiOJOeau+GO1GoaBjAkPKFcOcAWnUy9PoZy2qDwROK4B5l
XfXzEbS3XcKs1kZvfpXyjXqbdQrUptTfyCSpm95viEY=
`protect END_PROTECTED
