`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SRSqx42/GkYkmuqHj2lcvFZ2a/Jml8sePuBdkyQ24FwsjkDdnOmBWNAlvfdGARtJ
NUigW4/qH6MjnVddDmNfg37BkCwQXMAS01Y9zIFBSniPktQZnFMSo67gBIoRLJtt
Q3pP9YJsIpr/58CCmRvI1hum4kdHRxxOgan8R+hNqsA6/ZVNQi8ri/P5oglm9rn5
KQYvVXTROgiO3NDHeIlJqr03eXs7+pXmQ9VcbMHnJoqvSvBMwaD9xkPqxVci202j
uFlqdtH6bCDPlY4yYC2aZtG9tHrgnU0/oBYLo7w6UCpeAwdHWza4aisUDtfo5SX+
uXDzJuMgXKIKDDGMywrevHC+cfEMwylsN7Gux1sf00B2TbdwCJmLxBQnlAV+E9Nz
`protect END_PROTECTED
