`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mh5KXRpapCmgTDTbNN1yPIsNWBDvqVj8JqFP1I1Fc7Xi+0h+LMuICYCXzJYYtxgA
j0vb60X61ak/g0cf6XHhm+9KHioq/xxX8vx+2wkJ79IL+B+VXp3UkklMj10XYLbI
xV5H6quhtWVe/bG3UR+qt8nk+PM7jSWLFcin5HW+eACkF/2gDlIgOwxO76xt3Ln4
9K89+OR/ln7sg8E1qEhb3OV7jN8A/QdAEoV6spO0DqYjzFL0FboBQOJdI+zpO63x
X3BkiAXllaG2jUrDl9Kkf524lMrmcsCzkdyjZGby4PL86VU9sXZjR3jOyhvYBwKL
kdBLPFWeFxBYVyu5TWic88sSwhN1xhvRBPo3ayOIHZoSxmX1Kdq6CNbIPW2PCQyC
yf4G0UxpKp95GVcIEmk5rNZ0FZ1uttPxCjmREXWhkdlqYSxAYiEEGJLoJdHG3vH4
10L8X3yEPGOlu6Cw0+4nswPLaA0PkXP/ACpa81aNQzhTkLfOGGk/xC3qIyNTW2kQ
`protect END_PROTECTED
