`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1Coqs9nBevsbmIANGJY6aiWeHVIC+yTZk0ySfQ2CXudSTdFLhm0K5vkawCCRWi1
4nJpmohXJ3BsfWcCsIgybTu2UM1vuGU4fjC/kK8TgFXkwjGc1CTJgXvDay5/zEi/
wWIy2AB3mdjr0nxGzl0rTPp88GAiYm4kRfvAHoEtApPN+lSWIJJqgkJyDRGqBh+d
fOH4gUg0f3rweJEjz0C8p6r+eQrTHGpIyxRVZsjkNad7An739NTPtRYIR4A0k/Hz
lC2xg9M0f0EKNIxB2i6fx6xhbfpH7q2wd8aWV9NxxhiZMefpZq/YpgkSan5xiMqv
`protect END_PROTECTED
