`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vr4XrXXFYCkBgnXgJ2J+M+0xGtwScp8f9fi89te0NnudTwtSxpfQhvGw1f+ZZzys
MEpYnYk89FJvDOKkEUg8+v7aOIRPBx0Fg2IpGTX7YhneVR3PRQOQWDJUkLgZMFa0
02dS3b4tymsm0ueSUuJ///wVLJv9p3ZxSdHS89YJt0/EpZGYk+PkkU8ZRtqtUbva
OjW+JWvvK054CoLt8ELY+N7hbYett741C/E2RaXohVAIEs/jKRLG2eJY35XhiHJ1
50bNmyNLU82SyQQ7Zjr6uDdCOGuAjKiGuw37kniNto3lLbEjHZP7XnY6Y1XfTGrG
/EgQytBA5hAzJn8rr0Y2NJX13IFtQNjLLf2MhH0R7d/zCYlXOOW3xDCNcW0aKpfu
dXg7SRJWKnA7qFE1znfLbV7xnXveUY753FuESCy3xJqsp/YDV58lnZVJLg7fZDfR
xg2OhMtLWPDLHfsk4gi23tmvNcF1unn2ybw4669apkVfOU35ZOPCRuf7vmPnzoRn
C7kyUfCKNYJ7kWor70WizrwwFJ7zK8dR5tsXaCx6jnIL7z3TeITD5yLYRH5C/zwo
kRn4W6YlO3cS6wiunpICygbGiyVsHbmYdXb4Gu1lqzJ2VATLRIGqOaJl/bciEv10
B/hsc07QZb+hDPMSPV37BKmF9nqkIYpahoeG802QbV2JSimGB0KyACsidu/vC/cA
aKY2ti9BrCpc94NC4AH1dhFIqy+O/Gfs6hu0ngpjo+BriqGrk6PSUyOqnEvafMxw
SDidXHTK7jb7wZ6jcIq4uRaAfDRO+u+Proqy+pZ1vJ9x9saXlQ7eROtVQKhtVU9k
iYxHq2pYdoMZyUWGgvd6tDhJr/BLdVSEdmcpt77XgiF52o/rirCBfqfwuJF+BQzL
1PyeUeom3SRpN4FC4Ywf+dlkFMS6dQZNCL4hZs7I+5uUqdN7fiS1/1uz4myxVapE
GdlKsbQfwnXr6akqWrNPvajb+WRZHSEmeUnsk9d6ORD4a+vuT5g9der7ezNu+jhP
vXx+a3HnxmzRarskdZyLTZKZaH9B0uWC562rSxFmHPK2nY3LIVleA4i37AcQnu3T
QAGthYeJ7lQw+779y7mjbRC4iUsiDWyygbtdOY3C5LHB5hFGFx8s2/iMiUn0wMZg
ck2rAO6CgZ2GUxKJ9RiL14AVS66W5h8Vvc1KZCTzrXdRQn9N7/iHNf0U/1hbpih7
Ks5IRpEYzBX4WNg8S6xILjX+xzUjtrVFcMHMUFlnGvSst+UoMQyH+Iegc1lEfE+b
0YjtxL4T9K/pWXXev4M8I6u9BxLYuSzYPXUIefYjgSE7pD1kvYA5HgVU9wvFneyB
aI8quPd0WJQnaJJZIZTzFBtkHE0FUkfzW/iMWSZPlYeq9BpZKLnHlgWQSki2qxG9
D9wy3KLo9KpoAqyG7xuywDYyGJB6aGhbhM0Wv/18ssYLFGoa+koDN7L3ZGymTM8B
dAkBBE0X0FqghIMHHY0EnoH5tY5mCfraQTbFOh5s/EfOGI5HwhJjStMPZtOLQJNY
4QiwK+GaWzmUMhAIi7l6N1f1XdreakiKtwYW96A6jyKqUP+p+R53L537tRYVYr2h
5WafoUHfBUn6K/XXTITdou6Mih+VIKK0AysjuxIubcrT8fAipwCTJAgN26o5nhPY
Hb80OTsC+dJqonDT4DyPvKuw3hCirSc/yb6+6+QO+XdefOnjzVJ/N7vocel7vnmG
qlMpczHss7okVLozoFpEtF74QzhJcsWCZybNgYqyPl4CFfe2GDCoxBVkB7jfgcWC
fMdbsZ31uTXRrg/hge1I0cCBa9kbKdEpy6Ptrv5tAPvkfYLc0bWiOwlqzf3G7GIW
rqk2ZfS8ziX+lqBzKi+Fv6HHzita+5Kfi88lIr4jpIsEhXFPJ4z0EBuN7NTgkP49
VVyb+s4YY8o/g0bWzRl9xssUDqFdqhm1ud+Zj2knDcUW0b3Rv3ubo9h5YjyFlCYm
IV+AUgqxhEijT7ORzZRm/KIdJBH71DJzJ4/8dsnRp/33Zi4ncALNXSuht+N5cIS7
7sb8O+ebWQkjQ7EohW2WRAGItDhu6tvhxn8O1VBfzO844ZBWnS8h46Iv1loXnRt/
8abFh3u4RozjvyVbrYB3yzy8Tb1qO8Yohb1+OPKxz0a6RHA/cP7B5SV9ergE9ywx
uacN4XYkMDEjkgWmscoiDYBzQ/qzkADECJN3SgcvUuM22LWTyoo0XYy+A4hz8MK7
hyBirqhPSz5881Lou1kUCmnJCqCQHCPoK7egj2UQqIVZz9/9VZNQMR55hiWaM0yd
XXHTC8CCEbMzajOEN2xmBSl9HY7J8FpNwsPkHLhOSnjZILj1mDHldqdJU3Q2vcVz
7KG4ORX7udBp60hRue9/GlbgYYAn7bgloIxs3UYF2fm8lD9OcokxSxlcjG3826eW
jzK6i8RYIffg6gwevIfbmJ3Kvf2qAX0NW3ek9UIhV3PuqwcsEXygKxTdUSCteEut
GvHm8ug0VOAGG1jrfUpjr4dY02P1bAWvheTKkem9Zbk02IPxoeLZrJXfQ+Bom4ho
lxP6DUXfxfq0B4/g24xr4AhETcgigSkRJUC/rD4W7G5RkaBF+g+T2GYMqfW82WjP
vL91W/p6DZlvYieTzyyETprl+R6lrx2c78yc49yddlvnRcyPfDGiACR4tjDWHaxY
vpC1vBXFs8IvLx+Ob+5CTA//uo0+psFevIQd3sL1u97y1U3gwQmkHFEpAiNMJzQf
9DlCb7uaK6YoN9YESq6Ds/OimU6YQ6G48m/5zhzVn2V91V3x3xmxx8v+pCisv4ic
l4zXuNWM1+4ymkVKCdBHb8/WXPCC4xT3e44vPLfnXK3Envq0TWK0uj5NbMCrrMkM
f1cHyEYayyB9xYIZrQ9N31JEW1OajlOAYxs1+GHGmRqfUpHcHki8z551Aq7cgGpA
+odw7Y/NxsdqBDvhVLxmT8dbb9qPTHIZlL5K3ZYaclV+6lrY/H6nWBybq5rMnSVW
VJMdXaB96C/S/3ih/WTlGGDhwaN4U0lwWuFqRlF1PAuEaqQRMuD+2ZYT1yrImGaH
4jgr6duuPqxjLmPIAxnd8Zh55Wp/dYfd6bYsNoOzulkB42yr0+R7ipTWuDLUdvo/
QBUXz4QgZCC129RF22p/QcNywvGI1viAykhhfergLytlbMEUOj8n5C/d61DpsaMk
+dnhTxBWthSihqP5WTcPV6XTcemovapB7CEs+hmQUj9ZoD3TcVPQunf4HZKwmTYh
zeJ9pPLiPurLByxy3OHz8opSOtcEM1ztLr+vNLxIws6R7uwsphsXguzsP33/zykb
K8c+stjqEKT3KMiApZqSyu/2IvqRI5EfLeqJYKQz+HpnGUEmxGrzR7EjnRZu15/R
ci65GkskIVwnZBLBLPSy03FZFn2tFHx2YX4T8TihPtPpAj4u5oP78E0w4YxbBZwj
UPLSi/EQA9jqUKrB366AJIyPH2Efl25PETq3hrH5uqjoo9C4ZuP+PVCRklhMvogf
PYjuJOHtv99kLIqsZcW2SbWK5l1/nv++CYNacJyv5G8su0RUaaeCam5Zz5TwVXeH
T9ZvoeoAIr58SEYamMKVLSUNr/2deQ4zjONk3yVXNkyXyg2yQiZ6CuD38OgKrAAf
LTeZbTXNnLqj6R1yzwUOyfjDkZ7dqknf4qOdYGrQ8nF4MaZHmZ/9kHls6cLU/vCI
YGRnEAtvK9lmWGxOJu7ru1YrsYJCMR6MAreab0TmPLsO/BN1QEFQu9KbhI8XFgS2
Geu8DntWAEQmLDO1WeQ2hLk/B9/iS9jOPrc5+OEf701bsQS+6UsvSaHe3mEquXEX
o2pmciT7gvlo2upKe6k69IJ+Wx22x1LjcwYqz5WwAfWnzbCofbOYDt5+zm8HOQmo
wKQOTbYwZTWQq/aN8R/36bCPQK+6c5aOFlx7YGXX5sfhD/rsKTXyzSSYTeGpwPCo
GNZWYtSYBSBb5ZriEYgjPoxq8ituntLKvZ2+zuzSKVKUaibVaWxjcPkfH6rWF6bp
HrLzqaOA42YxcM4GXi/9YSx8vVA4e58ASezqWqx+oUnd32pGv0TEIwYH/IcwDlTU
UUGu7xmay0jtifFKGuBEds0Gr0EkQe/9LQoHNszg9GePnZlTufKkrGA33OPH8jpo
JlKyXvBETcFqerfjecTBlZWwg8UiI9tBrTsxWQBNDQNixB2uwIaJ8AvW1ebR5L4d
sHMfsFSiLn7r7/mmjKdJgEnkPc1npyDwBQI0UibbRBQVjw8HzHmRl4tW2ROkgAT4
4vwOjFfg5X67dtg+I74v2LtO0CpqIP8I0/JvszX2w0ZYvjZQ5LKL4ytOMkkodTUu
m7CFL2VI/kFH+eGoyGhkqu+a8EmEJJjFhzY7LJVyCjM5jBBOyFt5nTc3RlXbMWBr
JTEAVqDuNFSSHn3MbgtWVKrPq8c8/71mhtf1PxMrhIC1EeqmKD16sXIzozSWVdtk
+/grKGaetJDUA4+VrTrk9wBoBJ+1z2i0A3+0gEH1EHGJs6I48AL2DmjRBW9WorwI
ResLTDC9wvsAWYEcP6mfHZ7kIQLsbyXEyiJ/UbFrMu02Qb6/qcSoJzvf19ynt9hu
r3aahiijOTI+OkW1st2lwewhSxIveWVdvWDwoG5plBb3nXBg+6RPe6pfGP8LIaF9
SqG6fhytuHekHOIeQXYbR+THgoZpG+yUytCrXExaLdp8H7Zb3AtntaBdpCtEjAYn
ahltIy58X/FrPBJqpscEuWQm0Yg9cPghZaLbMJkZ2OBB6HSMzx+y98DJbixOsOu4
IxIASg+YJJeTU/0OLOqpwbtQr+uda87o7AROcnsz/JNe/0gldzLOPpGe5RjJ+To4
vJviV3D5lrkjH9bo9Mfx0tIWcbqPz5Hsf0EVHp8jvh3OylYvprRYlghtJsdpNU3w
MAR/YXk6ulKnpEemEaqp7yJ5Wlrh4ha72FI0PpnCOHc5WEGE9ximBlyAjCaNAG3c
TlU2nZplmcHEw8EvWMHTzvIydCgxf/S3YbgJivoE8f+GRkdkYEjhu0WP/TsXXuuM
e2vC4qVivKMSB7UrPsnIdSDtG1WOPlxRF3mNTCZ9TnEp0UqCw1H51tfkDv3yf2b/
ZJPKkc1U46sCIOzikjxTY0ELXUk7gQ8+gy9Q88aZ01vx0kblvQU6MU9jBqyPufrI
aPBRLIKElB+Qga3Cj5N0k+b4uGJ4gF2WtjRnA0HDL4+/jpPiizxKiK3pBVPvYwAx
uAAQdpTaB6DHtMzABLn/VVJxA/4EnyBrJPG6LbpsKB17ti66mjflozlDL2tYCUl4
y6kFXzdBE8ameok4BBDs4mFGnlh6kJiHK3t8N6HaxAb0LyYYe+gJmTfo10IjPY4m
CnRUPVYQQKAWEtT7BA13COdR4/xrp0s9I2CAyXMDoI0mTqg/nveE9QzYHuPM7Wwa
yWyF5yLBwqci9JMa73Ii8wy2WtTH/4IuIA2w2oy4OJBO/hQgDfmYfTNbj4fsIhZ0
x7pqiGMdmhF3AGy5K2bxx5tqbSS8E15Jg+Va2uPVi3s1oe2uUlMRPh1HSCLEVdC8
tKdP88b+A+8JmkE0ptGNUaij66QHb8EP/A7VE8JrvGC4EUjRtt3EjIM9ysqfi5Ov
OA8/d+GhhZtN4LzTfPeKwBt6gwmkSWOG7/Uc3Tzob7yPa/6V8oWLlaaw3itw6D0L
f0+sYrqABUAaMm7CjV2GwuK1d/6nAnGV/c9jo4wpnWf/4CDKvZX1+bbBu3Nlz8FQ
wWrwQk3UuNAO0FgJnAHHWkCmHMMs4jCzB/oWzuzcYQ/yvwWg9A8Cz8ylOJWCw41k
+qGx4JtMWCTvXpOiIFgVaW1m3nJOfm3rnW6s3pStOKyDReopQk9ku2Y6EVve6Rcb
/40CAePgkq2qRU+UZO7bkpuNmCR4DtUKXLzzsGRcYqlj1rvp0KhXe1RwH9szQfY2
Bzbf58WyL5nnOBlTN9g/9GEYUuZ7ccts3CFIRAi6L7539NLCdQ7iwcuSY/9AU5RJ
RwlaCx+l3AvCW2FqFJ96iLiK5A/2w4Q5JPWpHx8jymKe7AjWL9M5rQ2uhcbaZfFy
hDgw18kyXzOiLKTLUYhQ0bJa3ak/LoDMCVzFvIZz5NTIR2P/uWqaflrjUP/dhGbf
HcwZ3umHiAnikD12elYQtJfgbwSVykFHE7Smci1QQsz/H8f3ynfgVyW9aURaI4rn
KzcbouhWe1osKe28oYnqhgBPFZmtf+WD766AZ4AKdw7Q2TOjyYj7FsFe2GXIwQnu
okYKPnqd3mvIY8uXvdE5guqP0zCAmcxlK+62PvM85Pq4A6ph672HRHxHXB6sFjow
t4+63PAH/jVUWYSP4xan+8K/lFQ6iACUrVmOI7zhdcOOktOBRjzgoCAcIKw7bUNq
JsGRh7NzRXs6vx05g/WSq5DV7+T6xuhrVnRVEnI2T3QQhdXKWHOsZFHa6t0FeCbc
i8py0q06DXQvXoQna7qpoBBrtt34mTW0AcYP3C6hex7AtccMGhUIGQoINDIQyDp+
7h1lVIEdCTfbJrdfPYaqOsXwpF+8oxusdFqBrdqYiCEJtXrvr39+qn8RrzoQTs4u
i2cAmlxqCEp7wpEL63PrAjJMFCvomHN8dzs3GyY5ogfRYAmo/N28kAx2BiZhUyku
jwXNDe54E3xEZ6kFgpOs+g3gYG7Ow0xAHjmbuWLIn9MyMh9e8aRibbSv+n27YSdf
2bX9W9hgkpwautXi9ZXiGb91WTk39VW4P/jOf88rvZPZD2a4+sVMpcPSC296MMbC
tw/+f46pwFHmotWM4YX/SVyVhuf1wAeyxlpIPlffpTzUIshgx7/ck5YH0bmEtV5+
GW7zNh6XpuOIzsaIDX1S+5O2J3DwMj7qfPNRDiEUR43AGPeBkEiJQKLScjc9jfLs
wW2M7lh75E+/oRDL1VoeS3zSRcmFmuseW9i4qhxOVaDBi2wehGccH1fCZtakCfS4
XyBN2I3srbrUSO2ugR5YT/sgkLBrQwTCemoJAagEcF0lM8eiTIacMhRIQUQYvan5
AUV0KI+1Uv4s9XP7bQrMCfYN/iWe573E/rReVuI+6jI1uuH8vbjzRCpHhyyeMK1O
v1obFQWvw3c+LpUoneBHwVBOdkJzqJEZxlOj+CvKLI6O5JO/T0TlZEbfFjRPxcNl
/wEynXwCPx5RYn4d1cJjPpyFztMPmmuWvpj9qjp3nbCxMY6Y3ac+nQN/I46+HL9c
LQ7R41qnArW1MbOFjmy5vfJGog5tIqW1ZRu/Lam/fbZXEllDmKcJI5i/RpJ7keqi
EikS/e748xPnwkaNrMqIdfuhxz1ytnmyURbPJj+X5YClWyxkbmKqMyucRMUP2UUd
doIRb8DbeGrjjUKxX9X5aB5SS8b24BiSATanhHNDmdRAZIQu73fu04MYj3otZrSw
CshGCoZcgM+oXRxhnF+hapwmTWPjXP1hCeHwTIQIaTA51o728/UmHBwCXy5Zq1UF
rsKBjhafuD6JOL+cRvBwnfBA2k2etcTQk5w00Q+FasQD6vRCbWEt2IKJ02m5SLE/
q7DuszUMauVS1NOD3NAIRpF+GUYywoECMcv0gnbMOiCF6LZ32scBuwyFjdZS2iUX
vzdYC4dgU35coj9oCjHt4hLb5LUkYW4t3I6jyZnN94/YQ/6rEWw+C9/e20BMh5O4
Gy0HOO6WOcMSoMx1+XD+8u3yfjXN5GsAtUkKJRI3Z8BHGQygKMRmkZlvzr5eVA+f
W0iQCumWYcORgcKUn0gET+y8N2oGI09b6E9hERUcNAk=
`protect END_PROTECTED
