`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6IKhFemFe/Lebyid0luHdGcD490yJsBJ80oMf08zAYHaOg+3s0P91a9neGcYIpA
XbzlqTb0mJFDyIwAgUUBWTW/xPxxROBghLE8XA3GRplTYeQwIVra5mPQm7jd+Wpc
sOxUcrLDA7w4UT5BN3438V/7eRBISUq8I5E9rxLi6q6It+fqD5ZvUFwCTJ2C+CO5
H6nnTLHmUxbs6pWE+4Yt3+U6ApzMj7RbaZUIuFIj/sPJo/GhN/k1wJEuvGgIVK76
0U4Q97Pc94+AaBH5M/HuzcCcYJjDy2NMbgANICkMYp3p6gUqQHHdbBPhfD4ZUnFv
S0BbfaZPQm0EEhA/+rQtzIrs1N/Q0S63oKHTIdJuv5HNXVPqaOBzYlCNhZo26CkZ
B7yB8+C6mN2/nrikPgETsM9DqyQJ1mB8m3T12Cx4JfoZtAPAK/+X/ZKHRadFAS8p
g3DpE1sTLuzLYZNGSQn33TJLt/Rft7MxUYnchMqQ/LxHbczOoSPW6Z+jeriwyl2P
hyfPTpOAgLEZkkEGFeSc9ou2wmDxl2DjMlZD+7UZBtPu3dz0qNaOTEA6O7cu9Qrz
+8pH+4UY/T3Z/+66TAhfst6AEwyBdSH+rlwtsUdurANLdrtklhK5JlhvGhS10UF4
shOiH5GXbzV0yW/WZjJQbPGZnUb1tp6o7x/azyakzh1XseQskYEpYMEC6JhfBXSW
6anTaLrGNU24jkOCQkDAFeEDHPyXZAJ3jIk565b+FHkf2xznYJvbZtQeJS8eb6rf
Xtc1vHmolDyX7P9KCDw7+vTA/40gPbuUTOlF6JYvKKw6zd8KyU1U+HNPbC8nexnp
oZeUVNH3bkO85ZaSvqMpIpmyxsSVl7b4VeaAuTOQsmddnyj5E4RTa3VvAmr09Epb
u5H2Sb5RA7Q0Ef3l8Tnybs0Ufl4z63pUC77VN2tiNY0614x4a90fqaMYRQ+Qa7JZ
5q8y2eANHIfCEwqv1WxDw+xpRJDUVYweY+NmtkRX3Bg89KANw5jbjyRHVe443Pb8
nIfwjvINDCh4Q1tfDjZbMbhwIasMUE++XsBTWYTNcld1mhlmCkCVM7W7XS6ADi2c
zeB7JBTK5pMWq9Nj0VMxthX+/Gm19qydPlqaEViKQxoEmu1I/+LzzMC1HffJmdcW
HGH9jvczH4UnmD3u7QpWHcAnvDYbPSW8p7ThqLvOx+pWflA+K5VanuR6Sia+nXzw
jPKAajRqBHZCl03gFEJRsDg3HI6p/i32KAoDInaAlPe90IF3UdF4yTJNsVx6cfmM
5+cYWqtgdvTw/OCDj/ERc3Oyz+0eTmpV4uo2jUl82pJBtdvvscvwhKL0hXyjVYuB
K3LB62jlrxlpd+KTUptzUgD1c/EYJuqh5NprmFMCuWl3g48eS/Nis4lKBs0Agnrb
`protect END_PROTECTED
