`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fxLEsPaZITd1qqeA49t4xjQuQdexSiIM++8RYMBhlsWT18g7e1+s0PYlmIgu7rnX
UFgfhQji5UwSCa5u67i8+gJvOUd8Tybw1yp27AWOajn+Kn+U7ZqBhGaADrMZHvAR
iPWcAs1OPABy7dRvk54yPzWFLJrljgI2PN6/KcduEflmkLwE6VGADJazcyXy8pbd
ER3GB+//Jktdsrg2vJVdVd/mZelMVC2lrHDaLCXGbI76JaGUsDqRHR4PPtqDLVQ9
peW4C5AL5UjDfi8EtwaEs4XdecuS15wdCn/IckflAtca8OzGHNxwIP+bW8th19is
nhF3bIjrdsJrnmGnZk+7Y+8pGESf97Q4Vgu4yv8JIuHPvXMLr2kMy2pL1GcNJ+p5
QE9YK06fkf6phIdtd0K2sg==
`protect END_PROTECTED
