`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CN/A2ttBagolkmEydBnXqfEjhcPwiXlNHQO0dX7pd5uA4U6Ou1NCbFWd0wYUwuP0
+q+ZP2olRRXJ/oNQJZ6pPWuPs7T8SfguOxrsgkbayGgT0BmibSVi/zXhA9VqWBbt
DYdEDlEtJSYp2c/UlIhj0tLc9n7MZvFllYk99qIHkqGCkoLwzXTGKI4apqSAsigu
3cGCTILFb5ZP9QRvRhd4ZZ5NGmI0o1fG/0aygItsMpaC8gfUAsj0oFc35xJkykqy
+gaoWD+w6unu6CsyuvSswxeg8AhaEbvkkQM5+KK7EeiCmsoESjMwFvVHNTJtVkqM
sUtQNxlS8XSAqIKDQvqTNzg/FnhXYSciJe6yiOXR1qW8NqNvfzJ/UIW/nv93NP+m
Ya1myy3tbr/k8w3lfCgP23TBwXfwdm1JKa1zHdTLLqNrlmZcN86vZJnToQ3L7U+w
rNqTlKIU5UQVVvAlQUej97UtDj3AtK6ofHbyC+icTF3ibrSB/Pqpsos72GIm7Dd/
tL73l2nKR/7XQLcFLUpE5YFEFsMV0lk2cdOOKLXuXtRxWv8bS0HZv7qkh6G/W+eu
`protect END_PROTECTED
