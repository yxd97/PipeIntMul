`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvIiJHSWOgbUpSfSW11sGJP3+SDijdEMaWP8h4dEAv0LRLPcxG3tsdNW7CT4DJ6P
2nXaR8fRsJA0lp1ZECaJdtmymhi/G+qBMEpNMeFd2mE3pRpcK43pLXCJEFdw/xVQ
6sJ9wJtHTvV1l/pEFyILPr28vooArJtd/U4vgO6t8llhoilMrGvlAZRvyIq7P8Mx
tHUhw0b84rgj/RpCOg8JgGHZcbQigr3l5IdMGdGn2LWi67n5t3mAW65igLPF8WEw
iGIhR0l4ZQCylzm0CfSxuv9ISg09c5VL5VFRqpfgTDvM6Dt25l+2LTvKqWONAWqH
RTrDpXhArUtdEiwZLoLoo6eegxxxt0kQ81Pna5qeWbUFw9EwJXf5CZh7AmjePvsm
7Dh7aUE03caLTJ4sadEvZtMlCTvWBH033faG8u9LwTA=
`protect END_PROTECTED
