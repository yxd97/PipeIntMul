`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqhVAQfs3nvMQKYQuVQCsVR37AJjYQ/4OSEvp7fPhGY+mrNMuD67g0CksnAbqFsx
L5FPtC0Bum2Dh6cRWbQ7CcLLpVf6EZenA+IzDIV4iW8Gn0opvddzaUZrpzVTOvWG
50nsvkgiM2NHCO0PoIiVdqFQT+SyWkXQtrl5HmLFpT4vSb5iftWqidy8Ej+VfaVz
d6CObezxqYbDRTmRtKjqlUTWfqtS7Ukoh4GxVkccjwBOsRQSLN0UuwcSz95LjhLe
BERzcE3P+pWC5Hypy2JyYE0dueGMVtc0B7TNCBkYe1mrQb7VkI3sNXnAmrRCwlTX
FSXr/FgFU/ShRBMFrSIyVOmygZ0fQt1cOfXVIZZQlr5HS3xTs3h5nXO2jP9OVaYf
ZDiWnMKePXcACmeZyn6daF/Rks19J1SMYwmnv0twNC+d3gzKUuflYT9NasxgZTTg
FKi+I/BUl226EFMtlGXFqC99t2PDwbfiANR7dgRBQfoVZvq+lJK5xf+ybQ20E9Yo
c0JHTPMgn6ALZ4qOyYQ/50TyjWbEGgLzmrCD4b6mnu+JPKS+C2JdDjJbaPLLgG7K
RMNv9mVDVRwrPOP4i9HNrQC2Wu730E/CRYBa1kdJK94l9cWMRw75p6622Xm+wHhn
15giztQRdhpu0Wp+6WebY5DJR+yrF7KLKWANYIczSTT90LYktC/kZo11fjlxzjzW
8EMa8oa1n+c4QXy6jiu6xQFoqDKgbdcRzD27cOOEhZj9ugpT7V7grEY+/h7UoMEZ
YfeL6s3BFhDc7SG4cHp5s5sBnDYU7k3mNAMcg4OIXwR2qe5XQ4WafECxgYa5IDto
Yy52MHhFOgK37bZ8rpBnQ6jnY2mSsX9b20eSsfEubwYFYcPAwhqvkMGRXEzsqFPE
e9RC/6ndfdFy4YnebWT5d5epy3AO3EPY68B1MzxLrkr0/Ml3/0r7+f6ciVS0NDVc
TbwmfD6/wZL6ioXxgR+ugA==
`protect END_PROTECTED
