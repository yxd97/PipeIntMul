`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
du/pL1HRU6KJ2EkrvyuHSPRU2PNsToSw+zWFk2cM2ntwYsfpFviUdlIk36/lF20d
b3P8MYAKDeeT+wIo37W+1Ek594ChxWIWPxcGZbUx0f5L62Z29shZ2HjR7Kdu70Dg
ObzDv4kwQCmEa7hkkxm+Ke06XHJX+jKibOT5l+drFjFYLNhG0ZkVGTwtljccgxyl
3B+f1SpTttuvjS0SCepyM7Ik1ZwiXaNVcK7jcbwhW4OiY22fKsTXRJuv5X2Ndpl0
l5czvGwIaxl4DVMM7ctXTcSAxB9YX0U1Lvh8k+F2EnTl+yn93Y9mhT18DbTdHFrI
BQ9j6MqGo0n/DjSsICl0O1QcxFEeKgfVW6Y/yi4gQzelD0n05v9FFrdOO0gU0y/n
29HngjBVKoB40NRyKnzKvD5pabLVOkPwE58qry0xpcoUQj9qMjGPr1G9+vrVNB/b
tJy/e1uZDosuvCVS5xaTSC8hMA3aLNpKJsMkCTbRgidG6yJrS64T6ju3PRoOOPiZ
u0lH0LJ/L29WqeoCo8ayXjkqeMS9tmC8PxIJhxxFLq0A90TFjm9n2x+UlzogaKUM
WuHcnYjxSd39fj/Sf3JmWVk+kr5MdC1RpOq/Lt26x4bSdI2XCbhnc89uHSNeYQBS
SCfLx4cw2bJfHB/9HusZxqhsdlUCwiYBkF8wn/J+XSw28S8NsYV/0C9uEGY3BB/v
2n1y6ICeWoLata5mC7rnCjW5xQLm4P2rhab9/AzX6tZhfsF6IDXE/iR2jhkBW3ZQ
W9osWz35GHkPIA0pf/kOAJRSLZqm65FQVdrzk3i1p4gwAdugWO2mFhGytIgixh8q
4knMO2oqcRB0QOka8IPEMIlBhBn7CdfNBJNmfu3zHVheCfVoQFnURZbi5nRVrUTD
cTLCTtgHHk/lIfLEe/b1IwQ8MDf0bREdQxeyL/cwtRrWEWe+fAxdudRwDmnMB5QR
mgHu/gqaD8DqZ44gEEZk5DDq0gQ3pUQ3bHwyABcdZeB918ZhD3OmZeYdBwuMfHaq
Ecky9AI+glAk3mz4yiiJ3t6dGnWvZKC1RGI/AOoybcNQS1h0+rF9yB3+0EK47LNf
wT02XvIRlNUAFUbISi+KqwSrO9rZhZ+xtZeSFNlNsJ/XGUZc1BSuVo981C5OJPqx
EUwc188Qc69KH0/pXT2fbBf6q0wpjgmgy2upxFiytwnIy8KkX6vAdBaq1iLOLg+/
Ay40PCZsRDQfjA7Q3xS0B9nW4Cr9+kEj6zvNcJOzEOqiH/DLrq1+rvsa2ppNdpy0
mS8Dm5iISFZ/8XQA7ouZPYQWvluXcsg24pDODwvTW/ibhVsT0DlkFLaKZcAQHM8d
CFKlTO6mO8vvTHTZaS2v0JQid50WJoM0+tNdYTTHXPNUtMMp+5bI/yJXhiZ7957f
dlsPBGHokEw49pv1o3n9A8iPtUfTiP91f08OcwXUmoCMgdQPkIRYy75KY/cEicZz
URaq2yIpIwn0A+P1KpDhgoFg+CWKoUIIShrNDFw76UETpy2e+RDt3t9Xu6jfhyyE
nVyZYePCRFc2IXMxEmeUHsW+hx1BW+vESzpI5xv0GesjS0qE2jWL1pEF3mrvEa2E
GeOhmDNtiCz86uSLFA8EVKQF3bZEAYdpIpr3pgeUoSbgafeCA9IPeQRJ+H1sjqnd
qVV0kg4SnbXaCjOPx1duO9/zdK3j5kLaBwYltmzolbdfpnEgrft1eHddzgDJMOU6
9GfnwVJg9wPhS6vLyXyDLRsdqD2PgCRTFewwpCyK9W1UPsOiKInvpHjXRATWQCl7
P/TZtbcMIjqaaAxokqfI0jRoJLjqGBT0x4lTOi9h3nJoysD6tmg0SkmDk3joc6WD
qq+D1sxfXuFtLdUektCKghWHD/OjS0qYLeuOUVeMqEP4yKYF/VCrwBYOJPdkW8Gh
Heg7tJUd3GpVVqlDAomH8/AGnX+hGzBNsEVXjGS1E0gvAAQHthsb1gl2vJefhWxY
1Lh26vsgWYJvwukSiviIWM+hF3eaWhpXco5Z3duGxHHWqrpebm38i5YZugmXenfo
p/dpmgPxerZccfO+QiNmJZQbzrtBAQ1vU956bTE8TFy53VecwTyDcTIFgYa01GUX
OTbv3fmnfYnMeaNFAiXU+M1uYVLqPoP2yh/NkbFRXKCJrMBhBVKje3x55gP2nLDQ
hQSQJ0y5Giy3DwSM8NpjR4FWUeO4MueXDI9HgjMskf2gqVBqa1udqMeEo1TILdRQ
w1wg1w+l5L17AvU5zo19NE9OPRv5s0cEQdBBRU7lDNC0tq8Ksq9wDko/3l+j/JUO
q8fh2/AXttSt0XY3upwehYbaoKrn2QoXiLdP2KTCW6r9nV8XBVnSI4mp+8xPCCL2
6gXR2RKg3pfpSJ1ffrlc7FVhqA1QdlkiHq7cieRJiTJRwhwWESjoADLipxyZR4bm
d/Z6CpBWV/AQdf637ULuUkNvJyBmUMN8ydOx0bgPgdg3w5eSbLC2/VvOOnO7nCQl
MKn2+pmtzLTZp2kKPKhul124WUFoINP9vVYZZ40rsgxlDI2s7+WLKZSX5a9zzAB/
3aaGvFyfGIrAVOPZeowR99bzDKxUOPF2KDtpaKZ5efdd2AYwqpN6SC/3yaoaHjz6
2jwPwnAoqo7CQf9PxtBCMt7b0n8GxMDMGkVKs8xk88qynstTdpo8/LxlBGSC1M+N
0/KvizTJKbLdoqPyOP+deXLRt+xQGhdsyyfVVNGHqC8Z5Bvj5L1MNi76CM3/byAu
00l3Lz1nYPqa03VaXea1eu+eekcC1txxPexLNyW4gsiwYrh7VGSqgAe+qDmxEUFT
jL/6+Eqd4UYAjP+hcJVKX8emNN/xxgaD1d5txrCiSxz/aRqWZl65dE7xg2w9Fc3N
iD/Zex9+ukY/rzaTMemY8WX7Fi3SfFvVFc95+j+91I+51ZGjC/dYk9mJGmWvqNne
rK6E49e/3pYr6bE/xip/FjQqAHd4DLS1z+42T4eur2MaYd8nX1x4O7KCFKpxHrNh
0cdIoBx1hLRORq2ZLJdz8/Yt7ilrpFkWmvOLbOCdW82dRbiwSE+wvqDO7eIPECXm
MZt0vqnr1HFBeBFQ9u8pN8ONtqG3W8kFAyYVyNzfJY0zXK5IIa+B7fmyOnTUOz30
0YsPyZlNpPoP6opKEakjUooyoO2MW8ToGSVn7/txqX++q+U88bH3pj8ylUnI8r9O
mAbnqqpp29m10ea8smXQ+/6KhcUKG8kwO2nAoTjAs+kVzvBaIA4Wv2mU89gg0Ld7
W0YHQR+5pRgqJOktr/n5iXI/l1QWEW63AqdKHNZyIxRDOcqagPx0Q9KMd/VPs3YO
ex18PB/F3iLinkYgthyKAQ2glbM9qXGLuUGQy/gnniUvwiwBktKJiZ1AkMzh2LAh
2Df6LvtDONJsHR9fBMX3RwO7/zGyibl+QQhu/HERaT/KUlWo/gr3i0YUr9zdCO9t
1V/aeh/o4KBDeHLDgOjbPPAHdNRx8mguTDx0JgvVz07SP4wR5gM5ZwdTJYWq66dm
q2kDkwjGOzQA4uIyfI7P5LHkZdC5myFVI+I1fZvePsR2vmNigHHuKNfmq/7x0d12
fKmcJYnQJsHWhCHTZAZpahFDJUwbPbcHtTEMhs83gUPEfsHbCVSfZmNjDdfIlq70
RyKaXSe2EoXrPHcYG/GKF0jSvPBgLosnJvEVME8K98nVXg6mt5mCpxdPXCmDxwd1
L2695Po5VZTYcrlXuorjLbkxrJW0jny97crtnlaLvn5z9ddWQhm4mo6Je0x5T+gE
R7hgmY0BiUl/1XMYIkW5v8KvxdPGa3guNiWmqc/VkF0j7L/H6Sn3L6hjFSJB9RdB
YTUaW2W6BKOVcz/SOQJOO85m4qoyEWayFhYetX+89tS2r9ZzFIhnVdZHVFrlPIfe
/3RQE+ZFe46Pta1i0D8sCBQ5+Tzf2wArU089z1BiaAdYCN+YpaovhjOPv7GCgsPd
85r8UYoGr3FGu6tS5ecMKZpqeGIEn12txvwXQ5jyWPh6eJj/7hSh9QAJcpKmG2G5
KB/CS9XZpwr6Prq95Ilcfx2SRGsgDV7S3CMNzNu41kUDdGSdPJChwrR/PNHVAHoz
BE5B9j+PGVug3dqXTK5sUfowPgeeMrunYEWSqbVuJfOVB9MFo9IpC4fHfHTOhm7c
nstBDKmmLVEzRlZrD9FlUh6FLBIUOanH9FR5Su71b8kUPZpgfBjk5fABwcZ3pjBJ
Q+qkThMSKQnmVrrqSmnU6ilmbIrWkAPy6I+a225VRJjYSmNdCYi5Pcxwmjvz8ZT/
KQli0iWdI6Vg1BSDcawNcwZLQZta2TPCFP9a5iEskdHR7c0fkpMlO1RUGa6V6IaC
DZUhklhejIjPI+eL+DOMcsQ6VM6WAF8XOpF7hSaBA+R7nh/oHjSdDg97SOjFiGaE
ZboIPvhDbk/5Y/wMebC4yAu82OZqIm4gqNJGYGVk7ivwkoosPnuhV/QjFU0nfEDX
kc2VHYgwsaPKXwwToD1l4DUlJA9vlfXJynZ9K0XiaSmwJvNgoXf2lyGBeKoati26
IsAV7f8b8lWmBU6ZEU7qqVxkx53+WskhdTT1KIdzhSUEK6ltu7Rc4O1vlKJA7+2b
+pYVg5NR2+IFt4P3aeiE5awON1m8g70ivdPAuoe3BY+op3Q7DSlp6VtP1r4bWwOP
HjAm3p2IRbdrZeqXRpjRmMz4fkTZA4u/cd4Cd+w1YvTwgIOJoGPA6x0B91h9a41K
m+8E+vRpm7D26+k8uzvVV6lfHbQg/HfSXjWMDrYQ7W+HAwV1WxnaQgFVx9/fvuoD
fqhcTCCYz97OriEhItZeHi0Zj0Kv9mLyvLns5q8VUFq2crlDiDzqYo87q9WU/X51
aBzzhZEwrmPuE/jLZMMwCE4pozMfo0z1EWB//Cs2J5rBgU5JINhPafqxeXDjZrn7
pUbwhoclF43EgrDS32mlTSn0rC/XRRDVgeiMHY2r6NZpiGLzeahmBnRlCPVai7O3
91xAgytUa02Sj/CS5uMKYvZ3fgtLH2FDg0gnoNZxRa1fG1I0gInDkprGAEQfU5bS
NEsCjE026k6YVv5394kEJ4Qj7qruhbZrXg6QDORkC4Tv8KS88v8DijM9wX72wwWF
JsIt0pJn8yvZpVaMMzCtPt/IW9eM1DQbcPJM+17STWnA+VIe6U0TL2WsgNjNWt6A
7gycirhxqew1NtO+JZUKEdi5GcXNpfDzLkG53cCmbK2eFPSHZ3O9TOPt0oty1fcJ
/SyjHf0MsJUJ09YyOLchxUt2iXiPJIVr5rJP16n8F24gorPcXOjWIkXqxz73jXS2
oIpVx43X76xDhzxJqev3rW5XqBHoPTvoypCRZxwxNPSxrN67SEwpPz6P4WFxaWFX
QqDQ/BAK2VahyMR2M3SEVumL1vYRmh6RcMzLX51uORtkMSPdW8ic08khsdligHgA
xb7LL6IFpdh8Fx7o7983b/VmImpC7NM70oABAvurp2Rs2aV9Z41W16J3c5xjycn4
KLVOB6RgeXtFZCl81T23BphOP3dKSGl7Zj7w1/0kHYgUxOZmENtpasvPmN4TwSqR
0XBZHB3GRGnqC6xxFtgrPEKGG7QK9VeqlOqyCd3gOs1Ntwz8KvoBJVwkm+ttRKPN
zmiwltxZPwsaL3w6rQsK4FNNqDnxQdtP5TqDLZ+UcBnnEQqCsS+UJIimb9tJCdzC
ETZCLzi6vFh0imqHXou9XpGTq6kRj/mnt3HH2oNADCi9WgHh2kGWBWLGYDrof4lw
m9UO8Z6YQY+dpLsQweEploiXqp24h8v8kdefmRooy5UgyforCvJdyTyfJ7z63MPp
nkS/j4tfuGmJt7dja400Oi46fLMcusYX13BlGFy4R9fSENMEn0PeKkUDni5c5e4s
e/dwX1BpTfW5KVu5ImTxJ/M8ao/o9ojAkdKlpY+NykjJMAXdPuKFfE7Q7uchvcnO
pM0Kn7tt0ttDpPaIaz9PvC962eCw+694Lez0odwG3AwcPVpmFf1JASUKy6A4zFNB
8U0rsmZcQKFZUb2NJCFIqwzYu4cJXDA6OoLDZ4AXb+mkgp+4Wl3W9VWwDuTJLumv
aVUei7iWx+W4ADc3HGD+hKdHciGrO9948PhY4fpc+yDqXAlBjkuF+F9Kvtjl6wA9
t0uvCXmNc/Ro2+h6MR1SSa0j9fqItd4RdRX8lphk+nqwkZsow3p2C+gDjeKnFp4L
Z6QD/+sVWz5sAEEIC2u+Rwur5WIAJ1s1V0Rlw8cj+bMGl6vk0UVX9NnuVUbxwVQ5
IYrQeFZ3xOUcqwk4I3t6pXjN5Au/m9RCSaVojiho5EhN+rvnlEBCsCieuGT1wbMI
k9gbbLqCCELNb3/7F8FvtDH8RfZvKVasHzYSW5Vee0M0EJegwmDLHbBndyv2La0E
jA7Ld653g8usbZL52VK7XAeXK2rfA+gpeb94p+uJHogwjj0C83RLDJSpeFDAuRlt
tQkQVvx7ydmzo9iak8PQUbClPEXSxn+V53CU9SMjsE5hxyL88E96r9GM41tdSG4b
pEv9okbLYzz4T+2tWAHUgFJJq13q2t8TbrBgujr5eC4g4j/+89rqCdcisVGoZMuh
5z6zjwGlR1x2/VLf29bARWAphXb9TEoghiEywIXnlbDH/XEtgD75yfPBzD/0Wu9y
+YuNgqNpQv1nGD7dTi6XXLEzAMNM64SkX/XrqGgN+l43GHwssPIDNg4xHZhjnJ2x
AIGrW7O13LGTf/49XE5JJAV+Lk4vZDTi2xvN6yd38TLKLKjoFRRdjOlCQ77ckfW6
wojruCshRMy5RkylJRpQmjseyu1+JmiGK38fnfcAl6wRgkgHVZEt/VsOBKzEQZSt
NlYbD7hOMClTUV3ZInnIdlhk7BO1DOmRof5ce+o9nHKUCmhiHWX9PyE/GvUw1C5O
Zmu6R/WAUDfK4yFuiRhjreAp+ZgE0ys0vAxUYUbdZxNw9MP/ZJPa2X/YmkfJLSAa
5m2jHOeDz0H0Z62qNwP4PekjGPpW/R/yo4M5R6yZaYYW8Orw7yLGe4Rf5o8Vjpkj
tu6X77U65XYz4KRQsKg0to0N27D+RhuoIigaoH6vcjX+7V794IKLm/DGunLdsQw8
T9OG9TT8EiHQctek3c7oPAxbRLilqKHTKb8BWkFX6cKgyFC+ILSSAT198/g3hPjP
UHcAR3nxgHsRd07gru04+TXw0I8fqOtJnG1BwbiJEvlXO8VHYxmbQ28Wjrm5awCq
KCD83W78SD63/52KTmYu8evprKJzUN6TaV1I3ukWd8gX+xuKRMYCUe8XSb7HFhZV
Iav93ncT6NwyU7N3vRKdDdyk212oue5kfHq1FT+HmpNo/hqTz8Odm3edWAHtU/8I
FbrLCM7hchLcIKhHqw3srJYOOHpfSJLIxdukzRtGbEt1dZQmah6orGIBzAezjWLx
8wMVjl2CLYksnhOF74U0SJfQFGU5XP1xAHhW1Piac9t/4FWTKKwD8pwiiF61HZz/
vXYHXh9yTRwMkJUHbh+wMRljc7e6+6S8bJoHiSMIGYgBHYV/6F0jP2MhuF6vBNX9
cgcDGsUtyKKKCS6psrTryw2XkQ1VvTwPgdW8F32CC9pVBG82XWeFV9HmkZU8gp24
CjAhvezcDuitCehPEPraM7PnR2omUvoW6fepRoWu2UlbLG8fzFxGrMLbMsxj9H+f
9U1Ba6o0lnhoIUYuHOmRGxVnM7Ac9WjYMCnvmC+44/GVeSXmQINO2pmdTszo45Lt
vcRPNW9qJZtEkED0rrQWFcUPZou1vNdEClT1hrdfHfzyjPDDESTafNEflrotlw5D
hopnP8qjsyODaLTIH25+074GKsSL0zQ1h16RQaRf2ZlgatGI3Vq06LpIVNjB6Obj
nxoL7NZ+DD5pz/eg1VDAl3uVM5J27nAKtNBfobwhJ4P4ylf7GEo+2i15QNZK13bi
0S8tiOjMxbw59mU6E8c88Ccw94fS1tyns/vZutBbmXhjq5Whb4vszik1LdnftL4d
rcJuGBPXEr6Rf2dHU4JIEWN8J0rbyOa88H581nyltP9KYCzYwODUww05Iid9G2cV
6Cfn0AJQmpTUDTqzKxtTjda52jo+Q2EKK3EuvB7ENAm9XPiG4rfPG4ql7ZdRZjbW
N88haEILwFadDyG2lyrXlDXnhNcb+DKkQtKn3AXwtbAvap8VruBI+STgjPYVdGIR
qNtj3DDdKHBXnOpNe7bCq3jcCz+52DONXcN6vArMbf6832bA/hOQ817kLXQCrPTC
kMmJS2AIptakrFlUhgHe+pB9yOL9hUOySIekp5XAaNtKmzdLC2KcRGDH1qMSN6OL
Tcqx+MXDN3KN2apn6Ghvp1qBbBDV24K8mXXBw8mNOy3S0zNljMXGVtoM751JCPfh
EiXgaVwaplF92WahP+311qirseaPbcyvDzxBU9pWwnYvgTYREqwq/KH8gxXQlDWj
ceBfG9yt1EP1ueD8REKAnAvwvFRuDLxsp0+sd7vCrdAI+b6PRfVxi8o48iQOT8Hq
pNFcikEGIyhFUHU0nv/72Poi3E90+XmJwTasc7DzC/2MzxeAzvURYQfUQ8mQN39L
oF9ygb5mtdEI1B8rItAZI16bp7/AsBCcTKQUPgoAFhGZtSig/WZpumH66lJEqSHH
I8fP0qlAaOLqi8KGAVqLS8xS6PRs2t6YYHhrpPVBtQ+CQ5jLvBrkJAWG8WCINIeH
q7dXFhfS6fK3nmaaKz2Xi2EC2oXSVDyB2HURd7aURaknNH0bjgYISyATNGkaEFZT
95nXhfL3NoF+Jq5jzYVtqduSR9ErP273BMfnA0m94MZtZLZFYbykDHqlncMs42DN
27b9z6I6mVj2sRUHD/hx6NseYKFsAuq3UQU+v2Kv9Nr60KEMcc+wnbw9pIgAdSCr
80A2RcbPPF6uE0AFpz3vOlyamdPenvpQu+DtLspEMBTCKD+rPcCjliBT+Nl7VnGC
ib+4tN6KQPtqTV+sDbsNc+ZYJy4g5gD+KxV5qRIG1N2crkFh9U5aypOSa2euA4jc
MfWcuSAS3H3ygv2iVO/PCrEawEScAzHzI8sbLVG6l5jUXgK9NmKiaxXkJnXc4OrY
/jQgbbcCgy3+t5E2f9ytNqehE9+W7iUvj7yrO4BRxU3QMbihmjwDuYjUdmq6UY1Z
oI/SJ5zvfiazGS5ebhbEJElqPSnJzRRjQQ5voMdMlErHbovRpqDPwxUf0A+mUSIg
p6A8CiKTaNEWosykvtiq43318LiJi8YIRN4Otz+mIO9vx8qLFQqsBUXqbwTjzb3S
Cd0ZVakJD/Bdxz3TaFDkVcBwC/OUwpcJOnL1GDUx9IjA1vUPtFLY0hDT7sm7uhl5
rgYpN7Qg0f18pwGqeGCKYnU/88JL1n6TJWGUFWIjv33kLxqD7ucnPBVuLkrC97Gn
j9/nKIp5wbQuqk0bbWLdC/xQkMuT2gU4v3/c1ZA1yEr43MVdFr7JjulmmtJu4Cn6
p3c124JX1PtDVq1IpOZ7Q6C7d1+7HFIk/o+mnUJ/haV9Cp9LBUMNAWCkH0k6y6jD
WYFenUfdGSNmQBVLgFKw5YDcPSEnJimkSthmK/Mznvt6HIwzHIA9RUjCkYniIEtK
9TxrF6IgwDTQzMIY2VaSvohhTLwd75ql+mzFoH6aG8P0UjiIb4dWgWohIgnNCAOW
CYeIqeeilfW/4QdHu2PtCPOvzSM5ELCuUPb0yFrltIdskhiTh2MjzsAaOYjDAkNz
9Na7rXKmGkPyOzWP6hLTz3R6aKx8s6i+A6rbjkfX1sOTd9cKhjLU2EXAuh/Io87E
pPVWoj1Q8ImGsbaz00ib9QtVLggUSKvddTqsskABCTq5F0To8ahiQizRwKcV2RqM
eZ13exBpSUn5MKdUUewfoocB+anp1WAprkDIKNbu5wv96PGkyke2U35PfpiBSy28
PUrG7Q0po6Xk73iYvQxvu1zun4mo1E7EP2H2jTrBKY25Mi1xpanGh8BSGqsXwHIu
0nxUz7NY+hocM+v9/YUwhTa4hhuZKCfDweZlzHHOVa+mLHX41NVkkJcH0T0M9Xs7
8ldFS4NMEjFg8cRJzlde0GOFz8bwaj28K9pAVIfId40r/gPABPOm8KmOaYlvIrSq
K+CJvsSW9hVbw4mdV8ZxRTOsYkXgji5FTTaKR7wL9BXoqJhwZ1haZZAYIDIe/klt
CNe4LWyx+XLTC7jlcxtJu1dFUF3zei/VCXscR1OIzTQEuWyWXsHEMeykZmZNs/bq
9SR2yznn6wHn7utM9ZomhYsyMQXrfdQueqdQPG/VznKpwpVH28MWtaEuoJav8sbA
7uY1PEjww0ZgbCp4toUfeS4f/LXAyBIPOMCX3t7kIvPdbhz+tY2f5CYFTxpQuLY0
pVPKos2RLTGwyBiekRldVmcxsBHpJGC7ejOTY+b7NZ9l9Ko6MhPyorB1bIF8aqAq
wWMmBlAyC4ssAmQxUgxafOD2b+P7H22TALjC46r3wS9KfpfHBVHTQOAcHTwA/Z7x
HWEbdnTm546ceRplvCtexJnRWvL8iSjFgJg4zSxYOmn6hJ2tQckxLmJjMyPS8ci3
lua40LfrvQsQwvydhNBVUOK7mqOl13sN/0VB/jSYI6r6f5lMOppxh5ZrnoI+dnDE
62jQk9uhQYTrrw+PUgHAaVDr0ZOt/3Qj/PMHkn5sNl4m7TWZDaou1jhKMS+hJ+11
Zp4jzPkj4zXxiQVqE27q/Dl4hbIYiZJpl8iTgaOVm/MhHQFqzNHk5Bh9v2FM6RQr
2BWZwh9bAemBjkA1nz+sE+EFr6dUTzLZqn+Yt+EgxPcBdwtwM2fjARUD2YD7zvfi
DFblghN7LIOhYfUZHMXsbVEugoXiAkeRhoTNWzmip2iHtKeDHRpu8JZQnRNa/x0/
1iLfjmMjqtWjtwAPu1VRBHuoYO8HoxO07eejvHdgjO4BJe8vlSPfdwKmmC6pWIeE
EfDmir2VOUZPA7f+k5f+2y2Zjg6ZOUUwemQk56Hy7wQtt6tbzrEVs1M+l0WAHeJy
GNVyOupBMREOxMcdTtzMS2T/JETiEX5PCW+bxK0D3UEPCpIutN5S33HCEw9TPKLO
Oj0UtBzmpk+uu+MNM2AsnwteRVNi1McETPWaCTN1Qjw4yYSBD3Jm+4vy5vryT4Sf
dWzI4A13vzJIaVjceR3gPLHjHjZWHXJCnkMvr+/5SPSnnrnTR1gjo2nK6OlViY2y
Vk2es3fAXpVJ2tTwuoa2dOlyceMmeNmuY/TEBO+efKH8e87W666ASwjAGgYiI8ED
FQdhmDf3sYUcfYJzmVaqH0CQSl3aOu6Zr8JXXFtEBprkEoDlh0flv/VZFJGQiyuA
CFCHtqzPTggxmcy+je0lpMp+djCYYUh7IjXEb0RQ0TwtmxYD/4/AN9NYG1PWo8XR
CxjvXhc5WZyir5cObnPxsZy82ttNzZem/7Rrv+2XcZZw0ji2xdyzKhuP+SAfvqtK
aNqZgwQt9325qArF+/UeEZGY2Rnwqo+SkbsGx9IAGBU80kxM1iZmNdFiYcXmnTRe
3DqHIo14XUetx7fR29MUrrpZvgSMzm/5JesseqQKQxSAhsTamjLadw0nC7D/ZNow
F6TwWi50jof8UapmQ4ot3QO5obuwp5XOnzEV++2cbVie8XI4pvdE17q9r4JV1vIj
VtMb+z7Mvo8GmVWj6wxxKMIf/QCyT76iZ814XV+fNFHQ/XWUr+uGnUviyLk+WG+X
ajwbBDuEstjvOxmpTmeQZbgOwVkG/IkHMKRe68S2ay1be5Oc8h9+GVCXxu9IGUey
ihOShIOx46YR4RZr3/8GQlws7dSQAp6VF5ERoi7IWZ6A1adxWNR64EMg0cXYwxnf
ElxvBpUgnzAHngcI088uE32sj8KuakLlhtsko5a8w8TYbP3Z1z2N+tXrTyeojRfs
PItHpjHww0Isu+VKZ8tzM7HKaty0neCD3QDF3z/2/BlMXG2F4a8h9+4u7S969ia5
5ovBssz9VyvORUN3M/+jtwsqsk7EotsHrSR8vF7CBFx8/pD6aUD9DszoinRSfX2L
5ogKKvVmml7ws88yQCNbAKM9YckQGJUsuey5ejgaZWU+I7Q4vyoVDJ/ywDAzQvrJ
5vAwY1n8daNZHZzDfiW3xk9NG6e8FJA+IXhmQnVimYmUM5fVygMWeDXc3F7J7dpM
fxlcVRcpOSdXUwqDF0RzChQNy+rNxqc2cx56D7l9KIT39OeL8JdUIQk8Wppcb/py
xg4g5q3FOlglMhEqIzUY475LoS64l7SkW4Hy5bOXyc329DW3S/KcQ+awYTvwYw01
DZo6qS2njWIVY8BxUQWFFE+S9/kFM4Yf2C/BNDmbzvUeX6P3jbYMxjBTS49SBr5n
j5Hl+/Q0UnryMAqOjnT9gim0dVf5qze9WIUDo7IruPJbAHCZtN+UPPapymPCQBVt
ozV7ujJRGBxWnQI1KubGpnQIuzjorHNwJlv1jiOkjmBlTL2DQnCbAoeqdAp302dy
JBv0cme0RAAvKudpJEtAthyBfamqlpl/ReSyT856ll42CD3nvIBL/APz0VdJITsr
Bwc/Hc/PZNjCgtjZuhNTp3K34ThEnV3KzL1i/kqJEJO6K1eYS+dg7gYi338bdBrG
fSjMuMB7bYA3Ls4viIRXOwyzrQzt/Q1WCyTT4M4oyoix+tKVkukzs5CwUECTAgHA
UjYTpoKzfwYX6Wc72gDNVBEwU2yD3ANW1pME6Zd7+mj1rfyn62rHH8QOj6tTq73a
rm42+O153nxvGogfUwsIMnq7SDDbEzAQJlygV3RTBWy4uUMDXNUPTlqHF/ryIHv4
hyO7mOHCPseoIUHPYGMreL3asEiWWyxknwxI7nOW+67mNgq7hsdWaaW9HtIXY8jA
FruM283W+ETkr8q5NcMmwStpep1Xnbhg39pxt/9mp6+8wMuX74RwHO1Dv01hXl/B
KDLx5UfEDo7/FQYCm9SFAbJT8sgqwNjTSjCFwT3yXOAdfK/ta1z4D8vh3kKJjtjv
0rEDCLguh+e0Io7Kgy5/qNr/2F9fIVxAlVX0S880HoLvNso+54+7DY+LCUpXKSg3
BFB+w6lZGbBLpDu+r3yvRp94SLsbitXkF2pfBMPs4upssgYoqWD9uy2qPjMuybOo
AK+7Fk9Zh639+dHv93PQsit7ZXmrtcIX3KqiUBaBF70vVvFFcINiu5abYLCYlKSR
4NKIRmuAShXQ3l76Xmzz9e7qVpzE+ngiTRMZUH7kqapbCBbXUJh8+xIUpUjw8qwu
DJWukfUjx7pIZwCXnRtzVnTmvjWUJmW8xe8+WRKg1w7eIifjG4NcbLZ68Jdi6043
RlXq6l9HkJHsoETHHLUo+LnkzAgnVayXYg4xp2p7lLcfqpZC+cbi0BRZ+yrZWZSe
mtoq4F8RrDycIHMp01hLGnrvF2wjwLlwErtVIsaXDG8oBGc5hJaQOTu1OHp3nEG1
SBjcHDTpTi+tM3zIUn5LU1QpSjn5aQlGlmV+vIE7WJykHgtJ23YUmo5vdts1blXH
air3P7v4a/xp/w2kiJ28TujU7evFYDjCF45tje+5RepajKCSUASeHStPyTTxApRX
mlW0t/A2AE35q1ZDVDtEH9UfG/yi9gRT9Lc5x8DuvPr3d0bdo3gjo8cu3KRSBCVm
ftnEL2Kq0eISErOCqqdKXhphHx2/nYyhgAlBAWLfoX4MBTy8jGY04qniHRW7cM4F
ePxcN4+5+SzfiKCpJstkLMtsMBF34wQYaPCQG01cMS1u/sqBuoGFP0r5+8sN6KF/
CGCTWQi4uGzzAwqAOX0pDyz1TuJSfpU3eGqTrBfirasmbernsma2DZDaHTGkCg9z
UOC9dyjCbq6qhoDJbiZvzCXUGTmizIN54rBw315f5s3Obu9dkVg14NZjyrvZODlN
wzgf1e51x1g74sKgcCM7AA57W9hYKexfF9cqTaTS4ZufzCw0NKsnQ7GD8P0JqHn9
4PXWWeBRHposM7FwDQTyy6SVzPCJNGsgfMrbul2XbpebtUIKfQ/A/+tzhwPah4F+
3jz9+8pqQ1gPdDtsCtmVwq3uPFpGyNSGZbmezBwBTQTyCyMQS9Xr1Ex3Er8Bl6cQ
19Rixfu3pr+N4cRVoQw7bxn8sDrJ/IJGGHivqast5bv8XbSQM6073z+KWaDOXIRF
eybuEwGqTaFGvyHYS8HKmSAE4jBN3Do+xxUYU/Lb7NzoFMHAA1HyEgbYDKH/fhGz
TvCLeX/8F7deIlJJ8bdauru7662W/VUWVfi/q2DY/UUMEiVNlGMAQ26IgDXC3zml
CXgzkzrMgnHZxlgt3KpYIyIymsJg3/SCn3EWwBkO6FUshnM1/qXniPEfGCRTl0rp
3/W+ocuSf6pWKp8SWfWzQCsbW3CM6sdU69sMC4kipyeumYDzkO2tPu9iDtzkyy6C
B0JH3CBwBVYRgfD43Hvy5ZM/fV0ksAz4gmgNbAOBpkSYT6ddZADBivzzFvUwzHcV
YR184Ch0DiYlxoOvbGKnZv/rcvnMHH8EdPTqKvcKKfWqlpi0Cc9+/PUjzLx+l413
dumy1HZnwsqOPayq/ET/Spl8tCNSGTVXy2exPaXm5/hwfVLb9knta804brN/eTJV
XCKkD/TpS8D0AukaDStPcoGQ1dSmmRcUsbVSRRtUGuYsb4uTf2WbxSCCuQwTVxRD
hNjN0B+QiyPOMw0F+56p/PR585DQ9VdrhEQVE3Lx81s0Pyi1HkFfadjjx5ocbMrm
LL2cDSECPjEQzT+sJM8vFRD6AiYP2GT/r6Igh2afBFYKz/xpeCG24LmCsg4OZKTW
RJSdHTA59GP2HYS0OJ/AHxHlFG7+i781f70CQPlsmtKSwiaiWO7bg8el07pAL+FO
MhC8pWT2Ljt6RlvcdTbF6KaAEK/sRP4GdEMm3a7Wv/+LJMnuAUGXA2rB1jayCJxT
oYTTsS75D8kgTIfrcfBOeJ/oQzDy/XcBfb+YLs/p7vhWXC40eDmg2QLHGiLQZggw
py09e49OD45u7v/dp4s6/FGQ6A6HxPOib1URtoA8bIorS2QN5rxHxp0iSTvtc5CM
uDSnZ9PZXF520JONok6OHYkxNc3KaHrIACbHNpzUF+7MUayt5u32276e4NzUg7yv
Z4T/8tZTrsHbm6cct7czbXmPmlTHFpXKuez/DkVYMFuTgABi2J6IscGEk2GnFDj8
Q4EQi0OM104eGGxC8kBI5Gd8E8n/8FhAuxv5YxxFnc/amhRir44ML7ZpoW4XHBjL
myTcXPmC5FPDq3NrX+G0wwwfUhISooR2phP/sbE1Dc8PE8Y8x4eUZG7RNh+V5HnJ
eeXeKRhJ9j8+YKStSWDiFIphGFAgL5daTpidcfuKES5bTA7w17XZnxQLVSrMjBqq
xMT1Mf4aVK2r1uDihzNNb8sUqOHTLPxyGpHA0Q228oS1hNaLb7CxpZC/EvOVyzr5
32bDrtVxHIc8C623cSdFRoAGIuq6L3aj5GftjctFrxLrfTmQLCsF8anotzt1i0JL
hL5bus3HrdzZwgwyl5Jljh7kCwqU6Z2ogV5uCSYKKUO8+CM4jrS0lwzCVLHBDfOe
ytHHZfejGBsdh6fFEXvs7iKBB1JBChCYxwahWhywXVCBX6OlgwljQjAIJZtIKe1e
9KGA5A+5g7tQxCqF9g3/Tm3N0j/8cEnjTBnhgycC3TMCY48SxMsSBsik7MWPLOgV
o93NkwzBWd/us58JYiN568zccnI9Qbu3usf/HgRkmnx4lEbeiDoSRA+GRonuelWT
qMqSuiTMsgJPiwmmu3+ZruIHkdZkvJQM+vsimbCREEPM0ivsI4Tpkr1UHssBkqEx
lOGvEZG2uaIDaPQVB31jQMnxBJHZGs5QiRvbw3y0YS0sct7+/xzifVY/qRa8Cs/c
erykaV9bFH/mZFKC7BmvQ5zBakvPyTE1Ljc5OFwU7HmnU6JmUvB+ZWZ+njWPaABr
5xlblvH9vInzVpR2ek4KaGcTuuakNBnevdB+V7/0Xnuwx21Us0rQmzZYvs/zibWb
B6aFD9ye09BYd6nWNsRY+u7HDj2QNdrF89YsDLwcQ6LSvXtt9rdq/2hRulLUkK2b
/xaHm0IAzY0G0wi6gTRIOOO9n/f3XWA/aZT2n4dB9O8AQswCga7QsNSdtKY106Ya
Ay5hZzj1gxILuQHwAGGP/Y/HSU7XaxFrXVeXHNrgjZGyWcv1Eh9/cK/4ArI/NhPz
ImlCzibJiAxqhvVSrMhntuBILpf6Pw1beB0FEhqHnm7gyPsrETGPis4BjGqaiiA0
mQ5ox7OS4DPFKnxUNRVEl3ZyfEvWfavm1VBOhdFd5dFJUdn8rbvr0DWr03j00u0w
zD32MmlQNety3z45qkH4cSZwjm+2NqQhe2pk3HbJrUboZET2nJcusJj+yTt13sOp
JtNYzriHUQ403Q1iJMt6khVkWhsJaAsY0+N+p4ue+1azmPvc3yZA5JQouHs4LuUZ
f0fH33WovQHHOQnGyeVdGbEFhCuEaexOrJw91TziHvgaIFgZRRSjrICfQW1SCqck
C/cswtRRCU/rb5HuynQK2QvASp5MjsEvOIS1QuuSypYOT9PpQflZOLKKxh+bCaIh
yqn+IL+3UV8IFEYaDYwWzs/T+9bAIK5q7Jd/Pbi1u8ejuTpSYYgpDelP11xB3p+0
SdYIUjdKbuAuECVSk1nx6UFgnHqI/G5jTvW2lrizUI7mB5kWTx18K09MA/ySH4y3
Gv1u23vhFzNkZSirsfeC1UrzOQ7Oq3Ds6p6T/976wMn0VLuPro71PKbgNBHNXz5J
MTST9AyKfaxrsYaYasbvYDabKD248oqNu3bKkZt5b8i2Imu2xrp9vRdi4PcbjNnB
s/eWEBIsr2MELkNk3AlMB8G1ODzJPQlOQKOIXhKWJRb8eKh2cmq4PsTc9BfnAzXh
+0Xc7pNkwDbSvTPM9e9AmHAYrog3/pZOmiD5aG8BKfDSs0iQEuTZnSeEA1CY96e2
0BsTnxtWA3JeFW17jRit+X3+rdQ76r2w/5bev9p1qruoN5ro36fIKQdbVYFLF2l8
C0OMQYr04Vy08GSlW+Bwlj1fdvvkU/XjsO+H0IK5I+eIw3O1oMLGTd8IIcmDnCqH
7x1RDgxvuL0k1CFstNLLYGf8AHFpP6dEQQgpbQfoZc+61PJnQU6DR4fCo37YzWxp
il8kqjO1hdMtfsxSBGaXemm6dEkUOddlqZprUhoyVbHvcvsFUn5+1r2SCwdPWnGM
5IWZLasQO5hPmwTdKuEeRm1y/yaZOT35lJC3yWxnjuFnwTxupp7wQCUHnZjXjtha
B3qoqqj/c/utcySu3pV2++xMkokrf1kgsnG6leqQnTrg6DApD4AmKnNOYSIN/af6
6ps/cpDMP1ESBIKZS1bQRImEzNolQhxibxMdrhlyl0vr3vOO3UdEzCGfQFc37Rjp
CmMhW9oZxEFpbq4ImXRiRDZrpKJPcitt+dsC9zXimBEjAtbgRRpsA6UERVftHDS0
ejVPxOdJqz+6lv9IVKkfcJIZ+7RiR+elzDVCmaYxzufOcJcJRRmqRUhUo7aiN+i6
JKdpxiHnSY7AdIRy2/DSB35i2XFwJgrNy8x+fiw6RwVKk89zUA9PLUy+NMjCvubJ
uENrh10ZVa7uMOejCNj/YRx1h1p7VA7E/NzwGpwfhDT/N+0txmQ9OXol3DBrB2vJ
k33MrOX013OOs70IIDS5k53ctG3J9pT6HpZly/XMZakR7GZcU6kMQy6cprcyEmiF
QxG2eixjW6nz+nidki1aoBQJMU9emINo3ltfr1zMb4mUv3s8ncQVtU7H4UxvfWCh
5mPfqMs27eNHwTJFrfa22M430psiAlOw5qcHsavDo+zb2R0bqDku8p9VmR21Ef1G
wmQWvF1K9jxAP0SE9vs4CT9YmYYLUxD2D04DDWggJs5C2C2wMVvKqpBUpGFxu+C9
dLLmbOhFpqFnbhRb8v8ogvLfjAYt0WFh3msF7Wq98jwrxhWLspf3GryRsbhdNhsd
rcNaWsEHviwICJ2oglRUAWtkvUZG4ZempHm7A4VPoydNrS7LWIRBJBdXpcs9Y/h2
FXYPeFy4JTVBviVro7qy1myB0rPiqrMCAEZ4qxOsBDU+Ic2qiuyQQUPf3i+aJiuQ
Zbs77WovZal1JhRaKe+kipZdkED1JELJZpXUw24lJNzEe3OLbpq4U0p1qB3BrU/A
dwVvnj+/KP2vF9uqwmXlV9EYFvr1MnKRj+vO2TEWre7mnc+XkT3G32JEBv3aRaGV
P0DZoyMMuPqE3JUZIWiqaCVLrR5K/Iuq66DrXFZo59aqomu/wczerLf52VS8IpQ1
7gUJACYjfgtC31mVpcU/+r68/3E9BKvgc/jFfS80Itqh3eCAcYq/heEaM1PcT88M
RbPGT9A8+jXp/OmZ38mYyNB0YD9n/NQjOf34UZMk5BU2hd9KxguZ9bR38a9VFffP
u0GkOPhHFm5HSk/364cYs7jT6vYeTW5JVrZagDSn95yR02cwsX8PqtkDbORy0MCu
j2uXbEnkvTStMoyxnnzFzJhgQioisqKPzXMkyJG69tnsJ5K+8b/Mo18uoADTHF/B
tyDMBGWvjmPfAP+KiE6dCvDeuon41/ClNKDfqxy9Uqx0h38A1pfhBboMxpSmkKC9
xu8974o4UxeJT0kthD66AMP3ZFS4W4h2jaBZfjLR5tMbfNZ1FKvPNNDEqsiOuEeR
0dmwLi25lukkQdeXxm1lqZZRLUDPs9045N9R9eP0mhy9WpHAsfnEkveSelzdFQPz
Q1/5lDlPKEnqJVcUhGFQInSXlTbZ6eo16kMYk/ULncy1/z70Oj6ga69DCvPaPgt0
1uyw6iLfVGz5yGf0XKEyMANk24WFwGs5KlfRZOS1q/L1PB1Wbqj3wSeKS2EmAFb3
xPiJdhHxyNnDXZvXRuh0lgtSMzliaYE0Z/gqU3koNrTUKJZYcezfMlJvccM8p3ea
LvLrePUzRqoCqnC5sa4bP1i5R5jBsZ+AvtPr6DVeFQfIiiVcEJYqjycDmmXtqKKl
mil3967wf1HSYbuxJLA3eMPp4PqnQqPjqAilw0FgFbhkzC42WJTQzpxFRHt+s6tc
p46ym3nOE6Aeex7PspEQIxdSxX+kCHPTR5jMeUQTg0t0qyWB0EATsKVjXqbwjwWz
FufGYon8/rFZtg45O68vGbVkCQ/hZVfg7HJSKTDt9pLP8wqnJlWTg/BMoaaTO7QO
uPzKFSt8gC6z3xnVTV7fTzyd0ZgQ6DC9ZWf9Pw4gnkU=
`protect END_PROTECTED
