`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bJChHaaEuP4W6irtKBcwsAqiKWpr+vqcWfe4rXJodlI6fVFDUBbctGeNViJcd5g3
53GhfTvIi+7PTS9ecKCTqXXMx9dP6F3M/xD9mhojCoo98LhpBWGVizZENFNbWv/1
R1Ew40wXj91jc/OByRcQS1hlmBHFWja1Wxe494H/QuTKNBDyDjFrE8SWAw3khEsC
mQOmcPQL73HEN1VR+JnYYvt8MthJe67VSdUX+aY8cxju7BLD20Jm2Al8RyFq60SG
bwovcbAMcIGB3SCFqakaZgBNkimAPdha4GFoRALbPAATtW4t2dTAN5lZYp+Got9K
XqTTz9oSOduZdMovP0P95tZxtYNJsa0AvTiRNIZ9JEkoLxpJZERn1WbN3wxj9LMK
WgpwHUB4bs8uetdmFJn+lXYeAVuROah9JVQnDnNHNBxa1YiI+6O3mIzftDj4fKFS
hQp6fq5zsy/9eIXRGtQBX1sBFZtJEmQWZmQ8Rxo8/LdiPiMof5IALYB1aB7pyqID
75fOxYjVxV0rKcntAKxnkVCTwAG1XzqEGhMeLmw1N4W5Q4zHrVavgmh5g1yr9MdO
kZqTB0NRMsNncbnIzLZSgABHsYr/lLEcorylYrAuO4ES8gA4gihvoL4nabvY1PMQ
yzI1ZfO7xI9fsHWUl6RWTk4aUe2gMNQBbIEak6ZjD0bO6MRRIcXgBivP9Jt695aQ
H/R8hIaQ4CILfbdCvt4EAeKa0JJEjnS+Ahk4jegJWcNBg6jkKGKz9feZBoi+jnk+
xZ+HBxCbiS4sactFh70RG39KOWF04FEvwt8m2lqn9xDLa7XY1qXhq550jdYQDMSc
KXzsXHE3EtEe429flmKOupewz1Q332nYyRL4VqTQhNGrFCRJynQhoJiLH4T/oykF
c+KYXX7cLiEQk6eLkCh+A/lzORVmddNvtblyt8SplF6VcfzeAoGXM3GdZCrMqpo3
9lbRvi43+ChaSngJIhU1RNQVbxcC+lshQ4N2eHFKpTKD3GoLui21t9clmn7gjpQ0
gaigEFJ5bLgu9138GrU1nw9OtZFzyGo6NoueBLqRRkVIH3ubUxnMVoM8vpCbo02G
rRc4sN7nimi+KFY+SNMRGRS42X6QlrbaC22q7dMKeB0Jn0ghuv/I1bBfxYpkN0x0
tgqXSItkVGJhHEgZXiD4RvZ6Kq8uTZ2BnJiuc0qOA5b4d0AekVuPLZ4tD2fxZJUd
+pIk8TjXWNDlvJE9Qts66ScM9xd8dioDqQyg5UV9vVCcpbp73JzGorRMESuniyyP
bLQuHAP8KbTMeYapVH0ynV6jC8bOiwcYGzCbGTaixjOliq/4LKxgHJpt/2PGUexf
TK9F/u8R3UqDdtaT2y1dZnuDxF1r4iMNMhKGDKmKQ6bLx9r+SvTcg/LZoHqojWan
`protect END_PROTECTED
