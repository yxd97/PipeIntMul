`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3PyjJrUMedwbeTSQilrf+BuvuStdhW8G3uf/qWvnZQw/+9hpw/xn87DkcRfM9Kej
JL0XvZ7tepoAmeNRKrmYPys1AX6TEOUkJHhsIOTDpT1Xv4W6wnQ+GNYP6KppXhdZ
nJ0UeDMo9AXiM8asgCP3m+ERPn0mgyWQQ8yR0/SCLewTzJ8jMlqR0KLsvOtje9Zs
Jc0mbB5zSjALumNDXW7vWR0VYlGiUZH5tDpHC9w1zeqHDpQz9G/akS9U63WrmawV
88P/xuz4eufZb8GvGMDn7uozBu34zqq0c2TyndFGQpb/xYg212N6xf5m7xdcRYGg
VD06FDPs+/foJKWhFvol2BrQyProTCygsneQt5mLqFbFrWhElKK2fcQsBUgA1EWm
a52wRR+BqUub3jxaZGoJAA==
`protect END_PROTECTED
