`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZsyhEE607WRVN/B+CbR3Ky1Th+jUzzhfFedBonCkkHZpqzlEuA67YbEvWXv1Imka
wsedl8uJiTh5PJ6q4RoIho4Xx1gijGNVa38zzl5KSknxzvH34Z4axvTYUVUnQLiQ
9KC+C0XHoS6hTn9Lamf8hX3JbNMTYLTdM8WDMKweeh/Y5EnpTOp4Ci6bgXpoESI4
uqZjSEUe4LfMzAPo24l+aV8qVtKXIhorhagp6BD1XH0yFNLNqbQf6sStfxKZTbJC
ifsD6ZXQ0ddAsjUyGqAdLpB/a1K3ya55rRt/drtt1kMQSuEOKQc0txbyx5k0sedx
vCmXmVmlFAy4pFzDJO3SHGznLYusv5mcWpxSjobhFE8OAXjkF4CsPP+PwbdiZ3ZD
Www5wWy+I6fMuCuEc0wz6EaM72xzAaifY0RBNrE0PDUAlA2UdJeyW3USa0tJ65Pp
ku4NEGZx5sQMXZQQi9h33wfCLQNw2ZNFoMr+yrl1Swo=
`protect END_PROTECTED
