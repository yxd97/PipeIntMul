`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tmoTwpYcfCeHBLnuFK6QS2PccVyr4jPJcUZU88pzjhqQKU1PxxVXXndJ2HnSnmN0
Uc8ofGPDJIul0/4ucgRzRM9xsHDveTs6fxewXOLD7dPVvcfCfVuU5N9Xljpvxng+
1sLH1DDuFv9uitvoV/mHfOEMmRGmA+Td6i6nrayWsH+f5l2r2Bv0Zsthlccq5sec
se6+LsPBlSnWOfyJKW4+Y1C/tnbmD4xyk9gJdNvPQ/+YYT4VnOC+fqP7/klsBBiU
QjpbHomZjIkKRQGjVC15zasffBCIDsLFdI3Vq12wdfwlLFP8iX/pzTR8LZZw1TGm
BFA0vh2haILYA7k3EYlP3ADuXOuGxOpAE+TBTWIWxx/39G8+h0o+VFsfUgbGJ0qi
HrAUipJupCIjvV/kSDdMA4Vv/11XKXfwyh46ed8JZT8UN8dDtRVesvNa53bc3TWP
`protect END_PROTECTED
