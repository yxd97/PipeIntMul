`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6Ac4aEf/ic/fLgOkhnzMl8mRiLQL2pi2tIQWxddI2iBbCpG5YUd14HYowYAwBiX
k06sKmpYeXOkNq8avHxfaCpGsYW6mNLq9/+5830wPrQpzjxlY5Jst7XZXgUOJ7p2
P7chwhfK2YzAXNehEOPXsmoLbItlNIitDN975l03M6Q7zrA0p8a5ieAEvqwAZzW5
TZ2kjCrqV3J+a7LnlJZK3G0uS2u9btaYFCxH49Ndprj5DdJNG1a13fdOKwuX8qQx
JohkX843sis5pIHICqhz//a/sbcv4D3iTs4h9/e4RjRpsSnviPpCUKerGzqxaa7a
gEFUWkNFxDDgsS9SPK/0VxXGvWcd7IkJEbZCu3C8kAV4bIJTVpcgyU/kHE+LF6UM
fhoakSj8bqUlsVfdlmwkNjrTIzivUv/6R6DC9695xNXrDlj0HJiFl5LxZ3S70wBN
da/mG1ElInHE+l8lcKpcORt4eJ4jPCy+xm2DJhQ6FY2IDXfFkLJsRBQ1OduAmQMI
Su4JBw61ijQ7DLBJWz+xEeGCAMjc43qrEuIMx52VXRYvADKYo5waHgP50eM5xPkT
YSQuBQfCQd93lARBJL/O8MfD9MlltMuAb9FfBDfuOWsZpD/nGwSvruJRi6VUX0MG
ahhNXFS9Qyiw2rvc/CFh/XQYQt8YBlCH+y6RNcSMpv90/cx6IX3alD1zme6DGs8h
duX4XNc6nDIJ55MqjomYiYYdbNKmBPHB0XeWlHm927fty4nRbG7LdSXoX4aGAUPV
khGWVmlHCVToRGaHCjmAZbxd39WIGL/vYRiOanye9By3KHji2mcY1o2iov565Upl
lpEq5Q214MaBfjgsTOE45R2Vjt9Hq21z7kLlXhEgUx1l3mpKIj/DGn2fR6USyVWa
O046xM+5+gEWIpIir1c3v7UEccy0rWJzdxFIjeG3/i28ybW+gWm6r4iFU2QNQLfO
neDZCQ10vwRQp2Jemudl3TyCvlNP79OI3QCnLjaPSAQPMDLpJKXSqq+2Ki5xUv/9
`protect END_PROTECTED
