`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y79lc1RtPrKJtcsZfbs0CmU5pUNSfCGmFTcuKhuVPo5xHUbSauxeB489sAYVSpt9
wvLbHTXZ3lXuNtF9BBErwFGh0D0t292TnWmC+dIW/rIKJLtSXr7cToccn29yEAHF
y2EMtubTbIqVdrmdRiEwb1Grd/TK4qZ/3K8AaIWNMPhsOQ8yyj29HHIbZzKer8Wd
w12IMQ5I+E+iq49QEzlbaZ7gTLD0teHOjqkVgX3klqynnWq6HEGA0lseZRxA0VN8
9l19ze1p8IG0h3jfF7B4Gui3ZDUdy72/aP+TXocEU8mfp9lQ5s4gQlIXBAplK7ws
MkKHy2j7XKdSl5uebef3YzqAFFi02mdQ7AU9xhO4JjV5i3lPvZCvI9NsVTL+Ti8O
LtIUDQNt9lm0v8h6SSMn0reBHu1k1wbjxNaQA4Wug40sDmogHcAp2geDjGZLmH89
MDQGhN1zjDiBIT+8PkJEjQhxYErKbZnCZK8ZI76PxYsiNsUMfu2z411dkak8p/+m
6XT4zXSmHy7uGnVEmjlIJkDKn9q9ZD2t3Y56M5khnCz4RT7XQh76Bjtu0sE8SU/l
l45p53ft/Ydehng/FtakJTUzc2MLw/6fMZBk7Dbu4sv6aQeJFGLKOCxME4ajhIoT
tqtFgo6ciyf4W9YH2xbvTymUCfwe5BF/PJBXz6AV0oHOtIKPOWhXsVrZvY7wUv27
`protect END_PROTECTED
