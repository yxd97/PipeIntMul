`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nMTlEPs80xpjvPFeqF+tu5UInp9L19/2oTJLklpHJ1RwJe4LquyPq4kB8bs9EYKe
RpU0fNd2ijz7MCAp16cxJrRmOPtkseu7GA6N8nrMJDmt4T8IaKkJpb9FHk1jo2cc
x2zAqJ0AFcH+cPqjVKGOHos45ytv8Vujnl4lExOXy7lGxLyl8VDw9UY7sueZ4Eed
M9X8p6RI9l/CyULc51lo4XRLjQv5F6Dm1HkOKu2rc7PO0QgVR6oCNIcfQm8QkqTq
nGBgnzxrjB1EkfiRrFPxHBuDnnLfqgm9y4YfiMPbaytqGLUqAAwjAIUh37WovXDM
puIWccDkaJDQGJPw0TV6IARbSJxZ+OwVuNQAg/enWAb0MTvW3CKCE3EdIa9aa+SR
cFE6MhnqZ90DFSo+fMc2HvRyRPooebzZSgdHoCqP8y0HzvMBHlvSv9uua3BN+Uyu
BNGDxxyC/th4nzMhwgBDrhOe51JSefVeJZ2C+w/UAPjfJV6/Mxu3CsGDjA9Q6hFy
S7HBMgGcLOJiBFrEaYqHHYANEtQlOk+wnRbG3/Ne+YodwG8Y1C4gRos8D8wcCD0l
YkZcRiBfkom7wgmS/9n2MpxNstTMyHrA35NoQ4u1oGqy1UFBJWMktPzKNXd196QA
STobDJNDANia86brhMoA2B7sDB08kPuOwX8vr8A6GYY=
`protect END_PROTECTED
