`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RUI3geVUSbWpfz1loRP1Oczj01nAMPEpB77Ys1spzkd3yi8YbcWHbKN5MlxQ7nqE
7OEB1Z4XJKd4jruFVGF0o0PFK6ZYryx1psT2+mnFyD9uumbxYt4+zLVIO60/LHFt
yPXpKuGhvhV2RgzyBPlteByV121+8AMbxr4pxd7YcwjJn+2ZvYtKUbCW3GyOjOGi
HwGW3eGlMDDhsSRLimlFRCpSm44km97zIjN7hty7alsepfXmjZ1IBoe8CM2JIp+l
729YqCPCkBRJgT1GjKuhywZwNLMXqPmyIdpDVLSY0dXPvBtoUMQ3EshTZ+AaJRnF
w5FNbuZuayQpjKEsJL7pZSsUutNoX2K9yClWyLmI4Oyen+43YD6wAwjD1QX7XNdY
x/ERwDGQaSIok9dWnE/j2OQOP/xyDWR9ZOUyMRhmtOzBgPGqPIcQYf1FV4mz/o3K
wnXXiT/J4cURshUrur8SPEVrmCWxmeZkx7i5qmOM+2HgdE5KNioKirVvPUI7YYvN
P79lV76WUkw0NjZ4ln1Jdg==
`protect END_PROTECTED
