`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/IHpAyfvo8Vsn9iO/4a+3hAI1V0Zs1gFodCwuW9PRtpNxh5/Y8O8v/pSCPxlprp
Krx3UbhKUqilzgX+O4wtYKyQk5Nl5TNmu4ozbofM0FAJl6dUE1Mrm0Hei4vOKaDg
IL+IEq0Ak2bS0kXyxDwy2YhPvS1qxL5xsxTxFPzUsq6sCBtHG98DfNiXjhy5+acf
eX5fXYsXp5tzEXLGUQP5aYSfWVKFUeE9ML/DOUs9kHyjL0UjO+yWtN2redbtHyrT
oeS7pl+2aYwcWlMc2jFr5B1HfatVeW9+cLsWyB7yPOsAMnQyYk949ratRDQP+g9Y
ZXZFKWjW4VSdpQzOXBZrQYgWJe5JSFSW8F0GsYmutdqBUPVLpPBiHTVjGOcqZo4s
aXtHic8dmmWyWPmgHt6tYg==
`protect END_PROTECTED
