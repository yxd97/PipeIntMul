`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rwrs33Hx4aKjJt2ZceUG/7ShJSlFD7fPYccnuE3oRPJgDeQRZUx4nnAo5tguqD/W
xnzbuCfuhwPef2P++T3nZYBqnHCB+Er53IAv6Qong+YHN6SOy9VWHwAmdb0l6i1b
ikSGm9OPdC3bdk8KacjH5PUYCKw3Xg4EkGFk7yF9lnpr2LFLW1pKmr8P6m/MR4P0
rMqPyTqEaqtx28S1P4X+RTvlq29Ir/cKel9RJ94eoKbSfW06/MJ3QYrzErZQAmKY
SNBBYL8eRut2Ar7PgphtfQ==
`protect END_PROTECTED
