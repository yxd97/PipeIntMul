`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P6XFAeW9PlxhdBQMDmIdZpvCq7g+qvyvrpz+OpbksPuWnSEmYd0XsMZQ+UNbhiLP
xDzjryoDt61J7czre5e0FoCUjYbNoUmRNiGFAw1HQiopuk2EIFSaULBVrwpDtT5H
+ZocxVUjKxvF7a1I55PB+LxhmRjO+Nxlz0PJSEShdlRZAAvtbeCUKe7cTtu1KISa
G5h64ht3dHxjgv+fkCuN6/LTzdXPM5SIfOSLtFX+cxVUCnHnr5hySOM7aQOq8n58
GukLGsoFq/1lf4m1SzDSb6dlZH5qO632k0G1QEzfuTEpACwAd+Rxr9SfeMZvuVSj
UR8K93/LNsgDlWafYzWFa3hfbOkZ419Rj0H6HpEw/GchPw2U/TX3AihtxCYyGa/d
zdHSuikj79/Up0dCkE8JVkhTke87JghzVuUine92tqr5JMobrAD+EM/+kwAR06Ee
fmQ3VUFJa/68N5IZhI/AJw35XIs1C8vtOZaGCqGCeecKsGUKscHSptX5rlhjCuO8
`protect END_PROTECTED
