`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iu+kZVgN9z0PLiFex3TwCOpnqpcufucoEWqToxWPyuyTCKhEjwWnsHQmrPKK9Zua
NSTbTpekuqRRgIRghuPIGI03OG6D7d8acejn9YvCBM6xQmzglfqRvdrU4OxTxTU/
vZkGVNSA+URNfEr5Xid0CCOQ829ugKKGSk9Hbq2uMkRClxiGDAPCq1y4Ldnv3Ew3
Js4tL4/JHTiAHKq3ZN5dc4L+pQ9VqkAEiWhJzjkOAxL4uhRddKFQscl291wdBwnu
HH+XmUF3WBUyI+8llIRKyQ==
`protect END_PROTECTED
