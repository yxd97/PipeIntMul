`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XOiEdgSmCaZ79cugk5N27MolsRhF5a83IgbpfbJ2RB22AUIHsGi9KbrmGgZXElRx
/ZkQhs1h4sULi+Mqq3ZPyW/Qrg9SeoD88CbRfNKsqgJHHePUBK/7xS8ti6FN4R3W
FjXyvOFnLVpszF/YEPIY2G1lHOw7av4zMiXpG6JKNWJCiGHEFTha4dJcmI5T+urS
AGQXP64GgHT8kRWEgmmH7Oq6OUr5CZqc9MyefrnTupPN7i4CXVYyF1JG9F9J9iwb
AUqjGjk4oxmUYqoDf8as0GG0TkFERV/TI5LCo3CZHXcbS7SrVdnaGb6qSq7djABU
NgHnUbDcSfuwgS9usnU8/dnpGnfx6fbGB8Y8C3BbfcXOKa9xFH9Si+qzzfbYmjY0
uwDRjvIjC8fTF0EPezx4CeMPbA22CkLNJnykcB804bzSOVEcHRFT//5puYN+Tdj3
GAxUOYC+jBVt/JR1Ur6/HABMb7TKxq3IAIumo4yXO01uOfeiPnYN5tZZOj2DDzzr
TlGFKdKvVVpULM9Jf1HSB8rAE4m3C7+sxb84GgVCOCI=
`protect END_PROTECTED
