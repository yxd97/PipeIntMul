`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SeOycPRJEnUJXRqv+P2OM1+8Ow9362t0WkTT/eMe2TC0gfHuje9HiEFaQuGDBk3h
wbUor+hIxdhJNF+JIKDS8pnO/6LdKDluM9rXg8VsnOY4vjFC87rTCt4/f7URSjWp
PUwNLL44eE0CpiY3LpLG7rnD9RdgTPQfRllxVoLjciw47uwUyQP+oALRnsDoG+9g
xyTvJi3BRYrt19sF+BNVFY6PTPthCAKQTYqvzjiK08HrHlcztwYm4cgDAkOkAy/t
iiwx09ePxiNsCLkHNQRX10gZltcomDNYKcPe/8kaqUG2w2tyUnJ9D+HBnBPKje/M
tCbczsWfp92T5jboTQ5DuJmwljeB84cgT+zTx0fAj5ks1FZzkCvUaOW8gxLIs4Ym
RhXjMy3NJzpauIxjYoSz1FdBFPHVFL/5NysYyIKLBtxiRjCoT7Zje9waLIJE4DP4
qnU62uGY6for9ixeHrDwnjGnTEfaVxM3uU09UNr3QQa4GJvz2yS9wy1PER2tv/rB
uRPvNVKBcWaQuEZOpJ0Rw3m2d++Cpny39d4EmQkzvdpIBRrQItIpl7vpeg4onQDK
3Gw9viDjWTb1W5xm6LZGhZjtcc4ktVqRPVjvjyObtTdC27IS4bcnj9RkhU1PHtb5
qIl/I7wCSz54OrVEcgoEuB9tmcFOxvVVj5daJi9B7yTBxMGtBRHaFBzuMzPS+V13
tHqciqVI/LuSbmgwGPzEAsdG8UNJYhk+F+E7etuPTfA=
`protect END_PROTECTED
