`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+bb3zlXSZs7p2Yp5zf7fbEi3vT3cbCZv2bsOBWWx+/Zuf7U1FmdoMYhOmrsu02NX
vBsWGtvGZ6V+cKHoAGuyad9t4uyu4Zrf+krh2DggLkB3H6dcux3mEYZgd7fuKhHY
AmXp+CbkNOxGLRMoUG1ZaoF9f5lGZJQOXHrRsRJsVJBMsodN3kD0rV9314zVn0Bb
W4lCLZIQ6q6x6fVHiRleuoNv3uJwSxHMmh1JfHYB1j4SfeANZEnlkefaOyKVXHSJ
lEuLMenaaTJbhuGkZaWu8OYu4fNVvZ2sd76eV1XNyqUbUG8BX1mPGl7fJdQ2+fLD
3gtJ0oaV2/bW6zkjmP6xy2FtVGu2Xgyye2nSatuccW2/LXVCiWoFIsRzE811XTjv
VJ9oX4+FCCipPPAbesQ38zp0ss8FiHjWkP5Wy5vrIWE3E339YFp75wtacmMNZal/
xIKYW+vfxyWDm+Pq5PxGWSF5wvZFtr/mNjon8CLKsdrjPh9xy3XSicaO/OdUJOmB
K9lG9P22gu1RuI1MKxrgqYe/sOlkfo7ApZi5PcDOf1HNPWJFGI3aLLsZHp7JNhcl
aRhQs3UDrhKNvbnspsQFZBOTIT5ljgoVmtrE08vgdmnR5NgNBLYkJ+Aa3ydqLIfn
RwUqhdGNJhZtfP/YCZ6NTvJSnJ9O2VlnS0H2Dx4Y5DSitn6C7EUjZ/jBZVZhuAT+
+usO5F2w9Z/Q/0iqjbc6YA==
`protect END_PROTECTED
