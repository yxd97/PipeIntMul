`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8nr3A2z+ZvKB2x7zzeyydf/pGrDROSiM3bnvsWpyeG+l7O4QteoLT1YqMcZNoLhR
g53OHQHHYMF8uxThAThWuXPNBwpsfPuR11lOVrKAbyvq+lXeLKAw4HoZRiOWU9/V
uIBQ6nccCJJN6mzj+KshYH1KqRAjWCiQX8K5sAr54Nl/l9ZKr3Uopf2wvEafb+C6
Zcpes9474yweCiaHLAYZf0p7eLyxIvAYYwsWXz/oDamZwBzBR+s3X88pOTJFgAHT
l+jgdhE5M6uWm7Cz2Md/LTQyMNuGQuh/0TzvlVU6anvVrMgkOqM8N0VgLsI68i4N
jyPxB8v57KvuXPDeIUbBTcddXjpSiV4Myptr5Qgsd4MgHu9arqhM0lYHr4oZxCoH
+/U7cEHmIVLUXKMBfLqo7TrFWXY4okpY7DJvn+nCPd19vV9MBMrRHtiz86XK8Sux
vEMZHTfWvsn+zZRau/NLR6n6hMSkSsXjQ1LNZr8Iupt/7lzyNc7c9/zhJz1sEfJX
`protect END_PROTECTED
