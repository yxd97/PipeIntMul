`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hh9qG+bq0HiV5LHeZBVX+AhNlJ7nI++w8rmHqCEjWZAl8rmggqJuVpfyCW7Kc5+O
wOCq9ogJ4EjmWBwvybI/8Fb7qjz+rgNyeS9Nyg5zdCUAw7jmKUNA5Ue1Nu9y39f3
YhDt71q/IPe8KkORt2/4UBRM6O6fzvDU0TfjMDe0UcFkjwuWccdCNnzhRtp0BRvo
bMEQwaK4wc9HXDIGkz7Lb42hn9ucl6YHzOC2ezTP+Kd0iFrRj5oMkexFQJh7e1Qq
+8dFsO4pm+jy0XMJxuW2MBec0hL+8YH9gf5vRHHoqgvrZ2y4fOZKggD10RmUQyOW
CNxuvfPFlaeW/Vx7e9IOvg==
`protect END_PROTECTED
