`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsWI4poE2SNAWZXwuJQjHR9l0TQd68F/MLHkZDM9fmWJxK2DfK1aNMFL6Ip131ty
GK/QzEFltdNuciN6qYhwR6dhclLOoP8RaT+1bbc5nLLluFM0Iln+aRMBEVtt0XME
CIDHSQS8b3HDdGCCpQDM1mEvIm4hLDMM7QXqmRdpNaJxHz8r2UQwTPvnDAoW2N0r
d2JuFJQBtmJkq2rc6JfBAdqi5tBMFHkCWvuhKs3V9O3k3YVDugE6ZOQxCGJJmcuH
M6W+vp3AxyoOQ6Borpe8nw==
`protect END_PROTECTED
