`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhlldhP7/7KbhUOOt/R/u6817GUIZHiUqSfrURf00pqPkShjqW4n7IIpwz+WuGNI
TC/itoG5+50mlpbgZuFS8ngA9v8vg5LCUFI/hIQhaNkhHbVi/HHaCLN9LiI09+pm
zyAZTphK+/kqCR+84xhVWtObg9LBWtvUqP1MUQL7EWV63giMdEPDkbzOT9rtizvB
t4Iaeg4iB2kkh7xsOzgXmfPbrIjelxkxTNBsKozlJUQ0BarRrH4jKOl6vM5mqkgX
DNfvR0xpGdYy5r6u7H4aXu2WZHvpPdoRgmshkLtiTBNppdqKvt24SGiTA/Srv8ZB
x/ljeKANPz4qCKKydz/PIYz6DYfge5GsRLKW6/Tpix6DC+yxr85fY7kEKo9RrhMX
NdZHRqGqk95I0kLpw/pJteKX128qgNpHutc+s1ALPZGm8IUy6R779DxSylh55Qx9
dEp+c701HV1eJDzoG/r4WfGxGYMii1DsITRlhlzbYT/il/C+Yh5ejEMHWT8j4kqZ
qx0PgPSg+B3SVND2CH2FzLVyl17L7IFliekQ7aB+W4nXok541y7AIyzIq6ZSrpfs
`protect END_PROTECTED
