`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gujBzSalJ46UTS1PePn2Sp+oAdRrZ4ZFDu9eoRcFrCVTq8ytfheGhOHa4WNnZ6K
8m0+bXpWgD06THn4ArVkyp7f0Dfxe0Wjqnz4G2+wBRHWf6Ov60A1+BniiE2ewpeF
4h4xOccQRYMh0GswMo1gSmrPiCjlnaF0ov4ukGPccDFXT8C/IKaR7BfKAz4rSCL+
SM0kvXCmujCYDz/BgJqR124ypragNK4VCCyzHXJcWJRZFy1jmWzNtiod960kdeaz
WpD0Ta3ugSzJtcPnJ2J7F5RdF5dKuRdWeFl9wUqBXaWnsVBtDfeDufS4Z9bz2QkZ
vz7hmI6Aei/G7z+dZwuzoUmtJYMi74LNN6wOsTOJWlRKGrNB1c1yQuVeo/NHZIz/
mdXd/yP69fP3MyadGOnRzinBghmlcQc8/MKKyxmmrOZVD2ctsX3F+zNljY0P+f/1
3RHI1byvR5GGxd3Ku2siUrcWq3Gs7ke77F/zGg6SfHNv5/wcbzYADWVhp/fbKsfO
wNVtNOTCv6q9e9CF6gPrT1q7SaJH2lm2yCR65TiJFce4p5mel+Tk6bUW0vKVBrkL
IMjmN8HSh4A2IJpXHo9v0A==
`protect END_PROTECTED
