`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HijE4ae3UnKkqvoP3kwVopCoYSOkGqSOypcwEgguCU2Unxg+7tQFXR0QwfhxTASL
0xd6ClhzLENHyqCdpNXXIfrqjdu5ZLXivDZbcFvyxT1cuFhtGUKcEohExdMUej+I
TE9NdY0DwB1l6ux52EDeHOQmxmvSUutUCzzs5KkSODODe9Otpb//dKvaT/uk/Sdd
/JJp7AyqojP3u3XBWuhF/3rE/yyBsRncIZ61fbV3nusxXAZkoMUUzlhon8UTzltg
uNsaAAZ2qvz1dpRMKqur1xy/y+EVyJE8jITuXFfmF66rdOApPEEcjOjD6dz//VSK
fTFJqynWrI0OFDCIUkGTRHSf/Lqcc7G7g2L8IgtaJr8Ui/z3FMPthqp5wvoHSeWC
F55Lo6A1qX4rUr3pGQpQJafHg3ju7Hs7bQIoKyKRzceeydzNbF45TE2chuiGrv/W
7Q9AFQMtXUaIP01cWGvy3olV38704YggnW6OzMyXJPE=
`protect END_PROTECTED
