`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5RELuqEVKoNA6LM51C2BJjuKQBsR5AVLsdSN/kNHA0ChZ5hvF/Qdz1bMBEqAmFlb
pAjW4JWvgk6j1qFgwGOVOxENRCJ3Gei7T7xVgSOy3WbXMjPN+vPwOGeOtJadITNE
z6F/40vQVpbvP1dsgVgdVR9fwPZCEDZwd3RGoUB9Ru2SDvf7B79qR6ydcSFciIhl
4ao6rHNkaLVt8FNKyKFewc0EALH9bnaMgb7dNGFuebj3TZ/PzbJ6TzZZidPCiU15
+mZTL2wPLvDjyObFUA663FnNQTovmeoQ90Pj2zFX6wgBHmw6GgfNWJPuIktbIoao
JOvF2wqxjDIPyYQUeJocLonnWwUEl+VVqp07YfZeLezjSq0bHHoyIRBk9hFt/ycA
Ah5npuy4C1Qs0c5l3d3aTvXNr2Lub6xRMHXH3w39gB1Ht2PUoTMPCXf0uWER3ts+
r6aUjSr2alwYuhloss2rCxHVQaeC9tCejg17pGpE/SggFZgvGrpZJtf6Q8iukVp5
54hH+DixhQJVnYuBb5rMmqKTGdxJufIwYjAXnN+LUqI9gEqNiOL8IX0BNW8h02EL
2uJt6UZTnZpm7bqltF7wHyKnlu2/4nyY9SKU5ZDxY/Nc/f3QbnQGrINkK5hhVMzr
oAWcw/8wTR3e/oPGi7XSXeWXSZtE+TjgcE6G5Xt8pzA56LVM4tDYLu+ufojpoPEO
7SB084l5gnOPiztFKkCYTxDlDVrO+F0KN2viuohseiaLUqBgwxY6noqqjZeJSa3Q
A997GRqHFbjppiiRX4N5osrTz5tww90sK4NDIo3C6Zdja/WoDcZFxB4kKO/nXDkL
iGzaXYEs7Wa7eq6mSQC9Y3EVf4Kz6uq+1wZPepgb3WwX2bsWUbN+FDL+mzagRERW
n6+H3ndZ608Drn8QA7IMAjsp+t7NyUKNaCv8iQznOaJG/X89e5F1Kinjdb4QqWCb
1NseW3vZ9ynegUK+gM35WDi56XREW8KDsRojE1/HAqXRoEqbwvekjzuWUxoJptEA
DtazRH9K6+Sr6zjV3lLkoua0z6AE6IVzAJYkPYw8SrTC6sdtK4MyJV167GhoMxvX
pLwxNUxt8UjcGKc3rCf1Tf5eRhY/fJDgcW3fadkHjFP6iQLHNPMqi3vMTGDIYe87
Q43Njvt2m7KOh4HX256LD4r6BYl33tL6oIJbpWXclijI9y+x9FZz1LXMreixeFXZ
7AORtV583LeEaALvrEpWj2qQ7fCqTzD9Xk+ZeJ3Z7aCN8WVAy43HYJwTldtsFkw6
dmTPuKVaR4HJhrTM/sVAddj6iMg5qV2ULAapZ7GWOSm7OCfwzEFQKh2vdaaPFRr+
o9WRHpkEVRWx0g14u9rMWQcSf+BFW2MwDrfxd3xB9UzHQLMh6rVqUyK18cJdV6BG
GZoHNsIgUr5NTmTC5I8QzRuXlJRzoGBgEmS4B4wwCdsrIMImZhvw5oTPLzA04REe
bpOqI4ecUCiQSRJ9jgket31j2RUmn8tw+O0U6tC8AsetHnaXuYpO6qVY+l7VxHPx
1tDLsGnjF1T8//uWohO3myRf9sqHOpxgSZslJeOUrK6JgUV7ODWu9wyhvciL4lT2
jeuDD9oo/LOBrK9t4NYB7T14GZongAo5vtXmtdYEEmmrWUhQnMHQETZIReWXoAuk
s/yeIK4UPdTcCDH4Q58k6BkvQc+WhetyV0+AdBQsRL0zj3q7TfJIqteBnw24iY7q
g0RjYmFZ8egxjz9ecvEy4FY5KZHLZpZWNKWFojzrMUpSxavqjFvp+fsBgmwEN0ol
k3pkAfsahquXaQzbPNJe/fvXGjHwJUZdXywjPwZtCY6qZLttRKkSvwCngrWCGRAj
+UPTOn/1UNesrCmtBgGF8WPTm5W+jVAhCiCP1ak6xVY5V8CmG6BTFOJwvnpDxq4e
50IJywcfyFhqhh/tn+z2Sgwvn14F1dHaQFUOgGnjzlIm1ittT4zEIm2GtpgkU5Wa
GneuK6NOeEijrbSRxQV56eicdhB0x5DDXYSo5vrUa/0gzCoei0qM5GgyQnCQWRtk
MLtYzr08XFwzIQ1Qcom9v10Gx3n+u/kAwUVERN/gAFCy1VMhW78fDbY4l6RUvvQv
bsVULZ6l7SxVbN87L0u7vlLm3Y0qu3IqpsEzJcG2OZ8IgjRVqSnwqJILl3QSrbqq
5kQmg2W9xv9n1ZdIY0w7EwZ08C62LYnaPg28wzFD5CJwZPR13AQ1M2tnjyUSY6n0
0yo2Y7oSr7c6nb2UabheXI/q954UNaYyO4En/WKctAGbegIK/O+q8TThl0cQyJNk
LZp7+1GKtUXVMIA7q5YDpVaw8b3qHf8HTX49srZ1R22M+NT7tlF0E4IeteENk0QM
YtM4Kn+djcOUHPTxb4umKLm0ABPNV5mZUYy9qYugPe+jQBBld6Fva2iPJiBLno3O
kslC/bN0fpQB88lvIvWSkv4LtdBe6vvtZ9IfgsbkY5BEMgQoB617vcd2g4ZSjLsB
bqTtIU2Oe9Lydiy5ibKZ7TGSkWKucMAsTxL38ZrFgojYoEyeBuauHAqz+SikPrqG
KVKRtulVldjsLBkeKtBt3Sfa6pc3KqanU2xzhk8EyQtwAb9BJlmgj2rbi/OIvzZe
XqlkR65yNI5CidJBcRCrDhFZSpWkYoV9EjxCKjmsTb8Y7wQLNxH+x/WDMWgVOdFP
r/ptJ4emDaZL3tC8P77lVY6AeYRsfrsqzHhbAP9Qkdeb63wnkF0lmQOsnyla8Y7z
qNeq3x735yHjMO0jHcSybgo4cTIcpSqeJtoGm4ce9661i9DiLiP0Zh0zpRnK9Etk
Nnf1fqfjDV5pVgZV05cKMeJ/xyNouDE/OUs85km/xXwGZfrd/+IakvE/2LKQ2J4y
Z0X8PpzKDFe6LXvgNSvlKNJVQIXMwfjfkTY1L8nulf8C2x5vBfMaBcmq6AHv5FmP
Y04hfG6o2EaZNE4VPuDg4gdFCiLO5HwP1NuFLcHMwoCj64s/dLzkzj9Y0OJJW8LQ
RZE2Nu2S7eDrGYY5OpOZBeantfxGu1dpQiBfF5mSMbC9cuMCSLjgib+KFgpW1cEc
W0DiOiDYwxHzwbhSH9COFCnO0GPVPOwCrwllwIYh9lxOxkRcs/4FE4gH2bV5lOfI
cUuutsWQSA0A5XnPQ4tlnL87hs4em2jEWAKjbhIHoZGbiN7kBvOYqv4bK8kzk9Ar
rXptalcCwvn2ewI91ppFPLcdAVH9lehJcxfeU6Vf+U7PXAwUBzgmOGuwnusvoxyT
bHXvRSY+uWPs67E8cwFzOsMEYYcD+H7L7wx0mrLrePLYTdBW9O5GyYqiwYSqfT3J
`protect END_PROTECTED
