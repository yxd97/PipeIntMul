`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ry7OiVbLTerRjJ1Cvw5JNzSYQ4S2lBNn+crtUQnYh6hyO6VY4QyfbYLbTuInHKNh
i+HIwtxJ9Js9B1CsuGndGwDOHEOWtfNNL4IPCDlDzs3gNPZfsyVr+NvfA1JDZFhd
pE0rFfm8Dcw9QYPBU35LOLyRQA0xlqmam1CC42UrM0+RJz09WkQcsZ7bVgAxXUFU
qIJTXeEGzdHcfdbN3VXuXa6hV6IBy84QEFK7+X6rqYjdnOJ24UNqynIwkxy5OeeB
`protect END_PROTECTED
