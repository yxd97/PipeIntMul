`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3BTgZ7RrT/4Zijz5UWcSW7tXUgPzAGsIwpSC/MCeItQgAswZiqWeIuasjlhxe/WJ
FXZVGTHdrVD65NJ2AdNfX27c6lupDF4OepJCaIpqTpfETvEdMkBcoCnUqZU6Q/Ht
aRkpTBEiClcSDosziCTxQWx2aL3E8H24s8TX8yIFA8pzIUDdWhGDocpXjTSLf+ab
9CVf+5zQy/jWtYl4ezNU0vT0TNT0uUJ4YG24k9BRvynEfAoXKj2tkkwQIwkZ3jAz
YQzMRH69Y3aim8HUzqAQ36xKcR6dC3j+o4frhDYPytmzfl9s7+Sg5I/4RD4JEJ5a
GpJJbCnBSez+Cxpk+xjR5AAeSO0fuJveuonQxUkg9TPaJKkWyB/7qTjhg9Vjny7m
6JKxGYuj+qTWrmj6o1AetSW2exyQlJYPL1wQaZSrjACTOZNhjFOgkN5KPo7q1mU/
R1bUuoxs8cSpqwPEIXUisvjnlfBtOuZQ7Qtgpl6ICRdnFfFAQDAS3EqshgysnfLL
qq0rDssmkvMN4tniGT5/6gFHdBb82RSgXV9Bx9W6uarDbOQPJkdcJgMD6vXRgCJT
7FoeZO5Up+LCKqNU6KW4NGfwRJUPCJsCodsPCiqBz6KJ2NAyTPWjqoJ1f7drpr3i
B5C4HV/O4zqYU+iqRRJb1Un3rQk39o9mdA8BBRbG+QmtYln1vFJbxirih5ky6nNr
836V6hKrchB2usBHDldlULAgqHsiJ4knizGWSm1z8nC6CBTMTSPg0FW+9OwX3gi7
hv12TNBhsLiDsUYc7x+hgI3mD/JGbZuXhoqfTkmNuhvffQkeS/ajurPHgCp7EJAL
a7SxvY/UbbEw/jIlH8a5QYueovk3KLGEgPLeNrCQpNs/Ef//IdxCKFdCdSQdkowG
RR0glRFXGsdo5QOlCqGAMsDgKnyB5Yn/ch/va3NY4Ge2mfLTiiLoORAjTH0CsMtJ
wyZivuoHN/9zaCZ0nCihURAjRmjSYuMxnnlX+r5RJEnHIZjjFW6tgV8Zbr+mJ4Pr
y0LfGf7+GhJBSO4GH8zQJmxZ3ai3t8b3g2E0KSycKltGC9acSWVAFS5IT2Bdv7D7
TtwhDGk9WYo8/dL94I4LQ/lon4Lu01zxWsgmOK2KE6nNE/BBhVHDhW1lFTYC2qEX
FGrbaMjI0wkO2NNbPDy1Xu7HEAEJEnaG1RD0iX8kzbt5xmPA1hIZJYuytnibsUzd
FgumvLr1h/M2qukwj162MAWG0REllvEUKZYUfL2nGTox7Kd9eZw5TlHW+N0P5G0f
1HrRdxYdMIOapELHS9WIQNXGBC3El2M9P7ZnObLiAyHsyxUlbSGVT0cjxred7plI
S3uLI+iqcf9Ky8fhDqNqXYK8tPM6d9+ZWfGCEFdisTeVXkzG+mkrjR/BJ0BaOZTX
b/YBIw17i0OF1qqm+azQfjODK5zSmlxsuYcs9wcFJILkBkqeHPxjGQ2TI+rf3BdV
LmtLbd6ENK70+cxSLTNLeh+XgpsFKM0mNnjNCi/TtxnWW1OBHVHF5D5r4uL7VPMJ
dq4/kKMVVlNvl8W2MZ8Qgg5zSi/1VjfGl5E8CJWoTek6VquzyxEcXblFl+nbqsfH
kXNsFHryApBbnJ0wIn7O1/eF8jbJ6savhp7YOYca7W1T5ZYaX6i6BqX4SvbIlTXD
sMpUwqpRExuOesRwkp3z/8x57rmUKyaTZgOFN/VCPLx3E8YYXPI8qQT+/acrHC9V
qyzJb04lnJufCDyqOGZTecxDDVVYC/+wRUlj4x8YlDPDqHBhCsmTCtZjI/STYilr
/K/tr82NcaNI9Uxnr9DD4lKMOeL20IoIlgD1IwXftpuxbHaGEj8FLoB7q9ekOaiX
X/5Nf2bA0ai6crga3LXfLcBI1W9CRGEbstjYhtZSXIb5TFHWsMxS7MzqkTM8j+S/
yEhkUEx7dN26Lg0ChE9CgziqtfUyRpN5QZX1e8n1TU/3tdlMnVQJKAHDQx/j9Bg6
5H8z3zg8S1bmy4Xtiqbt3MVraOHSj7ZPDjIEbZdHUuzk41FvEWr7Qw+ah0inihm6
84zKaRuOZU/kE1vf4gRlGgBp2jiD6F0Lcm+EibLxvHj/i9eMdhGyhqVYh/fhQj9g
Ni0vPmLqTDKYfJt0mS1uFWUvLrRqQLTtPyhib5SBRXPPpcam0QdcWlmvdy6p1Q0Q
q/wwwcs5ykmfEoT2F4IgDGbwhDMfrz1XbEQm/f7pSORXjiSmrIj+wM0N27KgkHYU
JkVp2DSirM9tblKlFLVip38Z9XiVKvfcYGYBVEUMejRvhxOHvEmUBCzakstn2HCK
69/VrdI9JOE1sGWTku/oPB0XldrmKOmFUkM2603Oi2whkz8rOMp0TD2oK9M7IWsm
6defy3L98SU6PzZ2zXWrzHbKxgSb8gTL6IeL/P4+jXt9R3QjcW+p8yCoUpzTizN9
2iZBiAwqBPP4frn9Ff63bTDYRPajUV/RL+Sneq6Ja4zoCnWBLg6HdfTVj8yenfOf
CBTYV+U3fLaQkgDnaj4UwDr/kNpOAOndWxGKJdN3W08ySoz9QqvxwCU12Hv53az7
HL2OpMl9beUCrHz2N259GA5LBsNL+lZ6JT+Jf3f8FLcstiJtA99XRrH/Q51m5h80
WRLoz8hWBQI/aX+ftH7/ZrEfQRoj0HYoT2EntmwDmX01KKD8RfEAwwdRynQLelEi
ZvEU6Yf86FIop5WollHsZg==
`protect END_PROTECTED
