`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVHvZ8E2gXWc2Yv7Ql40C9N0B961mHU7mVor7YdrOYp/u3Oa9CXZVVVRPX67biTh
yLzoIMGT37OA7V82b36eTmeA/GcxxX/MdU3W/hH1S+KorukcRSDSfYva4eCanXQI
UlNxK7bAFA8VJ2RMkPtO9FKPaLxCPCzIs29aLhWbi5UQcqnHQA/uYxy9vnJ/Sew4
Wx4XshHuKMjmWLNqv1PC0IinV5PmFlQE6bQ4lYndoFazeIM6+DXEuKjMYcZJC+Mk
omNHJ4zZda0z0OsT+tm0+M3s4iaa3BgkfKURfZh5L7WvHoYiqs1vYqd+yi1ddLNN
zb7Uo89ih1uiKn2P4KI/bHkNzm7fLnSTzMkzQv/J13wotXSq1bSy/l2orAqZLgAY
xnatR4jPAPcOkm0oXmfStvRQWMDQFuIhgg5bSI3Jif8cT5CM49r9q7Pz7Qri1/Sp
ZE9qpqRHgMqKlLCN38fgDS4BvF0pyCpWvpwqhU7z6+6jF7VX1gAKxMKCPw8gXvc8
yW7OPnhpSSGFetJZavaAKh+emrIwEZtIU6znSStVAr0=
`protect END_PROTECTED
