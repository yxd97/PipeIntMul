`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ec/gEgJdZjMNXcY4kRiV+S0GsaIyTxYKyy2V9w6PYwJY/GlxElrfMD58X3CqVI5s
SeS8+62XO077+pcx7q7HTxluEsocT9/o+cvZCkppKoabjCDap/sgbK9mdMDh0O/L
XieNbWKOG2lA3MkVtlxxIOlqUzQF0EqYA4ANSOlNwq8QxfwXrd6G95WJ3NuTybeF
TEAUfpnGZUvpDsbZ/TdXBBrZKaXj6qUddeNYajycs6A+RlBiBoDttZ/4A/G3i9oB
zIib6nynKZBhovD1NZFb3JpMnKpEr+5TEsbLIbgGM/OFE5rv/XizHxWXIAfqAf8C
fCvEQRwiciSfYjnPh6f8SOA/Bi6FGz7Tn7aruLwjEbJE0qL1xAqS+zUywkqmUI12
z8kYHhGnp/e+40LAhSGixsFmcasJ4hFZvrsBDCbMxrrJS/UQIX+asaTfplqhkLaL
CZD1b5JrvaztebAHtbmSSsJJAYs552GI3Yrs6gtBIkPI3hKdilc8pgBXmAl8w/lq
vyTqwCPzxI+N1yFsuPNfUwM6xAvRZIcQhgGOQC2wey4PkYL3fqEbMNTg1P2XZLhW
WeDzAX5H7B1z+yoEmNn43lru5gZ8+rH0CxW/BDyjsPtTOl8bTiNKliBhwwDkUrsz
SeA/4r6Xi/kfwcuo6vhOEnJUzK1MJ3Yb1m35kEMcSCoxW9DDbFy+oleCwcFEBUUQ
yNNeaHHIuLarMJXZ26z1tvCwcX3cJsoFbGw6ux07e/4hKsLJPP1fQOF0y7MfEJ0z
P/kVXZBvvRNQX4Xar/qoGouBhAcIneXbgbg7QyevxpQ04jvjoEnV5hTPPfLuNANv
biiCJhWl/7DGxH0YwhLEWmPyShq48XXU7rnvVe6Mf5M07JFP7+s1HNw17HNTFAFq
VwUHLNuoq3o+MTMGDMLrsD9Wqi7cmnsls32vMZ6THJZ6GXctJt0RhYhr/koIWg0P
tDFLGuuS8+UtNUOnpAHLdy3AIirs8gDpcVJ+jMEYktW0cyvc3BDjMpGo/jnYifYy
cvruJ5U64OQulSdx2lhs5pV5/wtRhVBlI6Ibe+yjj+rZlFtZxfCJiw43gmMvPoTu
yn6OuiMvDpIWarUJcWgKsVUTQa6mkBEiJ+YvVxJsRSLWHuRtxxCraOnDBsXgHi1a
9aabcnH50pqsPC8Tc6Z33oCKCeTROZauL7rg87k8vh/LATerKs4fzcOuNUsa9uwt
1K/uPvmYb8en45pZSdc6prnwXrxbjYfHKYjI77vjyDBLVZ91Lx+MgwL0e0Fc0Zr4
hpBoLiNUQtYfZF37pWTXjl9q6/2BeKSlkOw8rZcpx4nzHDoDgmi/hsOTZr3WzdhC
dVnAEbxrbG4JSlEmxcUZ/ZAEA/tikViQ8AmU+tU71Q8lfiXc2XM9UNa9eyafo/Lq
aVPDVkW+F5RZ+xo+Su37u2+1yL28Q+q5fmRKBtDXp1poqzGGgnzb7BAtV/TlbIRv
8bjNznsSKpoLrI2/HwW/DCOW05Z608n/7ZLQWrWqxGkAs6UlxAiXYp0igMNDZjDs
Dff+ROskl6WOKgUVH60jvUpbIghFXZvTONtQyIwMyzNdLtyMENv5fFqsvPG5+nOT
ISpTKmDe2D4RnAVy6pc4/Tn1zTEzZIIKCvZdQmBwXZWrDrT3nPkyERijHqLk4CGY
tRlYlFCyjxZiKp+zL5M3e/GoPGHnfJQcwgY/UBqS/A1DbmdzqNXb7xZ5gf2r3DQI
plVJU3o38FhygFvQz7IUvNgRR+bexSO+3gTZ+zFxy87rHNPjH1Rzfv7z+mxPa2e/
zlRa371vhmc8x1p3HgF1TryVCB4vzf0dDMJHw3oUgOJWCDxafJigSVTj+h5Flo2Y
U6p7NF0OHTjtFfqc5tzyROpYdd41B+05IIOZf2Wg79Pg9o5D6CAVm4YSqziVlzr/
NTTpHm3bs+8MXHMfvUMUc7nK7FH6RdRM2Dg+odSVMVx0VksyQbGbJgQrVQ49zHYF
8v08B+5/IhQEF5H/M/iB5I8v8OVEgE0yiFOni+/3BoPqcIaT9lkZ7itN0gVQxRCu
nKYkUzcFL4ogShD+1lAQGBP+lEOt9FwHCGJRRPoyW9C3GXVM08jkO3U1aHkbuT37
SysUv7DVEiH3BhUjw7BcD07usuvY04G5AIEH/zevXKwZWQJDWUXsO3CFLBGpDBa7
LYwuHDMHIx0SAh598c2Zn7nwS6V9kfUOOBdGKXKtljJtlg8bTIm0Ofy7lMwOfUPV
ZHmiUCtbNvje2Y5BYvEJRKfKHP4GibPACXZFu298rFgkXdQF2i3LvtxHYoYEH312
OJ4gkBwmfFOfAHr2+BvuOghI2zmFTv4pASTh9ZqRYQTW+jt7CqtMM4SR/7pfeMzi
3cCH3M0PV9C4pzcBTYSAfCg00squXvry4YQ2pTAwhkvJjWSWUYHSHNBnELBVuYQX
seTKDSedO+50zoTFuExohKLtoDLaphRkqnKXTD8QzNGdFGmFasIkkP/RTg0bCH3P
F+mhChJKaEiIvX2aIRj9frcFq7LhhFFSQ8pIxyXHa6sZ46UcMwpM5LyZ4iP8zqvq
vy5z+KRnSV4vhJn9LBudvCFonkB4Y5Pgv2JsSd/Pq1/5FK4i/wGaiEFx2UiXIkaN
LVVjH2ds0uhLLnf2SglXrREmyAh0K+C6K6+mIkJJlSlmns3EfW03nlXtxwtp8Yfo
UfR344AUEtkRg1AQkY0bXAsewzQqwyGKVTy6jJwIKiNLAd+gfwpfk8ilBhsrfM1o
GpooQLiZPgyZ2qaZrKxYIgG/EGAotIEazYRSXMlsHNoA9xVzwe7zO7a/+RhBgFlN
pxA6fyxuDWwpJftewTI6Y+a8xg7vV6pTd4rBrJafdlwmgEfjP8dP6IQEJAWibd9M
W28Cyv3+8cktsGf3rxGibx6bI9yNP4LBrIEYK7Ne1exyxviCKr2XJmWdm+a4xLDD
2BZqVgrP9Ni6ZbqXYCQp+JRH/dfyk1WK+OdtB/eviERNnjbNyarkFNkbBns5CXNH
HAdEms8l8SRsdyvUYLeM0+ZDh/LMkRldKMBf3sRSpBwFnnDkhZ3LOP/xdf9py0eN
981V3GlmwobbGrThXSZ4bWk4YmDiqisxoiiM3BAZL+SThv8KZWGjB9r3FCEIQhrt
rrmK8dtPFmaoxMBhKxFj+L7Xcfi+fYaAwH2t2fs8MGjA4OC68kRBJDtiusInk9Fb
fHUMQqXOOLUnR/PZSEfPxLSFChPp8SNbwrGa0NWOZgXGZWBq/fqPcJX+JRZKtbU/
Gkfv1KA35PcN3/JpIjW+dOnBzk6YsysFbmiL5qqsPALJDElVfYlzCTmM38BRP2Uo
VwYTOp8GprhNbs5Ns1uHVx6DqB55TBAdxocv7jgv81J52ncXjrJ3hBlEa/lkUJyk
6H7X2gLxQ9niKblLkhSHm5T0Flt5p/ERCypgGrOp5KbNUlUvEQIPpm3fjg+TYAcm
z5M7OYAzCtR2Lv/izz2cKsjCcfM68OUcXfLBZR+ER66MsIzoXdQcnCEFGbaRoZ8S
+FuUWq8AYt2DOiZmaBjs0ubg0eYq4bN4iut4mTnh9Ivb/LF7P2AWgb+gUCaevsWU
SGTtv2AXHuACka6kOoIJ/6siX/PlTOZsGV12Kk86E9q7VyZGGBYQg9e5xLp/whNS
dDnQtIFyiOm03Oi0MXdQv2i94Mc6myxEO9nl+xj8o9X1zmPtAurUGU0vfcm1lkXj
DjFjX0Zj6cu/gTdtPUSmxbsPBh+vmULSmLkLWm1ZerISamXdYm++XZHkP184AEe3
sFlTmlL8PQS7t5seqSNR9tpGR0gtz8KN3ZwuMbcBRG1AElK6qA5SX9KYMLL4PuoO
aRUGfqE5wKpBGBuzNeRdPbRIv2yrUAh3dB5T1qzyG4z+lg2pgxE12fVaE6s3YQrO
Iqm7GWsQ+6X4YZhC3jUKMWHbXbGV99ihPb+NGlvPC8jhyg6bidD/XYSOnfr5xySF
NabcXf1NHgfDY2G+SVSjFIk72A4IGJZ1YPhWETr5HYEeFW4mRO73dIosHF+BKrXg
zYwdlz5xAERCA8dJBLH1BAhpVb1oAFhbBiXgUQnq9h8QUTeT9cISIAI1KNkTV/I+
JXykanB+HMuTE4VgFw5sTF1sLIVR9tZPue++CCm2tynkuBUXJPe2xVvY1+Y/Wuvi
8cSgwuC2bc87xHSdDxLfcDWhWor00Gqtcm4yzWfn75zue2ffzEEPbfP+bWXeUQi4
NrazI+SkAnrRglaMTN6XHjUUjxqaw4BGyXu/VyvWQhoaotCk//f7S++E6gBbG5Kx
Pv7Nz3eS/XMqlsnvgNCnBU/+BrTYPB4nJsmOPVadeyp2CXw1GVInC34eJYPJI9Vn
U4WPaQeqHVjLpFBzjBCbKUjCh5YjjoG5MjDMFhp/OSUFTt2sFBI77CtURaRQ3U7+
nN0lBlNH18N6Y3H5Ka9nHtLnpi2wJcLjkRMPJ5tAk/Hpf5e1Z7WRNkNzr4lBaYAj
YQ6pmMMPeHKH/Gz7zIdAb8bcQOuzQFwqaeMG3dGlmUFVFqb+WP8m5wfHCVeFsvGG
xzdOn/S6Zc1bV2anpSO8yHpRbFncfmMJa+VTGZ5lNy6RafrKKVezoeCLjfEmKl0V
211GxZPSPfpA1MVXW9prip/fxq8t8BycvioX/qxRDimTbZoOQkDsB9HTRGqMSxOF
9k1mV+bhxAOb6UJfBaJQ82YXJElqnleFJ+OuJ5fje0Hjn7KCqPV1Jd2qCZbs6nTP
u5KYZ0hkWq8lHmsb7CCLQ5adPYUEXxVjlJnMPEXI8qpbhr7cjEYPFkqku6nsOWMz
6OT/2lvKh4VPK7UarlOQ6jUDUkhbQCYqjZtBvnerFcA8z3h2uhuj7q3QTIxgHIqy
01jAMf/4BK3U/nsBmgEO3fyB66xHs6J+wV8+JEI2H0xTuGkhQN8ZYi5LRKEQ64Dq
JNc7pTFjjPgpY9O1gECzp+lxxuGDIRU4fy/wwEVqo+qv+DixGvgZ7hGpFeOYlzq7
bES3anVEbOFtq7QPOVDooreqNZ6TDYJfGeB1LD0UhDXN108orK0RHa3GWw06WN8U
ThU3D1B6YxWdOIUN7aRs0Z3fOB969dgEl7wFiEYCWG33TfG8ZvLSc354Sx9TwzWB
ffvY44TglwMomGMRFrYdmSgv+RrY+wBoW65vW8hJVjHvWqg/ve9R3CLQ7mNTzeBg
gEOdjxmp+XG4Ma0M1ksrVtZreFTU+QF+opxvHX/a5bE2FQuBNlM8enRpUSFs+uVx
4z9lc6FPKK/P8xNCUH9EH/OCenln6N9RL+mhQ9pOg8iC3tpzqL8V6WU0FMQbjOkm
Ae39/rmh2yY6qx2zaIPGAr1OCr/hz5Ayu7S3LfFb6JIMgVrd+fIJQPEuvbwRExHk
5b4Gfe8w8lNxssxS8sRsj3yTioXP/WgJv6hPzkg5bx6aTmkpyo2y3+J0VaE1GMN8
sdImyCpYqJ8tWxD3ZlRVJCh+a5bb/iV9KxeKT1VoTwDfFWRbyL+3oaxVpCEUMQLK
ph85eQdRzf729CqUVS6rsXibHwlt3TNJKOQBSoBM2ZQwILIipak9SCnAMgsO2Fdu
9Ilgt8evepp5ucLcr8c8ZyC8z0MrYQfwoHHN1qQFBhLYhvcFwSkl/hl1BAEpQ4F6
aAox4SzkYebQXrEIqSPemRW+FrKRxdPRV69W/DT7ystF/tsxZqc3MLX9RxTPtAO9
KHvc1YzvSExUazSISXWwrk5PK1U223FRmRL437u7Gh10e01J0oByELCoP4JwUqaW
g6ouhAAxRcdQMnSqf36+YawM557fs2Nl1FG8bdxmz+zog4wbWoyRaKmK+6RFrWFC
wBwvj3/j3xQRdYVEha8ohkDrYJ51V4txUzndvPF55QxhNcdoq0f1IUWaxGkwcKA2
8RfnRja//6LU1SP2hRNONsKCQ5jY9KrFXd8qwYj3TJ47IKTHXPGUIU+gdpJ9jmgc
QO/a4Pzj8vOV0fRW8Yu0Wfn5sQoiBdOQzIDmqTHDTdG9fRdTVc6U/d27/y/AoZPP
leAP+6Mv2He6ZtCufh9ehCc4UZLrV/3oh5vRygjjP7vTJHvKzFZDimxzOSknuYhG
QG/yPP1K8RYU04ztOMP/eAd4RopLOuCU0zansOr2JggpI9VUWT32TKrHPRMzwNjd
YR4MTgKIS0amgt1AsrmAqby7IXPBf2R1dMFLjsu3FaxM4veTW1gHvYI0JBa/RDbX
5xLxwf0E8srNajrhal6bwr3lo/csbMw6QZHh2opwrpTCJvhSGmVTv4bSY7F0cC7v
urVxTm5FinQgzOAVvLRxhYrmZrm+0uvXVHEMlnzPcHLsnzxaZ0QbbNU5U9WLJG44
RB07Lcl1VseibC3p53HV3eE3DHFQRzZ4g09gpvYmPoY4ZtUQUhx3qRtHGDOL4pze
Ny9G/veMefmL06IavNkaHFkBQZt2+g0N3ePfkvXHdiCHrdvIOpO547WvAjSJblKj
hqdbtNd1bevNbf7APKAl/OYH8NXO9f+nTLFlFezB2faenwRnv7QRlXfSHb9QX0Av
rXcyr73XLqT34ZX8lxviZsq2dfiKheR2R7bRuToomuPVvpw1tfj5L8vXfLp6piHs
vG6BX8+lQat/Vn4Sb3evp8dozNWDOCNn5ozsbTgmZtuPfVsU1mskOlhP1rXUe1Fk
AyIboXpNxp4l9YZqyVf44wp10kTiDGd4JV+adYLSKfh7/VplE/lghuQ95eJ81Cg1
ndvTqCI2qAWrsaGq2V6AM3tsgpVPRL2iXmX8KLZ9uRlaQMe48wrcoD03YbM3dRZJ
w3SsNQTaEcireHWaF6WohhqFiN0C1r+k7uxRXKjJLHrrqmpACs4ZkGHyUkSP/GWW
MQ7gCHkKW6VNexhVzXq5qiaGJdcSFURGL259TDr3Ctq/5ZY0wi9S2d/th/2SmsFo
OT0yTuSCc3tfoYeWA/lNPEEHMlfC6zNGjY5UNzSBoQxNPMSXJ8TOhJvm8JQyzSZe
KYBjDsz/XGHXE+4il+kENfjqg5hJPrEWDhTo7C2SvgOyWoz25UVcGcNJMwD2mX3p
dW3F/WUc2Drl5qKgTxvW/ibtsqyaZ6Kc2FCJZ3kFz6RHTLg8dvV8mZPYqWfgQ/TO
cTgLc8uBVLAjyAPY7Ucuj+paIGrU+enWGOpjV02QrgNzdhcPwK1BJJ9yX2nkffvz
PjrE3lycLsG8OmW6HvSAEZfTM2cPvSS2A8N8iFGKBI0vCl3WPg4Cz67aWvr/M+i0
i6Zaq5sai2fZwUDFNrHPgbK9Pnxot3VUh1shInT2B8kFmRC7iuB6zbUtvXM+x6aq
Szc8d/GONHNYiuKvXp0nrYFTV056IafZavtYgdkBrGk+yUEYeGPzfxX+DpGbcMR5
BSUdEbwbz8l2u2lVCyW5QSsiFmIq9TIxYaTvh9XEJy6UjXfo4jvcbyOLyyOw63nE
iWrhVi30UAJiZuXH2GNItV86TVsIX3nWqJ6rFpOWWj0OGqBq2SXboPozLK3PNczt
qZ/M85AWsTF/jXtSTHNc5P5HfePJesRtaa1pC4jFKCBQWtoixmJdHdmKgLY6bweR
HWnudXqg0X7PVqDg8gQ4ezj2O+5Fh9xQd5asB4ifYnbP9iY+0Y1RTAx8P/dcKvjP
G932wnxr4Mfhec5mL0smZh+bR3Lg06Z17OhnFCLrLwr55ZQfaplGWZCbRP3aURSD
cJ4hvpN8JISH8gtt4Ox6NGV0zPKVQQkJ38BjawgBdXVRulonfID0BDOtyFGj+p7b
xNm1sw6vfGhg6rO10Y6GKELxNMOVFBEbfsJ6mKcjMZV6mwFkp0F13eeAPmRjYCC1
iRbN7bf0sKwVsy3syveaafPMzpO1lb70ijidAaFjDooJsFBIM6SImqYBUJmpgiYJ
YYPmSk8fEPzYpFsG6Fj0hd0Hx6i5Gt9IPki56sVRdOQm3v6Y6O9c3Wr7jalhdHvo
qIYqmkUGZkgv2e7Uypy/rqqYaVTFBJTlkz9RQ9QoUjyai/KfRRI9KO0GzdtqA8d5
apccvWzG2rGFzYXuvcFSAxrTWpyvsYrT5vwuq1WAmCgyrS44R1lphxJhPrTtJ2tE
29ilgvQDf5y0aGCirUuW4Ar7Gmcv68lEk7k8JRli7cyonm2B4wfBOaJfwFs9ohrh
+E/N2Bfw1JKoucUsnmAWFffVt84SPXKKaxXMRpBSYO8Fxae7rjFZWK8XHk/3whqy
JDiG9F1YArXb3vKCrjUS6CXrtOuAOEDtuPUyR6ZVBcn71qzn0TS5xjjCKitsS0bv
3qRbcJiPlkdfLr8Kbm0CAqBeQO7Vvxe7oLgRDk5v8PamaHRnvVXALhuSg6A/R9z+
kPmF+BrBoEBseomc2xecf/cLErhOg/uzLM0DmVwNF7b74GLFojsxrX/4a4lfjKbW
g3g8ez2off0yQJ75xeH//2aM8MFqG5LeZCF5O0Vq2oIf51b+gF5788UZH4Vu/Mwq
l1mmPYgaoXTN0Ke5pOQUMmHwrEsi2aGisFyVy+zfQZ/g2kWMgfF3L2SIen+Y8/r8
6YwQVE0OBngWzRj8xxT52V+4/xE2N53n8lIdPow0t7EdTL0BbHiUhkbpXYfGz6RJ
mQrZ6obR/IEHsYxcfT4Au9gCZXnjUJxDXeVhj9ANUQRKWwZmKeX5qOYfXj0EoXG4
oxDgE5bPEhtgY7BEo4fSvDStzU0hrRoNbFWbXXeTDUyWGDp2XjEJwVMvpsgCsx01
QnFatXbkFE1rugw6u5Si8yWqbVkqF2WuWz1IYindw+mgcQ2CpYUpL2UD+9UBDZE8
vDSi25TK/7lodgCpiyqA+mbZeGaCciOj0w6u2xkNISp2wMDRG7L1xkpR5MEpbeSQ
bGboLW2cppAFNJEcOFF8AdLWkLnyOwl4K9k6Uet+RIpGjuLQ3Ufw9qvpsKVNRSmr
WeMIIuSnWeyQuoGUrvO939rgl9ifMlb4d/zkqsnP2a9SQfbiY2ZWcwNbUUTq6BNK
mxTgBR2V2oFzdkYYQlS/n5ewp9n71TkiQSPo9aFBq2Oe8NbeL1bSqoi0z0APQaVF
A5PECH179pgWSHkq3CnDAaNTAQPCICHETXczqI1nQVzYHKDk0d20ky1t23r7bsF8
TOaf+TlSSfJFOEHe7HTOTtBlqSvJmVc+G4djKVKH3fFgGtlexzGpd/Zzrwovwg1T
jMgbAEceSbCZcQXzHgyaFRsFRPHjy1MWrbLtgAtdrxMB8yTdKQsqVT6lTwEu6sn7
gCdYYcD2rerk0y6+KCTzenGYTHyRaByIWeq1EuLP7Y4LnQ23dZPObpieojZD23YO
1yYsdW+4Ep2K2h+wavjyrYK5dYtESyoWJ7fJubLliwvlKkbJqYjFVadG6LrjnwbE
NmOfyxYlSYEosDEGDMiUFD08ua9KAewh2kVL3XQH8JSjbrtMNssufNO2pU+FZRIz
8dnsJZ4IfIS9rxYPLkxANYBOIlpAzs0ZZW0XOxfyJ3ecFCSXeNY+EHyNTzSzmlHh
oM1zDyeDFdzw4Wr9ApuUpwPITZufWVTnG6MjM8H8aXSLOylJuWoWqLphNf7z/QKk
KxDKK4BOEatLkK6rt4ObYNJ/UgigL8ruAAXPs7DGYIrdlHBBM1qOFvJ5eJ9rKYE+
5WYkLxLVL3VcyOD7Kl3KVYb5peQglipLWMfLY6H3UAL+EcaJL5SL2ORDAFtByw91
q/nifN3J/O48Bl1bvHu4aAsRmt9d78xqnyNlXj2umYN4DQdU8rnVSAy0dKZekO0s
yOo9UUIVsXdADs/QdOM5MFl2u30qz2aFo0wvSvBtfyLgAwFMBYKTSKws7MlUY6nN
sNAbCFzGUPDZO5LQdVrEL/25KadbxQ+ij/tMixCUZ8jD7M4EeCIaRXwOatH1vR5a
UVCTuNsDcKu9BbfBmjHl/zW3iai6+fTXoN1ndxGO3pGjDQUc7v+UGE+NzLrBKpcb
IF3IaV/LCwUIXHzvFoK9ueZUHQrkgOHqR+bhP/sUiB5FrG35ZgE2gNclPrMWm3zB
75Dk+bo+4XAMq+HzHz6jOYpqBWqZrmqg/HzhgtoA9sZB7D26nPUMHrqeJj5YuFi8
ZqTWFbGXUsiNJBgtqeKNAi64bvSkMH6vYubmHLLlzfK6SWAGLeF+FiP1t+5hQy8b
R6MfNOWaVadmip1t96XMRmSh1fPrPjPPTYa/r1VL9oK5acDlItoi3DozmNuvDMjd
4iuBh20duHVwSXLRbopA/h/H/YEUYlGX1TgJHChB5gbkyxSZ/KGzra4Waiwr1GOV
pa69WnhVCadsMfFWUrbT5JhvjYcW8WHu0PkJunSkDwxu5N+WLlwzFbzKEQ9RnLZ5
H5RRB5L7kq+g2JDIDcxIvmezBxHi5lAFfywo6mJUouwgdUGgIL5qllfB2Teu8ZiH
t6MWoSuaZ4PkkIqf9h36lAzHMkN2L+86rj2CEQCzDi1W1Kbu4nRN2cK0v5Fk3mw7
CbqqFYzoMddfl3S+0A23ddWgqoCpTe6rs8bc/SYSJo2vo97uoLaFZtvuUYvpQG8a
6o/wH53/J8ZkInwjX52aZRfk9nBOPPMH1BF7qD/QUnoM5QbS+ObZ/pHNZInjo0LO
eMzA7A6R6SRNgByXjL3WoJqPKQRkrKv0OphAFGV9MA5ZRfRkcVbG982WEuRxoFDP
KTT73Q/syaiyTqtMmdwZw9zw9jhBGJqynjHzlGrqOOhlpAdcmM8sDBPNMIWanMGc
/KSs7l9YpLa3Eb/Qv8yXnZywwV/WFV3f4OfKNvjrMqA/B+lxu2sxnJ80Rzf0PFXj
Ulr0K4qKU+zBXtoGK31J4WX94KkDmMppi/tQ7XLbyI6r3JAm/NqiPnT2YfJx/L9o
NTCa5oD0E0O+H6eb2TioDZZIgs0Rawscm0VEQ6wDs21AH/wpJyQ7Y1D1gSj0Q/b2
lWEMHJDkg81y/h05Udro/XS4BZyFPyiE3mpuCIWtmAXwiy21i0mOU0u9WVv8qkaE
ITWgFTXCIrkkPiV3NDUIt0cVATC5q2wUqpC9iklTHeVUxfeZVr8uSgrzB1zkS9kk
ZH3F3U1Yf28a/0oqdnILV/udLtHL8gimfUF8AWrYW92nq/B3iYHFhL0u5OhZpCSU
jWpaaNrwySlJl9axMOwLQx55sXIRYoXVJTlrcGdDSrbOYiullsehQzbJ8rB5NZE1
tmqK8nTu/3mXINu7+CcO2Ndqua0XO0Ssjay/k+l42o6kCcqh9G2UfGYq7ow9/I4g
EL6tMdTa8D4CGGDSx6HOZfuId+Bj+chFyTizsxxeYvskpl2vuslW+sZtoRvjFt1S
UykEtmEK6jgiWZgZ9nMyOo85iQHbGYvGeNEPPBS9jAPOHxvW5lyrfOBuPTjwz9rI
yIE2GxSeD4S7D0vLt0DVdjnV517lQZjeVWAmhqLPgqvI531MHFj5cHw/yjsVatGR
jdb9+X+5mq2uek5IUA20KUddwFE2dADlP52HX0qjGYJ14mDCfKAIhVxgwqIqx58i
JbobDBRzaIcaOLGnsQtI32YClPJgcQGUTn2Ncex1qiaFhHBnHQGpgndCHLQIa4/u
fZCKFUEojQyZqcgZNKyDDDkDYEUrnoFEHl7ke9XEeV88b2dovu2XePpp+mASfvOC
s1mNcdD2WwiTrLZb75HclnPmiSVk2kmbnMAFJhUH/lUizgR+Kdm8B4HCy8J4nxUl
cg7Kaw68/XZMUWpk4RJRBAA/dlbwwSt9KF+J8NnqB3NnVywIZHQsaintkj4ZoPv9
6LybVnE9zxwbQAQ0HF+7T5EmcdtU+gqnoX9RePLKse9iHBoYCtC27t0gTOsGNZu2
fd/NKCwsmxzzHsgH6QzlrSk8N35FBtt4hM8M3AZBdOBPw/rWD6g8BuTzBtaNIbnQ
fBaheqHVJtMuBveaXxWYl4bKTgX0UgHftZS0g1OME4A=
`protect END_PROTECTED
