`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zl3lWVRZpdVv79LKkAU2WwRbVAdQlCHwwMugyh1n1GV5rnSJ3v+6mfSWSUjh37dP
nb1Z2MbfbNli8u4caar21KlYb1defQ5MS6a8Q+Lj0TnQTAM/yYW9Gu/OOImEmq6f
6g2EPT9WIY1mh2YVuznrEQXlBUBx9pdonSxEODwqT2ihw12LE/2TnoGlNeaoU1kZ
nuVsEPDkvYKIjQgbqeNg0kDvrgP2wveT97XPXaIKKup+q/guWLm9qiY0mf7uTs1S
siiMDM5GgdgespPjRAwZPYrMQfHdSkG8T0qhyTXA1UAq+lRJeM1pKTAvdeljj3q0
aU42KsY9A2YLFCRULYhmu6PEAfHFoxz9pmeuWNx50Dd+FHc7z+P8W4SFnR2qVoeX
8Eza/EktgyB4qsLtNwsFB0c5XqCi0l6rG8ty68DhrE5PvC9KbYuejp1zJDFd84fH
HbmQGH9AyiUhL19nE9gSTjv2Zt0kxjY+9C/PxbZMLUwa9ZLB/qjGQax+XEfSsMNP
gFq30yjigqwbSvaExCv8L71oA4lXjgVLKjlprBnyJ/7YjEj4ywTEozm7C8Wf03Sv
pyixqiyrywdl8VPXZZTRUXyPB61QLFEi78SuEzl3p6ShqJOHrQaVRrSYHqeqVCYa
C8VIrBU1VoCdqfV5rRkKlINGMh8gBvhIqWAJNivW77f8eg6O/ytAfzo2Q7cFDvKT
gJCvEDw91PVXf0q+Q17INYiUnnsprLjIz+qAkp4RexzKfS0WKxVFHl/8BkYUKTa0
U41GOSPrrXrwy2TDdYjCh/2j5kZQOTY8yTD7F4X4n24X6jBBRab3urQHHMNxHm8Y
OWkgIHgLcCwwxgWrYgSYe79V3h9R5D8R8t+Yiagp2HqWxxAtr2HPwRwirVJulfI8
k2D6Z9orRiM97QzP49jASt4Fn1O9rPgoOnVzoTLqlQnjBhU0Dzc2CS8Nr+UrmtyI
XmsSXGOGP//SIDdr/wdTdYrfwM7tl+93TSfQ+X/NTRjTJzDZE1bXEfZdFUyPfYFQ
oA7McluzFVX000SZYYE9QT45/wMrChwAUqcnEcVwAE74uMfquqpUrEnFq5jbAqyA
N9Yh7XzpFDDBLdt0Js+khKMQC9IvqWShToDy39aVx1giXmp5gwuZqPvFHfsbdISC
S+KbrZZCkr8ACGUHeXIJ7iuVl1KxJtbv4tmLc7bhGqSoQZ+gWBcQRC3KNB47cnUB
BLPzcleorbDVXR2OnXUDc2k3/j2PLkW+S9UZVWSai6RcM6egbXesOxIJmxqyjiSP
8U5C54BD83LYhyOL2SVzZM5WWBdaks47C92pVNr/wZ/G8nwYebWRkqt/MsLXTXkf
NJMrqr4vzm7zmb5R/3DBYLY6YuAz/aF++VQiFQoHciwAsmQLtTIJLVnExnVLCFqF
GUFT5WCHGQGyQ9ICnbMP90N3b9JLOh4sDz6hqGtJB/1ISlzHnJs3JO1CerCLloej
pxM9Igmd/Amk2hzVCON+kN12Q48Z6OSjoSpNbg0LofIjdoIhNGYdO1RH0PwNZ5WW
39hEJYwzV9rsRj8oTDxMQA1J6OvIXXvHJIE6r/gxi/7SNiPP8GfoyjC21d+WhV16
4DtcK5D0QUKu48Eiid0JbQqTSwWz5cP3JT3drBOGYt8GgkJvLi7tKarw1ge/rpJh
2NzMKdoxz/wCjcwEy8sgPE7CBelMNxbLqxpfiUa5yRz+lAIDmKduYMUuRxwYYF7w
Rna+WvVeIcDzmg+OV7WQ5Euy9DC5USW4Jv7ys3qcTmLM2ql54cQuFNEKcrI9pIa+
BXWm6tMFEevbrJT8cTc1Wsbq1NB1EKOcRRs3dypOIJ8f6Bf3+toz6HXZC7et1z8f
FUo08j5IVuDAe/E6jH1zJ4iK4XqLeTv9Bml+WCwDumyAoNUovZ3s8VS9YOVSaaHb
r+stO/7DJRsvXb+pzzJiNC0Zf5b2hA6JW3a2Ez/cj4cmoC35ahfjwA7nDrfstDo3
VOqOSToVRVKM8vHOf5kV+qcU29DRXRQXX08Y92QXd6WG30JKS1K7VVSjRb9gjp90
/ZAAI9I9hLrqMX0y6GhQ0gC1RYGeTnIByCs3UxRUnReS1qzxZvLKzvGe4D4xVlLQ
4t5Hc/pdgHsAWA52Jji2g8eQVKUXH7YJGr/vKM95UDBUi9tbKel5RMFJ7InEy5Bh
PkV7tUWsdpl6eZQmp2RW8C8Mk8CRysyOq7L3SNA8Hcm/rMrR9GreCLlrpR1IYnJW
nMb0Vw4Hf6kKX4bgDTQ0B/WnX/zi7EhqWlm5v1M9y8p5GrDZF8z3z/1knV6Nf8rv
/6McRsBg5kpaXqxtsCBgFbzszTXHAQ5ocX2VY9lY5/SkezQQnIb48tcA46DohIiC
7ofbq5CZ53WbCeL4q18dvV+aWZ/ggAiAKQZIZhcqA3D/8gN0ry0MQ1cWQcZkoPYH
u9bTIfhrUO+/TmCTGeoGLxU9BD46Guo+Y22HHVJT/tL5iGBGp2YcGhqzP9/3sJHE
Yd9elVN9DNRbLrmI4t8nxmgXt4URC/bw6an1PSLUGRMX931C/JvWudrhKGZfIx9G
Wx8Be6T03jrdvQYjFBi/V0Xv1dEgSrzPMVIX1mHdAVtLlgDgBo/iv9YLvrjDkTBy
3BbIGR/Bh69JLuzFHKy1glu+c8DB3G5VGmmrev7XnW83NUiYORfL3ecFqdcz/Etn
tLku7O8ShqJfJw9Nvr/vI2HjwndywmW3+gKCKxjDi9dGHrBm8Jpa4IguOGs2AV3L
UytJGJ4lU6uxAhS2wSZqYfSmK4npraefGYfhfExKvnetRXuZBXmOphc28Q9DHyvk
J2LTCGAoJrawFFm8ao57ZWpWJwIsudaKTDUu+OsmpsESFPiftahcPMll80gTpO6y
Tq9KmBm/oPfdDyZL6cyKQwiMs+0OiBmGAOXfUS7z/8I5NUtif+nFy80e6NiJab9Q
8YaIDNN+EsFOFZoYskyT1yOowzU7ucJMMTFcxJHtxjrxGYtBXRHCHBBukZTvHVHf
841Kj43uLTW4DwjaYwTOdaY2MpmZ47LIOn5GDKG7BOHuv937pwzChBRe7avz4Bza
S0N6zaOJQaBKGn4mxnS+IpHm2ko4CcUCR4Oc3wOKKhBVqqByfyRAhRvKbc+4a5qm
D1wf4fFgDH4Adgv1r3Q8cptRKsGvxgTIltRjMC636O8E0HMqmm7jOsDGPZhHgsMU
Apqc73OW+C7VnJkOlSd1elNaeCkd/hD9q9qINpTf3yY+rDUIaZouwlHoenqbKc4t
pCMYR2E+g0oj8AXQrJMvmiFaSF8n1ZJoSZk+8N/63u87eQOBygRkorqom6WFkg37
e8Iqp8v2rQfI5+VkKtaCppw7jVN3ozr6NEiAp2EU6gR4ToLzoirOJ5mrBnmBONkA
Ifzi1Q97kGaUWSyTGTSxq1zP5m4IVbyrqYgHJcP+odwYy0pVSO8PwHNRuZdfUL1u
xoi+XdbBvop9OQtgpyoTjWUW+5jASpKnfCxrjEQBnlDlNKyhqMKbUp0z5UlUbGfv
/t5ng6tSzA4W78VP+77hj2rFENeHScpuZM5ZGKLYgcNZ4EkAl8d4ikVjCaSVYVA6
m/Oluhtv+MOumDqH6mK2lYjSb0FxzTy7RLP2h/BtQ/gyJzOl87rEFidErg5xpwMf
SwfT441YSONvfE25weldxhmIeiMXLrK+cjO0Sd7gEDd8B33XGK3FcXrAEtdL4ICi
Kt6m9bSljCDLHmVji0e2cFuFCduP8lhA9gCOTL91DKaDGHTplXBQvCajWikfbkLx
wk2RC+i3M9cPDQn8K8hdsMEwKmh38JSdZzM9RW4cOx9KklvVXpZy6gCyV5SH6B1K
tnlHBrrzzCLuJql8UdL2q/vXZzpkuixOimqxfT5qDXuUgylfGBb1E/VFDMu51uGH
5ORNtu2j3jf9gAnguZb12FeJIA7K1p6eIwBAemUQoYDem/NOab82TXxA/heRD4C+
FxbqPlA3IrqVtRr0NxSXQuFlGRfc0Za2YTy4jbE7vqFlFZtRKS5v3mNQbxyurVAH
TaDRdtCTqY9w/iDN6V9VnvLyLPlOHoPf4jADYyNe+O/tSjVi4ZBBo9HjrbjJCRmL
+RjmVFUWiXOoNRr9f7R2GzEPFfEBaW651Ny7cFnbIOEEPP1NatDNW+hIYY7y/Gnj
ARwDrAd7Ws17Kd7HcD46HpU0Z/CKO6J9UNlDka4tYoJRGlMwQ5Ppc5pC8f2yBoPT
pFjVgmrHmaGXaa5iN/9zwetSdJuxxC6s/IOXwjGgMvmt/I3GbUsmonbdONmZNvzp
hxlX0x2Db1H5rbylSeBAmXeOnCV/W0chuZaHBdX2qqLuvOGVzH1weEmOp5BHsnwJ
awT91owyt0wOSx1keZFHpj0MHYxAHiinXuOHsfC9VJGWSvcYiu6dUIg9JJc3m7Y/
Xfi7+WUyQRHD4kzk+k7YW4smT138Z2HUX502n7++BNSRJB99ZTJ1YpmyZkyjiHfn
5KmiIE4oPBdP2zEZMUO6A9vFcPcakilYlrNiSyBWCqd8g8XbQCaDbmLfzPNUHxiW
RO8WxSFGR3Ssz9LX+rvwRjp2661VkAuVlYlQgw8DD2EyFLbKoNkOxBOYe4b+V/Li
OUt+5aREQLdRN+5rZb6FflLxPMpOF6Mk8bwhhIx6XPifF5ngcpaGCwKZsU6gOSy/
FxcD3iUjW4QtXkMWuEryADvvjpN6zYVr86VaoYjzjE3K+EybFI5y8duiEa4UcOAj
wp9bbNSWvZA4lRhpKQ+8X+uHzxTgNLjKg/paCoFbAwLsZdRHTjb7PkK6z38Q1i5Y
H2Nfpsfd76EbkkViZfdO7fgRK8eRSQKDlGLEfooV0cuMihFHyHQMgSsktZsncuX9
wEwa5rUH6Uo31lJNO2BV7/QyNB6wXSXew2B8suhPAoePwIdHCCSqHLr+Ojil9uQa
oHyc85KhyLBaEu6GqiB+M9q0y3ZajA5dGpSvH+y20hvwncOtcFoD5lRnSbFmvZ7e
nrLQWZ6xz0ltcI/OXv1LGbIKAOXICbOTLcVK5Lp7zbRxHNdRHRahy5YOfmm/ruMJ
mJIP0osryCbUBjdacUUcVE1K5OPdiCorDzMxqggQuJU7+6Tgu6HFZuLI4jRixN+2
h6yqRJuDdUb9+d3yyN9M1kYwEJxM9Bg0YRi7EY4bToCOrIGhtQ+bfWf37tGqiS40
BKu1rmUAv3LxYOzoQRi7tlT0heY0hZNouuLxXbmduAlq+zMHp+7iUPJesoUX8E7x
YCbIHex3zBLDq3L3pHo9V7z/6/tSXsW5HAH7K7DG7OxTwSkIeV5j2dLHJQHGdEzd
p/wL6RMNUnRbCZjzKKVa9OE3lFr4WtE+IbohattsKeBSpu98kNc0ZmZySIywjia4
/wLagTDwDJOTCYbwdBy3qhpQesuG7aRozodWc3X/O3IxdQYBAYwSC8HXEsZ4rIYi
n1LL31Mm5fzp9gp8wDI06h3CetMJNBerCt6LvAQHcrwQZrPM1O8B3s4Qx8DGBMoW
LaxKbon2j1FcXXpxMQ86qXbmj6DV1TuQYiM/8xZnVqRf0ZWByy9KVNnQgLymcxcZ
KsBQrkGLsQW7uB1VbWrtqWw0J9bSOhV+9YIIJbTcR2AaEXh5cibno230kviZ68Px
3c+zu3GDODOAnO3g0Dyu4tODok7RnGSbsqK1vC0VN1NAqYDgsCNQPtOzohf+WbH0
0f+oWiU3Bw2XPPE/NQONV3GEN8QYq+JVmh0GBMVkdvvT0Wj9LZG+HdCXY+AIinx0
MVNudO6mraJ/+Ig1b0RX8ViUp2enzcqMwdeeSTut4naNX9b6V9wiggGWhnatofzY
Z+c/GvJnbWVTpcSYp7JtW7kLl6+6Rijja5l+Hbh6BerwqebMqv8NPrHLmHq1JQSn
ham0K8LFcZhnncFWt5VKevzxhKVC5FMfdK65GgUl8uHMSSS8UVEygzyoK0ZClR01
98Uj+qmFZZjIEsICNq+n0fy9Al8PDZmaKzYA5yPURtOFnYkRHraeMhgQMwuf/tSe
kG0CvrPaU6keDIYmYd4pg4XgFFw85OXn3ThniLvnysCcrhGUfiiUi4dLBb2HVMjp
by5QY460t/dWGQZElDMMI7+8tqX/4Mn34GN/OhqgRm0d+pzy9obZw8VksrUAdhlT
ooY4FRTkS3GX0dllLAUojZU0eb2rjQ9W3nfJYMyp3PWfg0SyorrQxdtLyteHRM3W
762ETcLLQVEJE5kDw96PK6P2Jgx6vnjqg/2cFPxLw1XeaA2KQLtypZE+4yHu3vke
9FihKgUG7bUnwSagKkNOX20UeoqwLLfuEQR0M4tedGc3uUDXSBV9CFs1q1D1hOco
TQyuwm0OByxXYhcrhjGlh7F9qUFpTY3PSzl+qFlXkKEIz3eZSA5YEY8AOtBrW+cS
4bUXYHbUPc/D+FvNaotfjgg2qXzY60EB+vbo7RR5yvvn6W8T61d2kuk5SuyqiJEK
M2rRAWMa6jMGAA2OZXm29IX9JOmyoK/cbVqrEk/Wd+FKHgBVRhL61d8kCx1mhjFY
Y0/D8BsQ/a96ZLAEQwzu3JD5qgNWknvd5HtJ2BQVWy7TA2ZpoNSILkIUy3R8JcLb
teZ5RTl3bYggCsU/pmpetyLt+PRaz9q24DVY8vQbXk0uVfTM4XZJ3CXndJlxmXEF
9CpbwWW8xRbLfSBjLSnI4NkLk5SjGUtdFF+KFHC8LnL51ivEw2tkGqaKKizKnlCn
ai1AmuD7+2YPfrzHO5V7IoqV8KB7C8oO4D7mt0GFZ8ZEshzo70lcnSZZUp4+MUQb
dBjBTJHR10PfYR5dQHIOfepW8n18vytFOhX/i0f295KxBdoYUI+npmN9JE7sQxCn
OlVLpzrX6N40GKCcHn79lbKo+xxDYaTUCxZDaLIs2K34q6Ht90g10jBBW4CzTvVZ
KvTJphMhFlcrfxkBff01736Hs3PQdD7w4Qpxg7kzbj0ut+Yk60buhcUvzgqO/ObZ
BV4V7YHvsRh9DALQcyqT8snZYBGRzyPB0KAlSALY1GXzvcJfUvugLbt5e6gZjfgk
NRk6TVP7kW3OQgbndWhiNd4Jgn7OZ4N7NZ+dNPARI0Q+fUYaczRizqDtDPhR+/1V
XPBN7Tk5OBpTrORNE1B4a+4+1GiQ61zi0GcqTEyHq19F0b2ZIJQ2iJVWNhYoS/Wy
RViYiLW5Fwp1d1tShJIfI1ru9Kr6AIOnbLHq9JGMt0qGKBUqhrI32fjICuGvghxF
BcZL9fGrbWVxth95z0ZCNjIZy57Xsw+HaRfcAwCO/fHu8fp2F8ucJuGnGTPgmwNh
UQk7GOcAugX9ZfQYltIXn/pvD5LmXbhPoEm9InJTClc=
`protect END_PROTECTED
