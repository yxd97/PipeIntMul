`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhPHmRe16KPWRSp7gai0atjVJbWzHHRy3uDpSEbn0raTU0cN6jqUWgy6bAy9CGOU
lZbFb8y5hnO332LFRCz60LLG70GqQg8J6R/7lKoBzwR848eyBFPg/4Opa641IF8Z
GryEUKeqfqXLVGHmZUYwKeClksG6Lvf1HhpxTTdisOeDMkKtSwEmapRTg6abp55q
UTI+nDw/B54wf35/rkLICXHRfBBUf+mSX2Ha62IN9dqQTkJyXx6g2Or5/J007aye
RGn8GljNf5il430UDFhq1mPpur5IuiCFmqhmlrkPibGHWgxg9k46IowVmhxvUF4S
OMkG8IWC31pd0bY+hF9yJ/Zf9guAG/kgb4DWWpRCUAZA5cexlNvckkfMs2++1oSd
KMG2nhTCwts8wicr/IENbbXHShufx3QpqN3wno4Fhoux+Enjnh8NKv8wT9l0VHsD
ihkP26ozEvltSwzz5G/3zDj7gzV7vDQvMa+ScNSUf5TTU701JF59TAy/5Qzqe4X6
XnQYgkd7KTtpB9ep8ldUuXTJbtYRVDgy7K3a5k+GHaTX3FUD7zbqCz2dB5cizS+y
EUhIbrHs7y0mOvQUPG5+aqeyPBNnhDfQ42rjA7lpuWAwWWXYb4GX5foT9CJtUWce
jt7cSB0BaKxBxK/JMDjqBignWESyejgH0nZyJoeZyzsaflreXJLRUGqmhFJdNYog
AVpcbp+UIX77oKS7L6sbY3PdVJq0+fDYX2NMwIys+0knnB7oENvdmBTsd4ee2wqN
qgEDw1yrT7aO1ddcd1+CIbThKq1tBTC7tuHF9mm3KpBuPqj6twwDgf8lMzLn0yP8
03RbScIxEGj+YSCAT4H5zFxqyuYTZK6tYgUpHKfkraGtchx3HfgSuHHKRIQMHQYM
9854LjJHsaTe42brJOajG9QBiIyx1Xd8yRGJGRjhL2o1qcDYg8/VIoXx+bLEzqFO
DvXo1wWepZ3OPwtkK9dnm5H+FBd843WncIHVMexD1xBuibw3MQIBjS2s1xx8KtuL
fZCgf19AePUrXsLP6aMjH+qe3rsvUQqJ+QjSgFeJkqrHg1o8+HMf0iUNc8GJtVJq
fxTrP6vMNSmSCv1EYldWxBRAyOaKg9MY4LeyH6K+1xsewX+jocqg671zvv10oGCc
`protect END_PROTECTED
