`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKWAk6qtFktVHs/Ha5o3UVQs3cc4Nh9qEBuBt3p4QanXIk7fPvzMcGefJsXlzhcj
VgRvzA3UNwg4LyEN0zx3qSo7fFIoz7zaAjx4fTJbh3zIWdO2tlbx+lBqfvuIcVCb
hWPhVawaYKWFnkI/WwouqEFf18r0uUJjopV60PZxWaHf/22ptQxjxzE0loHGZbqj
9ohiWwJ9QWd+CnohWTZ5AinPKjhpMzQqplHJpx2wRVbpswvIBEuDXdBxVf5RKB3+
1Pmzc8y3lpOjc+pVUEvQqMfRXyb6zcIn+N67jjUGEl0MFwOZSC5Oe0PyTgwYt25s
GML+i6WmBvnZUwHLYBdRqt7Jkn/z6jWFzUSUFrNR9Q2H8F2q/RlSTOWZArwrxm++
4syfyHGy5UwlXnR6C0s/8WRYutXA2ovhonSDA/703hOTDF1Pb2WC90+r8bTR1ot+
y+891bWBnxzEiDL62SNgmM2FUrMFZZ3Ogl48ue8/EWGa9g7Ka8ndryVjcDst9t0k
myjkWLggBqbVRFiRXekirhOvZWPO4EedK30/cOMos/VAnSjAAbqp0pCKEDQBoA6W
JNpPPVU6qs/5y0VV+rAqdLJxzcWZEtjrKUaa5tKlb5H19BcxenA3OBQsnY4coFlV
Rd8uzlES1YIMMD1IwpHIhZLCqCZxCtuViwe3WLNIhmf6jWsIQMby3jYoel6oJsgY
jvqy0k9HHNHsJzc26kzcac84RYNi9ZLyP35BmPRpoFKiHB+lMgCDDeORcu/Xiqev
DnyhvMAwwXwJsJxCFarHxA==
`protect END_PROTECTED
