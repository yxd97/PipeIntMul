`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8lh6kc1Kwjzvgdz07WT25ePl+CX/WnzTEMJZSU6TQrRzLhSxJzlXCqMnb55OS8Me
86L5hGsosBofcaJSbT3H8ojEQH3g0KJWn8yRQT3VIk9YRdZTA05nT8P8B3WsytY0
k4S8xdNhcd3kX5Jg04xZH0/ma9Ra233AX/n+AhmOS/umwiLJSITkuC7fS7o9Ch6N
JTy9kt6B0izT5duvFErtrIbNxTcQWb7FagBNwZzuFL0H1ltPcWNMY4Yr95+ZbG46
pY3wn2hV34GcQx9qxCFGiVt/xzHIlCSudMI299A8LpHTm9EhgZN+eNv2KBfN3bgJ
NYywID6qPqalmPIoTFZp9T/LKddoKWHC5WV2zh8JRNQIIJGUvChCUW1iycPM4oWQ
ETOFAdqBWy2Va8HfQNTQsyU1fU4HVKvuoWzN38k7HHp+eI0qJiMzw6/5y2DkUIav
C2tEyWMLanq4AD2rELhpWVh5RmQr57CpYpcC1Srss5RGEHE7qw+4idQ1/tbxQ+Nt
bliE8E4UV/WHGJaJxjKVAXzzDboGK+rpB8jBl4KpBpKlU6A8uObjwbrrlp0M3YNk
1PSq5Y4uBPGHHzRgN0ZN+QaprVajOmPIdB/PFBJicQxmXsEHnCfTqHzj6H7y6Xm+
PYpbbxP9OLWb1O0Yq4+kHb9zIX9nzMY4sb4S5/9KuzwMpZ8EVDcJd4wvbKc67XC7
ZmCkZNrDEQfT+X4PbKBKdcrhk1k4HcSt4eqsYB4M+34eyVHZyK97d3cR2RL5HJ1h
p3bGzaN02LL0748lLJz/3qmfO78S163MK/f2/p/CYnrCLmuh742RKkbwdiV8yooT
5n9Af7DjDiaUvyFMyouVmDMnqGVp+A6NCG1YeogR6HpnNBe4FJy7a38Pyf1KT9Ke
wOY+d30VG6OD1YL0SotD1DAQne/S9oYH9GcrSXOHKcJ+KCTP6gBsg06I5e4aaFqf
tWijZvUc9bkoGvqqF95UP52uL6MYdGb2yeQyMePdOl+WfaHbfWDNn/UoaNrtc769
ZCJGNWbkQF6KKom6U4r6K8x2IX3ZbV91XP7gemPDkTWkD6+dNbYAF5+9z0tW7JG3
Trgfg213DzAfwkLhXkuYfUBX2at2J1CCa8bSPBEKynFOSLQbn1V/ukBWfLx9QFb2
u2E+lAWx/+k2AJoYr1uQ+0hZ4Pt9d7sJcJVKt5dJHTf9RJap8TU8wPM82MJQruJN
LlQEhShrMsSw5OnPWM8gR/3zqpichizoJG/e13BSfO1sLdqzRs+3RkDbrb1mY6aO
`protect END_PROTECTED
