`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJUIztodDaNGiKdDRMcAhGJeDPkordrsJD/Z/hwXsWg7nWepkyfYMCKx0mh+KLtk
qBhfl+Zh7xxny30ufuAgW+TZOTDvptfanMtCE8KsL6E8qTiE+UZQhb58KY1Cj+1O
VOXrHqQLwiRL/YqeydgYKeE95drnbXyGEDaQXjndlyW2hEZPiaaO1gN8T0X5txgU
f6DDelywsrlhRsOHkVhSO4rxaihfV0uzhB7BQC8KH0wBxcUgby0MgAeFJA36/SrJ
vOJxBdD8r8A5J6UFKkM5TbWFQd7PDrM3KkpsYN983o29gMtGSxgr2yi9vt6UYwmG
1n1ki/whK+I3cTZEpuFSb83hlsO5YmjMTc2QxM04O4/529ecDZuDPGYPIHd5lavF
B3gFlaCdurhi5TF23qDzMpPDfzQIibM+gEigLKbuCO7HiSb6HJAmwxlkQZg19h79
ZluY5zM8rXKdx6Pjh7pGSVRhAfDgBFrKoAXl+jnZtayaygXch7ZoehxKLHSQZt4S
cIaisOerj/ZOV2pGiUv06TAV9/GmfRvP+t8CqL+oLDVTWHBEkxgzLSZhr9TjZqXX
+MymJ5ELm20fquYqb8mdq08RbyZSUMn50I5DpTPyvbkgDrkB6z2mta69YxNCjNUU
yCw4QMvsZok7UIJ0AEjigYt9Sf/TDagWXvm2MNmM6nCZS6Z/S3t4JSGC+z6Nwxwo
SqX8d/rLqs3U7yJmONux7s71A9xTVLGV7urCOhmTzOns/8jReFn1D+kHKFxQGC0N
+rP93Q8rfWIRr+ftjpFaZFmPZCm7G3umJCj1p98C0Xc1morNN6vUjZ3pFtC/Az/R
qkERgX2UdGxNGepjaHkp9k4kbY0jMWgM3vfL5HsqHUeKKHlKpDIcfMeVJsxo2pqv
11BhhRihmt23P8jF2rUT6/nNP8Jmn0LaYYxGaUax1+G1WistWUR4MjsxUewfCyVd
XQeDgwvZSfl/4Uz4hKpnFmrZ5IFZAOXjfsAi7KjwlwAfEK8Wx84IrLgdZWBuX1S3
S109LTNr2ZPIh8QwWgi720lFYsjR7R1tj7+DhUQXO4OcpXTtI8bhHB8r4S3pZ3hE
XYj2gPH9M5pWMm0nlWj1VqFr8NEkqQkkD7LJFXspOmlo7iLRvjfalPHhjR4rS+mj
zgRjwzQmvZ7EsGRL8zsMl+AeCJ/nyU9tLrSTLucvzkjJeOywkLczVqf8w8uOaPdT
z/oSXelnaYup6ygmdd2TkFhPnH1r1rPGrT6Losd3R+bpbrilyslnESwuBVAGuWbN
YuvcnF+Jq3YyxC5apUc4XvRJCuUxiNUTk6y+K+bXLqqj3Ev5juirUaK606b8hb1w
z9ltJ5ScvEk8r6sbWpQKjiPqM6Z79+eLBHPuPm3PIxPzdS/2gFEjBl5diy1NlJec
xKQUcFT+uiA2FHLzKH4P7M7zODUoDvplUGigafxrPXUmCvUuinvhWWTLYXn6w/SB
wbpcBcagoUSdTBsVuRE5BW1fhGUSQY9rKn4uiAMOcc3efz5b9XsEXyfH7jlrgJUC
cDVYoFNccNhHTAABRSIDmfBN8e8GStX6vQ7fBBOJyoOVPnULubUrUXSm9abRVIeK
IbORdTxvIU3/BzSJg7mqyXrTXb3pjHbNBGGK+c8dPkbqILCXjS2BEySoX/CTO3/p
HSfA0YbWDuIpsw5lSRuwJTNJL3iP9ZRZKOsFmi74hEbKdbyvVCdx5CEOfljp2bP4
b5MbKAL8OMkAfls+URy4++2cB1TKPbhZ5pP1lD672omzzOW5UcFArx7E172RPtwW
wkpRtp473LOUpNSG9jbBbN9LAcXN67l9IVZ0S57naKRz0R7TZFC6SbT5+0BjMDkQ
eJ0iam1B408jyWCeHM/K+/UdmvKQfdPN4kH7EBiXJ+u/0dg4OVoQ9dFKwi5ZAugP
bpMr5bKfZUoTDlLn6TLaH0D3skIgm+30A+ycgrfh1+1hDv31tAvKNmpxCM7HS9DR
8DjbU83bHHB97hbNOGbJs8roEelNTi0y8D51klxvYM9EgayYecCLkBAuFlUn8fUu
JFa6WdZbzcwEa/EBq3kx2ji1NGAZAjcrRyWOFuCidri9Tn9oZ/m5GIG1Kcgv3NX2
ZmHNRdfFI+ZxanMx02XQN6/t7y2BiawrKWhBLGaNRTL3omkQFSybjMvaSsa5zriq
IYn206Ha/g3rZalDdq8wRdeYSWNzHqD4VfiHz+HY/lgM+X5CxL3HAuwctm2HbZ4l
tvZ8BE86Qcm8O+HNOO7c71oYoC/3XRPKFDjqhYj5eFUiw5r8QYPkb62tmHbuFSrg
yY8VpCo49VTDxxFDGHH0onk/gD/YrN+kXPHeFCV0UETH5/C8mS0ND7k0Avnbf2Ez
oDfpvh5HunLaQX+cGHKPBjqU/jTTj3aCvq3tcJGlndfUiW+xz9eW41QfHPN8qxuh
SSiaku8LsMG9fOuZTGPB0hRU/CjMMLhbk0zWpI4E5MyN4RI4uhXxRQaO9FMOACIt
BkIHYtd9aPZoCZrk+KTeNFVKrRRSmO5QNhYp4mZ95EtNhsOdXxi2GbVHBWneLW1+
7ZX9YPeiFkItIgdHpDJRx0PeuErdcHapbmzPHIt+9q5jxGiwh2ySmQk1CJthD3T/
k8A89xsVmBZTKEOZJd94G3ujK9BngWd0NuXfCA7yWM48h6mi1UA6MFLr1HCJj2dH
RI5w4kMQY/OFkYP3QvD81Gepkz4J2r1lbHF+/Xb/bPzWKW78d/9aENMIOEN9LObQ
QS34VQiYqnpKm4yLuhROJUjykM19p9yRfg3CtIUtL2iFa+QdLHR5STmQYdPzKmFX
zo+eFxNGBUglCD1Bkk2ZdeZHvETvcVGVHfzfWSlr/7GdcOlR15fiKqE+Y7cD+i/0
ycZzlvmepVK+T4t+IXGgB9gVA4htYzd8Jb4h68hK7VH/fzcy8O37n1HlAA5XSYCC
sKrYWauup22tJKVDNZMRMQHS8RW0b4Y2NEE/tvtqMil/nku8s5RGdTTZ+xaMd6ju
U4k5tUtD6/lcJVu5Fnd6+mrIC0efpXQzJztvfnetXUce2dL283tqPGy0djfoXjA5
558wWJVVgGdnQr3+0mqee1kCb1IoZCexodqyS9TSVvTrwJl0QGdnPacLnFtakpLC
nC9QdrHctyK43LK0j2NQJg==
`protect END_PROTECTED
