`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJBIc3ULx04W4qAV6d9UslUrKPW6hHLdbuFV9eRxZBcGV8Ac0MB5khMUa7PNDufJ
zKdyiObvPOiI4yYVgSvCG8HuxNgpQA8U2uP6kUF/JY5J3w6EP8LhkC7vLrfWmAdp
VcRlXBl7WGapejse0LMJL51iTGoioigpCZn5XFir9PRyfJoL6+HCh0RpSxHCK29q
sZeHWKbmVoeyFawKx9x7Su08XnCUf4lVSSasCLrbOMtltSDu/5JwIOE8vM2jf8g7
ZzExkZ3K+zbN7AIZDzY53it9HxNsEU/B3bFFJrHtvqA8d2Do4swU7XpbruA8pZAR
/HxsCYIyaEMA6tq8adGLr67WGWJ+cz0vbHVxcPIH7XLB59K1wbMYmuDPA6UM1Rvg
`protect END_PROTECTED
