`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h4cFS5b/KVDylalYuum6sG2fNyEvboWCN+aFoA1sg5mU+AAiTm6Tw+iUFC7nkq90
xZ4FeB1oyDzK56UXnoMiuyW7m9SQiNlWC5fCHZE40eUqHIj0C8wwkjMgjcswHG5j
dDAsS91rfFGItldfH8+YLK8nHPhl5EeC4PmhcvluQO0zh1gnj9jlEhCWklEyFeqw
vrS3etBFSVZ7pt64EsdIrqvIvR3kGuOPnMp77VuE1sUx2582jHLGz6MQEyG7R8xE
y/UmYAYSEz8RY2hQHwsgWbwHZZmX4YuWMgElA68g1qSYg02Ox6vDiz1iOGu6H30S
RLEos1hEqy8ZCWetu85so/M69i6XkQMRze9H7KASG3YrrSRAjZaMSoUbYJX6UdnZ
ck30U74xB8Or5FMrwJtf7frey3tNHOCa35/Z2r61fBgjOReaWZCoDRYWLKNtYtwY
gHJM/ADKzPCaSAybRp5uikgUPRFmQ6xP8irf1ei+nma+w8zRXKFART18VPCzIjZ3
`protect END_PROTECTED
