`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
846ZHt7VgA2YtaDXH/KcisBM+Log6ApDRDNb5QeziGPvOHzDdX4iSYvId0APw0oW
9pEv/1if9Krfs0WHAPQqZ/GMhUHscPFH/tsjpef+eWDjmZFo+AqyLRaUmJcAhM/y
B7gs7UXW66/3VmSMlsHzkLNFhbwppBMlpxxsB8zUNz3ORDJUc0aU7Tox9u4cKqUg
Q92X90soG7tq0Lna2XyepuzGMrEtxWYNtGisbhvzhp14yTErOpUDiaPNLHtfOAb8
sCqEVyMaCDzm8HV1pskQ0v7cnwZf0tYg9P4MhrU/hZsP2VUxT9PgEdGzttvlIIvO
EXP1JbN7FojMl9W5V1lUKmSXzZFvP8FGP0cfVfijZKnoE/a9y47JUM49SU/rxG55
vMMwnrB+rDaSoj6ua/6BBXfwrjCrsapOflXY6gXaq8lKRwqaPUV+6bppJeFQjlth
zblUxOLmuThpW7FZm54zmvM4ad5tb8fvVOyvHnu1/FV5pEeWbgl/tqcmjkSgyYpj
CYX1M1GyYIpBBuwajxndoFs3uEym4S0Bdi+FiWCBtQagnpWNDGW0uPanLtdB55l3
VkofOpwm1u4BUn1IMMrlVX2u91vYph+uDAkk+CO7PJWPx1RzQQnBTy1tH3X9n9sD
QsMjF30lZ5FCHD4qZcZ0xcTTaevUV7h4JuEJmCOEZr519eJAUevVsLNplPdKbM8E
3gAxpzjnRKko2VgkYJ+qVbSPO0k+psfT+A8aH2Wtc+9FAmIfexrtUFJSpIedSwNf
9WOvHpCA6uNfWXkM7C6MM1fu0EVs8WZaKbfqi4ttwXFrfHF0/spAIBcAYeHlCnPd
7vxoB3FTx0g7+o+htXJ54RyPKAxbZKcff1fKrUwhIua9A7afDHkLbbQnTdYyde95
JuP8+/eYzUPkmUgyst+80ulOSKpdr/59Vh7APT2y66IV9ESG9cXTDhQq6dIzOz7f
qDBaSZT92t2sY4BQWzwA91rp9bpaJslAaX1tZFzRa48s2KF4R4L2RS764lIHwmxl
WBv+aB+f3SzljpRQqHx7vVFawD+gqso7gL29OtIpc8ZYEmhWJZqZ+VRRDgPPqr3D
j70rBQSzdgAQKfSVgOYYB/RY3rgRb8k4vq61kjZhQ6znyLwqgD0TZvLQugnXHsYn
Y8QyEGqVsfW385ShC8Rg+bIj5QwcG1/Tnxg1BHLg6X0NAEsV9KNTymJUYb5Vn0fF
97xjG+kjRQmpPgSew6e/nh+z6Ukvr8kU6dr9jm5YGqjNggyBUPdi6KmUGZ+5rAER
MIz1y5VGzrqyazu9OwVAtNZcHdIAk4/Kx77XfsYniqHU4aos5Um3lsnAQTaygccd
2TWmxkFbk5AFpmQMsjjkwwMWm3C1ixRqgobVbT/xqL7BCWVNEZ4ioGe7VvHGFs9i
cSLoRpmOvk+3xt0/3tZkX+YInSknSMngAIUBCD2Fosu09FlYQt4mTilegQDVRrOV
Cl7b2kG+/STfktWb4fbs1HS8gsaq0pbHarfgosCIwafs0/MA6WM7uLzBKnvNz2k8
e+tyEkipQlr66NlIzX4lui4GlvJeyvh29TQOCOHjFDu16ASp33Fxk5s2lEizbc37
uyfF32rmffz5d1w5hj3xrWlJ5D1CXaHhmIAmAyxPHD8ja9gAlL/+FxSAa2ZkVQ/n
GPpaukNqA5AamgCBGXUwr5vQJ/mUtX7nYrVaMgb3Qn+Q9enMq5zm32j82gvnq/bn
46f9HDELCAgqXwUnqsGRDkkBhApLIX0DG358+EwrIM16dYBOtB2AFwle941ihIrx
bdZgTpg2cXsMRuJm/J9IRR3mSGsvKFdWYIS9ydvbNxIltx1xCDJbmcAHzarZMp/U
ivzZErC2o2iO4RERJE35zpAnGD/uhpIETUyenhQXd3dJUk50MBrGvZBb37rReDm4
RAJaQtoAQ8tB1YgzmQ8GRaYSCDYoAxop1IvKRF1npOnTvMwoyJIh4PXGO1+QE0i1
L6NfOLDZT8DkxZb8C9dpE+WNzp5R8XT/naeiNbQIhU57moawwRA964DqzVp/1iRw
VTKmFawWB3H4ZlF25WMNXq4mUH3Mf0B+KKVv1rpySLOASNDo6/XacbaA3DuLERo9
a1PofCpXWxleotiSDZY9s53XMpbPtfDiI3tIPNREDtpZH7n6+g3Ktd9tO2o+Wu8K
vruM8sjh8EDYk6utZjW9ZaSaPnz4FilI6fFvyEVIri5HnouvectQEmS3WvMSq7lY
d7LPf16Bgr+f8FrC+3mX/pyOwWsbg2n49fWIV/baEyGfaS0baZWptZl3uKKlMf4r
HQKc8pckvIW/yDRCl1zs5XhdpOaZytrly9HFu1qIGAyGKQkOYlwvOD9M1D8STo1+
U/RSaJp//6Sp2kQtI9QSpihlNhRgE9H9M/VzTybBORNLIANVfCt0aYGtRyfu91IP
hE64XGf3ooxtBCRl5XXveJ1W25/t0xRXMHALEqKdjJMiT91738PNVvZ5uRrHP+tA
OLW/WStkJyWvsgAgPNXdgVzFS9NseGAR72XzGD/Ait3QDp64amqM3sjg0aNXhm5m
zQMwhtCPZGpIM61YTna1R+MbMx+mpfWRUidHxqKmX2KBKZXXxtFs5CIp/gufELaX
MZe50VauLsbSXOUqD0pqYs5/CpSvi420hl2PzsbM1gU0sAq4/K5aCAtDmYypCxp8
NKoh87NqH0dSMLjYDvP5CTgzaEe+ghm/Tfk61yV/ivQmZJfkkDQ64Mf+R5rARF/M
I+BhYmbbOW89mvpaOPdvq8iZbrDdLtOJXq1xG6hvEy1gZcFO7cuMyWd18osdIjw6
7sBBml5pGEwC+8IRFN3OBg==
`protect END_PROTECTED
