`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pckD8OcHyZlObrQurFaD8uQEdgAsG0N90EpdP+o+PIUEGJZ8IXqtufExL+Uyai/A
0X1oAG8g4IHsC/KmnB5at8MOxb3a0MMJ/tLSI7CsYEb1EX6oEE90dphTFelI/0og
3OJvsFHWR9kYafhZsYb2F9EmoWzerYXNLxeZfc8WpCqkKTDtRzoC7zAs7WaO87K1
QNEWjo/U6n/GdfCNS/0Z5j/+A1kuV2CITRbiy5B4Hq57dwi3LzBlpCB/cj1lQcGJ
25pFUdr7Y2cirPzKkiGIzMAvJftE02LCRDvw/mYbsncfQ/NG5V5BPmQykErU4qx1
Eglium0jzdVBvifVn/izzLbnCXE24ndcpTdbe110l+34X28OUSKBvhexm8z8Bn3X
IJStFHy4b3nC7nm6KHUdtcxv66jk2tWw1whYUV+Dn9d7TfY+0/rByxC5mHakQPPW
`protect END_PROTECTED
