`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KVdBQMcuOehUOtAGEHNklBd7x1Jd+htlPIdzWJcss9vvZRvWIKsj8NiZxhVAY7k7
5tstGlME71uW+92cQiYYJ6dFuA+yfcswjeSnyOx0OVpMixRoElqhumiMVtoxUib3
LmMYTMl2D9dtNrSEYbNwJLzV7G8M27/3eN2Cb1OfgcFW++LMAo8Z/NlOrVMKAvqo
RAu9oJqGmEK4YWiYSmbAgWwFqzagT9fcyfuwlnMNNomr7g2PTnbSJZbc+8nvgvWn
gq+vGxCZRnsX4WPj67Lcku6Llx7qo19ygQlsBfPnqSnY+nRLeedCPXpvwc7ZaKSb
d4CJ3g90QE87pn7is68viRGoYIa5X1NALbnnRuIDVYVy3wY6LnJBHvjssfVHNtD9
TjJhSTJUK4xwXtoLwZfQDaNPf9kOGbm8zK67iKk0Q1rP/KP427fVXXYkD5Lnn3b2
dbIvE6YaRLyzIcf0okPvsvwua9hdz5TKp5BRxdg6s9F5+mkw30QddlTqheNBmix6
xsDN5iUzOGHR4uDTs1ygdX3YuZuvePtswFXuMp0812RhJJDzFie7gJJ3ztdZQIU+
CrzTJy0MUqT8PeI/PHZatBk3jMvEzIIFKA6gNpGhmv3YZeiPBYl1+pJD23xQG9EV
9NumSh9Xk4W500UTW/HNOGATg1P2HrojiYVTNfuuakI=
`protect END_PROTECTED
