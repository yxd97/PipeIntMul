`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f59OYL+u78M5ZYNi1FAN7jRYaF0tw6YkB6VxWreTIQhroqsb+Zo7TcdbNYMM4tB6
rOOb0keM/VtdGtQ0lDzLXr+QOh3+cFMD+0Pkk8wIL4pOGc53fkIV5E5f0dsjj3LJ
7G2LJ/c6sxVdVHyHF2ZCGk1sGU9lY8yzCnZyAmDFi1LqaxWUF6bTnEoJg10TuMEm
+D6mU55+g2ebzcVAZeHgg3Ol+Gn27IuPjY/sVfTtipFgYi7SZYd3W6OOXTwT01S1
fOkDCb0ttaTwiyuGCTT44MdVR4zP6nfrr+d5zO9yGk8mXWcFFWNqAkBb4kJcqTRd
F63S62d7NBpWq7VSZZcsTcY/yD20nTG2H/wIo+bWDOsZJ9jNysEzO4OmB9z3vrZ8
UFVxIkxPpK4e6zn6U/yL8BHm03pZtk5qHRu7c8doBtZv+/nyCfpFGkt4AfOn+aE/
AqvRXEDWLSgczVd9j/7ooHBJnOndUhvl/RUIGO2q9D0Flzg33OYzkjnVZj40okQI
`protect END_PROTECTED
