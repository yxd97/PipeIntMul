`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
158dX6sMrRgcEQmTPX406R1d1cGZ8iYz1xoj7G2cUVVNuLZ3MSK+AjBChxiRrIzm
XG5aLQKM5zAosS9ubm02mYKDZgXEeKxZGxvzwzhxX5WPmPD1qe//l6wShMhh+stA
Gzvv1vhelAVae+puwiSDsHn2X4U8iL9cit310vuQrR6LR88rSiAsf87KckrDF1X9
79xoIT+FHQAFJfBiHFSG96Nm5A9escptZ5IySXrM+LPL2aNHKR1OIp2hMBHKJs7s
yADKn6pqV7Gq4gercpy+m3ruAcH9NvypMTpjK/6TN4ohntRb9w7Z31IuXzeJjC49
ygZcl1MGPPEzl1bCIzpCfdFXBmNNtBp021a4rEqJx5yEaZtv9sKwPSx6/o8gD8nr
yla0bd9ebuJPos/f2TrImiJCrmx++4pLlPZ++BnR4/c=
`protect END_PROTECTED
