`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ainss7K3H9jY/j+gg84l7XPxbnHVTCW1iaRhWC0y8/oAV7z3m/9baDZmHhBdlmoI
x6JFalU75sFTFXT4VoGEgXNtqXdMneaimgQVARUDPG2Bpuaq0XlN+6TYWRnAYwju
2Wde/ED8Ge0z+G9+xSXu7MmiO6erm5KNy1r9yzlGEgAgZhjHz4E7wpJtJ8xmroZt
ZUQOqN1YplP9DlI+DQPu5M+MaepyCtSqNJWPaTM7IC+daFQRoQmVT9bn2I959Bvf
bDntiK2iKRbARajLw68gL0Ngef0orEBd964afzcPnz4JCnswVRjEBJ+ipFOyIcoH
CCggPaOO41W8prbyrxuBzkCH/YdC4dEv524YLZPI92/D0F4NniaCRUqEDWEYm6Tn
HE0O9g+41KlINstgvJ1NqJ2EMSnLe2Bbnq0CVBaEs1lLA+bgkOxlJZXjOKXNo8UY
GlVTREK/rHa9Or5XLQWefHHv3FMFPvVLWHBdMwA7YheTGm5EtzNOghBIaneM72W4
MvyTdwkFlf4xoyGZKMlb6BcGAitF1PvTTYmdqNvpEhb8BhKjBp7nal88uEdc9D1c
nYZG8AbIWw2KfSJicAskxa2g+HRKzoYrA0OMXXWqxBQZVElwTDBt647+WWlk7XWJ
3Hz8azuRQWMdCPDX7wwV0w==
`protect END_PROTECTED
