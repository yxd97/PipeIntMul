`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BOlnPzv+2FJ+h/CR70bymYsnQzgyaQM9MPyJYcN8OplYve15vd7K9BYwxqkaeN9E
MUr2Cwt6GjIlY92KJ9xIQYUkrM3OiL/Cj7uraLj0fXlrzMR/K4KWYi7XaQCyxpuY
h9BEjvZXp+HyN20/zTdZXR4+XNoYneEMvZ6PjvL+tkYW/be50RjC4XMToO7lSrEX
/21AYPVtzga8+7dLfy2oSAX6kWGKew/uxWp5414flnajfcbFLkiBv2tTepH+NTi4
YntlL6Rj9JdyX3RPWK4aEdOta9dbPN51Ll5smaHo2yPAh5+VtH4G3mKPGWRLh6OZ
h9AudzNvUvAvTWoUFqBYzyZ7FWl9SCCbYbYwq4X4z8GJZYwhO4bndGm+jF/krvww
IK2IRX+p3Q2OahqTVcIlG8MVztvy4nAazCbNbHdySfMqf8d4jU+UlWPv+5kq7NBL
zyowgiLjNLZgmhXfZMynMmmdKWzuvk3YgzjBfRYMvFuUFgkywdJ4Sf3XXc9vrmcn
kquMILgchjxJTtU7evlgQp7OEoJdjmD9UHnLWr1OxTAA7APhVjsV4gMPHgLtaV8s
5qzcgfQarDeOqFwPEr86muR/pbyh1lZNu09R+Ie2bcQCk15r2AtqHjZ6vSNtB0Fp
YA8EpJjwK7ezlcOhvs8ged4sfAf0fDU2Uoj33Yh16+fNQR77KOTlyG4n9rsh9Ejk
gvnwJ53oJxCr0zFKf7NSuZpdF9U6/sd+hEkS3DN5nV2htWdGUtyvXZuATteXjq3/
xqvLMreWSOfVUM0BNbDxAw==
`protect END_PROTECTED
