`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vz12egYTiZH6Cl6zvHq2RtxWLz8VOJ1iadXczIoo/0uWab7azQpNlwlN6Bf6ydrA
X/KNToKOoQz7tb00t2G7jdazX+eFEbNt1gDlHsO1l7GA0GUvR2lcM9cN7IFymObw
aUwKEgSDb67HeO7ooUufLO9Tm8xmxxjePXwa1m+2rUDANzegiF1no4fu8l351qiG
TjQ7wZUGlUrrruytBUsZxqVsd34pHF0+meEpfU5SH3GBH17RLCgoX6At9gkIKuDf
0EE7zqZHBoFlyStC17LUHXayAMHyDtp1oED2l1V9xEhR4DyDqTPzDwsV4rEkxcU4
JS0DoM9b/gbeDE7zkTjnmdQwcGydyL7PryliVaD3y+ElDPR6LVEK6W0g0VuV4O3v
d0FlN+a/8h22gHds2EMraV8nx0y92AuXtEsteyRAR0hjQmh57HoB7oHRwfF7kK1i
JYut823DhWU4y5pRGseAAc1VfcSyLihExyYeGQBM5CVZ0D0dHkn0QFegoRCYCQV2
0pizIAf4CVaek2iGo0OF0Rj55cmYX3qYHHTSgnZMyTJPyEYRCOSgPnssofTj+lE0
J11W1f5MQp2vLzb5OsqOZhNCEYkrtN/7e/sh1gxHhP8WzNDUJlqoubMpOVGWfYun
mALxQgE+QJNl8ZTqaJe5KyamJyUXTLMR7WhcJATppZmrLXPJs/c/7MZdjfko6Tm4
AY4Qb0N1Osh5SLHjqcQBz3H3l6e5HYvD4kZIsCPn23I=
`protect END_PROTECTED
