`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIYstp4x1750kfT54a9lnEWnGlSyXscjQI5TjfMf9uxhyZXk8o6dUOpYq4U88RBx
3OBXFzK5hB3/yzw3dSfymqx6K3qTJRH3Xq0G/kiVHd+nxVB/TdzkpPzETDiv7KG1
/BpeNQXWZ0X0Gv4M+4uLN/Le1XY7ba9ziNqIejEsVOdFbcFrj3b2jPN5N0PuopqX
o2tAGIvYa/NIUjlWy6T/+GCxCKPEhaACmuuKn3GJJL5BiLxX8Yed/tq6K4TWpYpS
Bib9Pz822HADitbeDgqfGBdQi7xHgUbgcVEPCM8EIG6yAuPj8V5YQG04xc8wfLHm
IG7kQN65gHQ6MIVeTlmoiB1pw/tZdbbJCLSjuBbUXsphXsZdMQalAC0hylDtqTPB
eCK8WD0MNjcGtfsidVs2hlHXaLLQc1VoBzWt4OST7zng4282adidfEbKJqbwdDkF
nVWGvxVQYedJJcnnYWoKD7itAml06JdHf2qUPNV9exN0OxX2fcqWKUoE3X7/KBvf
m2WiyguD6KNtTyLFehISdw==
`protect END_PROTECTED
