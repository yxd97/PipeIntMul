`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
heguxcHb8oUidxuSk0qaKQVx1a/YdYTdn2FiZ2Ygug4IjjmwCuMc5XkTIQ4233Cc
oIcHblKff6OGIepl8kxaXnJfObUcUh3DGHkVAZFtevvlGvqc3hzzJYJt7K6KHHTU
bNovcgh3ra9oSk3fZ14sOSvy7eSlHGkR3BIAyGj1ClMKbaJATqU5KkGCBh7tcVrR
wfkY++pzyb5yWWdFyb5u/QeX6aIZEUDFHQDkUV2a0kc5Pxfhb9JAruftlI5ki4av
xrzVKv9i9LXOvimg0JJW1WURYr/2kxUP37W0SaxneZcpYD3CBbJWL/K6fQ4Hekpu
Vr2JpaPwiS0kzLfPi81t7GKyvgT23OS551IVyI6D26f7k7Nl5jWqmYDU1xf1iSbQ
`protect END_PROTECTED
