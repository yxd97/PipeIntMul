`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sfxk21xlQMXSESvjQK8LwuDDnTfUL/6V8RLFKyANKgCt2iy2tiV0tx/HsbtIakmx
s3ECm8h0KNXIdKwt4v/9eBf2WZPp8e7vYvLcDjGrQfYWC5DKQkEi7t5BR9ox9+7L
ZQbnt609KWMiXIzyijXDHoL9lQY2T+hnhKZ/gVsxPXzgZG/UJDzdQ+ldaMEjnBjO
PFB1v6rwW3NIEbErGTkKNWenaXC0f8hUFuZMtAxizFRBA/NhjfthHdZZ0Sxz3cBq
dWd4rr/jkDZmqNh4dYz15BQswWZ+NABXdgZKgPwqB9MCMRi7cIDs+Qa5UfMiuU/N
c5Hap983ADuxxfcBXxX5xHIO5IckV1MJLu6LBiOCT47TpfJlb2Iv13mQTzz4kdIa
E+VJ85wwGVs3O5x9GqhmofLeKJ1qZYNYjJN20rCcAfwtaVeLGSyJRwOxdcA/+7bb
yt/C21Z52rHaxyN22BYt/AtuUEG+wUdUcyxgblnWPeFWXgwlvNJsrcwTVsPqLfCh
M4hA+aIYYn7S2E5jlI1YM3v4VJi0ZCZ5vWBYtxaEFe5i81bvzDRpIc/9SJqw+1PF
iFYMe9TvZ3wr21gG2jwm3soDBUNAvsbQjhZOY9/eHGkuTxtjUMJ9P+JfJLp+tpB1
ddG1F2XcR6iBWb/WdNUmj5wXe4J1w0Lz7pB7Z2nApcFqOkLcJoudj5z5rYZ4n8x9
nsLf/UuqNKQAzKfVozg7VijpC/4HbxZq3L04CnKyAGjn6sAo3cJX1jhdktaXNg2Q
v+hTYEqyslB4SMuN53JCJpVOcq79GERw0NyprM03HwWDDoJwZbgdAGpJMxW3hEvO
lyRWmNXQZpze7/QhMyvpaO1NEcT7LCJNP/MKA2KpBR40bw2zKTeaZxL7O6STQqCg
tH9qBvhdLaHw5bl0HhkMIimOwaRRwfG+DYZ+mv+3+2RN79W1NazIkS8OcL9KkMOf
koqqA0cgqDP/s37SQKCHuJf5Ar22a51bV9QMqD7HIh6/6EYRSLq48P33FIa5Y0+H
1x0gWj10rdGH+5liEo4UyuvGw/3QyyFILqMshf829ZON5vVsdDNmSM+4YfIfk/gi
3q6RQs3W1zNF3ivAy+sszdOLzRjfxtdr4NFlZCUt6w1zkK92XqXTO3A+qgXCxIGL
DSvu1l1nPWpDrt/8jOhwY7FaSNdHUp1NzDWqQZLbrYkT4f08qv0UDYA/84EDrljO
Kt+T98CgjPrCnIGjyWsjQvtqb2NNW+qXV5D2Gij2Pzne2JLf05k9kHuE8xXZPOu5
t9sL4u0l61X8PwVI97v+KEzR7iqUzgiOOZyPbTZRB7bwkt19jfV/yuPbtZFTzv1c
DAPb4YQNNAt6E4+3ycfrzOnumxTFVNUK/aysNAqJq93PEhndPRALYh2yGhQoecBA
KddNqXcz/BEchtA3d4Ds784jQUS7OAZ4OEhlVIl2IMacgOPh2tLB8lnR6iJbiGHI
gxjtf+4rtW5DMBSMjWzee1Y/NTELgYjK9zDw3iYTQWecTuYkK0rnzlCeHQwNVLRU
TydDDgNxIJjdRlZCEcMQwLjhn8oxDjFRLA5N2kRohjLeZO4gj77IDNd99TDu2+y7
M68Adh54DnVK07gpBewrw8/L3+fQ03czp4Sxem3Rz8AOGzZoUl9wcpNdlBtqxE5X
iEgPd08aNEkay/8xlH3Ckvh/RN7dYs76wAgIpuNHdj3KpWrrSQRmxS2v9/NH39Lg
DTsQ132pSuWXa0SEd6UrKPucgxWnkpZF0ixA7AN0jXWzer7/dLLD8/BrntiDh1GR
iAdqCcp4VDALLjC+9+4IQL5Ho7B7pgwvjuRLZwJyuPvrXyAjuwelDUZM8zwII14h
R3RUdXZhJ5Z/e+JP6VdbmqCJaQkzseio5w+9EbpCxy2RYFDXpYgtb55mYloUaiAu
gOPp2fxdnBJiQFH4hHE9MFv+jupc2tQ+7DSgOR1T+Rwu2gjjAWX0vNvYTA5t4axX
O+HcQ0hclANkqQFyJi+E8+yB03cDAKcXjaUB1wEyabmzBj0nsc8/1EQQunfU7onJ
k6T9LFp2lqRaZSEEIu97u2mBwRq2+8LiE5cpU38Z9vCaen+TBRsyFWEGPEShbvJn
NxM18AzL6nr8Obj1Zex1Z+ahL5XgxsHhzgaepQr/qGvsZKVNsXietpusmDKDOenA
ptVFkmLJsPFKzfWWMsCSbEwr+7j1ATNw5bGHjEEL6J3yPE1t22dbMFB+SiVXc3dT
zxFP0MwPhBlck1FVHEMzobvVUZWbEj7HMOJC9S9NpysgNzQzKExgSdpcPHAHTDrj
0TB3nHdyitJmvTHwBalqcxw6jp+ySAZLuzSn0kspcIOalXbmInzsaapgmb8sQ4fN
XSX7DKOQjcLZiAjRREvY80o5UAvL7hb43Wd286cJ+VYKKiXDh5tPIPlCEcwkV6C8
jJc9nStMHPiF+5d5spihwuzJYUrQlYvK3hcHI/iRwzMX5cWO2fl+lq1JuYzOy5l0
yL/YryT54N5PPiGzlpgjl7mfTcAflUn1ERliFpxw+hqQ8Q9YgAB/kHgUDYbnvnqc
UYpBkgHzD3R5mMclBIb989IhIC6+kTceLIof/s3qkVDDoRELTKuIeaXbt+MYDzPV
pAlXNFDmKxxtkkiyfnXsYpvBPl5prfUivjkz6QATE7pZZa9XnfvXNeylr69bLsQU
op4TZFjqxXcEvDrnsfDMAUzTpteRtlZQOVF2pq0S6BfYd8qFtLi+wIYVb0vOvn0V
QOlFdKW8oXSusCETuAlViLVArW4oIEAEJeBm6iXNxbsurQmjfbG4avgrdt4Eynfk
I9dxViqrYfpS0rL1HVwnoSJiQ1z9zyfQj0NLf1gYAtb6Vo08tpaNNkS7ZrA/3ziJ
X6kXMx3Iq4OQzliJ0e/9bTjnfMAfmYV8arX3V/sVyPuea6GWGtZXi6GxJiSGNOxE
g+Kk/hkg5G+1FJgSnTDzeSdt3o1XaWIFA/phqF3OWysfU/K6ugGhoNybIghfIKPl
A4IUvT9PDhH0LjEFO9bL50IO22+pdEmy8d7UDi+SWTP77HyhqW0OEzn5yQCueAfX
lVtVpXix3OM3iVkU96/8niAD36FExEJGCtGDBdWQwlCS3Wr6OYx9O0m/FiI70kfU
XMFs1OeFwlhgc2REyFANMckwkq7Z5cCt3EFmrQypzvTzHHXF313loJqw94ym0vNh
k6N/IL+YcbXiSuft3KwFkGnHeFxTOYv9N/fu1gS9Ks0BCTV6U5KQ/ysQwidWDan1
6NiiEaAB+u92kQ+TBgW8+GelLAUtndOUjlyHs6AZEIvtPZExJM5h/H0Czq9IPy0v
hBFM0wkIJDuhoA/pe5atmPEKE3diJQTEwSkASQRIsAPM6HpuY0VxZ89euR40UUQx
qOyjj1677sMnHdfakmvxiPLpuEEYrve1g7Z3m2zO8JNAE+kQyAGIpEdWwomQdfiq
+Nc/75UIho6F3zA99uaE1zw3g89oZkGf27YXy5o7AMZkOG64JKOz9AMknn6tpWzY
EAckWHTIPtoWLXtTg50WMX9TIVClZJCb2uFa1feM1z18c4VWC1ZrvPxYBKw0YaUn
jCWr2llGuTCtkzBwXaYb6AmuaHa3tAZ7dHhjawsdslAaUiI/qxPogfmrZGS69fts
7RUJxC/jSvi7qkNlGwnFjfj/RA+bfOlJ7eqt5RD4HfM8mNdEqapa+PFnIwXv/4rL
oPvRDz5wSSPbjew1iq43JNecQl+k6R0lcbjpnRY8X1FM+itEW/bb72/nOFuuo6Ql
r7jvtmgCnySAQ9eL2GxfoAQJgRqqsUsjrX4HejTnfub0HR4KIkHQv/tvqQeGNj89
xRCb4XhAFaLHVL7/7HFYIelZqrssnX7tEsSCzs0iwNHmxZ/GyA+3VWLkXEHZzjqE
fdQmTwbbWfI9B6H9H+rsXqAuWt9HHJNhdYhHldM7HoPaakxzSAtUjEgfWyWehPTm
8tcyG1Teuvvmv1yf1NNAfYNa4JvivIe27XpTY5xeLAvQolHNW0Oauilza3hQOXXP
LXX0nujvlX6YA/9NDmZ0Qk4R1Chs+PWpi5IQXFNJGiuNwE1cqdaKc2FAigr0YZWt
LZs/Tz91dFvWp6TBlmulUPuejhOmQS3AqDt7iNaeVL2aYFMcYl3ZSQmNZ1hbuoF/
RDiNXNJ3lLFsaH/whyAFwrQww3h/sUixZz9IjTqNrwX3fTcNN/Tm5OFmTM96hL6w
v5OzZ7pvXysNzxeITCRkLPgZcelU0QQy/TzFKgLfvY/t4cgjf/+BBD0NS6Z3rgvD
jxOlb3cR6L5fJIMfacDSgDVfy87B7C1MHR9KZv1CdSVKBLiYlsncB/Nu/QJtpGse
1Md23kWaN9GRfdNTuUoGkFL8zvehDzjoxgApMHL7rJed6PzggOF057+eoGFRdGoi
Q71kD8i1Co7DaW+ZwaV8rdSEOvF5MLezTGcaJY2NjfpGHkRU/MgxyOREq2CGeVV4
8rrSZTqKcpUguH0Fc+iAcfkQo5uHlLCw1SZnH9c014k=
`protect END_PROTECTED
