`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wLdpJOIQ52xg/F933L/xRFCfGyP2ZqfuVNqyRkuFTbtPpHwrlDHpdUbcYYgu4PT/
BftzlqQhuZfNbqGZJugI9ZRfgLCIW8ol2Ss8h8QkOYl2HN8+9VKhet3NI+gcFHFo
NGm4i1Ddr0gWAnXAir/HxlKrlQSF5D5alwCG619v6E9Lz2FXKnUQwOP+uUKy/SFn
lJl/2YxjSbugSpt06AsjGcz2rlmi0JgtiG5K8onazvfecizoeSoDvOxglX8ibaBL
Gjoo7nWVyFn2Q+U+VBYp6jrfvcKSE/1L6wAH/hOG/eCAbPx4ULQ7FOdNbxMPg/0a
+UIhVyK+UTjhsWInPM7USAY8LTMo8nuKuicoijkdpK7ai1jPFweDszqdEyKjLzxK
lhP34zJlwwg+ZYp8h5M2AEkSulo52r6yfMRd848uUbg=
`protect END_PROTECTED
