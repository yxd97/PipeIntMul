`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mxcqJYj5h3hKRNco3gV08+Key0X4h1V6hQuFDRjb+Mwl6RfYdp2dVw9+8sAXBu8y
c/tW2VUu1KTA3FKsLpWVENMwK5JYXJurEp3eNezXjecjjlwYNElhneYb/xf6o0tX
oYZYosjJZBknaXmvcVIj8uPv36v4Ba99HOGRQBvHGvzlIuxAnCX8JCa0i7+SDbcb
PZfo6FfxJ1fdVWGHDcN0EBLzSU9tDs6wTzKqrNrvy3SeQXJ+AX4C0Ee25MPgVAaR
VX3xE/WQb/WafXg6mFMFFg==
`protect END_PROTECTED
