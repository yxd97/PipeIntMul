`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdC+yx4SM/l5j20jB8eVsV81E5OHcftZ9AFTAF9NxpyCR0GVY02ej18rRHR6RFyh
eDxFB7oL1izwlZu3OkB6Wq6piJBhnqoauLWuebbjDceu6M+c9D2M9C0rGUUypQxk
jH5dFkWWLJ+WJpK+r+rdkLy5WXh9Ey+a04Hd+8RP2wqtiqXrH7SmTdzKuV9pV2mP
deK+c7wB41BQytDA/S12rNMaxa9WNfY5GaRYOmI72DxoruIriBaUqfJmnsFJ9D1/
VUn2SFv+9G726ljAZUSx/RkKkxfLs/96dboo8QnxMOb80/neZmxa7b2/RGiXKXxW
2hJbqVsdIMiRd1A5EaC+vRQMnLtUV3sZYXNLx+rstrvK8ysahW3IdypbklZ7sY/3
fygBV33cGyI5uvM5/gc1YSGugJvTOARfea+9WTl6vs+grBqPBfW0no7C0zqUyid7
KZROBwUveWJs8dS2OzQ831vTJ3tDElP8h4Opi6YeeU9stWvEz2yrJsde4Po6AMO8
G7lfjYHNdDzMv2riScFlmggR/5FaFqEH4BskB4Iu1rHP2Fq5bRbyB4rumq49a5G5
BZKW4XpnKLAmHhSlyDiFj0VQn0/MmwtC+lK8ahaT0B5eKnXlr5ZvbRbUV4HgUyZ3
j60SDYKEylT2x6tODDVwk68U4GquhCA/kAP96sFxwEsruDA5giXA3PhwqXCc5Sid
5Ld8rX0g1qbxloQ/82XIYpZ8EUDmOhjuXGeaJI6aEZC9K7fo7A28S26YkX/OdrIQ
/LxByyYetRf8GJQSPXEuXYBiXDf4HknHh7ad4d18BrotcvZaTEetCvYcdJ2d71nZ
CYZdYEt+zV6QhSaVaYi8W6O+DJu+Zl1SWKZoMAQPOnHdqxBU+CXjFJ2wzLmMx5Il
2iBY7nc0kOb9A5HNk2/Lh7ccNYPiB5fxo78QKfU7mDhTig8QCa1iT8UmzS7NBBV1
JzNAIoZAQXasfhUN2TPE3Bqft5EnOqKeSXOYS/zQ48fvtBQ88YmBwSXo3xlsaOcc
qzO36oMrN5nNSRdIKw6Bf8YJUVbQKVTHCRQMnDBDmQ6eRiRrfGzCManGGzM368P+
ow4T3wLA9sXQ0e5pAnOCcSdREGYps+NWogN0M2wuSJ5pTiCARtf5q+/XLttp9oDo
0n+b8/Ii71oI66nI2Qx6InchQactBbWCJp/OOM93mbxJIB31xavFZDZp6Y+D6t61
LgQB7EONTVV4LuV3w1k74C9YnHqPdYmVSWQSaAy8GIeq9FCKPsqymfEav5kUw+ee
Hnzeqr5VXode9Pi5Gnwkpv8WUdT2gpDLagX6dNBegNm5tDjIPpRDAtnlJx2DmKWG
pHH373CnOQpzCVhywM/ReBoWoYv/4whAAD/ef/SS8d/E+0DeLgsm4l7pikoovB6o
FvUcf5hYbrSz7YkV6tnPK9b5dXWnIIUL9p2VmpUd89aq9PlyDCausPzSCDL4B2dW
VCMlAp8UuvxrtXYiiYNdwJX72Yyx2wijXnRI8kC6nkwza4KF66BV/Ur7dyvhcyjT
5gk/i2zoacNnrZiLQOY+lNm14p7fCJ0cs7+0HeR0LDssni+9iutvRC+bXTVEyi5c
z+PT8NMYFCOUeHqQocJq7CXz93Ub1u50+2soPI7HVEnHKj4/inOiGvRWCNR/hkhG
6RZw3RklOmrlV33ZC6L5xD5n+gFu+pm+pqZL5zlrg/5nNOGKiZaKRkj5tti0S27C
ys6t6A9qq9xMveYc9TotNG5l33/m0mcJ+vOtfIJxnM53aYEmMCbt9L+xy2J1QyOF
4M1qRxnJz8cA68qd7zO/h9FKkhwt4geToqMyefHgQVXNfsqY6qgRb/q1ptxWaBAZ
lF4IHpZcxQ7SQDAOgoAwTLypjgevpKJ2T6t4rTQQTnJFw4fu8mMU4r81yxIsPHNe
bkVlg46jGLurKKKj4bnnZ6zxuCzZ+4mOMEkz7euyRFlhwwhaV6L0tApnxOpsQu4l
T97EpAJiqZu8MHMJm4T87ZoRooVDuetLNJkqgPP1MGU+s6JEOIrXMQNUPZsEiXPo
7Ze3huwxMhmLXIjX5STOVuGIe2Rso+snGRJ+3NlFWwto+v7yETQnHiuC1CSd70xJ
m+MXPWqa3g8tgqS1dhsIv0TFTVFVAb42uRD7Nl77n2UpoqTTot8PP73Mv7Nt8POr
4DREl0HJo59ujtpIJV88DAP8V679+8ixzS1/R7OjebeZVEOyZZMSOXStTxliBZhu
buj6znWSf6kgB2oeHTfsw+rffl1uS0I55O752dWNvKh2vUcMw6LhB11TU7XIv1PI
Xewq37durTXCTP1ycTonFWLKBJkVm64Wm/OA/+HwuAWOz7dV9rW47oGxcBTd2o1/
V8TcsE+2JTji+CBIBtPexX/AmY49tc4NZhi6UUoqnYnpe7OnxJ7gT28YMoB0rLGe
/08xSNbYcAWJk8ZZXnVuEbKTfzjnotA3uQOGUm/c+yi8F8mFB4aH5IwDlv1hn6EN
MEhwfQdaIdqWwolPmGGdgbQbZBt8tcScmcjV+dwyhnYgSIPXuw0vPB9pZ7C7FPqg
7uQGjeaiiFMi3mXfomR8hK8z+g3fvvJwW4+bv3pvMGR6r4QTMTk+eDoxs27YhfuU
FJlweR0ywiRoxXzZ7Rpp+rDd9z1WyA+hFdkCMv3eZRPoc66rZXNRznuhnkl7ocmS
TApioQ+TsmGI4Ci787Wr4oE1Rnm0fpLga+HsBOxbFWr/vN3JTx/Zf4Ruo4U65bBg
PS9YOKd6DG4rAasemJ1r3RDgskv1nxS5HRX39xJhVW/z+GB9C+shleoTz1gvd7U/
8IjiMaTRczzb7uGgxOPfiD8AdiUmp+2fNWVQMwXv5t6hHMC8gYcl1ne+6B2anB0l
Bpfivmeuheq2Px0LHPuOUtT0Kv8udfaLA6MgNIjvg94eax/vjrtUgxaHyPu4JrGa
`protect END_PROTECTED
