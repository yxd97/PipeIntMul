`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wm9YDb5rS73/XCFwzUGQEYzrK9WtvxEVo07GVNOAhEGc5a/zc5MWucfb7coXWcWs
oifk5jAVRdq1dgX25WbEyiiq5Iu7lyPW8dq78W7W5Ls9mAXviNaPXyfrh0oPxVyX
DMMBhBmtRMtOOp3LQW/O5ulLcf6dM6H7nacD+TIaalcEKF2ajs1Fj6DtRduzAwlB
CuV6ZwSUUbSOy2dYKEB5a7wlF7+BQZLkvcIZ2IgpWhrmqXcBUz0KOd1h3HFhdcLs
EsZTO3H4QSscgD8lVZQAgRkjWZuqjWmyz5JGpfJBRZ8PfWtmlvNuGlC1gzTnw24W
WvWsXNt4cE9vohR7MuetwzvVUpssxHU5U1GsqQr8tFQP7LsMUfQFmItBlOtWlZ4N
P63fFHQylDbkjVfwgs5bkgzANrZjCJI8ZjsJG700D1baribrxlIvJt+r1bx2DuEb
GqKrqItQAogeN1ohSgFh78ckz0Bok4OO6KFyRxXXODZVqRqPTZauh5zR6ixP5vTF
`protect END_PROTECTED
