`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7/k9fxPOeoTSmKrhepfZPjaI7rFxbCw3HdSgi/DPqtf5CCj9qR6uqU+yLCzxEPE
9wKZFoDwlGNXRgfD0I39zl6iDfejmDJpRmMXfvwaIJBWT4lmKA3hNZjZ2QCy3hG/
jbspfLRGN7y/r/Eg4cqCntWPLWdeypCm2kbbYIkT+z6npYsAhbzUbwOSliIZLMjc
G3iUUMnNQdYpZ52/xr/SsTh3OYGdP3Z1qINg91IPbmvk3Kuhl/04jBmQKMlEAaFx
3XgFZPVu3+X8fLcg7zSc+n/nJhLEk8SHF65vQmTMtoaoQII/HtHC6WKjr1ZQtXVU
LshhVbCi+pDSJ60hGEECR02dnqfhMdGQeO1Bp3s4k+wmsyKE/ejHNkHKHWImCtSY
RAKYPAnENcHipW7JmpA0FjPusXDrrOIKtcL9ldhN10Pep5WZ8ZlJ2vFSmeZXRYdG
du4Bu7KZfiDkKU+Av90mkRqtyCqe+iCuiXMlhBXjfBd5++B9LRWTrh52MhjYySBz
2btKvr5XfKBUilxWImwAtVN4WOvajsylsZBuUbC/2XmOwdtw2zuIH8R/r1gtKp0e
OObEFn2oKazQZ08qMQKEP4Y38tjUS12UPYfKX4r9c8wTrgxTFZbwg6KV9rcD3fCh
UorlCTR0nawyfpysk4oTi4/CdDfb2JJ/lfJxrXQNYXZM4zzdBoAxli1z0nkuOAYE
lxAjdrHXk9fYAFIsjT4V850yi2e1ObKD4Y6JSiUOuLynkOyuqm7P2xxsbBIniGGo
EzWQCmOUTCfp4bRtg2WnQT9KMNop1zOK0l0ox+pWzfkKKcZ9LT2eMi5bJXh6ZWeZ
kfOH2wWuKoOL4xU0O4xJzwuEi2/8jqxo4BhYkP13t1XvitHzpR/pSgrjH8N+cj0f
R78ZKIFRW7cc/AtcJofit/iLJd5+Gef949AV8toReSLuegJVSoTHrcRAkGNw86tJ
kQqPBFZN61aQso1E+ku5dOhREb9/u1oL0DiNXE3y0UrILbcgMbS7kS8uvef7IYhc
BPzUu9RkoGE/7QCleEi8YxoRSA9Noaq/tVLRMtDtXu5c2r90UVKTNtqq9L8jRuiT
Sqg0UEaXLxc9ydsBVldVziQdotx1etEbpI4AVI775k/WzrSUs9xdRheojlw3i2Dw
BHADhn/vnY06iEA8hxi0MwYA0ephObYUJfCq/gs7ml3GXKYn9EKjzE7pL1jhC7rO
XjuqJxBjAXTFibAXuS7xYPndBk2Xi6ri4xR4JLC+WyInxJjuEgi72jIgooio/LKY
9No6X7FiVh9k5KdoscT0cE+t5LN4sMCCbKaK/aVRhFf64PEJFr8a0nylRzAWTSUt
SF6WxpiJkjRv7qmva+gljly7gp1IWGEKzWqykUduFI2RxS8F9SkyXZI2c9TyIFp/
euXmzS4XlQGBBDRB7aF9pRENPdXTQCNbnVTaPbThKnaxhITB4NyPAlo33234cxSN
uyUJSJPGzzEGp7ia1TdHE8Yr6Rc0X+++3bb27cXBryiWcXyrFhLRkaKOKp/8zkT3
gkKZVXAY/ooFnln8SR31A22w+dNQjGwfJj0e1B4PCzNV0GalKW+/MNku0dZhhMgD
1jJZkZ3qEMuuQzi8H/wxxr98O3+QyY3aVREoVc3JRoBpwjNmqSYnGHiPodR8OXiX
rU6qG3sF0i2FlIfXUnP4Gy98fnm3B0/FIBSrBEHJFxtzjOnansMJyb17slayDl57
ncqmCKPXlQNdjbbnbetXz531bA0Rd+A6Lm82gdeTHSa47I81mgP75NDILfcnfdot
yWQQhI9dwfXWoXAULR391nMiuXW7BtJsXdsFUDH+XL3wWEqgzK8CU+eXqxAzH/hO
udBzl8xa+P9Roe8E69jMXGpbdfOkLpH2JsrhCf5IMWnKc8AvNWxIMQmthYt9eqJg
uKO9Q1dt+45xvlF+Lf7/EcddTGPEhPyz2EN8SdzeyNYY7aivGo6ep35243WXcVPG
LYOTOyMmvTQIOHlnfOkC7ogZPhMo+DiLXyA/0n4aHbNURPbqnLsxNmEY5hIO0rC0
Yc3r/WFGU+xWmUO1MyuH4Zq/pb3RDX1TFXvFlK+PfIE6zSHWesKLScwhcMSnlzkT
FHqDimik6T+g8/HWdy4SrN8aUXvvSPM+5kzLqAZLQ2L58czo4xsckCLkoF6reciD
2tZvInVvHuXybsVAaPYmCfMQXNnGG94Z1GbTzMjKnULw6C/uLqBO0aLfbtFxjFf6
HW/w/sgutVdEQwX1Nir1n20WI/vVWBxK22KaVaw3tsR/Nd6k1clCe/VkW9/b6PZ+
BtPWWQzl8I88fuu3d2357Wnd2T6EOSMU23OC7dmxdsFBGNWWBhOGSb/0uMZiMAMs
pliGqM2CiXfJDPvDen5oOIwi8jEWKX/6zcS+GmBEsQNBHLl1pdsvbvLcybJ57aoe
ib/ytVQnwCiqkzJQCbom9Cc6P2wH0xbr+a/LXIpAMsKZtpW+pm9S+VIRVIMzHCVj
wp+wRKHUmNds9avfq8ZjE/47JVRuJiTFdmhAFfb3QugdzRnfPluugBuqjiizXKO8
xeMw9IUnsq86chiBzHVDtOvgYM2N4RQmJZLIqvdbQKzdiKZjE1rouSn9k4fpQ/Ne
OUg81mbvimzIUK1NAtRX/FMCgHlbnSuGNDQyf1D5XM5l9tVnsRy3ABC5opNr1hvf
QLY34kax9oUd1XF+uK4GyFYs5oGts4tHso4/WMwcLWv07fqY56Fq39bEg2Rp1ho7
5Pem1wzCQ7docqKhKKJVXkM+8bq1a7I1wqroCVibQWGjvcZKsOgrJvyK3NspBORW
nhjKVq5kZ4hpbKOtwYbJW60M2hrHiAMBCkU737L9JGLqSqyfLwX53zGDlWOwKGM/
x1sQAKwKFf67ChOs5wRXWXRAO1ZpGv1aIVwJaICEOiOifhYNrtEmyLkBjrSyvs7m
ocxfbCTzuQD2iEVBRBBFUmuhTQ1CboVT3dO5b/CYNOVC6O6+Wpbx23CSqhxMZdcy
QhoYNt1JPDP3x2iWqhaOUaW8lJl6HQ0e/2c9EN852pDZoFJtin7UEp1rQI5o52jv
7HnjtFDWkObzOQcFrAlKcjN7vYO0fJmXkWobpW9NirTY3h68vRdwYe4NrU7cIG9S
SY2K9Zvw80+K98199IyodJCk57oECKz1obJMsbfaAm09h6yXrkQj6pi4XYUug1xr
HuFjAetScSsMiWnOjF03dLhfLBcuUmxTzPNEFD9oUuATEhNxITfZ2OAbx9Hz6pFK
aSS12ZMRKqZL/US0Jn2+Txq3rSsnsO9XelTCH3u5nDxJ0tHSQnUrH5/+ZnPhvkBj
1YT13BPooeh6VK6+3KLMKszMzt88uD1xDhzpv/0JtmqFT2F7SaurdtRoQL5B+nie
drGgucNLcquJ7yJDBR9lPXro+yDf24YNaUDfTEEu67EuL7MA2aDeR9H79AFOMHOy
Pd0btl0YqYRPnngecq7RnXAg7FdwB4sWVZ97C4RBoRh38zlYst4dlCsBJBRhqzjc
nRMZxVxEqplfhIqryeC8sOXQE2tN2oXkzvWnyjB+idx2qKULwif/yPIG3Q4BVPkF
RmAvI4olCQsn94jHDQldsBneDvIMx3eVnqdijfKIZ5dbOQwsPwk2rIRI4uLkfcj8
8R8JJ9tHjiYdD4PnBj4O1CIJWl8n+KR0gF9EQoiwsj/FONNGHFcXiztzE80pNHPv
lCjcM1e31wxbB9naOPzXVsYd5rKKgFHt+4Frkx8azgk3JkEq/LMXd1T7ZBwgj3ji
6AQaFU15be3r7RZ8zlNIHcPO1sqYwQcPd28lwSqLDM1PVtELUyPy1IxGpz9wvtaE
C1hfWIc4vT6XCcRGIDOPce+CPK24uP7aIQqIzeGGtl+tTAcK6LsHzGOn+ngOgbA2
o0SqTIW6WQlVKUw4eGDqp9fbjglTutpuGatDJCcRSOxeXEQsVvTRPAa8QaOE+5vt
KU9LXHcFWHuFc3W5FlR4KcbtfK9tboviUQZi6ahJUE/1Isgv6gRCMvn0LvmVq3W0
aeObReA+C0ElgDG7vGJkuqRl0+Cxj3JGf4aF9/qsLzC8QiZ4W8rcZLY660ZBdAE/
MI0Ok/E+06bSyOGrYhZHzL1F0bW0dUlCw1ieNcWTawlCJbtirInvsaLTkaqaBIwK
/mr788nr4gEAZXVjMmNhFtYkJEuKX3DkvnRENVnR4fm43KwiywLBUk9bFTZ8/vWa
6LjRcKfwH/9gfvNkzqaJPaD+n8l6ZsRn5+XFBn1PlM0F9I/nyBm3VpZx5s2MjcNi
a6bjy7Rn0K+ayByAFwtckHFka/noXgDJZEGkcg4xedNr2GJAwHkHmdFy/4u0dMW6
JFfDRsGygUGWNcaCZ8xQ3hNzsjVQjuTk+RwZGpxpTi7P2c3SLXX6d2CAm4pdBVMU
HwYHoYeO5j0DVm9ULPH9TLn4lXH5Q8Ift0305jSvHgJfKlhp5QcbS1/1Zw3HI3wr
Avafpp98M6XJ7+I0VgpjyE2DcJQIKRum7GlDp2B3cRNhBA5yFwHgZ16nbbSc4tcK
dsJDzcDdOyE7RIpVq970xVUOPQo8hVDFdQxdjKkP/HhBZ3e4epQ2MZOKBUQtmiPb
xOBDQZJrqjs6VojJOPPlnJ6LNYhHrTGRv8f+4rQhgb1FjNIkOKnKIyRl6RrVpmME
NxVexMHj8ZPxy2mtRlUO7NN37BqoUnvbdeTxiV0QEZAcEr6LcwgfS3x0kwa7eADh
bsiqmHUf5iU900r8qrzbVIEMeJLzXIp1HuwAPZa7h+Rg/0sBuyta823Eay3W08sb
Nj84RtCIIP5zfbbgwGDhgYdVMwSnEf39L8KvSmUXlm/RdmlfVuUpyGb5bJQ98GA0
8LySg56E33hhhMy7CVP4GjTCH5Qr64LU1Pxi5AN91GjbLDQjQNaHTgQw+i4QYWiD
P/rWa1386qebfNnhjDiCQVA5hYsxopCQei7KCgsowqyJtyks+5CU/143LdOI4xjQ
95IRkC7E2bi1JSEJl5K9WheR5ZQlxf09oRTKxb31StiK8SEVeYPSol+KXFNt+E97
xdlea3QRPNSNCxksCUKIyk22nQx9ynQhUIBcrmb0ZBXXLXLeWIQ/GRACWF1w1K+G
KFqaoK3N6j9lRWKYi2hJMJ6Dl2qr0ywWY6gXOV1mvWWbzf2BwgTGCX2Zt4fS0K4A
7K8XTwECT3j4zLqOdb/NUNX483TR54JgQR5uPiPmbR/yugIp7Rk0EA2nNvT3z+Hs
rQNzWqQ04xgHLj523gLJh+q0fKCSw1BrvGUrnqgu9wF3azHNA9Jxa22zH5VYEbPl
Ftnb/imynQ3t0GfpzDRdIG4Tjzrm3i763VTwFdILmjItZUrEquqhOCsB1C0ggySY
zH57vTeACvOr70EcgV1kh+oY3qtDLbzLbMIuI6fYqKi2DS35u3MERAa1sQ7wFVBi
dbdtiqE/IbdKEytiPVZ06YdUVjChb95BivePRKzqauQn6hPdgvNjf1YItOgUcb8Y
BcoXbPEvR2FkEG3+GXm1zUw8ekLR9X2PcYAaebJ2rRmhoThQDnLRXXtCofJIrvGN
acvLh0m6SmsBEsEg3m9xXF5aLALxGr5M7EZsnSCsUAaqB/4lVIIDmkHYfTVnfqhn
3v3jxKkLjqzPUd58qmEJvIV1S1snOQ/v9nKxOHSK7gTp3J30GkDLA0H4+sko5Qqr
5kR+HjKTiXxtupe76cym1iVUOGUZdIHY2U9/iF9lMw32++25T6L/uBvm2kWSMk13
Y34bHFUosq/00qgR2uL4qFEM+Geolp1nPPH20Gajbrzwk5p72ydoKK37ZxNen9Zp
uCh9DRzU+wLMPbU+NF187mt6odmkO4jCZQsIJuAFxFo=
`protect END_PROTECTED
