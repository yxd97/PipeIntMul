`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJZZA0c794jpjT5jTckH+Y62CqEq5NXFzV9zTFFKmB0L5o9i9uSeWx5TsOBYe0sG
R1rz/wXA8ErfQVqkJVMQpLpI2TBNiysfU3JVNlfuO1GrXbtw5tuNLg4diS2ksdO/
a5lU6mfEGyPgnr2v4YDIscc2psaxylE7cmAXEynG6Rd2xakHzjl0EoLezQtUth5G
S0a4EAUhdpXReajrNmQjYhw5o9dbf6eXX/ff8ua9Vj//4xFRBE9LPoaH+SP1rflD
sWsG7njZkQe9kStQrVO8cJfhB32FppGL+aQcvby9/kXZAWpuyOrf2KY5LlH4K2w7
eBVjHfkUhoQhsx9zgIgkUDBSTfkJ0571JKkbmFWuHdSuSf4o9qnN4r+hY+rPgLcz
`protect END_PROTECTED
