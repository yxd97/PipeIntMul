`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXdkEpehNzByyBlkgjJdJFYiEv7Qt43B3MDhPH4SxrQdRZKUEQtzH9cnW0Klg6xp
004qIZKzUVl7tNbgDXuy73RltGf2a7c3hz/NtdRON82Z7f7BKaIxZSF1vyg9jUpU
P/pOYI0/f6mP8/U772o+SWCHIT0vayWQIsy6Tsd+rhsAOU0DjdRaLpOvWG0aKCLz
GFJcAZ7HLCyrZtR0PItaXaTc8RjKk9TA4viRrPozNkLsHJGZgP+5VUWoHD5t2ope
T8mrXf5dFMBq5i9ECtFOtcDEjOq1VyWqrKVUIC/BvQW1pcTaoIe+YSaCd+coDEte
1iUQxRW/WmvgZMuz5+eqxALGHW1DQW2NVRpQ6hOll3HLVFVm44U70bYaCj8h0mDQ
R6YBRTX0+0Vv5+VWDu8w3R5USpkbsERXYwwpZhXEfYhb+sqLCigeR/gzLyPW0zPG
d6hyOhmwfv1C6LMtyuK9Ef2qaIW+EFelUh60nPODODHPg+UuhoYxOmYsf6FM1AEW
UzbFzV+G3+IiMb/YFD4fmsaFeg+KfXN+N+fOV44KQc0CoUHKDuaNMh4YOlW+0FL2
lR1bkGSWrEPpGJscoScnWHuFOVoxQM3xCJbr7NbmlEiGmn4rAEWA7mQhCRM97IEd
t18pfjLrP7pzUT6kaAO13yBMmGbG+d+GBzHE2bbHcTetnt/Klc0vz5vJOBguHJJY
iaCW6Ji8nEM/5ONQ+LzvwK3e3cWlLad73az3FhWQ8HD9EdEz2I9kQ2cesoNJvgny
UBZHQYxbF9ACxwEPuLZuayV+r1VeHchfa5a/YsNKkmXEH3lvX1X6zRUMbUwvWLzt
i3/CBSvqvFFTAEmYgF9mLjJBG3s/rbGvyWvjoqlMp8lQNhabyvCUFXdBGI86FiCU
3yR+ZuZ4v62y/tOfklahjagMGarjogzlnvJPoJGmZP2QK5PFQP8LXxKlAvnK9J1p
/j7YZgFgdzYcU3EPtRrA89lVE0GDOgxze+3e1EaYriUt9kNouviYzcgeDJo1Vq7V
owZzO12t/HnV8VmNjeKlmKUrju4zkGSfrd9Y/WQL0FawxhXUmtsN4l3jDSP4USN7
men5zUQ0heFM+RZV57OxZXexrfDIkEE6me7CHmmFHVzCqIWRTaDwmqYNerIGEiCH
3wWxfglHsdFcwEojplGxNfi4WelFbcPuqQch2mcskPqHFeLcTfYzGS1EsT7Bp+T0
wpI4k+B9mRmBH3xLuR5J1noksC2oFJfbu3MD6FK/4ud3rVQd7RkhqIK0Kdsu3lyP
FNg+MGyyh4+FSZT+ioxmx2keV+EH8obvzp7q3aH8gEL96Ycof5SXl1uBjYAU5ESs
MUy05me5hFlXBakR1x/Bj2Gr6RB1COVptIjvjcQhu2x+uPNdspLj0Fm7Sn2CEOOn
VYN5R48P63+8rCh+vmWPct/Q1jLo/aWce4p5S3p3I6bWE2/yCRqWkCFPu1Ug2/al
OojfWjNW/OQY1FNxiHJaPMKcQ6PcQBVI4fvdIWviI588pkguhfOmJ4O3nRs9hzSA
OHv/BWFYnQNbuYtrOAG4fklVU7FghfPjZL8CbtmsatMauzH6ovErMo/61mn3M+EK
M+9WUiVGc2ljJu4hcZxEQwv+k/rgp4YMSq3LK5rCaBPtsu2S/ZYRRL+o9QW0YZGr
CVxO7+jXHOgghhT97ItnrTBg5gMTtPb3EhUG2DIinnYTf7lkfMdb+xHDgl356qLg
CEGg++Z7MG6rdHz79AewF8aAoNxgctPR4512Pl+bxueXjxR+egK1xUcKu2HfwrCK
kVZdp7cfwsuIEK4m0o2M/ICjyLSuBtqJw1XNKyXt+dr76rfVsMa2IGPWg+1YfUrr
6QqXwqSVdjv50SThlqLU+mEk8v+5NzsS+rJCrZZn7KWEWZXBQPv7k2WO6zJv4Z7e
q69HHiSSEe9tUEPPVPfguYwSTLqaUjF0WYWOU3+8rw0Cb99vPapy+y8Xw61RwdKX
CYdbNs4Sh2+NlOhGMJsuutBFk3koiCFwunFRUlLC8Lhqu8qsO3uhyLW54oEKrFnN
wpRwJBP39Gb7bhLCLY8e5+o1XsB9gKu/JwXOD9VCw2KCdyMvLzWxon66yAPqvg+F
SlUaNVQR0vPBI+smxqolmhrDd9+4niEJeAVcaT93L10VTvPCq8IlFZk6kEA7/3eD
f0TaXY5e0QuGROkcAnUXul+OZyW8jNByafpoU5Ea5CuxEuVDaPdc/M+BMG5r2K6M
gtcYxBYNI5WwR28mFdJfjyuiMvTMranm0ErbDhv+2j4vUJOYCucfktdfjmNMNEN5
RtsvaBlXA0QLouM6GpRqrDZfQzTuuN7Fy9v0p+wve43N8OuNPO1DkAR2Mq2BLgfc
tYAXIXDGdq1Gk83bnXMGYB0j2v5OniBvU5Ix7NYkmNS82+Jud5omfqzYYv9ogs99
uDss8H77a66h0m2bQkh5zukbDB16MvZiU3A2I35v1HljczoL2kjDdqol9my+XhTc
V5OaVSpfkUAWS4IJM1+g93dGs8kESpKdpZR/hnvbAfJoXPTMjO+CWHk31+bXH1eY
ahPesMGzmDA1g44ecLwrus+rLp7iSXT4RXuJcgarOtkOVvtkR0Xg8/f9JFyhbaPF
qoE8muYLVzsYoVic04Yacb/BOPWZAZQXRfbjst3pas4THlDTkhAu+tJg4Nf26tpz
V4FQa7g5QMC7W89UwQ5LGNUvRtXftudNg0NibSIFP2NBowyEyfIvGs2d+f/8bqGD
wJGLWiti0q4lhBvHEIGdN3R8OS/bjR9I4jXSq6Lfvr7sgSnAyeoNPNerteYA/kd6
Z6CJyTti9wW5bhkBfRljsq7Xj9b5yqNU5nkeg3ZKl0roSd96RHD+4fgdtIOziS6+
dWqw8s92QiFwkmc3akbKKtPETdnmDwEgZuH7afKXlWklH6lfM2o6tv3c3sB4C8HD
3j1Df0byv5wGneqd8ENyOBFdG2YvRCd0K/8cfgtHYCCaWC34ogTBvpHw9PYSz6En
ZycyWLN3RfSb0adlSF3h644HDlenPUx216D94ZTiDHPMe7Heb+7Qo8ieUOiJAZXI
yHRDxkMhFDxeqDlSgj4W6owZfa0Jy0xAgA+bgAxqXYMOjcI26r3fpo2hlnU2ARts
gtF61oZpu7Fy0hSTezEW2m/uPOaIy3dhj/CH71XDQ2fEuJLy0tIaV4wVVzTYb65q
b6VEF2KClBbDH4YjAxYvpRd0vh7cwgOYmn0ALiRznRn7LTfhTR1lqc85IChWlhk0
WOzYHu+/C42yoEB1eyV67bRiFeQ3uIGsyRUuS/oebInlpqZ4QreOU8FcXPXQq5ww
6ZCgDVP+UovFNOXKLedrnjV4E3TEE/2gxdO5eY7lv9PFQDnoCoUQb88QlBO6nRHo
0m1L6+WLTDNXIZyBXofQUOTUGpptVlPxrul1RI3Nv4VHOKBDAdOHQjw3JJswrbXv
bhfGkIBd7IZNIZHQpc//mXqAFIqJvduQ7vDiFLCzIRfSAoeOGn47zCFHKRa1wf4g
cvTq/EkDE4iz8TDUry/Y5rZjvLriOZt3V1RbWDQJ0P/h81Ov7UrCNqJwFYvcQ/yH
dHLXVpkWRv3+rIQTKhlpTAiYv59oL3uKNE9mu5/xeBSgIYm+Uj5B4fPePYcMwT4C
SikfHfKgMVT3Qy4aK0H75MSyOdh72Iq1QG6t7aPTDyssincoTNcPyBZQqj1+wRB2
yzC8xyGbSb8WFLI+Ja+Lvlxpjq1+MpO9Xz1spgVaeML9LnM7L/XkJa55BsRCORRD
E7Qc7/Mqybd9m4fHk8i4clnzQPHgVxNKLo3Q0rKvWHYaoeDpHj3FeBy5UO3tdLMw
ImQpoCW081q7jydfEwehVhpc16tO0R1GYHfvYxWdRp7PjAcx+WOyLBZ5ZBFLPGsj
Z6WBbvDraKOENFFBcRxbHu9d50TRy1/1yGnEnbtYirJ8cQuWeJlTHO8G2wh/nZze
xha1TSllSNH/xiMUy1ss0W1P6BNh/X0NcoaTtfS9rl5oo8oorhFz2jDG/sSL82W+
0MytiPwaIEljTgGGNImxJ00f7QpcjRpnWQwPhq1nLUFOyngAlfz5+4o16RdoRAyZ
R1XyKP6hopW+AtkrwdPsLYdbMMBgvjqHtkOHJjUuSZK7oqIg+FJTyaiNl7Sx/W5+
i8EbnXKkXAj/rocuBv2wW5jL/HW5kDC5cxKcdBf/yYEKAtDTEuQMFJh6inLCn2/m
3ocVF8spKnaJ6ozGQfPZCxzMxF0V4/noTOdvGz5/U9C7fIRATxvmpAHymzDH7S4f
kMI6WpDyFFQ0KFdDwSp720eexMu1A6EY+kVUzkfO/RT423JCNmSXAI3Quljqd6nh
5nyxBPG+zOf/HWDCjEX2xRnsEkhO8nH18bnSgfuiiVvot5sWrZSasuuaOYCRYdkL
FFF9fbXyz8csIAE7fo35nDjLxkXSFfF0SpGpoISlvke+kXNmvOxrnDdPyq085nIU
uwGUCWJc3oT0D4LNL6RbH6tfuS8j9pmgl4+grAEBJ0SqM1zWDeevPUb/+bsQo5Yd
xoZOPIeD+U8aJQIiPBmf5D/51P7lWxXXc60jJE6MvWVvkFdC1JoVdglGkBAJQZM5
oboJHO//8eThwL6u6RR2piLvOyTsqXlyy+E4o0/1AcF7OerTd6a0SJrfEIk/IUo8
nhWZjaAfB2cqnf0i38kG7nQRtT1BdBK3McE07w1mZ2FLMdygGsnpxqIXJkGH2wRD
xV4vkDVO4VfNTmpkDnqD98ZqcJm/i7dzYKEb41oAE06qgwauV8gQt56Uh0MKkl6M
8gfocmGhpCPZCq8ZSInJHHVX9/RVJCjPVQPcWMSilpQpkzpaFRXPYFP8Xrjj5dB/
FSqRwagPRgHTfHtqR29yFOzp/SWIDL5sI7nRMuWvFojMaD/sPoMdqzYo3z4K6JWm
SUNAHGuT2lltyvmbT56Vs5OZ0h2FbS97uKWWqKAOGmiiTLGX2uFs9e+VANIzJwJK
CX8mJ0pVPviRqWOwocy/O/y8bFSVSXw9EpcqgXHeQDG8cgFMQgOo8xF4QBYz5yVf
Hri66lRO7BZC79eT+PDQRgLGBhkOXVzXOI8JCi1UHgBt9Kue1v5lCVyqyMyS/pgI
FgBGOWyoMjA7KsgasqMXSJHAuwaziwB07FYFZ+NSF+92fDBNnnD33bx20w1kNboB
T3AXTdG2d17GXZkCW0U01fiCgH/cJsgRWEIKS0rGQGy0GWSz587JUabFl9qQ3KBN
c3+qjXe7xcYhXNZmuKyIoDL+Akjf6+Z0lOPbvoY8CUwWFRwIZ+EOqZ/aeEqe2NVB
l8pXx87s5q3g7FdHsQXhfxdCqsh3OQQ3u0vUffxH5n/+GrAxe1larA0hrDQEXXuv
XGwpBBwnLke7hPg7VXAOQKK/kokYZBl58a9Bn9RmChQaKywQ3C+OhGFosIsZ7u3r
UcqPBXDGekEujiVAaZPiqCeoA5GXD8jSowFXX5NnVAriEOk5lIlhAWAGosKfv8sB
5ORJ5n/d6DekBqAmDl2QKiqyccTlCG3nm+UHp1J6+6DJ6DxCL3i9OvlhrXI+KH6z
eFf3keySvBWrxMheQsOWWqO8zx5Dz0vL62tcSVGgM7NCJE2dzaGIpUt8GftmKslq
aVuommWqGF9RbgxwLA3cjYLQdevOunO7v7dleMvsvcaXll7Zxv8AFlQV4h6GCGRR
QvFb8jzo2ZZ81vw+Pq2nadPxb6Z97sAvLIXWzAxyAxxAnSDmnZnuq0+jVjV+SN36
gcBvllWThOOgvsjGc1UZsq3FLn08IVp/4l4HY+ofhWfG8pRUzpPfuwz/PDHCR9n+
Vyaae4FEmxiQ2gfmSGz3i2BlMmv52/kdSaxfa88Iy4Bs+2R1yqkj5/HB3zIdWhL1
MPkDqFuE9UJdQE+J/vGh8V6/eFJwHetbW26BNf/MrUzGkNWFcGE34QhjfmkZmb1V
q410zqK/QR3gNVGv/scOB+rpcMqY9ORhjRkBqF+QhhiCkjanWx1K/4xHbFSh4sKW
m6j1WJJCd3EOd7VA8iNsiGc68A3U+uUtCcS62q+/aWJ9xpAKJ1hHifs9TEAwGYv7
b2CP5T2P7nqUPj8fTBMQ9Z0KUJ9mmaM52MYO6wbpvK27+LtO+lPWJqqK/PTDY7nY
5hloVKva1Rv7yizGix+OKmprXWTy+XIXTZSLgvQI+Vvhb6fNeKeBp8+Z4EiF8W/6
/d9czjXWXWX4fQqzRsiBktVLb9UBI7OvAShah9wxOe4xjh8KGGyseQXyUePsUU9z
Ddh9qKIVodgQU/yGUnm0/gVbCBFMuye00Oq7YMJ6l96BN8uCQ6FnMtlTxIPrn2f0
ZOO5kSrHl9OnGxHVK+mJnnhEHoRxZmKJJdBP960WEQhk9Sobtxh0/NjwsOAVSV5T
a2Vu/vv+9vbDSMycbF/IlSEiQfqzv1v8Xtu1leQOSWnhht7KxuLXRq5IALCxzYvl
qPuUJr/JsZZXURjjrG5oEn6uufGGHyTcZKQZ4hLv24slInnnW/Llpu0FevIp5V1j
4Jd9nlhE2qpBvZhJ8frxGkomKiuwp0BeQEMneIh9f3BjqTmNXoGTclWy9s/+0Udm
9V6okjkHy3sVDCajpJoHO/fp2Ifv32C48hDVYVt6sHmF8VrIRYlzQ31fbJv2vNrX
SmU4nM7OLcCpAzXz8H20yIru5JngZZIGWXoQplEJXz66lROwY7/YDc1pyTl0xWzO
BWIdAkuOQDVJ/dSx0/vvwPnbfBw9FgkEI1l2h3/Zs82lmO4mRmAtuXWNMnPaLaf4
HgFBeDcior4dhl0KEPxp48OT97IQ4KkcyoShlOgWWIy+XS9yb/peF4dTOZu9wA3w
MSOGX1zNCZ12bPpk5/ByiGkVvSuRVMPCaVjGh7FVlJaW/DReFQp8fyjx9bVy7LC6
JxQj40NqGG75ypzxydcLhP9cX6VzLhwGqXHAzPLnRj1PfvAZ1HAOO75pDk1h2l0D
qvIrVQUQUmLpKhCpkiGs8naKHbZF0JGXXHVh/wOTTeNF/rO/Cx+76WYaRsAfSs8x
diw5GIGukjL7ZpNeUYYkPsBE8JDMuYR03va80Koa0NwS4tmRERq75cUIsg//Okqu
/00WRb2ZWCz2fiU2iTQgWyWy0/UKJYlnyCvmIt4Wj1YIkXHHEz77mQQhLDUGutO8
baVWhvGlqjGIyK+RtsJxNRccYzucsIEaW4DUGgr/CiNu1peqZKuouydf2IJ9vBhP
jT7h3QWgNDc+RDtrza/tDWMVqUGuP4z2brpPtsa371b5VgLIFNsRUlxin3zUQ2rs
2ljpHJ69PGTvzggywasMql6Enx3DbpYnzuGVWPa5P6CIHQcftzVDkBpf5HZL9hiI
mckoM0woZs+jBzyqZgGiwAxwZcQgSPuD8ihuP+qhXvP6qi22hIWckfB52hSzY6uP
F5ovlixJPQkVJzoUzd6wRFpztvdUUXld2unXcAAXqeKreNo0+7UH4CMVUZ0bQzOp
lvYmsrq8zV+vi71VKECYzCkAei7ZvbI2Ly9meW6oW6zyLf0o6UPpE5CxlvpGtbxU
S0UOWD/DpS+Y/7wK7XJvAVoV7Ea5nbVZymWPm2jO3O2I/8B5EiS4VTZrYbMDYlSv
BquYM8aUemHpcvqmTDkDIOPU0n6s/N2MgzbEXFazw3hkEkt3b8bynO9K2C8QhWo5
N4l745gl33+NALfcC5Qoz6VeQIHHgi05aAuksspHUUaqTrb+CyYNJ3oz104Sg4Pf
hE5bSmVXRzzDIF7qi6rN9vHT0FeB1i2dssq+oJjJFlJNrmm0du61uuqj3pYIm4OU
ZbHI67r+FoC4/7+EYvXEpnVCPhMFbikwtlqIa6FtMZINn2uG1GwydK11bI7eQWqg
jXyHSP00SfTfR7ZCOIZhmWnspvU7puv3NuFasM3taHcVpYNpNtKUSpknBESs9kMR
WW6bf7GJrJryNqel3t+qDb+1HNk4FWFklMC0xuZVp0PNoPU0tUe7ZAoI24aETPCK
BGxfV6ubJ16AE5jDJjSTO9uYMeft7F3PyKVFLPXwtVNEIkLyb331jNHxM72INw1S
4Uu3jMT/JO2/QoSCISZdo1+UXPe1sMNMymw4V6zQJn+EKIIlMV7gafcugOcpWqpu
pM/x2Hafqujt14PzIjTUKzBNtW5oqAFqp91P2sOoAV+QK2iVJJ6IWscuhAWr0t2m
t9RNFJvgk2Rxhc2e0NPemv6Eri6sWGePkJy43RiuKNt1UI919eo3KvjgKdObgcyI
tPAFZUaJ6Y3qDF6ZOZIk4JMYEXH6rCes3QaMMzWja58S1lE5lMXC81VMEqtdaCwp
v2/luP+zFzXZZv0McOeos8L1k8zJ5qxJdgmsbL5xEn0DMavQ2TMwH6wWPywqZUwT
yRqezHkzfNHBxyKuCGAPjDdaSFayD/ZufJDSZIaOFzsADxhuVrNisUi8jr+9RmZx
yUTayRD5HcZfrwMJAN61FAjpQGvxVf4AbQWL+yQKgih05A/pgPBjz3HEXmTHZiZs
1wl90+EtBsZetRqfTt4f8sA4EV66GiLczSHB4ffk6Pa6j8Ags35r8U9NBQceJy5p
eA8BB+OSfBK0T49Ab5rthc6DlV9r8/FZ1rqE5BZQHdX6kRFQRVA/X06EuGJ7o5du
DAd1bnOenmOMaCgXXn/l1QJtG+Dqs6yck9AaE0JsK3kFWNfHmDdrw7GaQsgAqo8g
0/vvJQV3CxbWYmrFJ/+7RdyJ9zv2/93Zlquph/pStjrguOBys/RbDd2gTwZUUU3k
mCmZRHiUC1SOc0J8ODcW7EeiPL0ECGDYHYO3of0QanoV29+MsuYXbmV7IYh1Dr/7
zCX/zvtNrCldHZAd4/aI0VAay+iHHgrn/b8tVunXE7ijJoxmbMoZCFwdULUnHGA6
hXxJ5eYDax/TVuW5kat3PHlmi3/Ja+oxgC7v5MnTq4G33+ll68GzaUtMF2K7g767
atHCognmf3VYf7B53zrxERQWwDcYXH545b8lkrTYFS9Gbpo6VFbUw56xxVveAXOl
TmLO6TrTT1rpmDVmqnaJVFVX9QJCejHxDw5vXHOM43tnZijC8nr+a+g0BH693Ah4
7PFbrji1+PmKfznd+7XvyzZPBsQATSKQ1pELpo4n6mSdFTYZYya51IEFcfRhlQst
r7ZlYo7ViE9xzXF/vem+bNSd16gQfRj39kda1c8qCZqXd9kKb/2mktw90xkG3dc9
Pgp0KK/lMnArU2v4LUaY3xtVGH4In35fhBZ0Bw33Hw7cRSxk2OyXYrkoo+TZdSvF
P46CLx6aqle+z22laBLPKHELzACLUi73ZPEvvEWXgQndP4owUZHJ3oXkkiipU/Ev
PUmfkJF++X10csaVeB+1sJLswLiTc2gDv41F21WNF3lV46obpTrxWjmlPdNLyk4f
AOvGbw9wEawSEGRgOi82JtPx2qznmiphyc8dplDY/pZzHXW/orrXX7JGn/XBRUqN
NDeiDq8iUgYvSTj0FwULF25qTAguZoGRcrltYuZ9NJyfk2OvhH5EtN3HmoMYzXqI
zzecrEFduIw9niACib0JwS+ZRI7Mh4SjMq7OdhoyB6Fczn3jA9m3wqMSYslw/gJ3
eucn5IL4Z4YV+bd2WVz0LAIssFnIAe6Em6pJl6tfDXNgF21wmRToYgcfuOJ/F93c
AjZicURPJvcGWjU+bn+33UkTZHxWMyNwDShxLKvOpJ87GAs+kSaEgawXcf7uGbt9
eF+v3rM122V1P9Z5Lz2vk9Pi6FPNv6NVGQg6nuxf+0nhZ3cFV9FtcOnqdkcU0zcr
/r4J3Gu0EfFB+2q/Jrq6Kx6XTT5AJH2Z8vqgizZuPQ829agmsIH4w1bjZfiBkQHf
Dh2gxwWCPlANAzJLKfAq8jJo8Z3CHLQQdxdjerLL9isKuPTNptLxmjldENY1zLch
/V7+3E0DnoT/yuhGf/EsxGTWSh5t2yaczYNZ1eVYIhrA9Ditc7Qde7hPGTYwRC4M
V6DWWHD0kP7sYUSlxm2XzRLC9Bbru+fVACeFJmWqn1B/CkiaQoQKApnSyAcrWQzx
RwxrdJ6GDcoVn8ohxj1QR3W+xHqZGV2R4HceiM72QcxOhPdqFWB3SUVBSvX8pbsE
LPCTt6NWdDXSEjnZk81okD8hFY03RhGg51/C2kJGueUWAULiDpMJiNXLPDM7pd31
fmFKCNWTU0I3eORx3RYCNIsWzMjGpokuv5GnKIGS50YyHY2mrAFXw8DkFIna2mIo
pqvP/lGFpYB+LpVckTz57Sjz89FA4QUXUSuZ6HaTgsPmTaMM5zQCpojO5EDy+mF7
6OQbEicceu0tXZWUY9bELt+FUbzxax4b1DkG0YLi+Tm4a2vsfXhuJGMW4gnSOeJq
8CJiK5BuM/CNzE2kazGRRv8oV14iiyJ9Y2zW18Jd9hxM+Ic1Ndz6JPBKat8V6/Jw
jSkfhuSqEgsmT5Iqnz5uwIf2X/fH95SzdxfuqMPbumGeznsUo5wluiN257uqHcNz
HQZcK0H9M9b6ydplFLbBhtJIk1fIxtGSc5aMXfrE4tAy4ttEsMige6LJua7k8oii
dll1QhsJGDND42N6/TZz9U7572QUS5N0wY2O1MlOHwI5wWcVowbK8LPVdhWpNkR0
jx/Y+xYa79rTMlQw41OixNUxBrlBitPYjSDkQUvXvWhSs/YILrzXMPPcLwRunc/f
YQLxEgAgVYJrjM5teGRgXF3efHuBSZ1N+KuaysTFmfNlwa+SiJZyX3kcRxx4GkOv
UafL3JK19GZP7/W3z4CtNqIo080iOhYlhnKMgguY/E/sWGYXyAGxnsVSsufbzzwe
6VDqUctEKilLvuORYTgIbFaQE6wJs3R6eKHKa15OaU9UsZAC6YZWZW9ZVvS6o33Q
QFAIB1m8mJBELh1kUCpcnwKM9fDAmIsFIua72jBWXAPXv7BGcbfaDoqZCiy/NOQx
zcBgqWyc39vGnMZI4If8Hv9o6GSW87owCgm02f2d/LMmFElF1cS2z1MgQLKjr5Ng
T72kRvpeLZha55tYDj1kz76hYtMaFGZCewtJ+RSZnH2WD+A4BFVeAnL67nWdKajO
JKqYx0wL8MOSPdip7eS4YB+FwEjAT3ZfI6wY8CsBxSIIpShXk6LFAhuEidsQs8Cp
RQKDk7BAFqp0i7HFxKmQfbnJngYqW4hSL8pPwCgEvlWPtveIICwIOnBAiVxkpt7C
hKxu0xOmt1AOxJf1oA7LUgH0re294rdMn9IFQFA4j03cl5tjnI58isZ6MVS02V9B
4SYW7NME9YUCCcLAUMcxTAPev4mtkcl85bF9EHa+CVf/E4H03XInmkj0r92hzLME
yo8Poxif2k/dIXsYv45fEzl/CvkiqcijQcgsSoLwX2FYFymhrQmbnKUUzUL9/EVt
ehdrC3ewC0YRqGx7HbHAIk0QtqP17wz8Tk9R70nTbLs103fVupkehdkIhJ6Wtcs5
grma/iFQBYsUdl/R8jt4mPgZvpeqD+oxKPtog7YOzAeBHDgSz3T7kVxkfPc11QXO
eINsEMUrRYRIBHPN53cdA8Nu+/HSdCbuUAF58YP/MfXC5iDPWknRSxp6SwdzS1Ux
qZemaxipltfvmY+IrMoH8X725kXpvjbmo1eBfX6Ns1VknhbV8eLShYUm7jdNcUp9
GdxphzkRj+9Yhria1sm/oU+DbBvWIBxg4QV+sistfwtbproV3jCmyi5hNlzWCQdn
RyRmTPWnxogCOnNjKDIzvmhB3pKFaZNTmYNvbPNkyrxVQyPqRtpNdw7D+3b3g5Nj
XKpr9a74Flenun07aDcNAgrSdh1Et+TzloRjy2d09X1ERRjzdo+zgQkEWLpvcsds
6f5BV7GdFO4yPh+VNI7zYAms9HKRHVr6hfGeCY0vp42KmA/bZA5E8GK/Bgrx+VOQ
q0VP0HjBc+q06Y8wxbiORKyjnyMHlRZ2zwbQH761Xq89lsuPpoirZKDzeH5hwtHy
EQOCv4Pz8F1PQsdrTz4FDRP59mp4+E4jYESAdyIGlgfOiVVbiXc52tkkX3tJVgeE
iX9Esmej+kGO5fUQp6aHN1HpyfRhUSjezSjcw/ndiR0W4eVwBRFX1RA/CVMfTdx4
u5yMolI+TX1ag/iPaRyXOhGGaC7lM02piVK1+c1xLk9UBirbkWUYJbPjhmB2yX7n
O7RMO5FU0nq+Ow3Ze8NwEvk9QDmq/KSVn0TGfSVPnAJ/lCKA+TmxiX8IM8UzMbxf
K4JvOkZQ6eJr5AkmDLYyPhM/G1meIevtdHjkaH6lkBROD0GWk3Knm+FOYB8suPBr
23vhVEK4yaP1zQy/kkmiFJ75rgcWWDXNXKSF0+s6XGd8SjJSquQeyG6zI+iDOkhS
R+ZK70Pcfo30SbimEub6BkrQrki6AQ0WPA9o8Si89A3UMESlU555sMGH+DC02yip
fZEGsbUhdW+hmnFylYur0QFpyjXYcoyW0BEbKV05fLIoY+hcN90hIBtGRCHv7J++
+myvPW+8PYwglX7Ir7yLQvg5ha6Tdb3HSfu3TF3s6AHAgjxi/tB0sIi1b+aztk+4
YEFjJJ1hz4KN5nXCtbCDOCUPSs41QfAokMYK8awoW4UMiiPgXbOJcT9JdlDn/MGs
PvgOUkumxH5X5BpdceO5NBzlAndq7DE8cJwJvZD+UIuE1KUaK6TteW6vWXgcj2qO
zs3byY2+LJaft4IB6+RNYMbE6u1KzU8Y2b3e8RkZVgUj4ppxU84IYfje1lWBs7lw
x/JQlWhT7NqTZqK1QVyFom5QNly8A6yKZaKQhJotRmBYbSUoa482zIA2wPf5hHlx
Go6yJo2f85VV5A870LYsWFNzR9glokgJOF6PhukUssbmgPl+qWAoSs4D/+5DVSy5
DPu6HTiKHO0Vy0OYtou4lfDftgA1xJm/oYj5lnt6KLYY9rsNAu5cFGa0667YVjC8
oSz/F40z7sGCFem67A8XGLKloz+aSAtmMPHwtb4iZjxGirRjQgc2EMRv2Poul2OE
1IGGmSH2D5OlOv4puM/iJTaaJt1i9zkv5eTXiOUtB6PMcICjWTduT6MiOiHgo/DY
yXzULNaAdh216s/moNDbVDvIJ12hPP5qcgX7JO6K1X3oqGGsZ4AquhITZWys+Lyp
aD8oCX29sU33kIaevu5Jd16y8OrzmZo7A95DhQJPRSnFU5fnjkn+lvfJYyE32kZB
7N4GoEUDP02pKWXPUuZdnYlDUDr/HiPOoS7gYVpkeIKR512WCCJe8WeV6Hez0Gjy
MQJfm8peXUqPWpY9PPnYR+Fqgi/pGKZC/P3AbqUEmOd8IcbOiu5+h3fqq/Zn6Vw4
yEvHIFFXuOhz9OPYb/nFgM/6n3kGk+fkyYhg6x6Ss7fvhlWT4vElyWYa+2+DaaQT
I6IbdY6eKGVl48a+DR3ZxIRBX6VYdGM2hQZJFg+7g+B77PVJyH4tlO3qNRZI/r/W
0Pm9cUIMY+E25/rJBFG5sn/41X08PWk8i+NbccmFXNPpWoxuzHpPC5W4w7NLRdxE
8LJciDwj2vCDFC93h2IoQeqBmPN2YouBwvM0r42M3V6akzRVmY8nRMbJp5rAiqBq
mWyA8X0u9UHuoczjQqHg2SUsAYHYVnHXusWk/b24/mVCJsZPn+jRbVmnF8AuMJGY
Hxe3MRN86SgG7yTivGDSt7Y9yvpi1KeScM5uJl1nZlrAOAQKUoD3nim0Dxan1kYx
DIMI5E9Id4o46bdsuc5SsFCt4iqtC1cleFz6QNppaB1psuTUo/Axbz+BDm5dFWtz
YwOIT6OnKtROEtHEx6tZQXg7/Oe2N8ehTmlNabKl2jSHEGlEZgzHws1wnUMH5RN+
bQ6W2Yoa2EPvXlexYuY6RvYf5Wx8Ou/KKTdQMHEAGxuSSZULuW8JDCzPCUVNwvQ8
jLF/i9q+upPGJwbI9ias/FgmGuC5VcyHnyQxujUx7fpMi3O6MUL7iJdd7fJQQdDZ
NcPX+buulEQIP8kSeiKoRJNdd7lFTV3VDhtM8qq8UgMx4mP6KxdI/vCiWfRzArKr
4pVeymBRzPC4T3ceZzOMnmBAz6+HzRpKlJYO2hhm4mLpTyNKLPUqZhSueki1chf0
T0l71it/gEFjAmnZy4PViwp8OEWqXKYY2sR76slrp/IE0KfbTdjnZ60Qj+1xRckd
DxXu1HNn2Efu4Ca6TkFmDCaWOm9E4shkmN16xEXn1FGkRCvKeSvXwHVKGW9YREsu
3Z1mYsdlQ6UdMKM/I8B1jx42K65TRZFHiEFInM2bj9YX4PfwN+tGhkdHm9/k/1n3
uhmjlgPsCMt+d53lkOoFEPU+nEnUzZPlD/PuZXjKEo3wPDbVJZgAR0Aib8U5bX75
55wNtHwcHhyjLBC6LyEMEv5/xODx4qF5LfwMNNuqZLaGTXE3rcLor4stDJsXAhZN
9I6Lh0WgJ4fxTTtkFM26v9A4VmBSgL9qJjWaLyBswJV04s0Pfuai4P6jGbQo6x70
uLiass7oqa65BlaJWkNFFaqt4KCZpl/yrKhBx82KzenSe+sO4f2mQmThHfTNpicH
LGdaDvfaIQ+oH75mo5wF8pMXd7E51aryfIjP1zVdoKqIf3Z/0ejh+np9OSFxdOx4
ke/W9XTBagCzdBi4ed6Esiwk5GM10dJmrxWnF1QMag9yW5jgVanlnqgt4020QYf0
nFdxS5iUn0b4o1JEHYIVSh5EMBG19yFLUQJFDwl6+ShfEYEyeRnMHqbzRbYLyZJ2
SCgqt07ZbeyzoV/gBAAr8tS1ZnmTCEXTf7BrhTZiWiPsqqrmPXssZxRe3XyK1rPL
u1Aig/nEU/fUGn+FDxiwxYPWkRdKX20956FmF21RokmsOcfGDelmOoGjp7x7hy7h
dXzrnLn+q11fYcIFmRZpVOQl94Y59J6p4zxUnuhRxEfGmtxauZuKnJMPbzwTRZCr
vJekt2wqXhTB7ndAL23Sd6ytGZ4dQBo9lBzHCvSqCEPWnuPOhItnzXNbnB9fr2PW
xuZC6HpBgGJfVhcoVe8CCkQl/hWxw2RKaYU0crwHSPTyMPQVbpMTnhY5qFAmiH35
RH7bP1hqmItKlbeArxMHf+utm13EPzLvBhwucbf1V1pGQPhw+a2Z1++cD/YkAQ4Q
x4PxMkSqMCynSwJB9aw9agis24scig14c9GcKosiCvjDpslrA5wq6K1J8ebPbEE4
sq0FF+UQN0P9zlvI0jXSfNMvLUXqDavCUkrdpXNCc5lMxHtf6J0eHEx6p8cJsup+
+g7LPVZPVcyLRehrEcKDx2I20CoVkAxzSNXDS9m3rnAJCR9ck3vTDvDWoj57rHWR
QaiGD+tq9yAjDmSLM0uE5jp+t0VyAnUex+b56AniXjXxMH8CE5gGTuCYrIDSCem4
lcCCBPRDTOuneIw+EHg5LElqoHTVhhPi2ugz31H7Q1741xxN+U83wwTGlaWptNJt
JEh4l2/L56GXr58mgCxdj/EIt0sTDG9IZWUVY7If3w+hrQSCMq6MLTCvthWU4pRi
V3bh6NlNYwf3po8ct8gdUyYpO+rmRxoqsQ1v7H3T6HR0zfka11h7JAyeuUo0ixDb
UqYXSW5LlOxWdzbQbutbAnMvRm0zxbnL65qTKvreuc/o+w74iSscvjsuJUyRkNJ1
1Nb45mM4ceOiiEJ4m8KJTwQ0mRKjLI0FOZtLcXwvrxF8VEGVJf+XLAdbxpsg/tUt
niRl1WI9HCakpVuX2OiyiRBVIQyYmcE5kFsjZuH2O2QWKEdTL3RRDbYE2QTaC+3I
lSO91cAt0rx3w84/MRf9TrrCiTspA0m1i0EGoSTJc0kapKy5ThPSszwnEzcpSYq+
tpUbnESdPyXvr/Q52oJPWsAlxFR/K1Mn76Ct4fiMdunXNd/h1w9HF9Qj7lWyqRzu
2nRYuLhkUUSm+VXXD6A4yiA9acFJbxTxy72890TCO+x4hW8O8iIFGUdYn4yUVsCO
nH5jsEKIfeudHAnziWs5q0nY6kJAboHLNQTQNe12/mXYGMVov5XUVOp8r9t4rPMj
boF8QeCE1aCpDJ7+WNv5XTYw7GJkVep4EwSK51ZtGDqYGYR2A2f/c9hOBmSRaUfz
nm2MqnBgGRyHtLtPtP/6v9jeKdc/qHv8/dKLAIfvKhlbVev4doeeFg1b/ctnlXav
4oZgb2wLZlWAXSlqAS8rBrqHmIpxuExHjqPZGfY9zJVbWywKCEhHRvr8v6jPkP1g
xzDWVeBpRtrKg4jJuw3W4V9Evket1WVwNZ3yPqw6iVCM4+1osVdxjvXUOeGrMmSG
KtbJV3lg50e1VH7I9G4XeWoFTJDmNwS7luCMdAE4s3bg6Q4H0L034fdJIbPanoDv
IoyBf+QhXnH+Mb2tVknFAsuitfHs/Avk7KfOFky9YhRNYQ0h3iaoWQ1B/ghApGfM
nTIXrfsIUtLPE+1C6vHkyMO+9OY2Cdbesj3X91ePJPfHfuAt+t512aPX6m4u9WRR
j9s08MhNKDitGwYFsttXTQjhslyuzA8mYtyJaeDcL5z9h7n9OBojecwG0BHD/Ygg
+phViuWzUpE5RuBQe4YRiv7ilnPUJCT25KfGkivhmK+M3rW+UyOc1mcsDBxoqVJn
C+IAodVW6rsp34e/bP6+lL8Q54vsGFCMd9mhjg8jVsfR9+g4szSm4P+Pm/JCDtuU
bRf4yNy7IFjofAmOdhC0wZhpE7xP2lEEWy96MetFPstaB9HWsB2nPNF3OrVpaKwR
qhU/AmWM/FZAb/T/MqZr80LdoIGkpbjk8/Wa1wxjwFRsP1yjx/MN24kfef5csvwB
bM4ySo13yHcJOT/V70XSCI3j+yCjTWncNm5aTm2SkR+55zr4bIkceVLGAc6ozSji
3MhD7ngGjr4BgYHXwpYJupQ3oUYwYvaKxnzByO6DScZg933obR2qxCVIr7bv3EeV
xwjFD07QWhDabNijBqm33/iuv3vnetC8GcOcqDDH/XIIEKLt/V1/ezhWzjluIpsM
IlmmoPXIIhXU3/XI4L7JxJNdKJSDXBjheNYNBezCSSbLEKW7i5WKeO9Xpj9UcwA0
cTqmowSNVlvGYivsifdHpnoYDPYWhhvsa4JNYXabtsHfbsMvbh5aXlOz9QogsEPz
mm2HjY8mmJ6M0A6+L6RW7xo3VE6P2ps56e4+bNFrc2F34XFKxdvBDmv76cVk/r4J
X5x3ph88MYSPIefsa8qai3RGZM8ADGsShK6L4lOU85KHFJ+wHdze49n3iyFaJH8w
6kRwU+r/TTQ0cl+9p2kel+q5W2HggsF4gcyNjadrVccLhWfA+zIDlLVrdpD0Ulxz
BBPc6s1cCNOkJFVR53+q0rqRTzCKhT2QEdvT0jvOnYnd8OYbbjs0tGmM7s2+qKoc
zVplFwhUr/tInqve7A+iI1NpzUPi9leI+iGV+pGfERyHsbU/I6Zi2oBEKNE74cQV
le+x+jWBhf6OwUYTqv1GfIYy4foRg44rGso9S7aRTL/MzBQirNYvbG3ACu27aJVN
ufwtgn8FDcz/88so7Mtd9mxJg2kBLkF5RazEpobINnDKE8qkI08b2I5w1wpWImBk
zUNRuxC8nq2JY5sBfindMXVXgm+qsRP9kzQPV2u/ZoiuZFyhQQ/943l41wFo6bPV
VqwdFIUvtCyArfCNrBKG4U3xjZdDGfjKQIF1qVPlvebDrRxDM9m/E92O+QwmKR5M
qlfGPsYnwEQqdvPPXlvkNVO0kxBbKPAodCdUZVbqxHrflte2ECNnjvVjM+gigHCV
+kO0p2vLQ3YZsaw4a3NE4KAJPrng6e3cC18tF2W4LA55Y0y+uoVvE4YappEMScMh
GnIG8Ji+dM971Vy44O/VIIacSS/Gfce6AqKY6goUCKUtmI9/jyELb0ZQOgr7vm99
J7nGdwFA7xtwjOq3Hwz3U8kTESH05t94iJMR16DrHBoUcjT7sU7D9V19Fzoib3zp
fLDjl94KrM4GTPhWK3qb7tPMKGO791nKmyMD8dAcDtNDTWS4J3C1MSq4C+EXiUB7
wGHWTgh9A4rIoSggMLWWN19eljvNoI5YQIWOYqggsyaqJOB03opm9yVVDuxsBalg
OCmsgTQs5W1P1RVpKY2shUa7L8X3G/RZMfovVUPf2+EwNz6Cx22Wz1agVD0DNMZH
Ln4rLuHOHTlWCRwDwMmqXrJRs5Zh+WT4AtDuucfMzT4HGjjnjk/OlizhV5wMmFSQ
86hOw/BkdrOy+Xb0h+R4Bs6qyfBLovqMpqLinbxUc9h9sgwqbPPDcAFid1lKv4SY
71+/0zy/1kIQ2UtRLBHxUhIHmtxmogTmbVkdyUG6OWH66MXEvr5bMjKmG/SmmObH
LHh3/AoflV+jMo0kAqHPWyx5C1zGgcodDwlxipoLkJEmryRXqfCkAI6yoTdpMH9s
4S/h8a+w/OZSGx5ju7mBJVue6m5ORJK/Oe5khTG2BafwIA+ducpmKaOYFxHIYWr8
1nNLtHb7jrZo4OIpnn7++36xbAi+qqiOpGM95/3A5y2vEcJMRWWPom/W8HaN5nJn
qFPIKMolaK9OVPjdq0KdrhC1oJQJbam9Pd/wNQBmFSx5Nrp5CZbYz7+UwXXvcmn1
VB1R0KBsbhj75moAfmM6DFm1xw4uoN9ZnEzrib4822Q8aEq7hP7N9+KFMevOlrM6
XCv7Q7Lx4cFfLko83Um7pt2uPXEUlpRniLTQHJLPWE7FFhM3PJYIJ7pgJR/jC4V1
06TZRNmaWWrZaqzl1Hx6NRvEcj2dcwyjSUjgyk9i7MqJLUSMacDBNizPxOzIwawW
COUep0CA3GUMWt2AOj6/9lYTcrG1DGON8Qw5VFR6O15/VOXzfKGbVrQW+UyH5l2e
DCMvgXhchaNA6D4+aJWhOfzRhZjarYaon09R4uvqFu+Aast2cvYf0HpQpeBHWBEt
V1fHuHTT2wjy4AzA+CH9obxZiP3Ie362vyUsZ/fyeJjkDNFagT+snhYEBeN33WHR
S8IQGb98EPkPua7cF8M8batjCaLgYq+REFAXQn7iDrmHB1xkOPtxIDIC0MzcGXMi
yvh2w/RJoh08xjkqnhBCdx4SBTDvhRX9w3e3VwtaCDgffuiW8fWWqVSd5f7p6nDe
81IPhLD2mJ2jgy5hfvV2fnf2LYpXt/Puel8gxxGB22+bPJCpeC/QCYDby0+NaW7a
bav7ItlF6nA+Fx0DxkTfxSp5O2eEdqm2TXoyPDe36tk9z4XCyTJR1J1CIU+Cc0Od
cNBwN/1wF6aN6RbM8uCoxL5qAl7u3Ebpv4R/s2VZw+wS/suarYDdtwYAutk0VZ2p
uN9ceHKEUbum9slWht58vmO3hJEsMLanUGhT+PLmVRvNCrUItDktwDytsiGjMn4G
W32QOv3urqmTYKFiUYEDgTh5Qr4ERFEkKyrjc0eOJF7FNW59aO4qMJA1O/+boOnT
qh9bipSVDqNAd8VhLEEt0atsvGeOi6CUBUASsLmOJxK8A0Zg1Wkqa90hDkSUWWxJ
OVQ/tk/prAhlHYT4iVRth5BHAQoDxKnoP+HXBpP3nfFgC8x43eXlOg7yGpgzuppq
5pKWFwnDrGCzDRJ8E8FEStn3aOb3bnqEJO1qyeNOYkANl6PyuDgnDSYsFNI5olqC
8NIiJlb2d2YjvSMrdSnKYtvkSvFBT1mN8yW1oYhUQ8Ofj0qJ/een5AmaNicf/uaL
FBupQKm5Bkveb/FqPSMFGm5FDtKeagy2qlPaRnie6bz+ALB9exIHAjKqlOQDDj/V
n9kOCrhOEdKiMOTYta4/Knw7ZrVERFCwghnhWer2wKA70/7njo5VHz2Bz83FZXg3
OI1QNBNmxT2D5ngQn2ekx5XeV3F06ycVAnocXtynHsZktBvDHhLaXQ8ZzAgdMh9c
e3IQxeaVNZZQTfA6zyIfxJ4ibERV4kW+BVR8N+sXD8rUYhBaQ5I2FCme0VWUdofR
U2oEak2aPZM/4VXIEvnwZRjDjbhxLmKApAgbswYrqdgnd8RXujfzwjxANO2oPvuQ
g2EJoNsbJ49iNJFeLr9BAfTEl6NKTB2HT8wkKALn+Wcz5rg68NiQwsubZTGZwLl6
tEWZ0y8ymlzZJXVZQYqWSJR8HSIF5elusW0YjhcqvyvqXXJH6NGyXKzaHMD65f3B
55ZaKKU6gO24o1e9/MxVvttIe7K/o1jn7VVyZP+jFWRlA28dzQbygIiE9VV4hj4H
+C+fTzCdgW9B5i0DLFUt1jsrMGR49+3idM3uJ2oGAoTlJRMKPtqFv7H/H329lwWw
ViKS1MGAWxpXO7t4UjtIRrfbAJ28Udt74zIa4lApEgpq4zJOuA2cdifGijJDByeX
6VyXYvKA17/CAgghsaTTru5vL2DDUzE3bQXg/Dm6RlxXcryatpvMlZzwhmpVVVwr
XYwDmWmOj4U/S/SDVbC9tiJtBdyD2MHMEriyW1izbjBAs3yvAz7SFqFWtCmx0z2v
+EKdgBNJkVme7KRxkhfloQ37l481483YSHVHxTaJkWDan9k3YFovEPphBFMvHM1v
v0ZLSUadE/3FCUwrjG57my2url66p/STHzl7WyhxnRSikqyH8si2fdj9c9lecVjh
EgjirvCnAc6E+WLcY83G/2xm5b22rNWVBxJjRScuM61u5F6NK8qJAMd1s0CYbibb
WIA77YZwFsOCrLhFqKHSaYGLP3VQ+xJN1bVhYFyi6YYdUudyCabd3TMMsX9FtnGe
sL+HsvPyFCyTcttuAyGtg+p6loWZpPvpIMrJeSBINW06pEx9TxjCmf5nbxTuUN4e
Nav4PAYR6pGS1uw6VTb/qDSAsD+LYZWKfmYLHxAsfrc3SM6AwEmsrzqQi4+r4wKu
4Fd/kULMzEvLp8AX3aK4w9FtFa+zYw4DjsTqJ3I9AOonb3UzPDZUbJ+K3doDSaNc
zKZxXbU2fzdkHj7I/vwnWIRZIz2/s+5kQzEnmsZPLQqXl1nbQms1LR9X0M8Tu4gy
oiRPH3iAAHPX8SiE8Y87arCf30cxAdoad1wXF+J9duJML9SHxTh3Gvh3Hdck/9+2
Ny2buGpqFOxVW0eqYo2qqzjvrY6Fdp7wTs0HrnTsdEL7qdpuu3LGe91HxTzZB6uq
jwF+Iht+TUK5eQ+7RBg7CZSBxuwpltWANQz+ELeJOC7YQykiG13kRXZCMvZFhdcJ
/UceDu6+IzFrvSrwunbInW7Tjrc8gNLqjwzBZv9EDRUvIXPMFmMDGkvRgBFPKnN4
bRCP5qqUI1IH6m3XnfWQjPpmcye6tgR//bRgAKkDuaYwvbPHhajYelJ+U6MhaN3v
3XNi2qx8BM8tzsfBJ/GwhNcCKcusbpzbf46tMaNrNsZt1STxDqVedtChoaTzUrC0
XrDJmYgrs1OJSIUo3HN7nZWVCsZSRgTWgPNY4n3dHHlhg1DZUgdALwUJBgv+QyH1
1x4TXvengr1CLq77QuzqO4OBEkv6hih/PmcMMk4amCn8A4EfKrvQpBp6iOQb50m3
Oy/kSAfBWiGKzw5U/qQbuS+kqcHl1xZHyAYAV+kwVfXrLRSbrwXP1d5muhcPnwtA
duL6q3V9VWqJ8XXuJeap//pOI0UlH4sq1xehAz50FF+ZtOViElmUcWABQR24BIpD
v51+YuPmwbZxcJGDnM1AqnjYxNtSe3Cjro0/IYFJ4VdUys9C/62dKptKmXzyPjD+
Uk0nGAwcNnCgmIKTl8QH56uAymH1cK2dth5gKRJDk8UTx7xE1OUMLV3kLj8YoaMO
XKEvglLGNjaQTdLqcWncGTfHWs1yKhsQJmGiBWRrT8zQjI6bxCXUz4Nl1xGnEupE
pg5JQGzREyMdxbAl0ANnO1Mnv5+vgCIj7Oqb1DqAU5V4GcVUpsOKNC4UdB73Xsms
XjWDzmPnGVCecYHzqcdygQjsVjUUgCQQNOxquYdBpsfUNqM+NRgAN8TzCIqd6nK+
wQE86brenOnx26HDQ3mMJ617jaUhtcre3DLTy9rO4dPPA3fJUDm/YxBSKtNPaZ66
15oEOzP9DTsX7cz8WUmfPBKn8QcfL4VkxBARrYaRmCCr+NGs0g4Vxm0xyxs6HlzD
NHTxxt/W8vfR5sVbnqfb48T1WzjkHpeTzdiQfEKPWVXSBH/VP6P9pZNGFQihHfHK
dGMHHbXSe8XUlgnWUR5cR4e7q6HlP4+s/YC0oB+QG8pCj+9ec1nbYwSn5Wq45zet
bci3bygUj9wQrM1S5zZVy5EFu92ghhEKnLtaVmiqvsqmZSp+Ej4bePifH6BrSats
X/PwBJH3fzufk23MpmQgFy/iITnBbN6RmjwkfyV6PaCiIWV20dtKD6lNs5NpeHmM
KJk9BIp8GBsmlJhwXyMu+LReCOzsUT8chrXp8nVqYIPlIBQTUVtboikprsR1xiX9
lrJ21DkoQ3CyufIDj5DoJrRHIcAyidn/RZ/H8OxZdpo+XVgj9OVgOjsHNfWKy67Z
ur6+rmdcrIkm5xzr/FxY41CWeN1bxq62OEMlGe8hqa5McXdMTN+BV/3QPN1DHCBf
9K6FHJ5H2RSzNiIF82tEKsfjOlZqnOk+aVbqPCr99jLvqTQtuV5y+9o0alIfQXaz
sxutgzSp7UTh/2aywzAvDEWq5pyzN2z/ObUQR/6NHmD0heUfU2EvKtZzQfywL1Ro
8Xe/2Mk3uPdFfryuqDDl2b/JIH+eCNidPX+Xh4s1uwlxdT4M6hdILmbiGlpz+AXT
NLwXGDsNE2CdGebORYsrQr/KzrYF6K2hyL6Q7z/A2QzwngIwYqdrxCHaejl0LzYg
5UNejm1j4419LKry3KagNbJhL3bPm6aJeJw/GWOUSHmmLTQ76OJTUwWX7TrMkEQ9
p+FGqqHN+V/NRsXnrspFcvTkGrRAEh82Bb4SE6tOiukLYOqM68QBkszezPzCnrAU
p7hytQJG/I4BPaCi/0VdFnYraEhQL5PrEXcc1svNMDI6Uc4DGmJxYtVCSTWVbfBr
TuXk79AryQ+yywYSVJW+E9R52pSoKpZzwvLG0OcL68LLeOmTuBAE4SMnagBqvikY
YaS0nUIfQuuWpLuOA4VGFP/SFoQt/sN5qPY3SSGARs9dQStk9bAXdpU9bShL4xC1
yqVZ1vxwZZEWryzIMpX7XfpRG7BOcQDuuAe/welg9I7pYStqGQmjs4llWAObdXqa
Qzc81zBhVFvZ1fxg/VKyoO4pF2kYl8h23+SzPx1KMnULNyf8asfIkiM4mp5eYl6g
lScU0XZWR1yTp00Jfje0+h87P2g31ICEdIq56EPD8yu/AXAwE08/CFwkLe2nA9rz
CtleGOufpvA0Lscv6vsEmJAaxu8oXfG+nvL3B6jWYYe2MQl7syPi52yWO2HrAFrB
4/f4ghItPJKmQlVIuJUXJ5dGPT+Tnakm5gxr+sYczhrYhumy7lpu9yL0YvdhHDj4
BgMJhmOvtMe5G57kl6Bcjb0vtKJXdopYDayYQTZ9BI9JuYtbaEWmJfeQCsDRgJm3
KfJ1PthlzbZTIAQy7kY+YwYFWoAokdejzRteBCKOIgP3ffV8kXHT+9uIBAK1zhfq
EM0QhcrqtrwryOYLzo1j9HklgMe2MYuxXqzLwbIvIbtU0bZC8Ha01g0y2OuaNHGk
kqiG95h01tvDtKQZ5FrpVU3dERVEp9+VjCcCpOaBVikuXkVt++nBy+Ee+hG6hoEd
8t86d178XsWlmKZVnepf2tOA+VdeayjHJvkk84ZTOP/GIN11XUivX1qZ9yy5ZbNa
yZybyzS8YCIr8VHfoBQ1L/W4ylBSsIiK0HVG7zuFZjFXpjTldGjbdwlrUfpwk+gf
JZxURHUjDwWNUz5NtMczPCdVzDnBogqB1p87WlfZeg3x+pTHTzbmCZlidG8DMSMg
G8DdMNFYDJP7qGByM8vhnBVsyjN3pzk5oysM1tbbAHV8SlOZvGnhe58GW93+I/aU
pvRENAZHDFeFy2n7c6qO81NbqDsm9fOslyQD4Ijj6YZudbMVmrrxgn+ZQ1cPbyLb
WxJbc3RETHZhnPYbVkt0gZ5e+n2zHJoYIWeI39mU2lK+rfbTxdwwg6EwdZR4jewZ
D+2U8RxtheE1xEzSZKd3Gu7Xvh4MsuBgeVtET9bQWkwyEYD1bUIPQF6GRFNNhehs
ddedHaBVTPBPp0lFbZRn71phCObECkHBc8QjpzAdx7RuBabFXh+TQJyjoJpIzCXr
LU47mFgMX5K7eSCFAhOY39TIAoycIU44zNTBQ9JHWga2pcgHzShnkxAMmHFK4ZYf
q7ds5TAQ8ikJX9gibjhsKYvSFvGfIKvtEF/RhAEGQzgCek6DAZyrBbKV6B41dMa4
elQzmt5WshNJp8pfQzPK5GzFssBU86iiABy8LmTJXPUC6CRqKc9C3WHHRCHw+qud
CSu8TKta0d+sa/XoZC6SiiMvr3SHcgizRjbF76cTG8gG1VC4Gfwr9V+X21cqNJod
pDq7cLWGtudYvvYzx1+ysh1Wm5bPENE/zu4IzgLx0UZBqxW2/9RbNeglLNWocysl
+sWBTGuYKMFhj0ejNaut4iECiEirCgfgtRCn/nT5jmAdl4LV8BVNpI/E3/1HPrMo
nahjdDx5o281PRJ4rETY2BmrzVB+SNbzZ9jM+EcspPMoPKIlnMoveGZktR1VU176
z8Ofz2AIHW/T2oGI5MbuBvGIW8exRqdZPHe1oLzp3JAJXuDvzewwtspCmQyyxy7r
NjSnUIkoTegqadeZw6Ionn+Gg4X2dcJc/qsE0K2WrWZ2+hEX71+oGv3wGiNmqW1z
UxTDN3er5Jslcvys0g64HEa3f5VIsbRTfDH6dVCjbrthHD0BeCuO951+XpRaur0f
mQV5bCwe8/iBoLeNHDlR5ouaOO8wzfdQzmv/BZjHfzbc2c5pmIqlkAlf9MLVskPY
JWTWubdyWk4xhXiCEHEqCT1fRROclhVqrFqyLjawbIEhEbYmBRlc7V7EY18OAISp
c254Y6Yb2Ay251Sa4+fSUxcX0BpJehSLkAJVI+zbsERlPhzjBabE7OG6HtnmamzK
1GGJcdQ9Rt4qgKSeqMjlI/Yug+8I+VLU+lmO1phvfl1X+glj1tqPIxBBnUEdkVhu
zlr9Jpz2rm+/v2J59M/0VG2v7YakoqmgXfMrdPTci9ORs00aJDrsDkFrdkfxCGLO
WNAod4OtHQHx3yPOOtsEQ+Ni0GFLHaThchfo4z1dAIYbKx40+5YIR7SZJO/rWot1
wgJubo1p+7c4ONbjQeOqAfPEFGE1H0eZqBRbHL4CBK9j3scqYMIEnljwG1vdS0ED
IQoESYQSm+K/k9ogUO2uI0sb3kjkAyewlrpST9M7LFjZC8r1Chkcnj/YvjeH5onX
O4HwTbjc1REJZ73AlTsH6gVHXeJ+3Ux9KTnNKSLKLVC+1T9MrOrwrwBgKZrlWZGj
XLOxpLZUk5KKYiDywM9m1LkyXxWmbJePiZx65rdVWupfOAf2GRAQpHWBoVEKCP2y
DKbW8PvjcY0Mdiw3Yu+oiZrqBAvMphlj47SlP3LV2xLjlmao8bzgWbql8Gw/SA3N
MH1egYjCX0bKH+PO5Xvxqf58HTuOTjc4LRQyXxq+Hn8HJuCE/Na5HWAfVBdeEqcY
XCnB5WCFS1kisAL4BL/qes3KSXHmhZtRM9dT5kBLqwUdlWZN/y/3JWkk/H1fr8oG
CUtSYqhGeOlkaZ1mrRw7kqvDz4WhuOF88F6j8vMT3EL1Fv9UvlRWNn6F3RFI1qDA
VIatJSAu02F4TiAx64cAtJoPbuzvBWqvX8daPtIJgq5wMvkb+cASgX62ZdLjOu2G
SkYLCvNFtyaAkif0miFcWf4ZbjW/y0IcXEnj9bcSUI23BItHoob/ZrVrqlWtZPyC
YIXT51ScJkcyOnDZ6E3C4rz4iAdsWpEX3TLjVppPkpn8AMwPNBrbqIJwBDHyMv3W
w045PMDWlBgZD1Se35SgKJLGElVPBTj9EjC+MXPsDRwzioe/qUzRvqfqhI9ewlw2
nUeHzdVbZ60nGawIMjsbFrWRItsyaFTHuyhCoZCc+V5aWgrpd5bjhvMD0KaA4f5N
gmkjKpK2DxrPbxGzB6D4xMrWROgLtFy3aoqCD5D58Cknih1wDC/tQiH8bQgcUr8g
IyBg9VcS/Y+b4uYsRME5TZ+0xHdFeC0/Tcz4c83dTUP/lRpX0srwO/Nr9zGIT66T
Fv6FDxtXspXblzULOttJtKCeaWa7awzpwIvZngk/nPcDacoCnsuefCPO3wKfRGPt
fx3Cs4onLqvNZ6vwdQqN3HoMqKFe5GhGZCNxHFvp4rgZkh+YPwSjgimKDmRpSqMP
TDvAkr6/aFhIsH1pmC1509CxvFYH6snZz86GbmSio+GiB02JAZMH0bN6xN6rcwsC
XRMCKHGo4l2bCG/VFwMO4ljFHaK7e5N3P8VQkoDkPwFe6lJj/HXa/jkh2NbIbjKw
S6RaVJ6fHFhIk/Qon/r/0yk+9HefKP1Z0acLBRH//zu73qZ+xGHp0C0srywqKvC2
w0DrzaU/7yFrJtfBSJ84std75DH+Xl8QbqDrcXC5CUTQk3PiWO/p4peuUW1lNMZB
T7qS25CbGb6x0N1aquS+tl2180ZNtSu3iUGbvEldPf4NHkUDTwSIQ14Xr3Ye4ylj
YUjbFd+Ut/FeBoMB9YtVjHI2R61lvWGOZ8lGDfrR94SZ+bvk+8YLijnfMF58/qUG
Aax5PcQGulG8tClI3NLAScUT0SPrDMHwAnojxPTWGcN4aE0Z60VrZtz8dpmN/Otb
n0eJCWHbRqEnHxvXeyhhgEg80Gy8dmcDFaDSTjxP6u+lDqGgpqqD7xSBocl4912k
mfZ/oY1A+tBQ0nnax4U3baUfo5MAgRnwaCWgYoxdYLamVTH2JrmTFRcC347KM7ka
dCByY2cdMVjEj8n2vHRguRDmsq6OrKl7MMN+rOLAfWY+LOtWorWXeS3DhzgNElN4
iDatK1mNPp/D3+EDGPgc4acfY//mK570c94i1iE7tah1Vy3kVjFhlxY+hWYk1xZb
+vG2zihtdrp5LbfcYXBw+i/ySxOUlBhZO9UAPRZFavdaDlwxY3NVT2fuYcCkYd0f
wyG3wWURtzWCwQ1xDtDKvFuMGpbIhEsaR99WK5zEF2FONh3yAFwaeBakvGIvY3u2
0ydIEc7sE/k19OStIY2+kYRgZcVJqTK0N5LQX8okTYmgj69zVkwUeQPopgGa5R47
m3uAMS3mh/axoUwfQWaZL8UY/Zypbe4N+Lo5TmfVzzsXVg3ib/LRZ2Dl3behwyWP
0cQjn2b8WR05QFzAK3OXdxdlrPipveHMm9rmOOcJNnOEJx0zpZ1uAYJKeCFku2+a
P1bURU5hwut5TtpeAEei1bkmkZvnYZMJHdHfv4fMleadzNqeUrOH6VpE26Ym3vqQ
q7LeixRLYN4QHNeEYSYt36il7tkbuc9hAlvH1M7GXkI3gEaYxLxcfG5FO3aNm4Jw
zlcv0EIuvNV4UzLZ4TcgPeBsZjP4thA+QN+4bKpU5aUIpBFAbgh/r8wOJLQfYC/f
E/LI33CUpH7s9NRERfhT3RzrFLXHj1qbAL0znFdC/YnYtdfAE6bARHM+wU7YPpso
OUPbhr/4NdifNyeumwCIG6k46/HrWgLwLm1NJrHAvsif3WFS6YlECymgrr0DX4IQ
SLU1L8lfrLHmr1sTN/zNFNVEJK0Jj4zZGydP1WOy7AqUcDZ1BwZmnw+drDJ9Any7
fAAtR8LCdDZqzgWYSZ3A5hL/nkjveJ5YO9oX8qIQ7l6+c6wK+dI2GweAwmefT6b9
DbHzk4+mFQHClC7UNlZ/NQCULRPLO7FY+08sfl5mM6SdPbqhMtFgdaTcUauEl4aP
hFxVG5YQ3OoSBXns2s0A6bwZCM5viEEWQibVAmzkT3in/CXOfoKigp/cWlg52LWL
0TUti7eFq7pXmpFINWzloYUsjA0AAvNPurBUPxCbCYj/AwN7+7TqzxkuHbuwLMUt
gfQCGdKPe8F58Fgzr+yWw1XseYRiGRhowHuVRSU+Bh8E1BWNqFWAKKlxPqUn2IIp
wyxkHQ5kaUjSr3/1QlD48T8KmCtubbSNb15Xh6x+WzC9oXarARD/0rbri70fM/8e
o6V8uCtjupNy93pZCXF95P5/KuHxStUFGM/Fvt7cujAZbM4lJQMJ2x7wW6uAXMOk
The9MDqUdxE5M+R8dBRK26fecjQPSsjWUQVIYvujnf08VY5NXzoyO853nibQKib9
22YMh/EKPvGKAhcMMv2BUu2cS5Jedv/s74FyPL7mPVuTWmfBHUX9IWoQcaeHsQav
MqgfZwKnlltWzNpiz/kmckCEIqxOzn5nxQYAeGe3eZpOJMBF4tI7Zj0CCUSxBNuu
4emqEl5rxGHQQiq6fEpKQ92GiXehJe8BTtv9kyzWHlQA/sU63Q6JUD3dnE7/oPHJ
YKwaVUlRhES4WjBCbjuTSAXmbc5g2SyzKuHiuVE2Dvhzck7c4xTuNUxW2Z+sZQmJ
XzbScPFUGrfZ8K52blIYnKmNMMAU06ez31zOrMzjgkobr9qnOPeaty3kVESz2PUa
dl993BD6Xj9wMyMBk8kSvygqyvowFwDPsim3wtN3MNDeN5Z1s8tpbuMpbBnf9wEm
kx+AEqaHdRjmvTYGWdLj2XhQmJeSwRAfJhDc9xMHKY+2Cy0xYPBPjSfs95altaG/
vNunPIor01ePB0isET8+FxtIarF4iAbJ9TvE33e47DBe8IOocwQVqIoV0W3Jm6J8
2bTJV6lPR72Sdve+aK1FumfjB8BSMZeQ4iHoxSrr/HgjawhWuLGfEq7l0OxZYYfn
5Q3CUDcRN2Oug8P2ai04Qt5iL9MZtSr3oa5lIzAD7jNWT8ew8VtfIsX26j8c+Zxh
++jARGE40wNbnC6wnh2FFb0rMGAOyDCBuBU83B4Jp8hW4Z8kC1CDCepUOHKaCh5p
7NKfGi9ylm59WalrnJtL/kV0eTx5ltHbN4WRw/MhvoaewiSWmtoe57cez/29WK3N
STfuNv2usA7psxAuxlt1bg7ulaKPNEVyxj2N19aSJQZdQU7snAXChfvqM4Gng/25
IbgY/f1QHuBRumrHYcrbczjPNqMKXvUZhZbFvFhTmHsA6irjmlthzY/1WyvhLMtt
fwcD3yOvJAipJm9blgdjx6HS8SyWJr1B7trCAQUfOaMSTZLeAhzF8hBbsXYp6w72
+fyiiuIh/Y9GgmjwNiMM6+I+/xA7KD6mrgFb/dZmtnBoXtZEcUlA3SH9UmA9viL5
VIKOA+pKSJKWD4NQvhOMyqWnSR1aRKkMNQNYtXrzGyR3zawq5K78McyqzkTSaRQN
6mAL8BdWF1YbuVdDToN9IiFT2B6cn0TipAwl/wuEuXSGZKh5E5RIz2C9LiJST6Dy
LWg+oy0IyJ3iEpTRIwyMfDM8tcymkVcbe7C/2iwhJTQipaMmqxxjEbGFF+J1y2Wg
ENf4chKzXpM8Ib2XtXiAkp8JfI5dG8QYndE7kQUN2mXRefyt7KwSnHVd8L3Eynd8
zc1+mi9wzKq+oXRCm7l3pgbiZp1YIu04YNjpwExk3OL6ryIk5rvkjUXMrIUMaeCT
0CMz7ZXPuerlpSZyMw4VFh0AuFUiC2CHocMx4t+mLcQzkFN0T/6CykOOYpKPVJOe
9W6pmwxqCp9rDcdTPpCueYKY8q4ucmghriIafuNKbXNdP12UseFP8P2+l/9YgWar
Rjr/QvdD7PFOQF8pYSSM7jHGXGE8k226gRSLw5IoEztwajxSYC4OsF7zRf2Nld//
7vTbR8/6ogfnXL9oMHTDKk/kJsLLfDzOOAq7XJHBv2rNgeULsu37YRGj7tlUoKwc
RbPuEp8syjDi7pVixCXriaJN5xKpMwg7RdakrrWP4ECccO2JbqnBiFMFHxhoYlur
5BoDdBwC+GyhYea/P2/b5apmc5BulYJNdlr5LvBBJdqkTVnMsE8FfhVdP/TlKjIj
7ejHqJNYbOfBeZ9q+09UjnQUFLa49r9Xq7NVuMyndII8VmptwEJ6MRguSecxGOnC
JUuMDnxaWEjNAe0bEYroKYy+LBl9ASa6TtwZudN7Q0NG3SL7kL6N+Feszd2Vjl30
Dp3ggoRCfrONVjM8ghfgXpO+J/hvgzFzY1RYEdzZODpH7MQ5pmV28PaFcIuGBGOR
ZPxy9xMXc0fgx8MKDDiP2QBhYjHTd+Ko+BLFiftYkKGgdMwuu+n6a2jZhjdT0au5
vqF7oYoQM9vlpS8jIYU2OD9rqVfBqyW/LGwDQKQaPlx1Kk4uBxHQSyHfXLplU4c0
3HriAHNU6zWXz9A00yKE7zQf063XxYOL8bM93FKJrRd/Onaq7D3xRbkO2KcIEqkv
K13ro+ipkYNCftPkV3fdURyrazw/hS1+XqurCh85MKupL5oesSbyBozoFhPI5qKN
6P8UPZcwv23n2PZy7XG2S0cJqP0cx91498SAI4N+6GZSF8dRJNyc0ixnSP+laVr4
dtRsxBiiNT6kzwgQEqN2XAik4oeU8Qt83rfSnmOBB/AS65sjH5tLuEM+wN0FZBf9
FDkxe+rlH+AWAszU1Su+Q/yJ1Hh6f8t+0k3QDmntlqJkEc4Fa1QZxYx02Rj0jYZQ
Vg8sM/4nUVHUtqjmxicfMtrBf/fzTNcaT7ERJJBIahqyyTkoKbdKJujX6YEK/mr2
YyEnZtt3qSEBZfh/T+BpCmfYrbpwgbRO6pYBWag88b5+RdGSQ5I+rYCT9kXEvZB+
/g5YrcarePeO/5HZq+TqVb0LFSr/LfO9s1VdG1VfAysshbQjjcp4BMXAqUJjfuUF
s/d8/92fSgk4Wd4FpMSsKAG1MTY6r+yPPwNrvHpl6l5LxBePktVsZfo6b4og3cdx
2vbvXcvtKNgHEhfoJ5dWCWdiuwJmbs13hqIDS6iCRQaZpKo5EWCwFLrGw2d5YgIr
acl3qW38k59domGukLp9+aJVdS3WkaC7Zfw8TdsAkwdNem6C+ys4fb6pjmtxXd/W
q4lLE2acVsDzDc+PWwUFrPjcCuaiDJTX7DJLIs/FPxu4C3YNzS90Ng64vKnVehVM
hYwzVZHBO2ySJdblh83ry0j0HWrF/E6rxcty8X5rWL/Q57q6ERIjcV+TzQXdtOmd
OXbh+ZMp2Too10bWxrwc0nisr74K1EVwJ6zAgnbw3L1H5I9jYs/SJ8jJNVP4JbqE
HXhpRhPxzCFHx4PLtpJjQmZKbmHNr2MBWdkCbrEQkdEdu1nrq1RT7IYRHB/gtaMT
a5SJboqXSn7U3GKk75GK2g==
`protect END_PROTECTED
