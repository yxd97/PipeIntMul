`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+x2qzuJO33vVcvMu4gxmATGMZtEovjTvLc/0yTevraVG7OaESuHBaeQTbhy1XFVL
3AdR3OXw8L3u/cakashznehiJr4ASqyoGByoDuzmngOlfvHD0k85AF5/R0npFNdE
cJ+bT3JimT2qp2SyoTlvz1WOxxBLK61fY/UhIrfOTfWzFzMwFCRN5X8/sWbdigmK
rV9w7gtu0Ten7hsAyW0jdD0PW6TpnUcZgbClcSybH6bfNU1tU4L6JA4k7+dDo9o5
tHQyzXKZbTW0LGR84pvFT0mS2p5l+HMX3MzJlwgZDcTCFC8n2xQNgbQ7hyltzy4v
DcFnkJeIiJL2kSlY5ttpmYZt6LnNNNDT8Ah0/zUvs3V3ZfqxTcdXgxqypuiUzDIO
Ti3SQx+Jfu86Oke+yb9Xxg==
`protect END_PROTECTED
