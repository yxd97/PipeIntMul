`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HUcx+pP+Bf2FyvH7KM+6ERe+S479i9bB/NH5IcgN+1PkoDDkgGshwURMkln2vTT
sIHP5gerMp7hG/eZQ8P80hSi316pbtyJGXs86qKbubtnZLzJr3NuIFALWbd3rHE8
LJEGi5Q0pKKGfu2gb+/C0A3QiHsIT+7FJehIl+KkCccAaJnnrSBYgqenHeW9Yedg
KVq17zH2zrwsb5GU3ExPXVEzWLOQnJ2Mk6rIqR5Vw8XR4fBKV8X6zfBVtSq8LkKr
UfuSyO+9VzSNBkIbhK2xqo9ohJT9eolsRYYLz7dUZHdnGloO3lAnt5o+cSMiqhpI
OaphHTDUoWIwfKJRPVxYOFEODIS3KfQRbmLN5U9dWDk=
`protect END_PROTECTED
