`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZkkF0WX9E06M/4ooiYFXtZ2MXkR5nJI7/NtaxegPBmuZT44EsBhthlVgxyI8AHJu
X1X1TDb7LXCfYgW5kFFhwJCQytlDKt4WzeQ7NuYPhWv8Rqbme3F3tkzwmmaWv2c+
qNy1SOr7DyGlkXChjcQedqAz3UocnVnUBwIL1SZ+4UMm9vPmEHmCap+M5mvO57GQ
8EajXNHHOw31sLE1IGwuT2medPENRgSmPkf01k6v+FUpzbvnhu1kpPmw0/l+y29s
EQeBh7BC2KsAAnqEtZ3daXaUgQ7PXIAiyNTnaixkgi6duKWkiKK++YoWfLSDredG
8Tf6ZwwohbQvdu2puT00odTh1VRamr0wDz6LoI6ttRsYmsBguZsaEGpMMN12rceT
/4k63YcIUfJUsmp7Tb49mG3oOhrReMbRKlOr0psT+x1+hSmbmifp5UBUIivm5fRg
o7lzFigs7th0zoIH5ZnvWHZMQJdzn4FuL1jRybfpPBApUX/H3eibPDXY0Cbm4u9+
zc72N8geHDF1T7a4dkORAw==
`protect END_PROTECTED
