`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXN1PeNgjHcZtZ9tmvEeoE2OMOy80fVPMNTngHTPJ6/9olvuFBh5rGq4S2Aj03HZ
LBMlPBU8JA91W5QDPjY2oe8Jx2aXk5OeQe61A/Mmbkl6v9gJkbMALfb9f+7bhmUb
VbrRSwRicqOYbmhB1sykd2V/b2ldm3m6CHyIMIOf3enMiRg9VFTM28CbWfPZnHE9
15E3DNDprB1aXBcPumQrM7+Zmnyyyb0i9x0QFt7s1rPXl6h+BZo0M9BaEt9m/uyQ
uZItOfqRQjW+Q9mswe/N/TReuVIgpJlcTCAmPwGqcVNVV/XK5BM7aupIkpZRURqV
1eX/lfUYcKP7PIGczEXiIzgsPFaAJR52qyEi6cfwjoTDRgfjQ+k83jmUiBh1r8cX
WlrLzTGZIJkcs/hRn1U2fCa1nEcEXUwyZJe6WOrKWYTz5kzfRsvmukpcBxZIu9Ik
sPOzBZIs1gzCzJaagsqMOwbK2ZDBn3JUk/HNPvXKNppjbKOtOl0UIJt6JpJPZjFv
lWbah2qcBwulXe+clHUGKxnZsY6g+QzWG8hGVr5wpd7z34iMKCkv20Sdkp2RKdhz
1nMymwINrm+FU8ixUUL/XE/aWmb81+QwLgVd9/oTQmmaBle/TsrQeODHTEtEa2CJ
//JekQW9z4PYrAq8Qiud5kK5QcGbdIllCdtpfI8s9c6iyTXYRtJsbeH3cu9Gq6lV
UDoziRWEhm/VqmOZmxwaraAmxEc9WrEuadj0dMXwj29rjgAUNTS12v+5taRYatiE
8UYmaxOmPKag+Qf93ZPxk3Xx0saj74oexQb7v2FKd/MxAJARc5IrqNIM79Ld4qFt
+LRuz6tkNllxJAyj0yq7qByWSuLTTllZKcdeh3gyLNOErrGOuSB5zpiOTVdpWNGV
3HV1TC6h3rfVJgue6ADBAEmja5Ni0ObtCVFVCOi0Roq5QdD+3FjfUmFcH9Wg7LCg
vXRm5oY49T8kLOTsQBQngv/wK/TKbmTJOMUP1uXBLV6DY6y2rhKDBXobNfrNOGp6
pGvcMoPm0yZcrFBpgcCkFSiYXfKRd7YdQhj9f53rrkYfAfJJ5+mzR0SM47eWD5RD
CQG4rNfATs35lWQrI6YCmF84OLaXl/PXlxx3HxxBXz639zi0yFdAIKXka9ykAdjq
NEwbeSdjoZJunP77zVnJjTBnNi0oDzLunmK6utZKHkc5VMqNV/iimWyYADrqJSv3
WEURduqFAppGK0XNRjEc1HxDKLKlQrpIssDq/rs+p36cFcqquJARGWvv9ojrVCTN
Yx16iOtBnPd5WOXo12pkeeAy0jXY3dtfTwprkMyjO2rI74hI5yCNFusmNIYxfBJU
bfmTtMgc4WW9YdqqMSPnbV1ekrN6KOoIUh2f9REO/GSCz3W8c96+9aRZvIXcH0yC
jdiDzrUbqOZZM9IUUB8rbkU629wOzYFusMKiVCEx3r7VoV8ShqbFy3XLrddyy4/g
pEO0x2k6TykF3kZjCuZdVrD4OqUyU4+WMWoNKaG0ucDItJhUcOsT2kmQJ8ilS1XD
QHnBVQXF4aYXqkqEShEl2TxafL7Nl9qDwyBHTL+3dqafrSJOaGRcpERUdObKaaeG
JDzOhivUNR3K5QzPj543xIqnfoWVZWTS0LYU5P0kRoATT6dqtWFjgrWcvjEh9OGt
UE+57meNajhx/0IxDO016kTY3SJa7pL4Lhh+XNZItOS/Ve1gxEOH9icCIjCo2A+i
BXoe0DFjKgIjCY5qW3pKgXm9HzFNe+lOjNTLZMlAFhN+8wI2LpTV0K4Cb43O84ir
OLrHVBX+1foJSoVGIPPK/nMS1ECIRNJHh6/fXnBV6z2qMEwodkFlU5p4gjMiOnGs
yqKrMxYzqYlvT8iqi0kpqZuEF7/c/VXsGi8R2LXjSwQAr+fcgdwL53ZBYuSOrDEU
cl6fmCuCYNjpY4+/Rbj2D/Wj+PWE4r9V9x3iZg5VNqd0HyAgq9hNjEEIQWPc0ZvQ
6MEmhXoAh+AQSZU7Je7T7oGNpFjjjP3TZLztdJYFk26fjOfQE4j57R3VaIVMuKtY
v4vBdt0TAG2bey0Uf9ecwXfOPf95UrfbcOW/tUDEm2mkzziBMlu3CPAoxoT5Eoke
puTkmm5Z3KlmNqAwwuoEuqNw8ir6Y604+ar4ODZHO8dzwSxXAdT07/OIl3rs2L9v
4QetSJSZXUTdnWq2LiSdSYiXuwhRWW1CoiLtdImQfmeb0vNsgwGDJ741GN8AjMrY
dR2VyY3JnNfdCrK+WbRPvqYUqsX7ZB2xFQgTTMdeHbaXf3Xill76YB4pj1GP8g19
uCh9ER78Xajp4Vt2JxUAl2H27K3dROGMSRjBjdbBMDluAoJas6mEIs43pMMi5q75
Xs0TyBv1nHAhp/X5P4BUGT99mFJPUuxkpyNVCxpSC32+kWoqW+dZHPAuNjjyFGYy
VgWqnrei1qFaJRgXl3tzorTqVq9DDVhDAH6Iz7LLIerFtQBGu1aaO957sHfswXD7
n3aXcqa8aYuigewfabecZ/BmQLnzwjfAwFU1iReC5JJ3MgAPPxUjUCBZnqy6Fjjv
ACgHaPUd1UWrgf1GBtvQ8CSsfFngy5jTHZhpY+Lje4HKuRKHWvWOug6bwoPizWeT
3ckSmnIfiAB8PKpxNU5kyln5mo6fWkj9IiRunbusx3K7qIXb6o2d6ZAQI8sxtSnW
SnSe/+5hgocwvSc3a8Os8aicNUVdVx3nmnM+xHm0PVFzKCWWKPGx/0gV5+hWczsq
/3//E1Jb4mrWpHk2B1yJzn/Swqd5pm3THCl08C3s0XXBI6UXmAS8+ZtRmiEtr/it
YyxEIOczqUCkY7j+0i2iA9bglFruasbKHTLaZyHj8K6m7xp/AJFijw7283nUpy0x
OjJYF6vP+p/D2n/1okAictwTRFc3c8N1r+4iNZXiYLZ3j7/8J35r3QzgzIg3OwWL
/RfrSQXT6+ZpRixinb7tlmDOtpdjP2DEHHoU+CGNi1TxAXZH/aSZ8k3yGkC2fJPS
IwzrT22OPI85YAwG0z9fp2J5P+a808Yp7LYK8Mbc+9K5ESyHIwZeqQtclRjqf7Ec
16EsA20Z1BmI/5WM65iO5d+w2NhftVRJx3o8J0HU7XM2K9piiWZTfSCLJ6CgCKJM
zP8Y3meokpC/rSKtHJfvQMpZ4i1hsvntp8E/LQYP50Cux8k3tEoApUx8oyb53dhj
phJZEZ+31rU5XvknKFIyadkjZCPb4VuFRz6KvBUf45DIalzAwrJNORnEKkVWLYzi
/ID30E53w54d7TKHzxOT6nP7yR/sXGY80Bkmy4JIULrp3dTPlXOIO92/9hRtBr2j
Juaaaj08pOKsm6ZovEv3ZxAPKBcPCua6h2KrPruE1res/MUNxYPmEQP4H92FBiVa
FHmOOfRzTi2EEsUS1GB1p6IhKsHk/T7C80Y8RulXyrq1JL9Pd5jjxMPkVUkqZXWS
msjqs/Yq6GQsVvRiFgs+jUOxRK/zcje6AbTQvf1MhUMoGDIV0jtJ7xzc/+gLrJqg
wTlbkd8UPfkHxRciFoc9lqgN/moTubpEnYUT/JwfBqef+fWYbp0XKd1ypA4tPZbA
dFQgjOOZnv3ekXIjSO0qW7Fm1U7ehkCVCz8ft/sFbl+BHYiwCqa4MyN6u/pjGvdq
jICDkwD2disuTa4uLQEZOXNetKSnxc3kZjhdSxCjlL+RhKrWCUEzrYZfHF/N2jM6
XfqtEOtDmeAg7OLex0VC5wGX8gPDtrH8CA0JymKnBD7DFO58+ZP2V1cGdvPn9AIJ
phCgulTFqT8sbl33ho8p582Iy7KNDXzZkBhuBcWRZ/QY513hXe+XiNhy8rC98EdA
w8TIEK8rPOEbTKJtQ/LCGa/Ppeh2kFaLKAmyBFyTEsKF7Cjba0T9MitVozx6k9gy
hYTAMXUfFW7SErxaMDmGcuCIQN6YOd6qUQgsW7NLNin6DixsPLMdz3i4xhqouZUi
21SC08RSyB5cXswFd+hWHIBef6di+ZIyqwN+pEIYrnLUjhe3x4j5XVdF+DJ5EP93
ujMoHVGxDatrOeJDizRge9s8W7Ff8RX5k1od/RbeZ8LNUleYGk8WLdxj9tmZFXkl
XRmk9lF/oj0kxyfWhcw7C1/A0MW0UmptaKL8JhtQjaQQLcfnfFPKiGbljfLdQh5b
E7HihFMkNfKDbjAawB+JQYzYTpeSZSGV0B5SaLEdDqEH9EQ4wscGdQeVQ1Er0VTr
znZ1Faf70e208HnBHH5ukejP1noYogd1ovcwn7X+k1yZ+EiQNbwWVoZzaCVtVF/n
wJcA/ZoO5MdojFSgRE05KVznY7JSNxGiEZdpPTcTcHaFnWxKYs05KAvyRaMGe5P+
0YqnPzeWjTDa+/AFz3w4HSbd+fYJ296iq3G/Omai6qUdpfrhyPLsm8D7UntIEb4u
rIhSV/lb4VYIMLXNFSZcTDqia5Czh5/4Fg5FawbHRPnEwjfPm83MUx8wDz9jJTia
gbl3ET4m8e2mfszEaEEzi5gQW6ux2IwGhLlVKMfA7fQQMugDHgQ8ZENNiicJw6hD
a1gDEtVSo3/CI+FNdXlDOf/LSJrvSHoxMwJIyv8Aermq9ZJWDkkcp6K1nNIiqvRj
Mhros4HHs1fsD2R7/Bx8NS+PWm4+a3xHnbjz8wwc5sXV66NprzBDK/v/czhs1R2u
VvlZaNuCYIDtzHnk8aOOg/nZlhh3j3rbx+83hrLoH5lgD/I1+NIzOnccdn46LlAp
KfrRKfRF58pQNBGSA9gwAKRepTCS5PpuGSe5fedNZC1lNUFsc6rcv3ADd1m4kdNv
a/mzU6DfZn9T5ZD+FktCW9T0uBdIGtKYRtjqm3S27vka28budn3Adh+27yZwSMLl
bxgif+LBWtZI3TArAakEMA+wi33WTsFmvFbA8jqAIFzzHfV9yY1BRdbiFCj6G0Yd
MUm8UXNneKhrP6k6ihqbITwaXc5usXr3zzMzbOpZtBDQXL/sWb7/uvMGIFLIsta+
Ih6KrdWOp3FsSoALcoufN4J/8cXWpZCLPQ++KbJg4hfeBiycYgTDNGyQZX9z16Ua
m+2c49tOxIscHYUadScajstZwThk3BALqak6XvMttJEQemexWkKTrM5jJmhCH67e
bxDA77eFxVFXrnwtU85UQgS+guIEufCxFNyI38dNgjljQfNiT07VfTp/vaPuU9WV
H7njvG+14+RzYWSJy/wbfk+3SyZ9TnqmUCYvJkw4WRGQ77/j09JDezrHhiuibYXy
zQhCSP/8UW45tijj2LwsmHicGk82V+fHK6go+UsgZfmJLyNv4vjxdC6UghKFcQb2
E4Cv0tNNcwG8nsd73DQoBGrpJdAfmsF0GeJ4R9fJUytztYeIjUYU/1ldCdo9fzzS
BnW59j3K04wtUy8/x+dUROifg5Bmnz6LlN97jrRakAwr1iFQkj9vVnwxt+Pd7anL
QOsxg+hfHwciIM3EFz8r+59PpFjCnYIousArK7+nfN00LrUkRYCDxpHM9uflTedl
g7JfGqTcGpnuV6eC3CHrcJPVTFQ8XjpnbwtaA7m2BuNzobGVswnYZsq2xhSsb5Zx
Rh+hm4h7rIxNGarL+CKwAFmErUPxqxntF4I2OzWYJXQsIeoUUXWGRmQiTQH95gwS
uZVYNY3YP3NIwEwTHmSV7NIc86SS5UvEyuU6KWCIINweVJim1Jeh0hqAOse3l2yb
s10f4O1StQgdN3LwxlygRooZFGqC9ZwvJQA0IHAGBTIj9CbnJeEcaZ8XUXJrSKTz
YyGTMdhWxkX5/tSpkt/+nBCfKEdzgSYPGDWYCCFhYD0hJNenGVmAvodULW1Afn+C
44FlidthxB8n77dqU6I5pL6az9QjwtRpueNsja7KgVOIjYtDcxzzAIYNHlxuVrqI
cx3mlaq97MgF+7rWqMHDm5I4v5lThM0deoY14CcqgPcgR1H1l44dhjdknN9M+PF/
ByAxofQ85hfHIAI0noRc/jwsOu00FjdrASyi1bFyoRzN7XbR6XCuHE+raJFB3QTH
kEPAF492beiGYaWkWLuxRQtJmI2lRg+c0lWS3l2YrkTurT9oWhMFi/kTF0EG3fvf
Ubj9sGjOdCzHUPDxg2dvEw2WvKXyhBra+VN90ekWyeOQTF93dVAS0aOEvp4ckVmU
OoYuRZ2wqr2goTUl+Eis3DcEhy698GBniLxiaUzumPtiwFH/4f5vHc4tbdjaaKjm
X+tDqVGIfSzyJhPMoONPSi5ch3pdwfk62JX7jeSEcCmfmapNSRUQhS6fgSBhHQem
+G0+oSDMN8E3axJojQG28On2dEcDL3xPBiSN1VU6ZhYGzxYw9eXyrlRNL2qOyoWc
HAA2ZM1zeISETtwobg5fnPi3kR2MqaFqXIkhJuFQ1i+jxz2e3JKUb4SyzgzahT5b
9oT7VLtccrLfNVvAT01c7GBlrw/yLWP1IkQ4gdfuCGChSk9kQ5YpQT5kwdMWHMy2
05B2G42fyEI9TsL8IfaEVNfxWmpYRQGai2qQwKNJwyni/foIt8XC4Z5tXRcCTK1Z
RNvcthrmbwNvIWCFVLlu9y6Ap5/zmf34J29efY8+9Hl7XB0wK/OZ1JMfxgGNdyCL
taCeMqMZ5u48qN54YcjWfQhn0jFlWL7H2tTj7Dwv6XsABS1fpdJ+gAIpDInWBT1p
Dry+s7JGQuprlysC9cUHnEtlaQQHLO+H6noztzaDeQLj77io9JDJ8MCgis1Qd6Es
TRAzhyPlM3+Hozn7t58MrF+dvFxEKPqiMEWQGsLiDoZRhbwDfmXl9XCMQiUnOVQI
nrePYYuA/aDI7RBfrwX9oKIyXYD3aa5823s2aHWzoWqvNH0HpsyQIX6g0EvfMuon
rzRpVRqj63CQ7p3132g+0G64pqmYasQEwyTHkhFtqyqrR6yWudf61VNpCDUURhuS
DJqOfTcD37tulGljbUR928sWknf0Slfd4n0fgdhIeRUr/8zUJSrc4vimOphu6KHB
Jt3fHM259gdTb3KNp3fXHAMGtigJMqtEJIRgarpTwD06qO0QTnQOF/1y6k33N8Kr
Fcr/o5MXP5zrXGddOjkMv+mkGdNsYdVghthE+opOp/zgyKtv7R9oBMTjvR8vA+Fe
VhTxq0Vc2evUNMarT9qD2zamazjcm3pbit/l1LmMDhT+oZClopzUeY6NY86ZbcI7
VmaqoJ86Zn6pp5OJxMDjFRmdGJLquSPvuIGiehPCFEZAipftu4dfHEaBQ/E97MJe
qmu5/i2yPsYUF/p9txeHycNyNKcrps1opmsgzJu4sWYFVGzGsmUSggWOHMdee8Ra
ptLCu5qidRN+r9H9k8X6/wBSwVebNxgD9FqKLYs7FkCOQHODlb22MIlvdmpK9pb3
+J+diEhTTSn5/VGr0HnUrF/ePOIjEPl5S7GNrvXPXQv/tn8oTjLlj4W9SC8JZlM+
BLPBwrdssku/wL2kzQhWm9h1TIvATu1sdBnHlTknNAe0UnmzXd8DjHZLizQfUF3k
8elNGl2vxFZ/HOopn58w8lmIwk4JmB1h9jSCCMRdE3k6dT4aYATVIgDv6gBhT7gj
ywGWhVFOQ0RjQCfpaJxjc7vBXgL7yJHw/bIQEsHePS47a919xG1AIzeSrfsfuNB+
6dhn/waxxNOWoGJRaQHw9WUKGeSywD4AsGL+8VlZNG44W/hNV2dQH1MfRWDdGj1E
XQ3532kSchlqiVtvD/L4IU6HwapfqbjJhWqAny/exzPTu57aPYjaebtUQ8bvx86T
pVYSICxlFjQ3fzvwJL0uWsFyW2ImD2DDGrx7xgMuUa0JvN1CQahzfu7jgqQ8PH6M
HtRehFr0FTZhhB7vexr4dzCexjGw9cx/DEn/4nrVBdr9YjCcbTSqs4nGLzgm9Sj9
kuKehK2bnOzAr6nUy0GoXByGjB3zoAHBgELt/ueK2IM4brHlgcwpB9eDVoTcpn4z
2p9yZK5j4eAH2pItF0i7elCwqIRb6kfEAN5CxJCbtrNYZZF781kcex9OsuYnYNOs
14F+7tXUBi6ow4T5dZWpO8ibzG388D4XWcMF7Tf5PEmsm7V2HELp4GSYmadgli5x
KbuaqBiatGMFeREvnu8BcLmSuw4DYQYTf6TMApgsjbyqERln+RP89oukZb4wQboa
Rf1n24XRfgY8X0/z+Kyz5gqcaJPsDTxJaIz3WiFRVK9z4Flr6SF5V4BmqeOml+au
xr4OAUqXMounEQhZb/eYx6sQe1/y39TfOZdmNtz3AZnyMmo4XUnTLk8TykGG0u/E
JwlhyCfmvlhZXpk1zig2p014qv6fNnl4nmSVIaNmmOGYomVoQmj9kBXL8Hzk5FHb
Xx4VyJQadWSeZjpN2ek6LgY4OQ+33rLEL53Iy3gE+isASXoziJiiLB4+knhQi99+
GCoNI13uC7rmYS95lxoTczixjoRZWgLePfCL2cNyKhboFssjzeh32Gj8Xr8l+qjf
4i9QqkfqFxOSdXpunpgV5rzYhG6sGm8Hbe5zvQJwrsyUnW3q75d1aacaT0YdyNie
IUNG09TdRckWVz5g07LCBx2eMXktlr46tjOgs8/4QZzMnHZoOM5W0HX5hLc6trDB
DSys51/IMJneIudNw64m4p89egdCIZ6MS+1TWtBkmcd00yGSlNO41OSDyR9SF6Sm
SOGlAilMhgzfX42wuHF9fwSOYaQv7vBHy08f8WYUrA78pWW/J5AXElsnZoWkL1TV
ig2WkLQY56b5Zxw15Ym4GELrpa79B+K41TWPk2fnkNL9krks0v5i2S/4Fv7EWOX9
Ecmx+2uh+gAfIJZ9Xr1wc6+M8SUvKkijZxMp25sUAF4O2CuZ6VZZgoGBtGPFwEJw
cMUP876BgH6cdDAzRj8ukMn6rdsfQSvhM7syqZGRlyTMEmYLr5Id0oH+a1yTfV55
CO3dolT9/xmUpVmO2N+0qwtSWZ8DrbbN1xhIzsFcuEXZ4DPLzsNjF+jePU/Uu6Je
YtCFQJ5nYF5QHQ5lWGQz0sC/uUg15jb3+8lVkAgQmz5EHgg93IMAC1gNOuIR6H06
zb3m7ws+Zd26T3UVrXM7LRsHTqxYaeQiIkqN6+SX6ltqiw2y/u66QlRv+SmYvGTd
K+xyQ/wsQK2PeMUqwThKHz7AeyaEv8aYxZTPtBdY5Q7L0X9JtMZooI7sDV9+Nw7q
6VAlDxVcxlqWEBhQ+eVVCvWwV72OeWjugyo8poKX1zuWlCi4EY7UAlVrwTCtSiqw
uqGKbpz8k8rtSrYUsz1vVfwwuPxAVCdF8VzOL1Q9y5gZW2uC11VMt88KuCzJee1a
4TIvop5uTACGy2t7o8WAtK5iW1FaV5ZL2dQoFQNjQoEuSSYBRmJpK8FmizM/53il
ptw/2NPZ1FCvhFtxKfHND1kjrw7NVslJUcYq7pE82EabPubFd3VQm8qY0rY4AJkG
+4C1GzDjlpI8CH6uX/qAKpq0n4+J43efmYwAEuiPTTMspN+0PQpHmHU6Fzr7axAi
xi663m0Ot922Xpn/wlJXri3tzxTlrWWvFXyo++PRjRnzuu3QAmi3QfxqovaW1TPo
guUqftZn72GlhPoCCx8AXuSw53PUDONGw/ArlTwaScsIppnSmfOVgj5GQjhxi2wk
HFvtprFTS5cnsDeQ7V5w0bB/0vUNsOV41SbtkyiYqiGxp8zEISgeyd6JmU0KkLMm
1f1uKNFTspFhrxWrO2JZJHzFzD698n0raKg6hS3975XTVmUYXs+3DwBfIXTgVJA+
PnTnUEg4SuX+j1thjMWSLo/GruIigF3TouLmgovVG7kc2o7CKJP6a1ccVlvWhKAB
Ux3Bk4160jFKfjIqDK760VrR3oA4q/G2nTf7I4HdoWEYT7qvTB6bufBPvQCj2MuT
DkEwh1Bol4AQWhzyF1CoEa35KHYtltONaNJQMjHy93njc7wfnexAPxxkakhbqaI2
nU67GyKvmd7kqmbb0wRqgJHY6qLHZKdmOofAdoWETLS5SfCFr7ereNNJh3t89U7R
Wqi7nGDnMdoHzBCaefQ8zBezKz0uMBe5f9WDUVJh3B+XTsGNyVplFHsDHL9iK5yv
kutWqke4NdTu/DXhQV/5utr6L3IFQE4zJ5ZdSqLhgpSovw+bC/FCXm3p9rxcMRDd
bO8rNyDEiZmPmm7LXsoM7bP/DBNHstPfML1iwAMwD7O8obYtySQpiCVRmdDhzaX3
AnYEAFyN6rDZt44v7pH+PZjomgMfKkJW4HfnEaEp0IDx/gOcRXhPYXnivBYH6+sN
sFYiKQWwYw+ZT2xJwDOrRt62DL5Pv0VXLvrJdE+pfZ7X5FlsNIVk3mg5ss0z9zrB
NBlMpeuIXDOqe3TA5bnLlhlULRGkdom7O4lguTRcwwWCVDNshGd367J2M2E8cngx
DHvKwqjLPodous8rMy0wDbI2ebEANvzjOxZBq5VQAhTLUMCezjEDkW1Zbk1MPO32
02G1GsXcyxZgPZHhiq4spSLLSFFyvoRZmJ839GMr4OfUeEVrJrN6Z2UFDH2IXLwO
y8yMvIXNDbWkkC+53OlotAeuBOiLZV913+3rWjCakKgG1vSFx8Ckz27b/TLQ3A5i
Nr0L2hXDZI4J2rL1r4g9KwFdPw0f1sy881sMMTtyZC2KqeC8k5CBlbr5HuDpxT9s
+bvqvrJhOJ15eAfsjc4/IytRGjYU2Lfpf9c6Pyh0a4zFhKmu3Ezcj7upycxfQW0C
0l6G1YA2Cb8DfT7fbZAmS/QqSht2gzv0c5XUvPF4p2MZJsGhUFE1oo0YFP3H+ZNB
ULW0CNAXCCMJgfdCoaeRvx71KHDlPa7TPV850V9m8a+p4yB1WnLWRuTYyFr5Dp4O
3BOnK0psJMu5M8f7EhcbVZolgxEkwx5+2OtMj6H0JAR3ZhaFVZEvwnuFObULVwQ1
kYoXK1n056hhlApILDvCW9azXkv32Q5BK97xy/m3OiEdAJ4aLKvcXVmIf86S6lHy
EJ/nDHC2uZPS74tKil5YyvzfVsKLtphZpp1yIf9htYLHdxeQWgGWzwSafhHA/e6I
/rS6AjicrafAO/M98LkBSG8zcjjvK1h29NoCc6g9EobC4g9dOG06rEpGZoLXSEiF
vdqAVN7IhSGIXfGQtyScy/nZSvVmiL4ltq37CPKygJIVPGZXb4LuFuwp6wJ1YwOo
GgU9I8qP0a9KQ/TiNb5N/0PeyNE8KGLu94ESSbnq8QV2HLmIZ4KCh/85Xp9VHddY
tpmTPcpZQYMC0jBIiCeQF74qQcjVWEA4KlUX4yDV31w9mbIdrM4PwEYOVsgM0hCe
z93pt+Pcd3FrGIdOkMMAPsZrDFZNjqhgbdSdGQOYmM0WNEf4sKbbRZTYB0Xjs5OX
ik6hXzsNE20SLl8/sKqiVzPCyFbh7ydw8eAoKExKaGhZoUekVU5inxAB7ytZKuaV
BEck6niiKExQohz0foXNvw11EZmoBcF4oMPA1GNwHV601lurC2IHrQu4m97A/Yfg
iKn1LFv8MJAJugbRNcIv1jW8qGak3d0DWCJEABebL3YeFfttjNtOomWGftVFDyKL
J01qFqLan6mm3IJgsRpvE4aYPtXbUVPEEYDdiPaCHa6Ol3k3vU2msV5BFLSxltlM
nR7PpZ6ztmKTLCPlqNH8WrrV0iBzOGZG0GbMJ2DzuM8A04wfkO9kBwBfaJMJZLHW
IdGhfm4UQVv3qS/q8jYmRTk9trEK32qjCDYDx9do6JBWePfShT//7ESfScf4Im4k
6bG1OJPl4qsU4TM6e2hqrhGKH0usy5G8Miem3lc3uuDTRfgXhFPr5TvOvSYCXT6u
zdN8bIk+cLC+kEKhmtWk2cNJn1CR5lZmO2Nkp2+Pb8W9Ogfuv51GBknNyif6lMUw
sW8+onwkRHw6rYyO4Eu1gAj//HNFjD108FCp7z+TogOfya0QxhBVNHFABbxlIjAx
TTeo2GHQAfgc5ofEXND9Pj1WuKIqGjQ/cqOAKHN2UWB98+GkFWYlypKM+3ZORDPG
+Z0HpLTHmSUINNcNscBaWDEKzElUX8gtfDrNuEAVEs1ClkSlyeFLV2Rg2UaXbGdP
r+wIgaEwvmpM/Kc2KiEVNRpVf+wZtdLNL37zpQ6APZpPl/Mz+aSsQcd+5GS4s8fv
iwJFj5g4VJAN3pNcxspOwfp9QrpNsPmQRR0mVJNMKYyhjZh5AYmn7qqg3PV+kfUh
rao/TcZci7LbSVrz8wHfZEeW8gGnqv5cWBw3OejL9VrfjQMU/bpsAe1Y4CmMfg7w
7f+OQcChdaL2Picfkac6+MrK1Y21NB4vm66Pm96Pq6TkXTpcj5xQXfd7AZa50keS
0TXInV1VMxyLhRcEhwIZHbE2KPr2/vPhHoRBslqgydx7RSTKQd54ilpl/gyKj/8H
/+9lsgY6vlU+S4pJzRkyWfd05QAtuozmYCU4F4ONeClXgmGoelbiAcEU3GAuUe3k
6nqe4saBuQI4Tjy9vQ9ALue6mO4a7+oSamTZZyyIpNCQOBz2E/6qFzXIsCoFBYDG
4fQrHBDqzNbGUSK0qCfeYDuwArjdYvpEUuV5n5O+G95+eMBoz/Z9X2twLK34le43
P6bqU2kSLbY0w1vPnadV10JmSlk/tay8haagO3awyaaRgAcK2ifN15JJlAd5EC2M
5pE8C3cV57tRfZpMnUn/UhgTmeqKjBIPLzacUEFjxshZJCH+CKNTAExI4r6FJ4OZ
XjOet7IhlKv5Uw7nHlL8f8ZgMei1GqJegjL0IZNtojudanDw9k+xh4Q+USQop3Xl
GDGZwzfDIz3kJsbHgR7/5PyXUsEzILSxqN/THXoC/7LtIAqT1/xdNKWQprErRg0D
upEjK3O/cMrnIuvk4kKvoWfnY70iZExlkRKiSEGmZ1CBWrCK1A92XCztjzWf+HMk
wC+9+Dtgzke2iP0QFrQU7SuXgmz7RGK7avQC178mMdxooELaxl1+8GhMeSTcq47c
hVPPfNr2GvCNv2+hw6EywRSVnCFSbZDRX9BNV7QP3TVNvzp1cfRSy7pf5a20zuUh
/JQ4q9shLYxyPsepjbYX+HC4YBA+QqIYW27oh1bxF1X0lQRHeC24VowHiCNKWaa7
9+pKU8NkEXv6X6l+rovLcUi1Gy/mxl/Pf+aKLhfxRjs/iRyHkMb2vkp6aiZFcvJf
JTmah+SKfpZ/WJfCrtMPK/+z4gHBxP7n+ut/ZVC2PnUE7eiOQ1dzUa19zapkdQFW
ZWkWocgjWvvD6GffnaWfJTbRi/Nge6mtwtuvuAESEcJtgq8G5pssbCylXqR8IUw0
wHFxkp9yIKx2mZHAoieBtBdkTHSsoZbT0ZJhaIkipLx6leVh3hMtmNLZNYADO+pq
+6aNZ+waN63fwKkd8bop19Y9zK9SaDIlLeFKJ2pdJFqq6ANIptHEMMBFvO76mf8i
7Cu1rQGEKk6cp09A+AvliyJTFp4f8JRbrWh3ADcZSLJIDA2t4NLhGMnKQo7dKGRP
grPGXOMTiiH19WHnY+oewXM2kiHNvSPmkZF+deiNQ6XGF3C5861TfEeMG1YEZK9T
mxaYF26S1VyNt9c1MY87cyajMeITe1ZWHmB8nEkSiNBNbUG7X2jBGb4XIdGCl5n+
yz1J8hymA+ynjYTewIi2ILv8NPptMSeGv41Li/Cuuv/l1cP7DR8C5L6fe9cO2G3H
qtMneDchmDAnhoPpdnckIwLnlJxHkRxOSlZgVFc0BPXlTsRLkJAaauTsF/KmiM+Z
l0heuQuJjGpUW1Ace2Xde8Ywipjs7yId/AUQP5LpPMNCAweXSfFMoO9TVhmZ6pk9
fqSHix/Hs5cKi6/kr1qxibYXHEQw6YIWtlCqQgxra6QbUMGyjBynLXIL+E6rcm3K
idi3Nkg0OD5aEYmWu8OK6+m4ypxCK1lLhRtEvPFM2nsvCLyL2Z/KtH82XxFDwq7T
YR1SgS8veo4g2LtgNLFN+5FJpTcUZBciALCEBUlF8+DIb8AzrrUrIgm9Mf4pSm0H
UQ5R8Yxwh/p16Lig6lSE0Pt9Y2hKDy7vEHPCq9s9JD6c4Ff6hrY2W5rWHxZDejdd
yZD+YF8EqaYjJTnTxyWtz3X6ziudXjTcJE/y+0r+uP7U6Dtk5MExuWnyCceHmgwY
FYS8681cAMyh6R2k6upFbfQWas+LRmNnRGnknMRdxDsW6GyBmjIdRerf7JnExL8J
K2Z8UBF9qUEAt8lDDZeXWoeioJhRQh2WhcVWsDQXPLHXzV0d38lYK6XXGxlRNgbI
`protect END_PROTECTED
