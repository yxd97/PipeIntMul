`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bqBwFzddjupasMa1bYirX9Tbf5F75mYn7Cg0a/UIKceN2ir4bQEGo9QK7XPmHec
/O+G0M//AuPyYJTiM9gFXjTgQqQIpW+/8NYOv2kSr15Nzn6pOuwMgyJXRmbY0GKB
0ux9wi3V+X0+bG4wUVWTQ2eTV5tC0XJCLlRRJEOK1rJtqsew9sMjQW3TT8o4Y5J9
G7UIQZ3Pb24Qu23sYNRCexTBImH6G1RAFkhWSjxd57Op6AMcapGMaJsH4MYSM62y
xhFeYSQfjhqtH8H6i1o2HA==
`protect END_PROTECTED
