library verilog;
use verilog.vl_types.all;
entity OBUF_HSTL_III is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end OBUF_HSTL_III;
