`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FzXMDlvr3mMp0qxSHLAegfCYnVSO1XrNztuQLPGuldsk4jp3uZ8zFxgf5wAUF54u
YHJAbXDQXpeUj4+JDvwYQBARKyIpUlANpLgsn3JtODGgpTKQqTI7XC4D9ERu54fw
jFzNemD8dVsMPsi7bJ/85ZvIduBDdvYP5FR2FKcpVfMy4LSxrjd3A8qTQQbPy0gJ
X8RoB2uRm4inAOvyjBanVPmlF/M0oJwdmN5hW98h4s0cZkV6MXcdgVxx6dvjjMRT
v79y6+SLRd+lJESoXpzs+ZPDjkvbnUvQDYCnLTyA8pACZul1/cgw3pSrgeOuP0f1
1/HNu0pEVbqoh2zOQ24Asy1SAX1T0RwQHt3lYKhoewRxuoyxXMgPiokfDemolxVB
MRnHfCxkRz12lp7rVq2vMQ==
`protect END_PROTECTED
