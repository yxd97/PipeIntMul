`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYlONv08Ze1Dso6ntJgvkvYwEKbQyYXhyfVJ48MLdpss4KkjRBB9BSG18HEExGgY
ZAKV8QuRSu05idPXS4UqSR6h0/EzjEaRFTFL6nNxXGbyF2ynpTiO+FlyJnXrX164
pvkaUbNlJpsF3jYOaOvGNX9yi34jc7xRacxnJSDkXvqKTLheP/ioR16uRg/xrYf3
HC9ZqXkEe4J/+ltwLyZ9cRlBto+5+45WORLrCP7jj66cjN21kYwcMxXITKxqraf9
eSfY7Pbwe94R6P4/HYkIxMn8PxVA+F37VywA4FSlUz4yBiOwvDmFAUpMdfULi/Ah
OnYbCiysLPaqsEtUlsww3mnXBPRZ8U0u9gw9U7Sn3wo=
`protect END_PROTECTED
