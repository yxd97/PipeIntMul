`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ePsbIFMAlMYy8De0bU+uisNM9JE6Ke4d/IW4dXrS+YVH0pGBIS55J9FVXWVhhgaZ
Jzha7CUE3N/zDIumUtskBFnjlrMwxDfOAKMlL1UBc4Abdcona1AvO/oGuVanG80P
xbEfUEC+OxKxkn2JiPQj+EgBz+RB6AhYcacGaLM/JiLZ2K0rIscdbd9Pvj4bnTU0
4ot+y6XQ4OjQzwi/dxLSnsC11wW3Vd8KRHKRY+9I7dzoM6uvVq8CmdWSuMdMzRE2
vlfyjgoQfvp3W40GUTJYwQ==
`protect END_PROTECTED
