`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g91Nh4KqaABI9HGFXgLUTZgXsyNjzfwKLWBefMVk64JFoqsFTm6WfYnB5og0Pq9t
JQHRN1oh0NWGTCNhmPqG7IMgKk8q+J5Lsn0N21OJwOw9EbRK/2QqiQWKKZtwmVV4
sv/BgJp6CbO04Mtjnh20hkPhqUbbOHNGDGSzETriSnSPlMx0pQJlahw+OxZSCaCI
XxoUZCJG9qWnw7/iDCJV4SjD5XLvmMirdnkqKtmCX1RUcpJvU5S7dsxftGx0WxNW
vPlXxP8tS0RHtfXKMwPeTtCjvfG8BRX4HD1M4LL038pzSpb6kwylkxepQUgNaRK2
r1BghpzgSUrwhgVktQUdfzNRrBSIA7bWYJGaDBxU1kSAUZfh4O5K5ptyVVyniRCj
yCQrP7N/W3xXuC2C7RxCd1fE1469kAcpVufsx1C1slA=
`protect END_PROTECTED
