`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VoZP1g6oADnmaRQXf9c7bbE7ngT8Zot7pulENPYNzhE7oJCI7fphLLDVxIQAtGbi
vX8Ra4KqXt4A9YNnT33BVlUj4kZqC7nvZ4N/HZNPlpO5HREw8SnNdepdb/PTw4Lg
ZhhBNMzo6wPw5wPfe4QJ9sBNKOqN2JSdw9A79JcZy6b3J4XOODtx8Cw2jcmwVeGr
6HRb3WrzbR4v0bF7coCSrX4DZd8M/XBb9Y3wpC+TSPBqqiQW37K49lkyPWMGnAOg
MbIxsly/ElMmYdrapXVLncBbU88CpGsP9q00/yX0zt/1w/r8sVRGVvhlr6Y4dnMi
JO40KXTywegXx9UOdOj0rFaSKve7ZPCSHuc7FGzX6wDRyoVZN1q4wugpYApiPiLu
8X1IyzQbRtsT+RHXRrsvK5lWdPi2cd4IphiwjTyQW8wg+FZGYiM5urujafQL2O/r
`protect END_PROTECTED
