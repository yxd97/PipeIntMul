`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
avXf7E4oXJi4ufXJrnL+8YSc9MoGD7uG24FmRF9BZQz2OSYhogu8Drj6wl/lBrDt
gCdrGzsfhuglJcEPXg62jGXDAUsZBRKSvp5upG5Zs2a24ZGOcTLJm4JmTSDQL0YD
2IHMSpvsTBfxPX7UJ/0GQzcmhfz+T8CSvyzOhciEMB4FaYgSWKG18tnuYhVO8kdI
2a9hkNUBDny6GsOUvBDWESRwJMSg7ev1hFML+pOJoS5jCrG6xtl9U5zSIs5a4hNf
O1X4QSaChtAPC73qZW3rzg==
`protect END_PROTECTED
