`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgithtrS71KmelAa2twzDh1mzIRrBnL8u0IKlx0zauKUWLzoPx1ukUnAi+Kljs7z
JRsQXz4uUFIo0HugVKeuGH/HhF5gvCfFnBYWJ0pD/zS8JTieKVPIlVZbG1e0BhyG
z96FqA8Iso3e2MY7dDoOoRJk5kv8D0OdohnL0qyO22z9A3NmKzb++vm1Wo77BGW8
MfOUMFqcQT4AVamVCqS5ncXVSLmLMkhpaN159c7dV0L6mXTPjMjBezfKPQ4xoT3Z
weYOppPH2U0kZ+Q6wCenkQ==
`protect END_PROTECTED
