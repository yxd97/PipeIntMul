`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rynZbF1iYNEZTU6gZhxsYrpGvt0gvQeNvZGt7oYKBFVlA78T2XsfoX/evCBrG9io
oksudY5poC3Wa8xj9dwv+LRenc0KI/HfCbz8UDm90HD8jSgdoyvSkpi6eBYC2tsI
t/Azl4ydF1VE3pQcPhfQNmbDucG6grJV/fT/y//ZrXxWsPoGDSgEyMockm5HObu2
EkqPt+IpYy5t4s09swQdUC6Q/UvZ2h2foKhaB2zxeiogqXeZfJOl1RCPCBgx0HIA
on0+SdD6rBgSfN3aZBbLO4KplvwhQO+XK6zoj66m+WpncWBNmGmb3cswIhkcFqpY
FHndVQpuByXK2O+8cyc9yQ==
`protect END_PROTECTED
