`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
434W0BbhXuMJZCk4T3XA6n/jEy+LN5kiKty/7XoAT8RQo962QIpLouO22zgMorng
e2aND/8SX1vWe9h4Qn0kA5+BSqgFAnpKlQKxoABfYHZE3BHgSl4RPERrbDhNyZU6
2kc/6UFrMZNg1M9ra1BEOy1eAk3OeNe8YAX1tMZQM8z30FzJJ9zrSCx4eVFMpeiz
3uxeEc3s0KY+AZwqWLC1QKudCqCoc2SX5bti489aUPTRyh5lJEQsd1xPCoWHlp3F
ZZQCdjfWoNJOJT/yPbLvhDwVfWQkri5BvG2iPEBLvgLhdxOUWnF3owwzuGCXC7WT
vd/K22Jjj/RdsI1oQOXUgrxwCrBgmru3xQudkxfRw6mb38EcdWL7yPY+/LBgONht
GCPo7MTVVm7/b/kr1gf7W5Kfk58Baaj9K48KtfkVN9H3NBYSbiNk8fKMj/6qJ3EZ
`protect END_PROTECTED
