`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B12FL7FZPPF/Rs7Btue20Hk82iBDEXXi92z47CvOJzavevLHTgcE7Q4VNGnezmjn
bRSRWSiXPisWd/6MZg8KT4POZLbkoWC52g9dYMdq3otVgXtZX8aqbxgb8PAk3Rze
wFI5bO+O8PTeGzi+Pib/onso+m28nb9bjNwd50YRgNa2Aopgh90e/G8MSH0BM32F
w91zC74zDGc6sYy6jE8LBY1UPFXVpgQxU0/Dorz5SBgqSmQDI839p7+HUYRekbg4
/XsHsyxaObxOD4wLl/15ZVpTr+8Tu5iUSU5JhYXeYgjs7Thc2K3BRLu30dZhediZ
nYfavdCUgqcARWu+JcuKBfsXzYiNpp5Th/WO05CNogwGbxRHxCA62Yl4dgsTZtO4
CAVFM5V08hQSQzp6NgfksKhMvYTvRTa4KBQpI+rEo0Xg9w1PeYeRLXmVchR4R3r3
JNeOFF7+v3jDjZztBYxqbwJb3otIKyi+sdxMnsZfQYk9NQOL8g3+8XBO7rZCvhB3
`protect END_PROTECTED
