`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFN+SOnoV+yqcgC5dXWhV+IlsyPDl8QpvXQ8SyzA0JuQIG9IxidgCeLdF+sLPbvv
4B4RSz/nnK32UworqxzhKUVjzYvscDjy3LRdYQeSgJ0h4E15Ji++MyNM+NbH/o+E
1qJfZWBu6OkhWEvprCuiR6txTs6WqO5F1qSnqXUwAzdXAF8P3auMXMmIdkBGCDbo
sQ40mSecPCqNzaOdQYBkB+9xPqa9gOLKTdg/3UUgyIM/FOnLAlKz5EtWC2scsygA
GXoDIvAqDgMfrsp7PQpWZpXoEWMhY2B5ZECNIj1sqLMRWEBCranA7jdsDkVlddym
ORwvVXuK1F7VyPia9eAWAMfxQiHRHf8XChbUSr7g1WkBJ8ols2MDeha+MebvqOtp
RcCsPcZ/wuoyFtdvPwF0CMoRSmj1Vvk9bFCXdYOZgYDQjLazbj+YpB/75eNRwZW7
OSAY74h9VeOo4nKZ2zzCEnKxtYdo4PLiUUJTv9YpNiWFQIcovgfLKAcZTJA1fmAu
`protect END_PROTECTED
