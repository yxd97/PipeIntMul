`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KfTqhyv1b/ypHF4msgYNp5I/2UCombW2k6XvvkE/Tco5hVAjhyf3xhhUSgxsyEnD
RkxqJlIzHm2DeT9qjgQcIuyecYZHQ69JTcgNZsrO7xlL3MFKKrU2e17Byo3gWcLf
mGpj1aj/S6SYbF3gZaBzA5Og/Xixmk8EjIWjrtqG2e3yfvMgcACcP5hdgBGxQqiC
2BGMf1bIkvZCZiWvnl0HvvXSAD3J5ev/XRrPKPjUYk+LmwqnPmx8ynYrmi9JJc1B
fdMP0sA4qmbVUDjNGg592800jOE5BvLdwlx+O+TDJiFmPaLg6uHZO9tDc+MrIK80
rRkhpySWqNeB0O2QcNuMnsljZDwNGTYlm1BaV1RvaTiCAN79Dbxh3dxyTYAg6Gt4
djUHHijliHGj+HquciI8oHYp7kmS+4lPN458p4T7oI6ishv1KkDhO5GFJu0voz6t
WRrzK1nCY+n2gNUGtPdEm5D3isvYQMNtXiCQnbAfRzp6YaDyFW+gjpg0wsHW5ukG
ZrO7lvQ17FRp4cJUXPMGj1OPRbhOgx00DoUrbawyoyqkK9Gmqkmu+HEheVG7ANhN
GY2mfcwy3zJgjitjTRMe7Wi9+N6Z/tYtZ2rkf67rMV9VBpUk/6QlgfLs7DKYLfRN
MbzmQJTi5nXy3nU1x1d7fEj+uD0GxXmFxLlZ8vHUV1g0+/NkHL/dxvZObBmADNqk
KzPd2cuzrOL2UmWgWNXqKtmNap7/RSKIYmeqGlcrvPQHG2j8Q36gVDzgzVqESLIF
MPe66ViocjhdLXW3rAs8YwRrvATwIRWLBmIC078iu9nYkUBnBCHHUGoV1mJ5bSam
1hK+zaxsKWaqo2d86TH3ce/K1YhXC5hxNeN729Q71waeVY2xkGzEStiiIdEaOOHx
r+OXcsJXWwb39KdbtcI/UNyy1QEFWsyQcsbPyvcPfAz6boHmWhffpPo0/Va0zvXa
Bw1EpFIm2+YNSTiKVEM3dve66IEJneepdexKmgu1JxQeFzjI1yttVEoEklFlDkMF
EnaPTsSFWWwc920D7WifDBzKWF9Y/MXMwkO6NDWdVgRyWo7g4P8hOp2PGRV/A1CV
z2qfAj5I463i7oEkTGMk0gDBmcPdxpiWq9ltLnrXw4pQOHg/vGgo/cqw6x9Qlztl
EJSYcpFTzWGCooj0p8NkdyvFbUpYsnW6o/sfI7QDiXcwZwMxiN/c7Y+7r9ycy3c0
tPDkkEqQINEv96/N6WOFXEtlbeDZWX1GCuSE9EOG0BVwgPHtKh+W76iyJJ+Jw54h
1eE4cxU0HvMrAbQCC6O2hK/YpiSm7gQvjYLlMjZ78FDpOCI0LdzrbX67P5mqaQyo
ui7R35U/0lZ43AIqRH4J5Ddlce6a/miUVfE4fqU8vxwpiXnll/nKFKfEkoPKqvot
c11UqPB7wB5+5/WeiWWGVA==
`protect END_PROTECTED
