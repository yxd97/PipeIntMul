`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uOjPXUAJbOdfFyvBsNvogUEQIZtJ8Nt2TImukNz1gHLpjx4+Q+5YvfgI6EcMMDEU
cBvntlB6oSMWeC+oAE3y9wLrbqTeKAocrbKmKSL9hytjcbWeXNFPw2jpiTn6MrQk
PSGgmdHm+s+JtghqV7Hw2futkyn/coNX4C/LFv+u7kRMeffdSp1I1QbTqRygZtUe
4+YaohRwOw/SWsmJfPQX4UGukwr/haCQj/q8CF8D0EcHD0iMQQm4x1WW/92EmN/X
t9wyWqTMZmL/efBM9oy2/jrA2C9TmpRCvCRwr+FHufB0trsjlg4VuYoO0FjhKMbI
IuVYAHSrppAdzHT8KSBgF9FtCxqhww0BFTwcAMrgCdxBJavdwltQP9z6y72mxOlS
bgdKiKTLgSh/9bbGEX0s5fvHTcBpNtHQV1YhL8EC/Q81sqC6kB0/ljV7oMqogyPS
/efD+gKSQ940Bo3N7Wdc4r+/oMgkcdyRW81g+6vYl7O3A7nMkVe7hw7GTIw2p/Wp
rc/nNBddNBE3GyVw+Xd86HTupjtztdvIOvxksmjGpBLsoXc0HtLU11oqdcPtldzK
UDgUnut3qhZZ/4JyOSNhECTcWxywoyNQEtFf7m856WDv9Mv2VRFMBH+jTbG70bHJ
CsF/VQ1tfs0+g7hnJMrAL3HfeGI3RWh/9mijsTXQYLqhUl6vm4DokGXrRKZ9/L4B
VFZdBCN1lqR5gW2WXIpmXwGELLmku3kS7EmkAVCff+6iVfJENt6kuaVR5MMQfJ70
wpmYRai2aniNuXxFHwGUrMkJElqupDlcwYxn6ANcNhfIx//mr/nswrXROlhQ5qDk
LaObvUULYChr0uju504ZhvynBA0MZyzmqcR6E6LpXJAM7A4ztdLJ+enQBqlGxjWu
Ydv4VprtsB9Ax3w8BIGLAGOCV9eDPQNO0wi3JIzEqBIOvtGLQl+s/EaMgo3wyXm1
LJFc8lt2M0im+2D3apKrTPkTjs8eQFLfNhDbk35F/O4rf4S/EqnqwnQtHfF2yVko
NTiO2n2DDwqo9o+0mhuUXJ/598WEuoM70QHJG9T9U0E8SpwXfMCJwltQ6tC5pFUF
1Bccm73wkkQbtUcIlaFzv3kR3nBT/ffPN14ybzOuhB58XsAOFCRRgExumqHTO3Ym
`protect END_PROTECTED
