`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hswz2syjxo7RbNhwZfb1zqRw+y/rjxas0HbgkogcrZFeV2hR9z0jAvMweuPrCo/E
CM0ljWwCTVqBr100swArVlbpXjYTREk0QxUznzn4VmGdegWX/1+TE+SGnWoBVlsI
/y3HtXZylw2p81YxTGwYPeD8AAuP5vF28yBfwLidgzY56lUbJiLDQlgNOxyTHJVT
x+mhVKkYhbRS6kq3C1M/Kxc8y7m551L84geAyuLj+GordNF5mZBNpwvMltt2tBGp
A8IQw71RxLIWPQG4kY6/AO1iGnExHV3BJSXzQpKmzIfzpWNa1xo4ZqnNSx3Prk6z
ilrZ30N1GELe5iCXuIp/oZTR85W7q1xMK0dYE8JSXwFv4010D1qOcakVapklKOtv
`protect END_PROTECTED
