`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sRpkrK2kH8V1TkXaAuh4ot9L/PrsTAlqMURYEWiOKv0rhi6q93eFPE93rCtbGCLS
pW7mQEtZychHVZp6JdKOgnUPsr8FnKwW+e0yoYPJfXIR11J3lLLUu5MmPQjFv+nQ
+g9EWHCsGT3gGPxVr4Wnb0QMxJRoQpqwmQrFprmojdxNu7vu84hqGBs/nK4Or7mQ
udQ8tkGtWD81OvUn/unqdLgbi1R5Y32XwR9j4ZVUuA90tp7+CF+CI+Fajsj1dqkR
rZf0aIB/LRd5LOrAVbHufmm1Xa2zRgHzByb9tSy/1kRhwRMHws/n5d1ItpUSGIjw
4kSr8Bk2Q+0Eda5QxeAgwLbeYdKvyNugE0dr88Ttk9fwNflYfkISu6jiM7bwU+XZ
Gc8YiI4c4qNQsPv9Xa1CDD4iKqBr0VOrz3NaG0wS5svk26DyccABdd/2UCrlBUAf
aam1pKBBF828xl5Fm0ch6h90S572JmCoEMNDeYVAZLl78YAfwZb47waEIUbhNyi8
0pWIjeRfLQk9unY8xTp8lQyh/7NwmmqKTUnqb5geKACDSZoZFcyKjSxmqAmAReOf
EVLfjk8DTPXDwbqSqmPX1l1I8MIrXpxKO7YNTP8t/req4mrRx2MoCpBzjR57Qjcv
kGSRKsiVcwn1Nq+rZicPCexGfZoDSWTrweeXIg8AZoW0c7yz+ijKCD05RSzp3Oc2
CCE5IvuBoCHhvormc/JF6cqSLyJFkzc5ZJR1mZzMX2Ah2FpTfPjPu+pxcebeORNX
21RownNUAlY0qilJ7C4kOmncAJz5ydcg2DQCnfTHT/X/4Rax57Wlbt2USciTK1qF
9vCQ7VvJ+HDepKuRaJ6yh2WE0/Gi3q0+ESrdo/jNIGMwE9TP76MNdsc6hG6ipCGR
k8zGouTPHu0Yf/qf+65V84OIP3f7oPFIjU4HLGYyTuw2+PchgL2iOlG7+VqFUkuB
k5dEONT0HIQUY5oZXQJl43N4KKAMCZPcSoQAkxD8L9RpMwCvZ74TikJyyCxKhcuL
iB0Xkkqjfau1Tq26pTuqvhuFK2HA9mlXCS5O1kDugFSaDhQFRcfp6V9lt79qcCn6
pMovKVDjJfDnOwSU1mWFpiH1qST80IXrLjgNcMBXWniu+mz/Q0A8mIJpmMcE4tCX
r5xnh9PdrM7uliJ+2V5caR4TZR1fw/2pPyn/iyS3HjiteHPAefgiinTHNfdAgq/N
Jy/MRin67M9orFtBOn1W18JM7xvZPoI/cwY0kOHkCDBK4NNjCvrQxOo5/qOwagR/
Sz2clyRL8F9rXWfxe4sEndrNJqbsfMMeOjqYUFoV+ugLJpCGnslE8UxfqwMKEsr9
joW7ilNRHfqJyX5G8Y1/vX35QIFd222wH0pasTaN8Nn+8QHboBrqmt1FYdkPnbNs
Wq9Mrrh6m0VXqayiVI1fkuyA+W48TBApADwyiO+s4dXDdih1DlHPt3cFGHQSZzMs
GhCwYk2AUQ3qHysLOOsnwoRaLfiIBvD8n84hD0JOL7fCKlsflNrHpaGVBvNL9bud
THG+n1PZb9r2EnvW+IZ3LkX0P8Jq0a3MfH1ljvpUbW0lkV0PsDGyoF7Jru4I0Ujj
PxEaRpCc6WYIF7t6EQt0N4E0DXCpAz7VK7PB6OP2aFNK4d6pNt8YxVOrGr4dQm2G
1RFrvJX4LhQ9Z7RYMXXamIY7bAJ6p2XorfESVHJOTNjIazRbnDYr8zmmmLLFLYUc
tZO8TN89hqALO/zH2px/4Ewaety4Kl2Q7y8o6596IYDVaJ+pMXzId573JiXpq93k
NpMtAbdAMdsTq+KT7niAF3QBjhQaJFth1PtGW4wHU1YQxPY+l9i6P0zrSKHiGLRn
jC+/SNZ/aFqm3lmiqnrIdZ3kWA1fhPneKKFFehJ5EeH+2c5MoLDdaNgwSPYZawon
YkZ26Mz/h7059SVMEIn249trVSghjVtoPqRONrpuxfp3hQuLjx35TdH4oEhCJaMs
cGxVz0PYdVURcppDTq8x59uYgcGAG8NnTv3IKxd/XvN83rl90UCcyjua5qv32g3W
3eEer4XNe+51Eom3C+PBiG1XQFCSTnfuByz0WgW5pzkObuAmYI+IrzJ/9NTzXtUD
snsn1hUzguAOgJjzloHBazS2YSPkH1yBqqQrp8ZkA8bRSoh8gOqeLrcjLWg1+YaM
YUxV/sliiRI6lE8NgQTkZ/cSNzDuacjPc7Sn7uc8arECq12J5A2h17V3pnnAuFw/
7gpSscRTl7wFG9/+n3oxGFECWPl7hDlpbD4V3gfvtLmxKNFBNxU6dUSjvTf5a7LG
j3Cc2CAF7Q3XyNL7aFbwhp3Ku4iFWf8IBUOocYv3kgZqvaMtv0FrmQC3Go+1nfgL
eaF+bMMAkaMw0Js0MqKz8pfSIdTataecihpHhyAZ00nmajBAVcf414WsT1uChs3k
mPvXitxOAjL5k9urJlSae7OL+U3/D4B/hUdHdrEvxDHSKm+fy3i4OLSHA8Y/AWqL
IcGFRuzsIKMuyK31Gv6ODckhtOUPH5DcvyXGhZMMPsF7OVtgvmTCkCWyUQtuZOgL
tIhSkdkfl4X46Z3XkdOBBc7Ahzu+/czj/1VuXN6WFMqb6oUtEnS94VBZqIpV7R8n
13Q0fpJLEYe6KmwZStRPqdP9E+tFjlySbcbBC0LhCp0RJ80J/f3smSpdDJX11x0o
gqZ7iFos27XZTwTYIQDh//kuY1fW/W2I4x3Wxkt0962CMmOUGg3nHPenEUVf701n
7yr3Nx3uF77xRsMt6/GlIHkwCYm7aC2H1lJ0Kb1sbvi1osyOxHzNLE9Njc/T80dU
klx/XnVu+zxsCXxMG7GNShdafdLpk8jVWvL1AbBy+I21iheW5ny2FyNAf5o5l3O0
VWOMAQeS9C9lkYMYe5CQpScGIGdZY96b6vLZMTRyR4tyhbs9gy77Y2RtJ7pklIFy
g4NW9k9Hxru7X+dVdFKEjKx0Izf1N7qNoJ4UMzfQ3AokbfITFfaqrODpDIk68ubi
D4sCLSuNiL7t0U3BUaS5WOjkvn2MDHZfTHgqoelxuFRDMX0/pLOCZbC7XURgvApf
OLWGbPFh7e8GIIDVgBMLNLnzv+1/Ziz2T8X0oNxMcLvC79pifoxUYAbyHXmiabCj
5j/HSSpNCKXwfRn3/5iK5KVIZL6buPnkATmIIG3+Zw6qh+A9aWFP6i2SR0FFvjBT
tGk9RxCfkmk2TOgFPbmkehecsZ5cgzAA5QI+OD+7atzoBObj9j1aOkeEzl5xVTDM
OE+2/4KoSCIeXXo9Di6wUJfjgXAUvh5C6IITGWafrzfkUQ8jYMm66tI5yrjWFHqw
LQqgC/6uzloEIBG/B9KWshBR9yT40f2gc+HMtmTlODJRJ4JcYUAVdd7ClxYctHWk
Y+L4ZCesC+REJIWVSRZL2q5H+nm/uFMiwNo97dedk346RQV7TLxcs/3X5rfnkE1s
9c6/fA1yUvppVrTspYXUcEtu2xfwbzDu8FTwKIlmabYcCvxOAXWpgGlCBY1McRdn
E7rBNFH+CXmGChBOwEoFVG/zAM9/mV4VP6+KtP1z2xN5R5/LKXGHPNcsWOfpjxkT
NqW7Wpqz/eGUVjj2Hx08WuvSnzY5JZSIY6HFciJJbBPqBHiFYM8lx+KVtOOx2JS2
XynyK6U02shKOhiynXEnvzbYwFO/fakG9Aw21WDUJU52KlF8DKkjtYHEsRe4kv3i
lC+aGpr+ClfcVe/H1SbvFjsSTqxFxSJeD+894TD4xvhLdZ4bYTnAOdRFtDT0U4AO
XUP8WdG3NuMqomt0jN643DTrwN+22hZPQESgGBeyLGBiukR+cwoYfBe980gZ+YRc
cvgly6Z4LSCUivGMHa8UpFjpk6HXd3Bg6DXpfBFl45E77yFF+AScL8KDX+gQgLNt
uNluf/RG0wrXSvBjp3yMNObzR00A1TGnFgRWs0xrjde6VknOfh+aihzsFOg9lht5
W6V/6K531TYB/OP1I17ee/stYdB/ZtZtPs+DozNZKBEPCLdyoHTsZBMYVJMiTdMm
E37JJdcYEBMsstzZJ9ToMvgCzr2UPk82QWhaGTCJQTSvNacBCzGMRfsco3Wc19jJ
cR93/Kp406p2NLfgy7V77F4L3SJh3vsCrjURpoHFNfVkBXW+BAJIs5TRLlowjtZJ
fITk09fymaQgd9xN68joCeilze2RbmKFJJu6QPc4jf2cv4b+n9383CBARCVb6c8o
3LhuZzNxgb+TJtnLwCKdoiUm+gUC69aTPVx7sCmq8ETMbDqA8I72PR+t2dPBDJ+z
J+VYowBKqznIGT8xfAHEDSmaFW3+31SWQ5pyOTp9PVR47G4V2zz85Qe8ENMHQ6ys
vIWQmBK9zXaCJjNHv3UmE3iutYbH/axo6TFrTVLBAu3hYMWtmmGjlXjSorXD1wLR
XPqaD8Sb4shzH+EqXHB3IKpIjRnnzW1K55ObSkKxh7mPKRQn5ICN2Dim9qsOIinH
8PrlGsRD1Ze0PsnjC7w8Yi+JFBZ6ADawPa6/TGyKpNn9MI7gOKwwKluSJaEBMM7m
jOnrLI1vYvES4enVyQnnnFuhbqFE34TjICZUmQ/W4c1kQDdYTNFClRj4uryxOAQ4
rJWV9PopCY862mPBzf8sImfzYBEKo1I3Jc9DEyvvrX63kiU15eJ9JtRzd9hJRuns
CGTMwD9vOGVI1E+vNPQj/Tmq607h6EZoA0++jyXF6sKkxazz2sCNNJJynIe3tqLS
o1kl6oC29uCP32PDbwnDT0lfPyGGYe1hwJoQSJlwdtzQy8g22kUDbBKtaytrBjQd
F45UvLIjBACs2QB/W/fruyg8ek3Vy8927d+8vCwz5BBy0YCQ1WdSBJ1Yo/mfzs7v
WF9IboQKbfqWXgrOw7t8axGxW4btlPtmqlHrrMBSsl5AQYGspzW8fAKLkMD7+seg
ydi32TocsyVZj5Dw9W+o165xesoAAukKVjlNECRy7qqSLqVBpe2RjSDxSyJi3NGr
ZCaszyFHWTYIQZttHmJ5iubzWi+Qd4Vwr9x/N7DgyBQcGWnTCaDGaA4yD92mhVLF
wDVOLDW/DhbhQ0W8zkY7Wa6SHC1pqxDpcaANQUcT2lHc3uFC4WT4qJFlbN5F8vFA
2IUfcaCDoodDeWx+t6BHcu1T4Kz4XA3iv7gb3QyegW76+hAgYM0Y++s9SBflnmFX
7zlE4pZQPOQIaBq3JCyjQv97WiFYEy6IXegy6ievdQnMV7e2xPUT3X208PAuBjmG
Q8iio5WQQI2aTk/uTf1inxb4k6yYmYOakbE9/qC/mP/I0ywvu9ceADgAYWFmtDQr
jWLKOjh0CaJon0NyNf7/pMXy4DOlbXkSrLMW7nYdxBVukc4SbqBXk8vR9KL+N4pS
2HB5Zjkt0umN0Qe67kTzaJS7CDuQGmRArrymducL3Wu5kQrPK9ZSi+H+EW0cH5Ga
qUKGHt4Rbxc9kjcACgBd/TJOsfXriqznE7PbS7jfq1bu1kylEnkdllpOUaW45hsD
4as19mMVFQDp06sLDy4mNA==
`protect END_PROTECTED
