`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HhXIdhTbFcse9do6iwdpRGAw8B39LyRqnctf+yAA3ABJizW29aF+RHFhu01ogTxT
vrFLJ5TWiEW5+1smKiAZgVy4lcp82VPWpBXBWN7wShPSF3B9xF9XtmRLuGcRNkas
oFSzwCvKPrZt5A+gplGNi3SQYAf7/JaywOgj5d4KDJKvZe9jQBtE+/WFYgNelXgq
BdNuEAenFaj9/c+KACgGBLRUBZSSTaJ/9g2u5Eq220pntuUdor8r9Oom2Jc0bP4y
kbGQOf6RZMJz1k8dnDQ2/u6dtZwbaUOr4e4a4ObgG/jSlFYTbzJmJNscS3m2z5wx
ASvDihEOB5dKSaGRx2VUOg==
`protect END_PROTECTED
