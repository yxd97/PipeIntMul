`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Us04gK1aVXJ5+UuqQOlqW0MoiPpXI6uRo2uU12zPG+9yKZC0ycRrKO2/j1iC2Orp
jtYriYRToIfRxgjqbhEnsFsqpoj+jVdBhpVA/EyY+KdVYZdfVDZB8H8xA9H5aDES
lFDoep3IEGSygwvvPG3T+/bPskD9tpo8J/VzrUb+nU3HE0ENh3LEcvylmYxNpfLq
yTk+APSrkHrZ0nXhdvCOujtgzdTQUAw3zw0671ocDadvKYjB6FwaLsEbbZnMMTMy
xduN2iyxCL8ev8qDvfsfetsiw5WnoaJF3zqwyLmW97YF9CHl4kAzjDULnCzhEkSV
EmrpbZHPIEcm2eK8WatwRTwAbnJ4OmSys+YcFHQ4WWPo8OZ5U9wz/zu/r19DqakK
exzP9YkTFxtCrCFrlkbXAaEyhd/HCjv9tnmoMF1N1z0ZPDIshrC2vfCpcxTcUcUR
dAd0Xorw6WmyB0/m2bxqTS3AjWex+f0wDsJeOZUTPKk09nahM0tfHfD5ETovUKOu
qvZySeYZuU0B5fKtCvlfmbB0qd7a7ZnzYdh/1W4lOM/ME9PCmydYEWX3SUqWlKX4
3oJmoIHBY8UULTsLwmb+4QC6lYW0aMzc+y9CMKxFLdsoniK6fFZUkEG5G91hPtkO
fgF56biebEMA4nxMbDmpxlNh7CB9Snfw9wpa7XrDwoU=
`protect END_PROTECTED
