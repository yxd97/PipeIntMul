`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VN8qFf65nSunig3YU3NspLaZR82Th+SI+30v3Xv/ndyjzJtUuhUtw55/SGCkWCtR
rB5Xt1whyrgawAM+mdl/gE8CsSVkhcBGYV8rIVejmIBTM/uN56PCd36K6+YTGVoB
O8RQbocN0b1OoSmfH7+wm2s2fRcy1PrGS8TARt2F67shnWDExZA0g90iaWDBFaMO
GwHdT5/FWrrU5GxXGxuQTOr57Gdc0s54yjd6NZwLg+kzggl5Hi3kwfdWQAytorqG
xtX2Nyj5Tc9il1tGPPjVUNFFTEdLWe3wn/RoZAG6lH+aO92dxGGMpWKxbuPDzDgL
7UN8AtzKcBrA8Pk518P1Vp64ZQWNG3Jt/1HyuBcqbybmmni/wv2+mVjmd0hbo7Hd
kS26Wlp8edzNH3rky/9fRRfo7dpMd1FQdUc6cl4hcJJMJPG9u/ORi0pmMWgS/Oii
`protect END_PROTECTED
