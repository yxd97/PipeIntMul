`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lbW/nHG6nc2xg+7JyH8Lbx2tcbZlBnr1urrkAVpKYcOYx2W94hHeRIMpA3gT0hgi
PvBsP/xhNTBRpVryHk+YTzvmRM8xS5FDqz8OhGvmAWgMOkaBRhsY++fkKPuUcLP/
FI6citQovL4fRHp1UhFgv9ibnn2JUJFR7N6zjTaXu/VsC8lP/OpgE2a6hqOjC7Y0
YFLJn4DxtzrGH3DQHMzBCRcvNdG/ieLB92TBOA5rPWPjPS1e+82M3oFxlWOLeoIt
GfbBxTEuXMVQsluj5S3rS7vaeBv2mms5ekmtrnM93zpM4FqjrR68/bMdkBmJ4Y3z
QKii4J4PVtQlhrt+j5PmSEE1mg38MCXUKbtR54yiFBw4tahQmjoPbR3PStUe6Te8
6Y7REdG9bEnwN9kcSJahEDAn/neWMPwrVjlnrjkLM9QF08WrM6RgysmrjRS14mIC
2gm488GE9PUd+5QU3ARdwCtXelvqI6Ovk1NEByhj5cw7WMKNkPVWdM4pScbNLRWO
fzPnRnzcjM72pgyipY6ZyW/2CVjHp8ILA/R6uGW8qJw=
`protect END_PROTECTED
