`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BU3H0N9CWT22S69mItLCrXyEklc1+whaIasyVOpPoCzNT2tIcvXggImJLWChtQNX
PvQui4mA5emXxN+DtIxjiTTFY5mUmcgrIqgSK8t/hVFPhoHC++OshB0w2nYZSWFe
c2Q2Pw4fRacfS/5dJ77Oc9GFAFrmvX70HgLXrl98/f2h2ssqZzJTXy85DrW5/XMi
qi3cSo8SOycRAO/rKREa+YQ+SorVfzJVEvVk+if6JYEeeqUOz6hc56sLJJHy7h7K
TaIHRLaZJ12Lb+MYBawuzrjPBMwnFDtjLsmSWWH+IBdDARyjmDCLT8l/fCpv/pyo
`protect END_PROTECTED
