`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0x4DFCAvE27Zy3afY6CT5WdPictXLRyT2nBjO/10uDXGBvoGqPgx2zShavzllAOY
rBc/+nhkmiXUiZTmTQg89Op1cUNUGG19EGoT6tzL+AKKNz1b4M2BV59wnJBKI7YV
HozOQ9C15yoAFAk7ytrdX6AOFcKacbTeJmLtcSN2iVLa7UXgwyFRHO9UImlw5pFu
WD8DPo1o2tcUj4KArKC5exypTpbEF/mcNH6Rgfo01aUZwsn9GBZ/Y828dwKz70FV
g/OXFG5UAoDcmopOIvAHN59BTm0UCbxBVaEmC4qY481Aq+VE+hycjsz3F8oYFYQD
7SRIoudHWRjfzJatnB6Z/EyRcw6PZ8U7WJ9/fBxh4ZsHazR509m7wW/V7+W1y+qf
PoyABjOGFvKTdbw+cGovwpZPVtVq9WH+7GJz65L+X3q2fYH21O38INtrw6KYVFXD
GB1n/PFSPUgqqCWs0cal1cjnhsyNBho8duh6NeM1Oh4F398RCZ3YzqTjkBiAukPr
IbwmepUepWH79CRULkuZ1vmGO8TxhqEtZ7v/H5PDQ+5faMNzNWXeodtOhsBea7P2
+JaDKgTw9DWp68Gnxmb+a9gfKLGkACGUjRNArORGQT9Dh6aMkUy7gOIDi21XsxVh
BrlkuNVIF9DP7JNM6DA4hBqvLKCDJ1Biih5I78dfzRtkPUiTUP4iai18jW+Nx7Ut
MkM6lKZy33njh6iJcjIUgQ==
`protect END_PROTECTED
