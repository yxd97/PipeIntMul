`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Ktiljv5RylHrfMwoc1AJZ9jkkKgGnojLJck4rBLJLOAvZPzVK+wcP5wzsnIyeUK
a7pOrChpcatgUlhMtCYKBZveQ308HaqnS20peSIdw3Pb2X+xBqvHa9aVQGxi/qQ1
2k9LRNe//3PPxNOCY2zdw+/9V5OiOlDTUOlCGxZr3j3gQYNAPfaRziOpLs0t7m/8
I2Wh7nAm8yBcjIB0mX3JoWLmqasqv8j6UyP74tEsLgvmHR+KRXtpwJVBGryjqKuv
MV9Whp1zAJpWaR9A8ksNSrvC97yFMJDbO53x+btFh97GcsGcu1YQMRBkKOvYqptI
D7KjKNpcp/Z6AHxMbZrEpVhHp3M61YPZds9oM0K6DkEFD+UIwKaIZDShv5i69bwT
mrNRUxcPsp0U6JEDSiLPrSRLNBI2aLVu453MFTZRWUAgcw59Nd9y/YVuC+dGoVZo
HJA7sbT7UsAnDi/zRP8SC+XmSlB7tpS/wDfz1XH2uoa+n8hwrE3x0Il3TXJYhILP
mSfmipJroh2Va3okJhLMov6WvVSKBvdPjAOE/SMmDl+ab1SgECQN1goW2yCYZ/vF
27kvyIPExgnsT3yUyz8Lz1yxieYzyxqtwm0ZWDpu6e/ch2f713TQAhOtKheEU8Uw
GUQKGZmwPLe2dlnP/WRVb/5R6IeaBga1F2M9y2silGnZqrUiBw/lA5zZeGer3KIc
6ohOQdcm+ij7hf+HOC13VXazlEvLDVwTCGjqd1nMnnJblHHDfZZV9kc3dGUehPPH
yv/niwUQwLAsXt5XBK7CB/JW0UtD2EWL25UgBP/YS/INbh4oH2l5idiMzbaEk1Wd
4Irf+6wzTMKWn4KCpXX2QX3bnUdYRvmCSZzW+qeyQqOhFUzhFLEc9JtxSVDyh7Ps
F58V6BO1fFBxNZMwcDb6yfo9/4aoZvWu7o7etgbVZ3Ph5Pv7+qE/23C8a37qcKy0
+ieIQAROADSQKow4vexzdTYIHEXhTAxFh7Hui5BxGeU+VLYmggnKIq1wgKk9Sei7
sZCEhycDKEkVIW6NeV66ghAbLJDQhyh0JoQ1WR/1LxvIzY2oxeT6hD2lBEPnqwv8
0wDqhvI/6W6RBO7Qyd7gcXiyO9nXIREoOXbEzalqjrxcr1YaWkABVw3pzan0MaFc
b+LrJxuTUoC5hM5dHkVW8Km5GEzT85sogPw7HcqeLLUTLPxDCog3wq35Nl+kIo2h
iGVYYZ/wE8qIpeWglciEiyyen9A4C0x18hyhru6BFgAnHWVkrwL9pDl+vvuCL6LQ
JlOe8WtVsn84rDmi6SfUNwVqO/CaJ6mE9ZsNIsN+bT5fKW4Qv1CHal+B+67KBctD
MQ3Wv+7h/pvIsxQdGtFh0lKh5+QOkAuRBlCqMz655X+ITcT8M3yMPmlMsj6PWjAp
9cO8skSbIVBQ1BtVkyYRweMOA7vmqGPzZysQhw3JqkXkP3MXyVSKwxZu8a8asVr5
xWZWCzonG5o8aMfC342SojcHj1dzb2PGCvRKosB5/sU+ZqJyMTHqae95qGbhcLgY
BugruMVNpNF606Z8N3hPdXREkTHGhxD7rZhveZjO0ad+Ai+l0x+8fcpxrsdBUvY2
UHCJgEE8D8aeAUD7JjauRNBg2K6V3Bkz+Xh8D7+vtRAb5DQJZ6GQACy/PIW64yt0
k3TZWAZj/EFY095S9TDifYTPJ+opCUVR6Mt2I86o0D4M7tNpmpq86s15FAs+JiBs
LwXNkna2C0tJ5G2umNEAynH7flS8d3S7vH1I1ZqwH10h2HTTcfY2xcId4oLppqS6
6/rmr6AHMiILmPyVEy8xDECb+6IrY3utwN/9Er4WxYfwmXW1VpM96UtBuw/ukpqb
ggtNaSrSHV/i34uXMK6XabzEaY9x7VZeNFEYVDkSPdTXH8o6Hf11lqdGpm5dARd8
HnEUBQTL62p6k2M8zt/GtvcvKPFJ09uHUMFp2Jc5zClBB3gcHo7KIyJjmXkZWMYQ
xLwxkxozC3ZwPyHjvRncIml+q3kJPj2jJIOZsyf/sLJzk96qJTCZDVNjsXHNXamv
J2VqBzLDG6yYWaBeh35mI45NUcOX7QNSNRkfBNZlAvyeAtmF6pHdnwUzGuCMXR8E
2rXvSP67D+3H2UORLm9OGxqrfzJ/ttbBZd4fEy3nt87wsaJ6MTRMf4OwLHfH0XaJ
rqsZQWErWSFWYIzlUXgVEm8wQtCT3fDPp2Sd4SAR85gdHA2boURtE6J8ZlnzWBGV
PJOa8s1aZaC1poz7nz+HgaUUPXnbjRGzEu16xChx37m5gXOWpgmBouwdZwApMU3x
5MI/sTJGuD+V/JQ/JamSVR8kL4nOzmIJ8irFgE04NfISStfwY3/hwiFbjX7WTQJO
GLMEzLdPsohuhNJKzRWkcVYGm5edOABXdmYxFnuYQq7oDh7MHyK/0pL8FwA91lYd
9aCkWXR0GfFZ29S1AhLlh9/u6CyZGjEwJvqqF0hGCVYAJVCqQltHBKEasAN5S9/o
pKPgBM1NFSgiLVTkk+WM/ByqPxwaWwCuLaHlBl0agt6doIgAO3/Mgg2EV25M4G+t
hmEn1rld22R6lIv0e+WFIZer7KSm5cX3dDQfcr7hBrB+e0gEzPpqTpWBI7VezvKF
1bYndC9zBGUU/rI/kV6gzdtANASDlC7wnrJR5Lj3/OjYW2PrTFUZT53ihQswcuyR
k145+PMA2oUIByPhyJySshCjWT8qqIz3CmTMxyS4CIA11oPN9djcVTDGjvXkEJRx
5pficaTn7NCLKS/NqyPj0XCT4Sl6pwMQSwnmUIzyw04P510S6SsGewk4WCRBu88o
UKoNA3nOc5jpqAOc9hmpPK4fW/1BkpwQ3nmkGtDuKiljZaZtaAWqfeBn8PkEd5g7
XMu5A6tKleQurcytvQM/zK+HCCO4TiCvel5o6IZpD4EIpoLTz06sl+hJVNxbIzxi
N3cND3h5TO6N0JnehN8u2E/8AD9hJ8CzrRkTa7aIYpj62Q4fz/kcB9eBPfr5pYlh
XxuJUcBmsPl/Wr5ag02TCfQUa7ysJQ1Sa5QsThPrYCudOuQtViqReP82g/stA62e
3H7lBtAHvZFVMeKORBjc/6M6Ft40e0xTUveEuyc2XRtLYH3WTy3AhKtFW6sL6MQm
7wvFXxriRl2HQpCi9z5OH0L/BRqjsn3xutHJExCc9R4ZoZO2k8ce9eLrI4e0zoL9
PprpSparrshJ3725pgnrY42VK0A0nKkuCke4NMdkovyAnYN5aS2qIuluB3gDUq97
BixPQpVDXWfXpG6DMPX4sWx+FBFw0wMn4ptI9l1kk9vn11H3zapYzMxVU0oVuCwW
i/HpND5pMHahWQsJH0UK8bi/udGOXVOzKwjA+V61tFf4uPCNW6hcOoqj5YizsJjC
z0gPJuO3vu2wzHJQmvnVlp47d1C25ND3sBvpA7AKn/mA+XBrbObbIrNcpe7ax6LC
0efwdIq/+NK9r93AmpkXtQ6RvZFx7EgFOz6f0uJlGwZhbwlH+YGo34h+nzaiC/8z
aFm/V5YpqFWkJs36ouSKcWGLbnobSNka+mXSfSRqnFsXxArL6YDBwHhtatZQT0MX
q7oqGXsmQeoHqeCzSX4KtOg6GHgx0xzmbAeQU/hRr/WZQzzf13Jyl74ZwuZL9nAh
WPbQ0pHcab1Ih9n2VCwhp4ElXcdzobdvEyPJ5y2c5efyYFB+TC3cDtMZ0NYddY9e
bAv1loUCPmJYWhMce9WPJJFsvJCmMab96PJF5XK4q9muj1tQ5ujmrs3xJIfPqasP
3PNe1qBv/8RKtP1mLFJ51dQjj7pqpcJUTEQJogOBQ6IcCp+545vqqfVHcFZoNSuL
SxjSWv5hWtFFfpOZrb6ZJtkURXRbGpFCo9ntt4+rOqgT3G9male3ElJOQaolw7vO
G2/0EPKbXJtuhsNWCaza/qtGKM0tvwG1Z34iEDbrBt9fmq3k350ZZpnzDmM1eNrw
Pb23n4/ZY5zsW82KwkcqYIJ6hWmF8wsKZHJYQqqYFvQJIr+8v91G8jmwzwdYifkd
KKe6LOhw3YnOT+vE6cI3tsR1B1iOF4rGsFUVF1fggF6ru96HdoTukJTj04Qr5SJl
MSJCs7+5SbDgraal77XyfPAe4jIILqdFt/v4nIh0/cRpPiia4/I1Vr+bWhkPxVxl
+MqI/QGlxVvDWqTprAFyNgJpkZAwXMVw0ZrC45jd8FxHBmkl+elf7jZmq3gQAVPt
yf9c79+GMew5eiAfdgFtaytWBURFbiLvUyiq27Yq9yxgQqZpUcqQeZWbOpm31XpB
HUJDpwukpOnMSjdbPh58dzo0FpyD+Y+TdOXgd6s+wjwfa3JW1uONOdk6YU6iP4us
fWQksEVbLm96luYzg+aziIe1T2vbLN+mYuzFmTv49YaflS1A36xKpCumB/iqqoUx
EH9k4IF/pcUEneyd3rSmIaMtJj5r3hdoVz3FOitoc7ZVSvS7YbAtSWBGjyoqcJoR
YY0KcE1ztAFygLEYBdjzwZSF7ehqkhNMpUWyt/MpTt9/XOHqzJediP+yJuz60bjO
EQbSlxbdgrTRciYTP7EqBxcsAhXl9I4f7L+O+qOFIMBsthuuMFTRUBPqubrX8VNi
1OT1BPLPgIMmFFsNwoLdI6S8TPFXFn/rCkIesi4gsgbI2d6igMU2z5TqvMH8VYLx
0yawzszahvIHZUguwnWUMtKBBxZXqP3BNOXYMGjmubKkdtmoyu+ZXbLIyYa80kbX
ziliLntnuJoWTmzAxykcZ6SmXQaD4O1cxCgPVsZvBy/ny7AefsJbotHVY+FfboBj
Zez+66o2sy3LntCUYkZ7O/Z9j17ZiuNTklAWa0x4TW+vP3xlV+fQ0gqt+F5X1BVz
Hjkt7sCJsjRci5gYfYJtrCAYmIvJC2snD00euKYtGluLnQfSlUyDUvMpfxLZX13o
3qDpMBGNKBVxXrLTRs6ZWvYCRcIoxXvjXq+biXy85f9Iw2jXZaa/YBuT52wVgmux
0zrCwAVWr/okLWMhNnIKUvh+dDS64wfalkV1WRt2W03OShJ4vPjy577rDxy2GJhh
xw/OdHAFy5PBHyWLWOTaE1AVr9/dLHfchcuZT0Gt8DYCDbJ2WR1ilNwI7FzNgmrF
SVx6Qredgwj5p8Qra71u5FS0jg/JPlWeHGPj4Ls9pE0vWNd6HHFWr21TiQaiU9Js
xU7bzYxT3A5RIe2oio07BVMVwl2M4ygbTccp3+ND1yH0i4MwDJzwbEDELIlEbrM5
8TsOAyqPuQ4P7yL1kzbxAPZKw0BpWZ97gWH7pBKDcmyvnfsBhU/CyrR6+ewNUsOa
KJBhV9m+CYZtF0joiMXM2cflfFCmUoJfFEGP8qqOBijUBwgiDEmOPJ4l/5DQ2c8K
pflOeH9BHLwPju4c5z3Qsi5u2cu/OjD/5NU+wIjxkexVUDiyKX1VZ4NPxGh2BQd/
ercJzbjb/VN316WqL1PwREqrxm+gsutt+ywTOQJRIZQjLvYV6dtt837cfUBZ/6eN
TMCcBx0KibPM9dipCLYK7ZzfZYJZ5M1NipMKGbMoJHPA1NydemiEqlpIzd2X4KVc
Pzek/cGUWu3NjojzjmXxADmKnw/B/Gdhj3Qfg0/DBeyVjpWCj+ntazIVTw25hEIp
Dr/++XXfjGXH3lsOjAHcLhv/LiNZPWs6x1N0d26ZSg7gYOSbvBhjXPoX5azgc8NA
aBboYnPEqzoWiM4Z2znHDA9YhljOs7aWMk7VVAbzviv4dqApcSwyoOyq22N4ROX5
iQ+m4sGIY3NFIB16R2/bNEXW8+XWntrFPUirjKzd8tuZHFJjlDthPHKophDvQ4eq
AfgkjrFpDtzAiuVPAuhvjnU7ihCJ57PkeLw9fXGhiPeFQzm9/VAIA0ILLADajgN4
7MUyNPwevO+Tq7N/Vem6CLvdT8wuMj201cx1mh0F2kODJuCXp1N2fF3BTghiPq8f
XGZqpk0qlGwmslI/2f4PleuNtJIA1b8xGoD95N076nw0aH0z99GM8jnYuPLBhro+
HlyT9EOKaEciYa2WkIF9QGi4kL2dYWQYxpObovCUIHmCuztHDIRuAmMPWiw6zBA2
KbsBY4jOoSBfa42fADOaNCmQkjAmaIP1FXGPJoUKSBC8zpT1n2oPAOdqCxFL75a7
KCm+J6UWCBgdSWrRjK2y9LvOs8yuMpCUNiFFNcJJ/iNlwKQIpglP76iVDny251IU
n3pQ8GFaFs3bY2FWkRP8ZeCP44juuMksxySYAoPZ3WMAvdBDx2Exa5c6jDRs6Qyn
LqX5jGvsMouv2Wko+kNxmIyDUhh2mN+XFLZvqGh0qr+DKp2/Fv8RPtg9gkzHiFBV
SnZXO9qyZOPos9/o7n9cH4zwtAj3jvKRx4rfXibRHmISLiqIO3yT2ZgQk5becllt
l4Ecfy5dTR+qhz12GaRLXN4VSaR0nRLXFxhqmiZ+8wuiIfDkm3gnuntpQE3qbRIo
7j3wvIVl3VO8Brc4UfE2e1SCo9MSt5VEkRcGdhW+fTjG+qsuq9hBiFX3XhF3l2NV
wAs5CwPH83+xetlcKIdI+DmDUiAnj739pjLdUEusnrEfo6jPsydrnsf0KlOvQ9NK
5ClpA4+A1A/IiGE/AWf56zF/X8tQ3oivYhZsk5JiIZqg2iZwgRI/qCrYJ91qDv7G
95FzWOA+1JZA3Ka0YPJddcE3SeuQaGUbr87mbQ4W9HqNTN2e7ZEfWGavcGNyQ+Tl
DKJM2V69Pmv0ti+uevuQ1dskx8Riy0xL6AJbC5TOAX7gOTvAHA3rZ0+c6I8W9D+d
eLCTEWUr1O0+qGeltgXSbCE3OQrkOu21b9GopRL0P8L4sL4l97TcDQigWtXw85eB
v5P6VfqfFhvWFSaG4tnzwi7ewYic13RhGGO6ehveYIpLAT86Fxti7ApBxkzt4+yK
z72Zwirp8HfMcq46Lmzx1l6Q9XrnRkfM/1/np9b+ojVpYqxO9Yp5hSh5+XS9wc87
qe2z6I4FpD4MqY3GqCWy8XaEc9hfPK0WBsfvZAldBMdMBhB3Z/eOeR4X1pvz2/kZ
DCCKdHgF5sgYROpbGPCJcOb54DW3Azib8d4QDcOJGAR3CmdGejN5SrQc1VF92KZP
ltbtbgwcTPXdblg3P9M53NMFbh547nA99QP5i58K/oSpRbTYeOsgz7pkvi6EIdPF
+IShySr4ianpEKIeVW6u+hqwbiEwiw1119Te8BS9wkZcx9yvfNNs+W/ik1gWXGzY
ygEw0VN2xkp731CpI3qQFlSBiGa3tCz5fVC1cCu8fyI0sYxBJFRt0vzdIRWlbuxW
5jU4Bchs34upU4cG913PEBPnZTXOiEwKrgYVN1d3Aw74qyJBKaKKZzPWFQrfa7tr
Hm+H0DEd40k4avnbPD0fOiif//vkt4i1oGZCZuj8O6Lkb4ISTHn/W1r+o17d36Fj
dXc2VR8m58XBRMN++9w594m4uysX6wnacsIhWsaOzjqeFCUwegDxUmBbu3/Nojkh
76HGT/pyXgVi8iq5na64D2nyrOSXfA83KEhHGfzoeZ8nFfTTd8MH/KtIXLHTQuRL
e8DG6u/sFSm0sPyhlf9yUIymIM3zjZ8K0aU0HqPYM81uVJ8LctoLyc0JrZdMngg9
saOgOYW/sKGvtobolOZCj6ilEfmrYBRnBE+lXL/v5wCgQqE2pDV5U0Ka4cGvWpey
42dBuk2XZGtZpx7q1WI1LfR38jCaD7ywlCGJ/Vbq8W1p2IGamtPwEKs5I49/h6Iq
Q+81gopmFbNQBpnhSIlBfX+b1K8yIw3cT+0naFcOvGo9pC10TqJ8ckEccBa6qqS+
P+xJEHyBJXmO2OfM41rPAOn6GgBw7PeWOoaxF9t1Ez0gc/Wt6ITCZJQQ/+YM/oHN
eQ+0/Dyh2L/3qJkglURrP0Y4Wos8a8tkKeTve4ecjySks2hX3CdunbqpAos+xB97
ErEQApRoXeMHuUWba6ksCfmisLogndC1xHnv0FgL8MhryhWoETIMIgjqA8QKJ9Ek
jpQ8F/GVUDxed6sFLyMU5CHjHEe5RZrfc7USndXNdUBl04Zv3suHyPsZimsr4pNc
ZfwxmTuB7DuOpDRwBZyy50DZF8QjDCs7JbI2WJHoEsTture8SpnFQq9tfg9JFASv
ko4C4hdv75v1JhpTc/jtgeYhdSqgx8y9ak1xAQ7MSDiym36VNm1vlDgb0nIXbUhI
101uyFV4lrQC6PMdkqLRj995Ii9Sbc0Q0GjQqjVGFoXzUoNRSKAck88oqNJpUyfU
78LyKNwRrg2Xb1sE5ePrfmCKdYiTBJvwvTIApttK37ZZ4jzM1wP8LT8J8wzZihbq
7oLpJBnjGH1KbbQzMSw/1V41nAvj7pRP1TGeTMW/bd6+67IBOE5ChkZ9/2qx6+5/
i/G6O1NzAVneB9dVC1RoAjgNLwDg2/2KSx+pAfq442UV2q/im6TEFS3IMzKiGqD1
TbTW6ZzEFKjONrMcJCOusKWCzXhzELg8dG8FuK6T5CeD76wKBNZ91bKcLjng+aBU
bgcnPa0HjCK8HdrwmlPgtpukmgrDRt6U5MfXGThx+qdnDem2kJu6j4mB1wDPLx7g
xxh2jG4d91Wh5uOAuX3EFrF+u6sJz3vI5Fk6XQk+fR722fK9SpCEDLOgl4KcABHG
NlPj3P/zXBcQARoDkrC4p6sx7bwmzCZDivK98LfiBLq+Svpb+bxwvjOGBtRyhsR1
tT54lD1vRXk+S4hYc+nX3QQlj6kDA+QPJ6iYjDlLaLm21EypNrIPVi28pBnxeFeh
ioEJemDPpnSHGVU0BlpLKo9u+IYHIRCDkQiABT0ZJiW1kIJcJLhGlrNVhuJCS60c
CbcdvY+PiMpC7Rz8/dXPN8Yvu9DEQRJBuwwzmobhj9j2Xwai1L6waY+1upgNfnNk
Wul+ffRohe+fDnrE1XzUFKOpI3UjqiWDAn2HMAOSn/oEWrcavf1S1xrePnUMUnA2
VL882j7cHhWqG6S6K7ORKT98EBfNjzFPCWaq26BycTUjr4Zn54iCVG5jdYBIKJm+
qEgIUnTmwrdwyg7wZ5iMKxLY6H6F+fm2PJ1a+rsf495PE8GhU7LdRmz5OfiMI5yW
Fu1YO9h0uAAFx5nj+JKgGbz85a0012FWEoMR4vE7gD+ihKYWngOqa1YNuQ0ETu0h
UfAZAeR6hu5gTAiWF6NUMxJF387ystLgn5hYmBIxGJOMcvB1tv95Ej1paRWdFtab
Q2IdWc2r52x9GXPOsCX1dwutdlJEG1InG3xCIwn4Njpp0w59FWZEK/abPThcdqPD
sDflzfzv0c9fRezV5Y5ZbeU1F7sCSkvigLTKimAZFuYL22ZptO8s5nU1UZddVsvQ
nL3GyDX7p6zokXyswTWijHDircTy6elm1Tfu9n79LfbX3tTQDIRpFHrPPwFwYB/4
ecC2krMgdL3S+xJgL60E1GCf5VKB95M+dHkG9MtkGXIAj+YXvkWhZUmehIl35pM2
imXpvVKpSdqHEfu7PzyVGMpNldLs/y2z7e/N9/K1vX/uIr4nMIf7TSK921YvrA/N
jOdAfz3hmNBJAvSg06ByD81SHqmnlhjsbouWBispZ920sl1TXv1woPb0nyT8JkVn
oLu6p7Ygo60Gi3jL7OerkrTrAsihAYP4OJlNKwEYB+jdkJQ1Sm2MCCVu2aSjeUpg
Wsuli3vxe6JJeLylicTqS6oTyLHwzwhvvvCrp3JPcP07jXi2QzJFKy7jU0c5feB0
poecFIr6XLs4t3GS9qDRn1z+vrpqiuC5chq5PbcfO5mczqQPegvS7jexBsAgqJ3d
ACotd0g5iTwX/X7aiwEXhCFwf0XnZ+ahrBTYUTO1VhE3dmNn1FVZ8XU8WoqkVQwl
Rj+8FpXrwrxUfP9bJ1YiVyGZF4HK0v2M00QxkBOOoiPQ+cSG0n5ssl6NGx2V5UVm
5hHl+cKImdtTITJDbkgBqRiAQX3kc4kvSwXCoUSW/vI+gVhU+9tmsKaEY8s3n2ie
JRX01auJldSCjkknaSZUwWYxnKoFq0Q4LKD9zcN1SuVNaBKww9qFisXehVkv4FXe
utrC3Lyfn2dOJTBYbe5LUIirNTy6WAxbfAVLHroxefNi1kYPZGYlJfhQDHV0fB0K
T34ptUQ7mJiozte7N1zuJvHS8zpHR0rwCASnA7a3NptFB5yEB2qO9thPxx+fIQKa
tQBCFpBqjdaoqdHEptSqCM56cyOM7WCivcNnk9uAURD0hZxrbBl7B7UDkybmWqoT
4L+uPTtI5HUY4EDUHGoKVWOA1D5vAsh1WniMY1QKmjHZckCEqmH/hYYVARc44Sbx
b4CuqX6CG9UuwI3jQDebD+5NVR/dNeht/yRzAzoup4GNOxyBwoAUdcR/mtY4pKR8
dXDiOgY+piYsquxMtCW00LauVwgGtGtAkl21ZPtI+nCM7kxZCYOl3Fd+tQzPtbsx
KcVbqBXI21TNUTxK15+KPn/TXHAA61lfeo7G0QJEtk3YONcSLvgSP6XnIK/Pr33r
fMsP02obRYPcP9yKX+Y+bIEkn3qFZFjRkgxW1sjn7S+nZyMR2lb468U7F6cDtSG1
eY8uYueirfutIUzyrnttM5zIxzTF3jBsa0Cld12tUDKx0dggwIDK6mQvhIA9cLzy
1CCca/iJCEABpc+srNSf7inc+kuQtv8y0QFG6mbl0Jkc9fjSvKRslf8boYxuUQ9o
Pgdg+AD0ROoX80rVRip0qHrUB8u+k6wqbSAw1GyA58AjyeGA18HeuHsV9Nh8xyx5
p8L/s6jNuV6+evYe+eEOl23b5PzOAjhap6l33V4zKgU9hlJnDJ0DBG5i3ODdN85A
/53PTAAjNJ9/HZHJe3AmGqiUiJUyAbYn2kn6NU0JqhL5LBhQKDEOGoV/S75Rxaud
j7Nd2Uq0+zqpvEEJEFo5k6lRu8QuvdNhdnK7caReNMKIevbUkkmV8UwYzTrQ6Q5o
OV5+9k2rges7CVWxBvmqL5EmBj4+iis8jQjMWQaUoKXZZpct6EJgnwNWWt2Fxks8
CAkoWRAvH7IluOjJCV4w+jwosQCQ4ryRY5bGmrtfN8VWuWQsc8zb9Z9sy3booofv
xSoHOUk7TdidOA+bNZ8Ovlcf74GahJ0piMs8dXaKr6gz/rnbEKrfNu+Kli4ehzgv
e/nhWaMhjBHIQIfm/JoAoN6G6Cd1W13QvVwubcANxhd0C7Jj1KF1+0wBSeF4mMXE
nMCMBbUpEJ3ApsFE0m/0MJ2HVqqXuO/zdHGcI6RCHepHvJM7oNSPhbOEANuTLcrl
PSLbz5pYn5yKity5DVCi5IdYc84KdF67rWM740OcJkFdy2wU4BKm2GnVDblXJmlt
Pnboi18JWWsNozslawwgVf2ZI6tcJwnjPLhCxgeQpSXIGJpZ55XdQY6Y8+zoeWYW
bIExzW0MjBC97iGSjxEH1eMnjipgtVzERgkY8MTxW8hEUsgkVsoMLV8fav3x09iE
0mE0zijpFj6r9SMVMMnqhfQRu48TGdyBqNE1ybJ8dUkMxAvEJCuSNjPQhsye+XBl
4BxpRRVl8J6QkZ1pfMaFK9KsMu30vboNVfmmsFC6T28Q70CMop57dmfx4HNvoB9R
fjRWQf3ojxC5jFsYf4cW/kZEfvjMGDgl1MHV7mVXVCUUGiqDE/Lf/OyHXBrLUoGn
Zk7SBHP4osYb80z+ai+yllHWTGJvWoonC+wUtOeZGA/tvnFAndyc5p8Lf50YRfyT
H01q1yJxnuuXUtiKeh+wDmSzeQUv1Q5nb5Cxu7fKYFKW9WMS6eVU1NnzFZ3whLUT
YzsdwySzwaeYr6iHRh+0FYvGrHDXhyVK7NKMI0dR+nLufFN4JHyEz1SrC777l183
Ys77Gg3XzzOAK5OGfB5suxvnckTvwEfAunCAB9PcO0ay8/739QxnfAZZ+o6y38sP
ThzOeRaYVODArJ4BqE/Rmv3Cn4ChSw4vYAAsq8SWUL5b4Wwmat+VfqvhCNYLczEi
TcqaAZOmFpPmXIPekUcj3yHDjgUugn49GwBPI7BmPWJr87ME2ridFHeeAHEur2xV
KTsyt42qIbcPS9bSWcyGD5fIIyOgUnaEppmg0Jy0bwjpYYR4hdN+FZj8loa4VdRs
kkNNQHuePS5cFnvEfB6Jmk0jFAm0ELWmHqZDHpMjjM5GpBO84+R2Jhdf0lvLlJBz
Q0xev6T7qLlk0he5zSnfORZofgWWfmTP5L7RRtjKMbPjMg7ECqSH4lvpXtO2AoXe
Mc96gEYMagbgtDmdseOIfs3B48MqMzCsdbSxKtFj/hGoXLUv5lsBOG0ZNFxBvDzo
yuK5x8GvGp8glw04ujNwZE85IIbMiZhqSBge9Fx4Sf5FiaA/+DHKsjQFrsJ7UVuv
gq5re7CVNFtBX1YpgfypnYSNdhmeVn3f4wXjoDt+nCzMzLo4HOUlEQKNqtRm7z1h
SlUPfsK/kKS/a0nfGeo63pc6CkmU9BpzZ5y6k6RqwNy7+Lhx8tnxwwCLY5jfSEqD
peuLgeGIPg40tjVSutR4fuMZ7KZByG3c0rKuXpbt5GuWOybaFbqkZSLo35OxHUgc
fOu3bwMkI9oYWEu6P2sFRGQ41f7bF82utErODY0rDaPUt3te7PKgknrYljwYG6Sd
fKYM6gUjQWf7t/1ffe/fcGmj8TtpULUiD1YkiigPwG/SWzUloZGQx6eVi+BPkL7Y
/0YUpdV7PTGgQID9Y8uK8hs2G6dEV3ilVsFHdnzsnbEu4h5jBxTCkRsiMoxhunNt
Aw7yIblZxL37XmF81+NeB6vuoJsaa6uzNFFK4D1FxFqw40j2U707pe/wAeUsoHfL
OvbrfUjr5eRUuYyGo1GeB4VTWihny1U0d2FNccdt97tdzzTcP2C37FL0cRZra/0j
fF2nuxonn3ib9/m0V1ZM9B0WKJ3E4K2yJzk3JIJSwtHee26PfH7fMdS/bzjAB91u
But5zvxlfXTfSe0nfVStfLC9vthm+nVnbIGN9h00tAxz0ez8WZ/fxiUKnSkMi0Mg
Xh2/0jUJo3cimVdiPhG4Prokpl6LTlhnVwwQxbdBy4Qd2VAS6DG8YyKgb5PjMLp+
bG86oTCRA5fAdkQQipIMvG5ZnBSYXDcZkHMByr7QASXh/WQRquz7qcntPCRhNI5r
tB68hsta5xukck+EMygMUTndTIBBFLJdU53uubsSlhnNAzt8y9+IN9JouFFyaC30
jjbKzb7Z3IO2OUV9HpfbsAyx1Z8nz2lXlExBNSdKboCzCnbFAYppew2qsxaaq6+s
73igsHk8WLimPgSHOYaxFtjKM5w9h0ky9RUPatvHTOUM+tpHZg9ETyMeywDQ5F/j
RcjaNenoNdfi618aeZcSWD00yNcf7zuMhzyDKmCcF8I5H6Vh9e86KhKliuXZXz0P
dlHLlbRr2qSFrvj9SKc0IFXwPOmJI1YlaCyxLn4nIXQklWartFnFwoSpeNUo9cbl
hRsrSZ8gflDakSPdgCM/XyDe21iv8wWE4kvA5EnpAZEL9Epxikqdv7qjh1YGe0M6
pFEQykaaskiRc3IPYXIcaaMRpKOggF35s2Mb21iGf3vqfXHGrd96BPJrRad3f+t1
HHruBKAgFwqmHt1NOXVD30a7+UeBJEw8/nZcySGsugcHD9wZCT0nM2dGhxNHXmv0
GKybYgtzhXGx5HGqoiNuU+ejuZSIJm505W2vjk89ZAqpaps6KN/4nbc7fCn+m/wS
5AmdaeslHdi7cdCo/OYFqU2oPcw3YV7/StAD3RM76nI0d7h9C+ZYie4x2GgAIoBJ
j2wKgGUBWB4pJ3qoBEGllR1SMYkG5l4ceUOj1RY4VUNGHk/IKpuVgEqfLjiUGHvk
3wP51hCQFLYD3UqZofReZ0el9sCyQGGMNLvPdkbyOQ6hntAnfj1aJspfKIdVPg1F
eVz1UxVG87gEy5xSv5eTcLnYovScXynfeRh44Bl7JC4Ptq9q7OD94zcXmTk8etSJ
Dc87Lw1SGMeS72NH6y5LJxNXH0TMR1sVEyBp49DmuJO0w+dFzGX1EmqVMMEvTtNS
G3y/6l+V0B5vn4qto+84jODkRxuKuo/4Mann8cJJHOYQTyphbRf0/9k6K7LzDWMz
gocoe/4M6F3D4EzYDPyN97ASDOc5KImud1a6Gj4b+0mzO1F5Nki1VVd3pkiYeT1l
+EZMORzv2NSaSw7n8BDI5fnAiQSv10kO155GNNROkL8S+nAEEesrbHxNErQO4Gr6
rbeCbYeUBazc0/vK1G38gjbi+riSrtYhHpSZ2jutc9ot58WuEzeAB5MpXf3qEIqQ
sHSMRscYmK6WSBVKCzdboBzExAo/dPwnsAixN882/VWAMVHikxQ/haWlCAWPIlPy
lu+YaaS4cfEAghU1vAEM0Y7pbkvrVTBLDT2B3l9i5v51B3WFDHrt+GUcrSMffrSV
vvhTMv6msR3G+oMaRBj0OREfvLJDZQ9kYbuxDav+gqtSB6bbc3R3lTYrWtodCT5z
hEG4CB87OGYrr+0jk5QZXrwWvpTolIOGTsvgnaAR+1Q7s9xoyVlxHlMOAlFtsD/2
2pKWDfgMTcD7z2HcPm4yWm23P5SO8WkEn/ZuaObLKYzRH39+YKrU5Mov/2uxl0va
jiRnmKpS8FGxJ0eQ9Zlu0cW/Lg/QazqMUsWmf34eW6Z304u4jD1XJXsDtKd7L+Hw
ZY0VdovhXYxe6atPQalFr7q17ce2XjZS1Cf408J1yis+oAKbQ+98o9ZL3x/xZJhI
SgPwo6yyGta4JV3XuyE2X+TKgL0rgFstmZliGAZSATVbjf3owpmYB9xafFmfK/9L
1/2HWBA5IXd22xxnA3UFwVGOBzZHSYYI16TQcQVGcl7rjy6f5K1M8Dn/+35qeJ3M
x60t2o2isPPtj5RFHL07C+lipXx5duobrHUkF+cCVa02NO8hQVAbW6rfHUPbJPAq
GtHr4sEWWPD43o6JZ1A6v/OFLhuCgXfq+QE1XVz8uWtTOznpefdIqMeAB9qgR87f
PvXczWT4Xum5FzQbMko0Fk30nzfyStkhalkroJMcoaCFlKhswrfeWyO01hSJDH4i
fIWi+G62seL7glldvLA2ApzuFzqFFKNYU8V9x+ETeEK6YsX+GSSyL2zfW7Qc+59A
PA1eCCB4B62lSTcY6S8Sh3apscICZylxT/2M7ie6lQmZNGU3GUZBaOj/RnxHO6ty
0JroW2nvmm6BUwhkxm+1KPeMTWQcT0Ks3FaqQtty8SM+ZRZZPAoCEp10rf8d2UMf
kRpAN4tXpy5vydp26xwjMoudiztWQ2kfI9L1bZ0Jbk0ZE33rNgbKeZJPS2kgRQyW
KSz+KLvVSpsoW3RB81GbaLPeFG5Ne3/hsVIDF/DviaSeiKQRoAuo46ihqgfGLnGe
fRb9Bh2ZaF/qdCdGoDFYNmoL4p4cGBtimUmDhm9IUvSoHFIkXnd+k55LpX1VnwSl
mcg8Zx5fKOgTgu64gGFMbugYzBG3iNQNeOyu1BGYcrQwOU45Z7490bvgHIM7xRPH
tQqEVR1IVH0Uq0KHF9aI48FNZkDOZ6KkTN+zgSyJnZNyesqJNe6e8xvgw9uIVu1u
9fQpxWsWf7seFvGJc6UIyzRg6r9yUm675ZHodq4vkyMuN8M3eV/PZgjDNm59+e5p
3TKNavkrSP7w+gJB6dTrsLsWpUj1tFmDtyUTwLvPPL0IYgK1Tb/RYXN1vLkU6dSp
vmoddRowuw59/yaBp7bXjSvqcX83kZj+eHLAMmOlyqntlASwkA1yw+fEy3HAfqpQ
YMwlP0q+ccKRsut2xe4tGED8fTwoy+//PFon2reL/36rVpOlibelBOBdHpcTctHt
ENvkuXHiUL+BdvVnO4li0pKPK2bGJOJCvq2+e0KaTd3ZH2z6zVXPoyJ3yLICOVd6
nZ+xPRCcYN8NIwFlqFXkMvzliH6wzVIbqize+nttjCYPRjFfnfNvFJJnx4/VT6Vr
6kKwKiOF9Pz/iJay/PDp7Jp+fCAjuZZqIZStbJGwUnkfYRIP72RK6+qYInLoN2UE
Dj7zCtP+ZvqCjfZf/4WDxDn13gxsZqqhEndrSIXubfcPLExYVtK+dndXlRtOKv18
QVUsipUeCZ3xNlgF7zRGnpACwBOKRByHuMXWhbywAi6yhgdKPjBgxkhXMdvxU3KL
KOO/2JSg2GGIgfHC5EsM98iK18/3K0xUPSnY0omQ3dBMk1u0KAXUKr0d6llM+jDk
D/4Tm1sJqVt6btAZDDu01+9mCKZSEPK/bIlO20zEZl2nDHfDUhS5ruK4N8Pncq9P
xkOafcjX16hQeKhpFMNVELJKm5Zo4c2qsBU6xlx04oEYFIk2ozqUS21sWvztNnfI
1I2PFuXy/OwZGXz+W5MNIyeG/+fgMmh3azUT1GZCffMfO0gd5mPzXdJjLF518oRx
BsTsLXapqRyKYb2eDFEmLbF4RGxe1br5jwXm8u3X7m32agubByUvhATHCxy5vpDN
/JrWBN1IshVvyGy2bVFbdO2krJTnxyhGI3AQ+FCBDUZzOa9WzyTCgK0y/hs9vSbt
YYdbpJEGTg8Kju+sLC3+P0opEVVxc7fr7NIvKYykXeZ3dPvIoosze92rPNA7bDgE
gyCSqJvPgnAwIxB6D+n4cMSoB3KpcANId161eim1kor5SxiCXi0esqJqOOndPH0W
9XiaSkZPaXEs0itenMXMuvhYyEFRS6iEjnVzD3S3wmhpDIcgIjTSSt8Jx+B077mk
GJ1UkZHdv/Qq5mclN7iW8+7EkITY8Bsaxue85yP7cHaHWwkgGmxfLw4X17OdGobT
6AdK60u2FwU6gJJnYmw4b7Z92zQU4t4uk6nbTbSva53D2LKidvF0RZ0PtFBhuhny
Gqp+LbPyne3rf9ftrt6K2iaSHuntv+GzGhbv98paTNMAfycaiKgCltlLhcki04HY
S65XzJsjAX8JHV6hUMJTjzG7Pp6eji1uvaAOGz6Wn2Ln+ldTSjxz0jkJekexv/GB
RR/v4WskYfj0pGiTVEc0+s3KL1POyIzMu+l/+P/mo2OLGchQ9mcPmT3WkDZ/VwCq
mx4mYXpL0YPTcfNbg1VDom5ibpDn2tLXt+lkV1Tqg6UD8+P0vOHtnk7I83P2lskb
hlIQpJMI7BlNj8IkMfyn1TaloEzy2DDXK46rlgxE36ybWpIhXOUoxnJ6Jr8wYay3
nKeRyUmm8XwMgJUuPzP1ZJDTrNvoZuVEnW2f9SiUPx3OO19BUal6w6h43L00xtv3
/kyyGGElUlqnw2wwua/XCp5MbDd3sNngu0+C74Hz4JGACWgl0Nqc3E99R9cUCd/R
oAy8CtOvA5xIEe9UbAPcHPd5lVmW4Je7jJPyEUxQ3Nd+Bud+Hsn4EtLtcCkw+dWf
oqkV2+IOu9wHP9riTBnkMHqKsZds9JR0+OpoI0h//jcuCit0+YI7UZgI3j6toSk3
mSju/yy6+RIbvoNwcHkKbHTv+pJ2wnBqzA378FuM9mqojMPSH+woyU0h311eoedi
SMQK66UI0JvJH+9O+lsshDjOsBRxEYPtEhJTcclk8LqAczedQfjqft9Dpiw2ABcW
Jp6USiUXPnIyskW2pQjFVEp3CPGEJ4nm8ktyP2wQrlkTg/MSpAHjCQG0Dxj1fug9
fGTboSHMuaN/O3x5wkZ6DnjOlw15ToPkKgFKrtNn2MVSCInah3xogALwGxZ/V8Rd
tJ7SAUXK0dIj9pgx+OawWqZfEXuSlQzkYKinCgFMsDfuHZn0rde1rhVLS52I1zh7
gtCWVmsfqXAyK2Ij1uoRvibFdsQSNrhsLltF4tQckrdc3LrfYCGVrrSSiBAcexsp
c2GtW6V50aK5X1U2tMsz5wJauxVXSZcwp9d0FnCdT+tA6iyzBJEqcxwfwu2SCMiC
HK+ihRTyctd53QMf42Jl8ZjGWalIth0Y5PokcC9lw3XpaNwJX1MHW4H+zZKPYAie
ATZxQzWvT5oRp6DSrq5glscCnmIu0jh+Cqpoy6qPIGBTvbeZkQkHuzfuJccklbk7
w96RHUSV6X6M+S2RGK7Ps9Dshx/u0SeIzJt05aSIaOskrJityd9TRtgYJ30AMd8i
PqxJ1IBCIbfI+j2iVEvT1jf+R2SWpWHMWjG/HmvLGpQSjmaLs11HwhRSYKa1EVG6
7vIXQJ4GvsjDN+Xfigdox2VpsQByxSRoL0aZpZNQtSTzlY8rUsu/tR/z6s0TX3/H
Q2IiOJXdvk/whublJNfkd/0D8TM7zr6FMWQZA/q19fzUDLlA8W/knbmLncGPhOcz
de+VX1PMm1dSW9bRkabOYBMZw4+GxVTycurSbPLpvOUdk0U5vLqxOxKGOwcb5/OR
u8pjYkvRT9KvTm4kY5wQ51/CB0HUdaGEhQ66Ko9fWY++WTohv4Ku4osBCB5TKxWl
Qtr/kdckPtfgdHjdG1JIm2i4SN8v6IM6tulwtpOTSzR0JVrWgyu0xpLX5E6Jnbsa
EkOxXLvom+dlLXSQozLvGk7v67XJuDS100YXm81b5GnTfpiBTBvX/UL9tYK8g3Gg
IlSdY1pBGV4HEspb3yv1rw6Rhl7Eg0d9pKIoONjiQFIOrFSK9/07GtmFdb3/uIYU
qjqdrsv84i5d2tPHkH/yinN9RJKDHyd9RJaWFu7D26CzbABQhrXCq1jDPExCiNII
5Rj0VIQYbJfYyceJAlG4oOinyNGoFxRVz2QMNr8TR4BxpGVXBmZN8cx4n74k+VXR
ApOw+40hY/WuHDS8wPmqyrvP33XXcBWmKPTcWMEU9abpricBUk3JFHZpv2ZgngeK
nY5CGNvmDk4YTLeHW7P/MpFQIWIb3daN/06VrHiNIUKFW6fAc1znYPHSDFXlX717
NOidxrNlF0DRY8OFiLFA27TSysYN8q016NCAhQUBZIQgjk+4ikFlCwISR9RyGTIS
tlPAFoZGq+yk8QPeTTHbK3Brxv0nUXLuUVZnQw0kUXZ4Q9FEw/WsLBsrvqEVmg3O
pVFA6RyapC6MdLDY1l8PEAPkmq2mr9y0Y+Qw6i96FY/nxFazXJS6JOdOp0dQZ1bV
qXpMjsijfOasHthH1nlg5ceBBtB+28QTHDyqawPgotUNZ5tDgTU7tmNcrE68rArU
iVIK1gqygozOfcAZWOuCs7nsgmfyUEsLQn5d16jPdR2a466jVUg8DVGVjcgjzMAD
44M5oaDa6IYIosZto0uQjwcNbvRltcOs7AJy+OfGBz+tCv7LPfhhYuOhaUv+5uL9
I5ibR6+5b+x3QhfOhnmggu1TCwLCIeikeQHCntuVe7JiSWgE3EZSWb/bkiC9SsZv
+RHlUUuFVye1yu+uzxREEtaw8QqY5mOLOBMy5U9nPgYFSjZDDTmz+ZE7i5bmk0J1
AXL1+QqTEo5M0smyqQEM0ckccVAUUnKsd7YwIBO3XrxPkZTf428cauALK+l8zh5Z
y3twP/InCHRB2uLzieZ3ht6KmL4CLNRzd3wyr4crbgDn8W0/D8YL4zaLLG/QTqyl
IOCG93e2iamzvqC+v0rMypub6r8o0WPn4mA/3u7iDRUT9KC6Zruz8RxLX6tTClQ9
rNvdq0zToiOuQu3zjw4Pdmf72JZPb6zHpWKf82+T3jALXgfBoa0KBrJYDwAsP6rE
7t/WiTJl1TFaKIHv7FgogZoWMq3oSMUmqW9KJqgLITqlrL/sNLGBD+2upFb+epzj
NeZRWvtVFLhVfw4rbldZIyZJyTYHAiG3Pl3pkwLbH0BBW6mJBfShOTAJlqcuw4vt
asOvPHmTbzyjeErJXIqg/Q1TGejt3axAjCCEHAXBE5skwOoVmhok/ByarYWEdhqG
PNE9pL0HCiOiJu8FBxdEbNUz03agE+FtGJ5N6NhiYbiYuHfiZ42BJ5T6jVtLozbk
laxMhpkVrN987e7hLX+QjDclCXnBroWR0C/Vm51Cc6YIqp861hPCeIcGtzFvKjln
QZE7x26mqRm2/uB0R2Fh4InI1y6BEuA4ySpvD5FECSr6uzrmRluJ+dEm6NAcnP+m
7t5iSz0f4toXcWEbNgs0pAuPHcNgoC5XiL+QQRZ/9d/PX6xNAuOEMyLO4IUWMXWO
Dr9x5k8a8b6ARy1rstPlqIkqjc0aSnT6hkIyTjuGgEgwIaqS7XrUurrfzVVciu/E
lHbd+oGmjlyJqIQVoh+B/mKn+Y4T89VmOaUq4mLvocqIxyzdpWaBpCaw0HIjRKKU
E+8koc6DwgtB2RNenH7k1+ppEfrQpAQ18pM6X4vsXFMdVopQPD0xt3jVzkJPJcHq
UopahZj3mq5o/UpDlIb0oOZoO13tZi8GlD96uH6mD3+qoXQYhv+x4J9jUiLdGqOJ
yjz5MbkS09Dmt1LS68g7SuNBlSlwc9uMDf2g3CRFXTKQE66yjMftwwJce4J8i8Vj
lkaoNh/RKaI5zn5/TM4Wo1ty4LzpChQAvckcAEy4plONhwZNRrcGM85yHQa9vzfR
538ZC7PGXoYHAJz51YVV+0WqertYUtso+J8Pt1i3ef5SHn4zS7MtxeHcUpl9mV8e
VLRfqqRyHdlLPx/DjaosgsgFQ5bnwinH7awZUsXFXs8kRLv0FKYar80mfpmHrVNb
pm4NRpX3Zos7893Ln5ugaw==
`protect END_PROTECTED
