`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BUzjdzhOmq+eCljELF+SgwsOBK0Jz1q2edmAY34/6dTtVfaTKnIAXHuBWoaaq+G+
f5pQ75U/MkzkikQhNEwBFPetn6ba61NaGo9VzGfgNAKYtebnisyJ8LP+MjRHupWc
quZ4UJfWxpJaKXCpXGjaWEiryFvEHBZlTnKJ1dXhjzmWoiYlbjqgEN6LMtulvcop
HUzEuifYT0sL8yfhn2jTzyt4TLH6MYxOL+qSXr1RoL9nE1E+SD7gxB7IcP077cVi
wyVFehDzfu8jvQ7COC01Mk/sjHvUrxKwRpqOdMOfkgdG1DARzr/+pqo3d+x7c5wY
CIPde+ffQbbDvB05/jV4ldi1u2YZxX684+UeQSrOK/X37WDmjDSXRfBKOwjpNUEV
Zs2MbpqoOvPUSYxoGnn9DGknVqdgEUV8vhHGZX812UWfjA+mHOrn9k1cpA5+BO6e
S3Utf3Vb7zWRRsS9tw99cIIMvf8Iv3vwJqmjTa9dJygGM/Ochv6kubPnG29kwqP1
J1po+8G54VLgbfFzPcRGvVtN7XL8exoAUq3GXA2mPsYXcrk/Hiua0z2yBwr4gFFV
3DHPynAioCpDQRrLfBDna+lFRdqMikJ8QfcyRpwXX1KTWWZ1AjwZieEa4KRhaon4
q9WX9znbyHWsgAzW7ZjiLPpQKFb9iVsmdkqNsn7xyqzdORvc26x/kh/F/W3YVhNS
6N+RqhGnVuH2OFVZTHVVKkZKQQV5w4cTaMFFIOp/1ecQjmtrdPpbuwabypwF/udG
Hgy10apnk4wRzqINbZ6ifQZCN5NrzL5YeDd5KKeQOw6Ik+FKrWuVNCKsrLb5OnKW
DLwHCLCwmDp0m+hc9HIPlOkvuU76fmv91j4v/Iu6je88Vc/FCHERn5utdz5VmJlJ
B7Zc8zhE+mJ+NdlRY0tmNECBLpFCLGW0mNgYvGj3s/GbOFGf64/HDUKOOYSLDg76
VERcLerGyrDsLicD/XoMhzxbZJ1C5SkNeWfm3vjrq70Hv7MY/tJS8UvBu+EBgY/c
b08eKbU6ytdlZrAot2ixgiYAmacL6Spf+wzYtIcThVKUGdx9e+8XLv4DYdZlfOaW
Gsxphr2HOlbXvNDHXmYa5eygeY5ChcslpnjRAWm+4u1dH9Azo/+xLdw4QKnati2J
xv+SlgSda3mYwlM9ZA2wXyTwVBxMV73fhf4piRFZuXZ3su7UwgXdkCdXtZynMnGs
Ws4KY4QItleNnhwP0mZSDjXyQSvfdCxcRJfl2tnNhLQLOqWAHnQaqoZt8xP3viHR
mL73+uyeUScvk6bI7Rn/x4AxKEA2vFHafmB0b3N2FEOi5hg2ZqAK3/J7hZUBJYKU
OtBr2qycpyhZ7g4CruU28X9WiwuPObHP9jcaAGShNXLIm7Dae73ICumeprrztg/a
Ab7su81h3QBELJttRzXI/Sxw5Wox0Htw7Y69PMOwaywARLbyvBouREzD/oQLX/Ea
3Sq1KB0wNvWjSdwjQiWh6DF1A2YmP6JyEQi7KHQTzgYWaa0ur2Dc2cLXmyqKk0qy
FAfRS8VFL14znq53EVwEuKBFxL54A7nQm4xubLkNzY/QJE7Xrw52wBrYEqHNLLZz
+nezV/TetdQoj1CC3dKgLIzkW/+tYwtxg9k/RAcYfTtQk2nPDxNVE5zcg9shZ3rt
XDj4Os2tGvO90/nu0DnSdcFYnrD0gUxWBY1ZuIFClaXoDoeeLt/UTBbKy5533vet
Ga3C6X/Q9lwATZ/tZLXBJLZmF4t+9Wc6sKCgR9vKWWmMlmmEJGJgz1jmxq8jfccn
xIn9NouCSUaf9B7+ZCoyypBc86rM3CDrHnpvuqsiAmbnD4OR+fgWlz8p0Ee2ALE/
lEVyJPXcb2Q1YnXhNBi74c77zO4CIkNqMUCjKhmw3TMxWjr/pOYfo7M5f/3mCEz5
wubidGyK4nLFvmPrg6lTr5uhA5WxJNew/ybTE10nDbQjQ5lklB7B8D3gbo5Ef5NR
7qD2Li6jRHJZYYuyztWfj/A7eh6K/FCukhsi/i4ujb6GkcR+k3cUiuTsZessF7nS
eb4MSzvN24PI0sGP2lBtPcYl9OUKatR/fe73nb+IJupdwKV2Wj6M4Vc0DVKpcn6a
JN+CNKIlgAy0cAdF1GVMMvB1rnZsLwijt1PPREegsfMa0uE3JvUcLy91Xb5Gylp3
Lcx5D3ogdTDhljmSKbnmwpRgLvLIrhxTmjFA4gaLnuCjC9dEzJ8EtUonycqY4hVm
vzpvLL3qjKVJPMnYlHH2pYAzSDRP5bIeByHeuwTVyBTqKwGNI0/Av3BfijiOlZfM
iT4NK/mzJd+Rey41fyTMOZhh50gHvHV9lMCRW+2vGaUXTZH0oC1xACHhfLsNCvQV
jEQQUVeJG07zXQBjavhOfs8sKk+80VGk9wgHlkrLpv37dLJVjKFUWeXFZf+0F2GF
kOsaxXe7vc5sGV2rx39nCdHYXG7pu89qQUcYiq7YSmzDGxAUAFUu/Qi9mXB3FFsF
BZZnfQv8uAOV2lqJIqCGKtbChe3gOfuJjEQqNHRAXr3YM6lkuPaxlkFzjr8Ey+Bc
mw3xHcAjuKglWiuLrEsb29E+1yJmvammoOXhBDaILnTI5Ga5OlZcuLuCMPvzB50/
bRWUCZiVN+tI/M2Ds4ooO7bRrxiJqPUf93RM/5tWeHZHm4EZC0PefHiKX6oXoFuj
L9QRVE45Wob9eUVVBOB39dRB1x6kDe6ja878qPGw8vEvicMMuzcEqr3wRXOax2Gx
ZLyh8x5CLETrHsjJZXqCleUVN2dRYi8C+ve00DhbcrPaC7KkhGJgH8TAOWWpfc+h
oPu0M2uksskVSzYwQY1tqKYC1Jeur2P27GLI/RUO3UTraPj/3IK6ohqxF4JCX+yX
Nigl5Dro5bFYOOr8RyuFQiSVpwsvHL3jDotVV7iB0N9hPa8PLC9y7IYZRQReXg3s
c/ALTLEDDMfWBFJ9bdpbEbQCnKj5LKRki0H1nTh4upx9jc2y7+N5lksBo3dsLmLM
fbAebE4xCq/KZA8HcZlg3ia/lkF9M75LVYv5tHTeOHZP9IYW24OH5gA/AO5Rd/Ed
VGtFGHNGah9mepUe8yzI8fkY3mdFkHeJ/xey5UnMvTWI27VzGRScHB2dLMF0DL4l
wdtl/uOS9t/2hho1rIQad/gvnpG/nvelsg8x7tUWWv1D7FnN/d/nNiZ8APYWrWlv
hTRyas2AFi6DoCIIunYtjCTG3EomXwSHJZPD+rS889Mr4+TBKvkeQFJjINkhU2V3
W2ZBA7XbuOczioHOo0Uqpcuv7GOcL2IGsCdDdWi2IauSdY1l80XJnUaRWAcatZCY
GYOaSP1Aw3kzuvUWn84avJBBnXsZVVmwAGHES4U7QtUqdi0mnuOsYqxsiowqtavY
gQLj+PZgfHbjEzySNditO3RM19zA/iPa1r1MlFuQzTdYD91xz5RsA4W8ic6zIQfU
odUL/sADgHwfSxryLbKW/xI5F6MkR/kBR7zcUQEVtIXQcyD51wAGEQOKaZOZCx9j
8PJMronRAcIr3iEkqolAlk/BTgDDcQC2HFtpyt8vk4FFdrViVcsFt7wbThWQoFgF
YtBhXqid/JrqzTIN6WA136V4AsxRm3pRmMv+8f7wUPwXBTYK11+wIfbEek54TLAw
8IC1j02StB0X/6YjABTdBm+62/HLmye/YJvCCb4JvasyTdI/cqmNdh7akjRhvK7L
4hgdE9Yf+cbftRu4Rm5REPwKK/dluW4fWZitUbUtB/yxJSvKZWuMk0bH1RSAFO+F
LJbWLXIFJBR+h729p0zk7CtXPxx+V2dV41pjuiPFh5r3Fv4EhWAc+5rG8YtV71E1
YQ5b/jeMRWuQ+2qZs0HxpF8v6FJTXUG7OrdGrhwy0l2AuG0MwH0dTuB+vXD9lRPv
ZI1qaFIuB0zLf4sSGMfpmJFOupvG5n58Zf2LbO9SARt1jm/Acu7tlqofBC6fFFX8
dA1PmY6c8yL2CF7eJgxTxHJ/aw9UIijCUstPCMrVlV/h+3x2yWD1XC+o3ecvLXrL
pMABRFiqmn9RQfb4Y6dS2vdd16d60IJ9Xg5Fa/lP10+vxHkrWAg6gxi7c7K5aoc5
rZtRdFlmLm5FLfBr3fGZJbSlMJHNBXVHxhMugswOHd3RoIJ8JiVurYyWeBazWFe3
JrCQTPT3oz+mAwsxCIBX56sQKDBt+PEj+F+iL6Im8Nqeq5jOcpvsQXo46vuWFQyG
ZP9BFJFBrAL+ibRBXfbv+9Zhtw4rc2ou0xJC0plQRsET6v9KP60BJuzAQZpG51Vt
/ZmGLN/+SOXPKuxBkj49yHhPBX78pwuJqbRKjPPccOFKXMpqelKmD9Kh7a6QlI0q
pSguuBGlwj9zRs07c7sd6pILlgC9MvssXHe4YH78bvOT/i3F+O0CbE0Yc88iKb95
/N5988yivut/bOirpoC82yFbmL2PF8WgZEUcMktyBZeSVnZZLpuVKjxulbYRnKRv
W+BAt3dsJUMlM1Zi11egrpQXYuIGJusR0OlTmuAVRFXJdJTsqiQiOlWoMTUVlWic
wLgS8oGqVU/cn4U3a/GSOR50aZBbT2YmO2Rmw/i1npo3sLYzr2Rr48qJUpz/Fh/b
HIfSENVjVsX5wdfAyi6+qjHD2o7uX5LjzEG1oAHQQwR5KNEE5SkLx4Ki8HQHcJrI
/SuHXB+2l7dnKBTt8Frc26hIjYTelImripKLY0/nJ8rTdOIkfWhu2z6pj7kBFIo3
I6426fhcJH61r9AMBIayT5qyBgEMyeERoasrGUW1nrEEk/7QqL6l/bLluyMgfwpy
34BFrhwHw7wX3fhR6BXButU2reqLbU3xJ3+4kRHl8XxDQCkWwiCzLl4ptcW8/BfB
M/AwJjadZDkIk8YI7MhiF5V6Mmhy8l7Evb/6VtcxrE/qoOGTx4pnMc60ChGCr3rF
0L3jpn47QtLF1yRlEIK3i591nZu/qqFveIHEQmYYJZ5tH43G8ROT3tWHYt5pevPR
uR9JWVQ+OeIDHhMg6wWq1CAHUzn6CT+3cxD3lpXpJRMDuj17EQSejOQfVjB4Mtyb
bKRnmauBeL6M3BVDsNMDhIldjf3uQ/wCpGaYC4o/l6z7wOCBJRIyU/c2yLXhPVYW
E4civgHgMPTJrVwThnHO7PgrNu1q5gkPXDSGzQ+B0siRk1PVbx0sFsJqEvWf0yLJ
l8zS2IKsSgx77BVC38DyJCxkFs3pfbYL2tRt3QbYaloLJ8goNH+v/MuR3W6Be8Zu
+FcYI19usqDFkpxNWqIMiyFtlOy7ge2fizirGqdlGICLeRkvrb1Vna0xgdhVrAdo
06bOfgt9ZLHBqR0Vm6EZhJZWcKeYn6pvY+TNMyL5+qQ1b7sA7Ry6JXkjVbVK42F6
RKTkfmjdEfdvKcyT1fXp9TqYflqKZog9h9QKTAktFRACFFmOC8Q3rjrRouHrppzM
Mdp9/a81iR+btWaIZStMm+1MAnIFKLxM2SPraUcFx1DrUyH1/b9ac2ZWaPAmBtAx
JEfJdMUx3X84cImic64evVprCkUExD0HwvqxHACqFcVHLMaUqPNJjRYXs3835p74
U8WSyscXou2vhWtX0CqB0fiZFiX2wevTiYku0nhvlxnnv4SlMV9Va1pNfbtQVLuu
NKAfu0VNHJF6fA89+ym28qfJHVaMOkQnCwnru9QwvO5NUwmvJTMlcmvqX+3lnlnw
AAMyQLY3Nf14k1kjcumeueRETGzm3qszCM46bsy+H6Kl/y3/L/olquScXQ4nPw2j
Vjf/rGpA/43h+mjC/fqdXwQXYBa+pRwdcOKYDuSa2yqbWIUAQjuBg8rOXCvfDUni
MlYoedo6G6lft8uJgvAPEwlS0l9JABz3xXCVNhcqdDbaje0jkRSfwKh9Bf8Hl1B/
OIvlQ41ug9qS/cv4Re6QmRfcCS6PYVhpvyphoyEyToFiP2xBbebITkkMe+iKb+j9
sPnWdj+Y9lQWppDL/obDo6vEWVbu17zM6Ipf48jhhE2enRxzfEhC0TLj+7SEaThN
6pDvaFpIFz/dIwx/nTTGML1DdQg7vctfqXZBNBCMLMYQBdVP4EyJOY3Iqz6uhnUX
atrxREUD37L7ZUkJPoSBr+3kgVZX66fbIAJjXl+1RXm2/q6Bd9I5BR4TsOPYFM/I
fRPyCPQUma41QNGr35vYcTTSgH+xh3eXBSJ6tQeop1bZLmmN585eDVvL64ydKdk2
/4tca5nrtn3igzT24MSYZZzXtougjCW8JmkZ4txHy32s7jXLtIAh21XJhJzNcQqZ
VPqT0YUHY7JDkJzTPSN4CGMbdlYYB4JUFvF9AWuBQ4wIJ0B7hIh7eCSy1jWMN5ql
MJoWuAaAVTh9tkYlJxhKH1DPej6bYQ+qh3W1FBKkP5DyFcOncLGY2AoS4D1fAWfb
XGlDLWNlAP+DRAhBySbk+aHB06r7G53Q7BDLztotUJvqEmrXsh0j+9kf3jFWxN5V
zviYPpLqEmG/xXlkTGS6fU+7DZMJhbHGSIc2o+HL+49okEZCMcLikBe+66kZhyME
U3//CO9Q2cxvH6IDXIfJuuYj5BmW9Nyk1Er+GrB5XoWJQtNZAoQHW3tHu2UAmC6i
L1HMFfrcI0boMwuNNvzaP7QuJ6Ni2lV/hl3hTjR4R7oyDSxOch802A54aoALilFM
Z0GipnsKayWzjm0I4TcnHrSYPcDvT6RZR/edv3OSNTrUvQJP+BgeMzklPBP7M5bC
omZXQda0Vh/7wRg1kjVZhguONJThAzbKmrxfVWxOIoxALpZPN2SUg80ZyozMsUuJ
SVGW44CS36t5eAeBHa/k5VZQpBRWN6/vNDZn+0XNtpDPSfZkbJNS6WwOTGuTTR2j
vbGcSSNNnf50qaA/InbSkP59LD4tUVUegzGPN8YMiLWLMVJ5tbspHwgxplJNAhhu
FPs2NOOpRMH06H3JxH4duH46/pqbYiuaw1js4/d67NKGW4vFuAvg1di9HaS9V8Sc
PaP+K+OLGKzO4cO7V5HkKHCMfpbplmQYzMT+yc9hM6/jP46+J57Per0wCdArzNNt
48FFbUyUiMv7O4nfrdLso7m/k6M0EMId4l/KbE4rW6VyiQ7sXSw2elvWxVBBsi/p
VgahLdMizyK6ydjWxx6gIoJ3rn3Bh9QxBcLHG6yJ+CEaDsDBqz1jLtcJ1Sx8BVK8
kLEG421VVLQBtsUHHw6ZpSUyIBVvmWe6xoBdBwzHQFE9x8SocHhotjUYHY6uKR6L
/+B52YwDMV+86R/Dat/8FD84Vb4PeqEF6crbyRC5jicVQ3spzJJWuTu7MDgofMuj
vx1ulpOALz+fpT/En8ozXyN1y91wC2oRCS/x3bDo0KXJwTRHVEdmj9+Ayg7fRbWX
Vibt6baEuT/Zpj8zMx1OuFaDHHCO+/Rk6Y5DXVakIvemt4LljdSPEbfd+eXKwS/N
uKJPYkye1LaGenmtBp5Z3n9Ws4umJFPyhKHrWW3nJzbO/t+ZVQx0ipgFttjiwkdP
Fz5Dc2PfRMVRjjy+Ukth7KsM0eENB5+QU22G488+6Bpi8nhCzqar1AnWPw1iNI/I
TK5HRvJI8tD0RBCStn84pwKcUuFl2jknarGf2K05yh12nSvgyJRauWw0wmAbzZN7
WwSVGy6i/5bnh9Ix8fH6GLKXZtJT5bqu/Eb7vJ/zo+YZMD63h17Y16nN4tEwrf7s
6f5i8XEMXjWWy5VfTTX+vP9oQW7QyJwnu/suQUN29l/AHD5H9NlsMyL7CnAIRcKY
gTgA3EWrooW7CV0iHO8DWxKZBvNJR9m1x5ojhkVRd1f6PxYJm0Bagpdfse2AjIDv
9x05esByzSZf2JChXNaRNpmDqs6jblhadFHY8KZWPoJwWBzzZH3aYsLBWm4NqJDW
6mXAGgYjfK9srQdGswna4huh6z623ugnABkK0VgYl2S3nVpxdFbO3THrfxWPkl5J
569Sos+T463vdCUSCyyXVSlMxMHTXkHVrtMnFXUjmEWei6eHJLRMyCJtDIZYsXW0
m49O4rDjB7vnNGzKd8yQnTU/SZp9T8EyxsDQ0NfO6JJg0aR7MJ98hm6r24Z0yd2f
zpXbkR0mloUl6StGY9rrb4XjsaaJk8aGMj7Ggeef9fQUCc6NJVj5iU0bqZSv4k1J
vRf9aXFTdxltBIogUkOfmCyjjTk5krsFzz8uAGoWEkRCqfiviX8xLdpFzsRMGUGc
2cDhqCkjnLnAEIrnwS2oVgmHrtnbGunWhRFCccn64fSCPhb/VTDApyXAXmdvxRQu
gwadp+uEsDAUYEZa3K/PN8z1BEJ+EcCvWHQ7gEmkXiYvfpvlkxU9L0LbuYVxnT6c
Nb3QjPk88bOMp260koXZVSX1SUF7ftq0IoBaZ5o3zkyN5X4OJpAkEya4F4EEB/gN
zHGcti5du/XYUSZJDWSHtDA7ykyePmmcKX+iL4/dXw01xj0weOtUD11VWK6D1GBd
zyerHE9CDnN7DBimGd+Blc72eq4bwCwSvkMSDNwPhQ0H8O0G3Y+d66VxUls39rpd
6NCDfciVpXLKe2+5Kmz6+D66yYpucpSgF72usxRZCCIOGMJdKVV17KnvO1wXpTAw
+la1R3hs2RIgDoYT+l+YB5go4q7gIyXRWrhPoM42TEq5TwPRYfrl0/qJtfiOXpfC
l4dpqEUFw5G0x7RwQcJVtJgiYFXDsq5KI66izH16ITcBCy9FH/JXh2J68wvnspdx
478jslzIhEiZmT0AhEsdbWQ+oBgXsRwcHS+iB2Ye69HTEJA6OHrDFTh1IMDNpTT6
JhC5Wel4iREo51s/on2LO5Qoh71VSz3F867SQVc3VPJXpIKpsdnr86fvVo4lbdsN
SRS0dfK9odNcokmlAhULH7bgfmqcwCPhgVM2chQwOAvtTnx9GFJaLgUfzlBE6zQc
2G4hV3kpdiHLGKjhDiqf1q5Ki2IjanILUIMsH8qve1yJOf7aoISXZ3cPjl/KGz9a
GDRhjjk3f5JfiTSO1Q6ouNGRdeQrvPhTEVAPB2AHNdw3N0/e/6sBEu2+vV3PYFZb
72Ypb8ybnUjFSkIN/ri65yyc7cgajct7KBcos7RkgVgt1Zt1twI9vkSur0uNnBiZ
Mf2psrna8G5Rx2T26nBt6ma8PTrSvj1s/zC3u7sZMVJ4z7Pp6r25S5nkZ0kHdINq
+6B7fAFWL+Mc6ZkRL44hmeW4IAiq0G7qJGUAaaC4qZhNbneJb+IyloYj8bSiL4GF
rt+tsp2TzIPxKGdloOaJ+VS2wMHsaddk510wbaKJRHCoGNzfooBQt442MLemseVr
wpmczrsF6TJnmCuphNen3uT1FflqDIF8LktxI9f3g6Sr6SdmeOT6/yirS3rRwAco
WHHLZeZfUoc0zpjcNIfc01iXuDkvh/8fobWEhUh48wvad0HdICVBlhxceKsWKCaH
axueFCy1HesiRYad1KaGpftYdmeZCAT5PezkxaBQn3aMcZtuLOOjmwo7qVKFmDVD
rft5XiOiZ+UmHyCFQNdav0RZIBTvs+miDcBG5bR1xQG5hVV2BSBV+QKj/y1ye8Q2
7aaKd99+vL7/4QI4nrKqMmWavlSNwoqmeSDzYtGg45V5NH5zlOHXYgG+H6QfDfuW
XoqQEnY1mSm7IHBZkRG7uPxjeXhQPl7ufZgX9GUVls4yELTislFtzpW7KxHpvSLV
oqmBBehMF1JPG1qY+U91rdV/cCs1dlF3OHA11QPVDqa2TVPIEunUPsxZi8xKjrH0
WPDhsj1dBy04jvDthr6AUnfQRN4vnTRJYUx+91ltfaB8UeyRINMcdKBNgZcJHb3P
F/LQReuEjqAeVlz+60UysEL2vLPmxWvBT/GN2qqqDj5Nc3GYZ0X3kgQDhVw2paoN
MbwNX6yDVSsDXNPiDJo+D7NJagIl5y2wp7b3kLPcVFLPE3rp1u7jDXLIR1N2GZMJ
KzVRrb0sFHBn6Yeomyq24+5RpEpGqxXJ/BvcQnHOQeygMT6IQfKXxG7oVAW1TgHK
/3An99xd/xlUIf6G3ji7giYcy82hzp41CehSyWbIkrZPgUZK3XkgRUtojrgq/+5f
yAsHgPPmWG5zY/Umy+a0Jkib3JL7dPCBBfF6hU4PENd2H1DtfuOLcjYjhMh6+why
F7QncPQ6xukiJcrNh/Ih0f70YBGMTM4rJMrY/LE84f2wrm0sHb6y8hdZc4RyIYG3
/8odf8r0D+KPrnvZ35rGTERitLMulOOdR5Vo6DTy1Fgx6U50rbwlGqeNdHOuxlvA
35hHLE+reKcWKdoj8cbkwGSuEHHvSkUzmqHNHMKsIUMQ8z4Hm2hwH6eI1NRAXoti
wYutO+CssQqu3W/3yHXbm7wT5CVFNvzG5u3RdlEhvaZtjVGh/ydPzU6RvicOhJJU
W5z+dEQsPolDgbHldkeNfL35zZWur44a6G07jWj8t/GvN6sLLiUzKN3VwtiAbHZ3
L115Qx++jZWqEutj4cofjoU7fjw01HPkEXbbstOovTEbSLyFaE5AJI82V2A95tbh
mG9eqnRUxNauuyAvUHFcone1n26jqE/YfcLF+StHbdwi2nVgHfKg6IOdA9MbSGpy
qMu0gYe28+WOV9KGC8x+9LdeRQmT48uhVgOD3U+t5kPSeWROVDC+vCe2XM9jheAf
KeSTeQ9m55M4D3xEWYSrOIFvjeX9sVM9pUQlNGbdrO3vz07dDKgLVTFH8nelD6Vr
MPGeur1iQwE5Kp4ISPs3ot5oDhj8IR/DEjrSswFhc+Y5be9UEyIh1LAXIY3OcvMf
oOgQVNCiZK1q+CAG8mf9DoD5ehB0TJvRrUMfS6zF5RKTzzyZaE4LNGa/zW+CRfHS
O9uyxiG3F3kKoeYwxaMz6pY2FMD8qeOHrm4MaDoxOGudv9kvJdNzn+G7kWpUzyJP
OpHod+fN1IhIuejc8gGBvm4/cIs5QZLsXlVu54GjU+v94Z5G9K111CNNRxWyVhZz
x+VUw0TVujKzZUdXCK0m4tNfErRahSGy9gQCCkhg9dguqd6M1LgtK6oTD2t9984p
/yRX6cctI80m0E5BinG6BW4MgESdsw/AuRCTr4rSEvMGcx6TzkDfFmWwDD8pkCnr
QrFkq+Iqoe1v3vnDdZXNAbEtv6BeUeGQSDbh4ZIZljENR9qs3uMpn5cNRPvok3H4
9V+rJK+CRM6VHXDtsIibwCYX0jLu3xdogHkBTRpPcDiWP18v7fHELSMHFe/2LBls
7jupK9iGMFrcSa6M2jIOKawgp6g4URiEe/h4b9elOMKAlaaIOt5Vh2a+G6faB82G
C8vI4ZEFHuP3nQTrdsULC9Ic6+n0JyaeTWad4JNaLwNsRzKR98OKsSRefB5kujh+
WVdoF4xSo5meJgFT1khktt3SFJ7yYmn+q5Ss38CPwfHY9CvuKCRsGYF3xQNzUFZh
Jht54t0nzRjFR1nF2W3uz35P6sjpDePc8OeWnAvcDvI3bS7RHGhckUzLut+idSVb
cVF9RNYQHAKBX+Yj1OCD/pcm6aXtXHskYspgqAXUTgF6sTVT+e0ZXfCYq+4L06Dh
ZaGFPyO7MYgXepEMDy19uDz5OIG+M1+0BUo3DUN2gMRZHGnpL9FW8vBSYgt5UgVW
a3cE4NmxB8GrrlsI4SuleK0f80v0c2cKp53HevmicOw2lzu6KCZIQ8vIXH2oy+R0
wZB6gX+NzOAEmZkJL0yze4oWN93+tXuHaAKCH7JHM6aMXPgeuurwzvPu2TJ9obyt
m7Kma4RKIxFroTt4zftpzLJ2+7zucK+vAD/bYnH3aXeHl2nLafSncYrcd3rNzCnG
UotOe/FvJ64zL9ecdEf20IlOuRbvKtOVvQyEEvtHl+hienpOlFaXkRuFGBp7r4Mt
OWQfFy96hNZ1fZUD3h9y4d+eZ56gj/ucnC0Cun3PVITv/SHD4NjQN25Lag6c9pjg
0UmFEHND4Fp1ZYt724OniMBGhOtvLCNvlV3+UxZtyl8qlczkrtuJRXjVgnAIffml
rc4lacsbdroTCSF2eaF8npB/WmRN75D3GHgiDCEu2k3RKU0OePUWVr3o8n1PIZCu
3ZznGnZ9Ru+/SzXNFI9pY/1YJZnxGOcOf1Jy76sQZnojZM0U+i9oFVNOiohq/YTB
ZfiLFeHxc1CBydj08WimNchx4WhCCTN8zQcYnp5Od50u4UquvL9HnXu87slRPN1+
njh6pj2HEi4q7PJ9Dd2v+6S3YonvqPLu5e04sskG7SR8WrmMD0kzikk29UO7bvoD
3H+tJZnWL6vijiHTRXB1AyceYYMblds8zi5zrLlIf0+a+hzu7j8I5Ak3YEOoCFhN
oItA2/lNYWbsXnK/RvQejtvLZ6eD5TwX7nh2NlwsggsbZg4R5ZFr2NL0a/CnN2vQ
L5skasvmWsfXQk1wEn+52XLAu3jVpbIFh9wNpKZIutO98P6ua3UPzELU+oAePyAd
6a5Xs6M8Br85ze4o8FNwteuZA+lSWREfNOQLHj0JsnKwBKFrooKpB+tkTiPJwYv7
MwZjoE8vA7QKATdMTgztbqt9xe+Qt4KYkfnYqiy2F+akRPspgTvNhoBTC4vBy0ux
13IzylFptJylfPqHruHtF8g8aIKQdb7pKzIZTnPoiv8tnUrPJXKwyAol/L62Lu/M
0IlpbX1pupHgn1bxVePAg2n9NqGBEKYzIk71CeiW3vGqOYfgcMXPZVgN0jHFH53b
n7oh+LeL7LACWWc+pstIxFfPYOuNxMaHch5c3Py+Exupr4YfqPH1sw84xXFwz0iV
GJv5tQNMKB5sO4scGeTXj7DCV48FWQXQcJ3o7A2DQAVXAYHnjM6es9SOqX3Qnd+g
2k+J5xS9EhV2cOmuMkjQ6LdeIyMI1ojy1Ry8wAwTQpI8Sc8XcSpFWGcyKv6KNNRA
AeWfbU5hOFJFg/Uqv5+k+C5k4FxtufNqPT+artQHnfzD9vxFuFXoCf7OSaxrTM5l
5+9Oa3O9F/RUg707Tmr/o85iBdw1LYmLWH/RYf/NOTSri+qdrmAMkWSeLnoAa27j
R7Iwo5zuHk/QrcqNPQ0W4Yy1AwQwuYb3qPyVjg6Zn2U+bHeWxFsWRMsRc8zrrhLi
Y6jhZd0U9Aft7oPAs0IX7bRqLKW5UFnNT1xr+Dk/6yoy/JOKrd2vQJADwXcEpZPV
PmmVG+oNvi5hO6CcTNunU+syj3aULNJv7yEE0Tm2j5P4HvgeGxq9KzZAAGtX9dkA
nZfzEHnHC3dDp+u8pz6b3D0HQMqGwmescOgdNr74TS9lCrv6MbxFz2Zfk1bdf67o
mC4I7qfvs4ALNV1gbBPDKRF8DSAC+O+CGnEZmhSLwhP+V/yh1XUbXO/x2gn33NVH
HeUc1iSkBRjMTbNPx4gAa2q/ICzUeTM+M+5pDhtefOL0Ic2lmzUWeM+2zvViKCQD
AMofyHBLp9i/LB1dzCcGIe5L5USqqxpJ2C+aFs7b06PNVI/1lP3JSQV9FkD67Ls1
gEXZEfV5wBLk2LFDArV40zQZMEfdY1UoseV7R9eXhmGnYlPbqmZdEgXc3erRyOlc
nc7UpSvMsQp+axyYEbqjPbgpl3tBHfPkFe0JEnz3i0doV18LHU++MaAshAOpjMTJ
vITGgHinP7czyDyXAja6xCRb6Q9Xiqh7P1Se/qaxCvQC04IGPum9m6EtBbbX1fRi
f+u9o3obVpOzEVReDuDFoQ/TzsxdEY0Q5MtKruw8vkqiZSW3Ge1TDSF7FQRGnLDz
Udp9BxOVmtjUDeKNLb4ozwgshx129BhbsT2+NBX2D4ydcA8scJgGqJCXdFoW55jg
0eZuToB5DazmWJPnr4CZYd1Fp3pnFKrnDXeYDh7JytZgOZx91M6/EycgrpXAGWAL
2eyyyRr3Y4QvHaSmiCZobKDEV2lxqBBpAalcvfJbFZOXxeSbsl5F7mHpUfbw+GYw
ZeRq5cOd63UHOivtXJC7h/pmhslnL1eMmdpzQ5rCJjLiOx8InOp29nNaahXMBS2R
ZJLq/4eSQnNjDQFp9hQY6ZyVfopXQaVkWrCwVWShU/MwlMwtTbEiTay56InnTVmB
T3wmU02Y73iZWzmVojiM0xtgbTtsKWxF9YbjWX7wLREuuvgGq5oLowRhUiLXTaWf
i4w2kEPaZw+jpJBNmKr+qfsAMolG/+Zod5/y1+nS7oDfzwIxXQC1gaAVtW5fDgsv
yt3fZeW2pr3WpzEeyTdJ+uDmE60m+KuJV7X4mxn0Ivwu+bGolNMmWn2kGA6f0Meh
drW+jYEyUykyjTlsYDzSCixfy59UloNrycblbMAdNWnR5L9heOEhXiKNDqzcar09
1yUrhr1jZ3lO/1Nyjsj980GP9i5E0GX9iy+KLSUqHCBsFUVcFP9EL/cs75I++u2t
hcp0MmNGWw8bDaEXhwplKnc+Fxk0/mv2lCCGsUyVMEEmtpMd8gkOcAhcucsmeeOY
ZZaOkM0tN60oFLKgKQPLvnhdVDG34lXi4g9SwZKFbCozY6xT6tLzzsg9GDiV4amy
ERR/9OmopyffRvaERu0gQpC0Sin9BiZQrl+x+izgRc1ov1UK3JgYE/zkfEDhRMEN
x5s0ogbK/5BrKePB2P+FGK+yaxLSrc+0Mpj+eXo5Asjk0JtR/wcLuDuhgTgdb/gr
LTF8TY4CRBna0Su11jLafNccBCXUMZk9LH6gCq1IuAOoPfHGfirCKsdIxozzl+xq
R9VCKN+wVcOKSB2semw8ALqB/Nk1CnNPnMLC6XXcmUAeIMJa7dCtIVFiVEOOhw8F
mGWta8WQhkNkZdXtPzyx4kLJ0aKWvdpA/++6GngC/2Yqt7PKlyo0aUhK+yr8T1mv
SdS0GkjUow++T0kf+flsWFEwB17qUIPvUfJTqGWaEMGepXZY1nq/eLjPWmdUd/Xi
M6/U8aVTUhPfc8PPuQUEx3208IRDmoU0dM6NV9B+EJ+F7sllnomYvvVu9vThG7ct
fFbE5NznNscBzw0IHnnYsvxXj6gqprivLrZblvs8P2fhwU5oYEbuwcUJD66RnZkw
598apZ65ZyYpo6aXe6nUITB/cp0CnT1edKVusNY/D1aV7nyqDPAasGjmhknvOo++
1cqfsCE6cbHc1aadmz0ZqrfmsweGqFMfQveAeyDQAzAYoTgmQ0ug3qcI8gb5mR4C
3wX6uHcGONz3voia+b0/mR/j5xvyyIP0nOYsrUw+V+/iHe1Ppn8bsaD6vigO6b00
lbhHPAGt4jpP7SEY2n3n7wEj2DgZy6848VP6wDkb/w/+9CWOEWtlKnJ1oPmOIETS
SDuNWOVR4QdpP1RXhBiAbpSv8tL0MvVSLd8IS9/Uyj845V1l5fxXk2FcpDIm3P/y
xZCQBhj4lxCHm3a03n42KcaXcAIxzOWjDATpLVg+ilS2Hl2En/LHfT0jA8CxtIID
mkxQlqyj1OnFC3+dv5vMMOEQiZyt8WAnRGk+W14cuUQE1H5ZXNTKtfz6AXe7zptV
9YzJRVifEuOsDjwD+fpyReQXBhII1gu5sfw+pTu5aW+WmfMKSU9moGbal7njOFXW
Kj6GJLMcKSde9fyfH0Yz6hEJ6waU8LCCWA+IxHt4nYVSxCzRQ2ln7goOx5xS0HYN
lsIwD8vOnjjy1H/O1J/2DFW0ghih1KuEBDiuB6QsUdfGzzRBaX+hdCTLUTrB//SR
LMQRun1bXLpQwMjD3kO5o8qU0SrEGlCWcakRPHRYcAc+L9DbJ3v38z5//aQq3qsb
8d2LdDE/sCHqe5ty1d1KZDndpFfoGfYMEvzUKocDKFYy4aRgui8Pp2UqxO6kABwH
fQ4NHT39EJQscbMtV8xCryIkiulI/5NPQ9FcZutHH+DsG5we3+LhwSEFYa9cdzPK
DnW2tf7fCrXtPVXt4FoMauKMlQmfWxRlEblBaHHd7sT/NstUOYGtqnnmxLIQPFJI
QIBt20axtuXaLgAFfPORMcxInVZGO08BqI2+IjuNVHQUFAtj0FuR/HO746/Z18Jd
0zuzpPpg+oT22fd4Sj67d5wAukbRpm/D8YpLoJLhWPzlKxVfkNeEUyStw7AY9F4+
ABtH8U6mFkfBKjiOd46M56vaivHbUMwKtYmwYhEHmwNGUdIGLFC3BJ1BYafYE4wH
YSIVCAkIiOdZG39nSWvJMdv3UYESsgFao+rsF1dWHr0t+vYJ+4tMIPeNtSTHgQNb
z0NZ2FyViepMQmzOwW2NI/Q6krm4UK11jOWuW7X4KCVcvyslc8ucteDMvVWsZCgi
bBxN/LzfoklroHHP1PFQ+DDmAOYbKuGiWx95nx4mrHfOldsTj3RcX6NYmqAdunCE
y8qr+6ETZ3lyAmzBeFlQvSLm4awhTBlFR1QUTIyoTPT00pU26l7ciHpJREw7KBHQ
GfgqUJ86mNLy0EnUMkj5KZfE0lU02O532HH9Mi4lSG+R4wehgw2HhBhijaMeRkuY
aOdQgXNJx38NIEgk5VqdEf4KpVIctWHNj0gPSH4Veezr7QYJ5RAYtNm99VjpD8qn
xEUvMjS78CmSlIt2A0uyqaK++9Uv7THA2bVjo2hXVAw5q6DCBNiAEYMKn8Zwf6FW
pYye0ebEPeP1blHjBg7Hc9f8Lsgu1NXjrQbPEVjP5I8F013nHKcxjHCg28CIUWut
2S9NXylHUDxX0Cpquh7NUVPNGUPtEAa5IG+O2AESx+u2wapsidD3COJNHqz/sBpM
zhxiswbLPa10wZ/nc04rV+Y/UXgg3wbrdZoylh+nlm0W5/QkrBqWxNjvdVjo08xM
bacgTXv+Xym2nAoNbXDy53dUHf3z0Cs9tKc/moU9+1d0x0JmAW7JU/U7R6A8owzG
eO+nFWPcELcSEpENAV6QDRWhI59dDjCbOhof/OgAh/5KdnucfUDV2v087mzD9E+R
V6E1pTKH3DmxbBlUz+Xyfyeoj80DC9y97B9BsMw2OTgtSSwrRCXBlhHZP42M9GMM
bzNBlAKBWS6kn9wM8sBqoWioFvkrZXdo8F+uAogu2QL/KKvyuE2Ynj3zY9oK++UY
V3VeeaRwy6rzFysgm4yUV3cufGT6CT2gXaTaphD5S5fvTypliJKqeXXlBlijeSKm
/VqftFnCUTLTQhByyK3l8qXGJy0+tHaHhMXZniK52l1kgvcURw2fw3G69cIjuFIt
TNedLj4Fr9OiUKcOO7GCg9NyF2QcSu2wk9dzJlk+mOgGKzR7MCmIf6IjrnG+cW6/
TU75jErsPzEV5VSQANVOQuIWLSctU88ecCTUXeo7qV8sRBAmU09tgSH/f8wE6naH
JSvqDx8FDRmCnv2SQzhsdhy5meHL20TVYo4p0b7HKKYZsT7myERt1aaM9GdqF4tj
1tQ1QYRQ26cizly7TkUaUHLyYRvNpWlNG/w/W6DC/LsSZIe9NZToQVgiHU7FS6yJ
Da7qNyx8xwPtbMJpCDTTp936VrVl4AcQSt/m38FJiROjaScy+Txotrpuy+5I/Mpw
4JGzq2HgVLp2n7VOWRit74jWl2BPi3qNGzoNzSZvBUsIUTBrAsWkrSJQspNjceLr
6xnAi53sPaRMS8kAntlWUd3C18siuDFc8ZEiOs2/zwm3bWrK0MblZjHGEpmMrtom
sifCgzBGjHJOJp8AujYmOYCFjHad3WXGcqb/jf/fxd8/sK33QElXE3125N7RJxjd
zixhi3GzEuHGgnnT7D3pFUZaSy2qF8ZnsUbjXDAsq3lPJ3dsHlNblUMUedToD6YR
6nxrh3vQlxucJqJ5+4JP2i0ZBY8YZVOIrlzEEYaJRZGIsN7p+pSac8UkGA0SVbqQ
SBmCtSqR/zVWJP1soMdFhi0cPKsM7lpAUQdYMvfhUn+VL9wY59CeqCMe55RydyAl
W1nVZ7mGJpKvRdsArOLFFuKNYArW+gSQcaO/NjbpOVwk10XvkVl1Qe1rO4MlRLA1
SpA9nDkjsnfktvutw+nsBQymf8jXEIn0JPeZfirIjq257knpbvOJ2cvhlByp1xGG
h6nDrCidI9ph6HK+R/7ppQTP5FG25FQ8F+feYON0ww/CdgqXxlYb23+7RKNKNbOv
Lw/CFQiOPSwtAD6IGwgRp0+DLm23VLWIinedpp+93Z0/xfylkTu3zsbRZqsOezjA
1tniJgafmNju626khU+iS/boV3t62lj226EXo08zihtvIpidrYF85AsCPAukdsUB
A9spFgg9Diwdhw9P4u1ufgll9Km3um+8ZR3WIOrb9Yo9FZ5GZEW8rMfKpQYfNRuY
NzZPpD1lSycBOXCjC/lP6EkB0U0AUOSLuHq838+Ehe+9BZF7cufPqTv/o9w5meMg
G+ECjBYlKUL0eUnq+v8eIMzN1beMRDFYMP1mcgplAauFzJpXub501R2ikvhl7b2Y
b8fAwANpcIIfBTjZGhMmheO39CBb2uiM39M2BWFcKlYR+TPzlQwQAZm1QheSAPnj
lRNYnnahdhrpluo+EFxACxEUXEksSaRv2VddwBS9O4nS7kP89Ixx+OTM9uw3gLd3
QepC6LdBINtcEz5lLFn8e55f7qMbL0IEmjiYOwQeTW8M10uX9absOIsEeg6Jfq5g
kp7lP6VaBD0cRAKgPEbs7UKoab2Ot+n7MOLFhKAifXkkXL3K4DJhdQoNJm4e0CIk
HVZyps3r7rAaSpOktQ2Hs8WCjQgEScI5rr04OQO5DqogOcAXqPXzSzBeQUnTKCmV
Et0k3VV1xAEwMVzZ9YcON+bPt2TYlVWmAjW2MS4I8SMhz0fMg6kH4FYRGDeK8Vfq
3bKT57oNNg2IV2ULQZ641zizMct9Mp2qhYbr/MlPDsZkHPYoMvS+epLRJSJLkDZ4
u0VrJugBc99Zt7IPUFkZ3f3/0EFCodSQMimNqkdj+/ZHu3Y7hLMPjUuIh1hWbIYP
WL13nc1c6Fo99sRA0tGkXVKfxTY8rKWbB7Nfsf2FeOOSA3NeBoG1igXd/Z9ioGKu
UDvTMWB3Af7kHQqO1ttcnA06nZic78na2xPVQMfnDKWNhdu+afbUeaJnpxXzux86
hJV/PWmjmi7hrXgM//0JbAgNT/4IIcvZLHp6mT17RDL/QdmXYxoLK0/lUvelzlaZ
jiFgUbbK59gkxxa9ga/gqnc6xjpTqdKGD3ZA7r9VPCtCvb0oevjTTfzxFGBOTQHR
3s3LcB0JXqyAx35VQMmzQcPrxNiQ7ZSnXaiTRVfPs/2YQfAsxOEA0yQatMfkAeCV
3zs+Bz0XgjKQD6hAJluJiUg0BCVyyGSuf9qo6xcT4R/c4ZNBcd/uMYBmrwL+0La7
K2D67KWyNs1FdMLbpj6423ZhYsr5Z4jIIFapKMvLUPBNmr0pdS2hUMfSrnsvymH+
XHtJ8qouUe1gPkrj1vDXXJACZuqXwkFDKdvPeYpoEz8R3AETW52KDLMUoyiozn/w
X8CSMmANnUYTTOlg4oL3FdsjllFo/6NTxcNQkUaq3ZUfOD9XHTLFLBZjpxUjAYDE
stMKK6ZwCyiT0roTylwGtmifybVVBpv3C9X0/t93u650sMGOXb1wBPkBGpWN6lRm
6NolSJrf0cX6iNCevRtzi+K4r5UwiXd0XUiIYHhIo+x/8M0vHfs3PAFVRIrS4Z4g
6uPRk0xtWTLzvuNzUYLuUvFVZ6DkPWJj/1ukrO4wG0hsuiZG+TJfx3UefqDd/J5Y
Z8Jwrl2hj0dP831yk47zIUdxiHBLXtDtUL2jKE5XM+sCCjaoK0CMrPXM65eTt3RM
k9czDFIiU+MuVYI9mvZhL7VNtuR1Q+lEBGY72BHZvcwYsN/XOgOF18zlNq4MZtbJ
V9Y8qsU+LSx0Z8ARfoeseD/1P8G7ZINUWUF8CcwWy6zpkzBYekTWiWDDy3jweQOT
rctHv7/ZKw680NiKhmsIRGKpRDn/tw4p3Cu/SOtbeqWPvYA+Iy+iyAfuQjAz6LJX
6RiG7SREWONNnoYMAMvXCahfZnWaNvgCOFIJskwIywGiSNrgOlBY95cfdu6qrUev
Ql79Zov/MqWAJ/VcPvWu2mLakpJQ3/LZVelmvHGw8AGiuzM4uWtvYgpecIb4gf62
24nwsmn5kITWrsQje8eMGu0nW/RaQbr760n5uhnQ4iYsZW0ZrAHgO+u/7QVBS3wt
UMvNNcDIrRXyzl7m7jqNfx3vwuBjhCsUcb+UApWuD8YhCOvN18vUE4xVOP+WtvZt
/H5wxaGJn24nqgKR414uxVayaF8Q9idEB+h4HmH1Hlb9yWdUuF34CHaOWSTf9A9x
OxEU05mMH/aqnZ53hwKnM+wtjNUcenXAuedUiy56rZyWz7LzNagBN7yEjbjd2uoV
4ar5y7SdNeu7xV3RLsGIr75K4/IdIXngCro4PafLow8cTEHYlHCwigubfQ/Yzs+G
OjoQRICNvFUjwmVOXHHdfJ5keZ6wQHdyY9LCZogxw1HQVhq1CpY0B1DktpDfOoFF
AQfzQcWWixx0SstJeUoKZvdbv9UVPwYkF7zd+2eBcGUt9U3gBA7JRwnJg+0RrJGu
p+NggSM5ANfiIzym6j864ekLwAB5+EwyqjP40uU8hvFXdyya2o8DlrEhSxON8uW8
OI2TvN8uLq+/8JckM+N1IEi0f/IxKLdisrVynVT0Rvy+UF3aKtwWj91nOI5Ah/wy
OiWhZXJpxUBdDhn9iWaScIgK8/31rR1+tca3yDc2z2CoST2Hvg1iktuRWV+jq2bn
1B+/DVXMwcUDs0Ngv4okEHoraFCsWxcm5ZcyzEoGmtPCwZ5ocQKglOq9Dzxjkg38
STKeH768/d+9CMnv5Hm2lwo7gnlHHJYPUHDGtKxaf0GFD0i4oBbae8I27Xjjb8o6
vAe2ryfJku+48Da9Gk/oLu0y38vB1XwDd4pGWDXwPGoVdpYKWNP6MMLDmjwVTdgX
a6/KEd3Y6OOjlTT77JMqEqvfxVeBp99yIQagAumLGMeJZ2/LqiXq8JVjMAPSEtH4
p1TfEak6MVu1XCuqUHdyHE35oMF6V4s0lwdyn3YQevnV3l9kAH+JAq51HIiRtif4
Zf+QIbdqMm4X7xtjeRy4gU58dpwT+08j42QGYSDLEISG1YAZy3z+vNgkwoOL3cK7
rkBNSb3rUNHhu+VXsQgulS2lw5xBxJJKI5KUFqJ+pkp6IP2tfEwFpQ6gUgUcTAeR
xGocLdp46bdltA3LmxEq1sY9rcn5dAo/ZtZajYq9ohAhVSCIPndPltKSXdXrOMx6
9DBJIop7AivvGJ4ubw5re8OAoQSXM7W2mH35vR51tvlzxRgI0z6p81aEDYcpxkNL
D1Nrmv/GeN5D/0hAy90OBVNsaFjIzNfDuR0yKLDQ+3Oz4HqxTiWGs+pIqhMzHss0
kGCW9UPPYlTGzel10AO/QUPST7T3MGOQHWbujn6gR+FGeDpv8NvjbxNQ3j/xv0+G
m77URVQainvs8yQAdVbZpmzfU/XxOi2Xg/8zBORo1dtMh7tqCyTZh8MpaNDsPUHF
pS+KVqgrX9FXB5IZQwelzZIbt4OKI5BlRbhkgTZC7M+hw5cgJ0L4ZMfTmMatsuvx
j7EdNi6lbNLIJCFIN2PIEeWi9SbvTXBQBDMqoyPgDWnnLwOx+7+veOKxKF7JTt9i
u870x2bu+kyy6NlkNo+htFiw2wwZRIcwtP9W7i+yAINbZ5STPLrbJXzBPEbHejNr
Tz0znEcKGEzneVO+KUcgkXpMcAPal2BqNrR2Xevf4HtgZJPXPTzTnlYS7hpHSYST
uo/SPp2LelzOq5YAJ7/DS30Ecls8cEhnZOqbnILaUV/HGPAM3s8p7p8bLS54m25Q
9od/gbR4iY6CINhtawh/EmgRPb3QVzgYYVW8bSk3rYGxd8htYyjBseao8ZS/Sgxu
D/6gVKFdmLSGEFgmwgbgJr6HFNhUrOzYbS31X2fS2ozSLQRYUbeRZu4uOoiuvqd4
xr73h0kGq3YocYNKRIgTCtlU2dz1ZV2kFVydGr6B6zcSx8cKmljSjxKPoL7Zq2m9
kcQBrPjch1EwmJ/VYkPDkr55EDXcPvqOVp02N4AEYVBPJKbpsPD/WF+/mzXqb3+z
FcBDl3jybX6jWAZIzegi2m1G0j1iQtHMoej2p1fy+nbhFpt10e5CTo0TWhXXmiY2
lXBtP/9r1U0a75cwa5CzFFBu7XbCl/9LuYqkHmbT5E052RYtPcyAnu5funZ4b52S
8AkUyURka8GQTmYyaFJy+DcozaL+PL5JyN/XlctU3dYYr2mgTsWmfj4Zg+XqEFGa
3AyUc05W8MLEiOTpzoM7XkQ2l5qz5V8yU3UijLgkoHuPjqDb7Hn2VGMnb8KvXfvf
eNtC+M+0YzJdSO7Q5lHydR3V3c4l6bH7QDUR6ajNUUzA2DCCqPYW4BAH8MWyX6oG
59Khd9TWqE5Z4oxRBtIK1dz+zERbUxt4wXt8bb3EWxott18EXKptEXfKkyhD0eND
Npr4VScHYl3evuKHX61jmC6G+0e8AyIgyDvxd/+DeSAV/zKcW/+7sDgIVwopWPEJ
aAUtuXCIVUelMr6Vx5v2IT3u7cBxOkl+rc2qfk9CJA76sIRKXW/g32itsdjpBjMo
Qr9Cvyr0Zj9VpJBYA2XQaib6yEBtTdzqznB+ezuz5y7u/4YcCKO+1uugGJnXWXZv
nyD3VL/VGCZRmhqECaIVuGfj8D6SDFUYiFH6kgg/3vRDJbl8oM26qKQ6NgLwpQC5
Z+aX/xyn19rFessn5OheEddjRDVyYLosn4P/3sehTyT9JW5j7p91OF3wO1Y1QRes
EBEVJXgMYg45u+dhBhTwTGrzug0Zm8G677E9mPGoWqDrqkc39kEJSetb7BNwqMNO
gM3SJupXzxMXlNJJHXR70Ixph2YqMKJYQdRD5wOjc/qMMbT7oS/kxuMubuE07rnd
ZRL25BOchVkJPm+yqjCAhYsDrGaPR3iHB28W/bcD8fAg50Y5SOPiw6NB/op3uWZw
IXsTy/Vy7Pq1Ql2vNmqdiQYmw4HlQfz821hyDxGNhykXOZaLUdhaDOhDcz4qLG7o
KscQA3T1EnrJbIGO1qCT1fgM1kyT4BQeCU3YYEqRf+MwrN25izRQiJ9il4wODYqB
rkVe1C7vweMdI7DUaquXbSlc8QntP0q62lGLp2Hri8Luki3CiQ2MxDxo7i5xzcjU
u7PDjrWMg/Ml+B8tdFugO720LpVaHa/h0rxLyH/GlFRQKjnoBw0FBAKJdp0GyI3V
U+ojOBdqH/MTQTtHZJygQe2gBYSBM1wMrtrv6zDtpNxpQ+EXxIdJ+Rz/jquA13Sm
X6/jxuLyuo//uNIN49s4qFdTQbzPkewsSaO/PoNqbc4Lg+veJMykdrId1c78Le6b
B/u9jksIw32APO0zUpn64hNEiOgxwQtkSMTUQobvmQ3K66rN9RzEmzNTZLk9A4qF
AOEjjb7tYfwN3aTaMDN5F11enDGwRT9F6kNyxelnt10s4tepES0BU1W3mAEpYAUY
FzFeuPKXrJ/PlrrM0I+dC6CIYJzvEuWJ0EpZv4eIeYdo4SXoKxq4W/uCsCokxiS7
G2OUOZAg0+l5+yEMhP3wCV3TXpY5nBNgcz3rVGr1mGtYg6u3ReL4OHzPjfMGU+3a
C2N3a8LQFEQmz4AYsKU10axnqm8uQhvCQffE+L57u3cx2Ph6HE3DRoghzUzId1H4
T2Zq8gJnhybNkn+wvbaqpLX0ITHshkxSAdux682+Wm6GN+l+j5mth2olkZ7Dk0F/
/1NWDNsAcsKLgG9fQwRinfo3KFU2QKCH0nJ1GZvIQihyvyNRXXFcFNy4kf4zGFHB
ISdmiKeornNk5fSDiH78DV94ZKV/+CisfgQYn8kkXAPL9rJ9jMcJ3wc+bTp5mCXS
NOudRfPp0K2EF56Fv2EevJt14kQFio2q25HgAa9dBrTHqNlAhd0pguTnIozSc0uC
WK2KVjIeH0b4/4oCuL3Cvcp8O0Z5+kP2Ul1sJZ11+Uv7VeyBH6cBd/RTXgSEEGlk
hEnCy318eQWXmn1txfS8SDmQ/6sq8L4KWyI2DdANvHiL0gCzbIIJPSEARBSRY11+
RX8kEt4FeuGf8mmkt/9KVuo4rSnnYrmnkEMDDN9g75i2Fybor+HY/kN8yeLTNqvm
PNfn1cs1TjIZ2ClKMohmW2D4Ko2aAMJ9RpMvfJhvnJSLeo/x4KVKxKBwfgsm7R9s
Pv1EyjejyWpUsaYZy+F9QCbo0N/5Qmru5/JtQ+UOPuhVZ5aN5a8W5VBN00WvALnR
r69tmqykvFHoEgEniM9RjKfk33HBWXM/ZPzuW+07HtiEZnBHuI2/1NPpY6+yvCOT
iqNyZR/qcgbHkGwuW4xCHSFj7MANQGXVdroghtcFAqwVeW9xA4BlpTeZ3jPhXU9n
HLHW4+zR1CwdDHxYXRjpdUmJzZcRSDI5yBP8ZtfkH/H7oG5qbLIgpj3cpxj/lj+K
Eax1X+5Iy29ds1Ww31i+Q9+9yETkOw4dpTDr3kiNANnojT067ksa13ZxOaWEw3Jd
dlsJEjo1V7GQkAf9DhtAdKsBrrhpPEKnkYi26de6DFBqRDqsjYo3Ve7QGKzG5PEP
Z5gvtva9y0v189+6vFwBGuVwvEBkd2yB45akMuofQFkwvxtWKnz6NWZFwgKSCd/3
WuIekFSZb70kctmzb7e66tJ3rXBYOBYgtQzk1cWcD9bPPhcZYgmZiO+icOjhIXYL
pv+GicAHeqp5MdRewEuO7cDkj619qq6+ZHOLOL3JZUF9cMw2p1O3VGfmg1Zcwu2s
ys2OBU9OuZgg4EOY4Nxes4Wd+s/HI7T0ui0An8zNNKqesbpOeluAU98A9+MQ/wC8
dmF0FOIna5eYOFelHMuPjsbEdsboTG4Tt1j9a/mnSB4Vq73D1leq+Ldzs6Qtsw1S
xvEaDCl3szeOqXST3jvUSLuHy4ZUJ6UTZmYFv1MTcuItAjOz9qjpgFWPTdXUioH4
aOCunC+15Bx2Mw16eouedOkvJ2QCEy9pPYToH1uB3Yr+vMsN2170llWSQ0Kg/KTm
7qCgCWIIiw5c9md9iXGY7N5drd00HZVFCdbr7FAv3CQTLfwBSSf2jQtjo01eDxj0
0oWs+IVYjLWog0VGvPr2UUh/3fVL32YcQp7lpGtXFwriW/KCw/OItVE/9NidOdSZ
lYPJQhFlxFSGEE3fukRaW3/2ldz2B/OT80gglZuCw42y1EOM4+TUwflKBnpijAwE
cZ89rIZ9cFuKjMHQBUwAtEiWGZ+qDeRpnWMJvimdqRBu+CTEB6IwL8BurA+WZ5q8
DuNzfjhScGqddrpHoLEVVRRc0qLsaybeoCRAOhIF3VnNNFKwk1CP/NY/B7ORmNOQ
xG91Zea0Eaq6Mr8bKeXe58sLIt1EyYkbSbmaLidABlqxRurZ9grVy/sEra6KqJPT
qXrbMhkSRAkKPqH9gzD1Oeddf8hntQVUaFYohQA4Iwv7+IksYzifp3VfU0DpWn+5
WrKTvD1lfVkfVm03/eTgbQUwufOB8Zx9iptAjuA9MFfumLlkf5IMgrya+QiIePYQ
QiA2fSg+Xlq7f6n2p2oAyX6T6EVIOPcMgpDVFyGLEmW6buo8mQQWori5ImvVKz2p
3npxYlQuHyWr7MyFJwe5qZx+eKbrtpQw3xUm9SQSCqmMWMVk5F9jhnYZxIBsN8xO
bKvDlnvzDN7CpB3xBQB1dt1lf211jJm7Y8AARwNLE8ZJItz4AQtRMG6Zr0XM+Xhx
Q1K+NKLvkZ6j4d452IfpGdWywt5OVC77XrDwbAAlM4z/OfIeEU6AvS6+DgGlOdme
GlU48/96wOKUtoEnfr8lKuJ1JrI4JmGlSwF4NJZoSkPvcuNeAJpAe3BmBokiaIgG
3PWFagSJcRex6yraGkA7eAwS6KJCJg/K+hh5Yc2XKOT7TjiP1+CkYxXmyT73lGas
N0nWOYzq6Zz6nzAw5C697Wd9VnNAaU4Fo0T+PiWda7c/KlDt+mgcp/MSMHfVIPFV
bDesdnHHnnHbzRNPdi1GIiPfQKMEVCEmVcDLnqIfvmNMejqB1FlImJc0CsBF18xx
KkmzvF1R5FY/1F3XOqejcWOc/V9cge/BQylUupzwgG4gHas/yaIV5hNkDxejilJi
VP2RlDotGYRvFibARZUosBjBjk16w4R8qSFS/jhxhXNbCgRoyLCyoU2x0glb9keo
krMeH3OgMsPigdMyZ3vaed92btUIVlbAN924/aOFNecGonJ5luj26E7589e7spwg
zq61dg7RimFx87o7L+xWoJqW47QM0Pmkb2PIm5P2dDx561NTRk1Atti0kVAWagMI
gToaNjXQKV6E1Vp1NshucQwe/nreuU7Z/JJef3WmfvHGs5orEgdK13HDXTvTrCcQ
FJYG4GRJ6Oj5ifHGduSU5EskhtB2xRziPokzHY5aV9X5gsKC541rOCdb7HrGuFEv
QOa4V+dQ3NBZ5Gw9e7dI8lavZvIcbyIDtpw5g12+segSKkQXXPCwDDMR1zwrnJ17
wJo68JCWIeT/QQFTIqUfOQGeJJtl/ssR2rVFiJCsMzLrzr4IleTcSC7QGdLpTW6J
AbsJnq7NvNloY6EKCi3JpgdexRT6DTldQ2hu0/96W7kIXs6tG2BEUT8XCfzwyoG8
r94v8IlLA4KeTSPVa0RYngwiYxUKz9IAIUBPEYpXNhubo1B60XynQYQESxXU7Zu0
ypYS1ZJczY67VtZx1Gi3JRv/fbOIxCnnIpAAjwJHp393HIOPD5tm/sBN3GfgVWVx
uNI4GQ4pM+fezjBJXuNP143OEUbKQIJJU4znofh4Xn+I0okPvsCfMnbv8t7fbsjG
cxf82X2rE2UTLsUfJwF4ZTkg50awZ9sVzNzt1dGv1QYBgGtwIq1oQmho8oFpWkPP
Xpl5JAyQuzn6pybsVPQZmtF5LKZq8PB2rI4rq2NjDAX+c2SSI3GHNubGkQHboMwg
vE8Mjs5ekGGXj0FF3KRQF0p4hGuclNwYJfQ1W3vzY7dJSwj92HNYNZUe9rdQB0LL
1BVakBXuMcrDvR2lvTl0N1axj1Hyj2QhOQqPTaRhFaMiSPLU/fvVgRXbyeBvf2zX
kofx91+bCi+6XyxSzMaipNwwJ4bpJQxUui+M71Y4/M33osVVhlgJ0NVXXqNUyJII
Y0Tvq3EGgb0hwIj1tg+fXvVVzyELgmk01eZn0Gus2fLsNZdks2y+RjYvTVdX8uVC
2AKNDcHphfUR6+CVhPpDfX2ng+8HKuR9ToqdyrwhIbMaryugwIrQHQ1QF+Qp2Ry0
Bg0JImdKMejk/wXEJmsLux/MZaz4fcWMgcbYECJrpH01CLrGxLxalyQl8kMTqgh5
lu7bNy8kmGSvvA9tL4PGjhGAbTKaUJOYGlO/Wzq0cmUCQ6g1C4nC5Qwg8emcRWkh
VxomyLWVtTB3JDUf+iRoTR4gpHL4Z30/poW3w3KIfgQoESwUs/48CP3qSElrzrG5
Y46t8xqwGHlHUAtZxu+CM5yfVq1nOh9CP0BUTX0Od90qZCZ96Rhcd9QRaqW/t+ys
3iq0oyAu6lZ9QxPGA7uNt8Pqp7eCjRrhgPomMJz1i1jYGQFZ6OKHqdD57O3c3OH8
iT1KI5ynqlnUAgYN7QeQH1zY8thRa8dFYRIPC+yefeCNG11MNjIQPD/4Z7zSYq+L
h9bxCVhw1S8ccn0aNb6rBbLsHzPjkUkfs5M3tszvNEKbz/yDucp0w5W0cNM20q8P
lXwxbTJk+2AYlLU2G6YKErHyKp08KpZVM/QZZKbrrIcL3McHtglamBU5mHBTEbtA
hX1drYWdlLhH4v7b7+zJ/ue470DO2h/dyeCwG1HtWQqVc1hMq80KxhKTpaMtBgc4
Bzc0FfNMAQ6AFvsgOwWQzKlaNMkBuI/ghPUZyQCDYMqxAn+ItnR0N3qDLqEwNkp4
rxwXQQwFX+KMaCe9mY6TCFrSlE7RAPd0jnKw4XlwVND0pJMI+x1UHHMgAvGaTU9q
xilZJkr9XXU04n0SFDO1+5b5bKDKoxlMVx6iZeLgc/TYx9qc6EY3VnGqadyta8SM
Z26lViKQtdbo3QbtaLK0+QXgjiHOdwcFN3FjmybyB4jCg1v7mi/X3hHFSqKvy2Ug
RqV9xbzDFH1fzXX0yElJsdjgMwurJ5392YxYiBOvorPfWyMMCTQ1t7a44xgcRoSX
KIcXHVNN0B5ktrb9XH7eoJgnnEmQ4Z0xTKXFSTKEROkHSZB7XdJpUurLP50lAzRv
6h2yKsuCp3xfP6dtNupsRnIAt8VDtYwBP2kikEybk7xxRqDigYro9YcuSdLSZTZG
gf4/E2h8do4Hnw8k5kyXQ66Ju7GmgvCfKB5RDgOe0JcTMa8Wd5bD8WmPUfPeJdZM
WG2OWHvw1feTbyRPJfWj+cWxm9rsf4odtVIrlbMRys9GwdUKCsASeJIS7/qPPbE4
DeluQIDR307fji6H8aUzQnEh1y60LJ9MyYEnX+q3sETtDZVvOZmAC5FA5GPDV9IT
yzP7OWercJ2Quqb5KR4CJf2S2yQum7j8VvM2mhI9aG2ZEbHYi/yID++yOftN6Yxx
q/gedZA+hYnNxGZlI21IjQyTEv2mUvYQoHmX7hUsjMaXtzrR49+XgvYFv8VVvTqT
O+NKrHxpuZgdcvLFjmWePb8ARr5ute4UILRIP7YM/7GC43jutdwSz8w0DwF1fEEh
iEAXQlQKQkKQoKnKGJ+/wwvT42enUzLQ0oWYaqaipZp7UVSwep+Cx7rPNHIyNukY
D0kVDUa4GATP9Vt4ctn3QAkGR6Hg99FOpzwwDqc9bVyH2APp5p5IzqUz4ZcK111B
Ctjx0ta3hc4UH93GxsGHj6qmDt6GYgMPqZrzCtyp2BhdnyMDFODfBiK6A3GA5XVS
4GmeL4DNvqWM7O5iS2KCt7dA+XRJiiKNLsy5/Z6LGZ3IsClFiL07D5NP0JL5Z2Sv
B25IAZ/zIjxcAqbUc71lEj2JfS3l2jVGDVs9J3BkkwdH3MDTKw40+JBX1WYHqe/E
rkjG7CTBAxX6D7ntn9PXAoRZ69vwmYVQH7IgepSll1pNFLZXY/IWm9jUMTwfZUD1
/ysR4t3mIlsRHrlGzPwzt60L1kJe5j8jQfadH+tTrxltGTZDm8QbozDhUTCyFQ8T
FcQ2g7Nxggb6qZOLTYW+01z047yTyQ1qYB+sY4QknquF+1RUvmYI0jG87UGumzE0
AnzljCXvAI8EzvUDTehQhErt9TfSk5psb9pif+QAp2kSCXMuxsUQJjdAO9mEB2KW
Nv6C9ckbTnOVZ5Fv/Szzic/aoUD7ZPq8+oDiljR7lPH5TW0GCZ/TyaIISGLCU6dn
tCzq6VzzPXZ6C/K6Fefv4lAHhUzdsn1skq4m8F+S4t6cU4RuMdFFUR1ZCe+IXZan
cLCbH0vzEf5YWnFQfsMiTVVoKr2ZX9gqnsKo43qAK5kUwSRwQQW/Y8+zctx1MpNg
H3ndDlTgfLGNkN6K8Ojod8X9qU/u2VTqjFypYvD902vu3tTUj9dpu6hR2xtUyBPx
4CexCKs8mbf4YiJVGIWHuJUWiauhT2WuVD0dyH07sAWwASpIG8yrmm3NwCeC1xkk
I0iX8R4OBQ9W+bCS5A9LKLraSXpjoQVgnTBorIUCkNWJpMWfnMoPOyWBuF4Z5UIF
QhpAY3DFAtmcvnDal0ZvCaiqZj7CeqDVX69+3j+FVd4578ZdF2+MR/VVtBelLPnB
czYQeAwIr2TIfDT8kBtt1vMW+0EHa65EjBYZY+Y11AJ7Vg7lya4QESw7vFUFP98I
ubwxPmmTqK3Ohr5cuMEmv4RWExC0Jbtq42jRC9xqwoX98LSFE+oqd2/t2My4duc6
CEyeRXRzjaDYFFIjpdh6Qs9H7DWW/wLf/uD2nuTVAHXhHY9iSapkNMbkSa+Iy0rh
7nbTa7g6GUyl4PrCgPI61aUzd5H2UD4wA8TrPZ5G+s+1vXnnduvwP1FSMWEQOQnL
/DuG8HzqS/x0skua3LfekLvVx6qyX8pFIBA2HJZuRL2pzvHBMVBCyUJOlvB9/QjY
J4Dz4R/iR7GvomYHQzBgpEhpKX9txTn/r+h5hrjv8ebbaVuZUOctLcllR1nA4xMm
mZ579+K42K82SDuhVvVthQBXsxafK9MiLbMrJhPDHl40UOOs7cD2EP8yZZXKUgiN
OgJPlAW/aGycgidQKpmMM2HtK0sdUpahz5uFYmYqFNyG4h7L3THUxxxF9HM02rgT
90LOYEGrMkloVrr9W8zs8iYc9j4sFG9b0yCQyTwLrMFJKNRX1XnppJ6biMSV7XBY
i8G6vQzCJ+n0XJuCxy8PMATBqLNu4cke1OPR9o+ErfXB9xk+DZeWjkLCFBXKuT6g
0Ykm/iQ7xzlWOKlSlE2giweuQ0QYH1moeGTNCWu0dGFLWkrkfm2Jm35EQm2yB+8k
APbuVwcOuZnUpNtuZgeNYcvCjrcIRaHRwkR3o47UX1BE1KPqzXU8Gbm2Fjw3QceT
pTp2AL+zgEbwTK5IMwHOucV1ie0ZtYHuNfeMAJiN+HvRaf0hIFSqQ7DiVu5z7FIY
C7lWi5ursyYD6LxTMu7zFAATzaB9AwnjxEPA3zePdAlZGb2BbHZuU3w9MAwMABbb
/kpy71Gucwo4xDAWWliFmABpVUy/VKB1yqjSTg5/sX7omxtjZhi6Kd8siFt25v1d
TebKXV5nkTQ4/hcPPDxSSyq3pDxxyyDaR1heeTIDzn6oDC4R9x3/e+Li81yedtoQ
3brQF27wR2nZq58kasq/fYv6zbS1M35pFNxHWCqcP6ZeBP16hrKUfJjQXTUq3vx8
aQbPojshyOOaa7G/vOZQfCzpMnD1lxJ8GTHrqMzfWov86bB70zjiU/8SOBd4fU4L
NqWTGmflOI9C75QgrRH2WCvWxF5uJFnXRkqaKqytSt3ZszjJoLj64CsW2x8diT0/
Ex08bO0JgCGWBbYYdfEfKhtYzCNKjbtLzifHfaxelhsAgjAXX81JQFBxPC2x+3UM
Wjn9X2OE5HzNAotysW3FeuKlIYf3MVjYoGMz3kD9QbZVCkrnzuWXsUXTDQsCzLZO
LbKdb6eNlWEN3cIce1WKm+l/bhu19CPLq/IrsMdLFY1rzRs8rJw95YAjoUiXCNuj
Te2oB5pBNoRz265Y4CQf/ZzY7SpQNvt0Un/gdLyUQddxdDbAQ2Nv4Wo1UtzaGQK0
0VyWuKVKpxr611Y8FoyakUq3ut5kEXwb479BmLiKKXIczU1r64kIj2uAmM2li4rB
t1Jv77OAGJihxKXar2rPte4xpZ5aNblIoV1q6gvDIbE4fF0/eVXh+k1Rw26mE5p0
c8xMuiTuuNwWQ4qaGB3jEG3Cfbo1zl2KQnJvTohUhvQjHF5UAVrpdlaw+IOq1Hl6
3VEHLekT0yYgDeSnh83n838iTdcYkPBOWB+9bqaoEGVnBQGVTiOPzFgUIb9nVcfO
j/m/v2lxgmxzjQMqZ7nx7rPGL7shKP6H3i5Ao0qTkLB3NUYppftsiF7/X+ArXVsY
0nj4mZGvU/BgcZvWUabBg9pMm/aaXQqmzVIaPpOy++s4aNBIqQmnJhQJgsF1Hqp+
WRnEL4c3vCf3fBT3RzCPT/X+el8TmeOvYcn+FUMmj9qHV9g6W9syQh7ocgJMW9Sf
bZV24KxqXo68lw7E2tBM8pcTyPCtfCkd2OecFN0G/aHl2AkPoOZSSrrUWBwbUhPr
WsuzB5ICw6FTO5E0G4rylLs7X/xM2y/jDkI8oSEeAZZB4COr0YgoddMYZiJb9NUh
nyTz65bAHeSe0/Dbr9xCgg1p8KRIYkPPt9UN/5o3EwSOF4A+dMiE5jyT5MQMjynF
kSFkA02jRTUQbJ5ifXxpmwL6VozpLjMKBvxvwtImYzJvIgJ4JJgxqKwb/reKEhh+
nvojUNbw4Q2aDyusdMVHmhgUSenacgQJ3tu50mWIC/mkCh5+ncbqpmLng/4rgTbc
Vba7KgVN7gIBggZyzRICA5bRINtR3N6cWpbNprsklQzWZcHnwmA3vUvJ0/9MwMpi
1rK4z44UiaDFFalltBD2JzGLpBCcnJVguUDgFZi1RYvWv/ghIC/1GCamroOkh+9D
oud1RCBndq54gJ0xokpeOshvPzWaqB+HccQMxNhBYH9nI+MoTkAKqkWxh0M6S9sx
Wbg/VBnBE1J+6rl/Z5tvwmcIa7IzsgjBg86EBJVq8wPAm9q5EUCjJd2w58SmpxdJ
xiNh+tvkpravn7p1MKrFO2o31YTwVdAUyLgxfTfVgNd7jczuPKVzyLApDzeYUlpK
kRnNQXz9hopilzoNKtcQiJl3ZTNE1J9ilKw4Q0h7WF7BCbZUoMu/DoIHdxIkr9ws
jHyViHCT/q7eKtNA5C53OOmua/TCt/D4BFuyq32NjGkvEmUrBaWtnaEUVDsiwrKL
gDfg435qBYg38NrHz0hrVmSjy5huwakAa8CfPe+xVZhRZMhXQbZYcfoT+pu23sh9
QFhQyNNynCRkQg50//jn3LFgZ3YV11SDLZzPX1p2L4AQpivtYyFLHZgg3M/e9iu2
h7ZID7SO7PcPXknnwRlDXYk34fjkXHhuRDOQfBlrJhM3KoDVf7CR9EIn4nozsU49
KgnqyuHoeOVfaLtdBkXfdeOg8h2Ebuvn4jAV2N5QvFTH2pf5iL8bPn3uR83lzIOC
LrTnrqUNoguuUDAC5NW7GbO/5VLBhvjJMixnPBA5oLcXpdhEm/eLF3g5AmfXgdCa
Po2Iz6z3GAAhgYUyqVJpOJKDzd+rFGSfh/Eqal70lLfWnUryztgnrQ/qR2SXcL6v
Y3q3DCzSscC5HqMv74WVUSisubprpV9eVWogvqMR6a7CppoWaO/Z69Hf9FElsX5l
GQuOeV2exLP2W+w3KEypY19p6A4tdwguYvewD8kKk2eZExpT1teVi7iYmDc8Kwca
BSdeRwz2Td2t+CXy9bA33bEuiexvMuamAG6ZwcY+dqj1Urj6apoSF6jWYeeVG3hS
Qj8ab4DOz65sO71Cq9R26RfswkhOZsXTOunSLmgHSDXjwzwEQZNnCz7nWyCvTKBe
EYccpo4ffF8yGKktVAO3tJNqt4nKJ/KGWgvpU/Vi8F7QFpmIYl/1j4R6pGzZcxlg
9uMXkrrfkvLw4XW54QovUkgy4V3FpTQ/Se4404rKUz1IQrRbuuzXSzZeKX6pyVOG
zhV3k6Z9i23/i6Juz7GhHydOS/tpEUdCC6tCzAhN/ewLeUlySqzDP1YlNZc8UU34
yjEFQTg2nitcgkCuz1KCJ4pezD50ocLZXSIBnyLQmp6yVJfwzbyWRl97OeTSaw8V
yP4hPy/kvHQMFZJ4a0WA0xxsM+N8PGKqNjiR1ZUfreneDzlwf30eUA3OFA5JbyWo
oCE/1i8RRXOI5+G44iRjY6Sx5kxg+T/LWCtzVlyjXpPFt6WXEytHLrFwX85bOsws
O/57PAYY9kQLbz3cnngHs4MQFHkHo+kJ9Y4yCQdfDVxWRhXXCs5WHtVit5ggTiQf
soVJ3oEnvrJ1jYctLYKweSxp6otDmGnIR35YRCNRrE4yiwSAe3gMqRGIiCzgAhP+
QvKwMTlIrhmXX92rw2/3xUwSJw9oWC3jd5V54NQrE8gMHhYq40K025JOKJRPg2xz
ZjKn603+nRFg1J2YW/mg1j5tlRZdkgw9//H8lPW4P8oi9ZuoTBe1IYbttmRTTxIh
ZRTgzrlCzeywQgGEdCM+9NVly+BmODjoP9X/Xxi/BBmxCXbb+/0RrpzoerPQmSEf
Ou4QVDjfy0KbZ4qJSKnAlbpCBRTuSOH+/MsmIi5kMGV8TT+DZ9p5sD0PjXSdtZvc
yHoYwnhlZGEzyIidsGjKEPF2oE6XtevQsvaytt8kFmpfVyBCvYZaBc9wNg5tccBG
59iNb2su4yEiu4rsK2cDHTSDbf2ubK+Xjv6COczk0OEgTXGxepSZaUC6VL3e7t/r
5a3CGMwyq0X69u5ku6dzblPwCjQKWHx5pq+Ai8YQnMhz+i+PNpMHfSh3UkRW/N0H
rOSYFKyrPCxQR9WSieelhudQSaYCN2zgVjYoh9tvrgS/QwrYzqEgr0noIeecFIUK
TgpT6qIeBkfKxOK89eM2V3DIegB8+GcNd4HJn2XmkLykD6w7TLtTmU/xJaSRcTZd
hYNSl5olwTaUQhLAMBTYMJ0MM3j2C3BF09fgpHVm3t4SY55NovrwV1HkT2D9FcKQ
08X90m//N1poxvZosHujjwcEUQlrYPe4hWdidwgepQTENsxhzNIQFdPBmx63qPCv
WykKdd4KCiCndTPyPq2DfgrNwpv6D+pk9lT7nQS5h3rXP0YwLdl99hfIMxFTfd5y
TcmnBsmapgOXLECLBJ/YRLG3OjM3DBfwc1TQ7I8A/CZVqq3JkMSdfXhH8/hulVzX
miYrj1dqfCBUbJ4F2+GkI7qkveB8T8ANCXKqWVJd1QzMDR9lKND4UWvdSwZjVdeF
ptQG/DcRwf760bKgG0DslkQrckBmdEOCGoa7DDU+bUlKeCMAs1pCjWarhNKcPW8h
apRPKvFnG/y2z0ooLWQXGmflvZpdnD2toRCWC5huJrPtAz9x6YjF3gZYliDphRqK
2VSMjjSsCNlVh7nriVkNikGldqOgWreqsVtFH2fOYrvrocARuJiieY0KBOPsxnqa
qFuHGb2wtOspRUbHCajhacS9VYaot0Lne5q1PTokAbFTfapwB+vUYrF46ZkymFta
H3YHMsYhXNoyPdCqYH88d8FxaxUZ1Tr/B+8Xksu2ZKm0dWrYJHf1L02Xo/IMog+W
VAbT6MnwVVUP4jwzy77O5ynsdojJ815x1C1oprr8Z9q3nUqn64DplXkZzgmixHRm
N96YxR+rlFMdWND1ro0Pob+t8DaFqfN27RptE26d2zhLl9HVNlWx/mnhPqXOiPkX
tNA9Wh81Dch0ZAXsNZilnItHqrqAGpK3JcO6Tfc+xNjHaOopWs8Q4oz3z02hF6m0
akY3SHtLpz+8CZW9IqUGVu7X6myhzsCedrpd7mfxIodlCsE66+rSWf5anjm5c/rA
kLz/Sb4YbPd+XnfAZg03H88jlJSYzmk4A10y6Fs9MhEZ0lldBUWIpt+xQVYEliDh
1Y2zQg/uztvwvO/rq2p1bWR49l2QzHWeJg2/AGfuN+IUv1u6NrvFujo5dzl+xs4a
cMkqNW5kI9+3Ns6XGvgF/qEG8l6OTfWEbEWErAczcjlCNPAf83Hb9dg5BzxlbYdT
2ICeeG0pzYXNiAd0d5hhaqqM8B4al3i3yY0MIQkrbRh/SoyRuUtMRolZzXCyXUtX
Q5D+/SDpk4th5XiL+5EWlzlcZOstLZ2CuoHJPRN74+s1SS0POMjcMQ5S8PVi3HVc
v+n3L1Hza2EYotolMHhRZmA6T8nZ8JhL9Oln1E/E6JWLrih+qJIxiXe992UQUEBf
0sKb3Kljowdydoacrw3L4A9MGd4s387uEfnoQpfUVhgTd+LsvFD5CRVkb6+Gw06z
WsBJsRPk97/lPfEteEKl29NMf0qHEqikSrZfTDfUEGwh48pbOr2Tb2C8+wN9ansM
ZKATM7Rh343l0Y4dDjydDhyW5qOmJZmAe7iG5RW/rH2lB6fSzQe3WL5r9F4QBPaj
u7qEU+5qRV/8PDN1NDEHEs8lNHv6Wkl9W0b5JZYn3XfGffA9OrSsgqLwXq/cGuvb
W5FkeZzoj3kZEfpFZOtpMrhiC0WQZ8o5mkhbCmIRrTbc0Hfd55XGXDC6tqhC9hjP
Ip+Fmcct5DRgRIQmaDWlEidCxO0INkJMrxNiHp2Sl7oskdyXtJQISmvRSzRfzS0z
kM4v+PvglA1tXmBQ9IUlvnIP3LQ7cjifotVmB72DIWHoW5O0OYT67k6tFh55rL9u
EJ6IBSt11hrq4kbeFRgYcC1ayO+fdG1mhqcaAoBOS5agIR1AmKw2xEtzq1udNvPR
wj3Hmrao0Eu0mYkqxBavtsJgFxaCMTZnla0yhibPK8kZs1WE/cl8DIBMn+wmiR9c
bP8+CNywY97nXvjuBPWhfRp91HLJt8AKhkMAtkyzVjb91FUD/uzbRH6uYyHW2Mly
snIhw3hv1xja7qaWhBXxsgXPvNOC76fzPzBUK8KMdVgfb6t4EBK/9xXTkULvASaT
tKPS1BKqI7NUYmTe73gWKdQ1JLTuky0Q7ZvUSI3jMVnC9C+ol0M4zlxHWPSyi7Sh
4xiQB48+ypQ8a46d4N0EwLl6BphE95dgjM1xoWC36L33LUj/YsGm+GTvh0QaOPwG
WJRY3RV6ORc2wgUrR1wdcLbI76jYFBYaauYPQWFwNJ3RHUW0aqxNNCdnNM8Qdxc6
UFJDcUQO7GMJJUZGOJZ9De3DBXTYBhnVX4IUaRNkW4BT9T8MTpbjttBxr5c05Ddj
xTs1lXjL/pBN5ONdt6hp000/tmtU4bjSxzjzZ3frwFcw0Y4Y6v2ZNVyPRzFQC1Q6
uAf+tHgZWoF68TCE4HbIrs10D3dRJ/JhTE9pFZ5KKoBMcTxHso1uQu0Ht/pKlbBZ
fbzjxazJ2t5VXHvMTjNstnWmTr8B9koGqFcwQPnwbZVeynhLD436lRfDNN2sjEeQ
iMHJv4/QjHjebVifopLGSNQ92gNC8Xur0yuSp+gUP4hRMUeM2G7OpdyqHViVhdkv
lwrwYeDEgEYvzz7K6f46oQWouKk/1k71nUbAH649v4LuNp5h3p/AFXeLbDqlk5qY
CAT8Jr+R0cQ8QurGRGqKn5OOqKBxAQThyJKnobNyvRG3SPyfRSN3O3RbV2qjUFRT
YaLlq1cSHrSm1C+RTxvnPABjuLD+LgZ4VHmxHOgwbNVip4V+gLzJ5dbL1ImXzz3w
DUCNeEF/hIfU7MEqwv8EnTfg8jXvo5jUjzHTb7wHtCG+roBxuC8M6f41O9/Ptwxt
jmjJLo64jn8J7BQMQbO1A0GUz7ku2vFDvghnO2aS37Qt5AWvKjQM18Ol27Q2s7tJ
wdmXDvswdYDVw9zNMUQd9vBvs7hR3oyGjdpjmrGxtU5Fdxzm+OLdGy13U1Ja3skP
GmI7yw3x7ouUJICj3Gwc6uFg3rIPBjhix6nKaYT71SKvBMm1WcBPkC0NeXiDxHOT
sPJmlr6A4AvOF0kd0ibm7cyH0wI0VhUCf3hp9xrCX7V9/FL1C6Mw/ydAtLGdgLlF
VDR3/qV5e0HhAl5Zrny9D3/UCn75rO5GS5ZlBcs4Ngp/SjEs8Npuw/oSQZfvep+s
iHxjRY7zGVhWmDn6AbgMQKVBHpKPzUUYx4Y6rzBN9rV1vNzBxjCDfAxhEzgFqphG
rMRF34uuiWQ7jnq01D2EaKvVALRQbgJOWnwmMv6rgcoDvFIJ7Toq36vhGYouDgU4
1f0ZL5vx6zAHaGfqha9/QC+v0l8xESVc8XDIC3O0OeXalSHlSD0urSrpDL2vx+/f
sO/I6iXjdwviRoNsK3nZwB5kEVjIE6qb59ascEO3y5SXyQFRBOmJ5zGzb6zGxbDx
fTTThL5qcSlail/rkq6VFr6SN8h/tapnLBjObP8ALBewQ/kmXz337HdsubIE+kxf
SxVJBjI7YwRrQ4bT3fVRB1X1R+PSujsGmHfXDj/lAcxgUURhzN3IZFZK+ud3wBfO
yao5US7S51yEf/gLPD4rEgAcC1Tg/RCw7DhhOp6M42K69mAvumWNgY5kmV0GCcFw
Gs7TNSOyeS5E+IC+HBgUX1YeFdSpOm6bSFZRJHnTs1+itKwOMJKMKZ+BUuuLeslG
iGbgihCGu+m/ZPaRDlPkN+1CakWkfAZ7V6424+mts9ozPAft5mJEQc/FQlUuyw+9
Wljl1aQ/mzdc0O8cyiaGeO8CC6neMKiyZzN4kPm4Mkn9vm4tec7WjLp8oFG38Qro
WXpe+EwLrVaaSEEDWr8C+kfDlikNvNBa+zOPQxTG7UeEkYy0iJlgw+tzqOD/14ax
LiEU6cFfs7GKV+3FOQBLJq561YaIO1cZwH4N8SUwUT6QpF6jRCeD2LGOEJPl8C4c
dnDUzprQbyeXb4vR4bbpYC++rQnyKrLZfIAaL/qfTp+MjnklaIetzZKboda3L5h4
TRkGqpXCEbsbDfBh8HeYM52rk25i7jx/7gb+KBAvB7gMNfDiQlxorVvLiUOByCYK
TgALLpSauoQGdOBMuTiWNUyv4yaxq1P5BBXMy8AU22io3BhEo++Kf5RJOKGaquTL
hXwHlxvcLTRVdqhZjthnjK31M0zlAU6zw/qp+pquUEM7Xs9FkBe4hlGnQDnNKVTA
5nmpv7X2ZTc3tYSBLJfR4EPEeyBxvNQVQ7b7NWDOyx0rIL+tSeDGOrqO8SW1CbOK
LwLn3hBbPwHq/AhMUrYaXOYhgTEFwmGQqSdJL46KV2NTRTF8qFlw1nTD0AGaYlmx
aXodaTGXwgt/piEotWoesuTqNH8SueIEM/9sIGa4aaFx2K415SeBsTMsRvaM12m0
SulRiVEfG9+3SqaO8pfvHg9Yg6CzSd7Bz8cKIzA5uNy3LgF7soieX9wAoGwbd+hN
sMqwv2+6XPzloNcDAG/8bx6xDN6ANP2xY79zBfSPmsegvYmjvDheA0DghIUiCVwU
RVizHtRdwJqbx93dfZbdN6UoqHRHtdpVeEuj+5VrJcYl7asP3WBiBsCLpzeCInlB
MqceKg9hPV6IBlNnsy3QjGAYFKXey4McnrYEwWJUsWx8XgK+9k5d6MVJviM3awdN
BxdUjAJLp4XFfNRq90mkstm0fjyfdN2Wt/Zt7YdgZ5iDo9nV1t34JWrNj/c5s3S3
YfeB6y1oD8v6c1THW2EaLQvUqHQsBGJxKJIxmg0B4Qs8LpHO90QUTldRfmW5gkia
m7E9/4qaVxGB0ajqdsci6KrjCxkNv0KgXrSSFxXX/x5VbEVTsq+pNsXYyaI0B+wh
Gt065GmAJwh4nSM4EVxbTu1VFOvyova9PXrBAaNVDxh8cfz13x43+CmyM3DRaH7U
FFuw/9AkkQV71qJOCLAkgFbMzljwMzQV5E6N1LK5FgaWahBTslFCMXNoB3ZA2mbZ
cvJwG3vW5XvqnzV5EtqyaH/gBU8i5vHJXA4uPDOZh3o4yWesbwcClIfEEk5cS0XC
2kr6hGUAhqeLuGpyzFNMknwkJkmQtBQsvigHp3Rpkj5bz1bCMk+eBgFrF0VItox2
B5CVtEUZkKwCobhyHG1U1Eo2nvs3DUTtrXxasV6+DjMY/TiPbfSqpahLiVLSAgmQ
klPQ1PXtB9H1HvOYaqgFKynGJ+yPwIGRmE26kd47Dx+cP87lhI2mZXyCiaucltR2
8S5ATMGowXpI3g6W3vHwSSez7UlTWRoS+VcLd3hwUOvvekDg1cRHWuDxIYAjcvSY
dps/PYWqsVXlXslm5XUpHaE+GgE/pqlqsuPNXF36rJU4Zn1h+DzC+DquTrMpcI62
lhKUhTuick6pFLvMHlabbvfQ5HnTAMS01gtjOkVAPJQ1GbJhc773qn0IT8rW81LP
qp2K9zvwiWcGKaMWi9fntYSegYv6CkLV8CPadhDNElWh/QZTp5EUS1z+bQTuWUCr
tIF3hoHU5YL/thYoSzJnzE8GStSGcQ30piTLg6nJ63ns/OfrTgpT1FUNDmQaVyPy
4/Z6ssXKHUA9TQRL4ClTykziSUqtwP5/Z3ggVc53FfUV7ouzUF3/0/K/UkZXcNkb
1WECpYV76ZSK3I7zVzUTZFIf+ySElGnsQ3O2YSfzqbVtZGJuF4yGEDtSVkOVBMBj
LoNY4TjKbQ63goyOr4nG/d4PxnWsiioivGmoWFcfyeI0+cwMgVvFrkjY5LNXEEPc
9mdL5nk9YTy79se5Ksf9D/NmXSEggx2VsQWwbXxyzsKOHZuSYECievZb0WreSi7v
al2XFpOffRMCfuoYDE9nYfa/yQMNb+0QnKGuJWTf5klD2VyJMfZZWsWnDmTDe3TY
5/nhv05EYN+aQ47JpOAkfllflLWddC/A+Uot9/xCco7AjrnW18/bdNTzWoNkxciA
RB8PUopD9GZjcMUn9wul3iQlMZ0s0l7vHjyObYMqtcfiSPRlH9U4PEuGJnf6R5vR
b4YGdI2sb6SmX2J7Vb/79ETdmDIWtF7Qa7u8WTfMKdI/U+D2Ypigc9Qx4KdH1LT1
oyLLVaWNhrY7BJOrccsBiQn0J4zyxg3BAUD+pm09rN2G0g+YPz3cxy/N35luU2y+
/CY+2rXKjmxS6TM2K7FAuusomUf/ebMq9bfUUGMA5gzg1afl2CqRKGqHyN/6q5qm
h4PvIFS/TY8kxJ+URTkcwabEuZaFSgGUthwHjna/Hnte6zcDRaC13UpwfZCmmE0z
n8r6n22dpXw0emhwtoXuB/CVpO16cHkXdVMhlm1QZYWinR1+QwI/q8Qm7xAfBas9
9Bs8S4BuWYlbksWNMd7PLE9RW69/JTWppFeUUUt2eDEDHzpMx0nX08BYm2eOY+RC
+bMi2Uyf+v/4FQ/j0N5kprTaVkw6WUnRDcizvSyfm27mmDVkyRN9hWiTmG46C4Bc
QJ/phw7Nlm7l6D7geo7GRBqNvk7yTFogmTQBjBG+sf2wIZppd68N2ECmtiKQ4jjY
gNU/JmJD2CRE3aLdFBJ5nnJLnhATBCXn5rgejEZaKADd6/kgBrOhNFm5kWMqS6Qz
UUlo+A6l5q1tk89s/U0w3MGaxta3LHmXdaOi4jPE6ZQafv7gmwIoUaBvvGfPXV7H
sRKiRC+BKdHqSjJOriuYzGftQ5gbSDkEIWjrgrhAFW9xYLBpTFAAIJLZWJoKFufK
zPanvlyG2OZ9GcFtgV7mMdwizx864JNhmGKjk441Vt+4JCE2sRywF335LlV3UcE/
ntTZAVJqkWtpb1tSY5Al9fMl76EV/JV+a4Lag3bZMmBerDD4hF3DdwHs3dZcEtPC
4htJfQmQbqDF+EuDF21+mBjIkcq8Zn5db+tWK+LqSKQc/vUIeMQx8nK47VF+U2VN
xH7yvxzOpohI//ARtudw0cC4ZLGhiyn2AEmVB5XZH/eQW1ylU+zv2Ski2rP/yhIh
BoyycCXmX3JD2w0q6mXTF2sg/IkmacGGVUMEbDCHI9C1NS8DHOimd72xVC+0i1ju
sj45I2CCQ49cRXEzf9ARLVcHycMOUmMsANsP2+Nr2H+BIweQR32PzwNSf/9R7Qim
eUE5dKZyi7ZmZo+TqjUXKSA2rg2iPAp5+o1czA5OyGsk1bdey4POr5xHkAra5GlD
gMBwcRBdkwevctLA0emMxotWlrTAt8e8MkDmB573T//MmOUC6+4OMn5sOgEOUsBj
6ZFOntFzHDBYe/Ue2TFRuvrVrixwhweaxevsPmY/SCbivV4KuF8h8cfnTDdDFrgw
BbtooZBvbzQ2zvzOsOvgyqR5WhPa7LG1nTPgsP1F5DBc8JJZRcjabeNCT1HcBlOa
toKQSG5e8LJngDCwUqZdbmMiiad18Tsh4GX8g+PySoLDokHQKZbQZadNeLbfoW1h
ouJWqo8KcMFF63nADiOie2DEAC1E2OzN/G+Z8W6dqBmAHNVDiw2vt7zAk8nVTLZb
tZ401mOemeik20yI130MwaS887bPVv1hdIKXuM95fMflpwf88K2L0Te25Fb08vhb
YCGD9JPWmf1n12aOjnE1M83G49nyTi+QMM9lu4mILWr8k60iYf0swqJU4VSjkFlu
NFai9RF0SWhkrsidS90s0Xck7Uc6WsJpt/gy2WBm31Ww76y8/WSnbFjRvcFZ6ovV
mvHMW8Xmj+dmsyX6sglarNayvZ6bL2wLhsUEvvrqU5tTQNAjBBiVG0RK3WfO5gHI
ICSk19CHy/AYgQ0pkMhc+dS/PR3Nb2Xm0fuAAvugg+QfmUuMIFhoCYWiAYa56rp+
t3SiFLmu7yP0dph6IzKxUNTiGPTXH+R7dRpJL/QqrfeOefCxxmCQvVMJOesaoaac
6zb7lAzozGhDtKTrzEr1yY0sWuhXGlWhZbvaAtZRpbtAk6u4Tclx9X3L1xro4D4Q
Z3RfMwR53ZYdwhbLL4i7Hzym5tgeb008gtIahgTDzmV7rq8k4nyMwv1YQhSQtBfG
JtjUQh7GAjdS3UtyCSg5QjsOCUWYMekezdNsdlUnX9Eeo/AKwg2J42I5EX8K1SBd
ppYeC5rltybpUQxr+wkcXR5Dr6ia8ouhLZvJ19bTlA02B8+q9ife6dy3ehEV7dcD
duauEEnUdXa6fJgaEt6n1HDFYemK2s525KVVnMIQVCe9pVNt83nEgLhfppRslK4x
pq/+YRX+pSskJ/CWdjGanHNoue6mvfatv0najxmPU0YQsM7AR6qs3MenDwqT0ePq
rVwdPxTVXZZW3qUphGEHJUBOcrXxqbmUPF+6x8YtqZ5pcGpE0lKYyzWSTMLkzYYq
tSkr7LpD7wPWD7oA5Nj/2oJ5mHKohupHbmZA4ofiWNWQA5NnNMMy5B5PksPVM3u2
fjBx98qjHbSTXSuRD1/8A3RHTUIolReo/a5Ii/PeLhXpfc1atv5KFqEU+pBQRs/1
ef/yYjldOIKoH0wk4u97lrUwYqaTLrpsNkPFPN3Csq4y2JnCFGM9FBCzuUAbFU2M
JvmywEohD7LogeeuL7LptphhcxxGaC0yjg/GNA64m3sOGVY9dszJkeN8qf1QY9lN
TuWBIVKKd0lVs+U2yaO4r5VZadhSsYVXQEP2vM3N9ZoUK/2Fv6tL7J6UzqgMcdUa
LB6L4kgkaqFZUdCd57Zk4nIgA1tWsHB2SypabcVlIfIFl1Xilg1WIrgGt00NvIKG
4oln1eCkX9s+5oYPYmDu4EInRfMoStQNFgZ43FnoHOlTNyvfPUUhxba9fQ39ij/t
k6uINSr1+dsQOhAypUY64Q+KojYzB3vEcvwb4yhEmSFcQ31yDOD1RL/Mb/hILW0i
LJnkBidpKhxGy+Qcn7eTudk5G05vrVDdL9U4f1sgt3Jq4G1gd+iJY8rqKvguxJns
swpw/RVma5A5Oc9/NrpjEEmYq2BYMoKedM7IcGcmHhQqQ/FwkJBuXVVwrv3/wSVn
kdR4dbPoEI+jLKp25h6IRX4HUtBptxAaGDs4L7RGiIgnIAXR9oB0unmxEfS7MAsS
5dtfqbJJ2NjrtZEDDEpgqHIl12/CYDYD918wDlJixxYqyRlflDivCouM7PQAvs2T
QwHC9WCRmtPAkX8AQn8ZrwF/Oa0vjEgvbzS91TC1SeGo5EDEHhUdIRb1BZCjs/Oc
zbouFyuG7g/mlXlk4rqab3cuN4YCAAVoUCB3pEmOChZqaPuNI6ZrI1ZeZFjHQDzC
wFpZtlXbKKVPSt4isJIsVMFpd6Iu8nxjb5LUX3escZrzSi29mJaycSTqEf5nKuLj
KnbcYGm5DsjF4OCyypjIL146f+qspiLQOG04D5VNJNUnKKa1GigTy9lvSkjGtGkK
ysawj7b4+rw0RHbS6pBIX8oDL+3vTLbpS3ne2UyGiAjz668cWTxzqirE7ethzF8I
P3J8mWmbAPLdHDCFq3C6cJQ+lN3zFoElydvY90HxSr1HS4+Wn9RTeAV2qaqJ8Y30
tw2uopDNiQOrUZXWdGSpEs4XPGJQZMS+oYAR9VRjXBlPo7JAwRQXpWi7QDnzEIww
ADvReamS2pGpuHscRdbn5VlzQl5FIxU57jOMoNNyGFyPT3gTALCNgwfLtbm7Kqid
h/QGMHsnDWbOAdWtIOQVi3glaafM20EyYq/nNdBxsgcRZJmENFHdayZh6bg41x+w
WXiZ/C4aWmseVKVZEGfflvKHlOVk+URXlPPIAiMybuxu6WGC8F5pc6vX1qZv6ww/
+kYsEbOCWKQWhOVe87WY1ugh2+KlFUO/gY89XNlfAa/xKbidyTl3UNBdQLLqOyjN
WtDsHVsnrP19vZ3cks3GwcNWg2e5GWMxxdGAeq8lK3NW/dq7vN9DnENfVc3mkUz+
HNKaYMJ9vbUPs0pLSfi5u2UTCHI3S0PLd3STErD4k5SVRugS0lM96aVeSFtcRUqp
2SesgmKvuZhtWtB7q5V/73WLkVvLPpe+mnAIcgZbzZBRWdI0hnTTRNpVbyftZBIR
Np0qfslflX/vnmMy/eHhm691UQ1+ZRfz2eGb2ug0Ke3w2xiE4pSf3EKlJdDvDobw
kkZnyHHTLRoGbLvNXcW9WnqB/A4ncCTltxHFFN9D29iqRxy+0UszVsRRha4rfDXk
7cdPyGunLw+pxVWEmK4qvPLaqwqkVSM3f7S6aXPSUqfqqZQIgqINXcUCYZ+6j6QN
Fm9Q0KBdF5dEqq6gpNf47RirXHo1rKCFUtcXbUAeEVrWMyPMSM3tb/xZeBoLesl/
gbZdOVxKuVTHw0n2wode65t5ppUAq6Nbuj3TtwgyRqPHdfz2qAWQ+AR9T+r/HoR9
Daqz+whP7NQAmk4kocO7saUIY9cvSUyQDSgGRkoy8tUm5aC5QiCUNMemw+7pmJLu
f1QQxqE3/SPBfba//dofJOIt48I2M8Vv075xLQYzNPWS+peQ6px9w9jfLyvgiJFh
gqIPp8k1zB9fts5g7MeWa9aeNXT7DZiYRrSguMCmi/s1dG6eqLqiaV48giQ+kujH
YwUe3GuyMGoFZpogvlwUmpnvHsM61IlsZXKFtFKfuJpyQH0/ra54TTuFlqyjZ1Hz
WPn4vkGox1h+7gWqsyWG1NuYOpEQGmEKH8tGzqiY1VY4CJ2bemCTw36nE+gtTKBw
L+03JifjDxq4N1MPIj7B8XACXAKwtTSuDBI7q4TYx8gOD49iOtw6mFi+GiuUK5oc
OGDCjrrxH4vu7iF7/YKZCarKxHDiB9K9xZLq7avr+dmXfh4ECm8B0RshhxeRtvHD
ObjTtfcvpZ6ZeD5J84BU9/W3nek9GyicOuKZw0QECzxq4Nz+aaH0eRgKKc0FfwSF
YAMOMaDdv6BdyojLWWcIC8kIMNEcBiGyR+p0Bpo5/bSIz69rJ+CtLpx/iPEYvJKW
/Xcg9VoZh9S9/shjZVGwqKx3EZWe4ui676C50YWrxVm/OwzTgFa/oynAOh0yqJH4
2PAXcRkWEPkzpG4bQuTqv8eA3vnGshVcs1nhEn+OHQvE+xRuEm4wpueGe8pufydJ
7PAG2y9lgCsUCyLMdjqBQPVSg2Pg/JTb7K0KctBfkLipY0OPKknDInh9MgXMwyHg
mAZhGVOKnN9D60ahfzx0IDh1Osy3koVYxw3wHQCRBeF46RyQRJA36kcXWshWj95u
WhIdHU5IQ5sA5nE9SECdlEAiUCUuTkTN2kLyeD9n/5DSAbUpXEmgXeLPPXu8k9sH
FQZkAQCWoEdO0e3dk3U9v1UcvAv4/bbCCqSVz/+QrFHF4vWmkX3PVg4BbA4TVh3y
HafH6OVS4WkvlJ7EbZu5KWfKKLQJp/TjFrwTHV26FnpiRxAMBWlHVOtyVf//U104
XI+JrKYizdRP2miITCoLAskyhjtp+ZXftRBFlkNZe1oDMdzi9Xzq/lKT0SiL2sJB
tX47eEJkY6JxXpGhnphp7BbQ4GmrXP6dpvxAE22LHHpvt8siYwukei8uxASjNbe+
iq6eux9EfjqK4UWzwoqJ6a3i+0F2XDYWCqd9Q2+N8VOKAKbNRpxLzIZSAN4AsY5+
kwRhNZ1SmkQNELJWk8jWOfvdPZgiX9b7NH/Eo9wPA6Df8yc0CeaBJOZ7i+bmRPLs
sRf9D/EX8mCijLmA2ZF9ZlTQlR2/x/Bk7sifXB/1lgBc0hu0aY+6M1lTSo4TAKWV
kyELSBn1OB4a6TegRBt/5IRB7X2dE/a+/DGHoCA35ggrCuMTNvMbhvTsZj7kDdxG
CGMLULD3rII7G/x8o6IPh9NhK80PFh2EuQF4BaTM3DurbiIKvCMIW6BJYyDJwAFE
i+F8TEUUxyut4jgDSk9AtIZWWG/G42vbJxzFLtXL1irH1Q1EefMO8GBWqyKaFXNt
rvPSYE7VnbX6NkEB1TqP/jvdKUEuQ+2B0qDqKNW7s9/dxWRrEbAWbfNF56m7Au02
ufEpj7LQo7Prdz0MDNaKZmg49T/DJ70N1+AgWttfJE0CwL8p9Cl4wHEK6yvXX4tL
WCpobXnMdX3r/GeDivzTGMLd3jyEX224cPRhsNYybWJavCmFKB0K4hF/rPQMqkrL
Ohy9y2FTpAXzY70biVq1ULz+GsoWBWD8ReSkN57ieUtS7R6ZuDn4dP8X4FJliNw4
+F10yZe0ypUH3Db6O6hxEpaGmqpmmmiBtcFQtgNFXvz3cKWkCx8B8i8d2qA+y5eZ
JcgNXrB8mRFZPS0zGei5ukrv+8H4DO4lXDnm96nOd9hMKilqbP9ENZ8B87uboerd
dBDdthBXl39TXeTXnlOBKGhCznvM6y/71rN/2jTYiL5/Nt6MuSeqzwW7Zj2EKRqA
qjaACrlxxOoApLU8GDlwSHSfRdasV8ma5dBXhaHnOUckrbReLxcOZSQDcJ5OM8/0
OoOSsDBxvn7qaS3wJIaqGqwLgj0sw1bz2Z1iHnOX8PnUB59PJF4Za7E47ulBKp4S
Ec4Zp7vGFMyVwD9+VrpkvOwq2Fiu274FJuP5yUCEi1iLS/NdZKELvR4CwHufwLpY
wjJiArprbY/chvpaHaF1RMGs36tp7s+U3iAKfmvc9e171nRs32eAGpsfq46Bnqpl
kLISbMiA+nxZYBdpaBnHZtZaAqnC7s+4JNTN+V0d42ll2smkDqmMdCBo0INWOyG4
5YbA7dGfrO3Nr0enRBS6vDD2oo/kzVMVqSr3ftg8GgqqR8kpm55AX6yEaQhdCk+e
AgNTi4g2+pyOGUqOwVUgXObR3bdKZJF2RqV0X3T+KkT9+AbZY/2pGQBbKq0fbVDH
nZVNzFHHqosa7TzKwjOw5zi7Fvjyneom9zjJx6HHUrCJfvD+6m2ldLWVcIf8uWt0
ziFU7zSpbRFta2hKa+INt9e71WMdQCj/+qtfa4LxFja+qxTtfsDzCWNbkTPo5uDI
MrOQa3Dh+pDtrLZsPhME/XvMByyqreVoSYs0/r7WX4dvuwdf+K1ilaStrwHFY8L3
fLGrmIcRaoWoi6Z77WlNfrDAo92nE/co4H2EblYsDp6XCcgBNQfVB2Fg9WSwBN1O
i8jZybov9yX80teJXHt9rIPCzXa77xJ8CjfMammsLqkgHpQSfCm+ztilqRwUsL1k
zUyNsCosciP4WaAf4xHh6vhynGRQkyI2c8hbF+cT3s6Th2dCLklwwjnrLekAhaV9
koLuVW1si3fchkH/gQXzOTbgZFDsg3PxeJptEy7ADoTeHRsCwAXBXbHrKk6rOWur
c1ycYCRlDI4lendZg7HfT9T0BbmR2wPntZJhM/XYpNkIIMgG0zxMWdfX5/l22mla
ex/7pCopaJBDtTDDIvN4f4N6fzEAyAuBo1wrXbY9hM85up0ZlzVnWW/D33ZkHM5/
yz0Z8lvWr8BLTznMEm2B0tBz1SVz7Y2gRkcOI7Sa/7PJ6kqOBJTHv1qz0fiGl/ni
bqTy+Dcu0BhtyEyVo/9ZK4ZlX+YqZHbZuy+ZDWrIfFNe6r7s2EyafZE4vdSfQ4fc
G4zjlRk1ez9ihNhwRowpFebAKjEON1TfpgburhHgNtOIEj3bDJt8CxWg42L4HvEV
c4og78O1urz0h3z8KghBU703TtIhD9NK4yJ6kXUTlZGbC05hkcjpDvRXq0BMOcmO
ip7lS5PZXdiLDicmSBOzPLo1O3MrtUJfHTrWNbTp32K2po5HtAeHQnRcnFBOQOZ0
mg/+3eqEnfz088quwxPOFTHygOG2JUYsspnmMPojjk+HTA2xhFFuCef1pWTDf34C
HfwrLs03R+kVhwKdUQcIt5g2V4eIK5m2P3HFh9deuwSP5TqLcnrvnjLgW2fe0j7W
lIemmqhdyTKHbvTvxOMJ513NbE7GpNV2yQFeJbiLqA1nE9QO9m4dHuOGRamsvyIG
+MGrIaf+yS9M0F1NQwuMwOUbZzWQfEmHtTDfvaAddjdmTcDFY3+hVggsgRaRHgER
2WaS2Z0IkD5Sm5wCESR6YAIn2gj/erKOZIxp3kHxFcEH1A68e8cLhYxM8Rs4wADy
7ceP0gNuf1Zk52PpLrc9hBNKHQiUI9x2JI1RqiiKZ2L1zK6TibHTrCdwS5s9JUr+
SLfOuh2ny6XfbLg3pv/dKfRUT1b9QNuZ0Y9UXW1oBtLZy5kOtsGHrALtJvKizMan
dno0oSuILatcxBYrkcC1ltWfsijqjAbb59CA7cE9a4BqI7bcgEYSl9b0nbIgNthX
JJ9xkfWZ4w0GP1wyTh4QUcNCXGOckRzoNZNdOn8lfAAe2vgjBE/hpPukyV22HwZW
d+rc/t7uj1ovm/ry9K3zaXznApEljpxO5w1BJS2s7BRTizlA4NcMeBUvYVQvLWL0
GAE1qJCThOF2oZi0pBEGMzIrTxFhPVpQ9lsdPAyrKaGxI2zpEIXcvPWNVWX8cSKF
hqOYRnL98+J0TsdXIu9/IUvjLPkOzemitVzgmAegdJ3VUQKsz4inMXPw2gseQYTD
Da6BEnJN9Iqgb26vVRnDjonbj2DxHyEqjUYSn0EVQJbur6l5P9M4jtlkRICUnHGt
YNinipwpBP9mwGzHwwx3hWf5+YMzHceImUno5JAZvBggBZhDEaWRKni2HWZkbuhU
03nSVFepvzxJC+utm2SBoCe/D9OLMCEmIp6pMJvOa9SFl6CyZiu/0j2OLOvhMH5r
qJFVoEZ3GmHQaLzxxoZhuQ1EEJ+WUcsUqIylLVhGFk904C7IZNhlOaSz2a3nvaLI
3e7IC42Te6pcf+f9rD1AWgKVqi5ec7M2fagb872WIeUl5LTuVn3o8ch8Rv9zD8QW
MnXTLVuLbK/vZQHUNpCqRaJ+LJJF0vsvWPvCzBewtTEEivoKLJLd59wfVshZ5iCy
nlt21iBd0NTMlJEe7TynS+/BhdVvkhtTwwGt5hRx2w+RQsjQ+dzmB+rR6p45LyLy
VUC091v+D74PRSKyS5ZuDAHrmjqi55n3L+fExLKPi0CoLNrfE4JITuLxTDMAbK6C
HeH0H8tayqNN5RM2S84NSY8oEP4xuiXu0aGPIqv5bhoWebj4UQYL+1lF9Aq9FO4f
mHc1ZdkUvvVzKaWyMXPrzICfRVT8y3E13TA5DrB+68aOYVNb2VJ8H/PBZGoEsV9z
KQRXX2lgZL1LHephfww2AiY2ou7qN2wwH2gCqxX/r3U2s1+CIshyrkUY7wV6+Yoi
Ah1h/FB7hcm3h9fcOldMo6ygzXeGR11JjvNGn7jktQ9yrcIyzgkac0PinJpfMkNP
FlFd9abpE9dQvLa/lN81q9Hk9I1fg/TC3BMPdgmERjYYg12udwTULkr/nuEv66qi
CGgHSke71w0x8o73rSJGKnDqOdlAvtyWWA3kIBGGQrS9txmxw0pzoK1kdnfjoc/m
v4ZOqVriZLuOLCSLBocKkfD8eqYsH3GY0N5PSg8ldGIteP401BhNHKJ1cLPGAwpo
QtujDM8HwjzKp4uMpgMnmSGLYOTIzFWDownzoOOcjHZh88RF7x2g5iXpjfmVu/XT
KnGbNG8v0eg9zfV5SW37idLDYRkJpSKvcvP2fuZ964Ff34kE0D82Gs0EK5lVlp2N
YImKFckkV037dkIOp5yfmR3j1KzhNvPTlBAPpQ5ae477WrYS6z1Sir4ejtq9e6zh
RlWVTVXehRC3STG/qq2uGaml6KApO5dwlfzEpBZDiZIhjqGKiDrPRR6qFp/q//70
3YtXb0PpSQt3Eju3WALQZ3KEnvXrfNVsLbep1+hGoHwv5UJ/M1w12D85z3qs2KBo
CQ1AFcFgaAaUtNlPgYYjIFpwKGRCmvpuaDRs89Z/4jOtq/Xu9fNaCQWRdSO3A3NH
xaGFvX1v8O7dAKBnKSeLNLLiSdL0OdsfNKLCr9tfcXWD6oGNT0BD+LhYjGneunJ1
77P3AEEsq0W5HKRzDh66ZSxuSr5kbHec4K5ZS4VKKGkSiGvzPtyv4YdGm8+oh9P1
2JM04VlIZ9FtXRdq9neVT6eK/FtaDQ5tH15p9ry9EbJYlGd1suPteg8+NZIf0CCt
8kHN/U8orNfMJoJE7iRybDQZh6jWXCMZPQRCWQYHVEJLRgTczzoOZuk8L9vuftSH
7GgLiBl7nentL0peNYmgrVCrn2jooj6c8jMCHmXC7x+h9sipoU4/p1kP0CRMnngY
Cp1NvcxTL2g2pRsw1dIBfcp4lr5isIysWL45DPLhP5+459giVEkoMinSwGBMC5n0
o9p52++oUamrM4vHSdU8dQQ+vQL2qPDwzQedP/tZ8/ie8YcR5N3SVkl5X4sEgXOz
Xh3ckCrLX+OHhsiPbZ7xcxShBm1L2bw0YgSG/ykXyA2bUe1h9W2geninvF/oQklX
6X3A5ZjUVKx9mRJSR0jlowYBF7eLc3j7FTL2gZAU8K+8/sknr6QIc1ux0mJKybPt
+Qrm7J2UTrWSGP9iMF3a6DPo6TYs3lFEecLeyE7zUdAfeBcRSx80Na4SGrCzBswp
Ug5ejl74PVTceEh4PsEF9CoTHgNXvdxQBgywdrP1n0ccV5a1Axs+LEKzSWXREWF8
3dxX19U29vHWWEcR8xfpGymRPmtxh9IgH+7Kncfu5iV/wERzukiSWg7Bw7w+an00
u74G+MQh763mHDUKAhs4VL7+p3HE23djYsShoQ65P3VyCMyMaLTDiwHNyzis1M63
Rb1SBx1dmpTRPY8smYvTbL3iArFvD/ERpcvqxqeIepJVMw6JAhMEROEumjQDUlEU
E0hNhTWiA1tLHr3uhiHpZSaZbN1/Q5NNWeM0K97uN9+JX8jeLPTIZ2fqL47h+h3H
vua3ox4tmhzuziniYASiCj9m6u889pfSAagAnZMvuWNvTLO5WtWx0WBmIkycSoO9
dktV4EQB8G7L1irXjOXbBBpDGqI492f0YzthytvzZF5xAxgNjlNCOWtOLHBK9I4u
/MQv7XyYNX9ya5cHZwj+O49BcXPmKtHE+niCOY7Lt7pJ/w3HBVQO0cDZGFuxN6IJ
xtruUPNarxw6HHq8b52dsOG0GCaEnkSs/AuWZFPvSJwe+Gr3IO6iCFVZjzVmIpcm
pwLtTz+nIRRncn/gB+LJuDJvj+gjqza8IkfVcFNv5Ldy0Oi+3xRln5rHH0YWdFXJ
4iF4KIv8smhPYcjPrl8tEzZGLULILHZ5S1C37tDuAxh9Z30Ves1cX73TGL/shGwa
4fkcOyOgiy9yqV72lFfSV87fgWp8C+9lMJrehXd9S244myZo35ONDHEB7Bw4TCxd
bRuG8T3UL6QOfK7UBz6/y9rKPgd6vIfHV8M5fwS7vYniONGSN93ouqLu798Dr85U
QAJnBSA1ZjYn15J0bOt5FVnlCB6yACXF4QZ2ukHFxsYABgn2YnKIC8GoWxq2mqQ8
1GtUYvH+nrPZPihGkuo8Y+tSYV84JG26mHp2kXIK1KEW713eFJYyFQYoq8oa/35b
10KR4c/7R+0KGmzLY0fNJxDLwJXtU+S5NfI3nTxiLBdIxVmnU0MmVrccaRvpvrHU
3vMhx6LzoDUA+aXJopMoJ3ncVhUlO6xXw2bQ3FB7xHrWHH63dbyqsz07iYzdXdrA
T9iGM7lZe66BvtWUzJ8JVgXm6Qrb9or5dNbT4umyivjb++OCnNHxjhLl37cTKwtW
cMIRX/PhsUH4d/y2O+aMHa7OD0Y51jtX469vgn224hXUHB90qoK3ClMbbCSGIEhr
O42r0B6MlF7RcTGukBTp7pPj1Bdga/jNW5WLIN7E79RdZULtRBoqUQo35HQ2oO78
7Jz6Ai6vn2vRJXVS23cKI+eZUW4QV/kyvnG7SWN38I5pjP3L4cHaF9UDDlUE/2Yv
10f3JTz+fPT8uGPxZC5K5KOxM956kqWttHL0EfidEJfrYbWp1NlAtQ/vVKzuWH6G
Jvc7uYR9U4zGsRcQA/egDDPpkfPlMU1jNdliN4b5jI3rxL1lWTS7ltm+U6G1VHhX
5u0RJrLaN7bk702r2RzezTyuqCQhzXYMu9cas236tIhoB1ufD+2WHdbWNUDM+p7J
knnUhCvken4Ad0kGpaHF5QzRAcvwE/g0b5OkOPxGW7F30qG+NlbP6u5gbgwEYn/e
PmfKiwuK4kTecfpg+swdnw1av57tUgiEqBDq1T/1LtTQw7vtK6ErDxt8XaXhYq1z
jxcozPxVn2z+fJ3TbE/X89vdm1EK5olZ3PnWknDOVmO/Fn2h6H1gYbV1YCmPzasR
nQScFaRvg6wOxFpqDr6gtc5XLYmIVpOUFeYwImFYW4x9RBWz5FmEEQf5W5M+ptm8
BypQaX+xZDEekEpM/JyJLy9gkh/H1dwCrmuGTQ5JIHh32e70Sg0qNhnOiZtqPB72
b11w6PTOEUvGCoY46HMmfHTpyq1+6+cOMl89dq6rDuIrOMwYc3c7n1ELgCAhtCkX
Xe013em90dbSbHniM91aEYpx5smfpOyOAK6mofuagKx87PUQi8kTWEPAK59gP/MF
Juq7Tfcdp5PUEvKZafq1Fd//9naOGYo86wrfCuTJAT5gEl8F3GwVfXVwpbCo/yh9
tCWXewj8scDXXLfnpeCs/PLiza9zxVgosZb6i+3Bjri0iZp4oK4qg8iyfgRYI6E1
5WDIQIT4ndjhLGicq15JM9X4MnM613Lc7zP83kZ1R2ig8PJtmEiMJ0tSKRie4wYC
JWUDKekA1Z3jW5//fy8LUxKGxHLzw9TyeJUkTiS3yeIVZhGyNK1iSj1RuD1boKrI
J1IABBfRLbf8GBPEiS6n76sLpH1fKWvmFq++P6Od+hlVw7pCvJCPkhKYV4aLi4Bx
FzeOipbJVb/aDeL7qZ50WmOHtEZjABdj902CRBTpt/6d96UIdFDQmPJM4a/7saDi
B6NtFpAIP1BaesF6CyLCjxEUySrk2fw+vWU8REbeje4uaI5Y1JmHvvtaHECstdVf
lMfGnSlZTVem1kFN8D3geyvYICvFZvl8F4y9G3+Thbe8F6Lr49hUOD/QOEJvF+F+
XJMsWBQqoGXPnHq30ZyG4hBla7QHG4Z5BG19KLwL+ed/oAzgjTRFxHpIMLD5ZpOO
3ieZ+HNS2AmQGoU7wBIkPXP/ab+l3bJbss8HfsrxAi5iJDAKrRRDnUCKz7MFMpO0
89UkX22M3zhunjaoUDd/dRcZ0lo5q4qglhlZZmM7jAX6OaURSPBDoEFPmqTflQ60
sJEGbdGc2ToPm/LhgBRjsKh4jnHO7eKo0pUeqOxGb/txq/gbix+J42YDbXYgNa9i
s1W4YF5+jmM6W2ZdTdcqpfHF0FyyeZ3JVTFCxMeZPuwK4W2eDwe/cVEznodUOocn
sOo+wmBo4Lju9kN3Zz8mJUBt8LPsxSQLiJ5NLdyHSHGH3MEfC4Ynx9UEQTHO9Lh5
EWX0vQJn8AFtA6v55gRBahQriQlVEP/167agpgLcycpjYwQVMF5PVJgQHRnuA4dk
RlLBztQhrZQ6oSuDBGtNOZnOVYQIQinZaCcc+Tzrbd8Vu5GxG6aKZ7pxmiEyp67U
0oO9K9FKSzKUw4W0J6uu7P7HE16AE3CQl8041paKHlLN8OpRXvsCKPovsbPSF9ql
odnd26xCj6YEleM33v8LFw5kboXJMrj404JFA2lCn4fkNd9M+Y/u+9HQ+fiP9stb
loK9aAa8rhHbNruixLuzVOzRG2fozJGyMgT0Y3uNuImAsUv7nmcG3F8g4ki/rgOU
b80nq2cwPJahLal9HHZJPr8UdIx5Ay29OmZ+3VvqX/R6oufPBuM3EOVphRPPBUn9
XBQVdb64TqGjvmDjBlJqqTZ/jMB5WMxcLtN1r8sWHEvlY6bOB+66cB+1Sz8YdWlV
FKKiE03CiQNYP4vkhNCckNCgNIBscYPfh7+BcvdF7X93L2dqkJ4aWNNTWKRbkpPW
MLUuEj39zmfZAZPMxEgKI3phOqRyb7KArFXd6xEb8RcTZajnv1bPcB6y/pYBe6Hi
dpGcvj0weJOXusd4Rx0i/OdNjiObSks/NHzKIPlgyjXCeflbwZ1KJkZWuDWwcL8G
RUPtkpMViE97libXg7LNekAXbnyLvRv9lR1cebBmqd9LO7XIWegXpBN91RoPA0ag
1ThRORSPUHRTTLX1BpbJa67X0lHuhLyJOVQY+anWqJ4Ny437V+U1IapIFJdpgwiM
MG6Yb+aVbD5Y+DiXOPLTwXB0CzOC3fnWMxk73T4vtPm+qfoHFHG0L+VB3mDt6BVO
+QeIJyh8huTjp+y5zzOOYmdnrKWr7VAe6X28Zg2p7aYsZvqwpBl2S5wvAZD5E+hS
5ieONXcreKpkn7ah6QirNIgwcZSIO0IYFPAo0PlAyHzkid5fgJ45TUhOOap8osYV
kkqGtC8fTEIkVf6/r4IXIbmOHKoUZI9dNk0kN/xV5DdBqhi76KUjQR5m69stykaS
O80pW+hmMi1O2OlkcO4D/wyjLoWnppP92Zb5UlHTYiGAMaqqWJGVcxCTL4iEwpsW
PgLNGkX3FHVdJFNu7cMkeocoL/n8LJVBKY0m0qMJvtbrAwbU0p0+uH0UlhMVXXir
8bv330dcvYeNhF6OkN2kHOUOzivBQprZyA4xRt4V2i5ZRRa4hLujgk+GHPN5oVvy
YQuaQEDCtE9uTZxOQtL27BdxzwuFM2LYXb3oaYNfqpGPlqJRPitL3gKc6dfQEp0+
+hxFt8gPsENRcLNym8xP6qfU9xpJ3eAHZbFqUp6qIeqmODPtByVxDLQqpsyY57rc
ISKwAU09Ui3/YXZIeBUcenPVV0rQHLvZhhhxOWdcjxBjJ1QURcLuLzTiEOUXMry3
vMLxUXG9XmuQPGlmjwgLRLst0aeNW3BsA3MV0OjeLfsNXfJyTvdGEYNPBd1ESAKo
/OCwgyn1IuxxBDsx/D8f1Q/VttailE1g/OjVeUuK2SIuUphVi9xziWO0LszDWyUg
uFBn8frQUzzkNApp+HlpGWMaFXpFybEPxAGNghjBJZ5nXIMFwbdXk7mAYZUhA/hm
9BHpx9WquXrYQfbC+Pa2e8tYCu6xJu1gPCLee9h4/BebrOFtV+mhRkBlAe0Oj/TM
b86szdbdrJ18L8dqvIUd1tL1UiZd3t99UODdTq8jd3Lx4kc5tpU6zR5HyGr+qLuH
0kTBfj5VrPEksVO9lv4hmGdn/XVEaikZWHYQ9IeUdwIvzFVc/336NUCEtBSILyTZ
FWTVL6dktZC4zkYrmwJVoBUZ9xsbLtEaHs2PwZdp2CkC2KKFkJS4FDosZ1YCAhbH
ykRk2fGInQjUNnor90j4Iq//CUe/GP2bv3k+aTxQbVW+UBl/27sOirmNzzA2rWiM
h5GQrw5OF5t/e3uINyStEI1Opo4PwP6iVG0j5bUh0R2yTEE9Rsue2Ox+CxGyWgyW
PnbbyfcquT81cro0PVJ/YvIVoAJZHALdpSDzQl6VdHtOWz5G76dbDtwEF3KDun24
OUkR07WapErTyeHgwzwgbh27+d0R+HO2W56juqKxOqQc+YfGxM1/eyg/KLh7E4OQ
HdE2ZCHxF83Mwt3+aWAcpYqRlAiF4AHb7zkIPycHCJmvw1uS+Nl4X7I4moerzuQH
7/HrPB3cFtK/HmXTuejqTJdwkWiJViuQBnjQmVbs0vqaXO63bpoq2FGYgUGb1/JB
hzKUDMnqU6pgvKFLx+tspH6Q+srQPf8gbL2aSPxZIqDcJGrHm7Qz3yyUIclUUZuo
aty+bBUJIcnLSKKL8q3/SM51s5I2a+Y+1AyLoSltwFI7VDtx5QNMcus/Yv+4Fg+J
dkK107e5Gr+46YKY3kq1ohRjMl0+8WLVEUtae9J1oqtWH2FW0GDHc12rTNLIZMjp
s0c2lNuqXHy1xQFn+qZ1cCZTkeaJBeJ1V7b8QQZmNYcuI8Pk99w20ZIBXE9ZgEf6
hQ55NOJDH8rYYukhrZj71d0ueXRl16iuMIXguMZUZ+USC73ukNq4MI8Ts273LFkj
oVgemtOk5B09pyGNrFWfEjqghSi8SGAp34e+qzw98GfF5Tw9gqLuEDW4L+VNzICs
2oAXMXwTdqt4wZIY04PZKA/AxarU4hiZHIcCSb3b4c09aW+RL17q5a1Pr76k06Ly
iDMMDIv7zU4+jPniu6m4kkWfz6ocNNeBf2X/mb6zStkJHf3H7Z3X5tSiKTMsyeUb
+lWZ5mWem4hv/F5pgUP0D9xgldfhk1Hy+tV0YE2Fjk63QkLJq1CdsD2kWHWxj4Ji
dYiPNII9Sz1OAFK5a+vMcdl5WWqQszHGpchN23IuZvikBQkVuovmAsGDrckUZ2SR
I0wsXcCGF6Wtg1GwbXYVDxGTmW4MFnN4seiA1PI9VeUPKVs5vnvKISoDzEqdS7vK
ITKsYvGopIOngw+rVYv68nY+IRPw70moTJcHzbwaPscDaluLjmSWJi+sc6yTARNJ
+bupL1w6mG2nwhEqCAiuXNpTWRTavFtK+4UJmpNLVhJEJte2NKs6LOF5rB7CdFFD
HsYf1l3e2ghsAhsuArE7YlYxirTqk7hE0q7QjDUWJdTvgin5hVn59xaE46C/W5/L
uSGiSHHC5D2Mwboaws/7FrYYzlSDjF0H51ItROJgK3Nf9S8vGsOmeAFAm2kt1Uxt
iAE40X3lHezLHnjqKqznNy0iTYqP7R8QyTMmxgIqoCYANJm3Dm6O/2ErS750Madt
H1E6GKrVPFteTcVcJepxi1ndy5z5qWi7Wx0AF/KHnPNfnB7EEoj94qvCy/FRWQMe
3g/m2i5jH4x9Rrh/18HYbyDHmyKxbmRwEPPTdR6+fuz9meOJ8fPiO86nqaKpa2pN
0leoKy7ocBnrjC0GaN5sURoXQJ0RV7GTD8Cn1DzLcPB5rFYP462KfbluWP4h1+Z0
+zIMKWtRyBD7NQo7Zw/ao/l3fZSVHfL87PfpN+cHCV10KOES8EyeB9V0A8ZEvc7J
+u3Hs/KbBCOeEqE1hOu/M6R9QOYcgpBJ9BZ2f45j2TgQ+0SJuxProNwWKuCreIIX
fZhGe3azwbkyUDYv0OTqUXWn1T9VH37uPTtsTGn1Q7iyOumxt/UibLK8pvPwJzTS
DDiugqSPW1Yr/zAXPZb6KsPmKlYE6lJ2Ta3wUek2OaeqkUMVhtKLkJhbDgQrDvbw
V5DwZdpbAezJ4JQkJEAmzhlnqjSsh38918KASpIdLNJ4APWmRJTKq8J7IVNm5yfw
MzI5P6QE1v7n4D28FF6yrEW+apj8xY/vdcQthcD5p+Xi6IUjzYQ2Ezw59Nuudz0m
QRtUQI8OeYi1eS5m16k3/Ijw2aXgIYpMukVJ/s74tyGTq+Vctgk9GXfsDz/kW2Bc
I67kOImlCEuozU0zhVQe7U/UuaO1bEJrqcbZKVhGGxXBj4g7O/gr8p9qcNWYWVB9
WCWobye8zeGIIc7jGCzf+JeuTNB15oUlXoRcDKxc1L2Q/e0Y1VUd04srWrmLxzwU
+F0R6fHfRf1IXK45AHLK67S73p3HN9Xg0wSDVrqFF7YGDxlOdVKe2l657ApNnqKd
qXWdWW6oUDDI32OrPVi7knLhaJeCs12a/0p00kRyy6EvUqKY/F//80j5bVBqZOd1
YNj8C6MjgyGJ3+w+GsPv72Wid9WFHPta1yMCR99yOa3EgOU2vI9+Q+zc5GGE+0/M
CE46tvM8UGNci6vpGZ6+EkxuZPrU23rrvH/vfBbjsuMn0j4zDmQC0TnTBclIFfJG
WwNwmAgrBXSiFDajVlHN9vhakwKONy7Kr2KuPpKbw5JgX1+NwUloAwGceCW3eaFX
Klu+bBDvWKPC9VKJApBeWdnADoM/xscX0Qqr+N35WBLYaYjBL6mHXl1J+E46veB5
NNA+j+BeXsbN6whaGANFZiPiOoWSxSEcuVR/pALijcrPdQC6mXnQIPcB3W6uCSkF
u4OfKlGGO0aQJl4WD0rtQMZ40YPCZ906QIT1GZnHwd0/M7sHWw39fG6ONujXhPb5
RPmNfMZicgiXRZKH5reJqMvjxVmSJwHay3mlQxN07ZRm3k+E3Ivah4rGDYF281qK
IuBw2xGlwPFE1MFmWdK17qdhrIBQr1ebDLApv7zzfKmYQw3uQOGGk0VtEsMgtxdK
4V/LVfv7AzTO1kwRe02V0VmWImpcY0MgqkM6520c0Vb4wW6NYRuhPimCNleSKY/d
AgqN1YusPTQ+LDaLracHOS6IFJhP+6Yl50jWs0wWNaiEpK0utzyzpQ5yskDCb3eL
FRQvJ6yRm72FmniQixvKVJ3zpAMPMGhBDFovIRO34Ku7irKyenrhouVT1sim00RV
EH9kJ9mkK0RcqhKNTcG7Dl9itgP0pfL2FzSBQFkjeiUnnBG44JzOBqfmrttQDoDX
mtC76y7INB0BySTgtkC17CREn2/Yj5i0ivlBOPz/LDRQWM7qIAxnxHJxcxntEoxb
FCEPS3o68YdHK8diJ6XxgyhyX6PHUufqWG+89O0pZ4VJs6yc43+HcEVWzoLN1MzY
/EXNbLtemEb8tTdaa14+Us9m4+syYRG21G2Xu1zrnzsPWxJ3m98zpP0PjM/eKqX8
+suIpgKrZsaBwc9MSkSbil3j4F883yATUZ3XICU6m2FFguiHu/72drWcgS4GK7b2
3xMZpmnB5uNnf6c7Am9z88SK4G1BzEuQ2mKb0h/gE+s3/n6vmqZXGpSkZZ2e7kHG
ViuoWmEmlnj7LVpy5a8kHY1w+gyNcoh8p1+SWNwYtwTl3xhun8IYbAxyUSpc0D2O
WLbD/3X83qEZ8JICuclTUFrTqNCK3Siyluwkq6NKif2yaEGyk/oYyK4s1uPpPqAO
7lCFXpgHfrCYRgaYfHjJRrNA/Lz8FR/qOLm8/Rz44LMzQ0zogK16IuS480+8wZgu
+ZYcX5O6ej8TernQgH05Y53QJIXwveGqi4G6nkFpOHuu6bbQRBJBaUT5gPRcg4nW
r1qflieqVYeiFmU4tcRu1dfPmXsMBh96j2/kd1RbvFLNpOC2SF4mHzpEV5ZL+8u1
nnihF6EZ0N5WPpHQMwlkehnAi29rg4TYtlqq9+rX4MivsSBVpaMS10EY3NWMbQGY
7FJoLcVRhS7qLkAfaefB7fV+4Bhb6651+qRqR+rcOFQFXKoVNEjEt3G3tYb3T3MY
p4BcXWiI8aw3bMkt9Vr0WiWdTTvEWP+hnstlGgNfnVvh7WQlX1I5mfb18EalyWEZ
qUBZoXOIj0N+uRYvS1oQ4Tpj4IZoGSSjbTPjMGSnZ8tO3TbwoSqtl2K5I00gkXpc
0iBtTs6PO6hPUYs5/StxhyHYx4Fw3E7V8JXLk2kfZE0O6lsVgdbQOhhaw3gm1ehy
1gtFt88LlNzxIZtzjPXa+akMutBXD1yJf6CfwJlu+3aRgsoRrPX2uIG7A5yklIck
8IZkPyjwJjmpNWBH7S3/ywn5r5xRzx+4RkkNH+2aIPktzWeEM6l7bGP3BUIsP734
QHyO3IPcOOvmT+l0TYu86zn80MYx5FHXFVeaP1glyCNBiDP/8XJftOe/NGiXZqVM
T84CS/75dIJuI2eZcxaeKzamPnFsYyCchY14DKZFhe8CybI1XSstBgwNPxnrabt7
hHUjYJrTvgm+gUi2sJEpBxv3ovtKJBRQ7YInWsmIHCMZL2boPe4m0LW8xEZBvfMu
YedTcamqXPRPWF3Zy8UIX9fJ4yIt8NgbU5Anr+Lml1UzcTWujqFt7+soey7G3tH8
npJDPtNI2BZjUOTG0neWiFYkkqKJ22jZlniET81u+/CSnwiKDD8HDa7MpD/TGVNw
BY6txaNdYP+0nfSCOsHC3q7h+oznJL0LLVEd8qU20LccezT9jQUhfcz3ERkUEDt/
WaGVK0XgR2osW69htGJKbULDEi7sUMr+idPsIEJmK5dLBitMlGvLVy7NF5ibMBMj
dHWd7P/HWTYCEukTfaJbm8Qvp2IPjWwm2ui7yWTniLEWoo4yUYhepWMKeoV5WGsf
1H9TzFvZTh9uApTVlFXtBBDPZoa4eQUjXEe6b9mGLcdmuBBHnTU/uNFSmb1unbdK
Vkb4j1J2jq1H3RZNOuddQ7Q9t7W2Xb4/wmN+Sp6gULHi456aJwQZ6yqT4F553xEX
htgyitMFm71KPPUnLBqOzAsvok1ySBgGDhu9iuhNoyxeP8hYcpxGPAFL3jlzHc2h
0JEv7gMS2vJ5FRndylMgDvK2xYZnhtbUul7YR+DXhWfDvv22yJuVaYuZw/zZK6uj
m0TlQ9EFgk6XKGHALwpowZK/ZK9hkVZ+v4L4AQTvNWnnEjVJvTkcdzW0mRd0XBJ5
ByJDHFl4UtLtZ5NCjKYyw7HinrBKvWO3Px3LyOmpalpY6cefd9l8Cbr8s5eYze/o
bUWFM9FVq++mlLjHJH9fdndeNWcTGlWplDimnM23C0QiLDDd/Kxvg+LwX/bPnlc1
yoF4OgDk0s8dFmwjGx4ITWK8UDYGBB+dKR0CqwG8D3JAOXy/c2Mv0/Il96IhWOH6
eAR15HqWnPcQOs+nCKw/zSQvoEfAFfh/9KHl0RNdjUEgCOvo5rWd+VpM3RjVR7TV
4oLsfPZkCOna+/Zl6H4/piO6By8ZjvckOyZike1g0KR1yU2bc0abKc/hcq1Ti8/Z
qu5ieq/5P6+q3L/OjzgSgcgRpCb8rC61lm7Md9jLw7pwsEgfri6W4g61T37/ga5N
RN01OfVujMozr2uShMB1/MFC1atRIQLKO4q0Vd4in2T9pf7XcQu17z41lVytWwXc
2BlUEtA39NjDoBPHmTLK/Z5pncnvqYuRNzu8EvE+y9frqLBl//ZDf5ngoA8OrmQI
vLzQVoMlJHGIkHtyf69Qh1fGd3X8xDMLjPjnBL/Xisat5oGe6tnElOkG6QQdnShs
9IL1jWTjF5i7++gUgoqTOq1DLE5KKXvUG8jbc91kf/H4csotA0ELV4DBrSzw3sCy
f4AP77ikleRzvze8ZINSG7rMElvUOhsOskrJA6tvj/HVae7yF6W+xSbwznDMtGj6
Iev2BKhBM3ecOloa+3xNJUJgwXAn8IAqKrOtZOCiwuinqtRo8/uE8Viq04wEsnpw
3bPw8FroztixXQBKdl03HZgwMnIj1cscZHkIMeFXlx6dYqvUtooSeID1mPyr+8lK
n/VtZrmeJCS1o6tQCZ31URMpXb+PwNVFzUGFb0PZVEN/Isbd++ORCWnUMV6qqFUg
TlhOzuBd/S6jfZhVfgZKzqQg5DISSX17CvK82oH1R2VnELVTqQcW9u4nhEMKDdyJ
qq53H5yuDCe64vYUcCqkkljwshQgmvpLPobd5KboEgGpKhh8q4v4tKR3bO6Y2Hvi
c3ZZS1KpCDw9tzCLvUn793r9/DPD0NS9Eg52UYMvNEQDAkDZM62x289bZxwV/Nwq
1JVQh0dR/KuZPxnl5fTs8wZ8S9S0NABTTk3zKGp9X8gLhvobOUpL9a0BpYCiHfTv
fcqyBR3eoBut1+hWZHAU0pleDRnvf3E3TiIs73Y6o5sof7g/C6sibqK/RoxZQOrV
o9WlylphO1Zht6k5FoE3nTk2jwhmLHxmtSHU3+D0hIcWhLeUakV09CT2/hgAC1CL
GzcWcc7JZHjywJJcYvSvsDl+DAsiOrxPBpo7fQAtuyroHmvJl9dGoj4Mf6yK0DDG
C5Slgimkv4kxie90IRVPNvMyLWO+LYjbkCzPRXCA0WqIukriaHMn2fbfPf2CoU30
xeWxhO4+ltsFhOekH/tsg4mp0QjD3BrZEkWcOnWsKiJWtnFnt+4PKA0iBy8QS2VK
nTGrkKEKiwdc5/44jHpXug0FCdKYT6glsRRtVjrEehK1w08Q660OiO+1ZyoBt7CV
g5FJU+zNbeD8pNCkFwyj/AaGCffy3MGsfGNqbJke5AEON5/H1fjGg265pRvxD9as
UosMuSbNDVeo4t6cEiYJPKY+PHDH9wGY12lRIbvlzBwf6Jp96GRMS/B+X331lGHo
H2JpiPNRqqrcetN+RPVosjkA+BcfZEhZoyNb4I1x875SlMtnR2phFEs1X218UPtP
De7aKGMxVDoftmAOTsK3dqQwT9+hJx2IlKcpXTyehCcvHL2S/ipRhPoEtT5xme4h
hCCXoNlcCuKPUnmQ/sWgOKdvmWYS6Pc+NpLH27bAVF981ALD7gyIFB56MVHJcnH4
D8Sgd7N2ZidZa+4/g5hWLkWKD8KhPizVw1E8cnXix50k2mxUdf0tx/aKd4HxID74
eMTX1r19WTUF0Qw2ITloIiR2IsyhLe0OnVCeiGgyxl/wRgrWxhY3UZ7xCJA+Nqrf
bwhpkCQsy+Ys0n7sjaihOw9fL731VHZxF6b8dMKSwZxKgUZOJcI+3ORSzGYh8Qsb
e6IvrVv/HiREvv6OrCbcrd0yaLqdyNkHufC1sf+d/ZGYl/IVLmX1/HsB18h1T4l2
wwglBn8/ISmLZ6gbc+dHdQGF1DlRZzRYtlhhjlA6scH2yB0XTXBf0xxLjI5yr8ti
o5W9Bh4o2/68KFeAp+eprjoC0iEyLdIssqDHFT2eCcP8uqunBA5hlzy1vT/b9ibq
v0nbS4C8MbB6Env1r3cZl1PslkiKOdI+RUlNar05ZibrsDZ92Oa6Fup/LJ6Jo8Mf
rsHRbPaSgF4ZjLeZKk4WhsfNKD1jCTUV6xceKe58/UOPaRmcqaf0AspQKC1J0E7f
o+N7+9swKHmWbZPWHxIV4TdjzPdYy8Nqm428WLZh28pf4B0IXrzxFFhu52L8LWAL
87ncisPcCXFtcNEfW3ao5i/ia0wVt+IDIuffVLJ0ODM6a/f96f2my06vzywI7o+R
/AM+37IM0N3Mp7LIPEpJqApYAJaQ9v9hoycVlPeZdr8UZU1TM5FssHSYEa/QOlDY
HyDHteMYXc127t2nS/exfby+nKgQHT683qJ/kDiEQn5Ix5iYiJdxwYUE7YgqdhTq
gj27JA6gbG0WZ9PfgTWcfMM5Iu3ZlzwnO/qCtcJJ4/qGrelsMp6qFZZEc/yXIIIH
IN0zQ/IJ1dR6CxTdXwrk2VaWS/s9huHcwgGHvb1TLzgmEuvMCl5wM8f5+pJWcXbR
Jyl66D7UKu/B3vMDfoCgM8qD7e7zDB9znr2Ne0h4YwhXVN6McDFGYyXOBYo+M/OZ
rg2m1JB8Yvz2JHVrk+TdhViw0jtcINxNRXXuzkHjMeaj1ldmsAtP1gGisfyuzf8U
56eGUV2B7G0VrMJNtc5lL5yMyfy5vTqOeibGUwuybsi5a3PsWJBVXAcMxKlOI6xk
Q8oOWH5Sne/h0a0wXZ6fRaL+Us9NiKBDsoV6l8YROXb4NiVsJGgahddkRD7XHjVs
OcJGg5/9IBQ/9W6GzD0x+NL9ybSkhY21OORjU4yx+ym4nHt9nDi23hoBjziujJAE
QbdjpOO4HbIutUV3db+eRC/2C+ZbJsaWuo50pM8fqRiAHPfIXccq0GoKI2FAlVek
tJ7vWkcUEXszQkmYXzSbrxHvZps+lwuUY9maj0dGZClYINLgaLII1B+cOTl5y2jS
QdsdfUy30UyIkRYJcQsaiLT4umjr4n66PSC2UILSgOo=
`protect END_PROTECTED
