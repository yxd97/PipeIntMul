`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/qx1G/TqA3Y5hvK/COx9d9zyYlnQ0k+ZpDcCvW8HcMz2sQuKqiq/BPoqxyKlHhW
5uTAmcQZiHmXob7uyE4fC9bUYRPk6RgI46uwTv8jq30LE7Fq9CjKNQUFAWqP+Qyl
Y1Lrl69I4uuONbWI8ojIpxYRpadobXd57UklG60RUiIL8C6V+bHTrxo+6oEj3IoI
TOq6MJcRkF/DEmKnDqgKEfSJcSVDJ9yz4NuXm0ONqTe0xSfPKh703IuDq8ds5r+q
B7D/NI2HzUxHjTviVqcWyAVJdxAp4TO7NM2eCi4J+eA=
`protect END_PROTECTED
