`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u62TX/Z7KXHSPI9mXjuyyInIfqhq/g4FoeCS0ZpuwTvdXmhe28IXV4A6ju0kGsVC
qAD+Idbqp/a+VS+O5dm5mKj4whascKGeEOh0OrK1OUKYa9uyxNyP1RPk36BZxFNs
PtMP1FCM0wuBBW7/vGCjCUQqizFWCKRYG/VfwU9TYQlWaee2fPuspubnCHCHqZZf
E/nIfdcOFR8j0nF/fvoGnWjjCYL8Z8+enQXi9rBfIee4PiNgJlao5O+JpcadGb79
V0YBWMIW5LD0jxkqYF2wN63BQ9Rkt4NfiPH80OVpZCEFCyhV6NEAbPSD5yFDq7xN
VtAUGnDs8rG17612cONV51n9AFMMDpHzqd29krmHbA8a0gBiBZc5yFJ4pcyzPmLB
V72IrIOUI2gNd6VIr6MEvdemkdxgIut3M68zeiCWno7x+zkwnB4lJfW/F4p0pB0A
cuATL3Tv6AKOTWnNM8dNV7Ot5sWtz4YGIzAL2/ENvaAy78gLED9VCQp/3DlU+HQ6
e6qTRBEB+sEgChru43yW0Y8Ol97kz5tDTNfO/mWW+pS6jEucfMR9RbAAusoaVNHE
03DiajSzNiri/Ct4mtnXEuApV+Cvmpt1Km0++UbRYy6w6lFH5IyThsA2GavooKMu
PaMTjZLjIbKShRcSznoPt6ke9wjFPamtBrG+jEuXbYovFVI1+cDAUJRZIRKHXfHl
a0ycogTrzTVar/bKt6p77IdifeJMitDs3mntymf87OjEdrIDLARWUfsJBlUEGZqK
V7SRG5PlhKwFFRy3t5jhnUYWCCvtit710MX/19T1DuLEMMRvjlG0VfvrKi7q6XAq
jBY6OMzEo1GNfQigekxc4OPCBlR3i0Odk983Lqxa5/HtCGH4sSW48YL+55btg6xG
YXXRzNzRAiqNgcyy0yT6TzUykslA8jbOIsE1Q19lKD4RLOpsyaUiPoL0PKaehK5L
`protect END_PROTECTED
