`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TGt+78fuU9DvEhSQlqY5gVUJEQNMaqw+C1qSbpQvu9Ot9RJoORTKEFV4wVNq1nY+
IyN3VUTFjmuA3tvw6l4zsMzyxFUzwDj+4+ehbXOjgnNGILbiNc+uQhtPNkDk1gz5
tarHCZNoiAoAMMfz8kOXdlVVFKO/cXFqTNuU6L+67DGHizwYi5egTs2syqAO0bWN
FedCJfasfOl7aKj4IMUOnKfrrtcD8m419yggI+/6Y219Y4EGZe+ANx8eIfk27kWZ
VNu7efRcuJQrlKdcbrap1g+LA6/AWv44r77YCHqmke8GYz7SuInuofDuPp2IgzPE
ZY55mgYa1UGywNbdY4eCDVTlgvaQuq/DIW77BhFsJCJtVdlx2Ih6o9UD8SE4H9hk
bqz5HQH8H/PiWz052MQMMvtdwbg1zbqD63Hvt1SZUyMqrpEGa0VQKL8CocGn/ttx
J3Kvs6PR3YVg/yClldy3DJwMcD99/CVL92pUeSVAvmLjwTOE9OaYuJiXwJW3iNb5
AF09PnJD1WroweLtI8+pgPp0m43lAZHGnGusNDRUgpEFIZsKenV32mcrwUB4UXqL
2BnlSmGVlzhp0gQ+N2hVRxfru4mxlAcHsynkzev1XcYvOfM3HA5j2kq4cbsEDiW4
IcyDl+B30BbXrK3S/A4lCKSLlRqBl2Tswr2ERB6HRT0ANnw9dYBgiy3QJKiVD4z/
4Oa26pKtk4WEgBANrnvdR8LcKLAWS8w3uBY+CWV9g/Dzd+u7caXggCj+LYGyyn/M
Iv9zcKUX4xclPnWgX4n1qyvauZIDC0tUglcyQs9En1yg9OlJRumw1caBt5TVKUBe
HFcWz6OVlsBu23P5uQqVVVrH2huVmGfhp4j5i1tR248=
`protect END_PROTECTED
