`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fHeEPTEr3zx+WLSANESskVQqSmh0G2dxysykcuMOXTrIX9hVRa6rSjPH9lSajaq
UFIUgKDj1m0rQdfH9eURUpD+XbbUeEF+Sm7xGUkoOdTyqyxIy4DT3RQ5YcxRhWIb
zOddJOPuAEu+5l5T+1RouqQMqb8iy07QalxCC1JwUDsuAQEWjYqanIL3aOrBs5SX
eel7LaCzGVW455tFi8OSaBx5fsXUgkLWPQbThVy+44EEFuy3fXocg7QZ7ObDLrOg
ZkoXnoMypn1EZgbS/JS7O3/z4ziDPG5yj+AaWcTCJ6LPL92vdtqXfad+FvxLWww0
SuwBM1YMrjFht2c9VAPq45mc/3g1uohksQ3YIST3KbM/FvX+EvujKg2HIvvSoBMx
yCi4qotCQnXaBC9qKh8lw+8l6GAvszIo3MXzZ19eXI6iB9MJo8R2UYHXxnk9Ej8J
uniuwzOevpzN8VcdTQr7Mg4DTSPTxjBi7/2KCls33DM=
`protect END_PROTECTED
