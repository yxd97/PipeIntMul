`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2/v1k4qcLuUmDaLor0el0mcBerc0ABWhh7KECA4fZcAL9QdTVzhCB2d0hTs0MtX
JlbiAhHRgu3V71l1lfZpQEodlDat2peTi2t7/T2HqZq61JBN9jsAZdV9R0wQKjjr
V2C1MazOzhKEyVJspnHS8pF4v4V/wi8wScJNSISHgSJCby/fC06JVX02EdL0p8zA
iPpRtuhKUdUeChPd6JvtUM/GGXjufHX2rUCWd571ubTpmyb2CLmUdOvELlFYVfVb
AZ+GeWBTnTbnFSrdpDJ9u1FXSY1hgykVIBbDdzJYVej1zN8I1ijvrNk4jqXkQL/e
pQVZXOyHAcDjqRLUHSoYDknAnUilkOEDv1hVNg1v3uLUvN/9X2cMs60HONZ9/q5e
vcOHoHxPDh9lV766jcWXu+8Z3rL1F/0vlcmvVBsDfTx9HQmB+2Sfkv85ZKrsgr4f
`protect END_PROTECTED
