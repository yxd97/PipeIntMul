`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yzew2rVSN4sWazMj+BIkC3rcR1X7O+DiDvR5UXfiw27f1vqaxNVxuWWTiN8YtCLe
q06dbavZKqrhw6zRIDugWEUkJK1Lq5iHQunYKo0+AKJ7SERQWK4W7m6+0vzZDOGw
YLFinfw/Shx11G1Jam3u5xs2UO7H5cVgHf3ryQhFBdQYXkQl7QvT6SUrp/6lpgKb
WdQMIrVq98rN8IwH18yrqdvEljCWjHPxAEWry2IqvpIrJqySsRG4CJYC5VbsSeqC
hFT11wBct/pL1yXyl7ajrODXICORJxXL49zRg7A2cA6e6JU/TM6u+dQr27+gOZkR
Th4Vm/tWiCkXc8uhgEPJlWiyAl+VnFu0wqnemnQ4Wfn0c2yXbsFLvnSaCNQt6+cv
`protect END_PROTECTED
