`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NdTV/yQrdmSyUY2Gscirgj/5FlLFlSALIqwxiEs7nBB059VHMe+x+ARp/09g+Gk
mO8p4galyN0Hso3v8Jh2qO8fLujmear+axBUl7DvPebBZLlrJRlj+nsGepd2XD9b
wr5z7GkX2c2k2mfnBksDOFe/AHw4D4BP4Zc8MidmzeJ6N5hve7dEhGMZeyhays6h
7R00TWXJ7KJWR8rrXCOwzI1tc2jqgXMiG7gLLEQFVLIASsPihY9/cXP9bvzCWD7D
WTBghwiPjVVeaAzdRLSZsw1GCCHIclHkYHzqaIIK+HtgwzVuhzSAX3u6QAh+j5sP
c0NRLbVY+LHKbOz0pFGcHw==
`protect END_PROTECTED
