`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6sojFEPUEwk/jkJR6J0DwgKmVVQoEkiNjq9mXlrIoss8gkygwCiH2RtSoXF+Lyti
V/a3EotQ3moH44G/O0k+I6tFZSPf9SD48l6wMHZ2Z2fJQAt8Y6Un+A0cK1F4L5t0
v6Trw86D/YaqKh0JDHn4Ky5mNOmaGtYCZXWDCWsrFwdTBNKaThN39BKZwjgzUENQ
32Uc00oOCvckeRdQEH0idVXJz+kMB69p6A4SbYBg/+nXqOzJFGQQ3kcXnDlFX0Z7
`protect END_PROTECTED
