`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IlYNmnRuMkDUFWAzocUWET5lL2s3FQrIh1lBwiA2AjkCeHOHhFCl7TVZtQ8jKKtl
aHjHIyYQxpeUIXIgEYPNLg2y6/jx7LzeslArVQ09rIF16b9MqBJQs0GIi4F6CcT6
PiIlIvqJblIL2BV/7+3VRgsBHLpTs1NXFRkqwHO5Ae4nDnlvLBUUQpp0KlDddqHl
Od6uckmXUNIjlDfaOhY9DHCWBLt0cuVR+AxhLaiPEhk6ByWfBg0yoebbXW23drFq
Ry+8FA3wga0JKBMN1jswjEOWXmNysCadmyYRmN45jHtu7ORqxen+x0TejVp0d54U
TL/PBlewilBJP7sqIARQId79yws8S8S/sAECYOprnHNkrzQjdseVtPvuI9K3PCka
pZnX8tEkZm9lUEPcXpgnL8jdQ4+Y+NHkE/BPFfi8BHpUiEIHlU5+H/7JvYvnGXzX
zvrLRVS5eGgfuhzBKyoS0mlsByfqeCWs6kk4Swz/HgsDCtDZZJJHGpKMZ3R9GzzM
xslpF+HtY9BB2Kwm4pDPN5PxNw+Fhcd2L3GShSOzmP2wYaC3pZ8KTi10ltr693BG
Jj7ggMH35S5LM4gcFxgnIbk307RZ59+o9LUddpJuw0degh53DArNhlx96zXeShGy
LJgDz+O2IjUDpKvv3zPZlyYakUckg62ZmauxIlXCHFV930e1SswM96J68+TrGVQW
UkjXvb2lfRKYJC7N370XWgMFbW65wFotbMPcijbjQQgUG+RaVzdwG/3WUlBP15iy
`protect END_PROTECTED
