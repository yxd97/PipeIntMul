`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8FCMqb2r73FVwCJWv4tpkBubucxrbcfXnA/S0qjU4Isx75LzWqSI8sB70Vf7Szn
RNe7Mv+B1aVK3cp1drhrgIEpxQ3AB9NSrWm+zq7oEjn+L7thYQBQk1/NMv6r+odK
xeOm5mZl0ishLQWynVeeeasljh3osmPsLvVSiRF9sHa14tOHC202PQdUfYsqWCyN
aOa6TQgQv6MIDbnE0ikIL8BdItEltTc7FTt/jSzrk7HvDMcei33wl9JSwMR0VN3S
9KiZ5M6AzKufkkSqqKBPZ+ok9oZIYVTPSBeGwEJoVaHZmcG7u2FcfF0y1L5XoPW7
mS0gMSSbdmT5ahT/lgkkk1qE6LT+zzpmuaTRMy3O29OuMndOTYK+bYTbNufE7dv1
pW9IAPcI5F2LRr0WshJVrLQ2ijKCWMkinZaxYNY+qcgn0rsOqWgfG9W2KVa/SggD
5UWCjSMzJ3EOar5GyYTL+aPik75e/0uxF0SKx1T3aHVqpwJy3XQF2OtnvDYXXX+l
rLigJ3bcw/1jhfG7JkJBlA==
`protect END_PROTECTED
