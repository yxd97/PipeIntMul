`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qa0NhLEzDltCXRhQ+g3nzZElc7PqeS6SMpmqaE3FIyMfwIPohxhm3RP3j2o1IS5I
szQBoQB+9CZnGAQwpA36mOobo65/hd23Ic+XIq3RNgr+gdbLwIV0kKellc4XgWXn
StHBCpBtZ4PC1/DPMezqV0gqIydyqVwnWrf8wRfNRCfPf1BbznG3PH7i7NPmTS/e
vWY4rXRcS5Zw1jgAzgw8Tw66nRYJzO+UFGWvvjGe8P7zud4q1WNtCtTKaMr7OJ44
IBnIiwjfawxNKBc7BzsNq3ZE5/QixgQlewJ1XmDmpjxXyQfiRF0Fg8CJg09ZlNCR
6IssLhXdUNIjdfQv8W2uusJkjSQ28T+E2kk9DxCKgjZxz4/yqO4IsOuvB95Aqw6f
T/I6qgCoeqmQiYvXtxVDhRqKvVsl8mROjUGCmyGN4sOCExVafhPQrvcMd4h6VO39
uZc/jNfzJLmfLz71Tw2ngajf8hGKiWYDSBHWMpzjEkDKkKbjCB2V7tfOS5OwTGZZ
`protect END_PROTECTED
