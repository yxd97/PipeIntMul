`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBMVYCA6a65iiWuwMBKI8+Gt8kOubdCyBwvCHTX7hFvMBMyXQAKPbVw0aaV1z8YR
2zxb3+cy5x7d7MY2c/hg/AHR74wehZawMv9Iygbo6JxPYifkNWqZFaRrUKR7BYPe
i88fzt2VJzx83mwmvAGP0L9v9ssjNPZMCTV3sZsS6gbR61aey21iCp4NsHFm1bfU
IoTK4zBu6DQPD72iMdvmf0cLhIgZCu9cZ/cBlM6fqAp5RNgzvxeQCfl3vquCW9SM
YuJ8lc4zPjk0uP9s2EaiYNJfN/5ijo9npvJJzsqRn43xy7Nu5Ia9hc82EgRY2G63
3xd68JuEdgDLNjVreY1jw72H+Fh5OdIXCHfN96tPEonxdq3m0pbmepROSt4BvmIz
Inb8W/rtFudsG/pA3CxtNm/TTwgfoNtLpWUjNI46YYI=
`protect END_PROTECTED
