`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yQhP7L2VBp4PqRTpleUaskX8lRavI35fUBI6+S041a9c+mk11gfT9kSRdVQwvz9
rCquCQ97l8rSwfGw0MpmlKnhw9G7jMoqDI1F6sZp8fXBef0TX9oQqG0IU1MuQONQ
JhKyNbhLyLfBXFEc1gJxq+ePDKmpqvuL0e3Qui0/n58mMSw4/o4vx6SqGZ75l6Nb
agIvpu+1LQhyb5BCUbsAh5oszrHJnu/rj5OJOf/VTJDU2DSOXh0hbwH5Qq3k3VKB
XVB39N7xsiPUcIMihvOKiszQVS+s4X+GGn+qzwOliCOm3kkZstAJ1903nBOWb8zE
`protect END_PROTECTED
