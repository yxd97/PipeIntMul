`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7M+VhwfoEJkKI5KwCn5JcdF36qvAqUUL7K4rRQ+/U8vQGwsYVVB98UrqPWfxbTA6
LFyEyln0dPH4zo4MIko6X14aKGFfjNWlDFOW2n1lcyiqvjbXfF/hYMPHlXLAOILB
FqTZmqBxf2M2Ein7qrPjn8CcTFLhAqDdI+82EUfWVgL3VcvLd45xb728iul02ItV
jSTNFy0Lq2U6m19qyh4YLRlwfJmoj7TQCI98BshgKDZpyWxT+HNaUAR8xVwSc8gp
6Ekqt3ZzFYdrDEGmT8Uq4aBu/aulc7M4h8+6dGvnlQkrVshnY+y1IwCArvNq3fFr
khO5cOolk0UueSBLzs+T4PvpJ7N09ho6r4rmaX1TkblvW9BpgUiVYVZDqIlhK5aD
DxkvK3MBZyFNOOmS4mtgxA==
`protect END_PROTECTED
