`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AnCKY6qD/5Ay9oIBkYzrW+UsX0uhYSbkyOIpr/t4NAohIUd0kxppsWKu2mqX7hkN
/m+Uh4ts0gMr1BUZYWVHnAhYpdqGuHy7J9DWrtbs/YBw+NA5sRvEVGoF6q2T88vm
rkwUZ97VQz06m5UgrcP7DC0fWD+i8/rAmFAF1JmtH0LKFC8mvUEohm0VwM6Q2EmD
8Tx02C6cGC81pTuPyiMraqizmWfwsIvbFtvcXP6JlfvKZL+UIAMMl6k+ktTK6dgo
zt3UXZ6D+wb4RvaIScRX0G28N38Znn5v/M9HY79c4Gg3vCNNxla35bk/nDwSt5rr
cADnTsT0o2AGQmr+jaXtDFoNFZUGzTkFfBLNFclCcPtpyZ02yMHBkYhNdC7efMzm
jGY3xCbk1bSRzEvOUozjtw==
`protect END_PROTECTED
