`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4lUZ/KSfSUr6f/hM3+C0VteSattNCxLLYoxyYqtnG/8RvNFvxhBbUJimKtkPcfN7
jgOdu99GcEkSnZ1f3rjL67j+qTUHeL7tQuOssr8nlSqgkvaqokqlRqeY6oYf6CA7
oOh11aRg4Pn/bSf0gD0vg9fW4oECc/IdaBoKfUQGJF03q9ArszaeFRiPqtN+/Zi9
+yY75b+y6ufiBzREF0731pnFNeqPbMm6Q+Eds8iu7R1uu1Jk8g1X1DbbJmlbmdef
okyjcUJ44tliKVSWNeHEQ8Tyd2/wK75MPIDqcB9r2rI5jWQBC4BjD6IWW+6sm/qA
LO3mTedO//q8Z0jM8JMXPEitjLPVWnQLQAYfRSJ6xOLFzTYANulC5dEDy3uT0yBu
HAb8SUIcfgRvE5juGHMvUwyUilL9IURNezPYI8YsAiJjqDwRR/Ti/DxnUb47PObD
ZOzkabULG+CsJMgez6NDyO3SRxQ644/CDK3fqmSg43kTy3w1c1+wwjyBXehUOS5g
Dm17x9MSX9nubOGgY/0XoAhEnCyP2FS7883QpnVqH9R9aTWLEpV1vbPmd7AGKxWb
qyjGQUMZ00egRBqZYb3bWxapVEyPsTj8NVpaf2AeSLcSjvYM6Knta7D2cYcvanWV
10IdFrQLHWGjA8RijmKHrxqdT3Za6tHMyCuSP9gofy+fqM2MfT1Hmz3upeFo0ccd
Nx7ephQCtBuN5Ehxn8F8FRhkoKtar7PReouiYh3LS/Qtolu9U1KBfhwtj+FGrM3y
CuUCtuElcGzKhCBBSG4g5AZ2EKgGbzgPeZtp7nxMj/ecNhaEUNePiClKHgi/HzZo
og+oJvGMA3Vcuc6QDPOlLiONq6FMxdSwS6ZtM2CkVPZqNWx20novApi7OTQJ5S2Y
G/lcBhHO1BuLveK9ytyrUbdBRwRTajiMWB87psXjIF0E91vd2OEdHN9vETXMRkt/
HcNv0zQ1N6cr23Gdzh9RayJpM6yOMI1EhMbs3eXBQvtWgDCG4shyHSDbaqBHq0sb
Dy82+PfHklhQdBs96usI+Uu99HxdD2mw5DWiIF1qBylsLhUp4NQ60dDoVm6Pndux
K7nyL/LmYBjpH5D7BVNIk71w93ukcSTHY80To2JZ3l6J1aWdanLc/MsQonVPwafm
GNRtG24afOqfQDOyVcROoIHFrVZ7BenhdPkI6MSEgu6K13Ack0Kxa/LV9MK0vHMk
tbFK1LbNYGJVFPS5KMNoIDQTiG1MbK+R8yD+/Nsth3TE58gthe4VND6TZsH/WSRp
PDixJlkK1XlSFqknHWa1rzqrXf93S8IzS3ixgS/3OqYf/ble3byZ4zy9GyN95Rzj
egxVskBBwX7qo/vlQnZy4KLaDxr6z8WHL/s1MIi2f9i3nZXfv2MEZaLeb9mW5uQA
P10WG6NV4bJTZa0fsBNNJCbofY4Q8DzYBjuwI5vtZL0ozXvHurax+s8n/Loe/Lvz
TKg2NenkdmqZoUalp5YUeSOnCC3XhoVTNNoFWSvkmZiHlRdZIfU03Yn3oIpx7O+x
bc2Dm5AbD2fiZIBJVozLswGSe0vkx9M8quT7CWkWQJEx5PzFlhm9aj2NweBQQSZL
0WSK5hR8XjwvAoSqS01CjfLcG/pL7dpQkrNyJ0yUgnBbq8Fcexyh3/Fo7b93wIKf
Mf/6d8v7ZzsTp1QEKgpGQye8MtjAqdOtOaaji9cEA9ZvMYZJYkze0GnGui+PEmb/
Ms1Jwxqpn/ecsQa3yuveujTh/qfQqbMX0DsJmyyA5dXzCEPg51r9dIxQ2pLSCNar
S6V7ugcYeto1/FamhFhFkAhLRWWRVeUdItKxj0+Hd8MUQunFxeLX06EEXmBa8tFH
zEyM8bLnfVXm+1COHGtPox/jiAHOpZY7YGHXSrgz4Y9Z5D7DlGBp0x35ToIiSfHC
5L9q+y8YtCNxQhM9h/jofCVFq0I/SiYOS11T3CDp7NdJmw9laWgYDYovmVTRYLH/
SBjbtN/VNOmMYTZkz3tlujXqign5KGI7byvf3UcXFYt+jBXsMuIVZy+Fdwwu3cWx
hysHOWaOV250kbs5FfK6jdHCjWghjD9LeSn5+2JILA27RPeVGVH4INoEF63S8CTO
EnLnvmjT9iuDcigrVE21fodesShg0837aaPqH9HFJpLqEv9rDxZAD1VrY1eIzFln
DMvwc83Ev9yTbqwXIQil/vQ3bLJnVqmKLolXLQ0MTffM/g2Q3FpSfLzuYXkZ5h+W
542jG2BV/xi659uiTiZLqel8nx+ocs/lj4Uo9E5GyLFgl2B94qwB7ED1jrEewD6J
r4bOKne/cgM4RPF9W5XmKwlrPKJSm70kf3t5izAd+0KzlfZBO7V8pihzjIDlgjBJ
PbQmt89hSHGRpt875t7sLQaHJYSjZiziXr6fXB9z8mNZZ3SdQ9TE0IiBaCq+wh0P
4EPNpuMqkzGpMbG+7B+vVYVAtRO9GaxynuAsNd0vCtlUOd/XKjhTfUyxv7KbH7k5
P5BSdwXRaBn0jybYO04q2E0LSOzzLH0kaIw4CIBTfxsnXgiBkD8u5v7OObk4hq3d
N8ENgPwnU5HppoKL5WTR8o1ffIMqVDPFPqls5oWuyfpIIvzDtvHSpL1V00ZWAGGm
K993UqRClyvbt7RqdeCAYsIeRz9elJYHaiQpWAcMG3aHLyKEBTR9YX/9ZvxswAOA
EpvvaGZgoAbh4j5oFfjH2YYwuWL4ecZ6Vmgns4dtXkXAdX56SG0c1IZclS+kwgrV
0UbB30f3vbyb49pOEJG0ejqUK3nJoGrRGvTmAbiSG/gl9SJVy9u0mcxyBp3IQs0t
WO8dP+ZzK8dxBMX3Fi5llQzqd379YXdXRflrpYtYJFilLKpprI6nJV58LeIp/9ko
SOFuPcvoRu8713NJf0WxnFtMHvwxDuFv87J69t13Po3cmoXimqWU9mGwHDBMd/uI
WKQlsohT7Cb+FBP6j0TqAVlHWmaCDm7KD/hdh4i8+mg4U8xtD8JqwJq6PVLQoF4f
AJaFGqipNv0hgBBMYTTRlEw9ImcpfEQACgvbZelW9j5zBCbDksjCnvfz42z9RwqE
g4rC0Sf7KQwSZZkbc3Ukgef/tMilN1s70cSIc3ZJI6DRzZLP/0HzI5n+4My8fbxp
rHDzli3bUpxtGyHb45W2HQmNWtF2JI2U9T7a1vPoKAc=
`protect END_PROTECTED
