`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vARtxDIn/lNJGAY2AlGf26KU0ryCw5X9fDhBHUm1K+7BC2zRp3O78nqhXGWHLp7L
HW6ZfgxeCxRFDsD1VgWmLDhswqRSqOoAfitOvacq9mqaVmBM36nrmPRRhnFJ+SeW
4Wtss2BecZPF5SvYMgr4UfJFJyrJCI2mpigh0P+fJ/Tcw9LwffG19jfFg6j+xIJP
2Ouovi9dOQKHKJAHqOWcXUnKFCatr1oE5JkFZXlaN06J+BEgMtVd3M3yY12KpVXs
xUDtxxZe1DRmRzirhJ2pM/YlPxBTvVj7ZWCHsoW/TyhkK4Lw5KdO3/7ttVV9NmNk
IEm0bro7ndFbIMDm3jm5DRMW0oQwdWz3NFx0UP3AEL3o5IWKQiXsosJ6syR+o0u3
Ky+KWXWuDq2Y83/TFRIr8iU9/n3APljwkPjCbQOgZKOhCw3lfAXQ5yA8u/4CIncN
0YP/XHXALyD/0GwidpCpO0Ow4EydTKzVu4CUgCO2xpLLTsnUi3qkHW1BEfXGeyfU
V95XjM6NesR9fIuq3G4h4PRyzvqKj3Q58veaF7C9u42MiupbTZfyS6QsCTvv0+aT
xSa2CGe+a0HlDpHQhgy7olO3Fz2VSjEI0khXMpIe1FSPdD6koTGhdFpe0Jy+R4Ss
goHARUdOPB3tgmGRu7QRUNtguV4Aghm4JjkVKzXR9F9+IFLENi7VbS+VX/LxUpzU
IRM42qxEnujeUy71ajAdRIkpKdCB06uYLX3lEbCB2Ys=
`protect END_PROTECTED
