`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JhOkHkcyxEvnJgz5XFzpfP1Pj4JnzL5C3ZPsgGui0JidaZxjlioaBS5fzl4pnc0F
JWfLu94qSX4jujC05ohWGK51QBWhzafvXsznjUmIFXICdzLB2EnwCTZYsrW2XIac
5bEHs+oQMkw2q1nBHI83848ryERQq978YGS4SKiBalgLUPBfRvFzEAJ9aE/jHsiy
cniADtEYX+D/BG5fntaKk/MClAvo8eQZ05A/98GR0QBxyH6WozVbqs/S68UmiYm3
I/3zWDXZo4IqrwuhOPdevTDKZJ1bXnYsr4I4OQtQYuWwWO075lsQtphgsD0soM3r
vuQoZDjl89Qf3CmSS+b2jrXzS1Dp2bpWKuN6XnPnVbo=
`protect END_PROTECTED
