`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OnMoTmbQkDvUJTjNvay+ml+2QPZkK7fgOM1Sh3BPglyaEkuKT0oAysL4WVTj4F2+
j7Adk1iUxtLMFFGoI9mrGH/9wlqfH8i4o1F1TJYg8udWnoI3+lwaNA3c18gSuOqX
4AuCVbCg6wqIN6UeEQHDva3Rp6e2S/mL0aCKdIxELeapJjrtqvqqDZEYTxyOuYYz
FMdGH+Fy+ry7zxX64nybLta3G8K7pTvIokepwfAkzLxb+yMbWr+q9nJ8DqCK7wYY
lUDTC1cq53XlmXN0XX2Z0UjNjM7LGpNJfntFUEVF4byERltMGmMHIE89BmbTVFbR
GTQ0KJZS52jD2Qg+uAkHOdg+KmOGbeAaaLmgB7wB8pL28UyucKo9z38aeNKJIYvQ
I/OZvxlfAiYoYHKFusj+L3Gaid2iuBC0cK+wZeDzTRlRhOjsHOBOqSIOby1fh2Pn
yO3T6mRc8nHZsjysibo+NORljXbZxh69JqvLybubfT1kncGcHGmoI3x3EpL27F+8
`protect END_PROTECTED
