`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTjZpiUpWq/5Z8bRMyGoH0M4eSIa8Of21F6L4PriivyHg44sD+3i6y86Xfk4v7jm
UzM8/DoqTUrQ/duMWznlPxy+qj8MGQjcmHrldWaFY0IECqYF4OCJf/gMKQYztuNn
rIVKnmvvuhEmjYtLyqtTyjw6eSv7jQQtQaM5EF9AmFtyTUCqCu5EGLGqwplALttv
qf4JpqNeUzwqZ2Hlk+2H4SAF0iYWL/pgkRc3oveePLv2+9hJGBa5bN229Hj+PQyX
V0Jq3x340TfW2ldMPwi50CvtRCdYL8q1CitHFI8lu0jhbOrW984Lh/KGuWxQk7yX
vp/ha1ILR7trlFEGJrhYfvwFBuMrQrOOrXY4jHFOUdSvp+I5C2oAMJ4nYqilhrby
tphlkua548d6T63yQmyZ/e/GlFCyHcBa5lYE/LcJauV8QhK8TsBIVc0XelD56Thi
qvv5l86I6jV9VBpyT1ZiTNfLt7hWKYiaprZuzvG8RNxyutDvNhwLg+PUjKgO4o28
eFEprEvpHvBEcfMbk7F6AzPworKUbRiMs9wWhWpS8XfnpzgHB3KWPMUe+dDegGza
gAn3zGE9axrjMcRbVas3prNb2i2gNfnZcIvIsppPxdYWXbypzZ2QaU+37ETR/OMJ
DsPEdzvYN0aG0vL79YldFA==
`protect END_PROTECTED
