`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pFu1Hv0Mupm0MkwCVk2NO7rkjlMdjwSK530kTDd8a54gczW9/SAngWXlV926gMqm
fydiDr+iYCJD1N92vTrwRW5SPGwvD0Vekd2YOl2RY/rR4SSK/2CPdej/uAIfRoOl
Da5a7m5W1h7gYWoqLHTh3xo+1FDgBfjEQOugs8EYW2ir8PA17FUd00e+PvMqGzSq
M4jEh1T0jz43DkmT/iNlJ+Noj0qx6waCgwoySUNYJSrEwRFZahJCFsqMWWqz864p
rDfTUPK89QOc22z9aDuwNvTcygugK7EAg0WfzpaPUQrlInqAUlmM1Dgn9dI4LXGL
VIiZwQLZishHpHbCvC2vtni7LMnmsFlCE2I4m+s9EDQVjjz8HUE9IUMMuMv4PgCE
1h6BYf6HRJTxrDnEEEkEOiiVsEks14mGRcykKFiC4LRFrpoRfMZRZo/RFzkpQKII
9nPb4NhdUjF7MJrJN0EG2SBc+zDi594Tr6B0Ebs7Ae8lSgKVNI8PfYaEN7PIhf0c
iTkIhvIrUah56Y3XsGkdE2SHG54RIRfPiLTXjAyLraE=
`protect END_PROTECTED
