`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JKHBZPWx6xsQ1I+9E3l+RbW3DPLYTIaQyv7k18XCeD91/NInhQ2ISJyZ5WTOR94a
Sty+T1qlGqBHMwWdpZgyvTqCIuZfYwGWPwGFeqpyzjw888IyetUd9O6dOVE1wD3P
m9tQRBsD8GLsm2/cBlL80HlOrhJ2ldr1TMCTB3QV6aTnccpcj0FbIeYglU0E5Trp
HaBpdFBvUoXtwtVyGZBZHdSufYxuUSIvUSqiWjpSrjl9+xhJogJTI0OSQi+LKoDu
5HR6Ot0o7jOkO6qXm9ecm/d7BQj7PzYHzvyz4IO71K69IdLqFn3Hs72SEd8PQOoi
b4u4q6xsgzG4DYDo/NXnYg==
`protect END_PROTECTED
