`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/oZlylQFVpRVNd2+F8wIClyUeIuG+TqaeuBSJW5e/NWdKiSRmHIvYLnwUrElWHAB
xTHgi7YoIqZKoRVUVuu2Rvp17U6JBZq2FkPThhGzlIBrSN6H5BJLoAEbPPbNhP+8
8Jq+WjA+pZ6tcXKTbic6FB79ZOlA1MM0K/v/zj5u4+/ebor5BBkdomRAZzveAnYB
GWPDYUE5511Rbgl8E/UNQUoMZwQsJ13vy2lvDbzCset2tTGHvo/tbb/51qKoOU6U
KZ4RwiBcHW6jA41syKA+gnkdMqNKCxtec9+aiT4kOyxzoQOvZpMuM4youPdF5C1r
KgBYHeC7fRiBcbVx4XDOzIqaLfzZBB38ypJ40Vdt4Ov8vOlj+mqQZc5+VzqBYMzf
m20H10KfO9I/fNooZ3kutwoNI8uOlseKK/WET8oWK1g=
`protect END_PROTECTED
