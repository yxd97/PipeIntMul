`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSHjodFHe0srAbQDweMoDDICARbuE1f5Bli5rLuWk75H36z1v3kXm9HbyKAqj/uL
RnvMAOTjQyQJXEAHH5ab56wxEedWm9K+zFJUC7zhCj2amXyJU+E5ObHtFKACwhTr
6FCjExyeaxD+OTkQF0DhTMlzJirlp0izp3AQVkDwRQ0GU4gRBA/zqK/lCPWqEpf1
C9frpouknVjLqfhwgnxMCjCgZNCGKfbb15ee1x33Xq9rlZa02iMeJmlmPFE2cAwm
+uqIqad3MFmYefqiMNHH4q9c5hktcSUlmK5TU+vbNH8TjLMOzzbox96QVtSRtScp
+JxY98R3mcdCH09K9sk0v36CoudEyw0OqIeiG+LQx+OdtdXrYsF9xSY5wBkadTnb
5//x5taGas3me6ZaPZcZdxJotBY5FFNOAmSyRV/IObUG7TJR8+5XKFnZ08HkGKxj
FIpG/IqyNcYVJy/ljFZWccYITaEPsNW8Cfsy5/MEbupPOrzSSd7yYusWPqinfOTt
DWHB1rbhYohxqkXNaNsPsA==
`protect END_PROTECTED
