`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sieFGkwExwiPzFUnchE2eljWgwQsXpI3ZITQF4olRHxSk204UGRjO8FeRyQGGrKw
5stY7Ben8TrCA6VDIb3Y4F/liFu1/FJHR+6jMbte4ZgCALXZgRdLHOJLEz3Ea0ZU
ZdKlVuRpjoIEfhtn4BBKmvnnSYST0O7iEIVut5Zgd9HfGxrXM13wNgnB1/mabkr9
kmhREApPCmafgGVyAdQLxc9NlaOPXNKqgl4hWTVCy3EuYPmcTgy4CCnUbRnemfzV
cbe58egug0T2BXJm5+ITjMkRHsjPIwKV/MSrUXEDCz1QWHfiaXU5T0n5hp54EHgz
5jy6dgJpILQK0Bhxa70XrbchFOwKDLZETE/XmqIbEuBqAnSOnhJydhIwJnm/1c6C
YaUGjN7kLaEL9aopLTA/BpiKSMT+g/gFjazzSK8Gp6Rbs3snZsOCD3fhUJInGljf
wtF2t6CbS4Oc+Yzwnk+CCZPMEazAKN4rA9F4BxoNxjVnFWPYXGOkvMFZstARu1Gn
DYJswn7QIIwxouXXZt4uN042RJ+LJEa81R0GK4cAImgOdflzNXCMqKBq22epXU13
8Ke6Cpuh0XKq9omXnTz1GxebECZxQxrxURu1dK1rFOQAelqMAL4chnnNWw3pvxU+
xESIqwjVkNgXuVm2X+rd3mE0VKt9hlai6bDmoJoQY1oLl4sb0dhWqpOTCEUw9+/B
4RIfKkn7ifDhXWqR3VBMe5oXe/eXmL1lNln47+f7RJPx5RhN0cxVQC/NPry092tN
Ub0cgDPcKiwHk8Sc+aOvLdRbD9gLe9cf3QXnPZ7a4t0nmjr8C6cg0dn3lnxuj0Zg
J4WiMVueBX/P9EVKuhXv7+GlrqwJHaAKrtFu23NISECruybTzxLnZO0FIEJSvRko
zxGC76QGeRy3FF3b2VADjhleV1wiYVmLC16nOet6VFRiKpgBhma0SpaUUz6s/lHc
rG3MViSFLpgxahXQpMP+WiM2yo/TfzLTt/2T4h7iQrGT/yYbWpq3/U1C7eoKn7r0
xWALXo4cyWaaZR6eXGyyf3DTOCHxMrXvAqO0dCXePMJj9smiZGs+lFaMk9xvAbpn
uQqkkgWhtmEYbidntJMk0Lz1ZW6X93bqx/vYxl0I/rLyAmwyvBZZxcyviTgHgPYM
DolPAl2jIGOtFmdQeGJ9Nx80YmThb1Lt42JoFss2AQBT/pcsyi/q9Y/1pWhvk2g4
Q3ewLrBS/KA9fd/OaZ6uzYroNhMLOChB85usauWd57rUAf4QgrGIpak4D9/lc//s
JhV4auDXRxYVR6uPnS49U2BjJMIDVl8G1V1f9KAcavwA42Cw3hGEyQkquk9SJkaG
HnEZc874wXdn4PZODJZZ3nTjad2pDkIclX8fkATkT8fSLzvu2suYobsLixSf9LrW
mXzzGYl5FRwvSiephQzW3czjUmZKdJX/+1f3QfBN84VpgmyBFlO7wqJuX4esG2Nn
yCFwQrTjIrFzmxbI7/FhsS8rucOqeQa7SHSQt18sHJvBkLoth7VdYAU9nJR+Lr6g
tSByZX1vP0qLVthZFnlkJmWMkhqQC1+WTsXp7kcoa1FLl70uyRCF/TqG1b7T/IHd
2c00LFSPkNMXNSD2Wk3OsDP+QE/CeXYnh2VMhGyRevTJs8ZZ7pjDLOobIV5fZMOJ
5/0/+d0CXkYtFW7jRTw5b0EOOc3TFdshCVry1B91WFMg4TChnrV9DKKRM8xc3F75
+7wdu9AwgSe0w02pu4xTrmyu9BrOce11sKcF+R+QXX2eIBpxSWFDnrSNYvh1ZiD0
8V19vss4rNB+rVErGh2Q8kYui2mM3itQru+w7KG1xcihCfZxYUIXMl76cdoUwF5+
53DONh+YG3rUil4UO8hHTlHdYZN4QAUsfBLBwvfuax/fnI0Y9MKCZu9rUiEdBoE9
op+FAG4kSqiZEwGwo696ZIT5QwTqv/Qr85M8DwqKMAeJ1btCD4j3P4AGJAjByX+w
pw1TgNJA9vi/GNHEzeRpwO9M+SebE9OVvu4LQi32WirKoNwLuQUh7TV8DqachWdA
ZCCIz0Y1zfkQeidZfSrGvowRkyOcV66DLBPtaLq1WPSVQ5ganM1t5/s5w1Fewq+F
qO6qbmHxFHC64iVACNeJwinsgysYBnJ2tofLoW731/+pCCKhjoMPoXh+c0XCtbtV
92s/h+JO0FZLzfEVwTLNElIUmWQfauAT30trkoatRNBRCbT44CA+/+ZOy7u262ZE
soQXpYbZEMSrHtAgGuC5me0UPFSdoa/COzM6b7HAdJz5Ya4b1tWxuIdd2NGm7Xh8
rslHI2Gg2MfZrbq3FG6sIgA2TJdaBmyeBn6jUdnsbfI/qnAJCT4KVEjoFh41iCOV
bDxC/nzg8NTUjLVyfPlyj0b2r/leBxjE9XJEgjadzKWwEhryZ/8JlgqA5nAEkCZ3
xq+n5GchjDAj0JrhSScDeXy8xWI5BmMWOwfB+j7bRd+JavKd9LpwgJ6axhi6XIQp
VlR3cB6H+cY6jWmgttWFNK3Tysd7jVfYyFOvA8z6IBQVwSRD0M3+fAKsKNcSyaj5
FEtoRwmFwbUiA+3PZUmGrPDOWGw2MJX/5OThZQe+tWTitti5kJmJuf+6eTrzqWxV
DukRhIbRbFIzAUYDMPrIYxa3TryoIlafc9u4+TvI6cPDMEGw/fXFSQBx2q2VId4U
XZsqirV0xOfSl3hR+lfuhoAjyIppaNwAaICaj+MXFTQXsGwpfYoXaiKTahKF+oad
8+eVwwF4fEV3NPGzUUnajG8VbqZOQ7ipAs/ywuDhgJzGWhEGqZCW//p9+rTmOAt9
qmw9HG+9b+JHNzZyjDal4mcTt/atfjgf+haeMT9WNf3NqR1E3dGUITkj5fJx4dIt
Wls/BfI/hKR5/I+AgakOhxqAbRfRp7gq0h7bj79j5Mw=
`protect END_PROTECTED
