`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SvYIfpj5xgp607wqV7QFC99Xq95W27n+/Sct1emFCnplBpcP6hYXzUkkqPtMSYd8
FsoI0lG+b+u4R8sqkNBndJ/qSn0Z8Az9A7LmWsytHbcR+MXj9x4M2bJf0Ou7M9vN
9XaCMeusVqb3XIj8kxzoR5TujLjAif+0J1j3LwxQP6Ra4ZdoeRGH4elV4HB0oT+N
sputVaaOsJCH/Li/1oIOS4HsOXlwzYSdJ3D2Lw854Q5Jd71ak9/VieWleXaFIX+s
J2XLjeEbbmUfHdBC/pGk50aLGaR7xg5oCYS+SJ+G/QFBuv4/N8iYl5jy63fp2L5k
qYz48VqNEdx0V6d54WP8Wvm3H4omM6Eo29cjMbcsX7jEBMxUGDGGaETnG52h6b/G
mde7JmDGOQhVrU6JyczzCS2M2TR/XJL/dYvOhauZ6S3sOTZDHjwwXKt5oONZK7km
22d8+cwOa9TyePosFgeiMg==
`protect END_PROTECTED
