`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MX4aDxPpVx/T4WXSXDA+K/gRzo+KuXQmBOUgDHxoRK3sL0OEUKa+NyCKi4w69UJG
9XT6UALCZSwqjOvxR0yb2KXCMR/4Eq37nmFxbdgWAxybaUoETqLxshOag3jevaSI
TB6PHHHuxs4TMj6XcS39OozYT68lSlTmfBbUTRlYs00KJxd8wch5dG7HJSMWcw1o
Du7EAyrNx/4jC6brpGw3a2hDJS4wKLHffwn8v/r8BI32RxAR2xi6n9/p1Bd+QGNN
Y5IP9fP6w3yANJqcgUVxgeovjm9JPwpMrMA7ykEUSiuv6AFjmrMItJG9esN3qIUO
HAQXrK8E4iWV8MDzellkZiKWwVB0qNI4/SL8eiycCVQ6XELnoPISh2sqJCFYt1WR
xE2Ayf9TLBfeG34/o5cl88QSunCte9DWMDxMiyOOETWbJ0fyj7cxZD3gFall9jS5
8LrME0cElahg0VbDmqwLI6LbiMHzL/bQwR4Y1ZhCuNdf92cqz8/7aVDRCvfJpXvd
VB21G3zykU8KKHnzuKBHA6/xmJupOq6Xdv9PAglQ3LX9dYJKrTHq8FbzxUt2MyRN
7tQa0NNpqOffGiKe62Z1e9Uc08ru7S+IZ1SlT2IeOgAgUUlcTUu4Nlff6CKkoeJN
4V0bNkc+cWvCKNFu4mS3uR49n5w3lyo37ElNvmk59tk=
`protect END_PROTECTED
