`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
utnhDjuV9leAY2Bpsncz2bAbBkNcMgmr0rsD+emtjCMMU6fYxEfAerB1U3Ck1FD9
U6zJ9tL1X2hyGLfvVNaGVaOTPeMTsjdHrqGSHLJ8Occ1GsDDDID33uEAvXNh93df
DFcjxd188txoUxODG6O6RMyb4gTKYCm2BD2R190TtQAuIZ1u0q7YvfKQWYSDLDcV
zYP36KFNxqQ+ZBnrC+FbVnY5RHrBrbNRn533cbiBqWQH1O4xkqg8krJQdBl9WNao
BOHrvIcHIPdGQMP/na1e/zU3ju3o2WVtFycTI6s9GSBZoHrxEgeYcxc6YT1erTOe
bVPlfWLMRHicqGhksZT/bmlZXHmuZTlkgr9c83zgBOf07dV2iFAluZiVL6dG+t3S
S8gdq995/Wk511B1F1gjmuEHeEmzN8/wOXaGO8C/Tidcycr3hZF9W8dvJNx7+CLj
arpxFZalKFtsPX6jijPh1MuMC/GP7+Fj4XSnRfP006Wxps/eJhgPj2ufAGH61j+N
++OzCJjKUWkR2FKh1COapm/kx3h0+bKBV7gw2nuU9TlUgXZ0eqcBczYf5p4GEbik
vKmozQ/rUPy+bVd/wi/1MUEYY5+DLIejbRRtgl9WAlpUfJLw5fCQj44+32WWWTHR
p1NGTyYVDlfQdOzT67GvyoeAoCWxJisv/ypyeQmOOCbx2BKpwCv54N/u/OnE0xVO
sbY8hl8cFBxdPKVjANF5g1cShY8Qr75f8ghNhvt1lpixor6yZqq9L2RmB6PPRSyk
l+JUPECNmkR5cV8AUTLDgA==
`protect END_PROTECTED
