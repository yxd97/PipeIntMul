`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CpN9ATIAovrFYY3V6BZB5fQkILstLztnh53TsO+VbJkmdZ+6OiiT8IyaMMhArrMc
AA9cIf7yFIgu2eh/B+bz2+7TGb8/0C8Fe9Sso9phtUzrGM3Zjx2Z2gLKHNX4HXYH
880oKBS+VZT9pasFDUuifLyO9rjXWrUNtXRLuLmReWsrux3kewZS3p/gp2RGPoVx
7saQqljEPjHdCwSmOletak054LfSLzSChj8nFn7vqaYurPfIRHwJii0oPAMonMxj
9ueoPsoNjkr55kM4fC+LeUZ2Q1DKe4JWhy9djWgcyGdqq6QjFoKAjwN6r5bAsBeV
0uHRa41GWVZO5qoARAZmneaKThY1zjI1yv7B8GRriYKNcuUqdTRYEMRwPQ2/ofsD
zHPFhGyJ8qi+9hgLfBRstYS4ZxPTsa/v8omVup6dQYxhMATevQjwx03ZamDLA8YB
jfXUvD1WJQbJ5cAPeLMaaZJC6EW3Udvt1zcxx2ifXFlrE8Qj6iPHuACwC9CSsQ5E
6knWaXRyUWngA0894Bypjhys18RLJR5w7lKSJbo+Rmf5fjwqQyThSChhjZt1gsWQ
INblaRMk2372MjaDMo+LlAwooctNEkk6COO2YXU5km6GhaKCZjA4vEAwxwb8tJRN
UUZlbwC/t2VVFkspeFWISK3PmRbUyuYa1OAbk1ZQhlDP4+oT4USse67Q4BFA137v
shBvrS4Di4Mh08xmoPFuEvfbCGGl/VD0NahmPQjUyFh6aolNkLLSOk/6Bbfq3ChU
CrMiEcB3XwoF6iCRqg3A0YOso/iWFuDRzD3MW2cFP0/DMgmMAFytoOxfNoXNoY/4
ZE/HWATNcuhOxGKYSUC0yP5mrFz3LrudsCkyIB7Miyjgkw2USe+q1BCM5gAl6qyX
Ee9ZuD8BZtBszh0SHrDGusrllKWp02eWzZZDyRbxXmc3EKwYOagIvwlAHwpbtH+I
K9k7yNRqXYRF+a2hX1shlo99givAadIlkrMHAZuzXpQpBcN+pnQW/l9OKFC7lDSz
+QdGwEensKRG7XXqe1aFFr1TfWwDjLLmORr1Gw8bP4hCqaWllCTK0dSQvm+C3rxw
rVWtE/qmRWh+WatrToAClCaDqRT8kCinn7jz94Npr7pGixIQFN5kLVhgC2MLdmi/
OckSsUOTkpCXQl5dl94q4Bh1Eo44bh+AiDy3JTWTtD1AgtHkcKyb9N7Iyl5iy0Qf
Vkzi2MNqNKgch+axUzARk7blNDEbYzmOGYtIClSXI+zS3J+toraleO02FzaUyUVd
oFO4Ew1peOYoGVsdMEmEv//iPFEVwwHWvkUCeQyvGRkYBAmHAtYbR9f7ew2HZFTZ
b+jpvnVKcpA/jbcTVyev76IONZOn6uoV7z20GCXFX4WVwYivte4je0EuwLoju0GT
YtPdmaVtpt3Y3/ixKb/xMkoanmA4bK/WW9ujigRCvUlDujrE3ongA/kJz2rGWCG9
3cms05vRLgPNDuKDrj97gUSdRNc1xkwg8WcI7WUoekSWR7wCrnLIybhjbGIiR5nR
tJdGhv3K+gG+6NuK2Ry/kxwFAn1ChB2nNHC+gY51nuTOJPVmZW05F2ApAkcBKN6U
ceK7UVthfeI+r/GM1Mfgt2RxnBSlvfjT50zploQmBWhAtUNvNFWulQ/afDPtM2v7
H4q7+hkA+9EMOoZugRcDos1UvzEtbJJm2ZOe/Xn6Lf/7s/GoW5deHeW/pX5VV7R7
LqvoaT99KqhHPAZYNdYZNhNlWlDeeOqDSq3yyoDeL4MuRx5q+/5Om1zlgmVi3yXa
sc0Vc2rsMHyS3KUTNShvyzFTNJIzWBr1jIP92hFWER3i408TC/tq75//i+ZjtuwO
ud2zxfVu51zjNUTg/MK6pSiuRz47dVggGWjVqg1UyrHIReBNH4v8BJE7nOC2PAFR
sIDO6AD5rQZfRHibjxGqvfCqXvy6VHNpGY6V/nUqNNCTvYj6cata4wQ1DBWUQlbz
kvQ1HlA36gVSetsA8Fc9fgDzrRwKcRlO0Hpfy7quYc58CsLiUwhFXtA+La6uYLNQ
yiG4f9HH4HtuYeNVBY+2AbBJ5kjhyJRCSRj/FRmBNByO6UM9dVYNMxzngbIf5Rop
OJqJInDIMNw7m8EHqZ6zaS33+Ri6wP7vj9L/Ki6HAkDrHPXZ5o84c25F3ZLZWbTv
F00+ZGqbEl0661oRuosDtUNdTgZ1LR2JjC56XplLB7iQSprbkNVprBQJPfbR2eiV
oZA9tXcvTI9r45ix7GvTpUuc+G/qTVymJDNbA5JWftJaMOG7SiPQCfOgBhDqPIbd
L9k+KSm0kUU4Hb9sQXWeg1dQir+88DaJr5TzAPEMm90D6mjra49cLtOvKdyqAVod
LjgigUKDHooQzBpiS/rVsCDY94uWbNdag4bm7OTN7WDVSrG0RV4gyOREksWAZ74s
o91tfxqLyP1RKN4MWD4H8xlJDM1rF0p1RLRqNMsdpML62cZ5/wunlognew5H76WV
doC4rh9pWFayxWaCllypDGvH59kJY2URFFz2HrJNR0aghj2OupWe2gaGyfg3OcuB
eJIAC465ITmjQCaMDV3iWWrBNg+/ReTNCqfXE9Hz2+HbkEV114VVXjgGSNl10ZwY
nn+1h+QHbrxZqrRrg65u03IqzYezJUAKzXGSj7CoM0g62mTDiFKQ3p1WP1qUwmVn
acpIKfwnG9bkZKDIN78V+sd197VMWaFMNC05qI9HarFeserDF6/0U3209B5AaFbt
j2b9DeTtEyFGDmwuvA/BayEMtolNEep8yPWdLWfrMdM2pWyiIGokHxOqymXyTQnN
G3f6sorK3qoM+UEzyw6Pvw2Qdf0boRxigL/bHwHg4UTMFW3Io3bflp6lAK3n7qO4
HGjTeqgynNM/WMk3tegeB0bwfsMTst8Z8HN1dD/KfYiOw9ogvameWPRyUOyfIanz
W5coFDL4jL5cTnRaswj/aLfvfLaiy3WEeRuwx80UaGoc3oGRj/1wBi6KYboJszlI
FOdZwDC71xk+HNij6CydCwTrzY+Z8jx5sdLsTXljwDhYGaQNZ2FBhpAl2Rjuhwng
a6QoFe2dpUDVADUSHGAjbQo266ezqvRYqeSjbK1kJn/UI2VN3PC/74ObaW9jqB3v
bCDMVb/asXfc5cbkDaLXl28mz5TgeuYEw1D/QNXLdEgDm1ndPvFA0aAIbf53zPXA
l3KOwkYRkKSRvyIICQ+SSOJRGZ94DfUxmgk4WwFI/4+ezmOKN9JRXfOc73MzXqMA
UqvXAt+aJNnD/k0IMrc7MwMsBbTEXzKX+3m/F3/Dqdvg+TpA//IB7zJPx2cBWyU4
TjpAgh3DfLXSdnVyBFsEUa6mzK6JbpJZyqix+LCH17VVNSVOLO6LSt7lXH9M3sQu
RhMwlIbnLyVi+/TIaJg6MyAFd1Hka2l37WzIab8zhocYjnU5M8bnN1Aegi6LiMGr
kdsmyBrzdwpJ9HA6QNPWUAIOEfWlIQO2akLJYgelH2Pp2UOVDsCkQWJCUS7RKVry
oOyynlnSyQtjlDMWdxQRx/SdXoprUXVwW1sCjSmiiXlE1XBjMgtCevMkPZyBJl6Z
2WHtAvmOaPS+GdhYy6jvP/khZWdDKn4FSUVfNNH5HMoPpQU5xBIylnm+y7F/Fafz
eOhL53MokMdoYST3tqR8tQDib37c+nEojxqp/pR2h9tJ1D9HLu2sjn2WJX+I/4yV
tpHR6mixtkTZVHM4+XbSIBL/6+svhYeP9PG378smPnFsEfa3tof5oDVilSGX3R8K
xp0V/nq04vr06CwOKoXwBYSKELN1EPYwGMtm8XQ2O/PHTyFYQN0AQa8yGIB+bNDI
boKxbUPtZflzkEfbENRAQqLeq/M2iutndFWJlmUwLTF5UAnMophL0CE1oIMqRQQA
x+LJZH4Ofec5/KHe57QcWqDc0sj9ig5jgJmsc2L78LV3ci7PnR6NjNYTeMmdD9MJ
5E+DJA+1r7TLWf7SL2Y7RS4MkvR3gjkkDO95C1Qr3zEzjztYN6RZ7sQd4qmGxt6D
anECoEY5JW8u/87qZJy9Kca+iJHumS5VQiRJO4/5gavZK7vV8DpPDgXjTQR5WAdG
8klQeJLhePHJWIsHfrpOzI/PXLl4I2SBufbnPGHAtOTtcLpOvFbzDEgXzZDuMVno
`protect END_PROTECTED
