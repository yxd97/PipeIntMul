`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmA+hPHd0UijbNVEcM0PgB6IrDCpbmeEHqub0NdN2ipHZuSX49DZDeN3r+xdji/j
BPpNkmlJGShQxJYoAmuJrdn83F5gtgK03s9cRUXYZeahmcBEAgR/KkJtvt78mMGE
gq9bZsHaG5hwk3VogX64XP99B6x8fqxVqydEgSQAnRdD0ro4IwQoogGWYDcUaY03
22abxbAhN76N75FckAD0k6wu3aNyf9gvdSLYhOmMiAWLAsUor/PbyQ5DyCFgSBgF
zuRAwAqys7rlCc+gHpsclr+idgDL1KmGvMaj/s2bfdFhCZDRksctiQKNOFeqEkqu
`protect END_PROTECTED
