`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9BGlelCpcKYoFhwBjrbbbemqeb/6INI1rYMIaTq1hbA6sJCrx4aIkUh/g5sbQ7Y
eGK1gfyfk8MAwqZyuXHIrp6SH4vnXWJ/XstIA7E6sn3PgEiB3u+OlWpQ+OgTIdJf
xVmrJC8/P+ZozFCRIrAtjRDahRJ6OFul1e2btsGuAf2OKppTTHOXD1OIDFXv4Nb3
BGTLTJ+zQ/3ggZkKAEHYUKQtP4y+8AJYbDvTSX2wDTjjCFmme4PeTaYZlm+PzgNm
1/AlEos3TcWga8qdteWwjbZJegWX3HHPgcaMoWDU8ypAhE31LzmkpKib90gNgUi+
NusWaqePCtmAVN9N5hiZd3+9nEIyywVieG6MVQvF1n/LXO7scwQcvqZj6c+UYW/7
7Ej1eEhFvT4JU1A8dUbMl4oXxdVBHar+l3+aGh0H3lSwecO5I66qLD27yu8ItW0l
V7xNl70gQYKpMaGx61G/706rphYVvNJ8hLCFeEGXjANLA5IAE7IM38CAf1L0YJp3
0q27GXRwJPXr8AD5R0CBcgB0ASjAVffDH93x5lAEVmNWVgK1Dpes/dJ6b/3RniTC
nv9eHzkHBk2ksAA1YZHLNUiehP79GupRI8fiHuQTyXqcEhqjYRO1fi7WCJ6o8HIm
3OV293HS/LvyB0dNMrJ5x+eF0JNJkGAwfyVzjpcFA5Ku4uxvYM0bpFoIvhRTxe3h
7JzvbNT5O5RF5ME1VsbExNF47e/9vv7g9BYR30hIOsYKW1Ucy6Uc8GzsWpordXSD
JzDwfl+c0Ie3CADLlyxs2lrWnlWtdFx3Pp4yTFe89s5eytWU1l6AVtw8fioRup9V
gpCPN/v0sl7E6H7fTq4HOhes5eb+QCWwzbX78qHsorGTa4SI/V1257363GG0uhH0
RyHn9vDRWOwp3bg1m22LhaW87ZFe7f2DE8Rf+TEuGXy7ISu2o90zGG2GPVS6QeFo
jhDHCdnr+SoMn6sd7r4AW8h87OTGKa5v63UVdBDtNHuAbv6mv6eSegLX0X5nNOde
7tPbOCw9EQ73lEGqbknjd7RQSfR6ffnPmZmKv27Dl854ACXEXARof+6D/cQWJlye
`protect END_PROTECTED
