`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pI/rif0cR7nff/PkoDeisrLAMTnAbQeiSR0OUG9tYIH1pqNqhVOaRI8h6/UTf4yd
gu9wUtWMC1f9IaUlS12fdCunBzLk2EKmpZ8F3+hFg9NyGzPz9kWENt2gfSiwbPfe
2RVEtzEJ05tTwuvGxzOB+SbFtaqrRO8Jb+9NoTUMVXNlaAawmmrAZoncgPrSL5/D
6dQFH7+wYfDKK1j9GGdazk2prjJ26gAn3+FmH+TiYRaFaxpAnwDxRSue4ssgjgRn
dMlwYf3EYhV/9m+E9oNkz5HuEoZJgfqhnK+LEzBw5VhIGqe7sneti+6nR8Lvmy06
HdT9Pnp56YDxBsumOjMxxBbZWJTop0J1M99zjoDgnhWxRXR4Wner0Jbm7QwQyx14
`protect END_PROTECTED
