`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQhao5P5FFPeKcM/gtLQP+SgVLM+o1iIGRnM9k7CYRfeCA9JKi74rxV/1JBCWYHS
ctFoDKKdZFaF5L79a4INAF21VK/DIVmNTS2/jSBMjKiM3ZhRm3t2muI+thfcucFy
MlqbAN/Uk/wpCNBimZWie/vpPsifu81rueWIghRNRFOjewzrLRGh59oL67BLSJdr
xjh5jvBIPKeibb6Pt7vmXMrtkRsj3eVE//S6KLCwNMGXEsSprBxwYVyiM3MecPpW
3KMwoGuBOj8/R8j2vJwV8mr24nh7VNTk4lQeLC+s/atujoyr3fXhT/jHmTqlx+7f
wfAA5DU/mpNDpIrA2uqg21DIrOuJKN4Fo493mDmiqBZqcYikive97LRonL4+AnIU
FHIIo+nv5VikhMYRijSTdp16nORqkZH9sKAuGfcUpwLwnS5kUK9U+CEbjbm8GEPc
EpY1Vc/SMKT6hFZiN61DPfvrA/fPwMHlObI55prBLrAJf+xglnWVvxnL0VM7UBMJ
XlWbrVEuFfMOlDFEKXZnnapsbVYaHHKzoK+7DLE0mEmmurZLn/RRUxX4B4phNk2n
ZCxrm39OinmlTbv8fuzSYXFf5cmma0bH0+0PcSmMLuDUqWpDY1kz6RUnzex3bPZA
TtRbw5dnqk87/KLG07wv026d9DZ3IkyF4G9adSl+LWYl2lX7Uyr/T+Dh5mjg3hcj
ImGFkryzpntU0ijCr+FwNX7H/f34yg3U41t1afd7NKnj5PkiwiiFunBsIY6FPdTt
QYLuhyn2QQWiQtiC2iuyyQpdbHK4d1GobjzAuG24bVYJqNw26T+qn1nxz+SBNj0X
U9NP5s9RbM2mo3p4lQ/xsQ==
`protect END_PROTECTED
