`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XkBtohVNHWVYwsnqYFRLD26s437M0MpkG6NyZ9CYPk3QEB3oNEuQuoQPFZNBWwLN
blyT/CRygLh0vNmPNOHjvvSm2k33EfO4+/3NZut9xXDj9qSbRlMiVxrwdFnQVoiF
bAc/6Czs10Xhb9OLIU/k3Wig7v9kIf3lBcNsTJOT4gSjYXa3ZKyXoENoWpXKy3uq
j1Ickbs6EpgReB81SWo0/s4Jp12Hh1tAkTSetuzTqCVsQMuiS3lx4PWvCHXkP+/H
AZSTOraHm8HazPL4Fvf/Ne1DT1uHVHWi9zX8K3GtV286R+/SwT2GSRKYw2gHTZJ7
7HEtqMaaMO1Bi+RewFRO4KjJG0tuyrZdkDRIveZJbriB7Hxr1zMiorF5xe/0D/rI
tclTYj21tUbgZmy8n50YSiTELaORd/BO5xJnJNuVSKTLpDDd/9Fb96E46Yrn0hIS
HvpHdlBacJMe7LDy6AoP1PTGcKgTOQG3hkSod29hysDkhswvCerXKnqzQEDYJa7/
JyYtlUfySu9sQKvReGsWbGvHtPYPmuA5lYSvTUMyrm53OlbCE9ERtY39HKYjjA+j
LEQreQWpURpWlVW7rLfIL1OM6y920o1ssvvPXRdjHIip7isjcgXcfGaWnOkWH9YV
3KFCbMZyfkfwy6R4R2BnnDLOmzv1rpHNruTgHrmF2JQ4W570Zpr/ywBLz0TQqMFs
BgFtWdGdsWrlJjY7GD8BPWFj6GWqerZugpGvp4BBGBJ1ySmHBr3uBtGjrvz0reUV
Au7SrsBg3lW0lSi1Uh8cZLK4foZQQftnQETCF3kC6yZIyb7fGa9NXrDARnThQhJ0
g/V2bwYyUggX0Tv2cwVPr4QmszNZG3Ak/a/wcOVumGcDXoGEAk4RisA8NU3aMcde
hENd0uqI3pshvdFIw4rbMYh4skN1+LCvXUhIJyWrl5BZTF4aR1VdSGDu++JcPTCZ
+LKuac5ne2CnIn2b7KQ5rbmulTf2dm41p2X81fwfBwYrCHmLxICZpa49p4n2MECL
o33UTjLVXQYALAAv53G/1oc2QyuKHr3OEElUtHruuySSIfwPFCR9O6BqHmOQaRB1
ySAP30FFu0kKbKDVt9uGA9NvFocBrf50YNMA/lxhrQ7mBt420gyik698/EkMq33n
MMnO9MuvhV3A2/OS8tMzqfGDaL3X8ra3U3PETwhcgJy/ZgyZb36u4hI4jqXNwCca
s6F1As15hT3nz12wn2H44mqK/1iG+rjzJHDbmLkFUfkIfaviqB6EL9+ANDXEKsMb
Z7jBM01PyVkWPj47OrGu1bbhm/RW0bZXUiQokQsBZjiNc5o7l4uXvSqdwEhcExLR
uql5X0Z4trt/Tmb27qX2dt/a0pBXQYZ/4hA5I4V1iEsXsSg+3edaNOjWQlqlvbqD
UIZjO05MHVVzWNwhEG9QeYARkiJ+GVItRD+LEOponPmW8puG5rHW/7HoIcD0Um1C
wJn+I/1r7KIx5YbonC3ha6tyyp1KHfhgGGwOpPLJDxIVvBuTP30U7iF/fF60P3i4
muyG05zBgt7dWlixfMhq2S39M7PsO3B+bh+V1fXRGfj0A168wngKKc2VnJkH9i3n
AJaMlJaue/n2IaWq7KgSjUA/oyvceLRCLv1nRCQysN0hmjHjYTnWZPVfnpNarJNE
n10ZzYEtlxmOM8Nht102fg043DEPpxBO5a7Iuts3oGpyfzRUefyJKGCuPhCupayW
gHVQWt1ZvrBBGk3NPaPtnd2o8jiOCwxrLw7TED1KLAg=
`protect END_PROTECTED
