`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QzvmByLL4z4YA6XKT2mQy80M1EWiPYMkpMAt3NjCivRwQsO3dVCRpKAvd7JIlUzR
swMZX0CFIRMruxae5pCRNOPIm0pJsJOs2VNPkhZrPmLYkhSWStycXoY4G7nK+wlZ
JedMLlKHOy1MMaRrmkIqtKRVsnIz9HN3nBFs85Lu+CAEKDD1tgdMr0bK/TettwJ9
4RTS2g8EjcNJeWnPnPKtsqifydmosX8rMyBGqvkY3HLbvzNB1L/TQc+/m/kZCdO1
eSnGtx39VZWJdId0CuMrlA==
`protect END_PROTECTED
