`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgQn7A0zz5iGOSRBYKak/obdsHhqzEYVsHiCsXCfOWenpk6wTc7j4uuOATmTmlDK
sUJVx6DMq+1DtVZLD08rKPLhMCJJgvgpIPt+9rLmQcUMzJdub8Fa8BFTYX7jbk7x
YimlEE36DcLALE+wklVLVs5pwpgKlLqhcoou/ZS/LkE6OBNSLH7tEE6h2rGx1uaM
A6s/b5Zl7VrViSWILkrQbTfTKC+Jv1FvR9ITQ76qe7dXJAWeKxLgsgdHxlwSbWLk
SWl1efSsaxDKT4Q2e0mcQMcT/S21jWApkqSaW52iErsXYr/6Tgh51z35M3yhmBOl
lKZ4gxCkWYQGEV1sobCI2FofwTuCjf3bHpdO58YjnmOnA0oPZgK24I9gjgCLRtji
D0btiy7VKZv7lR1DraP5tIK5pb8afw8AmbbsYn2SMkQqGTLUOo/KnZmZBatn6jbn
LJDtFnUVpOtXQDsVYf//HTfjQntqA4FGuYPWggvrPXHG0ZZApXtzn83v0+FPYob0
`protect END_PROTECTED
