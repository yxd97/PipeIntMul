`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
clxV8XC7eSWwG+Yq+ft4g5ZoXVb+Maw8sKCwiDnbIWLpXyTKRe8wamIA7CUa0+RH
IhqkhzMadU5MOcAHGIYn7O5IYDMyrifG5gmCfk8iiOW39Gm8Knqw5DuDV6ofANET
l7bwjNKxnv18gxTyMJFDJ8gR0pC+VsDgtv1b+uBvrRO5Ie/uLCE9p+2nkx9tiAoZ
8X+LiCT0gO9hswM/p760xmu6e18vWeQwwiPt3sfVpN8PAt86E8uG91N369XthaGK
bsaPZ7Rs8I2wzKdqq/rs8gB8+vXQhFWmtDtW+suMj4a3ALj8BRLQTFwUHBDiZYH9
lkhCU1VluEsG42k6mFa+ILRjeMkTC5BvdcS+N+vx4THC6HxhOSS3zkL/UNmOeDSr
buu9k0L/9CiheKHHllhbcuv65tJdV8fR0WSA8I4GOcO8moA3lYxu9twVPoPK7cUw
SOuiAmcemBVoWK8LmWkXDVNE22SmQmj0ie5Kx6Mx1GKwJN05x/6A0UNIhiEI9GnF
mcCgaDli1bZzuPvIXxHfiYUMdz/FpVd73jTBEDzZOHG7f/CCliBGXkBR4gzBqQyz
7qn+KvXSJShf/vomGoE1Imdau52QLldbUFCE8iJzQz0fGmo/Z6fRiyIbP+b4/EA9
UIGZf2iqJF10h12d4OE7SvJTz8qGQWJMuZv4dIRmrEaWuIqhjgrAypEAyTlRWg0B
C7jqAf+vuzarZDNGZe+J8cpxXjmMZ9cw0kjVen5EljZEGyKIBQCQqsNl6Qc3U5vA
9Op1WCrju1sM7bliWk4FuSyyFGJFJ9S6l71ijDepnfOapfdwAJYqdxHCSFGPlunW
K+EZKxms3vQt5t5fg1l6JhJ92sNL8UQ1p4vdHFTSBMSY7cf8cATtZVj64QVeLuAY
1kaYuMZMYT9wA5hN09rq9ubQ3IdCF0KPCPu8C1XHOrHMu//V4FdZ01Vb2hv/nlcy
9Twu4StOc1L2i3yMopT/RIlgrDusWCrJUglUQMH+9ni3GhmEo8tayPIu02xisZSq
F7vDPdy4wMRo7QKs0SAnZ0x8d6Kepo1Gs11PpH1NM3mMwT1OAm0XNcRP4fTxRy7b
wLTDvoVqFcjXT0XYXTk3DkaTrcDOpd/d2thkQSVMk1WcIbgfieAcX7zDr6MJ443C
7aTC2/iuxp/cARdUnm3w3z5Dfio9QzddeTGjeu6/PHSWxgGcf7XcQTYcXze1ng7p
Acjo2E4CPe7+7HOB3oMMHYxh6BJ04oX+7GYyI9h468sPttptb5EJYystgZudAI0h
dor+qM0fULab4sTY7FAhzSTx+iXfrWZ6ZRJdG00J8hY68ImP9JX/IyJi9wqI/n5K
98QRKhul83wdRxEFDkQS4zuQ6y3+rchRmihCmO9UeSvaHqCmKyEd6qMcQ8aeQCVx
wa8cKCISqd+OGcfk9UgJvbaLGcPRMxPBuBvjb+cGVvQtMZS73F8wNIK/+8OX8FBM
yxK4xku/ivFGH4unt7bJmiEXmTwrF+H9kd1tlOcu+smbJel+jfD5L4YbSaogIHRa
k1wwxBRynwLq91NOmRk/SBoGHd6hf02sxU4oy3aCQsBadyGzay26mqVgxx4Bf4BQ
rfKZ1vK9U9ql0Z/ckoyd72zkO3ByspCAdLgIsLy1f+iee9zBTFsBRuPnbwuozlLc
zImvBlT4xVY9t3nJtd/Pu678qP9Ljr/4KGcuDZSR+US9ZBLSZmmtlW3ftaLHojP2
k7w1JlmsK6a74bQk3ibMTEC+gY6reSyAOOxT6T4lGUZNLmcrUq8eEfHBF56Boesl
LpkgWA7kz1e/mVoB7C8zdE3KcetMDxdn2dXzom3RWEutKgVZfQXcn0xbKGr0sD17
sD2IVGCV+ZZzbRzzONDkT+KmMUoJr7wdn3AT+/NUYBq/NaYNRp5QsiJCvqxhaJbT
vwgo5FsyMBJKtZjTlGGs6x0+N3H9MQJ4MAxz0lLYTIHDf9bhPXfbHlnh5YkvNRK8
thbVcUMC4ASQpD7HJr13M9Yov0ysoguuPEx6QCj5J/mHEKYvocXAzze+IIAvHKp1
libdWIQCrkl4j9C361KDE0I4xTiCGq6qpOyoa0EM/mWSHekDg2Z5qKRHfM/C6MsS
To0D9FgO/V20TcBzJ4tSc7Vc98MW1821WiETJhret5StkksFbX+g81OD7k7iKZZa
7MvC/9fhFpVDPZjuHFtcENvbS8sebabtyi9B84iBNq6yNzIUIg3CWyAKlUufTvld
GyTwWMphKsMd/tiDCUSTGIIUSmXf3TafRmEsnRfsVuD02xBF85iR+UfpIgXWWLKM
NgEoyXx0BKtkZ2sowEqZ12aOW7B5L+ZhCKKKyMp6sIBeY9VHYc0Uec/OGyMHLiwf
ZGXQk/HbuVEQRSv8n+DMomrIDR9a9JHISznZV8L6OgDgOFHxndWxF1cC6eVL46a1
OCPV6oZwkaysa3PJIHlUMeh2TLzPXoeLxHpPcMw7KqtdH7PLukLx82QzZgh5ImmT
i+rGaGPJxIDASY33iunAWHqYglr2plr1G9p5UxsXp71XS+nJD99FioqMLeBt0KTQ
xzhCvpkoORzFUaWovzifQEMEL2GtjX8VYQqIRufXso0kSRzGwMvI2Xl+/6d0U8lH
dEbxlYJGQyJ/fm+RvRpuBkPi3B3n1E1EJ7q0eUXsFynFXW2y5pCBSReHUSBdFmqT
cse5/ofc1hILrQHhlNfIjLoTN4tbeFSDqdiyfxLNS3s=
`protect END_PROTECTED
