`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6ic4lvWfSI39UeBgxtZXJbkJmKbau9vwyMULAmDVhb82ZTY3tNME+x2PVFQ5TT6
/VE4KUIs/wtsfDINl2eHvQw1659xGUrQzN/Vi8bM/MOzcXexg9zmB7VBOdWKX47a
4uCxxQz6/KmU4S1ovyhZNG8C2Hdfn/MMRPwhTn67VCOko1zGHOS7zY8eg8uzS/19
GtE0I6jTWQlsWiE9rpyy3ctNUnEPq0nwEF1Gcm7ufcEIIUMKuR42bgQS+Z/9o5ha
0KfZ7kQu5LuQPShgYL4NLuFGc17QmjvdAPa+aqO/206YsUjl6edzfRPtnfVv517o
Gb/8+PybyoPI15oCy/FPyLyfittjUdaI1RqA8v0tmB5l0/3JE4+RqIBmm669K7Je
RoyjkL8ILEKurncCgssJkiopSgeXAiXTuDs3nu0IMkzaidpZjLULoyeqikypOJ5E
/mU5nWRBBUKjGxWzHqi82M1HN/r77LKQA0NQWBL/AYgrygLTjogZ9HHYMEj2wNpi
SGVlOkf45s5RpFOTFwgCdcjdYyOL1vzzfgJIrvGAaNFVceVoMjazL0DcStbZPVDw
VWPCVyYXBprsFDxey3NGpUAb3yvX/LETiy9ajjp6OSe0vQjRw5Qs4VyFwnPVn4EM
GD4fDjIeZwA1E7CRA5kiWSSKyifYjZa7lGVyGmVlioBuANFF8YUIxnofoJjY4py/
AwYonUMMBVb7QRLUGxfkqpL6vB6SyLCOMYfVvSRRP5WPP6flx/+V1w3GEU3KMJ2i
huIslR8t4tjlXQarEmC0AMpDy5uJHS4ld4wvuUMtDuHi0Pu1cq0XIV7t9id6xE8N
WdZbLiyeM+fR1hIWjDGdgAGvowlf+5fHn7Qs1DdWz/6X+YhV90VI61inFECFVpZJ
RhoAgTvPtHaLoqaTp2GXIS5hTMHo6+pRCMJF9FP+HX4v9dNcl+csm5r4BvHssgHo
YJgmv7wS8RRUyT0X5u58R4QvyZbS+UHmLH1Kupih1fwpwInrI2/vZeIy+29CbAr4
lxLF4rWUqY53RErRz9yT0LnaK3YhzKsKnFEU/yuliX63SfLFEADe3KiHDTw1UMf3
Oe36bSGi7SuTdJfHCWek23deZ4NbYL+9HeUx27Mx8P/LHVkbmsVZFXBe43cFGXy4
JBHPBXNyIIsdyLxnedSOMk8yJcQyrPqzlkj0JZbrP+3I6WhBtUp7ayah9p9nxhH1
CgSc1GQfe1bzHm0+JODRdmfMLe/H7qjSnAJcc40Hr2DzDRUXhLZHWtH69S+H10IN
5u/M5OHAc+YqlphEJSgQE3PJGqtPkkhfJW1cS3pPTHgxxGX26S7+Dp8tNlFHYPvS
LwuEy1aGurjqnXW0wtIW/7+3e+esN0KHCEj466ISQoRejt/tm2t6d2TCSEiaeSrv
xTQPDeAJLp9RUwQwImLYLE3G0FKK5ayqldUvr08VXXvnPzkqtxTLXfuHRtVJn3qd
utV4uSAVDProWJTP07pp/RnINtnqXoaOwN34c+UfzxfbYf7tKtScCGIKccfa88fY
f8tPPcgs2Uqq2stFw6UtEhXiLEV8Wl8dFY4caZGNEDl4a8wj0klwifGuseT7OVG9
qBrqLhjr8qxtbfv/cisZIAl+4fX9j60UG3bUHwXIPb43e7C8yrmkEd7V/E44Upk4
TSZQLnt5gLMfkZiTFjHAkj+WjBIoiX0jPI2ANEW+rST4s0RyYXNW+8woRw4PfocI
VI/ZZAKI4LUlMDm6oPlE/h/4JHqGGSJoDuvFZQqVQZqr6XmwF8Q1Id6U0vcwhBgd
JraK0fshfkuxpA7lpaOwn84d3rSgXwKpV2eCVJ2ZN9m0CmRWt/9qxGKvCi0sJnWh
q8UrA/kkdaAbbpDoj2Ok9S5RioFxTg8ecN6e+kcsN4/wMd//NhQ/wstcKnBo0wm+
ygPBBPhW5SvUDI2ZodearAvxSDTDE079hJ5TmulXFktsN4+sc2DGrXSe2GGYp9wD
VHvDPCV9qT2NgZOhP8pMoo4djBJaiJT4DhQ6L4f7DRzO15wcWQ/M6hMUFFb23rIN
c0va/UHLnRGOq7bUJCpi7Oguk9mKnatlLxQ3WpKFkNi0VaATfnzo7q9VjSbQJuqe
7PWkN5LRf7k0p9FdWInMzEJchmaKdUAjer+TwQOpTbUApLKkMLNupiC4GHJNhBw9
PnMSPTgCiVhBQNULvSL89mfuBshI+iMBJd4WCVSnzDJMspWzBxSkS8b7waZJQ9ef
Uly81kZBZRSkjP6CME4MkCxZTwps+RKlm3tnVXybhnVuifKH17twK+xxzKdJtYHV
jZQ5dm7Ish+xAsJycpeIU05IlGLCB6YCCdcZY7fyfjCJMuelIXmt4lSGaIq3/uKs
rEU1PehDo3J3A1gW4IYQTpqdmwN/rMVhWR1e2eU028ufoBfT7PnWobSvG6c5/pMk
y6nfbMajqGQLanSGRQz/qO7dU6dDaDWW4ggI3JVXhl15fKpARYXb2RFDyLK7ybm6
siOLIf8DOAcsByz345pmbCJFf/EO6d8Hw4O0tUH1kOi9w4h66Ecot/FF3lkI1aP4
JVTVFZ9MSequL8KGNYDOGSLMnheDmzbeN3ea8XTd7+pGmTcBQ2MkPKbD2uo9hXu8
qi2R/x0sht2llrZd8FNm30CfFsYQTUPzlCZcvUgovLxRDRbuITl7zLU62JlvhBbJ
hQlc3iA/otkwUPpeCqV0TLxdfCpXRD4b55wxsUuf9W7mNmPt1WS18WGv+65lmiAC
noJgRmHxLPquuAhw0VoWAnGvhOMs1dOT6ynNgxEIIu0qkHRbXnFypW1kF+E23l5U
tvDpYUErc2P6s5fOUICmR6Y9YwAYp3RCEhlkLLWlBt7NBhKCI5W65HWwgLigCc5O
Np4PQ+y9ZzaVE6+MXXDIEwmcF6vGN8THry7WGRvynxpm0WfDCmoBK0GV7vlofEn5
N81PPGdLRKkhvXhQ4VMI/S2hQT/W3nMtgVj7QeLi/beW+zZoowZLmf5ZjMXOi7ZA
u/IrGiSTtMU55AyODKkIHwzCiNoPRkMf1HpmNkRyDnM4qWbv54/jD1/SkgARN3dp
roIsiXFqeszI79vD8Iy2ZxQKLKwRK75cV1KlnBJSOLoi0b4ayDysjk3yqux02IL4
yK1ciNOoIUu8KMXWmNCqpkB11i2W2/Uh3LFFHXihXhYYZiPcQOrX1awBP/YxehGo
fsgGGFJ39R63oa+di7+gWhbaCm7A6sciOUw0F/cgp39cuk95ylqtkJ7l8fdtuLxt
KfmTtvWPtiZtzJHvSTKStjsDMUAJpJu+UEs5MxO5iOmaT8IQwcZhwAWcr53D44YH
YI1DTJft8bAaY1shpwnWW2j7WHm9aFvXuV9bIrbibGjllA90+PxaKtCtPZsX5srb
/hCH6iSlwAsoJo5QPDKZ9Zok0juw1GQMnuE6pJY+d5mQzwkFWg0IZGl3kc7Q9WMQ
xbLJx64TJ28Q8DcXz35DJTTGLVGlXSDYppjk4cbbTZU5BSd/mQlsPEurrgxEcOly
sWgUSzdovjH9K66LnTwpBdFwoQdXhLmzmeQj2k20encm3OxjUWh7ic0KcU+nmFvP
eDETV+7Ha52MWZiXtb6ugltL+g32SZb+CLSXyFP0P9HTqJpT5FKQqsJ2hiZ8yr84
lFIabLvs8CxvZccaLWSg60pZDSWdBaUQjLAZCxCmfMKCPR8WBkBh1GB21u8ks9z9
K+cJ87pOFFruYKOvEFhPwfOJqNq/x5Izg6pnI1YfhzcTtm3wGolUL5eUBw9s2Ga8
aP9/NjttkQ3ksYEJZ87KSDAeTNpp/VDOcaw6Gxf3EIriL7TuhdhfGW+NGfvAS6mw
yyIzU9lJEZdlpi6o1N1narKzmRjlH6SNTKCI6V5g+RgLLgo1NLhs5tKn6VJXiUB2
hOn6ob8Wj3rsh4ljvkD5OxIknTkUcksEWA+meS3mwSRlPTztQ+zi3wGZaYjyfBFk
k7rTOgJcSv/0dWpBsckWLBsTia2/zrmCG/TGkQ2hDEfkBEeUgzK+MIkFoZkxCk7N
DcL69h0WDpweVr5SFu14HA5/i089foySbGqqY4mfMirHEcH9lkxK4RL7QgUh5vx+
3DTKaJlI1lnHoW8JQ3xUERGAURtvkkc3U1/ifZY5fjrf93mqfzua5Mk9uicDkt0u
PRRpK7h6WNt/90P+85dcwLJKHb6pX5wrDzNu/icVLWWjHfyp/Wus8f4eo20LOrEH
PgO8FIZef9YSY3GuZ5R9sNyqjClGGxme8tfJFo3iIwydOw9wB0KgYK7epMVgqGZW
GgRmEw9tSDTVvPChiW0yLiQf+8RS9XcZkY+mfcKItTZW79bYs6wA97V1vip5mKjW
hatCr64j5PZpZ/CT1me1V568GmbMevsEHVWdWH8fwOEXpSjRZSwz3JFc9tU7vg5z
cYuILFG3dg5MKewv9NLCcE5L0/+bTihTZWTMxmKVqr4oCkJfMj6eIaKrfneCKpiB
E6K4rp/Vmg4gzW5Mt2BHVVt92ufkSK+u/mttKlsOzfXiekLkXyPLiBUMRCQDvWF1
ufrwm8Sc8W935Tqrq+x+VARR2yhcRSJtblFhpRvGGXI8dK5aKKhTAc9pZkKNDSxk
wrzqdgIZEDmwkJ9XQgbt6KqLRpqpCScml+meFlqqYqouslVGJTd41kjXJITN7dQg
vjMH7xckQmxvI/7bqAA5o3WX47GDE7aiK0ZU+fMJxipPHXo5WvzJTGT3vdDBGAdp
p9aTiHUOVqAsrn4bwY9cJuRTCiCnxRWs6avFdyGVS6t9d0aY3zUaLbLDcIdOrsFq
S6aav/X/GPMUtX+m2ioT9av0pcLjfMET1mpoXvxOKLAl7it3I6cHBwgx2z/xl9PB
fSckx1AIL0P5txqKHNnyaD+2IXj9wfN7kvv9p+YR7BVI2LNHkc3w9evvt04Qc6Qd
jyGm0YwX4EXpo/WKLs+to+2Smi+xHT9MtgTXb/FE/Ar5E7ELQy0oaS3MQSde23Gz
lf0oa/CaBwzebFcGyC9eHMV5qcztVpluxa8Lb+hSvTvz8RBz+iMYiT5+GoNclYHG
ShlxTKQCa6wReuWa2UeJwOSzqYpp01LO/oxEOmsee1Wm5eZM/07IfMuhXF9HJmAL
kmOB4ZGqQAN0xS4GOHJknW2lqEieZC0WdwIkmDyCKRhokFvM6E76ccnY2l/7SUtc
/Maxs/dZmi2gQlStbmnK8BS2Y1A2xosJvETaopn4GiuDU+i/jot9PBtE17F0N2UT
EbrqzyEdYkk7xHhHIbzpv+zUZhYoGz2lhFCJc8FJsdq2pJxjwL20qu2MP0UBnt4J
Gpz4JmJ226Fi/uiVwRMqiBaAIvaP57aA05l1Avx+WUApJve+FjwVPTwMd2NjUS7k
i+S8H/1/jmOhHlVRFjJGMUwK65TP4398dKGuXmXN/itQvTSNQQVm1hpIE2PHNGqs
Rg0aAgn+KLaV4R9fDIVYfUxqwIDAUjOvmY9yB6mFYdkY3qaY8mca1NJymptiysAD
t1e9eBymW/pYTSQe+4a4diNNim0fNyMr3c7XEweGOJFHdN5PLVqpHcJSo70169xr
+B49uEu699fDbxnA1oQ2kGehvNxyzlkSYTcG74Xu4FN8h9wby4V5/nj/OkmVAmBa
kaQXuF/LiuRsr9dRO0gZ3mwaUb5eEmJ5wBi0waR+LGf4LW0HdDBvObgz5ODYdumU
7rnRrMbeGwodXwlbD/laSeNYsRQwjdnSnt2ZuYb5q6dOb5kqwYfBAdJxza8iAc0i
sJccFeyYqipTtrDiurRAuJpCceCpygX4+iQ8LpK4jF9Juvc3EKEfA6bpm2TrEElu
mJxvahB2J/8nYKFMewa/r55MaeweGfMyp43NQOSH/IThqaZ9lxtyq/LlBWBRDrQe
2OrZhKNF5Kw/0JbJryTEzDGvn3/N6DnS2XGK0h6HJ+2cj7oFhCVrmSw/89XwDsjM
wubciAxzpwiwXyUm7wR0gJlEPnQ+1UxijTDDS4dkN8puGK6LYCrOThmNevyIfVmf
6emUsJo4t/qIy87fI/6P54/mYPOpBbgTiKbMS7R+vwFkLDM1XgOZBjywhlJgqmi7
vffgLYiDda80Mf/9d9H7JX5sHIQFaDw8+tyZsOWSJ8g8tdNMdELQkLS2QJsIwz0r
EmZhDEhZHrqIe2hzzi3KChzDKPjC3NuGfP003hWmdnupBm/Rf++cUbO3n7E5GwRy
DDCQMdMAczmq9tg5pRrqlH8X+jVbx9e4dRaFjHuc5ZcPpuhM0U3XImBcMuEGRKdX
ocOMzTwcNeJql6KpOTFlJd/fxrLM1OX8ZpdNkOzQV3DZ+QCsx8zDJbX/e43L9EqZ
BLHVLGYGEvLT6bNuLHsh1a2X+bXcOn6sifrAMevs96YWeC5b7nspRmtSsVLbss9c
UtHJxsKilAP53oGGTrX0Lj3Je2yeLorr6oP+dRiRd5oFYel1I9sxQ116Mi+PL1Ts
4DGTDZhfN5a9L+BX5ae9nuFaK2rVEzUc9/rFE9T8X9lcI2EJt3MI5nr19SAbucgI
lVgKCotItUx68jngTXdxJ0Q9jY5/+IlAgFlRTyaB5A1Yg740OXAbOjKmppD4Mq10
paYZLxvclACOgw26sWbJxVtS/95n8A+S9oPTF/VIYnIELSQk+URrJp00SqathLMO
O4H17/dXNMZh+imbjF4aF6uiLHWJ/RL8/y9khckqMHLnWl0/prmEq3IBHKADTc3+
kNXnuKCrf4gyQ9NA+npAdRLBH4RzRsYckiH5E/5vVw9dZQNCYRjlkhFrxoTvAXd6
jgr3PfPj5g4Xmzy4dkNdL4kmH824C3pDlu4XbtN2hyHXjDJcJJ5PSyfqdG1T/xal
wZxvQPPFeZ9GzeOgdfTsH55ZxBeOdkYK0JeNxIamTrYlYjVbmYa9GUDwsGWxBDQJ
INrZR01CRFqr7pOHV5k3U3XIpTTaGO25PrB/Mhuz5OQx5de0qdYLalKeeJzNF0Df
+OsBKiej1dEOHzGtmED/3w2UGxPqXsQjDXqXjFUx5kRwx4ETFRTnzaA/MgmuPYgG
JpJ8fHXqvIa8H9bGfr+4vZ4BUPsH45iK+6AMlvrMUagPnkwsJsvuYpDkPvgW7vAK
TXCsyuvxMY5I+uZa6bJF6+sj7iFxjeQZh0vJYcsykk+c4wvUJO1Ymy8Zln1PJS3H
Z9Buj6S2PJ0bjmGOfjfIhqlMp9uygy06eZCvPJ/yD3vv5xyjy+E3WLCj/3VwDNFQ
Qq+m30tu44arEfsKLquQi9vPrnlbbXeAiq9N3QzkpMmH/NHQGsMImhv0dxG1I5So
R+n+W+G2z/P9OM81VcM4WpvYR2JeVv52kSuUSnEWDGi8bt66gkGpy9SLKlKkFC+j
zbj6GSWyTMcObyI7FN+KGu36hwD3ndOTE1jwqAF7u6DmGjCuSaCWFb2NqrRKg4bH
4K5rRgC0t0ldNNtEhHXcuHYbmBumHL+cC8YpC/JN+EKgfITrXsHT8V+3GbYlQ03u
ySdhTfivPi3zAx+sjq9qi5u/UWLuXRGHqi2ojZrGGwlbLpNpRLkIwJ4xIwma7nGF
14UJ5UkpcEsBSQmQS0UJ5ibTMg7evw5e5TnIz980ST9UF0WHYerTcpHZhNXL362e
GCtfsk67KfG1bdXUGascg4og8EoLtOmtYWkrSX0t6aKuAsT9EaWoKEaRW0xUzCcQ
YYZA4PPdMq+Kf3YSecwOz21ie7u/oUCR/26C0jC37qBJLmO7fRJ7oJ1mbjVzY8uc
5n6tUFSDp+ehG7q4U5SMpVk9iuyw70LB1pQmVjsWhsUUHxvmDB2mqsGM0Vfu+gY8
FC70k2af0Y9IKYQhrxY2KLLEY/J7SDzAVSwDIb3yodawGCJDHx2+vCiGc5YMGyLP
cKn5MyKP5Y9arxTD3iiIUcMe2QzvhhQvongL0f4BbXK6tm9WokkKgr90COHmL9UL
L68ys2bv/eaTw9iPCYvEXdVEWL8A9YsW9XQCQYaE1Hp715hT1MTNWn+LTnnbp4BH
7N5XkE8NrZXSbsuuuNPtU+nVXUahgg9G30BRuWjmUOJBZAs3b+4+lUWOj8Ibvj/L
cgmhtiEfMScp67AQZwSOltHyfDYoagUXiSgIxHW5fnsYsbATUwkV4xTDhTqk8XpF
Nx2dGizyyLIHwjj3W71htGGTlgi/KpjyOP8pPBGr5KJDJ3njkFt9+puHR9LWohJx
AWyt9kAYyuAgKZsHbWr1ChblGPWtflrwQtviQOasZhN5PJiQf1yi9NkK+k1ycN83
BtHRQHbVz1+QIlmM6KObhdcgctsvAybn2hxyMDjMX6XT0zQzxDE8OVnjSu1t93QN
c0yEFKaHI+/uS9PyxBGTqRisOwWwziJy5zMQW/D3fiYhirByWhnVUAEvrBTN3QiV
GtZBjsFNL+dG6rx5RZfBqtVxGz9vryVk9w+ULcbMcrLanZ/VAdBWBMthYVHXqorH
jGrk5fYfrVdyBtpKw13h7PX3uWFdmT9yGhnbEqThwE7Z5kNFfUjiyz3JXZY6Ytt+
pZTZR9ct7e+wRr5sPY/vds0YcPQObgfmOWhjU3SHDLmPxnPi/s3VE5gqgK9GAg4I
0LLtke29UoyapeexONWsx8GIU9mn0qob3HDEOKOGi5razI7r5eA99n0Y+agTmChH
W+dumEgWsp/wE9NixBPWR4qjOJ3Y1OJxGT79UUb3rT4xm3+TH3e+oEIoFaApcehN
SC/IDyLndZdjpdaCePbl9Ubcx0b7KAH6/UxEJlPzLaLDVxfrhqRuHt7OajwxiBtQ
cbTGGYtmmwaPJj70ELO6aPHz9TAHXAgY+5BGtZBUIv7bxOaSr+e+IZ68x568jWwh
BzIvrgOJpaM4r4aXpZeDHVSp+iPAQ82DmnmjZm80e5au3P8ayuTVYz+yqrgiZfC7
pJMnBNh3rwIILb25pT4rs7Bs8M0H8vlVB3bFhf3sNGgBziSCdSCfN50Kb/e3nNDd
MFQopVdiAnr80AXkSnERxHnGVfVjiOZYhWvgXacm1FHwTDvwu23v4oSdw7CGq2R/
hdWsai/5/U14BqA1kjXTpEKMVo8ZL5mfRwGl1tHgY/yBMWCzTFeTn1T5WqP0mbya
K1/2gYFgVSusC2zRB+3CYKkpmk+qbrZZN+j0Q3aElnrgksXXpIkz/PfmD7TTvnHL
9nq9LAVJ3q14PPWpNuJsoJW5e5+NVwmupltM17IN9oXX/zQD9fuNpfojdZFWSH4J
krfJWPDUstRISZrf3qni1Jjup8VaELLaAhdfJ+WrUcwNBi0eaEGIEB6L4x04/qPC
GyyaHEg5NQmbwmGJHqAhljMUWuC+eW+o8g6JXlZf4v646crRcAGvuA8xCrTsVK1T
gu5hHNR+yJwjg4lqmP62aRZfiw5tate++xXGJsRgOC1QxuBEeL7ZiTj1h0Y64L9M
lgeEeCo7fCIZAvMTCoo2fOcpvXB2IBRJOyy4En0HSz4XPLNNjT2rb+zHPZx+Mncf
5SueAbB1CSVML8zhzBRZlrRsVLpYIB+NnzkHOYrgUEw7rZk1KxC8D971OCYgbafe
n6ZYEu09QqqaT+XpeZef5zOecgzlDxSBQn7Y2w7z8Oia8RJClQ9HqD8/GNtcMQPl
H1Ybtr+L9jYrG+UY8oAhbRt0n6vv8t9s9+IG5HuIVwTKgmN1nzrR1FghDKW5utZ+
lfnyRxJJo0OV2qmMjAVPK0KSVdZUjFTMnlo7tNQeDRJ0rtfaLZy9uSn0aSnBWSwF
gtct3nQ+6eY/DDKiPvhktoeu3mNaVVuHWs4AWtRgeExYr6o3sCwhz8rX1F1FTw9m
/17ipFU0GIt6WWtIEgNfpNldIntAogYsKByhGX8U7/S5k77AkGIy2NzLIvnlL2qO
4jKaOMBsskbs+dNIGR1ZsG8tPiJzipU3FsSHov+1xBp/bwUCTHRBXjZVA5ITkePY
dIc752q1r3HVxydjcCpeZmTueBqjBcgJ4pqFJGAQkq5OdeKer0ofvEUg+E0eOm0Y
I/w0jZkgTduAYznD15OsP9kcxNZ9G1qgVcqgHynrUP2TWrmlk3JZDTompeWb4yj8
aKJCN64L/RCcZ0wZnPKZV0X+akVY7ud88vXFqpDQBiXeM6jF+S7Ly70R5OSulnPh
KcJvP/v/CbdK0hY9RXfdHohLovhTfWv+qEUglr5KWN83zZ3fOObHwH97SMVYQwP6
mI8YW1PJIlr0fRKfdZFhIHsNc+I8zy5aRo1a/Y/q0DCwt26EgjKVKWPYGgzzxBfQ
jt6BHdLMlYFHSgPji+qwLkD13wu8nIRXGMdR1aoisQ1ckDyU3rvZBEipYENPHKCO
NBEyof6GBRntWXUtFMriuJeWH3irEYqDTQ7ThjwMjXR/mhy1niNFYEsUaS86FYFq
1sY5X38BkqTTRV30kRYYPB5aBCkeltwIM8d36aPZTZzzywLweOfYHp0dK9mCeYas
JpDDlmZJabXw6o3lMiFs9Dtc1QkPW78uDktqIzhrOjeyDWYy2zYLD+ceZ30zc5g4
NUtS9CAgVCyWLD+eCos3IU1iuWF3kKdibY3SkuFuU5Xt5JTAc0k8Rt4vVQsYMrG8
bOm3yE/36K4y+VBQ8b8Bpwms5qMkb5usEJ3SAhitTiWhOTU3KQhgzUMtR46wwRHG
VLXguO68OEwIEmYCuKfX5NMD2As1FbI5FsAp2J7cSWyEyv4VJdIUcU8PGm9cVjsl
NYrhop1WIE+fMAgStyYQy9FIl+ua/4HVwJjvoYlJSPMdTe2YNvVXJmQPBB4t44Ho
ZGczEkQ6eAOO0MhAL+On24WABql3QNJUsTKgcC++P8ijegsZ6sq+3qiamoh0515p
3Jmgz8VJ1vYSaM8oosTdz1d67gOEuGV4UsCTDthp50pAltH6JifqgFW4eEH5bOSB
XMpL4oZjaeRZCkmVwL4oFuQ3Qgu+ncjm8vIxdqFoNgD+3hBVvmU5jSxyOXXn8x+8
wUUlrddIsI8oRfh3FESjXst8gpZ7r2hSCcqxiut/2HBYTt0bTaSza2wdQL55Bvs/
Fd7tMbzfefqsxtbqs4jjMn0QrxzlXbdbihY/m/W6oMP0AnzIQZcN+gO3+TMqg03w
oZyuicOl1JRyJ151i1RYf45dmt69nipqEeJaUVQWPRza37FOq0YG/lN/i9QlDZwT
/EwkacGqZzvFPLDrr7HHtbM3yPH2RhxHMg6djXAYWopUVHVavzx5sN/yG2wZWHW4
1XYZOELQ0gfwhMGE6MQviImeVqJhGmGmFzW8cGPWoiqG+m7qBP8kdJ7wv8ISFJt7
RXuQLd79mFV7dahwejCkxy/k3lMXNUVKa2rEH9XEO8ooPfuaTfI3Lqd+OJ0qhVrn
Zh60c7BDomZwwNIPMkx7RdKcYMdCn9jcufJtiKTExnRw2JSFrnnArzLVB0ufvcxJ
sI8CAT3Xp0/au6lygJG8SQzDxD8//6aFkXjBQA7oY383eqiV381IOGqeqj89W49K
wGxF9SCiXY0PQysrqLtUhIp0uRIlPcWymhI7bH7RavpKRQtaK7FCB7u7wxptrGkE
oLwOQBXOISzqwFl1dhzIUSzYqiJNrZ2eedux+BhE4qNRhtzKIH4JPuVeUwEkSr3W
rtdB4JSnhVyYx9pKmWubGfxV01uZ0gmOoLLyYznM0JoSryXq7SYRuGSGF7XibkQD
V0VJkUE5aFvHEaZ9h5LgL1iUGFGN09T/KoK6q0D1UPEF4gFd/Xhmu4m6odRgO9Jt
Az42aOW68Y6JEhADGReUZIO6WniFuhtqbissv0Td+i5OhrZaaCTyvC5oOka+wlbS
sR/6asvr+4ydXcVfYtlFfIyhjYk2tdLTkGzXEA9ibGVKHMm9E7vbUIo5ppNtCt3S
9s24KcnuuksMCX4zn1ZgwQ/apo0P9kJTVff+CgUYKUCCQZuVxlWKGOtuKK97s9er
Z/RX/qclm7SCSAdOs4oAIHqGcLoU6bchK/a5vAku9k7+99EusE+tASsMAmJqokCa
kM1VeSq6gGuApwwIVF55rhHuipJ1gzlDZhXPcoNEgCQ6AXqz8tp3M59PfRhXA8vQ
SLcFpMALYBhAJbXHGD5uteRkwhYvv/MN+ndxAV9Hytg7T4mYVuIjuBWb0D9UrYrQ
Is83T7euE6qlMR5qADrJNpwLj3UH6st9QmuGO1zBM3oTPkKVavEywer5MONwZa95
8lXj/MPaxv7SX2Jies9aX5m5Vp3eVVBb6w414nzOh6l2ONHBdYFyR5Ou4K2h+1TW
Ua272mbD0voH3DpBeYri1vqAb0pZhLbqGzMk4l+gJCWG0Gx7MeFypYaaKX1F/cgB
+BuyQsitvLFJr6KzQ9rr0ilsMmNb9plEzKCHd+Y049XX5ydzYFJ9IdaylMWIE4vq
MtUxxCk4LVxqUOoGz3ZIV43jHVA5tSdavUsz9EbAIaIkTpO/IxYBDslwysT4hdXe
BqtpYEkH80psTLB8zg5jCn8wEBA7aD6acLvYUpKiaW2olIHkgfmYd22iszBjWlqQ
wqLQH7oX5Nt26r7ziY0RuVKl+/khziKVK59Xf0/puGuIwJG69j4abExziFQUI2tn
KkwPpF3RK2p20WMVxhEfuSqbvmnjudr1nY4i3Wp1CQbLiyIXTnDaGY8l66u9Q+hQ
jnjbjox4kDhHFPvIgRag4YxrXLUJQ20L/EdkWDTnYFda+K5oxqKIAXXBtasDEp6r
HPKpy9gjxqItjgZNkAPWDOQSui0beLMkoqNVr0+hiInx06CbAHz7Z6xxRTRM7IGx
bn3xnM9IV7k/stAJ9U0qwGJxP+Te2p+PcUgTEs8OdebVCL9ZSWZccmdHX0drtRxR
QORNJbXsZyOFWsT3mp0RIs170z6srKGG8MZVnR7wxeFiZARzuG1OswHhcc6rxOAK
DSz4PNrMRusKHjyOxB+IT9JGqHLrhsO8w4cnGIH0bRaKZ5YRLl9aqpamm2An6Jth
2NyIcWGgiR4GFUIm4n4DIoJenIC2scnnK38N5AzJR7QifogyMsjNY1ENMJkatf3p
CfMxfrG2pLyl1iSUB+I6eTmJPILOGlib6nSGUT2xke/1pVJuhkZgP4/ULMASnV6V
uw/Qhh8aySIjA8SZsBWK0cqdEOc9L77NWEOplCnyNzS2iNhGsVsM+n/4dAUtH91p
3u/hxIkS1+H8QkESqO8GLwG3WSj+YzEJyumNIMVMXfwkJHwBLcPqBpxjxDppZT1q
cDeWwZFADRcXol/LCDkO+hUfDQRp7TwEI7HGIsKVGX3h6Tq3IPilo0mXCQL5Uqpr
TQFM1TrvMfh2CYOpLg00O+1H9h3px28m+rHQy2D/12aL1vbM9cNnwn04OXY7iuEV
gvWJxADVd3B08X5SWTfutLsaHBLvwwj2Jfs8RW0zgnV05FXCS9MlMSDljoiTMwES
Pj1XxhHeZJB2kvFdllcGevdgiGRT9ut/RzOHQnvRjNLrPP+EOiuk9S9rtk155VVy
4GvdHnj8FW1nf+iJgfQRkB1Rdsb9CqQZctwx7i85EVkxyRBtIM6U/gWtj1JX8saA
IAHIS55fXAIPOTPksKIrQGsNm+/8sjdwqh69kE13TVSmLYmDlae0YoSwd3qQDCeV
qfeMtShZyJ8oV2aXE6YaIpQH3P9oB2ZTTnMnIDn89Ck2wWWHLw0DjICkocMJL0qH
OD0Mjr8JqwrayMIagRnfN+g1Q1OBL0dhdC+DrI+30w5myn8JjCtDDr9qbyCG2DJu
8ECJxy2k1Z4AvrbQ7LHSJ571FiZ4BzlAgkV07OYy1F4XJqLJrwpEtlvycCqS+qEd
hAISZQ+ESn5vW2W0FDy5d26G8Ja6XPpXPbzjNIDZR9S3+HxVvmK1tJ7DOvLjjC9J
SkvrES97y6fgyMKJIXaib0VTGyQTODeeGBc5tUVH/AxyAJpkpGZn7gl6BaAVfL5U
PLNKmgtCMoKeQcoEYjUS0QIAp+mwrn8w4SGqX1rT6Bo/BMluSihRnSs/hh4nVmuz
xnyrt7y03/EK8SbgSZpvChJUx9ksWbcMudpI6mv4Mcqd/uII/l5arSfWblDKvMOY
hUI7RlIob4HSM7QPSUyuuTRVJkKMeUCoOD0PtftV5D6CIJBk9PvPDSU2mw07jRUE
fZ3AvmNYRmzcLzsKYjkf5qas/XOWw5EglWeep+iYxpenV9PVQmrKUv3xVzaoHMyY
sOZTtRQMz8kWtTU1lzkZTusNu4R2tAU3M1zUo39q0Hia3vKd57bxFrh3UhftxJCC
66cNM0Ifa9SnLBGvSFnNpOzVjEAlVW4po0tPfXUv3VDFVixcNlStxeQEpyGNubDy
pwrrGwiTUjrPFZEeM82oLVLyPFD0n6Xo47Bls+rdRjjNkX9axgowzucHGUf1rNvm
O//JjwwTkbOz7Z2Gs/o+x0oZESWGrsgLfkZ0bo5blxlbYVfNaTLFzBYT6RwoqSnM
2rdhu78W8gLHte+bAGAyM6SxYmdtuvfny8vLGxos72A7L+3KNxo/SSdF87YLzpip
98pQeIv0Ih0qllz+cpzU0kYnoTVSEaTqdnYaW+CTEYSJjc1PGscdyHSzsmHE3RhM
5wB5m8KD8+YQ8rSRAx4yw3pz+X/3fmsc+fO2Bs5LwGUqDlGxlCNDU8B5m7yidwpu
cXirLLpJ41IirclIvwJ0H1bnqfda4qFp5vX7wt3M5jwUXQXhunN6Y/B05ksZcyR4
w+2033rXJms6Mg0rRhEtf3Qx72COfmXaZxYBF4mrz9OsrFPKIttsd2uqX1pdFSjk
64zpvnaGg4bYnZfUY/CtTFkzBvqhaJc0p2lrxTbBtD7kmX/QZ2nrUvh3fAzU0h7a
Uy8Pm/hSzsPbt7voODwNEpVuM/Sl8Sfg2whrCUbDiR5H6Cd0d9Dbenl/m4R/Ljco
1JVf2vg6qUjegiRGluThtkAWd4+Zau1xjS/a0FzFtykMYN50lfYhKZioYIz+k2dF
fQeWHPg1xpdfZ9xD9DHp6LdKMIhtOyFLzWpQbDsgzioaQLmigWBbgXZ/DJgs/Fq2
ZVjBfJsR8Og3Obp9DKyPcTkUG7mbTWN+xWXKb6C4uZ2G3uI+QUsGurU5G9e5rP4z
qV/89G51v2vbI+dcL+/WwUXDFz6NISzrPxd9L/oYxGLRMLbtR4G11OoVt8JOqz+u
2YpYMWFnV4ebJV7uE9vt3+6iQqYkewRBcRS03oHDbXUq+FjFD4ullRVdQq8AsWOs
WOiC0GnSEOom7lb0HjatL8WLwoe0MoK8vMB8OwpkINgUSz9UwfhHXdpD62yf1kbl
sGO4H3WqwgI3FTkTNWcSKNf16iaISptuMxZfZ4kyDcvJJxYeShR9JNYSrddhTuDb
CgnQbCc3ApNnaxGFtOlHYESdUSEVHkHPg4wMqvApZ7+Hj2S+0JsOaGQXCmXyMFOt
Ohk4nLj6teHBaohfbcUkZwA1t/SV8PCCTd1i5s0N1ahwzCvwKArTy/5egGNxzKPV
e6vzwFFa5vUqYNzEy1AzQKALOlO3t6b+8yhllxjnBGSNQktW5Kt2yd23jM9eSdmZ
GA4Hj9Icc9bN2E4sqlf4W7eLDb50FwVOs+01roRcH/JTaHYSVfaYzviM13pWPSgF
VJGjULYLh5my6TNB5g6J9PLwluyzVu4fo+j78Tp7UX818HpFSNY0+B9cICbQv0OA
CBuK3GC0pBeVBeTafi+lONQdn/R74woC/GYfmOvT/nx0voVDXxEDNCMlU+fCNMUB
eEcZOkZcv6KUCUSK03MiayPEoRxYOJIZaU2pxoHP29fLMkejDsWoie7cvglrq/cP
BZzmF4MMxJ9P1Ulpe3K1e6C3ptGj6/T0V0awmsQ+9PIV9/lOmfhDWnfyVPDkf+E9
oiM4E0EKknHqSCcpN5xR71nMEYbSr9g5RoCmwyQeWrCAAAokGUbZKrK145JVRuG1
7l6FBcz8Mt6kivBJF6lpTzHtzeeyGMtag0ygginzzbCK2HGtYQs0rWauS0iWK4Mr
oaVU6jnHWPaUzwY8fhXZbBZ0p0BlAce2mNk6/t51yzVzeSG6txgjkr/g/QdjGAoG
mmF/lhhT7n0lpbdK3jPFPYHHFtv+OlWFTEtVwaGNvfXrqVRx7gFugWBcTo7hxECu
m1ETpNXKMF3SmPRzRmAddI+D5MGDROjmhOJCct6IGfzsXHjRTvoPwXVK41tJfVek
/RFeAM63c2NqkMJSHZq5zZfx4LQLlin6AYVB+pYy52+2pZ0Y0GsIBa2dBZDqRasT
IHbxYwDZUKsC+wqtznUjTjxMG0dRI163Ud+AcCNsp2TImqrZOsXQ1Soe+ODikNUs
qypmP9l466T/DjgA7jf0txwqNNqRvr1ywHP7gifYbvuj4962IhWiCvtBeeBvcYlf
dbJCRlAOGb6UYksCkn32kiJE+Ai7kipO2bENN6o2eL1CrzWEEFYs4mipt8PoES/m
YiDVLfFW5xF2Kz14mS0qNO+oyeo992qQFdGucOzwRFBp6arfUNSAfIIrOUT2pDQ3
GuhJc5vKV2yVSn68cF3Cvi9X6vjU/lH/U0xmmbKoX03dbnqzE5v05bMrI9SundRV
GmasdqxrOIjUbbJgxcCAWRCWFfRlnR2+FhTuPPp1KzgiTK1L1GhX0c5IEHSUhF4l
XKVkJc2Q3duFQzGXEP0ydtg2vbv8LxGBT5mD217HnRrMXfT49qXTzlO/AtYnopcj
B6/LEn28QwuX2ZIRzb/gWtsOEOcnV06bWOLAS1rx0wzXpozH1cwPK7In2VbtQ4K8
SyprJqmeZS6iwBBa937o/AZMyhfnpInBGY4220Z163sir058V9SYyUEID8jwgmLc
sU0em8Rj3dhOyfNZXjEdn93b+/EBXxUywJGviHLOww0I4vasktuLrjNqNWDv0dl/
PTBGF6WmJgBaOi81hwSOeax4Tn9IFMKIWJNfkMZytTKLp8Y6tsKZudCylRjgXL7s
2U2/62rionUp8Otgnlrj75Onlxxq7hgxbfLpUKRP5UA8TZfoFJzjlmxO8QpwUDaK
S1cuG41lCGRFaWx5HRRuQEQaUfO9UyxPsU7c3DXw7niB11Yq3MlAzar3evh7wMPp
AjYCyo7uvoVZA6+ekgoTjQ3TMc7E1y5d9agjyJsE7UrYgN5oFrFSzgTfPdmc6ixR
bHuxboLbcrRwc0y99zaG1JHrGq9nH6yBSnexOZQekWtdpt+pSjR5Zq8ODaTJ2zra
2DCMo0IflGtDk2rGTg0aJOdyV2ArWudQuVHUNa/i+x1/BH0yuZdL7HqinOreGlhM
8uu8YBSoLKTsUUnn68ywEHvhHhug5FqNicagdzfN95VKPL5Z3cFDqHBDW+TPaADl
nNyxJLqHHhdBrmmCGjlm+vjIPQ92IxBpR9bev3J3iVm6+hVxbTWnpCUQ5igZ/4jw
rxvDKuliwa6HLA0Nr5npVRwJNgt1EDBpZPATOwlOcp02M/6vJFSbLdsJkhoQBh4w
DMSlNJH5ClxK7Mfu8ppPwl/XIQF/g/je3TgxBrnNLcXSlWDmqMYravj03IXbHrcx
wQEj4Ip1aWWfUW4x6yOV0Bjpi+XnqdOM/RMD2xx8k0Rfi1yZz/viSnVvGF59t/d7
G7GH9OtAMhVh82x39wrZhaO2DLP6jeXNaYideIQqpsk4vdYjp8YVLTgAatzGfDSc
oQEtg0kPXxGeP2QbaWFBqCRSZGZEeTsMKhLSJ2IrDSyU8cNuafHslhsGGfpOq+Pr
ND723K0sJ5zC5VaiWRhcO/5Cegq2pZOQ35OhcfZ0se6mqlkIqcupiHvmO28rWyzy
YwIYq7L7SDMZxNWdb5hGjSMbh9TP03YduN9zP/qFYyMcGk+0XXnuPJtrNzSFJL8U
KCsckYcIkyOhQy56UOxUytFYu5noQ/tmPfPngCNRCVi3IJIXi1RAsRSrm8x41B2F
WdUxC97yWJ9C/LOfmxSPd5LInZYdCgbnymthzKF4ZUlR2ztNN8kiFjWhvBbzVpZh
Si+/vxquMThU0TNlWnioTUrrS840wEcD4BqfovwpyJ7U1kfJR5SbfzGO/DoUWPTx
zEVSZqzZ4ced8Ji07VhCZcjBOqcTQi47fzAy4gYrXaVoKhbnV9oPGs9ClkP591yx
MFnz4oSps7Xk2ojMApYCMH5Ellk13xAgEQVR5KuriUg/2mRSUM8Q/dH8tdzs7aqN
9OcKawhdqNij38ZVUfgbKVsPBQ3+rs+c9xp2f2nELUYnLp/iGAKb/bx1c/QCm6r7
D5AvdrKyAJ7erwfnLwZ4xhyw/XX1kIiqdWR5i/cX/56zYIIKr6GlKgf1XOk23L1V
F4gq94TFr9x+lKGIvC5obdsznpjPWGiWXKOdcGW0SUhKUkHYOrQY6pTfKCOMdC0F
c1lvXWA3IOYmfpa5UAo+mIyevz9y7QrnffNisfViw4qp+xdRqX/62QMEdxG48/QO
D1tY0DHid1+Wr3S9HgdnZhu60SxxvNYjxZg6WZzIr6FO84bs39vavcmYLop8cHno
UhVscGcg0vgs4bbjbe8OUteNfjJsWTcg5829JbLaDxu7ArDFrhArgtGPIevuY9yG
4ZEUBWQZTBDSTvbvx1ZCozhNbK8BgA2G/T66boUYLz1WHpsv1GyaoEmjxlnXnJ4h
GNzjJ1N3scNmQ+Poaq5NLI2DH4OF9tlUHZiNyUA4C628D88SPL/k2A6KER1Hqpbt
CNHUcPrQnVPEGKtNDf57bCQxC3CBNRv/srpGChg1xR3VqPc1xU7f+PVdHCUqr1RE
zdTnEfuj7NBfxegsvIXu7UNey4/+VVXz57IxY1XOtG0nArzsyt6DF2sPAucaaSxE
q2deuXlpHdKiM67Zpmk/WPS2HYb0/3ii2bRCnCx5Hhpq9Nv0kQK8j1icyLh/B27B
8Ob+uIDZ+cAZcU6kS4SWU49d+6jVHfxwfmfDQoOpKt5LmmSalm0Ru0F1Gb3t8fJH
4/s27HrF/ekECz/fCnelf32DTAr22T2hZIaQ/PjWEiA3EFt5nRd5/qOXXdRulQ0b
806GKGuYWw0+ThWbZ/JmZCSABtJJ8W+qIX7cQf98h6qWOsr96YCHc+KlVjLPvYHU
0lNL7+mGr2XWNfYRU5riSWw7PtBbVCm1eU40FcZDYQz4BbJYbFQ2GAQAjtkUwRD7
D8Gyw/b2nVko54HD4hHDouDK8jisoOBN0wfVnnaPqRXyGX738kU0/qWq+YFW9wPg
gZfpKrOBCs3Z05c19+BU9urlR7oG/hSGtlJXY7YGXxdzaImZzDF/3gPSf17Y4Ah5
wS9lGjeK0aLO9uEfaklIExeDOFjHQaIA3AagMw9DJJ/wamhF5doJ5y93RcGZdSKk
otpp8yEdrflSiSY6fhODDjtiBNdtxSA5LtJb0aRvB36jd9m/1jF5dIr8eoodghGA
5DAp0aYMux4E6IEpsgK8e5EVfFO8KSCU0fxwmlFy0fHS9cyGNFvpBMxcvuVyY9Fd
3l/bOZAW03rkHl/comHt/2A6Y5mRSeGGaSGkUGio17eSlLM6AEn0uq2/bwzydtaH
Gd4hDmEq7E19AbceDPyoyNPgk2DKe+mLzx8unEhJrzTjln2YE2hN+pBCvLMDzmt0
u2LqH45zTGYrbpTagFgAvImPCaokNoTmbjtyT2yTMGUzFtdenN0eCqTbfLgZsr27
QNZsWxx8ks+4iAj+HyeNTWT9IIcSJL+WfqVnCB5obW/dbKtes2w+onxvA/ljlnrp
tMhLJf73a3L0xZTeCzjS80A268khGew/gpnwwow1Ql2Y03Zc7+ZJb8SNk7ZXCECz
Al86Jx5gQL9tvoPOylFbsa1UurEQF+SF5r1/KvLtcHRlKwi77BkclSk9ms6Rhb55
opwo2PcMXAp2yLWqNdUjAp5rfT2rgze1/DVxM08CA1RfGvALd4Rh/auIyfA66mtY
q5HjeNRHxQVBbEjxcv4GAZD0E8WQ6VEwahGe/DPZF34/yOr0zKnxflhdaiczbtsS
tikFvvmu/VANeXb5Ves4JMz1MFAbNckgSHQebn4aNfkxQwVHcvCBNn20s9XRwFWP
OUbDneefcA0pZqNGICDLT8q4HMFJh7aHB155/4+c+vmifhYhcY/x8LBzMFQoEiHc
egkXAazboQWqbO2As8F9Awnfo6BmByC+WDRD2F+BMgQViqkduConjpdbs+IcZwil
9NXYftpMLKwXdAV365TgVvL7KIsQRgxulJ1+egCUr85g/ggqmWv2EaHW7dTd5Znv
0JbXXkwIoWILH2n6gFkZWOvkycyIXpkJgkbGrf7EH/BASMko5kLtvQdtDD3NXwOi
kaIfOKJrvkU7FCuf65ySMvsPJRiz+HqcoEHYis2VSmmJ5jI49fARjPKJcCBepQtw
kC6fNvDwe150tEhzx2FeOBhwJ/sWT02haF/wTdiITLh4VH4I/QCuI/Prw+59KyEV
ojEyG2PEAnJ1+mTfrIXEZi8D3OK13TJHu7UOXxcKObW65ViwLTCRf1+qzpl8Gyc7
ovkVlUHSH/ICsnCklbTOgqtPG9DFC13HWCyX4PyDg8fyX8Dm+ePEOe2RIS6xnB7D
Cil7sWMbdLYP4QgPas3/32eMo7U3y2LhHfLSmWVBE+P6X06RGnCqXkGz6cztTTCS
jm9hyjiSa+zxZP1dvgTeIlFl4yxHq0hSAzdPbeAMx16CX81biIxXXalsUQ7GXOjQ
7/3fhGOUQqtg1DahoeWJo/Lby8wAkv8orNPRWzOJIEPWbbvWZ9ubkRR6I184cN94
nqSzPBexITLZGpXUux54cUYEfqre9ewdCErrrcp2BjGM5aqeixMEfCtE9pSIIzGW
iaelN28jOll/uYxDMFL6TtiEV/Nv/B14HpulucN3R2DkcW6Q8/2Rw3N6K56hbOCJ
BWoy6nU2eIzttcrATtHhnvqYb6AuJpbmsW2EyfvRkyvtOaz/4kyM84Sppchnrpe7
lIFLLtansC/H39EtZU1KA/KJsdD7IkztqdFzG7QhXVwnela9xgybexD3mnT3A+bL
mhanA+RxoI6XGwu7IcsMkA3F0DRWaUutzhcq28AyziHVVBZ8zRTxflNP89/kS3Cx
eCJDKOXySZQAVCz9qWSaoj8ZUI+MhClo6DIL1gYSBJetark2uIg0Q4SPKQDoRfjN
PF9OI6R+F8rNUj+SP2rvo6BqJPRyf4kHr/MHakyXPqngdjtogFwmSKEWh/vfbf28
nQZ7W4fkiGRXnoJedtf4k5FeMnsil0/ZYOTepwAT2pBxxvFoh2LilbgYtMQrmxbP
4xnoWR/DmxBLcXVu/CvZumUAxtKL2u9rmrKxK55ChjCdOe5CikVXn+FnYZafL66+
90LDKPd+kyjPXkcTq0n2AYMgK9bjm+jqjOYPzupt4epHm7BS+J9jEjJGSr1sPMSi
EAgmR5QT2GxONVabrnaajZXJJTNIJS4DOCKGq/l9R9SNarINHGnSVekJGIziXgOA
7aA/eG6eGdwyuyZDnM0W5HrkugitvNsHAXoJj0EAGQOvQ+ZAo6eMmQpUgbuMhId5
fYPrrqSjEJfQfOxGWg+SL2+0lCy1Sck8tYnUHJbKgwOHTgsNDyhSAWvshU2Zx3fn
u5bFaQvDyjZTx7XkLxGuXGzEhMQjumXeuYS8zIg35gfNU5yksHnFqP/+IPZkOzz5
ssJFmfABFevRNdPTcCXRvFvhZJnnFmrXcKSaqZzfPxDac9+1GgKxR7Tl3RVAqrWz
6gBqyASotuu34m0fHf/FIdEU+RDOC0k12hqqNWKS0B2g+TjL+ATCTseJZELErHoF
TfA2AqqEB7m03ECwWBVqxvSb5m6BkqqTx5fb8tfzIlnRmGOGT5Q+bVAOQc0wUo6E
2hdo5yYg1geniaRQgl/bfPes0L3pCavfkV/iBlLXqYJgBmOF0At/JhWnLnI6jBJ8
ct8Vdiv65AByW8wMYkfaPHu5zk23R1ZnH7hAMwaTCIMfANA56qMMnDW01EXCQ2wN
wLypHFTN6/cMs8GAIVYuAX5mbkL6Nw1wIDTJNEtuxLjK/bELIOeNQBgwY6QJs4gZ
WbQqF6JmWTtHdpfRoBSUk6pKo4WdHHHjjUFX9lSmXpY3zJVuMd6+t4BnqvCiQ8mr
j+gV+SNHuoJyO6tLbtLOax6FMCJSTbSkxHScek0pKGQiI9TigLL3Frv9exuE4jsb
j4TV1tplkWjVwlb/TcAHy5BYvJwDWRGYRn4KHwAyl7I0i2unQnHqWeFO6msSKG4S
nisC65OwmVq3kteQbxuLNnkSEKwUiFODXEYNCZju3fYBoBmNNteAT3MD5iBtbivA
qPwPLSr/mTFj7am1fKaREe1W2ZI6MlNrQJPr3HO6sbQQX34XuSsqTJmUBpvPczVp
LJZYERb6gNwwyG4Macg59/iRuo86Q7Q5iEF3VIk27WLDqC+ND3Bfv0u9yClZuEfB
6efYeQHt+7Zcy4a9h7GoR4OPCNSs+WT6/unhy1eFpgNzLom1bqv2wHvp6xJWIWjI
lmSi2aKCUKNudE/nVk1XDEkJxBSOHotlRNBb6peyISaLpp5FkVqcES3tHXWGgNgM
Zc4z8BbkJEjabLMhd/JCD0XQboTtzGUNI4B5WvKlp8ukJ7rrpxTPZ7ctc+yPzLig
5eLlGdr+5e3TETqy6auoy66X2FKKYSbFmgSsWMrsAHgDlm39iyJi5J5iZCkYn4eA
ELOhGCp6/FJldmCfLevjOzUX4stmIraB33yCygp7OQ75tKFqpCtvqtikCW4PJGvC
uaJB4CYqeyIqG+QoZWt0FMuoTbekEg0Dkx0Tj1yjXUeLKJcPibFW6bJp9aOJMwWu
o9c7veoAllhRO2QvtnC7EMhwf/6t1LWBZHJui0/C7XqwY2DfIbgqfZquj88wnXRu
mwMCmHhoJ2iaLR+t/J+oqnw3pPX64lsX8oAkfm58VdCTIjrN8Lps+obrMCQyym6v
UthMmcPqAWymnvumvXwXu3ewYVR4bre850MJfpEEyGuRPWKBtUSEH78kPgEDHuA5
dO7TzRsPWZx3ZB09Qc07eI3Gzh3AEWsxl8+B5ehb9Px7ThozIuobp5ZzA90Zfoqt
AA0+SpsgYHbpKUtenAMD3reyFqhD1qw8kiNv6BDQUGLj5JQY0oNkG4fq26YI3B9O
F+1zvrOvrdeZdSAFOz8tGr0ZVQpn0knsKyT0pulKY9M41YBLA9izbsAXidmhxV4/
NTU/yrY1Eg1xskR7WlTmicHjDzYpcE0OUj29cIZyv3uLYPxp/0jESHinSxqLhydK
FmV5EpJAJ76IQljiK0fonY5dhaZvG0Sua0f6hLjLvjh8A39pJl+ll8nmiOzkBPeV
vGGG+SObxDgRtVfsl/C0b8781yUP7v4vAt6LXyjKBobp8RYDN2KF0cd9WeSYLcB3
80eWG57liMA6Onc1536+WRzGatx5lv/ri7EKuCU/vF+mDcqfRQEhU0sP1hSINgew
xqAgwMQ/Xm8qxAA2SDS1pGLMTyBZc+nb1S00MN2hjD+TlUy14U0Bi/MaVNp3K88S
LAHtExSkNfAsF7IuVxRhVWPwtiTsCIv531gg8GckB8D2aXXen3DHyTfhis5gGAzC
HR9FYzekHJGmUOFYWulKjhyYjXDJEwAEkx0O9u2AZybLPkaz0KTu0/xJccFVEuMf
En6Jr0DT4o/E65BfKJkjh+FpahdNQZej3kM7ie0eYD96cdKZy8gxt9s/9BiEv24v
n1qMv+/VEY/q4UX+Lwnvsc1CPBF57Kla9K/8Ms5Hu1PAtCcFH5eCnC2W++ttjvLB
Dix9sXQt3WI0N+0M/RyMfdJkDrrerxO3StgUzkxLdxspxAelQ3FgsAVLn1hLOppV
ALbaWen0ax7CHdNecMJ0hkpmYvaZcI6DjxpRzliRK/z/8Cweu909vimRQf1uERq7
Io//LpjBgsRnVHxHwdPky4EaO/TnQ+EBnXNYpyUtvRoBoYTi8OxaclQlbCsjqAT/
yqxCHvw/TJNGT+ne0z04RiEGkL6rDo99FfTfMkQsiwPcT5SQ6YjPODqaHLl2eCtS
ewQzeh2Umy+lwnwiIWa5+Ll991Z5gfi0zggUpGm6RK96WxT3yQ/Vk8zDWpHkMisc
nPUnF7aUd4mxK3WJHIUvGQjNGmJNWdhC/pW2pY0QPsri+V+a3wXA4Bkx3nnAmibc
O7+p431K1QKRamvDigRVilX1E6DCTcYmWN7Md7G2sSGmtQruDM2S3l2dvTdnptGS
iRvst1mtWnBz2hpHvnO8hQCTyvtcL/K9ANM2WUCxueAJvEYr+W6KuCYXEanVuJxX
Hu6cU0ehWHMLv6++zxtyXJCgwTGekGM0GNn41qbJtDzbNsMmftvRkoAZjJAXpzvn
umLnJy85Ri8ouHuWYshM+D6p+lisNY5yoSytqrq8lB9FSIO111YXz2cYXBsl20/L
iLv5QN2paUY4BRhb3Q7h08o5zK5xi1QHB0JLL7nhWFbWmHK5QzlkBbUdS67kWTNu
8KJm1yvJH8a8dy8NFqcG2+bZBwtnCRzC3seyGYP55gvu3nEf7Q3CJAs7KWRyyjFz
MMHXnZZe9Qriqc2jm+mTW8csxLNyoEGeKbNLouBmTSKVvpOFOHahobEAu/i2a2S9
32yGYaYQ37WUqBjGulMa+DWvDnrC7PAbUqAWG+3LR/nkTypWL4MkH1Sv/Dcm1ozV
Mtf9sMfsZaIG+59iXgKWeDc6yLT5LWGAazB1NYzq0mFcJwRpC8t+91TK2EFDG9TL
MARWXNoUo8gmvFk8D/cQ1ri+Q3IKphC6mqPxhMNp95UzKdl0+BBq+6BXZrIQ/xF0
ipfyXoeR2+GrzIEKId2mCg+7L7SnC0ML2ptTW+UhvatStjUAJNonZQThyh5rjDns
apvfFyOkUAwY/a2WBZ8/CpM8d5qGjRCObWTTXF8Edagz84WsM/ItlFEMm+T7mvML
TKRO0oh59a0IzJllBYqsEpEhz8GiM01H6L7vZ4V3TWr7QTAoxEk2gRxgdbwaXt83
KIT/pey9fZj7NmvYqCTZWXuaf6/7YimZMuWKdznrDJ68xfTkrX1MC5ee6hCQpVB/
i2WTzNvAIzTM233ngEg2tLh8Uv/uzFiUP8k/xFTETH4Wn0PYfmMVCxTo59aq8Qn9
hJT8SjUe9mlekcvz055BZV1tD9gOPoHt0L0J32IE4Wi3sSVMUzlvxVuULOFJxYDe
XaVYzUo6fqpUdScGnpxXhHysY5YcRJtytLOzwpueVjgMXWhKju3usCcsvzGIz4iW
yheEQy7s9Ep8ae3RZt3wkO1c3pkwldB5L5qkqbhQKE7MKum09c4vYl8uWFIyLXWD
qkQfR84f2cUI1CCr8P2FpvoeOB6xIuh8abQ2nD2oDL2xNhvhhmIOHnu32cOXbvj7
oiuhNlhy5xwazXR2ytPKizH6ey9kHZVzajivK6eIR/jEe9r5IS8t5DFdP0Zt029Y
amfHSRtCMbKAZjJHuECxmLxzd3NAP8zhz7Z40qxQf4Q5FfEWfzKbNahp0ZuFqAr0
DrNuuR1VuFeAtmoAWnkeMeMsj+KtfZ8rmg+4KVN4VZ810xp/87KP2RaD1I6Fr6EY
9vjVwc8pKz1NHvVg8iUy5Z6g8SYGll9aRJjU0Ue/17/JGh5dwzAh6hWWXQerKS1i
ChvlAaVmvBDX78t32c+PTxeTcdoFxBNVujfOvsVfaKStgMloOJ4ZSVud0VX3MzPj
kzNXZZrPPOUw9bO9sSmYgqYB3m2pPdC02n7mSRmMHy0JUr/mw/Zo/NL9URtwTBza
Xg1NNnpjkM8tRlOv35a40CG5bZDDgPjhgt124M9Rga2THRo3eRUzQJHZyhW0Ud5s
AZjOu86X1UNznevLoBN4zw3LrSkmClCQv+A+tnJeWEQ05QyL1BlEcdfLUiO0/QJb
CJmo2bBOsp6RtRBVZDHDBI2YKbolTM5YkkSRZ4aBE6zt7fbvvRqnBN2LWMZx7TNq
dYRLpYmGiY9ax3gAe576jxzKBPvMEqHN5i5d3ySDyxj8NwwmjJK0pWyylRLjGCel
h1GspOfcnRNPICqeYkLAwHdQ7NTi9VFPbVbNlYBlgNbMdZBAadHOoIdCmYqG2b34
YqKzSOp5z+80Dt20nygRQqdgjfXm2aOBZjXtpCsn6BMPQQimV6w55Or16+htWbJI
QprJ+HqBUUc2HbyNMu9WjoGcAclIfpN6V6edEIEUvj+DyzYpCxDAnT7c4wVazOlQ
NqK2vtxEB+vFQpLTf0HrtNaxGSixcZNxiwnV+nPh/LlJXtPWQ8fY4Ubsq7NOP1sy
UtnxjhASnB6MSuT4b+9mrZgwhecUNg4kCcn4kAAvY9Vvq8wsIpIRzyqX5VN2mGK2
MDBzlwEchVA1Z8WX28gYu/Gf19wQjvt5a4jt64kQvZ5JcavwUlz+AqJqsTvGA47E
9Q9HH9ZlYMVp4ShBNF8uzKUy77A8r0QrNEUGEdGobU8b8vG/TAif3N9mIjKVpjDB
hgWs1vd3NljVcgQ2IHlUBzTnC4osXST5V8zf1dc6pl0pl+T8fyZIhyzty4iTLbW6
5K26un8AuRcqvvDwm1nshrdLeL/YuNovfia1mAXPNKYp5XaCaRUqilKjha4pttbD
cTVeDoAHfFPD20kc5OS01UuYehYEhsTa2z0bHz3kjeyqJ8DXahI1gvSvdKdrShHu
PAV6DAwPHnLj9jgwD0jvCTMcmVIq+LwIKx8bG4lFDSB17iIe6gXv6TCyEcZfFGl0
b2et3q/Z2Lgcn0H7/0DcW2TkP8eOt6Dy7w1us8fSRtyqW9bmj9xn8KSYIf171ZBE
OxxbzSYnVTxdNO1sLOJGiaIACoXsPlCM0Yp6yZ+slbFmjqK2DTUb1+xfDHJpcY7v
15O90ub4JNqapqgACt6e4ExN57t4XN73zAfWGitdzhM+7CeqrihDi2cD7xebP8Mb
OP2AWbBFWZ66IBcK5ik8vdU0r20qTmEWfqfj1rEQfObNm5qX4xmlKLl9BM0ZdHsD
GUWU7pYToTosaKRNvH/E35ElhWa1aYFXDQM8mSSiTem+nv3UUSihRz0pyznYGJoh
oumZR4tl39POce9yjGDJvMypurSbzSfB7o37vzgmeaYIcSKCS75Pk/1raqgP2M9H
O4uMFBeJtsZwtQnaZ5mrhbopov+lCAlb4l07TCXUJFZmDk+ryJEbKQ2VqrOl82lQ
QE7ihTNr1Gt1N4bTpEbilOtKTJStwBA+zGcPwZaYvTruoWvqSLWxN7KhoO87AI8E
snGKYuU7IQnNK5SexRgbNMCs4CmIhLhVToMFzKgH27EJ8wPTXZsX9R1bXWnmcbju
qSphFzft5Ek9i9BONqaBThtKpjxxuS6g6LlTv15MmdWAlS2webLSbcCFCX+2ZVMo
h4WAIt0HqPNSnwOrUlYLroyKHceZ4lUA5kbv5U7nshvmjnNsbs3dryNDaPa72v2C
K/0tGSofX+vmjaAlxcbX+UNtcQTVtcZPF5QgqN0Mfom8yyH87ZeuFz/YuOATcfo1
kngeL4EhWg5JR1U8m943FZyuZ44f8eqsxp/Yb/tkEowHoo+ueADgJ5oqSXIV8qNJ
NCxriTIQzbD+m/VLn+zDePfsi9bMtMB71fkGOEiq6ONnACYxuehYvvJy3guEIq8O
dHl3bx5qxxu6Sn3A9P/ZCBvZx68GfRhMm4+/ULq/QwTHRpmZ9GlhFKmUBZdi7tlB
eef0IBN51I9FqH+14Xzio6KXO9JGfboKXCkEQZfk+jg4quyCAsv0eJoY3kcVU35O
tkvaBPCpacD5/BH9ywWGkUM8CReFmji3we8eNPye/ezZOarR12nwpEOCADFK5q4h
h+nGpl2KLd4dsi7bR6Jef5RQvJG8jaRlsvpU/cZsTL7hkCIxUQNUMcpE6gD6OtvZ
1Pw4VebhCdYvQZvm/O7/ED4c0CRp/fjsjnbyWxn9JZdeZLTqQJPfsnA+6cFfWi8O
bRLTyBCGITIVvc0OLa3768wooDItaOguK6430WR0m4d3Hpbsmdlsv/Li8JW5I9By
vXmupzqASO+kg1WdovVf/8fVTaE/gHrrpi+tSLrEjkA9r+w+70gLhXaqKScda3tl
QEo4J77LbcTF59af1y9NBPLAVEfH3Ri8xCWbn0EjeY3fGNU0h+LeKMUYlA5QrrH/
tJ/b8dZs/tVz69Qltx33XbWtDBLJKU1IvYY/p1h2TTEvEyjcu264DBw39sf2E+8v
QnPo9cFCEcW+B+glEr73RLxjFiyrcadz/flvOfTwegboL6QoxRjyZ+8GUGL7I+mc
dpwFYfiSR3PsZv9IUr/qMzbuis/O/zxVOhq3ODYY8GJB9awhbgwl+6Ga/bRe9YcM
yhHi1tkVf7jh6IGCYcdeOe15IBlG5wsYUQagmBv09etTQ8fEWgnhHO1w2jq9KlDr
/VyfW9QzsLnmyTIkSvmItHn3Nk7lUUF56kFcK3X8cj16LBAmOUbZJq+Ea3qUrYL6
n8HR0Z8Cvchn4i7r2epJ9pWxfbqdifidNbnG3g5gDwE3KHWpV5jOj6cBzM+2ERHV
JtAYG2vzE3qKmrlWEsGj17+e4k/2TzCR9VWB4nKI1mS9vCo1VaOfxSqXtD0uDEkO
YHfzLnjUT6D6OEdiKnC1EDb2lnLO3SvPYnd/2oUtj6Y6BNutOkBqhu7gFdsojHqX
wfEMzv3yMm7+uLLexem0zrRCxfd7r6KOnAoxPsKZxFTvMJ/gs8aLe4mZvEmZRy9A
eeO6h/6+4tkSQOeubEaS83T+bJTs9MT5hsdjvkiDzuMT3gGtpvaVwCBZcQFNc282
wNPdOR2R5TOqhU143hBZG5lhfShZOYJoBSKUFXMzYc+hAODzA8qF8IBvOPuCYZb2
TIEpJFzJ5PahspVe42LJEU9xv/DvcmPStAOHIvbm2lG4nBDC0DmvdbHrAA8qJtJl
2K1MoWAiz1jeD4LT09UQlbcuvmwCPDihOUk/640bHH7dlV5KN1F8oKwrKuOtgiOg
fyK7J561rLsxwNvuVz+9H92FOsjApTt1CaUYe3QVCvLaqAloUJ5InfOqzocVSfZ3
GG2RWnoZzymnfzGCdF9PUa5kD6xbunIFaIy3u1VUptsfNIhYL5+TGt8KE4Wi41lw
kbY+T4Er16LXp0m0CCPQSnHjgHlI1DW4qbPrZL+1CHLHZNzOzdZKbyRbfYFOCtAr
+hprRRCq3Hbb7FZxSd7gUf0cizS/jlBgk3q8RzeGBzRHKCq+uG4+qD/VcTtUBILN
nmkl9lz1KX8paCa5O1Dt6gpohz3yrHoQ1fnvHN8actBPZzsXZocdwaayko65o5ih
taTg50Bfic4Kb6uoaM8rRc8d/qWL2ieJBoTAhzaHk9XWCJnGH9+TyYDI3GgukVsi
jzlj6zPS5hXqyU7HHbkTAZ5AxwD56an8WasU8Feha+k+syFHE7/I+hN9oFrngCZK
s0pbfsjluviJ/JJ7aXG3YiIBAz1qbPAre9nyiuafLzDCeJyvaqncFbZ2zlqBoNm5
9m5BcbE/xOZx8QiMgJX1b+MTwUwg0x7PsYY9uSSZNmKb3cOOtQTE9A8xGPxA013b
afLRg6Jq3+4woqXwv4f767EQPtr20D/7ubFpZq/wCLcjRWQ4jAjG+sKNut6NAclQ
lqvhaNtLj4IZeaaHuK/ZPXj5mojcEXzq1fK1ctIcAJ+tRR0NZUdDnQjenxLAwwR1
ZiC1xVGasqg/BSW7Q8AFBWOFO0U9YhHoFpKlnBbFTE9hDOeUMyPq9XgWJ/8iBaEH
YoxNG20yPpE2SB6P7TPlzBfmmY35Xxehj2OJllmwarKjlb6pKPfCuv15c2w1zNjT
HmVK6DJA4H16CIspo0I1GDFHYVdHv1G8T640JVE43hb0JlREHYRzbYvXycw1FaQi
Vb5glI8+MYKb/GKmDUB+2oPCJaAMP3TCM7vMAy3+xayT4T6ASIDYhcts5eiw+LDT
iEGmznfkAcoJvtK0Tx0VVtWeF+Al7HmKFuoUYPW5upl0Rw5ufB7aX1DsqG4laKx9
xcwg1muJI3U+72SOn0mod+Y/aPeBMoSLhj+jGud278SRnmsXEscQBmytNy6OCDE/
EyeHE6JCAUEpIj+kPDD3Xlbit7siPcSLBVV6yIoRpjkTU13xGJT2ew5IjvFPGN9B
ehuPvahLmVSpLgBHCPm4wez3pXXQdBQj8DSEBKCUcwKJDTH9mp9zVn95qzD1q30y
v6OSAhyM3/zhbxT+3G9QMZPpxk4B52KcskZ4Z4bxUc0ScAb6VoghEZ18y219Sssc
keiuCvRV6ayvj4qWGP2IVRcwq+78js+AEPYKS6dbdcjDE8V1LDHLr0QSvubPCNiN
xrc6yQIl+nKmqlLOZOLEi8BV1dWFzUqApP8WguGgjhHoBRxRNYgFOIHDY8irI2V/
jcgkAx2XqOiGgpxNSHQ34E8+2jzFlrcJKk2SJL7UFsXINtf/NEy0lkges+lMV9OY
8KLMEKbpPVO+z0F9QwuPREnE3S2Zf/+o51dTfa1pAGn3Uh83lB3VmUoYdhzyOaDm
N+pzw8YR7Ad6Oy7RQ2rSF/kD2hh2wUiyLC9c3nHiYjH8U++ZVI7Ep60P4I7AcFr1
hmNF9dc0sgzcB807zX13sAZkBbUIIxur9b5lB2kU/1DLCePnVQ3ZefrJ9vdSNytJ
CNuu3pF3fsSy+xSIYVbTDax2FdplxObWYL8D2u/UtQIvyxOSLo4YSntMQH1R5CAl
jy/o8g/XFUvuJm1rKGaaZHagM0Z4y7DkTfgo0n8vZi1kAwCGGdj23upHPlHn1zaq
v19KLlYZSlvypRBh1RpPXNf3MsFQX5Oqd2IoHUeKQOUN1g2V7yPfkC4PudnZNDOg
ipQVql0i0GM/jNbXIgbBRJ/V/55LFsqqmj8jYSgH2ixhB4MsxE1dmf5Cbj123EHG
Tu8kx6e52hDw6SWgUg4or6iAIGah6XuV80cHSdgkMpm4cgPmFUGguPlzrfQhX4T0
BjHi8vdceDmoqM9hAukYIJ3VXBpvM+yK3i92HX74GMBj5epeQy3fyFFmuQ6zpyHI
TXwSOz5KyJtgczU8V+Fs6yc+tCdkCxC9PIaZqWlYIH4hWpgVjUBC5wBobLYxONcW
AL0rjGA3YuWcq5L59FHYpfEwH3GdcMIYGljEUl2mhxPPER6fQAfTAdJme27zl4N2
vSFe/vo0Jc76HLiLNdbp9RlMibS5Qti986uyudvp+1p17CE8WQzTdSXxOxVjMmeu
wctHxJGSTbrh/NXJZd7D6zaBzxz52RGh7sxDyCZBQa7x8haB/oeOL7lIksCfDVaf
Ud6C6MqURBxpktMmfI2YRQTPAT1twqSOi4yaBJXxM4OTSba28brGSP+FLbad4Rby
GVnq8H4PiZzKsj0SaUQ5xbf0SGFooY6sfsQC1vvs3sFO/7T0CGyrsjkMxFnEtRrA
unaHh+abOeMrqcJBWVNYcShQ8roPg3pk1EdGtNz5oQAQM2X7nHyJzaeChfJa95fk
Hi2Vq+h1Sn+r6k4C0tutn2fxv4yKdq7dPtU5RAAEzhTKW1qX4YxSYxB4iLLW0npv
8MyNTyAx4/QwSLdoOv0Og3kJeStdKYWuwTH1yW0v/DLijQWY6dIFz3JfM6kiL1Mx
ygv0w0N5Zmgt/iF1ajfHvn1lDyyJoD+Sf2dHuHNg4hoyEl7qfem9U4H5dmWPdels
KwvUnOHcB3UVuBZrs1nEuSgEQFyBhsHRjOMTJmb7eatjYzTDDCJTBrG8woFUBvs6
/h6vagpOV9eVC3kakYGai/hZ4+xtigTmb0rxKjBECFntQKCX4me5WUR5FKCczADt
G4rN6Qz1bFJbLpAcGWDCVLdv8zhefMbd9353DrmHCtMDFQ0D/ZjdUN/MvYsEaFiv
O59ok0bbzXwQXsKxpaNXo/tpbeO5HB30PCMWWc4mZiyZ7e2SRAa62EJ71y/WzSP5
RDBc+0x27WLidrGERB0VlQ/6L6WpgdD4OU2LYuuXbY6DxY3arTjzWZ3CbXXfdEXH
+sR0vnbD/BgTyigzcJi4MTFfT5OVafpMYF2gQWSjN5yBN1dC87RafBkgZaPYW+aB
1c51ThuxhGDWB+oapIiEOucvsNyOTqHhLEb4VfEZH4iZCRNCVi4MG+eX0yXG6YWc
e7hZmFzSevQgdDbCWOkqgv2C/hqLO2N9KVV/GwyObxD9CzlIzF6c8BpMzjySNCAH
jqD8cK2KD6HAJzfJ4ynOqIi2ta/xhU0h5FLZJ8FXMx+hsNPAC/9+PLv++YGN+rqY
bnzYAL+Aitzm8hnWDpyOsHL5JI8/JSGZV4PSrQHyUWpCnv46gixID6gH2UaJ5geq
Z8dDsF2W3wLx2idjYULOhG2IsIAHLtYaR/zTAvqcamWvnU+XPwFzVfR+x7Zrb6Yf
Dsc/Ck+Cf8Jpe/CBgquPTmca4YMbLMniecyCzqIWMqYF5lhZB7stkkOqYGGtBkOT
BLgbEEzfvknqKohfUFxsOV7lE7CR771Kx/f3R2quxwSnNCNIcjCRq/1xQK3HaEEV
7YofWxNh3bpjHVRipfDAOkLsxUEY84wAssY72oSJZWGz0nGoKIZ0V8nBsk8CaEqq
As6Mwx+EDKESEGTk3Xz1fLDGYSILto8fO6o2p5E8tFrNjP5zbsKaNM3oaS+22mCT
JyoIuAwxvT7qa661F19BwphVFI8uuLfxAAMIY+9uQSi3vES/rOFiUcuV8gawND6H
Q/HfDMbQa3vUJDxA220sqVlMwVnpBNP3Mm7fHKMBQ3cW2C1HdVI+jIoc1LZxfWyq
8YH8ipBCkrFoUPEJn7FpxoQFOhR0V8dD1Os1qCO+B6+HRgxpDHSujEX/4oyx4526
VLVLWPB0Nc2tp3VR/ObVts8UDBW2UzQ9edrmJdhQbeAj6CAvvUTJV/xXQqjNnqlx
b2765UOfFChAp5QocJar90bqebsNg1UxRl4N1PlOTrd7QkMKHOKxQVpLE92yE6RE
8neRkG2yetD/zIILBuuYEG7VB3YexmXagWOk2Yekb625YF2bwUAkTBFlD2SPzCej
2fRlOIGIrGfqYgQc7oIfEzRhO2MN1FTeskvzyOn5ok6mHiZqqpbS+kDgZPPHuleg
FWYDAWOc//9AlhYEp1UDko5HPP5HU6a8kNE0M/6SZYvEd+bfqq3xivnK7ZP1OQiO
4PWmApKXt16s77uuJfK7gIiOS7PD10PEh8yFF2XYK4ZLzTraaPjw5JycYYwhPhQR
WCBdpR+kdHqtqJADPZWb9cIG6ktPWYM4t1+RkqTQsrkw720p3gwwG+TbN+h/0vyB
Kx81GkutIsHOHREw0e4W5Gc9/8VIGHTT3nYjAICzTU0jTJVo9pB3DKBw8j/+RZV2
4j9hwJcmaeIjXcFZhkTAJDvYC+0MgJu/COJapZzUnxxe3I2nN4pQiKpvHEL3NKdj
9yBn8ekPLwCR0efq6BTDSag2oOSz/inn9KlCHv7zyLKuD+a/kI8DWS+3lBUz3S3G
vbiv/5yNcUlm3A57oh5w+rdr47LByql2/NptBOiFNZcPG+8G5z157mxfFns5zrtH
AT2J3sP+qhJY72zCz+QyNfqRLc468UtD7tVcWbe8YSiLLmN96crf83QUoco5cEyu
Cqc1OxBoFe5tiTI85x1kQUGR3r8OBhR7id1XNSPW27Hgs50KrX+mxX3/XEUY3Ww6
YNev2Q+Me5IOrE8AWyZMCDXC4UZwLShaoItnAWpKGjGsaMD+oucHHmxRxdghgLE1
rNrQnIZwQ3q0SQKNREMR+W8JftFvAdMw/5vCU/7MYOLutDwcQoo7L8q9LRL6xHky
geUsAwH5r3rvzPfP1RZTjTqH8Xr9lxTqqklv66oQPuYWNWaIpMv4iecX1zZVmgsr
GCwFnfG++Va9NpCTOC9WlPuW53B938cKiZRmpvI8Fl0hZttiZNrgSoS9FN1n2rmW
fENEo8+UFLYhu0ez762YDm4WgdBuaveRphkuRSpl/2TpVQp1tzgb+m1oW/Jp9Vmc
ZPxMo94hdwRNpQPE82YPExRnUhOnMftct0yRp+pZg1MbUDK9mKBlLEY3U6PtJGbK
4e3bwW3Z2D/XlICRjMqE7cbYvZ4O5y21Jw5UCUikM4KUsHFqVGaVWK1Z1yu3hvSp
W4Hx9T261TXUdrayBV40zDwmEwo7YLD4Qma52RVb0A0bOO9zNyB7pvV6xM0DJRpL
/3ltA/tGAeGsSf+dCuvhyVf3Bw1PRW+d2uvLDejcokS5E4bGnB+qWUhIPFreVjlA
yFfrFWR0sZXXQcC9jCRTHyrTRyn20Ekkqcua9+t/u4JhkVcqmk1ht1LUZX/A+/OB
LKKjaXQNiilnf79sPzeIWoanOXUykXB6NZpOSNe8VL0YMXEpQtX9c1MhGp4a6M8b
kQSdITxABl++FPPS4CbTyqgq5xjbnZs/qzcb+/Ho6HSG/U8F+uX9NdbBGnRtWzzd
rnUh1tA3VxAUOBwLIPcU8eZDP8Lsj2rVks9TdfwDQcFsc3CU9mgXmt4mcQ7Av+VB
mI1BfO6/YSy6L+HaBSC+w2d+/1e6B/4VUOQglUG/2XbJUAB7haUkyRlLPu+yurvN
qmhnriMcB7go+t31zwbcEyjrwLaR90aCGwROXJt1q9spveV4LEVJ27IrIV7uVoyp
ByjUEUnzsX2zk4GvXQFQoIKQCaEdLgIUpA4GP7YgkgqIt20btgQY1a8p/0RR0Hpx
uckYcj/Ze0H/nl91UmonqsWAqMtO3ksXQqaDDBBRyxySCKUqvq6AWD03sC3x5nB+
VK4gCKCpaLvap4aTjSnpPUFHkxwhIz/nmVXigpMlPXL5qKYplSxwAsSjcwd+cVSN
+k1NdccWUrTtcOCS88rv8T+9Lp9qJniNYsKP92Ju1gru4p6BuxcEGf1Y915R6+Am
xzlw+OkrtJSetLlXLNj5N0hfdBWHNu3gu2TGxoUMUIclvxtPLrBhrG5JjSnDF/gX
Xdel+Qyd1sMzbvem45uUy4YK0AzKvXifp8tg6nkthAp1ZrWgYQ/Kie2v0xlPO9kE
CzcbU0SM2zBb0EIV7v2jqTti7urqqzRWrya4gMA2XJe0SSPdVC4cq1ghYnCDL4PS
VC9EIf05Eygi2yhkvcR22/sWLPfDJ7Zknlu33bvJZAMkR1oC1ChEFXd7f63koIWR
pmEeQo+Q6oyvbyJoe+3h3dUPiaY2D71bs0lC8D7Xy3WikvJHFAgs4Tfnk0DLo8dk
Stgm5Ex0rNriMyjYSup8P01B6LKPTY74Kgc0c0bK9qjd3q2XUjjbSErVnp8wIO0E
xUQu4Toq3J7A5C1l62549VnY0anyQ2BQHhkGyDDcGa49gKrR9Zk+XF3Pj92QUfW7
xQHq/ix+YoEee3lfzTTnyGpXXBfKkdPr/SoEWbnQhU/4bzP6xrnLF3y2nF5APoLO
6TGNPEBITc8zKctOCYW2rM8+7Zuaka/U24kmfL7/q68iLjNiXXou5auZQQHPT6Cl
Wf3vN6U0Xlh6Gg7YWUU4/Sje5Y0s7q34XSsXSktKSW9Nrw2mi1w87LLwy6oITteo
fB0Cz/L6u00ERo3YR0H1guMIQLK3dswjcuhNvvOmQozBi9Ejq8qFmhXFdBhKwn0V
KG1pdqaO+SwLarJiJwHssHBHh/UaTX8ojV2SvhVhg8vVuGKQZSxrQ2XNqvy1NK/q
HFq8Sv2HiZ+OuCDmJUUvVGDgPnmmKRsZ+0sbqDr9Tbe8BsOum+8EADKaP1Bw4T5n
u6YxTtq9uwZyttOtABlIRRLoDhgtoNSidVxwLClyaEKnMSL1Dcu++3pwhL3kVJmO
QTSnS8kh0dccRFXs3iaAdn0bpEDD4jxWzYJDt5idjSfY5BcjXbKqsAmDdf7b1Waj
nnVeC5yIdqDhbMik6VwAi6YNuPIKkrtWe1+JZ0l8HyYZqzZxLTw9vFlk63HTyrGw
EkGzrlytVJUa2WOJFwuOCoFHzXDlsjr9gzgo+ePoUX195jUeFGMcCeZapcx+Cphi
dfjpjPAtpGeisgrdaqZvWacDJ9JRo4PJFLqpzpPbCmYf4a3p7WNquBk7dPxOplo8
Qrm9J4CKeTp5K/TsWh4BhCAxGNH1VR/GEZfGTbJ0slooZPlRTH2YUsKDXweELGLf
agrPDEFzLD4ZfYtWQv60LTnNSB79plQPuRKgAdIPzJ+UMmuFDJAelrD6yOfZEwJN
g2kvMLEpVxV6Vjwx6quFXdGaxfmw9gXcuUzEEgV82Sw/FYmvVNGFKhZgz1VS5Xqr
C7M7z5N/wHbArQXghQj+FwPDbxRh1WZ5lJKnBvVxKAeVgimqJCUOQyOAtI89l8o7
+5hFuf3CZw9heH+922TPeWrCf4HVqcifjtJr8qaxrECYLe8o6Q7KF5IxkDhtTNj7
CyFKA7Kl7UaWz3vmJDqDuUq5mg9nA4QD2eipn6SilEzBvZ56Ta42Mji+7IUYZcIH
1ylu+6zskmextA05aF+Dyp7Bi7I0kFFl5I0TqSLWEAuW947Ms+7k/Mg7g0a6wRsA
IFrCrjULQJz3wqmW4lKqFhweqhBQXwfcxK1nfZddvq9V0wdi+pvXZesSPcQFpAxU
/VwPpxozEUFgZ8sFQZbNpRceOX7gQBXKmYJtSpj8a3rFctJnv7ViPG4c8YRvgqNf
fekOb8dj2PcqrrO48hEgsYT4dedSslepDtzozSD0o6Box7BOSbXcu1Wo6I7OonOA
EtmJbKpp4VsoO4dTn8NpaaaAbOxnAa5PAnbyn2I2Lywu0C4XoY4e+yO4HVFXAE4+
sWKQs/YeOR7yXSKb+CLcqKJEyHN79ZyhVvI28W/ozCwJtKQpyePe3x5Qa/XXaTv2
bm2toLmTMN9tFGIuato79GBxQ+X81T2JrQsLtmV5uo5zoRRqmWC0h+B9QCNZK6Xz
rCuPAzAZApO+5F7bUo4nPVA/ClR0L6ybOiK0Aeg53E8KjCkZuWnyoaNZ5FCzuboW
n0AVXc77ZpqVa9g5bGHvnBX//KqiFkw+WucquDGw+r8xWsdXqXqkdwzB2fPGUzn8
AeokHom3yZ19ZvN9NnmLv40jh4aBFzpmwHRHUqE75LSbsux0kVtit5Wj7qorD8EE
mFmH603skHYpY+ZSa5KOdeiTatwIBO5t3NCUAoQ7/5hm8juW5gSlZ5D4h3abconv
qm+w1UWq/KfdAgaBP/SBHWrUNoCk8lNcJu1DCUVQ8jvrJsOQsIEkvcInsbIOdWj1
8cBcGbZIfN8CVPDiKcU2kJXMlPEHRroJgEcjx0r5bdXaZp62cwvLbBxV8o5pwQH7
h0q+UXiV5/OBydUHPYeYx0Os7dAMv5PbuZPikKdVdyHxxmrjgfOq7cj/CwkZ6Za8
fiN24arIVrsme/eQKpXWYBaxZhLGFLFWjM//Qmhqg8E9tvYwIeR/5SI1+zmFsBj3
Y4elrbp2g0JhcVeXTEHuxagqnAPfKwW8zAmCafBXV8ah6FTBBx/DLMBT6Mhg4m9C
CqNEj0/zDHW3cHOgcOEDYi/X8JFB7khl/15xp14cKZ0KEfQz4caJdR1y/v4+h1hi
D7SB4ohSPdL1CbBysu5jqZWlXhpTm0Pjv29ERGTzx9t+WXb0/xQsjvL+XLffLZe9
teWr9KNiqavFKEo8EZ87LQah18Ny/F7/Uz9yFK65leTRIAMpJVawHbsN0NvD7DqX
cjzzXQ+Pv5sAFjiPJ8Sbv2GWt7SSHlDFEVv3asRdwVCZ5SWuoTTZl39mOlRxIGqH
Xov0d7Ha3GnJQ3C20JzZ64LCRKn5F4G8Z+3mb7Xx7Qi+3XBVIIjiMNulIa0R/qwX
o3zN5VK3lMhLiDCPiz2ATJj0CYX86nEcp093v4sUDKRLhdoXfIQY38SHqezZB9JK
eKc14kIzNUmHSwcv7GLiLI1cJOK1RcyhD26f28zApC/wHxwlLw8kjXU4NDmKs1A1
/Ge8Fe3mzgMnMp5EOAhj2RV1zQy7N/KgkA1DqmbcI8A/jsvlwlrj989lAIlnord5
Is38qj7jDmGcjeoUGEVes/YzpneVHtVP5X/HFXp9MR/XJf95yGeEl9iJ1iJ7IWKf
Efz71gRGRaJLV22+zFIvA+onN6iAakfKBfd7E8BOPIwFF8lXu2gEsewtpPHrH+jy
5yWX2+OOZ98rY5HfsJ+fYbOY4T6O5HJfECBu3lkjxl9qjE5uhT16aj5wxeKPrRF6
KIo5FbAAL7svKvutpVFYrQ2fcTJp2wWCmXlN0WvcsITnWvrOP/NtOiwkj86SpPba
1TSpxmLBNwAMcE8LPlA+LZFiikvsFgLLXBaZiEn+KWhWKxYzhWgbzU3sFQBv2U6i
2TKd8PklUq3wI387PgjtwNxeP9VOLFN8n/P75xmZrGf8O1jeumA+FR6xPmLUZSiU
yzNUHowS3vJs3iZWAeJz96G+fjgtAeu4yIuyAVddkVSgB0pTy7s1/GPhSKSlBRO9
z7DKf6+pA99MkJbTQZ7EEQTw1MOf6DSqd+0YBUxuwiIB2B5qQW9XB2pj2qbQCaiw
2Q6NODU7bO8ubjOtHZqFthJ4Xor3BlNpIn0hW1KHu1JDaNebqYlbgH6O1wkif43V
MDzIWCXTuPGoO8C52jcXoRbwe7r7RnE3Kh8UQ664vRgsuxwTUEnPmC1+LtadrH4z
pFZ6eTAY9u/R8Z2FFE3ILYIyKr8JOMQkpl1GdIzelgxRZ2yeSCGsOSNOYs/OdqvE
0BYi8s3KhC/Dtm1DuM/XIQVIQdEs0rQ/CSgz7+K4I39VFp8Ktk5zjIZ+FBvAvQBK
0hTLadQMGngEQsA+msTTSYBdtwEYe7e5IUIEVvSQ3thVzRuknRMj1+nWGUbaUxfb
JHDzH2wP6XCU7CSJHu+bBtF+S2FijPzoLGl3p1CjxzIAUYrZjKuo4rDI+NXJhq5R
daBv3tXgAeustF2Rog7neLoJdttf83OWOz2L6QnwGjVMZiTibJtLCQ5PkiijUQqI
aJNkVcB+ry005B8tQc4bSVeUALUZpAaPgoUO76xU9uRRO3zMCBPu2TuaRf5mSlNE
XAOpRJ5htFQKYiY8XDbpv+/TjlPiydz1BuA7WAmhfgcwTGQLQhypIP2fHaigwwwf
ej392E+TE7YgXb0HOb7vgVtGL42BZBYr6dWuiYwmlDClZ+939tfZGolfHnbLR+Gu
hwJVfA1PrmEipYylzzlCdmmE8pomxsHp1gMtzLAoVcP142JXsSU2gD6YVM1i3nxO
Srzjp8CZQ/Wro7fIhsr0wYGNzWetF/SxJymwTd8uMnz6e97GEBB6x6li/Jxe+XNN
neWcE/sOe9pA7H2KZV2f3pC4wH+EdeUzDtcsfGoVj3kIYDSyyXg+mtypg1senozh
cYz8wNEUW8giY6Bfrjey8siViM5lZfjD3F8QvELXXy9nZTs9VyhUEAJa0V3UZ2LQ
yr3NwQO/MX+fc54DGnt53iBfTasEElVd1+aI/DDYX0nZNZgcwyO3vDNFkJ+N6TeR
5uabNY569tgM0hEaFhoFwPJx9dsj/WoskFTPzPbor4mMfk/pzs6dy3w5jHGWHsGJ
LRK3SXNt9VUw0sBtI/Mew1E1mQ2ADN0Ucy6YM1XsAoF53loMZgk58bArfVM1LZoJ
OEEN3IPu/S/1Rz+2Yj/bjhUETG5eYWs7kkrzH9Py/CjYmwWlHFQrEq+Jhrz9+Sog
oMCFE1+NyfHkVLT8i31bFkJ969pc8zTBTfgBW+FIKMaXhy20bkSjxBPC+UNCAUT7
1AzYJ341dwk8GoVYFQy2J4WwiZTNiJyBfGTV9gRlHs/tbRCEBBk50UWNratM+EKp
6wTZIRYo6IU8JfyFqBCfQJgbEV/WQGhdORQ7A0TiBA9nk3C+qcrGmMqwD2SwFhbd
F8PrwqQJmhzHGbkf34zPp5uO7Op5eRUeOrqe6DAb7AaFD0R/Q7Qo0suy9rPRqzjh
9xCFt0wx6L8EpTeu4gnnjXxnC9uMpRoVyrVkkzN8gyb+bvJZQo93YNjxrwDD9tg1
X7F7g/KdjW7nHXvMqcI6YpRLFl0+TaZ7//5oWEX5rtxHGhqhww98/0CUiF+kLwG6
gwbG0Yw9f0Ur6mJfS0LU2KmPHxPI3A/dQ57nd27PiVu35YnbNTmlRUY4l94hHP4f
yenGjRsOQGQfsWj7gIGVawKLNl4hUvDb0JzXporktAr+ZZJuG2MJM+Somskrdpsb
oYpvWXnZVgQdqnNKIM59hw/wOazyxgd5oJL33iSn5pcbcIHDuDDznopNeE7G7hmj
AjaRN0zfFuiX0JnBMl2yOZLy8bLzWBxvJB7IAw7QkxgVUgzjRVrrsa3LnCeBQslW
6pWV19JzRVjDnitC7oBY3QZgfmM5o/milCfJs5JU9jbDLPiN8U9DerKAEUT3jz+t
Y7uamC/JCYsN2C4wXsMBjO2fcFlg2WDWO72562qTDeOYWIssrYLbedZ1af+Cx7ap
Y60pUpAPM2qKy69MDUl4eV1K5+8SqbNRBPluabbvUqKG9ijivtPLdWVV2owpGoq+
BKPCVRnep0Dn3nzYHwO0fQ5i3RIAAYPnS1QRrys+lJQfNsI1c8WGHF/Rk5JfGuT4
4qD+kpjUUdobksY0/wHxFGivho2aJtailZrUp+Sv8YLY80I3sOk/izHRpr8ibkpi
GIfDW1IDl0GjocCFIZsnqK3pJ1T+v9n9+FCIOUv5KhbAGIzyrfwzsjzxmWlleqVt
CJVtAfORWsr47u1+lg9OnsmZ7uAoNGV3aZZZ/hDoao6T8rAzxc+gE+FrYwZEI7av
velYrzx1mNpkBbCgeaot/WTYFoSwmmJxiV/9lKPPWiyBk4Rtz4UbCX4PZ4l5ZpTn
M6O9OnkkwEjvX4N6nvEylasXn99fY+sKGEtdGVvK0qkePhjd16Qt9BZpZbWOyYer
A5E0Zo7MKJONAiN8dyNI2J+WDIR2SLLqOqu7uTEluHL9U2Sa0b/k72c1yx0nkXfD
wcMMJVux5TmUXTopjc4y66SKIoeMgwZcDeM8u+g1lE7hZXfoWNQCmQ3XwPttdwsF
4EEF4+EW5caE+xiNxJdUsU54qh5nHiZ2rfl9rULyH7u1mlf5GnqS4M+6cF8QzxlX
HRRHLyQ7kJtx5k8j8JeH2FRpMzk6nlDiemZjO0CNC6R7cKcPd1BcSiYSWR5huPmf
o0NmuE/wYPo3BesRc2G1RGpKiFSW8yQZysCMdV46gRhBIaU5kTqyDcUL9eIusbJM
mzZtw2/0Shs3/U2l+vC8G/BDvnQwJnLca21eImHcpx/meQbzzIEnK51xvX7rYI3/
n3S7CYWRRtZ/vA8TWcB3U9JZS8BfGP/Ohhc9oeisJWn07OkujKVPEJefAtb/mnKG
6dSYYg4EyAJZqDFpVVtiNha1b53DpeBGY4LCragYJAFwszELXpSVukkoNtIiJYNU
YMloslCNSXvqf5eSYZ6ugZE5/mQXA7/B00WL1fFKneCzM7aZzxHaUIS89oDxZz19
8S/gMLN0xitU3CQe032peGO2u4aw7YlfUphtyK67iyXcNQMuUwy6cvmCdczAkjEy
zsW5TFMiLQXTPUaR8GfMHGsvOsXKARFyGJb8XNqwxZjtiBq7I0Lb5Q3AALk82z/3
zQ1LbY3wfsNpZLE77XVB+hNUOWt4d4nbH2qzQRKFbLsiZVE7P0SHfXDmemtf/vqP
a//d6UddWFkErwkmzLRuUSUYg1AGK7qlAGxlJMxOdo388gacphXd0TeCJ0NY1UCf
2Cvg+q4ojNi5s3+NqZmMCcbX6dHBQY8QTbGypjFE0/4U0dE6yabgNZYEuOUuy+gJ
C+RBbErSwBeJL72q+myNPNFblfu77qSlCyC0+o/dLys+pMM6JbxIA/eFQhqcZG+w
4malNLPEa1LmhSSRE8KMU1jRlCcpdimlDBwWBMfCzjkQMs3FsDaGCXizqns/yZY5
WHvFXSrnkLrkIrNXFTrAt88motGqSdjVnPoPyVZzlNWw20VRhev4jBTk3KHyyanZ
vG+hQYp3c013WxVaoyA2Df/SJcWwq2+bANPJM0eI4Fbr/OBhcNe28i+GMXemx6xM
bhIdID3VWmQtQEDXRjcpLkwCyGa+cjM57SBxjJizKFyilHTiBgdq7goj4nf+I39+
VIgQSGjUo3ha2ATSLz51k2JuCHXYZvXlmzNlIxf2u625kKiBXikclJfcSXi6t0IZ
bS0aCCk0pTzwqjgXuCXD6KtjvCf234W14OweRhOPQyUQyyCshOX4HD36p91xuMfq
rY9oiwSW1cYdtQWBjlpwBVto0FN63TLrrnChm+vgUoZx8dKBUpKBgiWhrLlYpYHf
YfVrr3ErJ4DLvv6F99wWEY1diydcxFDj2hVWGYxj4qY95J4pyn4zXwVYbGD1N2m2
j8l4SK1gh+po0iQWW9Zp1djicv+hL2388+8ggWm7ya0vB6TvR+twkbNEbDke4TJS
ambREFHy6T6cZGBs/sTKZRiRI77glClVGpMkQdS4/5GLBjBoVUaoDEvX8nQnzSzK
k8/lcikBFzOZhQIRb6osw3jYC8vlIaQtJ8lflqLoOemxBjkxkxe0iZloKXwXmpd/
IQJSIVNULFJR3jSg1I4GWmFPMhCG/j+n4IXqkZt4S0aW9KvV7LOnVGOGcnFIaMvk
GKyNu0He0gkaJzewQdcGRjbSzZuVPQoou4Xf8G5ue1vH4pqWnbMBt2bwN1zB1s+N
JNJs//5YKhOAnopAOK82Ku0xlEo6Qx7a04mt1fOlzTEqoYALewIAkfAwrWICNmnb
6aS7Ua0DKZ3j1Qe7cUip5jW93ddvADinjpiOCxhCEne+g3sO98UffWIlBfpNko2h
eMGdD8BwNpIxOHplSZZ9XtwoS89MNdCeJG9xTRBHTzOolwUT8ZHMPFiZ/R4TsZfD
VDWj52wuESBCLnL+r5UUg32LFfsU5CSXbF6SbQNLTvVR/7f35lt/Pnw0yNPq7HSY
0icYpmjJ8Sm6ne8+f03fim0Rb6U17aBSnEQVTyty967QeJAYkwvTQOG/Hn5K+rQW
pmDwsBaqIGM74xqwvQl4q7JyCIP1rH++BfoxPUWjWE9GZBFr+JzQABEejQ1+OOg5
Vpu2hksJ8gaZKi+3LzNDuke45mcjHcV1cA6qBfgmc3e2h3ObCyx0PcuZJmVy0DkV
E1nN2AinL6NdDp7wZ2x/1xJWIiRlNAARlQlQ8dbcCqws+MGRdgOXYuNwBIH+ocC7
Cl9+Wc0mdx+Xql0SDlz96kCAn+1Y7ubyTZ3NIAm3GQwBKMlk51q2pmvDMKBIuRmN
QeHF2ytb/6+u62hiL/9H3ElkwDbQmCa+o5BGhYPxZCyqsJr51rc9/UYjH1UW/OTD
xhKkJpNjaFyjgbkg881gUyvzUKNfb5500rYTX0YAe6E5VS+xs8q/I1F5/QTSvlMC
l+RpG2HAIC/4eur+l3OD6qsuZ9wMm9+m56IwMNwRfmk9U+Jr79BM6zhSNXp9zqP5
gDhhjwNFbQ3V3Duoo2WLL5jC3yPUKgGQkhiwp706gAAZlXMZ84KMpCErlrNJYvRN
7E5pJrd5uLybL5XOVq10F5c6QtpNLCvONNfr3MiVtwfIJrtCpf4zsERgfS3uaye7
hp14u2c7IAjYP36FnA0t0nprsfHsocWDK3BR/YCXhD7FkS8nc/jQfVtvyOu/W11a
aOxT08mymaag94umbMAH7K/tLLZJ4UPvhxpMnx3HzN/Ija9SnkRszuZhtluUVzO8
4LoxDj9krU7jdEvtF36wkD5vuq+M8cr0dqE8d3S4NCzuHH4SOvA8+YVwEbprADSm
Mf/MXjfrKAphiZHUj9Nyo8YXvIPgQZAAE40Y6KyksUuzUu6JIe4EVtsMl8A6n8AW
hW80e/A5o6n+6x0q+W8TZSf5Rl/OmutG9RijsgH4YDFuA72koCyRS3KzNYAzt3mR
puI3ctpuWD401EsybOp3ojMx0TPId+h/7ctYOZv/j9xyNLcPAvl+185VMIDdzKEV
GIKk/1f0dZ4zMLdvqZMI/HKObjQ8iikoXVKmExPL8s0syLdmLyAzFVMD0R9ZQUY3
iMMJgRnnELgg+orUmpwwwopLeiOvAeEaJF03ovF+cdhUvfJ8O4Nz3cSFk+9Pwbcr
AEj8Em79PIRRgCLCQyrMyDGsPSb1esgmBeW1agMRecVw0M82EiBkZXyqHQRGAdbR
8vkIde/KeSv+T2/k7VXs7//RcdjOOKvA1yiHPigVy8A6FXeill3FkhCtuLP+CVYg
EJ8+FQPyAhvuJvM4HbrMAC/SNczo4RHtPKP2Ni6Mj4/x0xE4o7S+girGWL9zo1Xp
Oq+DQekbKlPcVUGcmbDOhcSPj1nB8ZaxgBTW2z3Gv/RarfSWSUIx70SLurMVxdun
vRW/Rk2ON7vt+YQBywQeVjk7O/Dekq4sVNl8t46oGWvWhrI8FsLABAWMLeeJEFvd
2YKtk3YIHW98o3k5uqo0CyZbWyQWRAefBZyERdHTZJYGxupwlcOEvRLupSAMXAEm
Yk6s0bLgNkz197QS+JwN22C8/01VGYUxO4hEZGP1jnaQw+eJ2XElJEbsJMCe6sgc
1YZkEHnuepBvqd15aQuGPR0PeucBPthebNvZs1XzpZH/v/oVO1p/uxnhssy0Fuex
t0VhsZfIpcC5XycCNqjU3w44cRDBMpEwWiz2hhsecXdmPs4xu1HbwGhVatZHJFwW
I0nGqJGPX9IkxrGRdfctGI8B7G6tDh4x+4k4nbqp9T9T8BXbSU142RBKhDwQpppj
G8V2RUmklk+R60xuioBe5HMg5imyuhgAUyXjVNJrifG+8JomO31FVJ1JfIpjy6VA
paIsxZMJ3QnG69rItVLar80FEQHKmZaCrc0gUdOB/qIBb3jO4j/Vupd0EaU4zj6z
qM75QkmqBMaHjeP7hWMGnja3Sw+6iMqW7iNMVCIJ0QB2ufyyPYzJBPZenTjA1QmV
VgYImZGJR0E/rw4PXHEG/6k8fSkhLdLpNRd1CKGDAtk2TeNHDBpf0JURXkaU2djP
SaFAbhALTZ8JZZVewtUz8JJFq+lurHkyzu5tZKNIK0gVG/1eIG2cECWfyym/OmLS
KiWVuySrjjPEFSB6h/v5Kq6dwOvUC5t6d/hjydfy+potlNRPHXVRt0Nszu1WsTGY
iygPrpgrbh2sNnvqLB9EwDvl9gyY6fWVp+owBHjlZHag2UIlSVoLsLtcupZx8rjf
Z7jZ8Y7eMYMr3Hbb8ydfEY09g6Dpy7pnQmBQIgtqu6/APXi9QtDnO1+/m+YG6gxH
JADRu8/fS965ERDDf3XO4E0MM+tnD+MMGPxP6tKYOhf1HyEna8xjtMxPkzcNEptD
A1oJvWsuXveLsHaqt7J83nJ4KCk59IpLHCyterqJSJPEwx5N3KkiYW9wNwmv+PUN
er+qF21QkqxAp6rod0D5Lg5BL9Yk6SWkDXbScXeo4K3J8d5fO1jcSLQ/un8xaXYz
KPgt228VbHCnUMOXYO34QofGDh1kVZRossQRE/IEATNf1LjhpdcKbMtXxt8zr4aP
g2VnilgRO+XR84rMqBYBFwpU98jLU0VQkD5ZPO6wMKKag4jVCfTlgwC2JO5WIGMf
pVPJvGvqTdteo+U+dsSS+Xa3XBPkSmlq/wPYkRc1T4Ps0KJcKWo7qYkeAvNgZD0r
BvOt6hUe8PqHP5NuTy7ZtWAMgrQtokylPAifraDp9S/pdMN08RSJFQCIDF9cJImb
85L1dE2BIbqE6FjAvpGR81fpCE9OtrRfOFk3BzRSOLyPZszs3G17q3SCr5iN57GL
RtlgQZF69WCZeR8iMKEctji+c8kzzbBvqvEmwjF1PT60OFD1PBy4nu4c4t/imorB
7xburwAzJEC5fID/6DUBPkeZnen8s/PJx6y/V8yrp/Iiyv2k9K0n72kQwi9bKM4u
/drn72AXKC0NSj6Z16KxEFFKXF6+pIO27MeNNeDaoGTgDvKJrSiYweBJS2vBzBPz
KmBNF9TjrxCYpZ2I5R9cCWHH075JGckp3aGUO8xE96VkKzh8tNKDo0ap7Zd9Ml+F
VUVoBownWCBaVkjHHx00TCjSFYx6eeHFRl0hO6er/LXchDSCH6ZJL7CTuhTpgROG
aDI8Nhln1ipGr2EZXnmyeTTBYEEroK/L5qpQqhwSTazm0peNoXbTBlxZM7WGpixW
uPqjRpXQA5vnpZqmyaTLAn4g0Ht2QzAs7xHZSoUQIdiDniRkVb7beTghxDMSb7Un
8CcWvp3VupxJPNLgyG6M2EYbO5zCtPfmGLFtqs63hQmRXCSNAyEveaexIZ4V9GNg
Fs++1O51V6arrKQS0Exco5AskJkU1mscvReA5zVgKtbioZhI8jjIvP4UEGtTK7tr
nCxdE/O9mdF5hRDvrj1ylo8nWfpHPNMVL/NY0rhyhL8nJSH9d07EI6xZjp2xGmfJ
vn0tz6kc4SbHSkaHslRA7bDFuiRyhHDVLDXmPciuE2IAkgkT5jXie6eCnd87/gbK
2saLA2v9VBEctNq46bHk8mP8g950p4PxOCDLg+z+GTyvGJ+TERhTHQdgcNxiKmSd
f4WvBjhdjyCrazEcrCH+9p26hx4KO7YrWD0Y2EbF79fm4u0zRk3PA0AtfQ/3tE9P
HMM0Wn8p4LgwOp5zbSOhhJgLAbO4CK9lJhJczdOH/9pf90fOLfJ8FqEbMtGuVl9c
5FvXDeX9iH7yHulDb5DldgwohOxD8sQnyUQhuHp0xxYUflIOLQmRAuIzemCJOM1W
+L4h1d7MA4PpJMhVk38nw8+sisI3crjBBiVi19d6vNG0AGXUJV4DSitWLbUqPI9A
IIRzZf+2Z2na2PqmvWiXofAw5FoKNzsqWj7eyc0L2bewP0fxZYQn91vSUn/2kbTe
dRDXDE0lLKN/MhErCu6v9Q==
`protect END_PROTECTED
