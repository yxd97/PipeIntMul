`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
be+JIJ4Eq3ldzFqgwzDc/FSveI7UjmMfgMGHZMibMBMx85vs1i6apN90XBxZxPRi
FHiJ42DikK/AveueNKDJvBYW3VN4+6ryt0DhwZ3wE9kKrMrFIuv6lE4Ah88NcLVo
Vwt1KNwej7PLm+AmXldPwfuVBrdCGvH80Q30qKH+KZagMI9zYn1b9nVMPykJDBu1
/9+of11ZX7cN2i71Y2S8nh7Fez2KSvlprrGqrPHSWTjvVibZGf8fHpZcdbAb0GM4
kpVaVImIgT0p/3R6XyeV4HE1vtyiWQI9S0f5qnTTIrRVVexk6FHQfA9kR7toJYVI
xZhfL2RMi+lJpeLCsIYr7y3buJve9fndPDkN1dSCSioPJrbKGA31XSMd7yWvLAJa
TfdH+C2+qCdSrHvyhNbr04tU2JC+jMDMeLdWQClK0I4=
`protect END_PROTECTED
