`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twbko9UmNNgSrbeZUWS/ngxdnDBSFNHdH3LKoT9+TqyH4/x6wQRlGumdBwowhcjQ
YCWeAoZNztlhoNNTQEpBB7JsLrtdMCWWHiighQi5tf/A8CD6v8cPAnfC5DI2rQxX
UB618tq/b+JHguleSMNDus3eyZWfdYHURoq5fC0e5nA0J7LVeKJJKAHv5mBE8EDW
SgVkD9oy5YtoaKW2tDQg/4ek+TDwjOX24F/RX5IdejRN6Xl1ivUT1FCoR94cQVnG
WIPvh6jqvgYmhwme0x42S0KR0KC+4wOINPLcYxyFndyobu9DbrrL2z+LXxKwAJ2s
H9HScHg46i/+LK5QtufZfw==
`protect END_PROTECTED
