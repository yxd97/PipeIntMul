`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMN2Vl5rNbgzIMJXzae9j8+PpOCJCuAR0jLt+uyhkPIFjHMvdiBCq13rKGvCzf6W
G7tqnrSkdw/uxkMByvrzug49IK9kecr1JiqwVT9mwUdVbYBDnwr6Me/IP7EE7xmD
R7LcOjSJv9SSZoUSXrJPX8n/nKLQVTEhOM4HwDxeR9vIPyLfI4m+Cibjby77vUky
ss8mekho3oSbA2BlbYslcg==
`protect END_PROTECTED
