library verilog;
use verilog.vl_types.all;
entity OBUFDS_LDT_25 is
    port(
        O               : out    vl_logic;
        OB              : out    vl_logic;
        I               : in     vl_logic
    );
end OBUFDS_LDT_25;
