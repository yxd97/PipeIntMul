`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TypO/oJNhkRI1+7NJ8IapVRR6mimWQOo1AjW6zfloMkaor34/LB1Gy+g7quFyyLf
+KyCCfRxr/wSGXcncE5FVMfq5Qe7udp4gvDnSDZQHUfiNNpS4dj27Vno6Ol48LUD
BAU8SpC/2GIp5RZD6P8PaHJI/vPsO1gZ0/2BJyirTmd93N3tgf8gSdjTMjb/NhAY
DjUh24PwapD3lQ0ecxTXOr4vB4t5Sy+WU7V2vwTFLyaSj4Hzzgi0b+iacdN2ZrRz
VawZAzLD1Oa91QjjJ+KnTV/RxEtSEkfQeUGnNw71l5tdfuDqpWClgU/0WBM8HUZX
rXq59feR5foXc7X+S+JBLZpP4avJUfISRAscCAR3usX5ZLdpwKd7KidVw+YtB82m
/Gj5rJB6zxNd+mfMWTq6gMatwZrqmMEL5PF2+NboTyyzFh0sMM42lR7L6AJ70jA+
MLKToLCgHxdo2DImIFhp4BSEfWzsSZJWguuicZT+TC/AdffKfTSRr0ZLseh4y3p0
U01IRDvxlMfpGIkC6EhDYVi4DYQrd2XqApTWC5PvKMSohq1mlBl0uN8dcNGoN3cO
nWIzDoVMvl7Z1ieT7W5uH6pCgITrUz9qTPzVGq/O7hjmYHue7cT4oYMZOjWi6UfB
cP5bLilY9/uyE4wPnT0uET4q1kQ8fibf8fZhUPhi2gc=
`protect END_PROTECTED
