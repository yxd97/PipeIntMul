`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2v2IATW+ebZOyehUbtWWRcbpLJXLCsuZ37aE1TSfbEx7qSpeBlatOeJdKo5P3NP
hYzFeFvuN30UxMpceJ5eruSJCtp1JRjVQCUSp7U5xyy+acAv3ggdh/5EfWWDhljO
Fn2/MJNIhCRVfkNikAdBtsnRleTH2WBVh0EPbss9taDB5XI9BL3hTOqvRnZm67mw
jZopn1bNNO3oOoeTt1/httwhmrz0KpJU5Oswo+BUPM2DpmwGh/CtbdS6D+016/FP
Mx1CK88US26SRovERVsdZynbRkeUvRt+H1P0AIpwEE4sczPAi6C5b7G4Riq9G/jM
O+RatBrawRyFNlcgQvAkCw==
`protect END_PROTECTED
