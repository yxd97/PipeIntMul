`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SbcecU//lPs5eHj4xVahHYxrtL6igMeOXrg524BZCC2q56xXviOZejrLVCFTYyzB
BzSSu2zfn+SS1lW7ZjSS47yS/kZ2FqD1u7NGHANok8LYHt2fhP5J3aNSsFrtKxf5
TL3r7Ac5nc+9gC2dvbkUYbD09BSAK8LKad+OvCG5JD/txS2TwC2LROymTtIwJYu1
CxhIwMLwbClXEnuAi4LWwQ4jT4mZ+FHtXO5gAvzMXknNPi+B+AxyT3C7T+BGPIHT
q333nHskO6h8rzif4G3bWXuGfQLeYGewXOLZrvkVF0wpAk12fjwelcP+/8+WjTYB
YzGgXgeawFz4KQmDafk/ckeoRWRaGpcinR6aoYrf0aqRD7Vg6J2BkHiPzh+WsaF6
Oyb4GxUhYaA11ChabdPOSSGLUbZNgarVFZ8gOcLfjD8cPxyke8ephlEFIA+/5zES
O3T4JEUU5Efj3AOPzsfqerliQmbVhNF1MoT8IfLBF1PWKrejtYQ8EOygQzVS5Aw+
`protect END_PROTECTED
