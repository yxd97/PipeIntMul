`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HE9czlcCjeB/Fxo2tj6ImPHakSE24KGzrG1Azmw/sTcuBYIH2ACpJaz0lQmOXjlM
grmkps1S2/Jbcn86QdN5nhB1u+0xr2A0SpOKqozZfcZtaximNrergO5XrhfcViO5
m2TdTQo3367iH9YbVudSaXGztol2dd2Fn0GCTxNDxKZ+jwxMmWPtbzZQNN7oHSem
5k5GdIYETkPaHTK6LsJyAHAbOdkcDDsTpifygnHQqpU23m867kEAzHusxgbKkKlz
W/tRC10UsZhOAHimcguh7NvOBo2v7GipFqEeNRR9durr3AuXuCIXOmoNYXRCjaT3
dKyN6S99V5adjCWLyv3Fqw==
`protect END_PROTECTED
