`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6jv3zdwDrS0/C5ueb1OaoaV0CpB+jKe+FkLmMH3VRFAJARg23ifYrkjiyHLFcQl
33UcZY6jidQ1Cv6xLb5S0wwSUdZKLGKEJzymm2xeVaAjn6cOrdpSypqppUEYJCTa
d4S5UK1xRqCiCF9eut5C7Ab5XH4g15qIDZ0A9GGAeGEsxQypbMOgHRyVRDIUxdX2
hb8ZJLwpN8Ug5dS+WB9rLJUtgkOiPkUNXhnEcCoIIjMYXyqTWnNaLwPgxSqM9Vxs
5EL1shfGfW1zECJTy7vAa6NVmVRwqCkBcZxNwKkMkiIxVa02B4E2oMchNMfDwkDb
eiH7NxNsYvD1w5YfPVgYtluipw/Llpvrh5oUIo/sxr98uWNL4qw7dC7eUEIExMJl
CwgpcQ97iYXF4bqf+C2j2nVItPNQy1dIt/7rgVsDHx7sMeb9hCWMvch3EuZCEy38
5j93OCvR3UIyaPtJoccHJxPXZQqsO7cz7JhhVm8boG97cW9v1JW3aNVRFta5wvMa
`protect END_PROTECTED
