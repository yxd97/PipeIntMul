`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hkUY1zNXzyjTZMZHE9F8JhtgbCnjZv1u5ff0UathYWPLBx/up1av64VWQiuPkLr7
XSn/4bC1KXYMU/JWHnEY+GGz3yulrqcH6qKdS00DSvb2qip56xWfNXRpv7ekuDVy
J/WGYRnsUzqHMSSKtNyJmKBho0F5d1zY8cgnqvryba1PcRprV1WG0JpiW1ugpHq3
neH+Kl5Rx5Co7pNAE7PeAFAJNh8mmGbQPmIjwrVW2n3Tu1xTJEX3D3ynGc/5oGL3
hgydxpM60LhLWy5nvWsMohsY1mXJxZlNGh3SPwR2PdOrna68eXWCBxZOY6RialTb
SD+ZDmzQTvwxneFYpGWeFDT5GWhJYz2YXUwcbG+jHbKs7EuH6uJdITRevnV9inN7
ZfFFNc46ZhTfMOdAZ91W0Q==
`protect END_PROTECTED
