`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5aT9QOIjiwunMZShpDsFPvTD1j1/059pLbr5XhsM3NTP1zODWVb5wfUsquKHZFvA
CMepXW7p4Eh8bkRNTNIrpaaur5msvnSgvlv5wYHETDyWwH00LzfcBynLVCqkajD0
POwmMiHoAzY/fe3xO0XQP2fB5zpV6czmhYGiVJSXtb7oaXGjR0b3HHLWJv31MJVM
XXwcTTwG0HC7ADPgIOeWJRTLDCFaqCmPHSgeuvycUyPSqAvO3MbPUvV3slPTtZPP
1Q/RQeceWBR/L0Lnh3tJAGLOw7yzsgMAEF7912qlx3WxO9V7nQGBmrzDP3OvACbz
`protect END_PROTECTED
