`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j1KS7P9/opiFF4bZHaAj6mPVN4LPAyOzjgZT0WNaXv776MVbGOqA/vHomanUTiIf
ZdjP3EqSyid74Yoiv5XGEs7oTUX9ii6Fxt4hnY4Hf3RJsTFqRzDeSnzgsO8EogxQ
L7lz0djHsc2XY6/4nIMivhDHgBzrZBJHA0VekOQA7cl9tD4zzrbFUYNcMP1Q3gm/
RKa6Zw8ZdXWsjE2oE/FfpWB69x8qcYQpXvQt4EzZH6/8pUkc+NDfAljS9acBIhvC
NWn9ZgLMMNgdKJ5kFeTqvt2GZlO3I9XwTlNJk+HjmPLcasMo9wAneZgCHZjaQQ3J
nEjyCRxcIPik07Y9AyflOpBn8MddZPYxaj/1QhW7mWN4sF52jHYzmx0MdLvrWKC0
XtIGVEzVLKnF33BvqXFa0KkrZv8DOe2lYDAs7O9eCYjQPjcOmTp2HgsqVeXSEeim
FLlrDUSaPYwXMARJ1YUNQaGO3d+ELP2EAPG2YOyz46F/GtkfgRK2Vg/UExzXSjHO
9AHd0MQYaGzExQ1SUWGp0ZKzeT0OQbFP7S2f3JyrHZpPeDcILx9LsTDF8JaVv7n/
pGBMp9E/Zvn95+otdgtZJFCrdkai/HvcPzyRCozqcjY5KK8wOWPx7rx2qtYuNMVY
sx5yN6bGfTXVOb7OM2q5mHbcjTrgeM/9BQnUgMW/JyGTsiHGdAuWOYtZCbjw3bH+
ZqbUnbRx+uDTJISAH1vvUJCd6WPj8REkHcapSJkq3yo8CLLBBryKnKFcV7s0xXFW
`protect END_PROTECTED
