`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EiGJnYBeaA+YqTTo+V42Z9jHs19/eWZl+2iDLHpqu9ZhY7XMfSq6aBcW/xT9j0F7
l+pfPPdv7ycaF+Y42PhJv9inPV9gvPZJqA5XGkZrZnq60bhJkHP1YYdPlru5Dspp
QOdKgn6K6BwnJjZ74VLGbmFPe0a7Au2umqH2J0sPD1o09BBCi7YDB/CThSDOZqMm
J/98q9Tn3/LRpigMQ2lSiLMNi7ktQKfMdZ1mofrCElnFddqZBS+Da4BNzF8pptOM
lLNa02I9ckDTTHEo67cjdw==
`protect END_PROTECTED
