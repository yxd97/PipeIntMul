`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eqhnYZT0QZd4KFYgjeI3+EI8pio53VrNgfCzykyvSS1gdGi1Y+kw09QHsPjNSub/
nRI4gwWOopvhS7PlW5XKgTsAFhNoCSSHqt/hxOyXvr3KWRJHxyg8NZYETzjpe8Uf
BzWTKBUoBBqP2a1bVQF03CgnZgaUMnc3np8LumGF6YR9I49H49DPRRFEeNscOS/W
ivd088y9Q/PLHo9yw+mjdOBI/BJhbbobegUDmMnPiNKXBc/vDXv56e9+PE98ZBNV
z/dpweqhlFTo2sX+Op/9lJ7KBMh5YJ1ArR6tzLo5UGg=
`protect END_PROTECTED
