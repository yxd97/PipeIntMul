`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYqN+M8MHVCX/6NV1Hkfva574navxc/D9g907WhyM4g6MbRh6NFzyB8glGNl5D0u
vBAUEfBoCMe7uPhCDgc0pIHMTBSdTPGo1dbFFMrN7PVvQhXsZrUoFIQ5YEWdS5GW
aR0/zzWf2EYqVlRKj1q9N2jMmzfoQQtm5OWVM5UEOTTpvTtymVa0yzR0kqQa5VF4
7H2qVnz/yE4ixkgdf3gHaunuyutWT1sMjixZuPd4Kbq2fJMFNQiF5zTxGDliVqqg
hkACooML7exfjVdqQVx4drPVcrCpDr3auW1NPKGZMvPytp7/D8codNYEt+k1nrf4
QB9uLslsmh8uxhSvGDOUokdLQKVauNfSV9pUarTDGehDvU6COUU07B7MG4Usw90U
9rdyPpNmgbtONrODJWOZ6/q21PgDd1BOqsSJ4Ln5Chp2XE1FNWFzl3IwRaoVng9N
5vi7ZoPRyVuzn3qWBzOQZFza4tRnCvNjEzcdhFy9OjgLUI0Uk+Zr2CpHmgSxUhpk
bOMz72m2nRGqvFd/GfHZVIAo1qAy5nKKEmGizJuL30ix/zF3KPbcX47IUFnwIeMu
ctTJ4fXSmRPzbTrE6VIlFYS5686vU5pooD98u6P9NCxkRJ+RmR1FOA7x4T+OGMOY
PavJU30hHhc10pxcLsL2ggZ/wFoIPXpK2tO2xxeirx/Q7Ng9dcEwiu7ZwpfMmgWf
Bw/Zn7Y2hqfz2S78cKABpf4Of6t5ia5qv0DFgu5Tgysn3xWtUfXkcWngZ9hHtG0c
h6rIJT7Cc5jvwKXTuwWmaZ+zxcmlGTyONqtMAM+lqf+TF73p7epdoZpvk8AVNEwf
B+BKRGgaYso8aigj8VHCALtFDq1N1Li1rIbAFRTbkGdN3MpMKKECxnGgLWN5j3Cv
ASKwhetFWdYQcHH5Knui2vNz6nulD/xpUOeWDmgsM1Xu3f9b4E193XnOSvnkzXMp
PgzgD+9QMqI3nQ8OE2C3f2P/DT8bK9OguLpLM1dT1mRilbfIiAMwT4sIjv2Bxvn7
43sL9GroqGWd6fIG/JLDA5XMRl3IWQUwOzpy9BJDdy2jWs3y01UMopee95QWu3zr
D8OczFmyJT6n4yDH8SLJVLe5tnRg9ATHoArAg/WZdMxuAEB8mpjRxV16RC3UFo4A
5UoYl6tpUtOhx9njFeOt9Y9LsLZIn7F/U9HSscwmbYEUdb/G7v0gKLPhcw1zRCax
XOWNZCkuSv3lhd+KmALUTJIV7qHZs9ElHd4R6BvZ15q/NaUYyEHgDV5bD7f4rxWT
KTiDex8XhglmEfl84JGbtchoWFudYL3CpeLtSc5DqQ1u4ZmqcEY93JtS3ki+yMyy
5x2IiSEMiC9QK4pzMzGRfqgm421qDxp+4Kx7vfOvSe18GnIogIBx8XWFcQ7dAPZL
e2w3C4W04sJSnvkxt3eMAKDuk2GIOQ05ktvYnzRng/O+sl9mVMV8ge5vixGJeq/D
DpZ0wZ8nVyPbse41tnt5OD3Zah6pcUOSpoYIpAkmFNAGtZ+rJbMxnuCOpG0mJjfY
99kcpczBoB02M6ojBxTajcut0F/GkF+AOlWRSkBDKBjduaoYgYkFEJ6F0BIFC+4B
IsaC36fLVq/tk81BYTfRW27YQk7H3PmgpdBpG4+O+nWXKGlNYkYgMBQJP6APRY6O
cR5xpt2nJeRYdtILQfeo1zjsbvFYAudIzbNyA7IMCbrS7PuLFnqoWB+OzGG10SX+
MkuAUei9OsD53/taU3232e3/cXjEqFfvWsHvee+f1f+mfV4u4cwvBRMGxziJs1k0
FnKFDDYHYvf2KD9QdQm0OrJVchRn8Wyg2H/0pkmjdEZ7CcyyNxEldXQkEJ1u8ZPe
vgWQ1i+IEVt6NNCvdzNJyiPPyKoc+gRkxDQ+Uzds/PKCZ46hFtOs3Z+MjNUbyNoi
IMeDeiBfdkDKNJPPL1Wviw==
`protect END_PROTECTED
