`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5f2G+PuoI05xJv42Hxs5KUcM1Vo5l2r6MsgvaMvF62ZkJ/pG2mo3rtT57S+XuBx
NLfykC9+Eej82hGIZjXtn1nfPAkB6Ju/kL2aVngeUH/DzSVX4PRp9HgEwpU5imUD
D1+qoq3dpcgdSlKMaIzs12C0GIYIgxOTo+JRcNEOZRKJlknbNJNIHGYcuE66gBnC
V0rvavNHw2pUdtvQo0XZJql29/W5y3Vr/NJ2ofm46sNU75QPFCYk7JXkOLavBlPQ
hwhOZ0p0kJkX7nyqZ2uB7LXwyam3OxbnqFholXpDIqomtCXPDoWV+ZNmWmMNVO35
f6EBR9UsxGsSJAJLGrcv91L9OINsxyUvv0A4EG5ci0ID8nzwzqRVM8LqrDfkI2Tr
B3aZKXP27p28q7ldwVFoEiHPOEUkhDximgl7SxDKTqJiUbx9uJ96CWX0+gJlnYuR
yZ6ohrwso+MF3UU+Rkaf5swQ9KPuEqmlSOiWqrXtKqI0opqMhmN569la9e7cdZYP
mKPEygYRRh3+gHeIIlwz7rSOmsvySPPRYjfFWaGJxXNxQ4U7Y4frEDuqUkfLJXQx
srw1u4dh7EZl5KgdzWQvcjfIYlZzrvnOcHnXogJnXrIzGO2YRY6rVRGW9BDpkLwe
DOH4yzzfZ1MCmt/Zl98KeE57T58dWL0rmSEDHgH4A+4rSE8k7T/B+rqY67nvu5ad
TPCUn5xRbK1yF9efsrBXBC4kKz48mHhd/FRCbNSdIld56HtjdAAVaJxOrtNh0I82
uyic1ys0DoM/OwzgAYdQ0nU+3xje3BFWNJmKyLVcNK6AGAYdPXLseF/8GGW6ntlI
HWkX2fbBPf8xnzAsDeQLXBa5UjcaXWngko9SB+tA4NXdiM5DhOTRbHVNXD5X1R4i
fZ0yjeSUKG3r7vaEJrKzbWI6ahNPSOk20vPd0JG4+HJ/i3s8y4tVvIrL1q0GIYLF
G/MpCkDHb9vXUxM7UOCHDrk8E95NpOcMMFAmg5xye7OC6uvkXb/oYLFBvISj8a8F
JDRPYLsbEbGViWQrLZLplUxP70NaZL5wwieeYM0JQH7y64ZO8qpoCczcxql7gA9p
wmrfAm0GXBoLn+Gjy715erXh/IOT7BPl+pV5M9QnDlzbBEaZ5p49OCJcIJz18aC0
`protect END_PROTECTED
