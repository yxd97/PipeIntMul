`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bW2d16AAAVNr1H3WfGGY6GuyEB7W4tQKBUA6OYzqiy5s/Ic+ZgQ9jTQXpOxwKxFr
FiU5/XgF+mfMZYAvuXr4nwVL+brCOS4/je8N7aeLrI4sOcOkckUjll4lNvzcLXm3
OZrwm6xn/H13rxX17XEeQQz+KCMBSPbWHQBaAvH4wb03kBpm7v+Xe6SgdtjjUrAs
LqJqetuJjLE879s1bfvEtOqY5aMIB00U9PtGi6N7x7Y62CDwqhC3sXxQLlTkYeij
osauzKRJSPzKJ6WnXmvXQimMPe4abJiQ3FT1HhjbiywyXNLjxfJg5Nn4zP2evu0u
yfGK9bF0gcKfqpE2S/Ti8A==
`protect END_PROTECTED
