`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r0FoeSn4fnQwReUtVLwUD9ciQi4/2Aw4tbvefKzdkG9ACr23nNaB4AtxCHqKsIfk
deUg3Zjb2R79iTy6Km858YUgL78yzkJ/PAW/sM/BnnfZR/W+tpVIZsEzlyMzJt8h
BAEo5c/99GS6jiWWISd/V7WPQ1GilwxYMjWW7e/elK2YyMQWXWI3vyNR8xQtHPB0
Oa/1whVBdZ+8oXY7euLbZOS+4fqct01L4AfBjG27LtsBqRWF+dS7tHiIKcd0bTZW
j8O8D5ePv2M6K+VK7Bc/digAA56Oun19JAmSgyS8mhmQzc28d2raqGUw9BcJ16wm
HEF0XQU8t9FqNzwij6Ubx4uZuP9mARyG4XYUh+BDEkhHGLVUr09aS3cUUiCa2TP0
i8R5/pf4H+Mti+dGRkNeyUff/xRbWh+za5p/nVatsUdzuwZBFjwMhls/h1AnS2i6
J2C3QcpNVbt5GZd5KKgpmqoPrtk8hLV19bMTwOBJ2rTFuEzajEGjIt269hvcnv8M
L4x/4ENFb4EaTFoZRBUuWN/2R7m5ZG6DnjXtCngF2e/bdM9j6zaSpmX2X47yNkdD
PsGMwNx2CimhTOccNfppRcjVOcIG4WnXnQDJtF7reBXus5GUExxUz6XqcFGdeHOw
tIGeOwuay7XMLUFjds1A8GBTALsRmaH3UdLkx43o0/HHxcAiTwEgDW2eoYqi3fMj
8iTyxMBAgC85TF7It1M0gzc39r7sRE30e08Zwtc9ie7B9fm7kfS8g0qwKvi4WymN
Gxa9eaCuCcXILL7ODBFrzdCG+X9qG9rg5VI6gMe0fmaKI5urEWg5n6UKCXswRCcf
v3/KiuLu3ywhZDpHiT4BB2v01qiLtTlScQk5vUZMZlf2dmrtCWZpjvZrX8cvgQLg
u5ydYZZj25d5NEgxQYbU007EOyexdC+g4e4KYCIBOUelJ1nY8TGRB3uz9unI2vxq
/wIwYSnCmyL0NgQOfbX4CvwzPpQ4mQtqasUXGIz14ELWqYv748ip1M1ZhPgn/eMv
zPq+efJ6Ye13zDaCcD60LS7cql0pW6OHybRzVh+QYkwAHkYd0OmK/Ujvnj9XBr0N
cqwiGKPy9Q5cs7QNEK19/HFnmgfDU4lpTgZmjF+epf+VPQtDisettrqvoQTUlvnY
449Y1Y3HKOEsQ8DFbZNGr20+19xQTkWLFnWOQf11gdU=
`protect END_PROTECTED
