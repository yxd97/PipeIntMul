`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xAvInUxHqcXmMKwGZj+F/BZgpmUdfFQZjkZQdcT8qRmAj042Nr8Zm7ZyKYjfQgMU
o1JgK2IgV9ryijPQbeA+84UBj2U/YFVQflh8LiW2Ie810e+epdrnnrpUy3Md691b
eWlCZLjkkJR16hQ1H55PDuGlhrQrkjluS5DIW2JT5r4U74VDv8+wQyKWtixNZb4Q
Zvs/roJ04BrKyAZBxKtyglyIzPAmFU4vgXBKIsT2gXpQejIeciLgH9zpm62HLSQQ
rUEGI/xzR2u6wZBqCqKzPOpJh0/+43K/KmFDhFQ1fQz0E4xTmgzrzgbjxix/jmn6
8L2JSnndLKBl2Ex4W9ipskY2/09fMoVpGRxeB+ORgpTERoj1On3E6e5jS5j7TShg
4lUfJB2lIWwHXsoZL0KoQkvnWOk+5MYhAUOi9rER1Bfqivsxiz+/gc6Ph2PiQuuk
Iw/cycKEqwUPFwx8GVeaRXnoc3A9d+BVt1sptk/JuXolGMyTQ+Fw1rdq53TNtmhr
P400k7/Lwlx+zsKwnsdDNF7PwRiPLFttMImxQ0g1QYsVflVm3GXLMNs7SQfnPWoJ
Ek6K+oJ0+fCjEEZnCBq/zm7//NR0Xt14osXqdDMgGrKh5IS+HXET3MvDumuxcYxg
BrPjx38uaRCShtz0b/hYDVPz7CjwWxXxvSygr86/ukfoV7feONqLhw5M3sLDYYyH
SVcjaJHB9cIgFLW1wf9jUfUOBl4DosfzMLi2yOwuljXRsAFuOSgfAWPofuM721e3
PMKyXnHGGJ4qf/Kb7Zvi7xStcpHLgSe/EIHQIIU27egWLzRkg83Ga3T7C40phatA
8G4m2VuPgXp5BpmWzqF6YWvAeOTJTcuFXabgCbQ5Gk8F1nW/CPG04ZsCKqr//FtT
3CWo4vWz7ySSv8C4q2v5NHG/J20UyZ8LdsXWu/x17IdQ6UbQ+WkjUXHUvaAy657s
vq+TTyunoOUtIjBWWbLiGRhvmKlrq+9VWsWpeHXQm5IA/sQA8bPlpE9+ClAzWrmn
7ygQyJAJo0PE447caWRiXV3EhF46aR+mMDtiLiFzpuzho6ihTj1s1LTBAGhvTcHB
X9xsmF/8GqAk5/gv5lWX+wmEOD1GWp4Zg4nONf8xpU3tkIvbUqbRgi7Ma44aM1wW
zilJ1DQNcF1yNYH7OvFTQnFkRh3qv5F0SCjHd7tjxL1XWB8vSRRMzMnll5SBPa+r
aY6Ya0KaGeBQF5lDnaGpxg==
`protect END_PROTECTED
