`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BLS4KMY91FKFLA9qfKsXcJdEp+tmCqz3SMQj6+w4erTEBjxgGxaZcpoiOXMz4VFl
RAPvpdxKGFiT47n3ne/WPvY0ED/4yDAHmdnJyYhtlmqslYkqcnX9lXRToTqMvFaV
/DKNJeYFppoJhhQzGqJmEvzBD/uHH2ZM7dzE9qumQ1rT+DHECJ8qnjRWoNTtXgGO
wvNZbUKpTOUMQVyzneh6Obd5GtlJDT5hyrnjV1/yIusSIWdtjxUpyJx1c0uWNFzm
Yjrer6DBUpoqASqHMJYCVzTDeG0mmG6/NsyVYhNaNP0V2Oz5YcuKPFZdNwja/S6m
cQ3uk23Ld7RBolurytKiA6IantUspjIIaLZxfzAIjb2SfpHKmr5GrZYI8bDF57di
hTonOdRBzo0WM6/bFH6FqFPMg5L43vd5PWi1MateiT4d63Ip837erK8/HuKQ4xuz
/2wBanM9gBgl1fBfNCeXTSr8Oei6v6y3n0SjbKRkjopqQEvrHkBHDFveb9eKITvA
KSv7m9khe1+nA60h7s4wU9spMe+S+RLmLqkLzdMdn+VN2hvUPoZj/QMAFog+Hwrp
G2veISptFZZGCrKv0cnSghvGF6Uwoo0Hfwyrbi8gZZQ=
`protect END_PROTECTED
