`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2BXbXBkhPaE9l6IDbNyuVy5mFqEfZVrtn66KouE69pdlsNq7ZkTo6lgvR4Vk43y
nvd4klQz7G2ap0s+6kRh+sFdG44DCcVXqaFe7RHu76jC5rIYJPTkFcquXk8ae1JP
HsUxKbkIIN8KJ1eePSecuyHCViEZcMKcNyT98uouZ2PDoc/VVQ39wV4a3WDBAJrD
hmNedOa1aPKusWzucGK2dVzLHUAUwyBCJQEsgdU0H5O1zsZp55qYqTfmMiWiRdui
28Ou1y8wOJmWwYdqweZctm79Ermj+NoCxo3C7BioOV3XGQKCe0hFDAcW2yKTso8w
eu26DYX3fbYxIW1nDvaEy9oKI2OG5O7N46BLwSytGQjlNGjkpTHycw7M4enwXU8L
WzGr7AJgiZyKHkQqKZBriGqYaNsbohZQjsdy7K/ZLShoGzFUY0z+4+srUrxoXR1j
32bx/m9Pi3wqKUTdjqM/3LRVvFFOkvGE/CgEOAfE5y7+XWXoDiHQz6xMRnpctdOO
c9D7w0dZ+nXR2v8MSZNAyMIIqOCHrZF+cSAGOLEeaktKfcDcaJIMJw9wCokwdIWk
cbXDkQ7irgIPAQEBN/PBZNyEZNbpuE3JjFRzOzDjgeqRAOmmmnXy75IkR66UE+73
ncLG6QeF+zxxodpzV27/9flwIDAh/QmDMhmAp/0Kue+Cvr2cjLJSMRjr1caJ7alj
R6X97Udnt2sjSzf0wBcFdYO022ay3wqGZotP8xnndj6JFjp41kp+mUcePGEM6wWP
nrHfs/ODkbXbM9oNwMOWfVyGdWxLmHK6rE6353ylUGw=
`protect END_PROTECTED
