`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKr1pp8UibINqsrzG/nzpnZ47id494R2P/WGIghbIWCyOv3t3kdwG705FpkgomrK
t2syu4kaGx0DohwfUrfsiGkIvdDwaDPor+wB8wJtXH3RTlgo5LKKot9vydHcQixO
YoEDdAGIaA+XCIABQ89ZCEKIdOj9x1a7U7NWyRQg8Yg4CxhvcqW6HQk0QObK6AX2
tWA/Xrq27YeSnxbeyLHfDjr7CnSngmKn3s6STGM7/wnJJWlc4gcS9aeqIkopuRSU
bmkyV9I+QbE5WRvac9AWIl6Cqy7rmgkSoZaG6kJJ85I3QM5KgnYK8iTFhBiiKEKl
Sm6ofxvnWRyDak7HjIDAgKCB4a6NEdd7r5t9KuFzZfbQUpQBP5rKpnjGfOR0oT97
UASe81ODi8f/B2D6+l0CH4FfXUo+S0t0808s6XxXOKg=
`protect END_PROTECTED
