`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xcExdukoWsm5FBA8NNoPDZJ04tUNYYrpin5bh2rDHgVTfOYpPvQ0tq/u8u72906i
kMhR4XNeDIfCxRSmYbf4+pvHJgSKu97SA51cybDZJWlomZkbBVHz23wct7xTg5GL
8XBdXEjtC9d2rk2jbUuRDSL90D5fxWyBgWaKnfVN73xeUnLLs2Rqdjr7Kg1Z9w1p
468KDlfhSpyVc08kQ4dFuROJtZtmzXpfwZ0jFVUmT01Oo8s4Uxi3+JinYQ6Gmdul
MbYBybmi/ZWe0KIyQdVAEUJge6f8NoSgYmeuSTF7JxPbySyvXmNTSbY9TXKdmo3d
R81T8dFTsOGA1UaX44QpaG52rwB0S9ffAsIOmaodRAqPkoCKCzA6fgiR7BhiiI6q
It3po3XngXKtCK/j6MDW5dxEL+NzlbUqHCOIzm73nytTcKhio+wRlxIQyf+pFJ4S
qcpHWLDcZbTs2BbPSGH3QPn7aSfy4559DlPFLYo0FIkjVWncvRoO5vmf8gOwTul9
iM/KuGKmlG7Ipqrwi7Ak973SRplXjNmzxAWwZMXSxj29OTLzgjbDTfIpVujF3q5S
8rSVATzy4QvPXa+qZ2cgnQCW9kgqSTZplt5wJ84IJEm4UjNeDJeHwUrZiTbvybV2
pNjL7JKHPiVRzu7Sn7Klz1tmWKXalfH1/ujrMKvqc+PwHUqGwn4V9pMpq9qCJgBv
D3Kx8FElrXPS8I8uk9XL0fHupCIG2V/t7eyVCmG9u2S+/27WG5EGO9vqyTpw1VVa
Ai5PLGjBVGzdO65F3rnobzQS3hmv6Ow5fafUzfcvrpB5q3l0kh0kQVRF9Sq187/0
uozphDBrNRu67mv3mNP3fjJHtRaPdV9YC5oQSv/IjYMkLc3aBEkdLMaZ9rceb+b3
g6bbXBUcsNBy1CEkqR+Tc5RjR89cE8Yu0zou2yzMrEM27x863FqtNAyu9oCJ85UT
`protect END_PROTECTED
