`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AePrhpHO8GGyRFedomg7vu6ojJMGWLfDb1p8VrleuWFXwZXihWht46ts2Wm7Op+u
omZgi4xvhv20foRsnxSMlZ4tTcBxt/LBjOSGM64NEbyOocGfpvQXwWnVX2ejisON
JDNjlggcxbXDyd2IuqORvdo/LUAgBCAY/zeH/9leJqgzJZwJpZSnjkOansUcxtJt
lVv4W68WCo2YVBmw9gjPdkWULD9Nxs6dIx82YkZMFxxP2HttDiPX/Z4sq0akBFJk
EDdSIZdPmhNONuqC97cNTRDFcMOxNwXJ2TVPDTJLbAXo843+vqE5PY/ITNM5Z9+u
Vnme0OAuMgtOyCQ3c77QccVxkBnvSLbod3LL1fnp91Ri94+9HKc6qgbr2NWsULH4
s4AQum35cnLmhgPKvL76XSjdTKCw1PCwuzQULYj6ruCVOfvXyi6GnwYaqtGhECkd
bGY4gcUgxT3d7exbHx9TqOC1eq277ZB4P1Ofly5Rgr75XWi6OEJFSYG0vt+hwyP2
vYqU0XWyiVBM1Zq7OpvqOIJH7UT8sxO+snik3En0B56+EIXjROXXk9ZrCnX4eNIB
2EWTouQY/Qw66bB6IFV3P79isu2KRjCcvY620zy/g1CNuEyKutk7HA/yGr72zAE/
m4b+LhwiapO23vJOT0qoK5BJhLQRel8A0qN1B5OT265gEFjCpi9HWqHK5/OIRpaw
RZM+Myc6aK4xOc68gyUG0ZiAp29AUoVyfQ40IJU3pdQCibZiMOFoKXut40Rh5xZF
FMobDvDLeCZSh2ubrdrE1VHEwv75JK2inYx1M+qCTBN9TnX3v3SmYvEAEh5HnFd5
0esIxIRFgumlhCtWIX4I+fFMJ1NH0oBAf/Ku7W4J/LE+70/mq7jAOU+SmI+c2M5w
lhlItFXs7Cvj/6CSzK2bFcw6ORmiZX/U8I/YR5hIqgmF7eZC6TodPj1O8/5E8uIZ
pYiuKXrTpsSdm5OQMyzScjIFkOLCUs/MAlBfUnX9G8WPT/D20gwNQKMfX2jLXJE0
T3dWjyu0GeysR7RIARHXFYSyCcdQ7L0ZF0sjWWBdLfJFfmZmWf6I4SLG289NDKF+
hdJ0hXboWVBS87JDCPD3LAv29k/iguJRgjFRJKQd1k+P/0j247IlQv+Aa25ZTzTu
nzVWztIwKV7abM5/rbARhrj1qe2CBjf/3ju7C3C1b5K3MZp46ftFfZ/ykrhFQ/aP
piEEhT312E/QpAa0u4XmzsoIX6F5QVeT6jISqw7lw5gCc+ChkJh+dBwJ6RhtGP9T
+r7J88AsDw0iLLV52UhowQ4nyKN3hwn7R0em/GqFksEQY33XJg+SqfnBtsQB9KDg
gzUYfElrWxV5cvnGw+iGUPoF0PW1oVtLH7cwna3UPPJX1oycZkowrPVK/5Vu5ZKS
H/K6Gu7/L/aXP2pGAucLbKykMvpnDqPLIuWr0GFu3ygW+4ReTjF57X9zeaY2ySZz
4pQdvTKeC1SbviW4ggQVTNut8nhJe80ia+Dlfyjb/Z3LunptzeLppKdRHGHcfFQn
OyHzn9t9/vd4bcb+TpGrJ4SQeE+6foaU3G4Y1QV56k8MxK4iTx6M2shjY/O9xCF2
OiWqHUhu0NLlQg1iulSYjLyueu3Hm76K5podChEVvHeUSHmE/+tbOzjXa0g4LDB/
GyEd2agr8BX4mqPBXEUIiUex0A6amdaLt/8Qgs5ZDa7o/PiqyicuDL0wioSBC/WC
tdtlfjlKEEZk7hYF4LCcbmSYgMlFcTQ3pnxt06C7X323DMF3ae+Cf1hHHIpVwLaj
iRh67DS0MY8tWhZ6atfjvft7hXpVt0iK2l/2fmjWMqRnUCovJhhlcu+o1bdbfgE6
EIDbnDzGY0fGIno6HX5IJfZAGo/JBEzQfp0T8+Ax3MByKFRyQwMMfEoGVipJL0rO
a+s7jnequeUbGdC5kV1I6J0EpmR3rLs+s0LzO2DLF3YnmilNJeRMA+/FzWnz8FWi
kAxGkvK+jWtS6dljd3kuuZM0D3eOMtRgYU+sQyB73TFtACnO+5umW26FWphRIczU
ht141RzuVaMXLy7syb9CdGPKPHIYZhm5awX0xvG87YdAJvT0r6wBVhvDxRpCYyAI
VE4T2dzEE3RI5uSHt8L+IAAeHlsy9SUOZq8RKslt4C6ThGR7MBlmbzYsgNV5RrLx
8+o2ynJfuSqkGVuBStqQgmLqDnzfLBZ3+KN6b7hbkX8euWMvHwIZGb2SO/2bFuQg
yoEiQJK2QFzQE/kjgJ2JQvbW5Sav4ItYZEbR7FdnbjuE1mIc9lbW33gLGOMW0u7k
09U3xRB5XP792i6xbUiSJ9vW0tRrFaLeNxa6ts45bpsxQC3cJWGrgFa0PGXDxyAT
CpDm0onR4HRI3xVil8JSiqlRXqRynlSFurirtoP6LIhY8TYSAel4Y/HwYdpyfwyj
oBc39KhzwziUS0xxwA1VVHgbZXoQDbfD2oJt25fLN0pNhNLijwvjdzf2lGILRVBV
r5Mv+mqZUsO+/W1oA6jV3LcVizq5J9FgoztU/sGckhtlvsxLH5+rBNzmsluSp1ih
t5l/5yMkDgilLf9ayj+rvwDnQBPMmMEI3U5oUdLwzWOpvIQEF2//FnTODIrzez2U
VX8K0ZqUZ/oNNTVKyxl2x4Gnx/Ay5lkoH6pwNodA1b7fXOM52V7sSaiPIm9vsaow
DnrEmmQmJ7Nfq9NRHLdZY9niSIdaPij7OLY+Esb3SzuN0dvVLHiPjV9qijcVbRBS
eYnx3pIsiQ3jXMbParVRFy+XjRR4HHpEmtT+/IpYnWLDClI6YotaAj+SUMk53uIC
/0YxDj4AnWGo9Jaf5KublqjRCNAgbwP7hyTsSkdi/nXHEy3UHiD/Q45m2GcNZR89
I0+Pt/QmdBtOEGCb3zjjJN2tkYE6fudAYrjY5cRNQ2Lt4f/oSpsk1qAV5r/oj7fz
19AXMlBNAAkpEHVsqH4Gcx92Im34gic9FJtZf+7hLnzFQzJfpwMMcpajFzDYkxtf
0ELbU23H1Ne9X7neW2pKU7cv5BzW748dipfG5X6mrtZf1+IIuGyVOuYmecd14vVO
36yng0lxuJX2Vk52zm8Pazy4Vdk79ISadOKq6zIJtucqlcbKH9fZo1oylDPXyNXg
+scRlsRwikksWyEJzWOOJYTURIm1wzgXR9lXMVEHCwKljuQgDonjwBOo/eC7+A4E
KIY6ITdLZ/RC/+lw5Lm7aqqPkHyAzSlKfVyZOKqT8Od8SXYEbflALN1lz4x0optE
7kzO9CAra9yrHu+KOyBuhQyPaqEeyL3Vj/rs/dgJIwBosTJRbRunJEHiyMu0DpMi
rBpOnmPXczUv46KnSbqnHPmtiAsknUd/hKVNbapRPPdrDw4jevw/9neT7xB5MFAD
y6bdq5cWV4SjWxstRnEtYtqjuRK2CnyajvHbSWdbiovkJUO6DxdSk/has9OhYlde
Bh5VwIY7Lykt6YSZlGCN5q/wrL7Kt5GtoprBOgQj85kN8SjydXjMCYbwk/7vyYPT
tjQuVOx8GSkvBXo/ARpnV9Cg/G2MGtLBRuigqPdxmAFjitupRL+c5xHwCWzqew0D
n0zdPBhLv8j0qYvkxk5Q/cM7Hr1xzDRCFkWl3XuN0hpJN5pJIFWorEQAdDCLYmmU
9H4UBXIRgF2C/8tr2BjPpH75B7o/HQ8N51nk1V6NsQS7araK6WPf5+p8UfA0NLYs
ld0ov3GIFSWtBAV06PMLYTU/v/hYVUhVGLC8iRp6D5JleNa7tFYTNdj5tVA+1RSn
ZeDTkI7FIOHrH2HWHL8/VNV0gxf+JPNt9TBxbtNp2i9dFGp1e50evaT6qn3rhImK
Bd9I4JGpqRKGjI0bTstiu9X1fAXi0e8trNhfPfpMtn65Gndh+Mhp9WgdXMrmySIZ
3ppD2G5I1sCU0IPmScOu2Fol91jwAU0lRbS4KivayV1ZtNlGSel6I+NB3jQubkvR
GrB4egAPabqQFodoIcW95wOXPsZrT0kEaa/egBcVA+lvXVdtVW0/60wWRVTlqvl6
t/Y/L4fBomCULxWsteZrZro901S7y4bUx0bC8UAoVEbgB6Fn29fNczUkJTLzoxWW
LFA3n8pbuvr2XS4SufLYVo/LES+qyQVC+ss2dqwk8FtgJLzjK2X5D22uloubGVuh
W0yGENTTyVO9BY0L8AZHfBRJovJrrNebi7ZFd4fh0pBxSvy9NXMByn6bJSbWR1X1
pcHU1pKXeAYjDB+ZY0ikYirJuOediM0LQ108KNYT+2RrU6eVsHBulponMhJYeFx0
c8I3XMiiZhdhRP5u7Y1/b0faH5MRXA608S4glYX04sHcZExBb4sm5bXmIHg5ViWN
Gyag7H5BWKiMzv4PtR5tQjhq9zD2Qx5WKi5RUO3FIXeYc1MXRbQRfnZ0C86wL0HE
7BNJLN8JEKjcz7JplAM0R9/Wr4vKONstPSmgN1qMq7sKWQ+fRV6yimMkb54wgzuR
iNf6x4bal4SvF3DIP/s+EM4D9YAI+iMU4nZjzjAx1L/HbUJ8Jmi764wccUZnyD+D
5YmnJ5np198/UwMdHsxDoKGtenYzLiktCMICpyPa7TaA4LawhQ1qD/yCZlT29y4D
M3GFF+FRMBBiNfS8LyrDzOacvt1iMe4aX9V4Mw1gilnqpbz+uAT55w79b7+57R6P
TZF1Oyic4zr0GoQRU/G4tM46pwEdv1RX6wNTs+aCp2xRUjCzvNQCunP0LkWxnXZG
zi8p8qwY248xMtb+vPY6Tw0O4UNNrddRG+Vbcefl4fZRyxJtr28ignQUvAX2oQIC
3y9fGBjvzhXfWWodZkEG997BWZjXA0OXZyLj99zQLMZVVmooPQ8GxgiVMXgzz7Zy
EzF1Q1oJT7W8sUwdDUmHpPbaVB/TRFBPl90CtC0O1VYIfGOLkvn7M0lvIzxkd68e
r0pHX7f1aJKyP0xXcunnRxMrtkrt76iEXI13mgTsc4kWBZZ4kmj12gMat+MPal2t
SueGp/4igU4Y+xlD6URZLnU6uypfsQ6SmIQ+s9AcTlGaPwVs3o2ld5ILDpImd4qd
kaXTK4DevT3SPUVXtZ+MlYB+ydljOPaoe6GD5YucN6mou7ZLhf0/ePy6Gf2Tliwz
Uz4Smon3pF9gxb0S0ILr/zMOebnLNOBgIqb41NYfcCe1PHYybkWNM6KcmWV5RVVJ
3Se+dMtMvoG01M9JMnVRxMwqQ2Qg8cV7YwLe6pNbE+Zbwo4mFoZHpPpc+HOVvlpx
OTm5V+YOqXcjBrzVHubWoTDzIg2xW/fkob0D5kPqeugk6nDMwa+/MAs1rzCQYq0u
+Ag8aO58+1POkjohOcIwgcdPfKOe38/T4zXaUd+WLr/cCkrisrN/ily8Cj34Qrw2
0gJ02/ZZ45NOuj/titg3aUnKSXyzpIEggPH/5fJJN5xoOotrpSjjRUzzKj579lAX
ljl6vAM3IHye/GvCOMWBPPzDaJ1YuXNseS082Vi6urns+r6wIOWPt/shUfu2Ygm7
l0WWfqv5dbrnHPqw6EthPCvJ4QfXLgzTYbPArNRk1dtn0u7xCilYh7EZdkae+10Y
td2HpqzEfwfCWHYOOk5umTZ09s32lG373hpPg2JChvE/+om4ztfErRwWNTrwinGl
FnfpiI6wta5nvgqeY/ROqhkpBbiadvAc/XxJvtMbCX2zx2YbD88H4uUAY5FE871A
vN6QvIF/nkq9SKOmbzINsTvEArsrhuyHCaoGcptc/6IMYxEFIVIiKUCgAC7LOI1U
4jZDpnd+k5f8+8qH0msV1pj2UjrFWZmrPlK9y3SIoyjdYZt8LlXvWUJKqd8lp7bG
/a17F0Mp367+TOXIMYL/tCu1w6bZo6bXHPdE97ziI9Ud0fHMjdq+YzjcCW5aX4S6
YJ5U9KhBlH8524Jxz2LijO0Es2yqULozMxWMCn4wqZGyhnqKfmnAXTz+pMATIhNS
UXIYn1QiMZ3/npIFJ/yuQtX1XK88n4MUmLlIxfnxFuxv1+5b9RDpRNW97ZAkDoSD
/KwNq0eJOH8oYxMGcnMMfY4ZFr9EaFaFkAmjen1daErstCKUh0vga1qo8B2WbjL2
u6VQeE7b4DaTUQrvY/GBNlMZqw0FJUvhwzpS/iziuCxyrz6pLJSPWdOtEGkshEms
Ds5qUSUa5PBdc4S/wzpFF1jdFA5RBLGwUG68KHjYac1gw9g0Luxubpty8TV6Wo0x
jxJaeZJR//Dckk9T1ENp+av5Y5SQKAszu93MXDQy6JioTvbh5OQvu4NiH6a8HHoy
lWPE5nQNYTGe/e8fmtvl3fQTtET1p77JkZStEXe0FGlSCZXq05rcyfhp3gE9sj+U
pmwcr4+NOwfe0449he3sUCeY5aHDSujf/eviNCxbRX+x0tpckt4mWsS9HfCl4rWS
HYvN79vETPeltWe5s2PUcW4W4SQCu3U3eZ0za7KpHx3AyS2obH2jV3f7yzo9sO39
5u2TIFJ67/U/oPOI+/Og68IunS7720nAqecOb1ZHyESO5yJp6f2Bb3EPQkVmwUk0
9AB4cMNQr0R86wIZxXyaTBfmxbjKBPFnLeGblqMl/fBW2ERyeiPAllP0U+XPKItR
eZaLJSRhwn8WLldn4sCGZ875fs3Npo0pPSiMMaPmSIEMzFUCvwXdcxDegOSW2frF
ltZI1C29mH4QzLltnVDpWAbI1KgKyqpE+QJumIeOy9W1j5Fn8ldpgs+JtEjH7UQI
76WRoU6BTKZepQb34ORJgIi3N3wf6WnhDrr7WdEONLwXUERP3uUBWlNtWKEfyrap
JBDlW/uDQHj8X1jSkqyp41Bk3k+A3ai7Orb3kMyxI+HI69nMvP3X1WlhGIbzI5lU
wDsVHJdr79WR0SBr7FiwUSApc5wLRd6iQntr/Uu5+kARrYWHT5gYKkfR6CyLjVV/
8A6MSWRD4hr6wS18OaqRgzmkqZ5DkHPd7b01hVud5NDrDWH056pdbWTvqc4VtgkD
x8zn9LBB8mnqcm2Y8ahUm/eR+jLKyuZ9AGCnkcbK/qHKaCj1be9N7ggbsX4lpnS8
JyOd4gg+ccec1uz9T6UghQc9c/XoldZ+xBSDTuHTG18DHTWh7ZdDKRmyDD0OU5up
k4ehKJL6JSWSW+Lvu7MhLS6p3R87nYADdLDh1/skcsukjgNdGXksWHzoWuM4IZFK
QsB1GuispHAg5eEc0iD6E/oTy8AZlMaYkkKMAQt0iVM0YPaJ/QF7uWd/rH5gfjp9
za+Gec+cLHMHQwdaciPCKLjAosiJRaBwyVSxychChi8fgdOVp40iK396JYfvANaD
qAZdtVC4p1QA/gNaKqx+AUkBfF/Tn8PR2voBh3V+RUYJhcVzraPNjV6zTGBo4N4i
54+ER27b+BW1/Y7tOgZR/QAi8QqjIdvjNCVEU2okWnmsqjQOieSzzIpkpaRB4HpL
44Opj+kdL33GEKJ7WPRio7pt9vlUz238teWmoZmerBVMjtW7ME39k4l9imkWyu5G
MJDD7jTZK/dq0rhHRM2LHOh9cOh/J6s9QaoLcjTLdzjGoL+jJ7BN0lsclMG6a5Lj
wcGz8naEJnc67zKZ0ysr1YPr5KnHWT7E6EuN39+85UwN6WW3lXe4gIfrqFOsYU6t
TqqlV5CLA70yxgV7tVUvn9h66QGo+G88Sdpkym/Hximd7Vyonq0U7xURxvuitC2V
Jc/wSbH37zw7fQYNc6B3tekmCuyoBImaiRq58uUOLP438NAfAvtmDKP3SiuhyR0R
QSYTNW4QJgiSBV5Y6A4Xwi3DkeW+z36tfahf5rzvliHC3Sg0VW8iwLN+0H/VXgpL
x1smNgfTf8HJY1dtHdnRCs0DsPvs8QoXqYIGSdrW6CIHimS/DEbGXs4UASIq/I9+
dd0zaBI6ATLlzTdYt9UO8BB/p1YTI+9m3tIp0IhEPzYy0NafgHNMXcLKtBs/3ITM
UhsuEy5+04sIOJpVt9fJbbUVqV+YOVouBR3sBpFkqCP1H6L9Yw+ZWuK/GKeBpDiH
oUyYAmqqbAE+Ss8zZ+QyP8UbJPmF6oNB6V4n0AGqkUlnJuOPxaMfAr4tiWaJWJ9R
0zxdq+uTWhAge/XC/GFGmWWsu429OGHTMEmXwfkbkY3wFHKIza9v9nBUV0h+1IFD
mb/yh9LLj8gwcaB9y1RmE3LBxiyhgRJoJTqGOccvBVCVRnFLQozCWm4ubD7yVk0P
/wEdLC/nnPpgZTfKU0gHPD4GWw3gdotVVCfC+c0AK4R4guee+QK/dAet8PLg5Fai
JJ8tntew/bAvKOB85s2vKDVo0sRO47Y1JLbFwGO4cYX0/NDLL94fdykEebM5Eizo
Ie4fkhU5yRQUkBcIlvQy0wl7bZQEyOSYDxlDbz6JmH8=
`protect END_PROTECTED
