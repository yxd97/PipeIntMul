`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iV+jXQ4CsS/k52kRmGQ91R2s3+BaV8Xxm7o2lGyp+I8H2F0+gGW0r2L/sp1oqhxC
pwox5jQ0vs9predkxTPsom/uF1i+2iW3gcdQLbKljVccPr4qV/z/BfGu56cqAMaE
hOMcteZgHabG9WPf0PxdULJEmsXIZPO7xQTY4MSGM7IvTG6LINY80lnjHq4Xygg5
I3gmLTCI1/XC6v5NA2qWDyfGe3fyB6L2UdROBuB5hZisxWK+6U5IQZwXCKV0j5B1
wE6yGqy7BYF2wA3Oflsd/lKuBJoaqa8Gblqd8gXHg7DLdk6TXsJ8XHKHKVFyqN6u
sURQIp4ruP8ZqVNgHM2CAuowQiD65JTrJ6zS1sE5ArPTyVmFmONczPfxeQ2Deu84
fR3LFPr444M659XWa6O/jfZBzV+FwFctw2bSCjBCPa2Wm2yRmUYoiZSMwNNK6OfU
Cb9wJhL5zgf8Hc+AsYdWFu2Vk/ulBNYlKoBUCs3JQmzQa2mLL+ykvvUA480zdovR
vr6Vq6G216QJtEZU3ntqdd44EBCVSVOc/e8omjTPpZDlNqnuiTqBNJPaBRRzQsaT
6BWH9FKCoiSzpzSdVIXjBG1bhS7JNHKDN9NOxN70C58eMWOjT2NL2tzZnhduWNiu
V/JWUrfcO2F15fsMmST26cNFGRs8sbSP7DRBo+t/f/mnSjGkO60d+LMGJoIl/11P
vCTFkaGDRzy4himh0Zjv3rkyaoi1xb5spoRyrkxlLvQe2WhH13oycmVYaO6YLVJU
D5vYNV+wnW0bxdSuPiMqu5SEUJeb3ysU0ty4a1Jhi+BdTd5J0Lprx0rqyTgoJNz8
xdRzTDg0Ks3ffu8kgiprOqq+WqiFcHxFYNOMvP54Neco0F+8vgkAIMegzjXcsWSu
qTnchZSDlJEtTb8kdzgaOQeWKO/yBZvuADvDTr7b9cZAPO7yFQNs2QNdsvMEQg27
75n4IpH5eoZ+MRXEBeTNdrfLn2x6wqrD7wKFBXHv8aX/ZTxPGq/NYR0vXej3le3J
`protect END_PROTECTED
