`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMKYXiYzXgL3jp6IrlhkbUMzXvkIfToy4821QM9GbL6SIx2ZODSUziyx7oMh1xEW
W+UVw1EPTobEgrBX0ZysOSMix69Gn77kAoIp5K1UpNGeDq2Co1CrDIYmVLrn9BzL
QQ6y6n5+Y0QnDVqgGMj/b95DuGPAhM40ScIkTyAhetOEU43LTI5uZBGy4Amsjkip
LQJvHh4LAEoDoMZxhHpGDBI3J+q7j+cUq4UJJE+Er0OLMH1eWV1Dvup5iwiJHWGV
9S8XNgTWO69U/6m7KcXFFt+e5aUCzd5m2Cw4WknvAV4ZV8PtFE3ESId+mzMF5d4k
JJTy2dXdumxdaX0MGZR67IEJjGDzyL0VJGvbGtCaIUSoz/l1VGvZzK5AprnivVn+
OtvYS8fBCnp0rN3FVJ+PB/UkQJyLRU9ea5U96u+wdSE=
`protect END_PROTECTED
