`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6r8NfzzBQM08sgK9oFhqD4uD6LLwcF11rQ8TZUrBbmnMAB4ruwSNqI2dQjWdqfi9
KMGN0fiUtU3bnlIVOhJ5HW/wDqfi9sdVlGDEMrfai6bniYYW6wc3TPc82CmcuYLk
51Or7/X5uh28kpyyEyWuUdeTJOd3LLy4Q8XF9WxtxVMOMbjX1YsaAuxaGmQyyyJG
vu1I+noT9vw+LXYdle2HXknp7OHg5FHKfXD6Pe1uoCaOS3kOnejTLL0QjshP2nrE
sXooOGbeXhPGEV0EuPzb2ji8SBDhDmkESzsPv+FI1so=
`protect END_PROTECTED
