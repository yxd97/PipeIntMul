`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AUOTu7u0PyBsGpPMRFvtaPKuNL3BEHC05x86ABDJpui1Zv/2Uqtni5cg5ak66xPW
1N7MHS8h2Ek/LtfWki0qrSVf/Nqao/VfE+kgmiJh2tNNiLJnC7Qq6NJcir5dEaVz
pyknL+n4ylLCJP425BLhMRZDcP+iKLx/6ndK383QHn+J/kc4PKbTIWw27VM7sOha
20l3En4czUK7OdJ4Js7EL6KJh2YdAxSvww566SEzqKb6skaZnRnt+IDUG4r1nyVH
jYV13UB+W5yGu3602sXmdjbRUODjQEuxlcTQoiaTojupdNNVBBPOpMORZGmUekAz
4WmHtJ7byFJyTzKShjH9Iw==
`protect END_PROTECTED
