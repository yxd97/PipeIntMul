`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N54zGRMx4rt8XPAjLfBRjLTAB/7M6ZP/Bhg+Kaa/YSly4QglE2+uBaM7/gkItmof
jzeIENp7QtaGRP+Jyc2LUhaw22vlvs37Cx+BUFysnK/IlxZ71A2FQtfQJXpcJKuS
m7s5pQv/8XxWgfmyiXPBUyZgCAycim/0OzSaO1gkdH+ZIoV+8ZsPhfItOWm2Atb0
9HXrKRhczE/lRtbKroYekDGaUdA0NfkzoJFADxWwTFyQaDPGjGHHp1HcpwOd4yp7
3pU+bPZqQ9IFR5EZo5J3XuoJcTbzLEaiK9d2zs1J4KOU9+uIP2gsYR4/ToDOw7Wn
pETUAOdPyNQqICmqu3nv0Q==
`protect END_PROTECTED
