`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1b5WJeV0fpP48wHGf3eZVmqHMrXSAMWVa9KzNpHMVRfKkDzLmlY1wJFCPyqyOct
jXIrwyex2n+Lqhupac+Tgtlghy4NCTkhDtdtqE0KIa3nyqsO+lA4VZSHLUa7fGK/
uU1KqDylZh+PMtx9eluBIWfOyXymKFZFU4BxAMRvgS835AtcBCqdKFtNMnexq28N
mZjiwHgGSZCuS0OCpg4YvW745sVXAAnYrvuPQm8rnvbQEahp0N/09i2DxJaspV4A
1iwBhPZaIH7QFZrZCrF2h/3ftpMJmfvSuSxm9GoyqV0=
`protect END_PROTECTED
