`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F7b1RQFIw4/zYrrrYMg5PxCNJlOdP+j58YYTgz+YpXgF1rMtySNw8l22TOBCSxYC
DKUcvdyqzcbQbShWaRZ47I59Uu7OAHPQGhhaobY6MwfwM2MrKC5cD2pzcYEppueO
fL1A+BG57uNoU+tdUtye6LZXdawmdy+sFP9ogLa6Rf19FU4t97fX1pRpGl88XNZn
5hW4DlAFzGBJpVbgJrIa+k03s4UDPP6+5yKmBT9NKtl7N3/3ToFd+xOKnyzOftk+
iFUV21IVS9SD7Bkvka3tQCCcwm+BHAPRY/fFTnV0BtVkreXjaoKrHggp7MvGVvYi
9+BAv2AqKc+lOrwlQilsROwNx593dyd7nmkgKorgwIsKYLwGpNr6BihHoDGFud9b
2qycA2zBk78a3yc8dR6u/mLuWQLESNgAPnu9VJt5GIxgjdLq0r7e5mxP06fL3jPO
7kaRF+ydlw9VuK6setDsQo7LRCH5x0rWgltTlA9nV20OJajwXwRzCHFo/Q4UvZ47
duuYJuqLiWSOTGhuCuoxt9w/AScn93Ri1o7Gkg2zoqo9Asc8dggktpRJ3BC+c+IM
7hQ/yS0kxRrXe7u5cBycDyT0RGOiyBCONPUQEzWlTux+yefDyrgHYDZ5/+IRF0X/
OjX11vp+lFNN0TvBbU+uLkrivQFhzIJzysl1PPRLsOPuinUSc0fQApaGh4+jMnxM
FM/9jNgzbNHBAMwgB9mq6ZGnQfTiQtS2vQIEQ+afKQpeBaHLeAKTu1gVPiYyMFCI
V7ZF5vAFwOvQsWB4ClftnzZeMEjTK7P65URSAc5SspE=
`protect END_PROTECTED
