`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
02sUmDxBk8KsAdbR/Xuho/CzXx0o9rCl2BuoCg+5DwajE5uC+Mx7qOZOb5J3fJlB
+hDPIF94Z8MBnDU7w+/HRACGRI/hjmIKvDUp5ridtqlbFL2JuzahECeouTTXcK0r
64eJjkvNDrX/hWwjV/7y89QOnMslsSKYLzFEF9mOEn8KsIWcuF7Oli5byfD2/6RU
GrQZYBfmw8Pylb40OyNZB5ZXP9ltiUcu2iVKAuPfmf8+bnFD/jSqijdSglhfmzTJ
`protect END_PROTECTED
