`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JNo4xwt7X9PPX18ofl5iRsF4LWfPyIJZlxEuNXiGUETlrCjkWrMCmblIDYUmE4dh
uGxrCY1KxUZKGksmqusjftPetYtp0EZ6k1UnHBPG1lAbytnLGGulR036XSZXo42g
tUxKScWKyr0VEBEaKZmEDuQSpBVEi2xdKXJftV4xXtT4Ye4iH71GvntXtAN7tfwq
U3JLtra6RDrLJz1rcMWIAFwnaVCi8JAgkG0zvhs/urYamdDrDOtSoM6m5tLB5I59
p+yAoiIRVlCib7orH8/VmkBa4JsER+P7xLD/VccPvl52pP0I7M9EzppgFUojsrIy
wxbOnI4isBWzGl0yALyyrYqeYtrLJkINXAzH33hYjBt1yem9voEkAy1K1tUzzeHN
B1u6+ZS0nXNeXOVG7c3Qc1JTdCkHBxzNaSlJKxxOM+DwEjuzzji1TYC3j7AnbZW/
cqXIKcxTZl9mwmBYJNc/0SUn0cx+2k0irD2oxEYx0kI5AmNl6xuOqIbtD/RnRyOm
Mb/yrMx0IRgqbwc5fUVRe7PBWt+XdPI6L0KxbTQ5Oz5Zu+lzu0Zxn4hQnvsMKqYv
49sKfExG0l+n9KV0Hv/MqHQR/eVvYL3O+njQvoVSROui6WXnRLLONcHcKrsEEo59
TpvqxdNneSLLInNV59sqEdM0m7k3Cv1IY7BmxnTWZ9nUHISVo+uUQiSZD89ji5CR
9U7HebYgdzhCq6ikozyrj4jfLgOL9qFNSbGP73GALegOQYvwwII3kka01Uv2h06t
grFEOWTBKZVnLeeFp0LR3NOW/ibbq2GooKjjz5tpcQFknGRKD96TWrmnzwXIBXuE
hb7h6XpArCaZpR2ZBU/FS4xtssC26dmGEv8urCvl2V4CohM3Mwo8M3NpKn83Tz80
GUHsiY423OdcRGznwxmdRhn9uWXUYU49qsmSOPGSfD0pTtS6hWNtWTp0vd/NfwMG
dbz1j/vumCtTpEJgWaQk2sPiBRmmE/MUUlKaTqKWubvrQmTpzJLdYXVXS7nILQ/+
P7ELsD/C2SRqpHoDppRqkICjaftFnm/hR/fbq7d8tJvTgrFT7tHDu1uPMR9sZa6e
iLet3+JwOBy4xOFOi6NyABvTjZV3PKYs+E7Ff+v6u2xxWJ7EBAElnD/MQZrVPqYc
cwVGeCezSQ3dfifk/BVW/7WBXu4LrVsEE18z0fSFoMNCkVmLz/+Z5HJfIkHTvZNq
JFEC0ATp+NvqbewvbT05BsZ9K7BP8zK1vkoeH5Fntsd/66AVjY5/yhFFI5IPZ0rU
AJel0Mi21g3sxptyrOMpdN/K/iDgK9hIJLJ5HQmHd1X9SE7uc7vIRO8wvlgqySUo
Y9gk5TpzkVtjMw4/6ef74xVBTPJB5PG1dh8e1GtpNVhASHR9MHcTsnybANMvZaiF
SZ82wcQcoAd8F8NFECMHuo8J3UrrG4Wl9lfjbExZbeuSeyR0dsBOxQo3ZBdo97Gt
87AfogKYFSazCRXdgbTYqiNv+Ks9o541GlIS6JNQAe8c/v9ChfCSiObMjtJh890S
KneBOm2tFEuZ/QkfUxh2A9PEj0DEpuwOBPuvbWq2pjnxTxX8Q03KPhelsNW24TXs
GSjKCsBfcwrHDXtK5pfqQeIhkg7Io4BDdx40HvV8qoBx6FtPqUXDV31Yk8XEQkei
HNyhPu85iZC4l/ryC3gAKnl2WWunsiR+yKpJGxFbL6QdEY2z3dyqnZw8oiOFlIkL
K9JHQPZ117o9KeW5dt+iAoO8XFcU+/2bHGSK0NyzIECkvEActOgrqN979ChX1Hox
4uQE+2nNvm29r8SLx7puRqFh2kcDbOD0mEYxZNWgoDaW0yrVhMz2q1qcSA5rNgts
zy7SPxMYi5TpR5G+UCt1Dly07QL2TN6gOEhHun/KmoAaEs5W2VWJlk6acemjLDDZ
Qu/26IQxNoQ6gT0VmDVoZd2zvzcW1vOrH2GXfiVZrMhcqNQlxqDveF+VgVvOysHj
v45H/9vzME8Vy3z/NTwZl6g9J1QR25wJt3HGrVWoBw9zLO4Uj+mi3C6epEcUMLZH
5XGJ8kBzQin2uAsIZMq38Ugf+FpNOtzvOeY8/goLjfXWH7OL+JaFRCQbIKD4yd4o
Xxn9IxHhPPzNLpqPuDSbojEXpRrEPVaQ2IcrQJlhOG9C7UpgL1Vwwp2nyLCqd1Fh
elhgiPVc/3korVZ+Ycse75d30C/XBf7CrEf4LUTxJNuO/622F5mOmv15MW6KEykU
AwOoeLFv7ifRS2AgMrCJuXk3LGe0qAARY5m3rc72n35TU5RQxFJOK4Hkvxeojf7D
cp/wnq0ofA6GKc1VBdw6C/xzy8pYHF1DWGow1sT4e2oioAgrIz+gbpa8XF4/7dF2
VE65ZaTI6kLKA9eWlquZKJ4Lu7qi/NP8Jt0MFs8Xme3gFOWwlnoK+zC4DMePSjYx
iP7w/aTHkI3YpfCg6ToPWuMO5k4B1su2sPJobvS8yaoM+j1vIwaD24Wb2LemSwYQ
S1GBUnMsMkpx13FJavXKSbd/KZ7+HyRAQVaKHVL7ccJpEYkyyRZpE7LDqraE1ekf
Ynu4pnalOSwXNxwoADpMErSGQfo9jxMjq7forNObXXv4fXOtOQ7eLp4/dfrIVjPf
hs6RQW0v7BzMd4G7on57/0ypG0Jzd58cnJPEr0KpnObvcIn0lja2t92mIRmVjHIY
5bbsx1sDw1yBx93dR+trEgIbtXoWfmWTASy9MmzoFP3d9w8D1FS9bcx+dn1jhnMC
+Vfpr2V/Hfplh9Tw3B4rz3aatS3RzLAmWkeHA/fzY1TTUjly6tMU8GIIHBECTeRP
fYcxzrwcbFbwTGNuqkhV9PzkIIIpPvXLQ9qkf/YnkgjnouALuXVV6RRG3DP2UgiB
i3EINrS70hERM6sxwAwYShNHpqhIeTcnf2NAeU5TPiiIsEwOK+EQ8Vv4S9E0s/Q0
F2uu/iPQU/Vz316ni0lS+W34TZUi1eUBqcsh6dh2MsClGKax53gyi78onfVipskf
j7fwhKUmcn/V5+fPf7jPaZL1TwuYdpAwRqTQRtMTqeyL84UtXeIq4s889FZyBxhN
EwbfKSOf18ucPDlrDeTDvvftjGMt7VpQqamLX6QYyg4utvWcL8CDGoUc9GjcaVvk
oVMW+9V73vzDlVWKhcGlgD585EAawBvpOws7W91yDDjRPsWRZrvUtp5dUZ3gM+8q
FntWNXLpXZSrTDXK3gFA9lnYuwftcK1/Es/nF9pvLP1Z4OdxFq+TOUsBmwzL1lEM
KF81jQ1nrI6R3sbtX0snz0E29qPI64OjI4ha+UE56qtaz2ZaD6r9wUvy9IcDgOL1
S5eEjpKOXpjgN+gWKl9NYVChnsbzEiTcTBgFZEn8EG5S1YqYXBQSE9ladp/P34bE
FgzBFm3x1ICWeNxEvGHSMdT6oAwtwEV4RWOD391Gv8E4sV9WLBap/jKnbLE0X08R
wHMV0hoMoT+h52zrw5gGCCh3tElDeBQcR7Fh5/fxg0q+sXQSD9QcFv4dZGF9YwpB
yAdwzVgt/iBq8yoJKYQWS7IbqssWrDwZIEhA4XDy54mtykvbZ+kNQim5q8lUDYrK
bb3rpaKcNcPno9QC5cVEmyZG1sgO3/2vc8e25R576D1MOM9qYaLrNaeYnXz8D6Lw
HlCorouw4kY7jEA9d3K/vyo20af52trvy9s4PDcF0U2XxagYAO+xOqztup+X37z8
pzEIvrOabjRWYGN7q0ZnNZajOyWhrAeRR3m2V/+0dYzTCiPe6NPh9len9JxROh50
oenJzeL8UuMAbPL6Gw/7DYBLsjOP7Ocd2/yQ4L21r0xNg89h2JY49bccUJ19c5E2
1vBwFLSDb++tkGZv54Jc+9OLNPO+IrOwhaX8Hk0c3eH+nn2szWvk68jj0tfDL09i
80/JXF1OppVDoRDIkApkTl0bMhHgnX/Ik/F3dAhMQfnnmbf6ijpwqOoGGB0M0q4v
MWBFL/gXvIMYIxVk0CcJN7AqCPXEPpwHL3L8vtKB13wT2vcnTrPUaMucjcsl8Phf
qMFe1Dr7Rifc5F/wveEdE9QZJt8vVKMPxVWfGzS+/U95AM+B4ULA210lRcn3v4XG
kPoYmxLqKG2iHTNj1Yvv/VssToh2AvzZ+cCSBwu3PBIOUONoSemVwcuOF27gJjbK
OmBIPdok4wVD8YeC88RC3UQYMr6v1iXdtOuLsP/oD7Hym373PLQCTbTqK55sRrvO
0msV0LAcWu8Hj/nbA8Ya6zLMiezSZ0tCMBy6wS+4YSetz3JqgkHSz0lXwN0nfEwi
OY5t7H4KMio1v/p1zxdM9zP+oczdmHQbvv97SLv7qSodIhHSDKQjcCxj+UrwsFXV
YtMCSzBib5xMP7zXRhkS33xt9qx5yOue7jtp7/ss8ip9eMI8Hutd1SdYiYGuLoea
EoHgrk8z4BhW1v8rSjvtR+URT0mxN2VyVSm7bMWtHmvhhW4E7oDtS9Sj6CsaoP/c
bLNRabCwOALu2gV2gqh0p6vrt9bXw5OS8ZDGPs1jF3ayJGtnwApN3Bx/arl5UCML
iNn9M1q0vZkVDtTAOO+rUGy4inlDkXzddNqYY7GjUC/vk/RLuL7NRYRJ+0a+7gac
08/ABULogT8w4QVtdNqMEK9Tq4S0XXjVTKr46GeUO3o9MeMqgnXo2GKQikefJ6s6
ThMeZVWrnhxaX2zLgSbSZxV50q6wK3TKvvKF4h9GF/9K23tI+G55zitaDMcuP6FW
NkSGTJvCfzalYIbj9RGdToF6O0Wzz8jFWtw58JOFQ0XIZqOe6gJf/cOUjAl9fBpn
C07rsmg2GIIGTw4QG5ctNDSijtuVHywFQtfwOJKaTYX+RlXBQwOQ+PkgVj61YYkw
pvYGr4WXgzIXbOlzkqfCY8Ik1JJ6v7bQh0LE38WiicJZWhG7VVC9Az4Ircj8L2HH
XEzVURVUF8JEbcYQ/J2bOv1zDLpWr7V3WnNMqfipGyAlNe80DFPuUlRf4UvbnePB
EbmacvkSmM/QuDHOiNMBWhrRF/BMTTJG6Ki0Bx1o3wyl3RLZ0K87QND5T49oSW9o
lcERnT6MLupaBy46Au5cYQMS9lMiR0zjaH5vI7jPOvcSI+a7jYKAfvchEEw1WOnQ
qER7/ajyZK/23vY3y6m3YOlrMs4N6ApJkftchg5fjRc4sELCZ7FoqTuno4vvNJzL
tbZ69zi9L1SBwriVpHeMpMsgM9Pd0J56yNEa4u5ylY3S0mGNYD73kyPPXIJzZZx6
lTBCWjWKoHel42CBfl4DvT8cT4E4qWWFFCCBh1jF+8JzS5gOQuEJc1p78gcULWuF
jKqz//CwpSy59BhTQCxpPxkWiMooihOzY+JdSUSaowGt+XCTc3c1UtlshmBSYyvq
/pr4q2/XH7WHxOmwgW0GF1X2WQ+2XYmkJRYp9MkWm1sM3RcIUfvgpyKQpYRb1qGC
a/JWYjrMicBhvo9hM3DNZmBx63G2n77QjhTEMdfC0sCDZSTjdW1SiHQEPU0swx1B
EYJ3dk3nUvEHZRQcIjOvM7nXiJuFGcncx29rAlVoXFxnNlZxbHh4LDlc75Ko9JVp
a7FT0srZxjDjZB4hKNFOXuDWmzwNczD+HO7bcF6ZA4Bf5HoX2hDonqzaWNm/2SYr
niIwD1igBGp37jeWYZx32gp+OTpVcjVDtr63q/ok4Pd0sY3hhnS0GLor7pQrptUj
hfO/uIToknhy3CJKGeNrdlN0lEyG1BBRFVUSoqp6hgHtFpCYHJuRR3j7OgLPl2+y
Pj867tVT17VjEPEwnIOuIxzrq4V7ybvRiudeyvVdhOBaTJrvrSI3H7tBDUXGmXEF
5ew+QqHZ+ooPPPzyDPz0vPTJkq7PTO0yCmBJLVOO+bSAK6o9f2+0uPzlJY1pUkwy
QKZlYj/UHWGK+7gVf3yO8J5UycksjcAWXZy35foo1ui90z+hBmyVTeVFjKl9uWGU
rF0/VHcgaVto/bTfi5tGM4GP8e14aPTEHFvwbvOaYwxDFEL6oavOEF9cbIVBZkCW
5PT74+LI71bJSr3KjHych+9JKN/vv+2nycqDRbnMI3ypgxzn3rDwVTLucnmTQItl
tSNhCTtg1enxWkBxfPQ00qWOXqMuFYdCT7mFv5xZvOa028rT9ocn2NIEmk8Qebuv
00m66HKwKL6M5b0VN8ScbxVbMsAibjPfs1XTtKmFJJ7pXnJNgO0jmSOGgP0hmuBK
eF8tUeQSpyxlD7gSPuCc9gswlUTUddm6B5fwpD5wkbP3MM0SrAUN5EigIIte4X5e
w78d+1xrPHCH9w+f2z/sr0oS/f8VcvOVlDaCY7qeWa3ZNNGlm3DUA+B1m2/kh+4C
JvGlfDtxa41n12J/aAGyxdPeBuk0mMTdCWG1vH5QKj5Dl0j4ZkQl2+Qhz4kq6KXX
8Ze7Yh+QzsNDF8LKKWQKjRcjggO2HxuwZifd1KTo1apVPxESBb/htOZQ1m3hqCtN
3raVwBS3tA7vtTAe8hbhXPQpouaOGgKcQrlYLWoCXyBVd8zJg/E4wcxmIY+FziOb
R9L5t3D16zmch/QwROAZiZgz5Dh9KG3DjNm++HAEg8WXwIGQ9fP8Nfb5+zQrwwUd
LjCjSCbL97rSpQQEDVL806/4ENB800M2spos1zX2IqipMJhIYU81aDuYQyHI1qjW
IIloeySq3K27p2lwsgfmSCima7m03PuNWBt5RH7rSpxQBjM6OGjaBSA3l5b5HiZK
m6MxQaE9zzX0PmDD4FnFlf+sitRlO4194qsHg5SnKVHJuFAf9sNzHiZbwkxpP2DH
uvwotaBUvgRsm77Nr5DXoGFsQ3Cbpf1EDZr3nzUmcinS1yvaqW85dRjQsAQIlIOV
al4O3tckA6qSTAzO0VSa1EjN77VPJbN9whQ9kRRDIfRL/G5AUBVMl+ScqxZEEgMO
B4H0zbNhF96mPfYt4tbfEhR5XT5G+aF+UThcyAwDdBTzL9Gmz/qIyGbfOCCLV1hE
e4yH8lxOM/Ux659jBhLBr9pcnJZuCRUQxSimRnEtkrSXjErJaFrTiK9V8IeWlcA1
TGmgAnRjPYFNKcaJ6qylBaErVrae/lDmAfVviNw2MsT6QPJCmS/9ZnLmt7olSWMf
ILP90QZ+dXITnFBeubsFis5boLsSbL1fCCuw2uywJ+YHQB0p/sK0NuZmWdhF7FK/
qakZA/Qd/V9uI0rDLSML1bg7xPXRjsOD2LRHyr4DMKiDqzIQWxyX7/1jwup4rOIH
cne/uVo7fA/wYpLEaNYz9RLBgpwJXG/u7a+JtaHXKAxG/kvuTQrIgjtH+WhTWdWZ
nMUAvktTT2pyp21b+ix85yhIPtNvAX5LWpvdPjmJrq5KTA6QzbojLZCugHZuwF4T
xTpfdd/2aGFnUWVTCp10823uD9HHmIgdJBgHqkHAn3lvODzDw4gIxy+zYPCMFG8m
na7RRufQ826w4SFLxJ7mgLgdx9GJ/xcXx3X5ki2QIqmLDkZCCdZYo9hTN8vtQ0eU
yZDObh0c5WENT4cFpR1CBzuCFPPe7Gt0CrIFe1QQDchRTyxxaqN7VG4ud1X8bgOm
VZTPos3tzTMjwgWuUegjq/mocM6O63tccvkTLX1LVoke36AGjuQOPWQD3kvdjZaE
AvdI2L+6IRVsBRWJ5KkRecJg5DvKyXN6N04HBJ3Qdc1UfjQTb6xcpBc1UIhylzUk
mkdWiZPDpvG5LvQg2ROw12DRMChJxbxCC6x3q4KxpjIcFnytaougZOhUbKWuUuHD
WqQ8w/MokyJDiIgrPeUaX/w7H6uNwOjYo+1tvQeaKzH/WnFWJVqEJJPnZUJ4Vtu4
m0MpmLsPXAg6BkVvwYUB1OtOg2ycyBApCYvtnN/HUGdq8icDIIQNr6bkqky6GaE0
T9/XPKpYM1OWgEdLmG2j6nCvOrc324NleZx9Ed0EYlPwLqHHbRoKOmMn0Iru+QgM
32f6yjRR4xb8fHp4pimXFR8/0fQ6fkRWYRcd/1aaVksVH5pIHr2I3iNHaqGYzo2k
193VVU5Zg02YwZy3HuYiLvAnJjl/jTjnzow5cnKSC2xpZ/U8wQMQrYU+w5vDHLkA
AGMP4lJUPkntuV9VG1Lu2vIp4kEOvhTKDjSTFvxpCF8Qh7sMqqNivx/X17cAmTnC
Xh4TSxObw8GoAMUynKCF5+TQsCn0RjSxG99IYL7/wWD5lsvd/Bw1+ZBZtFi1bx/q
MG3lLP2mM0GsOqmFksMVeS85xX28kyXwgqCW8bTZAWCd/+0M/O5Qq1pfriwB8N7V
wQEl4h6YV90Uh5ZIXxN2344H1yfhEYSnCOE1NnhgM1CJ3PDEf+PpeAIQC27bcNcN
ipgOXZFATbxwq+owZNDmy588LHn0EpRrqcrgmxgkJXkRCtsOLgxDI7MkZTQf9n6r
gduJ29tYN+nLlXgMs+zXtpZEbGmiRj5qHHkGb/C2rC1AjUlpRUYaL1qOvJehKOaa
djElJvHzWSEw4lKebzLkedFBNa8EFacYCl/W36vMolr3vUwSP2TjkcHc5y8YM1NC
bG14ZSNtW7hyJKKIqaZlbAa3oBD+631HiPsoy4HqsnZ9mzcKEbqXxT0xttssMIaU
eSKxsDQ00J4sQQPzLdcL7S2PmoC1qVhl9hVqsKxCrGaw0QANJiCZRA5iwTt5BO/6
xd/becALr4KYWLQPBHDWV92mZDfksrMtYR2PJ9ajSCu6Anu2PIf06FSVzTSoRq39
omdyeivepda/ze+psLEAo2iBistS2bB3MjhQ+xetWfoYaxeWBGq7PaSLIdrmCjky
iS+BceVfk9KaeQ2Pr2J3pi0uK8sXub+vlR1GVysE1FTUoqkX/Yx2Ke2BZbbyCzNN
geScWOzm1LTZEwerZBJPf//wSjmjBeV/Whx3fH7uWvsOYkaiv6RERqZTzS8yxIxw
+ZXFMLOQQbdqDOjy3J22Wu+NXXGKxFho+X0ow38nQmwDZHf/d7Zvx9BdJz0LiDaR
`protect END_PROTECTED
