`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
es61dODQStEZY/DoysuZ8UwEepL4UrSp7SlH5BHxI33TObiVaxYIgrpu5RFnlZPq
uiL17JRHCmt3y1SZ3tRche3+667Hw6lp2kd30Q2gFPRnXn90Vp+SywB4vcwn9umu
GzVdtsMlyG2Y1rtyF+Zh7jFnuEfeuWLMv0gX08Mq2DNAqad3apOje/t0p5MQ94UZ
0JAnToBARbul9FcuoiC32JVL/zJiHYzHLDqGVF12oOLqF9RLgcVVtL2q49ukfc3g
V8YLxWg5ku0+fqLb9c/su2r6DyAqQ+w2vkLNr/Q4PpPj6UqKdAVJooN+FtcMM6R3
1TC8azpp8D2Szl3RZxkbQg==
`protect END_PROTECTED
