`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
25lQvsQ77OmRS4qk9/Hy/S+S38gFKtv7nejLGBchJLY5bDl0mAXJGtw/wzVxoNuu
35qArcAMh2CQx+ccbF5G8oumBrmV+p4mt2bu8MSykQkNAPBj5kdm6uWQbti959Q6
t7mZU4SSAGJLQ/ED4lwW0LznHywS5jHG2cPyOTpjeVml6BMVeSKBE/TkRGfAOG+6
sP+SoSSDkUbIgd8nCpKqzpFseVHf54O7ZRV7ppea9bSi2pddoR31VHMB7kr9acsh
O5SkBi7VoGjBH5GEKAnKpA==
`protect END_PROTECTED
