`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ipkeYA1rkovx8zNuG3FKMHhOk5tHBZ+j9TzS3EDFHXFuX+vRDUMBvpnX78WmqWUa
wgKfaxraCLG1HllVV9UwGQ0EbVBer7zKdyvtTLpXQjfwEd+L5FPQYxI5JFxtVAjI
+5HiMkab2IckJzJ4jwmKB6b0d9CL9deO6ezblDtD6wlixsbtMX2iPaLPdfynTPcd
crGd0XbXNl2a84v0sVX4ZKfYR1J5bFnMFpzangs4YosVGRVXiTLS5cw3Sh7EobQR
/omyTJ/2tx3MXnUngH1aEUU/aUN5/M+vsnsh7/7L+P4=
`protect END_PROTECTED
