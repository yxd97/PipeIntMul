`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vh63+LpPd2cxtMHYUwPM+L40sEPFzQ3ZE3oQked3GIKCF5EREvFpYNDVGuXRlPq0
3twSlQzRN6XpA6OMwyx3y8JHUxbLFzOQvWSEl/1PSk4DBeK6jw80O6I3DG5wLb6r
shQqvTX71SAfDxNKJhjM2qi77NSbit7WV9/KcqmQlmo7BG0tohSNwCGB7SJckQeg
puXZHO04gZK1zV0q6xco6Jv4q7LpwF11XMj5fYmxU8j2iUCeOcNfLcIL4ldnl39J
zO7TGcWMcu7dGWr2Y6VulYRfXBxH0Chvw5/eHzYQJp+M/tYdHnWKOB9m7c/e7j1p
eo86ESySF6vzaivMmP5lBy/OC5Uo4UYWAlAD1QobGHDRf0n6hwJxmvH3cUJp5Jr6
vl3eMPF9T67yGyD3uDFaynVSYQnCQX07btNq/R6IMz0Xh01loOptsropyTjs6TNk
sgWoji9XEGZ/5MyoFSM9KWsspYMnmJ+axGplhayYo+hFu8L9/4d4DXiLoFxmN8AP
mzdIXKxbAXLDQBn8mX3M9/NjQujWKH8159kZvpH1pn4/fRKG/4maFsIWX5exsT4p
GePX0+qye27CLR1XWNeDPPE8s4m48RNnP+2QXJBgV0pjHBQSo1pezsmnVkkLyZ3i
3a5ZyXdTaiTOatjPXVETKQ==
`protect END_PROTECTED
