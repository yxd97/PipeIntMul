`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jUtbaZuKkm9as8AemzwijKeDBZJYc/lKPa4PRGtL0O8a0yoif/AU/H/tD3gDeLP5
B0HE/yURbYOksoZOCl8Kbq+L9d0VV0uYrNDTkeSPXwHkdA2aHgsE3vi9H4Y6nvxx
qrMbrAvGdfLhMMytA0+bIvX7mLw95qsDCFSo4WiTPFFPJsb/Y7Tx7jlZQRiaBSwD
ExDxbOaAHV/f21Ye+SNL9Zf0cLXnGEXcGHOCYULrfGXP0vqck18iT7+Dn4L8Pojg
Pd5nKS8r9NGRuKwVTFY7ZGU/Hphoo0pM30P++VeBLvgNFELDr8QUyJUUxeTcthFk
fZZ2ydsTu+7E+oXf+52alz0n6JkAtf4p3JyR1AfoOtfhLiRYAe/ilF2LYlAOB1Cr
ae6JTQo5uyHa2tb+vAt+m4Jo6B2hxIAg2mi4mpt+Jdlu9nQH+YRjc0tikxRRRK+T
VqfrT30Lydmx6WO74hCtQoNDa/8xcDlJ1ouUVrVQaoWEfPf7ccM8cp50i3b7bV9/
VQp7Fh0kGxeqU7JNwnXOsVv7vlvnBCbTXsIOyVy/nTrilT37ZUkhs5UgLGupi9pW
R+Pr9Pzo2pAIflO9CMrjNyn+jqNNgtu1dG0002dH4++ie9fhzDsM5pshKtODO1O/
78R1g/ACujixRi60ccVhJqgHUXF+9+ZHV3GaNCedey2SfqOhqdSnWSnywZTbh8V7
P+bWNblKLVLHjLSPm6HueSfETFU3nZmTH0Ah4XJ9L0+t+62hY9FOfV9juqfA392i
4+cmlwce8qUorCkREPmFroTjW81rBvST+GC7I1eE1ivneO/FuRng6h1kX9054nCf
Fj7YPsYA57pLpOgZGA0QO4Dmz0kade4MrUa7WDcfnVFgGx20vwoxWfUedtE5bjmE
2g7Ka//vUPPueGNFafNddrOME6tti9fJNjqBXB9vNlqy9khwTgoB+Yu8/XOp4WQI
`protect END_PROTECTED
