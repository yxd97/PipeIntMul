`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
530ixW4mkJUUUYQQQQ+OGD60yVeAlK39zuu/b1s7r15cACZ115WDZjl4LayKsliq
7nf8/uVSA8cwSxsmZaZmR1Wn50Ar8Nn4fLd7ppi21iXZ8ghKPthYc/GkjYUbmL5D
8Rj27ekXAyOCpMnVIDWJdEAzfjtXTHYTdwvvKd9A46OvavVRaKm3D8XF4yvyw5ul
uc0TkkepL8zfW5MaQ3HRZafulUBpp23M//B4fB3SpX2ZEaRpM8As2pp9JJ3lXQkj
u7Bu4OCjhKb6JDw/PA1QdOFWn2LnPfSd6rlzKzti7l4XHRExbuXVRY+/FYjvAqPP
W5I7D7X8oJL0GO/w+2+1rLKXPr596lhp0FQJ0p4JMtwzuMr6l+/mtKzf+XcSEZAb
sHJox7wXAuD6Sz5LBdoQEia20GNpAc77nRAwpE8KOEwlSJ2dbpxibaajeTPCwryU
dKE1yn50XwVOIj2UWKV1DBO8RUZabcFsHc2j3djF0PpYo9k/ORhapMG19RTGL0R2
mYMD7bY1ruzZOXVQyjVlK90vUmhRQwVCFp/FDlpyHywspFzA15UwSw0q9tEA/jzB
UttpTX5ezhiV1U19Wn97+tImCqlU9Of/7bc0wZajj4kTeKoZ+Oa/7Rv1wPdyJ8ZF
BOvd7BD63bdaRt2J6ZbE/eqgUZSe4n2A/iSDH+79u6F1J0DfQJB4hdAP5kjxg9jR
HF5rOeLQ32OXSF++Y+XGuJNuyR015EzKGeDzEUKMTP16jCueEdvqWQ0qLaER8yuz
ZCKzeGYEIFk/qI0lZHrsxRpVgpUvjIHiGcBcDJsoTJd8CDVgS9Nrr0+tIVtBaG+z
xH3txDDYCjQ7e0jV4Q+XAUqqi+O3yBihsmoT17Bw3QFeHcwoFiIR/s/NbQisiigz
qkIttnRbnyUdbmG6z0ySDL70nz2YDyp8DZVxVNKDQkHChB+NduxkOIZK6Y6rvs7p
MQLJhpOij7Rx729BOY6ez3KRHnt5cK3so+GgJuxSD8YVuJdvEkTyrDc7EJxIt+x5
4JBK5GQzpEgg0IA2pVVT+Dm4VD7qa6alXqhauUBN5pW6Hz+rZ7gSMFD3ZrNfQfHT
gBi27pmptKIrXFntgBNFmHDAqhSTIAXo6WHdW/oGrhdrJEDDP7M5lnTWSdJW/0wi
fbkOZswmaIbh0zGOhFsWTRYHumNDfo1277EKIWZpv5HUPSy8lpweljya3f0Fyg7V
boayfg148gV/uY9bODUYxcz98+KWWzJQa9w+I+aOYdfvAYiQfK350MPLw4+G0zvm
oiDTDwOEPmqQ3QDgy+05ze7jXrDtEolEigXD7n15qZQ1Rz650mficJPelm48/FbB
PT/pg+qfTuGoCkzkXKPlm4DT7WyF5YvqCR4Go23LrbqhxjYbm8r1fk/EQZgZSzqx
1gfYlBYqcNswbdOIGVFvOgWErdKGqk6BmLxuFihVugSpQ94JNqUxLLPvdJEhuiyQ
aLOsVKoSICUxCplJVwTSsoXWCaFcuZuRU1vQug12dRZEaIFog6HrDbGk7Y00O80+
q65A+tUV3Ud8qY7GQrT2tPIOPdUtInaf1lFlopk13zpG4ss2N+/W2w1kuXv7fIxp
XWL5fMIH4PQMFjOXx26iLffEvjdaZxK2VYxW0C1YH4X9Efgl8BOBNd82EZ0GHvP4
JFzGwJswcuwZcWIh0viQuS0VfU9Yxsn+aMtydk5b8cI0dI328ae/qsl3KrmlUynO
i7i65QeHr4bTz0Vb2Nsygx/gw5nVrNuzdm2JJJFOei68cG/l17XEewmuvOFXc0ty
IuCZBfDa2jPrLYi7LlAEDE2HkIYB2kYoMVwbNxgXjgdV5+l3blZhRFwMnIwtcSt8
9KfdV/e1ZjBC4Isf1YiROL3zEFY/OCGVZ2vjFm1UKuiWo7hT6Lo21gf8C5ElqO4p
0E7pCvFbYDU5EaLNMtpXnPN71Ha8nXqrUEEmmqtCsY7cbkYSRxvakC6AXLLkANz+
0qSo5DSkOnDx8ipllv8P2wrMaNRZOKb5+uwlG6T2GYKaM5jlms015CksKmDPSYWp
ycWwcYgTo2Bh4iAt6l6IX2V74sHIaMa5q9ZrkJvxxmePpWpeURqSQIdEOA4e25vg
PRb9mYVhBTMsHaO0k9mzNW1DjMWw5UTD2f0KleuWSmMquFp6HDJhgCIjOFHGzv7A
e3EwCRvLB2469XK1XxRtwVhAVkC7CWIBoPcuHJw31iDaz5WW+knYx79T7Lorrlkv
4pj/1gE97eCXuuPmRNRXr65tmjna1SEiprvpGyH7ZVyXhOoFY1RljvzhMU6d8SZQ
g0cYBc83LNZdTPVRGlg1tXTJJZXRbE7IT72YAfDRAyV8d+kSvvUwIIy/k6KxIrp7
W92oyjgroD+Ynf94qucSTYV2chhnE74TheDpt6cDWLEjAnZTDtK7erVAujNxcSj7
UlPfjWWI8q+M/udF5K8aSbMoDynK7XM6YftVjgw9rYFh79r5OQ2czWy1XNVjJ/lV
7/IWfC2Yn2+8xSKOIAQKw9OOPToRdKgi4/VFV8+DvpQbtspbEHFH7qQhSPRjCDgT
TLm/ZrSo6uGb3SXOi4f/zK3VYVjau0KMh/4hmGhXH+1poeeqNOBTjI6l3mr6erV9
H7w95jKNtxiOtiX63hZzAFzISO9H0us/QfJHpJnmc95TSJxVfHf5DEP6/ih/mDIo
VSXUp9fAJwI4PevilaunX1rqrHFshooRWFeArIda8Tm9GvRHma2udPqZVsV7xfLl
1pvxhAAiLRSn1mcdgJQk6wxzj2f0eVuLYcQYXjvS6I3AQMnvu5DbMw9Xhk4aLp1T
9eh5MvBWbYGo8JTPanvjeBU0pJ0NtdUXE351zzCuMRUhSVQvojpIV8HXwOFh+1jO
Khi6QfaTpnwpiLLX9ETG9rlGWWiUbBFiGa+i/QrvsIk6pHlLEPCZ6NU/N0aljWb+
yTplfdq5iGEsVdneLPxMqs/u5+Kbopyka1g5BJA9K33qTyJ02A/MA3yXQQEo44pK
RncP4pX4waK/3JfKeQ4mbMACzzUmvrBNBEq1QLOl8NW5SyKnQ+UOt06hfQzD5aOk
BOzYpK082f+kyuhBYTieHRXwFJUfUUgkivGJG1qpsrJTrP9XyfhDA9mQQEN8Bu12
iPhZHpOQLaiK43RrIviWjWyX7O7UEIsuj2aR1h4sR4uZsEo+Nklb+Y33CswamSp1
kICFiWb5Z4CAeovkPfRjTgj4ugHWhKuysbuoQhYiQchBEYd1aYiZ7d9aWEnuH2KI
bOfQnpVcUCrTKpfejCD7dRz47MiKuGWONqStaXnf2CNgCtGdMCAjPP/AeXFa8hwC
IfMCJBQdLhrLBEIdtGZ4hZ3loIBFWGxIczJGZCbT4dLaIjlxj4tQG/QkkugxFNi7
nuKuMpl+jufpJqU+YxaNEOkbEb8robng1/yk6uzIwmwZr47NwPZFB9Wtbc7f0QKp
ftm96Z1fuxhfgd7zGGTrRnm1xwLG2nEgeA0L4LlTPdEe8eFKNQIiIeJuPdBrIT0W
HGquEHCm/6ji+aS/LZ4dAqRfkWJj+bAKz+3F5OdyxdHWnXkzB/EsAzqh6FCOdA3M
xYI95ov5pi0KCzhnz5fR07te0qa+bUDFaeeKNcIHJCXUC7+I7OpAEoIT/HN8JY+u
vSO6F2Pk7MzOYp4WbsgeUavE2eT3WRZiZh9sBbh+HonhGM+nsT6cqVBM8w152IR1
OrlSwSUolaukLaXRGauf+x3H/yMWiT6flRqTfTeN74le3JsjVIo3y465zCCsIYnE
/xpeQMErKh2aZkeHB9D7rKKMytJXDIQ5feJPLLEHGNvJLLJ4zhHZQqzeQu9UkGIB
HYJBhYdmvW/fL/BeN2Vd9oBjDbl/9OBPssFXtPL5hxQ4999c9dXYWfkPAHD1GD5N
ycpaOG8YmWaXEvpZklCIAuos3wDtx80qlrv0WVnNqcCKVtWt6luBueC0ilKtSQzu
HsmuVXrxvFdhdUEz1mQAIPxPNFBtiDN4YoSzC46SRuWyrlduLBkA5XPzibd6l/1U
w6FiRuxITJA924lfKTaILhi5GbPjwipBP7a83/mXAs8ZJuXFBc31tqDbPWxjEXyv
wtkPXuyTOshFf5FKayQta2OjgLdpXrRCy5OjBWYgOR3RAGO6Bz+itWDuwdZXNLw6
V4m4yTZDpi3vVS+xtISQzlVTCVMdtA4SqjGb1j0qLlviLegGz1h7Mv0YaJ5Siwb+
4lvygREg79Gyhh2rvdmHXP4wdWmRCZE5+RbpQ00Iq1EzUDTVKh/HFwMqV4OsIizM
AXqofNuUeht9kNTSxAS6ywcJ4io8yZd6zWyqBx7NBjxOj8rkFr79gUZkZBmQLsPM
QH5Fm7C9reiiKWAQClg3QXkoJr+2xsP843OTSGTv7/M2b8gI5mIxg/C7mwTBKega
uI4mgCRKutGU1QDSP2Mxnkdu9Vk2Ael0djht3H+51wVp6NmNC/BQI5WGA3SZkeMt
3GZKOC9ux/y+ftGp4HGbDdaOhEo71vJJqbEEvryef3T42M4vXs/L382o7jgo1hcw
A74ffdZ3eBYRrkTLn+zooVE5nk6crUcNukHNGWYL/xlc2HOMt9KI+eLJA+Ce0ocy
Ez8CICwJJNMeUe13fj5BLaCjp+QqTvaPZkDEHYIrhj76lTypeavjfdmjIBienaxs
EbrBQyZVodLY61O4FaPFMwMDuj8gQPPE+BqGxPr0q8r1nGwLpdmb7ugBS3V+jEho
p+vtzcL5ptsnmOnBSiV+9m3j2B6kRSAm3yW11g+GO/CphKzNy1imB7VNBqpeYX78
QTdeegPNnsDqXVThXZCEMd7fWyuipnNIi8FA42VcXCjj6h+eryRjUCoro1UptaaG
sc+wXAjVZmi6HeUgeAjw8axpoVvmM00SXKabeGwgNiSBBC/eiltIfD7erUZptUnl
e+T8ASAvuxQgKERqXa4Wl9ZUVo8IMVeNJF1JnQbMYDiCf8eE4bb+vrn72HviwGb/
l2jpNxXE7FnzV2l0GabTpQMsg0V2yBf2INnS3E0idgv2lBzatrmYreKXVcexdyzD
aKb0WjNKfs8gWvqPjCeSo2D/DtdG7jNo7osGaDvlSynNI644p636m2BGsMFPrKWV
iMgW5IfBQZmbo3SWETC//LKTAdVOcBcttf2JaHw1bWDCNdO9dNuF9/5wgMj4K+HG
2/NMprbUPQnm8sJGGThDPMCFjfH13M7Rr1g63uTVB6y1J0t2F7JJqNsghvbcLgt5
/rOHRN0Zl2HY/va5+J3CTJlgeX1BZPycJoo7P3qZlYuT7QUbPaNbrhIyJ0WFffBI
FzxVHe4fpunEZPCJQU7Cq7DjQwbXKAdyo3juKaJxQ41bqcgBisrv82DpEbS0svmD
AXzPAg9gSfSfQZVbhouc/d1SmS2VB0H+htsaxyQxngwzZUuNwNGrddmgAXgKtKAv
0SVv6/IZXZf5rnJna8grZITq4rU0pSuhevyW8+VvfFKkJCNCXj2Ld0xPDvpXfeo/
IlJwbMErLMp7Ic7RPgfasS+hXp+LGNoaYYo9A6TtTxzATc4nqmwBZewTcBH21WpI
m3shEwroNcplwmoQYIDvEojsmy0mEqUEZCkBxo+ACoPLXpkbvxWenMocDkS4vKjk
ozhBdbAXiD+PSJehBcxKAttpA16nZGSJq5ZPB+ud3L4TCbG9llQq4/8qpnvXxTs/
cfKXYUiLctv3MK+4IHNanwdZBsNqzt76gKAAF3rDTEWqnDM+B0YQCw5VCmbAy5VW
5IhZdRSNMGr+37OnvDdltvKRzTGkTS9VMy9fInA5nwE4tVI4X+9b4nGpaqF9NsBW
S6pto8V4XkpcG7Pp6yvcfsEONM3ZcUOhMYpSHlbBMIoTCx71+xsdeJtPfJTxmCBD
auncnDcYnvznlalXoKPDXRGQmyYZ6KqQzkaHMtgUYyufuFC0+r0o6YYwkQS1llqx
iFcUNzZbkER1epZORrl6tJqqQCG2J/GQvZYqkqKPpyQU1W6pN6hQGd/8s59tXPHE
1Ni9wtiLfym1errkdma5xKewx0UNyimJ0vdPdn3PmlxETj749mmhGEhipCevfIzN
j+pirtxr680bm5UQEDMQ0WlQM6HDguugLmlsO6rvKU+w61ZEk7KcbRnP6LXF9obs
15/6JO3JBIb++i+l8hDWA8quRSaqDxm/26ft0tNyd4CJ3I115GZEP5d1khnCMEhy
Z9yzsgbstoEQeB8oM8OtOn8cWAnd7CdT25L8Te00yr3+KHK8qSJHFh0+yBMUDwCJ
uhD5wAUPXotoYlNMBKcUP8HcCqBpm91hQnid9EilNfgS7fSaUbHkSW3/Lsv/gG19
5UyZrdDTVCulO6CGIyN8beywccB8p8U6n7GADWbebWP6Zj5HbKxahXIhIDcTja/Q
SEFF0Rmfc0p/XKDIrLFUoxfbjx8DXV/LfQI7gTA5XtAr+lG+vQN42V/PgaYfQElX
AA3vv0zZsvEcZOzAgvhgtMYx9YxHT4R2ZOrrq9p/t0vmDbMnO3/KHZEQrm3Tovjm
q2uhbqW2xptZVI69aVC0uvWES2wZNc+5R0toVAaYXwjt7r9RlQsUuLTvVeI1T0qg
MHWqMWs/2lROxFH5X1FMOkIEYoe+DX6w6kliXoGlj8dDYTN1dflswRigJxCLudSJ
8IrH4lZXD/KHmIxTSZ8CU97ddCnr8t4TZRyfW9ae4g1PMlwvCVP441FvFjXAeDB5
EPgsPtcTPLK1xwMzGSMP3GuoI3jiPxuwkv6Pm1nuths0s5VlDPRlRB+OaRghruTj
YcX3EZd5V+9Fm4YxUnbVrn0Bry2/6ZqzGr8Qlj80gcLolrbz8NdQ7LDXaLOX0doW
XNWX3CUPQg8sPzJTlFkw3KMPuh6z5X49ckIhMB0l9tcvC8QqRfYFOb4KuLKM03R/
HSBvahBUhBgplaLRJtaodhOO9p8AATyuKijWOiEz5IFfR9zBW1+wW+ePmyl6bLzP
lNqBcez/PNk8SUgNzSqHNch3QniR6UpAYsPnWckkWbrLnGHR1mVcEUlQxqiCxBjT
3NzPB9aU6kemdCq4xhHXRMi9chnxO0wEOelCAhAvIw5ubcEmX93DunAcp6MvFAwY
CUXD9yeIEsESICCx5N8KogBA4CFH04wkzdc0/029ofyy8dGiVDi0ys2rObKhaHoJ
Yxv24C9fKqBXrQBdE/MYz9fKFsf4rJJtwlwa8xhcj32tA+noA12zsjHRG92Qp01Y
6rjlTjSeIWL2MGQA3F+Dy7kJoEU6ID7ofJOvt8cuJNV5EHReq5WoL72Sejum29+V
ehNgPkWbk7h4CkjW76FEw9llXj7ToyiknGbI1zmGX9vfLwhPmZ3SO8y67LmAHftT
qQgF/N2vhixVrCpa+CaI8VCOVbUtbqoZCyCpb/70+mdHJKmH3aLw8/FaBdtyLS9q
aDf/+RZ6Nq+8B6mQI4AnmvjKqzoMNzA0SdaP+5LQAfmFO4QTAp8nw/95LScYeoXi
kRr8UQY+XQOwsV+2SzUEO3guHTg+IHaTXPadbfz/0wAIArVw5vPkt1V12U8L/W9t
SnJe2Yu0gdy3gQdi8dsDmG2xoVlycFwt2uU6l+NsUd8mW3TItX71tgwmCAKqLWy5
RXkAAAOhOju1Hoa9Sy/1G6VaEza/QzKZMx/MvBC5E+rxB2lMuxXwVBZgaj8eG+dY
qqKHMeFPlD6W6ZoW84wM/JTgPrpSOPgzuj/FVp2KeK5XtbJQuVT88mwPu45Ausf+
wW5shrTZIy3vrBFOte0WX6g38k/lbO91I6GxeQr5OuggPCi/Tu3bfIaUa/xKWbjb
1HxccpHxYCeOG60rfsStrpOLYZz4uOz0UwwcJIP1eNqThCb6LZf9SGby4569/ogS
VLtwYNIhL4HPqIIVmPZmIQD8EIOIiTh13g79sdtq3l+qxp5Dgbv4Oq40OCnMdEMo
lQ7IpWGQ/zb/GW9ifFZfE6B/JhYbJa4027K6/RZK2UQwm4m4hNtK3ufUfYh52tzl
wV2wnJfq/xCB4r9k/kh2T/QGiL4wxgyeg1Zda0vv6SIco+wMn1a7aW7+TFFfd4Nq
Yy5+aYKXzFJy7vx0UQgrszdUfVe6kvyULblUU31AoByz8srDV/KcDZEaEZp5TaYj
PhJHJIF06k38+WzOfdPMwXpkWTL2eFrl9e0c6VgCW6+qf+oAJ7xrsZI23SRBbWdO
RAwI9uL9URIwA5c5RN4ILECWFEH8/OF3AVe2CqmIL6HLJ7bF1uaKaQiqzt2tpMTL
Xl6I5uvaGvZxjo7Ais6iINwkysjl52n0e0AD6m0qKOM544Zldqudf0JNNXoX1SDO
IAmo6Mx3Zn/axiZ0SdTLWeLAAoxBoBQdG58OwXn8x314Wbxw20DuKB8A9C8Ar3oX
UEBv74YzYIBLQF5/zin75dEaDR5dkVG2lIoq0LX8X46a+mLeSk6BbWDkPVArje/T
ihzsxz7AXGXxabhbco2Abm5iB1CebUEFvMUdeMFkbM7Cp3/Ri5z8fBxPUk/J4DvC
I6tFvoea/UPtOU7lsPS2fKzD+iUjY4n2pQ78/0YK08gTAr11j3eh4l0kTAjAEH5U
/VYyqN5qOzIEE9TC5iOsMxHfh2qRN6+bbfk7wrDg07xZ86J2v7rB7b5nV0izkB/e
5qqNpEOnwsA6pTDm2LZJXhBrKj6+QnZbtEuEKZ2WyhCa7EbfS1Y/HcURbw2FoTHY
s6TUbGgzKy+qz+y+yaiUxG2zQqJCCxififFK1aK7+vhpi14k9xkaxn9Q7mFmSdtu
q347wMlcC1jPYB2M+OLKWUItucHn+z4DuZFIk+o8sEEw04BdukBkRCR2N/g2LvdQ
HggBJUUV5BM3fMe/tUGvk7SUMWFtM/eQV2+UVCERRMeYRQZOEy3LCvv++/OKOL2I
b/84nCYJyl74bPxGkLW6ew+0adsu9b9K8/hf65lGv07UCp6vFNlpu9hGQHV7xPra
w06oWKNf5wjRnIwKMjhAR2168m/UixluZRdoBFQK/RHkMvBWshdob2KlY9rexhRi
ngyFv0A6oDcQQT8CQxdQOjonYhEsf7D7Bjc4kbFOve+nsgZcLaiUCXEvCWpoRsYl
ghM8S9oj0F/NBXNHFcfdnxGEfI9lp/nPFuCEsdHGjefnxRVRmX04pYj7yVL4cCvM
SNlwz8+ln8+pg4kqLk0URfu+om8QwVZ/NV+rV9XY0RLFAB53MNqaKVO0LUGA5yfI
TGbnfbb0lVzLXoiRPemW3lOgXK3z0z12GdqhHZgGu85vqugLAhX0oNxH7HwKbCAD
6LlP6YDHYDGUS5eLw/QnzA9Xc6PExZBAcaPNGsGvflhccCnVzuuRVkOYyuiJOR14
fuTzabVZT/ryEaq3Hgn7xXf7X/SXJ+NsUbEQpG/bwzeHWxxGF94sPqdJttYMHFAY
BGZAWQ4xnKCV1hvPFe53E6gA0L76k6G4i+ZifIJBT7Jrdliywqv1umeo381ifm5W
xFcjJzQPjXDSFHDkbNeljjogJfQj7j1JD8GzWvARRI38x2YzRBCSfpVKdUhpISNe
RlR0M7v8pPqKWGfusNZYo9JRJjluaIJ7TkyDnVogZGYmVoMj59RSoCGmBD5dlrkz
pRQsQsg11D7MYf0lb+bcKWs/Cus/Zg5Dn4Ay0gijOFgrYOVyjD4eClNPUf37R5hh
0Qh5CY/txd8L3BNMQtWaVh8GJhA87mlqTpEoJ5qgYxpOBZNvzW98MqrvbYdBs4N6
0Iv7remTw4EOaPsE76hgagNz399JGuwY/BqMxr0ywjbZoKTVQJQkNt0TOry1O0UU
/bdsQe1G4GUw4bvhlPOF5vizIvWiYXKAjO24c6CVqymV/cXLWANJuLHlLdth7e5r
6MSUfmv+T8qb7U4dFrfxAGn2TmN5gDlveQ7YIrgx8TFW29eurMPhrz6NJzLz1/2q
yyp0AIrtmCUKBpwxU/eA2iwIKSQoEb2znCrlDX4W62ahrWg6K/sMo3E2Bizj/CFX
nIMilDU+hTCgKUg+cK9agXZhZ1An6k+pYNFy7O7I5USZCoNJhAEgAvzbmreo3Y/z
+srtKKvM5NgtsiWX4X2JzhUfktF7U6ndQkNc9RHh2tZmLWvuRIG/Vp5EJfe/e+E4
3kvPI4Y41HTNrsMQ23kcTnJr836wf1A7wgs1gWo0CepgYMIl41aoEJ99yaenej8+
OvO+3D1s0Rxl+QIVWvpyMd+J2tUuDHtGFdiNjK7aohEu2tGI+48rccAvNSF/jzjP
iR3s5iOvCJJCBIJ5ASz5fyw8Kjoh0o/tnhJNzWJvuqQpFuKRAhzoCta0+uzUUGgw
VwcqZuRnJJYBvql5+O7LgkhL7sM46ZCCRyqO8zAprNkAWiKSALTg5p0DsCgsLexb
HB4nUkEWGU+46q6A7k8fSKT0mMxGwpNWIhDoJQhQ7L0IAsF/5GZKO2QlF8DU4R4+
XTpO3yLqGJXRVvNCTyWaGfqYXw8fQSxkhQ5In4MAwMaXlVTpzgAiO7nEzBLQ1YhG
8o0EXQfFMVsoHuoLjsCwelMyi0keRthJ/9N2FboO0+x+pCxjUaKZDSh0ARVSqkna
r0zormnTRmBrdMaYbuYibO1hF2ln/XpcPmwUQqLcrn5ye1XkfFywQqA5hyRPqBGj
5WzpyIyxWv+Xooa2RuUtPOYgSbok1Q3AvuZE3rgqJkVCIJfBN0BQ8l8rCLozj6js
Lf0xi6M7WjFz+exItrlrJsWENCFvGw8H6EMqcikUsbsKv190PPKsihpElw5mHJDp
obs2yLaPEzOG6/Cvb9DhAWuVSjO+/TlUeDp7HbS+cYT9hOT+9UjeDKLD3JvT8i+V
qn7j/TarWydz4bZJwZMLtCOFSyJ0cmHESCcmEitAEkqxiOSHzHv7HmR+2baZPRx0
LW+V0ee2e4WeKmLY+pB8svlQnumleISgRkIhU2Y0Q4KQXLRM56T8Idxocf5M4UhI
5YQi43DyBpG/NAdgxaBU1Ca1WQp21nN2J/q+Rzw9ZH3wKiQEE+GeSp5WhML2MVQ7
dKMG2lqWAvcxzztuJqlq8cEI5USRAEEDY99Xr/ve17jsTZOlPeFTFLQlqosXAtzQ
nHDb/cqfNmbhfp5SFJ3Q7Q9EacPrX3ZYtiprzW1u9TnpL5cPgPWT1Vnch58ZJfHj
xt8VL6gWKcwboqwr4uIKQadhacc+ejugIzDiNoygy7Xv3sY0fzT1L8TTjjNy6FE8
7k3ddGhvzw0v0YVkm08v4xU5NLca4AUmivgCOBYDDSIg1TPfMUW4GSgG5bgnqIeK
Sjm2syqSiwTJFmKvBdDnyJPjKaTczDgHWZ56KUR0wAbz3w0phxB9uECN5tVHWj6O
HY5+2ahE/oV7LMosZve2zWg8qEw7DpUlx2nTppqkyHzfp5IDDqH3u+sEJs+OhsYp
xmwKLXffUeJAeKlHQH6ZuzLc/ONdRYhl1D0omLRhILeCONONzJx7y36wDVHnRvZB
F+dmJC9HjohOmj5GwnxJ1+eCZq7prpRJJKmhFSU7/4YqNDTdTg/egh/zTsrwaWQf
+NUkzCqxXv7cWBa3fhvw5Y+xyLuNGLPfMc6EQwPOPwh3p6AMTNOCv0xyoxo0Rd1Y
PIecC+wUQqteG9q4mcov4xqkaep+Jpup7bV6AalaU1s7Xw6b2NxCXQnv1gOgkN3k
a+eOwEwOmtUykTqqZawtwuAluvxD7celPOvQe9qj/WeeluVBCeumMajXB90BzPN3
hZaGplHtXIHjDk5fUPXCuXUTvmlBP7Au+8+/SjV2E+2xVzGpppM+QAWH1U0YXrfw
Oc8FlOQcWdvExIat9SnHoyDOa3nuljGSxkkcRQMjTAS5PDMium4YgY8C9p8POaTN
1ge33pNYTLawBGAJyUQAs1u4l60a9n9Hoi3D216lkQOjc7nT1IbEs5KrR4Lt9r4C
ZowmdXy5QLdjkrKwKiwbRqOY3qlhCPv0aggEF39WP6uo1RvEnACTIYXrKt1xg8GU
duE2vq4JS9FqsYYYLnYxE/S1HjYZ9d8t6MJOvQ2TimqUxRMl1a0wjEP0NXYdV/dZ
UQGFlltgsYuifVRJoVTJUDDahRIUjhLhWFqjgiQ7Xr3o5RRFF+IQ3zQO9x/Sqv+X
y87NEdO9ulD+QAkE1TWkqOSEHBfbSsXWxYNbp3dyg4TGusQqTX/yUz9uNfGWgFVg
ga8NjBaQ2YKHacFV9OS0dsQSul6+6ARs428CYrxTPQXVQt+W12g5GP27hjYQ8PUA
EkQaG7oaJdwqz3gU2pfF1ZprTRllmKRKOH0quxzR7PPndwXbSEZJ60H+6rXS47KR
J525Tnah39ZfQ8WtdEIPBQHsilugkCrAPRCRZ3eyZRiKoY7kEifbGTZ2wULg/Agw
kiwieVeMW9YH83j58lDkCgDznry9A9sszNv21fRlPiNx0t2yYuOZk09zSHSQ9M2r
ZDc7n/ZTUVy7J2FOA4ncHjHNZe75Ymdf/HuuHamuPQaE/T5oLZLWJ09ThAmSuoNM
kSPxu8i2DvEb2QVPWj93ug4JjPVqTtJPEplFk4CJx8eAmhOBZira6fcLK9xEK6YC
YPWiGMMsR2zxma7q79gCYWuz1senMH+ya2rWc60lcCcHwiUMRT2sSkYOJVfLrBVH
pq+hGa0QrKaEyQKIt3SRTvbKXywu01Ke/X/rk0IuocTCYTa+mTDuSbpXJ5N6075j
cp/oLc3xdJSLg42FoJgdRKjdNVRBIwuV5CcYVsgL01b/uvRAU/K3GE4jzsaEweFE
z+CAZOvRUTrkPaANIru81Ci9I21S4VfORw3C9xiNoHqqQabHdjNVF9LILZBeNL7a
pbBACh6EgRwRk9PUNkDQdTnuGcnjpBNDR+RTuuuzSnJT55YT5MMgtiVgR5aw2kL+
oLwImulcAK0e/KqN+D3pZlb0lBvaHxPMB9Ku1wUCE58KYbD2vrbbXq56v4qsu3Gb
UNmsKiN36eaKM7aOswIKXaB0OHj0AUdByHNiDokgp20oyiu1h5Q8nEvno5iZqHa9
m0hEosANPLgRdNYq0zhxIpSAADQpqYTFHeqTiMxxR4iFiHDepcTNn7zWB1fuUZuV
HzXqnztBHm+0W0IsOt0wijOlvFUMBLP7SoaobXd4UnrGZEodJDef2/plLgsGwdYH
T1qlSru2ybgOV7HNnnTbPzzrKSSoacV+ZJluGKsiNRXsp3+nsFF6vkse8vQawzys
Fejiz4AiTAJH6q+/LoiXOA3ps3w/8XpeUIG2mgkjFX8W1HbdGLdnmFfQDO7uohgo
5msO4IioXGDJFCLIsxaDzuZYk7XHYXk5PYhTluHKdrWEX9G7RnTB9tgJweUpL32J
hQHsIwTLPeBh6imWskO/Z50TfEyB+Q+bmgVhfvwoWIvKn2idW4bzcHL9XcBQHXkS
C6XqPiaSMn+GkgEQep5K0b0FLtVwyhW+ok6yvuH1br22S5JDRCDKbloUsaQL2fxO
uOuWFnrWhrECWKIaXTvHzsjXtvoNmDjoEDSEoFH+0qctPVXYv4mJPnciRi9Rx2ei
H/QlYfnOpk431Drc9nlMMhiGltSUuvCsbYwE+8anrVO+BGGWHLixClfK7Ghtfoxc
tJD0TsL/QtsZp85L3c07m1eHr+1uo31oY62Hn/cACpe6L4b1msIxs5Lk7kSZciCx
cmkL+BboYLsFxt7A/2xzgm4JWDG8rBLFRL9GkrK4aRRzmw0NOhyOEAp0IsTq5w7b
harhlRKzrOUSQ2k7ucCZ44Rbd4TlJlZoDvMjStvM5w9sNggftFZreGQXD331gPtL
LcPN+5+d8Tcb95uyWcD5KkHMFKetHk9g9Mg3BryDFiJx77/B1zdT8O3F+lTUULsm
TBXDkXLqLr19+RQ0r3Ze27NTwyLFoJ3H7lFImHvX3wg8MAudZV/ADtx0vmTGb1+A
IpMU5JEZEheZSIRA9+T16uoQpOk/REvOXflJakubEEml17NL/5cmeAuMUGTxiUi1
CwmlCNVE6cI2GpusQ7ZSBqsBnI8tYJuO7Z+ZQ0uixlTxNT584dpcZ4jlZ6oRsuke
402PL4ww+UPCoDhB5CoiDZF6HKsft1N7HeSg4TpAEpzeHd/NixsmHd8YfJ3pnvfY
gwnWd+TenDVlyoTX3399zPXWCdxHbx9EcWBeCW+NOWALu7Qd0QYk7I1OHAI3g+X3
R9iQJ49qY2xvMNsfe98lTPKFSbbh/bRRPqfEXf3A6rOw62hhOkV49nUKAUF9iktU
olawv4F2cqkofjklFG/bk64AZu4eMOM7Yz/UlY/ipOwd1AB831khSFAb994DmVMa
rB/YIQ8AOchgsNxUdhtOeityN1VgxCb1C3AwWuREuTlLCpBM3Jh7MDkK0/RjQydJ
6eocFtor8hHf4vxtYAyBTEhKH0DclMP3DUey7CeiZBRIj+xwY+0ndHm0q38Yj8NP
5dqpODrL0m1plPSm5w7PJMpJCFLNXjLdwIPyqGwOJghCBXlxR1PMyi443+QF+SrR
agOih3Yd8Si5lXc9KFvE3qQQ8N4Otz8my0dDBu6p8Jg9SvyFPs0+No8j5tRFplDi
0c5ZGAmGu5JSr0rksUTs/6LPazfx9iFZcY95WI/4H39vf8EvB1pqRD5QYEtdhHph
MWIqL7dWIe8NWbPUVhtdxy8hb6MvfYDX4p4ctJOQU0NYGgEzdr+DgFjCvyb+HrQP
2XVieLc1YvM7UaM09AKvkXZ9vuzdcZSnOOzeDVXbowdfXgrBu+nxXn0/6NI6GxDM
v8JyOwv0JEIx4083nNDBqltvGfsMkA491QRVfD2Pf7iRWbKtKH16cYcsVOd9Bn1Z
sADLpcCsTEaCuYZMs0CvNoJS/9nWLdoo5zcK6MqASA/6NgPEBwId5wCNVzmucyn8
FWglzwp9RuEuB2MoUofsSkS9urT2mtBs9x5S0if8uDsqJTtHdkvKzXPM0VgjwaCq
9ofxXXrDWDO5y3SioNHp+YLWMWt1iugLpVBiUbWTytAnpJqk+Tq1srxscGp5pFou
Owl0JJVzYYFWQfAib+nlMANbYKN5n1/wxQbGKLsWRcfbiePCf15IvF9Gtpqo3KgK
zBYfRg5HleLpr5iu2zLEtlFctEmjidGurbkfBaJbYBj2FaKSS0UWgoH3w+6Qf3/I
IYgBacJW/6llUvNLENSEdVPlmlCWQ7vWY/g3Yh2HRjFku1lorL25B8z/LBJbcKaW
GZ1cQGJIyR3IeEvBKapyFsoLFdbrmnp80q+Qj0Ov+xaeiHVSaOEow6kkn4V7Ol3r
F+NSI74a0qjn0Z6BAo1CW2lnU+CK8FMTJKqFG3hJLMk8EkdYv474JrRw+XFGXHZL
HN28mf1TBFGI5n4IKqCLkw9E5WDeiQn8G233hlCg5oQ2/wh8/kRWAjz8VY+Pn7O+
3+LLHUOLZ4lOOA6M7bXCS7sZy2b95XYP8CSWOQtTM0mAmOu4jWxOscQJCuOjdPNb
dLn9lzE0oXzNJOfx4yGYrpDKzMyagUseX11cpC/QHjysvs3hKKagZFSV6W68XS/G
z7l8MAGSycZhVDSPts6pbppYSeaOaf15mJftX6NGuBzV3HCK4ZtK8cxIPMUDo4kp
ObJzlGwaxXG1/SCl1IXh3hECWKhWvVHyHBF+LhzffkYPMhcuPS/MTL3nVQwPtTh+
7f8W0fPexW2M7nnDZ9HUyQ9w5iRuKSsB+mTR+ad5jeoNYxOB/dKihSixBk13JqJL
Oy0I8TzBmPb4tDIBYZE0NeSCU5HcM5ueMKq4D/Mnz4A2r4upmaJcHqa2sfoiNLrA
Ln/sOIIaSLIfTD5ezgKplQgURqSCRfAOqZYzUrg0/Pnr3vXwQd4oVIW+rjOH+U+a
RcIZzBkdWftJSlZc6jKXhcLCwZZVWvSvtJwiwSOSsNR+gxmfAUSkHyNvrj3rSHNr
wOeHRIKdL0EHno5PTlv8DBj/TsPKlcMX+m53VAg1+wGrLvooJ4PMJfDckcdPbBjm
US1rQ8gO3MYX70xG7K4xMCHJl6w0yrSb5VpqpAheFSzvtThg9KyQqTfSCLXfvQ2b
PJju/pwzMQapmhLinlqj9xGjGJK55dAFnxadK+bp3KKtsY9lacW39aL4fFnWb89S
qRN7RB3RyBLy2ZoNl5OnFuO1Rm9tE/m+3yMxbb58AZoXohHEC8jvasHHlVUBbqv1
7LtKJiWkW4ZhYg6Jh1EYTmmGVcBV/ZO4wfIeWP0xqrdrES4FwpzLBEU7qXUKGci1
tP/My3avvP5s1LZI4Z00AHVj/p8HJuT2p9Yfj3aSPcGcL+GjThfXzDDHurxb0hfu
vHJeyupH9aOrc8FxLFE4QiWoYzK6xsE6rM+jiAWvb4yA3dRqHRSgY1cn46B7iRtK
URRx2fDNEQIWYVVqcUPea9zrFRZTvFWUnvpl4NpOc4CYBAWCpt/eLfK/HULjwivZ
zAEjP8qbtuT2f7Hr1XHnlTcXbZBe9KVp99PW5vrcAPfYjmNZ37qTFPXXY3vjgquE
JGturJSmARTh0GwRY+tBTzYcRW9mahbRl++OkS3ZRCaI5c/ktA8P10SeAtZoRrE6
TP7GcON9GVJmRUWOdQff9CwDRllD/Mvo8yJHUmoquRb7Au5d35dFQnx7LxtlyoXC
kNQNaLsGAzYvJqaVluXAIuecpywx+Z0Do1LssB9+sQtLh5SmbSh7g6KZ5c4JXHXU
pB9L0c5cLqOLVjh7a3u50u6z1QYPbaE7BESEDRXXMGHvbUuKXUctpm++83gDyZov
QdRvPijxScCA7QNUh6yH0POuq2BqjCoPWLTAGLrij1eYgNepHEqcWVtdetXg2cyN
ylF1q4S/fCyxze7g/hEoi7TyvPR1zWyTvXQNsfMj7ux86eBDkO0yI1fLoDXg50t3
yUFjlXsldCHKyfl3oaY9Us7Jg+Cn69wuN2KNAmcX64KNshVi0FteagLz+vpKgjqr
`protect END_PROTECTED
