`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+th2cQDHMinal8np0n4dzgEZDEbHdCwwBDHZEGDNnLfZOmr7Q/iNfvUq3qewtUVv
zQutwSdoS6VjnYs3ipDhxOzRy8DGn1qbSvmm+JuGyQv6U4cSoxSrjZ2u7twQHhOI
gx4Tnt75LKWwPST+VCK9UJrXiMf1HLb+BKVIeVna2DrHLx3pOO7B7mHIkbzGpCxD
fU1D5JbpecCYJUh/McFzzLNrMpWndsc7HHfGT+4QgtWapYB27jUBrdYgrtzt3nL9
Zyv093Xwsn6DWGbJitOj7mJY2CesbUo2lJsj4qEQIykyblZgecRYQukvJKj8OqYK
KbLDpxZW0HJ+t9nkemz5AMjEVN7qE5GzIk7lHzLaNldmg7244IuDYDE07R7MlthI
2gDy+I25YJMGsyiuVCv3dzLZ88o6C1MAZ2kTyvICwiNPbwf2hNcnNgSebBsIVNFh
gLq1bkj4zx0dJsZK9a1QkZjgQ0ZINSAQoY/e43tdPnWBlP4Usme7hoisDBdkwwlY
EAGEZ0Tbi5FHO36bmHkVxDtoHGqOQQjq8cXhObbNhVx+wj7Pd6VLHLvWwSWc6Cpv
Hq4gL/ePh0G0QMDx62kq12kiQpUM7mvtFJzcKTL3+w1Vel9sQvhVc8fTRq7qtGB3
bbvihGSp8dNw8c/XCYWgLqHD5Tk3P03VE6b6lkujR4O2yWZih5II+HApaTFmai1Q
dwvDQf/MSVFcSqUm3IGxXYaQxOjOF8v2R6q+E4+8OSL67HYF2yGOhQgTy5/GptBO
wUhDFXlMdQy0/rFl/wSD/2RiaIp+HNTk+NFzku6LjUk1FrJz2Tye6VShmIFGiy9f
MwnBT/DpHDGzI7xPzcorjw==
`protect END_PROTECTED
