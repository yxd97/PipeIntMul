`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZFCnt94T5xT6lOLuJV1Ak9oUiBMb+yvoJUi/bPg1wzjorym7MpKXBAPbHn8b1Rfc
ebt41gSnf12RHtgj+l5p78PyFydIaUWdjIO+qKnIGKJHOn5GTsA85nKek404qePk
d2D9A4If6LVeXfu2g9XAtCRDdiGWfQOY81m4gWRElj5I328iHYfHQhojv2Ugf5Yr
IymM93M8kofIbewXcbyheVGiVISd3mCzqT+/2fEm5tgMtlQJyqNviTdsKGuMtX6h
PrUXDYSnCcTRmwu7WcxyOSA2H037s5bY00yutynMCgtrPtuzex7Nfav8vuFX5uxM
qiuFDtB3FbZUnRQfs3IPKhpj1gYqz8nIYcxwDgjDl5IZ9ur8yC92v1k8Q3MzOCWD
vok+v4xKzQwvjI+FCkYrJtq/wJsQ8dJS1e3LPGK8+pFoMgqBabuH8Nmvp04/sVER
RbYbdU4M45LbkTiOGRbqbzA3yqYbVp7ZTb85rQiP/jbRR16S+vCA1ib3xWi6gh78
oEMBW2QEet01vyarH05SkV2gsDJcxaiM5ZF4jogT5cvTauuKt9n5sCDWNLp/NpXQ
kqUx5oULgoiet7LIt82eGrwl4a3iVCbl/MDHfHxvjJM=
`protect END_PROTECTED
