`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sbS4UkICrnhYhyF5Ug1cnxAzOB4F0qiA2VV/Zf65BjuAkSmZkyxgQsCSDLwO560j
G8Dbya52m+8SB+7t3JGLARRFnXydHqAY7efcIvFUn0U1EGBJ0x9e9l8fcJEY90jw
9jBkzFONsbLDYfZK0ZEhcTLzDij6P0dIV7yB/afMlK+IT30tf0Px71uiNlwSsMcD
RHaGo8ovYRsYP+ZHHBBYmXNCQFd/LleIJQ4hpcgpat9mxKf0q5ipcGNySz4Eap8n
VLVOoIH0x3gADiaWpxTaIzfVgcAJvgiq0kXh6QCjUsl9Duo+X4IbdjtrHX4gNURr
3wRMNtOl/yugVg3Vi2VPk3yUWynYqcS3Lh3NQvSaat8=
`protect END_PROTECTED
