`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TO56MFtTXeRdBX8eBiMEU8HYil1Zc6rHfp+keMEOsfK4L70QuTtZkBiFu9jTI+ts
NEqkTELhGG9jsfWN3tkCQMeMATofvb2rDPudp18iSqUQMl/Ff4nJAMwo888TgKtL
41ydSx4W1yx34Bg49EhzOHc+Hc1azCMRgOtvRIUf4wsNuLXHuczDdIx5ir7rfk8j
sMFDt3hAaJXjzBO2cBcnQVa9wgrGwvYBrJEDDzYl1vv6g0HNnZ+WCt6kudCkmQcX
3gla3ADf6xgwLLoBOUFaLG9n73uBfAQ1FVtcZvH3Svrou7k3YB5JCH+mMxcjoAwn
ZwxSyHUEAspx22UPp5z0QaNf60Sqi7PRSW9MLU+ltavnogzMstCSBUCeVUc//dW7
JXvlvmtVGaC7aIJLwDDerPD4ZnUnIlIYslmL0ku5RrDYV//PxHxi0MfCBvYyro8s
`protect END_PROTECTED
