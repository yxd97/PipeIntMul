`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qirXRPTGV1UKEKKOUNvVufaEbgAxaHwAo6OYsr1DN1+RWPPj/fX1OaoFn9CEV0+q
qd34Lvx9q1X0ZOeSyGC9f/Eh33y3+Etml2eqEU2xN1sdKtq+ZH9f1Blt+nVRTIkU
1r8YRucewmXmxaXDGLpD5SwTsW+Vceeyu9mx+7FiD20wRyS6yqENzjs9cDMwiMv4
k0JqTTZ2oLJ7NLdsSoR6GWWmDSIKSDBGypb1pRcdAwvxf55OLmAiHywYwAB5WWER
0uxZp0sMBMRVrvDbPZL+vYyCSto26NAS90LMkjbshHyh/sWpBkiiew5qurUMvDEv
bIHDfjIX/iaU8yQq6YdOYRCX22Juv0YVKkaxV1f3KT4UVaaBcUt/9uaqo1uz9Ant
RwB+MRxv1VIfpLJqZTivPLnpmKFEzkn4zDwdsy9+TpkS5I3VRNG8vsWU8FactR7A
fQ8vPHQiIAYJ+FMpZGDjbyhEJoS03bXU/8mEKUUbXsjkUm7mIvmAdnwCHZkspUM+
FMI++ldnSQaisk3+7wK13EIYcRbtydzoSZ+piIC6say3kPJFG3NopCZZ2Y+XpkD9
q6G2G7Gwh2hyUi8TzSF4hfwlQfR90XbE7rDQjZBcRYD6mSdk8udyp1L/nCxjSaGK
6I516+L64IcFYmBJEca7zgYVZNfXv+j/rfpeJimOxtKQmIDOkDDBRzv28Q8fxef+
kf6qUJjR4F3axNndfOGRQOpDh3EeB01QmpUjMfcnVwTGqn61gaZkuGT31X6EBRoE
/DIpvue8kCwEKEnE5hnBLLBWxByAnfXvEsEPqnw8h2bOqH3g3yTkyGUo3lpdpj30
KZKw+U4LLwgVwo4XyOP9sQ==
`protect END_PROTECTED
