`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjUhRCwyF0nxCB812jQBfEiRDxZ0EF56h2wuo27e8SB5gXSIynjN3cnW1fppCBmN
N6QZ4a+pgObSMbGR7Ud0zvGVwY9bkLg1ab7I3nW9+eYskPWp6jNJVygVQQ08Q9/K
baAhWTeue87AlSskWmfmCQ9VhufrnwQ5S2aBfUDPrcXrgPN+JrM4t93XmzWtQ/QI
meTYBR/CnUpp6XdEJfa1N1C6ZE5shYKmrJd+ODVAWOR1+Tb4J9k/Cgi4ErD4xS87
KD5jkbwOCTE75GRCB3yHAc6CEY9v+wN2QQXK3cgr//rCEWDSTbSPO2yhztTwp6T0
M+OpZOD1pyVGvXo9zORqLjvp0KHCljhp/88P2iqiQ1uy3qq6+S3BragrdpFQu61u
ry0WJHhT6+5kzN+9muCV7w==
`protect END_PROTECTED
