`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AjiBPaYJjkibUUCpRqSh49my1h3uKCSx6Zy/1RQf617SkGuMV6GV8RMNDdIk1ire
H1pwaEIGx+/YYPJNS1AKVd2TkP8QEajh2CLkkdmsNn9i/PnsiJpk14fHX2wkTGrc
6kotGoPjAYYeZ3SYVvlzb3VZPFoXyiSeDkxfjcsG+S7Dt9/95bO43JQfwBVIbpNz
Bz8aXWe1i/2Mvc15OlhOMQXCR9mlyUurXly1OIrCS5gBLDmkl79dYS+pufVq4qny
tTe19/OXeoTLonn5IzLBEw1mKmMl7zDX1bZW9x7ZBjjhy2a681FyPv8WAjtNzNRC
vM1PHrbONj5IBaB8TMAdoSaw5BVRkry23N5x/K2MGF6oUPcbuQSToPLtOj0pL0Zf
O4GOK05ygI82HeqnMRvR0Q==
`protect END_PROTECTED
