`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7oWPpQfBiFUBVYkYVNF0ceiyryojxLysrOILpw4V27eIck6ekdduuOidZXZa2Iq4
rlE4RyB/NpeeEnDXxQ6H3ps1DeVUiO+9cRodStXvB6eHWQ5KqLOQbB7sxRseg/r+
yj2CSoj9fMrXW0UKZsK6MwPGeJAdPlN9WjiPauIkoubdsHqI6ZCM+TgBIlcj9pKb
EW/oQBH/PPRm+Z6y5aGM4/MTNu9WkJCvTISD6wjR43bhZ/QSRtY960ilSiA34l56
v+XrkqZENpfOeBCuFXGR6AZUFUVCcbpNM8f0CRo0Pc99oM3wwtjDRwFrV3BMzv89
WcoWRWecaXQm8jfl2lIk+5oi9k0JIecRa1FH6JKqrAXaQsITkGdo9DJ+YEOcg6SO
+3NF2lgxGXWzIxKk5o7U3meoYE3AiJIfcoZ0b/C1LRtcDTUX2umzZT38wldnd+wY
+4kV1zr8eEEbcTRYtQJsZcOx+I/L2glH4XeTHYJSgqk=
`protect END_PROTECTED
