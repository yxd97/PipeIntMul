`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8X/zenwDPCH9mytveErkMJEUEROkO0g2PoUGGZWAzHSRIiFLcugWlR8xiuE9B8wc
C7ISIbyW3qaRgxMmFQ4vCSSePY3PXE+/2M0cnsh5w3czU6Sqc2PfMBoH2c+373Si
Su7S6blst/Q2CS21rWsHE0cCNLakoEK/63PeZna6YZfXEbSuZXspLH0ja1w69kyG
te1bSVpd/u1XOT1ZLtw7nsQhC/R35QSouC5c7zwB0Uiz2RioJD0SQ2x1wfrEbodU
pHWX8VpzcsTtgkX4DVnSflajdxiS3bTC30Va91Bd2UTbK0VMs16Z+OuF6+BYt8qh
xJR4PmCWO4B71wHkfrtQ/HQw11z7b5B0HteO3becPtw+cOTvXp+WTa260HcidwPj
1alH1Ifku9yUQX3ikE8xB2b64BjwweQTafGwzWKFG5yo26Ae7glnae+8w3sfUwQr
5yXNtfHgvoYuYzYHmhdm24cttUTQ5IWXCFgI8vCsKO8=
`protect END_PROTECTED
