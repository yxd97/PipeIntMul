`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZZEZFDRd/vUdK0tWe7oKve5+iIY/e1EmmfnmcPHvXLSoWBM+nTU5lrfwcAfObKn
0SrqJOOjwi73gs/9bUXjjbuEMZnSJNSSBJ30xu/pyyWMe8O32Y7JjOKI4x92rszs
GuM0vgqWrDLj3+1Xsle6hRLSoNNffS0+D6nQ/MHKPZqJ0HTXikaBfgwwGGzZhBag
tjZwLvA4D6m6aQrTdFrboipdSzGaFkgyG0Nk1S34w4Si1HPLHBGTG5UbJTFTgruk
aq07afwXUBvNJJaXShr1OK8ebCOrVLzm58AcxDBDhRc15UcjEV9LqMbxllekzCZb
h8Cb/RJOfMYlJ81a5tG7sCOyCTc+Lve0xfQW0zqpL8QBcgKs2mDaYcWqIlByRYLr
IW0j2TGUSexGfjo/pla3KolfenI82i/9wObGxV0IcVU7Zb1ZK4hKoi9QpTHJYFFq
xAuZx6KvhKN+W9OW8B0fmcPT9C++UEYi0TchWFK4vbJmRm8DXsbQCy5R2A6TLGU9
UyM1AvyflW9qki0SufU0fexC8ZdUC7Q4Gs6BhYHGPI6m/w58QIAxPgnve5WCYItW
1AVflwif6uZF1fdHHJkchuAa3K1oClEeCCjCoV3Vs20=
`protect END_PROTECTED
