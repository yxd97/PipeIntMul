`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7TJLGNY3Qg4hvHfLTUUK8fIUplV6LJBf7s3TkoJZBWnFMR/ZjXmaSpRk2lHn3D6
OEHRH7yiSguup8EQYaY8R5k8UIULCfbHrqnRklbgKh21lL2Oedsy2Cv6k6cXUyBs
71iMq/MpnF3kssT9B5k+2zTLKzk6H78aOauhu/Y8isvT0dtqNh9zKkawMTVQEx5+
sMc8njP7KpX5Pg+PH6xt61fMfroiWWnmzI8PsNKiFpU9DyFz5BGsWOWeJSZI7/E2
jqjk52sfYWWpGxThjEUAD3MU/nEXJU6g0BrLOhN3dDI6WwNznsX2N+BZ6sdl2JM3
gpx/WaGhNgCqfmFORzKfWwdQzTkWrKDeqw6uMvdV2djOY1uYhclhWsVFUzEb5bBc
joKDTicdP/Xs+yRQgAoCLA==
`protect END_PROTECTED
