`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/SLFnY5Qbg8LhXVAObAOw6NaYHmsUypfm/Sk9lf4SxxDSyYV5D8YllfKlDQ4uyBT
cqGE3OZqzqpIWEO0BzdOQke9rYe/SpinXw19MYaE8/OPO2viFx5zCZWnEOexkw+E
dz0CAqT0WE++7IdnRFK6AZHT2Qqqq8ieIwc1wxl4SbAu8tpNsl8Y/lLsDms5kiYz
FUDs9EE90Hm5eTrUSuh6e6wTn+L07uGrjyyUERog1fsK/ANsuq4kFh7axncofZUc
Rl5WKHDXpYdcMOvlSis0RSRyLcDoeXM74+kKLMzpQEpr+l4H/TBibP/vO3VdyZiO
FafBV5ntI1Nf/YpDbrxcwg==
`protect END_PROTECTED
