`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzmgE3rt2Z34HWrvgoKW6pzwg9YNe4Kazdy32PUMgUGe7rO4Xms1R+uBWju0mTF8
0TEA3/HfWXLoXIcj21vPJiQTWAncdHHmFnoYlYmtReCFgnXHTOrd/YYkTNaQO0d/
DNH/kDxeris+wTpfnbhkELOF5TVhSQq7bCLaQnmQDt2s67qy6SHajGnXyGBROdfe
M9ref+4SfyrBvqyg42e8TbXec2+WXPnqYSlg2cF0atL/bjJII5Qy0K2RlOpvMF8J
3DUbT0hN9aJ4P/4QRgmmwoDfeoWtpyMGCNar4eoyC8PEilyTJeTmzzo0Lcl/+mr6
2ZdYSMTG/laN5+mk3EfbEyCsPsj4jB8FZIWVjf6v5PKZHAR4hjha89D96fYVqUMy
GuStRHuTLC8EiyVBbLBGw3zoWZeJ4t1rw2rFhQ7Y13uMGn3fvd0rifvBUsVL/7YG
9jk041+XhyajFg15xs/8SDzT3fA16V/YOFqz/zYdHG3YFC+NvIx6fpIj/uaxGiLm
wmylVUOhIpzAD/xkU9wf4A==
`protect END_PROTECTED
