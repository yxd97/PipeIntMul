`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9ee25SfUWBDC6HLq932zdfWiProuiKh6CeXNug4wpOr8aMa8h0uYJMIpXlECWKA
LdFjEfXFLhz+dZWJAOf5yPeRaoI6FXXuixHMtbBbyzVg1KpnsdGvxm3GVnDMWPYo
/7ljClA6N3nKTqj9vBXVLRDNGjLUJBsJxTUKN/NU8vdWT+LntNP/R82Un1SFjmS6
TR8hPBcSJR46s/uYwgHS/rU0mpiZOWn4Nlg7d0Pm3ogEN+xfoLh4lbrW4ZFQyc39
N4f5wiA+baN+e9lj/wiQetm/O7XO4g7O+/J92EDLbGCbNZkqZfi7aS33aN6FeXbM
v2M3WG2k4UTIHSpkYdIgQyuF+SNl7ffoBB9vZtU4gk23WxjmSuYdPbIHcHDjt9hl
gnk3+q8qJTsE/61zUwaaNF3XQgzEJrijrnl2h9mPF+FL2EMoIT6LXbKYwssTIkdj
O3n/ee1Txwy4/D5J6TpgTiTSfUF2gzzSTAea32rGwV1yD2gO9UVZJyOJoR8iWgdp
PdhB6hhqQdOj/UpGPR/xUlQOrmoFCjTGPDBQaYKYkM+I15MYs/s7Nwtm7CM4EeqP
MKmw7FAHmad1qI2bxEfJkrdJ8VSnY8lutoAzZIEmniw4A4kDut0jlIYr1uf8X8YJ
iCP89z0aLTogQiGeMZspU+s+gdev8TY1NAEdNL+rsRbKEWy8sQJfBlwYi5YrFfnB
LtIfp0pu/GUYO7t6ADnO4aNZXwRE1IBm/CgPgDD4MAWHZ4JxHAMQ4aclRnckWqzY
jsXHxGAhiSb73RN1jjdVtHiewxybKFl8BdfJdQS6QX7ZVvK2Ti8h8U7CR8ktISJB
NGJYdozj0t1HvSaBVGJuVpbJXEDEFIzLPAbgU0o+vmwSKUyedGVqNi4X9Z95hXE5
ITIRkikbhlgGF5tHM2p9PfKnmBMwA0vptE/wj99tCQjcS1lDlpMGe+VKkD05jFFo
SkQrJdly9bM0yVSV5kVV5bW65NC8Bc4EtEzHgI6YJvdeKWyha1Jf0Bcr6zLqwyAe
6fooDfI3IFKX05/JqdFu6h1eRXwiRRLbYP4aagksg7pwzfhsCvX8eWfSlDWeskRT
VSxzrbo3XtVqaam3RPJV9Tw0Q0fecwcxZ/57jbuNPBAPdUuaSE09RaYSR6InQF+k
VKzs6eFDCxV5SePtXpKZJetyY7tY3PigdkzV1LEZTKLSIWM3m4c4Onz/uTuMLTty
LRuufMUwUQ4H9NXVtK0roHO2eTwg05KZryqol0t+YwOcDIR+dl1IkL2PxuVDPjZd
qbAS01gYrCu5GG8X+843m1GvdxddIIlN/fV3PiL8iIfBxpy4zZvEvP/3tieO8Thc
bEZkWw2iB9gQzh4lRmS6NGQHfvazsmkNVrBoOGfdIojQdqkmTDt8xbGdvfMu8W8W
cKwlAvv5OpyuZoNuzgLB7Aw9o3p2Y5iBOVdtj/76X56wwgypNfwMSekM1uWKw0DQ
vhMHydJnWkjg2CJtFu9kmqCKLhWQqMx8EQlR0AqdOucX8zXqHl2LQY/FohZUiIKr
uf2zFcqsGBxar3kyIrZaXpiTUhGbC974SAHQHBbWHMUOIAjYZqR4REWb0WLLIe5a
L0AcMgQyACrkah+aCVkwiOVVO7zKSbEIZBUGQM74tkdqw+berJSZ8jeWhtObTpa8
OAIiF3fyEL1aZ7YvIUALrJJKCQ4TtENTykhkQndfJVAVm7uCVUfB0QjuWNhgSviB
wqnsfy8rMyezog5Qve6n6+WsmfEevm58W6xrTmcwetFOYEVKnyMUjE0XkX7xiHMJ
PuCsfqOofsEWds/NDiqnntXjir92/VMAIsWkPhfFhEltuA+Tq9FUTIExGNDPtBIu
3QCTXY2QbVH8ayBSaKjJQQKVtt5UQs7xUQ+8i2z/yFT7+JR1FlQYlI4J+K7u49gQ
XG5jV03+18iOjmbKbEABexOyunBDZjjPn6zzfJhdi6yH0lfegy5i1RYe3D6BSPCC
WRr60CtWNrcluiOeTWsDavTV0o7ExjNSBl3NAxlc0qWM3T3KmPq6aOADFjLuyX2P
XQ60x13tc1zImea79mu6vQ0uTSBpQ+MMzD8ed0tB9y1fJHIUtw+K8i/jnxz0AlMN
2OrbSWVJzJBCIyVTrzRBmGGmquMMULiNqCqdCDzFpTj3LLMLwM1dyRjqJ1+RKH7S
6IyLVhtbHvAaywXcW6fGKfEnYYGoyQ+8Dm/wSbiVaw4Efic6F3SpCuusrPyA1XqS
PkWk54QYTE0iLSN58/cUdoa8p02JbYw1NfSretmcc2fc/smaX4Ry8ia2XrkfBZCK
0qRh006U5y6y8JL/u82XRCNGZVyGvOQ4xeHroz8mmjjXQhjZyJwzn6tgH2Z6niJ/
nI7lqET2F07h5hlEmXx9zOd2yZbAWK495OWh3H8fqtz8aATFaOZiNb+IPx5m+/m8
75n5roVcxIde5TR2porx7zhKqE+lS48KWAxbFm3uQNt4am0mJJJ5eM8YzpCf505P
9DTvRT89dz5RDeU+0EIUTOFWOEq3vR/IjSWzsRxWtR0SikwWgpM3Do6+zDxABy1T
gnqp5OIYPkHYvtBdxlf6DaMnCgmqM1mCMzM/TNvdoOXCSkKly71H5nfyzm23CHxN
/Jru4GRQYN9AJakchKG5pxNnV5o1y1zdEIJnllsPXreBqt14OcCVqXRMk+yzAtWm
N3X+r7LSAQYdQNgCv6x3BGFbLVygO8SUkd5KVR2x9Pv4t3cZ0MnAt/pYfArYFrd8
x5jrstl5DdwW1vWvNm4n/XTT3+UmJOYMJT4509jkbS1VR2s23+8b/jvXNm6QuNUG
1zTRwd9STBYmn33kNEhKET2Dk1yG13WkzIYOVc45f62OCWOx9U7gCUUig0ppB3R+
CZRMlnS/I0oIWn4vAYX1J2aCOE04KVgjlRbSHdVRLL6ss8SVQ30hvBEXQeWY5pUt
MjHSYH8DaSL/QhqDAVIaytfIknmsnQCa9TM2RBKvHwS8dsD2p3TfRmcH9a5A7V9p
UJisiy8iFDMtgtiGrNe+E7YRM1+fBFx6Y4YnZiW281jxM9y8hB+felHGAJ26JZRb
A9stxThN8cROLUArSsOubVdPj3hm1FULHoi1YKdgr0I6NqncC/QJ95xXQB90ogc2
M/yO+rduZ2LewDSCIYkiHP95z1l3fJgzz+HeFVArVomg7xJLqQFCqvaxOYNfzRJz
437eqncXRpsrDl/p1v68FEy01fspp8maTlJtqgj6qAflbh6opcO+iUG0Nby1lbD/
aqLtwKoxVG/mhqYsAbEN3KbO28CUFA3EFGR7qorQ/nTbSBF6a1kTviLZJ1s5IxRo
ZnhcFQGMCIEaeEvymZsKGbq844CQEFjrErs6dBxe3o4olwYYTThfj/ayVWc0MA9k
HCh7QxqfTcabXzyduo9Mrh8YXCLyE+0kaO9J5rW+Ago9i9PoqNrz0alSUbQ6BJue
o5tTroEh9L4tlFSXxFnx+AFnT9xtdnfnwAWyFmfhO4HrZRxtDqxj47gSM35FPsZy
FL6+ZCShKNKXr1DXyKrFnUqllqTF+l6LrWZ59gu/AcTOj2Rmu8ZN5TYivtRGliFn
nLDDfsr6RIE/hDcE6pC7EGBnkesDTsTGC2ay4n9V1AOO9d0z12+hyTZLp7wsUQ0l
VzTE4PsQsc2mnMuWlitNdoIzdwsKrUnVu5BbvGR2Fk0XQay+kL1LpMAghlyS6tuo
Gvu1gkvq1+REvMruefVhYkG7uuNiUyy40XY/2AL+AhJw8e1nC5lrI+IdjsWW4zxi
KhxxV/41SZm9z69sz0CRikZ7tzkIIbm58jbfMIFVPIaqzkaXlgfjkuhn9GF7hBD6
bEiMNfX2J/jyYiBIB2PWrepHstsst8dPpOmSYKkuPQInr2iOSnGKTCY2SdaNjvPm
UDNaQk8sehnbvMyVBJR2g01MKxqhdmM/OCJQnEBo/FWrZTzA4wnMnXQqBlyuqVI1
tpeiL6/8mfFWJONkz5NOXsVtRoXMm3ohDxhe+2+lQyg4PNsrW4CZeLEqygqo3Jkd
oHRaO2FtSM3uGYQujW9yfXsjuSYyjvfzL+3ohzlhthw3dpkWtkIwrj7RTqV5BN8/
qGVsxaLtvPctSYHg2lqnjUo/Mk3vO68NoUORIlZ8HrLTb7PDFLdYxGNb50xnEkyQ
0OsqYAuWNm30bVyyBItHeLgNVlpGo9x5aJyBnQx/OyhyRcIYVNl/2TWDi5zmBbix
YvD99wNj1cXyywKN0qe4js87bPXA2NcMHaguL3ZRgg0rlniaaGO4mr/CFIgOCHzW
QcxrqKpaOj4ff1bZ0XfpGMd4/Y5lJiyi9GBC0eoEG5SSik046JxWBJXonf4jeJz3
oNpYRk/FuYj9m22c093mnvDNAgPvWTydl5H86ykUoS6l26JgEcr83/CVg+aFI6U5
Juh3xriekTPyfFAm7g+Nzt58aQgO95FkvUIlE8mZsXtMWeltPRF8kZSes0FgS3W3
zZHodh2s/U0h3NvDKEz6nio04D+n+tauP5R++n3I8XrR3dL0B4nh7vhsrmtuCBVD
tDWTwr6XuXP6ntKQw1Z0qdF3MFxYqKiOeQ+OSgIe0fIk4zoqcCTMhOcgYOpofIHf
Co3CqHIv45VfoKSR/ZPehOipnzVeM5/YWeqJNDW0bzCLXK2RuHR9EnURT/s1HdNb
8bC4KL3ExwNvKgYhwg1QTG389xVxTVSGdV2JpjLFPS/9ozih6HFDsIJod2rXGl+/
6TF/T4kbwj6CnzQGcZYF/vtrCqBmx08ntEO/QFbtvIBjb0QHc6T+lZHb/cvBYvQa
MmOeyABPvn1F/YaxLsdFDa/fsKG1pWWtHg6mwqafEHQtO727XpaihMWXf3+NxiFn
3l1A5+1f3mjC5WZXZUwyqRJmC+HFuM/Z1T8HNLlWMRmkn5GUng5aJIkKLlLKS95x
usktwH2TXpCJ9GhyV8slau4t4kSWXlbMjfpY/tvd+RrfoC5OPiiiITUH3uyVLEj/
ECAFGrpo/NefIYme1j1NAL6jv08MQxNabKhoZItSFob9Qwil/ouu/TR5VnCbgN+Z
Sk038PALkNh68WpCHz4ekDrCnOnG7KkqRp9l/JlGLD6BAwdzNlmSLFX94EvtnkNQ
/Bk/F32ml+OQVO9Z3Spy0vA2Yov3g+n9JZX9htBO7TUGRYBThay/SH4kZ2EYxxPC
29rdfLmqPclTXh85CBaMn7STlcEvLUX8jKiwckaAAll5JQdY/PSXlb17hfCln/98
CUzAfBvKTr1XioswzAFo6CpP3FX45p1oCCKTXiqhXZ9IpCpyN2yrAKmghEUfY20t
ZRj1XGPRpj0uRpMMyAOrXcE6HLNN8750CbaU8uXQ09LIdbLxPTbEX/xGBr8gW8FJ
8QRH2uvZ5ZnnVgAhxpW0PoRiDASp3kKtEtR6hIhmU7gA0G3NBwPlzaOXUFeOu7ok
DFTyfxzcDk9/CON0LreZOfhRiqC1jiHCnU6S1R4wKgtcwhYPROLHJTEuXbORwXCd
oWX6hUP0M4lRb058d4HoowfhsGX0uhLycf8vt1qcVVkwVJZ2+BXczt/bvyVIiVhC
iOu44DUrkrv2fTkevuxsSDLxi9tlqiGdwFnnmXXXgvdZ4PNB3QBk0JB8oiDElfe+
yAo9/pu5KBnF/G5hAnHfVN/IKjkoJKjPT9SbVWWD4H9B3614/8sKx3MPVcYBUGxh
TMimjXSJEAB5ap8nt32vD06KoairV3TDZke+gk3N9Pq9Lyk7TUgWsm9ZY53RBYPh
ZmB2r5figexFYoaq+GM1Z1kk5LHOf2VXR9+L+EI/YXbxBr0osQiGyzzoAC5yvGh5
T5P2D0eu2uiPOi89tJ/Q8yANTIGwDPxYS5fqn3ZnefCX0K5OgBpOh7WIQf+FM61/
Osuv/uQL8APvcUmEXwkoWtTHjNfTlN45ZzVjXc2KWrx/kyXkKFLbFQ6BldXGF+Gz
q06znDALA9j+bwsnbWUW5X4cWlhR5U2/WSpfLOMdKHDjHW5T/WTdJB66Q9P9Ilku
MDnD9IhWScXqNdvQYcw21NUG/nvhiM23FkGXwRVJl6T9/UZ3fkSY1voqnZJgsp0l
L3uQO0nCJEKC/JdoToIvIw8hfTng5FI9gyDU3notKdrPJ9qLy6KVcj8Mf2Thz8ND
ZocMO9VAs1o9Qwu/n+7j69fhlVmU2aPaP5TBQoRVMR1MWiQK91dDcmBf41XT2+FO
9wFUk1jGyaSE191YAfSP4CVgejKQ3bcG9B5K2ce3tKszMceUS+4DY67uhlkYG9So
V3cO0oTeF9qdXY/vQ3Lbpk1UK9WuHOtB98M9ixdMnnv9CI1ON7NyJsIrgsmMfZbr
E1RQWpCH+2P2FSy/rz7qLdJNv37nVKBERcFdRwY6O4FnqwY2yXT/amU56SV5cRWZ
7VG17obXGvnxoJ5mVhiEiKlhHUOYQka03F/YKG79yFFqGWES2HGcIHPpoikLLiH8
sCAgwIFy4nv7tpKtJwhj4jq0yS7o8qscaPCIVvYxrL+I1T4DdfRsuz58O9a0W4c8
b8kun1MD+HcQv1sDfzFGvbusIwIUX8AdQnYmcAKN6ywIctO7OC6MBhJaEbZ4EaKw
zE4RUPy7QP190yToEaRlp2ZK82VbL3K0HRGb95O8a7BLT02HjPCHIoyKQuvVcJmV
cBVkqgY9Y3iU9DndsSaYSj8aeWIZ4C5kIZHqoxcv0yxVcdxheAq8Qyd8f+63b1Zs
pznFSCTnbjxb6F4N7OVU0S/GmNzCugHdFX+wRfsiN+GbJqTOI9OT4KbV+1AWryvD
sRlYALeWVr18dIam/9V5rIjKS0cTKXxMc6sGzA85ZIkgqrHMr9GISwaN8YTd0vSJ
yCQDxXOx+r0Ylw2P/sgf5ZZ901tlgSzONPiwHN6j2hD+tMSkH3qnyBjMDqOX0FAp
yIaDsd3gHzekXIVxYlu9aqaWvzjaplPT+HfA8sdAQ7Q1Y696V7DgIGPmcOhEVPw7
F8rUlfsCU+6l3RuoRzWGiW3LM1vJTtkFmbNyzhkHlF3jAjTUwmdFG0/Ts8e5kqKD
/QSSKkeXidftH0uoMMLl+ZNCze4TCoXv7p92qc6LCU3/vSaqC3B4ioBRSrWksS30
WJOaZWUhJHm2TfI9eCYThBGtdfreZ/YxC00+P3Gf0ebC6hHtrzhhL1qoMZVe6Po6
M6yUQfcijlGivYqW57iKoyRJ32AGVg4l8a+Y8XiP2hW9vu+O55m0ePp/vhElz2jF
DXkFK5A1HpBmuMJyE2GdLlVwbO7BVmmot3CsJ8VkAO2EPIELSlVsWTX+LE1foN/z
Anm/7mREGnjVAM1YbhgG6uHhnAm4cS7mrtu0vcH/mw0QjqOa6DPKt43FN6Q3r8OO
Gi7UW7KobD2k5p5Op5XFP/hrSOOPLin8goHTBrnDZ9C3wuQWdOiQpunplvGHmDab
5XNV1OS27r3nOlmrTzBMq3nt0FbNVsmNv7GkbDK0nMmKtAbzahC/UYM/zIj/8WWI
Hz3SMPUwE/+CK0oqX37Zltj0fFFL9BB3OfJbB3EhgHM1kpvJeVgwpxOMjlQn+Z9F
DgH8T3o6mWc5BAw+/ncWSYuIqk7r7zV5r6Sp05UiSaYuaJh7QbW/41m9oxFzZWRD
AeE0qbJaaKEbo0BVRbKQzt3m9evBaHsQAg87x+BO+BYn7Bg02Dk5w/yIDFBFcPAt
78le3YQ0pmMqsEWl1BCyaSB6216Ts9W2l2OcgU0I4uDNAE6GaUPq0CrPtjNXHvvZ
5wF+Z8WfPmqprpFbN7HlwS7V4pZfFoXBzndWufcCbq1OxB/kYfUyPC+HwhyE2pNa
qcDdDXr8LBZ6T9QRSiD9dobzAC6PwsqGFGsYsY9edKWze/q6H0fD54qVXcFboFB3
DtRM7syW5NXdzrQBgffUng2TTwbBvFz12emsy3bzaCeJ4qN7ZGdJY1TVo8b//cAD
RYOEdy/teLDB7jC5k970E1fpLCL2Mj/jc0wiFRMwM6QwsuolqV/N5k45zVuYA/HZ
9Q3qelbG2FXwYvDWM2f4V7UkTRDtNyRbZOjZMyvgshkN+ZVuvwov0k4wFW3uvxJ6
OgLu+RExadjXtcwRRbxMzE1Q6mLcuP9bezjnmJfIh6KpkU4xl6WvNQBdz1Pmaz/A
KgRNV7epHuXfPan0ES9eXJ2Jo685sPe2Cd3+uZkzrZeaz8H6O/MRJ+/FkpQthFMm
EhtlwQggFVmcZvoZSl5QqAJ14hTGr2KsFaxqtf4z50062k47MTWoNrEo/AyDMuFM
Uz/lHZVHaxaAHP2byVIAfR0WP2hptk3AaKou5rWtMzbBvamiJtfdsHtY7DfKE00j
6nCA2vOEnee7fT7FmHgbLPNPtcb6XTUbgOQDUctDXGiPErzHPaAuiW7vd7DmkbTh
bD04sroX6DlUU3n95xOG+yVgaQwXBwsnlwXRBDR8i6KRUCznsUSdNI3QCCHwXiB1
1Ll8usxGhyF6hiLi4cYKNtglHmgw3AgYEsCF6eu5LVsrZK7oz2D6LUB8Dap3ji3K
DHXFiZUEjTEwN+vUp+4yyjU4uPZ+mJdt4ufFcbF4z49jSW8nXL9TgwUjH2J4tMbG
tQfNKLpbwrJ7Vzgyu8xIm1/kjq2JhYRtMi3NBg2pNT/OkZv8HnGPkcW54DNoznfF
xr6uJ0pu7zxrkxwxMpzXk/+9zd3yVgGB9QYoyvClYUS+j/Ib9dgLFPjtAcGe1IMQ
3Yw5MRlEFuSyKryBBSCxjC8dhLT5xturt5hOV2Y4D7xQT/J+r34EaGP+2jytqz0F
rKJqXT2KHrVoovVoo1oj6Cgz85+NkLteOe4Pd7VrMXtLsBGQ3Mt7rhd44BpxGo5Y
oDrcqOVGNXqKWSf92THyIMo5/Dkg2X9pluol1rYJIGuQ85xkTA/W5Dj/dzZUPJsi
tyvDy1uoUXrO5UgyoN9JRFKWpTLGeK0Tp6BaFqeJzyvCoNDP+5SQwr/FAmcdUfHx
n0rG5MU+GKsTK4aPfrV4lzYEDJjxMU9tzUG5TGx4jipvfxJ2hpBpTIWwDSFVvas0
W7WJizDM5Ol6w1lXZb8wLvime3dWblHu2yQfAlYz9cBw5vZlhNPGhqjb0ZB2x30Q
mTSxGPqSKXQ+x3D+71pKmoVOpNd9p8oxlSF/nQbpcmCicxk/IkzqeQlc6Va4k3pT
K1VQlZYjAtNOUCBzhRa33AnMTNifs/KIcX4JRFbX7ZcecNG/tLjPe+3Qmai54PMT
xc1Y4RCtCXwJG6UO0x+12hgFJDMhQEhCz+Cdo0uxlStiVZoB/eY4C7syyWszPFdg
MILMh6ooT2phpTvxDnLUHClKzUEYI433oFKAtA6BF00K5kzAij/C3tJZs4wKd/qx
SKe6bePKUwJmauOLfpXdNCDvipl01vL3nEe4TyGiy+dJ4HtvGhP/UZfMH8bh8Kq+
6RboQAYhpocOS3fqfin7u57qKzw8eaprt72rqbi74Y8ZXJUo0hQB7f7Z8/vrIijI
FN6NB57YO+WKVQiY31AfFO+5IBsxhaZSdwB/QAcKvWQ3HM15WS4bZsosY9LxLV6Q
WewSejX6D2/GdcXp5pHeOTRilBTyn9ZM2oeHNNuQol8kjpXVFEQpNjj1+EPBa7ib
iXSl8vFkbzaclcDRM4x/86OvMeuV+xAe+t+k9g3Um/z7GFkbb8sGxYWGtPGSkxes
lGLGnK7Liy3MYWSt3J5rdBCSL/dGugrKfGLcwHxkgIL+cI0l5Vp2lR/+AjO93xYO
pHuYhRO1UzxmwEb9ktfjTFQGroluJcEGxkwr+8nMNjP2T7P+ExzfgVYII0nP57Cx
EDbZOvZWT89oGMNZ8ymYqunGMnFtwQ6ugfRDrqvWnqK4cnj1IYR3SRr3FRt2cuQv
6ZJg6U7sUtjqBTLLxogDNAaopaYtrtCk0eBFZE0fwo3IbeW4djSMGdAcRnPK1Dw3
Mmo6kMRf62hqPiRXeppM87/egZnYDO1b7cXGqrYFz5pv7sF4WOOOIh4cs8K9Zem/
zr0oUQZ3hvSdZ6B8vhYXsakXeN7KF34Li5fH+pHECp1DP1Md7wQ7J8JvYclS+VH5
d9u/uOuhQ7QDso66LORkwMrHJ7ZyO1jvOrtTrF87TiT4xvCrjwihDykNIeRO5K3b
0uiJYJpsHcZZDZiD9oScjeuyUzIcr12FV9mnZjZyVyxifs8GdFXe7s2gPcuakxs/
PMacgyLOOI+m6Ut4d/NzSrVOB8yrjHfVVNdpgvw/6Iv+fqYpC/LrZI8bOLT6N9Gn
HHQzfS8SZdFkjw5FZEqDoro1R638Dd6x1LYXO4ctnYoN1KfkZhm0p+8t+6+h9k7z
20x+Spp44bnfVdvrnWXBZ57r17yc/GLRzrFD/IyqzMIht464ARekQ1e4R5SIT/mu
nFb0G646zdEUCe3QcfA4pnDRNiv0IKHD50bpYN2GIr3qUCS96nmJhFWUvbovmZhQ
mwuZ7dNIx6Aeg4tC4SPD6fEzmUcBrdeqJiHWs7c+e6PdXrwENvlk/WZn6ZUJ4/MF
Hv/CB9uhXQtCgO2e+QGbKkdcRYIt33QTBJ9Mzy+xEXRwp2RTNTuprQxJ0vK93FCZ
UjLascYZkTWx0W7n9FNzawQsLj0KVkJfaVZ7OVIdx9qHHIHT3ZEwPgnAA43OF0L3
oHqyP3YPqVcS1M/084nh+NFU++/CIDzS8HfJMIfYBwAZakYne2fNHWKFlkWEFKMG
Ie1C65S6AJX1M5ksmRKKfNOzpakznxKSmnRIg0Lni33dsjayd0FJ8Ht8a3OUd9gM
UvhJ/saGByJhOBYD3thFWf/pyVjLgcC9Zhm0A3AR1g015UHTYD/KuIoSZMkajtx2
xDvgxJcxv45fB5Ve1i32ACF4jrC+GAdGREFoTNf442EaPgI4IMqUWF4Xh00qK2Az
Xkg147QnoGM2bjM3j+wVvMl02lLTM3kLbbEQVwvKFcY39kz/p4kxse0g7edo9+Mq
5R1My/MAx2fpc+nZPEd+TI50BLgLzd3/sR5op+oWkOyJoLynhVmaDNLnrQqH2QXM
lnx68WBr+XG1eRJSi50M/gfvnf9aYtCq3zZVnVEC90PSdSxdZBvEeTCybhbFl7aI
F9LhO1I4ljACNN5L8xp01sxMoZQxlhCcj8mGgkI8e4PV+1U7G5zIWlrZNocSPzL/
mpJ2EeLcLlobJiblftKHU+SyGSMtPxz2r1ncoXj6yKQoM9ZaRZp9YpcFftbwnBvB
8FZCkMxJSRKnJEiFuZZys9nGjyyHXujPBwBynHh+fuLWyay7LzZdH5hta7BDtt5+
6JaMPazj69BXw0gk1wYnRYQimvbiZwSCMA8VBd7V6XO6fzv48tsPDsRsQ5ZykTyb
8SWdJqMNUXAanFbKxQu9+pcJU1SBaQY86sHzi0oOkxa7VmkysYgaPgLBTztQbu4c
NA1PB7eleiRLOwQPIqo+Uyn30hCd5MbdfYhApcdQPR2vWlt8kRRYadQpyE/OYiM6
JMtNpfQxRVZhg+EaoVnIvSY9xIxm2LuX9vwvWeG7xImb/OL1xlq4I18mCl3wkan6
l4zNUYtI4QrIQfuWwaUIhrTNcdiDUa/GeC7+we5G8wURKSg/Yf9yHxxa5zbQWmp7
Mfw8JmLOsGaWD9H9NiyJE1wgEdbDHPIh1036tLuM+SsUzmqvIx7M9d41/BvsyUF5
R4JQ+lHVA8nURSS/XfkgNa2IzD8GeutjNjx4VTujGZpPgY3/473jkiyRc+qmW/pE
RT0tIqBufrT30DXOC/Vb5EqnR2WMUTzmmBLrM4N3mvN2bsVeVgfw4w7W8ytoAVFw
ltglP+Wwx6OMCXHnmJycEdwx/4MOx+mK03pBncA/LfZ7BjVAYRfVMt+AicEtDkbu
UqqtjJYkrUu5X5XPVAWSEeVwRKq8pxfv13a7ucYicEgNUZz0YYsTOQQ3vTkwKaUq
B8beVO+InYHvFrJr2WcdvS65iIh6IYZYbyDOWocfOtNv3Pn68PmRTEpDBGHrVy47
o06houO0I3oNK2lL4EfYqjzFhiGX/45Lli1OwGzJE0EBEK/2CfYrdgN3BLJVY3ot
BMVWDDr4iOctUWhqd+n0f9pGyt90cAKkkfX2QuDXwVzEiFtMTqwHMKCPFACcAF7V
kd2ViDFeBnEt9Q9w98pR4/S/Y/gThQXkIYyv3S2aFXwqxg40FFsIoF/idWZ1ytUK
GZqJ+Vcf9V+pSnf+WYaxJsQ2DMpdFPS2KYetnTIoGzd0ue3+5Kl/F5j+mY/dbPeZ
`protect END_PROTECTED
