`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2l6XaAtcR6tav8iC3hbcBtyAj9l2LOhxmhN9pmt/SVjDs5nwMPMrtpepfpgsbSPP
z1cAVk6yVDYTrswndzVL84b2e17Ph3YzkkPjtKWADhl+T24vpmdW6mVEeh/sq45e
c0fpX+mT1L5HSaSxddgMe5ibkuJezhGBYBoFkJFyMgC+LLWigVWehFIlPR8B6W/g
/Z7GI+m4u8kQJ499RNCUgONB6qyksFqc8RBQ5CB2ve616T8t80RsoK3FNA02/GAu
xaJnpSfjWPakWpVR4BXGFYp+fKKnz5BenmHbclR9hhI2k59zaMlW2aJ648GvbeMJ
iZf1z2r/lFRqaDVdYH0hrNKtfZv8dD4KjdbHgGyt3mIL7RBwPEqh17VczrwM59O0
/8Av6Mwtl9SEyMhagch+scHETNQVsySCtjmnj+rO3ZiMJbisR2d17TYMbIBjFeHs
0I5l04ALJAJqdjXqSvucH2Tf4XQnZy7OzaFscPJ+1rKxr6v6IPNC5v3CXoWl5ZCG
VCDhEAA1+vWRS6aGMH+RA44eFqKF4+Wy+mN09/ZrJ2ESoCd1XIZvfriK5cZKFy1d
oNlgxUg0vWagULfrdVbr7gaynJjA9veBTjoJ2AlaII8eV7lpIYJCqTlS6SgKfkat
PTWpcUnpFYEJicgXBkC198a64YSZ6o24jdEfK9z36kGc/G965yYMBc0b9Xs11G8U
Wb0YaK7kV7YtSnumbFOJnCuYvpdVOzLNKEmrRaAm90liNaVcEm8t0IJ/+wQ+LwGH
Hy6pOz7yXzDx2ZtJ2Z/CakfA5IuIEiXd42BoedlEQTGJE/jfhN/qJJ5A8lRHNr9+
Xu3MM9b/wwlRuqToPbhBxlb7RvIp8vVaTmaQYzOngS2unuCM2MtlWGp7cCgZg9ne
PJLrMtRuUqiTeQulE2K33UtCXL8Nmp8edc3VvLr0tqNWkYo+fki3tcfH1hUb60rL
LwJ9tQGhFQXq/1Qt4un4QfkkrxFUsVmbh1vsdWpn77372XYSqXoydjAc+HZxomls
x4XqdemI2NrR6iATH2rJQvqWvcIO2SNhlSP26BAKFMAALYsXkKuDeQMf0uXvYqW2
bPvSlgsRBlMtngr7B0yifNha2riR5Mf1LH5zjKK64CXeg5kek9p2fvnnPQyq6rL/
ZrjtzK30kg9NhkWTkezTl/JUnHmECoIvGRfE+C1ejvMNSGM43ox/DhHoQYhYH8ho
v7P7PxBqplogn8QnNosIDWKM1O4B+OOeXQNYcu15SkslBPUSvj92uiAaNh/X0pms
S75BwSlKmBaV23uYlkpIYDbHWwB+9GXGFvO5RGjx/xUxX90RK8hpljwWZy8Kehib
jmdP2GY+InVb7gk2oy4jEWDK9MbqY3MIiqJbvUMVfT4nA6Vjzcb80YAESrOF3i2W
xKJtCDgLLY8ZhnmZnDLB8bZIa07PxS3bljMS4IAIOCR316VU+V2NaNWbieGjuk1b
rgFTi049yfGYluVZsXGLayjZ0xTAxGmzDEKlVZxZg8TS1KpBuOx6kNnr6XMJ58C2
`protect END_PROTECTED
