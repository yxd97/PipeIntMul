`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IidLSPRLgndLDtJNv1CZDnl7U4gEI7KoPz9Mf+fAfjg9wx9hzuZUQY0jxiZvTZe2
GLa3o4Bpsd+p4/jDera4ApcdDMoXgHlPgnkoHrsORLlErNrA+whAnm/ic9Gm67nO
s2qRXPCoJH8mnWNHYqPL2plzvUmi8yYI7WplQ7VLinnofQwBekucaDIxHy5zxEph
+/gjWCM9m6schCqNLRC/j05b+5nDC3FIEaSGPYvDyPw1vH2gC2CqH+G8FgVxoxkR
MWgbi041zZ8bD97CaXjCBU7AUoKcRMT3vImOADzXcc4=
`protect END_PROTECTED
