`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xjJu7xdMWNgBvRAL31FWAC/9upDO0fsWh5m9IoqEQYHDHbPmksW5My3RUU+TSztf
4vjLn+XpRBtRY8BdemobImt90Pm/Z3+W2GZvrqP3alrf1owY3qL46USeG8TnP1gE
dbzqy3Bp9OqPeIn8xTSpQSIUBw7RHyn6AycVFoSswy2Aa7DOleDrRCr0wUfQYzuQ
hjec4co9dwUdz1B11+VQxAErkPx85er/g7+23WZ9qjwET1ibyR29nAfZDiU7LcPT
BK/KF6lDwG3ka9t7Gnw53BYoNylQBcd+HBY3aJ0pKMXkJsza1a030KoNe2JbWI5f
`protect END_PROTECTED
