`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwwZk2D+lHmrdkgUiiylcxFFUbC73e+La8UB/07cJJwc0n9/+dFmygvqACPZRTVu
nNeyhwBuaWSCTv2bfL6NTYDw5HQVOsVJUh6jbNzrvOlgTueZcP+BOePYeBLmKLjD
hnYOSM9a3c7RZHCkrxkB71EXEH6O67SGM1EwZ7yXr9/PKJPZhRmo7bba/Bwy27fR
zYp/vgKe0GFijxFt+IF684DzKBHsimRENIvyX+zWR1IN1xWIw98EvyTwaqDPq6ED
ti/o9EwFiMeVwHFXyA+bXpelfodLm/9cnBJWCagOKX3hw8IBKwfx0K+A07xqa8aF
jYAg+nbbd7YfKAaZ66hYM4ArhhH6xTVC5TXsB0YFXtqShv72fJsfPkTVwWzcDCst
4ubjF0rVJ2DaTEkrkc3YsbfQyJrAhPI97WdgblD8pcqvMFxFpWnPXxWvKjmC1pGv
Bh1QgCMiQSS9kW/0aqr2eDlue4fimXezGw7kdmbXJfe/84YNiRB/m//juCxp0pTe
`protect END_PROTECTED
