`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmpzepYxlMlAIFSmVp6t2jtegjnPVctt1fyySCnz6lHg47Gu1hR7bwiZornIznoG
h6pPxHFjTisVuGa7grhnVP5fhYhad+XSINkgeeCbheSjlKq/r/CmFEgctwni/Yzg
T6jrmQCVguvloc2LZQHcPb1vCat92o1+1etZfAOnYS5QldblZQzSgTJ7iVz+hlT3
cts5qCgCAzW1jW1iFI2Myxt4zN1OuJ4tUXQwc9U95t2Ahve71cEVVKu9NG+pmzKf
C18NE/MHzMwYYt6oFX8LArE6EVKd2/zLiWWNoLoVH60PMkdspXtiGj8DkIxia59d
JOW8sbgQ9q5jL2k1g2rrexuKWcMWJQq0414pwEjpDSzISkA10osC2EZFPqp3xPnv
EMp+r7qYWbRCXRC9j+7H+bXbRso2bvImKleK/x4FMKe8q2otgyB7BwEHOunxfaYR
vxunzvd3AbL41lc9MiQ3XlHcuHwPXmbD4uBR7LGxmDutx7tkD4cUUSoYGfGPJ3QO
F1MlJNl5FeLP9WCQlbBGBXRsJs+iHhsrYy+t8N/JeSmS6D24JVhxUmHYi4LNh77P
1FKzxOD8fJqkvieJzztOsyqyoV49NFZTU53AZGImK2LYXhvaJl6pkAk0nfBaKIh5
x4hmGAOeu+tlpYB9+zunOxsuS/Sk4Q28M+9grNDgYKypB2eL1xZNYz/86DozohcR
v68XTduWGZriz9NQDpdOJix8K0RMWkcPYpK+3MzSA0F5YaWGRSAAj0c/pqaseZyg
Ej8TMd+bUj+U2OMVNTeHsLiuh6pS/jh99K7UVKWbNkfCTaRv8k3jJVdDyrV02oE2
iWu0IuAwc83DSocLKoPtWOG5sBUi8joMWXE6MeLo1PsxaFDQryQmu+FaARnB+BxZ
WnCPyPSM88zPBO4Rujma5dc4GP2AXXkA1V5gR7zFChrjRlYo03e6esM3gVI8eW3u
ylZbSdWBg4bqGrLJ6U1KKLAFoWnfYMmm8qB7YttU3/PpoiSMu8JgXPZSyQuwkXFT
6cWnuTbtBB9/Ax56aW3rjnZCWLr6JjCtq/tBzMAWbNkNOjVp0Tl0ipkzGPYJGtY7
rb4e4ZaUqYYZSklr1w4eH77/kYlj/W/GaWXtkzYNvzQXfAhAIvB7GMTNpwPnxHpo
38gK9FEmfTVVc5aN+zkQO8UcNpd6y/n7chS8JGZJnLgP4DtAcRsgh8JOOT/DGyim
xdNF4cLCtQPiZzEFGCtNPNQn1P9OPWgG+Y1OdaV1PVJwOX5Lba3ls/6bbUGp3cG8
fI4+nUptDp9yG+RCWvCPulnbheAsRkJXsEKmXT9X3op2HNmwwox50QF41ceWywBj
2zgYAuUaqYxbjsVG/1N5mVKG3bGuTJtvp8B9N6ZC8O4x32SLi+sgCxPCL/nxxID5
Z/3lE05o1fjatUzglbBmVEI9lyDjoSJoMofXm8B8bpDnDn2qOMxiXFqT/zf5mW++
SYhp5SdXF0+QA1m9jx6/lNw9n9sGHqMSqeL4JTfaFObdATZlSFlt10CXGMEBU/Aw
c2jsxjhoyp1dT0n5if09W5C1XI+XtzLboschUnmUW2Lh5LGkGlyVY1NKPkR1ijki
Xr5f8A1pE5zsCm07PL/qodgzil1jG2TmDsbFLvn7rPoItZ1PgcPC2IWuXnInaDwl
tii0ul7u0pIwr1CvN1yzoX50O5s1sxZjOcIWNTEny8AYs1SdStEkiTXkAUExVt/O
az9iPJ/wdRNEZSYhSilYTXqazO05/gbSa7ALlsXFxF2Y6rGMIv7AKdcirVBc99cK
VOPypG3EN9uyx5pf8DOjxkzTCLRNAlgGU2CuWhS0C3Zh2jBUmgKRmOzsrGvxnnyJ
mhnr8r+xEIEnvrBIVlSCM0Uz5YijlMp+L/vqJ6nYbG2vfmpgxbX709pUX/Nqtpwe
0gu9PDGe+fuNmeK9nmCKzOIEF80Wg8LYAebAxDS2PqXe0S1gxMu2aMaLTWJ2smmk
dv+uIlvVhLCHER5OifCM/lGwoXlsD0EPPNELs49SIGTOCZAIbk2DhUML/fay8f6X
4UfiBrZwHwK5XN+NV23R3ikngvblv72tM4T2dNrG54OWiTP4BAgz+jENDsK2m/1y
ocI8lf0ulNZITf+7FQlaRdtuL4xA8jtNw6CgkRga7aE4o0JRqo3vRO0n7wfhsYjj
70E8D5VHWLZUIEsrxdYK/w9M0TB06kPGCK2AHyXspT34vLnWs5ae1dWlip0vAMNO
ldCD0BTkGardvouTeiRW911cND+HaDIM3mo/H4gmUt83aQdct663zzRyAaKpOE4P
X5YwXsKxW5xeA8aAjnkilXppHyZYEO9ZqPOGid79L5ICmUT13EdZfluJTpZVlUGb
roO5ANt29HFj4KLSMSFDai3CIZpGWlHpwKmuvc5/jVOQm8N5egM3QF9DK64GtvWD
edTjF06dlvkxKQgEFKpO++kLLcPFza6S5jSvhm/xKIIuFLSxHxGXN3fGt8yJE36r
u0WxksVzBpSfVUkIKdmFuzkzLCUZOvyXWJNGKv9VS/Yd1Byn3yyWOj3eOG8+dDkD
l1A34bNfJ1vsLq3hToW3rpJqEHl/if0bl0jGqFcTssyhayBG64zPNi8kEdkIg+Nj
EVX4kE4pMqva2VXXLXJ+Rk9B8goJPiVWWXY3oWg37JY8Sm6zbCTnSlbplSIreTCk
7TpLLi6V0h1wk/Qi8vDL8GqCvTh4Vn35YiKJaO7hiLEYGrPxRJMPVld15dTF2lfn
KEhtiiKBBejhDmv2KKm5fToTZyOEt/ltoyIKJMh/iUXdMWq2NiPTrn6H4s9fBUyP
f9JiN0pq2cE385RAwmWEyoobIwMbtHdmY8Ej04SQDMpw1a4uWtSzcanhYkaQjy68
7uHeyzPEx2F61EHSSQvHzE2J7HndVkezJBYKNavCFb2bw1I8oUAt0m5sBTKkMtxg
s+bzDEWHAXmGf4QFfrn7LHv+EwNkytR+1H/0B4adA6jYLU/ttfD3NKsweg09uInI
8IUWI/fSpDJnWNS/VumSlqqAC31/vYVZkQwYEsAUkiiGPEtMkf74E0L3GAfpNyn4
5rzOiYCIKhLm5XWOrqQF39EIiZOaJmHc6kYQRDRtHgv057laRXqx3taC7HjGIMt/
xIdAXGleX2jN6vlSNqh87zNWQ4zYkjHYRHTNUtws6vPrA1QPm/VV+UhwTmolCiDr
Cm6aAK3fdUpMaPt06330a0Nns1dLSHCo+khKOVBAiq75FpKdA//1PmDIr6Osjz9O
9VRIFLO0zowrxTMDWgkmKr2RoXgeTzPky/5kujYtg5thsX0fblCKWMBXm3Gi9zVI
TbYlbk5DUTrj9qL6pu7hxXR9ENtMYY+//0EB4rDDPb89MB7x1t9W+EiOkS3zluv4
3xz/IdBuaViOjoMnLncRSKPIrgyWLYDKxL1t5TTHq6oFQ1AOJgbHtzILfKZ9a04a
H5uVjRPUVigTm51+tbc4MbEcYai3QcILqj3GPFkoi5hzcFRRDfdB9Hj3iqasoi4L
qj7iw3UoPdmoiZiVE4A33oifQ58xMXFtPotkImSuGnOfQhvUPF6pXKSL6/vO50de
K3yeJ7EWCn3UgbWmjy7eThQGEmrk3YRwu83PLd4EcfSH6taFXQCHpfaR1chbr0RM
88uUdhCE5jb5TXfRou6nrqvodOXUHTbwR/DnnNmPkp01og/SgjpnkfYs9OaVnzet
9hRojAMOxAuuLST5FdthGjgNDS02kTnkxpeT+fSGh//xGJG4vbef0WQsnXik6aIY
OZ2bQI8rjlxoTYmkMgowFmZXbn+tpfKwrk91OTIiDJhiE2847A+HM+uwQdZ0B/m6
GhGRPR6Ul+v0NVWFpO/sWyHQPb+VDYb68qfR+M/rddw8dB6WFgwtiVyCroqA2Svn
5mYm2xaFmLJQXcQLyIjQak7pYouYhfBwu6HL8WKTcwJAX5oucOISyf2uHpPk/UX2
MgQHPB7Lgg8Te13TLieuwIZtZvYVpQUENpp0QWZp95sjdS8iL5DegleeBcpvu/eW
1TvYkA0CJSgCceBYITYvpUlByn+64QeAftOVqNemh/1SqO5lxh3XNyi2DMgDP4ef
o6C08GlokiDJ4mJh3Ky6dgV0FIiX7q7yO99SGrnEAoA8JZq/HM1SeAXyq+cW7QDA
awg5+R/jIHtwUGYhPNXHXqYWRTYSFTGmeD5MET58zTbS5/qMJWmW+krlXi3YZanx
b+7mUOq9moLetSuhet4m1iptPmhcBT4o3ev0qhTbdk8K2RA8mIXD3ShIQSH7u3Gu
4VOgiNlpFIdRN5Qw1SYL/JO85i7XSv9dISw0AJ167FEaqbkaiTnotQm3eF43cqnN
VzTiMraDoUZLL1kcFhlGSAbotg13qCXNmvF83DKt40H5AUQFaSo5aquGTaYjqh3Z
S7wYvGtgC0FbmLY/n8VYmaR6YBez80OQZJQGQ+ZDYMuQpm2i3DWmJCs8gBSdWLZR
znW1xge/JrVHR1XmZfHGWcJo69Ic4aPgRE2TYerkFyIIbAJ/ArowWW+sI2unxjzA
aF/JkrgZxn0TxBH1tzldRajWhdhqLRhMPoPadtbJccZ9HP6/h2LjkwiqERW028l9
QZCwzV2U3+7Gr1ughHI6AUVsXvOMqEw2XMt+zEYporfHmIznDq27vW2BYouTmeT2
mN1ES/31d9Jaiivb1lzZAZG1wgVfd9mexGQbm/XLFPZls26TxLqagS1V9rOpmQJc
eW572NVizzzsR5X3/CU2Kb4dlukodjcOnmCOH3bwSxS7mLvdAvG7XDOFkGvIvTIz
1801Jl5x2HXYirAx61hpe0gb1r01zPIo7UzJ+pyRNjU7ldQ6EuswiTbgQNpWeo6l
eAqK0I5KgBSVjCNWf4LKennYD/shcEFT95Q7tH+dUn/Bn6HhxfZ80JXb5QxmkoqF
QvVeUKTWCn1lfgDacyxqg1c0W+bpYyd7x8K7oG0JZUfaNwSaBM5y/FtT5J/8xMS9
j2e6j+FVejb5i1bhe+vW2IVSVUqXp2AWThXxVQJ59I86zUG6vOJ2YBP8UIya1yzv
KKE+wTBp6X1N8jJEdbv7odUfW+RPql16CrvBuqR9c1orsI/ytS+vw0ecnAIa6C8i
QN5Ew5rynGg3yftTMbVxkDa15y0+LvkQA4iora1EenfvJsMU4x0RznWuEs5TLKQV
U7xzRsY3dZPvmD8Y7nr02h4Jb2JgATBIIF1jlOf/G2Eg1zS7jmh6Z4jCuhzCLvRr
NtLF25zAldmod7REbOQGIpVop5JzT68VJXfWQkdBJKIjOJRNUbYFWbS1duy2xchT
/5GLyM1QVIMxyaGpyIdaMsp6M8O5TUEzfles26RfvIybe0CeqmvueB+70EWO97ze
AwQgBG0uOwdOYxTJkkMEJQlbP3BhAw4KDFCqkz3lhybt1p2CNBFZlDTbU/klk7Ie
F9r4BOT94MALKMPbIj1YBS3UW12pji1GIS9Rg98QJReCrT+aA4jz4ADpRmtasR25
faEu0ejeGkTwWTw7kux1zadDYYnKBK8JlH0Rftl1oCHaXSo3joiXhxw3ldsZa6SU
4LUVbkwkX3AvzBGPi5SAjOvOcLsKiLuvqQ3ASeby40+loAC5RGON6MCYcESWCjOz
tVIYYKvkArox3UrIWXvLhn0j8OiK+GAVeMebYINjiiPv5rMYisf4g8YmcXvi4VFg
hNohsniG7K4DSZEGQHSXQCqvaN1I9LJRz3To3A2sxa3sMSR4CBzVEDTAgnkzEQY+
BXpufEnW9zYhBEcYSN64c2yDR5uTieUmYXSRi0tH9cjXgS5dwuD5rUpLoABoh/O9
5hD5yDYKk8o2c2oArTVHJGiWXubEgqtMMa5H67BZsIg6G0BcQHzGkX8PGuL+g8rH
+DfXstMnKEfDsoUVyipx/bpJEexqChI+jlqUHRuhEIdME17cVQ9irooZhoKyb6w/
ooDyOTi/MkxRSDAJQxUMDbitqkmV0X6RDo8ldU/rWpnEvmPLmjDqS7HBqo1GM22f
TLQhLCn4Jl+FmTQV+lyv5KWs1dC+vVvi00DGCElHVnIdhMYOFO5dM0ciz+uOUlbA
Ju7QfYiHXdYchPr4Wo7R0dLyo70iR38ABUE8fD/3T3D0y5FCAiFNpe4gOxtAfKgs
ls7e7dYu4fHGf/mCYiHhOCbN4HW4PgK+OMotEzrYclNyE9WZja0AyDQ0Br5/CMLu
Od6vum2+z0Z2VmU6cgsBpsLhkVFR0TzZLDPeNbQajhSemsCRQojZ7Cg4gYFeZ3r9
mNjmUrOkKwbq9TTw9CYajztgfFXlYC+y39FAYe21yQ8DXD/All6WxArjSfhg+Nei
ZzD5ggy1mx5QUBSI1IctD5/J0rUBWd/2cR3gQ7G8lWNZnRYUziJqUE459d6yzwkf
WNU8PEqpEScaf2fCNAl8g1txV1YCKII9A6G66wBVNfEtQ/nJH952ARadXEpXHKjF
UwELUWfsrD3eghvgMeN+o0QyZx3t230U7BYLIbGV9bP5Wc4STcZffG+as5L4/91y
5R1tvAgHEWPGFYcjw+THwjasktd/yLjEhJgcdw8QcroW673lfVcps1EPKXfTMwoB
baTCu4VfY+2Qqn/a3r2fnS+h8ID/W/9/FqrK0tsFwQuho4JxBDWh45DBIX59po1j
ISpSS5aMvLPzDYdNt9/CqoKJlaDR69Yu4cGRraZT40WbLZiZwipVnnGZbUf/hqdn
U6ZVEBhRd3txz9YkF+AIVRdbGct7UyWykmSTYTrj2NUOQ9MWOK4DhXL4mxFJLo7w
wL7+4UX0oR3wUKfv112fAH1dSUHFeXprsfjgls5Hw7rLLYRszvXGKQD+G1qIIGEL
Ubahg7id7UvmMn+fGLBwB8Ax83i9RfQ4FhmX41jLDU4lvyKkaLa5bDFcmcCFNaWz
WBTiVSvzrz96aSObmgUmQ/xrYywtX3ywx++Ks39CCmXa3FZ9FhS4fnnHOsLOVxeS
TZ6MZgoMZ0uhcByFFECVitOqgNIU/8O8DtiCMs5MgJGJiMZ7q/6XmhKuvqM9p2dx
1WF7Z5t/3aHzPo4zLB2qofENKiaLEh+itffA5YN/iOokfM5iExxWJvYmSpXwhe2G
wLfaLIK6DYExqLjV+/H653/lRPE3qttfAy4flbIdGffFwwRPaLXJwqaJFtbjKKVr
fLptljHosbyC0mcbool5gA/fLuBbGaD9pjeKNdwFyTP5TSZk7/avhwg9zIEmTQhL
dHvr6ZtXURdIMkWJ+Viy6Twi/jm04YgCJd0i+u4fQOXAWarrc/Xd0orgaTEat94T
nqB3JyVkAWpwvEHyubM8F+0aHMIFz1TDSGBBRRslZyJmX5y3NPKnXXBJsmOYSXSD
`protect END_PROTECTED
