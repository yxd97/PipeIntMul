`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIWIehKjV/MKZjU9uG+PONXh6feGN6WzKSPteOVfKHqDtZgR+yRSZ2/9mtKIQKgk
7ktGYuT9dzlArTB4yXfTDMtQ4ZI66zjIKdfN4kWEJq255F0juua4dxy0ePa7Y34r
revyrN4yPr7aBLGpr7MFlJgeymJJ6xkPCUYl6TSd60Q9DPnDL+No2smOdQcvULTp
Krx8OXaHkjZfJncVzkRbz+PH7tzRUu1ChmY9919m5HmF2WS6fTybWvSk/9+oca8l
YYrT0uURhIeEIW47xvYkXSRSvnUV22WqXd8tsB0sgs8kKjlnTSWSrzTqI6YlwXVU
i6d7QUdzGVLAoIBkur5u5g==
`protect END_PROTECTED
