`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ADIGnHpq3jZ/uOLAenMemvYgG61lzzkNsLBo9Gj/VfclGA1sV14CvJxdzYpeoqAz
NmFU26q0Ow5fG45XjBV7YfngeYhe1ytERKIyji/KVsYyl/4JPqm6HGLupfBhqY7X
COeIAr4ObHMsfX/dL61ywXE7/a1ZSty3Q12P/BFZr3Ck/i7jtqCiQ0bGHNlXKUWR
v2aW0MaDShQkD/IPWn3+agEJoyZvXm+ogheBvUrPAEIVQ3vpUc7Y+PSLZRAfV9UO
ZMXnyEs/Zu3yUDmrxbFcFh0Kt8i26xcT9RuWTim7+LjZ7cyH8X5/M/pXezJcepYm
boUB3Xo1TDNM2BdjYbfTh1S3B2SXZui+tbKBFGMX+at3OBVkWvfywDMWhdPW01Dd
Mfywe9HzVF/ojjQsldN9zSLw7OdoFGWwBOvbemT8t470lG4PcEYDRrLn96/VT+sy
/aWc6WEENrBeMxuzuRto3nwILF+8qRUqU7W17JwvX/o=
`protect END_PROTECTED
