`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9I1bqTH0lhK2eJqUlZv0A8jn7/8S5UVRjS49gceF1hK+LdJ8gISVhSnCkqHk6UvE
AY60usN7rkcXGAjkNSCvg/1XvPwohEmh7ycI8yQCFU+/ot8N98rPUrCqoqfj3yD+
Ab4twwJZ63fvIE5fL6u2VQ5Y04fRQg6unhhRzHCft5G0ipRvrIj7NFyZ+qn98Fi8
DDWh44Y08yQr+oXI66oWK9GwX7v0YrMFGRS0Qo1ohPItJw0hd5Vxv430ggV+KRfW
wERH0xJGmtNaUvjSCdaL2S7YkEMV1Iks3TpnJi/aF6CXoPLzsaRodEYVMqdvNPRO
1o1Cayv4FBsznvpSxPJR3xgHiwKMZwryrDbxu6tXiUsRs9U+9Kx1tt/PKMR2NXTK
eJaCkCOtAbPebWMJfGl7hSuQa6cHq90AvaALOXRr4Nc99iYDfTU+yu1RZReyREzl
H1cJyPN+v+yuG3aOkVbHx6nYP1s0IctZzcIrVW9+JUzrEgMl6rl8u3LIbIaT9IP6
0vf/3jwhRvG9JY//4ZlxFtRsJsr2Rv3oJ+NYDkwG4XJC98CK+GoWPexayJumrMHM
C1zX9sM0wN3RdF5kaKaWryjTfX+18hYHo7U44rKh2NO+uXa83EiLPMzRGQfpGdJz
p4hiYRsbbUzRCXQP6kl3WQ==
`protect END_PROTECTED
