`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jjt+UVwD0t+zaw0EkHn1RgtenqrNF5yZquN1Zdk+USaBftI+o4ykvpDhvxbGozrP
EX4Xk1lF0WR5yptRAoFjUc0CDCfVytzHWt2v9voaP2sxEgRl9/4HeLv9QRXdsDqj
cczPP3TmFNdIssdBMkSw52f/csoUm8Vu1wA62WO+Rv6Rx8AzklWG4Z48dntMEs0V
Z3FUv4yQ4jEK598FIeexKMfSx7pwuyD7GEYPTy5JDsBDBn75oGWi8yixFCEIAyF+
Y0cjywR4idR17fAEmZD/470OE8/2I2VJLM1CM3tu6lkFhPZjCJELrzZDXRn/AW6T
qlsO/xo/XjOTCcZP3rn8juZblUhhzUjPt3crjSyW3lUYPaVKLoga08HB7czaOGCj
01Io9FuOrnV6xShZVBRoIJ8R/pf3fAsbCNSI5HvObOZAM3QenZnFgfrMuUByUraN
0SgFhroGo0lGYiUKDscW4hbMQvdAh4hmLOptpJQPxv9TfwMRJsGKz9rFhnb7rxTm
siMu4IhvJeXFEqHdVynpwKFA4J2K9l07cqEt4+Q4nWvbwTyplzdDfUHaDPnukd2z
jL98lNWW4vGpRuQR5t1modLbkEfGEnadsLizmZsZ9lP31kakWpXgzQOliaOLqTei
NupyUq14KZpkUWKuwCHPhWuBfk1mXYRvh4pkACm/s2ILn6N+JOkcppotO/RHTjZN
mAxkkGx4cA3oanaM14HG424Uvkwbu3N+UciBbnAK4Bzw0qVdzu582tpfq78KelM7
Ohwb8TIWZwLCQl3+h9VKncT4NOPpAwvRcSI4Cwt6lZ+Bczm+CxS9xikvQhVQwSls
mex2Uu4rPksI0sUjAHoBf+DcTzNFdwtkv16s9PVQmHW9U4drETo6Y/LMiN/BS/3Q
`protect END_PROTECTED
