`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLHPFXbVm90r8BABqIubRju1xeobcb/H6RdMmdMibMC4UBX+2n8F2XQ/xZAmBO7Z
vYttmf9CcB34SU8XstIMk0z3dPKb9bGc9VG2fFzm6sjg0j62cpNAmOJsPl4RSvI+
Y6uuurA60x4Te2LhrX6KtZX5tJbMM66FJOG9d9L7QViyRPDtBcC9WtQfSI3SqhJy
LKU1QREdj47DqeO9MCJunv6zToOdyePnF+7P52SR0f+yf7hO211DwZNcXWv2rngA
mNzWN627QhvLgbwLqsT/h5qzoWJScyqyShdprSxvySZyQpm2+MCU2aUwZV6DYltL
O/XBAcUXs2yNYipLWvWAH+F692zKlaczbDpXrGrE49AIJgiyZaNG4CC5nyesoiqr
jhRU98GgUJBkGQ2lQ8aGF+BIG7KnwiG2F4BXiYYwOHg4H2Gfj1XeDXau4tgnRnm5
uBu9PGSBLW3b1Ui5+H5zRZZjofg8aLHxUKzIVpnS3gK7p9uSZTOKhXzFDPWDNWYn
N9VCBmDwM+r9SvUWKkoFpyfHyKC8KfspKX7YkKJYfFfRPKYX1abttVdNC2kvSGCJ
v9GdfbTzTh6X0Y18Arln1n2KzCeYwSVw6nKR3iBTERk=
`protect END_PROTECTED
