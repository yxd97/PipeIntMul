`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bm+7CFo9Nc4/K2nupplpvnx6FbSv5dyMRiJDbbviXgbvDv+8efpakECv+PY8bUXP
Gt99oejgbYiVazTYKUrfpmmJYJemgvf2O9oxnZchs9gA63Wk2DS6FrbCuikpJ+zj
Fs4loWJ/Xwqopm9s/Wm7aXx7JIf2bsjYih6xhUgz0UT6XUmqSrmq+2PdI4YY35yO
iXmCDktCNMnwFIAnha8Ek4RrvGG9oSqHvDU4Ejhmg8P3OVCcyYCckIjzvqNRACrZ
HLggjJ/D/BmgRSDX1osRdUv+YifydRWjvU7wkQjr9M1SS9OL+HoK5nEQ02MQmsMQ
mTPOxxbX2a1iCDWk818OBYikFTt7zLzyKk/+KcsvqJh3fw747+BK/H9zsh2n59Sd
lcPyRfWiFZ4WX7qk5gaMr5Q1i45BihWbv394a4hVbf7PpnF0ZyNGP801A8Jzy/Iq
dkP67bnilM61LffgPaROdC0FW2EmKsvJ8D/cSLzZP9+oNX9lKHVkvM5HbnC1138w
0v5elj402u3maywP7aRfvvFFAajNuh4OUbvpn0ExPhVR52XrR038hXjbYzLfaEfz
BTi6jkcpaLSWsQuJFPyltnbQtboqHzJaMKevLklFrnz0S5HezFUwurza2qCF8q9p
0W+GsnuGY68xLgn6ckY43OYEYo43dp1PQ9tcKvUsGcqyAZFEFeqJAUEV785ObDKu
T/RBIcY3MYrZyCbJVyxHJi36/8JFeC1KdJMQvI3TQcQ=
`protect END_PROTECTED
