`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YYRDpxsNspNhSYXetkeT5mXbDhCrbGJQwhQzeQ4Cwddfm7QpzTwUoz8t+xOnSXFS
g/4+I2OFzQNAwPftSxa+c56rNKlzg6fO0c1Fz++ko+jhx1Lb5pJpe5M/zN7IaC2G
0jZaaLXAo4sxG+eGK0x8r2c+ItrL03Xd6OQ/Xp/TTdmnRP/fV/4FrXtr+D08Gswm
LMgEHt34ufvEUCWePCiacswBZ74wjpn5+92xA74uvsfvn9x6JtgCWiVdTnrBJiHX
c2rJHSdB9lhCsUswYUFFoipeyunXT6JQShBITxbbuAerifiraCrpM3zWqQCaEzkc
eBd4sEUS8e3SISvQ59fwbphTmidQpw8/BxANY2RGO221FO0pIZEKlS+I01NXp7G7
IeWH4PMrmCfrlnEWXGFV0FzKiwtoVHz2b+pAT3mUeoISaZ+5eHOW60M8YuGK+u/v
wGfDILIZk4iN45fVEXIdMqAZPI2Xp9pRwzG4xoUvUc7IQKFM8DhRP3H7zkIQG9Ip
29p1JKCk1mO7vQOxZrSD9lQkybmx1xXO6GDwrXvJ2hZJgKLcNT6nrOtYulAtzAyQ
wVIQPWcP5wO2j4KoDinlBjjoWEgJ6j5dsOqPIiyPfn96ijlTr2JQcF6snWgna830
KQLEvXncnYugmL86Da7qgTPhveJVHFcLX4a5ZVZNp11DP9jIFWrsNHsG1/M0i890
nOZrWHFCprS8JszfS5lzLH4GQBuF61lM7TCbCKACMCt+WbJctn44RRep09MsRi8O
pinRj6YuUymx20HBk988RS8EjYr9GUc+lmMQnLFyL2ap+4auY31g23ktOdhwqDaX
FtRU4ZxNGIa3u7GygiInkEdfx/p4Mo8Fm59gn+xBDyw=
`protect END_PROTECTED
