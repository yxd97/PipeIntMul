`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2akPYAX5VIHiLxa58guDvT/G78/JaMX7l2DI2rhgwzOWroAmjx1a6m++hjKhcyXh
7RMPAvJQ/4LhNOVWah+hAUpMNSGodB/KLLvw8y/74jLIE4Ed7YGpsUJuO/f0Sz6x
3So09WlSltRSIMuT4AjncqkuQJcXsNqTcizZvaPCCfDw6+ebAzvlPXR1XNHSGNtB
xQFaveZE0zjKTytrrTXueNTzuOSNL9bCgf0PFmKHICzNK9AmuBYUvudTumttpY3J
RFDi/D19068FG72Sp+1Aixvso/nswELwYOwJcNIoZ+WQicqM50SV7Pp0RUptcxh6
wjRApl9JtUqEx1pVLhRkcQ==
`protect END_PROTECTED
