`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuqxEcE40qa0VinvFM/Z5AKN6ta+Cch4j0eRwfQY/lvvodQQvVwRCX6UP4TgeBKp
Lx9T2dGv4unCKXxPDOD28iUsfGv0LLNhBDiwUOchY3C7DTa4scSLBZ+maHqjW5bG
1w5xb3fzJENsKKtEWL9r+c4JtHDWprxMiZ77okBk4P2zWYtf8sL0iviCbIR3mQeI
0ga31D/V2VqPvJFiVNCg3xt1JJ2J5z17Ow4dhI42odAF7ip0/2et5jiyZkbNeRS3
CooYXkDAwLgDq2ZjVXGIp2QemDVBKW5BYAQYxiDGTu4Ihchp+Z2rcRd+bGwz7jaw
/BNV0uKGCpalIb/rMoTcNyWdtGK/W5d6YnXRO5faK8sbrBHEZ2ct7hXS3yRA8Hzd
AdSI9WtzvOd7mQKX8LHSCikpZ+EkFulAQH8BvxenyTX3+BE0i1rHJocEsg+Zmq4+
dlN7fThpuNo/uKcErbD4y40trOseP4k/NmQowuepCsRrwhvf7a/HSvWjkNDjQCqq
FNwHKlnEahIRXVKTyDhWHkqxQwM+pInGr57bK/qx5Iv9MVEWJC4vaq+JqaINsmw2
S6dEsJ5qC4aTccxs7tKFDsIPLoRsfclkSxi/wz5H+re1fWvMnNVfusLDtaQQYtsN
WqDEP4OAtaTyD0R29wThm+f6pZtLyR0O0anDgtz2iGq7bTxPi2EG16ID7oX7G5R3
E7lBSOlAyWPaykYVLBoOSULxEkdILrhq6MMZhFGpCLGFFFRiYi7GcSKl6P+zQ/Vf
1V7btVLA6QSqOH3em0uZbUHmUxCT9ew8rFPiwy2kuBqQ6pKm8sr0VGaAqumHTJUf
G9Gaaid8z2+UFqSpBluFAdYVTcn1ZymPIaoq2rSkoPaBhQELtqrrE9gbYNH93sQy
VVMiVrxPFp65lXMmdmtJnLQXRFQ5izU6onGjXdyLH6VD5wzc4BXh9F2kzeFpFOxP
DMSOaIM7V6TuNxbQ2X0g1ka1Kka0DSuCMIvL/nGxKVuR1yBioKjB/GyeuldoRWf4
VMvaH4pzVfZ3WRA7mi0SK37O40L8OFgqHT8hQurHNl4bBElqRytPJdYgMi8u/nTw
iVUkx94f2fjLlqJa63lrGj9E2VtzB6SASJnvCgV7SNR7/dh9/sXZeLSQevi4zHxp
Rg7JRp9awMu6HwKBHdsEq8U7xhOYdMa9leengp9Tos7vH9OhA+qFRZ7WCaPLuAdz
9K/hubIRRfVEHIvb3q7BarcmxsnG2y8QHB2pJa5UKwFsYabH2qbrUPFz5Lk/J4RG
GcIxVKirrP1XefVvizJ1qm/X7i2wiZHpXKNaJP+yAo2INPnZFxpRSkr7ZY6illDf
QIFcnJvPWvUf0wBS5TIARS0CpwLY/H63ADRqOLEKOQ3FEkjPUuJG9p1LMp8gEiFT
fT6Q9y0xBg2yfJ5AaoNdzvHZnrQzqwz98RiQMFo4MBJ6e+Xnowi6USMCwcKioDQK
8mZxDDrpk6Q9Eia9s6RMO2bSmgA971NMpKDgXa0cp5W99R43LXDDwjPCBhMmssXx
V9jPHP+Og8TcoR1k9Szln8/AO1iC8A9rDzZ6QbC2W5OGZI9O6RVjT9LWdi5laZDM
Ma96dVh9YJ+tqSLYdIS8qDMq2rSdZ/8dG0zgfyELwAf0cnyxdUrauey6jijs/t8N
+V27QkDpmNPPjloSjebpsxcAFXk/LFpZErhBTmIqriZchNPoTnB1H0bPnjHEeLMC
mWdIdDuiZoxTS5zkJAneYMrnS1PnllKJQyOE2KndgvmwzUuXtBJI5IDeE/neG5mn
0uw3JFfWgKkbRZLH4jmAkP9J48JvhIg0Use4HCSHd8T5mWxOlUJPVUh6m4F54zLk
bh5I8gGzvCwGcKLzpMD4fFKasDEGDBDZ6EGk8PQ2PInNDgp+mSfCHL6AF7sW5ewn
F4+N6sjfy2ZZmJkGtHa/DftzlsetqWck5lOQygLU5oWgyxBrQxXzK25vYyJ0ggZw
FsQq1ZXKXZFd6NcAVsT8A5ofGeC350/KgiCqcm2hUdY75nw4c6soqfLfV3ddreww
3nhUvBDTRdnZ+RP7JSswLU/0v018Ux0DVsTRdUF0ztQEYlc9c+ctFGL/inT0PuA1
5emZCM7J3Emm8SfGFwO6sIrogephkBpX4UVRoTE/aPks3d23rV0x/LWq+rAdVHul
r6PMOCop3vXnc8NIesSjRsRYeQmcsWCz9IVegWjJAGzhVtYHua1a0Y6DhHHCpgGi
ngyi1VmXmn1f7svgNUyyCToEbPnNFYv46HBcezjwd8oQ14L8fZwsvnRZgLRe9NDL
7mWoybicG7/7WWWsXf09xJWuQdecOPoJhtWYcC/RfyrtCXWF9Gq3G1D5pQqlev54
VDB61sOTbrgqxaUqkTpSmFTKSNg6Q0ZCeW3qeouE4bv51CHUiO0K4hDiM2aq1qws
n6BPa0G7MwnIKxk56RDL1D3QIw+O5iBHlTm5NC9u8XRLfR7BMipzAjyeLVKHpZAI
6u00jgF+0OesZFiSP94fNFc7qWsCLcfIh0aKHCn1i9tb8UbqDPXLtd5t6rrc3ToU
/8nW2ETxEO5A47V7pghfacltj0UMZuN57P6ijA/P7VZnw92PsYc3m9KSWjHdCwwb
C0sL6mufV+te6gh7VFELqnhRyU4s50aq1wtx01Ha0tkU3jHJnQdcOZFb/sq1JD8E
x9jWaU3/8b2S3sS9ipbsUgjEwoW5RHDKbGG+8/dXgi/+rTK6+Nj4BnJK5cMWzaDy
g4i0WqzqlwflI1k9BIz51JWyVxgiuz+pkscT3fFRH9rvQtUX1Seoi793vSMioB7A
jH41ikDP3bGwibRs7VxJR/QF0U9WVBBWjSuTBYXSNsc4WxYT1mNm/g9kWk0jg5Ij
g90emyKfrYOHo0an6NdmvC9zSClOsid3WG3YhjEsmmPWGeiba9WrizJXaCC1dTO0
ciB2mmk5puBQbq/gEAeeBbHxENnZTAWXyO8sf+udQjjy7+TghUWt+pFn/D6g4Mv8
a7EpahrTcu64W0WEvxoaaTci9DFc+WMcupSbE0OtWZMewW8FDLItU+94mwAPGwHJ
2iQfi9fSkcu9w0RHPkT/67Nu0+WvkdQzTXKisGVmHFakgMqBPgbSfIyVRzEOaJIU
5i+2soP2p1VbVfv6MjvqitSj/P7OncTF6ZjVMbp1zd9jIP+nIwhtwBZZYzwHZzdr
EkI6IDT1DMLkrNFjgnSHbLUz5+0dhM6XfF9zL2RatQcbokHzkrb4tkoIv5nRz4Md
V5Clzu6cGcMcIwBI8gt3GCcAF7HMq5YPSE5q3yoSriy7+giERlUICwHhaxGYpKp9
rgUD4ECaU/UFEeYXPfxsOgCfHbwKSJcDFcDEWthKApauSRnx8jQTtU/mg2g5lYgS
UJGseBA76/12y40ibJ8L4ywmEz0Ks9pu+apFjdEc9ZklHSqh8waLkmosA6HwDjA3
Kgrf1q4sqeo2L6IwMF+G2ohwax+rqDTulkdo/dwHl0Iv6AUC1Tynv9Rzp17xt8of
VX4wnOvMxfR8KU/8iw9b/KsuFTXIUX3ox67UqGZPKncvaRp32jWS32KpEeZn2gKq
gPt4tY9yQcThc1hrowICxcWJUh72Gf5lhxtWuobto39CPRxeSevbGKzH4Yqun7TM
qVAnIElwVgVRhOCcQlGaljCq1BnIPMqW2qXSnGBeR7mYlq/sC4tmb0WtwSVrQrMC
f6hInodO1O2N6a3Or57XmI2sBv9DA/1pJEtOjvJmx00SRZy16u4rlC8Zo0r09f6A
wkBbcm+Ru/P4SmKTU8MeoYS3hhefy6HpFQ9rRnDZHsK+hIuZvUseKnKRpON+Ox3U
o0gUBU8/L6U4g5wsaqWMKHottN9IFrJwod1yMoj/a7FT7wyOZw04oFEDdSG7dM5y
AM9ZxWViMDqHH8mfu3UMaUaR+qp0CxnMCTfF2DFJcFXGZOh9hB99r3EXKljQNVgU
wy6rwabDelignG3XwVWdEnjC6Gbn1NG/mq6caaILZ5tlmdb1W6FBCBBZvI9ok82H
8+GfbfnDcwHBHKkcnc1w1RW/29fpN2+ZdJoYpk3eyyh95ikgUljgYsLkp5MRSeCQ
ZPGiru37o9kjZyF9f1qELyQqBK7LMLRPVEDDt1p5kENkFoOMLnD36vyb4uDbKpM+
Q/Pl9DSCCc/Pnhhj1ZSjzBJD0OL0V1hZF975xwgP/dXAjlTqttHkXgVVhizPkxl/
8GvT9yw1M0mhlby8ZLTns2+4amn01vqYK8H3mONdKV4STIsYB7jPZO3Z7XA/fZHo
RKDciYAkjHMRvpO+6RiiLbgvAtcc1Q+1nIMehoiaUmsnfJfuk04NXNXbEtD7POYZ
ApzNddQ+51bURkStN4NGc5attTFGKkUNvccrgIbsSFNHaWi+gKSto2ye686oVMj2
EgRfknxyCib8KC3UyKPyoVTMaZjoitRxYRPOaLyc4Ztco7TkhmKIlbLDV+stFgbF
XyThbOnn+WL/VLSiK+hZRMpiTKqwvWTcJ0EmO8mx0fpsudinHuKUm+wlu/0Sw+3Q
dDAvAypG+iWB1JaAdHafn17PyXzcQ82DWNp0yOadv9qr3KHLzH+K7HPqxJdGlko9
cqt2VRXawk30OtHf0FYRKcQQlL8vPYXfvth49S3vXIzcqr5ZhgF2G7EF4x3ZEIVL
+2Dd/7xFC/0xv+U+QxSl332oqiBPTvEdgMCYO2yRP4YHn+0z9IUBS970FEBQkf3r
k4zPmi7q4xFOdqQ9e3eYVep/jMpPZO8teWLWMIzqiDJzxZ6N1fBlsdI3ngecJYhl
gX9h7h3zoyXHrpoqbNbnTAiMIp8D+6PbTMKGzMQ0Uj8t7PvloNHiyarTFRAJoaEn
x/ZuD2Yfp3SMFWC8qE/H/Huvye0gHEdKcdA8YI8ma1aVlafC/nOFNeJV/4+TRW70
CWHBzxAn33WFCRISxBLaG29+AEs6W9ImfG7wxXcvs3f0mZIrKsUoLRp9ONWEIeEL
uaJIbvBgx9uq8MSn/Qigi0FHCETD4GyEAr81XzrrTvA3gVvD21oeIaW0ojdPT5H8
O36lDMn7qCrYqp2srvBN9JvUhFAUGbk6bqzBKKIs9cvpuT7MtuCWdk6exTsat4yI
Z8k3MVeU49TmviqOvtpnd6KqC47QbFBMJ7eOUOtVXiyZqnWYZyPB0HoQM4HGCeaE
E6WjlnWuf7Hg36+ihMlZ+yFQkY1ugvo+IwetrKQEH6GpU0zSw5L3/v+wXpzF/PNA
lPS7llKMlWJUI9LJMvrlW6zxSTv1KVyGgAyRW2YcYTag2ks6KL314Q9Qzxtd0xWT
1k71ee98mCeptJlX1UghFsRQE05r9+r1UYTZ2+FV0Dwy3HJKy4abLptfpzgMuCgu
E/tbWbXzmQ9AFaCcNHzvvYERuOPj79OfzFOL78IJnKxMKYD0EPlzyNS9EZ117Ck5
3axTN/5a4aVXty6qm/4mhvXTXM7GMnha7nZ4EiHTYpB4GU9KoBhgtjeZrNvGjyEQ
zxSA7rw9GaT3WFrp1e8YhD57C/9laAQo/F6Id2ICEBpFtiqUDbISh/Q4NKRR7ilZ
hWJAD9fz0/2QgrTF9rEtGn/W/yHUoot3FqKXBpd05xMOs2/QtDkK08U3B5gMumaK
Tf0GeBYNE6zjxB5I3qlo4jAmAyadUJ1yFGvYP9V8mkvvS6uG1YrxHJEaNIv1iJnL
`protect END_PROTECTED
