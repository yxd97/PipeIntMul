`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpewnVG4w00xvWJpTc0pNFlRQpdxdgxz6FqoNtCDnwa2Kjd8lCXhW1Qedo1zdUlN
jpprhnqhPE6czYC2US+ycSOs6VX/ynZDHaNoLSCNheZ6mWsy5FmIi1S5tezE0vVa
W+OTeQNDDBptxPqR5bJD/WoN0j5ESp0hlGCkEGZV9Hlp5CMEGxEre3NZT7CNzLvW
dAJ4V19a2jG7y9sGWGnx01VmSbXqxmFzwIH1HlZ5MIx845L6ogFNAWvMMPYxJf4T
2dK42twsfpotCX88Qrfa1bMewPIGLlxVBcdUGwRRTYJ6x2m6jG91lhkS7QJRpqnN
t55AJlJcqFb0LeVILnYZJeOin8sP0KR+A8MRx77Tnxp2+kM6a+K7baJXCMte9tqB
gk3pwYQ00g3/e46RaTT0UJX49ZScX4UoEaaA5pcVV0GFNH3z+8bdIEk55/eh0np2
nKUToNjyHChnHYDQyE5loFLLlcE27Qac5Wba5urui+61Kw2cpik9fh1sdT/E+3Kj
JY+xVGaZhz/r42FN3T1pUi9bKPbEgoaN5tlarEMJvxs=
`protect END_PROTECTED
