`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFQyFQ2YwVjjtCgxCzFmy7s5uVfe6lPu1HGKnDDroY5vQUXb9DSX41zfBStZg5To
Xvs4ht5GDrvhfS4umATFNC32mXNqukUVZkTzOA50VhHRPy7eBj7RDfv8QeLq5Vri
caCjhqK6YQ/0HyekhNlM5edCWteED+VOB0qD5mm9X3i8a4S2BF0ly+FqUWmMWuSU
+CZ52MtSg6SeieNudeucWU2xNvoQr7QdOrcvdd9M3QsKUgQN69kOJVV8MUMQ72aS
fR3Sn9KkC5XJqSxlmUosjrE0BC9S+fS9O8sbLQs/vh6l7GWeiwF0l+zE1ckd01ae
K30W44HeQlUXS268jbKEubmvSDfoh0hJWMpqs5bT0PiGYdesWZEx/bC5fu/1qyfh
FM8zO2HBUJPBJbcW0nCg+SW4WAoNdD2NDwsWxKg0HkWkFIAWvHROdM4MUV01NJJt
wmS43+QA+iBUEwdVTwzRb3XkDTdnLw+TV3CXNR6R2tB+isXBokPy/pH6KaiXA1sR
l+8MJe5scziD20kFjykCtwrHx6DFNJ0BibZidehaHvz/1XzLVLVp+ANt2aRTkjOk
I7PGMYSH0Kvr4o9B/gI117CAYWkH7W3r/Mv86YD8EA6YwnAhur3yL8IDkk82sQFt
WSMi28OaroOx5N7idTEKAVSsfV8cO/fGEj4/Fcf+vs+NBlcDL466mLpbETlG4NPB
IJNy8Zphsukczy1leN0uaGWFI5etY9Svs5rd+8pu/ihLiTn3buTuStYousqQtK49
7Wz/57qc6TzrvTlt9p9uqjkez3+oRNNUqpKz51W6sgB3fjxJp2cg6/9ct7D2M29M
B9aZzVSvkLb02Ocw/Wy3/xU4BJbnb4utbhL8D6Hq4GfqbcVj/pGMyzVQeVPbEsek
6FiE6BfRuJ8aV9YB2AVdbIBYFEU7OENzlELaLTQ6BZJJ7Rb8Rk0583zi8FxtOzvW
`protect END_PROTECTED
