`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
APpUMC3wDYxTmNbeFi02Q9zrMbWPINpxHJmGTT/gPNCFgRBanMwlMPe1Q25MfiV8
xsg/0iszMMKDWm34L5mhZ4lBS9hTXZs17OONm7vQynXoYlEiUnNngkGj1DY2vPU7
GSJ+aJHChBigx5e6P4vRwEqsMCgSr0tD/Sa3PDMc4UHDF71pO6oy5B+R03Qh9aqB
Uz88+Wbn+dPFuyqvJtfyANOlTKSE8kedJe86gJXUmc7RSUFTIiWJdYVjTR1ELDp5
jM2SMg/QoGjuPQ0sPcVHn8X36uYN7gN964+CQibf/XbpdY2w6XjrDYDzEgdPBY1f
ARH1rK8EnoyusxccQeIKZYadouR8+hTSzm42qenlAxqSw9UwJhv7DVgoxG2eqAO8
`protect END_PROTECTED
