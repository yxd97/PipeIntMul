`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4usmz9ijUIb24Lmz37g5zxW+qIahNL+vezW9GpbdabliHYLjvBnLw1SWTIRWL96
KBOcIz4mW1gtAFUhWvwfGtmS3HpcvBVWGX80vRba3CbbN+coVsfrGnG1PIB3W8sF
k+WyNBJYgFrFobDHhB2JLshEeaT+r3k7kUf+iJtdV9znxcRWIuSHvRpJbfJSa2nx
FZ3ZaEwb9FLZpzQ4k/16/KgoXs5SLf/z56TyS7MwfPXxq0jiPthPOawrh8z9bjdK
xjfHG/HSSKUUUiJ0Os1EotUeKLKEKeRW2fv9uWEH+0PyanxjT6cE/wjhgZZibbC+
ccUcJ+WbGD5suqZEnmkSFeMSFgPYWA2aF+xQHlnLsDTt8mfECriPJEA8FB+NuUAz
6lI7hq+3vL5C6jgmWB5EvWeDOJ3HabxpRsfZTAsFU6ypGnHAjnPesko9smDOC85A
QU7cfAJKSBPtqAU0/FGEAzhY/e8pcl6jdli/vVY8ua/K3ZtAduG4bQII79zl/7uv
w8m0UwSv5idsOGLD3E017o6NMNhWdzHyzbLv9NxGF+3dylJb6EzdDlg4qsT9rEjF
qYxBgaKlUnrKCq8jEEc9rg==
`protect END_PROTECTED
