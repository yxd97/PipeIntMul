`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFeXkHk70S/XTrCPCYAGnyW4Y5eK95iVdN0vG2SaCAK/55GifzGfJM8dNGvYMA2R
jBtZULv+ZtTmfIJwKmHutyekq59dN4MKkzftJ4NqAIVmwAzrz5kRhjyJ6OiFZg3k
5EAcdw4+hwy+BvfR8XEVvO3TA/OX/6WH7G8hLB22eIZq0h8DDdI4jhH4EGF2aSdY
IZkMiOxko73YMe0Qp15rNXf7AJWdfc8Cck8uwmQ3s+YyZlrvs/SEZfkKKI72EO3n
0TJpIkn1RmXIY7pbgzLeBQuqbTJ7vfoW7IS3RRr5Q+0nDKqLoFmgAVG419NOxL0V
PNpvEuURziMLtLYOQdCNWtUJDcLPUJ4TOQwltaPPYlGL1DwPzYC3qKy+R5fbj2wn
qnXxCTwd4lcgOdsmHWSMD1bSNPtzaOt7n+RAAN+of4Yut2jZZN+/WsAA8AHF52sl
gaIJOUlvNTExj71x09BPhtcuUTyTFug4+rycqhJva98SiUqHv1JlZaBlREkpw5vJ
MTzDFFiKpbBrlAGt9vz1bsjcTIpfQs1mC8U5EC7E+VVxSXMLOqaIN5kT5SrZXyCV
9Drh3Liqj1+83HhR25HMBxBRlEH5bxQ40BTTPKoqjMdXoEMDNmAJ53t7w//CpY7G
6NBg0ey/kZeTjfiGC4L19myo0A9BCw2qNtzzc3wBDcd8p1/YKAOjq3nsldZ/L882
l92ty4ewgXDw0CeVSEv76hP80oqPBL1OTqsxOJ7kuA+A2/esbwXA1GwLP45Gx6eC
IMn6p+RgXZeZ1CmbMvHo64+78NsQfLGkYjrjW/POKret782u7vs+bjFaz3IWbdrB
i2JLAUUtAnj5TX41kCDZxuzSo3wOxAz5z6iFfKaOXkM0w4hjEk4vX1CZeiHsCi5Y
kNCIv720mDFA+zTnwon2YWZUjai0j/OeDuo0Iw40v/Pku0V2QQ7G6o0qhtvzE/Iy
Ma2WmxQh2a56OTK5ri483ObD1BmyektMIgxPFb5LE1EQ5qPM2T5YVsDMPVmekRSn
xi2Ic8qY9gfturCBmtJYkBJj1tJI63VeQ9FofFrP5Uc4hofXQLBN5mGM90azSobg
4kb2hA451SejUd4/ck/TaKAXaRkqWkd8EqSDbodm0MF8idJoYCQ+FtesA3UIC8ng
Qu6CLLk4vGz2GbNNPeKsGmg9i3x9osIPfiqGTOxxEIU0pPp2eSApY+RxyRjf2MBV
5A2ndO8xhMdD3jgLzQg5ge3moZPSdrTmnMHlkPSeD1qauWdKh4AaFYwql/kmZJcy
CGQQszrnkhw4PJgoP/v+tSW/XkPVRRLZtIbLUvstfErZ+Zge1EA3r9uaTpcsskb5
ASaCmPXM7He4tEKf3gAGx1Xr+gWfIk31RkR0dwKuGnisUJ1GcqatMyYhHWpBqS8O
R6d9WDg3oUy41A3hsmxKh5QEbX5dGG5yQJ1DWZNiW471sNmCIlrnRZqnmRog+qyy
ulLXk4J1eHgOJEKyzVqpsdqC4gWNi2IR7gPSScjrwTvpDC/Mf2JKzu7P72objeMn
92Ti89GI67HMJ33tvLlGxBO8QFZejhjZR+Xr/M7NdL1b7AiLzyBEzHVyOIVINUpV
RkCCNgafFIXY/gr8v8DtzEMRfzzRWfCRtZWcG/3tWXm7nid6fFhEzQgs27nVPVcp
j5bCvVeG2S1ztMueCMYMNTUxww+ld7dNgILY+GZE3eeIrOtuydIvav48eR/FyiSf
SX6N0SYntdLYqLUrPvh3rw==
`protect END_PROTECTED
