`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPFGCJh/2Sp/8xKGNWRQdesWSPEBHrGlEf49jaoHI/7dda8jU1g11PSfYwiClmOc
MALSR24Szb1Mq/6u3UhYA50PkJBn95r1mtR+o9Ihyjh2YkHSSiQyooi//C4Jp+Bs
f/Qq3F5EwqEzaNxz/Ds6456/Nx6oSP9V7EdXCBpbc1ST8UuPLOZa6TlSPtxMDtNz
4T/Q0KXDqXgqrz9ObFDL2VmQjSwKgPx/VWIhPbK6Nwji1vem8VjFpvLxeocRxGNH
Q0goPANArHq9uSKSpZ/tG+ZSaX8BWjCQySxvhpP8AC3FiBFWoybTIl4eGkjOwVcF
1Z9pJ5SwYJ4U6GHYg+D52A+jpwUznG3Ynh2zUj5d0McVoT4QEbittpFkfDoWOgWP
SM74NFp9aNFxm+YTn1PZZK2AETOuromxhgZa8CURzHc=
`protect END_PROTECTED
