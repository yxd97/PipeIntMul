`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IqUQkMgdcH5cXZf4PX/19dst1HCsTKy3TeFYivgi1maHEhVYY0ffiJ+U1YfjgCRA
FUKmojsMi2p+RhbKXtpJ17/SfqLvUv26MTWjcbwqoEdadNwCanqRjxilYnGS6OPB
pgoH2LJwBG779/eXJtPJcTup2PsLx9PeWfuBl1sewWOyE1siSdS016lGNOZpPJnK
zkHvj5I6DMhrdbMHKUuY+dFJK6pPHUHrSrZVusWfm1RpEbrLW+cXQn2WCzg1ZENO
iul6srOlfKH+ImZbDImfjp1aiO8rYsVkDwNwRtPRV9gQt2sSnH556VxxPIY6Z5jS
WJUsEsm39odUg8fmzwvxfOTN2pPklPXAKi3jL12ibQAtmFwYpaMv5qzxDtJjhbtc
1nE6A/KDQVSV4qcjXu2o9Wohz/ZnX5xowaFtTB8s3y99oxolx4mz+Y5eaaCka7Dc
yApispFmSEkY/kaQZO3R4++stvQ6wqecglcRw/eV29qcXWkqcYSvfMlbIV+qza16
tUsqGKgtb2HyEaBVIQRV59z74QDNVBbZAIdYxGUyqnA0tkC1to/ZO88RHCk9YaKE
98m+PZnrN3A9fmhHrd0uoiPIB9LlsP6UgfQSp6b1KyF20oBg0mnlUf7ceDM7hGVN
Ggjl6jnGOUMvX9F+fXxXDUrYGru7CZsKd2kwM8Uk95Dx/yEldEtkWVgIT2mlQchR
mc/Ss4olxrpZn3xd2H5Jfzn9WDj14AGKAN9bGmltD1NPEa1dRSXc/vIMTBkqOemt
sQHScL7otYs8GDiygGTNr3GYEOfYmfDmKS6yvnN0ce4/aNG5EW+msSVMsHkhJoib
wv0EnDrvcLYArvyyMFekPXP7uDwdNiFzxf2RvA3I45sgAERteiS/7Tb1KhJgLSAM
EGtZdwRgk2GxutOK4A5zreIbPbiXjTXUC7r7V/xHW7RPpu7ow3r4nXGZak3lRAYR
`protect END_PROTECTED
