`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jnGzd/2w0gLq+jYAR3avwluQpN5HPG7GvzCIiFTH+GGRm/Rg9rp36nvcorVVvim
AdJO1QS4WTlBdWCiQWF2am75fuGbHyrFVreGGhC1ujmk/MIIOEDt6lK7ssNiJO6V
qKuBVdXzUcSPNATsPxfddEwAiqgkLUo1MThZDHlIca6KbLeIZsplPfvpTBeBMj4r
CK4kXnYEAQfTaPmq29cZ4yQaK3ZvUoPOQGKXiJeFR+fr7RGbgfCwNoj4Z2Z8VBW/
DameizkgUuwxjcv6pLz3DPiRBtnOJwkJry9zo1bSkrlZ8opM3sY8lor+k6tLe1aQ
2O1N3cfqJ8b6uE88IrurhpE3PI7p4gNBznUvOs94h3NgnKMFwMi9tUFlLi8B3cIO
hqNSqVaAbq2VlvY2G4nlDiVfT100PEKiQ+k4jIuQq+OFshdayy6cqfmC2b+lmBTM
+iStwv9SslX/qwvS+5K1qX5BciMj3vicTiJoIUmOhcPFxOGSSgQ2sm7NXA9n0yez
BOiFIUcNbMK2QND5xoZ+AX9hCUJu0eb1W5OlVCXENKKyUdcK1u52CubbsP3c5Bcl
inf3kJK+oa0OFdjwb1Kt3blWkFdn+4n5ysdIO09NnhcQhCy+oKsczLKr9AT6ocCh
Ba0IEyhLjsOAdHxMqVHdRD3Mr4zKhskGTqbpR9nTZyTu6X3pydyD5mjPrxhGVMk9
99QB9sUvgLbezbahbpw6zEZvZR/dbncl7ptzUfTX31/0S7BVWwpgwBXQEWk6Cl0n
YwAfDn8x8xW924cOxLjcXOEGP8JLjl3PdDMMaJqw/MC2GfyC0owKIT21RwyA6X+Q
F5WJwKEACw/DTndxZAHKoamzcvZAIQsDX4exZqjkrpNKOZoBpPv7T83Kis7MdNe5
FYKFrRJOt/ni4YTU85Iae3TQaJ3sW84tWGL7bHyj3L5rkr0LNkN8L/mMTJgcXppl
S4xwqCjQDjajzxuZoFsz3q6bseEDHblPEOkqR8d/iFUGnXdsGZ6qCwF24CBmASqJ
zwTSJs+FnSbTO86ODI90xTIn4/F1LzK979zv/eid4lDOf+Hlu5z+bqOfWXp4f8JQ
X9WqYeCe2ymB0l+ID12rpg==
`protect END_PROTECTED
