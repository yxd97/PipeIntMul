`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GMgqr+WNF+m32Sf8waGX9wLFpUuNc6nqJ3QsodkVNaUEDDQFXZosW3WB1YAXzLOM
QLzBIQvRpIxw5nnEXFWFzl7mAT12zACCwtLJZQQ56zEfxr5miMe1ntvLw02Z0erZ
AnuSn5MOl2/EEmB2Fp5D+BrpLU1hsR9Nto0o0mQ6mrzB0pVV2j1Hf/IOfxeS3IaP
o+krGxCGqztYxa1FS59skjDGOqiHjaKHMuvaY52+X8lqRy+0MxXMII5Xif+AZ69j
wfsXS29K2MKnw6xA9nUCaQ3n5KXE2uKn+GFnRbPaAfyi386JrUe0przfevC+TcXh
jmRwyCUhW6I9a6kIkTlOsCBlyW35tafa2fBtY0v6n9cCpClQpKo+tH/jWwiX4ht0
WRQpSMdrhTfQNLmJrIvH/noagkRXJA9WllsaBwjsEJt8YsLsj46Ramt1vCZVxVxR
xVpqsHApW9bEiCKbT6r61QDgVrE1H0B4yKUm6k5hRDWY/BWzxm80ftWm6RoVNjRV
`protect END_PROTECTED
