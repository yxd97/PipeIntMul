`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5SohXafT29JWyxrpj0oYotpI0U+pARzOC2DuuPHY0dGTTk1UTgr5sjcTwfDLkfx
ecVfOYhx2Qf3KRtXVjBA5D9UE94/4tS48Jmkh4yPssU+bm3bakReRBFfAQfohMQg
4Rz1R9fozM/YvXiaX7E3ZYEN7B9ePHVAG+t0qLVY4/zGS0C6a87eiWAcHXI6PhGu
+FH6xwOXXJ4eisuzc6rLigcAkK6sgPhDKOZ/rpanlGvZJP2kapGy8qtSu8cpzqRh
oi7CjV1eJeNnDT1vRhmjiwzvXrOGq2GepYj0cfMBnSBdjB4c8aKVSFSmKPqAO5jm
rkpgE4b7pgA6p2j85+BH4LcGSfTXzDwSxdhhwlIYvKtna59B9tLE+n7s0BOWrlwU
`protect END_PROTECTED
