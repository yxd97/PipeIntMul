`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+FiSy3ddJftrhPJ8YSxk9uQDBl575cvqmRKJmp/zVNXgWBCKXEXMVJKdUBZ+lwQq
AnnzobdPz6otPcD7FHuiDeJsDmEXtvdtCYQIEgU4sizlqn3XJj1fNEKN10OX+VoK
g8k5LBrCOjnkURvMNTIAdS7XcFVwOHuWVCeeIlht9kWdQsM6ka9jfaJ7Rb8JyD4+
zI3yu+xTm9wfhAlOBf+T/9JOsXmbrQQkXTACoFQn71v49A+gsl1VCg3LCxgx6d0X
Vjksv2dpjZWJCQwWDZmpHNFbkFz1YHCfv5dpJeE1LP2kWt+5tBgYGMbmDGsCPMoR
tAuqmbchoO4nTscTwVi6iQWAw+qybTP+aJFsftu83xUjrNIZGG9rnz4byhVi6+ZE
kfBE1J0kg5G56P3g/bJNoBMu6xNJRcP7qd9LjFimAlI1Bo+drr3VMh65Z3ONo740
1B5tCSXfGMFV58ywbu49flBDeMZ18kSNTtcsXEH8sQuKpxW/Ukm0oLu25OnUwDTg
A66JTxlX/S1+DfNqEenYhO6rJZ05Hx94SW8bzGEyO2Wl5WxHEUY8UuLXCHCdWHwR
6Xq8dBJBykmHCvvnIO4sCrfxQXjFe/Q+2oafzPqkbm8aFExR/QUlEzJfA6CmSo+P
FmV3UEZCK9fZjZzUQnJ2WzYGk1WtLNADzth/LfXZlcEyQtbzrHCoC0W9s/8QE5LK
nOpQj/eh4X+IDHZvOPwXEaPTPmbqkhmajPZBpn9MfR+NfZFvmfyXuEeTzW1mHVvz
ClhDoVAZeOZobBqTJHG6hP00T0zEGb26vBCkGsWwge3PtDjst7qpm/6FVXuH3Dw+
zi7nbCjHPrmGj0jdGHhXEYJWAQhUvc577PTcK9lDUdgayw6JxrMKFmiMqfMrw1L2
Xb35u1NcG0UEPk0zJ9kNuJX3I+/eGBFBu3a29aNsp+wZT89LeB4EgprQ60sUASZL
RHFBL3T5Dn/2C39tFqU7BbOGPt7DuUp9EuJ9CQiFJzQrL1jHNX0MxikWQUuSf7+Q
pmT+RDyypOw/UWNeJbbZNu79dHkaI6+wz7eM0yNNnqv4YDrehWU369zT5cbuoNjT
RoDMKoEdF5yU8HS0F/G/QCwIArC2JKki9rn8wJIPHF2SPX1o0oxLtVaxkDeq737M
oYushUGJ0vaEgGL55s6Oonm9881D/IPxQrucN8Ief/oy370jQFkwBC6yeqXnpyv8
sc7b56mH8RW0p0lp1mni9MoEN6BYkUZfvtNLyvYr0C4MBr+iVkiyQwUx/vCZXwuo
LdQsBuYuX3jj+NnL3yenb4cIWgkDEwx2Ih6UdxnfW44ocD0muY+0txv3kdF2da8J
PtCvuzyHxBF7CoLm2DPemrVvkoobuv7urVIpE5O2j9fRcbLHBt5R4uB36T70buWZ
PW5yV1vMNzS4x/SXpnTdMPztlS9vDDMl+r1/XyMbGAWLlCwDj0aeFlx4wAEUo0pB
HfOc3m9HdYbUeWG5pGv+sZvJHSRe3DkIf+8SC42r1IKfQyVxA9/6JnGWR9Il9i8U
lc3i6ibKEc57Luz9YCD5/X5AARifrEKpsw+gdpZemu2H7nE3uAfnB4zSM5/ePyLm
fQvagRrZf5AWwdmewWGWH6BuLwJhb/vAeK2gEc9Kj5e9/Cd8lZKxI29Mh/gKTmaI
eHF/TsP5brsGk/CoadBAYgo53KNuIfpmt1/ZiLV9BRqsmSxIzZjptrK1x0JEuVza
6g0eTyqrY/ZriVNTPjOWB2LjwrM2hhmcGy9442kmkcy8LppnDW8bwDhfSTqzXPv5
HYn9B+w41sCg1BIHM4FbCu/8oBaCDlql8ts8MViQRJhzHM6/HaF0agP4ajC58nuq
Gy+FHDydKkqb5/fn3LVMPKLzGadWH9AzLbKLn1rtbrrIKfluaDzgMVfbelRc8EtA
VYGRuZGNJ0YZXG3NOVE7+ZiThZeu2zcI0d/p1eXvwP5XmX9djQMXyTGIUUgRFFTF
/NgsLzCTcGwDil+upOheTcabdVRXWr9VqPR5wgfDX3MPQfdQhGe4xzNFcsVv3IFi
XnsM1HpI9NL0IWO54lbIDztJMZwqif/T0entHQxSjXbLbgIwJhgksF8IWnHv/b1p
EzjuAqPupf5baUJn0G0nJ2uQQf+PI/gCMJA4zP5a7uVCtCqEFnVrPyTLY+xjBJr2
8u8NCdwi0fwEipPrDqO/PGLSPYjeRdXomaK8fjxi1lK5l18uYNSxF09ynO9FTRlH
1XRKOYe5ilKXsR8CGb9MBUEMTVdHWKgCwZBJoW93hAmwkPIqSyadRvSBGD6oaiGQ
zh63HwcZ58vFzxxLVPQdRdHBOkC84vBmAwYG/reHBMcN6wBiGV07nlhi0HUStc9V
KkQxSpcHUwMN3Ts6K3uINIzK+cOHhGNFOfdv5ybAIGC69lpwh6PAv/Ao1Y1flZdD
Q0vHkS3KPskwz0R8i+a+l3U3LTFaJlu6bkGibRYMiRehlgvhrMSez8mF5k5Jmf2n
ZmxN+khyUaDP2Fw1rTJ6yfQrWFl27Tc5nsNZOPx8AOUWvcPONRZQHSZFbermdcCg
qvtmgqT7rsUWdNhYtxi2m0uMYvntHmdzpuGtVHaBqwjnyzF/xBBePUM88a6TBpZC
zDj/fnOb4/izXPO3POstj4oT2PauAc5cDins6Jcj479o42k3/fssODwq4QXD0VM0
QIDzA08mgQxFTbXOr7dSf4E7mKkzDXdgYKWLXglBHIvuXwW8YOWk0pm77GzXwMcn
NQNuXwxdHkSiGxd2y+sCbZFOHrexRh8c7LDKTGt4vkRUF5JTNm50Gkz5jmQyi2AB
P6yJLdQ/OLqMSN3a53Fwpq+ajFgPIAKKamJi0uTsi4f6RHWP35OzdMQZEMk3PqFX
PvtymjpICaYrG/7RchWuPMJ26c4KiQL6usaHqal+58BTHsZ0DwIzAW4XlPzESXHN
ltVJwENlkyA/fRXQ50F2Yu7LnbjpJTl99gHPUR1ig6Jh/pbheESDXSjuLSWLWSyH
RIzh01sOkcnPybBWimMQF1Hz6uoMOxhuTuACo0RsV7swuebKq70aAiVYQDn2rkna
vwTxNKdlBhnoXsRSY5kSnE70LSLAwy1E+SrMd7t4n5TbXNMnL+LWBZCAE52zFlN+
0uazXv9tpEji/Kyg6mBjGdewd3zmzR4cQgs3MrLEtJ7VFESQpB/cqF1H0hTolWWz
PurM14Es0cMHHQkH0tT6MopNo+KtLZaFgR96F6kdwoA+58hbMnDeP4aybyE7Hvs0
e0wEEQWvRTJjsM0yUsi5rQj2uxHrt1rbcTivS7y28ABWWKBKfmO+8XxDgatZJOsk
LZLoLwFHTp1LEfHaqh40ZEAmZv8iTL0afdaDoStsMJ8N3htpeQet01ss5yqm/Y6i
FHll9cf5Mh1RNcTDl3EePGSBeJkPcSsW1G5smk7BfupNNvPQE9qpmdpATzI/3wCh
WWOLvZ7Z/H+t614H0QLvyWKRu6RsGvGQMKQafNbyaROBgZfERlO2txKKGTWQkd0K
qXDpTCheAs9Yv182MqcjQT+hPA/aYZte89eRZnQQEk1jXLQsSgDVfmMSS5oZchZU
`protect END_PROTECTED
