`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ulkyPwJjUNLfgls6Ygj136Vqy6aKE06P1+5RF7KfpdWK8YUFn0ahFYrhEStqorr
jeZE32QfYVCnrIt5drvhKkaILZNqCOkRH+vJ5qa4DgLjSCSuplDZnD2Hd6PjzhjC
dz46p8QBCEZ1G57CGW9BxZpbaD0VjBmsvyWsGlAMc9uFTmgLqQuA9cheSEAwG02J
7w+0Z8qkOdQcA2/43TB73gnzva/juZ6CBuYmq4OUOZD6eTTOLmMkTMeSo4CxcwpX
jotiSC0jzUwivm1lS1spANCiN7KNQUhIWJ3Oiu7YY1s4CGt1wo1R633ea+XzgFrt
x7blkMO2/P9CmzWwx6DrMjPVN1DXTaKHx1+FH4R7DscxUpX4RiZ8ZzfFeS+ZDKHM
8dYvMo+OXJZVWmcqUPiT9qQ44GQ2UVQd0B2QoGdE8xPq8+dNesK0IBzROO0dnNe5
JRT3cTSpQLYWKpqspfUXglj8NBHM8OxpLlET25pxW0WSTZNxj5EzliO9DqGHQ2sZ
diq9fRztnGXzamgNYeE4EEaeNLhM4TxuugTLKmzfuk9SMaO3vSD7yORt427Cq8dX
lJA+IVk5SXDcWPXoYRbrqUda6vQHqE3GxIYHzpsQpeVhZA+qfZHLtIqbrGUJ/hus
CsZKsdH0228Y/eeUQ3r8/1bibAe/khTgvNppV3EETvtUtmzioRZI9/ejlJx33D9M
/33j3Z4CsWstgkGCIk5RitwfQT6cYwn6QiMyIfuf91kvDE/K69y2NPAxRXgOscgF
h2Zzv7iJE7Ni5EN4t//d+CKfInMfEkL1MaeCgMN8xhMW9M9ejmvENMZIj3pB35Wp
MPdkFlTmEqg6KlDdBFr5K2Fx/Er6FlzyZHjpgPA8A+cDVwK/PUq+vV+lnK4h8I+0
wxUhL62dKv9xFa9IBzMdGg==
`protect END_PROTECTED
