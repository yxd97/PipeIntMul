`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6K7zP8IyHZhNZR7UaBg4xujvYc26YVnXI/9QIv30PxVEXxoaRCa8yyTlV9Sf0IK
/xBk8S/GQq3hSUBwGYj3qWKnZy+9YYoD9avnrkWdcp0yvIsmjZfg5eNy73rpkdwU
4Gx5Dp9+aDpUz0qIwc9yZ9emcXbQKHalRr1RFOl5vJzB5ZIWHvUso2rWyHWi+E4y
qteZnfPC6kS5/G/vYo7hx/cycNLejnyEskQsOR3hYZP03WV5R81gSn9+orYE2tmu
NHau6vWagKb59NI/qd17a1lNB5O2gwkzCEmhx21I7GvzARW/FtSRdm/QD4RJGHz2
ez4YljkVH0FML9hj2nKRdH8Kh3KG8sbZ3LPgoHv2ekC8nyfuVXjRSDbD9fd2kASR
2khSViGtNK+GQsjARCGDGbG8O/SKoM39N05yPWQxLloeNlTuxmyMnbVuXMOzY1co
bCeeOyPz8FdlodMyeW/nXnYuKDCDlGD29etdZQUuZkg=
`protect END_PROTECTED
