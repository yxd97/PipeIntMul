`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kCXCsVYwbPiiwqxksWt/Wrb2xAwTju3Mo1x4/6oMJcX/xAlSlaasIow4CjQaCD6t
v/Kmp+WnSEHRf375ieNqv/+DbYjvpmWrhMUJwTrJZ41O2mypQkQoU+gy+Q5lWHp9
lgzc+Oz6NgUbaSGwdrHjp2/KnsH9AzKpJzEo5XE2lLx4KNLuOlYyUB1uoY+c38F+
32S6ibbfPu4VQZBFu0naX+GpT+Mp3JgiXKRwmd5Cqr3A2E2YPPBQmycOujmWww52
rzrECMgot2xeW8U3kWp2viLoCkmnbluDr+abRJhWddwmen5oEk+B8kHZmChzuQyg
b9CHsKZoZROTX4bKUpEWpXs6K6BgZmAOBUfboSuqcwTINV1oG2xiL2PlItxZ0nDs
/HY/Dk6OE5qlGF9xUVHOPoKW7qrj7FttE8poV6kQ3i+dGeI2luIP5OSx47jMuwse
vaQlOFXoJiWIvaqAxrxqOzEpH1DYIYBKo6EiiaHAGh9BgMFZEzvdai14XAt3lLVv
`protect END_PROTECTED
