`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
krjmGlnGxPF+zj57mBxPRh8v35qDbMSu/CcM/83g/lWaMNEZQSZh5/Gv/1wlKTKI
sxBs4+NWE18TQtSUIqGah93hsaGgQDKGRfbn20GAJqP/Q7eBMYagQJVl6x4W3THu
oLxAgNo3wahtMjdcU1f899Z8yvTFjkGOzzi7PspyN+5oCsckSr25TnqiV782eeYb
QIUPIxvjqkLDCq9E4Me6Yp7vvkYahEUujFAPRHBg5yojMFfX11ip1hIXvnBSumxQ
h5b9w+Ju5mjNeKvDS597gJqdzacc8miWBq+kJhfdO85I8MjXsJeCH9ON07PvSCJW
q5qPlj6nyb88BFAx4+t/dD3ZylEKBSPqETGAiRe3claAatPU55dVef2KMRsl+kUy
YG5W+oZsGvPcLx4hR83OrfWbahDUTSy2Tze6E7viSBeNoxmbP3P2EJUyprAUp+AJ
VIUdinpPe7LncMPBeIjYle2lnWYFlhRPu8crY+a+HX4o1z8EfDzVQc+22/PyorGs
8HkCH1thFScm+Pix/zP6pGNAUNxzwyp/IqnEdmbxaUog0MgbFq+DBqLyyWfW2EAf
+tbkv7GoouCatAb7QXYmP/ImpJfitPZ9lOeC+Gjcw9iu2sxqigu4BOT6TKtJ/yNx
7s7TFBMqCraRY2fGCwp+P1s0HC7uLVpGsXTBShvksK1AOcRtVPlUufwCmuJj49Qx
NK0e+bw72XYPcphtitM2n2R0L+HUS8e8VwEuY6a3nwHUG1qs8IgC44WB1dr+E8xJ
pAOGMqi8ck772y4dwMe801npC4z6C/dInvlDf73gWauLbmWamf2mGyzjWKClnU+W
JSl0xcNbG6PsXfw0XNUYQ4MO7b4sralqX2TRvODtoTOB3A9GCeLbr3HJQOIuozFv
bO3puT5ZK/ehElTb8PNrZYKXV6q04UE29C41PgcuCrM=
`protect END_PROTECTED
