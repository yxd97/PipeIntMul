`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yzYXNkJgxsvgQCKjlghImgJobPfGTcDLQX4/SLAkC5IW+cREbSwGyX4XhYI/hf0L
mLsGYEU/VfWuncljNG6GSOGDgGklQ6moB4Msnts/bhKFCbIcf6iT6/l1YmS1kGRN
dvpYw8bYvJHZ1+ipVg/5yM2FX38MrHbCGeOUXukXNIcPDTFODze6uBUYWp2O76Z1
VsOjMeTdO62yz4+xxq4zRcUVkiboY4coHrcSPH/LysQ3QiPeOtSxEDa5QvkhC1/p
dSTI3WOM3h0uKecScDpWkSiC1Pjy2Fbm4ugztBX4Nju8vkwBWzz6eM/pSTR1404h
UcQtsuyhGm2QrYLmYM6LKEYd4+nU9JbkHMaorJCwjVrnWUFzj1Zd6Ozs0rzZnftn
0izpFpmPvVs9sc0i+CzAe47eNk8Lk5f5yqzKGndKnRhhkGhglkHXqHa3StQe8+TU
gOZKNSDTQD9iUIfe7v47w1+2EghfJRTJiaN6OyRPmvayaUgRsa3FiNpBz2XDq0Ui
g3AvNJRIB0C9l1ZYEGclu0jO1RHk4+c0OCOuq6uYVXFqEhkrYIhtV2JqYf+CKQ6h
pNVT9SA7wzlnbII3IJ+LHxpLp0aqg0LrkN/QJgbsy1PilWPZeoKZV5Z/S9TzTvVx
WuJ2zIiw56UPLcsQYcwi+lZYsNKgQW0EQzjf99UrU4BXNO4Dttp2a1qleLi5mYQk
+KlQCXKkX3FUg0DKrBI7tLncym2CTeeP/6TDc4TPPhGnkKpOgmkJuahhi4en2FOR
0H06OOW6mA7HCWX+mmolKMF7H5MMFYZTO3lkYZkLSKvnGQDrKPEvzPj9ZqQa4xfE
Vfmi0I+6N3MViuMOhJqiosO8qN1sQsTPcI9h5LMpjGZwUzoXbLGkcgGdZki9eSPc
/hYSOvwg+DMTDiC3mog/7ZidMr5nxXFvjZWADKGVk7mSmqRM2UCCJ5DkQGLfkrEy
H5D5TMbyYC/wBv5g8eVYp2ub8vZ/++za/LDSQUtU2UEDl4dAczoI8TAWCVBs7QKg
55oOOIQKRX63NyZpQFY/27nHDF22tFKaJ3Fc6b1fc5JJOWzzxKj+9KOYBWqLbUX5
FfuOGvr6axD1COBtBwMOEY1EoVvbFp8GqMJQdo34/9Tc3UffiwjTmXacKw8vrP/0
+9vIDh5CR/cQobvC9i7et6OyRo2aLeGGH+UkW46ZQdHA7o6gn1CVZxk5mafOfcxE
5P4dAWwWv71qTlDkz2w7fVW32eZ6AWZCjGjl+0Hvx8VBKmgEiRvRkLnCRs29BbeR
`protect END_PROTECTED
