`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAdpYDnqW7r7S2ezM5PF/JBVyXLx/3QHxVhcvIQaJc6/3miEfrssU5XEPdw4P4TL
VQ/bslZoqsRJfni5UAFuUtojI35T/mVpGL+Mi4I+QIK0babGkfiu7C3dOo9lgaNw
bul6jqxJtx/NIyYLUFjQe7rd2+r9+dLjKo3wv6I2JGwEsrJFaxtpHu4/t1YQYGc7
gCSkgfNffzrp3xbkA6bx6Z/ZLXgg0xRb5+d0VFsMhO06VTATE7X8oVcyTUZQv5+U
L9oYtqjuxKoQIqD1zRwbMVJwcPHrV+sSPTyDL1VjTcu4DzQSZEgqXE6S1hsU18Q3
yZVtbigcPvuPA/WDTUI/RBUGiIX+Nph4mpJezxPHIFan2BTLATzARvo0pk9hbjUb
`protect END_PROTECTED
