`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VwF1mZnwY3K6n/P3+X4OLPhse7W6usfhRmq7vVJwosz58gdkEWeeifNX4ixrIga6
/aWILgqOFWh21NRiE+wzKyefMG6Wwo5nYMQPY3MMGhE2uGBUwofMvX6KNb5hWtYI
bie1gOA6fd4+bHvtY1R7r59IS/xPBPIh1z1X8H1YJUc1tpqTQZ4ACh8JHYCTtLjK
2RhKBMs1AZeu7GJ2nOY5p9lVfl74ONaldF35etz+uaLbyf/UxzxJHfCwfkvmTa8+
gKPXv1pmY02RwaGeiUNgPE2+IfPa3CYpaZ/2EfehfGSzJojrVmVFX0BHi8qMekf7
zg5u7pqrkhVqPRT8akPH9AIlhSsIYfocnrByrAXtBSu9w41CyMlsQwMA88cxwcvp
BIuav+qYNTcHnFmqt5rQBg==
`protect END_PROTECTED
