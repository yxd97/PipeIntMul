`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+xv5tesQ3cVgnuFFeOwUzHB3+58jUKUUCNGLKifcee8L4Ugzy2CM4PIFIDmyiAt
1pQ36aZESnZRovl9yYkOYEjZoRlc5mAc+q1SCXu8+uCPUNGoGBHT/qPtKN9dJZ26
uoWoTO3yyIEaIx4/AnuHWBprrralppr8Wi8LIoDrolA1trF9SPBBMPsMnC+SrMIv
ghD3LTn+zK8I3TwjC5uWnT8/kicv4EPF2x1rCS79hGuFZ//McXbGdQqhfTogM5ym
ATuYDd7fBMPjn3MfEBvXOPquKUzNy0SBnViPrhgHbXTBQWv/KLwH0qSx2Yoe3dOr
P/3mviEry2ztA9CS+qvLMf58CfyexBg58aE3ufn4KOoPxkUaMiuJVTIY0CoLOkPf
t6+QXQmFCuXQBO6NjDEyTJpOPjTtA9nSb06Ycz2HciPHoyaNtq/MMwpsa2VYVyrI
uQSkF2JEvp+1Be3azvgWo1Gwwy0CW/pqN20yU93e56MQmugxFCXWRELSzE2Nersn
0v5s2GqGophfBtfupb8Z8gjiFMwwC+IUyl+C+Rn2i6BXlOuRLGbSuTlHhvD1UbBT
IerodSU9a8SRrj8iI2FzJaakMARCi6+1T+K89bIyYsMlfrmAhpnD7RRB65hoZyMv
lohTZrR+v0K1xrwpbcevdZhxa+TxLkRiNGb482A113unpRJnKdqvCQLyW/nTebrE
Rm9ikLknGpujGV8WKBXdeSNd8k3haspiakCKwnkCbv3bMuDcuPi4cR7O31W/qTW3
h+laH31+htN39Ld94zC4bGUR0MWgrI5za9nGo994qyv5UMIdUYIs73VWbleqnpeM
ZLb98CBwmlzCW2UahIWCwntgIC9EUUiV1mBfmA7WSeEXZnXFdYlh8ed6DdhP38Ug
n4Tvjq+jPMZ5xJtSaNOcFiVn3lLKMIyH+M7HS/gzsSJ+TdEAwE7PYdO5X9Y3EP+X
gzGlSNl0D4kwpJuzYDbfeY5u9AWsCZ+Z8A4x2HUqijEH6jn/x9Itv8Bi/EgMMO1n
`protect END_PROTECTED
