`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gq8Ity2K9KRJBNCy9OZtrVlvfCoG/fiBApagVe9+j189aYJR2I6PlWvbixzvrDo
X8eJS2pJdGFZTDVRFYaBZ7HV3LVJlzcSkFYR+cyOOuPyXtycaEkZhW5AeqwhLt1E
M5khbn4BaxU+8323m1MRGVxNCw9A87q9wAzfboOWCd7DoSEpPlR4yksLLYuHp2xn
Lf14t6wwXzoxjUhTcO+A0Y4H3YN6Lc14iwgjtqMfMtQDCOufkcmYtnlr5a2/rQk3
5Pv2TJtl+KnKeOj5W39hwbkZZz55Dxy3Dxro3eiZrgDOCEaSxjxMlWyVH4evbpQi
47ZG3wvX77mMzbPsQsKL5R8PV1PI+64x4xS8BOkr627bPUFb26Ge5Buu3n2E4Mr1
O+dCUaRUTdA7IpYOuHNUxQ==
`protect END_PROTECTED
