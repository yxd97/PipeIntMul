`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBu9ymkNV/UeMpmcqWeulyG0mPOu6IQuSRSADili6X3IAr4upudif2FTGOIR4942
xOmDEwpqoNvya9LlqTz8PyN4OSOp63mMkz1ZGmkMq0jd2LZklC6rOZBJn7WhL3wP
TYHKFuFGFrbXHdhD5NqwhpjIezixIp9KLGGQE2Gju/GWSx3CMsMKINQge8MciRTm
vofr7VF7210Rv5cvDg4EWx5rRB+rUOotmxkg/OQLdPN8YjD71rs9JMCgCwiVzNZv
z0liWFJ//ZVK+Q3ibyvf/WyPmNFsIojRUdQv0QstJm3XOUecfBNZ6yBRc47nf+4i
Vh8B+v5EeY1SzPaLuP9jlpsX17agXM9nkB2wCCIC9+J4Bv3nXqM8xQN2H9XT5CKC
Eu851bPf4bmNcZ76AIH2gXMp9mbxFOV04VAIPOLCYk9G+cMCeOb5oTHLg0qvFaFT
xsKZ8aqacEA4hdqZ4UCFvAUNEg8ObefQIU+y+w43EAs=
`protect END_PROTECTED
