`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3V2yYx/ZLLVFVRXe8UdtXdDJN1xkmcRZZ+eL48xnKg6gTISYKeucerO9QaFuU3XB
Y1FmHK/ePrkmuQeTpGdeO6vgsEKE1I6p8c2mbxZuuX+uduC/fOTlLxKQeOgnNBvd
JAaiqNGFn8fmD2eYppzxnj26EGQM+xZF6hOUXEvX/fQQQeW97scOlom6rN3aWCG3
p4Afk6yu/fT0BgvMBluXw3EoygHcGpIU7RfAmqznFRCDBN6Rc9uiqSdKc8Mp0pBb
0LBbr1SEhWL1WQtNBoKTSjnvPZY305XVVHOWJxECWSlsWDHzh/2c2PJFQF/NL9Ju
H0s0kIO8SQM4r7eHzf9aog==
`protect END_PROTECTED
