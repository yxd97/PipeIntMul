`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
45oqLKTIyK7iAbb9PUqieMFD40RjlWTmGc4l+4HlPXKiWOu2Ge/6yxFetxQHvCgm
uMmJfBUQw4U1lD4//0J9OT+lrOTL7WhCoICeeYDMDoIKu7GWW0dEnxdhi98/nb3s
2wkS3qNkm4tYbV/+TppkjfTeGIn7w8nP6M7eeNRVSZr3i0P6dbZF6abQ+xr1X60m
x/F8IQzEKf2wkIWW5jHAUobvPN2dDLjIP8QyOUfaQNkEc0+2tw9EyKlBgeDj/iu2
y4IU65CaZu3H5WiTeAefyCYO47MavuHWpZ5d4phn7XBY+RkfsjsbBMCdzymw5+kA
hOA0mopgCFDIOKdO+bZZ/OOsnJKt7WHbtPFSBscsbtBer4aJMoHvF6oalk6KS0jc
Yhy1M7zNTgDWKrqSSff8d6+4wZOq5CFbVhlaJZa64Qo=
`protect END_PROTECTED
