`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rfiai0531T3xZG5e/Ce9H/iEHqcb/5JPtoE+NtqQYU9YPB2iQVWK3yMKJPwObXGF
D8Jm/gx7Kc/rGFLjLNXv2i7RnRqfVWBJOdEzmuC1ZabwVwU09CbACAOr2NlIPfdl
i7MnKKDMR8xGQ6ggxaU4InQt7ueE2F9n61tebkuGXJq9vIS9CBczNnpwU6Lhf09G
qsC5n6hnx8BtjabT/TjhH1r/zPEBx+B14Vm10oCrLpc2fosQ64gtrm/gOWdp8fFG
tNPB9ackWL1LAhQaKsxqsLiEiAHEJX67BvhggBR6oXs=
`protect END_PROTECTED
