`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kTfGXQGNNITIRfEpm7VTY1zFVcWCWnQtMBQ2CIU8BcjIBCInQC/SZLD3lP5FImU
/JpHiVk0Rwre1bArv95qtRYUMBYmbKfGj2HYPDlFMpEkE75FQ4i5nRhOsZ+rH0qe
DnQvrHbORhKbEb0+xyiXkq08MxDT5cNTRYHmXAymQUsZH9T641Z84/vCy7Uwui0J
WNulPr9CLoyriYTsX+/XKEcyXhxaJHCQId/AUBhW6h6+4GQvC6vH1wN47zpbg2Y1
zGbq/6VORrAcEoS6Q9jmteIKIwHwHYSJWXaox/NthA0NT8NrkCNKGuG8H5daM2RB
iYVfOUb/S8PGaiEPL5Y3hipLvBs/BfswFuxSUTbHsxbFhXKNOQ2su26fqDQ5gdkC
ebvGmkTJQzWaeDTU66AZ0Aq90pwk5Ug7Q1auOQ96vuA8ClibIGl9Od1VGCOD/bm2
8ZOck5nOQsS4bi5317W7W0SBspUf3tDmtTubII84VC2uD/KOBD9L5ZrkLNFDMOKG
NGCb81Drv23kxw364I7g93M2fZV1KeK05xhcVpgBbmc=
`protect END_PROTECTED
