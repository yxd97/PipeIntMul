`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ljV9Z+oZ1nVwQYpssZXM+Vhsc9RCO/+I8JQSegq/uMBfqc5y3is5vUeW7fxW9mj
t+JqWYmQoN5X/uC86FCfcPjKlEaHPP8qycBVCnQEOOmFlWea7sRf/YCM3HJyqbC4
8Z+IHyWuCtrryLvFIDF7nYUNMA6N4a9kyJQCvZo2Fs9uXuy9FPAyo1wcop2wNjSe
wIvfG996y5/m3Vast9V++Sd/Vb+o19rrhin3VtfUpFOd+3XZs6ahS8yILjqZQzYG
XolmK3Xik9Ke6uhJlql8f3acVkUNtsC6+Iw1Gj1jYSF5GqESgi/mQRkkUZ0IYY8g
bto3xix+VMtSG4Z54m9NqeG5TU55EHZ3bgTcoJRZs5vnKLlbYq4dnepAr+vUxfqV
XtcNlpTAHrPMN6JNx7jZAD1PzBNXcE0gEHf6TUWbqB0=
`protect END_PROTECTED
