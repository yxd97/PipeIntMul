`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dyzmc2jFm8dxRhvGj6eqcBoYxReNFe1flNkGOPLLkdwZoOHWiWJnPz/7DyEMSR1o
zB3xtllm5GRcFmdSQPvqHtIPVzBWh1y/1PHu1svspswIzxm2u5vl9t91j8kI50hT
80UXt3hwsWijplOYU/rXnMYcC9Yb7g5G53bF8OsVAwK3xreStQcpd5CFLwgJvY0c
9JVrExT0qtr/kC4cJ8EyqBH+bX+pRAaAHgUL1wYN0tpX+Fm1K8pLxqApr0Ls/tTk
/ViD7yqVT6GSdAsQK/v11UlDB9uvQKtyE/sgMcygTt3cNeYXt3NIJbRnM07/+k3A
BvRAY3rSUsGj7R0+CZNBtHajR0Em08zTwQ5vVVxXHjn5bQZgsCIfVth0YatiWwg0
flx3Lra567fDyE83iKroksbC4bz474JhmFb98fiJsXLm0c4js9dhzO6N9Hq/Troq
8vV7j+DIEx0NwlDwnqY9X/6AxOrp3bDXlPBAGE+hCgSd5vrIFt3TJtnWuOTMfgsE
fBKRp1LPxKVNHKNkslaMDYkN3x3hEXdhQGMbXqxnQsNKkaG9y3tFfl936XryjuP1
eDWQvdH6xDcg9z1mXU+X/FoVQlaer2278mNk3R9dd2K3NbivJBeNhnsZ98EZHGsi
GR0aGAUshhzqY1rFI0jFJgFabthWj/J0O72JX5z47K6P0UbQhyYTYX/BEhcdtjgv
2Bfx4VHiaG0orqXl3hbkGw==
`protect END_PROTECTED
