`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycOhumxyO3BorhfT98lbDCuozHpW4qUe73gy/Kgi0RSTm8VK3ugSCv6J5wNnbLEk
wZScN6IMK0n3vFr5yId0DTpkcpxQUq5Zda2Vi15nQL3zZD8a9zqQW9F68ZJin8os
koq1iW3LXAC4WZ0OAmzsANGFqdomkgXgksmcANPEO+ynCY3vk1d8NqSFiduN9q40
aagLztB2941o9o2beweUAsdbbx9ctSaGN/UE6nwhfyqo/vYBQFRLycqG8aYMdS4I
LAuI672VeGwSleoxUYWrSIWV+7BEsk88/Fl55pzWsgx0F7pMEHE8gHGCkx+/v++c
IM2DIRgSOOCkSYze5n0vcJPFIpRYuEnzMD8VDQqzsI7jk5JGvncD9srTwfUdIrmG
qxgy2wWECeiXr8LTghDLhqbYYJ41rDbWsPckgmMs5G7cMj+byeNUnUqi0hsHEaNq
`protect END_PROTECTED
