`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
87cPgm9ZBg73WNpr56RPuwohgh1CFZpKcyJ6RJ78mlfACB6hFbZwaViSzqtFQNVn
LJPRoXtRhjmszD8HQL/3y9WNYL6Yg/sKyZJZkxmZQ9ZHD+6jqTRRjGYuLOBixWGu
eLAkK0CcymtHgqCgtcosuHTwaC9JVw3kOMDSCmeKnrKKJC3w2uaNmEtK+9ivm8ix
FNQxlA3G5HclTHpz4l3saZ44VTMIDgmjxKT50oeBaex9m1ljz0kovl5pH5TcyXPj
BJqxZh3Xr/Zj64wg0Aj9tbogj5/Rcczi+SrKrDHV5wkyyW9vovdHgYhM7cmEWcWd
t/qeLmzeBv30oVf3YqYZpM+qB0mLv+jso7Ux1EtH5ZLsDummFyg/gtLtih2H4LD2
r7VjIw2Y0z/s1qpHNJZFpg==
`protect END_PROTECTED
