`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yixzDN12j0+rVrB9jL3Jo9IFNDlLl4B+LRo2P6fUX3s8XbBiRzUxBdGa5tknP6ni
R8KnMw/+8DceF4AXDQaax/ujq3RZ6ejB9WSM7Ca8Lxi5PGTsowSMkw7m7K7sm7DC
uatqX4qrvAorD8IPRORr6ZbsPjlPF7T2NfizwP6ByL+qSG3v9UnBuhfjUtGAOSHx
+vwTcgyATuUVrw+OTtUkRpLS80piZHbTrJ9tMhfYUn1yuucJluWs9fzF0GDyg/Iz
7oNYIiVcWISoR/bUkSVFBYKFqdUO+HdnAT3KX+h1Kt9c2+H+iY2UxOus0Q23bSIR
RGqUVk79CXerKg9gl8KEIZfQRzZ6fJc1Y0EH44DSBiJ0DjM8RrEQUoVYR8eFxfES
jQWwkJJIF6HeCGGQhHbRDD5G9LhFHrijUUa1usNUOl0pE/2DN6o3yPjp4FlpuBES
j5Hgej/uSt3ogWZXHfbH9+sPPlit6N5GJPYH1KgIBXsD/WZwK/r0Juit292eo/2T
lSmVlxpnkTgRh6ZRV3aYQ0I2m0i8hjVbHHRzodmmFOjr2JHy/AKJJF7rillXuLWv
`protect END_PROTECTED
