`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XAlrKHV8jRVlcGpTgveNpVNI8cIfO8qcavQMkV6k4pmwfJOHhsWhlovsz+m+CJWD
j327s5NqT3QUEF01OQnsUKQg3eFdZNvzhK01YAxQVr4TCP/RpuyYUF1SNIazyNa2
w4+CmsZ7jeyKKXmzuBdIEGDy2oe6tSgfsxWy5rVtFHImT+mJSXDxwCIF+wCkHMlI
prhwqL8SoGa+8glaN68dkxtUV6Tj3YwswGACZF6O/XkH5qXQiIOq2FLqwuo5H9TF
2QTX8u4+wyWBTU+ycOTsTNW4iDX24kGwnqOpl9jTusSE3QrvTijmHDSbGRZwKSy2
Hgu46fxFDyzdwq/PF/1sLg==
`protect END_PROTECTED
