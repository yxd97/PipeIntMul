`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0CUBUFzV6x5EOIK02HVCvb9MYOZZzMPV2zcBQUmiGOrxpa6NIZ8oiJZEutRJ0vM
UzPXsNP3FzM98XjChNlhVK5gru2evPWxFHgOe0aHu1sXv5dlunQ/G3Fd/p1ka+KR
gaVI+ahSU7CFo4FAE8mppwm/+fGEkzyT8zSbBajdjiaMD51glZiJw0EO/R7FypVx
fdLv+AGXYly2KlTw88xdzkFyfmmANUUo41tqYFLPzy7+DdEIIV1E2RXvtgo/6IUA
bB2vNkfxI2uFoh/Zf4vI8lAOVQ+CUrEYLAfwKnHYRmI8SPimN0ZbTSgzgImPPWfr
1UT4hB2GYloHK+nhWQXOeTELT6nPBJPHa35LDY7afRGzWLpGMKHpd0MMnA5jit6c
bCxEFPGeTqpQ5x6M6VImoA==
`protect END_PROTECTED
