`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wwss3WEalc3WLGrIqXcauvDrTbXWCbrda/zetmnABkmKPf65PP5TezfZIornuIEk
SyfCzwwY86Viik+ibv1PL9I+hSkFPKoykhl27PrA8Fx7ZpVD2YWTv5E+KABdGYji
KJTJ1mU/3MHMhf8MTBkgvqlqsdyOujIuH5bp/LX9V+eAxwtDg4xeWhgh2JTmcmQq
ZQWmRQpQFfR64LdQNyVp2PEOS+1kAKEnWiC3mX/pmnGt080zbq2ATXCd+bylrFig
WU+ElgUPlmCmESoUVZc0kJWe5b3MxXRaG85HA7qVcNkdiDCs4NTCxn6WTEw0mDQc
dOwgTYkfRPUAPIr2lh6dx3EHddokiuZwSya7wZMDRWQvs/WRdgCZTOQM9KBcBIEw
DR1xX64Xc9fZz4MO9b7ShAXCgHz8Al9LDk6o6ooPo04=
`protect END_PROTECTED
