`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bo7f2QC58q5UuWt34jDdvgzGYLDySLbvkjQA4FOaC9f+8Jy5iCTqiVV1aH6Qr6ur
7NpQli/1dPNSl5WMnWfONDkTLDGUT3/K0tTkqtUJiInY6JuIMEZNMcUMABMmZS4j
LS3CrGc//NGN5glYQ3/W8FFJW18EqhHlPIDc2qO89xBGs8DOmFnohuyrD7yROejc
EwW4MUopepx9d+UaglrOuDiEAEueN3JD7rT/MMuL+YfXVQb6g8NgRpc40sOQi0j/
ztroaunVwoavHOTsIACpzFEoBwW2KuxH0GIusC+7X7ishGOnh6pb3+m65eqs0E2U
nH/Q1ttdrTFXzNnRhYbeHaCzZ53kggizzOfOn5q5kEK9RVMWIhdnn0ht6eCWv06i
mGuwW4VsSwZKNeix+UOzYA==
`protect END_PROTECTED
