`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRjZn+A5f8FVFym/zyXb8Qhlwu0gZrWF8s1UfyL4PIy+HKTWYI/GhF/mwVlAI3e3
gkmxBlUeQOrdg6bb0hTqfQQL1MDZEQF1Nrh3ACPYdpg7HeLyMXTe+oJVcEMtE/W8
QdHCbC+ee/Hp12WUsakO1KpttCaXA8+9LLxoRIhE6FePXLmdDgoOQ2Ihh6pVIdVH
tfOCOPJHLzrTifqbwOJ7lFwqZ2QXMKqZnXJ+B1M47GXZGrQn5b0i2SMSh6W/qnr5
pe4FMAVyV034vtSMeVToQaqXlL6GGmJsrQ7ip9WA3di1x/M7wJD7YG+w+vxbHVlz
PxcFRmUPhFt6DU92l0S1oi0hdizxotIJX6eruIL3B6cYFALlNjWvFGTO429pBNUl
qRr55BXEcsMVinS2Y7MU3bGxvY1l9zKxFjXDhE46Yhdq8E3OAObinZDJiTIoZhB1
bX651tfJZneEzSqNV4BgEmt53xjwZWC6jzBAWlE+AJW+C4Jch6JkrbOvKjxNalRH
H5g4nb0lpUNWGikd3U/1Nqj8elyvOFzfABlTgQ6r83n8uxvf0SU9McbyKuRSSmS5
rIdz6HDQVXBr5GoNh7S5iQ==
`protect END_PROTECTED
