`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJ57cxvH3x/eQqwrijHLxP6a3LjswigJNSZEYqmt/JoFh/i/VcT8z0gzsqSykECK
QPvO2bZUijK7EY7MryA1SBf+TZt15cElCRI/PdzGv32/UKltO8I7XMR07x0Rjgmi
uWAgPjGY+9UiMsRfnHQz/y1p5/C6RZu7OY2Snv+9rh24L9sztkLoCcIAWX50GVmB
baDUiPXj+gel/yxIcW1+da7Ilb4a3lRY25QFcYYyg2WE3IczBp36xkeax8CJsLEH
kYRc6KzrA1BmIcXDqxclNQ==
`protect END_PROTECTED
