`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aII06pq5lHVrKl85maPFDrOWG485co0c+tO1pPlqVYyfAFFOda3l3AS3F+3iAoU/
ikVpzu/Ka9vUI9jb1GnK52Z2LPi+YLF55k11DGvDU2u0164ynQAjqBv+L9SgUli0
1YRAxhG5LXNzn9uXNkoH+oyjYGhJo4JG60sabmxVwV9P9zEDxonUylb9sJWphkwK
nyxL5MrftFvqHmAfRkkYYr1vXBMBimz/zdR25h9+HnJuxdQWaSAX3mxQZBzjuxbS
S6HqSaBl/gbeAzxuLyb2M1KxOEKBbXWqBivgDr8otpqCbwZGRwihJPlLHuUTUBRe
EMXojiUDbOVL96EB4JSz7tJJul7HbLeT0DnZmxE0CCkrAIuW39HjB0oKoYzOUnCC
VtpDfeHGw0L0SYHApVHLFPrpZ0fXtceBTn85vnm0369DMei+73k3fMBdM9qPV9yB
fRL4/+CcWf6xVGQ73+DNm3+Poj12jyIkyL7g1bzhnk5MkPXhJTRoTLmL441BwddJ
KpKjSRc+ymitZ9JaZh+aqquIpKpA9dYfvuSGVpn5+UczuoF2yo9ZkXaaGLIjWmvk
/0iUQjJnsOKDhTgZC0/s5dUyx0hBGNHcdMBxUXfAvdKDC9SHr+0u9lFub4LfzgW0
hgtK668UGzRtXVMsqrykwkcRIQvBzuvv3KNUTsAh0Gxq5A36ZaGSR7CGKdx/1i2L
SzBH6pV3YT4wC0VgcOq94GGbammkf/oPHIUaQUOiDPfDfqBrDUe1AvZ1QYWFtCTc
D+YXFVVdkZ+JAk0wH/R5AdFYfTOX+TEaz1qsQTmd09D+sgfwqzLz0aUig7QrlilF
rWT4MHvrV2NiQ0JT722VFYSYPN3W/lEIEnELCbxF1XAdM/qjD8rCoiaYSluYoyNf
iF4foeBatzShkiTc6JiY7RX8Sb4+02tLWTNiw1/OHUhCKARA1lVOoyywmj/LVaOb
H8GwYy0qB8QHbm1PM2gW5CgcZDJx3D2ZISpjh4bSRDtgY6XPW847nfa/SARZqoH3
R0/LQiJZjAYZxrbHIRbm2mz2RcPbspLq/19kLFfZmJUvPzW6KkMZ//CF3lfC2s00
xMtWrPHxohcL3OeisvCyIJ1isaIqxTqfbYQBkZKrpUHGOtPdK2zoMflpVGk7CxkV
9kqJHNJ/+AMfJvSp/Ms2tKMmGWklKPzUfruuqNMtDnFbDGVv/3lUvcXRWN9pqWsn
tM3IuiCe7Fqs67IZ/TbftfZWWaHiEqEpN6fcdK2Cwb1s97xMuSnzlEH3/5VHcFVE
CwqR7Un+v+IgXTH1zJWF8sGVmIdSsiW5zwaoIkdFDWhKb3YnxnKCPeG/5sW9gTjc
2vBUCLxF94/yzFzzR1QpHj/+8GnvGSk6CcFPbMKqC2Iuk3bLHvWTt8TZh7/PtlE9
wdf3Ymit+ytHI88nyuyx5ZYN+bGExkaS/6aHbNCilOigjoxQEqSglLy9rJnBAYcz
28R7a2xBgem8fuosqWeF8KehDyxgZzVsUeWiN9JpVKC32cE2Ut6qVgob3mP3keGB
N68/7jOhZEdbtnKqFo6eiLuxUdEO54fYcyVjNT0svcqwwdil/vuPRxutFrlmMULP
3UAv3z/kIg9HjBbG1S7Y25ikqAsdRVtI+M4y3v3HXySrKe6p4mSt6lh4oSAUcolM
ZHB6ucq9HWsU4jB4XZrvyIrHJN3kSOnLI02P/vdISb5bLoyMnhlzpBukq2E62qRM
J5ltBb07hGCzcaMMZKtAAYrtbY7BwAFKOkiEuvCaeRpQPgVC4ZSJaAc9ncsT0Zhh
UNSwq8iwa4Zcbn8MZH8YalzwL2tbuU8bfuqGitTUrfPcqY71tndm2gOd9S0Ynapo
9njkcbC7ZPSmYUUsqzmXgD/lP/75tfZKxF/3b4Q/r9yMrIPw4ga7nM0kARy93ZDV
`protect END_PROTECTED
