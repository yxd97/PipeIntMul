`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WHN3RD3VPVGf8JfcEoGWEtq9zpUvYJpOK9RRzOsH2y+S5l8qzY/lrgqHsENMjRQA
/SP/9qctHRMp8F9TGXiSMbsqB0vUZFl5E+h8/HhTcg0evSMU2Pqc+QcHne6Vke0i
cBW08nPb/T1wlgJ+Y3rBbfyn0rypEe0TeT8B9BByrr9dg9XhAh/QJKqMxFxt9yq0
0iUQMZCZkAZL1oBes9NYT+BdjKZvwmexVEgU0bzpi+PvHqbhk/8YZ6HXamNoAI02
8Rifw4Dc5G1dduSy5wfwn3N0yu4ZOFjzVnAcjcHJBeacdoMEeSMTdipzPlp8ipy+
qVzUdvbSSAahr1AbaQTkHKbNhALPL2QDWffXQ3QD5jqBsvub4h+XZzIHGkl06Xm5
t/qGYPKX3CvANMnBy2lqHUa7FiMXYX2gMezwuaHiyETuLyerLZoJ2RPihd+LKtpq
7mpMhb42mdhoCzl4gmWnYLqMnrkNxDZpzCFKLTIkuBwk9GP4hhLw/bhqNspR4B3K
RdCY/CD0BlU5v2kRfkrJ1Xp/uo8RZkHj23k7/l9qAfo7u1iOVWqU0ZvZ365XHkDk
z2YtJJHX3F0fk2Jipmjoz+YtnFBhvjv0lUH3h7D0f2Vprl8+IF5J7RH7x5w2mEsZ
j5lX3r56pi7HnTIynAek+xiACV1Kioo82Wi8ou9SX1S2lOX57O01Es8Q5tyQammq
`protect END_PROTECTED
