`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
niECy+lOsipCMaYdVDEuccvdifSbYAqyrrrMKwv9/LKlTU3P85nVoASumpt9g4th
M6UB/Xkn9waEmnIjyUVTAiimiirpx4A4XAQVym+KKtzdGNUOtOXnXNQXecwveNPT
6ng3c2CRkS07phrQCZSEbFIfuVxHBSyMCe+HtwWZDN/dIOeHraHLckVhdK1itzzi
yk/z/kjjFqsEmofap2LQmHLBO9QhjOEOwC0hKEQZWx7fvwwH2f4C+JNk9746H05L
02juC8zagQMa8cRenWC3fBQgD0bghW2Ml21K6+QPUTRTrN1peiy0Ji1OZzvAPZeM
P8QVVMPDKCnK4TAvyZUudpm81vuQ8sxfRaQtUTaZ6n9zzx13/XbMHiXm+a0zFYrf
neQTuARAJXWm2x4bXOAh+g==
`protect END_PROTECTED
