`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IgzdpZs2iakBlV5A8QIse3A1mmaFmFWAiPUeU6TYUiPPFA1DZRg54VU5pM1exRP
xaLgDvDeOHWkfBGwEPig49CTu0+bMyB1WrpGtkAb4uNu4LrSb2D18qzpSqnRy/Qo
NaupLN0wBUmkkerl15pS9Vhn7DRs+oCb3YjycUbzDD3/aRppPTK9VRQmrGjdkRzS
V2WPfU5d5PrqIGWKUEbYrB8nCKPrkurkV9sadw6nCN2jruIgbPgMSTOuDkGk6eGw
Le7cWrxykil0qGOV8jH6igF1lJDW3l87G+BUYhKDNalg/jKdIG6AFAlW+sjJvnw6
6ylvgGha0YRdRRnPNY7Ml6bKclT6Fh6l+QCJn8s9Qlk7GhTUKl8K7ambTvsTKEeQ
modv04wXR7xkGHKgXtzLhzpBqmjbt/VvdkfHFLlZy43MSdxI+uWzjjgSmIsx+spQ
V5BysTfZR7MsVw8R9Cue4M33Y+Kjnx+2Ygcbwo+Es5jl0kpq7ofBuJYfE8K27Jb3
L7Cw3DKQi21TeoqatpFKSmvT7CT2mY93zC+yJWtea5GrcQM3j1k5ssGoZZWvs6PB
qXFEMh8ycNXQ99CmybmE3yLQU6wlNyssVmYT27rVU9o4s2TKKv6dusDbfKSWrtUc
48ux9qNhlSNt3mYMLRpBjymZ5rdAsDa0CL6tS/lyEEZTgTfAkWzSWLZdbnyw6gOH
p83GftnY5VSaTmK5s5/F7Xu3ZMOTfCA4TOOhz+l9aC1AQwZc3eqKN4B+Jgi04o1n
QaMqUaFyNjiL4990LGZnCgWDTzgkdv+8y+iX2RFvLP5eRGqBle/lwkWB2wlAGho9
eW1od4D0iZA0i7t/TEuh0n3yKfzbvoNKNKnyCI02tT/OnLN2IyfZJq6L9lTnv0Iq
8LgvlyQ8po5Btae/Mt9wk+eQByT8gchhin3c6f9C6dOPn5m3w+x7pvYUBCqS/MBd
Ag/0i+cblWOFauxPz5Sj9FzwvgJyc57i7y+xHAjnREhhBsBIqAiUejY1Kgy3Q+PN
GpJJVIEcMR/9IDxdPu6dCJbrEp77xGMS3BOlk31TGQ6VE450sFlHWlBRPwv9SgLv
5YyakvzROu3jUn4MkdRF7lOoUATJFtehkTC4QsnMf2VpOXpDwua+DsYBaiMjX4el
9jWEeqyhtj6mPaL7om4oaHadrKVcNngeC7KYwCY97E2cxzqWxYAaCimK1Sge1fa9
UIOvINCDijhIWp4YlmXQsZOWDJmWSw6u5uctQyG3gu/hnpGV+AZ2ggNSt9lQKE7H
n4wadeBfdMCuPDWcXyIRWkOF9xEg0COC59gQViJQOfBK7ElkNfSDqBS7OL8lyVfz
Il2jGHNh2uUt+nVfGqz+3vUv/L3z4nxMckTRzM5b/WA7fU3I+vYi9sZ9S6+mEA23
88gD1BfjPXrTIy4voznhmCuayLUYpmoebRUWOm8PwTU42etvqM+oQNKn3+lZVbHu
+WvtWmNZuXrS5MCS3Zuv/G7qtyqJNyVGie6b1eWrTz3XNDozr8bmP6fJRC1JnpZD
ABPuC8Bet56Ll3U4lV2+njzYIOthVrX9+4mTNBkNN4Ub0+nc0I77DnUiud0alzlU
MIn+W0wbfgVQkCdlp2W2B6hYGoK6MBWvCkZ0KakY37kiQ09AFVPU1PGd5tWprTrW
jl2Ry6DSA6XO+6cxrGar4odhS685HpB58Fh/lVkwH8jweX/QEPfyV1t34VuyoS+k
jpzwIeUVivd/h7eL6vN5vBztzhrvXIwCygghSgmkYfGH+mGtuymhpJLhABJcvv9b
12mIZo/kO+yWf0RePzZkbVEaq4sx/Zm6SBCAZ4f52jGcQWaakDPik+3KeGLpUGWK
8AKVWWZrM5glsxlNvqXCJm8CzFKV5fTDF2/9oMSHu7RrX+M9wXJM1vdnQ2MaFC5S
rZyVFD2W5ka7RYH1IGtpP4VCCZqIZN7I78zOEiI3InfwrInytMUG++ibk4Sz+rqy
jK8JPdO4Ui7imyK2Lxs11DHpGX9bwEqc/wbPlt5Tuiiag3IZ2AQwRFt3Baxgc5Ie
OlJ80tRuXBfZAq8SL8Nkf6IxmNV4QtT64LDyJvYZblZy0Yj7Kk6G06twVMquj+Rf
62eoWSZrTwcwyeo2lCYjeosIf2fH2sy4eb6fgysDuC60AgmE0XIzOdBS0eB9W+CU
GKM5JCL0omuISxTTrhzRomg1BxTpQEFlAGyzFS0qNzRwH7lwfUqdCKAzHk92qy8i
DW+XGImm8mJYZvEQf6A0PZ07jlwbt7BSYrMh+RU1lsYLZf8twk6InP8WY1XTwacX
IWC6vPFSGc+KUigJKnep/GDo6s1hECdk2zklBFjfTgEu9zuACzdvEZxYQEyMobH4
qqnHZiHF3Tqq4Fv16o8tSNGDD8IatjShUx8Rl37Az2YY3AA8k3Cgs1iLe/GdUbwU
kvx5bh3kd4Q3ZQfacr+6Jc3X4J0bTrl8JGUheoS7ez4zv+FMz7UncPKSQUNWzAoC
0dsx3jac0mMSirZjAGNhKkAM5Vnv+DynOOMqLOYwYKinjBHX5vmNzJncXjmCBZgS
q62FhOD/PrTONkiihkQ52BXa2D1fEypWC1G4GyW0f8Tib+JB7nRJAcW5EjefHpSK
AYsaJq3chz0KoG2YW3E5m3n7NgokvCtSUgCyUNwTvRoxZVDPt10jf92al4snAFB9
7b8N8UIGXW4v7XVd87KnN2VB8AtRLUNZSJo2874Zp6WUOLMKvgn8WVGLTiVq/bTu
i6uuEB49xJnA9FlboQRXeBOV7KvFlYTK1nAs3yeZI42HNRHes7O/uyXqDdHDxgiZ
X2mfpUWCU7g04zuMt1msKsnuDbuZynXe8XQcZVSrMzmUXqOj1tiTfsxiBsK0mpTT
3zkD8eSO3yg9uhI+jKc+CeNRXf5Msbt6QE53UTgCa0bfQJLEVfN8MVBtDpdgJaQp
q4X+PeOKbVPpTBe/QraAZ0JX7BaJw0YwG5Y+mG53SurFrx3SsFkwNN5VU2EKkr9D
Y4WHD6KVoG3jnIApAkS453iRSDu/EoEC6No8xIkh+OrUMuRMTSbP19iKcY+BiV3r
Xk8+2Hq1yR99S+k27/c/PQFKU7XyEgbT/7O2QbTs/d2B+tyGWf4AvzVQkFkvGwjj
Cmu+ZXl8ydELTSwKWL1dSzvd1JoyOcngH4fTY1Mor+53X1cjN2sjysYxKgClbhZo
sMccIbdBqVg3xK8bI2BNmHPi/irBAQ2SzARvlOSIcbA2RVQxBSvTIpHEEsUY3zVR
+VXCQ9lg2vUqViUMKbizPClcrNChaBZHW7B930Uxc8xE+V6LNfIAeDELr0nPHOHi
RGF4S45ffzIRgsure9dAoErGDlERi1JQShkzw+HXrq9KbdvfHmghziE4cuRiiCic
5eYHdCjJs+O5MtcP/gL1Fwsj00J1MQRL8J7wkcN99WTG4ZtqaxpGq/xlnqp7lrK3
8E+0d+NSlzRSg2XdZHv3ihVErvbAbeFVkV6GANJgrl5G5O90P+70h8X6cpa802ZZ
vfOVNBHTguJ8XuBo2l3/hGMDUBQIcEv1XEI+ssLYnPYVA0lrs7xR1dgm00N67JYi
AOEXSX7885SgJfAmCpVwjuQWchA1+PTYHpMhesrqVsCp03oGsuBsR68gHvtr3n0F
V0G/sTk/N9uFuKhfH6PGCyDCssfRd1ZbZdl8lHxZH0cj2YlftwYk6M66v571evKK
QYkcUifvpkz7sCSKpHWHLSIb+brdEqk11YS+bXguRYcH+6Jhy3b8MjAkhxWtdHA7
8NYM3GDy2Z4xUFReiUOoziqmw56OBhOh4OTq92SqMlxyEts6Jnu2Ns/Y0rzQoCqo
OdGuEzXX+I0DsFXLIWYDrdLXQZdHfDPg1oR5qbYDQv0zGbVA4pUwtDAFVGr70nTI
/x3gRfRoZ63laNHxanhk/4sIFbx1fLvbZGpFn1wXOhrTpAm84cWf2JLAZLdCQkLO
1HdcYTUDs6EO2NWQlvyLL9B1XP3ANvAkacrWH6CDxt3w4p04k1+PEO0uDwVmKWRL
OR+NW0vpBsyb+8tOjSwsXQHB8VBaliRGKi1sK+y/NxUlKVJp4XcqDGXuiLD9WE/T
r5dfZXY2hi0ACXrr41E+0+wn3L0qCWH/MPeYQ7eBTXKNBpte1rtAqHBvSCH1IdS/
PiPLSylmNURrFsjuFqN1gziXMhUcxkzdrdYUOiKqxisxf+AWdFH1jTI0VJa6ifEi
y0n0dJopkleUlWkLN+6wQEA2oFGzrFHUS0Hpmg0PHY8dRYdX6f/cwEuCs7LodanH
WiuxNcEJ8vQqSuIeWvcZbumMfgFD3mVS9g/wc3r9dcCvyo7/vBFx8KXjXfjupx9T
0m3aVUXgU7FQtTUQ+jZbH8TpCss7L7CKTA2Y3WMehwkqg61qozmZMX2Rwu2+xTww
MDroOmGcnhF0m+0Td8J5+7guYa9ac5PCxQ16Qk+t8DLg9YiVlGNd9/4kGWuty6kO
3VtR7Or17CM2EbARFjZOJB34O/PCWKCN9mskhi8l/IP8HRMa+J4aWZSri87IByUm
Jp0CbTlPgcWoAP5O6gXjwfkfzNTxRcNvmRCd4wSkdr/Bohecle3ZJB76EAKpFhED
C9emdc38Tqxck6HuEwy/U8BOxSmgwGMdjJk142eo0OnjhUpILKBr8VjxAe7pcf2A
cJ+TxAFFUj//gkO98AlJ3G/6z8ywvQIDZUllz4KbrL4VJLDHQKQB9fAYAPgIv8n9
TNCJtJSQ1OTxBqMwNl9iQeXSyvoYcJ8CnsSKRt8nDDYpQ0F1u24rwtCildR1UKrx
tdxmFebf3xHW/2IP+LO5URas35EjhD61VGQvegi9p+TgxsIKVBYgAqbnfPex8/5g
axuzGGxvf0HgeRlxxEVJNC5aWJ/B9E7x11BuLAZN0V2lFcJZl2TXrD8NFDwjh/EX
dHWKX9Ykiluqp8Q3EaotqpEDq7/llb1lTnjLD2tt9vcaqAl3TbYBCE60neERbDKl
UJ2aPzas5BUPvzsWkegVZ2yydZeov6kwljH0W/eEAIryb93Rc5jsbvOJ1H1yq4Px
VcbTd+MZ8Muzcga3Vq/gLSdvo3Lg1tGkS8yuA+oK86GcOYwRsAU/jg/vbtTx04kk
aZwmtWGEbIPJCfB1Cqo5LWey54dbOwaHyIOSJJbCfvles9+0egAyP3Udk/QRaS5G
f3TYySQVzyi2QpBdw4402gZ9VaqJ/KnDP/iKuLXmju4a2/9sRr3Y1vk6A/Wl//k5
k9xQslG4JP1SXumMmLUFJ/L5kqg92PUPYVOtZGrKSVUuwFNSx5D1/8kL3jQ6mPC6
wKa8upAxvvEIQumplhEY3zGnbdNM+pk6E96FgRMmy2uUlJAo2AHLbOMnqiUrEnvy
ACnNLu/ERl1sdmtZ0qJyCHYY+OlzUkipkl0FTn3GTedIGdXT1jjKNzNELhlylsc6
Xh4LwhiteSRzxnTW/1vQQFLFb0CDUjEswAYuT9TYMPNi7Ma30dQ+rFrobQXlRynr
YYE4d0bEIYTs+XC7Tlh6M9B/vVhpDcg93TBxJ9lk0vS3KSG3E2c4XNDtJNLBL9tS
j0vWX7dRnfM1HLmCXlmvf0YWlsKcb14aHQKA9GKfvr877ciiFsH7exyDEcPmWLU0
LLoIyvYbK9ynwFDvD3FUSlgLXaprVCzNEnwcX2omWsE+eb9pF86vY8tG1XAm90mZ
5+6uElJXnEORXoS5Y7oxO9Ap81lQrw0s70kAIuPP1weZ09sGATCRHwEsTVGAbOJG
PoAvoWHwyFLizwgV8FO4UY/29mAFVrVfydCWbTut/0aBJ0PaCj/lOM/idy24G7su
FUh3IB2rgklyREbaHAfo5pYnwu4hyqBQJNHgYgyAystJrLiMj4hu11qBFXt3M+d9
mPA5n/w03BT78AUhRDqoxiwu7PmOIEz+mFmIqKQwANhoIu6Qm9+waU1Jdws0hMC6
bjmtOJV+Bgpu935j5JoeYqFDPvzJ91j0336d3koOwqYInCNz32I6qUn0fLUlCWG6
CH/6+W7eQxN1prEw3qBFy4/UA8vwJqEP1KkU9sxrq/xpSWpV9GCjnmBPQ8zSeFkb
u/5KsaBTeK19qN6zSKFhDk8ig7AuL7CKOKz3s2S0LCq/TVg+1hFE9vD64fsl4Ln+
pNSewX0n9MDR9vUuAP5or8DPV92QLsy6R+2PJ4CAID5R5ncEhX468FdnezZ24BrE
lExgJgocmnJ7V9peciNa+/XL3zKMygr83LtpLHoACrmhGOZw5iedaLDUvd7FJ8dA
OGSRwuwAel1oOWPZE3gdyhQqdNhfmTI1xfqGZiDu7pwVP7gWaqcWTSziFF+oX/hs
wgyJhU5xkaBQ0gRb7EljwLpqGQNqcIry0iHlrjyHUy8mGuBhBef1CJATH2wPRilP
SNGFTinlzq26X4zfKrr91gh2j+oJgQkWQrUNy89jtp0ja8HyGk73stmydfDdo6/e
Xv6eyA1h1YlLBEZcxAuZDn75hM1Ql7w1cb/ScDQmwt3jbAy3KU9fAr7fIF7hPaGZ
ExL/FsaX8i1K3JxfTuV4Lq3ayFHPIX17tbYjqWFd3YaPKPFGS1EFCeN6jS3rbYjr
ayLV4EtBib3n1actYuyupm8ZUXYhSFZzMtGbMjI0QbGfLoFQeToES1KqRaXBIZKj
mLPQvtHyhRHvWHArk5XaTtPCWtkgpkZMZDJ1ow8X5XFSDSV9HgjxVr+s0TGxB3Kf
UPkVS30RkeFdmglHOkPY7TAoH5B0jx2m/araWZ+afoXgxDCLpVJgbJZe39VhqezQ
CyJYnZ93Ah8OXFtClUIHuvVP4vsr8qsYcIF87IDPfrHpqw3seDe4laZCwABpAu5k
JVUdIBibuXJlMRpfUxmQDjaCFgF38a0M9WCj7j2TGuPqkJKd0zFBsonXzB0mj4wM
pxdWncv3UHKR1jdTVQ3pfJvzt3aWV9ItoX3sXQnrmXBDki278yx3aiEg+5RQTfva
QRI9urbpIscRN3nWWImdwAly1HZs1M6CUKbGgTNcq99WHVrVdmvMyS3n1/t2BuTP
cFfa51euqelbyowUb9FDVDhpCIgduUx2cmWyAevnhn+oMJZlELkM5u67JmbY9qcD
6pjawsv/w7KFBF6y90c2gPJBNjkrY+h0M+LRNUE02Q1VlL7TTIXmVIRedVYChdJE
k7YhhDawaM5fQecFx/Cx9jcB1SLL1Sp3Lxwa9JfHXbc/4PHoDlta5hPzNCHhyclY
1KqWZaJHulggKH12NJWy0pJPqZJgGGZEmMJRP2kBSZy6a9i4U7dGCmYEqrnIzEVO
ahnU8q2Tkr4mDih7xTrDVw5gRnlBZmRA6iW5c8baMNzE99QJuR+YWx5WI/80MYCU
Jv8txE/l/c6O/k2MgDy/1u5JFPjH1kgSS9chAt4jsnTt1ItXZ57AG34ciU9Jvz0y
E4QH7hGgVO3bBBGaOGlWsBc8/Tbf9W42/KBqKqtOF1klit0+D+DISpBy8gvvwHs0
Nr2qBFLjbMh6U200REtvZdYeTA5GS33//qAvTaJEW/y055QqJ7KOgZs30onMKBAC
4/ZhecVGa3miAmvYu4nh6Ug8TWrCg4gOexv4Y7V+UJ5acA9paPQryxcgyyR+Rx20
VuI6vcYvZthbb0PmBdVkcy/AyL8Elvqj/9F5mf6xWYEGAMz1kb3Wiwk4E00sk3Q1
inEGA6ZJhKE9GVyphPZXtKUVv0NhSegu/uf84MwzyNfGjV1Xv+JMhvj2dfFWYOeE
Gthm3knukGV2vaWU7oTjgbcVpwXxhpKhqm8eN3gfuk8HVfBnopihCysfHQBbIIQj
LHDV1vicuSe3bx+lVBj4nBDYQvNUAYiba4ZZThZl790I4YUSlmtesFDhdbvz9HQe
3BeGawwIsi5sUIw8ls9HoQLwlLhrgqzM4jtoNqV8LT2c6mb4TU1Xskj3FBeYT+sF
rkpZ4CFewQkC6DYAXexJwqu1HhtW6rz5MyyBpKkX0qrRltUx6m2VbmabajWE0YcR
/9/YaUnwTQGxgPpO7Ywhn6ZxdDDDxp5r0zmcOyERsT3tXr7xPONU3BMGkbm+yM/+
8P0wZacF4dZxrL0DBOAPsJ9Z72xndRNQVT50O5KP3ouirpa8NH+zwafBhiugqSgz
qzlfn3Zuje0yPBQ+75W0r8VzV9JqJJIeEQ/m9IeZlAFxXMGNrpxVVQIHm4olhHmS
LDwQLF2CNVGwtIPYAUnAiT6rBL4Qldy0bTGmXd6T1lefKeVmjFtbI9T1w54LCB7+
JMxF5DXFMpxbXTbWujRcULrcdGhuaOGbrsnqSuKHvrVhEJ0wHG67s0iPlhIm8ET9
JokdawuaE6x6G8HhOuIWTF0KY3m70pfiLHEtJmJNUoktgab+/KiTOcjsvMzQdTZ5
uLA/qxTe0eUB9uh+7zKlcpgJwFmNjN9Xsg7TwmR74b+Zk5n/0VV2TIolCEeILt5g
5ZQN93uhWZwdr46BX1ivr5ABz/on9CeDxpHKLqnfgbUQZlYygWsSZ6HW3tceYTIn
syJc43SzRWTeYFls/NYg6s9OcaxWTpiC+saduYnrvTJS6bgGA5ujYk4aIoEqlMns
hYCBVy4yyk6XEH68OhHpSuxzSTBm1mILrX9Nfx9RCbJyBjW8BW3Tb/QLldEg1Wuz
Rfj7V66Tb48QQ9g0G96Z5jOUzFPycCzL+YJ0GPorwUJC69AU2+21N0xLAt5bWqIY
wDM2D3kbonCAZPJluBY0E0B/leuD4Ys0pEszThGcVqe2Q5r8mStgf9qVor5Xe2hS
UW+YT8mQiFiZHMO1BVqjEgiQ/wTgfLgsyxgP4gwydwFObYZ3XcsInXcUaKGYhGCY
KWfBglZEVlhS/K/9RUK1w3EpxJjw50mZwleIWoLIlwPS8VhtzNYsbn7fdZ//sQM0
9bbI8onXrGyCVoZbQcFDgToDzTri2a2MTgqa2MUXSE4ACQaTqtN63MA+/9+sM0D0
JNbCESSSopQL/9r3G78Cr/4jpBpzAYOB01a2C7BpcKgjEFKbVOV+xc5R2QlAYJ1H
Nxp8hS9W9qjJVtsUSZCbBUhh0cUKVH1BRK6fwLz7XLR22UhqU/mVEKNX3tQp8mQP
SBaD5TQeTIXxlItU2JU/stFa97u47oI0ZiINxCpuAG3qyOv0hCVgmO5/TASxA9O5
t80jntgWeo6W9Vm5HI6JLjbsYfOnATDBI0J3GBx9WKEHvj/fSq3m57NjdCSQU1j3
8qXa1IC3UEl9gHpxZ93+BIU6yHx5aRvYyqgo2OwhMFklmOlGUsKTsrmz4yPVIH9i
ethI6c3k0c8aZTKnHnXbv0MpQs3ATz13FYmZmvj+pgfl5CBPxlJMLsnCpSISVXRt
6ZVFHohlQFopteLW0pDdWJUVaUwaSo/6AGONccrUYomCsrnGDMm9ysdliD70EA89
IYFux+dXimlWyPiDBTEj4L6zg6a7zAdjY5QsH/GG5eHZnaInCB/dVODySoVqka9T
37TI2Ckw3yJ/vqXz2XcUvCRcL5OPizBgmEbaUuqIjcEIUQswVBvILalhFLLQToPe
O09/TACQ8uhDAAbL5i2jdgIzUUG4qR00TOnCqzboQNAuWkyAhlkYzTchQFnyJQCx
C5/xF3RlA56ob2e9QenP0StaSjWFDWX87X8YEvLQrVaHKFeAhGTmvaX2WFwv33fc
FntCcge9oqF4zXPlToYGc2qXqm1rBGY4MeSCQRvScewgegSjR/pdNPBIz2pEUsyt
/L8uhmKwVMEALYwyobu4DTMWLD4cDIJELsNSNaXN6hs6v4E7jbUAEMZQrnRxhhqc
u3CIQQU3f/oEmZeldsaADaJyUvsxHeD5V1+GYTNUwZm3r7KM04RvwecWTsjapem7
zZ1eDiqeRHnSktHp8/5TR5EIXyLUyqxQ8L+5DFfVhKVqOlgtiS4JV/nNcXinHdYk
6eq/fDwlTKHp9nf/Bwz9wo1Lfrtc7FXyZ+U8/pUsquIH8l29+H9kvwyKVgSVuuDb
vWBfgm2mlxoC7ZQCKAX2Z09+2jojxtdc0INkWpkyB0vOjfKhvwfO/Co1qHQukta9
h6KRpXWrjFoPJ0vIw66wfF/O95VHLXkzxErinVL1wDSSei1yadQ7gg4J3ik8db8Y
BWqJvNgmxK272r5FTWdALQuAWYB5JkyI0UfKA7g65E/s+aL8Sf3DN06DzcBRquTX
o8+6ohHk3XEyiWdJ5flXewX18NmsoTFnxV/4ziVljFWq2sqKYh0dTJfQqBcORmFe
uS9fF16fzZ1fpoVX0N7aYjA7s9V3DRmVxueG0vQrFbVraADimDM1CWaM0CjnLKxk
i+A6GTq/Vp0ly+200RfCLyQyjvqvrIf2DVUBlo2Iz+o+Cg26eu1cnZw6PIuY1Knf
vqhGpYwmj+Vj3MQXCvg4owHptdqxhidNptuvTemp0zS7Wf8USmr8mXuuUlB5dEPk
7h1q5OOt3sGRDZY3Zwom+qz3OI6pnVqXAHMdcRiOmWxlQIusqVjUEgKSU0VPIZZ8
G7yu6M7RAzo7UHUtws3WnoxRlFv26wgttvoSTVgIzfSh7H+TPIufkYtsECXo1ewR
MVI+vw2GQ/r9RT6LJoyBxatG9J6h5fcY0kdOoUdR/phjCz5XMLtinQ8/klfAEzcB
Shr52MOpb+Bm9ISNJ/uwYmUQr9dCDhcq8fyIDfME3MHs6Izj0YpSDmvNluqhMYXP
Dyc//CNWS52ei/a/+0eJyRQy886sTXZn6YoqFBWNasHWh1LlX++X0J3AuBkRGaHt
+UZGWHYnEL+pJreaWG0cROsYBSyyHCFrQBftWswde9VcSftS/IpmrylsCPSJzcGN
JpP7lz43EeQ3YwCx1sEhLZn0AwBBXpX2qzs2F5QUligfpFEaLLob1ZN2LzXlYX4K
v9dQDCa8o/jT+3poVuvTcIR53j/X85kLxtK2KbyhMm00xG3GPrTbQIxDLLQUYJCF
FFd40PI4ZfWTDW3NsnC2TetKNjc0NWauKfSBPcfg7j4pbM0TfFFpa8cPybZeQyxU
2MMlx8WNTtCID29h5cPXCpbdOIq8txdJJ5Nn2BT8Ul++VuEcDbl5C5obNOlwO2cU
Ce4Wy0nIswAeNcbvxSC4s5VoDnHIgfeuWC/asgRzqmsEHamh4xx2v6MEW+iCdLbD
3ClOLmjGbEGW+M/46nyEBroIhctRSM7PFJMJCxEFzQDinv4kyJjBR+Tx7LQobiwQ
VLgfwZ4X+MmviUpMDeixn0Q1T/+FCSfUI5WTRTj3UWCcA+C+Su2nD0X6lmdDDgk2
xRXCYEDaeGuYLwGAVZ+op5EjwLszoC8ltXmTVCIG3/+BYTOqJUgTVEbG8JAqG8a7
iwDR7e5Y1qHp0tg/D6SFMjyPaLBVOMaCC+SaGxhAAfVeKhjng0aGDHrmRAzyAJpt
JlGz8O1JEjzJNKA0vQAEJG3WanHdK4sCSGcPq6mRgSVxAyU7BPfqOaX763UWbxID
Q+NocvLVWMD9otl0xWkqBkoa3iYVzNDYVEtqdevM1NKaISBZLtqqB+H28S1fSNtx
7aEKQqal5yQu8lj6DkkZUAvhwoUDaFUtWf3zyei26XrkDfHmcReAAGKfbZjtG2gR
YE2GKGAx4kL8ahdDb7fU5Rg1t6MiuX+ROA1smPR9kHxYJwcC+TpZz+rfButzQsKf
ung1l/mxcmfDmScZM+FJvQcl9eSFT79WFYUvtIVAW6M75KC4EpWYkT6KxqThA625
xDWH1ccnPwxz8LC3VBTYKzNGAcdvCSP7mn5EeiwXYJziJWjW7Rbcd4wxehh1nNmj
C4t13WLerXmMSIKDy75q8lW/DL/vbAabauLslb1czkvWm4393P7pmJruncz9RdnS
VSOUc3xH9f/AYNebrrecCWLZyHwLTZK8bwkHRYyKxGneio6aNM/t4Pukg76cFPjD
VfZ6/IEG9Vu8sxaWMVRco01Z1bOdOFIuZ+S1Fez/Ks9898de21Vti7U1Z6u9PWuk
r/rxNUIbQaX5K68mYCjZSh3Q6wKRPA7UxysN20OpEUoxgogVDFFJoWYabUu0EvGV
p0goKDSINixlB94L41dNcGV6jVuQoNU678i9SB1TMBF/Fd7CrAJr0wTJAuEkdNI1
jlWY7k4g8Fs+M69yyc0qZnAcHwLD/3VOm9zWSWC/3ZtuiyyAePxaOXGffspe0HjW
K/Dz0m6NIXCvvFKpc15cHL43bu8zouguQKlvYjmEsemjGB1SB5FvnMG8siIWLeZ6
G3Fg/yRed8GbnHUp9tOwFzskxGA6h37qUIZZkTEQFlNtVnGAxinK+jdfoLfepigw
aBuP79bRQe3P++6LzRWCEU2eBxJu4Y7S0rRYb+yrOp/Ua8/T1ZMHWHh73YKQaAZZ
btJG80sXW7kQ0i+8bYHBRoSrH4u6VTl1+0mFOOqPAZuQvHGGte9mmw6qBeG8uVFi
NqDZsX4FGpV9iDyB0b2hFGybW+fLIgud3kXKyvm2JvsFqoMJgnyeYgr2t64RXen5
pYd611Pd+sLSa8hMHyUfD0IkQCacYqYMpC2Mzr4G3uOuJsni9BZt6dq3bDW2UE7S
WQC3IKOO1w2mWLFknmCo6kQLbHvroSqR9GK9jAZTPXYri3Pw6Gbi445BrCobBVwO
CD6A4hUIKTzWEfhL4juQ5zyM8XzSjV6n4045qKOhjUw=
`protect END_PROTECTED
