`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3m/Pm7Q0d2DvZQOP0dPy9yd1VkKDqWIzEcfxkg7o5KI7rNeFQoabLUuVvWgbUXH
0agu+tCg27jbvRhMrCphij7m7Jlovu3QqGBAKVroODpkbaHze5qB7lD7hnkmXJ1d
e0W+RzfRhHY7JyACixedigqS79oGPyPu4VKlnObw3yIof8AW9S1hesS1p4glmfmq
reSazAcdn8Ji9e8gCVOPPDWRyYVsz8dW2j6IxvD0dUs9D3rHpViFpWgALaSQHvZM
na30/+iLvtRezbPaPydPfaqnjV+mWgeaxfUKit4ztW/LF+pEKE0jtUO+RY5lnCQn
stssady+Ys3qUMZgCaG5/iBb5aKSKyJHPOvMYf7odjak32ow0g52xBVgp5c92S4O
OXwSJ1zhkcfaucirEwKLcPP8Jb77jkuuUEDuqAignJdrX+QkvAEJ4TApao8CgTG3
j1eMrewuNIIDmM/k3r7m+Ay+g947hH+1ujsUHYZJE2oGIQzvyTOnr9UumxiKWkVs
1CE701OZT3pLFlOEVY9b3og4OFnwQhG85Ff9owjDq/PFJT9i1qw3SwjFONgQ42E9
xfZ+vCsJzAjyDFcZ+1fVNzdLkcdPsyNJ4R76qQW5z7nqTfkdvcNI0aviPNRvdHqj
bmYRNkwF9v03nEV16cjLzgZGxv7aQ8GJbM0elW1F/SEhVzYTqOGnUWHFIouDmJ2Q
8jUrn/WmPxfn2E63pHNlWX8HjhZ40xCMqW23TQLJKuOcRxs6TTnE/Xt/H9Q5Ymlt
18MolLd5+NId8YxAGTuoDPcQ4Xavs+aSyzcVFCAjcZVusQAYyGH7A66owCIGBQAa
ua89FxhFRerKE9WLnFjHekB7P8PRsYbNoYk+Q3UDKHRMMSbk/h93+o6Dd8QM0/BK
4iK+Zoy/4EtwI0kWJ0r42w==
`protect END_PROTECTED
