`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxOqMKU+U94ha7PLmxYfudwsgL1zE7jAA1WqtHXq1vsdm3KU5Lk5gP64jMUhXz/O
epoo4nKwX9ElHuFlVaBvsMbn3U5RQhrmCq+oACEtDPwwKOGHEs4n9Tgb/0wQZj8k
mMT2g8ZkBYYH1xkhfAGjvP3BF+6dGx4Irhc1F6TuFRHtsGU+gtGTWxN3Pmzf8MA/
ppJ+BMCKqNR4jrWzEIM/GbuMQiwHThhdyNQC4oP+9e4uMSdcYwvJAMIm9nil16GH
wfFWzrpylH4gwIrA8d6y42zmqr9aEdV9DPacP/lw5pkSG9r2H7V/AjK73FzTspc5
sk/qDmNiW81jUDLIruCZAL7LIzL1ACphFWzko1Pfn+gxnn7dUNh7gcmMuo23hXFN
9lcE2/4hdVrKamTVzFjgEZs79tDgmDu7M0MI1hRGv1+rz70ZQMv095mo0VEZoWlQ
8efiAupe/XLaW1AHCva43Q==
`protect END_PROTECTED
