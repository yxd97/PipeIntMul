`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDTEA0NU6e0uIkgXlBMz2kwWAOgEwwEmILoN0n1PZD2ca5Sw1FQET5hoTj2of+PC
h19ITNkgUOGDpNmgaR25KE2heUbWPuROQUxH2H3Au8qtPgNsgrFpRmK71qOebby7
Sdnx47ZWX/AN5/K+1XE5S6sJRqH24huIeQPZM5CPgel93CyeebsxT6OZiCvE+XjD
UQYyMWKxo1+lSkaGUXhhYTLqMpKscYgMPldn6xCTxAFMaah2x5elSkN40R0JbCgm
RZ3w6pFAEenm+cvhJKjhMJswFtUirV7XRZCaHdipJS3OARPa5taOqLHKDMMb9c0g
raem9OW06W4INQrPfLRD4RAuI9TuII/8anK0Y1iNOGfh5vPKNVjhka0MDpXfYOCb
KygWdgRd8+CbQos5zxBA1i1lNB/hBVMZ1wrQxWDvVxxvfHItKYD4aMiVNItAZ+tO
iairlhW+RcxLzDEFT2+jWAHjSplFHYK3j013RrjGIeZCImEE/gk1u9byxjvL6Su/
D9tcizua2W0K0Ign7uf3lrXdr40TaZa/ann2A5POmuu19cEDLI15YzB2etk1yT58
hT3CgkjrHBX3y3WWZhBG3IjTUv0xZ+6VIay0C1vto2g+eBDXGcr8woaGTwZTRMva
LIMtCrzdfLRB+L7b65lcfIDJueITYIyqMDcHcbzfzM82LTH8KnkBNmOFFowCAl6d
s/BJZIlax5Vnz+yDFXwzQbjBi48r4vuGZTqT93awlhmnMm+1pwkjXfBfx5MJ/AW2
ykNiUYwCw3PwNJNoG0NzKl0cigoU0Hbnex1SCkKn7Ir2Xdig+lHWNM8Gv3ody+Ph
HNOGSqx25VWqR5FUN152hxUaFRH32gjqUmvtcOvS7in9U4WyHq49jFUeuNNdBlOP
ms967d4wKW5BSispyeJlfm6hh3hsPYJ94oM2IjTuh2UGA4CvtVBF3laqKhkh7BG1
l7hRcb59V6wKj8YjLcdEtEZEPoYn66WTnFT6uGiTbzszzwWTJS3+Q3oSWU2XHWah
V4y7DYrQRzT3JC6ojTytt4TMzbVEHEXk7jiZ6D8xh8coBr1oYfQhSuY5dYSbFxSM
GNgSR2w2A1Uk6BJZn17VBstkVft3pLiZQFCvJwpcSJBOG3yDHIekY2IhJrvA+Y/r
IiwlCEL3tLJgl/HtVwwTU0RcPQI4d3F1n53Tgl5MGuNFetwB79VIZZMHHpi3a6r2
McpbcTKII2TlVyVcKFAHjeOGVhRIky5vBxfW/WrD9SqGwUqaWC1kJh213kH2NOsp
1ZWmdFOK0QLUMhStnOgTG3vAKfsO13XsaRsA3k4HklpnJAjk1LlhLgepj3ZaDRUD
XMthkwWPYYQB1v0L9uUEbGBcIYCVfW12N9EtP/k/RbFul0XkAT0uT/i+4dCHr1T9
doy2oTCV9ScafWTMn84jk7uZnBpWvqoDnbRlYS/YYJfKVa0WYFs8gtvfDkY7cQTE
t8wOas4ckYUqFqTJL0l1DQ/mgaJvFvVkCar7ZRL/7w07SO5+FfL7cKu7K4AM48Cx
kzSHP4DNSTF4r1StSbjS+zQduW9eOtAeUp9wCdM/YcIgYaQZ7+fcgBSAQnptJtVw
6eM0tpTmXg29goFpPP46gbQIGCenaKUkcSdnPz51KAW+fIJFJvK01D3YOr9uUuqs
zsgt6Ju3BKGfEk/wWXUceU6BHyJGutoCaxf2hnfIHh+gSmZsehcEi4HNesvc2Sul
06suXxsF9dLnJ0FaHFmKrAe4Ekm3dmvByyQm2Ej2P3fe0JbwTziatPM9udSEQPJt
f4HJZXPtgjFgP4fQse9IslKwo4A2uFCeYk2VT1HQnP5pY/CsGZQelZ/RW8hVR76Q
ZZd1KyBsZzolCIE3EbtxI6v9yTYSTq1SaYWgmRc+5ztoSTWx10KFjpcbKTSwO/cq
+/DQHsH7cpffaFe1XRIvrN01ApyubBJT9IuiaUUhOolXm4Y/H3IUruMX6eAL+mO7
ouSJ8FYMvUDdbCwNUWBXN1uir91S6WquVltiXfQ8bKz5jmvKjoLXfKlqRIDvFbO9
7bZXbZ0+GcA7KpvOyUo6PHs+nhpFTu7ElPwSjbeMWVfMHe/YyjHW8NBoxlvwZmoZ
Y8XeQCKWuLbnne7e4n8QAw6JezxKeQ7u3V70NZCH2ctQORjIJTradCQEZcbsRrVe
sTrKkh6udGLFIeAT2CyC6XyOMdcM/IeEEbntzL7erQ51IzrJGDj5ret5P5EAAN7T
mQEzimna38H9urYLLFA7VxPPWDeVBBdRVwrjZArcf2kSCBjQ0j8bs/RhwI/3BSvq
DQF4PGYIPzMgE9EHIYyP1yfAJ1seDs9yOk7QPnR4HMecJNCNmjW/tSRyVVJg7MPW
rUmBrX6VGkr2TvkabPfqnnazUw6yZPQbGoeFqvsWiz6satS+ijxpGkzr/SYRdHw1
Mfk3JQnVB8MVgau2BnI9m0MvXR5pr/Y2scxDwjc3UkU+IcwzxY8pKgEBZk/UIQQa
jTSPK6WUe45bWTw+Z8fjR/1O3yDnJlnBJLX7sG2gWgdwiFEBDV5vtaiwyVixDUM0
S00UQApwyuDdLO08jbmbQb7ZWiAjUqa6Fg6w35OL6HZGk7cLQPF6U8JalCmF6dkw
HBABH4UusO5EK0gLRAnMQ7J7TKVOYxLq/FyukEiAnov6RPm5UNHHbBnCaWRO6hP1
5ByJGO18Ffszn1R2gK5Ov0yZRH+hKDor/of4CbFTpciW0DjTG2qez/jZyAKXDPmD
GswD7o1UUrxyCkLIArhYgg+yyQrmdLwFr//LAZjpWbb3p4/DZ//r/OcDPra7zxQz
sgGE4uTmWXr8oujexx61IH0S7oil9ZHihJxxQpV+xx8MPxQwUPCg/AuUqIhtORO5
k77+8hkrxD4KrJ7FTwg1VLOrLWWrCsjJpMhQ6N+q2jzSdC8/pJqxdSqaDRO2GhEJ
r8f9gIXdXsmPkyATE7QXdJzOxRy1MCVp2rBDIhoC5I9iHfgpXadhej4xWENr+sih
umVjav9OfOzrjsLOYYFvKiQAdGxWcQLOSykpaoKiUCq6qq3eqYdU2vi8bTwjh3G9
5R2qTsuQ67THd4DWb54oTRl0WzZuc6bTfw7N9AxoL+E3yNah29vubQFRddt3VMDZ
k27uOM4dQEiv9SbJXW8UFJGWVMt8sf7mg0qGn1VHVIKS2cQwgl0ObwufDpGvaSxw
RX+OG2wDlrCCQZ7+5W4d1MGEvANSMB0scskIFs9qXNUgv+BHUqZYSv78OxukfbiX
SVDVItvQ3w7xq5QZOOewIQynEMRbahSyzKnfSuahsjqXCUcpar+UGwiiRTCknWP+
spUT3TX4Fwt3r5UrLwQrFoEue/os+ClqZZawLuJmoY28RdXT4H7ut9ab60vjMKdQ
WRhjWInrWCb9bNWBvlrgGJIiUCE2AwOS9Xo/jPlUS/vIqKa5axFUUkFDHstU22NR
ujHU/bx73wdBkanFUEpE4B9EKaPIZFc7j3+WkSGR8X4f/OBaBIyvUfMfD5+AZQHW
lzsUeyb6wobKcsJt92oiMn4HpiEXmA4GajMVhKuLdMLm6JK+mddvSSYqEFnOFbae
dfC0KGZn0W6DY1loRBkyadyd96pmdJXF4Pf+YmNmt3qIuIALHXx1s9huwYEv1fqu
Rpo3HHd/b81ELwtASqSOZFKhi2Gd6gVO77GFtqYSSdiX23gcM736xoe1u8ebeS47
TqJsO2zop2IWXIE9tm7b24JxLZo/LSlZvW7KUGwY4ljNtgnldIKarO5DIfU1/Hzs
AstNPScY8WRBD0cPTQNRInVBrWs3bUEEUxJNHqiVLf8CUdnRx0JIXIonVUlfqNVD
ugbo8ufM3OZbQVscRCV9qOOy9KWfy7lehXrqbkqPl8hpirwvEQQeNTxYewTNLl4w
rVgbf7QYSSqbrE6GOv4eecL5kbJrftp6kqY2w+13KJ6cnPHG+/98ksG8Awq9B9iB
pTU5Ouw1ZgfAl5659A1Zt5OWVwEQjyCtC6CFApm6p8Kj+1ELxO9VStX5Ena1JhMm
tZYDjd6ZlzSv/yS7wT1srnnofdcmMv2WSJdi3r9K68i4Tb8mrugjF2HkJsSGL6Uj
VFv9unF+rrMc+U7/RP8vwbkoCFTM6rZOq2avboUbrcWYIqYFdPZxGljs1mBBJKpI
UdRGqLrvGd32Dx109ffPZ6mjXaQ5jUIqqUqu07MdkBZ7t9wG+y4RiXzWOOT2/Bx5
rfSEg3UNS4ECLwgSvzONt+UkNxI5oTERNRzYrevxmUn0yaQcPsTbgmzvbVC9tMMV
msz1XxljMa54E3OyMKTnYxmBodTcEczYHIPqGJXkzh3CprT3zocb4jTo1G2B53Ni
xWe6q6xh08PtfjVPw9rRXkw6/60w8FqXMSnmVGiQtsb4X/OX7fskmt+Z9sJZqzP5
0y8pgUp+DyPauTC2GM9Yd6tc0EIf5B+aVMSJXzUgSHXqEbRmX7lTc50b/dwEmMnl
bDFQ/3QbraR8L8HeBW4RnkEoqjsB7aPJ1azSbQ6tVOgTw9KaTRlEUUsvcyG1xC6W
COnimZPEAIsyg7SNbQTb7yJTmBhcuakkAsiZ6GzRLb4CCtiaYcYzQeLXG72eREJ0
Fe9XJqwJpTZXix29JHrH0Ph4DnDB0+8ZKLQ3pYpArbmjzqHDaeohayvIQmxnqfRM
l4cH7vOk7WA2rxsGrvj5scuFvid8ER0OENdnm27Si2VDJIKpyvPogks+rUdMgcqd
blSGnywn+Bg81kIv2i5s2BRA2qDfcnw2l4AsvM3sBszJ4paD+gg7V+4/nTQNEf0O
fz/qyE5DUrZCyUZmaGJBDWBka3xjuJnWTVAQ+rRVq1YjVMNqLuvjLltXd457LUYt
fIeHwMpo769nnkKKAeY/jxEOHY+qSg9uouzlFc2sh41A6sZYi3WDGlGSaADbXepp
/Y7koa0dJACiRHhGM8zpMZvpsNorSQlAoMX21pm4NFPPupa2BRWws8owFsAEb3cQ
R40arMZS350sjUrA5V5MvtBKKtuP7JevSiZiAzwiVqn+BlgngeL1xl3uO+s77VH7
QWOZGWP2YgkmjojW6c6LLcRSvP+0x3KeZfu0roovAqYKJgDTdutJOgEjkYeg3hVH
zwpez+MXn0uKYfCqTZwP8KxRB3r1/3d/zWUa8nCNVn0LEXFv1hE8z2rTTPVdI1b/
N6SjETf/dR+gkks8sMoy46dA5lvZJuIOmQ9eCdcSMsCkBZqLzOvDO0AoIqkAmN/I
RjRWllyJiiIgVRtLYWvEP0Dpe8nJ07+fWUlvkzApLvxm4Mxysv5RFeK08ssWfmiT
3Yms/xQ9yhANkEHNoa58jOGJyPpE3IhmARyg3KCc79CEtfcm2zKNQSNzyYTg+4wU
2P6ByUYwiLPLiawM83jJ81qGiWPAwaDxN8r9+NPCkqlgRAgY1qEVpW0PwnB0gKv5
2vGbB5TFmLnwAui0g+miDmcIlTOPSucmm3eoiXN7B/rVZdVEktj/GLDZ2D+Tldlc
sR7ARhnSF99admXhms4gukI29FV/IZFGk0eZkulfgtbacSyvkIfQw/JbQ++uRYBS
6Hy1tyeeveRYUQr54zhPVwkSivdi8DMr+PviXiY51y1ZEIZ8025lxhpIy7L6gabn
UEpAKZDGD6xyJO+5a3fLUSvL85z/J2+DM9MUIiFTIw+3E75ukmEkakr+GNCQOO8J
EWIlFpgC/inLiovoy+9d18cutZp4DgyeIRIZnAqulZXczxHQ8ghiQsoEunT44PVA
pX3TSRM8aAUAq9ZWdwZWY0mgI96hBkvFJ0dTGOxFQ7XnZzCqFZ8jyKJgxoI833JJ
wzuQIuRQCDrf5K/wCcEU3SE+XqYGCrrbKoEagW7wDmXUEnBCkAWlKpmFV5DE+8A3
3tbDI1ZJCpJAQHFIUogC8K01LRbMOeqDH7bFHpd77oWEIpU557RxkvJau/2J6ZoA
NWYEKkhpV0aKW8uC4cNHv7Wk1146RJ+B8q5IbxAl821SnJ5d7Va2p0rQXjfpFec0
/HL5SVE6U7QS/x7gPL4vEb/u/ldtJaFi1RDyEFxBEBjH4h2ciizPEVEtFMMzQC39
9EwxJMWGCnTgteuanet7VJyGKXG6EOfvPwhZ1VJzHFuXGQDkpJlSzyzFDxTb2oU0
CWIJ/2pPdYC/FqJ/1ge5p5I2OY17E7w8WJT5rnWHFrmyX3KuR+5vaMShJVgjNh0V
jxRApzRIefEiFxYTN8dkX0tNMw9/cVglSDRMeGzCE02fZYAEK1b4xvD5YItpGQea
na9g30ZwA5i4TS7DHxc/iXFTuQGQFxCCbl80uAGGZR0iK1YFqmrhSrFT2EoBMKHn
M/tcSiMrLeM5zFs8IT6LGgcSzkRRlFN+uSuoO3QyexNQ3ciRKQhrOrcMk5b3EKLC
OREmzR5SxmEtjCNMAIWmsZIOmGkWU+vszUBSJdckV8H3d/iLCexJYDg2OM5sUGfR
My+IPZtnS9A972j/6Eh7UnWBud8eBxKHtY6gNyTMFVkniL9+VBAu48SPVdZXtMGJ
fGj+OXp9WHtyJCb3OiEpAH9weLUvQAEHKwRnFsSOhoYBSFdTLq4bhm0VwNZSkcCK
BMZhw+YzPksawARAmnk65GS40sOf4yYqYEXFjQIO3YpqaNp4cNR6lxOwG8MmjBWn
WXagSI34Ckri0ZHO5u89W0KU3vM0WB54WGIX7jar/nE+zixOEd+IHI2mLAhHvm7S
3/LwnGizvJMoIKgrlFRM9tzp86r6kyuzhdtcY30h+8CHp2Wtwd1EpGEIxNTgYeKr
fbu17z/L7PBfY/YCk3r2vve/Ly226MEWLzowcGGTpPJKhOHrmUY+I76pdW3N/fx4
YwoYhaQZ2IJvZLTrhUfHGH6FhjWw4/oRdrq3cGzY+mWQU4Dj2Su/SBcJvHy2q46x
8dtNRvZthrTQZG4hgoHAZ/WKnmp+bsp/UD707gQVbnKWQoU2uW5N+bYZ7LtBbt6b
YsB0Cm+P5DLzm83LPAjG30GNni0f64By0W+V8MZNSyVc6/iY6wHLIy6UZjCvRF3A
8X7g2lDZAr92FQ7xtSGIwOl3y9ro6twIwGfvxYtPzTUMCoLUYO2Fnci5YQhHKwpb
2ORuRHQASPAMh3Bv1LVminLqQnfJWEE3rxQwfpIGOfm+jYyAwwqG8BEP2D8/jth0
cZAdzntVaSTSZf8expxNc4W2JeE7ULnfhBhmNYMpGV40JKFVxUUZ0fAbdXOsj0+m
rImV+D0tHGOMN6xaigOb5XL9EPAH/Ax4HYt86w9wJyxqtyQPFOGV0yTWPjJrvwF9
qo4aockddOZxJhQ2MMaPZ7+Y28bUfh2kAfvtmEYtmY8rmjOcDu9ac+Du32tioCCY
6WxiriAvuVw2QAodSo+5d53lzJKQ6F9NWNEX2IBHnVCohKQxJOut5t1TpID65tYL
eN4UHBN/Sa9ONURQYtMWwym74uNHr0OzlHIPoZ1fnYrLFdxZyuWSPnHYPG3uyMl4
WeQ7xn1qkFPp003uuD9hz1ae5YC7vp/LR1yS3T1wS5uy5POznwSokKe9ionhdcw0
tet7HuNgPmA8Oh8G4qOuu/FroepK6dFlm+wyc7PPaAMG+nwIWvwFVzU5zJUOvKLm
tGnVEFdZ0/+fl3CDCWpJyFH3HR7QQzrU7QtcM4ZY01nvJvR4ocz/Ldwu0mjnf/Ze
Wpzop4+Mc1D8KHdSjVXtg2yan99hBi/v8R3Z5xSkHEHl/aCPjOobovbRlNT8Ut0o
C9njb/eL2Y18JAQ9EYJxBuUVNxD7eMcsNektimBySSQ+1OZqPPQVgi4q+nAoql5L
JB6Jv3L98PE4tuoe2zgcggWLCHCMiXW5hglAer8es2iUEeQeTeP+QEPEgsg4Ilyi
hNF3HKOIgWEFSUSK8wilQ2m76IhudM9C/RsmbfRmzVtgFfOKcYV2pXxAPz1rMVb7
OQPD7lC+jOCJbX4/fAY2LzvFAzbmr/Jo4RVtYY9Bt54gXXnAWH2rWn7LCMvwpS05
U+pCn5At1rUBsuKF3a+SPhib8PXd12aXCVUrVApx5j8RcRi67mALIIM5PuodotYM
ca680RCKvip4llpap+2GO1z0tFRprEX+Z82DgVGR3SqdxqlODYSuIbaFV3Ec+55g
GjX+zlI9tKsFmb7roqg8ldzuGxMnZ3F608LdwXP9ioVdVIPThgsUR0KYWyKl9lyT
iEBOhGrywa2HwQhBc7ciXKu28Gicx+vzxNVzWXQC9bnwfLIXsE+ZcjQw8WivkQqS
BTvuJ5mgh2mzvTzgXw3l2FZCqOvhtAIaXT6pCKGuhXtBci+bvW4ax7k6OeRfVXD2
l+/Ur8LU4nk0gL3cnf8YP+sn9S2sEf4aArvCQss36UoVgCI0HQRmunzFxjh6BQmf
yCzTeT3kh5lVfarKkZd4fGM76x6TSvh5TF5UaX3iJl19C4x00pIEnBhNdVrt20Ft
1JsO+R/kTpu1RjI42uz7pTeukL07c2IoGnLHWXx8N++QarQiyKejL+nf7+rNvVBJ
Kfv3wH+IJzjrCGPSzYkDi0oTpjUnx7t//StpvWdGR5LNGhiYfGjVyatOCXMbYaCV
FfLoLMWuuvbZLpI5F31oUyPXr5RzR6D0w+BjpTlu3X2DkcbRYQ2kRuYBlKHZar1+
XWCmRMAY6OR6QSb7QyVC3Xx4TAXOoVGEU91eEVoVVmyxYYMKObYO2eIDnzaeRVp2
xJuUFtFZnHXX8k/9xMmKKy4ypHre7Kgei2RWz3wslsOn8ItHQUxvwRrNxIba/wX8
5fyl1i0Vn0wygAudZ3UyEUt6IcG0hwVgsUXWT++GadszYJsREGoW/LSOfM4riJvV
wwQ3ARdsmis33tBdtn854YLw+17L1vj/9s+055Akt3VLVMqz/O9PI35RFaH+o027
rn1pHLA65jfhN3yXVdKLojppr8ATS5lz4FgqGIJ/bhwGNNDuIf/04RYkQruRW+qw
erRFRU9Rla+CD6USSPoCAwfZDE7rqs0l2yzn4/qVAl00MmGsw9fL29AYuk8Y0g3s
TD2SODaP5sVzc7VsaOrFehnk8Kk+m12+7AM7tDVjq1lW/4s183CtUnzO3dn0pTa2
1xQoreEoJexg1ygYQ8J4w+0GuGQOpuUC0RjxhxBX+pbE9v8edKdPZx+sk5ZCUC/i
3lUfqkBDHSROKXlphNVjt9zMyj/w+ppE3to4XLm8rKW929NpoOeBcU9zxwALdFty
ljKUYHZbSm05rxEg9ZmlGdW8ZgvXY6yRFNnY5d/aV4AOkiZxRFPyXac9zjBbZntG
5oLtCA9aP7wB9vwOQVChcjm7soiFK5rkcX2btPIMXmhrdY+JHg5nYSq2BlQclhKE
z2336Dg+E1hcMd4/CUlUdig6/rlREm2oQ0eqTdntl3Hw0n0E4IucnQ+qukcCmo8A
ce9KvXnRaCOLZQs5iZ6RZRGpksnWBAxqerNZyCY5SJt9KGZSnKWPuWvUg5+jHw0R
CFkfoptjhV7voUt2sNc/EDy4tOsZwhwuO8kY0YfbeXrNLl0NO+P7ZegJPwqKkZRS
LhNj8Y0OVxxCbjXArNrqJsv8q4lbGTCvmNNEkCTavznOyGlrbp1YJJrM8mBAA4/9
06VQ6M4EsCzb9ZzoKaCydWXL2ycAB9n8rAhTNDDJjcCprl6llhRGIep00RcESZI2
ggmHwU45Cr80AxrOXIvgGcylevOmdghiOvMXxRshZiq79LtApC0hkt8jzwqDS/9/
yz12kn60IaLailN1kkochJAVFHdjQ6fwuAfVyY1OHc52iZL67y66kLKMDL46FPRw
mfZPB2CmfZU4B7syn1wBUdfRMX+C2BbsFoNQZjGxb/u6F66Sfs1hzoPFCru2XjzV
LW4sb8xI+FBMtsRdzsWpuyxIungP9EPx1D1Oks/wcxSuUBX2xfCvrhUELrmPlcz8
OvdrwCXB/Yl1RxYGcI4U/V77a+1o46y9+c/zwuXA3q6clGAY5wL43xxgaDcdUQKJ
w1BZ7e3UpkGdsjOxCeK54o1RpdfZl/9dlCCDLu1C0nWh8WNT5KyvUUDoEj5BkraJ
SW3mb3aCayZL2pu3etfMj7UTOuq68Qm5bBpilNEUqniwmOzTQHyCf1TPflz/sMKo
WT0RmE5VGLJAlogLXbxWM2tujcQJTEhzBAGufEz+8ogRNzefVJkM9iyt2AdH5M6O
ccSn7euRVkPPPOw2SVtAF5EX1XnhXmrqg3hVgOtSXM7MBxZ2d4dLKF3XMpdZPVyD
/IyS4eRR66C1mhs3RYM6MYSgT1RyPn7z4Ze2vEHtX1Dp67QXMmZ2/vDJYbRKvfLM
7syogM6kREZNU2RqfmOq3VUWJPodAmTN6Wy3ly1s3M/IoX3XUGGIWyR6JUYYj77q
IUnjEQl+nZ6Oh5SkzB/u+IiF9v6cZhDn4jOP6BQ2BWK6XD3AZ8/hpxBGy6K+T0Vf
3echntIa54kcED9bo5NgBLdHNpgx3yXDxJWh9hXyvR0BunAdmP23LRNSKYko1XSv
w3eLxEVsmLKrxPleKRK3b1DpQRv/fMQWKYzQ6vTDlJNMf8XQUN3aUwAd02zZa3rI
KMY4Wafm5UEZzvlLuMy65hDVJwwrA7goaeoa4O/TL7Zrbkxz2qDnp+PZ2dHgZ2rt
uARtpaWcJsLiBn2SuuxKRQvRCcTzSL4B49l8WH2KlGCgm0xC1giUuJ/QBUM7luNc
0k+enot3XfjUwcZ4cq+qehqrejtnE50DIDCbfMJkKAMdazpf07tobKU5iaOBUMys
A46iYjc3E7J8jo+JhO5x9RZMKBmiTlx7iv/VeXQWCoEGTXoylvHvA0AstN9X1oQB
4GxKFfjKkzkBFCDrd8s7xxJmYVC9yvtvTUizuFHmxS36Bm/RThyz3JK6QcGjXgFJ
wwfDIjIRXyOILGfBINvpADYz+9kShRyZ7nXNERu1B6lDJpMvMuXwIJJytFKSAnZK
B9sLofBffUerM+ll6U/05t6bVb83xtH5xMUYqi/+yA+xUtyQIBw6IEX2hC4dyf97
/xatYDp3+kZY1wGZZl6Wty+jVro5xPFaFP606FLTT2MtZy00cdg4bAE4bhPGfhUe
Y7pCj88Q/jOWqRzOGw1vgvYvhwMUnmyNJm4gEt9ogWa5hymM0I3LW6iFs/OedpRs
K8CekHWoGES40L01/TigRUfsxp02N0VH+6HCmpugMchwZR2NtJu9kkQ++WvMZjf4
Dk/8G2eW7btNYRpHMaSfQiXwpqYzolkWRlgNeSDCRluiY2Zq0/9EiYYkv4NwNnE8
8c+/DI5uagMU2YAPxHRMXbN3X2UkorHmJAzAORJjCPvqBM3kbpJe+s1Re9H+gA18
dabDfR9SfNQ1fXbae4eZXeLPYVXgFazdOhvXAiXiT1QR9609hF1AUoBI+iKdrnxq
1ZKfK+blJzcvB4p8n6aSLFxd6dh4qE/LXqxuTTIQsLAOw+74Y9t86xhJfsF4M+FN
OP1blHa5M20fWFcHxrWhdXdeR6rpBbV3KzqrirnjBkITDaO32khdCJZDdqcLAV1p
CcI+HfPrXZFKhGkFOT3LuP3SX6jzTE3vZ8ofpgSuNOR/c+wvNxAKVV7YZ7Vt40xg
VOJ59RMicH2TDYa8KsXmfWlVTXmybNrRUy1hxACEpO9nUvI592z6TlzOjnNrsxQh
NyY7XHPm+MdwaX/8FddCv49nPwKqnu0TLG/UMNvjaDeStwVbZIRE8OZdB1JSxvRg
O5+XcoMBjlIr7zBqpxTA0F3Unh1EBmCgYSbBHbFpx4aXDtg/oJX6HYSS/WpZhYn9
37SatehHfMrW4fgc//NEQoyZr01zXMo5fuI1wPPhD0zERAqvvex6sfOp45DzTv9U
4fmNpDqv6DRoUCFlhohE3S304YBXJ+qbjBnz9Yen6YdSEVQ5l3B4Q499/gNcdEQZ
FG8nD/s2BqnKJCODxkZ2P9EVYSJNJ/2wjnu5yH9HmMFL/zeZO5SEyfHlLkBugmJW
8KrTCwQA8PTXSy34BHRY+s0aML/bhf8Sq6iTBnYXlE8JhfB6Nn6eg/FMsA5ZCtX+
4daIWDzjy4uHoAJ9EX1bZ2EbM6sjdjq1t3H2wSSvRYenxYPIZkRXZSdrrUJDKZph
dSe+jO3rq1h/eX9FUV7eVNUuesfiBvCb9VC0K4jcKrf9ALd8DORvln87ScMTV+01
Q0UtSyS6fuDAgGQ5MK+XaJmKUdY4/mjP82FrNlyy8bXuwdVzajzZdCQ9y7KOCn//
jPoUdqlLM4UDEPsxzmD3tomUl+41l99Vs7YBTsb77A7ZrGLOeKesWlf0woXxTVxC
+PKQe58K1yV+5Am8RPXS98wQLsnqJtpXQXATYtymgxuJrbY6czIn7/g1cN+q4rZb
4XAP5jQ2l8sxgms5RsfUesMD0mFUEc+45GVLYjek8/qiUX6fqsNLpLkpTJbtIRUm
BAPNTxl+aFLh0WLI8yp/9cMz/9nrxwp/5zHJfctxcwUb6qhW8KTdzXe2Tk2V7/ap
mdKao492Pl5X7ozLLRyD59FK7P15mvEXAdkPImio3OHREQ4I1rvBw3CzY4XiKuVL
Oik83ag1wDVK4hflqXlD9prODdP2hPCJIBXTMmf3MlzaibzzbEWpr+j+uVe85b/d
BXBFMhVSwWUertBJ3LBd8iIftZ8l6uI63MjNrSTOVO/HR7+nYG5GEGmt+zFZtW3p
woskXlwJ3RZt8kpx/GjbWAU5XOjCrIe+o/1e9Nhr4OmC7JwROUfvqpIm+QcR/5yX
XDX+CGFVObP6l/ZT33e8LvX10VHerO+jnb6XdAz8U+Igeqvr+k3JS8y4Bi3nTwBp
tjMnj6Fmb2YGR8k6ZQXHWCkIHiB9dKR5AnfOPHwtggzoRBd9hswstJQTyiYLk6Ln
IDH9O/xviKCCE51tZSPo3MzSaizTGAWpLarltwTKoexk2ry8ADygiPgW7p+aGfTl
vKJ+7Zq8PSJiCLvqgR9DtdXFTlhn5uOuxzTGtrPgd3M125Me4B0RpTyqd+rdciza
eK2B7VEhZStICH+zX1flWxMH1atmzQWnskWo8NB13MKaBTAQeDCdY0G3lK5hnByN
zEwc3asUgrLE5DkQf9htJX+tvoMIYtHo7/REGp1TTgyWBVrlylfWaVgziXepNCoD
LDzsUy+cUM4yYnj6ChIa+uWBkzLSQQhjFiGKZxf9h3Qtiq3ClZ2SaMtTKsCHIt5+
5gin1Eq6nS5QSgD8+tI1FV8TN2vTT8ZWV07YVZoRWmNeRWIkrAB4CYf0WQcIKj1s
8pwYfHZEaewR5y8n1kD+7UosihxBlPoDW+DYBV6/FK2Dgu5DCbmzHAHGbI9dmcLQ
b+94c+tZZou/whvqUQdXg+pwV0OZatV1XxtbdlMbxsFEx9Yr9+FqbDkLQOuislxO
zRiRORy9cmzche7hBNq2KUdU9bxYCtC/c1zdQw5gw2HhekD4BpKRxafvBtRM3kEM
MIrQQHB9BDZftQBFhUqjr4Ytj1wkXGJEyuQt++m9JkH2mn9Xa67VOP02iqVVFH1d
QX0GCDsxnPRpnzRxsYZpKLr/dru/h1/j76feA5j0RIy8/qePSOjo/Wv82QG995S5
obrt7fI7YVbLl/vCVLSyXR8YD0fmWIMLjv5hnZ2kxti/RxbQ1gQQyT8XYPQZWzgM
Ot9VJ4/aLc0oqF4sGQpH6mXMwTKXR3x/pzuFI+brEZrgOAuvGvvR0NU5+RkhwokJ
RXJGvrbRLDdL6JdkORSEkM2+dsNIihK4EOPpDg5UdqZhur+9bmBJDAYf7AcqHcS4
5V8W73oHfRIwdVGY9J0xfMfHmNfx87mPATrhRJHNT3Sr0m1eeNmblXV5pdQrdqnR
EDqev5x+XcGj1LKOBeaReDGD15BXeFK0itcWv2FuqVhi0W2Ep0AVrrgR/gr/GinU
VowkqbtUwLLC1RtZsywnxtpajqV6+FjN0UhgJx53LWRlmAvzG8SsdOBqgGaIed2q
WAJYCmU5JX5put0fUVy5Xm2PrUK9JRBi90cLVzDNJHLv8XXsIWGzh5KujfyPAwRt
NiuguYD5reSECbWacS5GVqQp1IuCHG85xHH1W8QlVQE50t6gUdvFz8j/IiXqYnIH
XFLLeq5tTZulxgEY9GqLCALspd8XcyFoHfRn+dAiTuQWBtSsEYMLRn5OWXmKooo5
3YhszackuI64qL7Rm/ILEEP4f+GQjicHJlkTTJCarsB/ftZnj8vLGrqgrCdvcqNV
N3ayHQC2rtyytrIKBI6bkCPz87sYc98ig/8oZ4ProcSDOpGHkYrOoOoqthpymJrA
tnT+/wqJG9GwEKeq67teJYILaH28Wo6/trozV1qyyGondeRxZ1unSQQ8z5Y2OcmC
+MbolGgpaMoUvYcJ/vt02lDniWCNMSE50SgGW9id5/FumC6ulD37z1e6Rqlwr0wM
erePQj4gf6vB4R7pIgcp5d1asS5fe9q5mJGfUTHwXNmNZg0uBDzT7PDHR8mgVz35
utYUnSJELxdqWG7HvkoDDLBX0gEGg5NNfSHD1IaWaXcablqCRE7+OJ6fRc6mQo24
G/2igkopY6prGu2pMcuGsGA1xHFNmmiudISaZAFLCxiJgsT69WYS/+A0xHi+29Ja
04NHjI5gctsNv9XLWuxmIofGASc+zu8qP/V66eYqCD2lJ+sX/iEUEoLKJQsRD5wL
3wj6tbWnxTL6aOJc+qR5UWWt6OQDcuD0KEuth/lKhxO+5WCjz7G0X0PvTD60llmB
P9kKGA8LCD7EegsqoIk/HJa+0MhLXlRlLC2yxaS0HwXunCkWRXmyRA4Rwim/5n0M
5jNl7d+ujCwkG2MMsYfwGft1tDl3b3fmy+bCct+wuOXdSR9uhm9IYkhff2/wMklE
AOQa3ME86otT9ilvWyAWqYua5ReABadhuo9lzBJH62BB6jtP23PQ5Z0s+ybiAArV
BOt7a5uM0w12CmONmeESzQzd5e65/ZVa/q3YjSUoZ1vBd2qqtUobIWwb4my/wkM9
qoSY209qQdvnDSkm3D5Sr+ZTpaysYn7aUekRvaqfwxHlqhv95CfjVXN9MyMiBE2M
prBq3hn+9zyLCMTFOoHoF4UAsZyAUSMgyJA8KO8yz6Vv4V5ZI+CabmHP4sCveq2Q
pVPn16/f6+ZqxtLhLE+2BSzlHDghsOWp0M8fwoMmR7YcSw1ue3q12IeAyYb2keg1
1WDUy50YhqdsB4XJ90di7wA4DEut0IX3XBIa8Ku5lAM7TtXeUKnTOHMkAAHb1LRh
gjkrSs8yQsisOV4jJLToSeuyA2pOT/wqJjXbVFm/B/wTGge8it7oQjVD2kCK2ShM
7RfvUHnMDteuezICzUSZpWh8vG9aRXmjyNXHsTDhIJ3nbK3+x0JxoN4+snmR4cQI
/OKi1A7m2uYg0FEg/GMo2ZNNoBCbqniImCtEt1qcR5KXIwRdmYDc+dHHbRre+zJY
T146nWh+wtTiFw8ntFwlbnbB0XcfwCyZXzMsy0ym6B8W8MyYTqGlbuLScfCqOvPv
/pSgteLueJxFP9XqESRMyHSZqNaZTTc+adFnr7O80SbdIPJozcX0dYhgOv+s8B0q
AdNRARaoT+lJXBKgaK5CoPQDhN6IOavF2dqjZno6McjjZ9iGrY4mAESjwWakNNB6
myDvQsRn6eCl9iApkxUtz2EESDsQBNItPw+xo8TBKwVwkn4wVzs31zEXuDlfBunw
vUdLqZH2YEPCNCd2mHVdGfUWAWnOpu475fTW3y+hHFFAII6vgopocnolzx3Ha5Lw
OJalC/JRTrgvf0HSiqA4PVXl7DHMg/oVXqZwyQS6DtAhMuYKwh62RHJac3JwhuAE
PMFDWMvq/3uArI3bUH4gOX0CKzB6ybIyi1zCvyzLWRnCG4r4ubZVh112D3lzdNUk
3gKGkfjOPDnEBQUQVn4MtcERcTZ5d2f521BZIupXv5f5m+X4HR9kyQ6F+62+v6gr
j8IwviOk+FpsnQKjctW4M2IDiCW+e5ZkDk3P7+yk9cYJLBUv+OC9E20Y8JlYkTpB
uc2WOyd13wDB05RKs1SUwY5uGYrzlGoJYSTTbQOkW66iJCYHiRfgm8mjcgi+Ey/+
/67Zpyec3VbYHWXiBqRx8QHcLu0F07uFtZmQbIhLPR0At5eBmRdSCCEMVTM9q7m6
Ce+sPZC4OZjyGrT1k7lgAYE7L44QgA1GSBkbbwZ/C611BCgyUESSuu8S2L0IsDTd
UvpsuZ54GQ+0NKxHFiVM7JM3xzU6PHcHape0yo67Vpb4w17J9iBq4MaKKCFf5Xu/
t8FX0+9PZ1K3CTdbeMiZk8QbbC/G8AuTym+D4D+eGLUtSjGLbJuypTHwWxbBs1kN
xOgY/6TnSMcVtVOwzmSF60CIeM62XbAoldvatxzTirRa4L+q6viHK+LbOGnK05Tp
txeIs2uNy4QD97HEn5eQi524wGC7v2xXbvd3v9iXY9D3P/i+S/y1oRXDKkrRMKlg
p/7Dy/GyQVGYAL2gn+3HRxKOLD4nHZ+Q5eu27xWubFY0ECtF51Whke1/TdJGYmZZ
JOmqhyLgCqHF8+T1UQI+mv1dr5uW+g7tOld55ABMtEdhL9zsAdJSz3GX++AaMfiK
1W/KOVYcra3xnOQ0cFaYfGQwal0ihrM9HTqXqsx4WbrsnjqsbI5snBoytyLxtVdr
PpY/NBSXpMEKeKb6CZRl3lhKg38c/uYDleE4NNmQgNC1WWTNaHvcHjKqeky+U13C
p+aZK0ptJiHhDczyGd4u5FfmUovq8frZUOCine9Yl+i/Ddi+1nEaTw3V8p1SP5q0
qJ6zrPPVJZwLpMuxzSo27wYfEhK+l4h21Xa9nNbs1hBNR4l40mQeqo9lRud/yVOf
mDg3PhTeKW30UwhY89B68CADraNGBjCHc05SsrvntddvqK0BkAtT0gFdainjhPKl
gbPV+J5LtI3D4FtPbtqskfdGF9NHQDs5Xv6XDKAH36797I40M4bJAYCQ4320eObb
yNuxq86jFyXD6ZdbNAjmJfoLwBq7UdQk4CrR2AXLGPU3sb7AhX6CIJv3k4qKkkPg
4wUHCnHF2/RpBXN70/N/23jU2YrPSXgoEYDSpL4LGPvEABYP5D5YV0UOwWGdXpOE
r3q9o/FcxIlI7tvxloaf9gnP4q8V8WHRGLW7CRyrGeJybcdM/cToVKEF5so2XWZT
ItwAMPb/GcngEZaAfbt36fs+GDvAD1H7IvHXDszDKxmy/f13hz3UlEDx3JKnfl0B
iIsgho6OPx1KO+gcaJlsPh2wxHUO8WrK7CWPdVhuab1cIYykvWdQWOmhExH+uu9J
Z0igERoqTTrXE7V0P6VRSuGWlWYBgBrMd67B9CEVjTrHKtxDdNva2OJFe19IcTLL
L9YajFT5yUmCD1Jyb757yNVBSZz4Z0qSeU9q6ZKmuMIr8s1gEkmxRTWce3N7PxVK
cPJ8fA3WzDtCzLqHQA+MmB8LyntJ4jARkhBj8KsS1NdOzkwVhcHZtf6baD3xkovP
uAy/cWLq2KSfIMZnlwmGi/ZdXbc4onAvxOKTBa1gQ7UGJMSRd/CPpoolL/dip1UL
Ld+EXBHnDjs37n0qP2qfvjpabTH8e51CvtHpdlDhWUmN3bvgBJ+7SW4Ub05ZDqLL
ew25B8pY0ALC4Rt3kex2cZTgnEnY5NgnH+zRQWC0yA/LLAPnynyFvUQVG/YzXVzN
93ad6Bc3oWWPqTDLAUsl7L7Kolzz/WyAvd4BSSn3DHdWbzNMx6NrwmzGwPAIfNcj
I+RFFoMrNagFrccblIlo6QkK5dqc2JipWx2KH+/fU+HNQsiwa+KLlMkWq78K/x5K
nm0yOLpGwLUu7iuGskkEsVHnDzZCJ+jLS7RKEx3Nv3hosiKLJu3eqfhdTvIG8uod
0GmgdubhAPrKWs8E8jJ3q9ZBZq1aFwZo+Uzro5h1E5BneBxuWvHUjDXTH+GeLhBJ
7PyUFZM1MIguEU7Bd8RCtKbVUgoCmfHttdroabD+0CZVtF5eGb74UK6cspNLbC3j
XSCJr1vUOiJfVgIkZO+Em2f9uUCKQ0WwzRsyWiQLGxn+u/yeFg/CBbzSFSJ9hBpO
J7MEmmE4gL3UE97P6v0eDE2Yve1004aCl1OeFSrakG+h3tDUpBFH76XWtE7xvAR9
oXD3zAxzxSyIBaVR8VrnkFbeyR9yDUjoN2B0jEGdxW6bcW9HKF+72Nuce3rUfZHY
rglCt6mqvr6dY0SkKszVlZnaSMdWYJlHJpGZgVA8MBctktKm1SQDVxbGxQ99cATJ
glIrGwuPejq21WDQngpcaOATbmHPEgpiLT0GG0+Y6neet1uVGRLW8gZciMgqTYPO
qBBbJ2s7Uu2aYoi2l7dfNcICa3rs+e2lnuNaJHB+DXHEiXwetNKpq3giWz0GlK6Q
fER901B25YT+WQwYJFBofBRYQCl3jp5zzPwinGeiqzm2ID5iwpFYECPDaaTyY/Ch
QNX+YmTHJToRQuojHH9Tye8o3d4H10JQfDPhRFnAFKZhh5wIXqMAFLn8oWdbzDCm
JRw01YxuQBJXQrRVTMqu4xE4vUs1oCUvU9UFlPWl7yFRSRkluy+rafuAI6ZI5VQG
dQ2ZTYgDULOAaB9EG5BES+ujkNNamQkaUsLY25VZMLmlAXbGs3fq4G10UIcT9UPG
Vt24TNtlh1FJ+MbkPOkGvDVGloZTPXASO6lTx9NnJch+2CUg0eW6kM0MUpfumIOu
m1v8ananqB/4DjArZvWr+Z4JMhLoVPa9A4CN5p0fWrLjA8nXxGwI41uMKF5tAAQ8
t2tSAWmNQnWS82oLgANpdDonXZjmvGjjq5hS1P5eg1htnbg10P4ZghkAkbq8/IiE
VQgw4TOba7uvkU+TMVHWTrSdbFhpxpKoHPHRpdn/2nuc44hthyIvVYvWDyOMQLZE
of6hN625aJVFfPHzskamTh0mPbFZwdhKCyc1UuDomR6DdNIaKocX2cSMLWe40OUj
O95hAo7x9BuKyfiJFZQGJvULEtGO1xkxGbChvAC5sceLG1764goS1MwA8I5SYRUf
DyJblYcXVIUsRdkSlM+LqRmXvRBpKQQv5CyMEDqHkpW/xh1EXqQh4aV32O35EAk6
LX33GjZfB7j77IVxOQ5hYurH+IgZYXZuVHbFtckVl8zCfEmPw2F7wYwv5asDplvC
+6JfM6CsDkhoWHVNyTTfPQ9FtMR/XFjVwUlPicha7RlNw15yUpTGy197y46KFJR+
I/8ASII0BLmPC57d18kHou2ZkBN2RXF249HQoQ0dfGt9nSoL+uZUhyXFXarCl85h
Alj86HiZDbJuvM9lXEm0imF6oXIZ3DvnYDyGB98cIUXojgMpzLnm+H4o2uJ6uaHT
Tz1KoPWrFAfNBOkBfmB+eWAzqxiDVxL86uoawfmUUWs9utJSQ9mSzGdF309lMNW+
QfM2V43SSv97G979W+UA7nn0GyGIdHQsqnjz48YbD6Vd5/GKY7OnDz922H+qGAYu
6nXOQdxO21NRqDxBlpmfVR36VH3XgegZ485PU7p4GFtvyNP9njcapRTxCF5YQEkT
hhbz7PnQRc4/Li+DzfshvmCiJKFk0JkcH10QyJm/+qWb/s1ezhk7XKyDm+Zo6GZn
cEkZhKNd+0e3ocneG3mZvRsKok4ueepe8NHrVwx3qz+gxv/Lr06rUgvHU/pHiMNx
+nA4/T6UvFmSWTrPv+ns3JRPxqgbcerf04u7SI8tZxqAYzsWIQSpmXCgBqQO6uTJ
KmIkeawcGuRnmIbJcHQAvnSlhaP3XiwnB0wpy1FEJzEU3qxvpJfRxvb6PkaK1lCF
k/bGJ7tQGlltkOVmAJNW66tHRaQYYl16SocUSMkWyxxwa3cKHWhcxyYsNN8uOq/a
8o6JEujLJb87ENt2mftswiS6s7db4kHYOuKrNRowVG0zw9QJtM8f4FwHHmhedecW
TxpwBxLIqYd7WXvzq6mIwrsPEuxe0fdM4HP8JHK8+DOXJMt0bCrgaW6/c3HRMOpb
hmq+4JaoJIpfqi61/3XQeMtKwSC/RFaKAq4oHaUPGZf3Iiu801c6WPJA3i1F1xoK
5c2UjCpm5Q1WVJ/ba/v2KYjhMmGI7II50sUZ3ixLENZQttxElz4DPHkkAzbK/E7f
mpccYy32mqGcayKKYLQA9wnsmBVfFdL+Vyjg61dwjPXmIsPjyxTNroiMZ53rZG3b
A78bF95iGyRneFnngPR18xd3tnaL7m6UxhvMv5bGEbMw6hSjVAjdNGJtcGTjHwR9
O86VQfw/kLOa7RxlM+L4VGJEcTHA2v4TqaPUB5i+f1y5JJr7mMmJr6hN3XNlxBgv
0LXegnRRybsvPO46YDTfPBLG1p9Qejexrjtx80fy1l9kVYLrL8NB7r0SS5+DOsVZ
21swajuxwIDkIQGkr8EvE510ZCKo8hfnfAGSj8bDBiwUBP+A7WizwWo3TjdFuxEa
BlFEQLg662c/3A8W6/FkoKyq+GcnSgyGTmFpt5odbYcSFjND8S++kyX2wU+Dedk+
TVPp2vCH99tYzeLG0UZDsNBp60ZqhGiucCuMHXkPuQi93zPzpIhQ4XNo85+MIrXd
2JAHHZWRFgM9U20g1ox1q/vJKmTg9gdAH2AJvhvdKfTh/bvP5NhpLMIdahGWspqZ
Jo3MBZTGOizU8g+osJhjy9s2TGV3R34hvZ3tT1lclW6ZlG1Uv0/iQMIutvz6ceM4
XbhW9j7hmPHAGXLnWaBYRuK7zeyh7pD5FvGpE8+Cp1hUBFSG2/GVi9iJRWB994qP
qh8p1tMaLsTHQ8o0Jxfww9SsdK513T8dz5tTSnrzIi0D62g5QCgDs9l+i0kfVlRv
jCNT9YkKlN2oYUAJdvxWst8SonbXGo4RpnM6NVaNdWIrbKtws5YnMxCarisLQXC/
OXYyoYE5vMN9Hn31vkOZqGytAzbLRrSE7QF0audBxcvWoqSN7ot2vKcIfD2JlxtQ
m5Mjsw4DYY7aH2LRVkU7APPG+0JNiT5GrITZIJbZ31um3hXDBVE8Tfuy12SYE9lC
FwmgSnv8EfdleySgmefj6NKpvvR5xMYKonfXksYIlcbqeeKIX8IL75jZDccNOjic
lQmeXFR75rFN7HLlIpwaT3PYHnsb5YkV9wEGWDxwrEGGWJhg5RBlG4e1KB8fDDpv
2mNeewcK/Afb1v36ScyErwWZMLcqvQzuzjtmTQu5ti04vjyXWpSEZNchWCHDbtvN
Z1vE0I44XsrboM5f3+4+NHGLy0SVzJal5MTj4MGj1bvn+bT9/UzEVdRUQRahujxz
ZEco68LwqotN88I2OyZW4f79/yi4CnUIoUjv/pRcDv5ZZfod77J5enoNEc6BMDPH
lJIZQ3lfNvVt+KUMGTifmz3DYeE0z+DUXuewGMIApthC8GVU+jHBaJx2GWciYqVw
8coq5ZsXlN8SSx5C8VM3Gj5jLrrx1fJCRTQHyzt6TWeBvjjIt/kI3c755fR64Voc
O0bJnUexj14B0FBA0aqTNS14ke+1QyA91+Cqu/W+RS1sTfEdxP6zEucxlY5lxE2B
ZQg82Q3v/Y9CKwo6o863jkPcUDam00X/fRI3yo6nvMATDDrHgLMQIxPiC7ycgf6S
ZtKmJce6AiIGP5FfyXcviTKEAMFrXkgAHDC/gPZLA4CsBs5DwSGw9Sifa2GN76/2
vYMByldKpjZwzH8w8fXCRE+O/ETKDFrIqlvqY/WbNgWYDCupcT+qVk6f4qX0wd1T
bVYVeaRMEKZb9BzO9xy/d7FE646ULoTMeK6KjvT9u6uZ+DMbDJ8/BoLuMU2oq773
PCEr6rAB8tt2s3FroNgMHb0U39H0/aY077DbmZ7GWwgrm3r+ss3bEsB1OaPOKl3S
f3sOf0Xjwx0qC8OBFklsUFJxR8itERjSoGHeqWNx73UkckdazsUTM4wgPuUlEHA4
jAjJ8x8fCT7oHuadzCkR5VuAGUPlW047vHg7FBOhSfd2UiZjiEM0MrlFy8/P7dav
xGW/rI2ux6wDf7uI1no6qx0qeVDMllELk7g+1TuDPeGXbRvKbOJe6huMiCSqj0yD
+QjY5fnnBhdqwT66VfEWymL9/KxVD27fWf0nTQmpfxvU6/WQ8Pv9GTv4f9m8TaZc
05dFnqafIcK4l1K23gWzIWjgisUxGf4/ETVo5s7MayVTKSwTbaxP/kB8+Us9Q4uq
aptKPtLCd9vu/EkM1HsM0AtBcq4wGNETShorJN18W8Ms11292LBl4WYNiMdJfVmJ
K++KZ8iUWT60/+rtncpzRTb4uB75+rVHy4JhBNmaMGZJXauiMcJgcI5trWe1KaJJ
DTX/G1+vPaguCfbyrgnrOx9yBYYXRdEGG6Z64+w+P+IDabib7Yalv3MANq/mDiZs
UDLQsqOcUQ6AJnsnaJUNfwVLYwTPm6ZQwQr+jo1i+UvypL+qiDwY5+9T+q8ZrH4R
AdGXY+XZ9372DG56+Kvkrz1aqwnTEd0Le6IxTQWTpGoGJohftbTg2UvPQAQFNg4y
sgYfgJKTBJy1D2sKST9BbBFTsJAS2wbyfCltfbvHk2ZCElpD64BDQuJXCKkhoi+T
Gs24XdPkSE/KDMxobtV2FyJLFK2WlH56oaUhp+GlOwPfYD1aRSrqINjWkPxOkdc9
qeRSHVnxA/ZLhE6fWe5l2Eg21bLu2AafMMUly8tG+LEjcybzGbdghaiTppgMuEat
Zo9YLkh+3iNc5txwkOmHqgsO8zMtdPPtGjHcsYXWjhGnirGyd++zyNpkTtNY5OW6
trvL92f1IDq2XsWtxtahV2rNoz+95FpiCRxnqm1Dbkyh1ke927Xz9P0vBzPezKmg
YhIYp5yWR15Qp3VhfPJ0w2xB64mH0bAIvMJmX3Y/sBuLEIW3vC2vI+cJcgMjf9Dh
eLC7GrNqDTiMF/CZTc1XoAfdI5jk60SaA07cvrElo3KZNhRDTcgTYEMJws1g1s5D
S5A0QmCD3RZbNb4WVmyXPOs8fFziR3pj8Yj6Z1ipaaRY8c3868YwUFrNg5/Y3d8B
2KJBdqnl3dmDmhMwnr0l6/GuKZJpF4MtdDXJz8JYlvfrnw/+j47SBCC7rdLEx0yo
yoZqgCiUESJxQ2dnnPXewUpEkHZKG/QtBlIEzXzU/vbmcWMwkaimLp54yMbut2fB
CBLaCQalBexmu/lJUisvvX9m4/iSTID+TrcA7NnhFwgvOR98hlIUTutfEzd0VaoT
5L4ybvMwwLRUvi0A2HYvrtLhfb7xdLc9LiDdzMm+EyWsoi/s4AxmMJUP03xY0s71
yntRWL/LqXOi7HSL6N9kK3uC0pQU7QWxKUArmIw9LVYKWwswFgnNsFbaowqVeg84
42fplMRydJA74Mh5G8SpAyK6sihmOcwE6yoZ3qHUgiLkMtlqISj4s3Jvh7xil2v/
3t8lru+VGiKYAX+7YlUdChhoG/9KG72qeRDXlGAKjQ9+AwjQfyttaemg072fh5zH
KAe9f1czZlK1zx0kW53/lMbIH1xkQLIZ1gANOAkfcC2Nj5PIeC9iY0BB3WJu1zHn
YMC2pOIzvIaOxZ4yisd2iVZ4iGS2BO5LoHVcMXYizICVkYXpuIdkq2ZffIiCmpyz
oIa+jPup1W1EIGnv53noWdtxwqH9SlNMQjtgxU9k58n6yj87AoIhGJz68SQrF2C3
SZwnUjb0DnUArwc+UexCXnrqco9NEjhpHHUySvMk9zBiPPcpVtXngcFDuEpqw+WP
nHTGnFbnFEJgV/co/9O3M+fn8JOgMKNhFLeQWNUIkRL5gQDcNkGaaH1xlbVDiNQe
uUimKAWguyILRoLhEsYVJ4UKiN/ZFLD2t8zaPUCGhU9qf062LzzvxIsaY0+ODcIX
OH8iM9njXdTlzyfSz0kDFeAw2r6klqwnrABrKDvhA1t37EQ861dNG7T7aYKWRBEK
ays5Dc37LiMkfe1NdyYd98Z2kaESLY+WAOH8nSD/fRkVoahLdBHeYAf1jcRYbPPE
+vL+vFQnK2NpTvNM+eBQQTrT+PLOZT/9cp58ABl7yG6e66Cp9u+cwG2sHLJdduK+
eJTq5dQdfR/H9aiin/JxbTNXBY7HDnELBXElVZdZjGGI4uxdC75Cg3MzYtxeeker
hC26zWKhTGeKXZLh9e61Szlvh9BETSdV5z8tR+FJ9Xd48JzC3ktUlBNSDuXwrg7N
ubp+SY+MIrtazMyDkcZ+wXQEiS1LTIIhI1AVnOX6P6rgNKEu3F4yzXIOXJnlrnEH
oU86uDtd0fTFDPRcBbHekiaIewyU/AGYQ0WWN2NdcL3OkKimm/LSUKuR4c9GkEie
NrqoZs6RpMC1Q7GTozJvezNixqFND9M4P0rbWsm6Cx0RoDSlbGJG0h/KnA2lNBo9
m1YluZl7ZBoBl7V+fDyP/QEo0Scwvzq9RV1PyzxRdBIfNgyOJ0btUtzy4Cnm6Y1z
0lkayRTrZb48kAKcuVt45ZWcmwVrkFop8auzivzPAOlSFZzXj0DpqUxgXBwrVfHy
5eUhR+vPNfN4sBQQkEwIe+JQxKdUFlYMe46uBaGGcLeYFlCnehAGRUC48aIQ3mfJ
6XJm6JMGv2dFDwLjEwgsF/3qLToDgolfD6yIk9q1tNdMTkkb5RppDNp7Zuvg/MDH
xKUgcGgQMfQlWsTgL/B8xmnA62atqzEvWqSD+M1K0s820JG7uH2ks9jxBptDvInI
58btNqQ7xXKyLdoxTpU4g5B0TMahX5sKGsKMxVGSL2U1mnh1T3xGKgB5wldwu4l+
2+vebUcvWF1g3gYhZotH5jiv5BH0C3/X5uru+C+qzRcJgZ+99m0Kfq3Hf/D87LA9
ca98zK+yp0lMQpV5dRs5XoQ4KnvBifWEpErO+9gRjW285oYN31aeJt8wVS4HYpY/
yiPNlFiXGehkKQlVRzSs/2fyQAGMwISYcdgH2KeqNTpoiqIFD8WBHTDjODvBsaaF
giT1CbGKxx6sMgqQ4d95dTbGD6hx/JeWCXpprl2bSoToOGuiyNvGH6yiMg0ilh6z
Nwjvuswe7qP86Y7AcDKGwy7B2ZL5MAGjE3NPsrWloem28APdpy+hdyDnG6dq4ttu
chHWXj4O1yTH95YPBAROwWQzRwLzNGCQ8hb9DGGmjA0Pq+wKuSu9qdJU+9vKTcub
8vGxjLqHl+JY8eDVWuCY9t+nUaI7o6dNyNOy/FriuVMpnp+rKn7hhMzDs8WQe8V9
tF1hQ5SAG8jJlYyBb0G9pWP8zegOOdNEHun56uFeU6y3wiDpCxtjjos4r7ddj0n9
PQ/FIjLCOMfL3/WfDAausNpC65kSO2b5jzeCF5dEoNaZzczHJqLNm95UPfZn2Hww
rcsZ0S2eWyDeW5lWuDIZYaEuALMU/cN9/8xWnNbZVIwWNi/0LvoWFfgjmGkfKwBA
oHlGFxBolWHJjhByCuf+cl5+K0HOOCyo271G7lvhmF+mDxdjDnRme7dxDQXrcING
U5bElEgZMdFKWNJnFCapqdG2uQi2KqpNMOAsridJaEeEaAQ4yw3qmar74pozkGXW
je9TdXuxwsCYmEd5045f9d3mz9u/fZSQGk2jiCOmghBlFX9U02XVqz/cCzOZCtd4
VAf+8BdqMe0XxQgFWgXy9GG9t3kZSSn2iW4avo/eTV0sxB+00X+IoB4XZeTnud5g
4brbxdp1uIdPUCwjWjfp0tyT7WdD58ZLPWvtGQEWye0Hg3ArwSCylPxeLHSxBxfF
5cf2b40k3y1davx0eBZJy3FW3OnD6c6wrp9QqHTU+ecfn7apu8dhiMec7xIl38FK
9HjkyHsdVwJAejAIyPIvHMFTABVDKOZaTEgJhu5zbapODnnIBQomkMV33mO1U3Mm
U4cU1/9RJM9m96VAVMJgasWG/nuqBsetwoS1iX/RXPtaz3Iw8l6sfbfPcWcs5Kzz
NOcV/sZnWmOnEmx9kV8tObJqMi+7zAIpzCLipSnLPk4sCEhxhjFw9sHsxMqvhoOG
kyWWzu79RCwgaKJY/TWem/mVeEeAqqAQTni6V8/p/7Phe0jVe7jmo2bfxXNHh+cQ
1gnZmDXeyhOuntDsBKw8XuZIjU4TfRHmz5xUQKyu1Mb1j/jrTUKqQd70v2messan
TlLJeF7V3++1P7+YCBGHw9Te+NO6kgZbgr4WfzH+RjntaO7mk2Q6uMeUgmZxps3O
mX25OEA8c6D0OuCILO2Ue8XoyNZGQpTWUp+qVHmRvFgh7JQNOfzzTFpkyTsxrval
SEWWFkQP/XCgN9brFm6tTYOnyEYNQ14fXIs2lN4p/Sk+AG3U4yRkmj0Ma6R1vYEQ
B4q90FxGEsuWE+449SslwKAu+2Sncby9VSk81HWzqnlHXpJg+dTpZf5Vfz+WdsJ8
kaEsJ84xfBEW3Xvo0J0tcErlIAwf+VQTSsSZB8HQwkMnxJ5yCL1Z2CnB3V0TfbIk
NPuzgfcYGoRZPF2IpuabjiiIq8U96TJxESvO4SjTlwOK5sbmBXBMuzRDAQJJufpF
C+SzgyGDeIkgFpkBllTeRfo8ple6zauGVeMlUER6kZRcWTqTHWlo6si1/PffzYyz
+pyr0iRsJf+nHMtfGviEe8vyXmrS0jJzhJImE0ToijoIiycqSGYB3+UhJ5umu4D5
XD3SUrfolLDHGHQL8iCgV2nVS6V5mt7zsAy122CF3hBPfzf66QNltWa9hOCEgPoE
r+kdGBeHYuymAQQDbWe4WDOjlwaefk8CM57NqoV5l3nKe4us6gqrUz5tboBsVWFf
rUHDx01GUwO2hh5KnggMuo2vo91nO6YrT2zUJ0S14e3po+Tbo9YDLkYvJUsFlBxX
3hqs0Kmd6LO2gI20kZD2Q0IGGbjXSTXJWwxrD78ZINaQsXR5TmQHzrojHdUZNvan
S7Mtan8BLeK6E4Nz+LGusZg7/kcuKGJFPVMOsE2xnzO3CBLPVZ/ISw0lhcqE0pTJ
LxmyU64UlNzoAQiV5IeMUoGSwuHglLPULXhy5z9Y8ALP7uXlddk/Ouaky9/UWMlk
sgeNQM0mMbl/0kgknC/yNnmMs9iSsswNOqor+YiSrz9Y6TpCeTrdSZw4d86K25+A
6ksOYtCMd7tn2ozBOtzZdkg4jNgjGOOjchQHFaynlZgF4shlP68wJFYxVPB4E57F
dF+XUaV7YoxCORJQS1sewSs9N+Qn5FEjxi088ooLPozR3AQ/K6hmBM9nz3/Zd6V7
fdEwjRGu+Su7+ky/yi+Sus2uYY2+xn3ahTeDt2MPPxiGfgawe1c3CNCY/DgjJ8md
Mr0VFofCRJE+aAIoZrtFjxOB4jSYxLOTf1aQ9CzEUMx7jPHcKxMmqTW3slcGCQPb
2FZPpX8gaRgh/A4K2bGXTyKXvQ4x9HnLa+paPZX4MXwtpYHWJk6g8p2Qg73wkdZj
bKqwlQxnuu5YaDYenjGQeZwEkoRYwMdWrbA3TllQNL94SBPR/s1AHU2B0DzZuPa8
DjfoTfDyKp08WfeHsDqZX7TzknsEIcYWhBx7qMFh+dGbbBXBgcFbS4LIFJJqJJ7R
AdSOTnaY/LBxkfE5rwJ9uT/pBOhZvoT5c6KQ5SpNHVyNMkRfbAEdATphLovyr7vZ
q1lrm1i4wEvIi7nMfQmWXA4LpXSnxEhHjvTRMwh/Yij5sh4hd1gYdRE4ui8mdMRC
ttqO8dPslCGMyXW2eGMvJA1TEkl+CI74WvEscUPWR9RG5O6xgjbABLgIqVTahcww
GngBixxP4jOhbMH6IoH3Jk5wI2D0xKNZwOYJ5WK4tsk/ucQo6AUFGfw9t6N1lynQ
KW1VgrIewFnrRIayAhy+7U0Sqe1g7dn4i4gmw7P/L9Vca+WIazpj4IkR4pXHMRGL
205/80/AXdljEjwIcqUgQD5AVLh4qgJOzKbcFB4H7HsphqNdjmXPq3A32ymHoV2Y
0Zp8Mje4rDvoGLAdcVHCwXOhyGeQgNideSw7ZLo5gQYcSqIEwFAfV6r9VC+qxek/
Tw8+S69ZRpEwlAK+miO4hQ0supV2sCBuEnFipZRMkiq2vL+0EGPe0Ar9C8/R3u7Q
vF1G/PQxvRDyRrcOVnIecJrz0HtJv1W04pqmUXdCwxjXdCt6lWLu+uCc2nt9G+9M
Y1+YGwxPOn1sQatHltZ21ah08MpS93ZHdSMMJKOLFwUYKJHeYNSnLh6lBZyBYOCD
tUZz+jYMOr1lyeJLZvocsmbe2uVwKYAr+DePy0YNi7GAdoAwAmARO30D30KjrIBq
/r2vZ3RnOcq++J85gyqhUFG+P20eFuJevD/xNJ+ZyTiqNhrRbYiJgkyaMDVWYHkd
lssmaxsKFyGA23VOpJHcmBsV/CjVzoslFG52TLbA/JwqUScoscM1j+ujvDwso4GD
6mYIA9jGbLW0Yye9YqwrWbfsRodHkEnb6xWApUzw5wv2cvTIKM+g8CNNrbwNRhXl
ScUHAWLnpJs2Gs0fJvw3k6Jv+y/TW2sfrPV/awHVwpSp0rs6wsLcgECpeuI0WWVs
RXE8uqCIt2ohuG7zovWPJ81qP1B2OmVGx3BohrKMHXU6NkM0NvYVFaTWlMMrtfzk
xfbcdGyDmlDyOZkMsk6c86o11RAmnVvIgKQWZZk17b9iX8h6nFpigjN0ArYtM4l5
qJJksp2NgmuKrjbEV3ssw9bqyFwjxx0iWGT0f78JTiG+W2lSB+tb3uIH/DRZR4bg
cQF6ygU7M3JE8x1/Ew85r6YRyWcyTqjOCF17/OuiKfwebMxqcC3sjVCs/rD0jTeX
DcmDFtjWzVADps2GmgkKBsmMeDZptyNWJDPBNcNdX5AdsIqUo6R6HlOTKK8veWe3
WgyKO82klR6o+YlAxmdfedCZADkXM30nXRxszo8eIQYCBQvFhuRSZI+wOZPbQciL
MNTQEti65ASVHnyoBEF30xAi3qnNchgU7mGQh7+DMy3E3X5bjL15trrv0AJzeodo
Zpooapv6DVrzWnvxwE3piiEHTXTlU76hIiWAPQYoUTP4UEBcXH6PZb/VcKIl/2YP
gj00cmLj5TT0BOmVScfqzoybIhc5X9pcIhAt5z/N/belSQY6oJTaqT1rIpEoMWgn
d8HUp0WkCqCBnc3AwvAOhnaNciyOt0bIJ9dSDK67G+wYM/Z4F64xkHFIYDoc+qbg
7STKPfsrl/ezviQeELjrbIvvWPed+NQMEklH8rcum+EDs6BhWGJRnmPYxnFAjwOg
ukFh4YRsLh8T6xY6rSuSCHcKW+XDjw6L2q748DHGw+O/jvau9cSiB3x3JEPHt/kh
vfE7W+ot1+75Vh9KY2mDKL6eLNDmUaEUaEtLqUXgeumuDgY9xTWuUGaoW2M8J13H
GWjxL2YpFaulvWgOIOA5YVNamgSEhbJSVV7FzpBkzjyVQq1ees6qtmL89zx49c0x
/bMxo52eRJ1VqXXPt9aCJB/V3H2Hqccwg1zK4stubFtT++YKuQBb8G6oVRaBcznz
16fSXBkSr0UA+gzTIU2rQw+IDukG0XepCyCefiKyfDRl59Z6aY4PjkNc/FcC6cr2
Um9Fm0LwvwRujBRMzXgfL5Lnl5UZhcP9qNo3m4bPqPz+PQ17x3wRav/IfY7uSRUl
MGIGtn5Hru+JE67dkEz6wsgyCtN0HJFsZW1JSkdVq3zOMKaTy/5XqQp3b6KxRk7R
PzZKm+fvK1/wbQ7Qi2qJmxI/0xKT4W+c1+KAi+IffKBsOhtTY8P8ELk3YZ4R1xoM
5gCPWIBmjc2IC0EAGBlgC38iiGMmZ3NqwJSjhCHmdE9HNdK9JQ3XjfsLY69s2ynT
K2Rw2kT3uASUQBaSgaH2lgLZC7z97l8D2hkJzEK3kCxkh2peJlsCZsRBn7Ij1TJZ
cmb3+evFzY/CY82D2vF37nxa1/Fp2S3m6yehvMN11z1VRBT0AH2QqqeBRXZeoyRH
FopYl3lRPWt8FVkEbMeQXOF+JDrb2E6TZhyKfcsHWI4S2/LXHetT21N3ti4JXWFN
edCFiV3g5sYlJlGvTNPM3K91yB7zDm1rzmIjHUnKOUN5/sUl6jIEXkO7vSwFkadz
17pLij8T7x3nbOyOEt/+jrEvx8TVAaVqJItzO56hgqABKbdJGJpzrFnsEmmlsva9
v7FARF14Pf2jyniqqGsGN/QARCvVs58oKDv7lMYjlkchNt8gThbrSQYYXHcfz3Dk
5AbIuKc+3DQggancw0lfcDq+4Ct/K3kb3idfPmA5OMh/gtD5Vg8MSEQxEkDTldsF
ScrWoJizOIGrEdPs5rj/WSs4l3YnBqExvBl43HqBXjfenIcvGcQyHCnue0dwEiAb
jKhiaXXdyKA4pkpwOUihvtnSw4W3Ad/tkjirzO9IHI9FWIh8Ddr1vOX08L6aPFMq
zviEc/6nI6m172qK8K7Le+k1huwySKq6EzYonvBQk/Xyj7z7wx0fB/YOsa3eR+Tk
V3r4SXvL8bfV6jZsiqVhqQYiTwakQfqhrdqLzjtpdSUbhjhUP5SZDYkdsqZAuYan
MQQfU8ql6xdQCGa/0OgZgk3rd69NInwYzXpsOFB+xKs4ertI25TbPK4jBNi0jBkD
08K0Vmi3/hrh1Kq3ruyZ5Fbvp79xgHffVgNVF1OaI1kIhYWLoSvJIXUl2zspCT02
iIqwCeOSP5HVr7sDKHAzS1ruBPZji77VuVC5LAV9Jrd0pHFI8FJaUMdsSPqkUKtB
QnXuxNKbocvnFWAc8q34/tf5pSmQWkINpknUJsbGtoOWCHvptpF52H+oBN8Di5gZ
zvg+7GmGFprLYkVfWwA075oSo+7MlsvXfa33MQ/9/oqrsJvpMk6l1Gp6HkZbYr0J
ATwl9Q3MpQzmLVigD16jJ/08NxeOj3XjchOCJvFal4GynQxecK52oywdeDwU7g/o
T74qeigsr1vCQ7BH19OdNpuVrmAf1o1iSP2vTcYEsVg+Gt38WQKH9gIzqD4tAhH3
EdfkjW+fXYqCa+6W8eMrO76ndvr2FRQR02OmhyQw8TB9F0Kd8zdMkJCFb1WRU9XM
K+zwBCR71t7g0nLKuzLEtEg+UFpwJQvuBMmA7BR+emSnYEquU0zSUEVAAgHQOF+l
YK86g/V8jrN40aL5sPf+zCZO55bHuDQvBucWylYyZA1ywlkM+ys9EwSco3F5sRr2
Zr27zflY18oLiaDuEhkRAoNni3VOkDA+2cOhV1tyA5kdQ4hftNurQeoNfMvHhWeM
N7JMPmbqWzr/Cepv47HwOuhXKuKqxcvzuTDJ6VOHk7u3F+nXNP3bz8g3qlzTGFMJ
mP0oYZXMTm5lS5GhPKLAi6Pei6CNz5c5UwJaJEyAnWs2QGeROfzVLWDYmXNRE3uN
/V/vGB7kpzJa15+O7kZT6kPnr7mXZI0fTT94TyOO1Fne/mehuI3wMSaeR3evOZGy
4B5wctvOveYo3wfExelHXXIm2Sf8/S0JbEUuq1Kd6MD1L6vz/RAahBtZtO7bVoIM
J0p2KdrLee2GB3gKIcyZfO1bvWfiGmC/k9rcOoSsGLlPLndlMuLf2RXKOlqYPnYi
7INOyNIlwlhkThHIbsHfQLRjyFa3RU2WyZChb42ZLZjfCcViLxIp4JVBH8q39Whg
7Xb5/ifnkBLgfViRG8iWLNUOfJSGPBwUsplEhqgveMMAsx+Vb75Lb1Q7SoOn8ODR
QxsU3gYY8Ka0m64SfUG/1W8zhRLAuQ7lbrXmDlEDijCjqrkN4K0n53ObVCbGNAhy
Z7y/DtRXSnsCA6XfoepTtt+8HlSy61Jm3Cv8oCyqO9tWN9wdXFkrhPkUbbATzsz9
+uAt0P+aqmmq39dhNYI9jH+NrMBq6JBUe/vznWXDBum+/gHgH6fClL2et8UnWWqt
swg0EfKAeA9Ze/5xQyoPdIsCkOZwzT4JKWB9/KRyzRnV20RlDNIEBOeeweSdFvAF
8NJHGiWUR1L7OlSD1QyK0PHI5sKhK31vIhUTrc6bfhaF1VLv7KynpKFZVi3XDrQe
GN2pFOR0x7ykyuOOcoA0mrrSlfQjEBZRNHgavwPHNI6voA4zlCeDHjFGUPNUp0G0
agIL/iIxQdWpiaOtfxDEpHcBGjt8MxcflWEcjxwE1a8WX+pR9WTqsf4844kNFfgD
BbrNYq0yn2u/Z+vEp4ikVnk9Zj/k36s8Bv9veEMXKefic0DncHGLFHAv4Ts9Ix8v
UMHhsFuhkZG09sQhVAnTNAdYBCuVuOUwHFnXXaCkPBbywDmq8yr1J3tFql5J4jzD
IgtfP68Hr8p8DvJZQ8Yl6tWfTTn/3CXv2D8sN4MEn2c9OIclbQ6k2ZKN1I4tmM5w
/sspdHJ1QaFbsNwCD6SCUWbvx3iet17qtqn4UEMEQ4m8Tb37B1cPU+eHIxvRoW4r
ojBr/7CwmBsNItvIh8YfSmJHWsy4jVzu3reJxsEaCusDFfW7uLAre8dF5dbnhGnz
xeUzYdA6uUTx+gZzjyeJI/HYiPV/Mv3pwQ7xh9OgrAOskRgeJ1Tiqm31osM3awt/
QTWSxpB5ogeRXtRvmLVhiYSUUDvbUjRnpTmw2bvADKEhVYWZLNKPTonOTOBPZLbF
rLtPer7pBKmxM7hCbS0KU/UnXy6OKhokSS/d36yAPa0pzbs9GGzcfXXLpaI5qSwy
lO3yIeiLcojuF8QPqd5Xvo8oV17lGbrRAthVi28TmK9hBQ2Sxg3GP0NnR40EuuMA
RtnU05mbyoMzRHiqgW9K0g2xvwUE20tSPSTgosAiMMEeXokNU53yIXZf5CLV8RRb
rdRu7HBQuYjqn69J+VKmS3cnKtsK6f/9uv5NKANZpVHu9JhBSvYFsD58swXoIRM/
Eqq9B73JzBomI/7eMHQ+wI/z4jBbLiB6wC42JaG5LIj4WkX96UmTtvnWg0mZkbmC
Oad18A1xRcMPbQiyCRGaGv1SG7v2gE0h/J+meGiozJqyBXIeMFrrPw8lTIdbYbnW
WPcOeBjMw71Yj6+7M7M6sEmBhy5v5hZVqjH4/VKUQI1NUcTEThaDddSfoaNQPOje
l3MrzT41axTRA5Zu76IQiHuwXIwNA7z5+Am7zMqF2dc0MMo+39BcjqyjBHs/pOzU
7rk3pW9tr90aImWGYIse/UCqD33gZ5XBNUlja/qKGboGRQAVmt/TL1hpuBrnqRjc
1wqZjuqQd0ZaC5R2MiujpIbMelKCrAeer6U+3NldpQKvu2G8MLNfISP3ylz4zqS/
AzlALSPwi4l2PpgjPoFqr7s1xX5NH+96TrKRoTNyvZ7+KhazQW/vzHYJ10LJz2as
59BLsQ2m1104Dk0K4KnFanHkRAJvEcPuwxOl6lthtlfOQ9mIwWZ/EImgmHDH9SHq
TAdkSNJ/9DZtMybdekg0+lpRTejHaJHu2szeqgJ17YqZaLiHODbiiJ47Z3xVvGim
nh6tIQ7qXbzgOsYPusbySEbopnYPZMbKk0fsAUKWHL11uKWBtchg0xnh6z2ute+g
zaf0TdA0n/ZZwTe/rf4i6F7+ajRVMk8vnUj50u/YC0SPZoIDVYBBQ91NIK/LkMUU
lvi8jZOnOYuy7b7iVCK10wUR/LCfotILEcShpib3+kiEiyX7eyQS2mR313/HwT7G
pHAswAC+gkCRrWE5Bu4EX64VauFSqvXMk5X4A5zgoJmCva/KKuXGsaHF7Uo6blLs
EI0Y2pvc7rXLZHpKjH8bt3sr2WLZq0BWPTn3vrVhNDCSXcg6LBE1qGOKnLeXdgEv
spS3A0/2o/ne9sJWKag1m+KzWa+HQ3uvAsq9pTQxoekLdKGG2uZTaIdPF+oFq466
`protect END_PROTECTED
