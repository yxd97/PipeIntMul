`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PhCI50l/qbFUoVHwhD2uJMsrsECNv9AkDvMJGbi9t3BIl+ZvrL4zfRnMxLLwkUAb
UT5IowzeSIx7GlKhly2QBLg8lv3WO9JA/FN32BQP0seU9wOfAQJ/qDB5KKJtf53P
Eju1kXepGocM1fiHoosBRwE5JW0ihbQtcaNMo/+pSFyxFrRApr+0XPUDDdSPVLAU
bXkjkMxXR0FdRa7YFrJHzkfeu3Liwj9sVWmSVSa+Q29z0z3z0GdJqXXZNMBZkNwb
RbJWNPW/kxQOGrEuaAQhi+1CmLqF60YKwP9SeIuda4IhwHiw6neaZzY6eD6dXt58
mS6N+Q1ATHONNIg1QNRqtPocqnnBqOkhpblhZnNkbpvukHixxb7aptv80bXphSJp
7taUxTDczugf26Tj+CQOonKb6+R8m76fqT/Y/kCKHBUiNklT3ASPdJMCg95G1+Km
W+Fxad3TXSsZFdLXLfgbOgwVa/mqYHI+jlYUYZHRaJqRQ5Oe5YhcnvHEX3jCg1HT
ZsgGfRq2SLcImkHtT02YDML6hRP+Mg4VqlHg2ANXggWoT99fLTDk5sTvfJaB9iGF
OcGZY5EyCuhaUUalv0t7g4e6HcilL0FWoLZ1BevFvIEQnGXcCCNMa8u6MDtKWOfl
EmYnNbj0QIep9ncP47boD+RK/NU/LPzmpcgRFrdOuQHgkrK9C/ob746sYmTno/v0
2IG+UhhqMyFN8UiPQPRQKps2iC5A2/wIYClBo8NmnlVfZmMBT+pdVLDrU7R4a6yp
NC9O66ARGRH09XyER3U1rE4hI8E4IgQeg7HEMit0MVKpO/lYio5u9E4C8oJUrGFt
Pyht+gAEaPTsE3VK5klV1pMqqae6S96Vn8Euk0jPFN3mKfPZkRTHyVgvP3b8PRYY
etBN+nO9KAFo+i8lZzZ0WEg6DXIAkWziIwKEZLOFjquhEBYr+M5dowfo5XZKca76
1AdKwnja8jcj/Si9GZj5FWEU6IW1Ffib0OE0RFoXvpc/Qs1fA+qZE+I9xhm13b6T
g8ePLioWVY9r+HIUTvOOn0I4pusN3l1SQgduKP5/aFHaYfcny4Y8z1YenPEvRxYI
OrGMTzc+ECeK+qoTiZB9rg==
`protect END_PROTECTED
