`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xUAsSznu3yjOI4N2pEqehs2TfOYunapaP96Ou48YCp7vkNgA2AIjA87UpDH+mKL
jJg6+5CTta5DkN91Ues57myHBesMTvojzgtfti9lZ+tAd1hmxr030WNkWQvUyOmM
so77uwc7/sgpORumiRiu7C40B9ZOoj8WAVxHRhLoAnbQUA7pzljZ8MTEpQsv30Cw
hBpLR/gRtRWEYKltknxDbEXS8uxhB7IBACgR8RYOv1yVlAZBMnY129hzzzNnkz3v
qIx4vVXzhWzwxA4H0JkepQ9f2my3K4DcbReJ9149PTwkRizff1p5UsXGrRui/pnz
Ta/eNabvkj6erEjtvtQPCvEwlul05MG114JrnGBnB1412zgFb8G88Q2R7bmtxnIq
a01rfw4Z5pJu3ANYvHc7tOH6XznSKsLKYOJ7umVEldtCwZPOZKxfOagiTirkVhh9
DiBFCu9NUF30dHvBJeeUnS2aGPvCPCxdDCGxWY9hCebkkY65ymYrwMIekHuYtx8Q
b8m7td5lGX2i4OuuVRv5+Dy6sVX0Pdov9lskaE9QAbzCxETPpAyBpYRAN4JB5xYE
HUy9XwAKV0REiumyKZZj76oH18aPQGD/kEI+gT8SC5gkShXYcMv+n3iJ2Dy5iQja
sKsmOpYn41TjWAD7KMu+t6sfBI27V1KLwuGahwtcQYFnaHkMbkwcZ3bKWzVnY22U
n+3HlR7yoxHO5ExsGi5fbQ==
`protect END_PROTECTED
