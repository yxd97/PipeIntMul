`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2QXkc3u0h/hMCgNcJsisy5SaBVD7/iFOLiRUfoDkze8mN6/mDWRwolMekPa9ZFiJ
zm0J7NelZUxuOKZfvdZ7f+xPy2zSs27NDRmQOmPMwcAuOtYi3kbFjQ0pZLDN+bz0
GUTFwJYUpyfZXZbnxILIfCbZablZn6C1AEWzwBu2neTxA79w08JXGzb88VUBkfQE
pimOO1TFgq9EMs3Y9PQRJLxthl5Z0Mg2uE6skpLsJKjGWPuWwvsddY+NxdsFBByv
KxKV6ROENHgXlDN+aH4+veXQbpVUCQ9oHSStfRFt/bPEAtxI2LFaDv99L7J03qrt
C2cFt/dTzuiAM+3ZFHqj5osgxVURky6GyUqOhtewXodan2mXTW+pJqFSyZGLXQyf
snKv/j5qhroxU1XeurcjBOeF9DJIcwH58vvK9r+ScLNcAf+iu8CskEz034CtdcgV
rP1v1hwpI1AdUq3MmKRulTj6EGweJTmxNDd1vNFKhwq5VprZn9EDS8mmX1M+slYH
`protect END_PROTECTED
