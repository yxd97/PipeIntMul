`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FCR8c3Ae3xEM6/sKrNWzmArmvGAAj9ET2TQX+8ioGuRp1P9iCLaVu1lCcnlp6L5V
wdBgx/fdrnbcuzaY1MAUBx1QAoQX4v6qSq1PP4IikT6XZeRB7IrszuoOlbt8zM6H
HuXTuF+BxvwGuTOoj1ojdUpoZ1+/eOkJsTaO+zE2ePQj9AacocASaF1SpGdcSWPX
jLqZqYbO+B4jdeWkEtrEx984wZ7dFtqfOxKR7Sjp/83OdiWTRgq3LC0lh1sCUrRQ
jfypfttlasuvDB3Dgf+V4SKvzpRwl2Qc4a2liWpJ9pjO/O/eyI475kCtT8304FJT
6KEDW8rc614wR60Oo+PEncCxsCGBB2d1F1oI5Y0Q9col0vHjvVwyoB3ePVVbaIMx
jV27cnNThbhrMJ4NFzasdam/oomu1hwQNW/FOiYZUTg=
`protect END_PROTECTED
