`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thhr8KvNhFpZP/aZ+5VE2afUCPt9IVRzsShlioGz/dUnZTigmRi2RxKPvRhDvwEk
xWXDjmpFVBoJy4S8T0Vw+cKWLosyjj4u/6jKdkn/1eGFQm3kOCIvh3ooGd67idjH
CAX3ai53OCIlJWlicLuPTAVgZhR+iHmuCmMIkcDGI5dFQITptrep2+E8kGBawZym
sBwU/9/huwsPmCQ198nToSQrShL0vdJer+XJK4R4d/se2dujj4M1gg71Dk+GIdsh
J/XIDfVGr+3bNZtB/hc0lyiJkd2efSNOObacA4TujFbN/q+LgBtmAJlCWR6LNq71
olVkfat21Rl36gqfAUDvKCHk88r2gD/Gl3sj0xbZxT/zhopnbwPmpGnOza9cg8g2
YseomfdAWoEDqZ8D98XD7PdZ01jIb9C/Sicg3YQJx/Ba0w83xJaPrN/i9VNYDiSP
nBNFCmdYxhqMNsLr4m9uYFu5AnyPK+2Iw1JabG+neMg0kgIIPorMO/t2oKdi1D55
ksZXTAcZJISbPDzQbO1YlzVzE5BYK/QBpTqy8vThm/OOYmu/dn29fuBh4quQjWvB
JpK1JtjSoor2zreqP3ThTVinpIut1Z3uHuS3PXcnX+fKaFLabl/OwwMalTPCipZF
J3szcF910oMRovSNnsHs0pbrZkYSMBFcdR4ddmmnq4JjyTj3IQvdovAvT37tjtjQ
Cd9cw9JCN7Oe0QC9nMwQJAK+cgGoZF9BQPpOVhXL661I8T3llj3lw9HybO4L3ZA6
1TygHGhgiIGDhWnX+1LfXoSs3NhDxHU3n32bmRPWMXsVvX1ZjeuyMAHwBD4mx7/7
J8xLE0OPl2C15u+vZN4x4I8bI5uzsPjt6lFS887TBa/IGxkAONAScZZKjJe8/IvB
++NkOwFHFotkwb/lduq+nUJ+rhTMxcN4EPZmrBzq7xDzImEA+81Zr1uIyC7HkJ4O
pI/QYn38rcSxt2157cpgSx8hgebKsJJszc1K8E3YjMzY9o1C3Nrazc2aswOeGNXh
aGKI31WZmPLMlWp1m+3Sz8UDwciqbKapokKR0W6z0ZBONeiNPRBHt7PdXrkcLrsv
13+lo/pr8QzgJKbWK6zqIvq9o8Xo3n1gqVHKWdDvjGI5tkeOQeuvW9CZ+HO9VJ6Q
mUTVxfNBnh3BTqOt2gDJ5s5n8WgkW/8kEliI21yu005Ge2yCrWQCfKfXSZBbCZA7
Zl5aPBYYuTVO7LCfzWcHbyCy13aeSFkYPrcqWuU2RzLVmq51Eg0lEUFgRRcp2isE
/LZcARNDvw9PsuB9R1byPhwkCm8KL5xloJ/FLgLlRRoLMiiANWwfDbZINkLVcPCJ
TUyn0wlK5DSpossWCokoxaXeCYvPAqw8/3+0M4+UBYaxCDzQLITCZrL8yuVeQHxR
J/5bQ24G+aFEKqD2L21tMIKCk8vgnZjQt4UUKUxY0Njs/RbZDbAjjxRzbouD91Qz
Dw5cUqd7li9TFC9E5DOrEHNKsJ9QKjVz6Jv4h6PGPmrDIpUN4WUXZ5VZ20sw3Q61
whvTmlpCU7b4xk78jd7lb5S09SZNSYo6HfGa8wZ7wlY5Bg+Ul3UA9aM8m7C3QtIy
`protect END_PROTECTED
