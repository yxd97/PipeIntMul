`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aO+g1G1L9cEJrrty+pB40QkF+P2/lpQg52gW/RT/Zd9EK9SI+S4huDHMYnDpiZL3
Ve0Nuy3If+ahYYiS3uo8DXL1XBbf6SLm9iHF2MZMoE7/zhKrfBcbaB1VrI+Vriy0
CiNZrY73XjzBLVXiPNHUHj7jyYaG+VcpXdE+MTNmdhP4iAgNzwvxT/tQFSx+aeLQ
pt6cSKLgIy79Z7wcoK5wvBbXczRR7R/T1dha7vsQ7kf/aWaOhBPZQ4Uzt4YB19Vj
4zUlrMYf8TaEbakmBgzsSsdiXwsNe3aE75JIT7SxsXex/dgFa8vPS4r3wRcEcjk7
2yRyCb+SKm4e0QuwmBgGGvLYKCh8tIXymCR7HXexAzq8cJgOCQJ4DS4yodyweLGv
u6QO++H6r+PJxtmaKmv2d2nQ3T4Z5Q+QYQItaWolbdGLyzI0kr6GWaTm0XDUQVes
12CbYqUNgBIOet0XHzlYrvall5o9VW8loUnhKyYSYFbjwck2Mf/FL/xQBOMysQBg
Ar3Gxg5o5Sl1wufbS/E371X+YOwm2iieQeWWHo2jz690xOqKZ9jEBg6YFpoedxh4
acwJUhY98J5ILurip8ua2NNCdW38nTYbxMBWfnsV64g=
`protect END_PROTECTED
