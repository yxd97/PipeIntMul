`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZtKXpDBdRPJ0FVuOoMZziYyvyplFDQW9eOWs/6SRFtt928vEtxFyRnJsnFA3iWks
ZLU0zuFpWemC0Dksc/LaVJFEvLurQbP/Dft2E+lelz9zMiRpk1vP2LaBJlOSB9/f
LuoyYJpj5UxAW92QQ3Q6570cE8qOqHR6YwRCk4T8aqL8QQNJjs8CHjOWZWE5MSpx
C65IGQyKNAVHkRj9HcFWjVSNQd0v48t0IBXoWINuNCPthFgMHHkGz6uY3iTp6uIT
QxLLpY1m2WTmUtZPHGO8ivvWNxsmW4IEUyTDWD/B7zRfpjNN7p4HaaZ8ABT2jPvr
ld7m81ybyEQxLZOU/AYR341nrXXhPMz0lbLtqevBVnKHc8VyKWvzFjIN8VZObgn0
ZH3sJ6lN8PSJWkQQ8IeZlMP2sA1nuywPKbNgjifhfDfDtZyGGcWphM/f59mezM1H
t7qqmukm7oc9lT/0dZP4RJ+vkUMcsB87JMEd0iAVOK3ZO/P7UT89nYwSARFxjVPO
nDZpQNeimzLWepU1wvLA9BobYa6XEq/ld6hSLe0gMNY8JWBk0Qyn+bUTxnGBVEqd
lkvbdQyapGVAHBQDFGR8vx3LPUpMiV1BWxEWqJTpn+WMFP4Zba9Gb0SrZrRWJw4C
AWCczRatSutuVC0sB1XFvwFVp8uVe9j/Qf/F89YJC4Wh7FKF5bvyNIP0EuUDKBon
e+L6Ce/OoEB0Ia5IfAZwi4ccgYPwk09TAQblGgsOSt5NoLNWCRDS+R16F+sT8XuO
gJ3pZmoosHsBXxHGr0bpNKk4QqKHIz1wtQGaeinLVYgmCqUw66iZjGXdYWV+OUHG
6DyCRtb93URElDvrstT8O7rPifYGxmIgLKrYptZhkAznPWWClkEUXvwQprEJZWwM
RDNGfwouPZhag4A7OeH2nnERKp5C9fedGeapfmoLA8elY0lmH2MOwyD2TZjnOqGS
7qWTlLwRqofTdY5+SfA4SVoWcsSbdqMcGjAHZLisiSvDc0ZUPRtlR3gWv3EPg1Es
X7pwiHvX6nfloSWlulJuyNSYjxFgVkquxDySi9vuTB04CrhdZNVSBOUQDp8EM9C5
J4AQRCXnwFe1D77/+f3Ct9dvTqeZrNCz1a8rF9bPH2QrvClgQYUKqf/46o3yvTdn
B+46OzYpnJprut5WC0tjVzdsdPffuGoJfmeDNtSUTHz3fsjJ8yNAKmpYQ7V+U95g
+YwQRlZGlXC69eHWQzE1h+2ffePnLxy/wWEh+KrJ5ATXgm8UiiThLeaQYTUtBlkF
/nP520mczY7Bjk0uyH9MXhxqUmxXgkNvtoMxbbcbJp8/DZuZqjeRn4q3qXmIcd75
gp9uUl2GYb0nBPMOJs15odP3QroCXz6ztu0f70dT+UeGwe7MrWvPJbwsKVD3fXTG
xA20ERsLoefprKa34fbaUWj1CkYdCET+nQXPhNezuhjAnh1JdGScR8cv+vCTsaMg
WwSwff15vNYkTsKD74sGyW2NMRLtvXHYRx4HdNgacNaIHIcfC8qRSxDi/GeFZoF6
ir1SuTJZHsagMqNfB8CAUKlpVc7ir4HQAf8qoWExJxw=
`protect END_PROTECTED
