`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wF5iEuRJLx2el8CHiJ60BnkFkOR5k5XbC8XwR2vf97Qet+tqLtWdhKQwEiLa4zd7
8WG8j1gSjOzvOz96rDqZ9Gi3FuaU52r8xbhl6/MKyf+KqkUUNm1e1Ie0QKx7gmUj
DnN/B6D8/+4hn3SWXq5ArFuAXoSvaUIk5YUDqaLjpg2MQSs1FOF624oVW9oIDF1/
nLsSEVXymEHJkt28XhkpLRfxroUEjShT5CHjb742/gP1H0o4h3Ath5a9TQFK/Yuj
smi3I45a+znzvtb59w5z8wmOhmPYbArKlzZ1fQ67yzg83VtIHWH53lVRmsS59HYH
FQ+FQNEQjGFKbgoURkbNprb0DTaTpOPndTAnyr2Mqe/BdutWEAuD07gNeBEVlzhl
vsKv8GIOzRCk92ZSNT8sLG8n4hn9O7rw1Mt27TGwrfhcBnOhnnQg97hm1B4g4zOM
`protect END_PROTECTED
