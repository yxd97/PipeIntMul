`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fGs86UBMD3b6xKq36EPCJHR9qoPixuv1XghW/Tl2S6GnPwjes31yxAzO1bs6MhP9
ZIf74NFFcD5RIKk5dVyQMafB4eWldTjg7UuERsnROeXVSFh/LHQIjK/vO2G4UBJX
BsaWTAo2Ga9kotnv2996WAyUM1LcSyCh8ZgO60NJFABxXfqWYCIJrqMt0tKEKC4I
UQ9TdsdYTLYk7w5/UbOZ5N5PPjijh4kvopzz1p5CGsEKZrxsrtdv8JD1dSX6/kGP
AKRiJLhQvg0MU1xA2ECybgaZn9TMz8mZ8KeGTfEjKoTrL3urNwtL9jclnUJiVnNK
Tgw1/4P9y0PCBiT4YtojeGedH2ZpMRGVFK7RZAFWyRuKbCPzpeNqv/995eWVL8Z7
ErZdYO9DrpYODHLNUFM+GDqBYhRS6WpnjkixiPq4In3Cr0ssaWj2pcBJ7wL2qEJb
uBbKt9hFX+DjC+krcyWSfXyMsXPjGXFnqYYcPOP1PTN6xK9QeDRtlJ3moFyz8KBJ
AmiUTtebl+l2cDAA5kuCtEZ1ny76H1VW/Sd0gnj9wp5pyFpiLk2GtDPIWBA9i55h
NbTFSO8uHlLKQ2ug+uiGUaoMUqfIQqV+fEI0ZehHsy1TjBa+LxxjvnjP3Zy6lc6V
J/JiGWyevQ2ABqxOWHzTVXLj5LJh0weafkEmA0yZW79PAOqMhUwgmjfAEIq2r+8n
EGTmyDYAIWHxmOQi/lzp389l71QkmzpqA5CgAsCZjcvd/FB5c3ZA7K2aVUgJC1cX
VYlvNFflcgYO8u1TpjEcZvO9iBwGKdLGEM6/kYlIVP3UWFHrTLajAXmGDOV4v6tP
ECfFI5Bjs7hodW5VtH1yfxTVYGARRCsh9Ru2Czh4rNQ406Bnepya1NA2BcFAeNEb
eZV3QaJWO5uNsDom+dlHRKfK5JE0l25CLcJ9L2qIdA3nClHIL/QmR6e8nh9hb4nF
`protect END_PROTECTED
