`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GA87j/oed/LrmqoqjcnNdtLZm+cVzXZ6DQYeJe4VRkm8t5pgGf+8IpynB4St+xy8
Th3S1BSc4kFcUU83ocg+fe/Bu6KKXq+gDJqqBDDKKMjYm5y4+vdnKo8qi8v5kEOc
koOz5YWndv/Cu4cOUEk2Ul/02EAf14qu6Ivc2zS9cJvPPef8jliRtygJmkshvFR+
FOvbt0A3t+kn6dePfxLWThQZyr9UVRhKK0lBbJ0ZyU0yJJUzij1IdFd5rFidQzbb
Nbepab1Dr56MANByZSK/I7pqR3AY5BSL4+7v78AdYwSRqY6oHzeKwU0ILqfHNydB
74AiWqzJflQNh7tnJvtGc06s3V31D1NBv1qUzeezOxpa45871afI1EcCAp/BxV9W
EGTd416HGc5YVo5TylQQ6A==
`protect END_PROTECTED
