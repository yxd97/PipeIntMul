`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PfsHGvM+kXpUaSsini5x40RoZllqq2O5mcvrS+3VGiOaRBTKc5tlwe1hwLTTD/s0
6UuVAjM/LCtDQakVVx1KnhpbQE1dEc0q2JhJy52cx+fVENMrbAyA7Hje24crOUpj
3rjKkGbk34MJs4atXtn9Q60okJRFKM3GqJBdcA31N3rljb4+5hI5qPpXSOOZiKhF
TNuQd6eLlbS7t4IQ+nXsT1YXDQgLQrpXOOGJORdrpn8NVtxxMglCIZzEguhfasyE
hxkYJHCYv782bX0XHCQqcgHnU/XNlmoS3sJUnehfaKTSNzSmxFNYWy+SVERNPxte
58wRKCJEb3VgPmm3/eAmPbUm+lWexvlitDhPgqdVVh3MihWX1IZONA4cPnYkvCo3
QyWoG4KSrKUSxCf/hzJ3YekRIO/sXnXOESTzKimO4BL3A0dz8CVcy/iTrEmpEv5Z
dKn3i1UhSZCDyyiWnwJyagJ/gnx6GszrxR016aaSsBVqyHoOqjaYrML1wvuhj4bh
xq16Notp9rMRFNEq5MZCBAG6QQA0wSRNlrsGm7g3/lqcId95aMNtAVO9o9N6kyhg
uw1m6ejTMFjb0EuZwlBMS83ZgVC5y9nGRg/IrIGiEJiEIei2WfJzEon1XV8BMY3u
h/t+vKxOpG2LvCWNjYMjqR0a27Sdo4qHN1L80KBYqmr737mxubBbba8qa+NE8WFw
Z6acr6OUprlpPLbfEa2t85+1a/uGaK7iOJt0/H+W9xFBEsGc5U7YUnOiXL9EBLVg
YabFP1oTJ5eko+Zje3QB37hrp/GJxJSqfu3x87OBJTNbpoJqrk46d82MQ2FZEefa
YZlZMtO7ypYeQzsLmiMmKJqbyDKjB5X5N8k+F0ld9+lGazOn9d1N/renXQB0+EwY
uRwSrcaXGRjsem+JnvTrzieYmlL8rw6ah5shJZT1M5eBJ0BXZjXjm51MJZ9JXIlv
6PXgHJtpXB4fPXFDwxnCnharAxfSkM1/vsWfeeOVwi5wu13MXqPZD9xlyN8V/Dgw
AP/38wI2n4aWH0OSe9OQMqmGNiPDoIMq/EGmtxKJ9H1yDS2MMwmPYSTnFcJidbDI
XxC7CoxhKFjQTRBSSS9UQnLktv6dYrZ8y+EHlhnPzGehH6OZ80iTwKgPR7/5fVru
NCQDYYWYfrnitE6vbVdKYIe2WXU28bQySAff2rCFTHE5lUy3xcMP4XLdZ3Ov8b5K
c31kfjTrXF9RjZqasnycWAEWqCr2XLC77xfZdzfMIRXahuOZ/UmYtRbU5BaVN8Br
ujuDgqwaPlpYOUfJdr1O2sT3q4MS7KUuKHLZMMnHZLszcToG4p6bCnxLE3T6nCp4
gyPFw6CKMPkmZ4+Vv4FcAXcItxFtXKOlROTJrMSyYT5L9VpX0OD7wfsYHsOuCxE6
gb/YtfqtIF6D/AfIvJiNV2Io5vJUhbllGm9a9PWR8ujLzy7aggFhfQfCHAQvLDQJ
xt49mwzCN7m5gnk10qf5OUSTjxBN1SfJLB/3JjQYkcRzrfL0JkGyojwom6xQ31NK
4bYo+rkoSCz8o9uQV9helMz1MNchGFvHpLf5jVlNlGauivdHXl+xSc+VBzpnQU0C
unR3FOpFJ+xGffCrUpULGfhN3OVmnAsZKEVwBeTcUQ6za7mTF5J8J2bUXfTnUg0a
tBiYrrZoo/KwLqTiC4cEmVZobORnA5m4pyanRpRsOYMPuLW7Z6Zv81wPmGznFLua
UQ6sGjU66EhX5gBqz0NwTaXyzqK2jgSPzJcnFqlLVXfyfHZB3Ihrj8zED9sCHZ5F
V9pTO+5eDJhqwNNwj/b8HCOijI6UC/DFjjDMvh681PzG5z7tJkQt8FLZ2JDMEMMO
NlI0YWho14KBDS6fw70KiOc4ERbchHVcjnBDXG/vBrs+x1GlYv5Za2292GGzswH7
rhJU5YVejOzmJUW7w7OKxVQsl6I7r/bOtwTsf1GiJkHd6zkNrvgQrIRNot6OgkU7
R71QyOtLRO61rVIQQoELCcLBaSBIk0f0mx/Wxw5OpWJr7krkJnpDefPwWB2AV9zJ
DzdMChONWjO5sqs4JWTuBRIWR7xhlSxU9kbN3XIudie6qj0LK5qF807LgiqnJH7K
IqlFVs8DBsNtzr2yTqR8iYhTYo5IquQU2sPQDK4EHULwgoyw4GFJsrgFbxk2L0L4
bCBqNfpHOGdj3c3PRQIUaVLq0sPeTgVsDig1v8F56OAdD1VuoqcSWdN0MPUHKyGR
PZwRTZzO3KQWzjGgV/Ri7LazpdY7AmWRfLGjDAXpsEzgqIyTM/o+qy+YuiiJDSIv
rogwIWF8FI6p/M5Q2VNnQvBoTPPHYyw6Q2kY3o7aR+kB6y0nhj74j8ZwHbrqeWG6
iK0c4uirVo09NvcvxFWFt3Nrd6tCFKu92HmjXVM471nlwS7mOr1ZwfoxRShOUvBf
RcP7PobHbTaSTBfSbpWx3QGQIChdthnoSsnb1Du0JohVyuBJzmaLUG8bnTeoQ/Cf
2sDKJf+Q5nxkheuITN4z8en+a04Csnkujer55Hh/Uce8J6lIQI8UQ14piuhgbPHG
uJGCN9r4Oai/Qbdxb9OzGfQ4smDgR0mgK4qYVHhl0eyzANx2qQS+K0NFXgCego0i
o9Q4j0L2Ae0EUiJoVk6LxiLqk25ZH4V4JUujVVJP+a10Nzg71iMBN60oFbHszVxr
Cf3xozQKJfMKL795dWj9R3zFaa3e8uulhE8xFJ+89KrxWcDL61VvaBMwTh/UlwQt
7jRjU8W2cqJQRlUnaeuVPSvEZxHdTuQnuvubNHkeJV+keHEKtDmEvryq+el3etAs
SBsD3yhQKAAO7Rx4QcIvCYOXImqhCR0KASxREnxvlwJFMnifuWlHP6rGYAt//5GX
nMT9omlHMRK5TiKU+L+Ddd7J7VuFKSMP4iwuBsgocBUTGh7Np2oGuZB0wrAwmXOp
Ssh6M+uH7KoQw3olZ7JJpjwyoiPp18t/Lr6R/iUKJ1H4BWBZXtObYZtDW489VWXb
ipMA6Mu9C3a7tBIw3QrNLD/UxOgkxnYE6ODnVQn0H6yuaz4pWWfRHv7hkV7lPk/o
BhCVDZEKtq3T9qWhTj1SW9+6vn/3DV66DEOv4Vgz6qq/lAWbDR4iSvtJORcjcrUC
ujckieKkt4v/HoT7UUhnxn6utpJ7uNzEbpexqYlkVrJeg6Xhx/MjT+SwN6Y9CQHw
f4UHpCbtDCxWKsTNlwslt0AWQGyWQDpJH/eRg9qC8syGvj8rNEA8x6C9TCnv+10i
C78l2LGhF9x4pm6AxHUvIekcrT0pgQ+j7FmggyNJccTfi4bIpYU0OAP7bA6+LJf7
JsBA6Up5H96GqDgb5nPrqN851VSYbYD93yxPEmvYZ9qHsasMSE8XFlW36GD3obV9
aPjZ18lX/ys0D43wwRaKvYIelRAwGPSlY4YZB/127G6+lId3jTJC/FGkYs5KMvy/
YDEMkLs54pxg5If7SU4NcAQHO16BTJ2u9Z8Km7/BRG769QQSeTrh+OHAmbpXUCDc
c3hNZs2j+tNAxiz3S6crntyZk9MbNsPc2eUO8+yZjOKuhngrvgNeSL6QIEzoa8VN
H6RfJFMJqpAshblMzvr5IU+GQnjQvJPQpSFoRzYQpxqnmmJYT6sGVZV5gp1j3aEb
r3k5XyrpPwOmxTjHtb3A6YCN49tezTCvhn1ersh3hGBnmdOEoSwFLbE788I3KJ0r
ydCKkaItIMshe7eMrip2C/WSfDasNhCEztxz/dn9tae8hmPGNvRzYUgQvdNxLgyt
1QWXZYamC38aKgRk78aGmy01uoZ8XueyctFdIqtbsOv7cyW/pOhz7xIqAZ85roO5
eG5eEAy4DC4ZULw4epCmuNxyM0uDW+/mlg0mWH5wVryW8csfWPPL/9qzMsZoIeDh
GBFnDXT1eHMiqh1fcKSxrX63PeXIAKnIANkkmQNKvYSM+yt3YzwSyWb6yNioSWM5
zQG+4KSiR6m+un4Byo/gzioRWx3gfJ8qayaAD+95pPMeZOgipd8wUdf/etUin+77
A9NBvWcuMBWBR8JvXosfZdBS5nA1+UF3K5J81laS05vb/7Ahf5FtUd6Usp3PS70g
msL8LVZ1l6/YKzTy+O0opAl48wyVU9HeWM7noidTy/IxKgNM0cNONFHOSo9vmP31
OpIsRxjM1SZrHQHGG8J6esKgk4hEJu3WFEbgVVkznwxGO7489BS+1o9S/PFO9c/P
Pofjrer8zbiCWRboFlkKvqvnwQfteP3Yj5v9UZkIhIWYyT0swW1Z6+7TW8SQVE2v
IYsvv2FNSrzA9tBivmj3QiX/P73h/py7zlJ9UPAnyIScnQttnKIOBXFww284K9/7
vETQr/XiqaaxVR/ZWr+w1iEbP/DJQSBfc5ESAMgk5x6+Xes0bH5bs8PBBEMIEWZO
7bUXP18gwaA3xpeJ4ii8SGSr8Iq521A/6WAdVaXjymYiIDH1mhFQnkmUmgtWEFsz
lVNm5jrDkzDDZr0AYM6CKD2ixyHJ2EBSODiI0FNRnNrpnfiDBOaAU9zV42435usb
EBkdAUyi7OXNYOY4g8CTy/kamhUMMWNX/b6Uihh5OT1jNIc2BHOfnc9p2SJdG4Y9
rfIE8iWhca2p8YCHHyY7NpesA/ZEDk/KA2//Dq7iYG0D86dQeuudbPA9NGGjzOek
4rCfcfOrC7BX0PcqI18JR639xYcv34Us+5CvFFGwe0GsE3LEVxNeNy626YUw5asT
m4clPL9/Q4vXue70cYuWI1+t32XduHUf4RZVf/6l0FdodhSSViiq1F5Y+8jSR14N
WwpoVNxObhyQHp3S6VqdtPHeRXL3NPpvEGb684lbhGLn3QW6UAbvgWL2/TUP99AI
YKz35LO3jWHxpcwSH50fpiyxC/CooMvymSJNo6dcHsFWm/JAXR7pFuPw1btbsvla
xNLK79jgGfwVJBL12xvJZMg2wV9R5gH3U4MHt29Y55Z19F5EMQ5A82tuA0jFvwd/
oPLERpIG+w3DUhXDdTvxyU7F43tNtBLUHAgWT0E9VWdxezHaeOqOujT07VdQAnMR
/rma/rO4B+Rihw8Ebxo2exQdTaJImHU6aaXktMMg6hQzrpm0CsHAwsYfGT+3TBHy
HjVtP9ghmcz1DTnoxQRWEjGrwpAaMqeXdJHfFx6khycUQmPRm1SH7Pk4KOUf/u2P
Q/Lcc6J/GXhJmP4nd53gIyA4rWlSVCV0WQOmnHEQFvBgPIgcVwEljkFEL0Pv6Y7t
+FBuvgSSrUysfVxLBd1ynjzkDeYGocLHBMBLg/648954sB9ihCF+4h1LrQKLjme5
Tvc5ScXsIrOedDD9pYTYQWTbfZhi5KzePSgk2T/sSTyASjqS6wmlAq9n8LnaXGpj
z0QPCaTbNFNKXUTgfcR9X9icHxYBTbs7U9Pcats572pcrqYL0YUhA2SdRWdOYTkg
yQTPIvl4y8g+9alX66fG3zjlRtp1V6zjwh61ZMpngNm/jy8p2h5kS1d09WEztcQe
LMSSqKxJxZba5fPq3q9/ElaHRgO79XY1PzT+z0IadLisn0qk0mh+056M+ZAcKv2n
7IybCppSne3d56EFTL6ISTOARk5EGud3EWzPci6cetG4lVpPgRorbLm/l/dB4nK9
MefxGgwWfODl1PEQEx33rMx6bVke4i1dOO8/1tbIq5BHlIxwDKqU2dP8GdfpxFw8
Kf1shkvcZYxnJMn9uFzZ8PjgL9lcfM40eDLC2lIOdnvOaftJ24An+HQw5uhwTtt4
TebQDIp6o28CtierdJf72dinlv4AFL0gcDEFSkr8gLDT96Feg+4eDIH91SQNnzVr
v62IXhsej65jYtub2Se64LySS4ZBLqIkaiJ3/rnun4wRR1gtsBCOSqfFfSRCtBoL
1OUgq3sgP0FnybaqRvezWPv+98VFo2uHkkJymVxsrXawnpBzVwdEMD2V905R432D
xzjL2JJ1sgto7a9u1JUKayNTBs54ntlkfQTxmfXtTBPigbt8w4i2D4tbVvnUvPzd
h//njymxzPTFJBtKHTTTyAhDFj5wH3OjCOQ4ANj+/anL1SKgubxB6FSMvZ3RGf6z
/jA4jN9ompXiBIx9sM7+MIKsbutFt5uUAr0q9gHtBbhH2SHSB9y0Osj2L5Hyg/0e
Uc6b4X2iZ+xTtU1vzeMSTTQycqdNZPe/ekqRL1giTZ4JdBQRZMma+v2rX1UlMdao
X1lAmTK2zsqyHtVnWCo3CJdru5ntIntL8gbdnV82bqwdx66xv6HEmSpvjn/LlESg
G0bD/2f2o6grGcx/dOyFTvHfzwqTVvkZden2aHA9n/g9gHcbY5ZaQ63TREJJpqqr
ofFKGRaA8iDKgCGFLpuywz5r0bRXokeHzjm08wI7M1lg51iME8k7n+JIDOnOEOos
7hkRGjbiWVPIWEuiRhGV1ynvCrdEKoKsa+ivMykrS8E/Zhz3+mJi0xRrIH39xV6s
IoBAmS6ZIa3zfvkK1d+lRiIFy0qofCNONn+KdDSCUhP2h3ov18UjQubi08CRcORD
im/RWqOp4H+jdjGHSVZa8fZYZODZZgXSxg02JoJxVGZcJxu8TEBoRjyy6opXrKBZ
Jq0ML7yLPkcpt7n/19saeN1ZEkJ1hw8R3pmlkhuF9j37KTAWXSaTxjbCYuCCywwu
fFGjcVpuaPOHSO9FW8o2LDakUL2PlCM0x4t6R/0WCUpB/xTvccTN+bFWpek6kmIp
awti7LO33joP5pEW1W6ijzH0c63+2I01OymPqkTwBtQ6rYR7/jHaDwYbAWhGifTR
4e130po3IVv7KmBCCpnOXiDZBD8TfhIhCiro0K9gnBZ5PIGf/fPpxRZYwWi8X4So
Qjvk2aFN9orv3IDdBnMnpCRcI6WRy8evD40DUtM++Hu6jQOeIO3RD30m3+g68QYQ
GKBDEoRnpy9neUxVig2fsO0vGNvy4l22LjcHe5l6L5MZAO6ixUiKowsAUjfv+KPd
LotZgzQuWzwk0NT1mVtbKM7D1XY/oTaRK1TZghd9EwJdHLRKjM3PouSNqFMaq8Fa
5GijUbn8jR9JdwwYk6VxPQbjQmvIkzjpY/U7lwlHLpu+r35Bc3xNyUwaDBTvnboW
9JmWTHC8ay2YtgKoDkfo2SHPzZB9qYeaIiDilzNACR7/KA8b8fAdoGaB2e8QKeT+
wcvscleF7aVfNWYAXnJeMfj1iod+kEc2kEx/hKtR4XK9wMyXQJUFvLVOeZx+U1LM
EWKkjkHayPA/NmsKcr/rIW85fx38WZQJU2sOCUPMLnpQRmODJIYM8J4HiiT2lhTV
9/fBoV1SEnrMnk5/iWibadLEbQep01WKwlEKEI8PYlNCJGZ220VU+Phn+vzlpiUb
QuZPb6mIHdBRRVZfpFsBqgQoncz6k9xRK7QT+TRJPW5dI3L9MJhb9mxIEHAlo2AU
Ne0IhaM4Q74tUbbTtDb/0S8KXdjNUNtTVbDFNymACsasPsd4NCtGYsO2+ay335fK
MG8eDZhrrRACjhje7q8srxok2GJ1Nh1XroarTuIjHdty3QnIbh22yoKykN4QTJuK
GAivax7nN/5oBJCCJHqdhd/1hbYXkGWMsrQdQuAW+xQCuMduvAVjC1AE5t4H7QWD
vbh+lOFtJ9qCDKy8wXpvK54oGWo4QCLiF7B/7UtLkrbppp7eMvg9nJTOr1s7/Tgw
hc08CrJ/0IHduVvOknqGzT9pMuPLUwwuy7XxJI6yk/k4YjfWFz9dyE/0L9B+KYPC
3h0ilfgUXHwvy+KaW7dkpBkFCFuwhetN6eRFhFWDMxqbh+XdoVOYIU9FbA5AdRGX
5p/UTtNFxPswtyLBX/xbHodz923TBYpDBh1vTqjKSLp8eJfpG5Q1m9Ym08GoRd1S
SH2yEg1spNaifb/LWSsBjrY1EotQKO95eEZ28YfG8XHtv4YcmwMSgrp7MCJ3+y/y
4bv6lLC2cKzpSSVi8Rn5i71l1/s5XMdKW+bf84lK+Q9Q4iKwr/tm4kcmfbamEjOn
wNscqREWVakUrdylqKtvuVjS6Zr+6HQHwmiVqZYpZtFHD3jbDhIUu5haS5kF8PYR
el7h+34g3lCtGaBlqS3wVO97Xxez2nEgBilnra8Rn+V0IE/sgNUfm1fpJY53UXSk
PE+i7Yo9y7rvTPqaaCyyz1Ygned2WMr4t2xrJV/3KBNvkejn06k+FtG4TJl8iCZa
AYxPcVRUhWQTPv0/BMqABe3mvCqbGPqbdEdHaKbvvK62lU98oK3V2EGDVsdIcgvP
DMCOWcQdM+Dl7C5qZnYx+Or2oBybL+2l4ZHcXhs/p7ejglrH4Tb7JF3rnALiu8O8
QcRz2FFWW1MRIIUhlXNFoms8hP0yTYVv+ueVlIQ9BeUOkJHonQv183YFTgNkmYFO
+2TzpdmlnEbLv2CnNsvnLJRmrpr5qWXzIoktdAbz/cvl2Nwjj23CthssthYoTeHp
1mrm2zYMbW0HnmuO9DmpNGkvYW2/OveYohxxndrjFbki4ne4iODeyEXOepLnA2oS
Id245XLPbSbb+W54Ds2y6GrrxzoOxiYfpJ67iTDAKjfJyCHVoF8rd9yy9WeNPGkf
qmV9vVMomyLvjZ7rTf0s5NuvuDGkeoBhGimXE2B1IoNIvkiv4cuCqjTSe4dicB06
GyQiNR5/LSjMqaoHJ/jkTqXCT2o3t/IPrNf1rkn/QI8dVap8jBjij1pnQziP9md6
2RHmhF/bRa5B0Rhu6AeP+HSfOCHyFV3K97qNqU9Q5EX/l4JXbCOeY0VaHotvNpZN
unuQ5tNpkAIJGxLrgbeafxuGDi/+XT/DEmfnOdH0oc1Thurb+phEH0M21uWWipnu
e3pN9+arkxj6kB89BTCm9XWoxxXYk2DRRoamhHorsy2sSXoN6WQzAkcF1u6rdi0w
5FYjyxXn3j+fzZ1sFfL0KbqjxjwBNO3tGNPDpTQHp5gQPItm4kTYzoDXFQFwMOff
K7m0xEr3WxAiLwsyuzsh5PUs4JgtuJ1+Xm5xki6711tI9kzBayROMoCc8f9ugYiY
amjj23FZDUo+CuehqhwfLwa+MfdgoGVqyKXYa/V+DHvU4nCWJhwbFqLssDTRHoyQ
0bPg6eURu3Ty1G1me5CaSYm9uAxh04gNvtb7DqPyBGbaygXTT/CAKznnXo1jBSTF
YVAfmHV+9uHLSv0muuFDPbyBLQZKP1NrmsWXouQe/s3i4i4nt8uHDVEo+RuLkhmv
7Lx9PzHPi/I/xhIa9n0U98Mj13aOrjMCvAyF6nKuDZSmEec7Fuh6JyF993auLN9e
3zT9QQ9p6t/bTrTv3mifPYGdQEa5IEtulskrDe46knN24AM7R4cQhYiRbshgdpxj
yfrbJOBIMbfIdc1e9Vv5cwdBOkZj8Vf5FMdH9LpYyt6UlrJRX7uxfHvHDPlklcOY
+QIndmgW+bFWdGZ6+ZQ9BIGlWMqRFUbBZCBoAb0iBylFWPTS6WLP/kAjhhM+2OaX
MZqHeFdBMH8mPgO9aUADPXAsD84z9EjePE/Boh+GXRzAusr94Uv1SC5fRNCFym+Z
YTAPbCEFqUfQ6BuobiciEgxsRf5PVCsXdTwCvTlLpfM5vrcHcvnb/KHj8phwe5Ic
l2gtnOal8bB86BD0zh/V/hdEoshzhWFKiJtl+GG9cLv4Z7OSiwIFuOSJs55C0z3y
a7XNyKDWe9rzTkM12XlIOCSwjBB+d5wBgdVGo9ImdnDk+bRPswvnFejKdhSRt6/h
x3Stz4Tib1IPmPwBQ1XTrHKnRZ/9pkBjfUZI+z7ZHvJgH+dyjRXFD3CAYpVZoBHR
h4CXxmoDnKRAADKF5VCgFTLaiHdgwSsUwJPoTwbOA3qdrWO4AyCUi79D6A4K1hxl
LAHt61HTMBu7W5qLfPdG++CKtxjMnF+Ch09O4IzVJ1AgvtOQW4Dx52y+dvcgYuN4
IbPnQAwO6uqKi9Do0CSGvOoHgQzkuN5U8iuefqJtjOQOGzvCX+3o+36ua8XGRb5L
mlnfuHff9xIKB6bBy7aViUHUmLP3OvuFoHmjY4zEPBxYC2wEF0DdKGLyj4xiU7ov
3Xt21dlJ4WBhH7gHw7Iov6+kKFcVPmx+WO6c1rxZkAp2BileJ9d6wccxgLcVGNjq
bbRPAmphxm44jDSVGy6o932WS2oDtJMl4KClSL21Z0o94mhJHmu7znFItQ7bm93q
q0vt9kDi97+15yWDcVJJeIReOAq1vBekZt8fZSD1GkkhT9TOVZgljnM7it3WNj3b
clmjRh2XYunYi8vQBAlwb3U9pvm7wFewvvonB9Tv3QnWkHYri9ZbtSJ66dtrR7Y6
KtUZJPkLBXonlbpBrV8Yrbsu3ozwI/ZROaMbyHRnZqjGZTHooP1/YTl4JZRYhfpp
ojSrMRPzTxWvNcnP8Yq1/nDgmGJkf5Fa/5tN3L4Ru4ZqcxfLmKWxDD8tw4gqzCKT
h8gayR3vges2zYGHRlL+NofCel8nJSHaKEfQP/0mnnafu3GCMU9YS63R9XAHUrzT
87rZqUt8rTW+P4r70cJKbnK5mlOEUOHXycgAjUBUVK1TUh5iS6gk395EEHIZccxt
74ZXncb/ZdwlPmv/n7Uin9whlNqiK2/VE9HogQ+n9L7B4LVSi0lPNLE3hXGg0R5T
8cwOTxm0X5bCOtKKH786ROZxnIS9gpKllrY+zIDvxLKSTsyCmlAP2qYYKE2MMeJB
Qp6ZnyylGMX9Pczze4vkLnaE+yGbtHlSfbY5suSmquKpIF+15+Zqq0ON3ROVhqzE
DMRdoFndIZxxQaabu1vj+r71IVUVZvl7jtvm3/67tU+nttt49rRiS9qpFTL6DGdw
uqdh41hH20E0uh9Z/n7kdu0BmlREwpMWo2ua7MjLATp3XzNXTmnRmcR2vBqfPpSt
k4mm6XJpDcgxsud/KJXqdXmUvOjK97aC1IDK9sq9c5W97SQkNOfE5d6jqhuw8PHG
9vXvswNEZWjTakyK7vZBEXGrleKMlnZUQVAHROlnvkKQeAMiPJcwhYaoLLXQqmn/
fgCwhxiS8xyIGcVtkcwH0avhsZuRuP2RoFz2xpfeViT50KVCUAukaffLMC1jbMho
M6UjvRbfrwCnpwJdEtRPKveGqXOeFXpvlTKUR2g6Jp+EFn2R+k308qYrrUriSjVO
z0WyIRD1C7jLyVVvqOG0nKZA1L8iiZZ6s2Q6iQ1ofBPniwHwo6XqItPgViTpxxcE
b4NtdptwB+cLB4bQWxn2qobNcW1YJ+l6shCToVtVfmct8Eb9F/YoitM8lAh71za5
H4ziL1T8hYUYxb2iNL11uTv4p70RrCW+e9HWZ5aP85W8+3HOIzQRp98O8koonLhL
aZbid78yGeXVpRdbSvr95lrs3G3CuJy2+vbUNudVhzvzMxxmFZNx7n8PbfZLvdwG
4yDHqxTBELcgQbUDwl11ATAwSwWjn7ntH4DHvp1JvDcE7sRE/n+a5vuvO8ZfwwVR
h+aKY8V12qA7yCI+7YYJtgeAptOn7OxWf0RuzjSk37wHS5Or/GZVH5EvKkW1jTFg
KwS5fhBKe6mM0j44w3yDxl8FCHxP32wYEAleUTMmZQipppqKKfnmV9g33Sxg7QPn
alFTYu0XEKhdurs1A1hqIRknNEThTQAZOPD8/39a6zpslx/L6QoQdnR7o4es1Ppo
lnRYUHiiCs4R5GlsHFhxJ5lSEP0uT2w/OECFQIsJQj/wR67oZ9OJSQqeAsmzj53v
GJy2tRwWeVrXPPMZ/6IpmpDA5ShsM0BcMPqIhUk/HY43FDMV4UspauXE0I3rXYHd
HR4jtiM0UStCb8WZL9ivVMEmwvltv0pcOGUV308ZPsrnsg5EIhyNh24RCh3r6dN8
T8Nt1cjyuL/aMHzzC3chRtaZC7mVf9jAIPeLmjVfql21v0nTK4R+/XpxviTp+itR
c629G/HUfygCIibBikqepdEiWYDocRt87jIMuisdUnIK7sIO7ZfmCgVcPFntC79u
pZWf7H1Zgv3BvVxYSTAvFmC3aLObZ+aPulPUx8pVXmprdfQmQB44Ag2H/HhXKIxo
Biu6pqnLApc0Wd3wNd9nrdJg9/Fz0qVGQwsHB9DWnFHT4tTWlXsiSZYChvuYf8Ip
SViRoKoCU8MbaCkmctTrwniX5U28OTK3ojH544pB/nsUvrOwKYM1/wBezxg1Xjoz
3DMqWcsu0u7r+fV8XNpSpML+pGZ7Y9MCjLS6iAGRyclc/oIRkbCPb8ml6dOiKMcM
DOfJ7+MUp68Mbbp9ppBMIQMDgnp9lt0LKSyUK8DNAPmCA9sQU4T5bs8Hu3K02CK2
2YBbNoTPQ58U5mFCLvsg9kTCShh7c/YyOh+dY1BuwZ/jfyCORyMoH4HiTNnSkTxe
zkCd8iR6yx8/z7vuPtAQX2icimof1lutFbncO7kwRutZ8R/Jvew8lcHKqY9bhP/m
irRDwW8X4FhiM9DRCyKHBJVCXyDw0u3FnFYib5j6T4LPuqEZDwC62v5dKykqhGO7
v+H6AXUFEOvTV7Kh+JOEMk13l53uczHVw8SN2IvEkOgsyZweUUcEQ5yACIVKIjoz
HP1xDZdZGjSdxCNzdnNZrmY2D+6gLT9IQ7UO+7BCL/mPjtBLXJLsD7AgDcsmmsC7
5u8c1Wz4e6j4hN98ajC/54DydCGqxDAih7hnAqSOZMRrpws4uHy2sIIE3dkOwnPP
OxL/qnGLCbIpho+SqWK/78yh8hOvWwGc4Yq3hq8nZJ6K5gZdFb/XG1w2jEFvE1lc
RTxrDXGc4xjY0hO9TJYANd5WMklSEvwWa8QZQYTfeW2Q+yBMvYrNxxu+ndYZUWDC
W10WDcpmETrZIQRnqA58JKJSPd8LB/4ZcOOB4LeGspnos07FZkr4N1yLLAhN0AdT
Z7ZFfyH6ORulhh0HWAEXuTXBqPW2lGqcg+A2eCL1wINU0SAuEtF8vstMNUjyBmi9
W7AQ9G5b9BwAK2aa9LKJ7ICD9PaYEQIHHeKuDp/3XPMe+m/g3nxrlyVoiX7v1xB/
GUoSMWjZjcgFImXG63T/SYaX5eyhuPuuz6ZQSn2zt8Wn5vbYXmmJ2fyFvBH8Wmcb
xlu5ebbmO0e4FahmzySozIbZa6kr05vB4nzKPHKynkwcO/+oaX+ZQ/+FxIqP/ind
VNw7ihrWuqcPLI4+8EWTPxF6ttna+hjoP49hs3/K41lJGXeTA4Uy6ixwocxgk5fN
O4ysB87W2Zjh7eIgFU9IJ9KSjACELBSsEwkFBVX5aHbRJpb5gJ0sDoTscg3vdtxm
k0HQpgxMkoL7WIIfVcuPXlbdrkp4rV4hQwl5xV3WghggxzRkvoyi1ygvUpiBZBu+
t5B+zVvajEXBKeBoD3AbSBjdpu9FkNViWxAaI0Tdq0cTWcQZeYBGgEEGXlwCUMry
+uXwSJj5d+oxIPe4HfrMoXJmosZdGRsEakkxl9TfNImaHEEJpjTxV4RGKczGM4uy
13+xvCv7LQvT3nRuOUcOwQtwosvMy0rwVy+yUIk30yi6IFp0PauBrYI7i+vpZ+Er
88drYvyC+5F4vV4nQJQhHjjm9wZSsAUCR/9368tFTUTQnpLgcNj/L+rW36AJdMwD
YJEVATE+s9SA/C5IYKUkWHP35XwTapS6vPmKR0yeWJoOh5qPAOJ7QroTCOxM9Nw4
wh73rCHmk3sRLfei4VW9Dohf/Yt36IU1vlshf2JRpVJiHAPj048RlVzOYQ7I5b9Z
h/1W66hp6zWJ3b2wJnuQprb4NqU8YfTCYHthYxQ0Ms2GwICrzcmmvdLYgYI3AYho
m2cbEPqHdHfpAr+UUIkvH37TbJ7cxD6SLeOOb0GiSgW6EmOVcrrrZonkrt653lGx
MPc45db6/4rqrky13sjVFnoYTQ8bCctxximmLBytgQ2emiPXOb+F71i7GMbWKAiJ
BzYbVj11x6Glp4pauDqAg8uzcfcoc01zg1wqikPglRQJ4ldWn2x/NOsHwFPzcOe0
vSqSFRduamSur/ORhegmDVmahovN4+DVmWISlkJdX6zHcZUmPuFld0Ggy6W6KF6Y
HwR+eKhFZ3UgnYfK2WY3OUHoR0zAIJrk3f9Q/XO2Z795noHJeljNhl/T3LIO/mNn
58GstEeazuyMzm0pXAWm9+o1jg0mzAquT579034HmU+/qJyukaHUMgKGdziCojJj
H760A+sVypoupzl0RWPtwwzLpNCelPqiH8Vi6VWFqGauUoJrqnGwwZs+oerzQxGz
mTVFxn2gAg61U8Z9O9B8UZ+GfjySXHmLo5lXmB5NZQQwJmbq6DdzvwD2V0ok9WcB
02NvO4a0LG0tqwl1gMxUiAuLgUsJ4iyhXDyNHDmluXoTX2343LkaOanha12VhiVB
Zf6FXwgihBLgWZ3TWxjH3PXM45avZpO9FsncSe96CC+SVp+OuTKdT4wI6fC/IlHx
1KcfdBnYN+4cnjfJBcXUn+OsxtnFP3bsXsX+6/hnJTwyFKtj2WfDMHbpWgrUq9mp
ERxMQsh5uXYLdRRRl/YKX0QLeohV/nLq9PpmJcBLgdWLUY2mohcJl3DlZO2khJ2j
cK/KKza1xl6HW6YkPaofwPftwEH8XQZ3m14ZhKIjO8wuNnWYMZIIsN3wz/NH5MUI
hU8Lue+hbvuz0+elJpZ2Lll4q7LF1Vojlp61X4lBjHnuQZO2+wIBfnyfWpVCVDK5
EFUfX7o5TdbOMGYc6f7lEoCduHdK0XIgV1UFFkLa3iQ/EWwdy7EJtChL0aFybt1k
lO65sgFAxYfuQoschqwr7K+eu5A8DmNl5xHQUuk1JaDoAjNOqs4PceiGqcalyn3r
vYKsDnHelzE1/0+S22AkuLlO9SE8pQCcm4JRTNlN8WtVfOnBKKyEkSSTEsYWoxnC
bFKadC6F4r50tvWahFz5wSkIpQyPu3xiYxEzeJnuUQqnCXZmA7Cb3uXQF4e4oNKu
9IRWkQgzRlkWak6dsluX0/jxyHXqNokXDRYdcVJHpE8oHm+2nISvOb20L9CQU/HG
ectZWOi4w317vHLGmIwyzYPe42CHVD/3+R4BfFCkbHdRUtC/+S73OGcHw2oHu2ux
q7csJDK5WMAX1qi0uuDe4O6FLLOCXy1oBivZnWeOUcmRsxiKgAuzyVWPgab1HcvP
3+ihuJ4Db5tn/76+WL7jgWYZ6N0oVxY8BIPsUtc5Xq8KZwbA/fHFsbTgELr9zmlg
ZXVhu/XfLt9tTrHUB/GFcPSfeiPzbLCcHLM7kLLQAP7sJSPyDg59ZWLxIAaUDfXA
+dRU0gHIUos/vMr5pDYX9zWyfNllJSCd6C3F0BLtUyqI+3L9k6oAgHAL5H3Av1B7
w6CO+yuSLTg46mdgbSLsJPsjlAWtMDa3JB7I2HRLaR3vVlfico5+Nksd1xV9UKuv
YIeeSnaXLzvhrOLXMacWXoLRYFGXKjjU0cUCmAqzHfV388XVEGIz3J4/tqgiLy4j
yIeEqSz0PHCgaYtM4PZZ5K6+sdnWo04JW2BDJbhDOBZnb3Uh0juNL0P/PrSeDoUh
vOdBswTsQAHH4dGr7qD9P9axzN7zyr99t59v3cK/f3+UtOBcFqD4dDaPtqmCxkZE
6qZZQDfFHtzMpn6IAnhZWruRyo1nWMUhR1YVttF+KZ5JfhdbM9U7UGpa8lx6nCBe
qe8ow35+VcPHXXw6bmrkVr6mCZf8WUUXNpRVofQbqzMrI+a8r0ib2E4Bb4JkId1N
o7UkV8ngSRszFDq8sQMGiWR/dx+16WQtt5exJqawDMyCo4Fs/CAjkkOhOCkW+mtw
y4M9Ufc/8SIB/YiYoxQPvBxHfTV3CBAXEN+Sy+DJl5pHFNL367wL6x2OMRCpamiH
gb5+mlQ0+kMhOGOY3aCLbgxfrrErrpnXDJey/oAsXchBvh6lL7Ve8uCjtaetrG0a
4WM1ZurFjesuj+9L6ytRoWTFXWeHOqBiZWREPu3Z6adaccQ0Jle/8HPCRwmmvcv/
y+L3Pq9m2mlwfJgufJUh+KdgVclUmDjoRd5NlM1OLTSr8eTXwR9cZ/9CxOuUMvcg
6ripx5wclJDbDxm/B+8GNvpg2vNeFKmawGon7UbRizJSH8Y+lhiNsFm1kdJvENzZ
F3kEIlRURUjWvLFYV8kbW3ZOAXMVDlN3mqMFBPFobkUo/XQCliRD9Us5N0UBqQlM
1j+8lgjVoWAbrB32X/0AOrwvuFjs5q7YdumhUCN2KFJuWTcJxRTbLo5x86DKbOw1
VpQ2Q2uQEW3+VUGd8t7noAOY9ze6TWT6w4dzduOFommavcTxZLaBFRpvyUW1dpwp
+GjgbY6HgNvjuu6XGZ75dFON8crnpqmfJg7BvzJOl71OhllklW//gKsv7E+HgSCm
HSgv3MNIJKG6Y/LqHfUSb1elBojFXoMm48HjCypRTJK1opd7AuWX3SSff7VEc1k7
ymt1QU3DEubbmR1reLeLEAWipMMEVrly7aUbHFiqm+4uo5iyzmsFIfwC87nB4e/9
37sRG/svkTO0ZY9tJAMAUZiVbVpe6ox/5yqK9Lq8BQS5ALJUHu/ZiP/g06kPYjwH
XGMLCDTnJTuQYAUe3V8ufB6B4c7USPVmzgW6zY56iwBHH9lULNgV1AP4C3MK4n1y
oUfmwPvoTwWdDhvLYxMCCzMZYzYSnoK67hu72pFvSf5ZWY1CoDpCn5/MnI4qcWCv
w7Ap4kDZHPBRbEP3+tOVbuK0tOG42w2PWs0KVxD9/5vHzBgfjXLsZgUwV7Yg2pPF
NuWwnUzar3EvB5KCkVNqsM7ZwadeHyTWxxMm+bXiEVtu+g7NpyWZy4zACkwQvcIn
32cnygrkZcI0uwvY/LInoiKr/gunTCMaUGyR2f31JogWASQveKUIZL/GuMkq96Qy
2u7IJxYYMcVxbhxakjlF0z96oO7TaibaHf5XsbXvwidjXyBVe3ZHGCmcA7frYtn8
7+4XPPAvKFGdbT5re9vA4a2nwHgAcsRbqB4xO8uNuIAuEQq6/3cg3mNej/KqHJjr
udwoST82cqz5IWynBrpBIV9l7Nb9DkPJ4vSMPLr/vp9h7xsc0rygzYlHbLOoFn9R
XqOYxh4RtFjeGCTTR6hlkWZg8yDe2pqdS1oiSkmJi7J+u8ITNEUteKIXDCpKlvDw
Oya+9lgTw8COox5j+kfwaT5yyw6UqFJDakdwheKfOEY=
`protect END_PROTECTED
