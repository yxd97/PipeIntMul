`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5fkCW9tvwtQEKjel4hC4a6MKjlO5gcmLqACTaysgZrLf2eGr6eG20sS6ktL0AfS
MRgwk+QNfv5f+Y2gXHtfRmLZPw5LGAmFceCSeEpM/upPjPResS5ZCbVWU/IYoAn4
vTCKX3CoEYQURKSWH8tz6EwlJy9wuvn+7W9jacOUvqDUklWDILlcQVjxc3M9pS7c
FQsW8+ZrfZmxzB97bKbHWTlZ2+3j4PNAx0sU2t9LRaniIIUuhXfQ2I2bvHE6JVf/
eEU8ECBD4S+OutdWQsTmgCqtKbagmHi1MaaFDHkwhhkh2tgrtXVdAHFF5Ol1mDMH
mI7menHXDW3cjzuBKOMXYIoR3XkzFGEeBDWn6TcPQxAhjss/dI2bUO99SJ9wD4I9
q6Iu1c4sYe8UCBRq8jY5G6BtHaABAGE1Qlh0uLEWB8OBp8DMj4xrgcmNiaTLsPbl
5pkgq1zRfj/CUbCSVAZyLfQPgIidf9xhr22USUPb08joN7apDMfF9GPstR0E1H0O
QzjjgRCj6MmgY9awRkGGxdVH+PR7LYJ9JQjAhVrqwrA7RxTljf+bNy051JfLNrtC
iP7YFvU8JN2EUKoPXMqlEQ==
`protect END_PROTECTED
