`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PvSH2iiFsDBufWB4EfJnL1azlzVmYoAPpeT4ZSNQuvlTnuJnpHPkQjCV0f29C9Hy
QVg8YgcT7t9l4rygxwggffdjuH1lwPJ4JRNNirSEj/eSZ7LWgnodZXJTT4Bf9+i7
qOU0zkd8eCXuShXsYbrd+u013stil0cZ0jqc3mfpEbMzTGiwTqQvhcoq9bcDsibF
eENOlga2s0RIvlTKruIzMQIOP0tYDJlms0/QH3jX1fYD0veUIMSO/RqBDjbJNm9y
UqijDxXJf5Rezf+RxH5cSfTngAFLw0kFoIeHDZphMIq+FbOSySkPggrFqZGGb/wk
Hm6LtcFAI7HoMovPNwtnY84Dg1x+FSgFZQcD5WKlcReYBkfhglt3wMHalFaABCSA
WC4/vCUPapI3M/eoAxv0nTt86YpmSwD7Ibb3HqvnM9I=
`protect END_PROTECTED
