`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6juDz61L5Rq/kW2W4AFBJCAxqjIp5Et0Hc37vgBHKbKHxgP6WfSOfNlwJ8QuUJ9i
Bek9eyASLY+CGA271E7Dp7TWmx3xySLFIdR2dLPKiPQZJ1Ao5jtKaZGMCgg/FVuu
1rHhGB6i5gRNBQ1qsi/VkzeJSWUvcTjA5AY0Us7Jh2pLXlrSyYQ1CR/fGY0iZjzE
DG85CVznxWj9PenHTbDK979ColSccsbZ8h8enOHeeQU7ETG+DMt9lgq7AWsVR+Xc
PVF/41Zds7XFhvcVw3x7A3E4iuDmd7H1eFDFsH5JcmimzTTd91Q19zWBsyk5Nfbk
U9WWE3rPADNqg3Z2vKox29zSbcSA3YsUCJka13xth5CclF0gYf4u9Zfa3tt0UmzP
Y7gUrP4BsiKolIKPBOna1MBtdw2XY18FhmglE+w2wP2C+N2WAIaosiaZTJBUnI0P
fMgg5ktHx7GxTcQLE488iPlZCzkGGBWYlVshUmkl33G83YxLO7fdTa4bWXhaq+qx
4DFJFohduqfiF/3sb6hqeiLQz1CtUStO7+R0TVrS8mJ3FxoDj+nzfIXo/uZxOaV8
qR5+kgfocUh0LZF9czikhzzH11UepFx6y7SVvtJFy4IhTLE/kTKyo169pVXANYe4
tigXpuzi/QBmE0gY/Ful3w0uRyblZz8ST1Z0zln2fXglIQHtqz38zOAHsk+IwZSS
`protect END_PROTECTED
