`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tqJaTqvnnrfFQ7n0HceLAink2moApBC9Numyu3kJHFD8JHmqQS0L/p4aHzaz+q9A
dioa7YCGzjjIq83wcUHChxie4z6pZYbGwWowH1GG0nl0/0AJHi0egKUxWrZK3lHR
uNxkpUUuZUBNNJn3dbl45CyYfAG9c+0mFP+NzvbUW4lTx+PI45PkMbgG9knsyMdG
pnVrTOLYjszj2Wwz0igXvPGGgGxyEMK3aho3QhqzNv3aKfMnGB6POcl067lJ6j+C
dJL459bxj5mHrDsAtJgZgLm+c1/nXIgxMglm/0lMpGrtdhhv701pU5bmykVIIgYv
bE6I1R9gYukSALqKhgn3jrKRzc3mF1HLhh8RpSmRKRcniB/2vfhYg4FcRzXGIh1X
vuc0QgjsBqHbc7Bz+eCQYmq6MTnYGp26JYQPLosd5IybsPtjWJK/G5jXlCfFZOPW
0meWEB6OSaTRlSJ/NDBxeBG/cxVokvjpvNnUir8y3H966kxXQN1d45nU7mEf10GW
wIjO3jcrFeRZ4h+gBJkSB7Jr1e5GnAn5M9qlmtoHnbaBO8KMC8bdkeYbxqKBkVgZ
6Ckbzj9IpV02un5EBlQDsTeNMIlk0pFu77w1Ojo36qH6WbiS306Y3yWbhnwc1l+Y
IhhnaL2PGSMZhskbnRp6+8thgYCj0AhQMAIFZTE8HD4=
`protect END_PROTECTED
