`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zW5di977XMhah5AKl2PYmtaJxQwF1OZkQczok6tW4r3mM8YKwgzE/BEu5tg0VcXC
fthuLNs+qOcV9vTrWakCM2d/yyexKmvjrGrVmJTs4V2SWZIjDM+3Mqv/KXPXKssf
sIZOYfIxED48run6m3YLYyaFOFegeiroPNDIw2mOw/pwMvGiuBNPzOeAGzjkmYpS
lXrozjdMaQJhXTmcLepqIHBiqRVyQQnsQ03I/0jTbLEKrj9JuYI5yzQKhVpxwIBI
KJGSgszRZ7RvCEI/VkTk8vkySnK+CGC/v9z3MI2YDoqNfrH5oP3LAvd5lmoIWRDI
dIB/6MVbztikyNvFz7LPhzMkbIYjmv5CbaFKT2L8tm9A+7Sh4tQUhWwT7dux0aha
yUQHozT0M1s6NeRdks0wsKlP/SVt/pNXFwbVeZsx1onTHqSV/S9MFhqM5eNyxfXB
MzqLTHAaMwnGJ5QuvElcfNYumThIgf3KlKvDe6c84d8vw/i7E7STMOlJpqdA5/m8
LNI6oZxExykS1udo/et/sch/uK43ylHXvS77Yc46Dk+eLDulJ0Fy7dsFwTewBQOI
Zu2X7SbdMbY2XlEUfv+HR4pYPl6nsRQn9UJX1/WqvIIj0xINdKARFzWvl7FWPQBL
E9PdBnQGwlIZZCnoMjnMfzX8amGKefgeVu0xpZEHOdrQUjsY4lFXVnyWJWgD9Qr0
oHvwcZ+SNt4P85sKZJ0iIJwVdA193fEJwVvgM0hPNcEe+rgEpPJgejrS23R4vLW8
xEdnao9PW/8SW47MR7IuwaE3j5zWGosTHj8g5ym08AFAmhGbssYzn/pn6rLybKb1
Eo7L1wnlUByM4aQ6RTquSpPTz6I6xt4Ls6jQPcAP0BUUwZaOhD0RntJ0P4Qs1g+9
/YYPzvrHR2VuVzFcyklUQ2nkwqumZGio8Ncj85tUm2NYUNBFq/uV+gkKRWwPoF11
Y3hUEcY6qN6pZNEVbo/wPmtqGFzuOuDB1cWOh82mku82XOtgHXbyKEVqf2PLUc8D
`protect END_PROTECTED
