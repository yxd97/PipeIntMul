`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oy3c2SOAcwPQsqF5kfgkHJYtbjfhRRSE3bz4QjrKouFbr2jbyLjZp49/RhHSh7oL
0hBZacGaAWKJ1yNFqTBHi8bTLuQoJhlPQqPQCUybFr4kZ7gv/1xXFM9qLhLeDXpt
tlwMVG3BRv6Pt4MRO5RLQLa5U3XNL7hrAJvhyzekQn4VxwLuKvvr0x5NTTeY5zEN
+TGAnm8nBDbrunpYmYkTp6aNYh7+oY/VR0xBu8JN2C9yi35sEpqU0iEEMza/DVUo
kxwxyMPdZoXCWycYaU3h5NQt3y/XIjAoJrBT8S2dttpYMlYvVQAX7LLpDk1rLPwJ
egEvDwgbquoxl9hHJppzKWeS0/KSy84kPcajhs1vML/Mt+iv4G7Sqq2AisulGaHD
HuYBniNDCmJUjtZsxThjirixBVuqX97TsjeN1MD5TjCyY5tz5mqheBh6FXMaub0/
rSszxpvW0vfNZ//QsrDWM+JrVow6dAj9CFWjtvjk2nzkwrDWhivOQGKDJXjWvc/Q
CdJfYWNFveOUSzLs+UKqi/kIYwb7t/GQL08h/4pjQcPkHUPfP8NAgk4f0lligBOL
jrzKDn77d3xcUx2UCAQwi3gl6aMWIP88GMSA2A6HCYM5BOp0N2pqTjdz+Rf0HuMG
fL3PwWcSqWM5FOtp35Vxh/atuEdnKbvYd6QvPZ0IWCkN7jewUdSJNZgdsWA3S8Fl
S2kNr4NlrT0UEW3Ecab2WnQ0Zh+lsmgIhkMr9UieF/b2R0GI8xtTr7Mm2XuBMf6O
NI0FwWRPYMVSn75UuR8MUQVHDYrhgTiSl8vwwsyBsZuCFFT2Wpq2p2kJ5tv2e1P6
Tn2RHAIh6qcNmLc5UYbUb2xzkBke+jkUVCgpk+ASNSn1PJDFQTSN20OB9O8nycS3
ME3AlaZtqfJq941mpOo98S3gbnLxDYraax+OwPKvmh0Lf9nPL7lBn3c9iiZN218u
xWG1+MZxNBIabQzYKWVt5QKJzsc6C3Sjylmet5o3L73Oh0VZG4oh6q3+EXZFXdaj
WZVbtApQQjlIn12hx7IhQI+9uU52qZ7GMStuISd1P2MwFemua/Teadtu6QbYRnEV
cDRijsSG1vMM8iV22v6KuvWxpWuYhlMqRCciNjw5EXJqjZ03xJseyG0v2JFKykFZ
wz5JdMPlmplcWxEYEfTPzSE27Aq7o2SsCBm3f+e8whr0eHKvmCVkWch9fAVuxvpL
9s4nFzUXMn0ddGe/NYOUUDMaWIm9dyzCiBrbQgeRLbtfEY9pM+HsqG/w1fYQpESa
dNSgmejgKjYp+miCIgqpFVNYxFdfE9HSxatMHMUacsKlymt5i9JLcps8MdPc1xaa
Btn5MhAditz9iRunTIuZ0j8SmfB6Jn1f7NYlr99MDPyRHIpmUrWfPehsEBak7bvo
K0EFCK3Esd+/oKX2vVFOWQmnNclfbYkPAOZUz9ByfLNYG8+S8/97/BTqdENfgjxZ
Pe0B62/MR1M2xwUSpHRDCxQH4/AzD+xBaSHUrylBTcBqyDt5t/c5ThE3k08r2dXb
85hYC4+1xV/tJLcA43UHnB6MtZ8TVWItAIkniVICgnf2t+msgAT6Rw3EeyUrryPh
XJPkxSPWPOKB/omQz4AUKAXTSu260CgDms+he6LyBJwT3ewkk7uYW11Dgvs75M2J
PYrd+KQIYGtObvwkIIdem+NoMQbqHcb8MNw7+mqJp4ZSUM68du4B6t5SrcdCTPfJ
TwtV67HVgI2FU5raPU0syH37/eIpINU7tSskOGlVv72lvUKLekWbdf4E/4IlcEVv
QIUtg7qihCJ3oaE/yMcBun4QajEaE118uMlkQHigvTBCyhYtf1y54Oreb8j+PQ5q
/Uz6UhDn53lWCoxqJB4Z+VsyAfb1irKg4SEGP1b+BLlnqdUe8UkBuXtb8R+rlxGZ
jbBq+zVQ64nV494iQCa9QuQvezIioVFe7aid240r8CnPzWrFNbKj406iHrIYok8j
l1EwttjD7UXetEZcwiT4ykdzWv2/ZIXl5MrwaWHHz0P7svxHptVrMaTX9ihkDnu8
PRbZwImbsCtJpTa9RIHiWp0ft27eOEQnAi0mug5gzkxSAlyZqtfMg1uULdqrk4oT
pKs+tmEI7w/+SrV/TJxZV+I3eOE+JRZNyhj7BLII3rgyeCBqagdjR3gYD4KNZm13
I05nuqUiMYzgFDrzFfm1aAABFQtHEMRmk6uiMTtOkLLnHr7pUcL+srLyvdejk7gO
PMkE+DErROMmoM+InKMSPcMDWK3atrbyrriK+oRpwfTUpMWh45KrsKhRBYFbyY6F
blFeaOxYdoH6MnRGWGa3AC4cLjmcvLqZxoH8819+ndGxhzqeAebyNHTLx2YkYm4i
iYP5FF/RShtp5fM2zNz/kz9qZv+DCbm6pLrC3h34MMA+fN9BXtOIyfXvZvZ34kp6
U1megKzd4uXx+7kpCsxwGNUoi8aGCkFxoFT+Pce5XF2Ai3o7EOxr6TAPotgRk71v
uhE1eIGAQwxaEqKKBqLuFblnmnG4N9FF6O8X/HB8j3TTKlcIUkZ7D8whOdx9+n8A
ZeqVSJKbtMpKM7vlFBckt8hoyQHXB7G2X04rvLdPwQwx47VDZnQDlwYvWqDQTGo6
UUV5RYiZuCKK7vnYgm9ZPXSHHjHNOndUsQjQgcNEwdqCA2QTR0M1kBwgzvIpCANu
GPsTdbP2/cBm5mzMcNWXU5EKcmUYR0AzvFeUclw/ByuPDNKjqSJqO/QtrQ65OJ9S
nb/KjtUe79E1pmLx8o/abfOQj6kQXbIxP+5GdG9TwVjIHJQJzihdPL6gAAJtYFVY
IpttYDQZg4LLjLCJKbmv/iGUmPz+3CKCFGdx9X6sBuIc3NdGJDToL7zZBNTzMKc5
dVXS3cHHbMw38xbJwW7AztD38fV8MNRjvXWVd1J6kiwTuBd+8GkoGocEVYMu7z+6
GMa74xBFk/288ucBNtz5y/MF39XIJ3KZZ27I60NQ9Suo2PQfiaYjaSm3u4fVDuZZ
7EOG5oqL1YvNy/y6zx+TZZbSLkCBsgU2L9yX60gMnql38+H5bPUBXl+Fi9eUjWej
sKplQ2cIPa9OKeJUAA7J+slk/4XLg6dpwx0gQFCy3J44yB/8iPWeaaN5Dr4D4yer
X0fAUEXK3HWWJ5/6k4TtJXV/Inn3Plm35GKON6IoDiBjNiaiw197BIAzZj24E8kV
yQ+YKR0qMfBhkfyolzkGj3D5Rwp7kwr0cfJAldNHtcrM3AK0jjsdWpW2oQAeVbmQ
8a1+XscE32pPpiEsa2Gr85ayscgqUu4rbdl+z/nkv2QJiQEPm6H6YUq/RBNPskc5
40ShHYS668iA4nICnOoJfBNLnnZ4PK9xOYqgvqRJrqEU7BwSbgUKBMu0mBnJVAKx
VkOsRjlzGR7k8Kg/hCI/yQefWhIi9LBhwAmMtPCh09GBEvrzhs9YYv77sTwyTjeo
NlrNON3npMtrGZGOO/SkuvN5V21OMOOXpFUeO68U+qQziO3u96QvnGrIbhpyHaN6
655agMC8FNbyHdzL62igoYjexq4d14d3g8V3HbFUwQWOPTuynlaky6ruDiBrgJh1
tonVxBrRFJ8ByrYMLMHokq413+ZEd9thkEEUi/ZBlJ06AA8QylrgoByGMX7cmlId
bSmQ3wNvNNixYFC1X1UC6ph+il0ypLDhx/+ieoLqs8duMD+MQWn2hjdZIHrrSczp
tJhyXjzXpzd+D6ZRIGyK9GHHGKL0T3hEwiVhuJfbjNUgYPSP1dbKdpb9dWQI6Qo7
5MZo9MVLi2sSyNEF2qrhCrY3McA+vKiQYY4P3MLVTMdMr2gZGIpjxI61gC1IzJTZ
vchIyYMBG07IR1bGOCPQH8M4qhM+VEOnZON8rGJsHKAEs2r0dura4tlB5S8sXi1O
y6msCAFc9oS50TQ/fqFkTOzcGrUmGTbSgzYY7ch2+lw=
`protect END_PROTECTED
