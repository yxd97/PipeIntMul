`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZmt3mdeyBjWlHduMx/Zo1SwPU1kkky6yxINvH1QOc+voBrkkb42UwZGYlphMkS7
IKCvMBnAgm4EwbhrQ9I12MW9iMqKqkto+YqkXv5zzMwZuPONopfxo4ETEDZE4iea
Htq29kexU3jmGhE8zTPptbHDaK2MHbCZwQZH+ft1v4P63pjexKp7temi/Z5d1U/7
tS2Oc1TQ23+AKT+eTg9GiPggiidkhgipdT8Z6KJbfqky3O7grlnGvfDLsw/bUYLW
/5IIxljKGB5f6TirJLlMq7HSHQHPgiv9OeFbNIOzwAB0ih5Cv5ji/CanJtyTLiG4
WI4fnF03bipB7DgY8nQlag==
`protect END_PROTECTED
