`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GzkK4MGYh219+AHktQEWgzjdlQacNDZfQrhSl3Er1b90SOPXC4Bk9oM85cdFD0Hj
2mujAwI/sqPa+YwQEO3Vv5PyfKFLfbYsjL5jJ/c+WKv2pqSqHLwThtG0xUZgLRRL
GuG/Lz2ioC8UBPIblmMqEZOwSE9d6+JKRguzRVMpP4Ek5qNOaN2fXiOn4d2+I4Ta
Ptk0LvL9Vh835yWwCgsyMoSaB23ZNhwTDxorZIB6+4x5Mw2vbgV38WzTSG8pIqAZ
j2SxiAPAU74U7nw28vQEDO++3G+8DlwSiui+phcBPFcFzDVtv/OfTGcYT5dipAjG
htm1RO/EUek11XpxzgqANHjpLuo8hCfDG2yrk6RWHXmoJSAc/yx59zYFw9gPJp31
Hxp0g1Wz+4K5XBKaane85mmghLtG1qrDOy/E4G8PMx0mbLRF0vFLpIE1VADuYcvX
bALebFRjKvQuASCARI8pp/vjIV94cUcZsltafCr4rADsVGmnWRhEQkwdwdB3L9mT
Rzv07R9YYxh3c5J0ooEA3h0+D+K9+26MBS7QvelenroRKyBxA5Pm4E4OFqK8eUeg
2PsGVP3CWULfKSqrZrwA6u29vRfewjejfpe25dSDbj9qTz93eXxfVbPSakFsQBWQ
`protect END_PROTECTED
