`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5T0XqqHJGj9RncB8VVowfTYUsK8Vgy2qcqQ7nM0upzoTT+ih8CqXuLiM65i+WNSJ
n8TerxI13Ok99E+VbYqQh0rxUmsSVE7Amb1QkbOlYnIrjAj9H+unUjM0w5MCFjjp
9LDHT3xrNw4uGdxUb4RuK9BfLoZyXmM08oh55WsKJW7HKI3CMPjSIVXdXdbdkhRP
pavAD77aXKPZ96tMutQhzpwHk4rPFFZ9vmiHQuAhme1mSfq/4g55EI8CCScF7fN+
zpuzzHd8hLHoXuqjkhUhQ0d1oMSmP8bCrCHL5Fj9i50P8u4Ibqqu0r3JYNT9i233
+3AobDyR5xu6fYqiJLf/tA==
`protect END_PROTECTED
