`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8kJc4XlOw/JieThwKWMkVD/7LC4nHOHvD/pZ4JUH5gx9H/LKjuyYQp7tMPE597c
JUtI9D/0sdG1GXGYRJHHGFvK7dNi4pWmTIfFBPj6GamkfX/nXIiuMPCdVSVygs/5
jeGyVnauTFrRsDjBkzMwwgtaFstlN7/T4uHCLtzyVgHqcj/lK+5iIa+VgT8fDzrM
aKsX/gkZvdRpQR7oODRI2JpFwHf5CLpFR/IUYjqLN1D3I/F0ze2HMajFB3SDhPtm
Q7k1maB7qx9MlPj33Aq8Mea3m+vJoRu8yoteIB0ad0pMjBpoM3gfnQkfdV04Y8/8
rr8rwYJ0JVyNroz+fuPNcDG6aSbsuKeH3taisFdxMuNdUohtgcB6f49dLKLo7YhC
YkqkwQMW/gMNiK8zl6+FXFEl1p0Sqj4C5p8Dm4K9cS9ir24csnxTyXF+eNoUJVSM
t/ZTO0NzFfNynaxVc9XmIxsbcF/WgHLBXP2SToD2kL4qLGyCXA/PKV8Dc+hpt8wd
HTlg6f0di2LPBMIdQkMObCnT97SrDSKsmTRdSEMptnjv/FUZXm5Ov1yOdHQbm2A2
jUJKQ9m+u+u+9Q2+F0MDKcVQaDZpfCTz++CJdvt0Yd+2SPOQlYiRIRvOfXr801LR
i1xzzcaHQJ2BrbqTUUr9iKL6LW+IIFBPR+s1wd2gTIs=
`protect END_PROTECTED
