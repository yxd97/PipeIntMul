`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2vkfFYzkBXSB0L4O4YP7rvzoIe01jRn64DoM/WPhubl0qHhY31npUFHnENgxE7+
CXx4jk/iHpMvHjOr1uYpvp+CByR0WR3gcdRZxicu6z4qb7wUzb9rN6nAS+wlGoTF
z0Yk5osE90gyLU1oxu6HzoQaZkKBXAQl+cXtZjpuNiTvvh0YlhfSm8ec6sk5nURw
5sIUyt4kI8qysIePInhU+YwyRO5ACbbZA/JC9PMJr3F5ewMHh+c9ccvEx3M0azcN
Y/hkklIYqvXVQHApH1gMUvMw6hydn4ykqEQ0vGoCbx94uj1vhiZeAsGSO23k7Vh3
OKYTCymuEDMeqU1u10568pMkxepIZ0xVIx2Hoyq97hRDBlBIvjWy6+XpiNRBPq5w
YvpHQbmKOgc021sthr8fBIUR6LDZl4tZF9XbZvw5mA7Zh4o6HjI69ytRbIOtp+18
YMIg0oVEvw5E4ig1H0JTzEcm47eArhGAEcOMuKHZNVNtZ7ECWyQkcWUAnxqhEpFi
3UVDKZhQ5oRwU6uLrg28YtEyElNTomMEvdyQfSfK7hUZKGGPegYHNtI7dBQH6rzD
xfANAV0GR+tahtB0jiUVEOzGjW5vKt5K8owal9/L25iZXQR/kBomM7IJRN0eG5Gn
6a8uzSYj4gEiaHtKa+X+mSopUHRNWfna1Oq4DQS65i9YIpyyloSCTTScYeyL8k1O
cv+TyzCXc60iplCNaKa/iSjXM/wM9X00bx77jx1e5MrS/6TjW0BZtEkQkiQDO1fG
P5YuhBPeTyWtXW0gEfeI0g==
`protect END_PROTECTED
