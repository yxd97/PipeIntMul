`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3n6BvsfjZSQrM+W6MCAKH0uTDxUgrbr2eKouURICUHyaBEAoPzcl5r6HSarruvY
OtE0H3sJY28DuNV9OhWy7q7xjugEvf7O6Wb2eUVcoRxtkM+mqwAbtmblqgYwNbLF
p5lLN3JV8jwe7uQrUtiPn8Tnuyt2qxLnHMIBaMGzPDi4coRUupSlpFGA4ZqfqLN1
khcRJlCY2ilJm0v6ehYrzvzAy0uPDQRpseGmcCA0x4VzWKrtkP+PwfoABHNaB5L/
ZrrAr5q/m3DWfAZ2LNMwOQAuXIDipitFJRz/lbyEziC1eEaNX9qK2CatHSq3nhNR
4lrFlXLG7HcEZCJseC+SvsWJZ/0sTo07F9INnzKKwenhWym5zVnVI+h1zsxlPyRb
KdGb+cNSgGKVx5XYbvjcmercz82e2Ah2Zvkf9TcNMZ4=
`protect END_PROTECTED
