`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
urFzgxYBC9kHZVSkRkUrpKK3wdidVaK3iruZlcA5YB62aBnxFTy7WzjMwDF0MxIC
+io9CYX3YBoIv5+oO/c70y+72xr/hlk5faobdeAqFHn02kBkKccjc8WAlA4vpsME
5C/gRWj3dDaopbTiu8x9zfOyu3FYONQFvH2JxpA5yZY=
`protect END_PROTECTED
