`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
koFeYo1mTrOpqxCV8lj9uDsKsHolOynADcD8Aq1cOE3lxQX/6KY3/EBcblHM0DLb
5TvUNmdIzuTulezRB0GH0kaKeKU5q98Wi31OW7im30K2MzCbzUNy2tV7oXS+LK57
ejos6IKPcB89mclXJV1v4aaBMorwirZi71+5jqyB9TjI7xOLZd3si7nVE7lw1WtT
7JoJpo51Dg4Ir2JW3OgvloIBRra9YpvevFKx9BFubHpX+4q2qmPzqEAQTo2/1gJU
kiZ0BfVGu8oh70HTT+KPDp5W6eSmInFd1F/crxQ4I09tqIza7qeKglzRkP28tljh
cs2WGiTGFO011GppEVLQhgAcpemF1ALskvH/JmxeoaSQW2kDRLTa1HI84IzR8e6n
4gJsvPoX0Ik6kcOjb4wl6I8+esl7Ev8jCLDidyvJDd4+y7q+KK2ibeiuIaD1FZ2J
`protect END_PROTECTED
