`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qEmuyGB3AA3Vy+smJv7UTbAx6vheuWwvhnU6awL/Tqxxiw2aRHlUqCvSE+xrQk7t
5aCBaxkaQlAtZ3sHZ+50WlCKRKn/K3Y584Gq1gVgyL0TnVIqzSOVATj6XrmrJX3H
vUR6832GKQTp/Ms34Nh6RIGyOgLLcjW6YNsrgqCcqj2OpCkNyvX75TpVntK0LsdB
hHNsjQfiCti3CudTDx+H5p3cAl+Sle5KiI5vaWbaWnGQnfAmauzYNOGL1AKCSZkD
ur1dkB4WD/kzPYvxXBnIx7rMSahx1k723e952JMUXO/bLVk4nUSmv1UcWHJ/WfDQ
KGvkMPk65vp+GVVgTUIiRLziIDn1bczQSoIka8U8bKOWLNxIPN2hSXpE+2D/t+1P
6F8lhKhsjOOOSXm//JRNdBF7CSHiGynFFpLnKXUiNV1C8/9QFv/QCDOVyDnKXf/s
73O4awpyhu7ii0334aiBnEwkVbo9/HxLqKG2Egc0wHx55/bi8/IeTPSmH952E1RK
9MAD0WSltTVgcpu4dibiQOHOc5R9/fhV6pRXxajMAIXJ1OQYHuGi2Y/WHPamym/N
kv6BOwTVSkHHstkBP2RB12T0FGsaIn/V7x846blf8zPCbIDyHyet01Y2ZG/QgOC7
pKsBSPfPqi8OMs26CGD9V+iioYBolQYxE387OgJQbqcoyZYL3eS56U+tZb+b9WdE
HfPjCHgqypEWp0e6QYlhKAPjhafTnTxKsKkT8npU61088PJxhTxC4VhLauNwI/Z9
VVeBye4WptAdptAyL4FKmuDydxZC+jKpLPqMGXOnOSOnqFykIUHcMZABi/0y9A59
LwtyStL3Rq5xEIUzutkcQy6YFscRjY9BXvm8R/ZhcmEZk/VsJtlKiG4TW9+nnFaf
6yDDcYcmT9Iyrzalgx0GQTZH2UGtH+r/P+CQArzBxxH1gTvMiVavl3TOWhoUbWp7
t0wB/OOXaJr4gArNG65aOK7WR9FO9c3x9J/4NfxMVCVrNZbsfgGK+v2+8xNbRQj+
u6Iqou8v3IX+dnPQy80Y5xtDXH27X/d2uxIellwAnVeGPW2hSV8nyx3szMpjjL9o
oMZb4vnSuFXzNUq/zV/73X6Z7ITeQaCpenTPgauyiFNhGKi/utyx1dTzjTVRHqs2
SH9yz2rq6QE6fiXpFwgivclgZUPz2v2b5x9id2E5cEOrA1t2+wa1e4nKCOtTrNQu
1PjtzTqJQHoWabfM8/Lfe0cRxo8bbFvILfj90HfwAOp+iiQv+XPHSxI/J1aGmfxP
FQw2Qfg5R6EwPZEvQQlENcl5jloKCUW5uKxmzHEYIvWEOEDSa0ZpvFf/jw57LpkT
qHtzteuF6zDZUDeNA45VeLuzly9QJsRKp6mx3yRpbFbMFZoakzbQNw+IknJH8pPH
5J6jwv8zzMD3FL7u1as1WRs42ze7qiMuWaCNUOjlsdle5FBcerCoRzmqZHJX7z9J
y+YJsphDu0UPxJ83FoiHoBkd8vqH8IAfdYNpqXT5DCs4/Nh2kGkBszxpQ3tf6QoK
d+TSrNdzlz/sHmCsoPLhPlu4V+hIgkUiCqYHQZeseVRJMEefS6fUU5SbZTwaJ1Ad
fcTatiZcKNEnajg7zZlcrLcNI5THVlh4XzW/i0A90iG0aYizoPOQMzUVhBQivdXN
qAZeS1rY24WwlAnfGkfk8YOA32XUOgha0wdfSlHF6gV+ShoGbF8uPAB1EliEXB6G
owlCgha7vOYNixeLLCTOvhlF5Ao0cErF6NWlH3EPVmuwt/pYNmPjmANpfdOWnmgy
wwvAA6X50CFnx+Bgw0c2kZ19Y2ZHnUUjAEo9ZuV/5shuh1rV+oA+HqGiW+Vk6a6R
`protect END_PROTECTED
