`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2YkKq8daYYrkvjqB/+JNZI156dIocAFNRuMG4Tk1caJCa7MWJt2AOtgVmzpl/DQA
5iHkErZysjTSCHDr/AVDDFGF/8k2z+rqNyT8YWxxsziV96D55EcmItpuiIAYH7RV
P/+Uk2mZxQtNxCA6koRezc0sBxnQ7h9aEaNYSsP1i4VsagTGf+2qOa5vxJ1+qXxH
9yJajqwZqj5rv92UucncM2Xansj/z72mX6XOgMK3eT7wOmBDsuiI+tclTI1IJJXP
XLqUnz8Q3kKKKYDxAD+6nSyZyCvOTnhhHtAz7sVC3zZZNNMqhLpQz44F84ODNwOG
JVRV1Ta6+jD6Zoyzv+eGTK/ysty5zIeh6GCewDqxf+0=
`protect END_PROTECTED
