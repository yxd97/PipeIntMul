`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MDFfDlTBYSnbIFVbUONw6wAmFVYfOvyLJ0AUf6pSFHUbroIP/hahWSnNb5ApK6u3
w86T4YUMzhgMgK4wqH9szkd5Qfjh+GONHHqFFLCqiC46eodMwWOnMe436BAB9bvi
SrZxN/GFPyoE1VF9wEHUHAxvb/6hxVVZva2tOhcQbeg84HhSr7kCgRMu4HAR+Z3f
aFNj+UrY9yVG/b81LamIuXlfwXoao2ovBpxFNuou4gOA8KQcVLwFy6Y/i2lmrZAk
OeOoXjFWh5atC7d9qdTOubgNbjUtb41ye6PGex2Mz4XS/qwu6en3HznN2vlM9gAp
nWG2HLi4HrIA2uJoobOj2tRngc4Gf5XceiE9xIt99T7/yV+EX/lZkYZsMozsMcnQ
WQ/dK5D7sACwjC51f4OJ2Rsd162Oex0TEQDao3DJcmATUcQ8QmNis7gK/oNY0nJM
fRhOXCym/tWcdh1cFgJStC4br0TLCP0xM3UepeQ7SzRaNLwWIHWc/tnXai+YHbrF
ewXE/Ckzhsf++MxausYXbGzQhXv2BxXDbEhcSCs8FOsd7Wsu0QfIWVrBlKc60Wn/
rw6qqKy0j+2xIfk/Q6xofPHmlmY/x1J3mG5gmGuMWlnaZPU90DF4M3LHGj/GnJgW
AZgRHubGR7kUUgEeHA59x8ACN258IhUF6t8XlWoXjFx/nGm9Cu0nsHtMO2sYzaOD
XXQWTW4sGmH+0qDhzo0i6/thHHZkn9n3e/BrSZT/7E3fi+mnDFKQgQsI5b3Jc1QG
9aasFF4MwvT4LsQQ5kGwti/LwCNakGE8nTx0bsr0FCzOoBFTEdeTccLclgmBjH9A
ndBYcNZHdd/nIJIY7KZBSU+m/5at/oI6+FY9yvAuH7i7m4fde1JoD8RlRLYJBpli
FWoRHT5II7Gq46l5naAuclU+6s7744+kXGydS/dp7Lat2mTLCVIBcZC81KG9H9gX
8c8HrYF1gWH3RxJFQe03pkE6I++M6XCYP+Dbj76Wh4QWWHsbbJ62XWB5RzHsRVsz
Y08tzmNR7NwAVDD79rOo2qBsvEKETcv/kPvgoLuTLNaz+EelzS0wRUsQrf5x3PQo
V1Un/VPMccB1wLwFk4B2gy/OlT98tbicMnZkaRz6unM4p71SFmthYDp1piH8Roxs
mC4lxNNTmzlFQUqR/YDnwfZRawTA6kn4IJ+/Hi/9sywdpV6tbLTMUDgneqj00zLD
bv06PxHeULHJ+Gx/KIl2eLl43STWLGYZfgfBwRSweL+R+MD++qSAGb+eHHYTa7ET
yZUYxX+hhHTBoMqbzSywbYG/UBQnvApbzoDzIaHfExCWJ6+02Xn3vgFK9P5OufOt
QR9u/3PPrt0rJqBNeT8XXTyRzcpoW1mf+2VwMTxqDZ5tqWL66LnksFKiik/T4UeC
jkVFhtpDAn60PRzVIJJbXgaajHc4W66ULeq4auioqaXJgIgkkeM0HoNwRg8DKhcQ
6bXJagWwv0BsgbGMXGWL/IcLVPfZo9f1VsYy5MUCiEwfmfzmgNoi3yVvPL1WWKPn
LkcRc2GxwVAPBfblb8VhtXPtuMLzcNIhVW0O/4MM+uwNDZnznDjzJVd4D1KdqzJM
vwACKEQXDLNAJb3i+0Vdjxpya0J/ZBsBFhGu/yf0HTgoAnjFVBfjllEPH5lmHTek
fnmaoz0HiyKJBxQEWuoHIUChKQ99NmYTgK/9osRyyqphbRUl+TtvZV7iFDxnI5Yy
W8y4R73WLvHdZyaBlneCh9dINFnMQw3ajUUhLfMEcZ2AU54LNgY72kjRsW7TFYw3
kkgt0V+HXfE9ErWhjyTrcEUqCesuHfH0Ou14Drx3jypr+bVB3XybNrqi56yJUtNg
HuI7s0byQaAtGh6/0JLVcceM+kwFViBRI6FP5mFM5jtXkXSSQJlxIGn4YbuUAgSm
XYMies0zyjBPSIFjWt5kIRFDgPXH+XVDHxiKyuimEDmnPhyhhlx9EEaR7pCX8KCC
OQ3h1QUV4pKjxFGRyOdnAEkbFDpT2/2yeA9Pig8ILDIFfZUFkzKRDY0n8g60l3Fm
CKjqMHZEJMYWz+GvuKSZfDSAusyw8fQ6SSK1vDfOWK7Pm+iCpmtbG19PTGmTbajb
LlYGEbzBz4ZDMNjH0ki8PcGuRFe/uiiLi662L5c7PzBxH0Ogctt+P27kXD/tw5rl
iw+aCnEdbmYAM+7yaTy82y9u8+lxKdSUs7/zkNhM4NZe8j6OoDswoC7ogXHe7eF+
Cgm4QirYpmU0ItJA1EA+f9KEHShhuMWDFfpbzNSARNW23XTCSn0fPHOm5ks2+qA4
WLQXNuaJg1hVS6f7Hin3pL+zrc+Cip0KK5Mz7u8a6Lip1Ulu/tVPgPCtbrrDcpji
Xf9Tj+T/bfeHlFloE2kVawkDeN+Ts2jRtmBSu6hWi3USwXbgX06oKl6131CGPfJ/
fEGxUz0+ohSRKKEBacad4y/woRUP4VuunHFr7ZsF9j4qMufJ+RyFLs07hWMGOYC8
SCdzu+vzgfLAleXMvkmq8QTsLTJqs09n9hQSICueLaBVuumqdKZXGI6PFv6rz366
co9nxKNjETtNF6hI+Py58qOz/uENIwyoqBWi8GiGGPS7Y303UpA+CEBG31urJgDv
e6pfT2hyz6vs2Tqs5PWaC4w2T98skSUkJIYNGS+dKZ1UITchDMVuI66WkjbKEfRG
CxRIg6qb9HRWvW1yjxxtQ5U2tN4waI9u0fKM/gtRCfWfXXBBLjS7bGR5cFBoDhNu
tAtoAB48OPdJwMKF20RY7tBkKoWinDU79ZldztUVl+aLKlYV314iOBoumY2cPEj2
yys+HBh6de/IjsNqWpjsLaDdtCGBHYq+OF2zydZ7mYFFYKoccGTERuWfWL27T6Q9
YLm+RTgJG/uTC8rX2nvBCcODY+OCJbWz2D67wdIENM2Cy6iGI/E62HS9JVmckRua
cm6NoO67x5bDXjmaVdbjGuvKzBxJw9XHpkKCzLZ5NLOAuLNF0awjt9tz6CUhTd6r
1OtMLwHnK4kYG0IrB8AR+NPSseMUQmtAELm7Ln26n6nzhvRRQ9tk9mV0JpAgB2bC
brpWvc951S/jg1qaI83YxDrQ8YE6409MgDXyL3MHdwKKFYxb5ggCf7nH4rJaV5/b
i/A99ya7812lpnHiOS69WUEQ9xVZ7d5EIRG8gA/ST/qcHQpdzX1rsJN6NYzlMPaE
gYs36adwRmeifKJEL3s3enV2EaE1sbMJ+mcpVjRLJyJJwD57N9O4Jcvn62tjooGy
sYeWvC+aRKH7fTSbHpbsXGuvr2vOX/BF4cMqQquw2UECp3Ajnc5fMljLdQr70iXA
L586CitRjllA7/1aHKS7YLPty/zne6bRIi/fxAkRfE1f1FNA89NW4s1JHycJ7In4
IyLm7mr5ekelG/NRbI8Bvc4YXbDxTgI6sUfEMkoxF96Xy9rj/KcFVH61JkscT5sP
TNlIxVz6elaxhfrUM86TL7nZFM6ajZR5+P1MbIpyOI9pzbiqFefLkOUQmBPkZHO1
1yOEGqAAi2I8skRE7tDVIAfCOmzNIN80PHjrzvf/8mRgCHtrDaq8lPwB7gYZ3s46
Of6Ct5BqwD3RRQHArsCzioVKpkaLBDt3UsjoEWeQSvuDS9XraedK2xLGm2tmkD0t
GrDDg/JwyuFU13JhVxtjCxC7UOja7BwzlM40850uvD1EPWU87NWRcT/PpwYj8ltN
jtUaHL4w7fUKvE6bxqtGT60wOovPbjCKc2LSz2EreLZ/vFKICRv+RHJx0F4AQPYl
Qhu8bBScNh5hpVzMgcJHTDIAhtolZsDmBKd2ccjqLTqk/OVTHoeR5y20lJqQawF4
DSkkG7lx2cNMflGJcjL3ipQUGZnags4hIktO6V7Tt3rIZlpV4HtrrsexCkliCtkH
yqXDnoYwSHDVe+qsaLhfXwk7fdHIRiQd31sQ/atpZGd+2/eXU4Yw3OnQE37ytRRO
0kYqnKjtMOyUsKaSGpKeTgVCITU/qUCIx6hS5gsqPh2cV9SiQ6nKgpDcuXO2xMvR
+Jwkf6xHmr7IghbOw4S2NmbkBa8ebQH24XRBlr7fCFXe1lAU7vhdWTYhujxsK9RG
pUUyMFPjnIEtRz0EdRDy368RzeIKox/AXNovZnkMtuxudZUKR359fMPGkZ/57aAe
1SFPVF1m9x7u4UxmnWxpXYo0yy4Ls6c18THnIdB6l+ascAiBgd7uBbEtFA+G3t5n
GElZPIUCSgMV/FW8W9lxc0aHjSwLem5rLvh2WtO7RFzqR7wPoOziJQTwtI0pe7ly
4T4PCnRI9OhpHy9rcf5mYh0NLyzj3//I9kZVgqr+RRDlTLcac907gcihPFhO+VjL
jUuyVdO5vEdt1KnVbFUUi2To1FfguJZPtC5TwcMNn7tZ1NAOT1h+UcqwhyidKAec
e/y+ANLlOpRNBwnW9RVs9kn2or8q8PGDAZE++mi8J2Jv99WGF8c45SsJgMQVPIBr
qi8k0Vg5I3jhvgyefgSrJtj74PEFsG8CUA9eoBVaIjYjGMdQu6KS0uMjevj0N74k
t0+FRsCNsoJlPvVGIFTWOco9EXiZe2TJequnxE8eOrrRPUChWyfPPt3HcFDM/cuX
a1TqJNG+gQibD8KVLe23s3D2P4nq7hn1HRJf0S6n/VC0P7sUc/1skrDil0ycbKnX
/MTmmlCdEiJEy7T6mwpCchLmOZ3XfhyuYy5iNXyvvUg=
`protect END_PROTECTED
