`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHH8qDnf4eTvHJs7O3WzMSU+2ok30vTEe5t7557yq2GauGNUwdHwlz1G68vHNqDg
ObZ81W8EG3+Pc8YnqP4cXIuNGBpVVv3507bepSH/iuVR2ZBpmrgNx6ukobBQKuey
C9bUfceTI1NdZ2RP/bfZIeSlIACybagXiLa5mtZCveejrvPkoz+fHfFArKFNrMdx
fkFHkX2A13So9On63RTWxp6loEluLdM8R1RHuqvvpi8wgYYQ6JhWGfhZHgmkZYUH
SHO0KgkyC49m6g2F0SG/jKPbiOCR6OiwoPVl1cmN7hbZ3nlmMKM6tL0+goq/qaLg
xnJLShUPRMudaJXQGhcRaepqv6m1VC1YEn0VNyUIxboZG885BFN/2n4lEylVr8Tp
BcGjZ4sVTve2ITAGytAVhhqjWxR6ZHOte2/1nYvosOXocIsO3CBTfXUlukDi8X2n
OJNuOvvyRSuq9OggrWgeeWNNj5Do1htUFl6IUpcAQlYZ3e7AZSxkj5twbYXe+n0J
yAPyIcCTVp7UEkL08mTzMKrL6VTCZayUXQhNGcGsqnKpM12c1z1+s7xXqtPD4tQ0
p8ezKIwVJZoQk7Oij7hcx6GOppRGq3DzRFjWCeiGuzbwvNzWtMVV55u4k76Jf2Q6
DhFGYhPCA2qXtAgj8T/9OMfUf7kYy3UEJ3tWL47UYZPZcghUD8ARytsQUhB5quDg
v+uQgFyqE/YRXKL3i/kvRYVR0P+h6jYjTfYdqd15fFK5dV+ZLwMsXQQsHZ0lRJx5
X4GjyTIGXqBaEMxH2Dm7iJU28eHmEUUFIYn+y7RnjPcVoIx5LLYsC8t9gkNRaIHB
ZLVfgIGn/D7ixNaqkJURlWeTbO7lOrrmN13uSAShOLCplyTXJr4AC//DHasU5dKU
O0q1t6d/chqarzHNPsb/38B5IraESU8Th+PeX9oVwMOIt6J25EUeQg0YEUlf/gPY
KpPEEEJZU3H5PLSMiE/WQVFHUN8dGOYZQEoyElzzMKHYdNZDLLCWdiCHe0BCEuF0
0OWjtl7votT31j8N3e2uZHGttFDvtrf+jJ+ezQf6czYoa5dcZ/HUVcj2hu5eM6Nw
`protect END_PROTECTED
