`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmBxXwRkJUFP+LNMlMlzeZeSvFGR20TsRJSsXUmFhdWfwA0bkx2TpHpn3BBOMoGR
6O77ERn1zCvv/auBEe5Yf5CGEey7DNoTIKkfFAlPfE7iQJ5IPHmvGZA4OtVrbjlb
jRwTxG88daoly3Cl8pAFZhZOa9XGs9OmgH5wlDkggczaFCfZ5xgB3l8n91qo/ng8
21BRn2ToQ89wZbKI44tUILjZ0RnfkKwr30TuWca5yGn4P3oLbAFAweKYrYzbsZOt
F9GmJOkwrR7YMtkUQfihk2c10ocC6LBQfQR83tiQqRnp8+6+zVVxSgIgKaFAG0vQ
FnUKNxhuWS1rTWqxi+Ow8K17duRQhSmpZVQg5vv29y6Wi7gthi8lTHs9awL+Otp9
iPKGYTg9SKg9D3olMTcrs+sw+YJS4MQNu9yh4oCYiGWjBABGab1fXMqT8ufVY/Ee
5UkH75sbWRoUp5zbndpdYZsZTydjcjxuQXkCTTOptcaxM6rwfwAnvr57EyBCHVAc
87cEwrDojuIJadHjMaQtQWNImbQ0ReZOXlJHLsSXE17cy2ei1bs4hVkoHBquL1My
wpWPQMI2P5aWdPH0KcqomAWR30DAL/zbIRDGC2x148Y2g0O9YeHaIiKminZctJd/
HZgt4yv2/Exs18AtdfvXDvluLEcy5jqEROBrE/nDmUxoZ4kHJkC2IvvT7AfQLom4
R2R/BGkEWAHDKYDtn8c+Ex4VJTDvDfB3u3+v3nsNw5ay+Z5TaShK3DIf37QOCgRs
F85i7yI6UHq6p7hFFwmzV0s5s2iqn9XBdFo8aEMGWVq4XipDIEHCuHogGftnlqF6
krYbqdj9ADDUP7Uds2XiK2coC2cKNbYhNy0ebfwdwgXKl5Ma1/JiRw/u8N/wPRsQ
a5VmAEXnE2o1pB+6rrkuNEbfG7k9Ae0LtMHXYjXMcUJ7qDZr/qUoONhNy/1lob4P
6iS+Wq0rlBU7Rld09v3T4GCLsHzG/BmWyZIYCaFBwdfxbAD0bXmmQnwmgqbrMXUR
1nllaeg4U324eE8a23EfSqHmD3yLNvMdf4DJ25fPJ1ARge6pSC+WlJFbs5JJIct7
zU7ZiEc06UGwQze9bg0JpSnyq3dDuMjYGyXf1VXb/Ad1nd4cKYrVheEmiVR1qic2
eF5Y1V8JJrR3jmzZOVR4WExLs65ie8BEMp5xdAq9YxB2uQioOe184JNhScw7Vmxt
acfyKfV/OTzN+x2AGcqDb76KwuKyn1G5PSGhwYS6/EkQj4cEV5BOhrTf0oUvYW5u
m40aXeoNI/lL2q1pNuN5oLxDwIQyMtCCWTgJYMVtxTyq3L3CFjh8o0v1XaRJXC+a
Cz5cHm4qV3p0iLxxrUbYlAvDe7+7fIGSPEOvSp4QqCwyam5Hzk19MkPSB8umhUJC
zT4qDvvIVtRMLkNbwY4YClM3vEDlc28xsfYYpP2NVq7l/kf1MInDzbGrTjBNwb2F
Yr5TVrPyTjpbdMNdSJIXNvuNWdaFWNKvy8aNL0bolbyR8XD3luzm5wqeACJwEtaD
F2uyMEpxMO9RvYfc0qyw0mg5OMuMAOitFA/QaAIkBthwh4QiVYaqGWbX7lRSYcE3
moGXbmxyeH9zIJTVKYqVzvjHKvk53zmyYDRAdE2ofj3+fE1nZW546/etTw0XswAK
la57NDOqGOd/KogATn/nN5zkfGiODYmJ4BCKwTTGObhHTTikdgw011D4b83XIzHh
P7sD9r48Gcu+t1wLT/YFJXS7Ea/4K2e2+wilFseYkZAZKTDxjEmz3EtrXJOJDxMt
DdcyhEVDzqTrqX0BclC5WeNcJWKgH5SJkddVcKUow6EIMC5LM0XkezXXZclZVFrz
`protect END_PROTECTED
