`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjbqTzTQBit63RI7IotGHdXFbVUlYPPlDNJRJEbu/pBByHM11XIqilSsyQZrb7fD
o9NBmsdbctlBnOhIctWmlQ6ijZogz4Vq2wC7CNaiFMQOiQnETQ7B+/5HPWsdx69E
+fuSVgcgHG70VJRW6ioqVJkm9qQMQxfODNh8JKKyRw31u69fYgHZeqKpBjBNv3Ky
ujzCka3koxTgCYdepfRidpU4LH8ARCC6qhINA6c2JWXwbwrl4cSV9ChRp83wyBKA
DwGNVJ4JLvq6YnnRbUfQs8XFKR9ut8lK0ELe4Z29+Qp2f3DQ1mfvmcX2IM8IWlmk
3X8DA6FMgfVOzVfAIf3SuA==
`protect END_PROTECTED
