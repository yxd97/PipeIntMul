`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5veIIJNXRZyW334zu2+R5w2NMnK+VURC/lvHa9vL/35M5Mkaw7AmAqF8P1ORWgs
X0r1XGnxLmJphoHx5HagAeJt9yK4n7ckt3W5Zqc4t74Bw8sg+y1S1kqGIy39k578
724LpTbblDa16YOygv00Kn2+paEW+b5mtHO5yaa00bn4c7+MwHMramWwKOSk38sD
YUSRtdcQ94GKcIx9PtHS9o+01b6KhvgwelRRrIXl1+xvWIbOib+Lgasv+Z2nG6Xi
gfpQzAE3hFiNfodm26B7HMecEPmKnID1AXLtrwwwg7qLB6cI3ykguOn63UhNyLaX
KLDqB0LvyJb0xhCo6W8p8REU2TWasSIx7NDiLRCkUz8IWV8NqaSiWeWJkVwYPFY0
gMWwQJduIN0W7urxTna2A+Nsx86sOK1/acH2UlOIODYQQU+DriTTXJawsGoMxCEf
HP/0bGK4l1KSAPyFE9wTm+zLBDwafDbe+jDFj2APCfvLDD0Tm+mLyaHtZUmc+47i
fA1qycoyJRddYbEONWB9uG4RTUg+Ak/Ub6mBkDl246cfmWZZsdEjJczUio/1dpDs
pIj05QtD5j7Jj39H/pDZ/6GO1ik+ayYdKmITExAJWgMe8W9DODEpcB7rGQ7Lkcfy
sQHK3MZEeCRgg6uF3fy4a1Xvsq7fk2gyrcKdDYCCm8aJIA2V/e0anTgRGGY8jYHK
Be7YOqq+758LQ3oISk5IwbW148nITCm9jzMrK7a9mEk8hrLuTZUn7jyQ0aIQ66/S
g5kLNX1279LOBqf8u2QGIYoSzu0c08CO0osI53ACFZ/ICP6tc/gnHebJKGY62J5n
9cfMUk1tcHXEFsLESBTBjdZSA+/H7JXFMWtKbzmRA4+9OkkNqfYGMy9s9hxim0R0
ggJAmcg87krFBtKraYPHAMbek4s9TIFeUyqeJzYKGLrciQyS/yKc8OU7sLsLTbZk
FYuOJLebOEz/Ui6GGd5FmQPdWGfcD0yENuYorpUwv4vWRNs8s5VBFjJQTwaIW8tE
QqngegyNWBr37wv/uEOoXDAWARm3qV/y1MXlD6AuN1L5ADFn7Qi1hoAA9fEYKBuf
cwcVwfgEtUKS3lVfxRGsXaGzCpNPvDOz+OS71/hcIBmZLlxNtpZqqEIcgEMo/Eoi
j65A6F04FblIgSWEObFWrXIZOD+oJLkKjN8GL56XrJEbkOh1uCITb0dm2c9kARZw
77flBmIBeacq47/uTGx9RSAgXMRiOftNwVmt7vIxyj7gC5say7ICP1nQZ0ytP4yw
3UG73vSAimD1KbBUpKCZi+FZwhwBABpqm5qtauk57feF9jx5YDidPsB+/V4TPTSV
JqO6hTodz9QNhy+6V6eQ9A==
`protect END_PROTECTED
