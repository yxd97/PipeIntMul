`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQoQSUa3nI4WznSH7n3uCb6x1STHghDeS7p/Xdh5t3tZB64GBtDtrVlNWYsrr1V2
VP2TJXzR1YiWurDfYcTDdWhJiV2z3NsdDO7urVlUjKP/FAvj+oBlq72iFmUzShsD
Uo1roMzp+TsT1wNXX8sgI1FL9k+rOaPXGljU3oYukGWAdpApQVJPQGRDTpxxajDu
YzxcpPBy12HtYl3XDFfU/UDApW3RP5UDPIDGgROu09GeVpOVxRbqnfzBnKMRz0q/
3crbWxryTkCdXUimDlyiL9MiQYGgZDhYW9OG8Yfyuij6lqUCgPgjYCzkdG5yXcQA
n/AxKHdim4jiB/3kingrIcrQ8hmNPm04CP4Y2IcUMVnNCpEkx5WfTyc4lTDHkaAg
InbI/J4lijOWRD37evgE3flKJu/erl0ztAnfQhMFKNRwFImR6DEDaXJkMTCj+EFL
/tbiEmJrrbpXkvT9n7wEfSYXgyIi6PdUCnbDnNEjqMOoGYr+NssvKWjuW3oxw9fO
7uRbaCbMQ5BTcoL/RKcIQ/sEuse6Ez6pgJjzpfgamwftiOYPRVV2r3bpG0iF8ylw
oy2o8aGO1wvy91JGQUmXFRrQQx2UaN11dqzKUY/LZzn01+yORAWmJAgLYQuY/1z4
7menCuAKPNgLWiFejcoykUbuma1mqn4N3oIY6nFibCcZ0xT0cVPZ4W4kbhsNWEdX
aHqeByTLqzJuNgoJoTY7tql9Ji4HKHxyMZZTdFGv/OU=
`protect END_PROTECTED
