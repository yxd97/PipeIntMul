`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYlH7nmavixcWEgXeaVayJjHx5N0sssyYRDz+Fe9ki41k2vvBvEjT6htRrgnMEpr
bO8k5ZM1QsbJnm4SuDe8DEEVX+T4imp1UIFnWZYY3bWi7iD6VsjbT6INNFwSE4E3
kFptMPHFg0zXFUJ4q2JD3hT1TWxtUY8yT9h/IUxOQDI8YTBrIi/opt1i1tFzOlVo
lTGZu8wnV8NesiQdlzwEU0NKrvTRjsx9CndaR1BqS2A74+zuJQkSsQ84TWhemB9t
ctAM8PFjVeIg3ht/gXuZU1azQ+2GfFw62bj8fuOvO1Js0vU13xM1+/hTEZj0I4vP
CiU0EUnKROEuVzrplCq9JCxv8ZJYXkZeEzm6QMIGfpx6Tx2ZS5Y3k0mon6XpE0si
ZYUDcldSH/o5CLl/ahD6TqcOOf57C8URhzgVkJfaZJLyRpj2Q0DR7jRVAIvyzxd5
Av5w/sD29gvgRutccJn41MKZU/gNbxwkEKHggg5Q2iKGBZMfu7itcwqJ6izjhgMe
3OcpodV3hCGQ5j7kXG5iVBYtA9pwBODsOcSzOAKc8iA+L32MkHU5I0n/zTR7mWea
D3CnGi0p6UDKXF+E9gis6d+A89gr3SkhL13hT0mbvcdyvzxboROGV/4K/IwJQQ1i
xJOfY9XVn9M13JFntcOCJg==
`protect END_PROTECTED
