`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jq8otpCzHIlkiiVA0s9bwsX1K9jcbMzRm+HZQRjiSn7x1SbpIRudddRcAwvsMQbk
beaSBEdhf+Nh3UnkzYU9VFq86jY9xV4MFBc40h2ZExB+N/Fub0zUI+PpkcQSX7Xe
AHyEixoWDPXTVzEOkh0mrwVI9gLD8yvhQKC1QF0kfS2wXjgwn6lDHKmyVQmUAt6o
9Jkg8dGQjlqIXAlA7JUhTFjGX5bCMuSC5UMhYSDGmwMs7pUY0vUs268ylim3z4KT
prPOPsRKvHTtAPnk6mhdoQ==
`protect END_PROTECTED
