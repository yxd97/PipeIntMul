`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YhdxaEsh+3eDAJr14o6ccFkKabaTp9W0Rd8SX5uU68dDIzHTArANcJSb253Sn06D
55Kx6rFbNxZcmzOghp117NKAu0q3R6tA/XeelpOgMKHHKwbYh5Zx/bLYrdEGnl51
9dji9JtExg6VTDJRA9b3bJlRS28yfu/e86zQPOZKMz2BhA8INBZ1MGYFbESbq6qE
4B6ihfD5BrxuLNrbXmvGxnnZFBVfPHpNurQQU9UY9Rmqnnf31Emx1zKURyBcvE9Z
QnOQRUe9NP3hXlZYqAM0WP2FnIq/igfwPcKHliBPDu2QZKZlZrLfy337ptg/UiCJ
8YqeYniwZKll1ofyCeGKConhuOeB+6dHhLO+esJ1Ba4QCsDn6ezgHxobyV8Jvb9e
4dmYNPSotQMdizLi3C2w9wsAz5k3YlXlqxWqoARD19N7lYU9jS4rSRPm+orUkOke
wh82v6NdZ3eh1LNeDf0uolUBwt3WM90l/mXvu+Qz391Kk3GMb9Z0aH8PKFxlkKr+
mtRy36i1DTNvgilLYd3EvjyskWUGkHvd5emM4AF2PncmgaScbJdJYG0qVnmv7ruN
`protect END_PROTECTED
