`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kYKiwUcUcYMyCSY71Cq+dWIpd7BUQ+fcctaJBfap58JATfGPRiXUbpxdD1Y7RAcL
qsdlv5EDSOCbgVtvpCd6jbAqDmI8TzsmpLVP1SXg4I1uVX66jUzec6qwNMA9+UDH
eB0jnchezW1mW6VZYzVrrrI+ZodhVHO8ErwizHika/VvjXkpPJrpB8F/hApY0xHf
GEiVbk54uzbtVByd1HSF/3r7UtsVo6e6Mbwattd6DfbmE1abJsipwNv/j9jRcVKL
UjlnXxKDd1fIyTc2jEH7X3vo2KCeCn5DH0uP0ryPixuEdfRU12ySIa5CiRjOAIHx
bQ9K0HmKcG4pdc4VjtWH1w25IbrKHoMP8ar6u7z+WrpL/ekK7u3KyzH2tmFG0F1w
`protect END_PROTECTED
