`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iwy8SrgkaLxvM094DKLCvd9QGrh5Nz6fHn3McWy/M6AVy9iOJ+M9r1F7W5sVA8bP
BWTMwuYvkfqm99QHiuWuQrn/JgH9V5s6Y1CwXxpapyl63b/I5HHPOIzfDKvuuk2I
UlJF65Uw2JC7AHl2hNRpdSsb01ezkiqKIAjVczvMDE0vGSrNXzVkFJ1ZiehCBZ/r
yRhMmH5+539+ZAMmu9ZdQdZPiYlziJX0urePpLBUyb2sDSZq2zGsrNq1VaC1plLH
Y5D6S+4Zs8s0cZAewx6hw0/QTC4e0ZEPupKCP3eMSNSGBAnUy32z0h/zIY/Z+/Oe
G5uyqq2B9roCxzI1oJ9fO9IXaMoOMDlFBrNwyWqpcQBu7/wxkfuKHkIXbHUJxw3L
zELsbRAWif0OirMU9xS3Dw/2vAuJ56fBCSnNn3PNwcXLQMCotB9eH2GtBYnk/jl9
kLmwQrRCK29MR/7jzybthio0O6g7o5K+uieeHy98sEhoYZ2nAuNIew6Ocvpf9t9l
tN4hWOch8c1MDZzc2uyi6sxcGHDYViTFy5bGV6z/eGQZM9s6tqoNGlrKkNeQp75G
DA8RMO/uhAAZAUDGR74XCxiKbdq0PcKKPz5yzRiSeAyM5SxmQcbjVGKKD7SiaEgH
R3AIcqnVubWZl7rwDd5obXjjj70QGHYB1a73l4mJNqIfB79Y/dQTHcTlWeZQmFBY
pSr5dY+Fe90e8kdKDVfsSNiQByflQgezrTdRcUpBBvlLH1KIrta5l0FEJ4F1q/f1
2OJKqXfSZUUL1+6ozpYfE9ln7WNhFSF1PcSnJVap8BVbeZdT4HM38lUV5N7cY0Sv
De6x4zCp7prbeXohThdd4b1eVviLznlO6Df+uI8zEK8F8LVSEOyVvnDWGamGaJI6
M3+uB00z7BEhxd02wL11oCPVvyoy12f+xQaSsqtb+PptBiA9ldZ4oepd7s6vlLXl
`protect END_PROTECTED
