`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBvUypk04jLdr9LHpyXa3Jn0NGKAFeA1QM46iuLtTSJlT1GL3L2T5hW/lVhaFut6
GqHPJumRNwHt4STaJTQBUia6QATxUpBcxPPoa4M7qGF3AOaN9KiuX1cmERL0NPcU
thdREPgVarpqOtPE08l+c7x+Lyyyza5RBmxEtZGQJkoYukRTPiDf1+T5o0YVSEw5
oX4hLRwugEjDMMkgwjG5yCT2pA7T1P9u7ds44jLxvQN2+nLlO0x/p6Oi7updIyfi
PqOBMWtxE5A0S28oh3dXLyYoJrH8Q1gA2qhBwv5ZnhH+g/Sr67GIRqpJ27kD8DG3
mMvShPX1CqHSIYJdZ8qazzj2TihCzuQGF98xfazIQooxO/pChfySK0G++WmwXrR+
RgBw94z7AUJcWARzdYg5B7FRGm2wE2djcTSlvoz99nP4iUCAJasREDNsWqQU2GeG
+YUhZgJMs/yZQqRIKbywV6102ClOdqjQzxLBfZgXhUY/9gl9R/WvkQft97Ntd9iH
1madfOrLjjWZhiia3LXlY8hOooYVBk/woyGXmGbp/TY/38JL98F4PKQIGDRjJFnk
LrKbfe0v0GXhidiKR4ZUOcvYrWd5NiEb7ZHJcK94xrNocTdRHlKuUnGL3HNB1KOm
O3b8k7Z8vBT160BFRdb0tNDbMbXMFrf1TCyUX2gdYlg=
`protect END_PROTECTED
