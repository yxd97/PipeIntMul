`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqGnSOw9e/BJlE8dc8LIrS9KJSqMo29IDPHQ7nH3ExquQRcwzhrq9xDO/XEuou9y
4/bjTP88zx9EmVQDek00oDvHcgakqrg04OQg8E4RtKxYlPkBXA0U6mS6MikTqdGu
rySbSopHSHbjFS/DqBn5/56weQHXYl89sJWm64ygKhmxlQ4cCKzgndCkCERf0sxd
DTos8QjwMKbUSOMlzAqfb6hGpLxqcr2ZeVyOBmRDZKa4jNQz20Hv0pKFzZtUqFHK
WWIvHNMpKYBoUAzj18RMW8PaL8npOSRvL+41+7SmLsNUk7Z7t2fx5HJuJoQ3tN87
GUIHid7tvuOm32DTrEJAw0b987f6PAPlNPfDKtf0Y2lnYw+yvqQ1Sacyvg4o2eG1
XqHoqsxqlQD3jBuZDsDiYgd0ZRz1QnWlLuScWEC8NaOFCgJvGogKb20Y9mj5kf/d
iloIcyXFT5zthwi4gnCHDGM4XTyOqdAEDDHgFNJMszpUUP27Lx5AEXGkDh9YVi+G
0L4Qs94ykyvZ2AOdS/cr+E8qL03pQMvU4KoPl6xc2JQhGmAF620ZKJJ92I+L/sbw
HyIxcdRH+eeZ7csgL+b/e0xDSO3ZJDzjf8V/Qhs2zQkayttLgBCJCYJGVx2irf7V
`protect END_PROTECTED
