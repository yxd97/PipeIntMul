`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
znfakUI9UWPgOtS5bwYnl/h6MJ8xzHHpPSzzLwqP1DawV2ZnS1o1IYJep0bEJDIL
f9X7YqnH/T2ZfaHlkmbeCIX5TYOWTj7mg1KmitIVRHakcSHO5zl6bOIaYOJpTYJU
RYNRaS2I/7FL/9jg37XZTTVIYd0ETne6UUmKb84qiIJqxrXQbgMaZsHUfkHVXulQ
dCC9rL73WA+ks7hGIX2pjhT2r8qolKeYOhdSQ+hnBJFlDCvF9zAS8l4PtnJHGSyF
GAr/aDFGJ/xafLN7dtbqTemjd/VF3qoLCqrbyb+ER6RhKk46eRTW9UE5qnPFNMym
PiT5TJxb8xtLKS3EN66eGAeTYYY/1OJO/6Txt10sh2/kDUFL2uWrSJHxThRMMb5x
QmRk+iVZyYVPnJpu3YmY8w==
`protect END_PROTECTED
