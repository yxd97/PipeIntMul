`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sBvIw0rIBEF9FHM2mqlbkPuZHf4OTwM2tghO+fgy4jL3PoZSnHCRtMNfSswY21j6
HJgXPc/Cw1AYVYNRs0bPlSlVqOWJMApiIXqivYsZjeLu1uWyZV4Sos9AdXJMSXEp
4OilZCXbGQwezmGJbnfnqe+d9cCa6wQhahaheJiVkPT5mtdZ8X5gDtbVcpCIUMX4
cg78a6eLN1Ua5tbzjEM+vzPrcJ8ReOp8D3M5ItgepyPBOsy6t4/+jo0+CzW4KQ+m
PzNW5UnrSHWx9Q5CBV9/kEVjG13Ye/baj21lk4Q7PCdHi4s/2k0x3o+u2EGHEn1s
OrNr8Qli/rUOUzi+QQMIMA0LGBj2Evs++A/Mw+/ELWoyaOsx0MOPM0+RHmDaW2ZD
EHq3L2vmssqfqSZWZXgkgGqEr5mWx3sYsHRBrt+8lGvQPeAp4GHWZvdWWVVhFF+r
bbNHgHOU5aanJLE7bulXWXVCqPhW8Ba3fAQ9up6G2X2ncXLD3WFfp3TbYKOWZu0k
B32RQWiQu1MMuCxBQg85B0y3aWrZoFrZjCH8YnV/XZiQ+bOHMYXaObdaqQX4tRtP
2eAgR9gQKQ4qNy4RkihgUIj4fjc4qZwhSDF+k+DGccylJSGUxSy1c9IoFogkRz+7
Ju8rzRkCH8wrf9kRbraxqaZd7JmXn6iUDPZVxiY2O4AvKxc8ynI3VPN6H6Lgxl4l
idl3w6PuXE0BBZ7r+bwqlCherUJVTgJCRk+AoSt37GWqOctHIttLYnJ1S6lu81pn
UzbtH8y2CpceQjRgeoxL2VptB7lQmUKAXHt3bJX0XfJCNaGmakfLaqODWxzogLFh
6sZTLxqaalVf1GY0kDutPMK3C+AaHP5bL9Tg6BcmfBFmuACrhbr5tLDVcwVkwj3B
i9kTEUTj53zjPeSBLQiFFDHDlzt3YpoEQY1OJm0fSSUDwylq+w/7i7KzmPbENsBJ
V+VejDsv1PXJ356j+OsyP+ZplcXbWdFTXhj40glXP+7UY/2jZJ9yy2NWZP2i4AcN
PqVQuzcG3cB6iJR1humiR5qqzbBng+OsVuh22vWsiOhq3a89jdc84GVVkkz/PAxk
LkPWMLMMKO6q5cRTOxM0wCO4JC8d3JtB4PyuioNGsCCudOZ4KEwIQtYjcLozuMlw
LA6y02/twUJrXo3ooIslqSFu1afM8LCZJB0RHElThbfUkFTOp1p+IUiSeB4eSBdm
0OkpaC31FguIHLnSlzoBYBimACHa/zzbIsMbYXTqhsd7uuTcrKSQSePxUpt5BoWZ
QiZApzcaaAmzxv/KqqR4n7Davy+eMOaz88eFtxQqGuCtfkGxvd0eIW6Ic2uZ4lAE
PsKNppSoOqwFTBA26hBRSpPFfwnz8Xn7V3AcoLLoZW6TwlEDb9anQglzB+bW2GdJ
7ZQ2aNOJsmnwgAfat/8E5TZS7tJe3bOwGOegz1E+ngkwOXvv/kInbB0cvjvE2Cgg
7H4xec5AOXneKCL5dBNuM/NIawol7k0OQc63dhh3nrGiAZ51v+fALLTJYkgbU6QM
gKGHZwkjASKaA/7ARM7KVHQf+dl83e3Me6dZhhjErqCQKEKIFGWpX/ypBkQLVEHl
8K5jVdkxaMGrpLDxba5hupr2Bc2/yh8X6lNwKH+9jTAgGX0W+WRFk0PpKgr2bFf6
JqDnZdC1Gpt5FwQe7nT8gSJySBRBD1xLx7pkgXQCGOMtIfC9XNGP0cDAgqBRJzzj
pmmsuroM6hq2j27v9GcVSHlonOM4WIDVD2SKUX4cnTsUVNR++rfGcWdS7L0iVoiK
8Pmu83xbywQFKhVnMIdn0NPOSo/eE0wmUiu416bVvuomq6ljq3G7W9ahaHESh5j7
1WmKf/9/hzABaf7yMxhTwVALMrc6h+LWomTdzrUVZtkSXCUtGVSg7TNmEuv0Juy0
Vh80R/8zCsJy34TDFVPX5LzUq4dwHf+VQldG4QMuOcJYOCOyUxvReENTN7YNONF6
IN8l7Eiu/A3grJRBV6F757F1VIQEF4D+zfv7wegxf4xIvFC6UNXCDXjzp/Y7UTXd
04xb+kEm/LUZMvlE5km6RiaHl5iQv9v/RWUTEhijhWMFbWq7o3pJ0Yhag2HXIiqt
LYDQgSVYzX6/8foKD6HkG+BRkpz9bZAcXL8eGsTS3SmsXTv/EPCbCNiRUdpLQHfi
3uyTifMkvG8zRYl1FS+RsAVRQOl1Y78noaipzi/6afjixGf6Qms0tJsVF7YgRA/I
Sv7+tEBpIHc11dX7LbFJaAV3T7JB2mIGNguRRM1Vd9lKn2SDDSFmdnLsoEVBEF+L
77+G8QK0Zi8+2hPlnDqc/L6tiqZm7h9ObNtbQ80qySyiZwRJ1YOOhEGYtjNSaRLq
D8vASMt8K2WsNbaO+uuRPiVMHf2zojGBRA+ZLP/iMmMxKwheI7MHtu+4vgZ8Vd/6
P0/AzZucjB7jCJ7lZKd6z7R8OTZepVPMQp0Bow29rhy9eEdfW9Dj+GIkA9ox8g/W
k+wLZx1m/e7WLAIQ3p+rEAzDUA/xdxLf1+ISxogLC/lrEw6XGGCB43IMdfE3cKhG
`protect END_PROTECTED
