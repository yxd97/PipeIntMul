`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxMsYa72j4/W2OY6zeGAXg5Kr9zgpeRPNVkWPrumfFVbNSh8+8KdukBMbEEVkTOd
gL8BBxhlc3mj8g72ubbqYUpR2Xp/19pHH7OVk5hPGYgVgwgxf863a3m8hET4ToDg
590BbH7i7SFuIUbOaQ36wB/lXdvmRoQYyRPqGjevCv8tvpDOpspMDNWZrXiahjK0
gKpuxjb8GqvGWQo2SbwmSYVAKYXQD5LLwpSFCMtyICgjmF2/ONZGplMWQJiAPFZP
6Gb7FL98lsNRRQQl5JJPafWcwJ/g7GLKdDmTJ1EMq/uUvc6yCOm8kzFFTAEeTYEA
G3flqAuW4Si6+mGvI5Ma20jSNHaZJ8BQ1DUOVSfb9ZAl1GgdJxGwxMDEI7utT710
kStvaCbscI445qnAGINskwBYg7DlA20g3kfQjjhTtwY=
`protect END_PROTECTED
