`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+j3FrimAZjzBV/Q9FTM2gERGnFNh3Tj8WfXEEanb5ehNH8KPX7ME3WjPIdFlOQL7
L5zqJ/iOGGuUhEgZNiIlmoFTtOlQ/JsLgDP+wVUC/CzBLiM72lkZwK5Isujyg35b
oq0VhA0vNzwsf0DGAsZ+DllJmkoUw2iARiFpEiOgg61PH5HuwH7SKlV/gVoGR657
dxa45PaPZD2V8wxDEjVY8vvxN//kB7QlsK0XHconbQxU9NXddy1e3XuLWVa/Zbwd
iLqQ3reZoU+XPrjg1Xwh2sSkuDeG0qryIzaH+hWuLkuszv29z2JplrSZe16VedFd
tiEHjeG81xANgSFc+ObQlaSfHK4+kny33r8UWzYPxGhTnKvBIcqrQ2pqJv8kA9X9
YWDKf/1bliLMPWgM6GIW/yTlAlZhvb7Hvj4rlP8DzO5J+h04S6DWuOiEuzzjuDfA
NhJGEhHQjggmXyldfCYtFjTXeSKjRLz+NugEHO/lgAXSRwGIn4YRCsIzs3DdCjTy
gLrkwGCGLadTccDt+JBkNSSlRlWLpWt4v1ImF7NIj7XyOenjfB1fk4UeYuyDaBMV
OhXG+EZm5aredkP7myBiNE2p2UEkRrtvIBbNSgfkT9rXWlooHGbRrYvxSqiAxr1R
bSGFIZKhdaNulnMRemlDBF/u2DP+imt8Symdf5qj42pAEKMAowWoAHOzU3xwCw/a
2KXh5CyccG3Rwzvzj6ouDCbKQQrHQRSRELMXBDehd4ObmHBt0rOnc3AvDvqMsAMa
6zSKbrN7eudzJuVyIL1S7eM4K/0F9RMr1nY4uFOp3V2iVgPyGawxMyRoC4WhMhk/
HXN+52AFJPJXP061Ad89SVh7MIBjrGjtFriVZVrYmf0OXU5s7Jr3TWBW13MrdeXU
eKS/0c9NdF0wQifB1054ZBkZGj4LsEqhQ9LbP2GoMwCSJgxacPl5cOlWBIY1EfXJ
LFaY1xkFZwe2bMyY5tGGx+fwkwb4/WYO0zk/RHVZXqhWeX6t4iZBMDFEan4YMxnR
a1QkFdnfPrjGn01ytukq8gpZGP6g13bpCdyDeNCOWSx5ornOW5rCCk+yKmP9WK4v
sg9xymIp6va8mTI5Fl8TAVBrSOLg+ZzvPYnVZ0oq92MKgmpGUzV9gpgyJAqf/nKR
9upVJXu9W/csJU3Wm/1DhZnC4vKpw3+ugDg4J554PA2c7O4xk9hrEVhbe9KT05SH
2FEpW+PvXld6gfi4q1zNCMkg9pDB+fP8rp+lZ6OU6pjiWvVAj40qHa/Z8WN4L/UK
zi9EyV/ivJ16B715fAn/fCSlf0S4QxVLNAca92AChmOY7WFgu2D7WLXnxVpeq0Vy
h6vVP0pi3li4d49g5fEOl61lOjY06hhjQgXb1IMPktCnG+Grwtovi4fWAW9A3YQK
Qka80TwrzYoQZk5jxuhWnAj0UQfstDbwwYnFJG5a+lvWv5UQYR4ayPoRRwGcDTp4
z2A+eCX0cx7rTihWUMeACpqJVKeLB2DT5dxbQA4ZY8yH6sTQbIByprvRWG8M40V/
Oojh7LpEby2fbDeFQ6M3277yC3tcEqXGHNy9R/X9uzPcrB98LSZjiytxVDEKWiJs
kjn4uSYH74zRuV+E4X2WDo5Cth4aAjOQY1L49keN5Asb8NBCVjW3j1BtRH58Oa1p
lk/mzBbjjQdlsYqU7OgGNFFfJX7ejokkZQ15Ixuxn1ZkSRS7llPCN4OtP/5EFCS5
J4ttI0uyLbFruGVEh7jtV673xDP/7mJ6aJvEELBkwpVLwQCp+OwtBlz5h+PsnsJW
MW3PawJSsxzpwtL5Wy5QJ7DCiYMSl93IX14PPFMkKEk=
`protect END_PROTECTED
