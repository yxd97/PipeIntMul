`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nmxi8HaJ4o0tiI1TKFi4aRCf9OjZdYNXpTMG5AF48fD4nRJ8EJNh8N1hzZziYPpZ
nM4pUCDbb/ihhKN6HBtA7lnpNUgS3RUBtwnrKlVcFOp6tGWN/dINPAS4ohMyXOJa
WJJ7/wQ+RV+TwVl0DW/rvBhBnecl4WDN+phUdm8UX9VhUK1aEEPUSvY13rE/y+Tf
pkdHYrfkrQIm/AMbiWzeb9l8fBeaKa7+BJZMfEHp9eiC3rCYpzg1YqF3BtzE3fs+
ZmjPpDdmX/7TIV96DHIt4b3K3mm9uwj6QUzpZbLnGx3rCn02QMyi75HhQkppIiJj
9ZNPrCCEdQMAQI3sT7+OWw==
`protect END_PROTECTED
