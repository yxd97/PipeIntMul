`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pc1gj8qWg9xT8ghFhWK0QFpHugSlLwIenpph+2LBLCz4T9MbFtAVGz/4XGtAfgOo
1zfqIGO3Q92kQ0xi7XOqNSBjiWLUzYinDZqdb+UWS0dtyB4cHWETb2WZMEVUytfN
nqpTdBK9mPBGH2LtGnAbv9Y4/ox03S27+xGFUYJj7sOEVXqzrb4c1Y89x/ihOo4s
ZzR9BwTvUAyNs4EAwgFm5owqF3oQY9YqooFsKHk+AR5KTKlIQM/EFMjpZYJ3nNIr
fg+PW2HZu7sL+k+yDbLws4pJzY+2+WcOJQIcfbKW1kFbyG+XRwY8ESpoeGiSXEzJ
ytTPDEp+LUs/losJo3m44ZpXcVMBxyfvwyWD0qOCHLPfHqbxROm+oEEOY+gN+SYF
TQqU0ed+LpQbRBmed4Yvb2clhZJFoddEwafY+JYKBjWCl9/ihfjoHRfx3p5ufarC
pOWZ2lurjZAFRXXvtdd5no3KE9GuzORi0N6OO+8iqFMOebBLMVaZQLqt+00GQ2rw
1i0DtN9+sjtnQnKyXurNJimt0K898+W2H6DinVDmRXyKXizGTod1kaJzMmXKnlqg
urIAAEbPTl1Y16tEY0eJW6BQ/k7PwNFwxviHrN7TwFbW+2rQ4RFwSN1ldY/UTIhx
ca0wcbX18RFRhaXEkQPTGfVnsYps8eytt/aWxkPz3bM=
`protect END_PROTECTED
