`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWKj5A09/4544eWg0UrFduldiCldz/2Nqv1b/Y3KDJ7X2IyuGqUVfjjg+gKsFYlb
WjAKXHrvw+HWDAHecD1lDOx/S2mkyKPWNLB92eKE8V/YoOKAtM23K5h5cWh1TPbc
a6CtkXczj1C3nFXCIG1UnlVXvKZqo4V93fpkZrtj8PGXmkNeuS0jp2+cXQ4uuQlD
cgxhNgSsIDSY6RYSGmrjjKOTTmpYxiLR6SR5INMvPHnVuKmbjcn6g3DlvDMvDgHg
jCV89kPZioIbSv+e/W56+mJ9D5z0OHT96lnmWCBIloJ0+2MSPh2O14ztICBUs6AN
x8kllbH0lOcIzbO+F8QtHtksfQ5XiBFd+KpMJePZ+pZqJm6Pc5NN0aqFOBp0HdFJ
6g7NTXa7z3yQFRthu9Msjb08zQpanyKK8Hz1R92T4L8aly9HiPW99FJXYquHBa2x
wVC76OcvFP6+rAtAOdWgcq6XWz3g1I/RT7GkEw8OepZiwvg9eeepIuxGIbR9saZi
71pioFGynVxJzHTKIhkJigm0WthewCylthfUMvFKmNI=
`protect END_PROTECTED
