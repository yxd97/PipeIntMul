`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohBOSGzrLHJMGccF+7DeH9eST2qcdlFlNRqrKu/xYrKlUq5xu4Lk4eCRyz5avrfW
UQM7doZ0YMAIdRf/Y/fiTuwX1PSdJ4hT7WgpY+QX3JkGsRMjvphdTOebpC+TKaz9
Oukrl/+Pq3VL+XKQ+ExxmE8T6N3KFQX2v0xvZPgESbl5L0KN2qNcqL5EErb4nZu9
ybpG8DlYhdDfCq9jQgEqI3zPa0Vqh2h2aA9krUzwCFUcJ2tAbMwxTce1291F5aNE
lh67TdZaDfOg2BiH6By4i89KfoAJttzT8ZnsJRRXE2Q1qRBsytTvRLy5kEbsqXhL
MpFR/KyCS9FP/8ADLKh9Ek3a7Qv3JYK+t1cG58r5dMWK6GIDSYk8ZfWKAd/YgtPK
odVN6qs7aK4nSxLdyYE8VOs83XX0kBG2/EkYqfK9ryqGWahQfaHwtASb87cM4YUr
TCGwyl0zdHxyfjUkbZo8dM6J82HefkIqiFKUvnmeto0lRz2WgNYG4WiSEOpgE1zt
KSXRFA+Q3p0G4Gnl8KCXweOChpI43tAQeVKMSELvwoxQj4TGIIxUFmc4Rjdb+TIc
1ZIxBL5w17OUEOLdPgWndFM2yuzwj2sfkmG3HmdSvpU=
`protect END_PROTECTED
