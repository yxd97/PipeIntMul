`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97MqG8/7QdG4wTZ7Gk1iu+aj+c7mUB6L5kvQ6x1E7RN+RUWliDgCFvFjTmXLFcKm
6NuS8WRhTRSb2+xgSeeRfm8utj9xTCPZEKUCaw4hFOHqarA9s4S331hbPzbiAxb1
HqIn4qFvZ3NlGa/TTeQ8ORAizLN9NLOv9YkqxN/8Z70QR5TDOGwR3NYOsW4dHJFS
urpx9TUdBySryLpzvOvcOnnJLNmDOZtBUbyaRtjtf/bKQuX8tg0Dty5Y5re9UFuU
965zVceLARFv5sq0eAdnIQ==
`protect END_PROTECTED
