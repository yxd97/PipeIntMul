`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eeJ0J6kSoptV8ZvwgHHYcnTjJQ3Ax5h7f0PCDtqsd7/1bXB2OjgaKVZWwmVg/m8v
zmuC5g/xa3sNiGbLZDWN8VpmG2bS1RTTFod+55m6mCApVKESQ3sUKAYuYkAcdSiV
dyGd9gC/53RLmDdkDy3T55JC+Xp++NrfyxiWKuqfCWs7CL6v9fD8DPp+7ZAeyGw4
8BnWRh1/BlmwH+oGEhyPo/UeaHms3XEw8m3KUpLRnubFdWRRxlRfPiOCUYC972Zd
BVSOITO7bq/ajf/UoN4tv86ui3pACIljn+i49aJdwIPpaaBPsPWqn7E/sK4ykjTx
e1kWY6RfEml5wjfP2gRBQqYiQMjyDzaj5giq4F8Tbji7YMXiNdD77aYo/1/8YgBG
PaOedXrgqbwp/8i5G3PZAWwwIl/l1TU5Tg0MqgQty1nEkHdHeieUcu9PNbZUwLDV
sGprSxNkSdyhzCWwghQ8ydWdzsQT9cY7uAHJ122OC7F+1toZbfjmmC1GjpL/aC2/
qzEi0W0YsOMnxQh7Dh5aih3MhGIEKTgfCoa2HJuvJVeBefIqj0k0G1ayaOOAsPBB
U+8VJ+nyZKhvtKVe2m9p+vEiOAte/A9VsoXb5GVM42FvgaLbzfAgsRiZLo0PgmA8
AEhD3hUC9esCHOrij2CLT6xbaaP1KBPj67avVhVTM3xgBay7IAXO1oWv2S/LS1+a
LkUQqz2nU56njebEuSfSc0KcZVq1Z8FUlHoobdjgfiyTE+hkMxWlTbqFKwV5MpT+
5qz3gFhtQFKdkPjRPPrhliB4kyfLJFD9nhA44g1vYmtzia7Nd0l02G3y/bGk+Son
KdtDGPQi+sZMt3sQ2flwCWCktz/K4Zbkpw06/n38DE6GPwLGBxfTcyn3xS/xgeN1
ePl0kBbmhGpsezg/EfzxMDbjiK1ISeQgoqhh7iE94nnxxJ6p2ViHeORoBKJP3y4X
CRczEmRZx/a83h3OQ/dNADU4kHDjZApe5yw+CLLp+x9arqDtMNjkHv8Dx1o2wa7o
GNryvNHtrrhZin0W7r0QOmKR3jxW0v0kPgfTKDqFhbYmSZNqqXG+vUWLNHGekS6T
K+aKTkntf1RIwNHddXCs97hOj4xKlgbMcb3qbP1RwGeIBhx7Z9xcr20YEEVZDg2T
jRwD8JklCmhwpQmZPeFeT/iqXdQParrmX+zZuBMSDoWg4tNH5DcsLJj8hWxGsED6
MYTC1X8JZbB50/vlI5FqiYM3FqNVxECk9qNGbWJe+it5Q6altvVQogzRUYUV64+T
Mgwtb52Y1wez9lhoDMP2Z+C9Tor4qVYfXAY8ZYgEVpTRgJxT4cwPnIz0KkQN9f6L
AZLaYztk62ZMxtW1K54iN0MrL2YeT4D07FsNm4fkQt+VauQLO30ScwgemdN8w55b
fd2/ZKQ9oXMiseJ0u8BBNLTqiPXHxJOYL7dDuT2AH21+qAuP6MBzmqgTTmo+amvV
gDoX3v04f4RgL/jRXaygyimyXqw1loxinyo7vDgTmTPPIJPi4S5SDZZeiCe/PJW8
EdtDTTp7jeteZtMV6mnjNyKaZ49SrkW0AfyoOeNj5hFqmeGXquuWP99WBS1UItgS
Nq0QwA/AwWjFXWUCf+nIthi41K1Is4f2CNqoXjfxPxNUNKzAiwyORAB4S4UsYMmI
yRZzo3K0eUNI2w6PYUh6k+VlFx+kG37a8yALTbmM4MPGvGyPwk/Kz7Owrvxd/KY2
cydusV4OS/hdlBGvg8n/CgnyICZuzjFOsj+qk6HoCU8s42dPmtJdhypUbjcBRI/3
ueKgZSPS8AhSfXwNoBQMM5/JFcEGdjBHA17lR1USePR4mQ45StIZ2PSk2kSWmvDg
tT4Eu4cJn8f+Znw6bR7PUvFeplBqWqVzyCY3xDlCHQmWWNjDGSUl3zg4Oc3fOzE7
Lpu4bb3QOVGhOembQgyP6vSnUFWMXzfyokzlr/pRpSw6+MYUGkKq8fSnSw1LxgJu
pX4IiJulH7lHlGqh7mVEPN5lLxozfnZXRPs69oZyfstr8++5JQdyo4osCjAdySG9
hrP+OzkeLx6N+duTyMPt+Mmc4db1SvYdvqygTYh3J/91761vRAJW0tS36ItFf6Vm
7k0i8gjZQLAEoBpMaYA07dZQAX3iLP/ZoFhu3LRy6AXg1CLm/SixnCzPU5UU1Kq4
GReZp9oqfOgs8lnjHUuOW9WyhyLjc0mDhJNG0qEVQOuSJIlqY/YSL/UVJVDxFAYc
3Tmdn8YaB1b+NmP+TO8PZ+BP3CqoxY9Tj+JhlZVdWLwe4yg8a0Q7tsfZLXDpiulN
X9LS1/7h4/c5LR69OYuheqHh5hx26Hb8sB4hbdNjsZu0fYI8zFA1rvrDQgFlH4FN
Ldxa2DuZhQHLjPcZ6ktyz/r+U65Cnn2BcpwlXrCqrRwiHOHvLRO3D4WtVv6Roaax
sfddjxgzwRgxolnNbW4JNwbpLPjwHuZMlUa6RDu+HpXzrT/Dk2XVIa7ZI6zK3qMz
kFyi2Us2DJdOe/w/wNz3s5TmYu9zImTnUDQmDSduBMcNqWKDmATgldImgD1ZGia/
2fSMDlQ/NUxGnN3QamZDP7Fr9yu8hSX1AtCSiJuyZBDIAjLS//h3ypmA4ARdFXzM
1iwzaH2QzHDBXzRxbmHzVJot51tNRdsSSHtE+nKzb67PoS62giOkZha9730GThgB
Jjni4TVQu9z3lEVDIfMj41kivcRw1TtPceaXzAdLDd014Y04+k2U6TJJZg8LohVg
wbvWPJEFUTZjgA3Vsfa9CJdmE1JPiLXRzci2GM1v9M9vkItJhRRByixBC4H8FtyU
CNFg8T3KAkeRD/4fL7mqfWVbi6+xvaBYiera6dkG47AL7MVl5oDahDvt0JU0J8vX
FPXkq9u05T+h2zmqZ83NgB97srClodkrBRrBOySMXpabdXK37v7nLihBnkLgSkUq
rFtAJIHIlbZrYPY1OriFptzjSRTpiF70DS6pRPltb7yWsZqAi4E3axKz5OZVWr4Z
ytoYIyYvFuQa9BMb7pK0MVeLbqoBklQFqZFjzA6Zguz53kzy1ULUDvPNLUsPP9dY
cPH6n8sZSB5zva0WB9XK9RZMEFXpD+Hd8xFLHMcd6TzmRlzWCrFRC1hIqs9ap5Vz
yhl5VEuW+gXwjONCQGTXwMqTvm2wr2GW3JSQQrzy6gjQf90BOs5uixyCPXsfliW0
MA5gbmdloFtTtR9XonhuuphoEAwYdLXAM1GgmtAfCv7aXCzq0vScLDkoJM76YeKq
rpyecWiquNuiJLfx0jnJQ20bBJXdc3sDMNqKTaZ4ob0OxDmZJGGO8qft5Fauh1og
onwPOz429KQ/2RgsiM+TY/C1he8n8V2W23VrFkYj5wK4riydE/P4GuCFv+LtFwa3
zFUnfX8Bm004IIuZeVBT5ODZ1XaucK6XXafpmXTqtJHUeJ4MezVihVhD0/iYWHPj
JrJfQuPHNXXztQO+qejqkc/T+NPeLfCn2HSLCD+4aVzsYvgwWE+pNUj3nZS7Hsck
NMTzGanoAXLnOUnLJZ+ARTVqkNTFOGNk/CgsAE3dmMg0bGggbvSXVBpaVfC8TfCb
Evbf/e71PUhqiAzovK8MrBY9pryfJuwL/9ego1dgR7e15Pvn+qcA9HvNdPmjX5d2
3UY5BjUi0oCboppLarsrJRMTt84JOgHITlfeUwsoQdyVhznRjueqWUynSjJYa6mR
ILhtqzK9gaQogb3H5QkHPFA9hsit4RDRUanG+WgDxMhn9m9nS793B1r6VHEDWeR0
McqzI974cNAEmrkL2dEZm+9rmkvQXjTSdW95VkwqMbG7jfiBLeD7WkkutePeGYGZ
VB6K9rZjOL9XAHJhv1mRW/XvGhH81w8ZJfxYA0AP4JJLlGbt9GkZtps0KMefLtJH
O/R+ld81t0cPOYG4DJX7ZPrMwDfGNnxBMdnn/ez5qY7JDvrYVbiHjwJthZnQiFDJ
YlqNvjMuMyvOrTPrUp3z/pYAraDJxsuv1fCZ0/wTbrfriTqJq9xhfUgDz/00CAzE
aQN00E+dSHfQPyTilgbkvIyRkT0CgwElYhARwRYUXlDM9kllggr9o7RMI5aAt2I/
MR42MP4sKxJ8gKzL7CzclMams9hTcLJ+CLZiH+QTUUBsmHyK4p9pKhtEJumrTtbq
PQgoUOyqAMtQzEkJ7HKZFYBpbOMFk3LWZQLp9726eKCkByeFt+v7N8ezDUtX90yD
rU10K0lbNQi6XH6xe+Qf21y1v8BHGCj3Dg9UMwZZ3GYo32j0ghgw5YvT4litxPoK
TQLAHUzC7LPjIoOLL11jE/v/H/3zn8a6LaiTWQ7TAu2pMdjIXBq1qpRY5GHTNriF
rlJFFTWWlMkSaYly2+ULzqjAoTSdCV3VxW2dhbLlrLy61i8/nfkj7ZcN9NP7CE/f
jl7p34QQrfTZKvNiRciS0jG0Fbd+OrNJzRwjYdWaJVp0WYBzROgyU3DXkRDeibDh
Y1zSmL5+VDe61SgY2hnMOhprDW3Q2L3NeMa8Lu9/+HE2yOTABA5yJrgdqkJQPRs5
kelHvNbj6op6dvzAa50+IZQil6EMffUHqPDDsD/I4KZKnqVvhKQqwVph9wktAZ1Y
p6jLzuYKiEOivtHN1aCEa/qypRwCMFtTB+xGx1PVKb9c/mXsqqzs9q8USQ7VWXEN
WuqPjiBtwMIaITkk6o6y9HfkGdj0DHdoQrGjgphUS5E4PZ1lP32ZrgtEoN5c2oLe
0x+lHERPlEarHvYk6SvFmwRbfTaCcUuJEuxR+EG6pSaPDHcWHkcaAhxdkpYowqij
cx3u2kMyDLn3YBG613r+mq/8OWj5yX+wTG8wrQP2sPCBiyydWbuJ3EDoCcVyHDxl
crCdx3TtqkL2gDKeuRe6KkaIjCgEwmFY+ZhdzsfpxQ4g4ImDP1yw6k3e76pjQ0XQ
i3eOVAE6L3k3XRcFK+AYbS+Tgqd7MTvcbW4YwRz1REPiz24wz8f/pPDgWnWM2pfR
Q+AhiVzVE8yLthlCKoOZ+h1xb5uc8i8mCmey5tS6ymZuvatj7zDiNLrYU+A/BLPx
rXflCMkrCerrACo3q0e+u/e4bJr4TcUpYK7tDD8xvm16i3WZKSI0tCExJtUhBFjJ
zJCmgy1GyrOA35nfIdH/a0IfmCkHpGeWtMiH2+DzBHRN3s86sHYtbh4Rf3N2Dyc+
DBM1nYc0KSR8L/8D2m+nTyqzBOYK7LTncgmicNUoKAbcBKQlbiPlsua4ICQiG0qD
eoQfWNBc/1v1q4jfUlhw7/FJTOmLmtLzaCJrGKxYw7HW/4KiwQH5DPWWLM/vIDsX
FXbBuzgUb4B7a/Gvuym7ivBt5q6tNSjLSxjn7yA+PmsjhvlVo2TgYDDzl9xoNVDW
pmYzb/neTXM2hqPrQv/HUyeGagI3TWJoFsaeI3xj/hWVw0ojEqEz0PdVmrrFrkDN
FYqRmAISivH+3CAZpfz0DYKcT49Qtl5gLXYOpmQidYm+lypT3ZnAitC94sKI11Jb
nGjoxX8pujDJk95dkmg2FB7smWp+/Nn9lukMymWmSxYoHB6IiMS1Q2D8vZDKZs9u
JE18fz2MAU69ahwKar36hc0Ha454uMnCQd9YK4vsrGHmfWQgU8NsfyS9ez1Uz2o1
S4b94d4z4N7y2fsc5cGbHGRcYDmMQ6YOhVYzABkIwhznUfX6IlA0gJgh3iDjy7dy
wVgsFHIBEmNBWuo9xJGOQ1bSaHVXH8jOOhrzT4lvr3Hai16ferLXgF3d5YdnBJl0
SC1xjRo9NmjO8nJpAhg+6OrrXqDNU7U0IlUqeTdSzahhAfirM4hLtW9Xjh9w9AjB
Or96llYC6IXoSM79nPrAU+nnxxAXB7AaoZfGruMspyvwgw99N1KSOwBAde022xC4
G2jSUq8Sn1V5XTGTu2LvAWeH9e5VgDqiS8KKWNpVqLojEiRGzDH4eXNqbw7HtxwQ
7TX7Nu5tCIOOTCpUUWWJTBk+q4UkETu6H1Tu4AHBWYE3LTRvAWs2TPVyJOOjWRuM
uXLJZvPODPWtNtLxTdKhQik1iMH+IRsV6ehcu68aeVoQ9518BRoi4oFprgv33t3Z
20rWGLpMbVya8EYNGDAsukclDTLP+L7e9dG8L2pW/EZdeGpDAJ5e/SoqYB5mSNLu
ooQrEy0ApMQyt4pANOWKc3gOmSy5LEDwzbVxFHAMjYuqCcXGlvrfhPYx7RuK/6dq
wzTa1xmk0DfYAbwmtGBNf2aNiAaKT8Ql4epG9PepGMN7uQ3oAm0qeuYGjgke+OJh
LE3ZHC1XW5R0Dm1lR8FpVSLkEKwUB9IVX/n8KY/7Xh1rhTJm3jBA9c0F3zOXXu+h
hTPITmQ/dWXdnZRgxBNT5nx7fcW/yaYtDVZef8Kqm1PbFahNkAw0KZyJqHlzKKSi
dDAeOTdDon8R6RrsNDzESSDV61mwq+f9uHlJ89cNZl/kMAxETIkHxKD+U+ebELI6
/WDGjkOlxT4Z6N9l64VgYmHdg01gEZlzM34aFFPFxajhaGGruDMaZDfRtc5YHx8m
ypGowr8/+CA0Vyz20ZAB3K3rmb5xFtahqoYYf+I5h0IqVBve+iPbj0+Wad2dGSfj
p9qY2OcOi3olNt/U3VuKz/LexUwxaJdM4Ye2j/Z+VwPrOAugNOzzkyw+DzxLm0vj
N0vo3y5hZVrf5ECCPxtNC4T5CXu83nElGeJSReqtvOJoe813tyHPwHTU/et/Bukp
52BP8VJxu5CJns6qJPTNy/Y/Q3KdX9Gyu96HN+JF8/A5hVONzkTM7m/eOSlICsVR
iB1bPP4bbEj2H5khCj2iqJuwKzXhuNzg6ryqWyvTdYTgcnOyAOy+GYKUfUKboWHg
1JTh2z1CTiIM7bvkYVNulmILdg5/Anpv/V52tiJOK1P8dm+KwNlgHilcrmIzvjAk
FZXobYihrg1zd40COfHFV14k2o6RXHa053Vmv1zNCJMrpt22lDlhLmpZgzqcYVng
sWXZEcVnqbsjfL0Hc7jfjqXmpsb9ag9U1TqAXtS0v2pOf3Vvw7EknoiZ+AA/YFj1
IlOkL3u9WIwJDID+bk+Yb7YAalu+Ob9ULiXdv9pTdJ3NAUNGn4ryVTj9Gi9XnBCi
7bHutgfPdXBIT5XECVs9E/YmR5jOR9y9B4ziBV+ZWfEAYmYbqN6rS3b3en9nESSd
zu/n4jTM4DTPTgr36eSda0IASkuNEqME9iJbmnhJf2JsIMBN88Q9+tzwgWVOt9Vu
2DTPONcoCNvWJVVNXQ5dAJRXulnr0mSKmulS/fhYto8Rs1OKciR8Sfj5XBNUqOYg
epb++h85iH5prc5Xl+HSLejrp0YS+l8Kg2PfqI8djCKuEY6sU8dFDq8v0S/j/iDv
mEfhsvTPvqHHveLW/PqJw8O2H95A9sGzyUiZr5euICc6r4zZRq01BRz55v482AWC
Gjw7WjwEQ2nCCgFVECqcQkiASDgdxPRbKgVro1DCsIj1iUQiIESbcte3bnOdwXZS
QMadQTLEmjdK7RXQr599jvORItRyC7t5g3rBaKUKSQ2ukgWDe6eQOoiUI7fSMcRV
lIqVffx8HOT8iBjqAeIWZkhZ4q/XaDEkmvhOEAxFuL2Wm31p55P21BURp+QX7C6X
wj3zJuuzLKnyK6lHm+Tq7O/IqjeaYLEvtE0NAtUEXySqK/cu/BEKYw8vVUrNtjXe
ed4CghAIEwTdYV+fIbvVlvoumKNHac74l4rPP6fYYy2Y8QkJeNlyobqbOmfINWRW
MF07pDc/AncKjtmnyxriZRuRIl/w58uEjYdkJ51Mu/2eHxCGFoFwft3ChIFy9Hba
NzJHRLbdXxSbjzjEoZr60Q3EYBhpQKs0va/eN6DZFt1bkcJYBcCKrTL8NnLCaPWm
Sj0n7X12zoUWTO8WFGnlVAMhg9hzKnSHv3sTYE1JO780ZWJTs+gBEdlEAU4FcPd6
ksEfACdWA4M3/nfGfixi2uamVYlB1DYqj9h9OxTMELeO2Rj3pmEFVSROLDz/Y3Du
W/rWjObmw3ZIOeJnNR+KaVLHKQbxmVJbPyyBwWzgIfB/j19fxZ1cno3MpiE+0Ezp
cOOqgFGLXFea87bFRf1H99i5HUuH2QX/eTjx+WL/dAblKtUluzvPtPeYCcaZfpjf
UxjBt/8MpPKZwzeeQQQxmIyziDvS6GOMl47GbeZXiR5y6BA5VTs/bq+MtYblhCEI
1Jbmkq5yTZQyByPA70Qy23lKJ1GsHuxbvPK3aEA5tGC2cI6pM6PmB5jECuUxS5Te
yDRcwLaEkstE5ASGogdXWv/0atdXs68fQ1rv6ha+YKVJynXPCt8bT0Eo17fIorNc
5FJiFR+8hxp7dJj6oqpR4hNovJgqnljLYkyTMBliwDjd2rk2ejre5abggRRKgESY
YVdrU/ikbr4YYQHZmaLAFlA1P53cMnYuMIdKdnRc9KPy8nlv7zmR8wur3BthAM0K
9Bmy72i7H2MiFvNi7nmEWbItKh0sgSHj0i+1t6M9oN8+uWZsgg+Uy3XviHapczlA
oELvQ3nyfWuGgR/k5nvGLv6x7JJxvNBVJnxCK0P2a/Axf8ecdPi2kSkt2m+0dAw9
6QpibvFxemfXiBIAFkz5fLF4Qc4uJw148sN8exL1IaF6LrS+G330ESl0eEszcNZy
j9JTPAnLtdVjWofSHnDfVdTuvmIbSbDf0qZvyJn4vpV4mYAfwBY6+LAb7GEZqhye
y8ZnjrWu5NI9L+xHVRc8x8RwySW3hhPpW/K5+fKQ/uu6ryZHrQmkN88SNOT61RrH
SxDYLKTqviT4OhwLzynt/pXDcCr1GZ/TUht1hhAIa51B0Tal5E223ti0q+hawinL
UCrURAYQHQCdx0vZjDu0n6snykZ0U8JtJqaBXK23abQhRw7KuuPxORJviuQ3CYbA
TYvNXgf5ft+LF1h8AbIMCVzKnSMIEfbHSHHvHmBAdLdKyUqCAREDVkiV7zwEIDvK
WQQMkXnBhxPMqF6LMUfFXY0iYfR5V+asPslmYlXWCzEFELvgW7l+hFW4IKm5fe0e
cNaEB8UBzanAVEkiXPvGifZpNi4uWOrFbC0f5RSFa/YbwnWjwzuso7IjBQftQOir
+rIh6En/1uMunbGRkHHa8mSYq9UtJNvwUe5nXMDwZ4jwpWq4Yu+SmOo1xKqErNVP
RHX8OuWtbXmMmwL6u2+Y2678P8vVPSdw9al+luYgEV4O8JNgpOdqIVlpNLtIa/sR
ElXaRKw+RWG8dArUt7y28t5phPYw+Ixc60/ald1UlCWBxPtYF9fzSQVuB25/YloV
l4MfMEqaK4iTYwDwbsuFw7j/X21MWGnzhq+9uDFsoizs/cSxfVxgddR++aI+xh92
7PM7ByzZT44lNZY5FsiJ9Iav19OxnkxCBfaLvNvECKnTnlrfV4WqweMN8XbFAM47
WDYbJic5rD5hoooeVf5B805VcuI6Qelei0U6nseT4FdaXfDd2f6AkmS7oVFKUJby
iwwEb4+MVD3zCB+vOwyflLJsT/69YoPCArcpdY7Wu+fEE6LwyfGwjpnbkikhFJET
X73tIc+FaoD3By6F3FibbvmYoXQd0nfSbc7hdVJfSmqKXTMo08xQqGpVIVEHotFL
XsD5O0gK69kN3CN/IV6KpsjeeI2N+cKueYpIR63k9Eg=
`protect END_PROTECTED
