`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+UOBdFo6umYoMjLpjCnnb9DoERO9XBDYpzITDDx2pW9t6uqLYRDyaKJJXH1MOHv
Oh6pT2nHpyQ9e5Q9GKPx4Rpgo5R3nrFy1b+AIgvUdG5Fs9Sb5NlLQHSdujJ+tABJ
To6oOOXqpLTx2BtfL2SJENX21zC8FHFrpSNSCmA8z7rMU/VG1B1LVo8lIUY1TajW
LYe0jYjX4scrOn+LkOZH78KuNBb6KKPE1PH/ZnW04dq+TvznvSVlXZFhO2mZ/c/h
adkmmyRdXikErhIlQJfyBkmiOLtdJ+Ttjuh3/bDSC0FOVzUqaAruG1IuJOVioI3A
PxtXrYwpJ3jicbYWSDDsBzLefQX0DtX9aeCIc5f8OKY1o5ajpBZaqPv9UufVyd5U
/iTXLpejWjQH9cQwj0M3sO7vU5mehaIJ6Nl1OLjakLN+9TOtRNIUpZ8AFXmsukaR
2921ITg/7Vl32sEHlS0N9Q==
`protect END_PROTECTED
