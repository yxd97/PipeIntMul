`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AQFb1dGeckU+f8pOKgpZ8by+Btpk6qC7Jg6XakPQ4BrlVbksSDWYAZGN6glht0kn
X/4Oh0fsXBBjLJF7fRMNEOxPOH0KuOg+MbdfbhhoUVNKdXhlMQMuZQYIb44ByNrw
mM7HqzY+CNKUtySSTdgtrkwSV0Gx1UUk80+c8MmtdzEvw1hLD/2RN0hGz/wBi7Ap
cmX+33gl1TvTXuHCNwBOgUqsrZEL785VfJeyX5Jy8cZBPvjBjg1mo2yYhbN3vp8R
921t0edMy758LKAEVIaEl9bg+q0bmXGDs+wqEu6o3ipAZqIr85ypfr5j4h0ZY5Qd
hUmI2pk3DlstnNhQniWYCwiKy11//k8phoIpDi4G4v5qgxvJWPivITphWDygjqyd
khRTX5xVfu7WNxItUwZ3ykqJzAuWqkv+l8JnPSgewitZ4y1e3Xil4gtXmZOnksdz
hxteCEwxnFqefK+RWaLABVv7TLcIm0ZEQ5DO59ONVVN4uZNzdaxLNKgwBtwjvt4H
D8iB/xvJ8lGkE+8oEAPhIKmHxWGkluP8cGG36R0BumJJbHGfXwckbo/BLIIeSeYY
uvjonhkyNMip2ih5uc7OM83qrmFfs1GoFUedS36IyfSZhmsJilFYqfk7icIWPNnv
Xj19AsInY6vYUmJai3qf8q1kQUfehmHMAZNeJ8BFc0DVlfFl8IJnJjQG/oKUYfit
jd3ELuOM4mJn6JodF/txVORIYO34wupiJpGZDSuK0KowU9fm1Sx82KSZOhkLP9sw
p9+Bc+N9h3b7MpBvfQ+luDvakDE8d74kGDbbwoBWae4f7h0Vb7tuCH26pvgndxL7
t/RBEF7TYoOJ3D+JGW8scn4WgW8H3XY6TKy6/Au0oCk5eCutjfMp99mmI5pi8Wj0
ldMa0pmsvsNyN41fDKbADLI4MKr/lS6HAwtQetOFU7swAaQbOZfZCzqzW4EY8oeo
JbO2jPsmkxUO3E/UxnRGLXdbUrSG/02lT7EqSEJlM4p25oG+gufrWzv4wcIzr3pk
Vho6kfBF6ubtWXlDfbZaL/5sLb0PtBZjkKOebl/2XgJmo5nUlCwgTmfu3E70J39d
jFXQDNuAnF0P4+k4MR39Vpm/N4/lggyUZ96mAROSAsTckMlZ7RFJmUni+e1i59RH
nOVQMEboqN1tq4faEznIlRYek+ddCZnEfUJqrIRC438H1KmR0s/hULYNTPDN1wnf
/4bVne4yHcd+mqrUjW55eX3TdolCJZJaaRRXpB20krcQEc/l0WhZGgHQxBptHHu7
XGqYGHmTdDDwgvqTiZOOqJrNMcPeF4qIaSjiC0cwJsAywyUq7MJ2I45tb63nC3Uv
7KjlmTY/4YuuqP19A3i8Pqj6hF6Nt1b4OIUXjHDFcySV2fXLCEmSDtuyJaput9+B
TlWxbQLRMFtSuxIe4XHGg6VzrJUmXOWXUN7JgakLF/LNWj3dCzbu7f3UI+vckaw1
xFrDy3ks7vMrqO7cnN1o+Xo1P9yLj25iwJLtzMosNtQSvV+nlHe4/WaDZxa1lEp9
7+Ym8AmF0VmhAA7zXpr7gEDJVoxJ5Vnvo43OKYLe2MQkP8YR3aew51iF+yGSN8BQ
YwqeMvMc8GKjUjWtcJlDypjlr9NTfIpeT4SPQ8WTzYlZQdFO3uJZdJOYQeFUqfgt
xZpRn4rxeP8AlBs0aP4dekh4gXtoUB1NCPvjwgZhidm9whY1DQIiDpZpl+fRYUzT
ms2AzTZEN6cR5gw1edMcrjjFWsszs1xMm8CUZVUdhXBebMi81sWdfT7myThPxSZE
Uastcl8CoE6IjgeSP6vhW2eCQ9cUbYVIVQsktcNWgEAdBXuBg50o60Wbu06qYgYU
BiG6GAB+TXEYNch3iFi3nzBPHJXNIN+CiYba6e6L1MLzJJn1QdrfTfKAbr0HKFag
JhS21OF8Sd/Ck+qnPy1L4o2N4IJx/p6vSItvkfF+VvCKnCor3Jmybokt9vM0RUnY
XaXbKG4R/8EdQJaNkgj37Pc7YIUd23LhWsCr61jstcyAMDDo98zTAZx3J7TRmY1R
P3YPkwg5ab9UJ7/Qce1jotEJVpnm66W3HWDr8APu71DecSvoANqVD4VoYM3h9bgu
mRBaCnZc3Ji30KEEXPb/aVuFi9s/XGeX66c1gE+AJc2rkV59kLSx8AMkzuBoL3bL
lEQTLaQWA4WuxPr3h6y8u0lpxHQ7aHDe8yDK5QdWNN8MPE7t9pa1wqU+D3YXalPs
O117kFkzMsAB5YOY+lTeOByf/oRxGyylkGBI/Yr7SaoP+zlVa5ksSVLwshpJnLNb
`protect END_PROTECTED
