`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NAOttb9tRaFuR435lm0Gyo+4UMN+niEguJ/aLKBSXplkiilSlPZLqvuiES/iMrUf
Z1VTqM/OOogBOGsp59ZGx36ExV9B6TvZx3GIkHm+UCOqVsMXtNjOZSgf1a9Hfsng
9+qBd4UAG61OADTcnK43iX7pNx/YJyEJaImrM4LMaUBVp0mwFdh1gyEaMW8Q3/bf
1DMyK0DizMe+Awggt+/4aoeBDaYerzQfWFGJE5ZtCGydn1hD9D/2vaGYikGQNMQt
4t28CYITCZ/C5swnlvOuD9DOqBIUXEE0R9ZKWgHeljYYKb67Zb5IY+IXgXuO/F0B
xe2YVWG32hRCQkgCj8mfYbGmayvRA+jKJEo2omiFGTSoGKRfPYNqvI67NVoH9Q56
vcjOKvd8YgTNbbQWjNOTduX8NrRM5KlF6GaLcUtJ6RSe3A3WGUBvunpwtR2M6nJU
GFefcOd61e77FhXsRoP5Sm1Kqce8o0AqkHPGzTnSOTgAKo8ZYammJs4CtUHi0GGZ
rZ55R+ovkj/YI3+pJcMhvpDEAZ3UYadiLAqAkNKR3qZozhkLtl6gOzcCjS2SjGmg
edr/IwaPb4dp96N06fKkmWiNa4RzOHaZ8Bq6jaJznHtbp257SbDfEeRYV44fQir8
esqKxi/spSq/fqpMiJno00Hzm+zlGlWZcj/t/qeIHLFgbd1sqyn1X0u4jWoi7QOJ
8TbUoQFhhjgreI2Guh8NQ+cPWPDxHQ5NiTEzVKYyP23JxpEP5k2GRn6ATuhWa7OV
w63TZ/F9dSGCnQ5HqGFC8j04aEx7I1o9Dawx25hXGi4UXxD8dJlg5doaoEHgCUGD
`protect END_PROTECTED
