`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mexf9jMPC09BknAANVF3ewTjU79s0rErD7x5ZLBDRUwchMYTYYrzk6ZlSMYRntZU
1+7jycpWdn7KfE8iJ3ibHQ7fojzWRH+ETFh/UhpGOBGijSdfde6hRJw1A2VCOdCu
4qVDfFVNttl/cyxVhcgt9ZsH3E6kn0EMZcg8cBLFWCTZE7ZYtKotbl8ldfmvT1BJ
wN8bhYBbudMBqQEfqCIS7ObEveXCFzvTHydeT9xnYQYLj7ROVN9Ojvq9yqm4X0MJ
ccNiViJgSGZTdEvrXhtQqWc3zfa7Mp3JCn5ykvcJcvfbxZX3oFvpuQ8wH1JgdTqI
IHuBCuY01zzqCsgRtcYyWorQbc7yAGfW1YhFDwXxDbFqtno9dGDpLG3qQZ4Ak063
IpYMzN+Cgy1C6Ohkn2iw1yZLGWxZrMYPt43sWz7+b3pb0eoloxnMqnUYMv5ssBA5
6lxiKaRdJfPnOcP1t+QnL4iC/SbC2wanvOWztc8S+HHGapcF0oFF779qUjBQNxbg
xfIJbv5yLuqE8rI7YKlIEfuiDrQW4d6KxMxHbK/S28mg4DALH2UHuXJ9gMmjgT5T
EvQp7pxzvkF0K84gPdnekdYwIcKkt3sDbRuqw/6IkVk0telxhDTLaDs/mB4Kvodx
W7RVZPeRFlvlyOlQaXAOrdvnE4XYyg/QgynXLuOKjP16lc2giSqdNAIM8W1wO+u4
BtpJSgQ+aUuXVMIEy4AkJGveWLO2QNw3zRSVYVwQI1E3reEX+KIrcWORn0av7JHQ
Mhj8YTXPkvD6r3rsM51BAT4M2hjTQ+mOIJjr2TdtAZNN/EfXdgBnvBA0XaLrdz+6
2U20bCaoSmlgyKjhZ1h6r97m+gz/2CUqAhk/a1hOUFq4zOMuKjeMYmJtpkpY1MhC
VEshDP6TfRIrPRHn/GsKECTe7zODM9yWf7dWuCmIrvKvuLTus2CQrIpCSdtsnAj0
ANXTEpcDMuAg4Tqxb+SvmrHgoZ3VmUedi+Z8sFyoU+eaAseZ2PaPBM6mef1cWUQL
Gy7R4mMvtNyxpapZJIq1ZJMMcfxuI4YbgCsHraWigNlZik/qQ18alGtpGLsVdC8M
bY55AfHizHD4sMhdor4OeKqHsBuYRESpMokcrj5jxSbVsheOdBGss1hiVYhaseDL
JRSrSq9kIef/10C5otkrMTgJ6PQniqpVRMZGldlFTxmoPOlIi88NkbfC7Cb8uGCO
zygpG4jQW3JH7ThfVUSsuYmmUo/t6mvucx8BMn5LLzdVQhVoP4lkpYPujteziJdg
Y1RiRW4vnDfRc9H3YUCewNBj+C81bKFeVH8bgU2wXjQ9hxJMHRxa5p39iH8Ij4VW
etHk9jTxsA8sgMCQSxbcEsvxuIGjK+kTK57KdDZFhS4+tsi+RIy3iX+kgE4qObu8
Z0zWwl4sSB8sI9gaS4NfpD5d/O1K++g8BZ7pCKA5nXMEio+KtP8raFsHaTsruYTY
BzPuxja2BVOTsCkHFrAnakbwj4T+pnT95Jn06UF5Yhq5HnJrND4NI9iRiwfvuDpA
afgwmcGgsZAfR9HYzMKqOQBDCdur/xvKWOLYyxkjj0a6lBnBAo92oRWgyg0CjWfa
/Q6ZNJAPpmMbD5QP73TiYlWLYVpvPBOoxIjEAGqNtBxN4hwvHyzptVxf2SJk8T7/
5lTsqtI4nFhN4sUlFbDgy1MQFBgDDtH6q7wsmE7UtQ149ibTnaxzQhiDByNdGjjZ
y0glhd4Xd1ho2OLDb+cNfcUGGkKyeo0kHnRgLxB1BbrHn+htuDXf/izNUs49lEBP
cxVmzBHSDuGIO/9lMaTT3Gi7/Sh2R/1a7APkF5snxRKF1TdKk0zt9I5Xm9nNTwQC
qaC2qRq5z7eIwZoOrnMR+F5Sz/wHdOG9GG4fToj6Y4wyEiRjmqhb0WWggfoRxiNQ
AXdYhTuJq0XB96581ixaNmOkXeuVrtOUNUHvjd31XFCD3E54OP4iiiAU8fIaGiU2
+ABLJwpL650P1k19yP6Le+i1JnofYKvFB7Oil8EqkhofZc1EX+GPd7a+WcqeROtZ
u+c3trq75ZRePzd7Jfr/9r3u0f8J41+X4ZWtIiaM7WjlAyNumLUMcFgfKZOdYPXH
YD29CFymnH7WGPgYKWlzN2WJoOWzA4Fpg0gVz5bW1GKaApmsVIOYsb5DO3pXm/AL
vrnVTsLh5GVXwMiSoHcVjT9Fuii/Epqr8aC6VSXsJCYe63k4tm51OvAkxJIgaHD8
b1X7RGJUOhXEQpaU4+ygZflV1P6HgxVJ+pZ6LHqDxAolpZtyLlAG7moPvvo4fU/e
M1bS2gs+dkXmjVI1+XItLEz61EV0s2kkBqkJlRqgALU3OMku1xAAu/r+AWPOVlRe
FONvSKPx5rpcdd8YWCckLCQqQXFeLBOh/EZ1ma0h+qpC7vLP/LjSY5u15EkjrQ5f
UmM9WUJ7Ux5+Za8kdQrEpfkd/2cuq2rj1qcu0LOTAUOqHPQEF3WQmBJyP2FvxP8n
U87BFd6v+GdAcpCiU1Aqmz5XlpDVgUnhZhNKtcERqZmRyyRdZkj6sFXTHPW/6YcJ
CYtwIRqgX1kJy+eNT4cAkTHSFuQzJuJmN2K2dAjDfJWym956FNXVf0TrTw1D8BmQ
UDf0T7GFsODWg4k76Bc1Zozt3eNcTpri2th9krIFXQIdkgasqp/OOKTPwqoLILZw
X/oi4fejcYydAyzw/NrYOmqjzgycNFOwfwKPQ7VmYiv1jpuVVFEdW7LfZrwRCsx5
+GsRJIilM8g5PefbpBpgZrZbTJGFnR5Xtx9hUvpVsUAiqUUEELqspNgnrISRohP5
U/PbyXejmezZ65idQoFn1YnFxvxnOZfXKniyjfx4EtRE3YhPfFUEFTL2i+CJK2ub
kO4BSlWzS8i0W0RfP9nkdBOOzOgggCt7lFAOcWCp7+uEnjMHXfKj5IZSCuk3iYYk
jCgT9nBNpSYmi0+8G02oASfBEDH77K0hMuV7CSBcBCX9eOwUrMQZ4JmAI3jTI/6R
0MdNnxkJJnTAnnwvvcgBGMs1q4ghHPiwE2JlTJEUOxeS1umqGiCR2bcXzNmWGPUS
aR+LjAqSGGV0lNwGOy4Xo3H03qeO/p4XEM+3TBIO9sz6utjl+JzgOTcoSJZr7TT5
KjdWUVevZiq5Gi29eZxeHXC/LdTnN9bzFbGEdTfN2cMP6hCdym6HEilkUFzWB7e4
SamLApx49ufhbya/S0esjNLK2iSUspV2017A6+Owny20PRt3d2rhqTsSb9naqqGM
HzNTMZY/B0wM9TNm1bmbKnb88lc1nFUbSyUBCrGxUjX0vik3ADJ3mqSTNLlnd/UF
bYgK6NUZO36t/flfhuNd8tS++0S6+MV7qgxa40v5IhL4F+g+rNvBZYz8yhX7SX4N
GXf/jS0uSc7EHjjxJiuHTBBlftd414HIPyIeuaHGbJUT/550Vs4uSNc04G4puJyO
9C/kLsZXcfs9nbNMj2fh9s/4knmqBk86dpUHghsjKAZt965tBafSQWoHniGYUO0B
nsB73wyoW5O4BdSHad7jq8tDafPKeRefjJO0Q10Qco+iONQXYOdmXsuf/CsHVw5k
nzwJwGj5JCnk6RTPNBfMip7hM1EpEd7blIqER0K/+Mh+HCFDwAoYHQe8ynkMATHX
+WIeiGMR7XhuqvEmAJg8X78+Susczpb/e0uI12GETAHxI+cmpUiB0Y1dA+NnQiXO
Z/PCcXAZ1LNp9bwC9f67x8alZWBRtt5iAzuUJcFPAC/8eO5L6caI+t1uCZTO5Vna
0GkmU86BXkXS6kMOYtlzh/KWql0XJ3PLfy0cr7D0kqeOTIjy/Qi0wXAJN+SRLenm
Gn6SBJxuPW7sejhVH8L2VVblHR2yu05BAYB6psql6ELa1tpuiyu1zur8g+ufAfcC
XtzsTsbX2KoKJjI9aYU6y78Smm1n/8uiALdRiaRQ6qodPG1fv6l08/1YVbnk4t/b
Lkw2l1IioEQblqpomn3dA99eggifXCATh9KOr7od0Ad/NPB3bnz5u9a7OmDjCpUz
SxJ3FJhXTxWSNZdkzDF96CaDpldbskeVFNJGpc80n+pvbZhP5UVilX+uOq6M+yFi
WKHgg8anlrqPYGGz1ue+SIArY6FgJrLUWpCAFiU+HqKKydX16y75cSqGTJU65tYK
RVm/l2ZbSKxtumq0b0dpwEDh7XyFIPWCTAxgSwysLXrrNJ5FwnJ+UhQXQm79RGAA
dPzjkUMP1DtK06HV+tCHdfe5B3UIPhUyQHsyKRUyrGsqJcqCdXABtYK9lDrQK2ki
FRe3+2FEDxUSgNT1kXRtRCgRXG5nbOFbJfARtdM3w9Dd5c3JtfxJGSqYjgeH/kJ9
36diTIXhLsmEsJoirhBC7rlRFeFGVNtb8cKFUMwggFa/86S7sahATqrm6JjZRzVR
ELBohLjkceQ63KpsteenhnviQZHYVb4Fa3JyESh9hj2MSLdaJIP9Y0eDs3j6CPpW
QC8SsRTtHSJlASr10h+c+DsHGWiN6rGxF8qArVn0ZSJ3M2p+KfPJ7vylXkHLaS4+
71u5e2y1ErFwNqndsX+2NTfE6pTu+heZ3kMOmUK6bh1VjN0l3R5DEXuZ4ADC8OAy
z2QGL6nbGxCkeZRiq/wwsI/N7MW0AMA35rxBLYGwXALApKlzps30d7kUsPOZ6ut0
WBwU6jLv9D+F6Gj1eH0FQwV7sf3Boz0x2BF/7kDgQIg6DuLGL44Wpo0N00FqlMJw
sA7v7wfh9TKDcCNwmMJT6xhETYFa+Fp+hJrGEsqI6kBbKWQaSvjO9hWf0YVko1Lg
VK7bp1+JnoqviBi92Ki1OrRHJy1OMxqVStC5Sy3KTeW/oNdLDLHB/VPRn+pNltN0
YK2CmzBD0RoLrx/a5oZ/fba96fSUDiZdxiWXrnturbP5iVPhZmSczFPT0sxMIfaG
aJ2IcAgrzybljXSyYXkSsm4xhbFPOFlLTwpS4v5mruUUPaFhDH3F39BCMEDP0htG
PbilB5i2APmbcPOLbtsa5vbwXsjrW8MYFT54D1/lxHVKRJQcpUqRCNmYSkgQ6aVy
AABHD3QaRFygWMe1JWVq7VToGDT/YT1Q0VumztZDgFhD78ZySAcZ675eQO1258Kk
fOB9ongRPujlIjYVRZlNoUHBdFd2wVii6rtSL4fWaDiHHKKUX0F7ZbznkLViYV0A
UL7t+nRGgVpUCCM/SUvsu3A8lHEAMF/vLD0KkfTcK14urxgv3fdxcGXECoOFkw31
gWbwGXjFn0ORfNPEikzSmrMcSDaS6hMuhcc9LW6GANKwa3RGpd48V0B1Pmzg+KLo
FoDI/d2A2KdZb/uCBSSza23Um821EukAqUeoBMSlQVbYOzzhog8ruz2F9YAE0EbG
IYwpimNrKja0YLehtDginh5DVfIMEYPf/TvjyNnLcX6gt4BfkyCmDfGgs/36THaG
JnpGACRVW82hJKTyWk4nFdX2YAtx9JOcfzw+bd153qs0oOd8zv21OppRmSgrFUeO
LYVB9k0nWHiKbfk6OkEkbOmRf1Hz6ZxAShQLrCjIAzfzPeqPtx46AHUIvdakGfJc
JNyPW1xpHecRBbMd85yI5w1v3MBCc7l5AqPi4xWh1JppJNeAFYFYGg55hyg3OyDy
u3nL/R4RNVUuUBCkEJqbjYaBk+22CxtiJ0jV56IraCPzP1RHo0ommk6KpGNI6Ncd
6aRx1KI3K26CO5HbaRFwoP4VajiXzqbo+eF4mXlp5smzF2qSHj+LTLqK8k/yPAkG
YooK8eGwUwImUXeMkgX5xVl2qIafoOcE5kgYZrderdBqnqhIURl9dFB3s5XPbhYA
lV3r/KhkE1m1I7Uq8wgUIDusfWl/0Hv0uOpe1afq103zG4en+bZ11Y9dqu3j/uhV
rCUl1uVYDMbnuinADw+GM9BZC9cQHrRKdhI4VJWTeIUnxlmQwSWhxiuYI35ISA1o
ItITIT15HMPwHO/zAJbET7iqy8suFtABlmI9FyCPa6q+Wjhf7OhYswU9l/30APFK
7LXPjPWSonQXymcjaWz4Zye2pyomNkLb3ZTu4nuL9Nmsu8U4Mjp8eszfQ7rpz9io
gDpji45Oa7v0nuheT8NaeADmhx+gnojnYWZInfczrjfiVmUTUJMInDPX1/IpWG3V
UvMiLURQudl1pxTYT7S/YRcOLDEnrFInTYA8f6hPnFakdjFS+Q53xUL7fPT/X7kh
4kUlrMJisFJ56rTTHovYxCrJI213FtyZGvKYEpj4vkOSVSlt/kROG1V77obZKYT0
nUYwoyjzxYXGXTAfB/oAPgHlIaRfcvZaOLZ9gxADGICBa8ljcEFn99tmopRWBhEQ
Y0AHBb1ySObAp88PtF7NmgZmvwkFB61shadftA3BX07fj1NhkqP1/DfATWl0Kf4s
s+NCsqGvf7RZCc0OsZcmRETbbDtOAw8KKnGK+HVTnqLzWmSAdSxfa4fd/2Paiq6R
KmhrMWaylB8CJmkaa3fXWHW+w+BP+QwQWDX9XbFmLzLGnXcmgH5s/bo22tgi9Jbh
NNcRYe9L7DoxJr0nLXFDJ2T5jGyZsHOEHaYP3URkg0xdue/UToQ9/r7TO+4z/HjY
l9iJsg+TUoqYwUmtFNUSPybkG+q13LYdu2Xz93AJnevVLry0EE2srNLSOclDCVYT
FLiNq0+5JQ6avpgGLTg7LdwAeawjr6JZUGY9wT5i59soDfGDSaveKq9bIXzmmOdF
1SVavoc27dSx7YI6V/s/0qRxPBMzDKSr5sWRz8dg7e8wKSsiu4Wh8HbLpoSzqlxA
zz3Na/VwoKAlfUop6L9AmdpOcW+2VxPROnEgpyT7/+Zd07e73ZVuSopOkxgE/B1K
HUfwS6klyQudzkJ/VuwfYhpObVXcrFO80P2+l89YXBgD6xq1Ih6zEWF3l+nzl/4M
c/y1aJkGG7Ean9sySIAk+A==
`protect END_PROTECTED
