`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PdP6ljqjM4sEVx+qWk6PSBVcfZv0gov44fFzdfb+CtZojCyMMqQmmX2U5+q3x5l0
32xcW+TAfpKgccZuZsiwSU7pZV8QKlkqjlkLF4bnwJgV3MuxVkEUMhrDLuBfv9yP
YjeJXA+5SZ5qkuWt87hDKw4Nwqz4GxxxCMOA/5UFBiOX4CY2ss0OEgJ8HXiWUeH1
gbUiRILvm6jypcdgt8OBwlX3rCWzJ3+5IMBEyDwyu+oGhX23QOZvwxFvjPxp0cjO
6JFC3GVBqzv/xz5uxyVll4qVFcZYKkcZYSr1JCwyv6JkW8VqfFso3w2O+FLcryBK
z9BvacPuxmDzb2y28aSYR1RYXx6z6YusOXOZc3Cg998z+cImHz+lmZgdfYe+TbR8
1RyrURmJxEW614C14OcMZGk5jvLbL9Q4FbtWpeSQ9khkClxl8emv/+ryKz06gLUY
9r3V0a7IbCWJd4T9t48h6dcx3uFqjncTMi86kS7DIbYiISifxlomxIEi8Gxy/RQX
P2VgBRV/dDWsBSpZOl6zJN2BCMuRDMV/p0lqVr8z4B+EnQI0CdQVoTio5c5AfqBW
xB2cWZR94/xtXo/ey3ZCdH0j+fU6C+ajs3WgJnhTTeiywNP7NP1Q45W4UQC4zSW/
HSzRlVDdC2VO7idy8LpQXl3uUKk3NEcdEv5nXWpQFAqQmsuU9xDke5nj4BL63qaJ
gYtjQnWyUrWFwq2Kk+OC66C5ooxb6qfxpFmLdPqhCTRenRNFgtJf01KpxYBe2Zxl
W2J+QwPYGhUfrXt/R+YOR+TqrmpG3LjLNAu3LGRW+VCSlq0Nqz+RGQYUGfBkouLf
`protect END_PROTECTED
