`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvUVv5OwJ3PqRz2QNG2glIMwjZIG8Aw2BH17u8cqZxXtIA9kjYyNv4GarlY1PV/o
IQZjAXNeTABa3G75JZgjatsjdyPvksWhkDEUxeXktzFrDM7h2w44KSr6DkEZtIEU
SAczrvr4Kr+TnF5Dfd/TTQpNPOyBAiEz3/ZluJmdDSFj75eMIw8eSy5OlZMrzYOs
aUDaCa7nZXSODnXVMRAsznU33yYS6wy2k/+Cc35GKuSA8o2UqhvijuJcogwbxzyI
dtx+wFYt5IIdsktfgRXdgqe+8L7421S54tfzIMM1awvxnCq7hMtz5ANc8m2QCELY
TA6F7EafVPPhrBz+ctPxCHv5pWXVwQt1VjQ1RMfjEuWEaEdQqLgyZ+J8XTiWfiZZ
pONEdp/q4v8e15d8btpaqUVhw0l7IKufrvE50kx60xxAVA6WxjUDUF8fP19wjbwa
`protect END_PROTECTED
