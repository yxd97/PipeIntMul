`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3tV31p+X9K7mrg4HD9d1sRrutX1/AkOJEXdW/1UwbFpR4YryK8XU68elY6rC53Q
oONySnEkoIlu97ovH9xELGkJKCxOZ8c0++Acc7SHg4B1WuR/Vskd90s57QI4v81h
TvUGB8KF4UYHmGJn0zhQKH0Il6KlDezDZP6YBfZKyKMvO01YdXAABDcXsVxVwArz
km5xuH0mwTor0AWeleoUmmTTsYaqTHuoD8tEYCT4OgoHYSxKV8SBL7mSTh8DSpin
fQ+1ydSgAqcCSJWWl6TYoaxUD/p7BtPz7PDdn+IH9XaNLuSE/oFV0bDgEg5nZthP
6LSGIUXcbDjZcg81xheZcmH7p3J/TM/Fubka93zqgs6PpBaoiybR0GHIc4TYvPiy
BZO3mt57TsH07uKxD0x1KfoTJuIWu46I4Wf5GdCXFNF+8RV09NJEzIi6XNL+2vZB
xuakrppYrJsvHYp2C0+jHanSIx1OYts+EfJcPjiyd6FU1M4mnmFiPXMvlIiL6+2/
`protect END_PROTECTED
