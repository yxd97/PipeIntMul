`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HSOjHxy8nDGFafblbAjyVZuaaqR2PQTs5OtiSy+Nb2BYblwtPQ+fjq8ttwDxaZfu
y0oCuga0Xw69lmdqxD/e1/9B4PmjaDEIvpQzd8da7w1z5m1OqvgaxBkVCDOxHGy8
ssTcjiUrXwBKG/K27/49diW2Y+taKanWIpdH3qhMH1U20+35NMiqRTzZ/i8KBSiO
Yt7srXosyTUURatMEPQW8MFISHbQm4jd4QSViDnjfU9cVBDirDQ3oYeuh1gITxsm
OkjmZd+/LsQFhemZufdxNA==
`protect END_PROTECTED
