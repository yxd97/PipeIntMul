`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgT9+HcXIGUvfeJr6Zn1faUGbr2IaxRCpSHRNBtYJ+sZjUShrpdo0gq3tL35FDxI
WMPMNHschpVKwDIhNf7qMrC4K7KUVU1qLBvWjbgKVXBTl1bE1HrXvyI7oNkJpHI3
D44CEq8FBY/IoFOeTkLMWIrnlqRrB5hUj9Be/vgR8J7SNJhqUu+mcGFX0ndwsTBG
fFotUOB7f5cb80QwKIKqFMkL+2vtPiwwZUITufpfoEbWhNyjHHCeu8Koym5j15vh
BvBs1LWzakuobLsWRWThUDGg/ZwJLNxDDe+PqsobV1EYBwDdw9sr2xOnpiuYJU7Z
Tlxj2vshbo16TN2lKdDzYFcKLmffehu/ZdRj4nsmuVXoB671fao88fHHrWznS6xY
YVruZQY+4EFAwITQXnfu3yp/KL0DPdGNnp8SqmIuTTZHWtKWxRRvyoVlxIwUr6h8
w2VotaWkDiL6lpkSIpucObvyDuJEZBWMr1TJQcQpMWBha2FTiCm17lBZtPChnVO6
XEQjc0z1oaBDBRuYtdn91bjegtgkP2dt9LlyXy3FqFrJmPsRv4cb9TucHAudIxvi
sDbUESCUIL71ab62wKz/NjAExFoq0JpR81DWvP+KNXugKjGzurzmg0rXN7npP21n
6A6MrbitYZ5JM0K8o75GtPAmdsRZbDMjdMxxSJeGmnVtN9AbBy+xb4UD7qgNDc4F
ztAdOxW3ygQeW0FRnoZdMK0BJAJzFNNzcL7Etqja9HqnbNJ4U1VnWHa53N0fefgR
H1TaDvahzXVv/rLMiti15sOIaxsPQXEUXrak6X2Q6VYvLLmFF7CQ+ZHaez8A3V33
lw3aXE8i6KH5nbBZswSosAl6Vs1PYrWGrgr5Hr+KqHaOpHpmte66Fx/kyATVJBBV
k1Uf0ejTlmq41BoYK+o8x8xmqrjSDPdm3ONdhBnCLZ3WwFClypC5ncG68J8jsBWd
fDNBfM2eRSlL1r9o2oCTAxzQfHHEisYGo2BIowgM28koqBy8oubFcw4wYd5vxN1c
j8iKLj0zqdd9rlo7Gn046vf7z9OshKj4XfVfhBrn07QnBAqVV7lhesL2NUxu9HQ7
zBAkPMN6LyK1pFiMaRXKPJEL4TvwmtqylzVU/nuNsumSzMsstw8FPZ9ch+DQpIPE
ueczrwk1L9D3eKnQfXAYKDDwsGPCzFpSQ4E2TUVDW+lJnxa04Q6k238vWzdIIG7Y
2LrWKVFQgtmmA96xPZERgiDg3+xPFpKgcA6NRh6przkGYoya1/WmOIM0aWGIUtK6
uBqzAzPD2X5FXVQIHb8Hky1qptxpfHRqmmRFPrG2pl4ChyMtcNFHpQuO80250pAX
qrc6tXSqNBtKT6JY+yZNCsy2ur1byvxZg8wb8svitaxUG5HVK/afLhDtt03o8W8L
kZHObJeCzYrdHlhOadftLdXdxraFfC0yPXlk5OGdl+VLXNZPCgDjDiAOMs0/Vg1v
4xwlsXkzbY40wjqTcHN0Mi4KlsZCxsnvrafwqXsGuik2bBslgoOGBEQHrohZVhOr
GRtQmVG657VhpErDfNX5s5BPVEGuuwbNdSmyirSj+UOFM91b2/Fe6NZKYpuQq0Ya
6uAt7BglulEjW8x4ZH8IH99oHDSkjVI61CuWjUn/IFqhzZCZU1Afv6k4tCjvSaBN
sad6Dn0jUKXNt+POvg4d4CYuZUQr4vuQkPpsD08cCqeH4zd2W2/vL1kkCVUyrTDB
pjiPoBjeeZNM844nvbhCdIZVUiReJR0UprYYQPzEzD4KLFimkB5VBCM7No1x/iBY
wYnU2IiVnNVP1AscJMBEoA1eZzr/9tAmwmi/7wc4L3+A0WBZB+MA5WtcCunCFAcE
LAL4FtyF09HPipg3kZ9wUKnuBc5/eMe+1MhyDP8arN1vRpa28qd/y6bEviryGCLX
2um6lPGdq4bLAdnuNfJNgsoElzKQ1uUv6GP3mqiEEwaSyCuY41//xn7iovvGIzsb
HOs5ZNE5W92szBC58X3OGKUQ43CaPcAB7dH+l/oWlLVo4CHMuEhKbpAXhFKBwocF
ekLok5+HbVrNeLM7PdxMmzbSKtEBt0sQt6axUbetwO3QT2DmWBefJ9v5sGa+xZ28
2mi3QxWYsuE1J5SPM1P+vgLcZmRaZG8O9w2L4LcwwesXqu69nYFfWlG6U0BEPJtb
tOm+u9w8a8ahA2nj15tsKNnFYfucsxnCwB3nw0XV7DsiYNVOKg2xRcJLNkOoJ8nM
z2g4A0N92J3/nV2xtQKyqBn57dSVkF7NWIYDOF4lmE9AYCmbfCvId39+7Oef0sVf
VnLqWg0skBBBADzdAyAGQW77OYkdO+DN1P+q7OgNq42HyPuLlzIwT+EgZ7kINzU1
r7qvE68mLx/5Li6eLTO+MPIoke7jx2j9X0is4ROgJCcZ4RDlNM2hNQwAt7uD+25n
7EuU0/C75NBX2DxDuLYGg+9ZXYU4Dtrf3/qHqQ5uY3tIFB4vFB/gftvUCQbrsQCl
IdhptKZskjzCLI0zI4v6+uzKjtFf6RD4PnYMz2Ao7fnpMkMfN8spv5GRhdCMHGTO
MGAYPLQO2y1UTSJ61KNAXdFZ2jX0oiGhK1/qfuHDR7wt0fiUatoCRArHKl+5o5Ni
AApn0mNz0N1lb5JcTzerFlMwsxhR7/8HrPIjm7lHN9AYkrggj+Qiz8Gn0PmCOqkk
PmUnVdp5jAOTh4m7TT0Mkv/1Sy6bymA0uNdLmX3DXupET4/kCd7caWj1QQHa8z3Z
uJfa/rqiRQZdClzKy6TEJjr7JgZJlkP57xUsUTpSV2q0/i8W+QPE5U7wmSrRpzsX
nbjHS9KGefcGWpYCbsytEBNcSEc8sdAaOIpgb35t6SP4oeocbNID5+TNzKP9BpCB
IxmmVT52aYKDnW5NqWeIaBVoQ8yGPXaFHtbxNdROS+dlUI1rRRXMF2tTmETLv0hJ
ctQhDbtN/3QzAV6RUI4AduPAOMsAlsmHwGuDY2i3W7B9Vy5vY9+HUx3XD3rLtFj2
34vS++DLwFgIlq8hUt1FwuMgxZkA+d7LPazenGIRNMDhW3JGXNKgRyDqfQ8++Lb4
dq/0T85MFFDYbhM1L8X9Rl9Ib2zFAE15mbrXl0khFII3999luivzoB+QYD/g26sO
R7kTn9dFHs0dKko2XpA5kw/paE7I6jZ9tGJ/84jg3BoOo4Ag59CFz5TH4j9eW0hf
yr/wT1/3Nd2PVfzodfP/X1mXDR0fRzhUNuxa/QGMmVu+Iks/kj1Sw5Cyp0L17d/e
5pfdNkMRb8/vXb+Kub7Un4l8aKD9u8FqSyd79nNNxdeobC5Ithutp9XUOjQ/odk4
8yyYINahgnhCjeo7JpIAYQJqRsN/d7P7YjFZMA/zMy0UXxdfwQOyzYuT0x9IcdFI
EYCYHnpzHr/tvIbSRsUJAW8b7FuOlCsOm4Yat+Ok+nvL+g/sS8L6mMIoxbWVh+wa
GBJCibk5O9mrY3zP4a/WLsMVkh4P2T7oyPzNTPQUDhtUd05Oak9CnnsBaSxkHUHz
q6LrVLA+68dpw1pDdIqFl0LdeFT2yS+/ZisSmHCvp9BLOQiFfmPtXtgOYkKT2RZT
Vtk1GJOLhTvDRS+piCupkDgfTmHHE8/Ixz3lSl6QFY0nCv1qywu0n6ZwE4Ky4zQg
gh+zmTPJpgRvu6eIAI/F7PXbJnzeAT0a8RsoiWm7dvKybvIWLUbsEPh7+JVQ3NjZ
QFAIhQtRwSM63Ko43/2IGEROOpGIX/F2wdiVDhk2rTiZWycKrbDEb+3ZzcAj4c7N
xhDML6/6EVXecf2xsT0rEBh9nhoLU88EPvMUpdjCvvRSNoey76WhiJ7R4XuYidXE
G2g9235MLkCQES/bQB78Sg/4YZA2CnQSbX2SvzoEAIUG7F/lbpZa6xCf0asQ3k0H
jTwTxF082+XqLFUPgICuTy7xfVDRd0AvgHWw3b6Cm5dJGUIp71h9IfclHGrhdlFn
Cl8PzUWenc99Wnd54adv1Q+wVVIId34LM9iIBCPrLQVRuwQ8WoNO5TuW+3JKcN8O
EP6zR3syR3qhcnXmZ5GS48M7KNDc36aaNzoO8BiFjWASU808ZuRh0sqkFbio+IQ0
bdA1zqp+G8NjTd67reX8apfRNLq2emZ02lxt8pOKXXFzYFNinfT/XYBQ+nj1myfK
sU3LU2jPcw7RrYLHo6ES9SFflruAdkXaSOouwxwT9eMqz6kiflD+P23bFO5BCBDF
pNk/4gt+tyJh/V1IxK8wDZJi4SoXW5cyV99jCuUzPMRKkkQUzKjKiDr8fI6oqJaO
dRr/OgDTqxQGDMlBELPvj3dcMiGhaSl1o2JGZ/QlNOy/nginm2KH5+3l1zR4omRx
RSf6f3WvXhoRr3ZcyTNZP7sL9hGoeQIZBoa1epqTBs78TuxyulK8zKz1bzn2PhXT
OIeqZ2eR9XtJ1hKxRjVHBO54BRPMH+KEfs6HcPJwI1YOFkIeglAEb+2gs+HgHVk+
h8bQHFqwV5FKvgql2/m35yZyz3BAF7/Tc2hMKaG47FCNh3t9H1NOgAiD3uVTuy6N
trj0Tu6XUV0IFcYGzjUQeXWIxLUb2QDpcvwkt798pDHI6A27QS441K+REDyGimR2
toNUxyUiZ6WJ9Bm02Y4POkEh7FuDoK5GSOKoVhSNgX/eZt5EmaQoWFr/qsqCwxuX
FO9Fc6WGG5lV53wxvHjyic1/jhGvdsWEfWEah/io/Tx30aII3zKaHdvJ2wABSwv0
hrzuoHYMHxjvwmbGl8lvciu/ZWLXh3T8u2BErgK/GF3HPo8ClfyC9NmhvdBnz/ts
96fWi1LDQDsxrxSxUEsaH2aGtmrYJKrLjNWgsCof7+1DV31PufCW9ZO+UIbhnFkO
ALjkE6ktWl14FDk5jVxaPkt1sl/dt4ZyNQYo4ucloyy+llclDzAR7RVRpTYPgXHG
pIckHYZqrRsRTygGBjXynWE47xxh6M+P/+Rlpf3HeDTrIDfmLVDR55SeGh7K0LET
SK3b41Rr4hVcWEC1z2q+R0gO9vpuoxB2KaK+w8LHijJ5glmFyJWoHhEZDCHsnoia
egcNO+yFcpOznVbO3WHoZz9cJBPSJ0I6+lOIZrcsudGy2p8V0utSkVYRVT+1jI2J
+dNfmVwsCSqIItQ7iWMp5/hL9Ipxu2UrEIRPgVRESqy8fe3AzcUIMKyL7VSbjrTD
UgZyFonDhbjxJWh2+skoyKL89+R59gMeQaXJUfpC8WmFXYB0AlEXOPjKVEMj2c/h
t0W6mWSyALwmEWLBKeaFJBNLYMuDJBtPHSXgdTyLLhdjU14Vfp4F2tLlxy7JCk1g
zv47IYpQ5QgIi/m1mOebBVEIClZb4eXeRTuvObfwwnkhTtNUTj0ATpXpbBpQsOyA
sR9aWzf34dtVFw/krWjA5lULtGM4PQK/a39uXDC/S0QjHYBaKLYhI3MyFQP+oWte
DYliQwIP4UhPKIsXeVEEC+/+/FqbjzFgu/fqNJPShTj4UTwYrDugianqaGtkVVRE
yaDek7oUlDBr2Hh8PktJTO7fM+MQsDc8tG18Ghwf+Y12ZRuiphedu/RkRuL8AXzP
GDa0ZYNILhODEkS7ufrVp1SLQLzw91V9EqGhFs3D9k8u83CUuzoEqAhX37GvJTfb
1zcAXCgXznEgIsUcgOkff9O1f7KK2enycvxOtsmtyu11zfpJUdbkdPqqFP1EznEP
uR9KPKh/keXsrIBAcMJuDOdMCj7xfAQlZ9G4l2mOvxzyFestlNwLP3W985GlJ0zw
ng4dL/ciuvMyhmGzmedK0TCU37JQquENk+RIOBj9t9ILPf4hH/firqQdQc9wMuO1
Df3fGMw83Z0vf1HZC+ou6mKyZpVmcCOXripiiid6HEFUmdlIaLawUihL3zTWUmur
d9h6p6U1uHhqPeFHODhKViFCd89E5X7CFWWoKPeJv5cc0Tn92Hw7G2Gwi6G07v3k
B/OnwOp9KLmw40yNIz4UiUZXRvV5tPT6sRGy9D4OeSFkB8XDmC3/LotKn/TXfQMo
OkfSchVjcuppzP6HwVlJ4U6XEzDjLMyROWS8VIiIPmc0PkA/MS6qErQDSVgt0a6s
GCx5+vuyBsQHpink/SFirKuJLgranYQexYCcnIHd9t04VY1q8auvdO4kLzRs2mx1
R/PkMYfnHeSw8v3QqD+a4m82RdwEJRItqvgoFZ+FrxIvD0J+34mPoMFAQx7GI98m
bzlA5FNwP+ebJCGc5hvgsMIAigvDtJVI71lKQCIuwEcxGa+aD/DU92JzrD0BORBH
uYyUT5eU/OztgVPoNjuNpOSrf2tTIPJRReHuv4cgBeximyXo0XsbvM+Cf2FlkYd8
TzmYYo8s6NqE8P7iQVk0sdDzP3X4hphOcuVeB/yCE+iSCcW4tY5azNoVEvwjg1WV
Q+05eFibokhqIfJfeJ2j+nQff7qYaiYR1Lx4pQDKzipj4mB5yZk4wuiri/+M7WOK
gFDg08kK5H7FxsNbpEvsFD7mjV7+RQersaLMeCjV1+zvgxLTc6TDp1XwPAmpKGtJ
UL6i8o6IenCBOU2HC6N+USMj22BJwAkQzVDk6t9ucq6KLcQwxxOvAMgNtkgkn05F
ptOoG/qD6SGoWXuFeYk+Re080/lU4p4q+LUxRnyZBvIq6nLAs7PB7JYFy9Nb/6ev
puFM7l9KdU5gyQOC6p8PlJeVmJsbLrdkCG+yBJjmK9IMVO3YMPQRAY7zyV3D6HZH
VILJGR3HB9rTsfPpvzIJasMA/bt8Kin/cZsXBJXEnbqs+/VutQ0Circ5h5Arxc0+
yiuax/UmzANAx8I45/Nx1ILp332oDY09cfoAjqTDY7bWFDyQeXRvugpgHN67BjN7
WkpB2SYpcF7AUPdrsxjgJuI2GAvKfhYC1ZN8io6GCFpWjuayv6P1DLG/8645Ub1i
PEivtom56CWhCmr/x31HhXkC+58iLpoNmVO0IyVxWhvGw20OF5ggvP4jUYJPC9Yi
LUZ+AA8r7sXC0lY2OeuKMVHbzFbe2pN/Hmnsy4mGAY7w6NTWDytKvbqnvV9G9Wab
W3PhL1+qKmEu6hBOOfOCiDS+JW8S83Q/hwojOtm4pSYkEWIdCJSd2Pd2lPUkFHZm
eQoXWn0yoVhuJ3YaBNdDw8iTX/LtpqRoZyj1ui7COdoXxtN2jSGg0u9zcCCy1Q+P
gO67yHSXTFAN0ybJCAhuN6734SA7c5g7ugq2hqJHQd7w7HT3ogLZlYozH35Ya2+g
BGDboS6zViwyCvkQIOEi0ou6XD1pVwh0zVVllTBv3QSa2mN7JkUXDiA7tKP3VJzu
g0w0LLLIQiqm6QvBh+qiB3EqX9IIYqRQzyojPc6hIL6iESXvAjFHy2vWZt+HmVLL
Adi5W1vNnLSfpyH7I03nle09X3J5ajHKcFD1CaRqsjDnyPg8Bxradypxi8hrIEpV
yYX0HusbhS2TqIqD8KhL3M88zJdDnQ4xSSNgsRrM/JGUarelSyocFYfzydvh/iLl
WYEI8uVsaXHOKu+YgiCo0SZY6qr64vT3xi8pJ6pmbcndna/rygxZ1cOv8YKDdxGm
dZ7iI7HCYY2KEawo6uMQ18LZpncazLThhEPjC6BMBf8pUcJg4Zog3rr0x1xrzyrq
M5TZTwZxJWn1Xi/IhrJLGtiz0ZWqEHXawq3ZV5iUjjkHdKK4K+FCk/AwI7IAQogp
G2ltx6zPCSaQHHK4yGYUCzIt6ScQR1FXDt0XtUrAFur5yf0c0BUj91A9ka53ZCNQ
Tjhw92QIfFvSpxojhlL7tbtayRpL45V/r240E6LaF8y2/nBsptlm/LuvjOl/6VYN
K8og+/BBMPU6/9RiNMHENb/60I+o9JbnQdrSh8QXdzSNq/n6a1USeGSRs9LJncES
dAcXlceZt27H0fSpJtsZV0D+2Qd1A+2QWXtugyQhnthXQTleJPoWZ0nMCgSQxM3R
r47ylXXkJuR1hdBwJZ3vSrxva32XtStAEajlFrBsegthGLmuv0GYSRkc/OTl58Xs
Ypo0FOd1CijvV58F2kFRIZGgWxgbLNi2i63M5cPWs0bOp9Wgy0pvCFs+FJ9qYcfp
hic+F4N2HThyfs8aQqpTg/fbyOT2jAChf1dhDnJx/c/bTlbT5cTUvFrviExhikWJ
tEZBiy4TXNgav/vCi4kEOJ6Jh3jr1Wuq8gyqzaufWc959q5VFkFl0Ctz3ZizaSIM
sBokvAtkFqHvmbs+VU0nm/uwVJK64jWXhEgwwd1qxkBGVpa+8Dhh4XDhX7mNtZAP
fat68C2JH5yPevU/K88VOX+xJzOA4B9AqPnR2468kmjm2nM4xTIpbrJbq4FGAvvw
pf9FYEhmcZ42h/5Rbj4sWAUvy73ntrdGuYXozyQpupnGjzrJeH0asKggLavr8TH/
0B5P3RK60kciH4XXkJyj+lk5q7kbH+YZ9cgnT06RnaNRReagvYnToQUoRTjoCPGc
g2N+bxxOpfJ7IKHex4TfKqZVXY8ehOLDqvAoApsT8nMx7DY/zU5NAnO/LkpiBeZq
FnNeBtfEBIs0IMYBVUtlx4PkGs2tH/48Ms8LHW/KL8eLxncir/Fp/E/oP5IIGKAU
WecXk7CXvLaCb/lqrY5B6L/SmOVPYHoTJyAGABRsg+gw+Ol7TZLJgYLKef3mQgQv
DQFK6dFHWVvCVtkNovjBbXKJi/ZSoJXQ8mr7c7dbnz4NlYh6Tmf4fs1b4UJ+Cl6n
37+DuS78blST2C47AKcryxxiWIMwyAOasL7trIV+7Cpg+kN+HG55kVUMTzqh/kAM
6IXH/e3mtshpo9oynHSJ9IzOFn3bWN8QmreUClQg3wKRuPF2CWcceDgpqngdGDIn
/V3pa4RXx1Ki6Ufl9HkJSWPTLQ7rk7pHi/t245Fg4CvFs1daJMn1Y1pMK9l3tDjl
jSM5/CCxmO4vfk8/iujFakkJ2eGDlX7Kvx/jr/nyEzej9c1uxD83FEG6lB1HMBrT
NxlF41nR3cFgcMwhOgIQfDOWeSelh1SUNgKhAYPImpEZnZp18tF5+q8yW+dv+eXN
C+PJiZfY/hAiDoT6878h6zUAvLzpIaMNEnzWkQVZzaMYFnTa6Te8kL05GCcpu9jC
csNwh64/PPrLtvCmmwYR+47DqOystBJehea/fKIBYyXRtv7xirA9QUp38VRinVql
Zlyo9iVz9jdGmc4kGsoJmfd93rqW+93TftpUpPsyJUno+TzI55TrTFyqVROcNvC0
83rJEM/zw6Eac6Fb6ayMti/q7oTz8DNXbRuO59O+gzr4rCYiV7D9PLmkZWx5qDrT
rI9nZYuO+eKZQgqF+8Cj0EeqLSIYYS3hR4N8+PN+aCzgDLAtTKqx0vXwKgvS+Tn8
MaviERrPa90s2kmTixMYwmBACC29ZKRUvs5TDiX93yFrUJZkMeT5KJiPW6c6UN6l
a4MqoI5v8SQ+yvrRMiBmFV1NlT0GkzvQzVgTEv54JEbgGwk5zQC+cn14MmOu3qE+
Ovv7GA237pSbZYZhd7bEvp2mWNS00f7f5MxCQNJ5QcnVtNwaMV0042YuKkJrt+SO
X++80AyvWBz6iEyLS03kxQKDcQsWtoNIpA9ZtrEmfYswQv2WUrpl0F3zSS6LZgQI
HBHX/Bvzv9p+h14coLux/gxItS9GPVFMdkwoK3tch/0Y7GoDS3udcenbyA9dJguH
BjFO6k9PwSHFFRI+PUqdMqIrtnnhSF8TLURWBe/eacOePo/udmVRiG4XUb/NPbhH
WX5gXQb1uVCOBjj9tL8fgBN1GK+OppeNoTrK4EWuKwWkzkARGPSdz8zL5N6lwUvR
vxvrigbWp3I3pXBNwyNBGQwwxPEcibozgG0bh9Qoq5bZ3cZPE7bKQp5+4NRIagcX
lcMfzA1egS2Fl2g5T/G82WRwBWxolJN0qLsGV/yNPV778DpcKxkGBvNCSiVvB6Zq
ShEgD+hszfRuWOIl2hJOyVOMrRVorMqXlaK2LDo8c8vADCTkH070owZ2g+bkV+Mn
AQ3ndqpLA1EY24dyJpxMDo37BJTMNcIfh0/Bs5zw4InTkAR2iuOS4nzS6W8HFSNo
wYQu/qczqGbO1GIla5ME2vVOLb44P4c69ey8r8lFiRXGPIw4bKUoWHUdgcsxHxCm
ET85425kUmyqPKNnKhlqW1Qxw0Ep3v4TdIGILlALkqi5Cbc/DqUdSz0QEe4UXPkh
UDHGnW3KJnrtLkXhWGF/RpLR/TzqowOX+5SXqNSckTB6tB3e2jH+zznkwxYdnkU/
6OY79T/PqlK1fueBNLun0tAxV+x7o3eQwxiOb2PWHP8izXoGP5xiIq9qlzSc064a
gsPtNoC0f3xe/kR/4BRU7t288IZcD3pAPV8Ae5ddu40EKNz+psoAOO4hMYTqTiuH
qgG/99G1LXg5wjZ0mxqNm/1lQQXaeJvWixlxDhDpZzl3ZPL4OdRzKXgpptAHA7bj
tkgvAjbkf8wlAdx/LNXkIpHRldrM1gvl2zKRdq3SMX2/n9Xln7EMMMI7+ubp/97l
7jLk171XWKxz3lNNOqRfmltrD18F1ri7oEYWajbVRVGzCKc49waneaeAuR+qkcbo
UzD53up47TYydoorx0LT3pC0M1mClbwCPQ3VnRNjh4HOp1LNfxqQOiz1BbjnYsJW
Rt/94rnj+S478h+944mk9cXo6iOOswf5nNGjZ6u5yjbNlMka+tlrMYNfYgMTihVa
PjnURtPkBSmW0mnyq+8eo3aZv9na2WTMXo8nSOWe6MlXBafp7fOQcTRGOiG8pOGq
Log7tc/zhJeRIK/GATskNFwMPDxpC+YhlKVkzppi4mbPEdMB0/6VoNg88TlTirgo
3QXh8GOOLdQmK0ZaLSBo7NluPHsA2oYz7o1xlzvaWj0h+VMyObQaLM90EzVAkJck
iIhmplvBMyIc9/0e4Ijhp7j77ba5ERgq9kOXWoMzMdDM0fusjytBRv7Otvs2m9Ie
YjeL9VwXrkvawTLaFUnXWmYcITUAtANMUMrUfWCp9g9BO/SxkL5lYisj9RVSE/+K
s5CawxGnFHASocxDhab9xouV2cdAZ1QA0/1eG/GPa+uLP8b59f0uY0zxA3Xaqwg1
Psb145nAlAV8Fz/S7OsSi7uGJG2UM8S+biHFqEQHjrSGC2ciM2Bh5qQfIIZk4liq
lEhjh7OSn9ZoI/hIvs4Hod8huW74daFwJje1wCArIekTbF/39F51otQU4BOZFiG2
hrvBBBygO6dw77XLbz/i1oy+H+G+sPVgJjloenpv4duRXsS/Ap4kJCqSXtIypme3
98eg3ANM2tgl4aOXaq2Uj8gHgxe6ahA0MiSjNtKVXZwWWgMRB3lvptbcPmxf7YOE
qgwIWdWfhkSS0JmNBEDZlkJxDx4/FiST8jVNhxHtl7aE8nLc7INo9sMBtxvw8DKC
9jWueltfM7Ju6kS3TRGEYefL6sV7YBeyGWN52hOMSxnsoD9OA186CZmTIPE4PUUL
nvdif4l4bPvmYpzn/1KIf+oxhNXw6mP5Ha0mdL/IHtmkdRniBT4wIKJ7dT6sGsXN
rLwt11eypiM/gio5vIrPPiyzv2OD9m1saLQqTk59JWgQtiXL9ZpV2Tot7VLP78PA
fizqerGtN4hk+UZ27uVnPEAvKc7UtClZVYT+Xho9w9vN5T8cuX49tjliPDxL5Wpn
jr1yjDSaM2HO+wv1ruM4zOz/3mOhCBtqcD5HQnQbzp9kXGKviE5cwQYiDlpkOI3V
j6b9ZPvSaQgkEl6cZQOysUkpwe4qbUb32u+3QfemZgCbJEoYcN7CcUA9TofgAfLT
/whRwr8iNanj4kZRmZ2qwkArvWat6snV+2STqJmKGDlkRD5soyt/9aG0BH2d32ET
ZuJmJFCQ1NL+Dj3SgE3d4ps4SuutuoUVXOgIeyjwmQPX378T7x1o81fza8K5HQrK
znGNGGfJmJcLgu6LiCCM1MVyhk9ljhHrEi7e1PYcv+xVxoOj0KtQ5veR7BTklS+Q
P1ipfQ/2hqhLJGkmjAqlVOfP+WuDMmi7+NnGkn5K8qXfafdDjfjM86/H+osBMDdW
EeqevChqiZtgHV8jN3JQabqDI0PIAsMICZt25Bl3fife+NdI2kzO8D4Yc0kiUC5K
YGpf0fhyhiCX6qHCLvE5rWbuMTYL/vUMG7n+lyBNNEpxG1JAUthGGKXdsOBnFWfH
+DS5brPJH1JRXqeOHFGxugau4f8Enz2rhwXNdMqLOeXEPM2t12yREdQGvcQRxh1X
iO+TArLtoRKGmbbsb2QMpcRLEgR1Vzy9T/i/7gTNdRl6U/gQgggLbPURrfZzqG/z
ci3qn3VnWI+osqnTiyiYCDtuF8V1+t3yzBcnrB85Kq7n9iLlc8I/83Pp8rf2sNIi
IQwmA31r8BVZdSvgI+ITH9/HSpB5yEY5UqheEHLWGM8XRucBrI0pIeALUezzkk6w
oA+B+ROHV1T3EF7faVQ6owg2z6AO2JQ7pNrgqhMSYQNQ8vMIpa3DyIn3UV1qugX7
MufzUFnT2GUFIViQrOqlvykGHqWMAWaGkMJcXF03IlAlCeHttzlCdZI8c9NnmUks
N1jDZY905dayuL7iS05Ru+gJmCpz9D1/Zs5rIwwnfZRJal+JpDBaTgjO96MSWTCq
HcyOblkwBCBlXvomvgtpBLxN9xwCv6hYqCb53QbsCee0ASuwuLK7Yw+JU7i9gtZG
CzmeTZeyyFmCgwMowjn83KaTDzNz6JdcjRa45UFo9f0RxonQQlMv+B2sdKiHa37m
kTOkW9iIhi6zLJ812I4DzvNq398xywrB5/5KRGnSDq4LXuLNg/8qPdAO27wPIQPR
v/fCUKe2pfzIXqoeCexGG9JUmOMOk6SR+1cKAvyfl1VEirUBVTzTJQP73cKt71ed
HgyM8ukFX8XkSXj+hu5O67tVzwtja24W2d9n7VDwH9ImU0B8DxFi87WqDtjOvYZ2
sfTWBKIY82POlSTPWCFYVOinTwym6URV/St5lY+VSvwswyEXGHkqhgi8ALl8e1FX
dju/R+iGIHoMpS/ZdOlkyeSAbyKP8JXnHybADveJxOxjHvH9rEFbVbvLQWN9k7+8
jKI4BpZyvlBPdyyPxsnKqh/y9oIRr/McqHTjuf58aOkbsVQIe9cv4Ky499hy+ouw
hAFr9ih2Ked7g3X6pz81/bs6ziFgOPmJe1g9nTWCuqk54JAbJ6yCPjtnl0/2u6z4
7C3aRFtIvF0ABqOrtVMd6jNMBqn9fntx0vDYD+fF1fMLU1UsSsEL6UmMP14Gex96
fHqbnzZanb+JHs6pf7lDyn4iuAFcVr3L9UmDzgPYZaDob3vs+drcZyztcNJFS/N8
ApyisHSZVj/0pcb22W9VHA8RcmYRPKT8cVuQLtdaQ+cuzHQ2fKTUWQ85QA/kyl1M
UV0qYloJwj8faAEoq0pQVwQUxwdV44BSw0USSrbyAPyBjA4+utYx1ZFQQgmmxEMM
qJ5u82IEBitOsXyya6t+76ADo/4rmBRDRaXYLMZS6Ddsux4QSO//7UO0q0WqoLKg
mGXaYax9Ep39DDRyWyAcGWYLh7MH7Yj/l8uWwVBOEPiQafHAJU6jSF8yHaBUf9mI
EKskBSuBxVvsX8AfNcGMKCQY+IvdFKGagOgkyR+E9ihIoz6ut63pHm21Dx/8K9GU
ouyS2wrNKjdestemq4ntGbwcZiz+uamgnCJOIasW2P7xvNdHGWxDWELDE5V1C2Fv
C/ddtzRhwj4srlhUlwuxn4YQ8LsX3DdEdM3kASwpl44pPy7nNdlnYyZ3dxzwOhFE
4K6RBPdoSXMWf7iF4AeaoGJ1+OY3eYwxgqpEJjSIXhDcKH7rPWCKLq3rynFdei6J
NKfWtTK7sos2Rlq7npOOXS6+/4ESpOXTAfTDbr0J+arQRJq8R/qiQPWwNshl6Y/h
NXaf5IwU1hZbENxWkeXf2nupcvJ15Aiib6bXiU3iL4DAAMvN67YPLEc9pM2P8qP5
s1vEAoVxGMq3gWq1jOdESb2B4O5gFYIeERxnRuqzAezfcTPKhD5NbMawgd6+b3MV
r6Q/R/WDVzdUxCHm3hTcCDxvii09btb0Gmq8AGdPKYPh4F+prFyl39XrIN1Zxsek
1A27+Ki07DRSZJJLtsHQcZHLFr7f6Hw3Z1F0FlkFzQQa6QBr6RofcDMDWuawU0vA
Scqe8p2+55xz8Dd/j7Nlj4PVmSKuvtikZXmD/IEzVIOwsClMmR7R+9abD23QQhCt
Qa7wqfugRTiud23H0CMOaFbi0EJV6fa1p036F6YbjjvrpdwZ3o5jj8IRMMGlaqmW
UAYqhvZJhgclUdBOU95jEGtp+zIIVP8vDoKFAuSWkZzcd47mirPLSqrsc2xekSSo
f8DGU3SCPDFpbP26EUgl0K1bnyLmyunMLYZuOdvaphJuXu2yt01PHLdTIsSxg7Mq
kQSaqnXDPHtzVhErGEzGnn/6JiL8rufkYQyhUS8GVxuhqAoN5hFfckhjwGrpv1Jx
EU4QWb/GMpmIORPyiXyBVUFm0IA82AVr71WmMVntnLNH8zCT7487paeg/ZQLrw96
M0bBcGGHIBdP6f5Dr4dWeC07R9MnfGg+LOc/fsQXbNSG+UvqlZIUM3+NELauJcWD
2nI1foovli6RI6+GQEh2bZA8l9n9j9qMk5aD6NxjemAACO20UZksK4OxiW4E65t2
TxUV6gLXEVr7+lwa/Im1mSYZlIb9QcKij6Fc6JthBKLUnLpxehp9R8tAFNctblcr
FIAojJX/9eAXEqHiOX06UGcgpAtR6oV2d9LXMLRaMDUZx841SrFOuHCuOuEQOsZ8
A2NggrGmwLXKS7W1b3pWCWTPYXVGAuW8k1d1oF6HKLlG5wcY1Ip7/HmE7SaHZBz7
dkMedarTh2YbPsieq0UxKF2KgRlbM7tC7B5GwDmVO4ji7V0WBF72ywLRPc71FHr0
EWkMbqrHhBAfg8mAtkOfYet3I4lwa1L8W1vzmbS7STyNJmlmINmJ3l5T7hFK+Fg+
1x1+aiyN8+OPmRElxKKXuoxvrqioe7uWp6LPr7itE5yYXFEfIdkcTHPf4gTSO82g
PDo1fY0pEaerLOBoa57Na/OXTiVN98MSsOV9FljZnB5nxgEEa5PdRMaEJHrAPzPL
cr7YuRGVkyVSUFzFrJCX4uMyaT6rwekfCXStzt3p6lR36KhG1f2DtbVi7pgNgQWB
zHtEGyaF9QtBzfUvmk/raJRqT1hNH4PJNnfsRnoiTZzht29ywUcscivCZ0IvPsBP
uc7bEzIh7iS/YyVSg0WajO1N67vM1DCkHbpr5H+VFMiV+BjXvsXJ14jTmbqgDsd5
QohbBt7E9/5CXtTUma2aQckurN1QEjWv3F6wxI4ZT4hj8qPLU4v26Wg31qy3bEGN
ZAT0jQtVPAuUJSOBbYz5u8eXPEj1CKLIm6DZAc7ggYaL8AaDg7er8FKpxIiNfEjp
osJqIJWovgh4fTln58lWYQvC5KR71/87qQSSIQsWhIjCYqnvE4iQPC9EhoVLzA2Z
Lnyq/u2ymBZYXF6fAdENBaJfDAM4s9F2PfN18uYnlX6s+oWSR6OpbtdDZ67VX2Y3
XrvSxBgbY+DDRmNy9goM1aBAoCsdUShw52OAAdgGpTrLKLI7p+WGTfUxs4p9JG6F
5o6D1555efoeo37ofhMzppvVCd9AlujlzeXUMnSsjmskWuYMrNUQ6uAl1j2+geNq
C9p7FarcqvJYnck+eQKg9kqNtvYLBf9TOmaABseNsKInbWBJF2QcNPLL4rTskAyF
C6fGH4K2aNbyHxLo9SStjDbdQVoWLeC3qjtx/NrdSmZNlnQKLud2Qlbv83hMD5Y8
5LEF/xin+I387F5hwhynd51V17nD5vy1079ShEe8zlHY4/lVKZwNAnqwPXGNmZc2
gDyC0dzbjwqNH94URljADA7kRG+C9GPtMwDiMU3S/7/HW1vDQZ5Bq0fhHARS963y
JVvGVTbg4QyKhbJU+B0eJNCjBaczGYbl9J/hqXhJEXGKmmb8houAzHFGii23+a7t
FOyWdpnBQfOxyWeJgISX9BdyoVoTYqOUpKzYdjXkzXDnehrpTnGz/TUhrEekf9jB
LKJgWrtx7rOglt2mEdOderNNN+d+/2zfXk6+fKBgsBAJA8a9l+liJOt1kc4Yeeq4
t2uyVVQKPENOz9VyWHizyfYuNc/Ie+gecaldDh3u0zqnhoN2sIrQ9xpns3pHqNZn
l2nI8Mt51WTl+hSfgMBm8ztGeCl/oCUlGKGPD8oyby95GMc/SSOtfRtUh1pOcQmC
IKTxbROEM0UfGYjRgU42ctXr/7QuJ+xi6anUCPB5zmueyXaZ9yuO7LElIVdaS3AI
Xx/D4yfF9EaR50WF2BGbggf0Sf5ilRIOrCeoKehraQ/xsF+kE5/Nw9eufgEYBepS
k7ig9rAINyXCAXuuwh1eEazPLhQww3amdQTAAvD15/9cKYH3W3GzrxPGsvyyDOac
0azm5ROWlW0K0xx1Dn4f23IKnOXRbok+MwVxqOC++pZumQWY1XJ+nVYz9YZS451Q
DCcJ4c3ESuctKqAZvK5PnnGgIfkBAA3vbxIZovRRbAdNu9vK83jyS+jUDbqdIojf
zLuX8gdjaeCmLI31Y3r3bxsLXJKw4RfNKFu1Qgw+brBNlrZw9kW3b43MeZhZCZHL
mkWr5L5ckOuCF/AYm7R+zQepLvEvaaozMAW8G7mjGhfphfc4C3DqQ4BDInu2WAq+
0rKDlA8FgaoYUjRxqPYGQibvLb3Q76thSk1pjJUQ7KejR7adtU0anwDejXelopE0
yHM+YZaLdFipYH89df5WGTTZTJbD8D0Cn5sYLAntUqKPGMCmf9Owu1RN9fvgREKv
QJ9gGfRp0nwD7VsTXzD4VaSoQDe7nU+D+h/u6cd4C3ZujGWyyO6R/wpBe/eOn1ug
f34KmHhYO5E14/nUv5L8Ia4cz2xivc5qrGmv4/NUZiY6eHyDFODArC4cim8DSyNM
PGmr51OIwEqFyRUDiNc4XghlYjAIt1RGl3OcxGFdCv1vhWfWXD3WnUgCpoP2ZUn5
RnorysUzFoDcLASrw6GJmGxOHgG31fgwWPJ5sdYfyTX9GcDLOUuE67MRIyrKqcD9
JnnHIvykq/9eDuCcktxj6OjzwYdPHabDhT2HrLkGxDIDyRDCZF7SIdQpB8lYyUw+
RwJY2AYj6StIXgC/D8SMizrk6cnBD7+2/y+P5EIwfailBFPosdDAcGR53x4Mo2rQ
kPQgSAQYEIi2cpU7qH9Jd12A6OKQoNzgYzlD2l2mVldm/M9Oyz3aDa9zB2RDd7Ix
yGAV2kUsWyUO59dzk80kjJM28qCPWbJTgq88PezPPBNwI/RqtVRu7LTdpVnppARo
TaJQd3qgk1wIvF9snMB4r0Jrf1fytbrt/gfzH7kI/Ah7MChGb9qLfyllwlfBnbcQ
j80zrDxRTioLwys5FVEJhbJ+eACcxTPEal9NFNu7F9uoNA6h9qy69QCB7nkmlS28
crL9YZKsNtJffDraFwf/QmTY6LLmgBbNCwRRDxcX8fQS7yro7GWzQoz6/uX8sp3u
/X9GIKXYpu/WhjqDmBYFlMdDQVkQny5IMmEuZYzDWLsEURAbVKWXatxS5O57kkrt
AjsdCpNtKpj5cWIoyfNJ+yIg60MTmHPtOrsPeENxghtphORbNFrfyHh1KWHnhs4+
V6mNjTIJ8kF522LE71qM6gJ+Zt0pGFtgBQCWDnY8RuWQ7zJRfq97Gu5oqCcd4pSO
mJM8UIGJ1g3BEaz1KT/gdOX6el1vNMHPyxK0FWTM7ysxoY/OfCCsGohbo3ih8Gek
wzHaETYKgK3OSJuBge1Byo59tm+ZL903gwJ1Vtm8wcM7WiPn2zprAAH+KKlkUO+O
+GySgB33Cf50hNCst5+yBwPU75rCiFN97txj/t1HIhLKMFJEPjl9s6g7hoBgipEi
Qu5ZtrN0jeLiF1QOPUzAYIQMWqb1DzMBjbjlOnxfAoVfyUPRKPOxOGYGTYApabM3
4yoqa74OwavM6YiEQKQeKORY5gMzbH+aaedyfh5kxkhi9fX+VayQcSex6dq+JYD9
TlbJ/WJ9cd0BPRj+cC/+cLVp5OUcmBH6Noj89ipe3/uyDhZAA41sg+GWTtDPND6J
UOYRolZH+xXsNjhDuixIGnSdFAG+6ux6U3lXOIH15tEBN4OOkOB6ifasMSyigOgP
bb3njvU2yqO9YbIxBc6sUsJ955Kt22FGceJjazVWVp9fbQWSUNvYFWDFOe6Py4ms
Ro6y3HHsNHOBXLoIk7XyEWZehpL0+imUs5ToTHWuP0DNcgFFCV40eLJt99Tm63LK
n29KHIWn1rSfTizldjmuVykNavYzvVOM3rVvpE6+LK4xYYX67/hLxlSEzWljt9Yh
SrufAPbEC1ufPJgU78zv1kLrTkNNMcMLflchN8QqTq2FSTb/BQ9E4ij+0xxF+Rqp
yaXFN9/VknmCdXXvz1M69PEz1dEu8Ds2cW9I+WKfz3nQmdvHgUU1qK2XjWA6w21P
T2+pyUmaMvBqj2QsrL7As/f0P+Diz/5Jm2752ycXyaIzwqHN5zyNOlEdizmB5l+u
uqVOFId1XuRZP9MiPFW3vRAOaSwwrbezUfTdgjcE/mAItMu/zJmuqRc/JPspUwIx
jhEEOvL2/PO54ZMTbw4MCScOcU4TbZhz6F3KxCzS0ecZtTx2eS+YrMp5dkPopoVh
aFIqI7DAmbueHLdIY8X6VgfHS3FX+8lbJTYL8Pl9oEQpxbUGlhz9pEQeXbqSolHJ
Zogc+TdjhKsUaJ1M0zZd45+n777/4CcUf25eSj4L/zhupdmEeJ+Vv0rVnpriyjdN
NIBw/ambcjphaJVcurzvtmguTrLo3iCAjV4KMeX2Ci8gBJS8zUJsybkDUUUKlcUy
RKrmqXUDZcfcJnmryBdTHbNveH3C9FogTEWa9N57sgAeZ9otHEjRL2Wr0FkDonof
EiZytTG9PGJjBWyRM8CBy0adj/jBsAfydUQD+gCFW+lzQC1uBOg5tr8KmQIUjyPg
90+/qIbXMiBJH+U8SPBycyal7/wzlFc62vE9sDYGxxTb1q5sWeeNj3SwANjBfmFK
SjSfipDameZBteJEjChodHtGdrgoq6/I+UL/eNSICQV+/B7c6gUmqMEuo38sVDXm
OU+jJDfcnDQvSyYUaVTMYq9Qw6QOfSwHQy7AXNRLNIInJdghrUnVvymOvejhstPe
gCxNhUYAAUapm/AjGzVuvSE5SMLRP/Sh0dbrLynEWki3YXXADv8469CXYMlf+GZe
cnowKUyN8pB2XI+iWX4MswHFMfknEOvVJr+MRUcv9ih+Dk0J4I62FrJinX+eODe9
7fS9IR/luXbSpnxcTwzgYagdpVHfPM6Yzrh8DQ5+WKw9Dwt4ivU0jjcIwOzD68en
0WaYL96solxC1CGCrOrJw7dmbCnvlfuMTI6ArCV/DfYrJ7jOZ87dhjoVVISKcxbl
y2eNDc5pbTn4pKW1ledHWb+Qstd29ABuXPkyWy9Na9pGiEAEBgfBglkB3sFpx2TG
UFkf0HPs32Xqe7ZD66l99jy5KDCWlycONPktxSLxa7eLo6IZVD3fPYdphvOWz7kA
IV0XEeVVfQsz9hMfawnG5JHH8Mq0L10Gq+qD6vUmzIiwd7Acbe6roB3pxVA7rNj6
QLI+j81/E40mPlDT4nyQd123ZRGyFPstcmxHHFKihDx9650gAqUTIYYDJVAiIkDC
fJUlrAbpWqIDytinacKbCyoTKvX+PrzNIavSMBn/M2JYL0A99yWwQceuBKpJjIJe
PgJkuBDgxldv7KNP9I/85MFqwoejTHYYQix1IyfXKKmYAu/TkvwEkVrd7JN2aDXC
amM5LHBDnWcR6MWuxV+HYa8DeC2Z2Yt/dyqyot2/R0lrd4ouZKodI+t3uCXLgOQ5
R47tsOwQogmb6unjnXioAODXj6uymsKf0dMD5aYSCZkIUCtsr3Gb4wzl6LG12xg9
gwc0LWVaphDhQzR9jiSIsXqUWXB7zm6NEGJrBT1F2rXKyVIdUj22gmKbJ9DURQMr
75nCcW0f3Js/sANvlQM9L561S3ILbWT5nwZfkRZFjutpcVbbnN+NTXXkZh1ZkeXm
2F4kA+UqU6lPZ64vjvMYeNebpEhnrpmDtTVYEZ0WtZobCKbpZ0BwyFiVT7yRP52I
x1BvUYcQZBcOlGA/6DKinR4O0Hi7WxVIeR/5bOn7U/UBK64+B53ZoS3OBnSuk5YJ
064s989AtwgJxxrfbPDv/m68tYI72h9xoltUqFW1EYgRqdBU4iQYXRAvp09ujaL8
lEwFXKZBZOxH3bX/CreuA2z5u9eiDZXoIWthbACeCDhgdL74KQHWYoaGsbPla0D2
gJLNK64SkOMeFA3nIthB48Lwf0c8Ur2ENwHpMiDl1yXbF/J/UyMiOJ4aJXM8P6zM
UYfrjoVqfN/rEb9AjM4jG7XdoM0iev3N1twkRte8GO+XrQcOWpT4kYuza42tAJZU
2Ev4jnHi7Q0fQ5D0gW4nE59f3YWjnbS0gyAq8roHHj7tLNNN6azSdZdIVHrkswRF
`protect END_PROTECTED
