`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wokae1zk+oTfkqa0TyVf1Dj8SUDqasUt0lfqfaPD7twZR5aVGnTjgA/Yfj9WI0VD
za5UoF4SDk3WO1ICnmbgBuKBxEISIyGAo9Ag6eT9bIO6lqG/0+deyUJ8mqBPA+TE
OVuqWYwglVqY2HpOhMwePsEzscswBOsATTTkxfSTfk4GlnTblJ+TWIv9zjYRdPWu
o0BRft9JhT/8Knj3gloBLhOvYwksx3YGuo/XZAyWxZQQ72xUOb73c8KDmO3BT2Cb
25UHU2sX+QHArItkdrZuWamKKGgw3AO7HV7zbP2g0epZVNmjJX/6GM/JAQObgXTU
SioySlF1Gfw4i4YhjOcHX9Vajk5PFQyYqFPCbI8EfHZDYK97NxS1LBFiRAr8QEKT
WEyTFfjS+SKKV0vhAdU9pg==
`protect END_PROTECTED
