`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KkZLlVFSMfj+SyAdAyvW2zHXuCwy7FgFhQ3jWvQlDh7r5/HdRK14JApKjsXE5jFZ
L06FnNQBWGxnAtK0X7mdkqduke/C0wj9VcovBLwijQA/XAyO1XR+aboD/2qZ6wzP
ob3mdIzJ22l8RRa9EKY41KVE3eNp+bnQT4Q7pDhkJv2xqBZ0tniM0W5+xhY5uI9J
iTn1Uepv9PmG48mKpEpYHssP1F7vIjiGtFK4ai2wRPE9Q2gExjdnGfWBcx1kcJxg
66Jo7ZgB9oSf8HoEKJ7WX1UqU5D8qri39OPwe6fSIlKoU2dXrVm/qSMStl/05sxo
vCxMXrZeM1jW5a+aYMrNRYTRUOVCHcwfBSJjpLswrb+TqXB7VtJKkgL1iIEDaCqQ
QQj1GJkQRM92LSZOjblElQYMSW2JJ4GNZ1V0yiVGwraSaV5LsfZ4D+/vIC7glAMk
iK1DB7H9eUKhNUjBqZds5LF12KkgOJWXeRKlVTMoZQBZk10VD3cAhXoubeyo+N8r
`protect END_PROTECTED
