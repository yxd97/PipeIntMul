`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ihVNs+Tk+H5Ii3I+zOR8a8d1/Ni3mz0au9+apdp8BneZ14VYS7bVpMyAzMKVf1g
kfRZaSJ3niNYSiB04OvJe5vnlP+d3K2DYm+NA5Ivl84Q8I31YFLSqJgba9KzK6T9
pNVRAity7EsCy1YwUp8gs/eIt7NjQmAr9xM/XRUnwJUIMBqevs/xtWYkGkE1Bu2m
d2VmsyD0ydvOQa8yRzuzykhHRYLBG8DAoKRj5WuYpgpU8vMcNYC41UOCuDzHSSmW
JQEUVtiZj2mPI18Lkosh7BSQCsJYJbajpW/h0CzYy9nDerShzFCSHPDj1b0O6xcO
pTiPH4xsbF8kzuHfB1+4Ier8MRvj5qXTpYCP8C3ICqfgpba03Rn8TxMLqxq5k7A7
8Qv+YppM7m7AHsA/r5X0MhNDzIOex7GFjFar+Jri7EIlCDTZtyB4PrATqpzeB/G6
xuJfTN9R42OgrMIo5dLnnaiV94zSff1J+TtKGk5izJOkimf2uEqhdMgYJ2IvQqJ2
AtbjZ9WlBOfdZIHDaM6frV3ILDYrx1WJV0tvKVv8OedOcjyWF+HShde2EEjcyiLe
mGmS7GDdLiYDrJZJC0mmMbqlTeYgbhrDQb5MBC7e+m3O0ynx18kwhA+6FWETUdb7
I+vnAYJ6xhf9TmKN0dykKMhUOGYnD1QV0nTO63djkTTZ9kCu0PHgSnTI5gsJ/2Fq
JeTjICbgFTvkgP8dgKHCoI1DrTmOw9h5ZRGKfyupSr8+mBRl2bulhUaZ34bvi7VC
i/OCY6MxqIXD6H2KWDIwzu3uB90uUWzGKJgyIg2xo1WI8Y12DxGD5SASwrnQpUGI
TLLJMkrFcQsK9kHU2Et5dWx7UmaOI0QgMuwjpONcNp4XGefFpn2tODfN/HqKNjHU
6rAM5O9thvUNFOV1/jPDIPB58RN4wBya8ep76pAI4xusZjSqOWvXe82CQGfEMphd
ALdkaeS23KfdMvomQwXnuT6UAH8U8TUMm5eKm5hXoLnnWqjuVmLTTLlTTb1ljzxQ
2qBjybyRCHabhr3J8ltfcPMpiEVD8Jdw049PZ6jM4/wn4Lwc5i+Lj2PnbgTxYv9Z
qTV72eoT9HbrzhjlFvNo/KRzhl5eQnIrx1mCNlI6sMReGZryjHG+EmzZThvZ153a
74ZRorNI7MEvnqGN44OhLfpdajomhRD2eicW6bgR+vJqkL+RPhYw4ZzwL2wmgeoO
pxkJe8HG2E/NB76Bb7PxVu6qE/n5PC7hPZOk9ewMJiju440SwHReMFYmZShAjKUY
W34ZFltzUL7CYof8eC+entsf+6UoRIgR22rlydZodtLBw8CvE8Mtw+wLaQe7ZxEG
yZmgVqw3gBH86gGqdzNrcE2Jdy2e2lgcTKCT5hMrXDBQcafBOBgt6rQKFXO/kitm
gXVpwGzwPig6e2yOB4IjGRM9zPvnRAZLqx6enyhHFCA4lA2ktKqg8MCX67U124Mu
5JR+biUF+ENLFnISA7isNt/Fdagyl5+HOYeW+ifce1+SUJBr3RFLgjOBVUzo8TMk
gdaTLrlVDnkwfKFu9LSjUDJuyn1J3iYxVMbVJiroqjh7EOXUMh8g7MINOXuVySbw
b2cDgK3R0RJr9vYZ68QXod19b/rRoCY8tu+PScCptQqEsZ2e3y1942opVGH45N+e
lMmc+7lPhIyHx4f1wL1w3439uwuCzq1dB6GWivbh/8xlDJqJHGaVwqOpFar9He/h
qFu79doke+AIu33sNvHKzES2ad+uJI9GVsBHw+u/TgSNS5NtD/pG2IMqW7Sf993K
c0Nr4REUjtYOkfOusQmkAxdazwMI4YV6zzM0lZxtBk/B/TA4nn2/Obgs+OH428Sr
P0AUZYPE8g7Q/DJ+4kPr9D9FR8CyqUF1wnIf9UbqxaJUoBepjnOe7i4CHGrksD/B
KRPRQsVXl6G80/csn734f9TLU4UtzpyO9ktzwnkxisAgUjAo8ww2iUgDUgHqqFvX
ARo0J0quS2f5M+dlmPjO1SxsUQ63RkozeGFz4v4J77jpEiBO2L7b6Op5wf6nOcaZ
ScAxRZKYRAy2QyOquCHWwJIyJr6D2rVMGnrXCV6J3KfwwoeG3sYUwTnsgjrcYG3N
2e7mb0eGce+Anvfh6ycRzpeSJ8ZfSumYA8ECy3fl6M4U3v2XuSTlqk/V1I/AZbUs
rUWZDB4DWnUqZerGIuE0I7jki/QKkbXzAhCfgLMxLeIWT3vQn+zmZIzcgDVfIMQE
aL6eajPdTeOJ/wh1IOdSzS/az54go4EySC/FQjQe/duFwyFo0Iwd8xIBsB9mNsqA
XCPt5yTIn+zROE07fUZgAmIX6Y1UCzL3kan46rgyH3bUoi1FV49zsS4K6GLyK6zy
pQbD9cs3uYhes91QFIDjvGQ4WKLSm+sJGAYiSPjE1dAPdnpEHrAZt8R15NCzjrVJ
wWsAaLPw+P1GpYsNCHXwOScmunbttY/b90pqSB0iLDqKZ4YNup5ZMIcANBvjfSYA
RUepFrJaj80573nRmnC9RaWpKKSGPAx9BNlxFYIdB0V/SlAY1IP/ITS3i2Jilwg0
3a922FG+w+lTbnMSO9om/i8nxY2lqdHKRXqVlrkcIKNK29+r2l6wXe6lXgBaodwN
10Ea/gad/pYIahnKxNi39w==
`protect END_PROTECTED
