`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VA/pWhvTj3S76A3/4SjVKSKhZKzBdcFG0xndj73twjxanA99HcBsriHfX1xE4uUX
e34QjxOL66iD/on1ZRB8Ed+2UWUYylgWZEjvKHOPzDqKXpnvq8+KCnqiyF8/axM6
cO/iFHcwpZ9GNa3lOnqBbRAKs8yFe5xZItVYs+edQMzlKHanuOiXNI/F4CiBECoS
pMDzbAUPU19SDdVfepWLhhP154YY9oMhkJGk2dPzdUSO3tC9YE4/AHRtFgVojIzN
RddiWCyup0+1VucoBqO7QJa+Rm/H0Ih+xkGCqZGj/x6tS5PDamCqRLxrs9f/UzNy
kqNojIyiO9HiVMBOx01mi9VEoxQunhiBCGiu2NMobqGFtGPpo4Jt5QJiNlMqImQS
woy6z+p8Ql6/UGIOTDHgMe5v4yOI1vC2DKvUmnr45UyIDKcEujF2azWfCrOz53uM
exTwg8dldukxMJIxZzd38osvOOulRoUFP/O1FDtVrmgY/7pKi/WbNxuH1rG+Jx7T
M1x5hKSqllP9y1kYSomlR8HlN8AeRN+KdDhwNLA9D0vOYRaGajbR0IV/jjUZ0zyk
2GE0lLzpgjUG8UwOFqM0jWSohweM7+tWbVFNRd/71/ALgCawp+g3Dxi3jsXxXzz8
YvD/xzjHRRRiugZq0iSuAHhCUDUg9R038v0DRggh6wxQMIKkJMTQQ78wH+bAbfGn
Fqhw881HeXTA+L6ijh6RLTVnvJ4P1T3HjFLtP79nGSz/2hS6lO67BPgY0JyJzjd0
QmsBn5TZAcFFESyL7Nw01pyf/hAfJ4zbvysB7pWYmEryCewtNDRxHuuvZUv2S46J
vSdZBwTqJ65YruDp8UzRLvfjV8MRFGi4NMdKALHbjunZiUtsJA4aWkMpT3WqCwTN
Od3DkfBT5s6JJy9dDUSeigZ1P8yK4+FZ/iYPHktPPv+ffJBSU9X4xLU0q8eml+zm
B6gPey176oKAX085KixJi+7VHVU625TLC4Uj47lnuF9pIfwqp2qUJ2/Z9R/hZBf4
sqpZzbAGfTkgtP78+/KYK6VLHBrXFR2C2jIG88mjbTLZMgkupUAej/OKdshqsQJY
9ITRDiMKVI7mQdBo41y28aWhl6SGvK5exUCF+2UhDtZrrMxts1DxoqMUEeGittc7
89JvRKJqFORs3T2kFkyZwWmQole7c0TWBf1rthOon7+8jOSgthDoR0d6ySyxTCFL
cokruvFqoEk1fyZVRMScEp8DUxo7F4eMtslLuyMHh3b3RJHipZXgkHzzxkZTRhC2
SRtAa7il1RA8Ch8KT1ZskGeZuGxFlXekl1qbleoQ4PmkS+m4AIOV1iZNx94/QHwj
`protect END_PROTECTED
