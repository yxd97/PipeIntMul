`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDQTYbnhp4BBfN2ZjuGaGf4fqvE+sdSazIegnLcHmVLpMCPMeWfKMhSGkqy7+6c0
mjFhFD2LWlt7592YbtLMh7LcHxtucF8f7/jmecJP5oRJq720WUpwwR1109lgDYnB
q/jjmeEVZ7R70DiP5kFdcYatlTiItVMw7m4QkH8Fzy5TGxs8J2WtYDYxk4xkkogD
iSw6GSveNfORqUoQiPGd8oVIXu31y21TlXd7u9OusTmlddVdR9xvyehRWKf6SWB8
rU0UpeR8DWauz9/aYQVlKOFELMYPlAUQHu3R0H6fACTKKWRSi1XiYrGllLJtxkBX
hScgjvHt4hGFSQvsLhpy+pRd2YGvvVQtLZZdvySDdHEY73AavA3zWr+/QUrYPPJ5
bi82KLmMdsMZcGnAFAy9p8bwKkQkTN27AXOMelYHvRYDdDWpgsJFmbwYLvDCgrTk
4awBaAygQ6OWb5/kD0yjUe/DxIgoe7wmRmKdE/m7xtDxvpL4z1kWPROhVbtQVfFF
`protect END_PROTECTED
