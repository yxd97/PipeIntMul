`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3ztophSTBtzwkbYQx/Z/8/sBjlXeMbjohhJvdkWw7cFOo0bQheJd3OYxXdLnKUu
QlHGRMecyGaRkfOTNQSiE+JEEen/a345bDOuHeBzI7PjiPyfzDUP8Y342HhnH6Mk
v9/HLGBEqzAWcDpp8AcGu2kx444qGya9n20c5E8qSXIwp6HTJTX6RiV79KL9aEk5
3g5VbiYP3xr5ixDcTWgIFSUGY6b+IqSYLtAAkjsd5ZfB52FSykj6Cf6pPR4L2U3c
FzUrFh0uY4zgucMjwoDwByjCpt+i9r/YokxAoDRtXMEdH9Td9c8P/sJuk8wAlWY+
lwJG6rjlkplteHKEn92Brf47uZTQpvQ6/UUMhlJ/547ViA2gyQjZOIFhpvtmCQ4F
GLJ+C8QbBnW1mc9a3AiJz8oSNUKmLOMwJ/X38wL8rUUf5EQTIeu0Egk+QYIC1Wgw
pYhC8vtTcluKfyuQFznkPkGSl9JjwXvEEPQG6Bo0ltmc3bT71N9OYyeiLWR+M8VT
K4L1BCzKyf+DdWSZagQxiAekxQ7QshF0X54mfCwacuhOqcR678gbmJOHQ17DK09N
YwTkKxAMOn+fusoEvLmBAUj9+jLcui1yJfC0NbYSxgkCXumSerSsGSsjOh1m5KqH
e0whCaDpOG8/naNZkqqylwj8HAUE2e8J3sy78hBeWx8=
`protect END_PROTECTED
