`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LR+n81cPEmQubrVv33JPenId4k5w3fEwAagT31RW2FjlB3aQTrSmyg/RHKARRRJ7
OhWtgku3kBLE5QPMp3ONcAj1taBPfHa5DwffbRNmqdNDSrJksEHeOZFQEO72k1Xf
0znK5sVIOpJKG3R3aA5VOSFo5JvxbzPu62/zQQEQysr/gSVQvvv82q+8l+yIxpKK
eRZs6aCIVk6Ij6ab0KRAlKqsf1dFe7jhJIRug3M4F1f9ONZXkNOSkRhFlE5ruanq
H/+W9o/xqSlI7v95sjx/RYP2C9fUZqSq3on3LoIxT+VCJgGJUFcb5weAOD9+UPju
84SNUI6jXT/lGzo3Ek+Tv+9Hz53riLouNqTc3nh8SmLBUPcwf7ig3WYNJKNzCsT6
9845lUMhZl8OuLr2WZ1OJ28fEPvwMsr7gikdKS8QoLkB8AGOHgnBiwPBXmfblw5r
g+F1BEbURNoqbumFiVHgIlUh2Iu4k2Zg6YIebLvnHI9d4r7wefYARZDB07k6Jbf4
+F1GQW4Z2UTjhajfno2cbTAEE3A3hzEb7psTh8cxpvJfXXDiXpi0LrLdvLpq3D1y
`protect END_PROTECTED
