`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sgmXZWOtE85GrygEGIEgBjd36GOy1BgVRANCMDFY0BqtUreeD/rlD+x113eKJ7j5
izuoHo/spgQdyXAqnQv8NsmCVwRhYbdihVLEz5hzxV9q/ibPAre+vKGCuuTpntXT
wdN0oOdrBz/Ssp0s6Yt+kgCAG8yG3j/59R/S7fhXw6AXSs9Y/GnUxWRpW4iguelA
CFDAyILbuPuFiBd7OgS4HrptCupSIssBi5Ua5XCPUNZCI3Des93XPS/nvRYO70e4
68/OZGUSe/2Ny+LcNwJT28ISKgdB5LXNtkNGYA+bG6/Z3ISx6ZAYIWz3fphhYgH4
P+rnrq7uAcsN8jANhcReOfhj6O09hDx+tiVkd1jEcvSACFoRLSohVtn6KsquOMzg
GH7IyJgWQc9/GuC5TqEGi67a3S9xOqgdI0hfCtwsiLs6B3uWp4UCp/bED0wtsEwa
`protect END_PROTECTED
