`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndVd0HcQIIN6A2aD1m1wO3rOSl/4K1C2O9qGK1pszpK3WpKeCb/4pCEJ35oD0KcV
Ylu6dpDHujhP5oGKCzT8UDg6Kw01RrZkyuUJ0FJQkDgZ1jVsg+vdHQ1kyNU0thMF
rENP509Qomjk+EiRJolbOyw58vBFweoqegbq3nPua586k5b9svV3X82HzAeo9NS2
XdBwif3n8Vv6t0ntSamUJZNau5lpGoIcVMgmzV0h3wDyB9ajA+uHAyOaCaG/hLwy
MA+qW3gzzrLt/AGZVpI8PWsVKd3bLFRwV8eLm0KdZ+bcSwb0wuHKB/f3d3dIQTGn
zGtd3Dvn8/Kf7IaVMy09fps9xhBx5j+TX0CsPeOTEzrEJ2yWvz3yY5y7ousQ7Df3
SYV7W47/TgJda+NliVI/dKfhEVaqxxTB1gyEyoxiM6tNP+B8E+uvdjuSSpe/Y5tX
9Szi+QSbY2yaFW8/YVQAAhPfaWL/7KSTzMuQa+g3QqrWoJUSl4I8xpBGWsIOdVH7
nlAuJ0R0ScX4ignwnXSZloiQdYu/DPRjDSs2CAVIa4L07Sq/1f3wSuOHaBX6BZh3
GbQML1pXasmCEDHri27N+yDD7JEWvoX8LfS0Iza49n9TFTU8rgMShmdl3cGJJp4u
ATwrkJE3bIunbQVXoG2c/w==
`protect END_PROTECTED
