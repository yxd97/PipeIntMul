`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p7+ZqbZXyy8BEIcwHaUsX/Tdt+dG4V8Q+zWahk4XiwRgwIiKd+Tdqvn7UprDU5C+
unndhjNgYJS8yDKrzwmZsct9wHLEK0BaplvJHNQ4km0wwkWaInVbIRY/5dTddASk
ftMnNW5fhBoZkl1MqFDAB7Dl0+CRWz4VQjIjRxpaR4oB4j8iwG5R9b6DhG4+pIHt
9imwV12Ae2FbVhHAfdiPvlBzZBWFrUWXkLUgMhE0iOL8NRqNVFqpoD1lyR0v7cNR
Yh7C4/JPfiMiyJYItGXd91/ES3MBPUvADwJMtbKrUFw+MLP9PnnexWFo4hofkrfo
Qj9mvuXdiMQqERGdOpPEL9A7tMRm+hGnAjruj1t8SmQ164QqVtUENjQimQoS1lpr
+b8PRhGgmlg/s65vBhod8YSQWtFKZ48jAp8oamgP9JVhcbotYWdIyWT5G+NaeaFb
nmw+BRIx/I5vHdtbofJv1bJOjppMlJtl1Vb9AxClpY1/y4HLQGDNwRuAmw37eOKo
CaF93PzBdk/BDSYNrqT/dHZtHlRjduakG6/oPihqjiNtl0jUi9e2hSH5Dtwig/d9
`protect END_PROTECTED
