`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+nHeM+EX9f0gjjRmE1yWfDzYtBHo/blv7XifCLzMixdgId+Aai+b/LiVXVdzAXW
KIiUXge5VK+51vvM5aoY9gac1jhPegvHUGF9rtzOpJI+9uwwAye1T9wR1L3qAGXV
u+2+nvxjAPuvQaVpWS291MnSiMiMC0pAMSrO2VnKpxPeFLIu7N8MZV91AcSNkjhn
birBrcbTHI6cZ//zGacSewSTMDNIzazg2kP8/AFUyJpBm3v3vUMfN0Bt6IddBW+Y
onHab/mfVXnqxkEWDrVlIypBnVVTYgVGdkxDk20EXQJky+VziPR/RVOWV5hmjON1
M48eoUW02sd0SmZmqRImKfmY5dUmzWS1f4K44BxSppfrxwvzaNBRPCvlwAe4QtAB
063tvpTxd4W8vHXCO2rsqpEN4YqoFX0whdnxhYCMRnYnpU993NNkSjbGOEQoD/23
OtJVEens/Q2zGVLoXh+Gykeqo+v3EftiWJNxEAU/jdWZttZrwYbOfj2m3VU5aMti
tvI8UMRh/IK2ltgUMdUBEYp5ftI6Lnexo3yYgATT+T4f5cp1M2E0qVH4FStfL3Yu
71OO0jOO/y6AXmIo1PhpvyLJt6cATPOAAVVn5Mx0seCsG50rvLFy2lb00A4JVwX0
G/bGjJy52z/m4CXcrMH1tsA9OoD2RvsXEE5qvb9HJSsAuYX4Q+MoRdh8PR5Hs8YM
XjowfSIH75fTgtbN7ygjsHrdqp5EROM9kLp6RNLr5j3zXteIkmUVox4obzL/6CHl
JzTZ/zhr+jdRbRRt1Uk5pw==
`protect END_PROTECTED
