`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z3iSQs8C84pBFuqmHtdqp3jaD/m9nML6YjKpzEGAzfGQesstR+3AtBrwgnhvg4rW
Ad61Ev63vspr6+NEaLRd7M9KvXA8brkZ9ZRM7VVUybIK69EmCA1t2K0Kf3yNC1Rr
OJJfe3kesgTro7HPe4ppHkYQwhFlyowuTnkcopTPQtaF+PZw1Q+/LnFhzEdO5U3D
2xBvO/0NATnUhgpmxvbCnrw7Lqbl+ST5oz/CzQb5n3LIBabFf6CoU+JFdKJ6TAvV
UteqY0BjDLCOf0GvMIMTksbonnzIMtQSu+MNoFXz5VLZoiIKm0b0io8FZX+RyZga
7BVA37oWYRWZFQ9MeHPYCLG52trG7RUj3QqZ1p/XBvLYrjHOvYUQqTNIu1q5Hto1
C5BY+Ob1U4loBL4//EzQdJX64CoFHjNROXDnD9kahcTLM3RW56B24plxuE072o+l
7I1PI2tQ1rLYaNsNVoub/KWIRMjBiW5FjEX+9SDcbQtftiHQQiyNC35dxIdiTbGV
YG46ckp56PxAvYMHMFejXwjCqa6lrExPTNRlrX7LuO1FLFN2pjM6LJ6Z7MM59twy
NLy8nYgNrr7jl3zCg96+NxoyX/bFd+FFV23DXvrEDiv+8VVHEp6HfMsCThBPI4LR
`protect END_PROTECTED
