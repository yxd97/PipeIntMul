`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3idRIKdYSZmwEjOsgJ22YA+hyB9KuLgNwrsQ4GYmBuQCFyET6bhulC6dGd5Ycg4F
GI0rp9UG/g3F64eafdOyuO5asYex+zj8QrKVd74BDkZIaEErA9clbqTPcOxHYqHa
SXusR6b8OX/UjpGxmaFe3gpOLj3Xy6fStLpqYLtlCi4YA8mX7DHsQ1Q2T6YxEXiE
TWOogilUjRmxzYm2+1fn7G6U/lTZZP9ldbVehIdBIdFx7Pw9RobXC4kTqDuMVUpj
dDKt7wV6+WGzQsQo+KqXMo4iDlFF/d3hN/zRzj+8sQRxxFAnUgRhVm9QTch0OXkf
mCqPTqxgysvdb9zLv4yld7JiGZ/BI6ZjVLA+fPuMmUZCYzgIa04xZtct6+I3VhTe
Gx5pnFN0sWagS5fGK4F+KGn7mwfA4/3Z2EhIjdBIfB23iXalfim5JqVF0LxC8REz
KnrQNEnzDbFaEHbR2+ooNIUJiSFnekwnoOOiodb2PBHyKSo+NzvjYOOoDkmoPFyi
jWbHedwrscJy4XAnPJB8zaho1rvVARgtIww9ZXqZmiWUZSisI9vLHRhtW9TDkGEC
TPF8EaSNzNsWFT6vD+dC95IrhNYLSw2UeZKOXsjz0wDGfdY7wK8Jz/WT+Oc7SAMl
yJMr9SKCxRfx5GN7rq5Y773F2Yx5QW0/CBd/aazpVsA=
`protect END_PROTECTED
