`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lKG66eAVDauvlg2fZhDcXLqVIctWgu5RU6Gu/412yQfQrzRZPA1Q2dZY3k+USZX8
/i21+HrMEHeDTgk3hKWjRtbGrY1WfCFNpK9aZVENiKguxtr/Iha1ry/xgOELNZIx
n98L3yfaUknUiqrFr1M8R7VW0GTPT8PCtCfBH6vy+C+TedF5C8WT0N+gs7q+x3dG
vcLAKG2GGOB5eITzNjbaC2Yb++LFMC1TExgRaKVqNU9EWo/Jg7bPkbH/p8VBv2u2
Kd6AkcqYghsvceWVr6q6Ldhr8WFp3NHxE9AopLCuWxztoFvNYfQv9/K5f6cbQXV7
um6TFdevvckVQsoYKgR8vzH4nGZZR5sfFyPYwmn4rO1KCmQaO3wfcbn+Abpb9L/H
PGcuDGJCuxjvY7y5gzsWY2UXMPFLZPI6qcD7/jP4emKV4kz96b2agyaLmHCmkjki
Gy58u28seSvtn2vHjhbuihABqNe9ml+v4S7jVzTFvTe37HBeqGVdUaew0o9TZLDs
Gw61uC8ewCjx1yK8BwQSOqJpg0Y/1u8i+mBtViILl1dg84DQeZOBTiyb1r2UHKhQ
qBQ+CFOOGq28vwULG6XcI/DitOrfFc/vy2v3B41DDZ3NmyAZHQ22Ush77r2U2MAR
bWeDVjdHPw9qYYNKB5jjk3OLQBkM38A5yuTZc8awD8j/9SBSp1Awoyvtn84R5I7m
`protect END_PROTECTED
