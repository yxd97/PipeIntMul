`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EM9jUufnifUK7cPpeIB62y8Axnyw9ny87Q7iGwORDiOVwHh/gI5PkZ8PULZuVKCM
pvx6YZ5msWZenoKnTqr0P1Gq+C7CzalG5jXt36NupSTMBlXTqZ8tdsnA3B1MlLK3
vf8WwT3yKKK+uPTeKUSr/mz5DT97FDpSO+IqCpR41UvBW8tPTT3H/D9VoaU4pdba
tiS6DHkWUjH6fiMQz2VXhMXlQWJjq8SUTQnqQRo5k19JwSg478qE8lx0xPPmlMX4
cCnE1DTzcb0AVUtn/cc1Krb0yOtkNj1aB5pg8EEuHWU6q5A117j1G4/12B0lM+MO
m4oihaPY8MNW5xf3nZX5oA==
`protect END_PROTECTED
