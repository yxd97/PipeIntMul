`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
usZNP+3X+fcEB7QEZB4QgnVqwasvXDB09Xnx9W05C93LnwJkmk+pFx+tgcDQ0y7L
UGlxlDVqAZdu0zi7n9G20QywYXFLHGILo8P2igEOkQN9ZMuBEzSEVvpiuwa4odEz
Wpvg3uWxq7W7fZF68Rh3GoASqNfy0AdeO/imxzuP6TZqgGo8p4YAhtbKtqXe7u37
cN1f8aHKDg6bi4RmLpYi6iy5iPDJUSCEmhW4xfJQMETU4ERsG8b3Tpfn5D/EYKeq
9HLUSolHL0+v4FD39E2MBm9EGY8jvfFpGNGwj5Lea1FDegglAAuTANgnClKOjjMR
`protect END_PROTECTED
