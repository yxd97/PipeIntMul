`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqSXVrtYoKMr3/hDQFNevJ5YsmAI2IYZo4BV+55wlCMq66784fYmqvdL34HN9EMW
pBO2GnxqhwWZoam8DIry0mQwfvI4Kt+wYC/7KVrZgbGjCY0JlN4kINXMhAf8C4mY
zTZ6PbpRrARcmWd/Kd6ilEtLD3HToQWTQ99vvgLAR0Ax/p99OzDdPUJrpeufWyXa
G4r+XAM478c/UfqPSvm1ascPTLy7hsLSsYR1pQlQa+VS2tIPagg7yT2SYPWgyihD
+cyLYVix3Y/Z+BDcbnP294mouuroEV9/Nocyxu6OS+CqPWIWP50HnXwghejFmvY8
jRNTHwZ7pnUCRmpmCbIueUqc/+kEtGUdjtv416LGxXOf/esj85R5X2AUiqd2k5mH
lWuX7E9R71GKCZpT7C2TZYrYasXd66MoUsL/4Qj33JbbODDHkcbJvId0nje4LC0w
cEoEHHWmrLpfjXHV8SWEesbxaNBuv09g6pVJ2BfgCo2IOHz3iwOqMMLEPVMY8M7b
6xUG00G6dQ8HBMnuKQ/PpGnp+KFu1+64EqK0iOnRxf6VLnIPSKKr2QVobxPrypCW
KdqYbR5he7YhJEYfM5efbvgctZJAcpHvv9rGogDnP1GpWP/nDVtxijJt+Lz0Kow4
MSwE+vZ7KhQ0Wh4Ubf5enqMKiYE+IyHLZcL1KjqXZaZrMIl5pF2BWXv+I20uLgOb
J2oaBFson9YSbYQ8ODsupTMgaDNMcrP3cPw5T/n5nvo77DfTQcbA2dfVVrhyh2aO
fRbQ6AZhFMa2UOfpg9KmJII1P/40qBzmnQFEkBZpvWAdMFEw0z+fDCLKGkHyi1fG
wcOQ0EWK6PEt9/l44qm69U/9Vp5Ng1tGNFSepxKXWpf7VuPA5Ta1spp7/069Havc
ecQCurgJBfjJLnIlrYcbEexra56QKXVZcOZEwxvWKV1KYbP6h6RayZ8zv6cGcnJ5
iemc9dfOGKPjMArLEYipZgzOsO0GkhmhY5G+wgdOKGwjsv1e//JdpNa30fY+1LX7
rcdFu3GTh9YNPVNWl5gHOtVGVgo1gYeNX8bsQWJs4RAv7aPedEF4YmnbstNLAq0C
Lkw6Gh7VqCCyYbrmxctjyX05/2YgEdVO0RfY+I6e22w5WUpnJI4is1GnPAV22K+W
T57xWPQyAFZiMyNgmlrzzQ+scoTHL8KvN1irQyT1Jmau5iVPG3GKkhRc8um5Wz89
GqMNDLWbdzI8JKjjLLU5sBcd3BepdzuyWhFflegZtYspq8qRyMlC/GVU+G/UPS28
J+wvlDTOGB6hyx8KcWJHWHW19FSyLW1CVpMRbbGiU6/NNxZM8j/5v+aB4ynjCaeq
FVYjC5LEoWm0wIC8i01BNOcke0sHOH5fIVKM/RzIzrasIn+BbzzQZbWGqSlJ2Tc0
3kWG2mZCxZKw7fz57thSuKxSQkBvpurjGq3C1rKzViCDAnGo/rEbUvJe5ss0R0l1
e/WQPERenCSC/uPdbXtdsrUM4S5MwidXpyslO7T0RGiRS0TrRDf1sC2xFR9CJPPv
vpxHbbXvrEdu/Njg0lAaeqSWzpLe78AtPkznlXT3/6Ig0tl5ogONRfGtL0f2cdZq
klshJXPCZulf9116uEbmLsxeF2+gc2mIhgvHnE2imlLTFiupKsQAuyrGDzc6ARhm
qRNYNVpsyjH9ETd6uuL3T1XeY+h7wY0uAtNQSs1JGQHGpJiJlSZO/CM+KVmzoxss
uITgmWxaCUGmSxQI/5pb3wMZUIZRfdiIiDBlrBhqCf+UTZtKFwD7VhvDG+JLXwgW
onhvxrsVL96dNj+31epjRumWuAAQeBJNBLYPeCHkQK7uFtnL7x/FIhwm7jKiSNHC
+kyZ4sNmhXWsT8SvYeBfPKKW0L++avhNP9sXbqr4EZWrSQ7u9rir03NgOS8+956H
peOXRDcaOiwYZsPJINPB6FP0RP+oUlxZD48z8JvhYtD812sSq7+bGfhNK/M6M1PK
tu01OIPWP2Y9RRro9PNjrembIMZh8l2lmCEh06T4rUYqOeemqbymcxsNccGrH0Gr
964csS49k0tpGxin+k4etYYy+aGN6LnCudb0siaMD+Sk78NZhcFxzpTfDgK5hKob
96WnE8U+EzGNU3rafEdyZd0WuZU9pYW8HqEaxJLTJiBKOCgaEoV9tJDbRqiWZggw
D44UWyrdk9cov1Lslc5QgE/+mwchOWSCD7Xq+ur9kfL682jVUfLmcbwlYPvZqCjC
7IdurCLJC/KQsmBwtJoB0WAgrWPbVln2i/jUiKSnJjN76cTxF2vhGMA6YMDL6qEU
zeRkxwBrsAm/1A8E63q+o/Els1R2ldJG++/Ns3q91J1mDxj+Y1VYHvIFSxGP+irE
dckiOrHtBMYiYL4k0zo39Eg8wnKOwvbQUhufvAProPYxRxyG73NQw/VPwMVgd1aj
bkx4yWgihZxihckNQZ/eqBSYCxiHD4TT/Alrbj20UkaQmATy+59ghDQXh6sa+mK9
eyPHWL2yYFxcP9W6iH+/wF3QoAb7B5X0VXa+v7wws/OdTtk2rnumjwXwg2hGOz57
mbwxxOSxkk9doVCPbugNGFuMEmSjygC6VyxuDpFLjEoSxtVQSblNJRDy67VIp15L
Kg4d0MhXxiGbZo2IIRKCoci4ng7pTT0xe8CDcLnuRJRAtB60fY6Ii4J3nhAuZ8x+
oX+QGKOCY+QarodpPxzP8PLx28JR5Opj5iyO2TberZY7bbwkYVioZexSs6DnDwyn
Xy0QnhsHOB//gwwx0IwCgRL1p3QwNo3QKuOuOMojjxEccPVIuhhnKGPUTqzNfRCk
l5RpjvbLK5XGj0g4xwz1Tkttt+FyJr9jccF6OHp82sLAKfSVFWrE3qEm8mJGSBdZ
1FbcuXW3xJoRNmF5JoadV74fF6goeKX0/7vxjy9UCG1SZgazTb4XOuP2YI+K37H0
zyZL/l5AM3Y/JtwKohRdNZvs2vycuZuQFxBEmSnrVE5eDs3TMWy+C065aEUB3h4d
QKApPu8QDPA0NF5aZKSmsBD4mCqc9rHZdFVgAqbN1GQVcW0XnPe8FbobGUAhQXp1
oA1JMk1Mqj9Z28w0CHwFSU1EjCs1qW6+kZ8qkVuVB45DjBnmnwwK0CArfPEhAj9S
+mBn5Kahf7prdd9w15cSOE5KFZKWNNvNHXhUYbnsabZJI36z44W2YmawhAz6u2+X
JO3c7e3R9/r4HP+V22EFLJL8xXfEiH3prIG4jDxlfoEzqRHCD5YEGmQkypoeKxLB
X5Z09gj0ll2fvMSChxYQy61KPdCnGY7aYumoZX5GtKhv9VZz5BXHoSeTwfawqsxd
yU1Qh1bKyfJ5ZtRAlscFI9PbyXN+RZWOrdq4rvx3Cxk8NpF55fpM2JsEDKRc9Fv3
e6rA3eABPivoctgc73DQpyRklWstq5/SELNUGoQBkxqCqf8CFD+OBMic7vV218Xn
I3846uksO8K3zZpx1s0BJ9YLIOZmqqUs/qgAUiFKnJetwHQbapuYVDpcHGvfb2OO
eI+7nQp5GXydDdasccd+LuehYxfwZ4zqw8aTJwP2NaOzWVBEGCp+84JK5esAgRkI
+chotvcJZZzhtRzZ5xSdEIpWlGDOu6jgAf/QpGuYBWInvF8nkPZdJQ89n8aN4ySb
saGWbVFYIh9ebv/FrZHpj4kAYq10M6QkzOYqZDGJhlSCYP09vODbfMxBiswpqMpX
DAtZBUmKPvV6aTKacfvePqNG7lEQoxjVO9amVo8FdJk2YD0ezOtqF/DWtrG38BMQ
Jl6tSQKIl3uJq7uW/ymyHX3vbBP+/PBF9ZNkU9JSq8UtdMfmeNNAqxh02jGgsc7a
JzGvRGA0Uozf6S9lKVaOjpc5PNUnYeMb74PErQIRJ98839Q2IS3ZCEyA7F6SPUsw
gKwtyrns3GitG++vavwJUe1QOaCrxRKRUPkyCVo81Wc/CskRhJ8A0fdyLQggrLGc
hYGSL/BFufZpFWB8DtQE8h8D4VCM8TFiuDDV2PvAsEQFPbpHmLwuasrHpNvDLp/U
rA8e5Y3iuvPw8HDdcqWHxeR3YgPnCu+J3qHST1WUXkFZ1HE6zfHoSOiHGARsDYA8
xDev4ltfLpkjilRLnt1DYxGXQLnx5aS+iP73hAEAoleOUCEqUJS4zp55ZxI6A6ad
HZOC1pAIaVC/qVr9TMfAWquUFZ+cBuh+1La6UuKJ9BSZNbOqTsk60q8xO6+AzPV4
a4hn3ddO5kIzr22O03QmlB/8FmPkT7IA7+P3RQrMEN9wU7/AJaDwfpDwydHBvBBd
b8mzPuK5n9GPOqc6EExL2Ibj68KK7BrWUiHdCSqwin3JT1MySR+gJ1Gf8x60Z1FQ
BeTq1TWImdtBoYywgBrZeFBJYeOFipD9rsz7CmGkJNEqsQonWreGikVAq8BpB7Zq
LoW8XQbzrKVw5I49Y8wyHPBYcuzuJifXyLtABBDL3c7CtMoHux3RkuieHsUs/0NI
245/P1PG19HK8MvWClP/snn6FFfMIcfrrvT4lCtEjjZpzZwLNJ1LqexQtdcu/aQL
BXKve5OdQIViKBCbn6QXKftSHh40oyJ93dKIq+iWx5UQ0r5D/4ThZQTDrXtg9I2n
/0xEUwJqbtdXmg1evTvtOQv6AGXCLV0C9CTpvxkpSAMFiMAzUzTa6CRd2vbe4ulk
dzQyfy4NrdZ8hDoieMumLy8a66McoQn2dPyHDzPtfkfgr4F6lOIjCmuSoED2iUcd
yUhswf/9GjV2RKnST0VXhgjMEg09C4TRA+NiJcmt4u3PhhSuK7JyGnK2o8InLlQp
12GkEXhW+Tt/5dzy9om0MdgL7/MzQhLhTXQ5Fz8ZbAlyJG1MPJvwpQIG2nL6ETRI
SE0uQ6Cd31+EBU3WczT1TTR4ZU0/nX84/cjHTHFKg0y3518ct76FtEaQ7z20iwsb
T5cifuhgG1bN7sd0OQK5jGo+wwBR9QYS0UCOg89FLDAHbgp8ECbcIXT5wIMNPxYD
GiythTDX4zh1yzOKdwmNYOu0OHOFjgySux1kpkpI5QTVfmn3S7e/FzkXKtVcBUze
NFL42KnyjE2pWaB8rnEgC86kyuAXxLagQphyS5eoCLK8JbIPLwdQQNyejYEF5xSv
pbWlfqv6I7NNY6Pg513/Ea4Mv29iakRicgAKdpHVGI1iwQsbh6fOT/NiI07z3ytO
7mjezEIawRIr38rRL21Kv1M4gy++c8DCR3aNvKBL3ChuPJB3sTWm88UAnnrmJif+
Clu5/s8XAfBLydOh9ig7qtXhAn7WBxmaYjuOq8zxGO/X/bqMdLhIGaM+W7799nwq
r/gb+0CMWJNSAncmQixW8vCzCPBFCIa02FUZfzMEkIhZHYS2+fCmLAaP1RgNgn2S
+0ik0U5A4K9yFESVuNzUYByS5sSOP2u5f8QuD6OaRwBGMtTeyoPdiAzFmemC/6+k
x3szeMomHaC1m3Bu+QigJUtrC6/j84jLUUEvZSBTa+dqMsdnwOTcmTf+Jih6jjxn
m1VPQN+pRae8Io/n2FLkKr8STjagWkKRNYmOuxAsGlkejBgdyEZUWhTDqW/+u/T3
gOSucqo918rydgtT/Qkdz7WJBejqO7LqE/N83ULlivBOqc4tbzjDUFx4CIBuf46e
yYTjuwnPkJFnN6lZLksn/9bl30/kZe+qLK/wTy7J1sE8U2F5URxP9+HE7HKQR3Wq
MH+TaSX7qPAabWFn+MxSppmSpGqs6WUUO9BENlJnFOS5gBhk9EpokmdlRp1ud59x
E6wqArIN3FYdL+JbPT70b+gBjurFpuPaHNw+SC07huDvsgris8GNeqZU0hxv9zc2
BnVr9dyWKdRzK0p7+LYFMQTuoOo8UTETznUqBC1ovOazzURjkkuuICNKHBYRBiNp
LJl/cBEZDhwodCdJWKfIKi2zGeroZ/WguZ+LMiR9U8XrSZGpoBXl4NlGM7iFwXUX
ILu9NgDBlmDWSPUDf/haZZdtdGHKN3wDwc3zIqLsTVh9E1e1ibAf8vX1wkLG50Wf
16vA0xZl53CIvBvjJPo7RaYiJ2JyWjJlqrgsL0Ty7yoYi6xReJHHwF50YQzL+TQR
deM6ZtRzcNNJiGxwTFc2VdWeWzMqJTL7vnWGoBkqrxa/Ksn3CF9K4NDv01hiEZjI
+5npKerajBF194i6ZFyp7PCczA1h5bpC1Wy4J9eiqO0AlaecTv/8mZedzXsylA+d
lIysSYVryhhPMH6hteXL9WD3IpKBmqhIO3AjqKD86avtGehFTGcTi/0/+8D//Dx/
oLRaaNIQ4+4USUFuRQCIsZj9GtYNfIEtS8dPGHQ51UmGaalEAqKJss22yfaHYl2P
O+gBXZs4d0beVuBJ1fSlDo6YA/UXHB2xDTrL30oDk1zqgtHvPZgDLpaMBXgU3YYK
GlFnKBlmt7DKYeeQlHPV6ifYuaCam3JRiUQqaeuMr8xGCkeJip4/x+wzCipqqxC7
LkZ4D5Tqvzcu6Ru7qPW0mpaJBgR3TdIbpbxTeVaqKQFuK6nd5cG00HeM3kPvKgfJ
+rcozbGVFHDnSuYFO6eCu5VCHmIjSYmrF3OdQeEh2cZbgABzN6SoSKjQLul6MYLz
UUaiT3e+K6AacRMWr4QvcgYnJy7rtnXEoLxEp2o6lfjlgnvvR5jQ2308x6L12s2M
dGMequ6/NsAb90Uk63FQCTtiqkE3KNAFhFJwwVj7TrSoabAEr56Kd4kcsTwrHCtK
fVlR9rKhYuxVUq8DMczz89IWg214xnLobyFGFVENVtS8SwEqu1c9Qg6RPTc+qEmv
lv+KM+rFpXTo6HXnAdnHRfg0bpVaJi/UPHsnjpT+OcDy7p0TvWBFeTCHoH/42hbD
ZNN7sEInq2jlOpygq+BqK7k8trnOn+SE0wOvnGi+8Q/J0ZPyNd+J7bhnpkTT44cZ
psgfN+h67iwCEUixDGhZtBPIGXCFhdO9ZCIGAjBw51vsXa8j98Rt74OzMHuQpVnc
oXRZ2shbpBU4TTU5hHXeSZDfhUNSBabt/JHnsJHeVvTEnAV+Ss6p1xVbQ4QRKqSf
YYppa3oXM5Hg6i8cvquCJQpGopxOU1SvJ4JlP2yNn72hx2XB9UzrS3EAq07vWNoC
MqwJ62DzMNPzh8R1VqIL81NtGT/ct07wC9Wgjc5uKv72lbyI/2yc+yGx92D16PHQ
nqYEiHp9jYDHpi7fVSBw5gHGXbXnwMJB4WfiyZa7uCrOArm+88+RW9+lIZfwrMxi
yLPyM04lQWHx0nE+6h2IWqEW+S44kh4dDS3OkgIcUsdqD0KhIVQxdcNP7Spr5OG1
eVv+kYSAFS79/qcz8TfNSjjS6iVCJ5+jjixdISwKsI8vxMSRYsHNU6eIhgkIUYUg
VOZ6WLptZhP0jAL0jJ43vx+zdD+a4wYtv0NRwRkJkT1JA7Jw6jSTZSy6FDUVqGQ2
Kx/VbZpe0EGUxYl1od62C8hlMurTP3ub74wts6gOGh+KqhiypwDkeUSkPYG2kdC7
1ezpw/fjXVaW6/ZE9Y4nLybAcFzqANxyUQWMinv3JWlTaeGGFnM9STqfvFb+N6We
28itNYcIyvGjsWL3S1bVECFqaJti+iTT9CLpSBaTtn8znsiRChuJ6GkagGgH91x2
Co23weiK7c+icsmd+gbWAMZh+DQ3oXu4+NwWSirhnWbFNP/1agf4AxsEDOL8i3+p
I3m1HRyR1dHGOmIh8hEEEig1oc3Z4aqLNoVuAwDONaxrTfGT45zpT/WeM/0k8znG
RnICR2u8I0aGjrKzey6vA0jmAC9ivAV+2L0gL7TZ6Q+1FrtWD2wZ2AaGVCyEl5+N
+JaBTcMMnYLgit4cI7O6zYpu8TTKIP5zMS6yqIMUH9rmMSlhqeGYPtBBzieiC5Gb
9U85c+eF6eVJ1knFTyM3rl6l9AOLRPGm9+S+b2I9TEESPFScWLngQr81Lr6ntdVl
0iIG4G4FAGoAZy2omu9iEi8aVmgXQeSbhPEfkcH90Iah6J61gDk+pFaOVrXIumm0
7YM4U7xhHZ3XqKQMTDd+IJjqHwe4i9tRPENKwqRv55Oppx+Y5Zc1GPO70JfEW+/J
vf2e4g1s2GwlOw6zNGYP37anzJ993Gh02V84ex1nGGpYmDrRjCulYggesiPH/Gst
daXzkH+FicMb5sthglSSmVwjC2QJRcdpoSFbcU9fSgU544lDPVkXN6w1NtDoBof/
hUTM+X7zwkajk8NwcouVjhrig60quXFFswEX0tTt6Vh8ScBUuX+NNVmBziqioAR/
jMMD+UiVnNevzbTeOzCreZcpCRzeA6atcGJ/ZwF4m6VjQhYVhf3Swd6gd5LVLga7
iMrxeNPhYY6BjoG0/bMrK+EM06B2i5nIjePtA1vHuc1+4CO/z4lz0maJ6HUUGiM9
6LnE685bnNVqksaXwd1nX87xuvy7ckOHoM3lTY4DRoS0qPQ38mOyCEIE3W+4l7eA
O9F4ApxjE4O69JiTl5wcimS1AaLWVencxcnstRJbSNZY9XXIFz30QptZPyNynviK
FJc0wnD5jYCSdPUaAekict+CJUxBMvOzglBao70Phd3SVxPR3Akr5B+cEpKHQMAD
k+OGUYNkR3cJdk0O1ZOp+lMX9TNEOMdcIP5htXuNwV+YNdjzzcsdEfWVxJcROATD
RE1wpaGsAkiuJB1VPDEnMBZX1IXQ5y038M/7HwV7QYHFmkuoML6oq8yVDH4Z/NqN
7Kja0aGBmjPRdBlXZSGXXkuVfPfTr8cFy9Iffc+C9Auv+CL/iFdtUVrNEh0CFjee
uRzcNobRDH2TtaB3IuPM/r0RMsX0KHl6GCLFJLeoB+76QLoXu7DzZRV03+FIORCv
//78R/aBcOuRkxXZC9779CWZaxfP2liowo6SP8dZC9LLXB7JLHjfcOMPgmaoRoVJ
CIaiGn6RdTZAN94YYtrr2As5O/ok6lyauN5dVhHbcl0Ytt74VkDY1xnwDLTU/5BI
4tAyG+ezC003scgn5Fr7fiVvCWJNJSWoiawd6gWAeQcdEtXCVj4Njm52CNnjF+hM
XYL778A5oN3fp1+wKvvAg5vQtdLVh1eNwVH+kOXvbyzam6azW6cwpShROzzn6nkZ
1JxlQ3Q3Iu2krn6gkjUaBY7foRrLPxE0fLI4RTULGozln+7Ln8/oA4yH0B7CWpRK
MV4bDdsX+nRo3r7EpO+TuuJIWHK05sD8eo+9t1Zwl/a+DsfvdOe0/FDxJDCc3CCx
ZEMM6BDjH4tg5GILRy0g4p5YslygcNjNM6/YgJ9q4YhrupInwqOLohY/OwJTNFkh
n4HN9odSd5S24y6Oty/rfO1Gh9yi1raKxc5wPDVYo0QQRssf7e21s/dFNT4Uq5O0
Ik1rsGTrWS/SBXfeuwbf3+yZszhJpRzuAYd5DbbzyZh9+4b1Q5dqXmO+Zbibz7aa
TBRh40Wko5fUN5QSa4W8N0ru8IBMn8Om/3JzfU8Z/G9kRWzRxPzYtaNARKNhJysT
BYcUcI5M5vgpGYpwPN6v1hGX6XKEDnRK3mW04voi75ihJBekfS4cXEiTXaEg/xrA
77Xjit634+gGTmwF7r3azcVsxbDiww7lV7Gu7D0GFxKrAwvRe+UVuZ4CW8g74Wu3
qchil01Xgci9+K9ZAJY7LugxIIfBZ2YZL26GXynFcSUUktGiuaRSQFpSMOUtHGHI
5FRST/+Awg2GYDsqWixziTe5UI/2H0PEJNFy8ia5tk//b7/yJGw0H3kVEN+MJS98
LRIVxCrepRXYovV+VB8r02AYfXptvm6Lt+/RFOQhJzET1EPYZ330Ji9j9qBAd++f
k7eTPcrxj5Rd7xYc/9ZGPTq1MrNGGVTB5GMQCD1xRfUifeRs70yi3tZOzwRcG1gc
pvXfRpPczV3IrJrEt39lb23I+xQ7c7vJYNxe0f+2EjQJx25+Gl915zYLysStjtOi
QdjJ2DYUEeTumo2lBzONf3RjTE88U5hECVjkJIcsG3OMwqXgSMIne1rwaosGU53L
80RPxzG4ihAr9PTf+JJYeBImhLlE/9Rt9uZ7v1NLmxDNAUJo8H63HT/aHBmEeSIn
f6c69oZod4ZZPcuiVKmKtP59MkPCsIEil8S9q1N+P7DLbWwBPufPnVl0vo4feKXh
qju+tLWUrZQP1EaSLZVTuipeGNe56BuJUCalgTIK+GZI37vwgCM65w02h7o33Uf6
6PBqdfRHeQ+VqMxj0cSZ/nTvwdAdRJ1qJaE4p1odPW1tX1JlYnwxot/2rk9MNmbV
haCDqizPq4Ma4q9yobwOUIL/ww4DyvegN2rwrkyP8YmfbTHOOJ8RjktVZSn2fK5D
GIEmydUeifpbYx5LV4jEXWkNdlZ0OaPaK/DDwd5ynEtn4vnm15lBuWM44FgWazJl
whl5rlDaDrITbMCxCXIaSlktrv3ElwjNoKrlcM+ldK8DFtDJeAtIi2Ye7USfLd1p
ke2HI38IsNuoFIlSB/l1ZXK2dNyjGU/SvqLnN51b3HffS5jI6ozRUqQ7sT4BbolG
ogUQh12ATGajkAQyiwPgofoV6yaQKDRoOnSyBVjwO4X+fhlTBYzgPIhyuvsXQFs+
MepNzg0CdPxvpa2vzl26n7r1KErZRc+M0ZO3fQ0sx7/gYkfWpwPeamkgeoFRpXnx
yxX5Cvxg5d2NU6p3uI+n1N61Fg/Ri380yBkGoZvAwwdzOmzr0o1dUN032N0nHfg2
WGMzaWvyvIw4ZzOsqjHGYymKH3ULx8w846Mw7qr7oexn/lgIOXGTLMFpn+ZiFynR
T2Qo+uz57qqxsimWfkv80tT44QO3fsYlyJD1qhwEfZv2UlR+VxhGaR4HZmC+Z5d1
azEzAiLEHFCUBWmjumr6yRavBxtI0LFy9FppSXUP2BDSqNN7ADj5ztfoFx7AVSmc
fKtwJ+k7mn64lAUja8vuV5pHQFyswt0eZlMDPeRz1q+w9OIgfTF7rYSYycNBlL0g
euLzVA0zVD9GaVKk5Rn/fQaS/18FiuPwB2iJn2ydHc/QKxy569SFU+Zz8ZLj/TwX
/tyzX+QfxgBa/V/zHP7jlVjDzpr+VlzJcvK44AF7Lh/oze3lVRUaAAcWHYd3IBBc
NzxUsUom9d3I4U3sdu4Ric++GZ4meOw9eeobwS0PtZIydkf5ZcnPpqtvqnphzhmf
Qas6FoHlCGqMrlkHr0xcIPpgPSLd6EY3LFy5TTpKoHCZ6l15eDX8FE5Qb1MXcmmr
JxyTIn+pPgMTEP/JPr4ktsTKl3c8FVbZXb76czh7r1QnE+A4Fv5eUKvL8yApAqlG
fWsq9wOf93NN4G7ccPA2auv6e+vzME+cucihEq4j9jKUxS6ytw7gaE4YrVdK+6dR
hZRY3vtvkFLqRXywOFYIC7Id/wUXAc/w3Z0mzorkLxeif2i6PHrnUkwKk8qgFzvc
9x/8d/laCOd+q9j3GgTJsfbliZVJmbFfHqd4DuZYrBz81D2D+TxZF38Xtw4HwZfR
hHhzQA7B1/dE5rHb5ZHz5Ew11g0ILP3NufUJlLQZBoY1UTOouQk6hWkO6feuRGjy
sM4T3iaXh1/+u1rxT3wNtXFJF8EywDbn61KIDEpAHzoHF0C8W4MKA8sxcwjQxo2J
5h6z78p/qVRCHGJtjMLHoZwr2DxM+5AFT25vVySwfRDNBrQ/BJ3zytUhNuwwLZU/
QdOnKWiq0L1Gh9kztJWr/vnfApz+/DjbLwiMAIq3YYASfCGS5OKOczM6UotXk7Pt
XN+gfJbMvDZC2gshTJaYc3IYMLCoV1ARLcv8DNqvC11SCVZJctEe6bPNNymPFQ3t
8sEW495uqm11trhqxT3J78/yb+C22F3BboVE9EEx/3XLnjYW3yb0jFOyIHyL6mgx
8CTfwyE7yvWeImtsNiBD9/r6I+CPsnWmxASq/WCfS/DdhFz/o+M9qbMwNu3qKzF6
1ETsiG3SlIBOl1c3XADA9jHY+d/0tlgAyUKVDhmvgTtGL6zf9qEJ1VqICWJ1vVVc
Ld2hfP0KM8G6iVOa1WNwYLnv6iGFXl9JjSfhCysXanIWL7izLQsHhR0jEtOQUv3J
//iXy0kf2DP8A4KHGOat0zYH2ESnxjwPE8n1gr6OywU9E0AIO5uDqCYFyMtmAc+a
eO0i+pj5EiJG0ehBFQIBh163GTCCHJzA4HyIpSAOeQGMgHpBqIKEEr9YxzF6hxv4
GPzJV3hkT26MmvLsIBKCb4ev0o6uV9TnjDwbV8gGxY1+4E4fatD2+ia7RzPCdjS+
DpgxcNKfJZi2fJdPa8h5F1j0GqnrbMnJN2mYmIGJUnn06ymHsQKA1brqduMoAVxX
7DpdrTja0H2EXOq4ct6Epv12b5vfU/5nb4ZAFzHnPSg2qwSiJPRn3h3LXBrT0eNE
IsvoFyO0VucBO+eGaGP+YPaDjI6b0BmuJOemFzExzMzgE+RJFcYPQdAC4vOLa1+B
3mdkv+VERJEGFo34Xo013C38eFCaFoXFQEHH2tP9u6lIpDs/dpQ3+qlxs04eCmNS
kGSsSUbg5v4+M8erBapHBBC6dubiafNJuiM7sFX4C4OLoBaugjwJ5DnSfxoLMnAE
cGnOJiYSTWjRrGP3c0i19dpkL4Kt6J80KavhTEqCd5B9YDLSu2KipNchthe30Lur
hE9mFka/0SLE6iIwqnqG78i/V0K9UQtOrlEKRcA00MX9riXw0S7JAOt07LompwpC
pYFJ7zVJFEI5bxO1XY6UXLUYQSC6TLqSwCM9zMCWktlmh3l59VxUzdWwOXhXjipj
koHcZWO1BQ59XttF7EZfr/nzo2VBoM5H6S2pvwpiVmShsG9sFRa6rvi36VAGb7BV
cmEpZ71BumXX/zPFCr6fmMRvfGLXkkQjqFQwTgFnCsi24Cp7JBzC2BkevhHyi7iJ
R3vmQCeRjG7Efl6vQkBjL1UkS3NTH1kQd4XyPrtOUHs26PFM21wPIhpauNeZ+4gS
8FYHyguOS6eBDyizyZhgTJykslfcYHYY0Zb4ED5z8V2SmzwTBJw+lQ06SBRp4Rrw
2stvsP8XN1iv15GavaGwpOSakAxr2mJPMnVCJzpg2AxnOivrjOqh4ATMc8T4jol6
2+BVDpx4D3KDNOLVWr4NKxv5nDG2hFdghOYhpRNw1LlhlVhqHX522xFnlD+ecSsw
asJzOQYg8xaCzrRfFPEXqrvwRrGMwpvsg/cf0USWGDDt+hwqukVn7NtIIydnZjeq
x9khk50d/qqPOLrlh1LyycV8pzU65bnbXcqWhoPL9Kz0gjU2fQ9MjruCsrfIwSwR
PXyEyhwaeyU851Lvzr1vcLauHqZp13/q7TWpTlDk8rGD5MJs4TpNTKCk7SDGiYQf
5THYu4sCjisEr5WRl4ClTD8+EVrNjFXdHrFEC2Gd5jNE7pGhmsvTWxJ7ESg7pfpQ
cZO3rQmQP6Sb0tUS20s1PrzClt+Lz7vwmP6OTJyW4SAkOSwRXqQMW5xw1SFgzZPN
HkQfonWa5kWeO/D3XVF0BvoW5CpV9xP8Le4N6pjvibkMXo8SiyKPnL7HnYvK9bQf
caqKJVngVi+d2Ekkz6yVmIbY3x+rVffjDrlXcMYv5khVrcQdETAyLE89tiZblg5h
9pYAkqPuyCTxc6MiNRapLRIrWjnfV5msmvi/3DtLi3lLpKaahyq4JiMSYpESBpmn
/vPkovSXRFmL6dmVB6ISnjGLnFid/b9+ctgw+dGeiP5ISv1rHoIOq4qkDHoxo8wH
rTLzAl1Anwbh/sT3m/k6j6yGEG7vzEKpCLJk+Qi6d8AG5gyDvFLlU0TBYrXWCPZi
hR+ovl0UroSMNt+jKPER842wzki9ycPBHJ6pGLZM6WvbG/e5/6+rEcBXjotvT8R8
CYz9B2OVV4y/7eXvFg5hUuUxURkDuukdF5cCH/RT4kRGmLf1U6cwgZ/2LqDtJkZM
KJPiX41ffhLYB1muSI1wPNcK0TBl7EiTXO3QcX18L5ojNAHrNk1/4NptIrXThMpQ
520n2pR1RT+s0LsqGxiqBsMhX/Qczp09ZAkJ5aN0kKG4IWXY6bJxcVm9pEg4dw43
nHuw9zR1WDfYXySKM+vCTNFn4HpU/LV3H7njN4vUgiNLXQyJw9Kvl/8akA1NHEg/
ZfwPXFbw/uSwPBalGxOI0g99+U+KxHHg4oszqvXMUjqJ9mTz7vt1SoZvEjbOLzGi
JCtf69VPuMMy+y6mbMQptRVe2FVh7qCgWre4ehVjdeMh5tnr0MqBnpjUTC/JIrok
TFcGenA01eYg70BXeNQJFmeoLB+lSdb7hQKsn6WvVZZOdchDHMAdcCZTKnCz9Eyq
fgAbQo9YgYFzmxa8IBuSfdYFzKxp7o+cQyy+5tYWGz32f4nwkTX2WFpmCmxHuvut
XUnp39TBKTa0FrJBTYKukbNS+heZpWppmYKBorBF1gIQEAg8YsawsLBvhwJEuIDg
x6rug/H/yJaSztymLgf04bdZPgEC4xdvAynpxUzaxUZaSwENyrxXWjiXVYEr3Tje
VgKPTSrYFyhuiTH9qBRl0uDASVyvBD0UluCKrAUyU+iWWTjvrBPpkhL6aSRFuad9
SX3LIkRonuLNJNHnzdwx18OxNzsQPRRo/O+PkrGEuIOschY+BibNOzaLJC3RWTPr
E45ac4HuO0oWRsHFXW/ZNE2eo+gQ2l6dOGsiWCbN2lAJfyT+g4efhlXbBplUYZkI
Zsjb0wILPpviEtzE8ryd/E/82U8KA8wMJdgBtI4vxSwyLh5+KKR1AGEFQOSC9YB8
j8dejpFHsuy3cd8A0+xExMO7CNUf6xcB0oFXn94y2lyejTToMRQEM0pDsX/AZ+eC
gMLVatZ0LdbA0lQCm0nk4UJKa2Fv4OH5RLDmlm0ihY+ALVx+2Qm8J3+kcYvfDKQu
QOAf2DLhw1daDlvEYxESDFFmkCLz6sRFNnw4ODcrvI0pozsUdkfDs6x6yWy4/72+
6lQN9itADhzCfJ+feY83wnPPFBcu0ST4rGuDlcZYioh2KcIK2w4QEMd3jUCP5jTd
0AXJ3OK4SH7a+ltf00OgM3AWx2i9o+DKwnFOtACcqfXrvIWMq1Nw3p57RieqDw6k
soM+P5mPTc7hR8FQwGLh7VqW0q0W3R7HiY2WhR+ukM+n9Uz/OU7NzLmCFRaWI8jO
hFc0oOgpLO9ULLjKuKcj/d1k3cPeqojNSV5+7my9wKMJDhVQnBTTmICYPYNc4Xbf
WQX3LQZhn1UXnh/kMg9/mQ/Qb4UibQmb5sV0JohqfwnzCVl4/FkEn6rg076oO9Ad
ZFeMtgbdEHwjBffyDRsH4QxFwFZEZ62Ur/dE9G5hokILqviKKe/yxLSrfkPXezwz
7nw0C+Ypk/ARbvQsII/oOFWtepQVQbjN4paGoSYZ5rhVtH0CSUQAB9wRrjzr44Zq
/O4L/7ijYae4mKJREjTemBwRYlhP1M432v6QDDWXyO755uNj9/cn0GwWZ9OI+uBR
wxr12vhSCd0Ya78qWRMEsFJ4gNZ/jd2U/1p/fJlgL89ozsXwuYuMijkI7Inxq3l0
8Tjuxcs2HcdSw+ycNM7GkPWpPH7l4xGlKIo7FY0r4we9nxdEU8H76DEspKQOQEF6
Ic+LYUPiwv0hDzFbx+qli34T6EYPzub4HFZDBWZGApyWt4HkHJEasBYXRvXdU+4s
9ugY8UEM27NgcWwahXsF11NWuceT8+IP7epAh+OXDieY+PGzi/TmSo/d7qtz4F46
4HWrQJ4AnNBUSlXeKerSARsH93ItjcXouJgIqa+GsA57akPE74aCM2ZXiy89UZ3X
1DQzjjdSpb5ThbcrbbPY1GJtIg6CMQfUfXIF2NQMZw9mqmlthySaGZNbyY9mCNol
H01MQNAbVVvUmLCM087vt23dd8FB6gUak3gXupWEDOOMwZF63VVrVnQF2brXc4mz
rIcQiFexJ0l1eYcqjO3/5lwwy/ibgnKSblUM3Y0FlXbAMsT7Pt4EA5+h+pQqEcE4
u0UN6Qcq6RVVxPTbMfr/VSfBqeQquX3O9GJaSRU2Y4YGhmyFwAj3CGduzDF2rKxJ
yUSb2PQN+2N+GW9Xcm4DOWRugqnNxkOX1JbY1Nubt8KMQl7T0Tt7olmbV5bigExw
VfAASnrg13fd0NXNF+chEnbLReYW427WWt3OZgNkWbygmKG4HOEjq5dvB2+XndgW
K4L5QuTcZAiHCY73irYXBpN6bItS+vXj4CF0QtFJrI0vt4P1h9YCObZ+goWYAVSt
8DXCEJMjVT0QFiAbq70VVXaatjNKT8lzHdUdTsCxiYBP/sz0H/ixZ4WHuFBV7xze
rngngYgOyREJr8CHJz6UU2MB2eCBnLbmNGo91UG/sfsTPWGvmYtD9USzelKlFBXU
lPzo5GvbfDagl6H9sqe8sI2M6ZpsvBlhxXZvyOcwveBtEBftZu3tLNeGbt6XZJ/h
ah+rQQPWAlHLk3onvS5YhEK6eWrTtT5AhFmSlGSd3uXYhWiU2PubmEEzC7AgyYpO
P1nhjXnplT92T6W036c2fnvUuOiHO0N0yoKhj63i+l+chtFkSavGS/8HCrRlwp4o
vVcNspszfzO4HEC1y3bYSp5Bj2E4nZthrohSJhw+LsYyqe8gK5oYiN5Z4UEzhDUm
pjnkrh5p2EuvOWjvH9/nrhRlAzrCukHQUB9Gpmqu7fLa02pNHwmaaOTlmf+G8sXm
Bscm+yGtYGd8pxiVI30hIfvXsI3BE8GTX0DfFZ8h84PWTcPT10HqPSbyLrEdrR/L
G6OgbmPvYF2Ia74kxAWymSKCPV41JQDE7gyAPvfGt+iI54weo/dzeAo5u7zXtUu5
XqGwk0cch3ABdBkApwZD9tGKY34j5vVZMBth45IgyjiUcM/VpM/KHRBQqVH33iCZ
DnmSMgIMOepQJgP91V4L5A4ksnWW4B20Y32gfF6Id4SQUfZ6ypElsw/H4GMeEPTl
kdc1E0G8PK0RHX525dRxYBxq0tBvSckL7eDHq+sXpw9xOnC82pHRd1BIGZkltwmg
Gn1Vi/DHIwvZiWDGsTdqjaH/OhBqCT4yBb0nHWHfCeqYsyHquV3FQXZrjWXGNurH
rtEPRYMtbBYFc1MSspJ0SZlDM0Bk3Bd7drAFwI/+PoIGbQ1B5wv9fTr2XEz3EvkX
mtJAUvxerxzHk5y2f9ZeBHFV4z8/CvIa3zcW2AtO7DI1SSWNcmfTgeDpkxmnYoYS
WgiKQKIoSTutQDyRMXM3TxbcRQ8A9ONY/3gVgbzwkQEppzKcwC7YF0nh+NMXJKaP
sRc1ixwdZUL69SvTbkRvEj+7gDlZWuZMk3jAnPJyllauYbdaXgunoPA+57qffpY/
CGq6I1hJh1ABQ1k8Nfq7rtEZyCz9eUBvR9bRtREcVAJodAita2OLSqSpGvcnde4v
ZHceiVPe4rKkFfawVenfiXKEMYzOHDy543TyoLHj8OrD5dDHeF1NhnCNT7BeCgIz
u7gQ97hCMJfmZSWKwiAb74yrRQGCLxti9tFgZ8Mb4HqFCSS3OzPu19Gpyg8G6mim
oMIMh10rsW863SL2lWNtkVz1Iw1xjzSmtxtTi7muttjWO5q+oQ4NRd+Ty4h3+hAG
89/4rIacsIEfqNmL08+0SUSwSVzwzc4gLi6aYqtNDiV77F12uE90hTkIETDT/YYL
E+JKvjtLbz/bKZZN96OaDNcx+Xw4sO74pohfMpKaJ4XqDpqoBU2CJxWTEB6UZOZO
EFQvmoZJzOFFLcJo4rxyhJGNYSiX61IIfx6ox1g10rq74mYGl3rTdswQL23z73i7
q+/WS0XXnK+FlYdQDi9KyYunQOQ2a0TDT64ykpdEWHiMizbeUng65zX+De4t+7kB
1C2LynJuHyLsP9rA6+DNRnYw5rOLkB8CvkoTQ/zOyFhKEump7nk9Fb0ZV2ZuHZFj
YtkWGGyfBUfw4A7F7K/T3dRahuec00kdn/bjClXEfnOKI+VLD49nTTr0CEVlr7IF
Rk7eaNwFj2w75LJjWPpBuqvcQzvon+es4/Z3tH7ibw4AG4jR2f8FHGGXaufL+U/x
9gueXd/poOpFI/8ZP586F5igsF4p2mly0FEZtwri8az/zDkNI+rZCYnORzZc5pIp
eTTgt7gel2nRvLXq+ktSOokmo2IalpSSxDB/ng6dmN9UGVNqCB5k00HKa3GVoUrN
BTFzrry/x/p6YGGjNVTeeMI0t2qvJWYCsQfwn3yCyRJN/HOGfrYJojl0TfrzuNeI
ARRxe8Pe4vMRdExIxyAKl+DAm7NwTeXPAgs07Tm2RlSm6rKYjzEPZuSOj52p7Qu8
i7GYprw0F9mF9n6HDEuvwdUN9PgFtJvDi4UQ7VULlMhLuMGhHu/313HSnKy0yeCB
N5PshnfS9adOgI3W0PGBHAS9d8U75JXsTNs682+kMPUi4fthFngUGuo7Y8726gdM
1RoEU/80Q/0CNJ62bEdiIc8PzTv0ZXfSDH+rndYKSjpmAwXZhNjLO2dafqmXP8NW
sDOnmlX/evuwGSAvxOUKJwfpr56t0Qn86oJif5oFBBP4O17RdKZz4gS7PGhPYGps
2PFbqTLzag119slL3fV4Aleh+20ZriLhyvYQVQtBBpP66UNodYOFodgZ+8B0iKV0
9SMTGKe77NLAAJLtMF5chUgirIh7jpD8mLNx5HX9zdPGQcY6m4iTt3c0OQDrZF41
pCxKf41y06HKJjDNKdPXhuaL0MJ47v8OIMppmgU1EFU32yYFVtNpxIc1rC57pgkj
LG6dT+sjlNxeemiJjuvd3mg6ph/Q8ixmt6Yp1KMGYM8vVMLT0KuhO/rQ4X2GaEvY
JZT06H7zHaxHVrC76DCq5t173Rpz0zG8DswpLjW94j8NINL7Th/ceZugz/9GKvjF
d+hRJRgE1CN+V+/xPdJxUKjAibt6+nzJ45Zm7tpqfVWYsCJbFwdL8gTuSSxOb0FN
OmNw1KFPbbDC1LC7YJqB0oIRMOH29BhQggSNi+odREgv6AW4jJDH/Bg/q1rgdanr
SEKfcYWfSfvIpoJza7GJrK3QlnlQ2C35Dux+W1+lnpwUqwF9OtD2oqz7dF15mr3S
K3hMdTnmMG7bHIFm8yUpTBBPiAj9tZrnlDM+cDipx9c2GjpelHGGPXd02cZTTlWO
SjZL2l6GRtUGE1awm5CHUyvc0DFfMEvsD5QzhpWxG9CCAg9on4EeROujeC2i3nsb
zLVjKG2+2oeq7Ukr0dQ/7WwxXl7fEUxlqGCo8MkBP/iIVdiDit/ujENJR40J2+R7
FzO36N9nBoW9ISwZnPf2+hpBYg1/bemmp6tVNoStnZHs0Z0EHcHwxk/E1WiDbM4H
I4GsWYMHgjR9tj1HOGM6D8J1fyECpXowNMz6/URR24SfzrF7cC0/BgI0+nL1syEG
tzk9mwjy1x5cy/9EkQpxicDE484iCgbqZAtxnO3zZi03gDrRaujDQ8cyOSrXBwWa
GK9v5IgP2BjnukomCsOzs85LowRVeyXYZsXIqwPuuW2veEoqzNf+rwz/xcy0aoDy
DvhzWNXOwdWzB3FAhieOlKb2OBW75kwYLFg0TGmjzxE2Gnc30CkeWCXT1oMrOb81
IJK73aXUDY/D7sUdlOKuDZDDu759FZSuF5k0EIDhlGlSYTytFWPL/rzGslf1jU4K
s4115XseyM0zksp/EEb+1BPV2qJ254TcKaUHyaB8mgu9dySIqkO/qevQdjJShDwQ
erDkK1mRdKnBYALVU9tV6Ti/pCx7dWPCCmNbvSqdRtSyNzIvItUA6cW0Ov/aM+1n
zAHrEuG0sIYC+KWEoMPvPQ5xaPdSFfZgl+zDa9EbIKMlOdtpmvnNaL1rgzMLciMB
87Eff0CPKZXbGLzfYeUohzeGoiWPDjKjglknVYlW4buBCSw4y6fZW7+GdUWN2dJ8
WIDIb2G6oXkeeoVasFwEoSaGMtN6RiW+oRa1mxvoenO0xsOFSWFjkTktO7p7TySV
xQmOUkteAY/wcd1EMTINNCzfn6JrFguaplLuKVB/WVdR4mMXpQtG8F5m7lLm4QRg
Z/majh5ZWnZl1rKrno+NIA11w+GdkwJKnRVFt4DICuJDh9ntxXHsy/4O45disk/8
eq+Ul64UXoHQQvqjW7hGqzy6nNJaCFDX/yaShfilEvW3Cnw7wtyABfKBPtPJWQ6c
x2SnQTsYoQyW6X3XCVwDlaUH9/5oLwKT27dER4EDmrg/uNmuD/CUwn+va2lMAqFP
L/dzOPTI4j+ntbGn6Mxv3zJEnXoccR9puHAKHsUjjM7zsQ7zflwp3/6qLCuO9x/3
fILwfIBmUTDAupXcfp7B+ImSdb46LNxkfJbF+FWc+16T0ToCMv7bBGQBJndsGECO
PuC0JnXN8kOmDr4FK8PoW/jcoPgmLbgUGB9Asiq3AU0gcowXtqdXeU7tJhR/9aoV
nFxgEjQy8t59a7KJzpuKDKSYtEvERE7C9V3/1/rRfVksWVOCcfL+IfgbnCSCXuug
HSChlnMTFzGZ60XmyGNOQHk4CogDXbG6feGCgQ4CNKtKu8+VP3HMcUfrTKxczDmM
Ib9Kp2N5/83gRRwX85/K9fR6ND/7k13prKkL/CZBPYBhVHABkMFaaEmUxcU07+MZ
DOndu4wsfG2VdZlXrBNoUY1FqxmwGEaeICl45mkT+rjRJqKkyeR3eaJ0d5XOSwqO
NeS4KXqkZTsvTDM7I0EL+5Z4k61NXNTQ0Ud3jFRRuiOrxswFCDCL+j+qXS4GF8dH
Tkjdcq9TFnqLQRfbDehO0esOs6cw13uaMm6uCoASX5mPUt0lq9xMBZP2XGNyNqf+
uM8havyoQUAwoPQp6SdbIPef43ISukHG+Z+kZPBdXGClqabTy1JHYYRjEbmCbmzA
11xeLvxO47eWAn3uATWjXaZUMnczXyfVqmMhnA0mmSKVpSIAWXpPhXRhuWHAJKve
CrUtSX8+mrsz4MHXJGXzVWnN9UgUi4REygCNpmfkVL1tj8lXo2UoNsLpfVUQpvsf
mdG0Emy1W41zPZ2rllT2LJXfgEpm0IiE1jZZySpK+OnPbkJ0Sm4iUJfLlTnaEl1p
a1d2/vPcy2uPUl3D3bzmfslFCg70N9Epq8pA2lln06HpZDQ4rjXwIJvSpkM414G9
QinGAIKd1XN3O2bRvi0T295MsFR+kGqkYo1Jc0vujp3htWsBwU1VWh7TyKD3iCEM
1+VMq37nfWEkS+q9Dps7WdCqv8YjMBNixpdjujx/kozBcQukHL14PxiAR3DRVEOw
p2LQyyOimCkqvY6A0Zri/w+M6LSGt08aGQJMak+Eh/8tEp5JOJQA3BffNvsrSa6C
nIYNogrmIQe4A0nu2CCOlepgHdwr3/hnhTGvpcaTjgQYyI/BUgH3xUx4lIlQYV54
Hy1S0/ur2bxJyNFHGIaTD3PvdqJFOb/OTnqRN19jLMI18jVIQ/k20yun9VqbJ5FU
K5LQa15yZkQAoWnJJhguzeaVlRdDPZtfDJgmblOzAhgSeXmYrNgzbKYM5SaTFSjz
x/dFyWf4y3qP7L0AlkyJ/vYJN06W2w2CDaMDiMniYkcTLs+0T3+S/PlMMRmHXA0G
LspA0GzOCbUzqHvfO0ScaIrUj5HdakGQ4qLFgahBrTheck/6w4Zqx4wJJhximKha
d+Bfa8OeTV4C5WEgxfObXgARr6i3RcPUifrhquCxuRAxqMyVQuXDp3s2/4qfCYPf
+T/e/vW8uX2ntrq0ITAeGzDLzCoQ/6VJAmzFKtWu+I6Z/05RAeqIkKIXYJ0fHDb1
F4tUiF/P09GBeppGEcdYnPWIf2oU3L862C62A03EHkm6LHG8AZHwsaz3ZIBsW5vG
5UdqXtagATH3CeVJw1FuUDENnbSz+5MrRUaq8oaB1HBgZPZLR5pHIeYfU95Fwj7h
305ZNkfIyKKUGA7pMKeHUVEVeqe8ujSPzGkStiJqmfDiTl1Uctq4sfwrjL7wzWce
sVUVFhLW58R3P79U+ut1FGRPt73GCkknzPmRp23SPeYTOB0QKeyxH/ua894RUT4Z
DfGdhQdYkacRaxMofDtZx99raAy0xBNB9nyas6Fg3eK/ma2Vcc0mqQZufv3LQ/67
QyecqQfsBIh3y96Ln2KKjvcDTfGSg76WaSgsFRP7sWECPDSLmqZTXiMGsoZmL8qq
LWZK5ARfNxImJrenlIiGfdTgCwrljAwMdLZ9kfOxSj2Pu/npxJ5Bmwim/+4tcFkL
O6Q8O1v+uW5ssVtjS+TbQuKpwHfZPrrrWRFE+1ppQCYe5EqReWiEXTJLl7pPY0KH
pFX/qQ4BSUmDjU+cxeBAv6ZpEjrkz/1pVQ3CLnaHjQnxfHgHjCj4ivp1SA4GZ3N6
NWlbOltqw3VS5QO6BpzdPrnryuYlhhI7lzJLzCY29JLTPQC9fd8SwvMJM4mxdv9K
LwgufoDPl6hi/sdSVklb/eGI3aPJwDJ/3Z4+LTIOHFnWH3kUXVQvOtdTaKtzn9qT
6d3DB1XGgDrtb4BW8W5RBeqY3aHPbjsKARLH6rTrYl6Ok87sf2yOLhSX6jN0UTgd
wgFtJArR0QGVxo7Jzj98YUGd8gztsSNT/2yKfF/k4kP4vC5CgWq4U5ibphHh6Aki
e7/i2v8O+jWs1IkSPJiK1XWj1uDbwJbe6+4Mb/3FJGNQaZi7ZFGNmM1p9aN8g1g2
5x2nmqZyzXL5XG2rHQkknLzRhtdXAhLIpFVIaAnnnq3A0A8tZhWIwprrQePZZnlB
lqMv0fOPSfVD4V31/XCf/QJFIvZrGXdQOvIz2ufGoLqyTK3MCb07K/qig9a7AkU9
DEKlDObNIKYXczkUDWmw09a6dgXJe+0qTra9LfhyXo86bggYKEGf3EsaKjqArsc+
n+mveE8/OHJ+N4UsgoUROtSojpv38du1ZoIJx8D5nkNWNPK07g73jw5hEiC+UMQX
XY+U0vAC5UVetM89eaUdYeu8k3Cwz9dfIoaz21m04KIhNCNz0QniQD7pir8fCJnV
X5abzztKv03q5Dl5uUCjacwOdDlPku268b/c02lrPpJym9y6ZB0YoSomFhrH8n8c
yBbq511FbDSN8FUwA2ysT0eLc748yYRwG33+VbDeZlkmyYair9Gnk94rnvQXmhiv
YOiVt4pUGHVutV/QGLGd+5u4W1YjBoY6wzblul+9UiFQ0HHxxWY1bLpbF4fLCgh7
JDH3bz6cMW/anqvJ++KXix/gy38P7sbsXrLW1k/CyssUvfgG9Irc2ZKIw1+3FoGn
ef3Yt3iO+2fmtVkRBA3usafMhRLrVtnwlrmkTzzl2bILb2ns+saICEKQA5cxyhPi
qoOl8EQ8bd0wPAdJOK60zMZjKgpYiCOvEORw6A43gTVDSEheUtLPRvtr1mVXnage
IMyRm9Tw7/gJDIgQSMUPm9iOK3xCCwIBLBCiORE+cqIN9yBxouK2xkBdBxMNXUrz
4n8Nb7TXg4PsHLjY5BmnCDI42esnuIGX+8CPh2vdeTSm5Q5UvGpKM6DSXvNbkLN0
DVpGND7lJ6VlCV2t9quKyZ/PLO4EcXBCtWpfcguoX59ZVyvC8ciaR7EHlw/L6GVy
kLn/tN18891f3YLY4D8dwDWpF6dW/xyyX+7EHetuHkLkKu5n4UKUVjMhmMTT0Ctm
nj98JAdOngCFV1iBMTUqZzCSSUtEEWhoT/8OVkpoLHHWqqDjwLpsio0b6ZJtlgpa
/Bd2QtsQ+ai5yDrN6BsKGuOI3RtQE+MTVogW6nNo3+SPJD8CGG8cnwPhINb49Yqx
3Tz+QEa6u7gxJZuwlP0nV+66l8HeyVtBwtUfglJiT0yX237PbbIpb39QGVh8ymcE
6AWk4p8l67ES06DXZ3cBx8X80TZ6p1oBoWFeJmpd2v9BklFYOE/nnrBqSHLRMit2
Tm9Gm/ZDtIfNXK11+ngMdOwhmYhCbuQ9Sjo9ZseVzwzwHkQ+vJKIPaGijpID00lI
Ad+/8pWYDYl0KOuywD2h7CqYkYbOU4namwxfG1gzhD2O50uXzj4sn23XW56CKpxU
NqU8LayMCR9ZgQBtIwjOPecCDRr8Y0QiMMh+tbSHyN1810kiAwJJP98UGurFxwJa
cJrcdLqTfwKv9oW/a1Jnm81Mt9rOY6tS5AtvOp+nXbH4m2SD0Fd1yTdvJzoZ2+tv
r09obEVpXopnvC5f6fWfh389OgoRjdjegEZPypzlnVKk3VXPDb4pMayF0UdyGaaG
RuUOqMd5NX66ZG0idNhreX7AYsLybm+U8t/prTqaJBQLf1paL+swQZifRbOlwUK5
uFpzDn9uUATVddnf7XCKHt4YYP78FddUFiZXD4ZUr2YW2wzrBZ335ShviPiJF7Py
CN7OqChR4j0FSSY6M7CR2ICHxmnSUqCYzs2PxlPInyLi41VAIrt4mGjv5vTqR2Fo
ZM/kMGNGLrBWxd4uGD9JbpE/dyjcHu1xK2stuZOJNImfR0y3iwkJ3a/uwsv0azfy
K5+xznYLqJ3hNEj1wgWL6RyfWw9/ERwTYGkXmpR8Awo37ghJivnY/K9iM1wKqz/t
l/T58JIprWRnV6TIyPN4JrJkXjJ/StduaxzYp7xIK5bWaSg+t5LseAdTbJAO/cvc
B4NFzDlr7MMMSubgHuEeFNOzEXjAS6Z/MWzoOz1c0SPMsxG09SqBC4iy5BiiKM8q
LaS4IYvdJCkxd5N1z31nY0KXfBg01t8uJ7uZBv1nfivnydQl280tzTLC57czmtPx
8EIAXFBZMsgULiAXiIvoRuLuWcBrcUQZyb4zfzz5f6WEX9NjZbqOMfQ1e+Cxr1bP
b1QEBme/0F1AzEkMXadvYYyI5Ggh2TG5al7qkyFDUQyp1RbWO0blw7g0v+Pk7kbm
+zg7b8YwtSUlDx43HtjOJ6YxN0jbSzB48+67/0aP010ThehPnVuu8JNLrYqwNR4P
JCam1MHfHa1RHOWPkWbXa28nNAuwPf+HbRH7SVUSwp3UNraEh7cBsNNZHZPaeG3u
apELKH9A2IfEqSNgnxBYI2oOV44ykQBIr78Ly5ObGMo/W17UUPkJO0TRRstp7qi5
+tZ1M52kU6wioEwgQCgkm7IWUcRQZtYijbLi80MfoTdADuEo/2KacWLf587gvUpy
8Rzyyc0RYlP/5XbjZIt9DZ1AAchGbi5v33somwVkdap1xnQeUyr6eMPR3e0CYmL8
jRSvnT+jlIBNS+w0x5N/lX1TQ8oPnIFwx3hBvI5zPAesqpUF09jI8CbPYlhDU4aP
w/Ejx0MK+eC5SCIkse5yHw/38a5bkgy8aON/cX2jgSgUwC/EiKWk6b/wLPUO02aG
pi/iVfuV1tFxIzRR2C+6A1slHDE4CMPkPtG7cRQJld0rnTmdO2JSLMu/7GYI06nH
vfE327cZ51x6q1sXzcRX5mXLXI+lHKRJ0YN5YzwqZsfSMkKg9IRchooVR1eYooNE
E9JwofiNdxMdCPmTO6dChf+BJhs5Kx1cey+eJw7S+g0Hm1tTGcQhjfqm0oSv1duv
FY/l+a/GrdizidKF14P//ZOB6dcsaCfJKXSXtqyAsNa2WJzU4znM+Wx4ng//1g+e
4vavoJHiddTbP9R/OUxqHTYEM6s0owViE9WssN0tbw99tOnbVYQulKGp+zMZz7q6
mGFZPhprAcZXzk3GzO2tpS94xuot/N/OS92His2R0A4nqP0e1zDIQDaHbCv52ZSw
LhH26ZLASve6VOQ99ugQrj98mtG260z4k9o5n4Joo8fJBOlgAaiwSKQUKVii4us+
fHx4ZHDuSlxt+ayS51dBmaqAHVLUNnrGicIby4RLgv/qnK38GDtfFyL7B0zezevP
OQLPOJ9ef0VFvEZreNsb69q3QZryzwioOaNOUDNevDJBd/Tq8d1ISIhjaRiWPHiA
buzCrKtaRlJVpcmTMq0FZamA3sXLFa6W7j35Ibm8J+659Rj8S6IuB3VLWhOEzFog
O8Qbqpp/c56Q9Ct/LOjo2Uyx18MQErb5qGSrWu+e8IkPWCYwpw2HeQ/wfYYyKkGW
XQqUzBeYjOrEhzCGon25fcsE9NCLrY3vrZnnGj1Nhw4HoIj3mk7T+yoxRPOUbOxD
2vBnR5tGb9e3YBlo1mpRQHA4DCgs8dvsr72vBVl8EHoo+reZ9nNYJGPlxuFg0hHF
IeQUXXzDpyv7ltehedSpc8wIg2f2vuKy3LlrLWZ0yRVbL4FGcRJho5pevmjyRJ2P
5UAPI1uMHB+fWZwUNS1wjdCUkGHAlt7aPh97tEPLKzs7Gar7fveAj8SopZarTj3W
9vmKUTv081Wzjg9tlKLZRa8FdEJVhXBQxuaKoe3dy9baclgn+oH9ZWX650jNncrm
w4jJfpeEr7tKVfPHYPHnjGXGzB4+WNoLQ3/J+dczxUq5LNmX3D5WmgrMxXmLb2R0
9iAgP7YLdpAqYrxSLZDO+oRWrSdnVxS8lvfc1xOJtNziI+4obn7qCdxhrNfGElgJ
EWOwjF2ri2C5gljiu5/b8AmCChjwDhCGn7lcUDxieDHCotPQSWKcoxRBp4ScXQGp
61vTYYRiZmXQRSJUG+4v5DKwcaCCT7HEJog3vR9dskQ+KBl+U2awJWskjP/RhHsd
UKhePferI3LGcw8FOYEWKo+raxTC53/IQx0NVOEgw4+cax+jyZcWFBEOQw0gwWbq
lreaBaU0q6lnV8a2sRg+tNrLh6xNkVm1B5+6LHadksNBg36PXFbh/PwuQIT/Sppv
deFJ0OYMiN/iLav0b0DvAsHMK2MXHm8NqL2969r6NMpeSM/yqNCezVNgRQDqjo0K
kHeSFjXhRaGEN6JvuZZjLjOGowyg4BJa8bADAuHHyDHx/BSJ4YfPQMZfTheoJVs3
Q48o/UxeZwIxGc/bC6UDQn8Hd/xNOlT1cr17Rymmaah1KSEf5dhrZ1LJQlb+WoJy
Skh4tF1XN4ySmtGt11OeiTsPIb8pXY6/l1ZgM49dbOrd7jIVIV94v/8W37sqNlK5
vKux4cibyk8tO0ln8mMH+uIJ3+YgoPY5C2XKR0zYgEIk42t1cLiX2Tj009cHDdzr
j7+2LcrbWd0CzAd0hDDE1nT0C9bw1s9As7svM9RniPPrqEu8eILmspewoa/q25MR
GEuf5MjPjFNjjhnGzcBJ3Bn3I/9pkW89iko3/aq6uOrxCmVrNizvEg/5XKNqeAtn
5TZqpzUmVLQQ45HV0cZ57vMVheWRBNQ7vqAVChdP9s3nC99pqti+ogxk9EzlnMNe
5bTmxMHvvQ0XvhMWX55oI5tCTU83pwLR2271KSxicU/WUOva/rUnRQgOGkjws03F
13KDc/1XDb8UWgcvhZMpNqtAoPOc0z8YzKKfpTzKV/ZtOeTSoSYowYXsLtYBdBGr
GiKugWebkSpTYGMShl1lJS6MrLoov/9mNGlNndRmfGSXeVala9w8Cm6vMj/DebGk
stxdduqmT/+oqiqYe7hVv894TSQGgmKnVSw4wdU45DcrZ8utHsj3oTpu6oSVLKK9
Y/+TuWOVUMHabIhlUBYFFu8F+OmdaX05GpMAOHghO8lFAVnOBTZ2BHdKFa4Wi4Oc
XFFlrL6YfokA9gwkEvlg22itFGCuW3oX/Ig4mt9QqKUuVeoQj9v70eqOJVe6dxIy
4OKd5XsL/ulcoLvq9iVtr8WRShYOTgyx37DyfPYZZMmZeJ16uJU8c5FVEWNqJMlY
agRZ6l4jOaD44cNfPak0rduZEMWavP5iUheKvsefC6hWBreCvaDos7lYZnztPvfu
J0JbecOnXYc5a+uOJDGPSVKh9WEMI7905WgF4eim+o2Nsi3PRKUoyH61ZSN83bnd
3i+GudenLjlk3PRItQIrM3a13lKKXniYrvd/ttT9h1WsIE0U2KPMwkt0DkvOvg6T
dolBkMIZkRox1qk4ttr/hF/kwb6f3BcJNVGu+UroGfnLw1/sv1YASAewfscTYuSW
a8JI7h7gqso4uNgI5kybAXzj5yvP9jvWqU7wJXaaQ3MR4+EaTgRmApeo//I3igCd
faFs0MeTu2rLFD/cYeJEtWN1kl/j+nZ0n2nAJvkdaRcsbbBnX8nE6u70vryerAIT
xmpwJ1BcP74Ud4XY/yY1nTwoCAtIadRdZ+jIZ+fR94Utvo0EES+mti+JzgdNhmoJ
SkELK3nRv9sQC5VVtzbdTd8JRotFpK5K+44jX4KJw4sG5bxPXoBB5lwP7rGum7z7
gsVFh99u6g3hN57gYSbqlFDB5ZpqzJgAQj7EKnxaH5kBneNJG5ivzHUOxQeQDbf1
OgDXsRtJq6UOyMX4N2FXEWwyhZd2+PCtqnqfkXV5yaKxzcQ7S34E38/kYdSi/5Rn
5N9ZngTtKpp2Mc1fc5GSZHeuHT2viVYi9eaZatjwtU4/bXYkUwU3L/1bmD6iQXf5
a5EvgFQtTMZjWBYoyLQzjC5xU51nPv9jMcTu6x9cV81Jg3UYzZmf/zeP2gF0Rpu5
96vRMMDQVEahFYC3TT9w3uIdD5Xi8khBWOTnuc9jIJnBU4MC55s7qfC3inIW9Y3T
iSC74Evm4pMt5bvdUnprzLiGV2D9ZJliKO81lOz30ANvIVFLy/mOlZAYBnrceE7r
EeXAU/exdtWkFoQidG9ykdlvNmp9RqvN+NDlsBUPfzbH1qVBQkWBBhWiyGuzym4X
9+UXmivzqLRaXqu5DX1DvagG7hmZXX9XJ21PzPw6KBdc5A/jpveNqDxYZgLybTDW
AxawBF9dZaFpTXtaEZNEs85Q6ayvTupHHZLp+eZKgOkrEO9BACXlCRY5aJ+dMHkz
QJ9HiHG+xCbobZcFGMQn7BkIrPnRCuZwEt+pvUJTCWH+hTBtMLPN3bM/bfbUhSQq
KqneK0zUqohBA8sHslW+V+k65B16m8PjOkCPRwkgD3oEqfR1L3nVP+A7vKxXIO9D
GLmQbu5nKSNy/3iQqrLpDWEb6EPE9V/l2ahm84tY/X8InBMr4StWkK4nJh+jHZuE
cJqcJtFgkIwvHs69AmFM7P+YyX0Owqhhck1erH8C8kPHkdqNZipBsxy2YACQhLwj
f6rL3E5ikmg6XmASD0LMakmrqyVuEWhzY5kh0F/+pfvOabWANeCd2P1Nlw35NAeE
ACx06L9VXuCtUSHntB1qfSVBUq1FmNl6UXelyLMJCrhlpPyu/y8KpYX3AEcmhjZQ
UCRDUlKTu6UdM7b4e8LxL4Ok6zzE3B4V6ppv9ufi59ct/WyHJvJobSkT7L4OlRno
5lr0GbKQZQSndI1UNkIIEgCPJZnrVGO4xv3A78TBhWw1H7JJrZpKcMD05dWAbvbM
zDZvVH0OXDWA/DuXnu2cqtbXZC/HLBo8lDKs09aGnObLnjEmS+87u9xDOVh82ZM3
Fd4hwlNLHIa2Ii+o3IUDI3Cz6Gd2xWJ5BdRsuWMfzXdd6SShj6niP54pA+vjdFep
VVBh1JggE4X0afKCktTscSmodzgzZixZ1y4bnrvwCaAihEjqjUVhNzk5bteMFn0N
03bzcyD4w1n5QXa3ElICo1yD76Cp2D6IsFJKNWAUFIu9qVfSkLXqg87fs6Snzqg2
ZPB0zzUyG0sjy7Opq3czjYvjBGQX/4gRN3RgvFQcpkyswaUGbXpZj3qsTZ4tl8tb
zEqVqRbPvuclPywzfi6t3uGSZQP4EsesIoy6bNzJHeEw9e2SBNWc/ct+ZGNIGaVc
hAKFqRwY+XaqzdxJ+1vJf7scO6XFCu2GMcFv8WJJq/PDl6QMhiE7UMy/I+A/n72t
FgJV5Isl66M4Qo7z5XmKzd/wLypZBNxx/qW5CBPsOcEpdAxzU3kjwUSP2k9rTDrT
KAPsi+DKN9oadbN+uLw6m0zo38c1Fp8/uvXwlaqZQ9e7Fhg0y4KK+s+TUZHp3SRz
1WnBK45zqMKSkwl8r2uOOE4n8WV7CXxfYZkAeXShFcoc+1TDnEdcG4fDXLt6iDlP
XHJQcuFgnwHUdK1ksLBfSMd1v/7CR5l7WsN5Qqb73qdO1efhykdjAoS0leqU3PSI
IB0uGhtg6bf3yLq6xIHrjw+taM9DtVQCjSQ1TNHm+d6rk90tsbiayWJt/2sSUSum
wmRfDeWI0qJnqPKAHp6rLlscnqbDRcrkB+mADqQmjqZ/pCkha9UAF4MM9kHB8YXA
uyxTXDYEiQADbZVNKoUnQfq7al2sITv5xpBBuTIQfY581ZdHiyr+r5Qwl99J0zPo
pwxQd/6p9LojUWxk8fgvgUxCW0FXariVegx7SLtqYyJFOrpznjI9rIeZ+WWTZ/xj
8KZ74RFAau5zMfD51quv3/IX+i8TY2vuK6ijWFBUMCXj39aqAEj0rBdcGmJRbNAB
s+zUaWr8MgIenJ+OPWjKlgi7K3+2q9Fq18GbI7iEk11i3qPXYmLbiGcOoEh8EjSf
jhQN67pABewS8NdkhOXwy75OINKsL7nywRknnGrzOu42fSc+2iZyDHAWqJLlG7Ko
0kN6W2lZt0xnuHIEyMyCwJHQ8bP0CnTN3la1ITtymCvzhVFv1miGkp7gs3EPu+Qd
S+6kCLJR3NF62InVtzM0f6GQ4aFZWI0gBYCvBhQdimsEsY5hccJvuChQIkstUgxO
7TA0X6K7jVfN0a6+GfH7EREgodDcQW7ORkrBpyUcXUbJyzLcWa7Qs6442gxB2AHJ
SggVgwGSD5VMb4LiGuEfbuVmC/zBz/VdvGDP/tlTrMGt5BwTXXoqlO5Ru2ap0+Q2
AxsTM5lKypq6Dvp8tS9NfCH5OV/3we2z4fziVYPX8AWPAl5EywNXv5G7xJPziBzK
phttskQcO6iFJcpK2bQm9B66UGepMQsv8ioD9rTvU4e9z++aPtJp6nEL0TNh2uag
B0KiBAKhj2EAZ6juVMF2SfYxvlvIrb6fwJT2gitPul3tGOAQCmf49ECqXkFHrTqc
RdJ+0XdxKphs7RMlGjMaJnD/TYxq1YBcOkClRpb5/MDEnQNPZkatG0y0yKQWr2VG
Fh7boxaZobiNiVPofuBcrbCapC9Y4W9APpAqx3d88T3wcZ+gyaMmZustbCoshPL7
Jxj1fuYVIZLJUly7S/8Fb7d0ZppP8LA7tXlVCTQzqv8KH0c+o8SdI8HejtBNORh9
rDW3bHQ+otMEEhRuJhLQ7IAdjl5SZ6KRtNZl/qWnUFBJCDGgOO6Kq3Gs0EpcpSX6
d9mJcY8MCsN0H+YOD7wTrOQeqahNUwKUScNXk3yAlbXMdZ7u4N5D+SddVQu5Olf2
pTkgMjFgHJbXh7KZLsj3LDsvE2amipf7IT1Dwo3ITZE0T/QvjOIDquSG4aFGnGQt
OjbpPUWuufw/BCaOggc/t7uxPUgTNE8b4CAzztz02qCSQQ48wlVRVvLlhp/mtx3M
joDQf58MWbm9dTOK9C3ClQnpzU0Ek0T9ejhlCnGu3A3+IFKycPHVw4IAkG5VBkZZ
+i94UJB9xceyrNkVop0Du6lvUddbDcRcII2niHAFyek8yNIXJ29lAstjhC2LOMSV
zhYYhGpDTro+rO04kKChI9iNywx1uRlh07u7IcQHcBVR+4nFXpwZdsfRkNnMH6nO
nkFbSZFyj8JUpFERU8J1MuGZlyl891k3UQgAvc9FuZZAJwF1kT6urDBTyksTeX/x
cqGzRaheH0+U6mf5X51pvvdD91cW9O9DmYWPvtRFfW+mxw72/y6zj/5A7NH2S7nN
F1ml4E1K0dwHphhRLIbCqwF1mtycQ70kWquwGv58xo5DH99Aa0PSQQbh7u6cmBJX
I424JRykCAA+N31rtQ7OwwIdWvYWXdNCPSC2qZuqNwfNULOHMEEimrU1/TfA01t0
TnoXgWI+yBWjm2QhzvB2E42S50togzFXeAdRhdbLHxd4dLnbNfXzUkVnxj5Hj9/t
30R70ALILr8mpJirrUaa0YeYqlOOwUOTeiVS+wOIqfXd0RR2x+fx1ZU5HZyU58Yz
qUlMgnxl4x23nys4Hjt5BRdAGRJbKqh+uYBf8fkyYlW4nTquhveSylt60yI4Hc4U
F/PZeLGVPlVfgiYEFLIBSOTr0cZouVbCfjrxntQVFJ3SQqmrxtjDsckIUjB7cVnF
Rtj+UPZdkXGoIQXR4JegrHmeYCYaaY0ncRL3n6Nk9uM/UEnnawx1guJWi8+VtRMJ
vrHEN8JyFwx3EjafvT+YrdTrlpXzbFgMK5eQmrNPGVOGItyllO88hPvoNV/GuyyB
sruJcR8J83v2fAGdat+cAcWZoCrYQsM1f61fE10aXBI9Ia19ytT69DIJy+CyDQHK
SjutQVazr/wUvfJ6Z8rmUy1qI4AiXC2O9ON8OWBL4f472WRZ6/4TiiBuI5g+Rltg
397gUe1RKLr7/nv7ku0egYZBn3W772bUWgOI8i9T+V5muSXIhd5sHtvEap8iywpv
Al1+uQ98e/qT96NTErM3ZGcJKTLHaRQ7EXpjivZmaFaIW0ms4MuSPq8rMI17h5CC
uHWsXOcFo9XnTTRikJqQ0YxI9JMhft1MsCaj9sD02pWxHkvVraxvhxU391K9d5Vj
Yr1iMoBW0WsKbXPfktWMEl4C3Np8nMaec8rlDl3z5hvC4X5vTPteVueWfrVP+ptS
mzE9f/4VHWtHPZPa9YOz9OYuk03r3fRdefHoyiVicHG5hY9af6HH8WmakfU1CQfU
0YUVMtquxXM5pQDz8ifp8rGH4pI4KxeUlkcMDzSNiYwJNh2wjDiRTSU5yHSgh+r9
+QSUmWTeFNbLRhheatC8ujIMTFlRSfcCLg7/JeoOHN0iTgQbzax9kt/5t2JXEs2t
hyH+3LjT7rhT4HVgkobJQmkqcCtEtiT/SptAb3CD23DcAgf+lijkNyNDfW13edE+
K3AcZ9764X7XDsdApXg6hEE3jj4A5EJpNupJ0OHtMNPLdPNp01WByRihu02WFIaJ
esoHBQrpb8MBJX0qG8T7Wnj2/laXJFj1dWhQKxSfBNCrw0ut3eDXHdliLgDibVBr
AaHh44oGHHGV5xrCylaUo5H0w54hk+7poTY39i1SyOMykWB+7bf412LZRaNJb+9R
byujyCOY0dmkMftmpCt6L5nAleqmDYsiG+akOtGruJ15oifGh9XvFZBwBWQqxMLb
I6t2H/bG7FMXPJaaYFKgcalI5XYvEtQpFiA26LO/iJoLoo7m3ZgaojC/LEOr1ksA
fxcFsHQi7qyEoosX9brxiKgvH/XJlVXdqbGnuHe+q3jwgd3YQ2qYCefWv/jd5+BX
DtlLbafLvHkOa7EHHw23HnC7sf2Ssg0DYKptElshpIE5fUNpeFAyxaKR65b8ayBt
B31giluMvxJtGjXYYqoFzTUnAGA63i7uBZWGgulsD0fozY+mxJmjS5cPgkaRwYXf
lCkDBDhckNZleEhL/wCflfAY5B+3WIemu998+fnoADAjuHD0pF/oX3i9ql/pOE1e
8iGxJLc8lk/9FtrG57WmegruEG1OduhgwCXlZUP69/S/ydflPc5bYAg57jDjhJNo
V0xVNVNgKJgpehY+pMf91WN3pEij/cjmktZvdpFBBZ+fZZPd5R4V6I9RdFBxaq3/
+7vLlupmJH9pxaapW1zgLsSRmIZiuRbi6sDE1wkw+SGBvY4oUaKRw0cRQJr3I19n
XLS016tPT9Be3NMzSLDLxCQ7qDBruyH1v6iiYB5VZP/4Uw+SvzaYJu1qBfI+NNHe
LCqSso3cGnIcxlo5Rc5CcSFzyjNjwczgUw7H2flBvXHwxLtjdOAGdj35tu/3ERTy
pSrG9iAqYC0xA5XTjuLFs1vnGI8Uv9+I5qpbzyRUgilcmOMxNSiE7YsGIJzo+r0c
skAqJamvhZ+dTVFJEf6HlaNxclpW9ppQ0G85kqlpOKsok1FHRAIi9RjZ5TBaRb4I
kz9buqDzlQU/4q2jW4FqPQjuLQZE28wOzZdVobLvw0SNov/AjcmJCDlCENEMkEru
OT7AmXuyDAa2eEBtwC17J5CWAoDyBkaBin0TwxXiSFgJh8tzIpj1j25j5KjQW9wX
O3tdmOMTRQ5K0/JUjl2Fmjk4buY1N4bMp7og13hOZfM2TMGyhCUdblfldJFWWtS7
T9QutlA2TMEA4TFDw5DrcyWmQQN0To6wDwxDFiVVEFpnjvS2haIbFUgiuc1/Zpce
pSdwsGyGDLWF6kTtsA9zcU/DFXQVj9cBqBooRbLAqQf2DIQf3s9owa2n0uT2rhB2
QDyKJspV7t8I6vczxg4I3h6QJqXr35n294q9PalCwbVynx1JUGZs6v5W+reA7COr
w0jVHF9OFCv9gW/ZYMjQRU7zs2gTci/GFCr2pRPtRFLtqB/DDsDQLA/lMT0rRxNj
6x0jUkYvScOMxc4CAmPcVgKTMfszGugFAF8mqOSIi95fsBf1Kaf9gLpw0Ex5q71A
FNrmS+RlEHGZEFxTZxewX8rSUh9P0lnwJ71RBgl0w1I2w0iN3kIQdVdBKwlFVpiO
7ysPdJFDHlI3dZb1qcSVepOcK+ysrmDhUuIXw79wHGjiqsAMVnjfq1EftEGucbGk
lT/IDaGYekD1tyG8OtHGLyfAQ+vby8R+MACNoBj3FFZnHvB5J4TX4Ir5mGXrKSu5
0eM7a23myorKIWortREyZ59zALqZHPzkwvFMXsengDsJiLbEHL56Vg+bpeG44did
5KV1zg7T1Bf9NsPqQfM7zp+2sYFvWJqWi9qPw0gM/FCxRHkZwonZyK5jxGQ1XCkr
epMhVAuo4gnGcC16n0i3mIC1k/xqB6MwWcTneGJ47Rav9ZO1xAI7Hz0JpDspEQwv
2sHO9lcOxm2I1LIXxNuk0Sl2fw3S9UUVVeub7XB0MvtuThXqZ8zUeEvg6WWBOdRE
78c2Elr4mXDGCh3wi/NknWJ200tg20twXK/rLDl7LOQN0vCiP8rZfwcLKJWVVmYI
S7tvl3oM/YAs3+nITJ71Jc3tDDtOIk62/9l/6KCQCci1X88NzB+1jyS/wG/oW97N
XdAbIuZyI64qxmwiF73KZlAKlG4ifInyN13E0nWGxOr9Pb3zZs8bPIv/K8ziesBP
JZMUcQpPm5QN6iz3k8E/xe1mfxpmS/LhTIH0PZc6amKQir3huoiuO1K9pGPbJJ1Q
3x0dP2mnJGisuho9mVg0iiYisPCi78HJAwIihG5ETojs5wo23HMZc3HIVm6cTFl8
m/lDT0ZuU0CFLBI4THtT/VJVqGIK5cRMRWRnfAVA+a9c5WbtqvKlxjYpP6LKnrPj
UyVMyG8Swz0+ZdHaAnn9AAiGyMS1ixvj6kDutvKPsbNfppaGcMDvOrxXNkfvyJKG
zYDfuo3H2RoLX+4bMPr4+BeNd39IilWfvo08I3N6bUROcIl/Y+/pM91q/bgfS0+R
E43TMjG3qUHdyM4bcSh/jm/pKNAfJCUtp3lqa66fBCVQ8LZFR8cmKfD8XrStdjQL
7FeXzhmWBEr93HkAoZijoM41t6j6TpCrxKN9EvKxNwJ0SIh+ncLzMZoIrUSmLpjv
3KFrGCqreyJTSHyxZxz5K0hsTa+1yMdYis1Z+Cuy6Ea2tJj5nV6KR8ic6MZ9W4Dt
YaxSFqaeqR8N6TZVCLybOcIcabtOSRCojuCgbw2MDOd3h4aQ73CUkENlC9MrtXAp
dTkeQpUwGxspI1CsI/cxirmMXcyLEiQjMrPSGzUd68XIHjgoMGjjzHY+LdLQ3b3V
TOhpBDcGGjF8+anrBT9gWwupfidnrcEJ2mhZvumOH0O6yWOtwn46v0qtEZoSSSqD
AYLZS5NQ0WNY6EHSQGvVd0ldbWKzAuaSUPAl236Xc+V223TOKfhiBnMmIiulm6pq
0/ZW/JtUYDQOR+f4V3dmjn7oZGi5KhRFcXd5XX9vfhlILsiDz0iObD8ETfJ1+Wnl
2ViSeLrZDrioVNGjdNKIy9r4AM7tUnaINOgToEuct83IGx4Zx3vfqhbDw6WXcnK3
IZez4GaPy8Wy0NfLv4j9fZZZNuT4wkK+e0cqqtTad91cMQX/v9XHflS+I2Trg0IW
riipktgVi8LPz5WmZrfx8nMwebuRQeZUENVJxJiLIr1bIZ2P1FmG/NslO1SU4AXy
3qIJP1kp2PdX67TAm863j9fTg1rt3GBCCMbCt1oYAfjUEX84z8/WRhOiSjghbn9A
9lSZDKc4mpv23A5on0mXMRauDqMXwTWU3cd9AjJT3mppiVmCfQ+R7VCyoX9R7zlj
GiT2A4cuspX0seIJlgaZLSRXybNzySTH1SEN9As7kjSU6i1Qom4qQD+BirOBGGrp
SH57r4WLTxHLb+6G1TYsFJazawh0B7C9zKzPnr8i2EW428s6EOgTgmyVXFwqOObR
BmXu19ud1teKKvtYYWfThB6jwLrOTGEQYflk2/ZvjeTccE0RAmts+rEVmbZV7DK/
Ez345fVeVk3laep3tTnZt4ZbvMK3z8ht/blvDJwZegPh9ZV1R2H5+ek7n9XzF3SI
u+8lShLzIUOIRE+KGwjsMWmaeHKgB5dFLFHJ5QSUtJhqnH+xHzUllq8/0UBYn62Q
z/pHj1G9uhb+MafqFaUFuTEtEBDgq73uXYerOhzrsPY5144iV0t7DD/JXuwgI5mP
o9sOQjtDHpalrWucjYRnxcnmCsJrPvJLG31Bfei2eW6iRnNbq68mopncdDRtjLYl
kIZ8c9evuFx/dCk4Dd8xtIFZYPCRCSSIh/DCZzOYT3SV4tZr4PuXTMB7UL+RfQwX
qoHoacuSn4R83i5S8WkhatKPjLQ0OvD5q9QPKbTZ3tO8+qJcfa1NQJoJxakmgjn0
Dq6ybGLe9p6KJK6aoywEPdCsG9sE9cU8daQJHgnpyHsM5Iq1y/Qbi5QzdQlTMsVr
rW7OOL7vt2RLAt2d5wQUT5P22R2g7LLxb+KQ0kJEsb7nEj0iXt8a0H/8F33aNUVd
Y2c9+hHzX5l8L5451nr+5iWy+Gf8KZdHtmt1c+TXDz1XQpSA9ZftdQT5XFVpSnHU
/CPlJ/SKBG+p8dun1QLw7tCxfUHeO4r3XCVhSiDnInHilb/dZbHpPo1lr9BYZjrT
jCjXXlqpCo7FYWjPgc2qK8+S9s6/keJs1i4XWVhfZMKaRg5p4kvcrqzUKfIa+shm
mZL8os1w6jHmL5nXObVpLKhZtZZRTfUJl6S/IvBWCVEVWRG2BIYnQlOh4+/X2CI+
BK9C+SlQsxDg5t5zCqp/Hbvint/7LiLyQ7D6WutF4MV5wybhWdGIZEM1VW5vRzpG
qSLKsPupDBdC107r/5J3NQfkopr1AjPvN8AkkSg4HPrOcjbhJ8BYAmL41pNg7gKp
Ote7+CNVQte+Vj4Phn+jJ/32KdAcyYTpry5u7o27WVXSQIgtPDP0z+MiFdGaTzuZ
4/u8MFTGdrOC705BLTWXg+Wp+LJn9aqvQLktXCYGuMdb+xF5w2Z/qJYRAZdmmTmY
HMhfE/MVVF1NnQ6u1uTCA54fqriqReOzD7A/U2NdCV06pgfNlVBK8pkmTqFFKr4S
g8MYBIZVOGkqyVpyGc2n56b//r2dSOW0thN6QFlrUoEDgnjtJkY2h7veXI6QZ1qF
4lgGo+HetLBo5WJeLXnAuD02eQoq3PASao4/gt1dkjdbY5v3TPxzZO+WaUhGn7yt
SfxgGcy3bqaI5HxWNLcBjuCyHXm+fVvQqUBYzGIjA+vRwUTk+00KChEHPzFjBICN
YzFcA+LgM5ZvZdyM5nbaW2FtS7CwfX9x3H6ANZLBqcISXtdLVCmEi8iUdEIQiNw/
HOjKTmwqKD8ixocwiTGGyXMRSyoHnOYpSzAfHlP/UBHKlPB0O7Lp9BkfopcJerFZ
uTDr/J9IMR7SaMdycsdO48jpx0/M/fDEOaZMnsS301Popjcn3VOl68C8oAFRSBK8
gpd63xFbpdsU8pbEAOHuydYoatSyyKYzkmnWo4AKURqsMyCb4687HDYiZsPraZT0
7irqBmbgNcA7DmKdoNyvP5omPLgTwRRMVnVnQl+MlHSjEgsZbMsr6Zsqkj7qZRMG
94LZbi81LtfiYxLZSZEpE6OnwkGQAvTUUdv9nRiys3k7R+zeLaviIu/Ca8JA1I4b
kTiqZWI9KUobz9DphmXm/DEEFF6PJY3+YpjQlz4nePFHG+jtaFunPFEh9sm4n5Lk
6RbE3HbydCOW1qClkRrlIF1SuSsr8fn6FF+vafNoGsNIF/vB8kIPxEAFkNfKdFje
VvkGqUjf+fJygV6D4QvlPBEg1hWvJLl9piMx24GQ5vtOrTe0/9qMh/LEYbbe1Xoz
ET0xd9cDJRvsT8vi+bV4mM4GjFLNQuHvoauD3nvL4w2iOCSRj7FVpOBHnRDm/Rnb
kyIcTZ0GZcVtAq2nNFL+xsxOkE71x1I9ehKq6Dbaju1HZrqg2M0lne5IgdP1z0AT
qTTUFEsLdCu9yrCy9i9eX4ekOuFtbGnrarQSEzgz+JRt7ZcMKhpSfYfMIGed/hEK
vjuWQ78b0YGVyQI77FNeVaqQ4BBOSZjJjDBdiQ08VEXLS/X4GwCoP0Nu3T7s9+Ig
2ExCkCz61eX4zQMVjjjufCAGa1/9QeXpoosVWd2K8exKnEcP6wJmwzommtsux0m6
pHrLVKYR6BcbXGVratR31ZfdIfCCGSpNmqut6Nrkm4sZrNnT2x9CHN7NAKp96pJB
oegLeRZsxZzLW1YLBhThkGJXBPtf5qekB92ZUX4+4ZqMPEyOnd6nDpqTekRzBzjY
I52s3JRB0lYSIKQTwYGN7J6hz4HJoC+5uUDeT7qm/IAMnk1P2iLUAtPgVGgl/BCW
RPovJtFFfmNw+7NtByBaPECIhJm5DiGJoe6Lt8X1yJue+AkZ3HAH8IcNaS62jL2V
XQ7N5nSGl0L8oUAJqNBpNJqEDMhdJ+BWu43Xy2fdy3bqKADZm3q+08GvL4n3XmbV
caOTDasN+wkayLiIpdmJAT8WSwW4wtIU6cv7uCoiRuokKf3mObVV9OJ+9evDQZiD
qFCamEsAijzOYdPoAIbNK/ztK25YsNw8AX5nUxAR+oJW9oRyV6KwahsbqOGwROsq
bRZPm/eXyMPjZO4iDt/C+c7tWDlVs+UIOrnczTV03OGMplnCPWpZgXTq9Jtnhlu9
KGj+iv10KmHz8U/8kx0Ce4Dk3rpXpWgv5lp7frEBfGebHaPazOLmKchdkCkvtwvP
emDjJzAtk9TFR2LETT+6uDpMXpJob16TlzHNkE/Dz2Wxf1ywo+bfIKxoZDnRXJGr
WQ+Y6Ts9E2B4JF+gRYqDWov4afLwlIxVkkax9gqAEofEZV/kinQvew2Jva5TDdI8
DqWuPp5fusZshhY6B+z6JmbnLcpV+ILbVhUnQW3eKkTn4oCU0yNRQ5GrRUKerfiX
5IPhzsj52D1ra6W22jxnxXgvzJKo8pV/trkK1VoliVhrOcRyDVUGjCQkhjPf0BfD
lCzMpDOB8KvLrtN4KuhkiOoVFsMO+/zKugS3raC/ZYXthsXKpQlQ9VWKtRVXo+RX
ueXNo2e090mR2kNnmfBryHGG0fMqGk70+qnDP5cda0bINudjDnn6ets8UgzjP9Nt
LlZQQr0MtW/UBmlJoPYIgYOrHw4TFD6Z67rgHGfOFEUIjAmDait5DlkhD93Bmx0B
ZfPAM5+6IZN0LErfz6WowOciUn9kC6CHBvvZxljYVEpeXGSUysB07ffzUmElSN55
f1udHh8DyXzeeWowUo06Z2I7JaZM0RLiw4JzfXeWIl7FsTMEIbJCgU+r1CN07ulx
fjHp1AQ6xo/YuoT6tD7OjSV3amjSuYeYaGpm0nnK3MlDg4x0kwyEko4BjIANSMBq
w41vDmfIpqSbhMoQTgV92w7bfJuBat8cQ7w5QBQ0R9PfI1WW/REzN2Xd0Zmgdw7/
vKlmc623N3YVBAlyk0HzUnqHAJ4eJgTps2B9cgYDm7aJFnU9mr3UO4uEDdi7AQXO
Ug1XUDUoAxOGfZK3KvRaIIZDUcmXy1yxLKURH3kVJ+aAJuvIf/GLxGEjKBBmiYmt
vEjlXO+eaRR263db+o3ZbIQnUM7iWx2D7MCc6GXgLi8YJV/PaDCm2WjVFUuA8NTs
8oSqck1OPVvZVxeTZXOIaM0E6n1o4dtfA30EaTuLY6g7RirQBNxY+OoSzZOcfJHu
F+jm958Z6kDobC0QjqCvdjYat2FyWB0pJLXP11JKq4E5o2tvV8K3POntqx78yNJ9
WpcUNeVcX8Iggw9LJZ0q0jrhJSEaag220y2nwcbLFX+XdFB2ERrZjaorrTxdF+7q
sojesG2PO6OQEjcW5C3yFjASuIop5L+Oug6JSpTCv5CFacfmHHfJywcmfyMssrOW
Z5T83gLmppXPjpntd1g44o6FuZvqCn5CaIdoCg56mn1/Odv+bka8+NumfO/ncB5t
kcADHUkUr0ITmEgzL91r2jPpBoTmBVh4Cdq3mM7XWOtPrZ8Fsb05Or5EOZjSmM1F
cCSnap4oDaERZUWEQXCqZrXOPZMnx2ZfKvdrdLoWQxXNddYW4hI3zZyOcDcLddOB
PoYYHq1cy6bSA8Fg2MG5S4cHzX0Kee8IjjKjpYG1ekS21MXHUy5aGHgYF+QBbjTd
IxLuX3vOwrMNPlM+gEWpT0rR2bZlmV5bFqhrIS89zADs5JJQzd/2ybcJQ15bAT+P
v5/Mv41ppiIMn/dexwHt4Kq6G/gHzh9kbLoe9eBoc60HjWgSiYO6R0NvRJ8HHOUJ
+BazlDZb7P/FuyGSwNe1NpO2V8rqZ2FHK8EnZnecHcSB8hvszlru4gSnJFT/OAbY
+mpzs89pjFRICSIvPpPwVGL1E3aD9+/P0ozqjcncjUe4gERNqjT8lnxSnvfJT5PE
XBYjLSw3IpBItyLSxPSOJX2I7LTj3Oz7fS58tT82dSO5MASPFbQSduUYxlD61rpe
sRf38xED/FHzQQlrMPBxudK8MSQ9GuPOiCftXH26+r7o3CfccKzcHiEXVBX972HL
rLZMeJGxjATZcJr9sDUmi14MVsfB7VHkK2nqczL08+Czt8bB5a6dfsnmM2Eoi2Da
NnAYnLeAIlLlzkeem/eviVBmGR4e2n094EVFc24t6cbd6ryrfITtMlg9ik3G+qOq
qetHh7JDV8wrbKLDOtnPkd5JJW5CDxXdXvuIeG4itPC3u6xuzVHViBs9HzASQkcT
1X3AEIoU8JD6LXiOvxaTzDOvpodvXoW0iCYq9g8rH9aj0tfFPnsnaV6NmubvFqFd
Dpg/S3W8ZmFQOiOzTsZY+A3Gx5PMkPjwkxCQXMlPKfReMzXALBvA/1DV9IHx9BUL
2Offca6rjaBucliYyNWoBSHXvUGh2YxTyKGx8w00/um3R1e6GmrfYPgirq79O+Ly
9lFfCbpKx9OoS+6aFntJ8X+JdB0e7n11o+eAHZg/WhffBNCa7lHSor6LtwG14+JC
/+4xXcsuGORqDhf8VV4GCnnHyGkhhYRssexByVaApS3nR675IQYEyjhVlTQ9WOM3
E8iOWPdi/GXcJk1zB2ZM/Z92iJHmH08u9IkMawWup+bph1QMvrPvAL2kbed8q8Tc
DOcKfzHmcljTPaS7h1bBeScsWKeBTkKHlcuUznY1EPBjNWSA0BL50aEasaK1Dd+0
xwDuLxXblQBu9wTW2v+rdlNCpi60J3OUS9k+7gwaOgPs6LsNMdP302Gm3eZ6mYF+
7RbHD6WUa5oLQ+tbHlici+npc5yxkdKfklKrYtx/x37Pq1/9IedRP1xTxQQVk4e/
lvJeZqq/UiTqgWVA+9r31QkUeu7g5+SKMGhNdfZLTXsxLBkh0tnxR+astMeyp+MH
btLl8LIxwah4JWnpvcax+JfBanzM3xlmAf6brkUdHV7/OtUYVGPG5h1dJLy5GVW2
XgQYkgU1vzFQFCnrwWG6wOKmy3Qk1nIzMjJm8jUCvKVBtUenPWP0FzJ1oyry1rzS
EcXkIB1vcdZYQtZnBT7n2V6dF5U6ieHVk3h+EKa5HxwlFDy5dSL/2sC3P9QCwvoA
BCh1URFpRE9lpBJlVQIINr67hxc8jh93qVpcpZrwLJxsBfsmL13j8EU9qc2sF84o
Qh7MNyCKrI+50n7juulxOZLxri7wnTCsFCzQhLsV5xqKcDDaUVSDefH/DLel2fAW
ccHpyuX06aQ6PJSSKIVZB+QZTnIZ8KXzA/24SCASyt9LhOATOz/wnJwhAQ1XpgHy
Dwk0TWOYAbAl+Y5j/nBRC8oy0S6ZimvvSXCKq46gTu/A2lMl0hndo5+ZSEbLP4qc
cuAB1aK829EeLcNHEPfEfh/zdMFukU41ioyKaDHkoZmpMZz5VGnEA2AarYy7QvoF
f0XlgrhJDmjycqZ5XdoAtS9H1WOaHAjQhtq0J4cqcvpsJYDj8QbyGuARXcZkpHzt
m+CVbddIYnjvFzrf8oHUeAdDEbLVCLIlFMgRAjASzDoYxwao3CEKG73219mv1ELb
6eJxyH2upV67oDFa9LSFxWsDpu7KW2sU96fhiGItPEeIhHTHv92+EPU9IbasQEf+
dWeXTP5peTCXyt2A2E80qBY6k12d6ofCa8uNAYjOEHm2N0g6ec91PMolX/XppnL+
ondleLuWXwXk++LOZEl5kN01LV2ZCMSzDFBEbD7vQszVN+e90zGmyQviFc6VSsqX
Kf+63dg+OXESEPZeOtHyxVhfWyrtwznx3vROOXJc3ziazoASKTBtENHYAEVAjrdb
Wj4Xep+vwx0Fu+HQ1zK1w0dWc6B9JHRZEo6I2JHvV4T1zAvMpqWfXugN1OQsIBJj
Ni3t2zIzoDlskrZsar6tXnBLKDUuBGoG104d1numlmJMzUhwfXmvC7bmi0Xuzg6V
T7fTReo1trJwHSmVNYQn9RbisqQlIZGbEYD1AnZAATc5K8KrOEe0JHHdMrL+kwVv
hZLmJAYlJLw1n82UaebK4YlFlPvurMdSP+1XTDcj095or7uKlCGmGWYJ4pG4TXTM
w0DdeOyQfL/oUvpNKbIKS3Jp2+CDc4Bx3aKLx9VOqJBoWIS0obfw+xiw+qbP/9fo
upnLZBV1FFt/xTzqOzE15xNkNk8RPtjDoNhhGS3VUV0z7TOmkseBtk4nVVCUAF3G
5zyJb/QVZt/wE3ypmzBTADXmRTC4StLnnx/h/X4r4nR2bDFdsKOB3ThEs/7niryv
8RLwSGia/obHY6a/iLQ180uU+BjdRdb0r62scs2HPKqvxnqz/pIPBzijCs7u8XG8
LBWcDDlrwY1/JxqnzGMSRHtay7kx2o5E7kAySc7hgSIbdIZIMArnZOD/igNSAXFZ
MATtJ52ypf3GBtGdANfKPVGvU4GRTsRw8dpthjZhfxtyqROFrHnelh6UdY2YmBg0
0rAhkpulhNX6GXNzdRU8QPfbQ4Yo/mPMQvIb0wKv68Nx6nkTUpSYEF971ruyhkBp
ugGJoGu1BxBfKSWOTMNlAC4e8ylHpJ2fs9fxTYjacvwEecdgvDH/lxEOjbW/HFaK
iPX5/Q4FapWh0Fg9i/RiubUFRFF8nj70OrpH1vryaaSRYMqFOZZbLtww7ct3eaPh
331E7w4QMJ5PM3jdixo6u7RhReYvrWMZDuSTq5Uj+ZA/HLaCZ6JBttx4/0kaL2BX
eDjaq3JXxYkwbROXequprAmAOYrQ2WpLRuDSb+Ig7N3rVmHjWo5QSB6zRRJo8dAq
n7CeJUSejHe/DJH2A1LOvQn9t1aP4WAR8pU7Gl5wbrC27s5SiFzD6VkKkMIdL4+S
UWivbwbEAyNC6YkafiYqNZeF3fBHZeMn7bdhU8barNNk4yl5hjDJyf3HJvvHjO7e
8tAS42gBxKjFZUDeYcLzUUFr38UmSW5tNMLtBFK2LkFlL3VH4S28uKcjdttRpj3/
IFH4150wd9q3Op4/p0GrUQNKy9qxixelQ1ICiyRXcqR2gFNsiu36fKS8VSMZphzW
R2WOUcIgsjadSZl/l7PSiNoWT2SnQzU5xv0ewuDZkPZubLab2mF8xRnG2TAUfjxQ
FvT4O34HP53V4HWmBW1jNv5hkgnSnQdWOC5RCbfclEhqpUmYj4MUfKqB4Mbr1RsW
vkyh2cm3HaAI4ATzGM/HEm2WYcJJdZoXETFWdtF6B3SPeX5Tjz8ZVVl20qwHWKLc
yqEleQZhFlyihhIXIMPkhjFuF2euilQc5SVxG6+Sg+hNdeOhtkV4qcl/W9795s8X
Ca6rA6HImBRVk5bnZZ9xGRpE9eKxiUOpG6ZehtrD+FOupmTaEdbl+s8hDA4C6PHt
Agr+yoyfVxpFCNTDKQ9IGUnSsbkR+2AEnyYONHrfH4lgp8lXtml1SopWs2nlTq2C
gZeqpukrZbUDL2sYUGIMkdZdqwNcP/qXHudtqotOqHdd+3xCztOj0ABi/ppOUbWt
yuo6O9Gud+NQOCs45Vp8Z3zc0ISKjMDSyjtciwCuHWz6F7RiDZldSaAhLwqEZnWd
MFcW7Jf4igvB3hdpDJvrvb080FYQAy5R5Ze7XQwmxLrDdUXeUp4Xjehg/m/le0lB
clxKHm8iJrRI1FSK3iNBN5efTzSk+qfwrMVeJsFKzkB3BuWBYfyxULo9fSNZGjb9
kfNjoVb90QZ1JcYProyhkkTqLt4sVTik+BcNMc99Wf9eyxVxCSIhx9bvF6i5YSV/
6xMDovreSj0J21g/H+iCvEV++CnLIEqWqbJP8cPSX1X9mHMRVbQDWIkxPZxbOElw
BAewuNnAcR7XEI13f1ZmvukZuJMogln0LQAVa4R7K5uvAxPnSqFjyGcg0H7Mmjpq
bu6NAvCK75iArlCFNAFrHW0PcoTbnE+QlrQI3EDSoxM+Ln4gLQWgEY0OpGRr32A/
a15kbsf4rMjlsUrF1KqKJ2Rtrk0hdRuxyE6I0O3MB+o+RjZP5urSlE0at0f+sEiW
KabG3fGcAVCFKG6HI+HHc1r4u8XypkaaqsccUp8bmZnxa437K+wwvHz48eSs8WFs
QRh8SckVNMdpIIiyW7mbfCEf04pNXy0gES36TuDIdpMZ9LI58kL4ATTD5mlmW4qV
+rDaD2safrJyaXw9zI8F0zb4obYCU88atl8DrTceFdh90PgSdE8lUFW5oLa0ZMth
TRidpxNDl7e534ZOUp6Zm3h+4/Ud8ovs6K7CtRGPV2D3ET41WvT1MY3HFlmvUyHN
heB1HWj+Ve+spIxfj+BGy6CON+Igu56y6Z3fhSuHmNwk+uvj4EBcfZD4BJoTYZMV
0f4OvzM1dvIpd3qzDMcydTgFmlshDz1hriLIMPKUrTyHl2ySPu5DTEme+u5JZ9Bw
J5Ye14xHMlhGwHNRcIIHwNJ+qbMJfOUkIu0paTlMfiepmYMga4RDsDH6xsAaXT0O
+udLFDhB4Z+dEAM9K03stVlCrqxlnNYOOZDhO/hG0eRQogQDyBMSz+OK5B1KXI+h
tb1Tby0Dq8Ugq7Gp9hhBTV2LMNkXgf7v471qfxsIMdbg4fdqYefmB7ymdeNdqUhR
9S+mIeaOROqJsbQ0TSzB0EEvE8OXA8TGFnzDT9rCyKyEnLIqWz9hbojbemdLuHMw
ZmHRpFrtFmEQnpQ5CbBBQOShTlQd0Uiez0Wt6GmuCMuF4vtIV1cpFmwKqcYu553j
BrV+Cv8etmNCR4OhFF397HvFiem69owGsWrFNcNtAb5r4NqqV7iaiihvPUmOY/Cf
rxJ+8eSpCoYK7qYMVu96zSMngM84Mwhoqp+CcAEFJThYDIdHd5iKUh5qBUx2wKQ4
Rm+fm4aPSTbGaYxwLCjeMqhUJa7he5hzj1nbhF/trDOEPAPYYvQ7cDlBDAeyHlCq
15ub+v97IqCvuzs2P7fgPS/bo+8C3PnmAQV4UszQ7aa4HzadTIo0LyCkBw6CTXEd
bFmzXlr0uRBnUuXjy3erMB5lmQUa/iknTPee2khVe8Qkc7xVkHx1PLdfz6Wc80pE
T30FWPi0buwLs13ZBANL9XByBTH5Efrt15jwQYJWC9phrhRyHGOceff9zsr0vt8J
6x4n019peh8Ty3gIbVbpZ8KoJXAPEyAzhb6u5EGzrh6laLMGrVZLSlGXmtJH8eK0
oGOuQc6bXytFLDo0iueaBIGIjx5Zz6q7sXnp/EvCEiLrGHcyTe1pKkiinjnEiFM6
+/XuQN0w0sNYjFefAyeGYEn10jtRgVF5D/ND2xNP3upySS0FyqFjON4/P6p+98Cw
16PNzHr1rX/Pmb+/UVrX/bdc9hGJix46L7vwCCROLNxqUyGnf4IY2vje+QWUdO2D
4rrTCLSmvJdWq+cg4lXuiSzFCoo+xk7ZJghcKpzBY8GOj9VPqwDdwXBx2JP5Lk2I
N6ixiKY56YMwcjhCH4p1K14iD8qbOMei0vCJVTR7hNSCiFklvNtQx1vQP3by9a5U
uI+jv8cr3bZBaNAF26PibGCHFM3EFH9D3kIUkLPGOyn0KZo4cGotfQgtgaRIXBko
ucRCChv0Xk6OIC+ELaXiBMDhAepffUjMvluIdIE4hxM5QKyUjjufykHZFtLrWQ3j
BwihnrjOkGoNuL3h5lakegDJcadq+/mYXiLcV/m9m6vmI3A9ijwpsxaWI/9aooQG
BbIAkWj6FQMS3z9N9uKQz9ENile9HwDVd0rfP5DzOkk5pegb4e4k7N4K8nKM/3Sq
t12r5VTRM61O8hUnAQ4eZyTLLTUGEAWRGdx1iMIwd8jmFxv1eriV+CJXsJb5f8+s
pGbcoLm2JSW3Vl6dcSIbNjYlqhrh8E/wnCIgrZHQfGOUPycj9ILjrjeOxWu86v5X
wHjBfccsoxIyN2eQIgJxZk42R81b6+5JEdM/7OQ8B05IOxRi23JX6SY768VNXZK7
UjGFPye9A5F8nFkRU9dbZIRPp7f5J874uUP25lctGH8CcUllE7TFPYiryoqjggTa
1z2dL4QO0HwE0ABgS509tomkTGhLe+9aXVXiCV6+0bQW7olB/+OYqlH7IS+TEkf1
k0mc1Z1wSs4hdCyXKyl7YXJqx72efrt98RjoE7MoVbW/zCd8+D8xaWfYnWCcZpvA
+ieb0tPXhATJ1B2JiNg9D7KKEgZyCfKBdWl1q8SlNBIB0a8DJ9D+m/ig5lTWMSZU
V0Q7XVYZ3zJMya8eEb7eGigilCkeh17gMedoK2xCZ51uVU7uoAdDrWkpfdMXdxqD
QpE+vQS5ZzFPUP2s1BKfSXjj4ajNeq8uttaSDaNj6dzg0+LqMF4RieuvvTuZEKqH
j6n11ZmGWv1Cx7eoYer25XKu8AdBMhtcVH3EUphJD8D1pBrisqb7XIPi0OnUAK4K
V5eK4FzceXkjp2ievu6FgAGca0eVyC0DG0MWb1mdqCiRsV08cSbAYQsxVzssO0kb
1VWSYYYphU/l5vPmKYIiiECYbqPtDKVtdY1ewAoallj8VjLpBJmlWr4/1xlRKHey
Qfn4sjtKPlJ8N4GkrSFIGpZ+Y6QfmJQg/vylIsIvhGbXP7r5ed5HGpk5VWjLTAyb
9IW5I0QsFQvV9tfFhnK0V6EBARAFadLIpjCeId02+1xKo0KHS+t8TCIUPsSMX2Gx
y+YrQiMdJb5+tMK68ILxeBp1UMwycZ23yc67mTzZJ2kKSkhF8I9bGP7gcfX2tyjo
JbjrBbg6050+Hq101C/W+u4e+I9MkzzZbSUOsVtB+UMvPvp8IJHn1zG73Rstnunu
L7Dln3xPLgOi7vDH73ZxB+a7mhfcYCrAoyObIDUoWy/IOod80391bFXgtkvWDIRW
keaUM4LDdvntB5COcdxIwLrR/o8sRaUIWE0mFxAHXnF2/sIfvsLrt5/CflBLfgpP
aajtNtMVEgN3Xa9E1FsmhvAe6rXrYua7WmRQ1ub0xCsekWXNLvYGciO5D2VOsmOP
ybdwKHVquCNmIMIRsnzArSUk54hiIO+uEh/h1XRAGGy/Z7+h+5RXgFAkE2hw2Z5V
THNFNLK68uSL+lHHSoJ8SScCyFSH6Bml2vyE4fliX9L/MjIgeGN+xl8Tce/RFo/7
ro7BcytF7u11kl0+nXJMVP21z0SGnFqSJaml4VmvnIUQcjYjek16aVdAczYz0G4o
+itd45iEW/2SXKiqd1a5697hCkeme6I32GbfsFg7zkfYjKIFY9spqlr6z7hsWenH
OmExcTLzGX6FaRwLtV+wpTnj0OoB4IW7V50meXIFbPDeveTnFMbtN8plcLgb5qc+
soqZ+4JnWNYV+fNrX8HTh3LegPHXPYt5WtjcvSkaPH7Q31te2kj4tM3+L5IDVsOK
dlwZHIUDqZLm0QD5qNpuoEzCm5VoKu4ZCGUKXM7l7+uD2UlPYhxKa95V7Gb9pmvx
KtASDCRUKU4LFTJWoVqK7sYSf91FUDVSBxLM06YlDQutL8/Eo2FDliLlv2fOt8f/
9Jy2SkfAq5DxSfEwZB3jNThDiQLjpl4F3f02EnQ82BDvaex9Gpk/vxM0fJ4+yQef
NmSNU3RWkefkuBY7wRcynO9A6jD9+Ouh44x9XdCTGYhEdxOO75vXeyUPnMBWhnhs
xg7MX6WJQ17wJU8hxBD2t7HTLIsHvOnK/D+lqX92mtCaPM0/DDl0WtLBpYbznYey
1s65i7hkAlBbs20BfhimBc8Svr09li7xJOKqMS8Bm8LhGzbOncAk8hTVexPdH5Ll
Al4e2gORfrURDEC722kLnb0yGMDVxNer1KRQ7LToEOAkzaCYRUt/lmlgg+qbh9rs
vrKpoiufIPUY+LbpEvnqQITVbkbzRBYpXnCLBGapaf1PM4A2rmrvLV8ESMSrpue/
c3TWJDjuvlbYb9QczdLhaIHqhhYSXmJG9z8KjxQrqlLl+IADtgQTXSsjxkzLdXvl
xj+ZXOQotxnLnwPOXRKBWN3k53/QJvRBX8m2uISr35CMoJIj+0N71Ggtz/9SACUW
mrSjXIOaaK1p1FTroHy3S2z/xeyTbVQeDfYWfjfXJUv06+wunWH/JEyOWHvIXDxf
/QKFWX2fugzYjYf9om2IzpuUjTM4EsASejLd4NI8OdK0iu4YIyxcsXTzLYPy/5d3
y4YQ3FFK3a5zILW3C3ADVtDHSVuRLseZ1ifzH0YH0VYdUiGIzXX/cfg52GQJ7xVj
lOM5BtJNGc8Qper3EsG1Fzv18d5cvZGXo0Be7KiPl5k8okBmP4mH/+iX8s1dBGf+
nDDll+s52rZd6n63AsGozAQdIxB88mhBBT4zWGsi7cGhF8Ruh7KsXZVakspEctTw
8okiTtJEdwoiRmqmYoQ/tg12eUNp28+0KgrWbzlEigkyCaspXRcug9LZdO2zMtnl
7FCW5NuJ0wMaqoYe9TqjeDGj0HjG5Ng/5THGgOneU9fAst1khTPyIclVbLwfVQ9Z
JsA3czwLU2vXbopLL9dyB8kGdbEGZDUHACYeLHyYAZqYQXs2Lp5X7QHoDQe1IjnR
bAP68ldrh3Fa7zznVLdjHsxu16+4zUcogr1A9+G9Vj7lj72EBUHoX13FHO94T2I1
NuzVaypj89bvor/SHaP+QulVm74pGkZXloz3CUzKc4vWNXaAR7EH/nTey7kAL5Fc
vq8yvn29GguzgiemRMIy4CS/ixisbiu9HIu+MtmUaQCxVfhWGWLspxMjawfP2YL1
6g5e8TdPK2sMxAAWLxs/G+IsphglDFu9y5wWOklRC9KypXQbGR6tCCaKv2fxAY0f
R5OqlPyrOX+iDrzsQyNmK5ogj2kuBed9+Oe18wVswgwpjIL7sk1XI6v/w1OPpydJ
vO7TSQ9BWBxuvKTK8VK7kjgk0iHQAvULgWc6Lxq0DQm0ADNlyzseSFpXDFfMviDO
GGFlzJb/+E6DQlYS7Uhp/W4EaDONTiP2phckE2g7uF9D4+lmV61XT04TlvslzQpH
vEdanA5fexpWq38dG1IGUKAKTBjyKiOi+yoL7Vlvgb6Cq+1wQqLGLqSdNPrf5Y1Q
HCPJ0BuOSm5GkWg5hNKqtnQuYaBRwdwJp7UCQRUgBnag5HQc5T1U7MpntqRIIQo5
CnblAruFRgkq7dTB8WAmSFNCbs8dh21WQ/GwLYA8SlvescjPr5NbYtFlYMprtm/x
liKfCFRzR0NQm8nArpxO3vU5ImVIBKvfxXgyNEr7M/QoGirZ5GtrAOrxAsWBkA27
nQiXVQyAcCU3Neb8xmlF7pyq4ZnqsKD8FMz02cuPGvUT2zjayYRZ0FmCaaOs/dwq
dfP3JzlAMd5EVCMbruJi619e4orC5mS9ObziKDYEg8Y3/0JDw+d438wUwglPGhd9
Mp3cK/rZ2UOOPQgN/RLc8ot86NjMq4zRT1dMTG1ZM6qgh1bi1Wk+YEeBr2AYQA5w
eiGxQTcyVNkroX5bTUCMgk6gEABpD1oKp4Mq49g0jy9tHxcbuTRbVahi6CpVWXAx
DB97ZPZYAAKBhUS7HHGjJsQ4HGHkM+dUdJT3igoGKo+I1gbQNd6pyCA5jYgpgm17
inPbK/vGMW69aZgiBhgIOAi6TwlqL2z5Sm1qvjpmgiYWY1ilGcqMxYLLjSjEIHcw
CTakbyy8AIaswavZ/U6qw1m2o+F4iLSgaJUWcWps2jLLGpNXDNbHvOEXb811Jhh8
ccjit3+JnXFekk+FQCIqwBMGQ8uz/24qcc3M6Hg6I3vXqHtlxo3+rg32u+sECKFf
+Ttehb+klB88gh2Py+qdpYndc95JXEWBpX0+8Ica1dq4mQyNYJr629lfcXsTLVNc
OpF8/16FLYnPqrNyKAxPZym79v9+wauzjYxACFs5DxWOD/579kXoVh2UZMQDTsCY
n2N5u7cJhwfrODOefnpDOGv1GDcvLqDIBI5qUYB/9u6G8/VF5E01ImVnpsAOBGF2
7NR/0wGg+J5O7/uGPaxPw/GxUtUdyR4l39/RVtGUKfVbEHcFFUzyt5g2f/Ar0qhy
0jWprpfelcFZOfa7+716wQr0eXxQ00L/SqDZqQJCWcGQAOmYYmMWOzc95BnytUkv
l33pL4jCZ7LE5igDr58J5c1iPDGI1ZD3RL+kbtqgNxjBP79auqi82X1b5IjnZAPv
qMfE1BKWlW0X1MgI7P+ZdMslbo6xShTtbLByz8+Q7lCFVXCGt7ec/y8673anSoyA
GFcGN244e7Holh3JT+Oad1P6gPkkPgB4+lCv6QWRgbxLQ+zbRSi/zHuTJOkEjcQl
5/ZRIoaFJPNxzZbOUfzfyeUEAqX1HIYGUeXNBU2jE8ztP3HEqd4nrEn+wVP6e1eQ
DC4frihZD9c75Bewb7XP7JE0+poDafW4+7sc1/PFVG+hgxKYlOehbfeJwEtIby7/
SnuitCad7xkIxULxpU/PMXOUBEAFetBMUUgr3LoyUQyuGJlBLne32XxItinqzM4y
pbPWtkBdIArlV11uG0UImBNSxOW4T9KADc0ziWY+37eyrqaacM2qPaaVNXOA2CQy
2CJy05g8QUU0pkk7aSQgRAN5ve+papqzLCX4dGSzz5ni41AkWlwvZgm7JSLK0Ct7
qxiGzG1op0MIYhqfpGXQFu3yDCGejW2e0Yo3dWyFSmFPRCcXdRSczsEbEGYjg9//
IMmrZRC4cEw7IbkOU015+9LWD3KBu8h2TGYaSDaleESGPPa9C5vR7SNGg/WrlkTV
uElo6Xy6YF/sXHHlgf/vcJNJBsJ0o+LPh2EdziL1JUT7uN3IpcosiM6UhRvleBke
IsBRGeHankMHCVOCrLmWDdTlRTuz3Yq2cuofPL7Yc5IQVXi6GX8kk3fnP7XqrYAG
FWKj1MoI4z8UnvXf8tQ528VhmwCuibfcxeTRoEHRdTb5XRCsRsVWwkQ+QGh3SDL3
h+n90mRJ0pTJG4PvhtHA4S3wMDHfa/fBVp5d4J50YHw8KuFzPM3S6BlE/cxwnXMO
Jzaxmz1VWmQ33U6UVGEZqCCFuLEqZwvNDvL5MFGliErgtfYjkXcPKC0Hq5iCb3Uz
iJ28P1f9qqGtqEzrOfq+LTrRmUclF6R5nOvNvNfqXpNVqyswTjjMtzyXuV+ECBSk
UZWnmeQWbOsEmHfQsJC2nayM8ng2rXDd/ykNe1AH4N2/CPlDrp0td4h+ZZeUQxmo
iupzHZyxwClnw45VKX+71UKqngiLxuTdVvQwkbDZP4r3KXHwg6/7GOOqIReOmbSi
076m+yws/h1N0RnMGB8yiNs/NO57VadmTx1zooC6YCDJhwo7Mt+HRudQTMHLEbmI
QI7+iKtxYxJbCyoKYq6JxdSXhbCPJUdaKwKzt7RwDD0dC1BmnP0GZQtO7JJVJbLJ
6R1FFZp4fSZ4FjWGh4tg3XpjCkynpVr2ikDkurkwKqEp8fklC3eh4O8HQRsB1ML8
gs10SPh3UptjZGMak/1wRhouKTES8FAMySKMXV4H9KSJCGRHEI1YZfxb/caDxkAj
pyUrsyEk4h1YCMlzejnespjF5K4O9/Vm/EvF5qucuZE0bpNG8v1IF5+OAuuV62gr
E8foivy8+TxTfQjo38VD7Wzg7arm0XJot3t+zDn6OXYA/0bY9UJAI/bVP4UlK+I2
9M7eQoDQ9TrlHkaN75oVYGx7PrFWMM3eSGiwjzdT9C7ZcdgxD5D2yjpQKOQdESov
BlDeM4joBAH+Qa5GaQ4nKfkwEhCi4S3F/EAHuTTGAbbgmkYaKRUaHD361ARNa0/e
zkwYQ6u6tF9iyC1qlyrcwO7BeyK/ajvQyW0jfmamHE2m4yiqi2XhNwC0i2iH5kQ7
6QT6VdYG2CPYCV0eAvm3dwb6yjCbkH7XCSp43xkBoYb8fgdv0TBqeXKhlbDJkkBA
O8JRBCwfjw7S4iwN5Tk024z1WWY7OX/LWl8ViFr2wplylzYHXtTENQuvsteBxbQP
AdMOnIlLdhngTOM8ZK8e3L1DaezaH4tzc137PShpjUc/KxZMeiN5YuxNIofCx3qE
268/Oacag0X6jOmC+9a17fnoQ9Ib/pdEczYdpg3NyM7jPLY4e94U5EX8XoKdTMoQ
sFHjS/o4H+vfZfTCI8c/nAwptUujE6tn40QCJdDZj7a5Qy3VBe/B8cI9Azo1MT4F
xYwtq3eHFbN+VmpIZ1YSy1XTGzqbkQFkAHVpO7Tu2WVZnhKWW6dun7hlyPV39Osv
0fMbGHlaFwkDLYfIpKn1yqjfIJdMubhkiA7yV8pehEg63KXcbX0uuG6JCHdh9/9B
BquSCzIyUKfly0XzNWqT3dWKU87CMGyLFox6meHXl2qpnMMLmLh7LvSopO4T7IYL
yJfw+qDfGGx2eXe3yX56N2N5O9ymw7xmASOU7QxfAatO/3Z3gWq6t7mTlhs1BXyn
9Qx73P7P0OYYbDHP2CCZ5OO5gopOcLv7Ix1xVFrW3HRGN5yM8nOXJnSk5L+x63SY
JZfkFiDN/vdwDaFFCX6YEtn9g80qEKmH71ybkEuLfwVInfmASE+TiPyvO1Hc/FAp
u062Z9++Kp+RQYEmK76WwtBoGfRAI/07A2OLrCTGknUbSuFR7gc/qU3gWivArflU
6mn0xoEb6gWnjS0MCIRUPJaiHC+cBJggOR3fqnMMcM6HtGDkegEcZfGoCehBnuEL
+5S2nRaUxK6arxqkvhXoy7ay4u5BL9KlKR1E3SUEw7ueaT0P8XLfgfFiZV9F9Li8
V1iTFaYbqoO3fsNV0+0iiQzX+f8vHbJbrPPRYGBIBWmxFnK1SWc3GC7M4meaRqEu
wZBgoGcPgU2rFuowJFNnRMQI6v0JO5fSHgwDZOWvTGdd776dlS87ot5XxMxajati
XiuABdIDE56rLFSq40kKWXI/ZAwG6S1c1JOrekbb5/9sPzPa2jT0VlQfv+ZKQZdz
PCOy+ki7svNwAm0a8nxPXEStUAVsdPxQ8al/2iGOKJ7DXTui2VA7Xz0+w0otTAPp
h9vCmlvkV4LBdZisKcwogqoNGn4SocydprTEFSUKMYjYXa9TPIYvt+XFUcVxzk7k
fW7sEOHRuPYSRwpiAKCGytInl/DE6jTWHvHQkyFBJHwd6WI0h19PFq0GeiROwq8P
hgHkPx0q9TPBjmg/rQJ53Dtvz9FVx9sadWMmSbK94z/qbELW8JoL0jMPpAEvPX5t
lXDciHCR0cofrtBO91BtDlyDjW9Aw0mRpzHjKM4/L875qP2wyTN6e2apz9QyXrig
a+kDy8lLtfVbKE+C/Uym4vU6ENspAEURPqMBAb60vStk8+ASrnNeOLQ6wdvzcOZV
6P4Nf62O04cL44CTIxsA1li3N2N/T3mGSrdOERp+0ByG0TnpczHtGXpouKKvpXEn
TMQEcI5ZyiD2K+sKnx+4OSZ9qPglZLNHdBQCoTIkbkPl1X6xfhSujNu9acZfnBaH
/x1EbVJOWRWl+z+rPHWbRTTspV11pfWzDCrUz3jjemtTM9jYYUdX+Gy+2fOGX13C
aT5SLDQE5b89NeI0bIax4VL5nmweq18uGg0q8OtuFTZFahLTeyysUnuXXsFeXta+
ameZrSqfDwJtYcSPAAnGQL5/q3Wi/J/xz4hXS1w/djVS7yUxzyWbPWjVUtX7W4ef
7DpDH/xNWy+f6zRzOfuq5dJBBGVy/f+ORTI9VYp5LHN5n3Zp7mux1aZcO9iYOyX4
HjksMevk0CmUKfvj0y6MIbA2C4A8inhjOHAq953ksduVBxCPcgGHaqc1FIw1HXWp
cn4JS4K4+YREKegLHd2asmKUCsrutzPX6IW7PkZG88/rx423NDYM/35bXicl1Wmh
hFDkN83962VXWxQb+SBg2CVv08ZW2LXna714ju29myNRD86zYu2+beGo+ZZpGXnl
HypapKsAoGg/0hR/7GTg6vZf9pQeFWmTKB8sqAqxVVi6GtCWo8zzQnHEQE81MT2B
P6gbIS755zENHoH6pC5rc5WwjpjlRwqFjdOCtmhdXrH6C+t4GyuC4K//HdpgFFUo
fdzHorBwqhk8JI2jpPbzs8dkHrE01YpS+xEl8GU0sd9gaQZq2DM0okBTqtl2Zyxb
jrYoIU/k8IyLS/6snyeQtxWzfy5k/ZOVWZtRS7wL3GOMAahmnQVCYzD39+77ocKZ
owQrDri0QANcEWlPOBKm9f5ZyEQm4o6lkz5+uhFgKFbA5g/5bH+R6juyBO/WdVZk
Pw/EPFh4soBekCeCPefOr0X6F5nmzfpJdbNu5plrlAccOD/hDc/jREldeNkitEoP
CfV+oXU9HD63NyetEqO1vckoyRAHX099Y6BdfvGaJZ2QO/VOpkGznT8GBmRyi1ma
lK0pI8EDM2L0wzY+GAGSNIKMscC/hC8KRHZGT2muwVKt89M5I8D16NfBBDAopbhd
/meednGdvzQc8roEExBzVCyyKQniV9oVanQO9ruHOJbQtj/EDR7m2+pj6lvKibY3
ROzMy++YH66PcvUyo/M1n4MGUvBjCUQKMBNJr40zMlQLEqZYyr7bx9AHrwxOV+R3
RY25cuKd3NIuPe5u21lX0XBlXPkuboQpxVo3nI7fOBtDfBT5DZp1tbMQZz3Fv5SO
hU//qtEnY3Js0xIUfXK4NaG8j4koerjUBmTrRdRWkJvmgHqVLibx0WrK6Q5Gt581
M4sLQrlMstP8zYsRCeSZ1/UKlqF81uGRjk95xQEY+nIAJNNuYC4ahzyJRYFDkKM4
1UOwziteD2vmMmrHkvT8wP4OhjVJkiIhtOUvYiAP7lnInrT6yIHtq0Ge4NtXT1Jp
hQKbrBgwCTOpZ38WbJD1Z4bwTE3EQnPq+vs+ayEnQ0yDEbObAY4tGpbmoIvLt68u
B/m8gNcTIxImKrBFjJCXGeCw6d2tG99QRJVk3LXp9Gij8TDTFcKFeIT4np6THEPy
votCW/cshgSrZvBG+qN1andBM3jzK/Tpp3S19jCd8Q9hBcrpqouBUoWw1TpREceZ
pO0iWVRt9mdr7JJkKQ3s33k/31s5tJQNWcY8XRifhoj4jOiIcBGBS+r/k+XKtUuO
Sp1hVMuf4MzRts+2/D7gCITA3rPe1qBizl/wAAqoEwN/w50DzczP7p93m3I92a0E
YzGJfKyR2cH8Lj0Z9aR1TH/svEOeNVEogmnO5+8k7OHglKf5HjrnoWmzuFkOArbk
n9k4eOZiyjZNpbGH8EL6u/g2WSMHcSeoarhfYdVCFa8sss3LR7yCmZ/BoQexqZfA
nOkwSo4UMS3YYt6yDGmsMA5bVCNY9ZIxbsa7mQG21BQgdQn4c/ccVLnqnohBHBFz
PD+j/DgrJmrHg6r1SXxL5vaSje+9ivqXdNDIGrh4yiyL0NyJy+oHYStn4Bo0nbph
ed9NkHucDJxtnp9DlEeITBKacpXFTp33tKL50AjIrgXbosDkbPHHne76hVHYvbqX
LWyO7dXZeK5ZD99aIsU//+E69+kX3jJanXsftmrA7tL3KRuVaEkSn5U314YwY+yG
yXBinSC/OzjcWgvD1mZsm3gN0+E8vI0nRVMG/jiCayGN2xUUzKMajlLXmEkryyd0
uL0BnIonM/UoC2XyioM9x2tkckB6D5LVg/F6F9EjoORWEQnFhnyW9W3Q+s2v8XKg
05lFRWTzkAucgFcbc+pp2At1c1GT6HTkrGS4/sZTd74X3MJPLS0afbDS1rmI8ef5
76wWLIQrCHMDkSCvXaJXGN8Y1gqCb5VFbEqQo8kQ5R6aq0x8K0lvJqM9ShwqlG+c
SyCIhL22c00yIQbJt9pTdVITfTwJ3SMlI+seVicuy/cXJDzLkrkFQv6I5lxSU11t
/3+/QomLABNEqbMr6Pe4S0xqEuSfUZlHJw6fPmgaPl5FJc3XtE70Vi+tH0yIt2VL
NarO39e/eRkdA+YLZi4Edr9417ZyFRFikg1UJ9cT5xDJos/+6E3pNDLDQAtAT9uu
5blxQpAAoZoLZI9Qd7vlgjpRXKP6FTWOxcYdOkPxmpUUd6ZtnbZpTdXYMDunl2rB
eVARnqujY39Rqhd3PXVlT/po+CIrNVUdjxps4G3nK+HuKnZyR40DTPDgViCP48kK
C/FIJ7b5Eg+SAMjuKmrunOiUdvEESz2xucE8SoMEi1PpwZVv0AAJGnknTD5KGlgf
+6L8LOBfmIp67NKb3tRx+Am24By6zDNGVo+bWMyTY6l0AB+Ud2CBNbiJ5MAUtZOX
qqgDOtAFklLekhxYwJZ8K4EjVJ3uizccCdw8igQTA8HODpCV78muGUFqn0LhiYO5
5EdxiCiOTJxdZqkoJ9mRne12bEmiiPwxQSdapwRyeGXPIp/qFtm86mAu0iapZLIe
RMnmc8NlILP7SebMh11G+sOvsA1tg5eZS916X/2YzG27AQG+pDPWclEtTTpJX/0v
v4PtBZ6PgrBtFd+5fiOSjiYHjjpkdZhHjMRfcUpjaIk4MdLv3BXtIdVSprdthMaZ
X4Syvi9O6a+7KX2zBUxvnrtMFhxKfX/ENr+CuDHyE6pIv6tsKCiiSdUqv0eihSGU
yE09nmp5zq0KJjJk7vicrV6VMjhJ4SnJ0Md4qtBc5aGbX/Z61FcEGdumUSmJgW0K
cU3mMgUFbaabHtj691sLzshym5n2khsNqbkyF3rvBtg0bW6Cw41vCq4P2Uc7NMA6
7B3DZ+FLFTPTAo81A/Z6ZBdvHp6d7hrRRF0hRHKLGdDBOX1h4lEvK/3oLoGkuz9x
VLw1xY34mndNtuhPNKadM0XupFbSZMNUbCu6HhL6Nbw1A1lVYKUVM8SbDWj4Dg7C
IF/P1jOcU05M0e3GQ4ikpwF2htQHvvrGASM28FQQS4M2YIdOlUQKX00+lSPeustC
B6l/t1UbPZzw6DL8JuZH4kwB13WGspfbiZusNE22lds6oYP1MQ+angstAWCa4AuL
rPqYkccl2Y0+9M4NCjED+gCn0WO9wWE0J6iO1B4jBnXPXdQNyv0MGK77MO8gF7r9
N9/YUPt2Ymy9hJZCVDUTz3MZnkz+fs6tdExojgL1WPrFnGxiibagM08+DIfKHEkZ
C9VZW5rMUzI07goXoN6kdmWLR5DdUA3s0bIRkwDRgks+zmXlpNs1yQbbQBY5uuJm
BbhV+ReRyLhb4b0M31VsEvvB8fZ9FKXq1j2Hb1bpEt/E8xls+qjk64C0kOm9ZiK5
yKkG7HHfl3i53x1kOeASFyAwY/+qXKGfN5suss5ydr/EWIf1v9klUahYHMLPCREj
Zj6Ovo3URzIwSA9WhuRH9yvyVRByILw0jG4N1xYsZqgoGyQzWXNRE63G4j6op8/E
Ej/iS3SolqUTszG2Z4UcFBbeYCzmhjkfyhKxbujGlD51e9I+KVBc1Yw+a2pgiSE0
16Dx/BaQpODovNMFLWERTzWeFVHkYrHsgGhlC5qFth9PVQfc5MkQWWw4LEFvuLCa
xc7Ytby0LFmQnaorVbwe7ZOYI6b0BeCpV/uQ6+B4WtQEaxPQl+xz/SU1lINw1eCn
rwUIaek4ofLgXM+ONlK0K0dPgj+SCEpUbcmdthMsG86xwxZxa51nQ/UPIlmxpsPg
6S8sis5HJPhezgURp4CZn1iKoiWbu8rEW0jb2KbkJ36lcc9ysvuhfGvuYOWwx/sH
PUrQW3qDtZIBfZzcfwf4yAgOTQAZSLSvhvB6w8f2yg52muLtlw1WoN6gTCibzb4Z
yF+4EBznG9mgaVJ80m7Stxy+gXCM5J+NkyLKmOdTvgAlLUt0KPMXhUgcfPvee8Vf
Fp0e5GVIoi6e9i0UcnkqV3WnI7x0DVmAAoWOs9Sg59tjYwaAkKQPEcVLS53rlh6G
Km4mpAqn/4QUGZgu/SI7akYx4Lrrdn47sMjZmIKgz951LQy3kxQBUKHhG9Bsd/1j
O/0CihkztF0h1DwKpjgGxXx/ECwkLgyyOBOKZ1O1yIZjQbfDRhN4U2GxHZ84gfWP
GEjMTO6NF8V7xDXMDr22Og+/CsQIN7f2XOijA6GMJiDZNgLvmTYfMx74MINbYMX0
A6sNsc4pSwxS7B5r4u+hRkEd/iHppZmoq40l/xyVW8ftyUnqG0FnM9373/sx1Fnl
+y6W35EiaHCkH1zMpQBZ0QQZXI/1B2M6E+QBtDioTcePZu0pcvLc3qIyt4yXCvT9
/MgEsGYV4jOSpqbzTswsldtj3rnywoz9vZKGQbDimLoMRVJJ0WNbrlaHt7E/qFCi
FkxxYiz4EekeE7YFi4pUIbBmGGrnBLEuvswjd6KSJ/i3h7PZAvudxrx8GTmCB3IY
MjEgeStE4utEbzugglYgr3ZkcYuwENwtYeFkhC74N7/KCcdsHsGGz0welAA2Mj5s
pk3xvWHzjCDr2W7sNyLVJMGAUI45rtnW0Ott6qZWgxeEVlWZEfwf5bbMZDBAum/V
eIEiX/HSsDIvPWs+J00VL3RtEt3hCiD5uJB3rKqMnFobil062M3iCR1sPJQvaZN+
qNc48A6ZoXP2tHanxylU62BSSIKDRGGaf15n/Lbkqz8nuZUgfdYw31kgUpRfJgxk
3rYkjFRWYGf7Hhiy9a//IbnQZlHGNzwBOGijjVecoWr0+kb5zgeLsI6UAla6OxG5
yFBNlWSZmznPMyS/SayZvwDTfkzeDr+tHr9KKn/Cdso+K9DSdymfEHTdEVa4yTQH
5iQPySTES919uW82++LL6eNNcXv5W9KR9vtUjmUhQvP49pS4cxK0tpjRs1U/pY7z
OPCpXDVUHUDWIyWKw/LNG8NzRJrWtG/I4ueoK7TFPQn2oaiXkzMwwedqATSxPd0E
NnofB8T7uiPV+jzwDZMIV1Mvts5zSYo7PAqIRp8MOjBS7M4Y+6D9b9lOCulss75F
kTF4xGe3udlvqshPELm7TUBSaF5LRW4Shp160KuM7ujbICctVUHTup67e27XeeGF
0xNBmrF56am6cvmzfWOqSwfLClWOGmqsZ7ohCu0w/PR1TSIoT+sPxoDRr1ucdEMH
Q0B+5xERtjhWKaQPQYpvI7oyOIAH72v6OB51Nlrk/UHROa4av0BjV/M2YyAXCSp3
HTJbY9M059Xaf+OaIasMuOYO604YdS6LfgAo8nJya1Vv2xRqrm+6Rj5XbHxlVV6f
ZM1svkIRul35wVcFpvEIbQhOgeDUD3RddpdlW+wOWWN9rOtZAp7uyMROWFEDYxmG
re5+ijzgmh5cQSp+e47IGDW3OS2JIEnXucdC5FkBCb2ha323cmOWB5+upKQ07olO
Bhaa/O2ja3aLTZjS6GobihxdF9qPbttcqtqOt0q05OufqzFdOZSqvTpVAMFCRW1+
v9Tn7jF/w3WEz5YttOVuRmMPC/jgfgs5/x4FIRhdUD5uhKIzVv0+Zi8jc6LqvH1B
IsY/4UpetXAOA563Mh3eCSJwpLBm8sverBQbP70NQ8l4/lvL2wJa8jY4eKhxx3Z/
DlBW9rQ2cf9rbGmtVp43ZtqGM0gnU+qOlSw8yDjfqMsW43Ux5X+Mgq1qYL8rO5+A
OStdJ686c+fLqJ59rv5XEGiECZXNU51K0vn4G5CZSApP591JKl2lPrzo0RnPw7sl
jU2kPzKWX9WfxyRFf8YGO4MU88fCHOFzEuwdwmzFMFFed+7q2AEJSazEa132GsmM
SmGHe0aVPMdKZzbus0PyJFdF5wnb5XMHzYksMxHdI7RVoUjMSe5d4uK++YTKkX+k
YSdMnutdVZDwESy3vSjy9JJsZ+/qDpV21oIdWKNT77I2tDTHyXMN0n0mO/nndOov
MWiZTJ0jqT1x/4rcRY+duC2vk0+jtmSK2XOQklB0VYx9kHiINgzCgdvfvuBs/Y4j
WjK5X6MnZKUHSBdjyZfy31NvprWXnuJ62Kde1Ro3dajgpu8JS5sHfwh9tFarOYAn
qY57ebYtpRWieKM194F7XBIpWCwrSgZ4dfHAvy200raOI3nHb3Rt8sR0wbQH/yxN
gnPTWmxltITFdUB05tM7L9G8IvsSgYKb9mPR2nAF0ptNN4yN6oZAejFV8ESDLdMy
bM0EiJQd/2Kh9hIC4wnqACos8wKVl4YyT7gTkAzvGseIlCHh/IdTHvO6XR8IRV8L
j5KxeAzQ4fS0h1gm0tEAvNqdqv7NMIgXWyf9pQ/6jzLlGJ3ZEbZVgEVWxiVj7p6E
EIHweTb4sHHPlGTCsRUcQI+A6KuLdKunSVxoCZW55aacsIKwAjDUzCtlz51qhFKz
mAZOdlej6aSKzqbq8MYcKjgPrrZ+eqYPvAglvHNpZ+t3osvhjKb+9KUzUWrz8KfN
Lt+3RnG67VrSimBVLi5o2WcflNOPqhNIP4kbAgtxYG8Bsn0EVEFcuzHJ7Wi/z8Yn
mibbuYOtfRD8KCX90wWHWE4ag+m/SNlx2srntroTLwxgLaLsV+BUz4U/uh596IIb
lVQgbU23mcYg6lHYRnl1vFJq85KxPM2aCRWIAAzzMdCHydoFeP/5FZM9KRoNPDLk
oV9Q8r3RJ3xEwzfKR7wq5jvR67Uaq7eMVFfNK4FDN6qAj7vMCHLiA41ppLwtC/df
5Qgcbao6wzCZnL46wNk8bjYbZ3xQW+vqgRHil+EO35hfLXG8AfMCnK1db8ttKSnV
GhVrx3LQ/GYuxAuz3enoql7edVXmtZ9D1QAx1PCFMJ11pRzQy5B1b2iSz1R51wtg
YqdRl27z2iPsxaqzfVoZ0K1//nAP8QsncPAK4SfBg5TmeDNXN6/fgQUY/ZqjpUW2
lGdu+dzpXmzneuslrVU3EotklB9cjA97nQFFwtQbgTzejtH+1Q8T+3d0wQMYzh/E
bBv022DPUnR1tj4e41Aq/EeMUjvBMFHliAZy8HRnD0IubzyOv1pPkjfW1GbQxKij
fMjOtKf0Km9ycWYivuUrpfDUrvFXAcbErV5Py0DZHe/cpIg4aNeCCmueAE1ehyto
KGFLPpdcTzyWtCt3EGxOerJFmaFXe6QeIbi/22i0tBfIdQak0wHTJ8dQUhNf/jGb
ypo0nJf215STuINLWr9Rhk/gMFNY/3Kd6HUyDoI8yg3mlQo9o27IliycpPBAKU4R
LxiuWyM1eOGRm6NHXvrmqzst4VNF4g5NrdyUAieBYxnlNIzlTiOWBOZ2B2v4VcVH
T1HLKZqWcpaJSv5HIqeRGcgQftvSecWwqFxKOU3os6ApWhA/apRx5kQAF4H3Wav2
CyiPlAq+cPJ7hO+XtjxnG3jj9hIPEJckeu/1heu6edinFMo0zyUXxXhhr5tyE4nX
CfeiwHILoqIF+ePJsmGE9DhGM52ZBNQHss2K+sB1qwGa+gpcWNYUnob2SN6hr3VN
nbtRG6GBZkQVG8IeUgnFV/GvkUBpwz2939yfjjiV1nwY0DiQ0B6mLPZBg2JWQkCd
Iu0SkckNi84V58IA70jFiPPG0XEEaULyw/7OiVek9QWl3D7K2H0A2Zc5BmhcWWtP
pf3cPIcjOefClcSue9ePEeaOno9bqdq5kNT5BBxsW80gwgHgK1JA5FmGhmArodBb
geEOOl/5zDz030/UN1gFiSVr9Leo4+ddTN27DvJCEC9AB2dqsHLpGL1vglvzyZO2
1agcocHpPE8KQXapl93Bu8dsXDTFzNxOHwXCgnDGNiOpLklTbb8iLLAw38fZSUc/
n0rWSPlICK8+ynMc8HBKnFr3PEpDQbFCXUPlYL/T6PlJKXZ43jTcwCU4yitkY1Qe
0k9ZzjIT769lGDpP1WjaETz/ETtaL5JdcdlBcMelRMjjQp6S3io9gJ0sQmAyKpBN
gbeRU48h6jgRWuUrBKioIOXgWA+IDklHhKszuPLrwJ45aRTVcUMgOS2aXUcRqpjB
1xG0LMCwxrFd80ff+koa02Y6rnv3DP7VT9qVeXWqyRxCIdK0NFYwW86g+vErkBva
2pLV8XUUV9WVNZPH6xPN0/v1B33XeSCYPSfNBz5Ei0kwvbHZO5z1YsiAy8S+qinW
Db2c+gLygxtEdMCWbL2usw4x/vqEqX2MHbI7O2bVO4S0bAUUU+9Jt9lfc94YwSde
1vgRAN5v1Yv5i3OtqWQS4QwMq5xJrbZ8QkV8SKl40IITyHKOQFcfRjk9+2pXctFP
rqt0/ZVkMpCxoSjGGXmrKuAyu+WxubNEnG6uKxRF2yfeTLNvspG7JeQ/2EwZU2vZ
Jb2fMbI7iCFBeIFPu62bBdw3kOf1Da6gKUwy0pOgDXDG5m2P46Fr5uq4apbQ5rLK
k3fPpXY1pkyqMk2xlPwqIF6zABe7TWcS/fPAEYnDT7EseRlPj8Ka80N+zjKqzai6
VIus9wjFF19rzOVv2GcWyj6pN6am61sLQfhRrrpaAQLIGPdmBAn22wK2L2pnrrMs
fxqc3HNuhA+F1eS2vSXK4WA5C/fqzm23D2ELSO0t2sjqDbTunEhey7HiBs07XNCX
1V6QITD3huCquomWtAIoZ8uK9l4kJu/ACIrFWAIzetVl7M8z0GeUHQuhXrDdubmg
79YXwKFLFluM6LSVFGsg0tW9Oq0UgtH+RQhUenwIUtrPU0CO4LhHgoiA+Ho9dupI
GKtYYhTjn9vOJ3l++IQTGSu5vvazhUJoHfYnysXab/ZTnMtuP1kPOo1kjeN0msSk
0o5jEaZ/oCHkhe3CFDChGo+bCCj9KXhSiwe3+7vEbI0iaX5z0rpNvDMQzBg5JlZU
r43LUZd36BhC0iMNCm86fn4Y28DSIMRZseEguEvQVVX0x3RgbbWWOat+CZTiN7SL
GG08THhpVVi7CalrfgvwaL8ZBSFLTZZZUuqDz/YG2amn+ASBBT94stUfkjjdrHZZ
UfR62xSavZe9I8mPpHJZrXoMnpwpfGh+Nfu4dOAPaYTcqTSW0ZJEvEryE18tY11/
KW9mLDyPMb4XrJBWCY1qINLQYlG/47fsdjT3axEBNrenn+J7kjVXxeK3R6M+sJZd
sTFviyo0Dgr+QtwnzKXz39W+DrC4ZXaO+BEtRByNEnl2dAd5zjDTSaufikE9511N
ceuJSakAQyKsD4jgNZajRpZfxdfd49N8JbKPgokm6NNui3TaBd7BDyY6SuMeok6G
6CsS3nvLY1sRxMv9r/uQ/UEOair2ldFHxKibByTKc/mFDYom9x7ghoNTAIuZCDfl
WGwgpIcb/5QSL+p+aB6mDySEaaLJC8bUDB0UmwN89SzDECw2VkZcuaoT6/Ffad6b
pQNiCPlfqJ3Ew37D9Do8Ix58nqc1y0KnwABb7xM+FJKd9C+IQ6G4DtwDx8fxoc74
V0q2wK/HJ+bc99pqW/LfX7kgqppq7x/ICFTtinytZKxRGPCqme2OGYSmH86OmvUI
rx3LgCef4xQnFUQWmBTQQf6MMnOqjeAyKT5QT0Jsb+u9pmZP6LOx6waHxV4GQECY
MBAOpIgmpiJkL0e6KUHbNiG0JEDKki7G/HRmB1w4AJxAOL/RbdoCIqmnkT5VuvWo
XQ1VK+zwjeOJEqfi8aYh7/t5itxCf7qcqKcMh+nb5NnJ02AVZzcz04jguIBSamXY
Pm8/29xzcLro+c7ChkymcUUlt0Edcu6V+3AgQwMz9cdziar72k9bLGjxuQ+UFJEG
43OaeTalqjBLXnPuf3zh9cb6c1t6nERiHwnXug9/LG/z5YjhxJAa3OI2fD7jxO2G
RkNQ56DDGNmFpwWtfb3z9gL1O80XktYUgD9UDI+zYVKDiwBIE0yZlHLPseHf36fZ
WRW6FUZouwtySoi1Vz/nyfuN15snwC7jneXWg5KxlpJP2nz4Uc6GDQd9wSj2Nh63
xURzVMEQBadRDrQhfrqaUTPxhTaW8YWVpOqDCpR14NjduA+G2xTV8WXJf8yInKfS
3eCCf/KqymBW8odf/Uk3665r/eupTRvMlOlXAXVh5ELlVWzltrbMyj3UgYKOye/F
huneCEMqOL7l/TIMCI2tnog2PE1E7J81kNjkVKQVzoEBRHb08ZN59YP4sW9g+pfV
yxKLmX43ttczuWfPTw/5buU9ALfOwiYB35Ammdy/p4dqhsUaFU4GqBfS/R6ynxdE
UnLijQWHCBBEgYVfoBEhBHnseCaN5JehU+VQL8V1esAeBMMPLiCd/lGqc8NWIUew
GQQM4rMcp845mQc1kU6FKasWdU8xYTJhn1ZWDVks0+UBcAJl0g2+jOmB/r/Xtdy1
x5ObNlNVtVc1PvhO4BprGfFG5M+f7HglPrZxS7mz5wL/0soCh3+WyPtoLWhm97NB
0yjZNjtp9IOrKsPd9PQ1lcAAjCy+h2JJdpn27v5l80cIzSSwgO3/99mDxLkDIkrE
qpsbqybk7rqN8X0RPym9ln+tcsHiX2ICt/dl/Tt77D7inlDrvLBG2/pEjdU6w22W
4hZzCYA0EvLV0v+zH+eXw3gmTCTiF7asNZN+n5rVzekr1bZ4X8cpiZlm/9jIlI9Y
0GvpheLtZ8yYC9MXmcqcvqVMiuc6wh444EoIjLmxuYSQAw3ygbb2LRzaynS+3cE7
mULfN+rNnP/Q1VU8K5odq7TVep8sIXeTS5lzKiZcPToW5sCPOVMQ1urQA/J/rXmw
gfWDg5I5ThY0yTtcll1r2/2SeDObsvqze2dGRvrIm/lV7gxcozQv2t3/sEHlOvbu
vsVtQXHZynZ5kYRKbRSw4/WlKZxXfYje2y3TjM4NCFgnjoYMwZJNlhZa5uQl3DF+
ems96wgVdIpbyqouEuIzgO6R8Y+Lp3skcsjp2ANaeEEdUE91uuq0/JPutYiYCli5
v8uCK2njg03meCMSnN0/+sqg3Mz0y8gUsw8etvZQgdVM/LZptr5Qye7/r7Lw5ssE
t4nu80H3SQ1q2oR/Or5QJWCK9Qj7wk46oaYiznVLW+jJ0xLvKMMkPgovq/q7TYDJ
Ltr1CoUJoU3WzrTDNSmEQb+QS729fFc5nglHn/o2VtAegec49JUK7WLTFdiaE1zw
A/LVVJaaPCex4jDoUUUIZCMseaopUXO5WUlxwwPwKRKoIcevGKIevcvF2ExC8Lc+
3KyPF9XG7OR23kgwkdjdOJlsa5PBvjxeKQ7K0fJ29D1YI1A4l/FRcbbgFhmxs4sR
047W2jjbiMKWAfjW/H2v5HbiHXTA7HwC2XftDmeUdlVTWvvLJmsFdS2TFXOKYe5m
jVBSZxpybbAfol5sJJx+Q/znpFhTrG7Q71BzCU+3eSEkYXbcAj48kr3lAMijVGb/
SEKraygCq0/Ut5SuewU+V4hZxlOFRwljyD+XSqvX517DnDajVZNCRE5tHY1AdwOX
S1YCT9TK63pb7LoWbD5hjXjSsUFKtN0qeosy38F++RT5MVimBnqwGyDiirMG0sZU
bRVMYAs+3GzkGdDg6lOI6v5Ra61fB0O5hi0j928a4uF/9liBRImV9I+LWHKsrXzu
AuRUlgdPaqrYtO8meOIAutTo2cKaJCJ9tWts97yKp0Pfu2mS41rwF5yNHX+hWzCQ
4IVREB6dtA7qWlBAzxFg5LlUbILV2JqIep57SQiCzbfFDG0kPSlULngTU8okIihR
ID6AqF9z5xkw0iIsnnreSFUoq8FNCYrXHDmqdh24YcyaPp34BkdCdPnSPaHjibON
EPR52XwVyubRs5InAY955mCLw5R7HgCyuCov+9ksVt1Eq6m6OEA79L6uKQe0Hg9M
kCl92IefYC8u9QzDurjGX3nbhZ7SwbJc06VlrcxEOqDVZu7eZ84aBOG1cE6f1h7h
Nwu1/f3ZcUN/M9nToYCRGNwggnCFGVHOnSy2vNd8gcLocePKB9P3Z76ghSUhbfmW
+oc82TiwdKK4jq1mm6jPInopdCsEmiW7ZPxxAdSuijh4ox6oy3gxY/ur4NHLrZxu
QyFXoTIQiGccPXQSWprambDRF3mQYfU1ifIyXTGv/3LXSD0sca1kmnbHArZmVfSF
D+4P8bj07FZQV5ajsCrx05wPo+Usxftnu5EpSf7GnYGlvrcwTbs3dpE7zPOGlbGq
t8vhO1Z78uuYx74Edgatb8WbwWBOgQKlNFgfEg38SpoDT5Z/ubInrv8f2JTtaEDE
NtWVu9je8G2HNguDbeEVbLe6hBHpdLpkPvkfVliVyOYPVDqTwl/hyNfD0KHa2UCj
m5M14lYq9abkgkqVBFeqnzq/hFjUeocdfcOh+OQxNcAXIOhSHUkdIvRmc8oxIvZj
aM2BuuUgafMfuZMz2mB7tf+BWnLGnhqpCfNSW88nFDdsAx96/IDujHyVplB1fAWM
DNg+rXI4wkzcQk10N1Mm0h5x0MnBf4kzwev1ojaqxIM1J7vt9fpOUo2wokYpLp8a
PFIuP5mgR2kJe7OtrPZlbbH3vxXUmZMxzImLi3yRX4NfnWx9KZjZabCiRgp+9wKS
hiEddvnJU4IxkmKkuENe8fBr5BBwNgoTQBC2ywbNbcTbrh8cXvkqIjPmJNye/b34
T1rkXZvQ2nXEc9Ne9hYdkEMTELL/AfqMpW0Zudu/TWes7hTfPt7LAS3IX+q/KUq7
UYYAtjusJEo4iaoAQwZq7o/NnFL9tIhY4fnEentiguR3no8HdtBHR0b5jfJlWNH1
m1X+BfP0irW5mIOG4UbURIV9HRuJhKJjgjQlBKoi1zdkO3/EkvSM+kDQi0P3t6oI
pm8W820LFvJbOPkzesdBSIAxER/KUgVc0ON0bVIyYBn6jLk6OBuX/EVe5f7zmD9G
ezqMJDG1Mf5IA5uyV6WB/TV+zW/j2czO3MjHRgwtSKwP7YDrvUSwN3cSjh83hi8n
WZSHuTva8Bm95UCix0e2TAO/oQVEcCTWR4CA2QZo/q4PSI1ILHVUMiiG7htY1emY
Ru0/Igtnd6G4m4Drgqc7tC4jOki9oDpOhKiWzDIcLrB/XjTciESy9T4ElOSKLZLw
GVY/K/mfCvmzAGozWrCtRhI92mGIAAA9jJhgV6ypuo9HLfNuj5elqgMHXg8/w2QE
Vc2oahIUt4O/zLj/LfLCr2v6K9I77Ta1vQTOmv3M6mIjaxqTBdJ2BffgFdqXj92W
Ip1dFHJotdUREMv8FEhp5zvnszwpyW0X+Sac/CFJnrTG3EsHCOKpUao1BLK2pAaA
MPbmzHyI0RoKsJNmm0hml/KjMbKRYyebtvRydEngIj0xjPBKUd8YS0QHSjy1cEZb
7ZD/4ZA9YmAvBb+W+68oQWifQsK6CrzTwLS2p59+ogko+R1rHgiZTQeJfMFEEnF9
bcbeArPMvwiSMReZJc5wWv7lx+2SscfVEEn0ZOzNyAO50YJ/cISiWOu8NRaYcqpi
KVJMJkX07J6bEH5ajdZw+kQZQg1Cf6yARGA6eXyiQLJ7Er47A88N26wogTYsVTWs
YdtU/vxgEMCNeUluczvtZAQtYgGn/1feP+3QjtN7i5Sk1NzpEOs++JWjCLq55fPz
yhhFctnQdqMOsWpJ4Y7XMq3mTb3SlqqQ9Z9XWrpvkzno6oT0hyIbhsBoVDWHP/V1
91lWEfh/wyQmj9I3VIQJYJNAo8Ibp17f2FG7Pgw19fVyVNEROvSEIqjWeMZ0f9gb
LdqFmk2q71CDXA6IV461/YrxXkCopTKETKau/U8Tt77WkI8nd6FlwCrnvDSPUKkW
TWhAY42TK+4icEc7KK6+LS3HUXSFvoZI8Qcm63FWr4gdYDALrxzvd6wxYZPhk2XX
UHae56b6hiwGj2ZMomSW4VPZDSHr9XtANXpKlrQBSe+o1MCKWoQMHfmanOifNxr6
/NIXq38PcBHZMQc50qVvHRx6eNwb149sidlMA2K0f0hgO/lsc7IWP3WviiIA5LeK
58K4ABqYXgOPYccWFAiWCBgpzZY+Utoeo5yT6prc+B55Ntd1Vmt0Vm/XtU8o8tdJ
UaOI7ZlSvMT9SGhzDIOEXZhrneJhrWO4FXIwuLJdVPWafBYx6TJPIdxq6JX4GPcB
unW5qs2b6mGSqiGMR0RP8DYICosYIM7w61KNfNu+IeATem/K5WwYyz6i4WEVwHvF
2dTHwkQ6uXzhUEBHmSM9famIOR1LEMCWjLpmvSewyvFrhKNpDUDCcxqjo0dJTsiX
HoUSMrzM15W/PQkIRv4bHdK8aAMDdBHaoC9gnbjXKOZ9iu3bXPRtdg31AlTZCEbZ
gKgYHFmbQ883D0Qgd3jhqU0okEwc23Ybehck0jX0wllLRn5BXv6D/kVaVeDE8vpZ
r1taSyfinegV5K7rMRiew87e9p6j6FIkRIUV5MhnYaMUmyAsCNGp/8T1L7uoh0fR
XoQhotQlUpHrFhbM+lO8D1tyfNvdib3JKRwrpob4Da/55b2uyah2Q8b7hMWFmx36
Lo8KaSV3E9GKG2kj5lYTOwJoKHT4TOHC8bdi3ImkkjLeMFgcs8B0AP1HAq7e1ZRE
d4wLHFfj8lLDuTR24S+VGhScFwBarQw7naWV3hNizOMCUAHCxlOk6Pat8WlR49Ev
AMa6z3YCAYLuqaFf5tyIoVH+dpa/B++Fxp47FCs9+8umXif05G9yjBt6+G7qUaAY
hYXHKkjlyHJqCCVSTC1yFP4fSzpJTc9tE74QCiXVN2BHqPqNbbYE3gRkjuJal97D
uCmSLaskIA09RV9Q1YcSmVyGMxMeY4Ov6NS8mr4c7zfBSgvKaOSCqSdBnpuUGDm7
ElSO35thzBHn6Q7VHYncyxLjdKXjxfbpHmwYOknnrude8GWjT070wfY3LsJFO2Gi
QNCNix8dKAWfx9UxK9B1My7DzFm89NbNOOQ1jm42xkBtko9eduNULPNGzZTqgA76
M6ui85c1vqx9MBcLew2eKWwSihaF5kjdxjs3nfW4PCVYCLpDeAum5WTFhswWGz2z
LP+xz2kaf9WTcN5Qwt1ht1Oc9f9G9iEVPBLb1/z5K9W3mpJpmQUSfcjyKp3j+zxc
Zyh3q69dnAlhXmuusUIFFLtOtGgwP3pPW9hA/0hIviktik2JNdPdibU7cTqgXXE3
AHv/dEb03IuAKNtfv9q/7QagNg5T7fJlvjb8afaIZH9WDgbs+BnbikOPBb9mmY/P
A3kNFSXWO6IPp6288t5W470unN3SJawiZRdrWL1U0h/2O4Jp5542iWmOKyklsvxZ
dA8JFkjoTk0UEuIlmZh+lws57DFQvNEhjH6etsvaGVnHW8BjhRKAVV1Fk8Nm9EtT
lKBce+4BjyO+YSQUks810sWkG+wI8KKtf17VxQJXBGGQWOXHVL1s1VjVofj+Dkiq
ORUX4gi6660MTVlmvrUB8Kh8a/041NzHkGMp8ycd+5oydXzz0GnFhplwy8V98eWq
BM/h0rZ3s2/oSnAxi+nzyQUGDDtbOBy18JKVN+X/UauWj7GEL8BPcrzxDSZuKnYU
4WZGtZLhGJJD1+jVSQcrjeFu17GAEPIiSY1zVzzrAkByWm/rxyQFf0jrBYUll/58
YxxcBhApBN4qofVLflyBV/WrZ/qNUcecB165pKfPrPOZsSXmbTVIQ46k6EsiLn2B
Knphp6mkCx+hUakQQOeAuwnRP9Gb1KpZ1CXo9rVD5m3Qj+TkVr658u36spgDZzIp
LzjMwpuhmQp5DISFWcNzN4XpKswLRzpQk+1t70Om4wRHCBHdsloSj8w5C6WqF6dC
F+W0SVNIcevmi2lEX6dqiCfSYR8Lxh0/da2G5bSw0iZfrLa93+fqYkFkFnSZKovs
zld76zM3caR5bQLPsU1lgJOK+X4maxf/dxP9WSP823goi2oNvgd7qDsxdXW4hrB8
X6VL/8uymzuSpYPGW+hfDNxubVzgvr7Pqf64IyAYAfSBYV1K+pFnzPjN5WMNgZfk
1P4wHNjKlnfZo1FMry9AYp9arf90lXZ6MOlzN3O4pPyFal3EPCr+hpgET4Gw9L0i
AOxvSVmBCzI2q1KYPWwn3be06iXY7xiPmnVqtPsBos3VeqtGp/zw/ilTACN68iN9
qwexSfJvTZmQbUFA8pCOXetvOY3etfSPA8cpPslmkt+prTst7Eag8Zt3oYTnqRdk
dYyPv6fmEPMoCAfChAh+InV5PzRTxDfXxPu07TTLjXaWfBqMV8Oi5CDnFhBkecA5
9/0UteyBccNRoK5uWOvu8OIiGv6Wuzfu/abKYcDkE9Ee9O6iW4K9DT2nHdSqF7e8
dZIdjLLOlaZ3x93ob2rikGOEhwdpkepXKKUcbUmCPCfhFWck7JGKGkQqrhqQOLir
Xdjey5nv0E5HzuFuSv3EA7dtsEeipPoiL8A87RcN0XjMsN26d0I4JqTndBamewGh
omBSZe+I2O4izMQtmjgR9TThmDYeLVFhRuj7FN5I1s/7cEvh5FvX1D1N/928ZRrq
o435OaZxAvUocEk94MsaKXCIp1wLC5VRAdz4l0SmSO6F+m91zXZVOOuIkLF0aWN1
+rHdzrllhKT/mLeLZXbtpyvEh4kvnr2GE+xcYg/NHjqiJzjGEvazpGtTHy1ZtI7u
nU7MZ/4WfbMrDBykAli372ib4znFw/rPO+j/gKDTeHIZzFXxBG4tLLWam0JDD9MM
HKMA47BXvc6AGlLvH4286+V6HiCA8Cz4ZwbzHglHQO1jCHAbPYzWqoNQpoezf3aq
Cp6KkFdSSZZ87mglz43tyVynxvK911wqL0nLH1bpRvhR8HiutRRXovL4PvhOoU8e
PbBxD79iUmN3lJHYQz7Kcdsq9CpHwQ1BxcGJp1j2+JbXoiiks2XBd83eIyryG87q
EpsnNaU10eeVI8hkhzxayxzU6wTsRCoVmKNt5wmQUfTL0uZFiwv0IJntKVjywWaM
vrlV7+WONogWI9NyFvQS+KG70xqNKF0NSmCiLup4nF2IA5ol7GzwZfs6NogyOKtQ
hqoJECSLmpHZ+hb2NimuflWCTWonjleltYkR4w9mOU7x0/Wz98cloDq27MPGUdPo
AmgpSy8ludDIJxavRUarb3Iz4Q1Fdf6cZ5QMeF2U6XEs5i1y4bN0QlHtlONA0eE0
8jZgAvAr+VjyxlUHSYDgDnBbte262tSLpo4rv02YsU19Gr6E012LmfdHWgD5Eg93
yxgyASl+ztM+Gj9v8Psndhl9ApwsEDC2nrxI/FQ7nzeqbSHLFY8n7emp9YTeZN/i
fbq0s6WNxdTuoavKsuumVVSzqMbQ9RysRU41bQocNHGc6scX/jtQICsVdxkT+g55
iViavjSi+PbTqb8nAvzOHHJyqXL3NmgG+aAqw8kI+Uu2fQJJ7SDgU/XsGxZaLk6m
Bfylh3d5mrt3O1EIoWfd9WRsUGdRH2nF0AErt9VZDNM15TaxEr+1gHH7S4c9yX0B
5I/WQODBwanRjaOmCkZJLBFZyEbQ3ySUqEsAigdckSK5nYMzF+n/A2wp2qfYgRB+
VAA+LkBpD0x7fN0vOg+WfBYmZZc+TCHjDdJbjbI+wKf6Z3liryy6eGfBUwHjok5j
EaYKmsU7ycoxCOn0QHJXU5wGmRtUC9WoDfWUOP8ALUns2Lw9q2qHRBG3YH4YNIe7
W6qXVWnfFmp355IwXIrwebbY4KFWBEykG0jH0+4q7irt/kZzJbcIsCzm+QdMq1ED
YoZTb4kxVip5VFt2lShEp6kC+jpMpxmeC6f7KBg98wbsLyLHlF18qfMae2Givyeu
aQ/+IY1txCrKGBXdi6OSHT259wLGYyZ1+E1YOhvanKCN5e2nQxgrh4FSpAn8jA1U
h7af7hXVcdmyuzAYVbflPLqdHszfcBDlOzImvPCgjrmSuaXW8QrcsLYbNyuel2Ep
gZvzHNqHP1oIQHB997vKb5yaszWYi2PuSO1MJPlQ9a3S8cVfJyRadiknANI8zMRi
s5O5ICKlK1iKJWFKi2nMJ5OspSjoRbnxUSweiHJiOaLQeYxtZZA1lB2JBxosrsm3
BpCLReaobUec+3jITFxf9b67D28wiocI9P0RfuDQGgpINWmaO4nk44LznjLGdsEq
zNN/rfgjVu/ClVKoa7FhrXC3ZCdspeGVv436siXYgYWsfqGPdjVxzeh8Ce5IwF6s
BW0CqJDa7sNTvrloCw5Jf+GYNjs1oO67J8m1uzsH+zhjx6jKEiJS2ZzavuNnCi+E
zk1ZIasw0Wi+wby9QWoBBC2qEttk0ZQkJSWfFGtLCL75m1frJKlQI8xO1QtYgYyF
uipimhGl3wETamfp3e71Y4ekPXQPtc6zLvi4hg+kFv/pJrVVi4Sy/GGPtMvMgOEG
9vEPeFfITyIL5kDd4BQEblDiSTSj2XJzHev90P3VoajG/DzQDjteC6WShHhITrhc
eQox9IUnG/MLzhbjX9MHbK3mv7/THWDxgA2vFdo54KbukiedS/WJhrNuWTA8ueBf
ndkSwac1Sx8eflqFDHF/9iIerPI/jA1Gno0C2ltvhBdSSgwwq2tnK7t9P5vM0c1S
jQxQm4chVw+nscSFA2AF7M0IHokrvxXp1uxm8Lrg3fZBKvLejbMoPWEoqt/KPRL6
SU/HcBBP57S2sw/R/3zrGbRefYF9wCspUOI7FqZfK3wVHzAGQ4f3zbSBp9yjurzL
R8bUXDxQubFpaF0aqh5GrbfzKmqAA7wHFtbeM+TBIYd2JpVO5TVVugA99k/Agv5s
fnoYNuXxGKJLd5pVRw1ZweaCLLTqON2AUWlckjWh004/jNUZoQao/lT3VrNGg64U
mZ9MPQ2WP+wqiKRccKaDTOqpGmp8JW5wlNFWh31rGxKVt/EvEOV6TRFV+6xVTngN
mOSszgC2r2U0dlw6Kw6ombtLypmnbeQoyxGZHkXVS68C6cmg8E2UJKJYMDtz/b0Q
Leld+kMJfbA2Th4PteqpMVtFJhUhUSbS6QrHTTh2cveyYfklDzg+o6TSK01nSn8v
P5ZPwwTh+DA5q5mP/vtlm1R7jAtLYsUrdG2EfbVd580UGw0WiSZraCKIT05Rrckd
s+6wi+dD67kjAGb80gfKo5H4Ki8xFt3zOowHZGo6PfWzLc5Wl+ZXDVpQizPhvuv6
mxBM6hX3VkRTLJPOIkF2MO/EgOXrTiXC6gnqYQtg1oeeHH5t4lShvqeOg32ccKDb
7+So+f8ebCgkeK6wQm3fZeKeYyUAq5BRwcFvCavVya1O6CUltjVIz5qLl+Yl+sW/
StrazyJVBx8Rjy+GGVhtc3iMoC1faOD7dfEOubjYxFCjXFv2cRNiqu4fA2klS4lT
/83qZW7a8prc3nVig9ji9m4D/Aky10fkCmSKH8/2Wsu2lZcmH0DRXnKsqmvCe5MX
FQvbNi8D8tVZ+GuRn/zOGGyMl9xs+pJJgYRDXqJOrX8a6N+dO1+ZyvN5ZgJftu70
fars2XJ0sil0JccHUEE214LYISGHY5Ex7ZJUw1BrKx5V6JXxRqICYQPckpGSJgkS
NvyOsmAs5MUOtWidbWtQTrLTEzrx4pupILxaE6VuT31FFEKqBPOvjlbOuU8VxOu7
Nk81985q5Lv5ZUXjVsOoDJxZsm6OA6ymMpvMECLosKk8wiNnaJY2d2QNn4FX0fmz
yh0WYW2bSN6zRH5+aEBPau8Kdsp+nWesJlkPZXM0DU2Oewcy4AsunZAEcsKYelL0
o3F5EUCCxlZNAZTzGS1bJaVfqYG6jYPa5B1qHtIBeIg8CezTpGECME1u5MJYaLB8
YLEwJDW97wsaTr+vGmAin42I7t8dqdVryJ2BDEX4SloUtb52Di572RhmKBG54Enm
tiepXnHTzr4InyuTidAAH3oNxP9hugC9Vey1AY8g7SDUdlR5IqBQaZruZGZw6CiE
aSB9Hed9doTeC8cSr0e+zBH63rxva21xLiT8/cLw84kN1XYGW/fguzJgEJKMcMQE
UHz2U5vdsEOmA1anfyx9GWOp3S+ZtuuCRN6zMnMOmVzGp4zK7x3L9CRuNxUEM4Om
KSm9AO9JrJn7Ok/Q3uxlBZ4ySjuPHznyWG4MxliGPZrwpTfxURgQL+PYYO0fKvCt
j/5FaGal1HDN+4pyZ8+Yl+qavTa4BP6ZK9G7rT2a8rPbWcms92SJpI8igl5beKLi
rsRuv1jab3l7jX2zwbygyMmzKCVwGAb4RLxh2inbhG7QpDpfZ7tXuXJpgDQg9xSF
mwDdHHECJ7kXTT2UdP3GbxjxbPdvvRscV7DniUlNAT9kJ7IQE3alBJEkq+e0MDpW
1GTNnvrU/neo7rTNUGwLv5O9udDuN/+CbZR/czU5EMkdO+UFyUQkr8DtO9jDaKV6
I5J4EZ38ca8Sjvd4sk/Y+wE6/XUCLovGCQDcQrc/Ri5GB2aiDpJNQCH17X6T1023
+MUGefi9fffwNfaH6jG+lQluGiFZehBOENzmEvFz8ii2vVfwKBbghUHTJubxcnMU
hI4VDEbcmbQq3NI3WGVPJpHEMZU4mif+jO9R4QmX3xBI3vsp5/g9bK2pyjEVYzw2
8eF3wEvZwVe7LvgphfYuB145O6qsD9WAQ5bkrSK511BTmy8kOqa9Bfxjzxwq/z7A
LjwIKLy8KgnXqL/pAtbNfo6Eiuw8Gn4KRyALaSEMVXmwsUfaVKSoW6bjHO27EJar
aB8RPLcaALNO0b+FVAf6hu3SGzUsqeAGKhQyxfQcbp3jo8l67/pwQDnIbVpFvLB5
bTKy80fYNM4D1PlqZnu57UtK6WfrF31BkT3uwjkoK7vmjagYgRwpm+4AXkWNeSEg
+lpVpbLKO4BCLl1DAIC16INoQLrdixXIrzErNVqTeQ480y8JbQhyRDptGb3a1t5l
jNhw7g+osLsGWDhA8AB2iBbDbyHVMMtPGCeLj1L9NNwqZqUV9KD9AGXCjYqrduB8
cKDVDQJcr+RG8ZLCrbc6ESOe6ouDKIrN9kqtLgppY7I89gKvL/hdzmd7r4Yh7KSY
cyh38htdCuwtDGZhZ0QZX4UzWQkFnmDmMoj4bMDAMzPCFaQoWvZUkSpWJAn47kMk
YNTUvZch2fpssviSEeU1fhqtp+m17aghAzk4DigNpJ8B67zb5kBmkEk5UFX6JiEU
QRX1KSMhyJeGdA12FupXYt3pD7q7C/4q11+9zjRmZgkI0trDLaQNHKvIb0Ieq3F3
TvZiFp5u5XUJED9PE1iuqt9pjzNMyALogyiGHrMFpl8E80tWgwdpTSS6kh1Zmro5
MJzM/AatP8ZeKNa758Ud2wLFLPZWN5hzqqaDrbqk2/+F0s4W+71gmN7COBonUJnt
k4FK/0gSQIJiU8qHmL2bO9cVeipGPzPr+8UQBkbgofw1fbGxjdftZt6s+LbGpsnJ
iXwAeu0PGBgIpLifsWxhJ2GMlsSMc8SmQRsG5C+TMa2aEkKl3CWCOFubwT+PZV3U
nVWXnVmUmvveao1wGREXDYm2JX6FgI2jQc+2XM72/4W9YBp108QOH0yexB2ErXuS
oZWyF8dqTfMvcfE4dMi1A9Ugrmc158pI2RZUGeXrbV7f2Q8sthvFOKTak3zA3m/h
bXbCp8mjIDUtw8mmQ6g/8GxjYCUvxHH4KD+0fMYbrE+F0iDeuiF0DIiHhQooZQ27
tJsR2xGnWvcLa3mlqZlB1ZSDgGJ8ukB1XNHUyPoUz7/1R18hwlsAXYGzoiiQCPry
Ltn+F9j88tiB3AollUJQ4bHm1szzF146DD7aH64S1JiYTtLjmq4V24iHnDnYrjpl
Gi93qNlI3ZFvJ952VdIcHFrutZhs7wyYtAKMAVyciUeKtUqSNVwUxyp9m/DlGZ+f
NHWRRm70ujEVB07YPiSaxm9qb8u2863RE0sfhsnFJsK2cZPAw/o3/BSWG2bdZE9I
LSZC4+ZNyInLNaUUE8DG9XQz/oi0VTAxxKG99UCgEXy3wH+gjHeDDJjl5soA8Oqp
9rj+8UZPn9FJRJte2LSLtlm8dCPWIFo5ypTp3achmxsAgm54MPqHtPd/1oeo8YlP
yT71rr17b09C+4/0r4kPU5mNfBnaqKDO7UGbFanVFc/egIlEcfHS4YFZU9M+5n8n
YUhT/glL2iYoUtvoOYbgy/6gyiuS8H6WHVdIMeIHxgcyMSyN8nzgoq7gztFRw6l6
jn81RZS0+BGJp4nH4RPoXfhDmohQamFhomKGIWQr4WM7BEQ1rC3PBxbyU5zPoPhn
MV7pJeLRCSjk1Sg9Ref85504qu79/eIBLPA9sJyywTc0YbrSGzV4omeCWxlxSWbr
9Nt4Og1bXjjNwhUitIVMOYWl3Lz7FmsmSEjHoA4ghGF5tJE1F9lu3X9PWJOGI+98
QCOLbYElgPzSYlLOfRz759VKxDF9TZOwai0V/jhSKcPlHtYQ0WFghFBTukur0Tue
jbau/nAYxgxUq++SpSasorgh21Ui2kAmyM7DDX0RdO0NG0wldJb2/zxMvVO+zTJ/
Y3Ra8Fu4nxZsNsRT9pRZv2rqp6+wkKMfi/Ko2rLj2xCfhMeW1LtCzcjnlrLyMa+Q
Sc/k7AEcHcouu4zXm+D2n6XTg0x19MHMwZy/qwrmfl9Ey/FJsQrPc8hL/afD3+dG
0WcvdxomtuRn5MUcr6uOGm7TPej6XgQ1pvGCOk8l7NY4jC0J3oAQt4l1Qyjy3bL8
F9MAVcu3sia/okw0zI78g41IImvLIQA064JXBqvX60qFA2v0ZurdN0t/o1cJKoW0
+qOSksbHkixy1touWVj3nG1pKbrH4NIT6DAoa9UYM67AwqoOtkYKmtOJgZvrqlEU
KPMaLr3p24tQqtmxrnSaZhDcZmcaLzKU10y1JRckp5xQjL0JlLfagGxRRO4vGhEC
pQpFgga8n5HHDc994sYbNvftJSERP2OoyPv5lx51jSoQWQKFtm9/Je2Odfk8Hy1S
a5HxqdphuvYriT6ax+F6/FxBKiYLlzXJqbDOQkS8+5UmVpVLrdHuIPy2Hj9vf3G/
6MHc5qaadydCYXx3F1E39xjv9sVxQ70y41ffWkHvBzMkCAv+TukiaOBtokMJlupq
OidEZrOu8GUPtS97fzXtI+hsohSb+ocJ7ExNFQlGn3Ph+eEEK2K622kjQomGDXy/
W7cr3uVJb2cDe2j8ctaGiAvdGEtUhCma+sW4rZUPb5WXwh0tqSXbZBqdiLfBiQHo
DSl9RC6T1chCGbcOUceuGW4/0EkHtx27IXcpRh8nQIIsz4KHyqXybZNajmwQrOTn
fJemajdYCpUGg+3pgQbdYG8RSe8EOzrVIsocD5vXqtxE/YMFLg2C2cV3DFMtw0f6
tH0AoJh8ZAUueGdeiueZszsNmM48/0SSjp+hQayXhTgXrMkMLb+U1dJ3FGRyHU5Z
wS+XO7+uZr5GHKRIKTQt3E7jAJf3onaghI50CJm1DZT+NqH8DXdMLGX0R/A8z6B7
FAdRn4tpY7sL/ahec5yPUoT/HD3dRBihJAFLkBDBLGuslnCE+QTGFL07xwdFou1g
56gO57QqaI0THOdCOGHmJqNd4m76E86WC+xxYLHvrKXu+1tvBS2CU1bH7hjSF9gs
OkEWXT74iQkmrsdKe2vr9cgw1zEaBKjaxWlwgYYx1obyEqB+3vU4mID0w+UiWBIJ
fIXV+HPrZTP94AiU5SbjVux63TH/EKwMov0OrI8lalPWQ3PVsGP+j6RLRLPX23r7
dYUGIt1T2ZLwHFJeQQfGDA5DNrPvHdJqu442Q7oPgMdGNpU6Z/qnk7ZRUO2NVrGb
BCjMYZp5QCS69Qq4wCJ3blEXjxH5mi1xBTJm8y9H1KCuC8zOTMDDuxenZUQ6EGtI
diAvVG9jgeWHv/zwwComiOMf7JfWM6DM0TAR4JNZ8CGazaTOGfIdCZ7xSu21TjCA
bsOYYvzbTTXSzp1C1tK3vFdfXbILM6B+fOXHn/2TPue6VclqbUpM1zLMKSWvV9p6
M9P2IEZFou26ufpCC55c99eLVLo3MI2levoB8VH92KU2F7UGB2TX+jRswKVd13Ow
5zN/wVE9SsQCXXqqJJuMYfotbVExuy73qUPB0/XU7SwxfLhbDgEh2jUFzzLJoCDP
JhcUsREnJtcoyIbFJM7W1JZKDwLidbsMmzuyhcMlGAekc7/gtgcaTBNWMSK1E2Mv
JKjxmVNCTj8/9ImCv4R0P+PrdKg/gtgwWuiSo+kjtlpUDUl0U8nQ7zOtcTMFt3Ui
vKuwKKIaqqvsovGoguzjT2GuF+DcBNBmCwlJvMiD6ujX8wDEBV7EoVJG8AbNO+bj
WKEGu0LB8AXmjCGanXsoUbcIhcGij8VFaoUE6ENLiLKhJcvE84lIZhGNX7Vl9gff
ppKw00FNIW9B743pJXdYzGFyElrfkE71eS8LsGVugiezS3UnDZqS1183SZuIHUlj
GkQU0npHPShHvaktSHL6vwdoM5v4eONHXR7e5yIilkkShSIskBN7jLplRvoe5+kU
MonXoJLdITRgtXYycqqUIj+UCXEBdcJz+cWlscdnFIvSJSH3MfnP1/lhfA6hA2f7
Qh7MvZn/Qq3xTJHA0z82U6G0aiad+B/8mLVyNKmsvdDJAcVlqVvZ5DmFzamMdXgi
Zs26uSpAsd9pAmlr2njTjcvnZleQoN22WXgR8FEF3SelFfC5gxi6nZIjKtYMo9G1
t3AvPXVhE0nw5wofGWiE+uErN514lcQ4bGsSl7rKFkzN0DPTKUj6VvNUYtOYGvh1
4vUJcmTvFPe9QuKKsLTu5nbxSG0XtFSvZPD0k4l1qa8QB7V5vdBrgrSNMaco349u
UefmtdIlOoQOJJdvW3KnKk+W8DiMPXMGFkHqtiAZ3OhqPo785wJXVe2SZSVA0bXv
1v8IQv0ta3g2RXNJcRgRVV5Uv9jX0N8scoyPoCmjViP8lwbmeJ9g0+vA80aV9uHK
PwlZh/rNgJAfNs+btAjUHg+QWX85ZWYlyW0D0t6aIgZXWzN0U77mBTPoOXK0WebR
2yRtDHCnVGjKk+Kry+oXU3KO+NiZwAkvEVZpWikMZPbb+dqCp3uOGjxBqfhsgGf/
KT9eIOmTSTq8ezupqzW37H85c/xKjQth5DDQZl+VyAgESRyMhhgEfcXU0xJjMIhU
U9+UJMxxHs/NHINxUWH1fFL12IFeaF15wXfcePpZy+AjFbJ0uhTk9SrgBWVbZDYk
eUmUC8RiRC1+0dhvwULaeM03dlwClJuT/xCjvDlK7VoqhC6s1Fby3+yS8+viBJPi
RmlO7Xzfb9qcD3dN+sxYjwf/6vnskRsTOpdT0kRJ+PNIHDbqus95s2xHTMb3tFAP
7XbD+MRQMu0W2HVwF0zmWlNg+5xvM91A4Ad8uXHXWbIbPQZsFtCiwPrvo4XG43Zx
Wavde8b2SZy2ak5eyOtaKwVcgP3UJf1Xa+2GifgESynHuBkHs0BSSjXGR+YrUxte
LuaS9jlyY8ZhVuuw5JHQAJ4jhLkqFT1HGE72rofc0mCDhbkcQCwIXd9xoe7Kr7lg
dBzuh5Is1j6cqPagaacdJC7N/HvmiorujF5R1pX530J4WxFaPmnhkb0D+nze8iI1
YV2rqRq14RbG7iKpKFp+S4Jv7eIal3cokwQ8L+wJelip9lIxoc9cWnX0WFiGKthV
2SSM7tjQwmMTcm5G0Quf5FJb2Y2E3gQxyQRcqyw06wmNEeptDUKidBq+H7EJ5kUF
qyMLX0jKOb08XebCNGWsMrfrQbiQ2Zo6hsC9Rg5P63iuOp9Hjjy9v4Cs6VLCA6cD
XBjOpglT0X3G1O72PNrfcqFawR3B5Fu7qD2VpjGZqzwE7OoMocoruqJxifU6zjys
XSwAGTwbplAWZ9kfBni0r3YfhXVeQhnVjXw0A5Lxiwocp3GsZYsMSI93+UEvrp/w
nIHNMwPdXcgImVp9VYbpx5hUNKC95/qVFq+ewy0mz5ICG6JN/LqzHQh558BuoJvf
oduLOAO0DzZRU1iX/rwDAKxbrzeIx+Zu/GTCmD4oGmd05HhHXX+sWCWD+sDDm/Sf
9RAMRHBURjjsfku/lMxBEP3DZtA1Jv0Xu5k03SiAy5NLpvUZO8RV8ruGpFEy8kt1
q6DQx1kK0Oef828bRq/3qVdg+s7XcROGRnpxBgFJJQlu2LiJNsGwfpmSllAUoc3d
r2C6wl6C7gdKpjHBu7nUnc7PGhTafkMJYLhGXa0Sm5eF6TZvC9VDVa0Z1Qkz3YHZ
8NB8lqr91uvag10coBZtWHFveCnS+1cU2/a8/YMKazq2y9e2wBDLsqAaJJ3dHMIS
2ZLrlrePd7i2wx/NXRSuatCSWywrF3uivSG/pfq6hbfsGcNLlf0ek1UiDfbNL4+p
lC8Ea/3FtXDC6ndQ8AzsWinjpsui4RThDIxikCrM0SNZaxYVthWrqWvO/nAZHCN7
F2YcDH7mi4vkGMyDyFINTOn/iBje2/rrQ/ZrzHL8B4wHqHcsaO2urwHIPg6pCHka
Zk9n4Wgl/00LrAVfyVR5/zyMD0/3liSXK+e9ay9BusC4WqfsBeb5atHcjx4qr1UN
svfGbK30HdirN1XI3Zv6BsLoTfM4eEjjhRheqfKnaOco/0Yu+wcJZxdgc404AiUK
khMQ5a9P4mKPKeaMdKJdZEt59ChB8v8Cfs6IJ/EgPgMDP+fA/FqWoql0hzQX/O4d
myv+ByY+puLTqGge0MiBv4df72wZgTYnxTgCpsjmo0AyE9K8i2nfqpihuIbQV/d9
MRsBhdZFnsz7xDohEFSK4/KIZgTWTw2B28eZB9p5WzettExLwZNsTo6gpClmCwRH
xnHIT3kjf1mAERtE8YAqPtUyg1Nnoft90ji+1yiGqI/nSYsq2NYyZvyoAHkUouPH
xZHbFOyqOy/nrY52Ta05Z9B1M+vbhlKj/IGg2TR08Azft19Bsp6etgVhLI47YMdF
u/x8Vu/sGfxsXwV7CswPfyhpaXWVXEA/iXrSlFpMrRnI584gEGK4ca9XOyOLHiER
4PM9mlCdjhyxerR1jMAr25injA6+DqoKF9caHwwLpo3iiEvlg7jp3F3OkYwxMh0t
y6ZBUoBgGUhXA0W9GZVqW5DDHwKhzb972w1WDKn8TVWvoEgY95A2XigmxfA6SYbH
fEqFn3HOdn+Wl/CrAd6JItF31j8eRCc32xUmexxea57gySP4jAfWbfr0pOMpIDLT
SI5LNx+KZpM1NgBne6GT7sZd5BES/DUBr62TCN0St5UpSV5w9Z1CLYrZq8/l5Rtm
NhwhNtBB+UL4pmzMmEOhIG40MhNXqToKEI9RGOgNKV9o4VdE0UxpElA1sTZwzkEW
tfW7gaVJvI1b5zGgsTu+up+reOHf8QQDDn7Ran34hNI2DiZEmpXMhevmlyaYM9pN
DpsSfrMcQzETPPT5MiMuZnTfgb01ybMCnefgTyDmLNPsXyONiSvbQVU0viJ7mvvU
kmWe2QHWd2z02+A3uxVa3nMnaYtuZ9cVjYKjR3YPArTLEstK4lrxDWmY9kkL9s9E
XCgC6VYTvG7zHewNMTnO16gdaDTWRkkQVGRcn+5nRDWQBjMlaMWdCSKtfXYUJdKv
VbWOOSJZl+jIEPE7pb38oCKeFyOwZZbs+kv29tYPzjswBC+6k30pOL0kzaeb3Kjm
V9eb3n9Nwp9pjglnhbKdaEh6EpqmfQJ6k8LujJbalD/KgqTDZc5MXo6inr00zkFo
kWCWAuh0ZLAEX2gYaXolZy7grniunoShChYONE5mcNiLdMtQWcNqs5NhhBMA1VpL
CYyaogYf+E4P8OR4i+GVM44ceS0NDlwLbMYR3i7gh9XqJqcxdTm5sHCHpJqkRtHe
C9BH8apdK6XBJINx3IPY8+Ci2/sU/1JtFYtVWOi/W14UG5/2gHMcqid66MWbZ+Rs
eaxrCh1ic17oHAb8K2lHoV6aY9+q4banLNDaSCEyGzHIT5lslOOTKdddlZ2zrwsS
I3Pu9o4dMtBXyaB6hIRHv2Q/RV8KgdaMrM93iruynDoickHkGxnVjbCq7cfsEor/
Slb2/QdVm0TkSq7A9pJzgmaiArSnGIg9f7kB8ztDNTQXlV1AStwhj82waipj5a7r
AjjVP9Iz0G6fFEFgfUcvTEP/Kz9iSf58gtKPKqNQBfbx0u8RU2AlTPOS56kKDWBb
5b5Tv+4m0dPRATNhpVePFYzjK0NXj0wGGtlvjzbYjeCt74l33LXUlXR+bwaPUYl1
Kb6IKYdXuNFKcyEMJB0WzGoRPQfOz2geYcdHQENU9wRbygIX9oszjzpzCyUJQDSR
cdSLyWHXnFKIj6bDW1QUr0XO01k6/fg+fnP4uElLcFDgO89RzsOJlclE0QHKAKbi
v1kX0+g4sKwAODrd0J0DQXQpSLO0i32ZT/M8zA4tQ4wgYQUgUVx4EFljsJNAWYfG
oHiuFswdR/9XLZNNi3gZ1+oKmsUt4NwPJbhTDmaPUSB4qPx/GYYyA89Ca5tTfTTv
flORo7uq9MGRXIzkeGf53dsaSA9FwDAPMwZVfariN/MG5993Cyq7SHbqRTNaDebe
mdefCdjli/+1AwD422srszLbvGZeL5Rtd+GRytQ/eTto6vEiOkAcKDJdlDJGVtvl
CyCLNCu3stgv6QNItVlpkiRTmUvBe+bAn3ds3fQeXuUrJcjWGKfhmEKRjYXwz9ZQ
hghJFVAgBer4QAJyLSKZ+H/yzRihDsIBH1gui2Dhf+cfqCjz1O9Ju5GEpUU4duSk
ohyKSWy7TQT+5o93H5KdWOPBVxwsNMt5dhEgZUKRSpY0TRfcF0DxgSiCYkxGGleU
0wNdIaGHWS3a6GgTFYjLkhWZx+j3ZL5bHjln2Yqe+rdo2DNLdXWhw9IeY0CnbSaE
VgXVmduSLsdn9aeCrg3Ndd6HYoUsS4CSVFkqkwundc6JC+n5opD4c4v5Z6mqEQCn
UPPxE/9WBajLC5u5N7rN1WVLQsnh1YmRcN2XvO538hLdykKxzsfkxB0xF7B+XRg1
CIpFGlBB5RdntZRf4sZExLCSD4jwo+RhtklDGZLuAXqL6Uaxg/05BuCnCm47HyK3
riqPqyoVTdXWMH2H/d2i52BqBbuSTARztihwbmpdIWC1vLHlo5dPrrtUouIDQ5HK
ZhWugUnBQr9eVm56wzOkq9sUx5HCKEbOYrejtWeAh7ikMjQ+uQsZCWbJzxSE2xx8
CyocNmBQfPpGKS8o1mrCeVqhVJ0xBGU6U/NAU28093BIJnqInrO1aHwoNc34dAeL
+HcGH72oKOXZBz8HZRFHXTiYQBf9dHfjK5zWJZ4BMHnuDHbVbxBYVeJbX87bCZx6
ZgaquJ2IN/Pg7qiwhmaoP8tm1jUHjF80w3A2tTHZzmB6j5+L6A+FVpIwXBc7vQXf
JVgV32VR54wzH+LLWwaQAPdwF281/EChlfYy/Io3DZYQfKTEYa/FwMLIxD+dZ6Mm
mBsNji9NNA9Jn0sCwitBabfwl6ReIsCLiJ4WmW5M/duQTOIPEzg7GfOFxEJAxQt8
IxxOynvPqRbc6xiDt4cyEU3T+mKorDwrKqxOM+BlN7tyXi5/RWrWjlkTHXfrxLrE
WAfUOHRyIEAJ4p7HvkOfY7nhipyV9cMW/3UvHzIR0LWSFJC+VT25xTGTwswIVpBM
0Eoszas2lC0N8vgP1G2XGpX5hSJbTNv3dpOMaYXJDfrfoSwIdxd5k90tWhxZ/dXV
uCV4LncD9VW0g96nUCPkBBALhWhVqMHDWE5mROC6m2lIxcO/HN2CAoqTvK3JibWK
7lQSthu9xaG6i6drqEEIrsDiBTTXdefgHw405OL8OrsDRTGaIHI4XxAa/fAbmmYP
w8rCNKcwiVLUgDWoxSlmW59UXtX4fdPoV+Y3wd/T8FZS+p6LtlLXWYwhIFqHBmIO
HLwUfqL8MyNZsPuiq4nHyKSxPNvHXpV+l0+I8WwlGgns4ozAEpanrnyAXNErTdz/
eA7H5jwS1V3+wXWNNzmInDTm414Why2crJPCRthzHql+6zd+ADFkmKdmqHdc+hii
L7tmkyt90m4H4JK7tDP+AfsSHOmI+t8/8MAMAUSr/m5mP6+8kRYljbfSvagDnsye
HVZfF4KVf7HNH6rE/sYWHrfJXPAQvVrU/dOWqV4ded8YzZc3swf7oG+lK4HtPm/U
OoTJG7amjgGFxJRkjPTWhv2w8U6rZipj0wM1iLiwlSIGoPekOBz990YPYvT/xOjz
T7FjewhtNtTyrFgMAmkBp+anvJtrKgiG3AYjJMNE2aK2mpAshWh/WiuyVJhAzojR
YudEXuG3SPuqWWHpWvDDANuHy92Eliyla4ms2YgFZzSC4/qMl9l4wKLMb5u1slxF
vfZ+vyvUQxtZD5pEHFonLl55c+AFVXZXwcKA7wQuecpxtk6lnQyMrXyYLv70QqYO
lSBJWBa6fHaYQGW75yEd/Ii/vT9EbCK6xCvPjmCBwN3HCX01FfgFCQMaDFvxA8UP
KNLjOqOycn9AJc0EaqpSAHPTLz3+4Ya76EV5UxBhaMNMzs0mYmTT2GZVpT9AnYp7
5PgfK6+CFhyTuWDYPKIEypeI/7qyfAfp4kT6uHspCCCSG7wys+U3Nzfu2ApS1P6a
m6mlxgibyVdz/PDxzrs/VBo8XI32hVFtqAMsMAxtK5CUkijUeYUGa0YR70fuSDOJ
oUqdGUdbDmFZAueWSsvwQXLTpgh/s2im/6Sjphc+PE0h4my8ECKiDQQ4eXhe3plk
f2Po/4oH/9gCDqGMV7ZgSoTuegNIbggawULjr8GfCxGZUhlVYcY+SRwx1qjBDltA
wC0+/j7JOQCutKgK6GYZBMjIOd+pN5eaLgX0v6rjCpmTgAFpmf6p07A8VTHlQlzE
5uu2kcxS8cczmnUIK72NsODoHENj075V6+MXN8inbs6Q0LlWUoQ1BOFrT0/1JKMB
cUP+p192tS2d0WJ/bd23tWRleRbmy4ZD3bz0Ey2fSQJzQkJR2tMJk4g0XuoVjmDL
OJp/gOGXqPT1pyvqe5NtxhBiszkFAUwSWMwFgbVhZNxU/3GkTuCbAns/yRgwLS4+
ZvcaADeV9pP7thskbgBiJr1Ika4l0afcC3fbGohVgzrZ7fZ+UImF5uZDYVTbKevq
S5sIlw2x9lfbznLKYy2DMeE/leHOr3J1lnviwKJej/HhxTTidzxWb9Q92T9ZOfUb
hagBKcARFeo4r3GFkhl1GMBAL4kPAxDzgyDVV+IYERxhBlfwoJRiWa0IqkTnGbXq
mt8HvjOZ+VLESFrqmLbiN6caf3Sk+JbFWMTPK1MIzDDh+uA9hi22xSYzUPDQgSHX
/7wkJDG9EgJZFVcuLC+5XTqzZcovcl9zgZ3pbr/QBfBvgoBX30pH8cKl7t5RgU8I
+O6A5M+Npa6x9aJ+TsNvzB25xABGAQvUwrAJbi/JcorKEWtpB9E86UdHySiAtvls
x0gH5VnFKb7GRAJV8f4HCJctZiBZ4okr9sSKCcZRrin95PejJ5uz1UPV2/vg4P6W
6UE++TjUKx4u9duBXyzroOg0KPVRMNAJn3CuQoEJwbnM+qSD4M8bhMGJvmv/VGD5
IKXXUgsmlHLsZC193pR/sXRG2u+0ycafXPdll6qrFxqcJAd9+/jZeYclJWbXhdHy
3xwAuf+RQFanWjtBHsHtITRKBTNjunya84thkvjGbQ+G2UX8VCb/i+8lHBABomi1
DPKfd14mbeSAHZedNIzmgdTy8C4CW0NotnItAawLSQSK2XuhgoKF9+xF0E+uCp9h
wG1PrikLRxYXhR/hWWCafYgVX+4ulUPfJYwSUXjwAqPCpVRrvG5OY778Qr7eUVfJ
gvEUUhaFywAuXjUuqduIUUDApbSrenSPIv1GcbM6J9JXwHThzu8qvA+YMcSzOWOc
Db759bDorADY3THngPRillYRXluestkqd8C0TMrcx2mDLiWtyoJWfX0ZRrMnJC5B
Zhbi6n00M1BaTQx4rV7aRsBz15z/wRJHkWyCyDenuEDNoXB4Kk765WO9eBvXPajU
irTTrRhNpZpPc/WpUuQs/gmxXoDPLTgsIAxax08yXYvWCCgCczMLDGfaR6F9iTpy
A57cYJxMQCsFsLcFYKSRb4/sU1hZtx4v1YVFcjLUwhmsgkgPBolF1Y5o0n63LkrQ
RsGBFCQm7pPGOLuCo0s7tdo+3m513EPaHKwQsKUx6rlrmXfnS/boKDt8SN61Ht2b
5HELt6p+5z1Djcg41uZPGSwM4C4surRp5OvrLoJ8jYY3CNfNlsMw/oPD7N+KcdXa
swDp92HDSbrOUPDr6m24s+OhUY0jIQWbY2cDgncR+XuCQ/Me2A4mFGRRL5VbX6eb
4O4FDHeWDJCi3ItO/QFJ56huGTYvaGQWq7wKdQSoDdlJwF4wd+90W7kn6AuOMbS7
rl/VWi6F/kakzqOeJE41cD4LChZ0NKUZu8KMrZWTa2z1J1q0lR4W6xs7ISYmgZFZ
YUYRX+9vfRnsTm1MzzWNnBd8vTrft9YuyXXxqiQZacjAVV0yj96D3odnZw9NsrWd
mXBHJ2E41hinVWNPIgMyNGBZRA89u1b3Dn2fZk1lJfjW/urJaqE0qeXvmkGaJ+ym
BrofvVQOGcU3pLLqC4W2MvejI9tJguni0hmgVu5GXaW2X/0fcF5+cTw1oj5FF9k2
lm2K/tf92G9pl/KDDRyV3niZLcHlxQzCpwZPJnMD0IyGt3DCeICXjL5t2Q4IjK4h
4z+0FuCkEcwK3EMvXjLMIKdUq47SVb+4YoBe5o6UwSs69ES4CXG3sUnaAyi18ya6
6tOCJ/UfYL9m5Y88KpDHTJ9aSfvkxf5eR6luGev+ROvumksdRUD0DDelMPiKKTTv
OwFXNYTAjfLRSFLjxmFs+TJ2paor5Aq7MFJMzEJow4Cx3tsQsFm8Mi4ijef4g8Q3
qCNjIRR7b9c0sOQFMCG/yyzH+G10p/+qaXtYjz2E8mNrkUPSTRQQNuBY1oIAeJG0
TukyNDSYxg13R4YyAL0RpgEdzH4tbUmqnO8NgrpvSWKcPg3bMm/NbEUBETF4kl3u
0Qckv99WZ7pPeGZQ76211twyuqVd8dGHItkfZ+ATKKsGgbpwrzfyvRxTScI0wXCu
CzbGwrvq0mf0PkPUfmRQMosk0GOfEo/N3zhofbpBg8NilqeZuiXKbAO3LlezqrCg
02NZgPKz0HbrdnBt1qKUVqo8ltdu2ILVin0y+u9oRNURLGJleVnNBgzIWTXcHQyg
IbCjEOxmgpslYRTyVdA6lvZaJhHVPaFYOgIiOeysOtU9CpDgOi/HUxTTFdMEALsm
uA9obUKtR2l+h3YIZc789GSz1emix21E8TGUn5LBeRjpCdtbZsPGTteQMZUUQXOt
sdC8JgZmE7blrEotb1D750Htf1cIy2+ehgaWtl+/9Ck7khHx3+GXwTLUeR9AtLQA
mzXcUzr0kiV+Wd/Dy3775kKvzeFTejpbtPIYStYoIpQzeD4QxJSsk0ejt19bHE1f
cVuUetfoh8ZqtluQaxq1OAj2CfYFW8WGsNJPXczrg8NkApwPRpws1anWgntQBXIU
3sYsy4qJct4CuKfrzuePB4wzmCmICu/GXWE1vKEYe8U3wXfIMa413O8h0g/ODta0
KZ1n+hf9kCIzByOlSq8iNQ3cEZ1LgS9xo/NxcWunnEu8YL3zosTdbA18vpsTYLns
qzr7/gSnmUvtnxGUf93PAwuaLczgqumFihxoTfgxvecz9sw38uNWIdE0q+42Ta2G
ju2LeKrL02VZkAWGG3vaRrssxhDNCa8VhhPWRPMf2zjlvFrVWhiTPmXC+CWunJPj
J3lCyTiH7SOuByQxInRQjcXx5XzHH09leechjMb53AFrnRWgY9ydXyCcwTNcl+XH
0SnUV9xujtfU/D//NZV7mYpBNTwQuV59LX2K1BUSKSm0zk94pdzac6JFsH/OG/1w
ZorQ0puDdFUWx2IOz0Nw+qqHSJkTRMVYAZyBDtueXrMzi12EaP99tvkWRr7pKv51
X1/KBIDUmy3hU7bEVEXtg1SMH5+Gu28RHNGPd/Vvi/C6Csi65FjzN0lKIMKb4c03
QViDVjWrwrFDKTJznLzx3zHfGuI81585JU7QXLC5/tqX5U8SOakcxhIVL3BirPf+
KkZdPskC7sSyUe2d/BwmeddCpWuVGl0d9qXwDUs4iesiHI6OJ4jLWGnjX4WsZaKG
10kTuclbbnzz2dh/qS/0MfxhDQrzuj5UD7o/QHFZiYi2+jmxAQWGY4ToRvTVMb+R
krD0qM/ebBANdDLHbjNMpYBdeTA6gzkGV6qrKShEi8C1ws8JXeh8JyJUwXqlaMUE
wCfSqt7mKS7UEWzCwPLG2teTnf5+mm9ZGj7PdK023+m1yppI9LoyhRX5r1oauHff
0zETCwwdVnmG6KFWjphXaOpTa0l659Gcig49zWiii/12UVeI3MYInM+smJgWb4QL
deM/4lKzPETpCAx0X08BhzOAk0MteNTD1DJWMd5EREqAWtkQsJ4tuE6DkiFZm5mu
wraTqTqmuh8qEl+9a8QtvH7nzpnWJo4of1vhN5WB1djRUV5dT1IIP6p206HtUGTY
XNHzww4Ci2fEUpOZQGB5lRRYSU1GuHlcyccB+TE0QshG4e0UFPc8SZ0lC/X1NnxZ
PcC2KLTPb8bZw1T1J6sywPYVEQ0jCD8MSI/HqDKV8mPavDcZHKKULzXa+cu8LaZm
1TDEGLOAQu9XeHANAM3obXJ/k5gdtEVzgC/P9Eux1KpbUQ/3GG/b6zTGUKQkbRmx
ZS2RosdP/4Jxlrcwzo122n+ddlMk1dWf3hN1+LnRkUaxR9YB13tArE4V2Y/4cFkK
E1Vp4hZ8fZloEATZT3uV4ek/9vXtgbFKrOK7z6pmj0t/0VVR9rLZEXcD5pmK1JEr
IMky6eSnWRXSGBzxY1feEFsMAHCeVcekSMLcc9cER4mE47OiqcOxqz9UqN2Wf3MC
aoolAJUwPLOfHcEwraauDIKMQpUjoT+DVC1TJn2gxmRnbopJZj5b7fgFwuoy9WsN
3hv2aD5RG0gyvpGJpMWi2fuHzIP87yM4EYKP4Qyo65kSyExv+XsK7wutN2D3gtQX
QzmnF4weK/BQO4W1j5ptffQch7pBMU+IC1o+G7p9EuQxgzrmtKDu8hFz8BFWdQJc
i3P85vQVIK1FU3zdR+Tr/coyc8SyI+RdyxCa6PeU7yRhqgcspu/a5OlMRu0fJ4tF
nQEcupsBq3KZ70wm8IfJhm7o40iAsh88jQojEHjPcLH/5rK49EO60YqIffDWJWRp
6ZYgcc8pXLxYbi7WcC+6sfa/YtzDQXEbPgt1VQdQp1gS1lvCpzDnKjckLuaYK/6M
q/7MXqpJ/VV+Fk4Dahh2r42FV1p1d1JO77+djUi0tOO+jPpT1bDfiwihpB6ghYGA
kauD6NVDx3Zk1I5miEfnIlh+XhI3UIFJuXUg0G3lEPPZBrK1lfSY+s8+cMjyfHAw
pCqMVOnl32nvExfcXldRWSEHTkYluhyqV9UNNCBDC4cfS4cYfHRa8j2FGM5Qt24C
jA3gafFMQybGTsu8f7UHTvg44gr2/Hwz0GSRIrV57b9w65y4Ggr+dVSQ9gOg1FlO
LffJxYN25Wud/eF2SQR/pBscDpKQGp0/MhurAZZBWNTNB/g5tKLZpn7a2FjVG5Fd
az11lo936U7oy6pnYQhQqdK6nOYeDcsVS4cJ0h9xsN/pcLK0+X8lfiEArxZpkXYF
6EMZxpBTZNYbC6E31aAlydXZXCA9DqtvwFmw0DAJ3OMAcwxUY3Ym01AO2qL9Ug8Q
pgl8d4zq5bVzTWvzx/NYxqCIBRJR9nU4ZMNEvph720fZgn2uUWL9iqeRQvhnvBbc
dzdaMViwRu3pr0oJW9dLJq4ns1SlQG6MV2rbDE/oYU+HP/nHt/a3bD6s+yHzqQB0
ynKBkAyjtPgR7D9HwJnLrayBXk5aRHMdNEEvMGM6DvupO1VlK1SURSC8nc8b79qf
tD0TYinTd2f9CP6yLK1YOy8EhmhBOYZcPWq/YMune5uI407aZ6xVmoL1MYx//E8U
PJ6RObvYBr6SFGjFNCXkZTUItcHemntTKw92WVmv5Z5b+28i1Qxm5ujHvLIukaUa
ZTl2D+D8lrkx4IKiOvVNU8xPYKEq2j7VUBQFxmFnZI0Pb0b9cQvaRWEbx7C23ybk
Mvghd2C1yh+z0Ff5giTW4Uicu69DFRWHE7sm+sMZxAyPV3An2vEKpe7vG8osyV7V
Wpw3tiwd6lxHvynXbqdVH6pd5/MOOYO+bepNAU8FbdxoAnTbt1sLApYOqXeYDRLN
AHFha/jbOQbAAzyd0RIp0y+3d1WikmvL3/d3++LY919Hz1crsqDsCqs0MB38pHvW
kwt/137sf9WWMCvTiTcZOm1TDOVn8CTH2ngGvdUvSnRTSVGCIYxgobuwvrDqlo2z
WBLiQjHqDvaISbA62sXg/np0wZej+EiLHed3OtoGw5SAPLT6nl7G6O2DYEUT73Ji
H5yc8//YCd3IKinxd3j5jgt2CuWSWBVTU6TS1gZjnFYuSeEFmRowdxSJrz3zyspI
PmHYcBv7ZfZJAbwvkMAbPcDPukEZMxsWwnzAUsZrt7hPa0yWcpfITJx9hfmXifcs
FxyySFcYsZ/yOMix38VbY/f6s1m31h1a4WijFBjHpa8a57LfLcE0f7UYLS/8I238
tfrSD3fLqNmg52g5a6DJXkytf0GKv6h3dSQLZfx+Gvx7efKdmGuf5MpdyBoT7dXq
1gxLCJo3GjrK3i1bNy5QvCG6bb7b3dsrBZ7wMQVYuWPY2CmbK3xv86APhVdsOodJ
kvKzT7JG0gHq7q9IzLM98N/skBATkCjIeOATOOlb4Y+HBi3CHMBYyZjjgmyI3eaV
E/bcPfvnoclZuFLbt2EyNLy1+LcUvcpsVgjwkjQz09ZBFeUZtq8VEA541twWzz2W
adPG80/qPKsk3K9egdtbhLJRAcrUuvsYi/zD3LdCxV30ZwmL3Oh341Lz9P/hdjYe
qKwFRDEcXa4zdK4h4S4iNLm7wtMPmL7bGYjALDRC5ETSdPzX1ZyDSIuBYCZtphJ1
CCh7Ri0U09mjZTA2qy4fhhb0Cc9WV6GjuELAvUGfqNkpZlLRF1x1TYAHMsjnJoMC
VAsl/Q7SPiPTviCuc8phCGE6hmQNLmnn/V9SJuO3w95+78EYhos9u2YIbSx8Cagh
2OViYtI2pSdNu61XPJBbrSKmDlXjeEB2CbbjRp0JoCr6YaB+9bt9FTCn7UnoOpSV
S+SqVvr/Yk2ANjQ/Zn61wGOCUeDdiD94Gk8FfPweN4wDY9TuN96ww1g5bPGTOrcL
WkniYFlkdTzqn3q4GspCtOpECoHG7PeVmlQqgCuoU41m2DkBNQNN9X/wxS/9Mg/c
OESNucJjKreu2IGh+98SxTBYpYi2jQgiv4Zmm+Xj1EDSume+3fRg7I/jU79pTXQl
uWTp4brTi4Lk0AnSgQo45XoWtUOaO3fGq/T6I+uVLS0ojX25SyrP3/fZFIPu+0Kz
WFqRlUMXb+g42dbjzzU1JNC1pyv1n4eBlXA7a5DwlizZrTWR39555kA2P1++jOoX
ZR0IswVt3KjFeXV2jEH/vjnpK887u+kVMeRG+qNzGb8tw3YjWmV8xBHaptfz/WJJ
w+VmD7mSAP/ZWuYt/Xn3LtUgGhW8bzrsM3Z5JfED+5n5cGLAd5SPZoOUQuWfzher
LPmS/Q1pEaIbTo/sm6QmAQQYzoeTMX5uFLaV4py1DYkRLg15jReZdL79n5A5Z1dM
BAO3ZCtJmhRNLmVSoPYLS8xA2TFjXkxhGRCAFTbSc63NqaOoGDxnKHsflU4zJ4yy
Z4UFxdjMpHQ7SW1h86SWx/n++ymqV3SQNlmr9JbICgNiq0A+YYm7Y9MyeinumV+z
q5lqkXGdSryvBEZm87njlM/1MnYFwtjGisIvLhauBUvMKT89ZcVGcfQeT+48aDK5
IsBuoVweJ/1v5LXZyL7Ixt/qjmHN7J/9nrHeq/A2uvy6sYwpvA2uXOOI+C4ssXKO
6I5+Ryx04E5WXI8EJyNbJVZRVsK3KBQIvSaTFap0Qdfgs2YAVlfxdvvcAi+ENf50
nCAUiBgfFpKAHWHbZAyx9GIELGJilSIw3+9SaQA6RPnwKF5DD8lm8Luqlh7mD7p+
a72icJTGWlgsJHZW6GjgZxwMUTFOjMvMjQvdKPWmy/vZrNoMnzc0J9s5cKTEJD21
fw1eAlp9UjGluHt1H/AhLqpB8uZab3R4k59MXrsUE5GLeliJBIKQk3m0frNl7Sru
JI3/HAEeHpO/vH3hdXeyE3EXWY7o4nTSdWdjcpUXLhn3frDnOB2QX8oJyNvfcAmn
xxhKKuiTrHSju/kxf52dewf8Uyhbjl3nz3SUfovyYLtFZ8kzjtuikquwkirDEyVT
WijdcqhgjTmWGm9z/3dZj4CcFXmLPmUXNsWWKCh9GEJj4irC/kHyzPMd12aCOsgW
5PJpo6QNn4weRR42ClsxnFLkpCepJMojqyMZGbNd1iebv/btvh2VZncsvvuwnwqx
IfhZ0HPhT3JyQ+02siv3iZyDQfLXyHzoJtuKdJDjYnJ3uXtjVkyUBKl5fzHC9qq0
7ecPqy4lfxyjpjC2HPdNZV26tPpUKrKBXzp5aYk6TGiRThZtJznWbqdoINXQ+MWE
RD1LHfUwiWqpE6hJqDITT/zP1fAm+/DlFbjYaTDwSzcR3oGG532ruDEXZDI2N2nQ
6fZTWqbtpaqMFugEwS80iAP8YUuZ6Lry+af678B8yfBMdXtJcmXdL0B4x3f4qORB
JKeCq0ktQRGsuL5X2ndbMl/QU6uxHKH+/M1na+w+VYKq5cZajG1UgwSQqWmNq7Hk
fACaqU4dTRwrqG/EpwbKBxlj5RjcZdECipSB10sUuNHbhpKBmCSsQfPFGfiWrQpX
/nf+0sOUckxYY2h16x/ff0v4wFrRDQqHLOWNBTbBOtSC00wgYUStgQMXaYIsq3nf
mtUruRYrakfteq7iy3Zz7eCfXrBWiYfCmuo2WqvjVcCrTKQbT6eeHSIyNUt5WcWD
I9K9xd3nn/MRpGBCekN356sRpp9g4YOVCVluMN8AOC8LGOnZ1R9nlcfkaoZlcYHs
kHiZRbW5lTmAppLRbVQ0dYT+pnWvsOncj0/xJvGg9LJOhQjCcP3HmFgGHRU2FjaH
9tLfRBCwAh6X+OG8AJDsh9HUd3+OQF8UqwjU4m0DgprGnWnyzRuOfKSWjzbxHaeb
WcdZnkoQg0K3IdV7WD0Xy0OyxUeH1iFzgKO4iIXM0BAFfbZzW+mMlSzx3lRDyRLh
E8UA0ZtmacdOAT0GMYtQL02HuWfhCWQQ8MBSrxb+y/cD3N+C6jocy026W1rnBl9B
F+JXSsMJW9wybsCqtQ29vjUGA85i4bbfd7d6an3UpVLCv1yONpEBJWOdioPymeEW
J/VMCA1PeG526yl0AU+FnKX4L6YrUHgpKgMtgS0cEVVWPXoYZMBh1WpIyR0TS50v
DbYFZ1uQRLtRj6iSfHX954mluxNDekepJr7ke9KWcbRch+esd1/vD2AZDwgYpDRd
dCHOq2xOEZSV57LT47/r7YOmxggGMFPq7Gf/7c/4h76cKlC5F4ybpAj4nz20URuF
UMsuQKuUioZ4sByM6CoRHE9gmnng+UrcqsxBmW+gBC2yGPObjFv1chlhLOqN5jkO
2TCIsbwMjnTzcvA1a3/m12Yo5Y/P8BQuOfDpK9IFuxxe6OG1Bj1B+NJnKMI6k3dN
ku9oZWkbKzrHjTpTnkYyGm7GyTSaEzh/oiQmVNxeyIkDcLBqzt9ZddplgGj8V766
abQO1xWm/NY0tAsF7EGYHi/mNFriHcQozmXNZmAgTNgvLojn6pjIbOTLvUDIh10e
3Kb4fQOqwwqld8WQD48CxSVsCK6ntX5zOHwlQXLqS4EBAWOnR5sjcK0tqBLTs3rD
qXaeKGax15RlqJ7e+vYPWMeMPou0vx8SFG14y9eTrSVrHO0OPymt8zM9rBMdapdT
3EDPdhzp+e0HmPTPn/cQaYZcTMFoEFuIXVgRcEuUfw85fzC2DnqE9VlHTcVsFuI/
YbE/anN6Gmx5dV6x0IyQGepwNdccG1S/cdJ7jroflo1e1PNiQzVYzONIMGbSKs4u
ZSisoGWPpGbATKskh6NojdsFzMbi9Huh2anPvQHXgt23bG+Yr1dr2MRUErS+f4DE
zaX+nthXsVW0M2Kvl0HtDzNjry74U94S0F0NAtWwLXdIB4cQpQwNThZ6P2+cfrhb
amTXSyFByxiMSwlA+1eMZnz1Adi8qg4quxha+JfXEVoIA9J3blRQXRgNV++cuUt+
Cu8gWi1xhjDfQtGI1IwE5uwRAt+yUk9QutS8d+y4M4nOsoJigTN0Pg/HS3l2z6Bh
5CIwQuIc7GYnycngAeAMqnAQY3jLFcMwb97G0onPC4fWdy/OrumUwBxTZkQQ1fZc
NZXck73p+7BD2Fs/c+eL4cA4Q6/XYbXEktiOlBuuEkj6rImLf0R7BhCDWQFpEOT2
O6z+Wzg/zjisblgOA9XFxMM6UxWYVT3S3A9i901MfpHFHF/9ZrEqovFY+9+dD5gV
B+hfWn7O1kpHNVVL+4FntuGQV2UksMSo8aapV9ZE+kPWUK5CpAHULbFCU3M5HQiF
ocMhJh36yt1RoYXTxiygQ1i6HTKqVbNByfZ7evGL7KH39Iag02+Jxxj8lnh2vvEe
Eb9NH7ug/isYjFdrkWozJH7W9oGu79EqvOb9eQ2suyiYavEA4JApcYld9QWgjAty
a0uzS77LN/bXcFgyAdX3M+TI2SA2aUjPVFaYcbei53hiOJ8DOmrQ/zn3nPVbnJwU
tVVn0tKlFONZLHSmZygxjv6FogCrht70FDy1ufE5/ytYk+pk9QQLpZJpsHuM6vQ+
X46s2H8MinhViusWmRqpXGjWrjOfDG3O8iud94SYJDS2/2z2StmWPAsJZJBw2ifi
qTVIYPfDq7BZ8STLBkQZuAfh1p9tpfxpIy5FMNh3FqOtPMSo9qgoXSd17AnFSyDu
zopjIzHXqMACpjXcb/3G/F4ipPgAORfkEZEY3jrMCrnor9a/wBgJu63LpZPm5gcf
O2xlFr6M1VvP6JXExLfzpDtO3IbZNKKaca0yZd0ng37RWXfkxDjgovNsjA7ZI4CR
2RtDLAS3G9D/FHstIUugjeL9XwALFhmx93fUfWLGWUiEsTbMEACSgyow/PqKjBxS
ZH9OAAlu/17llq4Y6JUI15im/oLFZVTeYG/Sy7R0+mQZO/fl9WJVBqtuISiOVjPr
168HfZ5qgRQ9Kh5U+SgvYv+I9YZm4KLM6AOQC8/ylddhQ4BVJGl3RpoVQaIiwu7H
/vEX4R+ha+qlUjtkXQJzWG6dWkvQBJzO8mjW18jGnDYmlhWnKO9kDnHGQtS5LcDh
HcA2fSEUvE7/l7awns85mX4emK4uv9s55huNmMCuNah/f1MdTZVgiVUVNTkgWU17
SHSGejtYV2e2kzf0cP4TPJyD38CDRuZLBbY48+p663vAmq/jW2fvC3J4Wa/IwIis
DDub20UqimSGuxyK+faxZmNSsOwwYSQzSCBxBiKiDExdGmB2rqaNeQ3MH06tO18+
tg4umYRxilIYQonpDA7AL/swMJSc4kq3HcbkL2Bw/K6Nlp1JUOnWQuNbxIo/JRmR
m09bNQHuTBH7aR6zA036FfsDg5+JT5P4KqDg4jMS2hYbTepetY7DTg9sHG+UE/XJ
OLxZXzOB9EU6leHQz+44hjUMVHJmKdbImlCo/5+5DLeq+PxUQ0MYZ5nfzTeLQuGq
ZGTR4spxGq1IRpB9Z6i/llmv7JbyAtMkBa37707i8/M62MLETbYy6kDTc7Lq+Mcj
/al30Lqmw3EFzHlW7seLmcjYgdZdewLTHqY+5kUd/Ei7Kuu34w9sTrX2SKPBCMz0
brikrSMuUiG9QkwPIA5xuUkQZw9cNCGJ7fVuDg2H0nRIDzd0pdshhh9Rn/1Eftvr
QadP66f6aYUaU4gjwcowUjpbD0ujGq2VDa3Lp1yJd+BdxUdmRvE4cqj2lMVAEBvw
HwQUy5VSWzF/T+D7jZTOW5b9+LwQF8BoVpFuOVieL4YBQXLgTEXZEPkE/IJTot56
j+qM4aNC0VWtqKFkU29COHGjK/sklG6Z6emqRt/bp5sFFGZfdpJKNCCQTTTFv+J5
djVjhcY7fpXxnDjTO+fIllxyeqlCJ3WcF+3wjsTqfn9gGXWkO51Fh+wx1+XLRjYY
A0zYOd1v9Wge7qGH4ecZvncM/cJLFZ1lENSsdqaQAE/RhUFpQVonrvT4tUaYxe8w
hgIp6oKUqnufHLv2M76DOqfDqSPMthKMniQhcZktrn9WZPEXwKDcDvXT1WlWu+13
exDdTFfV1Zqm5pyJaxDk+JkvXo77BQj49QXmtlxHCG77GoJxO7rX7rIf1/60+b6e
9iNmGAYBqX6tLT7eFVdObOufczHDRhj2gqQtaEQlhZbzqyvfQoXSPfyGKjSRnrF+
HD63vWU6EVsgNekQ90DM5imW+IpnAwl23V8n7jjx1+BPSK3vP/DBLl209OYOd57I
qSfSP8o9raGC3o6nhGoFq0xQN6V6Y4ZHav8onJN3cMCHRzcr35gs3IPpUlFnwfx1
40twy7VN3ZLfLzn6YkoPYOHZTGtWhIuZLBa3t3wDYP/HM1IpIW1qJeU+3DtkQ+zR
8Ztmaystvkj09U3LjNNeCOb88BWmzbzDI5HgP8jCBY5Kl7RkAGfHupIfeTC4wHCz
x0xrDdLhASHiQV/WWq/CtVz1qSD6ewu3pGv6CgQTxVVYI4O5Ufb2y2RSvs+8KKZ7
Q/1huQ20XCCYsISgvDqiZR3TG0Vxi4/xC5ptQB/xNTy/oMVTGDF/ZyPufwLQGcwd
3zk2WlFsF9JkQuRXQE6IXARnPCTVHsLY06aeDftAyJTrOu7SGOfpdwr77SsZ71cN
Lq0QQA5G/z2Sa/FnXbrCUkGCZ2POFj1+cVG4F1xFWgV/vHdfqg+dFsSXjPeii8N7
Xu2O/E2T7BDun4+ZU4/4UbrCw2kh9mEFK6npf8s+0uiekoIRmCu8om3fYOTv1mfo
UG7RUu9IqlJDchcVC6k7Abd1pTZ27MIxWJ7dPm1ml2C2AJuqeQcbO6WOubRB5AY0
uPc8CL8imXLX6DCW2pLXqMbnTelpMAO/1FQOAx/+2qy27+6oU9nryXlQMRod6j6q
6CB3i3NTPuk/268GOMHWitnGv2M0VCxhBQx5/5e0G9Q2axxLqc89eIVK1jQNmyUo
1KUCjDLh5l0w+WxPxyZNiOSds3vv+KeGDcamHfhKulIB66uIYnbkxFtGV9kKKAiK
1qxgAZHoL4X6LiQ6pAjYhflfeA1WuOBn/zSCuMzCGyxQnOfQFvOgkL0yIgNJeHUK
QW5V0zj2xhO3uuGTGoV4r/6sdyDqEJ7rveimqvfc7WeU4cP1jLJqqhDY6Ys/uSMG
ytVC9aKIo78k4x7QqmjTaRtqrVxKZ2fNE/0gKllSvia00CF6WdB+S9roCRmu39+l
RSUDK+abY9SeRG26SFCF98mAKsW77YufwRBguIB9YLcNnwNQKtehathnDz4/2ivP
ABlulHh9MfZgh/vK9eSWfU78qWadX0wkHtMaBL9nNIgc0dKG7VnqOOQk8K73In5k
hLs44S6SzmODg2bnyn0/KYkcYhgngDMSNzV7F0GBSb6O23aYhEW5WopXZiElNiRQ
1NkCtPG5t01XQWHTR/GU/r86kmABn7I98Vq1lpndM1GICxPyVT5LcurisJRpFgEx
D03mDOV5GbFpVB13Ew5Pwcqa+eaJVuQH2kZ5jE357kBJXHXkAfVm05n/9XTO/PJQ
HjMPrWQKAWRwPoHTLYwv+dstLuULoRmII0cyXB+Vkf5hFKgFbsyWI/KYHUfGqXv5
RdbrvQt6Rd6XGVAUC0ay8pQP6Ezcrubh9JIwJ1L7lcyffAGxpPGQ7SOeKEl318U9
luXiwXGczf6okFNkW04Xn99HNJ+ZKNvkjTDVWiut1ifMmOX5NoIwtqLJDdDiYfdR
L2+CsYZyMNGmlFS34792r2BxkE+DHngU1fFBdP1ByWdAXn9tq8BRE+9zNuS81yiN
k4doRJLmzExP/4oJkXXEFkUQNXcwWfabr8FCw3VmZlhr+Qe5lA1OAxqPEpRXn+ZE
7sQpEHxfWmidPkjeZLUa0lC948ZZb2m4W7bGs/Iz6tOL2QZwMwi5k2QblLXbh0vS
d3NG8w7lNAcoLvt5mmmm87EPA3n7a4SULEYl/fRD7zD9it5QF7V2pzDRHsDEQo7v
gvmrNogMpluAkw31hmaiuhcfs+a21HXLCDyFLCyYZbxTFGWn41HMnwC3ME+b+4yY
6DJz05KIPuIu4QcYqDXtJ875dw6FE8MgEhqj7qpwb7NIpOykOuSbuDipw4zYRKEd
kUtZHuwYpkTMCDJptuuiWR4d9wpRH/9GnW3peFMXbtapHUD17+I1fk+ohJM6GbdV
m3jcuP1N2fQLBR9+VN4/CLTyWAJXIxj8ThxEd55P0bQwZTDr9nm0SvqlMt0k7dKl
Zh1mO1I38AV4B2WkVke1q26wqYbwWtVtHbqU5ZiahRToE/ocS8wJn9DUYDE5X9vO
F1U/VGaOtZ9ELwElp+1vokf7LExPw89kjZ3kw6rU4hCjToMlTBZlMqzKV//IXLGk
/25NB938Hn7CzkTM+eIfIk+t8hvCj7237PXT8eJWVL1IvpPEXD+1GVvIEDf6D8Pu
EjcagpdTUScQ32u3yUdajO83Jpwg9ak4h40Fm7MCAGcF+4e4UydGLcg+1grZI1rk
USLU1CZhag7+VhTkLH3YjUwe9+/YxqLl37mL4ZBZBlZ+uOWdOvaJy4VImzVssZmq
IXOFhf7qOsYuEJMxgXM84qoRSJikNiYXugj9bbSAbe5uGf3aM6Bl7RbtRTYzZVRk
EzXg1vxBq76TVHzwWPKg774DsqJjs19rA29NRRRjnAYrmr89808oGeRnuEjnT/CP
BwNhNekL/nv64EusfvAqGyq4RAB9rLaPuEG6TKtAK3ihRR2ibA5/8ontt46C6cTs
omKlp7qVWkjtbUOaalczVY0ILD9pP1zloUVCgHnhsVLIc8oaJieaeMCZrVj7ME1u
FD/Oi+6XebEeXdikpwRi8ru4nweoGmoDgUiF82qt70qWWb9X0rEXRBTmwU7+dhh4
ObQ+oWOpbXCm4z+ffxjZj4XrJVcyifIsmWcd7UNbTTbfvhuSeBl+0Pn8yURY8XUr
xPPCYj38SoV34UzL+y4Ik5jiAwdhc3Ak69TItNmWHjfK72nJe0nQIgaLoNbQrFkw
b65BL1RQC8f+jLTsTeHLIPLJ5BMbt+pJQaB2Kp0xlZWYFuYqD/c5EfyCFAC3KUG9
J/ruxurSsQ6db7T6B34BhoDO0JO1URs7KenJiEf8g07r5E8pmHp+NRKxxYX6V1IQ
WqvmAh7NOQ8Ffw6XyVxK5t3TdGScTm+8hOpE6pvEeGEJPCk5Tn8lP75LNWxjBKh4
GoCn/6nYOXEWqClZ9GarUhsmtKAr9NBaQ3mlGc0MI3oKbnmL1kc/Sh3RI6XJELkR
JI9vDvVJTTW6sGmWQdNalTqhBsVnVNgrDfEmg+T8VHc6+dNcKgYSdUxl09XwavV8
CQWxl4iZN4yMBy3oXx2IpRZ/fjJ89PAES22YLylJMoNh6WFS+0xCwK2bxZeoWOZg
DOCMY2wf+FMtYxKb+Fz2c7jA1pMbCt6gR/FQfsrETqU3bLo/akx32XoP1xDJEMyh
e/OB7FEHQSt3372s45JjwSPyGaH+zcsZl6mJJImtQH4V/9e/WlR3gS9g07nGtEXp
jrpCsuFFjxV4ADZbShSu4Ks5eE8tYdv0YDlV/ClD2Z7CszzkI9i5IW/ctWVbwdFD
t8RqtSTxkhHhYmXjj+EheWwQgCF+pWGoin/Y/MLvwkknRA3NkDWzLm8iRspxOD0Z
bhPDFS+TgKhvDBPSH4fxjTZYNQFKvQiK+PC6UTedVgn768OKYN+SdzHbrYUZfpFn
DYsVowNk3Wr2iFTa1MRFEiDubnoZlHimFerGdtj/fVyzjixtQPSkvW6kUquTVYIU
p8hRJnzUe8UhswWIVcpyKwriCutb9RqzK4y301HoLsCLxdZcpaQqPRjQO/LMCP4E
4dySK9vAgklG3s3ExzEef5HnF8Y7tSNI8oewl2uV1E+mrfatz50YSY6QOkH1B8+A
6n4JvuF1uWjS1zfbnSyKPowwpy+fxntmws5lvAREEKCUqnKURM4kthUd1aSZzInc
3owCSW+dR/foALWXHAfJxso/MNEg/xEzU7jprZKgmAlIGza65fGZILglYpIuqFwH
jBsfwmD2E8oQgLN4JQ2+bODrNzLAWQHo/lcuZgPamZPABQOnM3gTq3bJIg335gf0
4noi+iNRQohXFtkbkT7Z060/BwP5MLt31WNpqckjo++nt93RRHJN2O2zNKCHHqRy
OjAXQee6vMs6WFlinZ0FORIb9/TrV0CeUUP7AHchYVe6Xi0uQvqwW2nKeKvjvNMm
MKrXz53ke+X3f6NhBTuN/ABjmGXw78YNUWMqJ8hCv9Luzr8c3AOJwy/KmjsI6+rp
x4J3omlzEuzIdiP8DJwMIztZuSvCs12mczTdKSAXcoCYvujmHWW6z6yYByvMyAmM
1bStIsQQhTHIapr0Se5IjwchBHr/uJXpB3v70rokQ3fiWPJBlfnr8cuFZw0ZkBaH
27NG+lfIvOCApLAK6Nw04Oouq5/1aqhv9yHyiuw9WQEcGa0ubIEj52maJjFbU0Hu
a4/4jCkYVtpFZ2ia0L6qrCRCYuIeuo3OwHdaw38WVRXkzQu75h2HPVxvy/bU/E8i
hFhF/UE1bTwxdYCEPEs3hwlDMSvVghwMLbMouK+TFi1eLFMOtPAk84zwha7OA1WP
g6BzHzhORuwM4XUEJfJZF3A9vcBGjG2ZqItgJW1iEMuJqV/UrtG10xanvcftrtL9
vsOCWluTy1clSKI4gflA4YKWh0ZpwwU8R14BbiXGJkiCF1ayHqZedd91x193sdkt
Ph9v/8METWiJBS13D8opBoJDFIjcjCWhKmbnWlDM7relNpbex+eeYGUp8K65/r97
8ae2xCnZiXyTckpZ2B7f8bubeQF8kXp3VuazSCE9x0VB2JXboNtWBii2QIanCSsg
VfNPBw8FjoTb9+fbkcHGsUMRmYohRCV3v+WkJVASiBMD0SJdQcJKMt0JxFDnk4sk
ftUlKxXQ88kutSLW0JxdmJg2i8yzs+Iqp99Wqk/qwCDNBPymjk+qVqH814YlaFC1
KWd/a4QTYGbTkgq3mPpRahHlNlCpvrBKL9IObwxkiSxxsOliEzoHk3aVZfrefPkS
WDK3vWnw22u/rrnWYsyZ8IGzWDpE/Z04OFv4uwVnno8LOm7pZjb0Cq0+GiIVbIsu
qh8gCeC8HT7AtqhQ79i0Ylul9QoypXqoaJzcz+4LbfdEwRHOMMI7rB3io5dg9dvs
4cpaNbK0kCNZ9WOhg0fgmnk/1PvZl1JXMbveKRlDuwjT6dpvSO4GEsWrxpu6bBD4
w5SprVj27hZK02Moj4YUGTEJmdNAfBZTAPYBHB5c+1vNf+lduFwrw6jQb6FXOpj4
z9Juv1PQDMx4AGGgtg/iMXJePAtLhVNEuHb8Hy4UW1pJ14OlRvc2cQEfcYMK4wEl
QRzWH7wkw2Pu9OBuVAnT404yQxIsZO0QFYD3pIT2pLQeHns7SReDBHfhgb4lv7W8
3Nwe/cNA2ZvuKzBXlzWf5AoGVxxu8W4MrdcSTFn1NRQc9ShnALGpt4XbAn7h8SBG
YnPyvbs2p0SRxkV8Y1OyRNxI7bEFjl6dO7B9/8mf1RCMlmK8KsfrJdQJ6Q1VoW9n
BoiJ0mOirjeWM0myp/lo6686ngc5LdpCgCLXk1rZiPaFLGW85t36g35SUkeP3Zfa
PvjvwRXfMTnIq91tZfmNM8yaTF6P4bmEFCtr+nSHRsF9rpcsVPSBr+5q8sb75j/u
5CsrNQiiXjeUt1qVNjCxUhfl1VfbkaX5Si75L8InKUduNvUx241Lb1P5/KsgTtpS
dJALZys6FVuu3yy1/FViGXP1FBxJKQufqqdRuquqoVW+IySAqOx4sMFCAiTozzfl
Lywa+cK/dm0qVX9C+0x3LAszr/31BrNZ9qXjbutteUILYr2+Ia31GL7opV85i67W
LM23fmY7LIqqLDA3aiRup8/oPXOKFUl0mL/MSiDyX24FeMMIPhN+gZ108Z3T8feh
9RtofrQF15EfkHgKWnIwMyst+ESoXbH4ygKXpOMe8C/uAz9mJYW1Ii/yKpPjYL1Y
/XFXo3jzsA14tXY1jozrHZ9jb8HNwFdjA71s+HzFelI5wn5Q2pcmynmlDYZOegYJ
zm2GmSdj+FwRkuZQdw8JUMgZ9NIOH24TPp/v9Qs6j9wh7oQZVctn3PRFodyZdBVv
FyXeoW4jLjcm2HxaFGhCsIPZVHqjXglqLKfsdK35CadJAHBoC6+wNaxtn75KliBv
8lqYsaE9uTs2veGnI/d8AfBc0vMP3zuxa3q8sQzUeX2hSEdBpB+o0P9QZW31myIF
vE9i0WuEGkg1XMbAZNn00r7FKjUWkHIsAkuZxZ//7jy9Cu805lUocOv1SMSPhXIe
xXO324m8xs6iZ7NLtL2ncmwYjRjU1yNdTFIw+LD7TQr1gOosivydAk1nWgPm0JcH
MHAbnSp/Nn8vubDC2+f2wfRwRH9yzRRpKVp/1Qg68vKC4snv7aE1MTQ8tKheWy8X
KIC1Ftv7Bh7Rb2KdORUM3eSuTjGaAiOrcRRXlHmECUnXD3X1uQqcqh2sJunSb5u7
cBWyCuts9MoG5lw+LgD7x6Q5MeEMFWLQO/kiOdLUIOs2+1tAYj0XQVShY1HGZvQP
8BlvYq5DRaat6SysJFaioghxaA0sux0hB/K1vkHcB36I5fG7TEIcpacyHaL5M8Yt
z4E7zsc+otVcS+6ljjmHCqjgeQp9l0sNk+c64TiZ/XGM0dImVwnuXT8kE/cZCfow
PsJtx+YYeq7IJtQ67Q8B7UPzKrnt1vQRqLanJZHSU+q/JdW6qf8HnVEbDZEVS7st
ZsS81rGvU8U1lsjc8mcmJgOCmc/bauCV4qoDehQhac9fPXnKQ3XNCm74/g6e6AAF
fSEJMfffsJCcdF7KLabnSvoAmpqtJABiWnLqCccCVqakMPZK/RnJZXoo9nskpnUx
spJ9c1XVzcKIzOjL6TTM9tUy6p3l9MEIaHHgiIHdOxDVOBED8rMxJDvRtyW/W77h
nbSQozAFrJCBdH3414a3T3pJ1LjiAG0Ui3TGKjqRfinEZKleAwS7xwGJlnD6aJS1
QvgDo+Cjn2rcN7bq/Up2EfXdYXUyzC/rpjW1QmeVA+hzfaw7Au1s4pIfi2hKJR00
0tQCgAz2i8hzKvZxMbVSjkCEU9+qTZ6OkNx0xWwy7sU5S7y/eLeAGq4QHwu64aK9
si2w/7KkZqjHelhYOt2FlsmhgIbefM5dDMMszrypDywg8XxyOwm350Bortl+dd0X
uLg6M0enZtuQNV+5T3sF0dXtStUZMupRDDDdFCRoQJ9XHOjJ/rJXKSQ7RZOIteZc
3m5CYzHQ+QWPXjRx6jFLhXmEos3xeyzCG1on2mu6t4A5vjcgxfwEZlOvfAGizDZ/
TYEWBS4V4h4tq8IX44wD8CMUSjKZBftlSFIfqE0UqtjHMerkeHVfk00COw3EtqYe
hJr9IC90vYkjGqJbb1AX1eOL+QjC0pRy+UlUNKHHHucEYzCvz9fhm7PXWOq/x2k4
vHkzk+jjZpff2FYm6zffBi7EyUt7nh54Gfo/lxPGPxXloEBNH2wC3d+hdvV6tFH1
9FigpPTbB2vtWa0wpD3JnYqTlcP64xPz7kIMpM3dK9PGHJHObFU7m3BHXiQIgbwa
5tN8XHDUE+o68y2GYBa+To5g248+wOTGGxKeZx1DUZtwBaxw+DpVM56H1a46Hd4g
qooG4GZAUJ2qbr6ust6ZlqgpyvhPcFE2NWbgWP8neVXtuzbqvDRDyzY2tD8Pla2o
uufD6nMVPCc2pJVLd+rEoBaIDbW0OBQ3OTgF1hnwl0KwUKnBnnKmAn6Efd54zFqR
KXlrUcHsgKqyMJNwUGj5JVs7DL4lAkb5AZiY3Y62pckAo1atPT31Tvhqu23Zk2d9
kXOvCGmyZGfMIgqbAdO/4SVz2lnOFj6qxNBBQl/A6RIXn+7Q+C1CmTGWWyCdWfz8
bUS6K7TUFDfYhOn9OSlDNOoAilQtv763LOqHZQq0c2xZYmSwktHtgYhR/doxY5/+
2nogLv1BGO9DsmLUWDcKaqmhztbB0Fn2eA/VN8Cy9DZuxt+IP35hQESgPmK1+HzX
+V2QaV+TRpKDYzmi4blLodtpzk/s25J7oNeT/69ORzY5voeP9YeNyXDzG9A7TvZ9
cmhp1egg3c/JM/ZUl2X5R6AXZdSkjdmW0+x/yjvQP0279wOPWdTIekRBdoVgj7Dn
x9fT4EBpZ5j/WsH3G/q8X+AaWLEsVhbsKMQwsGwQNDd9+BXXkuJJD1A3WgzgmKkn
N7LYx5+m39LSMkNPv546LwTzA9RboSY0zd5SSRbNlVSHcORI/PndnUSP7vxSkjlW
hooPH6i1/WzxCqRQgGRhirF4P3k0L7Ofw3sawWA7m9TFOmX5nI4eOwjgg29R3Ocj
xVoXCoi0W0/Kcxzpc+iZTAONPwRU14eqXQZxZjlxsAv84BWyDjWlX3xbm14tT5rB
k/JlyoZ7Z0XFDumUuVfSEJcNNSDnahMmD3M/vGbdRn5iyX5OGTdcct6UmzFnzh+P
xVfWX2jI2TfVdfz3Id0VBkoF5FlD/i0KBFggs2rkK0kppj63ykkZHZJfcKJwQzFy
ebmADPWF/kFWUgo3AUsWjaeBZrbJbNZj+OpTKpnwUSnftAXu1VnUlILfsR0R3c21
9PTPQo2mVnui/IsOFi4cMCUzc+Vy16DZ/4gFwZRvwEkurtl4nUnRfIPcc7z8EwVc
xdJ0rvsa6sQzo662Dmw0NbLvZVmLciEElBRchZ/AL2RZeO0yp54+eOASpf2VToQA
yufPGPEiWn48vmZ9vXQczcAzqI7QokAlUyrYHHaJm49guhikakS0OK5W6/+oUwvQ
6c6kChB9uVhgCkAy8Qrugzngd0Cjhig/GVP9g9zasjxsLoDYKXn4pU3+1KNHOlt3
Dfr6hThV9p8l1o94Mov3ORhI/aD3hUBD5KVrKVIV+AMjGxCL9Kx8YnlhaX4HZoLz
XuaemDWdcAiO+ikLBYoaHCmjzr67jtDS/3d/FN4zeKe5fod1aCQZIv32f0oVNTAi
rdKa3w+OV4jLN6ItEXmb5+Jde8lcYcBSOihTYsO0Ddr20xyzqwQDhcH0lM4K1Gii
uBaG/2M/3n4VOf3KNVBSW2NfEivKLSp0XlDervrinfubQ/bfpxu3KK0Pv1i7wItN
vVB8/dEthoWsXnRaVCfuu8/8nJ7DHRZzGw/AybySixmUM2oeY3zGyLZONUMgmTD4
HtpaZYfJJGj0xmnfHFgrsotCthdEh63fFH+iVGHYNyvq8P+x092JTMnbT0hOMzZ9
YGf1sfQfM3b9kE8NVfZQsGAhbs+VkmUqE91AY7frCI6EjIvejPAJGj9uNn00fbfb
7p3K+3LQc7Nx9UJG8vMXSBQDJq38bK/Weqw1I3Ha+pgoMmhx6as4CT50+SEMid6w
k3Cs1+tu7E35htCitfSODwAifjzMxAuMzrxLa52ouTUUdGPbGbhDYIqFslpEcXGk
nddEPOPXqEYEzEVfvdTy2mK2hp+nnkFVEb3bfp59cu9el+hsoBa7uWuc0Ck6wYuq
thrwPWoHMWIAp+0V/6hz8ls7uS/fF/Ly2QL+jXt3lwEA06O6XxTvLA5S9NU+5Ex3
X0Nxv7IPM4RhXzh3qP+7WITyjStGadoRMdv6XY7ZTEaILcYxLC4NiafngkTDt6fF
cYVXMNMB6S3tlE3KwgbJm++i3avr/Ku7BeZItx6DJo/7dobp/r28TLAjghB3RIEd
AQo31fH+CpbwBMD2ERE7Pi6b/4GVCpS6ldqYdR51JUiI9RZrfQ5fe216chMwqwPO
jJbhXEhgcqrFIZxHqc0F5wEBNUUBcd8bKOT/n7mdNuoyBtz5F2VHRn97q4KzvUB/
Y6BOtGdfQiLeBJo9MZ3bqHhYxRlzeT9XU4I55XvIiSvQiiori8cVlECi6KBZ1A62
LHebh9zM87nL6JAVOrg2alYLRViMc9C36SZDPYZK+OWV54qRgWhYA/npzV+sAhsO
Qis0fYkakpaAi3gncoV+aRkhm9HoGp8SwHMBiaCCcRpalYNRRGJWW7mPKB2EVACu
MhrSSLmimQ7Uorh0p8yWzwXKY3hd3g4e2CudZRM2/v34RP8WKpCGR5TxcOO+H2kb
dLR1qZcKZVjEJYtWf4A4pKFvntcHSizd3rKpz9ZJ8U+2LmCPMZRaUvpX36JgkB8X
eMDf2/o97GW+jSEwNCjEQDCWvk4+q3UMwo/OwCVFDh/JqFCpwVzRpWGzhELSpcIK
ncg3ANq0xv+LCrrp2AogBTTmLPzZtHmdtaPNehU5buzNpdAx+Bp6Y8Hvjm4BE/3p
UJMKKgKocD+Du49DGUzijyLWf4pxQCwLzGSyjCirt940dloxXFGNKw789pCmJDj0
Vn6E+pkLGcTrCSWz9xzMAmn+VxCWVK6c7x8JQBPmFR6oejxso7UzHpGSvLn2MITc
SDoMpOZwqS7BQaXGeopBiJtsH0TT5I42KYTDfYhIlsy1hSVYaUGw9xNayB1EbleE
paYYOtpL83PuUkZWe728DRJgf5WDZcY50BQ2SK9pANTHXI6LCPLH2VPjAA8r1pHS
yIt8yomYzEueHhzY6dH3WX7VP0kA+072V+1OvVgqp2lvE20UexMdLZVMigZnPemq
yu1tKg5/L70xNRNrkDT9RoIc84pNltHDOXNbNsy3Ys3CSclcIef48tAzClmPclh0
HIRd7dBsvkn7uOu0D0vCPVqeH9uKrkPYv6245GF+MhOTG9xW6Ou0a5fciJfksm6q
ZylTbeZxACOVCsuUOA2OrBq/9cuXcNGFWRKl/c7ef68Bsixr8FxoHxAgcXmYCInY
Ovib2geOQYQz9qOXATwUSCL1DZ6Alt5de5Jw0A49QPoqWx/qZSLlNvlej6yxqGJM
sZY36ehqE5Hs0WTjhyxQWs+t85NMDs97NWWKvvLVvP/zUu2YGeafFUUjM+bXwN2o
BYSt+T6h8w/uCIknD5TGl0jN4hvtDwklII5IUpoRITfuusoakh5zDhQg/6UboHf/
irvJM/wiCLJJwRgCvC7TIEyhdGu7/c6gxvZVFO3AxPZ60sjci+EbkKzACigv1ZU6
PfHOjmcEKH3Jv5BVzjrUkPABpEPtBgN3cbO3RQQhOvFtvMa3+9cML2uL7crfEB2U
6i1P7z6GIXJCE/jczAc3wq6kT4hH187olTXXBUvjADLwutC1Ps7praWlqcZdx1Ej
yKxSjY5Ji5bVWLwqX95nwhXDGszbu2bH0BpmWutH1hk5OcCoeEP1J16We5Tl3pNM
3Cs697pKwiAMfQp/Co9kbJCrEeqZhnqjDNlwt6EuyJLeN8MFygjrvPyNpCQafirP
5k/g1e1vru6yV/1TK4rSKgq8NXbpgtFeZVijsKtJdDPs23lAVzzAirWQAsjXGxte
xp1jhk+Ewr0Ve9JdKVLUQS0p9/UqMqgGihzBfko+RyW2Xpfc3qcj15wgT8jbIUgm
V5nggJgVL4vbGdWlLGuMPJN8c4sfMjqOy2KDe3mpf8P02kgLC4yq2ByDG42R00MN
vDXtTNcRXF6aq9DdtFFtqbqIyyj5PZnvGf+6sLu7d+Eqt12O1GEsI/w0xbNUPOUD
TBW9Ka6rfUhvcUR9JBMW2Js+F3nC0H4KyQOrvitBOaqsgrk3yoDbDmiqu3zUbtrn
vXi7fgy8RmlM0XXYm6OkYGvwVkgSMbnt8f2QUhAiNbJhOHO7+kVzMazqsXAXQCOR
VVdDAOF34mhgTAbLk0VGm+nyV/iJCcthTv9uBZesrG76/tcJy5zENLlqsFwpkC0l
rzlAglT9dIWp6BQhXWUapRDCRM/5TBjCbCqfgptLrzC0QI94mHIz8TDAlHMjKtny
J1rdVI8VuZF6wxHguleeaCNJGl9sHFmII39+TDEoD+YIBKzpPNkfWlHZcaARxfSo
Ew/IuGYEfPgbxzXtYMAVy6SlGsCmVuoBXhR6ESxU2IxaGsUtR6sfPlcKK4ATXGJG
6m3SMHpVt1ZyTdtmZKOiFLs0FvvjrsrDUVcpWwu0NqbxQQeyC2YQQwqSxJULFV0P
dkUWLC7cVsefVKUJv41v7P1qrQGnIhInkf7Tezt3hpm2HemCrjfGHVNnWNk3/xfQ
4GZPpo5mnW1AV6mSFsjuaKyDN0qB8At3HqZCRt5g+qowKabN59VmmI55p5TsIZI6
COSVz5O/jxiZg/Z5iXEKINN6yCoolcuyRVhzZzLidwys37GejW4H7kyhCYv1wC0j
RwRww/vzBURmXDVQLfAsEJNxLNMf903KMfkZHlV5hm67E2QJxbFJ+mFPE2Kvmy39
IBQxQeNFcoX4jngDQ1hVxNAUCoeBV6GfXGDZrl1gMn+IfSZk/Zf+sBAEYFFtfk+w
f50nm9EGP5Gb1dE3xjfhd23tOZ1LFoxCcxGtsZ8QI0eIpYzv6RpfpqkVqvH6bijC
0daJTyMMX9+vNsRd6+Izb7liqUmuyRCYqxr+TfKzUE8iwnBNcpngNEKZdQA6l3Dz
acvCZCsSnPoMyQa6519codcprmbFdNIvqsBqx/ycZe/5aUiyIHK735JSqVsiGM8x
x7qp0PTrALW5ZCADwtn59/5FIyLwsEauEyNFj8LSKYHCL++EXtmMkeQkH5bCsttE
0zKlK+LkHDY3xfi64mHGKydNn2ScOn9M3Ldy3mV1oKKQlmN7mbaMb+QeLFHH47dj
sf3bXfX+JAC+3KIKYWlqaEJhEb+yz3qEIV3fhApMUhhyPDVdI7a+rz1uxzDgk0T9
8p0PoYxrOOaH97Lgya5XnySSPtNGepaM4J9xMOiHwN1wapXOalKbP9EkrjaFvoCS
WRQKTk8pIeHNmokMYeclASeTNhWxidqWWFSrrgw8JOtAuX7E178OlrKOFfV6mA/c
XH99b+CAn/BUkk9iY8B/nXQCBPCK8oi99eT41qP4DMC5eAIWP31fBYOMbjZKABvx
P2G2J4ioE/7w1hGq6mpDWnhSLg190vUQMUm+54umBHV7tcanRlObtciO5yEFsEmu
R2I8HAukex+ev/99r8I9MBtTvOPk7k1XAzONAdoVK6oqAbOymspI4lNFKbnWGNrn
QGvbmPg5WuU6uZhDtB3eJ2f20SHcV2a/AAm/Ymnx/kmXSSTWAxNBNe+znAX54ObH
kYNqPuZyYB5aEfaQ746jCnoqmCmvUdhFDZF9BOUzCLa7fuxsCaYvtbPxSJEmB30T
STwVqG8sREr88LewHYwjHc2FcZQYUcmsTr2mDysEjiPqz4H6j2SGoQAsA6Yh4UyV
kbrAwgD+5MqGcuLOUnAPI1us4xp85syMjT2UVdyU5HZGmVYafZhQJNVYg1jL7wf2
HmOYpAP57H0OVq17MpDbpFKyeRN64w4Z1vdnNkUEawFpDZrfcAlvPvrP/a5vD+79
csaM3UPIQyDYoXN2g/chctD9ydhXkIJ0HrNC5iwW8TR92ZlCVluaXgcsbjSxRlMV
z3TyEyiwAF8BCqh0qM13FLgkEHx/U5s8TZuW4kkUS+x/J3rRODKXalgXa32XqfoU
bOvLJ5fE1Q4pBz41MQA0AcefZS8BMJjnNEsfwg65zOZmGjt7i11YyETAQ+sKJaEu
lVYJc3w7xZYeHZUOH32cgUylptrVZSQM/daa1OmhL5cNcYcnyYL8bm9eq9yQVkLd
WfO/88NABvl46+7aa4XDTV5rqt+jPQLZpWp44HFy8FBgDOxdelINgm5xNQLFmJID
KmtUju/gnf3jXmjWTJQuNfLTS0r2IyS3LpbdjTT+vKJjMkKKumPl70U6NGz0eMnQ
Xyc788AQ/kdBY6B4lG3CQdvCkgCND4nNPDWUM32vBdYDKjvVh2ZpU0ujBKDQ3/1v
sTigB3JmdjYlUHEuLMkju1bPZ/ST4B+vPIRVcIAxbDWcjK+KIWllct7Q5re1prZS
SnMMiyDCxlVsSncSOGlBBx+bA9zmLZy3DpNkwOAflAy1dwWYwGWRuNB6VvYbR07k
y0q1+tINyONMJ9mEhD7+gMa4HS8NVg3HSg8MVwSOWIVTZLaPg7DvbrboxnUoFuP4
GOxhXZTHryVx6G0//dfky+9JbOqfmx0L6WoiB34kGp1j3zgrTYs9trpcl5SJBR2s
cv9HXj5z07XC6GW8464GNbbjKqsVRxl4jeyqyxt6h0u9HtyD+5wPr+u3fUIUdff2
XIm9xNfY3xEBrI8ueT+Buqjm4vQXe+Ph59st717ueViozyxsRaMCnB3jqX8OVCSt
2hDKDYWTLVJx6HuzkfqXJEabnIzuUtcE7h2DAMecTbIWudvKIF/Vfpn3pFqgZNlK
b26j68EgAgh4TTWvQnhNtuBFZqjkD4/L0XxAH6M7iaskI3Y06hnX+5RnIWhck883
rRo8d62vFMNlyf6b+FtlumUrFQMJ/HZ9fgEcmEUJoxP5JImAYn5teTPkariUsHDv
0vX+vkBJQi7KyXIPVOX1CizNOCtIlOipB+xuB8Q/0r0sDrkyJTE4Tqhqwqz4HCA6
xRRTDnQuac+8hp8bJwOPeX4VtKQvggxbLJ0aCK7Lh50GThDsDwvEZ7yqtjPDG/uC
XaS3gppE3kYpNuI7rJUT58tjakRKPZAeTNufzwOA0vo5BzPcuVvrVj30ZsnF6GD1
0SVYwtxnnqTGqY8pvUvlq41IUYwysJSY5AG/a1nyPx2IDg4jiGkSFEA8rVOpL6/c
tA8+S3GLUMBLZO+om2YCglMG+YF9UsCynSZ3i0PMZTXXxwjRD993oxglpQG+tu+x
M/ZEqQjFdW9z8XmapQUgn6cY38Ym8mC4bqgnIzl4RJSb+WktPiEA1Ae/hNKVM7Yi
jZqn3YWWyV3MBU5V8SQDcgTTdROhNt4TnSA3C3W+9O4ODreY4bCNy8fvlRhtbQhA
kaps2L/1d3PWiLUaIDkvgpFm0q3ZemayZxaTq73hikL5nGD4/QfgQz1g6az4LRab
URgv1BFYrlXTL8y16fljLJeOS1w5qjpgdzKhuEkcNIYukopSNUWRifrriFB0Dd5L
tVYlXHWEGAkOMYx0cxBe0IL0+r4ESuqObOu/2N9Da/V/JsAW8t6odrWSrmy4tAbX
MW1Ho1YMo9OCmUE+ZqSkEOKB1A/siLn01u5x7vk37tGo1Ybs1pfudJ3eoywD2UMW
ZJex49i69o9RK3PojVa/WX95TFdebmzskJFvjyVG54xumum/0Vc0SsLnrko/vsIn
dE0PT9NNR0ETt6w62eWop/csqz/KprRv8y53hwX3osOjcxq0p2QyRl7OmO8YetqD
yUGxToq1PW+qq/zOxTbeDu0mMDLnZVPM7Y2SaN2txVsU3/BHKzz4XD/OzVn6t7Ui
Hlxynmq97kn+7YlSJepL45mN5j+W2ozFo7fccDtuitTHToeghUATbwFB167aidKQ
MDBFrJ1klzUmgshKpcrzmLqV4HAmyd0vC0+u6cx8kV+ulv3+t+O0QWg1ZPgCuINx
JYbt0EY3JKc9leE5d0fA/I5+X5ICbAK+79i1vo0iCeI/vw6vY5WjCACgfb/yiusX
lIdx+GPvK8j1iEbcS0ZJ9ym5XsGT4ZOyc9KGa42fOqV48eJcYcNzqC0Kfip1ZSQV
gU94FZUu6rb5Em4gE85g/M3YmdgBrG7brCPM2Se8YGL/GqMedcvn9L/Y6dm6FAjc
VjtFefMLO9uUTZeIIhKTDOSn7IN5NZeOu2IYZDPVbIyk+VMzexHpD1uTEQ5BoTAx
Ov3LK+TY0Cd/8YKRi29W5FjAOywOkK4QTG9ZWEwhdja8v72GcWVUoDwLsjLYpW6g
mG2EIqXLiPrTg/1m/s46pBzyVdPjrVictsP5XQGgmK5Js2XSV0re1hvBli+b4tOw
UtlOepM3N3bddNKTtxsbfjwuQd7SNUsVwh9G9X/YByCkDe1lG6i+hm7P5QLBRmn6
POxvnL2DpKUEUJSHZ5+4q3D6FDwfQk3Uj1KCjWaVPLrDv5mE14BktrRxsV9U468a
KbzDqmSwBx1+/fSvpzS41LgRC/0qx1eaRsJdCC+Q115Dff5Ag15bzg7jWNvgryFj
5JB2A56dhJdd7a7TmHbkpZ+1BkHlSx/Ypc6KZC9lST2sTzsQbNHIsHWpykdbOhzm
/kM7I/rDzwLgzKG8fzfOjGbnfSRNP3FBeTtxfVxn/xXhVn++bBwjLLGJPtRjSYR8
jwil1m+M5eRjGjWny5IoFEHpryeOkYQiL8Ah2XAEKOAiUMsmlvURHknqSNUaeW27
/9gUAfAAg9Ns/Jdaj6u84Km/idyl2jYJ1kIXQn6hU19p/LhbMIC5MLUFKwzdtZcl
RNe3L7MJW45UfMVrU0sj4u7nHxq2pQUvsb75L6u5TFCas6KKAT5Qa/0pa4b5Y4Cn
QsfMi++XcZC2gk6WUPtkfxcqUR84fsRTcK3DpL7ZcumZel75wnSycCsHErs5GJ5b
rt1zVw4EhhmcEYbtrFD1DmI+n7KY7PT8WK2N0oHNWrKkGl3fxjWU/gIZnmLA7bpR
o/8cyZdPcdbOg1wOo07MGO/Beduquis9VDZB2KbECupIiBn9l5zjfv2bXSyaZpql
kVqIPb3lgW9tMDXND8ouYT1mTbLdU2AzN1U5tSJgqtDlwRp/4yTcLLmP7iso2lqc
wcLkyPaApfcD9Da1rFkRMlXZI7460eiGKNiDG4t+J54MOvTkauTqoaLgET0EXFcT
goHmUZWbVEIYx/AvdUkR389eny+JgDdWAjnuxedirqYOreRHTIk4aXPnTFp2mWbj
GGSq6s7vzIPTtiOtGWYhG0U0AHv9l5N9i+xB/GylJ236c37TJp0ZzKenJD9l4+Sl
AtFr2CvRfzz665SYrMPPpxj35FQ1PLa89Gz5Sq9iGOxY5yqiOXrwQL7asfsOC74q
H0LRRZJhXccLfh7s1O5c1WPwDhPy6g6YPm1WZddvxMgsz0WBh/Yb1YZq3c73ttGc
QLve57s+gD1dIKFvTQ3nogKX0GbgXTkqF95/jXkGNIvANELXBwQVfft4qyttzpoF
GxOAGRogRFBcw07/gO5RuIpmx7kgBA8OXWp8jc8ljnvEMyFIG6Zk+wIYIHJWQxA9
lpXmLloYABnKCC7LjHVE7qJa48JjQ0Wr76qauKEIK3DVS3BhMtHjXDDJvfDIgSrD
+USAQKG2dFNmeLgOz0Zg7FOPSySjh44S7W+fL3e77cXmZkGCIlpTy6zEdtmDlT6Q
zbEnUtrX5c2htUUeO3CdQMcpHX1vebgksNzdJ4fFrOAOFTXXG7mNnI3C/mZEN8m2
lJ0pPHJl/zgfVe2KufeoLy+unpIQbX9SDDbzdv/s+fxPkOnvGmIjxFg08vPKFzlG
a3HYejIjjoZoOCSUlMhSUrDncvEvZONtzOoar+24v4KkbYSUGh30K/Y4fNruZiVw
rJMqEgnHBsxFAcIpNfjY9oKc6Mb9/Q0PrEQrD3iIJU51gzrB2VFDTOAPbxa4/lB2
E7Jjy50TIrxVs0qfbmMI7PDViIusosOhf73JVpMMR5LefFtkawohgeF0V4v2X+cz
q2l5k/NEWIGlflj3ig0Chig9YG+/1/pWb9otWxSp16JF1KGhgKIKaFR66AJijGFc
yfd5D+0HBE5T4QhOjNbPDis6domgxD0vvUraA7QgZ+aN3R2T/j+BubmD/YWD7f19
TLDtWZ0Xw8zc0xKf40ve6Pp1pQqehmICGaXYmtBhuZwr+t6OqJ0j1b4klw2QQGjd
cb6QL3GwDOu4aWWQGCaBncz0yjJmVtCl9STy08O+Q/MDPmeb5sQuxlbzflxYH8oD
uUHHlCONsIw9BK/R7gxfKhH1rarOgXaoxdpBAPR3k7ydS/YLfwjV9vwnIkzsoxXj
Vv8CjXDzn8+wUQm29KIAdMFQIdqZmMMaBKz0dBomcxbfHn8eKvvQNXN4AepZT1Qk
v8hox+kHA8cJXkBunAbw+eTSPC5Gq1WSsNPkATjqfZdmFn8SkyNsKB8ZZ0BjuA38
McYyL6SvE+ZvLJn1L+RF4jc5RbeRPZ8K8B73oGAilOt59sBuC1DiLZ21Z7GWFckY
PuIJ5ymAdU3HP1xDRBw38ynavR29VdcNTZIpaMvCVjNvC93Y5H+2J60N1TrMkDn3
BfzCSuaPbx3ayOkpPzsY01+9ViPOI7OuMEr6owb7q9swRLmaKpnqtsLHy7VBCW7u
MjZavkbMI2JkmyPyOJEvFvJALFr+rQR1NBXq05ZyVEwQCy4X9x2VBmHNQ+2c4a82
NcZS4N643DzyoUPCY9VhfItHBp/cg+xf2JBPAps5HkHsFZaOpgIkQDyWzJNVDWdx
UMMtmjacM8cyWyDJBHS2yNF0HgS7iguNcJ+cdgusirTuYjOghHwsB8Rit0EO/efa
WdLSrTdQUcjX/QuT22JF03ad3ErarsE3nnH3xxc68fpbVd3MNyqUqMmQp5evttzR
k/efxRc5JZNszsyP1ZsKMrAh5fwQo7bw7Etvb2xWFNTlN5oz8Q85uyAN/Gels0ES
Guhmb+IXkTOzCmRuGIFEkw/qr/jm7x2R8lUkNSxSAXemPhGH9fEvFrZmkibxj8/K
zpxZKa9xJ+iWtWwvl8HShEfMlf/G+YM4WKldgfFW/1aDGz57lXwqYH9djFrDfW9A
lvGv8hW62qaKXBmYW8o0shG2uLsg4YHP9Dhr11M4coBPHmVXmfbm1EtulX509f82
NTyyp0XZHWjmFmdlPznbtAN3VHDZd5wQvCny7uiDmAEp/ijAA2YptL8MUL1QRWiz
D9ilY4FtYw3lSMWImMbeyzEJhTQexTERM6wMH0+6+9QZ5+1MOiRVIk4BERPyXlPy
66ev0ftZ2JAkLfFj+HWmuF19MPOdvHzcgVdW3woo8L7AH6Kd0iKHV/ZFEMruJp3b
fZExIUJcFDfh+FCqy19ElTtakgTRhGNl+x03gVHbZGTapnRfGfhpkvQ8oZgxu2c2
PyqIgmtGErm+2u4BF+RywGbO+LWdxfAbMv250XhlPZ4bihoxCXHa4Mur1GVSOr/L
40fUpLPZ4QXyzOMNFiX5D58Xkf5cgoPt1ayVkl7mOZbP6OmqNn6oljacmTC4mJSb
5ac2M4ISnTNf/ZJOkFNslfB9/9tNGPmmgDsmumeWipUklZ7diIMKcFsfvELytMYD
bHjV4YZURSEXO83O+r+++tJ/ZR5cCzg6Q6QSv0DzAbslreMfKGrpKSw8AELDJ6VX
NKQIrnQprW6oYokb/19G4p74hHQp5RePlRlaW0Mvco0yMapogYhMQYDj0IEoTnqq
fncUqH7uIqqMsyQ3+K6MT47i5IQeJHTop1JMVJVXjREsy/cLC/SSATkYg1RmPanV
0+0pMGLALKeLDkmm8n2MiLPagkUrULO/J8UbW3lXAflyibbEOpxWErbbEt6GITEw
0qrSmTIKZruiqW3c1Dmmq+g1dE04odbIzWrGTWLoexhn7OCeuPME5RJ5FmYuCEeX
sdAOX/NvelJHrLiL8CDpgHw1FQKy65lfdLnkL/xiM3oTKLmsBWcy+Mxzld1bd+nB
fxXqqRNRsUm2LRcyObKXlHd/yPqQeInOlxioLYzcOncojqe+GEu2cySZ1F2RM/QL
/U76Tltc8YyNQd5xeZWVGYcQgbZJIDpPhFcdfrrCZ3Bv/oHoxBvspFRJyU1Lm9QY
p7Msa36k1zUTv/y7tdI+ZpNlbgx4MNUHKcCN30Rm69zKUV0E2hoN5+RNE7jb3YcM
Y7GX1KlYkPbhoJ7AWE5BepNP/xa6YIZR1OO/fY01On4SQKZ82pO97CoF3w2pYTBX
7edh1Zld5ArgcAzpwmhqsEpXHEmN3Rk1MJjGB36/bD3yd/0lLuJasXxMacxkKCA1
+5bqdmVQ2ArHpbis5EjXZoBVE7lWyiRUEKQ/SGC0wpyHra8MbUpXO/GtUK4XRE2z
6MHq7R3MAzA2Br9lnZ2KaJP4uYdEOengJrlyt7nhRkbBJVen7WxtwbEr3hyN8eI3
OZec/TFKkmanfWhEP0k+OwjGRF/XvEB7oNDvhYe3AMLkuj1zleVqjsGerW6BNszf
qj01OpnIWClslsdVPdSWn/qiEcB2PKlKzUGNJ9HYMV7QYAPjvK4qRFvaVStq42NF
dZFQyQ+r4rQaIRbznvRU2p9Fq9ozhweC1lEK5rE+aPfoAFegtIv8NrCQjIXEHLWP
/rznTeNTgSdcPxM4bzG0tsTUkxKORnSWoP8GG5rIohzG8vR8xrVOtM89kQxPcLd1
gB3lMsRYnUXFaRAoIksHog1L66AjLh5U2haQkAHZRvqfFEePB30A2L+fq610wuaJ
xF65wkNdUCTnsOHXycZ0hFE3b/5UI17UqlkMIG78Fnw3v36QOvF6pt0UQXn7hyez
rn2lZHvG9S7qr7K1Hs4ybIWmpmz8ab5pPB4Jny0P104ZOfKNpj1SJ6+PCWliNQEY
1UXeDsXSIpowPOf5DHw0K9Gyb/EY5qkehP2psjhf1ibfDKL/zM8VsDJpF6iFjkYa
5D2pzc3GElaW0i86z0yBWrvE84S5ed0vvBeOZaq0CGT4kRdi18zMz46y33KHlp4i
VEzWtuPsb1q9e6F7Df9N/Niph2nf5x6yM03uYj/MT5yDZwHor3eNpEW6aRbzS5fj
pePIfvDJFMtFue9jxf0kmei9kh8zDHP3dANPNPL3crG1SOf5MAXG1H8Fn2hhTbNM
zy2k8QyiJhLWg8uI/FvtYGPMTog32NSebgjbRh9f1o5TMAmcllHABvFPOD4ZWOdO
Fzmtn6Ua3YpNgRwYhM9F4HHUZvWI1OdgXqW1mPlAos1z6HMwuTVzkSd8t5FHNeNH
oWpvVFNjBowBRxXVLBGkIMrstVxcRWco7tuhR1D78+Y07tUqBeUyIWZeHHxCTR7P
fjyhSg6Z3UHO756t1dK6Xf4PbTafbmpBJcnVfFz9lCEIOCm2Lxd9/T3yRpCssUr9
L/MBPuH07VW+kqsITN3Wr7s1EaSBRE3xBxjFMU9A+JdggwOy5fO0af3Dbs9s7jtY
ATUjPeD3ZQSKlqfzgDGnNy4gceFtJ4ElAKOn35dxFRh7TtxuHkhaWQW9nq+bXlYJ
/irKiOw4a93nTOYGiCis9s9YvkiQeDgAhgNM0Dsxx8i7jFZZ73YFxqCoKG86rJwE
OsyMkbjcTBQ/m+r1UZAeLu6oK+drhOlGyi/WyHIPzJcuQW5EpNVxMQJtv98dzYEs
7pAngMFZzhUq11x2AGu+o/IAAp72MMnT+3FIDazxRfxAayyTI+yI1qnNc+CIs4nN
74VxwCUvDOWBO2koYKfJeRJTwxX+jMKugJKV9UsmCVtGo3EmE96VCDar4EqSHdLI
FHx9tORJgemZhisLEWRNp6kaPemNKalvYdTxLbs8nE/3Op/FFocfEEKplJFsWCbq
unxvrv/f4m4pZxXWTGwlTwd56qWuo7I51Gl0z3O6VecdOdlRxSr+MR14qfzpW67e
QNkJTrYs5CcO2JBKM9FzmrAIV3E2iTLUpstoqYN+ibTEIDqY/b/PCaDtYpNl1c3Q
+Md/fox0i+X08VFYBpVlCADLvEKfLs835IpLQ9DJyhE1XP0M8C/Tr+C9qv1ne1t9
Cqh4FBl5qLrDkWSjw+RWKr3RPvqs8WOh+LMdmIUSrgIl810092nGn1HUMZaKrFX3
uPAWbTXZven9PabF82hHlYUBTEEwjJcv+xtamo43dl/4zjliRCLesEld2WF3jY9y
/HR/jSlUnSTMI4yeCI3PQjvGwK4v/I4VWq8/alS1s6zhePt31nAJdyDpNcLpAdMQ
YxE5PoiSXxn6RissuEiJvfoN1RMNnfpPdNVtLvKVGULORNxxVQnGIuV2KKrMId3I
fupUsT0RTeM99xog9K2P7WE0lHle/5hnYHxOBLsQHm4c34jrM/PXERIFpdu6he0K
tNvJyPD19fFLdnojMZkBGwwX0ctqHbKP+IBi4wXBAC9CdHdXbA0MiilZNb/2kLXh
HaeFUnndXE3wM6meS5E76xR/b77NvlRmMKRQFG0DkOoIVKWIqCJN3m1kANNB3wam
Oo4jz+GmqL+fh6z1Rc9lxwXkmbLHkbuDglP4SsAg4WoH865tcBljdZiMb5cyzlXy
0rhGGpScY4wJfPjQeU4vAJLoJk9ac/a4h0uNd90q4lKw/Bu34GerBibg4VZqTmkz
+KaZeNvYA2qljLzTTWqJk284j3nURs7ChCkrLB+BDsiPN/7d6LlomXfr0Dcw+Mlu
U1FEExMQ5/RlMNNzX64jE8Ko8TjAzBddUK9t9EqtngxZs97IgTGTkgKafRQJZeNz
jee+mWWN0JW98qNzDUkGDfdlYUP5+vEGBClZTb22KA6/K4XijsBtJSJJdkBJLnnv
QYkXntdHvCANkYRMwyN2A195iFx+/lEKdfuVww6MHxbEqTAtzFE/6khHiGmWJgTa
/gADs58Szibgn/TlJRrTf9Z5aGPbY6CVioax1KRiw/w7L66c2JW1Dkv9F7D8IUnM
5o9CEvEXP86ni64Mn6sxt79PH4CTvbJ7TvNqTBHY8PSq05dSlFugpMOJKV1hv/iX
pJ2xOBk8nE5M26ZwxzXFK7XxvJfrT4yQ0YB0GGEHMVlBkWWl4uXdCzoi+rXkZ1i4
dqg2cut9RMa6buo9yXzCZm+TKpwoo+kFtVanJI5JFqOEdjDISw8RW4zmX7wNcghR
ru4npWL449/Zres2TrcBqOyHo+OIKK4YP6Fhfgtceiaz44ykjmnq4eUfVqdYcIKH
BabIixmIE0SsI57NEqiBwx5MnRHFnHLQQpaZf6vBu0+/gBpz6i0ywuK6fhoV+FVm
cR1US/cNd61BTbg7z1k+7R+8tAn5ZudFa3MhQ4INCGcbGHSN6oXHjTalDShBBQO7
59n2UKsOPzS/qRq9EVmyUAGDhG190w0m8p4btLxu7jAj/UW2TY7PTHFcsZb044kU
uVK1GoWVRbS2S4HVqXbmxVbtsQkcxWC4BGFz+MKhKqKJQmVzVx5H2yx+4WCbBHn+
4lGBTOOD6BkTPJRFqC3Wyxl7HeGSDU5IpFFzjMP4W9hwFE5fhUdVfocQ0ZOzZCmt
q24uoIgH17w1cTvHEZ6psLsFnpoEwBBH04f0tRUSVYlKRRkPU7+rI/mzmhfrKoih
HGMQxtKa8l54lH8u1OYPXjlaZ7trHkL6nXsX6EvJudICVS/SvNzTOr54pLvxWWfS
Sp+C1dfAQhsboRMvboWn8/Te4bvRt9M7svtWftsIJhsxSLi/g/3JJyhTwZdTcUNe
OGvKmbv01GfS4zVQPpOMy6a9QnRMDd1fLxHmj/MqY7UCCLR0XM3ebZqOxTc8nCC9
LearMslJfjD0bLL2c+OxhdBS6HMyMoPayYzvEZjR+UREIoGiHkLoP440lgp2lrns
gW1ZGgEdsM0vxFW5weTibFyveAlDRSHkeBiFyKDoSq921dqaKDiymTuOP4MPzreM
1Ja8JmWc1t7bIrhVKHVEgAd0pOyP8aYQYwsTp0cIgB+gQo2StmrNClFfQe8QNl/l
fHjRa8zgIQC5FzTGdDoA5ExpKufwEX/ltxYzt/7AWmMfSvbTmBRwc7l0TImQjkc8
GKqNiPfe5QT2Onai1IADiwKTWzFLr+Bpx7/KOp+pP2xVT4nvA7xiePhJuwFDNg4j
z9r+QGV0yUBdyjZAJcpejDxryiAIte2soVGAXYQYZXK6Ldwth3c1mw8cPjgwe9sC
B6NcmAAS9UmOe0QH1p1wcQ/26WFNOWkhw9Bl2oTRrihCyVJS2X1lTJEbuNWzB/KT
ThrMSjzXxOZ5LW3xm7lZQM/kNU1AD4JCPErN/INoG1Sz/5peUCd2emesbII6614q
Y8Q4iZoQtj0+UA8zZALsbI6ykORrKlT99HXQzFRsXwSLRF8hPygaeTNKeHfva/yn
qVNkJQ2z51fRpMagyrjvjfwAq3R3rMXz7W6PCLpbwat9kB2bI25uojsp+OglPxG6
FLVahDHw6Q5qbkBFWO9j5dSZdV7kkNryTwat1nMlswYyzXjG6D3M2z0JsETTxxdm
DoCSLFNdXgUOWLTTcbsBK05+j5JPTy+Xh9cbk9B95DkHM2rMLBYUR5azKR/49Clp
i7urWhhupw09b4IRb3GqXygyMLOqitfgDSxEaSTjPpXaYJnR00RL+AswLr0vY49N
TGS/hyINwImamA+PajZfEpNVXAWNlwDuf2B7Q3SceL4OKHftGgaWUITXcZYbtdZw
jjk0cKE4iTXtvN4s17oHXRpuwdSYSQEO9acDEzLqYJcgf9OPGaOZBcyd/GPVjOzX
GILO6wKn4Pn28MRFxLxKf0ioUv+RL11Y9GlWUq6NZGk4Rf79ONL10+lvTuPopotX
zbRRYlC1xledf7VmJXiZKdSdRBksqAGaG4u/Qa97H01p/CjJVVgI2k/wsl9cDlCr
MTxAzrQ0STUHnHogjlFsQ9+RrZYflucXUoomcFmBREAexqXGOSUrWawg6Z3q2zEM
6A0EwaLAMcRC7iIwWJWmAZDhXgdYzaUcL8hoBrUH06XckmuW2ot34qAzu/hjyjwV
QKiNLfcQRQjbuDNapd19d9v7+2u1VlphDYAg0vfkrciVYo7H3G1mchxV7ctno1Ze
LFFhppU1YRRhbj7QNTFVToJVfKKmbklqN5w7gPIOi7+wC5nViPJuMmVZqwUJHDFh
q4xOUzBh4U9+KXlI/mL1DO6Q2HdHes4cBrXm8Tu9nNEc+u8CbYD/bpxExehS4M/I
j2npzruKG/Krq0dIYNx9E6dxMAS/gk/WbNEtspJ17jW2vhMCAMRdr/avDWhwHThg
GB2/p61UZsPwZz+v//+CjuYnQP2HG6RsgA1wB9rBdl1i/a/D6DLpz7bbFDErmB5+
PXqq1sMHnZC+ropPZzdJgn/ctqLb0dYrhgy8eVUnyvoKjn0T5Im9kdemOPyp452H
NcNA/FbtXVXTKeAzVqehSaDFRi+MmKdEe346+gL0jcHPu7CtZUB3raUNCffbr9+W
N/Jk1uFPozpmyHgdU+ahkvcvaWLAuymktdcHZWYh+KIlZUJ1EbiHeRTeq2/arfMz
++932AEkbeXceRuWzqGUgw3uzap1j6J/N4DguHGnSLlVdlfFO9p+C9LVt+bRp7yt
4wsT8QYjSusM1iiG6t8EYepFsP6diI0BP7tK1QWrQXb6dwFJQrrQzR/GxETm1pS2
mplGsqRxE2u+UrWpf1iEFYjkczs6e2FqM/MuzN4TdRp4/SrGbh17RxIE74w2wVhO
VCY2sCZ4VaMNPZHTy9O0KeDThILkgV75FeLrxS/snrLA9cA+30BKSMVGypwT2SbY
WvGfXvrGsQDUOIoXQ+6ZRAWqSGYBTfPAAVLQoWEgfYeXUrQH2BMnISUPmc4E/wjx
/v+WsoDxNkUBTbhS/BjaXvHUAFSZe6NvAD+hh0q5zHPBH2o7cowQf+aGg8rn0GZL
R/dn0YSwDbyDhieo18bJ5n9ViWXfJqO7tlURx9G0gCHb3YSBqnhB05ldxBGbT4SG
j2980Ka+bMKfYYyhR+JqaLYMY4K0EHtqFieWIZiMfQ11uix0d5Z9Y9/MPtuCn+qC
dahl0/9wsKtM+1hn+pFiMbVgaQw9o6QWfR/w84c1Gjxvf/im6Wyddj7FfbQPPOAq
RHOTV7vOTAX5PDoGLSwN14V3BhoY1nRXN4bJNF9kNTBFnn9Ek087ekbqQN0XjQeY
CabSpJp/2oV3/jW9GgtOuBFE7f2i/5vW8qlHIssI82W+YvZRr+Aie7VRIOsDmm52
RpVWNDSxpnRWAFZ4+QeG63kqCxsYfvvF0aO+7rHxrSapZYqd/b/GkxnKnu3jfFTX
/1f44ay5+y1GlbPZopidsghxx3+WUp8VddUe+3SURo/gSBqAjAjihRoX/VtGeyLI
hphx13WTYgzYPJVRj59LyM45OIen0bH0S2YVL+WEt9ru/Bfr05FZZIxydcdHyT0L
PIU6wAmbVTQpz/ViPBhtqqKDU9hd9Qam58j2a2AVbszrx004zT6CiXlpPdeX244J
F6QJtQbl1gyZWS9ms7Aw1hs4bPeK4H4DFnILZAcj3BxeoKjuq1wN1l8c9eOJJ0sm
mPRc1zNL4+7nviqEV2UyVf4a/wzBfpB6G2GIvz4A5gH/lUJFUzsQc472qSk1BtJG
4xWQYBYUrW1XYuAFXpnWPctaRJ1Kw4TcnO0z/scc3XAGsp+3yVaHauZggP7ypsJL
`protect END_PROTECTED
