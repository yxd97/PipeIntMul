`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uDhw5qulLiIGu73CLFHzvCRubOCgpEnXeTiTuxRtcdw76bNa5bNI9RgC1LVBLMmp
z+E9LWjjbowUpXVaN//a+wthkycEgddHJe9oVX7qcBSB8hveUVMMEFCchRfyO33o
KT9eK+worEJWUsAX3PsYpu1FneKk+KPEYIXDKQqjBxf4jyOB94lLiFCrqXEZyeX5
E1NphQMpUdlQnWwwdBKTdGbws3f0s7dmpBPVt4d9xNCNk7hniNcy6ahLODSdeFmS
gbaaTNsuByd7VP7boxek4M6ABUgxlykAE1aOKIQA0svTksF8pLgoyuj6e5TkZwH2
9ie/defT3oBQhcD+PfmsN41UDhDpNSHqVtmGh5yZ7BksPNBWTsQVZ/KMmtBSS6H/
sgwsnsTKXGYm+z7R25wMTmbHj73K3VoaoCmU+KUKsY8621wzK9h+rsFFB4fPILWl
Dsmm4E51dL4FPsaeBnGUfD9k1LWLwemq5j91RiQ6CW69EIDcnCnAm4gGcvvGDoJY
kKbUy6bDuEsDFn2Ac9F6kFEwR317mst7SSHRUAuCKpyfvJ27y8+/BI30GcjCf/uC
v8kjF1yHS+zCyy9u6yHyHvAL81Dh/6i+WmAV9TU6/n5Wx/C/TVAtV7mSAT7xrtTo
gU4lzKxd7Xzdr2nQpg0evTXVLUZDMfFV6HY2QW3g5dZciTdFP3dCN58cITa2jluz
55KQ8PriQL2SL6FPuC0OE4E95lCUU3x9CPHY/JTkME3JtlIBnnfDGJt+T4/n061N
WPTw10Jdh0PgSVzvm036k1ONJn7XwUQpw6flvywsLq5aOvhrX9AAQFmdQpIH+6C4
0ATWO89x07ULeAtLu/z/IV/ACmkSuS05SjgyB7AgD3CEFaXU4gsOpjTLUjgALPu7
V4pPAFgY2NCnTe2Ekr21vi/AzuryRJr/uJTel8TWiWAMRVBYCnlU8rlxuCsElQGd
IXRWsKC+iKs/1nDBDits9dg40xZoe0H/PafhLClblvwlxdhiCCSddLes7rOJ6hBK
K6FGbimW/w+idtq3X4W42TjNC7bab6rJ4tM4NiT5FRQK8cPVnbLrofpTUWVJjbbM
di4dT5Uij96cvspr12h5Jwnoi3oPYD7Vos/6kLYi9nygRTtZBlgtfRCBeSRjmMCK
NsxoNUyY+eUL87c0Bzln7Bo/XxTarDSUbLk5hhur6Kki1SCMZnpWEudqjfJ7LN/A
mIlXceWgiHbsJqFC8xwzOaG+3WwccEGmekW9TZWo2ytkRUP854e8XFNBVO9czQyY
VrARC6Q1lhEHmFfjPcZpQrixQBepchXddJX66gCFaisVZiog5+QWTFeU129VH9Th
kzu87sseM6if7fINqOpYcjWmsS53zNyhfgfbJrOum/PTwngYzYLuBbfNXYeOwVts
bx3dJkkhmpLNCrZZmuaIUgOJuE/wPHWd7WfUGfmBEhMUZ+Oq5tz6X5xWKKtFu6Sf
FXobI4tFVevkJaCYUUS8LAtbAds3tsAND5LkUuICOklXQwJHB7i7JHrEFqx5eJlN
0mCwmiqixZn0fMeMJdhLpIS5SkD+9BTI1YprpHclgm8ASJLETKZ4mwmjSQ7iUphU
2fw6Id5XFJKORgW+ukD5tm0CjqUsk8dxrcva+z0SuRJ92WRHPqmDFM6hjcF6ZtFn
3v/CnDm3jd+0hMegkQpDn39zPz6f5ThmyyU3XP63WGaLZ3YaAo0B4mAGlyveDfMZ
gRD4U0bt/LneFy5IqWn0FFiK2hcgZvbfkcqmnZ0sv9T0oJS+rgNbtpxS1B1/PxWr
8HJI2iYi6F3VKlLXu/RPrFH0dQQWR4wZOynPTBWpePYbqoD/gW7owyIETqT+T0+3
fuN5kViQxpENg35l3nWxG0oO97HCVTPUe8ZPNfhm9ho=
`protect END_PROTECTED
