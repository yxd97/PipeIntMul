`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ACH6rTdf06WYgyr+/Ho5wZsvdrLphOUN5Gl6rVBEVf2tMiKS8yr0XgbKewYiAckW
twZimC2eYDvMAJyBI2sgXO93WYiM7L573JrYMk8RmTRVSgjV0mziA8ET3EFN6Qcf
hLZJn6XOrPv9n2yftW18nw86JYLVO2OpF9a0SQ87KRl6X2Itd5kY8xp424Zb9++p
HRQAXZ90GIZulg5+rCaEopTqcWvU0NChsmJlbbISfIWdI9IMB1JhSoPxHVZDW8qs
TBt5CVFc4MnHEwv2H+L7LaLLAQwKe8B4wR47iBX6lZL+XR6fiufl1sg111QhMx85
1sJJbTYmJH2dLBV3rMXeeChtLYJ8oQl9pXE6avMLdbfs6ncLtn1C3L56hTU7zG/0
8vZFfrL+zL3pE88gwXl12BVWc+mfXwWo3K3CD6k4gUDnP+C6cJ3h//lOSxSKUyF3
GVuuC+AZHRm+bW0yQsYpb/fS3vF+u9lK1x9jQ9kbs9A=
`protect END_PROTECTED
