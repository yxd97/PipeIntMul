`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ivTD0wgHqtpjES4Rbs3g/dFw1FrUyLgOxCSucea60NjSTHrDxp12jIdTOE9EGcdL
xKk7KR06SM4GBS4swzE2rvNnXLwWymUgK9dEwIEfkaMKmcK06rqN/iEHVXm4lZIr
Ab34S0fsFr/7Nfqe9xHFpvGJ6IPmBiZbGediF1CB+YI1EGaYmkknCUNx050N9Rks
b2sM+fLWvkbIYZ0FtxlpjclqtskdaPk2xywUfCa5BE6GMy98IMdJye+PTDKYsIMg
BQHiyrSwzv6v8Pq7KhZI+nNsFpZG404gsp+AraY4WmdxV4xwqmpDSerqNRtWc930
9RqkQ5ivRf4sthUDeZ7WO5UpmcpC7jfop13UsWeGqeSF2opJennuesqT0LOE4Z+w
9YkTLQangUUBawCXDF+GhiT8rFuCbA/Oq2/+/+Q8hi4sOYYZ6lGUOeJK5J8gD7uk
`protect END_PROTECTED
