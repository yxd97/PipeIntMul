`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFxoX2HJvIeHMTldfUIpCpIe+eisRDeQxG9CsKWNKFW8+RVdDw4Gpz2WKDsMav9G
lIjF/Szrha96/cNEXs9ctgMRk4jOpiGXz4ol8/7+hbG7i+6aiDqNul9we+7oRjbi
tppQ0YjY3GB/O92xbZk05ME0iym7u4GpdwksKnSwG9CTApnob/o7Opv4YU/8nQ1Z
R0qIedr1M+swSjYyG0bFg9aMqJ9UVKaLUAjkHHJByaKqszuVTwhdV2djYTkGvtyg
ro7IgjXGDVi6f1GZIZ7JHR4HJuoJ8er2xDtMWGTCDAIp7TjUa4RRz+GIX6tNpTxx
4m/6G9XnQZNoupzoWTRr+JwzEG9ev6AHpfKe4CjcssfKQTRa+FQmqMAwyFhZ9IV1
uSccJWfLKaMyn7O1jyksMcH55cnlQtgv5AYa/vBctw9jFUtJ4cfziNvnQuedNgKI
nElj/zpVU3J+9GlTVRvUTlclhCdAocUHnczzQM+dEkARKyvfA374fAeIjrnyZPlm
EDQR6K0m5qm2NLttaOWWp8sIETngMF3Im35gfXksjT3rluVIK9xpIM0/m7lAQXod
`protect END_PROTECTED
