`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nKlkIxS3XBDuM59vcZuucOiDDfPSQfgj9s+LtMhhTwag0yYMWAGwnGuZ7x11TQS8
F4lU7jA505hg7XiYMakbW97kvt5qKqXwvv8S4pt91e34IiD27Un/vb/u3xLuqAYi
4+BZunR9ZhiN4PhKCfup6n4mwhzMsLIaBzl4fURI9Y5JJXT7xuCR7j7i1/sqHdXh
yVn8A+S2F7qtLDUXd+eVnMq3rA8uuGV83y2TUVkWP73WwhPPZZeBn6CRTUJhirau
4/OOtw7LiTR/i2GVuAwEZcx3F7X0bm8YIOoq3C60kKQSmX+hRhODg77/uf7B3wvN
AjLQE2ASHY2UxN7I4d2SFoAc8ZMe2tlaJ89byx2xQxeqY4Qywdg8qzByXUsafSnv
yC0tFikXvmsjvatTy+ksrg==
`protect END_PROTECTED
