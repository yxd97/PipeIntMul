`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C8URQay8HSvmnzB+S2Yp8kajWSTTUHSSMZEuvOEocoazKOOBwNkz2faLMbsRN082
qIn9OwYYMeiTWemNYgNcAK+3mECWJWHDOTo4r/HXmng2IiGr1AJmp2ZgKM00E9Kc
wLvDNjLQiJSMZyXdVZHbUy1Yf95TF6MJRK+YbJgVBqlmVQX1rY8UQwNGEuFqCaZA
lKVDOMy7MmCbLKV4sCfEqlstF6/wG/YVeRMfhVGnCYkq8497rozOt6Idy7h8bh2g
y6OjjAEYBgM9uxMqByZougH+K5PRVpKNa3GfwnlKHtctmgxX+L9M4FTN/cysvOn2
Y6tyR64OnGexZ9X3x17mtZT8435hDLe7tMxuIUeMCaLPYat8q0yKHRsUv8OWnzKY
Rjhm4vRfGPpVxy119nC34LYPpyON/re07jN5tAUM7XnHVg1LkOZg0lNry2ToNoyX
4+vlGqftJmkfb/nnic0lkYgXLSP+nThYB1DVF1Yj0cYvmxn2ojdeOZuADan0eQCg
NUKVNkdMk/Odjes0swXqJqwIKxmDgF3OCnlQt/8xmfC1eMuon81SMzyaB+bO+h5p
7OvtxBAD9N1/9KskXNANQ3A3z489q8Gx3qX3sIbBj+eEqT5+GGq3bcw5M+dC1T2s
5MXZu+0dE9AYOChUZ7WBQiCEI5cTlHKjipJOtCSSmMxKdT0wQjT/HHQp9M333jUQ
+z156dlQS67S6+adegt2YzP5joEEHXbRiYcquVmfsgD+jy5KxdK4SO1p+3yf9Z3V
cAlBfaIDhfH9W97lpBbQQXquVvrLKNJOUjZpWygQv38E4b9JLGFuTPliey/RGINJ
k2CSiAGs2jg5YT7c3j1lJ+1g4E4A1T4R+U0PCd963hbYEjJgBmAbQuTWv+Qa9AOu
CNjRitBMB/m6wQ/xkCsX74BsQU/ndAAzcxsVNOFLZOV5z6nJznk4M4FC3WtjWjvY
jeOX5sL/4yCFlwe6fjvmVrG0nTOq4lrB94Yom7arwncLAsAQ3rjqjmenMWEObWKz
MPOIdzgQfa2pr2iPx+AW/WTss1As3IR0EWeyv+eiygWhrjxC1RR7MrUjyhrdoiL+
GoMN6/pYEohuEGek+RKL6XuT2x0raK/6Tf/v+hDqargrEo/U/4CKWxCXum2/2PzN
VVAYFuA9Po1WdYXRiqMvJL6uv3G+zXvN2n3KzJq+IDVf1v9z5HLNaqNYmFVn93Rh
buHMCqCuPPF+/WXYwdmKFWrUMEb4UzoWTjspE9CeoGEbtFWh5ej40DX//mJbrb9G
8QIyvLENWpuWUjTMAANHsfJ2sN+p8YbsL+h5XIa7TFHAseKtu5pGE8oOc4n4ooCF
3A5g7JFdFEcwLbM/n/BZ+jAK6yIsFcd3EN5xqX21VhQDTZzFd8n4BYqZzseQM+mV
iiceQJkZR0eAhMG8Cc35Q4rzPkDs+HNVw5xsUbDJ7B2F3M6GUydDmirxaEDjeErz
zMkR3H8IaR2oeNg/Bx9kRbQu8E32Ety/1hfm2PCxTQ5v6mMoM9yaFurWpNNtuEsT
EPWi8ipioJSW7VnT9fTL/shitjcxr8NSVuGukvYyrQCT1AdtaI62FFjPR1NPKO8A
TDEjYVcP+rSx3//zWSxVWp3379z1UtrFru6wwRyMjrABUeHA+mOSmY0TlmPXq+Pi
ZjfoFQf4slye/UJDALdfBsJqDZuGE/n/et9sdneciCL32dOGuQcDjCA3OrPcu9IU
fgBW4xzeOU4/6r2b8/JxYlQar6/9ubE+e5jUrMk4cV/AGZJCNCpBDT6PMflipiYE
KFavfT3iHL3nF2lVnSfMgbU4YbjIYhufy7N10g8d4pYOYN5dP94fSsKkIb/VMwQm
KqK3XBw8xK+hUYk9YG55vpmIf4uZp37RVNz10ZluJkTiSOQq5l/4/OwQZz5QJ2Kz
EWQ37Alv+tx61ygIvKzQOgulnpslRv7OrqcA2b1ah59kZwxvDwUbeW24ozkdYQuQ
J8azCiG9To85mPLugp2/xW5KQ/JMy7VnThnAZXUw3yxRFoHtJpvWytz0s24BybAq
j2ggAqPLV0K4I1Z6iRuaJvwQHNM0cGWejdhWCHup0Use+plfDtYuiL8M0Lhkx+NM
WJxf65mFreI/YOppIToIjtLaC6aGvlNF6+KVAS6HKdGI7gkjHmcJGl8V+HeJTfvH
WCBh1LqSbKAp5+zGkM7Obrc32lTT4bhk0u741QHiC5A05SKu621V5Ktmd5PEG+9q
Z8lMqnsjj3ChEI7w6bqC+OAQyWmgoCvCwCd8bS6T+mzYlTSQm+9Lony5Wekd5r60
LgVZOxvzlWugrY8yDqLshHPRGH/Hwg/8/0eushxyVJV3+qXx4mZ6IX2K2nzFO1zi
TKhV7D58FpYeJTs5957Byb1BUYT6nYOyonrlwAJq82o712QaIVS7WOaiu3nRVBPr
k+E+efXHUrcKe8zHoBM444XjEia5jUjMW6D1nKcpDxUGvKnM5DmsY9a2/Z+aUSyh
tpAYnOljutevxjukH7O/DEmYegRkqqxCfCbHnjzBEA0mlZdqJp+JCwlKdy8l3Uei
AFkFrO5Ulnucvshq7bpjyuGiS5KD4K7AZrRpPDYOOaiOld0O0MAeu7DPUk4HMfnV
pFtZYANlPO8GW8hLKeZJtnoOq49ylmVMmxVz+RA5ZblxT3sy7vOXb+Qnkm4k4BI2
Zx2ARFSJvXI3bggz82jHnuBUHtFsyUgaFPOQ6gyq28Cy5LMBQnNQ8wx/yogsK0Tw
deo7pJkjWnBzWL06IENnV6ae8UnVF/c9FpPwlw9j20o/nN2po84+bfL8Z1Yrd+rB
aBBoz5WCqCacuNpevQrF/snpdXtSXJgNJRtBlwdGcZe2VUXw98rQv8jTRCgArbMG
niz9cKFFed1FRF2gNqZsZHXkl19i5E7qZU2JGppEQBQUb9PmhAbMNEe0zsnMxA/b
Jlv3KHAd7ZKHJmf7LxGMw4ey//LqXV0EvAgCt0BXIMPZtkws+xvfGn3SaMvQSdM2
vU7vTvR7rntaJpjqWSluOwAgv8WXigAQGLYRrNfcqjGHGdRLNt60ap+VYR3PU3n0
IWrH58BtqksnqeWl6M0SXzbTtCUthU82RYaVZRJ/I299a7a28309WCr3TUn3iDEI
QSReGA/owRZaiuDqK6VDzBm/WCa/y13nAkR0xgCQYsRn4aer5zBWvsRkyh75FBkN
8y9KxvGj+eKreSqxdqN+I2/RBywvKmBm7F28oko7Hnt3wqmo9WD+gv+fKPz5cNAk
UEtwsfsrU3Y4Ga9E9/21feWeCjAfxkrqQMRI7wf5HCiUtgxWCb64wufB/JpWnh8/
/7zex435YtppOV8zniVA+o5WNiqtp+WpDdIsQ/xeeeroCuvUTnG6YAYuhHvVjMaa
M1oVYPihLfRQ/jnXIxyBQK6bTfChHMMt95Qx/E1n9VONjBOSDEpjt/Tx/a17kShP
r6OEx8htLKoq4es7IWsJ3IZUFuwdLqljYrHjuDgatKLoTbwkfrfw/P+NJ+7AxB5w
Q4a5KDCQultqyjunMKNnmaKUz4SQhO6Ze3SP9zg3MxdYiotY71cUVmW3M4itaWZg
rZkbTG0964QB1rQxx2MoQLrB+wV8s+HiRlnCt6glTHolRtwvj7C0PoUi5NBRrhMS
0tvsf0OPn9DGfy/1ESXerVzut++n9s9WG9k2jRZE58B5YPHyx4I8wtOFcaoAGHZV
8q4xvHIySNtRHq79QTzbtUgM8d5g8MrDlu3qI1NoeUcQbgQgbR+MZRxqD2R3TM9a
IpDCxl3Ng1GRy3eTaWKgbJCGwYzfXtfRq040SokjUIWAdPloEjGDM1P0HvAD6nQO
CoiAqYZzPQULSQL565u8GeEdluEN1AYEQgm7Un/5TKPSMZ5GoTOPY1HVo6Sngpdx
eMDGt0kLxZQJVQNXTS3LRUx5uPPZKN5CpL6UOFHkOyBnTgnSJYSbt3OGHFbNtCLw
MtPDikRY0t6oS/jca527lIIAswJykVHEwGhJijshrTyLV5uwIw6yiZ9jCqBNcF3j
arTWrG/FVfr1Sf+hYTQmm3YI9aQdgp1UoCNmKEEwX0oPw9ThqL8MVsxwo3PHxnN5
nIuEGvtJNxODg/+FbR1S+hL/QDpBDqk2kMeRxcsdaG1uCvZb/7chPjb1VMX+Y3dh
ZtvudZuWbEsIBRaxxq7I/Ht15eTXLtCsRRW57RVkPkUTSTETZcj2/Lta5OF21V1Y
MjsB+rLvAQjJTz4ZtdZQwW0wkGaUCFedoZ248+mq9cFGUV6B54dxwoQ5KzJVNQJm
FvViEMHLx3+uHVo9gOuy9FufyNfbLGoiZ8o6/Dt/MS9tzLAHxcwkmQv3cLzPETlt
13Cq9m3rR/cTH/33A4kJs5u8FiqiC8pNHUjBU3IWlPmPhXVeu/Ef7ipX/nmOiOaI
t4rr45gGhnItj3MR57KX3Q34nwxxhyHrNIaHJDyVK+gp43kVsvLLUW/KNWhhIFQH
xnDF8OKxkJgI3BzAK54KCUbcwRXrnxoYz3Q9Wt0BVOye2cC8UMWEAn/QMumgSu5E
ra1wTY9advP8PEwdieav1BqJkBv3tOEedn3gM1s/GZwDvAIst6UZwqQ6v7apb6W1
vgcsig1e7hCLU67Sv/dG7ZGVXtuj/xycvjRo+rBWAowie0Xf+FyDqTkzaLHnYTNN
94e0p11RyXHu376ei7FSNi5vRECfGXbZyoaWEMyD8JYlndRdUQHe6G1M7c87NL/7
HW4Hhe5w8811zkutsLjMqaFb6MkI7b56KKMdoQHGGgoReTj/j1KHowUwl/p+WEPR
3Q+gVBl93rHabgqcjB8vjahaZxfxMjnPBxRAgm5Ja7T6c7C8vL6xmcXvdFJ0cGdc
YDx73YERRvLj4ghn/jODf3MlMYq8c8QJGGHTXSQuFRE0l6bps4x3eNxRKnLk74qq
yH1AqOmGEKJdg7sHz5qlHeOBIxohLJb4RmjUP7Z/bdLfgR4/kMc84nE4PIX9e3G0
7+RYcCohqRjD7E9yUO+vbVOgXsZ2vqQqDfXw/sPpaqaD1VZF1segJmXRyi2OiXEZ
B4fkQWWBiyetg86Yn9UWeK5j2Z2PHVRG91AgjM9snUbqP7X3il2EBiyOmh5oqDnl
OwruudgumaFhQ+TfETR0VrndneT89ZpfcysN+Es84Ot2d6NL/Kpz1s7Zk6qpPr31
HXSAjrj/QVtcGYnnb920ih/IgLI1fzV1J/WrvYkTXS39rgcqqLwBVNDtwrmh72PD
2uuG4A9yl5JyRep9D6j1zJkDhm2J57PsNhUE+8ZqN4iB2Hc6KGGdkFRfD2l6Z9kg
SfEuJwobHgmLe1fLZa8guLOfCRe30Qiglr570aZmMyJGUsuJHE7+wd41lw27oakt
rsqjy4YcRi2oplchxVZS6s+ZYN+PMov0+mUBN1XGCnl/qutTK3cD/78GMHk1uzCX
TaDNyypzvqpJXf3iflQHsyd6eU8R1ZRs5r2WmhgEbbZQsaCAtmqLaY4KP+A/NhTd
/jpSiS3QfD+Eu8/iJGDxLxBkKFFTMIcZhSKUrNC9jBb4B0qx82un6Tj57ygKngZC
GqKaQshA0EhiXolvdjH9T9oIE/dSETE4VXmnWw0l7JrtTEqfoRGzQkO5aW6MmlzA
Zkp6eXDCwY8S584456QddmMLEL/jp5Ua06KmPqd9+blsYpWqWldcNJ/4kMHsf22D
3H49yJ/bLWm9b1X6zmh0S7GXbOWHL8UYt6x6NfPCUDhOyqzhXfEpBYEz+uGuNSFK
0cxj2gdFjqW+C78z9XUXbt2+c4e93kfU4HiUYqUF3OeFOqX/SMQw2kWpjythBHn2
19Ta7LMdETbu0ae59EBrtjnoeztiIWLqU05agkmyexXXZTb87araRjpOn07kzFPd
xqGInMPYgusgoe0EjFhab83ucxsf+o8C6XExtS3xOueZb3+YnrW5v+MhOAEqmiqk
5GCThxJhGbZyAtemGf07IztNBUa/LiZfmZZFrXwM5KNe7H2ys+Y4PEc9J5Hw8AvN
EutbuyK+9kNk/mzpOzaWM1f9MxitE33q1RzbkIExgQ7BUSxfXqE5cCjTTUgdxrZ7
fSumyRuaUQNuG338UHKE3kbCjRbKtRM58PbCw0Drt31P/rqpFpoS1h1lVO7um+nS
Yo1AitjB8OEr4rr/+RD8cNoGzY0zES9KazXmeh3hyDoGj5nC7+hF4Jwbuo2zjYTw
LL9vYd1t/40AtkQBIatg9OkRuQj2e6vZxb4TI9G7+kPmvWDK0Lsju5XCPWtColaq
hn+0YJRAXR8MKo8GNlT+2V8hzSAoGfrUzrWuvHG/EZePwbbNsIOUKVinIoIM+Z9k
3vidXjY6qlJ1Dzn0pdPt6/kL9/FKtQAB0mU4UexyM30s6ehoa8LXunpcfOPmlmzm
J8YFnlLU5EXj3Oe4HAky8yhiJhZ8A1Zio/1GWhrXeR4fsFXZUC2kmrBL4JZSsthi
30ROyWk3OgjhvYIlq35phvukYkvkNjJ6oMVgqn85SkHZUH98iYGfWTrgOEvigeSA
2M1bTv7NogBmbhCTu0KaPfpL0lmIGKh6KLzbktwEMwGFJpqdgIh8KF/1CdysRLtp
UNRED5Dds9/qwQ0g0iuUbpOXc1p7UCoQqRSL8UdFd7ZNEdTnz2KvnL7gbKoSIpnJ
gBz0ere4TQCzjN3N8f+A8Revz6BbxUo625LGpYF0weF7Klod0YfHm7OyfagZAC5v
KX2sf0kjCrTs27BR4+R/NnwLeNZg934CRNZb/i4oPKDzgUbcpv8x++M1Bs9wGVLF
xOUgbKHjAHbWAGmALFa/iPiKoCOJFz28BTzo8i0YwCLq4ukS6gjFASAjcwmTKJ1O
M5mne/yHz3VNWsUD+hld6+zfCiU6gx1vFCwJMmSUJYwscYwm8uk6yX3f4pdFt4v+
4tBHrAwHMfNRNu/HXtoIyQiyhDRLdp4+Yd68t7eCuWOQL7Mxob98O09/63houHh6
QUJyJRTJuJ0lkZ9X0oOwauTS/b3InXGfR0lvf9RF0aFMXCP+3ZfufplB4pLvby4T
RsrKYOe+ejTQwO6LrMk+I9+2wsLlikDz+qtStax+LW3jAVv4e11m+tRB5ikrugmT
9Hhh/+qdxmuqa7UaIyrTJ2woiPxrhao8wIQlZolGdpo+OYSUfflMGQwKhAZku6Bo
qyTEJ7i7uj57xFeyyJdbypqSgjAG5hTg8ZxWVk382Cg5WZTBAAePSD0VLHA6LUH0
tIAc3eb1go833O9jZu8h4kB7JNTpW3GiNSAsKwsqhev+DqVK68bPC0Z8YDldnaUj
oNgQDVJUaee0qo0/baFCzUVhBPYNWiSDhvFcW5yFH9bk7cz505JAh/RXJPsOkjbW
wr6JhPiYpJ1rJ1IT0R2BHVElYY8+cPZe8CCyEIpkf9zsXU9Y1CC6YykVr5VcZ+fo
eAdDWo0pWliife80jk0llNAWCZtWc0JjfzPnuf6KWM3Rx979ZHjMrl8bL1AwQzIz
QNEN3KpU28bMbfPSc0591CSYVb2tRhPiQoAgOHDm79oG5vbGhS4FiDIN+7kbo6x+
k3dEZ5nw323VqDdlZUQWDWBzeeSQEmhnFySoTWifA0S9jjayd976aXbESGoE1BVb
FvxARdCgyo0Sryk2WEUmd/aiaBJ5AUqrJ7Fj9X507hdDUKgrV3pLmhaG7zco5HGq
prXUB4hMtsPnhXbQUxV5/yiuAd8Yo7iVt6MRblTv2N8buk7JGELpQFOaWoJkqdVS
uBkpSz+FOk+Fvs6RIl6Nrg42ssPGCjZ7WVnKq+4+bgRFhEawYZZHBrMmu8/gf8rU
gj99wGElx0yon1ZEAOlC5SBdkVxy5ff/nt48GTu11HKjfPwgYSRih1GWuwbQw6rd
rJUZlBgl71f5juCeXL75L6FNzmsSJfdxgQli0VJ1sbNcBFUShaEBy7pS0HWp76Zb
FOcDeYqGGRjtb3IgcWQIM5k4DWIluj1OvmhH5080HyIisd5LQIW5Usl2riu3WI1V
HyV/yClKcVtVpo/P8N1Atc+23iq7v2I3T7GSGd/p0tYskhIgii4UwzbD8WCh/kfr
zYPMTQEHewFgWJFDdGaNIqSZTTH5sjXz51MSZTRaXC1D55C4unGzPkhNOGFQAS9g
urLqPHM4sGp1xOCowBkfYCWCUFLAJZU3AlTcqBShAjKHL5HEP32TalP+hQ1nW+Vb
o584iG3RdU1Un2zf/rB/FJTovJbTTxWcRTD+69rBNu9JzkweM1nxti2C2CwEbHHx
S74n6qQDVQqf5IOxR9fg7uy87NIykGT4o5+c4cNSS0vcD3ziFg0QCGOwxDOD3y6W
SuSaDVc0ABQ7ViG2Zva+B7Bh5WtECLSHPTy9b0INbuHuuoF6S1YmwxeL/btA3Cn/
qSJkSmzfnjJJqs65W7ZJIGbZ7gO76aqlUlTsychkCtrC3S7Zt881pQC59FR4PW9e
YBUZklq41bcLK/p36dt6T4fajvVc155qdcQ/iq+GEljQ0+qLY2ooxy5rMyCbkSTN
6wOO8PUj6HPKbg82jv4Og4BY8lGV81rDMHvGFoFDKHLpaJKWxam3NIIfHOIkxWfH
V8wQN3wz1yn8YME0XFnbtoAq16uIRA2V6VtbnE+s7EWylI3mXK26zzLqjCM0oPG/
Ad/xrHFG/KiZ5gQ5+Ro3drqZkUr/jA3fma1w54nZV6FXibFdlB4Pk0dUO1el+BeE
QHOdQmKp3I93fx91UMkZLT3NvH+afWnxtcTNbZs2mb7vp50Ks03guE9gXhzIBl5s
lNlNd7T9wRCtVOzZVjm5KMluV7cgqlLs0GEDU/Q7fatFQwLsURjNfxcW+zJSlBbd
Hc5ogJcTEHXeym8ISINKatdk8wXGaCEis4ch+Vck4iCYJRkXaRvqN2coiM5FOBxI
Wijd7/vPemPc5dOZsvukpEOtrSx28mcu1Pmx9ydrNxidwf/uErVVovKJsvLcUr5j
mWO0z7GRLoTtDs2ltVZMKEI8QzSyk2FsBpW9YXMWW2iRN7RRusDjPFwN+V7d38St
hUtBaCTOE9g2T7WeHhm/qZ8Ep90/8EyISdG4RF1U0QoPvwEvmShcDtC4Um5EVWGE
iGAGZf57W6nTF+HKc0SG/xISfkg4krQH8P0mOzZogSxzHL0c3qKD/IDRDu+sB7th
qMwXmfXLFFs0erJqqoTDvHMaav+J9vEoE0CuQ2bpKtOcr9EVcCCQhJMlOk8v9swr
uCm0RU0yjXqahP7Pp1ZxLAQgMnahmPWDfBjOk+DH3zfwJAyP+LPG+Zop6tRPVQ6A
6g2esqvOSxEfcF3WWE2aRBYTFTwouxo5P2wo9AWtKZtpAN6RAHSR6TlgRC40mzSV
LtBVgi8iTf6QUk3s96lQdxipv4oFXSfxzzU0KaCfyiQtYeKDNeSCwHue7C49mNiQ
qH1aRXfrZvev9ZYiy1XoPvSfKm1rhrDNC7YQSqWeH+DAeNJHNqYwPrcBvHig96aj
wRzA3ZW4kW25a99Lcw9EHeIZtd3+h1ZftmVhlp8SExDgdg4aiogrELXrf1UpiKay
IEc3KoctALkNd86Np4AQLfM6wsSDaGtSdrjj82BaV6apdVPfUOAr5eBRqGV7U1s0
l9Fs3yWmT7ldJRkP/+bWKwFFuCFWvJnFPSN2LyOJ7Jot8nFlxpRv88q8iDM3CoS3
7nWV+dWlKZCUA16fhP+nbE0JB0vU4CHV8AyKo0cHDj57dbkx0JRa/s/XJdytKyKm
+KFAHEDQ9cJwuHfwmFpW55M/hkGMs8Fm8aVJZNtS4rxQ72pFMialthKOxNF94SCD
/AuBxBlCmjb76gSxbGyU139wQ8tB38TWMLr7ibqwHJER9KcmHRwub4cC9JW5Wp88
tpXG8vv80GjxCTmJ5QR6elHp0kqcTFv/7HWnK3Ry5sg=
`protect END_PROTECTED
