`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Vpq8IuV/CjMUQhX7+CfIysNU5/3JztDUkUfRtqR3uIzKlGx2L+A9ucBqWFVw/WX
xQ0qiIiQ1PLgAdWsnMC6JXhps43bpEwWMhWSyP1jodeswAp5nb1SgERJfeEvcFwG
pMK27r8+qfRjgFFF3hSMLKDgV/BxvzohD/l3HqFt4QdnDA2sYNHkAmJV+nGXZLpl
8OHmCOl6TRs8CrcR1+BBQ7jAMCaDLWboFFTA005S11XkGmVZnCmMrK3mQTlTjLD2
fC2ssS3xoWTL8ltKJBYQTGQyKUhiBcQxgcx0S9620FNGr/eyxNYu1ejeu4rCFPX2
9FvbOeeS2OFNTLUELLd0Uw==
`protect END_PROTECTED
