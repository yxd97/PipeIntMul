`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L3bosPtE1vR/i1ASemI+zAVx0cieNQfwZR3NXJRFoq+mOhWU6kCExDg2ma1iB4pL
ml31E0BYO5JNhTzN77G7ZbLxlcoS/+tYJ2goKuff9/bZZSg8JZB/e7yLsxmYccTY
GuhBD+PJ9NjxvTSJZwhOLFtcgKnkr9ccY8RmWPVC/OUGNCmhv16ZX4HRtLj1CegM
loI0lQboDdC7Xw6N2RLTVgoXlrteCI05GB1swxRLL6pqF3UnJphDwjkbroYACZ7r
ffCKY67qa+R4j3CakeXo+g==
`protect END_PROTECTED
