`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/E0ehKilxN7qLQBljzo1OtNc7N30S6ZE/iUc+vBgoiQi8ihLzBkenl2tSBVzgFc
iXNJ4VAAgXONhMtTJLFaPI8kmVirJ34KH0HW81kjKRuAx4+nYzYoTq9UWp6YAG5e
8wXlY8l4dlxrOi1KbD+UDcLX8ULgAfyHeoytOq1dQG/vWitqGYa/jkTxMwutHhEA
FXrL4pyUHYRzlyQKx4NwXTjx897uNYxro5M7w0yVXiTKodaqgq8VWxAKeArqKO8b
eQ1yCv/T6iqDzgU0ErtOC5lWTJyq8vSdL2o3AvN/9cspH4nFZF6y5FTsNIDsiNFq
hJ3UBZdswEiPu84emBTr0ZZDaqOrI88++8UtV+fn9CxfFExekpR3KSClazrbJU3R
3bHvzoVkcsjeg2pdmAyE9lICeoZTZUIi+P7GtfZy5TQijEyC2DU5txJXLy5Ula8H
4fMyNhLtXSG6gMBXdqPozKJcj7QYLWlFZPTiY+N8a1qM22qjcXvuKzuDpU0xd6OR
I/R7LTwCYwq7RSKPnuD8030pK4o/uuUcgHs+w0VNkNqObewE98w6X+wE1pvra1u6
LhfFjXjEd7PzLditBB1dcDl/06fJXS1aXHnyJYR815qeq2s58EjgggsmMNcQXX6U
aBuh3H9J0tRduINAEoM13fLV45tmF3oeFpgFFwZlIsChj/l4ncOrMVjE6Xhc//Up
Oi3/Sp5Re+YVhCrLitnIdcUHkbkaKRxiAcUl5/cq/ClkIZ8sb8EMtz16MQzBgAqX
LjQs3gfd+rERcHG79wGI88L8L1jS/92uc2uNeaVTmq4wGgrASODCE47RZFk2EN+n
3TFFmGMVdOM3cRGeSMWkPMqRZLYOBh70q7I4KuBXKKowQ5FjrHFTBQLG/a7zM/Lh
b3dr72lT1xbGB8FRETdeRjd2h9A2tXtn8PDNwk59fgNasRnnsZMn1ajvPIKOu+xy
8PtyaTeE2dgK/mz0ZjApRkeFs5GbZfZCDW6RfN9TB5A=
`protect END_PROTECTED
