`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THivhMwVz+jp/5tj1rUFMR/JGGDX83ZQJCpf2uFZFQIubIAI0bGHwKmtAVq/AfWw
ueCHDGLgRaMFfnaCCOH3TTGEvNjxYODiwhjFXz0fTne3cSZKTO5zFrbmS2scX/M5
n4RNfFpki442CNqZrZb5w75pwi6AgCTE5XpNABUofiWuLBeYvKmTnsySvZFex0hO
XycUu4sr0racIE5xm8qFZtexKQTwPK0NigHqjbUrzHMXXPTNwTNJdyLc9C+YyCYs
773es18apF+V3/v8GXbUCdyp6f+WLXjxwUmqFxVuq+M3eADt8ZvFOujMXfUJ7uBT
e2Cwn5S8VOLPOUEv7lVVs3PQ/3OYHsJpBI8RKm05IU15ozjAsuTW6ZOIfRD2PzK+
VW+saMSkdPMnU1ETeb/wjOtwyp8WRcUw8bqpvOaFw22/Od6YCPW2Bgi9X7IMstg8
COUddhwUIzaFpsqcw/YzIODoLpDe1DmrrcVFNFl51Vg7zWraF6FsmkBqgxMECRPM
uVlHkTNl2TKh/9EIeMBx33GaDhXKMxq9DwUIe+2EQZeOd+bUba2qXCbig+bC+bSV
FBcOPRq5vaJkdcc/yp0xGW9ER/mB65exGsWprhhUmXY+nZyhKIM4G56jZJT9Wivb
m8IErEnq41Y6JSrsO1FgEKADtmktYpH41AlVN7hWmHUbVvm19XGkyJCNqQzbrUlP
MlwUtKAzJGSUBezNA8nS3wmKaycgNIs7pcbrENoPJ2M8H1DSmR7Rcos2HjRTI9RV
3YjFtThnaHtOE2A4wlUHbtblqbAh03HLvjNL96Dg9GfFD1BunGDOVF3ZkcsvCfSN
bht91Ml+dwavwoqMIflB+jcXEW4G0JRIGwIFAzrajBOy3dRj03cPNjPzHQRNo4rS
z1LACeJ7jLpBImITIKBcJQ==
`protect END_PROTECTED
