`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZNAjaJ76wCmwEI4SJoGJSbWxyuvmn0fzvU+1QduU90W8z1fcRhGMd0azUPVZSQyq
lErBxbFcsR8hX95UOTBvgMstMKItis/Eys+tq3rTazf6BlnRqm69S6VMpa8IUYA4
L8GHbePKSGijsoQfkN4NK6f5h+WXDxRKifQbNmgCtS+NMWeygvzDnKH6B9QFr1X7
2jztiR9UoBuXb1JVjczhue6s+hbFUi5fXje+ihqUVrKZhyz5Dw6JggfOxMMYirej
44OvCAKz9VsHva48aLY3sa1QeYzRZ2qdSP+ugoCsYU4DVWCW2aYa5LgQq1km3hqf
9WF/T+yNGPTgaBXkPgCUoQWBBkghVIXChh7aPifglEhr86wXrQz/j/t/XVC3bbRO
Jkbv/76GLFuBluOYE15qkb2MKC14yXxlMxG9I/K6ggRMlzGNBb4Vg2GEkKLnejAR
bRND/4368DUMAkbe14i5Fxxm204d3PL+mAhh4tGQtPn58HoTreyrJ8YanXrgMT3P
`protect END_PROTECTED
