`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmGrdNLqC+9tkiSTy0cM3F4usgaSW3cawdFKxnqUVVh0gJa5T48LPK/5aeGo/Axy
JfqfXiIYmVHG9gOvlZS6Af8qNxKUU7ALgLygpoxavE+w8k7mKDAzyaAsy7kmuFSe
tXtHoCuDecf60cO93PEKoPsgOLvVPxThCg45wO02ZyclVYCjFClNg+jy1h0r9ZFw
5ayDYnzs2vSsjhijaczQQw8Bqjmw7UCy9d3M6/PHdmupd+3No6BgS1Lxv9oMVzaK
S3A/NQaGV6d0nepcj6VMXV/AaUEpUuGInJhklBvmwfJnOaKL55aMiAjixFm/s1mS
bIdnoHbFOyso0dg+mb27sQ==
`protect END_PROTECTED
