`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t9mx1SJzDvSjtKaNa3Y5LsrAFQN1sKvp19GQ3prXYQHyIahjfUpNLPvoiDMqwfot
fjXJ6wZUeIZ6ueWisz5fuAuSVhUixi7d2hL+UKB2qR61u6OUYu0DiArYWHUUAgHa
AeJotffIph1Uf/WhQgKxtJ7dmg9kRUHSz045F1RZyGgpPkJ4y2Hps8Q97p98Tyu7
hFFqmLG03gaQfBXWq4eFhkwvkTestiXTmzHyuFAcs62cjCRVVKxgSYAkpPxXBrnu
hyuCkEgpC9oCO9JbnFAhbq7ip9upIWcD4+BQBpBmrI9APqjKoXpfEUAThvfgsPw6
srYtB2ddQ+DWiZkT5lYYM4m74dNsmgJK7jnXUUisX+Y9tmA088+0AYlsTlpp4CJU
2BoIzkIboAkGsG2nK5XGESzC4kWggGDIHgD3AQ+85Iokb65aOA+VyTRE6qVVewcQ
Uf2juOdO0FyaqZJr+CcYpJoNIF2q2t+4IBNa92hFNAZR3CfbvRdzQMtjE1MwcgPP
4AYx1iT/GvJNBYaC5Qh4dsHV7EoFWMcvC2IUQDPlSFx601PW5d2tD0rFraQsqomP
4xcV4ielKPchfnC+qzMtxtP9gAPtUCBkTiPAKqkRIg1cGe+/r4y8UOilo0Tz59f8
NjnX/mr+mUPC/qflxHXTsQ==
`protect END_PROTECTED
