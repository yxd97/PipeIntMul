`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6hR3AQxUbHmzlbv/m9jInWWiX3OLEiU+mie88lJJU5TqEPzP7AVwCrHiwKTIGBN
zN0PIhHwUr5YeS6XSYiC77t4ApT6SZImBfn9pSGJUkFooxTLujy2nUy6z9Oy0MUl
abI1cpAawNbDRY9GyxFm60eJb9qR1l9O0s11ZPNMXMwMmE3RziDzuJupeVn2UYwX
gkNE63uIcdA3nWONnd/45jWQK8bM/6o6O8UQyOlBaLE52tQfO60m3ZT3GTTQBBPy
XyrRxtjmCaj5b5PlxC1LtJyvj+Bpk3EeiEbw2Sv8yWg=
`protect END_PROTECTED
