`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MV1CReDKOJMI40tu9HSMSPgtU24ePTTt5fQtOl7iOD1a+sw5SmHP8nuSFJAvRHsg
SVrEL44hzXkgfRJi80KEVGQc3v50lFrS6+mjbLwDUpbXw43eCRYTeBl2XbVu3r3Z
W53gnc6Cbd9UhDqHS6lOCv/cc0wlK0PNuiAoJUXAKTnXSrQsgcOoLGrnUWOcX8c2
L1ZbrIJwtz8kikxJw3WAvxaqhL6TBYLmtDdVddAdtA+RaD91/lAvoIoE++bzTsPG
0SToneyj5UM7FGgn3vvUk4lhen9g/ROT/zUU6qDqaqhKibLyDkd1VgIm7zTlGiZ1
/ccp6rf/WGkxYRLVSF2UI7hPqFCEY/M8uyciCbPD285gvNC0dHTdQf40u5umUgfR
`protect END_PROTECTED
