`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqxOeCtRVIBfTZRB1cz7sb3uIO5e+qaxnJVonHy1cMScjzRBipKWkoJS1qXBa8ej
xuWAj2uuZG5sj0F8sVGl0aAUK19RLQqNpLWuFYdTWP4izCVTfrUQ31bn2aCfU0wp
7+Ybj1Kw5tVAwAnkRG34yZkjMpRJ04RgnPBxD1jvnHoitJj8EG1uKNeIBgFzEUcA
QtIjjkmy34ryR/nWpceRcP7gMVvPVw6IBzcOnyn/A28uA6nMgYrUbsl+7cyW6xft
j1qjH5HpX5GR3vKQs98n7I6SR7k0ccLog6eq/ixongVRNh4soFP7hzvt+ic68Fw4
nt9TgZR8fQIqiRAFhmkLO3tsfM38iRETLQXOFabOVyH3/6aDj0ku2Zk7tExPhBhH
mXNVnAThSwscr5gz+lL/wQ==
`protect END_PROTECTED
