`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lrfRZ9+00oyZQU/6PUKQ/hX2tL3uG9of4odW09nCD5NlYgPLsasRZOQJOeH7ru9c
3MZ4l93OrUfhS2HmcvCKG2mN6axxfOOIanxt0w97VWY3pipcheBvscaKLyXoL+lJ
5eGeh6+oNLJhux5gkhX2Ne0zDKjIks8Dz9Ybxb442nIa123zkMsyDMGzKkep+ox0
rcue+eXz9vlbkIXo1E12pD7Lpms/pINvC/Bacd/1fczRQSEATL2Txl+CjHFJ6xtW
LVdt9WIMxK46ucvKBYm7QKEyKFotsfyKODQwkf1vMfz56vK1xJ7RMm0+daZtxHKm
llEruj7Cj4fSh2Jt1/LB5whAosHHip6KzjTetf59S9jsC8fHLz08+AMeJkpmJeQj
38UBwXFikpJ+oBcET60Erf0pcaclSiO2Qm6g690zl7FuSrFu90xtyA9HydHV625s
rdN4zDAnJrXrqY6DjB1CdwBRxlIcnwibeeU9SAClL96c0+/LRR0qmiHCUHIBJAOk
oGIZ1P4PK8N7rktvK2HIOrQSAdaGtFfwMqkHPIKPUiGqq9WnOo5tYZBiFxxvsSSu
fez3SGhDKR4gWPeaCOQLwa3ubPh01f3HdTSMwkUnPFzkH0uEEfBOoxNuE6nTy+6e
E5Xhvhj6EFLd+kRP8anlHyZOdey+6Qaz1ER2eauVKhNZwrnSP9ctpo6S8UC13NF/
C9hz82R/9dGgzld1VQGyOBuqv3zJSR40NjiGK3WhAkB3cjIlmTOikGNi6aLIK42D
TVVwtegoYeElOV2GmmYIaHq1Bwo7A/A7hxxP6uIs++lCTMl2BsPOk4O17ceNH878
8j7/w3W5M2og0ZRowrM6WJ/QdAX4oyI78cNHu4ni8MB41T+WUsGQlj3LfK0u4iSj
5QTiHpsN3GAGG74NIjtUCQmWiL99V+bmwZHTAVBalzP3ctKTs4cUSH2mcGwtaGgi
J1Epfl4iw7mZFIJbRUstcPAciCuZg0n3bdoIq9sIgxwHSc3lNkjWNqO9dglCsAvG
z8gR6AwUhq6cj0qANY3DfeiLxWxYLxgb6KNVDx8V3MyE+B+98F7NAhaAoHw2Xe9z
bJ6If7Rt1DKkwlBDYR0NknY4NgiynJbx5LMAGAXly2xW0Cg8Pc/ubRiTcsexjjfE
MH30csKMjSK3fB0chew6iSooGa905/X4LGJjJwNc1WwJ5wOWyvezDokWKjSlrrLW
UsgN/6kURxosuJvwTK7FNTK70FXtEoTa/xAx1H/iSUoHwrLjP4rGChqyClJmuJYM
gAXOhViq9NqD0tIWRrpYk64CragD1f7oHE2NaVSw5LysngGi4IkzhLI2kMhr1Z4S
m2cyyUev9HkeAE1AQocFxers1dSBnOmJ/5e2hNDFJayZMV94bzjf4o3TA18Jn2JG
Q+oFw+iyi0udYETHhG4webkJqFncJqVK+SF/xLXx50yBhEUNOPHiuYtZXx2Jj+Iy
BiqE7J5TOSfGOiRof+RBkrKqE20L8o19tYOD6IATSkEAbW2NrhYesPYU53eZSTSF
`protect END_PROTECTED
