`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUyleDqhyc4Lu3ebEGDJilD/4B5TwciOg07gZGTvSE06HtFa5pkexv21D9n9/Aij
UY2pnIKEgprAqLpBTjMA5P/YEZFDjIzuvgkQHuB2sIUaUoCajDdRbc/JXdYsQRHa
ogdquZ5ggMSQopVb2/8KaFoThQYGXxcdPAYrx3Wt4VZSTnMSS7f1P8OcJy7PlVB2
iDZ3oHxuWEjYtKfsWw4vtIpLG+wvhMsnCBLnrdaRp0GCEPsl/kYUfYhxHZAM0EW2
wqLCUI3AwmUgS3/0/Hjc2k0kxqiun1RfiMo/JCsdzRYnHG6BKC0+ZAGgeDtA0Sqz
hYkTSxDmr1XDd0zipagOQuH2cpgA1AFwwfkHFWxM46kdiyAkVzWf0ykpFJ81LuLo
HGei9o+dP8fQCpHj8hqoiS1ncJYdSj3SB9WUcEos5lntWd3fNjDoTw7IDegK+aiC
IzrknpBpmO8Alm4eKpGYlQAyJ2/EDrAMyhFNNwXwhXHO7CsXlNChGlMVZW13feAx
`protect END_PROTECTED
