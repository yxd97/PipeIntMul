`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFUKJjVICcK0STkBuYEWUgmWyh4UFO1USv5uBNS0/KmA4UvymN5SiCgS/NIflHSY
HKd/Y0XxPkgTG3qnQeSw0V4i58Xp608w4SBeC5QYa9+yVRyjwpJDhgdb3mWA2aN+
p1kkTDuL9Q6za43BRuhxctGTQceTJAayoKseFjO/O9gOqRMplbrPvryq2fpe33D7
IAD66zpweA216MomAFQjsPe4rgVI8vpxuA0c3axHBzBnMkM5IMT+k6ur/i40xyjS
qJvMGZn504bMFUmcas5YTvIrE0WC4Bhcpnh/PipR1RA=
`protect END_PROTECTED
