`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZeuvc8lKYFgMF1xXYKTFRTi51syMr2htRpc2Gruob1ZyeSpGckUNCgFd+IRJcvI
y+0e6Khw/DyGfk7iH1lqneXQSDWSjZprw4nzYM59vWQhISdaZConkXOityjpeu7T
SpCJtMyifmFL1qXNArmkqhhJ/OEYzQdYqWSlYQzYoWyvK9K6SMRr0BN8GCDz41B2
vEhzkzGrKgihhKvvquY4VjTQ9+boQUZhlHLORNsZ0EGogyi+Beqhj/FTjZa3Ve41
3SmSjdPnO6CUfKuXIjmcmKuPM0tkWyNmsVXWNfjrW2oEThDb1gVAgzYbKIdr1tM2
Tw5AMmcYdkN3pbMlhaIHZ6Yw2uXk+C0WPV4g9i6qaJZyzq2KrdrbsfO+VEuqDf+F
i/eiPVfCSoJNswzqUZYzbT8yjuEycqVt7LzSEyYqWvlqoCLpgzI/8qc/oVe6oyt5
`protect END_PROTECTED
