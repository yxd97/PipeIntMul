`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r67Nig1xKUfLhPg7YZLzH3UZbVT45kopJEo/oLIqGCDPY7+tDDDsj/lYpMi2T+VS
ihVI4h6LczcbfVrb483znTf6Lpb0bpBANg03UvaOvsjGSW4bsydzXx6accmKcnHH
AvEz9U0Oww3zwFI2A91ZqcNXn3ZtnOVg0n1QMZuhMBkmcRMqo0KG7ENgjDuEKr0B
G+2O+Ib9MaXIJCiNXeeHTW3zW9trvReurL3PF3alxKnK47N9lcM9h669+/LhOYNv
RTpO5TiRaapFhtyT++XRqP2utV5REgNvjSqLDkQRoLMFpTSgyXCD8Azzjv5lcpp7
mZ0QWUPUma/9OLPdf4+93XF5U9suCsb2IC2LGlrNLyGYbeHxM8ASBIbHKXR/I331
2PmBiAisxEIThItlJ86rLZMVaMHkLi1R/VTmHXuzxffX1X2IE2UHokUvZaMlJ6m0
Y9eMBbDdN/WPiTA5E8yjhp72sulPT9ObIev6rGWxHgtdF29dsXbbqcXTVB3eoMtq
/71WkHV25j6j9OhkWgAd01YtaU0Q03M09NvMivnjlTFKUB5M46xmqAe/n6q8pw1o
Kt80Y5uFbuHtERPTqvoIV79MbSbLtxlxtIXzqpaTxIYZFXSjOk8lu/zvfVCY7eFk
Y1ug0M+53cbKENEptGnfilsVruBcz5lSKy7ZLcFL240=
`protect END_PROTECTED
