`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+RiyTOcRUS91LsX6sj/m+qf1xF+4PC7Cqb07+ffwLXWfnXekDZ3x/8q6nG/R+sfP
gSlbuWUGsov0v0IW6GLlscMsQlKzqvCq4PIbXcmyRYxgirAQeT+uspS/ADNyHVsc
5dSVMvPDNuitQnr2NQydsaFDU4bjBugFCGJ4T7Sr9Q5W8+2ACRhngDNu5gcgygHV
I9Ghy/byHYU1AowJUSuDxQ2gd0WojCmBXKu/GcH1HPNHLmqWYBSapCzpdsewng4b
5ny/wJoKwirzBa4WS08UaiRHmd2gT+SJZRfD4pK95L/dp820oBoGsrVNImRpO49c
VpyR5/qZoYvvn+vmNL0rSkTar0LM6kaA5jERAB0f7v9tJ5XObXDQ2tqSdgQmJK3h
MNxSGXEa/BQswzkcIyJt0R/JdAJ0fZrQARSUTzZduB0=
`protect END_PROTECTED
