`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y4MY9saxZ3DIFCWkdW1d9qIwHBQfWOtGrfeVNoXTv8EbxGisvv/silz1F6MpEtyu
OfXfKeaoCVeHkAqmxHDVTeY7B1xv1mtEE/33Ij7v04HvZqew3idXZ7Hd0l004M/E
xFf49ijYfkGr0UCQOjOHMDTGwn8H2EO3E2DsgH3DNmdydsc5UFG8rHJylDD4RKBh
+la1KAZ2mymq2deXXdMHWGMUb5YA17MOgrwEdWx8iloPDLyCcLXPF14WwsuFFxrD
4eji8ND4TCVKAT4LU9+j5H9CK8FH9byicJdfpusGc3OCnWBkRZorb0/sypIurzN9
stzj1cVHvdp+bPWdzBystNc3rGZMpZsTR/XL09KdSOMp7rRC4SZgsWximNqiIwp0
oBYUel19Mx+9wf6a8IaF8BPoQg3a9krqXsHEXGgu8hTSo+QdQaf6mkHv2IAVtzmX
`protect END_PROTECTED
