`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8AqBeLK2qfBkYYWjG9b/+8BuopveIAYbZA/JVdoUuD5YNxScr5fNtnmOnHHP8zs
4afzt0oWrFBhRKJ6zFbx7QWLXt7Jql32EeNnxW/0/m8Y1HSk6NPpvr3X6LLMdw5O
udVjDroIJIxWXi8p9syrmk757WjXMiiWYMOXaX39Yxk3uSMH689U71BQYIJhnowW
ADKTzZ1XZEUa6imksx+BxYHiOTb1WXw9EL3CV5jEOjpCzUE0qJUTrfk7ngEdVh87
JLE/rPB/cS6hxDXbz83Exx2+80/9a7KoklrovWI8u0cB95Fs5HYgsy6z3vWgzLb1
nIuD5O+LeFXWLib3+dBVXBDBlX3692i6Gw65PVQtQyV+dC0QEL7WXStImfx9a4f4
aia7Twk+m/aJxJ90vXheb7pqVsa/ioX/3/x3OVKqXjLfDIQdj9H61+mGIVvib16n
4YzAFL3A4mDGS8byFjH9ex3xQ0+CnxfWo7jUVgcXBvt1yxONsIrgtWY3bnPyYbhZ
R9Vecrmc41hAjLQsm/weUf6AUBrXhFh9oBe00RZ3oNyRvSI2BA7iYUwN7LC2IJXp
3RUiyWimxk1iQxHqTRhkoQE0Av59noMJqeBqGWUcfw7sbdB8qBXZDih/gqV0USsH
GxHyNBmGHExPqItqi4WhPAGPXboml1rZubaBKhJsKyvL34eJ9gyfAEUAnGv7mWVi
eoXYQFPW6k9fE9UHtbReHg==
`protect END_PROTECTED
