`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4CsFmzSQs3O/zAwpi0TO9fBWJgHuvicKYxUMmQtNa3phRX8MH3Uyou67Y/7RFkwr
OBCAkFXbTZ9onSE0Z3Lwmtwb+48JgkWIq3WMzr/ohb/YEhFRZPgr4eWQe+m+jbSm
d3YX3sNMItMdZf3TlFX0KlR7oc+XHvlGqoHcFAvANZEMkv4W6xpDbx0KC5zwKL0Z
Le7N322UBU+jm2jsJ1A7jKMZNlMhi0P8KWZIB+w+SBkRzfWazFjXQcjx2LnQut/M
fhTSPcAuOSgg7fMBv+QduJiFPZ15jExsDbafAk+KF+ni7gvSblMcuKqdZPZhpc+V
5AsA4hpL9jCq5tI1KtLQMsDOkIaq5oRET2k9IF/7WXqgPlZveeFHT85/hF2TSelq
UJdvd6sMJrqOvTi8ltM17xvDFTMHuplC6s84/+vbAPcnmaBAnYVAYSc6IJZ0aKve
Fd1yDuAioJ0DtJlMbU/Oq6HHoWs1yKB3bh24g6Ehps3ZqgN7Cp5YxBj2oWBB4Ety
qRNCVaVzuhQpHfg1ixJzd2fgHT4qVhw/EQe2m9uTmHTTDPtMO/wR4JHwJh6plNdh
1NOsjCt1qi06CN9ipj7nxKqk0NU43qbogYis0GRxtorucQ+uwsFtK/sPS3x8hvha
4pRfiylLgDRZY3Pz9lSXXYF1mhJPj369ZSCQa9YrrNxQyLvqa33vZ+dGaaKaViEK
RTEpNbPPvPJ8Aw2HeBE7/X8GNLV6QxJdQxjX4M4+lHYthM9Fn+15a/8fbsbky9th
0ZNbONp8eaTwp3vSXy1kvSDBTZHZntsuvuJTrXOzIPtIKoqcv7u1iA6v7Gzc8FvX
Sna61jLQDIGW5S39rXnnk0m0O9vaFPof4UA9I7+BlPYAPZHubve4rHqE+yUpM+U5
Un/JARrVChQum51f/c3kGw==
`protect END_PROTECTED
