`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmLMI51Gic6H9OJZ6W6z778ZLmDbqPBHSp09TjVpHRW2a0oujDXthIk49JAwRj87
jRM39ZamcleB3UaBTA/0ons6WXrGttWEM4FpIo7EkbNG8WepLiFWcvCy1doQ7kK8
D6+lS7h+C6F+ehQISbr5a430x+OBzf+y7X7u30zDZmjIU1TjYOG95ei4VcX2lb0F
ikKCgeMeHa893FKQt2C9tbJjzQBPVJxzp7QwhDyZmhSDqjc7nNGnuo4RgRi+yJCb
IjKm4VM6l3NfxVRDdoKLoGZFBmFxqeyzr2cu3hCu6yfwRFhBJKDK521EgYmaOoZr
8i1gx3JAdxg6cefQZBxn948UQMG7i7L2ucbJkqHtB9g1d5ORYAfF9NhYojtY3b3M
va51is5MmkHCclg+IDUnKjwOWDc3xJyA82SLHqpGAjdfR8XX2Zgd4QP01xEVqmnV
SYyfA8mhXbOA8/GUwP3CSsQcZ2owNCQY9JtVlclMoPcbhGdaG6of9k46or4PIXtX
Lg7ZJ/UnEO/cPwAjN5MxB3VQUrPhhIOp+L443dfdXQo7M6DplU7VsS9McsmeW77u
tR1D7OV00KvsV8v+EBJi4yHInfKE3V1YsJKuBO80nbF2s9QJkAPFjt7SgBwmW6pt
cAHcheNpFYOnMl0/UUon7JVkw5uvOFZrJc7LmgVbpYQeqcJ62jT3hOImJATD1GMo
C4IgB/NLf4nqH0n/KUR1gPxU5wfjS8uSDZIZV1PdHTSe6rTWicKuZFJGxUHrN1/W
f45UTSJ7uyX17VUmhivrAbxS8j+fEqeSj7K0vvlAggoNFB2duV+veQBRm3Bl0KDh
Au9Oqu8cQhpQc9yU4iheyMsR//GOQU36k/0aFtAOQ7/M8EMJm6Ps+YaaH/3FO/9Q
qlRc6nyLwO+c4+6RuGQ6/SKAGB5Dh2tCL0rbl0MpJsl2Kyhn+7HKI9U6ELSLbCAZ
gVCC3ubjez9iVBPmkphBIe2oKQox4jwM5ngv8iLVeykDuTquCkPK6o+uox9IewTd
mPvXBGauu7RoPPyuv+ZLg26LY1z0ZmadykAjbu7X/Hn2TG9sRczSXQnmq8KXX9VE
k5ryZW7jpVllLB1n27cuF7C4TE5DasMPdmJN6UaSVTr7EHEhYs4Dvmq45b1e7XSV
iDmgX7Va+BWTQs0+g9Zh7f83cVbOBh371xN2kfYf7RBSExboitysSXimjZfZpg6L
6sgGpNqxA7mLCEda5rxtSxBtHRxYhej4p5WtkITrZbd3PwjBlUsBlExHy+NbQ54r
/ir/y+kduIhXtSNg4o4ak2UGm9oRO2S1cl+OUiGldFrA7ebdO6y6B3D0C4C0fqj1
36Umub5eYMaoND73R/qtQ8wQYHBHW3DVwRgGtneVsiXiuVAe+jFXnN6cdGVSuB/3
LUsIrifKfZ+eLa/6RzsngvCVK2rdRqWQpThsvFaVDiKGu2oO3Ra5GODFv8T5iu+H
D6QHtuG06CzAdhabfYJwl3YgWWwY0FxrZgA0q8fjTu6xGJtgdDAMttAJ10xfljhw
n1DBlQuAjyX7y37J5PFdqlYidkgXASwcpqtaM+qktu6hJViHBkUKE3mb25jH5683
NL/s5Cl/RDBzHHM/2Y/3K9vgqZ8g/dTCSBVT7LWMPdlGOOnZRGZ+AyXVnSOtjK1q
x5d819a27znmoROJRAubB0A0pPaxwINhCInotTdBi/gqzVfNl87CBNYx22oSkURr
YKyQ65bNxacgtaHXwHAJl1LE0haBNFwbZMzYUDKG85NuL2sQzuJFPo9Eu4vULyLH
apJf/sOpHBNDV2SwsCEg223wXmnxlDi7WIqyPDIt1ZG7SKi6yXxOVhHw93FvD4M0
0KhLkNOPe2C7+5hrnVBHcqWA++OUTEv3qAonCWJ+yJ8ZTrb3zQBTd6ATHI336saD
qaZDeLZmSi1v5jx0EBMqq0JsV9MVs0M6y7RHpyW5Hon8wef59M8sddjGDCpmfaWH
jS/N9w0gca6mLOd+FxWMDAJ3gEL9OnYCl0lwQDCR3IiX7RO0rUvoOzqv7Ofp/X7N
pRka4zTyjyjrTDJOKoLg2v10AMsFMKzVfFP/Zax9Q1mAu87UnRVyuLQN2vk7HZAH
N+VH3XvTVvn3zPUNbpUiNWFBLehp5T+gHGSCBxeYbrbnI0OlSHjQuuV/lQOMZQZt
UTzSo1dePtQqQwt0h8OlCg==
`protect END_PROTECTED
