`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkliPcb6k4XkGbgCUS0giPH9kDhh2MmYAHH0xc48Q+xrHev+pFmCxuu6gv01QWf3
tRr65JobvWKWVDehisofOqimvqxEo+QFtQvrqyrz/lgNpcwmSn8u7jmeeTR5VQvo
F6FYuUS32nXY4X9LyJI6MldAxNENJ2X9ybTGUDH7EZoUmxxK7EmsR63l2Pc1fJBz
C50VELmAd++AUliNoETMNbvMcq7LKxPGXxYpSWcJsoej7danJbiBLrJpZ8DAx3Wo
sbYwNWVhBSOiCIxhIrCrUijedRHkS2UJ+ENKLWqTUzQd7fkz+EC0AHy/NQt5r6Sd
7y8/9wPiLFqNsRJQ+5kKDnNCKLwmAYSDJNkd+orJI6CbNgMl43x0ZEtBurh3Vhcv
kq+K9+8Z3rUR2V+1HkFEjiLDzp8Gmi6fqe+lN8y5nfu2UricbnYm+bM1Q3vNvFPS
NNupo0lm2/6oRBklJygz0bWFwQ8gcii92RINHwVroPWPlB4HR8H0kuDq2IhICkir
RGS276l+CBfYMtcMcEyjYvs12Uzqy6ef6eroAbKZ7tYkU/r5/L75yaiQVd1vA3gL
8AQKjqAmGOkTjU35aenmAFnxQAAL8WsvtSJRK97WgkNcCks9rrM0TqupIcQkPbCY
9sgo7P300zuI6rNNeToPQb8gdJWkBkLdj1hz993wny5xCELu8QxE0YNV4eVHsZfz
sx4Lm2L81b2hFkfxTfDTsg==
`protect END_PROTECTED
