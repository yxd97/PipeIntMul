`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1CzvcDrHLO7DvtOtlZ5hh4TPg3AmS0lPhRdvxIfFGyGQsRpo1A0kQyJ40SIltRA
hU6w6YFYzAu+HP0RhHF64nPcAAa1oPh2CFIa8y3K+UwzCFDVXQM+Ud7W3R5KiZHU
FoPXQ0WDAxNYs4b7b1+HxZ9nTgCkHXTpHsMpJdEzllqD7UGGsMlQLeI+qZOKXEAd
jFAw3QztIGjxPD+thO/ws2J0VRRtYd9B+GBvRoPJ5BtDq184ZrI3YJawBn6Iv5+y
hz3pJu6v+SKvR/OkWQPgSU/O8N/5hzUKl62jHDVSYVzvQ/BsT57D6SBaf4AT86wF
5yhQWU8b6ULhRPPg0spEGUG9XdcFysA86wjNK1mEaTraK4wVZoQmG0rTDC0Cfh7i
dgzPOFn7MttQAMCMlNBB2H0622nbqhde16K8hevd423zns0lTzPa5YmZ0+HH+Bu+
iY8ZdLivPRnH1qMMRErmqC9sRI+tyGjY1bsZDyYc4EE=
`protect END_PROTECTED
