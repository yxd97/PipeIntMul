`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFEZLHEVIWq/CU+on/ogPs7e4VDk/8gmUtsaK0QepRpVsbNMUfGrNL5oLEA370Kq
I4b2weiS/URqkAVc8/NMAUvRWhBIsHeglHqE3N431sBwwynR9X6oFu0KwVB5uCxS
aQJsEJP+wdStZcxXHMcKqq7CnaQi0I4b+a3+vritInm9Ya+4Z8x/r+pnd3LFZSLD
KkY63ke6nWQkDcVRsG6jAc60nspf5cR+hQJ89KGEzoc4L+c/nQY7J3HulMbPeg2a
HuEupvZxlg8pj7BDd28jK7hPLR+CZnNdiFZl3whI7K08lxmkT+JFM0I0cPrMChb5
2sNNvgVecg8Vt6N65bJmWtSNmYZAt1PvXBKwcu4WbgNFNA+Slt0YWllsQDyLxvCP
/MznEg9EL4XML6EA/Z9yIA==
`protect END_PROTECTED
