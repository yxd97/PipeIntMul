`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zLgMXMxPLB87nweCmi38NVHLfDOQm6SM2dUYevowAuqh2e7yYxDinQC/aeK61h/P
EL78rYO+oMo00X06+LKIcBKnMaI7zrFkEQpXEEGxbiSdDVv7N1svatUHHdw9gno9
LQ1qdzbGPNNJL+2nmKdLO7xD+Vr8VBZuyn9w/qTEFUZBtDoTvu5G2dM+KwV5lm99
Xrh7ZKOX7EMIyJJy0xNNZG5QYW5KbIC6Vh7zMDKn2TltwDifsw1CQOxOW0bGE/K7
nQNgCGYtxViFMROw7Oel4rI9TWnx4uJiZeYDqRqfGq09X0w5kOaI6oMfGkyr1Zi4
+KPdCy0nOGmEhkvqvqMkG4QPZcNVFPhfI8cBFAzC2DxwBJs9HCUpvkovnR/8bMc7
N5zIwPrfweoYPI6nDUPyh7OujTLuZ4J5Z4Ki4NQyU2qaiVOZ89+UjDYg87+BLE+n
wY7E49JSpMkhRzv0RzOaxOUkLCnQvI2K1qN9XjlhCOx1OrTVhF0FcQwOw4FHhNjw
DiBQ7BpCB/3F2v2EK51C1WgjU6IvL9Ep1jMCCVfN/7TtxFXiS6pe9MwfIjXrDDoP
8svI8CI5DaIfaw0rN1zworXyk2ecJFLwgszvtIE6pNMMsUv65tBOsbjA14UBr8e1
XS3YyC3+tcXXEcZoDmSd1li7VT0rgKGuWqe5lJPjHehBUSSJs56zGt0y5GM67+pk
VCFEwV6FQNIpc/CMcZ8FZhsA1UcCoCGwsDkuDCf/gQks0oCS2VeYG6BLZ5MkhWTK
zkHpjj5sTvKzoFuMjDjcFtIVW/1hqVnZt2RO1KVqt7gx7Z/KrDqtjay0m8juF5K3
YLvwYOiU+QYB/2HkaFmzZqk7ijyK9iq2PuJQvBT0kZEF/OWIpN+lbdgvazLexrCk
O2vyFj7DIWr2t3Rmj8TWxrjfeWDqbL20S/O8QIfiwViWcTI+/bksJb05+FmGYI9o
NflplIWWRd+WaabGFH3PDHMQhLpABZVV/buRg3R/mdyEzxPVzsjVtkFiV/AUolRC
0jp0Sj3fgoLMxN1GvsxXmSAHdLucwEJ/vyzTfWhhC8xjLr74TEngQvuV7+DMkwQY
QQz+qYri4l8bxYxcmNo9JHNSlN5Tq8WKrvqnwY1FMQmdQTv5YAiZ9lEqJC2Qsqcw
45uucHrD9QeWTSJpqJFMZcHpq8ec7j8mZd7wUA/vvBH8HYCKaE7/HykmTdoHUyQe
JJiK63IosA/Agw6H6/Re6iJ1yU3Vl7KMJhc8KaJ6dT1rISesyl5N1gzdDBnpM021
BVgu6W878A7w8FlYeOYrBj2SUja/WKtg7CdOPfGKyBUif8PcK0oNHV/9176CjTlW
fyxIM5phr8QAJF8s48xJzXWD1rJSTSKXtOZLh+VG0zt0B/NFOH7S3RWiuPuorBim
dQ0M0cSRwhHHmaIHramurFLOCT3mVjEqN8c4RNL9L5SBuZV5ZhzNv8j+DMFUZwul
U/+bJDfOIhi/ZRyxovBbhcW9r3YnpfdHVq8Y3+D9xr6rsFJvsgZ4Zr43jl73dwyc
KO0sBTwXrLMAUxHufv2B8dFDaSu2+yYmc2TwMNkT4C24Busd3RGKK9MVGcK1eAOl
uDJ5wSBpwYmGGaXCGa3w09P1J3a6zei51Mdh82Zm/Lt48POMYwxM/wjy33sKg8+k
YEl3zv+VJ6z9hqaKbApnrHlHD/U3AAUhlgOI/UihZJ1VI0otGvq5oCORoLXYx1HJ
TPxWWtU7T8WjPnw84j9WDHPEQD7GfNNZFa5pWP7dQOtmQT1DhQOt8VROAqmiXTtx
+1p7Ooqam+8Hd4coPBuPqBlv4cc6sV0sPVvK+kL6M0uq88gZm9G0vKh6ss8wI/yx
brgJcbsahq237Q6oxckB4Fk1Rurx8dF1ZBg20AgzQcpUh+/mLh7g/aNnLAmem2p9
`protect END_PROTECTED
