`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CzxdwrfYrvEEuvd1K3TfjJKRuohlb+eL5I6s0tO93W3Ts3Nou1joTB9GiKxjoWK/
e51VhLNA9PISfAzHaC0A2MF7n/TKV2iw3ce6y0inumMV8wyoE1pFV3D0AY7xtlQw
+bUGvGTq5f0ZHZ+8y1ZruS3AOQUH5/I74s9zHSsKtynpvDR7h/UHeW7qTvZ+3UmQ
iNeiGK4Ze612aUFnIz0nNpMRkPH8xDOW0uuptxw8xv3JwpsijRKOFe0Z4CoKm/jF
+KVTZUFfwI8/BeFdl7m/+ZauE1jkxgh0ArAI3JH/Rv9kZ6A85lD8edC35JDXZRml
9+2hq/JD+rnJ/WAQMQ99/1jcN87ABwYIS9Tcl+mijSUb1WOTNW9XlrVaqhdk8o5w
A1GhTwQ1jEpxHTgCfUlXqg==
`protect END_PROTECTED
