`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8KmJDv+m9KwOhjr+336z8BYsnsmTXEBBR32au+r0tp4aQnRIWO1OPO+0uIlfBZ/Q
sFyPGnWzrcX/s4QcLewNyFnrOElbL/Pe2i/jASFMNJWGmA9YF797WQhHp5piTJ+b
0kz+z7WgrLCbIBtWzhrsf8hKNpJ3IFQSIwSfCzxm+NYbKMf4cnNOqAczSSGtpT3j
Ig2OFRXkdt94bZAEkDxDkuWuF5zVYgpi2te6WSGtn+UpEVS97w7b52Q2I8maH/WM
ekMu9h2tWOnvfBApvrB7VI70iVMeRDjE+d2h8WctAASG0B9pL3EoYAATmwGlOScp
5bBhSs2bkW8SN9uF7lG7x8W27tEMjCDXw0VkztLVYt1n9U1VMMxwh+nWmnV2axRI
vmmsd+3DvGZ0/N30I5rGk9zeTb702e/CNyRNoyNgjsmzwd+3kjWqo8/zcPaYfBbV
PJgEXtLDYsdZK/a20hXCPbX362NSQpeX3JB/jvlocu1AsqJjsU9lxhtIfw3+fnLZ
yJMD/MNcQsB5wfWJr2BaMyeAfcTBquiYqXMtTHnQGKY+PIZVNh8lFt5RIF0IRkOc
MDAR6iSvBpmz5kPeQUUkvcbC5RvKDEGs9/vy+QWyonRsm9fKTDmLcNREYpb3tlku
O/dSTUEN4NYHptqaKifY/xEQqPmh97xe+5hoIxisjjHs0NbiNme8Q70W6mZbmvET
Fagmszy8Osj8GnvIJswMHFPCCr3ZduyC6oSAahSjYKWG9oTyRRYqH9qVvidmcRoQ
Gj6CWfrxv8XsKBXm06iyaNwq/8IEk4WlMmfJprgKtXNW1G9TsMIkP2WwBu+g2UEw
Be1/FOKmf9awxMfMBE3u33/E2uWwRwEZweYFEjv7XHmTUXAgNw5OeJLuLJZqHb5Q
V0avw57XpQpYkJGJX1V47HuTGD0gmAuSXFHDZGhCJeO96fUOuzvZ75LGzd2kDqpN
wUWBXE3+khWE5pyfNDyelDIRPupzotErscHZ0BVVHK2K60JlsJbKnGEg6UfsCzPI
UxXn1SRIb0U6gHeT1svCb9Y/suUA4wJVXjJQNvVBp6Y1Qg4WVcMvN5U1tdsz6+Ct
1Dx2BzUlMizyr9G8H2P/vcD0FPdk2DKwbbxzuPlvC6I6mX4X9eLZwPGQ76ZO6QKZ
+Nz6i9MXDMnC1dWkULH1UY2U8ZAV6RrPVXyQc1nh9jM68zVUVm7xMSXwUDeOZvcx
HERW/RdR2P5PWwfB2JSCkjg47CWMxFydR0chs0Gf7oICRfCxhv5Vcgc97Iq5v5rO
A/42mPfeNoSheJYW2iM7gPcK2/77cn0dq4RPqe1SzB2R7axUIwUw4GazbtTUKwik
BAg4gQx8PSfYo8n3+zx4zF7WKHKVEnTBIxdTJolUbOX/kdwVQBIbV1yk3nb+qzrf
bRoeM735Ek95+v7n7xJqTQm8sxt5vuHbpq960xNa9Etuk6sE3gx7dcGh05p/M126
wPGmj0FAD7/qMJVaMtiiPzNbZlNOYjXnYRbdXs3V3usvD1gmSU/V6KzDVa7EyrU+
ik0rBXkpc9QNmQqhjCUvmdqcabu8JT6/FWmJSUeHJEJXYWaER52yHCfRYR0KQTZ+
ZOrYUnbNZZ1357vJOEfdNzowETl+UX7Th0UwWhVqG6Xqhc4WboJEehtO0fxCVHrG
9QD1cMxlp1352ACSYQ5yQeb3xWoDG060CDG1i/+Q/Pj8JU0T5fB/M0Mf7X9anTkg
QVXDN7liS3IjxD8rk/4ne867CqH1LlvHs4QqqbxgSyP9I0Lh1PKBPY6jbB9u/XsD
sfeL9342Pji2UAJtWp+mS1BimaSOxZYJ5Frk3wwW6fIb3k0uQtKgeSW9e6NISiqY
P+p4Sy8E/NJlrCIS7hACWXIbW3RnyrFklGCk/eA0CBkdyOB5t+p5o69Tji+lSXN9
S/yWLNXCoN8RHYwewzEQXmqrtPH1s0y5QcD4e6Pys1NLT3TIaL7eVGYkEPQLlPtc
SZz853L9C3xO5hbFZ/BhG53ePalqBNpJ9go1ZwpMFXl7T07l3q7RfIIgopM44/eG
fs++rZ+/sWN0PeMqmrts8+7fCoxSBAlg9okVgcszquvg5b7IVy+xJ7KqEM8WWvfF
s/XcmgfUjBHTMoHuBevYTlOmOpF65E8nGAUL92btYcsM2QfHS4f5z3mkHmWtayIa
r5aHcEpVcP+o3qOaXoL4oZaNXT0/QJ59o7ZHCzBZG8oir65VD6C0qtDrjOcNPrKd
qXTXREe0M3J1piEbnJrSv3xvUtbrMmdxLfvstKgLMRnkhGzfqg2D48RcRpS1rwKS
5DYfZ/Z3IOoa3w8h2eOGefDLige6ruZHV1CvTcnASfi2MMLMVOOFr7ILDO7VcXvM
zgVGZkGebqkTgt+davet4VPybQUnuCjncmItYBL88nf0aFtnuie2XiIJoqUB7FLa
8vFMxLsAbFUJa59CsMOvhGXZVM+icIRr8zTE9Z/cqncYt21A+iYEyQg/Ok/+RciL
upckYu++BSbGN4W1q6xwaUTE4iu7D7UiRPj2C2Aqr4eT/gnRXJWYxc5KqovusRSX
90osCBiS4dbWhqeyeLvA+QkyFO/cEXhuI9xAXCXtBhbS4cR3qEVh37g+34PlyLjv
BZNKGqqGko9Kf5C79YPWaY+/h36f4L9GS10mwvNKKiIG8XER74Fi4tWm4vX18VMF
i9x255LFjyNTIdIqRfTs9nD3VdDaCEyEA2OwW5FNwvFNJDso1s4IxoXlCN+LjvKj
bRbrterMNaPJCSO4MjudSxrff03TyI18GPTVkOzy/HtGJDmDvrlmIkpMB6FTct8b
CUp3xhjafV/XMYmD/e4whP7KZHGa+28RYeI+q8/koi2hyHSjEPPnRry6aHqWzuac
lde+/u1r437BAHTeZNJUUIFz39KBR2SnUkBCMR8WBI0JiSLq5FrXEUCNURBVI/Q9
`protect END_PROTECTED
