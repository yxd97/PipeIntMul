`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFOh0tVwOq5vgsWOZOpU8S0S64OQnAG3fJdZKH5zxABuNVD3T794wVMcazWYfG4t
/U0Z8sK6OP0Xi5GCRbZUosz/PmeF4dC7K4dyuH0QtppG157SqJuOuZGCZ1lX1lSL
6ma8B7EuVNjKVTeL1Ax7iA2YJb3sSFOBUlDjajvoHU/P20AqI2PaWK7hWxr1vhMS
wsrddLaoHDyzffdcPuM1i35KQ+l49Im+QJWkRNZtcHsDJ7N/ulHIWntsn+ELXQ7E
vZzFcn8fB3kLERlSBwj7k2Sao5YW2F8nEgHYpeIKsST1/6+A7xnH147ZJGiiWAeq
VB41CK//EtumXhQhJLkR65qX727xbyV0wMI9DN7ahj1xm2yapZMc+lcTQO8TN7TQ
5Cp9fPTn+cCHYUnl7GKLnjqO16JUf51SrhUsaCtfRMac4XG00vpchFZOk+nsj3XL
RVO38owD1kDr4x0LiizRvViD8XyHGR6/WpGJRqob/m4aHVi3z487Lz+uYhfmhxiD
GXsKtifEU/XuekYzwzCKbjEgy6lr8zWtjI+ClGXWm+6WJLlzetFukzT6ApxS7EQq
r1Au9YAF9ufaP9gt7RUN/e2xlvJxfxVrHSHc7Mg9aUg=
`protect END_PROTECTED
