`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZMBKwKGwclXkixAVWzza+FwKWVqlz1m5yBYOcGrEYMXPRQQA36RzJ0JDCW7aG8bX
cFdFWYqZIuoSWZTOAz0vhMHlVQRQxxiHW7s7iRLU6/6B9ZbaIGzOwhyB2Q07jUOS
TQ1vWp6ZWQz6XtLLhp8U8o+apEd7QB6CHv+Bs9bUo5Ws7iU5oExFDKI1SdP4oRvL
y8oiChwiy3XE8Y4OADYBUjDThVtxkes/QGqTxD08k/hiqqwyqdAHwVY+qOtB3LHi
qdoZem8W7s36yeIIwzAnY9iJMoFaoYAGhUZ480rcyohCGCpNtnKQWCngsatNAmhD
4c5ZEDtdBwokfkCSImzSTGYRHm48fU4+6sKnRZ7MSVXAlh88jsjBUWfRezZ3lCQy
f7CSBY2Z0kWIR1ICAIEQqTGat1Q8JFD2wSFgPtylcjwng7pZrUGDfAdTb3UWnxQs
NjE/tcmkq60DzHbmg1EJRMbOuiAbxrqtpqC7YVfZFTkCVTj5YT74mix+YN2Quvgl
uHZd/c0IdLbQSEUjjiSzqwAoF0EZB3PdLBboB/h98uVf9a+M0o9NogaHq0xttzJt
+CetUwOEAdVJxaBQeKW2iR7+zKc+ZSx4NQ+nVs0OLq7JzvYv4NLplgCzpudtHvP9
t5olSv+JKqgGUm1YgJFqWyByZX4r1wgty56DBKPvXe5WI88QJ4r+8lBziLAT/dls
iNcxOOQqbuqgcHj+htrNHbGRaMw3gHEyioV5KFkmmabNuB6t991NeZKvD9Ka2cr3
iNJJUfaCRgmkG2O2sUMT/pZjZzVMxuTN1opPbWqAytQDOoLGPAb6FGQ0NxOPR9pk
BmCK0BYvPc2RLDRKpQKFjorHf9RbxHr5HuFG7jay66uhLoZR+9tmMhnKcEhlryfy
l5TYMVnDCfmADPyG774HvtESXEUnZC6WSIU8We+I/cIbMhdu9qWEcsRq2ncHhX7C
oeuz+0TuTmd8G3SxGU6B/gJOau6H32VynvID+MA5ItCVtbnmrLqJUDM81KPMM5vC
6iVwaV+hmOdT/eV2I+2M5k8ug6MHXMt+THpIzhvnu20lqKMiZ7DsewS+R8WZ55oa
1WsBiTcCjEU9j4vZCVqEExHh2ujI1EaHfXoZ/m+aZxl5GF8CxNzxFiGf4bFuX3C6
xBkQlBZ1z0MfsrlPfH8F6vQqZ31GagDg9VtlW7rO5qr4CiPAlWy+f2Vnf2EBBMFp
4jWZoQd6lMok3ASs2Y+WvgsiRlpdGSWnB67A5TxsC7ZELEar4L4qalYcxszrIDiN
K80LltaO6APgLc6ZshOSYr+z+hFd2Mv6NgfHLRnk/flb7aGa6tsXXbKWTEOUH32Z
sPsA43Iz+MBxYj+VnrpTjS5QxDOUB+S9y0zxbRakLHNFCXce4yyQUhhHBNTC0mfG
Al666RUe40+I8gsu994NHZODGdnC+M5EfjiTnjUQAHEYtHjTQhYhk0ut8kfmLi5g
Wx4ttzk2dPNS2qBYZGB+pVhDmOwudcYDrchmKYgiWLcn+Ya5Fd+RtfsAxRagQfJT
JSIwd1XTzeFWkQS1tJ7lUOLpZ4iZqrRAeTZV5ky4MopHraPdXuNhOFrFLdAR/JQf
soPV0mNqnagcc1WOsilbSjsj4y/7EaDI3kGjMG3JBGZbFot7xTG3Vfz9CcOpwGUR
y15ntLq7/Ee7uK3AmI0AECOIUtTkCI8FPIi2DPUhTUA9DnqW5Fx6mQ605SSG538a
A95lMqDD+XEa74akxcygNOp316URGL7BPHox6mb6K41GJQj0jCACB7Q/G3YpilBR
Zuw+fBpmsGWgqMs494aGo2NLemNrnG7E7AahNrqGa1+5DHRbaWJcGYtjXqHgB82P
5xYWWS9YvrGKc8TTNT0IRGkgsIICOLeil4fv+wbCrdVEUpnxX+K2OHm59/gCb3yM
mtsjPtruFHWQYLkBFUTQEA83ZHe+HPx/nFG/5NPnxC/5sCrPQQ9SVU+vk0ln2eoO
RnTpCzkjFyO+3E/qrrx6z21Uu+MUCtz+xiUto75r/z1Gbj87hTc5XRUiNktNmiHS
fbJIRUHUDye4ISuog6HMlKT+utP7r1gitmvJFZoQSmOXcTeg7EfWFSocitr5Tyun
rxxlTd4k5O/q0BeHecT0/l4NLwhCFIn/hhCzcSngXGaAW4yyU0GbTt+GpnY6YTx2
bjAncZaldXQlUQc3I4F4UjlXcnrN4DSMcqcNg0igJvxX9FZoPpuOaOkut9JxAU5Q
d9hBOQk1213BPo/mo/R0jwG0XemV5+Wrp40fzIOhA4SAeQemw4/ComPJxpPAkUYg
tFQBtFjGlbDEsQ98z1I57NX1HskbN7vWK7vfiIArnuugpWre7E/PVPY9/cK0U8sw
ZbxkoxtwRFmKtVck8o8ykN+kj+Y+fmhEJXkcGP2FoIdp4wWOiMkkv5f5aahYlNkd
sSlh7U6G9VUjz+VdZxlt06rYWHgm58pZrJR3cYN7ApePbTztN5wbLcHufjifHrfH
tcJqiu7SptXNXHGKIjHjL+psZjNRvnmO3+esJDjrB26aoXewahNL951O2DQ5jgYO
sU0QUgtjjt+6XghiQZic028tvS+MVUm0P7UHKPXj1RsxwKetScMlJiF4r51mUREN
3IpUy1XGZs18CdJfWK7vlUTtklgYdtmEzI1gEKFQfz9X5bghnharlSn+yv1evNYY
mQr8Z798aTjFxnEGRFAg2+PZr6KRbhZHP0VYQ9mZT5r69WeZScnRIHy/BIYTiYxS
`protect END_PROTECTED
