`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPpTROoHCYFy/sJEYgBq4UA15c+X6qkAuTa5XVMx9ZY138xB5NOgQDx6n8lXaAwQ
7yAT1mApuW121zTeBD5zsKxWmXh7lon8KSVfKMTqtZ0l6aK2PvigKAPwYSc/lkZy
jSGUW3ifjfnoPimwdJyJcF0jq3eCc4eYPLb3fo1f1rEaId7CgFKZ8HmKlNu0O/ub
furoDcZ6CTpkY/zsIE0zvc99A+1BBTBvvbU2VTHwAGuSAf79bcq9BOrY/wpPa5rH
HJARP1MuNISGiB8XIu0cTHv35YmqgUEh5lMnIsQcGDGqyLjBARLdcKbsvxC8LOdQ
/rmdIuScxGYRhbqBjoYP/QxDeDtgb3HhqFii294wi748XtCMnVg8g3j1NrMfceG/
pm8TH3d/5CyZuUG1nM0sFg==
`protect END_PROTECTED
