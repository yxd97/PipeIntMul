`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/WghP+P7INDW+SaLFIojuF4s2yOfaYes1qqlB10NY/g/7OLxJbhgmkdy1vSYVLwV
vjU6E/qB3zUxSnUKc10wios2bG73YAPGKgKlV6dQZCQBw3/a9BghokKEvnRgqKhm
/qaZWKgJzlEL4KoBDHjC5YJtF5RFIFIQBUpO/mVsJhqJkBDLQYdFFntKplDW+JWI
VxDmQMTwHuVeJ2dWqc6Axn0pYNd0Q6PrPNhCfHHYlZnIIzcGierafiOLnyFbwsLm
RWYk5clPEyjWv3Sgdu9MO8SAbEwvq8BONFIvx8R5x5TCPe20JNv9JGOJqEceLmvP
Bxl+JhHoT7yIOLnwFL/cCY+najAfwLay+oUPzUJcqYP2dPudCGNRkWNF4VWgKoRe
KyKfPUFda+eQRU2lM44fFNUjgiN0EWkViVpfWiqknZo=
`protect END_PROTECTED
