`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5hBhN0R07MkEdFNIaVaEEgHYfqP0Y5vvKPo1xb9S2OaVqVw85SWOPfmhZy0ucZsk
Z7nKQfd+PCA4ZGzZVt38NuBXW9VeBcqxcEiFPP8012xuguembjgscjiPWteoNhJF
bVGfE/XnEqVEXMMtqoyNOVKtgVTDMQ0ff+rtQwcf8Rhizr3hNBf+UlLcp9SOWjP/
LCWb3Gt7fNRxM5DgeW9Qspe7kNyt+HoeL/UTOAMmJRwKOPVXNWwZjBaPwdtRdht4
7B16XjA7u7lqp8uqgNIFlE59NiGXpF/PUIt/zyJzDmh7C5vILFNcCUyNpebOc6X3
PgpzUY4CE7LVQtLVr9q6vz0pYpCNy6nPkXyKkjGu+cydauJlykF4svTRywltySVO
6slUdw/vBaYt73MX0fF5zIN8QzAXgi8aLdTTmKmcs2VwH7g6keLFO03GNWauJHTW
z0aum452r4Uhc+MWOvAFMBVNgaAr0jiQNMie/SOq2hTLngwWf/V6ih+AnKfnFGGE
9RvDzSQPMKRobCp4gWodNwJ/xlc57Q76MzmPSoFni0/pqZJtFWZVZ5l6sWBzCD+h
zynKZlanhuC8gfPG1oBjWNJU/qzfOjYd/oeeqLIqOcXc+ojvTfYhUMnF9Ju7gYZU
F8cgHTv9u8IPCkjnXfg6xeM0SayTNXCuWEsX6FVB6r6QIQ7y/wCC/QlFM+4IjyVw
CLPZOrZke9SKH/aXpeQtn55F+4LuidsIoi4T6LlMFmUWR6D7GK8BP84ah68pBYGp
OAPtqYWZgoiGkEtCTD/mPJ0QVuTHhMvriPeA+RT9ftOQIEde3FMa7uLEe1zaQ3PK
aUDf9scMDqW5OA6jfk7QoA==
`protect END_PROTECTED
