`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ss2bpfO6+DTjAww0rSCwkNms/aTxX1CFI23VFNKv+qyH28iSyLnEavtMGI6ykKt7
xsr5Hn8Syss8fxjUB2BNp9KB9/J4Q7uTMtT4emazUYkCHbjzfJTYFcwTLFakcKJE
UTNJf5rnOHvpCXVIn94NTadIuO0dgryfIHpFisFUGsz6XUw305jSZj9cdI/TT56i
ieWkRNWN121V6YzCpXQSHiYYyUajjcRK7eXyRmQh9Okib/S1L5qQRzdwPJXUwePn
O7AHZeKMqD5TfNBluU209d1f/6neTv3+E6De+5OSO7AJ5S4GlXfUfxcEFggmAnY7
v7KleC0GtQJIbfehlIHxkismWQh9SQj9yO036hbGkq4sfht4sQcjRQ4rrwEHjt2a
XC8gVYxpuiq/m6gHzjqj4Zdjyajk+pKFiamnRMDxgBycT0klsjzFNdqwNp3Qd/Ot
1ZwDDCkF5CnjML+SOMLctOUU2mUHHpHdBrkVyszH10mDWqc7rmDWRaI9okQdaRto
0qx4Nat4VWkBvh9Ay/hOWdLe/L3vW/hep3XEQ8vAN/hllz5240Rr+gG1ZzpKxek7
KReZhgRmjHmZhDlmRrUNQzfHHZyg965L+PM51aHgvMy0PPXY//74fanx8/KiWggs
JgjKr/gwpOP5SBcTyNgkBdr0bglGmvx9Ia1VrP9b8WyB3KMlNQThWSVmJdn2dX44
FHgkk/N8iyPYftglg7eg1XI0FqDIVNnmTEjL8wK+VRD7PrY78mhTQohKTeCZQkmH
V5QZpLt9LsvucPX67hBuxO7hr9jVCPzUqoGpQ+XLK1fbnLqBFKNX2c6Npla/gEQB
HSAcFo7FNaKosf+oEikSHWvFuvznAXGYTrHLiZAZza9R1gHSflwZh/kK5LqdDjue
5IvoNS0QgLMAqIEPlaFhhCnfIJUcPkm24XVojyqo/qYnx0okvEaNYcF1IO580P4M
liqrjcrJMobIYYP4krspBy9ulY9PZQ9GHDVetuzr3Sc8J9w6JwS/HL+YJjqZr1JP
H3DFpuH+gxLJePKr/5qt0XMOSm4nKSOBbcHZiTHi9bo7EJ/HiECUKouN+wM6kK4L
dG92ra5WlptTwWntsj+RVQ8WsZUq2rZ65xymhqStM5om1wuX/mZKzBCyffMyklHO
HAI9kNazVQS5cAEtYGA/hi5zercEatN1J71FT5Un3fuSIzaoYkZfj+BajZgqg2Ya
Y3W1aAzvZk6XEwIywaJC2pOfiO4HUBtVxMfZEfiYEs7N0rx2KChMu63I7Et0s1Ls
dRxHpbKTdL/hRDwPMbPaRayvwnjgfrmnj0s8jncdmCGRKUn30EclsjqwTrEqBECO
NKCt00QdoGjXFSH4d3Hd/RBWAvzepTS9ednGmcmkl8wBOk8T/Q5TIo4EQ0FWYy3P
B8YwEpbQQR+0fsGbPsZbSmmAk47hcWje/lbhMtUOOivNQ3G3fteGCqixfWCMHv98
irk0Xejc6nXX92xLDP/jse0cHwD1s2HL0+x+qx8iaURhGWaYOeFDCEZTHx/o2n4Q
XNFU5p9UVwIZivZ2vDMBb/y+6PVebywswI1FGykdGRV0Vuzu3btSsofqnEGxAB6M
yS6dd9bVPwVZL4LL6apOH/dAZxE6GsL3rZzWmnFx0DvlsS5lLUHr2CC4tO/iIyzF
BkWf7Oh4a2xNN2JB1le9NzcQgOA8BDKfxE4XiW/pxiPBJuWeFtgVhyLGuIrJmoai
AY+wAGGYMTfZterM93+RbAscuyr/XhAo7eBZ3x/3B5swOn/G2dzOWkIgGnG6lbBj
mDQ1qlqvblzF1AeuFWA+Ts6Z9CpkRTg1RUVs0Lv9Wvl6m5YNsH+Faxs62MCfX+d1
w9AEyXcIsLBT6EOeAdcafdruVCoRAuM2DuiX96GQPsPHpNyCMkhk20PJ2iCMJ7h2
RCpAR8WMGMFKmLhfS9jyOAt3ZtKYNnsZOhgPE4OHVkJVBvVWkbRXMq0SNcnJy2xG
RSwgr3/TSBUnxGfFzmjFmjQIonM5mx20ujxMXyP2WBF9ZjEfRLWdizlLSJvhCCHm
aayUOGHFTDEQQRSTwxbboVRDW52V1m3ysFNGdONqh9JsmyUjegwwaR3Vj/t5Gfy4
XlV3DYFdHRHLPNG1/9Sf1HKLuqQ2u+j0tsVIdK5Y1l9s7wI/ck8kmGXg1oAsEYtE
Es+6SQxPPGKK/QcEA4QSYLfYi6CWYVhMd9bKYhVbI/9Rk9ZxiLkwZHw2Etuj7Uz3
XqaLhB4FFQBfwkbPsD89MlGe704BnLTN8GBd3fp3Ui8voGrLm4G/GbdAL0IFc4mU
5olRnwAPQZOBbrktQkZpPV505344mwuxomqQXic/gRqloZHw8b2LINi4n1YCwH50
NRcyMHcOqW/72qSXk8AnhY4GCcv6sP7vVslMHWu1oyFtXJKNbXE0YoGqCY1Yvk2h
dS9LXUVltnrsCNfseIAH3NE9JR1Hr9RVbzuIPxex8t61MtXn/k7o1+I0MRhiX6xs
CtgGoo0fIhbdaSzkFYDI5nOTpewTyyvEa3xPJOzYOacFxGhEvK5Tp4WXtnZ0CK1v
iAYEJQo5T5lknJqfHRNaTa4WLDmG97X7Z0I6DhA3VoSpIFeHif/0WRHX9pCvNbFi
3wy7dyGJ60CwK7gsfv1hH7fGDYJ3W9stwQuo2QKYybbPyeD6Mlgs17vbXArXoWPj
EvdfkdL4l+pBiD6Cem9asNTdtkmxujhBExfeC6Kc5xbbd3e5yx45lu8r7VSXUGi4
He8iiQz9s7niBybg5kSgTPH3jNU6PGUEeJLEJTJUEDe32ZoE3yLoU4+mNx5PUcIl
eNA8a2LgqGKifivsS0hoeIR/FU4YYQtsY+zfWO+SceO/wngSgSsDCu4EkcwspQ+f
J8N01fTF46WBUH880BjjAgIS+tdFoDGRHjMm3rkBZ9kmtqV+ZqKlh6e9vim+x5b3
DsboFvb+9H8x1V1yNQUL5IYWqLYDVEeEbf5m9DI8Fcw/djkDqVeCHSZOM5kQxYZs
xf6vQdQnJPmD4QimyCrFHzRR8lHOQLiMiyTJ1ZyEJQnkf8XkJygXtja9cFtjpZzO
ge9eWyBHmbzT+7JrG4/+Z9H2PLMVNWWZNWC/5QEeAsFA8/XXDrDQdqbrCM/y+GQp
NhOYkAasR/D75fk1L7vA0xI3jDWybt9HH8CwJKPd8xrEBqQHXHpzTPqc+jrY2k85
+ogTGBYWLwB/8xenjShibD1Vy6qlYK1GyMYH3cTOu0PPv0zq17A2iDo1U/micj2g
7Og1m1plim9CEjZJ7RYVwYjUuKLvBeCJ90Uo+qve9+7Vp+aQKio7s4qq+kHKRxnJ
vsBh+dkHyQvL1l4YALGkm/lyG7eD9dvmNxlmLyCZ/L0QonxnzmB5EL2ZsftK1nYD
OjBqFtkCV73dfyGTTyj/L0zwbmRf2I+lJ1iV7vQ9EDaVM/xuVvGwFGNWwCnmmJGx
PWCjEsXZGrQGCFHXsYmRocfIf1T4AdgfGiDGBbH2LeGKKO08tMK/Q54VoC4ckobc
p8+E2oHv7lKOfenkXm7QdzVKonaBUrFt/m/aBnEgG3syN1s7p3QG9nFlajc+P/eh
d1sHAOA/fzU5fh/v7GCEGrX8iC8KV4YDOgk4lKuEG9RBhi+1KI7Z8Ol+Y8/zTOHx
qkG9F+oFY4XrohFCWSI6YhhCc0pCCxDHTQdLKxEYSO7a103l66wj2b1UR8I6bgLx
`protect END_PROTECTED
