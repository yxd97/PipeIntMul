`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3CRfa1tPW7uYfk0m+OOUACsXtNKbqqeMp4LZ1Tk3Jpxx3ocDOlJv+VhgFHqoLz/c
Xbzjyv6Qyk7TXWg/N4y+zuDj5HcgbAByQT4o5v1aWFE8OgiihX9GYG5kYR5r262c
WGYTHmnBcbIStEk+CccKTUZ3Y+cL/93IC3SX1gDAkgvlL3a5b5RcKfLpdH+3coXw
MU4kZZ28NtEsXFzNtSNOtzAC4etPmNNVG2dX/cR0PDMzVKUXMiXqnokBlv1YJDJk
QtfiOQUEyhFs1a2cu0jypMVZ8xL8rmkQxIo4pHbz9ooBCqcU7mBQuR/QSH6cPIhf
2YEkZ4LcSaPLTuWP0DrmuMrlg0CsmrRDhy9DykvtKWDE5je4UC7j5rrXqtZghH+j
xyM0QTam3MUjW5lIOV4ueyNyEf1YRk8Y8k2u+py4ieEhj4j1IX+G7ny8L9wF1kIs
7TtYxS8QUV5qBmH8jZPYR37x4nrfJBnraHEaxhe2lZj2xlI8KX/bThPVKyXThvpx
KYKqqeSHLIcjIZ8hmssqy3bHgxaP7+08CLNJ5AC5qt5DN2d4xgDwkxM/D3NjyIrJ
3gEGMFAk/8+yVgGlIbUNlpwGJW7axljv8tZxDE9PCb8XTynNIb+ejEqSvFk5jnKt
DLKHTSHGVjAckTLkcP3ucOV7AzzX/lqg9jQJyEl/v4QPJ2313jBztvugRUAEyEy9
ltHtra8Zfr3hIVmdq03Y4hvISJgCjJoahm6z4kba6B0vs7NECN5IQKBxdEA3PQk4
jebgdPP3DhIbMs209QGG93g52eesyigUb3BpRomeaxMYr6Kk9NF+fTpn0ZkukaVd
G76q4Yeq+e7cIOu4Jp6FZRNvB+0VLYa0+lxoj5nXhL33JroKfc7iGPRMYqGxvZ+Z
fR3YSusEQAozCPm+K5EGfQVFjB0gOv7jawvaqHVXF1wMqyhmTB/34IkWyy6wvRbi
ym08NpJDf0gM9yiNNe7Q8kxlH9jrgpUVttbuz9ZcoaXdxunKnrUn9QGRPX7BZl9m
MiKuEAhlMBxgMTLr5LypRUQvHvaBZ5d8t9+F851AOtTFB2PlmyUVM0hdCeY2LVvu
/1vkwytKKTbCNkJIsBLL/ViW1Pd0e0ACyqnPpYvnwp5KRnMY2mLtb9D1C/JTo/K/
NuTjnHoyztAoLKX2D6I+u52x/mHLB8e5buzhyVKjH4F4AfwHsVFoDgrlauS3yn/P
oOAsnMNxVIyWezNpg8EqFC/heKecBkHVJ7H9GcPH2S7pp8gdjodMzD1dfScZZx3c
SB1BtLr9sgGS87WdNJD0inpz3wW8zkZ27YA36ZZmTdyf99oub/BYkMH0xVsj+4qz
olRvoQBQMtqz+rL1IIMEKAmFooHKJvacvQqNp75wggXbG5wg+NT8P1a6IlYwwEyC
EIJmbQyaH4g4PMzG3Bd8Nhd4vr4fWIFrUxmfxYVqxIaVRJ9WTRYqAm84YO4SINlc
HC9bq2GO9nB3mtYz2BHUN4DgxCbyzAPC8xVQ+hKRgTRscyhfZqJhBi1BY7a8niGa
yG4kw0eYpVu1JhNNs+lJj0WDFk8jMfu2tE3mRR+eDW61ru4m0NekOlltwlowM9A2
e3JBCKsTdp5jtgMUZSu7rCzP/1rkai8MLY+NlFoFACllOl8l2tHL0nuSWS9vo3Ol
xNzzigLOBvAyYgCRSCDLmknnsnMdXB7JefIPM6lIG5Yc/4Wein5/vjKGNjIVQXAB
XVdgZ+dnLmNH+CsPe4JzQJm5d+dSBLYCUcqIkOtEAcv1xTp5NpX+CYQiaG1Z+xiB
CV23PpuiZ76zphAPusUAAP045Wp6WnXFmnSWiaHBVgFTpa/p8gZRlAB4nb6Sf0iL
9/BdXPOHYMBZOANDfhb/wLbmu9x5rL0BJW/ECW06qyNrR5nYtXg41dP97997NvdI
heVD+9nY9I96i0aX85mfaze3nyM5Zej7Pta+cxMi4Xkk2p4J6ET0Q41TRSKtBNra
gW50bw2XNPGyadxDj9mTLB8N7cpd++K/alTlFKbCcnGYrP3t9RLVxtj7EI/Vm66N
ghUFxy03V5XzXRnd2mOsbDj2lyn6uyQB02sqYzibF1nTNonNUarF8iXoNNUEGr+5
vpfRox2KGZbuhZeHE9F3NVpncNnikJ2YCtd1aRj29AVgT+ryaU2fmgPCopWBmjhi
C78XKTTdhSWFHzxIzAoQgz38m3LBvOpOwbz+IBP0nBu+GSYYCMhK2wjr4V/dNHJF
e5eqzdd7FqVqIFiNrzg2g9NDCzO77dLAp4GYTJl5oVQ6XYc/Co4Kq8jVs/ghtNbU
JJLEhceUTz0DlJx71dluP+tzosYaIo8Swdi7kEmqCemqx0z2QIPp2jhPkh4D1LKZ
NkDi4Tya8p/O/k/YJFviNCUzY7eU6I3Tur3fdKBOGzW3x4RLUCT5SaaMhgTpKjV3
EDNv5vgu/WLvTbn8/g+CZMmssMcfqGrGOwsT+zBPPXGbSQai4uxyXxyk9uDVu8Y7
`protect END_PROTECTED
