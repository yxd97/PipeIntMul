`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFCtYHFmzEjUMCxphgIWmA7MMBAGizklu0TCrUhw1b0POKtBIgTb7jLdUohyXOD3
Ztb97axOiAJfZH+W07gAYpzybNxvHB57jjX7Pzx7pOd/bAVYQuACAsyYTdQyN68i
76LQ+sXK3FITN2OY5wWf/4gixZHXNCsMzVDnBinIGfo7nTo264V1/kdpi8uqpt8A
80ygHhsPdvjRtp/7oUNzCKOq1b5c5ph7Zy+ctQXn7D5lReiiyMhzSB1Z9T9AP7WK
wJ2W+5n6JVeIzO/EcJDBpxCWxNKJkX0b7MnmrwQpy+h2doVFQOOHxg5smXCjV8jf
n9Y8+QzNoYbRQorN9/YdWzzsmZdgITG/blvCHqzpY+lJSxpMfJ2k2nYomn1OZgPP
TsNiU3oOT2cYu96cH3ylD6+SFGnvKPbx54LpVcJ1rwYBpaucSIjDgIg8tuxUWIgj
1d7PlNgnYPPkArFtlB8WiJAPebjEpc+9TcPIwoRrGBOjIKRgz4awQB/6vwdIeYlv
iUYJT90OPsIKo78XbhMa1nRS6WkbDoPA0V1gvtmmzf8Y6J4E3MmasckL/bCOy6Pg
Zh7NERwR+y+m8AiIi4NQ3ZCjBOTTq6SbsVMhNvYFmaXR6xRnzWRw1i17dpssUN5z
8qa7eIHzUi/FMaQhgmkGZjvlr4LDHi6Gv0f68Z7CVQj4RBDhrCAhhCzrwKGa6z0x
4PPARoIWGSOf2JDf0nIO4hGOBsWP+J3YTls/jLAYxDQ=
`protect END_PROTECTED
