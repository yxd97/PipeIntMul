`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tep6hhK1EfZfReWG/R4J4heuYUKHGHYRe4l+ZXMSARc10W6LKiDfFBfCF+ilW8K9
Qq0LQNPKPsAVNTSW/R8EazXT7n1rUxWTBFPfHikIkAVNWdw5lBfnDUtQ7iK/jIrs
acY+POdIiSesqjZlg28BwgeMi5n9IovxmOq0NoGeVz0D6fcPuzszPR9VRYdf5sXy
AmPgEd5WuQfQgAdI9mt4Dw2p6r3bi9Sg3zkAbz45qlDPaMPKrMpU8vp3+xHvtw44
/S47CJu5431/RRc7hvrIlPjuY7/b/ksxvwkQbV/YqWgkgTFm1iPVyv2Fb/E30ILu
44ROxAd7cKJtldQHzdRqUGkFy5lcG9rKmq80yq1mnwUAkPoOmbu9mnTDKac5kmiQ
/EolTOV5jDsDp5OUJ6wI+3s/nNeyHnpQZ/xeFlWir0ZyLYIuImLYgN5KDqD2MPJ7
4zRcEXtCYMQ96+91S+ItrlhOtCGQNzAc0hL9N/O8j3HRrjn0FXhu8Lqhxirwgtov
RhBRdc0USRl7Ay4D3d8V+HzN1QcSLEaOx5sz+ee0LsrRhCQ/KU3GY6QKg59UUsPf
WGr2g5/oE067keZfkzSS6HKc0dnm0ITY6DqXs+Fh2EbTvF8QqOj9EoB6EQ+DbMhp
3g6Nyc0U4GxjL6GA1AwOndj7ozfArNYMc1t3zqH4xo3sjNbt9C38D88cf9nYijlr
zjDEwU1KPbPfZepC+dhBpsn/ys7/uHj5ENhNKCaWM1nUv4dyKfx8+V/C3y8BzH5x
+qJyLWOkOrdhe58SJ4XUyDZ3vhyjwN0fWeHEIVaLwlQhBotBQmyXMfxOn9WbBGKH
PEe/U4ROd6o+EzkFKo1ljO+AIGl61sNPl7K6uI6z6qwcY8Sf/ccJJwH8OaJ2jc3B
qLT0evJvOdspfFL3KI0EjLSd9TfuY2Sd3fKNbz41FfZ0nNE53ndcnePgG7man2QI
KKdhdMc885TzSq9796iT0Rxt7GXAnTiWZkkG2qBIY6maxGlu0rvJU2LVFjl0A4Im
ft0wNZRm9/kwO5BwUY0jT3ZXY2HfbyZJjISQU+6sxJSvPhv6sXRorK3ScOomaN+c
REGTSfAsU0S9KUegKXj9en4NevWdLs+FCF8VNRcrKem4+KfwyzAz5T4re4v/OdO6
nrfwUxnrMCUAiPlH3MzWWug59frA088i79JZqASwf9oEGZo9anssEiKlwe/wmX0o
5wmWF1yCsDhVu18iYS266OoNrslVbmTb3q1DDeLzTNZyqQhb70vHPH7D8mbPmZ5Z
6Ttd/Ys3sy/9Ud+GQED53kC7pPuChcRESI7yZ5uQOmwt42J+mT9Ic0r7/fqoy7VK
w86fGp0v9HX4c2rQt2ic6NlIl6TfV7/h75Q8X4A+3glUQM4GGH+X9Fj/wBHs0AK/
FeGxXqSD9NhDR6X6Nt1Spnrg6QLeVNLb/euU3sh3JoegY4Cn30Nprf0xB+/t9dy7
3K4iRN/vsLPZ1wz4/w/9ryahlG/NvwT9sTWRyu+LGhno4arzdx57/pxcCMC9wOzL
Z3xUyuj/iRtVBKNEsZStgp+lWP8U9B148GmVRzznq++b5rOgaOjQgYWek+RLvmtd
FeI7y2LLLDI3Z9Ap2gMLxGXwbefz5fyMLYVNUREYmuoGO1KO5IGbOjrd2O36hKpI
WaSwAz8hnqdUk4iD6HWrUI9yV3jcKeuLZSrWQfAghKgOKOBxjMyWW+gziO1ofapi
smcjzH5px6nzHOOvXBvWoUnwe0kw/2eHxr72mt1fiV+pR4NGs6qidnBOI4uyTtNA
czAX+ibCoOh/GrTWJkzNYA/Sy3qyLz5pfPEd7Jz+wRpSKN9BCa+3IpUhya+ZaHGL
oC1A8ITA/S0ocR8sVtNkq7Im4Gm+ebdLt9jzEYllnVtqShzRkKfCE9Tdm+3h246n
z0HrwAwR+kb2Q7vcGjyo73hdkvz0DYHudOQO+NcHxPtv9chqNe4UqFhgPa+zCHpv
tminZ+6J96X7CMSCsdSFRa2S5frDCSxmsA5/oP8NA2I4i0cLqIlXZpqzdtv+bWIB
6IAHuBqJJBuLQGqoy0rgZXaZ1YpwGwzFomsrfMPqBiRPrNlajbap7d8dmwhTAeeu
Ppp+m0IOqB+x637DXEyrBtTDTh7vPqt4xS72qqgWmoZubTgoLgET3k+zIYmiyCX2
J46QD5/5Hm7jBc2Co9Epbn/s+8S0ooRxjexst90ASxLh43kMtkHlY8qhRosiIFgb
J5IWfOoMriljAbaru/JBaAxB0SsrViYopg9piUUuudQFZA0Yt9bsQbjlKisDJtJr
LGCQI8hKPS8k1Wkmlg20Em6KzEE1Crx2eclIKR54kEhkzoqnGk4zLEVHdZb0ZL9a
COEnm9aCE/pDSiQIdxaav8Bso56SeqR8SqvIzIeB+HzeEDGzDgKwC3HJU4zxyjYy
7/w50l486f3dY8/m8qgAiwMtt+PBG/N3oYaZeP5gy99j7TUuLJ5STds6BVdegazH
QvHLY9VcPNngXw7qNWtQ0/0vGhP/IEJL8oqlNBKefyA+oNCRpP1mUdaQ8kVMYlJo
Gn0DLNDwZfaT6AzEs7TrcrlJTlzK9mMkSoHpCPcRBJrB5wtexb+NdvNeFSU0ghDE
HDD4W3JufeJkTkKG3t33cn95M8GNXMWs6vJmPjOaul8UfbdFTZATXqpCe7wJ88J8
7wSjD99yZEK/90i/MCsxHWB7Tp2qHSp26j3rwoKFqLblFhSfiKRSe4hieqs3xYPO
yVmsoGGh6zNDHxbuOOjX5nUY3qBsip8W/CGx52mEY3Rhr7uyL6bvYHgm3f4DRfTb
xVifoqAYPHynReg/w41u/w3E7d+v0S/YxxiYdGilEb8zeNKvfdIIUl7qt2H137sC
rnu1gW2QuCQPAMs4VHTEQrV+9c9HlE0UrZe9rak2ogHKybYg7gKNb2O/fjg3D5+K
n3T9FNdPnxyL4vReXJHl06J6k1nI632PWukpwd2wBRUuizIP38JmmHOFHjgaNMeW
3yDI1x6zjPJ5tCy07FszfmNb0cP7mU6i+gCvu2ykmNHg4xAngMGD9wLVUjlxn8JB
rWDJn7+PXYqO4UQkUZRpv+oS1UkdmK69p924n0DqToOHy57621UC5riNRjRrL82N
FwmbmM7hekz92jMGnle/e4cTeqnP6C6Tggz33m9G7hHuejSDcvTzVM2wW+Mz4VmB
LBqdrL6JkJfkIu0Wc8pTarRvJeEMx5Mu7CyXMCzW+ElOvQi7tcC4WiNxQ3iEUSr9
yzOLGGnfhVTUS6ygxNMU/0Bis+MTywGw2oLzuxYJj18Iz3j52Mkk/Ly1kxmBE4Mp
mBrCZxyPDVqvKmf3EiJn183tkQd7fH1C/PHm853tzOwZsM8CVRN3Vt5/9JU/7BJ+
o5jYLj5YKawaUDsrsADcOGBV5k/2+u9mDJQ2sLH/H9z5XpN0d2I6WFfWudtTNpjs
wYpAsb56nyFSo7yEdkkCavk3cuNq5HQ+xyJ3i2fJSdyOyGT8/I0cW0yIiEHbvuJq
MwDvuEl4rUKdEMW15sfGXIYr3YRNffNXpj6/i6fGgj/ddc+6ZPfsAOuRUV0rgnPK
nsyZSSg4mmlw8Ntvn6mtv2a9SVpmTIPnuKg5w1k90OSTfMdhxyIU7hPkcvkweAGx
bM5OUqevjtQwQQbVZDhDb7k5SBjiI4tCBm7Z2V0BbpJCsKqSGAE/QhKNClO4pAj9
VsGjTWa046f6hpgsED8KNVFvbyM7mcX2skSHzP7b5JHK9yBKvEvjiiBDc6TvGwf/
OovAR845BbWG51Ih1Gi65Ta/VBifmUMCgmcIBlAhTpqy+FSUR0FQ2686PxHpPi/T
fGSAFvLd8wAmD6qAgdReSTHMI1tyQlyQhgD/zrKxMO91HRsWOPFwVzQQH4nWX8fh
y7BN+buimp7+kr7/TyorpruMkaqNv37VzhN15jD/UW5ELzAUbJ8vUuHRPUCYdciO
xsPLH3zIuOBL+CuhhGfsVM4n8cLqrmdTdd+tb0j3Kk4OyVWHdvt4ibs5LInusaK6
rIBt0dJnYc2gOErSKytweO0PFsaAR8wW6eoJ49+p9qNZv8twmCUwdzyvNqBwu6Is
9i7QUhSmZJanImuwaKCUHQpId1VlMccNxCxBQOzsMi9DmUE//FQafTOwVzCFUaYM
kkBXecTHyCCVAZ80uFfVLM2T63bXWfkAT5H2GHxdKGej+/LLvrY1piTefauNXH5Z
+UnBuW8e8zVF8OdwdApBwMuI2l2Yna8brqfT8NSlaXQqp5GTeG+oaOp0gKSsahVW
Y0v2zWh4n8Le/0A/Zso7I1LtONqNsl63lBGUDrlysYKGbJ8WoxBOB6KVq3ShlOjm
0VwQSkLKDqCI4cVYhsv9CBnSVT+fX9cc8smIlZx49mJm4u0B10WclwV8KvBAIVPD
z8j0AaaBSdsqYy4xt4w+/64nfFbzaB5LWmPfyp+/91eBf8/8ezwrqALp9yGejdYO
ZsxTttg4z5XrdFYx0OsD9EwNMORuulaEequzhdS1mgzXh6jk3QEgoLsuvovljY4f
5KiKI7OOQEd0i3fAMlbuQbJ1RBHRda9C4YO0NCZJ3rSFtE1QCTqG3CDLD2M+7F4O
ZSOX0lFhKtXejZO27wIF5FNOis1tktOCVVS/fXl1jgbVMyMLzCaH6ShM/9KnWz1f
qJpBv8AVmIEdI1cKO4tVjjOlXFJ8j4xY2ZR9zBX70FIc0DgJ/QDMufgvpVVhBYNe
S3GO1XnQsW4JHV1m6ei98FLSqcQo/3oXO0XrAutuSuCi4kglLH1hgfK9zH71AkTf
5VzEcBbsVFbPJR+GHKRI21torMD4TtNRK9++MwYjupJmUvf/AXxmJdmhCv1NL6Nm
jfzD6HrryvOiFO7wwvTEddxEj0h2PpHIOU0srNCUubJ0r/35uVZD0/rs1oyP3/s5
9niNAORmquMFdmERviaCzjtQB/zpDyPj2FjXwUdN70el1w5+su0/nGad5M8PavOP
4DfJU93ki0kUrmPMvbQ6QWk/V/92bEqjdL/gFZsKbEagwiIEp19zel3srW5GmEry
zOsdL9DTOnJoPpeZIqLRRvBI46CwaftaO4eVtIz0oswPZ/5KvS5J9W0aZ9TRXKb8
CAr7iGgj2SxddLY2PtpPFSfoJs9paar7rQhOdKuozr46GhqW8hlmwtn1NTdm7wHE
jBb638FGr6F6Xq2D4Vk4RrfV5yCqrqmLcc7Ccgeg+vQ7NgKhxKMj6ee9e/AWJDHF
7UYH4dD4yoyAfY5J+0dE6TBxT/8K8B3MmXf6pTo8OunivPFsWN/pRQrXMpqWs+Cz
r7e0BaTnqDRqwuA0x4miuz7US93NKURFY6s5DJLJ9HFsxzRKIF2zlqWeMBwYf7Tt
6a/CIniJq12NmxEo5HDyfSDrtyaxh5E4qdoht84k1n0vypGJm1AhpkXqM1wpdpXT
qpIpV87MC245FD0z8m+whz3OVaMkFA9hvUwTRJ5pboQBX953qV7jtHsV1+7k9Ewb
Lxs5BL01tgilhbUHG5Of9hrk27ZtvoX0VCO0YNSFN2vXC1xiEkoPB5CbAmXD0LVq
j5zLuZZipgIA0ZtqrJrBhnbBja0FuyXML/5P+x9umxdR8rLzw3Kp9WB+ZX7dmVGC
iZ2o6OdXULUmQsXq0azW+9C3y9Ex5cIlsq5InEkncVnpsrDkCuJ0mQSQbMMr4Zg8
8xlwQHeFp1B7WFT+eHfJc7XDojg/xlOEdsSDZY5Tmmklfz6tGz5kPCvI+2uX4P3R
n1ygVS1KlwuYP5e+JYwHBeP8zHVwfieQ34dom3C5hbzTfEQIxg0V9sFSigRAPryN
cvd4tAt7i9tsUAWx/1y6G1LTdYAXAlu/Cc2FSkL5X+5XWxOlySiA6YwDnL2AmYKB
itMp29O0GUkrrG1Phr87/rcq9RpiWn+F6hYTrAfp8y7D+f7e0VSQK94KrcYrRe3N
8P49OBO75vjdTQW9W+szWOMfsW9mjQsjTHILFpDU0686lowMNQMZZsAC6bt8qBz8
/bBxovL7o/5kjYT65niYBOhywFAh+Twl84+UNhq2PcBHJ/3dg9rYmw3Nqy1SUYmp
6T8XEVKNfCfI+EqjCYWlT0F/BkgzyX5x4UlH/EuI0LNxdSlN9kMeKnfae6Bob2w7
ICMwsxZNObjky6JTaIkHjUWdU5XPiyTsJ8GfsZDWhDMib8x2qx3qYk6m0UzByHCS
nT59JuijO+3ZPIhZiFOAxkZ7TCJ0GbPTZ5zBkb76KAMGEu5dyhQV3JJIVx8JU6Lr
ywits9d8YHx+9SZ2S/5mq8Qm6lP0iNeuIEq4tDgJC61jyTJclZK7R6F57f72W4IW
1r7yfgimKO+R1oXAfcxKcB6rL0iIniGm3L7BP4H7jIoxtZtsE7DRWTTqc9/cViIk
6y5hbhkbxmCBXfHtS+PKzSAdZjdEbmr4C4L79ALOpV87BPTCCn+JMjYW8b7vRODm
NpQeGcaY38MmCtaNCv4da33mrO3IwIGDcYiFAUVJJbXRoVCbLCZ5Gz7RLBlyB3c3
bU4Tn146jd/NnxQBcyzP4D/SzqImEMsZ0WcWuPZ25GqFAGqzn9QjQQwIMK349fQB
iOLbDQsLQXnbQYemevGxQK02AI17riRynVZ/tqLVtXo8tJdms9L0Lw5De1kD3EbC
tmhkc56Ai/WhURPvNPw6U4JvnYQWYHZQ+5Vy9G+hNKLMooQNCBCBD7oHZVBgRAS9
5xEs6vEHG8jcDNFX3PR2KB1F8vj8CQL6Cp4F3LsfIGmsx9TCoxP5/PlCaTh7hWzE
pkzjz2NG72r/0NBEpZ208RpKJh67RqticMTiJTNJz6jMOlqdzjAMnjrW9ka6Gu1i
qglek4l7o2G0ZAJYKMHMrAraDfde8CUYxjjoqbEeIbKduiHHtdcETzgdXS4uBP3R
ENr59cJCWXNVjdywVpK1BUVe5xEysIDmfjAih++RIJS+Wjzghmtpz17VZqPOAGIv
9gO0SM3K0zcFH35YBS5cm7GzTL8W5bUk/+BCdPZ+/m1JwoXCZAJ3IB0pXq3qPiDq
RC/4cfQJCbMO9HmOCLIhKvG+aBmg71I0x4jXHOI5sY9LnRQR/UZN0TePc9zrcgUv
37n+7rC1EAADH4U01ujO2oxxX7ORUziYsLR4az/HRN8FRHKwMHR08krmCmJ+WkhB
b63BJXa+RKwzMpIp3XX37M7IFH5evPCKJlDmsI6zgTOlH8FJNlSswQqKxP1yvCCY
787Xvz1E9w9bljwauU/xfct9Nbin/U0GJzbr7OGt+p4jRRuXTDdKPQVJhm6GzC8r
lij+5qxP9lnOwdZHAE47+KyFVble8Bo0Py1D6R0gV6sy9ZdATB9r7qZCxc0aJD6r
kJVq04ahqx6RBFNxbrPfKlqBmtCBtP+hINGpgbt/NgTUPRABnTP3thFst0WiD/iN
IsO9uz5ExkqliYXLTQ9vZN6flcHR4twrfmyX95VUDs9uzPD0R+4ol2UC7RHhgpI8
8//vRadPy4X/aWd1UxNULDH3bW6RhXw2304LDI7F53wGja7Ntpje1xo1/vQsvOw1
6epxS699CIXQStKkiA/lutFHnJlRBzLr2jcRBsGnLQtLaqgL284qmzEtRa0WvcZX
CneJEqRyunSuxgKP8ZWiJjqE04SjvKR3WASVBjBIMNo/5Mg7qxjSlbJS9v4vRha3
13UcH2PGzTXD4909FIvIe5NSDpLuBkJdEEkPYO91KjV/SBqoB38pIg67PpyQoXPf
xU23hzWSCar4wdE5bn22VO2YWyyplEl3xErKIfYfEorIsqKH/8KzEpJk7SaGZU7G
RIR7XopWX/jV2+H3DBf6IveKtZfvCmdTTh3M+uyO1sCU2/DgZKZUy1hlp7GOaPDL
pXUGsIMOpyYLAP6NQKgt9rmb5c0vEtOzFge7xoV8C5XgFsTzBq9uhUboQwGoTwaR
jSe+D0QYdNW7U8o15XQfqCi0608FJv62Y9M6Fw7V67gkdv6ng8bynGX6/PThZM1s
M7DYnVWuO2tLvvMAt7pQ0E3ruzjxyEnY2Gnz2IR55Smr2Zf2AplhbpgIhD4vbPx9
1v1OeceFvm3UDliJkidLHGUOOwmA/Cuuy97L88wiIFiOScGkbw0aJrzmqmI0+cKZ
+RaH+DMleIMCv1MyizpgyQtwrMDqIRoz00idCy5RWsaJY9aLJ+YczypFpV/ey54L
8UhsqTpzkR9j7sD0TVLUT0uPFeX/bBqifBmWTNzxIeE4jmc20MiqiIch8X2JT2cP
5jdGq2g8WrwqRQwTXe9DwSbV7Wp/lTFDuSxPRFZv13/TAUjEtGRqOd0XSRL5vEdE
cLb0+L9fzphiKutY8jfZ1buM3OZ98EGEaITi9h1YgbdfBQ/D3aPuyz299FgbH6a8
cyxQ7n3EArEvM1O9yl+S8tMkASIkol4g3bN8mRMETk5lkLAB6+rpM+dTRdsyk9px
SFWMWxMbqDBwWzvcejbIlekuxMbBopcZYl8YI/xPUb+rDi+W1OQH8zF1NhE8SYSa
p9r1kMFtqDan6eGTea/NYY578J6IlbeXMo2cMaTluO0v3YIxOpfjbxQVJHemL/gO
QQ5sMXeQb4x1YT42YlMT67hjTc7Fk7vXOxpHdUSfRHH0yvXxzPBFjeTsTMPuBQkm
eyPTP96DAIXatJuEBSA7Nv0fNWseIPB9ZeGS3ehBA3AC8CDp5jPCpiJtlEl0/9hQ
2GSfbPApM1k216q6Qk808kYlYCB4/q7Vy0ntiX4+9u1+neOBKAcJm5Fi7eCy+8IF
VatjO5OJLB3LmWNipUFJgh/F42Zp+/ww6LS3zeFstVjaSmzsRFUZp1vuEqx94W7j
T7B+ooZM5e2kxCKMbY4Q83s58z4GOy+qZQP6ZPh4TqSE5Hgr0pmDJ8RTX/RH1G20
XhgWJz/WTeXikElZ8tkS1e4znUFeSNKQ/B0KjCCl+bFsyBrcVDBfVXyXiOmdCVz0
6vTeU0oD82e3LLUBP0JKMhWkZlCnK+Gkpxs9FeS408awzvp5zLiILyEFCzFXfeZW
qYYB9QHmaSRDuvWLz9sK1oT2RIzp0McTkrygvYcPK+DTmUeZwQsUroyLNvZefF/V
xCmd7xqrGberIzcuGzw6SQ+JbMTaiWKJ+kxDHzgwzGhiY2l0b2MqSF+Jm1lEjDjF
z0W8tN7JggKsXp5codHszx528peFkQOuBYHtVWdueQNFjRzSyYDvtfd9fWRDk5v5
uYR1qYMEodm/n4Se8sAA020SOND8pCf1AJVq3uURJ7fvE9PrPBwGxqtp7jIOgpsL
5H2zfYJIlmmC6JRqO3qsFk9rYMjy4nASY/t8NRVLDvmtnUK2ebHDZhXyAfXFaVyK
KFbPbIyz7HWSmigQ1yeoWIH8IEfQvxznT7sgpR6fhJDSDUFoF3mRKwoe0q8+lVxK
cvGcsN3ydfK6y1qJlI1omJa1wHy0W9x1QsNuitjJzwey9IiOHOWlH8RpdHbxLk20
qwQPioNPXjGxzz/QHtKkCa/MFdxctT4N2vBkIZnnPGeXYFBvWh0uNwg6grQk43JQ
mGgupBRw1j0Q0x6dzHtZNYI+jOMjqjK+gpxSkIoFyM1ydZDNikv8RrJdzybp8I9V
TKYFnTXuDa5EQ9cn681gshBBpXDfvj2deN1BatqbbPrZPP0HVpAGGTfav4pQS8F4
os/CeNVhnwFv8YIMw7GQ7cpyYhaNZv7iD1xvlqnvtzZkz9ouWG/2k6NL65GCuzAG
P2u2KorevaqIkzTujdcp5p7WHJLZMn1jpbqNffvtihI1j/GQPbxYk4PUEGZmzNZ/
SXxxmSYwL2Os2DVt78p0XzSUVuOH9U3m6B7q/HajWFM5D/27VWtduXrTD4m23Shl
pyTyUURq1T52VGTcXrA/8Pe/vP+k55bUQo8d7Veo92k0m8a2/Ea4QPe0+KnaIlqM
Yopy4nwZ1Nh10twDmWcRROPCHcyctcLiKDlrHymZlQLlTNFid7orNkxto330scFU
IN4BwukR0MSI/iO5CbMqNCF2t45EZxu8OvMl5IJfcjjtGJxdX8EqXSfQdYcNKYdP
RcX7CzI8vpDPIR0YimxQ8u507AOnfG0m6LcjCSoflOkL4Xq1PudmMwJvgEgPTNV1
DHW634+4WiFkUHh2NAzCiFrBAGJzr6HPw7m61oRENLuub99HBaWK05Xknx9Kngbq
Q6YA92CLfagN79IwFiQR9yVIQtRDVYCPRkkltp0wbt5GAId0ZiVRyQRsLwaZMy89
83ksISJOKce5NdAjcx3I1ORRu2b2qYfQEKWUrV/dkNqYDvDL/MrJpx1aJ/0OvhbU
aUXaUwxtHJjN5K0cthL4I98AMOY9NLLiMLRYWWvMuwWXiUorh3x7ZYjEtyVoMTbA
qReB4TGeeqhDagqChX+2g08XA4Fpinhs0fWpcijlcel8xbcvVaeVlDV9WZt7pldw
qSXVYQUCSatWJH0Te97aR+sZXP1yXEKf2gxPW1kf5y86C3Jr5aa1QR5csddHpOcw
7OeB60tD/9UU78BEq2/Tcb3c4wCrZD5V4RD5LpCTerTsnU6aaVeDgfcu34qFhL6N
RALF3ML/e/FF8pRQQhbBSihkHs0+pPsvfZF0HTl4jg6dVRwc9p+UcVQc1oBdJtWJ
6ddHVQuS11eyBr9315eytk5dDbuStXUIm5CD/AALHaKAd06zOiT6+Sa1NaROALLD
buGYkKUyt/x2XH2E748UpRwu1bbQf33Yqlslm8ioiziYJzSxCXp7MDfcvnsMDla0
rJ8hLhZkMErnUNuyg6QYaro/aZvPcMwwkM7qMQBQPahm48RbMl4eRi5e/JKQ+Z5H
7VtqVlLUoDATdtptcRRAbHFa4hqxEGIWP/zbGC0pSTrK+IX7+TCNa9yb0ntWDhmr
lboQovn55o1nmQChPMzAIjk/vVK13Wt038FwANVKecG+GLKS2qT5WDukRn8hNope
7F7GelS2Crr6eQDl7UErDEpPZQsUFE552SqnZJi7o/TVo8WjIw1UzkMpBWFz29mH
vN0J8IYEDzHj3Gn+zS6GuDPMP0Oh14HsjDEDKXIF6mSMmcg792JaXml9yaLcWszo
ZsifNZCtRMblFTQ0px1/w/tZeAQYvVhlowVi8HRVFcPt3lQksd8fJynb09NPSu2W
FzGETDkznD59ajtUlJCxiQHxEEXP8z7niTlegrZElL3dRBRXhL5AMU3dBJV4X1AF
8gB9hxzUxpacZ6IDtD7mfobDbuOqmhLnh6G+slFtToUECT46yvlQ04kO2vA6ab1c
t9s5F+UzXgx64PRgUHZ/ieIySuZtxIwOjnD2X5Pctybc6970Sm9bO0QWXreEHmJb
JCHmoSu396CzDz0BjYt/NR+Zl3HIUMAsjr+y4rCrmty44xhpjxU3B4+sUa6f2eco
zLU3cLYT2DEU09nqvxP1/V793pGY3wBwfX2oNbiFX95Cewsu2dVNyMFyCsLziwPt
Izvm28Jj3DIiUmngz22XNO4u0hRI0oN7u+VUqA66hsJngXK3BFIeYpMsWUIbYu4y
m+Nt8BfQDtD7P08pUq5hmnmqmvEeKqOK9qOvwXjvjtkrPUvRFce/0HJMQpZEikUi
g8FLsgPAZzLZgSRZgFUZlOG0eWfApjLlp46pdXnJLcOEVPAnrCn64h3XUo1AWWJT
i6g3f4qJgLuxls2D4p+1KKgfNuF/VE5QZ/DkPK4BW5CP0ynMHif3pFk9jC3TOiCP
ls8QDZMAFQZH9T6hC6i37qYOaqPhG7X2PrQqmJySWWGGVBgNrhPKdZVDblZODPMS
4VtqyBqmo/GCwbbSVVsWhzNG2kzpbVQquUT0BWQirSWpCapXdIvrtH9jKn7pze+a
RJpKxWQF0eGQkqyGay86k1QlrhMzhVb3mjseFEz4E+xNfcCw8k2pvD/G6EKek0G1
SsfN0kH1NnoxBnSJKx5Jb0q25qwHsiyuo2aauM1Q8Ab2dPoFG6r3wXrApXVLQh7V
NbcH85qsyImKOTZq8dMYMQeEe4Rh39TIaihOzOb0uhO22GrXxx6Q8zxKYrIxhg26
/lUU8Sr96kJrwAhFoI41mBnYWOVfUzeGlIENBYxGo+gbKPYVSfk7JA3ugIl23Dac
q9e0thSZRD2rFJReDMYyDWmiLdVGkSjtu8rS5MZ2ObiJiyqGQZjW605cNXbAy/at
wb2N3ZfvPGVgJJpfTUnTfRCC8728S34YUM/NxYiKPEadaN2wFAeNTQ/W0+LNXA8t
CU87I/0M0SSbLTQJlrM+ltjDpQp3dq4b2KW6WUjRbTyPR8e4U8ewQZAOByN6lTGp
a6rm4/n8gmA/80mjwFjGWJcbkbD5IbUW5gBw2VQBhhaGKeSmZYk432GZ9rYFAkq2
o/VUpvCf+hpC8c1DA4eztQaq+MFt33Y5KZ3nwgiG7B3RIkS1+o1SaWooyb6yroXp
UxNzd6YUZTYyOxVEzaNWyd0cZhmYZBBjQWIRUCfOMS16F9tCIpLKUA1SPkbGfgoU
xfTzGdisFJm9yc2+TK1XgfL3bKLtauaMMTCWJf9bY6ernKZ+45BbRGhmjRH8GVoX
mzfvkg7EBE1l/sRHj1fRbvVm1PyPdGgPbf379huwdD3PK9JOSxU8qb7qRGTbVlkj
yQdRKMYESXY5a4qa8GrciPqc6fon3wCxQRhS+s/+E3ET2tOoSWEZzyAjp9z3fCgG
98QsIfeEnl/hU4TlEhcW6NpX1UeftJUtqRDv3uyF036Xq8xT1++eXBw64DrasWCm
qzhGMRJJFOHW6+3lnZ4rBpn1sa7CPT5IueiCw7XIP1TG/Ae4PmjWunk0wNMqckBA
9vuno9a8VKMgdR3rT3dMPl5GOYVVZsQE4R92uswGkrcpq5n9mB0J2CKoSN3L/VXI
QWlG+BvRo8UiubXg9WKTjTXRPDArsarA04LFcOjGaXXBtLgDU5i5EODPfDHv+uTJ
vw8UJWayKwhAZ/Lgv7kuDhxd4ub3SkGeQujPJYx0run526iAFfonLsOySQKyQ4I/
X4go4AqQtTfi24nL5ljvV5j46NTOUoy8mOAW1gDCYEDCO0xQpfs0V8dSSqz9Uj21
SztBm9N2rwItdrDSgVouVoyeuZJwAG47xqR81ywkILnrBgtUVDzh6iGHIgn1wduC
xDzdBkUEitM9UirPH9zZjhriTi5VW6cx6arHVBCruvIzRsMEiYgpZ2+q+TbPy8Pf
tRmmNiGkYZHIT02V26Dozhpr/WRC/nVAnr97nl2pcIyzvEKm9lv5cGcwDU7L7KRb
8/G+P+wEo51daKmUmnDkvG3EBEF4acl9fmDKLP0TniDyy4gqIy7HJqH4E6CAJ0M2
porrntVcjZj3soBf4cImvdkXjJX8aFvMF0aQAJ/M8FgGEnbhCgiafMtULX2PIx1H
ntVWVm4Y2zV/mOZW0kZs6pXezWd6tOs567Ga039jdRkcv6e7P/1XOJ3MPhG3DnR5
zvq/e4A1gtNFMiLOHX4oDPUKuNR++glD7KIXmi9uh6RmDk6EmMwdLTcR3bzn5D/l
7w7DyR+xWRvRs7NPQ5tbJXlaXzrTr/334Y4mZk58NWNbkCzk70Uklb4973K3p5tT
ZhuGQwSyx/0bbC/Q2bVF/vJkJLf3qDK9XJiY8dRvYrXMRgues+RuJMekEq15Cxn5
laWTijmRwpts2o0eYN55AuxNs9ap5B/Iw9K0P95UMdrPa2KCQPYPS/43ql0YPdAU
0ncqIbtc2JY3+C0VILTzP295fK8NDdUnq0F5M3f4s07bLCDZisKfy/K8xNX88R2M
k8RC/776tBy409N8Xz3VYDtbqH1oQDomxAr7dTmpDOk5Wv7F22hcyjVon9/2uwUc
zlN+lULSRytJ1e9NBb7EVpf1ywDG4acOAHYvIovJRUUK5jRgCJNA4FBzyg9ai4df
1HilBzOtyA8RLSQlPnJrQslNYTud4UBrqfNAJzqQjozJ+y2Sr9PxWDaJvdh53yKB
dq6d/Nnj02gfWkB3NDUWXmWZ4jD+/GkH1tmv0y2nGWfy3hpx+lW7E+qJNFQg+TxH
izFNY9d0Ncx7GuSSnvIx5fguwFQFXifUx8wVgwge7iInk323TJz8QlSiINYx6BQQ
BAfR7bteY9S9FCT+80Mwq/NGIjS6gT2233QqE4+2iolFYUYUiQubPJPwaKJOZ5SK
gbzeGaIpMJbU0QZ08iIH81wp1M0aPnaljSx3PJTloWW5dcay1KMcsxXoj68lL9E0
xI6K7yOq649LlNTUeBGqY3KKD7BsB9kNFtPsV1Qa7uTSdR17lu7k/XLd57G4W7/X
P2xFXjMPsb850PrB5IF2hAq8vfy1vaxWQmxWp7voafj6XJ23qB1KZdDR989sjA4U
c3hbqZw0mMUTNEGHKQ4Wu8VX/Qnk6P1is4SO9Caak5BVYdMD0o0mPZRpJKASVbAI
hijWgQthrCStOw77hImR6T+BcarDEHKWhIWyaKN/pdCzNEByxEdav6LUX2DdTjgz
wx7G+gWu9VCYsHJkC3WFReZnstS+GVlIINfVw3HyG83xpX3WdzEkw4Y+uDJ4HsOR
TM7F/w1TJLAMXLlk/gZSLGUW2eGqsWZPeELlMf87CzY16TamDhdaoe30IhYAU+Wh
cHituFdWe2Zq6niJWxu7K1zw87iieK2KVI0W3LI+UEtmin/2KnhgJ7yEwMnzPIQ6
dJBAgfmH+2WagarqR2l3fG/8w88cLyNU39xnObfZivpgvIDqggGDeD8MN8B2QRYF
rlKzgpiPUiMqHDtChzarId3/X5ZACef0hz8+I5OpkPRsF43FWazI4wnp2UpNIYlE
grmWpNUyPShSUmrAO0MPSkF4aszhC9zvilqpxie5ftbXpnbA3ttPOyx9OEDinpL6
1sfVDFlE3h+HwAlji6P/i4brVqtrv8e5d8yPG+YpFbdmZpwPsX2nfGrv3mNuGP4F
aEeP3cuPZof4G8L09ld3XyvixoXkBXSp+GpjAtHUTbWmmm6fQpjTI6Dtgwv314a4
ftgUHKNGDtKvgJQbJijpwAkFXYt0E6QwIvmYhTMhGHf/9MG/MTM4wjdDpOKHti7a
cqtqEUwlBqUn+7xQZsXqH6B4HAoWQVHSoDlST4hUSdgc2Bhk5FP/+pd6fLbQR4h2
SBdhS4I1j9l+MKqZCtW/XqrbrSGhAKZoJHlKGTi9ibZXAT4NwRfj5LWfmB2nOp02
e/ofRiaEHJVi0tt45jKsD+puDCmcnvDH+en48nY5AFW4l/O4x3Olghx00sGq4Yvh
33q2TyIM1PKTD9gzppFnDSbEJYTmGm4b3ZEWJpMak+0lm6ktsBAJ8Ns6vaVzRXY9
E7qO+lVJM9LKsf0ZQuuIANd6+d5ZGXvZBam7MUwhUe+wsxChWIYTNifvNHLGpeaY
sgVxUx3kndmrVmRukEvqsJJ0MmjTffQNQT5XG7nXaoRNewJz4ch64u+BM0Ymsqq6
czeEusSCzZ94QKSv8f3HLkgPDIca9IfI+KVWZYcw8/qg+KbAV54VEIvGEW3HsBXm
DaGGT/NnfOmrgMaF1iZlRtynazvfRdXW/v4nZEOL0tniUyTCJ1MkDVN3v9ijvZAm
rBT1YxjBCoxUggucpAFdedRL8wK6zR7tU25MByDG08EpHtkEEOIGSkDaealuTuPb
32FfVjv0rjoFtHLA2DMUSeBswKe6TFPzJv7RskF4GoWPPUnCg4H1YqRzi32IarwB
CjP2HX7F3I+4CYH/IHks6xt2/0/z+P+cFYmWhukcSYpx3bSc0wONUv+EWYuF4qjx
XUfMCDcWDtozZwvxcUNtLHvR+SiYv94le1JV7I/Kdgqm1sCPcNi2QxD52IozCmWo
YtwLXYQydZXQcISYGxqsDa4m/jF2EIRcNBjHmAZ51cTtd/Z13MFK8svor6o4/uV0
FjZFTfEeJTcg6OYEvv97Vf00m+Q/h7InJrusJjiEP8RzLdzLnJrbiVdjGEIC3mJh
7qbDJ6LaLQ9yvX0gKWS3JJ8aQ+8/GLJ1jRdwmExfxImhEdYMZh6hSz4TDC51FSQr
nov4zWFOvxaahgeTuhA2uPKYJbhVabpQaloPOeFtpWLeWYrwTOeVqUsmjTDtB+kT
VNAlXpM3SKrcHhe6DaY/oBrGTepHKO2198+Jd72Iy5rtWrctgHr24pxKlmT5DLGw
XFvKo8OrVapHnZSCcodMtHePYCAc+VDz+3hlrNWKJOC70bxpU6um5sZk6PiA9o1k
5jChAp4ET39kJykpKLuolMLQCyjXPtng1/CKkszDP127jXh8EdTfFM54Dbegk++D
9qHPTlBj2AynEnTwQU2FBmGndIetHkgc6FauvFaixvG1++oc4R6DPqLmCyssbijl
07T4fd77SNTkCjM85S3fU7U3gP2+AFfei7SS6UVaRu/cMB+9rk6lrUj1N+zMMcs1
l7qWA4zqoCpOOjFvEtkh6cpmBNEaU+Fjul+Vfi0u9CAAVYP7LCcrs/WWMboNmWj+
XPUCxmSp5Qv2AF2dBhitUBqGh/J8mk2pNbyr3wAA0jUKa875KYx50NrPEWfpeq5D
ZQwBmWP0xqrnqlE0GuQ1E5XwWOEPmrChSk+FDo1NZsGuM4/qqf5Hp00n9eDr6dOC
YzM9UF9pKV81m+8oJBxGTK989Z0eS6XG9X+1WCRF/R9Yy/aXMN2FNovVBnXqLjV0
2dhuWolcfOhmRnXLR6qucn4aFVs3/+ifyUB9bpMKpCUjSzgITE3ecfIm3llVsOgN
Aa5DK3UhQ8MckkQmj0kxgve1PYqAxbiuVesW1E/byQ2NKw0t1p2mVRNqhfLcAdGp
O7PL7Lxqn0wLUtEhCOgwsyr6dTBmA8V7NJXf2eHLMQp7idoEPmSQ77pnMBHUJl3S
OSZtW3Xhc8zKicBEcG/DdrkhWJJw95KBSHf921hiU+26utBwePglDwHnrVq49VI7
IVMUVeDnZi6PfI62WlEft1OYHq/KbGPSl081lUS4u4oMruEgFJVnT4YKhvI2YukE
m2ehxk9mzcw7SZ17H0q5SY9TQ4dUClzK4EGakui4OeISNvxdKdelakW+8HxMqdSD
SZmPpIY0p8tVHlrIFfbLTBCrmVwOswkbAeS+VNV2M0wMH1FD03gjst00TM+q3oa8
aGsAdKFaHagWf4Cv24BK8LwjufoNomYcKONTDFBSo4xhMx2Kf+x/vXeIbw42XTTm
R8hyZrmIfjtzfaCULx8903q+eaHpr31D9QBlpBb8nny2h9vs6sp+Gb0hk+9sDLvE
Xl7se1T7Fg97+G6H2Gt6p/wKwekDoSjOsp4UCnQY8vLT+Ap5e6CZkmm6pt0csJ2b
yClCxSqARwbds/wG5cTAFRVM/HrmkZ3ROCE480qY2w24Zpt/G2f6n/fibmuIDDCh
9YwSgeHQVoixszIXNi43ju4nvfT5/BfByAaq335Oh1wxCORGymqp0mWMuxzPkX3n
RloHUVnVJCOp7o1Dqp29CKmEQSKHzvzrUsXdED7NBgvR6seq9Hc+axiVYvLlexhG
1aL0KO1rFqK9d+UG7DHi4Wtc3qcKn+b/B3XY7ZsTe69AFIyBZlgTdu8SfvzRe8HO
i4024IvVZ43oz/qwpP+1KXc7QdVwY0p03UMKIrSfSp/75MGcrZsHVwm0I/WVaKUs
rp7SjgRcup6BP4lmwYwwCRyBpD949i3jzMYwVbQDLyiRytDlQnw6iLX/nkNQcrkQ
lTe5iUBk66EdmDPp+Trjmg+93to5Ms+Jx8aaLCOdlgNAPV1Xcub9spd+8RRt+5wW
CTXejgcHz4E4mnCDf8jHmE6pmbHiIdDY4Gkm6pZ8YXepbGyyOnhvQfWSTIcFDd2A
5Zhhr2u1fO3sPaihiaAcDkEtVV1wPGtgbmfzomSAHcafQW/rPTsX4yqtxhKrYxIP
9CTEH7+VhIxz3IL8lbe8qYNqaQY2fbR9zIvEH2wiNEDJz9khyV4yD48HuXd6lc4T
pprcGAXC/6t2/dYVV0v5g319JMnkVGMTCqcdVUl4zzAp2oGPayyA3DHm+XmSw3iy
4iweO67cqUB+OoQ3j0eBM0FlPO8RTB5WJFDQnZJJ3hkS+LD+odq6HZ9ZXB87nT03
32ja0MHMWrv6v4pVWhXi/150QcF2ddcZ5eb/BzVF2dhU87r2enaAg5+IBYK+c2nj
Cl/xTaiU3XYugYGzPFVZzFPRy13UeYuP1zU2pyR3KGemlX3DlLUWuRnGL/MulmnM
75PtH6anG3fnAOIn2EsKRqWNma19HkebI/2buZ7zGD6Z7PnEp0PJy0Yh51LwGq8V
G/M0G7OHyg3MFGBWi/df4goKQ1D4Qlv1EtEVrT0UdF6rBPkMKHAQ5Q3Z/qjX49TX
MYTSehr+w7J+Kkeak2rJJB90o1uRrJuyBOsavZa7gyfCOUqOzhxWHR+2q+UIfJp4
qx2IfIBRNb+wWDhYTX9SJWB79tgwB+W47m4M+7s3wpk1jr064Je+D+2lMKquhuLc
M5qac097u83cOGhTzG94mTXbAz+sVkoCSUWdMGNCTZ2XTv/HX3B5+UuA75ji7wv2
SLfNoz9/Z0N2+HLX33WJGGhtkVAGmme7UOOojvFES3lc9nhjBau6KCfdDrjCyRNv
FlsQslxM4HkfZV8R4z0hFhs+XSaS1JSaZBUUXlObYs5ONS7LcRb8EAv2tfjzg/e7
h/YDgGZBZwtCJgzcOnhfXZT7PNr4WCBi/oxGqohO+gURN1AqzCzvAjBWxoCaaeMP
5FVq2wrx5sKELKHfmdS2mrcGC3KpACrZ4j6UbN/Nsp8gSpXLkKBKSNNQ2EjGegip
RlYFRPQ8iFw6ORo5hRtA2skLc+8bby1F0tUxZrS16WPIyS5+M0s1Gmkcp3MbBM03
zceFSQ9dKegpV0LYLjYNgeho9Kj7v/6qTlJen2fan08xR0jQZk9H601YsdG7UCAF
BUo+vEUJiN5zlToPTOleQZEhYeyT3XtKhTIxwfhEZWLNvPuK3Yg6+3zLnmk6ByR0
fhQQsZ9jQkWHxuW+QfwRoOCY67BDEDeffTW61si0fmqMRHpTpUrxBkAwHn9P+DDG
mh37habI2IP9c0EufZVwCIeawgbPBQc5ipfCXr93RSGNPj/CLQm8Xz8hJ98nRPbb
wWasC+Obb4sgpquMnYD0ZdcCl1R610HIr0ukNb7wzwETS1gp+kse4trsJJ742m9D
Vn4W7Dyge3R2OOpRSWtPx2dVlKxnwCYViKZO16MwYFVwyL2hPNGJ49agaQ03imiY
r0EcoI91Jt4FvK8Umgd01c0L2H7VGhqhNPqGNwVIRmE8J97R7KMNEgY3rpRFPk9R
8wJ5EsoLJYr8i6wtxko8eCYTHuhpRtzjjFpNw4uj/NRHIo2qFZMPuekGgdY0/PPM
aSWM5UqfiYFtRGPclADZ+ooDHn8PImIs9FtNam3iGVSOdcArWkyD7Fcd9ftL2k5L
RjQOsLkUg9Ju1KBKBo2ydsOWVt0wYjK83J7/+q4XA55cUAa3LdqoV6hddEaOW0yf
fTh9hgfkO9BOm9KUy5b/V6Ssv5i8iaW9wxnVNSK2qClwQBfAw2v8j/EJCwuYkj0i
YvDvzzkHp7NV5TKTlbAG4zEh7ma23mFa+ZE158u7wQeb38CvFwLhoPKSJ9S9qJrE
6y0LM68ow7nQ2LqhlY+nIGvcckolGVpj2TpTvMOkLDz8I/50onEp4J3Y8z79V3NI
vQbr14ib7IrIx+PBBOPITqtmxQ9K71iRlEsPz0crvCn9kCMOaOBTz1JJqcfsFWWx
KQLKN9vza6VvJ8dW4BtP1O12zJxk41KaZA0MCwJLBE7L/NJbFFMOjw3yzgBItqyN
1dFWcZIWdcgMDhnF2vYQGj7ZRcN5NrT7NlaQdYu9LEq8g8pWYWNWR5V2UbdlQ2ic
vlHdy1++geqRmbOiNGLpFuxxUSSbSXE1VO7tqS7M6wc2wO0UHfV1lKTeU0g9ik2P
AFtTmkYHQeKg3leinAYnY7yQ2iBxcZFbmQ+Aw+P+wh9b2s/DWWCnE8aTYguININq
YeWIUkcbpGYlGg8sbkWWvaNdGSA9vSk1wHU/AX77yWZJerNjzUQVFbDS7IRX9vGb
w/ilmYcxrWMPPFoHZhbf/kZyJ4uolG6L9IYVYgfYjoptFWHJYod5zZJ50zu7yat2
fjndydXjImLJ5L2d4LObstFPIlXuQD4r20Ju1Au62qvUv1NYyhWXSramuY3VXwJp
0SBC2H+pK8Yaa29KQNG/LwpnnOtGCmK3Rrm+4dv8TObDjWMOABCx+soANMCERtsR
oCRuvjAbqTgZ7YxOece4jPCH0lH1GmGt+qq6lfstx6qGJNuL7a1sqXVMoSdOLBEr
LAIe+46Vy5C0VIkirZYv2W1uDnrtRmjPzZiPqbXjxgx4vdWLejaLWyq9qSK+4SXP
rWDY6mwPGKyyomAURMkJ6alG924NJ/mwI9KbPYBnJ2NDHvBz1i9JL7gCd3SgSKMR
BQ0CzzZC4Lkbkv6Ffdt7kbXoPr86EgFjarfQp+OUrLx+y0V/HRCUU1LqswxcCWIR
HV9HfT4+Qh6a7yC3QvRctxt4+1A70WxuBR04wRPevlxT7zX/G/0p3G4QZpdQ+E9r
72ypiGPTC3Yy9nbewNSW3mOSpqTA50/Mu7ILzroap9pFB8UwYHGv9/hNz7/Bv4wN
odoMUBvZhVJbS6WOTbobCCLoSQvQizxOb0iTa2br3OqGh9+hj9iVNGNfN58PnkR8
fxJWT63ER87pIURvpJtcRvI0LqK+K9S4/w1HirQDl8269PQXRoKkcNLQtCwMGMG7
UiFdY9ZXf3bGI7YRd/dPQDl52jHh4T9K58FcSWBry+tXy7fyhVqqnU5oESENBXCi
zhzpVzdz1fEF87B+iZAM0naS2pt23q9fQVMPxMV0ZipeNLifw0Wmp1Kq/je9HE5T
kJkymhRLaUg/zJayal29cWWlxp+DiPCWJ6hjQjUrVjsNpYRpP1h69I4nqVQO365i
rXUkh76t9OeDLaumFuyaxRzJ3fTkO1v582H71MoJKD3p/hg3VvdoScTSba7s5Lum
yzoQLuD8R8fpdOs1fK0uQ3bhG1Io8tPqHWYh9FhEIOigavIavDOKzdhe7kZI6IdA
P6ob7QMPseNZ0JH0noBVPB486FZrpCpYXljRTNspJ8SMxfOnEeM+NgL2SesUAz3R
dPqaWcAcsw5qnDLquNAKSnlTBPfq3TCNkxeALdJ+oO5kHvSikNYJvU6TFLCbqR7j
aXwEFREFfwLvI/pRfhOzCmaXfWh04oDaq94QO+WxrYVF/muLSMD7CQB2DeepHwUe
T1SQo9YADdhmHnkak938NJOqNKe01kJ7IlfuUNlC333cQ3IHD0UlD/OFqYzwtxe8
s76QqTYOvEHQamAD6fDlZWdP+gFWaSQzIUr2uQP5hdGZtK4zacTU5qOsM+ehmtoS
o19VXsHU6SIkbwW0VQ8Vq+fzbmCca430vLqYhAdby3A7KmEeJPz5Thv51EKopTla
kgkvEnZvRq4CZaGPMBx1+lLdl0c88KzoiPVJuVBOmosgd69o4DdW92u3OOdzxqlh
dRHJYNL5gMiNLfnuO+y2gROClK5WoQkH+Ekc3jILczwOu375UM9jSDa7fRvfael3
3klHsoxYdWfPf6upcmAnPHBZTcJ8EPzmFlAfQU6QQ5cl+2Rm8eMaXTH8DhiCjyo4
ca0mdcZUtwD91Us2KtBWCmBtd+QHpjPEenIhRbdYmySIlZ49RC9cgu5diBLTiwzw
yjDo+ZxCEDe/vIq6cLCoiwkA4EJ2dVaHc6nFGQqaXt10v+WEkYFvkiG80FSe1Zsv
IZzZS+eR1PyuSUy7dMRWzq/qJg16EmxsJIBK+/cFiYpFFOAsdXbsFOvzayPDgSE9
oA9voiC6SmFKYwZSOgn3wgLMvJMPd/zJZzKNQAsg0Ai2mgIP7bUX3Lt2rLuKdZaz
r/rmOseeyyLDuC6Ny7xYKTP+bX/fR6QJFrq6Iz5WqtPUWCoMF7HKhtiJev8QcZVI
qRk4q+koR6w2fqlN2Z1dqVgITk5XCujZve5TKkiSGKeqcZ5GWpSWeyLmB9GPwZHb
XxbQt53I5F20pJch02+j7Dpa39a9P2sSA9LXGdVca1XVf1GwX2c4Tz3hWlx/OSvY
RGHNi6IcpotJ2cDEscoZetsayAGij0qwGJPRZFkna4u2MJ+d3zO8yfxJ2lZrWak2
dDdpyuXuDnqSP5cjCfrePML0V8LIdqYNWINFThu9+BEE653SagRBfnzi6xa4YzGt
X4kSiDxHriDT7jaziXED9nNwN91qqth09cWtuEPh/KLnS5g0F5Hns+d3JLqjGbn0
Yz8TH2qXzOnk3kpd5FYbMRFH9y8vHIFyjjm0VxVf71/E9CLL7qItfqPdy83Ued+F
9BNwVcibCSBDaQq2236N3DEyB+FlL1TDTDXX+NGFJWrvAnvyPX8SCtg7xh/kSvhi
t/Ao3GZhamNUupsyOShqZRVQ/1ctbsOQO3Ck/SPzeEfwnLcmy/+CZjhd19jmmbgy
FFYwXyTuQmEKOH7DlLIXsZOZaTXP+qNL4DFn+koEYQhlLSWD+NFt7wjNSkZBOPYH
wlHkkJUl01GEK9t5VxCEF29Ftu+AFKT+2qRiZslukc2AYnNuXgS6PRgt9+bKnJ6R
s9OcLZ8o+ozRxjmQIrdRTFg9bjb2+5UD0AVKLMg4GIqVdmsRMDOmPHz95pt/iLSQ
EqhIc/6C+MeOC7OAgm41IonSn6Z70gARMYhM5pP6rF8313cskrEWxWxwwrajlIoK
XSMhLzuXCA1tPtp9OQY3FNSrlg35X1zINxgJJY9m6i6aP0MP/PQ0iTSk3pUPz8wH
OHc7XqlJPw9sXMk3ZBXMxSFvYvWqKL/OlhafMDAfNhi/eYrQLNKrkxKMHqWg5TCQ
jgLdOCsbrsKs25UM7sNVk/r11EYaIeMm9JwBTEnGRy7CDG7xBxU1vK1wC0GAI9Uq
DM2xv3ViSCar974dPx2XEMRDrlPtA9hfLx6L2NH/tyDwXjQhLudaVQMuxwzCT1YG
tvCx5w1D0f9R8y5C2kV7U271YhfmYYNS8wQj7mMlaKe8hKAWJtoANVQVgQzb2AU5
abuucVRg1TGvN2AtLD9i2S9XiRtExud0LZ4xMukKezBGqWwV6tHROyhIn1uLL7rw
T2L4afxaKW42JXrIXFuX67L0zFHe0XMqanYfpcfVb+lwU1igJ1gwaowszd1LmCP4
gWDQr7PvY8K40Y6vnIEwyh5iBlC03PXGM9x8y2+GpC56JaFXTfsMCuRbb/YLL/VB
uJweHG3t37kzn1sEtKS+nKElau7qvYssICDLl9Qpgztnp4xZPg5gpxV1sAsDqQN3
r6fNMdhruX7nx/vKqcKP8pX+Ib0rQc+lMR7tIgryZIw8b09HYm5OSDGrS08H9Syg
DTrIWetC5wdP6Q/jEEqk9aQTyaLmF+vkYG2QOtP0toV7LqZ7ob4pnbkn6pmv1VqQ
OobXVZ5FS1CqY/Gp2JViNkLmCqr9YIyaAdN+04M8ulrxspS7Gu/d84wk/wNbfkpx
Spz6Tl1S3JNDyL6Z2OMZupujSXfElJGJsmLSATl83kVXt5CWrHVvPIHbDbv6ZHRo
7SYYsbl+ysPHoWImiqUtPSnzpXZvXNaxkeiuditZpRFXUAWKbyE6kf911rozop7S
YnvV9KpNjCnE86mB7/4BS0VSlk0B9OWqVmSnEhuoJio5zA3sWOXpxM6GLB6FL1+P
9X+ZKXkoDlCZ39zWmKcNJd8HHMW3Nu/t/idlspxecH/DL7FDs40ODvpHBngslt4T
Ou4ODtI105EcgKuu3R16I8fC65vW3riA/PIdUyaOOpMLfHi1qsUEfKKNbGVCI0KH
poSZKFUyVSERKrpraw4ribba9xQhYS9ItBw4dRtG5TzJOk+ucIddlc5qGEdjA2Dy
P03dlyhF5S4h69xqX2g40fpYVM2UUk5xbMP6TyrUm6gmvYvthe1yv/MfyqSyWYK6
mnAGU93S8t8yQ6BAcbRb0yqQPzBL6kca4ntn8A9rGb8mp1XLOeBmzHVPGL/S16i6
4qpmuVJHYi1+QCADEkfsIWz0QkOM/f3hPMFHmNPMJM/6tvUVGfvynXHkGC4eRZpN
tleZ/WBu5j18K1j9XJwhmEoIUuqOUbD1LNEm95XVLAHZRNMYAxRIOyNj1LE7KpWn
Hd4Ghp7TOt39WcDYEHqoRpFEc36uFFZXesZwtkZO4TMWVxvVbrq8Wg3OwnT0DDCs
1umLfuqZ2RtFr8zaZKLNR5mK/piCF7EQrX8msGqzGcWT1f78Bd+UDJLLYVcUwxN+
bDwHs/erNJi2c44o+mDVjPYA/s0CfBSMkRl9juayVKF7kN6KKBoNhX/DXvg8yXrz
g6qvlmaCY4sFAqkRDPt24osjEeX9COEdw/dwVRsM5kYF8XwBaiwLGL3v2RssjZSQ
uQqTB9dqwSnWx/uKMZbjBMI4fDHOY5LsCW+a1IPhQ4P1MUQqGOeXZ6wbOq0IAMa+
Vn9cHGksKsi3ECEDGJQrv7+HmbgQHJHJzKMPHwa4Qhh+vSufN4Ymqgk3M8mmIiMR
dZk7RB2bhvOVxfVNysnouMjRfhlgiKgpoVuXo/mmN0zAbhJ5lpKZ064SO8ek1lVM
MGkx1cBcL4QnWW4z5sE/NQadQacBD5nXJiSJ5r73a4WQzljRH9h6sd6XdGgxl7R1
qCR7v2SaYOO2etcCRjm07oYv+yvncGHxlNXM6bBw1WDi2d2oP4CVLDrJzEJZEE9p
Oydj66P4LjDJp+siMaQ927HmPlaQ373I44pydyqPVAlBfAfzVIjD1TzboIuJmQDl
DXLL9YsNfW1WOR1Fw26WatOUaCHPcvnoxjpOXQHiY7pvc0rbQ693vtgTIJpVqXMp
cMSA+iQhGSY+Uw9wwTd0qcMivIwcRSTx9YLXjtLAY+m+7+c63Y3gkaCQXwSXMw20
JKT6sDWlco/GuTUSoking92bsjJBf7hfei60aEco7FACk+VGzm+gmdKuQ2YIhNPC
jeivP41t8Eg3esMDGB0YiNC+zhHDRJiJE/cGW9pXr+yMzeuuX4SpkCoQe9D0Tkzw
eambNkjpaFNRB2nia40RcBXhDDPVfIEqlSygYTaw2aVACiDNHdAUgXvGlSRV/zEV
+m2e3T4TT9+GO1CaCJ4yLOLKeIiQAh37QhKzak02B0LLQnOgWR/PONblEbf+jjO1
NbEXHWqQZWD4MLy2YU3hOuH3kKk5CG0Ba8jOI2a8R+o5Nf0pgyW/hOyU7xT9W5BC
r9ooGQnhcaQ8vNp5zBl0Cx8WjlSKvkiudOOI6WYgdP6fCq+4qZVMmCzmzA2xflN6
DRk8DdHWTJdIcNtjLRtfpoIHo2IKwGDPh74iNs/eRSRLZntc4LXnthpSP5JmckRM
41hmw26YqsIu8BeeDM5J31YxceSV+uP5g15O74oI3ppDJIRnV+4UR9sIih8nGtt0
Jvuk2bvP5olEn1UwLbYCHkjWQdA9Gbj5K4awsNpl/V/EP/z9q1XFVASEal+cTONR
WhGXxWvvQlRhaUhEAj2mIyVYDRDXeD9JVHxiG0tq9uHU4gI/Z/5WOc9seKRrG6mR
wvaAOPokLYrvEo220P9BAD/e3Hjaf2MLbuOOur+pu6FV142+4k1SKymXztNxrnN4
xr13KI4c6Clb+Zk3HU+BQbFsKdQ/njRh4Y5z/b1d/pdlV5QETpZ08hB7OdSBItY+
NNh8I9QnDhEzndoutlYuzhpahJcDff4FapxjiUWzUQv+qp7i7r73s8332yxLorEz
a6jd7gpZnryVlzFyNrVA2nbVrltax+rlyV6j5ZQAQKZIYBn834J/sOX5LSk/o7AC
k7Afj/PqyrvPnwQF3bCaikTuyVCTC2Qeq6+UjkXOrBon946Z4YBugv7ZpQW6LhZ0
aQExXsKBw8ezvlCQz9Z6Ex8cM9lHeN2NR6TkXyZoVc3CKcd7Cm3b8EbB0ceueDH6
fAnul8Hdy9ckiuC4zjoH/v5+PNOvEYNKH/tEJsszUXZD9fhtJpzPnD0Vwm1fP+8h
6u8Pr2u5F8/TsrOLXTXebnxlbdE7CYUxncnD8DNo26VWGIdSb7ri5CaI8exY6VbK
OUkXd7ke6GGGgxOc2WodxGB0NnonufPCsq7c1UTdejUNfiV54toiDrhW0l4t7OtS
7vAW4zqT2aghSbILCkIDKVGWxqGIWgpLAfeWhf2baPcemJp5FXxOIZP4LBf06x0B
qa4IfR0Kx3mFH8BJUCF6hUIKrVoUP+1EoJih0OnArTk96Ykkm6jJ8lM7vwInjOto
gAYH1MgSwjRCDeCuU+X4Lq7j71MIf7DST8dvoTpnOt9WSarIiyBjQ+D+0qz0p4m2
P/GKlw8ywNuX+LeHs3cM8I4aFPr9J8gdLUjneXrFxmRynmwLVgNAPg+yWtcM+zZY
bqtsTF1mgig1Rj3yTpy0RveSBQ6qZkbwBtNnGleZQIYUN01xKYa2Wz0kamn4wKya
CxM/YcogLN5cfYcVacWPFHLMT3YLsdQmOLTlRarOZjpznjEnO119nLK10FzpvG2H
nzl9bu4eolaGq4lGRiAMom2PL01EoV7kjFqNOfvLAK2BVAHfpZKCWPxWsubrR5TH
BZWpyETiZt7B7Hn2F4XVwz8d7nw7Pv1SfsAtEGkB8/SQ3/gj8v38BqJhjHfQbir6
i1HSNecMcSftyGvtKBskhlvkCdPzhiFZZo+wlLOq0QBftsbk0qei3Ge2qaMbTrRD
GOtqTFDIFU76sFSSAZHd8iQm3jzRJQDXSv6PUp85zIv2isTKUsRv9oPNmqzE+eSD
VfWNoerM7fCK7SUwPfN3UP8X9tdfmGWtmHVy1APn64USzJRMrrMdw2w1gvoXwgwn
vWXrIqjGRaegTiEXRFLY8QVvWmfYZ64XkDQJJarFW8q44ZLRs2KFpnDysKCTzE24
gJTWdXpHeiHFi5dWvqwqMLnEcuHSSG5L/dgxezxl47wwPpwKFQVlJD4kx1vZrEcT
LA8z13Rplswcm4ijyjqMm/0EI2TKkYQ3ne4eK4tzYjs2+Q5A+4swgn6tABzZa182
imTwHUDR/OmYnTnn1inl9a78MeLYqKNSHZejE1WY7gQ1uXKJ81KO2+eikxCeqe7C
Z2ntQeRr7GaUOuPWo2026W3nKp7keA8oAD8CJhD/6u4PHAbcQWQCDRMCqmkEQtPm
KKeZQv/Kp3LNCTv9m70H+33dlS4724lV1sq0kbNctLqDiGZdbi5m6zjDeMZYqIW7
FfQUv1xLOt03Y/FJTDiCHMijOvUYbDYzjqOOyK6jOGyyFlMnSj3OROX+h3d84oIR
aRSDl0bHkCOqC2xp8h/2c6pHO0htk8yRtswiCO/g5Kogt+Uqvt03FlE1tYAu+kuJ
WfILwob+eJ/u/Iem9Z3A88T+VzNJRUg8VzsaIB699dKQRvTL7knwpirLsauO8pxu
8Vkx3VfMc8KpjwtNeGR95sHf4Czasdp4qL4wR9OvZI2Vt73GoxvE1vgFQjXGwE9N
MSGAaXGmcEI55hGEHrLWQ3fqB6BjLEJcL39sPV/Y9t+v8aP3mjbjJ8H37yKcTw4J
syILP0h46n5PPQq620DQJY6H7n2OAvwnXPqOLDJds1BAuMNPm8ru2JzAeN7GhYHl
b+QDdIg+81VaGBTeI0PN3X+rXqgVkhV/OusnEQtuHAjlxqSBVD2TbziqMZsDkGkG
O8fA/5u/xz3L3HFJb35AdbDJ4U2TV/dR+nA82Mdlm4hIHC2Yuq580hnXszhnD+xB
Ne9+NRVdy+rMi8VRLAGputeQqHYYz6x3nvm3bVUqslPNQHtfRTS57K+Vzr4Cg0gi
8UCfMUEYGWC41GPkvahRJ8xzBGaUZoLBrrC1qz9W4wyHyWwyG8naNzGo/xSwxL0K
w5ieoaFQUrfSJ352LCbOBXS0zgCF1kk5Hu5SSstBOer7b+Q5NdIIFWCK/UObmh/N
7QC/gc7peqV/Rmim0n/sJmNzbolXxMEjRy8rNcscYj+RALi1mHZfpPf+wrqiqgvq
fODywCypZEOEmwCwCFR3xC/QnRFaY0u2BLZ6GcwT0Pe1zvVAB5YBMhB9wq3xhkGl
V45LVfxzIRlgTJtGtQonx+l5c0taxx+hdvAWMKun3KdKeMKHdl/eKS/LARWWG39b
8/qQaSk3e2t6HWKuRizEG4Nb5ZCOdtU3YnJ7ML0slU4ZAGSDwLkn0zIuR4BC1QTp
SaT+PK5bAi9aNI3rvKr6Ljlu9XWbHFeDMOhfBgx1XmJxgEx+EIfX4JOiSzSXu3DC
NzleVq3qoSDkG40W6IGwMkTzr57tH6luWmA+t0lgoPflrghPZ8OHDohimSpj5rH7
O29J37yL0ZJosA8WTkrxJH6BO/C6UZW2iCfvU3i7tCFAbMXjiQP5vWjunboNGO4y
0lonxayD+Xu1uPid1uqaTtpsc5p6IWxECvoxHqZkn1mD603+jk8+5VgdQOovoWO+
gZfZ4LbYWcALHS6YXXKSgjMqYc6fLyvBXoSUqQK4SoXFlZcMmbHnQ0UWpAUTFpFP
ZYCaz33eu8SWhjSqsFtXrWreMfjvs/4qkYYmhVBsTA4j+x7WbCQMBN14rYbq6Zh9
36DwKmggolRmgKX4xD74nUdbwdSMvUuysvapDVnEezk3GhdjymB5GK7pU+xx+2av
yQ4DElPp7tOIU8nIYn6f9pDCwSysa+1KHPIgPZ7pqV5B8o5eSaboH3H4ddVvJJql
W3AdCTVFcSnke2o3d8CsMi/higQSXF0nKxs/3gw/VfxhQfa31q/hLF+2y9HrmJK+
+iz4U/M4BK8MH0Q5zo9VGEQucWTbzj3bXLjbUepA7+s+PPZwLYd5ixagwoWwqHvq
8HlqEy6bGjzlj5IeapXJi9++K+92s5f58dWZlJ5WKhaYExIoZ76fEQ+W9Bem/vku
bhVmYMQ1uVcMdsKgvAcLFLtHqFA4cXHiinLGrdJv1e9e7FQ1lWORWi1cUZYImVpc
JT72v5udHwa0i5abL/6aGKenDQqosVoX+oBxZWZ7n8+wOWjP0B9ZgK4TPv3m6W1e
Cz5Iwy/KzB8upsSqCKsAjbj9oXjJptSuAB5m08QXMDW7F6D0VnmgsDPhI89LuPl0
TM7UnGNBx5iM8CkpQF/CIqZpkFndpmeOpyEsJmNDjIH/EgohIDU2kQ2+e/H2bji0
UHSgbHMqINgQ2CBoe/1hG9A98HzM1uOg0UqML6oTE+jiw1KJmMZ/Vj9CbCJja8Fv
tyoeYHVCsC+qzcyWGb1p0qcKzAO3pESSSkuzKrdmF62SdOah+k4CzG02ZMBukzly
w9ho/bOlhA7ohWvn3ZfA+KSC00lgjTRymz23fb57WYjMS3EZR6gj4UF2YMx+EiZR
W4Dsvuf20V4Fwkt9hCLWeAHIQ9FOjL37aJUEaJdyKbq9TZYLiDNe18qoJDuII8mw
aet74CYx80DSwDoRlCTA+5ucOHztB2ng8GJE7A77zukuxtr5oLvm6ippmbfYBcPs
MavrkvXyVr8QbpUpS0iX+lecx/l6Vo9YpjINcVXgNIhVlZaW1OC9FUMpKYUyprLf
0Fh72KazJC9yu7aONWD7vAMGPYv4dCzTWhmh9Y5J4fSR2XHqkepTqHF555GHtEr7
FAxQGyVzPPXb7GLCjyK+7lvdcwnWsGLhwE4ZUK6jUwtJPqYB3c9mTERdz2xums4N
1Pb4GbbWXop9uAsOG09NSBNQz+9x1ysDZ+lh+tETFzEI23qNXVKjfRFkcfxp6gum
G+ZUKcS/F/LavzrCUj0W+i4ATKJPoJF3FE5Pg2x4bHRxgVjS5r0KWyHftZtG6dz6
7iPAbZ+GVj/HXktRuOQ/LuW4jHiRi9JCkBIHOl7erNIc2UXSlsJd3Gg5HScYCz8k
LS0PAlpsn+gA2SR9Uyt+OErIAAHppICQcZ1+jVvMbOM5jJ0n/CIaJhVEJsaHeW0j
ZMfK02sv9W/7e9HWGDr3E1gBalubhNc8NPiSQe45LvGlSCSC9mjBmGEYNStwfVOu
k2nhhaPvd8RUW8Etxo+cL4E9FMhNLsZcmI12O/o1se4ImlAK2IjKeELws2OoB5J0
jhXlvCD+kooPEofE5tlKnG861SfV43D/T87kerpSb09kiObU0BapEHbfBaolin8W
4rFDq5ck2iq7k6qk1DjkbQzNR4uc2yjAXLCqoFxP2jgthMoMkLNELMyKFXwlPYvr
CzRWrsTzfTDz3O9bKjUV7fKVsz/QN4MksK7QKu28fFm2c4pmRjdiy9iZaVEOokjM
bSd4gFSuPNWjOa9KeJoc1RodLLbbePN+4thygGit9E2W4X73KGYNQZ6BBPAsfkcn
dPVf41Zkx7mwmgnjqzXvCyDSg0dQGhbc4V3lw4923t61v9oXlgr1Ju5HDww7UuHb
4hSE630R1uo+qHtRpiYK6JYRe+X1x5n4PQV11uXHqeIwW8tFGO/E7yJ5EVMlrE5d
bxS4PgaNkjYVplHuGP4/LXjFjCXqpb94F1p7oIdd0+3WQjti5H7jAHhnwzKH/5fQ
A6ZZSjt8r2tUU+i5laGasx1UFiXuEHkanvKPxW1icMrqUczlLa3IP2z61OfxJN2m
nubv49k1mIW6W2IKCqEpatRbL7+8j/ddSAvTvVF6fKbXhvPYoyCqBScAcupsQuOp
xkHexFmnrlLR5K6BL+nxjYQ8ppxWbATrj+5xln/ZqiIdmkCT+omA+BVn4c5QlFaN
dyjKxqyOpmrsBR4/64rdXxzGOBV8RAkQYkH1eDL6Iq9YcCG+n621yEtCXdzMi9Xu
PgbkGUQ/l17iqxLVO5GDOeP4osz7nER0bClMG2oPggm14vh/9vFYbMY18XE6a98K
3Sh7yDKRycTzX4OUFUU74V+1h8SAJ5yvpbs9DWLPpWiqfRltmSxCnPhq7d2Mw2NT
EdvLCOnWZ30jVovnle53lMgjOhzjq/fNV6sl0KZ/64ascsh6+/Wz8JFB2Dr+YF+Z
jCpTJBUI8jEHXhFuC9mFp+nzTsdD6agTa9qZpMrq34Kpsuu169Sm0kQwOzWxgp83
dLrWikGUZPzyF8ErKMvRokj9yiJSCq/k4lytL06+uPbn0cWwhwTlY2i3HvsgtRIm
3e9YEb9HPNU91qoYetH7OlTA6OfuiXJUCsQXjvVS9LdnW3U5AeuVtcyoRt8qD719
R0PciIBQv+wPRNIsI4SOOO8dmpN84HKCtv66LUI3hfQnnPRMZWiFfZ45ra2SISEY
YY+1mypW0JQsmFnIbZUulpdD6AnikRTqM/z9w6B6Hb6AbU29Kne2ZHggExkkLPfD
kk0CiCLDrlI4TWrCxyJhlVbFBP6SD/mgg3ULov2sVB6LQWROGiOIEW2cxHlWzKbK
E1+vpxYMg3351MmckmnENG+jqvcW1wUA05oCRbnZufqj0AfDLB+VcoIUiEy2ZRtq
yPsg1DJD6CN441GDwup0X5ZFILTJrsAho5F1MNqt9PC14+uezbjdZH7BxBenn5hB
LgDe+saQ07YF0gvYmYiacFHREeNq6T90a/dFQAlVyywSPo2AYhVfUk/01ru1sD1D
PcoOqb0RJXYT7iXqu7utKb4ZH2ITAyxIr3z4DvgvrUzZb94TifhWZ1yOikR2+kud
ZH+nZb+cPm3Q/wHyDE9dsA2nHPjrenFAkGEjlZRYmCG3EEsfAigQn8di629q/alx
hQxMDKE7jtBfRjdM0TCe+pt8e+KTG+Y5L6S+L+r3TeSaSVxQ7hG7tnkzMPIfxtF6
/MeJEHZZDfJej6/OaELNqXIqkgEKKvm6T/z1jDMcmx3wtMALDyYXAbTkamOZmk+8
4SF3Z6djtJH9HRVV4MSqlzqp2FvmV9NwJ+3leDUwuLsQcQZqEAaJy4DMTftQmvK2
iJ+u/m5sl5p7Iye6s/X5yQygIqsrYd/OnHcxLa1sH/mH5FH48iWBvcS9TlIdDvGw
Y7eHp4XnLuJ6uslNHA6iP9lLbSloJYr6d3XwK0raJQCL63jQAGi825p0Wy+75N+n
PqjGk3BY20okdPCGDZUeJF1EQZZ00dW+yjrLRNRgqe3ClXoPvUNR0Jpz2zJluHgJ
xkTryS0F0JzSveKphkJMavxhCQe6PQxydukwifmF0BKD1ABYxDAXcoprd9pCOHv8
zsWOEip14OR7zuBoIrq+oeaxADjDkEibv8ttkfvKRCKDTJZ8MEl0LW48blUZSSCR
6t5uW+M4m5rtYcV4UMoeiFm8p/azdFFpfuvz/MbRdPZKHcOh7/eXnp2AMGVTGhfE
QmeWF5gPD0lqO8VD8RXn505MDiuoYIQw81EkO0GERzgoROPLRn3XFpsymQ0w2Wvw
fMHgqi4qQhcYYsPizP2cf4AZQeyOEpctLfqYyKl2bDrvyFAFC3J0gIiYAFFyrnYL
bRfzRZq2ryWAZYIgTkdFpLtVxb2JIw8NAyHz1iD7zKn83hgfGYZv56+1WHs3oTGJ
MfbXyiNinIAA9iwkqjtfHWccJdHUDuiKLjXdXii6C/69bOd2+8WiCu9QHyFcxIKI
YxG9QbySeEDISZ+OOXFOr94DQi+py2y2HyQOHcLTFMcpUbWHGHotarFV7wHnK/R4
wX4qQWvKb8T1gxU7/uJdvItcCNHOIBIzukqkw22KokkfkTjciL63zyxjqALhpCs8
9kPxB6w/OxqHKe3ffoH8oQwiun1Ea/0r0PFQXOuhLr1BGzdiorpf7LJDrmj3tYZj
iWlZP53p77SIwoi39vny6Tnzc83rZAOJlXEiZYebe2ykQvqWxPa7gfFByCTIZW87
ETfwwplbu6bR9GPLBXAaucWwyxXw57OaK5H6zt6kHTfoFd/nNJnDqpfbyslhU+iL
d9/nuDl+kIGscqUGDpl1MayH5xjwvgBY9KspGVAJZoZsg8rY7tA3guVv2LWVg2YH
npgTM7XC28CX6OGfYWuJ37hnwE7b13inXp7Yyfz4X3IpVgfzZfOEXyN3f/D0mttL
KNe8IY1nMr7JC8iqjA1bUTBRTniOyTjmR/eS/gg2WJPsX0YLaLsEWuIwV+ZxouId
knKP6dl/RjIyVhJCJ+2CziZLOEPO/z8AkbMSqpog6U8DbkKm4NJmfECics7Fvd9D
zw2dpxNdo60k7O2mCaecU8hRahM5VivKydR4Pcb/43TBgxEE4SUxQ9AqVhQvuvBV
uvtsnuWMdxikCC+rQbFVn+Bb5Wpc//opIUrleQOaf3n9faws75ObNze3qEIDRdnM
JPiyWIizCToDkBWiKv2hI8BPXNBZBXv+1HRRI5Hv/VNUZ2C6NRkJZ3tKIK0px+Ei
H1Yqf4+CTTf3ihO4O68i0SE2p++l6pGET2pPRqHIHVAOZWqf5pyNu8oDSPBufjem
Q4jhCDkP+q7wQxSk2aRNcW6rvwoel+NHlTWpslr1Ci/TKyYcBSW0z9UP8+JIssPA
PnoeJ+3/ajtVIX09brI90D5hGYp/dwECkEyo1kMzLxj7IkHTDij1ncGVoyqlk1va
+wNKsbjKuiOEQbRDSpZClbOk5Qn8n7kYHWjKsjeH0xy+jM6LWMYzlk4H1bxoNMx7
aMB7jnuCdX6nxbUkfc3heHCwNr0LHqwid/0fUoNV0+uDv+HdpYPH/jugY9Fo85hs
4TTehsRnljuEaEHqRjzJo6olgZxZQ9GeKMaGoG4zGWbki2TeeQ72Qyo29exdMVUK
4IRz56qT9TVYq/NeXIZDLj4g1ND3SkkbPyQArtFzN09R8Av8/c/1kb5DH6v1ILHD
vSBOa1mCmfU6hgcNP34gzmLvZpZiHjaqLHagUgoXa0esgopdlBrFHv/iLzehbz8x
H90ooYst0RRjasPXSGiK5/jNsmOiceNHWT0pi8RnZPWUHBwNVQN1ncaY6iS7/Dri
CkGGMDprftnP/hV70jgCtJkdQmKEkRLvZXbUBbn3xMiR1cmCHy8teknIpVCCRbxS
5C54qJCLECRCtIDMSbwKqa1Xv75wZZuUInWDWOoPOgIK76au2hwcPXs534E8l/UF
j3AkqBaBCLr2em1ZyWanhj58oRVc4Je826eAx9jI9VT3HL/rdkdV2erdxu6LJzAT
/EpoT7QcnAwxZoe0NYpt/PmjcJ5lDW+hlRsPCdn6M8eZ3tOf2uXYsTNXPl+MSjGD
U9KXabEjiECgbmIWbLl7QSD5Nt4LfiMZI9CgaD/c5DI0I/EyPob1wqW+uadbDwSb
gEJa8BTya7rdPdPywWZGXsM2Uu1K1zAGBn4joHGGFKnPE0ePS80xqH4hi0T2O0Av
0kMHwdfRDVwv9uYeDc8xYtpwEPQ+yYO7ocGHQUOfYrEqP0g/8NFHeeSocdtjA3Qy
ZXrcKuUR+35y4Q0ddwrUM8bCrurxH6E9QP+dteyCAwrA33ytSSv0p9nvfDPAm21/
hYkowVDTxwAd0kmtViy+5cgPgcjfxJSwGKkbvD/wLmzV5w0lH/8u5ptBfXH7FXKo
BPFSmikVSOn17H9Bx7VRJDW7I5XHvF0tt1PBq19pZz2lVBZCdh+ZHMOYq7PQ3pfL
nvMA8CN1QCcq0XfV0dyOweoeoiJDIJA5B1vwafpUdU+E9rxvuImBMqEVi1VL/bOS
WiIx4jdN/BCY6SgtyZ7v5lUH9VmenpwdJ4ZV7Jus/DrHvDVMw2fcE4qaluu5YSs+
nTlH+3oJQDoF1PPYpbbXfuFRkUCRrNXu7uo6HJhYLeDLFaIBU/uv1FcfUbIwv6Xv
2u2v9QV/8Bxh9Q0Gb8XpLs1nHmZel/6NiyTUPlJEQQftOGFRiJ3Ez0LrQUJ6rW26
gwhykq+F3vLGDJ2TJrFQ8+VsYY/uURc7sGM4YVhKs3tn2uZwBb2wSif9hd4B/1GT
Glra0oDyQ8h7kD6R9+HDkDZBPN6jKNR8ssrRaY797heXNU6wSqZmo4GXNeZ5VeIH
3pDAn9fWia9iiYyvF95r3wszlhn7+gAJLTywjPu21mQOKZNTMuYcNl/FJ/XedYHA
CvKEzmMOScVgKqKLZF1bS+H8nxCaX/P/uORCwgDxZIfOsFXSJb+MdIJRwD+xZK9S
nE2sVlCkEGz6KljpVOnoqt7gqrT18mI0zfv7iZOfj4VDCKMP5LX2IGnQDAkf1hyN
ZFbYQNHz2w2ZR/lIZTkL+HQkYbhCrMrYla4IsIrKFyJRmKGHjvQiNHJj/+0BAZro
B0RZu78CIKdg7m5qH4on4sDYzQySxChoCLqod+I5yFcqcDjeXLnnsSSXn1yE5l70
j1MKQxvgu7JnlQSuBmD4uMA53PFPIxuRpI2ihYtOvTw/m7xIdYr3JzA5SsbfL/Uw
2f5yeL5rLXzV0G8gE4lR38MJ/2G8UjQjJ63o5E+08vzrfCWtkYiZ8JT7Cmj+3vy5
/J580hnq/ablY0pMgvzatie50z+L6QCssL3p7nTOpSuPbjj6Q6E/5/+XKC6UPczE
NSZx7eEh8x/zZe8HOjlwQ0WMYqt3+WOP+sjnrKK0Kb5//HKexD2kRzWzJgvK3T2+
dcE425pi11cEMGFlq8OsJTYevtGQLF7CIdVhl/3d+A2Rm4/Oa1aevJ2OJ+z15sIa
B42eDO/vAlu/2/s0OP/EJLIhzNqXPfEWSCXaNs8C4DcDHTF+h0/X2LasWulPAhzI
55izsaGUI+XywiaNC3DBBQDBlSp5ixFB/dtpx3AuDE2egAX2R7mMvUJrR7j/7bFI
g01xKhP6K7fjpsOpLlI5tnpZ+kaGhW2Jndo2RU+LrgCAz/ZRUCZWCOD5ojHOv3PU
F/UCrubgFyDxTfD7NK8BP1oGNs9ZNBM4F/jbfDE9LT+8fV52ep2Hb6HoeDRHt1yX
IPNoGPlW6XXs08IpcHVpbQIYTemSBC4Jyk662ZwYv5BRzIFLfYybF8CIi20AWWHI
3nBZ5Z+BHppwonlK9S6OawVcH4BG/65Dwot9BBTowlPA2tRguaufqYrNusMdMXQk
K2xJYWfP0IsHYgJ2fXXkDqr24SsqAjEBNKNjOqs2Pcn2HxaKPzaP0LdAtp26cZ5c
z4nPIpf+VgKfvZWQ1m9RAJ6VQ7aYTSCxkVD2rPe9XNcJkmfRGC0HZ3Fqb4BKFgJC
WpTCXSRuJ5eP7ICKGyaOA+PYuCfH2Jw/HnkMiWcqWzZFA2S62KeGimQ5BmfYxzV2
Qwaqi+cDFlX79YBPZCD/rTd8r2gIklSIvQedg/BRauvEl3KupqtTCTxeFPmBeSw2
GXKMrBN4M5tBVAJPNOVb/Etefe7cBqE8HccCncZSH3cyKb8wj2aNEltm3Bbv2GKc
7SDWdUL6MkmhnalAYqKVlvuEDL3Fd9GuN8ffGslWkxBW3+4F8hw0p5xfTvCe5wDK
RaMb4/zxxk0XZKGGRjAY+l8jsQKH7gdYnxfIDKKcDMyk5gHp5/4cr0yRboVH8+ZD
2OhEVtkofRNlXmo7AbCYa5zMwHOMvu0uYCfy2pgIaiWBuPxko/LBfV/YOpe74S9s
aB59r7VKiHTEFNM3K9krOFnzKoPr+Y+HmIvst11AhbesNrLc4TL67x7FLcoWiTdj
+tFw/Ry7mYbRSQMmfPIoD+L6tgLahd5WEgrq//2mdogIsVe0L9jx5ymgEVFaaiv1
5PKX/A1lMs5ZojzSXkwSYhJ8zpao1Mwr2SBuI9ho9DwampMc2G7CJIV20QAh9RiR
7mUjduJ/EmeIUXI1M8PyP8jYeYXFhpPFGnG8IE4XrB7j4qFDyK18v/scILBwL/cw
CAhTbZDh3ovRD1SL8rdBrmZAGBiGx1SI9A7VuNqaRw1mENd7hmLB6iLHjwidpCOa
68GKUmGBWUBW3WqjP9IdzpofKp9qTRV6jb0uj+hGhc1x7poSnfOYoV+AlvU1B0HZ
lNBQB3gHy21OvLBlGfVFIWKsZXIXVWE0s69ke4BkrQDcQoyTO5QG1hbSFEDESp24
eg6wN09pYLK9fCJmxFUE14I1/uRPLbRNRdtwrZA6vFupygDoFlSdYj2D36bXyF+K
thyJLFNJBoAb701UhrsT8A==
`protect END_PROTECTED
