`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viSH/axdzPakIFCRJ1cKNsEBici1y2mJFsoOj5neC6SDQ39w8M0sIM0vMRZz3vwx
SB63DemP2CRnJIcWmOYB/rAJZ4cyjOWX9b1tF3s1d87c+8DHCpgVikgydwWEnGze
mwQgj/9vzwntgyG6eOxdp8tnCGwwkC0QlEaNK1IHF4sYAxvsGYsVSlOFVntwZbLg
MqajTasPTL7IKEQuWzuEuRH5ZRHWd7Kn7VqT0Vz2rLeMxNhRbdhu/5HiheUUdRh1
1ZQpsLyJ58VC1E0hHU1HE2iHKlATK/a4Wi9L/2p/q4YeGmU2vd3fcLlW+G9+wOfe
9/x4EzIca52t+taCa7O32QYuH97hqDkl9kNecAVnfNI9nzEoTb7S77ElE14HL5iE
JlkptVgJy6BfX0pE1FJUBFFdcDjKUj68foiAzsIu1wXVsLIJ+pdzHvEG6hiGYSAv
hizTnVP+bldM6ALAlDIFwKcWvckHfxrXr9Vwns4Eztm+gOSCJw0vpbz+oiE8EQNy
Ih4hHCbQ+sOrt3CwCwebjJ5zYvW6VzA3IMHMxTQ7iwqtc1jsdBMWDArnbSRi/K0Y
uCVJUZnNX9hyHpS956aBnEPSNo5OrID3sOrziCZdsVsl+Nv/dtO+rbv4Yl5bIyPu
Zyh6DSpAgFK7m/wG6BQCFcuEZrce5PbKrJJf0CapaVYSxDOSZOP4xhO1ex4zEnFv
K3bZu7tsWgNtCocnNvfPCcoGk9YGqdDErnBO1+03mXj1T29l6hskab1gYEBAigmg
CTAGVyyzTC0O0hu5XR2zSHEhVVjRhi4cKDC7gGVg6DuXLxBPmnKB71+rjBX9xmYL
f7a4ullk1B5VSBdh+kmvtDygILvUNscWJsbiIwst+JgYLU1+YCPcGhI8bf0BqF/5
6qjt0IteJ1486mw/AGi/zcYlUq/32lulhsX7ECfVmJlXeodd+2WVeQ0KseV1iV/J
Uaxh+bpWqfDqsVjC3hqWudQciDtblQlODzSL8NGQvGhk0optmftsYfDVi/DEHDHw
pwwg9JBu8WtYOyfUm2XyGikImOEHcINbKD/GRsnVnes7nAqIyFAEw255Ce7HhjoE
EkwlhWzx6TjRvBqEIXVzN+mBvMJYPiwWYZk69uBO1b8YYMQXYcxbOAv1Rlu7WrWb
vrxfPexC73RQhmJg257gGcZnFhajdSQuJDK5DLmILbRiKpz+Eo5bOgGyru0368SP
/GUn+F3Bhn0rsMRcH3jOLGyKljLaSdnzRWS7cnVlfEoc81ln/RIK1RyKtb+I1pf6
/eiTn4kSgZaTqTeTTtv2PM0nwahRfxnExy2BDCxWiCFOT2HRMxac2Kg8/FSrACqa
/cxgWbvBztb6ijwBN/AN2SxzJiMu8sC9x/0cFv7L3B/ftAwu7FW6p5JaZW94v+Bd
lL3LN7jj5u7L0n4BUBLSpnm0Ph99eQ6oXmSjmkpkP6rTkeYL3vAkbHM3C2yfpsDH
`protect END_PROTECTED
