`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOTNHSJxefvtmY5XQ3mKFDpsYaKkDvKXCD0yWoSTbnln/CRADTaZva28MdPvji/O
Fn0ZBFx/d4HzNQHMhc7D8Q4mlr5tS2vgeqXiOByTHxOi+Bt6qxW5PoFgIj4MWAXs
Q4izuu3K9MlDq7+8bOPZ29hqpjxQ8oQhBas7+Cqr0WvVPtAfMqzIH1vI9Dr48F2/
vGzaMZ5RV4p6YJ7zkfz0hXSwJg5DyCBRwjscvCMXJBHr1zIEZcnrw9nQL7ivwQ+8
IsTBow2Xg3X2VUc0oJL9rAoyvHDdD5dJAZ4ZXRi/x1xuCRfOADIS08dWe6CTs+sH
jx3HCp1AOJSplpnWtI9dUQ==
`protect END_PROTECTED
