`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZQlUqENuYSzI9BWQXcJgwQ4noXWT4bvTC/iE5YJBYqpNdZ8IwcKFYKTpGJE8PPS
fpvQrx7P1G5k54/Ui5dpusf0UJbyTI+gtTXTPmGpEzT8BgwtdrocnXT2BB0uZGwp
JQjR35QZgQ1dRa/2YD7tDbtVfHmXPNqOQ9qzk+mVfiDiXC6uxl47DotkiSNYLf+O
TNFx20HUu6DAtfQUv3N+5rhqgFKH7MTXD29zhZ4NoNKOMDNgTpl4WLyCTQnCTcBm
OH8iFV+1vNej0mQC9mx46ZH8rrQozfMbRECrlaT+jKmUXOvyuGVeYeRGC7DzMxXR
XDnh0cMBn+eBdoKLdD01GAo7j6Zu1sMK+9LgzRNTgWRNqqHHvYPFjzOcXDJ0n8QN
ywLhUsUbN6uefYMhfqYlREbWF1pk92hjZitz+t6lM0eZYmgAAv/BFYZrEpHrO14f
GqcSRAemPhwFWgHu8M4Y/OT3ooL+vcjwrosakI3a4is4r1ER7qZR7O+sW2FtAHZ5
pOBV7hIFDd9hSogS1QSRjE7z27IXUCKMQKYbC/3AV1mg1Id4b7ZirOAELK/go5pG
beJDZEmXzXSB9G7amEEX44UBkrMejOzacdyH627FTIp4ixAGwyhkx4r4oX7QdOIx
TjTb2Ir5O90lyk/9ueIucfHGtep1rpMCRo7H3G+mTg1FjpArD38rMH1jPQH80/YB
jD+4B6hNj1rL8+mlhHCCawNVaf8z+fzz/R5yw22NplibmhZqduM/TBZU8jO8oP1W
Qw9F0kGZghGMDaXC8E2V8vGmWyizCFJjOUYtRBCLtzWas8oXola9Gr8sDv2nPiw0
9bXVKMK+cfJyUSkBMuKKIiqkxhuMrTuKmBXaUnQyVyi00IU/8gQNjTm8MW1OvqPS
2xKhWPL95/doee/vqfup81BPSGft+FjZ3ATDwR+bM1hAUBW2gGCAHEoKinOomlsV
VodzshIsG/Tu+ZdnoXJYOq4m19z1b1tat4r/+jFXzsLRqok4CxWVMSSiyJ22B84U
BoR1920VGF+wB7K2zN50fAAA43iVgvuB1Qzuu3wbbXwD0egyO3aKzyKahGOv06UI
zL65PKEPbnANbHIJGlR7Zjrs3ADYIxjGT/gsSXXwkvSvKTRYBgVPOGA6bAcLwWZr
1J/R2cFC9QZj8eGMrzWZzMw7INhjAvBDJ0be2ZzUL9BGhuAuiGYkvE3qFuM/bpa1
GJ49VD9tnt6vzefZ2qobch3S9nrQd/FxisPK/YocDDoulVlFtcT6CXIEt9oXHwa4
DAZmdcVBZmSHRk8CszeWRpeMFgr+4buZkI2K6NL/HkDMKP7xKGzHg/ykOPOWM1yH
FnxsHZK0sTCtxq6OwAdiuObJP/QLe7o+u/bN47n0ofwnqrkZIrM1hiSkaLX3j6Xk
WH6d5TdZlW3VKU9WvPlYgkZwB9P4y8c9ywDzeOtN/i+QWC0k1mHqwLoTedkz83WR
VBbetrRT6w7YxBckL1BeYA7Gg2pyxNZtzOUjHB50ZjqZKQS1l1orhhSK2oJD+DGl
afEwHow9bIr4r19axFR1sNLi/QAEGkjwApTM6biFsVwmBdxeGJz0alvPcPbtdqpp
pfnkoGux91Rcit0/s7xLnwrNEq42MXU8fOYgw+omT+x8Ktib7Q8tTnQbSnH64Zn/
g8BlVAy7qqryDia6uk9ShuqzAhrkEb/P0FAVRHlG4RWnPNTV4qE1ieawzygV3yA5
GatIzWmEph5FUbxvr/wDUr/dtEmm3kbu2ej8bZue01rFGfOLH6bDDkQL4sLNV2QN
xEMXks95Ra4xiszJhZb8Kk1Lg4VzZsjhCJihC/pOUH9kuQaUMFCD2WWCFFUxS+uQ
+CZCRsm22oElcXXDpjrLHitLqHF7xIn8n259ZlhnLCjaDb7JXZXelzz19v/uIHub
JJxdb+QXLgoD8xsRm3G8+wXtQIPe8ZR+tZ+evpzXoSrl1thcbdyOHK1JBavvUMvb
tJ4l8nfly00fgHr76YLrrdRQ271cjb3dDxXp7VLlMT6Dc9Ur2NuGFagX01DmdX6F
YaNzhHriDACKm2AcnqEsazyQrwnKSHHmOUxukjJfnJdqumsnawJdDvwIRA3jaKfF
uVMtsdYKCNgf/lQ1B656fXaWRiCGx3mIydcRFKYx6y7XfIWEoJhIVZzYR7qoofD5
FawsACZ6Ie4zhVmlg84hpvZjmkWVB56wu924Vw29tw94DsN+YWbVXG1BjPTRMwnh
M44/YIFxfgYEimDMTIObjwxMqDvMtqlon0UKL2SAeLCfHnRQ58p0OeF+89hf9vho
79/SxD6P4UIhk1bX5lWJZSA2ryo065hpN1PIW4aLEfVsiweIP5A98v7GcuSPmKB2
k85VcSbXsdK2m9uAnkRDNsUqq3L/0JN1NhA10s8/wd3wxWZ4ywHGy+rdnLaDC6pq
hcZqO1X5umTMkK6g5qe/4l2NcT7yVanX2caR2HdNDmETda1pgyA1jQ3S0Gg4oIo1
nZCMswJOAT7zdlFtmHFAqERPY9wAJonEKwoDE9qIWmVc+5DJh7Ifa3OMdzPkQS1Y
+4tlBm7d9Kz1+CPtiSKzLFav54A09cRpQqncLLYshSSh9wnwcbvwi25dSlvAapF+
4cxzz4/na/eLC+BoLnzF22ETlb1v5+UsWip2WN6G6XFjg2XF+vQpDFUnBTn7bJ3g
FlaZt4Jpwr4yaL0863vOgJi+m/KqCrtkoNqHhTUwLpfkJTXVOpMbgFlCGBIyP5Wv
xRSUtWFtDJPetKsXEPijq3Ot437211uYsMfyn3iJGareQkerAajB6kek+dxbQkhY
UgSD5x1y6cJ0SrgHVmIaNohEbnmYS04FSStxp70PLNleNFSmMInNm0lWo8m096NP
Ghq5C0KnO6WyckBHqSAD3tCjsgRwToc4zsoVfq+yZeyVQekyb7FtJ6obTGkqFkFa
vJvDGJIXXbEwA2ya/WIr9EkPaX+CuoSiG5TDdB+sBDltvxcTZk6F84a/u4+KkK7F
xyxVkWFb293trgxGOi/5RAOhocTQQZxNJUMeoc3DTaGLrnfYlIdueoyuYN+0UyQJ
X+nSxXEA0+XtCLuw0q3F7G+rqdRQN1gAaTHyBzUl9V6SRukkoJMPPswcE8atRPe0
UOaolFp2Fxjnty/0x4LHIxda3WFU6uC6DVF4ng7RlQROri3IEt9QnLrZvN+wXs3I
lar/IPhrsTi4+B6KM55UN8MFBa8OEnsWFJV5vH+AqehtXHJHO3ZgWzOK5IKPLoH6
WLXJJWpSkVSmBEidajrUNUHv7K17EDKjreLSnZlzjxnbBKoTb3ymSgkBJh5RhBw+
J8D8/x1pL55I70ZsfX/iycel6bRFkTLdLCjQtBWnBcAyTBOkMcXaU0vXPTf49vpj
cTSCG0NITy+V0fE/hnZz6C9QLzfN0ne9aY6WRI8IIs4mi4enKVSdm7emAb4NJBmG
XOXfmpBuSZ6e5BZsYoAPUKBaYIzzuZ9uAJ+Gm4hNDI/1Sz+gYF+CRRgOglzKGp8p
7hBAoWjmCiosiXQl3S5F2C3VY75oVD/kJXGM2FToUqveRfBVXSMfJ4ALCltzVcxz
6HGXVc6ec52MOCUOZR9YBlrPdzkun2TvtwsGdd32MedgnCqU68nv6lVYf6nbWEGE
3apgdIPYyK+hxGtkHGvsQeDb40/kfDEkJRPiH4xh8m7zXBTKaJIvQUQ8HcUJ/57g
GAy0KB8dlRTHV/8YQ3HgwwEJMhTxcmUU3tgtHSgD+5yGeiuEEtQ6oAr9rmx8pv5X
b2nWEJSn0Vx5ff3dDfH2ngMglFTxDREcc9pL49tM7XBOMqpcTqN1tNK63dFlqHLB
hMDJGC/uPwS7TAK/fwiDpSgm9fLC95eaI5GXBDXsxEJXFKtD1Zt0j4MXVjZjK6mP
KUAPrLMi6I2lFIXrJe0tBfBYlQIsiYV9XI4Hz4W6/GzCNUMz4CTxBcaDYTdnOyBB
JOWTmllfVQdCjIAZkKeVOdJ/qfaOM+L+ZgxEUGbG6pcNtO8p4H3vHI8jWg0/iNaT
1WmEaJ1MG+EvIs2Jtz7KK6JptpAdb+JYVreG8nzvOz60X6wPbba19lwjrtOaDZ0E
+OlbUoik75QQ5yNfyxOZ+au09oEH6vvEi/G/C8CyTJwPY1CTPtGb7Q+/M138xAuX
EqT8nqigfWCHFxb892a4G0QswxH1Nk7uzm06570qeoUid3K+SecOqRdiFMdkPAOY
fgtFoDSi/zwkBNJE2lpJ08lU7ssk/BW4PI9duz8OyLxxD5vzAPvyb7ai4V5pIPsV
ustYUjY53YsRw8uRX+ESph0/QdfpwzVe5R+n5pFP8joA26etB0fYsP1PT6quvFB2
OxAXGBECIx8F3xRot4V0wU+QzuoD6fSEYErKd+jsWzGKtjdGFzVxVHbk1AefHiwB
tT88OF43RHh2Lngqa2gYWth+Fe7ntN7mkdXFTE4+afagiJ4v3P1/zI3q7ofylDOy
29KAK2HdFkkdvizs2dMO21hkUDmAk63qS5ZlB9ExLsgVh8FA97QDMhoIScwh89vU
OkVvaWyB/A6x8JYpcg2FkVuuFSDpPE7E/cKT8IBpKT/jnKp05XktyOa8NFAjKJ4I
ozrQYOaMoppmfgUAhTQlxDV71Es9OQAhy4Bu2gBpwABT1l88seOMag/390tHLKKd
Fcd1gYxUHkZxm80MZG/nzCRgEwcoCQ5W81Ylxi9WyOIjJedmAXaapmkcE1JB+pAG
TfSXqzXombVCKjt64PBn5UQe1EFMqp3VqGfIGXe/emLsZoy3sklvcaJtHDwS4ccg
W2hmltvuECszQdnt2HeS1d5JqCzAYSdri6g+E4UehZdvPRdVyrcnfWw3gt7/RP5A
PXmUUGPAKxWKGMaaBrSwc9RV6YqMGLWU6mGrDkE7MrS5hmpRkGym3n4NLgcNnm6J
mA6Vu642wWah81NCX5+8B45iubD0jjPMYhzaVN+tLTKlfs71QCCYnfLWDLcvnu4Q
g9P+lI32EFvLCzGsDoFLaGdn9PeZw6O0j2Ej9rqNoPxf/qAmRCouzwgPE4Qyy/+E
TUOm8tQK01U46ggl5qQ4ox+iWZvFR0dIcJi0YLhnCYmnf9QnZDCRkxtXaGHy9n+u
gW/bA079rSPG7AjGv/on3fCgKlAVyD06hDdZ/KRnUysCyN5yLUx6KbJRRSzQB2TB
EhScU39cUMZ+3GMkqSFKjz5eGzpUj+vp0MTnvErDsZOxE7FCKbBXhl0z6oLYz5I6
pkluZqqmiup7iSYKn7SUm1Oeh9KndRJZNuRAN8V9bfDZSlkLSfsoZ103blcWr84S
3xbafgj+fNKmKrQAISywG2OZ19yfi0XCIp/BS8HnVOrQOtMckYy/68GfSI5zRcVI
L41nG3S718pZDoEQsmOo8l2sOrHSEs8PEmOtPaZnCckZx+rnyZ/OwedVQtb58i0/
8tHpEtgD+LDCMpAguRsfGZ1Pe8KgZtcUryg0CKuSulzrj5sSwgpDm4/5dRdpdyXQ
Vv9xewsCLpQ3KgMUL2v9We/eCSUqaUc/eSeNH0V5zbPJV0kuCrr7kyaJKbVsSTmZ
tfiIEMHixQb/AnmgsLJ5UgUh0xxJigYpmmbC+/OE99AbHd1EvB9vQM0xhmun5xh1
tc05VswlULikQMbevngvVKn4gyBIQqZnIrKLfnqHaaAx8Fq+NVNK7jl45sWAGMW5
p4LHlRCVczOV3CVnAeJGx26xSjzl2yw6k7kKgmwJtb/XuacxxaqE3wH4NHEVdYGz
LPiXcUmAs7JNddO5sSO/UtlHRPu1VWMIVbHgFRSNeyN2wval4rm+J/VET56TK0fV
C5jo5iYV4mCpqekbS8fKxUBXQ7S5Vfshmwhg019AfBSCbcg93737ADsHKVCiT51j
k+1/nKTWaI1Jer7zfkhjwPidOe3W7GR66D4nR67dCEu/N9nKy3V4oNI4MxihzOIk
CisChqEFec06XDtuWa0Q3RpeQ9lceTcdWmbNgt7mMthaVfw+MH91cNNIxhb0UJ/O
1zAxx3uEsJvfol4RJXqrJpiYoxc+rj/lG6S0lYip5JEoKA6DcE9e5LXSX16DkFi2
rdodXUd/WdovOEM6sbTHeXwet0ZFfgR23VJF2zDOcyDb61FuPza6PD4O8x3UiX4X
/Jyi1JLxexlugluIXDEvCDaWpfhfMnx5baj2nTMOgk4KneE4mRiFadKdXmcWansL
bUQ0GYOt817ft+6bQ0CVQ+aE/hNHkigu/r3JnO4zOMvV13+cN657aDiOIcpQnn4D
ECg1u91AsT6MB6sLvJxzlCUDHXLdNLG/C7dnO245IIYLi7ov57CsvBhGuoEq+DYh
ryCkQUCURemXHZ/7ErPRdqXDiuMkTXgd6hfsJKyBY2o995Yluk8UAo1LtF9gAOQ8
Wkrtn0alNhLkEk2q36ZO+trFo5FOZjZb7kr4r/FU4BvQSnkJgPK4YrlHRQus3FiU
cR7+/JGo0SBQ2to1wgtP9bAALGYzXeu801IMRYq5UjADDTmd32lr70GYJHqQDvEw
yZL3eZ5nWSkMdI+oyBiS9t+FxCrd5WYXGWKp91vrioFN5N+QgNrWhlg2NrbrMcSh
MICaEdF9zQNePFp3bUyLgtoCOqK+6gKPJqlyqbEf+d4olKjQkPa5ej52/k/PbxDa
Gpwe1ZXVNla4Dec+Ndt//8S1yg5TaitqIMM/TMpnuhJY2UM1Kbdw+iwTy8X1bYIs
s83mGTXPeKLh4DyVoE2KgvOdZMw+R2l/id5qBKDAOrG0QG/qyLneiPaLUzCRKTgp
eAHh+Nd47v3z9J+H7z81ZkJHI5VCCLu7yoSiuDn7VQPFKy0Q/xAM/nSSfBSyZJQk
oSEZuIC/uqa0Drwm8x/56VY/oiEubBDPvnUAgiyNvUVrvpcZS3piKRZszoTGIqRU
LZ3iE1QKXCRkxH0oyvfwYZzcvcl1FHVkZsU1YkBRITu+yMtFJXrlohUCeU66tOfo
oX/sIJfexDu1GJOuMGJrQMfGwkO2ijGzggNQvC+ptOTM7X6wnbWoxbBQrq2zbT4y
yM8SaaTxP25Ii3bBVsuWD+bQRqwelDPuNTrRvJxdIFh9ihXsS2USIcE4NwNm0qb2
nBWnCsPyZsqRcoQ8PlPYAy1fg1RMrcC09itfqC3zkFBilH9k9g2D5+sCHdOl0WYj
CTPpTYXdni+1Usmv4Kluwvr47hJiA4AnhsEhHKoO4Q+lyL9ynCH7F5QZ9ju3aaVM
VMaqeKrNKN4oRCt7QEtcqCl1amC8WLba22Hu1lf0W35HMSVKrIKsTU7f5k8mfMuR
YbGA8x9MzSydhOA0qCwmFcmAFI8yCvhYb2eTwQcjtptGcuBkUM1yKIMKe++bzhek
PNx5vnJqO7PvDteNCurdGw4bXia+OS80qoP/yfhsKGEnWvhVhG7yPm9mrCmXxIy1
7EtrrL9jsyiktuKi5Lel7fR75pj4W1Bk57a3KGamh3DU3u0WiBDnrg5kZqS/i8gx
MfyqlKMmBswsn304eeaCocbukwjN0BLx+neUyMjFzKs4bL3v5JIaFeUses6Ewps3
rPFL/Whz9QOeEJmxTDW/DqennQ0qb+1K8EYS7S7Yi88jHwdlpoFdpnQ2UomK4mNM
uzXZ0aWXMX0XoeNR9Skyf8wVxJmSp3F8iDe6In4jzcWYst4V3pD0z4qZwPvSXTZn
qOxGeCprMxhcykReSM3GesqJl3oozSmK/OvL1buqejkT1hXWX6es+EkVtsV7kbCS
oWBc44MxgqR4D0ejI3Bi+ZrBjThm8PX+xCCxYONENy7pq5ax5gC0gDxRR3s5vTwX
pNfcUxObNEO37q6CBWbuXxBMKY3r67N6DExQyJv4VBs6sPcrx8v4dsLEDjSTYrnR
3evNmreXjEWqO4YDKFutTWI4+IN+Lyc8IUhC/bpDlGDJ6Q6Yta9/Wo7Baq74+RbN
fAOUvUwkiuBJRArAgvJpuwOOyWBRhz8OH1IZuIsyNXpw+DqJla+P9ztlo+K5Hm/V
/jK8eAZn7A74V10TUR5nDVnD+QwPYUHK8Dloi2qxAIUayD6u7iAxGRGQ7ei6ZJi3
3VKR8UBcChEoDiIh9fQH1OZz3XNKKV8xw6yeiNN3xbLaRfVBBsRBvkQRxV9xKW1+
kaG856RfesYGkeOqf2pNCJbn5sowPquj+fOXxXxybWNNyfGYWwF8393WM7rTLySI
Z2K4JV96zNOWZZqboRuCGqKyRhZ7eIpvJKuAu3FZn8dO+hezY1NgeX7zZXgfp5JG
XP2GT9ttFOmp5i7zmHFvfVWyUjcWKoTB5oZ0wOi1P6/KGhBAxoLBx78sSGapAMnL
WisksujkRX3fxDPQHqSY7kohwIhSK4nIrsOIlevOSpVYSSce4awona+oq4oh75MX
uDedSszvCCHdLb/QlCAl1v57ygbXtZLyRXY0O+YbHaJaeyoLIzviPI66F0V6hSJq
UKZwf2KG5+4baEtPXto0PQwJF0nFpU0wwBzesSVFZs1J/0L+ZKyjbH1nC8icVpIr
ax805RhMB1G0+gmgH0wFymPh8LNvYCdd4fn2xCa6/OBvATqGi4Cv4rDYvexaRwS0
ZDiN3iU7nF18wEvBtqrg8hlUPAn6qa6+ZBMngLx3cUG8q3VT4+7kCXYJU3qh6RwW
Pqi0OUhfOgJ6vDsKWMBg9shpOAYIg8WI6xEjsrkwkU9VhJpPAnxyGqCO1FKHA7b1
3NQPWt38AZM/D5VTTduKUrXDTujC2ofJMClZEVfBd14ez2GLWov0OiB6z4hjdqRt
VtscfWXu65m0v1ihxkft+REtuPg8Aa/iuNNANLOeq+n0lF0j4fc0VgQWF0o6kGgd
UdA1rrqHyU0/LVFhYSrGhXmTBLGfs709dpR+7x369221zwsiA6zmo+B57I6/KTnd
1X9nclN/PqvHa0NT8rCoFCVNKPJeaUMCH55U01/dghw7OF1IooY3c6FsKGz1X/aW
fadxSlyC7c9BczhmVLKTmgmabHggUSi8seoobdVRZx4mMoV6vbJUgw7KHptoLcX/
n6bykHUHAGgeQ7csdpYOpxZS54v4hzSUnHHXrhwZF1dLASO1oL52/VWaCIv8UoJV
iR02/Kkmj5YcHlq6IdnI1qh6x5AjfLMOSvtNbc22KVcD6YaeTLojvBNlgnxbTBBE
BSFuvemHdCUo9d6CneHlRsnMMyzgkpKb9otEMK7xJ59+PdlPxbso4//dPjAUrHhv
QkcMuCjDt7/vNMCqdsnc6PGLQjJD+aalTuIpbkuOD0oJifmXbc20xtCgMEH+N5MZ
7P173lwYCO3CzE0H6v5Da+4m9n9+g1OSWprwvo2kurVQ7gGiT98GEghxhZaueUjF
qbjuV+be7Ee68rB+qsIkTMiUo1gI0j7buyA6KR6TiMNUsKovfAu12OWk+46nWsCf
xKij1DWF0bbnr2FzDxFFIUwPXXPwzlaFOBLg2M/ZYR2EBNe20UZuorSEqfJ84HyC
nNY20rs88foL/hPqzgmOKUVhzThAFzOdfohgTXJ7KVflex9mBjjyFgu8d2k1yHpm
etQ4hZJSaC2c1u5p7kdlIWqNc95DdV3N5AzeKnZJsj+tAG2j+6/cq/4Vtn/q3QoW
fIvjEKtpcNXfnfY5iyfRs9/f02MWpu0FfpLCdNWarkOAXUGXeQfEG4JYDenpY+cL
JZ+m0npkEndm14Y3+5HiXkCDiYuuCM7PlEZJ6jAHWFip8LoBVVe9h70ujzeWgibZ
TgJXBUlilR+UfBiaS5S3XBFpPrd3Gx8V4HfII8eOpJOarZojQW44Rl1ayDtBeBjW
RASsc9IhxGa8Cxifa+HnxPH3E3QX+sAxaqFnAz8WP485CG+fzFyqG4T0c7ajIniK
c2qE5lln+Vq6BJKxZDUfW7JESlIPRoR1+az+oSL64qOBYdg2ngBHHIhmA/1Vvfpi
tbtkkIWcei3+XtCNz+BhbM2tzRoFSbKPcFoIKi8ZRWPeCvayEyFVMBnoPVAbsThe
Nw02Qvagynyy7FvNVqoDacrC8dy9ZOQnpw+Xs5lIHL6ZFALQBr1sIjZ007tSDO0e
Fsu9f1OcURFaHZmWIlzv+1FScnI3yBy40I6i/czQiYVYFp2YlKy/KWUCmFng2XrJ
7UvwydJaIt0stBam2hnOXB8f8zH5mAHCBw8ThgOG+oCtTiWbSerhwhbqvaNVhJbC
nZNlg5NY3GsIO0BCir16N47CN6W4ZbTiPCmIGH9x/2Rn1TUkm5aIBceZP8EBwHhH
osma/g+J+csdjcJMoLBNss1ay/FFW8HJoM365Qn6VSMvd40QiWjkhRQNNFNWfrhF
AfyMVgJ2Af99sZRn/A5dWs5ttMJba9rFvulU0qZNx0KhlDOjqUx06GDbH3nMnpoy
6mUUEDndXGH+L9sqEcxFM5lipKBOrAnU/T97xeL/sEbB4utxLjmk6TenOKn9EfPS
HTwApY1E0QemdyW8tGkyOrWXHrTtmsDxZHY1TnU58OWBvRX4Bf8aqTYzBmhpQDLv
BS9jNXUO3hGJT+K9ydXnZQZaM/qnRei+HLn0b+YfvIJurytWH43KQ5V7YpnbDBbV
0sT09XWcPjF7UcB/UrN0kH93VEnIsIrIvtJ+kdERZL1delZWTvKLlSmOZhDXLGgt
T8nb3lFFHkliyFybuwAvMYeZCjwZdllnCZ3wL5nLF7rt0UeE1g6t4q2G0obkgHg9
UWgWtG4oicTOrwrnxU1FA30AL51z42Dz0YXCoubSTVa7zdNWDYZ3KCoSQ44b3v9b
kf7UGvWf3WpG7RyAQr9xdnzic6v+EH8/Mq675gmljdGglysNMlGSl1Xqblk9s2Gk
dY4N4tg80aQD2Qw3ZHV1RIazR390vUuJGLMLOesTPrx82TdJWhK2Wbc02eufVyLy
OB3yOU8LSjU2V7SMs4WIBjNL67D+bY0TJc9Cgt+gdyeezespKTuSN0yYolza5Axq
VHf9Lj6rQC7Am/fnVS8k0007Fo839l7dVBlKCg89Pf1GFFcu5sUppFgtmjltDS3x
4zR1g8bVzjwJR7Bi3GlY3k1/T1jmy8/dEI6LMFcN5/m5rHdwwXMW0hZB20gjXb7Z
tz0xPaA+fprqQL3bvDWIUaSV4lkUUOAiTv8CGoB2YXg3iam50lcsB44Z25tn7KWv
VkUnd694io9ZYI1vwERvCw0uzvSixY52Qi+BwAOhFR6zNP/OQMYYFabP+Vt1s5a9
YpqH6+K0Q9ia1X9FESRk2bvVUyMQeUZRFU8D2w9A6iZ91MTsBbnn+mqmU1Uz8vUG
o9lblducJGxUlz/KXA3BoNuTsSzFGX1dnGs9AVz3AAqpFhtzrzyyPr1N2Cah66iK
0LUZcATuuO0YE/MkzUSATTtZ7k803kPyBQQu8D78RszOdJb9cdLc/aPQs6IL19/o
d1yecqPMH+PMPJGNYolWk8lMkVa4j2EnPB5jYZ1ZcBLgapdDB6XA48vOgT62tRP6
2gAHOsoHTgF0oQNNEIUPV+CYSRGjXboljNfHygEACXJrbZ62cRSRYUEbtqOYGDjc
tlfFXETHjy/mrFj3hf9vmtZVqxm24WZl5rnwPrnUMpSCuF8GSWoZeiDTnSJ+QZfP
Dfap3IdDrt8x8imOFv5JrGRIUVhF+KffMnAm/M41Hh/qU17zwZx54yEieg5l1eYD
BJTSBp1jS1SMXeq/UOc7+ZjBcxJJMDgDNH6nmZbm2r6dp6rziTsb0eS6/fKgJhWy
KiTxgte7q5hXICzZxEx5L13LP3Fhk6BRM3S1xCfG1BAVU9fHqOGX2+WJ9qlmtxg4
kEsd7Ak2ddC7jWuEnVp7pnrQnPPorC77+lMNzrz80scyRMqjl0v975EHK7EKgEH4
RnA1da+mwbzl6X1Lx73fMmXDn5qUxou9g87ql+aK53EUIOsOrUgRqBrtt+rsrrbZ
u7yOZiaV5CWWBiVOKjvokHeP/B7LWoI7IbhIh3OHI6TuwPA5ClS0TgCdK9VYvCdd
pdmJqon30gTxrYAQb+jcbNAZpTI/iBT75C4G5PGgjyF4a6Q7I4f0vwTawEKhD+RS
gLiOcPCECBxCQf56ixafQjX1D7f1JlOMESu0L8Ll5HVLNRFF5ifGa9BtgJTctoYh
MeSNbirao7Q1cF5jaGRNY51R2QxvN/KNRx5KAURog4jnvy8V5umzKJzTGhkGqsSE
PMl45oPmE3FabJHo+gCxF/+rZPHxl/C5WKrNZGul5vG4eF13kGBPxDtEzutgG3Oj
IOKca3lyh8qJYDeiZRjFz3EwnDyuaycHCHeiPu5RS2sULG+rPgijYNp5l1W81ZTv
HDxsgOgLWC5psAe+Ipqsyte+7D9EikGPQbH143IkMlNIHbHYQT4YPdHQ2JwG1GBn
7YYBlZWotXMAQQanfgchXh93Bv5oOXYVqzLDQMzJg+UP4bA2VsqP5PJfe0o1+lBQ
RTrgNqRGr3MUNe1rggcM/ax3P8G6ugRQL3YxHx+kBmOgl9Uz1LS1cJd71sqVVhK0
XWFS0wCM4LdZNAsvAcRBrhQbp2YD+T9SPB1bEnjLe7O7ojFWDL0nyx9WBrQ46EaK
crXJLtPd9Bs1C9N6FbQvi8pKv827x7KHnx4EiDBPPgKM3RDP5RrTNVkDV7C57Ihw
`protect END_PROTECTED
