`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZOSLPrh9hsDzLv/Dox3UP721D9624fsOwQcto+CdrsZggkkbUNzVa4KkfCBojvr
9oa/UtNxeXrOBUMkme0ZJNhp8vzKuRyNXTQ3fagUrBqcRohQ5L/x84WeXxrviwaL
tPaoZvyP6a1CNC2sMmfw1WbtutMBuUzVr2q+9B33HkAaERdt/CfALjXIIDphj6pD
VnVrQdqGUBadMCCuE+aLPOaTXymyG25hBrxYVNCtxjLsohboh5rrQ6hiCemOP7rB
bExVNrIPMIKVfkGjmLeSI8v2XPfaY5tawxXXblHfUsQUMD+wSYGqzFZdwTLr5CTa
hTQ4otZ9txAU8vdPV+ZsoPQRimjrDE8elGskVZO9LDfjMB1aca47vy3r6b7TvECO
GxfwA+k7R17z2T/MjJnhV6scLMvdDzfkEpFS9rknnQZY2AbcNuavjhZuDQDQqxMb
t6PZ6YcQscb0Qm710tKycImCQBW0cSXJQFIiAdcTZ+Jh58FbSNUS3Nk6U9u8LBE3
`protect END_PROTECTED
