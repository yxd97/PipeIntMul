`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jfN0VcGs5IlYssn1lO6KbnwBX6p3EMKa3WjASeoxtPZlPagYqBLy1uPULOxG/FAS
8xNTIcLqRb1USCnngw/DmxIqt/cpIaTU2HnJfQbVGRn0/Sj6G+dYmPRqyj6xCHgZ
fqM0fP9kvK4qA99+Wf7bePmbDd+ArTvFjlqGPaUS/pLrdpDrgNU0FjLiJFNbZVU9
XFK64aD5GyXstDkq0Up1ZVRZOymJdxDe3snxTxj1lvKSUxfnZ2RbZmK+y8QoiNaW
OPJEzuulxgftn+xDSjZ9Mf9J2yyRv0dwCUaKtKAEAdSQXckIDqd/eSnO6zchxVrT
XzdzNRA5lmVg8o5ZO41uLLGWG+5WRiYdIwuHyQMNsLvcXXKJoSwcOrQH+IQgmKh1
c2/nlvbBIMlKmANjelFLBs7D7uqJw/pisiUYUUj9hiMLPURq9PmVEojOqvX3d3ZS
eq7wcJruSA+WTlxSHOxLCp5EWE9T0QU98K7wrgmis1on9uCbgBSm2Fj6rP9Io6mJ
q/3gekBixmIILyCjbOaRtOjUckZgNOIDVl20P6kCIWk25KxhYMU1l1HYggc70wb6
f73jiWh53ADUblAc5kW5ZTNdil6B6Evn0ebQvpyA+QBO0hkea/JyxyTnF2JdsGFR
2AhSuK9huAnjJ7QwRyJFL1yjdGoTXtkS4CHVVevqA4c=
`protect END_PROTECTED
