`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11ZNL9Cs5HfFe5WSE8SxJXLku4E924bBgurxjBPzJWPmFrWDQOoaeBxWG5scfxtt
kowXQEMF4OyUwyQOIYcXodUJ8B2O17O/JRzw8OzBqXvOHWbqQEslRUSYPQU+sOHm
fbvcplr/gq5T/eWpBF0BVpOwfdcrWYTKJQiDK2A6RF7rT3r7uijmIoljvL3+EBl+
THbbfp0ALbfDQGhJbb9McweIeOVN0uPbDgxkhsJGNiuJsD2KyJhKBsJDGG8swcKh
pRmlnmTcro51V3kwPMwo35B8yMxqPEnL5AwXTvq8UGHvGMlHTo7UlNOKI3XBmgb2
5GK7+XiW8tUXr/NHFCxuxjuD5R+cFTrIORAMmcqLjSsSp6PqbCOWF+BLOfMpzRB+
h66WkWRgWmZtvU6kqEamvL+0YfPA3UpJeY5NEhZCQF5AVM72o6s1hjfbWb3K0qha
jGXdga1XKwRLGMprhxR/VycLUfnB9sRRNg8xuKgwJl9+WOSRNkrvm3H8C+kL1axm
nwsCRo8CkYUeBQu4pXltjzDWQJu6cKNoU8ckCKdnC0BCQozR33nAgHc2a6HC9DgK
vTfDXrDQxkpN2NVzdUxfHQ==
`protect END_PROTECTED
