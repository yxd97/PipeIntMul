`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ibQcoQF62vnVNxpUOzmIE+Y8WUCh5oQs8gk1sfewHBKSs2nb0bO0g5j8CrxB7kak
hrPOkFj95fvCVMuAIZuNg7RByX33o4MLp9MLYu/nL46lH3L1rOl29FW6Nwgy4w9U
SRaymVji5qtLvtdgBX4JyH6Cq+fTMeMi/sFlvoQYWTkA/wNFlvOn/j1KJnbS3f9r
y/KFVcWKh+YKAGkF2IpeNB9HKyRdqv84VHfr8IJONsx2bpp9gZ/u7fbRFiDoiFo+
amDhrpST+wv5QPQunq32qzlJdJkayucnBbThxAPi3J+2x+SX4vQLU7c5yg5niS2E
hVRRksZI7kqP+ECkS1FBmx+A/WVxV6gVMNULQOPHj9Mrfp2p1d2Dcrsfi+yhqW3Y
YbNqjxNCTflUs6/jVaIc4Te65v9DZvP9/qRVWmyORGxHAr1I3doQejgTEIfCdH6Q
AIpFu/EJMgaM9bfN0yFum9EhAZb2bO+01PIESQmYN3hGUyEArOCXyaUoocaxUQ4m
4D2yD+iJlh0nJ1QFZMsxrBal+mrcjZQayP8dV+ODe7K7gL8HNmw4EkyEKT6GCT/R
xQxPVUMhIHk+ZJAnvyonvf0NnSEFpad80xrggnlYkEFhVG1JrSVqk1EEtSJCZwRQ
hCcfCnQsSXo5OlMQ7WUHCliC7qKFWNH1/LwIzx9eSRUTo2yfi0+8CegHVzv4uHcC
TxvfBnZYtkts2pjP3LoJaAhhpFzDK2f4dKPHQFV58H+0cGpOncAhjdE9mayWKt0/
cU6ItrTlQmGutwKS4vJTrahrjfThb3Q2jceKSNG5ecT0E9SFmgXgjntHEdPLgPB8
No5iOFRZXksIzgIpdKY9Nc21prEHutNZMXqKn74htE3S7yNJ/Q9lDqzmuU2PkGvV
vP1a8zXp4fLQgKtvDIrMcNrIiACJv4nsbueh3DTs1GJfvuO04M1evTX0TYgYuIoD
0cVToux2CbY7OkS3M571+Ru7UCK5Z0AcgK2XXdkmsW6FbILKFJkjBV4NY4cj9Wev
7+//zi+PJt+0C1DsQQwA8Mw35LkCgLYCrLaUVhS5Kic5oejBSXYDanM0nCOOKaGj
PPXBFquLf/ZtLMXlc/o38LcW6hRpgU357UwFFsr0n6NdEnaScjQoRxmMbuk21LIu
pxb4q++IzZpG6mL6XebUKSCJ5K/0Yq5FKunjtIfBiL3OcViXExc4+kay/wgNVxUN
FYLEMpyo6Lv4ty1mtjcT0uMrLrEF76n/LKC9Gz5xpE6UeNHejazsTbHa6ztH1Kod
AeOuOPu5Y0b77Vf+s7Zf2voY+WBK2MSXfR9g0DnDlbc2Tp40DO2xLG4KMWwwHamg
dUJukq9Sb0yZKJDJa8JZRYTl8AXxLXrbJyYW0P7wN/fbBt52TsHbxR/F1UOc1Ku+
nzPQNTtPkFYG8eQWP2Bkmfu5tWCib/9pFhuTyB+ilcP/ai8IpWqN0hX8s2+g8t93
4re78/EuNZJ26neEl3Wuua6owBS3qJ6rSxxYRrkb1vGbMkN0U/UT58VAGu6apJWP
I7E11tXkEDpTRAcInmdkcueNrMdXFuWU5G93qFHq5NcOXH3vhMe0XoFQaFW39VHE
U/nmr4bXc0ijppjgxrfP1+CsEUVKC8M2yJ+wBSpYXQiBJH/PJU1tyoJUzPyOr3CB
KdiDdaLhw42M4HplIuaTaD23jeGk2lkIf/g0xBOSulbHDu7GIN8AFRiq8Bx0+MJe
yoZ2YR0PMYmmP/rbI+tiSsUUIRiEaE9JQsJJo6akmbi/oRN9pOoRSDh8C8XNSOty
DSeaXzKdCi9uRvTaAujMOIqQv9+KlTEQjSR5sf3lNiZXGM7DqBFc6lZX/idVO+PD
NzvSXuWRk3aswc9RgSXcFsgZum5FxJwDBjgbj25pec+k76NLqCuebqnd+gNqrfe2
JnEvEM/VZ1gBkyrS9gbs6KdUagyssq04o7USZn3BtKyw+GhwqjRL8HITDLJqkOM9
D8aeZfXHQx+bgSFideU1vlm68jR49/mgWD9Zi4Q2hwWMXpWdef+HRA7Zl1XNsbET
6xmrLmNpWejMKh1xqMsYXx6SwgdbfgPEoJHwMOFRuJLpr+CWIx0Ou5cKLrfYF3dK
g1RelMAus3rAq2qyTPhE+toj49CG01xVJ7JPM/HKiCH8yYmTctZo6Mx+gnR2h+oe
W2B04ERRzop9TySpIUHAOqS8fuWXymC1sCeMUmoGMRM2ARtgBqOaxAqvGWZzElgF
ZzkL1EzIoiIVaiDwMUiQY0d77tvrVLXt/jtu5JqIYWHFE+2clHa6kSx7vJX/OAAj
LplGxFSkaXZ5qOob/uhio9Nzh2Yf9Gbl5qiPYn3/Vbq8qP6pz6Pj4HK/hVfMtzgh
y8x5YtPoeKZmUiC/GO3RIJuYNqByS911ITLyqMyo6vtCbGSm3ud1NgkJDHvfJcnC
`protect END_PROTECTED
