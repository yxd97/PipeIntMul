`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QW9E3t6Zu0c1P9gpk3bRVzJ1k68gsPpZ+vVFQNdfozqxpCU9MK7TlS0WBD5/PsUQ
MIlhjlgeNWka5CqZv6mFpqj+n8RKR8F9ibYOBvueuyFFU1BeMuRkeOXglAnMxZgU
DIvqLaL2PEw2MxiS1tJBDyPSCRY4vhHjNjLlBwbg2irRC4Gk5ZBp04cmgKEXqGkQ
LyJWV8RWFP0f9a21bU7TSi6auKmZOjModwkgiC0Qz2m3HsYt9z2FP5TjwPz7u0I0
y13vFxXnzR9VQbflRv/HvMzVjHplFUbssCG19bSVDglUbrgUF4G/m0kPNIWNGne6
UxwBUdD8PT2sOEDbD7vOKVCHXod3u+k3cpS4MiMVKeUMiySXamggW2BdWdRytJh8
a87/2h0ohh13n4lWDJNZVPOXTlWnc2B+P6PzgS1ulWu9aTA3uMcIgGsSunkjz+CF
p7WPv37UlZ77Dlq7mabP3DsdRU7+1opxjVuDQRm8RhhZfsz3Yrga1WDzCTgIQwcf
jlu7zY11Y8QkJvGySUhD7O2IokZM9dpI1EHvTG0/DQ63EWQbLufNHumZSA6GH/4y
9La5YRkraX8xfA4vsu57fcN49+ZhyP/ZjfZPog9JesFa2N0HXtdqoFe4Df4lNTf9
hG7y1k20C6vpXeM6nFhJjE/UBMriKb+eT10vOtgC/7Qb4ss8QDvrgE1Y/1HmsZVi
YgkYdDcOUIvVJl7cQbdbAls7iqN8isnNKWXgaOBP1NHD9rqGTNtoLaYQlz9eiSmN
DMx2kiaezoWFsEerSstE0Q==
`protect END_PROTECTED
