`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0xmiEogFVnIRaH2KuW2IRTKwmUGoCONEfOWoyH5hDmU6J2Mz+UiXTOXA4QfcSZQ2
t07SXYCIpCFLexxiAu8PkjO3AA/2RodRyoW63Sr+rtuj003Nnnep5hfadAlMBoU+
nlQd3KYV1ewO2/r3aYsMeRMnM/CdNeZPS8sJ8PkD6y3xQ7r6AXvsyf1Q1fEfNQPB
L5adN5NnGs2MH1aKzoEhAJIbWjFlEK6R+0uJZIi+pP/dtm8KW1RawSlXaOcoOACI
qk+du7ELtKlBSfTq8tK8iF02Q/MKSg3actuMeuU7iJjGXxWdTpFGZeE/Qi7a37ml
fal4439AZMErcqEOZoFetNbfrzn4l5PG22UxoXRF/uJS/jaiYikQiMCoRDVnYKEa
aWMzQkULvRjebavtLCNN0xaZOB8lMfvIC0tbaOlFDV3CDCtdZhTol0RvAICQLCka
BAQ/Ffi7Eus1+5SyZEt6Zz43ggV4Wrpn31EMHz7sP+skBHaE5i7DgflHcT6DhiF0
wh/q5WGI/i5rSuKVTS5L4RUJBmaxtuXrjf8eVGDgWrmxK+MxAdJo4P4T+yauH86d
qqUWTYP2oqW8h0f9cRpdXN9/CnhW2LyzgLIsy1uUL+Mztkz/TZX8K4Zejs5D6PDX
s0L+w0Orejnf1rT8zJ31MAKkjpMtnNmW2wDpALHYza5P/eGKRq80IPg8GICdClw/
OJ+Reizou+6s0Nc2dajbXCQaCRvq3eN2WHljl+Xo+Y9MAWZZVBGQFhh9zihoxrtS
Cb6LjlyfLzZqzAHQVSRHQ58WJ5kTosANgOEFejqAOE+nshTva/UR2vcDcteGuLh2
GvltUsVOY3BPKPYNmQQlTUTlnMSwnOTJzkcUPmSJbTMZda2Cdbxt6TP9VvcK7bsy
kXDnBNmGDIuZpMHihjSr/hngmg/5qHz7mZbbRTV2vhI=
`protect END_PROTECTED
