`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33QLOw5IeNwLPJvBJR+WKY74ahCocD5PVuLcL49hF8Nrjg+PUVvqDaEDO1he2AhQ
aJkVfGndNjj7Nm8KHD11VjULhIiWxN0sV2xpeI15dbo4ITgSBrt/qfh1ZdKnDGmS
K6Rcae2biL7LGaDwxgjZvY3T+w8pQWGgos1gWobz7f4ql6B4XURIbZjaf2sJzncB
KGQD6JpEFn6pUZ2R+0C8WKTMJNqGdD+6pNjbwC7LFiLNxnSuPdL3a2XBUaQywZJB
IVKgo6mYZHChJ0kYPxtA2xYAWup+cqJpiVQlumCwQfW/Xi+S4CyrOMqVyFrKjwAg
+Os58yN3ltHLCzxTCwQqx+HaHsnuAgTqkOkx8heb/zoeatYGwcxhSIfJNqbEaM9A
g+DkAn8qP6lW/QAMTF9ioI/3XTuZy5XfslUahE72pE4G0FzlCZBXyNjm64vSybGv
4RGH3G0Dzsc1TXHxnx4B57ndQQsrR4AhfXAqP1zkx8CCsNv5vXGTOUqNn1xjGmmD
+0QraZtaA+tCPDX4+Zn3aiEagyGsKMgBR1u+zsTstlfl8QiuYDbJLZB8l8SeWIZV
B8/TwUv7r5FhU+InwmOtGkaPMJtnxdgZd8NJOnwBZ6ZM7QDvkpHd/MIb1zAr1qWK
p303yhUBmNwRB9w3PuvbF3xdJAtF7Dv2zsHXTm8ZuRkZaXPkylK+lKnNcG8CMRAS
muAtLKpdy6tlwtz3sQhqhip6QWjf3oA7tjlzX9M/c69HSeUxH8bFuhQu4g8aSt5M
FvUyCMJ8ynntGTcoe2kwxautALlTHJ90CYBe1gO1X56xlZfrMCe6IcKjG0EWTuO3
Rrj3U/UFHli5eoshWv1dYt026THGsAOWHY/9ZbrzL1P3b6Xqc02ZfQDzwKRO/lJr
PbYOfOYkXSnJ16cID3FzZjW4mmAv2ZYQl59lcQSDKE2X8YDHmyGuw2zJbXXOtX2U
N/dAPUeemt0oeKslJWkjj8ky1qRY7g/r5VW3Zp+ocE8zhxgPU/fIhmpuN01+oA/4
AtTseSuQ00/ogGpg2GiHDXiJqGIjHGPXskayqhPdRYw70/okwe/CwrkdKp3FM/Vq
srVRobU1gsnb/qiQW0DPrw3nEa0/d9261KmHp89Cy2Gq5UFyKY2cgn3qj/0IUxYM
5QQBZggNvTIet0YKqznIvRsNA4tH212jvwmfwlwOKXUsSAzmNbXIvoD8AyZ4El7L
2slZWAJihgb8od7MzfJ0ezgEkr6LwGr57Ifn3HZCC2wn/uHCT/kmmHff3lo3dfVQ
ZtJy2STOjU/Vy1kdzig78GQ2f7u8GJ21Ehh7dhCkR8E9TkRrDgPE3mwrT3mWuAl8
3ml5Zi15Wd+bWQfPyitEdD3haZyH4jJ5hWyiYF8fSxMjoUS+j2upk3BogL4/JYk3
7kYPOb18+hjzslS8sRk8idMIJbMtVgqOx+gTnW3YdHbAh2Sh055w/4SQxrdQXkHS
d/uht8/GZyQbn8PGb16WdhUA6tBGKhgARoRvKQeVymUBRqVWJkw5PPMpwygTzEaU
qYNETrQjcSXsFSJm/S3V7U+QkMW1FUm7VWTLayHJpj6qDGnwzMMYWwaIa67AntDA
PwxjLiVz4q3OrzwMrRX8nEValiSL3iOyEbYcOI9OMfh7cLGQyv7hK4QGc9sAbfGC
7GFMVkZvmkS/vvqkybXrg0m8VlkkiEF99q59lN1WvPsVjyHVc4D4mhyiUxuB5OTt
JudtXHhz1q4ZHR4MmdDNJHhiPlVmxjQnr0FJ2KRcoK164nWaPLcCWnhuItrB2FpA
+9mkUja7A5hh6WuwrSu7Air+Lqp9CamOt8ZYuuvRTvUCU+ux7Ehvl8wC/ISERvgM
EbTrwI7L/J0lXwqc6OKCKXjtu4TsUTbnLk6EB/YvHn/rLKIMWlcYMvgkAgrDiR3t
3oUvpQ5wyjc5AicBFQImTcxYCvVA2uXDIpN1+xIfdis=
`protect END_PROTECTED
