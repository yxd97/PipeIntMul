`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjjHcAeG0m9Khmmr0Yxc+Exk1hf3e26a944IN+EZVyduhK35iYi+MGqzFTn124pB
QqDNWP9RiXXWsRjor3MqRndJ1Omn7a99i1kxPta8L5GLh//JF18g0EZhKtGKS1j0
jc2YiASl8WQNsXFd4zdy5mUUIHqRb8MXl5NOqoFdx2pCxr6BnB3C07jzFFA055UI
pj+keyErrC3dsS/XQkMdwTFkkHfTiVZL+szr7CZFS091JKBDBe3HJuyEUjathIeJ
8VtP9SQ1i354nkjEQ7ux538m+KgCmjVivByIZtMRfYN7TkXghTzJ6M7KFQqt+lSA
MSLQCOprodtakL31jZeE9XdpfwOVGQjQRHhy2i1huYKNJqdjKNpckVeTggN/TAdM
8q8PJyktZLu8lzKeCNluIOb4CE8ieKpgu72ej5T44J7Q2aP+uRJj2uZds79sfMvX
CW3eg05zPDdXJATlGwYfVNwWeHtrMBXF0se0yb/60scTKYQP4yP0rcXz3g95mcUP
07NzqDfJ1UWJxfcGGS9wdGJZMkxS7AYurh0hzn4xjngyY7Nv5x9GYIAj8sawUl6b
1BbpJ6TxHqIeq2w7Vl0/G68FJi8lUsaHxX6WnW5kjnnC0iEDnOnpImxwThAVoFDs
59f/SC/0tAJK2UbfOOZaX1AQ3qDCmXxsOZB87j1N6X841rc7jBmMZubxNs76LAzF
lcs6wXRtnszmclLj3tSu+4J98YlPSQh7r32Ev2IorEaGKEnFAs3/RligjhCKcwwm
gRguq8kqBoewfNtRHRDqIIOFkmCuHq3vcW0VE0wjDqXJoeBHc1i93AyoGbAnrfHm
h8AisFD2CozyJMIK3r21pYDXr1Q2A39dBHMy8H6FT/0iuWjLqYojT2K6VX9HK2Wa
dcvHozam+cAn3bC9Xl8BDa3uXM/+WYd4+iJ4QCBo+SzUG2lN7NwPTS4Im4jPvTFQ
4uqOMUcZKW4Jpr/yagwp0cPsw2VCJCWKyRaDrsg1Pfa5DcJbnoWqp8IIJAe2rUTS
uBL1KErkKeAVqc36aAl5fDxubITwdodYGefeLqYVj/zdzO+Igv6Z2iVEvzJLLuWU
KqRjQY3jjnqvs7yeDGl3GJHpSKe5BotpmHvonjVZMfZStyX5KnQo/pk2e39y8jIl
Ko7ROvg5+h2vZAhUT370OnRJq18M9SgKSmVBvQvOralqZpdNvHfAgISk0OCBZjbc
+jX9vDVE8V/WeoMLxBpf6MVjAQ4GOkRHbXkC9LJHJzKmc7oTm2WDAByoiqpWcXef
j4UTQd/WnLrz3CJg22vyhZba4LtbgsAekqi6zYQZ2Kuvpl4MNoCUOeeOVSqABl2k
yJ3mqy6Rz9JP8bSYmELwiKq4ZuOLlAx72jYXuM55o+6OlpYIIwavyktasqztS0Do
1DpuGywUGhzU6nVZoeVyAMDOzzzrYcMr0H7uJPA59qnnegHmVKyjdwBmbuKGUIUS
bmwSvJILpy8XBZOL78VBjwMuVdFWRHhvPfrPsPS9NSpHiCVqpBUM7zCoGu0IKGot
6fbzUlpP188vf22SUzKQAHWEw8us28mcw+sIM8oOefkm8y/5YVo/+Er6bpzejtHu
1vKaocXHQdZ8qVSyshFF5IVlQ1od8+1Bzq3Wx3/DWK8zqwV62prEp6Zb6oo5I0wp
8m1CIVkDgEdzwoipyrSOwZsfFya9/Nw8PUrQVAbKtfX5DX28w6Isk2VgeFBMKsOs
y38teLQuCYH7EQtHSHGA27zi34wwpao7du9PPxVM7QTJAv4BEIbm6V4iJT/ALXuT
VskJvWMoBbGYXXVRUiljDCIWmgRCysgdJQQ1g+MQ1/pCStwG+XvIUJwYThRXdwzD
uyb8JM5/Um+qqZKgtPrTbw==
`protect END_PROTECTED
